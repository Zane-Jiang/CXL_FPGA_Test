// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uosQ28ZWa8L6joQLUn1zOlhXpfeMrQtCVylKZvK8cSbBoeX0thlH2E2ntjmB
fUnMEYTGPNj/0fOuWBfWrKRrgqwDTWwEf2zZpM/B5Birh/bOJwtVivrY6jy6
UFeVA+sr4DbLiEdNkMPch7p8lv7vUbCmI2nbj7Kaj+xqDExh6HqadiS0EA69
BkdBZT/J9KY627ku2u71QRkKnlRX3vUMuwJOjrLGUdpHu3NLBBr4GHcqXDOa
x6gSPEMPE2H91UNDBLU2xwgPsXZUH0Rq7R1wmCNMhVBd2NxsXMcuGNdDmpfL
JZXZ73RYzsoKNOnrJeuUXFDhrvC6xnY1ZyCw9vmbRw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YD8anBVW0za74JTFw7PiU2L5YW+nNqwzEzUaL7zXHVZhon6kaR2QCyRf9Z6i
gmCOOErDSbRvvk1wRbsgQaFPSmdOfxbGSZmE0KTfTTuOUwvYLalRUl73K5p/
3s5S+J6a5DPomdCZkb9OGKIwTXN+iqJPZcwy37/7Z+09+W+Z+Y1sf9hG5687
ElgvXQEw68DN58FkoLsP+MfAEHu+TCrNALSZX3aloYAY2V9aBS5JnHp0ppaC
gLpliThHYLDf679IuVws5Pmz/7XZ9MknEWW+ocpBiErIfuEs6+gEee7/Z/E6
dyU6EebT/Mw339E5CB/ysrGLJ6GQT6IiovySo6Zn3Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ncMNDbqOTY1hkD0c+tIO2gvZUH2G8dm4KhR5iFwsQHrl//n08PJdPWkU1C7a
IyrXJKcwLVfddD/984whKHrfoqwdHveZAEBJ4lm2FASUMpJbP8q90hI3qWqB
yTX9p4SUxVHSDgIue4Y2VoIyNRJ/npJ23uxbKyl7MP3ws7t0wtNwPhnI54ud
hxO2YPoJXxEQ9FI42VAGblJ2zKSAuBko0I2ZbwkprO+Wbg1fGOn0iHsLdZml
mX1G8XTPiBbRlQAXym/9inhIzb0XPmLCciO6zAUU8sCzBlR+fI5h22tojpj3
NWRhXmURkuVQAR3SxO4QiJYiTyfl1J8JXE6Gbt0pmA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kcnYRU2xr21Sk2CWRFtOkas6WA0NAKTbLNiQXDZWZ4VXunjy4DKN0kG3fvlx
G6uzImg93C2qy72ZEOllqrFETglPPjjI+tj4cB6HbKns3xTL9oqqSwSEF/+d
G1qEY5AlxW7gRMVy4U5H4rxNT6j/HofB6Dt8pDl8Z2veTnXgR/Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
X6iapQagooD6tX6Xkj3yH+5mNsP5N+Q54iqJlsZw6iTPSwKLcDPB3LJ6i9pl
LlyOt5FSwyeaxDXCpiX+CpN/BXqoGol7QvlC5N9x+g+yflqzy3s+PXkJW0Vy
rgIe/Oq1C7+vN3OxyLzH9siNwixpEW9nnYyFs7vVapzsxpSN7fSIOhlZitVI
EP7k6ytW1k8eBvXNHjeYkUDJh3xNLRJhxWSeTpK7N03p3fKkSU2G+49Ri1qx
pnacu6321ZBjZ2ilU7YQaJ0pxdGsq9GsQt8Ydcq0qatJ8u2HYXB/0Itre+uJ
XDU0TWmysyQxWwSRkBdcyGsSjoYdgjocVgwQEOWlHtiUYWhtcLz/ALqDiuD3
fLJEVMqgyuVquXlLUUczkjEFNcztG0r34x4IDtDP9VVyzZLQBaeLAz9atTTk
qPU2qq4mYtpNfIlLwnrW9IEQW1G15Ub/LDc56Ct5MkHUe4JDeQSImIOPl91Z
eMMmKRFYjJfuvRMLGXWz+dhxnHsBgRQE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CVgqMfk4GANERmOIKRA4LtL3rNcWjuefDwx2Ho6t8yaXK1Tkz7jJxNCZrKFC
RqgUtjvC8tCP6f4Yjvx8XexWJLCUW0u064z1KvfgSQHvl8m2Wm1HBI2mkwmh
Boi9UA0Ss8Lit0OceAYq6mtLESWoMKmvQmLLFPaZGxbc7DitY1Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tqKIUor1W5A5LycT3F8JnfCqf4RsQh+h88QvK9hk9DqBCdOD1nsWdaHdE//S
WSE9nTtVeNPz+Sbyqnzm3xw8LUXebjpgSjYAZImunNr+Z5OlXcn+8hc9Lo4R
TDSG99NLugLoX1BcEpvKvrnmp/u5ZaLB5mW/jPcfnEIsdRtTMF0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 536976)
`pragma protect data_block
ND+jcPwRZCUsoptF/WjkOe2DEeok3Xsy5dxbTuRAKPTnpLSORJp6u0V8UYs7
ZP0gLpU0X4XROMe3Ev+fiZSK1PFK+yTjDHEHUgXYTy8s+U3qpj43Om78IrPd
EynEB3mHNcmnCUOPO2Ut5gcKtFXQidHfXDh3chNN9YZd7f5xGDf9DT8Scfyj
OcIs6Vqd2aDqB5gRQjM8lg6ebq+h3wvtUl0iMzNlRpe6+Pvxo/yHheMyhyzy
j1HzhB+csTUptMVOcstSfiZgfVELhz+IfAwpeP8bXFaMpTJVslMa1su0d1Yi
r9j5GGB1wh5mnoN1QCe4Cs+e8UxWekV4+TFOqfsOwv4P5kdyij8j4MTQPgZI
U5nF7IXSe/qFHwop819fzoUV3J4yy2GT9WvTvskAT/TBxhjgfofwsL7kWASV
TPa9HqRBvKhIwA8W54ECee84coQfv88M44a1Hcd504hZGnKN6GTlPT9DTi8W
kR/+HyOKbNZSLOvP+0XcAKJfPC1UQAtCjfoeMYAouIZ8v3kVyMRnhcRTqd+M
ouClOXcm1o1j+qPDhuIG38Byzhv42XEbV5AxYfc9+yl+vMKdodenQZ3jaF4U
5/2vszuHJUIfD4gX8ZPOqjZYJK7NIl+31Cb3U1T76aOKZuZZIJzEpY+8CA2w
aiFsK5ZHQUkftFeJUNdHe7fO0DWNTgw8lrtC3+6T2s43cdEjYwHMIpCKktVO
8DxHLg/2AEDS9sik92kuhP21SKWS9rCfa+fw1PwxY/4sQTZLiA9Jxh0sXmyh
Cg5IGgZ5tZdOUm8yDhrM9ZTynZ/v/8o4whkJYzkTPk7kEL7TnTkjY5/xSF6y
9+z6AUrdO6fmdH8nNelQTBkLLoFyj54qQc/Kjm2uR5WioihtZXBAbLl2uDmf
cWeLnxcTOhyRF0YfObRULGx9+xh+zf2r4puV/yfcXL5AF+pNp3uZomzmCt5S
Y1zakYFQ57PpxjaFt2WJsvYqnjQt3Q3L5m+Zqlg7HkODOBQi0w4bKrqx6mDw
SNr5IY384nLkKGyVjTtfgty1yozVVhrHfpW6v4+A0477uq5CiOEVvPAqurIN
7kfpYIrIOtGJNpBh+lGEDtAoj6QDV04ebANj5kgvW/tTwjwTH/x4wJDJwWH3
gY+Tu+A0YPuxnZZXSbSrloCSvvcVWJhElo/1gbi4+aFqfDG03Tr4/ELRbXhu
cxnb1odXTYxR3eMA7cbjlv6E4jt97EyInDxvzt5Jgu0nt+NLFS44ouMo2oy1
JeL/H3dkq40iBwcRnumNnpx0X12ITvctFMQXBjyAyp/yof1Ri2MTvHNonx8D
9JdC5d6+lOUx1zezkSK+9Zdg6ah63krEcEKAHEYGdFs863IpQHKr59Uo2hlj
CMEwmmPkDyrenjI9WrkTJImFMA1OkYxsG2O/nkNH3vaWzc9zlrcmH84qWUlu
BpVUrd8EGAZjCIDqHxjB/kJs9iOMJ7dgYIbS7vh5X9KxetRmvpShvvrPDs1x
78WCy6pTRv/Q22WLk0EoR6pF6w94lfJnqY6OzdQRyarS8blOewxabui1/NTT
nu3yPsM9s2jhLR03zFttuwfvNR6812dY/V7FVsbGZjssrmhK14hyC6z7W7UG
/MzkEu9SabwkgZuLpj7WO6GAyktPhB/XGyyDnbG55rlYZy68s+3vGIPvDpzV
5nMWcVJw2hcTyv2pmlUlUdbirjsW78ESEKOP8+fyxqNel/0oeCo5dY37d/Xu
PYhy80Ql+6LuZP+1nb+h8gurjxJkZ18gyzrNamrH4MQz5uKehEmEcJF0jcbh
LwlpPGC9GE0YHUeqS7Fpc3gs/17k3c4IIIeOqVbfW8UhjpC5OIx6m6uI660J
2pN0A9rIa1svhfC31YVJ/bH3mpMCcvhNPjSxoGPWYi/ff10Ab9VGNxn4evX5
cwHHSic7H8f8BZWFKmXYQY9B99dn34I88iu0GOZ5SAdRBL+MWE337gDFVYAZ
DCviHue08mGTTnOpfl5kdigA1uSuGKuwaN9iW4mMMiFy5X34j0/s4+EvJ76Y
fJpJHc7fPxBjDYixd9gytoZt3TQxp+4BRHlQzQK9JLh7mNraNqQgulhWT2T3
b1pfVzjazGRWI+CCM3f/6U1sNWKpzzAmNNngjqPROFCUTx2KSQuKgezZA/+z
1lNx2M6ILaQNrpko7sM0fLynHfxeAhqLRiXt1vPLDbk76KRgef7pVMaonrxA
PpEAP1MxlwVOAPG+n8QvUH3qVhhNn+QqMJoI0MuwNg7ESvsjTHivxO1PamEI
EZT9mCUeJRX8ZKdARa530HIy8M+YN6M8ugjBt3E199YiBjgbvCTioY6U66Nw
tTxrIn7x713kGu5pWbb8F79ERCB0d57AfLBttLvVc2BK2QL/zFRtMA0on713
WLjJgZWPWxTVA7lKpZg+B90SXM6VjHA2b4cW/hWNP3kIEq0ZuofIxZfqR/7s
1ZSE19ERvymORapcDiVDZwlpO/rPhmQJoYjIzY9uhaFXcl5zz/AzCCg7bcdY
1SHBoTma+Uy7PrCiOkv2IsnygR5wrytFn/tCDt+ieoaBoi87EPhGF5JFRS1z
o/4aYOq4Imo0huB05E0ZdKYM2wHlftoFgmbOdhP55EqIGfrHVyvbJTql9ohh
DzzkJOAYXcvfrDx9Ym7OgOLT4LYuFdAdn44uM5YyPtZ9KVgj7wgakAHOa34v
u74Pa2xep/hjwruKEbqK1W2nAyH1zvSEzP3DzFpNQ6KGlrmBJN074o+7OZKK
axErKVKhU7vsasbWUKUm4xssyXZW5qH2YJNwDvFWIDKzZ+PUMYJ+8k+r9cf1
r+xC2PksAKSeCqOPK/U6B2AvajZWHRA+RQUq5jm99Ebh2wS/9hKdlLS9Vd+0
EkSPFwslMb3ylRqb/+Z37tKOfqpbAX6gzp/MqVj7P5hACwjIKjAeuaZNqmLd
+I4MJX2OzY4484RxI2ibsy1b1jQeAgYHEQp6lcirQcYa2Gxh4klLeCNAuzUw
5LnAAifQ95JYfd85TcXIsh9KkiwxsIAFadfH8R3Ivw4PirUgOKwxCua3knYq
UTmUjw44DTNhBs9ExUu18byNz9JtsqZsc/hwzlnKlvKGv6VmRpOPYFt++7Sh
P+mRPL658nOjUj7HHOROR/zJu2ktUTaZG+rxH2ORIWUc3vKpm2RMKy41WTR1
SeUb3G0upUCC8Mv5Js5F+guyJufb5zELHxHHUg4BIVb1hnsrapwDppwi7glV
3vfs3K18wrA0bWxYv0WOularC6OGtFJIrCWeuCLVcS0TzrxUuj01tsQAOxfX
YtqRxvraAt4EaKiEuA/Pm7xTWKNFMzONrjyQ3evbk+8oAPH5LTNbghd/XmRg
nfDbIkwwXoTteTIw+z/h5LOllwsNE5eLRn2hf+3p1k3bJCnTKtE5HM7i1DFi
PsGJcWR9tiYQDN8CfoWgDaQV0sT2ApyRvj56yGNkkzd+P9Ls14TT+1LKs9a5
KpydWNcec0VoYhuyFc9qCO6rR2RPFxEAcXhh4WMr9tk4gs617QJiyy8ck4gt
vP8m15KvuVSj8YZLULDoWd+0xggGdFMNJ07CCfhG23rAl3Nafn6r4eA3kxBN
K2yI3lM8CQ9FYwYJvdVecePPAEzO5XTkcbkBZ+y8A4PXR1dRvUZ2lfLBrzA6
QuVN0ZVD7aKbnjSd/PGu8s3fCqeU0D2V+R3+dIuICvAZsiRAwNsrNA+zZQ8g
X7WQcFLmZUMmOPLenPVG1ItwYkzjtcmXgTc9z2JnBXCva/HV4nalK+fGaFEc
bKRnqeXpEFBC9niSiRuXup2Vtwgo9iEZAko9/fMWSo9l0PgIzbox6rLiQzCz
C1uEamQT3wT+hnsR/V6nbQlkCvQ97wbdbV1ZFMlwYICguAjZ4sL7L/9kqnEa
UHwBpMerhJkGqYpTa/100CCwzHxlJrGQkf3dNW9xOx8iGqDWpfLKpjzYcbeE
YCCwOUtJsGsAFclj9l46SYMfGXWMgI6LloCsc5BuqJ/FOuoMQPhWJ176/HGS
PYur5e+shY9ruT+LQyeJCgr4QdB5G7vMOEqf6Y20i7gS+7q+3AzTMVcDEqLg
sCdJhSnQkchwoiLvfinBznze8Xy0qOnn/HlCG+VcwE/C8LmRpUfhj5GY0sry
VJNcowVMA/fb0xgk8b+WrzcHbAYuVXLRmQIvmm1M/WBmyk/fh2WzdL0fLJbw
5v5ksUE0+WS8BFO87FKhMZGk9bvRL7XllnA3vbtcOA2W/wIuXf7aH/TlCWIZ
kH1KhzQeHN80EXR1Xw/dCu/8cQxmWPTpjEx9hdYQADAro5LuDxtdiGuFOIIh
dsZoCkrywXY/bt1WksC8GltRfKasK70RI5Xjy6mqcVUhTm4gXCmMEZ9/R4M1
0baJAcolqoD8oZZVjqXZtM1qED2ag0E6z7NQFj1dS/z5azFyGUXtADqxsHco
dchl6QTrO6Po1maqUyC5uRpXDdVwUPnGnwheAvxhq0rNddcfesynBGfXOkmZ
LRXYATBwJpBaj/H3Yoq20CQsijWWX0TaSWAVMi17feJaCAkB5Bn0znhYONt5
0t4oAWDonxT7qdN0WhhdZx4poD2mKSRKjLFNiVYgG054BBtysxFV98nRE8yI
PzytSPY1nHPI7FZ4jEA4ynixdmtd+dg1ds+y7KnhBhuwZ8g1TaeMSUDHS5Vb
LUX464/yGrfOICuwyLeHGSjaFUecvlr+okwfl3rAn/vaTzrvHp/t/YFCkpBR
ICAnK/L8pU+6BW3Bc/giZ2BBsToT0wonDUHZ8VKDM0hMEAjsJIDUqIHN2CYA
Z4ZOYtjs9Z1V0NIoaMVEpsk2xY5LUJHabIe2EQ6lUWu9KtXfn3g/dHGCepuI
9R2BT4NSueVKKY1iHknQrWGYGmsrgDFeFI6F4kdSlqTy7peolENClMYVlrLK
Ua6M2Sun2I9TFWubd9INUO5sFB2k22bhiby+uXY2OcykSyPQe9l12CyfFdwu
15jBUF2nIj1XPgTesR0n1fM1WgrF7bZr1xIDJGRQm14pg+q+BhdnXA9v46R9
uqbxbfqNvQGU+nu+On3n6uKQnyO0EWCm/GMbYnVY1M9mHpkV+67uAXb/BYXF
YvbZX3Rqej7k6F5Vyf5nWlt1Iam3d7eUIxczg5S4ldpYrI1lOkKtKoyzP9qu
AEFXbrSB2b5VR9wkRdJLsTMnKqNI7BOzKBl/ON+QJVO8kdMj35/TeONiMmrF
Pm1SK0hiWSc50e0mokz0yQDYq8cRBbOQW2TqqmsvOiIeAyLuF2CllLOXKQzM
h0SVVX9K+5JdkehwGZ3tVcecktCNq0+ymHg+0GUTsItaPL64TDRq84pDWwkg
Yz+gCcxo53AxlocqXsy7gXLYkbOxeVsS6eUclIwVQuU2dsOp0R91tERFhj9Y
GBe/yvIEzrblmMaH0mAZn0dlNvyYCLR4H3ryGId+w3//ZTsJ4XQB/v7i9ztb
gZlQlqSM8UcrVgO8jkdhcH3YiHE5BYc5fUVq1ZkwX1Q+zlBU1BZ6rydwMumw
7kfb4P3OhyvhYMzBo0iSy2sWGGHCTgkhpSnavlrYcYGW4gkt2LcZKovbEgta
fPjnz7zDeMi03FN/PEHbTUzERdDlzwBYLtDv586Zn+fQp/VdT6H9tKCew70S
4ml/ZGx6OXaWBOWmY6Kq3MzQH5VbBfFgoh2T5sM4R44+xnuhjR5+tjSZWxIe
4urICg67EdyeBbm7gZ0+BLTJbDy/m0/D1EpLVRBr7hCr0RTZp1ecSsNDczF3
QNuH/RYWBqaz3TNM7NVR9fZ0g8EmlZqimX8FVxco5KWakeonvSzBIvtOb1yW
wmA9O+zR5KMBX/RC8BH+tt/c3o5sHOpjmsCNXjeqI6eLPEQ+ccIQAvrxOVMF
aq3SxVPJ34lYoZxAgU0kuE5g/SqTY1d7+GsGfyHY/qdRCGzWCxGEDOriYi+Z
YWS2n5HnjnZzgLIVw1i/tSYPiC4Du+aCwIktnmMRgAfhTf3i1UOPjv4Xpy1X
NO/FiZso15SEFEM/+ymmW+jcMZL/AnPeLNCklMyqmsYrIBkye6pZmIgwMyNU
ZCloIJshuRrxfJOoxzvORxoDdSWJd0y9oEGvz/ogje+sBb6Ym0xTBTsv1pQb
Tqvob6nW7+TAZi4e8/b8bQ5OnLl8ZY5GyciYcL6Ro4iqmlkJZ1EKqUOS+zsr
ef4L1BLrjJK3MR48ggoAVDCoc2fpfOLnJorqnynKWbA1YeIIJUqA4O5/xSHW
Leyw1pH/aFl0lwLOn5ZrE26EVm6eoynpfL/RzeJ7AVa0HjMKfdXbZLMxHMZl
Ggg5byKKGh0hSayeUblU7ZDkBve7pOQTEgmvLLQ39anznl5/nOxzAeNF8sGA
KkuCYBFwE8IocCjsa3Rs3KH2J0zLMJ0JQ3M2juQLh6eC+/HQmPQwN9lqmIQu
Xa0izgLvDPh7CMOqUcueHbCC3z0FscpTSGstwNmeNjrOEXb9I+2LE7cMq1F1
oBGOclNjZ/QMpegr5QVBJpCSNsB+qQ4LB8pneBMmSTXHvzx8S1ggAdWDb1Yt
QMaNjIdZNSfAOktlCaSw7lCJ6+qDU0tXN0xH7doa0g5bfhpHq/DUj+mtFD92
KVozsKUTHAwQ+5PjbKiVAznA9UC73UJ6TGMjPBzamuLxDlrKEKmr9kJ8jm4x
mEhDSLWn9SpulOsnY1t7F4VHzDr3mTBZNYeySDmy/6o4uC6QNWt37wGMoApe
onQUfzf5XV6LkmQY74P3RCyO4k2Utz5Plul3mQdQWLj9WX7P48fi4hkbZ08y
nT+3AALYnBQgvlHgFEG0ydFyWPgd8wHJPBJ2gYovu0x8edvXpoXFBKDdoFtQ
pv3M/Khbp/C5uu2E1g9AF/MRAdYhHP0z5qMwHRrdzLh7gxIyS/Dqgr9kbRXF
IKj5oHZyIXUqi5wH6r/mT0uu6xg7Ddz+gQcRvZNiCOuXph+U/1W+zlMdGGgC
i6CeZKoFPpc43qOfAihPcLuH+J6YePdSRJPgBbsqKkCGGwz3F0Omjs6xIrsW
JwO08+0hyEIQxPBRNSOlmgM9Ny2HFozlBknaMyogAlCLdyHMe3IOjSuPmGms
J7KlhvfuSoPEbe/8HdBdlvvElGjfYJYumt72Vq1cxXjS85SmF3c7XNdJ6aHM
t2HR01SQdhJnubg2HA/PyXVtVm2WKJ0omm5ZhmJ5otgB4vfE9nJAU46ehCCB
AbEw8y8LvzxM86daxe3f/MNH6oGCBEYS206WxaVAPsWM7hbEGcGT09laTAvv
u3Fy5w+gtePGZdOZsZh3rn26VoCz99Lr292gEfWPXhtd3wYZ54ajJnE6jiOk
TF1Bh0XzXRJx5o5WEI3sRTfKoZvj9bW2WZ+Vo2VUQQZSFrnTVCRnZtu5T7BS
oJ0d/PF0VeFS7jrh/PPF125Qoj/yT7NMjbl4Goajg+19+kLP+U8J32OoslYv
YVq8VeQ3OiHmfTooOABj8J3dbm7sgN2f/3/gog5BtxpOjy3Byp1p0czBrl0i
iOpYpTgIkG7POkdh45Vyt2x9+uN7ShYKeIvQwWTF2S4PFteg4E2zjEX1ebhC
dM0K+qkAPe9tLIEX0/pCl2EHsmbWqT0Ie4ELoTauiqoT32Bwqpc/tzKMb55M
7c+VUb4VfhMt27oVULS2Ibvn30UoRRrnYRZaFSv6PeYEpeu9Z2Oud40o0p7a
pluY4wjP0vdUZDJ1omCZsUorDBCpqoMcM7MEtvz0cutCE8Gp/lQdKjnJ3v5q
sXBqdv/tgqC4b03KrmcvbXPw4BiMbGIUlrc58uN8PonADAwG3bDXqWKNknFo
JgUJMAbjBai/kgUUFvl/d/Hwr7/GfvfA4UKKf961c3dblWx3nFBedNlfg37o
qsCx4d5vOv8hIPlGuMRFSw+3TFHcSS+rwvMU33/rll0JzKb0aNeQXrgqdYSR
37BiAmmZ00KOtYTcGSexwQByvn8aUBhkG3i0Trgak2PsCDZSbHh7YqrMNUXa
zfVq2s8XSLwlHESVVfHpGsaRByN+8Xftz3EnCZMo86ThKQFzgIXFz820CykH
cwu6PSG94cxbubcEJ2OB2S1pb2z7ZASmZ1asle6L0Mc1aQ3fhvcDF9ZBiVjJ
NOAJIM1OxV0wqHW0f7g6fS9OKp8V//avxbGq4CGvUOZAnHe8XSfr1op7IzhY
o5n4W82E02yLUWb8dbDnXJWDBaS10wn2MDWHCb90wQY3hTsObjWsg5/uai3E
K5RgJCO1H3X2iLnDAU30vIKu3zeBlIxIbmg5r7NhgT3OmRItxjJnFRP30ZAn
XTUq32IAtRdOISdv3O+tmyZyfIRWfwV3tfy0F6ipzfRfP+tuyMSLCIXtCptF
omDcZAEfSxpVfOl2yPn4aMmmPLeHye0vq5O0ZR8dbFcviLLHgxWJjlYYviEN
MIW9FNVr0ceGmgzRAnubbmRinHy1r5FCKb+LdcExlPlRqwg3cPGiAXHfxa+h
Hj9QFZ5nPjQ1TvVisSImtJsppd5XYQwv9cjpxKgfErCxYUD84Td0eTdm06rZ
b9Sxy/bPbZo50tT6FtszalllSn5PJabl6LyT0c0cYF/7Lajrr1IXkPia0JE9
AtgHY24BEfyaUT42ZjuIoCveS7OxKYFbiMKV5LbZaVOcEP9ORqh66oaj5RKj
3ETZKfmG+gKLA7gEnKuFl8ksnqiWOhnwQiPHQO5YZNu0CDZkMziVY3iOykIF
7Subk+bKyacrmr5mNHE3ZamRWyVZ5yUIeZAn27HcwFsU6MAxmUAoBhnuhuf9
B70EviYsEkso+vopGF9He/ZoYtRRDNzfgJR8fI/cDFrsYuX7OaNSgcwy9UMz
1C1Uocrl5y0UZ5QDTTGPTOOO3taPYnQaM1/vVV9qOQA71iOKKbUjPtgOhy9V
CfAL2UnLcDUnHxd+SRzYcdcxL0NTOCfjIcIT0mQYDjvgMozIAA1Z6S5Ikv2g
VhTpZvb/1M1X5Vqy7ysRKTGLBwEzUKj15mkQGks/djXN29IrRLwVWQRcnKua
/v3VIjYxAuJnPh585D0PoKL31dNNQ2hOVG9ax4xm6rD96Jf3VpcXyPGmlwp6
Ltzy3JypoRC6C1HexlXZ/ze+yATJdNAXx1SK9zLq/6SjA2O/prcCM3sN4Gfw
vBbYjcxTithOD7Xt/u7jPBvYxDJColjx4vYYJHDfRQyqi51e6J9DuZPp/gBa
ZZYb5RDRCRfFjwyRRddUvaly3M9KJh1WbcwCQlnOQ6xm3kQlrOarrG+KMk+X
AmzzE9T2AHK73UpeWmMYgid3TLujFuCJtJJecRxI7rzXbGlouPcRIMWLmhre
Ry2hv/jZEfWFP3JD2q8cTNrcsjWDKDjpPLzd6qf8aYZJiFyXPArTIfVaPE0E
m+Cw1XIUUpIrNzW7N+5C4P4e/lRlE1DBENhdAJFGv8IyrG5mC7nQOTqUR/zj
+7XSUJlN/oIOoEjrZ5aRrWHz/4+0BYMwp/tRoBxTbtS3aSp9JLfpu45QJ8pL
DrIZeps0QQQ3XI56204dMEE7ka/m/xcXBTXTGg0Ah47KrwpuZogOFRxzkqlx
2PC+IE51gYCUYUv0RMQWZ7GIddwW4wg04F/xWe9JxvN4cA36PUNmqKFndnPP
Pur6WllFpMR1BtrpXkL4JURMdxGCbgOYV1j3EJHGAljJpUVkVEegNn8v51Xx
XeIwO/tCyngz24uFrQlbV5uevnYb+NfrBDYviF9p/7543WgbS8Rvi9CjNOsC
gU9bTQmJhVlmJemKHDbjHH7KZ5xBF1KYvFw6j0FaJU5jT3807VXBkLN9j8WP
/6+CrDUGw4Xe39uLbQkQgG4VlyXAFO3gNHjxSoLd7WtB3JxWsZs0w0xb2ytQ
dtw7B15tPb1N5eVjWNLS6Bb9Qn9on/Y7cbk+fBLHbXODqI2Vu2qK9qjvnOgp
9s9xTEiqJ9ZLvF3uNMpI+7/bZcCyNsbY90dES1i9m4idXDb9e0aXnlXtBBop
btBB+auB7Pb6ljEDHmzN0Cqod5sEc9MLbgprRcjN0N2VcmleXhroL0V69q7x
b4glgUAlJYQT575zW/OZst4kXeTSrSKhlAhoc8H8it103zXE18wKSrC60ioe
+S2rxBGHFR5zhyxCKZ8qQszmz8D3eAdnPKjDDakmooDSpMzRM3MJAPvu2ANN
MwTMeiAJUyWVOUC1fXe2t/jF7/cvN8AxSJO5XZUh8mmdTCiuQrrSdIgWS/2U
Mpn1bvZrUKiMSDP/HoVYbEofa2BG/fMpe+qShBf6qoNyTAHRVx7bbJXzjk7L
/z4jwLYXBwY4Yq/O3jzzseobdfd955DcMdb7gtQhe4Gwr63IC45rxadVIfVl
fJW1AhyoMGRUoyiHJDwqbp9VJ6NvmIpze80NMxYnnbaichW68adJxf+khMHy
7jXYBkd0nWbWV1lC93O95ICcwh1YE9em5U37RoQB0jRq1z5aNiGtbpW3e2Ex
b3M8+sTftMTBI8GtjrM6ElpHMkAGWDNr3UeaUCvFM2U5cnH4w62FkOBhb0qm
aW+E52obtbh225l5MYR60EP3iE0YJYSfLioy8mYvBA8fOydMbv+VJiZSN0et
NVW5djd/SFEjaFl+NPYecwMrn022qh4SX5j5bxq4NfJOJbTS0JLfs3KtnKo9
g6gDLSToFuTh4Hn0zgsd0LOkRMKNWALLc3WkuTJrKfys9IWKC/2sBtX45+ha
bGAWaFjmn1XbHK5FIfE0aHyecgfo+HQIShsYHYkViT544Ptn66HwqkCCHjEA
Fv4IjH6FJBGIC7D3Qdh5aRD3919aCn9iJfCept7ShhXPEjhJm3q6xVtckz+9
MaMX5e7YRlL5KhT4YkGi/YMCfy2d2KedlYkoppuD0WYRR54xHBrH0Ht94efH
KgYywiPek/PLuRRRSqRN76Q2Y7PbWLBXYCZa/EivvXurfOVgs3YqkRAFhejP
dZmobaAHY23G4SQ3YLEdZLxXmYuIWLi+WlVHIobh9AMuzqi698KNCelvpgFG
z2qkwBJOG1BzAMUXXznlWClWnktCy5iSJE3/uRgX7qUaHNaPKzEB7Pphd1Fo
aAwmNwZfqg1ouND1YjXSw+N7VDv+7lDuN50OE3d0a6ViGM21H8MSmrzo8Cs8
qmaaJ/mGMvDdsEIb1U7KE65RsPBc6+KcDtyVxzoQ6Fns8c1bM6ymJ2iwMPEy
NyWfA5iVR2urfrAGY53eQW5DKzmv36EZg2Pe+eaJVbqWcjoHv/MpFqbJHZW4
jzEzMtzhfCW8P8MX6iw9bkIc9JLaJuDrpGvBo4HswzUCN/W3hJjNbSJU5DM5
V7hwWOVLq5dgaFrPDiTQqUcDyu4t56RljncMj/N7AF4egrEyZskR3WBh0Cjf
MMaebOX+DdOM5GgeG6NOleYsWZlNzJVtrUWDAyH4ka7WZEqJu43KngNGF31r
Ja/PtFiQV1gLiwnffrtiDyjZ3gT3g/8sTTgo24Tb5W/vT5NHKPJgB1VK3O8e
75DnyolmfpP4nU0FngV0chyzNjypVImZ9yJOosOHMfGSjqbOa6R/CQompp5g
RD6lUl/QbC7x1ZxT/eAdseAsQIYNohNVK9bU5VbxPnb+jFCczUFSMS3A+YHj
lvyd8+31cGVP/cX5oR+7oB/zNDQGtIiKhM5Xi3/pSgtwVZbJO7W9Nl3I2/6j
EpNc26Uk6s3W1FBV2Rufo7t2rcOO5Ffov+1pPuTmj3reM3FzXsVYNyc25lLb
PvliP06wSFx5vA0hnkb+2n/yZ51ArUG5GvSKmEiSwi0U6z+YX5j1qLHyW96C
NGCIJReIzUPi0bwAi1mkA78PyBl2vQLX0/ReTJJtDTWievjYxWiEJQMppp1Q
vjQ6WVNoDIA2zbt3Ji4Gz2wnR3a/avhjHQRl76q0heaSrFMeyqDvVVivEpvr
7qFrsVxTKCY0lscNXgkv+CeVPnBNPVNPqtOeoV2NcsHZnD6C+qmLCJUIPB/v
eoI0+zOSb+EWeaR13YZ1fNkh8PEmZoA+8vo22us4t21vAcAat7soLU5hFm1C
JbHuPIBCG9RBzyAqCdkS8jGyN+OYz+gTpNpDy7vfPs9YpCo0N6OG2QwEB9Iq
ZAoPfZBAF03GHFSJAQxyWE3zhPWVgBf5p2oIhQ5ocIvALPIAk06H91SSvrmL
vyOwIKZtyxrqz93WAZyKTnVDepUUoqahSyWPsbapicBt1X8RIIC3YV7CQVWD
ZQ+AVMoE7VjfP3o29BDAEksY2IKGGWsLjZUBVcSYh6ZApQN99Xz5f2cO2Oqs
gy0rX2G6JaczYmvvVKm31gFvFzmB3vIpGpIR0PfImPI33S700sobkj5of1k0
D3Klmn1IwgQwEMav5TJYsJKaeMYD8d8fHn3nTLEGjYXgW7j7LdGFyWx9h5fx
PxrkwKyx/JQdty2e83NRCgwnA2V7cNS/NdA9aoGmZ/iQNuOematAzlAYreWh
4pxjQMPCtAzt5IwekOxhfe5o13Op0boxi0JDZRcOWkn1pJwtSRVoxqcxwpFQ
x0gRNHVJ0I9dx8hlD8bAH4TGF8bGgEygeDWVl0bmI3Wjp8Q9lDYBe267+BTJ
nid69n5NBh1J0tfSEWh9f3i/Ab0XQtbBXIzXpUv5ji6zhXYRb73Ow6Qs3hC0
BFlO1D4IjfId7C1RI9rlPbeN8sH7SrUHh2WTk/h5BnOP5pQdq0K5s+QNK9Wo
+7YsNodlBXNO+2IEG/aiRwhGZBPOQGwW6+o7xZFsGlAE3Yr+w2/Sr/uk4bip
crd8O/OS0ZwwO36VcJNZoZ9hZe0/yLYcRDGKuYjflxoL1HRHhYvhg+aGewXJ
Npq6xnJ4qH+QjQQWBrYtWjOGsThM6XIKuHa/+BD+SHcgM6/c3lrmNt5qSHlQ
DZx1alZ8sU/80VBFLRCgIjS7OM2j5ZG6skSzcZlD88GH0cdvimKMj3EI4h3c
hz7B9X0J74NLU/JrPByDYyfGARcVB0SgLYMrJLre5cCiXT0mZOW5FS8xEoq8
kKQlVEzG9gkG4CsDFSRm+fmW3DAd1yAtVYpwBVFJ3kv5Z+tHlS9FC+SvoOnh
wTvLMQhQOr9st9PygB6LT92PWvDrYekrPrwjOhEGhv9tU3UAj5xsr+R32jiq
ZJaLJj7jqls84vm9cOK6wFxjrnl/E6iINivEbFikewp3davUqqlw/pIANBlc
obFGUOhPLKBjl3ByJuT5jUbiHeI49wW6PcB/sY/Pg2gJnY9GHfCq4rx/4euN
wQ7Et9r0zoyJUxMlb3A8VJpz3rru5Iez2X6Wrvy726Dbx4kMJ1+TlTvMbf4F
ucrnmqxeF8iiVZEfdOHzczmYBfhBCSFI9aaxVjL0xvqsL7Udao8yFLNG7YfD
LcBX/Ob0HoZ0AGTGTQLCYfvEcE/gISQB3Oimugg2oFWlVyQ7f+A8tLzV/5dr
1Aj6vhkmgjb7nTrvrRB3vX1L0ZbuRDde2pYhG1atjXcBoQU3vdCI0dqOevHw
gBOeIWMHsqVaNaKhOnc8HGMuzYSeWhGXaLai7tXG7HDi6GUdjagIDKxiGoB7
9yGH3mUeC51uRnGNZ8Fi92kDBi3jmoQ7Kf2D/KMtz3+D0K2LneMcSHns713H
SuD1I6m64LOpKFy8LNqD/Flo7lSplbt+akmYQc9uuzA2hy/Vk7fayglZRUE7
nadh+SEh8mKaUP8u59WovhTq7GM9V6i51qHsuYdasp3/pccRnLmc9PwT5Fj0
b5Ye73q9Hpma96/CMGyxSrJ8ySF8bABGSnNcLz0sPlfy/IEwxV0QDsmbs510
wTL5mrM0UoNZ8CNrM7C5qR95LMuOxzcJdvtEPJQf09JB2StdRl+5ujqCjKXP
DP1PMpF+K+qouU/5IsIGAfHB4A2pHI38ULYzbKjID830Y1EqIrf9Mej617k3
YGKHX4b8CVxb1P+cvKzobh++WFzvFP2CMz4V/TnzbJFjS0/GjYT9pfTD5O4k
Po/rBS7YbvtibeEJPodGNSbr/HLTzHvL+RcrnymzFWs2mmwnq+WcP0oQLkF7
XNqxabVm2eZ70UCMSZ+WHNJIfaiN5eCS216MmVxHBZUkDXSSLtQXfyALOhq9
4Stv/B/rBC3zuTYzMZjTJetD31uC7m6lO1s6aNAbe1G1jAkwySFCo8f3I1og
UNiI9dZMYBS1IzTY/n9p0KA2BdVllT5qZOqO8TdqRdd7rPx/URU+37pj1Py9
qcBJfFoBXivQK/lixKyew6YhqZer2QMZBZcHwvDMvTWW22UDx2d8fBQH699k
ew/2kA97fAOq63BzhDuD1cHOoA/LSi2utg0X4FAD557HugNO+Q2kLVLjXln9
+6mvgEo2Wyo5s3N9gecbKGEa6W6hfdvQeQZKIZpHc/xq8+h2+pQlIu1VfRA2
Du1lchMcILf94btIzekWD1GplIqou/El8vOqEnR1Zyg8hSZitAOolNL9CPcU
siFdCCrfaGL2yq4/Y2HuE14/j9SRjmXJni+W5jADjnbu3mvkbTqw7fEue3w5
vOI4dNjSnzSnQxINcdFmeJBTdDjlQqIuthuyHZot9eTffqWRnaY/vV2spTAm
v/I44Ty0LmPb4QGuAnYbSAez5UOXYJ5FkRN2c43AD31NW5BW8Rfw0dupKSkB
DwlTfvdQW6BhdgO3HDoKnqYN1prpZfGdcJz9mQrNsaHZiOSkkEYLR8TLoC1+
1Zv/QG+hPdmEtrodHeQfV7d/FECNL/UEFMwGlXIMQFMJCNGDw0vkZCRrnEDL
T+64tvT7yPpZomJkYF+KTlr08ydk4k9P9ZcMQa9KCVEZw24B2EwTIXTLTf6i
cNERzSgMZC4A7D2SAmhBbHFcWK0zoRFm5pj6oGm6M/y+rkI13Gv4kPHdaPJr
/Oj/kqaD69tg/Ps7X9cxIy++dCgyF/qTBVLXfO/xsoTSEVUO7w0ZlxbcSkgp
yxXkLXMcgS8XozVjAkCSiJ5x7EpuG4loSfu2eqGa2MhbO32/Qw+54zoROVlN
Ccibywp31rX3cMKvbbK3hrUvjj0QRCpr2Zrg3rhwScM0EVdMpWDMdyBvIcQP
X0HwV+dNWAmqbXLmQbFYLm+0nKvEg7MF3jRCx0mgxZGxz5nEKK4K88PuiESh
kdN/5jkWRwWZplfpPqgYQlX3Iu9I/mQGVcGAO2IDY4XzHecTFeTUgRrB5Vuy
IGZ9mL8eTpWQxmnl+e3MaBtERfWJpq1uOsG02aRPO0ejny6ISv3K9fklh/ec
bwH2kfIGZ0nhLvpC9Fx9ckBkMN//HU11gbQrMhxxaZLhGLmqc0c1ZOibhAeQ
cD77zrX1yspxbtPY2GNK8kUTM3AVR5BXMKYXupCYAs7reYOY/5nrqrm1eHaY
FDBA7W0q6zXwChoEpV4rFQyG4rHcdlt0K42ceUlFBOm+Iuy9e5WBEhYUTg1d
YDghdUJ8Wz15E/BEmr353qra7Q9A/L+YUk7x7yq4lV64dgp6TOQyJUz9Q/wB
xoaq0s3nbYMbulLRGw9qXONm9XHAynVZTXwEtbsAEkr1WgJ4XxKEurfdzj4U
P/NXeg6AioJkJziz+pra7Shoq0osE3ULjQ3cjKvk2CBlYX0sAtYPn9BRzWMB
mZp6VflR2SQYlkKNgHuK+BDlRh56APQhfXl6XGd+obbaS3J0J0wJtEyE29Q3
mDgqcVM9zzs42E6/VUPEiHy9lxDbLQJ1UCnJdn70KRx8ceUZ+ie9eytnQ95C
xXRwqYG68OIh+HFpzb00WiyaLRc9DP6Nir+JOdfcEBTbXDGw7b3fb3/aA1fD
iXEBTjtItMppgosMq+ahjAMv0V++iBSW0wkiyAlZLeA//FWAjqCuXBAb1qnp
QtUzmjoflkpmw98/M6trQfUraAaFCN2AhsD6Z3oqcVxBwJ0uXzDPDzv86hgk
xh/HbptlFLlDRP3uxU08d4faZARwJXcuFEwr0kbQMLAjjXM4NNWvIu+pD9Vk
XLtX+fGb3yC9DdxECowWNwJcrjuk/WugReffzoUVy5AHyNlMI/lzZSK3tlYv
NfOzB4tTaRbYKzEibk5j2mkqhhuH8ffigCkFhCjrG3MVs9tmUm1NlYRJd6Wu
8WZW5xsDetacDE21MPGZ7HIq+0mj6mYFiVGV7ktrCHCfc0gzta5K6i7UkavC
rJx9xIhVQYXkE2c9m7K0QlZVOg2KgWZ1VVlAWTDtpyeXDQEbLcy3ltC2wfN2
kN6JMtB0FIxeKZq076AronBancnkxHxUPxeZLT9aW5u+87O4Jmr894FBzPQl
miVAhNW/xqTo2qWC/feZpsgmd7LWVn5qKmemiCo9bFWCTKtkBhjbUUljz4/S
t4Vkb17U37/Rfw8apl5Uf5/CpPBqttIKOYsjiY/uMbaUVVpRetqKz58VBssn
BUzpqVdwZeuMUKKGDtZSClzg1JL9iCh4wND48Yqvlf1QjHqPA1tnI/aMm7cs
1/qnCLz9YxsKxkd9nWHtho9iwdUGnSDwy1jiRw9uNtu4BI50PTpDLCdvCFPQ
XB5snmUzGxoI6unuyx4dW1op1EnDYAn4iGdlaeUMxtGOEflHSoiuqU4tHIQa
WEXhtT2ucx1k6R0q1Oish6z3KyePZly4bI2Gv02vUBgl1THI81zsl/CApYWk
9Lx1FKSN8WQQQp8Dv6gUtlDNkwDc5acXGX0OKk2fE+knsBNNswRb52Qvp2mS
QHICxq2v4lmI9Ypr79jSqKt2od9Fr6zqy1IF4t4BA08dxaJrGnfcFI3vxw5y
EnloyAmiyFzbRfkuXCeO3+AK7kENWEvT05bbL2cQpwMBPrjl2XbWpf1D/0bN
57zzTtGx7lG/MhGje1mco43kt1I7WuF1M4a/2AzQRHWa+YWHpOFEZwlI/HrA
SlZOWf41AVm2taGC3zMY5dulKnupjkyuWi3fHjO+gPKUEF9PT00KN2vJkM9v
8EkCMTjVbuDon3PVzdUF7PQhrUr9Vrov+boEizjklquYfMOsefl+Wp4fLodz
B8uc+4s+/P6YfdIQcbkbozhKT4y6ASdlETSjbcUM3qQHemgJTitj0tif7EB6
+wrsd3O0Rq9LxrndOoAGVMONyCg24qhKFs9T9UWZJiBdU4C82Rb3sg+veJn5
3eJACIw1RPN4FrXhgxIOMcapjAWOC2Ss92OVT8S57lLIe5dD/paahzayTPt0
oozl4jipFzWWwFp1wu5VV4m/6wOwPdShHWWICfxywZpr3GYg6FzNm0HJhcsY
L8uTy/QW/hD2elyTgTPARDOtYIn6I70Jw0glm/K0TE7hiAOBmW2+IYiK6IGm
l54r4NvAH1LrrgdgyHkycg38+1bvUQpTtTn9p5zoZHNqMa4PjQsAoD3UyQ2I
TdXvHNUgNucUs8i7j2Yw/mwisD38dqBWgiCHZg9B7jkscDBaqQ5sjoZotX6W
mTHyLKPvoTLVxhOXiu0jVzCg13q8Jvi1i7KyaHloVjX6E11bTWqPUcQA9BX0
rUL4Co+e0lZ86JhwFpMwPKFF0driMW5QsIxy4JuNNWCeKW8cEIzYPZmalHAi
YbppxjwbeL7Ezw9zPTZkzxRYJ1AR6XlS8OGqfTpPMPqjkhL1QqnS9qWxJJng
Ttw4KH/xaNYhb/SV3CP5DLegHXSseGnoKFV4EKCyzrpbAaPyefkuKfrdfOYA
2aEn0lynxcKVSfRi1tH0O4Hlz3WaL4cuNRVjqZXnmVUFbRAzB+xC93Ztau92
cpfaD5MmKa9HODi+sC2B5xNA4zQIHiwe5vcU+ghOI1jomb+CLrRreXk+kuU0
T/p7W1J9x9SIoVN8DExxRXAak2IubK/uNRAsrcniz/X5iiowY9Q4gXgvuT25
xKdw83Q2yPeojD0gqHNBw3DQtsD7B/yBNBIEZL4pExb8yU0kVqyCfBP7F/sp
i/oyuyTxAPmggHaV0k9umT0gDW1oUawwR7e/Ba7N77TrdU3rkb6y5XTGHH7c
JXoIHjqHOZumHFqNxf5Y64NKai7YUFZbtb+kwQkr5dNFw6A37kec7mBDwH82
4FOL++STgWX0aK4NMGB/ZAyKkcJnLnUKJqm+DUZrw6QEs2emdFZpDg21t8Ku
1kmFyoDu1kZTiVdZ0XE+IefoEHIBp/TCFK5pPJu5uwfT69200rpHUJrSiRBC
Op2JrpZd8VHZ5oj+fG9YFYGzo65lnbaOMt8A+rj3WrJRd7OsOqJokuRUH6st
ywfsuZ4NKX+6hT69Uv8ghqZrLloaPAjXqUDS4lA6LIeImpDvrK/sC2X1Y7w8
9ib96bxcv0qlRSwKQ2X+HFCkIkTgncLltDndDEC+LlertBDKdqS20l4YEwwr
pt/WcZtPlJUoy9e7y+bl1FPQBxoC4CjaAYzjm25batWy73f4ENzh5d7DyJpl
7g2ohA1gH+6cbKpCedYFpdVNQYNQMGElsiJKeM1l1NEKYFSdi01xBlZkd2jm
w7fRw3VbVutguYaH2rnIlY287X+POtvoL41Rf47bbZQ1TU9yUlQZ4XfuWB+b
r2ycPZykBpzTTchciBwU18TF9CB5I0TNZmxEvA4OGuxCzs8zKNkGAQhPhI4o
m5N71FiYLbHMaj+gL+3ROg8omTkvIgbnMfPNg4vDCsom8KX2lDG7x/Xu6uJJ
OyYjjs9RlR4wk/gAFGiv6T0fQfS3gzQxDEUf/zb9ywhNxmZpR6arYwRgPTSY
UXDXShs+gJ8MeMZngZa0esDSx1LmEXNTK9rB/zUDyNXtqACTcYi61Xb/TW/S
RsNhdsz9xfz37UAEs3mWNn+BfN3YOdkeBbXcVXlQfX2MXBJdbsgIcuEyJuHV
GdClQFonH4Fjg1n/IjRpKCXKKrb8sN0zXwDU36Z35JYkhrJUCdiNSzz0f/d7
Diq6hYIN8B4MoATLUU+cp+7kea61mSP2T8pQBVKtpWb0QP28JRvaD6CYsbH5
a+c7NNxRTmaUlic6wYPRfNHKKiY7UIyv68++8ueonWGyq1ZnWmAe8Vih7jzA
yW0CXk+Vx+24vhq06CMt5YHmoBGThLn/wGbnSMtDaXuBkT00W3ZGGvdT74Ur
DAfammNfXEeD5lefCKcnwCukHOWobyQU+35SMzmJOR946iGqhi2EAJuo8vCV
IKdNCqRMDDGIs3xrGjnQRaAeZgR8eeDPDddlOwVyw9TDPVuXVKmZs0HlEga3
1nP38R2pIZcNIfgBP2sDHrB/0TS64KmR5R6ZGa+EoJWkLeHtBQ5LKmWYXJXu
qOhIm8IPjbg7ikKAb9CdKPyi5v8hRjjrAyF22xj6f0l39Uf2LMvD3rPoSbaJ
iMdieHJ4ky99tKHziJBmhSJ92v9vX1CqPp68bjRybkIk6LmjiMhADoD6R90G
A+gBGJY/Dq5M3iHTWdaWjZjGlzyoU6u/nZGLJrq9yYIMz1BEPRaEAmgcqoJA
72jvKP2TJ5qbQCIE5qjRf+fOoI1KJFVIZFz67CQBbAyZQgD+CJ4aKFOo5tjr
Wx4YQ2kAiomtc3WOx/tnzVTTwp7/b1hKZmM5z44gInTacMySxEk1rIdSd0rA
nBkmBwMFuxn1cJ8Sardc6p59SMw4E7v1IGuYFAZ/2IRwXdkRXhja4i/x84KR
9BzOtRD73VuH1U9slTNHmu+odmVVZEvE1pICwv7tLTkjtG6vFKZC3LGMfqXX
anm7dLEJlv2PohOXOLN0QSOxk0xrtqvOhKKWtO1/8vDk1o+ftq5bIuc9SYVC
6CVu+wT79l17XBt0cJnJLAYs/rMoYk4uBF8GRKeCqP0lt0d6ehLQ0S4Dm4pM
m1Q8opwRQ3uSX0scJ08Bac0Fo5xdAmUoB09ga1Kv6zb5icmp2cvfFG1CwNJ7
EGwhvqG8IEolaTcGf5ml/G1oKrUPTYeM2At9pOngVD+IoWGVxoTkNLqc2nKz
eU5FK8vRfbu7eeBSBes6ye/RpCpqTsNAYzkjEZXAiWTXFNOfToA/SSXdaCZD
ZWyHciS/GO9gdy7U9XRg+k0OoxidMS8mRq7zqu9+udmsf6swOWXzrN14TzPE
xcTYfUguD3R06pt0Pb/yl/orDZelZItsN6s66arHLpEE69m+cPWNpeSSrz7w
FXh9LwGDq26gMjkk0MSmzcmz83ckbETMwNfSFhWanHIWns4fvVJP/St9GAW5
R6g0HKS42FaGd9bKp3dPbaP7kP/VVBsrtP4HqbWS8dbbc+te9flQanpqztvA
s5K6tONgcdqvtjbokG/wa9uz1m6i4xHVj7yZ+UGF2NhanJApaa90bGjY0joL
Ix9LulLLMipwDJHfj1IVbWRqDJr6f8nxrumAZcmyk9b0iPFOTeKCPHo+lQBh
REuYVQBvoQxY19wl+CzaKCoUYLOO7kY5B2m/M4tsf9MywZTb20bKFOgrpmbO
0F/mIwFlhbE91X0saHpRiyOY27hgpb27joDXWcYoJTCPu50xTYORups5vr+u
nuwoccdgsSWZrRnUzE2zuvfXIXqUEwH1dHJTo5VqLddm+fdPPxKsHwPEeJMe
1Vxwmx9svIqBND2b00S8IpuH42FcLhzC9V6mG3QMU/ifc62q6vs9eOBHGnrb
/h5krXktF5oRFLjsWnfWrNa7rDSD7Fo2bHOOdqEN5POMPXr4q2CHBpPmzMKT
A11Uyhf6aatH0J1B9pKhx2ytMKflxImxW0U+6jBkhDGJmDiNFB3FQarpvnd1
+0IKo3rNpfDO+ER6T8Ztq1hn2UAmmh0poyO/fsJll7PV00nt2KI+ENb5EJqu
+3lHj84wb+wGQliJbPk2719xoSU4RnKfnDfCSN5lRuYSQZALJH0jHRU+Zf31
B2mCz6OGgiQU1wo9oGzGZVbx58Zypr8oVj/6aZOYvYbm84amoag79rrZoCa6
tEpj/gmrW4Ku6mlnmKzvkzMpRTWCUs9gg8MJ0FdtE1C7bOUmrJe1tqS3QMPE
H+c8uSygwDrfsc9bbKfng5z94WdZR88JK3tUtIV+LhjLOVtHd/vJYuddcRlg
drYB4d5krRlEIFHTeb6txmPXwxuM6+HSbCgcZKkdQzefNxi6QYvy6cLRsmki
OvmbjPDsqa8LsCQk5/OjBl3N/pG6BekJr16Hv0dqF4psP1bZ9MMI6I+14hE0
v/T+vNMmzggg96fDeR59MX4uzv+didEQlbSQ+LGqIOJ5sqoV8I6OWbsPGWI4
hYBrv9TBSqzwY0pQdBXU6FZiTNTFNYfV0uXHkQBB6EXoKRrMz36cbaBLvXKA
js03NnMbeI7zEAvKfZSbFt2BGiSmDC42z66jshBs9Va1yc2ngGfsfvmBdKur
xDV1Gcgt3nj031LxTRRx8J5qacTOvUysGK4U7lxlwtgtGVQdeXmgcospZvdP
bE/ys2etINmenCB4lwgon6of/mnkickH6W4fnh1nal8EX9m52ncdHtUuwqtT
aGWLnX96xR4Our/b8pCVCCZZYO/kcvY7JmAfsw43UkTBEo62NvjDL4R98DvB
ZTx5MxUYDlpWJWVUmSsXps9tV0w6qYVuBx6LopkB7fIsdozKAT/txVV/mI8X
qzmHMc3udCxYZQ83FVPhfsgCbqHgzsIKYJ2JgdFBduKA4MIDwYWgwi97V3R7
Isr/MWfhoQDav6oO1wJw8B4pgIlRW5ZjE7FUROXeX+bN+w6GHxNpTj8J9hPK
/jmfKpvCcgcaJd6FyWsx8HBcDb5ol+bKFGD9ES1C5Zm/9p0mgT5pnR4vEGof
3ZIPKYBafBFYPn6Py9jAdprmUEyRF3sNT4i9Uo2ATjBqueBckXCg3cC0Fz7A
R0538gUZ7560y9LkG/1TDSn1noZV6S6IjHvm5GrNSV6+2S91IitmbTskg1B5
yiClPSbr58QO5dMujXvD947wk+6e5bO8DoMAovGOM46ng9zijzfNsdqsGohV
MrELUFx6AuU8kTUYrCzFbPH3uGxYrXnXAMsqwKOjFkqrhc/40XnksWEs5X8x
WJcJLHKqZqxlM9ai9g9hVeRBC3Yud6VPk9XO+Z+nEXd3POn3QdVBvWgcxkgx
WApCEGpd+bZ5Uz43HwUG5iesZxK2RnLQv2k6EtzhTtPSA3SDc5Gto84ahKUw
2GwOjpR/VnS6FVTGcCiElFKW3HXUyXHx0l1ZmSd1tfUKiuL1wzSDcK/L8f23
6UIDApNqxjA4neCKBLwcHMTkKFKITn/tCFwwEHnf8hEawMtJcjBFEKUI+Pyz
yj90oyaMenwnSnHQ0dVis3HcqoSp+8oLM1WGtyp/euCIzqFKGVfezB8g4O42
5QPz7Sjj+9pzHIK2HdDp3Y1Y7B+qSyWvX3JjIPHTUdlXx46EQataYRNMkdBu
QwDzCM2w0mNs0cpZHSnytKfF5JNrqUghizFxv1s45+Oo1LoWNUhaWQfbg+7I
13CD/v++hmn2AtaXj1weliXOSI5BN/x9vjZAdVVw97+4fvscIO/Q/ZrdQUzv
tyX8rL5gGpKcSThRx4uYV2KiXb+lSOTa0sBU4Zl5gl43Mc5EH/hFCf/ERKE5
tutEVdcMjIYol/YPnZPV7a+FVcQH8YdA9NKT8DmKi0VwwmJQfNGMYsI8/ngv
l40XDdIPONBI9lyqbwYWj+SPP1YhUUMBafXvg2QnX0tGsfwqAHiJwP4Una6C
NkCwa6OpuUjXPltbD2NdaRj8fpyD3r1t63kij+RSwxlI5hSuvAlEE4jjOTQD
3/FiHr0cglJXUgtOg0Qnjr8k/NwJ64jx5FbTzD/ToTVBQXikd2G5j1JNuWb0
fgK3y3rmaQHIn29bXZIjXU9lelMIqqAKbV0Xah4eK9vZgAKCEsU4GjyvMwb/
OPsfQhFNIzyaCwyVDtwyfLv6kVP6/7IgxNfTP0t5U5LIXolnZX5jNFwEZahB
cGsWwC1OemVeHcpZBxf4EelE35GsXZxA3z8Yv/A+ZxUhGwkd8L0Mbht6SfKZ
xoCdw+5m088qZid+mGqh0B72eUXJYjsh+aZPLY1EzjHjxRdkAXgjIsDs+vMo
WWVKt+bpUB9OqVzEo0l4YxlB9bHO4c8foefQ+CHowb1suTY3saiWBKkPRnXw
Ic1ww9KSmMQ8ympE5cHH+ThrAZsPEmySIjv4tb/x5AMwNorD1NVJYyUv10v+
rfZUXaUYPlUC/t4FSB9VLEhHD+XQFolkRJUtqBeHFjsPKTeVA+Fz9CD7nTuR
g4sd/POTK7JvZeg38+TXW28rKBgx3bAxcThRLtV9ouzN7ZahxZSnjMqIbT4k
mG1yCyeEYvUXAurOr9WxZ1qm8BajPVIPDImGvCQvEqrZDCXGYK2BrMxmv91J
a5hY9kSEYHGh7NzvgUcine8nJv8NINEwvFemGd6aoNB0IbRnD4vmozEyFAUM
4nzQO9SRz/aRvcTkbAoz3GDoXfZ/pWylGieZXUSEFkVRNbMYQiiD2xbwiSh9
J6BDm6ZlCdxzaZsN9hYgD6xo3mgeRfwmwgszYNY4vbm/ELK0AEpXaVxak74p
EErkIsZ6zLk0epmwVx2OejUZCBpsxsrdvvnsEOu7b/p1Tkqdn08Uxtd2dRSX
N0Lo+jDtD/pAiuZsK89U6SaEQOEhGlp3//wn9/MiTWRIC7zvywYHzJkyasVe
Sscim/osOXHZynwA/V+kXThDFaq3LO9LFLDPCMoW7qQ1PHMOg0A6QWBtrLsd
PssSiUHWhQTfzaoiHOiSg0ZDuh8LTgaKDWj7oiRHr5XermDnKud5T4E837Yv
NEycW9aw72jrBqNKetJ52PwmXTbOZP3lxOqez+Hjl0v+8MG+2OIpVEp8DmrG
Lpge66A46G3NqwhoQ7zf3Ez+d7OjT3pfITCooC/rP/gqlVixUc6iVRrmGK8M
ErhllHve9sBUy1Ac+jWS2ifFry0lA0kcDxpYGFEsD2DqC1vPiSRbTcwVYG6E
djqVd1Z6T91gqUasI7OTOLH3n93AtVZjyVD6XLMSQVXHoBe2ODTI2dNmd7j6
LuyW4ekB/BVmdTC+qGVy+rBwlYzIRYZUROuTY1/JkOkQEL2a0kJhlfr+RlHd
+drZ50l3m+4syCceFw4Zs+R5jcFpOgSqgohBvN1FsVzzie2U0sSe1e3J2VIQ
pQX+KW6Q/B5ilcT0BKqycH+PgmYdIjaHTu0zBGJfXakZfO3s4K3qzjje+yce
08KYAze/ZO6u9DQ4X9iPqaTFAkS88O3yApTE2yI/+vaNT1RiuTemuvZWiOB+
6ByzHDZG2qY1hBBSkoWSLLeIaF3Wgzqyjcm/Qjcj/nweg1xM8PHmN8Du1b8u
wzn8FfpzXC7bvwFEgfMc8JlwPh/QPnPPCBKR2ndEUYqHdQ+KirnqOrDNSEMp
Cq6JXs62N3L/iV/4P5NWoaeEkytvHLaTa0mupX/kNvBaneXBXXnce988o3MY
hvRuKdJagAQ7QwwflYCDgc3WvVe8+n68LRi6TrWia/5dGVBUIPSoAKgtDnRJ
BAHfgXKb6h9mG5StzHpZBV96XhpUwnKwYVR1H2CCMG4HORHSbmJbytO3IuG9
cZB/gydtJltQjK32ne6JSWUaLfnJFD5r+JY2xnl25q4g/IVQM3QRaJ6Qe8MS
VK/D21dDebTC0KTPBvyxlmldh4tVv4wOEb0NBHgVIVgwQbOMzC1egkChLCa7
vtuJwEkcapQdXkw/IXqCqXu3EsvwpXV68K9tPlZ7f/3IXbDtcfnor7rztg+h
YRmKBeBFZ8O0tX/fDQ7hfF5iEYy2c1fSiPJ5GHYudaqwIo/2Pjkw/zhQHfhX
GUZousnSx2ToicqYcSG9YEycIhDsYKcZLMNgjCy6+CgN1NPaeJGB+jXv0b4X
xPa7hY06AO/dweMj2yU2ZQAAW9RUgGcS5PSVXbWn5S60nQAlg6rNShHB7pzJ
OQVKX/l8ryVCCpZ5c5pFwsGoKwmOORO9ztgKAHMFhNub85V8rh3EudGpsabM
pQC7dRT/RDpqCciKe+u/K3iu8TODpjVE8+vO0K6RVxW1aQBSCEfWTBmYsRD0
SXjSDZbMVAZGxXSFperTpFltFbg3aSBT4LFKoDqI5L3EhWLG6r+3BYTcvB+J
434pbj32Gjab0kwEW6H3P5cLfzxfrsFTkJFB9E+vt9cZC0HeWPtXdSCEPxzg
DAsk9KhpTRo14eHVzwoAbHKAlF+CWNlPqgapY93iyOr6JM8TpuXZnDkmuX4g
7Z+fsNMSQMcxp1HNke4CssjHdYqrNWvo8czaY5y6iXeTTDuUOU2hfgcyNC18
i2tXE2MuqV5EKXbJjpZ7P82hq960jFHQqSJmxje4MUax8VixueBZYtM7ePlB
bN50/LFZOY4tR3wwBoaIpmY1O7mncjW1dc2Zw59mdL9mWfMFnbP98mabUJwL
vbvs7V0fNzrLTOGmHcPcWAzuva+4yCcTb4HL8wQX42bl6Z4kdOZPUHDu7QpO
jZspek9hqyCM5lL1Zo6X9W5nXOrqBtNLuGpkHRUzUMwkSCIhrmGxas8BlPCO
R8gZWTNiJQQUUTDCeugrQ2leCmkGj+E9Sns1OcTphMNhcSMgWPdkgbbI4BjN
XRCXmdEy9fPKXL7ANO5jJDxROGag19rSi/iZsD5DmjLieVguV+6cpRUjvNXf
eHae7XJmA2ssOg3LHhLOrfRiJVlA3h2HaSnVilPDOj/MtrxJtYtqYV1nNaHx
qsdKRGkeB8gZXZfXGxjvWeMrUHT+PmkzLl+jsqNWKrO3+273EMFzQr4sycjZ
+OI6fnL59a0M+neob8n7d2GH981iPixYOhSRVYuBdMmKPcmjWzWY5qpLT6Lm
ZfNtqzh4BFFU6ccMDYgSoHn2g4bVIXPEHdMb/ftGnPykaYgMfOa/B2/MTVfP
mCeApZpx5YHbSQp1mvgSRh65UrNMgf9srmUuZhQ/vFYQxpXqs+pDmYSCBQw9
XDOoUsqX7DgcgCnc95FFCrld5hi8Z9egprYW67jMbmm48DZKRWWNwgyN/llE
wb6JEcwjcCus1jjNilhHG/MumhUtMSXseQd0SJTpDzJjl099HyCvf7YlAe3x
ZCmlPr/Q8mN6ooKBy4jpCZAJH7zQE4uqE4VEAP0MfmUqJK2sDA2ynfXtNExy
jv5AovcEhuntNEmUbBMyTfsZLr5Y/6o3o/W/Ak5Mm7rdjpiZmdQC8cAcSPg6
NiR2HS+w9rML4Hzo2ybB0hT9DgGUTuJRLA24gqif83sxN7rUHDlDP/BznPCa
3r1/TAt4Od4eN0exlI9qAquJey9z7Hl0mgemqBAzTJqLuN7HqXE4OXLXDTY+
SFmD0u2hE6u80qN08Asrfre92fZd6gja9yGsJ8gu+UjFKBNaXSc2DVKz/YgM
8BEMKZU8X5rL9No+KvKWn4KdTeGwaM39QjrOGumCN7/2QEQiFQAwV/H9beek
GoVzqEYdHmOZOG1w9zTtt7pg4fJC9lQ10EG9RmEOYtoQ69FQnmBuhX3imIk4
iZyPbOBB+4F8pdHZ3hxO5kyWEFc5kUumnGipAbh3HFHYAJXP0KE3/ElfYV08
WUQseMpYwq1XtQfF0Dp1YRoSk2gNRnLBHbdvTUSwqNlkpwDecktbW3a9Sfvr
TzKP+aBl76CcFSfiA35Fhfk5pgWMY2R0cyW1JL5KqG38HrcZZ0U0e/MFim67
3IIC3rYyJqQ6btYfIssF4mjXRuhcZcw8c/yXrqeTXxp8785Czy3DPJIINc7B
+dZbkJtSDPn+tnG60o7RamWXZpvIpQSPrwW8FpD+vzGNbVZzo9jFX+snZoYC
ZlPNhaTdOczBi5aJ/rF+abWT+zxFXxB/q6kuUtqSEzDsgkQQMDZVVg+V2sOv
M6vRpheY2mbMlUM4so5iV77DRhwkOXJUv+SVMJq32tZBKgmmWPEu9MXzAcZt
yNLXuTWegJQb6YeVx7yOdmaRIk4887YWPwXsa0/ca7kBq50xFhmHV+dB6h7r
brDQf55l5k0AsEefngxoOYOjSObUUfCAN8B1af/mCHZnik5fM+FYuwo8GhYk
eC7Z3z1dHZSvZAccSW2JJRf8YUdW3tLm52shKHDbOPMfgnHm5q//WipUJ3z1
jLfUt4lqksuGz0xUL0zB+yaCcLxMo05xtQOW+O/0O4gr9Bjog8SyNVwmYN15
pVPDmbFRpWjIoaDl+z/WXSvIt8eJuGRzQ9pISldGb5xpAkv/fwGOJIH1K26F
NFNdCOE/M4UOCtdTbrGP5PlmMGN48pze14xNHgA0HSTH+4wQNzRIYLBJZQhA
Xsh23q3iaSEDVw/HQMCGM4jPdC4EwIcRTywKT5dNBmesna9ADdDGV/9ptwtU
DpZQBDlFl83ftl9sr0OVOOpiw9t2OFWozou8ywxPHwr+GZ2iAGrqzygTrYjP
yO6INj6i0IwIvrpmdcF+mxuvcTkgLRpdmFiO6DS60fkdA0zyQxUFqtcsWmLT
v7cbqNjrn9M5WyCeH8QLq9mVm60n22Amvew5JrGjTwznSkGTn/Tz+L2DQWzA
QNgZWEm82UmpGcNkPnoP2pEg8n4cZzQOEKL6wKSchCHz7BII+GV0rV1nIuEp
lFNnxvbq9AwS2UHZYPnW3qEWleEoFPVkToD1W1/XGc/aPQeFxAJj0cDKIeq3
lng6Tj9aqXszjCDhmRocbKdvFoPOdJX0qJoqyf5pDqnmYFB9ISnong9HgepB
PKD8frByeZlkqbWog/U4m6s5vfC8Cdr2TfNdg8CKFr+A+MlxhFtj+zS3pktg
jj8EFR3xuxB0+elowlVh5/HF4coHYcAm30Z/gLkP23yae1NEZfApJQZ2+hX4
8J9FD6xfkJ0VkpfCmdouSnZixPBjiuX7htAPBaTtl9u0YR1bTyF2cfR0q+mt
6xpH1uA6q/dXF7p0RTp9MFQKhki493TRBnFCJP++vyqPPA5ub6ic+FLuiIdD
ps6C1uWN94EfcADFLQgI8bOf64l11hz4kPpwHm35aWDd4lZ3Lb1ZIqTyKuak
H9SsGfYicH+KLSLOpyWLMvLhm70Y71YKGmXUh7aX2KLcy/Eg5uibVQtVlBio
VarAzEvOHOCj5+oNy/IuiZynEzRAQ0ysDOaKuYeSdOOfqeIrrGmVfySvvNCI
+59hcqMk800LMgJ0bnyh1JilqrNSXqVONcguX6rF74Dzm7um0CDw7dsgsMEW
9H2EuVBboenuqyL3YhFUtKpF/G2L/d22CKkoI8V64aqPLL7Bt7jhuNY5jHYZ
wRySrBzAAgdI+nKwA5CJpgWtkEJrhpFxJG1KSbzp+gUwBYo9OPuU98dxJz8J
C5v8CkQFHCdAEqnToqvLnyei3Ax9IRnlYoSdG7MKF7fT/ZjRpPNqF3fhkB2o
2++cEJyV6sAAFNP6Sl0fRsD206e83/elsw/eCQRqgT0S6iMeOHQ93XMV8jaS
0GXT63PBwc1NTJ/I/RULx/awKUyxj8xF33/JtaTnqbgb/pjzuos6ctUSHIh1
0uVyFC6R5SzG9Pxf8DRNxpfjagGmt1WsYyawCK0tZIyGtR+RDZ9aVi8y9mtu
ckcAgMh40DiR02Laol5xBqG3Vkdd3X5eKFB+LZoQAk49BSfn/V06Ew6bi410
iwqb98INm8lk1PeCvNDOldnFf3yoHVs/Do325e1MRLkJ4gMY/CXp9sOvp59H
XekgcekmLqYK9xLKLMA7BJJKJM6Ek0ql1HdsaosSWY+jUXFPUVCEd8muHKLx
rSxzgHmppMzO/ykpQu6zlCeA9uI8RqbdS8jPyejzH3Orensq/JIF81rcTtV0
/PbL2f8wNNONUFo+AnUCa8ODdVHF4lKBY3+ymSiHUAhekA/lfA0npawqPDY8
WBbWeLQiW7tK4tLwwv7Yd2cDqY5EzCPBP4dFYyZQPpTUZjD5aXVMGW2QkDbL
JJa3J++2Lc0cNkg+F86cgE6JC7YE+rsHBOOFnliy1Pvvo0JW19ltTynPKZPj
5ovfJw/V5iYIti3YqiQFALNHiukfB4Nu7epBuhyaoMyijXZJYO2wsk2fGejD
gDJ5n8TeKcEljs3vJ4/D75hCNaEdvslAyqNFyRDNx9Hx/DU3POyPRSABR8HA
0gDPltaVrFF12mIlDcgo5TmjdySphF/HYY1+T/LjsOqc6sIexSyz4tx2O53s
SAnyH6l9TSm/SzmoQv63Su/WFVb34fXpUC1vxsEAP36+sLM+/+OjGLTS4ssO
PULKIdsk8DP/TygDYNW/YwH8IFVRy0d4hjW+ut6t/N/Cxr1qNlEepO1zt/u/
ZIgHrQUL4o0uKSblhKEIriYiOFX5jAvq02YbldL9IO+jfCMHN6SdyaiSHeFj
09EE56M5l1fFr0N5VKuHCujY1HNEjjHlAXekGij0FR5RdHzQj65s1y+adjYR
C5XL5iRlQUKJDA1RiS+fVvi4Jn1FsypKA9gymHNtEfbnOtug9T24Y4SLM6JK
OCMLPFlN97H+Zn8seus3UHxC9C2XASjr4a8i1CqT5vxYKdoOti6th7Lddb4g
uEX9D6G7AZ/Ey/GrxpEdcfeprmUXSEeLNYqdOmaH6yHkFrsA0BF8XX6APg4O
tifJzpAdGtHaxG26MJoy14hG7abCsRBPjS8iFvoCdnf9aCq6dLByizHTzt5R
0v7LI9REttdOFfdSP24cGQDQexipYKS9Y1WZFL+gkeLh4S9vBGnqYp3hzPQo
cUxtLy/5mtMMy9NtAAyoyIjNJ4ooYDX9ts3p9Z4MpY19LoEc79+6e8GpJ/cG
c7KUOSmE3mRwfW0ViCEzS36T5/Y39A3/1KV6UnaWVCtqfHwojlCwlrV9JQ+1
P3fxJ9f8ZDoWlOQOPyg7ik8yd/sZn1EQcFhtMjUjWShQeESDcH/tbUetCHiJ
rH31Zvf7NsQRP6W9glElSfg0KT6u39Rf3fKSEeQFOPP1m4ZYseD27YC6SUWp
tnBE40oK+QhJl+249LQL5CuE23cNjuLwoabyc+/EsyCbxubllglnFj+Vhlkg
2PVN6JdxW5ShOZ8Yv0Qq1xNdcG10OxGlehJByh6BvIzmDAfR+or/nL9iu30e
7CoHmiGTZILCrmeIvvQ3sk6QMCa+mPtEojAPub/Den3h8lR+7sldWajFP1Hw
pkSH4cqR8ca+Co/Qu8s+N5QoO9NLQDL1GpwSfxblSXgiYzAidb1A9Lw8WSCl
QYzWmozlowIXXwDjOlyuQtVQiJjYSecsqQDN88QYpnqtr0RaMO/heMcBOMG6
4dlN48Fc7GQI5xjVxgp0rt6j5200yLX8S+LplYo+E/k1uezFOVEH2PnD+TYU
Cnf8Kldtfqr30lPcR1yKoG9YOrVceVhGwGdXJCB5myLwWVwnATdCP4fTedt5
5Q40k3OaaEQ9WhcS2FJwu4FOPLFAx5VQnrF6CJVKIEd2UVINKvzp4iMFk5sE
w70uUqMlS1gJrW9kB/bt0nYvr+XX7tB1dDAHhT6GOvTwrsU6h8jHpNyuFe4v
cFIVTTB285HwbTDkwKCIEzKGCDuSpaSlCGA3tATnvdiQnTrEvh9ClTDUp4HZ
W9hm4Z2gAgUAcVPqNRkf/Xr9bojb52fNQirBxMmND3TAI0D914G4DElkXjME
wSLws6bm5DAT1Zc+Mxfvo3GQ3T+B9bGUaO9bpAO73UBH1Gn4tiN3McKGXKWn
81w7rNA1OkRYNvCrNfiKI5qPKxeAk6tJfOM6/SQx3QAtFa+luXebgEZHjCFn
v0vcsspipjOX4gpFt9HzUQn23wwGgWGoYwHVU3ihC217sz4Pkxb5XNKDs2GJ
tX+07jWz8peQ2xi8M2XtSXZLSIQ6hIfIAcx+ifUMBli4tbFqBUc2Y2biIeeu
qJcgnG9y02LsIqjyN97I2s3ELFbXcHGc8sFuQpUQ2+eLdyTNIXow+Jb6/lYX
0aC5UnIKA4l7ytgB0hXy7pG3J6GmaikLbgSe/a+ngPVSxgzPF4pw6MOIGZ09
M/0XPv+F5147CSk1L88sHGheCVrqGlursz53+WP6BLLFPl8I+dVBQGpnpJi+
bUNFNacxJs0dLSHUGtqarb9irqWqUfHFwDEIlbwnc2Naloo1h6DWat1b41ha
5LaAx79LeFvojt1K3N/TXBEVgpFjt2db30ohM+mZ/tOJKgpHtBdpYAtmrXAG
1ItwpM8oXBM7Kvkig6oRA7X3F8buQsgj57Ec5SlzDOp5QzdxQ31Lleml5e/S
AAD5KmRtnmqnL6YuLqrzJCIe4R19ykR9z82vpouW5sfjqWLoLhWRBuoYpnPC
wCdT7njKNDDZPlfKhimGCNPqvVQDyTyUwPsQbm1+235oF6+f0kCMDKrrE3SZ
Snoa2DLj/YR1AvMZE6Dq0rrTKvi2j/a2NCM7c0DnQ3dnrZRX+FvyCBHcS5Lh
JrtECdzf0EH7Q+g7xmIO8SO8z2fFRahOHKvln581vLbDkSuIlHJjpeZ96ygN
YrCi4xmmbSgvXkoFMDWxC1Nw8h47s7zMKhOYrXXg8lowAt0TVYkJJdAt23WM
UHfOaoIm3NkLeY8PlXyhYY2AZ9u+g9MMV4Wt+ywEQoade3MiMLCggUSVL/cW
63wPDzshjiuNFaT8193M4HUea2uS2puUqPxsb+VxE/88psuQ0kntZNSRA7JI
e76BAiK24uDxIRmLxnVge+xUwZCUfquejnU2K8xMACnq9szHiDF/+jnI/Mr7
LIk8qWfdnGScHNqJusXVfOq3Eo2hVIweVLfBZHiYm3lMTHXmfIRKLyB0TudV
AS/d0b7w4/7yTWsovCyQ3JMZrJoVCGTddYhaoWZ8DnHTqRmqB43Du+pmW5i8
L6FAwwTF/tiQstKmBZXS65i7yvyiQacBej8Haijon5W0vbCKI1kK1pwIRczV
8N84abfYrhmCISfDnozHXs2FUu5nkqI4otbo1d/FFtt1ObySMWymL0uNbPNO
Zp+XPCBj7f4pDaKnvwMQwC3ixnf3FKuAn2DbKTRYMsQVn/OryNujT4NQ7mKr
EjS6Wv+BRp5g+R2sGSxXzZaIWNvJa7axDtApcUDEbStjrVue566C/NsJ8HtD
mMjvcjKt4OQjm8TXx7E02DtPMNAQ+foO6WYAWAc0Czb+PoXeifx+v2CKiizu
OlipOTV0+Dd80dYYP4Kc4pequjR4NqvL0q7zwNqiEErnTsWXE5wfojRWZQVL
KkZtw4CbTzKcVw6ijyTHfrBe42Ng2PtqPBGzGfIKmE+5p03WwdPMJ+gCRoLR
ixTNKbciRTwI5o8pBpfqbLe/VUjrW8kQpVAenWQyYJOQLSdlwFlv4BgbeYSK
vKs9FLP1p6Jvmnv6nRDTloTl7YJJAJJD/IOdTLJL6gC0V2mURglxK1uNmfds
1gFix8PUgEc/BpO/OTEx9CcTV7IRZ9+wwgGfKRz6kAfTX37Jl6qjuB6PWXF6
YtI/nzVI1DDjpUeA2eBKPNLbcQy3kaf3OlXM7wk6ohQkJZ+9ZQsasHclqWO3
OMVtW+IbwE5UCnqsLbPaGfOoF+sw0Y74H52nUvkXt+4Y6TVyIRNNV5NmWbBP
pSc2xD5ncm2jj9udHqIZOOAL3uzxsLX3DoZMGYV27OnF1IZ9OnwY0XuJavhi
zVi8wZqSVfKHIA8Cm8yr6XwVuXNdinrJSZGE4vdwypHRPcUAG49u+WiNuSkP
iujYnO1MRf5/4TeDaG2n/SgHY3dvP92IriHNPbTuIrgpGyhOYLQMOQ62xdku
0NpbemA646alPFsIsNIVCWzdV5SkfhpAPFQjoLgfHxp6Z+fYDka6r1SuKTHb
nboKlXXmBwlGQxDFnVVLIQDCb7t3GEzzqvJk6U4xn7jlrUlA3yHW8O/gIW7D
3IPT57XZhjiOYVK8nwSDrNyvWLD2UJZc+NsFkycbuOSHyBBqQ2MKiKx1Reth
i4YnPP0XfFDjg/C8MvOyGELz+Zm+PGDUgJsIhLjwOjHJEvgTHAJ3y9YFpiVs
umqRpXXkflQXOiVEC+N6oaBoTWJTuGjw4n4pMV+cHVvFs6Bc9KVDUdo4e4c6
sxeqWnHqgxS/KGKSDPViApgcUrtkGRP5F6vktcuA1C8zsX9W4Mmwp8sUygMP
v/zsUUu4Jkp3sfJtFHKj73uyhU0jWkDbnXjYcRBnJLayO9Ki1WK1gMgjD1gq
K7ihpgU10vcdXBLQ10+IG/9iJOwGC5lxFYHRbHO1V9kZyHObrMMwx4Kk2fKW
Il6Wc6zNMh5X2YQllQYfa4fZnXiRkkWXOnnBEVMIZAINK7EI/ytuI5hJw7M3
8WQphykXn2LTC/gJahx+JxX5EheoJtIPK82Gx897TZ3PhX1Q4J0A80GOfs6/
JTrRDlLr2G1VWufqdZH2bQAFU3GxAf+Vrm/jGPkQETgdTodDuRzCn/twxNxk
Tengb9voQAwjTp1mt7CVoVnKIPvO8HaQuukz9A8jxdaLE1iZxrgyURCS5YB0
EKMZIRt3ZKdWowxY65pV/yLlyalGvO7OkmzdrFUnyY9+zNNz2auNQJCHEM0v
0W3476SemLRlc0T5vb9W+mVqk2x92AtW1tdiJ8fXAFb7a1VYMM9l4PVkMxcR
NfLpC6ZcBFgUyvWjKh/S4DrDFkKmHb7iy3aYe05LiojIqXZBYoKbz7+Ti9eE
eJpwltgwX6IKUpPFkQ423dCIHzzaSJ0N01yupsi7MZAZVSXjgQ/ujUiR2Bfk
hpUrvKt4VYSOOVEkCcn3lClj6SYRLNmR3Tvpv2SXbCXyKv4BU4YcPMkXqyhB
Xd8SdGgsXJdHjUdRklfgNlfN/sFTjleS4DySC22TAAFA1kSe0G6AcODLKzk9
NnQVMllb9wETz7r/s2hyasrvMHMrxjotn1YLoiuXVdObRfnlI/POWQ77FDNe
ITCsei0ZnL4KsLRJD92UxZN9WXS+GxIYwt0ZuKZy0rVzmCvC98R3z57cWVCc
rLZ5EZ7MdVoPSraKIcjqeWaFnZZ+RVWB0cGO4KtLgyo7ZvBj3Zt1DnDFS3O1
AlnizPz8XSZuQ2w4dc3AXDfTvzcXK6h/6TdZr0VGKI8ibzO/3FSrrkwDt7Sx
ZRXMV3zIPFxQSNU243AwL6NWTbyLa4M5dXJzXXhnvEUn5pHP3WMoprRVBrVX
MXkveHdaPhM8K73jQbddqyAABxif6AabgQfl831Ctb/WSmg3UZc20xR+68zL
N/aJ19FJge7KRQ8yr1TBR3QoQ4w9wrSGFY5coYQrHZDOSLTvfMhQ4zr636GT
G73FVraxnSbdX2HKsPrCOQho+JAKemmMAI/k2PTl+gonlwEP1W7+FpYSrIgV
RfD4ZztWXI2Pf5Zzk0xxRL5rxU1+Jsc2WYnD8EoOo4hJalk2bUrFEuy0Rm0s
id7Se+uVRg468xkQGxNBvy26mu4aCdfvY2kyQaFhXXQZ8Gi9LBMJEoVyfWP7
rt5m0iryhb8b3/l0CbQQCOUNbXS8Wz/tLJ793ssA+1CMHmjrBzawTOcT1P1y
L5mCmi88zD6iecEqEvKLbluM11RFG+HWEGSscq/IoHPOEKdZesvQoZwKSyMA
b9eTn0ZHevxkeKTGA3Z4UNpVyVOr7394prMaM1IyTvuCXQDITARDtiHIcNTC
fTgjQuKR9TIH6kzRYh6d96qHHWjFcfaa0Y+sdNCM4yE5S+NP+L+Mo56QCrc9
+pv7eqKSA7NiyG3hwTrIxP+qSl1gcG90kV+/iuiQGmIYKj7kLgrZ3H5AissY
kMHdr/Ctp7Jy18RnW3ToBShZaLieCOmRo9Q1UtUVP5HIoVJkxGnDb2inuwr5
vMPukqU3TcKQ15D6248cdWCaTaV1txz4sVWsdM00XPEUZyf3iFBnoyCzNEPH
sV7EDX+1M1xMDl9IcBWzXK2hTDPo9seYUT7og8ug9er2WsscBdfEgzCRRCg9
dI2Sv673XlPEU4mZYTd5Hwxh6iLZdWDuTj7gc7/SKWadZYQyHymdIqeW8ftc
34S2JZ1e1+qYghyrd0TE6Kk9jt38Yt99sJJJnlIb3CV5SUFcCRuYKR7TJCW9
5EBmwnmtGhtdHxHEPmsC+x+YnHErpUvFzysMHXCicF9EAmiIoB4AbfYLAblk
prYp56n8j4eVXKBWQ7v3p/+K06RWFvzcM4i9sYIvMMbW3lN2UvXe4SHY38JL
0n/6IM3nA7c5NvavM1+HK5SMDL2KGjnD1IaF2DErHF0kfPY9xjEO660YRc55
lZVA4EZCB4GXENOd5TjKcKIIVnMfGB7iaFUvmKqiwS/XGfOPwnvi9E3aMq4U
ar0EqpjrSlEi+PwNzlYEjs7MAOPu/+b+Gm6Qifcr0P/gYSJdZSUq4BUI5TZF
GZsuw74mOIgWBvwAMMXaO/nEzKeEGXkkBegArmMWH0YuAQrEqyLWY8Rcv7Le
Uagh/eGeVCUmQhKlNA5s4x6ID1VtTGWgXZNw/DQ2eizHTF2MDx6nzjOxmUTI
J0eaHyNs2IysSDemORT1/ls/h+ckgcqyx3HHkukSCYYLeLskrx7fTkNn0E07
HOFZfzdO4lZl4ZCesVfzQOQbyLZtgjVMesrIUacvbORUr4alSbHt/iBEfqL5
IhzqPSFZvdmN5kXYhoYRW6beRSKGOdDQ4SLAkMCbkh4SED84wLUS5LY/lTlH
tCxlPcSrVoOFe9BE+M7w4D9D+f1iTs0OI1VyAv2+MIRIguhCMPh+3ZCC8gXv
rzQVKQcNA4rqt/ntDg4cpi5JiyO81C49p8FRCQNPoqCH2ACWwlhuASrfsDJc
SCwg0JwQ4NtTJ8OaxZAp4f5FBwf+TyknOO7VHDxragxJAuszercf8iHPS2p6
ZOMEkek2fyOzLchAJ8285Zz2tHf91huKjwxbrC6EHQnC978sVUHCr+J0gaNY
ONucynh6C0r6PQLjKy3kUNc4ASMysjb9knK/y/HKjEgAJgAolnDdsD4qJHY0
D6bu0Bhgg0ieCjQOoNnm4AGKJRwg/MtYsb2MKauxJlwGAknXE1rQH7GNjcFI
gom6tdv0Ve0h0hMmw0atjl3mzxvv1vFOmXvCnt1OB5Ks4Le2pe2Q8SeOInsx
mU5vE9uoZNgd5g8oi9chLP7ZIQDyydcO1Ta47kBKhspeMLBfsTE3LwMreoiT
MAD+hoqtIX9jfuZfccfPJEG1J3oOcFruuBqSTyVm7wCx3Kt7WIAde4ZRrmFn
lomE7XrN3zTw64dwQFTBB/rHL7L8PvL0F5hBBtbmWQTGv/7lUQDp213+tBMI
7eg/yhXhpLL5zQn/DlNh/3xDH6LAScYs46zgsiyFK7TWH4FpcUR9tTVdTgPt
9m+v+OPw4NLFXCpOZFMYwt1UH7/jOJEz7YDtMWpEnSlRqJoldVRIY4s5vXy9
2W4vNV5XG4TKJI4jmRUmjMEgURupSwrpGqhH6QSSJNgqdKKLIm+sEFCq7ulh
Jp9GwSpdJtXCgpFM75fcwnVAD1KpsT3dfS8lgiPYgBrzGHTNXuuFQCPUQiMW
baxjGv6FTGMTezAYubgAn9+IXzMhim7ds3tiQSpt3x1cuWFQXvUSEYOMYjvM
aqc0HAdT5xsqxxVAuZtKmtFVLmxeNEueRRgswwJa79rklqfWhKcjuPGjg2wB
chGSV+8v4xQDWpfHzDZ0bXdYqXvQb29mNH7Zv2NXOkhejk3lQJ1hF38OKAV/
lWDAjR1UAgmffR0ehdEl2nOl5TWi51nnArwoWuB7jehzI5ESfh6Ii05Pt+B8
oAFrBzSg4B8BpAi6VzKj+07yNQTLQdAkUtDDTGAPXDLrF9wfqwGV3baVKiMk
7hvp3A3lbjwWL8NK7DYceiZaXulMAgbOBv3SqsFutHDSbRPcTSs7n89Snnij
eVSfSy0SL0egfUeP9qHp9EN/CVBoA+rxKA+29/Bp2O3wppTUMdFtcodPITqp
9xanimssRhRMsF4z2hZN+2GAQiJ2aS0VA6yuhXLy4upI/6yn7KdxEQMObY7s
MK8gnzV2dbY84twOR9crONigAXLtgKn5OTassH8tUUN3LFd3qCwwWZk+WmlB
XfoFo2l34TjUnhXmqTpR/e4BQWXXCTLdJVQOSuM2zo5rd7lZ8ZF7tbO9qpdd
ko1f2ipRMMRYC37VfuEzKlclqjJB51dC9fdTe9WYjRJ5nIxCVhJbPbT7nmfJ
leiinfNGjrbPYz405qtiIp6sjuiyDOcF8lNB14Av6mvxgBT3TLkKFZy7PxPi
8Lg7B9xyfD0xTyPQBBRaSJoYXiaLJ6k0caotbZTm8oGaUpm6nfGOOpTVa6N3
4dWF+Rjb2KwzJtMzOagx4oqB10HqSG1qK/nM6aQZdta+lyu3xitJpWu7dq+U
bA+b7I2G+pUokGbGEJHJ9ZMle6J42YzdyAq+SiyFu1togsmX13x29PhjOHnm
UJ+UJjBle0f+FPibbixSPuXmuvSr7WxOhERs3z071miWHXFZfzSvrYHf+dP3
o6EsBuJkHdUhSK4NLHzKdPTGRMPgFpsThOFOe9JZKMqRGgvOK/FOOWsqq8UM
wgO9anhr6BivelQA7VQqwC94t3mTuVe4SGaJURPbr2lYThvI5/L+pumPqJ1E
Q9O4mf5m9lW4IHq6lW0HFWfyZdnilesComVM38koJMvZgvfW8YSZ5rvkSZ21
huj/rng4GGbepSo3ok+m58YX8aB0GKP03bqzIvTHAJhkguTu7LO6MaBRiPHT
cufMA9r3NiQ31Q2My9qitcf6bZlYd4m0B60w/RkydD6g+c85ZocaIngJRrgd
qMEM882+xM2SpWZM9XLRV27fwaXO1NYDd93/dQp9KscZ+U6zpUWYp/zbd4e8
q+phjzIOVQwV+7KcEwFNHMi4q6x89ONnGDXhbmkMUbW6gpePqK8Dy1aix7Oi
PG1r8YRnnd/Dne3Gibr6R3OnHhIqaH8hZMlJ6Zgbl5dvR12njkHgy/nGtEoV
EzPyGANtb6XWtDJyylTZ7m98py5HF8z1V7dawSx9n6PUeMxLksTXURR+Xd6a
nzcTy/Ii/WVKktaEkoMh9b7UqN2IP91974WHz7luMNuDY6qcfKcWxPLxtjHV
FAIVjaLf6YlizAidifrDNbievxO2JU2HUq+JuTPp76R9S2McKA1l/YWJ3yC2
v11U+cDko/lP5q3gM/YDMV1yaMUJu4sfx4Ctb09oSjzqWreFlDESIQ8x3RA+
YlL9KnuG1WF7xpiPadJGMsS12ND1X/rKYks6l8ZWyZrPfwXgCj/L0QTgcOFL
ehuwHZGBaKxmVyymCkzpqt2ERCJGVr1hNPD7lhgXHh0ulHzpyhfej4PTAZa2
njMMMtr8ue2ILvlPk1Myt5ojET/w7IF2O1yrTnYsP78zm/qktLqyhIFvSV1I
UtUUZJDPHfr7YBR/IBeH6jpJdZdOLPBMrqOswpWrTDFctHMvktG+JYcL5XjV
Y7kf8kTNOAGK5SpXgVcMMNgxZ34tqj3L5GXNIZtSxSfrGEgZTYCl9oOAV+ci
yZm2r+lxgXkfPWR3D+SFnjCtXOGkXsi7lkPcTHukUC/+nPgTFFtkeLD/1Rp5
vRB+N/TJnBg5eA5qlHmcuV1ebs53sciKrS44B/H9xw8jAP6t82VueJMU9NZM
w2ZANrAvN3AEn6Q9jq5DwxHeH6aWaf/39+Wt/SbfXSx6HyFn6I0vS2RNESn3
cQz0yqVHSvdYFRRq1TEyTf0el5qnMFPLnjIbdoK48a1KL8hELEh+2uO+CYFI
O6dyW/J2LHCMXLJbDsIKR5DHNee9E3l7tYojgjspqNdb2RBBBuO8cVAGAKWD
fLdNE8E3CaBwEoCVHCLLtfWTqAElRTCevwoBFh5SG75ikfmJjVjZLrIBHRCs
/IXUISptRgPqbHfoobr295dC2e7iv20JLUJTWuYAhq+v1emCTKuah0IZBWQM
xu5loAgJZXMaMOW82AQQQbcLxHKK77APnq8egTY2nqBGm9zX3cydaCWsF3mk
vddCiuFFyWrxYAAILY9zShST3YcNATT8AB6kubp0vHaR9GyLc2eRlThVeqyd
ghAvSWMdkk+G2j11+cmDH/mCKppYxU7eELhxbwIgOXwFd8LZ24iDGcp8szjC
lYC6xMbSiNcprfA1jtuiCQV+tJeP/4lGZpmfcs9vUC7snV1oOLHNcr2akguj
/vrQV3h13TZ6NoRq+TtxA+uBO9Izu9Q0nMsmEJ/iR/Buq10MDoZ3VoVZuzrS
PLh364jG5SNG0WNKJfDYavW8gf0IO4EUUA6r/lcT2U3J1o9kIJCW9dDnSk+d
EmLSzmjCLZM6sd0QZehLTEOwIYIOPLKyMcNXK8bY8mJ9SqY83exg+cJdbjkO
dfZIi9MgJZyzhpiFD1RNp9bHCtLH/XWf2asSYz89vYvJMGyu6aXLuyPDhQul
a6whQVziNoL0KfmT18QHl4fuWmKhBruu8iGBAQipiXPPNZO2gqR49/UQHIyV
dz2T1luRpK3uXxZxIlznRcpvkFl72L1/7PlVDQ6TyYVjx93rM1qSX/an8Dhe
FqcmiOo69awVJV2JgaVWnIsI3nKoSTeWpg2dkU0RX32Ra+h2qwt33rIvZ2qJ
akM3qvTF6YiW5FmYfXTORTU1H7D+mWJok5+lHbnpMtPMUoSJH4yJv5AAeuGT
2/HPuQOOHaOHo1Wbce/mwoNPzwIBKCT250y2OSlYS8W5JiKtL9RaIHgVe0tD
v4UTkP9Sr83OQA2CXmh2oMMjtW+R6EHP4iXOoDu6xoJIhT1KauLVcWtJBb01
E9kFbTXxXr1EhewwTNJevENPp8MCu8jEEEJohPBwEncxsIE2TpxHAW0hGO7P
hBLr0Q4DETo5EUVorhioaGT7UBslQH/vfP62fdoWr4gI4xmf8FSt1b7upssO
Un4ubK8Bm3/puRJ5VOGripHkXQ0D9q4x+hPfipKWZx/fEFrezuFAZVr1tHHX
8+su7+CdFU+KZQNFANnOCf5l4mBXvu0tyCEq4X1/n2bWSByNUjNhdGIh6kwZ
i3nvcJct/7vkk2pFK/UmoUe/RVx8ckTvZ0AQybs4Cz6dWYNhjkfusJa+wGpz
rDVWHgCsVYqaW5NG+WMh4RK4tUkE6lKOgPXf2qTbOCJR39e5qsj3F1KLMUle
jCmxY2aLqwkFgVqRqGAebxJ4C/pMc9lkyCU/4Adug0xyfbHxSgI5VKhIDlrg
+Ns07mttPLkdsUuYI9fcCYG06IQGnpQpM/SgdnLOeac831mVSHqufJFcBNH7
CpTkVDEDdOyps/ChbwrT0OXFs66MVwtzH5z6TkqAJUojwmW2JpYFK2BCwYq/
y7LrbeMaglk9hhYj7SEGICpFpTEZ7ZhC/PkX8VxO1w/399UO2uOuwd2pCewb
hkon19OyBqK9M/qCn3Ew9a6IwPc3DFWFSE+IxSec68W2H/ijRzxoEtm4z/l7
0vploQ/1f3Xkn+EprTwcC/0pGGDey3e5vWrruFVOX9rmnlmHdVLY8yDhHVHL
a8ogjuSIc05B7TAQirX6yl4MsMAt/8mbfEXZRqYucDDnjrE/2+D5lrALgDkw
dmuyfsaa0ifK3F22oZJhBaD99PZwB1o6+9qrfl+z9t5bht7m1Y7o2YevJzLJ
uJive108/JoR57NiHD+e/e/Lq9mzbY8aknJ4PGVB4Eoanj/F4U2UewOW9iuR
pBh+J7i1RvyJNQwS4SCu/XM932G2xXdwuvaXpktU/5PIpl+yiCB+/fLzdjmX
XCPyxDXA+lq9HFG1Hnkletib+g8YtUK2iq2v6XPYqesevTIu9E8mCSI92t28
FRNUeLS0clTRLUaWEyCfvaNEn7Ei+PBcnIwXaDnIV+772GHiS2xqAN2/89DE
hWG8JBWOdiyQq/VkgPfvCKpYfEJkc80gQMGlk7U+a0hnaIcjuy714yF9446g
fTBxkeHP8hBJrQPs+4EJ0kmK9Wo7vNwCusOq1AlbBuRwCYX1Ma2DcqC7YmaM
NQnFhvrszvtdA0yvXk3BIe3EL8/+WdKpKdOOvcy+Et2KZrR+U/v2Uh3+gh8j
IqvawbulT4riXyHC5TRqFp7snLuH2Lmn6vALR5dDiaZchd/QRyjHYhI13nSN
YkM824Qf6l2HzyPUU0+AqLzW2Gq8yQrlq7sW5yg1EFWOr7WAlOs75SA3qVM7
9jhvs+ZLY6NfozDG1t/IEpHAStfJTqZCxUprWe4ZX11zU8BOY+lAeYa2z5R+
+9Au0wRq+2LfGpZkw6BFHlnZJgRDsqvhEHwjRmZqUAs4lTbQCFIlJNIxroPE
SyVcElMHGFGb7omfJPpHszwY9adbQzZUys/jlpN946etXOTDDb1uHvb4MDgb
nBIxeVlQanqfJ/pUhf/6bgDrXceZd+1StB8xn5vVbt4p8ap8yHWqLpIHtwa9
3g2S7xk1X7T72lqXvsdvlzKZT5YhyQ1quVX22j2ePVuNv4yPIU/Ab6VrUE7T
5ZNMr3tjbzgHi1ydZKVInZr3Ltn2GBTkbEJe9N4v/fA0bcP7SYoZdcveFZgL
of42DZeB7IqKrQTOqdD8M/Ibk9SDo7lKQsNBXkGduJJk/8PZ7hmxvOONCfEd
Tqnwu06y0IkXUby9s5t3Sf1rIJwd3pF6izMhjGRYZFSPWujPmOQOhlT8EivB
GuLYBwy9Fy4ah2hOjqniafbUEx92iZkpyx9HJOeeH4ARJxB/RPukYQrM13iD
BF5pB6D9OonA7Zlx2QbRG+Y0NAzDdb1nHzWgzcYpaSO63IE84yW2PK0U8tmG
RgoMJnDthGiSsJAWGDzbd6shvc2mPQcvP+KIrAlp53W5FuarVwFUGy4pkvUx
DVSjPr2cNGCtxu/6nQJslYuEm9wnwCgiJ1GjYNOKKwIRdj+Et/1uCPGX7i7s
iIydhQcVCX+urDODB3/fmvH3pEyZvSEgzgYcWdVcriGTJUAt7w50iG5eAvDd
YXWHpjEV8ya1P4ZD+WIGR927IpwSDBoSxOzNd93n86oenFEqFKY7gcsPJ7c0
5sJB6op3ip7vPPYO/nsCm4RJuBoYj0TZ9BkyE4K2tn1YmeneY2TdFZqq4I6X
Da/C0ZNu7AyUApLImgMyQiD2adwJhMg7iI/KJDZ4itGS1aub5DFzTs15vOEl
xkZR4a2Vw8HNx/chTr+dloyMCuNz7czQVkQoBOpwo+rNfEnKBC9/H0yFtaGt
mGCkNXekBdjGsl/mgImb3liPAUAX6YiQVR1hkL4447tRLqnFVCra0TewaIvJ
k+TlUbk9BU2874u8GcqVyaZ32sXCAmxY/vw07tq+wzOGp5a9aMplp20RD7Ap
vEwQQoA+uhQ7RlkyS+H4mJGWT4bWNvlS8lpm9Da7qMRdJ3YR+7m9qx6kOYh/
b7vDlGO9QKnsDsLqq7Z/lY5xsDvoztEL/NbpFovT1xwnI5UpPEMBA3Ic22Q8
qB5YX5wY4U1Qc55/BTgvaS3/S4j06oMZJsauPDi+kZJG+Uq1GMIBgffkjh77
4tcPj6RYYvly4U7B6hx3mITBR8n9F13fmRtIgx0TpCUtN62oyIls/oS8KirH
3ez2QhrFh+bm372EfcRX6dVPC1tpzdaJoOsfNndPKDdFaU1wKdknqZWu9sta
gT0qDjo6I+TCPlj4LHR77epcW4Xe8ZxXBb+aP3hg9iylkdZyiwqWayJ5O6iI
L0Tde0lrY5hyc469baw5VXCo9QEE+mGlcgdC08vo+53VxX3oO1fA8GUJrqqU
TzfaqOXY4C71+o7TcRZhmF9bTfKIZecL+ozdoHYEtJN8cc4gjYaZ7Df30dbo
5ynwX0d5LJEZcYTpr3XtuhdYx+UA3fEu1/1d9IxJmwvXUY2k4UqcHqlwyerp
aSSzk+OmZk2OBunuWF44gbHjDna+gwXXy9aQJ7/t8hgOJJIxfurP2r/L91vF
KjJFIU6qyH16qswdDaCt2IUkGstvgdVbjK2ILNS0hxEZkai9qB46MGAmqLGT
GJP+ramwSgTfGuHzmGjSmMrhwz76HsfUZJpQjdKUVHX8E137wScnfcHUMd/i
wVOqzQytT+3Z58t/9oHpjQv5+MxBjRkTLMc27kAWJTMU+LnPlTbQSBzuOB2T
nxt1CSXOgy7mIk6fE3+LuTGan2RGtFtmTtHMtY8haJsZeqiCygMjHfA8sLvf
vb/PTYNCtG4/5KcfquwgjBTgzgIXbZg8NMB+98LYj6iScjrBSeznvW8N/0yt
MfKuFo62c7lCVjYjzsjt4ofcIU/g9zGd4pLbqKZL4b89TYAR1PN1uEKmJ4sX
MtnqACdSyqbA9ATmfbi/pVzddHdfWOZggP6Gygr7vl+cFgk5gooCLHoP+vdA
FLPDNECQ51DWbmxpQNXenyD/V2qsS+E5SFkYQzP7fEaASAXpsQAzKg1t3BuE
Mx67Q8vM58DmiN/MgsPO8RTG9e5r0GdFFbgUBIkipxl0NLv3qWQEiItS0E84
4gn6C9go8WoumPwi9YhuFArq8OTNzPIE5Uk52wxmcm1vtn5aw9plpJ/aWRBB
RWARCIYm1dxZEqw8X84rXmq4zXnoYoiLQwpnrrq9JAJGtzX1sTcPkllf1/hi
RmSOHQ1uIvsFNw5i/edCxVI6TSIqRsQdIM/XrydYWSFHJIOLqfj/LkXdpkmL
2Y0GmdqDwBWCQelpF2InMhhnOGMuLHF/Mr34xlte6wmCK7jXBvkC7tdkvClM
bHv99lPgnZzX8C8H61H0ipelIy9FoNfEffO3wR++o+trevkk5K2+CJPytggV
wMy6w6CyJuY4jR724vmh1vjU+ALWkeYvndwpBdj2xRp2t0z5hRT/UQ5WBNqB
ya8F76NyKerhdETdGvyWUrN4H5LV2hHWHt4OVBJDuqgANmVxfz6yeGuOS0bE
n2nxmfaVatoIq+9D9EhhefB/OzZdjzlw4LZ5+m9Lw13CIpGboCgOQ17tmfWw
C9AUYz85tC8oXEo9SPn74XfbQEWTpHezKWMTs/koIYflIJqOx1IcA6vcDOnd
Dfja5gTUI8lTu3bgNsPF7g3FdOdTaZ6IgEPiJ9ku6YrKm0dSZf8AwVouUPD0
gM7BVSvyY+J841MPwJXHndVukmK+U2kIVFQMZ7dnV/bH7vXKUOKRnlIkV/1Y
DmvWdmcWSxklQga/KfT3hC9vbIUwcs2Ak5KjSiYwqr0ushgmej9dLd7K3nQC
GQ9bfY722uM/k/hnWB6Le8czM1HOX1v+q9635IJK+9919oZrNQp98Mq/oKDn
mBasoZbYpshr4nbKD66I14sgjpDARHNo08hY75/T9hXmDsfrzXu2aFKIjSCD
90rVWrFEXrt5TYAn2HaDdb6vJA8+50+1DNf83oi0l55Gms6OJSIfJhppNNuO
RG+r09bgyA/LawW18x1Ygl/drSa9sHGhNTvj+jfHJAc087LxL71YUIdDPZOL
rmps0bFyKPmUWORPYYlTC5YFQsEW2ZSLblERHr5L/PyiMngbgvXKYgd7YuFS
210nuYccUCVOC4tGh/NWD5mKq8XrwCkk7WGLg9NYefn/umh/qKXodF8ZI40Q
kRpOPnbb9g3HLgrX6Pa0O9QReNz2IwIzk4iS2+L/Ri9tdwlYoLIK5jF7FVz4
/w6/341llFwD7tnPGjML3OVXO8YxoML1IxlgfYDwqE0awnZB59DH/QcIlvxw
JFaz9vKY9P9wW3ipqDvX1on68p8aHlAo655PN0jsMvA/jgL9WL9bdu8HR+uG
9yWo6RSdCpJY1NhZpI4iaJ/z2ec214sT7LVlq/WMbmVhRByCqhBEDpkrqweq
I7Xm8G0OZuWp3jeGwAB/tYUaE+xLh3n70E5N1w6YlgmI84N75tFGMsT/9xd+
v553xOfSj0/PURe9D3bf+4yCSjjIitakriBaUtLHwh/08auS0bLTmJvI1+1d
k1z3+IvDxnFVwxk6QfXvSI8FV3DMQvZ/LQ9D7In4jnahCIwMc9VtoeEEcO7b
OKeAjbMYH7+cW/5I+HeYKgGLDsrm2tfRExmk6tyL5IAQT4rvVOCaIecnQpRF
3/EPDAbNWRqdP1HGOsphnylVOiUFoxnWOoLZgfkEWCx3B3V3ennbaTHla9r/
HpKNraub49H6BFf3kckBZs085tBYXygj29190+cYoZ6qYoM1cc7ULbgQVp3G
UcbOMh9X9qPsMXhrWI/czj7e1v6AxoBY4fLfCGn3+6jaE7hmnkq2uXfAUWVa
IcJYHNJ39Tst74353S9h5afx95BhUAr2NGcz3i436ymaLomEOuuunPbgHdhx
em5T4fYlkKFiRWAEt8I435mMIt+NLqmGW8vVPpMu1mkNL9au9qNpNd8zXU2I
vEMD6bEGDhKnQdkxcqJq+pQzDWd7tqeoZsp6QWUi0kQTZvFZ6gbzWjE6Naoe
PpYhyqaarKu6Iu6QhOjDL9REEaLp5HDoXS8hZlRPOtNIgI0LKWCNxaP8RboJ
NuA3oJKMwS5KNr9r2DCYpiZWjJ7Y6eUVtx4w+2hHDrPzVg/YxLzn80iGoIdt
Uoh/kVO8jX4YpZcr6nZIfU7isP7fLVMSexMdKySjrGITq8orC7rxpEmTwmlE
uDrOvFRJZ15g8XbBq8cmWbUZdChg9X3g1AFAtIKCKStcBiRen4S5g8TzPH7h
u3N1QEk0eidPHEYB3sP1wEo+UyzUTbkiiIDltK8z+6H4SB7Dr69B05A5xeNs
vjH+pzmPP1gKLPtTZVG1zlB7tgrEpRpVN+Ymg4QttnAH5PimLtGUDdKC9iHp
gwFZGReWq2Ztp09iOxFhHlCYJ4IDtKvn+iSKdSPAU4At4TkyY6SwOtcUpFVQ
p2HnU9HRq/LXvDReicV3lGqcFH9537BNdBPwLV4GYbJjCe315zM7YpaXPZfn
yjEnDojR1T3OT+9TC6pC6D9/Fc1gf9YFtlZ8GJYOVvksEiY5mEwFUeLOBDxw
zAb8mWzze7feP/82PgZlsML18w6DzC0mwLZwpZot5j141e/cE6rtHt3Bw4kO
u8vZeM1QZtXukoWcWTka+f38D2vB2EQ0bq72Bph6stQ7jlK8iCNjqsT2o1QN
0Y8jBXi3PVqkyBa8OZ8cJri/bYhsQnju5SKcYOmiFiEpEieQZyISHEiZDO/7
LTEvBMf0ZE2uzIyxvagG5vWpd0MMSG7aQv7OqyJy0EXAGSyP/6sY6o5nkjqj
bnJFHnPacB1LYFmSStuqdjN81V/fWUbQi8mJ3MNNBR4cQg4hS3U05pk81KHR
rn+jA20RT2yPUG3fIMlD/9IRM6IwAt9q1tbTrbt6fFJhm/m968V4TH/+I7BG
PKubBYFzE+oMzRhtBibFSUmEeqV9ymgSHnUrIi7bPGKiy0yONhjRPNCsX1d3
Pi6MgSmjiEaMkyPoZnCknmWMLhMukTSyA6jBrZKFsh3ddZP9DMrdcVb4q+IT
fm2cYSfIyMZgSHN1z3lgzJBNgN91/ZoT5HuP6AFzZvKrbZB9yXaVSZnjT34+
zbSUlQeWpZ1DUumXoqGMcUcCobHR5EnhS2DWg7gKsF1ArwP2LcEUXcKJPFvM
Ra3PuyQtjSMVkm6dImaFHCny4Q3b8EL0X/5poYb7PlfLZ49vD4lJyRKuNRbj
0krX0GkCr8Dy+m2j1VmAznz5NUCUvVwseyhoED/9yk43E/o89HhULITa1yts
SFnrtuuTBxM3Bkotegx/MrmsH6lG/tTUwI87YB5y9z2AxW0s6wYdftgcR+7M
BunlgbkpNrITLwClNiN/oYedBInZ7eyCN/RZzQ0Kj0mgWnkvLhTuBcB993Mc
S8hjQ853rDKG3rmw/QpKAOAfvs7zszOtSlKOWuiaAY8hqPUPt/b88G1muxmh
JiC4+qbM9BAml9UwDxQCBOz685UhNi5aNfA5rFq6Cqm86pdTQLSm5GVKNk6u
9sdH9ZB4OtXZ7fvjPLmg6C6uZqqucBixaev84nxCUChv+0Jf+3ZGtfTtLNrS
k9BlrZ3ba/6l+WoOaX978O4EFsraTXnboTbOQwuL6uuK8Z3J452UGuFMkrrt
bZWsOEsJLb09itwHvCLmKg3ateSlTP8Saw635P1btut0XWbFQiLh4qYveFqX
WP+6AkpCyCqC9JRuDmhm86XcPM/E+enWeSI7kQzGvzRe/FnhE2WAcYQ2CUnC
aC18IpnGfpgTbEfCzll28hYTYpZhvJRviPnpFDf7Mw8ojokezyA1MKhpvgtb
hkzhYrrAR4COcLcffnuajJ9NW0Hgv+SpYpQSkRDaUK6gdw97+kzKJG0b0vTE
DBoUbckOadefsQolTYWhQEpCdug8fA8TQdt5hDh/9LMH4DRl9STTjJ9xtWNz
N8EyekiAkqbHAahugxtW8uB3S6j8By+qaj6TU5fnYqkrjWN6RlmPs1Ts8PK8
QJapO6SgluYbU5WjEnWMAgb7GVasjChPhjwXPDKGewXgpYxVrt1VMDhXE/nJ
hw87gRU49VI7CENGJqf6Bl37yIOpMx1+R/6c78SpNq6OjXTDJd2kraP9yIum
0i+AuhBK/Yt1ARYxqWs0Vg2VtAtpg31Gw0cRI3dMOekps6hAyACQ3FqcxnHQ
mNrjdcBg96pY7g3h24PqivEIHfmo/8wnzpIYYO7vwcPBFlTVDX1ZpzDrJRjw
9RM1QzzOu53MghqPoZ/KddVPCIaN24oxIj4fxkOMM3Izm7mo1N1yYdq3/ry3
v9SNuehWf1uFZzbtHL0Kw/YbMpyb/Sfi06PBDFbWv/Nq9ziaPwoK57jLqPl2
8ZkU/9HcMGdb186IUad2jlI3YizrxP3DUUeGnTJ/tau1W4nIFJNJQRgq/Z9a
OqO6UcMQ1SB/2FFwqCSmz3C2UjyNYB7DON0rl/NfkTKSJdvr86Slw8yQsqqC
K8jz1ECxHSEn7nqiyBZYIabxX/PVlzUjjalrihGtuJBFNkbdybXatBwxIuf4
RX9XICES6AYvCjIdN0+jAsCSdpA634MwjMyQQccD9UFTy5Nc+LZNQiJsXUyr
xU5VcBBdSc5+ORIDhyt01m5txR5ZIjmISKcbCNKr9C+72saSD4b70k44y9u0
Rvt0JDsbDlDjqJVKflLePE+ZY3O3YqgmwsJmZsEz2J7LLqgmB0iQICHdpmJg
tEx7Qm1gfT3hUBAppSsJq7SfcAnXH7XVdWwmJ9FFNDEHIgNvXJKI9MYi0k2z
YzlREcyeuFtM6l1a6SayGeMH6vu7V3nGyaxVfq63m1fNxZntjiyOp2DVBDmy
nGoFiPx6BKkHLJpUmqZm9y+hleOjiFN7DXNEhFSdZ37XmrK5NaX7x9FaMhLo
me7uo+EwYYh48smKkSHMLWmbAAOBX67gFlauJ29mfiFsP2uWg+0c30O6NlWo
Rb0uOMt8iv51pepAJrW9anzk1KjbEvaAqc00lYn1JkpBffO4uKn8+/ekarcc
rHDwq1k7GzG+kQzcTe141NJ6Tg1wWjyC2+cqXN6WKqgBoiIa8K3Cir70/bqA
y1Yg2CNqOoIoTDbe1PxYr7RSAikX4CzKAik2mWFp3QU3oFjr9nUcnfpqwU48
zc2qpZbuxL8ntKbhMTPPKwzcda+xaVZ3vWG+WyiHvbJAvobzc16UdZRCDfx9
1ezC8d/ZqTRLZ8k7ApAMRfcruwCo/tw/zL4bWYaXZO2DPIOQuagDW0BXYg6s
BgtLuKrf2IG02x8EdRemK+ILUhDxLhyZAmErQ4P2bczFxS5gvWRmF4jZno5F
ICT5nGZzLB5JFBuF2Yzx0l6dGFuS7ohx9itODojIOA9zkTXAOsAOQork3v+L
kUHesUwJfLe4jh4IUCtaghvSTSlJxI2C3BXE+YcMJD19sI759dx3I9jfqQQ8
HnnDVAwzaIYs6bQjvWR6PRVFBP9Xf5ck+Squr8izPmq5yW97YrKUBv0HVwxC
98xrQK4Rb30e5zrbnibdxUkRSZdaJgjggSUFtqixam5QjbwB5gAWxPltuKY0
JBJIcFMdAS8UsYZzdPjSxhb7LQuPbp73X+XMg7qVgICETc7sfKCbrU4oyUkC
hdg0zcwA5z9NDJZ5O46LSg+4yL9Ng1kRJ+KeXPW/uhYhoferq2jMSOfulDd8
Y1VMejPtpwalc4AhDyt+2CzAaDfie/ulUpq3A1zowQ8izJhjDJrHyo2wOKbG
UeLJDlG+uzAPPqqL2asgkgzq3nC+Ax0I2mYq59F+6NXkDYgxx54xpFXb9WO7
VTvdGQ+I5Zozn+HfZRSlCgQ7B3pee6obuwzx1dd9dC3Dnm0PwEj/hDLeIBHQ
8vZj+yFsGOGZzZHmIWeWii2G7n6aSZ5UXJukS+vIKjrm7qyFo3KY4DDyb+ke
FIxisGqDWuvW9GMWFS3yL5Qqyh7Wx5nubATt23aCwDGf5LkXTxvd1+qvBbTf
sb5eIo0iYJQSVle0llSoxPh7FL55rV9WGNvuyn50MDUqK/CmlpQBF5f3J2ac
MIqrLcRNgACsDdQBwXwELtgb3Dr8dg4MWG0mXsuakl+q+RVGRW1AIAJ1Ay/N
TJ3zavPL160ttcs7pWt1QYkys4vlK89Kb1xYqRh+WdYdpl/icyvnjsPk/PYd
eJh2qwLXXRrYp700YB4+J0P7Gf2vfcKhNggB+PFzdsRRxCzsS5uYg0kbpTwu
A6ZRmqFrY3GOGRDGBhi9sEjeCMzPcx11fBkwa/GRQnkpExQHXos/1tm55EjJ
kKNfm8bXJt/RUgXB4KTAnwcN+rGxSF8mTB7JJ7jqOoSnBe7slIlkYYiroFhL
EfMRsfCdGzybF1jLOq7Bii+gE20arBkdVU6pkq2sZOfZOQ8r1AKSaLjhEuBU
YeBwpWNLlfzoySPicf00tfA4adxUikauSi3g7N9m/CjI6lE9SLSFqcH3/kjJ
TscjWP4q/SuvVngVSTb/y9NGeiMAXstqu9zgRD/1SSIMpFpdEPeEn0q/eVEq
Ymh8EPULXbQYTj7KLKAZmYl2dnbynF161LFM7GOzX3ojoTwgPJSYmCT6FEez
7PObtrWV9gWNLN9P5Ec4rPZWHVE5wrqL2yTCblfJXR1R8BgYATwBheH90ezZ
g9GHoXn0PRMMf6/IAM+HxBzgd92SaitIrT23QCKS7BFzVFNHoN5mE3eG3hjY
ux8h1kpvi17wl9lPc9ohoZXyO/8ZhM5nw08MzPac2/a1MKhKfBueDKz3DwcZ
w4fJeWRrRYPoXFQJ4bp+dCQs7fun+0A5lqosRCUnwUQ1MFVAxCtzbKNJxEQM
0c2Q8tpJwnmqiQYORmYO/lA9lR7UizjgvNuftDQ0Cm7q38yNBSmZMU8FdDah
EBelaGeZFmMrMAOq/lOUXX4EGuP8StvE3MJNOuq9hDgeIkew+yIegZo98bvv
UYwhwpG0PNcDgdbGIsapzZyltmij5em7pilrZrMCgW0H5G30inNvOOGTKB5A
cSumAgqI8VbQ+mJ2M0gsp5R1DxkJVy9ac51chF0j20gIKCKTBzxJM92tt9dd
O9n4tNar3KULO3BKlsJUYxnqKsEQoreZN4eM4Ts9s17KJ9RMgT/NxwFfex/B
Uh1k+cI8fRDdjxcpd7024RpQHb6a3GaVXdF930UpnVUF9PG8fUWuXSXOtqJ2
6rT2A40bYAyx7tLIhevdLlM9eA/6on6ywiH8OQj3pqJaDLvOeqR1wAKvEIPz
mUDZpl9kRJ1V3rCuV3Zfp4E2998o4eqBDrbFCJETlmYXcpBwyfsExmYANU0i
BMf1HywOr/WL3Dr81dmZhoAzH0fZoKu9ZHEr8Ee03ugsommvqcRLxo0khJXa
gkxkGhhvFYanrqE+KbYlVLOD4sw2JUY1oOXDLI5p1P3fqOm4FxRq5LP/1KbW
jhexqFc6hh/0aCdZJCGSBCFGgFqhwfAFXt/HLYHLWR1iPcGnOvCqwok96Mbo
AJfjOSxg3EP3azjogtnE2mjI3xPuvGIhc2kmdlqMFhX7ENI6vqCwboXvixm1
TKN2FSm7RwLC8MVvpTYx8htTz9fUX3pP02aySfITyWcM/2guBC1k3S6tubzh
m305WVnMqdj+hpl+YYQWyIdjOgODDIGz7LHw/FSR15DMlukrtcJC8lAncFk5
WWEluP5da1aXcWr6L7B6z1qjuD4mByz2/eiDAThJMVzAd20QSzZAy8oUe2kS
uRfjx+oR2pp9yobtZpAvAo7A3C0zIYCJoZtISDQjFhWRqlYGGcg+ZJ2KVJzC
r26lvGjOXg3Z0bd2keO9vweEMYj8I7ZaLUugprep48byX0uctUbm3ls+v77Q
dn1KqrxUCTbtok9NojkpRAxfgUD1/DooIWRXAvwgLTp2iw26sCRFk0hDfb1/
y+V8l8ALKOIuBzEOmdkzGglsbAGHry6eAWxC7ks1+FhMZArF2QA7MZGVvI2x
DStZ8Wjy5gagcpHsXxKkCzcECyEku5fTna44b1SmIyeXm9OPXYiTHglEpKNV
peG0bKIBwDtw4IRU2TEROcVXKHQbu4J4uZ07hkgaf0VO602rKkV4IcZbA1eA
q5KY6j+h1DsQJBJJxr2dLpPuOy5EFafv3qf6eLG/jztpslpFeUem6jq501S7
cccXw7395gqwxU0/c4SfmnTatripfjFrHooRoKY3kcjeoEfWMQFMkr8lvfve
ku9q1vdQ8IJRblL86ywdS6XF2W07L8he33n2VQMvgZvOPOswnuJecUaWaa6h
rBwquAFN/lwvzEeH2EH3z+jg71khRmPogq3AdzLU/1u8G6dUTX64qL/Hld4S
TDIYzTWQWp+/8auYbbQWJ+pxvHj6o2AyftuGsLwLgmAiEUT91hPk5sPFjtER
eguz21YbPQdUadi9/n1B8EUn388U0ahAD/uikBslUVKpk0u6XlSi9AenRgOT
ndlzUObM0B92a8lw60twE+BzWh8RZP859QCZXT1pD4pGg3YsNcmTtutC1Y/p
Nex2Or//1oFDL0yISjO/1pDxrztZ/w6W1KglZdEInL2EVpIeygqIvziMql/E
ZEu6BK2ewKbqSy19lL5Ps1OcgRXgws4x8ZaxPrQVPfQ9d036lBTa4aX5HrSy
r+fmKECOSGOteV8oUOQmNt+/bNy84kkkt4Dat4G466xwyneHtQAiYfJ4xlwb
qcEx1kY+zLtFWsaIGZFF0/7KOMPELi+13fIup6H7GkyanBNs9n3QMJ3m+9DE
NQLQMPuFYVRhrHwzhm/Jegvbzlui7MNKDhf5aXmnSvztvDBwnfmP+bqgyo6b
049OC3KwqhID0XSOB3QHZFZfenp/+bcxxhBpjhHE3aa5Yp9EV8ApbM56c9au
OClgf82yha9cCeoSueeOozYQWgYXz+TmgpvHLAThYHBpAJVGOf+yCuzDWBV5
4M7wA+ZcwHAzva1KEkH80iuU1pZdA8FE+QVhk+WHnUjYEVFcPVonM8W69p/M
ameZRv1m8Zq4XJTTxmeoK0T4uEcARe6jNwnuGEOS3jDgMcjV4Bjf8kS6K/QR
HUpVhTPy6AAK64Hy0XONbcRZaJFdxvZJETVpA27+rWDuvniht7LmF7LxqXWj
L/JuKCJNPyb8LdqDhfc5pwGUf5nIiGzm/hYvQ3HUBAl9oFDREC7q9NYxPsNr
/HT+M8TRaqo3FM0bfynjXOuXF3qTmQ+v5OPrmWide3/50er4+Hwer7hJVoJe
F79qXhsEnp7v1vHS2T0/whgfyBn7jLJEpJZFyWlnWFXsulePJ5sszz10jiU6
wlRVqr3gbf9J3PUWZdMjB1LFLin6m7UWYO6YSWxTCi6ytjg6NzalpPZydH/e
j8GGY71MAyc6NVxWYfWTA4vqgmT4QvIeX5Gm3F+TrwbYXvG9EIgRYnzXQQU7
jUieMRgz6tvPiobzHt/W1nkEjoRwWPLvnMfUHidy+ixL5ohKgLdc+JvQWaWK
COmUmtEX21NcE/Y0UUHmJ0GiAy1tEvSCpk4Ca67zzfhdWjzIgzA8zL5yAv46
1cy2fPeYZBFIWpq8JHpqWOpvuvhox2z9WIyB0+Hh82aHSEUioh7qjJg6OGCo
CUpIjGcDfhgsC8fURb9nMNo3Zbp4FoM6h3yjAZivN/JY+OrzM7uhrvAxJaZB
axmtD9MfeUK5s8BqBVeN+ioGTw9MY0RkTEu03O/I2SnuD2M7EiFo3Nn0MYpq
5TdMasVhs4gec27rDbBbfitOaucIL54TyT9XEbot9k63ZiZj64tCiTNOHqAl
PdTQP2ELcmBVDOecHQqltLazc/WcvPr9YyxLLu1fXRa3iF3NJMGBTE6dkeXM
410aGaJ6U4CyhKVP7XyhNrXlGxoJkytLXriu/qjPHF+EvZQvmI7HPF4vf2DZ
KPcxm6ZqQp/+h4lmDrIOCR285Aw0z4a0pNYniBJgEA7Re970SU1Gul1LcQD9
eOfHICRp9RWThmlqxu430HxJhpnKyBrUvYvneIy5CUbZkw3OlGxx2r4onudU
tZy+VOeLRVN3Kuj3vxq7TV4tIoR0FVscMYlQD+ONA1BcvbMjzCqPwVwADZYy
syplLykzBPiriWX6mGoOWJR5jVoRhZKNyCfv5xBlNsB3SjJjk9yOPUeue8Ws
z5CD1TnWg7Bh+w6Cd1k3g0cL8HNjW8xAXOClrCOUeUX6yVqs0S5bCK9+bUV1
f/9R0TCb9aCVSLIyCRLgy+Sy2T06PW0zgrJIJCipkWP9NNWBZ+Ur+d3voXMK
tX1fnnqNV0XekGkxymU/fxO1CUPK/KelvXkpFQi3aWSJ/2ItWpwrFDOnn9n+
oL/f+iIquAFRlk4yGkVB0OOxzgEkNPklYoqEE/FX+r1ECqDeC4FBgvvpot/q
yzAW97E2vGZlK5bHHzBt/IJ8xmdAF6L/SzblIdo/QgfOnpFg7hPqyYAo4eJ8
NVDfG/LBu00hTyg75//b/vtDoAVHVILJ6HnZG+jmLJLPsVLV1Jp31mB2Yhf1
JGMnCNv//RL0oT+VPjBPDs0sdHJu4Uh5R+V8zX/T9VulMPtfm4veSnMceLQw
nEuCDsjbvfCwz5OGFqAspwsurqoBA5qbhIkQWOe4yqf9EGeYWVenCI/Tr7jB
7/D2rOT5qEkgQcsY+GcWJEvE8THMop3AXtvEyUBpm/aOa+Bpr4O8dOSHHOcW
saIM4PqKgJQQ/a+4+Uy93bNsWGPtJUW4kIkhOpIocnzb7cycm2eYvYp3ryjU
kjyECeuYTZxGShPr5TxJ8D8UcY3LtFkpfm4wF6sHm8kwuvT2IcyTQeR+boeC
2Qs7J9DLHyjXPgLbebYk8zJbrTZs+KUiAuSN5YZfwv2cR7NP819BZnfdV0v1
3Fl9A4nxRvOE4pHIJQFfsXM+658N2XMqLxT3IDJam5WqhT7wRZise/92zNXG
Qmc2W5rdpVdadMjM2uS7RuGgCrL7MWovPMR6DtFiPeBc0dvl9dMfbgHD8rv+
vXOjTgY3YSBAdngNNLvd8AdXthN4iK1z+Z5HnUDxjl4aAdYUfKEh/M7aBden
uK8TYvm5HGZ0F8WNtaJq3BcXDgXiDxucyf2X0SRQvvVjm1nO9JDziPyIvUKD
QXVc2GT4LMeAxNVubbmzs6yZveFV0SMXy5n/gRmeTm0Y8Ll0pnZEZ5mTRHo3
rVLt8pIeabvFkz5C5R33PscPfYKDBqWqkQK6QpGUxhA10uzcpiVPXlb4wEG0
YlThTsvlbFHgaZao/qmT9KX7m6mDyEmQK3wAtqGLVY9zDLao5OUekvv6npD6
PRhJbN0DsCJu6O38+wcqcEnjx0m5hcZtW9SfTkvSq2+y+Kz/MsVFhE9vWWhd
egOdDgC5wwDPESfZXbN0dTBK9S/Ap48ajMXAjcS8DM2VEzCS2C/O1Ush3rcO
yjcqycXIdQFjiL+UkfHZrg+D6DHATATvsna2uq+cNWdeRAsp99S/GLVU30qP
Q1nfUqRUqJbfKPVzvQQPcB4nwr7zrJ9Km7SSw/m+jiBEqqiaadBVxBCFwi8k
wFn/GHO1w3Tkw7mb/il6AueBZ5OmHOT/0TAA1KPtCxLPXKuDbAU1YOE5i2pB
3dXc0Z/eT1216rtER5jwSPQJLM5msyhJJvSoH0RA+d9wgCoPJdrLr12kJTSg
T/bl/RfyiinYIKb7B2czT2NRCdcPelgRJO1SpUI3JfG6livjB4OnDB9ic4iz
S2qCnqPlYNsp4W4ybIKkS03iWwSY2nDYwMhccrQONOpP9hZTFC4ZB8gKhtab
kewxQcs2cYU/NXDb4jnSvGFG5Gbsge8yZgvKoFdOjO4cb0KA7Z+HfoAkxMdt
fdvvNFGOWv+AK+XBGwcLurRVvX4ydFuZ7Sdawq3+/eUVIuXeTqP5WJd1Lgne
PadSXrysOKKhY4iPczBLjGr9NlgSv9jkHilvEf7aqpC9Y0VqnedbwQqzqInQ
a6YS3TjPx4XylufOyvTbG15XVKR7oz0piCWf90+6J9zzxhZGLGAuJy9kH1uc
GMPvk+JePoJqDyWFU9QMMNdlrqIi6TJDmNqhkn+Vw9xe+Gm5Wo+N9d78oIq4
wLsLW4KE/1YlBZBidsIzlfd1f4RvPtolk3uuq6QXmRP9ZC8sGUjUu+f8ZLW+
9N4NcWYvw+P5OQLFgmvGNrE8DpHAJhVMYstyzadCKswhS05tlZHN4czYGwFD
9NTOMWR7m5qozLku6ajc0XuHDlsDrG589VQbIRrm8oS5bcaA/2LQOfm6HXZd
UoDU3Emv10HXmthH1CJ322CXximiuTayi6sQ0wwsLAG/pzIuIpae0kxy0R+e
llryqw4LLemSaZ8er2pdF+xysSa0t8FsScxRxKauBWZKl3UIzZg1U2NDn16j
a8n1yLbBHy0OJ1MNIqyqNJYmkCgzfiFOFtTrY7WItkJRQlXF3I5K4QUBXDeq
6zxo0Np+LsnhKnDkeGWoj/IMdTW3fIrE5NK7xSW37q3Sy3fVOcqPChsOP9nH
CAtlEbxRDW5ziGWqWClkntIuR5QAn3Pc2KWqnXL7v4MN2tcubuu9mg1iU7wg
W7oxtG4MBs7SnJoM94qc5oePYhyjxf1lcL+yZEQX7AULLgUj5e+lbe+aVMnG
BN6F9alcUzW9LlFZaAHnk45ADkKp1IsGzwZthH5Cqntl1N4ITn/L+nR/1fX3
Vgh4jDjD7kVYTIsMX7CWyPuW8ELoM+S5glKbPAzXbiXScVkEGJFjmRwb8vX2
aySLUXs+sOfPFlBHdvoWNTidl/vkw61zl9vdpeDXKNlnuwfGxBDJCtDP3S53
RgTI4tuX+XZIWI9EPwLCtdaFwzPwQ+0JTYfyoTnEOY7SEZb3E/1Vi4lQnLTx
6XjwdhDytCKUHCz8zMjQkX8cGEDeZGcvnYBNPSxwKQDEKeslUfnk8ktgVNxQ
VFz72ThDWVth1vrB+jHcRvOGlaNNgjXMcsm5MMBrh7o2g/HfMTodLN2u660A
NE4KNxUhzbGoFtB7fag+3CIeir4R33eKKYbnqkKz0S+tTXafuOyt6XBvqdpx
rSAR8NV5H7cdOGyzqPNnMWCGIJZr4nZYMnwri9DTy5W2HZrVhQ5m2dEX9nMV
3rff9S8yIHNpluFvaxVZZpB8fgXMfSp74zAchgtA2O3kH70N9RLJdhIX3ped
Y3vEpfjUByO7g8lAuS3xhHyC30AX4naPaVkSGG/zkqdtrN3bJ4cXgDPUfZT+
4S3J0Osos1XDx5+CujJoX20CA45I6mHD7UyG4Zd/vXVD8mgwul00cj1UcVrQ
ogrdCdDqXfLuqDBmLqwtsBYpvBncXpXc2f6QsYUj3voa8NbG20XZCYg90XHv
YONnhIrzHGyu8oQ9ZX619DjK6lBPK31dwUOTtRB5CIhpLYNN4Txw7YHLjcOL
qnQ7hcIlkgfYE2QOtqSJaXYV8NeEi0Nbb1ZX4jDZ2XNK+x3XQGkobN+3ECPg
0MpT9cAja2dpV3rv+fht8G0ztR6zMaff+nRN5tUCDEoR8aTCkVJ5tayiC5wL
a2+VGnB2cYROan7hkWKzqcUHae3L0e0TC9+0DpzEO7SzAu0UGtgZFUN4qhdE
wkCKd6S3vZB3cUXjB5qLVzosdjl3qis+8y0ggiY6zmmK/lZFEcKrrTqKRfuF
7FW6F2tYXXNr9De5Ty1HYCU4gs9pVFDpTPDHPk6NzgSkp8Q/6lcieYOtw3Gd
8zskJ7IoWxz459N5NuXfpCbA/5GUHTuaZ/wpt6C+kW5vvWkNf1nTfJNiKuj1
tOK67lp7eUfOIfEaJsImGr9zMNlbSOaB0+lNQnHguAfNsMXPBJeiaSWYvE1P
JE2PgGfY0PKGJC+LVO1dXDT7mHH+qKUhk+KwEZlZrWx2BF55LLcac1xywrwI
nX1O/JhkR/9ApczHiuNtbZTaQIQbsG3IcixLDpDwgCNuG8W79Zc/VcSSy7OP
Stopuyhnpl3Tg4E6b6BHyG+t1fPUpJREhaPZurdi7BDPIoGn3emLqZBfmVNl
3LEGhCsxuNXGf81fkLh4J2Y3RXqGG/PPyAk5Nj8ajA3iGUFL5gbmNRKvjDTT
eYD/XK6R15RpdeQW4wLo6xhCnzaaOu9GAMW7P3BLkNJLf2SjKNMeg4JkJAEB
eEyy+5TKGnEI3oJM6en+PIVvbwBPtjv49NV+miUuDMLdMrFKdA/QjDJPFi2p
9l52yG9LPdwUYU9RA8tWGqh67/mpWCfs6PLerxr2fw3A02p8KNZ3nXMhwVgh
f4MEwstq3+rJCX2V5h7xqQPhqIl5JBIM1IJhR8I04DblUTibmTAuuNr7g3C8
gZCQ9/WSDSqrHjLKPYIw/1ev/9sZbQJ2i+zAHJAWOlf9y5SOhwuobcanBn5y
gXdYtRpsK5EIiEYwRjS3H9CBW8iZp0SPteCpeuPXQMENlED0AJ85iUJyvyg6
pz0iqY2+zQpZxdSPd400ehqlSpdboDv/OpTxdBpMiRIZSzfdvz+wIP8YCmjc
yVxpDe9vqyHVoAjFehV5v78I7xLWSdvalH+5G/ZeqYQKkRSWL82QMTGf3gyT
6CxEP81qIEahQNDZADUazoybFW1nRg9vBz7kN6Sx08RiwnxQGQZxu4w2I3bA
bf6rjSO5inAg45CeGgBippovPgRjF+w/P76fcvZ+ZGwkJ/N3i9HweT+vzl61
HjXPcIQaB85DxcJG6cIl1bFodjWs8auWuKe3k3eukkOIVyUDgfhOrAt19Fpz
xHgC0XmIbgdWI/HRn1hx6pMAFGd1VNZsiW38AB+7jksUnqWIR2v0IZZESdjt
wURJPiajayrnT8Zol7jSUB5sx+7LC5CdB+diLO8tW7+Wh6BuJ4nzPryN/abG
/WjPMPXPkowegBU+lLFjrKwbdnMJecBjQEy4+FIJsE5GTGTpTkF45zh6v9nR
DS1GgwOHzsufBVM871EUEPr9xB15ckWVa01FtsyCVzQAEqYISv++4rhHgQim
jzS4vHVFznKvAod/U4ODHdhuT0kd4yI1KnLv0jLqLcAdgnihUiA3O44jc+2U
VJ10eKJo90AoX8ArFuE/x9aDX/g1HlPR9VshLIApS/YZixg/D3U4pnArnuRK
JGmrU2oE84iCr6CqP/oJJV9wHTOnpHsbT+vc14Sm+N0OT/xEte6qKiKKyTLQ
eVyRuv96eAlsrdbZDlgB0AzkIoHW1z0dVgmgj0k6tbyalojdJ8SrupDB1NU1
53x6RNG6LXVWMHw/G/kBNEIMknlzWBcBEJjjIQWVhODk6qDO2anEmaxXyxTD
eKjFNoDcKWqUnobcptmgUuXFEZOYHRRjUjjbMio6YgLOd+YDLmapu0mfJmCy
bgH++okW0wCDv1l5gAzWKnm6dLVnOwAXcdQV1HRc6vgN+EFlIGSe53L/9/55
DfgNBiBm6+11X2IWLhpzQyp65pknegjXGrQzeSlfYlfJzaS8AjX8Z3m078sv
+/dlOn0/CCBtpHAwU19SmMLJeHBoVHNiDwuklCtjxQd90bYtqSJ5gbeik2RN
1VMbu+zarol322Vpnu7JIn60u/a/GkK9mvd5Qdt5SttulRu10ou1aAmlqNv8
MrA5rpQ47IYPpyttebU6cTElawYqJ4XYITRDtSyfe8imUlPugLEck+uMWvTu
aWuA/z+3OLVEePlzdLhYyHBg5hH3ESVtmfAP0Tmy4zZNEZE1arzPXKSFKsyd
pl5LsRnFtHbyxptcnDhdwk5XsLgQhzQ3Ayk3cuM6iKV5J2kUeExR3MGdDiPT
JvtsAxABiTet4wgcKpxvfhMxJmZf65Kfv9mVmOd6NpfGx7nSa3dynNigC+AG
dD2cF3VF3cxAHQXFhiv50oCIwYTuJPSKBDz4wDmM9A6V+BmEW+wX6QiLPlvd
4CdP3ja0QBCwM3pEVz3BYsm+MUB60sg9xvMCAsUZjMocwyq9ormJPFtBz3Y8
rBrQ3lZUOyA01CytC+04AOJA8ApZcU1IYJpkMXIXLbZpGRp+43EmCvewKUKy
4GkOTuUMcJgc3gcIAChv+t7jXU9tRz1MZp6T3jSw50xIl4LgHl5zcDfA3AS4
riwVLOPRv5e9X4Q0m+bzIHtAc1ezpQzyn7HViaj6aQTIwEtmK14W4W4H7cQh
X4xHRifex+NDZCkenLaca2C5azSltJ9qWUxq8IxBJz2Yxc0rd8ghAP8H0yQK
6zhWsp2lrKMNT5jL5XK7KSmlzFRZtgFQ1/kjrrkGjp0b0u9ZpURcWOxCac2R
tEAu4DGWAbbjQURW9DvIpKIPMDAKXVj1hpD1N8Q2B8OIWiBgnOOSMi+7f41m
zeSVfbxlhO25Ek5l9r0Qfc1QNR6aLXASMHFyGo6Wb7p8lgljzuMSmh7IqQnC
sC1KexjMdYNL6JemxcNKQy6tfRFcN5uG2m2pV9M/M9Aw4/8MqE0KaOaTOyxe
rmZ+g4MQ4ESt6XNEJG+po5hMqz+dcDPiXjlcLjBIWyd2uu/apsx5GhsW93Qv
TD9TpdgtRh45aCmt4xFq47b2IKAe10lsAQ6XnPRQCXMmqUr/oBiMq4WQ63a+
o6VAn/o/Nza74OrKwXN8bWj8t9u0+NUHBAUb1xvL88LrcyhRlI3+1wHhTzWW
ugCdXJJDmFx6E4Tuo4xtd79H3iCae3UDWFR6g4NFDYuXU5w6F6h9NwMltHWu
i74hNvW6N7VZgqTGZoln6poWy7jtACx+K5WabMyVVM66TYn+mDMLsHsGmaca
sOlnaNlINBLlN4KPTlP1NxAiN56tyMbPmFkmEKncinjFGh09urUsYQ+UfyzK
+QoPkYl1zRSg+EIX0rfcrD4ravZAATv+VL+VUglBiMRcBWrzHgxuVPMF+9tK
BGn9o9IhrW37pdluJds0hVJcyHxq8fMpKX6S61wl6gFQ8BdI0vo9/b+0ePjI
sHCPy+8Xrm5VQMkWW1lEH4wZzJVMbDLL8JB4M1zB8o39BjXdM+tPi+AyGroD
uRscxEqZAcUgSzfcHWK1KUCquyqdyyJ/JQPTJlWBHx0k6N82Ee8NtiUqqS1G
BVN0K6tvBPZ6JlK+a1RNKsyQ5AwatzJX7yqSJ8UWFwhnOFjb2znxgaTt1tOm
jI7/ONzdmrnJC350bczO8u53ntWmDwQc7E03efnVQnn70clYTEdnkuMZmWd2
wOMD1CPbu8gN5yq0tKtgA21pcjZz2WCobU2T2M0RtQs+HDsQj8JznPyoFT+N
6ONRrlnwBIDGde6yHu4DcwXDKQpVJUDTsC1w2wJWNqDMSCXeC+VWuVZwWZ53
IBuOjdKaj2bSPqJtU13x5Wd/1QNBfWNfqCuA4g4QqbHgZr9pTXCdc1IKGlKk
cq+LQwGSyQjP3MndPSrqhrCkpEWIOrJ0qDnhKWqFFeQK7pNmCRtpJDGA/RbZ
Bh+SZC+n+IyAO79hh6yvMbk0ORosVVPNqI7XjDeaLgnRjwtTxXf1cDh5mDn/
UBD9JRfff2o+UvOrmWDQw8U6rlit9bv2EqtKm1iTLR8awH6ePItcfBnPucqb
z5h7w7Xkf/Im0Wwq3/3Gt9u8zN6REZCMp2Ri0nDKZ5R2gps9h6Q2U9DYztNh
wEgYcbkMr4Ioe3NqsGoIdKRPCz12Bf+6S41qx6uF3ViJQyUSkagPAKv7jxh0
5vH4EHvBpaEF/vcWqXQ6VrrR9KZCRf0eJmZJOzMcCZwtzpuWQHZ/VZza3h+R
rzH9WJJZajV3BLWDM3A2cfLYJRgI98YBPyhn5JzfOPoFQCGJb8VuvrWT7UPV
Oh9e97fYi6/V9mkHTTqYCkc05fdodukyBfDjsW4QVVBDXj4ohjwjGa44DCxY
+AU0Up9y0Gt0XEIc+urXIXowMHL1sRv18dPaVmc6pt/9Sretb1HSFFMf/YQ8
SfrzCLU3NsTIgpPfspFT2fLJ35F2HS/UTIj2BMvQJNlmYH3sfKklM+sGT2Wk
wqKOYWpUkrx2oMZOimc5yanGf2fGKIdnREl9SlynePhe2lbXQF76RUYGrmCy
fC7EbFR/jYFb16LwrszRLBNdf2V2QZ/HVk7/dDo91gSzWBUmaOqHdRNVg4BE
aKMVNnK0v/PstwQygZrSffu9ma5pJfcu5/J+Rb90D4x77cgqkp7qG61VlS1N
AuVdHN88GjJG91Y1Jlmc76jG/WYf2aacCOCCYbMHKoW4+XRA1T8lCeST7lzd
OTOT8gnJ9kaX3+9iaby7iQ+jdx2v227X01FLItihEnR/eIBwOqafBsciiK0y
a0FyKeHYkgbM4VL76Dd/SPwpf3tKUKPQ2slmGBDwQcDV4+egDLV6FiByPnWv
LSz0uM9D5A+Jojg2iXZDVYJewjpPrquNAuk52LcmVX04doZs0MEfsjWxBdmM
5IQL83gKAIHksvtwpW+5UzrkWrYnCRWXmpNbnnaPeUwJvb1OFZVYTpms/att
vtP+Zoew0tkPvcDeLvRB2M2nvXSJRb3Q1VIsF/qDO31v3lrdPRGIbEd1c+lp
b/ilztNoKauxupo7AY/SmaWORVnMHA6LquD0t/uExndZ7/a7s/rUYTgOqlvp
ninVFtIb18t3BqXmSymU4SLxwXmVJK2o6BY/Ynnz9RnEEn9PnaNDPwniMl55
DPjoEQLFRYoXnbkYXLyrMZkO5MFthdHxZSUe/ehyzA60mo7eSZNc38IDo1rL
ghLm6I2i/eV0k/hJDemcx6oJVkOWoVanWXZD0uIuxvLRLbsyHsm2sqle1Iyi
FKowHlNKIDzxVwYhyScojDuJPQqF28libXBBwqc9sFm8/29y/0wVUAZFTKZd
u6EGUq3khKA8WHtRjmleUCMhDQlmNQx3dzveMVmof1wrikyF2uPEcbgJeep8
tu0vJ+YGVxr5DQ0N7COKQpeQUa76Yzr3XrU9+u5w8ERouLujDfu6bu9ifM33
BgoQxCtN7diFNIFQQhQMIDPex9pPwqKdQqJXj45eYWZN3ouH6bJxqXehi8fm
B2zsQXm3+fyYh7qMpCa3VD0luAUgz8DJp7airb9jmwb64ESr6RBy79Hrh+77
pCN3rfL9J4RT3Mdt2hbrgN7Tqm/jbENwd8qhoHVOEbV9eGqmMQrX2Uz0nGrK
gurc9LSfeHYevO0/NDfV9ImdtooVrOwdoZxou93qtdrxSag3vbXX5ck9+5Cw
+TvjzDXIrQZZN2iL45CFHDoxbHXXCTR5Hje3u5ccN4CvaKYTf4M1SnHrw5NC
+FWik/8TGrq6GXFTBw7DlhknmVCWCaS4MbE/OzGidrKA2TXKzpHA9kFGcaUi
0ltmh3v/DcDf8UT9dDotC31kelsWfK0zo6m75LyyBimOPjNtEFxdEFvrToON
jcszS15F3CRXO85CUP+K/HfLapH0nN6Tttm6hl5/1LQRt0gYb1yOU1W7rByI
Eq7No1iQUlHzn1u6zaEdLzPWAzBhclawiH9sCN6vFIU0eH4LbaHAbB9xSka2
MDqRGpkbQuESE3j4TG1J3ammfADrLKw2xXUzSaYkUciGokIEYM7Cl0uEXsEN
6om/PFic64XgfPATFIg6R2w7gjWP2mq5bWZ+uMFcEIiVCIqmdIz223u9EOv2
vuri46xHoM0gRSxwsvb9XPtGdGQapoaoGnto5xQcFcGUluk+BPGmgA2NkGwv
2IAKy3VKURCnnHK3PfKXpbHvPdw912TuMogjAn10Q3po8V+oQE0Vvmda+P2y
U9QYuR1CKqcafGBigL8aKPT0nikDqHf7DOntX7ZbfyKA3RUQP4E763mho8dh
nPUNS6GWtRSKoS7xKfvCxmH77fmQQlOtP2/OmdoxGJycmlz7WlImC09bZ39A
/om1LUhsEZVvr7XSjLFbg/rHgNxZoyOLtpSqAbkFWSS47HJRYS1m6vfwtkD8
3ERUHTtOgFelgg+LFruKrSN287F0mDagU+y+Qv57OWZUw79MOrZQzgkDMFVN
yQqCzQnLw0WkwM5I6X/itKbV+ANMpDs8BI1vhB+vhfaQ0T2pLjM/t/+c1RPW
LTcK7Dc+tFGirEfIRRUe9b6m7c9eUx9MAJnWH4OlnoHaFf+qKRxt+v8RpqKc
hPQdh/CncPNMmPPSu/j2a4Dvu5uqbqojXIegR6cDo3ogovykXkAWZOZvFZe9
G3aQQ7D7ento1klb9b2QGY8ObhioeknOX+MvO/exPjlA4EB7bgmkVKsLLXh4
u/jHogMEfXyqKA273+WitXcBnhyssXsFTwk/nGQLmOsICp5I4wiJxkP7wt/m
5C/VB9qf8lMTMMFJv+YyzfQyja6NNT9Ob1IZl5ZzMHD5rah+voU5eCCCbbvJ
ZROlthRHxOl9okh2g1qeGRvWR6hcu2YJ/cos9Lz2VcWZN0aGAc+5me+reO2B
u42ztUY6atNL8xdkxnSpytEE2goaUI+Xr11d6V0O2BrHFhJoqUZjPV+MEQer
rNGB2vBFFXl1Iy+W5fudrObh+mwRr9PEl3buXYzmpDbcG8zRJRIUShCGAOPb
+gVuom1YSrLZFQV7u0Y/WmPQ7/XDU3URyQGKEaaA6/ZCZMjui2svHysSzKWk
xMpWtb4ess0ciBL52TKEawrj0d3PH5FJS9NisTuxKmGrrh2dvGuIkQ4zQIKD
Hri8jpg3xEYIQg5e+NLQAYu+KmRU9cIl3ItmCzAvRZGKki4s/FGxJPfbli5n
331ND0yqh6pnK0j4gbV/j4ADH/qJ4zJ5hX2lA6mJNyaSV3Pa7obGGMOj2AT9
9RUEnxqkHH/ULyQpZdc/hgtQRU/VzgyoXtbz89T/FeCRxV2jJd5etoToDUr+
ZysArJvhpSJe12/kXGIdCiQWHa5xd8EAkK1XbfAxUjnMPlEXRVDqUOSV7TKm
OEG29SmiHTgWbzmYf40CObWpern4CTwT6I5yjT/5ZALv7QDZiOzPpEbWxAEN
z23JDzF2YXqTAUuuDgbpGKQKWqOfQB9O+4TtAYP8y9px3snu3/oPmETKjR+w
XXXrW7jBa0gpugkfog7wDlduEPLQ0MwPYurC0a3qwjoFAWhoJGf905jESzYl
/qIlqZBnroFkMk/zL9nP02e2cPG7jiuQK/HBu8CC3GQJhUnNBRy4LjItz4mg
xyLCQHXWGpIo03qKua/F5Kg9rQrrTBQ71smmGyOHDy7ZA/khTxqgHPotLplA
gVkGKMaiC59B/UoCtYcs+eBWUYCY1EDJPWp7+aake4gTkDfLsnzYSjZ1PQC5
xBGtgS914e0sL4vk5rbjKGNPoygC3yXrBr6atNn+Lu5SRMHSASwOu6Pdlrvc
GCZ2kEvAqfB8lg6gBp5ZN3Khx53vr4y+hBDBdyGBSK5+Vta8AREPyq7vZi5m
Lge5gu4QoyuHEhxPI6aFOmhuDRllpVRvxi3ZCsUt1PtyM5CFjfxddtuXBO/f
NDXLc0tZtFcm7o1bMSt6VM0iLPXs3bjx0r9qTzIC0AKA1DUfttM1qC9PNsx6
An/vSxjqjH2VEDyq/1nXqMSLeD66SK8lyCiu6Kuq2cke6VXfq6zayYID7DBO
EIWGoSFRH4HIFW1YEWglJETr0P9rg1JFErwax5JBrEih6iKIFVIRX+Dokc+n
4U4eYaj8LLvYgwusyqx/8qJj61XUZzkGa2FkLlYOxue1vOm59sc4a+IMZ6Do
fhOWuCEvVa5qc8jTnKfuaZ8P1f2FlQF46WxwDAdoUAwd+leJe0okcYVEjKIL
VnAs+hge+nya1yaah74kzZ2Jc5hcMQiv8o88o1ZN6R76sszexpVsi4Ah9BKj
7HCa7UJUFJIXFPsc/11RWz3uiwAPwfPYdsfPuOMdDfzG5smQN3Qsv5YOg0qw
ArRS5EgE6BlFLvnMml7IwK17rkkC4sobmwb3o6ntQWwRH6ShDhZVfQ2QbCUY
5DuBgSTksAE0WXV/I8qVq0zyPF7LQ+rQFqjsgC/pgPyOTS1nrDbhrARtxDDo
PnZwsCNcgmMXwFSdlTNlo2w+IO9TxFGvNmIX0tJlHgRB1divMI1WmtdWNs0m
MF2GuLQxDbe9xvPGqCjQHX5yHduhoFndKpxjzBi1m+zJlR4JzF27xSFZlMzP
Tgeq+K77kvIl0fRiOy7yFPuQYz7bfpbLRkrTP+8pTcOvcOB2rDty7O0f0yfV
1guvH6XMpXF04+/Stvgk6TlTQM1nGgnA5jd03p1WFLAcO0/ek6XOatiSEduB
Q2ecrygAsSQpLVt5gPnZEbHyKtJVOw9YYWEJQmdM8Q6JxxPbUN4YFdXZ9vrf
pM5w0MdtfFtb3C9XcPZMrMrvhap7IFz3u7HRQq488jMUDn3dMUgQp3uiWHTJ
ZHCPRCBXY1amO6w04nMHgNvOySaGA+Cd3Y3TWGJ64dcAjDDsoABFKoWjuYw6
sXZ09e8EvI5w0FRS9bBFRQotiYzN5v54Ow8Ns73tTdWFjGe6wd8rCRXCyPUo
4IHOp9Jv3zFa6cN1WMon2Hn8sMpbA1WHFJ03ccVB5aDYa8AYQHcDw9iDGdvO
gbqPshDgln23S8Ib2kfxLgAlZWd2LBi5rOlvDKH3XXHHfm8B6ifarnj5XRgx
OPoRyI5h46Agit0UCqe9aaRnktb5nRJbQyVM981xhzdHQ3qP/tmZApT/B9h5
tCD7sA7BtRoIKiM4TcDvISxfuhWgj8M15KkaUUwde0xl2BPiNDGyYZMXVQWj
lbki8AFII87dnsmzXuSVOufJa7yYIJWlTwf/F3S8+rrMb9hCKXwKXEevQ2ET
ukexOi/xx7zy1T9mQI+WgPHDAql36UwMqj6Fl1HkgcorQx51DffgqojvrZcv
Hp0RF+n0ncFllanp2PWOqXmn8m+C49/JEQUPpR4cM3LY8GhFKglTnYTnKlgy
VGW3Z5HPWHntLtUxWtDlP4Td12uDZ/z6FLO8Z2Kyt4T3g51wDauKOn336JsZ
Sv1Q8AuOJi9+3DrXXMWZhNwRA9FkpER8b2672CFaUoc9xlHGSdF/ZWA5ibj1
0dS0Eu4A+0+/T5H3SoDUo3ZX3nEr51Mzat0rwKDK2L7JEa2d6CT+YBQ8iArX
AHnSjph8x6sQFWX+Z17HkV2Pe8jC4X8IyiEB8KMhWo5fBFawIz4njN+LqcRk
JFOHm0opnEfG6Kaer7mS79b2ZakAriDl2+5IKMyp7x+6llzntBQyWcxxIbQk
fMgSxwjybIvY7MIdBEZVKWP4qshAF/SSgixxynuCHdOM6IoQLt/h+P9AYVPI
ti0BgR3uU6CJTlIMTQfDvdxzp9T0NIN9T2ZE1amtZch1lxCxZe4WxyPH3c3N
zCsPDfhxk0fE1b24riyctjmcc7iLBugN+4Q+9SM6/P9+4B1iacbb6rWBK+Ix
/Ye9e48CUj5cv08lh8ni79nf51PxFs/FTJjFNNjFtNF1Zjz1iZDmCF3HLKvW
OpEM/lNaI6mpsGVviXL+6ES4N99gg+BYRJY/8B5WtvNb+/bPMJdwwWOsXFA0
xfA1wyzVav6J5UQbiTPa07uzmqH3LlqdqF3pPI5cc5clhGHgCEc+CL6VI7sI
A8Ak694pAMmecJ5qcq4EXVdeyfK1Pm2o9b7MfPd10Won+73iNorV8/1fIDLE
W7XaGPVBIiM1Ict2saPV54hfLcXPEpoNB2wz4+haaoSLRCaXLg1mWVKF/g7c
k3nHj7jy6O0HSdH7lgH56nAtr1O9Q6SXxCV+54D50PAxtTdDpJ1srBV8oVq2
DYsK9xuXkyOT3pEXUPPsBwoAqA2Zt955/a/uHA3zQFh/ccFOXNyLQVgSc4f4
HF33nAlUlbMIYq2+ldcb5KIsmv8LawBXB/thBmRjEIphFPgK7hXQT1JexUeQ
XMSN13Qw1JZ/4k/U0ZwKYil6KQbARpeRbrgrdcXp1eIvsJcqhKUrzX3AIdCF
5f85hd6rHpJVa3oel7W2EbhsW+rSuXzlckwmH0BwPs6InFC8vLahI72sdVY+
tpo4WSK2vMfPDJ5dNSKSBA/i2VGtvHxa6vLH8A6AFZdBc+CmcA5oApNLhQP4
7ILxjp7Be1mxJi4dVVzX1s7PKIR5i5mYDNYhWsb1RpAmP8dmKV3e1Z4D28wF
cu7NEgM0m1f4jlHhSuWWHoAwkBG0WmYkbzq9pDrDAUtz/l8uJHH3TcS3X3ob
HHakEwqedz1OKHZxgOcvtU5NCxFjBs2GQm3D3XS4w4NwmKhkivFmYM+1zwOu
1XvL2cACdAB2SvknMpKkK+SNFs7VyyhgKZhKpeiRNLW07FNvx2TZvPy8qLpu
GMt1FwvhIc1AAjENg5bn2JYKNCt0nvKrj8FAIhXsrfhUdnvl8U2XDfAPmFx6
HFuzAoQC9eTwuNrlGSXK3asDBjEHGGYSO2ACAu3NjwTKOWfr5SHB2zYcjl85
H3ay0YK0+65y2PlhJ27+xThPM6SPYyVL0kEYufOpcL+rC1VhOnpuoqBFR4qi
1ieJpuwu73ShOMO7JODBfEylvmTm8QIP/w3aA5hIBivwCKAEn6ushjcfJuj3
php+E7iRFib0VtiVUGBhngWJF0OxAj2+asipwcfbh1ciMTrCpC8516J6/JHu
VF/QEnkXCosADV/2bk0afG5JcDcBvTjXT2Z2f4vqgxz7MQDVSnklDBwFEZ8h
7z7lajxgPi+n5aTaPFpoNgIkb8Neqolc2GxltVQNfDQJ+JNVkDbUn4ocl9BQ
7mL2XGQUGBEuV4TNBPbN4+VaZmLQrQ0+5WgQNXWGmZJqHIUPe+kbbGX3l2LJ
9EDQJ+Al7tmFeRyzauskqCibWJB0MzjAMSMRHzINSnVREJr3ltxrzBnZWjM8
iIEbpWDuZhfNtAVTyG3Bj1RWT0zmVgxrrvUfH/YDK7YwthnmieQNb3gaVoLC
Q/tkLWtowoEnoMo9rnWDRWJ7ONQ211ktM21wKBIWTPv4Reoo1xwBM9nib0ZC
g3utzpAjTsKVAPywMwJ6WjLUBBAIr90VnkuyBq9hzzjycd6D6AOBH7vZE9Fg
1g/GRCoUOvWCTLDrep2q/+K6ED4HrmReD3OYFJn01ZA1XiFqUJZSXFwX9Xlg
A+/vtiIWVjl1aShvmh27O6YVdzod6AHtsOIsB1szUZ6vD5iws6vHOh9XKbtZ
S+vSBfjKfT+5DN0Feph5rl3wq5Rfuo9FtjnWi1iTPHZYZ/rIo89WJrqu1TZd
286510wotGyJ8TnFTM9ZoKMr10NsS/eRYYX/lxjZhQKRUyUTG2mpW6YFZ1CZ
/FRMoZ/pqfEBHYHzOcNH97jbakiCqlpubgt4y+1iaQuQwPrRPhO2ZTo9mYjU
U+Zle6eVYDXRH+jjsaK1Jk33tOxxk3/71+aXj7UKmkoemmZF9u9SDE6GflGR
/lcf5NMN+T8o4ZFgm9IK9DllIojfeSfzQukLT2lTUSRoWNqrzm7Yn2sZ7CC7
SzdDbqC37h8Vad+cOq7Jl5xrDNxJ9EbeQwCiBAiSzH5tLIJZjMrx0+9b/JIZ
i3n+1EuCO6DT23YjpDbL3MX407VLdq5Qq+D1guXYJd09hGV4wmMJ2ZuA+Keq
A1QRnOT9HScW714WtqE6o2ai3KfUQfbM7NFRa8Mqcv5galiS9WuKy4pSgpOm
/THEPDRqzxKv2vuylQb5ty2D6V+u2rLkh9Pr7niFAelwmbcwKexMXd4tEOim
kpxTB+r9BFH9RJy/ag/hJ8KsKiMeRIjwlFO4DBkhap8jykkRtw8N1H/eQFvD
8pHH9pxFXfhQ90OG6TDTCEfozF2vXG+A1f4a+IZG7vAHU0XmGoysfQi5BTN4
2V3xJFqhlhUvCBlckqAa7vTI5nLTwKTBjaNcCfY25auYIuvHS88SmTEqT+25
7arLk1cXtYmoL8S1J8bSUz8X9rPExGI9xsPcgqDzWDW2uYnSOAJZKBIeKROA
7PPEYU0Pt3OIDf3/Qyb1dfUfH7uJPq9hHcWQ/MtPCjcREbPmOPSbq3uxkNAC
0cwWJjKAQ915VHmuDgku97UCIBAsmGa9O9QBDzbMfI4JyANfb5Wlx4I9J1T6
QocOEmvsdz2XNJRhACYTYloQ9znAe8W+ty1JjQyIr/ap3TI5c87UgF5tWcQn
1haaJ2ijNiGZ6cnMk6UoaVNMr6tSfo/tdskGw+7AmIeDsD4oK38nSCEKbYhm
BC9282cmBljxhrfpXX2Emm/qY7TjznW4VV9Uz2jmbkRFAu3nQKwXA60RsMmA
0LyXX+FTsXkRAdzYcE4jkQG4X9rfyKB8SHmi9fYZSNRK4Xbbhxk7LNbK2Hxd
8c6pvJatMS4Vx9YkhJGG2ZhAJg/beQnaN8CbsxlKugBmIKVAT3Ic/wCrcFPr
skAk8OMhW9pc8DJd/ljWYQPk5F5f9oK/MqFTbvH7E3ieCT8KlTOq2WY/qcJQ
XXYdCHyXBJY+v9Oc51Brean2Ilz26GNVaKGGgadKCNyx0Gd1yAAC3Os3DWSs
86GPzl4LNQoBNZGy3BABohRgPOGWqCnr8+ykUx/nYJZjexSyZhYX/8li5ZKC
kvh3kaGaT196gsxf80xkkP+FcctNLCSN4Icxhcdst2Co3L6FIgeqKqbWO30q
BS2+S+TNPY13hnn4M8HfOzpTcQV0+xRHSOyF7P9itvp/qmlKYUtl8TgQQwe9
f+/lzDBMVh7YrUJSnNtEZ3gK8qeC+dXfT5giv9P0q9tkRyohBPM64SRHHlDY
aezS4UBPr8ddVALR/SvLTwk1upMwq/Zn89v3/rGxdLFqtqvEh5e82rr3uRrq
/d2nFNdw8xNK4MkH1Xa4a7dDDRHoMqFpLXMda136fsdUS7ZbbZR67N+h43fv
Su/Oqz6WgJyLwy0VPqnHepUJ/4RaKIP+mEK+SjeALdLK23Ou2nJoqtWHL6+h
uO7ccDsk3EORw3apD9C1L0MshKEQYkzJqfo2b/1nA5nrYAxzwTnR6bJRJ/wB
Se7LOIhp5aXK0LsuTATcW/UW51R9F9G/TRy9zEClQ2CvlC5fNpXd3cFwUPtS
1BHt95/UWDDEV8iap2nPT5DJaZMzwLt/Ja7H1gZQgLv8egfXoIOUGnhQEyGj
kZJcgOR096WHK72PmiTdspcVz6l+B7r3ZF6zXH4VpoNTZKiSaVEo/XxMLa5j
QtBhJrpydUvhflfR0A5PETk4Jz5xEQ1mbQ3upiTeSfszLIBrM5O36rRM9eIA
MsQb296ak07CD5ELmCS4FEk/1kCFS7TxHKvj3lNELmX3re/TVBUbXXm1ObY1
JFDT5k3MXy/iQu3KcURNisKM8WwKICuQmzx20nyOl6jZ7CbgJ8PQ9UnW+RpM
euumkUWdvSgoqsZ4MzwWBA1GLoSO++13kAtOW3yeSkqsqqMH/Pohg2jUvSyW
/TJZZ0Saf/Aofq/vZ7o3LWxN9Z4OCq+tcaSVrFQw5jkpGBTy1EVPSVxHWBH0
U6agkagym7VXfjJ/aAZazeY90Q4gz+XErkJIiuvxwRhW6zAfefADOsOnJOWQ
i7TUd/f09TdgkrXfndh90YWj2t5PAIz1EPqCpDcJ2WSY8DR2xUU3c8aKfYje
uhuKUggZPN8WMOeD4mcAKvFvnvCMIpYU8k0NBAN3XLTMYOUXVv+6fcODTEAL
NpFA/PnTUtd8Sjmc2BgiO7LJ4Keih6RIHFJNbJBGdEuYEQPjhmMnPBUEYhiB
A6HG4VqLmtxRA0ZoYTGtKiLfpJGWSnCNhWoJG9j0j0u6iHZaf+AQWiZsymWx
fpmwQ0hmEERqf6vduQZmIOYb/fYYZfXqKQoET/YiuIDHUpZlzqS9joEsH8KL
uye2eGOA+Dqz8YxmMvU1sbs/qE2ZwlKUCHcpFXi+ToRpNZuZ4Cvtonu7E9Ma
fqP7fxEth7S/VtKWsQBny+S8+Lp197lzWLTUlF+PT7rn9A1GZftIjiCaYV0t
LGhCB3vDAEufw/fhMvcDzH2B6NwjBt8DzLT31oVi67t+bFWajNH6cE6RFFoV
tAx3eyEemyqyqmoJirxJxEcpR7SlpXfU/y5BbJ5pmuItxsWvzEeowH3Yo0ft
t5qhfiRsLmcrrtacrXgLwnvJyKGZMvrdDXXQfDdy924ywPBlyaJgWNDxRNpk
lupkTwmKkJ5ShHkE3K0eAiuf4TTdApGGeu5gm5/5gEek2qKEJBMHBXm0oq06
slO06GTvEZH1IWRBB2Xd7Ie378MsU2PoMs+ctDDvhyo9VrZi7kWaCaDRgQwb
+dyP0UmIUCMpZT7NxPWbGOCnYN0cSM5OKlNhc7htz0NlerKtsty1q3MdsdDs
nvXq4dfUt0MlmUVvXhUfHJA6Cu0NsgJjiGBaOuyJS/gVwq/fPvFrEQTovQrH
DHMq28JT3yEiVF9psc7Ej/SfOjqI2YuJTMHsi8wO6P+UaeT218ZCAH0m4kOj
q6GqQhQEW8lAH2XWVh2xZvD4xOBBamHL0pYoy08D7ecdYe7cilg5vR/2EbbY
MmZJhYM6LqpADiaRt6ScIaSBnLgxapO/sVyMDNRJ+LNOVumDHSBNOtzYKeoi
fpXXVex8YaxTn4geTDhpCFIYpZ9XnBwjJRFVkIUMeXHGrVK/agLrpg/mTqYF
4BQQItjY7MjJdQwzs2CoisFLerzXe1gQLmvz1ZFG2X4ApaMPS/8U/zgez9dg
fILWFzLiH6WTUUziNUDqCmUOUQ7StFm5fTdLDdk9otUNptxzLTor607IS5Mt
vlKV6U3hlSNo/KgAFaOhkIwsXT6eE6ela3YMJVFzJK+LZD6PJAwRKRm6tjkw
yA0hpIO7cp7nnDznau4BfgOOkcUUdo7/b/NtkvMfh3WCemTPqY01AYoonCH6
CPUyySxQhBIYjDJMRypLdYCskkueQjvZLKVYR6wSwZcvkyfWHRHF+Taa5mOr
tktcz045aXTMTtlZnoV/lYBHvMPaLGUxwkejPKdB+VShmdTdVliIqN+AvfDP
zCU6OYNMvBGjWkSpwFg4ulu6peO63htQqGgfLinxjC0fVnmTDnBghj+NCrny
jc5quUte4qZ1o80SAPgOYnBx8jNBD37nZC1v566KSvPWx1k8oJsO9er68mk5
0RXNz+LAHWBBHH5Y0pKf2cxRTkRj7rc4rEhN9FKRDaChyRjK7uta3LcKs5x/
oqgP4YXsOFL+O3xCCnDktco7tTqxIgA5PQ7Z+lYCf7ATykhz4ezAtm5Y4kvB
g+sDVMiN7tOG9R0fSUDNpSbIhAUPZ8vI7vJ4dZQYsQ1fa6fL/6J+gZ67UaP2
KlsBcI+2veaRMY1hAOmhnf3GuViGybIseZe1ml5T10ioQz+ATnmuUwlWCUPc
b/mCzooyidnOtys5wCNvG7gc+tth87bBUzBWqOytOomd1snr9EuWHjId9kx0
eALYXXJi2k0HK/ul1rjOD9UT/Vdq7bUZ+k84J5o86LilCPvQAsCP437/BuK5
YG1x7HLuEtS5mrJoLtxrIugwgMdLBfMprbGokRKEnqAIN3mXuaLjMNWL3Har
ZBElwGStiJBYzxpl3VV003gRwkNhpi3iNtihVJ774OzKfnp8T//lE4sTM46d
tnYltbjRI+reGIJlpXCojloB86gm1sybZz+aLpRYmKQkgkLSPbWQK7STSdEI
NqwnFOiWdQZXOJYMBqhshnwPkWJr8dhQA48JLeu0kcMSruZkOF43KxKbJbsk
uVUs/RTilwsTJQlsoLKp6wVRVzZuwgCDamqs3Go/JLcbNI15j2IEYj0t28e0
gIOpL0rmTEpwJdMBildyu4LcVgmpL01jeFdQ+9OSUODEyaq4qf+d/ceDlI+H
6A45kxCWSmq5JaCjk8Yf1tX1xi0PNaZotygvSmr4P3BgMavy6BpIsdaMmxYY
qBkpxJYRBChCYYlIs9Z2NXJih5w5yFtl2VFBbJbplmiTo1lBkSqiLtztA/gD
nKmkE3U1YyM5Cqify6JoZYXvv3WnWPkHEXhAYpQWbyAqCoCk7VZtVg45t6h5
xX/Q/MkaMGnbLzhAou7LTCO9FaHUtDsMkdwSwXncl5sq1bu7lZ1bESGsR/43
GaiZHo/9K2bDZLyJ1gLS5p8MyfEqz5zCmyHGaAJryc+R6wbrgdIfSyRqoVvD
DnUPaguAUXx8Q7+xA/aqnFlsTEfdiPyBjF00E9ZZWKPV9xlKS0ABUjEKQFlQ
cDLLjlnY/QpLsHcyaApvI/SIQZWLu4mO1DUCsZGLhZPJfNqFaEs2cUpBrfQS
O0DpRBLAbb6h6lPIhtwNSzPzn1lJ2yQ8u/tx0emMWtqyGW5MVFuFZZc5QjPx
HunbRUnWsqXfgjaVwJ7JScn8q+mxBHQ/2Gpv4zKvoreUN0s/bwQ2mfA8PlG4
uOGPfy80haSgXJQ5lNYw2LoNt0UtgR0AGQmxBud+Bv2Xq7McdMEOu71tetU/
bItpJaBeyn1I8sdLQ0tObpCopjjGtE8cs8uwUJtn9Nwh0HZd8yEpR6Bkb+wP
YKLTletYDzw0mNt4WmeYUtt4QYm/7RI8FmiGHcOdpw3alP9qigBdJtnN/wk9
lWMoCgrP20BH2b6b7JpK4SS/lJxzv0sbGAuz1wr7/11NVSi/IYpNrJ4SH/PY
2XBz6XITGGlqllq538Aa4ZPRJINvRaHzDPSDz/+Q4QKUvm5DI8OHk4GwHJoX
mFqztIDPBx6e2jdFrtPR86KMfA7yXkp3kAJRkaWi9TwD+PDXU28fpmfLWKOy
nrWdDhxlKs5D4sLsqK8RrLqxKCZH8px4d9gTrjU/OXf2RQkACKszSmbtt7+c
GwH6HFipnrWL/xUtSrH6cYEezFi7SSbhuh4CijbK1cz0RDCdcIsZefPI2pcL
bWxFnNV9n9oNwUv9ilCVTAjjTfcaMUzO+CQlC3ziarNQs+3d4yp9wmTZIGOI
4Uxi8MCYncAB4f/kMYOKqlZHNqIiiBurI2kAiYnmKOX4/8GCn/igF+uGepfS
WtNPCsJzV5NH9/U7owHgNnr7SUtQ8i63yXQShrEL1HoQxWxZ3Pcv8Dy3P42j
DOXzNo4awEiRIutAHdGWQ1wu2KkDwF6QcHXoryEkLC7DC9MUgl/KzDklsNuG
THoxcB6d6xih2oxo8sEaalcOakc5nyVL3uXb4WUtIpHLLA4IJVze68c8CUnI
Kxvdgh1gkcjguHg0N7wwfzSv6zHCpqCCx8HASn9Uab3tOxnSrRAsjdXiqLYx
Q2UzY7iQv+KUJEgkhBBp1WRuG9C6KVmfK++RDCRFaHs6rZS2XeXpc0EfFrr+
OzD1FTo/s2/p+Lpn/EasgxKIZfziY6Mq0Az1whofqTKRozgDq2DLFZzbeznN
xkVld01vR/vY0zaKK7ZLKl3mLYkIwZIL+CIyBKa4DndHCDP6n7aDqEF/8Kcs
PD7YeoJMbqR/h4CUnNMMuiNHKBiMSyD7kKNHUPO3qcYgBehNh6iiiI50iUmz
rdPV4zygHShVJ+CTOm1yJ7nJvwiPfM2Cq0GsAEpL6EVQYxeY3S/LYjJYDYHF
KGmiUqmV0N2bvEEHbdpnyCakqSTV5dcemQXVVovNu498isMMSrp45or24H6D
t4opQ2XxQUueZcPzgrefPNN1opfnEMx09EGGaejrGpStM49rlbZajV6GS9tl
120nq/6P7+Upfj2lisGsSWQlKFrhBtmLZrrG+G0OdwDqoLLXAsi/Zx+B2RXu
IjB5fyW37RG2tG29Jv20mKI/9YVLBGyRzw7bD+0PaNx/YHwj7tpgcUE8sTt+
pwdHDv/vi1ryOFlaxFgNmYDYsdAdKZNmVDgKtcmm6wyiEYlTyF2lqYPkrIYB
hvpVZmYR2c+i113VrvTEYnpqN9PeDiji4WOOS4vJr7v66zgKRmcwqe3UTz/1
921/TK0Li8/+eNTGbfxDmL7VECPF6/WXvha0olherHPLOjc45XufaetGaC5C
850vmCp+IWrc5YpU+EAywbdI27s69uzJGkbhrWZEQXCVNI1ehL2tUx+WNxpq
5oRG9EFvK19QfdtOWBxTtwGQFxhrwRFQ/25Xk4av/FTK/+Ipbq1aivItsBK1
jUxnpujNmwA6dQCfvej6Y7yQjoebz1gmyZxldDAcAqhT2AAxaq9ILWazmo7b
WF7sze44BwNtnaeb2auwcteBLWpq1oGDpBhvq9Ug34co0d0Xf/GWFBRHj1Ly
g7q4/vf8X/j824tGHBEwNcpJ5xDz0m3mAY0favaqrxelnJCjRWZbv0sZgguv
Cbwp8+ixjew/mm3FjeiJxA9YQnql9Jo2m1MwtkSgF6AEeUwNiiEjUFtwyczN
1AiM0R39t3ltADPvoE+TAV7neDdafJ4qGhZ4380g1ncrV13wuh3hPKOfK3rw
Jmf6Z1a2E3IlF+CfyG12H/W1HjqKAmIZnKEU8NRzORKSFhcQvksSmLMLMVGx
WrKhARGmzQv2/AQgRrVE+qHUV4qnHZZ/etsyLc3V+AC91pWr/P8z80sbp/0Z
xaqHImFe2cmkquoc69FRh85TLQPBWs3r/kjb9pObgibLRiVcu98xm52nD0dK
lIc5bJT3pwZRGm4vKvA/RBe+ZHCnjHG34kawsTtvRelLqEn+LD4y6QYEIpSh
hIMO+T1cQFCswDcYyTEBtut27NX0YAPt0figcTg0lGvoSINcjTciW38lDnfX
Hmd8B0Ic6n0y6E+Ik5acMmWCuYvwpH2W3GpTImv+GQU3sEkbfAQf/VdcCV+W
t5h0Y5SF9V99KtEQ1uPXXqJl37GUxmIM6BGL+Wn85eqj8MuFg/hinhv+IgL6
LZfRmBCWO+81zD9mtDT/3fEOI0uhZYz8KrgbhhWNeCsTuobiUNfceoUeYSyE
PTWvfUGk149huYe+2Tr7ofvJ2DBptWBlwfuRIt82waqfkrQVTVZioad42LiU
h7wt9Vdbm5jBFaY/PD1Y/fF25O4GY7kr8LS0h1VvJPVRO/ddxXNnF8oiO+ny
EQCG+FGXbZIpVjCKDqH0iWBWPh5DqxZLQ29LZLL2MtK5GD8kyBVQdpZ+d1Dz
KO0JIApm0BSTPIUfp1RHJ4cgeWv83UgllB/cmDQlbhTcvrH+m22O6I8cj8aE
RVp38uQBV5opdLdfGJBE2hXd7VKkQnIBoygCYCd2ZfaSFJltWVSvk+fNwuBl
fy1Yptnkem/AGEe1lSKk0dQ5kf/bpWeLkoB5nrfu9d+ZWdDxYK+SiVTUaqoK
7XD1cVFcMTawe8e+ISo9MH/jFx82nSL3xlDLAkukf77uW35dPb++Z61WDDDy
DfTh1Xq+sNhtQouX4SVkQRSFYcs0VEs0ssNjSSssiUN/7PbWXUHNzTnS+Tzg
22JkJq+dOJulv0d1dMrp8wt/8Ax18sfIegixVFjR98OEmSh4EQjJrpBSMS/6
k/wJiPvyJ46ZJyVF4hHX9lDFAxEJGB+twbFdi2oL9J3YqWDuV3P/5PDBuYqT
pdui5fI2liiEJwwsDo8MBGjGHzgZZ/wW9LMJdhDdQLnK6aobLyhYXjZ19fto
U71s43qCWxUH7uQ23XkPiGR7eLWEG5rjWqqVUOOip1yMNdU/JGqvgJdwWJZJ
bury98WtTejRKqM2DHS9lTmb/XpNSPuaQJxEVf0ykhQ9HCROL+y2HQ0/Z6Go
rHyhO7552RK4WU/xeVg9tKCajfnZK/1lFBX7plGc4zZTssITue6Iir4pc7hk
wuFlbDbASGOl9eRRC70OtIiS75DDDCTDD2K9QYDjilhS+f5D2wTvUFvj1FO6
Jwihn12sKuTSqIAwvE7MGnKNgYiCMp4qjY41RlYG45tyP+2aRVC2tQcFqh1B
HojAUeh2TzB6BaJjRtg7k/VWHxjIFeP2KMYckr4TuiCsbNlfrP4tdZRdGp2Y
oQtsxd2NJEBs7xWnaxsBi6mswAmBHuJCGf0rNmxJ845OevYadQxWNDSDi+9h
BdVKmsq/vWNuYAkDdhMeGSpZhXP7HYy629nO896B8r8Uj3icdDZAklMhFoGw
8pAo+/a6Ow0HHQQJJeMB9Bz+GGXcI/5JR1VNxmNlu729B8L9NLheOEGphEdo
aeW4y0PP6KdhxR13kxyfqhXcyDmVIsT4d3n24P4d3E53d4sDQ39KNfxJ01fj
IqVQgwvpYQKPbrTmMZ03Tv8K3DSGFpv0gECRUKr+0SmHzRCQWJ2dscxkpPHj
C6jIsFqatLnSxHHsYzHeZlsvnGykOtUr+QPEyKEokIGo+T6qcVRxKxm5Iozx
yJPuV1jz1zpjZ087ZWgY9MtEwrnszZr7PfTysai1JsDp3vIeENPrPj/slmFt
aK2joFR4TXDeCy4GF9AkvFG/gG4HtQjrPSCzFIFt2F8uwqQ7RJXyLNg0pdXl
USmab9mERqu0Rwdw9nyi/7H47ToKafMrm/NrXFblIX0W1dBdy92TksSbgJwS
OcJhgYOTqaOswl1xxVXU0J+S8m1XW4W+zTqCFX7b6EKKx7c2rfOPoew5WlWo
ERSfzugsPSFkNx79DPyP97S4nDl2qcb7PKybfGZwFeN6vecT6rk/IJSfru0f
WH5el6SxnzI4G9ldCvpTyDbCddNl4Wz+toeP4hWjziDnNiUNaz8OCj9h6ybK
1lXNdj/p1G2XPJVxWooHFgKxgJfWFHf4lk6qZfoFxtgovsAz06xa/whwhBq/
5RgbndFQKGEEX9LoUXFB1m8qYgKd6rSSQSC7thZaYfnhIypY1ds8fS8jXBk+
3ZDI9IqHYW6SM2kOLQxnq1aUla/tDwgivro+Mbatb1pg1MVuQezIkF7vuHD8
qFiq3P8zi+FWjctDXyppCS2yOoPXJXWA1czZ+dte8nn64c4/14Tldy2Ae1Cw
+ytBwy/+IK5bRJOL5xmcNW2EOKAtrkAtgrl4Upons0xmyRgu8f9tI+7L3xbb
F7W9Lg5l4xnSlFtV/z/qUrYGav0HvCuC9GwPSY43wk+UdyFjPic6+w8KXDCw
q+5jofAqTHZNa/DdzxLPjd6pW91z3nLbpDuWgNJatvWWW5Njg+bw0tW9esBY
Wn9nKgRzJXb48/NC0D9UjiwCAchMDwNXyRYW88fTGneErPw8liArNW1B4esX
gWuJhyLXKBTipdr1oigFESxcCZXER2YOvTkG439zfAALXi9EdXDTbKsGfi2p
zfEk3cZ4fAx1O5bakQq3XA8wvNTn/JBooahGqeMWhZqv4tatVi2iNi+Q3hcT
0Xl7wwiPUsRygJtD78mU0siCUvc2DP2QisGjXQGJ61w0Hd8+O41ro1hRrxw/
/UaRzksOBHiwS2rIZBzQLys6qYnl78I7sCYi05AtiVg606sdzj7YufrT5lBL
e48QkEcvh3z8yeUm/gXIQy5625XblPLJmzXHay8dPofC1NPVyDFmcAH05iuS
yW0fafm4JF+EVAhRo0GKP8zkGjcbBnEHRu7/rPn2fukKvDUvRriF4AYnN/F9
e/UC05rXBWpB30kQ9uATxbRiqRu7E7et0XvwtupwIi887z51eb/qmQsZ9NCU
OD4Xkn+bJ1w0QbbDZan58CwGXEytsqRvpFg9r5GF+vXevZ/m06InQ+swBumY
M1XraWK0rq57/K/EijXzXBzBJR4FxabiuFeNmxBCufPwJ5/8K5ZA8GdW0JLT
6jHuhVDEBntbbsnR5qbnT9enTCkPcHd4P6g9L8891xmkB95c1SfctUislf5L
vytM5dDYeGEbZRiq1Z2VzK1YuAEVSoLkmij3MZV5/rpqdMB1IyBcwCzj+cqd
pm5z72cpdYqOhOPohIq3Fo0++bz2LeAw6VJMnkglG+6DQNetsRFIKknlibsW
XzdfTfHlsmRyFGVgz8sQxldunkPkLh7mtf+B+HxBp7ZaY3WE7VweBA9JrI++
yt2vqjbP7v9jKzWM4KRvA2YEXMkFYUnd4SlXnQQJmz0WjzSaf0lG6Exc6nfh
SJJCjtKfUXbtKl9INhUtqEPHfdQRhkpMpO4gM5zSKKxcXqeIa2QR5CPFfPNl
jGQGCLLYzIzrmqZoCR0G9sX/Mpi70+gfZjCgBkvuBcwkrwnK53CQc18gwx2q
5ggE6sfqPMn2Ng/jxJ8nycPRGV+JB6bV/TnO4oEqW7xBdtqAtnCBF6nsuaYj
TvDxJ8nr9qlP6fvkoNiFVsG8lnjAhx99rbLoXi1yqoHY7ofXVlFcveOGoQEL
D37KNVcOpU4CZcsUMChAga4aEUzpWcxZMv5xIeEtjHrUY39aKvZn3aGOR2Xy
MdlqBUQ5GU3Kn+3M+IxkOoMrNVQTTH2HcawF7Twy2sd3yY+GRQiyhBK+Mg9q
deGr3616QV4+9/PZdVwCQYAuA+1wEmtsRgWRYznftvYmrHUfH4yPbqI++oJE
QVeJCvNxpC3W722bY7SAnWPLVCYVfXYFb7IfIrD1yLujeh987vbup9UeyMGC
p9tD+MiippUSLYkMI1NbOeWfobjlc4vtq1t/NlDLduirqXAslAHAKkNBfsU5
kcUVfajoNRbcOPUGrUZeEvNjH8dNaABrguKSLR0iFnHNdK2MmUv56gvy/zH5
fBHAfQLJPZ4LWdHqT/LX27B/nMUAnuJBDDblxh3oet6qldW0TIABf+Lr7EW0
r0T+alyIy50XVza0TicFjRcjfrP+ujjFir9FZ+L4o9HmwSeW5JdHLZUDjw2D
pXCnS9nUtCpI8V9pcOClJHgbq8o0ISuCrTMA4KR33pGJFJzLkcOBtTzQ0169
kBWuHB51qq4/U39v+VJIjbRzxamYtX/sbmfTVG7jEDhc5iRlEKks0QRYHQ9A
sQtNlcWMbi10j7f7/7MsDpqe7dulMfPMr+VuYV9bM2I7ahjx/EsEBZs8HWcK
I9iz+pIL4R6NrT3Jlj+M+4mDDbWWxG0r05IPAZClCZTMe0gqwwNjH3j8flo+
DTQ00PaP5/JWghPYkmKTx/a9sC0coC0+z+P47Okcv0VjBU6KCvwuIPVK3fWK
qKRBzjPiH6gSiIQ3Cld+DVLNfnREMXhDDzqGU1bQEDuQBC7yxfVUC+ovCVL5
Ia23M+YtkfGPwnB93+xNWDp7euTfr3BjT8N+pqF4zayaxkoH3+f0go+octuV
mhmSGtcrdZeifAd/DK50GSYTGuibUcqvGRixOMNZE5uxSnnQCrbjZ1ZTDuvC
DZfmKobVVWs5jHGfYXAdrgHc+ZCbzGPMikxOtPk7ReTDifflfPKIedU3C93M
I0OX/O7tYInGLZbaMe/2CbfISBTfVXFyvk6xpDeb4URQHTWv2QAeUS29UK0A
WDJijcK23UIXtNN7WbCnnBhORgPihoMuHuX6dNMgzMlpqzZxYnwe+lmKSjPv
RCP3EwXrIlwZPloT3LUrD7GWj7aljtR2Pjuh1KDt5S9I7MQFAhqwVkCi3+F2
IhPpy26b1DBJ1Yrn3yiOdVTMCSNO8rBiGl/iM32BugWfKSH961vFpptpb4iZ
CP0a5jtQjNoJUfC8YnzH+dzKjxo+PQD/Hi4jiVeLNDgsXyFZRAaVxR1rUWNs
Cjxc5yyUJ2zgiRji0hTZMTgAqz7/jHaLp9NOlkwIt/EplJ8l0hrbcD27keWx
tygaP3Qxm3jytMRI5EJBRxIbJHY/unapLRjoeK0ByzJJHJlcRGcfrtjWjY4M
MKxcMz9EijFlWc/p1LzmQaXp43XNuNaQLRurDjgfTkZUi+IY+wTVcjnTBawP
aygjIyYFANsLvW2PQYs8AcaxbGkoSO5QE+UI9oRZ5eZ0DnX1+FgtwDhD+LpS
L2FES3Yv8zAlI0/Yzy5lAYiGC6T4xKsh1CrDJYZ4kbepqaR4Zo0zy9Z4lGLf
QO+15O8LsRKDmO5G07/hml7Bttsfp2V1YRweVq00ZiG+bqph8LA2XexI+InU
yq1Pb7DFyLQ8XH2QnPvEP1RCVpd83F53/AV3xCGjiFIXrWifOPEVdLAae/jR
SszJgtSd3/SYb43Y7Q8tWJghle3ynUedtYWBskGask3sDOEEAajdXFV4OO5w
MVrgV2hMLU0yfq7kpE9EjltmlO50lL3GJWYiCTVslFVgg9nQrAQkNTszBrbV
vXfEgQhLYzyytTLHmyMhHNAsE2A15Bp7EnfqY1+MdTk8ciFVvhIT6dlBmIJ4
1VZ/vtEfbYdfhofV5EStSESFTUWrZAgxZUTH842jpQj7IhZioSRequBh+YJV
KeIhscJPYSq9Wcg2HV63StAIPwXlUJKBwdm0IcTh9Z4KkdlFTq8Esz7wv2ou
ndt8tC6nQi24qBUo968scFjDJFOW00z/cngtNnaIAhshJaf5KMCo107Zj+3Q
Ij6/2ytr7FccWCCdjPZE6eWKWJv+7ykolP7HtnHPi3sctlrJPQhpqJ/n3Yf8
fpwWSzpauQZrfZjTtx4pg7kPghLJRLaWqy4nPD5ccSxcxxQSVG7bTh2OYbq8
rM8xFHTfOi77morcXPRgzQWYyhDrM1pa4qmD+bUYeTavikdjV2dB8lltsmne
Z2Yh/AzgxhRDoJznvY5BTqdskXlaTEyoqVY0pPqnXnJGZQ1Xnhqbxhf7A/IJ
NxRlhaFkQqWMXv+7h2g1fS6yTCEihjoqysBGOvALtzbf6+I6DNHLl21OgChz
r6bW0MnE84qdq/CU8wJ19/oGqnI6Obk9YLY9QBpZMfrgE0K9b1NA8XH62nI0
nonTN9yOhq6t+1yFXuRJA+/LUKP3LbGVRMSqhflCSMuhc7MKTRIvvWhdCIfk
dXQ90hCMBE1wQa0e+nsfdRnJXx8EbZ10RTxzlVGwOC+T93k6YV8PeB2V22fj
jjsdRB6gHOLuYoybQffftiiVtIpUmBB6ucRkvklYKeAsFUWpb5A8vQrBH3nv
hHxXO+mEtKMQ8hlFrOtG4pVv47Re1Y1+yJpsNFgZEHFG2yIVb+bTWAdlBGqL
78VuuJIrUN5FBL+fVkDwEi/DY5BgDU1eXavJJba6NIGpCb1zLAwMCiRJNWQD
PYGGhFW2BQiMgVo4gK3d0siYrzRfmJ7mFnuS6DGmXP1tU1bZmE7n1XkiLo47
sIM8HkoAJ/CkheXPCypBFee7zUoOTbyxiZJrfYRAvB2jLnbBOokUp+/XUqlY
HGyp2/SFAT7svC6/MJBp1nyGsDUn7pDdf6EajFHGBnd/eEtLUzTb7Wb9+3Sp
zBKoInIr5UR9l1VpVHSf7mei9yP65mAPaGl0ZCtDBMK7AqPx4Of0gjkhER80
Egxbgf+khgmX0Y1e3yLX4fRbIHIX6hRtCg64MjRRjcLIjLas6kNzdK1JmqWJ
pMX0ClNjxkBC7EyCwJL7sGV4DqSzgbg4fPTADMniohUxI+XMENqRq+yCaR/C
ijMIZx9mWvxYWPwlF5RtC5Dp85+hmJIOA3hk0RnCy71Z0ufn4gGeQ2wSfB9J
RZRXdloXbZ7u0l7iR+SzQQqG269GK/HUZxIMDtbBSlLTdbtvhDveq111JVnk
vn5HjLJpyh/0SGcSxfaRYQa634YxVyrVi7t6/L69f3Ac9ZCrtzc4lkNMHmQF
6w1VB3EH3jDF/ywOt8b68TgBaLj4vCiJrCzJshC8kT3PFOsCZ8w719GtnypL
/Ufy2MrJxQT6F20Sr1LqRN3hc71yMvkMXJw4P5ykJdC7qp+IOEmdH/4axYbO
IInUXQifoOkFd4rrvRfckdlfJEepL5QKbL1Ia/cSEfUEvsWribgd/u7H3YCh
mCUTdGRKk2rALyhm4DeMWi4GP9eyC5rs0kh9CHNLXDvI95qKLmErvoVHnyrL
ajtNMpcUxfyvN2QZiiO2QRm7GEJy9NJI9DE4Tb8NuKPyUj7MDvY6eIyUzOFb
7i4HWVjPiFePLnOQti6x+QFhYO1JtpYoARmyKGPPWPYEQrYuq0Hb2mYcOTAC
1UL7PqNpnDCAoWlhWs99a1RcJ82QDsVWPvTc5frp2It0pShLrZiJJfk39TTC
dBa41GKpEkpaWBQPkgwctqXkNadwYkD7nc2P2wwj8jsopy3Oei6H8z+mM3oi
HHCx+MULpK88ZNxVril3G9hKsrPPft1yvJD2JsdrY1O9BlqWdT+9QQskT/3G
AQGO+RQlBRU5GZNhPSU+znO8B1bXyTJ+gRY9HbVwo9MEbyZ2GFw5Vxume9y5
0M870zkBmWjxAfSMIqbM+agUvKcaHPgWCRwd/UOr0skGGfaMiJs+izD0Nu8e
NAE0KAp4oWpv/R1LjXPJKkbZq4G1IvhZM+2AHfHKfAQXApiZ9RB/THqolgtj
yws2bFVOaQ1MZv5fwCMNJEABwZM7MltKh42KEr6zmEOSnBlDM+aFU5WO4s3R
F+ZnchN7qajYtUmhDFlbdRjSoQQPQekWxmcOVmICSqFH0ozMZbzyUJ9lFLU/
3Iae4VlwIsrw4rc5S5m21Jdg1d6nzB72BsMVMFpyyg9yWkjyWMEpoEWyTX9y
WxVuS15YAeAEL1RbteyIOqxoPi1DKwkdCrAsnJWn6HI8t38V97g6/QPnXz4R
/nQ1Gsr7UANXuKA5dr2xNvGg+PHw7NAGCpY+CMuNvo+9zz0sGW2Tupt0kCid
JcJ9HdloVOjnr4WR1GS2GYQ/Iuo6Jf9iYe3hnb8/Ly/5unFieXpJ4yLXmUIr
SvR7+jeJtbVH6dfAcgz2FuVvygD1xFeH6A6K9H/YMTUhkVZZKMAqPakfTaAv
jBxQ3VEnhLAKY/7rEXNqAyEvSiy+uX/Ob9iVG05ev2KC5rT5ZGC3WLxLnl3S
PWJulH8Poj8halbKxZ4Q8gxzScwj3sENTQCPCKS2sZiosBXAVfgHGvSLTK+V
LJsG+pOqshVESdkPrOhRnRjqfaL+8CYqXhuq0xIMxYGFo45SHkZ0u5M0mxai
lnzxWFb2cuqskl4USNol6lyuEtXUvD0KPeklaSDDkumZpSb91la/mvXy4HLe
Hf6fi6Oy48YXXejIGkvSuSJuumYEFrwzPn4lHeQsznbwJa6+LeFCp9T68rQb
/RNU86hXetGVj8w22PgFjuQhV7vWeZ6OKcETnsO5TEWiZVXcPeidpi0gk7+0
V8xui1ipXPjnyGZQJW2Wwh07gWZ9NEXGu5Yi9ESQ4VG7i4Mw+6MoygSe2F2T
PrZ2gYpp8muXOIX8EqpcmdVv9XOgPHm66COhBj9+vblEdGkL8kIkN12b0Rwk
RThLr9MBwzVuTf/xdbCxvxh8JI6W/9uwZCpdwgQ/CfIdjhgJZ4N7nrkOatnR
PYN5t0MNWM+t6FNjRB0gg4Y27zuHXD5aFEcg4a3o7RqtIUCG50RRjH/t0gRe
zRnyq77PhkWOMhXa8nuLgPcF+vWj7RCVSy27G8/FYef/7wPejbpXoevDw4t2
JjRskHxZF0ospj9cwMGWj+lbkXhuDxSuNO8eJbd9HJrYPsekfnDEhmy3EV0p
Nyp82WecGyIMaVPWYNvwxyYcnS5WVAwbUteLdTLxff03BFD+GUoJctLzXpc2
gE2F6K+f5MIRZitPfU81HOiPlJ1/0id13J1jI5ZKii2oyZEAYe+IgNlFHgOo
eZSKq0BItzY/g8uh6VjSJXfYqH3P4Gp03x0F0yOI0uRH7Ll3N8YHl6oEQai3
WEI0gjWRQJB5o1fNirFd6t5avA8VOAVLeobSjyb3w1ZXahy6gp4wQI7gFGpt
Ffd+lF0ItTOKLXg+TYgwyLAc6FHIZTJQpUrqewxhFa03y8g6jO6gjFjOa5y8
ySG6Lh/4v+ChhkXQ6x6apubjGQ71/hZj6O/UbG2+em6Q4OHXFALV0bDO3+lz
Tbvnj2wmWZ6CruE+1qxsmvYXNm2Up/svj1AHfnJJG1D9WOej1jrBr46axhBJ
nJOeBFKMg6/JBiVHeHzGYGaMJzDGEsPAwcIEFI/IsPBu1p1WlLCNhEW+gL/L
VC//1SbPy+zOksoU0rsbLx0gJP+6z/ObnxS4VnCZAyK82B/dZ4BTi0lrKEi5
/RXyxcOYcScz7h0a59915lyrQvGn3mYH4QQ+o5YC/niAq1KdZHTyIocm3/Zm
VkiggiSyzutSPWM7UtltwSvWLMuEgq6fewxM1ryE7eNCAsvFOzic34vjq588
UjvoYnLY11A9roKKvgfj8FqMm06S4FAfziAD7RI//v/go1ipE7KyA3YxNwzI
xOA4tF7YGHo4Uh36Js/88pvQXe7KR5GCEFhmCYoyKxtCtdGJZbHE5752Qa1/
QS1VuOksAJwSoZHBb1DD2olI4GJviix4bNBHDhyrp8L8H3026DgzVdjcbqj0
Klr0z6OSY7vVMMD9NrSuBnEgC1vbxEKWTdl8vgkNpJfJw88fiMelqmndk0/w
/VlaU9gC1hXetBHYvZmOkBRd2g2O0NsyfTIMqDiAHETnFDebL+uPl6CPMkJ+
1OLEqxxCpBSV9D9z9l1cXGYCdim3NmYFN+nGVSYOubsyuK+ISYQ/jiNhotDw
/J7kyRvBkJ4gGvIZ1pIBiQJmBFrV7NY2yGgAR4VCnK6Jufl7OtAPNhETCnS5
6O2GzwZPggm8WytL4ntjIsHj0uvQsY/T3vzcrusCOQX6zWOsGoz+3h2Drd98
nZLFk5i1GjrT4om5X+jJC+ny9JTM7Pc9LgOA7nyKakjr7UJjkCJx7JAcXXZb
L5oGqN3oeBSdr9VeposBEiAPngJaozO1XK0cRgjsOGP9rWb8+a4jR1zzlL4k
r6sU/7QfQQLGwHGnU0hUfQTD6618uwiu/pqhp941Mx8JPcEl4vTVQxrB3mdf
BM+SAKZZVvTdRNb5YGPwQqFu+aesalMpnuqhvzVLSP0n5mTF0z1XBI7C9d61
6FRZv8fu/D7BIUkUyQRjGISsGE2ytnuBIBoLAsNbnWEBXcMYTPPuCB2LKun8
o9M5fjYlp310lDMNwikebjuTjECR3cEwQ8JWZTTI3z+8v0RHV8H6CGKk2uZn
FqJyjKSeoxg3ammb9rQGKy0XIBECBO27nKRthZif/oROVxf2LSIb0OB15kD/
trLgA+NUp3AvN5gq0Aa1h6fVLHH2JCaOUlcjj1W2yg7MUuFmYv9FM5NyyyOz
68PKxs04yO/ZbIUP9frvYpOtC2On33kjpMhqC/yfZkeBdSWW+G+HC7Ziz7oR
GHPWcM5eHNl7lEjMvj0lPq4O66eJHKpIN0dLOnWsy6eF5mgD8wRdXDx1SrvG
zvEzkIFqAv5+PdQDk9U4n0GsGrjgCMp1DHuESZHr052BgIvHDYcBxlkX6ot2
+mETtR+SlcY+f364XbmM0DW5PvLZ7WbkjNGhjP/Rf0AM/yAuVv5W5LzdzyCn
vch1Iy0FJWbBk/DwHAsDF8l7c4e/stRM+DGAXy6gzuW7y+CY7viPpCYyydPa
P87b20hgOX3hMzc2usG4sh0kY9/EKVU51rFx1A1Hb7GrkHfwiDuWA/KqYVuP
DPH88Jn/Z28WhV7BGIUnV+iDuFq3y/zasVYmndGwmME1DkobfKb5cwuoj4Kz
eUlJ/tjDtFpQqThOV7ZUZHx1z/vkIGih+H1TJhvLTC7xEtl++gauggzExgjQ
2sCjPGoYDMzaq1W5CsleY2JcOi7pXNpjkLlngnBChKel1EsRJjWEcltuNEm2
gW6EFcY2UsY2o+HDVvLPYMHuQR4RTc982lAgsPRaP2Nkjf+fuQn2a20cuYwk
j85wiHDYR6jFVBpucMHpXAZEPrzaK4B96i2Bem52yW7Z86mGsDaooeMCdhtB
ryblKY1HF2w9DLKjQwjR+rcyQr9ODF4g1Yn4Xt+ZD/zSOklHWrJmT9aHMUIa
Nlth4LPn2fFJVKLzk6DeJNYkMjL5cw4zaFNgNpbX7gXNSjQxvhemWDsjCx4q
/2P5jbRGd/ibdLXpvB8RYdHk7utPUcE6kIvXbHd+5T5WPP4nsdPF6upKHuc2
xWE4EtQN7+7q40Mcjgkp6JnkuQhy7t4Tiptu0QI4CfIZ0sm4nreXRrSIfolR
WlZGauatbIghp14bD/gZFKd2wc3topa/qTgdsG0FaobnsAQEeZw/aSfyMn5W
9nw5HClV8ETfxLtG6LMS1io118ExUQx/FM/mun5nv8A1ZF47IV3Vq3Ah3XsC
uSK7cYLrMgffAFC05daCWin8g/B1nFWGmiKbHaG+xolYCwK8OHWLXAmJFRzT
JBltipNMVamqHWMQOrYmsgABIF8Ofl0Zevn/lTAqiY/zxFazzyHyGlO/kKv+
FxxlGidyqwk4t1D3T4A79ENN2Y/QszkZyXRdeO4g3lZYZMVqPQqpCK7NeqlT
BGED3PeXdau9x6xfkBD0Js9QDMHMtkPjk+EZD4lk1NG4l7pvTq/r8MvaAOxS
2cbcHVdR9OoafSOzLorLRd0ETrEoz9IvoFAMpDLqEfKkATHEyEpWX2vM/wWn
xEZcMMXY0SRUiAzXnlm32XgXI+iJHJ2TO8NpMe9AtDRG6/f7cndnq1ARY76t
zje/6uVANYRIBdQpn0kKQd9ZZRo2M0r7XuN6y3pzp1zl40ImxbSQH92GPO6l
7DN2GHH/zI7B6NrM1+pRPGwJ2fs0IAk8mxHyubbUdzUaUZ6gTMGU0f7Hr5cI
Rz/aDEZYCn5+iw45ea/IIxINQrBY9Xh1CPlgU9cHHEJcgCFTXLUrd7aPZmMo
rT9xZK/5iSmXEMlgXEC4INTdYPod5WT0FgbUsVxH1ajtsizRf7KQNTJiIiz5
b1Dqwu/lMrTV7oOF/MDu6OIU4zce1XfNTamafBg/CxECB8T4C6VcWU1hUCaX
LPw430GTrnvV9WSfhSP02qk4h1Z1uhJzPz1q6Tk1lG8HmdP7CIa0Ox1IQ+Rf
aveSSOrwHP1WdTU7iOtpc0jZhLEu59ytQbxLSrWbEhPuptsyhRbeoYvPrkK4
YD+oK445xH9sBtWd+OGrKzkDH20ru4atpLxnszpXcBMn+bagPbWEVpMtwNDm
JXE25MpdsqBnauY4x4JfwJ+vIECL3d9KdQrpZzQZ0dYWDiHsAb6FNOzKhcVz
Sc4erof+ZGjfeuhOYIIHUJbWFmoI+S/2S88wgQaHzlUBm0gHGiOtaSshXht8
rtV4JXEMp7+83nvhjglDjt52erz9DXIfWaTyxX04B+cNfp5nGa3z6fX/K6Yl
fg3RLyidJcwqbPR6LbIqJQuq4K8xy150WeDsPSMnN45LAhL/3WsfX112L4pN
xzW8gakqcfsZ48spSjbfvSerQAQHioIvN2w9lJrdf1xnZOhlROB+zqJhgOg4
TzQFiVkhyc5mSGoyC1aoYf7bfofCgvlhfgK9pA0DiAIvH/O2AIpkIsRvzYYV
SaXoGdhob0M1f0QMxl5+tzW/jO2Eq5en1UuYGcVip1gRHt/JrIoT4eKFSAvy
n6eRlkgD8GK0YcO1/Ql4rLiywrZfzESWHfI7b5l2KMJlvEttUwfsklVHxta8
V7ThBcAXkLXBniUqroGCxD6VhkJGyLLUG9Gb3tkFSv7ZBbMjlcP2mVYO4y0q
SyXg7ahaT07U6Ief5FZtWs+cCWz7aHj4osF6MKxzuQR64yX1Xg9NUa56pawC
x46Ma0VjjOo/QzV7Mg/UhZfjnDi8UUv6d5ZXmv1/pL9XvCyk2ESMTYhPw99n
cmmlViO0jqnDl93JQ3vve/EwweEIldncPDQ4XVvQltFxIkBm3BNsWk4ghW2V
nPz0PqPF19Z1QgXoW5LqIWCoi0nQ1qfaBuSGx5+r55MpbzLKRFKbL+mGLGHh
KDXvS6ujzlmYBpQkU9DGkeCsmgxv6IcAIL9nX2Tm/MBeDXiTObS4CLkk6Jk5
1Vog5RSFNIfSio6v7UNGJUUd/0y3FrHYrElMOOp8Z105jImh0XLI2ITvRR0t
nxW8C+tsnZeMbGSgo944tTC3BhwEq1ya5N+b5Fw2wudly+pJOxr2FSvQOo3w
rX1rjRL41C5YPy5PJuvRAuZDd9cA40P2q8OorMisK24SgpKQul0qDDwKX7F6
1Aq5WT/Jx6OkJJgtdW7pJzZ4zdqyHsuYgYhFyPuqEdZU68sSaIQGfF2tqNwq
1smH2iDUjV4tRwO758wNXXvIPoC5kfTT1jFGp0FuGed4sFaHJgsCHQ+ChCPb
K615J6SEhzCeHkwLH80xu4pWs61Rcg4ixjfrCruUarYPKn7pR20Ciqi/I4An
0d8jbkzK7V/2d5jc2/h1w2zh8mnlm6EWEkHtNudh3rfy+89kljCww9tLlpb0
PZ+FAFEQ6ZFkVbcHkpUj8PpSCUbKvyhSn9gavHkUvbd3wk0/6s0QuLyjuBN0
ScWd+gI9tjWhKV0bJH0GE4p12rlS5HjipIgreehnWCwiAUr3fRZqsWPfSnN0
8BEtu5nJb6Vt1vLyqia69RlUus5BRcSVOKOjw4E+PIRCwkfirTae02pQaEov
qmMRsU5NmVG0rgrJWDmVrCxOxM/hQ6FS9VCT0mmxhZ6uKB3zV5Nd+7GFImcR
+czvOJLfpcS4+zt++eu9QACNSBgkOXf7QUzLPnKu7KbueB7i93NmLbGpFO6v
nRa9O0hZN7r7ZkFVhz/+vtFllxxASUf90UV+gieV8BNFl5s8MGf6MfPBSPWU
xIDwN7Z49tCBVy35igGfuXL9MRjNTfCVrKz3yTb1yUHHZCWejmjW6lWewFVo
7CvhKPyF10RiL40doeKTw8JBGi82LJe4ZxAgoA4NFag+8uEklNkCRP94eKHq
3/8ia9YcEEn/mGb5ge7nQoKZYn8c+3GsF4R8A8dvLwky5tEiCbG/XlbSyWB/
j6L0SONYvBrKg9XPcIXdssEM33FsgTeohdKYqBNfAf77+5VXXSJ026bZ6mkh
83zzooI2thT5fSc1ZZTNLyKul3rPMJWXlProWfySgJDsX+LKkkKCbkjeR4F3
UiK0D8v/FV6X7oqnHqabeaUmZJP0IU3JaKoC5ZFVPmvynr4OGhEFfRBOTTSV
GMSVXMxog5TYpqBHQxu7V8HRQ77AidQrWWPrNyysXEQzGXY5+lvQtKbP1RDl
7bfqnmz5u50jJRqawt85DC89xDnSmXBUVLQCUArt6PD/ey1nbjTX9rTfcUKf
66r73z5hQX27TGBS43hPk/Yq6Z0YUgwTsmNqc1p0jI5bBDJYIS4F1IbxD1V5
7TIZ5c0JFYpzXNm7RA8gqiFdDkuBZC6Lh3Jz2vGdQzwEQf1XqZ2zxkF7ndpy
awnAjSwnEl6vHOYgfTvUA5sbbnFeSpWq71oczW/dcU7/jmdUtFpuXqyHlOZn
NDKMRX+Ewaxp+IWDmTeU8Ea7ZxEYLiStybU1NzXiYTIU9k7H8CD9TjxoZHQH
V9M+xdch9NlIsBMJi5Tj84jFDuXpx/LUi6XnWQa6jn0FvVtzc1i/55UILm9P
P0JS5u38hCMKC302o+/UgnOKiw4aB3BPZAFXv39Hw+F33UO/lRozIT0ZFPK0
rvZQ1pvzB5diuL/lIIcQ+PZGhy2tiX943r5bLod8MFo+RuVjHjyD5UC5eSQR
Z9zG2zUmidXvf3fPaQSy/GLIkq9WKWPWlzvZEnTCmbDQI7c+u8IP/ZAbxGEy
iSAiScc3VEPUaMwjDHgTvuKP0Zxp7JDXrLvy2021dn3jHB5Tek5uJB8k0VT3
9dRbzufaVmJiCr0picsaYDKB9wqeeaBVStgEpA4qXAAUTjGJGU+8Fy2/ipR4
alD+Kf4ZAzwsmzMaQH29ljE1Dr3WX9etc/5AhOV3oNu4RxPq4Z6E/LQWInrH
4vhTNiTT5RoXk5QZry3qAul3yP/CLzDLMH0utWmBlNbZGQIUFyYo4Pl83GJ1
rqGJ+vNSGz60FGr+uzJpB+aJ/wF8zZkev9qhM8SyAJYDr1GJSB4h6PwlHXXX
y9UMLZxPuUHjj3RKT+D+8aGZoMw0PJT3A5zmjIZsr32rAtxo8zv42meY9bZV
v9HKIN8yKwyR3QBsYBVAmIWjCX7BOXtb54232AOntiU1XhB0hJRf/2p6ijMf
IYPCfJvn1MJUPd1dSxhg0fvfVzSQzzSmE6kmw/EA4WLj5d27aWZ49Q1G+E5B
TTmdJJ5Cncg2rpZ/Clc+G03Dq2dQ8Bs5RLLDf0lSMgrcWJllBSqit6bU9rwA
URmefPYtlMP/+iTs9lSroNHqXUHxpp0LZozJgtYV9ckuqr3eUmL9F8BTxfeG
zDIS6/S6j3ZDqn9mceHKkMY3+ZpAlFMvF/UOq/KlOiZAHMDAPzuQiAV2HYyH
Pqrn2S2+NrOFNYLouIQ05odmEQ3rsOPRSSlwy8vzmy8mWO0h5uodGhqf8DpW
xqnmXmIMdihmERnYDwjtYxhy7CZAYR+vtcJFr0yvLoEv/BlFQTU+dUbpOYZ0
fnRwTp1CogC8vjyeEXQW7Uvc6zdfmGf4MR6lpM7ldzpSFpHOuM/uzDxADnFc
izHCXLzAn1vhMOJXBGEjBdyQyGAPBrOoBHAVZOb1ZRca+NVYn78M5IcEGEwj
qBlY/Vz3nFXwQTmZlSwOGPmc+pg3mMyWsqu1IBehoj9lVNGVk0y4QxfaO8b8
BDIjvSqWsE58PklQtxqWs+Shmi30l3R2nSrmKGU2ISuxCCvGAk87yBCAHzMP
aY94Geeow12eEhHv75YDH6aGaHZrEUMVbt6W0bhWdJeq1zCW9C2ahYOuYMFX
BXFWczEhAjAmyp5RrLJBcvIHjqWAso2brSzUCDtbkG+SV6eDNKlS0X8qBTlV
Ywp3H9TXW/rP5lmAZ5uBw6I2Cn8+8nrWoX/HepQkUdjmRdlAVZsGC6PE7WDX
082QItM7UofPT7ekbj3fST2COjD9btQJeXPVpNdSPfJPS0q8cCcBhrVP9gsL
xjUxaF8Wnv0ZHjSuU7wDcmRaQBTmEVteDJM0HmllyuwCwb8u7JdI6dhu9+Pr
iGkApJ3ZgWS0T0M9Zv5m0g/TMd5gum3h1u6+LBZxT19fgsePdLUaGIWovcFx
r96n5Y66pR5WjgjxOuEsGsJ380KEWDPhHOAEOgPWwLtw7PGNfNFhuvYOfcL3
gw+NcVx2VbXjJ1U1AxUS9gb5LKrcmGxxWGA/KlS/tJrQu4xktg94qW6uF61b
3NcJWArNH/ARxRS2UVFvhlxm4MzgoYXAiSIkYjlE44ZYDrYIjoJAb19cySEc
O4dKF/IW/NUounHpc3qJxSq7iSp7qklGaikzR3sIwWrkY9gaZjeUBbN3+4Zy
MqqOkPZ87G9c0flzeWi9PSeHWQI89Zgpd2up50cWazsNFZWmDFu8MdhCDhaw
ma+tUtAzK5KXIsG3JTXlbGCuoSJAWDXR+zX8Wn45yoqaroEPjnVrkwaN2uKr
Wi6UX//SrFa95mBc1FCIwCDhmQEsEm3L5ZwfMN2vu34avOY0eOcweecc0OOn
uOit70pCkTzmTuK1p+/RlC8d4mu1XKJQew7+FPeJQNPn2PBRmtZPDmYE4wCR
lHv/hYwv6+qWUtDD88INHU6SI46/uh5GOKAhJzdbrEeIPju+YITgJXFHkwum
ORgsLQy3Q04XOFV37TahZ8FVfB0Hl4gKWa0q5RRGCK2A+aDcOcDjtzq37lJj
4roJGuS3iCDojX97xZ3ShBv1a7m8fiWFQ9FbuJA6y0ZcF0Exo+yv8dYU9vyK
ll0/mTlTcYhVn/SYBJl1QijTe5huOL78KM0nhfrj2BUJcwIhNBmTRSKlPE20
AIWHpFMbVp9XMjs7rxPQfVzFqo9Z23nmyZyfCHiXiE2SuGWWpR0hMDK+/W/m
/7B3Xrf4BQw5QWLBMEGMswWfCL0dS6TI4a6owCGjAeLd9yPnUaVbmN0SP2c+
wfzv46a1Iwmu7ZLeQ5QFVohFBc7n3w8fBByuNoEJQkNQyphxkrbTrUeajZBd
ZFP0l3hcEHVdhtdL/BTADi0WbsJEIrs35wiqjPrjl1gIFEQ1fSoSEhwNaJ68
oG3sUxll0oSaha1FQwyeSorEyqfeh/yPqT5by5a6oFjvkD5FOfhMJo7aUdrQ
tUJqAx8Rnlf5aAFP+xhgJbRQMuiG6FZCFiWqfWukYGAGgNDC9/6MWmIzSJOG
wbRdWIG5L8a45M28aNhdkqmq1Rxww/mQLjpg9oKBggwWn6G08GWWmHj91RRw
Ajv5tXwItNBKUsVX/gS5ccVtu3JIqgDb6+Bcwc/Gh9JVURw20pbpLvUGOcVr
ydXzr4Q6Lwuv89DCxJohvsmd+AUtiKxILfKuOiBMN0j6JEm46XdZAbxO9SLs
So1MXsjzf0DZgNVLq3NkbxBU6gBQO0D3l3fPN9XJ/cBKOd2Fn7s4cqNAHqgV
7pjox/AQ8p0gC9vKAybHgIiLTA6r8XwF1/SqVbG+A+P8Y99DTlyq6+tFa+la
HUrjoY+sgT8cw/hVD4oH0RKkKTyEZm2cnCnSwCFtURST01aN1KplEeEHteJ1
R77FQckR8iTpY8c1Hi/Wn0uqUzasJQtS10M/fTrqPHzeFybnE/kZ4f+wZAtm
8pxsqO/x5Z4YXkQSOf02TmS0ms5FF42GptcFEkKaqBw2E2pEk4UxsUKEVoEn
DFfTFFQyi25RKnt0pQro9HGQj8rnzxKOu+9T52WRsZaJzN3fbz7yXHwcMcvc
G630mvMjSzL9tVy1vFw5XMgQupyUfNdZkQyMGiDUSVtivD6+WJGCZfT11vTK
5GqVhB5meJkkpQzHqLj9qHb9UpqJB+goX+gxQz1PiMuBrJWaDJ5eTfwdCkBB
CMTbgF8/cg3Tz7S4k4cjY3I2sH41PvJyfgM9k6UePqDHn/0N6DHmrKvcXTOP
LBEO0Sw47zdKV2pyXx22S3T49fMjWS3YSLb0QVv0kM2iyP+rUkw8IfwDMet+
XKWPcp1xT+B/TR5EdAiQRRzOYcYUWuymnbZDeo1WIjKI+rvNE1m7riJyMgZy
Bk+FrwjQPhcbk4rV3MEd7vewOx0JUduJ6G16rsF/poBg8Ee6dkFSGOCS2mad
7VhSpH7V6Q10tfVgfVWPcSU4ZdJLqZzXSYgaIHfrp7K+BWIIsLPyLyoPtyL+
nzMUy6u58UgBXfK7NPm+ftraeB/tXrYKhHyqBRCXGjEQ9ZuTWZPQ09OQuu8h
UcV2dzQd85dBWOIRxvOI/EPCzl6CDHzSWYiBb4uVYV20ic3oFa5fMXOa5+Kj
RFMrssoLchxsWcUcMjotpvyBU2xL9u2e0GFXG0C4qgBsccMTRzvgpTnzaFAs
gK2WfgNnAQlTPDlzCGMSOopUTIeI2mpdoj6hO8vC9u2l04KLRCGBPyo5fhJw
O6Zysu4a09Vn5I6q+rNoK4gjds4LY3n1urYdvXpbwpn3CpuoKBN08Bu2tDD3
Q/kf+ix0oiwVaJ+9+mNspFR6IA0E6uTkZboghFrhV6yKCtsifxMgZBCum7B2
DzRgrs70fwJKnKJJJNJDnfM5Y7Ob7oHzzFWoS77bh2aNDrN0o5SJdqG6nNQC
uPyqeUFK0KMAWZnQ16KL1sy360ZwrhT8Rezmp50dWIpuClX+ePavSaDFnrQv
wR0BIJzvfWiIEMekh+z5wNvHRx9zXDd9Mmjeo/gxxzjwl2mKS2z52L+MdpVO
xL3Pm6JJSwMcGxZsDqLJJMpinERynasYgOmUzZptJlpUWUDs79b54FFxAm3F
NUyoKYLuuLO2OpwxtAKb1zDDMPOpRcgQLZsk1JiPrVxBgzYDBgoy0USZwgYB
Nd41hau845iLNZWLVtJJgV/f3PMuaP1uEbDI2ns2r0OZpfKyaz8qexBtbqR3
RJpwkeeTQfzKXmEViFwjk9hA4QOmuxfCpKFhtVgo9vGis9lV5LKipWwneV8h
R2O7sgKp7gWtwp8CEAsmAHzP7p9JVTmlmPrSYKiZKujI1v7OYLMtSzGjUEnQ
rZXtMhy3V7RVidtusw3Bn/L5fVTK8xk6BFnqAG83g3gCq0yS+L//pFjj0Ikj
sJvukyvyQhcCFtFEpoCw+kyjFjL+WJzPOeFUA95UszxZS8Cq0Nc2ygtUC3mr
1xaZpm3/uxXd5ZoXFJ/f2dlkxFaYYs2BEMgHILmmcJ4sKRs0zi3VBKA5Y0xx
OaYML0eLqyRcKEB6pobm0in/naxO0BvlcLpNYmViGH2ajnYxVAczV4LP9Jyl
BUUGJ8Ckf0DIyClQ6Uwd/78p8PUHGc4qd0H32QePTL7p3vkSGNAiO9rgcgHl
rBpXndaqVTZGYkJRkWz2saIECf/qwwt60NP5lR/xCNb9/uZxTA5YiDVdYJ5E
floq+IB2AGBXWBjseuFuzU0p4I6hphEF1lar1d7b9QdrcaelFNIU0r0O0Rty
PVlP53jgdS068ZV7IPzSkob6GHZ0a4k2lnzgjvERiKA2JzJLwxJL7kV58PCO
Te6I/n1676tSCpcaQzWDXzKo7GOBZdVIxwM+EoSAQBbwABwVfAPdpj/jA56N
HvpTy8sO9VeIfJ5/HMccYaRhwQmgZJny3wPb/XR56TsbWSPm+C5OEu7riJQf
MiVeurirThBS3+MYTvSJXWCaWzbNjefWX5hP87+Xf6C/tryvy9pSA6WSjUhy
kmUOTCXAwYw/1C+fIMnY9ITK+7zToddO1kht61nw+fiOHwpD/z6wfVitGzaw
1PDRR/dy/qW+eH0Bp8YhoGoOjzj6NbkKGkVA1gtWDehUWZ8GUAJUw6cAOCS0
0z5W4G5oVyxhvOmIIGPkokveijaRj27VKocNEE4KFq+xsMuOgxbRnDg9UGbJ
/9e/Qd6Wo/R98jLMwW00ogGDus2UBB9ZBxxC8J5OtVPZiPgD5msHAKTGMXA3
OHf2ITPGtkSyRxGJNrRP9ZHLiFyfYO+hY/o/pObO6bqitjHEWpODe4y0Mx7c
gX44Vst6QVTHe+hR2EIg0Nb6qFfsLUeH0oqcqKz19ghIulbNsInxraD1YMKd
neEqXd6kN+Av5bcFYkcQUYcHhn9zy93FMAwTfxFVPk5VDbRf62XDPa4x6RsX
HSjPKfY38b8gSEASe1sN205HjhVLYb3pHqibe/rdxCHstQiVsfn1n+gawKTD
JA+TnuP0JYBWhxsmhHcxBGtQEHdnK1+0b7V9M2WBx5CJI9zXaIoprL/ohiXv
+CMSGNKlbk4hh3OTyX8i4TIxysXUQiip8e9N4NGzWfipjhbrzVmUEn3IRl71
daEUfNVcZjoUWsYILmBN9AWuvjRlysbwd8MRtj9O0HYaBF9Fx1nq2YQerRb+
L8yEu5BxKqg7ujK5tp7C/2vQ4qWx7agkyuV2z/TmEjm2BEAR8q4yqdbj+El8
7pxy6lRzoa5XMCz/4dHRCORF4Ji/KU6LobD9H46hMXPPRFj0BADt10VhYBw/
ynJosSIzEJ+kR9/d+BPz+pQi28Xi5Ph48g1Zqz4wFuOmN79PefXP+TMk+FkP
ntvD9aFQRlQaGg3hseAXzlfZqcZ7HZa6drFzXTBX5AIQK6CCTdVP8qlk3am3
t1z+guOJlS15ASAUMPgVjbHgNKLZnRh0hCCKT2OFHXuDIofj56p4ryiyOuFG
proOc/zQEyQis4u3bty47MMq+r/XVnksjU3nC7nXXVPCJmcnT/kWXvVBPmb5
p+juKR3jajIq+2FDOeS0EoPFwoZp/BePmDLDUFL8XlVdh4mea4sZ4KMxGf8c
41nU6ufWzEe2Fzzn55y0P/WsgqdoBakJyB4ZJvhIPYNr+oOxNZlPX+TnZjRs
iQfwLaBagFoIxFSLcj5nNgv7VE/dXhZO3z9cvwKYJ1E80P+yPFVvxhpghSYm
SXYWFLaBlDIWpVBNavksDyDPyyC0YhKGGSI3UVeHUQAiLOon8EUMtHLNDoiB
sgL99yfhhfFT+odRGmH61aYQyJYMp9IA6cbgWwcLFqMzL7dA+KwBePcGRZld
fsn3h7u7uHyLWkouH2tzF5F2nXfvfxPMYfHC5Rxp/mx3o1Og6ZJWZVTpgUxv
hrAL40btclwQu69eePsHezHvvo0Hpg9Vt+7SSb6FCJB1oelwFtKJ/2GNvyDK
unywC5PcbGgibF51nR5w6hDxPn+F3itrk7UFoG0Ia68y2OX/Gu/Y8n91Nix0
UnZmgXB5SQM/F7k41WVI0H6gdXorQbKECO6AEqKTLrdd/cEoc0hkJlKW30YT
pU5XqtWGHaEFJozM/No9D6cdojrtP+TPPuhUxLGpKxtNw0mAEFBu/ixf2Sfb
N6UMqt8N60yGWn14z7cwKiI61P0f3hKm1hsvRI0S2zq4xNATQtWAojp13v1S
uotSGYNJ80OQLRRG0Ej9fByYYKUQWsiWEwPZMu0N4Zk2QHEE93SwgYiMyvRb
Qp47FhrHcYS5HxvbaApBjjAEviyxEkayXcuyJssvJtVcx8gI5riQS3Ed5hCm
khTI/xDNKAcDGGRFqpiu/d37vW2x3Sbf9wbWA0SdT884izmhmVOXHCHmdWN1
xGt12dazErapKZm5PrY2aNA6SnD8hJ61WrtU7459I6aCukLXFpNbYyBVa+i8
QvDIboLwzVDB++vpjAdxKpSMypRpvSf1G1e/vU6qGhLN/A/3kLuvyHYft+pl
MTOu/kMyY8tdzBFqQlzayzUucIS1q9H44t39pL8vqYCshSavKvhA+KvPqSg5
SH6SwBscr8e1Vl0XqWOmyLTJRvfvadPpuAXXG96E41GpELPuVf6GXMOSiPVe
ymDHlNqfWtY4kDVM5q/f/9uI7K1OpOU3v4DiR3kkD69qaSVHdEOjghGDQW1C
pmVOBP+I2tWcyCCFRpiyURqhr9tOa8coLtDCOyWOdmdRk1r0xILP703faUGc
rD7clWzrKfUUmsnFFXIXD0lcROEV+eRq9vQetVAxv3SAy1lvu0IOYxqxSEna
EsR4h9ABYy4en7eRgIvdzYVWBzYWa3KMSRGyVQzJPzUp/tj0CpP9gyvhfEq8
yOLhOkQ3vLGjymFjgfxU8gsPALn/rQLAUss+DvodcjM0FmVJsv9zWXLx6kI6
m7nt24YRP1DZYyWZgL+h9SxkoQaowi9MNrOIthHN9x1/946ICptTS7qa9CKy
H0VIVFT0RIgOuBHHJ/loeLKGdYCrdeyYyDyePCCdrFtRTtaPKM/EKe3Hs8Mc
EfpTvonA9sL0Ix74JhxFqLClnwRXHx7r0LqZaXI1LRSscOUO4MPhab+amggm
sPbVzPzYCKzvrytBl4mT+TnZcgDfB1IX5eNX1GhtEuPTwzqbjH66zPy/SVqS
57AHKLJdszvecAlmxAjmQgplbQd9GqRlA9Q2FvsavJielPulBaA7KBdZBHnc
kjzSXs6+7Ph5I07Li6oJTEj2J4PQOkg4SAxXrXQawY4RQAVYOw4RmlDDLIba
kvbRDxhHKXJYcAUWt4l6C3vHfC3OJFy0Xo4JJHvqO/lq37vBjcl2H4siI5mp
/36gfpe+uo07M4dpMLD74AG2q3SgPidXJl8g7H0LGpX7X8JqUvxCgQXMbLHS
5g47t/AeB/bX8hHBmAD9mjpok0sARNvzfCjlbDx+Z1PvpbrNgpDCAdTei2n+
N8zj5SKm3VTNw6j4cl4Hcoz6b+M0W/KizQN4Kj05CbmX+h0cWHbE+q/a0sVt
Moce/Ds3bfVw/d+8w2J2S2bhCrNYhV7M5+taHepbIQCfnU0q56QHj/4caj41
DmXyfdL+W+BX3J3gClcU+YvO4mBwyFeFITi2CJGdgXZJTPUrD+VRofll6bv0
XRPf8scnVHHh4o+H5DDKJUhM9pOVf0/udw77Wp5bCDov5fchqeOzg1KPBNoo
umWPVwA2LVyLXO8C+Xy+EVcp+3q9uEWKWwI5Qf9J2av6CqQvT3LzdFJ3fMBH
iPtaHBRJwxfLqyWvTKBt2lI8OwqWKuxmpcopgBmtSlGZbsSGNkL6mMgOcXxP
WBGMqVcxj6TPqBFT0yWrw1VCb0T7abAX1Tr7pVz1WQ2k+fuwtjKh/5zh/Qo+
GSkWv4cDuOB6sAShxjrgDL865vviSuPBn8vTArBOVVX/bgkJqLUYxJEpKTPe
b6aNY6N4ynlecemp07pBdRapNK5CXEiMyGtud4sD7AIIt6A7V67oCCx4Uzsj
8vOleDZ1mPVfGDp9dPEXy+GLROndCsshwmOGS/JT3jLpjpd2GRURZGzn3C5W
hlFhcjRWB9UdBPhUfYtwg6sZvwabKeQ7nEF9/+7Y7YZVU64ZRsnIXsppwWF7
vctlTlPoCkQ+5Z7OyuiRQEWgZQoJYvkeyapY6nqLEJUcqe9mQpXqZlZB33IE
/z097DOc7xvpDioVK4IFIz/YkEgJvT9k/D15g5oM45GWZNHtBodkNY9Ix1qF
tInkjTNrvUVw9dBhMWzqJ/5xXxmCuYnK0BEINjNXOgkUa/k3sIHehdKcIWUz
/CFwxdgmCCiRXamkQuMvcRKnbvJ8yT3wjuEK9yOOW3G8PuxX1Hh2NDi82UZQ
SZX/UjjAS5Yu5mT7gO/a2mYA7F6YO/R0v/9BQXuUVDcc7zvZBxxZswL+Zae3
K6ru4lnNdc3HhcZSaPC7HjshX5hiVUFhbTsrIb1YBpq65cyFqKW702feI54+
KWW0Ne5pD/SOPfJPCLJnkgIY3JzQbAtj8e9DR9Bqf6X9TixSo1wnp8LWLKt7
Z3iV/bMhQ1S00mWCPooyKe+HNfl3zrTRpuLnPqySURBChqt1g3qkSt1p9mR1
dn0y9WeMHuViZjZE7DMdWLYWBVHukzvkI64P8u0yTn3+JtOMRx5njozm4QE7
bROV0PVG+5vDymdnA457jxiYxaF7yzp3UGD3VpCNJkcGWPI/Sh1/bfQkjvgh
qnQzzuo4k7OQSmIZ9RvTmfsT/kD9WmZ+N4dhHbltl682SLXazc+yNemyl7V2
58y99YlunWMGg2hzexpmzuJOv3HthRAzyoxyckaVrzvtX5Z1BaDTOZ8eLu2m
KeaqKb38ixM78m9VX95AVV4gUlhNM10t8s0TL38ZDPodmqzj5GrXGaKVanqd
zM95aPvhUH0ANFL5T5UFj++hmD07OAyZasG8oi9yXad5LLLRNtc1efaj8mFf
NfXWjv+hvPvg/DULBekwqwIGPuZOyMZTNrplpZIMFATl2r7d3An1W5o8kEEs
OHKsL4USaRu5b41JJYb/MvAVj+CAHvjNNzFT2c2epakuYd5Co/1THpWnI3su
llERYWyvn2I4Pd4u16fkHHsrKuiQpau1xdehDTUOKbd/r2O1YYLuJEvdGzHx
6DrQFrB0Yfib7yGROhqLLgqarmJKqzS6M4aC1J8dCh4g0LbcyvFPS0OpM19x
T+dTknc0Ik/gmenOazAsqXvLeffuIgW2l/GmmdO/cMdilvWfFd/5p+tIZLKv
TtnLphNGPw573gwilYdzl1CPd2atPpMzNAnP0YtCELAnI6mc0qRVxr+D45bV
2puF+q4SA7AGQQApAgRVXF42er53OtT+y0LZlytW8J7Q1y1YhlvBjP6uH+Zb
kNpjdlW6hvK5wgphvJJg7ibPdQccXmTWj6a8EjfQpiVLhZl4h+3nMGYJ81oW
yz/jOpSuSDcqj/NCd8+pPOSLrIP933CXf8SBkFJKpuMWiyONVKCArDlgwtrO
nwG6j/JOBdf/qPBVnzFTG97OShgP1ms3vPKjZ01GGgHYyagqTYuuu9W5VhGR
cqOdma6L/pxZHVE1jNnJaBW7mSv6xl+0QhoNYklIaHN99K8Ztx+pTvYfeqwA
FnhF3qjRXg+i8G4QvblV2SkaZAf7th9Uc+CCTFHXWPpJPjFc5JmQWzExFIbZ
lQ07eRydXPnwRAXmKy+DVwF+5/eY4Amzt6TPn0XyecOlHvtztpc38I7enP/w
Mt8ZDe1rYMpSxsmWzR13w8Y2P9dyNJRQ6XsSgmn8tXYio5m9GYP8otbTfmqw
8gX1uoPludW9vemY2I87o/nov9nSACka8in7aOhrquDNKN1fBws5IiEtnamJ
OZsGavE5ZCdhXUMKDHe7ADDEGKFERbn3Sw/aGQVEuUCV6zB2YKgHcj0f8f5M
7elvKDwYAqd3hXWjz3sSWH8uonpcsy3ErzWnW0Dxx92Wbwn+z3QY54mv88L5
v5sK51v61HQA+QRvq+do6ICWMksOJaKti2MdxB5+7Id8WprgFQbCaS5iaVLm
l7DHdxsQizzSTANlN4X1x9IU9Ak3BfU9s0+tOD/z0gVhMBeUHmvdL7AkE9FY
8rtUe+d0CCa2vARn0o5aHhFPCAIg2j3PEa5+3qYyKn0ntbHf9tF5+PqHjyjl
GwXD2ZOjxmu+JCrHH/LCI+DAJEL/CyoBCCFQlrpwO55pI66/D+ecaoynt06Z
CgcH+Xdzaln2f5pxfSpKtesoL+Ty8T1onauK49zF1NOgCHi2Av5BRq0hqZpV
0Pim7kp6/JbLwA/P6c40gALPdphe6w/Aad3UNedob78j9c3PaNMJPRMU8IJE
OJ5+Gx/UxqOVIE8FMHeBmgNQkfdPub+5Vk2fzzidWuJAmCitgjvI13FkURj8
h/4PH5BxxqU5X5vS8geeKTbb/RLmEen3rsG4yA+4tPboQ86v5NDqqByX1TJC
PplNCmhY/h69XgRN96Mh/gr2tv0Jz8YVyLE0MfDx2wShZiXmLp/+hEaAWO/2
9SCU7mP0m8VczkAJ5WfNFtcJ3owa6X9aMDjSEiwiycWpwTdwNT6EpaYW0AQm
HOl3DGISsY7J0BeiwXeEQn+qK9xypAt3KbK0D0k4izc4thCNm0/WL7mPwrsb
ltyUrsayQ/fA9BvUC85PKdr59qIXH/9CE89T1Jo/mAlh824qOVY99DuSIy5u
6I4lXTuFdjb/SdO/RebSU049DefBQRVIoDnbFnFrOtfq1aG7rECQQSFophCF
frhB3ZLPx8YhBbVy2egtm/inQp4x3Rqg2yqcgO5VQ2LmhNLQkhWNdlcunVXh
3qPKqzseKv0PQBQxn18xz5/UzEdvt828betWl7F58/gPVKiBqTPpaP39Ky7Y
tVFZcgedvrlzAQ8G/wzLGuHVt/qaESkF2nmFPQKht28b60yVqXa3qnuZlVUW
K6d11Ta71Eew0iUncn42RUVv6A9X2uFCFHKD/I60mTDaOSyLylcD0gORi7GM
Fe04YdL/lykLtIzdwy+/kIsy3MS7UgnShyNGK9Bx3f8EtqoXm8oqS3dehmXu
5nYmkiYMbkCRCNqW56ifcQc1b7+bIBEzgH4L6ZvaWzOXxUVHP8PRle2P2MFC
8zANAtP7nirwQ/Lk7MK8BOH+XJxmxer4S/aSoa9N60EiEtjFbJotwKcVRtP4
V6yEtfgjyr/GVz98XxS2lXH87meAV9oWOEAkUuqUbSEUrBOnuwsPV6FiYgfX
Z999xpzFmrLkufeyP4smWRmSzBEOC+7IMDzo/GXp8tal0ZfoqocJl3emybMq
omePvr7EYb8lL32ejgiBBLTLakEsW8jvJ1KYp1DESPMMhGVOwJZnQMjo5wJn
SqIW1uKu5dEbP1lPxvT3Hhpkd7hEyo4ueQWqZ4t3bWmkfRl+PAetp5DNfChG
n6GM0DvE0xXx4GFZMBLa9A7Ejlu/cUwCsXfZKMoQLuiZlBqQe0oPU86v1Z/4
JUJ+m4uPLKHvnkVUbKxJ1Wlz/Ox2cl/UjZzOJKyxZMtN1XsWwt1u0Ar3viph
G2tRUGCq2I0LkCmgCXrwp5/Sr5BUFuauaGcjHd+lJYaXhafAsfiB2uOIXXui
WnYQ9682eaM+yY2zuFU4TKw4sOiDMYEUk68PQb3j4Qz1tIUt+HBzoKI/J3Bq
GVb3UcnTBRDYlsbMw/q2HysTWIJiMzDruw7vU+oMxrrG/ZmsA2SiXpkQPxEY
bNKgXcXG1sYS9bHTmFcLCEM7CoFZtqMrfI2BwxL1N2PJpn6QfKgOjmwwmb1G
PDw0W28n3x7YlHuDFaXQasGNoGV+7D6x3hUGKEEx5lBU2NjPinOVZE5knvlO
wfS0jELMDKgFikz2nsTj1c7D8TKl2LUCD5GNf/x93T2PoNyxcSEsjJpJpLvC
AMLL1ztxk5n9KHtpJkHbcXwaS+TF98x/JPA0/zvY1GQ3/HzuaHjiSh3tRnBr
rCwLnhkSqGRAuURkB508/jX0M/pZidKcSMwLmsAuVl3MQM4iutBSHwrEIgVi
AQ1pVZjsYC/Vy5fPXISL6EvjZ/UM7mqx1pr7Vc6Pu/nYMNOz2uFtj3k4AF/c
aCIIWydva7KZ7khjiz+Dv/6OBbMmRZi31ty2FSsy3LfpcqZfGh5Lw4yCemy1
lTQQ+O05JnvqpLvI/jDWl3sdB7jXJe0jeb3nBY1l1E7djATn4fjnVdxmSnnl
3LCWgY2lObw4FAZFLfgmpR/fCTAxRuN2fxzzciPhKeUv74Fgy/cncEPatyL2
BaYevKvA8Zx2SsgT9tk76PDPrBWoCqVv55XEcL8TJiAafT6ZJY1oehK2slDv
bUDEo1ab+7/PPN25KXBEegmg+X3wexXjDLVa2qb3tx30AX1EoGqMeShOI321
MMnVlm5KNFP4jO0FteI5Byix2ee7GkcBUz6E6+CUO3dwLoS3wnzAj2x+v1Zl
AXr2u9mzeqs9JkSjP/2ewIKI467CC6QWqPv4iHrlFhgKypKEaWBNVcAy2Y0Q
LmHfAfJy1ZwBNk+bqwZO7w7ekA8kLaUx0CaKeMA+bxSDYjnzmwjjT4yP32pK
ziJju6s7ZyRaYQ9g+P91Eq3Fw862e4Mg+e9Ip5Cx8JKNApPOj2GPGdYfhR1b
a2eFM8PKp02cG+0Ga+60jTspfmjsEbjl3zjaHGgy4yoQ4u6x3EH43h8STswN
g7WJpp/L/21F2MWSGxHuUtfEW6xpcmD0yrBpzZB1jy3rdnOV8icWVb7cGegv
cI+sT/VYd6EoWwx6pazzRb9F9SoQ+FfK+7cwxiN1F6K3hx9scLXQ2nEQa/yx
+KAZOSwkgYPBFf+RxUHX/ufSmyOqWE4r/ZEhNmUiA02hcL5fy2DtBUxplLf3
ZUq1jTCGQq0wtaBRCtq44+mo5+WpYNZ1Ck5edvf8bBvgScqlLBXx7rKKtC05
MfBxQLHIa6cY5gEI9F1A3q946ruDXnhsFETwNTWe22YH45GbVXppX1eVN5En
gHqoQmGME7NTOHIBCJpa8FN/FwgsWOX1PpDNQ3UpjpD7JpkajPM8M6yBHq6j
X2vrEhKZ/otIyLINWfwJ3LuF/SqVpTfGukPCkeSczkgtyTxk6Z5/PuH29ebw
gYoOCt9i+A6HxVOSAtBMBvZ4yYrQrclpln5bwBWAEIY0UsxCvLBOjwhK9v5Q
ttTws2ZRjAbHWaHCca2GwV3/cx+Nc4xIZcXiOupFwFkYOxAxZRmU+M9opKUg
h+OJEy8uWf168Ul2fiMp6lUzbM18SXUifGJU5TP/o+SfAUcFzwiKnMKvwZAT
upaQOpWgodYkaTSvRceXb+vmJ+sPCXJf66BmZXJlHr6ce8MvM7nUa4+5sy/f
T5I0vpOm1X03OkgBE304ATE1RDPXPIyguO3/WkW0oRoqJa2pbVYoNkImhC0I
B2ajOY+zXs63YRs7p+NJUbjN88/EDqhGGB2wMWJ8ZS5UZdEWAyaoMoHT+p7R
S3yuN4RXoKJIYgU9JbKZ96KvOXUmi3mtjUldnI0mulXZZk8knvblRL8LvW6A
Y8fDYrN5LqUwgHIKYXVjplGZy06aJiZ8xXKuw/TqJXF5AhEGE43X9muAIXD7
HOjLzsTlB6jZiT066pe1yVHZMNzO0ZvdcnJokJ9wX0GfozMcejPfY+ccvsW0
UtaMlhtpHLy0gCgLKW8OtxxT9efD2z1LklzfSlu7QnewRmCXcUoVVmPvaFiP
EgLA/lsjSlIPWaoafUxK813Q5eNwk+5TOcTHq27igCKtNQEGpSTBXHZKOBtB
lZKtdiJUZikd7148gOmZgZBVh+oao7tcE+eMY2vZKCAE5fc8k9a8pUiEopix
jWtsqmiduiTufKqeublnqcQeJeSdjO8lia99jGoCMeIe8n935tcv9Wl/uu30
kX5SbxSSdRXYaEXnxn3Om71xABepASHlwto8Q9WgI5v17+FP3DVHYIfreUpk
ViExo5ByRp3jE2DQI7OIvi0Yv5Ukyjt4T5YjxJCF13DNfG6ikJAtbnP+FAjz
kUXrh3bYos1mWmgNzgL1oXPSpsBbpnstiYTWjjltLHpXX9MPCwcqAWfjYW4g
uiWNh6Qy5Gs7o4igltklBxtBbvBfHL1cdTTU0OJzTJYOgJW1s0yOCybfiNkJ
cri0XOJTVU/Q6mwEq4IZW79tbdH7BpS5iWjRaDpTCVCZa6bYoX7uySdeM3Wi
xDUO2sl0YzXt0dr3rZopZYTWVLeJMzWFbDW0TmeN//hh6oCghSCS2eYfk7BM
x60owjQY7j+t/jhrZTsCw6RLTq/0A8tjSCag6YpX/dxcz9zsTvtFX5e+UaRG
wvqoxivELy5T0R9NNfF4SHnog3FLYt10iX2GsJDOCzB4LFjkSXmKtlBKGLy2
F8qcSD5aNnh2MbpKOCSlM5HMRVDEE/sAaplgmL+iCbiA/Zap/PcqVoU+6w0+
VfNJp0EsJISaYUIORaJsOAbutlNnyfbY+rVV9NNCfMuyX5cacBRCY13f+GvK
+8piLr5QF3s3KlttEmwCAoxTppNSQ9YQDRQS7UEIhpkbdRQV+vEdBjqilfAr
J7Jn4wzeJ3DCjKOcoNlVx5SAG2F6P+Ea0yB2tz17HrW3vMJMW7D5A2EnmTJx
Mh2YTaNBgc80RVK+ku2ltrsb3EKp6XEpIGRNUCJEaGElgecdELC9iDxx1EVY
PqmCVtxWWJdFQQibtTerndE6MqDbOHbvzN/1O/a1cUDdWLooq+OS5z+yGF5A
wiY1njsvwgY0urdPsGK+YdRqSCthF1LEfvYY/YVb/GpiO3/xhpmiAfhHozci
s2pT3hLrvZgG7c4HxupjMuscb2+I0s+myaJenwrs3xUp99NDwZe19h2eDhrA
vfFUfvLC4CxWmANUrqJ6jBGYh8/WbJA3slQTvJCNsT+SzJ/R12IJmrufjwdS
Qthq22TNOiQhTwu9xHjoqB6YX8L+msMYdVitsRhoSuvuVrnAyPPTwe6aphW7
7nM/1frZTuoWowKL2ghe7aktZ/yyPz7S3Lq1losuROEK7ohqgBRguXIAM9T6
cWZNGHErxKEr1QeEOeE22Iihtm8C+M+//EW/Ah9BSYXxTSImGxT656sllA6O
V+TlYPmGDX0ZKPjwASOerKpTZFDi4ODYkKbEOPiEWnxRNE+LUMLYB/rs3FXl
753SaTnYBz+oba8N7eXRlAw7r3NzP1WiLEK/8dkc1HIuumc82Agk8MmQFijL
Q9lFztvyh8wPyLMUWRRCgb+sTfaTrln2ec9OE+qydfYIeu93Sxci6yY/z3CD
Sprij1UI44YrLOT6AvnLoh+sIALkfi49n1yE2Kiw3GaS4AYPcx/IBl230mG4
Vl4FI+0eZyyKd4b83d8mcoPFlEDPnXQWAITUoA2TUjZ7TZaB0fnOVRPB5vCE
8qySUIr5MAlfP9Gy868r6Ba1nNgPt/dHHsjkyrTaN5vkemxuZ3kUQN8EHKG4
sweI1mF6WLzMPeobMULHASWqU/5XzA6WpRuD/2cWYaC0qe96iCI1OrVhxkPx
lPhrb8oPN9ZzsmB2qVanbid7qamSlHq/jOsCOA6uPyQN8g/E0hBjATwJTp4N
0W9yxyk589+cy+y7H6ZbZ1z3DftMG6hFpvo0JBMFLyg8OT2bbqeXHB8JdpLL
H7ejsnBjlaEDFNXeWOT5NCnHnxJtDf9ETrjnmG/fnezB+ZxeflAgro9ODEiD
EadVEFukKplu7+Fn6+DIxedD8WfjkWqlWs/r+WRYq4tA4bJcUP9DWx5NTZCh
k3DPFlLOuS+iLbevE2/noOcamgU/b0SDz+b2mzROa2o0Lh5rFrfBHf2/EHY1
kmiWU9nub5YTYGEowamSpvry7ka1SbhILW/uOAA9yOQiUHcaI3uT9G3KOB9l
47/TPsy4FqsEnXjRFWFjcyMwosO6AAn9mc8zsSJrPp4q3ZUjPZlQW7wEyWP/
M/rGE+ZIeRuZgCTxuqOVZWD1zEtCankb6s+0TppdAwbA7G5h2vTKfkKEONvu
f706xFdp0zwRsMa6mRplY9bCglQVrmlKgMkO84LbgsrMevGx5MV3HNtnE2ui
9yDDRZopSw1jtoMvTmxwAqV9Ed+0hm4wekNchsocRjNzeLSyQ4pUZkarBz5g
D/UfJBvHguFcNAvwFZSj6WDQer/vuvs2JxBVwFnQx09XGv6TzH4Oxq2dfjwe
5xfFmfTEe/gHPLNVajNK60LGUjW1EwZOYBUBD7D/ijtlrJKyw4qJIqImfmz4
UHpDXX8Yk3f8Zx1lTyL1k17CPexiiDuzzCUj49J0IoesnIk4PZo9VGpX4KZz
sXnWyZmgp4mRGON1XAIlU6Za74Hyfga3N12zpQmsgKYlMVaUdr0y5D+ALGKy
KCpxIOmETHExCfnxRkHIUlVMt6bm8xygJiUf72f981pXl7cRQgwlZGPA8H0z
3/8REoWgnWTrl/rS2paKw359cEeUmSuId5Ia4RjzUaOA+NbRJ62v/c3H32Eu
gq5DiDPQZPmH1AKdbGhiNHZW20UQ0Tt+UgCFKmg2TnHOtIs+1vwyzpYcWLl5
CZIntlBLaZZCJ+EdFbBlw2yXaZ5KpQQzSjGTWAJbmrPDgTyoUVHLmXXfys5f
wRFOqr70ODHgN0Kaf3r90h4Vz6BAS3mwWM2eqNQyMIAyKG4yB3tDXRt6w8g4
yUdC6ULMQa/nry7NE7betrZOcpVjIO4bsaMlp0tQ4QLlqgpPxJvh7Trzk8ju
ubGka75WhvQ2WtdTkz2sHWZyVAI5xvGPfNEU+gw2k93tcwVbL6eddW4bn/4w
f58Tp709W3zBPb900ZOCo+jJYBWsNW4pxgzAQwsmXy2vNuqnquUphPAIZUlh
3ZtDCCh5WDqdnziqtIjKZ88+ZtBaYPjktvkl8FOQ4NEypDTgy8Oj/vhX+i80
odWyT6lwTDh6E1RIdfRhabcJ4T/pajOaoPAR8ODTieSTtIA0Lmc3xhT0m0Rq
5l0UAg4lAdYy8zQZje0eyzmrvqp2FUMNyr9prjjeRNiVsTde+AGoiUJLaFAK
+l/BUY+6379PaPNW2lVVOYpm/+GVt2Krd9Q0XII4jaTRPLc24sA0algwFoV2
sahaHzGyBXrXMYlK4Q4GPS/l5LfCwV0h0aBQwVKKdoVEF5oaFgN31fHZUyga
TZIrtraTpYKJw+oNskr52moLo7ry0zW1ZL36GXHWpZ1sjAjunHfSONh9gBBV
nNdrtkliNTDtbBQFcSwNfmHK4PaeFnBIiJfd6VOWPZWVzjIOfFQPzWF4jHZX
QZtMAbwW7+e2dC5bem42VQgZiovX/r4JlVRYdycFt+om/oX3CaG3KefceXuq
LXQNRzbQToQt3k7XqB8YC+UWhwMP9I+OeyC4BbCfwA/WAaUTE7qzOGfksP2z
8Po59wyF8ghcXthQ4vsxpejMmLQBuzZ27peU88jXumyxjtY1fZ5iQpyPJMfM
lnn+MMYwX7qDHiKILekbzrZYAXvMrPEJqm2hXoeGOAdqU/p+8FjFpQM422he
Wj74td+TcogjZakeO34gdcK8rvpSRS9WuhdQiTdhSFE/NjVS8KNgT2HBa3wc
nITeoFM3qTKVoUdcNvmYetVZjX7Ug3HNc/uLjKwy4zj1i6+xfJWvsRYP9z4T
1ma1ieui857GL5OmVTL97XqR96hcoy5tJBc5L0dQHfdIg1lsFwWR0LJ24E0J
SGfbq++zMgpyD0qwo5WWMG6mWKXeazWTp3ebece+dVG5blD/PznOH1AwUiDi
AQLa9kfpYBymGKF62Wx4p/xche8DHfdQF1Nbqckr6xGj3fVBOTPTzcy5G4M3
5Q/32KjqzCmwFLXuRoG2Hh5Hzv4eNyLj7sZtospKybKWJ919P7MNAbPUDiIN
z/N+DZLLg5LWkb6iK9uk4ti7uDxt3ELcV6OHl87sWdqKYi3v23ASOT8zv2g8
Elkivqo0/1yyXhoWwJmTNuu2GXVaNuYg4VTAwbc4WoU/TRzwPAotQN+N9Ygo
g5TPUl+DTuhohb22oXAzhvBSOo2TS7vHzPpo0MLKYDpvXgiYB4X48NnpuZEK
ZgqDewQWmXEB/0BWR36PmBNGsM63NxftkBkX3IBfTxT/8GdcP6qGTM+3fV4h
PIowOSk/JGtHPsFzTjiaJ9KlsGmp5OhhlmUlQVr4cmni987AZFA+mIu6naOB
DJBObw1WQYG3sqg08Yk6MRJbvgW8CaTs9Hcy7LqsyqLqOQqlr/1+Dd5yVmxq
Js/AjmmU6YwOGVRXf4iNEe0LBW28nkzie91NSXbiS4e2pZDxeVrAOkIBbBB2
sVYi/mhEnFUYHpjgvSN5+I3eRHL+SYWUTpfYp4Vdekj7gkytsdyEWiAGeRld
2wjUA40jPSqy7t1tY2uZ7udlt6n9huSWXXjdHgmrYUK8oziRkL1vqxq74EGI
rLIerDwN9n/ti+3QPV/shqjwoMjhZPexe26r5PYcIkEDRf5KvNSUuWnOKsWf
s6nioLwz1ky/gHvIQlzWS7lXjLuCN28wt/oQQ64CPvMsE3Iy0ecEpa0At4FG
bXTWcCDd8U9qruzziTgvC7izDLgGiGzYwyxOp3tAfINoylLdjy+A+X+m8EEX
VQsh4sraV4ISasnnSZeQSD01qCesEQV+A0l7+66rKHw2xIgS+RIq646duqz7
s07z88q7efK7593f4dVRvkFm43iDMX2RvpN2OsnRq+JYZUFOusW3Z2Vh/l0G
k9o5aDJQe9gCDLfCqKcmu4dlmdeJfgipyk+CYS0t9ErAkimHp/pIxGhSxRZc
OfIK8GNU0MEnZG/OOZl7qV5cEWsAbWjJB1m3AMfVIqGgFe88pMnusCQfaiVN
6whKiZPiLDia0ik4Rrug+IaB0srW13c9BnFXCVLTD3hT6Qxor6cO7CXwWJCF
2QDi/RajPFdXb/P7YI9kpsc2y5IulHMSlne9RHA/B+W86CCxxC3QTwldq7rx
st97Zwz/tAudf+WzgahoRubCxbWFefdlYjkOzqXCuHVRDSznpazvkgZf98qa
qxN86xtqQ24bXLBlhjezqRUbJFnO6/PUxDixCWYPdmnwKmrZB/Htc82V/shW
Pwc0jcyLumksfhSpRcDBDCAnU45p7H+/OAu9xozr22J2xQCqwN7J0OSNo3Fi
NWKui5dSsuhW/QVN+n3hwnhakybNcRdjZuW41OCHlB/h9+rFXcV0LEz8ae8n
PgvosufbsKJHJEMKxYNhhBS9/352ef4HPKRRBsRuNu8/YlAS6YbESGgiimwS
Yno5Qjk/yPqqHrGLFbhj5jozlWTAwzB7w8vfok0HiSpe2GJokWQIZjS0RGb9
i0nBRtkltkYb6/EyQkNzbbi3o0sdahCXCKYf1d8meuatcFPeuhb9uJNBx8zO
nQlcvwlyaDx8zNDTme2GnKb+/iAe33P7B2sto7qYAb9TdAL/1sO+4iE5aLjh
2rSpgPKqgurZvLpXKk8S/u5l+g+OxQJha0trJd7G1sz38vqCbwQOEb8oqwVT
AXXqiVBjZ3h2CJRN7P/NrZbggj5V1AdQCyYnTFcJQbpWE/tzURDQlD9hGOnP
owfuYZTEkS7nLHhNo6rP0aSGw50DqMEpo2x03cpQCa0PAJirCqPuKvyzXFx5
20BGnmKDiWpoIjkvI1b+WzFAkk7u026fnywVsRi6wBzEN6Vf/1J3YGeZ+UZ/
AD+UlE8Byl8FCR0eaPhNSvFoHqk+f/nHr6eaWnTrzWrvzluymynoGw3m1H0x
OBYopr2awJ6OwS119/RK3gxyU2YjJAe5XZS7pUfw26xVPb852N3s2UQhxHvS
lXg4MNiB+nr0JgvyGzRsueY1I7EpvcQlDi9XKTRdNzG4eWcZpWQFgE1Phb6r
MZupAEWtNABJMoVT3PkOvrA07AggHXVv3MfkCpKZ13AW3O1BidU4806aEB4W
vPvfNWVqK2lkCXeqMqulnDlG+CiY0u8dZABGh9fn4Yncx1pV93LH2PZ4T5an
Ol7cVgvhoVkGqPmE4shj2jZDZy+8i/KwluyR/e4hcz1VBF/EOPc9S1aGlAhG
gdvGfeTNY+aIStlw7J/K6Z89gYLHuafks6LKXqRQV2NI5EayYK5zpLy3Jpoj
5IUR/bxoZ2P2qalTGBSyHfpwT2ZOgDhpk/OpKrZNe9uLUvgK8LjRdcsb+qCO
ZpHYBc2YS+D0h4kvo8CTAfxUhHAB8zyt4MIZ3gUDOcYZzdm3vlPPjbRWAqYx
/TnwWOUL2pE2ZA0am4kM80nmWZAQIxyt6Ihe1XVWYS6I3nRHbd7EsCJPq0Es
4Q4V3WixGbH0+IcFLpvknEyW9hJ9CzcN+CWyO6aKCPU5xVmgnEHRMhl17WD4
D4nYwrNPDEV5I8rCgPx/BLPPKYJgQHZKXUXZuuLk/7eATh5LP4n1f7hv0E3w
ZMX6OZ29IUv0g/rXuiLOphD5ZA37f0IR23T/HrlvqFOr9CsFeZHJGpEt6Nso
XJo5mSY6PGv2B2FIS0B0jUHnzmIWacf3UPjKczrBrnuhn69GwrP3DUTCy9qC
99QT72d0PpMu3HgxuxKqNsaEx/XYQqP/0s3gt/c3xvRqa5BC4k/aGDyMI4as
HBJwcHyNgZV9zsM1wkRoG8QIM5ZR4YSGRHd41xNKJJBu7eTiHZVDEBuB9kFR
e2lf1ml/Gv4Y+YphOSR8/+/pVL0RCzAbDbJ4tmi6tjTOCulKw3AldxOHctx5
IuOCIszVlhGgLlwDRIoYjnl0dZdgegW20XkpaJrxlSSlFpWHga8BnARnqny8
B0RfTZhPso5UhUJeneD/4cvYG+9KiRQh9zMl1Dt7Fg6JBJMgD8z5fEjh/ZMa
Metl9/ZJgnyC3fbZThAZSMCQM8AqM5t3r8uxFSBprOBjwXfBh0dHyV6wazUm
BkseLL8MGxUsU0T2kG7E9ZGNZB/TQjF2xZBr24n/iDrAmtMnmozumBf1PbQv
W2aYggOXVSXNJkVLGU/xF6WksKP84zHVvSz+Bgg2OWQcxAZ1aTQOpHm+EisL
oXVGcf+mkq0KWPYr16nZyvRhLDJwWUZBqY7DFrUxBL9F5JGY23+VZLafAtfW
l6luHaSuYBnbk4mwg67fLYmPrhHzgUpufaVjmnn+W3uF2z7HTeQx70yW9uko
g05j+1u9W2dSl27j3WxCIaFxeNLhgUTcdcpSaVj497nl5GPT537KplsKsq0J
dqaa5MA88vg+8zvi/PKjTF0zRh+qm+QY8QrRxRPOqqyoIGppw7aG0InCqQ3e
G05YdKn5tYrsUlaNHF96oyXOYsYTDIPSRoXhdWOSlsHLROScVMO2EbutCDO5
Nrl+zzrvopCuW3CxRGeR545pFqv6O84qamsxO1iPsVHtAzJGzrSlzv5XLwEN
YHjvlOxGN7lvOgas0lxhh58dXdYa1UsMLDKcJDUd7Z1fVTnW5jI6s6q/q3z9
LbVoNKnvzCheS1zr+YVcEvvFltYbGBam5I/fKxpL1TxDkdJhRA22gEbc+TCn
tNHbNvJcgBIz3XX2l7vJsLIW+r2Ij4UPG0oz9Apk+aWS+ubMOkwpx0+eCr02
Z4QbvhpTydnyPhQht073soaj5P81WW9zYCN/e5Irn8NZk99fbbuTR1dqBdkZ
VRqGbbWyU92wVaDgBATQ8Hct3TzbfuZH0RE3ET/I4IBE67f7Hw3+1Yu+WQ0R
7WKNsESU9w662Hw1HKHzEPA2ZZBVtJziUCDUYueqabkS0xrryTfpgeYSbUu4
mXCDTlSjzf6OXPh+Fqmdk44YLS/Qns05Gh82shXNjjJj7hSOeltch2/jy7Py
Tq7CHRJS1SrV9McAandx2PmfmW20CEXZPgLE0wPrIxoHW6AvFM+sviw2p32r
S/Bh3GymUW4G8dP/dmo4hc2emFWKnB/JmEnMV5O4L6r0jKDSCi2AUYQdAtSO
kwbIf3o38pm7TaJ4+y0nNF0BR+wnJGTr+mHxLnRPLgU0nHFoGH4VBH1lkIKP
pImfPR3KCbryXaR4+/uhQqv4GJYmNl9NNqEcoDLyionylIIcGjOf1knJPd9h
oluKp4ClRHeW+bAnJbZL4jdsvK8ngQoBjmTTU9fmY1XoCvXLrgAeZjPUmY2D
GYKfObG/yHL3czvfT7o0dLarf3yHkAdpUc2zYsFtuwAd9iRySq6VsFkkzn0B
KI8UwoRHYOvGm043NYRMi0sJxkl9ZcWSLz4NsRxKY/9njYWc0pvitq4oTgqE
8SKNFmSf6Q167wdzYza3G5jn9F3meh0yR9Vyd2Rs+8l8tvfWgrnDQd66J4B3
5VwA1AEdDqAZoJuR43lziUkFwB8YEILr5wbAmbGuW4k4n+1d3M3JOoXnd3eg
gh0DbVj8eCNKnmG+UizVaENZQbHY8XTktMdif6bNO0ORZG5P1MC18dQ1EK9t
p37CSdYeOiF4Fxwr6HvabYr3gAaSB54RpCYDcoJw5d6mWxHqcxzNsFnY6eYW
MpHPBIx47GrtCQnz3PJkmL/YBFwkJlwydoA+rN8l+cNtKMk58QZxt6JQVRO9
pSqZr5xGBWjvX03/H58dOBM9qf3Ei55D8KgC0Eo/Bsul3CnspIAHXPVSz0m2
adx5ZoyTSZiCm9qJN5owr2UTSh7qxzANv90lsRVzxus7BSql88Csav/+brrr
TFM7RCsOhp26EfhDB4Xmt/T28tac5BY34TGMP7h1uzQIZ6TjuQnF+e0XuWFN
4ys5IXOcKsx+93YNjEFtZz9dZr/uyAN2Ygui+F/agZV9VP/CTt31cnhv4iiS
5BJLVEFLwdBUTHS2UMqXZeC7QpPotofX1ADBWRlswv8mLgSN0Uo2rTQaR69F
AKpy4fxC77sMynjTrS7dRmlvdewXSluzblz64LwIwe7JP1PfuaMrbpH49OTx
vd82YtcLCGnib0xzEr277LK8GcRPbzraoNlWiOafkWqc+9trnEpqLmAAecTS
qtB4o4+fg4ymE891YxXcAnHParc99vkDhfeQEzO2Gv1tIUwI9EWtOtUTf702
xhJRRgmJkQDvNczOtednXKBv2nmYUPEf6VcoUwbCA5drI1vQGhKsgErY4imH
h8+BC+um8RuZFwZG0yDADu1VHN7bZjSRsh8FpWyLm9r0rOHB+v7Oux5kZ5sS
fz5//6Z7gHdWGwlUbWYEqG6RGzwgNmOyeW9mH0e0BIQgwMyRDGCiY8uwrVS5
mFI8P0tYUW467dVW3LCWVElYuMb7hhGaeWhhaGXziAOud9ZmnJK8TIeeiOS8
t1MzSRxqMkGXIxyTEVt3bDx+AGW6+G3l9raybGrd3HCMtyBEpwH6/T85nv5L
0cjtLsFFAdK8FSWOKGwgcQpYvWvQbZJo1qHvPl7hSCe4j3rgrqnqa2oXRDVv
/bdRAIT9R/x1YzuoxmAB3A1QznhNlX7GOUJO8p/+cCpKSNHmECSY/fSPc/G4
DkfV1LCne4XrRhEXOUEN+CR0XbNwEve7jCM/syyvSq0kZhkWS4ybIqQrdL+F
ZuU7OPsuKpto4tMDmLqU2pGkJN596DabBMfIKim3ckM+FBySWD12yRfy2rGa
6QveS3csdDXWZcPAtBAIG4nwR+Wq1vHfE+Fj/7zLHCf09y3j5adxyxPAn8Yh
XFYp8ZT02NPf8alqqXVtkL7WQ39uqZFcx7M4+9LYrOPvPyOOV6BjdkPc1K5L
dp0ev2ft/KwHKwCbVODZD+Rj8mw+J3dCD85si/HGYLrf0rBwqtUvwoOxFwUy
vEXQACVAXxdGiwAhDvfxL7OlZ+yWs96XHRSeoooZke7Rq5HUSNoOYbA4ExvZ
VazKYT1H5jslK9NVqzbtaiMvlw2VKe7QEPvUHJhuQ8puYNrZ14hyaPLt2l68
8Dk5L1JnxrU5vFCh8e5r61x8yqCwya5jmmtRzhgd2CUnYtK278GNfWjBmY/w
nez+oXmtWVUb5w+0ngrz21XCGENkEOmWIGRZM9kNS806m9+FwajRVwU5EXh8
brkC1kBqFK84KTQtp+OGXVMBtAa/aAyhmAJV2Dwh1MlCx4krjp/C7wZ+jcFh
YKFGEF3Aj4c3ZiGQ1dUUHW/Po63mFQiGNiLXH4u3zYin3ManyHtoeXf1lc1Y
7oxxA9b6HRzxaM7KIUw78NH+jCXBd3ZIA0a0FheOEHXpCYZXuPtDxxqvhWqa
5mdOdEOuj0O/86CjYjqdUBJED+hM3Zf8PH9G9t0IjP5GxxvhwBw1GTUuMd4Y
0L9DwLVObXGIraHdVO1f3asIrpvDC7Nc5wkarzYO2hJcISh/+hZczN5gdkvw
31lHAgXVs1UEyWjXZ63ni8h1k8ybRO98X+fd/j4+utKg9vM1VEcLTKtUtiKK
87UF8vnaoSjMXomLjC7HoZaouYVVAZKbN4UdF6R/Mw75kLBTs78WUXwtDmr8
3YoMk0NdvA+fXs6pisQXfcNqUKe/puDuVe5ZGw6uY/7ZthUfvyootShPb3yb
deYUth8QiodfWWR3EaAj+dsJt/1GXoLI2LBLD1JN6ayYCDaZBD7HUqepuvy1
3gPSNnafWuPoJNrYuqY+RDFy+w0Bi+OWKyzcjtvBU8slT35hG0W4alUvP+en
6h4M/AjxiZemwuc9pNp8jp/mcmf3aWrf/R1IHFDrAZvcJHckuWjuUp07r1Ob
QM9kGfzkwOkb+skaeVZ1q5zy2Au98BfruUJ+tldzU72xS9yqo3+XHoPfWGqc
WzNJxcQURpT8/f3LJqInDcPV7glzN/FWiWP5o/dTW8YzF4nFiPlouCTjoD9c
qHKLsddkVqjuWpSCTxDyYAivsfd8PJ/N9bZ6aI7UOFYNGI1RwcjxzPT0xQH8
+Zg1aF1JBZ/Rn9R8QvDb2+t5CLiEHq5jh9jIsEQwFhyV5cPTb4S48yA4nSvS
nnKz9ZSqNHlOs6gR7fb3G3gkXlj4A/3mLM6YzPpXpKTSWvk336SLBtrsgGI2
iQXEmziKdQgqVymO5sVIDbQzLKZDHkGLutlcvd/2RvjMqV41bJfeCb5+F9sE
K3RMfZktFGHzxCnjiG5Wk0wWRmmWuZakB4asu2tcxYX4ISGXkPeQLFxv9VE6
0MjSkdSoeexkX9z8GfqAuC8dt0QG7x3MLAjFYCM27j8r6ElvQSGWkE7KQPIr
j01m9mzLZ2BnlzhqSlHMCPYzkc5CPpPnpL//I2NpbszWpsPDm6+iko3bN2N/
DTUrPVDw6EoIj5sg3QT/iHfekmr32WqPOTYNsekM+0aqUn4EeBDvkxDZtunf
nOPYXjs21JCA6hXPVj1FJQdpReXqZKU0DiqOUDi44jWmi8wFZ5iAr+EVppaF
vhQYAhkrVoZ/5v6Am9elQ1imy+LymIxs/Ch8DdqtouMt3M9NAYXaHmCBYvJI
5oCc8BGmsYe9MoeTXsLdCkorDXIzOlVmrI3Noo63ZEuOgK/Dbaif9Ik/CwWY
/aZoBPYIcH2kO/m4P9Dz5WhYLEsyE2EhRkKbo6DY9n3JhwarDg0ggfhI0fD4
/5rmW1GAX/CJH+Lf8BogaHOd3QMQUcyv29x23/8M9PQFLkllk3MuvFw6u+hN
gFWMUk876L/07moCb68Uv2PmaxvPJrDJPFzh/XipxbDAndGr9bsKxT59UXAm
dVYW3KWejgGk+gruAR6/khNG3hS5HULDWZG0XyDyZ2HfpPOT3zqbR7wkYmyg
Q36GiNeBg98FLZssVe/AXrxBs5ZKoUHuNIAdT8MnaVdb0TMpgXmsAA3aa2jT
G85VD6kjq4VmyQx0g7O7H+NZ/6aoy0NidlxYDfOjXix8WkVURPoL19VFucMe
0x3Vcgh8eNqo+X9tT9U9QwCnoY49TeNCYGLm2xzFx/L1ph8k8mYtsRDRXKKD
9up58KUtsNxKji/aqJ5nSPBE/cTYLrGcgqqv9mywA64lDy2PbtOBSH4k8Adg
tL9lGbDVNxa1WT46bxVeS3ed4L3dvnytqZ1OrXEvgAOqibCWzy/B95DTRNqy
/0OMsA21WeN6UsmsuoslyUHxlhMzoGD2hBkAa2OJZhtSY9g2H6jLkwc7v+JM
iMGj76TMA7PbpbGDrkJ1pqgxx9qJYOvdI5WQEETcCXT/vyN5+dDJaxB1zr1B
YQuIgPTv1kue0YGrmrMYfXWkZZFz6Vx32IJbXARSt/Jn6U7r37HUulD7bU1D
i5JaqnvqYSUifHDrXXLh159tP9ElzrMZhXUfYhJ5TyYoryWuiUHPJ4ZoMF9i
B6gkPVhmLdrNmON8myXC7QwAhX94k7TI3VAkEkarAJFabUZofypzd6eb/n66
gMRBYRAouZJZ/OzctIL9z33HJ4yEPmzvZr25FADXIogQoSueuaRaX1Hw9Iok
rgFSIaBSOyJuCyuNrcC6zktmblkNcZhljaOr1QuAXreD0h1NcLzLhNNZ7sDA
FaI7QDx+S5SlafvoCefDZ49xa42SugfmA0yef+Liqnm6V4KUc6C1mYFeTfHj
ovT2HXjxPaKiJX0eOPwmrqTA8ove9lEpjnSs/srEGWJ4J9bZnTIeoGNReOH1
Gxln5IuPDucJBg/NC8vTdB+OVV0p05fMkn1JKXrEzN7xo1H2aKb2zpa1pIco
jAU/Qc8xdIJPR4XC+9UV95z9C3ImO5HtsLeb/DInCJzofYaXWxXNgU2BtNcH
KBeU/2mjuRxvLyl44B0BQDWPUqep9PyRteADTAKccqcgXucm3ui3KIGXtl9l
FLDd+KLXgpVv9H/4JgFNksx8tzIgo7YvPlrARc+4dFx+mIg9/juIbKRlZYa8
eY6yRa6HAxHB4FdScC+iS4R60EurOZsag+2Xa+6cTczwbHcCeOlQlpPgTxEA
pOT2bWTIjqJyTQjUVieoy96WnrzAqrpU/fp1evExb2zaa0OeGv961dr6Pl4k
/r0mbZe/+Yz3qjWNuKacx4p3j5LY30RIBxxTiLqbrPFVCwWqF7CqcwnxjO6A
i4ORHgaqK5CH9uJENRl2VCQndpKozyPq9tw1uIvqHHVybsAfc9zmH0Bn56dy
+iSX68o9gZn90dpOY3kimoIBe949c+M9ffvYd+oRKw/bS8ReojLIRIfd9VRw
I39uiRobqEYdzknXA3PIyxYxpgdqKkZC2SczPjZ4LS2NAhOv2Ghql3jmKAOE
H55P1E4z3cSf2Denjc2ZAjz+/qBkLZgPyfPcSDtx/47cpzm2zKfIjx+IadWl
FyhJxmkqDMEKeXh9m2ORImExtsvPKeG068VS62FFtbPXLiyLLKtb39DvCnXr
MHF+h6yUkiLPLg7VDjAqoaK363+A68PHQjEeLb8WxcBWd/Whi2S9eu8NFQ8b
wUYb+lEZfKaMaMENEgbvtGrOVv3hw3r7Ej/fQdguEyda7FDoqWtcKJwByC3T
Ffdis7p2tcMytKYNCD01a/DNY+T27Huq50K3VGLnU8MeVgjiYwvNUpIlzQEZ
P36ZYXhQPpfLnQ8/nYvNkPFlWTBjP0B8d8ggpb1lVoLNCOLTht7tcbj69dLk
n77a2VZCSKT4TiPMOQAvS7hbclaLhzXvot4YzhvoFl3UYXpo1gJEJlpYn9aq
XHYst/JzVKZwBl/cbnlP5brwjSqHt8R8V99BmbdftsHNdQUugL44a77Xrxfh
g2XjxuFZZoiO3mNMe6fmraAFB/dzFUDV241RoyWBe0A7ysDfcKYow6cITz25
hnfQBVAeA8T1DbvEpMgTIPxr9GP25vb2aNubDHlZe5Zk69o6rQKa8fB8Lvj2
baKAv/5bCLzMm5zEf5K9MeIRBDD+YzfVStA/RXXe+YbwR9R/LJ1ajCO50fkL
IvTm8ZvhozSHjsx3Ez4cKDuNg1qhRUXWKxxAwJC4RwikPpeAon9iXatOGeUJ
mB3Weegp0P+93OVKp1KFVAObnW2C80yLpPsxIfDa6pscmeAi/4Er5jUfPVWL
EMuJFDsBzZ2ArfQMqpoRm8FBn1FrtztMVEZF1jLilO3nAmEheJelt5YE9peH
w1hCK9CDMGqPxqPufUvfh60RmmtK0hyuQBTBGzZWizuUMfXdsLLtNw59pQRY
TwZz8+Org5o2CYDXSF2Kw+8TaL1XeiebGGFfkZGOhWJtcrZsdhJ5XLqqTiuv
DpRXw8usHPhKbrJBSDmyoXELOKcOQZsJGM63tzeUCnIp5fK4L9igq+WuPmTL
Nb2lFgXfd8JM9bwvWKAqW7TSKmIHglLEUq7StgDbTp4KtODIbYfQR+YiwXWR
xhRvu6Hd8gRxMil93m+l2yo/33ZGSXENruwPLQKg76Y3iEET3/TsZ7MC4owb
6XCTkdZEBVL/oH2quEKf74qttSsqYfsiU3yG1VJR02amLf8/nMfjxTuDbpJ1
GDR3wjRheiwJwNtzrbb+CBSG3YgoUxk4tkGHz7XOa+SA5FbHi0UZKoVZaAl0
mmTd5NOyDOgwOsV26XhMmMCJRNBy4LssoMAcVYSDZgiwOxpOwhj+Pt11+KXz
YUxf2l2vYFpuSaUbWWgOTAXbKr/s/f5YANcjRGQB9ezX3W0GyyM3g1FEJ2zh
MdmOcTMyRKc6VgYjF9ggnAISNoLn5KCSSw2AzIgdVNPr17LglOLcHxtfHNLR
7SkBH1N52ARRYxVRP2fYJ3rIB6EjJnieT5uVGFH4EC/CkN/+QEqr5AtmYCm1
DVPmbE+Kxps4PnlDmfWslxKO386b9dENszOEqSUtuqPDmHsfhcizEJxv7QYT
Coz+yLYcAOuU9RLhwXHxg1AQPIDFAoDqShfWd23bVcEMSNYYH49vTp7ghNka
tn7w0TaNJDwbgb/0MaLPvQVMhiyZORGLJNTF47G3jRauZoXiYjiUw21bBj94
uIriHWyKtO8DENcG6saHLO/OyTLCdn1j0pdupHOMzm0K99cAQD+UzoZOoWvN
B5pUv7UvZqgBidUhvvGKSDl7dTWdu1F1v9/PmJsMJb5Q0RF6ZlMBHAiNmB2O
+TBlwTK8j8FicTYI5c/TOMeb+AS81nH73kWq4waA6/Qsg49w8O0OthiLdGVs
q0KWIiXFHcrKmdiVEBE0nv9kzyRu/q0EnmmfkIxYjdYw6wMxG0MjHvTgdfEl
Nc8dbe0hcjxQ68iS/tIVQd/Wz2YmIgSULZYX9Y0mbaFife+soc1tTASk4TeY
pnJtMiLjDNJtewvyMYa5nebyCpqmBr87wophi1knCEatk5enQGmrZ2wXz2oA
JqCv7n4n9f9yklWT5QYORo6EobApmh8d6tpGvFUNahVAWbNGSsskLEmf5uaV
m+eq4pe+90mvh2xdOuXch3EVnufhkDkYn7e5tQlWvDiYnzAaTacc57vo356D
7gxRyC0O3+NDQWGplMWakLrA/yGuPfhNCH5MR4Re7m/KWksY3XC4ONsu/cKZ
6Tma7xQW/T6Kj9liCdtHfFatVSt1wI3brC1wBVZbz3SOZ0izlwargPwUWS0H
7zaBr+ZqeVHrk5LRLQVq0YgBFDx7/U0J+7fGHnDk9fVJVGmYeJLlD/wl4B0u
mwbI6kJrVvIgZuSIXMmmvU0SMStisof1OGkkkF+MusoLcqYmbITYJ27MSpxt
TZZ+napFh8ro6THQJ8S55ngy/xEqGnaBl0lrj0Hn2MdTdZKvPSpH/RCs1Ku+
xRMB3TDMb2GWtB/GEJDVitEF07FT49tzVESVwKDEdq+PR1j5A2WZF/ogCw7/
/6ybweJ87C8uDALjn9+yWoOlxKgP2hSoy1tA9EiXtQNwGVLCYFHtii4Fax+o
zeCrxo2dFriEzADU3SUgqc8qEQXX1oK1jpKFNyDZiEd9YJGjGFYSN89jmXWz
5QCf9r1oCOnQGIA00IU8qPOBNeRQN3zUHCjgDbJw8/CIJjOww9ZDnNh3WZxK
2pb4cBLAJ6wltgzyW06Cx1Une+aOw1VEfAiTNWpa9+pb6sCGw3EJYirRGKTj
Wja/4dic9wqauOPy27DEqVri1Rv1uaLvOymRaJlQDlrAskCMqoKvCmNL61Eg
FiYyp1dBAnPCoA7N+sIBKkN9g3Ayp0Uhs1+f0PDBrXn+CJNm3qA9wSRG/xFu
JRX2bklDREL7JB6+xiHTC16nNXNOSRTLwJbfTnqa090lNHx1QI745kVghB7U
4QwRrplv11wqCk9Gs0cS+BJMJzoTBnct5RA1PS3NTu7YdzbxtC3EehOP+QR+
JtvgsPEUpsOpSSZGgS/Ca8dFG4yxaCBHfGyq2NgkomR/+g845wRA+ieHiTy7
bly8wru0f3VlnBTJrVvYnljMYBCnKAeZHRYRwKDhS4AAoLSzhUmeR405JHwm
xPFXg9Dlcn9fmFWlmEMCQYhphpB0AJkl1RidtD1gwY0jr+6zSLxlMsA4VxKx
saYZUeRamABdA/n34mirLa0MKEAAHxAC1CKq7rHOF+LbUR5GxosFRUKM98iW
Jg9f+uvCvzFnRZuh3n/QACQXZvCY6ldwWGWdbKirFhpwGdaUi7VWnAA1c6dK
Bvio9NGHm8gpsOlO72+hQUMT6UNX+1GKpmD9WKihZ/qZLAPn7cnm2PYdbHaW
uBd18mHqBSI71prEAgEynHKOvvneVryge2L5ORkB0oWqsjQRKybD0zileXOE
E44YxbU9dns6r/UaIcxGSKGfLRUuWQqE5wo7abgwuOL6OD64E2Ul13lE/Kt+
SHaqpWSEUSMYSK+GrwTxU2LKpqaLSUcbdojPrR7zyUa/wPG9eh9YzA16kExA
qyJy0BtS3nhQYuDc+ZcNSPILkiyW5lAMPNlSUyOjsbIC3QLR8oSVvGM7YlLn
SyCvsqi1rC36/YsCNlfDF6OUOivOnEVWy8xNbl7qvNJ2G4XGh4mhhLnqy92l
zsRz3i8xHjJFLqG+Ua9U4c3HsHL8vz24HGfEoQCzUG+JM+Vb9z2nlC7E3GDo
M3bz0HM8/an+NaKIAfGobhQm2HTwNHaz40yd8+wcW82TxDh2pu32s4uWh82+
ar1H4sjU9TATMVKRpQImX9G2gN41SLaGgGqRswvcMrAyJN+4JaDR47Ul7gjs
nz3kThsA0/9y5NCpJQkem5niEsJtZUMg2raJ9Ko5MVOtlPXSBoi/VAVJtbEy
5cgzEsSoUUTVADJ2MjownhYmHL2RgUfJL+dFY1Fpumxi5XS5IGgAhYXpvA/8
XCPhr3CKoBmelxDdWl/BJBlYIeJ5QYy3Kjd0X/N57xC/G7yV/JKy0RZ/fkH0
IX3OafHw31ASohqmMqtMTRseq7vaNHNZVpsD4DC8/Tx1N6WX2kNvZpit15EK
EP3Yo3V0OkxhNz5oOSDRLNauyHviTE8agDl8n/dGH4i+99nMIswOszMQC3fO
DKOJB4VKPp8CNXicW0NL/WKuWqzoiV+qDQs71uFqh+M9ALUG2fkZoKHUw+d6
5LNaygV8m1fNK2zceBTDD/raCNniXz4L0Am5lVqmgRh6UWqnfAdi/OEMO/kE
Y+71hlypV+MbK2U/hEbn3UChziZlG+tH5JDJrdx7F2rFxBvVHS56B9t/jyf1
hlVbFsnUjxAlkOY2OsPo2aDe4pYfn+rACxT6snFh3OhHLWMZgHtUIq84JIvs
cESb+ZXzMvV5CZcgBVibIe24k29x3A97ueIP1x0kuInsWrM+UZtbUVGsCiLy
39gja9J/zjGEE6k7im/2hwE8qzjxTEG5aUPD8ftTo+1Mit0NCYwrwMQp4o4h
eWu1bYl+PwqNB0w7VZQ+7Ou/7D9frX9Nrkj0svjPfOmVx0QZZ7EO4s4poDce
OBrkVQ9XWUCdKMbEojQR++gfSlvgcJrLCpXIbALpVfvVDbGGLZPwej1nx4OB
7QZe7QeHdnpmXy+2nkQQ5ok8k2az9mu0ygzaY0Qut6S3L+PJuzo9vQeEv/on
KGlQRB3uujnMZtFYS663inbI9iGVriuVhDZFd+FqO2NrZispOuxdrtmS0LX4
5/6uW9xZVb6MgvhC6FxB8bFO7DBLwLKvqdeIrre7FldYixrTOBi4879xfZnV
6w4M7SnfCCCzoE5tXESZB1csI9tVGOpEVzOCgF3mtDI1pfE3PVZUhjQCS9bY
1D0Se3LLIsk+xK0oLvtbzK7jZLayw1ZLmCt2/1Jk/XfUZACqHqxuW3PE5GLe
Ms4pCXvZhkrlJ4q/3JVaEtg7q388XWwKBhSu/9K5XZZtlApyCA4EzYv+kSFQ
+p4+xqtXVazT2CDivPeyFkEGM31+Zg2vV+4CvBl9wroSSSi2RadMMujT/L/0
eHXUYLTEA1IeAYpDCet4SPKTAabt1rD5CAH2Sf3T2PXxw1wTQAIdMh18dF9/
xIaxm6pYzcAisR8ry77/A+2aFpqyZjyXUF/ciG/xEwYXg8/3kTHwMMawEtVp
LkYEOWsAY7ftbzzXYkN3anDc4T1Q17+uoJtunhO2MmASHct6NO1pdlm/Hwfl
nsKWalIAgruRoeq7Rm1TkR4bYrZthAtaY24TBQ2Hscc13WlC7AO3OfWLGWp5
Iz/V0zUBxiXLdNHOqllDIpKGdnkdDAVWgCkTRNLbKnLp9QBU7oY2g3uWDRPm
57Xf+4ZCGOs86DPlKQ+KNciwVCvEjD2Pw+3X2ACKHOWo4OYPSmzKG1WvRWN2
Wdqfhx+VA0KZnBMipGHuPP2LugOzEjnHYVGSgORJyoHPtfpyFuC1zxmPDiFw
bNb5973ny+1CQpQLTIufDtTJHdGIS7iyr9a/4W103lKyq1qotC3Az6lND+Qu
opSKtVCLGBnxgo+40ZhnXApgZEFlBCKu3sgE6Q6K9VpuYGY5lzgij/50f7Ij
3hYGlQENndAbC/1HqIIJqs9EksVfWHAeLbFNR15WiGBAuTSU9CjE0774qiBd
HicqlhkOxtvRP3qPrwut7EY2snqllpPpc9fPaJ9SMoDH6/fLpyQSODgEQdI3
4AfXlC5BkvWa1mrLf7xVvF3NZn87Fdu4Isb6Dkea7hM0CcxwCPPDs0hUJLW0
D+e6tTuAZtuhkJqbb1A4eCus/fH0HoBcKPlij0W5ePyxAwyszjhMUXgT4R9t
/Z+QLMj6n/Pn4A8m+VL5earGtq1msAv2R6NHMNnwBeDK8LQ70MSX4uhzTBV9
acNLRK8QxkasgsrkRfIGtP+4qozQ5lrogwuLU5lYNU+9d6aUHzfALrLxWHGR
ZDRwhfAiHw3IFl4jVFaCxQtDxJPAza+3lUOPR2PfeGyXM21sOZo4e96QdgKq
07VaE3/uGeilYxEtwNSxobFVLD2GjGaixUHONgIZKDN3LQ7R0W+4wJ3r4dSh
g/xyjLpxYoCxaNcVGHDG4MfQHIFSOTila4cACaJfJ+hwEfdyIkpZjOGA9fg0
a4UE0D6/MfaPfsaEAUTYmvP8H8M+H/LSZCK1hAqqoIT3wBqbEH82WcOMJwjY
hMxPgjIQdrT54WFQ+WDonAGEwd+u2XI4DUTQtuxsZry7cdEjtLQcaSmKSz9n
V6hn0iVBYpLv07JaK+1Jgm2MOpkYdjPGd4XF0+aBPQuPYIn2GTSwHN8/nNh9
NuWkn9EdRcXg9efQvkU/hfgR8QIlCCw2oJBFGp6wkn1+ZICJ9E1z0s0oyQ6E
ikRaKWhoXe//01ceL9ccVD1KuooIr6w/30HKVQFSFY/miiG2u/ch+k3cWit9
QGflTbvGS3amuCkfJrCKa7Ocw8v5AgUdMXzJQDTuMkv1CR9yaBTehKpjh71f
+nDLJuSp8V4ZbVvK6BErUsJ6wiHTTUF45UVfm3nORNWj4FLhFejbHOjbU7X8
LEHS9MXuHUUwL+r0c2EUJVnPDMNNOTRmUTnfGnJ7+GbM6RywNYtrAvBtrV+/
+w8oSyN2HANTpfs0gQRYk+eQZZaDNCKPtWYAmykYeMzTpeFslvxj4d1D38Gx
paunwDyjadOVpk3aF6RV+9xe+3PxU6sTw0kgdIZauzJzUQUPZ/VWtRUGYE7B
gD3WEY4bR6GTRv3LOKQ6dobvoFmGXr7T09Tz2fGMDuOMwlfi5njPxejGv4Eb
Huq2+wUqVFR9/z/ZriP9rrpr/r1YLu4rpZP1SYD+pJgZcTRpGkeREr2wcIBE
/p9f0UQs6U4A872iJ8cyxqcrylGe2tbyQ4vFU6styLHgYkQPVVY+Nk0awd2u
4wf9fZ2etEm0H2UxN8vxcLsDTqMD2OhxwWlQtcIKRagjPH3k9oB9rSpf6st6
CrCipvgac0Hv6qx13rs8yzUltD1YvsbvE/yZmskrLCP7eu6y9VbhGo8K07n7
aRd1+WCxLg1MGZ21Z0GvyWwXK7WAQmIHVbYnErsB2ugSXrziE0ABLpNxk+p7
54JBHt0prPSO4lSdYGRc/iiO62b/poPbeSqktHOpH5qmzqLMlhw4nv95RSCY
2qT3PPiI3h8sCtRJWtDz+0ON7jF2KcMG86HFbHQRVFbY5jF1Lz2TxrQGlUS5
e/8UDjbyKL6pLKd2ebtmnCjw3ZWxDJFjAb6LJTw7HkAF3vAzb3dzVVzZH0f0
c4T3Yu5Kq+Jy/qw2Ruvpor8CETv0O39tFvVICe9j/pOln5Az+3qPosdncvq4
9avKlq37IZHy6z80wl2dDk/muQHBnq5crfiWN1DGxAE8GTq1VQwtFQh35tam
S0SVZhbK8pluzWWqZC7PoTzhuH/IQc5dK4x6Eh0OkDeAuwJ5TBpExgIO3ulN
04KVZ+RKreOhsaUxdSN/ywGUlJDBT8dbxhWe52/HAUMGpyWBRrY9NJUAY1xr
6ShE7FJqH7gX0C/BZKM83Cz1QwsxRR0FRvjrEJK8WXT5mLnWB10zGOOllbqO
6OHIz501Rp1vr4SLEwC06vih9+Z3x3eMNtGvOSlKdeoIJ5FxYzqOMIZFRpSD
wu6L3Q1V+5LOwfymxTXWQy0UF2usNsychvHNxr2pLFBINnqQ+Ezzv8HOpX6e
3cllAi2esw4GfhK+2Xw0OHlf0sJG9BZcYym3/f7ozYODIQTrtyhlvpGcHUj/
I2ZCIHP0fS9W2nNhcIrFSrCO3Wq4rhJq1Y/X0VxBPqBa5AweZoocHEnCbveQ
juVnCHh+Fx0wBaDtDl0J0cbF1/58wkMHHEaY+Cls/L3kSJSrrf5uosUWy/4Q
6mz0fwT0b1BmG2/UUA7nk+8Pg9RrmiHVXQfBzb5P30/AkzePy6s39Ug4N5ad
hIF+zuP6hJLJ4G3iJ8fM3b17l3NUXHQ0cfVlY/oA6CakiUuRim/PZsXI0rPQ
npf9WhDUNH/J9eHjnhJGdCOOvC+Vraanwuv9L9D9jCwQd5ubts2JHtTaqKaf
goQ1mkaxCdVuEp1x3/Qxndqzwlr0LxdF9/yISo1BBXv0yUi3TXbZt9U67VaY
03K6+CZw+h/P6ST+2iHaLyv+iFpe+1Yy2me9pbiMrixmUoMPkUa2tLz3kIaX
VV2A3c6ari1jWxZUjjQCyRaM3vEoGVREHRewoCpwnWccUdUotr5Ft7Yi4n2n
CbY0KJ2f4GFGq+WZBVhFGdXALEA9QaTmA28GugxFEmDNmxhCYPka2rQXPMEK
AQfLUU5ODP1xaGthm0d7tby1ybVaErGxpqVpXoueowFDGyQw0jcJmm9AjgIk
tasJy1MG3NeF97U5xQtCQh2G/iw+QVDIt9wLh8OJaN7/Fh57winXN6Jomxw5
IO7eERhOlQ8mZDSkhbldUwcH4Rsd8iZj8Nl9IJO2WswKkRRwJ0uUitobH2ns
ULqD8+dEfEfzFzNONpt0F7XGWXl1sRTUS/mb0Ax1wiLLX+1BCGnblxXykpJE
MS5vpKEWaOOn9lflgN786Vt5QeMyUtJAO36e+MtiCqEuE1FEPF2lSlMPHsJP
Wh/x87uSTICh3u5BEkLysfDDAVkDzrml9qgnC7ulXC2EXebkmRrIvIsEer1o
YeUp3LeTYTJBUUCERX+oxJ+VsGuPYljykMEUxYGuR0sax8ztxIgJ1uR9Xu/e
rei2achkzeOLPn4FzwajNUf3uT2UWekNY9QGYasR7R8lnbpbasXJ8d4plSXA
toYLLnbVhUejSRdgIYcIb6CMJKXtT60ONtR5cxMZEydKSBKVQE/29IBWbPBi
CvRE5uxSilW5ihnft7eGiyojcMwAlf3JezkluIOVn6bSfkCrSb6ohZFPIu+T
kAorJcYgSsd7f/mhUUy7EIZeLaICvXnavboB2g+mn9YHFEFYZEwhiUSHTxWI
SqnKgLVgFBAVjs2vdeohlU7CiCdTUhdiTH9105UzvRfXmirKTbwQlF03HwEs
uwXNuftBeFf2Z0wegj2Hgb4zpr/AcgsUozLdhyIqtiyhwUOW/wKvjoqvXz1f
eFpjwM43+Smra2cRsVGy/h9vQeEDv8+g7+MEEyGi/YMpLXQ/RasC9XFOTSk1
3DSOk7OgKlVu1nMy56lIzaWOeLxfur+mGsot/fatEynNq6H4pZDRRgWKKKC4
245Im8IefQ5VwrwriXVeX1ZVSMZGWCsjhfrgR43NmanO5Hm3YkQlbmXpC0el
UpxOBZEvm+KI9Y1QJdXjQp4OXtgpLQ//f59xfV1WK8QBr8SpsTxlGAIyOcr0
4fCrboE71Aj6yNizanZD3vfv6rTBbidvwQI6dkmCfT3qdPs2qHjTzXBM3v89
7zBj5djR2SQpOxpHY3y06cjNtEIkhe4CK623bPD+8KiLJhl+Uf2INMxvkGWI
PmpE65VDT1SwD/bXOX4Rwuc5IvnqjTH1S8lvmx2TdTrGfMIhFN6OQStJUUce
/gtTKNN+wETH+Ic2XKfhq9H34d9Ru1x1c6dchHXQuMzrqFnLU+3wER+Xz1dr
Q5c/Rpc5k8WhPyrEves/wCFa3R6sFRUh+Rr8rPqMSbNUK6QmYIMOjkTVW/jk
FSYgTc+Tknal6mITAwYdVoeShkL6s/m15xG9OMi1rKr12bSsDQJH2r2EmgUM
0nLmxMohYDddDuuSmuugmQddHBLuTmLBlRvCIELwIey/H4OW+uSzxq465j6s
8OuN9En6+7iTBb3rF1WhEQzFL01M58Q46Y1LPd6TGANLZBEYFMXQFHzbxT9z
jnLW1YgHsDemogeOoLAWPRXDtVxUou0v9nwEDWIf+Sn9Btj3ArfEHGtReMz8
lF+SPU4T54gPPDw6LjvryZTuTEhFz/gAEYIdopurOV9ElnFPL0uOxbWzuCuK
N0exFzst8jKFdyuQK4VyOK2F2yPpe7OyU8lGy4B9PVttnOXbwL24YbZCH7b5
xaxA8ISbDnlEhEaJ+prZWpi8EHMJUpQhbJEdH+75OobI97fi/bpCWFgSJeID
EYeb4InzTFZfTF46W3uXjsG7SeF93JX33IxaYg+TydPFhdGrkgkyKI6CvaMa
GbbXeB849/JLxCRsruP4x2m4OWYg+1vsvCESm5Z7obeVQ5DlVGPqx7BXQVMC
zeyHF+NA1N9JduHhWM/XQlCl3OguqeG6jh2EkQaf0ECjEN1CIjNRM74QpIkf
b6c+qVoMRLSuyIxCyfS2PBZHH1mwduoSmTcdpqLmVm7lJcim+QuxM9KgmSUq
mJghubg/6GZ7L5t3q6JYMjAyH3gaqluV70vgBx/0WQFAy3FOO8UgZPyJbpqK
LmMFKcSo4UXorRk7xFPiHDA7oHor8rvNKLOPuWT+XRrJRTVuVBCa9cQ8Gg2L
JVfIN+MY+7d2i6h0yCxwDUf6dC+yb+CmzQoNKxIlJ2e/FS2ET2sgT4gINlsw
nvS2T1u0z22zCuawZ0DfrZ7AhZ/IIAI0ur1gkP0QbWKWWvLj6jmt7j/bR7a1
yuuQ0AxbM5JEnHfTYOWLNBJaO388MKNY0pM0tkd9+08QTRdsqkSgjGK7xLFH
dlpk4lLApK1vPuvLJBl8BZcKYkXS0RFM0DohNMYewVaiPIPXA/u8XNpnV4FW
xF+0ktjNl1Am+u8IAOTFQvc98IfgY9UDKUxQcW6bjAwkjklZFwYp34tRzLHJ
t3DHliQHMzb17oaco030JEMmxen9B5bifxL2eCeVp1YMY0ucg86nc/PFAOW+
To4XDHKdsieLK400qh1V4Tc5PJYJQzjLOGqsK3MX+uipVSRTAEBKGCWVH5pc
5MSS50QNFISeopDOYJFxU0PBhJxXYDcNW6VK8OHQWppihTI8bAPwIL1cANxM
XMS+ilwPZcjAAMR6nk3hD9JBU2tCXKO4XklzbjV/C3jribN4lf0pXqal5x4i
wWjPgMN8GyR6HVcEZuIIsFWZbZ1n0v8tCHR62usNCZlT1jH1uHyTOB9BtmnD
kjHB5T5GZyB66NkvobJ62hrUEeVbxHirisBvUWDCo6O5xJjVUzMN0UwfkOWY
s2KAO15daVLOGabLro1AxxOZ6VZObF5XZVx4SkXSimc2hY5FR8/XTAMNcxw4
Nt+u0YIxSokV+JWnBimcycS06AtZitEIRV4hj2YHxJmm0hfQVsf+jZigyrjF
cpvkXUd59rrx1ylVXpxBW2OLbRQyzZfc7lXkcvtCcuOtnk0mBXrdEPNf/8nb
Y8EdHb4K5lm9n96bsufYIgYVUTEc/MxP26Z9Vdv7UPUpoCtxykjygDaSZXps
aEjVi4LlVtu7gv8RKa458pP4NmWzB6WgoqPoPUxjlC2xo8oKEgk1U4Gr8zQH
Ztuc+CEKpA1CW4f8lW/TIitWcRpj5OCY8rDS/DayUssHxC4+d4UZFTYvHoD/
nvFRmWiTF+qyQpmmTR5xDsQ+t/7e33an28HFONj0Qs//57hdbLbC9lQVhVZG
pHwzKV5Wfd0MFRGiyqQJUeVnhr3SSVf7zoDQKBTdNRwpTWbExr/rSLH9slvo
ozPPdGuZZRnTN4pwL7xT7T88vCDIP6aJrNuzR7qd2YsPv/vREpw2wSTWhsIv
yzlHd0GPlA7Rzq2YfuFgMgQp5st5lQ6jiSJqTJkMJEfc3kI3Td2x+r3CNTRb
1c5SnPWh70LXsD8ywEQdaW7OO6r1eb+8LNB6VjS8QKJlPtYD+FTRxAaX/R7y
SpxOAf5UwI58T2X/NGYdl00aXBpxmjMguCmYZfi5zZ6t7O+fpQo9QJD3hNww
nfqVRSR3WVwuJ384NgAYXfQQczsmrN0ljYsH3lbqrUzHPG9YZq0o0REAUZsE
1GEpjVG5LXidmf+Zjs4M6pqG7FpQtSCSTTWDPBARJSMM4hJC9sYxoehKIlh2
ajtqlvHm4vXRW1yGDYZ10ZGOSMNITB93TElnAnhri+6EV4E4VgEvmXlxjlwp
RvY0fAxlLcyhMC722U3sOVMoLQLvY5KSBIMmRUr0kB96SuTSbiEP2rDxfDcU
OlEISMQo78gXfNRuDhw3Opnqa9KIoM0/0/u72h5pKEu9dr5biv8vAhs5Nm1D
KL8QEBC7zWvgaLpN3PSy6nABy79YEcd2D0zjHUxXwQO1kPqdCFyjbXY7b3J6
FU4hiWKC9N8brFVP6TENfOkyXYkRm09K0FViB1b5fRDiA3s8ZhSd0UJb8X54
hwOP/y0ZngcA1hPUjF6AQXVySPipZyGbuBQ9YHpBmD5saM1DsSvVh38SVImd
YQxylg4QFxSYd2BydolHei0FgAV6D+MS6pRWK8qm3gmtxrwx0WJMuG0OgmwP
BxgC0hceTjz5SM+mwpeld1WZxCBpbnFEG5ReaePZCVzy4eW0myhzrwSFgTTU
HxSzWzu8WAwYaqNljhMMplpVInWb1D9KEqxgKLp+JCRMyUGs38X1M9A9h3na
r/nd2kMRyg3NZ4dfA0Qn5k173uMNCcOYpZJjPsOqJVcK5OHQGIYmUC5p6Wma
HZky9Wg8dmNhDNrAVExL63Nh1YaDmsb/sSDM91kHGLRUWQ2KMx2ra3RgsTgD
uv1xTdmFpDYrLosoPQCPlvPGs38SZg14+l8vPGnDm7PchPJvRmPZ+5umC/MJ
LKn8f2skpfu0TN0ckgCoko7+3rjeukl1aYq/n1eyRRZOJJk4GdU282hUkWaS
WW8hutciDRw5XbBQWUREXd68Nl38z8T4Hfz7S7+zAx4s2xKkIzhEdZP2qfrL
17LRFyXk78T9/0TBkVPzazaoLLz/m++V2zTajOUP+T1NhWATd7D4axgOEsIl
jwObWa6CegbEcCjcraBTETZkg3GaS8ml6Gv4F5m0alKb1wyHJYOKxBeThnI7
MCYrF0BYGXniqYjOv/tJGMIZUk5J19GbVWFIgKZgyp1AGreQNrQ3XwD8rbDV
4qNxQl+4UM50qCLwYV6V0qqCTMTe7ypDnlG3RB8Dp3auPQfP+WV1XStVcoJz
i89eslo0nw3D8RPCpld5z054CIwQkdkCxSPVOs7FK9VMoPhRSbzHthU9VpXh
NEzOtJH96fEvgQRHQByZTenZodpYs6LK9W3n8Tx28hQsuhPaD1CM4qQkbbLU
JznrDAiWTu6CybX0wmAgV5qiyhEaWVIb0ja7r9nUMCnqQ2/aGkuQ8F/P1fXi
e5GZIm1KOymOCROgT0D6SMoruGsUmTNwG+78zo7bSPcYf319jSduc8uYNZvL
h7qvXFYd92ULNel+bdvuPEkGs7ndG6kSqtb/vPGowFT8624JXCxJ408parSK
rfhm1nojpa98FzkgDFs7wwqAfNqk1g8jtmNd/Ps/lwZQ9If5b7bkAF5VxJp5
H3QTHrKOu0b+98XcgEWrCgzy38SyKmnSAgQH6CiIprCklX5bsKcgTzRDKg2u
0VCQ7lkWTGVWF2cPYc7zOYAtNqUI2kjGMTLh378uQaa50CU1JSaM78qW7szH
ehWlLFFSKY4uQmOrYqn2W23xbrkRv361kkEVN7hYQFzt0G06YaTtpKEFuY4e
sZcGd4wcRZIdaE/qXGjhAxWgdjQrtmFFiiXCXP/fYRYy6K6tdC7VPnb6SoD/
5odMkoH+oIBJr8plKkpiUJRmj3I4awaWYqrylwHBaCpyaGx2ORjk6OIWi/l8
UnCVVf6Wt8Jmce/YFhzgzc81WpVeT7dPVFLeFaptmWFBSHjtmlWbEXK+NOAr
obw80UtoVl2qr3aAi3YAI39eB+Dd1taJALNc3FnP8kA4Nmvp27glAmLgiZns
XXb7pITJ4UFXMlOZEHrRUNb+gflIlDruv1bUe2f8bRMh6HTlgfvQqOH37a7n
odZ+e3egZXEhMfgm4/oz2Y4WTuGazxqAhBV9z1mnixxHNb1j6BwVKee73KkP
TJJwBxM+ixU5rADucLHViy8x1inbFCQd1XsCqXbw9JPdwtNQcHeii4/vEq0q
zXS1RHpBKKW16WtVKsuMG+xT+FgLGiSTOiz1zX1RpmUsnICPR/0OdNXOU98m
yFMKDVl0le2IA5g/nXaMjEu0gGisYqGeRoT6X9n4os64AK5gyuScfbWQPIA5
j8vhjveZPgRfuJTPtB0FWa8FJKbEUM6rkuTNhvz4ekGDY4taA2jo6DKQXFB5
WoaaObjxG1OKRBr7n5JbA0LyC5RTy2Agz7f6FyN3Nu8mf+Oof7UYpG//Cf1v
QhAGz0jGhnZ33fGYQy70L0n3KrPhIaLpEXha9l4Uttw8g4CD/4s0FHNZVXZe
kyZACNWbtUie/16JDF3dlFHxPFJTZTmI6xK3IEYPSkb6gIvzvEOLnPJAU004
MAAHJ+6DTGS2VNqTgN1HDkDBnsiE1h0EMTO2fGCtCUN+qNTwhagyzWQ82E5I
a7uBl3YPfWg6a1d5L1YBtzWyxd/lvoT+eBy4f/PM4iJGFQ7JhAv6J6Ka9CYg
iStQ5WHErVrD6Jyyl+AUAmY4zMP8m2Cmc6hW0lhbMVqI814S1Y49sGLGTWH0
cZJbiPu8yNbCvE+VJOmDIu9j4L6rn1Ac2li8+OkoB2u6pnbLkeVXrolkgVeB
G5xSVfdZrADNb/5L/9RXDDMaCmbBSC5QhCIz/P39x6G1p4n9LYEQkT+WndVZ
r3o7L0Wxw4WKcedc/bR6FR2uAUDBUIit08j8vV1BRual43i4eNw7dTSfFdJk
MdDkXEEgZ4Xei/1TDZ/I5qcEhk+pTnBe+/GlkIVYLt6Ep2f5BN0gsB51p1+A
Gwm6N2+C5s25PSMhzXHoTtjlx9NnKH65iPB/yvInvksS79EdwdpHcAg00DUH
o1L3KfYhGUh8ElF1xVPDZWt2pFMtneseIfeKYjCLys69Df8L3iJnVw6iX8Kn
jmbKLBY7nIniSKkPfIOZG32gHCdBxghbrUiB4oTh5bs88jw9TUZVNlTd91eq
r9CbTIM8JCz586BK43MOcRAMQWgGT6KbcqH9Vtm+M4x1znHC+nf2CLBir+wN
oIi9ah4qZIfIuUFHfSxdenEFA95TBd1fPwf+6q39lUhOmzMdkOr1614s9Vzy
TCtsRlFt6W/uW9r+XmpxtXQ31aIWQqr13ePqNzn28ogK4Dbdhclpvg2531Iv
+VE2w1PfJNXhpkdm17DxiIvrXNgnmQzSgw5fH+3kLHvLjLg8E1BxNK81TuCK
azKc9Yw7NeRw+Pgy8CWNfWo65v06EkLL4i7kRIHey8q/dMMfdQkEipStn92z
hFvc6EgXKmfofqpNJBmsfYq9JAwIPm7ztnGmwWyCyafYdDlmx6J7pJoN6Rf1
3GTZw4tACOuhi84bXY17FeROJvGJxhBCZvDltH77KsrnkOeGyrG7ofOcG1ZU
T5dBJyfFwby8eJN9BqjGFEvAqw/MlS5uYWN+186xw3I+xjeefRwcun6YDGu1
ofAmJq0324YapU5uR4V6ai3P+K8Z81Xd+sFp70QWaTh71yhcQ54Jnss07P85
HSD/dYCUpa1HEnSennImDHe4OIDtPnpV8bnG60MD0gwbbCXRDSCWjfO+ajvc
Iff/VuRSu2tIrduLx8WoCtcIbV910DMfZJvJZn38+/5gsTMKosYClzE+i8Ia
gk9k5sFDA0NeY+ECqMMXNV/3PURdBKi9w0JTvW1y+SJkglfukTNfPvXD913D
NVCdDX697GJta1RYEwHgocca7AmUMOQXBMPaNudKbhPGwF6Wq8CwsGE/dMSq
mU83sm1jf/B1xvSO/80felbofq7GYLiWgaoWARtV2TR7VlpZcxqv0UneHZyv
6Yt0JOdJ8SkvNB+wnYspgREIZXx7GbXY3DP7to+rt/dyk5p2wkZm5t0yafnX
pYwN7LLRbgbdGREJKm9+yWabc1UGBbaeSewTq+307GHDb4c5hUvDYcBx6Aog
MwHx3MGmtrKzjl4gGVGPjoTl+F9N9rynWxZ0I/dBhNsVuXWJjcL9rDisTSJw
rWn/7waDZuqeTHh0I0rTJ54dOqxJQXcduf/viJegCE9jVwFVJKv8U1RX9MSb
HoPF4bMkVGN1OCSem+WSr6pOhoCtJnTT31fg3aq2OrnbCEozb2C9tY+rG1hD
bgVlcvp7c2gWP6aU/Qesa5QthSmyOzVxVfg/YS4OutH5DyUUzTLqpNPzlKRy
VKDMKhGdmbxQy4PyjQ70waZ5wFwPFu/GhjJVFtx4zH7N00/kULwu6iEzyXrp
i/ZNcefJ0uZjwjIDFxBPcab8k8Car8EdV7tSWoTCSppZ/jODkkuLnoZCHZ32
0Fj5XZiPr95DUZBuX0piq7sp96Gh4FDk6p4zJ1eaeRuIaqpZflrL5qChu3YE
dYQwYpYYtgiqCBzVpxSKjlT3FGFxlvJRsJ7oOcLlpf2WrY6X0GbVOnkPkyft
flaMUZ4Wl++3VNLFUVgJF+5Ctwf//ydDd0sjXFRW+bAhVWAVCoIFXFuBBgHa
484sT2PfJZX7gnKZXo+g19RUpOr34U+4ZRlKyZRnR/91N081xO7w0Qnk4h89
QBHJsjg5EL9SMX87WRcfKlZ1JNbAI+kb8wp9Otz83wc6KdMPPm+uF6JZ5juR
Kz2Uvd6cKfsgN1/9O5IOdjvOUPv8ndEkCDU71B5iDBjUAnTSLyD6YxwuMjdt
6vz7ZyIDippyEhgcdJZwoYjYlb5bblVOZuTw3LRiokVMgZid8qarklxLKQbj
hGpcZXNtSp5SDa9qts5TKFNeSy0bMTLtvSJBWG6fLhE+gU9hWb6XZXeBaNHG
C1DNWopmNiGlCNdw9MNjfxIk4y9l0i0/eU7jUOKk96CNcqMNAFbGZBUAizCR
GJxoyi3ml8aPKDG2TP4WTyZEME9dtbuv+aasWLuFQmAroG0U/Tl2uTAPquLv
WfZ41lg8mThU50wIboL/GUPvUS7jpFM6swhIZ9beNS5eC8okVdaV0wZ47GFV
GNrkNuto7Bqqdqf47okHohf5OcI61hciB//ZR3Vrdu9ExEvylDJxBUKW2N/r
+TL+iHssUbpUa5kG8uq+JIZM7zECwtnuPxkeHcQtWBfC5ujs23aAKboO0glC
etB/3UJT0ydHQs8VUOlG7tZkMs0eIAZgqJNtr3DZqIgld1kWllO5Bet5L5ja
ppl9py0ZDADJCkmz0oWmvxGGpTjRnxFAc7DVELY7xyYr7L+no+QHADoqnJ+I
YrMWvQMIvoxB+LK6stl/5ONPIJvdeDloFDj1iIn/Pa+NGTHwjgyAR/Uob/zF
PnVYBJSZSdk6b032xUpi65vTGuy742EKIQqZ7LPxSpvPwsyhlFRBNruhtgWz
TbLux7wKusltHPXPPdLHkeyI/qmbtUS8ft7wlBdo9W4ZTzQuTpEV+6afUQsD
4KUf1BkF7vwso/O7yxamB4ePhUwu9+CHFcsx6cLvWOD35Fe8MRpD7AkARUwT
z7xo4RaUwqoob7yNe2S4V608TWcUlNsIta+PPdOzYOUBSV1PMlsDoq5QLpdq
nYRSBHgBB1EeETwFrX6FcbCkDdwxDTv5yhpRVu6XS2DtI532fLOu4xzeMOGX
DonuqPiaPRxDl6qr/btsG1RkgiDUXhNz5Bd2Nci4CuH7XbUYHkpsPj9ysFsz
5AuxQpLXdSp5VTHpXA/+XLFbfgRLawl+9isSn4iDuikNcnNkX4E12K5CSqxA
iyflyHD7TGJDsLBFYBiocQYA/7cX03ktLUAx/So7SKSBniY9TJUGN2lPFiQa
SiodanOaBlVzABlLjQ5NukIpM2vuq9WI8VTA0B03Y7rqdF3SwhuhSmHT8jQD
ZjwyMGLJI7vlwvxhzc6yLlmKpaXqS06ta1FeVLBQ6yZ3R7/5xvkYOsK4q0rr
Gu4d9oaPHlTHq8TSmY3/aawyaYZu7TU06pW/V6KnGWhVQp6/yDpRq2+RndVj
GUi5ARRBowRCpmY1ole6pJaNMvH8N2iBr7uFFv1zQ3l0JEj3Df3WrACN37wS
BPksbYKLdBd7wxgkEW5t7hyyRm4aAKIQ6qLpqZRuIuJHoJev4I9JkysTxdiZ
WaaqRwxRvAXMwq1WYswFocjmCob1ZjA3W2oo0AfYj1h1NkXRmKlYtTu34dSf
HtB2PHdHyP31PwHc7+2XtJlGS0uzam9SyAJnK4/6jrSlP5u+OQwO/bPgHq1q
wMg9dHn/fbpECLD+W7bJcyiJVN7YGr8OMP71/9ep8Mqf/DZmkD3i1QI89zgA
WX20mhtckuury7QpUihyRB6jx7XX/ztMD6uIi9kVrAWrml4BWPGtWkefNxFL
qxxbGltUNrYwWDrBGYOw+ZDHIg+WKJm3ZNEInC3YJbLjT/NiL+Tl0l2GgXIO
gWTchToVAW71CpOD6Ut8dvFNe6QWEE2epTWeWYV0PZbd5MZcNx4sUHCpmhwe
uEFwyp/THaLxTgBRTgRQ3jlI8nKTzLahHczitU5W8zucbS7p6rSiSajuD04k
szKPAMbx8RxTArGLYyXnCDmI/SeY7SDgmcHMyx459qTsbZu2WhBHEoZ5k6lD
Ajqo7cb/M4R3RII2w8i8fNkf0TTAtqDmHy3Ia4OMrDDeBAMvetkjGYKENWuP
EHta+JsuNO3f2Z/nXpFAYayMwrotigJwADGlX32fm+mp5Ye+98Q3dxt5yTBR
tCtFuHe8hQxxTMpy6r2DbT96atqPy5L5xpD+q8aQXJItpneNUurduA41kZ3t
kv/KWbPc8bXw22Igvw032+U1+o9cM261xNGDAcTN68OP3pk0FuirMP6bvhh/
wiLqf0H//MUd7cyL3yvwpLzqWmZK0KSAt/lvt1cBO+eaZfyFiglHdL0L0pOZ
nFBTJSLIKON7BYhppJ72NTHnVdd++SbdXOzHvHftiB20EjxHHtwn+Ob75FiQ
lEwOZjxnhJW/g1zX7h4bmTJ9AS9dC5fOty/QQinhjpojOEW2umrv4txxnOlc
hYhULofS6juOymAAKAHamERQCq7LAKfIusMLo3Wp616HCxYBtmE+zPujrJhT
lvTcgU4NqppCbxLW8noBFwXj0z6x64KRwBng3zIWPdPk4O6LLaw7bQ9MmYDZ
+QCgeDDmteX5zvky3FsNu7dFBMpdti3izA/2h+Cjw6mJHUTAd06CHmTV6mUS
tcGEOqcJFvUMwUiOGR3OI3Hfj/eN8jgOK7LtcLviQukDRRgT3nR3csCuk2s6
P3KGg28NUxqHMNJN5a1cI1u2HEoaYIIgmg8KZFyejs4ckH/xBXYfTF3GEjUG
zAg69v4N8ukJ3kkQfARdX8gX8D2+ZG2E3nAdD13vhLZFp1TXYbOhLpn3k1JU
t6Ob776HjUt17z0tMFRs2KBL8zjwrwiuS986YrYDs1lGBql/nU3wYyjC+y3Q
RhjN23l2r6Qxka421yoTsCRP/sboultxRnjvd0BBhsbsYTZc23SRwO1ZkV6U
47OOSZQFyykZvoutk1iDDyGsRFgm4ll4JhzbAjI4szLWxxI+jisCjqtcOnnk
YWFHe73fLBujqeTRTmZK7FEAHjL++g41im7ntfNFBYB/8AlUZUivHpBI1uRg
lkh5w3p0i72jMgkw2rrz1yp8xz8MpoQMqLalKxG1Osil2pk2b/fRIw6LiDSq
byC0RqlQzNLrBVjT+9nBRE/giRzco3rDIIwVOjM1hAQlmMbdiQEh21fhK2vl
JuSA4dEyWyEze8SR7nUUXzWqcvUalT0r5Oveae8PDKKAE10g8dpigI7uAvxn
QHawz4rYnn/AVuNsFKE5DKJbomZl00kfI1Opp2LwSiqiWtC2kl2yO5xRGZMu
gUeQBIFv8yHwVKh8aZl4ACRVx42bLEEcecKQRMP+uazJftWjozzLKLcOsIyY
tsJyuUpQDs+EjkTewBnSc9r/9oUS89m3PtET9jWYavjkKtDq2wz0j7eP0igF
5PpvWN7L2gNbV2NzRJLYO1/KzL89BOkg5O698eLfSEL15emAwbUHU1GhSC8O
ogS+NdD4FVOR1+3yjKZZw+2VRJP7LyH/i1I5kVrBHKVxc1uo01FyOumnE9gC
62cEV6B+V36I9Z7n5TG6Nw5S59lpdR2dG3sUHXhgcLlTQG5noP2ihOGKsTLk
td5ivZvagooWInmGsP6Exj+hSIzKe5HnNkklnm9W3ltbDg9h2E7XIZn9Cvym
GZ3NajBHV/vfwsMi/7BMRscFlp5/qLuzBmUtZpPACCsdcIPMAD+9GUFwg/Fu
F4BKOBVqiq1rRRfsNhOemt2EdcCFjHCo9YgCdy7/F2WQTIt5fuowfOG8ZVl3
i3bc+qVoUT9VyB/FSA8J2stny90OmpH8FzRIA+0hpBcYNLN64UlrNVnieN4a
jOQxwjpACL2J2C2nmDV5n8TjNB/uX1M+lbXYZU61C/qky82AwdN2oghTDSkt
nOxujxDMYQpzNojgQ4k0sm1Up0M4jcLAUZLmwd7VQwB7eeumnQj2V69I6gj8
I+GUrbJ/AvtaH5OU3Cds9nHeMblaI/FjWkCcjupUbcUR2vCPHBa3iU1FPtC8
yelS5El2zkm/Y18GQs8j5HuIAdTraUtRjDoQpSzigam7zmdKfQRKB6Jr5YqR
Kw2ENN8LXnoth/OFZ7y5ih4XLHQBn1FIJPDe2+awkKgeZ6g54VLuGZyv3i9I
mgYaFXumQ7Jqf/Jg9ojEPOtKOSfXpZi/WOco7uL/wZFQqAnO08fghLBQwBN8
5Zfl4RJbvdCpuC+k4nB3H60g6ZbC0yTbCslnEzDaF8dfD67CDhFCHE+AxeA2
GXRwZqU3pXBk9KkwL8R/hHOQ8dhNWfUyPiIRjPbATHqG/fObSHS6AnitFOn6
YoklNmtsK4hvKoiCn673z5Xe2F3BWqS+IniRGU1dES+OgBg4qqNrAlS00Ukj
lJ1lVKkR4BbdNhqm/bStA1jJPtWSoD/MYypMbZuf+GLZc7z2xIytTLDG8aqR
0o65sMoeTMsur/6HVGBm2V3ejIGLUuoHIoJlrQGVvXFjJwnQBkHiac3avigG
1xnZvcg99jUWDxZ4yo2/ToatLRwzUrrVavcqHp3jU2pm9XtDqDL4QX5BSG8+
52vuIdlULxJyDhcqQN0Z1HJPIN8uCA8nNXM9n3VrpQQUK+mQlshp+UmMFrWv
7g924WxCQw51a0U3dk6MeGrAc5H/9hSKTYXSUZsebVds7azpSZhTg0G6TEHQ
k/HE5DT3bZPeg7ESaU80UB7+oGhN8177ckp8n2tsqu0eatz64WTe/tDRJich
n/D+dFjpmeseFwwm0R6V6O3p3CWNO3F/0hyt3K4hlcz1lbn+ApmChzKHwBnO
aLHwte2g7+RGL6gMrn/J6pVSk2bS6OHlNInNxf9vD9gMyRIbfiCz1c3ohO5h
lFOfnJsKMfP1lP5xxCwZnjdUoXxijzOZIiMNtvawqX0Clo6ZqeUb5sDvcClm
t8BYNkx9+sv7FsVDI8WMiu9BbyYBKPe1wALJtz2yT9oD6Y/qSrW3e3+tNug2
dTy5xEXGoLbmb2xhe2uui9GQRcr7NSmgNrpJHOjNfaNe4CdMUgB8O41LRuv5
4i/xZw2AGTSgA7R65F6p/HHP2T0pn6+QqFDV/UoiraUY/VTUHKD4s9ooH2+w
05MvLYpOEnRprPSyGmuBadwFujXzeiA28nhcizmIdIf+XTjMQ+k1kC/S4Z1S
YP0YuhAQH8qHgz9AGk17E+9LOwto3LASNLiv/5qlPXnmnFmClToljyfPSzi/
MQJ9Agido0JyE57ChAY82wwrIrlUFg7XXgp4PhLFuh9rG/Ckwx/J4SZR+sKO
oFr4bD7o/tJ1PYTUJaG4xcnCdNfpsRh9L/8C26NX4n5KeQzyRGFFqOMdYzJ2
PCP3cuAMiOSNwwhV5X6d8WtYWLp4maey8X4W0nrwM9tcdltSLPVGLLSioP3x
euuDEeFlLahKHkrRrLfozKstJUYpafsD9ecq2ION3oYRIE918us+YG9oYNtd
4JnT0Gbzw5H95EuCnfBDOAMHV0LSOawSwjRTA4qsYKqzLw7/cYeY7OFhJ9OZ
uH/FbAWOK4xo4J1j0+UmLExPvDL9TKaRh05bFgIV7DbPk7o7nWISAOQqgOxq
TzxQxaO+7fViIm543RQFcITKiLW+77hbMVqW6cbpbkNqNdPZsHoXqaR2QeBP
OWuV1JfGr7uTJFH8vkcMZ+js+165WrcFc2L584moo3uqSXT55xLiz6KBAqrD
Mjb3s7DxK5JpcnOFoGsoGnT5u/Se9iIhdtZsMAwUnVR9ihxnYFZY3oE0UUd/
ZnnydzyphYAfphzoh8vvzFZGAwsC7sD08BHN+88QVt5eHmNIBDxGBjqNBifI
yZ+lrP0iJIWmKCMdJrsMvLnHYmlR3hG5Id8dTxH/CMYM3Vt14w8ON/ww07j5
1BLz4TpTk+Bkt/A45hcFoObC9BeW5cSi/Ioy0ZvUsMZwvQz2Hv74To1nt12J
e3atXidQWwB1/J08U9/ZazgcmkM+qOzWDT1JUeu4uBdy1XU5R+6Ub2Yx86rC
wHh+jzvCEYWtqpCfcmK0vwruklhZCVnXDrJSqTVmY4Nvl4Jg9EBSJ1t9bha/
cgPR4IWoq+hoMK4/4f4uo/5mvE1vaXoYczuB9yYFlreQ5bqUcXozc3wVEoiU
wPH8MPwVc7hS8zehQ3kY2I7XLXotYUIWs+8NOOX0rKYqqFuUgylRh17Wj+4D
ypFOTp43DS4TowZ4J/uH1cyiDewIkhbM6K7fpj0zYTwk1IGGIO6xp9SI65ZB
G2aZcHP36pPyqy4tAhTIA+tJne2kidxSiNCqXs1AO7JV9t4LSCEAPv/25zhU
mVsj0TSWTnOE+dgf/3t6AfG8gHvKi5TAfFG/Of8w0nVMF5RWU6QCzrokmf2a
E4DtgBpusPjjeuEMuxb9K9MNbQh0hhvSpkBHFMY9N95FSsVCSnw0yXS2poR4
i24LTVjC5/RBm+gbbKcvk65+KDPSRfRT5NSMHvUhiwMjP7UG51TV3VkSxqW8
o1BltXQOE1a9FTUKLdqBH3BI9c5DI9sdtkIDPM5pZS2TLqnYR1Ty+ySydNSb
V/gx95aICZtsHf6ohvGNA718iNca4WdxQlrelRMlXpQEiAiCITqTxtNqvhEf
YvHl/zZ3W0vJpWnbxU/Gxl6PvdsZTJJYi6KjWcvcchD3Q+sw8NJHtaJWuJim
iigJrbeE3nP/4eFNbKARoOho7v46gYWwZkiqTvaBFvCDLD2Ep8AUa5rvsQMg
scn441AG3f3l8U68ibrX6aVNy7tCwIVvj450tlfkJjVW9ctUkUtDE1tSqb7l
lpUWyMvITqwtuBrRjiG4mkI0CQ8sDmIawBBOXWO/zHS2VgG/z7XuidCvz6kI
axw/fbaL4A1xuZaE2C54WfHykMKrZ40jQlCiqrGJFajPWA/SNtqHeDtTCS7A
Soi4wD6zdyq4+z4XFWyFYk48+DzliQAfuvfTVMm8pBtEmWNO75/scaHPv6H7
Kmv14kD54WOz5lmejOm2prq5S39VZmyy3wHV8aHsXtNIoPoDegV8UiiM8QmP
8hzhHemA31bZMHSyjQ9R0hkQKpV9NEEh+/gnktr2OBZG730najsToOVQP9+e
gE7k+u0fBoimtIE02z4UGxySyHRPQNw6wH22/xSApImFbSoyQROBczJb9LdQ
zhgY0m2IMlY0UN9a7MEVSkcldRkSJjMDsboEISUmtsDdCRzKQjncjp3iZxJ4
U240C56dzj12c/uenOYbfM6tJix8xAOonzXtM4QEqB0/Z4pxRSHuJP59s8CP
rzVlrwEJ+XNKrM2CEEFVerq7T6J1xiGzWWiQt0RXj5bjY9jbO/LP5B8f+tzE
3Jlky2sU+x8Zt2sOLIfHsaI9SSIJKXfV0kLJxH08/uQK9/iWctI54lv94cPM
oeUNr9GZvenO6qCFJJ6prJqBXzPKQ9L33THaq2RsiSeBRqbs5fYtwokgKCE2
uHb/OQjQ/UpcpSIpxaVr+ySl+IECSFtNioIr+A7/th878Sj6HaYz9K+wdmLa
FiMqwc5kRJMjH6G9zOHkW2z0mz1ioJQ3Y2WWDriMJmRqyYifpk7ZYLVzLKsM
hl1vY/2H9w07G1xCPIkGF8bZYlBFwc5VB57vqM19fHzAZXxBfxCQ4vOhlNqc
EccpqO/+nGlEJXrF6p9pWlM3jwlvKeNM2W4b0tDLUm8MGMIXgNI3r9PokI3U
kwc3xkzEMnirNBORf08lkLzugrrUIZi1NM0MUWolgLI2SQR3nqVGQTaf0g9C
LGR03a2E20flZQgGu/0Jn9uIzsM4q+ybTH4RnVAZiFDRg9SmBnRA3m3jQxcB
9coblLD95PplcYk78lNv2KonOthulX4Fz6kjwuNlvfPaHne2YznHlxoh2Mpg
zhcCZxaWJ6Ayw8j3sM7As0mg5b1F/azvFcnGXxLcVaNaNmWb3KYOW62FSPd9
J+5GHP3GMNXMMR9bvz4AUmU4qJa3n7wKUSqOc4/MHUXlijGNsIH+A9Y9Rg37
xZevogKS6UiriOb3GCzY9Weiv6AKlcZwfluNpM11NcOEIU7Nsd5rJCABqMfK
y8SBg5CntNjLNr54TIA0aCplSWXn0uHyTmQS1vt/eiZEtf1OrsE1KL3uRtaN
LxSntdIEPzPxXowvZQLSt8V8Pi6ql6sJgLjt2QQgMx2uW3YUCJNoyZFLL3eG
Nfc0TmKGfFkH/Vay+jIlLwHcEnXvWxT7en6WXeRJqIEghVzLLa+bDtTucoPD
PXUNMtdUTdzxAjxizxtHSTE4C3/oX24Ew74TfhqmT8dOAsMQAaaRjEjrYNu+
ekdfPb2pWn2GS+aU6vcqB2yQdITL2tFneTrQc2p0jSoep4sTqovp52nK+8wD
uqfEYLoD+dC94r90H6Q/j/Fm2LftnCD11DJYsmtCKTRojGjLsV9332+356DU
usxDgpgJHHvtgOZ7BbLKPJP2BFqmEXAAZL0ngmJ1t/CB6Ydw4gxIhRRNOdK0
zfcS+rnhXrqJDHyjxiU9I7MFtE3jb0+c2rDwo89ESHeQ+UkwcmSrs200qQm2
jm7uCudMex5KUr+oul93nIFuN9+YLprQ1i9h4Y8UmQsuLhseZwwNKg3Stv2P
Nl6fS5bvD4kv29/AJWGeuDHDBYPpmEzXw59EIsbzZdYhQF5nV0ds7OxlHXUQ
LBXe8IojNYX0uHZgvdtaUkqRmTQThUbym2YAzqzcg/PgUJQlfhjeLrAq9/mw
onTDzonKKKfzMwDYIf6T8JrUwVOC/0XDyiNcTidm9sN6LzlT3DtktvhHOVNc
dARFqQ1ivcasNJ/RtcNErpcCZPoUwRXN4nv9WhaR6eNVORUJxEX0z2LhuHqK
aUgb9eGlkII3e4UTr8V0VLONhGBQbaB/hn7xZ9hBBbDi0id171cQAxyV5THb
tTnztIHFibGvXJvWDXY2G7nktZJgvELiUCibCW2EcVqYs0QDfFQ0EVnq6nYl
xPN7bcu91wkT4C+8kNJu0WalJ1Xr8/Cd/ws18mVaBFlhaXO9+fdaX2ZQ3BkV
170/bxuHcDBZ6RXw8BZw/v8mrKtc9/LwXV+4/cp/q/yUf27+EMrhRsrS4y8f
jlE0AmWWARa8xD/LcjQQ+iKB8TpkfWpKahkiZALHGQkP0+MdDknc61exNtB+
oSczOUxSqMkQpGAyBgek/wcaef85piUOLIWnQLBdT8JeFAw5+yzofISaf4lr
yFaI6F1WOlB5a1SarZZWa1Zp+0IF6ZqE42anWFVwZ9PW530rEBjyILHXoJCJ
b+t7ncxU5WllDCvrMURp5aInlUdosLx/BYVhyodx/lJ76UlIS790PYRTrKCg
puIgf+kWepFrZhK+upiiRbovmOGq3FCHboRVJkwdmloPvYoSHrVAwVHQ+EDm
/ZUMLndzg1qP+x+ew3NkA/DKg9s5slb9A6VoebXK5hHDi4ZKGvpQ3DzcYbW5
abR9b3x4zxxTfOT+1/LjwnOpPrYUlwQjObfcj1GhKRa0qF0eTVDAuq5ypxWl
AJyTkXGAcolQuq6YIAnQfQ3hymBnLf+xImtUm4Xk9A4aa9/VyGEiTrlE8opH
yRLkrip0R1NC2MfLTIJvvD8ADO+bQ+rmJXNu5737HF2wWjqGFwPpA/rWzB1l
p06UZ8JW5WYikWPP/NSDPC5ZuxkmsjrwXqPG4fRAtE+D+BTc7PCDd30WWSdb
hX2E5dxB9QVw9okSOUGdLTpRtciFf6MhIrYF3MSlLNg+1CTKVByRrrwK8U00
WdWck1+x/7aQDJ0lMVPXRHyBQh5O+ia87NSfHPPEUmxm/yC0Ew2sN4UbS/fQ
dT3C3U7vUe8o2CQ9H37g6jUAlr/109CeGswQ3tyBv68HdRg3+s+7FRek+KHO
J6wV/hH06bxCaTzpGCHNNY/dbHDTeA0fj2piJMBTJDs0d2/0M6Ri4i+4Xlv5
cAXEZgwr64ycH23c349w/znKmEG58aspTsLiXBPMa9ShMv8kUigpGrp3KTei
ZmzJsoVdqLEkpPwuMwsMzOFtrWxinUaWTrBZXwhXQqd0yfHaDwMn+ESs/Ewe
M4Az8kIdkAsA86Ff8M8LAxnzvEkOluwC6u4b/9Aly12yuUQmfPXkz0iYv42H
nHBSBtvc4Vxv/Amg3EUD6fqEbRz2PaAS9emziW8kUC0U+N7dxUSZD2CyMzX/
Kt0ZI8Nn7x2ybIsxI4p+S6WNuKtFAJ4j+ao7X2QvWjbYBO02proEqzTYmsWt
ISbgSNvmEPhNpBUV4zUme9kK2LBlCYndh9G1zRlwX/LHV44jQp00rmDCV8sS
MySyuxB0hlzYUffER1v8zIuR3/xZJAnjEwPc6MPS5wv65V/aWN410H+iOBy+
AJSRRr+nmKrdjnfhn8Diux8Zv8/WBbEJdgxXDe1cfDk6PIjQ1tM0f3PQoDyA
4w3fR/j9T30Oa3G7DsQh9CyV0ktYzLxoY9iP3SUdy4DPN2lgHoUEFiLzlaJe
Wn9LzMJOdPsmtyy+eNuE/yzCnOGNT0/iSrnL0o4rRSv/v+Er4Zo+LiJYO86c
MiqaHVv+v/LjF0UkMceSyIjxgsEEK+6IQ7nUJanagnMfgYE4kOagky+GGMxL
+dOx6Sfsl9V2I9RLqvFxChZA+nN8Xwx5XnCdP0TpPOZVB1pczmw/Jjxvfotb
BY6IRLh9KJL2HtcvRttyqkqLisYMdkoz0U7pxgLXfkSZKxD1Xw4lqYmPe1ku
+xxEESpi/BkV5KHZW+h9EOIbOXw4y5Qxk5JR4/AcL+v59xvhiH0d6yR7NYig
yP2b0Gd4t/hUF9sqL4d0ib16vl/5dWgbo3SVNgcqaVtBh7hHWHYDnoYiF2AP
jzLjpgGNXS36801yy095FuWICgGI1O1teHQMLhPZQdQWvbXfeVEY0rIDIcxc
CXRjybBZIY/svdOMQJQFGTFH7wnhOWWQxMqer2vs8R6u+brrNLDNSbWcdl3S
QL/W5+vT47dSN6Z7pawWE8sVSVTfXg9SfEQqylgYydxvZCUXKVsvZN/tBYnB
EUc9dNJHoEiDn5iqkvfyOg/XQ7OPtQRuXY5H5g/aouURetoa89vS7/QQ7Lp4
0D5R9Rk1soIz9M+1dU7UCwsccbEDGShQA9j9Ax7c5mEO8tG5J7jmcv77zO8t
7xDqjf9b+T8Ogw6c8uw7oeKV4moWsHIbFv5ezPYUkV6Ql/L7UsG15z3G+ysN
tSYoi2Ksm531pC15aI4y5E4lzgv6jRGLl3gbrqr5ZwPKxHp56z2ByN8WOWxX
labLCqTWVlCTmGASUKZigIdMjCIssB35PJp5WUtIauLEq53+l5+3bli07O9p
yN3xBbUnx1+TMjb43jYTBpu/B2dghUdusZ0PLcI+IirwEmReUqNhyj47Wc2E
RtS8mVDCvGI7McQkDtCaTpUiVeLwMuLnfccxgfhZn/rvylWyD6FiDV0qNgj4
joXpNFbV9toL67SlL0LuRb+DjGPhkCFtlScB9iK8S+zebIMBsxhCuNR88T27
9ecRCcAtprBXxfTXrQlMRknJqfkC/p8D0st4gQtaqPGoEhbXVavulBDsDH8B
ZNHw3PTSSlbuecKsYR7keeq2eo5aMaqs3qf4H57zLRKqcnO1f3x5ov8SMEL1
jc1dX2WNHxjr4bRIEaV9By+TU8a0cnfl+x3MSZlSqJq0n/6GEpnau58E9BI3
RKfc0vc2S8vjsMHaRqYdjnlRF88057V3t7o3NHyIs8iEM+0iHc1ITC5ZUaYM
4bKlCD1PxvQQuOZAG05p9zHJde1dBnzxf0ZvUI9GlF3OC3u0RdkE047DooE7
GBpbkNaU3yScOzrrygZkRtyB1cKnk8HmfelLD8gDr1OzyQ+VjKkSuIFFk1Rt
Qn8gF2GU60BqEm75NdXvYfBYvdj24NKwF+IQgyz4BHLicdSJXnx+lQ4ToRLI
MG13PA8ljhYAPX44O+zJJVFVs2PE3gWilbtgsfXwlHmUGwYCVzt6pI72B94P
9IQlo3XF4dVVN9qIeRcGhVdW4JUQcVDghRlrU438U4oPe07xYBRI3E1iyd6y
sbtur4htw/Ln21n7nky1H/dqxHIJLPe4ifiKRGmBSEV9CTi20Tg1Qt+ITWpf
VFhNY5JVndLUI5crm97GJUi6yLkhnU+eUj62Rx9K/OBy0clcRjCbmiqBG5BK
kXe+VF4HOP4Kj6gftpJODsLME0UqVIRMX5HXuZvxrFCYgaNTCHRO6jUSpzjU
CmOghBGyt1j7PPu1k+RyoSsuOZtoeCqBFo49+o5AqYi9Nzcincz3TtrOx/Ae
WDMZTwj4WUgF4vrpcxR1Zwv8ZenPBBTnqCEKfVbxEY30cwqZR7LPwGhvA1RW
mX3KZjjYc8ZwI3+Z4EkI54SdYh9evebMf1F5uKXReKjTdcMlfIrxhlLAj7q/
Ur7zMR1KP8xEoy0VY2TtsjAGCDLt6wGFPVXueHoMUZDw87P7QRRlzJBtvxN/
cgjSmaqKGB78TW9kfMsyK9wQhE8XINQHjfRcxmxs1Pc7OHauRpsAd6UuguDW
0RqL9pdQl0D1dKqa8ZckWnIhUgNMBQRFhq2Jbgfq0tvRHRBcl64rlGDdQ6+P
FjPY/YNbB29MFCJzBePd4b3r+j0BbqPDbi2BtvzTrQEhU8Q7vnoANN5yGLQX
e0t3eE0ppJc7lcHRIzEr5HvJiBAefPqrQqOeGlyRci5q70uWuNJ0RdE8OI+y
oYEFtyBGWF/eUjexouk85JaLzZfrCqX39ty0aIVDnjUlYbfofT8942sMAYYg
8eA0ACINWEJ9OzXHf6zc9a/l60MhdOI2q7AIjD9suSt5UvqS393CJFf/zAHL
n0oETUDNUzJWbnUy2BGnN2iYN4UTLPwqTKe6vtfvJ/kvAZ1LUMlPMLsqV28n
NvlYCAW4Jq/Xi40ES5L/2bGXKbm+T6J0m5VzqE+fCKayiuw+rpsaLBkgxN05
Oq/WxIzCtNTcfFbo7Ml4h/pLdooIR6/5QTnB1GpoXTJiVtJ58fzlvFGkc7FG
rZBm+/BREeTKhCX7JgVnXOMuASSPlk1klnYDrjDkb4LrEDWaEIzQbgMpaHWA
83YvIFFzIx0vxZFNVUX/lvORu5bm8jbfwC1U/q9UQBXa3GJH1qb7rf9hkAH7
JRgf0NZGwsvPyRdNZ59kqoqD5RzvHGGFexDf2zXDKdikTJQfiakzpm9bT6Yo
bHiusbSGtITiehLcdEwL+jATCoSfoDYAxJKn24VvlHhUqlOUMZA1CWw1NBW9
ArXz9yFEbZ5qfbiOrFYS20nNg8G8xZoWAmUtT7WrgWF9aMPSc4xSi0ILWLjR
iN1bskQVU99Rp+XbxymZRTI+zMB+htUBUko/A9pwRv42nSWYPFl52gsRI5Uw
ZCRx9byXn2AQdQgzGAl34jAVaJuEs7ZAv8V6nqvgfWYXIVeI1CO2KXxMQNH5
g+zUhWAvQhVEKLfdVO/9rMGZk7+6Dfg2XP8ZbdPgV2NDItEyPSxT7MUEWaTB
5CdX+cY9x2d3eVUEKGN5Q7x/BERWGdWC23SZs6K5Yqv2Lra8xWGTBTjS2oEz
KeJdl1F5E+Kb8Q3U0F0jMbCL3xtMjv/Nzh/dDlmbMHN5Cf/JX2d4Fm7xNBu/
ijbYdVbBT2LH5p74I8LvQy+YE0ug2rUeA3Hg5NPDihniqOvO4aeua5ixpxGI
xG7veuwOdhd9zGqhHJ+PrDvh6hHP+lJlfIBRtwlzqI+S0sgDv/q8FH4wUU07
rCofNRX6xIh1etEWTDxqfhJ64OV4hJy55ME2f+4qJ0IVhYXoBvhIzP7Tzqqo
F3oQ+9sotzF3dXvQWLYtRX70epPAwKE28Bf3W+sRWwMr18yzeUnZ+ahIICje
q4S9JZa3Egdt5mixdNHhT2eHj7tJDV5Z+ovp0jSitN7azJTvC2/TS2X2WNrV
n7BxmyTBGMvmlzwPOTLJzrNULoNXcUtVD6pTA45MEnVaiUvb1T+CDrTh6rgi
Zit17FxjCXHR6TTJ8InV+OZZ4sDx0jfNKwC+acjqGgA8eQdsqIbkohlUpenS
m9bo+v1LMHokGW8jvSRmK76QMsHRta/vGeY0b+pDka2B4a2ebWrvotDaCXwW
00nDGqRzpIxpzbhxEDu6EHXfT+SnxtCCj39aIYJeHnokaBOj34vf2zTL2RVu
j8TSiYgYe7MkRYxmQJ2Qz9BRan0r8M1N8JdEmSYqCAmzkhOcpD+5f6L99q5v
yjyMQGV2Jr+ZDkLHjELnJneE193fYuqsHr9QGHZfpW+ySFbdqmBTup7moUR1
2X+LYnxP/Kucxr2XPOIAXJMEpZYrn/kwkRT7xxwjTaRGG7BFDAneVFIRmEIE
HCC3oU5BaZgOe8jXyhFogtXbNCzuDHujj7uO3bOrdoaYFQLqbqOq2xghtdoP
gOgbwGKQq7KTdyUDCPjNCo+SFVjxMAvWxT7nLCFqVoVSAfI83oqzGmThY2+d
lQb/3g5DXdZGas/uAA7B0CPmb0bvPxyVAzIwEG3Zgfg9zHkBigV8cdW3XQVW
GQTEV9waMzGYpjRYi/lZWUwtB0Koujg72R3ETAdGmagLkNvp3pjN+R46uagz
/wIShaK6/p+wFZwmdiiTNUnRy1IBBzIwYhEzBEIn1rZghou7vVVzkBQ1r1cr
DNl3YOUUgMsyQPZUkJmHIFjL0GdQUCwewm3M8x5pbl0C/5X9ILNX2ZEPPrlH
/zotaVgzCk7h8n2OoVdKv6iWpxg2V0JdhWPiLAOmpZSaUpLtsbOddhX+zHyD
mRoFO8pSxGiqWl4Yl3ZxUTKMMIKN798Beoncs91qYY1SegDMJbQp+tQXAjB8
bBEX+JjduBS6R86UqkOr6+D5TgbqiZPtibLGoj1ogSS0E65LwmP7btw25YYB
8qHeNkT0SKVykSHyEVK69Vh8thJ7Qgv4DrCQtcSYbdd/O2VJ+1SEl9JTqkhd
81BPbXNhzfSlICWAc+xPFS4F9TVdR+V/c1m5eadBMa6RfxBg8eqS0CFVx002
5iKELz4SUJcuf+sFZ6n0MNYXa12jTjDiJrgfNGbqSJXMqrmdIKCTywn5tY44
/s3l47BLVwdBG/2HppXRsEVo+CKN8gubHlqyvKqSSsglNqwqXILGSi1ES6Qw
dPqDI2wZjGVNC47JMzWvyXY6TcI8Kc8xe1YkVQRweYRLJ3tBB5mUK/fvsJjX
ysKnZhGIfgVsjxudWh6Vdt3dcSXH/mmPeJ6R7ue+43yTbGVlvZerGuRwICZQ
Z3GT0FuXv83nk07yJEwfU5au8TO5dU61vU2wC+sVq6mod9jQfhHfv5Sy/OnJ
e8CB1H9s8pNK3vbVehAMy6ZewgSJOsZmXzezeqDKnX6UG8jFGDVOzA/j8T+Q
ddkH0mpZV9MvVmfNkUUggsNzvBOvCE4XDM86JzOPOigRZOzUi7nZ74Mz0adk
Po84R1aIQAoMwVb0SWqqYkS+A/+5sl5ei6HEZUeH6pq/pIFZD5IwT89Xc9fE
s6Zty7xJLOQ3jUuc0p6Jnhn3N8dPTrLn4oVq4E90uU1PILX3v4gd701MdSe4
ckMBKNjE/3fNc7+LRFRoee5TbyZxBntQZbfh9U584WaU5CzOEmwCZ4p27rnC
BX1oDzZhqUWp3lDaa9Rb+EsESvN7GoGodoJvQ//MqKKiR472LjAK7YOLPyve
QjUn5q7LKYv6kEwaLe57K9SGJHNfog6y2CKe+o/uiW4s1VnSLCUPds+36uXZ
JaKueoNxYg4hia+nj3TLiE+PfQOEYAhryezxWwmbDsYSkzQO/35oN2OYATdo
BJuTPh8j+DBWcTUYWfGrZiSI3m4kMH+x+U1gZO/dJgCmk7xm6xIuutGeuvpH
JhxheeLsGIZkkkKJoRso+rQANfkeQreh5cjWRzqHQPaVYrgS2Q7sj4oTQI/C
89N4BCCtIIbplap2FV7kthF5EJkNVizqin3wn2RfW0onaPddjLsOQ5MDFzJa
bNYShZoRTo7ipa3+IHLR5EZDXwdORAKodbczfrrxsxuhF1nCutxZlpj5m3vS
ULfEngqI0Kx9oBUKFs94d1e3AzhUg+iRIcc6TTfaRai7iisTCCJVLcITkEB4
zrnDGLO7I/a5zgoJ6+euYYpr7eQ0W+ZLFA/3KeaAfYiEIGlUcc3Eaxdux9ru
sUwVnBc5FRsKYCVYPuw04eZYmjR/FQn6oL0c4kpPGIPFKNz7+voYBqZGHkPd
esM1U0dfJvt7hW+De+kIiRdvfMkDEktBKevcpeyk+O/eVh7fpJty/bPz5zMO
XJXDGTVlf3FdC6Nk4U/7eDLs9CMLazRvEd2Eq80DrJtzihz6Zo6Dt2jl6Flg
g1wT5WYM2rb5tSKuLxz7IIxqdPGszDIQWo6cHhQknPgfwuanF5gfF+fTIm+X
4OJMFaz1/KL+yiSFzSw0OnFIgkw8XhYyiCqb1l1Mar0qk5rzQ8zl4bo8LOw2
Hjzm4fvA85PgVTj2HXPVPXdSZ1aEiwsrjy/WHem+yoAl+jkGsjKTApDP/stI
/Dwgdvo5X6Xmf0JIdGNoFPXhsJSqliVqg4r/7dYXzJVX5sV9fXBJni3vEIrD
/f8Drgek5S4QvTDqB5uIS/DwVZEGdDNU6B4irDs7GC7lHrAuIryxkgnuT+fU
AkvKEV7r+Aoj3vGv0WHzvrscODHV3Aqj5Hry23kASzhD4UwInMY+MMZRzg4l
lAznq32YuQhFuCe0zTapLP15CnyqD38hlDmkUTnlnrIvLS7HDJwh1Rg26oZw
q/7X7TJ0pEh9LRGSHoGo7suKJAPI8wv08pJVwrCXoHfkSRpl11trwTHocJ+k
IigP9wOx6m4TzR38uba2qccZ7bVZ4RUL0yTBmHnQy5JlmxeT7NEu2712j/xH
RaPeGJldkA7/NYeRhDhQSvQCqjfnChwFKOSe7gXRLyZ+qwyI3V2ruWgY2tO1
JfN/abjlRpoqLf45I9VdJTMw95qeeHhCLLUiWxTnBrgTz7J+mKwspMbPmkVM
gB1Ib+t+yJy1AM/NnU1hOlXcJKW/w1SEcntHdAA7zL7X5NhIFNhiXo3Ot6N7
2BO7BP0cFTVQQtVzNUiYBbo2xaC+6XL3lv8zCwfLQtMDG4RjlXVR2BE6RKgl
zAcPHGAdV4DxAKu7/v44iaM/DoCpKidoyJN8w8CPnLCd+33FjtazXKXKJIJV
qZ4U2H/GIpkJgDsbJEvYFGDEl79zwNRO/B/5JEBpbppBXrSrrvhge39OiM2O
s2GB3o8fFeVIyCIDApp19GbzNVmX9emR+aiQCYrvMLsevArh0oRb6+yHnlXs
7/SIQDpjI+HLC4E00tggITnPesTESihphr4f/ztSQ5ddPSPHh7YtKq2X8IhD
bo5uANFPmumN9kKjzQIoE42zoMsSF3LnbselYiYkAZ2mVkscOUH1mJfoVwbO
aKtWJC8yfEol5Py5COt3TbIDvqvukMZ8QESwAN9zJn52p3XhGwo1SgGgJDv3
2LDd6tYh3I5zE6yopaIAIfcxrWki4OSFRy1XUFju1XrCI46HfFD0BO/Vblec
eIiv8PjEKFUv7q2oxADZ0Lb5AmdkqVfzXhdwgXKqFv7E6rnS2yozAmRU9Un6
lN9me/eUkSOnTpmwhWPvUO7fVDX8zGS2g+X8dB9/sgHH3R+1AHgid3xRcE6j
YbIwXanIs5HTUuCf7DNiiuHZUnQI5L1y2jPsUnbtGc18I3P5RN53Kz1d299y
IaVrPpBo0vMIxknaCqC0H4aqFBDIoSnLozxn6TdPm67jWTIcAOEKwlyqPB+c
3OC2m50zSRUkHIihSccy1+4JUmsuP0srz5CUDHDjTYu3muUNCnv1kGuo6av0
+zO4a7ATCcCNijy4KANx+qbFZpYJ4BKpVeCrvE1SjgBEf2R0yJpkg5YyN4R4
mGoCcv0JdBWiJXRzIOQvx9m5/MGjv3HHq77wW159ai4TfLO4Q2xypmBuCWfs
/feb0Y5DZs/KSfNXE+uZRcbaEI4yZugL3UMKAiiR4RKd+7Fh0iVjBYgit1e9
8hxp5vYeuOvLg54WwfW11JjXmfu9r4Mp8mKAgAUfKY/g2wxLZJ1W8PXwSrCq
1+rG94Den+B7MLkz4r4YlOmLtmvUayBAo4RCf2J3GkBft3KIMyHTtP5vLOnI
BNFiFZZ72b+vqfnLmYPtfR4u5gmujJtw+iaQdv/Vudo/qiQTpjMj460UF3jP
S368e52AJ49YRlVh5TNqnJa4sBV9IQmpZ6qEQvxK4CvpFU+mR+Bym2g2KEeu
poJ0zTDeRWmTkmpyFe0kCuAUUvOt8UUckMaysC7dR+Keq5BDKvaMdjzPIv1S
+z/rrRwiuY/w/0JgKAs5y7rNforOWAiC3Z46mu8j+0iMV8dFmY0gCIGSLT8C
u7GZa8xBWHWA0B+4/Tqs4N9MS3nXt/dXcjSPTObQ9hlDkYkd1n9w9yV2EqE0
RdMJFXEW/XqEJvMEMxlACbdyTgsuyfhRQXXC8AedDEd1tf++GMYM5FiTCfU0
yD/cYXZgt+BcWx97dhJ2HHxsm0BNdtxK6h5C4e/MTzTUKDqMN1JaRXsobccy
dCD8s17OqUqEGtqFN6GSXV2OMoKnpW7Xhl07B59q1M4WXahe6l29GpgLhXu+
dQqFogDisq9b8raGBafm4hb2q4v81lHk4HZS54GETsYos2UwowtQLGfRasQs
7EclniXQCx5XkMay3nNkpeb2k9yeZXBsvy13tm0ElJWd7Mh9X6v2l/QwIdoR
pS8FTSW/Z2NVxnDvIMMP4MEVFbQKltFecZhC/yKaOq4Zd8AYClHUG/lSr9zL
DEa2pf1fD9m4bFStNhftCm+k9/I9uwcIUygciOIeH2H9NVk4rsVywsWbN8Hq
9o1f6Iy4r0XeTEJMj4WhSXhyA/8yenGOLsXuEgSzNrRYRHgqLg/Iq3S1+gxW
i6Vsz+f3fT782v+DTjHjcYuCrPLIeXcFs7Smffy/85jdDJdAbqTxM8ptsn1Z
rTLJz/doAX4l2IBl71Efd2i6IerRD8VTezeHSCZ5HDN6vUBU5IJWjnd6S/TC
EK34fTAkKCuIB04o4ZNJ7MWhDyeMj8/lWNHBNjWLDVqpBG/YIMN5SX8dz7MU
YKL7UEoszO90cHAKBJWN/RXUpiYIfrVIxDGMEmcZ3GO7LPoJXK/PfnWjbBzC
iPKy/TCiSf1B4Qtm9iNxeuqU1kbtqLAeINhZUn7qG2000ABr0jLS9SRIwTNL
8TdWBQ7RxB+kisFUYtx/4vNe5b+a8Jo1rak/9TTnd2h9tP3ZhLXYv4YwlBnd
QzuJHDKWBziZxGIKeTPCGU2eAjThGo/iggKfUwqNmKOLWmpi/KUflbUVK16Y
50nkSJkKYFjf05X5wa67DJvQlge5gC+74HoHiFYslk0+DYqJo88VN5PV331S
oDtUrwu2tvnZnpzZT5OMbRQj7G3FaM9lo7nHOeQX+eNa8z19JQ8ZQplUWWqU
ju3XMtJluYZ8fG6D3WkzylZvJV0TX+ePhqpalxydzeXocJNbVseWsS+kL6Jg
CMvT5LDH598H4XJrG/jC8qOAUqTwjQqxyzerf4bO64kTLXiN+KghIYMK/Hdv
xm8yW9vZ5QcXNC5vd0EZ46VhC38DTADuUTI7g51V/+i79AJ/Gyd9nfb9bjle
qkPx4YIW5fpnNekmmqwjOw3UU0yI+Pe2bi886k061HKO9cm71WJGtkRIbGQh
RBgnI/cxk5RlswumTbkMreS1TT4V5fgMlgvgbQ5Ne3PzsYQLV9AZwSVsSS2L
DQfhF0jtKoIbNGeXfneu5/+OhEgJzP+2pxAZW+B5HN3iyftf3/FmFC/3/cnF
J3v7VICIKn0Yk1+BLT9K+/cOk8xeiITS1h24NN2y6ozpojHV++1yw/9LHOgq
TkiVjZrHDi7mvvV9S0f26D2KJjzKnh8nUxKlm3QpeZTofzUpbNyn5aVmJXDj
nk0xXYmm1YiGeaOa4qp/vcMqM/ussKiqqWSDney5bYicinODr7G3tzgGQvCL
DByvX9/fNJfbqUxUkXHJsddvwPDuTefv+94+baKbTDiwxk6GYQUTEvIf4dXs
gMDIQ82V1Bnt9w/OLQP0rvNaemM95V70C+QuXm5XrrkK/EViHNlUHmBb8Vcy
rPoetf/zvbVzehKyx06gsAvCcissfBHMKepXClnwTOkRh7HFfegyjkI728fv
/afR9i/pgukSKD/Nnmu+kAeTSkwIDHeOa4YRM84ZeSDu09b/trWxnQvMhPjx
I/yzoaVLHKBHK2L4Y7eV3HDCf/8z3U7KjPpPj9wPTcwJnHhf7GbOXO6EEMeM
1QRg/YqiMmXmwd2xF3Gpr49jdW1R0n6zjDf+wEv7B2D3xMRn8O9505gQdrc+
8GVgLZbwJaUKAaF4hEnAahBD+/6gQNfdciddurSEmrvLGFsNXlAXIzdbbMSV
hgY/PmCPSieLqAkT5G1tky6ELLtkxG9A7mIiSNJHixW0RwwgttgcvhSDFkVn
74l3gol1rVP5nkEbxdI9AmmpcL5m797vuqRxUtforRgd+PN0HLL5kJNyHYLj
h7DqnjEtYwfAkKG53JdjPdRs2zVl6FItpDWj5WmEST9vobnSzlpx38SJnAoe
Kop3af+k/D0LbQeVykrTyEpgT/gyNXSF32NkB4WLuQXNHLnJMJuJ7Eu9winm
GGsZ2IzwBa7R0JwgNFB7c8UFxzKyiUZRPY+0bfAui4mxFqeBwiX6ROfqHZ7Q
5w4SgvzsNU/kLXlaNkJuKq1F0BYlH0ZBnl+UjchkrJMkRUCt8mEVn+HOBlvi
8vE1ivRDFZJ+ekIXf5g/3VAFcPqj74qHm+26KJ37uCqsf5npOlqdsVpyW2ns
TYAhT5yB/x+e7IeCFaYlaN6U1VagcpTjgLamc9O6lgB6YQxnznAR6xD6FStM
+wujhwIrJhjzj+sfCealLDOGLJiCHkWUKw6cObwzBRVpjHlcCTI/Lvq5mkBV
cFfj3plvm3z5u6AeY8B42L2kvTutqTh1SA72BrXWLraMARyxoEnrOESbjsug
ZdX7VmmszUDfoxmUMH3T1irmssIPRPIHFTZa2Y2FnIoftqJk6KPwsJMJF2zh
RhhOhVsDpEqCcwbrjaWrloziEKb0B86nlxhA1HeQCMvytBJgNZ/Ik48Zdhw5
elYBMnHNN0IxcXE5yIvwcmr0meRVy5eWYqCo4pspcabHgesN2zKgeEXjUPG3
NL657hpzGe0RQQQD24zDylLsP4yBBBw7LTZEbqdRG8hMakjD16WaFQ22SJCF
h+c2yqTAbYTPdfNn6GYXpqY8T+8o2yNB/awE8m9Jq401o+N8nftxt91yF3uY
I3ObI42EStg2p8qgSngJcEmcMJ2bcKlNNi4QPanSTUYAQp+2Eq0O6BLn8ixJ
s4TccvIjlq6DkHJEUWOJYkmzLNLbrUFKzYoY3c4WQdd22kyKvmzghC/OKWTG
6q0qo1rfyQbP9mo8eaD+yM+CnsK7+L/uLfoMWnvDaSHq+hkXcrHNgA9tBQz9
S+KEBq4EOaWFxPIhmVXnRit/jATNK1M/6bG6lpL5tiVSfCGxIqtAFyeV/0/h
PejDmicnLWCePBVtzeYKGvK+pOdbKzhrPUJH7Hh3/8YQiOrO6DctkM42pNQB
I2eV0tmJ5gQlV1nR+yAU8yR6vaLkZtgNbKAp769w7ZSO0EC/v4K0jGhrZrrj
4oi0If4Rk0vVDOCkZubi8sE34GfDuJmxwnK+UcJNY/jV0wygKBXeQKedhc3o
F0JOgCQCUeGYnFTKbAHD0bjABxLWifVSVFiq50p1ao6x+uEBqdc/N8oUwUAR
GpxwO8jiNAbVg0KaryueN0UhxIb7P1Old2IyEYZcxk6AUkNGd/jjUCw+xQzX
ctp/CCk5RxV1e3gwR+UrlR/dEwrZes2xUSMBREYWN/6dluuUBQ9+94syv7eL
BxKBsMCO5IGCApJbYui0LFV0oxxR8uCr5kBHswoHqhfSeqoisIGXhqy3R9Vo
fuig5yDg1QnHkFSAm4y+o4ouz9o8m/YnlHaQstGs0JHSexfbhsPF5gKUCbXx
jdZ/s2F/bTBQ4x3YsnPlCEoN8VmZDnuRtlE3Qd2BqVc9fTB9/XQoTWu7wsvs
yyc8q6b8T+hcsLZz3GCOFxwqisv+dHulTCldMrxipqV8dKkp5DOtYEcTRYwR
3Ck/QS9T6b6ddkEMoB4oMgnDi0PCyA6eYSQhu9izdo3BES0d5Kz5NaEH+20r
HrQKeZ+jWiWB7R9uo2Ly8arTo2WwUTknKe/o/Ay5LT7nyRasX8x20AO69GVi
GYiw2iljuVxivxUcPJ/mcAh04XN0L4YVNh6f7rKOLm0ujU5GML2aGWGBDZ4U
7xVMNYrgChTDhf/vlvtw1oHAiiCipHt7yJgQOLmcdLFR4Abtap+rgt3GSBdj
cCz0312SYmg3HSquB7IuJ5tuYSA6UvLIJedjK02+AgTkmMvPL3ZXgtaWEKJ0
H+aOTb8WhIyz4XuPSoSSY9MGEyXuHkitDyav/3/6o7Y7trDjJefNuurc9Hhi
kS7wV6ik6ZrNvTv2vMnOgIUPzwpW3sxu+cxxzpt7SbzpegrWg+BvQ9/nU5oJ
lyxkbM02l1nLrhsOgbe5lkqqUVW59tYM+RbpuSE4/l9M5yReTup/czCtO3J7
BxIcq5HVaEpYURLt7dFPlEwWPm/wyGrOXo4I2ylMBe9sdaLy5W5DaOO1YcB2
A3gb8hbXlIAnpgo8PpDglpO23f9Mku11Bbuy6w00dWjafBxThu5DxKWpgMu9
nj6ouIYrfsf5ZtUJF5F7kpSxfKz7qr1R3Y36s9hlRxuHCW8ZhMcp9e9zxwcl
+l8I8V3/MTE4abw+S3SQb4zFe49jqkLJBldq3Fc/d4a9fvv6zrItggT075GY
tiN6mrKdNMezpwplwfBFTkPIxI/+b2mXnU9ubbzlEUPFZfFBdTcA/VGEh4DL
1Vk6t+yJJq7ITKBIkdOYtnF/hJUAjUq5Aap/7QJMC0IOYOdoDm/aFOiT1Kpb
NKYMMyA4o/Lw5Wv9zpZSJjikgaVD9La7X9JprhQ9dtMI6Csc79mIryqWR3e2
k8PHh0EqKCO5HiKc86hdscOxwPtPsCMj9RKvmV1abMeTI9Nxjhd/bZszBEbC
S3IJugXauPoNJSPZPWr+j1lyMNdAEPE9hur4uEKAtYJrbXjn2PPwlZDk4mY4
9HwwpX54QQC4IbPPfMCLvOLjddGj3wVln+ecJMp45k2nAD3sEFwQndqQ8EVO
rJJmpuwIl2fiKIZAOIqQw4eYnF2lJ2MzWU9qj3m2bT2pG263kE3yOmHGKunb
vvnphxnEOXrYrQH92VPC8UMTXokCnRji/Vw1OdHNAULn/+NtzZZpiUdalU1t
X0ll/L7UgUa5ygIO2Zlh3nlP45KkM8WaD35IVuHFF8dqwP+tmVhCBr8gm1HJ
KCCD6w58Tvqf1f6VEvH0iVy/5PqZs1sGAwPUv53tv7PHXLV5zW3Htalm92f0
6EHPe0XnfoyBF3yVQYwkJAd5NkS57OPHhBZeZ2kIiyl81mmwsKdCFx3gQ/F+
2l0CrB4GycG1Z3y/JayAIfX5987YCJISbTeTfpWXugcQGbw4CRP/xUNSS1Vx
RuAL25HngWmMSX2qDVx40lc/+8lCCmF1wc2nwrXKAOf2FwyuuRPWkAA9Gruj
V0StQHIG7gnS2VcwojbZhi4pW/85sEezOK5M4wB/zX8C7tYUFrvpRJmQRL4C
Vg6Eq6zwdGSh6jBYneihiI3jz+lEXWO/+8Q4ieYxN6pwQgIaB8IPw2xHD5qg
xPysGhd6vvm46ocVAVjuksfoVEZgOYYZm188JJIahZVQHNFZuw/irpDZ23A3
azSGoFSWKjPaYSjsu15Jpo9UK2rG39ZLkEqKMdf0nGmgSPyeJvYc8WuBJE6A
s+NC5/RJTcw7otw843n79Yso2fT2PvLxUZtpLSx0T++151ghJDEVPgc282CC
cK8s6TJjophsyJGEXI5yrApeHw5+oxQQKyxdNcwRoi4uazEO69UFVLct1tWu
nMbjyypUGBvKtoOLzN+5WIj6eSTNQp65+r+Al4l4nBzt3Xz0xZqRbHrB9mEZ
FwyIM5jdMs6otRRcnPitfYp1k8cCxiDdMY01kfX480vHWunj9hU6YBDNCr4E
PQVdNUABrjgRk5cHOhGFUQoK0P+PBP4gU5XT08iVUjKfjkYuDKyR3KJW0NKu
q++Zbc7MKs3sOdbbv+VCPEbhzShyMTf3nttHgs0dXRKEbSsk01aVQk7jlKtg
1hDVsxJ9us4OiOsUhUuLI9veglcg3AT1MVd1gQXz4qXKzlyVGfh0H3/IJOu1
bUB4lTRw3anPSYN3HKdwSEKZDU9TKDMMwTkZLeh9Uyjf5ohk29r9KNfdycMe
dOTTLDLIfRbc0tXQYiCRvqr/gm9xgD9gh5VlPdyYofihq0G3DFRvEGKJyyFm
CUz4gvnyQ9gBwMc5cmF1jZhAmFa8iur2GG7QlWOSQWgbxXo1EVj/VK82/R/Y
VvgZL67ioGy7FTmy+i0JPQm5GGUaRriD0xxYPVTzFhTbtfR5nY/WLbtjGVs9
qxMLf5l2AWhcO5MExBixZtJkP6EJKoRXVfZrUGCoHyT2HbfWGjVkv6KSZh0B
ITdgZbtlMqIxbYKB96moSkFb0JlIxsQvbBHx/VvxIqxG44uLR8nWtYWnmawP
wTh/TnW6unjP5ak4hLsVLte7Di3CUIX1L47zs5wA/+XA7QC2OTY4eZKKWUGj
ksh8ououALhdVCNlBVxqSVXFQirxnzIH+w9ISDiRsZV3lArp3gneg9vXroRW
u7zy9t/L4S2BvOiSJJ9/jfAzVsuNm1aoetjHTeeqCGLdcEB46/9WAv+QjDqf
VKxfAlRE6JK/OyLIn5HGCK+GJpxlKZ4w8yD9pHVzBvdl1ny+bkW2+rwuiM9U
jVX2PFlG4fcLIQV6v4LZy26eOOdYaNJ2+1k0pN3SZLsyLnl92Sgu21PWuPBk
Y6nYwnoIft047Y9abaCaVsWDDh/UqEq7ifOPfYBniYe7pT0p7fHVZ4cvBEY1
LcNuCZtbuDOHrOC4Sk4EF3uEP37WPDRFaUKQNL4GvXTDJdFc562yPWx/bKpl
zkioxC4GqCVy/3SSsd48i/DtQqLSJL6CfRwlFjPFzcWT3QeZzYrIrr4+TRdg
754RYpbpjKroHkoC9rUT+vPppOlan1XwtycfQSy0dI1EihAbY1w24Se/0/gg
k+F+uUminHw9W7+2JkZ/AWM08UkfC9jZOnuQ8Lpy4+/3jdyAlhRnFNKodZhL
4zkKycA+Yj51UcyPAZGe8+CldQ37Jbl11XX9EJEmqV23ouvtrfvvqZxqGjjv
yH/Q3D8X79pFV4q0Kh4x8mQhvGdWEgO8qlMbka5Nd7G4F8XcfMDTm1PEvE0+
x216vizwa6RPj/ZTTtdkAaGPtfsnk9yTLw1Io0HPhzxoOfgpHv+ikNy0HtoN
oCMVUJsoP8vVdo7yim2pnCuWCsMlNAVm+j6lvBPPMb3ykZEONczQCv287pWH
LAt8NnystAitEoYBqQV5KN5C2d/JbfAfcb/idO3VKOWbtk7UY7fjZ8NoUG4j
P3odM+BV1Er4bHeReX4puTtgZo8/K1GVFUdxoEJiwysRxjBwtA9IuYkOVF/7
wa3rd99Jr8rcqK228duqBn6ZRBJMt7GOuoGuoHXH1XF+8lhph8a8U3jFYXFX
vV7Siuui+9iyS+EvEDebxU/u/4GVVz3vYj3tiGAzQ2dY3XHar2QuLDWFNBxp
xf607PQ6JoRVXTa7E6pyrfre1sDn5nB2XeJk3ybqYbQrrjQ+aphcfQzo1kKq
Jr6FF8cn85hw4nDS9QSng070GpuGLdMV6k63TNM+bn/rPxHOPni5b1pQcSKx
m1rFfnXKpTCWPeVj1ry6ABllIArNIXUq5XmOZxuaHNFSuIDUw177PvwOokh4
V8sfvlmfgbC7TzZaO9KN1CY/57S76ODbkUY6axKxeimaBmICfQHwY2HbhfFY
gIiOXgL5n1ncbo2iWDdaPjMJ+1okb1sOtNnBTEIo2j2oHrdaHyVTEklc91a1
Uq2IjiS2RpYcCgGamBqbpOrKFm70fjX7yoVGfz7rL++bZHV5ml8Qdsz8+LrS
a/FlZC7v6/trvrBeEu4uEzJl9ypCja88TvF2Dzj0bVXaBehxlUgtM5niQZkN
6/s9uagbaO7uFDfOmy2MQ81cDdK9CKbD0nU5kdLrcYOccSQPojONrLdR0PWx
o6cMf/QiwedUpR62AUiytCl+LcmNn6HK019Hu0kSg0sJ2VvxqzP6QeCCLaMP
TO0yK6xM8V05DLw4UaTDSkJD2N/uPwrvf73VBbOnzA51sIpBwN+/XOS0ld0P
E7sxc+vnv0WKZSauwUJEf8uDi0f5ze1WJ5D9k2GlmI3f8qXoLE9ORzTKzjYa
iFyGt3osQ0tG8sYCiQYgqd/E+zcg+McBgTCU8nYyu1yRPl84w5tN+Os63Uyc
0rksjQ3T6Jrl4iYBM/zfN8iPD4wL2fyOpHliLE86G4ZblRadRGzaRSCsGmak
/bcTptssSXjJotdeSFaVWJsoNwqJCKSuYsv6rfEWceKUIDCfJl5BpP0pUCaQ
+1pQWpmUpWw2/VTAH5LpCI97m8XLzgVQSGy3Xc3x8MPqIhcRSqpB5sYIsmbn
HBCOImO1WfkaMHTZEj63P/TVTdV5w1tT+ek+DE4/yGc339TAB5EOOhz68oo1
axIe8HnCEx5lZTE0aoOzyvsBAHL7K/Uqjt6IYnGpAuT8MfpKAz8VgeUeHPl3
ZhLNzwAFKSUookQO2lEtxD9BK2ie26YZnZ7TyVy3gZzYFE5dc4WG4SSm8WOd
sXZb2ZBC5ws6XXV8tc2Fu+1JMG5lSF0tpenOaG8gttfqZIlR9B+MNdYcPWr3
AkoU7xfiI7v5aHp5ccv9glkNn3n8YEyN5Y8vtmP1tJ3VvkhuVGTgITQoJ4YQ
HN3SReCYsYkFtterB+m1hN70r5QRFWUcsUFzT5MRkD3BXTF34aWv5H0HyIjw
VHqGYY6CcD3g5Ft0mWrI+2/qyXCWd8u/jCnJTiy2fkoooQTLMra+1jR1KekZ
uJEGXFcYnzTBT84KFYwp80gbxGINPP+NzIcJcDnJOz6fT64fgYsNfT2taxO4
NTyOekVf3XOxG5GaLVzMOPsZGP2siMymeg5am7p/pdHeVxlPNqC/4Ge7XeET
j8qGPtV33TMDVjBAzCi4P1hZAyJrqb09mSYMsFDrEpk18LK1pp7Mzo60wX10
SZXCzDfN3DxctYvH6KuhJ7TNy+XH48Hw3M/NY8CdzMpbTYGnY2DLswhdK47c
5ndQFtq7kkldWquhnp4Bk5cIBRseddpgEPLLhIbNiHAqjdYxDSw6Af7usvF1
Hdtz3uKEzmbau76eeaSAXk6wUUTm8in7QE2E2ZDfdu6pdHAqv4Hd0z6P+LMw
CVr+SIKejA0DGeGvjIOA45I4NFKKsqrZ9J19842bJAmecdQ8FRw99UyX87sT
JTSsBav0p7yH+ZuYlxMPxQW/Zcpy1X1LHL/sxurrBLmwbrofo8VnPhIrfPjs
cXIk1LNcfK04OFBFdNpilaQmV+GA8rUkyJ6iRckus5D8a2cY3QG7Fr6pqAUj
o6Pb9IYGytiqTxNj8x64ELkMxWVP5P8LIhfwoW2rkCE/DFUCC/Vyiev2xMQQ
IwCLGLAa0DtgpoMjjKsFn2Exi2ajOMp1d+S0LyZsm/nb+exWFi7M96ZgWIwZ
KcmJ0hqdU9YCYqzsvp316/BtzGl/yEl69Uy9KIJJi2JbnS9yw2Dsf8vTCw3c
TyEuZORplJfm6SbJo/IhSzTcIPmezB4k1OazNAf8TAwy59pWayeiQu7nrayt
3zTbL/C19wLsRFRNFSgGmvivvHToTAMefrvcOFvFJZQyHhUF2Y1FN1FYVxqm
ERZQ+75JMaTIv4eQ6leQx4Fv6x6swcn456vKkUp0K8P+ELXlcXbQjX5wjD+f
1oFy1PYyaVQ4Yoe8ew8O3Kv78wmDMPoUVIl6t5VPxSecglXJF8GWoRUhPzOc
YXS//wmJGVqiMyOG+YylVj8OPs81UIVE66aUl9qCILtPDLAM4jBz8eJqiQNH
VMdkidYMz0MNbui9ES1v1mdxT0Fsa/IKOBxap2/+HXspI669XKzHqNwuIFHj
jL/VVXdglwRB8QFxsToIJWkQpB37EizrfjrhcUEGqgdxF1nGhi9fKIsGna7S
CLBh1M7JZlfNZitVKqASpLr7e9vflu7xpBc4yNxAIQ/aVz6O9hgmeV+PpDJX
KsBw5ExvQKFPZvlrHx8wQUtup28izukX4WqHvn9i2unDDqOs3r34UgtUQOSl
OFhp7U8pmDEAHH9T8bAPYdRcpMCVT3OFMGA88H523d8Y0CDLuv2eW/Rx59ec
YKWp35E2YciPw745kNkV1Af5KSSWxJUQPAOANOM7jtI23EmjqWvxe3vxtUMS
/bV7kIPX2epT9/URAyU+lbNmfdxXMENYaiFSlegQ40xXWw+5CFH7obLe7gwd
u/CZtipXp7NQo3xYg/PEFKLUb7gYWhlklSLv3S5spMOwP4AgQ18MyHfdJA0f
J0bz0CwMGpa3YlfO/W9LzjDmhsHYcNKaQDM0u2zcqo5NiQrWaxcVXskGTB25
/ROLejAfgnP7geMq0Tff9w0BJcZ5I1M2upuEywMSJRSzZAWgO/tMpSLZ12u0
IK4NDcFg/W+fTE8gEdUzdYO03NXVAjaZKuJq/BkJvwBgm+OutR8kwW7QkGx+
OHgwijlGc9dIcKVzHYgFxXSbm4vcLJvN5ldZ5iWEYrqiknxZXAGRSTE3NOUH
MmjpJaubSe/YURdIrEWauU7OnbgD955JxJjaIGIOdG0ppEJkN5uRnMTvfQs4
3GCZa4bVZWNMqfJ8s7b/iFSQOMnyaNycLZ2sqOAlxiB9EfIkbgzhfWGMbJZD
VJaThJ9S8KREPXD4Cl2XhsDQ5UdtwlWx2uNitGeNYdrmbLjdr/bVJoXJPh0y
mISFayje0Yg99VIgdiVyQTdMsM/FVs6Gui5KkKC11yi1ZhaRKMLDaJFSO9bk
2g0bClHJo5mTFO3eBjlfTcmef3L5OksB0jmTtckg54UynQSlYZmxKi8ORMFO
UKkU2R9EPZRG6nhDuA+uY5o2DTIE//BJZdOOdI3ADkTQ3CMTOJOuzWJre4Jh
X8u6kXq3i2vDXxWABB1eu+/JaqznoUwUoxSS4ekQwQGvqtsmZQQuqyFvUefe
yXgfs3a5+yJu88FKHg9KZdfcoN+bLo1e+HxN/JG/5mzUpFYzmunXNGLCV28R
RPh1wDUeQH5zGW0AFoobLAHjdcRLFTKNfHJ1gS1UsrtZJ69tKnjbUhdneJwN
bvOn3sg50WaKaJgM1cO987RnduGImo94eYFrU4exyoWvgF0BU/+lWic1mYYN
vdHMzr2LtkDUzCWECVP9dSeZENuw0cPNMgwAjC1caKAjX6eripeB1m6h/wYt
exdZupc5muN5yk4n6DzNRMX7g3FHZ1mvSyESVtwe6ADoRn3JohyOW4Ibx/Ku
cN0W/YsfWXOqNtyxRVKow4JktZ5PIRHW+RFesdmY8crsqDMGR4WXTGxbKN4y
A93Qi4nbOJRCToVPOgGMr0gJXQ2fnghk3yEN5dmGA7q5jEoWDNtxxWKUNfcl
+LqIkzjhHkZ8NZvwG/vDSx0UPpldr1l+296OMFvYjlBN1qNpWBbUA3aEbLji
uFy76STekkYdFSKrjmfF7Ykq59JHm3boNLLSsVt4OJ1JUc1Co6+PRqYWzI31
2/kXq3+l4P22rhKQNNDYVSGsqs0fUo9JYI/sRsewzL5iFY5h6vFLpwl18Jlb
jBwNNR7SkaY8tkmK0wjVAe76MuL9IhnLuyEhIC8iGomwU8uGCPcrVrcWjSx0
vGS9n24e4SdQqM/S0Wq0anUy9LiE0dYEgynf65KyYmIRLhBiXuRzgNE25YkZ
CDFbDdVWM+WyuRChawCq7krTOYePnXr9ibNjAvKdNyNnV4hoeTR+l3nSr9Ic
bMzwBYCsUD8TVxdwVlCbciIqVW0OVHL3WLffIb4u8JZXLBXA5AqqMgS+n/lZ
nS0eGDaobJ3WSFEi1YOIndLR95IYEg1yGnkVNvgXg2wJ8KwaoA7qeNMrVLzZ
jYHihoLrJ8wgoFpfHbFXD8irz2p/LL3JC+DUL0zf57+k+AXjC87xuuqwH7A5
9e+RPyqKRguYaZFGUH86D501qOsGvcGfZsI7HnIaQ/4B+2xZ1PDPLAawDTH7
fpk8nJVZKOe92CVF0KBf7p7gWlLWEqOU+kjclK9LX1jp0kXHHGF2V9aMeA3C
tX3hVTfAuROhMl7xZ55bczFMOrDgtJqMMP9jdveVWXBa4KzdVohzm+kmn7w0
cXTZ+dWc+WGJsxoHvFLzFjFhdtqiSV2MaID8UDaLtCyYC2baYu041O57d0WZ
MoSjq02LhkH+P0+IgnD1XU5khEC2uWuA/UgWwQSnVaPxGYDGwm4PIYWFFYp1
xDP2f8EFrbKihzGtYX5egTDGOoclsSR4CKEgj0Xwb1wzttnZ6coUR5lE5lD7
ENdPZ0nTFJ8Aj4hCjT9Ta+mZSS1VXXyLUSY8B6dpp3xeDJiqpLGQnUN+XPiW
Dkb6KvhTgJ7f+GlU5VbOPAB5URq+v+ya0O2mza9c+SXxaPkMi8PnF5JzZXri
R7k7ceV/UK+pmsZWnU7FclwWTnioVnsIg8vddV5ppjIH76KdTMk0kVjenYvl
dfywfxyY49kGEitET7HXtD4EaIIdjE32UL1TZxEyhCGQaeLgba0rrF78gXPg
s1DeugK3fIB64WG+zIQP8RPK6xcFKMjFhouhOkCdf718t5BDsEMbavjyD4cY
KXjP3ix+3hjJt7QZe8GMT113WNcODK7+92m5jKJOW1LFImxNOMm+3pZQVZOd
YX+ptI/1NK8g/S8SJquRbUSCw0k5DV30yQvMe/8hy9nivDZVJUDtq/LSe+aL
DjHhBcZYXzbtBTO5+V7TCEX/Ut0gGoL2g2lj5XxZT12f866r4JuH7bqPW+yc
7H8uoLHpX8jUfOG6ePCaeE/wgz4XyEUtFaLZEikk5wzYzw5pt79gWlTf6s2W
sAwRmBdBoiW4nhsdffocmf6AQUMyvk/1z7arc0Y1GDuWTjwPy+/CaAV/iF39
jXi7cDMe99MeTfzdsLT0p6z7WjoLxWo9qaZ9/lv7PxXOjJI1A6FYXBcwRRGB
Meo2fN4GUlAlMESdKvQzAkkBcOw2oMM5llHW2jqwNXnU30IOhGmKl4992Kpz
6YwEgsiscQ1aXdQDuYczuqtrlhHU+bio+6wlKXf2rUktagk7TfZW+Xxo/eXI
4SeJmHmDLmkNfba5zDSsqsMhOiMMFqDU9kUFMNGWOCDynRY7dYQrUsxfR6F3
eH2ud5f/BozuGhqjO6sZtlp3EXgmgfG0kTLm24UuWUNV63CIn+W2CtyYLdMk
Vq8iLM6Am9cLCdq/vNrN21PMZa2WnOOiG7kRLfNuvTeYQ5qmtxvrTnRUkn2n
dFYQmeGM2yWFEQVIthS8ZgYWOmLmwwLhCn+NBXrakSgqxjxW8yy9dPFfluxf
riVLp17pboFwqh8M3Nl4ZQcwihuGxHogVzVQjZ8HXn1hvnno84ffp3c9zqPS
QkvW9tOlYvQDKsenkO1vonXWfU4h53OGmm6G+Tgr7Ne+FdlP0flPpBCXWWla
loKdH0Y2Zjrl3k/e8ppLdWb8pagaaOys0hnCCobAW5asnA7G4WkL2xbEeeqW
zn9YCs525a+/LQFQp3BVh3L4y9tXg6qPoxbtUUUlMNQlA4IWLK83PWEit8nR
nSnJp4hD2EKqE5H9TpyWJ0j/98HRZy7goj0TuYYattsRSFnNG2SqraD11wFO
Fr2aD6yc4C82B6X3TvNbLS8qi6f3xDarWu/Q4UiLkQeLOgbAo4DJ31Gi9O9a
DlYn8dF0qgmkwQ/ZJnMjkNirdnMBqKVyu1rjvWgSpdFuCdJYYP9FN7gaGOeh
nMViEJY2eI9lFd/PCsCjBwECusgOpxO+7QWuFEzorFIqW769DPcGNZdn8l+z
kJY65YiO0gZ/aVZEBVnLAPK9GyOjnKsN0kzWYPvHyIp8MsBZOo0WtgjBlgab
7mN9kpurGlUUxm+ZS2jGIw5VwdHbX6T341T6fRQsaLOfakJ0hisuoJ/owhNu
gt/QwW2/zrrJ9aEXfZPPhF3d0ndZ4bcXRMGVkJCMZlRjCWI48Minf7R7jLIQ
uUza0oWuBeS0gDLBMt2VZpwT+LzOg3usxdvy80Ke+75tyUt693tcEvcR51XF
RoAegKUpFIM9Wabf3oA5gBUHabCmcOSPAa5HD657NKVL/1yZrBiiv1m5BbL1
PdgB5mKQdAIHLTadEisDhKFp6xSvESwj6KtV8BbtuSKYh4wqFVQXhv12CUYp
HKvuTtMigs8jpjEqyc6Zcrw8+VlepgkT7LnZhjKt01/latgpNG66L2h+jdZf
4pPFaazI+7dsc3/TZ7TuIBviLgBnp+FbV0T7imbpJPBr5V+XUpGMbFIpse+v
NMXKouAMEzFUe179JJKq2SHhyePx+REc0f+OzTba9jzNB4WMCqfSVe8Rz/hq
PoYOVj1+RHxK4h49rtpGwovoQVyho3vcClE8baFLUdPNhLjYf8KVe2ofZEec
nkXZmAMqDFWrz1fdM6q/W7W9aKg+iNRvOSd48CdySgkvn9+EXgKMzFpseLkT
VO9JrvXwVX0Pl81bqof1MwPZ5+/XiYsIn8HD2jzQ9vm+Chqloy8dthJe7C6v
H9rGtr2LrW3d0n3En9AEVyvYm6XhlmNVM42t6ohS6xEnpPpFoKU5Xrsu4Evh
QcddKBZ4JO99BYP9t9AJzTKCOSvTj6Rgb8clrGp1XJ6grRqxdP7YGfMti6cN
FSNCzESQwokvXKBiSFPREFDlpn3Xv7S1N1mEgOp4Uv+/WxWpgsiSfD4+VE+7
7Hl92xJAPFZy9wH19IWJsUfQweIvXYnGfYA9igezf6vPtPL+abddExYP3V3r
OFW7PEMoiBhoH/NgQD5eWW4AChhV9ouzaHLDEujwaNQA3Qj23yYIoC0tMqZr
/U/uiyE5IWk1zH0JWqISAApJlWNjCyI1H1TkTiFJv4+WBWEX3dbTl6fJtqqE
9Grji9nWJDNikXI7yld4vC3uL3VaQquySQluxhYCZZmho7I0N6v3k/GmgfAN
K3kSPqa92OITGq31wAKg9Mlib00oCSP9m+uo/slp9q8inhFf6ZXuc8D3jS7G
ehI/Cw/SE2RdrflMQbd+SAU0M9ZC3+2p6qSsYCatK7nXD7QYUyEkzLJ0vemM
mWHWEGOOI34kqvUzJtpIQMXexnk3zzLUOAxtZ5Np2wIVeXyCovuPq4crtVU8
OE/r/eRL4egD8dD0FfOcPx/wH64Sn4EiJ6Ax+0BhdXBzjnN/uh7HeDqh3YDS
cx4uXHwSV21fXZKsqVkzvukQegdF5aa+hqMKWiK8pNz+12YgUCI7WOa4Oj9u
TzEDzu2ochtor3zSRLgosSRkcZpQCKsEUyMjqPQoEZZpLRqySCcRjZWUdT+P
ijWGA8YJ893CVBDj4ncU7gTiPMcPZipicDCG/X+Lu0aN9VEbB9/el/BAcn3p
Rb+MRQ5MYB+0fcJx4YIzrDZ/KkL7DUv2UjtsgxSNMe9kurc+9NgR7yigDRM7
e/3co8FPVbVhkAeGvxBo/EBoKr59Zr0Rsvzzg2J1Cyz1rGL68I4Bd6jZwsMO
ZJJmarZQZgzxNbJnHr7zFseByCh2EzpkilZWr8/iSCwvS0yQMngGAJZta170
RpO5nKWBLLUfsrRX79nlABJAe18XdSzE3YU1ub3mjl3puc0Bei5mfhfoxZjo
1mIOhjDkGcUy0CcITVDRZDKftbg2MXrRU40oMPoOLIORGe1riYOVBE8bQQmS
/wd9n/0hyidQwJepJKXWJ9pSpx02X4ca2zfwoS0rbhthb3aRyEzxjPWOYfh9
UHMjS42QbKlunrd+lKYo53CtywP4QaOEcqJcj996YgmbBrQhg9ODgE5dowJE
RcKpSwvEcJqngy4jnunBL/fUPmMWYTv52gish3oNFFc5O6bCoEGwJHF0HrmR
43ahDDKnlz6MfMqtUyQOYCHdJ2lod9mGw5mxz4PlTrFew9E2HT5z3xhYSnRn
pOvRQx50NFNi3KeO0obkkLGCLejE0BuumQcW3jc+9z8vS8co3APwq9BOfrU7
M1TsMiH/f+jI647iZ8x/q/uUTezmDoL7Gw6k572Oh4wBkGcuFQuAyqLNqY+6
1CQ3v8vzGf2I7W8iTBM3HEdBYrec6QTwQNEhS4TRa8y/or6jhV6w88XWsGvo
8uLdrsTxgpOPt+cRYMj4St7kOfJSW+zubuXOYd4UM1EFrQ0/pq3tAyeh6pyz
O1GcwecNDxDxFExlCooDvsS+6OsRywNEon7xucCzuhiW+E2loBCZ6ckQp/6H
riu7tuQe66oT/NysHqAYbtlnOEwJDuywGEO55Vmj6yPPfuei49DCbN2gkjjx
SoNRFc4Tn6VU/bbgQWFlQ2PXuNcI5nuS4Rr8+f2c2XZ0Mu9xXgLLC+/GryXS
GjUf0QIj+GcuRtqi55OViUsS3Nvu170Z8qInHkAwvjMhd2B0YxgQT8MdiWOJ
PDaW6FQADUEs5rEf8wMmGj2AVOQKuaEytN5b64yO8SjGK3/RnO1uJE6eCYeM
fEqEiXP/mIM6ZcoR4wrelb0+rFmfstNVTozAATEP7WlquZHuX8rmQyQD2aKE
UEhjaPEmZHmEdpQn4ZOIza8pG3r4rbsKz7kKXoKrFYve6bCQjal7K3U+ZnOJ
TSenUlP04+mhuRxE+ULgrDjtYdVSC+/WafUyT+dQAeOnBu5g0x/QsXm2jdJ8
lv3zfVk0erX9ZxbLKDyPngZ2Sj9xrE+zSvrpoAiL3ObNnOX3z9xsYwhAfu4Y
BnlzRe366bCz3N0LpLH99ojrFkNtYGWK+5yS5raNExXq4gMcom56SUMRm5rW
ZgIGC8y2PatL2RzejBMdzG6vMGCMIz4vmhR6KesOTt7cWRGTHeml4Y0J0Xx/
oWKa3hNekFWlVi18ZH4pBd2HzkdFPSkFn6yjohoxOPLb5PH2OwTR6OtIpTAS
AETvOZVt2IHXCH25yyzUj8S7q8Zoxw2mEVRFaplGl5BH1rZ9OH7MN/t8/OYt
cePZokvmD6TU4ukvLGEOCtksrvpkC+aJjNf+VdwoT2l6BEfdsS2jJJYhyHgX
aRAdR8aymeYVdhXaQVUcD6/2P9gaUkMD/A+8IKgCyennwBsCGpeA4u5CbxvU
IpiHbljckR0XmcC3AnvaPotGi8F3h2xa/yX19QzKoDY00GeSL7IpSTII9jNR
j0dQB48oI3FvyjPJz3k+Rsmiy8jZ23fO4LA77BXIVD/irQ9+i+vU90pnxKim
Z0ete90D3xmW0bKOBV3K70wwB19gU4UPGbom/61rICfun07gC/TxxqJmbSDV
Y8RBuaGE6YJ9DGPqFkbMM1hR7T3sIkTv6IoErF0O974V00rDr3VA5OcoV4i8
GBOEBR8xEUMVEkEvYMKgbeM8MFXFMUG7yrZ6biqOwXQJPG/+xPYhOUxqXyDM
gh/z7ybMObdtjk5eGTY/qMq5FdFvcQIsIz2dEY/cZqCM7PJzreU6EfJvbCKE
+j8ParMTv+rF9+4mZwwCM5qhLzIjdIYtNJkP32FoRr+E53wOpqtyxQVoEsRo
NiJdKi9HOdpCnh5IH8xcr+BchlNPUwU6xD5Y5UcO+EdDOfcKqVcOQ0l2ZZER
E8ZX073GlDJIuxjBJvrXRYy0byMXgcVJ2keaqwYG98HABQF0jg6uvws9NI0U
2X18bCpLj+MpEqpp5dk6LsY8V9/V8zcMpGMRyoDNUino+25PAclXy4TcC1si
fpMTdo1EkDAipor2s3Yi4OIJ+ozbZRJVR1xsRYO6i8BUPkSzDLfQlcKWBk4P
dppeKRbYJSULk3LXKzaTlqNg5Yp1b63yjmoxXEbr8a71WGcjPKJlql7HVGdq
afqWFlmnAQ9OnIZHiaKex+ojiAQTht8SoLpT5SC/eFLSE9dCRB6Bv/yLI4sn
kC22GEXwZhCcoJTDHGq/0RJNzbjzSmNk6CvoBFVh2a7kL8TWFJ0JoWwj2MRT
WwwqJlFpIGiCRjaP49pvl1MD4O595jY8uea0ivSIJgpTClLyMq7L5c2gXcyO
h2p9HJkMift15YSnZlHN/rX8LQvvTi4y8Co1ry470Gk8IXCdnEmp2CCMW3vi
0vloE2+08yCWf3bCZ3E/X3RS4RTrVfdmruF64scISr98NVoBydVv7FtfHZZ0
KX+PZSPbdohc80X1sTI4aiCMYm1Bi81o8GEd8ddX2tkTsKRwki0FQtT6oK4o
0z/8yV2G64CqDR/gl+WTOtp1yqd/4GtNDWuKVD0/eYCzPE6hZQAE+uf9rIiQ
fXX4iSIE3gbIf1PEMggg14Jzz1Ogb7ldktgIVZSPeX03GjD0747RsbEgYEDg
fAkoQjx7SgYm97aEZPajvia6B2D7S+7Nd8RqWNH9z+8PjrdMdcLMWQGXI1Lb
/rn5kK54fwRCAPBcHq+xc+4Ik6ECMe1yByq9cCgmL4ZJMSWT30aHor0NlZLe
sUqvEsrREln37Rivx99ByBzv0L1qr+NiLZn/sr0eb5NCkVh6FmMJpd98cUbd
J6b0Xrd35JqkARNFX+kxgx1AWfIPC2MXdrcfTF19A+rysKLHLTU1RZ5yNcTK
JzQmFTfb9DAoZz3c54joupZGNXjV2q3I5VG8zH6ZSF54/VJgyFubSt+oMIIz
KRU/5lj8mONyMdMG9L7u7cC655Fhttm5dqUXhsHOq/BoVXQmFMVJzgZCzlim
fgFZXU/BiFp9CpFCBFGN5UIy83V1v1RyI9uI0SEOJf05tyU9Bkz/vl14wPL6
d5DPjUgmCuYPs86AoHRkDABIwukNMmKkWDOrrhZp1gFPJKwyDLH7R01h637B
tiEX/VpjWbkDuVZUv3zGbqS0YG0J0mx8Cue3kZLK/jyvVjo3414pP6ehlREV
OYCiK2XHyAwFoHkEvM6CHsrJB0X8NGzMr6n2D9Ubbx18zi+nkWu4SSeuT6y1
Pdh4apFMfzsV2Oprhs8e4Ko6UAgw726bmkXyBSUkfoInhtVH/lswEdKfBUu1
/Tml7OezKwmjZZYh3Vihk3SodGODzBQc7xg1B3p8E84Kuz18PvMqvxRgEnHH
kSinvSTAbQA9MpVbF/J2Z1J44blmBgHzehMBEEyO2Z3r40NejLlpYWDNtEzg
+J2tENAS3ITxbstbnvbKKprcbhqP3HbhimBsnbQAzZJKPzeRgvcyfTNwaMMl
0fbEO2QLZocEz0LdgwN9wpXHdpGsU8lDkejypfDSWBG0BUIgcYJpu4CZz8wi
PyVPNT4j+AbtB0eOVm07Bfs30fyndBg79mgYDZUklumNu8jTNWsIJNjb4SZA
R3Oq/lmyGreKFtZPG73ssGJbgoHcijNyoG0digUpIiw1zZsnIEC/IIGsvxGG
tcoeGqi626xQM8WIz6ZRfjL/QxcgA7ALXfWfm+K+M1w9RwVIo+dsBfjux7PI
P+XgmnO4FGHZX4mF+Q9udvTmJ44dT9EuENttlVDr80oLYuSgsKMOCy//gjVP
AQD0MAINxz1/3JY8tvxlZlMYUDn8l6oo1l8HBdK1cDLJ58pyaAeFemA1/zzO
1LEePQOBHDNGZkDmOv2DkG1LLD4/P8+h131sJYoiP3ceFL1C/JaEe2nlqWvn
pHtsuIo88yEB+4ctSP3pdBhmMaXkoX7y5nMq0JtalYHXqGucoVLE1ajtOnW1
er9YhXD1mD7S2MxrMjHkJD4+TNuwEPrPop8BQUxoEbuKgLfiYasjIkXcUQZT
32Sj1QMffYf9Bmw2ybrclob/s0L+CBbCQCbWaADfKH5cL4s2q/vdhJxjvxWp
AfBM7xqpWQx+/zOhU4RFWnE2gnhleeEZou8N3W16mhdJciCY8W2UgDkUIqfW
/9DB/lhcA8/2UY3IE9g8VndWHP6UXlUEBbYaPwq+SGmicVgvqvb+nraEXFIr
tWokvwK0ipLNfClfW4lgyNhqkjunbJeabohssfKcZk24PLb1t4TpdG6UTigE
8CAWq0c5wsDmTJ5T5y5KUe0eHInadhCmtA2PzOpBSkS8dWwQXvBMcE14QyfW
Sj30e0REaRaWOutahtfa6Tptjm/5xvryYdsmoRwfKgMklKY20SS7nyeBfVqo
uZSgIywbaIVuTa4VQeregNb4A1x+QKMOy/c0i0LOZ6B2P3gTg9OknhLmqxQb
0bB2HtATQMMdGQLBk8mnTbeR9bVcOwZXOL+NZzpZ2skdKFlu3zB68b2ZbPKm
bVPHAvFPHc6OZDNmVCze/VAtI42hi/oYmEqwuqbby4Z2hT7mlEzGyx1/P+HX
QrkyjeYVm3mFFexlH+XE2V8uFfA+wrrBNsZGaBoayjz1r0cTR5lQTTqxPlFV
jZbaVBsjQTYSR8A9flwKn1s8kwo3hED1+xXBjUGhtwmcdhxZpmFNTBmVkTvk
i1LtOJOcoYT4x596/eAQp+BwFd1d688E3jMLKZH9k6lNyZ1tE8jB6L3HvOm2
PpnkRe6zi1xnaHrFRMAZ7gyMbvORWhcLmAAoVc4zyHwGGUVZeN1zfOYuW3ZI
yIOhbFEN8g0a2Ag86rEI+/BBFFXMft5IE1PTLwpk7tirQ3OM+BOfguQofbHU
jMsBpwkChcVNG+AGemXk2gVlRhwLLDMwB+i68MTCKqaQD84sW/hiS0NgkjDW
ST9/OdsR74jHlwGJJx2ryVUY8vWhfJWGjgkTj62sgQD7qcCekdiEiDplHvAN
ThDjFUyUkrphtqCExeikWUCPwOrpzGIWOLeEpOeAe/c5l3DTExiv7zrejGAK
O8QZWuAsvuXQhbW1D6i4hgcGrSpRckd8IFn5VBUprH+djVAkZVRFaMjB5/E1
aYCpIw3W7EqtEnqg0GCweXApqDVSmtdGy4HklBqewET1PDiEu0dIxlcivL9H
zdAFMI6AuU7JQinNM0rlNZK62+1eY5vYPo/X+diZq81cMJhCuE8NLTyV3I97
MBGolYdI3VvfUb+3ovz5fTsbVpGPfzD7DghosiIXs5VyQVDnbnWLeYDl7kna
ZfCqqCr/ODquwWKbU7mVj1rm20yBlJ6mcYsFAaOIaXkVpXk71lr+rWqogSjV
sFBomJjRbGULU/Y8MHdg02PbjMgs7v+KlRdvyaPgKQ2DoUwMMncguJS6y8B3
oX7GrGKnMI2A/mC3D4YlelUdJrDUb1rBQgzWrN3XarwthurdboKzLW8rAdr8
Zgjt2NBYdGK/bdXnhB1xvgtrOQ326omleILq4ya3+JSA3u3G0vmUz/vYXTNe
7Aq+kCEy7eFz6cM45oRG/IuTdHvtWsE/SWJ0bMG4wM6bKJBZuxHiwiJMltbv
xXnHUm+bI12YaGG9KDLt7mmQkIYsRSgNQB3CsbNO31TRnCTO0HHXN731Hqbs
1JvEa9cOkN5XqoG7bVYjXEC1tWnzl52mRNbQqiJOG315d0eVy++/6D2J5sDn
hIvGhsbQMaZR921PNoxWINcznr5YXd/z/Wp1i9G90/uaVcDUWDXIAzk4172j
wS+o1YP0BSgWkQtT+VnQuHbFFBQi+2qdjFt/AKvbelQ46NIqOOUghZE6ithB
zLxVoOtwNSbpZ1NNaM72APlLk3DCt4qyDcdKjPwxSfzXrr0HH1gdCq3cKjHP
b/eKXOi3WCUio14h8g3NAwgtSd7JDkzOc/R48tlTXr9celFP/QI7i9+cfJl5
AnsTErPP68tbDrI4wJWgYFAUy0UeNL4DFPhDYIo51KZyiweeSQK/WNJVTFUP
wbK/B5XK5DETwNykE/tLwaQKxtEWuSRJA8xWuf24JFdMLF6/CId2HJTilUWz
NggJATMg+r+dkkbfOlyoxhZgwhU+l4idwaGn0wFNaQCHKDZzm/KF9e+x2RwS
jEIlde3nXJ8zqW/nMnTmT4UZG9a9/cS3iDLzXPkxTSptNEHrDqsKWVxu/FLH
WUDw857W2YU7rHW6UKTIkfPi3gm6rHHqryjhocsVzdf20PIHnPC4OMOYrU44
1+6EAQE0B1OiIpuqWQjP/c5Atmsf5alzIQiZ9bgvQXSp5eiwDHwtkL8Dqi7q
ewnr9KqOqJeLfuADkjV43PFp65u5jvrZwhQq+UgEt7hoU4RhyHygWnRucOAS
T/DjIrzCM8AnhKkwTjo4AsmDoDjjWDS4YJdnxMGTXi7fyy2ma9zQCUveqKTs
iRYUxgIBvMromS/cL3NcdhUgmU9G8cA4XeKZktbAuIpN6W5SLHJ4xUtfY+zC
L7Ht+FCoPbkGUn/ploX2z/36hh/iy61ipzSro7v6YLjf8RxA6nesXz0c7Ufw
odSNBw5+aS6mnmqECcy+V0IwCJPvpLW3mdfRvuED4CnEGo6faktGR2QMZ/Sl
4BvQ17G0xf3VaGgINhvoyCUhPwHjOhDKxJIpg6SWxNBYxoLRDXe3fbL9xE1W
o7U8llCQfRYP0UxE4blQSvcBtNre8I6htKBzxuOJPTFcB66FnXGS7K2pSUiO
S0K6BmP8FpVvBjKSbp/C/NowFT87fSo/NgOW9tltBfzne8d/RE7Zdri4zhTo
saZZ7glwAICCWW+0HrJCLCpLbGRTPVtafhLnD+Y+gXptNESTME9oZ3m7pxWA
MbnisNN/EX7xsGci9h9rykMglSTRI9+Lolm1+CxnJHfFYohGNhj2TcgszfA/
rKvtZ/30EYmy/pzihI9ypiMDSml0B1Ci6+kAoZEc87syOwlYYBjNoyYJQNls
qHFacGvGsA29gomw/Y9KpkTTh9xDfRVa8i2IEs0qCjwc1J29Tne4FDHCpktz
EULToPNHCgCK2ldlEtkqD20OEVJ8Y1ByLua1j6gelX6NDF1R7pYJeg0IM/Xn
FAZSZ2yxuaB2Uk5jAWl/KuUTFkfzy8kPbbXCdeeUM4O5iL8/5s08lfr/aLmr
u9n+abe4rAjHqIVcW5UQTwEMMcVu4+C+SR+2OouU3sxtp3poGiQHps/aOAiv
AsF+4QoK86Idm9fliB7v83fpjv/l91K3hGET/nNurOGYjD7plbkrH2DJ5J28
pu1WmtLaIPdgZvwC9k+uALbvtug+IILwJCJmKOn+AkByqHZjE1ysrLBv4WaU
9YRO8tz3qzhbRptb+X3GLlrFdJx2hGFx1d5OkDxp80mdhyJeXnawLCyI7rxR
As55Sc+QgizVAWpT/aOleBwAAL0+ncM6pDn8QgeLJ2MUODNVcdppKc7/qEuQ
IAf6ALcQR4uMt7vTxUGKgMWIdXf3ZH9XUkwrfJLNE5a85dzssNzdXz1QKKnv
CGlgYrLiu9cZqHo5txTKPA80H+Zs8JXANICNRsSMzWlQYWH9uvGq2pS+LGuv
w1Apl76LR/mIlbTemByPSc51RrFchCwcyEL1Hi9zQ4frRe89AUgpGCv181e/
BJtHOPn8hpro6bwEOS9KbTin1OFkKAWh3x4xOw8ml5OjrDUdGxDGg5j+ufcA
zwiU5+Tym6pJ/9IADPiiZ2g1AZ1Z/fbcjhyJsTupxDU7kDN72CgQH9+JQ046
ANfKLPAqeGsoFKWrFLt5y28euaVOp0yvijTdpZ2gGmzTqnD2YPtjVZXjAT/P
IX0DQ1Lml8beyIiI+txh6IYaNMVNDxCC1JTtK9i7/fEHDpRClWNoPhXxyor4
Z3h9szt0wDM83mOU6rJjxto6xKuFxRonvKJhE4zw2QPo7hxYzOl7v7t1n/ul
2ZzVXQv9+vFG5ciNKCvZYA04vrLjS3sZuYot7v5Yu6K7RlUqanUWhobLsm5+
4W7SL811gdqlNQ9L0Z3m6V8/4SEyXML3eNLgELYEdKufnQWuGOA1nuMwZzT8
aQ8N8gL6mcfp46TwF9JUeAMiX74H3G7OuJCImtxZQXXdZfuF7vuCSKw670sG
A6w4t63ltfTB5REZfIJnDG/uK4THYWeDODn3jTMqg8HmYmQdTsvKjaGbczLa
lyMFd1olbtTPQW0ud08adnp1w/qETqdD2Hxtspoq7exfKDSQnOe4b7+EDx3W
xgUuMiwfra/T3mvwqNhjWmxhHySIhImxRD2pky1KCN0dHjeopOGErxsf1JV4
3ZPU+7Q+Q4GJQLEBof/gsS6DM1x/0eiV9sPhMTaFvVkBficAQLDFZcnZDd2p
lyPbjaTiB8datn02dADJG+28qHoUhAHjui49CCCCjE6ppWnWwNAuwekogHc7
I6Urb7YSYyp6ngSHtUKMdIytSYZPHGydEmh3r5lV/wBxC1/UnDUwvx48ACRc
a1c+vdf0sS4MJJNbmz/KjPjxmwfppxkNdt/U7IymNx5s5GIgXLYSjMkmZ/8v
jYNzZ3Mlvt18RW85uBHzY7/h1SYzg/zSm1memSje6bMhfTstax6GOrAjW4JD
W/mkMiNkTT6NnE1GRzAustA59liwa5koFhiMNYXJCyZfrseGK6dB++gx+268
3DMr7ZocqM5BXOh6k68Funq6UiuFxOcQGsvLa+yhkAmuw0j/q3oaEIm89LXJ
uULM32NBWY3qxQsoQXLSlwBUoOr8CKsM5oW7wKOxPVddjOarT3A6ESv/C+dD
BorimeDIogzR/uD5wxdGWvjFnVMZCNXOUqG0hEwKkLeNZAwGHGeLCAuXRCU8
Xt/pp3hTF/Bkzb/VwJwNtF4cjKoValxz76jvBWr3hxr0LSLpoU3wr6N30+Xi
jDFP3GAF6ui0ro7IZJjCmW2zJysgdlKENCQbSasodlknbgll029PcU+WKklX
T1lcZrT6d2pmJ50PiBmjFJlP0ynp0IRVX+A916L3+pWqBootRfZXJLQghhKt
24wYe6i68OswvwiFvlXK5ZUzaegmm5mv5Gu8mDCpNaGy4oqNgJ9oRMvIWdsZ
zotLO+Q3GHWKXoz3Uz0dy8EZVsY0+7HImvArFBM4z3odD19WH97lHHZymPz+
AvQ9o1Uup2sirjcPfzTqFHcZEbRuOzeSwhYgZ9YgPT7tSSkOMqpCWg8bXZBh
0Sm3Jnpp6vR5kQ2niVSG+AKQzn4CwWbBY8rbI0CtGp95xwVD1p91K9k8Q75h
akCMOs74T/gbmtI6NR+lkZH5TaqPfcZHE1I+GnP3d4JYjsrc/CZLapv0Y8A4
Almq+ymMyjf72oO2SzldRoCKRU7XX03O+jHWwdQV9EjH/tpTkxFUcRLQ8M8G
2euvRaOQVFTCNbxB8t3VPcIp4bU7Gil01nCUQOvmhz4DrlBZEpG9vJ0EtA2X
Y/yoJR2e5ddeNKZU9NnrN0D+22JmTYoeU1LNLD3If+i2bdu5zTciiRMsZQNA
rNhvc30eguQpDOvHJ8rEaDijRiMRPrgKPSlowEShfs/LWiIVUSckg69hR5iq
UOuUVJN1V6rkrzoCACZQpz+vYm5J1SUYAhH2UoibBi9pmzhLQ9JEuLsinH3b
Ht1cxzcStsgP0GJ6kkJyffaYCZG+eoxGhCRA8b6nhN0ssbnEs1k67k0nJ7dw
Pzk8CpEARP5F4Je5+aTnEtMxvx8ZcPExuZwrmiDB4O8Qaa/1A6UbiYk1hb2z
2qi5ROef5R01gkWelYg5PqzExv9xaVv687pX+0cU5FpL29FijMVB0cO8qE83
XKfU1uPvgvcMdildOrjSNgQ4HQcCi1lvTVYtzSMkhk1GhX0iXvUavERi182t
tvevSgWcfsQitAi/XWOUWi/SaHd+OSezJo1l0AnG7XZu7zAbwtZ/yIiIRiKO
uEY6RgCpqQ00Q928j7zEApjpHcHMisNB7LJGeNX3Rq5RbsPRX4bmvZOvm+SU
rDnofJqX3bqmU7+Oz5qDBPlj7S4F27CpfPO1AkZF9ok3XIGXPqpzkE2Wdi61
Mk+33knXWx96KtB2c8rtIwvhEPiMNVZ/G4CZ872wonwDyhjZX+zHxt4GPiPF
9OyLmJ2CGgX76AkKampyee+MqHuKBp5q5hkPEkQ2lWH32wu4rwATbBuFg/a4
JDcMmFh0i9g2Q8VVRYk8dYoH9CEkgmQXS5V68GnAkqwlnnMohHY1fgzgGI1q
49DzNnKp7cEz25aFG4zzjdk+MBS6qTMX5NSfu0FYbJ3t/9oL3y377GuJA7nD
5A3FK0X1BZblMs90wNIaOtx1/BVwuY0DTI4R4hwn5FeYCVyfQy7kyjZa6Mr0
smrSlFV8Q9mP4IfQCB9FGUIM+cQB7DeaQfWd4+/QMJJ5J/m6ktCEpdCQWMsY
hl9flSNGx9WOetUT2gaECTdYcZUsKTHAPiJHDC4xhESGRYYyCQc8uPWGzGEr
Fw3Dn1HMF0/Opa08R0dR9r5vbbjnr10F2dCSJhl2mYVqWOxi4SKQJFQKtOBo
12V8AN7aJUPIJIBmZk6ljuw0UiB5PvO60eErOG536utbOEDPHbhLQYloRn75
PvgGXktMZBVy4d4zKiM9PB/qfX1DmRu/lbGrbEwRXb6jLmO6OYxnsx2vfsZd
ldcdlfXySyVmqXZJ1Uli5M2ghNGbcAQlmLMhO8p+QT8Gj4fG5P+GIkbAxeSx
QNHkPlWjT2mZm65z+1tF/GpKbAY62k839pdVhMs67nigVc/c04YqHk4SBa80
hsBx5vNnFvENs2gNSTp4He2o2Hy2/1HF21Yh7XVVIMKs0lwPPKHAyi3T0XHC
FGSzeHOkhZmrXwSU+7ccm3aVYwadC6Uw05j67wyImuHodJ438ASVaeyum//g
3iAd1PpBAnLmKdtV2kN2bpVqDD+2euvWrL3Y1nTxOK4EVlwZbzr6yjGtczL4
eWGW0B9gmHKrBiB1AOxsqvCfKOsURPE+XGMh0aX0dh8BDbu+SS9XeB3eejGl
zH+lj4Vu7D9gCdjHEKR9F37UKMYgsSX5E74t7CxIOpMrnR/FjiMFIOxwL8qz
/1hsgmzyE+spNvI1zzjk8Yf6tMKjN7JrmycAEQFAqwBkFh1wly7eMN6RNg7v
ZxDYlGDsDq4jJuMRYZy0t0y3OLdmB1CYmnwf9i+cUlTtMt+TBvQ4Q9Db5Mo5
7s96h3uGZABup7ZLzvKoTq8Yo8FG3mHYDv/C++MH+a21XlbPKvB+3ia34uxV
Vimwhl9SaGyruQiMf53qRcOlhEgNlAsfq6d9prBajCcQFvZq0CwsjVfZMTms
PsIOi4MqZeLuxGQX02QtxerMgX8SsnOYLCkVAbmleECjlUrmho70vVIwm8m1
rUv7aqkcnX4i2xqyht2xoUs8I5wVb1twg0aRqOvIBQjO+WazfXcl/ukFjLe/
/tjPpaLPrT5OU1yuy/bBnkxgl86ERC5sMdJW5z/1CHxAqdqUMwIbQK+Bue/B
IC5h2b/deMkwp9rPwo4XeWVEQEVn9sQUxi4cklWnKtF+C2v2uuwRIuxLv1mi
HikRB9Ok7vmpviafCYAlhIQyFhxa0bBr/38zx59O2fp79hV7zGsqg0/9RGRo
lMFC4N0GCph71DyZPWt5OHMaxf9+Z4Xpr/gvfDfjVqKkKBrB4q2d/T7+kC+E
UQHWVleCm/kAz3+l2bKVMNUQKbI91tu7LJncLr+XWg3pVxtOcn2kw3GFzDNE
F9sMJmTOUtmgfXOGS9hVMQuGAiCgPiL7M98nIw+xXVzVN0NOfY5SpkU8hngA
Ue/Hm4S7vzNgm9XYTETo4qSBeC9p6Rv2Y9oLq1uzFaBQZhEg6CG5t68AvZqH
JWsrMaKiFkfWbc9amerdJBxjNiOgwGhhQVZgLfjp/+3zRBX2Cv9YQizRDpYK
42AZw87/bnvnCLI9gs1RPo244WOf/5MP5LmmSwRslXOunnPWw7yDJXl3fa5a
zWSGodA5rjhZkH4U6zbTPfo2+voFXLHy1uiVcrpbh9Y7wjzOcPI0iEHmGosc
9e6dlLN4B94PNg08gUrIHZUle076XmA7FcoyzON0QOiyoFKZhvJCTTBfuzqV
HOvOKRJ8e/qH6mcLU5i6DOl524MqaqkgCqm58NxUfGJywrtRUa9IgI8pjET6
pUIDTFl3h0uHfd7ksy6jhKjHs7+PGqI8HC2FdRXr4j6YLwXOr1MpcO7na3tH
3OtqBkDz7BU9MeDq90aqExgxRKAE5Zatgm1361NTNR5mWhiZG2Y9SaIgnSvP
Ktm7HH3WYe+R/cmhdLp1nqIBNvjv1Nnt4a0Ykyh5v7lGlRhn+rc95s2UaWG9
mi+u71V8ls9ui/e7M1BWROktng9brqEw8W3G9rdtRdLJFs7lDOmFrPKRrplI
PlNtMYf1eI9QgV39iniEbIikpnV7E3MkkbJvRfdqRSF9t8Jf0auTk7c9z8aq
ydNOwGNFSci1RKIssZyYC6W0nYudwG8P0M3R13ttqnwmcDwAHJa7SgfaDp7L
X+Kdl4m6V3ojOZHt6dLU+84pEg3N04VLMvjfPdnvPOlniKi1jP2bZ4v25Dtf
nvMxsRl/MNqiC7H4KwGgeBwwjTQkVuDDYXSY5a/lAnEQLixfjxA5gjJwcM3Q
jkr3bzDTDgE7YRDzSwAPy8A/5ce21HM+quYs/ZiW6oHSyeCNCfl6EX5Z5Ck0
BI8FafA0U5lMduUkjEGWtxXD7DtnPAGC1SCgnSN3OPRtYzwvfigalzBpf50W
GYZjx3kf+l3aFB09SBKhZQA/Pix80PR1Z5G05Q/OZIiZqNN8g8ykPdglUfTE
IvUNi4aChUiWDvKfcFMPQReuk3fXAE1qEew4YE7caKRzCDWb14lgT2+JPNW4
dWjjMe3YuNZSq8Pys2f3mgFZxOvqRZSazo5Ky1jcwXRm+2nRY/ncSidBjwPu
l9CruVMEUI/CrHNEMqYX8FQsL9sftz7MTbpiDEjz9whqYvRRpuKYl9gnQ0PR
R0b99Z2oJsiq0VcAkv8VJVJSFexI7Mds+cQu1BFC83f3OxU5ApjFzbONC7vY
qC9twl0HwrWn4F9KSQE+VzvJh9y/x+CoH/ejW2lux3OtzDv/V7XCqP6w8vLJ
BWm2IRxZdQBkRU8kmAcjmDyomPrDjzP0CJIht19OZUqniyPvf0jOdm85BHVJ
jGG9o/yE8MCIHZ31GEp0nddXv/hIiAiJfMW+hA5CpPnn+rQEmb4D216IRAEx
rfoz+wOPlBYdK/hDICWloWgvfYTY9fuNEX6EBMqcz1HrAxaQ1WgifnBuCH3+
HjK2MB0ef9PHO3tATY5YT3gnegJAabq9MDllAp/mEU0KZWLwm0FzUnzN/NmH
namivszLFE4NQL0j2MGlYsLhgiRb7vZthI3CJE/JlC1sJuP1jB5TJZHOPpEU
6YHzXgUSQ46cx3JRZmTu7SustcJUlBeL15f9NDUO4V6jxyy8YtCkbMH/SqIy
+9Gg5o14zHFYwoRo3hj4ISAf09U4pONIq3eCfN7Mssix3quKFn3V76UEYxJN
5gLkgL4yAlO8THloLMMOK7nmciqtTbBl/rIngRV4jiwOYptzHUNVXig80SK2
rgLCzP8KpwqWqQhkN6CQ5BnMt73dYgloPdR/l8t0hFZbMq+LqRqVWZdc9y1b
pzq+v0fqMWjv9PnLtqevqARgn39pdIBUr4R7CbTh35tc2Z2aEGabT50YSdCY
tkDZmhctTKQU99mpiIzj6hpCGYXZJ7V7lHSB+wGOwJKmEh/0rnMPQl0UETcE
NHiAKqzbR47iTOdZDl6e+nR2A0grNyYmXz4p3gTggVyE1rfI3kjsIpKnndSL
f5grBJxN9+SKX8DU3T6iAoSoYAMRqViXcynvXeHPg18zDhUKHIUPUnjd5JaY
DPCp29RIvRCSi4uJuIqGP+nQxuarDphI2uY+gywbyKz5l3jQc5bzn1YwYtys
5tk8rHcP3drIDnkaivaKrjPbyWPOFXbZw2RcodWIq6qzlM4veSxKVOT468Lj
Yn1iuw96KSsbw/BQLbaUbYl9lpepi/5DkvvD3NMPYhN/DBVfk5XKlnFgnVw2
Z19MEBBg1dqxOICxa7/Q6kx9IJ8yxPczRICl3MjXhGlIz44Z062cUeua4MgZ
ucq9W+18X/AdCCKpOnTv3+HGMr2kGezCKVOQUpGaWyaMsJHlynzPyiL0mYP8
bbMtouh33ZkKHYya8k34Zl2rNgipaELFw82OywMAoW3V6bNcPLZ9cxk0dKdK
SLZun8ugBseJr/1BLMwFssOsPeZP/n8kOHNdJROGLv6W9y8K0WsiBzGDtWjS
DVwsChNMQPDCkX/4RNdwY96dUBye90ODXbxyql+dRiC1ywj1DeV30EULGZRh
mqC23kEeW2Hy5ztbu6AMD4HULdfvixbVKGdhQHo6ihfHSCJ2zuG5d6CJ25Vj
nQgN5SLCfLQteFzUIxykh36wlKU3RUTNpc8D2hFIlqT96LRj8R4zFEwPNbDN
77C5QpTni9/YE+6PgOeIqHWqd0j8YjeowSwHOfY+H2T/0kv8BxR46GMvN0Vj
t0WzQOzwZqYOSUJ6F3PuEnkfAbG1mzyHNm5KFwm0b6Prj1/XJ6zsXp0TbCYf
xXGmwz0NEqPQ76zqiFClntbdYKFVrhJGE2JiVzgcLrhocKCNLxVi/VO8+G+c
66Y7QBPHCJoFwoKLBrS/E3zqSDZ+JMvth1pXUaczUd9wgm0Nvp/KLxUaI8r4
wGTMm58AmvQsOOVAwnjEW2k6A3N3NPa3tI6DtiEgmVifErOCAQHXJKtHSQkz
jUAdGIs1c7FG7+n3uRe6ClXpgyuA0k9xGlDIiVzg7hb7xUlVxgaYSPNG4mre
FA1Bay8HEp5S+FvEAC5QLPlTkoBIRYCVX14LFv0/kc0454nGitx/DHZJGHXY
K8gc0BlKSXJacn9b76fD7HAal9LZiTBRlD/aLrUbhqll/57DbPQYRvMuWoN9
q8jgjXV/wgidWFVTkGcmjMd9xTfkRF7VnbybT0Y/6vkIwr7sePILiDQEh7xn
fPauWaboeIFi0hcKbxQSlZtbcHOT+BnK/lIvNKUiqigf/kYFF6+kT00dJnNl
TaLmRmuS3XBytio9gNj9/ZiyN/YBt5/zXdOEFhUay712Sw7r48DT2gw/3eul
nJJD+kpBC8UTCA/IIF4i2bcXb3E8iJerQZ0jyBqY8AyeVhzRkX+qf5vxbalO
7BfREiCVi2f1uamZ/4LgPLAZD6M2FvJiBk+tSuJroy2KKrJC9KonL/1tSI0K
+8ImM+Ho3O3pRY3YjJux8mXNthZd6jxPmwrZ8iJDo4foqQBnul4Rr76I+pib
SKN+IXngzXwctQAHuy3jH48QTCENNo0AiEnmd4mmiCjqM26jcE6PxSUTJLcf
8pvSUEIU3GwEOMkJ1hlkuZFAxSor1rfodLbj6r2tlQXcgGvgGs/WDDNkUItB
7fOsNAGGDEOR0urNWqmo2z13vgX31OQ9OucoL8u84hGTziNhHo1jhHK1L3+t
rBlH4blHzt0YlDNXT6oTg/Xm1F66iEIbg2qmbNaxovscH6vpGXvZca3A/K1U
79eEEydijhm7B8uuRFEentisC7TdnFN0+kAz7feQqDRpuI/vyiv+Ailz/6Ab
9wI9qUzTYdfV1IzQAvWSz4UqGDsj9aI/DWwIxmvkJIPi3c4m6w8iL0f40orq
iSfoNc+RspZb79R4tu6nQmPjpV5i9uchgFDvntLjvw6QJy/jqIKYkaZQaAQJ
p1EECt6Xp3Zr6U0hs2J2NWaqvdsDJTlPPfJIos0ynW0tTbKwdZ0aApx87BBz
ARkHs2yRdoxK15RRogrzg4wWZQ75MC15R4YT41BnEB9BKA6YkAvAvSktOEnw
+xfR8Tzwy6orpagylLOuHJ0vJYTwEuiGqfdygck9dbpwT5LHeH6RPk0tkzHz
i6l8d3LcPQeGyXlKtkb5qn6o6eSYYxj6oWTLIV+a0z0NexhM3uFOHnNSJZAo
8f4bb8dowVvhG1xUtig3wt7JyaejBo0ftSL1EtFstuXzbdJmzdsvycNylKV7
jVv5N7HwjCadpVqfd5K90Ljh3DjnnS6E9GwZgiYnQOpiwTRxA30iHbku1G97
HNN0WzMMAMoQleZ6RdzxmkHXDB5Wwr21C3RIcUGz1xVscEeje0YQlJCFPjs+
3/XCyJHjYjCZr2oy8JvxPf8vksExXcCpmajHbtETKf6cD/9GNrmzAf/94mAN
E2REiJ6O7WAxE7QxQ2pgTjYbGtPJeuDIQANBZPwstla+0UZ7q/DW1WVDyMkB
85hyCICZX1GE+gHNcTRs1rOkx3adQbbBNcGc550yE50KGWggs+macU95zacB
3FIVQ6keDudepsrq0IrCZfN3fFn/NJPvRyMGEJJiINFl/3DTyJaf4TecVFD5
FlhbrpXBvuR649wiJNbmNsh24kX8wnPEKD89n0tR8Hotj/XDXE6UOoq3h0GZ
pU11LYulTv9lZ/W9L6C/TB7VH6fOVXALVE9dXkQj7oJrUy+D/4a2Z/qxeP0S
PHMhaO8qdhz8TqC9Sy9WTf8N/jW0AV56zJH9uq3sG+aeItEHBkSWORbi36i9
EKfN6xlL6D5+DrvZI/ExkaW3EQXxcuG1fBa2bxYyK1WDmV2Y2MhZAzp9dYEZ
r+J5v0on/wN7l0oF5y4m1xh5KlrW4M4K+jrdF4sjbyRTwHlYEDeverfbuCep
1yJnMauIEGF0o53RKVaHkQMGUZZl3edD1b84rtM7PiEVQK8EAm22ixYWnbmS
+HWY3DgIjyD5EUCFpJeHMU232SBitcMXrPgoDW9n+AyJyqoSvn0n8uMTB6i7
ViGP0wSS4GdDBmJQ+J3O2G/cG504a/X2CLNMje6n/jwUW5B++zovhjAlPdKd
R/9nj3HE+404VfJsk8aEpZLRn6EcqjqScsscmpDzbff4l5hC/+xFaTpd0rTF
YU5FKc70/vzgDiLyPfEokpWZkMfVaS4hcZbmFt4m93FG1IqdUnNY4AvYx+c3
w2r6kL6VVlKJJUWI0ZbeRhjFjZy7JXPWrKClBGBuKFF4n4Y/GjUBJGwb8+9/
fmyONYNfmQ6k7HxVNwgsntrQ1zpc6pj+x4a/NBDwqz8rTjDtU0gF5mqK6Na/
+lBATaUzAgmi/tXSCpOThXaj0LtuzJT5mrLgY9azLHyb0GTTl9Il4C9RdhOL
w8BUZMA22mcsIQ/wOZB+rPZWcHIO0XHXc5PpAdY+AFMdhV2SpODW7ouRx7oY
3sM4VqlfqpTeudg2wK4YWV3015j8pTwMLB6l+/q9FJ1yR6tOQlpQqvNY+Vui
hdq2Rjwu3Sr62BwzZQSMPCPmoYdvPoTLGz4LONbes3ORjJlaJaTUaTPuw2Pz
SHXGSp0c8+CWqEpjsDSG/LwNiW36caSeyf7R2raLxJagNAqZcn1+vZgKnDZx
89Bg73Y5DV4vLeAMNMSkrrDacI4Ch4wvQuD2bxAGvj4OspVzty0MD5H2Hz+/
iN7OVz9tpwNGCc+J9dmkeUxtJu9AnD0YXHCJYB47IMfjKyDtY9EyYjsDN01v
cDx7sQP0bCIo97TkxBxRbQ0JHZWSlIyV97e5Hn/5mTcZsh21CYHeKMcGv9tz
a/G4uuYSLVlOI5Hnu5/6QZfnWnoV9UkOipLoi/qxr5zK6b/wz1zWmVIKzlcy
1V3T7AZsxBp/0Y0VwP6ZWiJybPZ7oaqq3ixTE19VjrXDkx+thmOWiJ09DC6d
zYCYXCp6LkiaL6f0EpG1Hp5qCM0TLs9OR2dfp+i6QCLD0VQyuXyuaTkE36mu
GNGbb3gi8xOHWaa72vZSzl70sN9jZzkaxb/9i7m8AAtDATT5Aj5ZhfnSf7BD
fWh27+AU6kPHN66D7nmhnepGTC6RZzD0W+Y9pXaIg1tyYQkJvEaLnFT95pAx
7a0f8tPPItebkv2fR8GSXm2gvhGJdcPSDjtHyg8SRRmxbrDZvUwvXTRGfNoI
ZRrfPgARG5lekKXnGTelNTv9PWOo3FGB+bcv/L5iZTYbGu1r73riiM9Gt8Dw
oBrcooTt9B6Io7T4s4xRFnsQVebjyvlA8pBLoIgBNs5OZ59wN8WHpzvIGK4H
rRvtM7hywhof3yVMBHP0m2NmENs/fFCIccwF5ZIM/SZ7THKiSt9XNO9fWiS+
eSDALgWyWU1ZVlsMWnAB1cL7wQaJJ/V9lO33uxSOo/KU6B8oAj+ufX4XKCXb
qYzxzeqEeVgl9QTHQE5AqypBMVD9SIhMeeMK+7oEWmH3j5DDYTN45i84ncXd
qwyBiI2K8tsMXAJuuVPmlo/NjesIySEH92i3vZv07Fe9O1tks4arJFlnw7uj
0qf6HHuL71D2k34ylBRs6+G4wZxImMXkwBNC6r1Aqy0uawV/eQYKdoGi4+rM
5SFVJOVPiyceNxDbxvZW0OxOhcFgCjY2f0pLJpBJ1Mcq7HnlUfDqLFZIkzR6
rsqzo5Q+1yMphgvKnC6SGuEtYP5AyGQ2I3a7elygD9GOtXfjLWSTOU7EeZJt
6J6u27qw7jzxjT61NQytf+HaOXdqT6Dqq19WRYvpM3yYgk310F8h+kV7KpFB
R7tt8Y7KJ8SRYETB+rZF6vn92okeJhlrqoMXrCazdJbsjEbXPhS/Ux8NjcMt
ZKSLXnfHBG/qIRFw6yw5L8Mrk59mOE1KDcKmxlzmtQJEZyCG16R1C7I5j6vs
xjC/1HcuPUJPhfjuJTHQkiDXTF6Y3fPYru1smI3oH3J3LuVYQg09nvIg4zFr
pnD0JKztHcTZncuhwS2nmGsJ7cdSOex9RDJmnkItNqpNfVSiQx7lTDW4iNwB
yllJflZLfvNkc6cYPwNI/JEMwMndWnmO8S8vN+5bReT+cj3/A0PqQuows+lZ
SZJoDHdPf0X7w3EYJbc62vcF6wHNUMVun9c9yAIyTMNvW/bJZBwzczYW7vCR
DlSN0psKQzA1tQenFGhh8EPWHCUGHmMv3c88DeCXkJVf33GbecLqiyFuuQzb
5ukeQWYCWL7eWXvuvvbkDACWxNh57Jpk249pQSaYbIBCHrr7f4eq+TdjvveX
Oy7AXy0LPBfY4Lm3OFGvX0O9LU6BaDLL7F2PxgqGw7+Nd7IFY1Yo9kumoJyX
djtGXkfkffVROBxs8w/3t/NBc4J+7pcv6HAOipyFzRbmYZM/QBh8nnoZPx11
tKt6jJD/BzUJ57dpZcjTGShvw9qR+2aYPzTM8Vsd/Dh55w/hQpN+ultDSuDP
wKFPJQOnbu1QnbEalXpJglYOHXn2htN48pmDMqnkiH9SgJf2+P05gxnRxWaj
Lb55nB+VWyDbhwt3mszlmkz8bp3E1bxp/n6ApPeT14oJWRAUreU1mdDGYCou
SuvJg+oE+Kh+fqyxPYu1cqdIrRrp1tafKymVp0otRlofSBB+hwxk8PayWBRj
dYFSirEvc1z6TZGOiUO4ifBRX/XqPivg/mB9WVsieAGkCiGxdtaaFKCKDg14
QPe1i7uzwzsFm14CoNb3kkAkSeFcOUI7n0f57JmZPs3ywx70RpX0TdT7HKVn
7zzZsPaaqKmG1luhg37Em5tiIKFaCGorVuum4Un+EX5P0LJEgFQpTVqKAHaX
aCSisMZeZDc8yuXLWPeyZuLV673+EdCYJccr2AgyClVEXbGTD3qT0DN3bsiy
V8fH4ok8XsBoaFyTl0lqTASv76DDmv4qCnLWY1eRLY5QQLjLcd92RfyTiaIw
BwrgAkoFZk05TxPsmSozNyHZ5QBCIGuaXZJw4E8SpuPxnEFdrvX6IAHEPlOF
zqi41XT3rMHxlOcv3glda51dHv4ED0pcpm4nzWh/AVdjDO31MeGTBaQ0nIZ+
P3eWlJAHQLzuzYPYp1DqonGWfj5Emk5B2nH8lEMMIq/wb1saWZZOqE8DIZOF
MAzOXc6oOwCWazthbNiaWIVa0gxrL/lQZf+aK+91jUVOZyUQhYYB3KKDQTs+
MPSIGhjid3gX2E6Yin/26P7J9GubxFUxGOw5tfHA2xANiBh/S4dMHSk0iIu0
ibxrQbmnWNDMIAgMlA+2DZ2Z6z/z8C2HDmP5tqglNDGUmV8dzWW22s9EzBeX
gN4fan38PdwO+hZ7yY4DOayLID13OdlXtufUpdam02nOLxd/5rQYyGC+WhW1
FNuMgfPLkx9/PVc0RN2mqzxvoGjarucN1tClD5rkTL06UEszpfNaEUa2WIeL
gGevy/9vGy8MhUZ42VUXsRqPDSo2k3eodcDOUvaFpoDdiFK2PO9IQME8ITv0
Jv/T/ONvxLl6+afzxq2iPLZXjp6LXddAmNgdwPwjT18MXqse20YEnDw28Ze4
kCDP+FGnuT4O5WmaU64hJQOrGTQvbxU/2Dr+RRu8q+pYR8Okx2ifbY2L9/nP
PcdtmIK2RJhUe4pwgTq14wqqyv7wTBHQtqeVUXIDmc8KcMr5LQRLYHKsZy2t
SL0V/Yvx7SClGnHxVceoAvsTSSIH4jS7eXEEEnJHG42aPpEifx0JCnVAQfTl
fP0GaEHME+5sEXqbJlCuESqP0TH0VcNpKc9NhSso5uXvE3yQJI6jaKY09vr4
I8QCrsAzS6RNHofbX6t2MDgMbA2gkjJljJ7lkk57jcA6pmjRcyItSeuxjf+s
q2T92gv9cT6CtHepw02a2uvuMn0XLMbJFLhvt8IWw1djr8hEc+Lr3LbFZGZ4
XNNjeK7sP+/5Q3qKIYzhzLHt2Cli3mKM4wMn/sHnFqe+aLJ+jHg+Oyp+oGe9
LS1I1njmgdbzbtxBfwmSbPwGSkOy24nrsNSFel1n7CJt9fxlXWhhycGerwHe
ns3MQwX8+6wvA0b2WIZfAiuuaCxGC/n80qDYvBGWnDY9TX251VPN1hIyJJwK
XBIFlks1CaMC2eDbe+P4MVd/uYP8S4839buo5h2MaxVGo9Mn/RxtmrWdLQCQ
lPg3x7fFzMB9FGokql8Zj1KTJ/6+wLerUDOpxYCUohnWruINeDkSNzGjYLEP
O+olu+bDXz+C7PEZXCjjKpQ+fdIQPeWqNrXUpUhqdRQs4gGAGwxd5fseJN5i
ao5Ys0FPTIhCUBm/q1XYsjcZaaQcMdtxjI56ixb24NJnJUDuhiGSGZk05zXQ
WGLrvOlfT7DNbmycFDqiu4WG04w5biIz/ve3tRGmsPkIhynZ95Ajo3ehTiuw
Ac0a6MChv8TMoTfB3EovDdJGAaHE/IfeS7mTJJzZO3cj27yZLu8ZAnN6LoZi
OlwiLJQaNF/H7HSXM6+XBVajR1QGTivCAOCt3slv4oujIbJsLUe811VicFaP
dl5OrwArgQtWgKczvje/n/Yryhs8HvdwGvvXmJCTaHlTAhpwP8amAwFv1tnU
izfW7zSwS70gUBCEU3Fa82ZKS4wAbeuF4KO85b1L0e+Ir1wKIPkc5O0RJHoj
P63uzBcK65SObO00tnnfOtnogDeCFY4KGRdKTCTuQARrGq7IFwCPQw7buyE2
uI+9gBeQkNkgW/ESaiexKsIU1iVFgqSN41PtiwPlWPmKsyRxGCnLZ3CQpFiS
CMl9bJj/V0Zv2iHhm+BheY+/Cxl32qhdmGAgyvZYRPPRz0eJuYaHl+O7lJ5D
JuD6mys0RqGsa4YUaVObdHnHiVk4sLMRPzf5Pik91gQTGiDubH/ctezSWhqV
LS8+b5vBZrQzq/YBATehNGREJgQPWUmmvuMGxFtpwgpknKsw0XKE7ozFV6jk
79FoUPs66c1oiCLnRcaBZUjLyHzWSyfnk780pq2pyXKaYEzkNivBtI3KvjpR
emTyC1U7VEaXy18rvgSknf03Tr/ccy/gUbyotBqpBgi/Zn3BYa8BmAygan8U
hM5UiKmPriyipmARm9kSbHM9quneY4NQd0U3Z4E/YX2Ytc6ERInR21aDciu6
2K+ob9FrQO7LtWk1YiShKKeSqvifJ4q503UWtaw4Xz0+ksKJ3ht3Jb5ysNy1
/5gRFtG+CGPssoeEny0LfBVvIcw/U4KI77ERKa9hcNE09HCoZ8GiaiFSfj2v
Nh+vCszwpzuBPKP9ZWnsIgPzoTOZoOkC/HSHhX1BIzLu7PBlMH6FYa8vocjK
aKYta+Jx+UL0/I+bnjzoum4Lwtfu014FqZ1e4Vjk+vWry6y9CWJj4xXs0BeR
lRJuYWdJ+tHeIBRBKUruhSQeXvHNQrnde5mbF2ITQGOFCybXpjz2J/Ar9yXw
OlzOATjV9PWWEcPUX8k3QwuWETK2wfTBpFtdStEekcAiOimct9vMihBSfIwG
6YV7VhMVE8KNtprMmO69vk5fhJa5l6DLHhkqdvUhOwyVRFa4+SATVdwA66Wn
u1bhloS1lEc6XgAMylwWMyjbAjplv4PUv94y0KJdLZJTlVZI3fme3uQ/ny3n
fk3gAVgXcQFRq73NM1cvNSJuk/3yfxTpFQA/+CBkOwIuJ/YNLdd2zUJzEM0a
Og1o4e60aUMipT0+G+FEGiL4EPDXrfzaNdzUwVeFSLFpDx2UFVpHPv+TIduF
kyyctWsWJ36noqovLz9n8ul6U0JMhV9NB3tws2QCqgIEwz7B2hcGqT5ie82W
XvzPjVdDKJzjfHY4kuzosyt4NqlvY+TaprVkh7lmIuOJh+pa3JJo9gB1f1Gy
jRl6BQdFZuK72oMuS+K5bDUQzR5O4yuo/+Y98vp7seay4h0POsxmA9zWcMqA
k0fR68bE60Bdk1/5eZzh1o/NUfKSdPK2opkYSDGeHjDckll3SmxI0vuNs4gF
yrMd9qgiG5J4aZLPEXda9g7JWHz6eV0QnVGEo+ylNIN0rjQMEGgtMXjYRWYM
8hGlWC7cwOmFAx+kO3MDSPLUyiwDrg7VoawWubFCdrVEE6Wgr0wiQUOKuyr3
QEFQ4qEBgdAe1Yt9GeIixl5wBGP2wtGzp/HPs19tfbLjJxDVDcES6Kiuy2Wz
VdvbAVmCeZX4dWnnvlC26RVfhRDj8JcLgdLlIld9SjFykXMDJFVkVoU2mLNP
J5zALpfyc0zqhUBXLPXXSajIFaqaddhe8/y3gI7HT+rzj+i+7uZ5hxZn2XrJ
uu6zQa4P3Di0MDa0Gp5Kcv6BmiUQtUd5wf/fGnFdXCZGSHdT393yy4sToG9H
Qz+BuCFB51loOwoJjR9Du0PQQBJgzlRrX526Y4NYf+BXGSfqU2amrQx9Btoi
Zh1HBedX/5b4C1JPLyZrdDsdGXVy36/gGvPySbn+u6jt1tOzLPKarFdik7Jn
lOpXk0rsQMz/XVhzuTHmPPkGRspFEyCETjRxATY1daad+hfQ2QbZiAdvpKat
v+C8q5oCHHoGeicsFV1HlUYv75uQYs3UYRLybyC3RLha3gx3qRpTLAtzzSjM
AC3/ttPp279tEAstdWXjeNFbHyZQLcl+44eWL/uuRkOpiMzc+kVrxSFQaX1L
v7/MMkaGIRfzP/qSprrpVngW+5iKqVa0WK1d2qRtWFzXt+G4Gsdcrr9YO0Ne
qxwyPuBtbqlyFw79mpHpEyRovqRLZj5SfSt1Z4dCtvLeM9eQnEDviYVXZ9CM
7yX0lzzgHz+u76hUv6FnFZN7in2hETOB4sIFDFY1PaqzeTCnUtkG7MFatA7J
m3YrYpqUu34HyZ9iS67CxvfEdDMGyp0Ppu43wb1SLwYE+d7uai2HBHtNfg9m
E+bGylAitih+jOMc1Z4HaN8Jjzy+EGojsPI+I0zLxeOtV+JoAfe60b4wyAhB
xqpN3Rf/sZwjIJYRul/1q+PF+O/r+v8Dm3HSDQV3ENVmTDEbthnROTdagFSQ
xuma2vMZFXO8UL4MPdH8tAYyjaXR7QGZkIyA5WWVJCbaEaZAZIXn+MlEZLl1
bbJuKv77mzGNE5dXKD2JwAWr4oeWBzEVRwrSyfCMOEmZU52o6jw/KwYAz8Hy
KO6qvyEPrjRxO6Shhv9qIee3FYMg1ZapT/wiiYyk3UJ4Fw11BIFNtuVSB1W8
9tu5lUL8T4ez5FoO9cL+KPJmkBfuRhQn5/Dku40ax98TEMUs14M5R86ZSsLh
uR4JIZCpHn/eALjBiqpJhV+P5XDN0CuWQdpzQcQ3u/VY5ERVxIdD2mkzymfb
wSiFE+KNRWpPh+RNAw0ytYrl6HKH6vByDp6jL4DqfoABcCtD0kOnreLPl+hh
8aNTR904EY1pNTswGi7P2KI7PUPMOjr3jId7CI1RwYybkcroKE8RUQrdkKWr
su0B2Fe8lTAncCEWocKdWjOfi0QJaLXESWPqVLXWDAj8zwrGLVrlcE8zTFWQ
Gj5mtYsOX/i2Af+9S/4friNOBDEGaWKziEhi29FG8tf9pTGwm4UpwDarw0mf
SAIpmPFSgwE9Vh3qEymcharlntzPBUNlb2zkPpbJ147oHw1mJKpM98pipQ2C
nuYKrD+UAMlHC4g5Bpt8KICRWkOlCivMlvgqlpaZQppngUDl+Dc8qQF1i7Zd
cnl9b13rreqsfAnKU5R4VhfuJmEHc+9nCKTth9qxNLqk6DWCo+SZhmCX6H+Q
+ceXVf1jKCfFo7voA2dXxQSJKa4Cp84T9FHWVhNU+KzgW5SDFre0P6HmfDQp
aii3pQZ0A1vJi2FF2g3mXxyRGXyj8GRmGtRxBnzj2vUKgKaWEKMfYTJl5HxW
8C7P0sVlozrtbpEn7r/nIrrzzI9zX/ak/CbgiUdGw8/65oxV6LviBNbsLqti
AkkftKCUrxMv/udSSbuysIV30tQaF7beKf8hXeOzVMujmKIJ1ooPQcanSWrx
hSjob3y42EAClfWr9+N+trK3D/4p//T4xhwLwCADra+bW30KaAi0bMWlkTU3
4XPt9s/kepxS/He6t4IZuu657Z663LOEB5a/xRVFK43YpJXDMAFZxEJ0L0PU
JPMXd/0HwygwbH1yLB7ww9lHUQz3E1pNOf8V7c7ehOJyXdUl59UCH8OMc1+V
gKb677hNI2wMfVmurldruwlqxFAd30IL/GP6AIH3gltVJ/XOF8Jd8ha2xFrw
g8D/ws62AqV2WPkUmdVp4LTyGHX9c7LjHtwZisAOGaf14MmDc97sFJNFyv5y
w2zFN/xxG3GX1rwSGLya1VuaAfT88lFfsnfIEW47MUm2MWxjA84K77hgXLOc
jU/Rb2tM1wyt7/ZZc8R2Gyd1R7EIQvTaWmzG1a0TWgpwPnTOODLhC6uioKAa
6u8IpsK3HHCE2Fcqo/iVN0AxafDDkrLPF/uJvDT10CCMtp5V6o1JXDGgGrDV
d27yHwB9ZP4Mok5C6dZb9+WiT1CxTXC9zHWc2VhFTYvLWb8j7HkLs0lNg3P1
0NJctHE+3eSbRc+h2QYFa87lLKejHlcLbtfazt5fofTe7vyzS+A1wEb/WxuM
/Z100lKYblHJyFgEvn/IqScpLjI0f7ksxIOSb4Lmsuy2S6EBl96jjBdnhN8m
BThp1xZN4adDlEZ9X7AVa8ybEYJ617q2TPHC61MpfPlDDZr7gFUWQJ1sKj5i
Cl69y2r19JU5pDgmzP9KaCDc2s7mD3QtlsuUallheBNsfjJmiCuEwGopXQoc
13YrRXIhmuLWF+wmChyRBF1pIeLQL3hGuZMhpAReDfWS1DoJNEJ3DdSCcRJz
iRskiCHpCBXr6VoJts37ZSeV1gbMrRAdjRy/ZNMWbVSitC/c4O8QkbxNmOMB
K00vezGZNp57pJo6txe2DtH5wDAMaPXxOMECokX7ABw2VxDzf3vPs1z3Cgu/
HqSn8VauekngAt5iv7pRGJG/c0I8VcLuOVgL7A1pxyU0ZP4tO1D7CFeNPVIW
le4rfr0eXQIxTAG87DerkFZmnlZyglZj3Q5oTUytAAkv1RVWoK1dY5py94jI
eoKlUL3qfJM7gAYx+qK8KnuOre20gCSFHycENWYLC4ARd35R1lYKIAgr1dgC
etlwjtnnDJdYpxMlXUixB3nvFsMm12XOe3tObTfnRgagACvVU5ylx+dGMEzG
SWyiu3tG78tJNqLhPsqyqKZC61uJhb0NowjYdmqPnjPNpUQEt6hece0V/ZVK
J7O0V/ol1ojRK963pq8OkeMajLJ65yXUTWxf/uN+1NLOg3izm2+dg6TSJ9W7
lvUFQPPMY/TtfmsoIF60/KqAIQVSDR/dQVI89tfUDdrlBB4D+RzFGU4QBy7X
suzg6k9s1BR3GT6Q31sHFcwMZ+j3yfTHXtuUFl3lCq4MvOdkSmaSBUsWaeEK
N6eAqrXh9TXP4ExWXkjY8nE8Cx2QgT4gGVInpBdPqhLSY/YbIlkmT5q1hj8J
e8SJSIQVcWLth3fdLS5FgM85NOodPO0JZfScwBR8UIz6e8KoFeBp0NE9ggGh
GFPZdxZvSetp82UjyJldqu0Mht8w51MsK/dTPilxA7eiSAfRzsGW18rx3wZx
U2NovRam9Q1Ptbd2It5qdUNmfgd3dETPThXUZH9aWUBcTkm3+77ruRsEEBHx
3MDVLUd7KG95WHi2dicOZZIUpYMQgGnxzfHWlsakuRUOjZpkWElYROzPNcYT
peM7kDJARFo2c18/F+MvkMC5FrwlyyvF2NqupYWryo+2sftnD0U85S1WoItG
HBkFWmjbrXYxsB2UcA8WXumQTQUvQRBYoUbfuUsRm643GO/o65wnaUEbMJtT
S4UKA1/IVhWjwUN5dXYJFOwLN+J7gQRzAQOMn3NiYoOoYXnIrQ4n22jr+Gsq
Zi43Z7W642D4IWWk5U58PLv7hjk6cnsBawyDxRl17LsVAJODsJqAJ1aHdXKc
fGZlzBHPP3Ok3NkeRDbOzp+bSL2GCbAFFOcA+rzQi+L6l8i4tjYG9cv9Uwg3
FL4lWJbBMfOeubLjLk0TzebJLQ/TyNqDXhiqelipRSVgit+Maok3xIosVZKa
0I/5Yh+yqTS2U5hsqPMCnDbfOf90FVSrOzVv6kq9zSVJpV7Ds8ISmL5O5gqx
n8YpNFVaj7KBsRUZ7FZg/Kg0R13GzM5GDEZI8gZgB+iCDG709j089WMCnJpU
bwRYyqQ+03k1ZrrEPBy94QvXhF/dR4MFRLc735T9LSqREXgHv5llkv307nyY
Q+pisfPkQeqbX8rhaM93btRfQpCXMqYGLwUSg3f4I9hW/2gF7IlvFDu1na8h
hg1hYXfpHfN3/xBbfZUo0oVhH/2iwF2ojAdfIH6x5mCGc/Greitxw/1VODAF
8Di99XMzroEBELpfxTp46saW9tMF7D9hqbMIi8vHjesJakqnM4lJey6NmB90
1H7pz6qY76jK768efgY9ta6C+zyoaAhK00C7G+byAxZQpncOAnQOPP+he/iV
VMd83OmItiWHQy9msWZoi/PeQiuVzS4pu5FHfm40FqCBwt47mDDcPtSUFJY8
UAJl3MR7sX//YMj04ggAM4WTupKJ0E55+bsMCDjJcSxA0bfEWm5TlZ+BSqKm
UMAG3wnT5uDrrjlFnfJg4s+51IoFAtjpJjtjml/Gbl8WXl7tuc9RkiJvbmHL
4FGnwtva2RZnkMeAHE97TjhTAI/7w/o2BqSkLHT3Vz6eG34AfDo6AHcO2Hlu
ITZTamGLVFKLx5dVuxZvV9QjFidsZzHD0YEPaSQ2tqaVHFWJBKcUGK5PWnkx
VXB8qvVMCbO4PRCLT3nR1hVIqrVL2d6drJK5wXI/fgCMLr0itlKNJqMKnd+c
ispuwQIXOp9XlaY841WSeCSnxp4HrR8w0cupZuX2JYrj+1Ju90YKd44JhHFL
W8ShHHpxTihKbTZYFiL//Hl88DSa5WGV841zQPOem579fFSp9xbUQ6/YXhcg
PMIHFv2PWe6q15v30ZNqCgVIljfBWuzIcy/aQ+8Sa/wVLa9lyXttVhhpYrqF
UTyhyW0NkyngO6/JwDPKBa+WNRzZr7UJucUjOs0NmW6OB51iLXjDMDSME6q6
NAnTFK/lmUMLXNoqkiH8v7iaZmkEDzAPKZ60/BVmH8XjoKyv0woSXSG9f+Qw
zegxneFR3xZGkK6iheJ8SdnKwluAxipi5WlIUt9mfCh96mCm0aToFEG0b3Hi
7aoLC1raN+lsMgkZLmKNBi33m5+4x4OM5EJ2+ibo1MImvQ7MJVPzrP8In3EK
hWKF20wMuL1iZHyn8vj6GN0ej/RPXVSxt4IRKv2LLfvMBbcI9+JC+wxfRhSb
jlHQp1PXHb+1JJAtq2p00qH8cO+tddYQ4YmjghEcZb9mSwVS+Y0ZreHpbHsX
B0qxD5APtSUrbL7Z0VStQpYiOgiElCqLsfcg4Dja2K1yRS62r0IhFT2HCLdU
vPI5MtAK7TAmwTtt2nJhCYcE7GvLus9ocag+nfcB7pmujaynN65i6KdYDOrL
25vRwi6rJj4C8VPpdRrJGVl2ymN6r/lmQWUHclDmrAeeBqfZUOzDQcKnQSL+
DedsA2tAbh8vHbck45jhvmfhattI0hy0M1JHezHXAInvngvwTaHW1Ad5qTHq
2+7QtFkCv+qRkCtNlVxYPy7YXOVr55OH+sHynwBu4Tc2TC3PvsxbkHw9KgGU
S42YVsucD+98pvJSfNbK5HOqgDOmMRIq7FLzlcIvnZ9D7RBvgl23r1Qtkeff
mas19Foc3+Nu53L85ARKSPMiPaZvVbueOSJ4P4KHvt5Dwa7uQykeTwGOKo5/
fiyYqSXyUizUrQsYT+k9c6YkBFrxbWj+HyJrmX0O7nuHr/XsUwPOboaO/LVr
QGoTeabnRJxbZxQfoiaJ8Ki2PyvIfNCPtYvUG5IJkFkwe3jSp4Fz7tiI0Vok
JtNI9n1FQ1NYVvqQw/8AiaatqspdtQ5QUHUqp5NhqqMjBSa9NKLSo5fFMmeJ
/Hq0OdUQc9seU2Ahv+D+Fc8KahuNzaOwsncWncb4X/EahHO5coZD2nubV1YB
9sVbZYCK2kvr7Q7QBok6/9tOh1xFAOTWVvL+NbTIMMyyEMf2pnPxVGmgCf7m
EzHhDT9/hkNxWKE5vvrS+fwz3Qzd63vLha8oE+il657kpF9LaJ08xKfXJsCL
BEcfodb+5eRLH/iGaETsVDqjSWY6WKCBMU6TGd+W85hvag6XWziRvucxypSR
X1GfbRfbtn6JHM01jbRD/aYbcDRBEWhngpkjQcxfL9hB780vF4WZXUvhdHOu
U+dj95lJACadSPzH3ON2jMkYj5fdisLR7trm/P1gORgfwcV6Nunb6TYn0x6L
MKqvcqvRhFDZ0GLcGmPWtQ10HZAP7wuAU6kgsF+rElNtDAl1woehTRd+vz3v
Tb6dmZid7+fasalZom5rbq3CryNIx+oEMRLR+7THS6zhk2hoWaUq3oMbL7jA
G1fitKj+DMz+zz31if3Ptu+XV79lytqKgyUscNgFvDCX/cXmJUIRzLLAud63
sDbUPl9wAlUUxedVSJw5jj/brLBSJfrhSdDCWEZ8qp2M7dv8iglaPpMEo5OA
x0KBym/t+ADfd+aC65nHpSZ3Z1xn59Lppbs/3Wc3Q+dkb/jWX29R5lBqvd2s
NwgyV1lLIF1zM8kbj4DmDDR7leb7TBvqy5sVFqE2k2inROtaYaexIERjgnDX
mt15daSZijqIO6YhRMcg2Vu91Roparvgu3zZRzGHq/LlUDxKq0uoldjdZOKY
w+YeQAOCcxzDnXhwo7KQ/73V9DxVbAePi64sb21gx6+CCSlPpWEgkLMRw8H6
RxfoMiLbkRtniZO3bzjKdTE0UqLMDa65ZPg6EEF6sC5zqRuVaxMcTOdhb1EJ
vjNtBezf9qwZ0WHOjxVdrzpQ9hLoiK5GkLJkr3fMCKex48ipbOFA3/xIXy1U
mMzii3sRyf3tARMsJ/Ryj4BN3LzJu+G+Ocv4F2lTtylQf7X9KUxtlMNycyXb
/LO3RqY4BhXSPpQIshA2iAaa4TkKeQ30nICi0hFNp0yf+eFO+nFmYJRvqH5b
BBi7fPDnvxh3AFpiF3q7f2IXeilJ5+VQd12Ufwbtn5WuwXE6W7Ih5I/xcvrp
GK3x2fC8YBfhgZRcFs2iCx5dG4jGNZrIZNP/6m6kx6FlFCp0tOgFxb6W2S/m
KBkaQ0kxJ3uBbnGJwN2ekBBuvUVjvTPkB2QISxorzMZnOVqnShSMg4RGWwMT
i6qpz/gfRGGpYr849sQCs5PvZnrYqBZPPkTHgdX9Whv/KWImfVyPz9MtDng4
uKO04TlGmfAAjJQez5Lt6UXCbZz7ceKyY0EVj4ste4iRLH4vwc4v1+iFF4xO
Xyqglnb5FQ6IXJur2RjH20I1AcjL+naqc9mN7jfmO/KTcsQ/wNQ9nBhcCL/i
LXJNWkm+MsWVEsOlFsGXf59fy3iIyMgBlZltsnyduIRpOQCEUo8eSKksVszD
D+sW4DsMoIXilRq7VQ9KQVKp+JlMpHq3ZrLheX6dcVF+P+MX8qxSPguTOpAW
rY0g2CP+GJ27DDf30BcY11wKJ//I4Xmyj7LMjXKv55es2hTHQt97Om38jhay
+l86Dg9CGDyxTjR2dUkeasltU4JCMOKyUAD2iT3kGP+Q1FR/Rm0elElJomyy
QISQSJrrWUhT1ZjRXb0BSsbC8M/RLGD0hrtz50gSu9yf5V+X3i+h+ueZFF2r
vxPM9yiNFlZuPPWBcrvd1DbLsR43eOuTQ4S0HiTPNTnAJ9GXCrnlB7RnPsqz
+S4sAcrDVzbWRqSXP/g0c711/qzE7qep3xXgJxqP+yi6o/qZ+cPwXaeVDA/S
PFjV99g6mCoLVOmYQbNx/ag17Mgb5IF5M2ImbceiYyF0UhXWoTTpVFozdaWd
vvDJueUURsWB9oNRhrAiykAcvaLNUQrgEpJqzRQB0YjY6SRUNbPAwSCBBB7P
KZCthT33qdT4VVuDJVPlv7AN3hSN6+Ml8r6y5FZgzA+UGJemTnE/HdZ8nN6Z
m7Pg7kqAbpOsEV1uhEz0RZhdKH3NuS6x5UcZBf2EnisucFw6aA/fd9kZ/bF7
FxK9N4Oigcdj9EQYPbJA5iJBRT6mGyt1+DtnX6Xx5bVeJGSPFx0BPloTHYys
BM/EdDzR/sAhCu3APJL7uMrdfZgNoSLa5hJ2gd8N+pTKa9eqf3cDr/4YwLyQ
AmxQOEqa6PwbiL0xG7qYEYa3xapl5MSHXS3BmNdv7EoZIjjbLrnoIEODuknb
n4v5mYEeLWF9SeKkMiWyYsDLqLegoSQl/caZXulho+j1up0BEikn6qubrGlP
r8X9F3m8E38ZXcPwLx3WV3fprA/cwBH2BgnX69+Sh4Jt1t8oJodvuz07Hfm9
+xrBaDWDNSRA/KH+kI4/xLFPdtAuPjmOxdTsGBk32ehlufYrXne73iXwgY6/
bg1JKqHEwl6edw3oUfMRHIP4+4B7f6lbjgf0MEMvojYxTIFDzSoHQSJ3yBTg
5DLUgJ0Q98QvDJdpXJjyZipbzrO+hF4XmDtG/p+d0jg4MaGrikgJs7xcCGin
4HWC3KimxDf16GrdwdRLqXeKnswy/UffZZyrUpTxKyDrHCtwuF7lC11U7MRW
rS/00/MASSKMSTBMFCUX08YpSz310JNQWv8R+kW9t4pKgaznmOQ13LXgFBUz
ZR0SOx7Z6zka0q1AY0R7BSRIOW9RE2AQ+Oi0LUpD70EEkpKTOWeY9ijN7OTu
8uFGUwNGnoCnl/hBkOa95rj0Fgn/MyWYW26x2VTm1e5blDrrovY0R7rinsWo
8jyv4Kniyo6LrutCBo3Hw3SmFRQiBNR5AZvNGZu5K6nVUMz2CRfWjkQq1MdN
HPxrNGNLESFao5NvjitooKn0NnRBk8kKG+uoi1+ukwgBr0UitPNrFDRGoN0X
BzcElcP6Ro0aYRGh/36vuJ0UcIn32JqSqAdqQ2CN7TdOHqc+8w5l8gD/XHlQ
7g0gSIXbygbJ38eQnEul9lInVIodWI1uQ03ZlAct2gfTIMBLuNdDaST76TlG
am5/RSjpbRuXrV4ULMSzfihBKuBLngKfSTL5EL0i6TI8uSK0zSU1dPzXAK7R
TZDjG81J/RoSATGiBjOFSMUgVbRCF/+LJ9UN6tXlpQUNshm3ARx3nChF9WRW
fICQazCrbTeQIrugSUhAtOdCAxXumdPHXvovv6TN8oJdcdjArVq7wkW0YaU9
JHFrpWYrlTZcHPb/vyFOJBqLZyS2ELXppVlu/Ex+BK/uRcDKaYvUpsa8QDWg
kAAQiupd2Q5EfrvzQtjNACvFA3BXeBrg+Wat2vWnlaNBBsX6dtcnDUTtm/cv
Y3uQodWmBVKMiMzDU71OAvfFyNvBG5kfZY5uwgMOrS02ldUe5AqvK4C1fvhG
9BNPcISIhUsrfipJ+PQhyQrshgGfuf460BWwkjvvREC91qgJdNwX3MvWpJGW
Dq3n+vDSbwoLyZkfOfkDfKoIw8w0zFsHzxW6z3SI85FpjRncKcVCm899MIhd
8WsbfVAKUOcBQ7wnFwW611CjvyKAGyy2gh5LFI1pyKkb5w4uAcqBPMKuYiHz
C/oS6ZgJ/2Kr5ntuonVpeNHDqW4SqPHM9fMtyuRBV391jT+JTCbgK8R6STSk
khsR2ml7kmqb2LItTHZtqjqEo9UIgkZIDfHnuy9YI9mqbA/ZeUK5zXGHZ5k6
LVYtoxSWGZDH56ntAqoFGBkRWDpCbCUgzlAcEUQ/Wq+JJ3o5Ocd48oMWS6OD
2043/ma8SL4+CPFFGfAPog406697lVIwJS/G+P2lZTTbTPMry/U5wG+Ne/Vj
D7U0j5/yOw+i3EFs5HqSgNsCiZlxpHHTIP9Ci6gxfEe1uNhfuomwM138jHXZ
SCWkj/ycV0olF6xO3649NcXQ3ZwyT+cJPuoDP/1gtXDI7xgc040s3gUV5Vr3
EPmbCFtPAsGsHDATuDUfnbx5XJHlK1D89sIop8MI41uRa0rhcinT0JQtBwnj
EgYThmENt6ibXgIzaBEwr6lWQFLM/l7pyn8DYYTHkK/NHGR5vMwoOlCfxiko
GW5InD2EKOm7J4tSO9lOyMah3SJGgOi47RlAorTQWPS3ymNXRQ/JM2QzEqJh
RcIX1SDxd++Ocr+9vHxJzvcXacSGHFBNz1jVrTxBzGSsox7mGTNfGgPnGEiF
YWVSvqzlcpO83+TeWhMn/B/UDvvYXzsoMm+i8wGcIb1irG9tCvMLr6BxUtPO
hioDqZ6pXr6WcBSH6YY9MGbQeZANF2eOyihm16Flcur2/1PgW0MO1UDj5S+d
984CH9TK45NUvaswCHnCC+aKPjnFPzhuC3zC90W7B7dwBO2+jcKIvplimkGq
dzF0iy1YFuUelStEm7lUmdneyvjLtYwLraF4emAjgSygyVxeq8cDW/0nDIo5
XEHrFYEmMURRhf2RYBv+aXcwT8JGCTqRJMDcN/kMBgKYKXSIV2aj4FV25v4u
ipBwNbJ9cL3z5NK+xGsOj636woDh1QnIrDyxcQpdQLgfuMkrInWqZ2x5FpJu
d6T/Ihzp1gQELSSzRP3PdKSaSPDtv5rXwE/I/gegDDfRGOeIN664KSgx/qq+
clgjK6IB93whMOivbR/AJAdZgbrJX/t8puyclC5i1BY1qaYIz6U9wkKwubm4
j8xeSduKbDnI3P5xoPxr30VoNGb1LUSIKw3Oqd6/m2ovMcdpVmwsenuU1xX3
4ARPS13b2P6sAQR2PlBW+qD6JCJ2diaVKWoinm9R8//KiOTwdDTJDekQvqHL
Uq2V8WyMizDH/ggVOQ6I+LR8rbVYxSMpBa/h+ccvapAvjV9AH5q7VojzBt+S
ru9Xu3T6yC1PBtnD6DSkzzLFkpNixxMJsRNoqR063XbiRl2wp7oA1FYOyh03
NXcvFgMuLwcZAYjFbyjwhiAJXCWDj34PIdIAeU6NFH6KGx9zcqZNJnhILIC9
PBBBQR6RRcnCNOP+5DGuNcjWsGbt5Ch9h9LbQcOFNibeZATb+OtIPWDm/W/t
hisgYwSo6XvPgVlrUgVbZHpF6egByz8QhjuVih73ltDdN4CSx0SXAEcD7ux8
BtKcgmlruJ37zi6L7NWfy5cN+jjhO4lmWSjdQqMCeNypPu7JnVEvjkDm+k+S
JTl5g09ehlqlpwDsQCAMka1ZH+qfPDlV8BudsQXWjPZL7SKdC7hc6zuQziJz
PS2uEevAuCyJUpTauPcvWdsZWWBLe7a8+enIL+VSa6Zb0NbV5w4/Uga1hKgz
DlGaUj8vz1GKDbAjepNC56W0JlWU54FSDofGMwHsjR3iurS5/yXS7ai8e/T8
URpWy5bH30EUKit6/EKxWYYo2VH9k5Tsp/1+eMFKa9AQaO+iDvtbd3gCG6/O
E/zt68u31j+sp+vQCZuIIhFaXaGHpBgt4kVWB6QgMmEKSmlO+L5DKU0Uhzbm
NbbjpmjPvEBIbBC5GTvSUsb3d1GC1H7Dz7en7a6DChT6lRdIg7mQY0qeBJlI
eOtqCKQruFYlDr4HDk2fgACufGZW1LTCRuByLQw+Wjia8kgclaIz77YBAWfW
1IRl+BMnY72Mk8t3DP3XuDPWwG8y9KhBiZjvFyYgONSQaMOiyaw+BzWOxDlV
3JiEDEo0yYNHY6CSu9pzAAQqKRw7ksodPxjTwD+wi/zM6NpYfIx7wIUxFGW5
iaCeBnNun9RlRz1jlHwptnmursn1bU1uSE5sF11BVb1HVlzPB9M9NE23L4Qn
xD83SeTTt2W/pozjRGqil4ulP6WrYIJ5ME33+bhTK/dBMYWW1HXk0MNETCsy
ApECUuhzj5P8/6t0dRMecZ0mj80nSMU2jnFc6BCkRtBpCQColYWjw8XSokXt
ir5uOkN3xxeqLDk7h55uAYdDu8CZ1Vn5eQcAim0H7FTJv8ieSIqfyWasXloW
hDe0+ECB48Pe+K6Znpyew79f1lhcxGSEHa9ctYiI/IbVV/EiythgQVjHfC2A
cV42gs6H00w5PiO6vwxIPGDXp1rsYGTA7RDTL9JZMLE5qyJ66XsfBWLz/Xhx
n8dqlxCSU+FFOKgkQV8Pipjnv+pqH0wyNC14K3/vytG5lvU4ptFodESP/os0
JEPxsVpCV6l3UlmwtjaiKbNzXoD5fFeeg+2+bmECN51M3iHiR7WLPsA6hh16
Pb2591Q8CJU/1DnvRxEikkPmuY6cbneUfO7hsGSJZ8/GNeRElSDoTOVchjpC
I83lXNJI/R1/ySS4Zhqe1ZxXry9fT0lVsGk/D0Z9DoAB+NZZBBm6JVv2u6Wl
+QgWtVp7OhN31pe0MTsZUzu2qEkw+Yq6n1AfRnPFhQn8kNBiuaf4151XS/q0
FuVlOuPcNJa6wM/BA2aYzBXPTJ06zwcJCwN0DqIrw4tQMJttEJK7s+cr6Fcb
iHUkbGDgVLuESMC/UKA9D37d06DIaqdwg/ZBBjPMvUpYE5K/5O5LGDs9xjKk
JJ0xn7llYPWbfzqMq/8vfe/JfzvMpBpwBtmP8vLEWd21syWBTrU1y02UjX3f
quiDeRaaCq5touY3Z7XclAd7Y5sqZZ7lvPiAvN0+sjd4tjv3fb+Dclt92+bF
KmmMWNuyfICVmxjU699Obb5ub3AoExirkwZJn12w42YUoFePVPNqIFjlb8WT
xC7gr2b8p6MX9zUHXt/qmTd6QaRZ3gnOIz1kOBy+rwm1DYQ2vw6Qd6Yc5odf
8QQjaPyjZapPOcq/nk/hC2VFs2xih3fZvHpgCFwvjTdxrnapYG2PRTEf7JDe
KigOcAmuPc1MNnvOXFRaynBMe3bn6WwR5Eet7/zvAlCaDHC40Yg+hp2egato
LwCLHRPNt9kKTIzUkmEyWF02+8lTqPPpT8DkdU7ZZGzVKdAhvcoSEeyxVEom
8BH5c0Gua3a/HL7TRSdSr513iMMaRC8UeVe0pe3lsgFKI/07k2kc0Tzp0Rn2
XDXEtynxt+nkwMjtBa0c2HYP2w9FAsYqjrHqTYUoX8T3scE4oF/LGhHsT5Fi
p0XZtafvs4Cs+kT9dHa6A5yiDoiH8s7vmq6+R6BCtoObT5/8K5GlYA9P5qq6
hfDfOTQIUyhXPv8ZqNcSgF7r1A0r9CmCMJG0HfEHpixHeJCKw9F0qfVRlg9y
WEs0o1dQXIA/F7wqswUkxyf4FhollmhwLcq1MRT5ZL8zTt+3FNsKJTIV5caJ
6ltk+DW76JM5ahYxX0XYy4HVvvl9YiuRmIFDzixFhiP1OybfXEnawy6cFdDn
drY/aF68XpNbIAXhhU5XP72hiuszges7Ur8YwoNqI1WFSnAWsQfqk6ewpKiG
mgtb0PflHj6Iz53B8yGh6OorB1T7/f4x0AKbo2MBdcKLINuqI4N7NGo1ZDTw
JTHL1bQOV4IPqmuO9ifX+XSgBIJJCB1x5WEckY14IferIp3L52coK1Bm3pmg
2GHQp0G0WFvpU5qvV4zyh8PxtH6davPMefaVPihiVLHc7Kt1lhLiFJ/yhip+
AnapsaIQAh2WsNMkUpKdS4Y6MNr2h4f6cnbUJrepvbbro0OhK/TCu1neJXN8
oxHPg+7nMMF8YdsioL8oAJMhoaZglyYOQCMdEcBp2w/1N/3WxjvTv2u87WiV
UzxpwOSjCdFGJfkyf1qvSxfP56QzEzhfEaxw6CRakUL3QJFybeBgTZgGAv++
a6X/1fWaKkmPd46AkPCAnVver5k9DStqTkgqcm4WsDP36UWO+MbsLBAFaa5I
aNk85F55LRMoSaeNV0QjwYhPn7tyF1nPdEU5yuk3nr9JWq57pfvm3TuQ04V7
GWMMUJIyHoFDkzFdvdSixHpolA3qQW92u8Wtr8fMXe69tTsb269QWvfK64u+
ITISU+M+LdA0+P3WNnI3OI36iH0LS44T4C3zW7JhneNR2gv7URgEaNrW4Hgm
Wcin985VMkkV+PwBRc9g/FtKozYoB+avrMhodpRvMANDXMBXteel1mouM6ks
ZY3WPKk4yf8eDBW/c6U3VJ1yW75E9ic5ocfS5mTzG0HAgUphsI44vR14+lII
vyvWMdj2dTuhDOVCbto92dYWaUuxr+1HkFLRGKqZYwpEtw1Hl0R1Ur5DtuMD
NDdiGjyWYn2q9c/igVrozpFarnCVx/JV4l+4wfr9/Oc8MxpximcPMKQ/5UJG
JKFMF99IvgFHbVLm2r86BB79XZd7pGc+8cZiTw93p6DjLsYcpgQejyso1Nc5
JlHt163du6ZmWTHDfdjEpM5RhkFIg6AqTETh/3lM6LpKu/oukquei3lUmD5C
Xva10m2rb9iqPzh7pg0PDeIIAUicCPNW/N95B0Dpp9RMnEf0pnd0UM6ap0XS
oeFQpl7ugw3wBLCDLSXG5ZkTD/hwbyZW7o7dLabQd+QpHkYsBZin6x6Cd8UQ
bgG1pRRRqtuAcNg/rMz5Kc05gYs6CkXuabzg+y5wXEWUOZ9pPTBPMaOo4kgO
SDTHTA4joU10NNpeeHGXmw3RQ6l+HwsPbCxMhIsYHUy5qvVj/qlaxmz3dCcl
Gc9NwBqODXs9BwazkrFXTZ/yLeNDg0YF6XwzMOKs7TuVc7xkHt7wT8eCAU8A
oXdi/Wn9xhYO5zrEoufSVhBYykb1tvBXVhpv45PToWPeY3wquH/SiD0mIJP+
6B90SMWk1E9wsyre/2B6Q4Yn+xGJTuHLQvt1KDUr/967H4/FYMsRCNqqCcTy
IPzHX5xaZvMQuCH3bn3i2CYGOUu5L3jpBKYVc4jhcZnnVjeqUhWi3S10EQ+F
NfEC1GwaLSx2s2MOncsdTuapjKjMUik9aCAMTp2EQxHswko08zUkjOIgv4pM
wWJya67tJkB1DBQFS06qf5G8w2dINe7n+RxpfPYu+p73dNCbrAEaCFi2lYxV
H9MYUUr/3aZhhuLKAW4txhuzCkt4Q89TPW+uWBbmiXuxpSmW/Xbsc4eZRiRi
D5ygQfD9D4r1yNIHaoUkNnQtjiK+TGLnCGvuuUHNG6N0gJXwyKHf5CJ27iNT
9xJpFDUGeczVuDzGNAKWYC4rKa1v9yJXeYkfMHBzcGTH1b49VJy0sZPcStpO
UrDMzvjDFiuYjS3V02ViOSpK3UmlNDVpahQ1WbgNGkRhuBTjxAxY9V9EMSPl
5wrV5cDnDVq1wG8ozkYz+DYnrvOg5j3Q7QBPYyK1ZW6iOCAph4/tDu2MVCkf
PMELJALDdfAGH8xEx9Fg14UiOhALagx72zZz+/E5o9j324/yX8acnx3mhKtO
++S0vBEONhizAGTq+Sl2e9zvYZY6yZ4Zuvs4doJxfW9nug1GoYcUFiHby+vq
3rn1sNjpHdLMbWNVgHVr8xXdYFcqpnPYBkGWC+Ddf+/Cwt//H3sVI6Zb23wj
dE4OwutjC4gW18mdPuc99/5120KJlokabOn9+v148BV5Lrb6dOLu1HqAMzjN
GXWuFsRL6aoPd9c58/0QjlyFYmnNkQkV9XGj19OdfVaOHnaPOQ3EY9tUiaK7
lMhdXPQmvtpV2N9hy91BiJCrT2pGQns3HT5rdJ4yGaCdueF7bt0mf1/C55m9
2sZcf1X1XLTSZl43iW1/Hbi3cDae/r0TRFPwnsK80VtpErK6ZZbSewXjBs3j
5DnhI08uqcdIV9mBNndlg5+gi/nFMVmFVYZEfF5pwNNYWHnZYEne3fKpy/d8
alP5c2UFJHA9spUQPM7njcyn7/KL+5qJmzVaSssYyOcsInGOyX/4n0/bTO3p
Dwm+7DDwendNzGXQKsYZzPUOVv3z0AFaAoub5EAQYhhk844XnrlhHOjy9kSg
JnCxCRiXtGLreXZ7YW58ezdoN8wnnpn4LrznlTvZTht41V9GMtDscNngCi6s
OXdTPD1Vh4fn+TN7MpK8DW5Vir2HLNx3k9wUw8zUSJtJhXmtET3NgKmtz6nm
i1A7elzj7a3krO7pDrBlcruY4awgXIn0kyhju/lRCUXvMNMmIBud/iZ7/5uY
jDFavc5GQ+L7teaM4ORtxfqZF5BWMURgzqowl6MMIcjgAqvrEYHSjztZhNq0
qW82Nszvss/AS7IsMB+gYNbmk9ekkT4IoOrJpYqE9AqRs/rT8H3AUd8AuHaZ
4kyD8DNJxEtE34XOmgXWpv3LhQLJK+3OpGI2EM6GZKjXik2J0PvxWXitY8B3
Bbq81dY9DL8DZAJGovzxYrG7qyKPXW6ICiUWx2c1RNhs5OGWKtDFTnuFvr7z
DzzxrDPqZBnUPW3iDddN+b+QLVZEAKW2hsVG9zu9d6GQd8RZ2NXr3dCQskc5
tAqPeyfKMuWv2r1OXq049mZ/T/uAXFuUkFGYcypwpYAnw7HnGI/didMUHoRl
EoYi2broa7dUgAM3zY5/Hu+jxf4cSAn8srz1l1/i4ydFu073GJPXGfG3R0Bc
rjrtcienaRRGvTs4/k6jtTYKOus061ctaKkuuZujbiMSj1zEI/6wb7qrQmz5
uQQfPgqkCYlFvv01PQkg7bQrqO4ZtFhtR5vgXfDozjrmmA3gg/DFluzdR5Uj
JLru/h28htk1n72dJcXIQXnr4uGNTj95EVvwarSbHV3KNYcvLUQODHDVsmMK
NMDyHSE0Yn40PSKE3alEZISxKL7Up2mzn32OfhUR8Bcy3kiUNi4SA/gtcuLa
aPnLSvsHK7t+jupiXAFqwyMM33hZJF4jzfuGuSlJAJ7CS1r0GeYGLseH2svy
5CLb5lvajYcGs4OsdmnEo3Vjtrn0XkZn2PqnDz7A8FEwMunaRjGQv1iFFv+D
ENMqoETFmZsPreIfN2eCItgye0KS3LkpQGGkOUCUt3La1KK5b1jwTWnA7bzk
qLvSCTJu9tMWOiRPedIxZzuy3B/4gsGRpZ086zYh11bjJAKyZWkL7CDm4Fj1
G3+SAIKJurMpNU9/mgZ7kQHY4dgkItHkQhPObPGcizmELKtXR5juySu3kfew
IqKbQZTm7ICTj18M7Gk3qF+VsNdrzduW+U64WjrMW6r1AyoLLN8iyKFXbkq+
/Joj/kkxdzmROegCod89AMUTVaFX2jxcVNNFTGh1N8Z4gmqZhOHHyIntGyLO
7ipThL9vokAw1eX67BHIwzDKLu7pArNnZM/iXr5YXZeQm2p4uBRhU6rjqeX5
H4407Mpbbt4AmbEr4y/NjE+psSA5+l4uvKMcqMretxHyFhxdzPPThmGm856H
x0UBCCsMAZj3+WxP1edicTIlxEC3OKXb9L10PnW1L3QkI8Szidlp5Tw3JUai
gAygfKiuFRVaVheiXokoZrGwud5ULICCQFY0BZ8ReGHR6tIUa4AKEH7T5QEO
UV9KbNlFcQVNh1GwCvYMFsUfqCxpWzVhESPJlty4kOSbTW7gEGn4M0B0RmyP
MIuL5YgkQGkItB9l9rFGUXJdFgO8Q199pBACPUrUs+wtzftD/z4XKilDeg/h
VaolMCMEW/VagTHB6rQgVlrBbB6Tz8GTeUFkLiknVGjJiO1Cl6bTopbcSO/m
p/SY2OMunnYbWWK+trV+rPyIW8PmNfF8g00N+UGk92ivrbopvegVkRfIYBVz
U5lAskmjc4AmuqKay3Ft7j7rQla421erYDOL0x1Wa2aUY3pNXca8LbpzSxBM
2haASvplKwY2pOK2ofw7bYee/toLeWhzdBc09r0p5AwDMOqeyGpHEp65/tOk
XinsyRgVx/cG5ctYiVqU/7o7v3kLKFZyPN7m0Y2S0DAW3OpQBVRoTT2Px6GU
RYcFwdIVwXPveT72KwMpGRV5SAeeXNU+lKxv4rtYYQhpktgG5MnnDsuP6v00
raIQRDN55AkA0ClxkORfGsbL+aJ1xt04jxGQuQeDQpiGyl1F+yGFDugD/BxL
93kow9DC2FnujEuslYzwUFoxe7k5CsGR7hKpU29jZIjPWUnRRJpR/dQLBpoo
LYfCbCia6QhrO4LXYvrBVrHV/dLkxRN7+RkIGu1+5/luysX5VTagAq9S6dn2
NwXe6yEW/rJ3GWT2kJtEr3634Yn0rh2jsjwyP5FRnKK+TxbwinuuqB+pI5sX
NmhJ9nhSN9vAe+22Mig4mKTzwlo90xoAjrWMsVRhnIz3XTNz3qqwdmBQde8g
Ruzd48C5lNyTqBWXHhuuxbvhVnXe6Yc6M6M1KkMi+Hx2jP5dqXdFPwnMsvwM
DFXa6MX2zWbUuDPQkn4ctvzKmzV9lhTVXsVkF2U54QxCXz7X7CqNmvVE+se6
XPS4gAfGUAEnwpV26/VXyOpztQmvcpk0X7ThMWerCD7yvMCrMXRPf+623tCq
IF5YpwMTRETh1+RmY3uyNCKy6oL1bDwECxRAh1wR4UMjfReqiyne9qOBmTUt
LeAmhtDs9Prpl/zecakJUSTAtdANVzOrGvZhX48WNzTYgNOIW1diiYRTdGjw
XFSTIuxVQLeHIKo+vSxDMMojB69SyZ/VVX7A3SwRsJtiy1tsuxaMW77Q37/Y
U35zyXmkVNZShbDzgCf/vrsBqUISNybxBVLP3/K5U/lrOeLcGt3Zhixn8bSB
RhE+ze6o0SiqaabuN6LbZjI9r777ZiiFEWxvY0xU3cLn2c5W346wrKuIuf1W
z19RSMFa6ZydL9q3Sv3GztQgomVdVZXDIL/Q1IIqVnKXjXDD8W4rlWp66nkd
JUIHENjKwn0WQFw96nNfpFHvVMBRUsz2hluo3W9VFWNXbnhOwSlL/eBKB99y
+n3+BQPHCa6Rj8vbScJeYAutUrp1lqezcKqkqNCkGfmDc+Sxtc+5Hps4ql4c
pJtlQPmqocFZpP3OvavUCIS9Vl+C/JQwjIQNVIMy/ynU3clkNtKMA4nRg2LK
590lYcUj37NW66rdSsDyTCG+bC/TWj+P2onadjiqsX3NsGgkiMnIA/ZTrt0R
Ao6yd7HYAKlGiQFlZ9Y3R7UAo43AcZnIg0JYCAvAR0MJu0OKcAT1FjspOMO4
XTAXOOZaT+rv9X2UHANPlWTyoSq6TvtW3TThmdd37tYuD3lVWHuN7L76CAe8
Xhs+REqu93bbzU/PesXyF4xHsimAwcuA+dsb1NUr6i3O0XFMk65gl/BKYhX8
SjXnSlV+MwD8D1SHY377YdPlTXTg3fJarLlrSPgpqA11AweMOALgdHePbQHj
PSbvw+JJz0oOACz56cTjQGbDe4SWUpLPNUimLdP7R3qWv1WQr6/tBr7hMxT+
y03qys2eWcQF0cA07OuyF7xc8m/jfVvNoQDSRz7erptkVmdY6q05vw3LFEgx
B1HtFR+miUddjzN+mwSbSjM1L2hlRfsVtqQjKfW3ovOcR1a7vjGGhZR6irJR
/Xl5eD3r5+eCPtdJR9iMIDQBKuVn2ODsm8Ifnav4v0SALt1OB77MekX9Zw+m
ao8xWbeMZBi4BDfC8OubWcClYY9/owIDHAK2ruT9P6cQp0blyUdieaw9H2EU
Cz6/mkCWkuVOCkyTjNX9ygBUJKp5puzlmMvovuD4TyKFS8YATEWz4esj9iY9
bbeD76qI+v1xIYrU6IKh/RG1yH/w7rTvhGJJaFY2AL4WgAzc5dAPw9hZJElN
XgjwzawH8hqBiDecE1NGl/efJ5OEU//GE3NvGHFhPVPGRhEiRj+qB+EBI8IF
lfsbI5aZhv36MyBos4megNy2ieE2orwOTve3R2x/no57ASklRQMoCP5tOdRk
Suy0Gp3QYNLjQ2tg6Ep8O1Bdltb9Fitr10SgYsn+BfLOag6N6eSEnqFKEFHP
s2qW8GteQSuNJA1d5Smfm3gnx4tlj2Ixi7WTB8pZV50oBWH/oJIb3vIB5XGH
pZXEitjZx5dw5N9TVAeUQt+Yy3INkcqlVfWwcKSe1AKk03XDHeRMMxnP/3eR
nTQz2Y3CZknhZ+IGeshHFnAuGp743vsnW0JF3LN5gsEzkYKiXUECwzfe3WuG
aqIJs8oRzvfPk87VuMHdMK/tmbxLsgS7FlGtKGKS35AVNLCrlbh7Xo00K8/K
55JOynAZ2SUXcxVnOoSsCXPUMB7JPnZbg0SbJ8boDTJYJ7MqtzCZnKw0UqBz
Prsrk8xFQ1BwWm1J4RTdyrckhCIvqr7+tVDZ70630ay9/+Q0BB+PdlTQku7j
Xpra25ZRaP5RgbabfKv6sNqo0VzaaCBJRk7b/PEviXe3iy8qySlTvXYZeIHH
3iWhzMp2eX27XoTqBFLIArd8Wcia+M8nAXTkYHCeiWZvVj8F6aU+PwDcfr97
ePAOn9sGY/rYgcARhleNQRJTd7KfioFCJ12ql2D0zi+xYwGzSo6VQdxJYTkM
923KgWR6x0aB+iaysQDR1/ctIUBYegRLRrcXtGkuxJet3zq/jGkLJoIsMdRD
hIcMDgYg5L3sXdc3pIwurMxJAIn7rj1oQ2hHSpxxNPt//QXiafhKV+PKqJ8Q
3pMhR0OXLMhUyk3aT/911aSLw3pYUthARgACoi1IJ7DJpa+uCS1uzeRIwrwx
H7GGRMMFS5QZGQ2xhnAUV+IKdkhF42g7aCr6qURIiw3ce+h6e4vCi2Sw3heb
A756cIMX4Uvsa2EejEkT5dgIVa+Hv9Z92rkoKQ7hFfeufUQEm58XlZK1Qvn/
7kEMiwVRM4CeLdaNV0swH4M4EvmvqoyWxKeP2VhaoD20u6YIicjSzlzXSETJ
CbTVLNg9xJGdlzbCcPcFjfLpSaPnmCXFwLuq1hPWluRFXB6XlbGoVWewZOSt
UfbaPatEqt+9ZsZ4OqYqFiuhPcALVp05T+8wjsNQ2fQf7aFs4GQ7xfLTIKea
orimbbinwLcxCWTLdUrGF0wg7WxVPY14Tl2MFbIBiD0EdmoL3l0Ez5KGV9WU
KO562HkBHRoofFSpAje2SgcJO7woaGTcog5cWnmRcDvAHf/TmlgbTjQZGd/p
HMBlaJIwSr1eGcM5QBO/6Jigr43uW48EN1pUj1+cuRKnlDX31V5sHlxjRrBZ
krJTxslNfFA77jLR5QDkrpXDGbKUGfX/dPBQ90zaFZs8ZW3cLC5pyF5NDfKa
MdhdKWVjUNsYYdgUpMzReJiVl02kSpgHb3T5ZH49EQfRvO+uAl2SIRMeH3R6
nkgdSgg14wpR37t5q3XHPu85Kmd0q9P6mp+FfGSFcvAak/wjUkSRoWc+6zLD
IET0HDbdvH73nbHZi4Y3sdzN68H7/eBDn1sXYp9LbGmkB2+PRSDVEHOb9eL6
C2l2QTSJQH0noattO+RfLaRXKVrK82kNlHQaoqCK9ZZtUOoB9SNdF3fwmcBH
vzkwtQeeHnN871LhG3sG88OQJzeASR5QLswlT7QlnvTEoGeKgwVcAsLjAZJr
pFnTroPqncCmSuMuuKOcsWUKMCfargXKabGQNRhxkT+NlKBK5CUZnlKcEmDu
5/jPBWDvIYA0buTHzVMkoD3v/LktxBc+UYwlV07H6K7M//TJmVi2WJJUn227
+cH56iRVh7s09dbOMzcmuNxqtrhPQCecI/hhsAZra12XgCdoPXC6h8emt25L
Lzy5keFFostsLSdnf0zKhDFQPQOrNBjVwfzc9s5Si0QliNgGBakTgeWy83/n
ZGbRwBtFNVF/0YiEpifCNPSssCjJ+Ck4S97yMNEwNBM2BM0vMhQ+mnKoxyuP
+BNZi8PtNkyLIZExbThx1HQ/YwSiIUod0fl/HQpI4LJjxM2xBxc2PdHX6fqX
watrb/jlSD8feKScecqRPWasiQkHC5BtoQR4vT643qFCGbaCJHDI1V7gVsNN
39Tku/s3WI6p4ATDrdh7b8vj5ZGMQMCQM0y2OBge/0vaws+qDTs7oItsNxD7
TzC54J/TQBT4VQtembZCi57V7Of69bCn8j2ZbIP2XwasB8kdXpN3BfNNxv2y
H2/mmo7g2As/bv5wd8I9+tjfPAFdeR8+DfQ3SyrtIPzNk7HZIgA+2FcBu4PT
dtHL1XbED02nzoGct1O6t+hVQdwu+mm4GAnQhstLDVqZWOsJe2ksnU2YC+s+
dOQNPXV3bPFasNw0NB8vXiOFVoa96l2VvTKFrcZdYazWIj+ed0BepUNrBCMi
MtQs56b7Z5UST08TT6kKHi3k9Ws4jMqngpYVZfq0pBTpZXex03LcM0yVho7s
dpntkCvdK9FIcUKDuWeMSkSBKQleVfsyI4mrChgwtaQGKrMof87euqDmHl3V
h7fiTzseUD9d3dBendN1opR3ViTzz4CaAQkCgQLFtgQ+kP/oC8Ym+zX7eHB5
t8s84T1XTkH2QgqEtW8oASlbi2R3pEwZsUzWE+iEGF3NpnrW7RKIOWsfH/Qw
ppp5jWnnGjOk/M7nGA5DGltrFo0BSuF+2tDviX6dC8JbQG/eTcinjO8v2tqO
4z2UXMJngjpPVYL8KaBQLocd0VNXfdgcVERM/HDN+0GobknlsXIrLXacFazB
bJMGBBmTEoWVebFXOGUkrv02D2P9mJ+zleKq+4gCNuA90mBkGEHqk93b034T
5OO8w5H54W7lXCyPrqwbgUGXIhyHm5I5GMvpcj9Rxu3UaZVyxEde76bCUNr6
mArbSLEht7aPfzLQ9n2DwhZExnxN3c+v7MPUy+BwF5Ld75VtFmhn5enxaBOl
BjIPHBwzDkKxpkwnLcHvtd0oWK1PXJQ6fbCUC9Dx3LIuPTvJe2AYrHn5Wzs8
ej8nU6VWQqyS6rs0BGrmHpcpkqsvHNiBpl4l8zO1SIXKrC6sbI/4NSNDEjv8
5zzzgcxVKmtui8mUTWnnrz+sQUAAFb9zflpObhWoArCdBZ3mih46jdVJJBHL
995gIcDp8fcVBXSICpUAMVvvfnjtAMuTrDy9YfsRJJLYK9I53t+oszqaRGPN
573Op19xVdxgTwHrru0teGdFOBoVjpCNJ6XUGeIt3QoiVfW/1xAQBTarRfIm
nJOwepjj671eFLLsvP7RIQCve4fpTo8bq6APzQmT3MeWccAg0PVOhxSdY9kR
p8Ns6rlJFp7Ull2QLWj3B/FkQbjSmTqNwL0l3w42vX+ZU/o+fjCJxvAK2GTb
ddZoT91bX6HQMz86eqARGhKF9VzfdDIdYyrcJ3MVtvdRkAZzN2A8BmxiBz4h
To0Kz1TD1+vRKk8iCcXl2Mpqo8Z/9LcntcIUJbVeq5aV1GJhUoNC/0Y6pIia
/jN+38ZdW95rRCLpAIcQMiPgpkZieFS2aJ3Cc/FEOqENPR8hgJDN4KnxeKe4
no8t5m1Wb6OsNSoMMr6RHxFEJaawNGERxhgOb0lBMy1PQ16o5ybm7aD6sXVB
Ma90wXwKvZddrvQApzrd7t57THW29cIrG5mI9rlmv72QgXZnU6lhGrMfwkP5
yvjJwroFDM3LGS/k5VaPg76fGX5DJ+nE4tJK4La6tNqwg/fLGuoAhOQNxaOQ
COjLjl7uYIRkOrugBRSPa9UzSqIpjV03m+dYCU4l5h7gzTqs/ua8Q7RcepEC
f+R0hGT06lG0DYb7Y4xd+JVYAJW3vuqxTJGu4EkbqqsRVzZJT+M6GRYGeBpp
Q929cXQYlrDTOpsIFmM8bVuKVI0/a4Wiz/hjRAat2rHanxvKkVeRNWCzPMjG
IAiLR71sM8raJFMAkh3jtysw834VB3k3gV5ddki6PjrN6Tg2mmESUO4ewf3B
J4hbGW3eyxOzonlHKmZWL+kmHlMeIDYcLNLTMKCr5+CijozwjeUt65O6mRwR
s1BQbdel38suJH0ZY9Bfv1jdte1hra0x85/8MyZeOjlbnykblAMazsjZoEGE
8xBuOWSodetSEUDSetwXCJ4zCJ8yMzUAbBAJ7R/UCyW2m/K4c82+fq0mokR4
Pf4dIiHyK7blLEXxhB4Q+s2bRPwXQDl17MAFb0d76PN+2zgMHW+xa6KIqJfC
NsowlChJD4lWpF8AHUIcAe0UJw/e95IMP3DwIn75ZOTZF2v/I6/uSNf85A+E
RylbsmX+zeWyepMWtqsep/IJkaUX4x/3W13PZdsAfSooCRpn0j2Z0Lp2E9NI
DKoXPs5rdNehYTV70RijnxWKUBYjtd7PJM1TOpOoOviLOlzoA/eH0wuok5HW
KfvJekd6ZoFYMfJwIGkyRkOdtpVKOol1vQy2rFyQv/xpybj+FIoEpR3U7MnO
o7Tp70rTpqJR71BSXvlplcW/a8tociwBRmgIFBGQNKMZdSopMezyoDlnZDlI
CF2K7BY7GtzgItW45BvA6iBI8X6WBzvkDmL3dIzHG12UhBLZKqlX2saWB22M
awaWEW0YvGgotc9MEPliVahhXkAWWdvpfma9mkFfJF5nokRGIYqzsQtVIHzk
dvHpduAk3tNzM0gflxydKTu5ro8ddyPDyISaNnQHt22F6enuKaQ2bizWZc6Z
/U3Ed27YMdUdKW2cizMc/j782pIl9K/p63V/Bj1n4hDFli6GGG5Uy9Gi9l16
GOZzshgWzbjSb3jqwesi7LmajulomUwMFiXmg7pJWx1Jpce4UEQ4oHUac7NY
WSvsq9BMGROxXu7hw6onblVhONocDIzNj6wnKwDIwxCdFybkTxgY885b6eew
JIGq1IETm2q9ZXCJeokmg6+31Qh+LFgBSjWRuIlJ6kFO6CpCSIotnE+OQ5lp
U1sJUfd0W8wMHL+khj8imzhH1RAcvguCNwRRcguPdrfGIf+rts0Bhp+BK0/r
dhjz6lSYIczAe//CapHnlY36H58Iy6zLV44yE9VbeeL8bQzR+zeyvQI6ezAX
9knV12dzRbx3S3b80dr+sCr5wq4JRpzI+WJj/KIB8yeSC+BPIKAJjm5U5MjX
gLHk/4P9w4vhJudKFR6HP4Ytx4Y/6HUbD5rePZjBEFMkngl2HSCRDoDS61+b
ZJF/kMtieaDhnFN9pQCVtweXUkLecWr8eFoFcWtgl4w3u763kaStmBaxeLIH
x+R6tCOJKyOP5xr+LEhePHl6V14cXgnVH7pC2dM60O5mFT3U1SsALjQ6echw
VbkLsTpyTN5SIU0zWKkVEM4+rWQl1w4rvbxECeDJcJywZgLl3QZlByT6XRzX
Ew39xYl5m/vvM7zM0bx1rLhcaAntJ/W/4+onlPpIx80MJWAUhwK8z65Awy+6
OrMJU1sLifiCA+T69Q2qQ8vWyVR+oZo19yNzCthKzyJ+mIGWQ/nZfBu0PraB
NrnrgiM7fez2oruKyWXNRzVAEybmbmQ+z4ezBMVSdi7eOknW/zJIRC25jP4b
9e0Fj8B0uApc54sM++aGMhqFqehHDBUpW1f3ZTf3Hxotv35YQy/SH0+2vgUi
4fz5PlzroyjnK6fYdWuiFk4/lJkQcbbd9IrhbUgubgTiy9nBLNLBIlNS5RNd
Uin0Dx29sZtPx6MUiv6P0Dpe3hXjM2+kFS8/IJVvAaH0Lc1TOgfhN6Tc8O/H
DTddD8z7AvdoGeiJmGkAUsOT80Tjrw6VPQzPWwk9ZwMhdxF59ju31d2VJuZb
KUm8jd1lLkbbDNnIRUgRXg0R26B4rbby1nmgOXtVH0equI2Qh0isf0ZaS8fN
k3RfOceuFQv8iW/VQOtR/7AbFfqLdeSiprF7HMOUqRJ05CIX5OUG9P1lDBfT
wL8MQo88ah9+KJ6jNOH4pInJjBeSCCa1NiA7RhSkXfNj/lfndkzt7nG5Ay4p
+c4gTTUzunZRxxKqSpupB5WVPJvZKY7LoWz0lUsKYIqGJhCMUCA/67y7jZwZ
KSHCciZXs252Ll9Z10vApMkTnJ+hpCrmIkZ/Bjo7YXvc0B1OInr9jjSDLgAy
JLoMmZNzw0wkw0btG7UHm6h2FmPJmu+uFcnb1TdvMCGKM9ao0JDhTS/eyPKL
BRgxKlq/JtFfTOZvCXHA+fpENhM+6itE4DWWqi+cZsLFMvUX4Pt9p7VeaTwX
+3Uas8ozXo11k8dLwk+0XhpBdHTD6v5A2+3/WsJYgBjye6WMwvQgZZPeLAN8
TPsuhTeGbIXUvZVfnTafO2fCLbTzTcjezDhR8QQZUo6eWXOe0HyTQAoXNn7C
gw4LTMPjHyUW+WAdGyAefLSn6R4eUoNjh1U79/z8crHQmpFGqybnt6teE9Vj
4dg6kCUNgKUcsqJR/WpQP84EDfBb/1gkvbV8xTi+JxZEAGxy/z/wqXh0r7nv
Z+hdD7XSGdi+tmyHb/0P+AyJqiz58CxjrjafBQMtLheAb7GBpt/U28WsmTLp
uZuhuUHUmBtFtFjqRlV8DJn4CdJSFJWhu5XA+JK7o5iOxwd41bgngDc35duS
kjaEbb3GtDKmQvmqvFak4NZMDAyJZGhbGv45gTCKaQhCQaBh2fONedpOSRgc
yADxzuhOaKoSk6vp8d8hOMLiov5ICS5k1WxWL1ZnHFMvAsWc/5hgQomCpBxS
wOD6XL+92xD2Wt/aXVU4O2VSqPcfPUk1qwKytuUh21bwBBSIFCtd30SZcA70
kNJXttlRLEN4FXpbm//TcXOA/4zX1V6gkKp+A/nwXAvCLLa8FLP8FWLwaF3O
UKDsq7bsjOQ+O5QZs5RPCmtNBjZzfoOJV2i8doatfbkWA6aEnY/RU6WiDpKl
Iz2Dw8WuICktMsu5se/gIW6R7b8slUOpaPx1kqYmer3/75BUEe3xy4/bRznE
1uRyV+O1soDWxKzLoCyh1zr+cDOxC4hwy7rkdEqNFY9I9fLlOXj1ulD95MBF
HdWJ5Fq20kcsgxB23aKC0A5fJymtxleaYuHTh+ur3+IWSn8l0vTxLvVV1Wst
i8vcD1Yp42IOT1zMcw/l9e9aHLndS+4WstDo1gOZ8SJ7JHdT1j/1ZfElG3JP
q9RerfCR8lUqoWTNH5c1L1p5XuTdRni75FSIX5MJf2YqnXDmEsCFStZ4hjgw
uK3CHte1LfeKCvtPmFxZ5P8U3cWki0/iXul66bjPBzuFHrsnMQUPUE4zpVaJ
1lbNMcpNl9R9JdPUPIlohBmIwIeRAc+/i6teQckGj96RTlITkcsMgnOpXBjP
Lh2P/wJ8sDxQy/MrFTJxvJxEsFFtvnqCKg7gMj2wDawMXoyTsEcfH1rvuFrZ
qjYctco+JjrWRWxYnfblbwVDUtbx8SPl8ioGSiCyDoCzLMmtCTE2VIcvEUCG
ccSQ7C0ZpSCTMFoWiXiQwncMxQIVMqZV5TC6ka+hL/zlHV9h9L3orBH/N6up
A0FyvdjOMoLxz7goqRTmyu205MB7WbOyAliZOcJf4KHWeAxujEOZzCf2BGip
IVk0leMVdu8K8NMbvxD40veGGWWBxnetT4IyVR1Fz0vYxsvhFTsHmj9JQPwX
rfxG+yDQGkt06/BAMsX8elrMzf0La1Ljz4/GUYr7N7d4lYrPTxYPxH3w64Jn
tSTCF0RBoBcThPZApHdf7hJiuBkGo0bz3vkcGY19+0JAy73reIcIgFOyXsEv
do4M/Gn+t51NFQCTLA8NA3SxD3+7DTiyE+Cy/iigDsLElgN+X2Jh6RUZu4LA
I07eDAPIzqUHwmXcy1YK1IHIhzZQ1ChySjhPs8f1y+/nnS12hFyLMwD0cEj2
FYUNV3jdHMVX/CYaHmbPuZVyhlfHo5j4vzwromECKX4euurvCeEOezmiFI6G
HavJ92WrlbmFjO5Id0lLr+UJSghyrAsqn4U938aDqcDiaCTc8Q+z7QZPu4WQ
g5eEivStIOJhX2YGnozbpx9yiy1W2qF8am+F2WSXvl7OMvKL+sfIj2hjFCme
IZlhQRuFsA99jzTG7wTlgu/o2m/XrdDLO18l/dnTH7bT+2wWlg3rZJQVI/2x
mXZF1VwI8RRtBOkQTgxb4pdAIB3bf/asMyVDLItu708DiMX1l3R1tIWUodX8
TlunknEzUdJDTJM385LkoiaiS4KY/cv0oLZGVC8sJFDbuyuQXs+YQXttqMly
Bpwv5sDdflzZao457s2xkP20d1QbIY8n0relJjLb34uQf5AjDYdl9fd140Wi
VsVYCFSQC6zGQJEKpMovgz6PhvOX2hieOJfRqT5gcMSehA1iadBCBPEap+uv
2UqSavG8CRn0c3QLBZUTdLVCKZmkdH3rCMNnzM17u9Wm4kkmLBwyqf4RYqxj
2epD/ISQJOxgM/MrEFPF4KvJvDXhQin+29N3cryyO4gP7z9NVIyAeSBcz5WG
PYqvV+PoglKBm9NqOJB8BCGoFGtDvQe1hfGxhDZnh0lwj93zFAKtmYWKZJBU
U5WV4+0l/5kvBXJ+YhTz32Yfm4pvgVgesWIFe76PZ2wQXePqwv1MDTt2Qcr+
yx0ADdWhuHxk/BuoIc4/J+DESvdwjf1CanMODUXTmUp/lDNyS54u3AGZWSoE
8ena7aMZ1tJtiZsPAn9ZK/m5D/TxRxXl5wKQalkKahPGvWQEEIxiUrOBnQhY
7HvyrQwMojkwMJj7DEaRfkd3FW9MEAIjciGD72FA0VRDxXGT8Fjp6/VGN39q
IZcFcXwjDY72oCjGL4vFpNqe3zNaJ3/izF88mSuzNziFxA7iprtuId3Jn8eQ
m1FYlO93nKoEkiI6er9PmGIL+Aoki1hOvJ3s9Lpy2wOqtVkpd2qUM3wvmOYv
TuTwgYeQMUB1elXWEHapPp5WVjZ5FCurMjBXYFUTPvYl818FHYnC1JU23ONX
hPkSZx3cNb0b9+ZJsK44dLk8PiEw8hNC+MUFSWrc6sfi+eBeAkNwY07v+wio
+kvZJ5C02zAMSg4HbL4kIl4svtJThGEaoFllLKXtkmGqwQhCrkRTx4ygb818
HTiKLnWG4DuwbuoEZXcy4MVXLSumLbllRX1w6yVumPUdavG304Xk+qZs2/DF
p0jGaJun2CFSPjThLsJBUk8h6a13GQvp9BEKkZTnfQoqbTiXqtC7k3BIS3ww
2KuJcZ6cAwPCiRLcxCsQ7eoRKyP2dvYTSa6wn6NZMlFgOVlIBj/cSMEZ2QlX
DNOxEuO02Jb016BU85n9+wC9FbCbeKyvVsZJtIBvaWvNQ+TcDncCeX8YS+DV
VcBuIMXsZJ2KXjPH7R0a86e5bSzoRpbBRUtsbBdX28d33stW+BCw9RbOoCtj
GNWKoOyf19/cLFlapHsiwJqwvMppNQw5xsHdlEFN1Pawj9Sb++gTMnKHtC1e
dTd7cqCRmiOOTGwd7zH6ZKAq4JBd2iytJYQhuj3W65fza3hcnqgyFqg/tJom
oInU+UParXii2zAMWqXUsHMcvhbsMLFORUUHmBuHq/ugNpxbWb++XAHaA1jA
ANg+1knV6E+jZk4WlmU56s5uauTWYSXghTfel1KaUKlBP5uhbLHYPeMa8Xer
sB2q2R0k1Uncjlkm2NHv49g877d+dK74Ow6Tf2Bwsm6f/CLWAj1DLSEeBO4+
l4AcYc0D8APBvcug6F8IwVDBv39oMcAnNCi5REP7ExKR15dez68DlatVJGrq
2o3pVtNbaFjb/GZQ5uQVdmeiaHY0Afvw3QrPAurS812AbuJahskOR0RJxCTg
Ugq+nqgxeJaeTNF9HZeRqMbPbWy/dwdii4AxYNAowCc8VTZhkkFuaxETLTOt
doscE5kh0/T0AGvBiHqlDdp82kOiUsNB/VfTo+TbgoUfeOGefbrYJtGNE1r4
CSE32UARMYptMO+ILddpEsp9acfdbe5jtY8huA50Fwblicz2kn6ohIG+O0zI
5yb4OI2+qVObbgdEW6he6nqkx5AftJyXjmL54rOc6F7SrbQdGW+CzRZFsTE2
DsZwYHmqUTcjO+Ff2VcQYGvIaGMkA6b/Zp2kVKi+seWuzN6UeKSh+/2412K2
IzkW5Wco5Xtyfvytp4Lx5bTicTA/CEZct8PI7n+Z2QlAp83WpL8K0BYWNO7N
0RlxSdPwRJ/WCxtlTcc/tk+aYYeIB5qdVAxxtchWApH+kySQ+3yYc9ncHX6d
Jvs+OALZN3yVnnjwxfNUI+9B9ajW/rQ8pl1qx5iSN8ACvN8JONY1WqOtMGN5
epLRwY6L4u8xtykdvL1zpYPIQLWbnWOM6Ny4jcFex7GfpdqL0ceD8DzwE8t6
YMFR1mknY507jcfHmr0YafLx6TiQcRzr+7GRIimm0ihhAFANF7GJyvgE/L7K
hOPXI5Rv0+cPgbarJWDYuRi4WnOMZwu3viHGCad95TOFFhB3s9Axxgra4Ctg
erb0Iici7jJlCCOZJwfdz2YnJfVYE2b2S61QqdsjYzo4XeuQLKCDmz8vkz/I
3q2BbkUM/4nPScdFSXERExb2xm4w+YCg0fuCDq8QPM3VwWlwHTnlGP5JNu+w
YfQOTy72xB978DHK3XLpb/g7DVEf2uwRmN1+lJfE1EuYn8+UfXnC4ZB2kJNK
+6TuGwgA+BAiEss/uB+6G6QhdTjp5TexGtpR4MIpfwuKQyTzV99Tp9xKCX7z
33gAjsN1NpfWGuz4877nBNUg8+hcpIfImePpFDrI5TO4fAp1PfQrwPOAUw+n
p9mk8zO+wqgYBgLeh+TrNaBGUAIgEP8JCrbsgKmZUVQHbvEqkDnAeJnCeB7w
tvIl7LC9zZnSYa4arigC+dr+ccao7NtWjnFM840OSJEEbifQXHldVslnwZpP
XzAznjQj/PrGbyNSo2ASiBEd9ijwewlS2Z2yfLcx04sKRTXzqYnS/ZjaE6q1
MM76wp7KtvqhfFDZ4+ae1G19N1foN0K8ux/92Bus3aOrbQO/7N1CNlvsQu3v
TVDq3WRzVouGfwIju9lYojSEBsnViF4q43nA4OyaCH+7t8SBa1DbnWst0O9f
ndHFH96AOQe/A7/yy9zUeSfkEIex3rYcB/dbRrUkmL1fxvFPgKdip3WhFRmU
Ke97u9QHCqP9AI7S6OmanyAyJOFCVHbuL/jrF0a+EVAb+iaVeHh8r0xb3J5w
6t26icu48/yo7wedNaGY33+JzAG2w0c1Bc0texjWBClhfiu7ISLxq5yWtdcA
pYD/PllS0ffIMaJvPZQCx94kvWs0TU2qzUcj56EmyMe54UlarcncSYj6auDO
NrfTNNahGl8wggxETMKJevW3D6/x5TsU220LdS/wHY64ZYu24dT9SGxMNf05
240zEJmQ6fW9QLlg4p0z5IdRSBJUtzeuqfhG09lSFFNwocD8vAl33E6lQhqV
u9Vcab0FE87Yl3TYZdNv+vhehqB3Cy98tQAEnIJpGUqW7qYAJsiX+HE9fO8b
VqgFDohmYTugWmL6Q7VI5u7+QRKkhidHNy6DA9CXd800J2SK28oI1Z6vh8dh
5TZQ2mu6maGGIU3nnxAD+3gpLWIbPUfXp/XHL/PO9wmnIajBvxJRRzpz1Crj
RTB1yNUAweFHxQa7V4dnSElnioMZogogNEYmZqvVOTOIWQ37LCJgH88xcGu/
OPRkUuNQceJymXUKhxi8TvXg7rWaQAlVrjwbEDPddwKTx/lm03ir/fYZnuOL
5i/Fn8zK+Mu3wjs0w48Vw1W4qJjzB/d4UZ4RrfujCXI914CBnejD2PPBjoNM
+Ft7ObrmIi/buWQ/Cf0Nes49BhFatO3U/IyLv76UyIr8jgo15cCaO1RW9vBy
dKDeAMnIyIIO71dOsUQFChyNSFPA3PIUCiztAoBHxszBlCTs1d/eq7PqVXui
U7wGWKBWl+6Y2q2hkGkWwY0abRc0A1GjxXUBlHiwIqt9OLSOSR4qKI6Wb5Sy
4494wq2nSuRH2WsPDKzEZez94z0zp5S+BTwMDPBRItxfk22UquhHFD+u2QGx
q1LLaZnLq+npapSw9sIYVpcT2krt6zJNuH/pIe3+4hyI4fg2GlAbt5+ZtQe4
IZ7e8NuV0L1kq+kR5StohomwwHGyBTpTT9k/7X3LXj8U8m+UQYMHQJ9mr6zL
8jZEtXqRIBJQFC6JLFjgY8RqGZpUT/DjblX+soZHmtKMzodDaYzKTK2ppAwL
wsyk6q4iEVfogYWBuVWdefdMbC0tJXiHLGaMimJJebvaf7rf2bQNLPG0z44S
n985EOyU0OaKhW0WESdul5SUWzujJj8wAkd7r8D/0xSKxibfrsSBG4BTUVTb
5TJfvmUKMS+O0emqwOuEiKUXknrLV+0LKvK1icEed1zaSOQy1QND/l0x2rTl
MdaTL5mdbKdXtnBScu6Xdd/CaRlYQDNP/X7W+u9LrbYiDg6PFqhnyhKX6/46
glzWPgkC/NbSdpRmiRRGv9hA8fyct9hLH2UWqZ5H2gM7ZlqeJzDE0Vwh92Wk
sbwLuIVd3Ghd7mbKQYmKufWGXxOgWGD1lNoufSP5coaNUF0lkn49EmKYVw6C
q7rEwwpusj4NemVPjpw6B7kdBVbcAy1nOqQKHacL7jhmktBimZ7sNEhQ0pNx
FdFXs0KUsgGY+Gy1EI+jjpfgs8wUmk0tAbn4omqVuMgZEYrvi5oBlv8ZbqEw
x8qVrZCak2eGZ93L4WycUl/yZ+GTVZr7LoxCG0GgmE1+b6VFk6aO2+hTN29u
Dat5bhBJqR2W7uhRwbv24x8kdbVm51BGcgh4YGZpwjxiFW8JUwBlFik0e6vK
wMA3+DX9MvE6mGaM2XA7QnamYQZu/QSqdTSe5L4QQpg+1f17BMQfSZaHrTsJ
Gwx7JpinALve1A/iOvVz9o1DCb0dEaKlXdw2IOnOLQrAJk4j80mnEHVL/QDI
vSvSaYNVp0n/e/l4Q8Z6AnlpTm2jwfasuguPJClC3ChD3dMPI3tKaaO63hF/
8SiWe6cYa4n+E3IFj+Yp+20hecdnf+mFHTSgpQyau4hQJ5zbrZoUOoeWdOp0
VL5Qta+zcsnlVYhtYQ1o22GUwJOyMBSmC9jvEUCWQI4DuyroDhdUysksbzaB
+aTL+h4MaxRUEBGjdRToyX/DtUEx51b0j3qfcQNV3Q8jkt6XWIOhgOzznneC
/4kO84cNYgYfaJ21Yq8EBNWfQHMtxgwPmbo6RJRuaUX99974KeMMvhSDu+BJ
YBG1DaM2t5xVUFCVoq7c8iTuuwGjANknz7JOn1Cj/tugPjM9Sx9vHh51lMxm
+06tU+Eulx4H8+/Up4rVtCWtCBUMl8oGvJq44AZHi0stdKZcpD/c2y3mRMe2
3e2RTDcVh6A9xrSprwbqz/TDxMED0Eofz6VE5FhWjRUVpdkKR0YXdHxcg6Nu
+YwK9uTwlpq7wVp4vlIGSKImR3HAHt6Vy2rrnvu2sikSsKK0kAkA3lmAlBhV
9KNLRInUm0ZC6mt4VxqhaLlnM5vf36g61gwXA/he2SbZlqCc+hOAYn2Tvt1l
bheL5WH128lUdydSbclK1qvOhTxsUmzlO5LSWl0QhPctHsImqrZAh4qf/ACJ
dmKm2E7roQks1eqI12ieGBQjPbmqenVwWIuDhELKT9QouR8YHPZPZkzG/EpL
zloCWcAiugPcxBkqd7D2dlVBFVLHtf2MlmdH6f2U9AYUxiI+cH1U3qWuXqRA
KeVJKcl3y6IDbRy9RS5fWpAS1kli4g+iFZrcl7gvTaBQ87+ubK3LhmDIByiL
yHYuMA94sy5uYHqDDc+ZUHiHzLboezOVsWBnW9U68JkcgQl7f0Z6qQf7X3Sa
4vTYC3GA1g0Uf5keHUuZauu9AuRnxZ4CNUjq4YtJUHsT5JrU7HOyzkDk8DGk
paSK750hl1qeAR0LY5Q85u84rNT7m8He/SF5KgF04gZgg/wp1tpPm/JfA2mf
qGMe4SouJYp1oXDsd0bYHcvIopv5MQMShWwZ4543z3pMqqSnGpkx1pcu6tbQ
f6FlGTUSFdBHspVxATBMuUCQ2f5ugQ7f0JZ9qi9fHbPSfbBcddkhTJHxQXRI
TNt8EH62gmhMp8TqDwbYAGLHAvx8o6aon0pIahbwU0EvqLfyzuawRfNaZbCI
pYzpBSaJpRbTupyk7/Qx+pzaiWN3VGwJD3rDFCfxCnFiZXRAKR/bmTMMfW+N
iml1Khy+RyNWt4hTQ/Vf0JYkhHAd6oaa5QPQJbwIwDF46yc4hfJd6rrS6pTX
2h+SR0Ps4tUr1FrkmYe8rJvX5l9rwG4o2+wVj32YeoJhxZkujhG9N/+jXaxK
dFj1JbYDrjzQ4jBFWzHXVywd14StEqa8YGVu4qKpvgMEuP/TI7N/jAd+9Vte
7J6uq+8UGz4sb6DN0bshAxxxyVX/N5mxsKZsP44ALN7NodxZbMxKBOlyU2MZ
fNWMnt6dd5bsZp+Y/nTDStC6e+FfhFsWDOrOMXwgFWy6qk5kby3jVY+kJEVD
bZIMTTJPZi3cbqPNQa7vFkJggqKgwWgx6YwLGs57JEcLYd/FIH7ONnXG2Mzp
7n7UQcOK5MU6OFhDwl+RiTfSiB5R8245Vnum0PjLpOFM0ZZfCttRmK3+C6Br
Zmk4iS59WOdh0RyLsP71+BUYx7xd03K1ZzEZdrK+HNXAFznDQjeXJu+rgfx2
Lk4APvdXftwzDKB3ULr0WKdYwDYeWFJ8pTsdPanKUJ8FIX9epITdgWC6zF5e
+tgtXNQe+jv+6q4/pgTrkLS/zB3FpbGEXf7DsmyUVzxi4aHzR4FlVs4s1v9K
TAmmzwCVJfxe8q/8WOTOTjcYhYTXjtjWGSL+70MsHNEmgocHnUudAmQG6Bix
ndWnJiS3SKsj0dMTN/guy8jZT3IXYMNu+PBFZNBAiCPDhRS631TqHE+x+JkT
bkf4neD3RvGoH8X7nCBYsTnNzMp6sgPqEH5CNTpX5cvdD0IHGNHapmKkj/l7
KaPPA0iz+6Y9J3DYFVvooZnaK3ePNsfIn62n0zJD3L+/OAxmIoIbbhgd4Idt
5d83xgL7m7rfZWEY32xs8WqDIerps4XN8XHZ1bSkK3LJTbEP9dra/ULVhZ7F
rkupFIFx0ZxnQF7M5DQzHRZ/rlaSRnkTUcYFDLiMxBpcwTE2NrnL0++4imXM
/n9jWECuekTShmXIHokH0MAnmyWNx6Ad4YWQERXX2iszwF+U3PozBvLnsf4R
37tvIKn1fXBtl8Q5RH6YDUic5VmJZ2wcQVaiYF9fgLWJwHCIThIEjmPftPEm
NEtuDkBLeJ39IdOHgEB+QZNrVEfdsquF1ik2+tTRupA/UdILmoqFI8pmz6eA
hguENbZS/hx9W3AS7yQ0SmAN8Ts/EKe7dJYhOk8wcA43V0uXgsAPLcbmA+Hw
OewTUwjILN9vRDGP7bnt8h5zzbKebYrro4MRtP0ovbxawWoVCIEqnNArlOqg
QkMKHZZIxvrPuj+bwIq1I301QoCyRaBYHDc1TPVQCFo73T+tYs5XkY9Twan6
iC/Du79tbw4DS909cCnL3hTGJ2fvqsxNoLBr1c53B5xCLNb7gk3PCweQHvN5
JtXkmcnAvrPCVdBqlytNJdqGqKXf7WhnMwXXh7dg/kWhindioCq1pLbbKR3N
k/wp/xnsKvD+43tSG40c35NB/M3WGM3BeH1HpBp0sXDCtZYASQymOh/ms20c
pERKyOiz9xrQfFBc35ZKss9pUEe0p8mxzM0tM2eyr7snSAXjiwmoh/0pQsi2
9MDcKo7E22X4lDItpg4sXqdy85GZjNWKYfJVy/mbuyi7NvyXeMKakMr0S3MM
tPK5QHnOZFIEK5hvjc5NGb9xkI6VTgT9k9QGbduiP1y2aLle+88jKvS2+cOB
IMzHiX3YEnoGuiUqddxbh8DeWv6uVxXSr8ILH0GT1qUF8JFNHYI51aSUJffP
xL1YjALnPmtScSPu3oreIFSPzGm4CfD2TDdLaZLLmzhnXApuuY4t2GR0so/9
MN4kNo/i+RPYI5rEV2KzWOioFZzbDkkzNuNtkH22Sr7IZtdAjEnzpPD5Ew32
NJXqyIbKWAghXksoiVPL12mvithnzO2PABz3rsWYhhD0BKuYexyBr1QRIguA
ZRYUqobyM1yZFGVAOotXsvMQJNlsylnuS0mUY+SrbIkuv5AVuT4hVWhatNaM
58S2Qnxbd4r37326LOfVdBumX8fS6eklRUVQ2hI8nwkJ1LBFJ496eKjxMx2d
yV8wTu/fxx3QUSrdtAHdFqKhPFmoi5bFVVdhOFmhKPS9feeRyipgqKDVlgBR
668Bxjn00CMm1JHWBVoAXQMYVkzqSSIjZsfK13dkp/BMLAkqQOG66AUs8g3M
HTyA17Hf7OClKtPahzKkiTyBJ2YT8+aj4C3Fq7F9P/EdFNMHeJZT7G/o3sps
FvgLLaOga+4iCsvayB5Gr7/TtETuY+KmaCysQb/Z0toc5YZLe8l632Wu+wkc
DIfMQKuY57t1VzSoiRdxeFAfe3GgnNO9y5FrhclEToChvKp/FnUtJrdFVMjk
IciwhU66nGzT2uiMYoeCkLV+0fevXSzyCfYMHya5gpo/J2al3qilmYFxuv4k
CfRjCdkBz2rLeWqx7UBXmS0DNaysFU6lPzd7nk/wd8xRQrzlJ1Li9dONN34V
U2uTVe4pJIYbhvQCQmn3FAzWEL0CCcMYC/mOJo7D/E5QAvLjCMAz8i9rjfNG
adzuCFb0dBSYZlk4eVMUjqWGBs+XaqS8P+6TFPhVgaKmJuaCb0SABU1wxxQr
XN2igfXf3i/5K3oZ7yTmOwZYni9P5VQGxMuDSmr2Mh2k15oZFo1MiFKNcYhO
/9CK2ThgL39iINRvcAuoyahDmZgilaNYnkoVVWLRxfvWO9FPvWljWNEKauvK
flRXtj/srneKe8hicf9vNlQ2y8kKK53p16BbNI+w9T63PC5rewEKOzkjrIeb
ySXfBVxv13m54790T6I5hwqrOEbGYQUpKBirR2MHFtIEGy8Jhx/oMfHLOAY2
16ChFYtN8qMasS6AwOs/yWj2nGY3dTucR9SXOofAGpH2vOMwKFqyBcpgUop2
tmOIxtQeE4XG3GaG882VRJGTGtTJj7TA4dzfCIgI7dG/fs/W7jZKhTHjDSV1
EzopA30pgd0dP0y1btgmkhynoN0BTHYS4XpyZnl/3lfV/ytU5EPE34OmFTbv
kY0OhCiAMSeg3acQJdsyYAiuqcejbo1jaLei8gzBcAd8row3Cm6UTL7ow3m2
zpZVzNO9r1DmCrBhegZVmoYqHwz9jNHGRw8i3Yb32RD36E6zEBZp50v0KZgr
cK9TrZnDLO8qFKQGLvW9UK1u0es2yvu2yuVvmh6tjzDBgvOQ0JsW8VfzIqQu
Bvvlkj5UWg8nkel+NSppvs9epW+UMlEodN3LlIAyLje07Mzt77ifsL8xlnQz
71sHfcLbIkwCKH3S95PPgOXVNGZV+8RSvLrzkj8FPGPZoa3Bd+l2lUZlIfpb
AACNEKCBkzazJX7dT1h/WoCWNoZl4ZWPszQw2A7un7HvkrDXTpFw+UnbnGFx
cHvthCU7GSD31Dmj6PsoLFb3+mTAVdbunA6sGCI1CKAp2dxeO3AKELPlo0Ik
dlR1XeYuWNCYznIhx7q/z+HZKMczHUpCWNZ78lpASjt8N5qXCEf57NcXZSig
Ntt6QqdsbxbNTlaejB6n0Nor8ZmjS+QX7cLq4Nbe1PNVGdlBJXjNFLnC0dt5
ZOrUAUek7cjOwrAtnH2uRwiP3NyZbbM2bmlRB35XhqFCGApTm0mcyrumWMWv
MPd5Ko6rBhqW8gi66lQce2ZxehDpZS7CYKCrhsm1kR0N2xLLLTT5O2U64v3f
zUEuV6LQRd6+B+0ziPWBG2oTsj1ZZ0uv/V4hBCyY0o004VWNlWW+kFbmryip
+osc4zbCn5Xzzj3LDTMJekMSGv0AofEBcOBJEEJ2/DdKa+50K3RlFz2F1/np
KIxL8lgEUh0bB/1eebe4cTv1CzZTQ7JJyL/DPNwjJoFgzNcf4tVgTnksydRs
G/cXqT29aJfKbWWs6+MZB2Sj4srwsdCehW56oCYyTQW3Wma/+AlxfrIri7XS
dg6gL8Abr0c/0UhIP6eHqbni0eHt/4jSfrH2+6Kl2bPW+PLjvxv3Xwfy0A2I
XGWBqKj+6lHVGFlXI8bTjv9k6M5Q+cKMe9zX0RpKTbSj5g65Vz9dY4EV2WYn
Qxx+1AANHnz0+MWjcvPEv1DendFZhmCsbemrO65JLBbt2eA+rQeMLzkbEbyY
ZvaCQmq0H8En/Sk5so6lMWINdX5M4cBDAarqMVCBK83DCBiGuZtjmQT/4GIs
W8Pta5ddeDwILBG3NYif0iwWy+WFfZmyIFuh7E33UsrCgPzOl0xeXCjQZC+r
JqZDVKdHx2xf6UWXdmJZBrvN5uLqNxrDLpCfxtl1Jbc0X6c5TWk0l268IHfL
YNSy/MRUTtjed4vUzMStq1xeBF3MLUkZux2O/ZDs4jRqIaNJ6E9R3guOi8O6
Gd7fW5jAZf4vhCyXSb/zcMtdTufPq/g9knetVqJlaEbwFQLevzkWjtIHSmgK
AlfxlY2mSJy7qtKPvMedgttdJQLSY4ohgZszfj0/37FiPiBQmNvmoy0DXh0c
v00b9K2t8Bi/0/REsanRSSSwKufvcSl6FRT7uAanbGIQyAcX0RUPhlThcFsM
LqYkjeS5c6hoQQTVuBkBOyd+pPJ8vp9hie9hvOkveYriTWi2m92P53V6WS8J
E6+QtlXYlZTtjz8o4GeXtcwt96EbFcbufizT5K8Rk6H/XVrnpa9v3tUvbkwR
iolp9V165F1jnYfZKB0NDYBggCZD76rJiwOPOND/5hCFG38KW42n/bSMNLHV
Fk6BG6CZeLw6vcpBdUDeFV1i82wt8w4Sym4BNslYw0GlH0szOer9fZWNxY12
CaN06+aVqET/9WPS8r2XqDQEuccC+sIBlNGirw7gIY6hvMJcDYSL0TkpKtHo
p4pwoQEw2brtmJ5OQh/PqPmjZOwGG1vZUvD+MX3odFMfbqCx04svcvuBPyaD
Aem1QclMJmTuNv7SiHNysbai+aJArYd/Fs/fIAo1w/q/w7vT7C4Vx5l+mgxx
42wYbmP6k9XGU4qV5urjizb36RGJdZPoE49xZrwd1IcvWe2SoUzwXsaaQ3q8
LNsD/ofYhz445z0GbLlwpmzEz+ma1DYZ+ebLGQrQinntHpA7CslX450n5hZi
/6XABlvjO9KRL3NI0HmxuE43QpzRKbuFcbuV+5col/2ipBUKuuhdSnZf1u4M
5ksWyI4N862sDJE/FBVHfCB/7kdU+s7/R+HTNiXDunZSUwaAdBAuDTCTBY0A
IxAFrvujv2eqxy919GJ1iP2Ixs6mjfLGivweVbJrE2BiPkstFbVYy8YV6fNs
kbnb7KbXTIx1It5tou3xvM6i6jAvqr+ZqPXCZGZp1N/0V8edT+znPrsuh80h
4H/6jpK8CT4sE8jmxjwm4AqTFPQ/r4wLo/MhuFrxK1u2Z11/ezjtWgXvr7OR
uA/c9OzAM5ijbUZRIvDr9aJ5f0ZUFADYvjVSbnoF9FjRs80WErBGqHvQs437
aHxsC7OimDTPQQnoue9Wo1Otev7XeckhEITU9Iv1qvzBBTFM54VEWfIKsF1C
izXQQfs4PGvoNVnmWnPloB/w+fzXvgAH01ztBHFdHLxGjIzNUfJycAHjjQ6m
UwxL32D95dK1Gd1pOkfR8VsW8cM2MvGO58Ygz9rnb9tMFrW0V8xnAVuf2P+e
Jzwmfg1MRJFM74cWNjQRS9YtSIU6Cz56ctKl8bXfKgMA1Kd/S4osxWnFM2lB
/AmBfpjEymFzcHz3HZaNXIYlnz0Sz5AalgISH9KpMqOgq6M+ulMRCg2csNno
FNjA14DfnJVgkANbM4GbMjSSmu5ieLLd+Ad1e6l0t4LaEYxSGhJ4ybJg8Nb3
z1DKl4JYwJ6LfyCzJ4oDEhB27Zz77SHVMVnezZWmfupGomUfFrV518q4o/rp
yQje0Ci91LsMqcB3MeBAI1jveuteQFLXPYsj2CbIQmcspL2eU0oNs1tTgvXw
nRVtmiZ1exxKMKN0ezNLBKiGulZRoOSoL2rqwcpn2jkA2Ciih2wcyB5v8FLu
8h5NNuiHxnJvMvbUD23mYiqbHzrizBSziJV3swSxqIzpcRmlgroTnZAVqBep
b5jGjX0Rv5FcY0BX1dn8e5D5C9AyCtfEMaZPZMd+SjeOewct6N56Bok7Sd3n
nhBVVpfrsygzWxG64hFt+/CAo1RjytRgO0XD2iCW2vLVhUhkkO2mm2oGW6+o
ZDOFrutQFikHxoEnpHV9PqxwJnsmN+TKG+nOuMDtX++UUj9NywcOilC5Ypd/
vDHmVmc0MeSwIfFOeyzPF3xSvo6BIVyKb9uausJpUdvEyKeoPKng/2tD/Vav
APV+Gsw80fAtfSEQLZlJ0gGRK1VTGOm6XbHb3u/JGb5akfVXVapQTAF31qy5
rKfof4egHp11tFKYPjCT9mEDRKHGIBG5la9WJ+JDzc4CHgtsAlo24N45cSHa
x+wWKC/8SIUQbcJME9DUc7MQSf09Lm2sitiORoKnpoboCGnsTYWRzKCRLDPw
ikEhrOlkYx/3I3qLqaWzjiOt7uBeGzavatvBmrhc71UTToqR0rNyxsScONaA
/R+rXn1YPvAWegobMj7FQyHRY42K/AkUH3QBI2CVhCK8MBDzdpXwXgZsuJF7
TT1Zea9CnQcZZMZr94bQo3cKGL3HdQsi3Q0jB4tvjk6Vqc81qtFuXE3zuy1E
MS7XAdMjAuVhOTo2FxsCysL/jo47I3vz5pqGneawwZUeAEKw2HOUUQJ1dTsb
Up9QkYEFO+NNJaGIHMbEX55Nh90AaUO8EcY3331SjJFEMxF7lpaQaFMpI7sg
9WMEJoqiTx8L3ikdMtL0dkAVkj6nTyYc7crdqsJrBkdGBEfIN56EeAC24Lox
lvNP3dusiS179C2eHcd5zMT5IjnLDtbf+Xn1drzlSZu8+nBBnVUdAaj0+8Wu
vDFG1WQDY67KA5OR1h5tiAy5emWa68uSbvrBgeyf6Im1guad2AgNWkkEDyTS
z32BSjNjUg90btqJ7buc4N/opGuDzLWXAynj4nAH28jb4Rri57supZGgWrcN
9UntVOKSttEPI2E1ahBcgwwj5VwkjPrCD5pKV2rUbiDdpHA7wMBBWXd0TRaH
AuvtmA3yDtgy4kbOb7+2/XNfwELNXlPKfZfFLE7Zfpci/5HA9Mh4tFowM2W0
ANbwNCSEmDBF+IIWbFeJZZ5vAN22ks6pDDE17ZUolM1qJ98RrcC5W37ADw7Y
DJPUYyqw7ovOvFAGaUG3REk5n7NJ7bBDzzXsNk6w4Vq3rTxWT2SpOlJba97N
XlB+/ePkuuUZs971sCDJKuZAXzz5dOqN79wbSLC0VvndO4RBhnneAnwBHlIH
kCxtqiTFeVEy22jBMZyxZXjJ6y2fLV6RK7lTuLqhhTX9Ngfv4sL3KhuK6HvP
H4m2zclGGnCnQSvr8cEUvYNnc4h1DEs5ymWktRjVVg88PUjvnX0oPekti2xV
S2+dx9y1zNXi1aBKO/NmzRxZNXffVKNFZdAtE6RNKF8jzaDSRkSskunkdtgi
0gDvpWK3QtCX7F9Jov9jD61arzs4K7Atbowpa31xwEDcAP/BcGv058ZsKBx+
9FGwCxCTp920xRDW3y9BHeE5L20xmt5sef3caIbmZ6XXpXGpUtH/OeC0y4HI
WjlDxbWKYjoPkGQMrdaiL5cjEPFgZ5SrDpMJuqjAtMfeHgFtG5nNC2A5R/jt
RnZzgfpuhQnIiK2MPDteLiOpQSGNpRdwI8S8nCe6BB1tlDWqUa9Ob/snjjod
HV9R7eTvyi23gY/TgmPrIzFWoBv/EL2eJuLLEBBXTuS6sqgA5ts2d7Dq7lVi
BK/QuNDysH/IGILEDqPt51AfNq9dvJiRxRSbYFbvM76ZrVXUcoJVfyEUFENO
7BWgUAcCeuZ7G5psNS2IZlQh9eSw8rPjYIGdSZnCvjCftTd5cvDjtGJIi5pz
5IX0TLMWYCKyu5QZwrNZIbpxNMKPbZKNUcBPUT7xVNKO5+3DZNLlnpnwi1JS
0eF/vAjhi3t7T8c9tZQQnhf+4HQEl6EsjWA4gOISkHY4JlMVFt4rEJ4LICav
wqc8XxrbPqezC/lgdeC1tepGllIJL96zlOxjNaomQRIDM5Zi5pw+E7pcPLKJ
hDz6sbd6b48+/2ONHkxZ4gt9tTS2xFp9B7eYqZoCv/CyrG+DJ5XRWDYpoc7D
Zsm09XuTHADYfpokYVtaOFgaIL0ttrN+dLBDs4HoNuOA1ZB/1YbtGDiNfdwL
vTZhHWGtG+xeUg12jdnPMdifcdGfoj148FyPlewtgrka85Czfncibggd5c1r
19Qu1trKD43BNmGDJpuDXWLwmyQNpM3BeBvkRrtrMMXGz+PBj01ff7sc/EsE
bQHf059+b62z3zb04uayUnPzqarfqQtIgdAYwQ4Y8j31RJt/6+7fiD4bGszX
b4KYPYO+d9TjwA6AKsTk1vZlS/+XY4qI2KcvzknTYGSoEc9HTzBcxzzevH2M
a+rOgSMtBCv0FDXDxNQZpDorMZeDi+8J4Wvdz106WQJTECFnpYXn2lbk8FG/
GMKTpNksiJtxQKayVY1+77owJGVhtgiljDFeuXY7GdHwwdGErXUFWzc4Zq7T
Vven+B35MbLewD2L0rIafH+YlmN9/J7MmOpvammQq+OeVGe0KMCDneAC6Lkb
6QE3HlHp99xlKUYcfhqpR/Xjnhpd6a1QMo1WsT9qao1306KNZK2xbbKevmfr
tMAgDY02jervYPtQua8jcao3g6jw8kvMBrZhJzf8G5H4gislAgoRBBJip3cx
jFpXc9YkaAjmXJRmaWvs+goFP8qj8Y8hnXz9XVf5Yq197vxQs5wIaH0r1/iS
wWJFVqFAFz4aqjjJ+QaX+0EEnl2A2nAvoxIFB/ELDhbZkxv1jz8Ozz6N0UtJ
XB4Hg5sJX23W/Qdd5YdpE/kEn0D+gawgmf9aixEgOQ3jL0BSHWfF0GfDkSzo
lYtJbOAR3ts/kU4oBML1vSqMn8I5FgwfnL/zCcMNmSYHCQgRBY/kpGy/eDmk
7fyqQgZ7hDN/Eg5tt30U/VJbq5gLAdPoliQ+bd1HeI3JbG08fioD1Q9IJKZr
hgOY1ke78m1u+njEvuNDuRKrijh2DBaqCIPRri9xhnxzP5joqGCt8SFFbOc9
rCC2BSlq+F1vc/DPDNHav1leuhyyvm4q01SH438w9bzSVgP9htkJVZN/MIRk
LrK1XbawW1sgZlU93dhYzBIEvWukFkW+VZDUPbW6kpXzuWs6sI3Bf2aRpsqw
Xldp0eDVgACJn9IRWsjQRjK4FBxqxUPN2jbtDGnLpufk516fsJXIa5aePe64
ndVmNbyRM8aOtTdhZYwVw4pzvOzqifcY5Rv8Y+1QO19ZzBeTRmEKVElHTtO1
hG/hRLFkOsbSS5r65vC2P8qzS8T8xo7hs1ULUTQHeCbSLkXFHejqZu2ozB7h
NAPiq+ne04ggQa0QuvYe0xEidH5vHECz2pYQp0jLOGiVlli3PKrEZFiUqQVe
WEP3qasGmqQxwtN7jPVu/fx8wHoT4Asp5kGIYvhl03c7W1GA04r3u799GU2R
TsQ7uQoWwcfWwpo0EWyT+eF/9ouEcJBQzNAfNF4ha6tmIMkmhiKRq01Fxcg1
3DkiORAG5bMEBtAJzm1dy334g6h/3qYTZP0J6dCOjIMPdDo95SsCYFVt+lPt
1uJwIgZJFrXEMBjuwxUoDaoOGNxn9TegbiYaJCdik9biChDMZxwx4mNzeGBn
7PtU/yqVaVENG9HCMfOHVQu7uCZ8hc8esXqNTZRhLbEHev0kE7pJVy0OCXEn
dF9Mctn1HPXrBMpYAKpo57DeEQa8fh+0mXnfFHPmw97A7nCQI41EgnY3BuVX
rXZ1TWe/7QSTuKxH+0+zTF+jgD5VG41JYy3sPrUPeN3w9NYLxLL7A+PKzvfp
oThVSnzzQS1hSpvP7SPp1+qFoJ7mL+axK94/c/QgHatE/MWIyladKG3W7bwL
Nb8r9hv1/J1fT9vdyD4ISO0xraeegzCoPMLpseikACgwCi83dryvrDnU9l62
KPbshns+MtIhjvhZ2PlRj/x7EAsSxaL9n9xp2D5xdeP7lgCzMwGQw5tpLvjU
zM93TBktdEo1y7GrrqO60C87uD7OtaH4xMSpkujG7cQMfjvCxAWfLZyq82bf
cNB4dygqOy8Ckghj+H6H4eJ1+yvPra9Vj73kHI2ZP5q2qEBGjSgxGQc31X/f
nnmg4qENvIO4/Zwg6/MPQutIXT2TYKvyQVi32LHBNBmCpqM4j+lpv0hisP+T
wJyjU0xUC82KsR+HeZB9vpSx5ZmWb5CnZuxy5wCens4/P0kywEMb+IiWqBAN
iOy85HsW+UPA7HLUL3pQRbahrZv37efVTaxNKkaFqmTzCTibWPBRtWz1Dki3
SAX9mP2Oe7uVsNcsD66qqCs0F9wXgYtGGSMiBvSchX3yzLYRTOQ9nBk4VkvK
+O8Q5VxE3NRfvTIBKujthZzFieinFptzGsWQBMHsKThpWuWmrGo049RcVTMb
6VQcpHGLyv9RYejUPjU9Z+KJksbdLngUdj9DFApYmRQ/aZeXXjKQaK+xtNTk
FDxriVXp+c8rrIPrN+Z6row2hWQfwLYJy6FSk1Qw64YNgUelnKzRzOWytwFF
oEkEG2Iesn1sNIGUGmTDd1ZzbJb1txNaovp0+qFRJ5sWB3TiPyALUS7sNylk
48i9h6hGEkFwhFhIzGV6pZxT642ihRGIUmcmeIRsEdnLzICjq9vuqx3NbYew
nQ09sBHH4Q4v7hwXK01ijFISx3uTbSUzM/75eqFsK7oUkeC4y9nGaC3TO6fR
LhghkTmeHVtwo9ZtX6iv/cR8ZVL04lAPMmMmDGsZLGW+esTJ3d/xwdao87hU
nP2J+vh0aHXau3fDSPPHIjW9M7eZOB0eIz9XN9Iud9hGy0oRU2cErPmiSDue
JBhMUZ9+lUEOCZ3DkXv02c+TBghhGLU4Hw4wgfZFWpTcjhbQBC90BiS3QlOZ
EsjY9q9kYxKWxaeVR6SNqVAJLl2+zV2ErZx4lneIFlRn1lfGgaTZXM8Go20w
WPznE+8rADLaGbu/xCKXkw8uG3EIESOSBuO7qE+Stn9BNdGcNvifdnWVxlNB
P0l+bakuNk2xRjZJoSyO5ob7UfT1GKzqV+5tnhsN94skzvG/I0gVqs979sZ4
7+/Pbi2ppDPPn6Y2JH/XaDyv6cE25v5hRquo4c0HSjbqFdx7VGErLF0NONSr
iFhSQ/CYwANZCmmDHZuukQ7chkBTbFMC8pwx+tebz6BTS2rP0ZsofzENoMki
a9Rv9ncJ5qzXBrgv75mSQKCiraGFmA+1xIPSCiaa1CCxJFr6fWD8IExVv0u2
ZcsWP/gXzf196O8Ku3ocCfkET9LdW7+0gGkzeqcuAECqapZVu6NQb5HS6uHE
bfMFqhndBeh/v426qh6rErzSxccZuWHv8zojxcbOdEBwsZWVWaABEMjImkqd
nXv0g/uIn0BlFZaFwrEa6XLqZuxveKCcmasW9NuptVA2A3nSEgwJH/c9A760
Jbjs0QbrJA+I38AOr5IRJObTE6CxdfYF1QBAbAH4Uec/X01zxYbBwIuTfmx1
99TyKYa0T5Kg5MfhCKg3xRy4/mwwUHqV7hPjbDp9f2Is4Ah+Bf528QEOVjhN
Z9msMKdqJQ2aSEPm1ArugqLiupRpVu/h+iZW+8S89joPYAyvvBnTp23pflWb
GnnU5CJkiruzGNz7LtZF+iSXVziCwjOBcclJNShYNZqWTxKl8itXqe1N1C7v
KjwO3jtUIR/FT1gZfh89qWQH1+h43uE3jk6fhlebjd8NUkUYjcgsUxXBXszd
m7s3yUPuVZDlXLMp/XjMaX4aGMOBFIb3zS8noA5bNNlB39M9Ll1TENUJhG97
SFJnkh8wzouERutuOUQ/dYO8TNs82DXjR0yfOfgzxBCyWi4CsV/78DnrAeZs
rnsgMEzgwvmOm9cxMlB6ToCtOFX4mKBCVq0lsUwIdv8m0C2jg5CYW0oIqrJz
/Rr3rs5ap5qQFEJS0IFu674VyuP/2QJDRvuCEpKGFwMPC7Sqfga4pghGtinq
7gYtqAe19DKZutxh1IZ3DaNBB4ctgQ3tGPjI7Xo3ARgimkVaCxvjNhhQF1WF
4ILPy6xjmYkPif6oi4t54W1H+j6F2qjNn3GxV7BblE562Wa0KdxSmmy6ZUr6
dFvt1HR+IlFuKAu21uPcdycI5Q7mA3DCGDoh1QrGiqOly2ATvIF967311lOa
dyMjdF0Yv9C15wEV8GlyINHw82aQlrQT+9f/NwxGDFKOha53QAaGh1bAVOQX
zJGHpreTzV0MXgw9nvv8ndLP4Z65UwmpqnHTYWgHS8InUJsxIJQhRton2t+P
vRlYYFVGcsNPvunKDUnYJhHNAAjmKMETr0CfhqHGFtS5P8BRD4NXDIIhqIBr
AV8Zuw5AYH5f201yHYtsJbqAw+Mw+Vsi0JxPPEgJBtMFjcP8Ek6k8wpAQhwQ
cC3K06s2bjhA6ahal1Ml4PsPKp1d7pzwsLutdITMtwo/+GhqmId28a/1H9vk
U9WI+sRmnWUkAankcmQ0A+ZbjCeVg7iS1nAKPs2iqH7D5LNFfn12kFxA28Ca
YwPT7Yn0MSIcol+K2dfF9C9wuVOSpuA3Rkh6rLY2MS/K+RV8p2sBQbRiaMOs
bxgcb8u8QIE1sCnGfsWUdrVp5DdvAwsEWV6df+mTkwtKvGGAkGCfm/mrQXHR
ap+hwGndxNF1Q8a2ox/24qDWBcXFk4ysGcNrGZ1uTtFTiQ+muQLqH0yNQU7Y
KwlNmsghGnQeEDVrUk+XRHeHnU4deP7k0qLhB41ZMfBOLYESrMaxB+Hqcwt5
kzeYWzdNDskJe/Y9diTNLq5osP3BkvYYrzr98fNBMC1c5Cc2GmT/rxeEjjAY
uYPnuAD3cCQVrcogFleZX1JVA+nDgPow7tky07Gb7kzrEFzY2vcTfeNt2eSK
Cr8voq0dyIe5MQhl7pC27R5H+wWusqjq/+qS95njgIqRwpy0A0FR5ZfJAGl4
1A78YOKeR6NUQgbX7yKQZ67SMDP0nMKkw/icYaXwSJWMcNLjd94MbL4rEyUC
MI0JWx4IGDuxldmGmvaGla/XxL1zc3jeEZrEmCXX629HK9ztrF4utfDHjxSF
bQ5sw7XDW55A+oZOfZRmNLx7s4L0nKarPoz9NDunQkeBLtkpdRdpXoRPI0oj
mSzxWPxnVFK8MnTYE3WXMW5aqnsS3CdZBkQlYlTDYUWkoaIiF87ExZKBVJ4/
lkjP9G67d9Tc2lHj+QooQEkZCt23FaPilONu0fiWeDdtvP22OFW6gcVx6irf
Gxaf+0ILW2g/6X9ERfeKU2WuseZ8vP0BqYi09IvIFojFQbwtERZtInNw2sRf
hL1yLU0lB1RsblLVOlvlcjYTP3f/nYBrXmYBDbkchxne1VtTs9xPTs+rxnwg
3kOqJExksHHl8zTznHx0ITalUHrnH2jusAKdti+PZaqvR4iTlaupcPbPeHgQ
lzIhBGjFqw7GjUBQWGoCycfUWWqxbFu4vgmocDkhso/vZovY9EQYK5E2Eovr
AfwqhPn3I3WlH6COIQNM/jVgBrZe+FmyG9wTvtWAckgvTuj1DOJDUg3Dl+0h
VVC7tvzkdi+/ni5iZzuQDu9p6/to92KKgMDS4VzruNqF4UVENZYGLyxd6egw
FqzmImwDGzdnWNmArEm6NzTWPvjIAcQtZZBTqLtKHOzsRyNJJv6itT7+qcJC
m1sp4bkJfONKCIbmSFilTQ0R7/uCkjZuZej36SR84dEEcoFypQDK28HXRHEJ
3B5GY4RC+5mH+LnphYBI2D8gRpkeMdK72k2wXGG5R1sGnEHu5u8V6YHetD1l
iXumiJsfwC9yTNGenXvvs46VEddJhYt2gpceXli+T6rzIjbQoVKEaMtcFg5p
fmqigSu1l30NueuecYZlRdeUYFtz0wpr5YnZnktMarHlZXEynMd1ppzQwY1a
lLkJHH2vGpMHoDC6SOaXSFaMkP1M0VqlyMny2kXbDwhyvoRq9lmZkWRkY+Qy
hHN/dPwsiBnh6Ufg1Yr8BmARKKcwc6LKFcxM104e+lQZ1Is+LttgvglEN+Pj
uAvk9RcVAZ28uB4567RTjR7Q+K3QvIuy36AWxoePx+mBu6sN3CD6lTFVYKa2
Yy9zIl2gbKV5YsI/bK81je01ioSlJ7LQv5mSUkqgm+Jp2+sN7byuyXyBzC9i
aqOATdeRPDw+CSlrn6lc0kF0KjLOIxjC6oY9Ks8//lyxchauJNBlOwx1yGUz
94/uMPGB26sk0s5Fv+OgMRYv5fgFcER1op27Y3prJrSzYdj18VD0rDpcbk33
7HtBler+W8RzhZiwkJ4b43c1H/MFUhwSPThmoKwjsNyQLV2atvK8iNIn6J62
F/Y0oX2+iuXQpTXy7o9NpoeWEk2zhOz1yk2hg+e2kXJje1nLNSR7JEnV2xft
hzpGv6tU56XJQoDOqPFe5jHObTm5beDmVC37XQtmfJ9HN4xY5iOYayRnDLtd
zjybM1AjEm5L90yxKsbkSbXzLKCyII+mJ7OKMWgyI3EBUz9xadyJ8GJkgLYw
FUl2W9dBvHhVH41G1F/CQuLr/N2Xc0qKw7j3DYfwBR/qGF5BCSvmtOdhKmts
wDKGrPEyb/20gN/NGpZBaMNS3VyrKNc59zTQ9OhHOCzZejZnkhj+PbCjhsq+
EH3geNijTyn8LnGfw2dpvWFBjK1T2abO6EzIOEYvYv0a0E/hFatz3OzcaCxK
dU//KpMf4NLyZhXbvPAjga3F6ixF4tyRROv0QhsPe4EDfpx4D9GC0X+ktdoD
RzwGB/tc9nN/dDXU/5rONBeelSBykICtzPwrWoH2/2+bACJmrx1OrCXzOEwO
aifqRCwGnw6mz1iBGfeQu/Q1hTgQ1UbnyC76blBFlztZpIsS3ri1uAAut5df
ey7qnwE+RNciSE1x7JgfdeYzolRShla7nS+PxPSUTRxXygzERnpnYKGK5oAh
27oG+Go5Lbe7/Y/3mAhPtnnH1dYS/ZbiGd/B8cdP6wH4Yvz3DibsuLOv30Gs
mPiwpz1Q6sKTKwBrhbTZlKA1KPNrJZvkqGr8y+/+psXnumarUyxtUPcnYKh9
ydNTiVwbc/fOJ1zMo+89s8v4JNWhvD661PsvO6YYyBjqeJ3yxpHTpTet0KHT
xUSpR97k50GTaZ+KhngM5LzXrc++Hb38l5CYSkvWT3Ktkdm2CErQ3gSzVOlT
2F1x/bqiQj0Ae7b2hfgHICmWNmFN2YVU/WvJNa7AtpRhym5D02NQBKgSYioY
T9hcUZiyWErHG496fENNm7AQgPtWhOllenjDSSSO3Ym6QOVb5Af7tXNh5eto
ntsXxT3Y5E6YN6k1I7dbaKsaZ1Iz6dr1ZFCxjYQ0sRGxbP55AKzsv8wIkrRL
RLeHRfOfSk+c85QXLpjUt5pPAYC6uDva78/ZMbFv0eS8mdlJKQk50FfCG9bE
15+A1rJaJBLV946onhfqqp4hAZhqNz1bXG1OQMhoIly9p9A2OqVHvIVD4Ks6
+mAdYieUBR4ufY4f/5eCTx66FGXvfmpmOOyINldvsgdweUL+IEvEqBYob4yc
uB2Eit/Q2OhxnMusNTrunjdelv0q7OUj0LxoK0JjpXvt3gqrKDuHGqt1y+yh
N+Oyk5qoZ2tKzHinyxaIjtGJS/jbs9KG6Z1J4vFK3GmrzHRr7s0LDGKvYpCt
wPQ1eKbI8e47TBw5z7GCps8gqPzhXjLx/qwx18WI7u5aPc5anSc91jS6crpU
73NChWJ655w0J9hROXVjon5RoVm5VJycKxPUdiwZzR66PKdzJE1UgrqFGLRm
dwp/B/13hI8XRZhNP1lv3TUB2M8lJQmuD455+zd1A12pgWPcoACotRBZyMAr
tWlIhtAmwtzUPl6d9YMdHgPUiYZVyvFZLIuIT3szFgXgrK6IpN9hXdBRDuY2
7nvIKckGrdXBeMw4ZerDHCEZaK4i7/wJghz/VxqP95SX/L2BPtl3sshFeAsq
XKJtcTfBgzR0nCnUXMM+aq3xSIqq29pO3mqDL/UZiNX7FR9OJhKxKUffKWXX
6Z0HFdbcX6AKvZGgeHgdd/RMvY603ii/Q1aF2GHikcfdiJjUO5+pPyjHPpgF
O6b1mT/BMx82QgrEqozin8HOzlU2TBTn0u1zMxsJcR4pMRt9Rf5GPVN0HCVZ
UbCbAxNiIxOmRhSJQ+0+KOiOA7C1p0lGX89XVAo0X6abLaurb78hds8ZieFr
IWpXHve1elmVq63h5P+GL9mhEiynAmM11ttD3hIWCtp4GJbq9wOgQr2mSIvz
K8UD9wiMbHnSgvLZ4lRbwEiqb+0e7GOBL0VzPZN03mpPQt7MFjl52bJ+vllO
/9e1sA4Adfh34WZzQQd0HCtH10HGo4sfu1e0nbNgJ66YkP/iGc63voMleIvZ
Ts2FYxf+0ZgR/i8m0jHBE4cMWHxElKZR4VOyWq2z+GX5As9zRAiPqJuKdGqK
UVPWfTGJxrovYAjXnWxOfoDCkZ2rGqfbt4FsaVu0h3ES0o21lBd7Dz+31Hzc
82axifYkXJLLGS1p7W+66IPXWE+UFlJ84hEsXawegxJxliBQlP+JSb3cY+28
epFXhl46pg2RU2brlPhr9iq/d5iQ+Bl+NGjiHkB4je/pB+obyEqMPctfKkq6
t1g6/T3ZOOeBtXUmaOgSmkZpr3kpISzjHS4w8u9legREEHV98XByrWhAE+4k
757OOzRPN2rWFx8eNDoL6pDHaAewMgANS3KQBziJFmgUqhGnKYDP++CPqeFX
qFzYu1yVwxlJtLuP37yAfVrXjiOajhinygz4QSIUaH4LaQwZ92C72xCIl48J
K5hOL4jFmbecbInLJ1gUCsEOq+gQHhqieZPQzGKWb0JombC6vCDFmehICF0g
89gewjtQ+qOdhjqrqsFXOmO0R5l2kJB+EGmmSEftdgELfCcTY+CuXO5xRMZP
/bD517+ug4T0gn497vl3zqgrH4dBdyg17EsL3QpWavAhgO0AImjn1pFd0Y0L
UWz5yEMyJmBb6UIZh6NcwFR7TYsatXlQZxZm0YZE9dH3MVUNhnvw8djrh3GN
3RJSHRJsAIjhnsXJl9KfYP9DAjiTHalZgYVniOYdNg8t4cJJXNrCw0K8Ub5p
2ML7+OLYlVEN/IK7GYwNtwXpsDPBvO+lFcWs23EGlwyuA1NcclZiBrQ7mg3k
8PHT09HdsSsYr3HMcXl27GWBfiKHAA5XeHNPmlLGaf3X+Omb32nPM8p/RIKq
k5OaU/rNtvlf7UgAG3jVOeIMa5p/5sHSy3THZzwziME4WOzWqLELvzNAS3SO
IE5g0WTAasZvf1wIMmM2C0Y1L8Qm4f3G1t/ja6nFom7Nk3aUKhXUwa4kSutk
GgYHjJtWHhPcifyEsR2OXu0D0vElzUAXk1udfzblTIUcn5LOYnG1UFIVZl9C
tLwchQ2jp+utGnykkbEvirXf9fkw4zyBgcfWIomQJJAe8OCRYi6nHAa0s6Zu
HNA7mQlTlj5CRynGY3HZ6Zfg+JEA7TnKG2dpew4arfe6gMoDpzeN+LMJGcPC
UlezKvsffYOhKcUtPUHZna0ZkXBoutPO8ES39ZyWcgzsuIR241dmo48Th1xz
9kpWAW7yl1mh9wYZqqRZSJda7f2L5azvo94ew0d42xi57PamfSD1lfDBgZbM
Gblxr70+B7DZg6B/08NgyGJ8ZNWtCtRy83BOxQX6p6Kd+p2F4xZURKN6d3Vm
plTeYej8x9u0deUbpTmFT07nIec/55o0940MtHq8kZ7MFjwfMAei6eWQy3zC
nwSsZYObbn4jaxcmi51hzHze/y4LBVAb5anqN8oXc4X9TPwFag8QdBaiFhhb
tYrLixI6t517Zn9oLMJPDRsAK2sQQZyGFYC6YyJHWqcVnveS8in6f7pZqudt
6fmw8rB0Pg8nU40fd4CEZANDWKMe96tsgp5efHx7j4+Hthk6ad45AjdakbDS
4eRNs9nY7bejHbzRj6VHjVO2VnDi7wutrcXYPzJQiRTnfvqPFc5wlS2EpkbP
+SeFav+3y8QdwRhmtoNyzw1pnLbaKiIjNYaxKCHuPB5cIvnfgC5o1cv+JrE1
CfQcdeFEtpQFG6e3WtdnDZh52yLlGNgH7sUTWDbxAvwRkD+cGoKtnUYZCaDF
41voXJjOBeHSur/UHMcuxjwYfv21/FvOqrPsHTi1iGyTeAD/MrkTMO7Ou6Tz
JoXJYVVxjiY2sAqx48CycZRHdClEz7Eby6P2IRpeJA2KTH3dtmbeTseabqvq
5syLtb7d5Jbb/z8OU0FSfcOnumPgPpejX6P9A4064jqoM50UC8CvCWZTAZOv
1jSXO6/VON1cL6nbDQ6CGM4wDHjYtKdk/ZLx8I0odqRJKdAsblkSiluHdfit
Wt0m67zESti6eJTIJc1X940CRL2baA5QJyGZccoG1v2H3+AddndSIBMqij6v
1FnvOCfdpsiKUTgA+jCzR0FKkRQFMCobRgYw88/VTg18nwmgh9vmSj7Zxupy
+OwV/r53EjS8psB6/h48LGmIxQHFhTFQlTZg9TE4Qec7HRrDDOuv+hAEjAiL
WYq92k8cK1lvUSQNTKhaAnuS6T2pVcYkVJPs1LngYdkDCAdnNmzqd4q66vSl
ZGjycie7ACEVBQ//c+0Ai0QhLRk9whtao2K/922M2ZV3l8yzqdTVVQ5dMIp8
3G45xfxkcOFED/1mGnRGaC9mS6yCc7+Gohg5dbbv1GY230wSpBx9doN5nE9F
XqM8muNPGthP+TJqwiOsnE1z+dNzyfaU1F+7s8Yh24yLbzA0hBu/xy5U6reL
9tRmfuoqi6BNpJ47RSWnlPC2HYOEeDK/ty8Lq11HT4xfumFm5eeC4DYfRJaI
QRnCZtEVt96C4GzJSTnGjxbkqLAFzRF5NnEshBM739zAqaIzNSEEeIONftiq
ac6xOHyis2Zetd0639RRkBL9kr8r9Gzgn9muWxoCaWdLDCgzuoqVvHKBPgVO
GDkCPR7XnjysSe/+L75tMIXmV42tLpOS9o13hDVVd1Jx2wKupcj7kJbLYLxm
hsxdahRKd882sj7CqYCWL3chcQHyY9ne5czZBV5hWR4GJUojc1mG6vHLtWrv
zHpR80ejO33TtkA+cxkA+CpaSfhlsx3uZOWSx7G5OUuJ6mv0tOpmPFWkNtcI
ITf7X7WrkrawOtjupuBae16BPG5eorMmQhf7XVTk0fHdjec5/d0s7Zfogn2K
ovbmOTdmmajv+FT09apI6y7uP3T+Vei+kGBt06DNoQzXRuMp4DTpxaRTt4+G
71zuB1usW41v9Lh4/hqZPYi7f9HmN0NNXjVquNVKM4MNxtmLIFrDbnI0mKh5
qsd36VaiCcL+iS7U+y5SlKi+axWEEhfJvnNFEo69a8LkNwI9Abw1sdohmn4g
b1yC8Om2Un5T5UShu6EA344GNmGR2gJb2QXWCzJ7wjoyYXyEzjoLC9SeHBD/
rg8n7Emn1XsNfly7IF83F+i0CeBotF4t4IixI4/8GnQxKRs5uFTRXPa6wIcX
cOjUFIVG2NK6H3K6tZuzqrFPE/J47ehVDsjPahEm1CkGAHLCOwSiErQd9OAV
QF/1QSJ9ZnEfTAKIpGsh2cZ+F5ySlMB2HPh8oGegWLDKVtS9SIx2TTsSGIi8
VbKzLcgFiG6csnURJmnQAJ98Dp0U/zRhw5zAnrDt4bjV8AIHi58piK3IFn6j
5NCmXTCzzLMKqRoy7exdwDaptnNmPhNoDkjv+k8Jj3IP0qwte/mXbH7QUn6q
peoyAn1Zk5HvFbWn5Fnq+pG2oLAcEiRlfJ70y07I/gtZP1Xb+Q1Qwxu3goXp
6KzTqHsk1aaDWWKWyuPm8vEwFofdBCOaJOBdmvROSfiz3wpkuI3FUK0/c1bo
xcASd5D9fr9keK/5Jm0e5cP7LDWgVGz4GAEP1VdEo4+dFo2yEwAn9FGwBzhy
QAqME1BS4VmPC3OkYGQ6qTNTO4J+PWuvtDMVNWHZYiBGftG+kotkGgJUozmS
Xhf0e87Iqtf9LjaKX6lMigMxy5ELZSn7b/OxU/DyuLFtzo43bn4dpVIjeUDP
/x8S+G/LLn5jfh7Jc6WA9PcP1TYvqKPkRtg4P9cr3psg8ly9J1IqepxJ2eDP
LvokUoV6xnYCvlaIukUnAeFuA8tYZ1cyeOBGZKnsVoTyq/+qQ6giHO88puf9
rKgUR/YSa7vIRw3QMaLb5UYnnS6QNcaTFk9Z2dmDwlvjj93esAofbwZT/Ttt
hZ+5ZYTZXwr1Kf6jbsvme9zWAvvJHFHFFmt9CTaj58/a0v0B2adD2W+KQW28
eGBXNu0Q2CRk4056F2sSlmQO1NO3XBN0Iw6ujGsL2TJk0j66D3LNxcfxilhW
Uy2xoVlePeT+33S8AndBepWoiEixGnvWIrHkWQVGN5jnyps1EnN0bbhZWpjN
PuVKlVp8cnPtYH+UBM2lbABaJ0zks/DwFFsyxunorEqQnjARFmA863W8DoXW
qH5EcZgxn7VeFOWtpIcu3GG7/eyOishYj3WpUwCZhq0G/pda6W7mft3b6xVR
qb1TXO0x1rA1MRiZJIH3rWh9QFOPwYXNAa0T/33USu+xj/vMLAYVphoQKixt
IXts1RjUl/bMgH4DdsTy7O8TxRcdn8PAJ5UdYKsF6Q5NiKRJ4BNVJ5A+JTMJ
UZ4WPyP83IIfy5m/vlwgSyiqw7+8GthdtYkkRQ/vWhpfIU0RCBR9a3qNbkKC
yAMREPYicc3yp2XMiq3vIlm1oAEStr4cD/CNcjdPKLg585lH6JrQLQLLplPe
JnaQkbtuMhKTOuKyhvrtt4X/LcH7NOYXLXMhJB3wog924e3hBx43qQ2TMVPE
B6pF62mIHKjQIR2CrKnHPpxbuxv+cuaoiyna6pBtu6VGoHFBoFdklk02Vz72
P33uVOI4N/iTX0qLQ3frygXAnPAXGLS+aCOxdkjKBswtHl7GoGI0KKdIAB8H
bcqJzQt6EBcBefYU/Xq/MnRwbbeDx7F5mq8yjL1Y9oP06nSTwRWE9ymkr+3Q
Jl2dcOYHgQoc8mCzP2bA/HYiWaUNS0II1nHPO35TVY8YGEhjqVL5PsMoBw82
1fplA7q0kUWt0eVpETQak90p6et8OAAb4NKlThg4JcowAUO2ofibCRNt6vrE
+OFOVS+c6drpnF9kOs0ZgZGZ2t2MYb9yGxeKWTcx8vih/7IY7HguC2sOq23o
+jX3vAVJ6/BMV5xl+wcl3uAUkKZ1L6Kp6aehv0jqQ+YugaGsOHM+y1MbvQ7Z
zdlr5dNeSPM1QXvs2zQdEvdeOpPsO89oEzChBlSPUWnZWhkEzXMySQT1k7Is
0+lvI1S/WaQgrIsSjYS3wedoQBVvfNjWWNB/gfJNukGyCPtGTf7Eg3iEDdqc
tg9KSRwyibECbWo3mRYmoy5G/ed+nBiFq10MN62G6MwGmVG0xnmPFJKwKvDK
QmTZ17XsZq6vfMAwgiu0jHV/ASR8UXNZuq4WChNL0+y6ubB43q0WeyoHBPCy
wsX4p3X4Ukp6F0NkRI06tiwxhbg03SXEYkufgIrmVVqLGCC84sWixlhSg9TF
NikmL81EKRMUOJRUV84j+ZBThy9nP8tV6LwrXrQVdAam4gcJ6m7bPZiqrh++
eWPPoJ21kOLdCLDkp+SHCiG6k0erlH4rcRx1VvD047eksGzkB3MouX26k/3a
laS3F4mIVyoM4M8YuTAajfFhv8l1VMHRrgSjhDwX4CEYnIbbM2/4VeWvYqKf
Nc089dyOezzUVO7E5/vD/rRtGAYmWLIk0GNTia3Aqx26bcrneihB0IHgAwNo
sTQFmRKz/ZQ+XVIjz9+1fmb0SolU4KnGVlSJpLXUTdDGFL567HKJW3+kStFy
jycsIgMMmOW4dhTsw6cgQ9EjGNWK3ujtgbA/XT5CZ4k5zS4QuojZVQu5mc3k
1JOl2Q8cqHYovJjx/pWq4SsCmeR1RlQpmEM6EXWztoA45M97E/WNwdq+Vyz8
04CEuptpEjekRuEQwgtFr5jOUrcRHSCWA7wTyHFzQegL+csTCi8vq76T0iKV
AXIWEuCrNT3xSEtkgzK1sgRB8wyR5mrpTgUWP9B3svuFEXJ1UuGCGtvrV+Fe
O3PSr42z/V6IC+aDcEPUoMtsgaS3Sj6JKXKMFnpS5YeoqB+qUbcJOLHGzvm/
VmNSqXST3yzQGdtDkM7GN/aWGCofz5GJtoKLOymwkC7GqtR68sCCDtQCYB1/
XlGiynHrjewWAr9FlaMNbXXj/tfxO4+Drd0AH5kz2C42J4bQat8yBJ4AQPKL
F4eOsI+0F+k1mkpoCe5DVvRoF3kh1DQ4YhEHNMztetzIdhpquXHFcjwEztwc
e+XUcdoPqNG3FeWsIf3rueOQrZSboDOVrEBkolFVvtRKBTSlgPnh8e7v6o2K
p5YWqVGDBsltbpNf1PlLZDwnqIxbS8nKoRItiKJxcSdUGA1b+bUaBIkY2ofi
4SdLwD1Y6i0Z3UQ1d9GnUua7URc1iK7krpn2DgNvsblpjQSWYLK6tEfSf+3R
qjSMeAux+Mtpy6qLsp8uTIyQHwMg3kYZiYLL3tudCBXh7KFyoLiJJVBaeFwe
m/0LBcc2PRUNwWahmfa/lwKUjyq6iGKvjxMWD5Xaok+Bxa3xPk+/08tcjMv4
7WYGVHmTFbA7EehYwRGXqFbA05HggscdjznsBo8Z4iTa41jklYJ66yQEly4T
VgJrXB/AUpFpkXnk3iJvQbCfwsdDrIFl4kB10oWL2crL1bFPuDLoH6JrKwwV
zpmrF0VlOw12m/Id5xaKPHfXEMOqoR6SzPXInoHT0VzSPk9EW9vZpWjaPNx1
6Xh5VQvLkWYat9piTzvWU2Iw5bx8NrKwJ7sZSnYN10pNXWMMXJ4R+ccpqkEU
BSjIU2cmiANBLlFzwDSEfZQ/zMyuLrshSxZPYSpFgeizs90+ouV8ku2sQcHJ
t29VulvD17t+JinoSMousPDUJ5IWG0NlnGBFMnIc7CSZJuRXqiCaWmeVMjW5
uYATYJLphhhNmPqWjxgXCKPEewvZPQZCRQaq2meB0QrFXnVNOiLU3g2Cw6/v
ULKA4Z9x+KHERUWl3838JzrL7Brr4bpNy6pdAuwWU7DvFwcxHdpPtx/k6tyd
ernBV46HoT4/SCiwSSGTpQhp+GG9/T4CT5STRDlaxOQbdjoCskx2pI7xsiUn
MH82gd8LgLIj9m6Cy/xEtKlcK70V/b/Bh3WuRn7k1OTiB+X2k5D2mOxNRG90
E8C7TL1zKUz0bHM0bRyTVC0voHgEJw0Jd1m1NUOpgurk13Z+nQGhFJdgNIVr
dvtj3QMQ8G+wfHKyspkcZtyLsZ92CX1PosBCpUe0ga0A+OaGS40XQ2qt1crw
A7+zl9X8WLyUwWHIFnaxmDPlvNwvet/oxzN6W9NkPbPaqPZkzMgVVoEe7U3a
lF9VNKilxjzFUh4DY9YzIcu8ent+bxyPLkRwWAh6F8mnFT/q/jy2baLJ4f/K
whRuZHppQlH0nYWJ6KQT1xiQPrlE8GSFTgiZ66CtSgej5eSWd04JEhn7Rv8w
S+AyH4dvm6q58ls/UMqRauJZQVtAeNf4KHseTD52zKPxYZdx/rxPwTXKGq/R
JO/o0C8HLw/9fRrRqDPTCjzZKYkrkyq2rRURw/1OEltdmFSYu3+EGzXBRo0f
wKtCiNI45mns75xEhvjjOYXHjLABwmkkwThzehkPSt0bg/RJg7Tbm9NTfKVB
J32GZHG9/9ypD8cJTQ0rbCwxUtxOCaolChnnc5K58QD7+cFS3A8pU0OKsYll
Kljeq4bDaBSmRT7vLRSLfFzUpsqkeiTp0zrwPIMWP/PdD4XtKgYulG0rv5OF
UN3RhY3OZgcfq/izWREfBDFLUII2XTi87PlGS5MMdvChNHQYv9GOQZlMXUS4
XRjUNjvQ1t/+8rSACGiy9WAxfLFBAy4cJ5d99KzhPtyG2MB9Bg9Ve5QINxg7
NEGGV3v2UW+KK2PtK9nT1pBtlxRLpqhW0O5bgZ1XTyXY40e4iONWyTZeaF6n
3ovr/Hh4CmbNwJKOzztm0Z2veA0fyrj9GYFTryJPScCz4zy6pNgEH937Wlvr
cjdT8c8LrIeZq2jxKBIr0Xe4QY/vjK5+lk+IBCShrHr1cIjthHPrqZhl/Kmk
Yz3262TWD7XH3hrbFE6ARtYP1SxG7hqMxxXzPeRD/TPoeeuU1/CoaQnm3dbz
n+axiCd6bTRzWX2HuZeU3W2dq3UCy6F5rNuyl+fNxCWuOKpHiX9XZR0D/bk8
Wk0xxgaiDoYFgiOWLK2YQ7EJRFLXkDFtBEUh+YAGXQe9pkhGYEZ7anGDynbA
wMJaltF/wU4tZtqeDvBjnmPK95lAqb8Kyb7uu8QhT2G+8FyCY7i0JTpWEr7c
RPNXoz4KQFRc/3RbYj3DijeKks+pny/a3Ecu0rxGIXI3fzTE+GolfqpJ0Tev
IyJzV6bwGQ/GbHLHBzu/hvlySJUL8uTXpO5TjVOey722YTCS2yxA10R+Akp4
Dt7CYQp44ELRlQ527QAM905mWyH20ZfHwN4DtO2RW20qumVO8dE3B2dDipvt
lv9nk2TdTQrpugQKD8WkJIrqLAWqb6kf//Ej82JU/mYzlLnWyMzJ5j7VDHpq
TIXuQtR84ROkolay6/mfNYDRN9k7vyWE3W2nI+FHJDnsGL7MR5ecYF3D5owu
h0dCxo0E1C4RGwCSDNYQDWvCTCOMHaBjErFZmfBIsTceyFUk6vlyaKtIqdIk
UKJzOTkiTb495FVbS8p2OYsi3lKkQraWkhYn9MuhGJtg9w3R5ASgkL7I7cqo
p4ggZZyyS2rVqUQCnDhvMyEXSXzGkfThdZQ8KoiVU9a7sNXKH5Ff4Xl/iqpr
jFAkgzzoYvjyqD660qlqwLDjq02RVL6w2MfUqHCA7HRfjZHoIznn1JPDO8gQ
/8aqM7dTI+H/iQpal9pz1cCEn/X7PAEGhuGq6oHVxXUeK1Uzrpw6XvUA6tfy
I+7T6l8uWzwTKewy0ao6e4+NOJXeBT3AxEZI5S6e0b3SI6o3QVOR4vrRc133
BMi2yMx297Ouhdl+EAmkqayDlSIFJHXl92tLVjrUs7ZfpoSOGFRtRtohw7g9
ha4471rXh3rpIpWXhsTDrYQm4rN1CXt0bCw0xwylf1y9od2EOvihBiuyDH+g
Nxsx0SWy6GTr5M4TJ4LPes3fy07TA+a1DeeK0SJvbADpxNlwUGyJZ4X62wnr
9bPVkXCzGWeI9e7sjfS4Mzz8woNzUsdJnmCerAK7Ica9AKmpALb+7U00wHRO
KZ0yO0pRus9xE1M7vjDDDa6r359Ql9FvUtStk+EnP2xQO4T//0vaxOyCDUpY
q/KH0xjTo7gnWwX3k5wKsJc4wDul/z0pwXooAqc6j/A6OFlByAXADdD+7Ahz
vXAAr8Hm8pBebFJxwwVJspIwfejecuPizaThSQmmqcIPtqyHBkBoULUe3wZ9
S4uHPWzwJJ5WmtYYrqcsMB0xiPBpRbEPbxLKKi8HWzNX7u8rG2Sw0d0izM44
pbNWyTtTtgVNlGb2QaGqU9M9P609mGjY4D+2rH7MqDOGmmTiJpQJvMg4Vrm0
hpW/M79uAkzPBTF6HxwZgHizOndcGiB1D8I6/noeU0EC7yJY2INbnZL2LKmS
xOpmSnFcA4wkh/Sos5fGoEHblXN3fsZAjTaEBaMxjShW5mcv8tRY6aTYBZ+s
sYb7hcdLeUhONLaXw8Nv0AF0W4dAbYzWsxdQsOaD1n6GlluCZwCkDpo/krkw
Bx1s6DSlMc/bXt4YvQZf7kmQJG8TrF5BtFuNWAvP/0qnFraWbG6Dx0rWnQ/P
ALEaNkHqEF/WArn5El+LZR2M9AOKIqeI2r7/mDVzs4gBO5yHwF5irW9UDdqG
0vqJZQ/visa1ENYugd3BrxxW3tD145sYxEN9LCnEYy1bd14ElcsASmBWqOPw
NbiruT2jl258EBzSZRBafCM+/dRVk79e+zuKJ6jnJR053r7jxli/88r0aSZR
QpZw2m5CKysikpIxR22phlog4fII2fNOESGaZOW9PDGZXFsLQ5YigPd1OPj4
iOUyPsXlmS630gLh3JkYO2b1UhYNwLGcdX/5WTm1z5bp+bwycT4ZmJ8d7JMi
K0TGUvYKqbpPqN/SQg7N6Za6ORqm/F+LDxs5e7cnVQcoTedhYketWcp2ywMH
VshqN9JWLLO1MlAN5Tt/bo0jhrkzdQAJi6Cp48tAOk9IZSTA9KJJy2Lzs6aF
77M7Db3BRjovQ6Ad7+M9GgnRT+nPB+WwSoAsWf1mxv5k7upNv/EFugF+4YDk
2K2Yo2cHlP57eZLaIKhBU5/0jGkg4/ujhj6ZVxarzLoBitKWLI2U/rVvJNkF
iHmCckggShm4XZGVyn38Ikp3QY0GjU9YPF6CSM/INOskGhTqMzUD/4i1+zSs
EFs++Bw7gda9exAbi86Ki8q5+tRlAJkLP8CtQHx0hzeIql+X3CqsS8MbR+V4
d9n8c3w+dEVmZAAie2TWDB7SEyRxQoEkF8h2X/Q9zKTIBFex/Sfhi7LmDyj9
2VAjoJD0EECXdVau+Xh5O+eQVvBNuBSx0atx0jcAmJaeZVi56xTNFkVv/9rN
KavsS2wKJnfitNIUDArfTsahz+IeWcuDkWf/IUBat9Itt1ID/Uw5y9fUdCM3
C+Wf5YkiYpFIHNCwxFNizfR1jUYKevgDZuHhDQjSnXXczS3fMwCQPa4u4mFW
Vk7uKJ+q/jYVTrL3TNTYPDa5xSBsjZ0VeoFrMjTzJP0QYvnJnkOHS/YvTSK+
02nQ7T9/dCG5fE/5Ph1c5yRhKUI9VZaslkxFTZwzYHhAHOEN64glnbF4b7Xv
hgnJ1FWoL+F5CHF3jPXzquwkO+NF0alncAQUpatjcvmKX3EqqFnZPbNrCk82
AtT0ef8Kv3Z4G4hFun6djlm9rrdNenq4JpT5h4OYS+TF7aTSuG723538K0pd
f7hBeZXc+RRhnWjdDdvip2QTwUyAbcTlGS+p/4IFmzFZ8oMVNtTsvopTY2nK
5j8vtSkVLh5AXkibjFztvgZgkulwfoLrDwFssYMSeSnjyO7MleN4AjfxFrAX
jJlH9HtOLjxSo3lpy2sasmZVBuf7ch715AjG+FTtu9Dsxgi00F8m3o86wFrX
6sq3Ns7L+Q2OhYiEepWU1jSXOAAQgcXZHqSDD0yyp6UUzYkX4+wO94E0KTIL
y1bDUFrw3ILEq2mdYMrRKd+t2aNm230jJMxf/J9qM8ISCt+3qhpHN4EhnqZ7
SNWDmSx9ns6WBAt7eotVkoS94ZQfj8aQIlBNuSXieQSTNaezG63OR5LKlo6e
5u6JO57HVBXvNqkk736S1cRFhfyo5NzOzXbQ/WNXKbbJGvuN6C7AcqWrARq2
lf1VOU9BcM+HY0UEq7wErc2nxX4iv3vF90pN0Qih0VSl8aFNIu7x0Ut0ZNsg
umanOLsRgoC6s9CbAwNz+mYxjoOJKzugtZHek5vmnonA8/OPBLIvTU1JpJ8V
OLZyvYxz4svJAhvs7ZNH3Hy4WjPkrmPJ8cE7BGsapgobBjngfycvsZcqIyzN
mZBWZgUjsVHLsnx8I8bRBT1tHf8LFhliOy6EjpuaneQoZJoTOSPQeR7OXFek
hUlCRQZB0RuWH26JvDnIA25t0y6CfkQBM+Gz6U7RlEt6wYiu/Fm2vzRdu09F
vkF5KJw16pe1dgSmGY4F1q1eNxx3Ue30S7tT4hyc6D+ZCtMuqypyzsr3GesD
GvGSg78SUsXj5ZTI6qy4rZwyEXCIdI5L6ekXX7v8EceFrtbkIHrfv0qPLfAT
xRtEdogx3LAMsHizWoHERSBI2rqYzm7s6bNwIGodbPeUCtIaKoIRKe+I3wDh
ITaQeT9VNkyB/svg9P/xXbJXBLofJT5uVF8cygaR4xod6fqTEMCm7kKQ+dhU
XrnQ7k5ySXkcAgOkFMqlHveOeCZy7lg15nJKNUbcDFjjuQxmsZm6u00sMJb5
JNtiFAqEeuKXTJRS7mcSv58rZVYyES/Rc9szgNBk+F/5LQ5Eb7C6c75z+FM6
aZ3ObJ4tMmffEGoia0q+28KFLsSdDcb9WmUCGzi3bhxOE+476SXvq23jWTkB
cH4UXjuOU/aHyBJzVfzXeN1m57a621x0bzx7PzzaoPcLAGqE6FsfkYCWzMY0
yBJj3FY7jk+Yw7iAYd0Cl18tTUwbtgW4OkQ9K3Fzs/vpK//dKwoeN+B85Fcu
R4s7kRlgK+cMLHJZ9ZHr/8i+GenhTbzEoehxQydWslVwOf7LQR3/I0LAVt2w
O2Jlfh3iowEqclsW1zIfjigBTmAS6ygq3wyE0CkIY1Qs0hL8qG0bTRnyL6vK
d+cR71tHsvPCNyRp3nuSWhL8DpTwtgFr8GYKunZsaAY+xH8SAmnHLMwLSTL0
ziKLXoY3alCf2tLAiN+XxdQH2FkeZH97R1bZ5hlcMJgGbjPz/pvO5npsENpr
zY5c6zdO4jJxOboMsWru3bnh/64vxa9VkKCxZSuunU1ZzJxXdkr98AOrvWvW
JP9klyTuhkpz+CkmyobwkTiSub4f4iRplKpicZJgqmECmS3Iv/uMBo/KOo8h
vHyJvqMoMubSjFOAtNdypEkSDAr+KWbjjFuOz6tgi9FVwT2EbcXJE3ZJGUSx
vNM9f6xdx0+m1Rr30GYkcwZq3MsWae9baqKvwCU2cxGUNRTvOUd0t0Rsz3vb
WhlcTxs61pYopGjoMTeJF/o7+aTOWZxflUL0Gydc9Pk8WkgFK7Y5GunvO4vV
Z0mOr+SBuchmDD1iVq4/cLm3e/IkuL2B/afC3/onifq2ZNYXqOhwD8Dr7poO
1ftTlHc17cF8D4I3jnQ2Ts2KR3dL/mTesRL1FUFjZoDXaDgtNoVpaaL2kXcB
6KXD6WZMvQKOzjwvJlQ/qHd0TWhmQliHOj+Tvo4hlq+Pe9bbBh9VGeer8JhG
LrA32KAp5cFAK6ZNtZTa/Vf1pbdwFi5Vk5Wnr5t0xS/xUuKYhbrDDbaijiNM
r2lP3NyDad3p2T4OmWoK//vfcToPnGHGnHdHSGxz2KIibagne/xDy2XBtsgs
uvhhlAreAB3F8Ll0g3j5+zdrfLC/8cypOC5m0LJC6vK89nhx5xBsr82y9iGp
oPdqCtbZdBkTrBGWQKxbuhWy68CBMtkuO+yUZgGI6zpK0TMh/7V/KtLH9Nhc
J75VIu31XxToz6kTeIJaW5FG/VnSGlDj5hiNm4VX9n03WKuN0V7ZNQJfuq0r
DdP9F2rFrncMyF9tqyN05Q3KYPhz2dpJftgMyt+qRUJvErIAsBosjdIwdzl1
XOZD9TKMUBKnxcK+LKfg5G3TvVZ6R+4DHkK6z8a5/FZj2iwXZNyv4s9ljAus
MAJZtHPgag9vRaqlxIWZJkBses32DXfi/csjNBWEILQJvo5SVeypPqY6e6SM
+RV5xjY5DHZc2gKaNGRWTUU3Wiux0oTZARvkkQ6aOkeXaYRfeXwwgQ8RNlWV
8NfP0xvNaUyqvxfYPV6VbkM0spB6A1S4Cf1sbeeUsJyQJOdwg+StxRypNyGI
8Jdcop0t0v+teZazF4GfsxBFDkaCcUU2iEZPWqpnMsGwZYVnFqzj+snY5Nax
9xlZARUD7JfovmuDdVHvlEQtDwkZobeuC3iAtuoDFSqOzHfWYgtW+6tYc/7k
NT/Fs32RO02VPoZ4f07Z1wTuIR5RMW/CbeD7KCDTc8ETTZqUPx3O4ga8d8W6
S1fJsoKPok0tvA05JU7qbQJulxCRrKlL0PxLGE6qF7oy5VgN9K9Kh068vEoN
BplHusyvSohkooQ6V22Fo5allR6h/zLA4fxDUFFIjp2DHpr+Rb9yL4dm1MhV
2FfLd6CWEkt7DxsNuUVlW3lVeFBhxxjDSfPtWHO01uYIqL6QJ1qRHWJcFXPU
RR5XdnrsvHjrjJR8P3XMHOXXOcuyI3sjbb7Unq2Cy18aAOt1yS+MAPURuJIm
6TSnK3hmjsAw77Y/XwR6eEnrr8BEzZDxR/HuwqFP3zPCcqVN1fMNd4jxXzFE
/r2xLRszFvg1P0j0EvhP3NN7t/S8qal480lYe5x5yMMBsD2X4MGlJi8qCGSy
tWuXEgvg4yYkWzonfs1HFq3jQm1TlLBvJK2hxXZO86OL5SBC5YWDEKxvj4L7
5Pqn/5CV3JOwSBIDGad4TEVV0Ct9BuGlDkSYhrXClgH8WwR1aLJe8M45+7nI
YcxetieEA5Vm7XtiMkKxSr4vcIo20fEd+r+Xtm66ckbVbYSUgCPzzB2WXSVG
YfRfzLUxLp323t7gE/kame0c5dWgZZeirxxwjwHsr/TQ6LbA6QmxHKNTxaBj
NbT+IQIa6m1cX4nSrNmJpIAWxNV4ib2WQ6nLGgnCr3pne/MPX8ePKw8JqfKL
IDqbH7LRKJ3DBJE/NloZ/MWU2x7CF/bH+/KjdiK0t3LkkHC9yUMva6MlM3SF
MFPt22jNcLN3f/VY/2OalyWJyzeqgcMv6EA3lxT50HbX0Ykweic+B00jdcm9
OBMg/f+GGZOvBGqu28ewWtJdo63bT0XIztp13D6di5U7giOjkMF/3Ak5hsjq
EtJwRjpRoWRHzfBWJoldvFMqeaUgrDB0rOq0NboZqhhtYxdEllAUD/WilsZX
7FiQtqm6dN9UGcZWicO9bWUBLk5hx8KMsaXdZEyF8UtCnGEGyKQXRvZhSjT+
sxq3e7yyZoJlJ4+488JpqUs7FB9e/6Q4mQdJUNABWJRjuHxw4B2m2CYsgPYM
ayXdRFp+kvXO0yA0w7dorAmc6eOWBE4F5YGK9vciM6Ez9tP1t8+eUXVbB0rl
+PMTZF4b5tQllAX4HxSZURi+5HnikKGZ1vd/+OW4iFQnXeyjklNmtwyU2mAQ
1ccN/CTA+++yFh7WHB0yj/J5SXqqCBtzWWJk9ex/GHGbAHBb+nbjMZDZFRgw
tZ6Jla0aU7uGmurWh1fE4fODH9LazT9OaNXFPXOJMl1uuN1Y/omBTEmbt9dY
LZ4eHlipBPqztRcqdcmqAM93uwLTQbspTRTQGN/Ahwx916hCDp6K5kas3PdG
CMRR3wT8CIEUJsaUxKUmG0Z88BlrMc0OZc/BtsypwgOwbo8zVUaHbvfzwocl
wdbofz06rRH/eVRT8yxI1r5QfbvoW0po2WVVgTLS0HqzxXrk5hXgaO0WvpXL
WaymZLgPwF2lhe8hQzuF/4b8o+r25aNijewKi13X8hQnm1msGeED8pe+tVVo
Yzk9RzuNCy+qmouA1ZMXxYWXnHK4EmI/NbLw5YID4kNZsiDNQgL8jfpnSxCO
9ljxoCHn5kbX/VQk+e2vA028AGdcYNYevA08OoGsQK2iIZpQtPlh/JjjAwFD
w2wSCR48zQpY+1ytXSFL8DSfxsSh7Vg+3oeIXvcGPpR1FLL19EMNUA+o4VHa
ZJwXG9yOlsQe8DUI8Z2ocglD4YyguiFQAgxuy4m4i7K4otBk450J/QtIyP1T
3Bs0weJP4fSqpOHWd2LpSkm2vRISPsjTMH8+Wjv1JFBUObLgXC875LIYpkeh
A+Lyt1CVhxYlPMytyYiEH4jRr/h4Fnpr2AZydmL2p7buQ4UDA15aB9Ngm2wO
sxubAfyFsFeI0qocS8SIOawgVd1LQEcl9mhuCO6Kdg3xcbgn83DM5mpWnmyp
VD9Pj8rHVOvh8oK6Xj8+nV6SlNKrlBDbE6MBk6wdVs7HO7cGEcchqT4qpEUf
e67yo+6q7Sk78pWhgWcGlSxON89Ejb5lvX5Sc3Yv6eQ4Ym0xcZ0SVTkTlGlT
f6CpE7BJ/MSmE/MjUugwD5KGoHyTEMGXaadsHkuXfUmdosvOLkhNKT7nCXv5
YJu77UXEwzAsexdIGGgvmxIwieiPA5hSvD4buV+dWcZOCI5HVpfLa1/YcY51
+mxaR3WdFdTTnnPB45q4J/azgB5NVh4rYAjuWgI1dPJCuKXVB/UUJYq3LI/b
occObaZZh/39PdnnAFjcBgGkqdy9wz1N71RA7R93kvBiapNOgKr7mtknzxIM
vqO6InAcn8m2a4fgtU5CChhlAIkp+tkhLjzCwzSKJO7c3vhzFIKhS2JQQGHs
cSd+82NCJ0zFpzbpt0FkI69u8IgOMpCRdOV4hbjMxsZ2fSoDMABb5TJUvgP4
roYBIHv7q1BoOQMj1NvkgboCD5tcQ7r/P7YqzcjTcELH6zGL1iV4wvUgrUXi
m2Vx6ixI3a/x2or5+1xwNrV1YEUZY0kJ0fozmkE2Wr8pViKvqN3BD7SQ08KV
Kk2WxX4ZWTfcjxZjLbgCWdtxCV6q/qSyvhQXj7eFsonOnu0dLsiwjwn+x5fv
T/JNC33FHgjuonCkLARkvSLZm/TUhuIvYkAdE7KxokSVw292TCLwsv9Lv4lN
Swe0+HViyqBvdb+737P8S67YUWpm4EUvwK7LDHqYM0qqtgU72v/J3xiynhOc
BhEslZxn6yr+T/CRun/cCV3OZo89/i7jIKzUXcxPFk4I5Jg81AZMDbGOWhLZ
0yeL7Tc9hZcnGn+mWGgx/HqM5HmfnBfJ6zLJEr2vhKnsav13ZJL+FnyqXUGe
XQ/sX9znIfTLgRqnElB2iSEsqB9oJ/b5Jp5bWIa+mvdLuvzv6bQW2IUdnunb
se8CQahkUO+kV2HU9mPNwWBF5Vhu7yBPeXH8LHam2LkmgEb4Jsdk38ImDwM4
HjzBaHGmP+OgrNF3HLwC7wIuHQhLoCeWAjKrfSIWpSxGv8Vp37MKLa29ujgq
cigO49M25iCaOHhVLHtbbUAfgMtpuPBmmVtUSZibLhwDzFFcub8KOGx9erCC
f7P5fFNf5bCLx1O6UODDYk8rSIvUWyTq+2M5VRH89FQlkCn6Mmu4tYx2m6gO
Mzl0qKID5jl+GKTcefOtlthKIo+HN2R1sYi3666YutAbsTgz/Ou2RiRW6h5x
IgR+2t2lmeuL2IoPUOFoatfYBO++g7E7ZjRYBvCj/k8pPxi2Vf0L8Pol1TYR
Tpav7iW/eoNE4LsOQf5TrK2VTN2gYGhcNy3aop6H7KYNpYsK//i7IYMqbhW7
/Fyo60vbS/Qm1XX0+IMrHgI5y/Kn0FKyusm2t6CI2ywFQtyRAJGueazadktw
4ijnataFXKRlc8PHcvTzMnVMU4Uejch0eaVrrA3spRJjSrzvabBs3d/f26cW
kvP7i5m1Nx4A+bnS4K4M4RJO6W5Z8Ez5yPlLMAsDNWjBx8PdupYZTncu4Ei6
cjSDQEPDknD4/ytQ2g9ti7Y7rkjU7h77gVIei/TCgyvmjkxyfHzoziNP9pre
YqSPNFORtAF+Mk0ZXDPKNLUWjU/PmHPKOqjvjUarEPRpFUlleSKzDSoxQsqU
0UYova22Q43ZzVq4CdhW4khKSXOhCJXBqBD9bgByr0bqd9I2ozv3jav2sHu5
l4/AF1IZR0w16/5/bK5q0RcjOcRSu+P64gdDNg9G81PQpsRiJZxgEqheXUjw
xnp83CtN81tAYXw7ad3vP+gGg0Qubtdu8KhF56w2Vgjb6X0dOkMFTmURHbCp
osv7Z2BrbGZAhI1bGCHgv+KRE9TJKvzsx+bfih81yXQZFIBDdh3bd2efCrO1
P6/TDjYp7JOR1mWXcXdoIf9Sj9ghkeVqUieHHQUtT5DXIbCQIUIdmhvp9m3P
Qjok7qzHH+ne4jDszvCEKExsQqulQ9K0YycoTofsA23N44zeECnOkX7D2VAn
4htRPNb4liYWHjGf/8wxb50MwhpKSoFnjrfHD1BF5JxU7Fde974kUjFqS+Qy
WMPSRNp+NcXvtIV7fBIld5j2HZBMpJ7e7LE7jguvf1MEECAheZV/hj5Fo4dM
Z8mhnaBFYehqkHzdC0/BMrPhBNngx9AkvQSTFFNZhzkMsYGEXsgwXMNudMJA
YDsFLhrNy3lcgLOMl8pJ7va8Y4rNu5WZD1vvHnyaE3p3Fox6ZjVkXlhyTcA2
5gglPCGSf4IocX/E7qgvOzvgiR8kvDbVB5RSUbdW9QbSHMTG8xuGX1XBTDyE
Kp/HCxDeq2O3pZLcc8NTj0yL8Txf6TQ/GvdzmWmLDUvIcvX+v+/+QDuktirw
4AKqdL6nP57RdXlwC21wi+DxCpknc8MNs5OWo8aYoECdBM0qhdQPkKY7IV1x
YOcoeXD4ejBIKi7pNlIXPEy/ICFi37ZbBiNY3pv2+RKQ8qumSUX3VxlzYMbC
jvQl41nA6sGXaDnc1Z4KroUgurQPqkLauoBFCrJGpVNJKu4LDpRSfZR3G54v
RUPtVmCcYHPbioJijbdVZ6DSkmsTMRwoB2cm77tHGai/ViZZRZih3wvR9nZs
XH+OJ4ozxeLgZgW2tCvBoxRw4B9NQ97jF9GO/QPw6HVVjBOKshC+Ar13RHBW
8XQ+Egx1+zS1hOoRRnEG9T7o7Wzso1lvt63d2HlUTdpKtzppk5M2BD7wkRf7
tA6zWL+s6OwXK4fyGbD8J8JGvRUYXtQp6M7p+z9cgfGonwtVEX74x+otlfZq
t1ObvEIfaNsQk6aaCIhjcG3VefskP5nXSV1xWNI3ErPqN45y5YNlmw+WO8Cm
aVlCw/SdbvfCoQduJz4pnptf+GdJ0343sblKHWmmE01T08bSki43HmdhMboM
skfRDLYhd/+XVtwzT6uhBJzSnb1P39J6sx+5CRlFsn9WWh1YnMTIH7LEeNKB
mxsALc+e0mKpkMEDNwAiwqFJQ2onT7LsdUSr/TB+6A07PLt9aNAbPQbfSmLw
WuQU5XRAo3op30DnwxUklVpYqDxLaFdIJUpX3vOiYE43v6/aiPWzqKX4xLn/
5wGsQ/oRtckLza6+98aG4CUEnT0O+36f74ZhU8qysdE2EfSZz0wh8ngb4lrc
Wx1GW2QUB1AMe5H8lnjYDBQA7uCIzKjWPCxOrsy9qRJz5gkf5xk3+ebSufby
9jocGkLBvr95E/6CVJqb4Nfk6MPLKNOBKFpNDwdkbqERpVGxQ3rdamTSGlIs
S85Mm5+DiP6RZnjOvfLjJJJk5rmRk0V4+0RrRdx6h3icouAkiPKvVMV/ZZLY
6x6vmQNTA5CmIGo3RzV8qouW/11gJYORlHkTOwRNaCEJ8/pop00CTFmLod7q
F7lgQn7kKLLKtNLE2ziNB2tI4PfJGnU5U85jgKJ23VRXJyqRYnIG5+4bvpMI
ze4f3+SrmZY6K38PrYC2hr63qXTnhfwYTwwl9xP+LC2sksEs8hb1zPE0WF6+
+GakrDgLSm+RJVSy6jsej+CESvrUbOeE344tFSjA//jeurnEFWDIKWnhZKs1
uBMOo6otXCdFzkt6XktvZkrgkPtK3CLPk2Ellrazxp6dTPZb1XtbHMOwf4XK
oeq1ags1Fkuan4q28ZX4f4SIKp4pDRAllLRiVfFDK7j6vPhz3hM1QI1p9bxP
cXVFWZ54vaUEYcmr+LXVBTskY4R0FsPs51fp2A49FfoRvL3diKXmRXmthPTl
uVLLBFOep5gPBXkOkXcPZquiOrC80tNBS7HHWqZKdFKoBWbrHCVlN6CTeUBB
jgw4a0eUa6JRMQqCsgl9y37m3Rx+GC+apgr7gRDb2VZ+Rx/YGK2upBrpR7KZ
dmahZAGWfRBggSIVe6yVEHGi5tC9S/95U2Gqhi7O8SdUJZiyFkJr7khuhrAl
k3f5Jlt0USqVUi7HmSbj3olji0Q/qsNVJiQWfG12wCCrYuEw8TN9uwRCG265
oXXC+nx7oES7c1cAWZEOjskYXSVYbq/0eQHct1q69ifWpBs3I0t4YqdrHmND
oj7VzHYN2XOjiSeehhuVb26YRyZzorwNZkutPN46Fkkh4/7428MIaR1tNoiN
vy9rgtOjOZ1WXrAF9MscCDj2BiaAHN6CuMwOnYzYlu53hTVn8OIbELAmALjD
vaPFv0a1kWt5AOMr/Z7pTILEHGqG777mcUfX8lS7NkcDXpc7SgSQPZ654mNS
4ISL9X4Ahlk6INQ7J56EcOKZAdZoyQuINd4MWzoP+egq5keG3s5dR+5i44Kl
Z1NgmDX9uVbeWFc2iYPto6HIj9HPOXjWB9tRZeEBVxRlygh52asTHgEEPhYs
tzyLGK/JjQVKfm96z7cN/bfv+z1MIzSiyflEz7060c98Elmh+MeVkycHgApl
sGCnXdQHgeerpl2m6cqHYkj7gbszqxfPb+u+d5Cr3bh/7oFTu5ycc/lh/XS9
1L1ei1rRXNt4Es6D4RBKVySNSHPkrn/lZM5ISrB2WDRpvK7bFfSQtsVg/AHz
F5pNuPbkiplxA+2l8UTezic8KblJkgsasOj0L5pmnlb2pXcxSielRXgVmZAd
0qWSqhZkMmbKoqRvGvl7BTJPi/RPdE7KdF7DcIPLZSC1UydQxjncLVZ6YGm8
IY7X8RxucnxJWtrKAl/Z8QE8/eeCKsL/fku9gHc/87jlLIMEflHSKOM2bldZ
rTuFHbzzu/5tiZkeHmcJcEG9937tKCtXn7gD7w5NZsEAsiobtE2c6QgVuTUJ
1q20iSBHRryWaXaXGp8/V5VZrGM750eENy8/6wwCB+lvlwx8hafs9c7ez+tA
H7yF+lqeL6n+zF+fegn+koFVYYFTj4vU8gU5GBxuMr7l2WhQotNcclPR6FRJ
rMrhCG0fS7qxOSwGQIJKL+ecUw+YPEytfTwg0B2adIVLYdzavz/oHnWlJt8i
84fVE06oMWHo/9bfXXF5BN0ZSrm1C9dVoA5Ujg0uI48iJHTqAHYBWhT5IJA7
t3CllI1UPtL9TiC6Ce7H3DlT/TVG2dzh6nbnHEm7bMJvH8gnrgPwxstyMNHW
DI6JpyUY0RY1wLxZlzv1zVrb8smNWULPgjvvkRKzyzjcUmTMdgUc+iCn7bIB
YdxWejh3CMr96MEMEH4poRcvqaVVgDA2n4iSCestqmpD9ZMoZN1bLaC+6Lnk
tlwlZHs/9apZofPy0ECYr66T3Hlw6HJcza0RKu3bH9jnMcj87cOUOKLTFZSp
EUSD0S5IognbsCyaXX6u6Kj8evmfWsJrRbH2wkG6sgBpXCCm8kAOkExWgpSs
XcrkTTOa43tn1Ol4L4cIntJN/oMBV06dt6RRJ2r58b3QPQ+QX2GRkE8BQ/kr
dgfwFnAzNyqA5Mcprpf4Z34kHnJX8j1gscurRGy+P4aCGuk6H1hC98VZiKeF
Jkw8ktvLHuiF3feV40Hks9AV6Lo4DBQwQQfNGjnyZ7Hllsi1uDlX4+x02BPR
ak+U1V+6106Q+/OF6HguQhCCqXwg4acRIicC7h4X7DahFBqC7UE6MJRnpHeR
mrrDvVc7lVvnxVFXEK6Zrj6QXgD68xuzui8vF8Jzu7R7Mk+6Na3IbD4FefWj
OXNw/PZBvoAJrHuV2a0RlozJt1fo+srD0zaZZ5GUTzlGXw6Siw9yq+x30ck4
Je4hxolH6ayK9MS4+5MF7rfztC6ecbuA9XmU15WSJ7mAx9Loq1bkKj1UdILw
iDU5R1CxlUsWNxRBN5KT5YqzVWEkpifjFL/cmPPUJgezzgpWk7Y3a89xeOtH
VeDV7ELwkShSECZi9Hw1iJG/J25zG0beVmU1lJ/dAvrPb0qmANnzhf+vUc2S
qAbK7xVaPPSQNlPlVKzQcNFC/cq/wuj+r6byYxKSnuXMQGBKI77A6eFlfD94
dzlWQ7EMosBi2EqGyUliV0emb0bIIJ7b4E24Fzp4Et/xzSqH7naNLAr0WfSm
jnRu7VXcVd12rhy+GoJWQFh7G6Rwk16j9ow83lQi/UlCckswuLvejIwIC+2Y
ngHrSGX2bl8vxWNfoG49Cn5FC/4CLonlTpC0+I1RIYdsJ/sE8b8XUXsx7QFO
cr1zYYBLKtQNSH0MsI+NDKiX6mPgYKvIZUNL3XyI8b8/vfCwi7jXhg/s5nyA
sic1tq5eWj1sweZEY8kOtxtCsj4rxE8ui/5RYcy5QDBq+wlneITb80E24TnN
De+CAQ72rt4eLFYZ2IkzNvpQbuY6WeceXBKC7iZ5YlIAbpeq6/xq4agM0n37
1PaLDRF37/v6tCXWhFuINvi9ELBd50Afv25sJadPH4SDF/saODtaraTP3nQz
CaTmNEIhV9ExrMCZu4mS9DyhmtegxVPyrSBr++pW15zyfXVcqXZSA4gmAOuc
MHfjfDtwDQrMWdPJGEv0IowNTPlw75ZUpdi/KjVoBEpaKSeKRyuuxxK9S4ck
/LKEc4TCg0W2u2vU1uk0y1kSG7LSOTyuu9upbrf8XoIFlH3e3bwoMQx9qzus
l/n3cGvRJ08q8vnLeI3Uk9LgkBjSOqBxNWN9EtYpOfc8OK63XVAXaX6Luxei
eUWPDHz58Wf93EWqLFUe7Pk/Ey4cZKtPhOSNMC4Hk6l3WztoPe19YpbXlUGG
9qCyEoJTNu0LeX4dsAHs74esVGae4yIjkPVsvwKpFmh7M2x67hnk7yphudPa
ApkBXZC/3J6xQltXNWtUeRMOR+/e8hRgHtem6nOqW01THXw+L+P5MSxG5CpW
wrAeGrQr2vJ73/H3EI0JtuJvadwGblaLIOWvFLMy4WCGIAcvmclFb6NidTft
MpP+ia/+7SNNeyXnge1BJ+sJCqA3KjRAqxqfXtAuaIQ6BW3tgT4jnnTsE99h
FfZqgG6DGfCcBTKJfkVrFrDB9E1WBGHW4dlyWNnnwzRc7vOLhzlJyKc1K2vW
Pw8yI06OIDFaDsB8CcaAhUKLA4R6lHGJ5S11Zu59snu50S92VuJ9yNJi4ovN
yC70Go/Pdf40Gi82NdZhJXnjEUOJpa+AyFoNdhdPwGGWuA13I6eKG5dS8mxr
7CVaQKj1X+YbnV8qPjLynAQg/W0ir+TuqyvyCHpD05oTuci50wbneNOIO/AK
5O9Gh0MKOa1fyl0gjvDeFLtmACJ3R6w/95ihEPml/4sO69UgwycQdAtB+CZY
Bi+vIREMJgsA5qamHb+2BZta3vjxnizpOfa/ZD+YWelh/SbCcI0U3EjV7hZV
ucVhaOAeI36q+vSW5jNCQSmxFwD4WP+Si1aEiPHnQc1sZCGbS0LyBUD9qFZk
3trisz14sjeIGP2qtrESCuUNuyjiIeh9eTDL8hY9UPXcTTJVeVbQSLySoZhr
PfJD4KzdaojoZvl487/ZaqzKstCd1GusbsLW7zpWcX4j0pM//puhT+M8weHS
IiL6oQDlv2C5yAuB/p5pRm+j5ph53N6CKywevp7t7+vlztbKI7HILrevQujD
Liv/C26mAY6uO0gXwVuBd8zD+UtR6rucr3+NPD6HqbGZnKpNueHVPBTHOMZk
ybqwQf0GJbsAxWfksfIYKoTPuAoLYbZCfwTZg5/g7mIqSo3lk6MiCAM209Sm
V40hcWLdLyRFbmaitvbKkjqqYWbCWj0/QQLisu12enGq9tvAOJl5qBHfXA43
Ku1aowwJ3kEBfeUBEvV2HGcEDsJJYKNfjjnjyVeFMHPbFZwWCEtuJ4qyfSjE
cYXImNhQBlg/qnHWKDSyzK0KLr6Ep6ohEvFQ4glUyj5s2IojOk7dKFgo5f8W
TEPf7xEFh0Yqop9p7WsJwpW8eu5ftNZ0XEYdtPcHPrPp6l3ohKo/nQfPbBtB
VG+Q3yxAYEPCDwuB8LCCKoCtji2Hn6B6t0MIQ3ks9EbaWkHBRctdjFHhT0sL
qfUNFsP8iQDU3wNGJPb499RNvIu7bcH1DZ79NmNBK1s3WIcEh+M4k2LWzj0U
xcnys8FK1rPPQzXim3lyF8xY0IzFu8Htct1loHlEFaOeIur3ZZeGpxML6bDG
0ErOFFR0RUyxZN2/G8YenRsOfTud8MDl9wWlbQV8Th2dYksKy/Zk3MT8jSxf
ClnFRdBR4e2oZxdWoVqyPM286+edBeHPlLeBO3AoQPNSWlcqxPc8G0MSEeLo
0v3ft2BFEfm14ZCbmgGr7HCK11m0imywg+pd9yXGevGFjP+fuFiuCLt0Y+OO
adbQyTGOPlmPCI6dho7OUBPwsTyi+ijgLqFMPCUGa7whWFkGg5w7N+ApPzcF
NWJ3UIlcyXQ7fDQOfaX+eI++QJNESPHQ8sCai5RD1a/nz/0gugtynyyD3GVA
RiXUjD06O903/INZYgTbgfIslpWZTZZqi+i/BGUnaoxyMaECztRtJHD7QYvI
t0keDI3u3ilB//jy2/EZMvWvwkoUO7WpCGrv3/QmULPJif9hGU9MOPVoYePK
RYf8mfG4HwntcJ7lGxisQO1WEB2BrrGdcDN44vHk1gUeEDN44S5+cV+03hSx
tU22xsN2ExcmKJ13Blm4aANlOyGrEM1LY/12u1l5yoF7LrD25/srNnheOgwi
gauCcUnrNF9cpoR5mHb33/aYfg4N/W99hgFhbVv2nOGuLs4Y8Kb10QVfnMhL
DiE8qUwKqEJup9G3BpEpJHk6dVWRJf/BM7bumlw675z3elw3FcH61NIs6F7/
pclRHkilj5HTGiEj31ej+8I5SXCq02v5gakUxSxHA8qHdsVHJgJv75rhCFdn
3qZQgM8Z0/mIc40GfTtNzS8OVOb7cap7Fl5cUuB1aNO03DO/wV6neqmy3F1a
uBlwvrCSB9nKU0FTL1pX9KIZpDpXnOiSByoyBENz7hbLMntFqjTDFtw2Tdaa
A579Q2RogofZZDwSpJFvKjM7yercpQub/ILv6XjYclQTbXfH8B7sp4nrIIT/
OsUE3Wx63ZwRK8V2yjG26lbJIPCXtpGCYk1Nf0eR/aOXB7k4KOoGkBHGue47
MUuEPF4yi2/cH9/SjrJyHJKHrSc8NIF3g7SXqv4IAeRYlfye6QZ+uKxaMB4c
y24QNhZrg5rR9pBVWtiWHIYFu9pmR3ofMwxJnVgVJfBrQfdxreTGJ1YQnBsy
wvvyLtqYI//Foh4ucWnoN6FgJH/oZFJozK1EbPs8U9BiA8tNl52Y6ny+H307
wgt0tRQH8+SkZ5Nc5n4IdB2ZOOhxyUIrtQBxS9rOfUw4nGz3H8qS3/LTKPGD
dX1lDpsLMKNn8zNrSxXEosnmmyHyrAkdPuM92hrMANqh7pBedpXoC9lVlpEP
E98pvT86a3LubKq9Qx0z7BeDqgrJdc18ukqHjXd2uImGTnfS/Kmfn+SnhhHa
BJA+O2IfLhuzD/58iJxjOI+zeIPrYouvdIWbnR3LGPu9C3qvx4s5+sAJHY4r
ET2AXa+68YQmz52Ab505Oize5BdjCr4PPGftSNtAmNhgfikA88mvx7soeVkA
XnEs3ecDNn+MeOWIMzhYFmaSHno1n6CNpOa9XJsb0M1V7jIqdTOJv9i8YmzV
jtWcDakNw0HiVBdvWpiXJcM8l01VEeYCS0flsaueiXT7R/O0IonGy6xl4pSn
dh391QXYYSJUue/roHhvJqCrwi4GtMw0kq8zy+XzI8yPVT2g7lyqXhSCcsCm
6AkfiBSo/H7IO4YcZXqG1vlUBX8QW8hII1Eh86x9Q/TPcU4KjN30fJVq98/a
kXuAtyDKd9uA16gG0PULDgD+YTFKp4HX5M6k3PVZNbWf2ZZ21iDaJov/Ll6P
2Qn4GBbHyY5TD6WJdb1GXVaUlaZisM75Oo6oKq/GlBKAlwyEc2CYGGEt4edK
2humkbCLLgTus2tI2xWqOks0rCUH9yPlKA198DdeuLHaXvSKBK31CaRS2weI
tvK7TEtPQLhf8wD3y5UieNcnrksDVwtG0hAtcjwo1bEqi9h38kcCVNQemceL
9K/JXgDBiqY1Aqcc6AC6uVCd7Wlm+cPU/8v+C1f6lmUgN8Ck1SB4W7niNJ/P
kV6iIoNJrBHfYO2dFyg++wHEbLGYEPkk9ZpDACcVWunXOHa4DTpUNLKbeeJ2
AX/Eeb1XbVeYj6mRJvJREwiU+htrbmJU6BxqEu4p8EXoJYaJVT13REtN8kCE
cmrFkZpJrY11RmnwdSUP3Dlgu4injPt9Rbr4XFhJh10HKlANut6kncm2aXjP
ISIExLO+Rjy2ywEY+AWAGj+IO05VATfBqmtupgYAsZEsvjyYBT3rGnBDYJgw
aZX6o/l3eMqkS4oWsv+n5uGOTzgKnXaO8wiBKz2c6rMEZ98hYX4o0hCnanBe
+Be5BZ/UU4NEhvv88DBIUCmgb/s4cRnfah9+85xFc7C5QagU7NDBz5oOkGyh
0WtIxjAF5R1I/MpxRAW9UFnapz8JrBa1YyyicQ1wobppBtE34vUOpMyencnJ
/T/IamML+Qqx5G6hJxYjhBZhW2EUDNmwo5Bc/zxAFVL53lFgkca6/IKNt7X7
Edyk3zPBkxcJK6tbACrVOrWyXG6/1EflwHELqEK+0D2zNZ5nFQ6lLyj7WGXp
V86zD4538Zo9Z9MHnKI819YmCwZF5Y0GALoNZk7CYC6+Z8PUvXrJi7GVFLOd
cDZoXJVsangbPqmKx/C/UxszNfECUyZxmxqBJeUOeDmRnsVgIwoNlySPNIaK
+tQ9C8D6YkH0szNPS4WwMVusgUL8mQ1i7Tzhn+WRMHrvqIcEQVSSara78Y2r
u455f/2sRo1AxMKVsJp9c7zSg+BY1qoWkL+wVzhewZUJN5FbxDOGexgHDYHa
pSYs33FaK2KaKtpZzftjyezK8CZzZADi1yI2O2QqwSNkQLpssci9Hy+O7tE2
u+4uWtcMSwNDR2VRXdnv2xhKoMGJm/De7XjrTzRPxPSkqLSjZ1bOAsxT4qB4
HgywBZvvXv8iRHjdPJt165DtziuSVxzfmwqS+E8mcYlTImdgRdwSNfhSfNZM
99uy3A6ubty97R8JO4WML3uWLm3QWQXzgnLYJKWbGO6IFkEXtiZpoJBpDCCl
WqE5IAfdNW6sTBMEB72/01Tktxz+yrPlMCOShZbfLUf8aACsuo6Spbi5GEE+
7A03LU6nh6InGyUHDxMbV26Z3256KtoRekfFP152AajDNzi8vJqlnFTgk8fm
bMuSwadCApLOKv7eOm8sOip7VeNIbl8TNFE2blt9rk/DhYDJJfVyy4LEOzF2
7dyNOvqzeHjB6WMz3AdM0Vsq1ljtm/mlwcwyi56pmUNftILVfNzY/QmLoqfS
X2wN4Nx/NeskNX9ne4fqFINuG4ppQ/oK6kmZWABxO4VniuEmSV1ZuJb04DUm
UfGhoCYvRqz08OFqi1m1whp/BtrF12r1o74DOEVjyTJrUPRqZqipG8AlSu96
g5mEwj2vjWTjGpucYMG5jZREG9NLAa1FazF66bgVsd9F+ofpianKzO/jRwrp
qzMSNcMPRIYyIZSZ88k/u5O/kjal27wcBGaCPFhJPqp/NHut8d79IhCDhLSs
VCiv9vNjemZSzyt4BIoYKSB7Z8sGGb1F9U+1fG+ho8rcp0EGX8FlMNRz40fp
gM6k1wS9dyRrgPwAPM8PLKtaNRYeigeG/gnn2RU+PEXazaOw26IAOnYiBvb4
8pk0kQtK5fT5nBFTws/0k0yBQJjaxakAIfNoEUSp7AUGFr7H5uRAWwOPDLEv
6PMHFxPdGCUe7sldVX47ebeeSrQ7+2hl1BX5dMA+Pe01Amd28QlyrRP1NUji
hk01cOsb0Fo90T4u1CUDVlXURAZZ8Giv97LghuirNzm7LIWqG0yQCotZjHbU
yLUDXl7hMFkfxKrPpQa0rehD9QIgubTIMLsQzP9vAujMuWnGBhrp90FDEL5n
i0VPonmRQ1KvoF8to8nTyuW2N5dyHyzvQuLyJHMPZYa3C+vU2fL3vtL27DBz
7DAHQsYg1J3+JJ+MhTSZ4o95Qti2leHlLlAmnDyW1AqQJy4hfGEvog3+JbRP
UaINvDey8XhWuGave374Mf9wwuYdLyLjOnaG/SQs2gDNdqahsAcxbtYXvby8
rWU1zDN7ako5/O64HQXfSz3j8eNMWYsHS08DfIKLcEWiqcp71WdMyxhB5jKJ
cFXiI2i89s0jUzKRMne8AZTkDtebjQV4WF+SyZBG+9460NwOWPlRmO8wLxkB
U+O1rfK2sl1Q7QFzblUD0V5VLMJBLtbrT4xJf6AkQxOJzgigdV79Nrs4ot2s
rqGNYyclacLDTiTXAxkcRuZCB2NmwtxR9WTxygWPozqBrdsqpO2gVERic+Ek
0Dibs0Us0KRhDZVzhX4RGnvIKTv9vhgMYIU+1vRJvikwozLl8lmKhnifOBQs
pvIz3Ujwb7+6D28CieWNTS+SaYLIXOuqOzlZFqEFjW0MYF64qq4FpKUn2SRE
RY0k25Ira8Apy5YK/GZ36jUCGOeel/e5fql8+6d2SwWMJ5VMMvVehz95mCWJ
3RNlX+J4GbZQlQ/lZYQpd4QKS3pv0geUDJllvf4Mfw/6qdjfMR7vGiDTBt9q
ZT/MOdN4BBg2i3rmyJngC2rupREmd5Dt9cBWRI5o6/SKMAPXTzsB9/i9Jy8o
cA72PVnrA5e2MrJWg8MgQIgH8hLUNvamUZlGnxfqndedazHh5X9YMiU7/7xs
PPD2lfPbxEI8CN+Gb2cWx8BQY63os00NUH4qSvHpXzXc5PJt4dyp042uQFOY
dY6SJMl3fd80B4D/AGyOdkLnWzBu8P0SAMD13fCJX+RVJ9RdVpvojmvgH5LW
XicDzqDSOdq5Et+rb5lX1S8TQNhYRJD/NmKBhxbqYMH3rppw/wmqHFI8/sbs
daOqTkUvsiKcHPH1JXocoT/ZXObHcLwF7mt7hoYMmrnPmXBLygl3KI4MDwOR
eKHf7yF7lySZHkVVv3oI23gTB7Frhe/lmOlaUVlkpAHKsB+/Z2zu5UXzJi1M
bKRxqKACArwKzJETgLBGnygPATAe0cx6j0eSKdWlv6WtAscPDVGekNcQdzmU
xfPBYgW4yXuvxiVI/t1AL5m22rE9iydok4IkQBM1VBWx+07cMlJXG/X2HaOr
4gEceDOPEUqbB+hYF7WXrROrOPFwqyQGeyJVrzJ8k+Ch7UJaB140qom7SfdS
xZo98j0bEZ0yrKvTymaZz2mkXO4ptLiV4Dd7AjbUxhblSkxBPy3V66/9Hri0
dth8gd2IXxwRKSsY7Nf7MVkO0siy8haLPVfxs1PiHLDTGO14tSLKjUWDckKl
N1nPYTxtO1W8OwF8U3SFyIy+x7hE95/dIfQ7OEA9bOPyKhbJwBlD3Bb/jOf0
SbZYS0guBuBfbZCkl1cnBtRgGfN4nJd0R8j6CrXwdsTAXZynnY3LF4xGcBYS
LHJoLT6KULMIqwEZAPu0RAuppQspVgph3GbJ38HKeQxavxdB+/vklNXj+N6E
C3zSUoHE5yU3gkZFTNgeOg+axsUov/RCyPbR59DMwDAyn9ESBux8Co49nzxl
ukqY5VdS0be4RuAp4mWBipAvP7e44j6khCrzu8PUBI+obySpW18VvP9wkovr
4uS7CpJAKt/+cDo1JhIgPQRHo/b9PvnIPeU2m5g/Q/KWbYyZ0FkWt3sgBkxc
pnKNZdCpjKOcbuEQgPRztG6NVgMbBacZzS2/pLH1eXXg698lUzryCUC7oNbQ
F7qxvszcKZsN57ic+iXrH9n0L6at9qd/MuQoh/iURtFHlHHaldADLqRYNzu/
M/votXs7iRDpNFehMHa6RX9DUit02J/AyWEXhpy5WjJ7MyUvpXquffbxYJUy
YoQ31lubHZ3/MSw10uyK2EeAHgIzpNHjChmbbfbc1Y7/8gvieXfkHtEBqRnv
CNlezoWcg85ojuXSWZUbAyknP0bA5XI0aI0YOyMgl4U6oLotDwvSGs/Br3Il
dITsEDNmuzsBHUXlc0wJDZKIyxr49F8BUccKwLiFMZIjmHyszf+TOIse/5g2
v4RRPkmD0rA8D5Bf+b2mS+glIfnChxw/5laPk28Owae+ieeeeK6dcH0N1AMW
2HZNbRIU7hTA2zpTTUsDK7JzyA2I7cqU1UUTetTeA7y/udMQiNk2KFUR53CY
Fno5g61CosDDog3SICHn5B7ruK40zXLqtwSZYiSsHkJqhjBbhh8m7m2BkDaJ
I+0em8e4KtOlVerZd7m2bdK7gAMdEE2ouzaGIXr6JkC8PDIJa7kyZ43Zo3w9
MSmy/nj2TSLmxvn+/ODwA1ZFV5V4kMNmS5gG+qiEMWTfXrSAoF9tT79DNmoC
7qqXCj1WJolvOJI0qXWFxookarUGaz4AENAM8aaaiSb9KhvDxfuDXVFReMwN
SmUbpRyYV7CzbkmQi3wuF/60iF7q8JIGrAno5RzS8JJ80Yaict+bPiKUW3Li
k4T9OxxCxwhcVXgzBFJU+eI1j3z2mWPSOAUmyFQp2Or9TJlHwrr78lmV05Hl
d2abGD/R3riTqRk8BswZFDXD9+S5GEQ4z2/Hz63yP/fcQDfQ9QbBU7NcTmMz
7xQG1hxdCRvt28OEEF8faIsmnOK6/6Yyj1OkPxGtB0IYMFUEV8yMXDyZuotR
VMV5DgX/BBVsi2B21l7MK8ISSMveXLuhjjR9gZFUGJYKmet3S4lzB/NxINgS
MvaLqX0aWbDUwALunAuXrmkVstWbdCj70CnCsdT8tX6/ZhQMAtbhZQkfgsHK
WNXuj0NVEyKgHSRTU/IzRgej4MxrQtTatz/kAC3AbSaRBLCH+ZB8vLG0rLJk
6a1Lxo8vLmBN0FPprVOhzZql+AoXbcxrt4yrkWrWDuEOtZPVtmtjy4Lf441o
5gZVSoLlS/fwsDIdAo2wlSwoTt/Rf7h82tTZV0QvWdZ9JJGgKzY2b0DUApZE
hJ56T2S2/UlQILEhHCzJpDEMVj+YS3pPAUsAwnIl4NLLOLnveYuRkUnbqCuI
f7pwHdeCNMl+zy4vEu+hKds+gIraoY9rX6dnG5gIDaDVj1BkNNJ0ekkaLo2e
8iwBvUh5ESehlmDtxoVQ83lsVuHbT8Ha9hCwgcCx32Nl4U0DbVMwhZ9Ynmml
qkSW68K798+WZ6r/nfIDrVSSfhIDISyeuzFXX9ApWdckmIiy8HqZOMR/UX1W
OYIOFpwDbre7p4ql+wTZcWYPz6/hEtWyHbW5M+uWrVsx59q3jellt3keJWC2
UaZB2ok+POI+XN8d9Hnq+a7c61CwCM5d8qBcpEOIHm8Y3qhjFny0jUK1jtVI
F1HuLekvpj/OudKQSkqQ0fGUSUX6fHZhagPJiRECoN7UdAlTDFAIQY99YLtr
dxTKjiFrKILOJPxgktHahYk6Iun7k+82npcHvHzpkHNgl5XB5UfANzjzM6wQ
C111BKv39OgVL2qtndwdNVzv9wt4JhDZbGL5MB1VIrOQsSSE+F0v0gPd+Gn2
aFHFMgfLGtOuPbPdiDn2dXfeXIRPe5eXPHHAiHV0EcwgDHZrQs0UOMmSFPbe
dcOClhuAwyKY+sbpCJJkrfdHtHwlAocHoulS7NLBTQjwKYpXeIMxLR3LlpSK
B63Z+j3KV2TLuCgt1gMG5O2oleqKAyRBbP+ziR0GXj2h/8nsc+0ZgBs6h5ao
3vXfZGmrRrLzkaTwdJK1bMDE/ffFqgcC1EkLWLZIbsWdLnghmh6d4MbDqEnM
Oaw0SdVnj7Gh6fgTFPOKF5Cav70+VD3MmaCH/CKNVKoY1Lzps3yBtYlrqKW6
8c2vYpHcHwqsRjOH5VFSuShYDxV5SbrzoUTiwjj0DFmzUU8A9LD29AwQRl+v
iCkW4/9FPX0bCUzE/74Xs6M06lN8z0Gkm9/tpVBBY0K8B2YelyiT4kU0glyr
RAnt78zvCaRVvsAl5isMUSa9+5gCWox9OwVncxBLUXaHjDJDzxZMP7Y/HNG0
UXpUKNCRbLf1lyeIIk+Ukdyk3S4romQogeLKWgfjkQub1zQQP5N3WOI0Ym+o
RAAoM3DC2BRFKyMPUR7IPRZXiK/1pHul0XpDS/lkfw6fTi5PaKdHCmxsuNSM
bMy1f2G8O90ajT9w61hZd4Lyx2uoHY3X0mc1QMMhZRAmHU40VyP5OYwYgdRm
pVu8FHGEQWb3NrboW+Caud14fSqDux8qt/PZ13+kohBNpdPN75ZastsfyIfc
p3ZqcCuObxv7yigBh/Zk9nWoOHGqNlH6Fyt6k4817m8xgY4wLT0Nmf4GH61k
lRtiu4vUV1bZuG/Oqtpb2U5+8s/rlD13BAHn8YNI0QQ6IPgHRt02gS1fk0+d
ZQlV16YiBwC6TMjzCDbL26CsLZbOuRVVGBezOtwaddHb3vc995il7bJtV1An
PxuKZH4F6oQz36O+IiCKYbEZ9e4msJSWwZuPUnAWlbmM/fDK2IvjOC0n0xFZ
TRWEQB2+d5m/89oL97STkCcLLDRChN5L76d0/9XSFWiK55CmZ6hBvSBrTaSs
xTqYD9AMz5erKe3A+CE3iWdDWWbgJHQ35fHhYFCWRvsqUIPvRgOzmOIBxKNY
3ptTxPr2GTwRNaWRdmaQLE5dUMBpQsqpJaF+hvJ3uFx7nB0HxCTnT9e6qSfz
XPuRPMMCTIX8uejN75AcfRwpgk8Cx0KNQ0nRp0OMUj4hEvLdmYycxz6altxl
PLPqJlMEJn3bpKqGdYShmEvS09ZYAMTzUY2KKjqKWI0suugBQYi4x2F+mxEJ
YM88GRvxDF7GOf8dYqTdDtbZCOcURtFEBKpWLk+hRfReQJ8hTrD5z5MgmWg6
rxn0s8+An8x84h4+0nVrti0B8JV3JgFLCiVVuC4KlovWjvRGb57+ZchPeu13
alAiMcupZBEb33j58B5kH1p4Q2iyUOp4BgdV2KDL068c4ARvNWAVQaDSCHBs
XmVgWiqvswLON2CHLeTuLWWulRoadtYqqEOnqh/+4eDMtoC316BuJeOqm7n7
xs9mj71bOcegH/r9zKXs+spnqw75MAM9vDLHFMWfK4nwoRPMIVPF60gcfkS/
2gOr+pER75UHhLSRcC4AOKLwUQ5kAxCK2+BBBx+jodngBQa4VyF53dHytj6s
Rj6D1LJmEJq5A+dywr0XGMv9EXuHxCd0GpCPCkY22dtvvn1q/c4wO/dw1BEb
wrC4pQbHqn6my1Rnm9Yr5Epxd7zUJEP3pn0zX0rMHgVRN4Iebebs7l3ffLjx
gl9+urLXCRNTQ+maawpyeN/wLcYoNEX0IiGMDNg8FUIC+K30/4b+IqL9wq3M
2uPvi2X78gbg6tcQiM7bn0TigUPpfYxKhNnppLStevHh6Ws9C4mOxaUj90y0
U1V61DZk/cJfxP8Zexm0657uR5Wv3UXwi7z08oNlCuYxlqWwChIhPemUodE/
VomG2+TO6472kmmiGo2bG3BHx265PqfP2ki0/XsGdSf3Pp2qHATHqf9DKTi7
ElbDJ1Ex2oxG7aaLiU5EleZBz2DIA22ZlXqUBs7OYreXMKmBAFdZbRWhRUpg
KMiAM6sED7WLxuzUzeUsZWcEBP3CZBc8PxZRjq6IJmRmqWwRIuTptH7hbSlx
CQmKYFy7FHqot8Qie2k/8Lu00KJBfU2J9yMD052LQXs31WtScgfXVlZMyLMx
AOIWd9PCBcPxVE2LaLPWjQ9bd1y5LGnY/EK0V2BSJ732xhideH+9ORlyNrDN
jAq6DcpAkNwKfe9ifSag+h4mc6A82IfYJmdYqy0th36k1GkCRqhMwVcpmsQW
b3vV7KfBv6eVdeDGw2Akm5OC715xwokmyfALkwnI57nXLJCs3+QLSYWZyZJb
k+/n0oGD+8UYtNd63VNX8Z1pThjhw32WdZWOdfkQ8GoWODHu9kSt8ytfSj5Y
jqgQE8Z46E3bicqnGqB+d/SN/cAv0F5wNjjA+ORcw2QsAiGV0mODGbtAWLVo
UtJSJlzPYUuvk860PVI44Wf5p0wsUuK7ASf+tZnkx0dvv8m8hb1tYi1y/zsr
2pCS4RhANqrbaZxZu4sXf5iK+/sVsxX41b6m6TJva76aitp8LGFxy+PJQgzj
p4Npa3/ZpEvLJnYqARCrMANkKGS/tkXeCERvRiC/+dU2hxTPbO4shEV29HAS
+DhL4S0MxodHYPVn2EMfenADtkdjCin0c8qV1XXrmGYpErRAPSWCJkHGVz4v
juntoE2ts7RoBM2/Ev1AgS21EkdZBr8GnJCx5ow80bIxzfRGqp8gJ1U7yKCT
loZgQu8zVY4MljCXFnR4LpXcasd0T6UZKvDJzCri6c1Xi3rnUp89vwJgLmEb
2FDn/qPoqOmLMlAdbfbU1afdGZ8xGrgqc9XmCJ9mAqtF7dsutpdUQakxgbYY
F0KbnvABZWJNEvAuGeVPTrKy+O6aTuijZq0feVLKOHTLSKuW56hpWhrVkY2k
rCjsdntWrjbikV+mp9bLxKVAnU+/RmtyeCAy8QiPD5vrPw5IsnhMojiA+hYQ
enGw3jcxs1rGcQPfBrkb5tXcysf7OnKXFkzELORQxZ1YOCO2vdwYIljGbDyd
Od5jchrwpviTsfjm04Z/ueKFsZuk3yrvzKqDJ/QrPQJ1qnqKZDuzW6UIaBJR
Uqm7ISIoORjlivfAVrhQTsy4rWM7+19OdFbFHbflVezC0UgZF7h3yV6Cg5SO
t6V3JJG5RX9MmpCktSlBl5So0WWmClnZpjuQgA7pVu3bvb4fCn68lXUmoxBU
4EXbYsTuhCliZfqREWjBGxlPMQre0J/8z6xQkw83QRmhlb868/rZsd/k7jVH
BQcWxt7iHl/QScxqZTcwAQiCRrMDqMx3FFuUSKZTWDtDU/LZUNFlAE+YRkUF
5MOX0aYSCMGAotO+EvO1l3g68fJgTF00TmUWYpPZcpx6XkoA2qUOhn6L9CqT
/NFD5Tv4eofwz20oqB6opJ3ABnTct8aMeDqXfl59Apf70zEAzmbf45hxObAS
UxLSuF67+oFmmt+XQpxqiWpJDt1FTO4Pwvg2WDaUnXLWv8G+uVQJawdTO8PR
PF7a+1ut5LL8XeCS9KDGMs8YvgzLwsvvvgDwa99ynGhMClCcw7r/hBgeHJtE
7E1jdK1eIK/p/Su4nJbQb5kjBMDeEHzwWNlYrJVNtlhXYFsVLw0FGz47tl/V
Ks1aSGxfxDwM+4A7v9tI/vfq81KpFN56QwR08akMke0t0GuYDNLvpXrWmjFT
Vb0qy81Rf7vLK+Z25luwbi/IpmzNxGUBOHFSIpHkYSzXqVSA16G82cs1OWOU
LdRaRZ9ovPNKRIf6qZvNsOtoFR28XvHptmXV0swaBU6hO4jbPVhW5pGujoxQ
z7bwbf1i47KjbTum2Yf3t/gLCW2z17TRib6UWUNHrOpP0quQYJ03wB9F0IEq
UFt2gueahGl3fxSzHM8apZIKGEcZprzon0AlMvX+Q+DbRGFSJgqng9dht+WL
IH4UpMf+2WSgEwcRxxljFie+PIYdqflvZT0wie2QOPwGspc+9mz3YX7kF1EW
KbCZp6Zl47M4Bofx2k5N0g0YX19MMYK1Ko/pfRiiRkKodjGcV2mWzNzhtptj
UsWs1F5nt80FcxR++hwb3GxNi66QWKW+GbNxeeZ++7FWEH344uE30bb1XKhp
glhAQbnlgr5pvlS2F7S1IjgThGtZkXws18SF5Hzr2fJURH4Hh7MFlUw41BWl
cp5tfuwR8As/jPZwG0st/0gtGWH50RZWTHwNn1ay3v8MF4x7KN/BZ+WmdLnL
Ery9XoLmZpe4WnDWXJJgybLlcBjLQm+JdwAuhS1qI821xOo11TaWcgDzR0KT
jy8uBNZAMs1OnMHXqmW44PQRNjm+o1Ay9c6HBV3KpOPLksNmpUjDZDkRi75I
gSYV693F8aTQmIbOgax41oaUuBHpsCScwoO7A3G/F8NUa4rLCaNrADMbH1Ci
oBsX7G3NLRypt27cw4/6GVud0XL5JD8T4u/f7AF7nJLxvUetFR3lET63Kq0a
hLEJWAywksmT1DNvkcJkp/IqxVZWGlPudaf+7ioSczyWbt6vyYXNyIxQ3Jv5
LRmEkRVWpm3tF4HpcALxgdDpC5xL/8FGQk0CRq1b9r8KnliVgn8esFMqEHGS
v4mSwEBM1mqy/nm40W5K2voAVGiGW4FGrbLqiiZglJciS/fBGJmis02FwZE+
XcS/pDCQPZTryJdpTU2kbtrbyobuWJHcbj1JdErPRMJzYXUkZKHov/YF+qBw
whSvyGVer7LYXfWCYHXmnxAFVxBdRwzsg8elBkLKEJKxfjeldlNUsQPm+c16
AdpL/5wqVr1TqFbPjqoQml4LRTB0B+lhwEozmYisx9gLgkJzTyL6g1xCgn6e
XwECBQmLC2ytN3MdKkBOVMcpkqC0ELgnes3hP8LWdKUJhhg0PJH+87GqSkX7
eCOvqDqp/xH8YTgUbd+RThFC2ta6YHi4oID9yQhl9nXhL5itdpt6Lap6nMtS
LiFdi2/QgNtZMVg4eF8xFtFpxEx/1gjM2fIamuJ61d8DlnEXeiqYPyw7hrAQ
006XVYI4EowB2GXE6jKqwLEOg0z2KEXFrx3RMm2MfCIbxlHOC+IgGyRIyggm
wb/ORf3Lj+9okFqgCrlTWL5JdCFYk1rzKV5oaEwiEoO1fyCwdowGECcqLw5S
cLszDjEXrY0TdyaqPxm6Ie3oDn6TiJsXyfwoCHfOdHKrjd0e5+f448gB7wXd
dXPfJoVempr4qQWMN9qkzKPpwbpDUL9CEH27kb94oobLlszhcObhXaSoqetP
kbTy3NhE2BEZzJO6uEUih09gTUzZRvUo8Yp/t98hsV/BQ+xOO6qxcUWEcqhi
B6wRZH6HUa6GdRXQ4dZk8KGIecrQNi2U7RhGs5o1iQC2H8R3N5x8slv6kL9Z
nf9QYKViD/2CPnDuE2/TZo022j4/V2X5DnIbvL0W8qNf3EONVVCimRzWFlJb
vv0L346cKkICjaG3/RssZAmmNDF6Q4+mG9BjAW9DE+Fz2XpoDWUODZl51q6c
SWePT/0iQd/vz4Yri6BM62f6pBEqOwXsOFNGtHXNxfWBwLoPxTfjQW3HKMXu
dMWXJ51ubHInSo/ydO+R4N0N+QUCMKD83jIO9geGRGkN2XqdAKr+AbgKzNXa
r4198+3U9tSNyGtP0QJLkhFSPGcVbJ+GgOxiTHUr3VQ7wZTe80DbkUyjZxaf
2U9OdFNhMCZnqIkfMtRC+SO5f3s48TMrs7psVN153axugXs5Xag2c8b8cmus
pQXZYSdTxD9g7O6VJPDmyWCKEijwelasfgDHBfXg9Ol8Svnqe/wkAcBJF9Wy
T/Hz+cNaHiSYTZv3Q12CwkgHXV7YbhQBCqJQBomTceoFn9iv+hFt3cUJwcS3
sW3J0b/ST3K/2L8Bv0AgiL+yJem+KEADI61elbUN164R5vmh1MoQf2tWI4ym
mQ7uEIqaeXT8qavtyHktmlbXjUODpsnL5y55aDIh5BXygNTSAxAWe+R1znvk
bSBg49tNrX4rJ2zQBAH4cgSAgBBMRDRkxJhCCT+aQzx6Ytp57/3eAYF06+Nx
sYGH4ySQYhPoaStrxFH7cUM7/tCZyW2oaOV2P/jZufYG/8BhOKr8bvXyR7gy
yjT34rrDTWPj109UgQoMV+NSMRQU1P6aJpgtWGuB0hfYj0IsKbTACjbtjWdU
a8991vdyMGN6lBNjFkQ5OhsZTfjkCj3lbTqAwVZHz9AVpwU8A+4wARL5pq7B
uz/jXZQSm2NsTzijUpXMjIf6Xnv0FHefRgzoqexDgOzKAETpHouPBnpK/dJv
6B2Md+9Oi4slUCAkctZS2zw8GizfCXUTqE3rDbKMB3o6JSibxFAV18x7Y55i
MJE9zTZrujYEZc8Ce5Uh1P6wDmfZRhcLj2ivusc//1QBjSahnD7nqEr9R6l4
e4yBbY1Wz66WMqqC+ImynXA4lTiHhaZ6BS7rgYZH+pxqXeLaoa7OLUf5JeaT
J+d4auZTMtYkdLBNQ5IO+aOzuvo3VsutjSZQpWQCFkHvfiFXJcc2x9rEnx6f
0hiGFO8IfrwzN7gBqE9FIZpgQYx2AfKvr3ByJ5338okrWCYMnw1+VxUbPNdC
L8PNjkiOS2wjt4Ni/r8Y4AJt7Ynwvy9UTKaKC7QN2MKACeCPHQAnUfoUha+R
zXf7ov0SS/KhGXJ8jB4ET6pcaL4ZZAoGEH2nI84exaTmfFhJ4TPULUUneLz+
wx9L5opEmybjT1xrAjWH5YEWrn8WcWFd5gVgVcSqK09V8dfkLvWdksSwiu1k
JA7Nn5igwxsb6REluB9NvwQOHgTDKTTZ6QKVXLK+oSnq/b7fjsoLpOq4KmJo
EO5a7RynpwefEPkfE47tQriSVKXeTzez5WEd7ADBimE/vF9BLwgnLLdJ2yuP
yPUq3mp0K7vfNYtNGiqrJ+u4Xgs4JcvrJbf9EhJQXduNSAQGJeG9ffp4jWLU
MrJjG38iUoY3oqkf3IBhhbeWC5t4KecPYJ2CVgt4eWkJFKjR2aF7/5zsiQ4C
4wholfifx/PerCOHKGLlg3MAJ7gWAdeoACaYWba4OyUadNjqosO45R083Oc1
at7pS+JHJEV6Pzhb9GoNkenJ4IFkpLX8zAy2vqwlJIkV1VpYVZnbtv6U7DK1
eJ2bCWfejm/7WnSoQ/pxfpJYqLs7DK63+p7RmM62PRTxcGkd89GEbUOxh0ZR
sgHOddf54s+rE+mBBpV9GNJz+cvDQsGXeg0pV1ucGnUv2xpZQ65J1NMunNj0
6qS6jMjJNm9nYB5FTuCPNhjGJt2N4hEoKWxyHBGZV+B4jxVpMMk4+I02FwtX
kL3esOfvcT3gayyxykVg6yOxlMiamSkv3NiuOHv3EVTkkDYbqV/CsuZguzr4
9S9QbEJjMXsrzxJK9viTDwBsixtmH0yUkIJAHtXPzGYWrQ3w9Xp0lEJhrIb2
BdKHsRoXexak6VGbj7PJfqdDuhmaWqQYn9eTGLukJG1plkIshQzq1vfls6hs
7SlmO/7WKytpfK8lYbbD1fQNCFdoBUQbMMzLGXq8KpNwp112q0uKYPuigTPt
FFhJI/URQW+wH/wBgKBxCqtEB5FSeqmCM0fAcFwmbM9nHKENqdTlw04Dvg0+
9P3tRDl7/XYW+DR+NBefqjSHRtlECaDIvJ8uCkyhk/lLN1LldrcHbmECggk0
YFYp4xWqECSoPuYXyAi7iXeNIioKNyDSx0l754fh921wCxiCGVacTbwVJ2bM
X41F6vvh4MT2t+jjWyguun+KXWljYmMtf1GkgqnIjxhkwqp3jA3ZuJ+yuNtv
lKQ+eoBzP810L4X31JiA78/h77ALw8dTQdS7bRWq5N3E7WjsLdMX9FZDGY3q
0Z/iwc3ubTwq7pOhG/MmIgjb3Owf27oM1tCrFaEwa+fZW0LPd4gY2mzE6wkz
I2Zff/WIJOKHd5kGohdIwdcrJ4t1o5K+Hh1qZEAS/nvMw1JOijbFNgK94JIa
Ww3hGsVuwRgn1uWoxAOUCSP3q5WjM/wsuTebSda+0VJxCxgUF9WE9cdg5KLl
LdgTzazW7vYwau5yQ2VGO0QGVyHU4CupNJPr/hEWo5uDCY1IYfUqSjY2PHRX
r5rJwTRcgPWmgPh+LOk48oyE6WfeTGRWmPzN9q/V/R6oF8Mh9wBQkLt4GdH0
7SDBSfhn+dmETdMcxQGO+M7jA3DJrZ/NVvEorjQtdCheQhC8bQPEHoM7yhjx
y4lu88ODytw/TYlS7T3Ef9l1ODcEXvwLQT/OykNyQf3pNO5eBWxNwGugQQsf
U3z6iF53Kv3oIn10T583/jbPRFTPY3fpOhA5MMsHWjkMu2sxrvhCPF6/PjzP
OHp7+4stBuUwDslfwFEED9NLD6O7wEwFj1/mcbJgdV6oijP4xkdLIsKBvOrp
MiDLq+tWQ7gRiVvCWKVrzxAxSDR6SDKZPDqo/IPgNQN4DOvLpKxEywJgvUdD
z+Ih7ULdMAVtvlmKxtqmOiJIG4LzUjoPzWTsiOclL3kUN4UnPgKZpvijjEly
ggz+RgF03AHBdYGRlIkzYYcjZDiyd9RJ+c/aY/RCxLmRDJ02Bm9+2Yxn3ucX
ckOg+N6ULam9smKaeT9WXAlfS3QOynoHIe1QfjPeQwE2SUygqa2+Zlv3aB6C
Tfr38E5uNWwsQ803Zu4Zr3WShzKKwF3P+f6YTH72gp1LK74CFD8VmEv3DWDD
GZQAK5BmHtB1mygX2nqhto674xITru8ZS1ntF0epL3WpiqBV2DL2Arm1q/HM
D6blgisVWtZZh0778ZDgEMf21I9oSXM6eQsZfXOKfU2DcrHoa962+EwpKj+w
2YBl2HSMg7N5N1q67Cg8vGbDCzli2WUuVraVbPxSh9Re8B8ffG1m8td5OSHA
JF44fJQ2FZd3KW8SK3eN5hmeGI9Z5GQks1Ksd9vhdXxBwziBkiY6ZSisvOqP
8Sc3o22eH+RdvgEPMlimYX6AaWm/01LCGwygyciqd9J6/bazJZoe6TTv1Cp9
+IgQIriEy7sBhxgNcz6mBZJwDCtXFlRGl2n+GMTUszQF4JEEVoyQsVC7u1KK
iLSh4V3zNoEp/mtaq+cUoG+qdjCHjP/xIf+oa8xp08Fw2kjzf+X4PZGQ8nl3
npdYCJNHuw3xjA7oLoEWM1cfHyZoCoEaFUQB9wkMBKIxoUpURr6KT+CehOqN
KWLFz8n53jz7fHu4jQ97q+xVgIS0c5PCwsOxC6qj0hqjFn4UO2NJi0juJUUO
vHzSdjzIZogPQmXmjgVDXlFHs+fCPtzPV2NCjy9732WoiEPAAMnSWDXfkMj5
wf9nwMWXARYaDVqcozoh2wqVhSL6zG6NLY8IvcBqGbF4MEyq7aLWSHQ3wSfI
bcXuBzAfoPt5KabgtHduJARQaNlAkNzODdmdMeLcwiSZg8PU+UvJDon7qo45
44gGr1Oxa+kK3Mpoq3SfOrGHApNUnU2fGX4tRtFZ1krh1+ZOId/B+mo5SVlY
ZeFxVVinKjASNBfOOaw7ylDbvC/jMeY9FBUzFQyxYUo+msh1rSbph2RCU49a
xxKwtq14llBSgS6JcgEWQTR7JchDrGZXZ42G6SxwAYzgMyR4iAElC+Ec8GWy
ONy/Qpc37PpYPmdS3Xyiyl2UVVUV70G4qe00ooB+YM9xIJwX1aMJzMc3wllE
1F0Xba3bOp3fOI+EK1ZRzWBAKXZTpCmQFA2vr0G0pmoSdrKoYezNEc2uqkBj
N5dZjWviMaufoVicivJ9d/55ijZ6HIFtI4Lv3xvU8uFF920EtwD6FSCaH6uB
ZRBanxB0Mv8X5cZexTgawVca7d4/E6CCy+xYQF/SN32qYsjWDWjZ7JwE+AgS
Nedczzo9rHQQo4/HC7D1VB9C7+MiX3wETciFYny3JTRjnv5TzPW3RThE/GZs
alrpZkQthTxAXNj1VFZW1F3tsUCp3ezPexTW4QV7BFisvOsYZx82YnN6KwN6
1l8HmBCLbX/oTMCD87zXrosQKHDP+c8wQO83qGyRJh94x1J+IXIz/7btFAAp
bcHVLU0xcMq5Dm5x2X4Ht8GwrmxQ+mZim2YYXH1HNOAIRdFxnwh5OLb7gf1l
6+JNhiSmTs0o++DS6cdjvZ+UVV1Nxz1lhFdK6piqpcOcHFnp35o2VT8mTk1l
Ldg2BNMLMKw+6KGrHbaR4ul4u+ro65LWvQHYaUnj6QnrhkAmeptvD9qRZDH2
MwHyUIaOrSXYUDkWLefmju3IwIO2LAprQeYjaT2/rENvrZx0ylsZoLm4BCu7
OMRF55hw1JS/VJzItHlzo71L+xuBtclmv+3X564P96PNDF8dbb3+GXVkJRu6
6knoycUv61WXqrvfN4FKefsAPI98OP18spXqzfAV6YCtUO+oi2r6aJjdhlI1
mTqjp4alXwNYNSFvOdMOQ6Mzq66WbegDeezJ4pcRujMcTr4e8CPKPbRNXBtm
1OaH6BijcAC2Bw71+JoOV+x2r5LVt+tS0ZRrxlWR+cl6xuJBU1/jHdi6ZUP7
By1rsTpBLwX0XMAJdWxMvjt9ZlA+Q1uCK9MI5qKVpKniepRDwlyBuAVKZr5r
/ijGgVQ/EfbAWvRynK9EYadtoz6euXqoAsrZWqaE6KHvoKpn8xSxaYwag3QT
GIwx5FdacOQ4C2sJBRi322uSUQH6fFl2wLjDzyg/cWKGSrsTqPA3NbTjt6gP
y4kGcI5eAlZ7a1fzp7bRUTo8QOapHtFjW+4fxS/vFDpkTZSv0x3rICLckdSK
Uy04D4HGi7AoL6j49jMeHf3lpFgB3xjknjmdJO03/SuZyYiZW3Cqs3kCVpvb
gAE4RNf7Ced+OQ28FLzV4dH0r0Yrs41nP9yFjKuBS/0DKmTeQE1LEEo9CukD
ul3bj1hpqmvuOAduWv0nP9TRFfc28s2ADFBdDrqX82FM8vAonmE/ghSNKWQ+
8djKH5D07E49ZIS4vwCR+x0DGrHBKlARqrgGaw+x0EeLsv+6zo4OzLxQ3QXg
6lP4zSs1kB8+VSLq3zTtPz45rPRTOY6AaGMqWci3pX1Ri0+YR/xWnHi2F1ow
h00IyMpJzhZJ8pucldA6bu9E/cTlrvQ5qepu2Fdy2yB7+gUntv/XKqPMpcaw
EnXGkG+AKiyaJ7fa2PgfGss7Tsnv7ZtsNLB9qblWanZdtDsxKh/uQcq2lUwj
l5jpy/6QkP7bjbkAL5kAWbZ532+AMejG2TrfC+lQasNgq5Mz/3eSdGggPdwp
BFq0tpYR4aiceZ351zvkM1NHKS1KyBdYgIrKgZDTJaxEfX0qSN8vX3MWgasP
lF3fBzhGT9wFPABZx+WDjveATZg+ce7XCVb5DOFcqXR64+3tycu2VUHn3m57
64DKEksx6lbxO77rBXP9xee7aTrzn8YpyvSKCxcM+kluDoxWQyJQp7uuBV1e
xUGvh5pouBas0ErwANCLkCWqzpshpf2UsCemeNVwQMOFGlJRlrllWt4YDmGT
gpLZ0BQNrXOIYfISgvXtAOre9XvOha70iZoFWad/qlYWHo+0aQcT/a1K49rI
qGhpdfwyOpSvAOJVQoOKlmGaaiSE4kRRfDHnIDndRb7csl8IgvY4yrjY681k
/b8ryRcV1gKxF2mjDvEBaODfJFftMLNQxnVdb4DumMM1hXRse+sVt2jdpk7g
eamq7TdcEDX1gkzjgqlLc4VW4IlZSxToK6jXwKMKV9T9cHEqevwkH5/qr91u
oz6Zultbo3gxMckKMDccCJnuctvPNId0hFiaXgnYOHlZpeQT2qS9rwrEdpTs
SJW2UIAVOzVFcl1zzJvQ4eNlYe0+BtPJKXPHpRKSzragTwmCcNLixdiMgFnj
2tCPFoEvlPz7Hs7vsZDOV3wrpQj19aeTPsapodmMmgLgfidzppnyvp+D7zon
CvHeXQd8Kd+PY98yUBP9Iu7pDG0KZYww167Rqq3dBKT+P66GWUXrRMIdLjqG
0MzhzF9mGQxv/ZcKGhYlZrbrnH28enPAMsSAKDYRX901EkzE2O0yZNai/UIK
itQ88cJn6PHUoHIPQ1lcZDLxumS49znmL3V8lmefGdI+mVT8GHEkQC7YuDqc
zBq0G9mCTo+T+/cEZwuK9BeaEaTKXhNxdHDhhB/Lwghv/f92MrO2khRxEEHD
3rIZxLnariHh04Da0fY4Feqy1n++3qHpFz48ce2Mkp6U0tXm5z9CzFtlxyxg
MihEIX7DbOoQ8lTHAFzUx5QfosKVDLnnbrtxut5z67q3mjao4TiZN0xWADKW
j6NSeL48mqZejlj1dCiuQZ3QVOC4bBI2y1yW7YvRrlPEuoK8kMnXMnuxTO/M
83SUgLyYpOdj2lT4K9uXYHZeESF9TXhoDfSRV+//h6s3lDmCUUHydykfeoN5
b8F+HncekgF0iZOGWzFRqTkZCKZ68w60Fbq23cV3BHtd96ExB9it5uGydvuq
c3+DeBDU4wH1xZOgGL+ihSwz1ct9Y8LAploifSibWJ6TWTwVK+uRCEacG68Z
m30jyGVXh46r3otZJjoWOHqzcaqGc9tWhFnfUn6+PprWkC1lwhKIfGP7X3Uv
QgVVeC4MPG+8uzWDc9o9qrqm6Qk4xgbslwpoiL6gVPTjbWN3E4C5EQWRwN1U
Thbqidvt9RRbNi7rL8bd/8UCHSmHRvuef5ZIXuMVxvLHKCXP2FJcaVQ0MOuj
wkgebqQW26sAeS4+/GSpotEFP3/AdCMqj5GP0t4orZ/wwmCsjzUlGMQejMoF
5v/AlEGY+bhTvJ07Vs0YEWLSUOmgZjqK5LruW0rKSUHNU5xFeHKVAZOY7Kts
WfwJg0gp0c5ZlXjodVWeNGe4Jhk9r/TMrxleMf2oRr6+4X8JUjtT+1OZG9Y+
TBmFVrSr1OnMSBcPemGtw44ki8Xz1kRNkTw3fh4wUUohx9HeWuxAQR+yaF2O
/QEruoVKH8iH3mJEFqTYxPRgGh46X2leMVEi4dOezXCjG4OpNiEHgOz9RiV6
lZial1CwkdMmHDPTStEVxxGAWFBh2KJxvlAsJL740MSR4mxDwuusLLoLaGNq
1JEVpj/S1bt0AHYOPkm3Cm2N4xbqzYjs1GAnNrc+4yLxwoLQfHvWjY1a9/U8
CAduOowZBO2B+8lxQpg+kq0WxeAy15Jfi7lnOlisVp6+wyeP8FyqtNnVk8g5
mQfmvcxx/4DmM/DvIZlOCvhPjhe2gOGwjK3DNwDwrkBgNc6eaGw58j/y0N67
eSv3fJP90u46u93d/zWkCHXw3/K39Apapq88qvrDPI4iKgv7oIiKL/Rbt+ns
IFNr+al9EIitwWw1UHq6kzIvM0ncntBxyIEDpjunlnLWrrH5aL6YInYc4E4J
SCsyrtUEdYX4zx7PTrWqZI41kX1Kb4SKQWfU0ZlR37iQgZ/YBUrS2jU2XrxR
5CBwWP1pUCedgDy7yHK6DAvbWUIisaLVngB0eoAvUdW1/6b9wXStM1N/xj8Z
Jq3OREkUhxd/5B6QZ1F4eXUfqNxSTSFT/E7fNBs3kqExVegyCoqPcBC5HHbC
6NmAT2a7fX6uiVt6q0RybN3tnT/NbsUSIprs8wUQNMiwMJRfyQZfeam4EVfk
BKjQbh9RADaQBens3c4LJtlH6WlFsgLKr8W1sUSjpnNWKvoI+IJFJF0uLPX2
4+068kIM4so8pwgXUBQGPOFv0JrzO3HNB3YiT+McQHwueqBXLBIPVuSgQtwz
Kbq6ZZ3x97hei34y7iHjND0T+cEXqjBidGkYNvzHa/wJPvjh8Z4p6/GLfxia
N9+LhUDo++22eeZ7TIDKuGhqcSEshsq5ZT9QiycgaZN3Ed/NwH73YP57yMkj
VP6eqv35eXhdGTgy1zWanzZI1r08al8+jGItXcDXR+p0r8Q1viIxmh15Oax9
neav5T2YZd3I3mC9pX7lm5IooZM0mGXBeL9f/jlhjPANC0Zzf92tp9q9jEFV
aFF342HfPBDbKxMxDmr9bL8xKEPhul60nvL++gmcSKgi2p8Y3CFzR1f9deU4
nWGfz1RZZUx1yZyjphTIRLDWFw5qDHtXijPgl/pe3fuZcdIl5rLOthNPT23x
OjoBdZtVvLzJ/B3d1apnVRcY/TNGGXt8I5jsG3AahSAGWgHlNboK9Jp9rTp/
iwQ9TAyoyCHkmUPm+bdeGCeGHBYLLX0yqPUaoSmf274ItPKpFIwmmCrmLyz7
KfrOylPWZTF0hdomiRT4MbG08gPBuhaTiUDqIUIycldH3/bbQDmFxRAM3Wd1
2G9hMnpeaKiLAlrcuogeCdhCabGdBiKmqapt5kw9c0eP5gLCCb0a8YCP79H5
VsBwtNg77xM0Yui6MJaVChlcwZ1ONUahwHQTmqHQvRk1+MsQMIxO2vTXfYpY
qRHzcsCAZ7dkIvjrKq+yl2jxmtqNtG4tPMVptSprouqBGpVuD15ScSBCA+zI
y0Oag/EwHB8OzM78n67MdQIOPTv/64vh7GhAivfIa51bt3iDl89UN13drw4P
7ox5Cfh+fjOf4PFDWr4QzHY3bEA576wODMd9GxaTG60K7UKnbvEnX0jNphTZ
g4Iz+W3sAODOp2w7fMLcb/eFXFJXANV4sqYwH7orNe3hk/OV7gp2BQy0fZGn
f+B/Zv337P08y915hJ9Fy93bwF4cc+CYaulMuZNR9N12rU1ZE3wgcJwgytr7
KI5muzL/XEFR7w/Lu9znvet0U8ACt/GrkddtTbWF5+jSyE2ggbj+kqC+U6iC
g/otFm1vQzQa4Y7PE8JX8Zr6PTEgm1ODvRfex6OyY/S+rPDvz/vnnIV8RoWN
s7eh/yb18HMKSFz6eKJ94ylR1oGcnLtRwzLj5jVhn1b0uTLJAr4kSvY3GKTP
bF542Db/vUuNSekM9AY+wd0X/PtSRFNzq6KBGo5lRPnb8AQAb+Jexj4D9B6v
9HxFa4z5Sh26FnoL9to5/Gh/De2wlpmf2KlqTMwmI1IGfyYx3RVpG/75QS+n
XUsPs/2TIwypoqV7L/HRxUC5ph1mTLhC9aQqN8IGq+zdcwW+Ko8OaAemZeeg
0N1h9IfKFhfQU7ul45HfRv5FOZ5mVX3wjGHsG8fYxFQCuK7gXWP4vs7l5hNO
Gn0htPY2RfXPxdybmVNpJDgy/GK15qOmOlv/SoNJvAbSHWX57m6nDuZC3LzA
LV4DLR3+YcXSXzWItGZyKmNt6sjdFqReEqL9nIBv+aK7kganSIqp74Hx7Mk5
7C2qZGmsEeVu6AeQnAnm+bJj5BsVoevJdMuiIUy5hoZUszYlNYIod6rHHdJz
jogE33M5aktGkasH6EWPo4Bz3zauWboRGjQmAWMNxZgNvmk1fD62YQxjVI6Z
/h0bdtyxc6if5Byb+aPu3dJUKZv2t4hLZJsq82PKBvNj0LRa96BL89f6stTh
CQnVNCO9jbv2bCNR294qzEWC07wRirBTprd3zSKYB+BpoLpkKxDtvtT7CspO
nBqTLY9p5dV6M41G6tz2P5F9EReQVtHcDtALQsovXO/GyO6eyhjnwjv/xWlt
d2aeBERzd1zLr2uytwB8jkgexkgutIYHlLiEw4Psq+YwWm8n+9Znp6333AGY
vrGl5hz9BMMl7t0ciZ3+NM/uAg0yznLvCTiPKRsIt+huysRVtQl84tk/EtqB
5pupwBL2f3XYEqwSME8ERKrpVzRPpdW1H3ItqHDe6/u9MoPKvbrqZ6HYxfsC
SRd3C9xFdeZaTT99jRzx8d+mCh4nJfjic1OosDUBhsD95+AbeLZg3JsvuZTx
RG6tSHiJJexFWX7EEg2Pe5BntN6DaUtLijVnmVIvDRwqMQx7dKBmum+YQh/A
F7FrA8iCPIoC6/kNvPt2m6Wba/XlxxPmXD0WR1k1cDy29jITeUtW08423dU+
idtQERHGUv7CENdiy2MWt/BA2ypQ0ln6ycqUN5enAzB+lE0K7+HhNSXnjmNf
97uQ3Ev8+6x7e4qNeVnKGwqI4U/pRAUwVtit1P/0OKVfBHmj5S387EmRHyud
MoTAUvMnnN5ia+EIp7C900WkaXy5vQLECTBneco69Xmz0FDfRk6h43IfVGmv
6VBlkC9LPlF4FEB/NaR6kM9fDeOZQq8e1yX/RWDCg5EmAGxD16UplfjlyXU6
gIKcZRqoI5lAzKrFwCnjBkP4lERtQb2dl2lt1DOAab4Vbsgq36/lCmnYrm64
vMq67f9HyUlk5l7VxcAsX4J5zPlwqmefjiY1eXdaJMC/Ngr+Miuca1chIsvY
anhOkky/XHCwH9RjJIkx/THVCfwwEkifcvTzeBMXpF9EUoNxkKUCMHHdFvIP
/A9+dBQgTtE1i+Gw+cKu5d4xgIOHYxsHjtGCxnIuKKGnQJzRpMi46HztN26E
i0dQNXYfd2qPiYFqYcklMQO+tZNjiQemf7WTl5wrJKKFPL0y+/ztDK2JoPzw
XGWvOtE3OTtRx1r3vS3mPyRcZ8onidNysNo3F1UOcyEeeWsl5v5uK6wp0Pxq
FLfSpWuZFsXrNU25HbPvIPxpeaua/yAkXntP/+Fux94eA1WJdnApO3JzoZ4I
8vNeiO1VNxghJljriP2JnAUOc2IrQ/VAOFPxBekxN8aNq1NVYoEL99ugLeMf
Ngb/kscBqEeSL8Atv8d8lW5L51yZJGrIAEmpOe664JgOXywoaQWZmi5In9uI
LDyPPJhOQYZTm9WvB8aSoiEwA1peEDdOrZSl+2gJlTGp2tY5Pq2OKI59Zh40
Xhew/tAUrNRhGi5OWZYuQs4a701hrrtwBokpUvCh7qcvN0O6BwhGJQqA8p8v
uadTGHGvw+hOQIMvVISLULuswk3mQCwrR4qyJiq0KmGHwjvw1PBXYwrxriIn
JfzH9/ycIMYMtUUf7RyqinUrgLcSqx9j5wnCcwbiEyKa3RTuZg935Lb2de6C
LB3AE+rIp99w7+smS+DEcV4bZzEW4iF/gDxQstK7CYsZ7oFhrDeogPg2U178
khJx1cyHaewcagDXkNRMzC0FNwJysUXTX5h+OvG8yJDjdYo+uVulGWgsaf1o
qvWnMHCGrkSUk7sxPfIFIHvLuyoaPf4isa8WVwiIZoUdOEknGM9fS5BKuev3
g5foLXCcjwaPf9GYyokKeuv08lNx9/PMnq+mYI4Y4lSq6hlJ+0up/3+6IldY
ulM+pTMIflPdI3BoKqb7TOWGivun6C8HfsOrIdxzpYJAhSLWRIEUzIFSrY0I
SotGCb4m5nxiO8xAAvgD7JTyJT8Hb0iWvYQm0h9KJxGdManIJsEC1wKUL0je
iGlxF3rZDPUzCt0TYZ4D6MPpxw778OxikWN/OIbmKBEbkn6osishsIjEsTte
vE2R9o4kgXjKyEM1QuL5G4Xr+XXqDFBXspaqyP+6HYeT8cpHumnI+4Tv/bXZ
/g1TXuZRvSIyakhn9SdeytZe/7kYp6H27ePOwc1ikJooST+Gg2MdgF+FYj0U
0acq7FD6Owdcqku60VY+Hxst3SHh62lqzfOywh9YTZQP11AkG5c8MESMabFa
CqeYJhrKjgPwFHQaXz8kjBv7Q5Hsb04q0HLP/WAZrwpM40O8w0xffjyBDLJ2
kVw1d/HXjT3isH3t2PDU1oFaNQh4U7e14X8E6mw01DZzb5O0dj5L0hUDV8Qf
B+UH86kmfLL1NfkJr/TXFKUTV184fbXhRaKuMmrip5Nk4IPsAyB9KXUKBNy2
27E2HQXYrrXaAPuSbMdnwynfjlNPphQi1ligf2/gU66OOJE97MNETTg+nw0h
TPjCw1bcwXOesFfD5E4iqqUug6UCqbDhkF11BJsi/pqwomz6kJ56DkcA8aPX
SIa0lIqSVseBqiATpSDZGeoS9iQQQyWAOhhlUVp/zzIQpMGlE/Ks06FhNQy0
fe86Z4o3s7J43Afh5wvTFdspDzyK3LSxHEYiEYSyUA3rALLA+WxL+pfraOjn
7l0ubDWG1/6frdn8SxpFwkwFB5XPJ/6fmd7kKoP2weYY9w8QsFreS2+FXYOf
/PraUidzNw3xzSKaApchF6RXqwaj3r5lP7s6x5ee2PtH6ExE3244X2aZ8qkq
W2xB+SkN2JutuXXjQnq8lIigQdpKNO45h45sZS3VKZ1q1Z50FbtPHzvXN+Bg
OjeJS/2AufulQk2Y2wsIVbNdp83YjAP+2OaPJezmJSJQ/UPoY56eOLG8Ba+S
GWtbb/+NdZKbgHCCHqP2eZSwnCWTy7DqRMQr4C5xB6htZspXn7C50+9XPNHf
anAgIAcTDR/jBffy5kSXwN353kiXGXsHV+QofRnK3/NC7bNlEWljA0bGWuZ/
KG6x4fTFQ0fJ/Ba2JSrGT1ZY20WPWZnk4i7iUEudAJ42bw87UmjiI3jHopaf
EMpHwcU/ReBPqQufWQVK/DyZzyXSvD+wpY5zkXkQH40f1f9ayg3KC6U9jmbR
08TVJO5Xh+AaxhMDEQC/gqLKSLJHArYlG0q7oOx140+HJqF2Nd++H2WfL94g
6mf5VONi4FCIL7OPVI+CR72uE5sE+XFyjKpnewPCnkN8YzoFA2YnQcCBCgbb
QU3GkO9JsSvwhJgz/TV8aDJ1KxVA8ADzm2wi081wodJiRYzDPIKh6iWEPvzl
W1AOXPRdNc8pT0m7arm+pMwmNSN3jHkOKnePdSOG1q21udpQpYG+GAPkC+99
9b4qn1K9SHbyyDzt7liO60Tahjg83ip0/HlbXTNZY7nDExb0GmtiA8yUj0Ww
IZLwY8Rm9l4lmdXVGW0cTMeJ+nhZpjFJlsXKN5Vu8CoOMsCKbveZWvLTeNcd
mYJRdvW2F19o2G4/4DbtxmplSWjRubzlOH8knXT/Blv/ocKRA/jPjf0Fc0VC
Gdg5V/+qirt4g8aCEVc6gdqXeetu1q+pH62uXV/8cBXNvTmN8k1aRoBtrAEs
79+wosASZyr5FabM5121DUb2bQpmf2OPC/Mqq+sTQzaDCFRwVuSwhbytFntI
EgjNJmq20btcgbwC8nuFSB/LthhheiA6wywkwEz9jKgiiQlMCGVDnM/6/tRM
XD1FL3q9eqOfEs0lEJib2JZYoxIDYJtYGJvl9dzycnxA41dBeWFk4ZNd6AiO
yxwO7pSRAFrpF2UYCPw2puR2xx5ue4n5bCnWOlz1pSXxPToxmTLf/I3NXZ84
/DUBfaMJyeNQACw/T8sshq/wzUAuuISzdT8ZfjLyAtdcp/rBfUg9bLjWbZNh
HrrXxyB/HxE95Wi7pXpnPJS40r1KSDl5ORcwnltZXPP5AimQroU7T/gHlTgR
qa/LeWD5wiRGBndF7BTRNa1CwT0tT186jVk7yjxBkC+/AuQnzFrteNur/Qum
j/BXR9xk2EbrE6AGg/4P4Z/OaXjIzJRLb7fwPeXe6Q9PDJgIljoNclUOFyjZ
4zYjZjb14EPsho/xud3nnYcCbmKXBTqvb6knAxWBhOU4wNTrt9Rw0YJZjh/b
kgtcFo5R5NQg7M+apbBy0fvwbz7bNwh47/6ABNrvt3PqfAQyEpEtrQEL5O5H
bDsYF8YskTTzQ79Z8zEd5B+5ZCJHriC/cTFFHfes65Kcj1m2Vr1HbBrURocJ
hJ7yXkD4CMdtOa/RofC8cVMgoKVy5KTuaDWPam8P70ZdvwmW1fVv6ZdcPy9L
WNi6awun0Rlw80zUG14hcolwe+EyYVvTg4uAXWEfW2xKpac/Y6nSaXtcIPMG
Bvvpiv9EjdmdtXYVpJV7IIXiR7BJCJC8ec5HIjCMIXu7RvM/BYi98eRW9EKg
6qxdoGUiUZsFOo5z2ExNoN12Y6weTULtptytbAZuQWFbl06kj+krhjdnoZ6D
bkerwsFBK5ZxqrwvGshAu8LJg/Upa7t7KBbo3g/hDQc3CThbvmXgxJy4J0bF
6f2x7ayyUKwAnuOJVRkZTIDtJ1j4cd2aYk3vnDnuojM5mYd+0X+4sadTnwAW
/57AMRAeyMhbW7BC5F/+kAnrbNZnbtlnYeQjMcQeLkymoDKRVly4I+SjnXew
0xCMICf+zdr9lyR0OSzu0OZOLDH8ZEf4fFKae703Ft3sx5HWNNPzOmE04w5L
n1ThL7l9DuxNAqYsLtCMHpRkQr7G9uHb8qV3GXpL4CIO2Z3TPBLGYfqSowND
aVaaOIPRqESdxLTZd5SzVP/WminC0AyBhCx7IXdM1P+5Z5tt+E3ssSCEN1ts
jE7ESH3EZLbdp7D7IJThVZVohsaVtLzFBk9uVay9xpXw3MDB1j+9g6drWVci
d5aPxeM5Flj1+n6TnZ8n0fyILLOEt9UJByNNokEAkr7PqlEMrkHyXDotBeh2
Qo6O8QXf+BX6tzfjK4QCGky8urBTO7X3LffyPKCY637i87yze5n5Rq3ci+r5
FJvPAIrhv1pdt0BdisD1mFmOBKQGBvVBwBnYvnbzhi3Cs7xG+qK0+ZaOysn6
V/kO3YPbxwOTPn70bwR/rfIJPFRdRtP8OR2QBMZEF0KAD4epqmvMlo88mcQl
k2rdteE95Rt+NTWWhVNG50G3eZdP+ISia2y6ekQdl8MEl5ihLr0XIPDJwXOW
YQTqxL3rraauZytLIu/Ji8u/TcRGz3ZygaT26OFSPUaIx275WvVYZf+UiG1Z
LYAwsLOX/1wBMoF6LXGVRcfm87hwFIm01vA5BU4ZRaK0wzd19evYWbhjVAL/
nwLl7Tzo9wraMFPJNgzh8ZW5uE1v51cCpQor2Ow/lWLMl5JRE8+GdSeadlfU
djokXLfcKnQ7tIbWw6Ey2p1aAKAN51Xkxr5d/2xav5eMCYh8GoQP1Xf/+BwB
Ole2r9cJd+/aFrC65vvvOsIMRiLte6CuAUzQ4FBezAqwdypF90UjoZ4q+A56
bJW7kIU7OJ5AVc6D09eJNGQkT4BPIJcBZ+Ncoa9wdfF+6th+rRPXSFjwxsUp
s6GssS5zDthaUFzccGcUT/rN5AUN0iIN/rs9QyduHCJsPbi0hIs5g07VsfRM
Ep3hZjNUjwiMGLhZUr51pidpZxXsN9fgN/XBB/OCkpjFvUbhuCe1gl9MpAjZ
+tgTAnQcXOXgU+Q76zwwDnmCrMim6Y2q/9TvMNi8odksZOzhxNAVM3ZPXKcY
io+/CghvXbIqIPqs7jMv4PKoL+gaZSxOF9CGdWUrBz8IuAGBzaiTiwUONVx0
843dMiIJRuF4J5mZ+16lpLefVkQwktMf7dgrZ1/eOeY18dgLdcD5baUuguWG
2JG+6rxVCi1+pV6A6jmV/SvZa7u87z1UbhyJC3tQSL40p4gL/frSUit/jPKi
plSbXeeDExglr/KEEMRUSDbX9Vcr5KXI6XBe9RK3FbRb9yhOuwg6WGVlkERI
j8TAmM0yxc4ym/1p5QOeQTWL3OTIleE3qjxyfBA4aSkEweWhdqNlBQwk6X/J
NW6MWlcBjyDwHE49KYz+zTYEbC7fmvvP/gS1EyZ9oHbIOJTZR2q3Fxl08BOQ
TVVS9YGuJ9/HX8jnVKoWTfRXFPczIDEAnP0F45Gd7XLpv/KH+6GbxCV2SrKv
m9XAWQ9AxDk3VrBF+r6BWM3zA7D1//uLLTMgDvrmYom8fvm+PoZacJLaXOir
rdaqhXSeVfpaga6GHwPiPSryc/vUrkbX7tPfHsP5px+d21hcBeBq4iX356e0
YOcAFgw8qSWtTJMovdjhUySdIFdthzoOU7eI/E6V3H/TV4TOseURsZbBITUX
7IMBKERbqQXpA0QjSHhPPHjX5A105k/1xk/0czh7gOx6U/2YEVCfwgtuLqJG
yhcexkg+Z1APEq/a9FeuD12m53xFkJN/9AjHf9eON1f9dLDvFZf1OuM97vnN
YRi4+MeVYKgZPMCzmGoYEpC74XmUwcliYrQcbTRBYPF7PPK6La3qt4NxfBR+
yRTstnZxszHwUky65oZQM8B1oVtE62FBx9acPnrMOO/6O/kVe/R+GdfMvWLP
ffp6TalN0+Fj03hZhQMJhkww0qO2GryCH05IBvOiELf2Xv3vnr3SGBd0pp3i
YVWQzQXho4/P8SUwa/h9Z+QGugQjvi8vlAwhdNGDmW/8V/Gbs26A9QCmQGOT
khifgUtHDZ93k7RJTKOijeUUzUlC5Tqr2XAIAda4zNThyusiRf01EJWbDJ5q
8W54u33bJB6XDufzRSC2Xrw2RBRTa9yebRKs6F33LP7EMH8WI0mWuFh1pfyZ
n6ku5hbU9bcDEVXCvAOxoZ3xD7cKeYgaw2GdV2jD9aNpJJ3OWWyVAmefCP7C
rh72rIVG3pSiFHXln7lZ2R9IGdRBgid0T/QJGi45jIPwhtXxvlVw0xVB10dZ
U3914DMzKpsd+nCbEfBsgRovrVLres8cND6QzTUhqYYmowSLqr1cRF+4ki4f
TZcCwcZkSjKKvLFTnBt9WPaZvfheIvXcbRo8D1qehmV23yh3S2WJTlD6//z8
eQXEn2yPGmJ7Ykwpbqb8XbCIgOYHT0hUU/D1yEhbjadiBOC1+EbKdy2tTqog
MCGXFjmzhbl6Y6EMbi/3NB6L6kjsPTTUwCtC7/nyfjxFPadI8AOnXw7294wM
z7MySlMXB9dpOo5CATgNf7lK8MXxGucRI9pn5YGORwIYzffceuGCdle2cMax
OpYxSYBsht6HKjELiu8blil4/iMGH/IfhTRrnflGBWZGgslKmRviQWvisfh2
dwH+UyWvJEZkniZLrMfjbyK+Qqu6plzfVPcM066L9Uc7ziVDLzYRUiaGwgkv
KSQm7jVUu5CIIziBy/LFYXechk3etiukSX74rWKTJ+gZ4CyQ/59NKUHddOBM
EqajXEInM1d85sVbKUcDae5Cd9hPEtoD1zi6qMv9Z/HnqefDx2Vr4+AWUEKc
Rv80xUYmPQlDWO62jPrVy//SQl4rUN47srGSWooZYE4odKzkx0BHsQzgNK3y
LxfqVWzMEC4WMhA9JgGZNdMB7A4BrXLokpAr9AbHPGu5hrns0s0TK/HU/siA
oh5U/b2MEgWSwRuZW/X5X/BaMSw/Z9BxkTimWfgvy9O/DHB0pCU0ANJ+Ugp2
WLYuUBcnji2sAdJVfjgP99+mk9POf4t0KD8KwkbgMbb9oNdfmnHcjxLCXghn
fF7hZNmzgm+rtS+AFLUKU3j3Lck9FDpJ5zdMcsskatAC7b0PoY34G5zPCooV
KQx+7oXVEiDMcpBC66WEL89XUvvMNu1JBj5tu4ofE/YzZqm6tNTiS+zM0zek
Z/FNZ7TVJbQG+A9JX1WOclju4Nxn6FziN78sl+lPcQV54Xwsawfis9uyIJPJ
kvlNS9t0aq5CZh6AW+rWkPl7I94uo45/OCFxrjEX0WjVwk9AEE57T+JOWQYj
sixFoLTzv5mnWrm2HHt8zRr3LdG7h6E4pGFCTYCSrlXfjOXd2lx8zkyEC8br
nwt1YNqo/EnLOtr6eWrSNBqL1LRuzjSUZapVFZeU1LBk+VNT65BLqjpfsM5d
Rd2rO5Ku8brdXhOnaP2uZn6zZ2wDVvHIt0D/zcLdOzUXL7j7z00EFZLWFQn3
9k60kRURSJcSDExw8pI/TWAgRSOZhc0/ZlmPQP2tnRlBTSiik8/BQLm35Aqb
bzyI2bc/Gwm6VRVv317qhV42FjYIZZok4L/kYlqwjS2KFB5O5jgNQJqowLtg
IdMZbh6hEQf/LQ5QyskswOLaj++4Cu0IdNUJpRn3c2BP+sQrHyUTBUwlUtTf
XvRR5UcKZUVAobkKqP3E+Mg7I8xQdbyjBJ2WwLsNlBKZTTtdR2Jo2SadKnGS
VukAUXpEMKA9OtUh6I3RadGjbhVBUMNTaKPmxQOe/rkEkF4RUfb96IWo2A0/
f8ScfHEePvuDagTEil2z+ZLjTDqmNa7kflyznXy+Ai2OmW5TPRtQD62qtPUZ
eJsgHPoy2UdZwzivKZQNS7opDx9oUMI+anw5wqh4Vtpb7G+/p/8jBsZCltyL
YmvHmv7ecmo49j0BfnSBfei5FFzs5gqZZnaGNhMBUArM0RDp64Ww3+SaL3/4
uI9Vb/qgZBY8yLlb/bUrGDjtX6rabV3fNva1FWMgTYj1XUtZpZgm1Xv9HFzj
NEsCLitBrNlY0SPYx5iQTifO3PHQ56jXv/qCiexEsxdtOjZPVrYrPEzhNqzf
bUeMCbAVDyi67xfMVyiQf6GfDp8kjgCk/8ijSYyfW3YnL53LL3W6i02sLU/f
xe2rC7FquiZmHb363DAPEOEiFOAQ1qqkhMz2YKXTAKUi5I4kQv1zg9JniGQM
WMVzFxrH4sTwJSJu4IhtFvjyH3D3ZrIfO50fcnoSnMvE3uOwYT/Zd8BSMdgS
KzVYX2r9sgMi+vDUd/xSAY8RplBDW78M2UWViKZSn6RfCnO2mqJ3AQkKgvg9
zvqhGrC10ouQC9sGY02O9/f0zmmAGHdSAgUUSw+N4nibb4Erhwb4Q+lZZxLi
ajwYjj0AYkl0dE9VeeBW0YFwyv6/ul1E83KWtW0f1MaojoVcz2yo1BETkti+
INlNWPrCtxflcneP7vm+grF3/WMkJFpmPD/jseWCZL2wWyFb3Hu/7tyhzgeG
kNK6Y9nVXp1VwRuwC8MM7nIPphNNwaVK/m0k1WZoeV3KbP55U/cvFHrkk46G
kUdS2l4TvyM47seVjJjh+qy05sYQGxKIRNAslK2FIcN+EoPsCmvip/vr67l5
wawMzuR1ITboQVZElwZNj0G2jy/anx+QSaU2FmgA+m4vzMf1KAques6BHy5Q
TJpVZVKUU+1PTbicCogyn5xHYXMz/2imkOKTPNysKM8kfq/dJoKa2ZYMg0jy
J4fblHQaT0gSegnDyodQcpxplgW7ivNoyKvGhfbCEBiP1LUYyC9mjBwxeSHb
wJ5fEB4o7yNIHrhPQrhyxc8ad67O/o/UhjDSeqhpNTjV1IL+nO7mfyrqmPrw
mdLCgQ3wmNLA94jTcYUblvBEhStKUUNZG4VHMLlw9NKUHkG4R3zZPu2rw3fG
a+YS19qVtW37GQ5buLNlpam2ZqD6cwipriCafYm07bcfU8hAYizgo84aWNmR
tU5I9ki6AnCzx8q0hj7gmX5d5o0T4OZwF8RX5odBBE+okzEMvcsQjZlYh7t1
mC3GUzBYwKv1M3SYr15Rh5E6P54NW7KNZ2TG3Prl0xf//SnBQf+DkyqklL/U
tsKruu8Q3Hdgibh/Ilg6z0phABFtvXPh/2hu8iCGnnL3HiZduEC9huhzVoFw
yPIZqU+RhJ71/ZsHsuaDkuRVDAOiL7PEuWafkRg3yxgugROLDBgAyWLl0whj
KcSvvSqHrBBZhSJ03R/MwLlrfHHXP3mWC22Riu6Kf+9hFUQVdtfpFKc82JYA
ZQaKguiA+Q06ybZpoLOsWq2muuBsTM7hIjqVVO4B5AOI8TZIv29EQc4b4GEH
CWbWTNqavNjkfQJ/B/XNiVeFyQR0TLr+I3gVLmNQAGkH2k7im99IEn6xRMbm
Ffm1t5YrenS3SSv39qiEEyjFWm9sUo3qJv9yWws2yjYEbEmdfnFQ2SlMIp7j
xOoWJf5ZXxqFTzdjYHQTUjB4QBKb7q21LU5bOTAzQQWOf+p8FnbrPJ3JB6/d
GHfCOBR7b+Bc1xSMyqLp4TxNRu9Ww7pG5GdoWbY9M+EuFoSXOCFHZAC5dvx7
APXZHZtZ0DUOhtUIv3IVdchOIBbIiK7EDu7XGzwMACarAcGop2rQ7nKzEGYa
oxzgC1lXNwNO7s0ZpvXK3vysYDVCTPW2/WHjrREW2hoUET3+scMlY3TietHS
OmNaiKzwskX1FQ67OTYFyFANsbUhkWVHll06zkShU0FWmuz3edp2OX8Mhbtc
A3LTuXDMU0RmiUZbGySVOXRNGeYi0qTNjwaDtwnldPTYTJ61gtI2EaGzB7vJ
GqQYX5whxIkzjPkIYmsLXkJS7azNkisCBqnoCSSxTSd9nSX4fXdvH63J1aFI
iADrLnM6NdSdxNJzQjd8QYpr9EekXpXfejxM0VIGGBwi39iLPRJstusUtTKd
MSedR+Gf+KhsBJqNpPKNuIDOwcm6vjgYKPRSZpPEzsxFuxFTnGy1WCebkK/b
zm2AT+xKhWiSVK5rOpPULXafp+fskqy/gC77acYTuOAOWP8ktScsSJVreDtj
fUPejUYLGp5thr/44YmhlPGcBUPzbqlEbrGOqFlCJXjW0FOhtFe+H0AHS6os
JfPD0nU2j9AmKIYe1ZHgNlLKLjxEQF9bX76Ti5h91GvAk+H1qIeJmSyMqZlA
dz7Cw/gkOl1mToGw86c7b5vv59MvJPe7DwU1k/d6LIjkf4IFXFoJmfDzjTwL
1Ob+I5WbPev7TkQ7Btt8CPoC+nxz/7JwDhi7q6BzfHg5j9pf5qxpq2GIOPxY
PCyt/s2udAdU8uiGwZPqwbTbq4dFzWNIFbPsIow5VikmsGDpU7ZcbM2ezEDl
p8xlZc1vaSm4nq27MVfbjblLpUnTsNKfoYU8EdS/zAS80fouOl7XpnhS+CS7
TqAdLTKrNhiL9/yvV1eqFQlFljVxNVqKIe6RjTxscA5A+c26oy4k1InyEl3n
IdyzQRg3ja6EkUbR/t+SsQTl+VSOi4lfkorImnhr/VwEwuwCrG3642ru5ZN1
AAXsb/RIJr1JYzBJCE7zoO3wdeUY2PyloSC+eI6htZ4OKO9oU4Qqkrq4BYyt
xbaK26jdo9DfY8agl3gKx+MixS849LtXvR5LDUv7xxshrD9wjaxdKorKqV+X
1rTG/L/zByqNzW6zbeRGX/OFS7Ekeu7Tva5c95oBUOZHnQFgSWfs/JcdE2Mu
LchzyNd0eJcK3KDY4LprUtTSpbwp/w4lHXa5EYJ288zIHN8zVv9RqMSR5MFK
R9bDW0ERI64kZg+1ycscJibPH1ClkMvFmlJ/JJYFDa32jghPaHxiMddjC02T
Z0hBDVhwh91gEE71h3jn6k8vgftQbmyDcH127b+bkB0weWggJ4XQfsTMvtSb
GaEQug+G5jN4yzt7z6PEdZh5Kf7VG1FyYuZIysuvYQbRrFrCeFifAm4Irw5T
iI0gLxQDVD06k00XuRo81nFaUlWNNHiIFe25PJaySE0leoHBkC5f1pOtaDLs
0Dz//quOzVOf2LWMVKHdnu7xNuyqmeOg6eDcni66pbiqxoH6TfM2AYDmZj4U
phbnU0qml9cA5n1sNBCpZFzpivDJARVmdVcGzggHUduYXL2EMo8N735Oiknj
KFD6NaElmkAm/aqy+4fFR5BImqOsozW6U6+Z9p1vBaFGcdNyf7P/uOP71pRu
5yZZg8JXXsb+tULlmW47tuSarJPy9+Ivj+Thfw8rr3Bxg8jusjwefBeLL0uh
5sqw8bnHTDux0y3v9TTv8MuCpJv4KYHZo+nT4h78TKdfGtUSVPaFo3zJ8WxC
SY8ONtLvMY3jiUvwsn+oWnqn1kIrUh/6+6KpvcFKaD1XYK5euLj/9FwReKTx
0j/bv4oH1L3JUv4NLHdCRqSm60NH2aHNoe2ckl/XRU8u2bw7qlpeOaXfX1fK
wg8qHLfjTtrWCSC/VkA9oJAkkPPhUb5rf+6GEuC4rcwk8ggL0Apbl/np7vXY
hZApY7mGVK9wMclSU8WA8HSvCmEndoXeKrokcvcTRdgLJUzvQWIznZdBQey5
xlWO5P08Fpds8KE9pjsgsMb1TBhDYuwVYAy9oiYgCJ1kvhlMNGT0tk9BITLX
EbDmp6TY9A3KXr1ju/zmoOYojRr6NpkSYr+E/pZBssUmk4icNr1xMMYHDnBW
LIlQsZdEEvg2UTmmf7eDoB1zmKKjWdMVciKVC0NRC63dkzSfrS5UE5D9jX6i
50gI82v5d3sTjKBpiuuT7lv/NI422+BG6cjANlPVDPfSLXttRPCdbyaHBOXU
7xaotf1zqdzO5X4153+vMLLXQgJwHWEBlael7DHjz6PSQoJ1flbqRcVhH0NP
Ak+4o1Hj6mLmNS5i0V2an8t0UH1hf16k+sOFci0IPrz7DeFkMHxywYqk2UYV
WGLBSagMgcA9UV5/jarVRBTGJTCy4B9aFMRUV09teHZ3oDyKqqaGT/L3WxXN
ViabNKXCqil9bSizXDROZKi8ml8blGfWECKdODCwIFwemN0b2yQIuZup8FDZ
Dg1F4HbStpTL3EiRovmNOifKUOjOJXCVPtjWkco47Xg5fMPT6xNLH6g7Bfle
42BD0AUqHvEb8mk897BNWOruqqCDotfSQSvcXrwA3LEQ3S8b6lKM/ZTt9RaA
u8m4IQejvxysdFGTYUMtHNAHGB1OLooLlWJlngKFtrc8uls1btGqliw37Qb1
eVn7fjt+T6y5N3l7XsbZXQAYNm/Wf95XE3NUknDunG22hbgUUpv/bE25fo7D
yyiCSVuxiAj3+2507GedLDSmGRltgZj8SkOcutz962m1XaOnQSDfjpVX5oF9
pb++RzoLOLRCrufUxor8BmA3Perk4nPgEZ1ajMzMi8sWZyNz8BdUlaVi7ied
Z2qs9IFIk1g5CnLvjyTg9t6FBg+DBGlerv1mq+KTauYL6tdi4d0Vg+eliPge
vzOBWLiO4byJ4GUaWDRNx33+Dug5m60T1P6TwqmrfI84Ws2xA3jpxrEKCe1P
QB29xawlJDn9PtY85cAxHgBdgOFqOJJYYQ1oV0bC9j6JnYHhVj886MikU6VB
pn017LKhNe/0c0z99RY4wOrUDeaXBdTZPBG9ApkRURbtomXXewT9W4spHTZU
bN3vfW0N0iKQu/te4i1wOJ62VqpOj0c8fEOpixRJpENuA3Ym1dCnu9Wb+G3d
4U6yfXCOAs48hBFAAa8ZBgPqSqgT1f8dJD3JEt3U1W5oC1hzLz6kopvbfLXT
2hGPUtbtbkdAWpLkxxIsh3bmnu9MbjSnN+4PFgggN780C4GRSJ3aylhNHCaz
zMIs/6sBFhDmyL94/NW6huSiL25eqY5vCHf26zblhxVTVm7UnN2HI8RrEitB
QlmKkONsdR4l14P/tz5IQGp0s0+CRC21aN7j3HYz8TABMnQ+Xfculrt6NSI+
AVoE8K7+FFJaXGDG2Ifxqk1PT+gHHNilvPv+/2m327G3FD2kuFTZK57owDAV
+yqvU+NhkET6+4dd7tskAoLlZ0S3D6MSxs2lsmOZvP51Kh4afKQg/jRtZnco
ffNO9bbggp4j3+q2Sn3nikvsqubfAlIzwbGQERCczdIDkUyRAlX8DdaSPk4s
DaaoNu1KhD5C6fZ634Jys3o21qvmNl52BtP907UKbrAUYzAWBhA3FByddVsK
pYUK4T79LNa1hYjdvjn4DTC8yXW6/e4AZm/AW/8i4QfUL6Q4ngd6YME3QrI3
v4T9+i7WB9hsOCIYVhIFFQ29lYsxBSP+l/ABOz0lDkxyRV+X+E8lIyXYCJmM
8timK6Cjtg6vPv6hyMsuFAe5JCo8kjTgth500pqei7u65L7C+K6ovwNa8UfI
cIJmDLalYfwHL7GlrCEg38xcpi6c3YmcHRYyKtKSpf92TMam8htprleE+1VJ
9eQCvTXy8RcIlH0ZuqjjJHJhAe0sTeZ6467iHa+yUpPqZD3vVlVtS3PSmEGg
ZY4oXhbuB7MXxCSToYc/yZV7BihGd4c8VUKY4gA75wGjl5xQ4hrbvFwWDvGJ
niXez1rp4XL+5adbJc0ne+GtFE1Q2Oiv2XNScx6Wy2jKAq/9ZuEZtQjZtLcx
IYnYG5R2Cgrmt7ciMLnUEx0bNGzUMGgTL8LC9h1Cz8WQvzFW5WYWWG+eaYZc
CNYJHaO+67kXAWbVLuzQjKeV8zPgTZjbDVyhm0lrYNNfwHat6goaC4hLkdJU
kqwESfTL0CWgHM5EIdCCz0c7ATTQtBKR/HXiBIWRFMlHUUXF1wsmBEC+MiXM
462txFi3mtAfE20fOtT3Jm2Gg/rNov2zwlwnrRAMLOPmti674KF4PxRzyZB2
HrCrp+u9FQa3M/QQXbG3veVyl8WNLud9tKadXR/mdPq9A1LUwVNE49D8veNr
KruUxLuv48vFCLKDHk4H7PznzKLJ+yc6Ybjy6T89N19jJ43KVFi2mFQn24LC
Ja9x7k5N5xepdOjL8X9lWjlGQvbxwuh9bi1l1VSwdjBboAj8N18GBBHAE7PP
xdWzXUiYigVaFq2Tem/OylZa6PRBu06/rOlYb2cjN9bTkKPcCLrZdMkGRguN
h/00vvZcuesKxTM7Q0GQmJE+Lyonh3NVh7tji8ejXKGv8k/C+dD0zTEHzJzU
TUNSx8u5ksV+jPEosPGX6XHn4qgufF+cLWB3NzRJwdiBblaZgZ7ZKL76u9B3
J9P9MjrnJjs0IF6D+Vq2dkJgYSJ7gUQ6bX27opeQ8h/eWKJrSv1jOcJi6XLs
JxGSG4nwFigolBa9InpW3mSUIjl7wr5U2vineSdfi3SiB/gx02ponLAvClRb
YTpMHe/5W1kYURxjtNNDsV9WRY2nXkQi2OhgOgCX1gH6luiHPuHWHqpG8D3z
54jBJbzbi7kPzJW/tz959HTlbfSRQj9NhDJFT4Bb1jLuQGn5HDncGNXKbTqc
M5HYduxpAlVNRsaILfbwmHsu9wludf7UIqnEQ5vC8VktqP+7erj9gmGfMlJU
5kVqr2nuUxqD+E3/g0Kbet8yduwIVOTFccK4zHq4FK5unajfyZ4Qi0qs7c5A
l5K+13tHBx0cVGthixwnw6Gre/8fGKBWp1o+MLnTnkU76bG+7ST7uWb4C02t
xSihYKbG2GRK6SMQnmwUc52QJMP2TAvlWUjruEl/JmKOL/9FIzikjC/Ig6pk
luAHbadLUuK3qR+Y2lHzJXii9/B7Nz44NDf/5IaQWyN5+Jb63+WYc2FIa77C
6aohp7yK6eK53z82nghK4mTTy08kVw1fm8GbE6ao33/P8Orx79eLJda9Mko0
q5FxDQqvXtbDj1M6AQdKMeinGDcjnlLCbcv7wZPilImQkOexOw5GIcSAko81
OEZAy3UvqMUnzsxtOLo2aB1HBl7EHw0XRPwMJM+pZn3SxcB8Hfj66UTBlD6y
6iaimOjTSiqa7s4pv2oAswlYl9Nrdz+KbK5vi12fh9VEmcGZ94IDVBZQ9bqa
MC/Q3SV0NO1t6JG4uoeFCtLwCOjf/unoVmAJ66DyvhCwVxfTe87j39TV4tmU
VjVw8YI29Sndwn+FFnABuUG5mr8z+/ujtTlTQ0w+bGOeU9KlmmW2SIKLyQJF
HQEQb/hBpfqIbIVWAeI8Z5Y9lAySr3gtopdBNLnlFgIS2KPNOQ5i3WEi1Waj
qbGylrlFkPP9g7895yCJSfY/l+sVqY1CBJqwsFTIo9B6JRa3zGbFf/b+w86T
e4ueYwncogcijpXL2qGKOV0Y7Xdjk6mEm/+KFGjUUsOI/qT4fYcTaFk6s/Rm
s2YL7YiKV+42Hh7aOX3CuRgqMNzBpvAilLxVVyx5P/SZ1bfNsgX4GsjlTGGN
nhXz/zHS2n2yN7Qnqtlw/75MW3uPlynWeQ1MFWxw5zURGJFnACP8eUlsC2vu
BTarinPK6cjj4qrO8K7llNdTEpXQq5GMfwQIXFfVBBgpXNQJjUGOJj2yWLK7
njF6RFvepBX/ox7HSaXpLMr2RgT994oMCpQ6wicuoj9+WBpSWliocSEzidEI
cx065Kcjj31xuXkBUBZRoqhZoLLLXmKqNapMjf7pM2JxNXYpALsaLDUw+D6O
zSILNkXrjvYkYVN2F/hlJgOn8JjgBmiRT0/PQwFQxFO6d/kIaqmcjC8MDXv5
iaHMH09rkcb5d+cYIjaRIbJ9+83q3Y6U7KNF5mQdDCv8s90u3wt3XJsWz3J0
CZ3DjtprHlscsaq0lKOPy83nmUigA2Tc2npoIKHT/ByV2Dhu/oYaq5APka31
U8xj2tpxwRPZFRktEFsaouYY0+c7T50IqzXBmBGifOUycH9qG2Yglvc/lWjI
caPiYGPEGFCUNjYBTIosuiyeoobhyYCyHYEnsS2aSPAwof2sw9vlkJNe59o8
+7HyQIZbcUyLkDC06lwNkQuBFDbEzZyo0H/+W3ypMvSIh+T/2YFzyCGPEy3m
zeP/g1r4FavKWLpoWvqt+WApmrXhPZTNdUtaNTTFooSCEyfE0DK/k8AAz9tw
err6MKFDc40vU9ahgutfA7IDizdaPP5vfqGPz/bLCUOIHdsla5alJpF1VRGf
nAh9O9aOvY/N3E0NUoaspZ6r0QaFHbZ+snO/5Rws8h+4KWgWQFT+699f3THp
/d/imIMbvxTnTC7JQtGmJlgaUrbRaAEzF8XHVSLpLi/wORORS3MD1330IK2x
CCQFqUAQz0lIU4D6o+Lc77AmzCJPFnp6bZoaW+1JMJIUOjpXWb4/lhNOf6AD
ckP8RjsDe2gdLtPl6gQYARKniggY210Y6bjfCLSselpAWaQtEmqOEhnVAYe7
lCsncWGsewFyFJ0/VKyGnuyeT9R99yMaMk4Ze0ihAWGP1+AurQWt3TD2OQfs
vP4BSQ95DQcF17DqdDLYDiCSGtfRIt3OsR/HkvoxFYoNrj21NJbhbsND1mnp
h+zq13gTR5yoL7AVd9zyKpBCTRATJ9oPeGvdCe72SW0bcEnYdM2ST0vXd2JU
SsWO2hYxkEzA0I2MR17F3wHOMARddFLEZqsjz15TZtjDnbz3nXuKrO7jHpGT
dc6u9BjdcvyCSEm0hVzT4UP2Sm0F6lj5xvewKwUuPTkej9IlLxkngxXdfWBX
eBlFresHisp02UFoOgTS/AJkjhOJYVDSkvN33xojX+4QvDjqrXKAXUTJhNHv
Sr6kVc9/Bn6pV5rMkhod/44PFYJ4S6PLXiO6wp605b9ht499SnLRRVbnhkuf
TnL/nfMzYL5pOBQ205Wd00qaqbFDnDSsXZ85IudZE3culgDZr+tJHoubq+3Q
pthDMbYH64+bkNAXnDWL5Z6Va7cJ0H+H6mOdofp6Tsi7/yq0aF4FSSWK5zTK
KWbQj4UQOAOneyAsDFuMHsenrwWFOP5wPnS24SDzgA5ImZx4cwHVljVUkNfX
FSgB1j+sGWavd5FuWEXXjRC5iz7NVg6VYP1hwyp1WA38qcFVIX9dKURHLZZP
X+oBcMYCJ6h8muk03CG3BU9wky4Wd+j4ndrjQpfFO3/32UkjQSBvet8CkKoB
HZT57AHoUVSQTUpe2vykZ4Vmts6gym9Ie+2t7/ISdu0V64/Vz1wfxcnNT9OE
88YO8k1PO5C+omJW4RgAYOh3u21ayaTvUJz+4T55ZyKdfrj5u72EPtUSHita
+1mB6volRanlEBIj4CQuNrsXYTx4c8+0TUnrEzNiwnA4ORSAy1SH0qjQ3+qX
+lxtz/hElTm9uJ5FSrYDS/fn5h/wgifGqYa7wBCRnYLA7yqokbaWQy9gF5VM
tkc4Zsy4w3DENVIkQ/1FJKohiEG1GTdn4pwXcTuhEJ+71DT6FyCdLmAiTOGP
Oubjy3LxUysLO5OFdPWG7CpajY3sr72gtkUPhA7UU1yaLl3on6jC60s37jDD
dI8oRCRcRJn+6X4i4/RpzXi/ulBxdeFqGZfixGnzUw+KoW42e6S7VKpcd3tM
QJwbdU66f+lSvhqAIS2/Ae/DVPblbu881T0YCatp358/uo0+ITofMlueLlIY
avHSdIQaBhTzvLKr0Z3jTrtAv2juS6Mmx/DK6RNAfWIwwuj56ok5usGGoGYu
EXo/v+DeWhow5uUs3A1eEVQv+oFQCd//befgJ0u+MbtXGXtHdihQ5kaTyqNu
scbcsVkAeq2abzqMo/SNiQyaVykE2vsXMnyEXDSsQHBzIx2/yxMIEvIgtBbx
xXoY4RF+R2Z/N3S/iFba35WooymcwoiFgGsrfopnSct7LWDoywfILdj2mXa1
5OEPMeSJ41tUTBkelLvJob3R2EZp+QIGdw2E7ZJGd69qPZwqOr3D7nqEqYue
Tlna0l9WUZLiffjPTCCTNFeZzN1BP+M/Dqu8D31QVxkLNE6d5IoApQmdVG8s
U0PsB9xu1K7MHu97QDDj7opzEciXXzEg6bvjR0YBZlhWld6ghh38CuSCw/cu
D7+z2lNWwD880ACtEbPDaW8VQnqckfgcxQypFCDnlzB7XVAcnNffUcZwJKSP
ZjkmqcDKPeZbUps4IyGUORLkmogmPfR26G50FIb+6RYz9nHbE1hvvsnd1+vR
2wsDK18akjf6KOQsH55bad2M8MDU5CoEmPw6GnbCWls+EItGQ2j3aO5c7IvE
dyXzE4VQIfHI15JAVnkIxG3JA10cjVIAr/aU1Qti5a8GPTLk22KlNHNCI6Oe
ava3vxjQw1UEz7M8DO4xOWl875YON4JoJunqF839giueDH5KHXklY/M0t9Dj
BqVNmfJ6bmhuVDZQE2GCVZsDwslmMzMROHi3CdWp2+MpkfQPt5TIrSnp/p64
mGvcoJoQr6E6GBlCXXK8QZrtrnzmKwJ+0VL1CQo55dVqFpQDc6tyhfY4pgQU
bUS+ZmSDDJR65CxlyEKwy6OWz0iWh0E0j7IRF/yi308M1qkBhWb79irljvtO
cYRdsKmvI3KS9Tb8UACP7t82n81Sx2k4kT3VFQrnAkkMzKduVNs0rirx5bxr
FVqPvqqUFT3M1yseFdLgxK/VJ+JLmoBnbMJciP84I0kh1g5W70o6lzQqn5Vo
kqupC58wJ2hcTrguTg8wHxUDwMWWioqDW/ddnCYxFZHsjERiPq/4OEiWCJAz
6nwKbNiFZkZn5qmjMMYLeX+ilyD9BwpPbjw0JFdrkmSFmZhmSZiZZuMh+WNv
eKAJCbvo1p5sHElC//NeiardPvCHb4+MZCaVc6w/T3z53tuVjf/aOizFTR3X
D3KF+mzl2aad2o6qcpvZFHqfkGzf5xbAEQGNGl/h85LpM14VmkN8mXXydrFD
NwIhlZD+hOo0vsz5foOZmYtBYJh/bfzfdrt+UX5irOv3GTHD5pwtV5oj9Zc9
8qSnV/aKiznXzaP9sd91fNKFhCtsAMKfipHY7vVnHEOjoK80MFqYUK6Lz8LC
t9iZlpa99yDxQxmiPA85QQNuRinMgN3PHqP5HYIAYk4XY8oL8JfkraAI22tt
kf/zoPBFvGxfiNsstPt5zJ1iYUyfeiPdsK81dypJYrp8qUMGCPZYnpUVk+Ww
OSeqqReX2N/yOuLHHDG1XZFQe/pur+nVC9/bPhDEgdJZiSFboCCzNh86JWek
i5WAXznAGQmIOKbB0k24y3hu/HK38rLMN26tkjXPJPMc+4waMWOnDCivC0bo
4G19kbrVzi7ljZEE4eb3ldaZPrilaRWdZRSTBGtBd2NUnqmcQLc4umlVNFCz
rSkSkEmBqQFk9khXYMA4gsyAbSWCn2VzdmuakH5xja3BfpR2KaAObubzTcYS
Fiat42DSWSwgP4j3CRGB8MuYj90ScF4nHJNOa48RIF8+BzSS2zy1j/5aEnqR
3GPAK7AY9p6BzKZnULqs66dgeWC612wwphEgdEu1VEjUorw87syGq/u/ju2m
oO8aKoKbhKKOk6fLTirIRwb6beNCv9bJ67xIi++JGrT7DSSpwmRH7E7VZqzY
xoxLAR5iEK/oIJYoalsXdm9NL+H05W8GAqHtnMlzcScX6y3k/EUhzWwLdAlg
DJ8ijJpQtLfbIQtREPZkx0omZ8d6s2/psreXeifjPP0kCKyVFwJsUycSdotI
Ov2t/dNrd1gZAiJrGlNe4tK8/bPB1Sia18iAPQmQxEFK3yh/Bk3pUwkrw+WT
qoVLACnG+brvPnGy4HqQp3iKk7IoufVr4/V35unLkc41CNx+FmiHlmOH+0Nw
IkuEP3FpDSZ9tsLBP+EXvcYYM081wtwWhIASnAVIuKeH3Ghbf3NLfZ+hAtgK
16S35U7WKSaMsxs81t6d6IeIG9Axz3MgNNntHCovIN54cI2EcK9bZ9zWa6Rv
NyfFBe8ZkaSFXgu7mXGpbFrQXschEi+b+ii9lyRkCBjDDmnnEzuYzPlzwS2/
jFIVbLvMRtMZfzYrT/fZVL/E4dyacmYc/EC8OYttvMuVyKakNd/ien4899Dx
+8coVKPYzSFvNx7y8kJb+LgdFVTOAnlGammlja7/3+KyPYLy7uQEeojStiGn
4B9QBRk9CgcsVdxNyAc+4f/ghSWIyl/Pc9vBYjhkEDDE6s3OfvosD/sxPrqu
nBdz6Rwud7ZanrKdUqPbSXEONDfDLcOtf5JIMX1nlUT/zrfvlSEDBQeMzQOc
rCDacCMTXjy5stZU4jyXONz+zXhkYmCzZ3JRRqST1jKk4PQSgicaU7qvujD1
5FazO2j48+CQmvgJ1wNQEQEq5vWY+V3/iz7cuNfihoGUr2niZ+1PxA8wtLDl
DugpzMLfZBrRu0fgP5qXj/rQCcv5KSW5sk5SfL3qsUaKKDkQFJKAO+QcFRNU
RNA/YKE5QlRGBJLlXWGDWOGuWN/6Ka1nDdUEvfgXrIGIxgxfaodX6Kzuo5/9
cRo/QEYophFF0gYtEIgtWZB9fdoqPYlDdMQ2IYb/cR2qi7Q/IS24+ulEOnl9
x+1leaRrDgeBka99VA7OvwLkjVSp+5pcgnMQrv0d+PS+T8AU4D+13OtsVbgK
FecK/fs1srSe5giWVrlaA4UY41jxl2aMflo2T72ZpgJA8LG4XAyJ5RS11oos
geXldJ5QI4imed+dzVLSKQ78QFqDB/JZItgXKrd3CmhI4PGBzRtY7TIVDk68
/sBo0h04/k6A1oVnnrmhd2GX3o2KLg+J0zeEDFsJpJipOj9d+9nldGEqhSiW
LnED5ytvgOCwVbGLPS4bOxE1DM86/xzkJzPoG5evJsWZXUF2/pWwjzH3jakf
s/jFRNieDRaMqyDqLTXB2Pl2XPSsnNDcVR2InVZGC1nele/DbAAl40hUiJRq
OycWlcc61kU5VbqPLVmh5TJKyCcd8OHSF0h/4/zEL+QxUSDJh+qlPSNqvQn1
9wZJz3t4ITCkc1RNp0rkOsjFP/NvoztGrzrd8yUZ9kba2JYr/QoL+/jLYtQa
gXpwzbhKWas/5ja6QeGTATLwQgUGHMp104al7Fa4wYfVVzDLdZngYsTt5TQV
vQEj/Mp9QGkppVk3wdAkise5oOEOc/+rpkMpt16tAQK4YhyQrsr/2L7xEIai
BPHFMhOjypXbXfj0qkIiG2upo7AoC7nwLgtkbn7T6pPmo8YGkk3CJQaI7HTc
rfoEGSLfl+Zs74rB5webxlmecuQsR4aDEtlCeS6EH2mn4dQOP0wiH9J/7y/B
UkvBY2YFSF9hU97TOfYtd3XDxKoyy+dKEK0jEub5iYemS6Cj+Aq7gbmORdYg
yLhfWWz8954hTVdn0aNBqmA9ZD1gdBCK8U9hz+6HzHfPdm/wjw8lgw8TJ+yE
vHprM5UouOe27LpDAmyh80mKONfpYnoRsMrUERIEnutPH7W1YhHhjRdAVRP0
IKLqvEOmOcAMePJLYX7SD9QEZPpeg5tVcr/Ze5LajjGQ8sKkYREJNveraLU9
m9IkWiWWRNnCN8YzryW/E9xgbQqqJrfO+He1v/tEJWlLzi6D9r6nJR2IvUKX
bKLUnWBrI5EZ+qMN3lyWgWbEbcOdsUCuh2v7PNVi1OrUZFVFgnenAaZapNhm
wLqPDWVZSDc3g3DiNoFivmNspFwJ+442hvI9W4TKW5KWFriDZfpiKOQz5bNr
+7EctEm1dEfxjT9S7LUusmAi3SQbcwfy408ugV7gbNMhFPuF0VberSlSv330
dbGtOnROyh0rWJkDw47ZsnCT/w2XJVsAHvfafLQ6RRnMknXtHJzyGlE4+7Eq
f27Oc5UeaSClAh4+gsZ9hdIQ4sy0QIU8Ibna0LnAyCGiw+Y1/03fuhja63pm
rB8NTddX5sFmntkD1iME05ph5JuceA0FjbLkq3FVeTxKtJTe66UIbbHmrVQo
TJxCo0/KKtW3Y11TsCfu3idx6ZU4VNTzq5e0F37lvv6D1/5eI+dXvobniaSw
UO4IeFfEmP/h108sax+yG3YHRjv5cBy9U4ULKQs9nw0XtQzEB7bsqIrCA2cP
mTVRL5GS/FmvPsjVEvzjj2ezBGgCjtwmEYyLpyK0y1Ko7m6I1/vj71Dbd0K0
aru853VD+GLk7jPXzrGflEjhapVczjGRyaHakRHlEjm6yJX9fbpw3+VKC0g6
gfxUlasZcs1moywG5bEYy75rN4dlgG7qsA6DZqwBe3g2v8G27Ju8Ml1lIXA7
SfwhLhyZIFKUEs7cIANj/KM9dpRlvFm/KHJ/EjlNFX+dprtzmNMfAEAbXEfJ
V+QJPE+OrPcP125e8JKfFSFCgBHQZM7h2Lr6nU7VyGRqrqU1cBp6vdwFVr0b
ZCCNl1TicLgapgBrD9NOd+SPcpMloPvGMDAtkrj/DkWEtJwkYCrwncf13o7e
C+ScQmAsds/4YkahHdavjTM0JMHR2sDlLAv9gUO+4BzYY+2bp/s0+is2bf6h
Gr2mL1p6K7pcbbesujFbqhnaRuJ0JKO4EyG4vA89GRdQKEEak6+SK20+3xJB
thWxlmVJviUkE17xIC2aB2q7+bqh/v9G8Zqd5Gvny/H40LL1fgTkgcpWnLWC
DdmDgQXWvR0otGn5F413aIroPdF85EsLOSc7sqB/1iBLjcZAOS7zd+dMCETk
f7CaZlSTcGE6FKXjFHrcShy6eoAglLJkyYy49TdYSUaNtHZldf5J/Xvo5y6A
uOKPSjkF2tNXx3F2Gg24JrhEVKMc7LoMOMnASOxHyscs3W9/iPxzlyzfcvro
uXBymqjofLvVqRQsrC2IacSasd/k2f91HMRQxGuSd6eMTurJWF+2oj55gJX8
FSefWHSVVZK1ummDQQROv6dlHTv/j25BqheFaGqQIaKogishXC+BRQRZ9qYi
JCYN1Ozdd4wyr1gSMYCC8TCIIsJKA9x2wKfzslVptBhl6H1FYIN+NBT92Dmj
wY5AEmfj671IqoYLbIsUT6NBDspHkAGbuXo1ZgnlLSe/9EZJRKMvFIi1QuuP
V5a2qa9M3wkbHjAZ3t5RzdE+Gp/5lO9ejv2sEsP9kpj7XIXuuFYzJ7jaMdPY
C61tnZHR83WzrbRh+N7tXI6PzJddSswAO/85glx/Fbm5bPh3Ne6c1t2NMqY5
RVrcwqFOo6FkO/Ytzc5f6Ziyzn3F00LHRcz4Px1A/88o7nKtkk7/L6dBoJlp
bSjKWAnyWgEGsnhI/LJjf8eygE5CR8HBe8PaAaParogsEQ1kq7OLHaUcCsL2
lzPnresZ15jYb0TI2h3FFrscb9DMdvu0ytiX1+VFDzqpZ8ljmYVGjHhSx0lm
Y4Db+Ip0YJXZ/S1/u5Mp2o4o9DPBGCi3Y6Sjaxm7Fickj6ahvFP54C03CmXj
4lP6/wRwZet/Fe2r0GOfM+lkuXq2CpCxBJqoOqfD8Kt3Eww73y7PnqDTKkOT
4PowLE8jJ96z6henaI3sTfGMVULM+PFBuWtks6FEPL5gl2bSLMApaRqwBPVh
vaic0KRZF02oHD2so/q2axPvKsOKvdOmLl0katSU1xgjCGEneb7u7tcYnwvl
C0frutRrOUFrL5Wj7CHQw2arHhnlBi383RM4SJNBHNQDtmR7tXjF1M1otlJF
6U0MyoGb1p7T5ihXAThev000RbttxDksqxPdk6SbXML2H7rxkbc63n/tmdHA
ZXCIck91e/27t373hz0pbSAKAlOrE/W9G4aY1Pue9FZew9SWEfwKuNpTHojf
PxyM3kuOCRsP9Ie8NGmDFVe+oz/i7V2OqdTpixN7yyO+0YYihzpwMZfKkpPw
HCdR+de8HWvM2lffqo28rsrxtb24IWuMCLYGgnOvcWkI2dvhp57wfaWoOp+X
IE/DSB5o7zAO5pmZv5ARZjFXnlcnSxMHF+qMwEanAT8XNaQUhPb/LVo7/Gh3
6Z0eCYzOuLd8V119LwprqqPBcl/OURnVe/fC2JcDuIHw5ROVivjHGGNTmKqP
wCrlpYaXQqjZSy4ehv3Nb6yANJrbfPNdUfTBSV45EoNjUdbp45nly0u0CjTy
3T+EzVmk9SQo5ExMR2BoNYbllTdbLa5KXI8Fj9sHbKLeBom64aJr2deBpIfs
SANGnTZK+AZ0hheejo84aaDO+evOxSlbxu8FJ2/HAWnRn3OfgGtnk1I9kvuH
tLfKRNx76Fum9G+ixTMkGqxZupbUCWpWOnasLX4X+t1lnHFqMgce3AYOinay
3AUXZXO0cpjfD+XzBbMfDdas9HiijMomKrTJlbzk0kv2212ExhgEQ7KzUY65
3oRm5NP9cKOw0A4jdsiU0/FlXo4s9PkLCymDhk1OIjgvmCq0qTmfXEM5gQml
Ch6caxfNFlbOxelMBISBlIAuG4E20jNly3SUfMW95bM8n5dhLSdNFtUfkfja
dvrZBZngEDa2PHipgDdVZIFpjQlMxj0/kv0Hj/TiJr/w6Iz65IVBJcu4LXRO
+ogrH9KxJyodaG/jSM/iFIELB80bRo60/TJtzUpPsE8cWJdq6TUM3Pv4UMCa
KeDMnk6pU77nMq1CFiOMz4aPtjdS2GRwjQIcvQpA2jRhizRjodidWx48ySeM
94V8GInRiWEKRPp+yfhgUeHhoHRuK0WY2GI7QhmDyAutYCxuB+T8uav3e5gX
q9K91KYN01Hx7GUY6E/SnJF02yvWbo+ZKqn2k4GDUm3ZBRIahjGGkOXzIDF3
gBW9+G1akXG9hEN54JgP0zy4NZCeN/GpfwdUWjuATJMjg0dF5XTRxZuv0Vf9
58HATTcXEw6ebXkJ+LiZvgoQZue5O4QV5Dd3kBUTR7B75eiJ4nzuvuVnG3x2
Be5QktmkztnMNTr3zKIbj6T/5J1+TMkYm+LfgpBuDUOEpPYOGxCj2kQfRXVE
80yAalMS345cxxZ0PTVswBjIKR5REGLX54kxglz9BGPEX66vxcLaAjIPcH+1
1HwpqpQ0SavM3QrYnxFFy4fSmfWsNVzqQxa4+u6kZ0rwI4YX1v+Rix2JwsqF
dvB1Bti3HBxCkOe803SrgJ6rqJIQPjvmb2Fokf/UtqS66RLNge0+jKmAZ/OY
Iw4i8EjFGJixyj1Q8xr5Otl04e5687mp2wwmP0DecSnNKN5XUTZtlj+XFs9X
AlJ4gQglRAGExNy/MAZF0s3cBz7C1ecWmXpRb7W+CeSFdWNq0OZr4rqnPKyw
qJTXcRYKRkrs6uIMw0QwRJWg7gCwSZzFQFNILj59yWJhWv60oJV57qf8KL0g
NdY7NENCmERh2PuJ8LSLPlUEjZV1TDZVXYR1EPyYaYLC9+deEM5/pCodpN3D
eulXu6/0V41WN0CK6eyg83BSJzyysLsDuWTOOXDPAy6fh+gr8wLzLu23n2g9
Xcw3zUZsn49XqsV4omQjkWemh3FDSiWzY8vJev1jfSsFH0jf/J6qCQnp3wZ9
Z0Icjdp0o1BY76RE8EmNW4WYDWECQc44B5A8K1O1SqZQ/91j9nezHMklnYrS
Vn1SaXbwTWLmV2daLv++/HyQhk+++l/lnUvjc6YG3NguMvV/5JWEodVSo5oU
ShpjWQrMFvikME7YuHnpRfhWBhT+BGuto2NPj4TAqA8zZhQ2+p2D2Gew7iS9
xEfwEmavg3fynAKKIxl5JfvVOC8T9UhDuonPc2xv1/eijkuNC2pHS6P4E6w0
+qDXQA93QvMrEDGrh4QFFRoCmyarRzLiqWLK4U+KXItGj12E8ldBOAkHL2qs
rySq+jQPAEKF4rRlTZlG5uQN7gsoAnqTsAsdLpdtZARGKO6N04x9eQWuRJSU
0CHVP9HpuDSspulKmOj4HFYsAKimKwjq8r9G9jTV6ioVKJ613e1xYIl91+J5
lvcKpTcMXuUyFrPaQPOmLwaIGU6UGQoFKQWGJIdd2SGzQ25jiOhv20dsVr+c
bMI7/FFmT+OvE5qWCC/H6XGyxSYdaFicwFrKUCZhHG5t39LC4BeEFOvBH/PL
ZG/jicJFRM7DOimBvQQDUqY9yMfn0XwydXyqreeRBT1u8ECP43FMzeJnHLeI
/H8b5c6+dqDrY/V4fabSP47LBVSXDQyViwxQBopQZBS7Wiga16t8TZY3/P/P
FZc5sZZUKg5Ub6f2bNhCtSyVZopUv5lAH38tZJDm1z6LQjGqRO7D/e3u0fTK
ichhN28/CSeKnYLvUEEyaGpOPNP1e5RwCh2YN82iI96yfD3I7fik/EHHmOEg
5sht4oMV7unKIX+5Gv2/aZu5qvjGRQoW/ThCBwrt9p/j0FlrcNfY8WvhGP31
oOz8h2S/FCG6Szl89aeFTIBEU9E2C19YmYogjd4/0z62qH1wQ3NjJ4noJx1j
EBySyIBU8lPADIt50Jw2P/1RKgaDF5ZTLMrdFWFDWInH2ISvKbo/JzUfNd1S
KmIp0fqNwkSXHHQCSMCbkn4N3EEwhC+Om/FPhOJO3XZ7nD9C3zE1hU80CqTX
6nVIsY0iTXEzXDn9XWnhYmyMXPRnNw/C17xkpafT9yOaSVN7ovnI6Nio9o+2
5bmH4jdE6IhZ2TVy8EnfyByo3NnDkLRRnHZLE3kO/qQHdpFymrqo+Dav0Dk8
jmO9LL44h3/bC+iRXeE7OMR5L2J1wH+9M7vM5N13HNljJeEwXwRn7wEeHz3E
XuOXZNMNRLmfiEpR9gAR5npAsfsaJ2JB0H6E/pydzou7BKHrHYeEOcVfPPkx
vTw6Xh6RTUL0x7B3OaBCyR3QCfOLfhD/vMsdA87xT+qaj6dLbwUxXqgLxtOm
r7Qq2Yu9USAK1hQoZZNB+dj5Bxh4MplzYssOuo9g2k7+C0Y/Cc13TxprfEas
ygXINva1J/NGzIk/KlWbD9FiIpJfpJQuAM1F3gPA5aXUZFFKWnmtvrUPcrr7
HxP2QuPEGz8GvNdHIVwIcivB0T8XQ162vcVDDorcRpXOczsC3uK4wCMtAsVB
pDXfwKUAFKRKFMEpUqCOT4qSA9KtJS1UrSj0OZLkhYo9oF+PNvLnZ1ca+M7O
lwA3fkuJH6KckH/wEaQ464dC5lFBcuwxSzATvYAFtYoSj6aHi2f4CoqHlJln
0UQuSd0Vh3atSwTnW2/ht/GGmkyvDptpjPQ8uHODc2ck8fvtZQXnQiKC3JVp
gjNvF5Qnndd6qO8nxuhBZWcP5t2ZMhyuZoPVOqM6vJ6L/wzh6rX0Nci30e86
w6+ieDVZ8W+m4EDZxbcGlEPJrO3eCjCEEHXQkvYrQGwrcjm9OFP1l+9pXHlT
wFG7to0RMzzxv6D1UI7NbmUaj/PCBrXOeviWtEo4vEiKEdCgR7qplBkkNgRf
zRlgzmfVozqK559qp4YNujQSvBk1bm0KqGbAFPTwoaAUsA+vISkjXzcOuHp1
0ACiBwAeaKX/zpyMSp2GtLbPozdEDLpherFJ1P/z9cJko3XWla5jcqSgiVSv
rpBgpzLdlFXpE1s060ZUQ9mI51Y1vbjYbjBOvVGWK7dxmgwkpjtJIY87nrtx
CWGxo+ycDNSXlMgucRErFOjH+p7b+xnawOoOq1L0DNQIhU3LaV4PPTFTHwk0
WsOjfoLKf6TfRmiHtpKcG+xae+8UJLhAbYz1NEGy8f73H43tln1BVKxVsUg3
SjE7QSbNQn/g3MLt6SulZYBRwDjrhaG4K6rw7m4haC/bKz5U2bfhqA0V/GTF
+TfSjEXiWUIOioQFc52fFUbNen/sXjKb4c++A7UrRFr91qupneEeDtGeTxc/
uneffCV2k35lZbBBsQ+8lLHx4W+VE180mdhutIJOU1hVh5mqSzDFHocO6vEB
aluJdLjS0cCZE+YvBRLBN7te8ssRuzkmqH6m+6bOwmDNhtfUYqcQJA70lmUU
dfShpXOc8g06i2gVoF6iuFX+POsEJ4JB+oY0nj3R3SnM946IL/nH47m48kNS
bHkOuFqvBZ7iC6P4TCfvTKClPMTOL1bEO1IdIT8sAX13NePrbbhseFoA6H/n
bKJaSo58AsuaD2TQ6Y3M9UckiXSpWzf1UYWLHbOxfyWi83Mi1LawggVW6pY6
g2BPrvn+NY8KgvzEIVPLnsKoYtQuv/tIIrVTXqw1gG6F4IP67rCdKIrQ6CRU
0tWzVfzuuZfAOszuP9Sl/8TYrPw9rOc8v1ibJjYPr8cQcP0P2ZEAgButx3qj
X1VmeyZnLcf2lqBErNp/E9ndJqaJAZGty0ChiQ3O9JxuzuKjTAf1UZSnhdpx
TMpeeJ7bvmMP/cCr9MdO4xyO0lmpKeMrhl1iZkuD5gcRk4Vuni5yp/HfHtT1
Hz5Uloc9prNYqLJhaLv5kqGUCg8oBxPpfTvZ8wuI2zZaaRgibbtKTJGG+zmQ
vKTjo8phfLH9EcJHiCIy5L6MISOipLrBZRQeI8l1ZvIXYDtHDfF85WG5qFzE
jErEPpDehTI5xyY7l1NcGL8XZXjXCeEqtEtW6TdKLrGpHbGfJfWyX1GMDQ2p
vhpHY/YahvnDcu+RxgiPEwGUA4QUCslATluKln+kHapGH9MaRQKo7LYRKMMy
o133OH8F/QprUuMq1bZ1mnpsRME5wMRZw48lXPcFPN84+wRgDBXHeYaBI6oc
c9qrJdfnrEQxozsTVHn0TxzSrCy0ZU9GBz1FfTbz9xRQo+gqjaUdTVVpox3J
cqWttiG1qco/oFh+WWxE+dVGQvdh3uo3oFqDHwlCk5COQs2BSGgwwFaofxWp
/yR8mQzuxS5owuxbjFvMXke7IEhNMIBrC9uKuuzYd6My1WOXfPszzqJTD2MZ
9x+zG7c1uWhusb+FMQ6Th827NXNo/ReFCnfeJqwDm5+Uy1D9iX16m2WH5kat
gZwjUvjQvihClB6bLA8PpZeyE7uYl0bXc2HKQpaI5VM1IlVVmdFOrJvjmY0q
M+bL4VDUizYhyCv8/I59Kk+ugi26bCHrujeV48pus2lIwtO8rMr010/esCNL
7SKm0jZ2a35dWCOh8oCnpV2IrT3L3okq/MVuo8hiJKPOQx/eNfvggP7QfwLA
65vZEJChZMjSBZ1aUYb0qJX8uKfDziEjCuQfGda8BTkg1RDsGc6HoX8cU3Ij
R4Rptwjh2QAqq0d5Od9647F7BKPCtrVgDspOgafh2kkeknswpPacU+EWDU9x
JZ3eieeWJMRazDud4OUkRBlzpqaJTK2UiQJ7PvZexevs0pGMRU7wwbvBj0kn
z3gICdzyjaUzXGKH1yVtar1JjmaJZMZ5/fUmPeBCZUzKww1UrqXhIqHz1m96
iHV0NLXn107xshtvPVlF0/+lODmUhHnGcPWkc1IGLJYbD9MahVhYFDwnsmkK
JdHg9Hbl0hSolyF/wjYIMJNuiTkAPOtuS6PWQ+2QAJP/BJpX5A8cmw2zw444
ZhAVSjceHnCoQJo+Q1WVxgwDYdjI0ze53OG9WBtrPzch9G8zd1VriJkvSaae
0eLBFlxfIQJfLRQG6l7FSeLBHiDqyGLHYMf+2AbQ1/eqh+IMUA4bxChWeX92
KhWGuRmIqPdIKeV8zzNdWWyYGSgoWxZIEwGqpVwjUGQbTPQbwE7odukW2PlB
8zvsZiYx2V/Unv5O7ZI/SctET+xQj2Pn5D8afAjNy3y3RHECCgSwFrCsXGcX
Bt+RqO7yBy9uvnMbRhbeRGqtQSLX46w5huRYN5F7ChG533dWd3QIjN8nmwkD
YSvNzX4vk3dGH1Q4tWrDamxp5r2H0GYI0B+oc6uTCpIp7VjLTvfFZmjPlH++
lfANrN39mEvhdtpzdwb3uigmz3t/EAiA8BtYwRIPQvYBOkshvmLFmxBhauDv
HToghIgBuxnjjMKx2fXVtVWNtmE4cMlhKW7sq+hX1fuGAiy8HXOgtTN6i7ad
R8HvDxR4ZG5YqUx6yt9Yr+epV4tCNZqMbIraGZ+IlD348Q1UsyKy8Wrx8hvR
DzsvtaCz/JtA/uskQaBnTI5eRXqGl5POsJsdhl5XPQzXg9CNjzkCTLpNTWwM
y538IV40dUI8/JVvxIgcb+CRMMbE/YpcesYutJATv9rzLzANfd2fFTyWvOBV
hv8yQbD21PVIJ//wAZ672ymIbmhDSlIcHiyxXEJkDPs5fN8MapJfq/6LxCbL
tD+VKLTWa0F5AXYNy9PXrqoXEm1NNNot3XaFQ5fbklp+XpI62iCd56WviN/F
ERVM0PEsqwygW+SHF8CFXcj/mEu1U9jVm8U86goVsBZ9ZfCMAuYHe+5mbavk
26XPDqb+/dHHkuq+2HsYLvrOz2Ob9b7m8vcwOiAM+e+n5Hx7D9nBhzyPBWb/
0faohZP/o5/a+hFzv2EuN9Le8RV8sF/5rNHFxwz/PjWBy+/XL3GjOTl1QNnp
cwAOa9jZr+U7PjGFCzeWim8QyEcpytCKGdMy7vpRky/XUqL5yvZH1mnLV5Vp
Vnrs6/2riaeUcu7htbYA5xXtMmXVnbsaLeCCs7FY1XYYccK7XNrEuN4HyCbu
JPe9V+rsOj3Ho3f3nULBx2ePq4nrwRFjYMNS8qZjLSMF3Fk+TMkSxbTy9Ndd
f/3Dey3HtL1vvW9Chy25JFcYTJFYiByN5HdS6SlPrrnyttbve8F7JY61Hil/
hXlkx09UxLZ+Efhh9kZdsL08X0gp+43QBlflL6aewKICh40MgZLwrFi0GGyd
jO6WFAZJxPLfIf5RJt7PEXN0XdgrYUx+wzzNiFXGgW4fqyldX4E025025Zps
BLMEYWD1UVvqwntRJ48NqVsN/vwbquiktQ5qCawBlnC4xEyQ8HYM28BKQ8d3
u2qfb/isohPriV1tRZ9AeOCtU4uVl3X+9uBCuwTOyP5EeqJRjt721JoYA68r
x1SbSwb+kUq2qh61gFvTDsAPwh9Y4YjVvbdGYpSrkOzNx3LQ2I6gtTDp1G5p
hb+KLi4L79srrZFTZ4IbZcL0YamI+YzfOwkSZqcLhq7EJ0yitIeV9d8xXkNI
un7Wgzy+ADx1Xd2XyM7ejkMWrOw12YhixfCFM32siKwsQ1EKvhxfaNqBJiYH
n6+w5Je8eMsUKBw5OI3T1L7BkZzpuxOywvRNkLrs0ng0GJZyk1wA6FL9G1vd
hllP6ns5Gd5f1+6PVr7B7vN3dPON/Yo/QpP9j3QBlz/8mbiPXVfVAhef8TVA
Wr4SQf2tun02vyufpgA11PUzIAF+eofwowqN0VeydXMJRGnNOWTnY2fzIvVj
vZixBBqPOqu6JBnUrfBEVCfBVZyv+0foZQzigOf7UMps1Kerlykeg7O8UCt2
8tajQOtgTcSuk+sO8iblwstDWTL+DlDTaVTIGidftGtMNYfMuw8QVaVyamuo
UwxOCYyHys8NiBT9S09M2YO109JwbU0ap8Pij0TEDfJbQuAd/Pgyk4LiOFpX
8utInS2EDH/6Ny+TUTcaZdNsTlRUkdMgXkul9Tco8RYJdt2vGajuB1wHHUDw
XEogLNkRvQ2B0c/lSwPiUQoybnsTVqeFcsWfJIWs80yqWHVo/J9hguNM71Ex
6o9L/0UgiKlj+yKx0LvkX+mEHVC1W4hQjaDWyG0m6woJ1eIceWXMJeTeoq90
wiZVoUozKHuXePFNib574FAKoLrWbCK/+FG9ByzJYdQn8Vhr6AMEEXrpKhdk
RGspsAmx9uPsZtYnMcZA9Uke8ootLQ+HQnJYHgoDh67ZIaBaOLS36N875PhL
Xm20Ir3G4K+RH0QgBUxB45TpVpWYL0hpQ6zCwTEwgEdurrYv4r6NwVgjxrLm
K919+B5BgLO8gGmylrUqmJvSwlf72f/7XRQtIlvgQGgt96NC1b2lZhj4NipE
XfGdlJs3vGMVn82KA+biskBoLd7sm3ydaoDj+ZxM9uNGPDl/ZNz7s5xQm7sy
zcZWr8B4ZQ5Tdyj9xUZkw79INnXFQCevVaq9mxtDb/CGhvv34SXqittCAe2T
b0yMnzLFYyQTq5MrfkbRjHGdzcnkXrN0k0JMxMxzAuiLlLrk1VBJ+yPI7cLG
XNspd+of0hxdaXYbiF7+farkO1YPd+MM8rsEFt3CgalGTXPA0z6irzynF0k3
BBDrsI1o7CnUNvnoYI5U6xR2q4jRbvdUPPk/9VywwizGoY6uH5eUW4l/0Vg2
EK0sJuGsoBXZSSAekPHefiiovhbuEBfojUAdc0Zl47VszcaWQ9khdUszQby+
ZF5lSf6cwsyYZ//C7sxebMq1xOfbclnTde80AzvRJ3IhEz/2/82frfj8pkAc
1C/QE9MScbM0HT4X8KglmU2NvzqkwlvdCzCc0/ZGGJKMkbqlHs32snZoueBT
XawZp9R7NkaisHIhchM0atw5k1wwTJ48BZvev9Qnp0TidY+LhJ3Hd2+b/bN8
ClGruqUI0p//c3U/1ESA9fqNo6otf4RH7oSmg/1bFjZGe79fs/DDgdP+fbXe
7HdSq/u5ZoS1pC2TL/bV5H+RO2BzsY35qbc0l1c8pp5mUzRRZEHz5b6wgX81
v+crTf7zv1bs+in+e/K1BNI03oQ/0q38K4szQpP7TL3xr6FA9Gn/O4Yqs7+M
W7wCbqAtQoQwhs8F9ZbqOXuPveBIMQRMRSpVdIHL08wofY5ExklSbzKU/Zov
GxjG49ryWCyr0B0VS1uQExvJH9qSsbfZfxPy8/otTBYefdg4otNI+CvU7XpY
RiPqQ8JUbq+tCNZHTMTsQ9f/RcG46ZfeeGW6phqkZhDe9tdFq3fFUemT0RIk
TDBPjbJS2E6+0BaQ7dxSTTZolb8UZHvpf1XzIgx6mg/2jONz8rcbJTaw8FZW
YqKmTIMKku5nn8HPkd6r0rWIDSnKKpsPNLu+HwAXaMJ+dk8d+9iyFOm2rHGN
bGL6eIa6QZMSjBQmDT8dIi/y1WNATX+vrgNmgXJb58fvHNdr1a6cyTke9eQO
S/8nj80hQ0E4O0KSKo8vw5LRfwm+C4Yo3M7OprUbGVHA8kNg23Uq7DquuD7z
n3l6/6+sCh9w/Dp/Z3ZlyfWAXsuJCVhcf6FjeZOKBzS2wfvLkHr9HNYwVS79
4/LDONkuDtwvABXm/U50sPOnBco93yLygIBT/HtMLBYZE2yUWMM3HyX7eQ9o
gmrSDPNwMRcJaS3gJXTmLkfbKFNVMShQJNmSRPAtZZWuGtzPJVZdoYTWbi2N
8Ftj/hw6zhcnF6ZA8ykQ25hMwcaSsqUUpVUYwdrbteL1xbgLAPBfQvXC0suR
7PnBZAfmWHIN+RBUsHdg5yBhOq3J25PawfhKD27ih39tVQhvL+1BwrQRyV4C
xPSRP6WrMDb0ZA5vODBZRckEvMF6Jym/7LyZRXP8Bm0lC6EPJDr67P7AzyPr
VmWOE9IEKZeOsrg7bao8IFi3fes5hDjJm6Gj+CoGvidyc54TNNqy5+1lAv4d
CiJJ3lXxU67VppBgSAb4wpNY1+GuAq+wsHdooLHSAdGgRJ20AWs7tzLRGQGB
byrh9XG9ChIIibk76pLRn5d4TN7vN2qUc4AIlBgXPEMnPmpRsQ5locYydNu/
b2L3hA6KqPDV9gCzQAYXUVfQX1x1uQa+pAm0rwtnb2hDRl4XcbJVDAOG11pj
paa+mz4ca5cQa2SLmyMkSZzmkt1Zjprzxf+TTc7YmnVuZ/6Kx1XWuYOPImdQ
xUIpSUIDlVhMb7hSuoag6q7gHN8Ub/Y3sdN+t1wINZW9ODqK1GARVWDHfNXJ
gJrkr6zCk9tfWuIyvtQ1gNFPtD57gSLPrA9d6sGQgNgo+gBVqt0DWIzP4zNY
Cb3yhkPF506WofpOhAt3VhDmdDJjlqCVZaW7HlQWgSIV1sxc57Uf5SzDXEwT
NJtCnNViZIgGDx21fjEcPghz0unFHncTQMes/EwEQibcQW0rnaLpOku+L3cV
lVTJLOjfPVOMa9uVQcL915zG0/qn6Xr2SBwzxaxZc5PkfQ+vBnrw2335QG8U
4FsqB79FhLqrDbYrswgxW1YyMqC3ouEjxULJJAF+5Ykzf+ueqVrRF6I04CA1
+77GP1wIhBQio3jtmtVmC1yb4uFeSaBLJN8bPXI4mifqjul2L/2kPSAiLLof
AcXKeypsbRndOjiXXBXiUz/MpSBQbXV0kSNX5JNuHD9gm9MS+TKdmZDIa6pE
uhjAPJ0D4VeRy2j0zYUw7WwXDp10B0AS6JIGVF4P44MVBALUUKW4J+uKewrK
URp//DUifNOBuaE1RTQ5mrd/hM7kCTV4myZ9DPIYXqDkOqfFcdwXnSfvcwB2
wbNvx5+8pAZ+Pc75J4CuPP5tlIjFvU9KOT+NCcbdhBZCoFJ6ODm09hgRaVZx
YrhsRGYvCg71sFOvhWPecmLsZyS4C6weJiN0zc/isiRJYphxaUpx/PIBu5N8
hQPX37bHT24jifMqF9LluQ26fNEBMkWxReW4A9hZWipLyaMI1LVP7u6FYkgx
S+O9OV1qcKdxZnZFnjn735/Dz/K2/9J4vDkaKygR+b/Ca2a9C301TavSB3JQ
2EZ8kS5ICny+qFQ0x4/CKsGnAnKkTkcU04Rmg9mxKweyJ9m/K4OjOviobf3m
r9SWpjsrVhvdfmh+YUkUxf5EeSesW2acAJBwiACB8flDvGrWts2/Ew/WT5p2
HU1D2/h1+/sXomv0r6usIMcIGmrNA7hXWTaNX8xwl3Hk579xEwInJLIIHfbr
XRRe3moyrze0A7+iLRGCj8Cfx0LX39wzOz4dI/mUDrAS6k8H/QMPqg/J264n
9owF8Z8VompnBkaXeqNixCbs++36bOtPmwbyJyNoOY3mpfj7hnECpGe2Bst2
z74rTcBRgvCqzO9DnwIQde2ItpfR6jvPMXKuIhLAJihypY6pcQoKuQNt0UOR
t2IWGtjgLWejPIlUaGfU2PHeoOkF7IcEJv/3Pr76ghluTzyz4+h5chAYQ1y4
5egjmSUdJkUuCMdEwIZERJEqWETIxb2x1FnnBDLDaZt3b6t0Fafb0b2HTWZ2
e7EPJG98lj6Bh/MszE/W2amNyFfp6ABC9/GDqRIhyBgWf4Qzd5LLqPOg9L65
aH0bGpz0n3wbHDtxCAHgSwW30zn7vOIs/3g4euLrzo0a8uIihTyZoX0vo9IQ
9hULVWd1QkJ4RxKMRWOGegAJkrG438uHc4uXkiTRu2sHpbepgOIydhMAkiat
I62UdhZhCuxGHlf1BLAD1CDogLqxpKbPVqmj7p4nvo6KqJLK0ldVKmlUAOmr
I414iVJSYiA1rQ0V0MDBpR7PPxF9gwrwIjbZkAVJsPFfp5BPoNBrVKXp2S96
Cdy+i3LvU0oHet3Yvft/X8OP3GtXYeAma6KrZfFEXR7h7YKCjGy2hfn6bTsY
Y0rcBbtEK4wZ22VIq7UMutzn78AxhrmSKOxkrHTbwar8V5yvTQjJGlFfqGnX
CAGA3+JJM88K5DZMi/+PfjgplYs37otbcV+38FbtizMF2AGRiWs3ui0JEfwY
HXjL73Ga0DniwxRTWlVl/HDxDABbqhFTSBGF7h16zc9rOR+QbmpIoEw0tu9k
j9Tc6n4QJHKC0wijp2pMxV/oGxjllEZhqTRlZx0aXzRD+lWrLUHJnA0F7/EL
wpERxiCjVr48Jd+pp5X8zLWVlftCF5IZWK/g03hYUSrcFSR9z5ngdShveIc3
4k+y0foGWGsr+UuX12LrtWflvgO3mYT6PlEvr9lM9/sQvsko4xw7iaUi/Tdz
KLXqY0RajOiGmneBK9GBdfSBDba3MIVrWUvBzrr09d9uhRtsWeCTEbc1IdDj
uQ3MsQcfIpd1Uq3lZp7wt8kcVwZxPOscKlHUosQp9jZMfQel/h1q2BggpTVV
iGIP6UljKrZvNNFCCAFK9LsWr+5bioCb4ifNqH5bGporVfS1qPHxi2YU7yvS
qc+A8ttkv7Y0nMKwec/i/OUObcdn0SC+t91KQdTU4Z4IT+OoUQm3u/YVPjBQ
mAmj2ZYhOL+YlflBnNr7c6VgIRSM2mZUkzrUYewPES3NG8kdN+/TtzCZTDrF
s/PSK70hDwIkS/WWpfXWks1zMSOw+deFLbAfGIdDVfquHTZ65JHQ9YMbtAS4
69yPBOcW0B1wDr4fYpVr334wNz5DLqRZvJGZn8OE0zaeDjHNQgEDrlCt8eBf
nqzB5oVtfCu2rR2WIDUR+3jjTN4kvSmGlY038bqHuKy3v+CUsAzGNg/KCMKr
sLnHHYlKBoHXmy88qVgVDzoUe+i2M+mO4F3O/NDt9z2g42fBHIjaZxmbVtDN
IfaD4TL8zXDyJJChf6sAAVzL342J0wEI03WaAAMhbTtvKi/ejfNDPaDLM1hZ
8vwzQgVl3pbWC87hKC33C6AQXeZOjt3P/Y9V0bhdEpvM4M0V2uLPyF1X3kys
FuPIeDntuurlVvHcKTGRQxg+BHQOwFgGUopd0oU7ZHJr67g0P8ZoCOTU0asf
QCLVoKDjCy2JI8JcfQWXunpmIrylW5hF3tW/0bXxJgYRiTkQl0+4jQO2ss85
Ztyrby/MaBaMY3kZcSKm4MkIi/Z7S3+b+TOzLHXfV5dWxHCcc9Q6oKe5QMgz
vaY0DFNszPqAmYjEvnAUf5/Rbs8YX0KmWPR65jpcMFgua746gsFCIicZKWwE
ofv/brLz0L3o6xaXLQBmXebYH0YLQTyTAjG6i70zX6WgFWG7cSzYMBhAw3KL
mOkCPTt3ygwBRoYpjcNi7AZXmn8rTtCoNptH/IgDghu39aU4Akg6FvRq68wO
23AAZiRnb7lO/gQMuXVcOwZpr2KudcNv9figYwcFl0n5TmCM0Xyc2AcXL9qL
0Sl/nnK4aO7Z64ZXzGTiH17PJnd1ChyC5D2Ga6X9p2DwCq69X9vYNUOOZ24b
UkEER+wX+1zKdB0JOGayt0HvEGoEJXwisfOZQouSMx60w9smsZ9qu0Qa3pVE
DxyrN0SMCJBs0RkL8ZolzNZuzohHS+qWgMRREDwLusEI99G4utStecs/wK01
bcnRo5P3XBoT3Hvtw6vT3+v11jZxYZ45C8/CLecGVrKk2tJ7NXYPVxePe1EF
rOHeCdoZH4sJ7NHC6TDlgAJ0gDS9wny54nEXUjuKI8CpnLSJ08XJk0IXEWjU
MzueUiqnU2IhrQxRs5SNpXPlrKxE9z17gNdDwFaYZOq+jTTKuexgV7qq7/5V
CtFC99AzXjA2vc/iR9LeqMRE/NzHS762jwAIR5SOjGwcXWDPppdmZ3FO6rd2
Z8mEd4MppBw9JTUFY5ML94xr6nAm1GhY74HSjO0+yQ5yH5wTAlmVWSFGY2k8
+3BQ7igXxtYUezeyhb9ueg1XvPfj75/l4b+yrz1Ix55/rL8dHZABEnc8CxIo
aPb0OARVjBm1MbjcVEMSJJ2rUV+D4cRqcnYNAbpv0xedK1KrrPh9Ve6CxOsW
k6oxPPOfyspJlkbQ7r1sJ+HZWISaGNAZQMZ2R/7rug7FWtYydPKtvpORZDMF
aAM050fYnftKlaJvty2HGkpr0IhgnVAUSm9mHSWwd5mFRiPSHblDTDoDVQKy
aDoAPtd3S7W4tEiSnVM0v2CLow+i0jX9xXqo0EbO/es2wsikgGA8r/A3dJpA
WoBY66SPHTVI76T6VefAooSt2gSlkXI3GgcnsrJoOSmsHg6lAqpXkrAhl8D7
9FJlENd2ziAN8vV7xp1mui9kqGCJSIB6FoOsUI1Gbe0NPVjl6JElWgJhbprm
9v8CJG8SgKjjyHsAckMB4Fq5k4a8fzEqsGA1/cxE4NaJX07Qmqpyc+BbT2el
2eW4fxKrYvvzwJuYMWv40ZPoYUSW5eOgGnoWqXgm31y6WEqjUIJbkOMM0WHr
SLTasg74cgJkYbepF1aTfQSRWcw/6RUl5jWjDXzWYL8XWGV9nXYlsMy7aIvz
V5EH9sppdVZNS1QFfq04+ZhSqJBAF9cXEBlLjo5Jvn+t9TpLwzRx80xdi2Vy
N7/RK4e9z8mQmh99aDNKRAAiL3NTZtHZzhNiYKD3NZ8wvzZJS0doNEkhGNWB
7EfEHyaz5hMIYgt2GZvJqTERZNmoGdhRSsYzCv6EQYO2YsfCgGmGIL2pgV6R
boaIcQXSiUThSvhuikU0qJKC/Q+SgHLh36UhbotJIi9JsIZ3pVDsRidRPxxI
0e/akZ5tN3/mLH8KumY9oL8i+KkCgkAjfGteuk2htlKbSCl4Sy11rE2GAxuT
vOrsYEEkPId5Fzhx5AIB7cB6GBwIXc7J8pBmuK0m9ukkQbcjCHKCVGpn3CRZ
eMbMYCNvqN2OI0qIw4r9fV4/tDSv1C1TGUEWOIWMZxk6hYQqqYwsEREU7mHD
X6Ccd1eo1490P1Gbuyg33U9JBZ750hYve2hwYYt4kIzGIaylPCs4qXJOdLaO
VFopNdKRspw6GGB8sbZJUtq0SfJJoHWH0zBhbPMwPS9Zp5Fx4RfH0cDbcNUk
XmiO0JbpoPVgf/Umlb/0VtM/oCeHf9TtLbTrIcfG79IsrZAkl7SnUcHlIWif
kBaTBBhrEkz2ZxGMizjt8YYAh5zWNmnJcbIN/Tg05zGwSzn6xgIhCMhXBSqs
+bYIq8IOHyv+YEOitHeedvx1ueYTtP9HWwxgg9RVl3F9M6io6exMTFi39qnw
MEpBqQTpXvZj9bn1qGQ1O+Ykxjc0QaDJEQUowZ9PTjH9T64NfBUf+dG8YfkG
lDnWhf6RBbx0CO2K7gsdP10J3R0WKSeedO6bQGl/hh1TRJ4CvFdJdelJ9Uk+
tKqkikhFkSnyhIJWBbF1vtpXH7U5XiWyTKkqeSHSFg84aaq+iqBk3ZG4RffP
AfswrLXfatEUVoFTkKzO5ocQt85gtvIVJRfFaQVwrQHwuAxvGCFBTM9bZNXj
HtzqmHky2bZg5UnIKhu6vkZFC9Yy81+v7vmR+M2vz502qx+tAGFRiI6/Q4d1
o0bqgn5J6l17U93nON751lOnhyxHWEZujT9VvLaTGMmtViOjGFcZLhtZ2Nja
18z26tm88P8tQXZFnG+yuBi0jHOlVVxOpCt8Vl79mXTaZ3V58TlRkHG6q8r6
Moh5ZDMkE+vCujqeCBz3+iSbMOuCD1Ite8kHmCoah/HlFQVqqknAOR0Ia7nK
4IpfoQLlW11Qrwm1QSGr3zpCg5gz52Ouf4D84vOpn79BH6HCXn2DHwC0MQB2
q34BizsJoG5AaPnp+yIcyP8dW+HqxNotfb1LwuXZvVZvQBcS3R20WIE3WZ4k
Dy1oN6uOpvnsMOdVpQy1k0YCdrAb+P0/uNpLP4zijAjJtB7bs5tn+UUWX0r5
WJB+LwBEKnwjJyTWMuyPeOQ4dEWDwDz8zug1dITxiQ/9YU+0TFD3AtHFwhTb
TTLlrxQQ7d0Vzsqs8BGdSd6VQl2HQDOKpdeZ/0BcWnPc9WFO8GuHBTFF5JdZ
o2IwwuS7aLVrh58pmYN/7+8F0PgaYF5j1xirTGwxbbHfnnFkcbpmLB0P8sJC
Pc1taz/KAiqayIsvv+i/pmMIrofxlq+EbhrFKz30qPtwaJ9cbR+Sm3DhsPFE
IcYFtM4wmD2n95Wvthhpv0xbSSh5mLaIF/M6Dh8OlcUulz1VuTg/XhxoTKVE
XbjSPg1+4OeDw+b4aiD7PZA0GrNNxdbZw1YcinsFdx39lu8N/B+5/YQe4i5d
GJWSsQ5h+roEMCCzhFB1MLASMIOuqWo6w7ng6wLJ12zHjQCOyZgsq1chMqdT
KMM0VDHNO25sxSA9Ouwe0seudlzsAyzGLcDY0LJUzEhr4cFPSynRelkE0Gs3
Pw40SB4qHkpOcFC1z8t+AOytwnJBtfVfuKlaiZlwNZoM0dulcIHxOSGYRkRW
2GxUgjA2a+aI6V4EF+0as8b2xXJB1wYBonu40HE3VktI1dELhfpnbzJeMH8k
Of+R7x6Q0SjDbDHHukhaBXmBbQvwF6gRjTvNk1dz9G4gK3Xcwu1vr+A+7DBm
uru0hJ0bVcZ3lRbMfv/hrnF3hLghyU1H7jI24ZYZSxILvGyy06+xzD/4zAI/
XEVJeYoUfcn8rCASMzJCm5BQZeGCIS2oQKAKGGOK+nFDJnmfdCqz4epBl8+W
UyFyrhWhss38B+yOq+qsuD7hWPijklkal53G5smZu9lFfYH+Ukl5QNlvL2VX
qJTzYctL1R7y7TU7PStXs0nibDPCtG4POe7DghMWklRGpWXC4+xzLLRikqvu
CShXauymefHDWtkva423fw39AsrSK2j/y9LKYmc2y0RbpQXY93/5WNUVNx3h
VQ6yPAO7TCqcu3q5AgZehp3IkRIjdeMB581XbiAHeHZ4ozAEWy+KQtrKVJt+
HnbWQd1jXZQOOp+XlrLo+rP49cyAfWRjzsXIwDYV6WgDDu8dPgv7WZtJQIiN
qqbLtZ1IHHWBCyLj4TP+InePXYR2/JseDOh74SrCF3tC8O+K4PC+jXVgejqr
XvP7w/qztD8O0PayJu7X1fxjRZSig6DhKqpItHuekM76XbjqPm5nOyhW8av1
iOG44yaQ3IM1Mrpb9wZqeqZ/xpwyfrnGQlk2Z9nMRBkD1+ZBq/6+mv3ck+UC
W9VvmvnKEOniuTYRoPrnTmsnsVPned8WUYiJM6beICcKUl9gL412ivCh0TjU
NY0N32j6ofbMbzJGCWLSa7wO/axv8+2E3S9leeAJE27zLhf4nUtTyyMuJjVq
g6BvxMrIVdBdyQFZBv1TVBxdwEEsmihO0SAsGqOVZ+Nkf11coO+bOIUZYyNo
yu9c9nch+goNBJ1TbCfxjDsF07lGxnaC05XdOBwoFC5Pmf+QNhWaj9kitCZZ
wbn4fbEr0cE/tfd13EH1gueYK5Y4QWTjog8c9CepTpJuBP3WGiRsufojXGm/
5Skmubl2iEgGWSxylQkLvP1zdDFuvcMwsxBujspDjMSwGZHn8/9pwJJy5nTV
Yw5ZZVcpam7TU5lHWvb2s6Is/V8+2mKQO6gdpQ3agu4J3tUIMcQZk5Ti1iU2
r2S3IF0bqHQuoi31WHCmuxaT8yGiguxFPMuyP0eqi8y7D3OIGhvB3Taq2fte
Sn459vN8Z1HKZ25plHt2aRnuhi5l14DeH5bnz/CeVw/WnQP/p35zm/iFhvPe
kuNZMbnMTnuOvHSUPtOKxSOIor23TrKqvXmo2pC7tbbtoDw/+6voPNKy+842
YFeIB/Jh4RmWoG0CW0XV5vhsKAbEC/7l2WyvICRVCfN9fRHN8FnaYQ//B3Gv
lcLQ1/vhCPUUo+PqpTxSxNSegM2ZOmOWjm1omy60UHnuTRwPhM5FrmOe3Ycv
qrLZsb6zVo7LTWtOnYlMzgwCIbuLrIB+IkxHtSZspQ+Y3+pCZHZkKVohUfuC
v3ZGUa7YFGH8hMJNMpiuHIh9psIbB8f9HUPZAgDdQLNR0tP6beUGlU2LdoOq
2ymBp9wM7DzGvUSjtwakYZixcLdvKo+fNg46Zq/nMkp+Gv0i0sNTQ/4e6huL
AmZygAMK4irf2tpxo3A3oc8cckzUZi0VNBEeg6zPTx+61RcRD6MjpUB4p3FV
siVcy++rmblSE2vOOprZ+o7YjMSqK4k3k1gmmsB/24qeVlcmaZ5JeXa0RgQp
S/JA5UzuQ5/nbNkqF2D5HjpTKdV0WVTR0V/sLmSc19sDmhe4dbXibUI6Wf+A
sX0Naza2fMsLiJgZ5g3/iQ45JTXvGssMVzpNrlXlLacM1gpzp6NRXTJMYDBw
qzcZUCUWZVmHaaurQ3GcE74hBvEgE3Aq6xEw1eE3D1zjmQSvZsWOz70IrXm/
7dyOWBt+Jpw8zF/bUW5q5w3GR2eFJPky/XKwqsZN9fIBlD8Y6FhVIcF2tn7R
X2n53f0+IfisMYX2DTGW/1GPk5Ui/sTrhKdTIrM48WrCW0JASbMO7OUEc6NM
x+mHNYvrUIqDXFOzM5z13TT2GRQpTvHHePrLp4PVnqot760XpgfmBhXz5bxr
W8NBtYdtGY1GO10gZyeL1x+yw+PaTL+bLP1ewDj1p7ipCMmQi27sr8HFQT3V
/1hzZg7u30wlRYx3Xpd3rKCOuMcHGGsBfe6NvNrfDPvTZpL6zwAUcOC8sQKa
pDKp0aYDb9D1E9FaaGLzD6YTrKbaOlMlZzDXm2idiLu6JwHh7yNDLDoUnkwa
+DQZD2XLS3P/NopDl2jwNHBGDM3flDurletJW/0DIXvg8bqrQV4DE/HBFuvg
kslvQ5RXOnVqfANkg00TH+enIy/QiHHj+UBe3khyvrNerJNjYujPghflb/ly
VRSc3otC+2njZN+ct1Sx1CGUTXuzfcY/9TPI6MtnwarDc1W2uqdgw52HXwwT
9It4Udnp95hBKXri6H4a96a0iDzpTqdItW+mpH33C8dnHyDo4LrXn7b48/ZY
9m0DogkjyAuk+P8ORwxHlgrxjx8DV7bkC9An/GULVjiOA9rHiH9I/sLlCNJ1
Epgxs31iqR0OWUuEeP7hSJzZXxT1hwsQlc5dsmd17FOUroYz35404Sw8Mh5O
eLiNKqooKI3/i4VvJNt7F8YnDZHE1PbaePF24Yv61+yl5tZuiOj2z3ptZpPy
pj54Jx7oNBk9sP/aRzGKkKbknvPXkPYk3jGbc/QtUUWCikvCEyJU2eSjEPOd
Iie+qpWdr405o5U3fYz4+9wuPeFYWam2KOX3dG5WGhGrBCLTzlBTSIHuq9lu
P0K3Q0L+QWs6sqDb+62L9tWjcayvhHJfRXtwxpX5SmkU6qnWJnMQbMNFqUKt
hZy/Z+c5xJwzXc4iu/1DlHHSkZm9AlhReENyY/yKskRIfr15SHdUps+J4k4J
XvdHTBFYda1MKndLCwjU/bRKIUJiGqo4Ihob3KTAb952zl4TXUEcuLWFdhQ1
J4ywMmXCDhd7w8lEfUu6BqzpVTUGUkkAslEGaaxYx7ElgoGJPeQUrVjZnC5/
BR96r0AQepFcliudpJ3AlYbwTt69Sp/7mm1DSbyl5qxYG7/mvtTcZ+hqjiDe
d7H9lICPRnDu7fH8edNtmp6X0J4wyvEHW5cO1mQ/NdwMDJg5o0ISAoaqlkuX
eFxLMsLzbe91yemffAYJ9dPH3/nni4weFQCIshATA80YY+LyYyNJoUrly6Ty
29IZJLPvEWJcguphELjS8n26QV77ymb524boYdGcGMVUhqP/wkm/IKSr4ZFj
/ztqO9tjtFxyA7qP1TYJIKNbvFWO7Q3yGNU6y5GD3ulvv3J5Y8tttQovizeQ
QS33AMTqJCqEZgqCzX1Eg4rL6P8URUSCyq4WztuRUaRfniV2+g4cPf1nS7Ng
mVamKcNwMq8s4hzz5o1d4DF/953AfGXoQCP07CTWCLcdhv/QnC7ts66w6EKe
HqELd8iE1vWeOg3A/sq6C3pUUas8LB+zAvNnHdBcZY+OODbzvaV1cRpg+HSw
maGur31ZC6D9uVzCQIDxmF03uQ9VTWrUVpDq+JV78B92LGO+4VgJH2SCq3ih
uVgW4PXTEYpQ77cYseynCaTwCpQtA8DnQEPs3No6In1tP0LVBNti4+KOdWjW
ohbX8xU5Du/40nQcZUQaOu7Q24etbLhk8riAEZgUsK4ASAf63zDX0P0pA+Mf
OvUtnv2mSMu6t9A+3gJF5AzHt/ytFhxRebnuuJUF9a2BaI9Z61qILFOAFyLT
aFmkziZ42EXw2T9kkGfTSRZLrluGaLhMtZgyen+RC++9kZvKsggrMpydXOMK
9Vv6ZaxSX7inRrqB0a234Yx15uuG86BbYlQrED+rptzf1Obwm3H4NPY9BY/q
+Th2Q49fHvzlqUwRi52hZwaaAIhgKw74g8gAk9aZ1VrtQGgq1avmMWNt+ubz
765+xpqCGMQmRuoo+/r+kWFSON/ZQXfYPwFCdEW2F4bDFUjVUzWlF5TQvTI+
m9fyW0WS8hu/tIoMAi3aYncx1eaflTnAEKEGM5r23xXEwWVNU1hpaiWexqqA
kQhEXrfAxFVTvSp7PDIeviWz3lWCSumHjAKO7DbfLhF9pFi8DqTlUxdmXbSh
Y3sbaf4suoZggbMGytSv2Py/sDpZwZn1UPyVIj2rybRf5vb498n7poNiGV/M
ByHAJbWRwSINC35kuVi2Moh0XY/WemMA4ELDazr1CJoqM9Yu6XcUAVpdjJC6
mZ1r2sr12uukcfvcc+PG1QtX8OEykfIutamZdMPjtyu8gL8+txAnHOum7QBK
kcvWAnXfxmi51qsMW48H59cd4HgXylRSX1cpW+EVSDEDeMo6rCBQF4Vl6rVx
iIGPEGq/TEzez5XHcdaZ5zBTdS+UkV8vRYtsaqri45VaU6V7CEUrQIzj8ZM5
bEgB2SH3ZcyDx/YPhZmxLWkyvI+//+jH016ztbzlkBEApWcaILQpkWIZTTRL
zmEhJKSuFn2RAYPcAzqp/7nYYqgj8ljG+J1TIg8T3Yqgc0z3JNl3DnA3dQ0s
2o/AzjAmsgsApHSHbcVSkHB3g0qR1Fucjo7+RmSqAPkcQRIYndWCi61RKOxZ
sp8odVdIIwdCqr9jaZOm7cyCPD/8ePhCnImm/ZePIdnwfF9Tiynwc5cjHLqg
rinMgBk//crn6i8GB78kQvmfV8tyOm10NyU07jetC4e3VYC24TAi032tA7sT
+KLMxXF1MhbKhHnPK2CPu9wr5ZwUJFXpuO0M5Nej9vniBj8ZGY9G2LXHjLAF
oHpj0sxuDUV9bHpSVPVvoNS80VZIGqLHlThkktOE/pE3p0KpBILmUFVN0jeU
ZBUagEYjDwMII9FK4wdUDcJNV1HdhbXEVRPobcOpteg6AuoC1PFZNfdarico
uKSzne0ojtPML7JGftzTyKD7XaNoD+goVFw4wGVLujR7/L09leiFDExakyV9
SdPTNWKx4+qefb+rg2RpnzNkMy5y9npLDi1LNlIlbxa4ZF86Glq+v7Y0kWsD
AY7iY9nFl+GrRb6K0pOD1ZJ+r2ADUHcXhbvaoyDTCf14OsQXVuvRkH9SXgD9
MrxyqM3dmCoTUyVuLeIlBQtEbF65PRstgs1DCDknPEVNtTPp1nceaYZ3oSCs
S8d7BRt9UkJGxWfAVAVuJ1gHnDYq9uIVqjNDx516AlDK+Q2mQsJJ1i/A59bL
z6viSesm0tqEo3fQArpfZfloFiFto58CDiEuf5pQ187LL9UI6bhrHejEKF+u
6EDdV8o4NsjmZ8yUuA1439p1uhXdPUOD3v/mDdlEFZ9ov1tMKps+GMWBvp6X
6ykFffdQNPPaa1YTgIlhUbXetCLQLHDKBtG5cpJ4rx0OY3ERSky9ZrR9DkH2
hXQAo5+eJn7ScGhXcfsjltJWqS99lacYqY4J+koLzYbZasBRecP6Rs+Q60Ao
ZZ2EKsH+KzpJhbvvkGcIrcYBvlDawTY98zh5xTLQY1iV18QlV5gY1dKHrDVb
dPQ0nEaIBwXgoOX4Y7KsRn5UyP/6MmD3RPHeb1KJylnyHn8/C/Qqqf+aUl8/
ohMDhoo+Se2qkBOuz1nHbvxA+/ESOcMi2G5NXhl/s+P2i+4t7wOLqcFk3MTO
1fbAgWPMKTdRhX0VSgZXDcDODCO5O3BL8UNXiseOcoaFMt+VLJ5+NokemLdC
jUnOxX0SpjaPYsZyD0pqzGOsG+eql0hGQz6edpbE+VSV5HoKW3u0ioIihOe8
0ZVAb84vvhdh/AIfbe9zHl1k/68S/72KCrmG14ITd+8tACQt8mXCrgQZhP/P
TNvvYhr7fF2ayAFpM/yWRux5w3jC5P5i4mUMip9KqFrWbZeCOWsC9IMYRcwx
qHdprwa4Ef3LtmREuBa9Cg3hvxYKUS1Y2NgGA6jbeh5grOq18lJnD9cUCqyB
1+3uSrevY/XP9Rii51FG+0SL1bScPJN72/YBkU1NwJWLuysWmX0zAMd3bGDi
+pc5CU0VrceEobWOzSxVIB73eUxkOTeXdN5hqrx1t0bpnnrtEeeiGrSnzApx
I7PiwE9VQln3HC0q8Vai1lDlIAphbUYU6TyuotFb4vhpnutXgjkdnc8WrkQf
c/CuOgM49fJBM8lGJeUXm2mYyczEXi/VPn/LBh8E3XQz58oLzzb5EDJ4Bxdp
FFy+LDcIbGg55vHVH9U98luC5ZhQSSJb6N7i/k7mzhJtYK0+S7Crmu7gcFuX
aYLqWn1qhhNY+lwVnnpu8cqqwAcK+G//iUKg4MvMpScMACvPT8CVPSCvflZp
b6pTImxxEZGeLMpE2PKrud8IGBqGS1XowG4r7/WpbPNjs7lG3ZQlq+kTJiPz
HUpGRyfIykz5g4y5gRrm6/5yKeelXYx4BH6cdfLsl/K0y59zqL5liIiKaWeD
gEN59cGksY4OUGTwKUkiL92cBxQ+uzo826B4GPVkwHWNT7Xwnlha506xF939
ndTmjAfWV4caRgV4C5RomGOEltQsK28jfudt91Q4BeHGn7bqDXmkBUxuucnx
ucyl4Ew4LHn1RMpG4dX5981/PRUmLeZggwQpZeQV+P2wTQEY6r9uk9bcwghl
BqTa0d65ukbgpvn6rvcD1aW5wcd1A8ft46uj/icH8BoMpcku7bF2nDUQNSlN
cnpLzty3QdpojjktUNVXaXWq4zuyReM6EKuPDna51oGnkplW1YjeCqKBk5Lt
GIkLel5jitrrT2CNPqN2MiHJnJ/kN1fEnL2PaUl5E5vK85vimR7m+Tg+AJBJ
heCLXr5HBXj2XBOjyLNmitjOq5q4CA55yVO6U5fL/ZWGUg20OKXr10v/bi7/
Tmt1j9WYleV7QF/yqV9Tsw/xfAERyywIPv6VjKMlibt0bY1eiOaYVtQmBtTH
PTDiagmyM+lNZq+MOwAdd8FZgoUrCH5OveljFQDT7FleERBDJ5V5+913SC3d
MA/q85cIzNi6mi7j/VDJPkYXrSR1udNpYL0zVnYheaDzitEqTtsCBptZzYP1
QQxvwzzjG/aPCEDzOn3fK0Fs+K/LqQD9sitABkwGug8lHGPVFr7VIC2z7r6N
0XuBzDes2COBkbvIOHBgQGOXwFAc0kTvQbW9EiyPOD7UPyXRjFd077J59Vna
vqb8d9bENCvi2D1PNmeHOfAbt/WWJcNciOVq486Ej7h10fZZJwFp1/nygGSC
MkKZqWlz+uYa91mTrSGu2RPOJXIEs1OUJjiOTsHSpBVNmidpwKuLq50Eyk7v
/+XixQ/KyvPicdEo3x5yNeylJbKMiZgNJZjQbFBZju77USTS0CRIgWljduCj
Zt1lmuoP/Rtprz/3UHbzotdb8xISXV8xPPfcJq3zxbgzdWpmtXBR7ffIBGFk
o6ISYUpQQkw0pJYVUYgzPE5SHdNlT8M5q2+cD9lbt1/xi+8dSdhhDH/jjICp
2UNsnj3I43xooxmoQjOEdntfQe8mGe1CtdU0HShXW8Ygcb2ytfkrkXRFsbpa
el6pYK243qVRt7Nj06c5+1mAgoJTbTJTRDjTJ4AKwo88j/3w935GXt4urF9o
YpRAcHvttXE/mAo2A4Fg90o3/hriA6PQ6kGDMdLbKc2Rz2lQ+/7waDEwiOWL
u7cnkfxq+oV+4EBxmgd9PseWlOSKU41oYfGyD++ey3SWgD9SJSaSWbrZHD14
aQPg0DkTLPoNt7/FAe6fCy/fCqUbF4DY+rnii7py1ICRVp+mPqo7RdjBhQ5B
UM/WRgD+1bfcFA+OnXl6PakvIgrTLO7DkxMyZIK/iPtmXMWv9O9Kl0iRHllO
0wbQo7KOw5iGbAG1kdbgJ/F5mWRqAvdNqhZoO6tDVrhqTWzIlC/qOnBagCns
0Ef5s6u2IjpDxP1PeSffel9wx+5scFT8RVohVIA+cXwTp5XPUPWbrOkeS61/
h+9sKLVvwbRf7UviZ6i3ibh5dOL91pBJGHS58Ok3rlfx9fUp882VpurZfLDR
MK7e6LFXlj7s9XpLZcG1/c5N4ODP9nngMCnQBgiXDwFBOYR6v0JOiu+b+0cB
V/fQleuTxvr2lQIAJI7hZveLKibremHbOjWl55g6dba8pFAEBzoTAVu8iA3Z
+U4Y4FPVBjKKM8zCiEKOINgho75MbhrJdhUOj/OKKSlr5V8N6yEAXXXoKQdm
tTptJkkx/YVr9uZygA8jOJAsMwAgcl3U9NEvQ7dZbRcwLbLquVcqw/HzYtEQ
Gv5lbUICfYXPaTnbNG3UJbsDTSEsqe2zCJoFvbNm6Qixx64o5WgoKkwZo5a4
R1XKJm0dzwLsA4y4+O35LuiNbZ3k8zxXLvJwU2/3lG3gjtcqSnS6qwOJzoJP
vnvT5FNeXjCt1sh11o88d4GUIeFuFddY1VNn8SPukhuwwqLRH7M0GWt5MWf8
MtO+3zriQmAOsx0185mm0LN0ULNDdwX0hXYHas9FkgZjO5wLWSEOSjcmD6GL
Ke2aLnCxtUjIBTAzFNEb8d1NMmbxVYIh7FRt1WOqtyhtd+NDwjwtRrN83Iw6
PL+CqPFHyROfq2KVCq29Z4QyG23jx7s6m2bz6kBXcykAgVzVvJDhCNEzx5+g
HdQL4UAykGS4bZAb/lpQ+DtMztOp6BTHYbo6ewbaKoe27cRzpYp5OJRCkve4
upZS0HKp93jMtzrrtLILWYTz9fJRoE8j+rk6+yotTl2aR2qWIyqyLaYAQmkf
NlRGt9zmHCpCLhYF+or1N8Br/5jRO97Ib2uUWFXH5ijxdMB3sKSW6AMyZkjE
e/0X5NIBqcKiOKBEighzCxOBOIP3vIwaPd1DJmyWj9HA6H3eJA6z4RjIZnE6
rTKDiSGZqcvUWfUqSJfZO/jVVWSJrSe2NqhEf37UW1Yu1aZ0IUugj3lTunrY
GsP51tyETdhrM/Dqmi4CNCVphcNg5AIrLu82317JobNe5VNVWjBd6a+Ui3xB
y9cbM/SPRfFb2K5j5txQbWYZT/MQByb+s9FBd3AEzGA3YIVQ4jWJnkarrmin
iWtj8tI9Eof9qBCwi+mxf/Yu5r49WUPDhB9L6j47eKlMXdrj/6TPTM/g38it
hX93YGAwxV7GIBlAt25wU0ISOcVAH+o3poNpOVrS8J8C6og/z4nTAcjH/TwA
ACzqgwAysEkuLFYYiJGtxRmwtgCBNWAR46EXLS7Q8q6s1khLNims+rKupqtY
3G1oBTKz6f7EXekPfE/hm14gpcc3L/4CSTdNXQ+qRPFAAUFKCuxQDVL5QB/j
8LV8B2TOgKmY4SmMdH1qNTNx5ESTTpa9PFujrQ4cYi6gqYUbtPVHf/wWeuLP
VZSymbn+t94zeWhIYzWDn4uR3A5/F7VnF5/aS1/cdDHn9KOXxh0zl/gA2WXr
eG5ty90/t7iU9xn+VIvQde3euAMgUr6UCy/X8pOOT2OCQ47D31Pk/eZpVxIo
l1wnYN+REG7YTmT94tce6l7CmTEHLswozYXcx6sYMcxsI6lbsNXMikvw2jSX
vPJf3NfLZB6x+SMeQEU3YJAE4+urAKDmG++OgVAqDQym159F2AfUaK7ETJvg
8PlMek79xUm34muQRIToLaAxZgZ0qeuHA4bCTyLr+dTfZknj87z4kFuWRgeH
7apxWe6rzESr/5nDgEH71PwJzOdl/3Lgx6M6UuK5GySxe5Fy884eT9Ufo1tD
jrKgctfaSfW0urEHd3m//W0/gcuf0gFINCUgs/mHcItw7xLgOe1g4wZ/3E//
Skw24CGAUAXoPb+UcU51y6LqjwWmofMhfKktrAT/QECLjfLaRgZBlflLKDbT
t20HYXzlzEtG21ybFam0oVxrXDRIsFUD6QBv8R0BqSazIwBquwsJWRh5zEXp
ki/KwUTjShLxISHup/fW+oRavWoZnVlsL/cdhaPGWnYFUL7w38Q2pbe0KJqp
C3SfWaB9czlfJdgQQFNDD6vM16PuElcboxcY9XZthvBlGDAlTTiQ1ljmY46F
J6UsQpLHAgMuJCIGAbQLPOafqVDwVNyOL/QaH96/RTH+hC/lvr9sJbngzn7k
Nk+Oe7R0NoAcn4ell+sBttSzYP/RDbx3LAPbWftMaaqBy2sOKKJ+qB+8DW7+
pYe0qk3XZ/rc0uBY2x3hBvIeZIustEf9DFlZiYZ3dQGwdj81bteEk9sG2o6K
ywIOUazJufW1w314pIEf7niKKm2/+lLdlg4BYVPCOqL79JtLxWnLu7YHI4M1
9MWzmQ29+Sw1psNr9PKrihPckZzdetaT8jA5SbNMxpl+LGWYV9u874n/jYbu
G4tSeqyAbJtxQr1v3UYl2biYDTae/1k6yNxhPEanwVw4VYWQcey7SwL2CfcE
FpIk5m22Xv6wqsjkNaEtcpfxRFq51U0iGf3XDCCqbPEmYArAGo19uLQWMkxj
6wXKk0Y3Lmw+Co8pm5+mhXgvWOThjB2n8yIOuTiwzvHsO+MRS10NfbzLcXXO
DU6t66vAWDzx4wOZ22jtz5ivPcLHUXo9LVsQAhDNuwYY/xRe/gkzR5onff38
L/7S6xsz8asrRvqTN3wTlH58vs5qkrZdnanUO5ezMDP5valpbKFq4Jtrwxky
rSbNYuX8gY0ThRjnmmlpdWexL+O9L958BuUMR+FmmuE8fNMOYgNtmq7gGeZV
E5/sUGK42zQTZF+yS81hzgddGfCf2L5s+kyVVDPXKgK9xe9mPJ7kQuZyDFFE
OddZlUEjD0JvX6faPdnL5uKwLy19IGRFap2kffSQQGeEjNc5tsU8kYepA31p
Yh7BJmvs8Ctg86u8bFXOZYGv9QFKvy/1Ro2oHcK2TOzEaCv3N6JXrlJCxuLL
I23pTzB2PMxkIztMxopzhy5UhWlLvZA6iHuBvBFvIKDg76JovOc2T1ezEvse
v1I6qXrt6g3eUWS4j6TnfSsFIQxp/wIKJAfGoCaAOr5pqQ9l2HVXrHrc07md
39ZfkadpJH5TLzHYrDrt9Rhx0ElICwD4X/9e/O/eu8+jMKTdfXMAyeKs5+mD
9h0GteXAl4B2yHVq5rjfORtHPFFGWZtwISd71QuounHw3f/WzTqQMBuN2lh3
1j5sehQHKG6Alnzv1RXIQ5dmJjg9Vf88ekouMT4uvPvzy/rKKUFxzvA7SoXN
vzrdQVBSBBVIFhOobkhFjChAVIONovedVbDEsKrTaQUaRROUQal6gwdEZFK5
0YylrnGuq0uyDCfEkXEs59lbazna5sJ5QOYDLympRNJ82u+DnTtjuGcg2zoP
R7wPZzI0gfn3gwLU0NwazeqjK/143eR7/y9JvOtCPOqmOyQV5XbnwhVAgt+o
XjUZ0aR7skjTGNC9RUMsDsW/V+HHwzpRcz/k77KHF9DAOdPT1Ry+H2LluH8T
TnP/oVz+Boc1tgceZ9dl04L8uNAj9xmCHJn67y1eRJiWnHMLN7w0cBNjJHgz
9OPthobBwgoASnWd8MQ1KVgKZJwwNpvjUnjmze1C0CCk3zXCrJO38YCNrA9X
S3nqXPWOXH1/vY/cE3bS96FOzgbQ4vdr6z84Z48/VVf+x0oLAac639uva7IC
8Kqmpatfkx+htrtV1gHJgL0uOVzfs0Aqk/ISDus21EW6Esook5Bk9D2zNduX
jAKD2w0oE/a3PdqN/AwM44K4ShjXx7dWAzWMrRtZ3lib95X/iMAHoZ9MfslU
LfnoPU27DJCS9aJRmRWmsDylZho/oym3Xy2orCiHqU7/Xl6bsAmaDVYnmDrv
Iwy+sk8DE3D4RNo5OK+QM+UbinVJEQp48UTGUXKxQlt6uhuoSE97k9492w2f
X9f/E8j22KnjObWfwhBIhmQFLoJ22WBdKLLvG9A8q1ZNG7q2uobavM1TBtQZ
+/K719v7XwGs7+JXXNe9kZDOChWMPhbg8pUtwTMgQsjGv2kS8gTYtwycZeR1
oOx1hr7mEoG6XpNVOOIoXsHtq0Ks3OlxahI1BVXFXALkn+DfZ0U6Sj0E4jHQ
L85W6OwwdbkdOy//MJjEFl9bDbPC0uFwW7zW19/xHINC+xGGZBGiprgaY1Yu
Eonkg+fLYTFcO8NnkAJhXb7UfNTyg5OnO/0lKgFGqyfS/O48rIzduLfsPlfi
AXAozo5OqpmnW2XOtoyKBmq5I3kmen/yJjqhbQ4vbftg01nLZ1svy1sLw0n9
LldpG3HdzR68C/EbojKnzmx6X2REtnUAu3nPJX/d5FF9fxZ1uZYELrs3GeGD
le7RUGV8zPEsfpM6EBRDmQVPaGAYvXaDz95qwXREHKjDJClsdStqnisUmVPu
nN3gT7p1G3xV20two16/Dv4Djweupy4TL4ak+V13IDuY/Z41xxTOdRGH7ukp
c3oec0FV98Q1bWMTC6ftQS4hCP4hy8BtgR3jjyqfTTi5BNc0LkcY6iB9sqP8
KlbwKiz91jIsDZ7n7CMh+LRMAiiIImr2bRHc05h/VSVCWIDbbgjLx9/00WHk
ZJhMvFGcdaue8gieBeEM95HfxtgwhXH8U9W73uBTgDy3PHnI4wTizwEn9kYj
l+7GDaacnPYdATByztICyS9jzTTRqbKWwsPEWZBU/okXzJnk+3A8GsnqVcue
ZvCULwNuKI8cqbWwlvLHR8AszYIPLN+mmih8WH4bpr933u3rBEg391VttRZi
haper4Uv4IFKNvUiPZShhRIw39M7eC+5jGFYLp2De/kgYH4DawJWmU5o43Sk
s/tcVFyCMvtHqEVTMlK/GbblxYLEsJQ5xnB3doLWJTp0GClJaHAKj+TSBQGo
CjmYonWN9AP2xl5Q6IDqFTHHDEhxmHD0iNJ2W7qcfr9LLMaNHi2wbeKrRgyU
zJ3dmZzs/rqd9QlaB2S4Qx0E8n3b0jNWLlYJte/LPwiortfL2OMF/JaK8Vry
SR/bAzOzARHzhVJxpI2Eg6QgJTwQJaGZySlLhTh74O2CHs5gRdEe1zPx8Suf
ziEwBQeIHh85mZmbvb27Q2KoL0EkbCsQ+TGOcB2wdkImnBMOrlhdH4Q7tFIQ
dpH6d1pp7LSshpT70xdOJbG6ASHkUdh2JJ5Fg8NN306FSQ4yBIEueJVfPGXc
U5I78Xa3idLTgWp7mJe8rDCG1C4fLpvTpDvLMF82umtc0OPIh3sJxQMDDc1M
MAh9JNnZsWywIKIg8lrimxhOfN2NOpZ5vxNtrFNnJmrogc4OLZn8DfUlfvDf
Ve+ZkTEYhFjTCSr0r8L4/00ryVw6ZKmsD8rrrjSTaElkN/SZcx3x/jm/JXhv
b1/7+elK4CMXSVzEQ3WUN6fp27HLw8Wj+NYg+VF6FD9nUjkbGV3X2qYkKD0L
rvr47onfVYgUFqjVAVQY6oNb1GG2uvx9Lx+MJGYm8N1ZiSW4TtWph5NfmiBW
gdCDL1G9DqJwxMwIjTez7N95uN4F8jNQdGVI5Xq1q7m0gEBQx8XXUtTruHLU
1fxtzgldb1KihyOrzS58rLH0y1PyRxENSVCUBB82+wKD/jOh2DCdlBbSIjGy
gFLfQNW0xr7S3cqWetQWmoB1oLzoPsFP5P248XAFD5mEE3Ojg+mD0gp7jn5r
jvM+jO3EBaY6DPM6Ln4H0ODyyJSTU9U6tfReRqJhwuNLBrFBsK8/tjgbqw4N
YtICx9nQ2gtv4OppHWdZF1KJZeIt1StBkYm1ooU9gIjB/9kDyIDDX3/813Xr
RO+aAStWK0UAIVxSLgX1ltMasr1lWX/do3YJ/+3M4dup7y5jsorNS9Jnew9E
gHGEYkosfiVRKnXcq/iWYWIy/stmay9uQQQruAB3EdfYTp9nHWOp9tOR7MSI
maJ5Xu3P9+iumY6kiixW4FQR7zGX/KGBUUkxOVi6wIXfuBrnuzLdTgFY72Au
Z4tIsN3hNG9fnSXago+5GCIdE//eUVf8l4RwC5OvK7Var1bCD8p+mQTzZ9AC
Io6i5E8RZCKVEDG1L8Iqzd8nUY1v9S7lS6UUnGExSa8HMJuR9HNOSEyecj1l
9VxCOHCJijxJ9q6aQCWvid7+UclUdGhJiLFC6abt+yktw0In+PbbdjxtpR9r
7YlcbV87n8xaYe9kGvmeJCi5C0WcWkxB9NqpXPg60f0rz8AAgeKiyax1E0io
X2mfq6HQU9E+LN0tNJZpZke41t0sfO7XfwMZcQpkXeZ5bqetV4aPCBQfEdxK
1i1p8xNFeQAA/fqgsulp7CmP1o6WqWdqsLJXP2huJBJDmZ4h3OMmkYQY4SYH
E/AqxVSmVPDy9bK9iVJn0coaRP0ddSwasb0Zukqhezp7jzj2MTw/AOFl1gnL
yyBFuPHfcenOEzSYAapeG+QA0IG0nvA3yHHmLv1Iw3WyuhTRzie1d/Ph5ujl
u4bEsDB4bp1AsBdRJdAlYSCUjFj1Mhtkm5j7zt5sScGvmyOdKRGeKEe6cSsx
8dXpuebTxayujNcUOmT6qbl+CB5i8jDt8SJEmvGWKHMdMS/B6pTgyIzVxCQi
jPnstUtCm+kjbo6qGibRYgfa3fHYxa0jYA7OhVc8fhhCmeKhk7KUMNpvCtmF
MEAtHa9fHWrpdf6lfX4TxvOnXOeayGsuQ63iwCM0XBYuvWmZLJmSXMuB4dqF
jQmRW9oGnGX1Roh+izT/+pGUjRr222WPbnPnrbdG6mpn4D5BPERdxMfF2eJk
gwLnc61OZcYqjb0u7KhSDaeOIgtVScs99Jmdmp4wva9BOfSFJUwWUtD/MO9N
RxmBP1eNfM5AjnuAyNgXqQM7HLuGHxFDyWabJnJlJCUl8VKcsTogLqPGv2NR
JQGo/UruFxveSqY1W+yTvjQFxgY5aw2Be2NaqUa5oOeCI/EtBYyUBzzRiU/S
oGBcJDN57UNc+M7B7EStNh09hPdGjVHJ5gZvtVVmnir5JYXWryGCLtK5tKMA
jw4lOyqejKvoyuasRfMisuTqfxzZ5Yq7xpfDebjAbALjRrFDncZJf9KFBENh
9GpLoPnpBj/avcnyawiYqNoEPt8fV6oXfA+Dz1pyPy79zSxp4xhZf7i5iaPt
2XO27PTTC//4szV1ixhkxcxmIdlwov+fnRI+9XWPA1UD+cETlXy/EqrPQ47l
l1hf3JKOOfBaHh31T/0mxQ93ilgnjhXu2vUhqnzqb0JtL5JaeGHIGUpYW2BJ
kVFpNqM/p0B2As12Brg47m7GczTAVPSDdUq6bUu5wBf+XpyCrbatslfitJLt
YuCKEWZVJrKwqyyaL5AV6amYnOOmXYriPBqiLnpByMGuN2yciOpKWYgP0EPI
+YGdfXCSu2FyaQ5+txQpsD/1PUu0FP4PqOSJ8IUworzhubgFJ/ZTlgltpye4
mnEjzpkcWQYYuZJS+lsoR6MwY0WK8reWsr+37IL06yAECxAi3zbEiOG133OC
VkvbXdkZ6sVAmH76NnLkTTryKmi29lFLXZdTayfuMEnbRqqDVdOa8RKmtSyH
wOWARcmDZRM4wiC/G3fN28mH4B9TEof/KqSVC+UUDEUPSvPF5bAOWl+al3Zd
//A+NXrM8mUkyKJ67bmaTkm0A6AWcjrnVPbHxym3QW+Lw5BIcVOWGI6Hxjlt
mC7J5fD8g4XmKug8VZrmS6NmV2dA28XELkBBDujHtoVMFUIv1hFruYej/vFc
AGqv2cNZL9uV1j8Wj1NzwfoCII1x5BMp2QW8TDfGRd6x/4LPjLXnCZLRFhJ0
6eF9a27Mb4NA/J+Uz21AGVAIjJ/MN4bopbsbP+ThNY5wobwow5D+nivZwd0i
fyRXrWluA1DO0jDAvoib9LKI8Z9jSTQfLSGWzHIG0s4YIFwhdWJGF0mI7M4E
TCzwHQDLliCKpo67CzqLB4WZHYmUNVKkBSnPPjkzsj9Z4apNpnPrV7IeRAvD
jhmb2srEYStgz756FApaK4tTzLQ9PSyEdBAKvMkRwv+QCj0FgxrnNs6Rp/FQ
KFrMja4PH4SPZ48+WrsI5gaFehI9WusCiGJRYja8/SSrfdiVQO38IU0ZRuUl
88y3/34wuCxXOLRjxXetKNdAesf1Igx/9UzUpBRR/BYoncAo86tk+tbqdfYO
klg9JIv9VMeuypkZ2et4fgXsQT/JTS32kNxQ1Mv1M3QNYwKADCGFX5IPx/Ff
Oq7leLLFbq9hoEYHLBbMf/WqagBY6U7gTBR38cdiUqBGF1ix83klWWLS1IWy
Ivs/zpPa3/nlxJIoE0e9beqSPRv3/S/YdeU1HcWfs+A0hdO74EhegqD3C2Vt
D4eTfgsLUH5dv0MPj0vt85h8P3FO6c5XzJj6jZqd809W2RTMXUUTxHUZMqeG
5eiCqF7v2EQMjucKWfOCGyWmzinD0ADscRTTuQ6YSojifIxMkp0dki7FdwGT
kuNK2cBGKxEmddwUCVsBvvf/OU1rLyl4EdfXSDVGg0ynpD02qA2uNf5j9KQW
WukI53ZRYlr4MxELSzQYZ4L6p7Qo5aC+WKUphaaApt3PL4b/hCQcocFWFu0g
+I0dzPVh/PB/Qwc6vUWZCxGChG2ht6wWigRJ9WKph2ucrq2r9+qe3I6q+csF
J0yYfEeIX20sBlJi/Pk0Hi5VlHmVcSB8hfsf5wm5ZoukhnAv3sLRMYr8U9Df
h02g4POil2TNUDfFFCCvNax3Ouwya21DpR4mKdYhB0C/c5j4YqSdiWoWRbnd
PAXdG5BeEVPi+g8PO6p7lVVQC6iobyeqUVaEABxYG+iNtCH/on6cjlGKlwkh
WP6ligFG9MRzQLANv0Yr01BODEzzRnTHT0ATYZSePrysoXiafA4IOpC46Oh+
6ltcOQhs5sKlg4ELTUSkVfxo72+8GqhfXbPwgc+63kNwTa/DggDdfr70mho7
uEv5QUixOiofCOuqBXtAvdV8ACZpUTyzG4MgGeX/6gkbrI98Oh/o/BP18zLI
aK9kHIG0bOdPMArXbzWbMT/BNcYoXzQzg7Alkr95Hr1LaUQKQP8QSd6ryMjX
Gw1gDP7HjQHpgz64fnWPSVWThTsPhyUfItQTlb1yOTH4IPWY8kMq6fYwBQdb
tc9YmaIY9gLCjO4g9wreoDy+15+q9pSyn4w/hJWXdz98Hs3ly9P9F1aEeqvN
UZtnoRD8DuFlNbrK4cWjY6fyumPctPjJcQGaHpH5uOWDw5TRC3PWUfx0O3xh
nIESJ8pxj/1IafjzdBfMC/r6Pa/CTY+ffSPed7/KsB1qDLErjHZRzvzZOgAT
C8tDsoQqUDHthg6m9FETpNl4/bNJMAHOX/cKY+ZoUDEr0HaCzMsQvTRakHvV
eZsBoPokOlxrS4W/UEdnKTrDkaryO6QTRgVmMcVAmuDAT0QtuhbmVTI8Drfd
eiVs25RSyu+BrqQzVosHV5cvf49+GepIWrbGdK1LZSdIUj101f9IpZUT/pLx
T9igZlwzZ/07+jsv9mh7+7v9ariJIO5xoJ7xA+qDdb2/Hj6W3xzz0OwHHTrr
ec+vJwbly/pbL4hPqcrOAAWN1stIKJdeqtRH8qPi59HqghlOC5hky1gARk2a
a3U0mx9fnNySjpKTSvgLxdWKxuBaZuD9r14Nvj70jOsgyvSuN22Z0zjZ1eXI
0N/XTmWOZQI81RKX8ZaSnbjx6/4z/bCE1OyJHfsHT+bqECTMqiE2XgAs1lGs
T8Vugsdp5LfRB8wpyFv1/UutAyTX2Ht9W/A2Ofd0C5xNX1Z7SYMk4GBLvNO6
Hc0jgRycsqdwnxP3reSgBSmd4VRYiD7JzJRc8vV6w7IJfLjaS8FXO6FS9E8o
QjOKAHhL0KUWGYach15pBpO15Qbdvf4vf9sl6GCv2DQOMfS6InsEzT/0NCtz
FubnrqkEQDuABRMtB8Qp8qqs/rWsUX33ZG+crx25P+zPtPq2BwXoMzwtExC7
CaqJSXzgvpfSStVPtEyfEYiDZpu2y/3QJQxmIuAGfONLmnHpcNyDBWK492Rp
aT2ezs4Uxa5WDopuRXihqUDSGvgAvEOuGkRs075tgOAmjW4/Yd+FLye1DYU+
DIeEylRNi5BcEfC8DT1fBc06sPpxnVnLmVStw0afhUb4qNMSwUakP1KD+58j
lRRBhvrcYUFRX/o4kB1QOPH+yHlV0UlUYz/B+B2ssV5ZXaaKCGb6+Ys/Tb0d
9dvGSS6sZnd4RqVmvcbXlze6HsOGw1+e81Bu0kDAih3cGKG5ZJixiABxwaCb
fwxl/lkxPajeNsaI1BpDF4fIVS7bCeAmKVFTtJ91NNOXDv2EF9M0AWZ+K8E6
o42686q6Fx+Z7jUCfWa99CRvFPjhGJYlcx31dNhEzIxZQWZ00oEJq7yWalOk
UBYtout0dj1R47C4sJbCJmU+x6cqdIaWdoLVxn74YmtX/P5eLXLit6WVnNxz
5L7jNWNbnO7lAxpBiWOrQ388/YTvqgdJrhdtJ5jb0ybG8kclmiVNfKhaBVhO
com7Brvsl5RIXAk36SPaVHv3scnhRTmInxfiPOSo6nh/wmnNjOIrFEd7g6ng
DHc1UD8zO7q8Ki3nktW83U+n0qER89Zl/8VDUDB6/g7p0yxqI9PCrljit6zh
WOCpmhuyQlDku/HEVzCdkY/1kReETQ3Gh/hQsJuICCJDaXUON0T0zZw9jCIi
DowKcuLVjF4FVZQQuFLDXmGN7a9PJ5bGyacKVeQ6yCjIEn+d8ZfdGgSHno3G
W33bRvmBkqfsPbXmPkkEmc/aTZLkM5p4QL3DTKPw2gjDvYNo0spOZ5mI8xNO
bUFKTzzJZ0xQIA/aRBW6qfuX81Y4inatBLEkRxS5CL21mpnwJf7sM4xh6uqM
DREPRcP6fFfvhMlFRVecdv+rJ+RTXAuECZcc6XCZyzXwhsQ0PEkjjauLYhTS
UO5aPrf/7KPMrlYBXYkLF/6iRn4ihqAfvS6pp37Gl5edXR1j5iLRPxJFmuXF
JD9z7cjTrKLtzkESeNwF38cNQmjqtJ8jZPcZW7BmBacjfe7p79UU6DwQW1K3
3bJoudGtFSitR5FGoQZtgDxhbQcax6mHGkJnHH6rswsD28mEdpHIh1dxUtV4
RczRcoN+cQg/00DPf3wQg0ZWwpTMoACELn2IWjrbkvU2RCmUkmA0ode7Ge52
LVgtN6Q9XRQ2pHF9PF7ICKiZqIPTddjNyXLywPFEqm3DDoTagzB8dABpNomu
nT/yfer/REnOb9YUDYS69FTTCVA2oL8NCBIsyZkbZJ6IpDmUTo32YsKAlq3b
0MNS6O5yTpqmwNKK+b5uf2F21V/NPQqTWx208eC6CnnYTE4y8UqI21XocUt+
ubg5cRPsWJ86BrUtvXnn/ZHdodqsxwvPJboarCJm+GjNCc+fiyvgsKDPK0jZ
3u1S02KXMDh0EdUlo0rzOiwq86ZS0mBo2lolPYv8rNlbVnVysm7UiCgV+DeP
Ql/pa5b1hkTJHUiw14Gc4C3qg4MRoAkGQ4mZF6UUbJYVdTxelk8z5zBZVzPS
NOwzkrvbimcEb2HWcElAWluhKRTPcg4nSGsw66nmGPOcCdyPYNpFS+Id8Fiy
c6M/zkMLOLVHENN9M++XsL2d9krPrwrzWvr/R1tWypHtd0qahPWVcSyWZVzk
W9vrMKxqeH+fdUNhJOUweSYbGEpC+r2Uuxx/GJNrtHSNJNK+HqNEUgo+JKeS
9ZkWYg817IW+OF2AYl7J7Yyl2heJp6N5G7RG8Lv16z2A7JFFcqodNKBz5apa
LqPWDn9fMc0k2h75DrZ2r12uRim98NuAhHiW2sGl2nBWkwGEVbI1l0X1AcB5
cWTcZdowZT3jEjJKoZdZCySxPjxuVPZ630ILj3RvKukcvGI3qoOfwlNglKXM
DzO8+0r/wkbg9X14A+bWRhnSZqtd4PhC5/2ihalaPWjtB6T3TnU0in2yK5ms
Jbwed9RGuZxoD55W+z/1fYoCVMCjEDYOaeYrfe2eCB4STG8ok7ACgYCJ2Im7
BKrUk/ZeLW3L5wz/ihut7JKP4AamuIQlagwbvcDUvViYF7FoojWX7BgreYz9
JYrlry/j8o51dCe2lq0EgaESuv5nnaWcp2mItH3IVp7D0ceq7gJx+zBSwYK6
07/LPUGDG1KVYFMrZN7smbQ/LohKhCldkQ9CMtHL1dgk9b1WwrBEgsrpR4vD
txtyz5ThVjH9CZY+x08l0okckZE+bEtETz7VDWA/rgYFsNdapxTotK1/CkVt
GNHj3NbS0pczKhkK/QnI3J40BFnPVRCMBT82VH0d7KsT+NL5mGGrUN09aMAf
O8xBiai0cMxILLP7a29rt4pnX/S72r9IedTkYnZ/R3Rue9dfq8mMWPWKG836
GvrpSwaD0+AhLyQuPIf/Azg46c4wQkCb5U2Iqjv+U8CDIrc6VvbvmYqMWDW3
KnjgdgC9bsi4AdAH+EEkNxjok6YS3k1bn5PwL8jIrnGXzUbN2wvxuRlXOe2t
kZyWAPPdoraqH+nEgsl9C7kQKaB2uj1WKBfyvqS6jptlgW4cJC5+jFa2Sa9Q
bcz/3tQlZFe5PJJzcKg/tej1J+Fmo5AC0iZtIv92lwWn6yz4nyjGDTeIo5jU
P2TVKjYpKp43w1r6CBYbhPhuO2VrhXIxbB53H+g6TNo9WxjhWGHjproDvqW7
j/HfxV3j8JD18FCbGluptaPIIuBn/LyOS1rn9AthBlvmpPT247Gw+RAHFTJu
6lc8aPHgP6gb78hksnl1CF8fbnTi7FvJ5zQ+kv8vN7ZCOnAYTANTErU2REUb
vtbG7ycQKYKbfmQv6brC/4dWJs/Ahlf4NTbf2a2ISqCf3wsXvWF9qE+KFoyA
feeCZEsyuLxaSZdkWRMrwdHChqggD+zWR/xx8YVRkJ7XPdAMuf2YSciQQw6U
U+7Tmay7HpSwd9aEhHrMZtqdbcAENlQ6PSIUQni7gFrhTUUIh9lh/SZMFbQ6
fARSbOwinjJUqHlhhlzGzRfa2NAtWsdMLzDZmkSkiYb8pSMOTUhxs9Avxec9
I6vu4oFwdcOaQ3G/BNTz81NNvR1tBAJHPQED1H2e1WRnYoH/Se9dOSzvVyDs
lFqCjbUtyihVtTlNfOgT3SrRHHYN8D0di3/pQNpTJ48UmNKrk2cs8fZcCerN
40b/fRSIQIJCFmAcAlPt63C3G8USkzVsuF5E02XK1NCJLExZv3I+mNZqvlff
dPiMgTk+cR6CrrjJp4CenoknHl+5YVhborL+enCnFfwZip049zTSgWNqjVFn
NtDvI4qy4lLi7SQOok07+ie0+3A8UqJ1Q9g/gNgYpdAMFuh0//gUgJUj/2l0
IAXvzqTHcVuABeHeyUGKgoXnteI5dGKBhtTYak0+62+khWglAbJZWsXmD9ne
wVJAypgWI69rsWyNuiU1iB+YXoqMxDkYz9nmZp/3zPQmQ6fwj1mDzINXhPpE
hJcgy0XWpEWfGNCCiIDUZQ3Yz/dYlrKvYY5d9iFhwChCZLoEkhyGpnUIqY05
HyuvfkNmo33IOE+OCthMPzfQ/9t2ZL4mPpwiIZtRMiViaxmzdbRji8rV6Xzd
4fv2YbGaUe18xiaiMGCWOfvW8yxdWqhS+VG4P0s+qv3BAZKzwh1ukZ6KlAsK
amCXxTN3qiuzUaA/kJSImVovYmwtvYf69G1IfBiE9Eu00RaXiDaLRYvvpbxt
WAqJwz0rtXVuARAAD91ghXYDUZvTe+GUkBlWL4JXxjvMP+TXghA3+goZVP+e
euUC6onrIRUtA6xSimsw4eHV+Api4CBX7TwQ+c4jiFDGuKn3pf6NpSwM3GDb
Vt22Fy2R6N6EAElTf/fGCTrhl27a6XCSbDypoP/Nx12ndK65hCFU3DXkgFkt
3Nnbav9W0c8vYar0/8CRHL0WibF0imIeet50UPjDn3m7pMR2fHHEFhtp2hm1
VOMW+v3jS72oMfLho8YXbuWamOhH4pURNF/sOh0BwuJNiN5ffyWsEe/Kxh9O
3NM5PZ65FdebdwMrgS2jaqPudyPqNZYpEL00BoGgDgU9G7Fm8Z0Dqf+2wHzS
yVNJjXkbVLdil2c86fPfYa+tuswM/peCC6Vxl+miawVr075tgbB4Ql5NcA0h
6W8M9WypCK/SWPCUj16Eftd5MjgT0ZdAokb+AWKJ8J7cZ0wlL9k2455wWcXk
8MJlTvawSP1gMWM8kpzGhea/Kw/AyWvmLh65kMt6zrKLXd0EVnt4lF8WVE2T
BawrHzRX+kXsJhJXEnUSSRBCV5irAoKWtQSqzN4hORVqPHFn6sNb4d6F2ZXC
ieVO5Icjl7cO0Fsyxyi2kGCBffrCEvO5QgxZKeTfz2ELEiZJZlXPU8wzWdLv
jCqy6xwVoalck56vBAGVmjGRM1ZluVqJ2rK5kk25c2PrroXOVK8qOmf1GW7K
KSrE1iEZ6nfegO0hqEVL4yHQ6nbpdF6LavLAOq6k70UdOz7B4VWomrajkjTW
I1veCqpZITzaVqUX8AdZUWpsyZpKbF/bPlzh5XbPM0c5URAvQR4il19JZqxj
Y8Hwc0aWyGJxopFYi6uEptx4UyjEMVE1jPvbRQInVU810l2+VW9xkDvYarql
jUra484zIni3vZ8CCuMNvJq021rw1ogKmq1Ek5alLbT0NoCM/3OH8Dss9AR/
1/fhJlxgr8KyEYbCj5mN2CO9NK++BlzKzzvtCmpoDeFzHPmWNv8rk5LOQjHK
ifwkNOEg8ZmGhvTjFLykzocc0D30KW7etcra9RWU885bg8joPw2YxCNQX/AF
K2W6zPw8qKPX/WrC0GdYGmQyclbjDhmNejUYss922hComnhE+fm1E8fIRMRg
E+X8aI0xMx5/oxUTXbrC+wLeecxHZoASn9vFhHhlFw8w9ie/srX6PTCKItzY
aByWOh5FCKwC06EQ2Cwx0V6mgKx1K4Wo0nNt2zbTOw4j5giFpr0a2MEbuTtW
BFw8qvPsejUoCpO3pWz5ptuYDneWtpr9F/jYKfxUmH4p/EAsGQKzNpwWN25V
BbIfspdyr9QeJU7sYl/yt++zcHw2VtSn3o0l4mbGsULvZUQ69mSAgPmO375E
lHMFR3tTdIYEI9k3mJlu7xv/vPhEmr1/a6ssUx5cGtu9m99v5JTSIWVjWbQk
87EJIFAYE+kQ+0Is547Z8CQn8L5ByDjnAmI5+z1Dzj7VsUcIiJF5zgVAXfQN
YX3eyAaDnqOObyN44UE9txH8kZFZlHUveT93Swx6ki7i9KNQCAlOVafB4QSx
kLebpNMMXKjcjMoTIEq+ZSWJ+9wJOIjGXWWr/I9Sr0XnQrzmCC20Zr/1kVAQ
bnOyTyHmoZn6S0wdRSYrXfCOhBg/tfXf5LYEQ4jsjQI41sBpv30hFawerZtK
fOa03L/b5s9/KhkYz8v8lbbYUpOpSXJIm6U8smWM35yxvUNwR14qsVO/Nr9l
fBcu9pZudo5XQ9u7Ly7edPv5EG5CJq++VWokUFfHl8LE4Vx4k+GCCUIOtRrT
puHJlDIb0fQeohSTd3i7FIEZL7eXR8BCgjzXGTqZbJBe2hJgcDpveyeKuCu4
RZJjbyA1lhe+hWlQK0HaJ9xj1zAJ/Rw4hqaYXpt+81e824iyF7YVAU0Gl6X2
hQTYP9224HP1DT33xsmVgtE3zP0Xs0SmhkjwyOFNcmpqaCu84cqlLPI+vcP9
FG2a4sz/7hNCqJ/bRCZkz9kAPFiiQCmWSj7ytPw8IO0ITSsTKx/eXcWM6Zm+
1bUqWF2kih1r1LQ23UVwuVny9Zx926E04x2CroOGEsdMbN0gfs1gCKSX+3VM
Fzr8pZiv05IFGLbumfiZ99zaCzrr+ai24VD7C61X2DYwY2zA/MlYvMvuP7c1
7ze9hbyvpK5dF8GPkLIaaTwHORZlvyxI1+PhWHDCqwnAfpMz2gLaaGTfaYpX
5oqjX1qM48spVqDXBuY8h8hPpQGK2worFMYjDPOpVyPgRq5R0AUiwAi5iQKL
7XazY7SvTCIv/cw/IZUPUPRBrByWGhNSYVG8LlJP/sWqiJM6CW5lCWd+hzlZ
Q5Y63Dqj33qx5Ey1hwg1iS6ekUx6s3IGuwd8BbJDSRB8P/Ohy0arOxOiVeA5
LZ2vRRIVZwtK1SYDZMhq0VzRVH87gLEk8ptrSAtJd0vVBr02arm4ZER0YB2y
Y66/5bWl1QU6nGtKolfVRFsExWq8STs2FfCz/ZoKjCMAtqJvynCIF5ajyzY7
bcHCwMVfws/j/I9lD3x8NLni39ZPc5DMVUMCAKI8mJX4gDhkO6KL3oeG0Bpx
D+APQphsbmaMNv23vXdo5INmIU3jFaTNOr08+SCfGEWG9fi8usn9lvQgmq0s
3da4sCDVMRXiagQ5gHkd6LIC5MdBZnTsaZyIu6SUYL94LIGihRHSfX47DA04
qaIbUn5a6PiegcjgidB3/ZO/jfrfnw5y5rpZIs1KW5IuDNbFNZijvMvHf16B
0xMRFnWJLkyim+clz8VYQ8NHq2mMwjrXZJjLZZUnHNAjoSg8n7wRT5qhDvzw
N74GmtdSXrM6czVrGXOSBnZLS1tDho9A41LBt32akrw6dZ7V3n7ZOATSH05O
lMhEOFSPJor60tnukhjhmq1OG26ZJHvs0goQYVzX/2VA6ZG22ojFbkC2J7kH
viejWAydCJTYUAqu3ZhVrkwewFd/LONqLgQFfjQSB7Erat7kA85UDiH6heIL
gz+eBm/EDoYjdkUyya9cZ9KwSAMLR5Bgq8PCM2XzrBGKj9XRUBS2IqNPkKQN
RppiQsqumln15GxPhePBmvrVTQxfRuqRq4/9mau6YaZWDn5DM0A3WoRGrFaq
OPnHdINycN1lYF0M99pMBdUEUg4gajvsLCXMTV5wtRCC9ZnvioZIA+27fVUi
c+x7ZpirSNvPoDM0mBMCi4GXXtbouoAUsWMRMnyfLUCLPqDtvE9KDK19CCBR
0DB40dcjT5V3uYmlabGk7JVwhwl4ui+kvro+3ML0bbKfp2CagqF7sCgSa4Ma
tFP36eBjIEUZRLXvasAPdp0M2gdCTVPXNSAqdvHpDIT9bHsOE/iOX03r7/tI
BFu7jMCjbTjhlN4eX9I1nWaBXz3cv1sPiZfwY6GeD32MGEI4abalfytTRcYq
g1QEBa8kl4WcRBXTpBsF4/26nd397kymXDAXc4XObPI4kwHQ9ftw086px1g4
WRvR+NJORam/8pvYz/LRUGbDQY+Uy/QFkd1pUeNxP3vI3Pv7SojJcUBhVl/a
962mqGvtLNWG3GsCJtJ+bA8saKvnrzTwLryz1x+F/8iTSIeSOvKK2GelznjR
jccdMNIqfWyXJp8h/sYfIyLHwBijwSV2E+K18eqc0s+XACSf5uThOzhqWEwD
Uggm3K7p5ju4mQZ3OBNB7KdxL/Mu5OEBf5cKGwYEFdHvbHnFY0yH07oMMyHo
QJZ6R625MXZYCKAZXUIzD+Is7zjrykj5l7VZAhBUP3E7Z3iCH9tfbrHVz3G2
6geJQi33J/+Jz+7C8wEyD6TrZ7U75KsEQI0h3zGWdHrmYN82mczJZeQBYRPf
JLpGhRJhZTNq4bdrO4mSTJ520Op3PQ4IXWD2kgZbFE7RuoSSwj41J3+TPjOI
PAnvvSgqdUHVVXQCTJvWyg9CDRySSMuGp493GUKRfG5C0SrV+wGB7ferKoNU
J/dhVhUV6FC3rz/QBBpe1DJPGOMYFejAL+KFUb7kZO0VcrAOG1fTy8T/6l7v
iaBEPYJ5CpINrTbyeitUXMolfcBXey2CbWAzJoVhO2i4rR9KQHZNS3VL41Cy
/PUW9o/fr05P3uXNoTRzLyuv99T3iYbwzua2mD3du+XieV8tWEiqH1wERlx6
TLS7bssjp84KsLj+U53GTjy4v5bNQ14VyFSPfF1pIGYZja9WD1CXarZE/xCn
xo/Z6PnLi/3rcVlfeNJr5aZHM5WpQNRyvh2vPxhgWAkbFUII8dTR9ipF0zFy
JAxNdRz5Lym8Sjdlk+rAGuh/sMbyxnLN21L2qqZEgzcAhKzQqDTJBHVZkgjF
WOkKMzjd21HTKm1h+Cn2LzPh16Lyn47cQnRPw0Sb/NSZ+6eWDT68aCsj86ln
dUhOcvjimMdJnYtM6eGAjykl6x4z1z5xYJinV44Hs4NAvfuTvVZhCuLXxi4q
LonxWURMAwdW9a7tBRL4vNTJlKPhi9N9dxkXf4QIQnbtMMspamphJPcxyREn
D8wJ/sIavvQ7WIews1UjPIXudKV8mrWPfrE6g7rhhsvm19VHVUIMqcUFmVC8
VUXG0lu5mJeQAhPj2bFI7ododR5xi3mlxasWc2pcq4hIOafHHAc21lPJP1bE
O0VuQdnlOZWBCnmk7yzOnMB+3Pi1eYgl/dylmd5wNPmg8UfcJqvvNjYi6H/N
HDmKmXbpP4CcFoDnqF2N2QtCkknczw8pLTm96bXqxT9ZoMdr9G9rPiEr6rD+
fIM1JXWjjWZYQi3ZsRMFtFj3TSCwD1edVX9Je4sjCVgTZDQDyqt4iZzi3Cw6
ZSA4dh4P/BlkvMrTEmKn6BnNZJPFNMO5ZxEfxsDO+wmW8p4LeP4GomcDC6Uc
2UNK6xHidUmb3TlJIOf/W50WLgCyHU4VAxCvV3FKato67h2L0xJf2SFyR35V
IWBDecA1YpA1fUlGJSjIDV5Y2iKnNDKzAvadits8B44x+upO316NDTYgQJiP
ksvBN70kSEHdC0EUPgX+pFXaHqgqLxE7vqzfhBr8MsHKgaDXWQ6kg6v4lxoI
8PZVtFLyT4Dj5B4/uoRR4j5YXP3l8eDisZSROd6eOAN1iSuCM+wDKFac1reH
bVragEgXr0wbJs0jia9pR0oF8mWk91OQNjjRWd/8ibFhA9wrVyOM3TViOSqx
YE4uBt7d3OTe1/hrs8/lm9XY1PqeB2gWKWbVDo5J7V2FnM6SgPpJJGiaqFo9
UNEyMXl0o05KwjUXav9aua4IbFpzJHtyxfGkptM12NSvWqPN/Pmzj43oeCrI
KqmzI8se4yyTGyIdNErTuvSeQszLAOUr4mXj6oAHlUYxOF+53IA9Zu7keUHr
Zbc9WDdPqMKJrF3qrbkWe/NFV2WT+QQj2SqzV0ybTdKn4UfJndxhRtMV3sVJ
MDY1f6V3l1ATZBUiO5Q/fm8s62z9YYjo93JI9gfC1j/kkKvYZOTmczfVo197
UajNObEdCs22TjNMsTueAH4vTyYSvxkgX21tVR2GePtnAfBEaUmHOgOEMXVS
MPd2YnZirdlEvzTzzxfStSzeRYUb0vOa5DD/BQiirMDJ6ivENxeR6+rcec+R
up9kibRB8CYP/lbXpOZRCnj5bCmXhks3QG0zuVM6LsuRBX3KjoHZQh2RL+j5
RWenBU9AOXkOX5OvlXTLLnoQwALfUnbZZ46o+zYtEqo4eMJdiuch3uL+Me1d
vKtIP1hVUuHkX/Lo7WtnTjHeO3USQSWo+mmFNjmUVxscxeapay+Hal8Zk+up
ms7gDaiaqpdbieTX99EBAI24ksYHAd4mMzIAZAERL5SFg7KJM0QeDi79e+vW
HloQk0w8/B+gJXVvrI8n9So1Wolzf26GuDspuzKp/jzgd5wQadXqodQMgL1Y
M5OMOHohZVvQo1GcX4MFjfetRJGRK75WRt91L/82QWUTuezFyEpjxKCFoJRx
dlQ+fquGKUNNSS2nl/IU4I29rcHHvoOvnKS8rogMoSC3zELqd00JcopPI1PK
ap3sibUiPhjlTLpcA178cDqwmlNHwcfk9uw3XUdkaJSeJXcOTRjiThMCtFTa
fgnSRLtInos4QVc3EM+bT4PPopzZER4WDSeDGY5TWXa+zMB2BSe/aMVsJ2u6
1i30b4xYhZO01PdLU6vvLC0HDRbG/y9ahcdbloL456Hm6AaJxJ8wHGd5tNFf
J4nLuIGDk+Z48ZdGeLQCtuVtBmVmXHH9rl3PjIrCNU0pkh1x+ywpB5sRgwxz
zt89VIDfdVOZgpnYhM0uxHvymkc9jMDWDxsu0jVATnhMXO4mCO1m6cTQ2aK4
0V0MtX1LCFquXwfqDFwQuzXJheSJbTnIxHqBrJlpepR11RFQdTRkjtEbg9KQ
QmfhGPKgn/MoWNxUe1nbgdkrzj9m2fEHYfMKv49f37EiU546jrALZOQ01U8X
3sFSqCLWeqDcAiqf8VnfjlKkZPsQVCKQLyn+yHN6nwjbvefvG4kFlZ9G7pLV
gyuDKBHT0xsOEEOTiPOhXQRTDC2bofw9ccXaVGpDm8Yk4E+G2QxQqEiIzkqa
Pg6G1Vxy51XQND9PdV/iRIG6FrbOyCWBgUQkeM5t91eWuzHHh3dDky8g0VEp
rjtvkGmz95PtNXdpuxQHuCQ71O169rQVEBt2jsdPRSkW/tfXGglVLUlsoIBw
nWhWgxuVn35Iw1XghFV2C2nLaM5zJPL7OmKKiqunOT//BImHBRztCvYKGb5d
o9GkKbRKrOmZHaarkYaZRYrF21RIieExwnfBRgP7CoHS24X23VGl/RO8zfL0
qH2MF1DHFfvpWkVNJCu2MMGZpoYuW724lrXpcwi5etpC55/7BqVdkFPHfezh
WY+negYRp/IsoIsbI8D6iUjKmROLF5ltc8avBWd0s2YwZ1k6EiGY1E58DhHC
JiPtNfZlESXC6BGQMuSsw553Grl1trrTi6E8gFZ0D45J/uy/oVhqzAh2Rsvw
zL/rg/HedV4Nh+BvLtHuCk7xhaNiIcgYYuK87NokwMMDBOSpNf1+sXvn5nQC
HzpxxgzmjgC0KDnwDc/N6QWwU2p5yfPzIMsQ+ou9vJRjAdvrzoDXmi+LawLI
MfAPuU9LVsiQzoCQzYW/Dg7XeZWvKVnnBKGdcTnanwmO8aDuScfH9zrs89LD
puJWyeZ0o2ZvQ5sBkGj+jbRaEEuDNj334HcMGZAmxOGnt1Ic/vHgYoE8SbDg
5J3u0DjI3JfDA/dFnZUG4tx4w/PBuhFkn0+bUM9rLdlXfAON6jB4KaaXTZu6
IctsWb2GAQdOHCJCVuBgraHZd+YnSHftoWR/qRIRvARkSst0LBQDPbYcWw2a
cx1KNup1ymi4Op/0ViCaB0f6ez4Mlwt2KEUYi627pXKZEWFZjgbxivE/3ndr
mmMsXkCOJg2Dgd1VcjUYVMZggTW4OfpO9jstl925d5IaOQmsyh/nLnMdRQ7N
8vOrBfKy/0oZh5qYYwCB8uqvUGlCKhmuG2/ajyTLV6DMdwumO5zUM7SMFkvk
TTgsJuDsinXpUczLz1AFqc1nlTmOGSnrPLRJvGiWXOvvRfLfIilHGWcTYMd1
A/MKeBtK+/uNy7G08rTJ7Yec4ruklG1xKn7n1T+1dIBsWJyNrC+M/L4ws/GQ
ABH4NpwTzE4vilUIsA0R9fSVuRgFhxioZTxi62S+tIDdk6f8sQN1gq8uBqmM
LgnH4himho8WWM1thFHQSK+zt/d52jmQ74xzDPKTdQs3vGKO53EZOSVA4jfS
t3SRAHDMzIHlLT82Sp+YZ3cJJ9heCNzZ0i4Va35IlNaLbJWGTHJnslfbBy8M
JJ7izP5In6JtblcmCE+E4mFQmZb7CdvQ12DcUepL2QbbVbrl5s03Kvlz6cAu
jlx1m9hhiiOGrUdQNikGDQ7EiwsbcqXFbDo+gKRwmyDp3EbZWRB9O31xwfpJ
6BckCqvjRWqT0ipuMNWBaH2BBFdLN7tJZ4ZoKLJPlt002MQucoHkDd9zpz3s
zLXzwfJMG/dVWKCn3laUrYmFSgAtJFdoSCijUpZ2r2zG23XfG2Arq/OsIlIt
wJz2g1+mgoFW4nYO/k3e9cuI1KcimIbc83+tbSFxQrqIeuAQXBgxzHFEz2nQ
FUJl5NYNRKswzzu+WjR2droLikfawpXYOQ7Tei9yStkM9X9q1ZsY4WZVZnb/
7IYF5lhW1GYTaI6ofk4QjlaEY8e890Fsq3SNfEcWwOgIUGwyzIeMeM9E9iU9
aAAcMj2mOMdn7J/UUDbNqn0yvaTmNonQrrR3jp6eLpycz49QefZoVVKxX+HM
dtn/gIRI0iel37AD1B/ZRxFdML9lrOeJR0pwW1NPzMv3zUxGFw7elwgz9zoc
6g5ULjrqTgGWpAhgtqihzGpWmCKw4S5GpVPFe0Jv4nSYS9/lmdksDy85fm0/
qumixUVpy6aZPoPG0vw07QNbfSgt8O0uyW+v7NiqV22Iq4lxzR9knasPusdH
OnhbGJucz+l3GoGAWwJGj4Daqn4ZNm+ES90FeOWeqE6CvgF8citTMsN536nV
fMrNSLatPl7OV7CatY0w0zrnZWrtXhgoqZmz9C8RlXKq6R4VpNfzkcAPo7NB
ur0SY2YtGQN04pf5GDs+naFD1trqjzFkgy1mSCRGPJKG2IumVidIH17WPHsP
4FZ7CJl3C7PizmO+tgUUZMVH8Qo8UQhFSW3CmNWnb+Rsu44MnuZlNnYsdiSo
jkMT3SX5cyDQZqFk4HgSA5obC6yiHJC5yKdJRfHA+MGnP/RwZ+oPHgiTvD6R
z7sWX7wcHjxjX+cJOCqxM+9X0YoOeE+WAWALz6UjeCWFs2v4xLx/XyNfUmIm
17Qf38rAhCO6wPXLDSDb3qxlEdnIJH88Z0uw0I1wv3PBceMtp6AT/AtFJXbq
BB+fTCbWZ/iMXsX5279hZT6Gwl29dI8oeA5MT+uspkYZ2qri66UrBqhjfMaE
27A/hdMIzsP8b4QsgBXcdgH9tY0gdwQoDR6ypsDLEY3O6nrUxVrORkmrb74V
WYpcjy1z9iTqvdCvExgQIOc2mePajHmIiiQZ4zA6ydnPHFUDDLb3DAZSVCYm
RWKlD5+bHJBl6Wr9THjKbsLKNcU7UIIu6+O83HIw+eghtJvmQYE6E1RNAGid
JUgyMpElTYuAQEnzwfWyh1/k/AdqOJCV1lOZn5gfU5uRJJgAHZVS1Ike+sM5
a8KW72DPjLvjvsvjalKpViX+iSPAGVutpaxWarym46HE24aQt29bN9bryuXi
+2oF3cm/dpB29UpNvxg4pxwWUNDICcyC60R0H1EQ5ng4Lp/dGRJ89Uv/wJM1
QuBAY+Di9W3GDxv/ZeHBuhY95TMU9pwGGJSGxvc5+XfkpjlFyTsq8BUfDads
+VosJ35H0W0L9bd5MidULXTQ+LeVe/9nQX63aNv5JHWVijkcItFBjbiXhFzf
AHYWTHpaotKUHVWwNuR765uwzx75pb75LgPDXUCh4TLVlBTyZnnmVo2lPOjw
i1KU9BGCjPyk/PDj4MzFEHVNY0oJReKnp9dpopxeqFw5Bq/VQtrs5eBCTCoW
j/rbq2qSVsCgaHenoD1HXgB9vzc07g10/p9p9yMayY1wotay5aTzFrjKTNm8
+fHwKpiI2exyisk8122bZ2dxG6HmBLkSld5/hs/4b8pnzBoDMYkp7MW9eg1a
M8YeepHgah3QpUuxtYSGzYo7r3Kx8BDZf/ag8d9/VMTUQrNQpGkc6hQja4Up
9dgzzlseFQ8lUJA8CjrPaCTWQKn6ZSNNqT1rvM56au7ZW8lVtYfuPJwOpiYt
GplsSD0UiUB6Jt7YgFHqGM+Nhp+srIoin3C9vkD6Da5gdLi8f9BXFsLF7aae
P2cwBNm7MciT1DS8qbPyN7Zk58naNLYEnuc7TnrFfpMi/AXkbm8oEvIk8F6K
ygxukOg+ytg0wxpDAnGQh7pDd0olka3cSuvUo7rBeTlL1rvZSE0q3TW/ax6l
wsOQW5EdYppmqtUt91iSAdgAVAOHHYpYPp5HqVP/I8tcOWPNPHXs+SViN+Hk
o3R93U4mlefL7reLFrR8nAmG75knhet8NsPjgeQEtsFYpYBPKD0GcXQkYrLY
Mo7ay+ViQ6v1pIZIWbrJYMYCwSZk24kan1KGfvqMsRQi7li1gJusrwCaikGc
Zo0SYRcVQvktV7wAPp+/SzeouadfWua9ks4rFcyY+tdlK9sar/WJAMPkgEh6
vyuSgDZ/1MXiovm56A06ponXNjXwVKlXJd6dLahDOQCZ+q1q0s/1EXCpig7A
79/cG3kdQqGv3vUGfY/Kxnwh2d8hLoUw8gYP1y3hdRs5o+YQb50JDXOo/mKc
5XChV3OqbpuWxz2zQxkDz+t2uBwQwUIV98IGMnhFWRPKzxivHcrgvUo9Wdw3
RIf5HJ43+3yLVTNApe2cefpBwXSHmGeDcsImOAvfpOSaOQsbVuX36S3a5x6R
5//lMuq+1pA5R1BhVm2t6PTMlF8NWfo0hj9pKhG+YE4gtwoTSz5hp5C0HaKF
WXIdTc+Rbd0VQ15NaCUXIng/9RAekXhEo2qDvLsgPWiTM/Rnvk0VECjbcOjZ
/So1AMiIVa3llDaG0muqZALoZKfq1iG+bZgDuoMBbKw7XcASXuyEQQ6jDd9g
i7Rv0atCACYb4bp870MCY1aY27Xayc7TfKhLDWED5k5bBNbuT1pKJmio5m+f
I4KTqaFTOF4qeJ+AEfn6OgGTNltd5/yuxtgIYq+LIw3duA0BwcnMQisA7kTa
UXoM7ySVwS/NqjakVE/zwPtZhXrO7etuE5cq+UHarAI/ZPkQTozJ1z1ftp5D
hOUpNSxuKuFC1JJXRmKiRFoTQV/RC6WQvNd/YqlkSeOe0NrNZ1gtA2zr9aOy
ykqN/iMVQsl4HIAf35rXTtgw7AfrKZu/dVAYzM6eHzjk9c4aYxqm1JMf/EZm
ADQ7aFn/yyPsZ8uRF+SkiW5VVYm1XRgZwm6asntawhWJ+srxPiGrhxMqXcw+
db9ZB44tfkQdkS8DqmOGBu6Wrhwcyqy8d4jodxK1tyiRlYhNwA2xOuAlFROl
tudGRlt2QOmeNfKZzFoKIbVIkiL0ObTnY6078NYFDVtSY5rMlTIRyPuGrtd3
ofyD2Q246SbK56HaP3qPKSHzsr7m9Gw9uyCOKBPWD9yatVieI4sJjbMAC5rb
zrjP7dxygbm88B5bfduuFaYHAJ3V25JnER83Qlld/+81AciD/J5xbm6bSV8H
S+oXONpbFilqsKkpnXLJHWA2A6oexVxGUWvYEp+fU75twqA6JndCA2OjM+mV
XqXqrp9k0uuCubJ/irY0ps2jKzhaOBSQcUcKiawogq1lywnt/yRhL0vCOROU
dLV5nJBtTHXIGe9jf5qAxj9uYJcbTOoVeP8gJK4bKXCuuO3Fy7FOvWe081FO
TLsMx4ndcAfY3cwiJqaFfoopLxdnBK+CyEqQYI775XxcvPhChsdDb+4rmMy0
XE7PN15lQ3erfiLXRiSHv7of+9fDihCXN8CPrFJNLGq4OMZVUv1JP+9Ize68
f/BG+AR+YfKpxq59l5z1u0rb2VBJVB9LzYLFUatFhYmTpucQzXN68yTZ0/X+
ZdYUJzYGIuiGTrTsOWTpcBoi0Sanma/stQEV9ld7wHsncrqQw9ve+RS7+1Xf
Thn/06rCwIcl5MbMvQBT0t7/SUYDA+hoheT+afAHQGWn0vcCPW/x8KMZ5usl
5PJTXBwIjFrA3LpVWAyWC0FgYu25JmYIOqOSIRCCmHGJslpHe+BOxE0Z74Ni
MA4WY/G/hexyxCCgqHZOYa1Ck7t2cjHUfKTONUmp1SO/Es0/q3duv4XaR4kT
6oUaTGdFBk0l1aPXvA58z2XZqSPrAJoJXOcksxhkI7T6peGkGsoPghTfn7fI
m0q02mFxtsIE2Q0bTg/lHCvp6Ev9U5c8ENr2gQlbAuueyCZfUoTaF7oQFhb9
M72t1ynir1vAPiZaJMpgk/urIwk9QkRK9/CkG568AjcVDJhBvafVTl1je6ex
+GUaIH+1efb+1RQVwkTtMSyIraYkqjJtIoFGX6bAZPKtkIEbQ5dx9/NJ2t+9
3Dl9sSVggM7Wol84F7nVQj7WoD0FfhcquNa5IweNxjXXXKwICMeJt3ZKD6V9
A+Z3sXxFbznqYlOI5BZFNPScL5yAiT4oobPy91gYVHfjVrZpvqckxW+Wtj4a
JSF4BoWVbWCrcrafNAPvwyEjlfYGwVQHC2oXbHGVpn/E9Ijpo+zt4H09/YLr
o5lu+lJ7Dos1vXgkqd00Mr9dl7ohG1a1VyRyFgvj1duYm8thMYunI7umZI1H
vSxQss5vdsZD/6AQVGWhrnCVruIcF8MJ/DCT9dBPb8sIrXtanqaHgG2TATkv
zLZX2BjTF5bQP8Pd3Zu7HfxuYL7HJf8Uw8wU07EEc/Q72RpgPb6J7f2KmW4R
+PNp7SDTn9uEYz455KXxf5JCrLP8M4yVvcoRIGKFSujJiwOFaFFuRbhIVv1V
nNH5BFXJBTZp1n24ioU1l39P68Y+AHCsHpHFkiSBngqn15Z3gqlvbtLKpjI4
+4LfQciOMtj6MO1nU0SMU+SxfHn13hCfCuiBwa/ljn28VB0pO/bZ9APOwMaa
P/cavq02PsZDyAREujfA4FG0LFf7SoOTcc9D/TEmtKYavdbIJNItWRQVg9M9
99QolwIszoS1I/mK0vMI27vREmIECNR9MdJF7Rc+hoVPMlku75eOVnRpbBDC
7gYQAC+OdAllAV6KEeDttNYQ0YNK2B7k5UI9VCM7Cuknu3q9nuMO7gQnyasY
tx/+LPTliRBwWtIztY30u4M0WhnB/GoeqlrmhMe1QBC5uE3tP9t0Ob8pIc1l
4uX3HgMuRRve5xY7y4ASXNYwkqsoZRjxGTPGUv+Z1J96qx7ude3I9SHri+zN
lxlj7ctvQAvRhOzn2gmTipRQPcy3Q04aSsqvPVz76K3mFS5wL7WLZx/NeUyU
Unr4psZFRJcJ6rJNdedfcVMsNGwqcu5m/olBtwcoNo/nlYUqugJecPHlivU3
opITSQs9e8SayreBm57mVU8TltGNyPUHTac7032pnsOmntKG7xPhpBNNDnw3
ZWe223sHPNoG9SHOOPOUqDZwTFazKZI5BtaD6Y/2DG0ScDRH6idHiNZ4J1rr
F4BISHrjRwvpDyYm1TCUV6kWob2zXpmEnGmNh3oxfx5uRFXK9BY8IO1lhQZG
+MvDUZaSXtJw7ZEO6bAdOXa9gmE0YR1PMMxSbVr0Y6OjU1SyAP4ewHrJRwib
xVMQL41Ox/p5xSetbZdaUrFPLYehFvZ0BpUJgnDRLDnIykCBYUMqcE0PCKC2
IMzzQAx8RHWtj3flX8hTgEThuxjZHhbifRHb79c2kByfU/a/UpCzKIqVAi4I
QNCiZWb6XbiibEIBbyhkcDmozzEvXd+GN1nGV+p91O4U+RoWlNgm76BJH8D8
cG2kGnjK5HpLnnOwM++1j3byTavZYp6Pmm1fCZ3/Ca9iKCD9Tjsxg9bjRiob
wbv37Z8+4PP4ykZVCC6CczYyB/RF3NAyXup4psdgyz+kBFrpYtyL/yDaPg7m
S/hjs15t8jR5tpYSz6li5s/9OUVwkFrCRukhc6DGKY4SYS8QUSkg5bqXTMR7
ysP08oXEQ6XM3rafbNXgcjl8+Va7/A93WfAKVBPUjWk7VZbaaOQxleLIMFMI
VluQV2VKTnPesSYxErmk2fEP8C3KvFqQh/GJFNvfw+8wAdvXCfs3xcPOsXfd
rB89zPtE9RbaJD3kHFJ4FUvTRhiDGx2fUq2D7NoDIxr2dU6OuepH/ctqCDBH
DarglidkPz/tk+rPLJ+eeZ4YuwKOqalIwZgpI3n+osvuZ0Te3rzk2mvIT9Hk
qJD8M2ZByXLJZset9wzZ6x1ZKxydFZZcZ1KAVzwcg+dA9s3TMD6D2ydwjklL
l1lJUhmgf74Q0UIQfLxR9uwxQEr4rTGDK+sRyMO5mN03tJhCLZiMdIi3C7pZ
hvym5JGkDUECYCNaFnKholOL+OpthIm+e51/HUWTH+0KufJIOhP/TjAFfnfU
ECV65M+JCe2A+O+AY4E1bmL1WXDoKlu33OK9bhAjPYkXIcNnk5JA7XJfwFCB
x5eYvgZHgPdxaXs4WcyByNNDr5eThrzIeMMdRVVJ3yDWDcO2ZuFVRMxWh7Pv
KpVtV+b6lfdpVp46WG4uqwt/Aj96cBqN+O/peYJurj/yx77Td3E8lZyBICgN
cINiaVAn2/6gmV5TA4FsGL7uR60pJsOKtAhSJHYYSd1E2RHMEPyn4x9hkHU+
9i8A7ckVx9b5bKhdD0cmjE+00/IKH/mJf4wx20ef0Q9nD7p8opg/oTxabJxJ
7/PWUTvg0SW2duvTWtwScsw9HKvOTz0kD4PdQfL0R8CMSomTVvDahHxmyyqt
Fd8VRfgOqU3SwZeAwcGWLY0DzhUc2r6/V16h5GVsL0X4b+As5uMRC3fbH4MZ
+gB+hyROjAC+WbvLpMgvnOHDEG+Tm8MEU1bZE9h235QtE78Z0Arcn9azQN31
ZGqo9uwaKzJl03aH0iGqfmn6f9EOfoPko/r1zePtxLKQ0Y6OOeYeWqLnhXhx
lNDyD/2z78iBm0itDSIqpTHYjRerbMbNE2sceeB6bFrMi/PPl2w84PcPuZd9
OeIOss1ZO8QZT6AV1REzOHlT4y1R+V/MkG30DLOk78sJQ9fOt0jHXHL+Kgu/
zv+KDV554b1XoqDTEN8ZlzFYCEEy+xLV3zT7DqgzfKDG+IaLSiIy/hvg3lAe
w0EaUrNvNe9qnrX+1yjZzeFgBGaE90mL2eHVlnBd47/cqNnUlgDomN+Wf/KW
6deLpE82M+3s2j54A8ApjR1eJib9878qw3eP+eQQqOKmHbBxw4BnhTQbO6YO
LIU1lq4NYuGKuKEBSRnMImsPuuFve6imdW8GGL3n5I0sxpe8ud4R/ATObqO1
7Dbf0RbfImP0jX6BcSRjR7VVLMdEtuXf/CAwwm5WKe1gwh0jgQVkOmTu/Vwc
Cwbk8eXEfcu8oJydnU2pXPSyRYq/xnXAQMroPXdWz71LdHLxB9UCAdPBgmET
syHrjM5l7hiRGZzc9UEYc2/WaBBRtCQdRJQU4mXjYZCEm3ij/Wq/2gTkJiSB
Nj3IXv8l3PkdfYgmX/g21bVi7N4P7g2xh/KF7FJUbqhHtJqiFhVKyFzTt+ww
9hQcilLI+3Nlc3uhwfFi82pc70zcYQG2Vo0bVy0sDslMxOqqhl08qCrSrQPM
akKGj1dsDeOLw2QmXbSSHTV+8FxVGBhEqchib4ZjaU8Ak/OvbqIvAIqJDMYU
W3XSHmnyYZ8U39wsh2aeoCb27WOnCDGUTAHeeMm9lZb+B+QkGk8RgPmtfhkp
p6UdkGcWm+tlSrSim8p+rZ0Ow0ZDVpW4r9kiagI3vLByR7Jx8p9FNv5M2C6S
2XhW82mrwWUhu7xhYAaVIQXwlnvzLM01ZslDCUQ/dtkWWt3lS5L/UqtlVMs9
IrbMbFJei0Gl+DW00UtGK5bFOQM8esL9mmIix3UMvLEZaQDmfp8Q+KSFis0F
HmVQ2iML2Qr9q6PTeU0+YM/o/6aPuadT66dolYoaDj+0TREObvoeVeh5BP1j
RldWV5au8gca5JtbltPgx8ELJDjFrC0R19uoIxzE+KnJIqAU1lrIivQdepyo
c0mZBZdasJyCwkOuv5RQNIZrPgKjIxxQBHDzpROBRD0weFjqEk11Q1nYrGzj
TkM/p2LMLNc1rfWQhuMSL8y5LsTD0zuP3r4GK7WS8vI2L7GJ/VD9TgDMvxik
2/lGOkh3QHu+9+tvrRr3ZIW0qhfc6CDbAbN9tD3nCqetUlo2Xe+Buq9L9quZ
svYtrfzzPYXEYtkkWDJaoNJseS1I7C93YBeEy692Zkk+0Z4i+ZzVbi/NLIwd
f4v0UdPV/3ksIubfSMa/NIcETx1/HSwn53zXrl5fD2Q+Z5MQBrokv0jbq7Mg
Jmt85oyQapdt5FIvcOAfzbTWhw0oBA1Z9rRRGxw9ZdneZNuOqrMWvY1MpsKA
Y5L9I/pAYBg/jZ1Pj3+WMvc0otkwgwQ5DGjYZFNAfdY+6Xd/wGac/WBDVFyZ
Xr4PCmmds65+MKonivLjcf9Ce73PLDNkn0wPPmRzwaxRYU/0lUruNsUjBtB+
1MJRnmSI1vfi8Anmf8dqCTiFqo/TFwhCssF838tFEPR8rvsafQIFP8kKOVrn
ECioovuh6vPJqcYdm1kXsBk5QgmcbFnmQ9QukazHLh5UeItVz/y2QEehVoxL
JtJPTxEInWcaZ05X+tssCpMsn8r3CAxlc+oHkAcPGRwV73SwaEn2EwraqIXE
Hg4DLG43kALfM+hwkrED2QuIsDoMOFX1mv1X3L3jtv68n+EMXVvt5q98fcwM
ogy7IAhLfR65lA4Dit+MJbLKWhrbJjZnvNFemah4p9N+HJq3OiKpFtQ1ii6I
srREz9XWfCBw6LgJFumUMW3XWDdMa92sqUKcZT2XWUKXFVdsMWkpfelBR6sI
WsoFEI5osRZd7nFKLq5LLsN1rM3VLzsZNP9La5M6nzOm/gJd1c9lj+2B0rmU
mQivjKOOzyBQ+JfIMfE6erbA0Nf3NVrkSexJjdc4yBx8iI07bPRjgGuUfcWv
SPOjRsD4dwVW4cgKjfle7EE8A9XpZiBrsvhrOlPSW480a0RvJRrvgtoRZrK8
r6/R5RKgA+STX36Te70VzDQfAMgNVXE/gufuOJ26KLNt5e23/vLLQaUfmIKL
yQLeFfWzHk2+8Q+d/oX2gR7Cutc+hha7lXtaOnpOdpeUZZO1qVelSrEAHjGo
jpmq3f8o78dPLLCTdTlAtRRHA3dx9vVxnVn0Wt4eXrQL8kV50Wyti8BkbSEc
/YQoLPGhFaRLjUlw1cwHo/SK+EvA4oWZFdWF/3LWZtDyD+uXXxMva1qKENgE
PuW4cZ6SfCpIgxDEe9VBaeTS4kzhGhJLrdJbi34RCM4cjky+7MePfdcxFBPo
ZUgD50RusYHFcKQoTbifuumHByhQfTkelTveeG1LaZ0ZhE/4zYvwQmYpAX7W
dDqzd0RYf0wHZCIQZgD9bX+0iCE/fe+tx3f60n99SXaCWnB7/w4/aaIR5Mdn
yURmsvdU6gXF35jM9h3RXW31pGFtQsi8FmFsVL1F0/REoFencsx0pT2eDv8l
qpoE8KPMqXZmtL3Xxe2VqnBQToTEPDbnPwMyP8v5BmPCpGf/AfSgSnyBTWfe
fsVp4PRpQjgttJuymRTXuXL1RXet2XVEGA6EF8N8B/DLQg5ShtVUq4HVZhKh
vp0ByRD89xLLOgt1QNAGbIzvDL0C/oQtZz09D62UPFXi0oi/6O1JRtrUtL9C
3UiUcrNrPCvrlYHcv1xfokPjB4Ot6K+JOq+pkqRCbNpt7EDouP7+w1XdZbiM
FZ6nofKcd1+h2tGfV1BgvVSjPJ82IhalBwjIud75aJb7Ua6WBbd2JKupvVSf
ZKdomSZnxYBoIGiWgLJu/bm4Xqrkzb9ILjdLN9JpP2AQX07h3kdCguglKAAD
l6SSCjaEOk6WmtuyRCqG0+OXuiSxghcjcJpfad1sRjW1g+rnZUNNRWl5qxxG
qvFG8t6PSm0S8MGAJGp1cMhzxW5C6+ADUF2V2HDBL0WlJmeX9aH1XbSDT9JZ
/tNGbTAPV9qoJIOmSTTOYx6D+U/p1//zh9rx0Nug2onq8SZCuLVoYS2OeVKy
yHHdCy8MKjh0Et7PzvIVZOsZRxPngy1YxRD0nQFj7GrEKrTE0VFTT1wV/8kI
jelmztAP/yfByXNzlOaWXyjl6t12Sf5E/cxhssFCb0okc3ETH4qYTF13Bs99
g3YDVWP0Op/Y51syR2+kg99Byuucjvj3UjKB/xt5wsnLb4MGa2n14UQn5EHX
iGfq9c1/ThWHiFJIWVCIY2rvoaPHkg2/T5TnaujxN6dJe/8dXwl32SRKJ1LP
bEwXHmnV6839LbMuifUp5ZGfEOvb5PnJqipy6qEPE4INDi0NJd9132O+hRzP
Pvr37mkTCbYArX5cMkfD9r4ZQ1/JJhODgM1xQHzEICSMm43+tmIP8q+WhR0y
0S6B+mDa5ZzhyCGNjwNSJy4FjYcbpgNO9TO0Qq83iN5xVOzAoyzc88TqBmoh
H1KaFHUjTiz/zWw5SjA6zZiRvwv0OItziHYxkJuVXBd2ZZ+R1+ApNDQQZLwl
PrOxCn0HDaM3oW8Hw3+LPtXsoXKJwOWKgZeHxa522dLRedN2etwYNT1ug+yr
jUnK9FARpMiHd2VzLpNbde2yV/uoDGjwUl80/IE2jlgPsu4N6iKXUqjiICQD
fBCXG/inmX2mLwfXEN6MZBlG5obTFol7EzE5neB2041hLJ1ZjW/JNai+BjKp
2xugl2YZUx5dzJyUwBcjwUU9d9I3mqFG3iATwq/umdUIKH4Y9YQRWENjFDV+
O8x76/U/98nNhvZpZx1K8dRZx9n+5T+PuUJye+E6QZacl0tqUestCNK3Lkb5
1JDqkiGVBqbat5mBrKm7/NuqoW99GdvhMyp9irAxB3qcSvnNMjnWFYPFmCTv
RXLYQNfhrhpC7e/KI7jiLyKdvjTfTZkFKlCgXH8bCWwdTpTuEiN3O+b3UOpM
GWIKVZ6ZvVP7CdszN1OKPIi4ZwMcsGeWerL9gj/lCujiMdKL5YNeVd59W3A5
BW1uW70+hE+ZbaVRLIJX+b02gKaS+UTBIZTuQks1r1CiZ1MZ/xkPX1HYhRk3
r6oXslc+jK0PByJiRImPrFglgG0lkKE3+eC5xHtkoEnOq2nxf5rhfUWbOipH
pAES8vEQoOgvdcZiWRqqhQZIN40CpXCtlEX7KPrINHSiuuQ8+685xQCHcn7P
neQUnDDnXdcie1fte48dT4c/h9AEELAZHC9cbnClB5h/DLiPeElTWn0L1Sqd
gZkCOnpvW/Nvilaq9nRwtsD+tBuNQL9mu5Nr1b+/GFjfLkH/ruurMnrpDbAY
DQv659L1jikCDtQCNp6R57TFI2w5r7104no3ylcRphOEdTp2hiCzSZPo8Vqo
I+iVzQZRg8yFtBYDOqvOT8heOSasgXHjFAsV0GkbLWbBpNxoi3Jpr/wtCMTX
NpE9vGIprrmbrWSB2cyFFDjvpI7XukqJhgovRGjZ8NvDp+p9I8QQJPUZUhsF
FiiQoxEFNJ37aiSUmpysD1bxYHa1NXr+hKS6abiYyvuI2LNy6xEsrMW7qztn
6NxBB93w9+LLBFqF9GIyV2kRxpg/YuOJ5S8uuCIHYWz+RxpDW2HFo/yAe6rC
xqVZLiLs95S9F5sN3a4hHFwcN8eAlg7jIWQ8nCyO3FIf5kpjb+c/QR1RFArD
7RMzTqibIqtCnRGLQnCsnx7tG3eFPSb7jIYdva5lS+1pEOSYCvly8qHoM88u
uPLFs+f1ZfqPcGHyknJkdbvsB7qe6Jm+XvL5Swxnm8Yj/k3mz1s0De6d+1XA
S/M68UwBL/pS7lecb+xNyVd8P+FAbYLQaKD+ANkWqfe6BwAAI4nb49I2boi/
+Pdbe+rROENsxvSY8Z50EqCiEhaMCfGcwlBrNmNVuqho7LH8QF5c0F3i5yr7
CSf1fp5rxK2iR+WVtD2+Nmfyoud390mstmpg8LCEOhSNdPJO41kWcOdygYFk
SKF6sxKwZemw3SICCB/IBWdYsFgjhGPfuDcxKKsdDkrMAiJZkXrWurws4VXZ
DWT45N6U35zlX0rsKXjUULyLdp8ZYhzDPv89IUa1PgnzYQnGbFNtb6hAoopT
+bAkOa/gsfmysPTduK5YJmTe99M+GZhfpgjQXHSP3iGM1lYILCbD3HM8hiFm
zhDV3S7MieklQbQHpSKgYTw1EmI6gIqrMEPWeJK9IUGPNUaEmP9qPBv3MgwG
NetZOhS5OIsB7Um2emQ8fRqIGAHO26Unz3+4tCDpx5yoSKldLliftnhRtMvM
VFY0SsMysGrylNoJ613wHBDgnkkB1JNVsmXBRnQfsn+mcxUCXwifcUX/I8dY
Y+I3BKSk79bVVkJXTiJ4GVVJxXAF5dXJm2rjFuHRtn9OAs58UTzfULiUHBuR
KSL0Mqsa9javLYeGiauYpte8CpjaNVAzGTbSp4cjdLSX/21AW1k7HJzYXqMh
eJNgP7HxiylFn54CCfB4D54zlO5m6646Xqg4zHku25qBWiXMemwobj6NvUfq
KFrhEvBfsu9+WP3GDiBWZzvsiGU8Ouewr5ukE95MPdNma+A/mAwHv3zrVbwH
Qt01kLgu3pMafX+t/8X7ArdEvmVzGqaTaNE6iBwrc0yMkKyiTsRzGi6VQuxc
w8ERE8hw9A2pjg75gyvSlRU71+uBQ4YU/wxitGcr8DLucBSwGjbOJ39v8PgC
k1DgTLL5RTZmntbThCBykGUBSQCpCiLOl4NdqvELrtSU3yRvA7QwoQq8oz9F
4J2Bugdo4GLPORifyehu41wJC8DxVORX4HT34fcEypt/6+GttzJ+LnkN3NsL
z/W25NxZ4wxYcHCFjnnhK62xunkvNHjTnxpoXdKFhsE4X8KUvnJQh6UvSI+b
N2BdASSZVXzApgjtjSuiltaYH8RBCvMwjsQsvuV/EO7Rq1xpifMMHePvf3qH
3s4CnNqt3uQMVTwMtKMAAaHzJ2qe/gRqLbwuivilzrNmK3B1S05NJgl9jwSB
3/LPYSLV+spQ6ZCfxNzeS3bleUgYDMiUDuoVsToTexkSYo8h8NXzTsJZ3VNI
2vQ7n6QqABg4ypqbhuoWyW1WVWcbDOG9qtmAdY0qmlWRRGFkCB8bu9Ozm7CB
i9oGxsifDuvpfM7hRP2QVAe4uZKCXxC/xqsYAAOBfPkLNavB+p1aQHq5gSQi
VhX/3jIbyzDIw2KkJ2L0DWrNmp8yDGLjSVkhIEzbrProXfF33e5z2GX6r7hU
vKq8RLVcEmHSPMOwxdUy66FURPa2P0hj3eJQ7D2Ek9tqnfe1ndIjG66T19Jy
qoAe8WwcEMOMIZ5Lis82w83K9bAJS1fsx0abWQ7cXkBUblkbvcuZ4IeKf9J7
tztZdAlgYYQyHlHAeOchAUJOwuXWfu4ADHYYJ+3oJB586lflLTmAeFMVPLzy
zSu4uP5V5FcNJjmvN4AtLuN+AbeC7nZzpFonbRPQkw6SjVJzTDRede8BRb59
+/Es5W0SfHaHhfAUbgagc4FVYUurNRTH09VEpizk3yKlxGWNiykHujcI5kzQ
Ob6QzmC9JwNQjRW4iUyb7oVSn3I9bLESbW+LUJV7WSXQblfPgLxnyGUScDnD
8RL5Zc/swk1VmZFiE1BHtvFBNH8XYy9SucNNrrXHSQLZ2nbaqt2XqYVcsYT2
uCt43nHCdbRjM4kzKwVg9CINbg8YXa/DBr+ZPlEzCu1aLeP08iJmKt5x7hq8
TauP1bpMkozTjRgYvKYj5ri0WW34lraFYMeFD9OfNr/dyXNCvFrxYB9dketw
KMKEKwJfcHgMKOsFWRlMAX48u1pgQhqGHLDXdiYd8zKW4vNsq4cnkSyHrLuK
/w6bhfmnIxQLZzdHPnYlKYPfwMQj9wRHtTKvvcHSnLoRV7c924gKb1N/cAEW
XbVqZvubWehWVfiMeX8FrZTrFYpaelSWE7PZdV/89BF6m0EF9goygWK9BK7c
9MJ9eSIdwrxtFYvM6MsVagWHKfElyEp89h/VqZu1iO15Jh6dxd3u4RNMdx4I
aY7mXcKESw4yBdI+mjRotk1/PK0Kmq/zKeVx8wA8wQK/YGP9oAPnR/5NJrqu
LfoC3d9Np4c8FZ7SkRB6uDppmCxjif3OeXsmfyMsUWXGdxEz8FwpRSyPCyIu
BPXkKYQ5N/0ZJvSZYTtMoKGIfyWmcu7L2+OWmdZGnRIa2114R8lgimxkFtvZ
7qWvSy/ZShVzvhXpCUsPXlaoX4Kf6Z6dWClh/JKa96L/8qXz8QwE19EiGyso
vOzBS2UFlNSyQEkfTxn3E2PJ6rM2rphVSBTT6jYCRIyErmsL8+dLf1zigJxH
FkDN9+BjK6BXF78aZG+nZY3BVMiMY+9fZDWM6LKAqbcg0owdjl4QoyMvUUtu
NQrDaGIs7e9WAHm70+HLOxb8GoEltGO46saezboRDPFeXwgOWETXsrtJVOkb
dcVOkZLh1IFDS8QlNZEb55LO6P1snAmUtJ46CSzShuxTW761R7Mf2Mxa76XQ
C2cI+04mJgJpK57lc38vAm8OtO3UL91Ds6dN9zuC+sm1gOO3jq/IbGtoSM+C
QQGELXj+nphuqoCaZ/fPvbSjes4lRBn2FSiWG2lXQO0S2ifUOX90UNkhu+DK
67l9PAaYLNpgxJDiEb/RT0ptY/r0N3k9fYlCYSFvPy7yRWJWk6ZvC7WOyAz8
0kLfXVJAZlrG0VE88wviacS+rOQkrYSLgUIhF0Uww7mq+L0aqhywMY30EzBG
D8Bf9fGFvhLTU4C06b5kIPYOjwO3o3/D9mduqKGGY+ICgRw1tDVbL8b76sbi
VPrKKxDS8Dxr4wTmV0FRjmy8iPXATPGt0MS7Lm9QuddzgzxDcyENk0dZz6LA
9bGAtVB8+DBkDiZvia4CFnUMwSm6Kl0q9RIovVJhuhFoPrxaR+o0Qg0PeSe3
63EJrFcf0XHIxMpeSUKkeLadey3mxWVfzJeDPN+f+1VeEVLtxD+wshrmCEEo
ZbKJki+Pa7Qo1329vjar6rkE7RRePTZrrT3S9pOVtwcH25LqZ4Rqm5jEGSQ+
o7uK5cYfed5TNebyhKb25Nhw3xEwlTHRUpFiIDJQynDVz8zGn0XIftcN3hQo
6B8C8NtiBxniV38UI6BtWMG35uniIClvQrcOEGZJEhq2pCYVctR3EpUDSk2s
r3lrq4v01FgXdZgmdXDUixpTxn1uH6ar10cH0crwT+V1qdY9Lyz3Vld5Afd8
sieaOUmzNNbPl4oD9URFIHaZ0ig7IrxduibyPHPiVVOBCbvlTyl4BR/iU6Fr
nKWPCqG99aaLEVdr/zOdH/HCZ70dJ4BLJ+65faKQBJZQdK0QdoA2/nfF27lJ
tznnqixNIKc8KMCHQFsjnZmirw9McIJPT64P6+Rq5fvXVjhyNqLNh+VuNKyd
8xkWVeCP7GsT88UuFM6+TYutIgXC2Xbb/GKPa6EWtlBtuWqMqaWg8PMa9Gwu
Ayobe0nLspIwpEY5cR9Sbm3hqkwaeJUiLY+xElLLXHWrPjhYS8gZ+qOHXB+Z
7jJOv9flnytwbif83n66b86OO5bRjal8M+/CCC3Nypyq3IowJkzaPcHqIU9j
WIKuY8fZvkwqA/xX8DgAkvz7W9DLszDKKgu5h5woviKky1BMbkrwKpl8GXqJ
sxyPIJLYwszHH8n4bfbEOKCptvux8UytUSqgXeP3h2nF9vAoCkS486MlTDLM
p4AEp9oPHgRawzVWAOArELuoClhA12MlENqHICKyx7mTMETGTpBJb/090hMm
X7QakteLCaAha+03pNppMEZXavCe3YzlIRQvu2jl8sybdNuOvN/XYaJsUVc1
QxKym7qvCkNWTtf6qaQCL1Lm7PIIdtsJJNyfyE5vW2hgdMLWGSJWhJnzxxMg
t2y2Lqvr0CwiQ2c5JRcppcN7HKf1rvqkjXLx6JxtwUrcvATuV4OEda4qXzZc
QcGyTZGehleBVgVeC20omEhMY2D1aA64XE0AKM9CI7fz7YWluA25qtOtstwh
6Y/YF4QDN2ov4qkBjuh9xLHLitEkJt7xeEYGpQjXMwGsi0sy8vAqwpO5bJNP
9aDkZ+6Yuz9e4kbT0Fa5fDULGH8C89ObeAZsyY3u/IJwihOoqGtewoh96JzR
jbqO+hwsk8sWYy8FEFWWhwzmF9Qrs3nVOn/BnEXIsknM+3DpF7LLxBNRQd4k
FFNP3D8UX1k2SdsXq7M8xt1VP25Cx9hLcwZ5cXh6bMJF5Lzp+/hz/2stz7qr
CvlqJ/PKAMKJuIls8jvnHcE8shTk7SFlSHcvZaGtgmTBXWnU+9Hrmm4nQddE
8+wcBnT1zJ9fXLRz59WXIjZrJwDI6Ejn9pbczSajl6nOq/gIxyks45W28MEM
0RXKlyrW+hoexLBuoqGuaDoESY/jeNLeChKmvhnU0gvxSn8LENxD8ASnUwHB
1CgCZJrO17gbAt2FjcZ4SrFb+p4uiU55U8NdFxeYQt9uhNkpxxYZcN8X2IL3
JZIgafvL1cgrZx6lOK24iGh40a8uUmTDqIHLhBs8A3KTLZfWlPFDgpvD4vZJ
8DUiwqsDi84GtaHtyZwyUJZZ1q9iofWWuh1T32p2qdHamNXXCb2ZkcVBm624
DlJP49EpXVpWz0EXlR6W6BBDAMX5agpVg9eMDAzfQrgKVRcLj2TqaMB8Bxg1
B0qenHjEsd/BHmVZ1jgacaxe5yqWa63HDOEGMXxcii2/02+++s+dKAH8Xaa+
kmVQndUs5PqSHfE3vKm7puEs/NJ/cot72nmO9k9VWSN12dLyuFWCrGipkTTC
K45k3gRdrfzTU91Qky5ir0psDNba4NVGPG941MyESzkjO7JE+7ggW15nTw/c
GXZI8LUtvmKcrlEUhB4L4XYKhDAx7VNJZhoayzzZzJAc9udwUWOZHpEacgDE
vGPnhT7pNR/DUglfhcabm9BIxcMNPXGEYUHS8jZCpp9nnXBMmAqHwXC87/CX
YwcpfFpi4swx290H7/UBvhcE5joqI5E7ylx/lTXVinkG2X/Koq8XxRzwinA4
cR261BzoD8H3SMC585Y86Q+jAW8iBa9TldlUKMv+QT+RQu7b6UsrWNQPoXyl
ROeR7B9BbTHGuOxahJQ6Jom5bNdcd9btxAvdR3n3BIl50Hyzdt2yDzbzGRJh
HCmdqCjBNrq/sy02cwMmHT928BHMhkXv3onleDKW5CMMrM+4/RyO0vizkq8u
9900lpb5qQOgpxgMUbYgTojqoSClzvFn17TW6Teueroic3aXl2KS0xiLbkoy
BWbjcoKIaMw8MvBZ6FbUdQ3GMdSYrU81zO/OFozdHwvQB4kPuyeLVVgqW72z
pfwe2uixVNjQWaQH8mhjGJdwNa9RAFXnu3UIFWaT735X/3UIR+diZZcbnK3X
UBu2RKtQ95wFKsayP4iXG7ryUFXjzeQP0nKHyXzHzfyOyruCC5rk5flB9J5o
x8N3dnkN3ohcr+rLNwma2pqhmqjLjBnKpx4UQWK4tPF0eeLD60ehZV4WbKRS
ZwqSxZ20BCSxQ6QnSG7I5mHzpUuYYfKHCNAdryytEAeIJFyGisclUnlQXIrr
8CxtFAVdoyhoe8Oh2ISB7PKYcgd3jL3Q+MRhujs9+P4WOG7vjmMx+L+pgGbh
sLAVKDNEnreCVZYhsivJMvMQ/gG4OqhHZPWHSEaXV7ILrC/4MDIpCTHktC+8
yMK8kE4ij64R9uf5FLHcIj9DZfhq6+9NRDXNuiezsXG0YXvha/vUln12OeXq
2xKiI4kneQjij9TSepfRkv2V+nzAuPdAmEiA9VCIX1yoSTBjAX+QX7Yaq0Wr
BR3NWCPDnHb+REEqxUbZNvFVNZcqotjF64KHEFojpFqaiK/9gsQv+mP/ux58
ZmWK46T/YNJIyZG7Thj/6LGiDmXHOyL+JrHfZWdM/kfvHebC6Ym0e0YkRs+w
iZ4X1gYhf4cDQo3oJXfGgwgEA+wqTYciEenK9/QEsufUyAQUVHqnvcpainKR
oM5PQaSt35zhmIG8+oUoCU13iaIIcu4twtJr0W1eBU+Cp2gASHhlmZHHrtpI
mmzQeBlv8jf0AYdGPrAzU8mJLIy07o91sMs2iKOgL828LOv475E2WtBtAhsJ
CVhwJD2G4leQLbwEmvGpwCZPkCvjf4lzoLNubSIcEfGqnBC23I2UEOWSYhwg
uohu40gzEjrd/gujzU8fqTIJH/Tj+459NYR5WqrBVSvluSFptyJnYKeaQmVu
qpP1n4JQ4IsPYlqfd63uHp2GR8gq8zbKgRkyRmA8BsBUrE6l4dfGU+hn3Lvq
BMfzNLj/OEqZs1twW6L/f8URM0worDllX1fHsOIgPs6GfcXyhdJrwugTmgpq
UpaGsWwYODRY8urqPwDZeijNJiD9Bq5Q8wvz6FkTEHKboUh4Ou+2Je8nWFni
+tD6t/mnPDR55ssu0HWuQURPAQ+DxrAIYmR+a+SSg97lW5y4qBPzKykD41e2
1twbwTLtbk95OCMrvz4Q8NhZV5YcIgK/UwBjYahBAFXP4j8+81jPca8JHG+u
KrywmUm0RFdASYVpwksGtN4fOcZ67zE3X6yr/1US04YSKQDxWiaIsWAWcrmS
U7stzonwlRKnNA+tJbeEIZIOryFJqVhvCnw9OVEFNG1+klcQ/iIaCyejTw84
MfFKAHFOokPGSWVWrbOApCPnQjo3qo3Zfa0VtC84WRCMwjOUq1OPuWxoykRN
OF+auOQI34c52QB5zf8fvSKPfzKXS3L6optIQgwCKRMeL3vpuqU0U3LbpC2U
UdQq+Ea5UD3JNRG3UM6vOswDH3iSOapdoX6NhflZSy6H/WTDEosgUi3FALCW
vQIyw0JTp6zcdhvWaWUSjlmGcSLbm6n5Vrq6138rrJV2VJgX44qzMQSHA+CK
1FhA94+6Mc0eilQkvz8+5CQcuiZgecKsoc1pzXo9VjaS41VYMd+wbK5OZs/9
195KG3TlHfS/Lg6PxBK7dwS7MraJFPU6pqzK2ACWuIhNmmD+mezrla0Wlwdp
H02UvdEci1rQZyb2yA/PnsbfsQT8gEvZUTQzXe41d3z5sCO2wcxGPtjiP6Cj
SuKtmM4RqrYdkGaOlinZ9BQFOjlrCoiDdN+7P9UH+bUugG3wo8qn3CBoalLR
djhKmTrc1Wa736nAZD6LpzCl3FG61Teyq9K/rVKdnlt/Rce4b6vEH+7d8G05
kb/6od6CfT9lD/lV7ylG0SBl9PCT0xRJ1FSSp8KXq9F4I6o+5PhqukhjUlvn
+5TC5iRkH3DVSQbbN8ois5CovXB/4o210PMrM5LgjkQqRzhZYoIxua2PP2GI
Y55k68sAZR2dpLfbox5YWv4jnerFP/ajLWYM8VCGm8SuiiNdl+eXzAskPwGY
ipRUn27fe3JrmGuKeuuZw98HPtQrUvRApeNJcfxJc+xZOSMt+5V86o0f+wL+
LLHzEkrd7NSNACtku6EREKA/8zpQumMH52nBFMMfTZpq9LBnFZjvDky6kLwD
hABquPg+Ey/4gajYHuRzbrDyR0Y7kcN6fHmoe8funu0mvoc0vVONoXl3cPyf
NoGdZW2PZ9I59EvwSI743wTua7vp7ZveenHxHUdTLXJDsJvclkH+OGwyQmpf
XCNq7afFLEat5Zciqp0ulGR0ie3zbNHlxBmEzSp8LjSeckzJ/NODa0EkQNWQ
1CQU4ptLvJFE0si/UkCsFgzAfRez8wRFZi1js0ZoUicvJ2ZAOpaPPIloFe4T
gBbIfyGPxLE0nvdTAH9Guw4cOHc8cAgI3al+DR1J+wf/aVEjvE+Biip3/D7D
IvDb56h+Ql88geCMaqAro8+BNgyzRmZD5UrbvK8TaVKWWhyOadpjEPV0FxIm
w0CO2KArK/PlEor28vgiu7TI5O46c6C9usugBiL6Bs0ueX52lHc3o0JomhWj
Zd4p6q7BPvLS96XwEuTN7fBNw1QGiEnUDDnaJtfg3vUX7eBt3KE0Z/44V+qD
Vjp5yB4Hl5x6xaq9OwTxdXrQ/cwrVzB4C4LT46GMc1yBQwMY9xPCSvwlB8MH
n+IFjP6fKn9onniMSNJecqls80xbsT2/JX/X6h9jtsTS025WiESUqClJXgqw
cMeadhyKjI5YfjdCoOEy8sf39Qh4DS0Eyhf1Hs+ixkGNUWauxmCSU7iKQ2FS
zSQymH4LYJKL3ADr6ukj2MokGvYJ+gBV6peN89YqxyI4M76btqeVBKPJzjF1
91l3mPynTc6bJG8BSNyIae2C7Ej7Cc6TGQqx2gZ6HPpEZyJ+FRwDeCz8UFJT
O7QrDKCFKEvDLr2ItvBTU8JfuJ5K/8Jiw+vYbdlJ9Bvw8py55ZhKN/Z3l+YZ
Arbf7oWPYYQ/wNpH9Wd4qVnpw9dn5PDigyaP/RP/Oyc+OrwD9O0bwd6S6nlP
epDGtIEAauSmqppeUzAXjrixWppQBdJZCLmQ7jzycQYCF9Uf8X1L25K/QsPQ
aEVMZLLDZhcnQli8mYBzKqD87+090HysbDr7XtqmqWcFlmuvUOMKSWk/3e3J
4phEu0uc8d/MrEQ7kBX/yCmt7iLj5H5tfdt3w3N67loJrsPUSksnB2YBNexB
3PiCGncZ2A1FvtADsjsPsJjQrIEuHFtPlcrX7qQet2YE140AkWPLpDM89Jmo
JqAictrKMHXXiPDBwkL4U69faeaE/lhQpL6sKGTFWZPkn7DT99SK0kqP++r6
uW5Xr497hUmDzCjtGVuxByQJIY/4rd8HH5SRt6509fIpQ5yXjvAHILAAiDlv
kgv34eWDUGWcDBq+LDPqHLRXe+K8bWAjjhcm2KoThW4QshZsn4f89emlfX5F
0BGoWAezHradnkxl0e7EibuBlxG00lOYi3D4hgyp+AAYw2nrxPDlccplhUlS
VBluu6WJboT0wBpzPPUEH8N+/JbvYiC8pwFHlrQutHxE2FqMpHHfo4S/QKis
EOmrh2RrkjjyiqxDdXgKP21pIpLZx7IbtLKOqjywLurg7d7V7JhbDWkOZ8Bt
2iKGKd+Tn1Fv9M9W7gSY+/1eP2/A42/26/S17afCZFLfHO/Vf06s0CwvWcvv
xq3dt+j14Wky06grYNrHUv/KoUooHndkQ1DzZPbW18TbVWGIqAC4TpqJ6Pxj
VIoYaEION3Qzijjnf1n/Q01sHoe+eC7qlIie5kVZyz2hgv07BDA92Cxhi0Br
d+pFIxDaC/glx11irk3ZyDT4bdajYbsRO7HHjkgLHalYVpCpR8jiDyDqVzPQ
AYkbE+ve5+O5aKc0KUPfJw00dl4qm2fT4oR+pb81qgjQUxTwsV+CdCBXTz3a
9YCZm0VuBLT/K+O1GHft9NhUYVlUnaOCR2EVog5rKyKr7Nw3LaQ0/gd+WJ1M
RfNFvW0LqIAspExL6ECaL5LbiDrGK+hESLBR8QLfeMFIzG8VVImomZkwzK2p
tvX5p5mUBAlPnzUXb7JNCKEYfa5o7w4six78bNVV97S/k2InhR/HpudCOADl
ZE3PMglMa7LUYZzGfFYjmS8jG8Mg3aFMtbGV4uQhGu5u5++uRqLZB2YlLFXb
IN8I7FaopaV5+C7PYbNS0Cn0l5tflwHMw4RpCqLiE7LTfH1xk9Xkd0HQKeGP
kFd2FHh8OIsseaMCJY6i2Ee3wXcZRzhHGoqXTPoQJJ+Gahj+QJbfZg0r5QGN
4lVZoAxFtxa60PacqHFmC3vybqrwTweAXW6HK/zzM/ap5PELqHS6tdgZ6bT6
rJv1ORxWssSVpfPWq6O9lIRK+xSAN3eJ0LKlXFOrIPzlxq+zqxaQQPSkVWD3
lCA6dDCUghBszmt06SEEaLvUZXPxQcJTXk9O7mHMv3MdBpgUgZmHKKUavywN
toTSHbqjC5oXnyxL6oZVWeJVayEJ9Y/9NIIrN1e8OPKIQjBPS/uZX2jDV4Rz
XtHXDcy3/4pwih2M3YI+JGwn1Sc3yK1u6CWXhdHdmA4Cgo1827Sbzfp37Est
HxkWqNlrLGpLRQD//C2uFHXTHfOGZu65IDpDRMewWglO9JkbJEDhMzkd2FF+
dJsefdXLlt0BGxRVH/ufPivuZS/rW2b77afP1sCa7GeJt9GtDFdTv47Jp0yB
CIY5el3+SwT3J1BxURxN0NFnjo4KGTyCaCT1gm437E06od97iv0j+3HigVxm
cgXYUoFjxhv0CJGG0GSCfQ6EIq1LW51uqaaDsp+kdgsO7UWspSi2Y9ljw/1R
2ErgW+b4mcxx1kuDNhPqeJfhnMXF8WFnI/29Uu/yWzLXSbu68H2hq9qDshWy
HhkXtMGD4JFJInKJw2wmL5eSWJnrWXPR4D5Hdw6cjW+Xc9nv53zxvOWqN2HU
yEa0Z1rPrz/oAQeqaFQs3Ox2g+19Wy0zkpYtZMycCxvDw5dqJfqxM6gVcUKS
/Djk0X0157va/JuKCIvane71qpq0YbtWHrf7Lu/CUG8YSvyBMbjsFkfGlzIw
Ss160GHLOrsNz9H84Yr4sFBNM1HOfI6S6UTe1nPlDUlWWlI+UkK3LcfE3GoY
0HQjvLqysHnwZiAK1XDzTq2uAbxFCWpWEB3UNdUbhc2rq98+W7pOKftm4dyB
fkx7nmum5ZCuby0zMIoVmITzOaby/2vnWxTp9Lpiqo5JLCT5GzjRM2G5Hii3
ii9JZpewrLKXCk4IBnSrDVUULu0p1zpzgxI7IAEHQDD4zP7vENB5Q8i4oXLr
mDWKihtje8bLgahcGms/kuQI0IXu0zFrd605YHKaxoWm+nxZ3eHxNN1fyv+d
7fUdBz9+18MH0fy74K/oz6bPt6vjy8P3FpL7qnZs8JmLgcA4a/IEyEXnHiW4
fCRMeUPDq4c62yIK2sLIcwz1squ8raxcfOCxltLPhmdSo6LOOgb+SaTXdwn+
D91bI+zD8y1oV++Xks9hlK+aQ53Vwf8gGc6a+IGvXiIpNr8l5yM9TNb4mQJd
figEMrawJh7kax9+BcfLKuMbaEDIrA3Fa0jiKT6CVfpKAF90cYbKuNXFJLOB
0LcYrAD4SCj1DEQvZYMszJDrkvDKgp5+DfFUYxLPnuDtrf78ZVLCK8xF7CQ/
Q1u30y9y2FDM5NjhRbfRmYezSGZIJx7yE2tJsna6rthArT1iTkskXC34ifZG
GuMtMdVGynM6vgr7Gj02VQIfoDxmjCdp3IDI7L5bRSE4qlP7C/QOQ8NXKXfr
9ThXwEUheV1QfI+jb+/ExL5n69lM7egXuqSPfT4qM6MOtv9fzRa9tRGSRpbx
ifaPJE+2Qhkbms62W32UZvg73lP4ToxyathDjUae+nrqkkBkRZdL3R1vSevO
1wUgNS/PpUMDUz8ohrCx/1ieBmKd/XEi7cjzM4YPzcyRHMmgPtLsNX+6rjlt
NFvtTuIGZQJa/XMll1nPqoCBeKHjY9i0JQVJtby5c9k8Fq9d0xuBpe+4ceL/
TFz2dJElpmf0XYxVhN78j2cJVROMZsXYUfU/tSGgjstHWw79PrvAFVnrZfDZ
sCdHGS43D5NHfU7/1L8T6eJk5fe3gdknCgpKWvE5h0l8YwGKaJozzp+mIGUx
zvZtvBBKZQhPzhKnAaHv1P0Ik995QnMRYPhBgi/20dyp4pahQUnCtxgDZQ7U
E23p634H4FW/yveBYVHN0Y1JFj1kpK1m3NTvU+idPVJU9EbiyIJ2Q5+iAW/N
lqWRuIHzfCZpZhu//8Hg3hRELVnHPTFFYYp5qZDQRtwcR4+d0TpDTXpK7ZhZ
DTnxwXYp6tLlLMxnwGtNpVpslUgdTYMnCtp1hfBEhHS62K0ugKPVfOIkS5uM
+S/L4ouaLyFG4nE0ZiL0OSZcD3qf9XUCGGADWOq8jslMHlxeaTcAXT/aVedP
TyTTMrc+omxY2+Q5a8q9eA54SddYxyJWfGmQ+lPK5AoY6kItbyV/0YFh2gJd
iS4ZdbHukhoPXS2gpXvWuZFN9vvqsR6MIYvK0zyJfkVqxE+AvUgyAYszM2oo
4vmnIt59DK2KC1qq//4p0TgTuv227nI+097BVIvhMjZ2WKNPRHpn4qd0eXeM
GSuvYevtNHLwmDuYre56NuFcnnbdynZoFOk0uqn54lluM9yCVSi7/kkbnnEP
1x8z9BrCUAKFOsazeIvvVp6OamWisjEAZiqudj2036v9xgpKIzaij27Gh/qv
ntIh0AYbimaA6Elag99Mj55mYr8A536r3x6sdTKmEUStRMG9HJQTDPGm/Nsl
ArSvCH7XpctT8zEZxMpabnjtnFMlN2k3KWknVdaOgNwfJl97NsdPCoCi/P/d
enDZQjWaL89lrUsbQCf/Qen/o2iA3JYMHKHsy53qvyVItIVP1OBDPMVnpfDZ
zSTKtwEK38tqLDJAzW7sH435u295MC0kyyGnVdZzUPd3smZfcmcZh+nBV531
w9IBzR1iiHX7h7IgZfutB3TS0d58f2I8QRZAiHnCvTPDMuIdwA/Q/JmCjK++
VPf5k3F+ER+clJatjv38E4QoJfqK5euO0TzdBNCD6XaYtK6P7T5VLo70577W
P30BVKej16abA7Kc1iGlDm/tmL2mTRGUuxmptYhUw8+XFj4ywWNqW/czhTZX
UybroFOmZ0AOPbqU9whdiGMu7o743FPcD0viKYSnQa5ny/x9sqFWtvm5jj6g
c9wJWlZigCcOhrX7GjLE/OZ1nHkWslMTwD1eirgIgIkK1qOPVE0ebKHVFkqr
qq5elhPYzigtAyKWg6KsKv70OLeJHDTyhCW3hnYF2Jz5bFvSsWvpghoy7T9x
ubwW/lLeGZgCCkXHQkca7jFO1tWdfSxALz79x6m4CFG9qUkhYF0gDKbxvD9L
U4yrUnLDkG72yhMu6NSmuG5VWKyB+kfZMlK79Wzmb0f5icIuBivkFKGjNrjX
WiZcipT/0l4On5euqdtQiPK0TruUDBprSFwbg1SUnJ2fXcXqEyYQrW/ME3ER
Xaoy8IBNNNzxJbYrB+rBSxDqt4pkdqLumFVjby0gZcin9p8CuN4PUxHC/qC8
IZpqh5xvNeWyJ8+RFRL/iBF3t7++PB1vDYEW0ccY+rlx1sHsgOJSIeBJCZNb
MnKG0x0H6pCSfI/1Tjbhf06paAxTSHJs5ZYLf2bU2YdSG1uxP3Yfz/+7gikA
e2qE8QGnZeEJwVtTLECIziX6GdBBVKHpzxV6X1icfYZpWV41fbpSQwvt/1Va
itxuqIWtuyQ+oHCE98Kzz8q/Z7OMH64MvIm6xSfg+VfoK5dG/hnk0URBDpPY
j7vX003470sDeFqcNyWzzwLi9LMM8NOeOavh0Vh+v4HpHj9v/SZ00Bre90dc
N0Sia6LwsWaeLApEtXXmRWHWLmTeV5LMGuZ3U8hp95ZheevkbyniAhnu+nhx
hR0GWQWXjIxlQU1sR+grPciiNj5Gee7IwuDqQ+KvMf46IXunvcrOja3yriAN
aV197v9O+6r1295TSU87nrmUOaP7Xxaps3v1PDYphFq1+rzp40xTkNcr/B2I
im8bCluHuVtJweCxY8SI3BeVKxTM7a+H8Etfk87qa7P0OH+/9Zc6s7fvXVem
P9olhSorIRc6VEFSdTBk6JGQSi1FTCFmwy9SIMyGM+BgllxapwrP/pOyBZ37
KVtvs5s/A+BWPMZZ4G/eYrL5inNinI8Rk/c4AICmvynu9FyaOOZHM3ntayuV
3LNZhpK3yTAjxFYSdPCuIo2DHiuSoE8YZhZYW6sKqF5+ZRf63xwkE7c0EcaT
b7GlY8vwPVgAnIuM+oDhtjXOBj1Z322nAkJTMQPgRlpEgSEYO1sttuJuRCqG
rYpQbab4FnICsAx1rnW85Y4fxablxvUf/TN8ql4b/97/KCWzZVJTg8JAQggR
R1X944Lol7FZJ5EH82e9C0xKJB5dGQWmLQaEAL1crOTbvzKJ/dSNQklHhZJX
U81eq9rLwH5uUYA9W/JZv1uWR24jHm3WLFgqf4c4B9SKYdirg8ADRNgV87+N
76rS2cstAZuG5I7But3RcLf6HMuOOrnaIeQxs0TjEHNW7gDy3gPrevV6b9ou
fOPoqCHgoQ3njqjPV8fw72mlSN2oz5kase+Vy42cB1gVynMPfcjs4edjxIzV
EmTOG+BTBMRevKrzzAVL2FboJ2SPMf/Y8AZZe6bjSx5drnvAp4QsIAFjk5cc
LNXBkN2d8eJkndv2gS0WA87p+ol5QlXHY3OiH/EmaJwFycWd6yWp1eRV1M4i
vgHjhyvmuITn0ftRKUua1rdORBYtgvSrJNy7OV1PgC4v8OD3suwOtft3tbRb
eiBqcYULprGVvKFrKUq2O76ig9iYJ33Jcyv/6cy4SfzUshAipX+D1GjiwoEa
m2WUKP5XnkCX+MWslxW50qtUkB3YslziwPrFg9AHqzyX39eG3iG6RbTLCHvO
LPog4ovpthqVqeylao6cOcqt1Gj9DQz5IDoet02OxU4CTyaEA3znW89ExvSi
RqsSsF8Ye6H/QUwnUxGvEp9vjCRsRpKeKLndjQ6eweJoh8c7l0Gh7m06/HUG
lZhh/Npz/18euxYN91dex6b4osCN3VLjCivGzMLlKx9H+HS8riLULBNQZEez
dNNx9SRQqybexgz7Dn+fq0AYF3jhjQ3eGaqe1K7Y1lATl1qZbQ+7KMwQnkp+
I4R0ZEmbdLY769chLQzS+wYf66yAsP+FgP/1d0hHr7ZYUrZz/Qja24luLNXf
CWpQZhcXx7WDQSsD1zOyLeQlJMMl4oBuzp8NPWfYC/f1dZVt7yCPko/TGde2
195OyRX5/NIXvGfRofBT2z4sRdSCkcfDgOZIAJwi0ERZJwF3sRMaQqZokklp
YeWqtWgEUpIMr6kjWwjFkWLPEG1Jh2h7UfEDBLGtjxqVV2gXYHRu8lJihwA5
2tA48dOmlKSUHeypvoxzmYYssAjO2SMsldNzEgVFifqu631N2OAj6Z0MjQPC
b5fILr/LmZjLnQ1+l+/K4jN/OpA050vayXNREUL81/4lmxcY79gJgaDfT25B
Vus0yOJO64W7toRYNjUQqtBeAv04Un2gfi+CjVCBiB2iCUnUnJex10lLoaSl
D51PizcmH1VjxI3K8PojLX3a3z/9Y1Yrb9HQ2N94uzDHoylATLbm+MJcYhhd
tyMakxNO3wWTS1NOmzA1muyQgO4AamkmRxDU85hyotBkxf3WpZzl+ya1qHAO
B2ffX53eHzAhaXF3tt6oHQV92WEB+equ6JS0dzS1Dqa3zM3XubhZ8dO4QPQY
jJq786e0bSjW7cXJ19TGOoV8DgjYcchVgeMS42u8lF9f62dsZZEfuGD2UYos
TbFsHmEiD8wTa76xzDhJ6V8tYzV4fJS7H04yKmQwHTCZs6eN3pmFezARu0MW
swg9KVLYZzAIAAkAqIreiUHbcEoRsQhBe6B8BUcOOaslE1wdmo/Wdi76GD7Z
Jzcm8ITRVwi0cpnpnloBcAumfeSkOHUrRFg2uDltnNtg3bidoB47pAYlHBig
M5lFd/O8CBnux2/ZF43kTRrvCJq8Xosy0r8dUa1J45NLdx9HZYQYISdEgTvk
dgoWm5g/tXSwVjKFIP0Z3fN7Y0hpwDZMm1KJiOc2X3SluBjuTBKoBHDnFNVF
KdLoghKyYXFoA4mYPubqZMYUYZgh7j6uVAyQlIVbzyDWbaEN81QjYrzSzV47
ZiQqlYa5kjgv8iMlPELQ1gFlXkY7U3jw/X3PHTn71WPJec2JpvBrE844SMc/
F4ki/V/vUN14+NcCLp5bhU5m+s/DTu5kECNUUgeMKaBxe1FoJvK7Psn+VbQ+
y1lPQepuYUFyj1GNaOZFDZx9Hxexd/9OdA4g0F+eOeNUsecggIhujkug9cX0
usq8XbvOAO/eRb50E9LFkBf/zdMNSwOtmvPLQWbFmk+i8/X9v/6t5quOgGkA
1J5Bz1UQFaMbLoqdukjDZYQiauuU9KO5ED5cBX2Ib1o4W1KRF8Q/lH+sPLZL
VJglKqip5V7k3Ps/tHr+5cNFAcnlJ0O0JKmZbHafOK0WAS9cTVq/ioOBicHZ
kAf614xEE3QVx6iH8CPHOlwQLVpfSFOlqfgRyOiqzqQGcAdHLD8plrK9DzFl
XQmY5Q6qXYJrnPw6oESr0BH6D1apP48zEPNASb+dn5a6/+0UC9ayx7UtOmQe
wqUc5WvxBJC7paHGERfanH5MrQDEBlYU7x8yVnyFBkRJUKkPGi5jnaP+Nti2
jU3UPFDswQ9pAkVxYiRkRgqhPKMaIdSnKOOkx1a4cPczB91v4JyVIjflg6sQ
u/Mm3cNK/uHo6aN5KRc3YbkrHL732dFhbLeMBuBjRbvc1j8o9f5LMNqoB5zR
aM5uvjzOCGS9iUEliFY+V+BPaGhylH3cpFu1acKHwLoPqR5hLRgqB8fNtCkZ
xlG1rK/zkdfwTaRkrKmJUURncEcmWP0ELBrnNq0L36fADNjQ42ehQh3j+9ya
Z+yX0nhYyIRDHwouL0z5E6p81Q+aGgt2cPUlDjCTM9WU4EmjQzYZIDGElfFK
lGYrboL0NA8J/k3QIyIv2RhkNCCOyi1pRfvVISg58xE75tFKlmTg+tyqG1X9
PVqmvklSBdO3DU/aQKQQskehix6lOgN/b2+dgqcEkCWseSgWHg/TOqWxx48I
9hEj6Nqw/hQqC9GmJy2OygvwXdj15vTRxIknZe16OqwJb4IJPD6XdjplNg9d
l4e0J42Rtp+6jZDREEZfrwL1O3oaevFsWj3/lGGYZms03PgkUbJ+k7So/870
quB/wUOOgbNJPM+K31gqS2euUy101ppZWyhx2kSI+vuH4ksKLDDMdRZXseSL
VaK5+oKTM4W4e1q+nQNH+eErInfd+qDfUPgRAYLHONPP3yM81/hu7yw2VNV/
m1jNXnc4mv/S5bXrmG6aFpXlGvg1aYbFzwLJKuJ7JyZDHnAEcWPWZhHDUYyq
5/z+8iMe+j6AsyYWL/E39OsBoAca1aUVSlJmN1PvEls99kzfqGQ2Qtq+kVbG
6b/FuJ1EUNJ7KJ27vQMZPzxa/JlfIB6ea0IGHYiSXH4QEn8J9MoTRpc7pF0s
PSx444aps8rEfP3wduMxf00mdc/D3yKnjdGG21RPa8buz6Beba5jApvolFhz
YPEGa0+C7cnuvqwEluLNgN5KAJnz3NmpEt56tllpZkf0B0YtiWvUlL/ODap1
ySFZd11wPT7tzdpgJjU13l6TWIoQMmDKNwMQ2TqKP6ATF6f7VAkz8uO2Y6TZ
Qa6VoWOUDB+3QiricH738PzWTF0tww6WTeO5q8qFY+gqJ6Qai+0pZOlgI50D
APlEvvbZAq+O2JumKic7RqO0Y5BYTivc493rvqjnmS0ITLHNf/yZ0qeSp8Ez
jcSXOqRwWBkGolRIE3KFgWH6NVxQ6lGlIV3lPPqm/2RPLAvIBY3etQeczSqs
AAEudpVsOtF/9yIWMEDG3YJdbDznRnYmdqkqsy7OUmRMf/TSEa3LvmoiIKXm
5/FuJ6u2yfVVBHkrVPiKoBGrK7X5L8v1mPH+5EcCRI2gObCcZSCU8JkLPpDu
H1WUFjMCU3Tv8xLpSI7qW+13AM0txfWLKItsQSC4GNWWiKO0O91B09wA997F
4Ia0tOlTlFmNxMALwd784GTyWwIkfpoItnDq4SoeNueuREJ9aQvoVqEwlMkg
NeuNq7GBSqqEwTJdTjAQbqpTp7tBofThRhBDdVcgSmSPgOxn+Li6eGX5V4Qs
xHh+Re8FJV59ILEzsu3XK8rAaQ3tdOiPuRwFb5NMSioWQgXj7jnYKBY9WaAM
PzBuox+qeTXTuq0YTzPPY424CGZU0EBXFgJLtrjvts7g+sTui9NZXyDOpmhO
fAgILdm3L9aYLdpr9+wWXLPExXf5z7D0ymf4HVmCU14fb4C8fjtcH69f+63E
k7FXYEfaJyAjZMah0w7PaqzddYlNqO5ue0u4rRqP3O/3S31koz5m4OT9aGjt
ItbAWCn2WaMCc2oWlMZ+1l3c1lu80R3u4Nb5grPV8w6rHaigzInDfBfIVMXL
Hbq5muSeOaXVGJyACVeYs8UE2Z0ENR6aDAXge/zPgYaEsPAAZUe+WwvSQY+Y
OXjGLRUiIU+5uIgisBMiCLzcP47oBEWiKzv6wlQe5QTR0e4AGcmL2F2jhiWy
/mNUjvdGQFHtRBL5+14WL7QFyBNQUl/Ll/OjRensBJ0EQTGjsqm0wQ14e6lg
PcrdXhQsyeBWRttd2cC/hLxln/wtJUNQgJlDgkep6y4YRHKitx0BgTo1Ie6t
i1SkjZ9jc6CnO7zC9H1YanVUSjWGfw6+grg24YJb+Esq6yvX0xCzTOYNW0sE
Oouc9vyZCEDVY1hdlTVklWFXgyJ+sLN/3z+G8rWyfP2spiXV/JCfF1Z7ebWQ
v5/xQX/GGriB/kJ0cpgJYMfgj3qVH4TKXFKDAUeK3vWJ5vLuWy3AJVJbJm0b
3SWeULh5XQVb7lcDdcfua640Sfp59RgEHvxfnpmuYLx3w4KC8Gu5/e+LhpUS
dSyZnzO1WA6/dXlyL1gqW+ry28u28nLD1+JlpfogJDxxr4SHFYE8gmg/+Akr
JrAqbWMn8mY2hV7CR02YyTXAXuoMLOTZo18VxhiWGgtFXYExa2lzHN13j7NN
fYGM/a4DpR++sb9jIHrXqW8XX3LgFrJTSIPXT9I/BNbNBrnEwb0epzCuqg92
epPJ+D24csqsAY1f72os8LbxY5663o6cUOCwMLWQKrgJ2QMOPUXT6sNYqplD
gYla4EH7EWjRWnYCM2tOdluhGB3xq/jKXQ4USE0zuMNKaw9ul7pEoYsQpIgL
fz6al7PCAd4l4GHg9J68rn0pi0RS+AgSdRw40u3cllbPUyEoyBGQQ1o/xzO8
wi4TilHAbYsYmeQYJsjJqaO2ZdJO/dUTdxUjv9s2tl7NRIopUcI7vx9eeBfg
CE4NirPoPJv6DRaf0Mdz4LXuvXWOP4sAX47pOb+szaWFgZGAKukciBGjFrtO
zE/fE4mdNRNWwmudoc2OfepUt6dMU6bq5mUXpV7k2EZaIvz7xyfi71JcZ9BG
AVOj4JcXmwiq1U0KQTuXVgvQw62mghnvMKW1QUIryXqPsrJ9Jrlm+EdqFlVz
DQiOEQhVXjQn0Z4NjwkwduH+wgXXVmYL3i1y0uOfLM3NvxGelYapSVIV2OoD
2a8zteWrFRzaQNudmb+/QNBv82E58uAqYiPozE6KtzQN3O7g9hCF7JWBwgI/
m/1QcH4Wl/LwpzCdr1vpzC95dQ+uNkdC4mEGxKRT3358qkYvXdo/EV/IQGR/
ucaNUffOynIoT1tRvfMN4gA4p40zpJTKhvFfJxy20ET6YaWMG/kXsDX1qJJU
0cDgOLIS4GXrQJunGNLt50zYLlRzbh1sqEZgpM/eOHYaI/kxfQ6y72Qqfuzk
mkwUBropH4B8wMID1a1Jg6di/a2hpBjBxHCtJ3jREyS6f8qnyv7n6kEz3c5f
XEkd/8RDZ7XI4U9XU8wmJjgiAz7u6i3i8ALgp7Os1imGuKPLcVY9afKq2IiB
vH+b2BBk1vi/i/XAt13tt+TewQXVrYiMbP/n5BW98HCRwxPeOpGZyXPyIfG6
cqMLyWdGlteh4xddCgeJnfk1rEIaa11jmtPnGU+vwgl5e90XFZK0zRsjLVCH
Reps33hZmdckAD1iODbCvTseVhN2p4IGsVuCHyuexcWw1Zxy5Enmgt8Ar04P
+P+WeqJcIXvzrIk407W6H07Z/dUKXhWJLgqoC3E1gZamYGNcferRYj4+8W55
7n2N7mvr2TThGrIXTHjsRzzxfG+R3i7h9QiCivrxdwvMKx0Ss73YlwMmmxm4
zyddUyxRXfc6jmSeUIzUpPCKffbLd+vsH5toLs23tEltzVw2+EHRGKSHbI9G
wUqn2lB99xED1+GmhuuQsu5aHtoUUL/ZCWadE4w4DZPpa9W9JET+8ovicGk5
cgchaiJOei8s8RcSq2t6GzKipUmT4AO0m/vhpKxe+ykF0wtzKWzpUo0C171I
zdQDU2C+tTrrqpOnPsZ4Tm52m78v9gB700OXbpJyonStaubeRAIhZ2nkSU2+
FfvGs/F757t8NDZUfHq3b4Us/K0r9WzPWk1Ct+GZfbPC2ILrEDOI2Z5KCDKs
ETlJxPUSAICEDCRxWCM08njFYClWmYIFdNOjohivnEGBldkheFWrDpVGIQtJ
lOLuXO+0wM7uREu3tWMf6GOdPlXDetrg0ENyi/FwuzsKXO7TTaYFSRphB2YX
eduHOc2vGwXUj2j+PR/QiYAzrsk8VQtYJWu9mJO0r88BKGwRFnuyfczkQr+e
hY9L3y3UvwmIX8fkxI3stSoHuJhFFyjXFzjk+bmpgjCzIV3FxmFmherNZuVz
rH6Ug/skdVEmN+P9k5LDK4Yv3KjI491nLKu9JIwRSHhBOy7V80V7IhwN1spV
PleOcKorydVh6wQYha6Vzx/opltGQIHilUVdyzv0Kb3n6E4XIdtJ80zJQysz
tAdO9/h4VWBlfWobdpwicFNCPpw2qNaMaqRuTz7zJnESYjvhtwqeCN5icUxb
EWWX7ZAw4U4hYzY5uPzxS4yHdJMdR5ynoKaHWCfqiproXNYmmIRMiZKL7Wg1
IkPT/onDD5rqJlN/N1Dv7EJpVVYc53sVNvQ+c3iimH+TmBh1F+l3tFfoYmYw
SAYdNrfPwef5GIiUUuugJJ2jaDOKIDMGHzWJPL2K92fNGAs8mwPtjjX7FLZp
aWZ3ecUzTnpd4r/1GyfQZ6gIfYXv8TSSzVSvSL78ixWFF4WD8wjpr5yt4gbH
lnNA2Ul1oFcCQEOfkKw42XmMS/hfzq7IexfgQqmeTKv1ir7iNyrqxxiMNKgV
5JW5Ubr6zezChQ/TpxSmZdhgzPXxL51sNAcoKVjLBQZ9zHp11yP3AkhKIUsV
FlHRsUDiOhHBWhqbynObLwWzeI3V1yDZH7QlYj9mMCoOxKt1sC/ToncGcw94
TaFHll0proctwim3cVsAJ+s1pzdYox6HrMRdIADH5XxJdcv6Fl1eVSpbNcDB
avVejAtV87t8pwMhklXae8xq2RcGY8W4ARAci/nCpGYnCkFhdDY4Q8SZFpvf
qqtt9bKJ+Fv6dSnicWgPl6D369KQUTwG1hLMb5J6lcfAtJ4MdIskowHNfDk2
dICd41z7y57j75YNd7vtQzHbVYcCbMZ8kqNPfHBpTvZqvlpdJ5TX3RFJcWkz
j6+w+8WF68Oe0Cj54M8mpVYyZUkQreG8WBotOhnDHacrYIvhIlwUVjfi4W/c
bza1D1S2MGz8YfUo84WFQ7j2SyFNovvUvQPfWG6Pijlas4RiiYgSVuF+lMKI
5eeW8X2VDzrSbkc78e332G01KEeJwtcMAMt5C+5Z6hLAAcmlKi+jDGRaOz0l
gGQC87XKI8DYCYRPUw8ZxLpkR2AvxCn1xPuaAp0R6Bv12YGEaHFxbDT37R5v
XA7ADJmnXoTjC7PxWgACgWvRbsYPYtyoxwQ0DrAJgbqwolsSvM6TlImM0DnI
SVQtgxOZK/CkOUlHPQuclEhXoPkPBtVDtb/jL6r6H+HwLEpZhwhhCdNoIC6M
+hLmMLtD7TuvIPt1jC2Ha93UAUdVAoBzahaCWzmfpF4b/FfQcmTZ8kz8vNFD
1kMfk1i1iWhGO7b3HL5AtS99A+lvv+d5soA0WwGEm3TmEBrThaV5aVWttSpo
abFuN/6A0dWv8tUx0rV7O+lcgk6mAIekC6bji7puIkqHh+liYs5qaRKxnB/z
4xBuL8SfdKPoLmtHFA26FvOwz67Pfc5zult5tzoLTeOOiFJ6n06gD6+B1GnX
8BKN0WdrjDiR75eeBl5TGPpbBe6d0mBrYGOGdPLzBYWBR7UZ/YYC/yJ2pbQn
6hV6seQ0qMBD2ov4f3ghhhovG4CjP2s7a2LPaighBYCfL7TnTSVRta2Vp8VH
buly/ax2ZZKGjNqx8ckU4TGlP41KUGHIaJ4YDYfXFrED1M6TXZ4JUUYvbAaY
ifsAp5gdFy6w9wW2XCpbJpkD822DOm/vK3I60jGmUF1+dBKYjiRI/jre8aIa
034MfWV1/Lgu9GqAsGuDFg4OUUXjUsB36jnbLzp8Pdj49BREuIOOerYShPzt
dSYcJK0DUG/NcNldnxpyqKoED6YdmaM3obap8r/Xc8XYpGgEUfcOQJPA6kn3
sB8b+l4Pd3uEawIllNKWXTHYw7QBuXDRJn6/3kH4soD+b7QmEG5AEKZ/pfzG
gpTXI83x+jh8QYIuuH/eU5uZyEqGGGfEK199TFL905GDy3cdzN1B/cznAPZp
OUzjoq29fBBztW67h375LnUjgj0lgWWoL4i1Br5t4WuYorBrot81QgUDWmu/
gYo05xscbefPawYEAxIpMYnpZw4lGydtXc2vTD2XJMUaQX4PAMlBM+5IkIvA
6uBjt9Ah0LmzjqDh2dbqPoknQlwDFeYRfc2dymnFJhNenjXSaU1TqWytvtM/
hh5oZ2srLjagrIx5oi7wYBMwHRlNck89/jWgz+sXU2gCjPSshEXoWDHKPCxX
I/7O8AbUlxXdqD92xnZ7qXtTqlfdry0hN+BrkicyOga5odzVnetG07MA55+H
FY/hQRjO7pF3h4Ic42ny5UJNdCphhsGINXgZQyCNPAYN8TLZhBX7aIFUWBwx
Na2EXjysbFQGcnELtuPfmwjH3v6oN7b2wp1psLT/8bAt3inCtgOeQy3b7H5F
LhGRw0LlaFkinltsHzmeXVasyrlyMlrdI+4UKORhd3CPm8K3XPfgtfqy1tuK
/G5QW9fLQ/Y76u8QtC5JQAOG12uD7EiFI7FiDpCQ4LlMVsFPgn0qcvI08nEM
csltxT3EfGDSisiaKTnbaKoxjyoaXvQ+FpEgCnHNqVyO2Dk7x3oIKxtEQx7z
FuBEO+SN61YErzDP7i3oAXzp8YwW3goQ6hT2o950+FURBOwIIsm1elk5x9fQ
Pfz5gIs2CX6QTuSc9h9JHqkz/BH+W8uOIBd3PqJHIf9upvk0io1QqR5dGGCn
ywNne/mu/0Dsk8LacfTTtwQhuDzKG+mF1VB9DVHNPFx+YvoYM6iZjuNwByBM
sBl/EYeMJ9KJ/+bgwTJU+672KzKILfz+1Zpy9osbbmdFIcbTSmKNKhq4hulm
ew/6axmhAqJRoqFi5HsnG0QeXFerJV4B0ndcDzHZxeDCk6eEpuD3gPbDg3mW
J0Xe1JLkfBDlHyRdsODsb3zldeeDbg00VVuiNmISJGnkLuOGJfqPpGAHHSvk
wAkZAGAUGySwwI4Xyiu8dBZQ4keYwjZd2BYRihJzF0f+iwXgFmjRDgQeuwDh
3Lmb7Wun0Xv0ASEQSV8Ndv4LBPZzQB1a2QNflIAzP4q8bWKI1Pno6/VYkcDh
mwOt6G/3T7OHK1dsRLC2/U1iLD3NNPIKMFXbtwvjZ4bLYbdB76ksMk8kAryT
o5Xdp2vffujBXLU8j8WX2l2l/H9P0pw1/I9739g3rLWiPA08lcoG0gjJ/dKy
I/w7J1GajA/x2wy3WdlAQT5j6pn+cgbVhrp6y3sizOx8tjNVIYxk3UeNSGa6
ixsNOWlwbJ/mlCekr/MnDFJDnWHJIbFCsJksDCSnBLujzU+lvQSTQU+Xoowy
Y12P4TcmpQ9KgNw5zFDSdWrGAFWC6H40YDw1qaQyY8snkNCnHGNun3A2ZX5v
spaCvw+OADJwvI2SkylVKj1Af/7r1ls3UGnb3udMj81TJ1+ioYHhsoeDIN8i
je/+S5SnewN9xkhzVygMYhMDcUEDMi3B0ggENVZBF5Umdo0JgGBkZXo3BHwT
WHvt45WmKqEgiCIaqoEN/0VUo0KYcTGoW0dmFxSsg85uVbz4MpD35VyyLXTU
74IaU+OD+AGxtLjNvvM16d3awjaUMEp6cUjWO8+M1ubY3kCseVO3miM52zNb
VZ60oT0CBwfk/8KNyF4WFN6MS7U5ZfcE6fTBvK2OjWb4crISzjhLCNu+nFV5
3nJxnd73/h7INostdJaIyrhNDGtZ0ck5YPpkO63UbZmxsVT4Pt2KzcK2rsRi
adNBWtl41oEjUSECS5VZ8V/9Ou+Pb//WsUXOhi0z355a7sr+9xWbqECjwbCk
SVaFa7iETe9sSHt/rqMG6agXoh0f5j3sABxaLpCURZA6HupsGQH3f9jHeVws
ICphy3RwZl/mFO8ZhQFkFHTGJLWUVP4Aq+wdtPdHU+Fu82pnz+cXjDXmc3Zc
zxM1dGwePmfqw7YIR/+41EoJWZnxdUXe7jr6Kc9Z2lSdKpxmDY3lkx6osRHo
Dx5Z2JIJ/83+yrD80wQV0QHbZWZMna7Mg7FA98kfaIkPZ43N1Vk38Ui195Cq
aCkKxrQeZ3Lf8wDTaLvENLCi59Rz+VJZEgegFXbd/sGViCVIfTgabUFkXTdR
A+BPGSerDbrgXAo/xZNEmfTu6bn99SdctH6pS5azd7fybr2ciKi2v+ps2HaA
TJ1oK8fQIwmsfQ1yWSDd1yQ6UoA6JB8BQ3ou3gbbG9e0zaVc1Ik7VbqB58QC
1SYe6/HiVjrNIBucFXK73iEeWjtGYwgUSoxBpmBXT9Gp8dyi67Mf4UR53IfE
VRmQuTbez6MblrNF9GgE5Bwy/4k483j8eHmQ+fh6WJTGLoyI4GN5EFwMpYje
rL2APuqAg7yQt0aLug+PM2s2lzF9nKdJ4jtN4yteva9r7IFJZDBNLhSi9tlo
1e3fx2m2Nw8U/BDJQC1luAz6hJyMRfTYPEDOV8HKYuJM4w2bAIqm+S10aeAx
YpYDlIhYZH1hSGR7CxUamysS6BFgdv4JaqWqAMScW96kqL0nyc9BFDN61Mwx
OEIoatdaf/9wZjLQQ+epBr8hm0vE3t9mj+GQExD9FLiY3e6pzAqqNURKHbgc
W7LraPnH7HZxDxjPUvBrk4dGRotDUxSaYuYxxmvN6rF9dR2/Uj/3S4IZPph/
Ke1yl7cYIi0bnddP0QCVmDv2pF+2mGgtzU9lTF/Bm3GrLA/SPnUJUsc062mw
obIH+Z7LmMcmK9VWuExsYl9r6kQLKefs35UoINSbdYvjX3FqUCqsG9qiktA7
whiv5H+ECLwpcxr4V2A+k7BCs/9CUjrqkspz/+X0r7KMjjJDs82/mE9N02VB
gxdjvmffB33WM6bEkQ7YRBxJSvHicEu50ifacqW0PuGcsFoalgSTM9UMeBzu
50c4JTK0zTXFaL71XWFHgpB057lgpDe97pgBj9+G30BUJF69hLaz3NO4tFaF
fAOw4D6VN2AZ+ShjW5oCNlE5hQYuKgS6MdYMULfPy6k0X/6lmQ8kTgyWLKpQ
blM1t8ZYbDzWCtvsI+5S1JdUTdy2VKx84H9pSG6Oihydhcy42VBoiIofsru5
hkHl2VjsSEoFLBn38AExatA4pW/kpA+tWKhQ79pWswmg1uycmMLh0umSN417
2DvuQEwr+UtkXTwvEueaSBwlVXUh3xGIu5EYtXwRtVZoPjmjgNer6syp0NJV
vuWpgmpETkMv1l63kfYiwlqb4wdBbc5lj2T1BmLVtRp/O85McQf0m1HKTSSK
hXM0Hp6bA2MS5lGrCUhgHnIwrdBVo9w+M24pG0CdGDIBSR2ER80nWP69M8K9
8ml88SPeowwxNO0xYLNNnvlV7gaYBle0YGyWTvFQvdW2F6xlg70cGlSghkO6
lHcMRlZ6hEqpETq9gZgvjtXbRlxUba4RlfL8b3AniY9tGPBpVVAoMOw+NuHC
EFUWybtoDa2kuoNgcdqfLrsrPCBuJjSdpWNK76xLSmqOp6/FhXlB9+jWcIGf
hP3uLt8dAnZ445Zc79jsnBYDXKdezs1jkUAfglhMNU6YwKus6TYj1qt64S56
lhzRkVMWXSVDoKMpsmdP8rXRonu9ou40I/H8qmpzJ4uhqiSvyOh52T6+jQJu
gYkNsZb3dzcjBHB5pu8mAmayQ04NfcHBrn03nUGqVIIk+KI0seiaxeneB6Gc
CIVwn4J4goBGfy0qKPnA0eClrEYCrbhEUeho9Qo5tr04WFwAkRtWosmNQCUT
vSGUT5fNm6c6QhModDkY52HzD42Bpv6CXaGDJC7vZr7tLB9HJjxvEbRIV1rN
eFJgEwprNKW8jFltucc1EttL6oAWcHaEROAx/j4Lqpody7ljOTB/9bPq56x0
QMCqQjcw9p2w+EcuCpeyACufLwSdQQZbZHW3NKCvWbsNLGEYT4+Gtkfi5fU4
buTXGe/imZkkm3LvLHX97UkrYzPQoOEx74qYnEbLxtkVwnVWWCE95JvrOEIX
FNqU3gJCfrGuBqgzxtIerPGcyeLBc83Ihj8MImz08Qhky3gWYXvifD1GZiSR
0rY2caTo6Em5FwyOakuNcLo7pdR9URNc5/9Ei5UBspF2qHtwInh3YLPHlwhF
EPmv7TMKCHkhx4RxiD+HIK29YU9Q7gQjMzkgCYjKsF9atBXtlIoz7lIF31Au
1CBQSv2WlYlEcciA+Stnn7UFwvdrHs1eRSsuCmTqKj/Ve2qRo8zfCaQSFAuN
iz+kANBE9j6gxeLMY7yNbTDA2sGJg/PLXPqOXtZjS7OpC6JJ6sgg9CyM/C3T
NuuKn+WtdQfPNhkJr6Aytv174ie9CwDCAl/R+jH5WBPIFaUD6PoiHJwh/BWK
5Ln6agcXKW0cljkXGAJ0bjF/X3Y/QRjmsIQtnzV7ezd1Zzsj3GFbFq44jRvf
jq9QpTMgvZgQq9rpwmNkT4TYuqtjF/XxIm8sXyNmf4yJu95beNHXr49wo49k
exVhHhITGrh4q5WYXogGciCeeB6mTMZH6BnFhcbq2CJRiRz/+TdMdgjBLXRk
0rxE9/aSxP2MQB0v3mKqXz8l2yhCzW7PBj2Q4GY9TlgGmPhEiJFbWvAqp81u
COm1XUQnRRY9BR6TvgDHQvUuAQaOOJRnB7TXzLfxTpj57g5wGEvAznSFT19g
bdqnkEOTgzGE+mcUHvn769GDkG6+EN/xjIVX2xnXcamY/pyCEO/KWqZa59uv
Ks/J6dqtmk9Ws8JL0WCEReXngzFfT41x51u7e+wf/vDJg8RePoWclhniLSnL
2PlBNCz2nWF7cWWXPpxkUs2Ig3KZfH+m6Lf7qNuwQzxLvnQFswWhgSWDJ+nw
jdGF3qGOgDmaACAsjVt77GRIUT1brEldbfFtx+1OO1ziTUnyDnaKf8dKpKgv
JjSuZuLVmX1v7tkIm7HMZXGoDSJeyNP/B5c52UVMokViRJXArVIgxTfezp/D
o7hEO1U/jFP7IPIuJy/ZuxPB2dvJM5IylSKPhIYkgzN1deD3Wz2m1pEkwrlU
SpVEtih76Zd3LGHeDjr7tsW9sMjxxcGOXrKNpzU4zmQR/3ZHLT+SmRLQ6tTm
lZBbdbLAX3EgSzXefggMlB75cYQu3w1pPilTAm90kLvnHcyXGUo5ddQPoMEY
P03flPwdR9dWBYHITzFuAT2jAqwkyZ7lWqTlX9PQjB/HQ+3Sv7Sq3JGbvVE+
96NfwH9CEm1e7SaGXGhGE+0yKyIrbZpn7LWnEs61A2ptHruFMuW034MB43FG
X7DdC2HPJTdnOy3phnGXMFJuQOroKmvcu9UrZV0MkCnVei3EzGZdpY1Xj2LO
xQJX1xehsYnpXiGCCB3bBP6StnYcvZCZ0KZpy+8kse595tYi8UsGJTfB1S6i
/NGoqhBrNmFUl7BJmAQo6a4rHmO2bZMxKXlxUXbSS1ax/aduAP+R9ONeLEag
3EjDfN2u3d2vC2343ZzIpmL9y7GT3mdqn/6GzO/IlnhsBO86NDrEzkOz3If5
IdlPnRD4P9xu91RruGDzmx0O1liS2UHzaeoSNDRTDNCa1ylCXnzwqb3B/uOE
0V9ALGHYZxyMl43HsTItx3Wlo7MXVr1fWnHCMm1FP+X5kTUwnFBtbL3qPHyM
PNtMOry1jy46lrYYH+7FWUDRvuPxRpFPNMgKTxUYMUJOHeTCEt48zReUJqne
d8hT/cdfweqjsS50szx0ZSIUCYQi8UjNx9kHsKU2d3tD7CdMUXeeDHReeSrB
RD/J28E5t3apAQPvhyXTBFmvJsyPXqQullAUr1XhL9tmhqbawbkuPzsGOXmm
nlrmiXmkcDV36nM+GeL3Ot0xiN01WqQi+1meggikB80Eczzq86U2jNTXhCVj
vF4BvrDeFEtdxW/4OStleRbk4bZkH7C3yV7BFvpDCN8pqnBts0jHwsnlk8yN
I/qIwSDBflkkXVwq/HQ1g9bJye8bNOoIptqW/wZwUMOY1/v6nsq8FCHALHGm
4xU4n6jmZhMMteTDoyRQwgf5H5MXzTc3FZS3vdVLScXIRZDahKFKGYngfhTk
ggcP4fiMtpjp4yrL0SQEeYQYiP721NMStU4H8S++znqy6wKTfmnIuOX0lFJE
AOV+AxC++jcQqnzkrnbzBpe5OIP0qGavcdiOV//HNIhloeVEto6kKiDbnzuQ
kVr1+jXlYUAQYJgd419pgIFlj0E8DTshFIZrnnSCLcV+P1LFKzyOYAjEcIQs
FbRbO7hgT6liAntumf8M38dwOxjXy0XWeSTo2zCHTqgOZd2S9ViNVO1afIB3
iEAZOqf15R5+c5By8J/+GCCS1ha2QbMYLG5KXNNmDz7OQyWhRVRe0Yb82sL4
NNsFcpc7QBBysS5dOxWrKB1R3l53VRJtuxRpFmAkV64AaFDpjt0djdITnsSG
0T/XNCfksXxfKmZ++/jmkbQDiMxfdctooiV6XoiT1+RLTHkIlBPj+eImh7oI
Nje+qi0GRvwqjYB23LI+q2NA84axUfb94n5U/11/ilemh/ZlbkrlbqJuU1Qh
VMXjmF68Zp7STsXttXZegkOjfyuSqg4pm+rPxURSyAweXNdl8kTwacVIVgi+
DdwrqtFK1QADzV83SHlnX4+i7x7FMnIAzNgH6RCUhwZSi8qbchjbsWGh8R1F
n/cp0Y3/lfPaSwsrZcC0OPNS/3lO/k57JiyitayYVUs/4bszdUrojXS9KzYn
4oEteuo3NXZO1oWLRtfuRuEd+AyhkSdo0+zXpW/UjYacIicvjFNmLcqgC51v
IpIe8NqPiJ4jZYzxFWFl3/NBd53pLm+ObWrxOIULyAL1nwHT7e56M/HztdSO
YcdXnpKY+oLN8FckKl/8scqcDaBvvJJjyca0qvtsj6WEgHFeiVr+YH2RNHaw
H+IgH2MOUmX9H+ZvGS/ljxNm1bRfy/Sp910zsXgXE6v2iASAmHypLErzln1q
fOrTsMQ1Z0vsa2mrQbSI/EFFlmpvJEayib98Tv0d6dKLDhzoEmdLfD3LGfB9
lEX1G3ssjEIYD9MSqbB6NIx6di66owP5RdLP4+2tz/agMHeh9dE0MN7urb2U
giMo/Mz47LiQmL/f7dUJcarAPApTbtM7ADb1EINRsftTELZEJnkmImOpIgtl
3jhHVR24rrA5KHNlPqSCT00DwLKYZ2bJmAiOa4oSJ/Rfo8nYnyvpeKZRJ16H
20Z1hzb8xX41evU9DSe0AmWAqOTR6mJP8f7Tdm/2OZwpxLMlSAyvWcvfKV2C
RUEouFAveXZwAVhEeWSYcMk82mCLSMSIPxVzLVFbP9NySzp913PGGsSSllBK
fR+uhZXnxUdIHywxF9K3bElggJGwI9WufQQmgHUx6F44UWqT1WasvF/mytyE
SgjAjTltFQu08V05SYPhJe/RYaam9zzt2kblHzpCWVeEMl1PXnNJPP42sXRk
W9yFgBBSLWWUX1dDZGjE36iPd4Jj7zzVudeNPtNebBAo7IJgCr5K0DL/4O3N
k6GkZLQ19KjGHBOZwR3a/BG9lwbxFiTOn8Jp2fmDborodeoq7p1wHFOz//4S
aXkp6H3RKFfgZPLYa3PQyDD8LDo+LM0NWSWUEGc7+ZAaxXVpJSIw9UjVKufA
jInRrPcsLUxxWZ6Jvfsmok7LUc/h9FNqPFUT9aT9oxrk6RkP3yG2ayIaGtzt
wNqLkOcqVE4p1kg5j+aSPAZhhyUPD3gXcWdF4MCKAz21apxJvJnBF8fF3IQm
AJbJByjtblvh7bC4KqMyMPB52pIuL3T7e5XuEynfpxKVd2G3jRuH6mqpB7iF
D4hqqSNe/+FN+8v/kChEaAqxtQcfIaioGJ4HPD9NL2BBk3tWp2zuNxi73ku9
V5xkfqPg8r0S01HZ5MpmfNYLO7J0vDBNU0if68foZyJlIQdYtc6kwPOSL2Bz
ofu0ungtfGAnCsK6Ki0F95SoV5xhuxxBhj0t1Jjb+8O4OaBXwvSRdU57hCNR
0jSekw+Acz3jlvdFZUsiuMtLYIllN3OyWKKEVW688pexZ1nE1YLK9FTUfaBb
FjGVDMSd/XBocp4naudgKxntnwa8238uma8VaT8/WizMKoQHVPBKE/pLvYTF
dL7I2oWkD96jSF1pcPAWA0JQmCQDu0JUfdkBcN1hR1LrBJxKWMeqW3avuHXX
G7UO3dyRrNCk12QdVoFrSaXFd5bBcvrzq/mrAYG7IzVd0gseaZrznzTCArGh
xsQqyOKbu4y+aeOEOE0+PRGbfgHgbpRYFDGm1JUZloYBjCsra0FynCSzKubL
fqYMnQ7oe//y6EGQXLV4wCqQyAT3KKZpGZsHaxTVlQbc7jS/S47DqWo+qD+A
7gUD7UDNUWZwkVipAelHwxt4zTp+qspBKMeLF0H3ST+zjZe671f1xvWE6LAE
qWE+uR9eJ+nkU4L+EguYU/THi64iRKRiukxHfi6yptDDsyaEd2VhpoN125vC
nKsNDZNC4A+Z4QeHL8JkAnkYaeTnUaUaeMFY23+KcItkyA+ALCFo2C3eWb72
Pz+HAtOTb9j9ZOUm+BHo2GKtYqYoR8eTZ8JufVsj3m/I+NkEjeEvW+eZZhJa
ZNLarzdf4hkOnDuHfZvKiPdivlNzDo5M4Ky0KIdlQfQUBR3+u3J4laDpH8Qi
oiwKUA229+c05KseQEd1HXXSwTSUseJVL+kZO+wm2+dt3qLLgRvvJTF16Cf7
zmjl6FOhRS2/27W/qUJzpJvQQjo5Oq/x4J/ltQlHH/FA4JxQHkp94jas5HB4
ySuagExy6e3bBJAXDUjC323Xya6075XWy71HT4d4wRg5LnOhbM5AaYOL0Gpf
0YOR+AnbfWlTYpIFdGLU8MHMJuW7S82XCmn3wmDiq6jynP3SnO8rkEAZWdde
Jv52awEqjiPDL+gXL3QJc368de3mDOqft1sTCz5i14MQepIgqm+A2qiOAGqG
GLuYU0Z+FeYYBTH3ppUzTNWNLCbEALsBHEMMC1oBHUEm8D4v9IasULSQm7Td
2cg2GjjGSWJsUYTNOL+L0YG8JY1KT+A6HjgnI3h4hpIB+UkLmdOd0SSsQPBc
TMX0VPhD87s0j6y6M652dL81H7A3SPWCAGOiS/YfDIgwf3QN4UDlG6zMG6bz
8hkUMbm1bT4hSRxkZ1I0zdFPnN9nBzSIKvDZkRr335ipzVyN/8P9bjUT4Nh0
TRsY13CuTbM9S4WvbKcwn0lSYcKkmAIEPKy499Lc878mzR8R+cYokWpkihjw
sZJ4sGtChMOojuD3dqGKSwNzhjlJpDt5lJmThFxh5aGY7Y0eJo6XBm5+7vRB
X/nv/xFlXDGx/Mn0Kn9nCA55Q+KcgISKrBJ4yESPMlNrKrl9/ZL2b5FfzfkO
OcTQhRv6UMdnwHo36f9oxcnuPV0szX/luIrNp6AGFfOZTdoS1os3aalXcp+3
RVlDSuWq7BJb42Wekl0cBqx3TQKAisivKiNJSK0ps16nAC+MIxGAo7s+Q420
nhJwMGKyaOwcYeYY/cjADSpg+8JktONw93k/qkbCx+iiUhqlFD8wJDt+tHER
M1cA5IfO2xz90Olzsg2cVpHbKU6IzYQGAakM3VGzLaciNnhPGt8zcZge7Cd2
1Xrh7csfuSx1xAlWYvc/9gRQQrXzf1t0T0B3cD53Kv/oPiM5XAqxs6CyOILC
G7DU3fpOlVSHrJ1lmq4p5ZikXBXOsBstKVFGSoErTQxwsqLesaT8n7o+iPhx
h9Lw7JcpN+iJhrj0cOBXPpq4usu64xvd2i/M5y7nLxY7C8bsDiCgAfq/skdJ
WqOWy53pFjwvoa+ZOBBXDqmfN1eFV/dMDn8lrXsQu0ZKnemLUUo5LH6FaqEj
Fi2OEVl5LNq3LRX/0bzRne15K9clD3mjgUeevukwvU19hQe0nbCV4rXsp5aE
XBMVfzA2dIMxk6oS3+m1nzzU1WbS8bIg1e/mqBCZg9LOWkl7t3e9leoUGlD6
xWHPks9ZPYPRVmmlENmIFrHcylwfSFa/aBA3z/yTc/jQk7vlW0jHJfOEQ1UF
357o1V4MAK0Qusf7DezUiuf7u4SMC/mc2/VfOtLsz0ICIm3gs2WiAZ8ysqXh
QZtLMbDOTIbeLbwrEMzAFjHqRgGpgdJ5ivNci4uWNnaZEhhyg/uJ1Fcu02Tg
ON6JaD0ZLEp2EvYX0/qg0UvwKTLnd3r/FYupq+r/Ov3bJg9hHxmvHTZsx/Kv
Ytr6b7aYACYR6M0iiwWzizXrRItI+f9pu8jMxsuc5yOAdlDl7l/qGjFiMGZ7
eDBfT53LHViYeVQ/KgrjweW70vkCVYrcMWR5J3sysrHnEqx4qEqzhhLRn3a7
BV4t+kcOFJP09bSJAjI2Jy5xrPV0nRsg7AUL9a2uktIG6nTqfaK9DGaF1s6i
9zARodf+DccUmKF9fMyhuURkGUZe8SC7Srma54Ivgn10KZuJzfwE/na98S5n
6OQBVlEgoAUsM7/kIUxBBtReqJNEBY0lwVOou+iksRuDPiqH+pcXVP01O+LE
b0nPtS/0mtv7U9BSve7YfBVcl+JXTswz68lYc7DcBCrenl+S2IrSZ/44LkoW
rHqife8qAwv3h/6wDkj0XBm9WV/+aJaUMowHbwx9dG+qnrvqrWluqvi+2ZuW
87u9NTRiO31K7EmL3vpF9HFtoDmpAGpqMPCYhs4mW5Q9f4edmLseL8X0yhuh
UUk+pbWk+5ETLsj68Lsl8NHMU5Sc5ZuWnZUKCebxSVSTn5UcOb2LksJ1M8Qr
0w0JctegBxHvMZ93Q0yVdfDTMBmAx6+7IOrwFoLgKhGyCZ7pbKz7QRmrf42d
1xdr/zB8dUG5wWRmHGSwqVoiOUe6rEZJ7wNIM74ZM4ro4PPwajO2psxpIwOH
l2r7ga5BJQyF8r76AIzLOoyhvvlAwnWkJ7Wh9My238hYGsDTBvoXFPvCGYHT
KFKCvuMomls7VDLbqtCyYG4sQxGgeFHKjWn4wmm0tamLVpr1EokK7T+/Urj0
FHoUJuR8gZZs3QiWHdnKbq3QZvA137K2FYMz+hcV7TbiFzpxxCCIBeG02JUA
cHo/U7tW6QM0K8csv5/PATYNKU6F5C0wHlN9ftaKfg/2YQrG+12Jt0L9ie7I
6qXJGoI0KX1tf6kAnYxckSR77rDf64fE6k8ESZqrbA7cqBAZzDXdoxwHjmdp
oy+XWVgM7wmqfDF1GgC+o6IhDPdwg/oH3PRLU+j4TpePnKVVHvZ4k0hYp2B9
V4l4mTVUdb5qsHleMaxYLjXErZOjY8FlOzYeL2jfDiIob/MwosO0+QwNB3w/
sbk5Fv4aJb8PbV8JZbz2KwyYBfvlW1aT/nxCTl1AsvF2J/YJrqKmB2bo7G4e
AtneBsUefbnMnMbQIA8/He4kt1igx7xuosYN9eAMf/lSg+zrJGPtJqr/JIUE
7mIyJouG9PBGPWK+B5ncY/uPmsxwR070ej8OGQUMqC2YL3HdlFFsSnmI4L7W
hnWnHv9yBAAQpCTxZpUjlqeBHQPRucSQx5Cv5Ysg7SGFo42uFBICf28UeMEo
INfZDeqBpatIPuMGmaxXC9G53J7mkiPpdd+Sc7vkLtLfKLnGFqU0Nhw0+RFh
tZSs1OvOzxh3euBB+6ugBrLE6QQtjVb4HOqS4h7b+HHCKM+CR6tudkOBfmyT
qLs3ObV5Pt3Sg0axl334mICCpPD0NcYChyqkV+kA/pKu4+aLhwS5X5hZarxH
xJpfqJIDrFv8IzCkI5KXbxq9oRFr1Wvmi5MHal4OvX4H4Ncu/cJnfgY+fBN6
pvHVu9o3XerVEfWZqmpgL/BYZChuzFcGaE5XY9hTQ2Zrwz+/gRxknqkJBXjv
4OMF4VoWmQVS3r/JkQQ2wWPg2fUum37RypmljcDg6CwilU7eWmvFDvEXE8Aw
39uuGLGyoB0fuEheULfJRQBWlZ4w9pb824g8ZpSb0JqjR2hnK+FjXeJRvuuN
InMi4Zl5H1gMxr9OgEYX5tYe2wKla/ZPSMi/8Ot1fcS7UBkzjOXp17TBIOHg
3AzaDNzUeULNMtQ6De+ME2wJR3FfD678lcB8cbgh9LQ0SBZq6Yi9rZGemlxv
mjp9thQRfUWTimtBdT5l+zVhG9MO47h6PvA3CnJmW6D90IoHYGYLZUxsS/gk
JrRpezppFK13ru8MRH3sE6eTTprW7ZL573FGQWOGkMSdQL0MM4/5/UnHuWMw
UM797IHY5/wnr6xq1lc5iyq5snyjrtQoMbkVmlcCQJahy5PGl4+UOfaAt8uw
vfAzNh65vfYJsPJ4hqzJK503PGAgCCKrsNaHBLEwsgi+1A/ImR/MczJ4A6Xe
Z2in6ZJkEB8sGTxw+G7z4fpJP5fy+EiA6pBOkYfb1n887MvgRKeuyofPBOKz
BeJu+fNLLRGzmv77J0ZgM2E6zf9YS5c5mG8SrRyZWiQUVbZrVFLzbDlHtsfL
zedp2uaPRihg/Tr/3TDVfuwH2yWtr1LO6di3RhVooTpJ4XqxPQSHzHveXCY+
F+2YYXLFrkq0weNncHX8vTmLASX/tZgie5djNv9XQK/b5dbWsxQg9pwBkpKj
2xxCpV33GmhtzqqwaxFwAxaDFBWhKDeXpQeejt/9sISHZMAS3kDnm3rFMjdW
G6V1CkNm0gOFTmILMcMjHFdi4hNYm8arQ+uc4WsJhga2qOSeARSrFYTU+XGG
ZL1YsirkgKh7NrIEMYsXwwn3rTh9h+ZKbebX0OzP3XF7G6v/ap4t2SWVnqeb
63n2UOe4xCtvUTVVQ0APcUhjQdeUuacj/1/0spkM8ZR58+1tbP2GhENw2Kfp
v+bECOCCu/Fv2oH2hqJpeZE9Zj/FDRqOYU5lXojEaKskgCMzwPDyAk5LBTSg
vtt5/XuyaV4J0wZCkiP2EbuktQ6PGlEuATVti0Ykd+ZbsawLBD1GZoMUMorp
9++ZO8HOAMjayAppoQixneIiz9tpdP5jfP95EMtgK8lGVCQzwm+fs9pBcqld
ieEPt3DqgXxl3B+Sg4KHdi6jcL0rIJTDWyLxpTsNZsgp61cNXvJk1o657QVt
ivNP9sTBwl/VOgo8rFBSCsJQ0fArjyEhv3Snd5BzszdFpiga0wuY1pEL/oWj
d7WSDb/DRzWTiT0///VTzvzHwMuOwpCv7oaQ1X36E1Myh1SH65pgb2iIeODy
LYagHhvEBYwM7FAttVcoQzbvtFs1l+JUEy68MS26rQKYZ1vuawcQNqj0KhPP
HL0JdVbn8IyYXlXBCQ4sDJf3x5lhX7Zuy4Qyzgx+dB3QdAKzUp3wGeWeVj2T
DIe+zEPzm8ABTpp3Xmgd+F9nXzXoI2EwZIWZK+wkMNQoV8QjlQ5I5k6qojT8
fNnh3YJV5o2JOftty3wblQBU8aK48m25THOeiYeB+GjGzu/fmjKqVzEkZBNk
x8T+6hHfm/tgD+ZqexjFsa79B7h3Pkyz1oFcFZpuSAsi9alb3qLBHAxuPtHd
Zq5VMn7LJlXkig4tLVO46goDrFEd5E7YqlR1t8xPc0A//aU5vHJW08Lt3Wmf
0kbB2GCcF/u4DGnUK5wUHY5mvZax3mhpprlf0r3ByxDJ/ZQ9ERvtpOJPAyr3
g7x83KQP25cMYjfHiUyxWNbDmJlOOFGA290QPcB4TxiKetaL3KiJ0ZLTcbPD
7MrgnfFD4jRNkvZhFbTAg8XOLYm9Qp5v1Vfyq4LBcKXDFT0vbI1O3FdGh7Sf
nnMBRjFnF6N+BCOft17NFCDE/PD8Z0/1EHMbM43tnw6xwt4dVX2iV1fc8EEZ
zEKNQWVoBq8WzJdMi7MTUxJ6m9TK8n0dDnwowQner2XVl6g1l4OJ3nltANTt
5b2Z+HziJoH1jrpNVqgFmpri22t5P7T+ZRkw3fMw+P6VDacwWzzTADbx/BM/
Sz21fmvJDpIlGmuezRLKCZJoi3DtIpEodV2zIAOABtUoBjSyBtMsZdyNQ+PW
WlnehoJ6wr3LdsvWA1s/i9FKWwecZ1NO5Q7Owa6HjWMyLgbDbweNIM5ZY9xz
GZEuMb7rXJ48MD4Mme+NkGHxrOzh37+pgz7EWJXWUgBPyXPGwKppn14DNhIw
f3jkfhX1Whra3AmHO/lHloW2K9GGb8mB7RZCNQ/Y/McE4EPtCC7n/o6R4+We
4UNcg7PqfQX9MgXrLU6A91xg6qNSOZi6d+RasYkOZ5jq70DSB7N6fB9jH9c6
C7uJwPQlz5sn+HBB0AX2gr2Y//ojOePXFe6nym1Z+XjyaEXoX4lqd7nF8qIK
aquIlvpyM2A+AaSGRp42lHTmHUNpW3PFkPSiuBNJhbKVPM6RkK511+Gz9tMu
EwA+V01qbeVdMG2VFKaEFzBm8S9QF1KDuupv07dXAeEfd4+76jP/FtrCYSIR
bY8clzp/1IlxGLwCxwbx4D5RZvkHP+22P/9u1AA+Zjwkk0b8JgIUTz175dUn
FXJ9FIMmZhTEMODpr01rPsLnYOHOm48ZN/JKaCmmI+i/XqeYaPuXaqUOnquP
JriglGiVtkp76UtPjdsHysYorXDMP54bmKb5UW41TtRgB8PcE3yQwSryiUuY
L0qnXX3VgDWle4RGiXYB4rBQsmW9y58MR/srVvq4AHIIPW72xwd3Iisj2Dpd
lxO1dNNa6/H0V74Xyb6YXL2l94/lWmEkye25XNQzjWfOwqSqOZb9+Ehpj+q0
JGD/KumhJ1gd93j//wJ14FMKJqTJx0P3gRhJWhM00qCKFwCQLCs64MBqEQxT
CZogmR3QVUzxEH4fveNdI0eTK+xFsXuK4+xhXzVB2tbbASFNomaxADQ9Yd6p
C1yBbOLdIv0Cl//pQWrtnJv1ib8srMdx4CX4W6HJFjoA5RCcqrnr/yoiDVMn
H3eP4/F1JQBYApQujNm0EVeShubcz0KPl3Lhmu/M/lR3JOXWQDWigz7eGGrG
CYaTHK9/1M7qrJAa9zPTnv54CQLb31sgDSYN1x/ItR4Jay33RUrXWMmhrGq3
ja7vgyPA/JwDd7StkH4dvj2HY4X9ErNTlEHZBoLfAoT+c2olyz5BM2iLAW0u
IO0F1O5JMfafwwhdu2LxG8I996rakfBjoTV4OMRgQiI8aoKdqWMhabJIum5X
8krNrF8iCrgNICg0quiQCaNVkp1gAA0v/7zaG/Vxm+ePW7SgmA+GS1XTJj31
HyRCmo8jSUrsmtsCKljgqeTfRaGCHJZEjhc9sOmnzsdz2mU0i/90CXUNKTtF
Tv1YJglzONVtP38ZbnQREAuhNof742p8tFk+bf7kqWpiK/oJJXFaKhGum710
g7477FwNKJqr4lx3WYAAYLNK2/EjsXwkyzdQs9NlrH3ubqmkQJW5R082Geqp
ffMMY7fElH1ifGCk/mRfdXUoPlidjjM+ggK9+cM9Y2QBXaERt3Xy3PjNdzNY
Ye3qs+Q00zPQW5Qg5ldLYmocILMy+4209ePJKkFaKIM0rQnz393Y7nmCTYSi
XBhQAkiPFrsVmjamOk87aWojMRERRN+OaknhH/uMDzQwTuMNm9xw72cgEM4l
Phy4ngSVN8Fg72e/mm2an/BHKV3c09p0tgboEOVm2xT//amTRQLvSugBaXc+
shZ55GS1nB7fkUPyPsOdalyVIZleXuTPUqjlBfVxKoC3xZuqHHaucuWUwOii
oXbhTnPXEvR2dzsxTWnf4B4YlIW6nTKZkA94hu8Vat6wYqBiY0yMCQuUfphp
po2EgCrvAG9yORCPEgEZrG3esYScdFSQiR3bH8SlPp54HNXIeAh/uWQrRqZU
M6E/CUYhxAioJUZez4brXzT0VmwzYO5c6VeCCO/WPY/j2JJIVGjy4NGeXCTP
FZQZn4zo4CntE8iWzBNXaKRJgstKyO3gQCWkdUd9dBwIo+phmFrEChojs7FY
DqcSODqm/ch3faSy/cqkhnVcayKFx/jwZb/LOVX2LZxtBi5Yzt3CFUXwaqMs
499gGJwPIDKzOj+Vcb2QkEDDEQZz0f8L4bbnhYyVMzlLbzcWbJDz6BX9cXC9
mD3s1rZCqHlLbY52q1YCq56p9TVcc5L1Zo80T1PV+oxyLuxM82N1l8ehXdMJ
m9P3bE+IGIZgDBtWsvrF0UtYzeCG432BoAY17q5rUn8MY+uE9BWwhtYnPWgL
kjqhdhUVHrfqwQwYfF/sZE636dU+mMWi4V5vt5w2s8qA/nqi+O3PmwWffps7
ddCx45yxSwKX8lj38xIP+H/ijpfLQnEybPnv502sAYjSgSauzPjDqr3RRKjP
d7exWCOcG4QJTgBLHeYhpFG2jq/4HpqZ/6J0qx/y16S0dPrlVzwojp3hSCIA
4A26Rd9f7Ez86zY2v9vCZyQX30ig+3qytyepdWPr6qwh89oQHljXZWlCEgyP
Nwtn2am5LxKywrDIXvoUTxyafV9Gt3J+19mKZvhWxmoBKTr2GGiXKJNwCx/F
s2JB68lfkuGhWkXjUcT6c+C/HApnqUM+c4PyX0rRLOcTyCQ6Zec928dFrh3M
i6CqZGHEugVy7Vtm4EBsaC7Ncs9N/FnBHeFcTROmRAUtJsXfXhdekSc9Rk1C
KXCv1jMTQ/4LkHc88Td7ep3Shb+LQmwUv41xDkIri/nc+fX3USYp9VqUOax5
uo3rSCDV7qNqO1GB1FePRX67izK5ZV/iOS/CV4y6KmQ0Vb3AEKXwGyTWDVq4
Ce9LTek0NNwr1KJKG/+4F93M8M1gqmO5+ZUSCzaKYuRizo4wpiIiMc0ObSct
xgXwsJRNnDG/3ly4Jx7pSAo8cJDQT2ne6sfx0YiSsGgUi+PTS0ICo8LyPadS
6dMTaoKH+7OBV67RQwg0+bwOp16ptHlkdlC/VznlZYVfbnvv22arf9o1gxDB
2mBnQFapePiCQIB5+NS48kSWvi9k86bs4LlnzXhy9/RJXMN/6oiZ1Brp5d+W
v+WgmnxMEeelSAZE2G3hTigEVLekSb2yAPKeD2MHdiY+hpNzJl/+iQgcCJzU
0q3/wXbXWrVLQBzFoI+0bSbVdAUo4RxCYdGp64itZ87YkXdWVpj/mvQte2LI
JHd+U4VRz8CWo4ajhv8YIxusTc/WxHi8DTDHBdQErfvYbU7ofmGOdH0cX2ST
fpSVpE3FLlUV+tVfjSl67qR1xwps4Q9NTgX3gFSi5NedwPvKngm4xYaMmNM5
xeM+IXxNaNjY4XnFdOCTd6Sbkmbsj2eGAiGmp401QCRHx50OXSFjEsXDLBkd
+0T4kLa+4MguE2eDfNptpGExbw0vO/2zQcDyB3qf+rHHBisEg3wfRVEeiYHv
CwKUG3bfZSDZ8gLXYPcuNAaALjXRFoBuzEWhS5z/x6WwvmEvBj9psqNlwVZ0
oowPDGyYg+t4eH4bAa0wDD0FpyUn2bLOm080F3IYPWWssFLyBP4EVO+dG9Fs
UwQ0EiBUx0AHYUHs3ggK455WWWtxX1LeUMQLoKNp0HPvI02WfhTAnST325Me
G/WLz3eG/ISk/cMJLeTEwaQuyoqyqLagylzaQAQPD1m5KqxFb548Rlc0EP3S
O0KT0ZztPKm7itzQ3NoHDkXcw6jK+tUlt79E/0F4myz1ZL3lhqpCzHWpNA34
foaCdnVxlJQ6E86vX4z+FtjjKoUdBbp3QfOZQmUtQwfR6NwQlnDfbT4wJ9Ng
htnLyC/P0ofcmoqz2Y445AL3WnCQpWctGWWZ/VNOVd7wqvPzHyr/FdBgHNDe
a9iZIhxiD9etjRFvnYC+ta5D9pBb16aj8WAAvqI3gfMZEWZthOHr1HuQ246G
NElPme3KxMRvlbCarDJp4aNQ5fa/050LxjQsmv9oVdY41CsC+3xkvLvwgS85
S14eoQ+G/laRXjxxxAKvFzi1j3OuZqWixAi6qaHDwPYT6wJGGWDFlan5QQP8
TbsAB34ttbSwv7/ofG96LH8knD9XXdglN6c+312NfScjZmmJ6g+dMXjMA8FX
vTG4qMnaQBf5RF/VlUNOvAGxP3HCObO7ygHgw44pWZVmAB0FTZAkyDge4yiN
Cq8LMylin91BVXxAti2Juur6SETBGGABy6PSTm0HYvuZvUobaPpbpKVSTgm3
hrhW3ktODcJsENqU9U2OqrZM0DaYSzhIahyLpk/Yf+HS0NpupnddDexJZbB1
UCUqgPvJlzqHrrTR0XZ9pEd0jxRObh5vkuQQLnxJOgxClYkM17kML+hLWR45
kAsogare9hXfcSU6pKkkqy5xi/U36kx9jpsW9UoFMOhV+8iIKI4snyXW8GP6
hJB63XLa+KSfqLi9dTkbapCzEMkJ1ypvABcwar4Cj9HfjYPyeyHBJLz6E9CQ
swM6JgLScJZB25uPwXCsAf9gmwiIrGLoNC/j1YsXoAfGpem/txiAVFeXWXM9
nj0h0MlwRL9sFsl7K0Qa/rch6qbiKaH4f4cYX/WesC96QZN4/95KIecqumpP
5WvZJDXtDto/j3Fod5Qb8sUmYO9RUCmeYLtj5sYnzmuNOWQMvL/AO8MAw8hg
sJMwZp+9u30Dg/bYlvCCxRkQKmVhmdSvbAZ6kFulju2HNsMGJ8cOcrJEzdXN
T3ZcD5sDDwj/ZeM10Y1NV0RDE9q3Cr7/L30kmKlosSZlU3vI0qK07gPoeywl
vFJPA5p93UPQfF4e0F3HL87Qd5+c+hraujPyHSWZbosRC8Om7NqjFO0RPmji
3egxnx+zc2dxf2HukODeM4fwybH2nDhkgNuUgwwrR1t6h9k8SJy7l+rbf6bC
YUC+/cjn9OnqMs7gfXcjdpGm9GUgiKTwAoBjYoheiwQmaCkLAfbF4rRIZZdA
+6JRFPQ+bkYcMHwbBNK8wbU6hdF8XWASgmcEgEG32Vwyjo7lAuVKquH6Yh/w
DO2i0Y5mQZVV4krMoarhKbqzacp18hJtyJxnTKBqlpovt8eoNDwhaQxXly2F
m3L6i62fEL8q8vBPu7dRyIuwZjqr/A6WNHaElzqSvrNGc8HUOzRBMlSKsqTB
Lz/rqvzI7L0ITrUF3GhH7KrfPFc40ykOobh+F6emrkQrS2qeBHPrVZ8DHXpU
jQXgFykSB3QkvFaMxzq9A39LqDYIE78ecq6x/yCWJ7mpTM4e+l6dm7xaXe33
cw7lo1GuS5KxxDbR65iQaN0DtPNrfEnK7KLopPTCT6OwO44LnFTs4Opv33+d
vUPSRkGJHBvWyINZvaT0sqaH+1acWWagz8ZVvxdGLykJUGygOYDwcl8Q0/OK
9IvzXj8z8tQbthOD+9ZIwCodMz5z9oWaVgC8Hh7044iuMyZYxxSooh48nVtm
koEaGNr2EUADqzh1ijUh1h5YrSCf6OoSsR0qtHEQGD67ZgIgOdECdSmQ8M0W
Xwsf2cIw9oxBaSMw2RpTRuQcMoRvUuPbXjnvhzHPiUOdr3DukO/rYYrUAXXb
mP7nBZwhE4umo6d72MdvBjl1xxKge6ezFL/KXY107lpGhZDIl61ndmD2oe0A
nucedS01moUrKqs/OUF+A51ll7z9kHHgIz5KFx0rI8QlUq+tLuylmNYOYyxw
jhfnbKh2NM8oxq2dpNCrLydXKhAXfxMhZv8Y0hhVSXiL94idPMItbI9uEU9I
hbflfWyMXDFEhRuU7VEL/j20zeevksGjvI9XxmW7IEfKjjz6+P96i4X19yGm
JN33pWwkjqDuqtNfHIQWzECUJ5lqRbKUEHCxO84UtatfJZxMw8NaN7RjOzho
38tLi9G4ptZdNekry90co2Yy5TIcp44Xma8yU4dosOpI9+SDL5ZbhMHJwTFp
kjk5DpKhBv3pnyKS404E4OX+S9paQ8s7XMgyplm6/E9W5pxufIP53B6kvEIP
bQw0ZeAexm9LY/A1fS+z98A8OnnZLTSwAj/t40FnHpE7LEy66OHyAM851nGp
6MU4gsBZyNc8B4fXCgHYgijipiNNquB3p0SxSt2El7oaD9jDi515H2gVi6HQ
ujRLX28IRmVOI2JJtj9uwTkFhU8oCYfo7OQDThBhYVVwwZRfiEOF7wVik3jU
b+95tLUlhJCHv7KaffkM8DtMjTT/tvU1fLfcyx1kXQ5IxrQtRqf+qCp8pc7A
wK9dbVGv11u+1vtXWvXBmgSllU++E2eCqTw/DIaE3KXOCtuhotlf9mLkymja
k+1o2jCqC2RTVzXutO0WxW4bq17MfZRcn61zjVTZK9fYvSkMaNHZfQwu9Q7Q
P3bJRgZ5zlMDM4Dd75xHQGnaN6XeY+As5Goy6YRe2v+ZGEjlkb8PzraQugls
XpXxQZqcS8igyzsL+L/XuKtYBl8HZMrJzxE43BkojmnvZOwKeIpW8LELkPvh
vzg7N1+Dur4PIZ8yoFaL6XPV9b8LJXOoVj2ER9+0PNj3hcFEPl5KwsEiECZf
6pLajhUkF8hQPqxx7AKQRPHSNfOZrVqP0xDUNh08AB5mag1za1aoiq5r6oFD
fg6VIn01Pr4XcNxmy99rj/kitVdChP62EYsclxLrBFYgtl8ImFpYzUWmh6co
Bydj/50DDtPkrxG+orUcvp9RVodUU4ij8S6wX6yRoLArYB/Bpt7tXGlG2An1
XKX6xAQ96UFdx3sQZ+6VBUiLj9vu/r7UxHEoTcJYOKk1N9j1VGS/C7mfgfIb
D65tx83wt2Pte2ZWkAY2rGaEqDFmg3+F94VcNC+BqfbLGpElbQi833VOPpms
CPtPYIngAzRvcaGpC3vBRHcinnzT4+tNyfpQNdmCGiA1VS0o9fMaYEWIWo+x
1o7sE5Yub0KQ7ig2LO2IVnbw+vDAFjQKRnw49M4XbXqLnQlraacqiLUxa7pl
eJlrEq1SmR6/TIc6xs6ZpoAgJRpk2v52CVr2styAT6QSfXpiClaQ9c26Ikts
BBQ00on4IQeiDJRtW9sOhW/2JXFGPCPdaZ/F2yrd2I7WrLt/Tsm94OzVsz3i
eWulKcIIpzyScdgt4ruEsQxeFQWsIVk8U0QoqLITQY/81QBYdoO+9rQJsGCA
s0UV8suQYgdMFEOT9Hel1qctLfY6DgscUM5bFt1Dxhe7aKUtjJT3xzJmCv8P
Eg39ZJw+JmwjaflDC7jBgSHcHsO1qo7TUQTXYYd1e/OmGicEtrdKhMLP7KKx
Yh8PgjDd/xbGbjtS7axpMw54M4ZZzSBj+CjjfJKpPTUmjhZj9nvdlX06JyD8
HJCxX1KUDezIXP4QTAvVkHRx9OqFHyWVj58HobjKnWR843JjwWALNaUsSzAc
5d8nWfudrLJCSI16sUa9Umx3Slj1oM0qv6JdZRDCAg2Ey9fBJ7KrlhyOHTia
8A10/6JncJA+BMlscVBzhnBwAAhFz6rWi7jISN0UCeb2TjJ3A34Nf0e2+aPp
G5BPb7r1onDIzyaW50PZcSCjnKxYujA7xFvBU/37S4Ni4Y90F8reSMQyzng0
NFC4OeSyCUEmcLjNEPuV/GfPxovb5MFRQE3ObHo5GnG/thm4Y2/U8p6Jzj84
PWidW7o/WlTUsC2I3/bDxM560qKfQPVtmm/HUNJ96R7him5zG21TaKdl5rWZ
IXaHCsb4i2+BXJ7fVcz6lrieTq6RqRVy4FH5yuZYSUchFkAIY2UfvgUsWJba
OPUUGSMdEchM4THmbdedd/OmVhYH83jQ9NQCuSH96Vi61XC9P4EraXl/zQct
DBtSSrP2G+CqptAvxt51ZyteL9EfJO2sZIm0CYvsjN1P/icUKothmjW3ZyMa
ElIF8eUrrhYUmySLSqOWPiBD6XQ5dFxkINBGcZyp4e/jrMSz6luZetPoZgax
lhxpfF+hRaDpEGio9KRQkoB0Q1pTutrpKMyYSGzE021ux5cFzDa/0F6+0V98
1YhIC0uvWANnznYIVQI6OHPOI52N2g7bOiWivcLx2MbN1Oy0mPOrJcwYnlF9
wmQJfrRoqXBeK7/H7oio1HO5aTeXzWJNshW8FrSCFVpSmVUprgoGUX2r5l5m
QCU/NRmZZuixeByzj3zxdeVHGhbW7ZaGwHGWlZ/p9GTurrVIsgVooKQ+MILc
IZSNLnSyYLFWvDTAk2E0ErL95Ms2bCViFyUPBS5CUsvDa5Lb7dthZvrGJeci
PSFwdEasCsrsSZy4p4hHOVJQhtju+H49+T4Ai+mboVs5uKaQwuQepYUGyVwk
DKGXzj2/Mrfjm45EDIFtpGbA21V2GvJ6se7UOPuMFswaPzmGnEFmLDxwjPjW
BmqiZbMKzC5NRqJPvNg/GcvOZ4Urz9ETvWoYa3LrUZvjS8byciZ4rYFrr9bN
dyS1ZOMkaRas/l/rAQq6zqRyA3T9Yd9oQthave5auWTpdjFYz3cnbIAhKCAq
yX3A8pA/4Cqx0pRl+eBHJGWmhuXHsKRGSp6b0Pg7CMoKf43a7WTrA4xrMms8
S9V41MrhFLMhJSskFxmTXjCeSdLC8GMc6RGglgp14YrIpVx/2WjxF5STFQt6
w2HTvJq2ievK59uADjyb5SmNwGchk8AZAVqffIjzoQ9r0QxEshmBJwfOldQz
O3HI+o+MDNdtZumEb5zgc26nb5j662EQr8IbVa0vNrtp8fgdFzcQPUPUOaM4
YSo4hJBAt/ZgbVn3BB7Z+gHiojJ1eLoEieWVhLwgomRUtP4jwenDB2t1/GfX
RUFRavKjkiI2dHOX7TK4PLaUTqnAQ/ykpUIpfWBz3GgwqsS9Nf5GoAO9vDKc
Nh2XoyPRg9fkYjVC8XTgzExrqLS0rBzue0Rg8+u2YaFrczzq4eRxgvojmYEc
GWXU1lgJv9zt6HZcFr9b0KfvnPZuC1PImYUobamJ/wmDhHWyXnJlMxrhkfkf
zPVTU3b6KmuFK/VS/HgC3qFaCiSo+Px5FLww3An2b4IAY9RskR25G8NRjOsH
jyQMWqxFXN//NPTnNUMxwXidkjr0fP9JraZ+TJqf/4dYuODlmzGi6B3d21ob
dT+zQMSZP4dTufHXbBKlEHZ4QZ5/BzgIQnQVqXwrlsul1e5ZzqoBc7gD4FPD
4VouelVhj4GvZr6oxGZRwUgwD2IY4ih6pJIe2nBOlSViA1Lnt3RtWg3pjH1G
3THEnwvtZHMWDcG9wnZMI89f07w9zQ2y46MKvskL+33VupqmK3kRSKuwdklf
qvk/jvd5VwviTsotgLA5IkywV3LCeB9/L7sqb9OSVkP23LikHKv1JU+mEfpo
YqtZFct+ypdrcTSduyRdytROa/LBYFku3kQvrzlIp7Sas70JAMPMY1irzN9f
NrcRCQpMmdqStDJlg//sqVCrpKRGQ4I2L4MlMfJ+Mp1HZJNHzlZ0nrXZUHz2
7QUtRfkCwubprsRbqFWq15vVuEO1EJU+RH4G0+EGNhiJNxlat6ycLMSEfy8A
bEC9+Os5A1bxImMbvjfHa/me1MumXws+Gr7UtR632nIae6TEkZgJBRK1m9Tc
gtS9KY7DGCgayNW+K9TFSQeuYI91EqZLSDbFlDo2pZfWkiT48t3l1kazWh6D
04XR3GyBsrmJ+jxBWm8HM5aNLMSFQFk7fvwd7Bymbt2W5URfU7fY7gLChpVw
9cIXnoe+KyL8xiiK6PSBHPriH9ciH+FVyjoreYIap5VVv6W1UscSRb41zA1U
Md4O0LjLfnLRn5ZcB0a1wumxUp5r/F7xRJ/sXRg56QYslAEslBUeAmY38JBA
598Z+8m5Ur296P/qCdFpWBIxlfSmCMoI8zkdQERvyrTx+TF0qvUjZhwnz7pf
3BvfEFL15Ge5d5qNoEymS3CVcuKiEdYjg2Gq9i6+VUno8u4lPG6+u4Xk1gwd
f3PSc3I0eIbt9oLYl2WMuX8bl5tb6n88ozikxzBwVeVYh48TWD4tKNyNXrZk
3EeV4/uxgMrt3VkTz31NkEL8qwzYKDH3Y7ybiZY5zQByG3GrJQaql5MU85Ks
APR6ABZh2G0vJmyHQ/NdbtjQoI1vWRkr44FZc2RDyywoULcuEDX8xLkkQAtH
X/Cwd1IUxcbV4OlA9ZRX8XUxB4IWxwJIi84U9iNdazZsGbQooMgV92mlmFai
wdzYZ+9ANrru0z1LU/aQa9QGYTeRK0lFOAyc7peLS20JVHD2KL+TIeDalLsm
mRKlKQbqlrIB9mStsKcIxdT1xXplne096opQlHupL0/4BranO++3m6na3CNb
xVh5fEOSVZv7n9BKXp+plgRHwgnfYOSBuNcP07ApUQjywL3nFYHz5XePkRjb
HgEYSUfqpBM9BpYegnpf+12PDhG9WltJlrs2HuFzDUd/qmUMxCXso7KbsmsR
qV0yAVs+U/rxH0EMsspxaFEh4ALQ5otDF5KSU8qZwFPIBkBoQ0VqAHGY48IH
cy94n+OpFS2TK7KT5nOxAS5rukHvPrtqdun3glFglppiKDAmDRQezDfHAz+m
Dd21UvaGQcCu/aAQ4soEvFiKAPFhn/GxaFAbYjpQlFaYHjoAQzDvhVV4aTHB
cNIXncuMEQ9gtm7Syzd3KE2EgUjaGwyq6PIxmQ/4YqwsM7onxUi7UGHd5ZBQ
z+cuKBncngM78KpR9lY94z1OnaLSOoufx8CUZtHF3U+JOfpRPd3RslITF8Mz
w9R5H8EDyduAO9xDGDBG3RNu5j+f79Q9T3nzY4Z4c88zdZEfO2KAa61wi/u6
fxNzAKC2U+NTMW4pgVWf2zTdmnoqteCXUAICP9zP6IU6d8N1OHdBNoQlUVhb
bMFItIwcvwfafOy9uZyRO6FkmXrkLqrVT+z+nA7kXfUP8BDq5ETRBO6FnwWn
959AyGonuAM+KlTnnSpu6YXCrI3zMPTFZT6+cu8GfnbILPkyvktxt/hl6Cq8
UB1gLyi6H2dCgRiEP8IxrZpPi7ESjw3kfshuKRXp5mx0ymm57caEC4V6x6uQ
7PpCn9r9VSBNon17sGZ3kes90xHlEQ4oOz3ijP2MCXevZ5Wk/vKQeuG5EFlg
UbuKYmKtpdmTEj/ym1v4siZJ9U/uULkADVdeQfyA7L3nKF5FXa5O++cYkSGM
19AQnPzriw7Sg0NzhtSAkYItQrLhu+DEVZUi/877ypv+IcjOR4vo50w0dCjq
En5kLy74NzIy+sO01gSasq5z1T29HLFvLUIvXWymuW+FaB8vM58/DH1rwY7x
3LaNL7IMHTUCk3R4uqTqqVEd/MYf09QCcX5+7xgz80p447QkwzvkfJee+aCQ
r86WNoUwYszXLBxlrDclkNzYUezQbX5EDj0CNLHPU00QBX9/vFn+e4mUkHcd
kaqhtM2/w5e2VMot5w4D4422ydhIKbxEGPtvSm4WGZcNqQA2G97GzCMYuEQ3
JoSjLRSj0KCBll0wT8pmk9ItTalNRYjtflGwLFuuPNtvlYk4aQidJNYONvw8
fjJ1l8GdJpPR3mwaQTd0zpAHfwo99A/9o7kz/32ZkyMABkHH2X5dzrW7SY3Y
Zwv/fqQfOX0s1QZMxPcXUCl65KV4T+yFOxWN9r77q/BFQc671xt+i8dlTmpV
G6fq3yen69Jg+DggA10wip7/yWf4sx3FzJ93hrCGNaVuOfNcYYeFr0bwFOVp
/secRxxK5Stu2/pq/3gJwP16wSLPo21IK+r44vts8Z+Tk1njT3fszwa+6J24
/56h8IBWVnswFX5h4d9lHJ4xn2ke/Ua4Y1C8T1fbqrxfsn9VFAYHFP7q4uqT
IhWMlqRoFXgbpjvCF4ABO9f8HmFDzDPa7CtNmyiUJ+RH6fqbUiRu/qSvzYam
mzLDt/Llie003wLUpzpQbY0pzZPdNt8zmGlXIopID4Ucn8GdaNWUoXyPMh+o
PozmZA6R2T/yoG4JJrfDSiV1U6i9Y1+LxNOHeHLEswvRhJVgwR3BY8zwnxUd
Cg+uKLgp3QPh2pS/pM8m/p/QyrCFk4izmxBdiWYDgFMu4TpEwypLj3E/DWGx
2nIbLR1f+9B0orPF7Fwh7yqO3YlGgPeYbXBk3hnCvFOW2hUOebjy3ZKGleoE
Fi5h5AvECODGNDcrbR/WHWA19aC4BfXjUlkdr5FevY3+8Tyk/x6Lzf9Z2S02
xOZaX0mKwBwEkvoUkGAmVtYnwbLqeQT4Iyv4SN9BHA88u/FH1WZWxC2TFa9V
oHmJq+rfy/metZBYIYVPZ6HYI70HvYG5Ta4vrWfiVr+hqhK/TfudQ9tQ5fRH
BM8B8+MCmTA8TsFlqLrnadEW/wVkP3hnniA08IklvD3hGMYZGFwSXDN3xHmC
UxkDiU8+0L3HACiCRZSo6deTlst7RkPiht9Dm0GgE6jEi/FropY8e1P+46Z+
zDPbxG00nZ/SQud96hi9wqAEK6rwXwIpG/FPsRxeJMSAMTwobgUHbL/avw1b
RAJ7YLuI+r8KKQCohTU3/7Zbbd7jwqCnbf8LnNqkjNoOR4rVAWJpxRL9Jso+
E1+l8eoIEgXZsy94UOonXToHo0b6IkBkq/M1vhcRcz6fdfqyPOKjoBpv4Rvg
Sr0xxolXtjzsYBUW/yiBbtCGZBp2qq5TJcA1KN2XJ5p5sRb8KoyzHLeneASU
bWqrsoao2nZ8OJkPBEN6XiEnkKA+EPoa7X60cxWwTbS58RvYGskFft103C0n
U9ubt5tYqRP/u858ZqHMlXrd4PZJpldy5sLBnUApIsNpq7vW17DMmTmDfWHp
XplCfI/DAE3gJlhL2qyA9Bxwf190Cj9hXhpxuMPxrCfD/1XzxGhnfF/wFTgT
rRapSgrs9sRdeltwiG793++I07dTOgG/TrOBDGOb1P8QLt8qNjG5vzmpA8IU
cmldeCQIiCncCu+8/gbgYgIpjjoVdy7FN/Hh7P4oN++VAK4UyUqCty89dzof
8xa/KvlF0lW09GzTb5hRTOSIXBKiGSPu3BvfyEj5o24h4mEYPOtUcOqES8zb
E1APYHZjsqH7TR3Mqa9TEqonFF90B8gYOXTf8rkl3g2UgAVMBRaGYvkcA+ST
/R19FGwmTBWoYJFzwCFUFW27ADJaVvHBNVAbZNSL1yKBhW4mnbMAybEi1rNB
3gAyIZvwYnEz60hT3pA7x74DgigyHahpdaOFvnK43EREydSejClwC16m2Bx9
XgYWG+iLQgk29SbKqLLe07MrzJE0t/SyRkPQ6AxlBsVbGo5JQeMTSguJOVk8
+vkfjTv1lUY+Nec8BVp/gdLuL1MnkAPM0MXEGm4haEEyXPuqJzCMUd7B250U
t36o4wj+A/RGc/dSg9OVzTmAoMjyRgRZ7NsF8g0+Fm9FPynf7nRKpOTgSgbW
Vwzi2sBSZc3XwaaM7mwJs8Bugg1Pnab6W1ARYzCC3N06s0nqyUpXdbPOAjAR
cowrUZP4ZP7+IIrXJCpho2k+GRl3FHhph2Ao9vM1YKwYu93WivkZP+zSr4YP
YeNXOeYdlRY/YaFxs0bOxnxPea8AfzminvW8GsPHUGnsOtwCNOPZdHQhnVnK
FAhGlCOJMDnpZL4+clpm43mgEko5lo9ZNra0be4VhgAWTgAET3sjVKK5Vgcs
AzhMQPrV/LfqPIh87BF/WQX+/c89ieaCmi9qu0NKUQlhLAzhNI/CF4auHcMr
CmR21dB3qtrJ5A0OTYo2kqFhs0Kg7LFkQgeg8fwVjfSINtM5hWUq69VZaFt3
daoHGTY2sFvIPdN19MSrgio3lq/wzB2GOgPtDYts67WiTQOPUeSiaZla1EFG
j7SwkHzNyUO96Jyuim9638OhhglfnKRF8xLI5It8pZUae4W4G0W2DTP+plsx
bH5wPXrluvoJ4eTBdXNWTb/Idg1InYZYAhPFkaFKuX+hjawdikr9UCojRAqF
mOjmQQKmR0/wqL83vNtLR3SxjWwy/msFPsmpB59phlKjbKXQ38exSMZD1o0/
xM3KXe5W3Uxfi7zNCbwWSRBebLyE0dJYEWoRgxQ+bsQqxAzjo15D2oSq6yVN
YNxeJuM/32frBSVBE/dvpKGs5d8H66Sfv6+pV11jjAoX2AOmMc3MDXfZID7B
DqhP3pM3v7FEonETjQDHfDcZeExpnWL+STHAsb0nIt0bWn5q/1oL5AkBwlcH
6JBjqFIkjU77UhuKuvlNj19wH0yGlhKbJDMRObLsi2R68aggr/qf+/uRPedg
Vh9SXlOLpXTJ4NWoXDsJBMIUo9EGr45s2KyF8+eszX3TyQ8aI0KMuriF3Hvk
lfg7vOiE9T5anMoOMjEbq2zFBQbfb69dZkwFoKLbEzcEMy3mxxGP0xOOVS/p
XWfGIdvk5cgiIqs/MhD+B/oj/FckVM2374ZUO+4P4pDh6ZttFv3qARmZWk9B
YdCx3I7zhy8QkAXoPIjday80nt0yiiCMXnVIkXErazEYSxTkSBxrnY2EgTw2
jFKFCCDLU59fxchiLnaSvRq0P8AQy9ajO2Eb3cgE4bcadbd1IfXfiEEqJh8Z
4cKpHMx1whfFsdHQkgoR56X1vYMLNU72A9yFHyOq3nXvl7/EnONd+++8ma+l
SwS9uw1c8spESrkNRGoWmAYj6WfFjXf7Tv2Thsrj4j61JtyK+Hy0hpxfiQDv
UgUkNSs5W1pvDHlnV+dKlJKokXIZAvg/XHAWfis+S5wEnFt8t4FX8uFr4mEn
Pz8fPLc5lVSPVctDdO19dm4CrKS54sDkG//Orf9gGUsMLnLZLeNs0rzQcsk9
ayOPx1Ys/Wch1YKwH8hV+X7JMNeNngHTx9ZL4C1bSpjFrTu77L94yN/oe6+i
9fNudcdfdSx8mERE5i3yc9Tcxydsit76xCv2qer9PtC8Niv+iXnySlmPBbD6
YVSje6hUdPX5veGl6X4xU1SiivtUxP5Y09UQJSILiG3vZwbtMmM7ll+CDF35
oClo51wSnFnjcX+dDEApK4taNLfd1u4ta4HzDeMLmkQuF4xXSFqeThodze7u
Duv+gkUdcVIfCI7ChNEQ47/waAC4xBsegVZru5R1JUxZz89uqg0UA4w/uYVZ
JvwzztBoFm6PVgme8ostKNRzmhEhgFAHoBqgTTqE2PG3PCT09itBYIcMLiIy
2ksvqrAMqTBq9MYp0FIptLJCvwoFdzYQLtKzkeOR/ZjKz+ckPfVkPenO+CjX
2HAT6X7t1nv1gjqZi86i+BGirBlFGS6Mharcwktp7ofrLpgaDiKvXhGwRupO
7Q0kS7EePAdZBdIeNKFisUyojZhJWQuBuK0dky1wcVO0TxHwlY19gplL3C5F
UvzyqYWo3aVRh/DJqIRZR6YneipWANFlvUBXpA9QzShzACrSEQgRNzKLvF2O
WXMLeYgBQnM1cyYkqy+1t6OCyxYPUSGR3Q40jpfFDxM+Wd8W86cliRHVTanD
B6Psy0ZjrJYS+1M3//fWmrxer8cqgAYSWBJ2CyCxoJ3k82NDtrP2KC14h+BC
19t51EWNitgVRp7atJixMEkyeAgwcJUamdNhYc0AA2JRm244nR++vFuqMJHL
a7WsTUxVGnOVmiYpBcwfvJvUG0PQSkf28qE7S0ajZ+7M8IBJG/9YwpTgJv01
qd55sAUznGjC5m1GgwzZUn7izX1jGZ1mCmLVb58B+pPmxsVyKplwL+BIxO1o
mHBtPoF4RKFzyAg/YPt4upfHyOO2ueQPuxbdd8OsyvN6ayNEauNMIAaarvbu
hdjPRwYL9Il0Zat1ixVyYGEBjqGQoJhpEKOnEW3h/MjqVU3/1Y+CQXpgfIEl
ypb+FzmLtHotfRZtQetC2M8lSW4SdYD8i7FK3M7JObXoDN24qPUzPMWBfPlj
GlX6ReXQoUIYD9e/1JhTc20uAuowDxCxME/tfHKmJmvEDvTViIu6m9oceRea
p/cdUw3chI9N9Y+PIsUWgWmgRZPE8OU7L93JGdZ3O2V6j3M3UYr1tSKSclNb
1w53zI44SMhBJRxMmOeABKjEtuS+ENpKCKrabHkpX4hqSA3Kf4T2gSNksdP1
4lJ8AKP4oQvjORFV4ZlRBAPB+fdNdB906dhIRMTPlJoLgm1N+HdyC6nFBSgv
Cnf6TS9G3QDKxXl8oJ+d5nkgBG2HS/P/AqX1AqhqQAAGPgbNOSAN05RW1Ih0
W1Qe/0k3nXWMQAxV3B2KpVggM8P1CBqEVoaZEW2Pug7V2l0HNbwgGbm7/WfI
SLKqwdfiuvswmYaRGLPudw6pcQUkjoaYJoYIG3UUjJ9nZ9QddUMoKZke6xNW
ie+n7uOBByGCQGDCarmhwBBXLIwlqUBs5lUebVpRy5/ZU3/yLhOzuO7S2Ue7
RNFQbaicf/ZqV/GszwucDedIdqhTjpE8eJL0o/3MzaJQboNoNFvOY8L57/iE
PiusnCgaT94lp9cau5D7f7rsu8f4crFdPWz1fGWj0WcahFylaXwdZnJIyJ8x
WnCZzFaZ+JM1YILSHIJ3nqfJi6vnmai/7kUgkWQtS+dkBYqupLGHED3ELDcY
NqKzZY7TVrrY4tyEm1ttfoBgMYfX4dFSuQ8frDBHb5dygN0sZunXiHSVTb6i
IR7w5t/t1qAYs4QMeSoEtfXTR/zNoMdeeHv7AMDicj4fMegOOzSsHJSQAGdo
1Amdr3UI1jTt4ua+Ip5iq+SLnKrbyUVej30WdlyvHAwYR603v3zqN5fitBAe
WMo3jRj6Irc5RexKI9H+94kxTo9+rUYLTGIOxaHkwpURZwtWAF8QlELKbQ9C
CIYKpt4kt4hjTn3NhtBtIcREXj0n2t91rG0wO6VmQsv3m6FvJFujakGsOYpY
bam1Y4u+7U5FaL8oLaNgA/WSbULTNh7Hkm4eE7VR569yVn1taslMYcHZWzyA
WI1SQ9RC/UZ5N/mH7l2OokKJY9p/B0S5nfiV2UfGhjCOv5P8zpJy1wu/bbZt
2bTvsJcMo3u3A29lvIqM0RylT/nkpeaeEuVFqS+AGj2xniXJXVTJ3/4xzgkR
tJHeG576xJrQ9nhggRb03SuDILWOMn70gBpQNHwZZePRVvnEh7qH+63H80qy
uqtKv7OIbaPKYI4qGLbfeLda3UjDR/qOrOqeeLG7C39XiTkkzmIbmd6Bsj75
JIluEXLm+RzZzwdbX7M4hHtoTEyAQ61cdJVz6FikHzRm/hB3gsDl0ZyLFDT3
BwGGUbMNuFrC40tbxaVerViBx9NhzSWJbX1Z3sqft8FpbGQ8zrrcnWesK2Av
gq6Qnei55wTyNZ4moJkKOiGoigLOw/JAyuN+1hYw4CIlrW8oQ/L9VRYh2zn4
Scf0WoTfir64t5UwaIXjj9oXiEf6qzZDtjl0iBr1rS2Kw5V/1nASt8fP3tK0
LFd71iV8v2LqaGhRV+mAveXK22iZMgKKGZyTyALEWFSOmziIjjtDIYc8j1VW
gOtDDV7Vz1H32iinfzg1qmkd6hrZKscNrY2uTS10XMfgZzF0Psben2uN72i7
KRpWNFV8jAHxdtH5FDW4bN/6BPpxrCp7KFRAYHKqHaa1eR69GOqiNG3hpo+8
9UVgBO5hgHAQ3DGhDmM2VPAjLGu+oE5nu0aRM2VwdYJxH+0FDMW5mK2adfJy
UoinbbA48hUJ+MeAINZ+awgs9GOu2fLAcJFj1XxmbgbokumtgTiN7T7xQuZq
MOCvZL65gXzSryhzoHtxQOH+Pr4IN2w9nsZ06pvT5Su1OypCUpxPQlo3x5g1
F8CNowlqjp5tJNf5YNTXjAdqqvp4G6FLUo0xLjPIKZc/bCQHbCec9FGH2b1q
4aGgnuSNehjrb3CXY2BMf7gjXM0xWDGL8NXHRzWXHcv/4ZhFl8hwUD/wv6YY
5TGlTdcDaxG2B+380BLqNYIGiCYf9BjzjZGkKdC/KJEpZrYCyo2IFC0I2C8W
pcj18D/zY+Z+sX+mJQL4E6Hzl4XlUwrhWEn7e9mfoNouAMobD8QduoB4Ko3Q
CTEhU/pk68oHlj4kuXZGF62c5ejjcBVV+WWVzOLkqnKuJGdpy0ZSxHcmKgYU
oJIHYhPBAKBohjzj+juGLGoIs/6omqwLcGhN0VBzKTfPae1x4IjgOukm3qTJ
ecHI8aM83V7mfVCMcFK9D77Btf7Ba3d71FDwc5KRAYxHYgiJ0VlQuRc1U/hq
wWXWoVbl1eKMAUXm30Rvr3nNFgGB2bVmKkuueLTHWkweDqkD6A4QIcdQY5Nq
mltT6lU3OxasZu4tp37Vbeu3APCLpD529BbFz2li/qfePLNm+qeAcrmD/NxE
4SVscsQV/Nhz868//VVcm6OB9qfrspVPnm8Pibn07MVVN3qGT3Ar+hvyekvh
p+NRj2HuoJcRC0bYZg/T1GkFOBPhhoobn79qHvh7VTyciIfrwO5T5QH1pndB
D2+O//RFmcEpmKvwCV1oBsXx1N0WW2ow4zLq0ocaQ+vb5NDt5xtUL+BYEvbq
2XQxB0MH9z5aNIMeVH+lgsInZdZD+Wod6wWIegbxc4Iucp9q3b3WvPpv48pd
xmEA3wN+5vbpCMo4awzhIYLedkTBWFLvqO/NFuFCPWAmysxed90Sk4qV8dya
O8TPWS1HP/r492kR/D2jvQ2/K/HjjB4CBgF9t6zs132UMeBqQHj3IFviY8PQ
3yL5F82IpjZNGklzr9ookbbGrdB5+AV02f+Yqu6vetUalMINn8Om3AJyybEn
BeS2RfOQyQOENd2ThX3Iut/m2YuibueGgtgQrz8Rt577tUfqH9Z7XrwCKpRn
uJLHjCN1HLPt8m0vG6+2Q9Lczj0OgMNFrb3K02Tq8vt0kgP0i/B+6AtiB7HC
Qjp2eZAHKktsviEwLPJRRIqJ76Eu5kogduiCaDp/UEnFrNsRAnmrbIhXjJPU
3dEh8TLg6OXEnlXQQYD2hyCA+7aDgqar2jG3oAseG7/pQxAxFVGMG58ix+Pu
9YE8hgVmidhQZcLxojcbfI6rcdOdsPhOYQ6/EFpGDTOzhWclb4OJFY6GaTkn
I5vfhVWBlfTPhL6rh33v8jPG/X7FxADGgz1aS4O5euNNYSrEpbQWdWYE5rHx
dZ3LnJ+K7RykhETgsjG6t7jQIRlfAIMk1Xnwu/uYAF6jFSAHX4Jzq8t102wy
l8CTLpdPFNikZFZZnOZzuqWd684ri506unI8EkdYLofvbP+WX1U83d0evxy5
akgH4Z6Vbc0wZkYl1QMRXm8a47FHEoC1Yl/QmDi0Hprdr2SfBkObDuzxCJEE
56TT4YT13+8ra7SuK1FgUCdU1QFFO5A0b98ou2pEMPdK1ZklS5tG2UJdhmvD
EAKToMIHafWiUG8OkOpH1iuhY0bS6H+mjsQIZ9FKPFRdaXKUOlCwv/yL0uQJ
+DvRIMcIm4lv4tuuKJmMGpOAUShllZ7GHWTdgVf2ib89VRxnsGf86TLAJR5d
ilajdV4H9c8WCpvbNcR57nln+KEpSO0h6BB5pvQQxNm20pkgjNDZmV/nqTWo
RZLs8LR5TNfWyda71NmBIn/FKo4SHwv+UQEQnZ2l3h7cu6WQ7TVdsHXPtuYV
uHZzFSAd45LhMKHagFtl9fNLRmgYTOBYOlXJF3vXLhghhwhfe7bhCcJg/ldi
HDGrImgOSLcy0shqeBMCdO9/XriRHvpqCM472CfjIEsWQ5tkOZOgIocMzlbh
P2sarX4IYPWQ13kMwRl8rS/IPyLhl6mRfRx6RKUOep/Qh+4mk69SoXrvJGm/
tW7SPvLgDxbm0GPXrkn6GMOhFMoLFEnZ1Q4rUOD+XPIW+T5zkG6K6I8GEd6k
E7WMMKQXjHH5Dqo+LtzA2yeZhRkzWSqKSTyUzYUu/6DK5gYzMIFqNDOyC/DM
MBn13bPZqTvLw4Hnc43f3plOaPlOV+SIlP07P3MyJ4zE+60usP6yA3si/pF4
9WjcPZjyu3FbFu0x4k7aNJl8EemFA2tCLRtnSE+daaAEZi+wD6mIGQRmXp+k
dqBEWjKBYbiB9wrhvW4D5y3ON7YRbhvlOf2B/FPhK4iOQkH9ERsN7O2J/PIs
W8trF8Lg3R3/641+zlLeM6lR9PExWyYb+2Lnk9t8nfz+1l5IIUfkO36jzMom
4MEJAp/vdMy+pNApBxXpf+qo6X364q6nLePI0a1Y4CXWYsgCcm3xUDGVPWi7
VnO3jpD/j1iVpMxhlAKsPOEFWL2XOi76GzFDRVKysrhHrE09aNkt90VNMHOd
7NGRNaH8mRs6cZh5FRY7tNwyJZRATHvXwaZgF5lIVpHGMMtjq9W1Xtd2hx5+
2vcbsXr2Wo4Pj7AGzG3a6ASRbc0aLc+vBtvPg7KiOmD8FPMpBwUb5vFXa1EQ
SAJZmKHLxmSKnqEdkvC3CN0lXXJSKgRmWOxD3IYEK2CEM3SkN/X7b4zBqdib
yP/Ja4D/h6HMesczPCkH0eSHkNCdtNUiGclh6PdgIgom9f3cCe9yj9c/faGa
1nA1fKulZEoapN2HzD5AeSBlQnKeIoRFSY4PwmA7vZf87yd0JPaufrb5a+EH
9/Bf0x0sFSQRzg+b8DTcpSz71Z+Ev/HF5eCcV6b7euZRrBvnp08VElH3n3jF
7QpLpusW0vOUf52LIXVFa8h1JcURfvmmZz+XO2TNvhuXCB/jHPQufBea6+EU
eHy3WtUsqCYZF2j3+JynlGX05MJJDb85hK0FcWQ17F1wEVN38SP//TsCC6Gc
1026CzsN+q30WrVpCg92LjMubUOB1OgEpPyBcPkcszX05spWBVdU1UlqLmHj
nTyr1WHXvXPpNyMWV0GoCWIMYprfz+NidKJrESzZIVQJXZ5So3XrcbI62KmH
DnNAm+B6/V8smXoGhWyJ1xNm8wHcy94Uu0qs+VYxXVpnybiEbPmywYcqDZVp
B0K2BpHKVtGjHT2Ve6fOc43Ly5uVaaA4EyrAGUYYS1qcOtxqxv78iq3dip5o
nMLgrgvVP6q1ApcJluKZjW12Dwc40/ZBeZv1wfobFEmt+COaGywqwL0e9jFT
c9JctVxkGi4f7ydUao+jQn4zlgFN1XLJg1th7xdwTPoXuXQm999gmfG+Fg5D
XKGHC+QVU231qwtCnS32D7EpzALGT1irsCfH/rrruhSgtj4qZdQxfMkwobL/
qRCPKl/x3j8WsUxj8mEnJYw8vp/GvTXHRoDX1xgoKJYz7emzmuz+BNEuwwHf
ahiVcR+XAhuwTwVI/XPCvHO1KIEI2l+rJG6Zr5mbuY9PXk8MoVxbJ7vJIE8x
1rfkWWHTQwjCkHv/ldhPI7+J9u9cuomKYGi46BNQ+3S8ZTvBqfhihFE1Ouam
JPCoYH+idZ64ebqHpLyVnftFPe/bmeBtEeGnkkiZj/WPI8bEFYkMNx6jLvFi
Z6H510KZ61SRjhz1IQ6jahjA8b+0H6uEJuW0N4kVsEsD2obZXXALX1fSYBeG
OUq/Jehp8R7qLWaXVgYiIv3uB4cViQ2OOqdSSquBuZ+Oo3GMdvrkZJ4425xH
TAyKnGYtU6shI2atUmDE3YB+wbm6ND1aEllhg7XKYdQJSw68xATJxHTwDtGv
LJkjlnwEnJSAXPYdPdEapR3dhfk9ajeY0shCF7MR7gz6o+/5wCgtUn55hyoQ
x4iacOAuyC0SYwprmLm32vHqTz1/GoxeuikmBrOlWHBiQ2EYdTsP+wJqzcmR
iPVOYF3YX5Ya+bXTgYYCG7m2b6ACczVdY8MRrQqF4oIL2UVFN5DdcDPdF11m
qVYkuSdZtV8f71OUQFy4g0Z16sCYdYCFEnrV9gGXgPVl2coAAZY8FLtSZW4+
R3EyX07OY3Cv5nba/rKZeNpew7omsi+E7mzgs8Flb440f2qwMuonIqoBYisk
xH06zaepjlZEjNfSKN3zkAWUsI4OyLRA310dXPt2W8w1Nlc5LjyX+uukZnEW
UL/1OflJxnEP2t/tbAgdnrjq0p3ozbU0DeHIeWWUhtq6Ycbgk2MyVtyeuQ0p
rRpB/FX1aV+Bi843mf/Iq5Hz9GgRr8ilDoY4KYoOEmbP0HFF+Cw11P8YtJrx
iijXjgblm0Evt5MfioPlikCQSPomrRDQ/bFQknvv6fd5C1WNXHi+jur7iulP
5rbUaz1OBRJ3o1cHOA2rfp0n7USJp4AbJO72cpr/aXC/QudsCLnkasz8OPHJ
b2PWZZVzaOjeTTt32M5/cAy2dPJi8K2pNY0HnXYQWreOo5g2LEBitC/sCRab
JG4v65hRdthqP36g4/yzrsyUKI41l8/mpZxb2W3NmZZ6Fly5zqiNxbqQhi1w
FSnQD5lzuSRWhbOjsWockXl6stjkomdH1qU0ewuObUlGXfwSCBMRtQOKRcZ7
4UId/7XqAmWoVB+5ZCnbmK8moPABh6cjN4QpJpGuqqhtx+TqpUW48uZ2DWgy
PLx540JcAkFwgZAfJL0ZLXVOj42LiMFXDDK2k+9f+HAxaDd+fXae5skAPx+Y
fV0wOISz1G1js3GVGECHgdLE0OjUbrTJf7XLr0clqqOI1m22UVQVHkm+YEgV
2bPOvuO4scZ+63Oe03uZnw8GvuxUfNTkCodvx/R1uTCHjMFG1MhJC0NGMGrC
etVxMeymUvPqheykFSkfdpVzGirZavCoNSl1bBlORH2Ft+am/xsLqkV69Kqy
3UOzNJd1Dkkpg7Tws8HE6FojDvLgzckX1FCw1lbag4vkM/d1rkQGYh0gDUAO
SOfPSJlMurs0cDUt9XFzybTMv2NpWRCXx085r/D7qA7REWCbEJp3oGLSZkO9
ADCRnw2D6JGnj+pnYH08XrcO/zvz+R9kOBw5TyXhUrzR+wBozsWdGpk0Pgtp
2g7ZMcFKfq8Gla9dvZhKXRe1Efl1gUTSZVj7v4zlQ6T3IRcl2TZTs+wZSyT4
mxl73l0JPU8G70t2D5++35Fn+gu4gUzWwjsjPi9SipeYfxou1CC5FEeV3C/F
VcXCt0zRBWNu2ZjNLDN1wFUQtGipzv9I8Aw5u70tTxELBhEdd1WGgDgn8D88
u64noxRtVfrHrM61h5R3E6381U/xmU660WN1XkuV6StcLJJHKdyQuYf66WZH
tmN/fW43C6H0CknxA8SKMloTW1tI4XNnWrXKDE9YVMW/ENqRkEnPHdTsUlOM
iZOeB3nfPVoNybmseW+ZYGZbsfko9+Xhy5MrFUFf+VWywmjBnSYcfnZezV8Q
5vKokibjG7vyZfyH6lOUa7Yo9DA+kwiYqovW1ZaHlLGr/pgh3ov16eLDCZKc
mBteFyva2c+VELOtHP5jkp3hbjMzIZVYaw9jIDOuDmXSKx9ym5XG7ZFxVPF7
qQAjTKQcdRCGYive5LspCKvrX1TYw/WU5XXNn2117njeHd1YM7jZv+11LpWn
5ef8Bqcl5C04zHHJe9lf/L5CT/+58iiE9Rd+evZRDy0M1mBl2llFP1G+RhpI
AIPVg0ki3R2nFdKwK4xqdDEUwRbpo3Mo9SzHHsmcs2M/z5lnoRMu5MtM93/I
fFEWCxkHUiTGeji8g+lqODdGVNQVFLq2WaLuKqyq3052NSXkN6WukLsyX6Ih
Po6KjXhSz3ugx7I1t0bEQ0bqkK3ER4zWQVu101+NUuAVh7IaOv+6lkZ9q7MZ
EmFu7yG7sBx8o9fvfcxTKuJpdngtH/pS22449jOXkBmh3ct0nKpKyFpvjOFN
bYRDH/Bu3Q8kLGuepciNj5p69aqnVRAc+StSgC2uHObu5sP0v4KXCtS8oUU2
LyedZ9kS2nwPhd03GAmoR3ffNPjAbFLu8LdC8EZlUbJtzuVnw/FXvk6nokeu
HE2xiJBoRMNvrCipbRnWrtmr7EsEyY9cYJzx/TPGCtX2Zoxj//t1sn5ieFb5
jXfRe7sj0AoDWFHzrEJvbJqFE6RBxdx2bxfieJUddWTbyvZlRpD7LmAv79xy
KKKoCzj2WdIaM8msZvpg9ME10XEnLO+XUNk9tjlXsXiPo77PbHlTE3s3cn9x
DVVV/9Aw8RJniql5nsFk1WfKKnQJfBPkbejUwEb3S8Qt5lUPhBzWQTWP0Kd8
VDmG89aschRhubfyyaffxG7lISwdZne7FaGXhqa4JWqYQoUKRFs2ND84wWSn
GWQzDlxhar1mQPTRrNi0ms/FXXj6/AqMSlYPdYsLgFt6CzIFZjhXUnDsQ94D
URjtcthac8cjeRODvFz7ZR7nnsps0I0Lys7dIOg7kF+UjjnjG5OOj8J7wTkl
1bYFEvs8B5U86EL4Nm3faixAsZexUHaHU4nrbxw5iLgiQlXjJkuMPJkczeqz
ELEJ2TOuKoJY0N5SsKmrY6tVdTdA2zU4FP1rMZFzIg8L4lsbwR3fv2L2+fp+
CK+kAR5DXosy65clwdU/mgnZweM8DRxjfS4WR+M6qyDjeDpFF2NrRYq8RQiB
pc/I9ok0StuAcMnCg+ey6S0f9xQY0V+RETpjJBDzSP8ONL6g5/hMAcLEghZx
o+8fYqk2bGbrCM3GJTh3phlwno/OW/72UtA3bQi9Z3SZiXx+f4WvFSDSprH3
0W4RWp+yJzLI9CtGNfZJukyPdfN3aL/4lr1/vePY1xJ4bXdjo+thwTVnRAjk
97zcIBSljIlZCSw0JBcqvcR6EACQAhX0L6XWYmPKeyaPmj3wj7tWAjsWTfJJ
MJqO3Y9ntvZqYmPLrJtUaHdiwxY7F/RD7jLtgNLKgzJr0SUsO500M0uNTlk4
p1IO43yEuEiTqqs9QCxmQq1kAj6zK26f2IfZ1Y7s2So8IJMJq2iNibrKgWqD
R6V93z+L/dbQVdQVXYcv4Vc06/au75gpVo5vdK7+WRP3S1X+Zgg7xDmz2uvJ
Qq42WAsthJLg8koIGrNXoeln3TX+16/ks0wZ2NyRAZcU+InUuZAgNEgjPLVF
Q97Y2jtQSaQJRvhfxNgdeLivlbZ1NY94V4RoSjZGVZ3HxFr08uddwvyNj0oZ
SJA2R8wRvS8UhdGU+PZWBI6ZXdBzImOXVB4ZoI2U/tzi9+iqrvCNw3Ule4Mq
zzvS8Q2U622kQRxvTb97z63DDbbQhj8lTbkvkdTlnywPLLTl7/pZXnHmIYK7
SX6AwlBPKcDUm43Sk94TcNNDnlWBLvct0fItxEZSSwqq7EsZZoU2hnudnCoM
GWYjSAHh7KfhKzrgjSG3Q5lqqdJIejAlajKsY0eaJlK1eELJ5i3pTekcCEZ0
uVYGnhB/4qYHfHrH1bPP1UoTgN/yIatVfSCuk3L//FnFiAXUtPJQbeF43vMU
F58OUU/+lmyAfKMU1eHHVMDS90lzWUJnlB/gnYvuwos8Vm7JiDcDIX/EH/G8
KFB+ozS10PQLl5OG2ES2F48mXynsbQogJ113k1QtCyo9DY0VpLBkicqPrEcS
ld6hJ68wusaRRj9kXtn4GhOaHLadn15r9vrogGg7yIOSGm7y34DYrEwTl/Gb
krV3BG8Q/nYRArAqZqqnyY2tpCpfxQvrx2U6fKty/Jkaa79Id0L/UIKeBR/y
q2XuaFNmK5U8qRFjiwS2zD33G0mKfJ04wbW4TBN7xU3w7L9+dCfHn2ypZ35v
0t4AotZ2maT1CvLYy9N6uRO/LpxpP/GRkAKI1YxSEIFV4rs5uph5CeJYnimk
yiuy/iHaiJwnzTrUuVwF97wE55dpbbQfHunWlpZhkxrDaWtJRRS+9lTkHJg+
ltDnhV+hFKzrMfV+Kp3Pi5z7HkS342wxGreITKWH+3yS5dsFSdZ4nmVjk2ZO
2dSQGvpUlXEuyYKMfHvaWEoO+2YTASKK5I0kTjIYmUBRHkrv6eGp1vD3Ypm+
/gwBLM2AXFgMAiKr335/J7lRGW4c1uLtxRNAT8cNYgB49KaluyZuJWzwscwF
VYvTENe/QZ8rLVOWWBEn3FFifu/+4Rkk/SYGRYP7ARItUF+U5cdECOBK+ZTQ
tlPUFgl73Wi8znFX7AucHNb1/dISSSBlQdg0Ngw3VugpG3e2Mb0omdbo/ctg
LHVB0o+DWp/K3nKA6bmWgdN6irLLvZ6apduV1nWL13/eusSvBzEjrLMe5lbX
+kDwIA1QEhwDq01stZFFPmP1Jao8OEo7QPV25UB2O9iwyxE4gUoq6LPoDyTr
g53ndtX0zwElnHxwIFN7E5UYmboGzE/ZcIYt0DpVb56WM8XAe3SRtpzfxD72
D+GdBgYlTwroii9yuZzFo6RhQ9RSrkyg4w401RGOUEIqHSUXKeT7pDl9fNU8
hVDBg9SW67PphDmqjMRBoE149Wsu2bULTJO/6suaY7b7ROszEiJVg0QcjaMn
F6ao252L96urnVhLUe+Kgbjr4aBQiG109SV/fWTy1t773/2Fk7Y+16BBQWds
aS/P2du12tB6APnAKTzkomuZCPob0iHaJsHiTJiwZ9SHUp8UJ4x0pFUxNDDj
dyMc+nDS7+Dr1eomOgHvnixt8OqSc3ufU84anX3GmqKnLop0HRZy1wQPKGe3
E6aKNWLlDBLryNiEohEUVPh+EXIYx9bP15IycjYRts+AZxw+Ld2kVprN9Y2S
RMS/zpRV18keUYOr3yX2Cz8bCJym05JFiYLvgcBY+KSct3v7SdIzl81Bq449
mKwOlXLHbLB7NSlF/sxnRNd5NT2vhMla1Coc42EDb+7aQQWOgxUE1qBfPJbh
hBiEuqYy2dytzh6l3Q+o9Di9lcqvI6LhpRLMQOPyXXEr/gXlEemZi7k5/YhM
ZqM/vmKe6f97O9D7mbUwe2MwSlQAZ1VzkqGlBLvRPJM8WdISPYgOrvqVbw32
UkeJU+mEykd7v5RgmiWPNNK42mfdRfeToIDVlKjaTKO153vTaNptcDajAbZr
v6sP95uvPbAAqfp1DUpTnzxH9O2+bxuFmsH3QoCZXF297y5vDqyawZ+5iv/3
GCq2D3bnPE8V69HsVOBlhk7YD8X8ipH9N0ntpWgvvyTaJuNRrihlRj12GRqg
/p7pyM0sWONEgcDyaq/BbN0tZk8I/VrikksRNSzuYsuKRyoMKt3j81QxWhma
Ain17+PgxTxwV/5pzXLEMkbSAaBS/Fr/8vXiWIYm6KJy3WkNtaX7DNyGA1gR
iQ4UaTSfvPSosJM2NX0tBpAHh65TScq1zgEgbd3UEMN8lbL+N1MCskimNI1n
M98xkqrMmzyGqotWUNog10PoC718V1o7BcBpvZVOUBIDlg423/4EiM/n3Ax7
zqh1lFq6cO1nu/ZfLrCmjW7ZLoW+CxOWy/wPHa3EZH2i/XqwcaVhXViv2amW
Y76+Kn6/ahVwMn/2eYBd34uKx8m9RiJJ+ElZTdoXSq3NM7WFi9wL5uRVzpoN
NAcwzLmME695AafN/HPb62R4ioNhOwk53DhgRXpDBxoUoegmNEE/iHIcKT2y
0XyG64XwVloxdgK1mtuYjS6DlVNF+GOAvHpja98bcq5jCBozIUM9tpBfDKTy
fzsjNct5CO2dc38U5PD2FFxNfiCBxqJXZeiS4siokHYLBZPBhaOck8xm3RJI
f99eqVGvjqSq3iDNVbzsUVBmcSlZOrF1OTjHeHPlMWdIXsKxung2dGTU0eFn
pVyjz2UT+HOcsRnIEYTa//OASyNA0noc6C4LYFuiYBERK7l5ucPtaL8R6+Pz
nmIJBcIsHT7fZgPaG3PwNBbgdNfxhk1Ov2VjiY1fkgnSwx6oltVbl/Id1nRF
4YEJyiEQL73EbAUcnu4ad5RJ2AM5K8R0PEmiPM750mzxnHhAl1YzkGDiovVo
OxcrsS1XHMg7mHLoLmD/4QR8nwI6fXjZw1rmEiJRQefAvPCcO7/EAEA7lKVU
+gZB5kj/fnROv2G0TH1ZsXSK8/aeQQFIs+GV3EP80aojh/5kP8e65dlRLdQS
YqghZuXgmJy7sR/90VHp0t8SSTljcfbcyiKMiFYZZeUIomB9fNMzuZt6Pv1B
8So/KRkCLM907PJIIsqaKiM7msUkzttrN5k0tYFPX0T04tgqB2T00vyTaNhN
5JzWGUaUUvumY9PXXX9XREbBzAaLrswFWPVhezTvRFwHiLWGKw512Io904HE
o0K93lgFh9AlzW+6Gd8HAR8856Vwi3t2sJP8Y2XK60m6XBS1xAtkARvLktwS
OzUMUFnun6Y6z1yZQsXSjQMQh8BAAfVeeAkLw1uyqfhyPPJbFc7yWkTiNj+H
tjSSM1aKl8FvKCiML6CFQc0f+PsQ1oY+0XnMiwBGnYHf+jvabany9OvxfQaG
sOGdsjilkkZ8sPY6FbTumIhZRRN//WUJx+GGezP47mx7k0QutZS1GR+AGwRQ
lQm82lv3T5mnpb4tYiYZ09vy4gzYVdfK8cyXahJI9OKhBnQUmyhnpwWMozPz
OMqnOwjtn9OfohAVU0L4RbjS0QHawVT9CwXaLoAuo8yJ9cyDfLsWTtJH9IUW
Rp8bLMUz73rlIKKn3V/+KHjz5DuFGrQDr9ezVObL/DVxQLyXSuwHs4FZtIJE
MjCIF7q/7jrtfmmKxsWZrAapPSsR63H71rmSUywMeoQjDzwDdgarOBSxqK2Q
LRDOsaZBaEc4OdcfawUjFvSrqNwGxhiH8iLb2AEzSd/VuTyNgA6fWoK9HPtt
LblFTitAa7BILt/JEstVSDQj5u5yL/iHhRq/LVAWpjWiPumH4aesn4MxUrZu
yAfCVSfLEIlzQ6o7ihV0mBsQpucJ1t1gZ5PpZLKkTaqtOqsdBLq/2NyO4RC3
Gd2gHqG3hIaogU1hCF180R01IPKRBJq464vzyHVToBEwPVYGf+iY7vAQQCC6
v8R+xEb+u29AhhfF6YXdJCMQT/uFm8dOOAlGejiN6B+2ZhtwkGfzbu0rijUG
WaUsW6ce5qQKjNbkgT1TiLFz5WJQTTaFjpU08F/botDy1fF5vr9+zX2b9TKL
mIZz8nTm8cFofG8Co/52O42EEQRANfMnSFzLyr49x2/DmWdrwOD4Fcbrw6Ie
UQS0dDE0vHNNg+yPD6gwe5eD8QBNgPDIlLq7I/+61r2RSssrXu6Wk5f+Y0iZ
i1bpnH2pjNchWQ+vEsm4qrBwwikViJyXTDDOsytmgzcJlZy4Ng3zIMIr5ZWI
kMqAc++AVZYKFZs2EfsnI671KkVd5L5ZsLhLNPOyiGrAZ1kfmjIFjjjyaGKu
p6qWaXH1nkW+RBmaXAFoMhPlx7Ug7Q9tAL4SXa6okxSxUUwFBb8XH6G+Qi5Q
SuUYLy6ICQMaFJYYHPejFFxo7xAAUZUyN03w4B0ICqHsRRi5KjVie91rwHWR
hatgGTwBu6Ml+4acCC1h8FW66mJmi/COcbGmcCaMtECvMwxenH5QOtIv//CS
W6Ritg2Mc3dM/1r8VX2vkJ86Xd2jubiaUEwYPK9AovQ4Py35i4iSKm9i1n0K
J4Sil6f3QwBJrwnj8DO8SDfYRfBuuref0E4b+p1O5IMlAZejpXixj82qC2EY
DIZQyCV2/+9cSezlhzohm3R76Nly0Tb7s+142p97eA36IukC+jG4PxjI3Yp1
NxTa7V4uQAIcSDebLwuXn/NLXh+Vj7KAmUNYBVVaVU/SfpSXxNN4yKsqdkZz
yTdBE+0bD7Jt/fUEJ4esk7v2zKNtVhlU5jdMg40QEWHKUaiTutxqYuMzk6CU
nsIHWrrW9xu0QrT0hsD9bVI8NRc/7PNC9EPlesOIkyYypfQuUShTUEEauSiy
BnEg7xN32jSpyCQGejfx0TuCDHpzkOxDIw/7yAVyFdO8R5Ofg9+BXkyynQSm
/klwL7ig4yAh7UeZ3qvkEwvDCJ20QQsHFeeJHuQo2j+cFPkoMFmI5NPXNK/K
wOtADmT2J3iuPh3qiSXZAPqUtk4O9XjmGCJ8sSnmbf+WwhExnOPA4aodNz81
KhYUCTFB9SxycWH61qvRvyiIftZFdfBNmm+lO1CCvfsgXWTaOkocpPKf0+FJ
cJm97yAjfS4kBhoaMBHEMKk3/vF08W+KqfM41FRzWd4FoVbkFsIlkI8rUluL
pCtGgJLVXnz+KWIb3O1jOhZnWEANNRXN8Gev8GRB22Z2tKS1v+4Slm5swJG7
6XsbLeGBVQOqxWzFmnlmQEKwh9ybbPyVvxbBfWay/g+RCEpj6VPTUw4gz2fc
rI06UB71UuzU1Gyu8Am3z8GyU8deklWxBCP2ExG5gPlHf7IV3IMqleMA4Vf4
YtMBricEmEhrI1C9iWPQ5PuZR98uKcmy9aHeWalzg5wcA56lbsU70cvbHamD
j/RFvR5uQQL/Vp1MeM/fkwnqniwLMIQlljPoaWHkAstOJLcPbZtlLWZo+RFk
yP9Nw8+xhgGCkgIwoi6k3mwv6NmY+Ma3JYPG4ZMwazzVftVZ2E88MxThMjDf
iVjNtLYheDe5Rsei6CQWrf56SoZ8T6lFfoZ5nRlsb0wChKm5art+EK+29Nqc
aPFOea0qEuPPObH/WMdA/6kqn5gCfFaR5GASyWnKHuM8JnpvRHyiH/BrSGyj
8DUdiFXQqGzmme3f4aF8MXdvQfpILFsj0F28YDxLQ94Vi4Sg3p625V53srpH
2tG1NXoLbKTMcgXSpZ/OpdY/KJSjFeW8EsiNWO3hE6jKzMA3PoA1v+maxEkH
dDBE1UVse1ZmX0oQcdQU5r/H0nMY3hhjo78nVxyPz2ivjx54bPwEjJRwishC
9QVT1N8PscljO5cXfT0+u/W21TSefKu7J/od/N3eS5UlP2ai7tzS179+XJUx
+WJ9RmJrObuiGOc4/ddIWJn1JjQB7sXM794JB4Me6QtfkzKdE04sd3WuSie6
afXe8xgOsdNhrZ0qsakQaNpuvtXHm5QPKioc+PH12qzmqdozX1T8YvrMcOmI
/Q7pXD9lswYwsQlxves5T9SiIMZ5pE1oAHnXbSmeUQdPH75CfV8VBL/iTo3x
lm2zDwTZq2/TtcWwGoMgfTYsrzcRQdDjK9vTyfgOPnRi22hM4WAzz9W3QLVk
W3V66+G4CUZE5hvuRolhov5gEIRUF7BgJ2jhWs94vunH4GQ3ltTjv77o/0Co
If7fRz4Bu9HnDxgHodzKnOxASsRkBfJYNu9u4q1vSUlZP8c+jsOtS2so5yAw
6GOevduxHFCISkpvwIiDASRGVrQjzq8XDq8wHug6fWAAn3anruuWjwArPYO4
MIMgtynbUk9wqRFvBcBQKs7Ds5186yO7HU4KGzz3HmKMdtzLVdox6mpQ1HIu
bmgyk2FYMygkpSqWm550BWLDxkv5u0VHTSRDXmmQ9w3OWd34We2MHZTYFUIb
QiGtgZSc16bnWYmWT2GtDiLJ7CHwW83+3UeAT5A58FcVv8YWIGAJi/1Mc56e
0JCnh+Etb966qyXvMG7SJ5L/wbeu6ZTrtmQeZyt5dvVbYK9aqxp1cEOYfeG7
K4bYleSeermDFzpCmHT0qPclItP8d8RjYrvsZkuO0CynO6Gi+HAVr9mWD9o1
q43Efm2sjYEBWINpvmqIf1UsDDjLVEYxxWYFhWD9IyENSy2qBNzlL+FnJQw9
ew4Mhuk3GZ0Y8Aj/GBZjn8tv6D3CjrJIwbSg+JM7Qb0E2ofQT43LpMjjz3T1
r+ZT2Aa6cCRF899njvqPnOu9GiXHR9MATybEi5h9heTyLx5t8h/5MH7k18R/
bqosb+Uqt/cZLIjEOTjsC4tqAIW8LTFVahziYojrl0tmsTbVToYbP+gdKqHj
wls9pl+OEXZw1yH1tuEIhbtMEXLN+6mqIFyITXqeUXXiegiRhXURJ5ZAC1h1
EoB7NrLunOnjRpDyWO2n7M3bg8ubC04/7zKLUubs0u0p7UUXti7PUJL5kTr7
C3MnArMasm+10Y0CsEVSpPGd/Tad4zorMBJZVOmDMUoJH13aWfMSo9En9dl5
4TROWOsHOxPktvO9ZFpVigIUpG3qtQvoUglPO2GlYIrYbQ8fCsy3A1V8dFwn
S2MEf7cWYLxSb4X6TGkBfPBLdXv5C1ry8LliUw9Ba+OZZGXQHKvtRdOC4KAp
pkiGJvNyScxdm4WY5V0xmyMVG5mq+M5eBSh0Kl6BsL3v1tgetipw5BIvn8rz
6TT5u0BZQJNibR3na3NcNixDzCL4ftQpRfI7fik+Gm/lNICfTN7NAYa/gw+g
ISQRanK74M9RX5oJ3Ht5VAMrAkCoBoqCuuMSC/TYN8Pi/vlMkIOryYQ8TnaN
o4nujfw3L+Bpys3SQJy3ppslHeopHLEN6rS7suD7SFKK5tlmarkEoPKjLkLV
7MZWZYTQi50jveOBcbPdCWsocXDSJVt2gEJWrc/sWxqSEKz3oBgG6ylkKVg8
FdwWekkWhPfozKNNksMRTk2rrSX19ZGTJS+QqBNLtBAkMGubpsewrO9rufg3
Yei7w+La1XzYxbjkOVhLjOzjDiQuyzynYg4yMgmNT1xFMcONq1zV7maaKfIi
Y0IQLDKoCrtr26DdDGEQznq/jBtpRB7pebJWzwW+HnybqzLi4QtaKzX9SB46
wKm4JMB4E9f2q8ZrlYYz/AFUkku4yH3yLtXZU4+kC07PEA/GyDTjXMitCxUx
lgrcuKLlkAOgqZmqQjVS4tiHGgeE8O+Wo1S0tLQIuLE1ZnA9hXhRvtcekmpe
cIEMmAcas84LHUPA3zwaE4EiWBu5U85AWdjAjwQBTPs9q0ZZBA66Xcd5PsAx
GviFyEylB+WUY7hK7Uhj13iPltzTqKCW4AgsCorRt3J1mDWIBTpK8aGcslE0
jG/qKppVOD4hXYwhXhoo3+hLP8Uyy6T5ndw/uX/OmW7Mc3MDTlggOkcp7/hi
SRl97E/6QJXJ7QxGp1kUrjbZisPvQyPaCsvIrnVVOMdn6kcw0VlO5gJITsei
MrhCfNk265elzGi4kAILgZcu+AQ/uO+6JHu9C0HJIchRU2hsKhp/ryaaUM/e
Rvs13Z7ydrfn1zmNXrLJ+2iivkQHN7/0KL9h02V8jAVgiXGfOfENBnwiLNHH
0pkPtUDo8DBPpwqQfvWjQE7HdMBQzO6xdECVwPr7kA8N8poghwTYhlc5QcBL
ecjZSlDSHx4gcK7k/gIU38fw2+zN+HlNakg4CugQNogLXgKUrePEbSuPyQxG
jOmD7/AGaarjAIC7dmDv7NMZYPbAfDEuFn8sRV+6lz9HW7ExzIKvXds1dIO3
sqdWGs4HXMn6ue6QNpT27fTmA3HCOjixgyk3NbYMXGPEJGooxuHleL980Dqb
dkF5oI+ZGl0AnRGjJz6l1e2Zy+7MV7n+aG3mzssE/EMnYlGiuVk9a/6rL3Nu
dENG/3TFN0CXCZxrrWzBCpvgaRSNifMbEw6hyjQzyqaJWg+wU7fMkywXO/6k
yceIYxBw5RuCrRMoP7rtNWouM4s0lnoJjbqD59pXIcM3OVu0hav68CyFTvA3
CvoOSyN7VACtDbQD4JbZrqsFlmzXV3MQhuAFDfYDTJ+Iv0fybsxMvU9KZT0i
VDDe141i6KdNcbvcKKKaR7Ojz1fvZViO4lRfX2K6000Gm5xyOTG4NXhykZ97
PuV66feh5DhjccCdmQTJEVjlxTnkh5hBec2ndBDkRtCT81Ug59o4dboFrnek
thxhYz8IqzE0sEAhfLYH3uMOlk2giiNtteCcqbqXwCcrsktYlyFf00AvAPkX
6GAXlZVeDINWHpo0eiHlU0JLqry4C9NQmj6z6GteyLCJ/LXQjZAIG2X3Cqnf
q7OAC0MOgJN+y6AXQO/l9gjhUXB+Onj0LqtYwJJeKRsys6EZ4PNQFq6Rvd3/
8a5ftPRZTa5bV1NKN9ADLJHZm2pzzJI5NE97aaSN3+m7kTvNDqpHpNo+pPV9
W6wPgCFd6A5kqgy5K2HaeewYY/Bwhq2CjNElKeCAqDAVPXRijqDR2Whp4Vmj
9/mjeosiDt92RfmW44rzY2ELl1pr+HsfjKN5sC9Impz5WTbGkOZEdh5+KVMZ
iIPpC8Carj1aEwoX+MoLa1hPKc/9eH9ahtGzS+2GTDYPAOD7X71vPA9pJ80Q
tS2V347LAvs6bpwSpUw0SzSrEnwLA3UUIHEDKDeeqH8fiAnkQm3mqGG60lU0
WkXtBRVAh7KsZGmoAJngn96GShVonmb55iKTb+PkJPbnIhwBjIyAlBWQeLhU
TGBwsMAsDUBZAYmyeFWnCrBWnhYnL3FTX2FmHGWfUv7WmQtIHaqzFvVWr8T1
EbMTB+xEDTaURihLPS7RSpL9teXXrYmVl8CsTwVqqeOxlCDDfFcMCKMq2qho
4F4mkZYtxAmtWN4umL/Sj1X1JBFErAAXdVxNKdgwHNwPdOvlz/cUKjTNyOtw
BEm+3pcvQBR+et7GhNEQTeR/ylwbX/nOJDnfaLoFpxaEBl5c84CEzOR4Cw4X
DqIJxbwG6U/O75zxxvHnsSJro69CfJl+Y0c8L71xCvWbSnji4Ddgk1mS6Djb
AjLL0jJ0Lsq0fHUYRv+/1haTw02CQ8l2jl7JY44c8oKpMe2zqaomeaX+IGGo
yBABv9hJU+JIRobyv19e2dfaLVIyPPf3Z/8PxQOlBUM20ORKkfAOfJfbv7D9
KNORnanibI7L75ka/ZcwFNAjgV0msu0Eua8XoEfOLJp8tLkbF2pm/nlEPo5U
MJx+uX6cIuPuv2Xxf9fa0Px14ZLlAnJrHZ359H7H+kwbOkQ2uNJLVsKJDmps
9Dr6kHhpPifdQl1CN8eVyUChx+g2dzjPzMPqm/QISsnmUyTUgAcX1bRrgxet
iYT+Ta3xYPEcRoiffU58gdWos82vGNi5ndIEkXiFcVf3GSDM7+vOAhnPDF5+
dWWM/Nti6DtCB5RGrQNwAFAM+CgLrsjj8ipKW8mqB2qB+P/gcd66TPD3GosA
Az3iknb+l5lZObNkPnms6dVZ7ImqcZkS67Rib1DkO3yPf66qo2cpJu2nkJF5
x7/JZXiiCkedZszBj3xSHGI+sO8aj+2DuaSYXKsW+6pOtXsZoaGe1VVj0tTU
zJLh+hfdPQlTNwaog5q5AfdxMHhFPAZjG3NAyslJtPExnjg2xdP7VJzf88mg
M4sSlFcSMriQBFcfPEwCt6vm19C9UL/Hb6wv4+s2EIfATGCqWE+fThR/hh9D
rfgaYYexxP/0ByTbYG3SbDNexiWgPPRcDdiH8KCDn+6QWDO7wqfLv2sxuulR
dwr0LoYFx14O9w0yBIuvCAzpWrFYQZyCnmaKoznTteWMhf2MfpyLU6J4rErz
vPMpiT/eXP8J3ssGUh5fAV8w8nuhtcCoL93UxWtkG/hoidcpCfC0ZT4C/bbz
AEY5D3Ij2t68WDlO5SdBanFXaE+Wu3JidqrJwv59TojWlD5etb2ZRgEehseo
S4aXZJ+PS/hcUS6U/ZsccgzzCGx63miD3wJWCI2hm2JATrAnisHxOIEMOmwu
aqh4xy8qdGoTdknkTjdIXWuIcte+IHvFdN6ZNabAlcpVU0fsGkAj9EEcrvjf
ppRPTd0l2CbJWIWHdfEQU1q9u4Pf2Zo/aK3dXXUtRMSUF2On8l+9kFsQKnuH
kXiyzngu5IrKJ3kCDO2AjWeGiiyaBdQj1jg/2wfPfOrp56et10LERvUzk1Bp
fJhVqiWyIGIEN3GcaJihAsk8MJdSXjWor0a/Ec4kjKT4uuQZNisnrJZOwG02
sbQTFF+8J9JgxzO6Ntql1WCYJWROkBzfggH1h8A2skye/8TrUkTbc36n1Rd5
6tp/99ASEgBy4j1FdGVL0mtiCePiLszKP1zy/1D1qRCkobuyT1xeX0cinkuX
SKei6msiI5JUYoi3xF/Mec7UvF+gbe7fgWoe1jZEpneCAeJ14eEFqPWSzKHG
2A6SbVNISh9wyZCtdU8q1k6ooEb/jsQgzuopm7JZbuSzVeh5ScFAG6ZxOx7A
Vk1FWxwl0ruEZXSlr5hTSbC1nOwdrDck0g/wcKbDFKyXosfhOh8ZjujlwWZT
i3bnlEJbm92W0E42tCkrQTHNpydXxIkNQTRxEfOln0dPRugYmyp9MoIP1hAD
3Su2dc4JM9pWVLTV7puOU/T6LLyUho1y5SWHRvxTnV9COu3RY3F6OvyM2MPJ
ApHpWGN4NNEnYIbhQUy1hh0Kqalk7Vo9Dkt8E0XE+eF96rzyW2d4I+QBK/Qs
4+IL7WPnRgYyOnHasEiH2Nnt3u20ttfVUcEf30CCpE1MzhWnuw7MUQUE33+w
AXQ0jnMq9RVCdjqcznV12FmZU4PTxzK4kdlBX47EBRsgLBwX/+NSN5DETo4/
fvsHCfGculqA4CYjTpu6N/JFAoKcbyqTu5CKekvGI5+OrEXnYR/b8CpUYwoD
O+FvaZuNfnaAC9su0HCZbuAVfrcs5/qPo9siAKy+GA+8DTHWKzdFVdXyzeED
SnQHdd4+Og9IoxepR3IWLYoGTBYAp1HdEWySjcEqXGG0lhOXWlKgy2RN5a6V
zvo4jZOj9cBE21cS+ILaENPQyLQGA4z69zlsg5Rxnb/T9WfQt9IaJJYiiVqX
0WBmDakgCNRkKt0vykDIyj6RmHHwjyvCcPYA4nsLasK6dRTcFtwdjHwTShVF
viKsIDvOQLcJqepMP00b3S5e+QyTuUH4hjdpbikjW8YxyU5TyDFzIWTTpU0S
QgqoB1x4XMDhMX9xdKaGngrYLiKosioKxlKLmVsLoqSuwQh/g2XeS6JBafKz
3msFmSJpKs50mnP/eImdgCi7dMcsskUgDk8ST9CEhXhPxnr3U2e9uzZVYXiF
+y570dOovNKlLUAt8inyZpeGMQ3I9HlazXXg/1XTZZ2Ewv3Hl+qdf/4SqzD7
UNBXAPpC/kPqmm/3MptzPinH6f971TnIFMZUjY8rnEiT/yCH0tK8zizK0K4T
xr4NDa0o/hcjBC98Q4qUhFDkbgHKeAPohHExZZLQP/a2aZVLFWdF458y+0o5
unDdv1LxknwLFD91a4KHgDoXyxTAxAtF5umh5Xo7PhiHRNSB6PMagq8/Kp1D
R5746yFwrd4htGXZAPopkxmto/063h/kiR2pvTFh4fQ5IqXGVSdhAMyhHCoW
zdZSD+6RVMOzci5D7RjH47b7q7sMkyxsElugyiV4/l7WXU63SEu/Zza7JbrR
I1SP5clQEak4GZHN2V65m0iGFB/4Jz2dalUZE+EM4xOUPh6GVGSdpCz6K0ct
1Kux02dC4gsmnnQoGiLBUN7yjaP3oJm2HzFegw2XBBRz5/Pan8DJd6Ri/Xhr
rUaFDMSKP5PvLOOqkmCbw8MwCeiRY+5bLczw8Zk0QidIpCy27dorSqhnwioh
l//hCBe2X0NzqCLAPaPA+Zg2RqfBzQF88ICcPsRmpyRon/1Nqx2Vn2HuaGBk
2GfD2Fns97tPbaCz+IJgpgv5L+uXzk1k+JPOfZpvG0EYfzS78Ew/zbNRgo44
1nNar/UWi0BwMsmtoA3SXriyMT1CS51+GnChoLES0wtgZSqXTsv73QJp7eC7
nGDCELlP6JDYPz2f91sxpae3LyUWXkhquzqVEu5MyRlCPMlWkfuQJTVemYuP
Poz0cHST2EINxHJlRs705sjskCEhEQ3jwbi9b+CvpGGz//xSDXccKNbh9xRv
TVcmVgrbAFoB1nHKJnDJ6AamQvnWnkIin1Tzio+Yxgn2SlGmVC0XRjoyiEF7
ODNEFoa+mcWncS/6hcCm5GykUfXJ0nqSHbSMdlae7s7bv8lvtODmhu1G9aK8
W7Qw2iDHEE9y0Mn7T/JKqHF9yN1cqfg0FKUZtjQ02b7TmObDRHQ9ayn9nT1w
PZcITJl4Mq0PflGUIGPqynNHKSC3udNpNpk0G6OFsdluYUN8nzB5pehXF4Gc
J8GzsMW1lUiw+QUhPdKkpacnR7ZqIVMHjWBoSfdlOhmhKq9zvlv22zvikN6X
x9Y/UCkNDPizuuPENn+BFjGEwwL+vc+UXhtWpHoQywstnKZ6ms54DQeUlLM0
ZriojuzgXtoV9YSQU4rYadtLGt3Cf6Qx+7Nqpyo6zoDfXiFV3V6U9cfX6JYg
tHvQ3auegJi09Af722gilDeLUICV7kJVjUmprCL9xvcmzhX7fRugnIEWad4b
0o8FlXgnk7t8vRC9JcATtu4THPX4RWb3/9qfn5X3EiFX8FLXVs7QGl72jCGk
2NRzheoME4PsN9v96cuqTCFjIlX9osFvuTLC0bsUoM4LGGQ+r6krY2U0tSsk
zpTWMAJJWByZuH6roYUodAaO8DPHmIBsqh30t21QCw1hQu1PkvvllRpcmKbH
hp3By6rdmOtM9MWGpgqXQcI3MWrAKX6eJfN181hiP5EGZbAWysHbrRyPUdRn
isUwyIhQ66EpeK3bn3IyzL2qMdAxXlBOWz/KXSsv9jjDRFO6YineJkJCaM7j
+1AAR0lklvDHwQ3MXsvfXulJVDzf+3cWaBYDjYJCb+otvUebqqQQGopKrSGM
X2PpQRHDCuX8B1QXu7ehJCLDZY/uQhhnpev6tx25tZ+XfnsFzFPV20LJQYyN
1jLgcQ/MCgZVJaRLzvw+oAKmTHRDVG/uIAe6kE8X/GojZ52bX6fNpuBQKGgm
4D/gBXiDoIwPJ1GorW0R75VgFRoLrdkzE3JL5UFEdjmiOpspkfzMryztpOOq
zVRcQBIkbx6tBJ3vTOXsN9ejOuWQ1umdSmH9YvNw0znTwm0b497PuNreUeu2
tp+NFyJQjmVwjdtl7Zu+E5p3gCSt+6/qWIN06nNxQ47gERQhKxK19Qv7lFOs
+9N8sPyq4poFWK0MVpndiTcrVjcyClSW7SNSl8ufhfu/FgtZz0z1k4OrojY2
BItvxw9hKsFMMqu5Zgg4gFb2UUFpNFB0M5giHIYJoDP85mbO+7DicHwIB6oJ
D28jgbxh+xVoiE2Wod6/Pfur2BjJJBB/PU77uMPAxylZkffkLeFY/afmDvRU
4tgeTrYfodslycm8kDS4WV2wAIvdwMw1AIKjsUMW0qNHxCXhfheR9n0HcTVY
8SQZypGzw74Aq1KJ02tayTfP2s7YjZwLGRAbybHg+ZRMU3tQHyfDNj8urYek
azuVkFAdAcv5Qsa8gs2CMuKnac+7xaT8IU+vbH8nYZaJOWfzTmo3lHQ2VS/s
guTK8QmI1bGb+JXhpmknSQurjAKu2hLp9iyqZ7m9JoOl+hotsUuFT6yhrjif
Jmxpao+EWfvWn9Qqh0spGwwYEiHaXx2KsmqJzranGXu0rB4b6rZQHEpRQDds
/Qgqkdr+vhv+rxfDaNI2jnM+oGKRCdXlkJKOEHGm7UGzsVtGJ4pIsv9oH7Bc
GmbQsYhqtKzQo/MLf6QbluUOd02iQXM4e1Yu4h4pQwsxhoMtI8aH/NkcRrtp
zylMcmVjP8SFf1c41ktUSeB+xjG0mXoF60GKbhpLz4sVMEqKb/yWFNxor9Q8
9DYg5C6vN7v7P4QR9rxI5IO2z6I27p8tJW1rEl80VCq+sx1DNzjMKbrFSs9b
l/LWZM58q3ptTW8Uskfg9GpOu1uMm3themAjxn1g5wMvHqIE9+yQuocuMVg9
izo+0hLiQTBMYygW59IXVq54UJTMK0cKSbxoIdnjeWSR8ZZhfqUe5pDXgCWg
0P+5LakOPO+6Uxb0Vdh6Oqi+CjHcZXiHGDb7PcIp7S/1eueWgHTW5g4bxpov
+3XdE5PRbQAJiqOrb5MBruDdC9ecVRqqi7MEwHZYbIX2ROi+Fd2Az9Orla+M
/LRxGS4KZqGImbEVzXS8M7GllO3MhVYeBlncUW5cbi6c/Xn22jOIwdgRWtKc
5yZVjhcFUNHPKzA6f0XcYAH4X2yMRyR5y1v2iG2fOSPMa/qvc2SMgWFY32eR
X3kc6BGfiXQFLb/WQLBdMrKMRKZ1P0WLPkyUiFuo5RufWs7xFqenUV1JaKf7
Xqt2/OvB8U00CfVXFKvO3k+JhJbAX0AG4yVWrZFyMNQ0KJQv4RPa/qSJ91D2
0g1LyIKmk83HLbCNjBc7eY/eLuLoAIX55KU61Ob/VbAejAkhoDMQoNATQyFp
xYaEKjVpL4hkTEI67fxD/YOYsKRpC6e85FIXOLyZg8nAJPgumxwgyEmwgDSl
yQAtDFmeoJLdUaTxcwCkvRXQvmn5yNUiIJD/io5/KO3w3YDdZNTuY51NmPCi
2UbRH2CEcuqWzm4wyb7rRy2LRAa1uVJAD7SQhlbU7M0DlN5J69jTpxqKApnk
yif1Kp6L2CwDejSI9EtVCJVXLXiN0zFdsHL/jKG/kRetL/kMA+ZcHlcNCoK4
we2WEJqDkrYIBAzwYMmgLJHDAMCVMwkd9fu6PIl+bZ6pIyid1+XKgUu1eB9j
tR0qPEFBumNLpfmDMiqna4yUELqtwiKII1muzJLT33ZOgjy8hurxeDYSQMXJ
fncExcVWZTPIacWq5siBhGnLFxmofMi5HgMsQGPZxZoNq6K/QxEr7ipKOpZ2
zleqxk1lVABoSEZF+zvF7lAJoAhfoOaMoj6CI1OYb37NUfwLXcZqA7e2RbJN
tXkCqg4AZa5rBfrxNaKfq8ptip5DxmhdgfDZmV/FhH+LaIGyDtrm/Xf9KA2c
X/OTO/YroEPX7BWEC2QguV3lIwQF00tLIMYkn380QvZhXMQzq/Kfl2obYiLb
w4wnZQPajZTA4tDQera9oZ4RzWPg9cfq9ymE3r7T3mkh+sDQe/noRIFKrUMC
gIIH4/+ZgBsuvfi8tJEiskvcXGEBrbw3uWm4+WVqdI56ZDnx3okA3EW1+G5T
4t2rCLS0w1ciiB7Q6Zddesk/oi99t5quiF+g1aqCk/Vo7x9oGfHsP8RWMbSg
A5BLwHjmea3gw0kmhDZ/8gCUt7Ss/YabHxvJWSzE9ORbQLPaBJ7UEJrcixWN
8zeFxxIZ6lJwXDy2/Lf9fejdUvpw6ISpv0pyj0A55xy00lwKD0sVKCWknadx
smcsywT8gD7BBw2hVpUg0h34OFLOKXEAKIQse6+m6eiIVhngigzCWGxe14c/
QMX9ywM+eZnO/LOwAHMCfJvFPEq21f1YpzAE/UzDK82VrWp3yAUQ9cqakqQM
XFHhPISFQtMnznUoIixm9MyF/xySeJ/+/su7lRdYwBpIh/Avvr3AqlSKFX54
43zD8+grXH8wkVB/ncZpAqAdDjaybn8ImojRnaML4TTOxPvK8BywrlvzQYAP
SciMSra7BdvbGLl9N7L+c9VCQboEjJjfFckBPGLG1GuJQhtSksp1AdH+T7c3
/dkPLEHHwGgXFou4xOLuCbXsX+Wt2WflBKYk421gxIcKIk7cIEnyVt0mLq32
bGlPsyi4+7Qu93r84zagab1G9QC6LYqA3l3vVt+mEBaOwonneAss1JqU9wsw
JOuqHIrmCgyHz7e8YF3ivKmAnyoD1Tc65GofQylQtM47UZwCTjPHXUPbg/rB
NRBW6UFRoWlegwCSD5cUlVf3TSksttHLRpRnAEy0LszoayfOZ5W7v44boFgY
2VRO298tHOyIUS2MmEu3VYDwpq9+RuTQQ4FIgC6CAfUWS0Ijzkp9duwfvDsy
lzCfKdjH2LHKo52fsaDeS5EYqI5PSJJe0omIcDpAITRsJlq/yrIdT1XDOMzu
RLXXTq/18dPwla0kV+lPsfuU4LDcWXKmBsm4Xh4ZTxoPJAeaseS3oYd/K3tp
xvRsqInl7UmDGf7rATv2NSWo0YKiFHbi2O6xAlvIT3YiRM+u0d1N4s/OmO8x
cmqKLH4foHPIgMpebER49uuU1COpXhJGuFs8KqYqdwOGKY0Jo8cc/BoOE6Oz
ABZpA8H1qneJvp1mqJFnHb0AOPpOnMsPJB3y540MLm/IXK3bnz+UH83GUVDs
6M8bhakPufDpWteQqdJjLT217l/yaKMwKockXdq2t8ItBi8VazBXRlb771B/
VD7gAgJPkRbwkvGBnAQL0NePiKme+DzUnJ529ehzhJpLhXf4vqTtLK6rzXoh
3CqDAXlugRYSO1W+1r+EPLrXgYL8RbwG34xsKdYIX0cjUriif0PF4foFijsH
dSi9eOur2V8vdAwSy8FI6qAK/+bouKWPauPA4oafu1Qzvkq43hBQ97Y3B3Oq
3tfYlUzqs6nVmpUE0AIq2qRjGmDOnCg2VGEnDuxuWd7OSDw8TPUWvvtwK/GT
DMo/QYo5F7j6RcBxGni3fNDfHtoFmWWKy/C9xiIc3qIFvK1Sx4oegRcFu6zy
BNiOjVhfVcmzF5fuGd8YcoYcjIkCbKD0clGXKjJz6yJflQcubWuPBDUiEalP
dz/q3PmSe+SozL6gjvi5qdMCH5WTdLYo3Zie8Jda329nPtsfsbEinDMu/vdj
Q6sYN9+AQo4OnJbAxCi2UVsa3pmfQbh0uzljZSu94o4JTduls1+hjRr2pMvb
cjOtkW/hXRFiiGkin8x6JQesR8004qRgjiXhSNojwR8gPtFOPGHECMkXaaVX
lseDK8Kfwpc2bfHRs8yS1vJ6Q/q7dQ6ozXDXNhFq4zW2uIozVRizlRsceqm6
6r2tLZDNb6hFc4gulLZezsjqRmHxsnmsMlaMgAZQA/n8K7V8rRTMBh31gCit
B45R2Kzxqaozcqxqf7th58O8hbdMjkF4vOcJS2TwMbNevnqscQyZejenUwgd
dXsBJWxa1k21gGzMutp/NezrHM+m0Am1fP5W9vsuwLqZBCM5mY0rU/HSc4k1
brIObHU3wGOc/vaVHOy0J3mLim9+pqVhLmVe1kbi7gyYYLy7hNR22j9IWw3S
ElUsu1nVpJ0HIvbeK1+n+xOkn4DJern956XmUBt4lbf8Ox9Zbmwqbsl9OKFl
VVbvId4QB0iGQt7Sh9SVywF0hsFyJtnJO13N79iE2FKL71TOoHCtWB1/4vYX
WHhr+xl5LlP0+o4W2a15ZFj3II/zZog7aQr9sQbrLSFUmXzH573MjC4/hSWk
N+JCWLyXGxxd4v5S5LQd+iOgQ+MsJ+z/+NcDKMk+M6aOYDihHsXdcY2CevQc
VaZ+MCyHacqhlI3W7P0muMcO5mFXWCkAdrRjYWoEOpatguDkM0xaKEV5ykGI
4ZPamXq9fTo5WblGxLrdvqEcw8B9tAsBB4usd9nRgPL5bI1RtpnW2ISk7/tm
k7gJ+m/tJXBpvEeXU/z/W9bpi8lm1gqjju5MZwtb4dHNSMLOvs2RwTxVEUzS
bdtig1YNLriuYVkANMtVilFyMDF5QkOaNDeR6pgbaic10Vs7gk/Sf9VTOz5M
guGIMlCnOaRxgWvGKTkofQkOXw970qg3VHnA3H/kx5Q9kNfpWZ5hRBsbIyWh
DDZtIMUWulDm3PKDHog720xR7NaeLnI8OgUyhScnJuucrZ7D5Hjpx5j4FEuW
91D+bK+/WgrNNLeLR4XNcG6+D3qMoZF0Zp9M29l5fTUk8sqe7R1ixE5N5pz4
lcKj0IfEBcZ1nWnvNqK37FND4ikep+T6R5h080lB1PnXoULzq/yr279trcst
PynPziGjB0kOOo6cZrdc8nBrQOAoTVr5KyvvaOor2rvtdVBkm/gkVzgK866H
nFHOC1Cm4VUIjvBA+jZ9NFPOn17yfHu89WJEo37NaCM9ZdWj5lleeJLdp6sd
6nOS3Ms0CS3dTRXR3CuGSflaRbBMlHFw/oycguzY+H2q06jY1dKAVRFVyKWx
3giGMfcJV/WTAyd91jfLLAvjdZLmUGIn+WCV0vDn1KhLbjid85C93/7zKVLU
D+U7tfZfghValM8ajCHgHSemzGPRws3X+Yr0jF2EmS8AfkYfo0aU0/Y2Ydcu
xHbgsgWve+h3yYky+uRWRxSaiu9w52lFxbaBLkOtFntoiXlxKIlwaW0VqoBl
b7+2RHfN5xbZoUya2v/b8ffpLGwWNh39CRhbEKj+ooL/QvQr9RN8tgzx95zV
RCo4L9KIwDNqP5W1wEJZnUke6Rkya7CDoP4z7W+j28Ix1yvMHi3XkDGuZUER
QjtUWk2bKmaxuCmr43/Vtvb1Q4VmClBZtvQTFPIBDeiK6DMZ5DNBUbSgSiAA
o+i2Rj2RPItEh1ejuzaz3PHokjs/l+NrKcAU8U2kliJY/q3IJ2TqF9LEkYNr
XpsMLkrZRLtJtW7goIDpGnvxrFnoVxYe4MmAxMsoO9u765VeerfRt3cCggHA
eNJcnTUlrA0EWBpWV1SKZFDkBrLjsMBL+WrjROvDpROnuYpdUQOQIucxBmOo
OBmisqiu3HBpdyUjQCR4p+yPoT7E9ayg+95Zqa2SOUjYycZ2MMWG8VgX8b8d
jh+g17exkawZzpkW3RWfwxbEt+CpWygps/sptdIgUUfST8po4gCzUKyJ5gBf
idmYeeS6jISP6gjG3HHNlp5dVEziA3BOAA+wQzvB1wo3E9Lh11Qe8isZ+eZN
EkxAsYaw0We/Qp1eVGLNcnD1wEfqqd6fTLH9nwd0yZZYRGRfno5D9fpWJ8NB
d6jRr1faJpY2eoYdtVI5Rbm6kiKVbCAclb9aVGZErmpWP437rLD8wTvW+2re
AFFCbXMTNOah71DuvtxVY/PrMIiNCs/OH+0RFsrv28pnhvIGDLg12DxkaL1z
WPnTdsqg3ParCl9hipBf1q2umO9kjHOLW/IxJNXnjtWRqt3BHY/0SrHAl45v
K0t4mKnGBjmpS63LtmbFYPFUdhR/jpaOyqfH7SeH3lMkIgK7sjJxiTHQr4dt
SJZ7tC1de4qJSHBAT6iVn5nLwIDRPzKHOalLxRJUNbLkOVpLXlNR8dUYWL9d
FZEi2PnflFh2z6IC+IfmC3R/TBOYEWcNXL0fVSQmV5B1W/NAw+xl5fkgEB18
HDN4M60Na+BQsJlOC1Q76bybTDgETI9rcnApydnp3+jIpDH+zw2WJEps3eyk
B86fIc9ufOVXNQH9vPdd7FK3BXEZIyQm3QutvQDP/tD+i1FgbBJer1PZhlnf
teBjf60aYuCNTvynsapOKz2k3XyGyMbRV2BS+6De9w98ivK9djbo43RvX5HD
gturIUeAbWXXJ0aq7Q9JbvALZ+breL56+7xeb+wMYWzWdL+HNJH6VJTGftiQ
r5d75k+KXEnsw5uVQWKPmQoGEflh8BhzmZZ3k29GGSt5z6cOMEFFVmQF3LyK
uPSgsX560R0Jsi+yeN3f5VsW8YK0Dd90SEXpY5Og25NAxC5Ypc0xEvWLWIX5
g6+/HifkbEdxC9j1+NFkAK22vqITtBNIZMdPdONHk7YF8oMUMc4Ux0n+bWif
qfg+yshGhGKM8hkxxWIXVsEcC9EdJkBRHq/F+Ws1h9ZwtZhRnxM7a5X9m4hr
trOZaPxcAfrPrTVZGVXtKex7z09Y58NUfqfcdTvyTTJkXBYkqrCLlSLCEb+q
9Or9D5mwcsxDJhVRNUBhLU7TwKGjCELJE24GYOAp6rDNY5poxjcj+WOad3gX
lx3ZfeoKPw3b1sQ8dO6oRaiFM3hWXlYjrg0XvGvMLfwqSyib+yrHRxTnQqPY
Z5JyUJU7RJA082nAbWWP9OvwHKuW/1HJadfzzmC+yqShhfY68OXxdThWduBE
H1tBjts49aR5AsSVz7GJeWT4CqJQCabNiFWLyZo/k9nDd1iBuM9OQa8rE+kO
ZEFb4JpyJpGPkHnfjJL2Bb9+DnZKlZo2zrBwdod360W7XwdcylbGxsYkfTrT
L30Mn4PmT8ta+NbDc566rzIJtDvdfpjbvDTbVuD3yW743fUihLzOaPPUxNjB
SaCOb1YlHNEOIQzVnlfGULLXzMS0MqwfgbEZSUmR8dbl34Hwu/63/JEyMuhN
1ooBvbko2W19qTW0kUJSOqIvMb0N04YUMjzPcs6UwU9aH1W757qzeyqc36q+
pGdj7F45Jq7p8r3OV841aOV/l9WvtKtkwvDlKDLtjYKGaXJFaH7NqmSEV+3a
HFyyfF8YNR0l1pGEbXpTIHcqZtwpWpjFplGX2heX7j3whQw+SPg35lBjGk05
IAyIEfg24JUkdTW32oqcJzO9LRMiT+GSeJrjslLaHeNzTO4uwjpgOV5UB5Wj
ZypnjJgPpPnkysdqFY7eGlA7jpnYFPknd4QmkYZQQK8nZvUWDq7ar4QQJ+dM
QSHsfV5u8KptGolpFfJZtFUhI9T3m9auTpxeqodPpY+WkqlvH8oQSXEroPNX
SoTC/vBTzMt76tWSLseUFDhx/cxID9OJ4xCFpqKv6YelG6Xc6BFGWDo0rrCT
S9D9Z/TkRNUjrkXUXIt7U0t2QxT1Vju9fKTF4XvoAQE0lmQzddTIzAqm7zHp
Ge+v99eFPa1/y4yeomA4OranbdgSO6LIcFDOjxv5YgWHr8KsdM9Hi3Oq/e3Q
H/VregpOTtnouNzfXwvdJp8FhX5M2pKarbN/Ra3vyXhIBoI+JcAfzv8Q0yJ1
OTIzbZ+31DAhTowvrbXmtsk/0dJlfO6JZ1nPUfGNJOTKot1bnkHQolaScLFo
BNuGU21cRLWZmKZJt8FcpSp17GXDeHGit019IX+cKIX4GD3FIkf2ypStuJ3S
N4GvR6tCVDn6eV+vOqKk/urhZ4ldgWYebNr4y64AALf9B05DOfH5gC3hJ/9I
D3NZp+gdrgyy6PH4jgbv5h+B4Jqr7tEZqvdQ2W+bjAUntDKK7tEZHYEMy/YQ
eK7ZuJkIgULfpndS9uOK0hF08WwQY0GbbWISM08jIe2uXsAZHUmUetVjv7R5
BbskTiqgBEt0aHfxTZZf++IJ6UH2iBqLhY3R5tnLY33GE4HAAJawVWaVDlRP
WWtNL+TKXcT0aLIwZwpxdYYBnKJfi+p8HB5o+KUI7sb34eW5QVkDOTfJHkuq
kEl5hQSVj5ficEZrflYpsBs2iCULCwcBVqdlTBO1BjB2hmCAfTVjMM6Yukb0
Yh2f0P6dJxPSlhAZiYYZHkdZcIqCpa7HEhwFgEDLfLmH7IeOWy7PhUe2ywVu
8RHJbeuxLgP9pgEkHIVgkTU9gnta08UhHKS3YQM2YexqaIJA3YvHHeL4GbMk
KWf5OrhvOxcH5VpDgEPK+/dVod1s2dTJc5cfhlfvLEs02wxOVM0YGRD1sL6Z
Ifa1ZDjMx7OoeU0sOeQd/5Pk65Vs6kHJshlaMYrzPFL3++Me+R0Bru7A54TX
4cf+Y4rcCE7r/xmLx1FjVmTcLZXB2iOPiT3shAHeJtTPdDFAUhTzjLkBVSUg
vUWPhep6/FeqfYgAEkHq+2YRMio9Z5wcZBdCXlSHz4hqHQuuOiRok3Sn6/oL
/+9LD7pMlliSwz8lPbUK8u+DYtbL2RnvdJQwC0plKLD6faUpSu2CV8wQg0iL
3NDP/WOxHAXGzHx+uDkq2JcFoGmBIIDgo5gi8Oz7mGTeCHT+XXxH6tabWQWR
3jF5VSUj7Tw+xmqVDZrWssAj5p6+jUIhC+Qfkndb0I0VvXoXpRs14bPCGtcv
9Te0gp6tGA3JGKuEmxfxdcYSZF+rINvgLqESW+QDWvl7ESzjCDD+XHUDP51q
iJya6uAs5o6Hx8oIwMV8MINOAQPX7oSoJ5cPdRrW9nF1G/dqbKkRQqVNrQTH
itmhBgaoSJq3+tHt0WTGgnAse38HzwCKICpRmfZcsHa68MtNiJ00/B7uWEbr
0kosxqGz+H79wRpA8g7i+8Nh38MeZ7F9SMyok8YLxyM3iolfeK/hXWGeB64h
kVsGyo4N6yYO0v19vrBmsr8gUQo5Gff1dDbe1GHHd6Fdzquu6UDFVP67TB1/
uDjYnarA0NgNjqRBdA2l4y5dL5gcQQy6szwtdViy6mALKVFmXGYv2WZQXANz
Q8J8l+6qIgN+rsEWwo8SU0sl81IcRuPH1dtJpI8C3CCJ/0ZohYZ7Ok9TIUzX
xxYSk5ySUegBg7ZKCLTr7qpnz7O8uXJd9BDtK9vhwDgV68kRMRGEpKyESGAB
YwnBa52dM3E5Rb4xOrPHuAWO48YVkB14cXJ6PMOSmRc57a8yWs1w0Ojeylvy
QZJM8FQgkASbaE5tuB184+0HpNQ47Uee9WKgCJ7F4TuhUp9vExuOPn57HGxC
ky4Km+hPnla59K7Xt+CboCbnn8h8//nFxWYWO2WoHdRhRDG8Y0qXOwXm2h1o
fm285shIn2D/Ial5+VJTM6T2tgAncp+4ejkf5SIc5orWOJkiHs2dDA0PjSWv
V/NX9jI3M2IsZLFr55TSwJtwgVKDU5Zm1pcV8x0xIubUd14Ke7Sq2k6jdlQ+
GteLUHp9R7AQy9bUJsanO8cjcWV08jY2/pXTEMBMlASXDMJtrKa2kXOcAbV5
4JWPpgiHsMUzfh44Oj5zgz75/14n7XuZwItakc7aZXEVok1Pcf6WTA/oaR3a
IaZ+tqAxAafGAnMn1QC+ucU0tSHn5NjcK59f+p0EWPtAB/o2Bj5FKE+4+55U
qTRQLTIQKIFkS6UAGI8CrsVFf5J/lv/jynS25+Imi6WotqcqFjPslOnOH7+L
pxaXg+GhHWEtRWU9Lnjov+ZrLEV6ZSARFiLKK8Cl/ckr3EhjJT+J6IToEmkn
+HKXT2LzMAQ2FP7bEhe9yzwN7Er9265DSxgNOImU+6VjR9EkTpXso+/KTJO5
gl29u6nrv7HhhYB96Ve4WLgCVhBL7XlcxW5JXo/zo2fIU8IQWZiXJbmktWwI
O4ok71/2aBC9L4Kdvy9vusDhm3MlhVqX/jLl2yTEG0IEsl5dvekh6+FpNp+Q
huoyGVGowCgwdopX37CcUCZf8sqrYwrr3fkRYHKp+jZrKkS7aL+6puQAVbp1
mKPW4UHsZObSzzG28RG8OM/P44e6Wye9OCBQ5ZfQVGhiA7V4xoF5r220R1fk
o2mqtsDjn5OpQU6qbfmh6D7pPo6k8wDcCH5JIFcL26LRuHo6FTgmWbJ2K6bk
DlAakItfjrLAu7B6znYDHDUx9O9xODhIExtjlsKULuVtWwgMy0VAYeZzes0X
+ryWw6a2JUH8WzTnKvbWzDr5+PRxG9Lwfn5MCcNDbfbqfkjn8NQrBRzaMNcX
kYfoSoUxY1AdErKp/TYRQCVW8n0OU8cZbQKVBST1h5BGd9cVuTlQ/Ffozbbl
B2Xs77WSGJ/5rsfRcvKFWMcXhIJK7m2CP3Bue0O/X/iDxy/+dFm0mLi6UW97
LWTbycXz2GcVpAJ+iJUGqjM+nRxbEiAf7ABfLEbd8rCMbAvXuCo7FdEFTcx4
LAPBD7FHBlYsGol6DRnZX6JL9KKfg71gUHMZJ5/7QCvzbt4lLbxM7jyxs2mU
S8tOD1Zw5jPpx4SSpAQ7tbcZOUqKyml4kaw1UNepL2rvl9EJ1lN7fg6ruAMz
u6GdOouZE9Zh0ZxPkK+0RjSDPxmHvRrYULJIIG8EHDPCcc/IKzNFgjjPM3vk
VPQdYS1Zt3ydTV7OTTSO4hqBIeiKBqL8lHFqPkpvVwnNFgZEe+d8UEeEyp9t
NxxoGGlCl/YzDUSekYtlbucrUCcFz2kzeNsHvakEJG+I8Hwgic566CqEZ4k+
XGlE1Iny+GcfCsIQElIisMt/LTm11PQwKVpYc0krQLqRHNslNi8M+thDBHM8
AxLABlO+pAJpMlqUSe6ii+1ckm1EAcX+GvLG5CfDqh7VEsd7SdgB7gEJEw0h
qtFkfyzFHa8nvkmAdjVHULi6QG63y5n8sFm53CctFXgQvejTZ1b5+shVcmep
30wmazQKflYp6rlGrpTPQmnEoeGBXjlCvB8zVMiw41O0vubtLSPIpD1tiTHV
s6bSEDMmOfMYJD/1yGsNI+xGs/pW3fKz3rU4RUqI+3iNfHuW8/S7K+FY3B55
0qXt8QS8jps/Ka63z0ydO638etwsC3jBBnvmpjDjGnDXh1X7Dq3nSTUIVMwm
D7F9v0Cvmkl4fXY6Xps0XY+N9WOi+V1xXZ7LrzMn6ytUrGfHpyK3wBskAF6I
GPEC4znbiWnC1ABbDTHRtcnbx8OZ1oLfGJbFGISbQ31ouqhULJaVCK2CA1vu
aafGCG9QtEDEs6LSOONuxwCzS8WIio3aPJzHpIABxes3GPGrc1jZ7ET6Vw5k
SUpwnF1gjkvCiFFg5nU+D7WqKQqWSAgvd45097q83xGWLa+iWb1PcbbCAHf3
/2hW+Fi3PSYD63h9E9fqPdwME/CcWRyxCZws9lrlnmufp04M0Ff2kpMzWaYP
GfwDlri6I8mxb+Sv4X5Q5EOAL2Yxd5oCBrReQmOLae6BPIGVjI1rafOEuIbR
ugZBLy+7jsRFaB2EjLKd0gDlftTeinjelxr/aUObFBG7j51ytG5BH4nTu+mt
VKM1LUXtxrxjCEpFGCeNRNh2BB33jgL9wMxuux8TNoH6X77kQYA+q+/ORiVP
CtzoQzH3qg7cernCdc8lAYz5m/p+qHl76EWsimmsFedaW5Q2i6Kjna/aExM7
SvuaeFqo/+/k1NUjka/1dEg5opw75NAPBiNXfaedsJQz6JkyHVYyZQMpgLTi
370DeMsqDU5ZTYl8lsWg/tJRyetZD5FkBohPtqXt/5QqHnsMdCShLCDKpiiu
kloFbhDsqCrrBfLvrW1A1HC6AWTo30gx2joiqi8m2MTnyMHzjlteIu1ImUTk
woZxuruNJB2G0XMADDNjERyEWS8FuMHfdTEf8hxWZwG23eikAuWnWvPgH4xt
qA7MAziGCqzcr5ichX5uFzOi8FhWPbP5X2TvsifJK6kNUgA0llRmYhmAiCoD
p9U7/s0Jz/jWDWeKwKGOUBabSomBnmc+5DtZN85C9uDCWQxv+AvVJiJ+y9j4
Hf7jXa7/J3a0rKo2N+umqPIOgIgIHJz16c47d0E+Vq10xf8zuF32RsgjzOKT
+kywBgeZqFbPLmf4djS6ILmUPQ/PzpV1yCErEMrBozoC8FCjHFGU9KmbAnzz
eu8el91JCGUHFIa4WEzZrKukFUG/zx5LMq6xPjK+sQa/3S9g9wLa9L5om5Mi
ktzTdGCbIp45m+dR8vWA/o5qWTUzckEYNWnbWmoR+JQQLAdpyXwpSHqeq+s0
es3noqovHVqDmCX8cGajRnQ/vcHIaZkKjI3m1zFqmXY1nRmZbzlxMqqz8P43
HBqTpRMRKv+zRg7L+BY8TQIxjEva+ZfOivZpy1RVtlKR0VYiik7tzbWk1l4k
7DQ+2Dz72OsVf5N1yL7KW0Q2e7FRmyxqQRrIo7UFLxCx5wK95POpDdLq51de
6kpaguiPZjk//6HZW/z4Y2w+alf0+AVJw0peMngmiK2wOaRf16kY8hu/7Gqo
nVKWj2UJ2UWlckIwJsvrU6ieSbnXq+SidtBEnaDsRFDxy4dzysL/y7uKvvQP
qVGIwg6y0kXD5dx/43uZxzeGPeLn3xLP4q95Q//ZDbCCaF1xf3xB6D37jbs6
zKOuCdLJz+X4IIP5dz1+iFYzPtYRwreLMhT2zsoClF5dLh34jtPwPlTt9hHs
DPOY5UMG8nmoRW432JgG1JumFDv3otIV/b1v0m0XMJzchGODrVBToiNNFqiW
n4C3apR170bd8CF8LD+i+wekBx9N/7ZueFpsU5UnvhMhzk86U0D3PaGxv6i7
jJmY0BrsRrSe5iRowlfFKzndBcVN6C3CaSELD8slWk2BFD7GAiqh0rdJ7A0o
qMTiZMOJkYwRAqEUftO3ww1OiAQ59ohV24Wuf3xUwxGQJAWvgJuUGw+4D1hW
CPT0rQhiqSjqGRFZMmenzlVRRfLwHS3w5kNRobpfhzk6QMiDyfH6lCrEYiu2
DqD1HKSo0C9hwS64ejILbaeuGFmGw/rytA7xPFbWuE9dyEYJJovN//d6CZhi
M7pP2C4v1ToM40DBGJqsx0Uwu1V7NJ3wQuzxjcewtja721ti7k6I67FpY+AQ
lbjpY+s7YZdKrTBbrDmyarb8nqcL0rgaRjusIWltasWW5UxSwbxrKHhIxkCW
X0fu3dkq5vee4AD14VBihek1hHsOH3IIWqcijOx4Nt+nbaFC9/snxgUu1oIL
OmHqZ1WNx7wOobolGM2U2k90T0i+CxkWadM4U3EfJl/R6NUWQDaGjtiPH2Vv
uKlyO7KYzaymMlGV1eFmYuFQCLjACBFxKyjY4yKUClJ4pHssVATmXaVueh1R
jrZ04IdFqVW452CJDzHHxB9SreFaZSfw4mRdQyGNU9uomMpxH9ASqtl5BLXS
xz6pD0b5agVcsaQOt2qGdG9TB3ksl40kNwOcuuFQc3a3YXPMTjKwss0PFrLH
N7+KoSOfrqQexrI6aAcG9KwaSDH5Il9vAkI4nZwJsgJUnPlc6PXL538+P6pQ
dDNNPsjdE9CMTbCgcUw+BLMJZbn3qwJFEIR01MuJvq9/GIQ+iot03kH9ktUn
WtG+rqrCpoWOCW4abn57lDiGc/35ckLGlgGDWS/nsmVAc9hHG6ThalGF/1br
VVey96/cw2c4KP+BnL60YPp2W8AdQ1WKlNM1tfV2tKredooWtVSlIfIf2HBb
Td5gt7MrmeM5QNFP2nveh0tXXupCCpqq+P0vzqXC+up0W3JJU6hOz2Cu938y
O/AecQr1hPDOVKwJIi+Ij3PefR/e538sn8XUEbqBLczBMLqgov7q0bnXPwJS
KTAeLZnZGnnabhbc4+qXKZ44bB4rxa5aQdz/RepZlKNkUvDm3NSNSJNq0vZz
OMeDPHcmOuWKWLO9wIiA1KHGaTqUhEvwgmK2meVk4u5c8O3lEGeHk0PHySS9
BJuQYnYrRwwgI9VLS3zvZaWqOjgon+WPkrxF7VF2WOjbkfuciZ4Fxd5ndesy
ToBHXzXzKwdNRZqO558HkSmj4UTjUhdeLfnPtUUDNapCf9Np/Kzp5v+heBjy
PcFYHsPI97H1VHiTyC1knZUiXcMeblzlZClA2/4uZ9jC1oBZwVqbPs8sC1zy
UDKFrCSKKv/I619UGq02vUvse/S77YOV9IaexF6phMqKdQGUVGdEMiG3idpS
uOjgv7nWo42PBSPp02dfmKWhM8ykkEpZwWr79U1dYALYOtrdyXcimHZQQAFr
K3jrpqIYslcOleClN7+6oO75XxUf6IGSG1uzi5nK/zr/bV9/l2pO0gtpldWc
/C1VVCFqwlAJGVmQKZCYKZcdO7U1OdTV7A1nuQ6NmsjhXxcveBHwASSwCLJY
KdG03ngpIsV6fEoxiRCw5Pka/3nsZtc4buIZtp+Ob0cp0TlrlQHXYU4NQwnc
TD9PDVJS4yVVp6rYowWf0CxQb/a5XhACicM7EnBbUyld0DOARnTnwArwObCF
BvYJOuDhNl8Y1Q8ktPUtw5xNmxhi2RbYwshQ4qc7Xb8Ib2LaloEowiUCgJGb
lVdJK2QFucunIxwJvwGZYSXDDtp6NeyXUqQeTpvzAPoyRpa2xXutpaghNFrT
X6rhb26Raz62nc7vnA05z1UTJ85MvY5al9M+z8r/pyivqJ4ImWVMAW71n3dj
iFfyMmWbZ2F3NFe++ofm/sPIBPIAE7Cbe3Z7MvWMcU4WZAxx9EwR0NvwBDT9
Vh8T8dvV5wwE0YXwEWm6MwMnwh1KAuJEPzW9Rlx6PrGYsn63bNPLEtrNZbNS
gFNDfseUzh5yMwtU3MMRinZoJ4wPQOzr074Xw4vTCEg6Iu0j/ET7TUec872Z
UmW32pgM+SKoFj2rsbFTPEKPff3rZLnfEk91N4M+5OEY3PMHi0WbrVsuT1bD
RsXST8Lf+KPriTXJMIPNEm/lz/U+JKMAmk7IvGV3nVvit/N/TjGexKqQh8xB
dq6rX15/3D51ccJEAQ5MT/uVq3ofJCE2m6wXkLTG1AidMxEtgrZztjISYhNT
G3KcOBAy2YYqAVGSCcmxrNfpclumrD8veAM/Na8Ropm4z75bJYvGf1fqf5Eq
PPX3jk+yLkdB1QMMw+oaZzZiJ2UDOh9y1aWzl0qaOBEKSdWWfuZK8hoRFmOg
TDwoN2VCu94tmC/O/kue0mxxOczydbolG/yrSSKkrRpw7KHJQxK9lzGPXxXp
lewx//8LewznBRib1dZ+xWgL7cwghT1ZFrse+57wembpigw9+wM8xx/qVzgB
YC58ok1mKfXmrVrljBeOWDrq9ddGo2CBJCY/cte0PpT68CsWv2Htl9QVA7+s
UdUainzYsc70pZtZvsEl3gscDz12w1JMGfWIK7llMY2AfP5yU+q4SVSyyIKX
iy+vBTRTaHUEHxIR5WKqryNF3T+Cx/C85hIEfDkpMQsD5+WZ3tEM8elt+KrU
jHNIMLNSsBdVRyyWoGifVr4cELS1MDBI5UbH0fCa5nNgv4vlfKcesVQaVpzQ
/v7kpge12wGcMCRgiXQcaHI2qZZHXthDquwt+QtP5WQHVMHqrQ1LDIvUk7H/
1Eg7/Soj1zoLOBG0/f2NVg5bpg5JOx3LO18qWnbQJ/EvGHsOxwSGPdADQZ/D
XWQZxBUfG8G6pFgum7W10OL7nHeNsAlbLhWc3Na5mi0lb77SlVw4w8klp8it
OlebeAPTgCfBVpvtz4JhOrV+mJPWp43NpBZhMHkb0IduCIImAwvIlnXvPioq
iJjPUGIZolrnWvwMRSmyrTWesS5jY9Gv6U6tNMr32Twz7LOZYhh/WBS+EMMj
oseawJiBpd9WbrsX7noXUgap4vKCHB364OaasbZSg0tN8CEUS8MF+5jwNRgz
GORLaOwpElSj5s/DQGro5ut1I4MWr9R+6Diec0pCdqpVVREyviZ5khTsYY0T
O9I+xjsGjhd3BtXxaq9fFM9VeRdY86VEIlaKKd5+e2bGxJ3vU01mvmV6/9YW
vsYM7pRUW027ZJpJ5Yper3X5fftrzDcR+ls+sBkyIQPcjlIt+JX9YIGJ4C5t
SGzLVjz1SyxSem4GjREHOMkldZ69U4oqsQxgBeA77ZYK73FvkbPh8UNSnGk4
J9IXoOzT2zaowh+yrI7r7Jq9Jl7mWRyYBEvxXKbzR4Cw3RwV+Y7fu7yuzVP5
4+X5A0IJ9UqwCi4onI9yYANWspQvTQLN/Zfug+PP0cYbMMr5ACGxoL4bg+Vj
HtC1acEUevKKCny3dbbVuK1DQlQ32Fy2Br+ycN+L6IgM1BTLbQ80n3+ygpla
sVcqgedwGyINmQauvtLjI4fvSrrc49tprz3iRFETBOaXa751ZgvLIPSorInW
eCt/KnQ+yQbtp3+2WpfRTE35fy8wdc7fqMWqmtzTDimATGhkppU9jNWmtZOb
LGVAqGHbdWWB3xa7Di/lpG0ZOYDv9aO5OuTJcKYqItH+laykpgsIdj4hWyqZ
tIem/0hHEzkEfs+4OGTswMXCXk0oWM2XptpJOuYZ2CMj7sP6IM1lLhknJAU6
Tdh+Hqg9M+1v9WZfwdQXTZDzFYWZxk2T6jCAvv/HG5JISj3JIR8W0ALdvn49
TRUK8AX0/yy9Uu5wsI+xdEnOxYaZr+WD5R/tqxgeYtQNQgc+BH7dnvNnKIS2
ndFBT2DfMrEYzOg8tzlZyfae8t0JE9U6m5nG7/GHrTuZ9ZHQ95ngu2xLj3at
l8pIKR51e4xkwQpYhmtK/YDUTf0IoCqePiMf/yShqjYnFS0n1sUYU7P4yNKL
WfSkZN4m9t2JjqEhpYgw/ehl5IuOj6fc9z7Rp6GwQixTAWm3Q3yt+m7ueMrf
0h8VhcqhjZiM9mqk3M5lHkgipLWcyx35GHsPq7cLulSg9vp4Ci2/6bkwmaEc
RCL3ESiZPhi63/7QkOagBfbqP8Ql3AVKDOCrXf13fLUUEWd7+NbFkg3tWDVG
BbCAdS1LXz6qMG7L+Qr742eGtDvDTViErMCWZ8ZTeGYS7urJb2NWsk1FGQ0O
1yzCLdBVUsIoJsX6cjJkTC+YTaeLfZCY7kL2Wkf1/YHjFPmgw0hF6WQXteuP
i1O/eYLq+e8LLS2Ng5jh7UmhHA2HId0LyEbEm9SEfNWPzrXGDT2r+LHbqXuc
cr0lPDczQKRHc8jXD+Z5MY4XGwxc6vzXxS6sbLrwWqisV0gXyKHArKEhM+MG
R4o9zcl3vhxU56gcYpLbOyonltuu8A3hH0FuJxs3BN4UfjNfr+dXjPbPcAXR
wBlLf8XDrk9H6jmuRCX3cDSyvgOR5QaQrqdxORqBUkvNTMpPNJ1K6KYIgKZl
5CBLcArLkZxPvvZrDEXmf+b+4vr+3MEQCnvQZYYVAXJ68cSbCR3MNZ6piN+1
Zq5uvfOaaJwpjunKApo0GXZ1hOubX+Nd43e+XTBA4T/dQE+N8odqngCj59G7
J3VVUxyWbH9NduoENuXmfBIdFPsQq8pzS60auYYt8fTSDR4y3b01ah/P7cWV
Rrr84GVoAB35LZf84HhknAagyRsJs4PTvyrNlrk2YG3xkZGBXHDUWhAt+QVQ
LHcS20evXy4XH+kQK08sW8GOMZwOBGzotzvYkxPpRQWDZL/uMVYzD2DgECqk
ng2rvNlG9BjAHAq0qrf/alDhiHKuWLeeBZpTA+1cfJPEeeqI9pyVmdhscZCg
Uwr6hM93pO3n70kel44kAkzW/tly53SuWtYaeEFF2w+DnC5NrHmr5EvsiLhJ
sml5o4+eibZl8EKtmlhPaIjNkd7MJHzh1EtfFpCwvntlwWX2JIJQPSXPYo1k
FFKcLJlMqE0oDpr9gZVKUD5CbmhAvN+6vFEtxtxRLWjVWlNiONN0oeVG2c8S
DQuz6jFvbxkIDGATLgC/vB/j1vXeNT30fvVD9ZZaHEnC3LlZsuXmrVRZsRa2
0syubzKkz17tdaHzjGTWNGy5avA6ZupNveVyn5a8aAsL+UC4clnFfKYmhF3h
GrhSP5YZ5KaiHVYmTl6RPCWxajFtIFJ8Nd68dtAYufhORZ5YVYy0U1NMNqUO
Am2zUV8iBRMjV/0bAR/U5xPOoS6FBDmlRO2fMMV9EAp9q2IKsc9x40xUW1TI
kSOyFEURuOXI+Lo3ZLcofrrUm+0kxEQM876xIobK/gNEGp4+l0ZDE2ObNURT
qVzbunJa+5dSwohJoqL1TLtDpp4XUTfvYeSMjFwMpSb4PyjfU/SwjaJoqxaJ
GibjLYnzBpgB2tV9Jt07sRGsNgiUYDhAKSChTwQU8XwFPhjLZHjY8NNXP+uY
/mtwsyybMSo9fUCvdLc6/QvBCS2Lc2sSewy8VOA9YEm7z/Y3d0YbrLZLyOEb
q04ZXkhMDLIkJOlSY4DPw+8572gW0t6kWCsGyWC8+a2rzuFFphT1PRHO3zp+
HmVswtNpG1yOgH6x/EjDq/lS++SzKW4i0IP0rTn9WSmXtogsicTrHYlq2p2A
/XvOWQg+9XYIKw0q+1yGbH+9ExHdAIw8YnivEQJN2JVMWIGl4J+vaswy/kOG
3IE/XZbATomT3qXMbwDTmTY0KUJ5Q0DTt9KvfqZ6i/vGgwmTqYz6xHmYOWgD
qss8RwsZg18xHZjFtjUOnJ55JG1sClDnkEmDjsM2m2YJcIY8mrw1a9/b91F/
MTzS2M2TLBgUfHOoTFLRShSd25SZCtk06IBG6YKbHohkjBzkIljoqDBR7N0y
4NqN1/Dor7l9b+6ZMNfC858eGAH/xJbmgFMEmHwuHC/12l7GOWTb/LH/MiUU
+eepzxX1yXyoxLUclEEA8QdAg+GmKnlip1eX61og0CGoZl/j3PpPz5KpDqCv
lBBG+6VwMjm+I4YXAtlZ++l6zchBzjJlNzFfbzVHbWy8TIm9T2OoeathgcLk
z9o8jtCjXZyQ6Ho4N4BNkRsXBHknFrW1Ff049bsdoYlJ9SN8BBKjycUT7kzp
HTAp036zBNcBc63PuSDzMEPHJ/aJjh53Up63KcIIXsdBeBRgg/d0c8rQg3F8
DY6ZSKsmkTWeabYaqi0hpQmaZiFvAvCLXsBKAfsEPYT9Ezbo0Fp1t8rD7TGW
bo8AjGlqN2CeLst97//ltGPy76rCxZ02pqnDRPrSWDJK7Mwjxg7BI6pFt/yP
d8X0o2/FKdz/nmRyepkAOr8zqKAtNHSQlY8ll5EXoA49PInK2hnySRuB/Kt1
9QMYpRR1xCSOGyNvr8uyW1UX+a/BzOrxX8ct6w8EMHGBYupwMUIngwY9wRvl
a2qIniByRkL4a3gLuwdtMjRxnCi/hWvFN+qwAYwOb6pAo7llyDalb9MqX3sq
D0LAbyJj7b34ptoy6VDmoNg943it59lybM65KIndnjGTmaIz7fWSUISenLo3
dhtwF0Cie1ecNLnky1wJnY6hXPRJjvPYRZ+TH60KvpAEGAovKxkkDvDaM8gF
ELFKlCXxLS/fmOjpJNnzFT1+s4AOa4iGnSSk9nY0giy+MvADw0cgVmkGI3FH
7BXf0jUXep11hbe8GYiKxZhRDwj9/jTg4nFaDJcYf7OHI0gzk0ePj95sycyP
V7/04V+gd+xbO00K+NMB9qZSF/NVnD8TbhswRyENomjkaBPjW821wir8LX8g
eldnk9bGmrInK4C+PprWxK18BZU2gdFVXWzRT4WIB8SEepM5hFiCekr+ioLk
KKIM+tJoqsSI/tNPJitaO9yJ8+SafvnqbNWClE5PrGTwzIJSJIruOecCawtm
TGW4ttUHHl5ZCpLPhRHuOYI/4VTY3KD4q2XEJnZJ5wxn640UspmaWNMX5rf2
0au4Wnw3Sxcm5Y9LGpSSJc3k+KzyRG8Gr13rhcRW6iqcEBp3RXB0ENAKkwLe
/TUvtPXIYS+z6jtxaPH6cmsXrjOpjfuHCsvMiZj10hzcluXk7SnxKBHMM+wq
Z6/O/hmysHczuzTvwVqoV4sSth0CBFwijk0mSxBFON/z4ZpWF7H9i7+KRtMG
IITfCge/j1A5B0QNMHP7QyKvfhszbv2g2gBH33cgYw2RBEE/UE+Be4PQ/9+G
/M25z3eW6k/gEHVH/dPqprgI769vi4RHkFvNKL2A9BietAiR+Z9450lslDcF
kfEQMptFR1FO/dfAgmDqHUuEPtkxW+cLSYXLmp7cmgmAcJxLtttK/DWIV57Y
Rs4dQAWChfVfFate2/JtV+ctuPkhpdwg0hubzT27HGhzO09Q3hj0O4rb9hkK
bGtzXuB0M5CRa8DZBjXPjaQfzR1E73VnC8TdByNfqi6HERXtXx3jQl5KMw+T
kK3Q4aoOuBcrtJkMESsNxDZtBvrdj8qwPcxnDATgylu1GzABiqwXycfktoap
B2xNt+sXDpCYW9WwFuB3eQWAbwC2tK1g4SrmgtYgQPu6U2OcQOrIaQV1EZd3
pTmPGVctGd6aiI4VDINiONzcC0nR7ZDjVsKiOQ0eE5FGrD9wF289xrtCLVwE
Y8vbjLH+DNvNyT4akhmuWwF/YNFRd9+3nkZv6H/16bwmd8cvXHgAVSOqEXDY
DlWWhGtHbMUlix9+TPNb2dCbNEtWuZRXWOSeuzkKMiH/sAURgUHnEaUhwlnJ
Xi9VbG4OhbSyWK2KeXqJB5EfpKLKVfzRPgKAvftYzt5TSgFpvXNAVw1s+EzE
vv6XHmgTly7cUxTzkg09etCEHJE9i/EoH8wIR74kfjC+5nB+4Rb41YfUoi/z
8YOEryZTUeem04z71NlUSGNz3ZeR5g8uawOK0fEUdwPrSfR43g3a0J4iy2+h
Cnp/qIwbDQoyBue3yZKCEARrj8mhvVRnxYh5Q0KWRoqcmmQCgvrGuHEjNlVW
vrzSLvu9Gez1gm3k1OVYBxnqBcfk2MMxRTixK5ZAJYv/8k+PehWO3/G1cz3V
AJvFbt/FQf0A+/HMtvvNKZwy4nyso/OmPQnzUp7VuVW67iDka9LBHAyAYbJH
SPl5Hyr0Yt1cMHquvrvP1rT63d1VuA5XsG5Fi4TRjXt8gurJZMzRYomcnPPa
WjCZOYGCocS3iex+0as1hKeAvuePjDb/hoM+vki71nMBWN8/PJW/T/kmQLP6
gA0ChtUZEgOGZnFJPgm1eJAG1TQLOdIEkwz5hUERSaDIO0156Q/yTo4ga52K
KceSCHijWmlZQ2DibiJOTpp4I+ZBvFfKse+RM9OmDCsJ1y+a3wyq6oFeb28R
n2i3qqoXGalrDN2bL4FLC2k15T6u8QQYgL4aF7a4CKOosar7nmfhu2p4NqNA
e5t75ZiDv5X6wCRklXs7bc37IayJ7JE6EaYFSUgHI3ck8bQbL+dyfMLCylkx
llk/aX+rsOUJyC10EHcbFqyzCW6jS4obT4Kov1xj15OKBTJw7RCYO5SCo9Ys
sHI4uGnCBsbAFabzNxWF0waRul52CGECnARRdb3FJ41AGjzWXUPiV24hut8z
KU72OabUhOnUheJm61ilS3YclpISefawwdJP3I+Ig/vMFGRfDKNnH7s8rdnx
PN1h4XNNE4Ib+PMgc890Hcl6zSjxzAByzSIR7+MTB8TE5Mi+QEnBG0m16qxk
MBUpTLaJ9p72llrPnpN+3wHi3mvSVQP+f19ya3r1iBgb9CVpXAZgFFh13vBo
5wZdxJBENYrROPNxLUUb0xiLVOpb/fpuxFcUdzc8Ka5xZAUXhBaIidtMssgV
rUiZMl1w455q7Xqv4OeZ4zQGcbu/GV65QVtVPDH7GFTcYzCFOVkcmmrmbBYX
r9llfuK/AWZoTx6rIS93FEpTkHuOZs9U2tyRVRIO0gWrJIp0JAukLd5pGp8E
7JAiXZbOT77qE13JD/1zlztXc0HCnsGy9Q2XkSw8NYFDC9RNScra4JjAuhE8
zZfTRPbpWCpwQuS8CVoHs7zRvtn7EcViAXSAGgIQajHFAIEpx1SlPOC5S+yM
iRxOWTysnSWUWuMnYATyB9opk2DkClHVd1VaGzkjoGEQkPsIEdbjZdQ6oR2g
Qvefb2NRS1PY0Sbl4T66eJPslJHEApKZnPgCJDvoMLLA6mclsFk06UiXBInF
/y8grlTrZV5VanzMB7jRilzNtwEuRSI7p6hBOObfyzI12s2wodbwGHOZhpTq
cBJPxLdJ7ICxZKAl2ZyETnhAEYYb8MnoNVVB7afYb7wrkeKVqvIH2Fo2/qmT
hX5FdSnFwLj+pyXXVPq5M3WStImxCUxFDq4y1KFXv7xfU1U1uK0bpEhnTZRw
g5yhgwejxFzMmpVijGalmvUbchwMsR+DseNdJb26GVCdpy80JQt3/h8mebd8
nc4I7t2SdfnErr+NGXeLspeiGT2/i0NLzEIs8qrOBVu95tqDayEE2v8+ocuZ
zTLVjWPWv1pyIRwFP/r1eNSajDx23XoJGvzSiQCs13kgsAZ40bKtjV1pRzI+
/BX/Va8zNcvzn2W8d5Ly/mTWGvaDMgp4win6CKOa1S9oBWt5XEs7qwLWHurr
iTUIsNRpYs2t4X990soj9cJXAizdyjlxx9+4XJl8cbFpL1IbDc1Gvt3n/p1M
tclPZcV+jhjnBOitqgP9Wb8F3VaT+QBIem5okUITojIhHZJRo9qcHNZB/Wvb
6dLM6POsuF8SdmKZQMeAeoI7ROdzcjxhrptXvd5LPrLFdsL6Ah5AZfGjBzgm
mDoM4w1P7JyiWcFl77HLLre2/QmURnt2GlDuW3jq0dzo8L1PKrGRxYBkDSUK
rkKXaPCTC8XxXvhowVbEb4Br938MN2Fl8VjLzf3Ie9VxKD7kmbansHR+42/y
tZSC9YCzjczqvnVwsEt1wD/ApRf6Decx7lNGB4cVunn/XI9YCatUFYz2lRZ7
oVM4KlE1Gs6lNR9ZX2bjbi4zybs4JOmHuVLWJd/ZCpkbl+VVQatjkEqTRDuM
RJMMjorJZfuxUiSY7JkSXg4v6A9mEE1MM3zWSnPjM+fmZOohSjAbLdsHF9o4
6FRqZIlmFWYIOybsnWJpyljfCq9OwsAYQWAzq7EbCwOY3Zjc4CliJB5izxXG
bf2diuBgrKYMz+sG4L2ORoRRLAdOgoeloortIxdsrNSTv0DxjfyAcM/cDX3o
LhETwZ6+5gf5wroZwIQ0Cd6drt194TCe2LDQ4rhUZ4+imZMxW7oukJW18val
gMEUmWfyb2mvutQTF6FFpRYW77BM2SJbyAlRGui9kmSCvP0LTvefYdN/A2wZ
jvyy/TK4QNE+PAQv0W0Rg9KYcBBZqbmxacfFZQbiZ9w/YCfI+Fdxe5HNam7O
UVt89jj805qSpkC/dwQMlmgJ0+/WTXTFKL49fxtQ+8JAxUqbiRXkOeJtDLuY
npt1a/Se5b+8Gj34w9CK0TMaI7j1Q4c5r53Qp7dITRnklKkdQ7GsrSalFXO9
Lh3QNf4HDlsBLeGxz7KcOJe66CzL69Xz4P9kJo0Wc/JDxIXrPUp7dr4+IyC0
Xe8HSvIyfmkaxEgwkynbgXEI+3vElv0NH5eOsXi+tWOjXn6u86aNboPYnYML
SQYB6KxPPLYBzB6gAEVfHKJbVvbaPP8OTu61lckHz3ZAjuZKvQYfzVN93Jdf
hVkSz3AAhO8MsQUGCnY/hr76p1OlFJ4poI5c7TYajDffnN/Gvqi2Gx5ZCQjU
K6fbpIhvg/jJqI8Yx+3/ufRyljOth0/vqPvhaPjrftlPY8dgoCsY4zvQqMB4
6xY4x+8E8kDYFP85aBCUlbzSl0PHoXq/Cc5kHfW6Kf8395h2eiJ0lIAzg44L
clrjL7sUG5Onxj+lmqA2LDRDL5AORF9RAnWsbpQjrsGX5jGtkZA72WGdnD6O
6f+JfpFJ4+bEw4H0IccX4uFKMLOZvT3fspxfSe9xbH9+6t91ShrkLZt4rKd+
ROOlJfQHNAtygO3XSKIU67NAFv2yGbkMkWDjAim9RhvsbYXnQh9opnFQqOHh
/TAS4GI17yEFnWMKeqTzhXCdFJN7ID4kNqOqEop8Q2MsvE7BR65Gs/kxbDLp
YbwCFo6sWgJGtCYwvyYlhIBPoNKlFkIpGsKtyXVIICoTAbUxK/9tIpaK8AxT
/I+WOqhgRR5zkSy0b/Noku/QOMd+ScumlA3PBDAA9FWzLixDqvQ7Vtap/rk2
rkyUF3LrGsmYhYpmmOi91AYee9GQRQ5o8PXBWbA57JzwEB1FlvXpXHaUdWDO
4BECrv3yl3w+sZ5hf4G+Mre4/YFiVUYD30vivD9N/38bNVF1Eum9uC7vhGOS
gSEZTEv+xjH7bzQwkN9zWNT1cqp8W0/nQeEuYrSI7jPPwg7Ve9A9mCXj0Kxz
aO+/mtnnwuNXAjhM0eyQ0IELLhZgxgX8fEBu7xhIZom/Rx5tyR0wyFnlcLMe
7KB8q2t5erq58WMCgE3lFU15keGapDjiwg8muxSjdJPRjcYtjDZ7Vp9Uocki
W9JRM70hBccmAuM6fwQN3U7GiS5mnggbhuic8bMgyXQZDNZ0QTpZb45+sRjM
A62grwpQpNfkEjYZseWP07Eg0Ss3+hC5KQx8bPGQezPEpS6laL8dvzPtVeW7
oAnt/sHLQ2mTJvJG4fTqDHOylpCpCqrY40gHfy3Wg6Tp9I5NR7kTJ+zGVRAM
04IG7oMcMCIsRGy04HoLs8pl/W67M9/eN33G+He1GqpZoOmgnHGH4y5YQPXC
2gQE7JvH4/caGQpaE15v6n47eFFGMdaBJ9mjg5ngXIUmMbDbf3pWV6fMX6gp
4+ZZPYQLUbEHCfSHkUBtPzsgvsxqQo0dl3CP76gXjqzQtu+ZU69ipdzCHkvM
M2I9cwTi6wZuLmh3Eqn3tNkOHrNZe0uthlY1sgPHkctoaYVtnyb3BizHAvKM
rsaaLIbaMZ5KnFbFQLfCNf+quh82mbtVXp3th8HTYMcduu6wEjpplvplrF+m
pOEpjhZzVkg1Zo7b+rKH4g8cnEQ8hlRr4nol8yqLbLMRFtG0w3pBu+u+31td
xGpIbPqScJ2cYbicpT7B8xKHN9Ts4oY5fjGQs/DPD9oxffQ+U7Y+88D0AfzS
BCmoHm9rcHdJzSB/RYJ/w9E/QCGKK7ZheRI+CB/u9EsGvdKlZOE9pyOnXgS4
ajJ2KX630YiWjB/uT4gD1OmnZ77aFRew1jMb5sN++W80GKB0Tdf4mjhyBmZk
+k5+yQTIaqlmWcQuxwkH7WYy6ccxQppbmMqi4WgDSz60NwS0nh5yn54rehDU
GAH82nPuXQcLqxyQ62IHhFvG9Q2bEMSJseWxc8zW6hIcQIrsY1L2p4wrjtjV
yQpmyj58kvo10CbphKD7KRTXu84qPTkKKzz1MSbnh0thMtt6/ZigPZy7Yt9o
YKCQspm8vjgDVy+tiZYZ7Geo/RW9Fbaozj7vwh3zZ1n5cvCt+MdKwsTaVyi6
G4iSfFuR4MwmWISNORtr8buDteClPgpYWj7+AbCF7iUvAEHO98jOBkjITjCA
R8BUfdoEcecpJmjBMczYs4y9uBv8oVIzRvfIfuY91KsITP9xj+R4Iwt5fzSz
8lSCWgjjnMU41LIkIBu5pBtN2B7+56JilrvBxwJ2a0Vxez2mrniByswsWJoo
YUwvrZUCKG/2wymWGILc3p1beZi/bTosezH8mSJI6gdqoilMPl8bIcCVrKxp
MIenYSeFyTSQ2locoe7Gjx78M+VxoE/oGAWd9m5HuTF2g9xfdHoTsZZ6H/kU
Nbod15PN8xIfOidoUKQrOyNLHlRZfQTTtykjh/alEnixlC5Tmehit2iUvFJc
uGwkVYxmPnL4EL2aCln4RNA2R2ZpFUtsiwPNo25Tqf+DKvWUEbYgK1vXVfas
YiL3J3VhIb1S8hW73tegjL3H85LLSJLnLevIMbUEX/CVI2Ekhq46FnARoDKc
m/21tKRKn3SeO9HA/pJgSmQjxSfLa37GFfbnq7IJ3jLyOg+YWQ3ex3lql0j+
Dhx/4hZ6KbGPfbSA0Aev24bCe+qcpa7kybmFASYoi2csdpdIdGfxpa2tJ7WW
4Dm0MMgI+Atkl1KwSqdrVsX5/sSWiE+PrL8LvqzGyJ7+ANrWRl5+rIuTcBDd
2AS6meNTnTK/5IQjj+JyiDL8KQYtbKFyO140kR1X2VEe8iHoVe92dCCzelzb
zO3smFmzpXURZIg2CymIRb0P8aP0A22jRnWDgeTU6dD4rvbmn3p0lRxVR7AO
YSYt/Gbg2CtkECxGkuh6X9XGOwoj7eXbxbaIJ5dtBGzgEWiEd7CzoWGkD8EX
tj6cdylTU4txKsoVccTP8K51W1PYbU9aBpr5GaSfbyIFnH5S0GM42P/7WVj/
pgcTxeRR39lp0knbR1OLcCk6lNWG1AyybADC3NKPvA5cB0CMWJda3kCfkggh
cwMqOx25/PIHyRy1T4WS16hlg2mxCmGn8+6LQja9g4ur97L/BS9J/tSPc90f
L6va2Ix8O7sZAq92h5z+d9uOTiFMI4q2LgnM5d6Z+/duYD5mUx8+7VU8ci9J
MkWKvw9wEV1Bo6rNqr1H1/aYHiVdy59WJrx9pttKYITQ69bVpkpLNT8s6nRj
jPzqAeuGzbjtA/UVNrpr9oH9oR5Ra4G4RFNF30Vj4fqngrPlcJIQuIhBLxXE
d5JYOZxy9DhcYGwsSO0bQjJR49xdmE/Tcd0L5KerbCbe4p3yk+0Fw3RiVZ3I
dOIZDpQ7dPtglX4q5PM/C9RQNB7vgGCumahO7qPTichfZlTcQH/ZdMnkpXYM
3EfHYy+Y094F5/fE3TZpVc4v9mXsF0XXnAqdqZK6RQk0JWzxFwV7ZklqCKIU
qLZId5OJq5uT1ZwiP7iFze+KzNiQXuWGAuY8+g9Wb5PTyUrAT4yNoD6xHFI5
vni6Ya5IZXWHVF+TzRkxfsKb+k+ghNlCCTEDOffH8Ee1s/cZ/I3g+FHIydnG
XiKbAVVEHaB8fivwRq6jT5wtViXQibspNJ/euQwv04ZnXA+AnCViiYgeNEhs
X0MYNUIg8L61QA85YUgwrRb48jDqfNU10RaNgBo2R3HnxsaupkicPToS0R2v
0pofwJ/jNo52j/5OFyvmGE5YnwRhsglBPi6aM7EY5D7ufpjhTnswVh7QedyY
K6X08kl/6t4N/7BxB8rUZUSbcugOdtdBaaEFB9OAB+rO3+i54qHHpRDCq2xQ
CLu9tZo/avAydyIJ4/GU8VfR9NmsVcBkZcnLLrHJ/sAl7a987CDHgH7Gjawe
I9YaqZZsyqKzdnmbH/26AN0b5Rkf74CbWP7riyG0LDx2ryPOwCxrpYJxcjDt
5QLoGzRmNfxzVQITWuRRkw0R84nzv8CDS4ZG1vHC55H5FPsGifQn+kJqAbzh
LFUyztEImUAC+3/mt0D1JS0InXctPlV3XwT8ftVCBSEPLm93zmJWEbSm+ZQ7
+oVoPypG+ldibFVzWFnTkO+QCEYnJ8FbAjDKajLYAMRv0zFSCRBHxva0YUkR
LhAASy16nFN/Md6L2pn0QWX+9oJe+7PBy8dtRX5Hq8afrNYpAqqUxVFKrppm
3RswzDj6G4hGiX0xhkhQfokr05JfKOVLhhc+4J21uhSLFw2BRzaQEulizu+X
ILXap7lCNGlqzS8UzVX0+9PGmM+uSuMGtQFio1NFHsfDMtXAqfS8iVrszL+s
dhfx8gIXD6CJd0uTScY/oSS85POwYRWawpfVqRs1/m8honlLD3dIh1XRu6Qz
GJeWI7bqHlJGSVyEjyWwhd7AEGcDl3qINOGCNY2YPH2kD5nnvaWR6AkQSESu
7ZdW+5rqm1VQf0cQ60bLWIAup+9QiNIR/4Ov8vTy/rb1OYXbPOwo9ODujXhg
/as5pbcjlP4oCc6LukMBgvUTrPdwTv4Eqz2w+Ssr7K4UitLVy0g+CRWtF9R5
MMarlKWfnG+/OW0Pe2eccOq2/o24EaF3b9M+yIb5XC87rYb+G1lHKXx160R7
fCfF5yE6C2Zc+ppq+7YrUNueUAxTfiflHp8Qd6S/PBXICnfsGpspRgf+VgF3
+kAvdufDESHoVS+Tz0G7DS/VzimWWrb7rDMzxkst4ud5BaVGyeWLVguzBRSQ
GdiqA5KVNsDc1u0upV65V03EAb5EcImoGnT/Dj6fX9Regv+nOMb8np3fQw5h
NuGKBgNnqsl5bcePZBftomLzJmAksyk7L1Jpcn/nZprgYHqiDX92hydednb0
V9TB5HyduovtLoq9cQrY8TiYJOpvp73Vy8PMOMoAP1PMLohTR4bIqYanSfLq
7+GkahtCnohynpe0UtJzUbe3Qh4KrpPRtA6+8uJOVcjflidT/bER1LEvkJ0m
CXHwRQCMJPyZwzIej4W1b9sZJt0L14QkQaaibHprW5wMI3CiBVY4JTySFz1n
flzfEb2p6FcFNcvdS/CDhXKoarfK+Ffqe4Oz7OXksGnBuOd/8P4lzlwtL1Dg
QvkUH5aAlC2FQ2n4hLQ5s9WqaDF1orU+E8wCYAAm8bQYPlvA5fVvuh0u5m8X
7GKoxmfY+3r0UBpiSxl8I09KY7VGgJU0+omSpNUfyxtSCHFc0CLIFXpq6Sj9
w4UnGOyQEtTd9wLr93EyFxu17eLgqCSdjMsFPTcsJyuL6Jr5edkRnBDQfLA0
tE2LkY2Y9lm9y3yQQObK1KlJ/Qw1iA2aSe4p6gr7gURnX9ODbdPFOlyjfgbb
RMc2DMsX97dN7OVeIHz+QGssS4hZg4hfWxYgAlQKtWYonzjJIfnwVy/ZZy20
95s93zXQk7xhcjdORknPwYJa3ua/tDriQs/KqGSBpN4vQ5Wx7dN0Na6fOEuE
sDsGVOAo9GutoPr8f5IeHUrmmoj0tBPOw5QfNRUvO6Avq2MzsXZJAmdX3RyB
ckVR37qEmmmzoXyyxp6YhaE+5E5Gar4OAFlfmejOhycoRPq06d+/D0rLNkV9
k+h5W4Nylf+DTW8kY2ndr+kQQv+/nlsaKZY/nN4ln4i+5rji7USnAb2yG/uM
7Kjuf+nfyTZZqgrWx8pniN5bBl4fFjTNhXbmTAwKovhpO6iyuQBqybL+LM17
eVnd0uuJni81qg3uK2LYZbS4nV1HA5r7q4BtiOFI0L8CjkLzsDG7NFDVTnha
mczdk3cdGM8/b7y1OastTP5tKofHsPXeuwrOvpeNR8wZCACz9Cp7YaYO8Z0j
2n7e43m/OJiOslE+SNHsZHHUDURJXJ4xh+kauXDO0eWIj18MxMlStYuhX1ml
MTeyKPQ90ohojW0WXbsV+qU32W96YAg3Qg/PfxGCXFHuAqnwQJx15NPcErc1
cNxDkIuL663PQLV7L92pRvf14gsAgX7tnWr9B8ac3Zu/PYmwduoKxYj36BU7
HJagzcJro/qkTuwychRB0EM9lpZoolwLT4eywusbwAWcttRG6IBWrDDy9R/G
Kmn1HNxdjChOh8C5QmEJQqBe3mXexzwu/0O6+/ZKCDJrMowFalw2CeehYMSZ
lbQNTEn9QJrsaFxLFc47wP4D58DRvD3VpYbT8TYTFtHhahSpXSkZOhjoXfkh
fMjfwioHDzx6wwV6ivvVAHPJaEPA92FMpiuDBXhm4z42iWe3zMrFfXUQ9svd
igD4fNs/n0L6HIVVXiNq5LnXXikPNP58C3UKj6D2AmAJlc/mCoBDscm8uVkR
ZEakjgKw3dYpdHfmyOEc3KM+cvWi0ChdW9pypJbhX4amxM1w71a0MlXlGcTT
rUZzNPo6f0m7+g87vybNx3d5QWJ0m92kd/lZoyXIA6VpUMspjiIR1xfgbs+u
69t+BhpMpUarhtlrX3uqZSNCbV9g7I2FRuIlJWarUyqbDxfMoha8kuSpozxz
Ug9F9rIB96PrM9I/+TpGebPnfqZm5sCTmrhbpO+KQA5QRQuQA7vKWdr1D6Ta
3Ns++fE86dIvMxtJqA3JAGKFnt8r6RPFqxKTMzQuyyyoxsIEI/7+vzOVisjy
S1+m5/O4yLPIXCAJEKGp5h7E0GX8iais1EtnFQBQ9xsx2K7FOFhyDHdGRGQv
Y9Bxm013yqsMFb8MgG8Knr0HA+yLgMOVUj2GuC3QbA7SOEQ8zhgT2r+2Jnxn
KF5zmd5i4IwieI0NOzJno69IWBqLdB0ZZ+BMn8j9sVhD4EHnwSfJ+eqlP7r+
HKgltvgaUtuDwuQ5vMqLy9naYTRLoabTPlXfmPCyQ4Cz4F2HPQQueHpAgKA4
OJPn2itSpnwXQWMe1uQcVkj8fOjzXhMbWF+eJsLvy5IJ8V4xM/8TWKecQ4ow
oDA2VKbt6BLr5cAJtYzThDIRuq57NAsoyI//lgwgCzq6IL1OeEbspINam0pN
e9kPvC06t3trBI79FnnxVCFPww+k7NCeCruc6rqIWevzYl1Z2HsTaLQAzmaG
FHP5bg7UHS93Clu4JRFwz2I5XxXcAs0A1Krqnq0yQ/GxAvmITLLRPkqBnAUC
4ppw1cZrTy9OIhksCtVpyR/DwbeM3dCkn/xOOR/bOOswnbwCel6T/meeh8Lb
yw9QSkVq7204W/XWv5PES5gjzFrrI0TSFqXNVsyzKFjMOpSjZoi7+bAZALzV
c7tmI3v1e/arIz5g9apIXyzygLCljzqoJhFOAqtgJiGCplQ6H6CZH47en+TF
ifpPuSS4rAE2x4V2IgIOapqdgV7YSfDL0G5RAuzRp16SEP4KOlTK2JrkQyKg
Fd025UGr+J7r8Ez3+kOdZres7HTvk6UelHJ8vCpjy6SiQ0EDH4LX3+FC04rQ
aIfX0RoTBpHoqoJCZBiOdmoChOlB4xEX3CnfN+8nFYul9vgnPwq53LGzSS2W
OZZLdTsyhNfDO8s9T1mDsxQ55DM9drLNbVBcS0Wi42vPDV/BOQun3ZWpnNUh
9obDHU91MXFk+ny4RpZr3/dLfIPDNynXfubUaaQ22+5LLJtNzJfaJux5Ec6U
9gnExOXg37ehs8GfOVXuMfwRmn4UFH1S6QUhq0TPuxmgXM2xCFUqf4D0ZtL8
5f3HIfysm84kSlKGsXPBgZEguvMWIsZ62Utt/PA85/LF2ccOsEeVUbHn2506
fD50luKGSM2Zk6NDnPH3Y1/5Hj/mE+AbnW6uwA4pnTQGJyDjyS5QlFD1yJtr
5YxNflvCkSFFazqQid+Q1/KxAAm5czau3u5TWABOoY6KjBiJH2uYVpWqYk6n
vJqr7uYgMXlgjQ7b1HYlqpz9S4w8Xkz//0Nn4YX3ntmbCF7pbiBtEJ1Celsr
q1fDCZPTAfmBwHO19eLzLRK7B3cD3HeY7TFFz5NRfgAVHlICnZCp6D+a9IsS
H1o5rsBD0Hod13eEJ6N+F6YoUUofSyiL+SwsdXVFFt9qjEhQ7JzdPlbRpy87
R3eODzjkZ/8hNh1dEqZ4iihyx11EaL2zSQJnZprGLgR2rcw9Odf2lwKiIfaH
XqaDWZs/71SeiF+6HAIkSoieKF4Gb0iK3ynyltXE2wLJy+X9L5+TKuDp4DFW
WD61Y/rZqN8XWsqRDJH5tMlc6sjywwF6o2InttSa1R5M1HDU96WhzpS6dAEU
puKx2CjXJbNEye9O/UKPe8vS9EiXRTiLvrdHgfbrF+re3KtTvjB9P4ib/3A1
NkZgIHSPR9CYHx/b+7s8/Vm3q1m4j2dDdORNq0hw5cJWcf3aSSD5jT1IXBEV
2fDytoms63u8Yri8dkmXfUJOkKIs2n78v+TB6qzorYdrwttQKM7rpfNg9Bab
tHnsMtTD9G+ZB03o8XUAemQNp/+yA2boq69EqgBCG6I8RUcaKZiWZfR1AB1H
dMl+O+Ib/0A4p/VzrJebhi+8+fs7Ouv0ybkDWNanc93NJUakj7lltTqY5DiC
JoepNUeuRBm72eCtkgnhdfOk4O+1DN4ODcAF3LSZzN5wypdapQDTRf6Hfc0p
TQQkJ1uqmGZ/oZxAVEYXTH9TgYh7pVZSTr7ur9XeMALQSbk1h3aHxiliJt7B
Wxw2foLJ9vyyDQqdA9t6oZdydaZYk6B+PqB9tVx6jCY50zZf7uy+gqSARm/3
la0apGMm2wCbmt0P5ZfpqKg+A5VTmUIDKXuHX7nxycF6mW/PjCU/GD+sRRe0
JzYrHTnSIA+4N+JsRcDdZlYua+gI2hW16vmqNmDFrCiJrr4zCkn8PywIsP9Y
y2dQpxH9vFDRUms+LQM2uVjhMYTaVsKJTIBYjX43YMwy28gWgMZb/soLgmCU
pZPKvqYu8G528dMyI5BpJNN735FSnSv6YBmG3j5kpSGZGsgyUScct6vlkVqw
NTLu6WFrn6RPYILn3K05DNa4purbxbQAbfv5zOQdQaJtcpRIgIW7glZtMfuK
IK6KQCVm2ZHwkApob8TxfHWrB0NXOkmg4WXr4HNkRcbKFDdklWD7GsaJvNx+
rJyj7COV6BEpcaU1XcpATjXTSIfu7x9dy6wXHk4btlSdq2XlYtJ7RYDs4L29
TDQIDXTYo9I3LFHJvVQLBOHkWk3nLFgcD9f/hYnfi/3sDkzj75oFOXoWy/mv
8brKLkhaUYVy0nvWPBRy4ex2eWuZwd7v0zD0MZMH+gKH8016rx5VQfRR9xRI
c0YpFbkmikMTA2YeFuoAQxEu3nTqZChHWFjabsM3INOEQ6ggmJdD5DrFltOw
iaYBGe195YmL6H2NZJ4hLWcKtPrUSiA3oAYfzUIr73IEaX1eHTjQmanwG30Z
PPO5aNI7dodHoyC650jvx+XyqjKvT5pZ+REK5UsqHq9pYlB+7MH5OQXBdQcd
t8b0XoZhSUkP7UyXCtn3eU1UYVetyiCFZPgNAchSS6utMmFl3StbvoK0cicL
MCqpP8n+ahLw5kz/Om3WUki3ZGfFbdUyHoOCshyVkTfFDdSBUUEfZruddASp
lZGU/oRm3Ro2esMguPpqe2NjRQqajD0tuUIfi8d4x4YV50QpXexMjcyuFlaC
MMpAtlA3/mExYYy4F81hHQi7jfI0VOixliCeDJoSMJJgzSYsnmlL1xOKH1/2
eHBjH9Eo3rqDyO37gpLYVrXqgtmGB7uF7KQsv+T/VZLKXLBEXTwCMEhro4Zv
zL665yB8VaHOibt4EhEJwwUJveGKvIEA7cugt2wKTHRgC1KYl+ABed0+1mCO
3DIgjBCeHNHdFvwbSq0idOzEeUvlen6dSVo3NSAqZm6YovC6J+t/xCPmIljs
DzxmMMnJGPC4pZYc+pwpSF/Q54tzlGZP0inZAc8PV7IN7yfNbcsVzfEcrriP
RYoz/lXPTzeB0uGJT4K+7Z8jenvPKF5nAYtwHwDmWyrBLj8nZemWo2hnLFPI
4DzLqA9Wt136SjzaB1y+W3RBFRY0QaF0HQ/A9XeGnH1NTX37vTGT96EIg8QD
pO/F22nC0zPwB2BpnIJ8XRuBe1iB5sxpVdN31ELpyMXb3D8VKJPEBnyi+Pjs
eS77z+XZga0vTUvWG8hdZWmWxaTnCjFIMGKU0lKnAQtPclfQbKotdf+Io40X
ZbTRtzprISukP4XwxcUu0Cl/q5yaQTyDAzYXD3QO320JG7oNVWoCud1cXh0w
htRFBRdJlVS8pxWKF/XP9X4g9UFsZwA5FH2ryQrP6C+7cxZeXEfzLvgFof3z
UQuylz8ZIdAeCqA4ay6bGAlp5X8l+5nEnn9dLyosb99zUdYyzC9Eh143cFdF
97PFP5x2Eq47lvyZYBpNv6dduXUN4FD+BqG+rMnAhjFvtSPx9fM47nMvR/VZ
npX3abdyFA+zNDHC8fWNFHOpDizrUA27ni8lTPbwlys0F6YoIiY4WaGRTc2r
PoEJ9lmLXcCxliyJaEF6dcwEKHbPm4fcSefMKZSAqlELQRQzkab0vImrZi9R
zMJvRgYW81rABi5QkuuP8jEbTnM8q5EmBu9s2GU7T40XZqpWnQomr2MIiPmR
yX+0NYlvKSpRkTCFXW6E0WX+2cMu//W8EMdKJzJXB70wK5ypDaVNIw62FTyz
xr7QuMIKnYb0o+jZw3c79+e+0D0UsNkUqCAceN3AWgIuReJ/+ygaZWhRF5JO
ZaPb2O9QC4IeRrV3Pi6rrsfIHz0PzVHvNhAXzI2BOcfD/RbjJPq6OXksr2/4
IEvHGN3cBhRRHhp/KGYC55m+AA2dFDgqoJCjJH9bfyUPysr9oRiEgl+yQRA2
v1SoLAz6BEsF/f1hrQ+yncxHVc/vNkedfDVhysuZeriXmWwWpAoT8DKZIPCu
w1tiIpaO1otV65G5c5yW8+K7qvjsswAarA+hv+YQtOWUxdKGaPDtdVkicmpi
ZBvbinMz3VhZV6aXi5dH5RcISSseX9Sz7s5BEySpKR4jUnFdpt6M2ftX5Txm
h5Y26YO5uMmKXOSuBTEZZkMrgmdz8oPeoJVQo1ThE1clh0XEn5Xcw+MN3et/
DnvghZGRZjfbZU+Ne+oizDz1SLKlBqRv0Z6brqkb6Vkj6r289vkOGuseUGJN
s1eD7N9/2yzN74FUmk4Py0Pfl6fm5VdPvxUYH0nMWSpK79y8ShNNhPWer2mi
XugnQrP0A7IFs5GQil69yFZdSMypxAehjCUqN2G4GFtmAukNHVhQym8vSS7F
HXfh4oONwi1OouVVIhsDgpweOTiO7kmIFCUk+JAzen2SZi3i4mjaXALWzw+2
xuG3nJ9pp2SqH2572MiklDcfcPwJ86JK+3GaLMiU6IIaXUPf1WPVbPHyBJay
worEVkM6/3zptstWIcmIAROsBuINkc9BFZVC4jaEd3lkmx3lpHIU0vdHIkxx
oUduZb0stvgsjbw6y5rFS88pYXbTphGMh46gmyka6DfhYn54x2LNy5CZunJH
bD+Gfz8fNTq5xaZYMBtyO1ATlnZsNLC6Qh/kFL2BctUsnus71H3cYj+Ej/kB
5YAJlPMc70vprHGTtmdulMhcr5Kz8Dlf36qaQ5xCAL9aGyV3+mFljwQV0MO8
t1BhgVW5kfayuneYWrqAPrfP3hbSTlTn+yM+PPdM6CnPwWlVUFpHjO+FSCqc
FGn/w9edt26xtV4zKZfb9rvzQdznYlVlbQW76tXDfflnh3jAHe/RPjVc6Awd
NZbxQpsCJK1VFE2FNYfg92QXDsAM1YLG2BXd7ImCedT/BhQcwJGvaWMVeak8
FP0gnb1ALWNuTmMYhn5h0NXv6ZC2PJQHmCPUD/wDjhWiglxF/1SV50/axi/H
gingAZrM1XkigkW3+1sFfDwF9LN+byN2LyGmSLLm9W7K5FAm70Z2rPqOptmX
hB47zcIFyvvIU2Hk2yBhOzMyWemkWEyhD/t/2rIiVdKleEtuG9RQUZadQcAM
a2NNoBtreZPawzToG33WOKvvLlphUDlrWR4CnaUkSDvjCWNjcEn9WPtrsBcS
OZp+FNoB+C94YO41ofQ4GJa82eXAqHqb32pT4oF8QgH3T8yojtm4Dnxe3N8/
yQMzvp8Kp2bsXx/71JoE4Vsw4jU7Z9978UKrZGR4g0z9n4vN8JphqsWPOd/d
0SNybq/fVkztYaAW1VTTpeO/FvVHGjUmkQrTX98HmpwNKhY9bM+WJUFNMwze
2xgabRvT/mcQbjZaDffVRW9ZBvP5U4gKKJhDsCs60elpse26NyDF+2qiiopP
uXZ0eOxHIP2uX6LiFLUldzYWtZmghdXOuzhrPbVnwvT3EzREDdAhv9csJPIF
OcJdNvtc9Nya1PaVhWtXY+mdR7rypw1FA2RkdXVsisavvkkvdRYc2APCtj0f
4g91EUZ76EZo09mzz2z3YPzhZMPuBD3XXvhrcXDxrQVqTdMizgwwGu2OIKRc
oRQg+DasuKFoJtHM+7sGGGLp0IXEUNh6D1luP3d1rwwRfA2pTbIqzerRAZD9
sJOyjJvrtdemeV+Xk9DOS92YjsM1DJ9C3en4C5Ia5g7FPZa0j4w7eYOsJcCA
nrsNe2EyyIl1enMO1DzllVPNtFktlk84h+DfAG3Ihyf/iwHlxMvkM9o7VSwE
kL4msS5FEkKR/Y7sUMsnbWFMcIBJxzRzTmZVWAxwkgeqpToXzARGrgHn07qn
QL2mngF1N+SCwceACp1uR4c/MjcjqIKoEoGVFTfum8ah7yoxNXqenEYcArR9
ozWAfz4lBpkuL6qQlCaPyU+AXGHKA15kdcKpjz8HmToS8S/lkzTT7U/kWrk8
GcmSxC+Fr73+T9Q05uj1JSiPedKMviLgQVxSxZ2QT4n9QKoQN2xho4UBDawG
2CUqpjWu6juD8ZPdrBS1v53ET3dIW3wU5/xIAQdSXhr1oTi77f8Izh6y+2g8
ublgMEuDP2LC4D2AB3RVKDpOeJYMb8ZUtCN130iCD2cFrK6H+FIkLYwDdRrI
MCsgnL5LFV1Gk+8HqqbAXAkeKltx7hhM4MZacb3a/PswTSfs9jZNPKZ28PTW
pYfNvi2VV9AxPMSU1DukVOaerw/I9rtyjwpTwnHfoCoNK0H67fBSc/Yks7C+
/f2rkHKLe/sW5yVVwhkP1QspYWF2MDJSMWI9ldWRzkeMXfo9tiOiSgAgRCFK
qHKaz8RwOhhvQ2reyiFHY2uZufy5A1xX5ObOtY9sdIf8xM0OfQkAcPgBlMBo
pg78lZX8dEgE3BS+NUvGlSKUcpAa9TqPlGC1f+myXQ+jxInmkk1toFyWSOwn
BECUs9EX1c6V4TqLKX59bWXwcgt0WIqyTJGr1Y0N/4+orCeUeQbAgd7+Vfoy
7zYfgnCqWqSyT5LOqZaCOsuficmZWhLf0T0kDRTE5olitSaovuQic+p2ap3Y
qkYVtzPRwRJyKd4uJBjCVSZCveJAqNcUZ7en/0zkuc7gLCCmyMx1Ja9RS2xr
lEkzO1blQlwAHPmyG7f01U3s2XZ8FdYuOJANmbqeIlHmM6Fvj91qQEFRlDsc
ZxhgoF+PLi4cp9Pr0f8qzeDdKaXRNnGAyVTg1W44QGSJmlsbu6Ukzwjk8+KI
/DttQuUqJNeJEzYuf1d3SUY7c7qfc5F9u7Hb6M0rHznbR82PCU41KgYZ+aIK
DunPstUzL6ZGNB9Z4daSi+94eXxYD9dMyoN24LyEH0BGMyxPbyNwf1BUXMEG
k3g4G7BURKHbeOmMZ5rNvM79lpR0e5UtnUzXZbjPcauu2rS5bj1zika3UYtK
y25yAF8L4Qcj1xxBMkDuivsQ8sGS6tl4Z0tS0I9KfKYpQuWP7Qx6arDZrVBw
xae9gRdq90wiC32zTjjH7yD/k+8o2oTp/jfJ9ySFkOULYEol/Xm9tfIrA4LN
fXsjpMV38P6JrR6AmVX/hKt7c4RgiaSmxErjlTy7IpJc75hN9U7K6vB5LP+k
/BuD0M5A9NAN/FJqZDc97N3dpMQZDuPGIaJ0d6Xt5dnCTzN40TxwIH+E+H4n
FWxavzoe1JWGfbuhcFF3lt1s8vrrVAXsrXVAtjmq1rjc7qddf/AyU4mQMZaS
TFTM4qaVQ7XkuYDduD0SPAsmXmqpIMOJHDM1RzdtVpoWAEZNHBHf3HHL8lMC
B6E/5DS5ggZCtAPJ9t79aUMwmX1173m0vFi1PlitpBdTgSs9TONzJ/rXEkxR
3/rrnF4/dmeUj52NHmc4MebJmcqOQFD9JiNGzNFIxJiB5fnhZWRCMPp+tFqF
HdZS5u+plK3hSMxVnSp01+ILMfYv8wI4Z8ZQk2Usor4M8qBXnBmjpKwZA/8k
I184lxmtVpkt8gZ7OsDzF8TGEHd+7o6Ma15RN6FeUzg2yO/b3dyZmG/RZBDM
9fKYRbRVlU4E0MZEHhli8wTJWKfPnmu8m9AiWNvnXED8wKiLbpZSIsBNycW5
FPsFhXvXF19xT73uLQvRQzJFOmLsE/Y94L+3X+5jJtDrG9s+ZIqcZQrlpzu4
BpK/ndPc3/xGDjKD8Lp5l4ooyOC3Hzhx9BNkhHk2zuxUqrg89IkkGl2Ow/Z0
cAEZiecZpOYB8+WZBivP7KGVUbDuhuzbEOxch826+IKUYxcnNlW4njD3Wxjr
zHROYPDz/ZK1/HrQSEF7CMqu8QSB0YXP8/pu863Z62Q5vuP5bCRMNHvxc66w
VfJJDcnvkD0809dsgCWBsGYlZKNeVWH+mPXG54ptNyIKSNQDEuqRbtpn02CO
irAnK3NrUl/DOtEoRES/SdHoCR/GBgfmg6ohoSfge0Nc1qOxUthTptzlz+CW
1Kl0ioahyTym7Bzw0C3R86/ybPyPpDL9T0zHJrYal1hHFkvcpVWTJVS5MHjq
3CVGszcEXkpcJKqFB+WX4LK2uXDpjiuVmXCQm08ZKEfHJo43RbXseFYQlVY2
WhYBHwezWFniWSh5R9tb/dXnbYDGP7Sy2l0mUkjK+G/Dz3/eSLTSxkGL3N5j
RsjQk1rV1n2sLL3F3Ma0Z6JONAyxYXpyoktqMBsD6dmP4BJ89Nn3+dFn8xqo
77PJuliUkrmP8+Axw0Qz6Ix7P/caXHpl6+82KlSOgVHvRzck3Gs6MrytvSB1
ZTdbEEaPg4AYzewLh56sAy+gmNlTSijt+huS918p6z97VTfwFRKutiWNjP4j
NzngLRxbvpqsUodQPKUqRjWVGWFb1jaoOqMv+/DtdNZrgnY2ZkofLrcv965t
hrikSij6T8PAqNv6AbByMpMP3Wlg1k7+UR0BYVlVivyJs3U+PcjTLD46iQ27
hlDQ+9Jl7CjAY3Io3b1TfKLcN23c2qaNtV6Vb49Uw0KBI1M8Z7EIOBmi0eBV
OsCsNCZ5JV4leQMqpgLJWcOt03rjTBzLBwak4k+sEa4qsyL+ajb/cEPmXxmM
JHl9iO/SwZvAI1JNaqyQJP5xsuMjayMPjJQbKZGZfouqtnFXGzkUsJ+ODZTG
Pa69twp8NWp5S3ZT81Qiy74/nRJr++yMcFOVj8vc155Al0i2pY91fp0++wOC
3fX3D80WrEjSNLP4tvKen/BH1ogQzwNEW4bRjR+TukUR9juH4I1vuH/oN04W
KhMiGz/Xts+odqq7L3JJvW8Kws4tcYfLyVOFpK3cK3I0V/K9+4jSsGmuBro7
dkh7s6K5Il475BYgUwILZF0wLXDwXH8oXB9s9TGCKuAVJYjEgFEac7Eq45xJ
28ztq/r/KHFnhsYLDip9ewHxYN7NZNRwjaHlnEtlrj9qj61ozWbIj0am05hN
ouBfoVhbCz4Nu085QHJuTeMOI4dDQQK+eidpg7q+MkgvZvOqHFmW/0MpY0G6
BY5qrtytelRvFx7c9sajk44NbpcGmiIPI1oKybpMfbp7YDs/E27mNPfDmelU
coVCztsSaB5o8lQFDSXsI26RxZFEh1UGQ+0D0S4x2SWdN7+J1AP4MYWMCib3
S5LIWimvCr1iLK2CA+hZwBAK7MyXPriVoKt59/ji0i/ZJpBzYxKT67WkyqkM
TlNzYDZTB8d4JaJT7VF7NVeOKUPZhZdfU5M0FpoMva0Glm57x/mIjjN6BN0G
YHUilywcj+U5jNFhs7XIemRlqmbyp5ktOdG9w7Jba1+J77OwiV6AUt5NeXnY
WWt+KsYKg+tClM6EHLkh2gOxGh7uXGxFrQWjtgEGgCcVXYJLIbz+p8Us+pBK
zV8ccQZ5wWMYb3fVcFXWPZ9IdFjO0ktbcePb3dYb7EZktlQPZeWG9vxLQuJw
HAjTyCnVy6oj7PrFivaVMYHroDQFYJY3JxMs9zvEYIGLVQHKBSS687dRD9LX
1ozusBcxIuAO72U+sI2JowWE/kP19iP2B4ded+xyoJfKSc0OBKITazLEcm4F
zpEfzT3E8VafmELBUfEqY0g4bIhgTbMHoemnD4YLqM6uTIfkQ/IA8Ot+ru87
TT75o/DAXGhuAnhNsDcHRHt5rz2TwvJu9JeaFlAhVEddHtqmR7GVrLGuD2IE
5gA/YoKYDqmsTzjlZ8+jkjoSxK643X88Qi5gARYdOahLU8VpCrvB8vva14hG
ydab1b7mHsowiT+lOe8BzfMjpX6rvJgzFTabmVTl4XUfqX7jfj7jd6Xe8io3
FKagbeOEstl08ZVeYjIf0KGB2LLt6Lx8kdMYDQCk47C3Gc1J1M6M8tzGApr8
FsgWXdoYH7u+da1Ro385UvDa5FdyPcjN24950dMfVlJgD0pPwy6mn9nR7ZLZ
NMtmiUfVoOxYIIrOd/A1TWGcwLUZM537J92yD3cqVqEgVOPV20lqp48+gBjm
W2U4RgXVmCrW85kQ9PFkDxknFJGwopj3GQMb5QAPME+QevavzlJK/3+iFZur
qNa4+WX5F7sGPfWVkNWsBTibAv7N7MxjwOR9sunj/aPLD0kUaoYPwqiKvmZH
M24o2+UEdRcAnQJXNhAwedsZ46WGVBeluCipNH+CnzLADr/dV9hQfcaDeYiU
hYxTM9EdHMMCksUSr4rIYp2gddSzIhxKtRnbh/TzElxZHMQ4xOMA3p0jN/OE
gmAy48Ylb+NT7yd6r8nm+7T2E7PwlKYEH7ATff7eBABbxpZETHrPsTwJ00EV
xcxj5sq9nZ/3N+S32lgmIsRy1uXoSoQt4z9YT1n8x8kvt4LLycmlDtI3h2zK
gVaqqL4J+UnmlqjEQuOjM+1z6q2K+bpx5HKLS4DTcdk+BIR5giRdHbAsuNLD
dPIMDks6TOHxK4DxlQKXZcj5JC1y166t8hX7uAMrPd1zH7f7gK1HGHsVAbKV
r52La8esvJFFHHaB5hk0MUNhzFkApvJBv+KdUbwlG70xpvps+tt91AK8DmS1
4RdBi6q9oHHoGW4R+h9hxDXXg6sPoARsrMxMx7hgtKTkodWgtds5V7ybTJTx
pE6fI63fwSx1v8nikLccPr7Q1Kivoj7Ejo/GUCuXbMBRZD1/+690mqOVeESe
6llhgIIrligyqU8BPhwSWxhwruYJP2Ei3V/9A7G5FBj6DzCSyOZjfhnxSpBl
36sw8A38aJp2Hq5duD/wbFJwcG7m1cBfoU68ufZWLcsUGqnr7Bt0COz+aSyO
tF7fwhPpjmZxGnNGGAYunzKXJo9gWBiE9qxAXRU+nmU/3pYZzlsAGsvRF3Lh
4f9zVlVaY831STEY9ovu0DJ/Tk44O74Tdzh/0uyD2unTCnW21XCburagtJWP
rpK5t+XPJXI8SE/05swcKwthgtb4/xyVOAW9bHOxVOAIFWPGbZz7oZ0jrNzI
7p6Z0kfX0thO/2ejf4t4I1YQsjL50gArPrePTLy18/UxOiluLjdJS6sx5Jxb
wi0CAx3yq9sloh9ftj5Nl5G7kKlQ1hg7Jp+fUFCbPs8TjfRCEnR8Dtvd8AC3
q5bIZdUwgfpZKTFgl19Jh9esT1UwwRM3t7eJLhVf/huaTl+Oca3rj0RD/318
mC4D/svAmI172rxKaNn+eZf7Jmyzm3k5hYreK8ONaJzG8pDp+s7mKeN3syzF
ocRUGhy0p3scQTfw4lCiXWACg3YZKnLCUbBjx9Fs/G4TVQejn4E1facORs7u
rboVCmvSpqUT9vOeHB6+ycyk6aVzTjKFhQ/ORZ43l/BS0gnUQNL0XUSY6QCQ
gNpsyCTTad5BQzGm4AY/5FbviwfDs9BLCoTAfFmR/ecsfNZ6se/B7ISJ0rqH
CsmPS0zrByxvWFX4qrRDieEO1k6yAsc5WJA6My+YxNlxThU6KPkzCOKTMlHT
YfwjZJDpJQDedqdyL+5lpuaRvMn6u8dgfsl7k2vqzNwEPf6wlZgm40qGtWha
kF+V+ntAB7VRNSnTngNCj4hJV0BxS4zOeTNVly1YzN0DSFc6nRN38sgYcwub
Pdx369/dqz8SNJ2BBrBL0m4i68ZKGWjyWBGrFfxxX1wQ1P12mA1XEvKAkd9G
dqNl3cWjI7xNwB/Zq+r66ek3M+lALJg0IapMUvfTN0kBTDtm25xW0EdQs9M4
HrexwPqVKdIk91t8UHsIWoGkp0W6hMMAeKF068QAGqXEQZvyFnA2/TuQs4yc
4TpW3ns6OEWFBHTE5Ujl0LVlDTzMcjv3oXI39Sd4zNNYnFV4tVbCOTx1MgfD
9qOyOJ9cRRJCvrQf/dPnWg6//hcHAM+jYHXFDaJRpxNlubz/CETtQPflIeh6
y+h2DFR2AgNCI0LZ5E1dnJt9iiW+nLJs0ZUKWO3lHUJWAmwjrIspfbYeFW+Q
dJdia+I4e62EQyqlUAWTZn9Utwc4cLbhKHEAIoCjjemZDuG7xcZwYkDoUowj
AnhZDABp/k0fU/rdQb46KRWYCymNP8efiEzN0mXr3COH2HSgXEq+hlmcPueA
WlCWHZy00mqjv21M069ZL2utyzyB/h6LeDwx6J30g9RwPnQdgCeiwsDum3ht
D6+i85wkAuM6TwE9zlVJvlLeb2xF695pg8PMOcQcT5y+bV8ZEWfhfZ/xnnEZ
CAHQc8b8g3j9Q1iAoneBYxj9dnKPVNWpqGJYsmd0tQGcSjMdpd+UfsZNF/J8
hwaKbTgHl0P61f2hdTNFj9udrIl1yzH6Ow6/oxJHjNKOQL77T1joNKcG1MEP
jJ2QjRlKnRm+bynwoNpvGvfpgSjSJHaDNiUV14RqRJ7hGfdoyborieCR4cUp
SBta/Ui5Bcv5qNlLNY+bxtSOe20z67eiY2ugUQf2+EHVbAo9fxzEb2YDTtJp
Tvqa0EEWxTsqAcYkQQOjOFFy09Xt+9r3rHpvg2/+SmwJOlzE0AGKAoHjU4e6
GnqmNEEwNPpud8zoLiYlwbeDABdh/qpuYeMXI5p/48igPn+2ql1gTSkJ6NU7
B/Ye2yNL/3DNfzCR6Ff6odvk1nT4Ffhl/LJjCAH6IT4hljeWOd0oGc7Aw21z
aqIRo5NW46x/mdIJLu+dZrQiN4Z/WtpNEyPUQeRYNj+/TTglm/Z0+3lsN54O
XdBo0uhB+zG69k6Y1RlglyAHL3yWOCI0mtcQmptLyQjXBQ+askcM7gK0VIO9
MJUS4EWDSNoN4P47Q1LMMdL5ppayv+AgNt4Lx8uCTGanYxuahg8CBjgtNmje
OJncBeajF5gWggjIAUhJyukwaM7lDpkBHUD3j4v1/lhsEw6hF2kYALpJT/NK
E9eKCUl5/oAifSbhB99RdSApm7YVkBMFrhhqBvLlTmekUpNJczz9Jyj6xmJX
MO2EV2e9e3ro5rux/5325Lgx/f/6kRFIXkhQ0FjC7terU8cM07Lh8GP8sYoi
VcvPVX+zv+W8vmgB6rgsZcfgpQKN9VnB/7/Qt6jz/zeMsf0p01+3ekBI5aeW
py0O71MM2jTfJv2vwZkSD9FC/JVG8PnCctOSA9TMjoRtDPAjRUnAdn3qeMXJ
11GQnUuw2AtLZ2PlRTDJZLQ3FVh3xsj22Ba7OONxwBP22iDiVYy03EOJzxM6
sghGzrw8F3SFeepojuJHm5UkiRg0p8nM/qLytvBcbwVYTMC3DdH1EdSY1gIi
MZiV/Htx69qZdmRht0Z406R7g9iTMT6X+Jw51Uv84DgGf97JUgioOuyarcNL
yLCXoNPUsr00U7fSZA/7k9c7ZO3va6uQ68NPfWUGkcyxMLIeggHpMZmZbMlV
Aw9aDak5jcFdMXGAsvPcJWJr6Nn+5Izs3sMkYE6LNQjlsyFHzf1iI1UCAbwD
+EQIrtU4zjepdBbZltyU6hTmAdDj2Dnssomaj3hFACYD46p05R7uUsWcCLLb
tiSDM+pECkKf3EGOaMhwaqr8Wk9xw6u9Vqq55sbqzy3/wN4eOR+ynxkGMO+A
cmIYLtp9s227ELCQJhpayiteMfUlXz6vHdqUZH5GM8gBQ2kWCiVAxIEfji92
8LvoZgsXLaEE0+TfjEP8kX7tC0M9qV3Ry82JUsdenm+a6xZ5DlosjohmjPky
yhzm0AY57Q4rt9S5zWdr8fZ2ZdszStHjstSzpEVklU1a/I1J8822PUejLFfQ
3F01HeUzlw3rXf62KGKrm0B6Rj7khlznTuzzo/XHKuv3jKiT7X1PMG65XgPA
4mI2H4rbJGwf7Ok+sT8hITg0eMLfTt/tt47iKMvc0LQ5u1PC6K8pitipupnf
Om061ZFOBxUMqKTBJIvKxl0dcfvHCKu2sIHqVEixnBJ305cEBFqt9j8BKwVM
GYBZgHhz26APrPYqMFeOo/LkBpsTDq/P9W8D/hNaPyllSDywENA7ZgNORvhw
8q1cMQIix4ISWc8fOOx1mqBoD5i0RGT3mvXPp8fRAbwPsjKxb10v4bM/LbQm
AM0JuqFfn+lvuHerFEy9k8c1N5XZHx7R4bBHOmAjYgeCKAgS48vyxzJ78GQ6
ITppIMcLj1+ZjVGBf6/mh2eI0B2NfRekLt8KL6KxRoRgJmX3Jm/o9pySe/6O
/dR4RezDHKi70wO5ne8sQwk71jE6cclTrlNA8GdTTqljFFCn95c2QtzZHM9l
qDOrSFC8YItlw7Vh4iq3Eg3p9g3OwQrOf0ieJoRdKmGe8FOn3U8u4lDBfuUd
1jk6ZA+Ppi40otXLdhTAej+TLM2aFljBkNX/TsIw+ZG+8FkiKEPsc3W3l1iC
an54CZU+IjvAWXvP8/bHwMVNcCwudjLgPHKZaWefpm8WGJ3acAyUDF0qhn9I
0vE1RXwamDM5XZYwn4nWeIscPjo2PIquIWGg1JN9x4ZgZbe8WHjjVJfa5jfJ
lWii+9YMDc+Vtb/IGYo5reP8vyQti8ASKTquAoyWF/AsVvkSvncSBCSGfpVA
FusELodgIqnpM+WohDc9whWHLWX+PYXinlGCgxmYFMwWVXlcbYCY+RdM6lQH
G24ZPPi+MUvNhODUuxx56QjoHTYpGE+so7B4QlV3SsBKSzs1PB4cwOtVKROH
zEcHvrbrUs0Ub9gcV62XwwRdpNVijcW/uDMpIJf0EGlfeCIpLW/gLdFAcStN
g7LX2C44HNr8xtdEh+a840La03N6+8rlUuOOXH59XyuFB0wY6wd+WDP3pW5a
TlTX/3LCdzUJfzM2a9Zmo4tTg/8QYr2mE+4MahDLEOFlsirG6oG4QuCtdnBO
xrjvbRCfAlU/MIrY8lXi/6crnx/1YyD4uJUYyw0v1hzWmS5kQ/Exst88x9n0
fsQd+XaJqY+b3MPey7qQ96yMx+TcpQMdr789k22U1oDmitINZmgc1xqSwlwJ
8icPigNXbAhR0NEZNxZ8kVLqNvzEgvsefzFV/nSjtIUB0Sfk48jJV4snzAza
kLs4nFN0a8yvkD+wa6baob4hkn7zo/FIoeRcs/lllv72dmueihm4UVKymqGw
KOm8jS/2UOW/RIGrW8heCG7O1YC3Qwio0Gz+GORDpLOWQ2bLvSwQcUHZHr9T
OJR+Lxx9SpjPt01dkKwUyzCIXw1oGnCcHAhjE4TA/pBw1CRb869xY1FKdhQu
sMssK7oB3eziRz+7P5s9GR5BRWJCX1KLhnWev+OPGxzYyjwkv6Qp8t1CG8kk
D6m5W3nSY3RntryS92rx1995HlfWm/86nAHCl+0unBNz8KfZkvji2kXEEB5p
ybrR+2XmH7qd2BbC55tcj9ZEF9xiwocAZDZplHwIIE6uSvm3N0kMXlq0ILKx
bvlMKWXyndml+Z+ai8b0s58WBdX5vVbp+xA3AO5J4IUg4gu0lHsP4jCbcIDv
S1uaOy1q21b3SFQjuBzq3Ph8y72yN7KfdniEZi7TZnS4jaHw/QCbmyDz6QhB
dp75B1OXsnNa2+DYD1fw8OK2zCXTAWENU062GPMHT/6XjqXB9Ru2MPpWwN+E
tfAeAmaBbqYbtU6YP12o0DajQ5Ah7qNJkgSr+vAjFmFsEZboWa4M09F40/mX
1giIGerb/pW3xx2MjL3mKnxNkiKHm4/zHOBG2OBg2AAsLBZ0AJNWm73d70qE
/YipnoJQrwFWTXGPL8nJdgTBT693Kc6fpdyRER/JbNhUCVe+6r43GbkMC7CU
2NKIrarvPjqZ4uRHIiEQMnBfg+WucdEtip2jOPMvQRQgtcllDnfSmFkxAYhN
75Kse9K2hJmqZnGhGxC+Hldzn4+DsPTR1zB95FDozIizq6PFn1ILhU0RMQWa
ALG/YXHCBcr56QZeyibXhUrCbOrWbAnLch2ms7gvwW8X5x1ZmQRkQC0SJWk9
WhIAdkqqreoTi62qlrVMa7a/y21aCmQ1F6uu/RyUZrZddyzM164wVWeKYfhM
uYKs4o8QjNFCn2IWVmJkEN4ljqfabsf2qZA8QPbqFNou2h8yEvbVjU1iNOhb
DLYb4QkGzJ97uWw7lj2sIbzyP5UA81G4dZtZ8kDyX6lG8OuPNr53dFv9WFFC
jh21xPaR+fgnFh7fLaEg39mzYanQY9LwmVjz2nnHVM/J7TFZTrXyMs7juO7U
1AcBuFpQTMDQAaJJn96jt1f3dRp5nvPqFw6g9noeSNCT8PYU9gtMhKAAZFl4
1vyjdhHTT3rfYB2na5rjAQ7Ug7wThdtvjsg87flV1jK8IErvSyOmWgJtG/Vx
3wCLB9+lItUhrrssBNOrpwU6nZ1pkyac1fApIAlCPheyZDl8vVqiqooSzafE
GRkGeOmMPBgCg75EjTJIKWPFJP4tFqa8sWG8RAMYbGakAbTZflMg3UoYbGZA
x0iipUhdKNqvvVoU9KgvypjZyDnUKJreFqfqkOO29ad4VlNdecjh0YXzTnzc
2LFwMUh/hD7GNHZ2mOxpHOYKL1N/fSO/Q49Vgvm2KjNOTpxXflFzyn2mJ1zi
KC6TuZDpuhVztvR2Za23zc19hfnJTwdCZ+ijy8/aHTIpo76k6zWaCWarLXKt
a6SEdX+/XVM6dAEC8P/wATJmzsTn+2Z55UNYQ6VbpYjT6zDLPqYcdujTYA7r
ckQcvbTQOQeTiiZaKUKrEd9aEp+aNHwzPT2yeZHoZbn5G+cdIOUNf1xu2M9Z
0e/iCKujJnHOP1JFG1a5lv5Y52U3yZin/6lyJtZe8PJ9rGQ1qFpyz6Pwk+3Y
7FIVdn9L8b0T22PxXjltzk1S+kYvO4ATOjRYVPQMsFvOyX8ok38tX48xPdrK
+0S3lf47PIgtbpiWAxoA3mnDR67fk5EeWOyHSK5Cfz7HmV0pGAaRI8JLNk1b
uCUGBEGviWK4dsApjAd/meAlV0xvFrQZ5vw6gXeeu/QzwtP/pjGcY15e1i+z
vyKzawQPumG4IKscDgNjUEdYq1yNz6YyhYk4eO0X69lovrNEkBu8Fq9EsX4d
MfQB5wPewODDiB+E5Hs1z+RN6cejUq7685SV8BTw/GUqWbTKV9l8wqznsIRB
xIljFFLbdnC9G/CNBPCf63AMu+0xNJPnXEGcPheKZA9EUXxXy3mnjO9+Ezxl
e+hRfXW1na5zwHOLBM0WIeXioSoAdOWpUU87x+cSyRWUijp2bykYdqLQaOkt
ZIrRq1lBmWpmj3Qx26ZrurOr/+LgZjMoCjM06p2kBIAE5RuBevKVALF2AmXm
W2F+xmTINi5G1nomS0w0jhFndFPXi/uZ9Ssqdb2al/khjN9XZVnkMphiUdFj
7/msdH//KPGd5tHB8ZmV+NMp240ieNmF2ckZEaCeOXvFDQLKjxgGEdkym4qj
wC56zgLpvi1c8vbgtCQKEWdVvmRPo8GxXa+nxNjk/GrLNG3LI9JR+Tnw1uET
l5YJ2V8+bzsE1PQQE7VKaLPHmzaVaL9434Qs7F+oTtifiWwNVfvTPfAtitPf
abZsAQCMos+umDdPU4t4BmT9nlekXXmZHLoxYfNydaHjm3empWQhmhEe7zty
iHTDBsMaTORff83Sf58axEXsrznzQj5EIrvOC3JaOC92rmB7jsWA+LHjeFuR
avqaEj23RcR1oBxDPFTTNdFGV92FD/JtVkSDEvASG4l6QN70wqJQOgUdhfp4
Kin2o2kYUBnkD4XNiciJ5FEM7gO9aTCUig0TNAbGFBWVqSc79amE/Jr2yhs2
1ZB1e9iAIIcVEb/DXpdsqrGCOY0mF3Kb23Ccb7QFKbYync5zCq7TXfhOr9bX
GzCxQzIYpzCDbieP90yOqEBT1Lvm1IyMC6tMJJwNYqqnI1AfsLL1Ir09TJCQ
Nt2o/AH7CQ1UvN7m5hva4/khoDWzuIGMHcjHZ8QOaNhV7nSjAlFb55kdg8oJ
x2CWHPNhRLY5b7r5KCvigzciOGLOIUwEpX6pDjjwP/NGeuzgA0oAE2Rc/by6
MDWInYuXYP3+eb3UdXw9nH4yuM/GnHGdncxf6yGaORK9nlsSTA8Reu1f352Z
nYm5/8eOcVVLME6hyTRfchGFHFnFKCblYKkxF6MrWfDwNSVJctGqxL3du5ct
i27n3R3hKwKcAkkE5q5sc1jofZvAdVw78sB6vzEVF+ciHwxOaZz4GxmcsMdt
IXVCXIoW9PNi3KM32lgeiMbfJ/UTuXGNdQbajn/MEcAJWUwpYiUT+J5o/DUF
PfEjXun3+AkngDitTdU9rQoIPZpOhqH/cVhwcjzFYaF33KkxgoJ9tJEMa05+
HNK1cEsPgXRm4of1os5hjX9exG84RDDdSpVpjcFG5JmTj2B3zR456iMa6iqQ
kRxWnUb1vffZzQEjBI14NfO9xzl1h0EtAyAMt/bwZA3LytS6Z2dcgBz270ZF
lTCDdBtWArl5PplEy4wurkvR5e4hIVOJBqIqEDdxz6PioqjQcHICoTXbvnKy
QaQ7JYgedNwnUrAuxIa3Qe9e0/6/MlbjGnDOiMqXD2Yo4guujZwvuKP78czP
mn5uFbQswHndcJUuD2us0AaXlfgDbb8xoUr2h4ns6uPDa4YV2GepFMS7MG1X
tNPpY+hsUdbC9ymNDY8AxG9NRmdZ3UVL9Ywqq8ilAypj9c0L+UpxvrG5leiN
WF25kD2+5aAjAHTfShnFprWArICF7xSYYhAQGyyQmV+k6KcfKV7RJVETPCyw
zLA/EQ9qcOnYduVP+9LDCTXuft1tUgljH071AMO1UjVkjb/BoHTnhEF2nR8X
LLl0+Ld73E5LrpwbulVQh4SL/rmw+UilZb8N78pnNNjWNhh8QcXqshFLsj04
4NFHTcRaQ46mUXWkMndzqXfRRtC7zHzkU7JnDItCfCVx/UstP7JLbnF0vvyn
tahCnru3kiIWMBpllDFXfILzdTtq2yv9QuB0l3pnnbfEc5tfqtH7OWwwMm+I
6vKJEXVCoXyn01ZdlRh5hDeC61GrvXkg7ZhVC+eMh1Z27bX6VNcL3oxgn/oo
jhr2gMWr7cxqn6VXVx2VtuI6zabHTmdgmLk7+B29y1Dk1zSZ3CGkUi3gil6d
/yy9VJAcGuRg3qgVELMwARdeow394mMHkeiYLuyr6S7zZNbye1KmIxO14l3g
8fi+Skw4yEoAsjqVrtQET2JOJMLnI1xb0y4B9FMhBRRp7bWi6XIZVNrTwy5a
8ZbnP3z/fTAyiJYRPi0jlydCSis2GHghbsNp0zZzMOZqlPtAmWgfXeX1u+1R
HZm2jpbNm/2vrY3/yuoReeDK5OIZLXW3vDnN5vkvSoBIUwA2UjauBzhHx4Gl
4UwGJqeyxeIYi1Cm/Q5GHiYoP5JTDJiJTdgsR84ao+wazqiKvWntZOnoO82f
K7WL3cmNFpDom8KnjTaCrdMtiYOhEXTMas/D9l3RNoZ+JxJvlRzmyw/fihY1
cErZhoOYAFQBxy7E6JONSlwa3chsuTnpwNzl6Dqn6GsJk7QWwsXwQ/3Yu2aZ
fXDZm5Tcfblh4m6NyaPXunv8nknZLdiKN27iv2t187cEDpf5THNAtK6qovM0
VzKK4llMT1tP3r1RbOi8ML8tje9wGG6UDXUzoTYef0Eqj/fPaL/zYNpZtIwe
QfGKFjZlkVLsy4Wex0Gv/QVinaHjQRQRuiJOewlE7ruWSF+0VcOgaYhlnNeW
l+bHGRei1ePmqm4Q/4fUNdo5gjgTnJf+6vhWEmFuuctt4Ou9e5mnDoIkwZYc
gfKvH92fbcOYnVwdbvyZgA1GnSyR4V1j83CK6z26hP8NuuOpPlC9ENiH986v
3cBVYQWGOMEq9BkxmkQCYilhFMxhsS/g9RR3lT3nSQBbbtla+ldDcQ6QLjU0
F/nmA4sRhrOl+zSCFVD6Ki1vjZU+R5pmL46WjZXc+S/mt45eb0PdMvzvT3bc
XCec4KyY7wPvbWhwO8MlaPJbsZsDwRZdSs+1ZzmH5ftiVR/aOJlnaDTSVDL4
j+vcD8Im5LiLTUaU10//Kg3AxHmgDYQ20PCrr22WqSVv/I4GCd4SkqwA8kGp
qnyj7ryJ8lPt/AwZ6QWQxEW/azV8vEN/OA366cT+sdgE6G2N+J767Re1WVNy
H663l5J+pFjh1IA3ZXBBnHv2Ri3yP1ALXtYEj3Gy1bozguLI1MhXeeGqI4uD
MLxZYmynnuCKU5EUmbwUqhwdmVMbqnvN1L/nIMk9MF5QqzywnBVsb4SVxwIB
TqdHZAbsIonx6QNg59OvbxVPu4h4lDBdGIoA/H80awl2yRcHEVdTMRQ+ISsn
vpucCm4CPzE4Sq7q/0coccJbXE+RXa/zOLp9FpcCxCXDZ+oyb9LH3EdusDAj
4dK2i0tE5jknPUZ4L+ryI6Y9KSmekgNXTEdpyKLv4yNXbj3exIRQOXnl+jS3
nL3BR0/3g06P1cbQOpQRQj6plnq+Ur3F5jemOPgKo0qpfK0lWbhqEhrefnO+
Ls2P8D3/0l6mT2hr5XWDfW6C9sNk5EKE3cvba6OGJW24NIauOFoG8B5gjbbb
9zhmY7sY6oJhHzIqoUWlHsfF7KQnA+oDWVgXCCD2NJoU7z0nD/3C5bArf0do
3U8omSNulHnD0U+wNbxmVw28NCFGTY33UcZ3jH9R9fOZGrUNqoqd3/F0arCP
GgVau7TqL4sBwWBUmA12vh4KHOs/ZjZAjbE0Uzz2yXC29uFLimwTspDcafi0
s+yzItAAmW4bbg24IaMOLNmGOXrvagIdNYfTKAv4JB8G9+sXLcZZNdMTY4f0
BWBipvflBiY4WNl39HdlHO0u2BuGry4aSsAUmAdyTJCLMhSDJwrFfvUHpiVG
SwOjGNs3dwaEr25/JfWmF474vx5A1IDdPhUe/XvisMJdiWlmu0kYxtzWgmsj
OZMSEQR936cXQ6NKrAO95R3Hv9T5XY325ZDogoUfSF0zTd/umUexSCvqK92J
AGCYLZjL78wuUIi/3XozCsfY8+BKs4BPZAYPvuXkJl1lZTKKsYiG7Us/dcrc
ILKtN4tdbs6hYjkXmVyGtvWSAnyaGnUWinFVZf5NjU1gm+rNsHAk3lu9hH8F
uGUXIjdRnLj5t2xz9EIaNEPVcCYUGi/lCCfDK94z2SIGzaEZ7Jztv06EKzDn
TT5BPLbbfMAcSIwb6hxEFPYZu8rDPPriCxIUHAdp4k2TpV8eXrSPVZJXTNvJ
qihLNlUk8VrEcxmxRWo5x/RAR/EBvBKOr4jnafk/8/0b/alcd6JI9Rzr9k8S
8B2JncvmyYVPC6m1hQj2sfC4UQSIgX1CRd9kBtT5NL+YSUM3zi60Brn/40V/
/emqbDHJwho8yN9SnwkuFzMe1WFgPDG46kPE8WD0GY2V9I/e8RVjNX0R0vC7
f1NUrVoPTHWBStUkrSCdLgUPOioYjSMTleDGk+hU/UBsBDNClFwlfdRGJYYm
JVCMyxqSSj2un+kO8E4ZZRnRSzgVHj1LE97JxWna1EBUAemnwopj5sQAA4vP
B8gSH/UTLDO9wZzsrFnTSWWMkCsZ4wPLtcq1qjPwMV/wl3J5JN0t3ZPpZkLj
Pf2uEBsBfUrlP15ktWkQWoZ68k2n5hWHiZUnAJvWIMJLVs+zyTwr2TzO6NTj
l49NVSR4EuKfw/L80fZT1/C0yEF9ZVc9hQztRBeL33HG2gOBuqkJw6vtY94M
hNzkXhspbG3xgAd9ducUyosWXq43HgTEr8oPOBlcgrP55H39SUOf5F+Ub0GX
OBS/4xzr7vaMsYGt0otHzUPhDWkHD4Trhy0frBqypm2Z4SRq09YodlzAqf+p
JweqEAAT+Guhl0FRzlK70TKbOtaR+eEOTv+kPiUZPuFBkGrikC5jb6vKMaxy
AMesFV/bs863t4xORyiKcmxSirfGAt92kxqs0z1A78XgiIRth/XiVilaPziU
aPLvm4oRdQZtaaFmNkD7vMy9Mj8Zit//hNc5Q3rtQHYnvJa7IdFGtceAkaks
MoKhcJWHLMJ2Qhq6A2yj+SrvJLxNr3C0XexcuX0h6aUWPSqUBD4jf5jRubhi
B8ECVjBCkqzn69Z8BlNRhq+F38AuxYneqOMUDEe1N238ajeOw9SffM+0Kaxh
Imy2+5+ZsOioUtEUA9gLqE4HbYJQeOpRf6+K0WXOydhjlQY/lGPn2G7nKKi5
Bg4qgxjOfniT7xI5aOQQ9rpuRp+Ew1QmN4en/UtxEBratgiLAA2CWfj/OxKA
ekHqj21/xxoYFP0n0fGYcoE/J97bl1MCkf0V+39B6izEFflbgtQHHseTGp64
UftnzUBVHzBI51iCWzeQxOFwLtGAbB/p0xmYUgMi/m5lVB1fz9klNJNAplMs
+wIwKX8GXjh3yzBENWudeE2YZRWhNSaLTzFlMbjzUUPaDQzIhZBo5uoOShxI
Ut0pI4TZNwQ7zKWtdgZBazgW5oZlUC1p4CLwjFYJR8tCJuis/esmYwX7mKEq
wyOtAAi6oMkGCSfc14H4tnj+z+qAySllA24SKvPzFFtX6vtz4oKe6voFNrFU
M3/CySB71Ow+5rC16FtRg1yA6tgi2vZ9PNdGo1TDRsJ2sLncJ9bUWeJ86b7Q
J0ezcDbQYeoRRgV/T3fn71cbjhjLlVXzn3DiMN/Tjn6M9gngT7dUc+uWEAwx
SCh74puyFkAnsH5vFiN4Wsa+jBBmfZQ3WebthlIkIiXDjgkNZ8zs1c3v/uMs
5oQToNIYOui5v6uy3Bz2y+CsSwqLsP394DZQbV5cfqHZUCJsMVh+EQHhw7jc
0jNBnOQs8UOK3Pu+WD61GllZzzTd/VWcOKl1vUthPFwY5FAs5xYLMjnqeIh4
/XfAU4aWgmtCZgfw7T4pkOMibkK6sokJ5DeGwBI/Ac8hNpKfz80H4zbH2OOh
ZZ5NroMq3NiqXmjrfu1wJHGujg08pO7FIT/+uyuA33i77PlscLH9D6ogUz7N
LtxjeIz9kgjUbbTBxsAohR7I9O1cY0Tj7Mf9K2IyC9o7vra9HtFgvKot0wJ9
zreUyT+6jHJ6EVeGML4sc1361qbuObh8keiLy3s0fDFFGEvvW1HbiQjBbFRv
Rtg/3MPwImLMOrM53BvJYgFAhb1/f0rs18iXmVUaaeEtgXcuyqR4Qu5Pg4ua
fEoofeWfTFGrp5dOV44YskPT24R6uzJoNgXdHMpD/uxfVxBFhkh9B7yMxQ8z
fR3oGv/fE1PDrvqd4k5ZAzDETePHJpbRY0f4dINMF8CPeigoZaHOs0M3ATwS
NJzk/M3rybpqGGMdnmtEMWMjTTyWGvg65kyKmS+lIca3UrKmTJx/PWS4Uqdy
h3M4mCgyFzYLS4xenbl573C2/bxC45jRqYu9DubIUTsUgSMoW6YAhQ/zgECL
j8LqiWqdbDW+DgpIqtQqu+cNKS7un6NzuJRI390tu/nb1AfONAQ3e/dcu0I7
Ri2TgfnrktmSV7wBSbviX7K5gpewOENc3hgP8miUhp7F1mHIfIAv3vT8vD74
MeTYm/I9JjY7cccmbz4skD9xq3GJUcEgX7OQmuOrcSKQ25Zl1+nFPURw/FsY
o/DKbEVnjWRTwiG24eRUB9gUNijjCsnO+VDa80TJvwPiQ/Hk397PozZvW5Jj
uAsYyeZlzLd/zmoJOfUf0a7qeORQROd44VUQDPvvON21WUqczKlsORnU8QVN
t2l/uV9uB8Z3PO3Mj5fR3JG8P3+TQkAer+MQLehyfAQKQf7Pdt8GWcb12Dw5
KrhIAype8kaAxg/T7IApaDQRyH7uJGX8wUYoLKa9DezzMzdPWQgJ6haks7n8
dUZrnWAj8LaVE/9GqnQAkorgzakDKBgLi+mNmIdHnVLKHYN2WBSsiSY9xrK9
ELQGZHlrQYaUPa6R3SicJUMl/yEdyfXzFALiqmC0EQBd9rsXuNiWk6q3mzKN
Hw5x/xS7QFRxfLDcgfr/i51V+46DRUI4GuRnxtnMBGJMcDhQh7T0AAjBSlZO
oJ79zwFOyb5DSqKAT7TxrdBxo3Gy/I111fJ77TwhBgyD2tCzHyWyutspg+C5
KCce9Af4gZcjr13RdHT1NEzkDUJkqaENvmFkLEcRzl5Hu73lJksM6AmtMirO
RVQGAp62KXpf2gl5K1/CyVk1UmbPvJ/qIYG6ZVsFIPyoLohiQ7FtyuLbKcyD
FrqG8dVAdLQAM5BMlZHNA1vYsODwl5kdwYpYp8DQn0PLNmfxA9RfAy++Ygc9
ZKa4s1o0BKjt86e6aZxfZBHgRcMWmzxQ1WSJBDpt8t5johu+ih1ivRCQZXk/
F/UPy6ym1yB9Bx9N40oaGGgjCZSpe3Oq5yXoyPWU7FYpcArQytw83BE7ylG6
+YTdbAx7Lt61atdR07H+2E/p11OumwfeH+qMm23ZWSPf1eHk/nNxcWbc9nlg
gSEj8XG+hnc6me65rgWDqw1iDSBkSf68yx4+WvNXu0fMyvcaSHmXN6U/WtU9
HJ5kIMDu5gubuA/PwwNsn/dHoAxL72RtTMNxrQdQzoHjjgIpE9NderD4iaID
6qYWjIHsw9DkCmOT9FzkvsBiseE9a5GMIur1lGc1/0HGtmHFV93HJjAYh79z
EqsfCmt258Pdu/FrnJqjZarykc7br6dI7PIFTVAax2oO/Ukrw4AIaY0yFHEC
NDb4CcH3SqI6l1oSo4Lp+00c2Gy53xsYVr93BJozuCaQS7VX+Lixen+ttpk0
ep7gvO3Rx9Xw+Kw0sfZA72096hnacyGET8EgOpxoSAR99ghXxkX6ku5N5Ipb
gEZ4z0v0tkSyTDezTgkxUcoyXwmU37uKkNeAqwd16MvENpFUHprSNIQAQiK+
hIaiQHfGXFJiMe69XIsaCZniW6RxYvrGMPJ/RRKs7qXqzBTR22VHPAL9kiU0
lBBl3+olfY+CHbmhd4aKcAte7/iqQdbsjoYt7IrZYgDBTI0hDjoIpqjGCLUC
HkhJtfINQjwbPcukGh1VVEwxyDeo7yD3eUcLddyRkJrW1eGGheVdMpeofJui
ME2OBtC7kUQPKlL+8T5kDIB0M8Hb1w+smyrNGu0fx01ho6drg1wRTSV41Pgv
7+8+ysmUwrUhhgrHtJFODPfJHPWID8X3/ZhagMqXK786Yf/bL75U6UtMWZeM
RWL4cHpneT/q3ZrSffmb4G4HdgBN//TJ4OhzYcVnNYMiAr9MbPcL29B61K3E
D8/vbdmv9FfPo735WcRD/bSp2bo6wuj1ICwL/DSAMcD1+12BTk5rBBqpFHjb
vuDH1NopuACJnUVAXWOv3NzhEfie2E2YHQE0dUAG19MeVLEwTuJW9ve+t8ha
3aFkGyII20chQaPieladb+EBcY3PqQtk5lJBHd6txozgHSbQK3DnWNct4BaP
BCjXX6XiN41MZxRgwurJ1uJmFMoha437bBucMbNlVsIi1dpYMsfW8bkc7gdV
8yQWoAN2TYL+UnsrMG+WiZ/zSf8vKA/XL1+a+0a8dITkhcP1ePTb52OyPP9Z
iY1FxHEKRuGJyczMYSkz0hXAUvc/V6E2D1se35yrTubJAE2qJMc8knmp0kru
blKKplCkYin/xfBxanitDtvFWoSShD3SybBxq254ezifC8+03llPVicjbMNN
L0X4+pFbxcNLAn+pg3u9Sk4lpr31cXXiCAsRzCbG91dNL1RbFaXDwPzbm72n
6nW53EbLhkCCJUp4QQUOmwrXLz52fjEnNs01I78cFM2cpvX9IExN8Jwr/DnN
IZZWp///BADvyDGZmSCeEYDJWHTkq/NlOBb+LHsmoL0ItYDzuHf9o7NzXqOf
rnWWjISdSK/5b3ndujYkEhUN0EjuB+9kfTRxeG5RpY3nO2I85YKXsIo4a1oJ
gGrdyQm8wlv4l0Php+IwGLxBzGnUjfkphDzB7Ye6yUKIq/PVdWrB1UHAyClW
XFPH9I2Q/w7OSjn/aMzoYfrStdZKckLVD0UF6kCZ0SBSGCAimupRdl4vXMMC
LuRhhTeER5Gp6GvaFGb/oaR7mAhTNeII2T81h/llSY2vAVGypp8yRCE1yakI
Qh6Xz+ZDVVIfAcm/71p+D9LqheOvI5r3UreYa8qBiCK2sMiru853OE57nxnP
p30n10HqumWv8FAoPO1Yqh1qBOeJ8PMsMijsYMP1n2eY5fNtpDbz30ioi+Cs
qH/x4lSHUEeP6SJLxknaM+n05/sEBlvJvqSWfeVITmT/wp8qYf397vOHUmyS
R2/MaR2BLqB1RtZ/L3rBvV3NCn6JgOI0x76uZGAmgXKBVCBXYX7yiQiTF7ej
LqVd+lv9tUE9Bp9kOOXaDsfdzZTnHM2/dDMuWQYlNSPCcUcgK7Y3rseYaHif
7DcmFx5pVXbpVSwOgiUlXIIquxuNUAvnyYNw2G20JoxW8UvNtFVI5517Dxvw
cm4ltVIApfNOiiE1x+99GmyTWrT1hUOmhVXqBZLI/0gSqTuCOJ0ANNlDlUL0
RnXsCBD7ZPWmC9dvdlWjSEzT8rKdI6781itsnGuSK9vqKFqfPMy8NBof2Vwv
oMjnfrgt5gc4ZLACJj4afZ/sXcuwt3KC6GKIlgGSp8qnQp/QE4b2EisX0WLB
Cacy4MR0bwhMKip15NmospDENQJC+o83+RgFDBrolyFUG/XjZzHsAr9Th4m6
wbYKUflfCjaUrMXls7prFapVqE1Yu4pddhu0V8lorjKXY0Ro+D1VlbS+GK7j
rkg1z4VnOrc6VbCBb86W1OFIH6J/UTgPda5jyyJ4IdE5YDqbM37sKjCP/z1e
UEWbGDuR8RYL9T+RPNrSpg0TXjptDHuvI210hQw7ZAPopgrpF0vwQi76xmJi
N2Kx2cXAPrFd4kFGzHPE1VBbdiElGk2cnLsxi4EcY4Nd+MBb5n3STzeOXMz7
P4ni/S6H/3De1X+UWxumMCyb4wFbT51eCibhU7S7RCKYnAH2F8FUVFkcPvLX
838DvL3OBCUk3PURrWbeyZPATCatG6U8rIHB++sliN5poX/m4RBjErZt4pJA
7JJftJGjntt36ML3XYpp2FmML9fuuGqoMzvTMop3SnPRMN4pw/zk+j30YVQp
DcXDcKwL1QkQfYxEEaeCy9hxWmp1+r5drFg2Yme+LxpJcbLZDLCzr/EwBuIo
wPHud00JvFLilatSsh0AAa4gKIV+ozdaCI4k6zQ7obykctGBhzj5Q3BGHpBV
nxkzs5izWJjPNTNBa0xymmZmoZkodq8ryqsKgI64kosNVSTwVFadK91tKowE
yQkxCK2iWFarkDBfI/ZPlEaJimryg93+rXnVpOLqtIIKOlPGaygTnmxrEZrO
MR5hh4HldUYJRIkphabHvyyvM78eIlNcGk5A68gMo4DGzhMI11wbyR1Grtwy
HT6TSZY8Llbn0sE3F3yOyDbds1bPCkfJmoVcyRBgRNyC98dgzLg23YoKWumd
q00LremyKhnWNhdWWHyIVK5RKA11tKg5JD47IjhBTT52YuyCVUdxBbhVl2gh
d9itNqhjT08QhjUnNtjCsDdsJcZuPP83NCuvPyidVnpys/TmUv8+ACWRYg88
E0svX9BkoFVmJ0iaXIw0qjJpfuo8f2W6tw0ydCk16ibMqiYtretv8qGYjVCh
wBHGtZjB5ubXUnirifBjdZouLLja3iKqUqPr2htmnDJyDE/IJZVuMSy1our6
T1mXqMUNWxCzlEzElO7sznpTL6Kg3O2QQzEXBpz/NVz0UsviCiltDYpiHNVt
vgiQDmkzXHAmNIl7xvHV7J9/v6HWrxmHB3CZcnTOUNXeF86A1UUVTUslYysj
4PDBUtbLiILvUW7Lht4rZImUkNGYZUw4L+ihTqjdPFeGvDwG3+4Pg1WsuCNz
H6mGBHT5/esOziUxFaao4SCBnvzeo5+2YD1oUqjXfjOXeo5RIGTPn1gEjylt
NNxMnPbpfuuNQ4pjg89Nk+tm7psw6NsXLvpNGXytpFlD/UbPvAIUOFl+SAHP
dKgxCreEFWL71ZhIV58D8q1anxN2fTlHnQz3PD6AEufRDPVN9ffn2C1wMvwN
10njTdhRLKnHpBNRw1JyJOuj4HpahEsGeN8U8eU4Gn5R61gDsjQcg2DveAwp
OWWIOCeE5XiB2fYzEA1E7U4Y0IilP+JI30s/Z9M5yH9aYyjO58P9OMRVeQZ1
Zahz3RptavYvsb3rtZFvuey6kwyoKdRvCbNj0pTC5mFAwU0AoJvjnXEJL5n7
uaM4+z15ld9ElVigYVuQZg6SZ79qxXMCUwlBuVR66T8e9g9fZIOJ9fD5p4SU
yOFm9fOcc4chKk/Ga9vXCHaCz3KusdpBd3YnOO/9g4nmmYE++MqCpdrbk4Pc
1r0fQyJIC2JxyWDIFgU2zGC5UWQd8giQ+hDIFXA0CVQ17Tot+xDO16W97Ncb
09RIEyFgAZ3AAK/ngB6qDYWFJlyxzp/Q+lvwUF5cephaGgXgHn3yoeA5B1xV
L7RgURSGfvQqN7Pf7LA8Vxop708cZPBkmDkIC6X/+f32lPok7dcLmZ15dX/g
NT4UDJ1W+7TOtQuLc6g9RXwOpbFhSKhTyR5tNH2n/Sp4/TpjXFOaXkFM2yVG
wNKcWDyektLyWCmjVAYqOlXpjaaseCxCT+g6ZaTJ2+q68aBDqkqG4lIZNHlc
6mPTdy1YIESYMiX1HZYXTZUbwQDrlvMqP8jqMKiK3pNvo4cnN2fJo5tfA809
WN5JcYgGvJOqIhvBaRPIX6s2EU0KG2Y7VVeJ8DuNWYqyishtVDhpIF8E7aWa
hfhOOglNBie4WJY1A/6KoemRT/flzLaaewIW43Xao3A43svDg2EpNxnyFD6h
DdhUHsoZzwqg9aPqI0vCLoGLcBP8CsslOZEqSZGs4O0lPXr5Scm+ypBDK95B
8Zo1rJK0XFrzmec5SPoizU4aoc7OU7XsbfrqyoFg5SnzU68SrQsQqTTeuJO8
4jTt9nionMIgTOYo5PR+z1IrzCKGiUqPIq6d0pBQWCygpuULzgJYWw79CgaQ
WRrNbXHkCcVeKxMEoYJn4Nw0Te4EiqhvzAbxZpkK1dNgFGXeGEwSrZoDSNI4
6b45Trwew3umTGoykLgT0n1au+3sLatcbmmPH+xhSHOcf3nNPfnekX2wyQYQ
WvCW7izxf7bB/eAjn+DGVCWT4zDBFawT7V/viewSoqSO0cH7mG8xbIV4wgwY
i72amTIqaZYzsDEwRfwhVWCdSc2lXxPPIYTwornppMQikh/mZB4O7k69KRaV
FdiVLzcVp1oU3sG/9WCCbNxWzaNVzTsn1xNcxtevN6hyyHN0hMZSvQTJU8h0
ws8KE9E71aYS3KNo7PlB/zHN624MT+61DsoATvHTZqd2s/KrdV65pZ38gfv1
oPOzuSudTA2N2waPfRXyFCDlOxfZlLRFSydQQJMd5IL07vI0rjnXWIIvTQOz
8YN6mwxxChrcWxaZz+2XrAUJLas2qtsPYdLubMPI+df9Hlyj2IjJVhq87zev
/K7/vVnM5TtVe13OwBosF0xuOr+LYNh+hDNrzmf/lVo2vxEFu7HBr/Sq08ge
CdU6fAbZ8Rds79jDEHNeNP+L8gQpDtTwi6OD9Pw5arVMJATn4KlIa0d2wsTB
CnXdKJ2CCm3E33fPksCYPcR64xL3L6iJI6RlhYukO+IGz/Dg+ex5NQOQYudv
IF96GCXqR1WTT0yKDjxnNM7HVw3AzYUpMQ4mm8L3YrnH+zOh18TRkUORL9tu
KPMMlZBivN0vB3pWyJ+L/9LV5DCsQLHTU/CbMGRU3fNh6/vTd36aQXBvwaHz
qdmgD/gOuB8H0Kyp8S6eKO7G5Bw8fwT21NovH1JBiavpGBLxkOHdFD1yf13j
q1YzTgIfxMdcZxSFxxDiKRfL/5BESxiNVD1/KLqOjHoVt0yiUrHlzcTmvR+j
0fjXVeD9MUlG2GDHE3M7zTF0xAVPDP4ANpKRUUYrFpuoZUid9XbFP1v7jdam
MjWykwCMFpic6uTeS8e0a6CSIOEvJ4yHnkUJJYxntJDXFktafJNCa50oqvya
mX/al78rWkmJ0PBim7QhwuD9qLIS7jQtg/pa29I0+5jMgN3yBO+y6AyJ+WOe
sSjd9Z10JZiNz1kQ7UP2XOozyMEOIWvLvsz6zIynXdJwPqU/B6pnD/VTla8C
Y4qUSs12boEn9bbbl0+wZABViSrfPKYDN9lZCmxZMRiILis+KVj8VJFc1Kd0
yvXWJnHbqglMVu6C3hmQX5JMLu08QCXqI5SQZKMH0MxNPqK2Qpnms3eRhFNB
q6koU29T5AzT1imyvDKxeKQE6J6u1q+QzKLKmuHaEpLlKrN2/Sy+R75VWXrb
nS8j/g4+YWkGzzXvbqb3Iy7RIgIj3TnFsqFgFcDch26DMu6EJ1s5UowfqTGZ
CY3f7RV36hR3xG87csrZuamw75VOGVu1FJ/Xq7/NDiddQP/oK2gjtQv3cBWv
m5IOc1LANWIpVVvfGqZsv4hD2iljoHwvntIY3GAyhwoTHH0AFAnbuDi0pGiO
xgl6+Meu4vXXMwRFF1pWV2tC5dp9LdPhJ52KTIMsQKPJkTrKxNVY51YrNbcx
oO23TdKsYtEnTfaX3u1o9KrS8UU/btPD1sENRlpnfg6+NWhJ6tQKQ7rqEMHW
4F+W8BeL7eCK3EkXXsAQyT6C4qZrcN/eJ7IgJCFp/ehcrTYY9BLQUAvZ8bVw
0zDJU/TIFb4nSRKbdas2mjkRGTf5JQsU0LAaukxfmTDff2hFFxANlXBe2Slh
86fKIXO15PjVUPcV/Pi47mciFq4RYGyEkpX9KwzZmtjlbiBIw6cWLmGAW9vl
/n4YMHdhG/ViimBgdOzYuVpWXEaj+qH65vABqG49GkxldQs7wv4qo4sUwq83
0h88PRFCKo664uRoO+SsMJWvndawJa6C7f/InxVyggnrPQvpIlyPH5BWXn5r
wlC5eL0dVll5C33tmuVOB1wXo6kwDbhc2ZacCdzzE7luESNJO5CxyOIOTF8n
cTKFZaXIy95jgHAkQTFGw9n9UFwB1a601TBuWZDbZ/OoYvZpfmeAJ+9wGOWa
VJlQjR2gcZrktg+kOdSAomsqfKpgmDt+BRTLpkOxHv37t91tcGZO0ckKS0xi
lUvm1LQdNn+bhuwePLYRqubVHhCK++53fGDzmj1KCvc3B80Y4mIn5JG+uJXU
TQ1vRA//wUSvcTaRrAQstvmEeQRBfp059DqY0xsPPW4sONMhIkrIQAUIaex7
HGHCkdAD+uimwth6ii1XMcovFtACxvujh7pYZiUxd0x972VjbuHKD6mUXAKC
pg07Ch+QvXkpkrxfnyAfwHzWcVb3fIytFFuplZ8BaVe9299kVtevuUVWEmzr
l9Ur831yQG2TenkDeJRfhhPEx1BoU7Vyhwm6XEHG/kNeIQHvniUuUW/nZHID
sG9DwC8M0vfOQpoSgP55xENYaZuYw0W+MnUQetfvdx7ffBUvAbUV/cxzcZr6
NMaHZ72bNKzBt8WffewcpxqTl/qIEGP2rQxxonp5+nq4tz9qUbX03I47gKrm
ObgbQhjZbVe1jHgf3NPc6cdTFYuLebk/G5lnATS9ehrZy7rrPdBJDWqwXPLz
0lSxuyLOtMi6BMwAkqMf8ZOPXlSPiUBLwieFCg/Ha0NVXlATGUvR1c+DzhOd
bOMd2DLKzeZNNxlecPdjfAadqke1/lT6j//MyC5Pq6K0Ykssp4UarPw8gPIa
iQZxjCluhN8bqxts6Clbi1s8beQBIPxNoiz1tth/ZUYIevGCL4X0GT1MNwi6
DJuErCxFHV1c+amdbu3k38GfwHjyV1HVggQ3tZiqULt7ritm+ywvbP348nwk
cq0AvmsVm06GvuSTpKyyeAoBjogcxACncif4P/HktW3lAf/LU2aDf0IOks5d
lifmg5XTRaEpPaUzRqVaOVdRTVoPY/eAMfQpmWTZ6YxbRlqZI0Vk0NY6NeeG
TOBnPCmy/gBvydz5Ib/6MEXVcoqujXxfoVFpbQ7z7puZyHfqPzbTV2IjeOkM
5erSteUf57wEs30OipoV81KPlSjYT3Qp24bYjOTZVgSSTIeeTmsHWP+t5CZT
Ebk2zeIsRl4K+riMIX17rxLAIjY3b+G9v0eejJCJ40s2bN4hSjDESD/CZQRs
VW1nxlOEuLgutK6+iHqFGm1uQSJ+vOJffftLufAFx4nptfPQWY8/iuQZf8aT
Lc34LlnUnf1CJNXPOTslrEgzpDxmGL4urFUSaW7jSp7kM/ZUyrOsIFgtxH/P
rPq0vHgqOjglMJr+tbR+GoDdBWd/JXnVlGuNJ5G8NaNfxoB43ta1OjKRjhqs
6qOwfsKoa1XTjstYXBQYJYG1Gf4MGMVNKJkcMAGhe5aM6k565K4fde2f5Tgt
wkcd5mjUclMKNQVDzcwg7Q3WPuMWS2pywvGDh/fN0X7J2WCMOXgNWPMkjKHi
9XH7lTLkVSBU8c7D2ojwIFuRs3yL+gYbkF9DsXuOUk0z7zUV2dQxvqHNYKXT
2bTJUPA4eyKPGG5KGkdxCAyPKjS0jLMfRxRVA5YtttXBZSvFoMedOiTOiXzb
C7Td9UKLzHo61NGpVnZT16WLlYJcaoHFQBdwWfurtoZabCkhVTv1aSUNsGy8
Gn5s8gu4wfztoDxcxGuH8R9Q04joQ3EnmSaoN9+7ojrkHRzSFPgx1itAEuV3
llrTK4fEdg35McV5rkio0ZAQrQtZM8reMS//a5yILDyl/PrIcLfZbDDhMcy7
fSpZaAWsz/JcsXjIQ0sW66taVP2GS9Bfpqx9NICptoxsi1aBHaOP1evo7E19
tf7Rtk9E8/WezHTV+Gz/HIJQ9YeRRQbfVNa76VmtlyY8Nm2GGwj6mCD01DlU
416MMBgjHFZZOkeJNnLQeAkWWdpis7KnU9q4QmJWNjjNogzxu4w+azL4D4Fe
SdOo4WEUeWMD0Oc1j3Qe37oqqofwzVUFtw4+3cVQK/dJgaqXxR5qZDzSHuar
vYl8qwOZVYgoJ3rE8akVcCLv5n5ywPz8WrzGIM+YcixVgK9jk1Qf3xg+rGjq
L/xDOD50EkovteoN7AdUCsAiKyZOP76OthECOW/k9FzXp3/ixJ7Z+TCskQPi
9jjYL38cW1T0Hn+0YS37Y3Cx2RKDKA7E/tVWExjq+dKvUF8QNpQ5T77qJAtR
2VJuE1XypauVaR0k895ux9Rijt+o6EtG0zCzkR+o8TXI3Ns6vSwJ+a1Wx4Ui
WG5BdMq3DazbTI2RaicsWUdlm6EBqyKIELYXWht7Me89Ib8CfwQdpNG1iMh+
wgDAsMRd9J8JSnxQcQuzZjovSDGvsNkVHZmZOZVHdLpXxJEKULl9DIwLtnFZ
WXJW08zcGQq4cc6eiTE2fKKl+jyc7w7QQVEtYkexWfrB9Rjrmw0mxUBNy90b
zH0Fj2GWEP7CDWxEXVbc1SkXU3Dli4E4t0CgsbZFcaBR2Pb5suNZqh3R/sjB
85ipRTj3ZoJXp/TWG7+PMy0S2KwlDvcqGYE4O84uzMwwuOpG/3SlCvnVTivx
7LD3KsuXiAgcocTP9n8V0e7b+KrsTcBkYwD+zXa5qZRuVS92W+I7WV/Qpbjk
hwN9otjhf7DPMynmTi1PeRLarPQq3qZiAW0jdkvO55oeFkgxRlXwx9GoPFEm
LDLZjeBuf/Mvf+LjX0mUM2PTO/7DOB52AxXaiNZbYL4zukjs2uoVKGhSe0KX
oqerFxGfwCGlsUxchl5k3QTlXTrC7/IHCFWB/B6NoWNZCl9lBMYla9lJmEwN
4PnP4thiuVttdUGIwZhLkFbMNqIsqSlMwy9O6hqsmLrUwUy9hev7Keh4s/3l
ImRXQdz24jOQSu5YmIWlTuukLffK5XebnQNiYYa6BBgmctGnzpCtvnXulr2N
n2oUpmylMd76HWh/wXK6jfxXl7pvTNwhfjq0gpHKAYz2Lo+WwxW6m4qQu/vq
jkuuqgwUzAaqyT2yvh52P+hInTr9qorZi5dx3wtOaiuQHdfE2+Xw5qMuC51e
bOOkplFuZenolK0cZIHED3wg/H7b76Q8Q1vW7kR7VtPB4S6V90yQREZm0YmA
gEZp6FpUacuq8yO9GwCdPZJVtcqZpTr7ZTgNalVFlvJLH6dVzfBBqBLvXtHw
r3RNrjYJ3ZrMRxH/G2Wbda+NUlDEi+aU2BApyoTD9GBOIBJY/XdIuea1rKpM
vgulSR/LzSxRk+xJ/7SA3Xm8pElffE2xZLRJCZ9+fh8u7AwBtkUvADKAvRTd
uxqhi6df1H22z/492of1wXP3XSim2teSsbpId32O3ASl3zmsDRQk/7f5zSJp
971agaNquerGNrrFnHuU4tlxDKTbadVDSSCGYdTxZIwFO+EP/+DWnN2ELJkx
LqWNnou932a0sKrgjGTm5hKsOisBIM2s5VYzyC6GFARMDoDWiWyT8DUa8Pkn
2rVfDjtaYB+lpgdFkhYXki7p+X56QSUleogKLgyCAb2vN2myf1VTpc81MWyK
driXwNGR5m15W9Tw02tcYGKpZKhlvBDsiFnI/jDPY9Cr5BP6f/SEUXrlbL/u
Cpw2xFp221x4IKpMkoMc3xvMCMOIBhQ+5uO8BxyoIHvvP5aiv8Yaf1UafszM
UUHIfM/+qsxIF+DLWI7PyhaLqRCiqpmoahgDX0evgwx/jpf6SJgQAQYOUtRy
qXqQGmShEKyVO0fA5/HDnwsCqTprsdwR6ovH09C7dfVZUyUZxAmjx1DmwWY/
6N4kbnOpNUCjbaFp3XDB/U+04HBNsd1gv1u4OSQurBAYFkn/qrc51HyLozsJ
lMSOBdus3pcNJPNhepuyiSOz8TjpBaEPN0B+VrCG6Lf5sOomS5h1zHLoKfDt
P5o+Ot/C5BN1LojNezS7OgBeqrZc8EEpmPn6duqa5qE+QK1MOIaOUvVhKH74
BagEYnlz6GPvBbg8zQaP74iv6sclcwmjOdBTm71jxUnfoBBE1lv24HlisHoj
3VBihTAxkbx/dAaD3HNhRycE+HzXX4XEfazn7zB80VBhggYL19x9H9PptjNr
ljLZBKqbcqmQix8xKnuDLslI0CIOtoGjemx+UrMKBWdkVwhgk4oCHu6d8yTz
pvcyD0MhPDk8iYenQzfDcU53e0XQQuQE7Z/S+zx2LOkxAih6eczV3lBHUR1w
OnRuqjw+GXQrCAxHaprNmW1x9TWB2J9jTHQwflurrK4jCqOU0mZBQSxl3Ix5
6esjVlwRI1qy01WvNEh8HGszcapbFHknAzc8yue60+MxEqtUQwvlXlNds+4g
b/6f+httUwYrwrk6bmEf5fpwR2VGXMm5ODk7LajEsHPKQAvv8mirVaAssjpK
7bjfYApr77dOAKv0faY+akLg8IJNOPZcPEvygIx06Hy2F/QogVHfD7MGwcMU
pHxBimusvXHPijRmb7zTx98Mr3lZgo0WzfVrtUJqGBewCLvvKPLYaQrjGnFI
MjZ+yTkQa6km8771xLUFaCuW7o1pjnzxse9ZLiM7xiUiNovpj6gmWxlLPEJD
M1n0Q9l7Eo4dELpDXeXt0ki2oD23A5KjfVHBuGohYvHaMGtNS/oSNPwTdaR6
FuJuTVOrXBx2k8nEnL5X9lmo1Ae6C5CFJbhpKwIPOzHrDCKOioytUJBR6RfG
vqaFdM3K3AHCcVFowjNoZMWj57CbwfF2b0OstKd1XEObdPOkyKGvjReXheRQ
Hbg4FhzS31TpYzb/gBAG64MP8bRbiC+F4h9ihWlLhcsy7/rMF9weNoX0IdHb
T48IUehzmd5iWASXqQL6T7A0VmzDUMspedJr+9K9o6RKFW0D/qlzvD7XuOjL
5DeIZKZLn86NgLWwAQXCIbF7sr3B4msehitoOoNlAI/ZbNatdhT/QMoYYL27
Zflgz1eMbcUz1ISyM+s0lRLbPbYXZTbOCINcZaHBpgDxexlOakEcrbi7IlOi
FsJbHmOttguqKMtTOHh2BwbE5uWzeJODrh2meODLSxSeMH0D4EEpujQH1G0r
IDUdL28OL+6u5H2mzWF4CTnzdCJl23BkM0bu4tqd3aOdot3Y6yGGTgdso9G3
eVtgnt91m678I56/rlY+C3OwcprZOqiEEfzvJCnnOk7uRl7tISrjTF8WTQxX
/9rTDASq2XSLhjh5pboCg2DRnV0k4m1G4UBFob9I9GJFE8TVvHa9IL8jFmmV
+6+bBpFsK5R85pmcKCriZR7NURw+u+iKlvKgMLnFDPchv0hF/xQi2MnwIsoL
KZsjTgUdAlQKqKo18+hek/8M11Z5M4CvxU8VnFKcNzMMaXv2NLtvPcnkg0R2
xNM0Db568RgbQ+pF4VYNDyQtFtcI9JQabemKjm4n12QbdSgGD7ZUgvP+fEnF
QQxYDz0/qHAUrIO7tIu0tadw4RfWby6LhGtDRjuGE1gBIgCMjohogg9A/faU
0SUMbUEI9oIT+nfVYKya3O+mQ4LwskYjAXvXfVtvxYkdXSBS4cWjIz7Msl0U
6UIVjxJJe+8MecvwkRNkkzfEWy/K/XFufMEdfq0STz9eksNxAGda5M2ug9he
H67HBNsX8i0WW8f9obeDDUxA4Uxl05+VXgWAw2E8EQ+0giJxLjPkIVTDdggU
Bif0RPZu+v9HqvPjNINKTps3NkSK7My8EwIhfe3n9x0S1LsswLC7XbC4Pf65
GNQTooIyAD61sZBnj3/zdH21SPw4noikxrNfhyfYVoie8jdchcWWwRj5eOc8
u7q1fpYB1piSHsx/TJ44hO7MKUsSzHx30Di+90LGmVAIuyxbzmMYxJrkWPXB
KLJSi21TP9gM/CGQDzluy56NhyDZ/E/h9d9emzD4I2QhxJjpGOIhQfn0uZ63
FvIpNKueScRpNqlDpGTYhsQ+9pb1a6ald2qBKk8CED4AMwhujuD1CcsqO4Du
2FuDc42TV5CH/JdiSX4HAGNZWTD4EiCkHnFJVo/TdElBXWAFqSuAJwCzQ0op
FDYa0p1A3oBUs4cMbEjUWNLY7+5E6GSL7b2a+vX+mz3W69Hd+Zy6YWCWINP+
t2hiRm99gkBXQKwTQb21rKl95OWaul8DqOKSCYPShUkYpYlc+G/z8kDKJQzi
uyXez0p2Bxwzi68EXsrRUgsVaoCznMDLmcxgGEki6ig304H+nom1Tp/bllyG
UvdB+dZ5VzNZU+QSwc4HF3n8gu1N39mUgMatiK77QL4+79eORFq8WuPecQuq
rk4r1t0FzVnv67TJoort69GWjsgdWLz10q1RbldnMMdz6wSOn4aeWa9o408g
1ZYOg+G7D2IgYezGr3AFesRqo9rr9Tp5qSBVTM3m+BEJuUQJpNPUixYRQOBy
Y411ULWn5rfr0xo6DoQMWZPWqRJmv5wuM4s9Ghoos9K0Pz//7MKLhl3GQw32
xtLEjR5QQkmzz7x50LXN3MZrBdAPVCV+3EQq3+Ltt0gjI3DcP5UB0A3+NV59
wm+1HZRpF89ce0qRJ6yNo9IZZ+mPx/F883MRMlIj7v0d1clsrm1a8LySgrEh
dOuhipqFxCBo4n1X4WgZwh5mx7ws6XYEMQgOrRCYPT8VBYm+b4/0edFfClW8
anjGYTs/YHP2DQ6hkQ4AgBT0hPNWS/SPPb19HinrlhRp41G3qx99BX1Y7V+Z
g93hs6XL/EnHL8NcjjfGsc2YJ/H1gRzDddUcbJKpfZ3Ml20UbfMlkkLJ1d9U
2p3kDoXkWdRHxIhMwQ+f7cvRpaJrYVKtskt3btOhO5JuyRACqOz5UrfSNOmt
prs0/NnauhB9f7kH4Etg7YD+I8Wjhheu6yzFCtCitJbopyMUR1OeuinFVdbN
T3+T5gLqpfBd/V7dN6ZrnFGIEab+yE9/Y34uP0kXmnKhjCotgqyb+q4YiZAn
JQa55QsclZ6oyFL1qhpkriJuYILKMvHqwD+aNMmM/10kFLr3UHwnIk4nwJsu
xHmtmK8jgUoj57AmV0TJA1u/+vsDCdiPbP73hHdW1dl/D3BVha1Becpe6OW/
BnWt0phH1t1E60P1DtTzg7TkCcmqvgM4MhWukHkcHy/bNPNi0qU1lDQxyVfa
KQdIa6d58xISykJjrp/NJMcRhNbSSin+xSbKUHUvAryn4hsTHo6M8YQaM4Js
Fw2to5GnZz4QKJWs93FzpH180SOiD775ew11nE7L9At9JsfbF9lhi0N3SIao
MvxvuXkAh6sivNRIqHVOy+D8GFDxiSKdI2/mR0uc2fIw4nhfzd1UjbebfmEh
8//RnUv9mD7ww8Osu02TJD6Wu73SqhwYSa8yXZ1+Bym+dlNc9iP0nHx2g/FX
ufmULZOen7eJGDjvu5y1ZF8sSYCF1lqyzl9MYJ9A6xhX5/4Pi4oBLCr1+kvs
UqhY8pvGuGBc979JdqAvz1wrGJJqVVKzR4lOvDDwA5VCeL/JMeN5kkJSFbKJ
/o8XEFKCcI7vDnQZrrot7XG2KmI2XkR+y5mfDusKnoqoMWN69+6ww+n0X246
55edb2Sbpa5POS+OIxQy9TBqg7mSHcj9CNhaP7MjvAkY/9CcO4VIte8IlBCD
GNIs47NDh7SprqorC3skXB17jqhQ9gbIt7YZqXudqZW6H63YDSUespRCeV19
P1vxvG2q0Y8/Cgj1eOOH0vOWWq1PrxS3IXrcjepYk5nJ9h7G4yaPvlygPvOX
Hh8BSxBkjW+x4c5M4KBNZg2R+PR75B5L6sp8+1M0K428edHYw0bQoLap/M9X
6GVL2m6+MlrQv8k+b21XCrNsrHbMk3G/at8DZp11RC1UDKMrIy0SJxeO6jef
j/Hnq73710taxzYDiEAgIXQ+pP/h4EgGtkug+jCRUK+CXPUAynewVxWpEcZD
bOoLRfMdVzBx8eaaSkTvD2XemHRXOc0PkpFmxk2asQEIUmDiJSZNLa6HCbh/
xoOHUTyWXVmgDZYnvrFUzJcutzsEpOEM4OrDm6kl9p1KJDiBgjowne+c3x19
bcJFI34A4oB1ul19CuCf9YHe1AtuHAyGxiyXORqU9tu095LBs5v0YuE5o+0T
++w1JEz4VZAOg5CPfOxzAZExulVdl2WnsgHMdbKwte5Itk9nJvuAeOSc7XM8
hpHzWQUqUGhBRWoPS5HftaTyXJfjZH8rzjrilU7vpzxRIrhKCeZgv1Zq31O8
onKDpstE42UJaADXfanyLgfBAxeQ2zhhF9sQBmD/BkSsbIR+Xi9qm1dsLdCK
2qopZpLyjBCn2tpkOSa5W2+MWbtV9ouxK+M9EIlTcPnLwWwiVTMrETIU/PHD
CXPe7MhSsdeC6Kcv3MbFfaK1NbgypboIgZ+cikyTC+Ii+7E47YVvhHY3wBUR
T2gReuZxWvI9CKaBBJkPomqjKdr+hCSRtbiHRnjTfpDLh0PNlEzF4jLDWMJe
I9trphFSE0Ic/Nh14gtTe0G4tf+POKasOL8F553enQ1ZVyqvurefWseT/DnR
X5GodsLHEuSeOZNX6YrMvRjcnOFtxW7hxjKrUcrn/NOVhi3zOGU9RlW1cULR
Px0R67nKKtdDRgPcbIaenMDzi/5mON5rmlQr2WfH4NzBkAEvnpfulPJeQOg2
Bh/cr2p/7mZeaz+03Zjop8WRk/UeNJKWs7Kha+b0fmJlgLhn6801MEGbY7nJ
jBXea74M1T57WEOnipforWY+IXw9ys8pzRokqTVmI/CLbeIGwRngqSwxgcQW
572VrCgeANQEzqjikvBTbDyhla8Du8hd1bCSmbIEP36NpxwkMmu8n1dwkEXD
ITWP3SBZhayBtltxs8/CxKwiGMpOxWu1VP2Nkzy/5hRt10cf4f+avWUPwfaS
mYkFZxxOLKEJclSx1gzEwkYvhddcJQlroD/ohGcUO8QTgkQYIbvp3wkqsqKg
IXCG300PPM+LDSftcyoUJ2HgnJz55c13d1QHTe8EntjK/vtUBu6xMA8gkQWM
W5j1A+yfwj29G0F2YC3Eb7NvflicSUqrq13bBSYlkRWjXqn8f7aQ6GYzKkjm
5NWj3EEHcLPUIEbNvdtYyJgzUBCRkVrCUBYJ9/QL3poiaf9zb1sWpnTu+A+P
yM0HlqSYxjn499BiCX9DQBJAjqNYolbL0wjrdLhIzgR7QBsCGYvwXjwvwLAe
ThTUmHgKHLGOl1KVub2NWWOQczmTgHPs6WXI95/Lfp47Q48Z/M6H0flTEgIS
lXqQYvibqj1EZX17jrJv75d0FmETuq6kKiX2MhsNnejUUKXSf7OBe8pClFOU
w4G6Z9ZEev1mC9L2Kv9sZzBJbySrthbuNXVyXDGGT8Mw7y+hdZbTA0fjKS6C
zTlp+sXh/rRZVBd9pAv9Oe9gVLman8tQITXf3C1sN6WkjNfJKWMCKI2Fj1a6
TCTAwIKpUMtRY4Re4Ru9x7NWne2VLFJhgEJSGwpBHpFzRG0iacxI9EKx1+MK
ZTSzzAsWH4SDWYAazk8hK/TpSCwT9fJPNErlTQXQWvCZtdART1eObu9HDcZu
NoGEAIJKS4y/zgwSIeXAVv5Z2dus5t+0+Gnq/O8dCIBGRn2TFPS2m6jU6+sC
AfYiIzvTYxQol8HN8zg8J7HTt4/1BQ0zNcYxuxS2MwjndQMajMcfO2bpQYaz
3CeRQYKTDxET+JtaXnlbLv4nGZ6sZTV0vI9nRI59coVM6PYWpPoKACJUknaX
H+9Nx4fJUzisP7Y/NJ83KK5LNJOF602xLNp/EH7iwrwh3iuD3WtnbjLIERot
JGTWIDuQKm/vUEzgX5bQAMFXWYOm+wYQdHfh5S23X8JBgz1VqmvfEnM03Epb
2rxqk87MDgcJSxgiVyTr0HA6XaSOXyJ+bLQAid+77hjl3FZLsmW/Qy+BAlht
hmi/3+1t1QQR3B+wEbCH9GvyGlyRPTEUQd3bDy+95UOUkvZs1B1CcTeV16xT
sff0iPKRv8VhAsy6GmXbnJLOWuwlQ7onO5lGXARuAk+Wl9IRTo7kbifO6ls9
I9Ly7wIdWG2ppW6LcAtrjKYsW6Z5n6JnFcmH4vGjD1ZXx8pnuOmnjAvfSpWH
uNj2ShRERrmI1sZU4Jrlk9rl525xCMYvJ7H6MyYS2EkSKNJ00IyXblNXsVlF
Ck171OgB6dwlhS1IFDrotS+d+OAbcNfhfOwnHAF2eDeDRyd5P93JN8cPGhV1
G9GeqvHXggrS9FNrlvibpn9r9W35cW1st9ibdX6Do1J7kWakyNUrduNMbloq
CbbaVeZKuQc6MWLgeIUsm+b0JLZ+VgizAs6oYOLtuLVYfWScH6kiXkinzDiT
E35Jvv5ZHSKRIOhd+o1kdF+9bXyyjUUTQ1MgiB0CCMKo/J/21F/sVB46ffSI
oKGSAXUHSPNFxP/+uHeuP8zz73qwO3jlOoRHDlEG7O/7m6ZWBkyZMHLVZs0+
veF1PgqNmQ9oyKWw92CRtvsxgDAA4eM+2hdd/6kzRQZo5qcbPtaJTNjx64r0
xPo+xc5zG2UM/wwWwPCzeQlANbIyDGsqD3zUOOtvKPot0rQ4PwJvnuXLeemw
uER2RKbZAOcyDL5HWmmdOcSYkXFIt4p4njNMDRQyba/Aey3fOj0H892KD3sI
42Cr95M9AL9/d8LYJWcEDpCo5TK/rWXPni+jjsnzj/OpwzdrU9oScS9T7B7w
1WekGMQ4bBmdJ4f/Q+RjHe0sudlNZ8dXlMXU9DIiOL3/aIOkRd6YjcGBeG0h
vIGSie0FG2FLqoRSRUilIZJDxsGC1nVHy1AtKYKRHhHGEYnNClL+zgSEhISv
iqDGwANC6RIld8titas8g/twXy2gwgHfSZ/LHpMC6uSGgcN+/z6bFadN+xuz
czQyUU9fMUpjeP4U54+TXNLp6is7fcfFyT3q0I3UluDzGKWIW2wio8vYSMxq
Zbt1pYnLYpDA3tF6ti3WHh75nOc+StyJymL1nef3P06Ik6vhWX0ZN+1KcyoB
kf0g0r5TX8EnTmGW6l+U2MwUcVFi5W1Y91qs0Zf9UbhfVFjvRRb7WVkGA6+Y
3s2JNJ48C1AJwKRE/7/YkQzZGsobJnC01q2w46LBrC4VrmmuQT/GbKo7Sthb
kvovco6lgH985lYmQkMKn1ht25MX+v66kUIjpKCv6O+Bb5uXKi4C9oX8t4C5
yQj31qJEnK0zj82xbCEpcsBJelKLe6UYzyG+vMU/iod005BiUR+67UP7ylPD
z6N1Kks8WLEN/FBvvERWGsPdkBfzLHo2oXuxM8FG4D7q3jAfEsfjjfsuwJGY
uMS5qPuLaWFt2qylEO+TfikxpjvlgGtQgyCbCAc0SL6VwSHicCdy4gcqXm5r
/Xrwj5i+KQxJmnRV8Qn8y8xmBnyIMMax0EE3Y0tXPdOea2PUXzjIZcUhH9+7
XYRt9SZuFFqMVDwOmEDSyos/Rce8Zrt2tSgIL6f2e/j5NWnk8IEZSDiITyGN
vkz3SB+lGWqZTsFYxyLf1owI9e41Md93R8uB6NzZ0C2kNoROkmw1RGl5ju8e
6tmCx9oJ9y5/W17SFMXNEbLwji0WKh1/pOfTp+82Dx5FA16Jhq2HBchNrXKj
0mWuE5jCJZsWRGO9W2Ss3Ih31x9UsULM5wrbjsl/Qp/JC4P+Ey433FGbDMT7
jhgi/3LolLp/wmMDFa0cEWaYm9O2/0lzine7bfG5vO0CuEIV82Do2XRik7Gv
RWxJ5IizyypvmiqIUjSa+r3l3/r/jGncnANMES9rkXws5uxAQ49sVb/3Kqny
b7vyYn3lHGN2S+K8owrgDb1MucBGZqA1buaXjdZrDSnQlEKA189NR5yY9SO3
48CWbFdpA2khTTS0bIUtsrgeyZpjPKxgOb2Mxg1UDMYpxzuE2cGpCp0iVs2u
4EGOq1L+jK4t28Bl6bkWT5jbT/aUqx7HTbc0xYJmszLsYWUFIj7bLzr3iiid
LdhlWnV8VgiAVGofWFWVQIuR6HQZ/YVowXloq9mzstKrIk+LY+Pyu3ZFcR9t
jmf9RaPTObnBUjunUd5t0Qi2RRRWn266KX/vmO3yEZAvmAWRGEyOYu1s8vkj
hPXo4tF8CefwftGcsNCbPu6yDx1SCAxoGrfIyUx/S7iFZS3dogcKu3pgw6eC
PkI9deG6tqoRYQdsEXUhjdNc4z1Pe4TMDVPpddta4xf2PJ/5jFlPjlmyqYts
C9jDRo3tIyb4ms5RPDtVfbISVyF3DM0ZriLP91olHaH5kA7DBfcdwFJ/XKdR
7UjQV3+39y69PfRoQWD9v3f/tD8UwO9tEYFNSPWNqJJAgp4xGGjE8kblqfmq
etOM6Nc00NHx1gJRNBIjfByaimjMn7aApIBpy87/GvjOe95ciUhBORR1hsDX
JuzBIy573y6LfHrstMjWy/nc/GyrMYNhI17RqMULPcgmK8tT2VA5JmtlnoWs
kWcmYjRpVLOnY8GWPryMQNWXGX+qUIhdvHNkiozBTnjLbpyZb6Zd70wIxUol
imS7GOix0vq+F23e0nEQKATq6edbXYHqFOFXyXYzdJdXmd5xdme0ZUC8qZVd
xFMLyE7lmGQEcqV5SDu0gmLJeI99B+bZN+bU62aPimPbtOsJCmPDjTmVCQCZ
KCB9W75Ltdgf/nKBguUjU1+j0rdndbE2o3xhopy0c24A0+Tzt6PuVLp2yIUb
KwIBS7jrA65A1RzJMeF6NRr9ntHSP5qtooD24k+3eZ49Ec5paRsIA0z4M69y
fYEeYpjH7BEIBuX2A5OnDXAZ3f8L/h85kiz5ZC8TQeXx+E7J3LnXpVpAskTJ
ardlas62A0UkWTFsJKKo5sEROyOjms9xKTo41r80SZZMp1DGLPqGhUrWn4ZZ
0FGJ4CwJSlh+aD7X0U93Uiw0KrggxdR6HKLE0aElMwvr8JAojcQHPzTC7ZEe
8aRA+/HyyhUhjpSfa1MVW2eMvCFB77eXUB2oHbkU1VVqIPvW+ntXZ8BNbpkp
pS0RLAOPWOpzhX0i2jB7AoEPuwM/Sx/aze1+Z4lru321lGnvLG6FIyaapomI
UaiXjlF+4W7g/tinnO8iY5HAjNiyRKpBNvjgyxW6VtdxQe//S5k0kdpjQCPd
dBGlHW9ld9hUQTM4ipVV4MkAHphDrrwLjvDc0US/GSqhFVuhmQrJiRqVWr6P
F9nXenlWCZt6rVgfqdgAgb+m5MIY6WFQcuLL9cVn0/F7ZygobCC2UGg76bZc
aNEo0XqDP0Mr4bk9XkM36HVL2D+Z5k3UqHseo03J5w7BmenjdAyTS9v/RzWI
e34dvIPs2LZKnETnPKntsS+Hteag+NMlq2hYQyqB8gbTTeHmol6+LR/Ee6jC
h8JZXBSZpHFeZK7NBvzeNFKMDm7kVD2Ki+99Pl/8xos+d7PlUOKGkUM1It8C
DfF09iu1ptgm3aCdkkzUdinEteQBbjMEQXm5HTx62TUxfceJsFGG73r4QmqD
aW+NQiBuvVODE+l8IGFA0NJmNo0i6jTln+zbgr7q1iiy2KrgQOJryAO6yxBM
H1Qm1Td+6gEFJ5M30XMXaVQOXYwmwJpJoOU8m2F0k7NnDsSNtB6CcmD+bSeR
8Ke6e6KDdk4p/J0DS/MUpJpBm1ydGeO+JcBNgiyu6hvBbLDlCRi0LKvsVnos
wGfBfmsngN0TftYC7rDArPG1+XM6GKXAbFi8g/mBDAvpbYCmhOc8Q4/NOhLb
DSAkvsBWDz99aCcvaEn9FiSYzOyY4pffMgpahhgXqTxSH4iTTukInUcrgPl9
lLMLrE3tXI6EouJpal3VDzvRfKu2Nh32w51jekbEokCqbbPmk5zF2o5x5K6o
b4JDNTe6vEJC+ODhyiFIGPG9i+8z/RR646ke4pecaqEp+cXB2XgEh1r/p6XL
CZ5G2lwgAOG4KE2d2ooA7nFF1ogV8D5qsIeg9LOsKa+fcljV+kyuE2yQyw0h
T2RM44YOENksd4dvsCP5VNzNxRjvdwmQDRIH6V7tDsYKTptyFJJbs8SLz6Ny
8I6zpJwMTvh/QXeeDO40i178hPaop2Bb1lQZnhzXT45geQAtMo+nwKRzPr5Y
WjLDH4W3lwFlzCQBxwMiiRnKT62hrgVEDj5NKicY2Jumc7L18J3y7P4iNy90
0Br5J5NAHQR5JjesWLAe5r6tV2C2ELXPNrAGhjolgj7EDM/L30cDfAg7+qiS
0BRpas6GqvqEB17VlBPq/B/Qd7MZY3hn6YbomH6i1TNezpMfl2skZL1jvZmC
NdWv+8YxIJcAM2gB9h+mCgLjVj1WQWgluMdjci/RGGXIOLZTbfN+GA0VZPpA
4PLfcvyib34SbEbAsPgXP9r/bxM/DNlP5FKsh89BEaWl+q7w8/DvXlIqtkBK
ECa1snrTz3/RZqo0JcrxA5K6i6R1BVlHChmCYvnEFh1uh2j56BeO92hy6gGS
iRd/GQSTKA7MLaGZhTNiPzEg0Oi7c2yKWDtqLTO8dcfYrgZFTMpaGlKsKca0
gWQZjOVsyO3sHoMlO0HzsUukIGJp2dY8KN99mhLzFn7ZGyRNTb4BmLxcRWgB
WubUYVLwlbq7Fsx9s/qSjP4RRIY/e3z7Mz9SYkFj68P69DHiz190aKylRWSg
xzBPIQpbKtuMj6dbK3hjvYNcs/hZUnEUChOcO1/zofJU8flsGQcdQCpOtHFk
e1Ebakx4ZUjHichLbT50JbxMM9Yn6IosisXJAPku4M5Xcj1KVfCdrxei+nnw
1Ec1IR8Zt+NZh6DGDohQy8AfhxOqMB8hzUK1mksCPtcczTjq5YrOFjszpncc
/UjnMmsc61xuRCK50ZVoz8eGmA9miWOHM/ezIBHhItldGWUWWt27M6pykoRW
ViNwKQDOPgBBtIQoXYWNSuNLf7G8JR8JcjVynSlUw4CZd8yTZf26Y8+ztJKq
8m/ilnYe1IYFdG3fCvCz840GDxd3dyx959weLTsaOdEmN9mFEm4r0Q54dC9y
NBS2GSq4xcaOZHBR7Vmk1GgVspQuYkBgtLY3E5wSDQiGwBKLELzP624BDVIB
6pPzPUsfVyviPr2XbHRFvdyyHhOkabmrIgaPPtJWj9UC7Gf7vSLNmi3U5536
ISepzzSXiv/OrLBINQgUXcgDBz96K8TOe1aeKnEmUfNK39aZQuL9+JI7/3Sq
sQR6R4GUXsuvxGJLw7LJic9mRBKU5TJTiiD7wWMji7YVp86rHTxRpGLKvJOT
ZfcTdHG8+Jo6+ivzDZb9spMLfcgEZ9VJ6jHSZreHQJ0bn1sYIEXqRKvKP0hn
8JorTmaZtdf8X6qA6w6C+jsh+UD22cpd/29YIrYsyKMePJjZuZIiA6s0As2H
naJ9Qxoz5+4qTNSqqUOSZs9/jGdd/qwio1GfOU3xvjfTsYIiGMSEQ2P0ecZS
dPdZa+gtjNaVLal+vgfyqGI0SOgGK17aUeKr4qW5F9CLX1keCtTNA9SzEaMv
Ma1advV5SRYAVhZFgH8b4CNP28h7lFH4byTQxFbpoU1uysQs8SUuhleafey9
48+ji3paQrFeREOsfwKbrjLylPqLeX5i1c7dG5qlzVU7qdG6ZG4Z/aY5fmqh
MhnD4yNEiiLgjKCogt2ucTz+pUMyhq0HXCSaHq2RC7o62dG3WXFqjp+AqIrs
42HG3LSf8YdTHSvKuYp2Ta0N6sx1C7J4bHBQhs0C4BIUZ/wjTIU7hxMrkp+0
Zfp+lZ5HaUf/vTgtvyAZFv9dRrDyrtO1YpYNgjefc7iHAkLO1WNqym3zRRM0
yDLf+qG1CqaeivMsg9nrUDts+TMd7z+YOE40T9vQalAIlA49M6wfBsdR+7Bl
kXSNKDLkvA2uFyIQwA1aSyz5a2gtTvqMRuktCWoTd3dUNomBfPYzonCXNgAk
gjK6/daRRsPYqubK124SEaVGAsNFKvretSg6k03mfs9bV61MBirOJuAK/RFO
cxmw0ahdcfUFxU6M5SeZbjVs0BOjdVESQcw/OpUXSP4Kxmhho3a/yw7onGr2
UGF1/Vtpx/KEI5dcHk8vzDkjNV+l7L+VRSu08sFvusGimA/1TPWKrVUpDMIH
wXZTJoxdqLVPfEFU4MY51LKUqeLnsEyrlXjIEQG7oBatvx14Gg8ka7yewxKH
gsjjy/0mRcx3aLPaKgBDfsOj3duI/In2QTPN9fhiwNZECLOBHnH0UmVba3xZ
l0UpClO4xrkVDdXDHed6xQcx+RPVOReh97tUk6MPUjWLyyBYQZY/IjWDqELy
KkRGHx/l32CqXuhc7f6T6StZynZmJiIq3pk4zvQUuBif0RKfOb6j46wsocx7
gYsjapbqtOJysMvIK7VIRHvUTnUiBQPyLXog0LIMg6OkX4UIUG82LzsJnzF2
swogzm6Jjzzw/1VcYPuxcfPJ6AhX/9OsWMGnWZCE5fl8GlxzEE6JxUpWQQnS
oTB8rdaxIemAe/I7NYfMCDNGTr4jhxTLIJuYJw57J/OsX2q4OjWbbe75jh3U
A/Drf/BpvMMpF6r1d45sw/5N73modL4c0mSN1TJDBKOCKZqH4yYPTfpA1GM5
VdSWvBTNxraNyokY3kZNYu5wD6FZXS4k9zi680om4th5LxdptRzfio3f6BGs
o2ORwP5dL4RnuNOzSkX5mL7ardMCTGEZAQZAL6/OSfoEm0zNpQYoi7bvLFCH
JPayOdP2nzditwzoa/epGT2CFOzLr/R1033S8xN6siCkfgwZuwHVZna20Z/W
XESYPwAEiSLhG7MRn91ghWgleh1iuuRNEm8nOweXg1xVgl6WseAX8CFmAD3D
58FeN3wFxPE9X7ETIDmJWdRSHZ3A9kbezgUZ3MaqrtEYrmnBgcpjySg4WbYD
iuyrRb9KVkDwhvVihD1fAicPEc2EClIlAIL2KAHEhdavPJ89rmjW94btGQSX
a0AIT/BOqGFtbM2sTQ089+Zlqly+0LHmwEBHiV7Iy0Ou+yss2doYoE6YkEu1
AKN8dRBIG0DSsbXx1BAkRYdeBSbyojVM7TrtEF5NBL86o+12L5h7XcPUtm7j
OOd9ldaLbKdIFQ46Ok7gXbOFwmsB0x1A3W7WGPP+VPLllBobD55+itt84YIB
QjktXA/Nfbw4I1fh/opLpaVXW01zSVkL2z0idEriBLdtOiyYSG8xdHswwFDS
ENUwwhxfpu9wwEIzFSz6sAi6WpI5qKjzQraGckNeh0LFBdBGDMgtGfrL8DKC
LhHJ3B9HnwnKUyG04brATGkbOYN+21/pqSxEE9nLCh5Xw9YaJLJDnciGN1AG
u3Z7oQDTaOrk3P0IPYorJQ/VnYjqbT/T6/DnvLywwCD2gAjC7pZS/UtTYu/C
i9domzmnQaymbID1NVlT42mrFdbdfVUiks7eOqXyIrdBAbBObHIyG09Yr/0X
fdRwfahV0OlMUE3Q9Sc0m649celCCkFMMFzqp2ZwiOhj5rvgtvXINQ9ENKpC
3YAwQrbkpEWVYnVnxB/CLB8WfkRx2P1AeJsRw3xwqT6/MOk7aJFcRJkyccuL
QUW25K2v66MP1IINxZt3KzMXa99Iz9EalskYDcQDpF1hQF7xMuZ1dumUHrho
ChDi1nHMIGcXDXIriflcN3MMkBBS/PixoDskUcE7aafIOIL9LP4r+mBFB47E
VJzjKFn9F8OgLAb3Ch4D3feWHm/8SY8M+uVG4wjHUoE/HNomOSxAJOxPrJo+
Qyoey2Z8+mQQbL1MjQZZ9fNIQTgg7wjKratx/QmUMVEl6EKqi1JsQXSl62ij
EIymRN3dBvl9o3EFEOrs6vB6gHFwNk3ZcSq9WpP1BIjBZYoa2r+ax+G+Hk9Z
YyhTokQknb4YIn4pBP/lm4WRpwjNnVP3remKeTjSoa5uNGlRTZTZz8YUrs9O
Avzmjf84G0iuUXKirif5EqXZ8UXfqPKwLuB23uT+wBzaKNTQb3DE4uNxnCXo
ohZNTH/a2NyJLJMybSIl87gxOJpO9mV4Ltf57n+oniPUi5qxtKbplyzzJCdA
v75ouAQzHiDVjni4mDVH12m/lvP0afn17RBJoIxzpn8ZDZE/pyO6/E1kBt8t
6S1RqKVhVzmsAcQzyJv3lnZTccZzataL6dOQten3J01LloR1QMPbyiy1Zwi5
Lo0uQmuNMm/s3x5Gq3k50yan2wTpjYe1ocX/3FnielRsypXg4RpyBxl5C0Rt
GizErFa7Fs2xL1ihZ4U7G27Nwto5ZM6iPi+iApTxzxbXtb7a6qRtwYU4Fk5R
3SPPF9R8a7nwGlK2nxvvEwS4Es+egng++09eAyTmVHO4m3XZdt6lDPIug+S1
OzoTvU+7TJHp1Qa9FFPB0eVvfr00LAE7+vNq+RQ8xVSEy2MfGpHroH/0/381
/cnjj6q/KL731CclHBdQGa9LaMSG8hYIr5SXt6Zrum6HkklZlalQ3L5p6D9b
HbaPojVO8dlc0jY8cvfx37g3haKZMX21BiqqLylGirfbWAJSZCJmUuzZ14ID
hr7R5PD29oxGCqG8x/A5Wtxatc2FvFjR+yPqHmC4D4pUqpvOGDofe+DtxYsh
CX0arj7TVFq/w6CpT88lelfMt/M2TtwG8QNzkaoeAsGIgOESAn3Tx+WvX2CC
fVOdewB0ei0FpoOmnt2xQzgVTerdfP8qz8p4P3rvNVuTJM3Ju49DWNPzySRn
2Pk3x+VRQK0nNE08Og1s0BItKDJj2kLJBFO+oZEL4mxRZvUg9XWsLx/y+aGS
/LrBVXZ79fNCCOQVGPVoNcI28TsjKfp0TuOB1IWZkcaAHhk+1p3mdJfpdXua
HdreCkO2rG3le2QECZ8e8xseZC6QTQF8rWBya/dYGjXPAdwLrGw1Q+Xu/OcO
rspFYAaVLQv9ezjsdWhwBV8y+YfPJeKHTaQK0Kvug2tnKJEz3CUETyuCRf3F
c6oe30dMLQ7D0GqWmPM+fi3m/h9elGrur4n1Lv0kVidbKmPo9ZkcYNcrkGuK
mOSg59KcHcbfXQC+v1VvnDjoOqEedMSpZp2iTh0zl7IKatcnJkOMNOuqm0ax
S51i++U5R9FN0ibuevvN4HTBr/rMdnlFcH4oKErMCxnn++hTZSN9bkwe4Ibn
HQ0+5dYWWxYx7CaTPd46qFHo66QSTV6M2SvCbrVPNoKK7QEvFyo1hhV1JoZu
r0Cf0opz+jEupgRWUjvKdMJ0ofjejCgFjJsuzX2TJR33ehPr4xqWOwA4Yqts
Pzlqa6j+SGWaWoP4urTyy1KW/jirKtmQoVN4oNXXPN5ZwKXj7NmJPzRzdtN8
lxwsYq70Rk6O5DSFPkjFm6HeF+KD0xlrYvPFe96iPFxmM/T1tSGoP4nhohc3
NCr/sY+m7q3yjuC3s3WcwAwPY4jIwmO9Cw+mF1X6609T3oZC53+vxeOPmg5C
GIcbTVhQzO4zeazFADPGqUh75a2Zry/yvQPSqophrLu5zT+QkKi3n0Xi/mv0
F2teFFoAeqReCmmpwRlI3WbQhhU3MZK4RnJzlSWAqz8tyXiA8O9X6Wq+nt7c
f21rrXewqTg1SUirCuIRW9vOg5RSxRuZ1Meur3z4v8JuUsjoOpiwqH64SSCq
BkZ+DeDof449LgV3xiVN6Wo1/VcoApwNM+/tM1G8uzGQjHHbe1YFBNCNu8KE
QJHRt8vFWqwOx966syOzvjr1RqmQ6T9MCtliaFhPRsq+xnZZ5sML+r7fmFdA
LvJGJzM+a86P2MbZ+pWGO76Tx5C3q92IuZLK+kBNrBUvrPK45I6W2b+sA+jX
zeyyxXDh+Fn9KIvtDZPhyh2XBoCfDPz4GunvIsAhLZWCBvzaxnq4zsyt+u8x
qJF+Z9GkRznfbH2exQ+gWVby9+g8viMorkl1cA9ZLCAQPD32AC8elUHaN79z
E7l9u3tAgDe0V4L9kIgFDx033z8UB0AvSlJhscZNnGX4cLtRZ0npJdw+jkzc
eJVFOBY81RUDVyIZWJmCJXNkTpYfRnyCMFVMc3ILL10xEW5jy2k4FsRqz3xh
9O/UP13c4+WVAmllv+uCczVMsgu/Oyv/IL1KboI4BFMzmY7CU6/37CbwKfel
r8Tr77qTurqC5WZ5Aq5Z7S4h/ijRRlnwYZgvYvuyL2ttpFsnX8oOZHJgoSAl
KkZm0aLGRaL4wn85ZBGEQqm+nH7FVLyiDZFHDxAux2L7F7sbGlwnPrLVRVUo
3va88cCnNHUu5aBVQ2UmLSvUHjMwmxnZqrkVzMgsecRvc5jPh2Lwo1Pw01Qt
kppCe9Q/imBjE3a7lX4cVbKMW6J7+Gj8xp6PaLGEoTYN2o8JYcz7C1il5AIT
p4opI8/c4lvrOs/bpoCG06GsqvwHlSRTnk3GMkbhaaOjHFZ9r0h777ZQIc+S
z5nXZyoDTl+dPuiNUbeKTQmYdLV0D6z3uwFzlhAYYT1Yd2xMPygwL39uK7hr
95Bg84i1IPou3+XcZOA8beBjAK+WlQvry/CdQnaim9mbw97ZkJisFxvoASgR
ltGs51Dg4EYtF2z8cuU3a+v41lGg5d9m2O3uZk5m947GvX8aKk//4LDfdQ1x
PSsczO7gZ7niaxj2YGXw5gf/6RgR6o70yM7JvML9nnf8641zCXbR2iOeMBIs
+6Cgjp46MGqoLA8faJ06z9WZcHeEFf9Zfm92ovN/PuLghevXR4Nd8wfIJYpV
zCDuWvB393SX703nWHYWZZD62VOZBFPeEVsZT7n2aFx5N616uAf7OWOBtqZe
7+JwbJrbBbpdVNAC1yfq/IWvOlKuVKmC0pi/ENbQth4byrzXVkLN5d3WcWmE
kMWkLKdUDIduQoWt0qbndwhfDRaa/G6HzSTczFolRuu70lxjzo6PxDkJIevp
S9mhrqF4ut+ev6StPUPBYsLy/GR1GmJps54YqAkTmNv+sHh7GmLSWyyp+Atz
bk/EhrI/dVQiPtYPrZb8qOMLD/9dtRhQqhGRS1dgBBr4S1dgkRH2DhTs8M3g
qe9NSymIKhmwbi3qzqRm86SHYu4g8Eq2Fe7UcSXhCAKcd+a+Q/lQwi5BhkYs
wkmRF/UuJKpFXj1qHME3UbtiYtIKQkYC4cEM6XoYOssYl4GWS1PjdtoBoEHs
jU3nPYzTZXbUD2rPU5uD0M58nrLT8zcLZie3EQslF4KTJj0EvDIaMGITyCo7
PhOMHEj9ganB9mf9/+Ku40SnCDIxS+y+Jyii1CTsQOyADblVTuyTBdGB8377
/5QmqRngSuQxpYVBg/C+D0KWV1DuJ2W/v0PGlUZ2DDxsA0LKktDqDyLaHfW3
DG13XpzvXlqWiBK0FprtEyPQtPBy6IgPnNVIZkU2+OGwOh1cowQQOnnMo2bk
kjXsjWdlnSsZ6a+3S0a4DnTqqJgDwAJuIcvfmu90jmTEJsu7YhA2bcTPmYJ2
HeVyMxPylO3q2JYL6CSLDATZHJAAnjbT/ARaz5gRsvZdR1Q1cGo6WwfXXg4C
dC0/mwnyUN7UR/kMZxeW03a6lXunnuthnRsiq3V+vWa2z9TalWFPhvxIEsHn
nHxrMUbYoMY5EvtqqO8NsidTwPOeLqc9NVvmavHeNFr3GhOPMgNOPNQLpgkg
YOBWXLbZ6o/xJZ0c6z41HhaVMKgqZ/INl0cCVjFbQy2CaueuR5D8qNyLvflu
ugPh5c6+vjZTvw4FQ/6ouZwTKIMG+LP8AZK6wJv8kzmCc2+t6pL8+FBtSugB
fuUWLdCZQLOrOYisTbl+OEYcTJz4fM7hSDPXq4loqwu4oZhLWIqWvqaMuOm8
TEj3cTGfZLuMNaeLleGXYvNxKhMpSg1It4Eo6F9yDxLpmoDWmdL/O2Gu6M9a
fRguk0k3xVJLdDb9S/cAeB5S0qujT7AlVm6tk2Ubg9MgshvI79MOe4qSVdNR
/zb9BXwQFtHX04Ai4Hlv3J8pjRnpqvAvP9BePq9nWkOa/EjXo0NKKuZvD6zB
6mf+bHodSkaRPOFiNiVkQEALLXdVBUwPqPpY+ncA4R6xOu3chkFf4k4YVOMq
GUwxgFhY3eOnnAUKnw2rwXzTZZuLHLs9ocsfCvvfKHc0m+KYJA1g7fEAJ/gN
UMEeBK/77lHWSEwxH7kQXzi7RO3gYpIkRgW2iOUXFZfJc4aTx0O4CYQqFlDS
OFtZSg+WP3zRj9dYlV9xTdU1Rq5AKmHwxmM0AoFkhPxk2+c1aG3rzB1r/zaN
1nRI/LnkL/DbN9lLJSnSKJ+Z4b46NzU557Kj1XHkRAjrQwV4PBTOEqD+wjTy
HPX+ilDR/Jf9+COwVBN+NwQqdrm3Z5x7fmA/dc6oCgEGVb9fxWgvyf9ZZRaG
Bd7agvwUULsWkMdGq4vqR/u8korKyMbriyD2Q4r6/UDlwECT6weUuTPHlTEj
5lrQRJSMjy21sYOxU2Nm6KLT6fX0y1W1Efeiy/29GjtrWHLV7W+DKFHGXyJb
IXw86ADIcFA1fV2jBJVg+vwlVi8pj6j84dsLNV/qOJXh69U61rMvktRvlDa4
wz5Y6g3zMIg6WlYq3MFnTWtV+yqN2LcgTAAG5xpEsTQPrgNuAPWiTAU8A2we
Hli9BRA45aqE00CIhlHxNvjtcXqOQ3h0xTnwP6c3t5QwqXmkdMq1UOAXfbs/
sRwZiMaIwIXZi0sfmMKqesOXeMqdp0MdAqiO9i2u7soOzp6TdN9M0ztcsfhp
+nnaZq6lmCuB8XVA5b1WZNNgLAQY0fsXhqnnivK+VkrKPjW5rnvqQFxLg/2K
ETLj5FGFR1astjdNtt3scAlTRioRdreWmK/N/mPqvGCjTpC0O7/eFJYalo2M
YILHhNVuBu8mlhBg++wm82c6WtxDh/fTFU79x/KjCfraZmRtvTBCIGGFuHgS
j3wH605ezsumU4VTNE4k4J6YEYx2681X1YmWRKr8CQQkadqc6GANgNogeGZF
JSSZRkVNPiI05npkNyHoLCpuTvn8ICYWkk3E7kvovjj6F2b3bfZ9ewL4MFIF
M4R+s3Obk1LlDBd22aBRrZ5dhK1EzBx59H3Rzh0iux4WsHjYlEzPmhm6vmcj
vpK75s6bsPdUd+7wCQzeMBRtNXehAktTlb5UhkqMjp2oPpk2czDsH2p2lN6m
8ea/0nPn/w3LcP4wZv4uLevk1pcUGk1glBDc2dT2lmZPNwEGsbiNs+w604m3
tPCm8QHyO9CNr+g1RY0j+MlcGAIkW/XE4+wjukr7CUGEUes1MxprRrh8oY5E
PCi1+A21c2z+au/wWFnt77TsJrclrsjd3YWR7Akq/rgBv32rYNEY77S1bsn6
+KacduouSLH0S5OX/Y5QWnA682vj84r2VP1Rt0kykGiufxuNzmRnj+g/wAB9
iYQa6mvcwyQDWM+pJB8Q8kdzeUSeyRNRX0QKFaNpKBzUad5AX5xmNLXoH81P
Xtan6d50hGsW1TDTP3JtDSmV9sIS0Pb419p9tpZr/DpFpmGvpb5b0r+XYVxQ
YdT0WjHSQpa5cxvbYT3C5o96sRQ+gn+EeaHfZmfD/ywUhvnOD7zVcDqbbfui
My8HmgkF25GCE2eWRqhbTxO0ATOfx000Wk1fIJPy9/7Y6ej8fsne8PQUWG0Y
hUXPH01XbFHuyCJuXy+9S9icAs31JHAV8W4PFmKD0sepsoQku4TIqF517Ntk
4qAKbOqVHl8Ab4n8qlddU/VWsnk5yBL6ePs4YGvUf+0eXCeQJViIsgMY996z
qzf1TyYjewR3RqcmUzxCx8lZHR6jayDS4gsrhdXDa0+Kwep1Nbejw6Wdhooy
0iy3OXCSeV64akm2p5ElwhssKA+6WDggc5D3uv5XfCjvpBVtC25zVfR/2sfv
mvd0fce+X/XnaAclu/CYwX7voRUI/Qdx0Thvly06ADE2g/+/+WziRwiix7WE
Lyo6G8aXe9lnGBsdGVXO3kTR1p+p20qZ5bovzmj5ISbS/lSlgY3by+n55rln
lh9GC0vlKzPyIAq3+0u9qVcjwEc3Y6jR97gSGxxm32Dh6DB/x7iUAY+kik8e
FUx2OnJy5iN8N928iiqkDY3epJvFz2rxbUGp61ys8gD20j7Jd3MBhdlTieKB
X8LrLuu8ET1s/kFHVr4ubdOBXsJCad6SrPGObqBuXtMwJ4wqVC8posqzASEg
OMe6idicr4bqPEz27NMqeXW0cMd2yW1ucDuJFV+kccU/4Gm/ojbva7I5FFZH
T5HrXqnnkNMIaUO/XxhEMwuZEhL0b+9tTYJsb68lF0SnW6tlaxV3KNBQf5yM
R+f1TBwgTrRupDT7/+2dTp2euUthCCx7tVIwfWHd0mbx47axsYXiJ9cLUdoj
70gMoeHvoK/9XZtm+im0rwXA8N+scNdXgeIaykXx7/EeHdAemG6LIGenJaMW
Yn9R9mxruemh9tMP8bXLFq1QH+NyaFKY9cVAfJCjtt+X44wefVqqyU/I6EgV
BInuX7HAZDqhkYR95KdB9RIKe+jvVXgNjbgL0wRReOL5HiKoZ1auRw2qYDIo
/VsGGpD7K1BKmBgYTP0j3GZbU73ggzEc/mTXc+Eo3SUWz2UATS9cLemDsEzt
lL/OykfUnlom/FWv+b5+dgp+Rhlkwif0Tyxsy7qTzF402Dp8gqoRUc6YrSsX
i5K5ms8yW0m248a1yTisU/NoOeX/CN/Gqf6BxVaTL/s96GFfFX2mGzz2+oRl
dpvq2FMf8M0/ZbMUNVHwvkUFvdO9OXpoZBh0eAdlwV78IrvXactUERCs33aK
bDG4u07MZLO0ZoZRevtJkJxa9U77iidhQvUClvO9rLbbTFiilIaWyF1ipfHJ
YkT434+8tW3AlQYxN3LNG3Gn0oEQzYRIt0fm6xDTDBfgWix/TUF6FbP3nlsv
da++//7hTOI0qmFvMB7GBUfbDi/GGCqN348UJ1I5SdS1RtpNr9/WNH8YNl4S
d0dp2MLx2Mw0ncgvPEWZ2arm2wk+2YdF85WXe0BfdRdte0PtmohqRvq4thg2
bMxuWWuVlifbrfxvfFWt9EHkgFecxyTduiNKsSt7gUq0D62tZAsIAWfS9xPy
CQsnfS2aCqjUGKS5+Dye9FhQvT0iLC2lMwze4jYIenKk6m5V5r7e+pD9WPQ0
PR2qHrtsqVelhGBTVHqUjkyb6TktJ4sKBRv1q2NYC5auyAEpTrkoNcBsu9OX
yDQBcysaA1JxHVtj0OuO3QZWqZH4RjyvVpcbA08mAmZz+QzPhSChSJHleIrU
lWTwVysaNbuei4IT7UZTLhGLBC06hRlgoyDaDEzcA2RFWzzDbI5HtU9lxyG7
g3X5hoWnefi7kv2+7G0cMIjF2XnvX1dafzJlZ6gln1a6QsBZchOgHY40Gd9V
nKTpfjmDXZy4B0A6J1hVw6LmyiIx33PTL7bGSj1sjKogYRDe/0bPyvJN9RIv
4N0wMqM+daWDx/dwqu15PoWetrRDG6mQOMQrB+vZCXXJ+zEghVGsKDiJ6f4L
x3I8HuU+BIkV9F9VfZgwPok1j4345mJJn8kylEz5bvB09kRJNWSIJMTIbUMb
O0vox3/dGhN2i53kwwU/9zkyIFcbbkD5tJfTtjXvNxYNkgmlluG+iVKOxYwy
JPPkSef9CR7FRqpYTSyhmqiHge70lhgNfHQJmtOaGNXi65zfozF/8tJReTOA
Dz+A++HEYKIcXYcD0++eviMDRbTyn4WHEGaaQG++9OhHj8TADdfTYOd7AMLU
k+ZQGRgbQ+NptzOktnIG26qRQGIduwjVkZkvDU3rOZPWRZfN7qBP6F2HTHoE
P10R1RWYPiiaBpU4TB6euMlqQ28/uitR4YjqOdg0TboAwHb6UOxxS0U+Ad1j
FNmknVDY4zsZDRhT2EyVZcSqrsU9h7LZ5gWi1TVd2eDpyGilQUoysyndEru1
Es1Lev/Bc+JMG6WWuyq81EkgOYWmXH+hvU2XFAoNoICzA9HQ+1BIhMMrSQ0p
O1CkDoEt/4JGjsS2PWAJyYG0s38PZgkn+s9w4puyp7zPKAiKUYDgp19txeiU
L+ISXNZX6ErSMSq38+ZkdFSUOKHjL0WTrRrne0AOL0iWTkaxYpGzokEspOeO
R7Vq6S+S78XeZZDKbmfAKBu8ErQeheXRGmzMS4uExCK+YOFkw8AeSldPzdHa
Ahdjzh3uslecM9Ent7SM0QCUCmzeO2cmZmZAHjYTa5XXG+BjbovJHjQ9C3NX
vL8DW2oWVHdiK3UAgyxnJoQjqpf8iZ1B2gQ+opkfLNOazAOmdTjUql3GOszp
/GadBxXtP0bz36sjOL6JFjb3dN5OWLghQlpiuhSGeZPwj9fSNz7175Bj5G7a
EfsSaTJcSGl2+8s1auOSgKtXc9Tj0JZh77f57xR+8eZZ2cejXSeIQfymDp9p
VUupJSmvZFMdMZQx4fM/jJ/72EQzIPg70zVOdkxqMLeqGIJkjtDb2Rxfw7Ht
caBiG/Ubdb2te98qNzfzVlzjJ2brY7vsYCyPm57UHUaY/mWWBhAIrBGZd4Z/
Uqg1kwCvr0ANZXD/n2Av96KNnNwmzC3xgX5fU0n6AQZZh9ArVAT0izZu6OZ2
NXk+Sg/KEM0VdQx6+LgLEmy70a9pfLF9TWOxsKMl8aBaRHmRVSIdNMYhW91M
SXg2p4ZKfZMonrZTXY1Z9hsRdK4qpeo9J7nrgGM9SqMZhGP5BEhjXB0ZX6Au
oqnlVBIjGIMoSnokuycknHhTcqiq0wxrSH9fDSdVjqCL8Vpljk1WDaSar8kd
Mcv2/mhf3UA1JCxUaHKkqoR3txlrC8qkPapoSb/qIZMQvFjfoVyKKDMLvP46
1xTWf7gwq+Wqwcos31tHtok1l1u95WbYtq4DUg23jP7yFlRZTOQnsI+HGinJ
UKv93uLZmct0Wyc8c8ZiS3fFUH1t0G5f/OQOW0nxjRmovqDoaWCqUBXiafEv
VunHr46uI5V2/No/EyOsjHbWdVEKaS74aVgb8DmZuqjGeEP/Dijio6qr4iTB
E5c+KqpAmdiuNditzvd0IRtbaVBG33qwbMPPluVFIIgbbW4WmwBkpCjKNew2
sidIBbkYwAkyrdcHTxGErraHOpetS/iTZVUL6yvCAb+5qFpEG9Dk07Y8yBF/
YbK+LjQiIK4vBhqzD86a389jmtKgx/+UHXXVCoOgyP45gVDWQ7Qha7bdnrS2
5y/4QHOK0sgb9oWfQ6A+mHlUEHt5BnsWuBF3PMpEtsL7GTtIIEqDePVKACOz
5YAqqNbykwkRCXaX5LyoZgkPFNo/svFSpYy8DaBzesv9nVyK/PrkAjXCMkfR
4RltRki/OP9GSBbEwRjtk0g16pjwgVtjoay8Wt9PTSBvWFXXyVhiKGiGrADw
4zdijRJw1AfjLUXhlDD4FAesBf7TMS2KLcl9QaMAh7X8IN7KlHToYbeCiIVK
JqDE7NPJPjVuozuF2KVuG3GSAF5NTGA7MmJRL6BMqXbuuFb3D8qSKCWtoSyt
CQMZWsm8jjb/tY/t4Uee+1bbsF5VLHw0RzoEaMnCn3D0fM3l2cHtE4PQkvSi
D0DNmJbYNvcvSinyUerKKzOyqsJgCzapYCaXD0XUQZDNTzyUMThXUJhhhY2M
B9fs+5LAuyro+MosbeFg/3qpZKB2p069aIRloYTPO7Dos8GBpt8PA+KXU2tW
8CvXG9kAGFL0jIPl38nySQ9OCVvPhVZ+fAfeJG9MC3laYEgfXu8exBncGTVC
AzcoXoXlQ5GMUQ9NbPGnythCwLQLaUiYZlUQOeITbO8BSMyjbn6Duc7NZpzL
tBVjOSzagJ5mPyrlD5/af5L5HjxmupCCYosEH8QKIgO7raXlO9eVaAYaD51+
B5phXSRRTZlC9RNbIanRrCDTgOOl2uolAOeN34xx6x4u8+nu8CYfeepEoNc0
q5xVxkoEoGyL4DEd4prZjqHAMW70memNp+zxFzWOBOeb/cZgqbCIXwfZB8rY
q+XhMyKOUOgQpjmIpqxN0ORP0mjNNcs8vcC0z5hTDpcaVTLWAprZWc4zuAdS
wLL9njT4z+sNIfh4FWVmISl/ME6T9xfYUheVS2EzAEnGDfcuiEZrQqn5C+MY
CqwmfNtjJyA26woDhW4OQ+WchLAfnME3es/eAKLUy6ZCH7aIVTLfEmmrIuKS
HoJedmnPtuzr8hW8mOd/tXwhaTFNm6VvkBQ7GV0G+yrr/odhQ2/CYS0lVtdN
l0h2aF6lROUYkuC1iC9F2eJsoC7RpfacJf/q6PPt1J7ZtFjN05gd1Sx1JIk3
H/uozasBkTiIHmMSmY9I0h8K+mfSZFuASsCBl95mDi/bsMuotvjS70kNV+nB
z9UCFzmWTnISnxknZxFt66GqXT9MPYCG0Utpj6B6j1aXfYgo8hOhOUPzVPAw
97Rt5VpsiWb0PErA4yNlXjDzg3q1+NFE2XgAnvSx+ctyN/g1QZG9BEDWZfCr
clbMB2/ECuqAHHo+dZ2WYi2xAOX7t+JONgNrZnyGBZnZ50mlL9YQ0mGkcpHN
nTWh489e8j2tacUVVSM1WxMuIo1SiOSY3OWhMC8OcZBKNdI3mHkgwNNsgzdd
BgOeVzZ0mpB6yz9UbxULgs0QtLBncHarbAMcmVKTgQAYwc9z/nlWU4Mkk5Ut
ZS+m+qupfJxhpQZI+rFRO4sEUe8F3gii3Fq1EbDwWDjV+w5yFqSsaGsP43se
7TdselYbZbka6Vl1aWAGI/gtllqUJxp2jOUAzjmu6uYXi+ENfDpv4FAtcHSs
F+QGaAoEPmfUKYwCChcyHzKAW2mwKqRofpIqXoWvI4QSpV72rB7w5hPaHjo8
5Rs4eiRsYioFIJ48ru2RXgzzXOt3rIanXk3OGTCNM6IYeiyWIt1SwY8pGJ6w
vbtYQtIFOEMZtceHSNW3FgJl8MLi+L5dsoXvYz1rQrn23n6ebVCj1pTZa+WO
cvk4HH7UinTCji/FGdCOdWCjC/y9tZcAUKQIvd8JP7HUSrcLMBmz+Ds0927D
rVWjKyNVDUq8GlZ42Hi+umiEFpV4LhasE5R6kxLCDapN4vBNqs4c2wwI/+as
gxVD7pIFXCqbEPVc9f35FjGGXZJpaL4IaqY9mN75zCnlgOkAmYijMoZ3nbLL
5Axg0dWF4okchan1rWDZJ9Dr4NFC0N3KdvjR4Dke49qs1/eAdt72U88JZyKA
Sp8L1qOxX+yzQUuxe2yrqcJM6oMQjfgQU2ucLkzkMXWON3JcBI9PZvoCEkot
/h2pwEvhduhrNimcJQSQ/pKqe07P8y1CObrbaHwtIeK8l0H1e6OwCtBd4ZTI
k9beDUYALhfhxuCavj8iGn9FgaRe28rP4b4zc0dKJvuVBV1xpOrXhi6nDQLx
GWM7b3QEWgsfVi9pzxSuShRoSox6rmhKERBG98Fn2JNt+SumbUVg3ZNr26LX
df3ulOqxuhJNERXWuVMUcgi+ZXZsHEBeqiYac+7MRHCDpEvbtrOlQ53lsGmu
qheXaR9KyNueEQu5gTGgtJvLqZV/Ou9kpt1a71OW4IziNAOwAkTz+t0wZUGW
YNVWjwPZrmpFnfBHf3k7gdYVzWYEyTu6k+D7PXpk/1HMyDjpkUsQeqYBduJK
x6LgrhUMgOReBwFOUIF3InLPcoPV634NRDkCS2zK1OTH24c0kMRtCduQTdtJ
GVqe6wuwxYh0Ac4K01UeAeoH8S7TYX/LPMy/aDOPRmxHNGggIIX4gzuoDDbY
q77Xgn0lrGwNRBxN2nKSoNIpFPzpIjoSk3edy3jPOe3WWiAa+/Lzoamb4hqv
1M1T3Qx1ugBRt6tA4RmZ6XdvAeQW5k6vRj008IX5lXEQAWM+o8ChlcMrQC+8
xzCIHczdUzOwcWoRNh6SvM/uctAXUTnxBgic0GcRJlusV9VdweCTvXWr94VY
B1ABhNlOHXrx/V/WJ07HkD6slCx736DEbmWA49oo4v6RZr1UMZ/aOk6sUH6x
DT+NAPFRn+7Hayc2+cbGiJREiUEJp9mvbLsa4WskP3bg9AiSh6BcGnHBprUL
wQM3A9+yd8UI2GV2ru3Yk5ZmyJ98iuEZi2cEd+7tjBM+l8CSjo2h3Bd0HACK
1Amo3YVYm9ip7adssmrJhfobMLQJOXWi6FjOVptGnTynaooAeYOQmhBQUgER
nFHaxVq5vpGAPMyJQLDDNuY1EpTmU0QTub/Vc90n4Oi48rhqeQmn2FKBw/GI
TJ6mfFmb9naMFMS+QpTTkHLS/R3C7p2evunDeYMK75ieGgNYZ6F6tyEURiU/
/NnmVYyCSHio4WHP8UtIj/L8h8amQp8MsTWudGFGaZqtztB3FodDlL63xRKk
c/G1sPvyHPhr1t7H/SxmAFlG3qP/IlpPB05gJNbVz56k8r5/uaWZGOQZvxwM
orjNBrj3FCLaftgsQLCPITzkdBmiqStkGz31iMPC/xxvqMGDZJ9Ljzrag+ER
ieG/QFapLwH+8UfyV97APCcGpHRLoiM3xndlptz402ZG0K8ZfvDbWtF6ueyU
qMu5P9VlBZ3H++rjTE+ufE66iPn6DbpmGSy2JoVsTA0saH5HU+TxYfpJtROc
gH8FBYfrkQ5nILRqa7Q2fkO5R/kPhcRLkQS+AKiYRBg2256vyqPlcmYMM/R/
o2UiLVJr5xdGzlIJatHF9ROm6c9g4u5Nn5Ghc5o2XQRjx+GUQoZfJth8kiFt
x8hBQbombMb9DIYmxVkWgpVI5N8a1H3N7L/6F5FXvZFAKJU6R5qUaHANqUWo
ivn8bUEG0O0WYhT+vGubb9G73PcLZey0kH6SCxUZi6sPOKyEQPxhblCBp0FS
cKF7gwTDouLt4pWMYHxZAGwycFn15P5KpSHhBglz0FHdeUE8EHplHoN+Mn1L
KI5nb2TY4Kq//DT8fj7pTNbLWja8j8r9HHoKBHez+3DAFuwNANj2UDnzoFme
fPEQm4+S62C2AR66THgdMvMZ+Zw/IXpg+QypED9i5CBSm4D1PJ5pJ27l9L2z
eIAFBu8Up4y+WUhwHu4ZRWjQUkOCoXYGc4LMXhF9e2E0VPk4YpwOR3Ku/pQY
hIDmKRmr6zokugFyezlZKOPQIg40utpgQmeN3QDV0unyW+1tQb2HJ8o+7Vwn
BySkM7jn0G/qA57b20V88GAXkVm/g4D5wHz9LwagFxe6frl93tnEJ2O8VCFV
Kky3F/D/Z9WiufSlSyvOcriUSjYCe8DBXbHizmtQyscbPq697lEy4aJriV5r
JS5HzBUVnrNY6RTHoTtpLsqhouwJ4g8PtFKBEEIkfdHSnMguZu9rZMvydQDu
EKml8Tr/D+kxmzV8BL3JTOSAWM2uqJmZsiCpeeEMOS5++3DhNHM3nddazLNo
YvtDxxHXqAwIstTBeqs9aiTkEntb8tC+p6dCNKFY27aVeStDIF654HqcmyfO
VlIdSKAeLlBUnv1ETAUUaSto424f0RQeLIYo5CehUkSTiGRQYCEt0JYrxs2m
qoTqyHibrbcEYqs8DvZNk4sNr8tLD18f9MoQx8odum5p01qZNIv11E3GP7wh
BJ95Yt5qwhUTBo0vyd7i1p8R3LVeVsYZwA+7LPtKbaLBWR2v5ghzp3brctaY
D8D0wI1m7/nQ+Iivq8gAyt/2rSBYgV3Z+q6WtieIG4a3BbUtfXYSdeIP72XS
FVCyI6Ay0WzhvUgyeIgEhRl7sNt8FsRqI56v8CYbr1VHXa0vAUMopLbQvfXe
7JTuoEci3ZplJBQnGSkWl9ypoL+fhzgzPhkQ0cHt7RhvG9b2D2c0OMLDcaKx
Z0SxP2/jejGIABKcpq6safXy83xvkBp7OvuzcnNQip2mcuLw0TXQALG1IoGh
8cW2M+aUJCcMaUlhhL2ilRe1a6+6wjUJA7GX4a843QNe7IOZUN2o0horRUYD
JlRbIC1l/zqhYhlPG2AhF+4EEzCP4YEc3UadGXmfVazQmhxr1ROEyqpIZoJi
D6b6fKxKadZbLD2JctZYoqe84MsgDZhCcQIHyXo25cPrzkaIElfVPvPJSsMV
/qO1WUrdcGdhyGdG/iUADwzNoODq1pJnpg1/uFxWSOKlrUS6D6s6Et2bRQB/
qwpBWHwE0gd+PMJUI+fCTgPUcyivc/TGpVZzmqtlPANHV+XNGvuKVicl4l5z
3L3wKlZTb4v6OecG7kPd3/MtQwFJfih5TzqWMTFEN7/kFCXXPhbw1vsfuXnI
1yl+VVEkH8jKKYKg0UBDDglN5/bd3/2qpjdK83B56zOIIn3g1cO+YCBVhduZ
EzN6H9MKOCy8sWsmEs8/lDiJv1tZ/qMy2xb7vqZ+fzhXk7ENURd5oKwUcNsF
hLRXKSn55RIMb1w4g8zmV3cY2L3Y1NHKtMW3L458fEm7xiP+ub1Z6rWzrLGf
XSsx1mKd2UPXe1GJ6uzS6eBLNQva7CrHAOHwR7lA5VqOhBaHAt00iZljnb+l
JVC+bZv4/jPTfIeOQfv0zIrpw4ViTxCm87r0Pt5+z91kY3WonJIjUF6lj4AF
gHkv211zWIPBZ6rHX4u4AtshSEoMxXEyEJlMEWoufhTMLsxsaSpVMsklzY9G
KD2I6WzAwtwNCmjIYKjadW6WYRLCMWkb+upZ7lLhhJx+d3Pm2dBoQifklpYg
pN+BBLz6DjcZuB3c/Z0uoJl/te/X3J/O2y8F7b2IeWf7ZVYribdOk5UI/gX3
iLqVvXU7LmUugcUgy3D0L7JEsNlG/ZlWbaF1wLVyi2n9KBvZRw+2OAeMBRrP
e+K8hSS0Al860GCFOTlfWewmXK13IzXq8FjCyUItiDa4sd6A4b5OTwMcAnKo
WIJLU2PtJIHZQ2ZImNjiaWphnRdBaemCqELETmaHIl7spXP0TecoQQ6FsPjw
SNKKQxR7XwqgO8iF7H2N7gHx3lwyxj99v8T1nmDRrSQQhzmLyfKo79ThdIrx
uMh18hZxo+5Rg62jykg1JE1RhUZDsId/etUbkG8MTkb+1BeXiDI4l9ZsL2KI
gBA4TM2IvJ8qwElDhMYxalUfWM1ZCevj0EZ09n00IBNSPUYAX9vzE3JOiHvx
85XOFS9NUW6eYnLZGWxlXsjxXt7GGXfSAqbtGn5vHX+NFhUN/U/5T/UZYaTQ
qXGACB20Cc1Qu1x8eWrrbKpym6aMX2h+/Yn1awFB235JMMOnuRyXDPk8KxXq
6dv+M5+EuWCfeBXWQFec39e0BYUycG6LxbzXsrgT7WDjYcKLM3cJBO7VpfGK
cYMpi+UvppJxRGqo33r1VW8PjZRNzqW4I1pNGof+PCawk288boY3QM/H1uX+
XnlHc7hBdNm3xbnF0rJK5wKtOeW6Z+QNVATqhZnYh9j8gP/EDeGXDXos9lEn
3IM3PQY7TqQj22Ec50M6lOwSqMOuRPQAfcToqvMiAGE7X3cQsFAREL1Seou0
F6uDLDdUdmxsOnw9FOqyZvEnxqA6x3VErI7PjYH+S4pHFVPTap8X5c6N7ddI
+/Sc5GV3JkE9OUyQ9xK1jomtot1kW6NN9TW6aT+fdSKnTamxI4SGQXOkZE+D
KT6SfK8yBvemFi+XU7ySb8f4Eme/u+n+lKUfwYiuICjosgXHJeY69FD/5QiG
1JUruSTFK0xynjtJJplarw1HTXdrGYiCkZkqi5b/IHcYd8uFuAtwEt94+uIH
/c5OT2p9Tg6sqlbQZukPmmwReB8LVjWs5/S7LOXoIgePhDM/CCQ3Een5IxPz
UHqw1cAMKa7Stl1WcVgzxrCZCMHC/Dg3J3WfHsiuQiIJ59H2LFera4yE0CP9
8cTLZzolcCGDUfEye/e0GTAp8XNC0ADXlvqSVolaErHz7lpdiz46IX2PS+BA
awPsdVP65cvCE3BeUnP05HSDwwW7lvrSW+WuOFusRf1BkOOWdpfC9DnVlIw6
l4+kss9gJFAKzJcsrvFiiOB3c/HoISjE9pKntf5hzl08F7Wcgd28s35F23J/
xTnupnDVK27xJ9b6M0d2Akx/fEqhDtrrdXUyefCehjhSbEjozPv8I3K0Hvki
6xugRgn9RpAONiOiarfDaorNNefBWBCk+fUYT04ZPE7Ioj7ATAhub4rFkAU+
E6brFqBLvzf5CenvPzscTGHBtIcl+0DG8ECT+NVe0c3afSO45AUddYbL7OLt
Nbw+JVjrNf5bvirtZsQh80geLyeOqzHWVxoQXa0WQjzpNHY+9uPuuddQh3zG
e2Zkla091EHFQJ6/XPQxWjL5xPCCdRcNQbt3GvQXA50G3oJgzjQn7bmbgmZi
xmWU6tQlrIWLJotyVMD1QpahknQ8yoyLQ6eCOCaLir1adds4+AeSruuBSvSV
mlLNRHx0hufPNO/EJmo+nCKgU7qHgLb8HHnerUeCv6G9nraXL6kj9LJvdW8A
+hKIV3F3nTy9QrA4rsxD4HyWcAsWmxIXsIXFucJVccOXRaX2LgPDG/69uRBd
gfdY+nKE4fxgwrCPr4QDG/Z4EvXYGmaZkTrhtIjA6iokgaU9KVJSKDoNYOyn
fPUdG1aO1SiOiflDd1uOhPhAcLoGe0YolPdYz69ptcx4o81vtcPsMm2sCi0e
beLYSae4jFnylULPz/VjznOkV7bovqjipLKDulWKbnwvY7Ys19nEKBFngtVA
nnlcxGPJRLtkMRa7QFxhO3dbbuqBgV0iqW0PC1MG2GhiYptR5J/LOPNmIHNt
CoBmYXRAvrbqUxFfXhMyeesgwbKkxwoKfi9mOSICGTfCl2ggLlpZm8wXZo5J
RXEVxUkIZcGtGzPXhxJF8+kYlx5He6rD8z1MsQrF8iEgzrdIXRxcPU6RP71K
E55T8fiFDIgOy7nQcKWKmez24L+oOANK5eoBkREEGJsRPDu4CQTuM64mtWd+
ud/4JtMKBisINSK5JPede71gootstHMLqnzha8+pyIZZln5AELYK6IhJOjOr
alZ3GhnljNC+6wjIXoKJrqyPmXJnRdWKR73/YwjjBTV+DRpuar1neNahP4/j
XHBhubKgnyGjJhwXdPSBYmYCH1EYuz+AMWrk1P4h20TGQoDLnU9dLpYd3vOs
l/xFYwAWoq0yJjdSug6C+nAI0yes1le0vRuYirBj7X5E0OG9vx8VJOcoqJVX
c6tyskR1+sGn+nuiMMj8VcgRMBjL51RJSpPGTl7lF6eFZG92Udp9ciRrQxK7
LYrkkuhqZcEjRFy0EA1hW/oV6fcZFk/k1roTZiPCpG1WVXZuK25YRb8Aqp3C
V+8tslInSQF3a2cL0eCsRYH2sg5pLFOx5SkKuZNL58iZvDkQeVi6ZkzZ3FE1
qJzrQ2TLULDnDhmgctI1+CQG8aJN/mWw4JaLmHwAWQBj+RoetwLGoR0/Da4y
5bI8fJequ49aF7iWo0ZVAlCxXP6kZdQNnBbI1iWAc2UNqO3PL+oR98Rcd8Tb
2cPxpOlYbdTRPkuc7yo2qPaeK5qg/4sJQghzdysSJbHcWc4QmpPdXU8v/qkS
uzeKY/9ch/azT5UJxoxo9V54bvZy1GvRsT1oqgiawEUd+Xe1ZRIxe9XVhwFY
wov8pi7OZ0ZW7uJS5YbPdEqhvmT59n1llSkv3glVCUiWLRbMn46aYQvre2k8
qzfnY3kJurZ8Qk+1L5bNNs5KtNmnoknLBTwPT3mj2UTNQwhiWMELrQZaVz5n
mPR1MMxr/Atfz+ldPaXNuux6o72KG0go++hk1RguWPVmS0DM0VJCDK3wSVj0
vrSO1L/7a20UYeVwx0GAzI+jtK2fokoiCPFTSIPHwsr94TqylBGNvbWjj3zf
r5jNuDe58U0QrZB33kU79QIu6ZZDW7TGd3DbEa9Si5KMLi2BThVLOv6EJfk6
X1utPDtke/rQ1cQOiJ5yrXc+y9a+H9nelWcJyHbQREEyz5sVq1k1gJkGa9Lv
20uTMzGv8OHQ65G7QArMnqoJomVd8Uf0iFV5Al8WI/hpR8ItdQsoYbw0Ubty
F/seNp9gcqeCRTb1uHWLK6mpOpBdc09d3yoesk0oNTuiCVayD7nedmg+g41u
xqqO97EBIXBsbfcG0BQtpRaIyjv9uDR2E8/+6giZVWwVrloastuNOk9jVbSM
QT1inL2rsBd390JSzHHzZVcbc7QN9WITiobRXy+Dchx62rw56smXdkOQsgLV
2BwnquB3Leh8MKOvF0K3c3HhI1oilpjTtL0/IHhktM5VuS4yj+XYx6VRFoSR
hpUoQyxJUR0lxj8b5EH2O1+gOuHJH963ehuuYzMJ+eTV8APoCHfG9mS3SZSw
xt9q9vBLBD1dwY6BOft7oZYbO2tExTmJcx60oPR3imtZYX/cB5Q/SF40uaWp
0ESToGC6Tt+eupCAp5+D12VT/5jZoZBz6yo65PQatCH4DAtkc7zS8JuWFo/K
aGEVyWarCjF0+iBvnBmIRUF0ep+hL+S7tNVm3D/Nu2CvXU/YbNs1mF9DuwNE
jpopt6I+6BDTF1hcrvkmuvl7Z4YHDncoNDG+IWu+dxT1BKYYinyZKUujAcSy
d6gFwWGPcLMENd/xBukdxDIxObfarFw/zDzXZ7VFPuvxDH3bvsYDAZ9ej6yq
2nnSFYTQGNmha1pM17JONUmJsLvTakRjhjW1l3VqwPqm9bZbxJJj6q69iNlc
zan5dseEe914ba5VFV6svxiKfEn/qxOmBi41iybzzP5dnHkDZcfInSMYv6SP
sybZGluBf9XFtN3tGJotHL6btNuFkSduvy4bMC8wEJR1tHaFsz6Cygr15T6f
FGpMAWUD5vVpWmgURsoPWw7i9fdConeNC1v0Tw4F/O7iet9man10JtwiRC8N
pODf5WCpgKINTYCrFhwff++cuH3+MdGtFdRZMxGLa32ShJ5cCWHUzw/GVD+r
i9LF/AanOTtTmI0PjPdUvDJZdL0pNWAqTyI+GKBMHymurg5V6vWmNvC3qbf3
mTELEy/G3X8jRM3dLiKx83HLx2t8EV/cekKwg1TKc3FhjWElWAZfryCSyWdR
pHjAIS166wgrKFLd7J+sXFZUwb9we0/m/UMA0T19tWVe6hhZayz9ec5YAK3L
dQOvJGljIsDWsHl39lLGnJsyLPBINz2hoghb0LuLX6iNtjirjH1RJtiALtMq
1EgK0uMfWX8pDLpyStRlae55wj+2735X78Wfn9dXEaLn4WNlNO48/CsEM61W
GMGwkV9dhrtuTRdPRIc3LJZf46qsvVV90oo6uB5+QwegIThYbuTXq9pNfLNP
T3iBOZR6oLvQ/WlEnqT/8TCtrbjBKvzZX7AYWkxW6dYQwOl7JkpFR/NF1TZH
sN6ZteDn+g8zxvTEqfpY6vNUH1W3w+Dp2Uz/zD4KZ0CeFkPlTncm+VWoFAs/
bYjxQN/Gijl7zdt+yTmKCrVD1gf3qTa0bo1PxX90KvSVaSuRBbaCB9wtltYW
PuJ4kdCxvmr+vPOogfGQEQ9l479HoEMMBfhQIUqnPOUnnCg7kGi1mECRQDdP
eq/qGWUNZ7RbVYxtiBtXUj7fgYv6LR8IbSvmn6x5SVgQZVpOHvEdYm4iEdpa
UiHX36NZX0bjplIpxT/ZwsnLK4JY9luLzNPi3xHKC5/LonnZ/YoEbxwole3Y
H88+sYv+AUQBp9i7zYN5jtFgFsV1ebCTyBDRY9VqTxQeBMwUdBlfzIjMePXr
reWkP7EhfC1xLp3Mhzqs1drjKEZnLsBQ7hbnovKvCnBmDwbU2qTOQDfig1FI
ffmpekKTaZXXFrrYePKn7D99GGth4oU/ep23jwCmiPZarK90fw6Y0SY8rO/W
i+Hsy3Nv1qDR+ehh6R0XbzFtUEPhCN1lS0wAuLUm6SGHih3onIc73baTBkGT
qr+c9znqocuKRF1wfMx0QP1pMbqG4Vjxri9JfWQMZHn/yOmGmHqTRK/BtjMM
pkjL4CHKKPOToJNIJ8h7t4IAVvFuxxnjqzDhPwGHjmP23TtV9R7elL4GBmlH
vzxyhmrSzNEErtCr8bovDJu/RaMVBmBre5XM51wJudTY2/hZ5BAblF5DU4gq
Uy0sxrCF7B1Z/Ypmkv56EfV1wI/aOALtfZE9Yr6BOMlsCvznac/az3ugXuow
dhrggNBVN/VFUSVgULOW/gNLp8mJ1PHQYCHnK0EqZtRmX/mCDeLPpCD83ccT
rWaj2a0lpjWYKkBlWNa1sHFeq64M6xhczQ0a2T7AbpuiNTQ8PH5bPsqtGbr1
KaSe66ZFNXBR3GSquRWcWunLk4WuEnVr9s0iAaRW69VenlKeTXuacIn4BRKG
I0rsEJ3Pm7ptDZaOiJYn4MiRgtw2jmxWoXQhoq9RTR+o7lCIypCVE0Ms8edV
gMTuFSwxEtQ0dLmVf8E6tzyCX2uXWwM32E1lNuuhPnkSsvdGa6fcbusiQou+
Hic3VCyq9TAuV6KqUS93ca0HPJuRUv8i/Kr3uyiN9hr3HV6OKJ5uj0mXlEXo
0sTvF004wkpNYFsPMU4wbrFofK2EAF/jDK1E6BFr52W1Ke6mmruQO10PuSjk
LP79sgSeFBlXHDJKogTHUudciHo300w1MY4uBPeTpv1c0bvzyU/keB0wqY8c
UxCZNSbuiu+JpC415+b05IU8dwZAhRV4XGnp1tdziEJ65Fj57s+H2ebBn3ML
I2iaQple33gS51cPlu+8KMYIi01sO+xLnHPE1JWlf2vLYrBRmITY7+dM3kAB
TJTgSzEPV4SvVa4ACTVBJ7QNxaJwl2PA+MHXiXreSsRJX+ghpbgw6CVDSyc7
ocZ5Z14RCQePMKSPIyggmV/esnFa1AyomAuyPIZ+dg+Wl0Ow56JWy0qA4sGo
9r7drT/G/cGAcLAVf37mN47vSh9g8zDKprO0SxpuyZyLEfNsMHS5ZgVqLusD
dKR56D+HV8hrds8/dtlU3r+B75I7cSudIsQU1LG+OQszem/B2524c4QBRBjU
+zt8EgYzwZXmiiXjWFe0N81el/+xcovtG1SmvPQTi0OFJBAFJMOPoFLUcLnb
Le+pqyPjnuCSs9pwVsgwT5vlswrDBBc1TLx9jWji/lEDr6N9WhmhkcTKByfk
Y47kLEzCDK5IuvNcMNMaCiJGYKwTlbtECPvTmibJ7m1NTUpCCkT8v6dvmf3Q
5AfYkiDeF/bcQ4wkGX7KZzi2u2SCBWF2dHupC5Tk3qaLk2HZrCsKHD6jA1LX
u4V+Z0XY6xJcoXFgTTEf58AgeQZ9pC9BPyE0d61EQUolRnK+CW38brMpZs3l
JBXUOR5DT7LWnksAwr+eYHrSIEghlHJwhhu2ZqmXHr2j3atGWyFkWTEUROWe
8fcdWzgycAQOV22XdRwX/4FYfGPvjFezWyF3XnWVsVlYKMHhVhodgF2+nGPn
a2/HG9+hERUKqZ+Ce6wXIO8KP2EoRCtU2xzsodAYYxJ3D45u+QCXXV3ocW62
DFHYll2TQUWWhTRfKBMJHGsvAJqwp3GqFeRMM/yzC67flBWgv54nP4shh7io
NbZCUoyibk3bQ6erHYZALIq/YB/xs5n1oJxBKgUAPkuvl/rDhNNmO4w7TAWZ
it2E03AepZAx3FEDRmvE0gQldqdx819CIuT2zDmdEe7Plv8h0wOgQPYsEXmV
+VtSsEwPUusFQW6d+Fc6u4+DYvgYoglX+HP3ie9VFbD2xNWifXSmM6XquFrX
5KGWtuuSmzPLpYWNscu/ruEoEgUi9OLnKO17XG3Zzhgr4G9Xlj99MXyButN4
g+UbjIH6LzOUV+3fhkh9MqsemBYCEZ2fMgpNHpAJk0880mo8Kgot3WqLfMj+
qg0YnfkM+Eziy3GPX4bG6fh1dvjGlEaqNsAW2M3QCgGSd/m0F4UvK/I/fcdU
ZyJV4s/JTanlRY11KEV8VGQ1XxB6tLT8plFU/wYgwZ5fGiadUhalPRhtW8q+
h+mHHCx9/x0YSTw4E99irYSjJjudcTz87Dn3nm3q9AvBto/3jcovaQ9H3S2A
eHAkTAG3DR77l/hWdePepJk/vIPM9Qoa9aSHUdSq+WNFWvwZXeurhjxENuqM
rpD8Dr2GyUcYj8DHdBEsPLlie1eBdugKd6wiivO7MvuEKaryRuhXJ5kiL4Ay
sYse2IVF1CdNLL6BTC8SWceHCxHcKnppi0Wnj4M0QsltQhIS5N1rhBB/0v2C
Fjs4uq1ryj+9Die2XsYBs050OwMOtnZJcJR6ar+9BjEzaOT5GDLVGD8g64KW
yZDrA++ddE99B+dP/p9Uq9wUnoXKRM0t0oI3Sw+okm4I7kcOV/xu/6+BI4tq
zdpuPS3MT796HGETeEBXGX4F/fBx0nRE0hNoP0k/HglL9po3g9HQDBmuVwjV
CUnSqQRAGKNdMY5vT/Pnz1LSOp4tTBC9VzhnOE59W6hViaUuaKltLbg7Nz3z
pmJiOlBeqdaYrqy1bUegI4jr1q9LBvJZbo7LPCKJoslmPJsSkspPLW3hRqxs
c08EVY73TGUiF0MpUZcwP+M8H31CypBcbldom+wc/gywQl8jBZvzxXzYaL+5
AFAKgYbrkRZgC/61X+qN4edaDniuuRMDYGS5hkGKdVqxDw/tfNRExJQ3DzvB
ugZot4mwSASSAfys2gDG/e6Z9NlZSGG9jjXTa/MpiYxmY2VeFGsCBPQjggA2
tywLnNwzh032+f95+dKmjHjy7KSlxVok6kzQ3YjyHyfq/49wbH6eHCl4D25S
N8l0B8nqKqcRH+a77NtUE6LDRXXKaUU3nNElOR37nlWBI2NH0RiuHD++m6x/
kZ+N4zJP16Hs6SKHlu5uBYFhqUXGn5y5hOdK6Rhz+z+hhAMoI+CPPUc5SZXU
S7Gj/Ir3AxPStqcjYO5gzJr167/anXUDDSxp00j5NjVBsEu8KVfBWXShh9Gx
Jw2rsfjMaeatdgqyI86hxd+XpDeey84h2UegK5SAMpn7qdAavvfNxJNdElfr
vMqm77FAFmz6r3NHNvO/vbvbCvSg1TRR+VCzHGdKZUTs3zK1JUhnMK9y9Hc1
3wZ037riLfuUWBflGf4IfecHuAW1Tk0gUuAKsdFUsZpCuEAlJGLXZYEDo51C
qyfHHEuTNUXy/mbygmIeIZen0unwYzPRZgtddi7nTD0ZFX/bPptvDujVxkdF
lyCuQQWPtdtNVkmpBBpP8IDrPtRQSqoAG/9F9SWphODU8UmJb1s3y4G77v9S
b8REuhxiXg8ApOgdUI/Q0Jf/nuOmx0nQ687A5YW3bh2Vk2+OrpD/vCcv9bhu
eed2G14G1BQZs00r8E2RMdsmSLtkWQ/rNBAFKrhtmH2V4uUrnS6WvWixFsnH
Lqyf6K1lNx0fKBnMXC7BljI6uafMH2d5Dd/84fW5dtHNDPBo3H8/QVN7kIbZ
ASByeZCBA/UZ4yGY4oqeO01aptiPXJKmxnK64tC3NXqzODclwMTygCLGR13u
Ib70hrDPq+ccv2YZnKOjYOvRYvoJuRpzT7VtUVZaFU4jFxPKGRWKQMTwG1Yc
e8DmothWdBpTro3tuAtyXPm35fcc4SYnbbPGm0ZY/nu9JudQkpuZDE0Wd3Dc
fcz+Tx2R3FIgsDbK8p5lrlbovO3T0WxXvEXxm9oMitGsHWZJuiegVPys5+eq
pocPdX1yoNzoMJZTGT+VXjbccQFGWO7xMvrXH9+mjq+KaqP+Pe3nzIiKSLbz
Ao44ea6a79Bdd7Mfti/cNvVY8Wik3iKrYAhjJWG8FK4PaAZswRsZiMsUQO89
KnZS0czhUUutV6ll++No7/or08ShjiN9TpWX48Rtj+bl5qTA0IPcplHBMtRy
LGmscNUxDLAtzjrmMotbgJUEHaPnOs55RAdmS6A+vJYvRx7g8T+VfZ43ae4v
16qTudBckKZBvEQy77J8JUQcEIwRDryN+zeEpaOo6pkWFw39Khe1qPwa+hBK
ZZgZo4AOymwatQP0cR33+xB7wL70HAO3dwIhYJOL0JszguOa0IrtrBYi9BY+
I/T5DPyHS2/8SAwcsuDWv1SmuxzsPt2V6ymVzcsH++ldOZdNHCzDuT136n76
mdiy11FKc71LEFv+kuxvLHUfLrEc5KQjP68493yPTGNpvr3yJVlBCuLFyJ8C
9kfHG/fD+XnjK84N4w01P3tLgOZSdpVHjW9MLjlEjyqwg5KtdWc7UGf1rxH7
CKtM9d/4+ZNykWHYD+BVLmb5LXh5IhBDUd5kTjffEmc1skl627sCHW8wgaTU
PMyd3LBeIunioMI7j16+1+PJdaTnMKX3Boaet5pe6NpyVALCBrw/8NU6PZxG
qQK1XTJ04ui5qFdiG2TyDtTp+3/+jvAIfDMrwEGgMvMQEySV/eVgZ2uI1Rrr
MyTyNkxwpRi5Ho6CghhhH0zJzZOlxhrY1ttOdNIO3JiAZfBWtWFiun62qvH3
MW9pbwIQK5FcZnY03nYKAr6O9B+j4C5a4HRRiwljlpx023hrphQXO6KmHdL4
9qhb/0J6CJXWY7PM35EBoo+mRTfIkUKC100maiFES2b3/wOJsDVPoaLlMyb2
w64qpoZACtQPO+FDoFfOKwxKRei4bim5kYe8YGYhVVXjnAJYZxcLhvIeVZWq
THgn71YRpWV8KK+nZuz+8pWbgmjr9x8oVdX0YTf0XQg3b8PyWucFh9yoonB2
W5KJFy36e/6gtR7Jh/73BXtzg9chz+VMmMGwVq89Nr6Ub/BFILnbohLgnhsn
y9ojGPotde4lkgXWt5gaC5oGa+8nloOyxlz2vCnSiiaKjm6kjIQU9VOyQdH+
C25UAAuYNvwWUsy1JnfufBq6oh0pYvsvn/GtZm3YBhkPn96YlyHUp3jvivdj
8hiF1KFBJ1DhnaRt1SQM5gXL6IfXUNB9ki0iNsRrnnwIx5ckT82a9yb/NP1G
KLQSIJ43hmGw9uQaEewuWC59euf5bzO/6TM/am0tlCUGOTSqJfsER1R9HqyQ
uilsIRrOxA7LIKCWXdOqlydx/j83dNXp34CnskSJ8kzVsgrf86ECkaB1fFwW
39GdDIduBeqtGERxBIdUXa3/3L965brxHkbICE2GfoPmMnmkFYrT9P9u/Jq8
fwnXcIQw79/veQXlG3gavrS6nXm3slZpUvrTgl73H/Dt734HbLIfhMZRY9qp
Vnf/RVvOqc2IeestFFDt/aJwO1tu9mYWDuzzg0H0YBRDcLlvZ4tkRCXcrSb+
qMjTxPFLsl0uYVi9RhzVkqGr4LwwfPNLCgDnm4IGAa6KxPkl5pRVzB503usY
m2ttpzhgTz+EvU/+fEfz/QgxHLz1H0yA8yZ2lQPvqseFoEJxcX/woDkLt+zA
dHYrYZapGT3bEci7PUxcBpikau9ISv08d5t1zF+DYcWPDuYgjaKcJKl1YIe0
DGbh75N2dK8oI7cYqvhF8QD+v48+UjCWF66GxEoxTjn+nUFR2y7pGUZ9uIpc
TllLHvb70pHafEJCZ9oABlcPhE4p20rpd7EsB+r26OntBVQH7QUR9AqQz913
tFf0ecWuDGwNQn4SRJOLxspUKXXuGmw5kJP2U4qebuLshS4JysJyoCMiYB72
HJ7ZRUZMNEN6I8AOVHKcqbxhBUBes19zliPjCaiGJEHN6BKFh3KVQgjJ2t3e
CZV18qOmx6byITneCrm7D82OBzSmCPpk6p5Hs73sHnjTeKbjldTLzrnI9gDj
4h7LwqllbclBh8+oAHYN1mzQHsUa0r842v6mZmgw7liYmbUsFahQmvwT/GUB
1TWx9tYPtbhLQILiyAomkk4e2KIArPrcQRyotitSl0rnLGZuaT1FxtkI6m4A
Bc1fqmjxSPQzVuf8y9s1rw4910yK+JiiBgjcVLwLxBYMK7IrluLW719Eyr/P
XcSpPpf1//mQQclwub6zzzMt0gCxknuR50ZlR4O585Mjl8UmCHfP7zIkqfIL
8iNJES9IfwyaSW3KgVpnBSR494bMRjsidebVFQJvAwT0Tczk3y92cy1mV6KX
EBPq44x9nO1H77DNxpanImnTCXbdPv687R6XFnlRwe/VHQE1grrjzp81oKyg
JAMhKA/W6PJx5fp9ZQf0z41dVbLV1mWu5hbrw2qyTC4WegFaZdo0d9EFF/ze
mKdC7fGSfL6ZVi0c0w2dybgp5bxqHxFQmyrW54JqtDmPSznJ+sMOZjEzFpmv
4Vk9izP0KBE1JHH+5qFvj6oLg2CcUAeDIXVJ6F0eJYI+E8RwE1xR8MKvqSGy
sqGgjpjHj+T3pqHRL5r9CJnfeZyP30R65WNM4y059/3pA85dp5N/xLqckXuX
ndOfejYPaRXIGjRxbgAQkDOpJ8ictV8/LvML9Tag2ADbjlD9E1G3LkopHrKV
US5Fndr13z8F6kI6Si+0YsdBgC4vWuhdWxTENjwIa6sEKMChbWoxXDTtxNLt
f/PIaKj+7NJ/JiSGCB4d+V2uDQYdn/Dzy9GpsNqpxT6+W2h7ALZsRiJHLJtl
Iu30K20mtYCsuwCeLXMEN1cyo/cSQ7LefUmEagBva1WfkwEusTL62ZRRIf5l
LGxeNfHI4SQu2e0AT47HS3ky0aMyO0sXT6A2I3+9VrAkVGpq9oeV5yeDxOm+
3oaRMqdz17A2SmZLTdecFlNHrSUxR2aLxKgS+d5AuimAaJ7wkdihtdjQPGa1
VC2P9Wuuw/D+PH4UR+NA4vKWLnk/1GM1UNELqzG8Li8GrDekb3IlvbpJ9D4f
88jQ1j5rv1SRVlkdm8Jj6dtRSrNyo89Jkxmbg/EiQ/c7TrG14EvLx8KCrqHG
lD1173sk7k/yH1VQBCbTsLsplY9Z53NBrwAW4p/ZAgRYW4DmLVJ1k2Zlp79i
bnYdPwORaxCc9S7Q+KFVGbIbdhcw3fLdboIOqGZWxzBHg6i3w/+ryBft5CBr
Ie3c8IO+aHJ42dSp3G58HfG79MkS12wvMOx3cA1LjtN5C61Jj2wo9Czf/hjv
w0nUzyYO6nk31XQT+2uQL6cT92li08yr39FVHUsY6Yx8NlU1wC+VLNziff8F
91zy2WUEi4dRoputZ++Xcpnzf7BzGuyx1H08F3JTqvR5LzrAWwpPrEb2iG9I
IieD0S7VV6BXv3XJmU+UuVgYNBYlWB8uNlazJSULgdur0vFfdhubNxALJ8um
WSbu4C1eEuBO2u8GnrZ5vX288cZlajXNr6iaQ3qw8SulUmqg9iz0p1CqatrB
bxB51A4EKYm057HrumDlMvBT05UtgCU97vqaFIF8pqpzxGzfEsx67LUdW/dB
/oqmOoOwU7mbwS51Y9ekzHLc3pJa9/AdmFxAAbTEatajgOQwi4KCMAGXvgVg
k4T7UvPBN1c7T4pL8y1L7ov/kU2KJCD2l6DTGKpXY8shge0n6+nxA0SHsSl/
XeefZk5gPg0h1YfQdP6y36dVGadVuEHCU0rtA620BkOIAhhFSVKu0dSG02Qd
XPGqxe0sF1AnTjbxANw/aEap4jmz11z9Okk68d5Pp4/qcyAjSfq5ZhRgfWdj
GjAP/Qz4gyuwSRQH5z3e0tNLYQaM2X+XHHFT5vvrVvekLV7o/BN+KGqIDdSv
gKvmJ4TfQiyVrERsmSxvQ2NFrk2agLzDQT9RC0CRN1OP0zmzPgzDE7Qsbsqo
nfqVsY2WDBZCkz3l2ynauI0dU5U8sMo1+lIyGKnrlf8cPs7zuRcVZzj/jd7y
Q8MDlx2PxaoNn0612RzQVrxjymrrc2OPbA8zZiYP1ZSMAbr7HRlp4tsWjiAR
7ctr+ZG7Bl3NM7rIWITtkWIx8EQpKeybMjgVbwF3XoZ+l2VZtwH2I/Fd6NBl
O2Q97ZNq8gmRyAoYfbY+yg1H3zzIpWkc0fzfhI7vyARgLttiYuP5p0dXBqw+
3OBTxOnB7CUqhRNAcy5PfUz9B7XaJqBqFvor8EJe58/tgelvFvGxCwowTplL
rx3uTmbX470j3BgHqMsVeC8O5Ez0ynYx0F5UC6fMd0kSHSbcOspr18UME9/h
vcYShy915S0g8HJbQI6GUfBcRlv9RWCbOu5XseGsmyPC3bTfkzKUIOnMu/6j
QyefUYzZpXhyoUUk4lyW7NS2+8XaNk8V1ZaZbW3vhQrh21FMnrK4V1yxF8NN
ZD6+KEfZPbNiYI6xl8jVIpkHUvGJwu7h1Zr6KtiDkaCfYhe3XFiKPCn4Nqtx
AHEPbuQpkZTq3WwlsSfowbW5WCjcO00aH3pOi2DvcrsjrYcNyVGJIJ6jd7Bg
hxGqryh/jiO0bUIu1JoSRFOqwhBJtP+3iFEp2SPg690k+G/aOvvcul86rBSG
bACsr+YzFvzXkf5T6COW5SsSQva29czWrveKB632b2XnqAjrStOXeVsoGqa8
ke1q0CRLJ3pD4Um3fl27xabiQS3ouon2iXLWvP/WaVaHO36F2KVZ17TZ0TQg
+kKv6BH59fA5S5pafXax8mAmVVc4RPFw/lhS5GYcJeOzdbQio5aTLP6xnr7r
DogyWCnCSdrHTuDPpyGWvgsXksYa+bu5Mu9WfJ9zyKJIHWZuNaa2SbemVe7r
IwOaKWrNRbKYuGQpWbJsiBnkKg0ZJ5qVwPmPR/fpuUDeXvQVqtBVU5CpMPO5
MmR/8dbF4qpAMspmKREutP1q+qO6x36pZnsw1PGFtuzyExreCbOjtjP7OOZn
xDiaPhdMITCrJctr9gSIjGWbg/bokT7vKXaEPti8G7JJnkUVzK2qeA4yOiHX
Teb47JQaUO7uChksJHA+tZrRpzVHXASJeNZMhjlouBupolljOXIRAsgGz9MU
Sic/JuH52nH5EnI1m9TwI8B5oHsmPOVBhfHsMIGz3D6xj+OoP3pe27JmecV7
kW2Z2HopGIMQRrSLcrlOaRuR6QzfRkLfx86zQgIeheDV8V4EKAvA+4IZG0Gs
SEJacNFBRZXjSfVrCyw1xuWuRNEWfkHSpOPLMnIdKv9ghIKQheTPL8kF+ae8
xl9sMyqY6Rx+eLIq/FrKKJ6BLyf3pKJj69SWUFJ6jCONuIkml3vd8pp1hyQi
1J6aHr+9dUc8iIvy/caoyYowBNTqbKXaKzhzWC5hY6eT2u7ycEf0YRrlpCW4
sRF4Pn8dHiZJuR8CAonCK+NylAuQRF6is7ioQyoT0K68OGw3KTVNyipJ7vvE
VeAhT5+wZJR/oU0zuezugfHC0CzjcjHxJ4M7PzYAEntG/n/U/efDHR34vByt
iJW1KO06vXad7DflYVy/p7ljeB1miCiRtEncilx+2hQqLsKwuL6sHrodbAuW
rIvgEx2EBMYHpuacjbtLU2OOmrEECVBHmNKX7edMFyycyGE2e6HRcKzY7RrW
7mRRUjPu0akHCXFEd2eNfqfQdQ8+/jWEz49WsJXEM//Vw51kqBperktOdxC5
TYYUFky2UUDQklyuZI/p5NT6IKCUhhA2RmfK4U9MdDZBBF9J6HJWa1tgBoIa
vle9lWPMlekURW1kKenwqWUSleNCRYf2yktzpGCVoPbZ2sXQHMlXA0IR72lm
AokQ1kBrWtlvr24liVNg8SXePsBz6Tts9xYb9UdmrB9I6gAqKdefsrTGNXF5
PsQprztyDIGQTEUtk9cz2ARR0wSR61UFib1H0ZYO4aVFiEBwoZyZS/ApccHE
uHnMRo5KWTzIHIY+up6vxG1wwuUg2V+ILxy4yUwIPuUXzlE7Wc65zwA0vNDq
ollsV4JFqSOldw4FXaKqNWr4kJYS5G03VvRs63Ss1fNZ4O66Q36ssdiaf1rZ
RiY2yXgu1Ic9U8rv2agMkSGHachhXlnEivZZ/g8yPzAg5TXUzEek7IdnPKYa
8LXiCoi24QO6bl4LjYcMCVJhKUpEf84G1TFhniSNMRDP0Bp6l5XWJncDDtS7
/3qe0tw4ssWe54m6NINcCXaYAoCWBQglvz+PASNBRAkozYhp737L6zxhjs9b
6wBML4rFhMCG2ZPUyiLD/HKyMUJ7msxo4hMXbQX9Wp3LzRlsnT4xZVZFLQb2
t8C31aNl/exyuWxIdy98+sGifCCCbUyiZhZlSeEVn0j6W43FotU5LYaWRjyr
NEHGUzd1hsGRjIrOoIrX25OrcFWjG7Bda2CCzTgG1eJZY1GhNW557wr/yPaA
4LYBhSA9Ol4cc6FTu6p7TpwJUCvQTSlBC9ec5hv22fwuTqhTcKLFTL9e/C0v
yGJ8zrhvgZMit47gLGpGTcrzwgo/tcuwsCAuIrpIPEd83MgoSDBhk2M72P2n
l4TT+M4lg6vB+Aneb33SqX0sE0ucRHTBZCqWr/8TSfSGHyaDScm+TyNdOHwB
mpbm6w1JjONuVuw/esBsAPvlrK5YNs64Pw/RnHE+7JI+3p7jhm5Fb6vzAnMc
GnwUrUno0ox40x7nvCJdHIRgmrpGBP6Qtd0ZNrT2rXEyZLm3RlU5oYixYAx2
/LpOgbuvqjZlMwTiyJdqeUAFoRF3iu3LQOsPVrBBOa+7F/KdQFvL5/t5LsH4
ZU6Wxz9/KVrggRpFbBwEqlkYiVxLgtPbcuUQmVCI/iEQK0Twn73Oz/gQFh1q
rSqbsg+75PBiyA6WfYRmOX5MpT+py4LVDQafRMtHscRG1o2rtZ0QSgKZkABF
lFbKHmJnkY3cMFgIA92ULwg41CuoTVPKQl5ZBlTA+AjXTo7wLPGbKA/ap9uk
E/3OGATM9Dc2OFOFHx7wN0CSOOgTzL+4zYdj1l3z57K0nrZta6crsMafn6Hc
dI8vitgPkappE3LfUV50hoTrFwD4c1fPQaonYYEzyJDEdIEFs9bF3oqC8Svr
EqVpo3kFgkKJLUqDm/fx7AhKWNgE6aEcs/I+DVYvCW81F2f2Im0+mS4lL7m6
GcfEk+ieq/jvB2jiXFBUMQG3edyf3JHUmoX5TWbXUPpzDKcOUyYkg5OQpzBi
0P2r1gev+tZrfHlfVd/cUwhRO7h5IP8lAuQjclUDDSC93DJ+/Pk4XKnWmXii
X5SdIdtV+UPLA6IxoYNgxAGiBhn76WDr5v3UZbnUEMUSD9PSbNiD27SfbKUE
UAoe9nrC6SW3rIUy0sOKCh1zi1KD+IffMTwZHQr5lh9/taIm1Pt81eoZvEbo
5eTZqoQVpu9PXvKJ2jZyGD8UWayJyC+QJU51p7jTLcOk/9/zDosZ5aC+GhEj
qbTQyj9VhaoCmg/7lByyhPA12z6TMpg1y9NqIWWYleKU+PuR7h6a86noUCnE
qV8ebDIENmihNsb3vHT+a8obv7kM/G7DU8LPGiJsbtvnZWubRStNQBZuHRXg
3xbwSrK49fiSW2FISob8+Ydhrqqwyjdt5gi/Ryj6zL1nvkkapw6MvC6eG9PM
kJzEoVFY4RNFgjl69gpVhqXw91zgmMSI6g0QxS/4jReq6LKeIM/IShtlWYkq
7Z/EudhPNh6qq622L4naHyG2BkLNrIUkApZayRdWME7G63y5wmzo2px4Sfy5
gd1dCYNYAmQSwptbU1i6O3hKDkJVKRnkd/AIaoyJjWCzEnyaQJ3rFfStQ6tK
yR5BvISL6kl3pi2n3zDfxGJ4IFiBMocVeehdQMqBJ7PD2tU5FsrE96nCcP31
5wrG2pytA4SPZ6ADv4VysqLU9qguo44XzzJkt24urFqIOq7ThsCvQPIdeoaU
vD2Nop50UKEJ2XlttfxJyuLlByww1NbE3XAhh6fpwi3DolAxQrJ6WTyYVhQ9
mFlbI18V1ChQuSYdGNHjGQhIp6BV1+vOtzGqU93/F/plXcMBNrjIGb0vqO22
tJJkpFsNItmIR/S2uII1AUdZ/chRZB++XTpShdFoQTlqDnJlCO/dqO3YjILk
ZYrNPT5k92xhs2IGVavyV2+r0ySJsxfWuQaUZ127IeO2leiHBx3A96Wg3MK/
lk6YCKC3AFMhgCNN2HWyIc0RcjG07mSiu14dEJv4AIvzusoYYvPC7DqUPRB+
c41RC5DM40+hYmI6nXWT1gJFfN57QQ4HuOby2HCqi7IDAf/VEmdTerN0pF8Z
s55Cudaz6FQOEmud2Y2WIomyLdEf2L/nRoodPxF829mtFJm/ttwx7ys1o04N
Bf/LDHYaicofZiDAP6lJeBSIy4NRxX2G3c7sXgaQXthj4EzibBX2NTAJnji3
7yEMf4R+0QcmTvCk+oLKDPCXy5qFkCzsPDeNT6idWC7HEg3nQAVR+coUGlH9
Y5UgWy16tKLP4v6AsqhrnhaorTmSI6Sfk1eFKfNMyxh9hE5f/3D4vrCvgK1Z
nGh5Qdnusad4oVriD1neaDmB9c20IXEdbsf1u107CQF2QZ5/dqZLCJzRRsdg
CIYuRgcQZmjVdD6enuu/3sv5KqUQIKmqLxTszI5t4Kj9ytd24UsCykMORN0j
QprAADf3+BES2wiP0OUShnLbPRAs7Zavo4U3mSdxN2qtNTb5QnhxZVmxCNZc
lBNT98uQKyhZhV4luAWvYy1lzGV5xI8mn/sU59hSTSAAMoWyWrWhwdumA8R1
7rmwfK69g15YJYyEwH2oZVT8EkkaaTWXSKwwACHhVejjt4f52XcqpUVAxmSj
7kHIKIg4Jn+pNHv6IcRjQRhh/3SuRvcoTejBkMG//YqBZTpvDQ5QgdUCnJw2
Zxv5R/txIGYyqYte1kx1LvLODmovINAEQHqF74s/Bi0zsxbwjDz/X9IbbFQW
n55ICvyVpps2M9Y+2TRdIq9JqAfEF4xQJlS6dc9qwUGfbNAYurahWCakt7K7
ZM5OkaWb7KCVbtE1QX0Og0si+40qib1YdyiTFpufWMpmkELsR86DagVvH0ne
IWEA6Op8tpr+NZf2lshi067z1f4lG/O31x1joi+cP3To8n+a6GFZquffL/dA
6SlI0kNZ3YU/CXqF4m+D6+y9YYz2H4gL2Fl9EsmBf+fvtCchbc8hkymMoJI8
N+wckSMql+Lfvkk3T9URlF7lgAMddLCoy+G7RC3ZOZcpugMiMYj2UudhCOqW
Nm7uUPQjAvNQ4GlxKl3zZ68K1XajJwKJs9fivTHvuv+O9lZJjG5PYO/4LqNL
HY4SYdTawn7Y4BcLHAYA+lM6FgRWk+z5KpjH66VDyUpMumg6geERaxNpBSvJ
HH+CYdRCj1aoICtNv7ylTy0uW/MK04UiP9uXexWKII0cJzPE4ABT6N7ft6Ec
XBfdndUDhlvSmsP8a74ITehbAwx0vnbGT0hcvB43UJ3Dt+ehOgJaMVkNkqoB
WmkYQrxu2oUgidozrMnXPH8PeeFEIdvHRDIJLKunh0SbJG+yRXyFG1g/wwyG
V6ewXj+6oOMjMKb8fDN3FIVLqVltGWyE5C9gkzatEhK5opVDcsBtqPBGe5Y2
SSfgHzF1/inVWIK756+wsZq/qXpTLEz2aitEMwJ9e6fc9FY8ZvwlNRR1le9o
XGh6d8umIBxHYdS98epOz67+CsMA4FqWHXx3RkZMaFpzPEQPGd19mZaOq86x
CZZ2r04SZCjaIJHQKD/VGpg7pUvhkl3Io+d12yDhKF7zVbFRq0ZbzHKTzCTU
wPEZxKANAAgEK1Kwgee1/JDvtoYJXYUA9vwYKcIFBlpwumF6f1XfA6zHZA6t
3Ahl+KLfny2MLmmNNT86jAR6m7QJEILMG58bgoS6q+P2RcT0maxIGieNANfA
X3oi2KB+MGu3MsHlYv1GOm69DZjqvWhTQLdMXDb99mMCIunPECD0VVO/8Pvj
MfuQkA4JOg0hHYIxi+T0ktQ99quCtK3+vMTx//eA4LwefbRTSagX2FzhzMvu
tQ3UmgrGawWvz+AO7NUHagugnEbD2gTSzSNXyQSgDQT2EIkcAAgUKv8GhHTX
yJ3/M09e61uxxgQstruo6tCBb0quJytEaV9t83Blw+ivTevjgjHwJAhnBJBu
Yg0gKGsF0C/ZtxE0MfQCEFRSITCa9kuit8QETmHbk+nblzmDxNyd7sZh1jZY
3XDPC8Gsuqe6yp15uwt7/zxBKUhie8oM02B2kU6dp8SmDKnj7eVAAvtm4HFE
zMNvUYZIYsVU+oQmrUFWu+nU2Uis94ZLSu/xDatE4+hYez/ZlA7Ka7IKBK0i
pXAolzRDNognBnIGrJZU5xpv7ypq0t44LsHLoIWObFCpS188Rl4O/ANF0b94
WQldhWromjak8P3iOSjL94+v9ocOPWzBRQcPBw7oybhPrGxacovwfxRnRSXw
hlZLVFIoEVfg1o/JZ8OlJqzAZ3QQHf6nLFpzGxCET46uKGL7XcV6aTozGkAg
CFs5TigNFtF3ft978YE39pqewTsqApdYUUJR630wmvjxc2Uw5BTk0XQZ6SCs
AJ/xu5fopMVmvAxCav2hHwpgrsn9R8tzci7u0HpmQScEcyo19FrVE9QLmehR
KsP7JO+cE/ktXCJ4VKMBQRUpmjrTBRkabK+RD80OMPHfigXpOeeFfKjMOugb
hwPI+Xbaax9z5KC3LvQyuCg7MCOiQjPBE6O6N6Kdadn6T1e0Qgkvsuy+hdRa
cZ2B/ePqxrT5+xEBTX9EENAbS2qbSlGOVqBRDDs6hQszuQO8JMsomizNbEvU
DfR+uzLx0k1BtnJtwtl/I3QXXTsuR1Y7FPNV3jumnrAZP9aGtxT8UbwSLQbY
GCeVXaryqy7C1etWmBjaWGCOd2Fwukjsi9kIYVos0kEFMUT/QnQ7TJEn3JoU
UYzFrMBIomjub+jUBBJV5SR93EdzUPMl+yIQ+wdXrX8pOy5LMf6KxaphY6Ww
LydT7l9jOtM+f48zqBhDiMJS7A6DqWOAgsFWLdAK1I1wNHCVoqGquEd2eGPV
lAFEdU0sPz8yf+p1Yi+3d4KziE/1VqBQ4Bavbv2ZJn4vXCsBvU+FAEyWfhvO
xbDZGRgARKOvuW1ZZ/xc45gxV88AmadHGwQR7VFyUpfIhiE/ETbT3t5dxMVt
cjz4Tdn5YamhefXTZN8godv9IoQdL9D+kJfEaOXrWwTw6ghuMxxpszoVoIDO
ZXbavkqOL18lh0hnQVZuwci349tH4c+xifaJjBRY/GixyvyAfpTUu1AOA5ZI
5FT9zKeYHgYAokkO4kRim/EjU3SQKSJZTHMYAsRAdXaxz4oou7U7ukjaST/r
oXpZcJXJ33jM3EM3KmeB41aVv2VoDSOCQ2R637FaK9ZSEhDpuNVwzldZxQNa
MrNVyemsFHNpAHIVFwf2R1ZkCzkV1KGWeDVkdIEMBtjhIgY9ecbRxKBoUH/+
1gCv4PjT+QY5LaC7STbiVBx4Zm6ijKW2mTqaP6x914lxIBV8+pL4tNA4mrmj
IKtAjcSCAqKHDqAy8KEgSLY3uz04zJCaIEZNT6H3SYUw5xpGjfyOo7BCpc1z
IS3tHkfbDks/Vh1/jlXAXd4m9BmIdnz6CZNbbB29XqHGHbBRGDtDGoOWK4rW
qjpor1ik/3NZodCu2L6f8j5kqzRDtEx0MulY30Gw55H0q44vMve/5r5WAnJ2
6WPGPWu809gmyN3mLH1d8HL8E5Az45hw4j2MyVoq+3ManI8tIDR035dXEpcn
jUkyMgSEA7oA28E6jEOMUK/cNaThKetO5zwlKsgiGibgC8omErTLbRi2rnjS
1HwGr7j3Ry7cOkhAOnlkNBprtQBbIOfSFPuTyVpDBUMA7n6puEAhoGpp4nE9
9SHG/stgZp6gx+uncUfZmASj2cyYB3ivVHmVesWmN+dIQsEI7H3BuReTmXJt
lU52agKYeHQDqP/UZ/vXzUN10c2OGTUAHhnkLPMJ/06ZlQkqvV3GjI/7EdYs
Tuen9bYXZCxswpBFDtwCL6AoVCNP2N0AmPl7LnqtG2efpMeGKdNmNgB3gkBQ
qf+YFFld4sVP5LMvUJ2tUw6p2RD4HJL/GTaaUGjc+JIaWHO+1vEoDLk20p7H
q9DsQJzydtbmrriDcXlruUkSAFMp28YgyZr9aCAnmortF5W/jUxVqxSsVoTj
BqVkirnFVn68/tUkEWSpnjcdTHy4UcKqlGRHcl0wnh0GYfZ3rqldTcNqa34e
3O+XoYcAdWAEANbJGaiZamWNfE6w03R4uvPG+OB1BPuHy90vDVCVVjKhjvcd
tGPdklUnpfvfgmCxJrcG8unO3MmbKMjHnnmF9CvlL+rokvT/ZfowX8bHQ1df
HmfbNmVTnY0x0EP5irxKY/cj0Jp+7lRZa6wScpiqSY4CdjiJSKJgP+DN+tVJ
AUJsbMXNNtUkw4Fg5B38inUZk0C67BoSjZ70FsPj3Su6/gxtrIMe6XjEQwiB
A1AZldAhxjXxHCH4vfrbbWKnbKOp3+8qqtoYRLtgasSlPOyqVRvl6Zvc+MDV
/ZN545DaRCBCNFb57sJsdIztKT1KE3qfZ2WphFFWm2ExC6Q4ZvvPv9l3wRRc
DQkaKBBoDgBlV4dLCbk75KMKek88uIzpjKA2hSmP9M+cn4ou9XruSDZ57jWT
//M9N1lSRKPcZCzIwPpO8BWgxnj4fKSqIKDYe9OF64fLbgNaYAeWIBDM010l
vYwYMT9HYxHe6V010XUiXdn0/hIHoyhgfT/EQ/XnGmrY46M44PAdTu3il1AN
Xowjyi/RVLHLTk0V8q7LS0k0pg66Q2PXmgsEy8fgSZqk68oXwt7PzAaJNvh/
D7uJ6YQ9bKG7z/rxG5ZryPDjVyG4ygCjA1xBdqwHj+lQvOINVp8YbyJfk4HC
DgO7SJC0XvRdnUtp/2CfSrJIMqsvTdioaMyDeqwUDN/80T/0jwNQa1C7sKTv
6Nm0GOysW4D+o0e1Xj0lKpDG5rmEX9Ij7OJOlaNLWrQm7sE6DA2k6m7klCD9
6EWeOo1vBspBSJoD/sxxeKQiteL5qGXzDkpp9JdT0MlXjJ/wbBfshqmJ9Gsc
/nRtIfAAspRC7F8YtA5+YPn0e6v5NPIQC8VeLiiRvu3QImyrSXRe538qEz6M
FBFwZ8wAAkcnWg67MQUeuABpr+m5O6Xw+oHLWDaDqYDICIMtQOyV9CRxOWT9
8ogU5M/7BhXBUKPKsYSummBcnIbqxfqlP8aKY66sI6hKWcDPg7qadLMJD0a1
iMBqnCpbSKPRkEyY28Iu2s+U0GUDBV+osFNSoSXqibplNJm7AH9dsyR5XxNP
yufG2Ibu497UlsuWi9kcIlcRUGPRQ1Q9RIkpNmizUXxexH7AreOYukBqHJAb
z5ks0ORU4HXo0SpMP95lXkkDoyUDoAbIoqWAw1e5ZBKa+cKbWYATnjI/caW7
cYapm0w/ML/pNXLXyUy8G4Hzqa4UhA5mcAD6hLQVyDdN9DQ+TNnYQco0SilL
nWCD9kYEXpO64otFIJPtlIKFyYKF0/NaKRnr9vET5GhFvCxJgOeYLvwHKBvZ
ojDSqIm6J2d29+cyEeS2+Qi7dVYfiYVJnqg/uBmDP8i9EkzWTQRDo5a2RArz
gywj0G8r0Z6o3dTq7xjiyMjRBBGHHmBhQQQ5PFyag7bRc6w/3aAsrW8PRYYx
/EW98RacE79JQxzkPX30KjPY3eZj9kBxoY71LWt2KOC8hplghAzcd1faEyO5
IGnSZ/9km+YQ0+Hvj8gVEw/D8KGnYRtRcbPvteZlO0wrLXMpe0OeD8i5JhWh
EcIiAbC6qMV7wpvhJZ4POmm2cEHZj7Qx44Hqfszn6mrkGLU8AV01Qpz1F0p1
bKraiqkefPx90Tk9l7Xj1oakWM4VePViX+NaDOwCEvJ18YUIohK736hl9P41
F5myM633taj0sBQ1i3YNTbfGEzqczlVDU/YacqmTa/+VQKPXbf9VPkacJEwy
rMcA3mdcY3CeR1OsPzfzkTlf2aNxe/sK/Ww4s3vzoedcTP/SqjPo2eVwpuVr
LASkOdNc/P/Ktdk/x/+aoNufVmFtP++7DuuqpdocaOJvqzU78Uo5W0MuwL1i
mY1Di/E6F6FCGyfnZGTfY1lX3nFErhC17u0YQ4yAlMszajdGJXwpcyh+AKpa
nWXxt/xs5lYFBq/rbSCku2h/UC9N6/ZJGiGpzUZlmbc/FfeU76A4sY3S4oVH
PQdjDd0wyRcdmkhdFZiyMnHTDloAICjMMs7cO6vIOf77qtdqFq2YGgsuNGtl
8N1yLoIArSzNrO5R+PiilxzPWZw1AyCjgEZ3/eutPQp8rH3TyP9TTU7ICuLq
key33wsosVd0vESsIONBp7fxOSXnh71gLQDk4d529WOwOgK1EYgW2tLNuuhm
NhSup1KU42Rl9p1aSUK441hROu7CFoPHRyHcZ0u4KYT4v4brHHxpk6RFarES
jY6Txsf2ETzH3+tJ7oN9Ts1y7kWAgPq6X8lFynYxI4/y1vAw53G+VXW8mF04
VdEqVriRyy7qGsheqlMglTDz3kyHEMQaKx4IwIorX7QN1FZrUSULh0yEXFxv
jKy+HPVym4niCGUWbCJYjzqayt2glwqF60ISHK46YEQXxearQNW+u+B83OXU
sj+PspAaHMT3Yz58BS82+O4GypBDAeWVfCtalrNMln9VCULB9sB1z1KoJwOK
WZ5iLXg/a1Q0oKbB2/kdl6tK1Mbbl1OkiD2bSB3SbIb9xCfJeWp5yxZur/rq
WIOyvSZOSixooUnXgXiBm0M5Bku2xfxw2alh2+3RVDPQt8Kdf/hM71t6Q/v5
jpj6MNqxye5G3/Hv3I8RLmD0dWIiSTvYaI/aQkK/3Woe9bCMzLipX4LT1F7E
I/G2Ll5wQZegG+I+/bYnfOkT62AFoCKSZCil3fJqiwDtUqcciDdVvvGekp2B
DGgS8MDzqxECiGdQyljbA1pX5IzLRzR0JOoLlwoRTMqf34fyvQwpXTjT3EqT
gFhsGJDay3eSrzt+z2tjeJI5Encxt0pnvpm3KgEVZ+hfKypB29o6Ry9NeV9e
j8Ciy5FwfA9X+y9lzA4ikqPbCS7PvTqtPTAXjZtRouxwB4o6o07bKrO9BYIl
l5qCWHisHm9h1X0WP8EwpR+2DbIv1ZWfivCb30qk5IWs9NlaSl9FHGhAGcaf
fDHJuucx372YdPe9WfuvawbhahxkmMus8kBaBm1mmJF0rowqppZyAIkXo+hs
fc8LHA4wWDn/r3Q5hadSDGAMU626X5R3pORBcZ+SUWP9j0y0R5LgzGBdnAA4
KpUjKVLk4gRoBtsE6XgdCP9VdAFB1OywVaH1laMGVrU/QdIsvekqPLzR/5Xz
+uiW4Ux+MFmFMUy0EzJGMAvk7QnwNgM2ES90DiktFV/bsC+ezvFikJa7hpRp
fZrm6q6dsqf1ba6SpqzBP9e30t7yFgD+0X+Kr/L0SCfH23ohQW5WLqZb95pK
5Q7RCHi3Z81HwHH/kbk+QP2m64EIjrs9I/s2Nb9HPlRzJpdjbef1MU6tP5GX
2YplI6/jI6fC2aIfYQVzpIZjXiMA9fh8cto7w7F2323VV4zm8Z/wD0R9ZwEK
LRea46nZOArLSYUuvdI8Ku2LwekYx/51t8H94tIQWgCS5UGOEgX4CaBsfklR
S6ovT9u4lZ/4h4kufS88sBONB5wZVSgKxTKF48wI0hBQra7g2/mFx95h7KYq
ldGjoKweA20czsfOWyE7o0/3NEaTq3tMZSdTUITsH/k1OufVUyDzYdz2bLA7
VBk92DBA5ffQaFFQr0Lvg/Mb0sx/5PyUPpOMLKlM/rjVKvxRHvMtcYPwJY9A
IDnXbzR4dKk+3saHYn90CqZ2stQaj+jniQsJQFB675iaDIgx3B5JNfrPRjuM
ydsUfIT03wFo+pKfZEHrqxMl/xNRLiq6hd9w0JGVvy1Z1sXdIUxPY9n9QkAX
LlB/aoI3kHSj0NVxXYZcJ7C+eC/0CNmsPfqfyFvCtNTC4X5BZuekaJ72/qbO
yZpVhQ0bSlkDb8pU7oVllQUKgeOn4vJTd7cmzmAsqdKclnmn/iuAt4qm4Fu8
Ozq0k5dGYLWI0/Kzaj9/yPoJtOJeVf3lcZ1QI+Lx1zhSNE4K4HIAXI5WKST/
zA1f7clYtVnw7WOnV037XoIUG+DSwS8Z33XkD2afaDOaHuzcVTHNlM9QPFb8
3MtOVYu2d5WMwdwzSmbc35RXojY4olW1dTBBzVuVNLmVtwGIC2yd1q7Mu1fg
CIpVFMclWo5yCvRD7u0WmANBVfvG75MN3pkiAtDJMn3htKMdu4QqpI6FOroQ
tmoh27eNDo6NrZXn2VvZwpZK8knUGQo1qdqw5msVw4B0WyOXLZ4d2JIeRPVh
q1vb+whTs6PSGjHmxceoaPANsC0/Gr+xcvOeAY+fscUEzhnqfEqgER38RDbI
rzOtqwQuAiTDBseIGu1oh6APV0aW39kUjxOPPYdy+8fm7xD9WSODDA5cWVPN
queXyjkKztjxPChwecev/XQZx3b8CVgHG6spCsGwNGXAqISrER4Up7AIQE1n
hxW3Ol222iI+JAmkmk8AhlT7TVPzevR3Ey9PVbq9iswOk1wjCTw7VbjOeNsZ
Ol5nMPJIBgHhLvtkKVxiIFvvKNVbBGMBmmJiLH5I00OCBNoKT08oiJtMfHFE
lLCFWlfcEeIvwd9VbKue0z8Eejb4n8A0QSbNfvv2iS0PZedClLUN+XNehm85
SCfePXKRYSg/stR/yNVV5NTKxZf7s5COXBFZQ/9QdBtHS3robN/KCwEauywu
HjXGNAGJW4LutCuJgPXouP+qHL6jMcEzDo8lM/EbwQg79++gI/29fwBI2ahX
hDZKVsizHnUPCPa2biD+l77xbgoNe37MOGBFEukS7jZUAvrxsjWxcxsR0tbu
lP2omyyeAbIQonq/7gftgPV1SRyilAF5ROlnTKPlPeXr+3iD5fvZxAL2PM73
WDqE/mzeP/g6hmK4Si+An8lhG8UXpWHeFsvkQPay2wGMjmsD5XGTPtJ9Yzwi
Jf0PI7DHUzcsJuyPI+/rV5lJdqNhjCRfECpwuIbRFD1oG/Iwsz+7ExHre8uF
1ZGmwPtQyu8Xpd3QuXj7GNs45EqbFLSyRdgmCgXX+9rTk9Y/IPzCoqDnO2RB
Hr3Ebd0fgprSdly/dR7/+X+0Ym/+412GmYeobF46WwSHBvxgR64pWT8+VVdr
otcWvjbVh4CcbQZ0Bw4gGQAjHl3yWFlqsXMQpNEonCr+XqKAQHmJQj0Vdv1q
gjstmvJqVM+4zX7HXNn55l6YsdEZDpzcaWA8R4EVG02DsbUGW4c6uSW9P94Y
nUA/PICDdcOZmNIXsDBIp4M6qyOQ8WssJs57asap60mZGGw65ShVYAURQswE
oHDeL50GAJmA8b4u8KgdWeBULBp3Aw9Orw6D4yTfdxcx5hJGz9TobM00OFFL
pWGwtxndwsCn/iiSGaHfeiloL+/VYsQ266fxKatoRAadh/QQoiHEuxC5M3Lh
ypyxkK2cMUVFmykw7ObVAVQhrOD4k3vqGCbweOj1YHwDVjr9cVONB82yJhwm
wFkcpd+CZ14k6l+5F3wamhuVYZcztLtz0n+vgI2/2NEft8kGHRzaUNVt785R
fsN+6FakZbbEkXR/7ar1rWLotImuOFvFLF5Ftwi3qOLw5RB0Ps4d6EfQTnAc
Odvvl4Shja7HllhJ2/e+sJ0JMO03hPLVJOVuntunqWrhq/2ciq+xXbn2npVu
3cw/ZEQJSO/XpHi6sl8oDYg8twZMPa7424GVXI1Hz6te7ohUXvHAyC5Pc7EI
JTS/XeYa6vVMna3dOnfGMJ+c3FL/4ld+fKe9WI7e69Pnq81kI7eAoGs0eaEV
9CzgGfpTl6bnjqbPVnOYIPCpuFu60gVussi06e6M9LKY9e0t452G2rfq1QFZ
bKDeNe8UHjuMIsJ68AMCUtEqQVjbZIxpLQUFhNQFfkmooj5WtWne7C7GguHj
NfvQkNuFgNqQ6sFl+/jehQgHNQhZPCdsIhI8CJVVVMp4R6j04f7kM0O32oK7
J+7Kcs8kP/prlSeLct/U3Fg9jpLmzddJQ3RlukyRta2HCqjN8/05I+7d2JIt
PqNIOZ7FbJAXOaOP5J9S53Z1qA8raHEHVfXaRjSrHEyAm5hLdwsozfZnPWBv
zMhTruOOf2a8Iy9otajMeALqVfEVSYc1dk8tjh1zzEtsnmyHeqwY0IDJO7rM
t2lSI6l/cTm+RRevOh+Ta9u8ZFdHDF1Np4jJLRfXYZaG4vRdvkf+daIszXO5
dd9g32B/BeUCWNckn/ZzWNdJrcZWLIrB7OTQ3t2sgdrVIFgDTBCdbT3OtzpX
7oltEs6bCWcGJIy+MOpm8u65AQWtZlo62Cgl/d6jkNy0W2gcKGa65wROOzm4
nKTwdgrF7TOrwtcpyJZuJ1XJF9hOuAv30KAGR0I7K9VE+bgAf3OWsxYBH//N
7eeKFt/zTMWdmEA3hUqxNOLlqKVRkX8pKLcTj+4HHqTjbMJwTXuFuImTLF0F
hCzByQxBco4DZJdQrdS5DzekcPGOBuVXfPUGicnqkqqDj3nERhsyqyBTEHiO
inzMGfmEpxsoHLQggT/xh4Pv3sI4x3tqHct03B88rwt05na9rr16E3ZQVRaU
2t0CbLn26nQfGaRevvdOpjJo+zXPs/V+/xDSqVTVLsTQuLxgYTIlC9Lr2qJR
R0z2n515Rmn7mewhrfobc6CI1yU3eZnE2sluUzJuZKqFla2ule/lUQGZgu5k
GXZhsdlHSGswlNiFvOqteVhqFhmAgzpnxNxTavxug0rza4Jgp330BFXVQnYE
3vmQ0B0jYB76Uq7k/eseY0sQWHEsaacs9fsHoLlC3CHcf4JNY4DvHl5nI2Sc
5UYUzsu9tl6WjsrJ0Z9/JcQ5QYGjO1nF7eEsBAWyMhR1+LbVAdm4dGaunfvB
pjdVJ3sBcI/OoUsmJAP8FXa1k2qiGncYoac9SpzMOzuclt8mo+w/3ydGNRIw
SUHgZPnkxkMAiNSr4y+RxWhcqTBOwA6ZihiBVFUF7VoaWnrSQ3NIOA74m3wi
I5sVItHOUdr27LN6RAqKirRGEZrgFGODOpQlC2ysUuYXiBziUVdUudX+6IYZ
9sBsJ9+TBQKSUWSjHzn64D8E0hUQDCfZHjpVbxMm2odCdwXfYqLwCLniislP
XS+3Pz0DS5GyyVRwSHumOC8fORm7efKEsieo6dok19/SsMjha4Wn0MHscQHk
wk8JhsWdizLNIgHcOayS5ri7uALUgk+yQN35tqLtITT1zThA/afjN1mQAYC+
vbpMw0L8K//ihakH1MaHwF4kmS0cB7t9L9/2Wb9+VNPi7MgdvfBvX5XsoCuR
FSd502q+eFYn4jZV72ul11tkYyqBozrra1jD6EB3w0rOpTuiAB7alMSUxb20
I9cagrFxIHFcRuRbnojtsIN7YyaMVxgPgXM9eNMhaOKwPc8r4YhE31H5Nqld
E3Z8oqSbWVLoyjHFYPknbDY/CQGYooJC7OKMmgDGyQYF0QzGAe/BRKV8SPj4
6ORArg3tNg/nMuXhbvcKWsfEkYi2btqfVJI+fXd3sZQ1r6BYHmqcZ93vgcL5
zLLXoTs2MCi5DsbBgFr6dIkjCgO6ABAI58W8GCcseXpvIiYrm7zc1HsaQtgk
YERZiUow2RTAG54ika+X1AvBMYsGPsj3Es9m1iLHz8JIL35AB0KGscDb8QWR
/20haIFPg+Ppu8kW2+p3ymtwANH5Xd72S+eZX6+Fvg6Jd3M3aS2thpoAgQ1A
ZgMRzL/kuUygKQdEk3DiWGo35aajq3v89HWplgic88RwHkBLuYOhm33T4oPh
4SVeLGo8eIq/Wv85fC3gBFNujwjrRykyFzRISydN45YVig2zPXIAclxNwxU5
Z0S3/f+AXZ9i6ie88iKIgQWS2nQomi2V3Ggu174YGHuoSrcRMTWDapfz2t7L
4xMB8PQaQpxuCGNpq1TTjq5SHyGsb03mQR+1lciPPscxFu2oYkvFjuNtj18h
qnx3erkOl3HoH93XSL+5sp31vwDUn2p6NtNvOsD3he4oba2PGLxAYvKv5C2h
x6uFQnrWFvT1Ez4M8xiXUK1nTtYPPUgKGIKXuyF6dRbvUU1ec9NgzsXUn9Fh
ImsDBwInKfX7NM9+N79nU/vdVkCrBYKkKqy/9Iz+oziBATr95GFdKKlghSmk
bH+WmxXWcM4dcvIqDMpb4kMW/QAxgPZeazv13QXYAUW8hc+v0MUUDbtdJMQb
2sa/ZhTqlMsVP2DT/ypxBYZ3VbcZBeWML+A7G8Uez1oM+cf3rLa+uqCXNVEU
VVcHk5h+xtATG6bsCGyZRwJACMmsVthbgd2pLSPV4kfNPTwzuN5JOFpKPSOw
QQH3z7+IH+tVWeJ39CXj1vo6Hf7ZXqr8+Yh1uq22aOA+Tr56msgoV8jMEn9Z
K1EP0mgOwItqu0yvV+9+TvfXt64116Y+MLgY9EGs8Qmp2RWqZ4bXV+W5eI41
Jf9o7IdtEKeWsnX2harNcBEac07/hMxXlsBlbUKXcqMXsIcGvkPAWdyo1geF
Yta2LN6JN2KkyR9uY/zjuukRRrypSkbWD+VItjuvFHjO7P0V5LKFmZ35ROT6
BNZEI5HHP+cynv4im55AjqDaE0duKlXmJpM4Jqe8V75FzWl+b38yZi0hQyiV
lqR9HqTvdUqlCHrKnA64UeIcNfKVuW6kNnBb5u7TcTorE7h1BQ4Vpe0p1IlC
u1DUgtrqT6enMROHfItA5B7dtiDVRToHaJ9yjI67u3GUcyWj1nUfFa2CVjr3
7x1lgy703gwVAi3LyFvGZIFvuG+79DaY89DY2HPn7SQsT8bTFjlf4DCo8G5Y
+Y7VXarPyBVvadf6sgGvnHxlL46bDyG2qCXRh18gH9ExbVrGvYTl8eq1pt9l
/ZdOHBKvnRimkjuaiFSIWfvjjo7XpB1kcGcF5+3faLQurCfG6y4pHpfTN5KO
t2xspbWmsOOx6zgvsFJfQntHcsn61qZftVFn1qrwozQH/+sq4xC0ePzen83b
ki0AeWvxBeH0RVCj0NiekUDusoau01JOAai67+HM6RBeSLg7aelDA8vdw9ct
oBsVp7SnHirZmsvYklFuRC1lv4CFFSXFN3gqx1gA199SRcjURlVtHxYykuSS
tVqgBP7FuedJHlwtZyiw2KAhRTpAeGq9SClW5i6WR1fQhg0GWKiJNJoyFXUI
66Ij0SETnBibsCvIcoSwf1eet413OzXIjRVmfCIUQ5tnmzPeBilALPykg5sR
gkVY29DvNOS5lsncfN+uwZZZSnkIXNjN/TlEANQZttmCxFuFilsNtbc4Q7yL
qeHwI1j9sNeu/xs64Jd/M/QM+Onm5RQQrgDfeMoe4vD7NZ67wZvZhycKEDOz
KgXBcboPwr+IJY+YrZFUgd/7EsVYgrapdPfXdFVBFXbZaLHErbHjSzDWtEZ4
Fp4rkZZc1MPcRPAvy+ZuQEIoeiMT3iH4jawCGXwnIuIDNxQ80uUzGB/ggvJv
9m+/kkvuQAiPok4tuAmcCA6+dFFxWI05udtD0N40CoI7QK5dVT0MYMOJJwxy
L2kurpikMlDb12DemUHI1GKc69UXfI+3X1KTG/VdVSSJpZdtt84aLyVAKQc9
iPj5WQm12ayrFQxgpDCsrPl84pzsezeIIpsqeLDVjYDB/jTO3iVZ8LpkB/xl
f4ImDaQygTpdf+rVDSA8c8YUZLKDmH94D5ygNdNdedG4PErLrNV7eeY2upj/
+TyV95aIoebhZXIKF9PLZHMuqnTj2qo5iXyI7MYMTrB53/19gAPPBTDwqRUS
sJ6J1EWt2T6bB3h6aLQdgtz/jun+2KsoRafCu8BbKHMPX1mLKGhBgBHbY7Lx
jv/UPufhlNk/bMKZlFUO96tLgulD9UU4iJF9WeN1tZiMMuTnoE/31oPaDTPX
HBCA9pkw0B3eSsSYd06WTyOESxGS7TE8LpEh1FsA7Dvw2dVkv6KXhZ/zKt8d
7WYbbhrF5hcuSqLPvb6ZaTN3kR/labpJ4f+sdA0D7Hmu0s7txmtLTBs1713l
++jenWMcedrg4tVxRokAaoHmTW96YNVy+fUCCT0es8pjSP9HSOTLA7mjDncW
7ZnPZ8MZfckzJHFvE5Xzy1J9oyEBf4t8X1MTni8QTaIHB+SMkj3YqXw0cNPv
tf883JJZyh02bNJLPM7/BUc8BPhcBlHprc7D4/xIyO5gdajAyYVYrl//8i1J
j6ga5iZvJzrpBUT0m/wtp2dqf57SAIrU0rvnIK2l9RkmOCmYMkd4fSjqV78z
fnpKp3iunIJiCy7uC+US4toaW3105En3IvRU03qGO0OZjhj/4kbwIAlJIgd8
DQlh/rwICv4gS7sIVpEEdvfiWVOZXbqdW0RFndDm0s6AAqo6TnAr2nQ1oOQJ
Xlhr4sTtl0thlZMob5KPYH5Wkf8/mXyjGqUADPtBa97cxBPcb16z0uA8ex5O
UGh1BnY44JlBWz0w2fKH0t6AGDLzZI3RyT/gR9mnH5WrSpUUn19pFfy6DyAp
5tcrpmp3K3RmI3wV86Y2icxrAnQuDlQEIC8UkQuycoNa9zIZ28tUTdqLTI3L
whKxP4uXuVSf62OiQsGoVW7nONV7ADXsQaWc4sNNugSWHG4+g9Oc30iGd/8u
EEy7Yhb0SxKPg8VgzdkCqQR/q3G6tXFG94aCHam27GazYzSd2uMn55Si3m2d
9EiOquhVtYWzcdB5BvUKh5DzYsC1oQMfLC/oLWOT01128R52jmkvMUM5wQx0
6Xm6Wn/aoj7u0eXbCL4tC9ekAJNv5lUxEVWRyPlMZ0r8Hn1EjO6MHdgzI5t0
IEv5jj80acBSyK0SfDvQf1Z3Vo9kIpFrUDkz9rWzyl2AEgcNyWPCSXJfnNw+
xO3m5O31MAqX+A0VpU0mm56REcbQx1dYMvsHK6GBb+Tyotyxzt8f9AtTQ7KY
szzuTHItx38PLIZ23HQ07IMohGu+Xd2xIO/Jb5RL+DAxIOGSC/njRz4xxatx
C06bvZvYFWKrp9JidT+ONLHokNWm/cxybjhVIX/UDAhxU7caM/VQt8E3tAyj
1/9Y9eR1fTmTRfBVjCKp9ZfHTgJlNuRmq+TPYkBHSCcig2asgKRK1mxuHFQi
x38DAspONNZUl9nEuxAZLTbv6xBOew88WoJlIXHjPt2L1aw3kfXx2un7S0X3
wsFBvS11Ik3IRhU3m668y8ah37lytGzQzjdijYZZRrGrfD62nX0CEUy2+5cv
VWyQmNKPlY7QExjNuFM2uhz0qoIdHKwP5ELENDekBLkBxWMuedwjG7G6/KOe
F0FIL2rzwmSZJXKffg0Sm8RDp/0nxUpR/cVD0iqqR3C/ICPsOZpSRvBDE8i2
Wd0WyqpEZlLuHAWAMdNsgNq0eZfNQ70uym515CZHsOJfZI5wryaQa0jTHBsA
ZTLhBSaduMS2HPADnKRQWaYKL/yFc7mKRuWfQazYx88qfaxjHk5tn0Kj0OC3
M0/2MQCrWLtn922GscrL4m0XlbESUXpqU3aCvgVzyqeMQodqEl0ChN4GJZAH
2aaxm60Hb341PZNe/D+z6bSDnUfX1wY+PPHqEow6RGzfRvGX/JkZnSVv583E
sCvGm/o8CM5IECwF5Ghs5syXUhRhfAAyoqRxP4rQBHfnLYCHNhAOV1Vj9MAC
UzBR3XtI+Ve+5dZpJgQWmENNPOIFVxO/Dqy/+NYIF5dhaF5VpNnXhJzUfNRY
/xpjyVfoOXZkV6g4Hk+YgUG77XSgJ5lga7wPDcoxhkRFaQJ4UpUaPNhy56ll
ikboZBb4m1HmukRhLMPiiQSU4Zv1eXe4l4UAAbrjBmpmVLvy5Hdcn94qS6Ia
JpJOm27/4dLw7mGVYHr0Xza9qPJN1Sy0dS9VovqpzVWLsW2JKenMMfhN18cm
yhEY8dZfTl1WQUgMWF6TRaFGshcWn+0xzUuxVXFli7jJzB4reS/IHLNTki1Z
RcYWQvPk6Q5ypHoTl44M2ENp/4ufXL77sWy/Sd/mzetNrDIAxyEFpNUGReNQ
qA8/aYQDHcHgIpP+OWG3o8ex+tnHu5GTde3gn/MR0wOchgVQxNHlRxz4b8WB
DgoFg0fn6uEL5gzGTM56wSBiIxTi/pLzdUpnCYyPeogxtafCBfxUEBi5QckW
+LVxm8qNHxT2IQ1L4tl1zi7arZH9O9tsGJqs34A25Mq9pdpiebsKQ5+NrPZG
CI4ObrlRebfpf6jIFE+TqOUIXvuofRYH3WJPg1GhujHQG7c0oXmOhc3xYKPF
Yhp5UbAL2on1c43oob7BdlbCm7YEOKgU4hxy64izfsW4pDBH2iTVU0q1gtd+
7Y5RK1Dy7jt5jWYhmP0URw50CRvER8qyM39nibBwzBKIX9cAuSGI96Ztq3/x
SelvBKJRL6MRTaeDls7tn1wEMo1W8GU/pDbhV67GPyrVr9WB/QGjdrV3Dixe
UuPy7Uj9GD578He4OEHFyAvRfBMFbldz6R/vdOOh//xHeux3q6D7mCDscZ0I
sg/tIfT6CVJHjUjjrpvUFs+urH1RS4nxe0DANuYce6RW2U5c/COGeeCCQj6+
meo29JvGslvmVmSz/x9bLwUF2JkSXEkn1H975cTDqdp9+qa7F/M3LFQZEF+Q
TWdgxBwKHFUwNWoGnS3UYeYE14WCnnu96wnniON0kactpoo2rjakClRTSpeg
S2GdnAKqphtSaYBmWElrYh5FRqGmWsLH2bo6ppfZI2UoDsmXVb2ZKUA0wDYH
qdo2FSivm6tggyakHZKXN2kl0BzcmwJkBaTIFsNLANeZz28+iBrKYDpIuslV
ublSuqFUjL17nbVfwNfTzdBYyUPKh7hN6z1DLe54vk//aNfiOkos12dhX8wi
+gUT4vFxaBDCzDTYfz6gJhG4D0JvQ/9xN1Gw4iIXJMB//1XXEiDhjtNpYXhm
MNYpC1OJZ1PH4DA0qs2iJbQjxoWNNBrsWRt1isWSitZL9lKJgUtb1wEuiWgC
6nosEia8HNTqKLLpKA8w/EJ5EQx20701VNjQ8cL5i4SLKAODA4IRMGt6Cqr5
KU/1seLFp6fZ50HM1OLuMHI83ubkAH7YlCGKQVxpMeD+DCGyWn3sh6W6AClC
YRtI2apzeExBydqxL/k1uEQbIixJrUdKGo/FTsPC82qmk+dRHgz5qEz6A+CA
rcY6hq4iFph7C8PFnf6ezmGUAFrFoMTvQ+9QCnFWU+bk2rG0N1LDyXaEQu7y
CPmKtxDtS2fczKmJ4OhTzSDlbLw0A3WB4PAa4rm8AJdc3s64eRYefzWEgbMG
ZvzRN5k6YtuxaT2FWsdVpRCESHCo9hvNg557b2YFHaHHgOjoxdP1pm6GHhUt
GvPwfVoVF1MC7xhe2BsZnVTkORIT6+CtzMNzJsU1VsHUXMS0t+kvLvXsWsQV
hv+PNUuFrqpgKVHkdPY6DMjSHrrsssszpu8rEWyPqY3eCTOwYfptYSmxu5CT
d5Iw1MZQa3q+xfIHaTNQxgyfrm3Ryd01euXo3SsKeEbiU+ygmDIEgItqNPVK
I1fyncuBxL0mUmFRWppVHahJMjwBNF4gxCUb0VN8LI15S29oYQoo+cza8Lux
34J1KBuZC6vTrc8wT0de8l3ljg6LPgDbwPRkFS++G61XhW3QaJd7iapyyIxZ
TLV1Ch55Ngosy1/ntpNBQxONi4TOrvVSyOqch9W0OLu8eyO20CwhdubWi6ih
YHoLxaKJ5NpenP9wfp0yMiPWdFnfLUeccB6M8WUY46nVapvFzl1645NURkOg
4xuOMFRdPtJflj5t89jSVsIye74ihRLg44qLNpEM1XXPHpSAlZHBcxw15A9I
QqYuBDmQVAZDT0q7CBsAiA9o8HAYINuU1LF63SFR80p8CIHr8MKowb4/a2yD
s8M+OJmw1DZiNdn2cKqEqev4QQ5oqQUt5x4D79ohYurSOfxPq0JSp4JC6Fwc
bnAjC67rWjHUA+ixZIZh3PqLVTPZNoAsY05U+kXFeW5WicERhs8NJ8AEjL+7
wFwQRTmgZeZEmLhUGlGWppLlwBc9tyz2Q+ngl3mIG6V82HkWVYdVmKk9w2j8
qWOkmD/HxsoMaYpXlLsaWAJOJ1rHo4vO27w3DRPPaBmuKd6EYMBMhVnbkD0w
UXIirrrHG2A/VzrPiIm+UR+XuqV8TKkmDN1QonEXGqRxBzY6EWUCYHi4RLei
XxVU4ps16s28l9lsProZLzhrsYQl2UG0N81Y0JeHf0kBJ2KCKVHPwbADb93D
KshDrxNOnxgh2YjXpKG7sSowGJ9QxtQSdlxtym69wLVl2rlw41zX4bKnOzB7
yPNimExCYQCSWBcvy4F9N9kpicfFUCkqxvt2vuBHAGquY3xiXJZBKkAF0F9H
M2wvzOfMQXdJYS5UsdVu/FW8UTKU95o8SX3fsszdoUURQe0A1RTqcT+zzFSu
RqHQjFmUWCIrZ32GA3iLbxuRka87H+f94CGCfwHV0LLQv8le1YiFrP/lObCY
28jnN2dKc9YcTAxR2P3UysHYsnIrASGWfPgHh4EBCHQFoIyOrZDtDMnXhPVx
0nJpNYDQSBoE1+PITP8DY+P9+vzIMV1ey8SeBSaowT6opPTd04+4J9QL9Q9D
sos+Njx2qRXU6TwMWbSlhJpi+DapL5p+JMhjor02Za+NSvuslQzHYzJUDPHe
zBm7PaeqRCvyyu5FKPa/9u/kjNhCfnkSd3JmGSNCpdZ4JFGufGTsOlyp6SZD
/U2W+GoybcOE98fEzioY5/8+Suhhon1zPGAeLfj0sJ21BSVdCTdmhhP3U6FH
JPM1+dXQhVgZcVyQlhzlDGdwt8f4U0PnoWllw4YLZPxgNx7DWx/+5QHzWL5K
MJbQVD7KbJRxQh90Fq++x4uG3eXvnacExxp9D1H90wnbyFBPVWqcQhhpwaGM
TzYkHD3yh+pRsvL//4DJ0HjksVvw5OvuuT2Yh/pArW4pcDDgA2UIyI8pttxP
IJl4um4GCx8y93KOc7I4tbHZ32ANkp/PmCQUkcFbiC4DgJRxVzZvrpJ2wj8H
SmPw1xOzSvU7YVdNIx00d1WnBrk6xCObXYdwU9gMpkvDAYlfwmbD/Sn5/bvo
vMT8+Tzsdh0T5eZe/nhcT0SXwzTJTUvPKMryz7HFX8E62dhQMgFR4P652sAi
ofdma3w1AbH6H8VklBoMGJn6auHlkzhw/zPR5+hxRUzvSNGQj+hnmEJdRNnJ
4wbcP7OarkeMQzk09hQsyqdCXAe6c6szxPDbh1qNQOO15L2xb4qkiaPvBb8G
AROfvJppLeUk+XwDMhBWpeo5k3+TJozDZE7h0SMAMz/Smvy5qZ+/SXJVFH7w
I8p2LWYJ0UQTnrP/shDOWC5c/FxKQ33JDPc63mn+au8LZLefLnPxVFhocfTa
ahcPvv7p2Uef3oK8CL33OAqm9j4B7/tnX3dVeWmCOAhezu+RbaewapmIvIZe
ICTEbHui+8REy2pYrCtrBoHEMzZ+2AfXJDpg156DQfLxpzVmxHspytK4Pr9T
jvYkJifpzUD84hTomsxvCVind2hWOvf4FGsp+HhSBES4IwbfROXNPnE2/dMy
cdfvY91nrwpzBLXGUz+yR3RCYTvdMUcgOvPZt+KhZa4hS0VvnXJRtNTxucQQ
CTL3aZDxvSMqxxHlQCa1o7Bgkcqu3x0YvLBN+WEtu/e7gDJcDX6oDf3kkWME
oyhoXv/L9fvewNzUESsjvI4XgukZtJ1jeTk4UOqLyvBMjhJ4D9VxARa1FeMt
Ky98dYS35NSfN8Rpz0+td2ecxzfXiVg7QkYFI3YBpG5CjJLfucOuy/kTWR8J
BWRONT+cN3jyIWu4L9ZY7dErMtkqRU3V/DW3Th39vdksNTmURdlitSCTNi+E
UO/JzgA4KyKM+LekghYpL76xBsYTv0iwqe0Kxsn0oJ1StMxwJammYE9xLDuy
557utRn7S7vcx2KOMT7ZQ8d1e+Tb8UYzqbmKoWRKz1ux9gngPrUq9sEovfGr
XKPEM9o6WFZOSkGxBEcqpRGYHMOJcz0uEkzHRIIXuCqvCHxOs0GvRk4ABty7
fPkE4l1aKzEeX1CQFZO3wHkXPe4h8QUI8EYxHUjvguPQLv9XMxbz3f7PD0YV
O8rkK00D/uEKDd6J8m+T+S8aZN+zMPgWFlhUwOQz9BF4l2spb5JCNkO7i8Yk
72ux6kI6zddmA5mB2jFaL3cmOCIw7g2KP2lCGdzhSlLsen+ly/XdbWicsoOw
/26h92LJd1UdZglNfiP7iGJNgHbENmVPUzkSmQvh84PK2xTRYPAm+QDNGzNe
gdDHdawVHd28afIqfhs+l5lreiJrWp15XqLkLAVK6XqJmGC7NPkJzdpO+7c+
ou5Yc9Iv9JQDKah6Bi2G7DDFSeS0hsjAKSzrQoROhued8+l/vSU8WFQzD5rH
vUyLPNpvm9gGrB3zTqUYcTVTgnhgBWRVrWO3/UgVZ+Z/wiSLZtxY10a/5dfL
I8AJqs2IoAP4LGBf2Tmgm9UWbIF7nuQX30qtWa+wxYA8J2Ho7pd+RiaR52my
Eb+kCVs+KOK5Cd/rVQOh1w4msAruz3Rbmy8pXXJtd3b1iGtjXa4F7BCAPrnB
JrEPiPjXddTIPYqcuepSdYT0KEIOpFKMfIlVZFlE7+E+h/CcJ0iXtffT5akF
Vx6OLfjpDKLlJenlC0oSH9lWJrMfsL8O04hIzoKnLD8OrCaE8RAkGbYRNIqJ
tkUemBmLrwUfrvvxNDKVWEWRBJQikaoSe989DQ8u8XBEVYtWCwkuVII1235W
40Xx8jrurDpVzhMQ7QrWGkJxhkxsMR5jnnfQV74nLmwLPhuUrCyTc8fjsgpn
TP52+QquV5dLaP1pxdi3gYpCPAfGZVi8/UAC0GvfWzlQPpIEeT+qw8ZXNbGL
inJs4k9od/5q/tPPoY5qHU5l2HHUr3ey1f/jbRFsunZc63xk9MOAtG4RudVV
FVdIa58OVxxMjTDj5Lev2bdfOYv6PR9xV1AFPGW9dpwxGB5nFPA72gC2U6/O
C7QPG8ClULk/0zab1L7XNeB4VRLgVt3fSXQaCNqRoK9msHHDeGlbbYP32miG
Et16NrgsD9sK3u9R99sLsITx2PUOG7XghILYf5zRCl8vwBLnoXM3wq7+UPgC
WE7f26A1jH48ukMUPDOcFraK7WAykjvws1UjrRzBznF/FYJAYI2Bu1c74gJt
9i3UR9WPY3HrtaH53vXiu97Pcg20mCHYjNoNUy2ldUnyQDkrqO35Vj31UJBW
UmNaVs0Xlfl4bHA30e1XpvAjq68MvfmGi3in/gMSfOLDdswd1e0NNNj7gIi7
JVbgGNqkidDIroIP0JgtHhK2IL46tdHN/KGc7GdMyiJzYxKOc9+gBmGGl6od
94sCIIPgNehObNwuFvQQ7QSjHlAmJqPx5zSlOPw7J40K1dkvGiGJguUb8AC8
wELMaUXnNpGWsEFN0SeL7wT4zd60I8Cxk1KoJ5CdS4Po83NVEkwx0tuSVC2Y
5MgukCBHyIGOPRgRdigKuoIhxTW+LGYAnrAM+GdK+BDy6h/85ZCwX7ARMM3L
n1eG8Z4wKXACV0ZLEsMAPAPNHu87Eht96FeliKOEdWmKKju1yMUlNH6k6YO0
l1IZ4c4ol/eODNIDw/3kK3c+NR/zsPWTTpMWK2m5lo6I/ZHaBrZFPHvLfOSk
gWIrntI+14EEfSPbUG7Ffumw0mavNVcPBJih4wo5EEef6W9Cblr96BdEaJib
zQh8p2iity426fcmHwGMCwZfpeqzzBa/Q5cEgqCtWlvUNVoCgi8QpuGDFBS5
GAP8XlcEi1W6Xe+4i6r1sbSFaRQ0oaVsAm5tYiiu373zXLYZqK6VATcn8nYx
rS3navgNSWfZNShawAYFOJpg6hgrByBsLrzxxGfqjp+OASonM9Tz+nH0XsTD
nppZPEXkaVSUG4vPPkk76vyJjmp+XThbQ57EhWRMgQ5k7SsooJAYhMpA1Eq4
Rhu4o/zwE+BlBwtVVrxGjLn3NKDmt9kn1WIzTHRsp69p8qG15vWCHN2G3urm
EDTkB4pFWeWSNbJPNbIXqn6KuqtP3xpKH/U8j1PT8w8A53NE/VOvSU6FHMUz
C/XWwxHUDdNXiLp3K/5acr9MGvD6RCZxBWkhYpv81vjvXMvjcINUIu1Qdbyq
b8lk/BlAc2Lt43R7gOg3Tp7rx8asCRldd17PK6PuaBj6uA22o1nwh6mt2YEd
K2Aia4/iXyOBDuGmnwMrnA3sdMkj2WsO1TA0Dpfv0P23h2oGLfV3fhnBQi3l
Tg/woYHFQatxUp3FPclnyP/zPBOpycnn07IXzc2G05ygHlq5ovY+LnRPpvzt
TKYsJU/BIgIJgKQvL2XFN0SVTZP5fIleMFlRBJ55+hiO4NNOlaSgN/GD7wjV
AKKhrvp7dcIudo7RL3pEdu3xz5NvS39tIWOldatk9dIQM5JJlLXh1QD8YhJt
vyE96zC0/+UI7e06ve55qigDz+pQLSyS3UselcNi3e2xtCruNQ/yi9Ynprtc
5aDv4G1Cp3vsl8ofgSe5O0RAh6/B0rv/CdTQlTWN9edCU5no3+DmBI0PR1wK
o1KFICnPyrMeBfH+nb0anjNq7GS4Hrwld8PIWqv2TwNunSE/JOk642s38htZ
kJWUDLq7i+vj5etIrP0qVd8DGg07vxD9sjt73r7opxBRYsrmtpzGyc0kqz0f
7alpYKNhxZnX0dtKWGy3xpRgXL8NVFOaIQSv7nrq5mJFKL0BQrGZ+TizdW8s
b1EpigQLr3F2848/SmSKKygJuupcwtjreW6RN5wr2V7PthGfK0gdvjq33hoa
iFROAcwZlGRI4xuqnufcS23TFSx4CAQsZep7drizefssmzUxRXXKi+CALZgX
g3grGNZOIkAMH0uKHSvl75fpJzKUAqM3pP/h/ZhUxC6+BtKvjwZnCjlBHB2Y
p+HhnV1Ut/lxOIF7fyTEtrIQMy7xQ+0BU7dpNo/m0UCRRjE4H1fvskwlTsWq
XXU4Lv2ke53/onPZCpCztUT/VzwZEn56SevaxUJTKEJyoN7hjh3Co0lwBJTX
lgtDHiJGI4fv+aVPXktJ8+mpsLFCRXug/Tk9zX206TSxm6sLaW2fnDSdx3md
3z6yOjYmIOwFSEYm2TMByd45SslgRhocovWb+Pyp1ywsK3AwbBAqqJP5zAPf
FQTX4Hqu2jnAFDm9jnbrRd7W/E9SX9xsCB6TnPpZO8tBoJz4+i7ucZCyM7Dj
WeBA+0T959gOZPZhrTr+PMZQ/W34j8QIZJP1e9YnvXuuq6NVzFq5RnpuUJax
oupYw+jI/d/6r98ikQfAL5j5utpF35lgYuFzOTuiaeXULeoJxn8vdpcokEmt
84/p9rMVuLPg/hlijAzlU5qa3FVGtfQ4X8E144uA/ybMDhxji+Ne1VRL9DdI
9+yGRK8FFfX0Rzdnro/AOMjhXpzUT8Bm61F9F4st+vxxEroAePX/UpD/xDCz
0hGF/WLH8sw5XzYh1J2Xgkncz8kjSzNC8mf+rn+ttjY8MjCbTRDB8AqN/JXj
mcq6SCtp1Xiz9gLxPhqFpGZ0c5+2A3b7nIUIy9bf78drjsT20O03rdetjaBT
v7DuXtq2QTmHEyP60WXqevFbcomD/59awv0Jc2Glq3URJgOZJIxvlrPOln/W
MdlSiKXSuSDd6KE3ERWAHJsMxiD6xz5aEfZ/PkHZWm0n9btf8kboNuBdHzEZ
UVDsZZI7721oahYH2iWxRM7MOrFSbavVBnCh4A7Tk4vglUSsdEkpiubh6MuW
IfeWcZzODNWfdg06BwaAm7scBJAMZSZ+8cU+RQdHiGvySR2xirLPTwkZABTY
Wq0hJWKWnVDfz4naXr/rc+xNU+TL3XOP5ZJsQsWxbYrnA3eXR6iEXKtVJGn8
ect02j01zl/GKczKquCscxwCgVl296kEmrXksmjk8WpAuX6a5XtJBLCIdgAn
xbhwX/w1HERjJZqD3VV7EncXIw2MVtZ8eF8fBkovqnTeB3vssyVk0VE+xJJ+
/iWgrKlX7cZH/5R6VdqlUfQlZ/XAvgqEHz27CvTLVCWeb78++pLmtMYJ6Yr+
07a9OpzD2Ze+2sCxH9E0BEsiYvEgbxWSv07f4UKYF/ZBPihuNT2roy0ACGlo
81OsRwSf2wrEPH76ZhGYfvrpIW+ZJIZA2na3izdluEv678eRqAALtLrA9MQz
U0/m9jJQ8VlOGevP1qPD+u3Xy6gYVUCbzA4uFc/BF3g2kcOG2hbIcHqn1jw+
JFsscPUTU+M+aoqAocQcplo1Z1H2Dc6WjK3ue8JtKoEZ0ibqIoh28z5e5RCE
CuN3hHuAkaqDiGJcSiGdZ8655qOlDk+IJ/Oco4YVqYvB97/5FBBsVtxOs9Ct
nQAsUvHHff12G5PJ7FRs7oNEU9O38OmhzaH9P0shkdWgtAX9BkhQ4RR/1LeM
fOhWnatHcoj+Kou1EX8UOgeLfTR5L/ZNUG6Njchozg5AYRxxUYZat0XuSR7n
3f74rOr9YL2dWSxzDZLgWaVYKjsrGwyp1UiDqUxlAh3ynhiYHiQzDfVZIOj9
SFlUUuf8aSGnQ9OHaBf0Be/Ao4prwbQJOJYn1EVK4MsYa1RL1VLPKEkuvlhI
g1DEBSeUH/UTCxirjJjGq3/0a9P813G6+eoSq02SY92WhZ046VFuN/jnuvCL
7rgYbMoMMlzWMvMKAQ8LguXhCSzxBqhbiQkPip2OITtFbmx7G7v41hGdmgUB
BX85jE+W5EJUaFwEGa5WuQNSnHM56GXFLbgLgAYNflhTLUCOK9AJF3pnNtSM
E2tlkUTLUiPC1h0zujJtddYNr/kk24QRK9JpUEVyIqepPpNparnMz9PCMgsH
+iYynb9+fo3m9hpHw95KNgCwn1CtYi6jSvFNcSG9QXH1Mkc8Z9dsm2ZXzup+
7V011ZGC7wfiKNr2kBF5QYSp2hwDLdz+XYt2G5T1q/sLbV8WKQtC+BulozJV
VyQLRkqfbCj2CdLku16GhxuYXSg/biwSd3aP2u8PxEtAwmmX+kVJy/NOh2+v
sTERa19ALmWFuaAmvFK7w1bkGsj3MIplsuEbI6W8NeA7KNt1/rI7sYC4B4nF
RpOgxiYg9YpBBVOLZeuKC/XAhf5TiFSIiNh1PzweoFDzxrmEWcgEoWYu61Uq
I374OWxu7SgZUG9ayQKAIrFAu4QwFTJdzL8Gj5r3kzhy7YFKZVNvVC7pMUdG
YmrdcmhPNHfzwjFQMvmqBYYGGeUmUI+TNlFyS83YQt2N/DPyAV3SZ/Fb9Wu+
oYZ6L0SydAsN6Rqj5fsfEjT2t9SVIxeIGiqKGn0B7HXaZkeEgsG3irkK71uB
V67a2mxigqQqe98uAy7w0LBrbTTFwXiwOlnQLnRvqo3VByXlx7X6ZmqJT1/s
AhiaSM8msMgbYjoBBlMFpQolpeEKjvPVbUwVXQZXvZdgLPMGBHXPlkdgseH/
S7VpUlKuAlHUeN5f0bk3BZJTgpACeqq/KFsL6uCEKOA9SfN8IIOP1p6vgBHV
zGl8GgcjRDfv7wDLORg/U9FSgLYtbsei1LPbxZWoBF3ufVdXpOxnl50ctp5w
zDxSa+Yd2zSTJgAmrWJ7uAykMK+6vbv9hlvN7iqjbaH1tFShN1QnIViWWzZh
gB5YBMrjfOyAkQIfhewblrIY8wS9syv+1qsYQ4uh5Y25xldqcLtRk0U157dk
IKgUQp7Rd8NEVI3uPLVLpHfwGOWtqprsh3oj9VJyeqR0NNr2h6u5M1xu3gSQ
4AHdZUPBEzvHQ0gyUY/e1ptaj8uiljOVpavXW8sMH8/MuVRlvbtbfXxAYPj7
pbKD0tDbFsOaq7E79aOLMAuOJC3W8UoXMEOfJ16++5wDjScCuetQ1vgxnbu9
wQoS+IPUT3G12nqXXzaXba/XjetVHBUf4befsLal2W32Eb9N/aRc2nBONghN
CvTBfq4GddlJKmQ2vyw7RlOCvHxaf2ACLrkuRDtf2Y9fZb1188AlBSJx8FJf
pxv6JqzXHR+NBImCtZf5NDWgaGBpyQNecSlpo3fajeKtI6vWM+4aEspGtJn/
UqNzLAXYlbi+BMKne1RahrqV70xQpAXj7A/Afc8J14DzJozTCchAw72TWRYo
KsPciQOMrnYivoEh/sZr7Y+Ve0DQ5t19Mc8jH3Gn7vMeoBE/hOV2LtDnW5Ny
LbD9xyfUCfZopc4vWyBX22MRKAVmuXiJKeUOpQ1UzVzqcnI7f5WnCL65yWZJ
vYPpZy8EpnYnuTHTCE+MXYKHH8sh1ri85Uy/cEIOiIoOpBMUiFOpn1MTnTO/
dgDPH0wmlIfbbBM3gBrp3hPSq6M9wi/cv8GviLoMYX+gsYbZVsF+2TNAAfTy
ETv0bFzelhcStvswzVTaByqGDzN+Npe1UcMYmZ9oOEcZVjRfWD0E7uivS94V
0F9PTPl+rksxDM0eg8Z2AkPWeEIcIFGyM0rttB1W46SQayiJZkGZ0bbCGi2Q
OzJB+VbDA4BGiAs2JjpNi8nsdhXqoINOkHFmdXes3Xdz8oziXNo3g+RQJVlp
ZonoULGT2zn9cKQPtVVurkhtrFt0OCT3JrpATMvF7pj/cvhNjhGdRjGWRwpg
a4o1ae6MdCG8D8S3TcEllS0cWl7ELRkat+HoaRweIJYmviSIkIC9vICQclan
4RISITJAV3GBR7KmLLFcmm+pkCCm1IP1hSHO+zGlS/EpKC2HTqu0Th4/9WMM
1HKm+7ORY1oiOtKSF7PyKpF0lPbYSKJ+8yzLEdyhlrgE6uSUsjWA1oukEp/x
hN0z4lS3aqKfuhJRJG7FcPpTIU4RTO1j/VOfwPoo+iEIzOvWy6Keszc2YVX/
FkQODtWabgQvs7w1kgAQmTtQVPTkrp2Q2kgQLcf4ZoD7PqHzBg86vpKA1Nhz
70YzSD6YygsGhDfBB2cSRFGUuK4gyMLOSEA3WBnXVl131olsoPjshZlworTQ
Hffk9AXav1J088Bjik2IwLnknjkSrX7LDDBp7emjhJ48ADG0IY9i+5sHM2DI
9Svwo83OhMXUWzqtowAcapPsRES6rvc1b5VZ2SmVkjs22CrzmJA/mHIWUEnG
SUXfdf4wIJW9Jfj4yejNfP8bluPQ+ZeTL5h0dLhZnQqQrAFYPpvyNoVhPfnW
fh9SVbe0da7Yy5hmzA0ietDsTIAyhSuMcY+wK97fel3gntYxZ6jRkJnjtwY8
SXbtq9johut7aJnkpteRKPqc56e6c9iBQZf5kAMT8Bjk38Eio2baC7Y8sywq
H3PBubEd0L0Z08T1YVGYkGk9FQfa1uNSvLig3kkN1a86E/8ArQf6F6Qq7la0
ipyRWadc1GbRAKN/DdOU3mF/a/7mkCqmtXY1VhnSgGpvD+D3vdyT3f3UHq45
dc8W+KuqRZ9q9O11wthXZvEkNGjEesreIsAZKy57E3LAwdjLN8LJRav2CFfa
9IpWMFxS9bnNw+f2LUAIh98EtTRMG68/nsGnMqqBfB3bNDVQhpovOXSeGlm7
KA2aDq0Hs73JkeFWYU3Vt/hnSoM95iAlNvsEZ1cFZpisqK21q0REPL4s+qD7
FS+5WzFFTl9dH+MHOjio7eCk5bb/q4Z0cXLpaFRB4NhnJgT8pJDXPvpYx8xP
05h53gOv3lRtRUpXFzZO6kDdFq8dStWCkjH9NCNBkaikIdA1/swqNfZvFEjg
6g44RPNzvyZPCEvhXCjeA4J643noDvRrDWuQ5kiLXv5byihEzCMCE6h6nwuY
9WtZIEQOnFZgYkPIh4DYC92aPZxj+IUMoySKEUs8yx8jDVXJEkLBLxHWsNEP
qdyw/8hW54e1HsTxu9Jkvd1xmZqdqiMzCEoXHKrhIY//hhCWtiY5RfPZBdF/
7Cifw49H0mQV7LKgxPy+WOhB10AWDtC/DctI6fqPxU673iN+GgLS6lrysHlv
OZE+wyQeL8AjI3na9RTdYRLFlg6mQ7k0bmX+YgT/2nlRKaaMZSeivH/B8Alu
PrbBMT6OMRrFe7XgXNZ4v03qqJbFlgOLVVncIydTrsUg0XkcEMfo4fzz1nAi
M/JMgKR2QdTi59wU7xvQaZdGxtscFuAiSe2XekqPKp0hbqXx2+ZQVEpcwIgu
wnSfxwKXKlvq4LypajTV3K37v082S3AOKeXSK19Efj6sIyI+GIev0uNbNap2
TkAp5N9mpwSdeSEV4VM3ZNZ9NiCm0af0GHzE+2HGSxdr7Wdbn3diCppVjdvP
SA/VOzYQKQ5cczO6TfpjrNjmihWujYj1+Q6kTJ0goANRZ3BFueYQYgYLLr8h
pZEi3qwCC9u3vls1QA0hCNZ1UbeFAsMltrHIDd/TwUxupFL6jvD9PbclaC06
fcu3l8LPvHw29OJHCZB0Rr1Xy2hhUKHUJQOcRowvsJuTNSmF6Az4xypmsKhG
VbIvYAW1Fh62+jrTXFzkDStjTRfP+xk/tJ26Muegq6SBKMK/ACD4u+8Y1dPT
/7Qa8/+vmuPgfQ6k81nqg1aFLUjK99XRbbWHVMo+en5Zpa3J3rG/NM8V/ATW
R2OZ3kf4mc1frgMdrHFpn9Wb14O+y1/4E1eOIBxyeDTz/DoKl6VZNwP9upC5
862zWVw0EwEIe5gQy6iOX7CQb3gnZVakNRCm4xNMWsb+J5uAJ/XjhrI2G1zY
JXN28EkM2311uQoF/4Uskfh8FcgT0Grp7UpHxoV7vW98ZGpY+20njbz7xFN5
fAgSK6RXkknLAnlpCVfG+3wliCPunkHcuWb59E4yfAptdzZe3M7QtReZm/NN
wdD8/Hm8T8HjTnxTyG1uxve5E0fNqawLOylRnjDH79z3Lmos1edZbjCl62TX
BZfv+Do5kzyrjVDnmZkOquMs37KZLpTQH64ATNFjqjGyYgCdtvGcepYG3fD2
/0ybIF/85kuA+FQMejHHvrVi1dM2cSVOCeuuaXvh+DteGDtoQAXr1+o74wiK
gliRNdzR1diKiU4UFazc2PiOklcNwNBRTkIiB6HGdbIUMyFqMyZFO4FUENmT
uqibhj/fCGNCA2HZmJnZ03FI0sZ9hnYl2HcuxooEvDx2iRtAx6kPccMYBAA+
xBlyr3VzysDXJoivX12sSp7BJ8KAuOYiuImbwPYYVjiIGXapy8YBZN5imvK5
ldMUFn6s5xTLXYfHNGTnvlHmLeQiqNPS41mRYB4iPKesyYnteZPPFgCxD2fd
CRtJE6LRumE3vYTJt08RXS4wOaP5o+ivuxpR4NFrofGnTSBI6htKF0OOymgW
muv+S3rSfw9DBxH9RZRb2oTiFFMZxSKmG6gMkn/bxrFtSWdsjytIWT0iF6Jw
bStt+pCIaV1+sm6fd3zWf/euTMfsYzfCVhq7/FnspnoBommfiAym40grAUH0
VX0bxvNAYWHjSCbbGRRDNaHo0UXxl/5HMtxqqawvnAvc0NakPNvnz5M3mz/S
64v5SH22oPJlin1HGek+LReBroWqwSBkyNgmjvfsS1MvoMFo5VcgId5Zf0Ds
wWiE6+1uM2PgZZRWQv9pPKwQahOyd2dF3j/BX/LowowW0iWAovu5nZUJ4lK2
63y+QT2ESOKGZCjG5JUKiQFHvwq7pCxvgC6RU0MNN5Uz+rV7dk8m0WiuOfSN
awqTZI7c8HsFx2SJNPZph0KsJFhvob1gq3ujpxYdC55J0uqd3I8eED28gThd
BHT0H+FFc6qcSqudm6gS7BaFQlyqoZoLWsf+yJl5vn/Nj/ROpbxDx7nvVGGD
WMvxGTM2uaWgY12SJcXmgb6rxebVLTRhs9MHc9SnuJ1T7h1wSJjgM8OKqMBN
lQ/EVbwZc7nu3w07qkWRaHyPDJhBm7ye02F9prrsfl7nogWm80vAUUF3u3L2
hVHoIYAlduJ/1rxbErPaI+mk5K7/ieRGjiRe+JzDxhRT6iTwVFH460M9rVE1
L8STiUSMjIeHFPYFqdXmctgnIuB/hzf8GMxweE9mXIEV19qnf0+inXQD8gKZ
en8MGH+mK8v7T5iTOSHCI38cxTgI0BGW7CUn24ome2ABEUYFcyRKkytNUZgd
YDyjV4P+nxqwK9pXdoH7P51/VhPwY0/SxzOvk3XyjghMTzLz2Y9DiJ6ueoIX
OEU8ejgT4MCam8n5gFGByyq+WGe337Pck3ZN+gABk4PRLAL9/vUkdIyHeNuC
YGLn2qdh4hitczQP3t0g2azbHNdRPE0anvOMaBakZX8bgTYnXWQWNKR9IFrc
5Ui6mam3Wpe1xgdV1wMFPkNbYcwAtnI4reCHAqHqBnbXrE7LShNZlPXjrMDU
WCv3QswYh4vBk30NDv3gf/a/XlmXogVIUx7ewUegoG6HeT6Wr2oGkXahLiVO
Ds9y7Vd26mX1bJLWlLA3Mr3GbWc50SIw6NNFcxOvAHGpJRks2IvkPQabVeGj
Fxad5kX2QaCzjsuppDWq6Q2Jzv9k5EvybZZzWr31P4jnQSFa7gtDvMsvgov6
ASX4lZ1g0flZMrdeLwUtYcWMvJPPqSnOW+aX++tIYJqq9AQNOKU/6cWGFS2+
Oj4Q+c/yxk7JDCWV0Vji9Hwnc4Q3jba+dK+8zgmMomyBw+HqW2yOHOM4XvoS
3ThqTulYCbHlzOP8PxKbNMSgn5Fra9rL1ql7ahSTYwexEInoGNxTcn/qLf0o
33kb6eh+c4WRL2TtUPbjJfWEnd8TBqi+8iIIFKQ2pKL1vL6PBl8sU6hWS5MM
/Varejt+vkD6mhhMOgEDa5yGZ81EfZDi8XBfZwoDgrCHJDZwKQ0yaYFrGr3v
jaifl7BGqIlQHWOvWTRvP2Kj/dTzQfm9/ezcmCHfRsvRe5hUcus9I+zVDjDX
UcMAci+1gKgcw6X2nTJWwHEsVcnX03+lav9gFR6wSEiGIhuCh1WY0MVH6X7e
xLHQ/mkkz8tUyMppmJtBQw/uwtWMCquXLto/WQ2upASUnWtnekUriXnvQU8g
/XT2iLOHEtH0FDvPgDLg1vxs45pPejcR+PVLanPit2Kr5T+2v/oT8ZwKnmM3
sllzprgIjp0MEQaPFKnNlqNtyYp8FO9G5qJ3fGVOhELOuy2K3N++cBzbJ27f
Rt5qkJ2Tl5Mu49bw+uDSffSs2JPh3lTANGK8p9dpfbm5gMi5WZIbL5YeHHPE
yceLAJFvDPM46Mid1GLzqiffybMNdAx9r8EpDXJAocYCDUxl8dC9LF/BX+ng
1NJeW1Vkvkf1KWFYAhkj1uXVtaEGleSJrHE7kZG9+3XuH8sx+YLB2yZlUnDk
1bdIL3ipSzqzIPxJcZ9GMVsUD3c7393Xlu1vi9Z9J7QLqidhnn+PxBQcQa95
Cl7BhOEDewqKMZcd42JcmrnrzyN48P3OEjHpX9xloN7GP8YRGzx7X3NvLo1r
2PtfwXt4YkZOXLvNfW0GiNWdko/uP9CWM0zjfsnQa+vWRq454aJI4XQ9zNJp
1qIQ2rWgcDxMKhkTiAymnyLzfQZ+klDGNkGra6l8VbbFIWulrj3Ka2qk85wk
6MN947gfQx4lxTELO6Rka10J/dXrwyQbxDfmrEfFv+hbGnmCA3vDMXPifFH7
dSRZR3KuHoSQNuH1W1AU6nosIjwvuGdP01pbpsuiiOBR+lWflSpShFdw5/LM
9uPIE4jl2OSRF1PbHsHOavEqI9kfgbPEGlGeyyUSqqY387/wEbqwabgFwSWW
mNUGL7oZsbWCigYaLxdSPgvnvE0jpPT5Odjgm1zMbng/kdCpq+sLem0fiiJ3
kx0rSTmwdmWeSywf7b19dPc4speQz1K8uwKbERNQFJRcUs8tNZeu9Il8sWiE
ngCwJ6zUeH1ftZEiKpFzmRH4JIi3FWAVeDzVzTp61Sz6cOqbenSv47Bk+Ymz
BjPy2lf4Cq+enD1v7C5DHcSr9xhfdFO8g5JX/as/GrZGKQWhhoIijyT1QH+e
Hv11meFBuCBbCIaE0tVIKXVkdPeUn5trM7+LE+NZSEZDXkXJM9GVgBnC1iYJ
7R5Pte+jSJvO0vXGy1UEuyG0h+Dn4R8048ybyh+Tm+YDOFDJMRoXx7xEy1Ig
lMKA9Ts+qLp7agIX9XCrjUd9nHCeg4Sfb27pCj14VMcjJSmQp6EVm/mzLqUL
i6ksG6inSoyte+YQN41/7nvtbqdP0rjvKTSTYvocM39FDVq98k2YMKxIl5B4
1UrE81XceN166YjVaaRUdRcm8tWorZQMA9OYiVPMOcD4a0mrjQXlUp2novGt
iuMgK+RWUINTev8T35VURSxJXLKuYBLcHp8LzBcAqGPSCYkJnVEu6GuLvTBe
rhsm02dRjalmhdntqwYMpzpZFFx97RuE8mbd9ENJ0O5CcwICM1Ns8hdajkek
i3P2kzdyyouRclySt0sJMEaELevjQigKACTR579uvSGiMBkKiSDR0tNEp9Cn
gdR3yoKB/PVehb6dQERK7nHi0FXBbi9bx5XXCZJoKWPvVMtlb5P1DY2EndBi
/E7XpM/Ll96BmZkVZh/Xkz1JT+1imgR2/lrfNIiK0P/4PWs7FTW9Z1a93TFi
VYbtciTPA1tOHX+gSMku85Zr/HPq3YzAntag7IMwc1E5PIa1llTNpsErDrIN
2kaPMCuhgheWNm+URuuvYhm+KnGKunj6o1vQ0ygQbjMYfF+0GEomNKs5H+LU
rAcvWzF6mBqAT9aXQErpqSP6IlS7jVD1V8okgkqS0DwEJV3P+bm6I+mwao4W
sfoHrWn4Rf3G/C7aSa6URkLnVROLae3qk+8R3lm2Q4EvpKSMiLknPCr9FiRI
0kAG8sRV7Z1IWa3eR4nfhGlCQPuLL3EVw218M1c52CgWpwjiNdoyzXlK/63e
Onp3KWbwFGjBNjJ99M0pCXxWF8RBTdHCizEGGK6Re5ge6EZuOkET0NDq1NqF
gYGVhVODUkbBgvl0tVYkiIJss1nfDjs4Uvrb8wFH0zGppIFRSMBmwNiXn7hf
7Po22SGHid6DuFJFqTlGJvxz8q33xTFbFlimbh3etC+tqZ6DAw71Ky82SWxU
DqrUYSnSYksjEE2yUWZZ9GE3ucxXRTPQ5MOPuYPUtr9Ws8rJlxjSkflSU9r8
k6M2JJ+5oDVU2ftQWNfJoFz9CURjm3L2mnWRc69kBcL12Xl8PeUMPR/35n2N
jKulYGKjVVV0IkRmyrFa5n32jL9ON3n0ZFxl4MGlvrL4CF7pqFdmoWE9a2dp
8uB3hC3n5LbWgYDQPQqyCnHIrfjlrDA5PwbRwPDjC1uqAz/iRr/D9bKAci56
Dj4BfY8yuWQH7Xww8bm1Wo/SSuPrhr3Hg3ixqB9Jdj+QMmSK2KnyEpODi98v
nnxiJRYONM/sz3jJMFwqyLhue3qZnXJkvZnBaoY4L3tuwXfEDCkI1LcwL7mZ
tTn2LwM80dGmXqYYWtXl0QGPSwJVbggdh5R1SaZ+/NzIH/AoXrFFoiKlqDZU
wVeHjmvLrUQgXex2CZwuh6nflGXwANDkX5SNhj81xEEzqQBkbMgP7XMYNaBy
CfO1aqf3MMPDqwelrH6RAPZKob/kOSPN1wMFsIJfOC3/yTbc8XU9C+4HkcZo
OlKhZs57dsO2FXotYxQHIyWmi3G6QGyi5tSaW154NWyqOiFaanMhLCBTFnqC
oKEq3kVSbbzgPA8/84YQ1Qg3T4YPY0alUa1wtT/W6LJMhnXppYO5dsDHcX44
S1smjty3AyBSx5SRC68wEg8YGsEXForlgciWVLZSTk+yYR6kyVoBF1b/Cjeb
WvVX5k23Q72aDxrzlKSEIHHv5oCrmYaQKkK66e9Y04A2EcjazsZ5fEos5shz
L2dZUNDQwD3znBhK3YLKC5fcs+vX5HNTo68SlcVVrjDhg9Tw4Mzoz7GAOQFE
QmoHno9RTF3I84b/gxqxGKRkXn00lwyv3jwivSXlKEvECdv3ZLjZRuSLLJPq
pVdjM2v5kmhUgXAeyFEJs1quaj20jRzq0G2yVlJxj5pdHJqKvOE2RkrKAHIJ
eLjTfiPF1T6WlL059OygaxFHHPdgLVlIvs0hB1jLOAIhpiw62+VrS/ww6Lmt
N4bFCgP0uNlobHxDx79lUOvNkYsINS8eLrgm97rQ7zqV3sAYxO+jY+6bj8Hz
WWFABMZI9mad0d2/mN16jjjv8088UZwYSM/+PnS7B6kqVuVb0x7EyZcn3IYv
+je+86GHL9SwQ2V3751zqzuSqgbTEeRHwagm57WHY4AcjXXezv1PUHgUhVx2
/muoSrwlyDOXialTjjUO3gB7F8KptgiIf0QvYUzojrbAoCP9+eNlwhDx6wqq
WsIdWjeZ6n7LT2g2CFnYBCy+cZbzwXa6sSQtk3IDe2z1MXsBSShBACZx/GQE
6gtzIWAUjctvOxrs8iCtFb57QIV4qi7LZgnPo4e1WBrPOtL93T1VKLD5ztah
rKfRqiZOJAnVrFtSK3NCvrfD3AirzBjxeeFDovkiWqHDMhaV+uiluVrHXLCs
ozLmh3R4ksA2WPCIIKyMe8vMm0U/sVSrUV7kGzwnl6lhvjYxqgeifSkGompY
x83G/qDz+Dl4xa7ySKXvWD5li2W/IKLouLJ0JKBKzQ1a25+2zSFwohDtHY83
hPD4ryZbzpKmAu4T0mQZRCX1LCMn9jCE1RbeXpj9MuWknWvWvntNDCfnFYCo
g2hu+7O7ZRweGN0cno9DHg6cu3Tt7RsdE4ze3JDJdAu+RM0Csq5oaq3JMShm
pe1EbQXONsgryFRvpZrmoucVmgmSUHMmbx6PfTaTanDDdII5uY9N691pbKm/
Ezff8XMiYCM89iJIjdUdArk7OSzQ4I+FcftqtbJ//HK4j5/jkxPLwpB9Aezf
hvA/y9xSEsQOY5hQqUjBFbIP+XpskwyPgvRMn3X5bT8oX9E8EyDNyZul8K1T
KTf2fFa68hT7d8tF0Wc31EHz9wwQxEfswjizut4rTk72JIonmSnigj2pEaxN
E18LQyztAA1j08B/dHXYP66g7FzWrl+x23UOAP2gIy/I8WkiRE33FzGS/g7C
op10Rmw/9RHq0//gCibmfE/hmHYfxE1Reayr5Qdv/i95Clkt7ugKu0aY6YtG
R0HOLQPjIH+R6jZpIzG7cHuGaLmMTt7Bxnii7FsMApbeX8HsKbr8rUJAzax1
W6/RpegIpreHuR9KXX20l1rd5/EgDWs5tlWuPqmjWoJIkGLeZvo4IDBB216N
lz8YSZGNVySJR+4pxIQkQJU8hy1LtqjcGtnU2VU3r9dSeJ1eutGvfk3pr0Wc
IJQKI7cAlBRk6dPu9h3j6j2krJMv0CLfOiyV7HLtcatcWTP2GitFvDlIobdw
subALn8rFiINqCO/TK7k69dq3+KmQnUv8OBd2KeXJc/qPIZvCyxRF6LX9jIv
O/3ccf7XwMco2aCI7GSWI/OM+ekeTjrNwn+TkjsvFSZ1gi2SBRcxhCw0XJft
x8Oz6qY3+TFw8mK+KIxvjYGr3DmrqCRvHpMzraTJ4nVQtyivj873CjemkD1l
mnUxDAHOpLzWsqQEwW4L1fTpVJtpnqomefWVzSYUqH9dt4xsWW85G6NPBV3U
dophnAUq6xWwl9nHzST4T1dg28g0kz03JmGWrmfG7BtttXRCurCXPmzmR4U9
3aOvFIxPOhFAF1eY0OGAS6FCfOsLKhyPZ8Uv2ZHvT46jOW4i2AQkCA+K9l03
VUT8lST5ZI+9uyVrkpZ3dE7i5Hg8w8wcdKaJXyyv5DOC+kRHXeH1zFv6SGkk
TaFV1LERrrA9a0G5MZFdSawzjxZmcqucThIe/Y2iRSqAFGH66xrWzMjXzWdv
Kxqu4xaHU/AWjVYvp3WdhA+gGLan62ZjtkuUnOYJVGYYNhjGFnLgOU3xrgST
zj19bxgUqM6fQIvVHpndHh2h3f1r+F3ewmZye+uJJ4hSodUTGP1fI5FVRPSk
pfbhoW2lB6FgP9oKmEjD5beaYmbh/Ej7lSzXrmCObMlavTYPg1GtXFKn8+Fj
I5rnhZDUBd/CmX9mFAdd3PYMPEAM0OKprFGtdhBMqZm02NzjncFfXi3b2q/Z
JXgwqVtKPq2dNh8btcN1HYBx9Srp3oWimoAhc4PucU9HtrA+SUk5zwrbrC0S
W17fDWBf+D479khlwIW5PW6QU+zl1ydRvPTxhM0HFjbXi6xZlfTfnJA0zyLJ
PBm1i+nfi6xFR+7X6uqYb8K6stSeXM3gf0qGrNJZWUuRxciwghJmH/08kyDJ
ib0xmRriCgyoO1oBG+mMVvcnofuROFuCZvYb8OiOzX0kK36YtaU0Xr43/gXQ
qJVJwDdzxRhp61atlv+PeAB+3mecY6/2E2WvqWp7BCuDSD0Y3K/sDNBf6TSL
QtiNfyj04G5ZQy8YciYrK+HPPmgDSeyjEAp3w8bEdR5Eb/Ka5SQG44HUUxlj
n6CK7oQS2Zuz2eVqi2HjZ4Ul07gviiocsjBrxLSuIOgubGMYLjtzgNc7tEKF
yROtnmgldPtFUGzVAVclWw4kTRgIt1oRUIh8DzDw+ks8G+CzzlGExfdSk8Xv
M02wJB+PxMDwHavKjRDurZ5OQwnBtsANxCi6qisxZZm0tHCDyKzgfWLpMv2H
mJTL9zRCGUxfj/6XOTqS8TEyXXI/TK60ibVn5lWTFQiQ67QbWBFY/WgEvcqm
7Z064bx0PYcSdLI6UlW+b5+ISIi5HGABOLN2tR7H3De/O4INPEO8M/Y2AiwA
1r9J0hcRj5yizKEOyn8uVVjpmYzbu3MGSCGzyC5YGQftoOdfbzbs+JMCk8k4
F5Mld5AqdBYkgtQoYR35eyv2ZdlE3PzmdHPwIqZlykUSkn3a9qR29r1/ZdKX
LJ3Fcg/iNitWDCl97dc6YuvQysPJ4KOeLLSSAeqJYa0b1L222QkQCmbZkaCK
wQV6+xpyicasZCYucCCUDY3IQdVw9ZLLp845B7QizoC2cBYtL2OkzaSwJqtI
LwwBwlY1eZk9ZevqFSccao6qEy89bfryegsyuGn388WFQBy1XtGeuTeWFFSq
cweSbXbZqapcuuWXfc70dT009KiD0am3O4DFOF91G1c5cHHAlt3e/qDRbozP
NDVDJLbb+jPI8zdiujzB5KOct1NMF95suu0Pz4Oo7nKXsK/V9jhPrfdyycM7
JCpVO81WtywppfcotSqvOoSCIc9kf3gmXZuhSOaRGxz8c02wQrS+YG4w/0Q6
4WMR0VB9PMesdUWZqSTirlUUMm4F2PMBipXGNrOqA4pqBdxqrxxoA6Ow6HKF
OwCXQOeFLxssNHnhRkJWSJ5N6vgLDC1H4V4dc8AqfxXgdxN4x/o3Ot0LclSW
VolVmlx8WuhQsgZz7uC8mVCDUFMOcnqnsP/ysaLq8AkMEnEYp3pft+N5L/OG
DcBrrsSdVRXsGzdmBh6LK4DE0opRUQoKIhTYIKlUbMv6XBPV8x29DviKYZrS
kWNDhDxIuYruQQhiuMV3M9Hq6JDAWB38UnFo8OfDsC7MwOEluG5dHH//GLHo
iOrPxJnqc1bPWApCibRBzP+qqKApx7xzbWo2S1AcKLJATRgxqPPD/Tvx66iQ
zY4qmrkNX39AxYPlvysIqQ/QjyTjK8bFKwcgGX0+BJKvYQ3hbeaouYR8jzlc
ZoVNLE7YVpG+Z7EnYQdcOa0PMCKI1zobiRhUipWfm3RsDbIJHC3IpkyYh7Fc
1JwSMGNvN1eu5KQsw0eNwBdtMbprrFW9KwVPpIKGU2FsWc2EJUiyjgnoewVa
xBTY8ZuK54TJOX9VpbNiv3twNqk/UqgsZ8HgaRHNPuaxZvyoctQRi6XA4uOt
i16YFYimVvAFr6WrwUF7hEG1z9qecxh+WRTPYj+NOU1D0WAn0I5ujmdafT1Z
g9jGRpLZrPi65/YyrC3pzOm5DrZUCirx0NHPMhAWoLLDN1upBX7P/yCUGGV0
vi/V4/KDG+tH7YjuPY7BReLeQruGVrDY1CX1PZxJX0SHDlzecNqmagdOAcSN
3Nr6a9GF6XyRtLsxc/7F9DpowvIQKFXz5wyDO/19YxdINzWb6Dc/onRR9nMl
y+RWFZ54J+aGzr/7fr6ZJABqfdIa6sjtH2z5kbqfa8Y1d5Yb610xAhCGpw0n
KAKwgL4qdWWs37zGfbeAbamBPW8uT+C06ROQYRRS7HOPOTmmye2ddJanEdxj
v+LbPMi76ADZyB4ToW4bwVreCdl9msFYA4m+LLjzNfl4H5jDifSy8GcjcoAI
D18I39lzmth7BcseypOReK8PLbXQCPf+QihbSIjhKk8jF5nTbAgwho2XJa9m
r12xiPEL0ighQWsSYD/N0TcalY/LJy9hoLDgvfQjXlus/aUvYsYO6s+SMQTC
6aldMhsPXZDE+0UcyQmPsYL6g3peE3Oa9B+rrRxCSVRm7xBUEIQfv5tgTbAW
wFznYcVf5ULiOBnQeJZtgkU4ovCfwDVG6L7jR546Fz9HWVMl4IYVW5vkl6Q+
8gPJ4PfBMbhJzzDfGBvQr6c+1defeA3kZC+CCef2573icZ7zfqR2/nI9gnf6
5XqsWaPJqgjAWfogwY/rSUVb9Qw/xfdFA08isopvo0IIMjyzX+Vrb2wmbih9
HK99wN43BQZFnhvL7ffMwGsc5rEivZv9cxL37IPdLE1hz2gAd0uEIR038eRD
tRDL9hcnk4ZgzGoTexIBKBh2Kvm2pRNk35niTnSFxkhFgvcqcAIhZm35s3pX
qncG0zAhqFc0xmDln/Ll6Txg+BnNCgTJQF1TY9yOPJMltMrlMM07Kbu1lMTU
chDKbzfdY16mAWOfarBbJoJFwDkJ1KBUC8YyMRDUYKHk+XT5oG4dN3xBkXHd
44NJRLL9MT0NEQcINSERXYSRMrrLjkuRt2/VVpfmFayH8Q106LzKv9JgHH/3
stZP70PtAaogyKhWFuj59lKNN6Jg8ZD8MkL6sqBGZ7e2egCyN3awMYAcJJR0
p56pj3HyZQXlJXMkVqcvb7Y6A49VR+t+ZzNA3wGnyHz6vs8p4+JeGodcxreC
qwx3afJFcJb4DYOn4jyRr6pWjhyusCXBbj9E40TDlGdPm/l/iREpHdM4Ciwm
1YdlFq2HFPQ2HHBEOEqPH14cr8iaiWZvkSOmwsFRMC6xrLVLP3ohbcJ0+BnA
oJHPZrTQOFoYPExbqQ4bmPvAqQyAF8i/OQ/JZJWTzyNDEUl4a87PL/hg1tjN
sj8f9alrqYBZzxoUZcfrdEXA9m/y/nBJoG5xfc3leM3Ul2Uhql5DQ8uD6eYz
ZhipNVdMhND1VBiSsMIOG8BlU4zpF7LAv1NYSCyFmESCFPhv+vnQwhXy3KL8
386l4yIa5lCG7mmM6D+zbB8lYr/etgeW8z+XlUoqsJemrrtV/UiE06wkMidG
jCgmFhe2Dtghm1vtYtkq/przq8QFRVDx1CsBwSAz5tKE8oubZaRh7lKk3Pee
gtxID4FTeOsn8h2n3q4J0GNFADSYlFi3WJNwZjbMwpCCOwpD5I/efMhaWqgh
iIg1uWvoAj8maLh83qNE3GU+7s1VKVmjEIk1aA7dpUMJqvaGL0Tk8XKpN6HH
BYu/YhjIiVPXfxtRizozUKaoseNYmbRCnwSCNLuFvg4E+FgP2V2iFJpae9G8
9g3uBU7ryx2Mp/xqT68eVwjqHoF+XuRiIJUqwM1X7Iu4pItl10mxhX1bYupn
NITkQK1VUOnfuXaAu02m6Wo6N3BNplWdkkvWJNoJT8Rs+49XtXT4+PATIbd4
GzmXlbmgXdq5lKuh/U8X3FT2URB2FOEdGknuTcZj7mhFhXaAdD1OJo7AzVM6
oQVoHEwYGvJHwBJ+dGCMcw3GD0Zsw8PrXN/6gn5V6KbJAO6upZVvtdjlVMvM
2lJH1ydWJ0klVij256QC2EgKXisNxWQ9W5FuGtwouLfmmS5Ze1POvXRXXRM3
P617b+/VXIzUgvcM0e7nIDY121lZfWXqnGRQHDtOElMMu1Xst27rU1JXdbOR
huZvhbcSqIYt/D94CIi6iwJ7c6qrODw5nVErQilk/5kOLUKp8fp/fUna3D5M
sHOaX+JGcUCjyF3vKOYrN83vniKXacJejjugY2MQhHf0CUHx/g+pgvnR/JoG
67XI5J45AIcdbn5wY4G9oyNMsa2GeojKh2u4gOw+cYnv0/IMQ8FXsscBT92f
a6aWpHHxNvEEx7+UFFBII8sPkKsUK9ik1Lyhxvx2BMI86/VR9TRPo5gy/RS+
KrRvL0x/o522/yQ5w6LfVOF9ztqYcd23DJcabSfEsX9ZtzCxuhDaWM0Z0RSg
T/Tklx4K6+L5X2wO1BayNzHeQpI9ZOZjb+8jECp/XG6yPn4IX8y7w78ew1XW
Q5de+4SrkzBeWYOFK9Vz2Yys5BL2rfGb8DmZn8Nyu8mOQHN76izOIMmsrUQF
qdAF5vUi0RigN3dQK3pD9kN6pAKr+21plcNWWgc+Ca8fYTTyt1vFMM7rry8x
nqo0+zVGsXWGM/4cI9KZ2kIAtnWDEBcGaCgAWVYBv+WnESjRAJqOtmdyu6pV
GyoN1OHsXhG6En+4ZE7xkL6LOkG/W/Ae5ojyUwbaGC62OgEg8hbVaeLltNNF
Frpyr4REcGYzMplj8zE+yVh/OvVMQ7zgp5Nlt28L5E6pKSHU116J/8gamq0/
/RCJkzGJMR6c7wLoJi8r5+iz5NJ7kXk+drh0PmziKDPsf/I594PE9elc5SmS
OolEoWw7dnCbqd/rCegk3vZhKLkRVCEC7X/bbUbZmafwFx/jjSpRrzO9KDPr
boi9xtHHoGTCq+UCdiZE35zANO2x9Pk6zHgSRmUdcVQfOPX0g8/SeqNpsRve
3LD/GyFO5v/bpkXihlK6wwNrSliuKmxXmwCnbg8iEKJN/+B3aupKBSLw5Sky
Us83R25kyxbYCdCe2lk5hAch+9XD+TESzAU3PL1qaNznTJOZ20eaLOV9kuyv
zcz98yu4VvM5EJ+oKaQEpDQhpJePEV1JCbIE5qHj4ayxBwTAIo5IpA9Q0OKs
8QOv/7iggTt0IIRp7ETWmB+Ad4mWTb44E9ratsKh5k4VvJQYSwDRFFV/GbzV
z7dUkrK+ahVoVSPAiwxKlsEEMqVtjA2KJxHp9XvU6ezKDb8Gj5MGAUsdS+EF
0Lt3ozu8tDOIvEw0z5gKlJdLH5UYbGn5VK49931eMInQScwXYznOHgZoDPtO
Y7bxWkFOZniRE6K/4NZIuv/joNQCzGCKRkIry66KhGjaJJdn9niEul9xmMDv
L5RZW9q62DLCPHGkZNE8HNSuM/AxXPbWCkGSG0wdboQYCKVH1Mngpdg6d9An
jnokllhBNJ4/bk1cWdyFaBn9o2giUGcJ3/9M2cIwrPDtySZOTdUlVvKdS1A9
YAlTyCtuWnJcmKows2eFWgxhm5RZeIlkP9aO90z7iWWsusRfUn7XztldvEja
hwfF4GCwVNF8Z4RB1ZjVH2Wrtrk9FNd/05eOO8qPHvsXsoNJL3EyX4LdUPlQ
vudL8BCnwMz8DmCFgS8rp9dlwUYwoWdeJ0E9KdlSGIH9DX2w3tF7x47zX53O
BDl8hiFesZXhiIarBwFxbllukSBv+0389xRZNZmKK6U4s2EN80i4eDZUc06+
5AEOkyRc2DxujLFXnlGXoci2+rdCjCFxO9BW5XmJATIz1q0RA4NZ4PGSEFcg
0mVZ/dQuamZZ9nkLfXqvIlVZLUbd8d/GFkU+tFuSEHs8iJZWdSPEEGgUNaXa
jwnhKRFcKTtx5fzbgThZZbr/RpBrE9ooml6ZSd2jIvHPmpqshRFvyWclSJUN
cBR4eNGormY5JOfZhU+dt7/BSOPZNgpV/cvOa6zJl9uiJYUerSWc8Z6nfv/W
h34lES8bp+RoR3jgFFYpxnNJI9XcTyZpesXsTcTP1XLLxTn8W2HiuaqQddKW
Z9Bp9TzxW2agwPVQC4NHS/yhEOOkKYI/LW4+MI54Kqyql/XXpm6xcmZkVsr2
n7k2Um3VMg1VgXl2llitXkkQDvido+OY0A1aSSJhlsggND3drkaDr7k/uRqB
XG2TqeVu8JjKo3/b69YAIpg7qig+dQupt4Lqxomcmylnmvq/nE15jVMO09Y9
2aeNCXDNN2eskFpJ3g08p8awSt6C4fe59o8VXlrzsOMuYpgJi2OulI3BTHS/
XDQEOGnrAwE8RSuYDqWHTnEnM1bqIpcNkUuW/smfzsn7nAeNNY/EyhS67OTd
Ae/5DEwA3zpi/XMWY6hhiN3vBxvKSImKunJDjkwlQJ19EFqKKXEUuK/rLMin
4/+WKbokvLY/em06+gL6qSQIADFVgLY2BN8nZU+i4oc9XINLHpSCvBubMJ1K
0Wp75Iqyv/tZqFRUtPl/ymrOrzMSV77Era0DNOyGwKSatJlIpeWBnMD90aOd
MVRutV81ZKxYvKz6nrz1vuvPUJyHrzw6g1ONd7F/YLd8MDi8BCtDDzq5KF35
WE2EltNHCYCZoXv+328FPTn+qVQW4Pk9Ze450oSAee4JT0CH1qzxRwKVoSrj
vmnrGPZ2Xf8/ClH8lWazUyqQuuuXQlcloNCVKDOXiwfe6Lish6WdWw335qHY
AJTY9EfcOlcU3ov4oKtIftVFQD+FjxahDipvjW1foRYW2Xnhz6k1n1jAVT5E
KVC0BBuZGysgrLqY4xEDLpqf2ETQQwR65VQV9KhEdmWMerG5QuKGLPsq+vkQ
AnSRxql8h4wTla6auQ1pvfVq9t7Wk2nfEn31s6Jbxk+wftmt64cxx8dWWtv3
yv6OSiB/7eI7vcelUb1O3pjFTbWAIUhh2Hr4cGIFpJGQSfnt+A1pnHNXSumF
qeKiKX4e/uiCj5fgnZCKFIZON2Mijdea+yi+x8clO7PKqckBdz7tmpKJLhuP
9vDmcrL75HNkYAQtvZkfLVpsA+4aYsgSpl2glSBMjW1TsCdTc5lovrT3TEf/
3O19SkhRU4JqOxT5iQ4Av0DDVXeDmhwKI8lfY7l4z+ve25/sjB1XPngDuAB0
Kfk0PemE+xaBPhQassf6NutdKLECgIt8ISYeyP4xJcCgNbv+lNksLyUhZZkF
ii6tBid1nQx7RTR7LVHE7j66yzEru+8fyZoBrlAmXqL6Ol/tAMkUZA3FV83g
H6F4THhDGVKqm+0GRH3FAgW3mXESYcscE5lJfuAa1daUovOmxhQ8x7ItQCrJ
C6Pgm8F+E44AlUnykjC4p8rda+xlav/H4XTliYQBhTnuDUoAjoR8rIIXpEId
AnG2aywGl2SJVmNPcbr0DKhxpHe/dDj6S5A7rPgEzLQK2cAZx5NyJHtyfEOk
hFMxsw+KYkTUi9DNYuxrExECXCyY3AQjCSreQ8O3Hn4fRuVMhNxLE0PScump
UlQpef46gMjH3G7yo7U73qn8dzyp6BIJyaMABKCqN97Uoa219zGM8gsNU9U2
ooLVd+grBBrOUzQVOF79NkunCF00DRl2Cem2F+1dxlYMjEdapvsz7h9UZ4Vw
pJnwzH6lGcJTq0gDCevmxQPvQei/aur+ckVcZZlK07YtChlHJIxLndo7QfBa
CGQa+EKELA5Bu19JKApwAUNBLyLeNF54uEOkKleWMA65qF5dAEuvL+HUVlyz
EGHYXwVc8jQb3YD7uaZl26edt3nlQI2WfYbDr5W9X7JdNWA4t3JkE5BECPH8
bN01aiaDd8SyrEMwn/mlcrrhIh0m/PKKemtkBL7OQa9GKWBlRdyyXxwYvmUE
pDeE/qWGOQU2SVBt/fx76NgAEBzqiP7XVQTZHcU0E6XmkZqMfEfHSiVddH0g
eJJqKCMYdvYEbUXcVhSAzV5B7PRhjFJjpWkj7f7CO0OEk0AGgZII/+wbz9pX
HK6tj7OBpaJyKf+zNbDAVe32b7msdtyN7qWQahGY2Zz0AIESBGNfZ+Z6PBlE
XlmScbfjEn+wu8bLWxliEKTwoVbJTFBuUcndt7LNDhBvkX06MCeU8d3Zj3Ve
EWiPFdylCGDgMQfCu6kY+3V/wI6oeTwaS+FP0grqeDGtDi9pszjrtmgjh7hm
24whAyb7DRUIoL+jBMhtFxitCtXCAJAFHhgvLG96NQMWD0KkTA/x+rBwx7LO
7k9Y45rBJF4Z2saCTH4i5VWe6YEOjLtzUPkyIeYpXv16mrfyeyIyog45n+91
sGNnMwN9gNsKCsR84PAeJhr86TUbVl6XvbWT4qvbSlYywIISh0Kk108RnzAg
ZnrwQjAsfwsdwjb8RaaN4ooMMDl57C99aQrpTiW7odHKX4mnyBVFp4tsxonK
3q/oQHsxdZJh2XT/J1NL1JWzWjemDgJ15nAjptaVT2wqApO1ah7Nvsph9EVM
nzDXJFGXR9/8rQefXt5YDY/a/o03d1LGUzUlA3msFRtcBvCT6Eo+Wo1bVe4q
akWE4mhGHQa6XzG52xtAPAM+Aj4TtsBPPEnUGY0o3pKgM9G5YhwxYe0oSxWi
PHGAokeNq4iTgx/f9GU8FI4SHPRZC5QBP/6j5J4xojm6z9sirBbUVHhl3BS4
OmjGhsdO/015EN2hb4gfWVGPUezuAKjWss8U2ulO8z/z/s4fD565T6qsKNtE
WvIJlnPpFAn62DLRIadhkOylfpUGa6/r5xQb9tEqw5wFNtFy7hHvJLZWtnAY
zIXTMLCI9iEIh328JXc4bdG9SccdvyPY07O3lEKwMg7ASfW3GRIDDMMhQdcS
ROXvSBf6WNw4pzqxhxNv0dIPVgDdQFsTOxbVmtUXU+yrYY3lcQA3GG2v4lUx
8HW7B5YwktPNjAyCmr/t9VxpsR5Ko4sfrTzaHUf7gfA1gBt5w8P9LD6FvW/f
kTeAiqvyG5SHp0ocq0PQBPSydgxlLZlvfxukJ4eN3q3pFHX7JYOTC2RIc9UQ
A2A0d5yAtt0wSDLpoTMgvgGi1YiiFfNWNAugLOIuztFDxqkztbMuSdoBuqZZ
F0prZhSd2/9XpsrISF7oC4rQJhPgB1SJBGLYb8Oh/mH/hOTjQpBRb+EArBfP
KjSST1BkcXxo/O+UuxzcARIXQW9CUwNfLQsrrdPK7FZymHm4T+TAM6Ish65o
U2JmRs2WUJlDh0/77XDLiGlPv6Gf1J3U1kZ1pB5s3QN5vcfxFwXWk3xRWh1a
ga9KH9t7LY6Gs7kY0nRWsrjwNEMry1JhH1PPtk2i9wxwFMZD1o7mu03JlVFM
JGcRoMQyC+AivgdVOwqKBFKFql95BCb41UO8DhOgsLfofj6ilXVvUdFKvQXT
Gg15I7U2nVQmfsoe8NknIF8iNfkhCCJKUTpNncIqNBpsKIX7v8xRIqwSpwXl
he+3v22Owb9HK1R1NQ+FzZRC0blswZqy7S09+KKZwhPug5SfrAhg+Z1z8HWu
ZBtr9mDqjiDNEUmsEdbO3uwtOk8r+lCjZUg734jQgK/fF0yHFIrbc6kgVj4A
pq3zxEeTQURtwL+TRwvH1zrCW4VQhOV7vQGR/kbdWBUIs8C125Yr0ZwicT0c
UpszL3OfurCBz+q/tR3g4ByVAb0JAHEhN/HIFcFEJTplXJIJ/3iBHzpE4QA4
QYI1qx4PXavjLHd91xyRKPcnYFeDqXCe+NIQ9r7Pu0lL674BSD2iKaN2XpaF
ILLlkadqI2LeDGHjY8JvIbO9uZF1o1LVUzoR1c7pzbLZyWMMzq8DHQVLzXpD
2HL4KLAIe1jMvGKbYPcLVyhV8zgSnL6Ma7v/Uy65Mg5MYngEwu9YHOQjA4je
YJXBYme+6T1kjisXKDtXqwGQ8m63oGMzdjRUI+censxa7UstUGEg9JNBdVUK
3aFxHf3WT0aUS7jRkPhS1SfivGk5iABGSS5AZKtcAgVdwoJExYUNviVqlrFn
2tVD0C8LZokSg15n7X8E1cb6nsbed6T0MZeBhMEl20UP410b3RorKoh1j3S0
EQsNFTXd/Bke/XhPZ8rxMMVjEbPUdvggPOxgesuZKN6kFhUWxJRL5HZeq7nd
hhTCQhC6g+IMveTDcF5q5tyW0d/1/pO4z+ZukwnNcK7uJKxkan1G/pPMxl6V
6KBmZoiUpoevwC3eRycU0d1T0IhiH85rBJYocMAwggIYf1FxfCtNDChRtvE4
8GB4CA3K9EO+NEW7KENk6WcDwq6zfHEicXPudaKNtv5l0YQ0ZflCxK7Qp1RG
JjUgBSrMB9Dyh4qLOD0SNmGzvtj6SMaUnuA4CA7BQ2W06SDKdzIqjjrdbprN
bS1CnYhAKKJcmdcPyuJ8nxauVlJDkdUT8SxmdL1A+Cy/8ZAFRXxdsIa3VKRi
POfimk0K0r+tfC4AZY/18Q4EhgHIA97hRSshwTWdannYackJZuGKrMAdouFh
vtqBoYJCL0NaxdmNnG2utz0UKQWm/FG4mpevqF+tt2YP5yHpZCwEPdY6MeYh
Ak16y9aUVlFagiWHUnx08l3EUNkBlMKBnaJyvYOZTJt+EZYR/dAwMNpb/VJf
6AQW1DfuMpNqTrIUnn3rbUlPG8cRb5Ap/TfMOcfQovl4qr3SIZx0uQfctXLP
Nye8576dfpeaFG8ZgnvaZxmXFr12H6BD7eW+qt8tgmOPKuLdgLLClDo0TLTL
OrOzHDXYgbIxHlNo7FUKz654rWLaTB5dxrDorOujdbhlO3xyNvLscvXDQqOH
G0H5fV4Gl8v4Edft6vJsFO8Wm5CdrNYzsQAvT+LR4no4N1frxUgmW+f7RonO
ahVWQHobjc2mzM9D7KoIGRiyzcJlBvj88yafCbQ301siA8wcReaB9y1CFzGH
uAUAoA0+tbGfu4Q5pw5n3UK4vl8g6y+p+NBePfhzi+9nRwROsVoFi8aeZsK5
F7sghr7Ok+Gp6VBso5bs7d+eciUN9W/SICEuDsii7LqeZ97j+Nr3nGmzxU6E
Eb1yY0rh66rR//IYbCb0VlN7b6W8wuWJq7ZMCF5UwwJSgj2c31Q45Jwim0SU
6hzNd/PfIlMsdWuMSKTHlKxE76U6b3BuviAK4ZBmipVzzYpIR2Yabjv94Dwc
DxEeBm38G/ZXXRCfKM96SP2L5nK4I0z1mn2GsUR1HxHm9T3Hr3eprOB2ueGF
NYtmJsDkBaI3UrPabBysRpHM3384q9lDWvJUH1dP6gpEGLCvOQEVb+TwHYHJ
PaN6QyjgdlEG/WEpPR/0ILHs8sQblu8z4iDGDuKPoiJeyXah+1OMh6MTfnHW
jeZdtzEQqQe8XOMwxyxSOa8rt5nG2mNRlLl2rbaPlLL+2cdO0Wc8AL0lBpj4
Qf87RE2s4STHmaWyTiP+FLYJOaBg6EM7JZrqMcQxZO3ekNOyiE1C2GvKSeFi
ESJA07I7kpovuTw4fjwy7sG+MwGIyZU9+FF5Icjm2PSNUX7b9bMR9aCdk2wx
Y5iuc/s8kAZIf0YpyAF/MCRoW/3LPTyn20Zl54igABkhjA8wPnbyKbXtWgr5
mHo+9ZbXb7kwvCcHt7btE7I3TD/L5eIlFJQw1z6amiAQcJaOKngfRe9E/qlp
VMR60+txzf4PVH58TOHc7U2Fp8f8ELmQ/f0u7XmWKdigAISNXbqm4Zo1ahjj
7TerTdRJlkG9wlTtMnRTXEp1EyHaTL50WyAE16Yj/KSuFSsaWWkSQp7Hl5/Q
4Qx/JhZb/ReYyXiZVRk5kvt7PKM5IxbGn0VSSrPz7E159YwlGB/xyhyQt1zp
vVK1IR1eyKCDyjunRlCJY/UuqtOsElDc79jwR0UhdNPdazoEkSr9i00G4261
0f4AbDn1o8yPPVlthKXF90A0EMzNkIJzxiYGjQz5gRbnbIKq5TGucZGyEDpt
z73PFLyB2lwwVqAmz4GFpn1apMiXf1yifNGEtrYxiAHcaNIlzoB9VRxsb1G8
WeS5V6glL7nT0WK7jIOYO0X4kekLIOnN//P9lkYlyC0ybvwIlQlqwbHB9QwW
ZKqLS+NrVfmvPxyVKc9MFhaDowEDzvlqNMJgSIg/zGz2AiAPWU0AI/XE+ILI
bsOuGyVGXkq4BdQmY2qIaJqdPHC/qdoZ3IcVpUUmNgHRtdMYtqXHjY4y1LCE
C5MHojeiai/+Ufa/B3BNcSawZQYjwlflWu8b/qcvAw5C/Zlh+TcuaRc0jWJT
tytDJvjo4LzJxKqwMgAkWigSSgCzA1th1PWZPo6dpd48223syGT9xJGhvHpf
2mwVG0KHxNqtfmhI9fcQXcIgipMghKzoJsnoUX4Q0f/obFlZ4kIAoB7ixnO5
77ctlH0ovGC4Y/2/A7bGUMg6z12aRrBhN/o9RebHEJSuyHQFUdNQzrugiLSt
5BXgBUUWVYdq7RdyAxafp5YtiyRMZXtyKIucbh7/ij6H29RihADaX/o4j86e
lKjI++kRANjCs2Z0cBU+3EPYSiQ5tmA4eOQB2YELsWddxxai7rcVc4RfZwpI
cPlyphOPidawrx11B7HRAvT5SXCNF9neJHaxtvCzeQ3v5mRPIL4zrow3lKF+
Ka47OnxWsiRm864nA1yXngBafIL7qxg7oEefRC6sT5oHNjCbwbWquAMSUphd
jWJvoM68tz2cZ4Eo7u0WuY7rMKDUZuNLQTjG5LdPz8azMTeQV6hMp4VMKSN4
uV3+6MiyMDa8hRZup08wIADZK6SMMlquvDaPpNizKD1lZzG9FBPwgSXijf/Z
1aFupZKbOwv4jut8+UB6TCyuCYf2NFl7TgkDrYCMkzqMyamM4hu7RLG1O2ZF
JKY/Dm1/BrOq5xuyJUs8sCczRW9EwjIS4yhVrxOrlhGrL2MQMQVZiOAMM+ne
D0fnmo6WBddhhb2+P1UhULYKXnJNk+r70DcauR7cAUGeyYGenhvNq7e28mXc
LWCiz4xB91keal2Z/1k4K2ejxXlibtdUd4vjMe1RDOzV9/gYOCObDVbeKcza
gy5cb7bwSLXGh/4ha36m3oe4C+i0gf5CMLBMxMwsLyjGpCJzaI3Xj+tI4dr6
LJZRLpQYq2Y8hiMO27bMCN0Yg/gjF3Mu999Sv5xqMbP1mgNxKsbuEsYtIBi4
wF7R+PxH3iaCoEt6GZevLhzvnWKlyegR5vBh1aYKZONwK9fUEGLu69tZvX75
alZMkqwV7o4HSW6qzdTXvu/fqR1GSSZ8zVXoclXRLe8VyDeWZdej1Ti2kw0+
3GgzccNUUuVTd7LL068LxrhZN56dAbn1D/QineJS5fYKdsb2f1+y/gX8J9NH
MJcWefrePFEJE7utwxE+yQuZ7h9XKjMoQEZ2e8ALnOWhKuMRZQtupIsBghbE
8E4t1bF5bPm2viRN3rCJwPlG56T0s1lhzXOUDhhWPm67u1IY6lrtj+a2Ts0b
9Ug8nlPgiJIe1vRP1R6RsZN0D3gAcCVpXRhfc9HTnzZoU04P39q9V850oqQA
LsYbYMdaePu2J8IWD1vmgeY2qCj3gj0AJLoYtpwixAuGZDmD3rELsoJEP1PC
rMd0DUr3GXqY/tfXTBjCRWsVMcmEvKhbPuRsrjYd8SAUtFdvE8xiXjYGPTD1
fJPeISeAKrY9im8u7zZEumm73hj4GmgvOX7rUEtX8wXLCHHutI7B82DIDQX7
o0sf+BA4BrFGMh8+oIL1LjMbosLo7/ZIlzUKHNqkNx4Yjemeh7zE/iczJhit
XRPfrCkARnCDHkbfDgeqvGXefBtBXBc8mMwQPgAg2iS1m3HmB0eKsIC2dnou
YZ1NTYXEZadAXoTs2obASRwTp4mIbzWaZojVkXrB7nJv44SV8BlDzrgHexR5
Rln5JvTlbcrz5UIz6Nbe3Yn5dmyAspDT7tMkwM5QyHedNsdhTgnY3F2Ev7Yz
b0wi/Qn+bKdPU0znXMLw7uTUyBUgGompgw1QJizbuOQ1nMCNkbvXQlNtNzCL
rNOu6IrzG7ZFEYu3kwuMBOW5sTU6fEmncRcEoR8NK+Jm3/LAaV4eG7SdprBq
vUsJtF9PTQQsu5kTyxGE1hr5/LnnaGbhBHNxDUQ7gzT5yxP51ayBOZzNFu7y
pxqTba18FDdE620ejWBd3UaYBv6rDxQlTNuC0xp56Y8BOlglgp2c+zjd6DBw
BKDLREN9t5xke1IJtwGQym3P75lImQQS6OzK1syKTLwdt+wxuRrXnpF1aCc5
Lszfi2wrW9sroBmdHgd++NOaadc0JX5TlxPoWXYoHEVVjIAaXFqIrKXMfOue
hsyj7ufWAGO936TohnG9MxBuwWcNRsngpp51x6w03W8gTd67/zNHPzZTl5Jh
kEI1zSnQjV3JtIQq/q49DHP6DHyRTfHo3OKKTIxHfxfYpNeTLhyf9F2WQWre
kLfAw2aebbjFa162IUMPQ+Ij4bgjMXpJO+zDlZEhSClTbuEXdwdnJWx4Ut6S
8cX34zBdExdgguQC1EP5lo2dxRQ0a3HfORPhps2KN16WXNfUOk0KzUcdsjGI
UGj0C5NxxurxEzrW7QSBJK8rmqJIFfsJZU+dGhF478ABziCeUoStjHjYXmmr
xJU137aYxe4Hu2Ef+8DHTDPsamQ38WSR3QCyySLl63n7MLMoY3CNv1kQO/mO
ppQOmTFj9sZymLVsVgQK2OX5X5YoAzkcwDxNws0iEb2ycsWQL40Oh0eYbvpN
XBYU9IlzJp9afeqj5C1Mrv/Duk62csMxu3v4bfx/wcvyr+qmnPFPZqvZ37+i
yOHuzWNpQLSOoMpPtDEr/FW76j0IDZqoxnb5tS8e9vBqKruIEAZsP8xh9b0F
8Bn01bcqZ3hAdJeMHHDniUn7BAO25bBQO1r0ix1xG15yxDPxmuPSZcvfFOGs
+dune3gbfXnVIQBKV+SV7G0y8pSiJgLBGqnY3KGVLL2llAUln22AMtA23wLl
gMHoyTaOrIXglZcVisca4hrUKs75lABnJrASffNgKZtU3I0JFkRZyNv6DaUv
JLGmh+7WZCSYh/mDanWjlO3SFIoXiYIfcb51NWRr5sH/Tod0ReYE1S/gjX3/
ewaqWP+yYOafEmcZMtEGawe29CWdWgat8/n1lGXtbks75nVz41Y/y3qonyZP
1NvfgIMmQVpbP0kCQ7LtMfEripsbWmLcsMJzXSVCHvYpO/lPWLGut2TOa7EG
SrSjTfOQacARHdPi6c3mJYVZBFtXdRhGHia/GJyJoLGijCmF+enWqkvvP3+p
eB97yErkDYxAH+6D0GsqOE1A/b/RRN8j5agWiHvSdVspfoOnwuapM0ZynZ68
geKLmw/sgA/xVePtfY9/Hho0f2Wy1EKAD5Wkd86yO5jjTXbqJuadjwvmjF6a
5XZNn+nsBriQDrrxHCYMCunxVO/eaDKjEzgPBWe9POE5ne7P1+dZZrqi3wdc
uKgdVTXhqjxAma3LJHSiTn8cUCtRMXoXGcm17zKtPtFSbnqn6+2AXh+PBEjB
5CKayfhFNiebisHNNMm1x4Sx5K1b0LUw1Hc1xwVNPfi2HN7ddGrXfvpP81KM
m1QXofmQuSmIWXuLFaeZg1WGdXkDn7hYrYuVnY2rf4rOtPllV2z1tImZDjA9
nFux3DOqFzPH7Uwt+wQeP6P1WjS62NYRK+pYLVm3dhJD2pooWlacD5acAzv2
nl+o9QtWS5YrLeRIowdMFqIdvET5+xEDFSvRQpMRluWR3E1gW25P//M/IEQ8
nzOwBCQ9fHasOwaoNpxjNwoBK4fD3gZ2CSpZlj6VeyAVAHZEP5LCGDyZ3q+X
FR3Mz3fBh6iba4X8Vn6GDp7+MaOoIB7bG4tupzLUrPQS4LV/eMpwUy8q+RxW
35CRAXMLZdyN5xQBhKLisVwkDVt/QBZ1pONicw3Vtw5igjb4JVDixk2zB3dy
R7QQW9gV7T+ovZUWdtXZnD3nwz2CsDhGn7bUlzEIr1e4LZXl6Mv/DByf4cOv
XJCQO1iyuHD6VGZ6mPk6w8ZgD4rTkqNuuCc59U6tZilMIM//arUlfU+p6tRw
h1HPDCn5vM9ra2y1YnZQtbbqCNEgQ7OxwEZLaHfG3Lm8GHprxTPouTyezQi+
5L/xFpFYGc5S4ZmI8CQMA8Rtzpt4xihER500LEPYZVXgw+NjSBZZgtHXA/11
IqcpuQATvNt2TKeNXW0HwKCBJmP3S7HGimd4Ua+bh5HK1GZYrc+bZU1eQlAc
EAewjociGygEdImDAL8rsQwSGe7Auu/4S9qLce9jcJ2IPAFRPkQHzCGpw9sJ
ENVoB3iZwtSK1KExTIiaKTdBGSbrgREdX09RpXY64n4y/jiMsXPEREz6YmcM
+CwtvAxR38VPMaviw/Vlnvgi/53YYbGxKNJlB9CulRD50a/FFzQ+EiAdflHe
L7lfTenIK2lowMLvwNQZalOhIdjLTCH8zX4pGoZTyuhYthnpVA+nEMjPnqjJ
wOE0AJkDv5hB5ouYwfmpJwGpKQvFft/N+YxkiI3MQa8ek9DPtqN+unp+blw+
DMISB3U7yVIu11VtfpguhWyKY4g3nj/sjWQW3Jjv/jzpeyhR7LWytIaKs3JL
vRK0j2tB6IkodEJcl7kE7HDaKmdR9uTBF1P/hd01nAraEjM1oJ3kKsz7PYym
y5DgytYvtCEXPhPhPnadW5crNr6bIhaLuazpFAJKhlxWh+P2ZkVeN8BcDEPf
tVJoguv/vIjlsRfBf0JyzCN8c1hTwWR5xjwgZIzKi0TQlkNfbC4Z7nWonXNX
BYO6O31DBo5TPYNAZQn5/RfzzpvRLjAs5U28R5rhVFl2dOZnV2OhyNlf6G2A
ftrPl5aGp6xOh/os/c12n/5o+jj41ae89VxPW2IqqZj9juNAXA5LgDxyZZPq
mCjNZf/qu8ywhx6LRBrjSf7/xoR/1U0ibSoGTpGPK7Hzn5de7xWIMyYRBxbG
7CIqRIhdLcdQGLrZHJ4ReAwSD8Hrcav66SkNzYRWtoRQIdROw+sjrqSSV8Xc
pKuJq/gdRkqE/0m2zolwz00KniplJNJo/ldIL9TSaW+hlewtXLForDcFDLrF
U83xBl7L7EWfyQkx7hNrtwlz76wHe/x+YshvZANDhSv9KCHyfg0xproPBdYO
EP8qC4zkz0c+kZR9RfdihukY7HKJkgH7B+rODiIXdfk0i5qF7yZJgHT2kCU9
e6tJDD6+rnT88naaiYTYzGhAP6Lct6l0wuC5oRPn2XQlEXGcowBxz1COejCl
URC1zbPBujTRgoHGsNn5Kafek83ahmd3ucbBP1NE5mjzzMiVKp/i5h8CF3wx
jmm1io4EjMe3VWj46Lo0gyxw7t8CKi0Sbje2NYAqUKOur9bRsElr3WxYKw7n
gN3E2oMpXR0+opzM9mY6ZlFvYkK/V7ru5p2ExCaE2ATmZpzSX0XmMux2/rFK
YzNIca9UFGU7hdxqN63DSMu5Bjyyde1uREi3s9vPKycxaHWmCnT8lGDlCcXX
4/CamMt4cIyxLMzui8HYqM9OuS4skXrJ1VbTdeLjPWes4ffWIc6UIkX3aHY5
PKrNc5DJbxTsd1Il/qbRvJ2c3zH7jg5FqJ8gZ8cw+a9DJwbSUqPPANP0iaeu
cNFVPLI/kxflo6dn1Qi6QwGjSCY1lqZb3hnl+fFyetmglczw+pt81JwCjIQX
olxrcR+vxRYN5hOrnn8Bs4rA2NFyX+EYxnZZFvrtTgHlNZRgvX954t8Q+SvQ
Gu06D9pqgI5FU7SllJqbrOuA/oU8IDZAkDAFRPcAfQHdabbjGqmtq9DFinHG
Me/R6+nX4gb9vd8LZIRoreHNNa6ElvJaQE2MX+RLXiDuJF635OCOl1CM+0JH
SrRjQN+F8ky3lMJ7l4xlO6Vd6m4vFIo0RdnrTz413wBKQapl2a6ZCaobjymb
ZJ13NesAFjl4epNsIuR5BiPfokrc+cAEHZx8B2I5rQafCKgmpVWSuKFU+iRC
mcqzItH67muofF+8AYnNzW/tFu74n27FGV5aoqBAltP7zMfrwN2YGC89tYbv
x5WDtzNQO0af16guOnFp88gAGJ70ZvSUSxdav72tKrygD96BhL+66KuCHtuv
SIL/pqUeEABrQOJjljAN5zT2n+QFb4M0uogvN+Rec8vm9a4k5kAqfMG9neMV
VzejZgnL4wIBOHrMIUMwvbe42gWfsLFMRQ6bRiGaCYcsmE/YnIE+X+wxQsXa
5lF5W/fJR6KUxWc4fzlbjsJTdPFjSoVxzXt8acCcl5m1BHZZXoQ8t2b/THy9
0ocPKJnkfdyR90A9yOzgG8iksl9dRznCNLN0g8ZBkOh0Qm5PbJG8+ALZTKCe
YUqy6KFX2O3gjF6LsXmXzgOXB91HIYhuVCmrrpoPJCFb0L9JVSAmP5M7OKdz
eAeP/EXRj+HaWyUqgRiFKBC7zv9B/XfckhoIZfLEHplpI4+iYfsWlZ003Ox5
32VxyW6Ovlgm36YV3moWCxgpL97qAYYgu3Sm2Bj46KhOHDLfmI2/NWSBH+IO
sgMMDqfvJ5GR/kWiSwnXhcbFjiUB2KmVGnsUP4/iGAwlmm2d8VY9nEQfP5Rh
PXuDeFsk+TRle06ucxcnY+XOMX7LrCQeqYbRIH6OhdYdJkO4hXsXZonj4Tou
PDCMH+9My0Wa7rnf/GqRtk8h4Y3pgfPbaIg5mCdXZsbfbUkeD3wXYKzdnHRp
ACxtThvnhUd5lDhSopUq4pnS6q1pmv0CyNyx6pmwoEsou4OiaMM+96mXacPe
Y1Ixm6vXAmxySsff4qIDLJAtELPMAGDlrzd2fCfI6nc+hkO08sBkvMZQjyPl
yfE/zTTV6m2bRMXdBZjzZDOqkYW14t6CBg34kihYReJEL/3GHpxUvRbCFYNp
PozBJ+8c/pmw+pWFGyhHMrPrnHA9fjaTa70tNfP/37VEInzSpfbrO0TF8CVn
gb0eJwQ5uxCzcsK5c9nr5dIZhH1yCb+CLDuhuEtcAHVW9J7XOLWdLVHqNNzN
EQACyTEhjK4FmxyJy53G4EK2BuPiiMIx0f5ceaJzrS3sA8VjLr6PVOPMHMxE
aWcLanDjRbRGQqmdfUxIXB26S2rtjawTvcU4YwTLExVDOdAiUp6sO42Gtwiv
I0v9rRYldzMIVT5YXWI2493kmUE9WQvSfCzJTEUdFAMjzVhnPLbjLIv8fkKK
IFmT5bzLIulLca87E0DcbHIzpuONKt/FQNlKsIp9sMWnH2XfCviwiw/+Ds2r
1dnI8GQ2X6coi/sbFzwheTNXEBi6OJDEXAzPJOkc48vEjl2WI6kFgVu0dkAS
xKLy0QhlTib2kmHY7raj4YOtzuH0PnSj96VBqR/azqJhISlyoU8csoMU5ikr
yYPWasB+pmdtyFczjbDmUZ8X4XZKKKWcNWWSfNyDUAzN/Yj0xrugQSHfdthp
3Xnj7Z9RMRb2cT9/XbmLYdPPIQ6tp4JzO96KIgN5aQG6Q0XzspfAj1rqOZHS
JSHUTzQgUiG7CiQ1K02mshupuo2F8VoVDVdG+saKpuv5vNDxnCKW0n3REsYm
QlA0S+nDzt4IiQKIDlmy5obNTzOZalPVgJbgKXoGWw6jTEvOAN7GncTXYBBW
JZNrHD+1Gm/c0aqOHfiikNS3tDSKFoLS8iWd3Hy7rrDGsoF4HACfX5FUVTCH
eegqrRDxmWWP3nEo4eVaMTNZUYkjLvQIQwAcD2/PL4nK+R/w+Tt7lir7OrbT
q8MZFE6QPqn6TBdwB4/g0d+w6bxIh7jIiRLLq+vd+xmU1uQvHNpBU1lXvPHv
1oNTvXKUQtRTHf3jJhNxygcZIwU86l4/UN5EXNuPkyZrRoVeAFqpbnx4eECk
x4yLBMIX95+jJxrFzWgDyYn/MpDqDUOInyPhQtu6mK8ugIX65H9eIuxQCEsz
FtLrLjCzB6oVn1aJ9wUQbmZRT+q4kM69Fsrmsn5aF9J8DleDtqC7Uw4kJ0Bf
H1QV72jFLSiWp72spWGm6XJdQ5x6+oee5Y7wo+E/G4CDFGWVhOjgql5L4u5r
QasBntdm28+8PyogGNN7MdLdAKWBtt3ZtoqVEwyEzfZK/IMY7enEdd1oeN8V
8pZyfdIemNm6rq5X/ZLDuWLIxejz1pw1eF5HkYDqoWHEEHtasPqKQUvAT7aG
YQUYu+N3LqnqTi78BMpV9S5BrzoEI21UsGgixR86PRbQwOENbfvkI4GFvhEH
EsrH5+PXirFzf2zRQIWv55/09WT1lQUDTyxSeRTMNrvF+8UzRc1aQJqzBKRx
lsWesArTnJqNGuv6sOQXmGJx7+qO1LT0dUo/FdBKKDNDPrGzKCNnTN6+hbTf
FkqmbEXiwZV4wZ2aOJZWvNOP2Kjx2lHJ9yi72ifGZ5OdCZgHLo4/qxoGSopK
cwQEMH8iFaLFEbK2UO+6TUsOeoZUBmowe5+/l9vi9KQuT216zv1BA0Cq97p7
jJqDtmEcTFkSN1rBOPDPRxUltp2xouirmNpKRfN4Xywsc6tDu1A1KvgvXTxg
FxktbdAG4rnzpDrZh1vodFPQtdybZuhVrCJU/osKhSJx/vUkajyoGfGPZSGw
jl2nqdT6RA/KgnQvPNpmRRxv9wok28Bw1BshVa1dXmP7n1Wyff0UVYdcM06h
LoloDo+++9koWwwRkxvA6ps5/an/8Y5wYj974axek9ogXRbzz53WhW9woslm
JYlqLc7+7+GjJYekNGLXVDa+Nb39vVDcBzOgsGikW4pogIkDLEooZfIPSmAe
tGwfel+ZMAqj1K2MMMvmmjWqn1XHpHGBaNEpKx9Dit8FeIx+/gFf7rQRMpFd
GMsP7cEQ+W3U/xsvNf5K5YYohr0AFWtwWx9ymp3dK3+Dta9ttJmUsnepUI87
BiDNEdCso4uzwn63w5kGrc3BFNzgKgAd99rMUdL8tOMpgVVkQm5InGwYG7+p
xEycd6jCjUFsYAWB1bKOwW9obcHsTSIfibbLz8VcJsKQH3krFbanMWDxaOVN
kAFp4UHe6KjTF8csYSlKO7WfQkPc/2321tpoAEOMjG+tCnoVsk2+OPZOnjlh
NJucDaskXlyB1Qc+LxH7+OmEPzxXZVtiQV6Lz7hTgKHJPXfGwz/v5mM0FJrD
kiNwLkicilgepQLeWgTXlRuABIdt9F6txi4J1oPK/YB8p12L0zwhQWvXFVi4
+YeZjdHAvT2NNa23r4vbHEUDOxCt1Gyg+piuSN1oZagD7a0YB0CB34X0Jnah
5p4OuiYfixDGUqUfgBY6Xbaxd92JQzsQOJkT3u48H4Ij5GkgWOBFhajPZxxm
9GBjK7GcIZKz8kqHg0uff7R10ESWcMQoU9IQNpTk19iSjn6fK6QjGMHoEFTM
4OSqfmnZ13I7ErqEm9ZN2bZNeEbHnearxiT/qglnlALXPaf0DrwejVvQi/WV
UY+tV03G1h4iRQCTUHafd1hPF/AL8DRKCnE97Spv73Z5/gsl0kZ86ZK8Y0By
DvhgR9+grdF1xCIfNnz+JRn4YVZhDrdnZ1rxnVWsik6Uoamt0pX/EqbbeesS
uPv1C6fFN6YblPoyZlIsSOhUZfyb9oX3+6U27IWWyFJOpXF+qHFmK+fiSNA9
thSnM24UL7wD8i+o1GbTqO5ik3cNqlzqSBQAc90AAl/jW7sxZKqM72hQ1CJD
oOqcpX0CN3VjqIuXWBgqZiOXi1LG4+sAz3oSIeovqRaWzpHVFQ+/OxaO5OnQ
C4TX0p6Pdd7ZHOQSqERRYHhCEgKml7Mnf/IOfaN61OuPv33j59F5vjwo/FPf
SxVSYrDQUKJS+NjMZadJXum9FDa8/FJdnNAJPZAENRaYDfkgXPrKgYNdv0Dt
tk4ZIL6PsSozhK+kEx+S9rIJjBI4rPiQM6Hvfw9/lpUJWKqtmxDWndBxS1gf
X/TyhLpmb3RrlVjiW8wuBVqrp/gboZK0PdRhtMFq70UFfm7T0m1je2w2Koso
lwPGMWchX6lmFSzrkbgUmedr7LUNXMJGdeQfe2XvItpMulVYlQVfstzaZHJk
RTgpPWjEykx2LVBUwnYaLuZodhhrhpqGN6+1WwLk8V3z3n/OTT7ehwcdFFNx
duUjD1TzeGoWUG0rN3FIubn/Bh7YApAEanAPuPJvPVD29H1qVX0i2oTCdghe
crxOljrSYNgz+sl9szejbZGvyn/ww3yVgPvEW0Fw7wezT18Okyfg+vcXyP3x
8Mrxop5P+dbOgOxxv06rr9nM42GQkSaSUdl3OQiRH4TzJ0OgknZarvBzxc37
B44m9rB6gmTxk27OaAo0xf/Y/rio7im4L3BP4hb3epu68751j4IlFrcT5nbR
awyTffXPKfP2V5m5RAloAYtdKmlCcfbEsHuAGGRD5ULIj7VK05VDkaY152Qd
nnpFa5B2bgFaJmsepANu6NBfzcfoxY/pnllL73YZf24oh5by91BUdqNKLnEf
d8m17vRDLl6TXys8ODGIqB5B9Qj0DrIs0qJCZyHI+j61Z82I2trf4OGl2ZB/
ke5uXmYY1+eFVPzAWbibcvpHDdV+k7QmtgTw1g9CDuRQlktTRN2uMlmbuWMm
6ctZozIagRKVLazrv/5IAk362T5yXW2V1sPHpmI5EEnmQIQbEdbHwxfHT9mH
RDx6IroEZMvgEIN6nkQsaTk0FRZ5eq2wj+jpUcdSzKlSSci75Bco1aYl/RRw
1VmvrIJGQEOkRlh0QQRwQQtStDtHPljDt0CncKxQPXqlDXV+tak2BMiJDb6c
yum4VQ0tagHzG8JRNvLlJqKZJMq1jnuFctQp8aBlaY3SJtyxIXyc9Nu7wQU1
mMG+7V68FhoLPFkiwz5BxWUWJhiHsFoi6apPHXwX3cLjodTKY0csurcn96LS
O2N18A1rihJsH77MY7gIrpi57eTmWGlUhhlxYt/OvR/4abGUq6hhaSZ04qJI
GWcptXY31Q5t36MRaC2QmdTTAhjxfLxzbCU3enjW49k/R58ZJYRQP4BHcpp2
S03EySrczilOWidXTD9OjB64wW5DhNyKs9O1u5O1SC9M9Gh2RMrL7mI/1Vmp
FbdzkoukovfzTOQfy6ufRke/WnruR64mKkVcvOsl9rlno3c2vEebwziery34
ZnwvDVcUxlfzRZOt2lNUwgg/TmgCQOcjW/fKtdwfPoyflw9ejdgJ+ntz2lT2
hRnlrzV3mH2XAKhm5zOq9vw4uftVdUD89YH61+uhUwCitVMT0WsHJH5lnux6
zqPB+u9doqXzWsyjdrkReFAXVf+weLvlsN7kGzxm7TliCWena7CMo9btCH7q
IAo45RRnP2coycBC6Ltq2rx+mzS1zAecaYYM1gZVbA4lBZy+ZXVp6eqgZ7d8
A2/3cZd7I5jh683PvGGvUaVHNDT79AI2qQlglXYYjFeXhRwmkWjFHCLJlfMx
by+r45gqGvWTSf8QNcDs63EQBuDH7ZMa5YdPG6fTv9hGlOmGPQ4iwovXKItv
QsUGpPXhIch517Qj+3V61XUiaEDHbDxBcCw2LsWDFRXhWGtKId+prO1yfxxe
uAe4miZ7VBatDJbGLTazpdbDAfogLynmqqv9XU3AvdNQ5DHMZN6abkKfgJX2
3K0G7c7f+/CqDcMtp8lPwQDXojKQi7w7KflSlgEVVjk9ppx86fHbVUWnkBL3
sGJ1YYjd07VQNGuw1pobAj34efWJ6qjhS9hVXhvyOhBgqiSc+4KhfVKcXv8M
uHd41iyEDe5pvxt5FAOQcgZ71dJIkfAVRMO4snV1Vquh1zDHChN44admqQW+
PjcSsFzdG4EV+dzCwCrUVG+kDsCiFjPNdgjMKjRv37GPg81Lpi6FeRIBOQKF
LasWIiChncOtXJyhk9uhuecxI/1w/PweJc1Cyo8kcIWy77Zk+Nvu61J5+mkY
fTclt9hLlgThIzxBJDbCW8giJUHUMSPz1NwsVBGnSvJUm+lokDVPfCWmmMq1
U3+3tCME/wY+ToymT4Ak1emQwW2K0Uejgwy5NCjdwjLDoLWwiWWF4cva6MJw
/TgXBlBBEiky4giBtDIuFEUF+e65PLZaYszQHXuMqluf1U3cgs5y2aU8iCwS
HLGngnykJueSsur0Pu8Lcr6vSIHyC7XN0ZPX99rf2yDzQQw8QJeNOcDG24x8
mK7/XKA7zWraPZcBCjJhgtbWBvpy44b/dMrBAtpxlz6adFCtDMZuHcdGGOmE
iZYPPvRADAaR6BvNRKCeA5VrUpSsdsZlUdcPsuipyUTj5Axq3Zl/W7ZKTCEt
yCSMKc9ATjs7U1mCvFY47Fwcu14p1YHNJVnCNo/qfpgWFhgGceBdBvniIelU
cN1nE/uLwgAopUO6wpimtvFHm1n2Hp6mitael/V5Y10O8RRwHo/vd1cquRXv
LMoBsU63zf/k8X2+2/LNqPHAKRk6/5vPqbNUHaM3xP2KQ0XJWvbaq8gr/2H+
XcyT1Ve+hbwbypU17ezI4c1tAbQpKXLYeN6fu24X9e7LO+BTRMQcg1Wgdqdk
/zuidFO4pMxb09a8WE1nksIJ57G2E+KY4ZYkscAhJMLKb+4V+SxYTG44gLOo
6ThI/oKeGgI6uRc0lbY/MTTg/BWWDAX7wRrKICf4H1kycP4FKPi8FSAOY22C
4I4bkArJxWnZV+YyhltC0SIvmVZk1bSIrwdfdg15hw9GpfWR0OnBVcWse2Ig
dpDe7VwAySILGhL+Za4Q8u4DkrwKN0SQRKNgg6IW9uHahv6ODbeeWet6+eHG
yL8bkDMvIcvMN1ZzIzCGpwrTXnvK6uuXe2kEIe9Woorezbpr02aPFYy+0rvb
guIpkdjj/pBdMBmfurd6bmXndk1bYXITqW4luThWPvlbBAf37wCPMyIdFuBW
TdPNzDDdcJw555pAcurE3sPA2p+B8nXyfIaXamvnQrKsKzR+bXkxMn0C+c8I
tw3gG3faxsrlBmQQ9Z3jqObBYY2gZZVrBknVtNR8dt1M5wK6F8ANltLBiN+Q
3ffg5MJxR8AC+ws0sCKJo/Cfjz0vhnsSV4zg9vE0cjtvwE7+tZbavut9JN9H
Zor0oZe8aFskfmsk+UInHUfWk5zs6TnxhqkeeQgnoQ2jTrgbXmc8bavYDukK
3IQAHhABFNf4HDmxEoLp70rY6owxn5Z1qQATSqL1mGn4RZpSRJp074sla8At
qSa73zdx2NNGiMc5r9O9KeehG3jpg18Iew+5n8TihVhX92DqNZxRFpBtZY25
K0iqt17lfSHDAocRLcrZNzgCejqm4lo2f5kuNJrodHjlI4d+tW7C+KIK9Nqr
N308fZbBFz5WrtA6DvGfI2xRViS96L/s4q2IrFfh7Qe4x9edL+/EYkAjiC7n
PB3Zzukp6GtMpZmjtA4Gimd5zZSNMz5pWNHVHA1PsCG5MACMXyMsgoxNH72M
s3O3fmjvBr7neacIqBiC2Lh3OweqRtjUejHcLDFHVvMrGTCzdCBbhoOdTzch
E9YOFnQJwUKZHtsG9kuD1j1A2HWQzEoBwiaRptQLP4TMC/EemDNDwEYJKVb8
pCKyqq/BEEMMkVhkx95R1R6kRtk+I9HIisi6V7FVd93Z/2apcGFwmSmyKcPk
G+tpDrcsWdYOfx7CyWoL5m6RR7ZduLMbrQS5+fBp33sNhXTtgDjbMxdfbNNl
sJniPmth+qRkrqwfSiXugZGOnRaxJkz/LKy8MtK+RCT7U0P5IqbwXS/rAtgu
kNEv624uLnEFyGpXyi9a1jKl3Xn1UTYMsMgse4c4HalBxANcKWSxUUz1WD5B
8AjHwM5t0E3gf0Ot3eMglRe/oV51WW7bqZ8nKY9sUMki3wJqL65GOjzaHlcq
V4KSNZk8XYTQbXpeNHFuhjAMlxRW01gdRBeUsAi/aGijRokISZY55rozD/tD
AK80NtjUExJXSY17t3PNb6MxBx+FjrXD6hUB31GwGfrtVIMks63Lrn7RQfYv
knen66enfmiZk4ARZj7XI4ZXDxMXUgM0PaqbXpRejAuWqgwHb+LahLE5DjPW
Hl4tQKICI00hXgELDTC0N7I1+jilJq7dHsVcty0QHzoiQL6Szoejf3I6jlrp
2emiqpb08GT2Y09ddOo9TmybzdL2oNacVrthqDDnYSgfQnvZ04nbY9gi7Lwb
zIQuWUNdedXuFyyBzJNc22ne3Ua/De5YGajkyImRorsVK/o6cE5bn5ssa9JC
BkHPup+4w00p768Oh2z38p0QSaFxnpcBN/bRc9C8NEFwFdMJLZUNOMYcS1of
paXAtKcmDu6spq3CZnWjv6gbvikSaefrog5jj6o2honSwgbjJk5xY4Ngka+Q
fjuUKWb3/MoEr0sd8Z3Qj6+3h2Yq/vbYLkCcyGepLPc+iayT6dOCdq1Mg8Gb
CsqXFbZ0Uwxgld05qCG9f5MK+3zIDgrQMyvHkAoqYRSdHX9gVZiIxd/qvLqr
WnVaBwdM3Pi9UrNiG16ZroGFVQ68rY+2bFQG91BczfGXaBuakqMgmWSL+CvI
F0w72dsaNJUPhRi4i7RBIFV1NSeazkArdk6jRGweG3+BLyZ2U/eMbqE0P/kQ
eEN0DNi79DNHDAkHb9sb+VT82+z9PQdm+XCCqtWC0PDvpNjkSqqErS6OfIjs
5o180adCkTi86fdvi5OzQ8+MjXKxvn0tWKM+C3teZxe853O2GP9tB+2FGG6K
qT1/ckHRAXm1DB9yMt6Vwmn52nrguIL1155iMlSXWtN7CVxP1iNvBNY+4iY3
10R1+Yz4HN/zXnc3f2aOqgj5tP05/Lg8KPCyQmYPeb6TWMKi5Lmx+9XhWNvY
W/w5OmxXDDrnlHiwXmgEFsnq4aKwbRcmefg2oCMfW0XEZaMwcQC4rDWQ5Fb+
SDc/Svt9j/Wc2s+TEnqYnGqVbwwGAQo2a/I/kvULBgcpIDfEl4z08enWF/Rl
jyZq3sHXjqcFBn3YMjD5JujLxT6+gll3Q5Jbs4jtpwxBpO3HnboyvtZlZghO
GrvSC5O0xDUYqat9hw/X07/LHQjpPmgkzYs6RbCYxUKq16P37DqWxtWvuYg4
YSE2o+9Q1+Rvcf5p3gN/rMLs7sxD+IGDStKCHjeJ5uUeVUCZb6wdT/8cDukP
iUoxQC6TaDbd8SsL4br8kYSdolqrHsn11IFn4092ZNb1uvVdwIczUi3V6/5o
pjBnU4Zj1FgV5N0XZxZp7H1ilDY0lcTyVNeCZ+0pC/E3RMpRwI8mJL9MrK3u
kx5/4NEVHMqE2jLxX5vDFT8HYIGwgMAMphWZqt0L+zBHoEpbrgIOYSYtQxHO
NL2fS+Q9oI7I11HaQf/grkCdgic/cp3FwljS/W2j78CTYKZCotGALgqqZzmj
vKzD7maAZqeC0IIKoUJrz0YxI0stngnzEXBemisBv5HChIyYFlFr8SRLRU0N
IwAp22RwYtBIkqpwhEZ7BYRYJdjcA23/QLrewwaNX3Jtt+0DbpoFmsFDkV23
Sos9vb+sKBoG7KPbQOe03Pp+ONi3hWdHELNuzro+KDPdfX9QAjGK/dM4T0Ii
4DPHqR2iENMAJ08XperXYQs1goJLq+/ALefO6yNrWJkIZ4t8tsg21FnOaXql
SIVjLvJybFY4a7Wb0CKF+mZGk5EthScfW9MVwhIMp+lHVOeWygWbkrC7KsrF
PYVF/yBg8H9xgoy+OWtPDQTNnRPGxj3VdCtuQYHVfs+4WcECCmEOFhWVM2Jq
aYrVphTow/oRG0gqpteN9B33WJetYN/+CgYHNcrylkQQufma1bu46TKDhEN3
kNnlxhluT+OBruygZ5yeAGHrB8oPiR3d5IRL8mB13fDMrx3rfiKeX/1pT7u/
5B49otNHvNHQtEabsh5z9MYaSaAzuf8FekYzc7vcOtTokXfi4L10i0xmq8BY
Xg7W2MfbRgHbH4iGEpMHcYrGTgekUwt8TL/WCPD7jp+oEsooVWUN261uOerB
z3V8wABnYvy+tLvwnVK02/dhT7acnG1yqHFNZJFpvdkmb8EUblQgGaEpD7cW
pOK/NX2Ah8GtADt/3k316pTaxU+3ZSSAq9Kh81ZKHDs9AlK4mF89q8irkg6H
UhZWmiEpWcF71Kl+rKuBCXdkMAkZBGH2MQXtm4tjkTG6X4pje1lmVhOAOKpB
2GWAh4COspd5a3M8MpH6AreZOiETZcBWvNFNynryjGcJe3dpVyRDY4OvVyYv
IftyNoLzSJFijpn5hr9xJiYudvx/jpz63aoSRNBoxg/YGlATooTACovZDeQW
CJ8clyMjIWg1dUseRBj/4eAFDY565Xpjcj+OIS6fDUkO+YvdlJHOTyRu79nl
/4ZAHQc94Mr/LQbS50Lf6lyha6DlgvTpc1Nxl74dBhdcTSPGrkUbocz4Ejz6
H8eZd8wJnmSo77P2C7mprML0G4uuk3Z4TJnPa+zyGcaBu7jo1qVnstVoY10T
9Euk9n2G4Og6Lsr9Dj9vi/yn6hbWrLfoOTvg00aR7En4/0c10xiHGeoT2tpV
U6WYnHv6ZHaUmdautFIiq3mXdfpdTDGvD0ZvS9jCNF41mjdag+AKjt48LeL9
ZNfRX7TTRQ/ZgWVv2VQTOby65+mNlCT9ICwsULifqcFpbpywCm8g7vFhfd6T
wFX4yH3Bb07HxkkNvcc063SVvTuWpIkcs8ptW6kQfwDRwaOenBixNoSU/9Cr
PJ3oqNcw4aalQdfOeFJtRwnz+8WEAqqnwB2Sv3pcgLSO2B4Y1gYTpNLYcort
J8sAvEWViub7zWHIqHkny3Hq3/np0nmhuC9kzAWoiQ/0c8f6e50MlWZkP87q
ctbZFSRf0KieLO0nsCTmU0o0aaAVTbaEO0O4KHF9sHKkCvdJxh1u+fbGBo51
ONmfHOqnc5qqU9+rkfDtH7Ov3rghtorNJ00i9wPc7/u+HYWZUSbhTdC/A21w
2FerDFQpjnMVYgoD7poUaEWMtcNnptLhGrqAvpfEyyMZ2U55QVkUizCbVH/f
hr8ZKeIREsGHRpSUcF7jdX9A0xzMC+e402nGa025UYu13ZngNzQBYiDgO6kC
4/6yGD6pJeKyfRd8MZeeeJBrjlNrAsmmnq4Rv+Y8Ex3AgHYosxr/ChcLpQWh
+hsHDuxNaM0qErBOag2FFiMn/BDJU8Gyh6trqQtJ/nJXZSW605VdIV+J3Rn0
tn3aUFi0b/n4klbWlNm2F2Z9zbGuDlVOUIkuNc8ZKlVB7IoJSQOFtFCKDZca
5Vg3IjJnS7fNVikFwV55YxP0tA4HLM5D/6lMYlW/TDreVyR9i1c0Cd9KFjU3
v1AoV32sLFeZmZx/zaRoBJiTr+gJ9O5WR4j5435sqGNezrbuLmFySDEPZXGs
E0xbITrUXH7rpKMeZ5Zg9nmqpWkKgQO5uAkNJS6cwErbVQopugxSX78zxlc7
fOAascP2aTGinC/2wIF8SkqNlJzLGKr9l1FARo4zbhC3i64MfoGCKu6vtnEj
YveCWmM35tr8+fOxrXrodXj+FrXeSHmMMCBTLYWjT7T/eQbGmuZwYeo+dK8c
xAByNm4oZ8eYlejdgsbcWBNIfw6yuocU5LeTiNfgNPhHZprwAppXM2MlodVr
XP+czJJI5qHr6MTT2zbiq9YVznFDj9YBp1SVPys+jVQ21kVTuDTCIYQHb1GS
5QtmC4EtPWoP0STPNVANg6cUNQyZDaHIzwM+8RfEnjwKjSv4eCxEvL40dPGk
EBklKVKzl+saP/T8/noWKPMXQxG4mFmfBVmQw2ApgPJPa/U+91zKTANqflHN
8i5LzJEnvcyFXTRZpJaMe8TX+J9LORLYDFYWspD/8y6XyjlSUIlkqwufH+D5
NIK9tqf0le9H+kldv+wBdfFCo0R36/rSVG+zB5NUH1bYurcQ6vmeGBl7HONt
2wiL78cjQDLSo60kWftfw+4iphyZKEcq7ZR3LV5wTr3kzVwwardNHemIMAed
bfWSEpnwsicoSKpaaeu5EQ3TfzAuMG2bygZlyyqtkHMLt97I4UGjkTfdSb3I
/FKrgt/MdB48dx7gc8b2TDIv9LrS84cK4Z+YCg6WNTGhC0QUf1TW3RIzTgVH
6XbY/ty/5Bs9OAEQ03gax2f2WPKVKkrTPETPOCf6tvq2zCQXRITUDQqfi/dC
gFz+MWq1EsKtPNBeQ0cwcgdMyXnDpmMsNnBL/Nn5rgJ0k3S6Mgsqf0ZX+xnZ
Ypm/4P29Zd0uMtvrWz3N6C9RhB5ZkkHHJZ6zEfBtAPW0SoKQ5gDptB7u3Jst
jy1HKwH/z3VCpmFNCMTE1ywTonL8FYn3UlMEV8FC3UprqYVK8c88F4G487PX
1Vl8Pr+e7yDg0X3JOfKqd2ebyjNLtwFANsCq8+ldRpjLnsIZu0MnKL9yMRq2
EJM1XggAroyoWQOtsa2+lfoF7mX2opbfr32aicZKKWEgbznVO/AswdHYgQT5
TH3sh91jIXOPIp0ExkUlmj4JSCLQlf2AymRwjiZuID/ngKeEaVBGJTeYTlLQ
pIF9uPzSi4nyb7waGhwYuB0tm6FMJBnwKxKXqOw1PCyq4JWtz/C6Zc/vekax
kSQdtTDVnqP3rULpTactytxwI+xWtab22blZFvQNQROwTLj05KcADngJdY5d
jPqcxlDspxYBasz1LoIOYrC7eaLq73yDIv2T02DgyIw8qD4CVPr0EssiZEOU
b1txi/5z45EPShRkuNWZcTBrRD8CgP3e7mCPXf4j+JxgjNCxdtjEllPzeQ/G
Ca9sg3dPDILbbmyD1m58onTsL07g8Ch7NKgPfhQOj/8Dr3Ma4s8aoulVPZuP
nxdlyUlGeddmHGQIlBc9Dj56ZoCi6J4p1G6PfGxkT7jYrcoSXuJPfg7bvaFF
jeyba4EEzTRL6BTCJCdZGW8GKh1cKlU1NpCEbYHSGtg+sJkVghJOphLtxghT
7Pko9p80vzCYpkHBKwSw5SxYyE0NsmB2X5fhaXyw8xofOo6+/w2dOVd2PRbg
YcIKfkcEe+89jKJ4Gpm3xloR4qgRsYRgHHQ6q0MxR2FAmjLoK/f381ln1uaq
cFs1T3jM4mLLqAD0gzg/odRRUzd8o9UWs5v70VI04sx8qZn+I8+MvtSfGM8C
v5H3VwWW+kR3Cf2BzMWCcSkJsc8H+TvoMubH+ApubALz7y6UtOyY3JCC5yyT
TLgnVIXM4+IlGGObtUdKrQ9fhbSRcnoQSHSHbSFYynYK/l1vmm6qsEhVWrMu
V6yyng8wOQb5FVqfcyPKbzJ2t/askdpQUw4cUYjRwioggh8GBxihjWVEPZ2m
aPoHpaJ9xNpEczx5DJNIXEB3J36/1PpNsmZhQhaUFQYYx1+PsvBnAsTDHhPs
57T3a95QaoDfkRUXSmQT/NrIGtcMv+eWkkKDEYES6OBlf9reKRQ3/5x9ivj1
349DLEpygBCctp3Kh1dzE4AUGECTLH7psXiUGWtPkF+6YfLZmHZODPbGsPD8
2mMfrhEAq/axXZ9OKx2d1CzFHDOTTgYzFzJllKZrXuzQqKJFJkrfmE80gKUK
o15cDAGeyq4bq7N04psrXN0zv63AxhPD2NuSlB6V/AjYOFsHfcS6MFCKVi2+
iGeO1ukLzcJIUYBQoU5NrTzak3lpxY6uruPbZX+c+rXmbR2YXEnbWBAcqj0+
jZtoSKPjW5wGMYp5Y21NC90bq37OwzP0Q7YqKZvH5OJapnEfgy2Rd0sGPeRx
34f2cJC7IMeeAEuWehB3Uw2mhCtD+C4PcKtcJ69kqei+Yl8+R6mH8Xnkizn/
Vy3fe1kCL7NRaobq96c3v8j9oaS2zPa3rh8IAt0RDUMqoldg3Cl4J63dgZWi
DW8qV1uOI6gRZfIJQNLuhihtfX1GB3lZpZe4PtJZozruynJ1Mh4hYeWuNWLy
mVD5tuHVMKlIgISBVKKymMGG+o4eicDWVtAJnkcRIFlNV7UwXmRWt22chiHU
KcqKMfXRKsr4TqQDT2XvuID26CiPx5pvYad9VuxVfiMPKin86JAoNdc3PaSB
/3GBLS1/yW0tGlNuugJyTT2FXGDdxQSafhYGOWlk9YaA8HG7uDFIAvb+lqch
D8SFmwVKLY49Uv+XMQtnfCFg9L5ojzh3BB8JGqfWGJiV9+CrKkh+oLzTCkE/
NGgP5FqFvJp5OpJCRecQeE95K7lJXmN61wamleMbnURw5vYzf3Axghrm04eF
6XIilwPG6g8Vmu9njKx1gOEIWmE8vFmkL+4zeFLMvQrxEn6DEFCJOE1A+4XS
xRFOpKSSbz0N8DpqxOcXo20oZ1LrMJ/stxCs+UtUjRlrRpWM/ltgAiCmFKzY
Y1pastpjRlSp/0lJJ2IDQs94Umk1tU+q6kJFHtkB5jRCT6yD+qgE4v8dt8fn
Ex1h7r2Ig8XBXl+bjJ5JAXNMqq+kkazvqLuwhMEWeqnDBLNgsaTk/zYITG/s
LpY4QldSXkJ1uckZsIUAr8Z8XDOXcFonRlrwY32NZUcqki288q97nghEjcPK
qbiDgNDvdqU0qxPJsKBgmiv3glJLpWEFGalavCKeNoFEOaAaLHlXU75HFrV7
qgQCbwW9W1RZwJ7QCCBOeB3pe47Nc5lmtnM1oRgp2PchcadEWd4TmSHeYLRI
DGQwOjVMYVK2z6ecgZMCQFlNzThTw2X9i/DU6Usji6jbiiojJ1QCMd+PcC7F
pupebRNgbWZfdcuX7/7uEvs2fh1LesVo0LfecNsMBIhj4BkfEZ6P8+qlcs6V
/7ZLJpBrevmZ/RgdopKL38f2rvtqS426MN9aJMIARRub1Qf18ZP6/bo+e0iF
UZHl+IqpsRAPZtGG8ohamo8s45RmBtDyRD2BeQgbpnkmxz1tua23UIsTVSjI
8iuqw+0y/bad09AOLKX+MFlBCzz/78QD1KXvcxPTIwXDxaq4J0OsMz+kcTUS
VEu8iu/xXAk+daHMIzZzTGZusGS8cOlqWA2WJumtZPBhYAbUw0Qpfp3v6i9F
k9QDPu3gU8bb1HGhVxJfBdKF0XyuwmUm/vkqk4Se/msY6l9SkRJNhTAfSf2N
QZEqZhlyWyWs9E46R/kW4df+gDhvs0Snp1OUsiz6Y6/dPOmqcO7sId7AJ+xn
gggwEq5fli/dyUIUN1oA0doifCtA0j5hkkoI9MoijL7QsEDJenSScTAVI5AH
Jdri+V2TGsPcUMKu7aQWr8jAraH0ydX5123bO9Jn80uH15sfdiBo0+b+prNi
KATqk3tT3Azvz251IKYLoT8G9QLbkema2c5p2trTOFqCHyMlgJ3WUBICuKZs
uhqRk/7QWTe8NX/1uBiKceB2F+4nwUp51c2q612yP1bUVJ6CGMY+0BRopp81
3z5cxOpSFJrK6ST5FgeH01HUkT568UnvlDYpbYcqZXgo6TvUgwwXuvbHplhv
loOXEGQLfnGM00ORjJa4NpjBJMpZoTxvwXY2oCuZUaClTHYUImnMc04R1I9+
v+eP4uRf/MXn3ayMyUZNwfXCsL/d/pOdZ9uwNJHNU4kWxPgrnDep3vVAxSHp
Bm7jCFIHDupl8XMB+STdtnnNgwD+Z6fbVSrwsgF6t31nbmMZF99/0lxbWE9n
fek7BLLKsbtjNNx3Zk6L5aZANhQFSl61WHRCyQCx/RWDFv/KCpTJQp0K//HP
L/hlYu/NMT98QZeMu5GG4cHtU32yY+94EjNy6SoWj4T+YaXyuYcoF4VxwEDI
6V+HGiVye0xLgBEo7/siYdGrKVMqzfhd13Sf0oSyh0yIQZhv+KirpNUhV0po
ggSUFePbt5VyawP59AVC1YiyVqBq07O/DDat5XeoWXEye5dnFa+AjBW0Um97
AkgoEGr5+5Yr5cGN6/5INzPMU88v4dRJkpLfNi9HjJnJ+8l2YkU8PBEdm+gh
Koc+CYUIN3TrmsS7DzlQ164oIIC6VtNgT8dbBMLex8dHsw9V0ufZXfhQQmaa
uqbg98IHieqAtliCNeIZ2UTVqe2xl2ICWs0D/PQc1xF+LsI6RSP8R/yOaeUH
eCeJtuSOHMq3zSbUW2x4DALs4WRlrElT1mjQAqxr0Ub3PeOOmlaRvB6+bXRH
5/SB6QWdXILgaj+AD8CKL3iEpUuWhyX6+yemCOA0DQghSIEz8V1UczIGPb2n
tccOPYBCTJfZk+84IU/UNWAxeST5J+1ijIHYANzkumoctzRLPtV+xjGeCFQ9
rRvaPZ9DgTlf1jq44Ge5s6e2Z/UVwWZxdOe267vIzZWaB7HYLxtOT0U4GTMk
9KKHJLQKqQneH8Kxq0nesh1VFaN73jU57O2vXmiymiVx/DHc4M0ZQoF6y7mm
a8HHv4B558Hhaty0InD+WU9PkUa5cIygYWID5GssZjhyyqisehYYMYtiopIQ
7LidSGGoBafU2DffDp8gFF0UP98ASLH/ob6INBQbaZvsLH4lHnrllQQb19OI
M5k+a1HV5Aaur8iEWjECvPS6RfpMXEp7dio2VeKT34eHOVneqk/7lMi9JVH1
pe2xXMJH1v1CB2ITqUmqzfVOa6HJAAe3Q+n+2xqtTXEWkKi+dszwUlx2BP4q
P3G/sfOE7SfkC7FvH9Ss3AtvdE9GSwh7EwsuEq7Ua/OEa3xznNq8CHcFCpNB
MarbsYF8gkLKMr16R70pAW0MVqX7tcycvnDoO23W9IWiFSSmU2uf6VlndTH6
Du35t3gXfX5HwtjzGskLrHQvSzPoBufzoh6CxjDFNLosPVhEoGymjYFNByUk
RzKNvDhvC9GJTVhi7PKdeaB4R5xAfonbX4JkFRCrS5/xfTtDjk+qvqz4OLpF
ujy/439YW3OjDXBTGBuGpSK/O6rNI8H9SVxF+QIrwSzXSZeh8EiGEJrePlNU
A5ND8CiIf2JZwmrP55ORpVgp2LwsXv9Begvcb08hDQayc0NEvQ3XoKiG8VGU
RpzHbQHOXKvQkLoBtmmAiLTiZTd6C0gOvK+hauRZzHlyhcDsSAPQJOUASSLM
nxRpfYVhGmRV/5iIfrB8xny5OUFm7vuMiz+sqBR/udzhE+JUDNFbRreNtOuf
9S/PDAicYfi45+iNn7F24vFt4Fmo+87q0DP+1shEKOujOJc4YmD0kOCbGBgV
+lP2nrYbvC+SLrvwj4MkZGsuZkZvXQMzvLFnr/3+vgqVQis/vBsI9u8Qvotb
pgu2bJRYlabFXpjUWFPAkMbAKLvtsRbSRtqur3SCx+8aa1kij7GExhKbZVKZ
y/iiYoykqnxwjN6QhLlPHcnHAmgcK/2MbtyQnd3Ss5hm86Q03GssfwbAGsXR
v2POAcP11kbFswuFhcOx0mfBcg086ZipR5e8PeRc9HbN86b6s4d6/3TWuSuh
L4YP/QitaXtnHLIXGn6eNDzDnGBH79WZngJTPnwwb/OYdo5vMT7scD31nwma
zSCevgt9YJoYzzoUuO7VyEWkjhTz/QQRvpKt6tLIz0uglB4SY+Gx5lT04AJm
FQdIxbxUJDLZ2xuH2HLNfcPijuLKd2zI1Dpd9ankaxWiOnMcnY+4hz6FIbo1
5Mh4CR3+XAY7N3RG3nlamxNWRIjKr4/F6eJQ5MokQmhIteidlc9eeeukKpYr
GzsWXl4fr21+2prIElUHc6Vd1ifiQ/XUACa9UpzfWf6Rte+wIkFrcfWm5AKT
34hEpnTYIQm0iY+Mf4Imx8Jlh8IhQfE79Ki0yMT/r42mmOg7yyB3+Y5nM5zq
l02AU9xrmqOevG8ITPKIz11bcP2S1QPseZDAv/e1CU1gZ7E/ZQf3XZd2YdGF
2ZNbfjox6st+7MKH5WDgZ71P7aEPcni83xOxMycfwWelGi5c8Ii+j8o4juZN
mirDYu1jNWCTp53wjF5eZ7XQC5dAGZ29A3aGra40wZnCC4hn/CRZYa0gzV8L
Qm6CgZp4+olPZ7o8pRz/Sq+OB4S4WQDHQ0C54MTIzfvllMrEY3QzglG5aZVk
CfKq7eD9VWrzQ5AqWXOrcjbvwS4Mfkl6P1Ot4IWfg3usoelSwLAHIGXj5msT
qrK2x+fEKphrCbP+YhKMzWPNN1Njy7ryedyZsgh9idfnl2iNOWJeVMiya79q
CE7SwWVuRIdVTg723dO8vmM7T9vGrYbLG5EZtYKvpyR3KmYpSU7wNNHwEIQJ
oNBr2qLRb79k6ixLiikvTLLBSXiqiew1kTlxITunP97PZWhopmnCrmvI8r9O
aUsx6Qz3Gwo9GmGxQpwCt14pfe7l4de+Ir3lOX5WzfCvAF1UH7QyG/joa8RC
KBmkCnGrtD7dx0VBAtQzo4p5TTuwiwXOfT5uoXZtjdEDaYKQpj9QdJTY4Se+
zxtCmbcu5RqyGgAuueu4hcMy5YQn9AlyhBaN05zZq/MMsCdKBv37QkLee/FZ
+mZUSXc2CrbDwE4Xlsvd8jh8yupaArmPU+4Wm79Ehl1CuY61EDxaOs8jYke+
tD+0pGUck0TUyjAOCKZE8noga/nxxqd8g0mC6QtNCUO7RA3UMlupjhCPOHeB
QEU/jwXD0zoFiEI9fQFsi8VLX7DLKp1aXW0w/MAgd4qhA/OhC0Heo0O/5WSS
ShVvbmUjxSb7/xh51M37TBIpPZyvlDTX8olwdgGJFUQBh4Z+riodWlDUnj04
AgED0JehQLcMSmTCfHIy6zv6WHNAym6tJhUEt/+31YHAOI/PUmueWvF4qh+c
PEFNuXV0jH4kVIduq7jNMbyUnvDdxkPI4UE8QDRacvNGi+TrzPcLW2Mdl48W
hFj59SoRMAR0XyhSkL1n6ru6RzOczj54JmVXO5nt9rHm+K5OzomlRKZh7Q2x
xho7wmvs1Y2fsjXuXk32BOvrsVuJlb5bSTkfCiy2ArvBVnqeFoxAvQ0lK8jU
af76wKnUgprd5NT1HM5uBa7q/Hds+xcYAhcnD2ZqhMVAApOai2lIYQFwvhR4
OcWeyfAE2dNkmXyxpREnhWSprQQJk0kx6/SRkhNYcBg+OEE9tOJfP31FMd2I
gQ/W6VH75iyh7HyJotLwzypOhhRpQ3jwbC9faGAFDx+sq5OpxGRg+gtMaRjg
s4jZxS8IY926vF1Qritg4eBfQXafwPws0xnsotjIv+eZ5tQQObx5EWEBMP55
v2tuXpAIqUiIR0kpw5fBGID97ckt0lCUo2KL1hINvcnvjcC1ikvXxtUS98ym
IhA4ISldbD+HEr8rx3z7L3Ki8cnB4T2M4EyXXkw0T1y3g5RxKSMrFQce16Ju
nV4zen0WcCU/75tuOdm+/WVqS+ZQHIm8FW3LS6iPM4WWqFpNEA8t+qlEZYI7
ZW88Szxc+leQODnYG152gqyJwWn96PR4pSOj2YpQtrRi3ZvdkMER/G8Wl9xa
JXaiVoilEPQr/AKig8+b3Ac8WZGYkkqYQO6htiKDIrb/oL99f4wOOhIJWKf7
jsHHw53tUYxbN3qMd9rG3LOBmTAMCnU+ABd3ycg0DVdzlGIzb4t+44KFFZrk
reeOtP3gOmeuMYFuLgs0ZDPdwFqX0EnvMjz9bf8lkDRP/r6ptfhhhmi1Z63G
QZvPIoVTd/Vid80L/GeT+ChxGQseBuU86ifpHkaZ2X7hehzSNeZOwiWDPGoR
Gh4h1MTmdpCqHSNyJNnGW5fhxjiImC5n63lZVUUDsmUGd/p+atmmJ8wPgXhm
NNwch+vIdXBiJM4hF/WHF/joY1HGdmHw+jDtKiF6urLfH6Z9wz302eBL+mBF
F6grCIduC6qRnvL6DDmHIEvIuwS1ffX5MmTzLlMKOXIMHN7pAvtAq2/G8iK/
RSkzf3HgiG7EWrcqB3szKgAgVGdpxi+Xa645WibSQhP6YKHlgVs0ZksFaEsL
G211cGdyX6Wtjyr/dMm4X4G5doHgtE4RnrLEO0ESvLb6FXgGHYKXO1dUy5YZ
xrOy8YxEzMGu37clbM8pvgCV0+7zpGzBkgl5XmuudEuyLjkXTjj0TUxY+R3e
X0/waT/CH5pzy13CD6uPF6TioSsnmFO3gmdlbvQU0QNgW4MGDNqjqbeb7HGR
1XnNmvubJ8IgjfQq2Ff9NbeMnHOaq5pFsLAqJYAeteTvRW+05R0hONPaDDr1
5lv+4607+Z/gZAv62tor0VB6XRAmDbTF3gZQKSceetWniMcW9rYh5dIFZZPH
u7AiRAe//FGU5fa98bGeXqwxwnvKOL3hUMT6ku1k/T2Lx3VYIg/u1AAW/Zhm
owzPri2pt+vqUbqZhJv7YzKETNC0Ov04j8PTFN1RKqwLNl+Sp2jaS3WbBxHh
aMurOxIUvEpdyAbUP9RKENdkoAf8Xoo88/TaVRtUKyTS1p5VFHrRr0No9ciw
3IW21xPLeiTq7nmJMZ9HnWQOMXxIkI//PpmK++jy9Fdhsf9uw1jPrW67OKDL
JZ2J39HFOcU99eHKK2t1gadTxwbJ7+p7dViO3KzDt4Qsj8NhprFgVKo40jdZ
xU0IUvndvPL8xS83gSdRnpinD6Rf/nC3guUovow8tGnmQ8BIe2S9GkAZw0gQ
iV3GmIJx/GvS3UmZ8pINEnseY7xqm6A4JJqEyifgZz8qE+8OBcnFcebmbxwN
DE11nrMFnHlX/mQD3za2IuJ40vUbB8Xnt/z6Rda9FuYN128O27ZbqARyGEC1
msGw1ponhLGFU+iyA4fWe89oWAKSEzyrV1SmR3SiMtCy1IDb7rnh3zT80frC
M+b3ObvfwOsfpfcJpY4ktpXu6f0z9nlUQQ6kgG4eiWOrzDnOToJwp6Ouhb7a
5NODGxgQjt1M86vJj8d1FOSASOHMHcK9ovX0q0YqeeGd7vNJUoTaQz9ZMozV
BufmixJ5IdWO7KjGyV3Ne97pWHAGd7zPslt0PmL3W1NRtWwIfznVSSJFE3Tk
QgHWypuBfwAdyjiNit2PitEepZNxqvfnqtA75VFpkajNNMrCx1TiVPcRNb8c
v7KIbgnRUOEAc0Zizyz23DeLqy6qC9eV5/ku99tgr1AsmNjdFCWKDEL1gStN
UKKWYkrZWPJNN77PQNVoD8yY18ARt8jfq0mJdKaS/lURyaWvce0t1m7f6SrX
JAl2Oe2KtEvuTJfvlh4OWqLZ098KZPxmON6NNZ+k+bb8bhdQvJ5Zz56p5S1K
L1C6mJo0YrdAjqhXJOqLCYBTETJu86xOq5tMo4PGLqzla3VDm4tnpa3oPqy2
s8kmiZev8j8PDnoQLSr+GlLxHM7DQ1XM8Rpn97NnuAU21wWx6LhC39I4XQ60
/eqXJcVb/juDUx9cmB1qBnCQkgMuQ1WMwlwX1oJNg6cpOG/St8mqXSUajDWK
vVX05SPLNm037z47l8vl6gZ1AfGF1KcWbTMvNVu+0N1IW0ff2eNN5Mmfa287
Bmov4VSEPwSA9qP9eaHnO8f9ZY3TtoRAFJh06U8H3VTQozBPNTp27KFHmpcE
cdRybqB5kqBXVdNhPq5VR+x5lJEsGNKDggtMdHNa4TkBmmYpBnySxe+f+0Z7
cpzk4lj9lHNbOACNziqJW1xnjNYM2Voj6lKK8ABtsfxlFnDC3OD0g32w8vUm
fDy3hxKMpvsYcq8lsZax1jfahnatgU/b6DW85ezfEx6Yo0jX6TRe3bd9tZ/9
LiexjpWwqhDToAefJwSY9bZfOn+cHWzV4QFIMEoUa9vaOlaZV23/Czk1bGnD
O/dkznArBvUUwNuKXLNVrpa+I1ThyfpH0K0GjXPp8PSjB3LtzzNvKvf6jIYH
Zz4ZCifr23bBADkM/1/uXkPQYj3RCck6+hwHUziry01+KzTkuA2BPCyREjId
YIEA+ViPjvWMh9uNNOju6jamhXveHXMaLLxMsiFS5ydq/YFZGDs1vUDn5+zf
jt/4O7rSpArWMmmiREHfit1uTihYAUH5h60V8y4f+Ec0blI2vnDR0P8zKEya
7MXSCptBd7zS79zGLQX5zgGqZibhzZB+u0pQvmM7SLXTP5kdM8qZVJBDkgwn
BQ+nm54/CJn9c2QTnj3AyRmVB6EhE+timKCADAvJLiga/2V9XxS1zLyrXQu+
UBLXtDv77pG9ufr2p7oUH5yXKjD4o4tHW+9nijH9rMv5Miij97/nxqofmTYM
Zh6THm84YzvRLBJEvk7G1tjmHMjV0Rf37s7R/MPAQGrEDdfz3Crat7av2O/o
oBcqeEZgiJG2biBPUS0OGI4mbneGiL0nJM+xxrnlviwlqLlwmFI5PwRA+K1U
bLBxbtkFVr1o3a2RXFwoIq3pPb/I8QW1Sn8LH0QkepU8lAyQAw69vpvpeNZB
gZaLIC8Qe4ZlgjO/aJhptCCeBKhb1SOZOYdAb3W1Xzf1VBbQ46+HY6mYtDyN
q+jgBDWGWSk6vhLqPorumXi3YtSzfuKrgjyZycu1pXQa9CnaRzoJPXu+UTFy
4IrRTYOLTuUgaYK5GBIe5o/QBWqPPQiyzcytZpsPVdwgLUHOg187hWJzIAxI
8T6B7YQQWQn+gpVvQ+M+YvHpES1tbLw94DKFs8K+gFe4778L44Ur8IpeJHDw
ZSDBt6BrWP4HD4JnT3InoVi9xvFLHFQT+wmOI8eQ6/C7nt0HCfe9q88Oa59c
08vu7xhVaPBxSZLFNE7//UIPL9S5JQtXcpelrvAuvy3gal3QSHKpwFFzUCO1
mFOUDSxebpM1dAnlIsaViKH8IBWC5uG2V2PF1IdrPHI0FG4qIkjsmba2fPsJ
V8KA7Y37mzJlofdUPo3WNOqftUHSQzHSG0PpO7eyuIxKKj2WAK6VZ/ElO0VV
kg8xlbH4tevznYjkdTDhBcDeQKf8Fiu+pcW/vUbEvRJflUzTwEvRkA9TF1mU
P8V2WTFXSykwH9PL89/Ky7sdSsk682v/Zbqc5BQ+pB4BDuSk2mu/Y5h2kJWa
wGKdH8u17kNcyBXQRa+SQ03VFM4MOluTZMiEX/oENtG7Hyl3SilqWYyKt9So
nX/47IdVjrQB9PLIVIgw5YLgABBD9ENTfyaE6w2WDdzEtVoYMK30T0Ah3D7g
GqDa4m5Hx02igwL1eV9ssu844Kwemkv3LAX5qEmr02U23vl4SWBOWYSImr49
nXTHlwoVZtmPOlhkXQXGQ3oHjxLEehDU5QeM5lqX288lx9HPah7UH5IwsJW0
gnz6eoSlqmQHmCHZ99OhnPjcMa+cUAoWhdwfF46sRuQ03mMB4rxAu1bECcEL
BZ5mQ2kSuPryAClw86wAiFFZLX9IjB6PH/o2BTA/OeyiX6U0BVN2/psxpnTx
mTLjAnCtNYQsmTuT9teT+OpMU3RGKUxHTqaMe/WE8ofaWqanwiTkhcZKUYa3
3gDUD3QUjWGA1NnY/Z2I9NZeqOTB4mTZmHggZb+STAu07U5uJpWg2J5O6qT+
bUinfjsJYuOOblwzCqMY2y88cOj1KEsAvhseAEhy3WF86SfdP2LS9NSTX8Qn
6afRDXjlu8UyphyW3p6GpQ8swKKlaElM9gc00QELQ64Y/1f0HtVWtUktTfEP
pjUppv2UeNVW3zbHaYjkf3UniRwN1mGJax1G2nTazxc9xqv7rQMW4NUWRzoa
xsxCxJipjhd3c7egiiWN3SvqRMMALTlkcqcp1DsT/Erp7URlx5n2Hx1WgKnI
uSGjVPpic6F8uLLZugN6vt1G9iqGUIuDcopO2NKLBNx16tU/O/qmTKX95dkM
nQFzIbADj684gfQFVEnZ1T717HVsq1dxyP96nGAOBShIGEauoG099ZWBGXwe
CYXa38pCG5kIiMTTVoCL5f6f0Zf41wKrFSq7ni9eaiq/DmugpXXoSnxX95gl
iAJdqoJqvo+i9Z+CEGLUaB11O2/+zxNOBi+hSjCpk9gMoROjStv0nBNu5VrU
a5l2T5+5HzkyMggRrQIAEd/Afq3H7jiMBekCEgZSBhn05D2bgJetGgWnTxy5
rkNoZF+qTkOGVJq9NCnKrsyQh751eQYF95tovOlYVgVDitl9/5KblLo2ZphA
uhAtO/xL5FLI/Nl8gD4bKV3xrejHKXEQxscPBj3kB0agQkFmbr1I/N5hcnTg
5nZoZ94T0IqmeleiHzTTyQSKwSyUTqCaaTtLpvUtutmepN0wYQVY30pCbAwH
Shg/Mz7E2SkDwihYTHqIwAEXgCYUNYe6iuPikZcZGs4/l2Cm7VVkAwBJmxQc
Ed9IrGmmi4eBOoJzfcV39Ab8OktbPTIxpqxNQiThxwlCx4inanykcTzbTrYK
GqQxrnqESFiuiLfsl8n+g1UMLiDJbOmn22XqDUKIwOvIvO1J8NYjLXTlABGp
2/hLiW+vVc14hv5MJ7PMFmv+uZIO/9ebOI1pGgP2TgxXW6A2N6qkQC+KnJmQ
8crxQyKw9qem9D0QpbgAKU7vpsc72T4A7VxL9sC1agZBq5/wAEyNtDDRGbCZ
dzrWDPbDT09Qa2tcsTkh53/2AYVRuDw+MIBjmbkZsDQbpIg/lznJgwycLCxI
WV6QYOe2HGxkAdrUG52MorBP297/5z6MNkSLH0hMTR3yhOyfLkB20KBafpr4
FnZwgXIWOHx1BdDo0wI9VrPk9KYGMdw+fJRYbdOEKBQrDnj4nOJryyfdFbU6
kiLPOpqDu9U6dzSetcfCJG/OSifCDeMVC2H6ny/+rFaa6TGZ1zjnY6DPQsfl
CWREmpcQqPMQJeJWqLFETT7QHUUZsD0QF9w+08N2nzzGJeQSLXCPBe70cWPx
VHsSeh4HBmKTJawrQnDc1ZO3Ub7uS0E7yeevkUvosb2IhOmIDBzzmeJJR5wc
Lr+3IOtPjT3YsLj/EKGwwrvDhDvOC58p/Zm7lsXaDXV/C1zIztPEOScEOrsz
Zv0fMJ9wcWIHy3/eC4/avMAb0EFkUiRypF8sM1CCanl/Ch07wEQohlfva4Zm
t0Aw+FxeaeBpUPRHP9WziZLt8En97vLx96mDrNtQEQSMWz/USQXU1bGjNTuU
EkhJyo73QoGCzHypCdRD6Mg9XhHEp+mwohrAp4JSWd+9Gs9CtY7UzilM9eb0
FQldrX81PHI3VQJ5G9IB6PJQUMafJjFDqqtq5FyQFDg0FbAWoKCUV1aAfeWx
eWYmaEauOPZrQqd3iXS4D+FWE81F6Ljm3JNABqB7G3KSEMbsgMqCZo9qaocZ
CDrFR2cyKIgkI6QozpMk4scSpozV4Xr55OuvRBMouUaN5/H3UOVioU8Bh6Mh
oS5K1FdEO9fnB3rq9sUD0idMjf9V4cn0fjtDf8UK+pdFd0cpZSsjm2Gt6dPz
u+PhEmE0z+MI7IJ19U9w8c5CVvXtPoTFu15sf50NMZFwrFA4eCVVKvPzBpZB
UKtIglo37mE3VXPUiz1i2TjvoQE1UfpGJFOhE6xXwQygVbP/ddrKWVsvGnTe
FGFWLdZHfrERt4T/zRRjhpHaRyLCz8A8hpFBLvInS8aVX66DCWqRhhubx92/
OumnsKbLBY6dumDe+ULv+FFCYBFAulqzJmbx42jBsspD0I8XhTBQgbWxGUnZ
CSAOcEfoJUFRQbEOdelbAgtKyBbUJdNVX2PsHL0NYnczXAraUOScL19OsBWl
e7lH6pdqUKui7ir21hJ77y89GE/eAQ99oYxs+ZhFwdZfNnJrHjgZbOrDu2hw
wTjVZNhtc0XvA1XaRlcQBlPA/muE8x9Zh3DVGAPuFcpOAIO00UUep1xczBAu
ONdVUtHIF55Ob9GZYuX74TdvC2mabJq/eIUSIaW0gCbPrWBd2a/D4rzZzIsC
IW7AZ6OCmm8Hhct2+RAmxncOSxp6+tNs+m5QGSLeCqoAMfSAKOfjlKN/JBMP
cpftGt0TFDHOHnxrCAsH83wr2ZrwEuC0e046WT1x9aWm/B+XKxF3DEY1vciq
P2HjhewH2+dJaFVjjFx3/JMEid4xaHlHT1Lltgu9dRBkF8TnlDUc1iWivwKv
GKqCxC0XmEURoNML2hN4MbGkTozulhV3GDMKJ/3wtCcoOiK0uWirAvy8hpN5
aRQ6aaCyKR3t4lKI1K/Ulnq5/cgdgARuLuvkUconFQyLjUYUQMOzbZOJBJuv
C4OB19NGwZ3N7ku8Vlsq32fBPBcrUk9Ocru005HvnblhbSy6bMUCrZ8tYEVq
0eJ1cgRelvpn7tBiQVgRcWFrxWDFp+GdYdOAgQ/qPSyIuyVpzDQT1VtdUGim
NEcHVojYW2QP5pw4QM9oo2XFUVI/Sc13+Qkuujazz9NmPDkrMt/5dRaXQd2W
AkuglGxyNwSLRIrbAJ3g5YLTmJtlRY6ZZDRWLO70/GBkp36g/v6KG7bs18QY
fem/Bb+646wMtmhg5+KzCEGQ0szMq9uLPIJgZ8FPUddbEOE4sI/6h/NDf742
b89zgJXxLuumYJ4x1yFsx4IC8CjsqJTHRxPHBmwB5xtgHl6+xvMnBaRU5M9R
61YC+Bzq7yU6sFtcp/hlvluuXRRXVNbuWJJKFT7YzoLshDkMEfu38G2yzu5E
bf4eayhvq+QKx0AqxyMZREoKVDHQJjLo2T9CvMji99PU69KuF6xhRuJLv4J0
XZceUAWAk3Im73r3uJ2YHaTXkZDjFk4MXHabkVtjdD5Lk/XQNa2+omi+isin
MIi2vfyPcYu5CmyriLOGWDHObY0n2WvoZdEuSohRlKGk7BaojWwitoM+97YN
6ARiOzvVwGGlgUhh/0ndRkiEvBY3YQpKZ1pTFwKF3wLWVVBe7UiCwmn1XYFE
QU4m9LkYcRoNKX7UwPvk85Y8yDzSkRRFoAwWAWzqsEt/H/Oigu8GcDUuEePc
W8UJ2nY6K9JUFePLUMs32oXSgTK3LoeSL8IN31parkRb+P2zxHPSUXgHl0S8
yDCECySzvM42uukSsqRKgbeCHU/LMc2N470sg8pNiS+EIy/JW9/DGzO1rOAn
6wFZrU8x4+IorSZAADfnDgiG1fyIp74Vby09n+6ramByTtJjIz985KzV5gmv
U6VwDQq5xKCYNjCOtIFMzzUjKg/EDAupnmwvBWqESNrRm6uopYDQ4hT6Mj14
hljg5AdSMOsTRg1B3SNaSelT8SF9E+u2NsH2oBA+TKOo5nX2apDhEHc0nKJq
+fk10y7SngvGmTuP3C7rbmFzupb4H/iA2C/JrlffRezsvt3uqGXOC7Gu+biI
bYJwMhU0pavFitMGu5EIm2yU7UNpuGXJtX7pLUoacI76fU5tmCNfRH7XXLTF
FLNj5SS9fGxTuwnfHUrVVcbJHTKelE6JGfJlVXxrENaFrAmn69HWPBhIQgYV
HhawFQwraaMk/KB0vHD8IQBFrnmQuGesQQqQ/GMuS9NG5gWB0sNITOStGkN6
wAI9dYNVg95Buu4nagCNtI+rxPtIDxOBmX/IgyhoTvX9BXxmaCLBPJRfnQcE
91Cboji7j2w/7WqQPNIjpyRWLIb6to9zwNsjKeAy94FtzMiQfQ1GQiN9aF2y
mVk9+gwgXE5GFnQC8uR8b3nkVqG8d4n+lWIlexIjt9MGT90934S1zGQYkmau
nvkHkSuJOZzX96SkcMyiQBzjscmLu5c9xkjDQt+p2vNrKPkObfRQ7xrIKuP7
fXJFkRWfYkV8lTO1H+Lig3+Zw/F4FHyLji4NytfVuO9bWuEGalLzOfg0AbP/
/SO8l4BeRQdFuuwllZTLMMIBT+yev5KJ5N1AoBBZWsdbaluVi3pfUYNedKt/
4muxXDWnFkdyae/C1Tv1VR6aw97sZrjPa1ZgLqBfLIX1O5iqWMi7jXKRDcIR
LFpyTpgj32DugKhyiYadLgn1lYmfQgN5Pe/LFVsyRJM6dSkcVEejy8ih6Qf1
C7H6CtDfQRakNG1AXi6gvwBzwAZEFTWPx3GtYGLEiPo+2vf2QAFHQhbDy1co
h17GRYeO1BELv2i72Wy7uqYduf5UqF7PJGLcVQAGW1TtsRFSQZdMeG12rDvY
caeFM4dpeyNejsrBOL8ayZb6NmDukIAMPyzA178rESdPe2075WIjPSxZNckP
vJ6UP8AANGvc8W1MKPA1BrEsSpf0bXAgYmV4NFGABUZaZOjPyzYlpCzOKpjh
99KDQYa8bwm6JVNJdt5Ot0aJHDNU/yLA67B7aONcNWgqqqRBKBXyQZPsOL7t
FK4P0KXjrW5ko7Gi0X5wUHq2ikqVfdzC9HPfPt+TD4zr/OVuui5jb45/DPbk
Y2fCsVZ2soDo2jMxSc4Uz2mUFUIokYJ0AJuy6cjCmIuVibNSdXJK/S1Ve7mN
A1BE4kY5kCTwIfe3cQwwKv4OonwTXtHfQWgCy89mZZtjFUs9JLSLCzouy/JB
r6AvZC/OKmsG3+nrSwylV6cWUARIEBAJ8TCPkzrxW/qDV3wNXjJffs84zFKE
nikvSYw8qE5sRYk9ExWfICXwkfuZprab24BtyFR3/XmbtkHKaXqcDfDDEK+U
tNLSPzSS3p8hZkwIBDgS0BBK7vOhy392y0TL/V7s1inW/k0C0p+/7UXJsw3Q
UWWVWccvkcURTyYdvnQZXpzMHN9SSfhqtg/iMenV4mZcRcuTrTIVB8xyrCym
k4tlRtpRCRmPtMZGob9w83UQ4jYcxY0usFa+i2GX7PgXOyjIw+dicT2hqXRa
OAckSlAFpzPnrBTsmFBrwTPn/y3ldd/QOHgD+nrdiPpRTJqbhfMBqrUZvOOr
aztKTb1nxX6gL2Ko7739HM+TDIkwGGCuxkK4iDFOa5j1sBGe6mmHjhKK9/8n
4T2jpYg0PtvdZiwx/giH7Tjd4mHvh/5/x3WpTGeykIejNHpmbSSQaHukRizr
4mMu5eJjaivTAquao2jpO+rZkWvu6Eroa0MjwNjLRIChp1fPLmPCLVmkXRIq
4ERw64QYEgeWJTnIUaSAUlmw2vto1H9Qpco7K9LmEuT1g3Gf/myJOqZxzEZX
l8/mLd+1yTrTRwOy8Y8C8mCrQcPocfep7MQsCI+SkjDdQd9P71X67oRKG/xT
pNakRfypiIcZgwLNKdvYw/zQOnTTXtELJxVofHOCNZvhVI1KAzHEePR5VY3h
uH5caMtaAC+i9UNvTfsaZtlup2L73wBW1f4XYrncrPdiqbtOA7k2PJfNJOiv
4MsHNCl3piQtW050YJiEGBoakCZTXxg5cqWVLA5nGNuQB+KbwH/v5tb27Mb9
MekF68tDzofapEvwhGHPUT+lattlgmzT/ADFwfyoGSeTx8EEyqCeqyFg/Q0N
zGGTe/nX/NBPMLeEHFEPRe/5L7Yc9vRVSDUhRbV5K7T/NO95kS5GjA0gN+R0
3gHxD1XRGyojAof2oAeNcBmCjgRe88d61D64evUnOhy7oe3HSQFgD6hOBbTa
gTo/h02sXi6hvXk8VsoL/aAxY8t3Wk4cXlyO6uJAL9BtVF7jrEH4sZdcoB7z
xzKAcKJNSYK81hv13c3YaIXFXbd6wadvjkNyJvpjdIuXjVR1d7ZEIAi3zXoQ
ofvq0AsVAeyFNFoomXDSg7ZO4qk0+D5Aw91hh/qdVoXG+GPkS+A49DH8V3ss
kRE/Vm4B8WrrKad2DKePlxfKqg/YCtZfNyP67Wuyhrfgc90sqXvjdvnnKX6x
HGokL7jbEOWnyf/jwy8SlGlc0nSfDbexCl8Iguqnk9/3xtoNSEUWm4AMkVMy
wkXdMCDu+FZziBlYAYIX7WMvp1WxD0GgUfRLdlZfy1U574UldLMT6W4kQZKo
7n2uGSJicdnfhWZ9ZQ4fyErxAWU3x8Us/RGRvuNPSyYA+UnayFS/B+0psdG3
ndLGBtetnmgayYLZ79vPhSpHK5oyJwfsCsGM/hQZ0zpSrlDiXM6FDSGXU/oh
WJKHXhRXaWY+LY7VeW1jYV9ozv1N+YZvR2VmrxKAHYIZ+UpAC/HyMtf/qkRO
kWx9SSgbQEJDAa//Dwi05/V9wxHxRbOote5ghUXJB+nuBHzqejri4b8mrXvX
+BbQKryiXYD8m/PA4Q5vIY5sJY06ZzXn7cL+OmXjwHpW1BqjahDqov+/1H/o
kqjOrLgjZumHpkMKDyA2ziBiAySsO7mrf9nAlLfD2BPXfqPhtIzfKyAioIOt
8Q2/+4cH5ZEXBVUfZigJYrXAw+ONzNN3HBwmYkfXZb1Fn9bJoceRg3l5Ix+V
c0TB2uDZetL6rHeKADqOm28Nvr+u78gSgSv4ymCyB+6iGOnykj5kEBb2UdB5
gI/i5rKBaNGhoqIoRr6FFRNFanEob7363OS2Jf0f4FLKxwc3DhBc13PKWr3z
u9oLTp1r/U85pA/hLkIUkslsXKIfAqFP2jXZBA0/sYWopeFGdGKM4Hd4LTY6
Mm9nDCtluxwlSbHVylwPkZVXPj08v42dcscNdyKWcCWjc6U5hf4CPpwV4IWI
+20RtQi//j2zNiKSY8y7aVNj3Fq5vwnWOy2KUeSiC+wb+Y5tsGX0pskNw5Hc
kCRuiO5fWQ6gPLyG+YOgnjJOvUANxAV3JW/xVfRElRozIqapnkdMWg9Exr5L
vPD8+eB31hvV6Bm5LrsLcUy9piZmCPPdKyzhuKNF/0IRBEGTJ209vuTVedAh
dKY1dCa7nTqM3anpWhoyMjK9+gMQZ1FpBkFCTT5hemADiQWXUeX0RUDZDNDX
BmY7k7etQkdQFkTXHmYGfSPADTsZYauLXXkByAg1mHwDCpdDBa1VU1GVPLNN
Scbvi4ET7k3Vvn1XCa0kXAUuQOrJvr5C2htIXsqR42J21pTRTw9S1lPz3iEq
s+U2ab3J6EOUFyVcZSthV+8U5hyEANSZWVhVnXkDFRiqQ78BafZG62OP5C0n
xP8i1ajljvbXnpiIOIaFWmWnp20Wexc4BJD+WpoKvI7LqeLrf4sU1PdVHIBS
y+YOhzXg31qtMGZshP8oFvJ3mpujFOY5/t0Sr3/Jt4E3j/DARA7ym9o1yqIV
JjUitsfQTJtPHZsLXZ8OP2CW9pMfrgAZhpqX18GoHTFm6e3dRRgUCQLz3p0v
/O0yC18gvjdfyrtTcY2npbF939U/HRgYBRjHc0Gg/HD4NyZgx+WuLZVdmJQl
HPwVOGT7JZyvg6LOtmPRyPqH4vjy2nAFNd/lf6CPB3J7YH3iuyPJmiqoPr7a
nGhaqCD6yoCFR3NQOBO7YDSAO7Lx33TDSULQp2laCytEX6OSly/nhlLsT/6H
7/rKaTQSAmVDm8ztnRt4O361rUFo3LjjB4pnALDGeMAXNPoHa+NYnAiQOfdY
/hKYF6f4vis2Wi+YfGbkH9ljhCv9eeQqkHtrIt5h7HweaU+B/hOcSEGoupd2
YpeoqCspsldrIvuqRXpjy8m4eaDhvzos+Pe3dAbNKjGyiia3kAQNF4I427gf
b7cse7eOD9FViQOgiPkNATgIZE1CGZVshjGHSPL+boCJ03QFQDgdDGIDzxag
x8T+EHS9G7fNKu8ottohzqe8+kZF+BAJs9xS+lbnMIhRZwwcsM1n+ZYIzLod
IT86/Hz/xrV0oCGk9R8Lwuz7CSBZhGTK1WPSQ9DMDqgeAaeY6TEEfP7VsLd+
swlaMVBHoRZd5Yqsfzxrc15A2BdjC+3KTQWpKos5xm8M3+b4Cj8Tj4nUpi5j
lRT2t2femfY/9Ks6oMU50zEx0aHNSD1jS7I7DhpAZfnKOdFot2qozY+PccAS
LCMO4cNP6YhOT870iYlQdjL1JqpvIxfBN42+sevV44UFRZxzzyXQxE8F12ui
bGb5+Tfze0+oZgtAPkNutKj4Pb2nUXjbNkqTcgDmVHAhMyKtql+OAR9G1kwK
B1csp846iQTBHvl/2/8TvUgrqIkYueg9gqyCcycBSYBw9gcEyvH0zAbnWiZn
28yZtyb06jiY2c2letmYeaVLITYkYO9h8gPIdD/xesHhugVbvIyS3tf24+g2
cBYN6wiBBEPqP2yG5SQ09zYD+049QrRF57iPL6iLp/OhIoNeGnKBnzDS1P7U
yTmn8J4hPhkpksgCs0OUwRG8A2gWM2PNDi2AT39J4AI8TeV6w6xm126u3nDg
JU6pJOqWt1MXoamRv838xTv0PpZE73VJBwPCBX+G6KCs1KQqxScKiex9qK7G
+bsL70LR+nUbPzYuF0vniAlQ+vhOMQ86pF9z0KnTMvc5wyYmUUMM+7VSI2ZN
NrvDTvU1TXho/umck56baKheGOoXPPCp6WNqWyV0Ci8ZnlpzsVezrF1WcHKT
PS1B45Y4DDXX2GDfILRyuFZRTKxwbDo0p/0t50JXuxhSK6vbWpPUNn+7JtRL
SfFq2GNKCGqBCYRJdreq9+UmNxbrWgULzoglnz4qZ7hw2S5VtzONHKN2QlBI
2SVTPWvHW1zSlj7mMRIPcJn16sp8mBBc9uN8u4W0zOjYl8zyLYesGFrB8i4W
b6QqasG0GCLPlPDXVy2MAiWN1RPyPxPRGr1muE3Ib9PfnVfuCWHtmYVndemj
yEMHwYDqX2eeCJhznajlj9I6w+qmOXkY8qXKZvq/sj/nqvQGZ7BQ719hFXf4
ivgqKw9TM6zgacaWK7sopf6Ex/lYcGP4+6jTG7L5deK58WK4PmmFwk1SPKBd
GjJnHvqmzF5EAGCsxSg1Qw26Lmdn8LkxfQFqsfL24YdtPSzPPfqR0mhQakLZ
ADr+7L5/nh07yVn9tpLz9CvmgL1U7GQdqVLCWFyt2LSe+BWl7M7iVrj7bsjv
kiEKLDjsIr/tWNGZQt2hxrdr+SMPvMsMVMKH3LWEjel4SAwLcxveNkKS7hVm
wwVLjC66rq2knpBCiK0Qc8zpVrSp6Qg/dn2jjabIDGYNIi0JeM+0de8f9vzD
pmcSNcJVLpdf9c3v2jI8xw2gz6lzrWygVJcv7AnbK/guKA3AxMUGx887YTC9
On9PD40sSBH7FUPnJXLGkelHMC4JKBxy4wETINzMxP1Z9kgjU7ZPO3RdEIzF
8R6/uKhB98Hzg3ylJfLhxbTPeuRX21g2Bf9lvlopxONS+YQZi394s0oLUm/T
w8vZlZwQjeSbt1cbelGU3TrC2LHtVH7I47LPfGwqIQQ73ov/YroiNiWs8yza
hB8ZRAI092Pynjh5DohrmClb810sqj8BKAjKUCBFIYLy5N4+Hup7tEDQZo4P
psfanbBFHyw3T8UiAo8ORH6pt1oNd7GgpBorJTv58jew3cg58EuIve2sz+/u
PKoaPOKEwG98mixmOnJUKvEW/byjVxInFiJZW4kNDkEpqFlP0Mmfp3N0K6r4
81bkJ/XBLGaAiLm7++oheS09jtQDPinwmUgPFYlsHva3VPXogoocV7td6+HS
P175/KnPdh+9vG7oI9aULq39kAU1pmagW8ocQdzzHupVW19Tcao0iprbPUuH
oxDQw0L13LK/5+rhj4/TNU26aX6YLQfMH4qE83/0B00Xz3yHj/JWJi0PDNTJ
m9OsAVZf7fvDAPFCGmZUEM2DRtK/6rV6vcHFibDoHY2e9FrbQAEbtvHYiPmG
kqV2/AZrR8eV36bP223QeXYkl6xhH7zkUSvHItinKsbRydTeao3r7dF4w8ga
a7sZDv7ZoLDkpwqxiKp9Yzwjx5LnjbC/JTneKODUYeEpJOrZSJy3kpIKm/Rr
nsD8CKjMBdahzedJBD8eBQ/ibiZEQZ3nOcVoL/vBDf7Q49o7fGIZthMSspy1
ZGnKmbfMcWhpuL2oQVgpVU67I8dDukZwT++zHtn1ZvbnORcArpuGccoU1idf
38SisOxZ2OPRr+Pq5kNdYBicpdGy5DHLEgDRoc7iRaDjqvYJ+Oa957Bzdld3
RJdab0ueWNXH2Ok2063ttLtw10FtyPy0Yf+pwvtk1slpEiz+QRgGleG8JZ8v
FwNlfvhTy8CuorZ1N/8wMpRMDzD602BfUu3f0eerMEFA0k4iLPH7GX+3bJt8
aOiGppk5350xgiV935X6KcroLK2Qu5o2cD0B4nx0A5ufmUnHHI4AmoksSwfR
ySMgSW9Xnu+Vzf9hBkav6dfzPIMuAqXVfXGYyvJ+G1Ig8irw7LtmAHburbT1
q9L3V+FkO+fLcn+kwHGxE14hpyZQBa7P380RfOziVbKGIcroprFjzoaA24Ts
rUNCBFbRcYdQA7SnD2o//81xeWhhA6yz67DFr9IWJxll8d5V0rA0sEJzOSik
AL9AZfFoxZreu79ikn2xL25JUwKOUfbF8hrA4Vj9RAtPQmrhw6U5zhwaJW78
7+2N5AhRfjtDKZ/OJ/StF9//xjA0P5tlhv4SpMVZIy05/X+l8NqtOtgO+rUF
xDeHr3IQcNYvx14yYqmMFN70EROflzD6xeVx/iM1AfT2oDQWcalGqfZDlpJW
2PhbmW9HB/Ecy1k8X4CgOgAgUS5iHVABnG11J/qasAHHMZZ3dHT4n8Vu3BBP
OHGaUpSDOC41OkaDCnMTVe+yqJdsa3ZLspulL/9CyUrfHrqJZl9jENjj5D74
ZjXUnGP8ui6MCxFoCZYqHjocGktX9/fOhFsuUuJUfgn1iRY+RPDIDEmg9hXu
cEfpwx4oVuYMdmRIqVPnfWBVOVETpkn8aaTKP4d6lwbInSu0RqWq98MPy4aJ
nHfsxVXblj7MXEuV3xytu3FL9lrlRj5xUMSARlOZwWTxEzN2l7iLWHYjTqOO
zojBgfv9HSWvODj3ntDFx1bS0ZwA+rXMnAwROAdkzvAHZJugdnFbesOffajY
foQdnudhGdzp546AlhcQC3bopIGLYTvqeNBNYO4soAFOQOwZmhAf6MB3ZbBb
kpNpQDvU/oS4UmF5MD2tT1Xblw/ch7uQeEFRYAhjULcAwYjY5Q876vLLSwGE
6mI2F5OagtdebffqbxO6oAzde4QuV/QLV5TU2w0zeWieeJsPVffHqHD7SFhv
DjGoXnqWuCNznrlIMzrz+Rqw2HMJq+U9JAK7iDGqGlQBxKS91tCNLxW8q5Kt
lTWVuRWnasJSUzBPgetpIYHEbPbimcQ2A8UHEMTTkh8Dt/SRvdXHVaFtAlX8
nZGHcVDKxatBAQuhUciCi5UnThUwcNmKr/2qfiFQpkSJXGQTDnFB5z37CEw7
szQVruAr5EllvI3wymRLpJMncL06bX3uboJpYE95/iFVGXyRuoRzWWaU2Beg
cGZbRX+o4yxIDjSEB/3AyISgnKb6q/XZZeYHoPfk9TXga34undDQRNqZ9n6Y
77rbBp/W6g+WQM7SbB4md/bhSYkXcJCbHDIvLJR84exZZRUBsG5ztumjehsc
f1eTJ6hhnc/GHRpeitAFa/nDz1pHFFTOSQ3OmFPqEBM4ucCS8SYylYEmNKdD
jSsQrwIhMwkStpkfpILx08jtgzRbm/miLXWGaPRdm20unbPF/BEWNKMq0Hgi
Ct5+cINIUorVR+B2ejO/4H86C90iSsUQfRptGRNS4/6nLNE3EXwNLyGYoTYF
QVQx6BMt/lMNb3shf8n06icVeqibfdnhcWmrgPJ9orVTPV5lo+Qyqu/D5nnQ
BNwm3sRJ5pg0lkZGhVwlQsviAWD9jOH/PUiANeFCDTzdKHCh5zv+/6F5yz39
Jgk9kzRqw3ym3RXHPX6MlMBd9Lk566jwbeFOG1uPLyZeE6kZgbZX0Assf0lS
QsaBuEPz+MSCvBSeydJs1suB/mRO1ie0RdYidLdUW+yMDeFJ2jY+XOlGL9nh
7dTA0aa7S35QdH64MEFnS2/Aa9wuAiYJWB+QUANtgk53tnAce+ETCOeW4H0W
c8k3813+iY4AWJ7otYPNEqT5CmjxM/Hkl/Mlj7tj8Ob3SaPXHrbVeEVA1dSP
BDcvWLG91ffVG0xwUt6fR+DguO/leHlAi3zmw+PhAuPpRs2EQNiny6gwrwnQ
qdZh2TzGMunzGxq/QgwDwMJaTX9Do7YzHVAJUjFpAxL8eeeVF+WpoBs0Xbvj
tJ/HBOuWo6Dsi0ugKslz1CnelBgdsIOZqx2arRGqOk1nz9yd3unOAVQ0VAqi
DvcFQ/ywmkt7DAu5vC/pahohyy7jprulxX6AbKp/MryiCc8Ok1kxnejnxlwI
U+aKYUjnVsNaMpYbImyCDot/13k76AFQDU5zjFl0Gk2HgJqFO0YvS8PFtVPG
C8oE4esePMhcVwrnNNb7V4xlY4BVvqW3rIQNzAFXCsmshcgKG/mCF3VvYX+5
pwEXjvCAd4EF4jOzcDG6E2QhpI57hy+lzyej6hf+e0qI21nWUSklUAa4mGh9
SeqYSJj7Iel8Dyba8ji35jxFDt1oxxVEFg2rEmbLreCfGFEgU3qCzz5trTbB
O18c7YPy84nSC+iLgk89VtwUoz2vSabtttw1EVJIVGQq5mKO3Bn87+xdT0K2
UU2Rtkw5eASKIsbbu+r4sL4SD3vm/7aIo706FfPPGWV/tqArQc0IEVl0TYW0
kcw+FVKJHoPrRZv+L3jMA7pF7DtzxlYlKJ02EvRHMwbqQFSVi87jo7XyvKB0
eM49+ZDweamhBOzysuIFx/a3pp3UAXG66d7cHi1+L9HlUdNNTW8OyPqxMgvn
YgQi/g3y8AsrnvFiLLlTFNeDMVt3P8gx+33pjPkw4lCqpxLn857IGYHGQwmM
YsRYiwcTid12fjsMx4FCcVy7YOZzK7YwoB3nOBMqg3oJDPFuDqBUHN8zXO3E
UNruOmQsJxKTaLHiW+GvBa7N4KDBOzVDmqSsn5z9bLDjuQmd0n5xnVy+nulV
gC8l3fLffp0pGV74Y/dgGDFPp0xp4k4TGOUiLMMvrr3TrfPymUmFpu704O8M
3RAOtzAdVwxfz7FALm44jU9hfYL0x6YUTD8JVZtVGheShAfaYNfaYtMByco9
y+eJXX64Nunl/iKa3ih/eEbGqg0BtMXcgKCm7tU8TiyRbsQLO/9eefeVlmdL
yMJqlnMZ8iOQLGGoRdh+p9rCfFOoZVKH6YcUQo0NetUktIdwntfYvJmbkStf
c9Ed8GpwDYmYKXc8iStkIJ2UOEcSGYygIfuKxa++saqTqx5b3aQ3dRZ1BTNg
elsMSGFmAgLtJX5XqZZI+MM6hBxAtknIkXToPciIaz5wmVYiN/BKwbRMSODX
E+zmd3HIfZujOkmca2Ezniy6RotVK/KjEcHFECYj5a2wxAJOYf/qZ8YLtWM4
S5d08yYrLBWk6YqQpyh+4RDZ/97CabUo1vwRBQhC0gFQygrK2GMyQL67+nde
5ltIrXqfoBXcYoqZa5UWIGuqCIp3JdQfFX5LlD/LJhZjW9UyIKsmyzOG82+1
Jj23ZiortTunjtcmFj10ibn4CVfwWiA5DtaibIbS0K4uXf8j/LZZq7TlgKpf
MkwR+3OG4e/NEgajuO+68Won6pRc3e0KD56qzVWhYaetMxbAYTHSrY5FEcmp
fmTUO3olCzwwfFKzpLiEpliqK782BP2EbXFSCu9kX60Vc7x6V2ryafxY/HlE
9DJwPX5OiDTkr3Gm3fbEvUots8SniU8fbtce8rzUR0286o4Ae2qPUYelUIP1
yh0aQv9/csklFCVSg0h6sIHnxwid3mAatvyNQbW7NMthZgDHi2ZY2u8ZR6iG
gq5+w2zUv5QMe9Krt/ZhH7+S/iJNmQaPX+eKpBd0JhNIzvAzg04w89Af/wC2
SsS43EYLsCY2d+wcUp2thH7ZcMl9lolmrANUjy1b83uhTzJ+XG2Q5jD6NMO3
U7GQ5TJL7rhgRauk0ryfs8rrpw7B3ZQphBGUIJXrRJLyut587YN9ANZb34bZ
5zDoYV4W6d+D/VwwnRCtLHTP7ogCQMnjDJv+KSQJttgqtwBGzRs3I9ARvNrJ
NoLa7pnxpUvtDyd2jwV2RWy7J4PrvvQw1Bq0MApHJ0g3YmTEFfus28YJ0gR2
USBAJZew80miEAO4KGXMsWE8RAgTVEGY1tel++4jn54TC+ydguEuDZVbV8I8
+5gDP2rwAYYaref84dCpMH4Yq7hbVnAdklltSwZJEHRIWsdQp3O5JRl9d+8/
7rr2N2vCKnP0etA1h2vPMTqtF4knnmzyFh2O+ZoPiuWfIZvldG5rc6iKTBXb
5YwszHT27dIAVml9lPPmI4Aev3TipvQpMxFXJXUxL8pmJViQXEy+RMmQ/dKf
ob6FjQDtD59Hegx1K2IU4fCbCIj3lVnNLTANTs0hqdpECkY61NJyYV2W8sOQ
NT2h+gf+uRBjHlK3quqOGblAa9YN60FXymg2RaZqyzdCxtnwv2hDDPeTRKZI
VXkmifkZNE0PrGLAQK/vx3OWA4SWyYdGszPbpVEpz4KLr95nmQrpkxaqpIZR
ipJGNmcDls4eBDQsTb4pVtxPp9kxZ2tt5JdOpj5j69XydOhWHzC66sddkndH
omcBngnZDryKt6Bbn4rMsyCk3pg6vOtRIboKA1W31XuEbL76w25yi/aAGpYS
KeiqNB2ospBAvDhwQ2s3nj2NX+Ss4+a7bZF4w8Ivj4SOz7yefzgUgW0zGj8E
yHkBmMBRxtoZEZDoxHdQaJoM0AaQwskolDLD14yh7y4au6O/XcqCyKkRJK3O
GBz78Cnmm8aa4i12clxMQsROe9tKIXVJ39CVS01vcNxLFzzgmWdLLhGVIS8h
77t+cZmDn2IIWnZ2Xo0p+/A2qMMa+MPr9mDmzs2SDc9Sq1AJyE/xv0Kg7CYw
OYTnrm6uYjRAHRiTAWI/qwCqDzto9UYcj+OIk4mvEL6cX+2XYym9tBB9OFsM
5VCGfYYc4X0X3dpJpPQCl5DobcOLAnMbT6tNKOg2JYBC89gBvKfSSYkSoPPH
keqqMY0bKD1RoMnXMmR+g+UQCyYGMnUSYCe6t48aeGDdchOZwGy3aGEuQ5G2
5JIPn9eqWPqtYTJIQ1DZmOevlAD8AacLeK4QSRRiRbrQfzdxBU/JXr/1yYSO
VDoI5BvmE10c5Igsx3wrfPTO9TaU931HglnbAN5EpW+vI1uu+EWotJIXcD+X
Q8VE6nQZa1NA1klBpImcbjUfhqIo+d25bG3WVFPIiIcCQIJ7X9Ub4rxEx7Li
rCFTPMU1OEo8t66Cdc0sLShVXQOpvf+TjxugGqy6/FIevru9glAaVac/13Gg
JUnAveeqh0k3oQ78tpwiR58Xu+zWZtGvMkKoEM5yjUSsHtNbBr1E1wRC8eFr
xnr6nm0La6tBUociPv1TtNOB1C3QBIdYAI19bQTP0QHWJQAGe+GbUsTsvi3B
+9+hBrhkNok5yUy6EhWGlT8f4/DhSWe1Nh1t6XWGhellaGWphMenGlv1Vd2P
6NkyY1a/ED0t7YIzZUb0GEGC4ymkwFV56Zat/aRuwuTInFirIyg9dCcmzznN
ICJPqSkAyDoAWhDqXIeKQvCl1sEieD+v4xsRzDddufPS6vEBC2ce+VwHgfpE
0AS5tgsCU50GiQ+w2gqWdQVPkzS3I9717bx9ovglg9EwWjq7m2xPD8Nveq97
6MtXQwwSDxRa6/19yb0NVzb2APPXIMzqivNtK83zbs7HB0Fs6KJzScnHZCs6
W5QtlZJFnCVACHA20vXMlnS2vuzqQLYlC6zxAlB3ZNYyOtcV/oyYIvPF3MpN
zPMst5w94nd/4J96NgnAX/jUGRjIElMsxOHHbjlQWQ2JDoZQ4/MPJ2zyPt8V
eZEXIPe57qgyt2KjYCdIIqM7LZ0F9WmMsXMEFFDPUbNFGtw1U/W+VlidPpWA
iHwAW5fdJFr3XU81PK77v1hnIsTiLRb5b+pvGn6PNXNLGq0QGdeswYFs63zJ
tGf9gG9mQaQA7WENsitzdovIg0t5kXywFiS1pkN3cByk14bCLJ4irePlpmlB
qLc+zWk0Sq8WU2WySMqZmogIgGOeDaJswkGUXGFfQGTASifi3UDqMKVo4Bpk
6LJMY8giFX52P2k4eXEZHdgkAkxVJt384c17AI0J/AHjT1Pql8XP0Os8hQsE
cgur18nbuIFHLcz6hq/y8+31C+NJmhjKVjGRIStk69D4cM1RaVs0MKHUZ8LS
VafBE5JhS7qCu8fqBPgebaWPPgWlNoQ74jtVzjRY84YUT+U4hFbh966Tt51a
n5J8muguKeE3I2PyJ2VoYK11TKF1NJofs6pYITRs7ZzwpL7jkjkLARKAcnvW
2i8e6DHxQ+wNvxqhqrw4a1zR/m+j3ZfhasbejaNKg7BEZjdKniINpayBU10F
EcdGiuowuWJmrUsLM+5fS+OEBXe0xzj4apQ0Pjw7p/O9HInWCoiYSvlFh1Ap
xBqF8yNkVz9Y80OP2zXIkpfGRT2stEkM6xTrPHBsKal83XX6VQoaTF8RtGnA
iOd9IPagpiha+E2+7XVgf+W+WGvbNz7X1q4ZHxOgXtbtl2T9jo1pJPkUZizM
kFCLR4ve1sOvun5e2rCA/2iNGj2dl0ai9SDC2bHsVZ3NH5aF+Xr0lvXcZiuc
1NNuwmsxtjwbN2DEeRNXEnXKVLeULuXnkUny8xrcxBwo88g1lDp6hDfUBEmp
VF6iX+XkocqIIzrzupE3MpUiiflD+a98hva3MhYUc+Sefx+/diLOVFraNNh2
0gSYW33+1fWgddg+C1XM3c11ixancCQnyfWaM0lTx/qY2mMnAFmDObYdJjGw
OwD69/zlcPr5D4eyY0QKB2MsR/vx0/54pvt8qHQxrwSs/Jiq1RwBJQuQkOl6
VptUFQKmMe42tyKzwpWPMMj7ZWyZ17ZHS1O5Yf1wQ7AbOk7Fu/X64BIHBz7C
6oWqyBAXYTBxIQ3Qw6c1cXJ5WbwTKH/5clWFdtn/uRzC+W2Amx0HUOOySJRf
bQk+zPNk3PWjW+eIPnf1czlJJjYpJGdZF26Zk50QM6F8/6PVjnfwTUeYQygJ
2rSs8mTs/12N/pI37TmjRexpRxTJh0sSUZl0tVfI9VU+zi+EkLBxCKg3FPcf
XQoxSB4ol6O3A4wx6dKY1OEM1E9y8L7DTkyAXXR8wIUrVFKOdMtVu/3807Fh
zBFaSAfocpvI6B7/NP9SCgdcaHsQ/u8xRY9vxE5SZ0hVAvo1ZkNZJCqKHhPs
7UVxlO5bZDlcDhH6AgEJ7wj34hsRwgweaesKg3KlkNGgRZm+nUVAlARiWW8d
nhTIdfRVmRIvLBGrvYZNDsKUcWcyZp6VuGn31WMNmJfeizS4nGvgRZwgcQiw
v5Oon7sy5MPtaU+ELCdPQ/EXxsDQzK1r9Rjjz33vIQj7AIUvX0/UOP60RVjj
oGhSFcgKrL/NdHpwOuXr6sko0rxQHOBcnFlFS6DOgfw5fZNaGD8UB5kPu9jA
R9X7+t/1IBLC7+fAlxR+i8thO0KrmOvW0UAO5ZNtCgr8ATq52MWKKQwm498A
IKIwPsTx1k8APQaOkptb7h5wu/vpZg2R2xsghOK5Vw0s2KVsvdnF6bRxZN0N
ef3/ANcEgC94d5HiZWeI9sJ6thIBK2WWCu+9TyD2tOg8dydLsu47c6+ooiI5
MYcpMcrPHx9d0yISjeTn5Oz8OBRlqk45oPN22vl7dEnUDrSyl0QNYjyHkXN/
oUet+KgMXUehJPUG+rRy0RtBoen8oBGTdVUqac8UTZwNfoAgJDvf2B8d7NdK
r7gSU4xpMO8m2eP+x+ySf0nK6botRc34t0nPuSgoWpBlPp3lEetr0EBD89nm
mkJGQ53ZZ1S9S8lUTQA9meNr5ook3Ya17jEEVhXyPatDOQBhHtpqdpnpnINL
rb80degiTNxGKbGFqm8yCPR9xOy3jEq/Js5bWE4Sx82X7FFaueHrniXoRPGS
T/v1Go4ktTtJPEWFv+AVrHCJ1rzaD30Js9kkWJdvUwUkwLCOwIu3h5GaJMZL
21/sW7nA/DZLthPITdQr25KMg/zXeEYNJ5FOZwCFlICMjRhinwS1IIfzMtv5
FqL2isc0BZdCBpGLrQFfz4aDcSjn5sztkpeM/F1cAaVst8Q6KGn1xzO6ECDf
Zf893nuWrhLmoomx1yKI1yDoAIlNjS4B9SzugXU3g/I3WBosiGnrSugaaT/f
Pty/AiOXaa5t6D/gqTX99NwnCjyW577BPnKg9ktojd1ocJtE7HdrkjR7WuZi
o6q15Ke3zRGypeLCR1iyzh5COtOV/U4PcRIg/voUv/ysF1cd+z5FTW6p3VLN
2k88qEXdVfzX9iEel/cW9oWietcuCFi1jZELytO0Fzj9ChEZXyZs+OJClSY2
bpSIhDuwtrBlqGOlV+9JYIeRcMfUjeFQcwyyBZsFxux1p/nXNpOzOrgkNWL9
Uynh70VxuTY9TzOODHMWDHrQIcvPmIkcYlR1IPyXA1yzuu4kdiLGFSjNEiEo
fORtyq5CmsN25UEHJd/XlHez7FP0jUQpQDK7njxPe7LOmpHq1uR6WN1TTDTr
psXAy5IVMXnDZW/jn4zvinLl/iiroOhbV5B5qnW04HGgNDiu2BE9GKQJhLKL
yJA41CZodY0n+ya9YsZjNZ2oWEfwScgRWnfS5AAbK2EhAfF5vsM1ZpWURzlH
V0ViZO3VF35Yz+WldS10Av29CI58RK+1A7+UoKkHIDOUAacHWJuVDq9rvOAI
XOJwG6ZksCQPWRtg4g2JiBvSvFLB+9n/wCsoT8rWCOnAe/IhEVhM9qv6/b2F
x6H0qbBqZfdiggB8AUvs2nMCDEUKy0YjxQetuVYXMmbZwtC9is3muAFn+GKF
zF51caOWDyPXkdLzOAhMiyl9RmbSFeIyTAnIGNKdTJnZ5x4uFoYBkdAdohUv
NpGidjTIFM6SHvn4rm3SpG6U/W+xe3b0R7cJLc3IX0p+Y8UlKAjsN6BWyW8D
FAIfCGfAtFYcMYk5Be1uvc0jPGpqChRJU4rJgc09mb0ysQ7qQpfoRdcKXnpb
jd0OISHzsRRfuJLjJBfOSfLFZUW0rZa6TPB4upceFxaigWdT+fdrM0Q8I9v/
tBfx/56Y3DTK0WD5cCi0052CdoPf98YqakdPp4L2BcCP0yBjUFORNILrIvML
DsLsTBDRBCyYV30rQtYs7goX8gBxjqNOc5NiV5COj8SBF3neElIYgTigmyQU
KOS4/O8/H/i0E9qaDRCVfwnHjt31J4gvxsnUX+wdPzceuUeKxIHgg7TPACLm
94O+ESWShV8U3Vhw3AkNEfC89wz58nSfPri2KvmNeIIGzg7LCP2Vp7eh8Dck
S/AupICvwcOTaKVjDqdpemUTTFO2D4ANHbULe0pvmxIae/OeNLs7q9wClDT7
w2ZR0r3u7vxJRqwGSiZ2JOcZZnW1oVJ+WWNOx9g7nrgFmjZKFYqvwcyLfAk3
4m/+PlwXEtjR2DypRIAAEAqGOSH+ymFirUrYs4Xa2eGPN5Q/5j6s2+9K6yKn
8vpexuaeKyjHiJZVaVGjkhhdtsLbjyBQ4SU58OZhXCEeB108Bt3ZfbnNWqCS
YrI8glIRWvb7FV3meg71bdd202uV9Z1zjTkzx/1rvRU4pXxwo1X1o3ybHVNY
3+cuRzLmLZOsfTVaMeyc/12fn5bSS+d8cg9N2JrHgCAnEeCR2XmA3by3Ml2Y
YApQiKSRjLcXNCpGvwI44RPm2sxHcLXlMHb9H0UNOEyH1iBuQBp9kz9obJlC
A+AC0h+DDt/7VeyjDUrLlOBX8HWNtwQIwff84+FhA4g4tC/A2+sgWZ7y3ljQ
vyV7C5g0zFedj4j4FayZh8U77R0ic/Q+lBlTkFr+2Of990YQ+mmxNhmE8BpV
gD/q2kO9Awi68frc15xOLn+QXmAUm8gtvAzRIwEmuIrWkxzYttLPlTyv2mE9
kMgb5++5nbyL9LpMmc2WZqgu22NObKAqUP7vsuaBU3GowderReS8hJ5IUHVc
0z+cVywshRa8mxACYVJkJNBN38WHINE1X89bkffCkBtmOq4HvA68s3n3n5vm
0luvEefwHicWh0Oa6cPGzjmVCNUgbeMWPqDP2m7oX7AF+RTSaVhRRWLfdW49
Y9XIwY5OJ5u1I2boOOAMuC+xKvqunfB7LLlQDQoXKMdjyzJ6xvxTfxu58pqV
SYzZjOxEnEWtENRrAYnmvllxjbO3wjpJ/SGr3fLl1UCulpnwFtGNmRHL6Yf+
8wAT5OO0N+aoelGKqGvzTUQKZUaTpzYSTRXnkJ3PvHAk02MphS0qPwc2dW+z
zzim0m2jp1yHS72hG4E3fvlrLPS2Gw3auGFThpV/WPMx2DmQbDComgAZjEYj
z/v639VUw/CqWg/LefJw84pdyOaCgSlgyaUnNZ0RqnNZEFY5UIUNrV9Q5UMg
i0rdZJC5GAMKZAIM16+BukfLCOoMP2snNNqLVKhigj1lvICukSqvxYuUZTZl
zZl/2YtNEQQxjGcKLAvpDRSGsWpeNvpK9dT/YrtneNm9soRXunEC3hvf2Xfo
NFqrI2eJHM/Am12gtt2Ko8SIs1moIHURNDzkS3oGJP8R4h6V9ZB0k1In+z+s
kZ836jfguC79iMlfQr4UAoxoWjpIL++5o30zm3+HDQSQMTga/1XGHKSKMx9L
cHg5IfWioZw/IBDDnKJUNGRVB+JwM+GLmQR9d8yoh2DFePL65DqE+5q9XAXn
htfWceXpXpEFy2OtJof24a5lmQoOpJsZMutBVNP1PukC8cFlwJAPINcEllZc
4GHQ/WpikdcaUl8eRlztU5K5ecJbC7RuHhb2KUVNnsxnX6IJjcuAmO8g9NGf
taT3UIHr8K8dSnfs8WtKX1pv37riasA6Fs4hhppduwPzzQ/7g/vkNVS0eK9I
Y5duJ56MRm48c7wYkPgvCRKX7pkCfFBn8QdFrd+oaE5hj0SOhSvMRmb2ED76
pErp06zu0hKrgi3O2KcTuElBQ4+m1hH/vqAhRtJnqriWunmreY7VpPqSX86G
Y4DshTYn6Qye4FbUTJnEeWum0RddJuR5WdG/VO257Ecj8NiSZN113t0qEkWN
OKU9QlJzSaIZcdXJCWcVmjr8Cmg6xA0fveMGCTvRow4UC03unVq/yFTvzfrV
zyHljUNMVmPq8iaJ+Eg6ljvMHemdFc85daBL4Hmm5JtWqqwlYQ76xLY4EVZb
+nRcbvkIGgfqDEcqTZ/rtc7Y7uExhWZvZMwZidzKzjUE2PGKzJAzq9weasWl
z+u0rZRazTa5cVFrF0VQZMWECXFLVmt8Kt24/JPqdkhTpWTz4z0MTOQcnmEQ
MKQrBRLYS1FqjUXJz52U+MUyxxIhv/4S/9exeLrrVIWS9qgn3GZM8hPVZnqM
hQ177ukmg/cSRZJy95/CXFPjNGMDqupMEGMOkrlRhaf8Mxos2ajXyX2lEMzG
bQRALkj8aI7IpilmGi5qKRsg3BqfcdUWAjpxeuQSwCxSxL9pW5D/7IYxll/J
pQO3sMmo/7pQGkUCROKqMUT5V/fGAVRHZxTcrl2F9xdMo4PJxu1N8y+tP8Om
lHa8HkTDlXudQKnml/jLZzX5IehlVi5qt9gs9MJfFAePUkIJGcPH+qZG+Icn
PXK8oSMM/qiBILqnwRfn0+LhawMSdyxdvS5cMpMior3q6XDzjfsA5dv+xhy5
H8wXeC+8GSl1WZ30xnqwjh+QN917DgqmeAqBZ7ID3t2OU4loY0xWmoOa/RJN
ixKDd+WXsz8CplOK2jmlkgDUNixTf8OGEXRrtyexnntP/nalGAvNtZtA8Fv/
H3bVZL4Qd5yapELg2MF7LLg8BWzWhTzw4lnbBNSX1lGzODagaGaEhFZurwqy
yIfCAtNAhbkKzJ1xFjL1C7nk5U6bpQF1PX1+BC3hIGmUQeqQyJCCEE5uPtXv
vX7U6vs9CIJKYqqrKN3l7j2nJKtFWRbbmRUrBT0yJ5K2Z4SxNoltfDic9T/r
5cRPUC0XvelVVoJARxn2mHlkOBVAbfZbYEuJJ7Q2YV1QVyd31BEYoCxa5x7Z
oTDCuaMQlJm8J6tWQwGUFtuGdGgYGW57Qc6Tas1CZu7Hq74UpTcJwz3kQjtV
Tmnjj0jSmMm1pZu8kON9n4aD0QdhXh2DxM1yr9NyqkYpj30zAPDKPDheOIe0
f0wHkvn013Dvq8D7j5NFSVzi0DaCZoH5y5nVbRJsJLIflzhJ95sWnuGbMdTM
bQe/WReTOT9r3Ut8zHhrPE8lxVdwd20iN5mnqBqEy92rAa/qLS+OFMXST4yT
Ut6fiGJLISGa8IPyqYXNSW7d/VKL4TG0x3/xTlKj5oYUdyfwtg1rkmx47zpz
RJ1gJ2fU/rmli3Z79j5uVh5/gAaTKp6T1z64jqzZZgRZXdAN+sWxdgZUV4KE
O3MOEmouQ394PO6zGGjLdPsG6y5VBzpKGDpYxmgZ+JnSTefKWIFcxb185b8I
EC2BL1SEIbw5lB+ud5QW6IanOsFsIVn8UK78/wH9YBxnzZYwQG82XSX5xJzR
We+DH4yfWFqCUDSNeD2NdyJwldwR+q27AWjNUx54FMrf0AiWaKpuMalCjH/5
nipr97lmTWfBkD6fz//SlsXtpCPcnILOksYW56Q7IYBh5yEpL7Cyj64+GbE5
nUFhUoAy0NU/fjRSqTX1DNugCcZDlLtSwVNIDp6/A5DNKTsJaejMVC5eyOA2
JI3nIzXCXWU0vb5AvjHDJrd1/fb95Kphtrfh1Wrl7fVX2nyfzCAG9hqajL6Z
URvJm9Ix8MfvT/+7wwM3Vg/JY9tTscZlrlllbmg9S/fBqchXAXWrgquBDiBO
xYEW036VOeH2nCEICI5BEkjfAws2jDoDQD3bboINtlq+6vKZ7xJWwkgOx6jb
njuNLKpk6wrjLdk5waIH1icwr2GEmsXkJgz/v8K7gll3QQxdaaUPDSxGeT6K
QqEcgQQ2Osc89YUcWRhkb/ThEf18sDMtukDu+BFx4V9rwyUXgskP/gZZtc0W
RrwkZIJsa/okouUxfYLiKj36BEY6tFDhqK+tHTUW3+TUUwURNOABAq+1zQCS
LghFSgH6a2yhM/geQuZRVEpSA88TyuGURbAEASYDyAaKES/Lf1O68Akk4UoH
mmyhczDWHbgBaehQnstWzN+Lxk1Ixe9hXFqA7WqMwvqz81Zo0SYMPW0H08y1
FNe+QUC9pFuwfeZfJ3r8ADq6LX7L7CRhODb16SKDHfFpAls3UmpWqlb0TUnu
YrPQKa39pJ/knpzdw7lWZNWnpxQ3h+VHTJQAuWvr3qkqqZLlHE8z8fK46fiD
sS/ChGb8if8EieIj1flxun3JI0GOOEmAA1fQK5LyPKHralWHI0ZMrrZqOOIx
pVADLlEUq9piKpN7uchGpT1hOQ/7h7qT/YmhEMxdQHB8bBpEw8XX56fPKXIv
wSwh+SpPGIsoTV60HgfF/vpZsMrXXowlu2xOnIAKAmDmV8YWJRObp2ETbb4N
XswlmMty1dZJ8rtlhcju4SHHmeiPOChOA/bKPkk/q28A1XfryYw+jqLxPCB8
lw/QwB2STa8xd3Sjc1DsTJdYu+ZgdagnCa8OV85NscKW9D9zfPmzMtqvaziK
xHiMYAst75iMpma6gq7tnOoSLea4uQdLDhbL9j2jyzcoOfs13Gnt9oVRShPv
nXlu7dMAIFMe3MeuiljgAq4rYzk/vF1i8x6K0aRn6Kqkh/J2n7YHXyzjgLpb
C8tRNyU7RGQQl4038QSVL/aIN7x3u+EOQqbQxZzuBnuCXZoyn2YGC1VVqszP
t+MpwyNS+QF3xTCQTRrGyrpm7lHaYuLtFycXiXwumzsA9O+5+MKOcQEpe9hP
PPtc+OyrZGagit5C4OZ19EhlllKOIan4j2yfbsUct0PvibkFCFayQ6eWGV4V
9y4MXocGH4cw6n47XwVJaod5uO7tqewvl+EVrMxuzh4blwH5+p4i+Lpqa6gw
1jnYeO8+g4Qe/01Kp4ARyU5bZTH19GHR/8tV4twRpm35XgoX3IWLume0A3kb
DRLcVHdD/Ixb5/ua5/45uY66KMZ029YOhpsKieh0Wfur/luJgyi+C1VDc+oh
54YqkGDxq5vGVw3LMemBhZhmg0CSvktmSbNDHwwYrjFBJMWzPd4ujLSN5Jfa
Fr/e34QdWFm4IyV3fb6xj59Umi9hJ3bwyagTqtg+jfswoU1D+/VqXTaRcEjD
MKucVNzBUMf+i31kxk7Vc0l2XCpeHE5Os3zOsl2y95dzYDQto6nxSt69OQyH
pDCJmjdxTJsjes/xGgXNNwKh4lHQyTTa17CwLsUvivEWNqlz/F8aRMnOqiFg
1nYCDe77AGBOlk4TjqTwKXmbptaD3v0uW2Ep9Hm3nYmyj/HcT3dmENJk7z7Z
3fl7pioyRxEY+rsfhyv54B5v8czM0TYihsQgy4qQ2e4qH2as9VehdO9KQzfW
RBJKl+Zwm3YCC6rm5UkCs1GfBcKvQG2Uhi6x90UDQM2sJzsz5EFAHKzAUT9S
VpQAOkpNwpFLybMvxIHFWy7gwYIEdAfycNFcX4PpDB9tC7HJ/f2pJrnP9pzh
M6/MdDNNA/WlyaBP9/MxvihJ5NFDr1wjMriaD1ONFfkbtlfkjB18mGbJ217w
88dQsMw4OCJkzIe3kRbasALFGXb+4n0hZSuWPmGLz+7R+Tu0nB8WKViF1eis
z1Exh95lRdbbfCL5YHk3Idi2a2y5POOG1Z2smMQFAfVY0IZdFojL9cmRfBfO
ZcGnAVTC3Gx+Lg7jX6GO3Qxzffc07a6aLDjh0Uur/XE38QSh1T6iL1COiA9h
M++RTqEm0hZShAJEAwEE18GKRQdry3esk1MF9040flKnswNUSPdW0TSoRiTq
0EePQezU283mlczq8e1qs88Vl74s3ZU7UTXcGWlTcPSznJfuKbW+4c8XQwke
ICvIUXByjnzoxIcKErAX/akBdc/SQe9oYD9s7nly4VmPzUjsaB3zYYFGferK
8J2bgeSd9lPsKH30ShEWx5NfBY3hZteisR13RC3fJt1a6FKOPOqLbfNkNz2M
PkNMghq4Mhe7M7QPxoyuu4xgI8o6RGKn/uOFwV5Eh+XVHq9lsa1tHXpLK/DT
pFmgrP40jLLRcHYOqsH5AnB+z5TpYMzz8y13OwYFg/ddmwg+kKK+Z3fPx15a
XwX/u4+UK/0K+5f4rNPhby32ORdxnWhXARMCYpOpDJ/Oq9UKArRUm8MsK3VV
fFP4qsGun06Wo+dY5MiR/wOtW/svePmDv61lfA1yNJGI7SNXbqHVevb2AU/e
oUrd8jhor5MEELVZ86trcY6eWp3Zp9RfYZhoW1kpdL7SBbSoS3JGFKtk8bNP
iyCQHprNGXFO2RHbISxoNN85g0kqoU7yl/pwTXUFrBv9/3JzIwe+yITvUtGj
eNw8yqdGVOAzRYvDWUxQ67AU/bgFJbSLxtdUl4iXFsmpny1ClYGprerT32Qh
fh3oqUDhPpJF4GVaxdHXkwUn3R12aRj9XJvwn05CJubwkCKCBq4Fv86BBcLS
+75fn7lQj6fxnsNVA7RgndkTJJhpxKLm46+tD4AzwRGtAFgICyE8XTvPcXub
gcstu1T5R9kAs3o+Gu9Nm4/PH9oiTyIXFwHXfPBnyyybUVIQ/bCtcAHJb0kQ
KeD2P5AKlkmZaOh9B37RPb8wXN7RPSdKScwRYMpncQ6KTWjjWhQwPdVy1jYP
SbboXitAkF8x3sYJCR7qQ3yWzFhKWmhffzS0DOuPdCNMNACaaRdMpP1U/7UX
kWo8phkdGjU/5Nb/f0U4UaQEkynvWma1fg+HT1Sw1c6mn2Yc7FI1/7RwKwBn
PmDPfh7iur5noOXUE/vUTdeoDnQcI03TO27cturWZ5J6Q+f1rxTHfuSXK8f7
WlFZ52+QDeBvgaBzycITjeAw4tytaQYpATgCLS6EM5vlLmZ/y7rePXBPnfFc
kYDY7Pb3DHPUHtvYU+tC16p6PQSbshjmYoaVv9M4lGXT0QaOX8hJu3PXZiOJ
77GZFk4SptYRAkqodwH5FsrQboSldzoAoZwUqUaVI57FvuntRdd0ZqWmPwZa
JTHIrSUk9Po6d6vYzThxqQbmrfgObaVg1XeO8HszmEgAKt259oBIFlgd5XLb
SNcj7Q3ViVqYZdHrtQzJnjEh/nFuq0jHue4GrXVdG0by/h4yU2eJYALYp4qt
2YRG92bKjaPkiP4BFw2wEzIa+ddGbkAur45QsdC3YyIhd9YZH53xV36FPaAY
RjZ57MJ05umHMwM0Ap8Q3+TkfJGUL85xN/CN1UzLEleffS3HCiJbQ1gu3xcR
cIzOCExnIi1Mf7R8pZZoriIUOPwK7eQlivZyWLri8wvMY6ixYaVbzbMVwLZA
HRSovv/+tlTW0/Fz8OOCQjs8i9q9CeihCXG4BhFKcdTcK52lJsIZrwe4u0ri
mqwcETLnDHCtZooYlcAyNE9LdRp9ERuXgj3oVtJvcy2R4Rmr2QHOi5PTgk6k
LvFYttCtqqu0WUYcmThVpa/y2CSOyTpGq/UdJpv6tu+IogBPlXxOTvPH80kx
5cOQsuZI/rc6m+14/+txoEj/wcIL592cm/BTEZ+jVPZJApFKwP8LS7nQ2+bl
8GC3TiQcLhRM/zzfKrsuVNQHPL4clGnDcA++cKiWZw17gaZEyd0s64eIuJXO
SVTV8Q8tMPXrMiewwq3ih2i7aqbUYoIJZ4dHEH0jAnXfJLmWgUkvVUFcimx+
HvNcgYsmm2GuZs1R4G1oLi0bwbHMtuXYRhadal4gXctDVEttX1C0RvHngdJS
MF2OFs33NCBmmuQDvzdvP62Ll6SqcxpDro1JXE2C7pYQyM41Kusrx5Ve7no6
RBMU2Ca61iEjYMmeJ2dSUm+BYQr95vehxLNOC3Cr0UMwgqwmvsxyexoV1JvB
itQZmk7ZcI+2nOnwoTyd1kNc7s+cbaAQwCv2LcpXR89waFi6aTsj1C2nJID9
9TDaPqsskYHmQBptxuFgcVWIK6U0vwWTDteS6JJImUO4ao4F89lNv7c5Nhpr
1S/gTCbLDONHHBuBXcHZJm0Ctcyjo6S17GnV/zoZcPV+fYWvnedTqPmakU0r
/Oz5z5qi8h+d0DHG00cPaVMXPfu+iUwcQxswWp59FLmiOTj+NvHmyN4nXFF7
dc208WUc8Et7X1PrEj03N5FjrQLfLf/45L+axTmE+QipijcFdMOIQjGIhqXF
UHEkIhAaaiu83QeHF09JMtKnohHfrKpNJcCxCYyE7VAecn3P5fOIR3oOrqHs
Mp4LU+H/ZA1qeoX9pOgbmS/r5KzecFtzTEKTnfQqPckp4UwJEnOtV9oLiMAM
9GV8iEM1Gl4Q68RdOos94OXLcgdjD4fn5K2mHib1xLd2g+NoL0wCHvhCsGWI
+4QqooLUSdsNP9ngWSILfRFfo4eGvr7q858IhwweS1HUbMnTv+pYvirqp36h
DmjA5fVbbGU3wWlgTMKcQF9DYxDVT3gD1BpVRrYwpsMXin0JJZSC/C0WM0e5
NlfZVA6/KqX04f9O1+PP9ZhDOvaho7qZOfKh/TclQoGIVUTfdvQLWX9ATUdZ
FVsKs0XX1I+PTrq/tedWNeGTlPzExe1Jradt/fs7jAEWd0XJoxSzVb4j6l1n
Z2uCroWw0BZDZwY4mRU36GK7M1QTfgXToJ0kuE4PwKB2KaMniTSoZT/4xvDg
0HFoh/IMQeVeT9B1rX19bHLTA/HPI6PG2fO8mHPwsOfn7MN4Swwzw2HMGQOt
l/wIR78AhEiaItM5BEHvkc38jZ7+mywFEf86cHErNvPfr4NdwEK6Jz19iY8y
o+NsCcE38F6QojxWpQHLXXZutwVjdkSNGM+icIYFKiJGMujt0Wsylpdqgmmh
aJxeTOEDuw6mda/Mc9aqwI4/9FhOMWgwy9GEGfja1IEurmEYZty8mHx5WoxE
hFEMXOCGF7iufNgkwbNW5w7Oqv5piusNaFy1MbsfqICF0sgLPY24Wr47PHUR
CeYXNzubCKdB6yqWC919xtLGyZ+owWjVrTb7VSv+wCHInAj5pYIE7F2k5pdK
69J1Ua//9lobtD84uuCv5w8PJ/j9vDyKwCOkI2r+1cXDIr3JCb47XwJsOiUF
hkc6jOEPAGWFaGCl6TXa/EZLkbJ32dSRHao+nQC4s7/XvBWAiOLjckl3XihR
vYuoopBujh4Hl/DWobpmOqvwUry2Gsv80NL5QWAelj+TAkgbhGRyC8ii94Fe
u3KWgA1HCBKfVvDHaBHfYj+554GyVOkZ+j4Vp54nJZ3b/X4Xi31znNCstjEn
8WQMwg5U8R9zFaVd7Ne/+Nr1AJ6FkAmSxERxERSTw2rIQV/vGwgiSwctlZkQ
qBgUrCtpqizeE+6Y4cmYOcTdqThCKFlVCIfI5xyHHmdSINEJN9N21hgz3sor
7yJ0vsh/vHwpVVz265kCxy+BdK1hH0TevyRO3zpYvPz0bwKbRn5Ry19cajRF
LW81fnxbqMffDad2OJfp/EVqM42s9joQRhGkBiDGP63JLWGkWpMFiqySUY76
63Q3nafsP95SFuIY67RIavoMPCz22GYXXRIVu1K9sG+0rv3kJVnFzWgzpuEY
nvmk907LkHWflEemvbaU/BE3U1RKVuPKl/1sRz5JRi6taGwr0zmLSsLk/+Is
QLYpYDjDHpRb0xRc0GHy/4PzMZMMau0be4QGRuESi2J0Unp5By6p7vzYtk3z
f0+k8XXy6uA0LITX7sXUrbyG/tUxuiD+9DGlQeV6wV+RE3GIwq8MfRfMwbKo
YbNGlBUyeEWcgiW+EQfeob+OJFOguAURJAeFTVSHs4yfev+aVAx88qkvLFZG
7VEM54AjlX1UpT83T+cMXDJ5BYqry4p1FZys18NgomejzIFIlJ3F+/fvYPHv
XRpy50RTv6QGP0c6bbKpiVv+jOkmciIVygsBjnbjYZClDFJTtplkvt3kn+ms
x3FwFP1rRRXZkjrkjmws26NJbD0qm99JzBCiDFZlNx7CGJrifKI/Jy4ILQG5
Z5m2NWdE/mUa0l5m2ewHm3JS+09uq0P9CFoBLaPmQLjRWDs+bEBfWmwbXtci
FFJ83I/PIvDpH2gzOgqY6fizwkBwOScES/lKfgbqqLodxTN6T3vctmH6w4EB
1dQs/PzkbML2buG+EsCtHBghhW3j5GYDxgmOOAyV3obgSq0dNSuHUXK7bBug
/uUhV189afJalMKi7vMQUBAeEtjVk4EKhCr0neY5DSHF0BZtUeQBd9qSTscW
5R61Z5MN8YufxMolJQf9H48qTADHrs111HsIeLxZlwB5i856LwTnIUcGjf/n
43XPAkXkd6YYpTmVVxFMWpoi+LFXZr2dhtLWyFEYkRt3NeP6+BEsCAkCgi7W
ZT20Wb87du0k8CTXJeDVFgVqtCv3VGzpWUJXQJGrpF9SN9izDKkvAAtOAKR0
SEUTXu0lD2tMYbxvIa/gT7ZIwUKQ/3kh8r3mUsP6F0TrwTTrdQ/03pWkfZfd
ANFIx5Y+4wbNfFb2Yq9ukjEVWapr7/iiXYYiUf/zs+nH07WmBosdCZNghXBS
HTvbVihbJk/vFJ1vnEKm1Hot37Cyw3J28XWG3001WzY+R7JndqqJQbCVJUBG
TIwFiVfyzVluFnUW14sWkgl8v/7O9ANvgXiCSoNf4faKhesAb7zTVpEoF6QL
FpFWaepCpW45Hs8OYLTy6Z3pSn14nSHTAElOY2CnZ291/2z83d9IcinlAynC
HQ4mfvExQBp8B30rlLkYVrE+LI4dASwckWiLNk9Z0OniwPs3y6nlxMIzTLkK
7ryV9vos9/W4P3vn09A8cotwrJQz107pZMgFneP95aLGLPHlYiBsEqfk2V6f
alad3RMLTJmHwatqhuMeYjaznUIl7bxeIla57HvR8pOXCxnhpjsCmQ0YnHCL
Q58A4L15prAl70sE9vx0ibnL8O244MzZfkJ9UwnmwL9j3p1owhUPLVMAs3vv
Uc3tLqr8drLHg3e6hjf7VxBZslo0z9yjL7S59Qx0Wtm7BRJ/u1SPSou5eSPV
cCDetdLwgtWyApTx6v9Kj3NnowJ895RuCM/oI66CjF9t7WbcbHxA4n0KHjNB
gaQqqOkU8GR+Y/FlTEyovoH3RtxhzGknn3co6e5uEEFdcrA4o8vTEGStzyUY
PnHPiIHL5t4eiUqTnowM2DstBTAUA7giTQ688kN7PBpi3ADN7PP2uAHV43Rx
6G02NsJV+jvsWR7myF8bYVd5ol/abMYerCJ638kTNWbBcb+AXu9J/kNe4qBU
XVQEn0T+Jcl+EX/0qYA9CV9uWWGyhakHTdVMqlbfsGHIOqxxAq589e1hC0ns
n+02m4v5VnQTDPEge6TONsg5cTAdUy7a3ITpUlYgMqRScuZe6ZcloleiiXiW
OX8X9BDthPufeQqAijXRntXCXZV63otjiyFeQEvoTt5QAST+hGEtUS4buRlp
Adj4aBOboAalXmD2HznVUmST5tMRFdxFZVU1Bvs9S9LQNu9i/dc7gNlJc9wI
eq5PcuRGdEXnp+mk/oOOPRsHbIvW87h3+/HdBxdJDTf/YHhn5NKyFFIlnuT8
TaX0iHBaALFVkSSfBGFGF/7n28ezP8fVTRDoccdTk40z1oP1iRm9+qqH/zRP
2mP9IDzvBsCxIA3CIJe7AzJ7SoN2/XouhD2MwByxzue9rxb946/uVmLps03b
iAqYhjwKCWYSVKdXVDneb74bL0yJwtVPBfIHvhMZvVe5L/u+LAtgd1TTssyE
cm/G91iGM2846Pghw9ONzJRRxdKXjYLltl7WgtEKy4/AW+XJ13r67EGUvF/1
ce3V/G9Is+3Ja9RJL9h7wds2D3OZU4FIaogX/jIaFW8SqSpNwJOFKiBexY9g
YtPpB7cBdwWbyERu5seZpC0Gp67EWdbf/uBhwO5JFRBuZi8SaWb6iFbsBg2h
+oT7A7z2D+sqc1+XCARI0D+hWuQEgY+m/CnQRsdv9ZMjSJSBOjWspq+afy7n
GJS0Kb1e0yKlTdQgynFlYRjKjfM8jtLn8fnlIvf4VuKOlIUjOdLURGIVIiKO
/AGaa1DRl7JnqYvnYwZPbOAnM0Qsi5CeWExukdBcs2RNau/QsN6wLS0OqwCv
g6dUSceE1m9A5sC6vBlOa49AHfHnPe3MMPZqL4PTRfCInL1rlJhnvkoEGWPj
VVdS/zA1A56M6M/3Ze8IL+sVTUrQ30DqnxWuTc4s2TOoLCkRaqfzlBMFkGV5
KD8paHX/KW8WmgnXMhv7uUrYyOS1V+6rhfZGX83o8IdPYo4Bc57cQeZswh2s
+Ybe7T+MFOGnJmkt3vU7tUxyUhJlNhJwFlo4qEWIa4X0m7fUIBJQl/9x5f9Y
EfCZas3vHO2X6/XPaFkmP9PZFJ/2pFLavhSKzvdxF0AIw7p0t11RJ+RonpEP
be3NnkjwKT7APB8cI3AKvmlAI3Iz4q7cCOXsd7X8s7+6t9GinUtEreE80m91
K0oXKZ1iS0Hn6ziK1E1jtV1u4RKXY3nqS8HXr//LKL0eC3sAskUJmEfbf30w
aIJcwMQ9R9ftlOvaWQ2D/2YnjDbq2WWsxjzI7eCAMy4bI3k5xBrZlpkN9AFR
/MmCCONXuNaEhyB2Ttd2IU6frMF9AUTMhtrplO/zcb3gfYMTJMqpYWYNflJ5
8Zpb9CKqNoBVDMnv2aTTreNjWvGnewbBr8h8qLQ2j0CSkLCf+dSrUNLoMTYC
pGQYL9zVjTkFiteegxFBYjZz4S9cNVqnY0FkWcqW0V/feG6gM7mxIH9Akgea
IiFjCuz7MESnSIB+hasDy9gucHdaO4volubkR+7lx+yqTpyW5huRXZ0hdNJY
66FrCys/QOsC5KhoixvrX/InOBvH2LcykCc8Xq22gwDkKuOLkdST4nAkuS1N
P3/hDZzUpxTofdmZ4Lwo8n8bCAi9AA0NS/vpqWV0FUrlVsmnFhS+ZmtDpQRu
6p33LscxFrmFh+eqMrOeX8QpeXeL1vyAoSTg2O5UTCJp10fbCAs/ZpD/kSHH
Hr1mr05HpkN2nxaUPW0hMky6sLKw6Vlj30/WXB0cGlo05k2HhRiyerL9yzHy
oqy6urrrYPOxraaICnMYgAFWUi585WQitOCLHAInfnXxybz9SK0CYngKMlmF
EyJ8I/ioojk8fejE4HeUklL+JWmgGc0/iaHgbvejYgFyBYYheUMyKsk0znmu
uXyG9yDDT9pnf+yYGKy2oZ3E+CKfiv7Kj7J7RspqkqPL5YvUltCmNC9noi2g
YiyNUgr3TXxEtYCwfgw8fUM2gOj2AxqGIJ+zl0NKGxCdnujD/kH9fTbVCG5b
mhkbZE3REo/ByS8x1r354HZsO4SqzPcxRUWZ+mERDXC7mi33VE4v/4rZljKo
KijEkMpOFiHHt+dkqIAyq9Qx+wfGq8l8Rd4i7OLuDrn2K0niLFu+Ju9lZYGB
Yw6RXMWz/P/0Nz9B2GYMIkkdZ+4ZPl4qXEPE9qwB82Oe7rpmVrfaz1TrgVuo
zs+1R84VaTfbGwtqpOiUu1k/YDHztop0Ydoxj+lc8b4MdK2H2+H116z4KcTc
RvTOCdsVKWsD1mStSRPbZI/eYrCRJ/mhj9w7ar7y9ok9v/ewomqxN6EFgkXc
sp5C5LgVZibD1SE+5+L3mAqIKrBmr5T49DYlaOdKNY6h86MZUA16GHxZ1ZqT
R/rpCXWiJZnf38RZFrDYBd72kVUiOeSFEn4dT+QL0YzcOyPtsd+ULhPZtqBy
ITEIwXFQ42ehWKBuQcXs6VhZtCZthqnkQy9aU19jif2QYlMt+ceqDKkiDmA5
W/n4R5KN9JWq+WGi6oeb/q3SmlVwEuG8WxyJsZjxkdL3avVNRDYv4CrIk4ZH
5IJ7+CxBMEmNVPttC7eoSY3AOQT07tzHBz+80lB0suUNErkeZi6E8I0NdCB8
ywVAeeWE8ntcwfYpxq1c057rLe35X97EzsBSFi0Q9pzrPVfzVQi8lVRwBw9h
64jELXoSXJUDwyJSuxEZYRCEHbGL00tldBhWFQsutEGFdw/et+Np81dhwObo
/VJDAPv9HhppctFzO2AzdY/aRSH86IvUdvImQvQTPHvi0vEYfs88tuwgbYaa
yPN0zPMjVlwFd8iPZeRzlk7dZ8g8p3NNqvSiTdOmHDb++0h/h4xgDk/cbtJK
kPZqqmdffIGeOovfUMVYMXeOs/pWQGmZvpuYu7YpHNb2qgjTjBFknWX46KGF
SX00Pb+WeLdQZZHXoHAR92XvZs5x9rrFr8dyj1R552mZK50uzkpwmPaV83Fc
MgaZ+WvILefkAlSvvABEpZFLBB8H4q8Ixz997kIdzGAJnuFicBXLPqC2T6l3
qiJsixkFIR88l+ecm2QRvB7W9fBcIekLROFgsRH++DvZNPUTUINfOHnylZar
HqFbJmvRJPBwUPkHAkwsYalMvK6pUkWVbEK7bfpKfkgY3jQypwEGF9O5353n
fd+tZ75YSgvysD8yhgMZZ7ilhzHc5XI0CDq8dAOHTLUrPSu2Zus8lcwzTCwN
YioxtCwuzFfjBFHnuYslWrPc7UWm4KXNgSM8/T72cRjDXmL2ug2rUUQ9/aDz
pa3qNATTo6NtdxC78lpvQ1sZiq6y1z6vqgo8RNyj5rGwdqclvK3FrMMuUzfn
e29oWjqt1NRiZtRHpM8+AQsssXhb1KS8bJoBEN2LNVBDpR9sgWrHLdveALOn
YlIk3u+jTAKi1GONAwUlDskyVl300M2nuNdDULDbneS9JwwXs2YdJrJxbtwo
QJxLl4DnCe9it0WWXK2jDsUhMPp/Fj54h9pnjnYD2DdWgTH9vHfACJOveJnU
BwKktfanxZv0+8rpmiW3QDxvq5Npnxovbvo6+33oF+aVhvWa0XUmkhny35qa
KxDX4Qb417ALM25HIOn/vWWLApHdSovrOJ1hU8cXz7JFR0FdlpJcYnXogLlY
gH3Fm/3fKtNy7wVk45TWst3dPzzst2qCtJHrKtJ6W5ET5TETJkmlUvKt7vvG
1u8vYUKD3+D7020dCVJPsjMRq/MN3bAxQ+zwMKKJT/hJT8/WgBndat0wfIEC
sVyKDaNhPcHhHbNN1U/kOUGhZdR+B51ABNyy/gvxUg+7rfBvhO8eBXeTJuPP
jNMthun+0IUCgMHHi+Jl0ltEbgUi6uHAtLRiQLX21qS2yLnIz1dzwAq9wix+
JDLeWzhjBaVdnXIHXmLDcXr3wywvDbbAPmtpBx9qxidBi2BQ3zrb1R2IBcJi
QIAAoEVj3qaqAuVoTQDPvZdaL0p5k0VBUZeWJ8GlKi7Rd5/tR+1eo/MdQHzl
BCqWXhz+kfwmHAMX3j5bk+34gXElv65pAz9dnyurTTCbZp7ujW/j5xlIe6pn
2bQwVPLIhy1pWc3P3rwNckFAsIHHVHbOxNBqYvarMMC9X2zAoW22BGt6mH8Y
k2kF3q43h26SozTMqoG2VaN3KgCqj6YpqHMuZq5AYeo4V64lRe0dPlVbvqb1
UnT73o4CMdp9N34uvFlSlX9FfLZ9DbM2LYCjtydFPCQM+JfgiFbU2ikq6wEw
jL4ykl13mnPweThdK0xlR2+C+XiZwaPY1rYBdp3on1+Q5elIy+wobgNNRspQ
9Jj78tW2fswwXpAd3koLESuEKvcMTT1mx0iPIMFQd7EdOO/U+5LA4Ltm4nBQ
Tof6+m4/NoXFum4HN8M8pb7D9SVndNIfVlgJs8LpRDtCJKUe5WHyt/XgLc4q
kK97J97qV4VtsP8AVj0ajvU3dfgDAuLkxwrTmkkhwdOnBM8bMECpHbnnCGjB
sh84Vke5bV1pzo4B/iaxL0qDdWh6ryvPYhAuAv5/W/vRx2grwEsGDQY2Syhh
6PSdQnP9GFm/WhPEhBO2tCoy/6duUCNOTUhwOtjBNvdcfjMb2vBnJJpP6Waj
B1fnTJvekOjsqoBvAKJVI2FgRbgMXcKlXC6NGtcf6BnQIL/yKHuiKRvZAUI1
6ABb3X/i/JtSzRgk0QTN0G3VLYX6OBsfVmwLU70GYFKGFpfVdK4gQxC3yRQx
nM9d/KZ5oIrPh24lJlcFkJcAlcHiZ0sTGjLvxZf+nu4MmUg74mToE89UelEj
qEZa6yxMStLT3pvSW0WwFWbOnQ1R5pHS4M7gRp/3kQShzYP2QcjDtE/qc1UE
Hb6PL+JcvXf9+hUC0orIfy4NRTLaQrumlvQkNCZmwId0yIznPAupoww5KTuX
3RQtN7ZmgHI0SRoOlN3lwKuZUO6g4RgfhXoP3UYoMXDk2gBXEEsk1XTnpkbX
Lr0v7V+5CmnVhLk2T2+WsJOrOotYShYO54mfVu4z+krwf6OT7VLGgUsS/Oos
IKwobDUXXOYrmNDuGyWUsl5ZlUS5KxVQun73Ui8/kkwNuioDdhwiaA4Dpoww
MUQUeu3ZJWply9qPTerRD7fTgLNZZCJtGzLegI7vWHWS6GCSoGmo0CIh1R9n
h3/b7/WzDleKqbF5Eo6iexcscIQJNNm3JuVhpCirugGE/kUR9Qk3KyD4oPuU
Qa1poj2EHlFpKIwKaLXCc+5AbR6M66xFNbK4B1BEkasxhjidh8gB4ETMZ2PG
IsHaGrO2cFXT/4b9js9j7OLs1pAgq1A3pa25WQwMZ/heECykU6uT8wfp3RpM
raMY3/jEwa1EnzdoGkVJYVDLKoLTR4JLNxzmfz4CYlyj7nC2xwuxTDRMIJb6
SbBoVCwCQrj7s/lycN/Y5kT0mEzgDBoRvXDUadKuy+wt8op858nYjXFkw+I7
czCMosDflDSxdnhbDvYY9Fk6amYnYaRaQsCY+T+Xso6SID0U7YEusejsN4r7
5qUe4FJ9eF1bd28goUdKZyMKOWGZ6pQu9L1tc6d623EvW9AV1g7KzBXeA+5C
nXYZKgDu8V4yP2vSUiXKZe7vO4ud7uOD2TRgmQzkAbJjLtcCVn0+0kUqNKJY
PkX4UmnkN8c+cHeSLYyrHr22uf5DRsNQGvhEyflPpbgbHq7lwYH4eHQPs//t
JlfS7WbobKsLYmqX46l9FyMamLXXMHCku7OV3THrZObOl9KU8ekR+FFc6dfH
ir2bUyrhTPNTbLPGJAaVedHzz/OxpxRGU+V+SvubMoHKmV1iLNaaD5x8D3ND
4EGUDCIfynBEsV8/lM56RNb1K+vNocBOn1EIv0e43Dy1COAmratW0wOWCfpi
shv5kUe1se0iEW4yL96xuy5C0/ClBbUPqcKKAR74a+jcX94OUFo27wiLDU49
VQ//NpYjCVruRpTwpqcwBmieNtu33FYnAHKMKSWpMW6rYvfIchFADj6rTqV5
TBIPXjGomYcYZGY81CC5XtRtjF79DQHxVSfk8bF4RcIWCb1eA6G7dzDmmMcr
ofPyUSAlZeGyn9Fia4CxqwvjBPTy1pQUvG+aJgFInVWPC3YkFQkCoc2mtE+R
9TEZVGFrJWOAQlTnCSuFihTRKx3xvhv3QP2/D8SEYLnMFgkIwSRDuyNlhsgq
e2VcdwZYQP851iTSo1BW62DmPrYuJWAnt3hPzK0voIO14t4R/m+xHxqoYo/q
Iotp1/XIgqu9YRpV1uq7WXl9HJkAoNnGDjm/fmhFTQzvkGdyJzf/ghR6Dgiz
fupfi7mHp559fAkulbJlTdy+UxTL3qKJlmI8Oi6qZoFpCFmkHPFS1XOO3Pb4
c8cxijYP4i32eNezmjlQkJ4hOkZKWa9S8DqjEtqrrl5HES7JvVndPxc73zea
uJdH/6hKQpGl18OAEL3DxkM8PX96m+t3ZiLUHVzEPNLEeowKLsv2204LAGEA
LfyghjLT/z3B0SyJ82mIw06Snv52gbT1zljuaesT1b1f5Uj7t75JQLRRSD4Y
y9gPrCbngR0u5eps8VrzsjIqizHpnUMO9OMu7iOtjcEjBQODvBqR1jUnCfPp
I1MooWxRUTd+lSXskooSa+ZowGwlNilbTee6p1XjXJwQ9HFmuaed6HVlhcHC
aPYHG3/D1PyHoYEdVtwpRxXy9lwTdO0ShqvAkGkFv4ylkzCNYpU/NpGU0499
BWNkuLU7TDgchLwHN0UtFBnW/G6K/POEmdYRhLGVPLSjqIvc9sowtzARyKGb
nN8Gs0kjoWjgFqfbJW4byIDvtkVaCBjssrtRhD9SnX05IHLyPBC138BzQoJI
dQ9bdikUFmshHmqN5l3nLc6z0Af4Rq+J9sBdioJxyxgeDCf02HtqQAbk84HW
sudMDzeTzKZud0Uk8tHeatn5+tAoiQFe1MpVd6BVUoEKj0WfwdyiCwaFEOGI
BFVldSaRZi3WCU5qLL5W5vPRZXvSGx+fCOlp9mO9wU1Y6BkYFwj4Aw64+kCM
ZjEkRPBv/75lP3FGQ4jqosMXPkvNGbHZq2I5d7bzaxLj03DFs/V2QwzD24+v
De/ieUWyWXPpJ0Iafi5oX6ThScp/AGhzvj68GWq2HnYThyKi1cG37B0lzrzO
QBOM149iTBwbNQLpqWpd5qsA3ChdOI9axV4Z7Z+H+Ex1mhpYD0Y8K9BsfIPi
c0T0kNIgNeUjOV9Fb2Et1sD6BkeODM0lurNzCQhptlEF8nlWdcG2/FwAPMwr
RWFkq4MBgwC5kON0AHeqNbFVZxJ56toIftV30ePvZ4UulvX5x2FFYqoFX9di
RyGhkfi1Z+lU7NGBqHqPPswA4Wo9VEha1fQOkWl3f6qDpRPXEwROwd3+s61E
qL96/U17aEp4IO4JcRKndWEpsyiFHkmkx3wJBOCoF1+eph5RQto6fbpvImr9
P7mDNDH6c0lz5/nW8g1kB5wzSV55EfNcbXJxOejR7h79wd2ueCiwLBIkEuvy
HhfPbOVQYrIHYH+8A8IM90aTBQRbazqxSuMKxFZ/QrZxeEf+JKpz3lLK6T4O
WfO03Gu/0/nbN9C/IZuZBPEftsOGVvp0UVDYFgyhAvtX9xbleXfEVtgs+IO7
JeKoLM+xPG94oNk1xYbHLomHt3fs6TLvBtQ2fqmfIF3ZrI2mShpkoCLjDiGg
NvoJhls/jqqqmWSelOgtDym0jaPwMacQqTs2KzfZi+QjZbZt1owX6+olaSU3
02L/94VYQVwo954SUtPAl3/Y6CVeBi0YMdQWOlYjPc/NLXf5P5Gd7gXOD6B8
a8qYMM4l9nr+/TivHdWMFcCLNBAvJT1lgRDsQCSemLr/IDhpjSiRIkWrqBon
v0fXMa+1ZylFzvja2967a2ZHSf+hiwJfdioOd8ssOIrk4oN3/6xXE10ucq05
BpUZXQkIZbrOoSLySbsLQuc5GXrCmLFKBj1/YSNxeh2Q3AKKagnRw/DiVv8V
VC2e6VwC2DutfA5x7pZWbkVXJa/y0zmlRI4bthRD2aCKX4400jFyIUaCtZ/h
TDzo9Xzi2/rly4JotsZ93yJPn/u7JujkId9Q8ufVs4zmkeEW/FQUADCq1kMN
vKuH6EPoYX06tz1LV0ulOHFZO9nxyVZJlMps7xXNjVjbMemNtLsYgB/oDxaS
JFRIHvN5rN+psRVbXUdrA2Ns19u4sF1EfeRt6Ho0Ef5TJyO1uG08FdStD5Ch
5Lkqh4rKqvU4BilDjsfamDgVVzb8lSW1hmw5gfaHlUs7/RwmJP9+o28I0gKG
3hsP0Jvi6cHXH7Ib0zzND/vYViO1wqaNdONvZnz2Jx0kt2LGR02OW88zmJSd
wfCkUYmNunDiIi9PvCNzSld4IIZBzT9hkpxzHxwO0kpB+X0zMna8AtuyicuA
VWuzL5zGgkAw6faSlM+2y7zhZS4zSY2e2VZODcl3uI/zcD1C3207pNhuvMma
MSWavt6ogPOxbYBBXl9UebJwkdXSnAmm2wMOLi+yHXCzP1loJbEMezWNQZZH
fYI25wjzorv2BPl25f+Q+9cqGnggbHE7bfpoaADXRcDHeH3dcReJjrsCp9iN
baxRfAUkxSe2gRf6APRObT+UoPBwAajAmFC0AEzMFHHlfNS//6PesPv1Wciy
WSb/MiSqSB/Y3WdiohsjGb1ehK2Si+EReVeCDe5dQLBSkou0iCr5EA2X0Oql
gcJizuVx4QTXno60L7oV4zGTZmJJN7qaLq123GwdBHrrF3fhtgoYcJkNRgVn
oxcNgBHLdWgk9mcdYIAocyx66wHjYP08fYo2FIlatigj0XtQ5XYptpxY81VS
/5oX7kePaq8EtHq9F08xUNGkCXICAC4MWAkjNjfP6bA4gRndKYSLUPzEsvGp
nI7ID6zOvxe1kVW+bKzEgJ/i9ztxfSf+Jo+46h3Ks0HPiC+1UteccuqCfCSe
Nb7MqBXwGrAqPRcIEo5PFOLTJCMbayTD0MxD8PuDs4gr+eT+J6FPo4nmyTog
jou9focfLLxOTH9gRCiTBL6JZ/45sb3rfhyITEzLAzGzX8MZh6qS4GoUGeki
w1N/Xdta4TsDkMbMHKSjd9rSvK4fKj1/wjmTihPdXvdPYNzdz49XUrAbEuv9
2M58FyWUkt0ZSRQU6izdEHuFBfrduSW7d8uK37Vnz5UQyCKb1SQYrJD4J8kv
6FXCox1JPDkjVak67WvRIn+AhxZbSB5Jwj6WupuHZSDdLSXifspo10OyyeYt
/mYjY11MGhT94+vG44o4XbujlSCsk1+DY1j1iTg5LytOVr+tPmKgtUpExYJ5
x5/DB7gYYngRHXBXTlfkddRY9w/Kt/zDKKR7RQwTme5sQhhXH/3O8dXdP89k
/M9dcn2pZPgn9stkVnINrp+mkdb3HbMCZ8OcIsddNAcIaFbfvHC6sK6qtA2f
akkJiQ0yLVHpsDWkRrpi+4mKNIOUgWLeCbzUYW10nFmBXCAJFg7GJuB9UmUL
GuRKUMnZtRatpFKCuwg6xodGm/1qYlui277AVHsS6ThgwFfRKhuwgJQUJ5Pp
7dcDGIz+0FOwNAvpGFI1zDlg2sMvtXj9mVdW/d+CLQj8ds48p1S1N00WbKcl
Ua/eLpfvCekybfnnYiDQ0EVLO4IbOO1Gr/ghFSbY8egZAo6826K91Vtf8trZ
KMrx8LYYlHVM599HPvLsg8pg/c5K16u6/j/WqHGKA9q/qysbhsgL91QpDriQ
lW21H7DTsXsgn2mSbuON4B8w7DD+B6GgXiSekZmEn0BqLsJgCXOMkZxCSZy/
uBHTr43o9Cy2BaGjtOxA9oJmjBswQBk/K9JA9iI2wO1YB2lj1lCJB5h2Cc4c
F92f9xuFZKjHFSrDecQLAGP2GypAIHin1f63nlCwmMHVHxr8stVNkhdfFtRI
sD0AzhLqCUOFjKPs+EBGw+VOHUrEI5XXcLt218ygII/Y/Za2LFRiON44JgNF
78iKxmNIFDR1HMCbs8kvgW4RZ/P2bF/waHyngHu6DqEdGeAeglErpfSIUqLe
7QAeTFktf/Tx0AxmfOrT6cCesb2Pr/EojlsRIaa1x1FH9t9jtXdT12V2Qs9u
Hu7Mw9jjE3LKD/tW7fcifEcYob6wXUmel4NtN3gTQL6OpG9DXf9PIkLr5EW7
XMSmIPBZ/DvS19KE9rwapDsfCM17fEahTb7kWCCOS4ueRzvqYlW6wrenfz1y
C+LpJlEM6Hpitc4WSF7WfDZpFKXamdMdKrMboT+FnN3eOqadku5v8XTdxuIu
V88uxJLwSyh1To0hVI/Swpkna1JNv01hDRhiW9LnEhWVviZS+aCWiri+qZ5n
11ZuoW7PSWOKxFdsE5laBep3P0MmUzTZqQoBcEgvFZHi/CDZEvGA1bPcv4mT
uyj4eKplc3nN1baqL33dn/QcCjZySoMpAUTlkTzFiFviuN4x/bHD7UqVm8qN
J5LwFfgJJazAh9bXVvb87Xf3DUOryZWeRDhA4e3GtxFEU7JsExh4GIbsBFLT
+FhBDz5suKQ+EGyPHhrik0Lm3rspx2TyURYxhbzzH2CRZd61Yl9jbbXlyBQo
U/nv/Fgl2yp7k6xfZfvwnbmPv6lZvrQ3A3nNbxLT1hn+YpG1xuNIzO8LkTzz
GWnaEzzkkQWp/PDtDDOTaVV3OosJBmyb/oSMC5gzrinCv6yUQlqgAFUVf9dD
HFyJ9F9q0xIOHzq3FdbkZVWGnc+WRkRP26Pv7YJHPl7DPl+aHbRMv3CzAAXW
tkm40Q7bwlSNdPT04Y8K9exdPLOoPL6CnhBrVGl30HP3ulIsjztC0CIgvKWV
brqbuiBolLaQpjgkohuvRc9mKwWrcac444ihUMUS/kG+mXvj7cRPjhooAoWR
dVixWap/1tPhB/LRN5bz+FgBpH2DSSU1YfD+e3EC2YYRC/PChRrWLIwJLCEd
O3yI2hc2BoeiY2j033YWuPGaUTpTV7WM+SIt4FxzQAo2zhk/AnhvdXKy4M6Q
kPy7BtLA8qoIKg6tg+2UhFdOhqhwcuzTiMLjZRWYy6FNN4/UUhyJtyt8XQeP
XwShn/rlc3tNxapal3OlKT/Yo39Ab8Of6/aZPNlnSRaPPrTQvV+4adIW/r2P
rtRJ99ckXjNaxoU3/9t8EusnYQxpd9+yzZ42kH3GRrhMiS1jIaUI0a3xiNHA
awHaZbAaIzjyiF6gwh2GDrat5DoqAC+NUuq1PtLh11cOV02IXaAwQ+5vYaIj
3xYVhbqLbyQIyfO63F5GTkhymR+07WL2X8z9hoCY5wClvO2tBppT9efb8ZdQ
0UlH/+9HGEXkMixyEINAGbvGfXrTO/i5kRmww4GJcZrs4n69SCsAkqjT24nJ
SOd4VcLyZpvVcZzxqUP537vryquuLM8OgTaaAQB35gGEosqil2FAEb7QYMpA
UNXUms/jOrfhzkg0dwaSoVPd6W5TCVenwt49R6FB2SuW2OQNx+d08O3XX7og
chThhb5n93eVIjw3EvugKqGazkfRPgIQ4vUxnR7iUpW1OFIaAouduXm3vt1v
oPUo8n83DvaKWI2VVdhJI5SItMWAzfP0DD6UFxbSUdfV4vQMugpzjNvuEuCf
cdP65BH6dfKiwAgROwaBzpc8hUgGuN6decce5LHL7iMtdVqYcIcYHmu5J+HQ
W63Gnqq0xWgnQfXniG/+K5QybaL0nrwKC2J2KgCXEceMEB5sR0JAQ4onW/rt
HkzKhR6Bd0zFwcM0sbAVpIk1l+ChTzMogfqOmhEwCwkrJENrb9TAah7n1zC+
J3+0ft0kVv5eleSSJ5dSeo4AbWdDRZvTcxMt8na/wCu/HfUaY+b3iDZ7Mqk+
VUQ1GYlYhGhwj1h80uc6F9TEKTwTHQ0mHs7vjuEbNls+krAfcwXjnefZy0Rf
n3libV3MDC05eSSPOz+Os4jvAoEfwka9kLwqMnUb94tK9gfoDG3mBoWUch43
sxepheBq5WcY6jb3edT11jVQXcSfvDf0drJUmfoUOiHVgC5AxnJS3Pp3Amzp
0pCnOyl93qlPM3c8wibH7Vh9s6B9zF62kzfuHtAThAexKXoaZQY/ZSkDLKNy
qZerh+E5Y/zYB+Z8MgOhGn7zkRhrguQrxg/auozgEdRVzyPkRafM7tpQbJ2J
wywXLY14xJyL+7vbzqyNvfZisxhbayCPLoD8SoEAn/AYt3u8UdFrhOEyKCvF
4h40TKH0n8UtHUv/zoLcAUYvwSqZ8LDl5GpdDc+/z3RsklvlJYjspnd3Gk3a
KfMfvBd5HYNLjMr5I18g3bkfdWxZWZdpjJdWgaECVjE2Eae4I/XSKYe+KYAK
bY9k9k93fbVkMpOEk0Z97Wd/aTN5iUL7w7X9fLlQ9Sr/+FmUQ7ml2P4Ze4cZ
4VVGi+mWUmSQrLDMXsKH92r1yk48oES2Ji2KFNT6aYt3zR5yGJIP2ZZxCh+e
ydp2elmhtlBx7ONaK+d6BZMCL55IWZ2E6naISTn7oIeOXfOsa24VjJoNUjNU
fHSz/CDStiitBZcHEBqmFmdu2wme31QZ37xOAqSOpPhAw06/rKjA0FQMXiGe
ZN4/i0jMI7Y5MpELAkUEdaYvgPQC+VO4+ak1sAqFlD3+JCc46RI8vzKkGqrr
d2ACX00m4J50A74WDQdzw9y7dAESyzEjgP+22BAb8/oLW9l18FNpL2M35l33
oWHVWT6aEJft6Ro/QdgtVc/BXJXQPacTjGZ1YssZnLdbcbLaFmk8znWfJNqc
QHq2jrPDeDEMgW+IsDh3/56g/i8jUQe72POmonBMmFCgEcneaZms3tHNHJxg
edV7+IinWyAmOvA2z9N08ZcQabgqEBhfQGXS9wq5x6M8UQdVZ8jTSpwyUfBA
wgxXFlFINemOEOffJaAsG/0l7ErVdjCe0qEc7Qz1/2INNilNOAEOI2Ajt0hP
NyzkRCV1IfLTIlc/sLBzm+vMaWushdkUk5MW3cq//tmeiY1TvisFAFLn2lYx
/dXNsKz/Z6nrfSOsRnE0mMhDRA8HphUm3H+FpU8d5Z4vmzKI/NX8Yeb8VDUM
YrxFLllhQIILVIThlhf4ua99znV3qk1XaCLu4Wa0IB4VHgDbavA1fRonx+zb
m68bboN6uL4fZNp3qeCZqxLTNCXTiLg/5QLByAnrIx7/dsI5uqc34P1EC682
LtsKeLNP2oi/LwN+drzHL7WAqETLaF4BOFft/0jwGUCP8DKZcbZk3u1T6maq
pBU2xeAkOxsi9KXwV+e9JIrrXNuf4cDKRIcDUni3d1WI9erDSt8U9rY+Pdmg
ikASesQVFE9Gqi7/i6BbR7TfcKC92BeJqNTwnl+h2a/SFOqziTwh5yxArgLp
WBdkHPKZvgz1Oh8KYc8oGLrMAH4MqCe5NoyAMwbyuLUQNlQAm1TIuqSq4Yk/
50YQHxowyJJCj5h8cU9O4mqiqhvxJgIDFC7rRf7KFr9zE/b4nYgoVTR/HK9u
yXYeryMwhQ8nLQb/8qCPCAwiobApCpzCWBpvtW3FFCTJrNhEee0A4CVAYcpi
uJE1FYTH/YXM6X2qGiXObPyty5WR0saNbPEBsFDC2Y5yQ0hObalYnHCkj/lW
DVD+74M7TxRma6gc/6UBnWtSn63Ci7RJcMY/uj6Kw5R/1oU8MrEU0fjCHurL
hcNAeUO/+rg5r1TrY2kv737iZPdgfZ7j7L81ydyrg2x7vkQ0a0Nnwwg2eFXw
IsF4/eBfk1tMXQqRLgO6T9sDXRBSQKpFZ2wj7PexHPhwik6oZJtKVH/6wCFI
WLA3asiVD7uesxfKASgFqAuu301IR4Jfwh9Z8F2zFJrMy3ULbViDeBOSyOSo
Sfm8uhWRLM6LhQxLcD+ub6PjDzftB1TmFOD7SmxyHxqPlLsM+mMxztu0dYLY
fLuHYbNq3NLhk2sqIRkkTNi7KgdYMknBzkh2+Qt6dBptA3YGSyWTIdC3OkjH
zgg+Qykhcuskz+mNUkmmRaXe3C7A5+81BVq5UHyNoH60D/x+lsvNAewJBiew
7CRbrqNacxKhivdJrDggSi6r7PwZHud9v5czGXGttHcK+QZdiJZMqQDdTz+V
omJ01tFawj3UZEyPtF+//Kf4Us/ZGweGE9WVMw0Z5eu8190RcVdAYj9EplQV
t3+I/njrZQYNLc1Oc8AGyp2hcPQgckQ5MQcbhSUzGqip+/7ZMRHPExyG2ZRx
aHpDSMDt2+HkBZrSrr9CR053GLalDezDFDVv+lWepCxj5hbcZMKOoEqTwgrR
o3DDzrbM7Nbv6JaSqyPp3nyenu0mOVnWQzL0N5hexBfdyehlOY8jG1R9PTtw
74y4sRXWl6FxRQw9IG0t+wc+C/Wdwt3O0VK9lsFq5pxUpa2yq5TTS+f99hjF
G+8rVu56yjnye05bdOrzaGQXXGb8m2yNyqO54OYX+lqx6iudHiehtjG/Lfbb
ppBzTIwFFfO3d3S5XlRnAMfrqB0dHB4o7zu0FruAIPXwQrjDlqtpLwB5C3vQ
3ED5cn1sanYMvFEc1ZT6a5zFt0s0teaJnjTxsspDXRuk1gxzxAdWojrBeK+F
QX3nyftMD+uND0+gmDmd9L5Ur1+LbWZZimQw0ipgq+RxXRdI9CvK8n0ZNgZQ
sAqYlHNACwjXrry4qDD6Mxqpn1Rqan1V2qY3K3KTnF+APAiwm40IReM1xSGr
qKAY9aRC00YscoVq61Fbvyx3+pK/9q7p/oQJwKyQmHAPIznrE6QmZAR/G9AH
rkZkrlwCMccnJEkIzh0t6htCBIpDISucI/oXP/RNimBInLpPKT8Pe3RAcqxH
sxBFZgQgmaySLb6gT9xFkt8x7GPdyNBe1SIqWUKrjSj78F1Vva8smLTSkY6T
5EES0mrdGnLbO2c6QbWJrIHMMsua2J7B138IzbkscbpZ+JFipCcc1HGpfjlQ
QFBBjclRudsy4AmwC0uAAk9zQro1evkg2z3eKz/QiU0IA83l68p8DFX++siY
GeTil15hO5a6OQig50hgnQFsJxLbdmVHpBOONs6PoJaPQtWxl7LTzniZgayN
VVZwJCSLBNC3ZNIw6w7ic2ELYm09BJWQUAy8StFgQ0C0pbYy11zmeJG6V1TL
iV//v0q6x7yJEXLUeVJsBE9uv+ssY1GJkl7oF17pdvW8OCGzZu5LljJjyaUJ
2occPeguGZUJWygHwt8eKeCqAWnWhswlsGal7XqYGfA7jzkjrnQRaBDmVsbR
ASQCRIre3eAiPvQXBJTHAMmcPB3lcc2dU2rF3x8VIHUwLHHFsf4xpddPjOfg
8ftLroQ0HrU3/rkoUQVf/qKqPAfz9TAq/7YOoMQFuN2nzyKFh7TzNWPOWiR+
MVzjbw215HS0NZWKUUq+WwBjj6/QBQztqqZWGusiqhCj0IU7sqgrl6FZ5K36
F64uU4H7eU1KyY71VOUdJvUPbV50kP2PfoqcFacT5hvBCLaeLgasPBPil7Xr
D9fCeVgQtfKrZzRpGuBnt+yOE14Zc03qSTKkwOxsMz0Kxs4TwPWIR4erVkJK
4kwMETL8/TFzqgQKZr1PPTfDjvQM/3s5DeWeTzBvfQirOlHJBORrws0FxKEc
Y9ElBDswdK3mak77T+MrvaSWN9Qet4uW1mkQd3lqOSZiDMgnvD4jj5cQ4lSO
TZv7yOxl2gypbUhiSSpy6/qJtJdxSsmwDuLS+WESCViT72Zwt3MzG1nbScHn
6ombDMa9yOnScIgQjRdmVorA/B8GJeQxGrTvI8K+1XoM9fGTj1d8tXR2ZVb+
OvNjyTD9jQd35yYbqv3LzabM/Ee7cyRBlaqYVZw+qWKjaVXg0g+A7JR/rVqC
wfh8VHtohnj6PDDcUFZ/5MRFrVoCi2jQmwQnIXeLumbcdAN3TebfpkCSENRj
2iqoZes0xaY9jCo5H1V85rRbKLXf+HJbf4e3a2iRcHgbDXxloAZ8vZQkYYeC
obBC+i7phnYxErNvHQVODgKxKFNjntcj4b7YfP4DPf0VT76EXA5BaWepbGhu
fSjTi9czQiAMJzqOKAHiGTFW8I9RKnEnS/AeFAu64fVf9NOIooqPKSIEOLCS
qfRQ9yVbuRzCrMDfOil856ARWMrneWN6q0L3bJsgZ9nWWSD/Fg9kQswOqGj0
UtqFfew8co026m5qT0uB+WrSA5T/Mc2iVPIUa348cOw2sEM/nocLHBGXS5IW
8oTwLsoP0g89qtADyOBKawdnPPQ4Jw0f7rXA5r8fYCjypLVoEa9W5zNWv21h
KAF1BPAPMGJp+YYjCmE7IGu4Nm0u9LRdgv5VRjPL1cNsk2PIyqqD2GzmfVaw
1AYzJAcYt+1XKYH61nfSuJWVJf+J5eVqTimHHUKh8W7SDSf17p1FE1i4BBsX
XRe3KYHKr6xoZl1XUtEpwfW2odJI01KQ9gRo3JRPUCdbPEJqcBLHzOtNMoiH
IWuqbm8IsBeDMm7zU7PL2iDPfPLyJF4cD8x2E95UBA3rWtSS83ouD8scbawI
MQs8bRNRhZOzL16tgpvyiqaV0dGJzjWrtU/rgpA2mAzVnH8kA3BPny1ALFkN
1WiSE2j+CJ9De5nnGI/laVBiKYjYeiSAKhtrOivl+stnWOVCOy17hmXzxpfg
uzyNtihTqeFlTEcsGi1Xx3EbxgNP0hdNILkUxwNJMiV6yFdAYTt+yxoeqO/M
H8oH8ph/Ypo8jtCw9wPEPjdBCg8kDWvxdq966Lvkcfr6EM8SbAiNuByymXaU
VrbLKJIsG352pYfXsoOoUEdQgInwEmT56J8wwNNjQ8QlW5Lr5uOPb8ROf1bR
CR5w87UGs2MDPombhrkbar22lQoX+kDxNyfOh+725tHfxQAdrHIFNAmwFfzj
yHPRHE52bTfaB1/WZag01aWItxERHTUtmnsr/tb0+ELDljW5zVo05renvM5X
SxIwzmeEyNK3CGkGqQ5FdI4S9z97xQKMVgk/VRMGOj317nuD3V80YuipxDQ3
xf/DlsX/mRxQCFep/yLMEbDabEDLAcZgqh9EcjMuoaIfF4DSe5RM4vbvdntv
kRlSByL3TqG4DHPMCQ1RogqQfiDKgENQy6/oyKK0iwuunncz9B4hX6RwkZXK
z8KDNrgFXR4PspkXQ94wMGMt8Bt1Y6pQpQrG00GkamYb3zEJb3cHM/fW3bl4
wqwYu22zsqKWso7feQ6Oi2guiAaK8Y4nvAhyJby3LQYtj0aebhWdZoNDza+F
xRb0g+lTJWxQrUZAdwzPh7G1KJ1Ur7COd2OElLmBdBK3BSZ+Qbv3A0bR4mIq
ExwjAYz2MnEzCiRD9aaYeRApusyFsU8F32R+TGLAqfqkBwVtfQw1mJSYFoiV
L7eyDvzAPboCQdo5jJEEvS0SMww/T04KxK5e+IW3h5GD0ju/V81e4+oOZn3R
PX9aL3jK1FRF2C/AjVPhL89F1NFQaXrCC8fX5w0P7QRhVN2eFwOCkyut2IB1
31HLm1IeK03sSfX6wzw6q1h49Wsw18HvWbmMEtjRK2VFt65XYoF5Cngzdzp9
kT3Uh6lvYH7z+ATGiO+UAB/t6nKHB/ogbF33AarhE/qxntQduwLkordxoznN
ZGQRJcd5gDRPq8Hi/pAmp/esrmwdPIb3QQ2maAJO1hornF5KOH+C3/OIUUUB
zDwt9pr49Viifrf5Wof8tXlTxW4TI+QmFLOa/5M3lpP3Bx65o0qnqAhLuNTP
Q5xKhHasKMqKLqesL02Edm+usaYJERwAG7fwU0EhOKp+CYTJRKslqnQJfPA0
H7CReSx5s3gPlr2lz325I2CWV6I04eiyHvtuuZ0WusnHQS2iYTmP4KNfz/J7
FueFEOIIZPJjz6LyQf/9DoKlgjJG7X2CvPVsk/rc6ILgUL6McdPtKbD67PQ2
w2DRCIv17MgVJq7QNDAUlkeLkN60t3iRKpHqSBLc84FnU9orsRdGOvgWA2PO
JvhoJCBVkdPYB6rMpZCzhMC7uY4Rz5eaT5qVpFSGoO+t00hT4LM/4sdaCl7U
GxukKEQEv2NLEBVa4uVQ0EeHebs7AuxewWy3uQYs6SdobCINyi7MZ94m09NB
fUp+ef84O9zrn2tGKEWPomJXOfE1Phikb9jI9OQkCG7eWpDbUlJ/bORZJft8
ID7ohG9kNE+gC6lvwsuAM2f9tpm/Z4TBu7SXK4BV2rTIGA/DHn7KTPXHI7H5
oe6YDLJJJ/ybF5E/o0fQzJc7Wty6q+siQLL/mDFOTwF6HWw5zrTAZDDztQq5
j1/bs8NO+wU0F3gDANdPUqD3GK+xEoxiwtpq6x1P/fFgnu6j+ExAjcSsoMmm
4kCEWzSkwKUBUXemHIQGT9/JgMgCh6fGApIAsjR25fh0573IB47Czg4rv3v1
+ddkzV8mBuZbm9K7Otlov3Re5Z/wP21sT9ecw3EaN9443P3B2r7zaOi+s1Uo
svbLeHiVAw4Y6d3GtKmDBL11BsPJrsrY0mP8ZVDvZTdGnWzlRAAMtLUPX0Pd
WsV8dxBVF2kuB5CTGonKAoMeX6LaoyMH/M25VeXkgwkoDDOIeu79iE/IzNn2
GylcHmu5q2B8pZXxESehRTJonamxp0UmpvPkbDbH2qbDLE1oybMmrNayXElt
xrTTQiW7I9PqEuI8bvpAOxsHJFG2+bKfntfwR7t693DbnWGLa9p1WNe58jjM
akQDoQFhdD/ljHTbnFMxnh6YsTv1zwj/9ygxP+USxnVyOZ+2cgG/9T5sMc8b
MgzvDZjGwllWPhvq00rAlFRCzQ+nAKMsAmTCMkdOBeUvqGyWzDS2ZD2kkvGe
D09Jwd6b4xgJWgu7ThdFgEHu7wbnJJOqZdr86KzPzLheGTYiO2kDm7TAP9EI
o7V5X/op4QjJDf31shZpMSoWNbgDzFDjzE4OopUJjWGYuPyW1OcHYLyHHFuH
pcDhjMGC3hmkjf772a5+hUS84tp48dvqpQnQPn9bzMtp64GtyG9knRrrXipg
Whu/eLBs3womxgcZOlV+zesgA9LXlHMuW7G1aRk/xj8iSfs5XqNezQiYEqum
iqBiYq2w68ta2x4A1sJWsWTTEZguOFTGHNHw5ql0f9eXpBKKK1j1a1jkH4ur
sTeR7si+/hjpmgMlgQ8NfbYNrncTZq+navp3TRAcYkivgiCMWOl+APQ3poEu
9eTRzQ+RfK4gBC3Ak3Z4ylvMjn+Cq6OWyL7NwwHJx1M1Y0+vElNgsaAnRPr2
6PCTAZv6xqa0LBOvRQ9QblGVUd57XZg6uLinPrIXv1mxK/81OpSVssYzgJQc
8OfrsZigioD2gAt3Ve2m1Kvr9XqBPG80C/fmcAFmJqxvY+N5aSiWmFrxjUty
3hN4UYIFhdOowoH7pZ1miDXVPqB0SeK2ihfXwxdUbQeuU1GJHs8OwfZm5lfV
CBCYLfkrdvrraHDso4bRl5tjoMKwWloHlh0qk+kQoV2wdTe5wBexRrarM918
7opHwFTnQ5RRRoDES8+BvID1J54z04IS5GwodvOZhNk3NS8/jAFy0+owky0w
4tkX0wYkbzMwrWCfzhMCrDp6t1C2rIlnJ93GN1e5Ug0GCHq6AoKqjaI1tIGz
NhuQRyN/8hCGf4d1+XG7yXhCjStNUxlaHAqHL/78MjpVhFFgGVbppf16TsKY
2zkzu2MK3RAsXaxHdfoN/AWQ3O1DdlmEXLtoOezchoZvFsOot3MGe4Z+x4Bo
VsUvumhK9TGZE96zdio9RGqI9Xx5SD58KiCK6LxtLAFIasJOLtm4YiOxLglu
7lSrJPcGePzQbpr2Gc1HAnOakteLb65sIyJX/+64EysuFlDzNRZl6yIzmIP6
7NE5fhYLhmuSOJeGVghBiRRbjUExHhagHgIXMwao/bevOujDvRsWBm5sfftk
iX+wSO2C7sEt6TFf699ZaadCFTL7n3OrCjpqEjqE+gfpY0LFdw/kX8bkCbQx
vPoYPvgE5tfDB5eY5JAyMRnWgTdKnWg+fkgyHI8R+bKk9d4/7pi3poguUcjw
3DVd2CCMpFAAj4fvgS2sAIamWy1E6iSiugCt+o4g6ukgAO3V1yn/EzycgAsX
WKSBeeobunIqGhcYG2RfkwUeoAEFFOKMUwjpbM6vZF1tuGXKlRXhRSAjCQ62
ixjzYMfHx41om+dj2+FqkoDbWqkPSjkovsDrZk9CVC9eymDx32xhdS5w9MPE
Kj5qEZOasGqWRXKbcPKdqp4S6uzDuVn65knZFlTuEEWA/VWIDYy7/R24PDga
FREoScsPDxsfOcsqDzUVxR0JG7bovL3xqbGj9915BMzyPSyODP9G4kgKC7vM
7Ijv6lh2rn/7IbOCLegn//7LHFQV+5D7pKPU0qB5trMBpyWFU5SRGhDiUvX6
j18X06BP23BbmLtHPmsXhd1y1Jd+ahkJVKyXfGLnxIyd52kse2g3USJ+f4MM
9NnSoteGei5F4AyZowXqcFokQh5c9RXdmSxDODEiPG+z04Y/nsmw4h5QN9uA
BiMi8x0PIxTGDciDSr/KAl0GPdHgR4Yzxpgqv1rjLaYlnlJIYvzd+UUKDzBZ
9fuwRAvzWy0WFarxFxJ0T9z5ZI86+rNU+kk8qDQUe2uBZ9EQKhNTUAP6Dk01
GLTLCGLX3memcFG/ZZmNv1Mqo/S9HJQyo7yV3QC4M0u9YhRhVuCJ1FLXs8Pr
ACNHpYyVdKiuOmqFhhyieF30o3O/ZqlHZCX/XFBCgLA9EXdq+kV2mGpZLgqW
KhpZhl8O85O72NyELQF24wgOMcQIyjvII5JzMhRv/GwiIAO+PxoXbiU/fqtC
GMm0GiWq/AorEnE+TOFZ0mktOGrx+Dpz1N7F1cTO7Jro6jda3FMYfXFc9Nle
ahqVJnopRBokKPeLGC48+VjDQK3dNUCTJ7OkEMNvp71m9m0eizTN+2H7FwYl
JietYcdWdMXAo6iAWLSj1cdJ+lz3cPcryMYssVHqLT6CHucy2QSOyTqGjfkg
FV5evYVVAvfjI0LbvJef0KJDMlvg31hYxft+d6GCBziIuRM1f9RftkChtukh
LS08NLMPTFxg7LoLtrT4yx5TsadKaI0vH70TgPPoi9wVSsXP2Z2s2tTo/ktq
HcHVUohDmDq4sTo2jMOI1fnLxlgviDYEwpcUAhQxUEN8s3NmmUHCx9WrPy6M
fxGLSBaFXaJJFmYmfWag/MRYUatUpwFcTk1q7aOGtodz7plnYLlT05h/hZ+S
tXCQLRnMIt4nk5WuLJakXWcNqVLllB+dOyoNT0FRZu/o6gV6DYw4xE3IubtJ
pOQHHmvTvTQLGohrtinr6PC/Dj/qB03mD05ufCR7EYsZ4rD94nj3AQYMthR6
zP9Sils9XxFtvpKNCwGL/Obog8rGh1tPJX6AMRoNxyCTTAmyHB/GOa1CNxs+
LKufrnzrLVQRi/lHHVJYLD9/qtfnPfMSLokEfFiiEhsnfu7lkWqbRpOeUjt9
v97ILHFshro5HJHbP2E9UZ0Um4fYauFQGnNeuO+6JW614d61u+cgliAhiEI7
szBuXeuJbE87KAXTTz/JCQ8JUB7EsMG9lBoCT0Gl8Y8sG/MKRzn2BveOVLXr
ZiAjB9QMsh4xGnrZV9jhZCSL4VyjqcjfhwMqoQuwWDMiuwUu4//JEb6V5Ol0
hk2TLtEWfjs/ztwz6jAXFED4SY/xgSxOIS0GMfx0syoW/HdtsTECFrwu0xEH
b6MX6N6uaqtAgr1W7POBnPY66fvsT/6tQHPPE6amvuI9Q61WUuJB1IcGH8CH
niLx7TEcpChBLu36JlAsjjs0N85Y53oVtKxUYiO3mo0XEd6wK4aj/wlQZrAU
O+HwawMhKJVi6z0+bbZE6YHdWp5ClbXnOr98CVQSdvIDY8zSlt+0wBsTOV+2
Kz+WooOPKpcq1Cz5pcUr2jemGf62+/5fJNI+bsJDvrOLO2XctIIg16+d6iH2
0NRKJFe9GEzATm411fqKwXG+eTCC3gyPEDw1j7h4KZ41JFxKeHW4q/o2UvnH
H00djS0oVRhCOwiOAghsDxmy7iC8wGQ0Z/uxeSnw28LGHQlxq5/mHpdf/UeA
fawcb+fhRtmXr8dRmG4cUtfLkDPLX/Hsa1+bNJhxmCGjEYeISVlJsdXXuQiN
qPI0MaITxqoU5UFMi6w6P07lE0Cnd68pfs1HgXDmnTyeHzEwMB2k9TqvOZhU
oumKyibK80tB73NESm6pKskyQGcsWEdWHnohilqcP+DkylyKurJ+ysQq+EUL
qIabqNOMpUzhkTxckVCInrO6V2uIYkcy4HLKFCOUhyu025Zwa8n5Dd+vXzZC
SInz27IhY9to0LSTQ8dDuhZBYUvxiSz/QDjTEH35OCHFw944u1izl3ilEWrX
/+WHZCvHfOaM4W+6lhKG28RIEIaRFUkd4mE9E6YBeydOE7eCGrNoIFUeUzpO
L/vUBf7eo4pVkI2OYjLkvxyG5cDTekCnyxfmcldjgFrAfhaDPn/Q993l5KoT
m8WOSQ8Ut1k0wYxzNUzQl8jYtzIuv7r61NqIUxAOiNgJl2QXDFK0JtbWAM+B
ofPuar1bKvZBzF4O4pSBRxpnVq/vep4fm2+gc0LbF3J3dzdKF/2xhrrqFpZh
I+7pt7gvW2hZZNQ66dQlfZuiMQW631hpk88/77tjSx2RvtseC0AipqWWtGc/
fp+TT7AVOJi3WImeUJDZjYuHlPv+mKfB5I3jA31jlZJ+LxJx0zbLfVp0FKMS
PlfMvG3temX5ALlUagJxW6HSbHeQvjAFkcAtSGXSyGqq4GPPVMydxIEsyWnD
klQ5VklFE8nr+hRfkzjPuA/LN/XPGfYKeswY2ApJVo1AJNJBolDXKWF6+dGi
1wXzPi8jOuHyPF8iCrourSUC6jdWVA4gHNuxOgMCBJf8NgnGrx3hkQl1KBCD
6HuG66f9x72+5H4WKjYWDaDu7CpZW68NrMHz0kFYEzP2332/crlUWCDPeBPi
vl7E+if6B50ZhFt5dRDhm0ILvgn4JQn4Tl0MzTwbGv4GbT5t7pVBOENp+4Ya
UPS2IK02vLRvV8lwg7iTMAInGBWplL4tAF/SU/eyYeDN44kdUvhl8ICHN36Y
+ncxZxaEcQy0Qe9B4HUG30gL1v/pqrIUmUA6DERdFUhLleXagV4N0PqmseuP
s2noCpjLBXi9a+0iP4ac6bGeLxTUx6iTUJveJbyuQhuCqIzHeTdhgEyBDqFc
b/EGMDvzQhnaPuvCv/GLNMxBJoTL8PLfL1GCEqCGPkGjbHAEDe2PvKswNEZb
lfPO+S83zYvLuKl0OvEH3tsnwX782T3gFih+mPG8zVLtl9lVw/r1f/zDandg
dLnU1balWGwassgh/xhuNyY1A5E6m2R/NRbv4MMRvm9Qm5Se4IhLNyjB1uaI
kDXXsW6hsK9hccbEddM+VGya12CaOEBaDDzwd77ACsGr44IqwD0b6Vs4poXY
HsTYru3+P9bFbQ0Apzdl48W0/ldfSW5+X4UokB59UY9uZTX7wvDSRzhpzHlU
Cu9K13ogxg2EnwlJvY3onv1nuSHpl5heIx2RykcBXJxiprNqxzS1wCCW+GFc
VL+nl3wIPc+PvQfaof8oK/PEpHghV9N7ueZbIptEnGU9xVnH8bhZm/YW2nWG
ALCh1HtRyYwIGFu0cf/R1R5RbFV8G1w05zhZ+Vx/aGKrSMFIFgJ8iFSgFZuJ
+L/0dZJ5C2geVxBpdfhKeFN5q+WHKYnD/Xb7s+9mIhUyoSrqPr/VSc6UgSaF
wb423pL7SQPLXVMVGb3mp6+lCwKjoAkAYMpcJQGjOaQamIcUfa4VsNfbEa9D
x5lJT5rmbHKMFlJcWe11qcREMM6aqiYseqrB00fVJCAP4Ah82b2hl5o6sx8K
u+Pq8a+/hnKuEConTQZLEF208gLqGOqk57gP6i4mkiFI4LsYeWYm8Vddko7P
V+kDeJ2qn5WKuxe343qugOUx+gXhnFWBz5NCa2/lAp5Nl3tLRJBl0wLlbZ0Y
JyelYWpXFE3dStohBObj54J7AUtknj9U6FSAv1E+F+KukFZjPfTCaG99wnUe
Yfh/BJhWUVzNkT81dQ+/s1yKUx5AfxFaFXFLlLKOXdL1LhL+DAty4wL5/H43
b7NJfYR3+d3obBL+tIvyGlNXfVUg8R2fpLr39tgRIjQpBkFCIFxOCfnKHW0O
XT8eN225BMZLsrhMlot0QIIZ+uq6EMZC6c0MeFgPAD2W3m6WuNRKxSW+VMLi
szSVcVi14VUMIyHkD8hgBXHBm72s9BzlyY4LHbVVWvyNtezy26dgIeYNKtDn
nuNdr+PW2pMcDMxJMmE+VDXi9H8Kb+OMYQvhKNUK6Ayi71qjownTaxSCTbxP
TCU68CsWsdoUk1HNqDlVo77hCPVrDZr+mJej0O2oLuCODQpea6BaONyPjyzf
EloC7R0MZ8HfRxCS/8lutHSoua70uCoJqPCTkOKjtTtjeEGNXr7Mm4ylJSgK
G6CBHdo0KaKsm+Is1E+nU0gFKg4agxFb6sN5dyb2s/K/ZmVtIIjAXwKdm6Ai
DtMoZ0ugIQHIPIj1am5uqQ9Ds1lNqfNjwmJF1znoSOkMao9w7rMIh3LlRJQc
viOwp2At3zGCZIBluBCEHIfj36rSN3CGsXAOniPT0J+Dbt9dXRXN5q9hs+4K
ikgV/LvyoVXYEbfX7ZGZdQAT28iTwDULpAco6fjGlFhlcwGfnxrRQUE4oiWy
4V9evIzU1d9fEyATohzB7M6XoiQ2WrTf1If5iWtpGBz5vCqCjCLOUnlEN8Ht
OHlwU99q5NGkhLRy5VBUZ3BoBUQuSyMIT80dLaK8m2trPENIN10KGytws2BA
9AURPVJ+sw2deil9MJB9uJG46y9NSPpwuEHYQs6dkd5cC6nbJLcP4kLDQlxe
IegaDD5Ux46S2iJyJVZjYsmOybrUXMpVfjBjPw4ODF7IiyQGpnNOnx1yeyPT
ZpfzPUL1OVFhHfmyanryA8urf5LfLh5FoTceweyS4NtrOUjBAb8v044kXzk7
IdjXC1+qsm61u3dbqYHCWogW1deHMSLqScQ+OjtT/PqLEWw5izD2dtb+QO30
lYLWMfw5VO7cFgqcuOmViUtIUzAMVd+EUHCRo+WROJZuFZzZEJGwQ/VbSe7i
C5RzfOwSH6DH9wEFcC6hnhBWhDqtvTOvlfMbusK3ptHXIxwAwsrQTf+V9201
E3xC9nFmG/FknpfgLr8NiuGmTkClIkNtH1bFGhFI17eBxDFdVkMWJEtgBQ/p
gIhRG9NR8gHfCjTqVHmV/mmbPxz13/CzjLf3D0wProBn9SnWovtusiytZzOY
fmRc2xB/LDfYLTUhmYUdt4alyg9+LkAal6w9aCDm+rCipUTSQA0/faO4UP6y
Ez3BElc6yxZbBjxwqw9npiEuKE8QDGqVauXi6kAKWESlCsIbDzxPSaRO60EM
8sMwX4x33UOrDJqgGcrCRbeENrKPtwIe/w4UA7y0iLe54QhFyyJU5fLvYhKq
umv80mgd8A7pXC8yQuYzcGr5O1JqtZffDGC7Wobx680MO77UVT5eRacEcP5x
qsFRkboJadkjFdN85wpR5J95A+BvrgcZ+2R7jrbfMZj+h7vhTeDqVx5gChI/
TGpu+dEQAbX/ZHaK9kmsmjkyIdjoSyrbOEcoTvrwsk4LQQ4xBUGll0vRpGbi
tdRacc/MeQPp3w2CHQLGT4FvWbEi8AakBjL8qpGQFXUWqtHZ/22yD3kb7jv+
FCUBvHaWZTOBiBJ05i3lid4lCLOfceraJuWjUbAqFYbtGZx+KI5d1LvkwIlA
ROb1ohvjItf2440ZBz/O3d8s+iyWCKLfoEqEERaG9FUGLmruX6ACcyNgr8py
jnCICYwESoGOWct8Qrd3pIks0GOXPkF0x9tIfkCFrLcppEpdR7/afQbMhN8B
hzs1pU0EffpN7BJOdX0LY3KhQzBr2qQTLESaWCw5y26gU+iwyY+MGTUBrhPU
B+QHX2IfWbzWfJmaV6jspyUKOUSQQBzgF0Vy25yQWh7iaIhd9mfHMHpfUcpO
vHqDLLWsLTg6IQ+kGCE9d6EOJ7PUasn98vxzj9BPn89HhAifeX4kr7Ngokt0
2ohUFgge1wWMfxawxLM/W+TNrmHF2Q9trwt7cdTLrwFv8uq/6yMMIKqGESDP
k/05cJtbdUzWw/HAwJtdHtY7f/Z2ErEFIDpg15PxAajiGu3i6N9UTiOfYFpv
6SgvID+bcvBoem5Q7K4+Sy46TTjl/qjhhfbpRLONuzu3b52XKwLXCDLrFf85
UheLxLWGMwu9xlfxDDZWNA6uBV8pSwhjxv5NfYgYmoNZMWIEOw/Au+2hrRvH
TO+UOQVhnds//Bxl0BS0yxDqG+1mgqz3oZxlrmIK+bBj/+tKHB/omjaxW6fQ
zO7JefObsm4cZZ7RznYuoEwctHpsy3nOSCMRXF7TqmvyaIXOE7n4ENSOWoVi
WEJoYbEJeBWrMF+rnqGhOwp/+IrOQRObzn0ba7r/w9aPXZZMOUn8pA/rwex4
5wFgF71tAL0BlVkFJLSV2Bv7uU2DjRjA/ypWmx4DIijyA89hog0O4UJNlkCD
eVGHlj1BOonvD4HfS7wDqKlv9Twe8i1NCT5yNQ5BL8AJwmSzemHdfdDKOp9r
jb0A+nxpmlJdyYnuHTDJGb7bxo6iisu6NteswRoUurbN3S2xJSOtaQIzhoZf
tBYtbatIZpvddTxrPtavU2HPBUUfCcBN9v5+U94FGqUU6E4FxEPS3NZJ43gr
tN2XqJhbpUPX0LUb+k7fPhRxggBNyjL2YUc5oRyc/yzpGrpQH/0l8/E5q7TT
BPysg24xme7V0j/pnpPeKMH61fHcGE/G9PThM7ivh0VUrPIhUB9KrAd6zmHw
IApjLbOhvGub/KN9bPBdbPsEaVCQcjnraoFdbs+ido1qKp4jFgDT+uJIKVLe
Dh8GFu6qaumsbck84ubxgXds6k9DnkJkoIEB12pi+sYUp3qpTVCZbEXXHAwg
jHQpgKXWSrIra62GQaOzEARa/kNAnxefwZo11JxxDVmq5zhm/TrUUEfBOczG
+VoAnctCR9Y6S62nhdVf7k6GU7tMZk5Rx25P5mQEGGNYt61ilobXtzCsZfKj
/5hw5n9wrD+Y68AqhXFo2LehzrbAnikI6I51cJ7pk5KtUuxBBnWCldZH0aFG
scADST7IPFv76WIV3v4gHV+pZyQPba8/MZEcWYx8oDMsgQm5gvpusgMOjcdq
QjDSpcN9G72xwaHfVNTRCUD6DGFMUOxC3ddDC4JewIbI0tX3QJz/UirDdk/N
rQOlbGNxduSGbWp+uME6J4ez/itt7KTVO+/C1NvUE3NvzTFFrgr4uetqkyR7
ifeLabCC8Dlqm2uZMRfpuZ+1oROrK400Vhc3mFOAqKKYauV0jiKZkgczMmsr
CXM4xitBKUYz466yFfjsZpJ4iYGw3TWW0C8jxv7HyWH6rfI7iYXKtLOA56PS
Sy9oABkYjU7j9r/cmO+GRALBE9yYvegOEsRQOwpZcc5SGXnOYkA1ASP4wnZD
zREjHNV5FofgwgcLXT9LdZIOAXlZem2xiUoNsJA4Gtob187afjIgc53bdUfi
OQ4KyDdZs794kwYtQrYfRfJdPBLHmub/lE7pgl09qBx9vETc1xxKqng/5+TB
+sr7bGUoAQ9+bTrotsa9+WUZCitCgReu9u/1UMpEWFlsgmlB80sFhNkx7ffM
ob2zEYxaqQzw8/fk1+c3gB5Qa2KR+Y4RetWQSy3tWDWZpm31Kq2U6wPGN953
VUurYItwZfn1Mi3WL+p0ct3GirGYKA1SaRRmJHUFR7sHQ8XBIaQIGNdVnXoU
vCYP2714oxX4h6GPHrefC5p1Teie/yXl5uaZYBO6nFxiPsZyLAFotpvv/Wpd
9pUqDUIdZ6gmi1sdCg5hWkAej6r3c99xFgAmskRvtRXjXLMox4L79uic3kny
oAOMnVhFmo1N8Rhn6Ec7qqidA5sNEx9ZYEeVNDlNQ8MbCkbAk0P6q9BAkM9G
iEO637bvHvg8TQNlLLmDj9jzwu+Ian5MD3xVCLU2/rVE49kSukDq5OEwc/QU
ktRiQmtXpUR/5zQ7sEFJqt/SVx3qZNnn0NUZL24uqFIbnjGsDOTCUewn+qLo
hhix15xPlQ2+lSCSCVc4jp07UAPCw44z7IKUpd3MuzM/PnTAnZcl3pYgLYPE
86HDieGNu0WFVxezmW4fAndI3IG1H0k2Y78aWz4ICGatKqqrNk624SiYkNCZ
YsWrkthyLc3DnwLedp3/ieXMw8KbmYa+l+rX9DB6Swv3DywUdHVGjcXMIqfq
OSaGs7FekUZ74Cyknmy510g1H5b5cErOE+xiOcQ9jgsH23gXkGTQIrmVVbPk
kG8jjDOkd4DH41Vlx2XLVK6EuIjIzG7EpiETCnmzWBj+KosxGovaSMICCeuF
cTizf4wdyNUMfumWmRVrYpIW1kLqyh8MXtSQnNlU6PHute4QXD1UUie64b52
XHHbEEB57abh4T6rC0Tr4xo1XOWrEAdg7it28/ENBHWL42PhE9CCcmUQU0KF
td5fuDudpm1EwbChOULg9uw/p6SD1vCU0PDu5wDN8T9VV7jlEw0I8BrurHL5
OraXG1/P/v6BgcfLABIIkA4ukSJsRt+ilGHLG2M+J8TyBqB46jVtKSnsurL3
iFo0TXd0wfoRIf5L3rbga3UQpdyIZzL+chCAoba6CRfSlBhoKEMcOzgq0VY6
C09n2eFrzSd7969qebZCl+5yPFPmA0n/smYJL3pw5uNLWOEyUk5LpfAHJzjm
Mv0PNcGzgAH+LjnPyJIniEySY2tjnbHOFDOfgiLgUMpJTE8WMWoc8lGF/OzL
5YRK8Rq8VfFBuCaG98w5Qnv2m99nNx/zRRrlTeYZdLUpv4LJ0lyon9mjbJnS
tTqyWIg2nAPvvdxddpIhp7CVlpzE+XhXcbbdR8Fx2HY5FaqZskCDzN4yv7AG
9qRn+M/bAtVvvrcHj8pioUNMR8fy00JlM2niY16wJG+hwmPvuk1Dv/I4GlDT
oHnEv0C6jbz3axxObbbO+on+snYcHrT68kLmpU1EVJOyrjdh8w5z2V2zjrjC
HC68HmCQzE8v+Y2vrHzGQLYHfLbu1RXFqFihM+mU9QvilyvtZZ75jqnEE//y
bRba9CfJKbws2OfEzqxfZccZpHUltO4LCm+HE398nmsMNjy+MtpJsfLXuCZ3
C+V7IFvsAgFs96FLKqdiGMnv8p2ULkIAiVq1FNVPZ9M0vifnsQ0u3CTS5dXf
Ic39vpQOavod7Zg5jnUcw6IlsyyDx0ZfsG2TYUmYDAxyaj6wqasEorsSXq7w
GxutGNrVv+luEotnKpJu6hTGwaNCdQw2UJXOJD9R6wvU9SY+R2dfBWSSbCUv
tSn/lunzBF7StUrNvhL9Y8Gjm8SAXmhf0qUpCEyhWtYaT+aRJN5SzeXne567
Lyw3QHCHxuuex0mE7PP8hKIBQ4SUbPgPdWjUO02y77cqX2ZZCB19WcJUJnck
Vgf3sJjsGRrxDbAHMzk0EpGVVVSLKt2/e8YjndQQU5glOmamDnpix4zyBoRj
XicyNjnpEKM5kuwHT0dW+leGgG6SWN+AuSLC7Ip5Iec58Xs9iaQ8AGFUtunj
Zq9MI2OQqi3yrC5XnrFw00m0huOAw46Aiv65TOToqc6yJ3FDy4mioDS9ufrG
DTkwkBQxI15KA6JEOPgrQg8iMz4fUJEIA771yGcCEWYfvd3B3oi50UQLqUDo
X/PhQ3JuMC9/7/Aq7fOkmvSkcJsNw4qm4m/ycZrdOLQ6w3uJkM3KhYerGdps
g0Sjc6eqZ0kMlMQhwkHbc0u80vSopJmVWFV18o8CpHRJ9J17iYpG1M8H+hrG
mdH0ZtUvR041zBapr9VX7eb/zxNtxDRO0Zjedze7mOmP7uAVkiBxRI5jja0F
aR1TCc9AmpR2Lsm9bzqwXKsVxd9MAf46AWPOmDkPog+Zwdm0qkgLNv67Gfi3
hin7Xj78GWcPYSrWtMxJVvQzQKkkUh+T1kiw18ZxrV2PNG/DH11pbqp3Th53
MzvcuA+XJAaQWRSy901hDE1nvivjd5sq5cbv9aBXkTRF33Hs2MCRWjsdu+cc
28Fzdnc2kd4U/d2h12SIBOnNKPJxUX55pTBugfVATs9JykY6gF85PHl8yCSS
+d9WfeSZ5wR/cID5A4gDiv4rS0rH7y85zCBdlZtoDJwQIyWo4Gq9x24npsJJ
HZ/tIuS6QsqFHwUJOOnFI0tz4jG0Zr31nehUeCt2asbCRkjtXKypZMRBz13e
UEE1qGToGPJR4maeg4rioXCcdRrcxAj39jM2yj8cVH6AFwpC7XdE1+wtgZyK
p1iDdRi+VCL6Wp4Qqh1s75ofSwDeNo25cSyDQp10SwNg1K8jf2VM6Dj4fpAT
uxAsWxnbN6gKtAaIoMfiqDDhVws1N1ktWR9YKKZy2cV8gRZSeTUbx0aIRBXC
g4OnpkjVpOIzV4DA2ETNuLakIALbh3atD7jRh36pMepyMDrX0+wQNPfeo9Du
bV47QMjv6f3MiAEE9oKZdIJofkb9tKoCmaBcJNYKfX3GUpw7yPlAKNui6mGy
4oF2EUS+xhLP5hZTigLHHzgD9GiMXqLXqLRvam2hBb8ntLdBl5077zy5qknL
rL62EgWhMPPTcXr+yOUV8O/rnNtbtbMgCPY9dd6LNbt8+Fqr+vmJ0D2fCAzB
LaLaEmRPdosE08aWJ3nFOh9JSVK8nysatTFs7YpcW9Q4cCwjM+xREYkmySor
b+vkZ7ATPIG5v7uP2emLjEXwsYX/RCbnBd+85BLI3r9P+QTfMjluMQhovzrR
yHvHfg5BGzSQtA/4+AcwgXkmbeXySSo7fFZbO7EmlDbpFJyWotitJSbk9o72
jOGSwMkUUhz3Y7Mf1o/rVxBkUiE0LIi2TiTsWwGaXZ8jSx0AaGaBWTkUAqUV
FFf8e0QHtffkSAfsd8zcFSV5/tv8KKhuO6PiCldEYZEbNDqeSkk2OBpgKKI0
chtSJHpr5PtEIhSVKX9pLtZmEiMUcrDlF7EVxVN2BKEHyd6s+6CHPsyTSxzw
1xO05VGmarUcwzClrE5F/O9q6lypH5YLBnJxno9Ij4D4SCee1uOPLqxU2QQJ
g14lZl1Y4k/VNE9J3UnDvVRLsB2demK2OWO+d3r+l2yYRn97RCcemhAOKaBY
CsYZJokIz00Y4XWJ/37dLOagJdQ14XGnowIwdxsr64UBXOC9JBhDzJLxyh2G
aFb2fITLYM1Yjgihg1Lf4V+i/bwh0/HsUcTyCKJtOGKp5+R7DqTywpFZfqpB
rccvSd6XeYfQaVVIPrqQP0t1HA7jjE4xuq4Wq61YtqjQAewg7VJiRsJ4UnIV
K18vK4p9mBbQi2PGLoWXg6XiYuXtfjPLGKUULn+SoNwpK1kuQGMdyR/8DHnz
d6j4B3SZ9jQehCOvh85U5+ut2Lav1hrqsmmEErogHm61EWn0C8ky1OGbz1V8
6sWKfwiu3BtSqajcmhxwnlt3QfHwUVYCnF/PZyldADHnGiXrYVptb8MI83or
zFoP35hqLeweH0RcJNqIyr5eluARj4wEs99fLi6DUlt79+4Y4TCPqs21ohl2
P2/cdSFEdAA42rKxtsZ4sC3vpdTaN85cnBmF5pQUej5wmxJeHs+lVAzeKzvF
PCcapJa66Q1Mn7IzbnLz3/CExA75l7CrSz9/LERyjjjictfrWxTqn6Togqhm
PovXXDyyhbyuDiApYN0Xxu8/OdQH0390HQOn+D22/j1mfqMOufJI94NPmHpF
q+wq7r+T3V52BvsymQjrwzZPomtyhfZv3BiH9Jq97C259TL8MsfIHBAwPnL2
ufPluZ4buzhr9GgaEeM2tp4yKVf3byKky1Th3RqnoOzYGuCSBKpQXJhIfWXU
IYyFTrf9JAfUJ0JJKp8kMXAlN1bdgdgmKMjizoYDqgSOPZZ9DGlwgtKeBmW5
eR/lKh+UrbQPzrE+8S22MFebO0gm+pyu/cxDQ+9Y5p1EYjma6EoOU0hKvPZo
TgzLTdEDJbDhVLLaH0Sg9/w734lnrM3/mBaZ25lqPo54H2aKS19/d6otuBBB
wxG/Y3Hif65FasmIDhsBJTH0T5i83Y3aJOysV7AUMMtQk/0NnYIhn0+Vr3Ab
MQEtuOFTpf4avNpB+tND21iVJ+BkP5IdQDoECYyZhAkCLFp1FtaHQ6p/FKyi
cYVKQzgLGNc/TCZDFiR3BRLRYhoUg4l167Jaor62aE+DVQzscqP7mJPDCwmu
+9tFzjazgllGwsGXo8j1yfGkTmU8lhYz7C051EJe/gxnvpLRCfaBqwcPK+Hk
Np9gKDFbjv7Ej/w9V4VTPMnrK/Q8QkxOHmmA4gPvEz1AiKnrRnuwbgFLDILT
W6OpDZ0ut2fmO1hObljmvYMi6cA1Di9U/J7twD75qEVYRLudeopovOLdLIIu
PDlrYBVZF57BkycCzQJMjM88ustI0y0czwey/khMAGk8ysUvqKR+6G86CJ9G
Sl+hBONjBrCJjjQXfkjb34iqSF96E3fnF1VOIaeHWMVeTl9BHmTGr3+BVs0a
y6XyDMCOR5ZAEQPTZHA68aGacjD/o/hdqVXXbZTfuz686zIHC0e7ZRqLpmPg
M+rtj3rAvRoMIvQ+cBypJEsyFSP8i2075kxINQF9A8sS9efVcMhu7mD3nv9j
DgTvDlc6q+LiRu2NBTNzpoIfCjwtm2WiaWgb7QWnDmPYT3I4oZkfuBFZadt/
THyxvy+T4qHs3DbI2waWjPT1DwLl8Nu4yapfESg2q9xtvDkrc+Au8G4wDdp+
kkK0W/AwPHihAZsOAIIM408gqP8atfGoo+9KHLmKoEzISL/gRwWgTGEUcFqE
sIXL4koFNlH6pAiZHTot3yfrwGFjt52OY/ggrc9PSSMQ99IAVOkABUiRB8aH
kOhgLGmPA8lKKmO4CAoH2eutM+XQbwfdcnzdVMiWYYvAO0TAUxT2SYGktKD7
OeqX0HcQhl5SpQJEqQuaJZ7s1OJzwjwSJsFvIpobfunYUb52odNXU9Qu/ea/
DKvLA6jztZpOr7aKW+58nOe/wnEvzF4WaZmv5UmUMt/9cq2sAr8mEcyKLA/J
K3DgHpOx4eASh0V8ah3cwAKdUdvLcu0cpz+RaU6cYE6nkLozFsQIwNGWSsOa
VRC656oqcxUe+JGE9t7BOOAjFcMZGAze5LqaR80dY2+cz5LA7roTRtwSaAkf
OBTkCSmUCpfRQdPrR/oNJqRxJJwhbc2nKoYvfnJgUnAoAJPq6xt6MThCgfrk
dtSsuQS3s/98CtevLWP8nFR8FoERSPiZYLZ4vSns3ioe7dN9ZLQLdXog9PvY
ciMyHc+YvZSNgBJEcrPFcKNL4s9TErwhtJMXfUbaUavNEpAlHU1Ja8JfQ2DK
dZzsZs5XCBI6V49d9k9Tyzx27IJ3/Hcoh0hkC9tCE1oazFfZhh5XkeziAOUx
V1iMoRPVOudWSc/+SZm6TQnDC/vnqRBgeuoXGHWh4sjKyj1feVwDepavUb6d
28D4dpBAAKD9WnC85kTRgC70BuAiyLx2wERuknjLWgGyCBMU/eWGOTpO1tZq
g8i6JRBUuF32HaMuGnXbv1Zgm75qewwoXfSKuvzw1WcZlCsjtH2Km11l8pE2
gZlI/HVphQiy1AXRwpAYSKRInOZYoPYJdA95Qwh4S3yXo0PzPO6t/3BZ4Ykl
4mNsiaGlA7f7wSeLNSBgDdvq3UrycWLyCgASj3QoH1kQJzuIwDWK5mzLso1z
GYRlftRoAMMwM2nVCGaDOrE959sj/uzdGjkqTFDD92Tb05yUfYqYWAzvPoH1
d2/Mkm11tkTcUIwgavZZDKJaMgwwVqMBUA2s6jofKKqvA+WD3GgVsArrgv6V
YLBh/1arSbhZmbNiMjkitb60epAT9i/ZLe0SZNowLCIhS8FAwDPCj4HQvA7/
UY3BnBS8QjtjMj2XF3HZU8sCDGxd0kBhrTS+/JnQ4FP0w8pe2iY5quC/vt0F
xSJWG1kgHrR6vUfKkGxFN3jPM9GmX+QHtjMVc5sgYSXuIanhWF0AuzsjImy2
LrtUaiv3IAApbl1EHhfSTGot3edlLm/kUc9Kb9xBmfGfM+n6JwPSx7xxtW0S
d3gdvdeApV8nzxs+9Yq9mOTf1zA8+tz8qGvPXy48Yqf4SveKn+U1bNCBV8Jb
8H1KchH7wWcpIsEQFONBP6vCQRHyb8XApaML2t82vqEeuCl5cDk7j/UqThVP
s4Lql6fEQsGCmOFjNeNlDDIzTFc1cv9YKfYioyNC6iSu99F2n1xi5UK/uYN3
YUfK/mz5gNfBiFoDDCFLGnsUz3hwho7pH79pz4xj9EtrC5YGHsWx39dSQL+P
FiLebSQwORDNAuFHAWFs51OXyjzC44tT8a/M0+hIzgps8byR7mmu4V7T7yWx
ShvKVaWS0uKk+RF+aex4Kpb7wD+AHYk3jrQJlQ0kf9wbQ5RkUArk3VvcLmwZ
4yoBv8QbC2UT4YnD3Va8xyh5AeoZVwYl+sWdwjan3gvxqNI1eUn/oVJqVhSJ
y/C9u9dOjU8Ms7dIJYwUQ7NToWuQSzdwVUZYe7mRrTndaehC4G3uGZW+XmJb
IF6PInBLiKbsmjj7CSS2WiO0S9clbEDEtZ5NBvvyUQ7zwUnXfytzuDPLRfqK
A2uf4tO5ua/p8pncDFZcnrAeovi87RtwYMAynENfyZW/reGtxHprBYWZ0VaJ
XkhNATYkXp4pFoiLSflch6nnlu2LglPlQzcOPPaRVHBasO3aGJ6ZbipT5o3q
U1EB2aiuUVHOKu/2Xz0/Sh2AFwagyGewlVq6zO+bKjxrUJYfQV5GjSyKuJDy
C833Iw6VtM+AR3vmkyzcQOmQgveCZduEnb3XavsQDnycWQ4KC/fdDN703T6O
XwrDfA9PDWzeTJlbttooclyjz7bgPGF4HIzU3PvHxxlrGmzxPYDqfrhuRkFt
7mucINX76z8MLtLNTJspb+DIp8DhGSSwr7A2qGyRJ586ENUxQgpqW3Y3OssL
Wzz/YbGV8sXLoxV8XZAz23SL1Qde5twIC/XtjfHu2CUC2DfUJ1VHOcNMgBLO
7ykYIOPO6+Mu2Srr6vNhzvYtwXjNJmGckNIy/N80kGT93uVphz68bBSohQBC
YKQ9yDAIDE7d62Q9//C5NINdaBZnQBuyqG4ix/sCAVysSfZAUkOwfAED/sI6
CXeo/34OJgamjjz1ZSRB64FOAcMGcowFc0gebNdcuCgVPVpktJpglFuka5li
S/c11CW1kAFlouR1Y43guwNwl5dJbVVSR1ijNjCTJQ08ljuhmMO7SV4bi5Ne
PfUC7ekefalJJgretHPLkx//dnEOyXBkcxchaGljmFQWC/c/0n/bDrL854NN
1XVDUiwYhyaIZyRjr7f0c+8Z9GLRVZpsBYCuP83GC2QT0tCwmz6alubzAy9/
7V19IVR62vC2DtBs4Nj6w1EW1bIancJ3I02ApAj83pX/FAFRRZ07skl2zsIa
aeTtHEcKJVmXsOnVbTuZD8OUG2nF6zdYoWv7VAJTKN6YAVGIBKDnXxbRX0+3
gtjAViiockLeZRWPK4Jowr4bDFHDExjEdWOva9mpeUPEjXCndN3dL4GOAtjf
cL99L4tMQ6eCRpyhDIs4Q/ZucYG+MMFqHbrx+Qls7vBVA/pmwp+kjyoklEna
kf7Y1ecYcB8rnjcGYtnK0hI9AyPgKVIX3BieMYyBvcRMRnqdDT5t5qHMwWx2
wUJReEO0d0Yrywa9BeoVU99WquFsP4B3OT3ZEip/By8GjA+JaWxI50b6Kwcr
KFoHK0VlwycJPZ1SEm7z/hn0m5BiMcmkiC7VJ8sL7AV5yWPMeAuNYGndFbF3
UaPuELxBgLYPRHS7ZdIA2g6aCwSmYkcRwSh8zmL4hwD/afP3RW4TnJwt7hsc
8wnISFOeh567682Uk6hehQF/dcc+8BnN1yOWBC/Zipy6MTHGYLenO4ht/oxs
VPVuGkpSHP82kyQ0uQxRxGK1L4EMfNVOLtnK+y3vBzAEF3gVmaLjwQmpkJP/
cl4ve5LWEPPskeTG0dWMABXlI/W/85wCagtKNdM9Ajej8ZQ/VjqAt/XBjggP
JILxbrTaaUQDo6omTlNjK5RSX0aVUoPBFaF9piNK5FoAKJad1PsGadOfanGs
GJE4OTPg6VEV1F0ZOPnRrswidB57iKTQo4CXur+JynN65xRrTLs53jG3O4W8
zKoDPrXuCvvHO4Fe97+Q8Kji6N/a//z3H276epQmOdZTPeA7byafgJKpIhcw
b6f9yA+LQbgcFhi4zBjNkkgORLDES0e0fwVyr/RRB01q0VanQ7pkzfjOQCh9
X/cTUF1hvwK0DszmZ5d1yZ2Rqe1jippCEwMQT7R5giWBezVBwe42s3jFOR8E
7BI9J6+INmfqrT5frS54mGWxo6AFsXbxib6hOZ+WvOHTrQfTgXrtBDrWRDAB
8hi2FZwAtI4liHNUjdGtKIG3YGlM+2ojuy7i9gW2NcQ9/yiRkwbO51E9ORQU
p9i+hzgoKweAlwf9AQv7GIuzeOXWsfjseoRaVjskuiM4RD0eGErVTDz4T2Q1
YApRZh1a3HBlbMlK/NldLbjHSetkZ7cW73v4d3A6DtvyFF5LX45DdNPpiU3C
cQ1CkfC8nRRv/p0nYcd7THnItrqLHHiG+GslUpZ/waDNXpDK2ndsCQCHiugE
ftklUigJqR8+5xqqP0ATz9Id3ZJdKkeTDMMXKTUBd9Ajkf55rj3rRqB/h/iR
tM8XwYezcsZpWwAI8ZgL9RXf+f34JCLhQPsbpqRSgvXdrXRmvUttolITcuoR
XNCqfcOh8wJD1hXzamezbBoHtXKzEjU5O6Ga8z8MtEYZLtYK3puyR5JpBT8E
NIdG0vyvIIYlgIR8ggFHUs74vq5PWu29sBt4W27YWAG9WuleH6lYTrnxfQ91
Cp8YZkKjvchnC/sRAVXNs0BRftLnS0JjGOVIEuQ2WgFpzOji0QeK/Oj/flgh
4aywNVsy1AuhpgzMgWByS2XvzKKFembbXudsVw1PUOm3uJlT69tmt7yGAGF8
alalLDdOKOOiPFocsbSH3599SAzTK/Iq/vT8xFU2hSt1jTGQIG5a3aYSZvAH
1mrK/RoSf5cU+g8B6o3AAazJcqc8KjiUYxhKCzhM5c2V3yKZv6OQ6V42yT4x
JyzrE4hWQgJiddERIW1GtYGtnFQoIIZMcfC4jvyRx9UPcuB3i4B1Sxem6rDS
NVGVcQ8rY+u+1BG7FfH0MJRk/B4+IntfazGS9A0iGWXA+KwY6bwllwtXZfib
wgCClnMCf0X+Qs6K2rB7VL/FF7/epS1XCSIpcMwdldcEdziRYU7fbBNDMwU/
In1041QQmSdjhirW0NGMh53zPpszYVqyzOewCjQR2J7lIhw20wy3HZiOvHCn
y3DeXhYB2Z9H43/Uz0knMIGptiTM/IFatov16sgsVKOEhva6XgvSlXDw2uS+
enbpqo4bMCfHROeLLBIYTioYl3szu+wkro3JjOTLe+Kt4MRztK7qQZXPX4yy
HF301prMhCnGybCL6YiNt9fzSvFowi37m7j5GWG8ZLVXSTdw28Qk+V0wsNjG
7R2DLGYvMnXjLwNo7iFLFI/7iksBD3XXpReiyK/mIyHnOq3atmhvdS+NRcPh
1sW3mxfUZH6jTo67jZuDXLn4HoWRZNkB9ibQ85PeQRZEjMUrVonvZ42SCLL5
Q6muwzohQtNDM0HQRzQ1PNXiU9b++F1caBgVo7d1O8CbvHhRykgv2y5h5x2b
H1CRCXhUPDcBcmD11okbL82rirK9oOahAngGkp+K83QeAh3n6qOhwl+HfuE0
727jh9Qi/vyTmGH62aCE/MkJy5gFulXlHru+JYp0lsv8JwX4YUCTvF5vhTlL
XQ1/Pn+dVKIbHgQVFi+fb1QSQr6HH8S6nSKPfRE+9+UzjMEvsmreV3e17dkA
V4oVy5gPGmOXIv3mxycG1z5uwWoQYOmSV2pRWDRzCdPG5ugEoAiTcGLDJHxA
87SeWtE765b+8IZESG6YZ0pAH9Q3KCjD7lxOOQB8dl0NW0d+rLSnuqM59inA
ON4AiSC1Wv2ZOzbMvAtjnx/6MxzOKr+j4vz0gzv4K0HrwQoiPEkTHKdfsY86
6hHoqGgjqEFZQvm3PJQr7y9/3pXp7fQ6j+UfZTVEiLI4pD2KL47C0UUz2FYW
Uf+TOmI0lZmjxrA+aMQi9FPVpidD/Ryw10yQ0z7vihXAnpZWNSstDVmvG6gw
5hyv7sznEc9DycoYGrlMDweClSVVkr2WcPZ7hwhS5VK3sFVkTJMzAwaXvSR2
4lnWJ3LosE24chMf9rEbV4u3d2lOSVcueOO4NEMFxF6j7ZCz1PaA2QuIIQY5
0rziGEg5J/uetBUlfom+K1DjmPX0bEKCP9d7MhLL8LnwBSOTfktjcsMp0pbW
iL0pDQ9/WTEiASFL2uOIn8y/N0AK/YzyJFKXfuDQY+aWBPaqewFYxayj83Fe
2rapjekP0cafzabBXv40SXuVPH1xHr2mDWFSZzH9frT0j9fA7hdjKeEMymlj
KyEc5gmWXIXzEesFFV9rTsF7yt0T+HrMidtRl1ygAAsggNaM6YvDpoTqWEzt
PwdWkpXPoBzRMo3qxSCwD7772Z0fCs3ckxUBoGvPZ4chdxXq7OeM9CtH5FUk
O2R1hTYiVej+QhI0hh7yzgo4LJWTrVDmq8NtN6dg1M48AF65BXdRmSNP7PL1
l+FbWjvvx2t1RFvBHjbvRHZWQRAte4aZ8zgDvYbA457Jc8j+OCihMcDGR8PA
kPMD7OuWDjtflRh53+HQK7wzSZVuMK05wCS2ro5I8P4TGmVzy+wzOTdyX9+2
S/9WfvEvYzDtzfRs7PqG0mJysD6pQp+gDm02f8e2TAMiRr0RREt3YWpZybxW
f0BVNzlCW/SgRVel54yORLAeWugV5sXibanhC1tcHZSwaYWYSge9eWfZZMRw
HDCS46lt3NuZBZqgEdC41b9Mp7Vsg1oNRkhb30nbLqP0SA/smABGoKNsvhsu
K8j/C6h3b3VjYrdPQk7B5EmOjNzThvGwImG9/OCLBrVr3L1xCV//uJ8vGM3n
YRifk5k9UTM2jJvLGezgKpFz4gqgDAPm2T2i9aCMKPOeYX3X6AMSOeVkfgx3
Mh6Jcu8tYxWvoH9XzFGtrLf+k1uA7lhEsGvmIbxYlnh3aslcvgx//ekiG/LG
LjpxuML855U3TDIsP1SjrQnGJd0xdhf3qzk5y1NEgem0XNTif/D/5ZQ8DZBO
+/rGMzmp7sxyTcBHK906E5aPOWOnXQIjwO7nrG5/zh7Gob4pnpaaywgTBG0C
+8KxjTuiTr/zfIqo8HokH2HmPk76xph3S8lW+Ufd/cM1wrckDEKJDEjP1AfO
2fGMbTJ7vPqKyIpNIr9qL75pVhUIhfJvMa+ytia32qqzt8ljYD6keWud7/PF
RgR8H8Yd542k84RIsxpPTWmaEdMohQ9ojLHLjJWYAw/I1w10LxodmAWbq+CN
EAkKbPQ1jGvtATdpg3lXQcOeLWP0QT3FqWiYMyCGzcjfWjxuL9WrDo85Tela
keVNwNcLz0Fz2qws9oaxc/RsIl1+7my8m2w3yqbUgI5e5LX7TQBmSEoC7/mi
4i7aGErx5ehZUN222bUxlTYYi4Skv3UV98GSJEi5onG0bP4ODvuXbhs1ohHj
mbw7iSi3fRI7bWmPLFM4KCP4XH28FrpM93PS00w+2m5IKSH7eI0VOclGbivv
UvpUwV/+FwB/awVLrvEqI2rFXEFYHdQicy2J4nPLw17SZn7EQPuUrVA0kDOM
s+GmxuXvyFCJU0lWrlC5MxVcSBKw3x22670IXBjfn7vqzLXA3Mc5Ggqmt5OV
Ea+cXDwl0/rg5CWTydUZYiP4FdpFSxy8A3w1dhDtEFfoLPQZSTU6tNpOLkFN
SkqnAhSWRgwMrssZZ4LEbivOWH8uoQRugR/aDTG1yodLRxNRHsCIltWI77q4
xjP8ikaKlVCDV0QYcj1uNN1BjMJ8I+ac5aB1SSXBneAU1uu2tzY0kIYiDc/e
OLH/6BmzL3lDUXFUsCdc42iP0PsoWY8phdEWkGA6Aliwju9zGBwVt1P4kNF/
Obbq+UV5dglojXDJyq5RLtaI6QNvccnyLl4W9cTfrr/7iLOUrv355kEWyFqR
3oOR5cKgDeME9SzQqgrHCd+nftRV8+YKFGQiayOdDs55nYjk6R8KpFYNOnEU
p1oipa06YNBruIlPYIMVYnreFK+dgvIF9kCncxNvTxXk1Yinaf7oZuc3c5EI
+PsA/jarXIcgYI8WgdILEf/tFpCqsaqXIXcqZ0WZwcRjAADWqOPhI1zhZLF/
xA0hTjBbVEJS9XfeecfWD9GC5oU25tRLTQGX/9qynaE0VOBRvlkXuPaKWapl
hqBaxHppigW7FNDBAz/1htiaKwz80l4T2pzIb51kjmPR6AMeTt2KuGuhMrRH
2tBcw8xphH4vYH2xjVFn2FuO8/GLcM077anZ6Bn9mT5425by5DmwumqMgbRn
NFk2NBtAzBSh8KTBgPzRmH4vYlhRaZ2gcxst0d5Yhh9uGtQnPKo0fpQWEav2
RbVoBQZXhbWfkdBgNUM5g369JlRjeNELlgX2i2BM9CcLXMUDwVXb6S3dVNJ6
FE4RIn3k4VuB5mhNnIsexKhAUPxgRlfrjmfK0Wom5L4a/KvmUjzcEQb4QG6r
jmaEz2iaNxNnXxZ/kY0XsSS2LC2n2aAU+P6EEuxhPLTL44yEe9C6T4C0m7tX
QdYsTEe9jAbOhIuyIG7GL6nNqBulP1aL9SBIV4GP598Z8liTy2UWoH8VO9tw
Og1yahmaM4BgMFnX3MU7mf0+3KVCxlyvmxOjUyHmhGMa0mbxjGXCG/1NdK8k
ttKJqELK6cXTby2QnBSvXn4EZ1/eHzMyKNLxpRu9rrIftFRdYOJ3CDEhJMCO
gjbFPQAFs5ZZdEgAkK0Yqgu936GXpc1lPbOaLg/Ejt95CNwsl+PTs+OIbLqQ
/cCjn4bwTeR3P9ux8q2k17w6bt7mQrzKeDYPQQbIxw9G/X8PbJRBIp5hpsr/
zCW+bNAGkcURFkfayTomfiLsqP0q9QUWcVOKYh9RyZ0uC+vXBQzZZt9HJ83r
GkAMAsZvZcGXYQlc4xOx5D46YbzuY1sdCsTjXGtIRRekneFU3gGGzio4vxGl
BdhD95x5nTH4SIC+yJulTLAphrR6BSiLx0X8GwXHrvgjnxLGXRwuwRTQI/Fz
NCZ8F0mgSKUP8IK0Rku5Tkn2ldGLGsppfnaRJxsrNSbqEkl15J2TIcEWyLNJ
BF2kbKjyvZwTbMCp87UZr9N2pxT62Xel5yhpdwXiLPqI7Zs0Sjeam5zIZP0E
OdvGhewDvEKppN59+mHzpD9XEmL/ySHBjkgFFiRsn2sDal2lvSfkpheWpa+F
42Rrr67q7gNaU0kvieMjGEbEEghwMvbJeLdkvqaSmTLkpfizR026tnUygwJa
4ANsOI3uCrCPjMhJHxLpFpxFbanRgbwPx/vl4KJFwvCV5v3g/V02TQtFzoze
njUo2jIEh3j4SU7z/YkmThuyHRPis30siVZTk4ar1Oujmo0EpWrhI1MKZtbV
1C5sK5CF3G/3cOUJ4OWbdF/7zfZvbqdBHOGQDOCFDqQ5W1mdArPnyIO7WRSY
rr5Ai2CUWud1bM7mTW4ZwVk4Fa/dHqRClU+YBTOALqjVMRIl7CZ8PRwdQgb2
0IA8AFwhk48aCo9j6CQD26Zzmqjn1+tjFPd7TP1tza+QB8F/LJK+Gr5U+uHg
D4qt08TX7M4KEoR0pXD11MDWJa7Kxhm9sq49UOcVrUpfKNyW0RPmxfIiPTIF
lxctxI9KMhs4nXx/2wJXLay9BafvddcJQaGyHQvOF2dge9GgQU/2LTldj3MJ
P+5S2tWpthdA1AzGCtjCIQxvVvOxalpHxRVVpnc4eos3Sn6kV61HEt6ZT59v
t8tIPlSVkDkgVbp25DOuWBdP4c8cZej8q2pGAq5y72QuMjRAmSkE/00tigtq
6zei0RIysVgPjZkQbSKDAkxYPceZaiEIUp1CEBT3exHNwqEODt9+NlBEQPry
LoWc5h5ZhZQFkzY27mbURgs4EFzn56Gn8sG5zpTez9ph4q6KOrzznzTQzg2A
Qrke6JSV+wrQRxNYNcAroZQi/t1xsBnxMIHoM1+Ovh6KtNDoMIRDdyDUdSvV
OSvrKggo99NdJfL8wLhn9pOISXVtdEmneArwciDHXgwlYPzgVk8v1WuBkO2+
FdBKBImZbJKEdJvRGPoEDoITmeUGejuwjcZ/qGF7Z4Emy1FEmM+HO7rUhLij
49rG7NoldMl/ZOihbOb1wLee2QYeVvohbv7092iE7CY1PwFGR9DIy7yY6vdL
ESsBRI2aKXxkcQd6Z5DGhEUlR0JZZJf2ML0Jj0bC/DNGydWv11qCUUoy5yz/
SML0PNM5XAZwM2qGYOI3+lrAZx0IuLqwU4HbpMccCoYPibLim6oXTHe9qdd2
1FFOLKeIegx0aAwP0dgiVV+LZ08c1aRJOABhPe6HWGaYGvEuWZau+DhIrqzR
YOOK6uiaNtin1RGDKMO51ZHdMIoLJ8wFlAgHejutJCHD7Ti7owrTnHm2VVhI
3H4ASHpD4fJCCW816M1Rmnn4vcIczbdsoD47JM1iaxm0XgGvtw2bub0Z1S/l
Jy+6rL6WD9cmwoX9Nd2fu2YEz9TnNymJo/pRkFWqLv+u0e4VO9bUHTFPd3Vg
h2D49XxghY+WgED3LEk4KYbV/OXr4PVvUIfeij4PfW45FPq9vbYxt42MYlbF
kSJfGYjf2yVm+r+hZbAPVxuTG1LLOO7474yKZKQd4/KUU/2DnHm9xTW7RpV7
QOm6cxlQ9p8RhXo/N1KvdVUBaRE4WIQ1c8o7ongla06+UHG7cEqGUnRA26Pl
L3+canqol+Gmf3Dq/yHkBZXQ8fuX4K3obsrr0EwD93Cz24bIQ8Sq48iYqLP1
MEJcqAiMqBlPYBaUPtWle6spJp6W0yGlEcwmr6h0ZxflFhy/2nN5WzlbG/Te
ILYieozbDpQDhwfNXyGPDFkYygRChvcMNWuicd+7L8wpv3KvR/CMR7a4Zsq1
rivohILByIyye39Ph2x5zSeSj6hmaGw5TAX+4TpJALlfJqeKwje6dMo4kue7
jhAp6Fc4R/JsA9N6+FOUzO22h1zZzDZFNOtfDN6n++BiiSGugZROxU8+kuKn
9mzeenyHAbo6FUq8xtt+aPTmNejWnTpgcCLS95fOLR9YE1anNqErpGKJ+a2s
QsQdYEgiMLB11Y8pAPGqmg6RiTU9rk/8v3gPeFMJ2QFEPSih5jjayzDunz3t
doH2odNliNWGaHuiK7nMVGzXFD5Iu2cLHwhLscQmWkU1G58Cy9IJ7IaFxjqr
DeopM+gmL8rwmpyMg+F3dCVS76RvAWMo/SL688e9ame36moQZIP4uYw17ffS
UvAcdyNCbCqHhf2cheL0PAqkvjWlxdHcnjrbfuO8T+bldMe2L0NStj6hNGNw
gCHSnqriaLnToNVa51ydcVr6YKQEPYZs3PkCzrMygcH24SCMVt+JeX2EGu6C
OJHQZFdxdr1SPFoqk23t1VAQtGPZ9TomSMTPsfbjWKCREKvmuQskSPhnPIiv
iR0oxCUFaqEyoZXFB89AJ6KjxvEm++ZVd28luNuc4ziwGPyC9uwe/bL/0XvO
Dcq0fbuL4b7lTT5fRPmgTwdXjMkknicvkh2tJOcjUf256cMge9ADmKjmCplX
MWqBiajf/r+PEFXkbhpdT+xWkB2V/SQGKiEJR24MApxOXY5QqWfFRq5pgqGF
msCaumUihwYstKeVXE+2DcZgu+roR8OYrVX2jr5bsuhWUJUKXsibJNFtrEE9
o4AHzlrL5qJilPVKIxuE8ZhRiXcUnbPfbeHb7ebIaDd5kW0T46+vLnNZJgjR
hlIs0SBYDw9uFvMvBiqyvh3YDS58ts5m5JFFwQYzOdZi0ClpzNJcKDJqLb5W
L/yGPTOTBa2u2pTUOLSMK3/SuxLFzUqvH4Fz4G8xEwHBe9DQu7q1Vr9DSOH9
N+rB4YJyoc0x+XInlSbEhMvQk4S3AKHV/feuc17oFU4ECsjVDKiJLvzFRCM0
IOpNPo9Y+2EqiUYvaT0DGrQocMXC1OhKw6wnHfac8nzSmyxhR6O7N7Yrc1uW
bPLC1foO56vIFI2muy8bDCdY7QMk6xR/pBpidL2ekPoO2ocoN+XfF8yvACU4
wjja+zFqAlOITlf5C9wAcwwMdRfyC+ivfbDBrTyDeLEorHzmIy9bBBf1nwcn
NPLAvG5SsK/9atfRL+nktr6N3SDdRK8wzJIAdx1Xuk68gPh6TOe9Q2GPmQqB
fVqFghDKOLTPP0fDDvtziN4x89GLkvC79PJF71bpznzqZ27mzNeHiZgcTgQM
pi4Z2TMBMNz0hVsScIlFQPtJUoCqzGXvQhpbzGKPpQw0hYFXwtQiqVGgh/wu
q4PDVOGq0lRLeMXRbIJ3yJP/JA8dDqcaQWHd9K2dyfIoKy0BkS02sQyKU9WI
i7O6FAgK/8sL9ZkuwmVdS2fKDhgMaSn2fNFxvKAcseUMpHbQqMWJfTVinE/S
f85yLWYm8scNys+Pr/5WTf55J7EU7uxcD4GOI9Z1BDa7vsXtj9cSmEE0pBjF
5UshBqVgqVyEADJ4zf4N6tQQNbPFz3UVT08YzQSfmnhQWoA7nZ3ye4NcCbZ8
pSZ5UhApgx0DLMWAfWY2/MDgdyMKYNxSsAj2PdbYXYiI64pPgOT/scFX5muH
9SwyME4EsWXVs7mOlbCVnuOgKcHWEGibtgmsR4bazSBfmX3LA8BorFbPPMyY
4yzlpf69+UA1I5HAJPeYtypYIMZ64Yy6SQvwRICYPdx5stlB6CstpAHjE1HF
AFUd+XC1lhxxbDgsNeQkTTMo4F+xZxrzfn9YKiNdJCATbiVMvdTZSnognpBL
sSzB7u9L4ClK7GVL4EYnePBRi3qFJYE7c4JWfNG7axMXms5HYJ7XC+41urrw
/0CT198LFZ32JAjmNgrTXO9FC/Bv2tWC9SGDmi892cF8abe/+jTjspHAT+3N
Rmw+Uwccf+YnhLMpFvhhf0qIyaE4pskAfGs2ZoXXvSjhcrdnKBG2uszBBrCq
TxeuMQOyHrbB5OMkgsZUj2ukPtWjZDc79y1V8Dtr3HDYuX1f8YL/n/UERmTO
l/O5sMIyxPkga193t7QvrnE2CxLn2EjcTfztLUK71iXMt54Zs1e8xQvVLOlA
TpODAKk/HmRJDBZXPXRKa+hQHydqIpLriueuxBoSL2qg6If0vH0UunmqlCWR
YQ5U/YFvWGJkKKb+x6y1sEer1Lzq/2hcfNExOR4bKW70o2MsNmHlvlKFEtu5
Bntl+XF6m6ak9ny1mWyS02M86eeTu8ms3+78DHZ25JqtnnpWnYR//Dzwo29G
tnF8NuaqWSecuzORSafL2qkAFtFdYtdBqhZv/MxagWVW4I6ULR7Jw0x8JZ+a
TOd6epIcGuPhkz7JT6R9G4h0OvESYpUxbcald6H393cPvbX4h8c8aCtAm5dA
Em2XFFO0A7uMRwSSIOVDPBqrK89rh5huRhoHQYcY+qcNlfhkbJT/1Lv94I9I
2aEyU+H260ovQQ06+yqChHP55hemChM+ROGrb3HZKzl+k3pwv02iRmc8JMYn
mb84gUbD1pv7hGGmBNRANph/PkDspZ0u8jCQDrjhdKvS5Pcq1+PcuJtG3cMV
GM621JvCbiMtBYKD4msU/FwNZOTTZtVFAMrV4sX0jleRzPunBvzydG0mPCIV
lDNg3xj26oAySmb621eg9mYgy1dKxkJPcUlDpa3KMBMRs/NFPO2ketBQMKs4
QMoyaaAKuDUinMsXXKunpQn9X/fAL2CxeQllwvFXN2tV9q7YMb9DUDyEjwig
/QaquVO0cKy5o+nz1NppBVqLbOCuv2WhUOrQDGG9lWuAeBUYA6fPMiItXTXJ
XpT7bwcGJ5VMLfuUyr5peFSlWjwadRbUo7MSIdux1HWk3eW2d/zzXPFYGavj
mLWy6nWySTxVxq4lSD7QwEeQVRXEZNkv9TyI4ZbrP7kEyNpNSJ9oMuZw8Ly5
/NnSdpBWcTOyeSP2gA55iV6E+YRludtaWlRMSq55ba87lp6yYE2bII5Gt+zR
W7YFJgnb4HUFOC6IYK4nvLWV6lLpNy6Pt3MpXnj9Bcx2l00p8fXUbbu0qcmK
hDBUejPKyD5GW5itLRUEr9nWkvpjWYo/SocZ9TAPxmTfrx9VL0FvItS5NeAG
a9IhQDlMd4XXws8oQi8fWIfFcOdvADYq1t2t+ZQ7RgqBV+XbZfqiAJ8nEsDO
RGZ8dtlGww7eJYDcH9u+eirf2XC1ck78A59fKY8oyO53jnzHyGMuZOSFCYtp
Wy5eGr6VkCaxGCtEfSbzreAc0Qi5lwZxQ3NnNws3I0KMpEwCPRL9nh4guKTI
Q2ROX/pocvvd4N4nmzeAfpmq8gX9weCIFDisH1z/krs5wAt08wth6VReC3Ot
CX6bflEqDBVGoEYu7PxP+YSAQJ2ypdiOsfLjvB+aNelEkixd7HyWJFIGQXCA
izyByS0FRx0UxZXkdxUUTBfcMbx/KD/T6hwFBetGfzUy3w/h5vJdeAvdXsRy
9kYukwRs/eAEco0l2o5lSfApp8rnFsO/5bLMvcm+J/VhP3fctb0mezuxYSKL
YZJsQ8fhCJuyQZZZDZZORG7M+/Nj/lAO8uhkFqHUuCQomfXIGFBNJzBSvGZS
qA+AGMB75XHG0MJsse0e6BQBEcqD8RxZ7+44G/8tD4DHbMIeLfGZSN+3zQvo
7fJGONRjAmmuWFCIldIk/UadrjHes2iYR6Fb82OSrgAnkR5rnFef1yvNmXLw
N4jdJuUZnSx3vD0f8Bs9aIViCEM9CazQYG+OEvdR5MRp56dnSLLxvoNL+CAY
O3OaiE2P6SHO6NSvgPHRzr71WXdgWZS4qtgKGnLk0NaPy9K78hUanQf63B/x
xO2qO7Up0UFCOZ2XS/kU6DMvflU94aOtfYV2+GwpWroa8YtY+cSb0T7tktGP
zNhQx1UVpGnvPCvs2fUEAFyCzDKIghATRlR6VVaF8vQfSvYOpSW3ZogRRQ4A
rwsDuFB1c99aMhK0Rhnw7G0tASSYRIutZmuJy8vPtPhSpXfIhw26J2lBculw
4Sv+tCunc69tidfr8j++QVr6H6dV3SkqzO3NpQM2AoNl99NosinGvEqtHBLy
UvvcRoDuCHaWH6uGl74eMBVVJkODum9aisAZIQOEqmFTam81amckmvxaR+8R
dE9nm2hzHS21QRG6X4Uhsd4d6gAqbeN8poU1PF4zdPHH2bwrNL0dCCvkDI4X
xmSSRntiRixre+nwL+QdXJgeD/zVr5B8MfJ0hbMHM4yXA2Xb7YRqRpuRF9By
mScBQTVCO1x+5rfwV2NeLU5nsJd9ezU+zq4MDbgv8yZls/WQdx6v8vzYWJOJ
CmIDABV5ZOgLvjvwuCFKeZ8VoyTkeWM1gGkhEVDQ/iAKfbvl/WE3AejeC1jW
KnUs+ncXgiDZVJUK8s/nSMF9u6tZXivMyONRthg7YS+BMj2A1KRagaakWTCj
rxzt0ATPZJOB2lB8VeKav4OTwIYv5Tp1LhZ2c6VGT9qzbQdhsk/00LfDyMKQ
+aUR7LTfoATRh5Te87LvCOkX3MRj8IIC2PzERthP6SdKad/et4D1qttBv90V
OPJxEFKzOMUc53QWZaN/sbsnwDItUM21EfpTWis1ONSulE4wlEeN7h8DzoSH
lGit5+S/uoCPzVlt9iNnDMX/IHnZrAqiGrrFNdkwWtSB+0g++F/OVxA+ZvAc
3+7Pev/UiqF08vFEdg92pZFQSc/GbuNMAwf71hsvrVdob7o2xJM08qjvUsag
ZtDV11EZjAXVTvV8xNsPOQHe1PlK5XzAjUcXdIsO1G+8XrbuDUBNvQlbzRxU
6brCIsxTekntbIA2RLUvNXViyXLATGlTjJGrg2fEQR+sOtxIgK1t51MbVAPR
IdtSAanPJNy/8Yxxb4pDgfJ2Tnt3WtRoHlcTu7CB/7SODKJMO0H7MUFYbBlP
YTo3G2iKHmNFgan1hpXZe7bCZfMy9KnUvbYrTmjCsYl9Al59w5gihBqMXNZW
dzWyRBkEl+S7sd5RgUPylFnYyeUbyBg5AxPM9DWhMBrbTw4dUDjDwgj7Iy1P
IBdXePThkk24dxM/kONnLs8aEzYFZfZ9oVJDFSqje9cc6e50/iCTEmJykc8t
Xpe2eWEyZDY+1pXh4jC3Kz61/395lljvRhibk8sDKCkrhTiyRqZ6n/CN0S72
knV421wMQe8zS356AIBupLdyquTTdxbb/JY7C/8+5pe1Nso/XtjBI02bsdRr
thizlxamzH3HXjY8Lp96MJOUGFJ/Rr1HbXkeiG2UhE8qnvD9/6K6p1PQ9ZyL
tKwkg4FFchFJfkYe0PTrM5bUACeXP3xihpx6t/yphq4JEhZawIeHAIdrKkW7
qZihJcsaMDNUtfReo28+UZuF4m+MQobpbtZTGYj+d0rlConIOHYAebSqn/f4
DDgSMQNurzqIeyJYlqdj6VLJVF5g8KRJvpOh6iXx70FghBCUzROnzks5E9ZZ
6FFmP9lNds3MXI2PwfBlF/efVpwkEFLUJzhkboN0iBtlhiB5wQ4fvYiPIYky
bmYJblJEPfZ17rXtLTORSftaKiR4SN/FqhtDzG94VRFj0NvXo2VpqvadC3eT
mCXQy0TrIXzZGyxrvUhItdAcVBSczhuEAPSkZ8YxAb5Atjm0GA/Ys7MnYDMw
fULFgIfr98BlGYKOJvb03rdjLSSQTgQlPwqp3HZhYNK2jIv/Az3oNrvpj/9i
SsKqwShsx3tbG5TIn3I2zZjcXms13cNAoJa3EKHTcewUbBZuDlZJ3KouKEac
QV7n7PayT7+cxqvtPf4W1wIvHB6PMd0nDDAfkemp9iaHZchVtjLTNHFbn8OR
jWjaV+AJVE5Ifo5OUqlH71SNJbDvGH6oIvNzaCfiFOf3wYv+RivrXN4+KoTQ
Q0pLpjiPh+7smuXEANbkjRnHdbbP5RbrebmymT+CDRiRJkFhttdWUlK77gFJ
vzwYlMyggb7zW9D10Zo2sj79gJ8Yt9zv7AlCv/LU3Wjjc0JboDBcOtolLw1V
m1h7FkuRZqohL4YSXOeYjAZIme0nIu6eNXp+JY7l1WUnRFqCczRtl3uqe409
OecYp1weUR/GvPtEbIVdGkLFpHaY14eHU2AG2YUa2N+zA/f7HSINDMaLCab8
zkg1p3P/+MNdxmXc+r1BAf6WsizHGVEviB6gHZ3PwKCqWCG57ac0ecac6RO7
lywOSG4UroxOrGs3UnNFDr77+ehLdYE/V7OKohI9TfUhXb0NBcBYDvEGL8tL
jTF9nm4q1dzqGDM02z7C6HBKcTWGNmiwM9kUpNS3gumy8SWJqX6wJ1dZk1vz
hl+oYUaU/OvK4ZfJG6jLNuvRv4gXZvcV0wRzt4/JhCm/KahJ2IbE/6XT40E8
8fykeqkXZ5aqMKAUk6MIn4Oscf82XymfI2Vb6eL3J6yvOym6acmCSDg9LDt4
crKiP3BxA92dLK/c0x8WQPK39ETQYYOmKy4+sB2xm62g0oNTo7K7j1OnfNTH
REkm8XoLggn2Y8fHtbDdvKQ39OcgqMpKusm1jBkEF0Z3EM8c5+IxH0sAnAOe
Dfe90o7m4Ar+Mwd7Kz6dHZDTqDJoBQEVst0OPcRFvbDtQsFZkqE35V8XbQfZ
Wnw4EIYrJVjYnPrl7ubithx4z6EdrSOfrQMVRFMTVh9ChJxZASRsV4fnAk1H
yWzC1DVjwiAn4+M+LuSWhVTXSrqUr5ho6IjGjeWSwMGAtKae/0VnDfYFvL89
wX3CpiUXPdXiI5X6GITOLsaW8UgUs6JUouBy8lXx4rh4sRrDz3X9a60rrtJ+
Ep832NRvNmW6vbtMiRxbmYqpr1WZ/Uu9wndw7h6MSHKbi6jmAQBg1KBoCMl7
EqyT0eQy3vb9CImeXXDSLWwf2zwrL1EjyUJOrfiIqiVnzeHke6WzuSMclWoQ
Kdj13gTbvtndZV1L+WweCjrmVicGfozmSftBqT21Zg4vnVEGKNGbTrvq4bBi
GAISzEw23CSyhjDWRQQ4O79WTwSFMjfVat951UdjE8ZP5CEfc4KwgjBc5wgF
cJKm30mRZRyJa0zERMpSOioO5+7JUPpFQ/fNfskLWXOIr7u8s7vRlyhws/UH
BCC70DarhLcoem5lXT49cXp32GCPm6M9i9Je5gTa2KNJHDeVQKHjpCO5h2R2
K+ZKO3SPz7e/jkn5JFJgTpMLyx0MWsaAFd2y6trfHz5Xo7XRI+BMsOOWv7Ri
05qgW0KUjZ4Wqfxy/Zjky1KyBbNb6mdcvZpfsNDzvidPZFz0g82tb0zbPBR0
t78RrVUkIeIv2MmVE3x3QNIdiBis+fFneCbAvSMBC22swU3bSq3s/3tfVAua
eabPOBI3txWq4fLES3D+oXXVD79CilGw68Xd0ta8tR9w08KJhJntdDLSAW1u
YZHTyvNoW1IbZpTpffYPgBDFXKWB+zF6dpQBO6dMDp6UB3iqAWSScVzEGEzn
DaMx/FAPmCVXWRozNxfuth0GZU0nEG6FKThTAuOYJRfhS0qmNFnb7sMJ69we
XRgPN5gYv4ISOEgBwl+iJo0X2bheNVX8IIZPKH51OJUHbZKRiukDFcwzJx8s
cC7q5CSc9i9nsm3BFNiII0UMgK4ePCo4CmjkpA5hbTLiXyG5rsIwsH0s4yCo
eskQ86pAllgW/2gdzvVqZzOpvuAEjCqxcKwgdrz8PQ3GXings/exUgHEj2BD
0ecPcI2P1zDEQqkd+e44ZMH/bEaVJ5gzDqnOWIomoAEUieCC/DZ1RhY6T3H6
Z+mY4KdIi+8X4WGD7/XKDx8l0ti4rT9pDlDZ2VWZ7M3D7nRHcjmCQCnjVggM
yahT61F2vT1ZiGq2jP8OmzSq7sFccuC9gHiAlfpMe2pfFKdC/D563HxwjyxT
nbgVemNgcFucwgkLNPhI1u4/QgLyar2AdpUQwuhEGip3GqR9mENM05p0RNLg
fQK5bXUlfoYdd7nOwluKD/HT+LdH84jqDOk+SFxVS9ri1GlK5wyf2ux7ozB2
zcviHKDs7na1H/ExGLM9q9250q6bIyaaTuFc+bZml812xMylA1G4HNBsG0FU
xTZ9jvYTi8p0Ey8k1+Jvfl3D0YNz2jGiVcbn1KAaaktFwX9NwPqbKFYTa0RS
PjVlsitMene+VUvU/KI85I6DJzTGWsq8K2xGoxr5K5ZusdcxR4gHz4IeO+h8
28XLOR05FbmfzXxDg2OfMjpD3ur0UPxjmimyWSVW9j/gh+KVpS+K1XLCy/r0
j/+l03r4jsvQ4+5V+dkpjsAockozyT/p/KMdNP3wVZY/GIoYz9RyXmPezJ2y
mH4r+8hmcpuhycaFX10Xqj4pVarOo79Q2xQOA5pTouLAbw10cjJ4UMaVBwaG
Q0tJ2ZIryR2vycuaI7CTdNq9itslMuegDcop8/OIuvlRT6w/nJE0sKbwawOh
Pt2eCPohObPfQ5VZLOXyPBwKES54r+e+HzL055aUtspqnxW/xRyWCLyQOrBE
CcZ8+qdpcYIeAjJUIp2Jykqn7hSBG+N7tDrQuDtx80nhZ2kvcyCcLYfkni0A
/JMkX23QtE5djl5xS0lucUfMYIFPQsEuZorw+N2AzWFPQktePfV0iW1ayrXt
fqRvoqz0+S43LsvCzyiNshVKE/VZp1U5pp4V4WxTY4bY7zcWeJQhEdxmNwcv
Kzt6hJQFx4Xl/VZXl6OxcAPh+oxV0O5TJoPoYuDGIaIHgEhJPgjVcsF1QrBF
wzjcOhgRDYxKIUP1nvzTQBntCXjiDEam5iFA2qePHt+YVzi0zmv4073i/OlM
oEuJvC7KD3PzksxPyVVZPne1GmYrUX4LyM294NK3tfC3515oHjqq0nqBqzbD
G0UUmC0WYRX64mDNu3Apq2C9kRNFvDc4Q+cgLHMPsorj2kHCfxHLCiWIHcf5
A0zMX2IOoy6rsvRCpf3GTNY/NqbqJYQRdGB49gUUZBTgrEdsKq1R3gKgbYR3
H//J14E8Aya7g5T25BaVNV7cD/2v/4+quPD12szL2c1F+a+0vQxcHJVghZkv
CJTIok1wPhyNVSpch6nqYwBUXZZsW+rdwWQ6nysbL4mgbN6J95lUNVo84g7C
NFauJ2bf3XrgWCnrAcZqevumv3PCVuAEb93dCTN1W/LppPKJGKy55yszBaio
FgJ6Xup/rWhyeyCOxK57rnvLKyTwxq0SIeGBC3nOFGyGHxtS3+LEhSaN3qP/
EpqjhthA0byM1Qf8MsH+QnCmKBVcEOH21vBRQrhTcbYQt8YnvqO3D8Wh+oAY
pX6G/D3BotLRh0zZzI/vcNGp/fISEW37uYQiDP15cpRToGP8sCynraUarJt8
l0YSMkimWg57H+no3pbBmcl1re/NtAPHtmFijnC6AUmj/agUHIbGI/THcbe/
FF0eFC5zPTM7vbBIMKwFwZC14ontNaUdBnyx/SUMJyMhpDMnNMgn0LRWTbve
a4AwFhV3AD95lAajlVvSP/NG52FAp6jPO0bEXBiAVJlCQV15jTmpSKwWW85P
GC4rwYqWyoDxQokMAWz4AfuTInvYFOi4zToqH0+2yiIVgyY1bwG8u/PNXpDt
SSDVkwspiojcNcfOLSGD3drqZcqoXVogbgjdRs0ln+hfJWs+Ge6ybXMeIO8/
vyYIhpxTl6RhlV53FgiDB4lX4928jH4MHRme4jAxIZNwhlGc5cJesUlQf4Ux
GAyxrS/YXB31aXBWupi2WzUu7+hIrSLmHnYkLojvbSCAdlUYla3GfMIS1ryk
1w9VxVfevT0rSqv6AY+hvca+RTQPWZgnmLDV2JxNPAjzhD4E3TzOvVJnwh6v
poQ7Wz4YWjC+7aZESwHLEmIIi5ojuOewOiIqVvut9M8TiLQYCZqoB0VCceZR
8TZh/1vHP7/XMTcOplIm9Pmc/lEglAcnhuAoZDthJ192LsYET6htER9iyZnH
dQb/C8mBwDO94wrHB1ICutPln7XFtmFYDgcxZwm7kLsFjzsUXGgZBPPe1sZA
lqWfR3MB1BSiQP1fBuYufdAo4YTBlPgr0vxozAkGIYLaiNZRUwf5Xb/eHyDM
dWLl0hpL2AV7EuDPwMA/d8ag5gRozsNmC6Az4y2Zk9SOi/SBBybPMtXDK9hM
XW39nyEOoVqpS+xZkYw0vEH4atTjyRu5BdXVRtMekGjeqUEMroRSdZYPaV29
8L29ywKP1Gv6mnuLJqkqfaPfUuj3Xfivv0l6ghFZ9Hl1/hfS++TJPYXgGjXc
ieKSKaqbJzEiLtk6w1uT5L5pZtUg/KR+cb40iaWYqfhNSgF4Mf5ocXtXHXzs
+z+Phv+ZeFBpvpH8vBpbuPzFFUdrACtK0dtGDfBGUxeVo69DKhNU3grMcQbt
bIMPryeqdMvnz4n2/+J18xA+q7nHekTS6S2ic+JKKsHdUtzUHdZk5fHBT8rr
W6I6vLG+QWMp2zInFehDL/pgexeFsYtYudxxNg/8y+8kFDzcY2MxPQDhXJTZ
lfIAbeXadej5EJF1AfBINtFDuV3MpbB1AU0aRhuFJFnic24uQctMQxEWn23K
rYC5iqlpZUexEkW2SsG06vdNVqOXZi7CuSvOGtoifQyW9RpK1RxR1vqR4HW7
Larz1U44ldiTdq0z31mT0W7euaf2sZ/2Mz0IpSmfdU27YpECPmfyal11A8oh
r/9CFgVitHROx8MJmqGh/rU9eYQcxzEIOjarURpdqQBGkBBJbBf3G4KlO20n
k46lx4vDCM2DTouv94+Sap/KuJY48iQyYTrAYKcCCeyAUgGbjAm5nlaLpuBO
qxSAv0Qv7NK5boEJQKdm1kt33vcdhgP6jK7/6FxiOBnKHSJcCVkEMkhSetck
sYEXgXxddAZjHLPF3PMajzRc5lbQ+S/FMi5Q66E8RVunoUnWEBkOREjrjgen
x4cNUIKEL4FOIGFNizc78o9t0Juis6AsZqX8ZIh3bMsu+imAW3D7E7VGJxgg
ULRn0ZPx9C2pnKq1YxTQjz4eOnzQNfe+3WceoG4HY0ir7wi4z36k9Cdlneos
BYIFnrlemn82WBI+O4U49YrHmV1wmHQEo4N2CNo5DnNo6sOqdZbJJTeKch4p
gzH38800INWvB63Q8ZOPaOxFRsAHYrZ+g9Fi2A+/p86LhZ6AE3isOZnqGaXc
NlM1XA5zOSzXQm1ANWtfJcGghJxSC2C9m3bGRlqwuinrY49lU1rnCbGT79Dz
VlQKf14UGBlXbn76KFy2dOed8yuhNNKnui0pJFm6YSNGcZummrcXsv/FnLsE
0yxLXn1YAGu+dXGJ9dsdRh7sO6WgQIm3dC1Q0LPsLkCRrlvmuQhSYWBxagtA
KcAorpRbZf1E5hyZj0y26aNpvzIWOA7lz7m7QEfOGhXN2f8MtUrJR6uaItg0
nrQgvY24ezj4WKzW0Ftj1IfoOuz2kf4TYukXDkd1t+Lerl/SZZqvb6tG8VZm
UxG7LJeCPBISPzCCCOclW6AeVBljgt6TSLkrbKd2i7q+UeVB+yVIlnQy14nN
D+i0OaqWX4dO8foogreAPrf+x9juWuzgabRkfTHa8bipDMSFfKlN7bRTk42S
EMGp6HL8ufwCha15pW/boDvGNye0pBm1qeifGwhCBBgs8o0NsssZZAX4Q4fD
NPkIRzYX/I34XFk/IjEEiVpi4gbhYNGcbiYGGur707q0KnmX73XOCT5LOQ5y
IW9O8ql8yN0nXl2015Xv25Iba01UQXy3arMAI0eBDCsp97Ge9190RaLwQxYM
pWXGSsJV2pB4kuuLBQ9vAJW+71Y+1Tkl1uPsgWYA7iMtiuEldQ9I7Usxzlom
QTplqfvHF/2Cv6GWXu1lpdJ+p4HG2q0Kc2YUgBU6I6UNTMaijPJx++60CqtU
lXDJnGZMZWl28tVWdfk4bj6O0TrzF8ICZQWgv8WdsopvDYFif9lDAq7smrEh
GekvRcAJdXUOKQPUhLHg8ffvnRpbBJCT5vIO6M84CZc1ppjct8gtijpTysHn
LoLW+Q7paAtr/hAU00SlNx4aVvF/X4POH9IkJWGN8bLf0MsFSS4QZPUu78nz
axGNnDwQT91y6eOuRJELBViNbCPs8CrlOvV0nQQTQOojIn9IaYTPJewnwNkQ
gKN1nEN9+v5Zo1FY78P8Cv/6zMOX5bBlWt+M27nCeZbirC5bNdhu39N+bTBQ
L6ploYT+Wt1CEIhGOEXPKJX48iK56oMwwHF95na824uV/gSlurs5m4XGDWQk
CBurrW/ISTemSWMMxSpdjtUC3Nih2ZirjJp3e95hdflBA2azx2P6QASdnL/d
OQ08skf+NFs8d8FDmn7u9PBHty74Cwxsz0rDxiTenaGhXn9uNG6WbxE4EV1/
iUxV6DCw7fTGYVnb3D5xPWDnQGyG8WE1UxZtZab65JUjTL/AHq6Jg8CfxuFg
cFY9YV6aGXRDor4KIxZyA5jjO9tP8fZ2PsZ2gTJrqOIOgeXGz9Z1spQC4o4q
IsJ/ONVLjEVnJGkmjlNbcgMeodV/aH6AOmA5pX/BqdJWQ5zJraklRXyjyIU+
T5I69SIJsGswCQPSoZR+e6ZWQbqgMcOVi/ixEUAhkIqFZnz4xg21sSzYVXgq
oTI73emgSOFDF82XleQbhQSllyaHIxlnMQ362DHpulQ/r2KL4dzyTME2pTvv
6eodtERYmQvoXT9MBcO50ZY6i6XydsXkL+h+kH+w5RUmdTuurGWAqUaioPUb
P23dWnDcY90AKSR3bmqEEP0q2MlY7mv6BbApdParTBieEINkhp3W+DbZIJxl
AkwC0+aMA1dA7B/l4O2IRXDSv3lHLzm9GRutXh8O/K46p573RAnbYXIpcjkJ
VOYNiPIZKTIRTc+Hz3PIDvvdI3ZNeicDP3NCDBGOFum8yiL8WtmG1oysSM2H
ixFSXuJgSU9ltv1DQuozRvG2Wgrp7klEGSYh5tyfmut6l7nL8MQjO7a2jG5d
zBCVKgDKYElbVqXMpd7XJvWjAObZAYGdeZvHIaH4EfaxbYkHm7PSd/WDpcWZ
7XZD5sIngs0HZY1HB8VxLk2qNVwKN6bIcU341HCGXYqfEBDwY7XtVXQvJmkF
0gaZMldTVBSadPrv+VwryzM9z9yfRtPM6CAcyKHbd+zspGg0xFJmZxW6s0Rn
hPiD1azWZrBjLQ18Ib9ahutYIAj9FdqkVBzee9caR8doPzX54RJb9fMz+gwn
ac8ORajG6lcZ/szKtvya2GBGAF+XjhKGUQ75PRfpbt6wozC2ZZuWPtd9R0Qy
eNYxrjRlK2pBMV0AVSOA8j3xM/rKqnRuN+dQnY0FU/6yDTZyBFdUWUoddpEi
Vrm/vK2fxwi2sIEzw5GscIh8vbdcNkp6LT4c4gXBgYhgFMJqP+zZHHVBs4qC
ok1bIeS5caNw3RXO7foXGgbjZ3zD2giBnf8IiKe59IvCKKmrdPdtP8pyc7qc
1x3oWMSbi30f+Kl7Z+8Rjm+a5uT0vMDglT8JFZzYfvQS8g8cLfw2GDKZ/lYz
YLVuf4vCm29/j/vpgc2GZEahE9mrnkS5mqGpIhORzpYb1SANSi0FmDSNtEKm
TLmeefH450na1uD87BVvLl75LzTgau7Yo1Vn8y9jztJRIucyQldUTrz3dlI1
e6o11QHjefY45w1ToOIBg6BVi44hIKZTiT2AZtK7XXTh+0MTnobZUEqzz2gt
KwTXfZvjYMAp9B8phGBVE46Et3eYXDkE0kbrEk/YJ+6Zc/x+cMhtSt8frb/d
gPsmNxXWjVyOtmeXsc0IZ5MtKgiAuwG21o38iE7flTH+h4ewksa2QQyxl87d
FEU2reANkHWcQBGEq7UmBYh6/KeyHsPGu6sm5FNOTcO/m0UmFYs5UcmeZvaW
KV+IVLEmglxN8/1Zv92oJQfNEFQlO8jhXadLch9PxjoaIixSeJyLTW9utgNH
uo5ecVpWX0A+Lnr9zUkeLsJWlQlbenKRHkI5pYwJPts+ZwaMSc1WhE8PoINS
Gci1oB+Cdn5lXLGyXlb/y197OGQ4yX+m2uzNxdPcfLdg3HEOab0IyVLjDlny
nXfXnhVAAaxu3YUHehfJ8y5vCWKNwqyZBQDRqZ0qLrqenEeELWcp2iwmTB8n
SULtFTDt7325f3CJw+9Mj5rwIzSRd2mewiiftaQSP7xUV9hBdPOwuUaYFeCu
cvM6cQeA/bv1f89qjJlSEw0jlUJXnEFugl77Wi27GdyWRgMCkhpV+Kbhw5ff
UoHVsxBW2ci+lehDXrM04bN3fArea6YnWYrnk/SbOEDO9G44vqKebZ5deRiV
Rpd2Q9LaxL3+f/GFLGw4pf9SnrT9oQ5NGQ7z2in38uc/jMqd

`pragma protect end_protected
