// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
oVn/0As3kqiJfc3EjbdbGOEG4DGwuLx7NgcqoGkAL35g6AmbvIXTlBuOw454nSgr
yN4Y1LSCaEwtrpjGGvChBxbiZxBycRUpXRqX2IukC/LXJWwQKkp8KMHZkSRy6pa2
pytLZE7uY0Zan/d6k/nSnzStJmEmcUI2JwBWmBwBr3k=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 18752 )
`pragma protect data_block
a29vrisRSZtXYYktUzZuqotRK4CVwpLQHdMf/ang8DFHm3J33EFElUBL9//LcIR0
4giMx9SqNdlCRcn8ss8iJKH1+jYYFMWwXwzyCArtv2UR8hFGdDhWM3Wg3JRnfaGh
CeA88Fwpk+cRzEW6XxexJ+vKGL8arOHMT0xQq1/9hT8GFIgP1HqyPmvPpA8v7Jmd
zPNYWxlGkPbX1rphbSs+Urhpbl7TVjJ3Ds5+bVRtB7CDqkYNO76RyuG6UwO+yIiY
aEMWHJvqjPI6iVfjVzYB14jan9RHT0tF9FMEPlA6VFjBnPxgrfe1adz4+/ZdL4mm
l1ud7F7iT9fISxGVVgD+cCmNuk2a+7lUeurY7YsJBo7tdu7mh4WtAn+pPdqxSoit
gxwoe/6BgP2m4DHMPmlaepmR/9KfzGVv1fA3x4wbEovgadstSfvIF+VI+eZD0QT6
/Kexmhc1slb8vsx5Wmtl6vpUT4lno0/q8a7IMPyWiaZRT5NP8cFjbK+6cvoY7f4x
pGn5DGkIsChj1ahcG5A138EkZT7N6Xc+BjH+wmf3j1YT1UyXhftPE0HcMK7hrJx0
OgP8dghj5QSmNHjG7gUOlCrizvuoB0a6mdnZ7wblyChpJJutQtpp+LtZv5wU5KVr
cEecpW2ezhryIx6xI1JpCnSv+OtjsiwxZ3gEXEdgr7w5VZUqcvTc6WEbCxQZ9u82
vI7g6PFAJUFo+pPZusdRVsHTGRfPwhegtFFzIGNDpfakr8bBDez1fw8ad6H2STC7
ZAv8kX9JiGBWA8lKR1ZzlT+xDZfRoWArZ7kjpBWpAlu31bXRA4adR13skmow7X6Y
cqIm+cSxHPef3fwvCCLjQPv+WS4abhIE9kUYOfC8gaMWmWYfl9Zbkaa+UOdgfe6m
XycbvqJv2Xcad5af5OmhMHpMlw0uF03gIMHmHwNwwe3ltO8sp7w2BFYuyLouujIu
sHasFaKW9uDSzX/tVeLB4P5GminbjrvD7RjsXiqPwmLp5gJAaStp7sQWhRjqjlFK
AAeGeduNU3IAGhNP2eBWdHsoK/GRk4Zs9zQilV7Ul/Y57xC90+Sx6F+8ZRBtSRlM
NJdS6PA+JbGnSsdXHMLvWkFu0iLr+d8kIvqotS9jmFhy3avVHedDC72TVphYOG23
sFkg501pllempvo73jMZjHQgbROrgxt3OOD3LT9qFwciuuhAX4oEIX8HqfcbIJ9u
n2nTWTXgz3VTwWn3Z1gB5wSWZPq+WTvyo3Xz6L7jZIIsLSTQ3/RTK6RpdayDyRyJ
BWdMM+F5qiGF3t86lVxkPoyOlhjA8ccIG/LcQLdkm2yesS/v4GEbH15sPd9TfnIy
Ur9jUL/JkQX3+jbONhY+mGBVJa3qQGDMnQG8H6WDxCNBF0kVSJBXWCkiO2ib2eh3
/KO8rFHJeSiOLKa5GXFdMTH8Eg7zeiK0ujQkxd8/bjk+4ZaMNxvzbaFVIcCGFbRl
doy+YCbmzv+3OdG9M/LkW312Ls1YkQTl1R1N1qJOHkh4ly6KZ29J8X7ppoVfPCDQ
VbD2am960Tv1HxRHObIoIbGaEbYYy8BtJ0suuqQAlyr6zSj4fhXPjT6ADLN5gWQV
zlXsAazoNgciH68/lop8EKoPUcZ2SvtqVGkieXeeaXZ7r/Y9K0EddfGDthF08Wr7
bUgTNiXswHPN1JLPCJn1YESpqiGT+wd5ZlH3MPyTZ/6AWvQRqa0FKfyEsz1qh65T
yuvUR2jxryqGBj2r0cuvw4bKUh2IbegtKzRcP6NSLRH51I+8aJmG9nUSXMQc9lIj
+E2gnmHYeSaYf86LftWwhnh20/j0V9zzhhcaS2ym2YZFqW/29O236ArjtegOP+oY
LJx2dh4v4tnBA4He78WemCkDllxBNRuUT/CJlNCo9BIGangFizxQvFLTaolfSmuF
V4p0No+CUY7cyOOWQ6v6GvGVHOC983V6HKkjVuMznn3V0wxQ85iY8Xn/e8yZ/djw
V0SoqKTtnWWK8KMGNMyA/0kTQDuTv/135d5BNAHJ6iG6RtWJXQ2Zwf6SQUiUJOUb
pT1yZW6y9O4bDi3wc0VwYH9a8AlKuJ4Evl43DZp0eXZgLzBUgnOfA1ClzoWQ5TiW
/wgNgXVZKoP50aO+XwIZBKH5hw6s9vG6dZiWR4niKGha//UJA1mkmE7ZBPvWyGlN
JvR2kJq9eDVxTX+5VE5DosXDx0tOt8IQvtehBwpZVzR+DI+t+mrQwPx/NHBcYfSl
uj8gckRGjTnYClh7HpY298CjU6eYYIBl3y0eJUPQzkMF2YCCdc8r7zw9fGjo3Nsc
jITwq5V7YsWRNg+21zovf/SmMjNHyvf73AgVJgJ8mmE0yBXfRRvBrdMQ7jfBZY/d
XeLfQbPgC7pIdWNIph/8pn8BHhBQkfRVTZCJqeyuTd1lZZ2kCc/FdT71VxZPBHSY
Anz9ObAs4obIdE59lid9iSwQhaFOE7knCFtfcCACeDV6bAlvjCKuHObJ3/sVGJDU
I+XU7y/p8BbENMWmrltwag0+FPygkOB455kP43wrZ7Tv2swElScYOsIPp8pth7NU
rGmoUeemV1ANMd7TGsvaRHBXlZg6XDqIqrrY4eNkAKWJjmeSd8ibdhbyXxWbK/U+
vgfs5s7X6CiACSeZKwY5+US+7P4q/bwyjFRZBovzuQaQeKQ+YWVXULLFONYbhYQt
35SY8QanxXMPfuwff9DRmm+/emmMeSE0Gelpl6rW3vqNezcjFVhpOCm4M0dES4KV
MiH5VUxDtIsE2ljNjPwmTpU/T3onErNknpbtl73aWC8lGGsZy7mpc8Nu3OIh/xIV
nV7Daz6HDwLqM3FzLL/YSaUQ7DgljdnNprC8Noq+PoUcIVrNSDD2+4o6BFPleqPU
+hbWbb31fXQJzwoxwJ524g+jnA7IRHF6U4rdioiN1H02+gL8iDLe16yontJ3UITm
SsbsIk/6RnX/Gzi3lDn/ZEw5qXodQgVs3kAsbYyCEWOZRH8aiDrYPNvV6UnpH4UL
B99pFCXmqkIQifvzuQ2ipvrxbds05QxiI9bbRiDFHugNhI1OKaqJnUEQR/xFrjsv
82wR1ELEabeOHAloRNFO3v6mg9jvFsCJ+1lUip6Zp+RNC/DKjjky/CY0GPy8qSXc
nwRyNvqf4yq/bs7NIZkQbiMzX6zMmW0w+sNm0f9vh8dZDqEApWEMjuC9hrWfdTcM
jAWehFGQDKO8ORJISXGudk4av1vTU5+1nnRFCKLeb/tnRhphn2Peu/IowHyhKml9
FKLl3VgLAUQXdfgeLKtfzOckGvMRHpZy5UANe1dEUDdVR1Ew35r4aLN0EsuTOrRB
hOvsiMVdtxPvFHPckdGGO+XbdTNFXnRQPHjYkvcJNduB6ZyoeWqFXM9Iln3K+W9x
XA3iOCwCegAcmGFhOt7dt02nmL91jdX1gESXQW0shhf27aXmQtxA4ov74Ge9fMyA
XeyXveK4iRhuP4AJJ7II1W9zmWSep2GnBT/PwYspsr6FdMbk0+Debm9JlzKPRzjW
BuwtGk1Tz0FpKJk2fM+uyYhMN9zd8kFqZCVKPTVMsbBeRkHWraa/3Q/FfwFDpD0I
tu6amQcJyctoLtV0sNT8UtSqCgx+LQTtJt6CfsmH8yd7EsPrY1ek4XvrM2fSgc2U
+H+VLthx+KOm9elU+MJOAm7tFBbpZS2BptxwrSMgiFGGnx/idUJ+WUNDIBYkfF9A
LlTGApXlhwYevBghHGKJXnGtGGZX74VAJJ9Dco9i+0CuyvIFmSIddK6cIUyGhhJ2
ehBcYysPmMVXU4hqu/zTgQWqrSXLiD9f5sm4ClkuUAtgrgBrS+RiNVmzN3hm90zX
hw2lvMDeeq2uoucE4O1L+Qtp91o7+m82s+uEgxLA7zjmWMZHpuWUXSgh9RDy7OOv
AAswq+jZhk3pvxUa+7JG++wJqAMGBhsUuMvKRY0KXbo0LduHXSx1I8MtUMcZXz1s
lpTxy7fwfhxwy53+1NReC2v8IcC9zr35DYfkrsGm+cZyfgHeAsvVzKDCdSx3zC5N
ulabmnlfNJutm1f5LpkcBgQSAI2ATacYpKmwKxRW168TmaUeuYF/fiWTvLhzO9BK
ToQ+3FgsDZ+nT2GMzCFkvgaL/aaN9yz6dlFp9i1/xVu6IOJ7DypbMbfIkwuSvthX
K4K4bYHwVqa0sbtJPz747E+IVusgiWLi9P93Xbf1kuTt16/5FFmYY+m3A6YoaVEG
B1Dy7c/nLSjgHP/hZH6CXYytLd5QS6OH5GMTq8kaF1n+wDhyygKb0omL+0R+Ul8h
7TByc+ClH4xouDAElRgtJ7ZBQvQfCREVT8Y2axALsEjfH/ykj/Mv3Oqn64dpEjQO
a/lDY81KOW+L4hCCuwR/PUgzd5bwF9iLSnIOkRgdCzl9o68i3ihI1LNrOgKa2cxO
bmVUD4RSdL6K0bI/LcnH3nIUBR6OHbLAvsBrm6ZBGuozsRfECmnxsKMtnhwszzCg
lnPWckJAMczVXDOrw0SLOo+6kJUgAT8DEY2cMWG9g+iE2RQYBs8yXIDtAptuV+D8
gFla0BG7NxrC/qiZbJQZJM1LzeWqxD0Qqzu+sy0ETkBU9sDf2gDSMGl7DWbBkpuv
Slrw1XdcdxQgl/MeCOPqEliyNAVnedUmuut3UEV6feTxAOrDe13Rk07snVycY8qs
v7/Ye4wIbSG8ik3qc+8CFWsiqUPUVFiy69I+Sdt5Nsh1TEJsk9HknnU2/20J6MLh
zJWYFWPFoVFl4qf6r6opveQPB7vdWt5sbjOsIB804p+PyX/tyaL3kZk0hDK/qr8H
eoy+tsenlhKpkDsPHcNVEthZugHAZ8qtjQxa8x1xGBhzrRGEsS5AEGMIzonirJMv
oPrhECRIxpSnHJlB9wH8K+kvej84BvAVaA+ng1WEgVC9PEzl5/jn9D+NLFfqR2x0
3x7NmoEur5T+Lx766f/QOydJCSpKdWdqvLR2nrcomqbUC6KQTVqNeH2SuJP2zFMh
O1SbgC04NHFQn5CAyuXz4YdR4f5/7d9d4zikjpocuCNa2k1akhsYO9cHQ6H0lVX6
JWAyN5aQVB+LYZq2cKP/mRra2dlFmd2KGxOev9jPnlAWletaR99F2LGd2Y2Tv37d
I4rVjjXfzSFFw/QDEisj7F6rQz5kC80+E7U/CfPN7k/p8FHHrFr8YYve7E5PEo50
2OexvLiQX58ChuC+4r5AUgtHsMO/mlPc40Q5SRtbQCZ6hYwsdg7qCSBrZd9GA+Yh
ISPiH4iN9FCWKaKIY/pjPJ0XtEffw0e03FRYmP57w7hxV9O2EGfNZ7g5gW+sNeHP
B5OmwmuOrdnpZDDsvUJvVJoINGVRbB6uBPcPuHREfZYm9fwRjiXfket7FSiUmlJ8
i73ofAwkqClW9DOTvW4nNPbywzarKdKslOFRw6WSpU9suIhnS0n9gyC8qeKXSCWk
psbnqQzpNRhLzBx+WpJVSZIWwcmD2F87awTgu8F31AKdLGsBHm28r/v8lc0p+Ntk
2vmGf/vvSw21wByCxJxcyi00f+B6urhYgtlilBthbCGTUezT1DE1ZJnqrD0VDRRZ
riWK3ftoQ96oBG3luxuSWLqo1Dm2cSBNqRwCSasZmZEdgGrAwlt/99MN58PLotyh
sXcoXWAr0TAIlZN3qEKQyE1aBvx9aILbGlUIrJVi70i/lNUiWf93R8W63/B+pZg4
CoKxKR3SZBltCrSP7YS0+J+lP9yEkRxVbIfHVsAXBVfOyTGvGtSDSB4TLnydfOPq
naHi62b1FB3spEIIloL1hY6lm5orQa2zQdhRnJeg9YRQvWFJbdMrrlPPRhnQcIsV
HRVyKCQb0PFpcNicDnrdiAFdZbPTqH8Z2S6BrxqWkwEQKXNZEXJd9FoedobrjER4
fxqJz4/Y5cG+Hgf6PH8f7mLP5QS5ejI+Hgoq9y7T/hbSMwKwhDn3cF4V5b3rJR4k
f072ie0N/6hvyq5Q9ezSg1DYcmCd6Udwtg8b4qoSm3WxdoUDJwmMu42vQLKqyTJ4
CEmxWsNzZ/VttkD2P04VisKWqFAsJANvI8qEMY2WMhO64Fz3azdWZv2yvpHOJJ/k
b5fc0YFIgX5GAyILUOz0/hw3O4k+kkRbUoB4neaZqL55h+EQGUzmclRazGuv34Rj
DwCWiYQCEYAnxkJxh+9ClYQBkOoEma/oqFoDQqB7g4ybQ7dXnoKDphjeFZ8f6va7
GgqBXPU2tSO0y8VYWK5CB6Gsa8XYW61Kd9K4l1HECdxPV3VCQ6XwbL0c3fPLi8oR
4ALK4Zyq49834D5T1WVybOeOYhSaUQAhKFTB4W+p4aFVsV3kLe008TX9XohzL2uO
z/RSuHCgjqI1LvxApRjCfDgK467tzg6iU89n4YZRscb+c68xotf9a6+kcueVObxB
55D3n8Dup/bll+bJOGk+mIuY45GVvihcBfmM96PTtGMVKgJKY5/gKaI6d0wIj9SK
t2wqGzf44H0unIjsSj1xmENMz3ZYruTAvpvIFJRRUECyjSs7qJnYuKreGO0VCbjT
sceLHpkMX7nTuVy01/Sg5E+Q6xYoyH/Bdei7oyqWry8St5v2uAFhwSYZSpE0OxrV
3kDNkTXiTQET9QzPh9apeEMEz4o2jfO9Yo3sypXRLzREz0of4cxuFkMotV4F0cMc
FBUvjDE8GtBIVdmGwBAuyFtqXGp5qpM4eXaK0boFCAq/heDa+PWzH20ODHTLyMNU
nZL9QsPbMi1mzTKu5WsSTCjqTk9srk2IQFpW5HUjOrg0n33SgoYZ5m44H9fNtQBP
XqV6fDiBDdjWTEy2ZwKojtDBeEtICiGqaiF/pFod2qQJ7zT9YaFJcpvkRgg+SaPs
1axnm74yRhV3smyRYXlJjOJ9/AEdvV81LfNb4dk5uTrWxrUCBQhSJEI7oB0yKQ7o
9xD/+mCpoM4RgIBmGVUwILSaDbZJdNeP16q0vqoHbcwokBtsmqt/4WKNpqOZ8OGp
FI53Emvd0cLaPnJcJGa1J91UVTH9rocAlrcrtijFJIU1Nx4BGUXvkHnZCv6DWmka
BDtIihHaZcUorjMuU7ZhAfodkxS6jSfinXZkVgjcCW1Z+m5jgPKNDrFMPuXHECPF
0Uu2/7fcu9TO1yWHU+3CumCVmk1/APKQTsZO9WI+/46E1rGDFHIQsTayUrbLi28c
l1uja+s5plka+X2RzsbZKUEkTlDpORB/AK3c41nHAM8Gb02cdCb+Fqm/lac5qMhM
GxtmMGwBX+q8Fs8+0M5BW7f0wxqvq8MNaH+QuK+FUK58sLRrbsA35MWEqLePaIQZ
xnLT28wbOTe9KVmqDWbWCk1Ofb4lhC3U7xPZNxRzn4P2DI/s2D7MlLOvEuJNwyIJ
Xd4o9cNB/XfpLCMjt+TjKtQuIUAkYYiF19JKDoVJxHPUnEs7hdkC+M6hP3C+vcj2
v/fHcdrs4tsjOwKi7f8ssSVSdGI5CdwYO5i6THxx9WuVMIr+4lC/i52nP9mCaSNh
7eOhVwN0FQux4JOGcx7g5NCbF5b+LQs1z7sAZIC6dJglSAe7YXLvxAu8zGtq2/SS
jWsV6mvs/v12G5fk0bVkycr6llTQOO+8QILO+NXSXYZ7liVaSI4Y81/086vRS0HM
ih0on6aNtYXhOy8eY9NJUYw9dSNLx1tmhe+kFmIbcDh1v6jnVyBPlSN6Z0XD5lnR
AjcrfsyrOPEtdDKrRNjprAbTinwaLbNm5RCIewugnsSUn2hLx+i1fsath+aSTWOn
ToruL/rYv6GgYleTmTpzVJZwu+ysXD4G8FosA1ZGinObHGykNAle6v9KGV0wBkaR
jmXwx25BVH8jT9d0wLraPiyqSNknEpZn386aSqxdyAGwJQ3WrjU6uY1VwpZ1ypVr
SlYxrYxrbizlr6+SEIOVrWdPo+5ZFiBFGfc7gAJbv1Ubpu/m7T0rcAId74LU1CEf
3FuvX28TWS3tJJBxSzXkYhSLcYCCenRvS2R4/r9Lun3cZIBwgDlJKsm3XQGkz71T
4HyDo4FER5vcKq3bhqY0lhFBMd4BKnfGIkWMSnr8HhWcTRWQz/O3OyjQURdnPKwJ
bfwWBuJXjT3tVmC2L6KAnPmWD35Zq61Yem6nSfkvepqT3jYJMpl3ztB1YaXyQTEn
PPWQGL+YzqQc0qHOQu3VasJYJ6EQYN/34K54HSFE3n6jkDwg96p08XikQt+t67bq
c1111Hf7Oe/LjPwDLHAPNG9hGHhrxP9fsJh80gbST4KQz89g3+IuADEQ2whjBQiI
yD1jKhqjoOO3eGuqZfvB6Nz/ArqMWX0wITFFDWVdg2JVdr54ozU0sNhrn+wNh/WT
aeFgrI1nfvIONNW1vyppT1hX4HgthPd5x+VQdjcvix0IUiQT0gllMjeTmS3Lkrbf
fgMR1faJbwi/8Jpic1bmElOqF5jgQKo/9g+fLFy/QGGbZN9qc8jGUrTyHdK0oTVl
G/eOpfIJcpk/Wi/uVG/2KvoBHzRwtNyFG7Yna3u76O2cposHXzPM5hgscdPa1OHx
QUhmVqoi89FsS9MAXArYha1mBEnvLh43S326mRxT6BkcQDmNTdQctwzgfAL8MA/X
4xTqkbuC6e1eOhCrpWrzYAjWDrtndIbNK+az5aRdCjcbKHJI7bEEAVmZsmiIEAtg
zrKteSN5PJccEerm3qukLnkx4c3Ix2LM+JpjFaddwVDKNfnSICKlEIm19A2TPOyz
orMNZOHKbgENryM9eAgp7yGviG1hsRx7xqTKlo/ppaVBbcEFWdY/XoXVBacEfEFI
wS8bbH6KlGkygmJgJvC9r8DzktDRwKVed1W6CZdeWQMiioqKKhxCcEZGsLCE9+I0
TTjrwKqCN7jwuZ+UKPbbaHMivA00lUJJgTymzAd9qVMlQ3uEJnAlq8nSJQ9eO8Jq
9izHM0mw7EBCCp1Q/Sh66ytYc9IT5v0zruZmAS33zcx1zD8xh2eylXSKQfHwweoF
HiC+uxJgds0jzJqntOjN/eByhU6/Yw/PVGzQZS1hzBbWfXF04s7MEZVqZyt+7rpU
l/3Er8WgExrRCICyES+DTA+b7Kwjku5lf+sW0qSNGfpl91ddksWVL7bJplpOzPEp
X8FdGko+mqnM2Jb3jTjy7XJm03792d35BtxXD4bx4Yiou26GdSh7b8Q009+J/iOM
lI6qJ83Ql7DwazLMsnuyfPfMqzqfy5ttTJcMiDsH+V1bZNXe5cpSCdk7MuKicyz5
IUf4i8/TAQZ0AtRdpvOCDvtRbsMiBBTO0QtmDC4+igjKkNOwrQDc+h5oGCqTvDRg
4rjCeur2dkWllVLUbKvkl8OUiEfD03KdYcsBgV76m3lZtxjbngKTQpV0CJXCQdNa
5hVC4L48B/oTb2iUNc4HG+4sSWQaEjJ2a9/U82ps4QAkOgtj4HViXm9FeDng628p
fN4YPKbK+/R+xQ1vh3rq9Mbp18g+QLSsrCBi89p9CSt7GmBEkXKozOyI44OLYAKg
YEnMU4k8S6XeQALvFyvIvCy+77HSXVayteWhwKbGk9J3c24AAaiaHCcIt1oUBDYD
a6144GNklWdBpR8Qd9Ak4nXkcGP+7mz+goq3mHq1FknkTHdFO/2ctjxfrF8r/8yU
ASb/ftWtHvdeE+s9CTrBiAcOLtj64dEj0r7fcU09GH/3xScTz8UBnwnS4SHPW0rE
oBAkYDlUfFavxckBP8S+wPoeDCXDvs4HLvmH+QhVaqizijvoF7w2PjImq/3HemOI
P8qOfIki3BZtMMDoqlhQ5p2X98wdMdc1qjentGIo6W/TShqnyZbo06xL7+SPI/+y
hGeYiNbCDxgk+ZAdFTjP0k5gZRYSeinE2mfgzfCDNe6QlgpC5OjDkK7oQyskFAwv
sHuoS9N7aIZ/E/xz+THN/sfghul9SKOD7VkmVYXRcg/MGRhYfkYNK2+VCI69t4AZ
oynExEFLTlM4A9WrfP1UxHh1kwgN+G230YvrvVHYbQufIgf5u0awQZLJ6wFXqUBp
bQiME2xS7/yFdfBHR7J68ndrHYTJ66F4l7bkpOXmzyHM1LGlUomQ0T3+lnoVinWx
Fl0fD4Jx1CoXSKcD8bb1UxMgfjkCA5RQN5rUcWoRERHbmeiIFW+Smsv6MvJtOipL
BeAQL8Wuflx86THAC6ahvsM+sZkpIl/i8AE5sabc3lSJVmoXNdDuwkWaqH3xNxHp
wL3gv6dpeuvE2kqpVfk1DNP5JFFRToIySXOHWFN1WFtF8Cd0XU/+wNKNBC5aRGS5
/pOwP5PWiYnlHLVyi1+KvnKYnTbNfKQR/xYDp1ZnV8pRxTH08pvY7HtnHMJpm5gq
mCSZzelAfmZH6KeMPYMBoFXq17I3/YXNEnVTinsvH6VCQC//OU2EUqaYVcKKMX+N
RXeR9mtmdVKXqSc5NHbo3ZgnM7xN0LII8LUenslTVDuhrHYTdzeA7JmcYqBHVD05
FeqMpJK636P4/pcgxki/2dEPUFRc9HSGC9ozT/TqGIs29XeSmQE27XXkjpK3dAmA
Zk0AizvWw2jRTpQPHuGvxvZtxMRJd3wP/iIeUkqnQKSRw94ECI5WyglOUywNFOfq
RNBAs8xMx1HXJMsx09OXItFDIXux/zX7S2Hdl8mvHB367QtH4NI3W4+lClt6Fv6+
XGGYno310JtD49MddV8a7wVyVyQhs4flYdDeXALofqeyTXYy5pmPUv9Y9JoclFzR
QwfdMeliCfzpsvDAqWK6d4kSfxSxprkmZfXHFX/t3x9pM3ViO6aJTTU450IksAXz
FdCQKpVUhI2jlaGKYxd/3p29GH6bxhrft+7NGeuElLtLPvpsRj+pjFTCFyPUGzOI
G6rLSRH8KhyVqxsSm4WrYvdeihSn0QyNKbO0z9zep3OELW6K2gXqAvmAw9sLgz5k
qKrulUx/Bx3shYCur9N1EhBIXOQnhrXoeDU3I/idz8jc363SmwyVFHXA0kzb7WFN
c8ajA3LCkxw18Dl8evdlGupR2/1fxD2YJDgJNETCM7zzgagnRjxVPYDkpBrRzH4o
qlMo+B/92sr0tzFw07NLNaoV5Q8VBYdVoYOXI9AVUqlEnKy0KVIEFBNn4nctpEe3
2SqIiZEAs7nkCQNkLMdhAluoCxfF2OcQLP85wLI7YincCC45UgS7jXATEugnyMnw
SpgM8b9eEXQJJ5r3H2Oa0gcPh0wa8iQPQtg5wC8v5eQTv4pZ7q8fVlEI4jE5NtGn
74aGTULnGxYh7it+hBiC5giC+OndKaEK7FLR8UThImH0PnIvdyoYAfeGfhyyDtZz
YQ4biq/+aDIF3trYy2n82LDd2Fy/y5vI/2Ed/4FjJWGXwbrQMRy95paLagHvIXRD
KNgiStxYrCiMG5u2p41CRwosSOeS17f5paA1JMfIlbl7pC6Yy2Lqjld3Xw7f9F3F
Zdnt6NMlm5ekMDpqioLKBYvqBnzDoygXX30EYMbWBNAy9iJmiu6jqj1QIcctmLdT
X+QSXnjXlIQurwvaAA1P5U09l7WRoNznu6lv5eUYR6OjkFi1ja0EdJkKfGOqdL9/
lu9oxZLYTu8r3mAvenRqtnrJje2FcnifV6MkGbI/BN/3OaZdOedQRJDrs8XEX+/n
RRlMUGvh9IWwLksj7hA6YFh5pHqfS0XKROzyvEomGW4ZFi9bDDiocEJzG/JdyJXh
FyhJrzcTBDkaLNuiuiWLR/SWJ9BiS4/HDh02gfEUKhuihVAnl0BEXn1FMZ/jfC4U
lfT/2KpoIQe34i7VMi7B9TGnypiAxybz3MCUe/yHiTbiSp/aVfSFmTQLz5Jc4Wmv
9D9w6aFdzG8i8N86W0e0aXSlJAFrFF5F6kXxhAb53vqAqVNKHxQnPtwtxsgUb8Rc
ofjcOhFmP/wm9KndpEoHqT63/v2X7bn4D3WWKWC1J+oSCyc3hVur+NaZBG7/o5Pg
2Dvs4UvaI+dzdCQlZKBu5/NzwB87ZnJaFdlE5udfk9bYInYckgO5i76ktvyqQ76X
XQrT09N84wD7FA6XbW2EK9qUaCpBRjZARX+aVBnnPV9hY3SYx/+TFZieZPmPngIY
WNEEHx181CwCNOzPqFlryq0ZOlA3LjowyY1jSGNpci9BQ/9rt9zjgmL3FYYvHeox
xYFQW3kdNIn9wu2i25NH1p2Y/3nVeq7qanaPp0TQWxyTR3M4OQs7cGWcGN3iB5+B
ti1sQivsri0sdHiu4QX7TjXeaeVPwnFzu0AzY1Bd4RQopX3W/n2XITfYx6ZzNSS7
46T1cfaijLYvTWXGQ3Nu0Ql1l6Urb68wocT2dPYDdm7L12Nj590mbwtHD/tCHjiO
Qp1TZXQWER5+1mx/Bb7lC29lsLF1KClG1tMWzAVHQJg0CKXH6WQSr/GD7x94oAsZ
B83eATMyHaxyD7rpQHYr7Fuj8ZE4C9Oi8Q3AIjO4YHMv8aSVkzjvHqWNYwROM1Bl
6ihen/4/JtlO29MFLNfb6oOnKJfdyUFw51fLMzavo9X7QwpMyMqhfs4eIKG/yxuh
8+f3gzLBLBCSpYYfHkXY/5LqA3tscoFAcPQwlOvineLXdyjkDowsTsE77RlvIR7N
dpeqb0Jf3EUMXns0sF3Gm+ZyTo2Dmf893TzqPZboDJ93XNQYmgYDeZtX2wzwu+BN
H7qaXGl/3H23beSlvUmdy77VUedglpXL+bZ0ba518aZr5OMxfu/GSYbPrdTqIryl
E7ZWEw9kZFx2+px4IEmgWxY9lK5KaYN1DU3m9E6eooD8hwI+O9ZZZ5VL+U6KjwVQ
941F88BmwBIHci7xZpeef+WU6DdJ8pE/bXTBkOBrZ7D2NWJ/YYFTFchIxFdYExEW
aUCrB3JLvEDlN1J02S5pwgjh97OSNcSoo2mrNiVtOtM4Wgm7OxzKMlA4PoLdtcOI
J4cd+nQq3x8uWQSOeSXPtkSz4NpzLX69hML4e7hbUsqoDj5g9yz9Jz8JmKxYJYBR
Buo6tHzcpnRm1JKaVsCw8XKmm6R+q+017vuYvl7uTv5fU72+Ild3L/ZE0I3xgkKF
Oszx9C3YQ6KCIZZipOzZfd8f+F8ZhjffOyRwKw3HEvMsvj/lkkzDCYzPjTIXfU+o
K1V9Z17x7XLJIxslTPTiijTsZWe3kwBWRwcovX2+BsowEgREWpotaJdUEqVNiUYA
9nf1BKABniQAVYGR1AVMe7oCT51IL1LtlH4+kstAI++rptlE0a5zvt0AiEibrxzu
OK9Au+o3McRBI2wxgT17uRcEoJxKD9JzBwQdyyyNJgc1cZn/N1H3ZdQ/xcrUIB+F
JofFTEFde/fViuzWpN8GEoErFd5notQLeirSPbPnBGzDyGeZY6Xy5XhOc8IXRvyn
mzg9SIQYXg7qL/whg6j4CtzeEMoP3iT3q2B4n+Qw9D9/A6swHsRBp5ROvVc3gYzk
R7Ay38Dh89hg48hQSml84XWLMjXxtiPTSC6Hb3K4GsO8gpKRFjSC4RWdX1uo2qTN
cMW5A8LRX4qY81RhNGbnhODpc76AmRjCEj9E1160w1j0+hyV02i8uSWUjmCFc4Pd
SkY7/y8AoVG2us0rlVyOTHWOtT4QpAkRHzP7i9CPDUaSpGIrbzchp/wlu/7vVJMO
VE04XYf2Y4ohWn6EtXw8aUUgeTc6XLc3JXtfv+m6hPRuR3oS2H3RuM/8wVlTlWWZ
7zr3gMOlzXVkUzNKFOWw7TL2eC+be5YzOT8TpomDvHpVitnzLnqQUMtq8gLexsNk
mvLLEUJrYyRrTGntwXDd14mj4aGpTAwRuf3MMsZzTwAweuQNZJypVlLwasKM8EF+
hP3Is6+y3qMbgSxWbG+sEnJ1enQdKpgCUHHM3Ze60NA2apNVv0OHe/ziIV1q8CpP
/9J/nwNNUNm1Og1iX4+uX2sM0reyh9+ZxznOMaBDSsv7Ib/1TzWO/YFXbk3DCXUx
XW6kVPJJF+bSa1hD/5HCU9CGYnkBJkBU9Bts4VixO4b6XZZTa0Ic6SZKdOMBw2XO
QVgnpEhaZ+6Z9WA+HJAcoLXrS3fQxwkMoDRAtShTXMDkh98E0cRdY9v3cCEPNCV4
AA3xz0kNJ1O8qlXbSCXX3EF9GPUxAf2soJ4S6ckG9tIQFlZA+LjtxIOFaBv+RBS9
0qOrjmF/EU2c0qz9oIct3AvF0cQdttI09UH3+zfs/CyPM5ou6l9h0ZwV06F2mNVv
i1qbS97VcNKiGm1rtNR7+xTFADUj4ylr7ziZMJzTMdlRm2IBXz7Q2W7hNdO7YYTc
aNE9+OCxE6jGmsMdq/tPdtSaTK9Rm/gvNSoa7cQgsOZEv5qMbCmC7fUjwFF8xeUw
RibQhClRHF5i1E3/+8OoDNT6CbUpxPmzJVk8N87txrG5cwSVjQOWeDRQTr6qLys6
6QKPDgcBu/Zx4ypRgSyGRef2bmDX0ebWr6mo0a7ErZvLovnHclHofPrOXIoHTcM9
BuYm68kQeMbHUFQ3repKoZT22tt1Bfb/uej3u/2C1/cYXXVZ7KDQamrQPMdC/q4O
+4QlIGwvq8yYOkPUYKXY3H6EZs684/ClfSH+78Pkbgm00yG/EL/KwWaSDM58H07S
f99AwexDMLPQz6OZGBDjJ3MkDz40+/SjM4qpxTOgrbgKjtlua3lLoK1uwuQN/ban
zEKk1BlkbbgZdwgJBtlg7txK/LGC6dO2IR6vNrDlkCH0djNhnd7WS8xcUsWzBUa8
CoMQOSYm4L9lGoBYelVyZMKXRcqCn/fXwopAIhMHRp3WJYSk6eSYqI5/pi8hPffJ
0Ju9Xn3mYnWGC0NYEy5Z1J4OuoJ7tPMgkEBS+ETCE/AT/s8P1q9w7ep4XEfbGnCg
6r3w3YQw2t7Wy0ygTjNCJCl2naAWwVw7i+BsT3+4q7+cZw5WafSdypJzbugFiPyV
khlm3VCpcTeHaMUvKff6vnmwDxFkExFOi90ccjMJfKHNxhJplMHNjlR+7tFOTre6
Le6KdSVr4rygFtmPtrjWr5XfWg6FyyaY4kb2eK/ub5p05HsTzAriFd4Govn5TlCv
yeNGrldeGvRGRghSyLqlQvZUP0ZHt3syhQRrFqOvIfbXUaTJRvD0+Kfh13+32CYw
vVsfwLn8AGHRFBxWIIc+87KV5tVhwSlPfVUVvGw1CaK2gMoC8LRIDO/g/FcJuSMq
bKvsyicq4gJ0zwOxHKFNsMBCqpYdklNOQ03yP+cPENI5+cJ8LZEin08C7Xp8psaT
r19DZbq4JWd64NkoKsK77ewV8+ziSKg+F+5m0J/r7XqDfUAcJ6YxQsEEsBawbgXK
VVKBmC/dzDQtb1eWrWxZC/O7GjjjyfDAKIMp018gMckPD4f1gyT6J1DjmBt4Q1RW
atzpu4InuW/NxmiSzARb6mM+hKTGxecvBbvDj24YjWhMu2OX/MOFlGs8kI/AdMc5
EEkrViEaeG0lTeBLUg7cVL+JpolfykShz1IAbGDFOskIXUKSmvBQqPVqP3M59Bfa
l37cOlPxXCzOyCJmxMvo0BUp/Rpi0IB7HeJE9SuvjZvAYnN4DGi2PpLV92um0Mg4
OlFiaeFFSPdcealn81PKaSRY8nGwIfQmdD8/VJPlJsxw+D8E2xCZqEhpfw0afHAK
6raEWzzmG1eyiQO02SfFKgCV1MrEkwfg49IJGZXCURvd/q4jw0of1C1F+oEBsY2I
hHcCmesg1tPdJ56nXJx81uSLf2t61dhnnOP2wT0i+uFXJduLmYTiHG6Cx9Fhj7D2
5rQSctsSbmS3ANwxsxq2qH369i5Mq0PKw3v5YONrQeRLtsCDkLXCFPax6zhKAPqO
7NNt6o/+u8KDTWb7cIySe43rLQFtWR3Q9oh8Vi+iGxFbkfqxkdXGa7cP1g43pRW5
POOX08WujjpRKOqlcYZiryKYFaT8MhNIZrPQWft+lGv22DQqTlGqGF5gs71UkIx7
Wvdn2EMAGYb/fZL2V8uhCBtQYexMVyoapQoJGoX5mCaA1akhhJln06bEUGYXyyZy
ug5YNx7T9OwAxdSTwW1OSLg+blXux8OXsvUHyJo2VQUUVAgAGoNNmkkOKRoV5fIp
bRmfZg1G5P8RHKJCqC14IzOyTXD5ExPw75WP74q83Qrg/iBjlkMJdrwCWsf8DYDs
UA+9PiT3hBos3K/5dfmY9OfHw3hIc1gLAo27DtYS/sMQRHp3FUMVHsewVFLAgYrz
0Rt42eQGqLS8u5NSPj+6UiTc1TpCezaQYvXqnUXNj+S1+i2zGn1Oa8kTL53nPIHI
bh3R11zZB7bbr5Ve2F4DCgE6il2FjsPN9cRRq7qRRdaOsCwMHwbooUnoGIqogThE
gGdMxPKOTBOJCMJ8tuv8gfN/Yqqj7Z1fSY8ds5PmRgA74LGJoETxX1X6yxgR1TYR
mcEWkPQxaG/f9f5fAnEPU/kRupKWLpY06pnhVCy/pwKhhqI7V1VGqu+e5r4RzfVG
+Cr8+DQJh8yDGkK+gkHJJUe/gmAEEK7Lw8XZNlUzgZ51qlckXUg3HNVRG1HJO9/V
+TzGC8BKFf+ifRB7xV9JKt8HjH0blGC54qSIDMblISeNT5MBoJtKbLe74W8IR3T1
CtXee7B0GKmKthnwIHk2ixuODVLOUUImHzCc8kwDt4d7R1Aen3H/LfDKeSmyn0Qe
h4/cMHrwaYMMYyrV3IiA4an8PijOZwwaSIB36t5cLg+pOeEtSYnnD9Gnt9OyTKnm
ri/acZor3/z2herfONliodBvk04avoObp5e9FmiHJ9cgRJ5D1L29juanii1j1wZN
Hq7FCBXkDIu5J9lbcfbCJIaA+wkaGrULnBMdj1/cgDbj4xGfZryinSf7qEsoaJxE
QeY2CVKBwzQQc/losALJGHaEfaqtJ/MEnlNyLjaA+lIe7VpiYPud5pZxzboqHluU
Q+nen7UwArz+LGmfVe1QPqe7oefkasA0Mzld+5MUQduhzJyT5q3KWmqz6uahOsAN
PXZ9de+gXc1MCTAma1J+zxIMydiQWBglGJEmsdXPsPtc3cqV2pEyJV2vexoffCPH
JoLw6MUXVgxltLZVwxCxV5rM0y4ABpUIHZGc3TsHKIbRG4zHP4DlRZNbWkveeYHb
vXEKAlIfMveqdpnp6DUfH5KO4BnDbpqF5OslkdXrOpoXxkRZZNMlewRNLqT6bRSz
P0plpZaThzIdyjSij05VYl59+LlPnulL65vCUpZ3bWcFHYCEIJX7V1HvBVKMoRAV
DXBeKGMmzL1RItnmFjfn2yLEpZxNFUWUFRgPNhcKuUNI8lfmnRIet7Rm8RYdKk86
k21DfVL90klB63RZiSxRUxxlN8B9z39dMF9VSSnZnevPRzZK1nvwkyE9m2k7Ns+P
KHL0Gvsbk0/wFr4oq8uuCYqQ+6NJ8NEPljpTHMqoetSK//Mlpc8GhyYarDAiCRni
JwySBis/VSNL66AWD2CygEI2xrN8T6fa/j09cA78m5qSjGSOI7InUfJwKtj61ND2
uoV0bb7Yc9wbcL8UNdllPQhmGcpgZ9iCaYtnEXNY3OykfFqfmVkO/xdyD9McgJKL
8Chsr44K52vzPhFReJmbDuyWEAb87wDBAxil3usmwlBXhFfNnFim+IWRirDzi6tn
fU7KVdCqldNr850aG55x17Ts//elZ7/bdFhgkBvE6vH1id6CnXYcYIhYmThdORK5
XZR31YpGvxc1t7EPAy0tJot2RnvtXDlYb9cnLbuvG2vHim1mHqpDsU7w15PfOM75
ukqx6bpqqThXoO+2QeTX/426EzSK9CK4hm0yxTUBThB0o0D1qZ65ISAHj4RXwe6W
p8O69rU4LPIoVHWI3t/Dzvc0v6ZGuL8zPKBTaOWH6yLE1aFHXdOnBwtsdv41bsRU
BKTWUrrRKV1XDxGN3uFqLsAHhJh6V7Dxl8CJquPlL5EeUt8zlRkYhsfrgmR7R0h9
8tufYyK8PB4xfVJDYe14/D3y0fXRTUA96ZraiU0nedt4MT54HCkMdV+yp7ITzlA/
srix6MKsltVDV3iRFCEMdxjtudmy17lAuuQPQG0uK17hPgegqG/ucP0jyqZD8f1S
hV637PBWWqNqA63XJW0X0kdLI/mQ3zaP0YnyJqevMrCyHCIWTa1nfoCB9LmwY6s1
o2gm+UIwi8xQOJ5xlPL2kd4q/acyIhVjpM+fyrwCI1B+Owh103PycqOt+XtWRVzd
I4BH6e/Wtq1bUshOpzDi+6uYl1lxHAbrro6Toe/8AHlKAr6p8wmzn8HfIZOx8gOc
w73EIkS2LABWyFfr7MU7rRFSxFn/TplloiHYwKRFjDuezkMCTvmhj2hiG1ygwavP
09jukRUYnZ535oR9D66joszkK675ILnukTf3qiwUnPhGoayKS4iUhlWu8wyM2c30
f/Kb2D04mVNApS13ka4hVfxnWwqhqHSa/jnitWR6o8mpjf2bVPsIpgbt/LBiNI/H
RW36vQhNkmO6kmMAOUlWotvaWq+tPGaxiYuQj97y4QscUYl9JGuNHOMjKlxcd2Ax
6yXDzQ5GoIR60d08qBdzS5EROmohp1IrDMDmehmCtTwpVq5LwCE4Bf3oajcC1btv
H53vMYNTNTwmIhsgmaTJ5mESPIj1VloHiADGXbXlgUcH8faqkuzfGXLdXIYHN5/Z
3zo06zSS1jP6r3l/O6dmQ/pAtBUFCF9fOdoBwd3AgyEXtcU5UEPUU1vp3qUBYIUH
wiy7cotuVC5h6JKF+bV4ib8JGlcwLgS/w4S/DllVMLaD5qtQe0TS28kXbdto4Bhf
PpUIg6BvijS4+e5KLJVBL8u7mrz9Ln02exHKGQTyKqtdA5L+fVLYI7fbeiPpETz8
ghqNg8stpg23Ovb+S00r3VdY2flM17P/4x+JTE5mgwjLR4QPn6OBh6xX1npFmu00
4feljPxo1r5POitbnuxDmq79lRL/XtWRxJA9e6w+wIyGGTgM5I/bi5L2iokcyWnc
DFcJjmU2Ll0aCM24aW5vbk2QwaG30filY25WsGUmPrL1I3BvyVIqf0jljvzWcbSX
DDm55F/1xoxG8B08kDY1JkjflswIKzjf/ITKNNlGihp/CnAe5+JCs+ZTzJ1oKbyh
2bMZSb7wx1flw2a6NwZA2wnwnaeL5oL/bY166XFvPGF8UPbCuw9e8QAtuhsQXqBL
LAm2PTQzuej5U+31mpDpsDiiwiTbwC4qrkrYrAtvtjxEJ3fqKJCLY2o8ipbiHEfO
urx0v9ZGh4EQVa0uIg5B+KJp4S1HU2u7MZ5qeFLjAl7un0/K97dXQ01/VqUkRMfY
sHjnLX7n/e0gp5O1S9G8ii+VE/PjtSCGJO2xBlefZ4nBNQ9MztguqOz4jMMhEmqq
cyBzkONzluUbTQon+o5KCKtJY9nlteniqys42Q4Asjk8O+sVX69RXhyvKa6qAM8A
akb7ULc9EKqud7SrW+U47AzINAGCEYct8DZ+g4Ca5PQQBKVVxOpQYq2jYUcH6Ipl
/ztlajebAYwYUmbT0qW43j0AWuaMwROE/YpSpWLCfsKdBKvp+6TE5QNUjTWvg/Et
FC71IdgSjVky717VC7Xsdx/WZoVsNgvuBgzKX2vZiwMhIvYfWTMcL+EAeq9lvB/x
s8Ia9MGOEKlS8IkNZUTth94cl9GZc7ozI8a85lM7oTT0uwkDK9YCGIOT3nclmMUt
b3ouybMD5fU4HnGrqLOragp937bK1pSsFdnbXV47qPDDk79ieAsdgOWQgTwQDna5
7l+1V9wIY0ByfFSpkYnqKvcCSpV0FAOGiw2qwnCfC7iWRk21fWlmljz52JMjaXq+
f7I775bjPEKZ5XX8As5z1c2o1ZbEb6PKInFklQwqFhu7/P+dERAxkqQZHvHrx4ke
Nn4lm8IvbGFt181I/OAA7ohUxmAqghpHmxlCrv5POcAnHsfG5izdUXfvkNp+UF8f
k7k3CZmTCA65C3FP3UYT2mldtsmWnsHKUU6TKBbMN8wRCwWUfO+4wezhvuDDJuPE
VCzXdu+EpjIapxzhfe1S4ZCJvSg7eWku39yPiU1tb6UfZHm42tNaaJs/OoLkubuA
jvfK9jiN7YItpEjjv+a2KpWkleorgfVZlFr3qSzglnXbt5FYyrp3rkTs8cg5NgOT
K/5So6aygKuwIuJU1C4geOVgPLA/PYfV02bDOypwRzyOpQE882IQeOarfZM0lXGg
dJhMr76SVX6rAp/6DOB+cY5b3Vmpj5/DclfF/7m+6/vR0PrJtegwTqEsS/NLCU46
NxjncX08EWXyeSmIzSo8ub/f0LfTw0dS+3X3CuBhPa+W1I2hYv8Vk9+mi4jcvf+f
PS85W475XYDASywasxBSh2xks3CU0Ec8cQI3D30t48MU6LbwUIeDd34X27AUMP8e
xasxUJGSB0+FXTlag8SWOArX0khdUjuhN+pfBOclFL27aK1QwEMjL++Si8HRTMrs
kFuGegzJLQu7iiYtQUDsNvh4+7Fu1k0gFfncz0pgvVm2XTNPMHZGcxlYdlZNoDgx
QhdfN4+0Xpthm7uBsoiOWYQwZfQZI7oVpGWDrWDvflv29kLAVCbIu02YkoDmkxKh
VimbxXX8D1IAxKNU+Oias56gksYLCsuMAwZeAoP1PxfUi6+CnSA0fj5GtpxREMwS
AIezh6/zjky7IzKmQT+wmITBwpDVSv3axvFUi7B8+fp7wFdeTPDZ5Mxd997pqLeH
+lczxEg9h+I8fkltUDZzNq7NTirIMje7RJ5c1kqHszjUJbjSTtvwDM+WbrynQirv
zIPJNrZVM2tV8b22SWKnEUYJZe69ki8USFM8fBPE71wN9/bFlNtIxqrCcmxtB4CG
nrv+LXrDB6bVTcBnpPhAdBwo5tLsJcxCMplWkUb32LAKJQ0cQigoxAgKqPRKyPEo
Ijaeyhw530ZLaMHDp0zkhA26Yetw5UnN7ZhQy0UxBe3jZridqrR5okNdS6pI9NUy
pLPfFNjSygY+kzCZ4SB9ODUOX2bhNUZm3G5Nvs+c/qo73zq1NPtgoPdgV4FI6QVx
j0d+hTypE4xvpCkdFugIYnlug4VbcY9UA5N6+xb4cp7r/V3/mglu9uxkhabRLv64
vwlATxYhm8co/Ehtskxh1eZ07oO53QtNMoD5UTrVlHyppnVCEasQi+JpktkQDxed
punW91lztYJeNQwXkOqvU1NRC8RK6tVAdNtimM6eZQ0UKY5Q8HYLq2MYGC3IAlKj
yOlDDNbYi2meiYPYPYSZJw0E56AlvjQeTUvaohu/Xudgw07YeG84P7UfoVUpYueX
WgbQQbFH40xIehZfiX0/vtu0ugR+7na5+WPNAtzK2Z04p3jHGuTYLU29hXutylSM
k0h3xYMYlauPnyCeSf0yYjo2Fe91/99yLITyx6W9TsRY/+DoClIoMeYIG62e48k6
1pvECYS+97rgFjaLSFlvvIKScNuWSmNB3ikXnMlTUQrNcU6Xvz+2rhRzONOyvGux
HW1PLhWmCt6s/x0RiC35vS3Ci/9ldOE2wHPD51IexWklue9lE2npD2JctNPhQV4t
20o2TZuPDaS1JFACSHPMDwIte9EMKedwraAEHbL54Sj34HlLuepUi+2srdN5R1FO
lDgKw07ii8nSs/1I067S0FpTGDeo//tiJVRuW0Hh8ZxvsBnI7NFe0VCNfaP51klB
ppgDutu+ABX7TPK8iAzVCS9kqEW3GoF021QL/8B4zTpEi7nxwu0ByjZGE62PGdON
Gvp2HNx1I+1Fi6J01t9SsfiKBrXAbfrup/G08RaqMfI7goWrMXFpa1ZbGmeAb5B3
kbWwfYeXe/fdi+CFuA3NY+twnVCGPatKbznwPIEHOaBy5GF3jRvNF+jrWvHNZBb0
nRUn/hgrDepoBZFF9Orw2ynMnStG4UDg85ktVTCNwoAvn7cWSI6E5V60P+WgTPxi
HYUK2Jijt4IBuuxQLd0DdVgCgqKOx7KSozkZlHAtRKFGRTLBmcu+IlxoUemy7T0F
euISo1/RnVApB47mALxOkwLcVCGkxzmYXWC9qwuhlhCwlyhI9c7vbWSNq7MG7WsU
/3sy4qOylHEPP0j75KG/YETF5Knln1SOm91afpkU71IkagnCP+k4C9R5VHxaK5rR
4mEQFbHTFWBJCnuvbZQWY138uW3r/Hjk9Jk349xNYM9aee7DBQGxcMGlhI3PtrKj
/aKh675+iJJvlZNemB9Mxi+H2IepwBg/neEhxuv4USHPrK8uQd/TqSSneZhIsxhr
Wcgo7/txGzS0QAl4lJyNqemF7LuinP5h0jYXyCXNbKw0omPVxA0KL5TtByHsh+Vt
EAfhCdLyfPBjcGncagRqoqkRft5uCe3tEFGW3pBiDaEY56cAHle18/T+HDouNhiL
ZyxDwN7GgIIRizpJZrVRLPV/lUUsK1RLzYNfpL/ysXlvu+rqAkZdhGKJxXu1EKML
a+gXjqU3hGHvLGQB38a8hn1EI3Me3dDMCu2zMpSKWkW4gbUAsjuXOhCxasmkpbZx
htZi1UCat5FfFI3bvVH60xCfehJOJuLr5DnVzHd9Qwbo6gUz5QYPbET5NnnK0+Q6
COQCJrFUJLVGLGc4htqCRB2MCkcQx9G4Km9EHQe9RhqDki2au4bP7YL6TgKa/udO
4OJadua1sDuI2GREDUPAfICwqomh4gg3xAW7wqji7Uk4l0JlLUHQruqT/qQ5Zqzk
gK07RycCkdnAB/K1hoRVB1zmcoKEllA5YwNMspxq2uKQI8L4EHRbfXV7bv4f8/bA
4Eg3p7HF3+Sc7IGnOKIE1rlI4OhuPpIqKlczHMAwQac2bpB73aAhNxSPdKA5vExA
Nu7LOw4/b9jmeb9oNHG6LqCvIA6js3FhJDiSCfNno6FQg19fW+33xYVx9g71Wml5
wNOusW7dQ8V411EVbXbfrWwYVpJRF++VM/a2mwQe0FR3YMq6Etv/eEaa1CokU2HQ
KDwx+ChxnfluTVKZVLXnQpmrGQQ/0ySh7mKaoXgjIFviiH+ZKljZKS0qJfsr3P/d
YXetQwulsei0HXymMpfP/AQEcW2MRSo4dmlNApcaeZ9pviDYGwt14pPaGhDNjkrO
Y/ge/AwNfwEhv4cz6sG+d9fpGbK+mittwIDUgKbZbKYNNPO0axdp3FxBsLtG/SN2
6g2WvSw1jYjJRNwwokeoGxFzn2efG2ocJDZWl2n7DooR02gnRlCl4NJfEIchYoPo
/Sj3JLs8zVsLLv5VmX63teXRTCmR7F80woSwOUGaFAl0BhPr7Th9QpUAxv8gduzI
s6OIWeXkAm9G46QzW4ZilqgDOGxE6b1fVosnlpnwFpiLwSMYMNaB5bXc2qiLXX3C
NMonzkIuAElOUn0+i5DPnbqijushMPNfycjkQNbcGF7+GcGbOL/Laim9OX1DCT9f
YIgUl5JsJjuwlikzltcUuja9ezc326hIYNlt9zF8KC63Rr/WYG5uvAQuV6IXaTes
HBmxL/Dh8d+4miDTI5ahaCnulWSj3k4VME+P5QufGV+WixRGp7Eek05kzW8p6Dtq
LQ2SHzkubIMtJdDLdibGFjr/OsWLZDqBZ1ld3luAIK30XaLYYFX67NVR6aqry4ut
Ad4MT4HZD/HSMkcPAptst8rHMNPFleh9bZr/nSL3eigBnlRdVK+/GgMO1VkQ6ni7
eI2fxOkw8TqK8WyIML/ykDJi4RTT3kEYIHTDaHlt4sS8EgjX/HiYnDoL8C8rjh46
U5/fz473FnK5oM4Xo5hcRQseJrLfHlcq+UDTKS5ZVxub8y5Ee/Xxx1zavYPH+lsv
pHvyr+xRjOnSCAFIFLCI1dW2p13OkPse6pX5f+PcuRBuDtcrbPzeS3z3Cgd06pw/
nBv5ksLwhhOqE3KlHBnyGMjUXqi+Nvhnfembt1U54Qt/2KWhZpJh0fijFhVcXqAU
elc5kuVIfBA5p8XXjKyU3Uv5F3JfbAaQE+0ZeX3gMCSah8wHagnSTSBGbVtO61fU
JQ1fzQMpDdukkIEKdZmCv6jOIE4EC8VoboVtweyyCAoxnqca49dEwOrCTzx73uui
4BQssz1y6jA7ujGf61lBj5bOjfa9HaEDdBDBbUY0pyfx1+rx+IaqOL6omhTfyCkc
C9K4lMUAy67Rp1MofCu0O5O4sY1zRBRaYf7+JUlkh1RD1CcJk7szsrSTHIAr3ou1
R4m/Xvqb4+8WeFQzzUDipqmN62hlvBaNCUbVC/H5hE0chXlosoAWHLS2ft7/p+s+
7GyoOp8MbgAbFPXIGC4InYFUIQJKgTGKoAAEfCHmjua9pGqy69qgSAxWDXvS5sIi
A1IvjBgvQWt1fAbxwKx9Xp0agvwUOhWPCtPgSwGZR5Mw+nwL+79CiIlX2lfuqdvp
EDF02FFpJPs5ljPBZm2+mVopX3DQFznwN0/fVMbbvOwQlVHy9tfY4TnAvhWTIq8w
N/71SJEzB5czn3w9h9WgqmO5J9goAnqItqsCQ01CKepKMkkDx3/Jeb604QvWmWIO
77FlYazT2Op2bg1yh80iQZzGDcfIljh/eAKCK9CY0jji1gVekmFx++MCqTB0jMlb
qKvtn18ATAo9jZhkp6dW3/PVw1gg0eQYpTJzs28c3JCRXHkJewVYgLun46d52K6u
O4y5yC5JQjWJv6cETJlJYOtjZxHo7PLM5J503PUv7XWAZcQFu394ooakufi/4jqC
skvMGDCs87u7ahoLIDW4kN5QVsnWRMngUVbxI3KQL5zAIqWoshxSX4tNTLTaM/kc
vUDp+wI1AVVrpPaHhzEEygTPt1VujPau0TY3uht9gfXMXf5LIgfOAfeWlTUAe9e7
xNNAZWg4oHJs/vGeAwMkUiJRhwlnlMB03U44R7rPmy5eeA4CqEPEaaTOY1/8WcDc
2nBOg36hzzmE0EC98WiNODCFuhi1NdLEozSff4BvxLlhwdq5i/UHZW5i74Dmb2uT
/OCrGhnolmFl4R4B679UyZbX7gbLUzSZMygdAoAn/K/B3T4jKI3OMVD3STY6thQj
UgOpdjHbXXwc/k7Lml85+x93YqRlJW8Kd0p/tiMQokJyTqaXR3ww28XBFKYI8Npp
QIaLcCjV6mw3lmslaPQi7tzG+Q9hXGZvye6/8vClDmM=

`pragma protect end_protected
