// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
N/qVvP5oEWMuU6kaA9xgmmgIyvgqD3h92nby29to4cUnxwo4IJyQZl24tG/QJuCg
MSjpVOZWxLdgrJuE0xxh2wjFZVBd0B3zHfgM1WO08VxthvKfRsVLC7rotXIQryl7
FCOj4xtzhO4Mt/9tHk8Ak5Wykx069hKa/9i6ZYb3S5rtFXy0uqVU7Q==
//pragma protect end_key_block
//pragma protect digest_block
SL1YVk3Qzd5z3gbk47hGLQE8MzA=
//pragma protect end_digest_block
//pragma protect data_block
FhnJc+fe/Zp81OsRKgWpB4dDzQR8EzwWmkL3y/VoqW+hRGJpqceg4HLrqZ3bUSvJ
xkDDLDVTk+Hklk5UkutOk/XCa6XvnVJRa04CgRgqCGJ7RdaHnojILXIHw87sKE3b
il1EeV+6SMXDpyi/pMNjg3Whcy5sbzoOAA5ikcLyxe+3dCthaHiEx4RE2HRWeor/
RL2lnYVwHsZgroU94Zz0nOYzYqWMMZpw7zAmPDPlDJaW1IEwlOjHImNJ1kEgvFCp
qzqdzDJpd26p9VKIH5vU7eh/jCyiQS+A89WulXci6S7s61qdtHc6yWbKNSclA1qn
LY849ErTGUqcXOWOxmNl+Kq2BVKDKU0iTrcx2fbng1yCR7GJXt36ujd9nbgN9eGJ
WPHTkF20J7eCHCF0pliCX2qFsVvC+lPUkN2gyd2BiztNykzbgLYXS/HXpB98ujUZ
4JQuJ4h/RWXSOBtiCzhMUCy7jobjd+GSegG5tcFgCnRyaQ4GL+DtK92nwvyNFBIj
fuLu1GSs3KAUoREswvi1USasNnKkX57qJ9ydulqP5nIXOSkRdxq7B3FU4yIF0VEf
E6YZDzB582WtcwFgCZnIZ1pvPVdLkXdDn/mmy9X8pvIYIXBQ8mfPdhWY25SNP4TV
7Y4UVgtVwWM1dOQV6nuMvcFUMte4DGRcw1uOkWRqHLW1zHOQ9YRFEvvAXW112jCY
PGtVYFlx0aQtiy7y1k1FX8PtbwGPOdBz0QvdwvcVhbQwft0mgtsqxY9VSBbomoox
CTj3aBljOqgKS/1bNSW+EgsIiQBV5yDujZ+JHrxH2cLzag3gYWGLqJqfYkhi/D2l
jBQp+p9ugc3QZI2uXQNy3usvJuSm9ODbLo7uFS/ukqV3S7sfMgEznWLxnyrSHIJJ
rDe8RB48tXFAxAoX8JiBmkT6jCyoY+fk9Nqo4o/sOLdCYrBmCLlM2BE6ol8Qc8aB
DRrq8uOozFoGAwbqnaqabtHHsXrKVpwZe+c6dvnne2pAlPTAZkkzXqX/eh2JPuHl
2NPYP2mPWbBEntf4TLKs9yGOPzcs496o1UurV974ZUqe3VOXII0augp9eM4d9D7U
XJ6TOc219acRp5aYiSgf08maMOzCiS9a+opht91rDC88S+gtxa4OHn1Ft3PibioB
ycVm1ViCjeq9WlAUp1SLPILTJv/VwupWoTRE85jYtvmkWZeHSr3zMfrlcqq34kHU
W4tO+0cVxkhRvgCqGoG/ub/RZHQWeUdueQpSQpUHi+u6hWBDxbWR9AayDBvKmg3G
pu5B7xoQXXdlmDTsxQCr6kRwhy89nBUiIqyzoTQOD9QP2ibIlyD+HkVuS/Qhc5Pu
5p133ueAM79MjMlXObsx9UCH4JyWyC1twgSQswdnCHyi9fzM8affusbkrAtdhmxY
Z2DYRqiJs1fSBUKQM0jiyYotK7MqPZwMe/UL+PJGTGJYSSHXNbBNXUXjS6N5aoiU
pivpkCwgvN590KTgFpG430uwUW7awdI/87uy+wJXeHHiebhUV5vLgNkrU48hxRpo
as/lf9iq6/JcSMHfouzdoiNIAeviWzdu9CUvwLPvRTnIGhqD2LsgbZEpqIziRTFS
qWhZeUUiGA5c1353WZezUWs/KSduDhFwztv60ygZRQvQc2mJeDXGXNIjQOpQ+/8x
pE1htUSF7qXT7vyyJHqwdb1M0oK1nim1TSL7wrsdt/Ql5Wp7/S3C+N2r7IbKhF7O
4lv1CtHCRjRUdSJcthTa+c017GLcjI3MHTMJpFuxP3tfDzIH5joIXIDEk2w8o4Zz
LzDS5mbjyD6EkkZL4fLhImsZ6XSd0CQj9xgGUl9QXaQZJOc1NlJic1icoJt7QZSM
wE2oswjFwVhFdWpYrMEXYPqizh0nYPdGi4zpHF1HIMsSgHk+Uom+V17z1Hd+GOzE
n+RQK/0ZBfttpmUPmQI80auto7ysXkiBdwqwz6ZC4RYPAh6GNEa9p/9soJLiKD4L
z0v6TTaxIuoCWTWg+tDGs554E1LWA+lfOYY3VroEaAR23ELJdBQBEefpQqOOhIw7
KS7iQ1thgTu1GqmRX+q0p+IT1gHcZm0Jl3c08KUEJfHaEuL0qEkITU6o9GCiu+vH
Rr3LtO64Wxu+e3ZjlP1Z+T9Y85Io8Nes9K2wRDcHWGXIyV/rYzm9q7DfbTLyPpSa
cbQnRa3hibroe3LcsfxoihLCYQyW66rW0x0AEGXAeXkUZiJlKdNvd+H+1wnLcwnU
Tf/ppgC6L9cL3VcUXrUsI5JN9+ypdS4Y5HSWS7uQCQPRhcijJ8hqWICbmhNsrANS
a7s48PVWK/ZSp64iSg5nQeg4u2lVH8VT4+5HpoEh3QFUKoPhzzobfwbrHRodpFU4
v9Zq+V1XJsFY5Og+0E2Hg8KS0qR0D8bFIFev5iqTpIyNbmEpGyV+rOsWFRlsae5V
bed+bWcloJLE2zb7eH0UBtIoKosNTC6CbC1GwtmBorR+vbr2aDSMoSoj1aOdqpwe
DinxakJmGjO6BPy5IQAcR4IpJA6FuikZxN9wM6fGS4zgvpk5pBERKhy2PcsluiY4
dIlis5b1rcgMnXnrXyFxvcsU1M03HxEqVQVhQnP6vxzES+UT6axrgyXprwokqqw9
M5UAq79lrEHQyCipj9hxgad0lent9XXj9I+M0vLeE9dHcA8vI2eh/+PDo8sgpIUu
lRUT7bU0NGS54nA2kCRc1KF6Q9cAjtqE6gUdBG0hNpXM9zKxcQ1+2YfmDP5e84Z7
wn2m0fBDHMIyITC5w46VnlooefGiYqiwI+f7S1cUxTr26FDbrni8X3VxcqD1QGMy
40dxYtRJLB+PVGMDbALZkNYHkdK9d8R3PEv4qT4P9/8Kde31OoijSi+Db+/xwx/t
acKeHE/W8ToWpB+57liLdIfDbbeMp++JTZIInIAEfZfMKhLgZinw8E8CJu2XlkHl
K+xNdn/jjl+zcfYl+LmOwov4kWoazdNeKhugxm141bVOX4lpJusnDY1y2lOGPtSr
k9Y31fqccZKYDOnG27DAWbcUPKCzXv7zI93kYqI7Lv33VnyNQaI1BhIlu4U0LWiW
hPkHty1yoSh/liLG6YQqcjgReRxTBcjP8upENZdHi/f5phChpEuUZmjcTqGv0IqC
b+61XOcnK6oTqjoxpWkF1dy9Qo8Lh2Oe9zLPDdGPBFkJ/3sfoOGbH7kjNCAGfzF9
QiAvFBQEgNNdmOJ3pGc9W0F0YNhCYb/6NjZsTqGhIvEpr2QZV7A2wqnIxBz4oZlP
Fd2ClHouIzzHo9dJE1voHTJTRY+N5/E3D36s2GD0lAm5ojCaC5bmeI0y4iKBDMPm
uSzp74ZrMazF/NPwx8h2rslxvqroFJQ6X/NgCjGHqQp9I5v8Cdznrw38dM3EqgAS
sS3QWldP9nfX3XciOumfZFtnDY5LAEbfNto6+/HsJSnDKeEOUp50TKlPjQZMNZ6K
QGW8s03U6857/w1neOaF3OgTOp4C4AV63yVqGP0aymLC8Xcoid3xMXHCJOzZ4zCO
n6r30wQyZ4JkDjK/wkqk2lKK8PJghhuEx2ohjCISC51CZprsY13cx01gSZEfSnvW
j5CKS+3JAdiHDNN9GiwwIfqbs7haOJ9bjFbJq+fxYt83SFyHiGAuK1oq3DKmdQ2V
hTF/11Ad2+vN63+PMv2Zexkm2MHmh6Uyi/AU6coSdrq07OAvPVOFSfyXLZwxUpKY
6aPsLBmnUQBY90Eyfe3RNm5RDFdwSwOBpLZGFBkoYA2EMG17cVKOj5C1bpbv/IYc
ZOVUPe4fielvnKdWBQ8phHqRYhoOkXExw9eoy0P+LE+uVpVQiAIXqm3cPbliKeZA
AbAfW7epgh83V1OyP/5up7j13VB0xr8vzjfxz7IUuFKAMTrHPbfBKNbbKiIy1ni4
DrTt3SFB+HIXLuDsU6o2PEwPENOMlJo2KTtUirhGc+sKrIynd2sLWz6u4gCdCJGG
Jx43DW5e1CPX1x2FXw1UlnHZsDr2dTDQPRdE7MEVoRePBS5oRvy1kb8EPKGa1d4Z
jInhGuLCIvUxjL8fJtcWRVSjQvueO62CyuZqZAgNXJvnRVzoPcEP9jKsB/ERCPm3
9k5SsZ4M+LoTuFNCcgHjvWQlNAEvOc8pR6Z227hzrYymzEloJYYVXnUWByNCn+sC
eZHXIkLrT1hzAN510lb5f+XMkOJLOjqYRp5VnbWdQsQqyvcd/chaHj3CLyOuDWRx
bgVlbRNwgRmShWXVw0zKivFg8fzYqwQCJ2kNAnRbP8T8FARKugDpg7o3FjD+Ajmr
7oovU+fx1zGQrGm6QSOxeUj2hhH2RaIxMivpMJBudRDbKTNWfo5Vg/x+tqGw8HXa
njTa9Sav0ybuFB9+CeaVYvFSntuO795fkyrb5W1WB3wU39bScsxkJvl0sdyb9dDs
8SqbJHkVE6G3CA6j+XQl65GPOuQovKSinvWp7uDOpj0CrLPFtEN0Ip+DzrjwvrxT
T+3d2ZdhgplyQc1FwbGmKgr8ax+hgB6Y0lDnQ9goNSACj1sPYZOlZpTqQ+iQB9pL
8zO8K2cq6kZdXZkLRtgx60i9Ob8oVFU+9WkoHS5NhbxfqXR6pnUTedUZW6/xcxuX
K+ye7I/7fq3va7OjdPchuI39pJeavSy3lQZ2FCC6qpt+I5c1OSNLpI/s9LyqI/oe
3yLUmaWIS2WedR0a0PwvqkswXBjx9TjyiBOO2Ty1OyAtl0YoprK9C/nyY7faaaob
2uQvud0+0lZ2Mk/8hspP9Mo4ZeUtkZw/56xo7PSJKZ2rb6Zy5WV/HZFxflrI+mRh
Cd4vRfnlj62yyfo0z41MizhrCUMNJB2ki6zxkX3ueA02L+/Y/0c08T7Ur7QnsmAD
Nnag3avBezEUjN10O433ssgr2o0ZVJunf1iCIwgey/e+4xkhnd0LnjD+tqjWBMDE
34pW80LJPamcjZrWwX7+eUggLRQ4+hVBYvUdcEBo/Gg6NpvARk/sgfpas5wLpqWR
yDtnQ7975D5ih+IUjDIiQdpVhAN+zV3Tp6K2WY7kL9/JrxH3yXJ9+DKv4HTrm2N5
f7iwtC1jcdA685fxyGgUteIM5Y1Hfzqo8yfckCKnC3lAP6DacdOSWHbKSvlgd8vI
1CoaVxp7SudKO/ka8+nj9y18Iv+x7PuOAbcphBE/EtGmf3rlOJZakBBG9A0QPrte
EySX0KA8TlwAEwMO5fkvNiSyh1NRT1XnLMQuE5mszmGEU10uYxbgVUePT9a0KeNk
J++ymOIp8sYbU4BfxUz124MBlyEQY9cCfAflZUgZ3C3/9nGMGbl4L54SabiXEZpj
nGr1RKb7M89DqVAoaNB+F4aweeuR7LP5bMEaBIoLlBTOvDUbghByLYgt/THHEIbu
rEJww3qMgL24kgyY89Z72G0yLeZc+FSYvDaWyqqZnp3uiHITTVUImh70CcTQLoMm
nvKQ3UBDrB6sSpfJj4DK2qgrOgtupm9MLrV2K4dDRiru037vJJEuDkKaBuVBpuHb
NE2tzz3I3DN/c+/6arCoKXFiYg8qqklzDodCWsba0IbI69iSXhm3vUrUuUnB81vc
3gNWg4Cs3OEon4/+TnxhBeYmFHxLTnmRWNwoQOA2PPd+ZZFB8oh+ffrwxiTLpw1E
ULVl5p53n8im2zsNVBGQaGrTV6NSfbfhaYL+j6kDiu4oQuw2uqipKgbJNOn4v875
vCMe/B/9BaTKlM7xTTe+AZhGGEHZREgcgAn9KeHeksCn11jE9+SafV9xUXTBUvyY
XtqOnxeZX3mfCHdeLHBpN9fqgd8Cr6fpspdMq1nMnC/6KlExupxOUkkc5kuuerDh
ajluNPzlC7ISmQD7l+TNtds4++Z4IXFP3eqDfTngqbAJcSo9ks52gJ9Nopu9vvAL
H8c8Z/RqmJgx2jFwxmvOh6MxW2t6bmiSwbBpvFzcgDFvbRbAM4/vJgxCW7my/a0U
Gz85Tf4KafHQradrl/KNIe4I0cgZYNClvpxIF7yP1YZ5snXI50Uxo56Cs6b1ZV8I
Fb5Seb7GSQQtyk3xWKHPEHaz212xw0nE+c/REw8mX8YHguqVtoxMDUszvVbTKkAI
ABtx9PNoGozuhKjMA76Eiu9fE//ea1dSt9TxultPGOTQZpXUVyCdDNn0eHK+pLcx
N1rCVnexEgL+Rj7HI5p60hMhozhltx7dRO7YeJdH0hEB6jYFZ1bkNx19fn4VR8Ki
zebSLN4/EqpWn/w1Oznmr2bIeI21mOXO9yetMsSjU4B7RlnRbYqPXV1TuU5raftY
76dBbwO6M/Xfe2FMfvN1Fhuoys2V3WH6xLbCYwY6CCqdNgjle256JwpYWVVu9MFf
qUXGUyjKlFa/a/RhFbk9RSOc67o+UwKwGkGLwP+ZM0fZ5DNrSIvc69nrDhlwpa8X
IzeuUL7QQZHadUP0BoPTqNk6XAwZzFNMAfvMxh2Rb5Ca0cvw4TlfWEOqyMllRtyG
7WgCim2FiWGz86SxVTInYTL5vYJlJwhlA+GiqKu6TSYs0nDpCCqy15GP12PlxEHi
5stDHgXkIbZsQnPII5xm1pZB6ZmArWLCUD9I3tQyDRsoIK2CgMl8lzHdepM3ylpu
xOGINkAuskcUjTINZ7Top54kvy2nZMELaoMqI5ybIaFdsfYoW0xWg4h/CURDFfAl
H31uahjkxRnrACMTH1PsY9OeEBkVtmJ8SFwFIm1FsNj4lyUm16x9PE/OMRkiKKGP
CVmxRu4g23yMA3IKz7rLaaw9hoWUzvU0bT3H+A94iqlcNUVYylxgydBX58OIHOaN
ZWdSf/Oq5p5LUFm1nn1sw5j7gvJYt/4ohDAQGVsivkJhSdyVL+jwFIc/Ga5qubN9
5uZnoJNXzMTSo8sBqMzFVAfnqeLyBymAj+PX6kW+sf/yOSGaJDzqF8AZzZa1i03F
zentl0LhKreNqJMFvcPFw7c96v/wdc7UXiezuf2fJgPAjwuafvlIWicI662fSsjN
qNXAmAjbdfxkbFklvYeSfTTP8h4lMXe/yPr/kdxV8cj/5nvy99BKWrcENRxtSPps
6q2TqmZXFW1BJrahaRPZipWu7KfAhz3JUPGSXpgUKWhogGpAae+w5AMPk4Gz8srI
DiY4B/oyZRZFzKxMRFdxF5MXp2sCo9CtLl7zPoKy8zMmuPPbgLkO2pPemHOqs2ZA
ZuziOfQXblbUfO8SOSSsDegbLnX7SmAHW+rb3rjwxPvrNtepPgNZGX6jbY05gRlY
qdnpewcRMY2KHcUYl+6lFZX8jTU7SFxXq0EO0123Yajvun6sA5Mv5RuWAysVcQdD
ESPsFx3XpeAkwZ6x+LxhMdwtbvuXQG70VjVNhvEhF3zH0CuIsaz+bEqFXQsRoUv9
EapjZGGKvwy/7qTehW1MIK6U2nGO6jYHfkFAxbrrtNM5QODtfkieSAjHkf3U4HUK
B1haju/Cf6mVLhh+O5P2vqBwuFXkW4r/kimW8+EwHBNxwuWfuliSSFxewCDnRGbc
nHqGAj9wsW2qwVz+w/NMuSsfqZsGpjLCyvmi58xZOlfe4wJe41j+O/nUN5eInmmS
G5ZZTpLF5E9/edwHARXjhexJQwK/zGptRCigNcBgbX40PIaw4pbTBKaFhKKW99RY
+ztLaYWNdzT5m/uP6/f5B6Qe0tpXcnUqwJXGyjMrRafc8hY5cmKLJ10l5EXNUC1E
NB85oiT5pLxBpS3xNMyW23vrA0dHM/GqC6J9lmChms4PFZ6lCRUnFesUj/bxno4p
c3K1PSS6dJ7OSqasKL97U4IfYJqshMHeWE/Q/AVOVKqXvVmYLckGabwXFJs290p/
KcpfE/wSOjEHbDDCTSmIz2dUuislMWCEv5v5jjBMf/k11Pc9tVZpjgY4ZuxVVyDn
FuvxZhXvEfyfRbExwaJwZiCQIDhajoxrdzevM/sCOR73QA+/5k6RFtdj8k3lAtIp
enTgm6MSaZsNz+Ktuv36YlOrHxo3yXgq4N2uGNEgCOLC5whOsQiQLJl1IAlwOsBo
RjI5OIeTAFibujx0wtjNLI3KNvIALKlemp2Q+pDQJHmKARiSUG85s2m8cHZoyBq9
2FQA05W4zEh2XBsiK6B+PbCRkQdA6JtBqy545MyCjLCRyEV6yHpH1ZmRav/P+w6D
m1+mDcaSfzV7gm8TqvfTva/HFD/o377LiGrTTDmT1unP9ecqCJP4n0guUjOjWB2P
+OVBZZDAnfE2/U/x/LdOpaw6OarTiqjO4NSV1+VtyFXPoQ4s1xlfNrIvF96yjOJ6
99n3zNV1jtMtgcBzsstL2DQqoB5cP/JC3CUdU2GoLeeYaJRfM/2SqwTVIu/Q3x3q
yr2RRn6aWn+cyZIjuLPJFV47T1Ej/EPDoKEf46HSPlCTKzHuQILAmVchWmiPzcXu
t37JlI5035wdsA3o2Cq8Qo8SP378VEkalk4gXTPHhQvMFUkw2O5SnDsRmfz76lEn
wlTo0fBoU5pgHpkO57LmEwMFh/oM+/Rt4ZW1GI/lmhzpxmWMzNhB+ZkOf/a2nzb2
mlulJiJkpGB/1XxcQz6hh3829gAKGVTmQPNKPo8bfy8SXsFxQEuZ1o0izsaMNosN
kDtC1Bws84bFVr1e0oHWO49sWV3tJPqyZWy9hlhHSjSAClmTDKXXkJpn1cweaDHc
GuRwLMwwTzs0ldes/QjUVhsNz1VJmG/0KBNVZorChlwJ2qa/5VHGL0dYhlEF0cvr
0RXb3gR7nWdj51mv6/v3BJMAaLAxHfwVvspiGcTP2hPdH2s/HYTMFZmZDcUIhEhB
gijuR80ATlE8o1swEjeKstLQKqDGQfmoPaEhLCs5g+XOsdT2rudH+stdCXVCJnDK
XH3wUT8xIG6hP7GuOgIC38CGNSSSy+PQvUZ5OjLYWw4+vp2zjZWk9kPYUJCqXGjS
XkA1j6IK5af9ytHWU//3I4k76FQQp4yAfjGaTmU+Xbc8dXC24CfFVw6iEqUHWZyX
PMolvbwp+oz4bLaDw0iB5u/n5rdQyVfDkJpxHVea2KpLpRHGJ+SsyptyBWzyf9xf
2/PXQ2X8EuQygbtzuS8pKhpTJ/qqPgKg9A4Z/sNDVFd4mk0WMXnq3cWDeiFKSNOE
rITkGEvwddNDoAyoJ85dXQ/OWiIESwV9JsB+oun1d7e2R7yPnZUcubvQrJkDDtlx
KhYrgM7xV363tZ8BeB4cJFpovscLL6H1xNWxJaYrz9gihDa69gT70xbf9vOl2xKc
8akozuGMFt975Acl9FCVHd+RjswabStW1/FgXVhKchM+je6wEF+cZUttT1T8EPBC
qZwth4BNOaYeEXSbmtljffwyZnJarSmsYMyeX60FOTMb9uhb3di19Y//RJ5rfq20
zRK24f4TB2LTVUIngzgiJji6GpbYjl+kPiHBTdaRmLqm09V9Cqb1MkAH/t24Z0en
1K0IROSdy+N0KjjA61WzKvaeE40rm6ViLq2HLuxQKF4+bDuYDSvY1UPRGyQ5RxOF
4aCPcfXyHkVWirYOl6LK0Re6BddV/1GSL3Pj8YrmVekskrPrmrPASthsOUoy2cM7
i/8NU23+3yVyj30zkebEhNeeeL/fjlVKQUPE+3sKRT34WIAM9tN3A7B1Bj3lE0aA
MIpYPCeBvG+zQIpwmvCGYN1zkNkVY/tSoRRJf7iud6ncfZcWR9QtEF5kTttqntQR
GsxCXN9TYTI4lnS01fHnI8LgiHmyse9nneGS0cxYrW7xqSgMiEAmLbcCa4Ftb64v
h+q/PTC/BCWTuU112RKmiP+tPs/OQV2sgEJRaVUjhkw7oc+3UdnC7GrGDkrb1xG1
ecMzTYzvN+zf1hZHHtPbudQqAA0ABB5NMkTfpy/z+l0f19xxEfuUUOoOyCfEVbJG
TfQ7JkwAK4NeIxCCz/iGZ5yxAuP6AyjjiX6hLxP3bOUguD7i9EsCnoerW5GLMsJT
rJujzk4QVq8hFwq/FhO0s1hNBCIytUoFsUZo//m//T4b4yunYr9MPpoSb4ugiqGK
maWpGnweRMGkpjANuzTY8vLuHsnbaIiRXlMGctow2z2gLpFl2AtjM08zwmiXOqol
ef4+Qg2404UBzutkA5kPXODTX15ys7+dC4JYDP0uPtZ++2H/uQe1YtqumyD/hfcr
kQY/ag7qmRqfjLrfdWSAQOV3Rgo406FWzCyPDVTD0PzcpG2vPD9KFJNbjC2bDse6
rmndDQ2eLhbUtiI2HvAS5/dBSJ/JHxRL2lfLVpiWcfhatfEuGluLwWiEUosc4Gpg
8tUBYc2LF6hnY35NGDEbuGltSf7xR3nLqn2kraM9oGLU4ECC4AtWHZNwx5yHpsc6
uiTgJWJM460wSe3G/bvRvyZB2J8FXbATt/ZxZGKHWTd2Hf5r15yyoRy616lGc2tX
QAtkg/+tiXcf53to9vHD/JdLi5N8a6GQkXb0AG3Q4t8ShzWtEyAVTHrfjo+iw7a7
fIozTXU2t0dlCsDkDpIWh0yZ/+a2NqcCCr7VpsIDw2CUfrp0QA9MlLzl68rxA0of
Y5IKuMfQxmxYK7stdkhHW8kKB/gBClK6x3V2HHKIwFNkyVPxw7fJxY3FgnaceDFn
+5NBImiX33T7L41FPlkSKTKj8oOGEuZoSS+7RWNJYrwvqMGK2TIqarcrAoyZ0zcN
ES3zNkFdsAO8ounjQLZCC1KRXaxw6uTfrZ3Aa4gX66STMN5bDIqPTJjoqQceLPHv
Ulwb39bYsgXsUEtfuSE/qI04LQ/lyoUw+31IXrxmXKAlENKhULG9GollIO+GxfMJ
0bVdoTPnYgTWItziIZeMwIU1XrooH/M3TdlInd51gC4KRZDIEygfWpJA8xYx+3Td
jZ0NnwlCBgkA8NiQj95Rj6+dfx4mC7TxYyOpNcWOJeJxMWJmmZgcqyvOWsQqlfNu
CENQherHyxNkdjw1MaJ5/1mROQ+98djBip3/acftnWdzW75QeIi/8iSD2xaS+2/y
kHOd89Voksf/wDAknf28ARs/ELKp/zGnNbkwcw/txI06fwIDbZSIQEUtYoAIU5Ii
YiQBaBxDMEBbx/moVccv/tmKvIzk81DLfE+Ru3nETS5kFj9nY71MvuFGy1UWCMpK
KJ4ebw2kLZTLkcjrDKnXBe3UDvilxVzmI91BbA8kIwKVlu9wiMg7wfzvizBHxGiC
9yJc2Nfp7tocsJAJE3HHs09j1WOu7Gb65a8JLwpk1dUJLoPS9iwATVIWaYS5IVli
VW8oEDaZ9mTtBLKo4YkvPKvgzhx4d7PYoJOCEa4hIoPybAW2pO6cfOIDPqVP2CxA
4dYbWesp6YBFwiCo3Q/1fStk9haFBjB8uXh4gtnOfwYD8YPWQEou6mKleuhGqzOt
1aQi/nv7xAM+1f2ny7qDJA2YHLCoQak3fgyjroHnUCof+rTxCPfYkREU2QBWEzm8
mxlxzYlp7Uvhw77/8v4XywJnNDVVBdkMdW01hYK3NCRxim50nSsBLs5QY6jlfY+Q
ZO/2taV+lLlCQbaLp+GZfN9QC7lp1+O2xTdID/+tJTV6ftW1xTJDiWJGmInwKnvl
nidnhdktfp1K08TJIFbivjSIDiHH9kXxmoyNl4zDDu9Yu5sivoUYlo3oz1BG6HIl
fEeHCOQ0TV6ZoU2E6I+dAT5EzT8SzmloG4qpPuQ9a4or/aGrxNSXKRLZVYRQZ7gO
W5zLjBT4m9Brb5tZBbqzwocp78sg/eJCiJzH0DdlpQIi8eGUFfj+Syjk85EzO1PN
3p3ceVrjbYiI+83xWq34O4/7J/HgcqZRcX3kLgWQufWNhrwi8gdr7ERGlGfmvSWC
8PcQ/oVKgiVTTE5b26y+Q8BYK4Q0FitXUhKwqVBelg2kTfw+aeg5VWprUaaTtYOx
b4b/j4MBLaYKkLaRy2VdRPyGUhyecII7ZGkqnMDFnLBo69k/Wd7vbocRQIKamVFl
hPBzV9AiZMejdjv5RbzH/U0W+x9G7es07C3/jrKxVvNK36ThgqZ0+yg1pqyU7od4
XQ4auXKqT032ViGyQVg75Uw2I6nskfelvREyYaLUEpZD5e1LjGYdqI5tJFwAl7rM
GHIEaOhTK2ocZEKlA83tZWCTR2pRcjvZHn7TmCxUVaqXZXLqf0lF1wEQnsAZuEWy
U3dWQLGVuzOd3oFcipCSo20QLg3YP1H/NwWh4hygeY9+6iqraIpqVcbJEAyMIcir
ZUrxvY/9dirnmsdee3dSvzdYpDeXVb7Q9oMxQ7K7+yBWfddbeEM5Y/6pxF2K78a0
m1H2BPwCBG73Mavms84jv5lZ94JwhzdGCehmkcqg1A+ujlL9Ta/RBh8c4ZgfXsvf
kq4F6e2hBkOZX87YuufLyO9TZErrmeVnkSU3eMQRZlX3al7UuH2/6tIZleHlcQtM
lZnlLf9Nt03et1CNwVqRLpYg/9nMDv/li9777U4aUL21+gHQI+4VD2kvhfICyE+9
1fszRCnGOXJd4dPZ0GJdOxiN5nPm9K8EKVXzYgx8M6Hyu6okFmo/llK2P4VnY7E5
w+LbaovlK14Vn0XQ/gm55MNziy8BVEM0Kl8ZEhXs9auf94V6r3ojrk4qsQRbcIFv
yTQ0NvvJujmXWNAGJe0Zl3kgc4PkInrZDh6LgxHjVXgOicPo+znYsyUwiU4ZMMRn
GSLalZ76gz0zZGuzZUA5HBdoWor7TjXzcm/5vlUTUAyNuYvis+JYPinIqYjMw3Al
PPDxcrNlMryyU5kBxiQ/ZE5hG8kE37OwTRd5UZ5O+JQ+x03AffVT31P+nOb8dFWk
CmtPfHL0cpIUICg7nDwvFTwOsisJATNa9LcWKVFfHy/KLhslDAtjy0uw2KPJM+VO
jd+oxcTzDwcs8j53AnOA5iIsDwrGYlJ342aX8A+z1WHuj9Z6lZdY0l5WPpJ9Za1o
jmRoC/XMVRvq6fpEjaO9zOErQMxWrO3+ZQAd+ZL4Q0TnFaJqUYRs1oeApJ3H1Q/P
U6M1hWKJWdHIaqsR+BG363tt28ia2qq84gM6v3qKXhAQGjHC5+dMtXYeaWtLUtSX
QIGn6hnXpeEDf8Lkb20RnkHJS2FdanY8G3FUHxuBxBeRSaVsPTJo7JoMJdepeSnL
uI3iPineI/89fRgWpTwwkiQHx+S1USfWE0EB+4gkAMvnLkretonNK5MFLea4OAb7
g5oWAyRFfH3SetghjAjVvuy9rg56UJh0VbfjBQpk7wuH4V8ODokdMwiC7SISl01F
vYHxW05xfMmvjLC7Ja+kxLM3PP0shZ0MtATyeJTNQPtF/HwKnznSfKWm46opZvxf
/wvjGMTDgxi6VN+KALOHVw/iifoP/8nhwj3SPYYk7vKY0iT5DNCZfMX3SKXeZJPL
K29Vxz4LBroD2UUtZK41EChsItyYtLwuSPATgHmnqG2zvNT+FkdI2wl92MWfu9A8
aRsngxgcEDitCiewJ/XsGt8AagLlTm2T4d6dVzx8xu/w7DDq3uGcY/o4Dd4I8vqr
DpJeeVqMk5EtOEitFWtpIe5qNW76sPBiBIE1BuplxiCX1sfHo5o475ZxC3+pGM5z
WMP3JYN6lgOKKm7C+eYPI6bhvfdb/CU44n+sYZ+MrQh+eETpRa4jeL3imWFF84yO
K7lURZmeCB7X9PTt9PjGICzTuz3rcLLltwv/OV/K76v0Y6zdJm4iX4oRILd1PKZR
Y7dT177eyyOovYnpzTiSyV5lic771l9EKqrTQMclFBWHcZ1/eAYCW+fQ6H/zTks9
WsShWgBJdYdLGH7fnV1/FZTWFVK+LW2sDPOzpLEc8aQf63dSYy7eP5eAa6Hx7KvY
xLsBWPV86qKXEp5eZU6Fp418IkOov/TJ3w2rpHD/LkcYwm1qiS5UoVPDTkEXKVbe
m2qXVm3gBy8W1zZ2WUXMrVftCbIK4CddIiJ/80MZLQpd/+emN5cjIi1Oi50FW4Hj
WvRS7oQPGvCNYSxmvdGTkjIQJLSB6R63eCcTfuEAYG1qMCPaOZXWeqd/bQNqKuVG
0EdAh272dDP9FPsHEOeLfcNlZPa9npBOYz1Eqfy04SvWR+gtAgQcELL40bSzpjGO
28+zmeYKX8R8ckfrSvHxAnWfVlvAqqMl4kqYljbtNG5MgSBS0zk1qEyCdE7h9BOL
DnH8OZnrlGDinCFb5FhfXJIlw4JwFi+/DLXkT3TLtYC3ETgkfyVAIQjBeuDd4zqM
2pDiEPiPlrfwDfvsKKYrnRsC8c+tEz2v4hv8jU92AmOZKamyNXlbWydqq/GRhOI0
JD4vt5gmA1i1uL7g6MFq0MVyABPyrjoioNgCPmGYV0Tljn1g/xZRu6SdWYhu9aYo
NcPG+5QzOPowFZTHb0jKVqI4hPFImFynFXPpBYm5GB+rJXTx0rdFBEKCkBQY8bJL
+1W1BHIId4VyvEKUaQ05dSdR4q8elrIn6bD1a0eR+uEm9ZRQ4K3Dpm9DwzL5+yQA
QF5U0n/8NrI7H6/XuqK66WwvhfAQjOCXknbg7A/H6fyzo100NHeL3B2Ah9M8Tj8K
ebCAv0ou9Ehe10JL/NF++Qfj5sXKXEmBaqJ/Gmo9MUnDq0MBZOh6LI0zsK+Lm1aV
EaGg0lUYlwtKVkm+y7CW0yGESzduSd+GScOAgsiNRDC+ZvR7CryxAMC32zSvFlkH
A/e5GOiIvCWV8hQI86pIdsZzLZx/2YlmRX+Ya12KBAWfJP+UcezUTQGAqSIr41Io
6I8XYZjZ/ZkFNUDcG1MiPKJoKshmMVrinonaJWxQrgV/AItEZA2M4BT7pSrXID0i
KLCT0q/TjlxkvOhygEHjvLbeNb0zkmy22/Zn0ScXM4sjhu16rLIQJfkk5xUY6fe0
cshoxQgr2EpBo49MEhTcfI9N2RYiG/SYuuPJv3BV4kriEpDiMbBcIik+KiP1FgZk
WpDg9J/ibJLHXnhcuBrjYP90br1GSuLyRidZRovGJETS12ZzM9GykNvGfBsDndY7
ZGFhIeq5tOULKwiCaWmCO5yDiz8+iC0yvN2gISHvX29PvudVjTr4MdVDIPME3Y6c
LhTroRsB/qhFFKR1AyX+pnVPxvEriBOk5ZTfb/WTQICZma2Ljc3Wv4mrzP04crFk
LKoLreEo73qvFzpyJxUxo2iiYChHx8LoJBPcsuek8QCpnIsFQjDRHAE7yuETEZRc
kaG9X2aRW9OW01UCZb/DG6iDTcAVZ2k7mZVvJwJeYhQmIADNd7LhM1EY0ASfR3nK
y6UIHj+FI28mdsZmXnNd8umZ1K/C5BnrMTvo6hnOzW7UfVAomDWPrjTdXFma8OBp
fBRFhyG8gcrScE8uVbXm4YLzcI6YsWpnXkpXu/u+CIJPYgs88iCZb36D6X9CEr/3
d1HuUZ6SDoz5u/8keeartLqoFyf4/Gm1y3AlO2LAX+tb/ztHLJ99IgOxpKqvBlK5
gadiguoLD+/wuj+Y3iCwluPKCGbnSv9UP4HaLp0Mb/foupISC3JdM6wFQhXmkUba
YJvGdmxXZWjqtP1aSfyIGGMXhflXNpXUj2oQA4x7jy8/DM67EuZD4r96vVAngAKr
q9k6g/xTpPgjt744lGwoBT3AFPa4dwL58Ws2n0J6vQduUqkAo0xYwP5TxKynClLc
G+vcRAxbe2X7QEiUc2bTHJCpQYQpOPKdxBeXNS/ur7nshG7mwqeP6qi4MTzaqPXv
1SC0qXp4nERXhf/QY6/r/RBvBYNubcgXcgUUOrYaHE5ZBFQJkuolGpen9ZVGbteY
pCNr0oj7qCUPoSurHs3H+KB/HFFcvC+O7W+ALhWmF+G3D9zM8pLdRyGQ2ov/RxW+
uTxL2Ow3b0/dsebgEHEQ2bKZ4JD3PkRO1086rIwWYEkst8M1DK0iZda4L6GpMNk2
z39Ab7pl9EyeridYNxsdlu/+x/mDutL2ge4S+msIGRTYV+M1kH4fFz4QUDtj3Om2
3OdV/Go5gImMPoqfuFrg3tJkNbK++Q8v2CFx/UcBCepAiw6iMjOFqU1xWNKOVDpL
CoXp5MxEckdXnQ4HpadhdkCYoKhdMjuNzUNKkt7vkxE19gkAUijeRlIH/UNFVXqr
fMyRwhbZ2Cq8jmvM6+kLiSXnp1ZVNiWoP4m+0q3MTzKqxsj00qsQVmZh/nUiMY4m
QxhcHG85bC7ZKDL4uTnPVx7VM8lKsauo+NEe3DKoNLZRqZvVapw43kly670DMckb
Qfbz6LD9k7r3zMNYepkqJ6P7Ssv/FooeTVAdxilVy/7gQ2o+FxLGbGTTTDgTGrSg
ZzytNMTI3Zfn18Mn55POXKeuc8XwRw/X1mvBkdPgNFo917YwnWcT/Q3kn6YaTL2J
+REeTIzLMAhmKkpMAuWUPZUeT07WsbvK7s5xoQE2p8lnSG7hFOXp4Dt73RpkWbzp
9hDg8Ke7+5HkeWdDOc23dfY11jC0gW8M0etY7+Bb19UOeDgoPpfczcpj9ioLH2jj
LENqMcBKaln10RfsonYL2dmY69hP/DCQg+FijJR6AADUNhWgXpVVveeHsLz6R1bu
vq6MNiEEGovEWZIoCrmsEshHBm/LLgBC8VwUIxz5E29ekOnHvhrWXVSsyVVe7oD8
GioYmTgQWmGbVwh8cBI7S7QbAJpwZBGkD/WEidcVlFrrvh5fIBXhZN98bUn5Vg7D
gI/SVGdoKZROQakbYTUcfuD/LnOi8wOmIvk3qDycCQfXjuOrFVa5U6Rs8i0s35zM
4fNeFI5PibumMDZbcl/9cKAWQkmvsKVE3GWkT+o3wTcf4ZmJfoVxNA7KhTuPmzVZ
07orECkkTZzX373c3rBkv0sHB5g1sIRXxTE9fDXfWqmYLnaekdO7xvPVL9cXXj4/
gcEF6Fqm4UQuUzeFXW6n26ZREt5R49sfr5aLA6xCYTrjFsiLHYqbEtzLM1ZrRzjD
wF5JpCFJ9NmtprHbXl3cy8FB89JUxxzYwliEsZ+6WONBM18wVuHe/2IMFFXFGtmn
kCo4P4DKThDtMQeNiHvqOnN6nj4q4fc8H6Ttz40SYA/Z169801+dw9E3vZS6Le7V
I6qJP4INPoYvG7uhg9woS5cvDRrkCOa6+wHDN0kXFNdkuX5LcHi60snXwWAW7uXs
bzfJ3t5rCzjxSrrz+bkSCR9vWhkKbNFPvbaY6lcpjMBxgFqMUR5qWqvJyNPdPL6+
k3RIRwei99IP4EVf1sITifpa5NUfuZAWmSPuNvWc9B4xpFD4x77jQIKs1u6+oeYL
pl2GwYXXBtalChVVZpLRtx0xbgMx0/tf2SajCCvLxR9zBDCQwzbBZ6GnFk4b3p+m
TDYIqVXDtOiHxu/1WFiGJzJavNZ7uwDye3DUwBXU5Pl4eRSUVH9lNvTtEN3LrvPy
Jp6ZryisnZ1pjt7ixKhJuYK8myl/pHX6JDJM135D8hhb14lEAteG/PhHSJYw27kf
cJBdbeXAtEH/SeZN3qQ0eJmsw6diIDYVZP8ZhoPgMxTPNlEmIv14mXi7IyR+mBYk
faD6ecqR7FzrRxyx5E+tlc9fDUp7GIuUMRTJsj0+L9fKgeRi1BUlAxlIcuz2MYRM
LXlMJnaGqhRiuWQpEp2z+t1+qejYtEW2e3tgt0HpyfOV0dxbE/dNv3GY1PlfHCr6
NB7bTvG5dnG7q62oT/cr7HZUnJ9lKNpzpRxTGT8jbo+pOTfYEPZcR6T6mmjGjfd4
IQg72ac2MWjoOP0Kv++NKqqB3a0Dj6E4SduFQrNUkfvVNLH+KwMB6Vff9eizWI0C
tSynyOsCvxE5uIJn/SKldyoXOLQgA2iOWlCwwln0Yj5AKR7K2dFDOBD/P2fmA1iJ
C5ChtGzO+tX7BVgLYOfIZGcJ5lg91Yp9gbciYjPaTJZoWSoWPc5pz1E3KEDySlek
C/Hg92hWuLWCDHOwtoGT7AtpVbbpDUInvxvbUH5gGl92ywulnNqY7P4VZ8NXF3xx
X8k91Q8ULDnXOD6E3fBzlsyZlPm72+op6aGrbW4PtrEYw0Puam+0HDGFKbnl2zYA
pt2x8r0z8B/PQ89OEMzLooDgC3gYaibmwlpuAjdjnfWFrDNQwJu/SIp+dI9UEze7
KVYg/TI9PjuaiEROJvtirY010+0SiKEB89TDHDblmRrqqAuBslLuzXCQi1RYXKcq
akGFME2CO9rDP3cvnjmnV0eYj1Kdv6j7xZwodbklmJicJtt6Jos9fSqH9CWdRZPY
KQyuN1tSWE4JvpFldGJYlQozaMrXfJxSSNSnkZzQZQEhUla8uvnTh4yZhtYCYZXF
9YEL0oZIrQNDBqdYfiah3iWEYZFKt4fhbl6T1nF8KW21dezyWjtQ20vHzIenj0J5
/o1mO9nRUykyIb57LXpWJktVTl3XLgNRPK+bCYbkIHMkPcwwe0mldgwhqY2ylXx3
6suGUxE9aqY9W6AWXHWkraUISAwi9vmkDPNsWYrSrTxEX/cVcgeHgHsSFy2SLNel
EGTvp0dH1rf/z3zo6skIInrLsthC5JCQ8gaxfE/ccyckQVyg2aN/niXTEOps1Dij
nw+emryoR8tc/BZbAJRwxLqNyyJQxfMfjp6j6eZONqxC/BJiw1VAOmxqqPzr1ygk
f89yYr+gnAdopfdLlF0H2vFIF4Lf861oB9Em9keU1KzRpXpBiOi97AaPnkSUC3so
0HQLXxzLWpLo9O1aXgbovnSPiOinowZ4FoD4xmU1j8AgDrSyB0Y6wgS71sW2g0V8
Op/zy/EzcGu3d+J3bKEJzAALMcGzwAEjW5QkKwR3sNJ6xF5g9kDixT1iOzWjr0bN
HBr8RGHi1P0rEmb3mxwO93cSgMv13g3SElj64K83Kvn/nZQZYqh/G9PhJuwGQ6bj
DdREdWu8GcvMmEXHHi3KT0o8Ky9whI/0P1MBkdxLrmDLqzf8ezUgaKO6NmtQ/69u
f3MbrjGjs6pUnqIt9uzldd693NifoeDureSPtoEFKvccMP2BY1zBw3zwrT3F9FQA
qpxsWnvDCQ62a1MKQepLnL0++Sw5wZ0OUoVyHSrVOAFChLe4UwmpwwnVY+37h7jV
grVV/DNB8Rc0F/+JPb2c/HV3lk5bXMJhaWLFt+eiZUr6pyRqAr8N7kf5gDzNwUeV
txtZT+k77S1M1uc+VZ5ycIJou7LQ3p6e3i707EZaPG6bInbLND0M7MktYgGLGAiS
vw/j2lUDUPScbWHWXrnq9LP+rRzJ61f9RSr7YKSVYDQ/eBp03gQmHjzl1vLQI0wE
EU5NZ7Ns23Uhjop1WkjUAitpQiBkPv/iBdGuIWzJFJD7CkanbYf2HcnG4+400HT6
0inMlfUs234+RofRaynhDwgQBiEWS2K2QuDnK23UNQCcbbt2sxQzyUHi+EMFvpry
mN+0e6xkBU7IgvZmi2XY3t+Cj5DnwCvoQTHbnvXal19o0KTfQB2SONGtCTmGuzOl
OpsCN9ZDqNgRibhTLnU1X34SA4fjKPzeCHelWalDnJO9VTEYg5Zg0JVnAmVPDt1j
kTf2QnQ5NFe/ruaLLtrtSuYbqPzFOioT7QIXZcJ9igKIKPTIKPN5+LIj1LKfrjUn
YptEitpAOuTm66q34vIBnw0+4hO5D5ewL3cEFZYSpZPNeULM6BzPTkThEV+54z69
f1yRrUE0YP4Au97+ICPP2374ASSq1XGHYPFzERKhVnb5X+oCMXzh7auFg8Wp+Xjb
HA8aza2OugmIKOJChDLvSCH+icuUlsGOuOapyTpV0azDs5UmJjaWbKpK1q9FS4AM
pFanYrbmuA0E7f9JrhtUB5KK6AAKw4ZSK+swEN9HLnfk2expc5S7qnFSrVOhZtEf
Cm95H7+3Ta1WJXwxXzAuwDOhQu5Vfhp9ztAHevJ5eBb9QBQVPOM6EeKUDN366k6U
yVx4Xy5zLd9RAmKSIYaCaSwQM3iipEHxpD51XyDhvtnhPCN7Kj/C/BnL2jrSvaDj
u8iCwN7yFQHlSPn2C5c+CntfZupsHwjeo/jEB0NkTEshXN7d8943vBU7OPierslk
yS11MP3/uWYEIQo0OvnAgz25VC6L7ipVUxJJcazMOLqnL0n0dO0dk9SWYYSH0jWR
pXyOJdXR68tzuIjhVDFe+aQp/0abMGpH8b0owRaKAPx0nqkhwLdJtVgmCX7Xhku+
OUra/98XTNV8t9uJ9kdbMboWtlTkhCGvy0Rt8BuoEZcXubJc2kOEqkl0HaOqcNA8
mfZWbAOpmvmR2Gv0qDwLVlqif41V0NzYm+qQJ3hBKx4iOjqsKlXFhFLtKCO4qFXc
PQ3laP/8MiOq0/1P47pGwL+7EmmE5944Fcg9NJCATW0G0aK/1k2Frb2rG4N2KIs/
Luhharo37RYzL6NpV/wrA72JE/NLA1vt5sVHFkodLuKcUdhnA1UkDUm1hz9nJF5u
O/9PEWvv7oIbR5PNn5R842TkPRzcDDj4pIWAr9l7vxR/9BEbMsWh0mAVwJrIZe6a
2q8uwzK3LOFl72KG3doggZepkQ0OEFY1ztjLy6f86mveyJDXSQO0hSsq43/Hea1O
58HzyIL/6nxdfN8vyrdYVlmVoS33HP8d+VyFPXZnCV+EeBLJDVZdOeeP8KzcKR6v
qxpLCiIuLigXR5f18Bc+QAruFX2cZb65ZXNrB3/eKxQvqfugQVqVHC69VcJRIzJA
pdRJXQrK2lA0+tM1+ybSEGMOX11CyPbmQPWQ4DFgq9YZnlkMdKmNK7o2Qd+VBi1W
MGO4nSpm5oAYjchqvsjAlRKXGDPCc//C8u49ZOMXYXQH0P0WGj4iiZJVFGLTlArc
O6Oxev3b+KcYLzxPKT8Who6bPdF41Z/FiI7UZxj67JT1xYI6AGoN2YVCeU0dVPQj
WtAEmjmglCc8AAbn8l0wYxAusrfG8JPkuARac+Jn+3KlcbiAGanocIB+4XCv6SNh
dCR2u/rr+2/eh6URmWf1PSaR6fL9GJPMfBGyMc8mOmGStrUaEjwz1C8psGTAZmUr
+hMkeCL9uQsF6DuDiSNY+o9aMo9J5kFXsYxftVNHxNsVdPswz+Dr4g4s5X4KBSZH
XtAoL2/zsOtGeZm6as0nC9LdJujPKdDhrny++YzCTOqOU2ciOrwERPlEZ+NEDhYl
F+eEtHw1jcRfJKfMMomNJungOfCMsBtHFiA/IRIjohwGRWKRY51Mq6Noos+ORuCu
P+Z8XqZvxZpe+y6F/xA0mRPEV7oY/7Lub7gWLkCxHxPWdXrXC9PpRVI7ubLNoIA/
bl16ErZgr50eOXSp0ZQovfd8IDqKdRWWIo7+9NSj1S3tCsrm/maJ6q5JPtX7bXOT
Bnso6H/waN5FeU8ljd6t+Y/cHxPwAFb8SOLPeTvYkzmVYNF4RnvZjvRme6kChsaD
8nBaY9Lhhej/dKrJdS2GbXWNgsrx+iTYkXIVRvkUx482PjK9K1kX6Cu+FLse8IHV
IKW+qftx5APb3pR3XVUeBhrAk3jr9BaFtxQnjRiQCNa3JDia7DwAaU0rQumx/Gcm
YlX3rs7zYz33zkuhxEVrkyF1eMyvAoiSa7CaEifvVSXOvKdcSTVaSD4AD2nYnhRE
mRmrBzEuIOz5BBvCwlSgTnyaseyO99PMWhNnJSiGW66/PtyE+zjdKxC/SCpuij1O
Z/MHvWTiRpXm3J59G2rpSO/Btnv1Hm3Nzwbk9TrguKpz3zrJFTNK7U0JC77/PIKQ
vpdHdUDWJuvyGnq7iqYgGddUvkV6AenYU63I9an1VaSKFG5+8HZRu9eQuAVBc5gu
Z3psWaCS++tEkNi+aBTi52BDcdPNwUGOb++SwYlpZykhbhjn+oiYPdv4vwZaO+Xc
r28qV1vrNRBL8OS5z3oBBm4CIr5DmoKnyN3h9vt/qEsKghiwCHzd/jn5mMj7LXi5
YQFrDS/fi1Dy1jpJ1IlE+4C90vtx0d9ZXfAVDiYl5G1WP1THZDGLmsqgLoSp5EEw
1qM/9PWxXXMPeQ+7UnJedAoCQKAHmo8GaaR4fMS1lqrxe4NuzbcB3KVH/XzprRhX
Qr+EHn+Vc2Js+tMsXbdZU/uM2jNtPGB6rNPYqYugtQcUgDG5QO3vQydnE7u7lyOW
xwmelKarwF23JP0rbj6fSh0d2gR6atqDV5Fj5jPPwbVQuOQLUiwwa1b/61EPH8Bu
YYV3J/sHP/HI54HqiWfi+CRjh9pKGhnfA4x0JNjjaQNw+h1sTtbFeOxCnKRZ8O6x
bcd9Uml48aKv1YBIBpAk8RHhneiX8Mw4qJKl+wSyYeGPXbGWwKGkIFK/m+5DiS2g
CZPl6AT1Xi02j+KH4jqipa3DfVN25D84IFvlGrB9g6Hhb/2QG/J4hPffVm8Zmanm
t/7byg8/3lsNCwlmVQYKXEX4VLygw5Mw9XmdegWDWv63UqZG4MG+kkKT+bm3lj12
OtB5eUsmBD4BRQSX0ZYjUBVNUkVVQmG19VCNSotTrz8GnO+BBEZmzmcNdADhqvLI
MzCCv5w2PXJF7oNzjdj0oGkFqE8LLeU9SpPM2T8m3Of5L1ObP7g4llfg1XBzEYFu
912x+pn3U2kghRRl+fgcikUAq2iuZXKeSFB8Gd5QyRRJjWSvqIczOuBbC054ONYw
asNVv1RziUnXb6PDtu5UXdxbAhULWWVi/+Hk71ww092qiJrxgrFSzk2ythDRh4+i
mkqeCj845bcLS/rh3kxdmJVlSF2aag5g3Jt0quYQ/aoCx1nbc6f2/XxFcepuxZjz
dLD2/xakAY9bChS9qMZ02rDBwZoaIfC29xa6YlbrlpQnPshPOoebTBJAONUMcazQ
wApK2Fr3SKywd9P2V2/twXsitHSULSq+Xt39v0iDH5lgowAODxAjI29mbLvv/BeW
SdKch2rV4q+UbJAWDlfOWMM7Awd4zO+0hhcGBntP0MDItvnbw0VmQSW6hY/8l3zL
UWYbz3TSU3CMFS/ec7pPXS4TSVDeu+G4TkpY9aL5/jFT/bqyliYx5t1N+dmWbQiR
rHc9B99eM/NXa1KAYF7317QLX5JjQyJ4sd4bucesiG2mLDUao/QsKDvqT2G2zSNF
xrz8eD5vkxBqwdHJQB72KgC5A9cQ8y6E3kl1f7lqtVXcO+9OSdIMhMex9LTPlY5+
7D+i3+YvOrmXM1/6g+qR1+FP9CvS6i2U/yTF1EhGRS9aR8pyPyGWCpw5ITwp98Fb
ZWdUu1nkPgE4GnWhKRyv5VzKE4l9MR5bE31yfGTa1Br6ZRJySwBvhH2NOi8RTc4O
N15d2NpTcKnLVaXMWe5fDNN3yPAewnEq/0YjK2Tq9ZV8m4pw/ycw2nYNKiW5AZSE
MNrcc+PnGCyulbkEC6QoZZ9TmSPsk0MUX0xm76Dwa6nsc33hjnoiZtVELVzsSp6F
Qc8al5nQfcozAZgUDLT1cmNe0uNKPo8+f5VHEZAvLAz0buxtwhoIDbvzOihDERiN
SdsrPgEjVjdv0nWWVJXFn4Qco5tJGTH7W0T/lNv/ZynIGx23uC8B42fvE4PC6wLp
EPZBMuX8Fk8FEpAlIEFp1xHrsdiIRlSIuyx1hmcepzcJJyUKjIY0h70aCTe26jtg
fLDyUPWEe+ztShgAkBa44ivMfyY3KwjbhRU422zDVM4OZGxMD1/QS0jdpv9RkR7O
4PBCeaE8w6bowA5rH1Jfw74PkpsuQJVryE3o5oIjwnhRyBMN41f9juWkrEBBFThB
PhXrF0Obkgr0uwjKuRKnuP/gM9JIM3eSV/8mJ7h5115Hzp00fIu2/W2Nvgeo+xyJ
lLAPJKcDVOMcxgxzIPo2ifMaC4qcfTeNg5AhKdQaKW+cWsb2/9NSU9NwiPsYj3xm
8rJclZmbxU+0UVVpeBWIbVVSZz1GaJ/UQriRyrK717N0gXOYUVBcPzQdyBgHsjEt
/WAS+1KTRPRr7+KNaheW3qMs/rLdo7nFqsWFaGoJOQGYvr3tNZWL5zomgKzo48Ul
OiHk122UUfpDPCY0H+IssfuOH6KBuinwt1EvEHhNjAfHUBwboyXWDSAXFPIE6/iT
5Ap0RbONzDm4NmcrzqtSggzO8dJB8tjVyfZndI1rnxrA1NhWZabJ2wzLBTDH+lzs
Cqboh79NxIOzXFaHAchuSCeSuRXeYoqymbIWZnMypIVONUT/tlg/x4/xjXEYdWHI
1waRrqTO0wHaL+850fenyBnawuvsuG1bvpAkVEDyxciSfmGgVRg7xcyTnXdOXGs/
i6w+tYTjPm3gPBGanVaJyA8U7VOdNuKZhOPiJcry2cx3dv9KTr+L8TxZfoyUZO+q
REftxb9ED8cjGrLFEDzjhSJkRUs1uTJnAVHgxsEprapg9pDtZAnKBZGKR2FF4/mR
IcjeGvlWKIcwZHO+ZmQ0sySTXd1H0eYQNaypvQJASeqbnESFESsrULYbJV0TAuof
FFoWlvjBqr+oL23JBzxps+8IdUQ47WNinWWMFXy7PQQimONHxRvvPTple0Rz7b3/
PwuVn99kxo8iDWlw/PSQ4RDC9njvnzOnj9gjASGfoyjWWCdXzx5+HzssmofKeyxd
Cz0BCuyJM4W2LX4OwM1/Nrwn/YIAmxDXFQXe2ikPDoNshBtZW/Mvy69NQzr8TyA+
rxiTqZakzEzzKy2CGRP3ElK5wvvPDi2WheMqC683HLqTDdpNUozjVVPbJKiePyga
tfHwBTUTugCbUEjhFbJl6wwaZre1fHSKRcWS2Mlzp5QJtxA3auRHJlvQ/nAwWkFU
cFZ/Nagp9i3wRgfkXtgJJXYXcwErIll059reiMTJkH7CXUlRWS5OkyA/uAbBA/Kk
z0IdDmwTWNL0XGk9BdEayetHgj5Fdnj7d2cdxzXMnzEgLc973G0gf8JVk5Sh4RZK
7qiNanzm/wkZtqGNc3s+JrbkMEhNSNwUEjIPRXybbjet/Z8uussAMNLnUJWNXGOC
nJb/JbBEQn3MIH8FNqlNHCWxUTQETAN4nWO0/ucZSDfXWHWfvp0ZgVf9W32+mCQv
VaPa+DZFeMWCBOIyG69MAUhMDjT83E7jI3I6GF9mj5vjE8eVcR/11ZqLJlXM1AFx
GZkj8AtE9yMjTKMMzMWCUVkleT5J7qHO5cfnGjUx8Cj3i7ZsQbfajzZ6tIGpLVqZ
0fmxSWodhWE1YgoghGbxV/55XKfYBms8HG9rRyCSK54NuJRfABBN0VZ7H5+wo9VG
wuIduMW93TDpXUpLtAuZrBWRQ7cUGQsdJz/J8j88SnV84wDUcctdMW3U23WDZx55
hFB06BUiT1EwdhhdwjPwcASOptG75bDYcPNML7TUPlwclVfT/gCeC0Bs+AjYHViT
yrKHP0/LoNXJ/PJ2z6oYdw5QQe7QtQzal25ci53fU0yIr+MkTNqLK1eNuG/4zCt+
sN0fURdBUIPsToHmVVOzJ7+iPQZ9amDy0j2JDJhZoSUeD8o/rl107SnpngwHDoA3
IEEetCOjEL4qFrrmbULckO1eXO2+BRIGwJi2fy/JMlF5lKn1S/OnjrkpcQcvWtqw
3Wa9vk6Fy77VcQDsqHlh/RY6K9/CRLq2dIhnLvHxdB+UxkEp1gZJYYCVE2JzJd7w
xv+RqfZLa/oQ6Ab+MSamGSp0oaVpTMtZkjVX+avQ0nsz/vh9iBoVrRT6iTnGPXFQ
zd5KqUn8zPr58Fb53mASdh0KcqY+fZ/XxAX9lChimsGZ2W67r1HkCJZvyeP0sFzw
fO13Z/WzbX7/v6eEZQfqiko0gG7RAVK07dx3og63bPF6o8OS2pwdYTAjV2YNGisI
7HhT/Bu8Mp+TqZJG7aO0IPkoaRw3j5ixrmGD7nuPopaxXrbrsCYp3SjghyB4TG8S
AqhokSnP1a7WGlUsZMqLTJEXgHiOqEpZ95yLDbhqVHa3nbjxOb3LB84OfAGgWsew
JuRODwIIfBhPjxvKhCogkZ/XYuk2tYRI/g5abXIeghMBTrnkwwBH4OleftQL9+Gt
3oxx7oi1DRwHQlNi1+J5g6ll35mypT4zxB73/UOwU2EnmYpoPeFmLG7YhjJMPUsx
kd+r/UClHIPZqdQpY//YqGikUDUw6+EWn1Ct7oa0dJWlVLijVexzdbSgs6z3396S
d4npa7j5gfBzmdKZfakTPibbE3l9wbJ9hQHmispR2WHJSlygQSh6bX30QCBMVp4N
2K6BGMJNME7L1NFw5SOFB7qwEC3ihpTvy46piuJj04xtpzjEUyYYLf1bRwZRAvA+
Sx2SQBNRPUbFo0LFnr2XvRD5zpsJx9RhkeLdCxT++2Iy+LaVdkVFRMAA8GbExvRh
EWUKIYMMvdwHwdiyXCwFQRAYYtSTytxD/kSy0hVMnHgN6aVEALrsEFPOOVN3hcCd
+zq0JcUZerJ6WVXkQqKUy2nNEPYME9OOuBhPPpBWa79jCrN9g3uCSYpc3WjJo1/y
Nw1n0wRwRLNUBIGKfdkImRrnyYaCRt5BvWvaW/+9Jt3QzxSoC+/cxg8/dg3AxVk4
3ZuzbYWVab0eJweFcNpCBgq3zaxX5lHqbfPNQsfFo8Wts7B8YZ4eLvXo+9MOp+Lx
QZ3g337BMn3MyyQbdkd8RTvK/jnc1+jNLJKxn/0l2W9Cis8X8rNwRlmZ/mcs7y4L
mhMxtJ2tf7E65SV8zPcxeY8eF5q9xQ7Z645M9mlADHOhTqFyCZ0aQd3KWY6oQZeb
ME8z4pLNRd1Hy5XegAPJ9RYCLuGlIEegAqk8vCB1YSF7+2j24HjeUAQWgZtOzVxo
3bGpoBMNVo6eHXjGgE291O7drgbQt8mOfNaBV6i4oMkkwIzOOoV4qwfDAfSDjcxN
rRXB12bA66Pn66kCCBUz4nxomaLYKWn5Xqw7PR9ReDBxGRNs7Mr0ZpLBzWza2jvT
3YZxXsb+/W0ntaJtD76wMjbU5HyU6hDWxXoFqokqCIoD3f5HfkiU8gW1Fr4In7m/
J71i8409kvmQ+Yv7ArK6BLJLXAIrd5xd7YGBBLZTV5rOzP5DCACVXh6ZtUariRul
6rw5m8zvXZSPpypcbpa8nwrMYLe9USJy5Ga+s3WVc70bmvjsMSmj15oZW7CY+cqW
jHNulfzdyGUfUC6Bv9BKyOysVgGzHl3N4gckyIXbwU3dO3UAflE/aFVf4c+ImDKn
LCT2ZTAQ+RlFr1weqNPNsQBraAH51eHTkLL1NLRovBXnGoOUJ2WvUMRyKsllAtrJ
ZOlvNxg1rQ/kWxUwVVRkrPeoAMHs16DsYnOpluZRCliHXZ0zZu/3bD8+xFa+SMim
zQrdvNNgiVE+doG6O6/+z49Hg1i7OfRt2UeEC5EWDl0d/IO5wNG6gvKe3qRiCoJJ
zpsQafxxdFOgjQimkRGBC6+L01AyLMoOYXsfWd9oww2t7x2TzIhLNXJQ9OlnYOW+
mxOetrdOjYkEQq/byHtoDgsw/XSGNVBgK/vWK8Nk5uCT6Svhzm5EFxPWTtUXlxEQ
WfdvMOV19y7PnYodvF2sqIpmaPQNWSizFkRnWcUpmnaFh8KCyto64Xg9udAKop17
Q8JhKgaVjEODVvsQmCFjeT4+MIVXi283wYwpo5iI8rauCs8js+52bzJgNgCKdOe3
PTROFV6GTQQ8+zY5iAuI+AQ2KIskuvBApUijEWrvTUfSGR3F8iz+uJkXy+UgFfs+
7env0rFg62iPGnX7C3l5GEdZ8KGIbuU/Z47p+1+a2hthbkZbt3wv3eYbZx0C7HjF
4LDXAdi1dQyfhLQwA1NKoCPhKsjHaK0OtQkyfF/CC+Dn4M4o9sVzRkj3EO/05aVW
9Tf0FYxj5mFBnymMbaBiA286/0b7ZgznnSZOdFanH577OduV85PO3Vv1W/q2jc2Y
8bg3ZvUBCLBnC+jsQ6jUM4CazYA3yFBH5SFh5+xEAWoQG2Ru3HyssG6J3SnDLslU
vNNQAqgf6Lmvj1flFbaMliabi3ax+w4n7sjO4+eY0MpFDi26ybd0zpkaxWs9EZM8
GHxhTnSDZtNO90C/CeVu5/f9Jhb5fXmhqeXr86K40YboLg8qZrgAsgCUFL6fw5yE
lDUcN9OTPi9TUgQSQCrj7qGYT6VD8JRTxbLP4E6PgN2GfaKrcFD+vEFpG5qoUD7P
EVnayUZl7OeKBtH4sFtIg8AcNqcctDhxEhPX7aCrR4F15ow5yRcvU7Gb9CdfkC2s
+cWkqutIHlvOCHXLXpxX0fVVDl2byTEuFYePLOWe0n+RYJtKl+/th2MCd7YeJpmA
ybr5BxZXmlPaibt97QktsoY2xFM1zpV+Rbdxg1qjK9ZLYIAKLs4LzXsK4NGiOc15
g+mfTctfEkhfPYtv1OtWHTEO6d/xoBiEgN06BPBL19doWaOQuVl0fB4WotMnkfHI
Fb55oUPWyaocxLPZKEQMbTieb4MIwWgvIMAbRiUPeqvg74Md6lnWm5QbOx5S97Px
DNZmpualPdPZCXPXoSyLuYTTAVafoyMDyjkEyQlkzy39/OfcVixhLF/3BsHLDu2G
5/ZlrfUctV2k4MOTxWGeHlUJxQuUC1z9ky/z8EG7EA2SL0pkvHAPrASGdvMl+ikf
nGIhxak6i/eZgYayLSstsJJStbOrIbukEAQRxROmDfaFFHafRpXg7cd/j5tU4e2W
QL9lZ472i5V5YBHUa+Q/T3/hAQt3AjKT/AQXWUk41B7M38Yp/wQJgo/4eHuzftHm
EEzh6cILS1pwZMZALsrQxXkDtiKj8YQx1ir5oDiokpZK0dNyjyTqpbeNUN8KQstv
ccPMHtkPMKVxbyIcJr7pC2R1/uJCljWu/gbqb50SM307bCNe/A8O0I3CXerE95oE
nxQ4D2ynFITp7lcyg47SiPeeGMYLM94GmXkMg36laIUvaT0y+xAuYBux7oYPREYU
EdfPjxYSeJaHbmA8pmXzOoWNSVMTZdeD2hOzHZhqTRCI0CLKlK+iqvEAhdqmC28G
Qg7KhH7uOGHooj1ShFKP6yb5eB1yIZJF10Q2TGSMN9W0wFKPh4NkICu7a6icNl/9
8xvzuEl+roA3zRA1BWe0wTj4/PyVm/0j1G84OeXtT/1WRkWPYVhStzPwv/PoeF7O
M4jeFAncjNYP9Ceysb/nmygxVwNSzafAlFsxxj4U7g2t1FEF/r/euBOORMtN7noS
TLgSYGCmCMnxcKAHdwl45VLLzMrca/b0WH9sbkYAoDRod8Eg5eXMkY8j7cc/eGld
pc2z8Lb4HRXfVU7dccgT6zFdeKouGv9bqlvEHBQjb2vWEvArldUC/W/aJ4l2/7Od
UALkOHm/Y3ALn/VT4CrkP7ML3I7q4wQTU8cTDwU2S/l1bW/MSSYXTe0lXPbMMSMj
T+OUmmXADYziGq5xjCAKPgLyoWTZeGd+mHk0rVzYDm9MzfBVHW6MftUvmtIHKcz8
sJABsx7PKjvp9EmX99XhjaMxpsoxO4GrxBWqkFyRo24YhSYDfFQVbQODoeq+XhDs
m735ruieTBeX/SXyP6h7GXY9qNHAlFLTa7tfSy0osFJn14a/sQXDSGVmbIyOmKQe
DDgq5LIYZcqEpMd8bw/GFGDknmXPAD1m4vkmk0+6N9PJfP0cToYiyTP/S5IwOFcB
iDcqOZHBr0M7uaa9eHzFDtQ/m3mHwBEx/tdtnvEAjeetun1FuCAbSt+sPC1N9ki8
VIiOAyGvpmRsIaIze9l9q4oiQz6eGsaNSXIFdTxcawdN/XtT9LpsGrocXZTbCsyI
0sy/EiEg+Kg3UNhfhylHrbesrIAXUdKxtLxxQZMv3UVL0GRfux7RlG2bj/Pks5As
chG0uER+6YR+PIrvqTPpLcArZzKifcWue5jQyhXVSztmtHaA8bLELs17pZSDGaWc
+k0PuPKnji1saX0SM31pJgen3JMhclHnnuvUglPhWt6fmrCWxyJ91vvvSWbb9vgG
UhAOHwQqSuzwBTdpfFGPDbUwoPJzfFudnhBcFdN7c42Dp06THYO44o6R8GHgrTFv
xcI1FctVgA1AwgolNaupASS77JUGEY6YBwB0P7j2Xa4cNWxOqWBv+uspUcUaG2WV
ozhHLoY5UH4bJj9D1IDyN3uGL8g7nvvaBUKlp/KMpfhXTCsdJYOpRGwGh3iJvYfH
zX8oWQOu59KtyMsM/Qe1LMJNSLi2SoaceB1XepJHx56k+uut7A8l26bx2vMMJORL
H27RB6H7gHVsATMacQLoFPLgidd1ce63whkHsDiMy1wV6o3zN1ayJ9pH/JaWTwW0
P61PoJ1JvNCnjCp5Lx7dE0Xg+NsA46cAC8ifLzmlI6KrBReB4RG5CmHJw0O4A3A4
ZCjQWfiRkIg0rzezOh6k8TRsEkMuYda92D6be450XW6DYav3Y2PAbr1wovWaP9Wm
vVnp/cNH7me2gbVNNy+QRtdutBHySegMuuzy4i+DRC589264cUaE+yCrWJr1vP3H
SwQDwxgDzZKiPX7KD8IgJPrKbH4Nw/8aCnFuC4kHO/jxSRTe8TSqD9lJoqi9Ci7r
UFOBFkausXdR6M1gyBXRbdStuvQTo3KFyQVJfwlww9bgnNrk3LBIHetnTS0DcMAJ
6ugADb7WC3XPT+tK1TgK1vc2duxcroz2QV+Pwbp8eCARalR9p97igza7sz1rbiWD
dy3c6JPf4oU2a7S5m5bMvaAmoyeKmtxzMT4bkcinbAfPDkiguuECwBgviE0ZmnwP
pssdFYEyPd7YM/lY3t2NZYB9Srz/cNhVaafs9UfFCu2kp6AKZg2xnmf0ylzUHUpU
Y6iredESJ3XenVD1Cp7z6zL5UZ/YoDjb/4a2/ua/L7yrGxd5CliZnc5Ff512R6JY
mN7hesZ5m8I7WlBSFswUps2S8/pcth3fQT3VyMd9z8eGGj98wosq94/IJI+SpON1
dDHYmX6OZ3MbTJEpPtUOL+s4bx+2HQ/MDzDjGVzyNvgUaSF81pFxotZHfK+BEC7d
5RhobTLDahpp6DCl1UC7kDnnYXdhCwJf3PUZ84+6hb3Q4hqHddo9qE0zTVVLMSHJ
98NsUMrowE5EVxRacvbf2LK3sP8/UHGK8gQZ2IZ5kipD5h3lHsI9t+r/ku1Bd3Zf
xvxYznMKvXw9gkMpMSEXYrZb5eWWOF8Z07BDoUTGixl94jYHX2Bl0mfSGyJI6OG7
a2x4SbB3bkMXY5vFo8qH5iTho5sIV7GgKTCooPJuTTmdHlGejdUBSWAPQHsaHHiV
AH3zFbauw+z/zXZqKMbl9VE4d+JLFrpTqXMJkXp5O50pLzqvL+qIUdJqMZ5WDAN7
cV+RW1Gd4LO7cmsbad1vh3EudHA1QoDvFGk4OeR+ybi11brN8pXBxIfvyUlBl4M7
XXqh9ILGx22jj0mzvUZNYTqaq7w0pvGcAAGCN9XBzyLSx63BCzFY/p4Qc8hSV6TG
G9oZmVqlHiER1gjt4s92dN3f2JGRVipuXoAHa/uKo/igtLtYNyzHHoYi9CPsAqHF
748PghfKKmXH11b+3RCjtxalcwcOfOluHcnSo6KJ+GXSLCTav/oRXL6QKH+Scp2W
obCjQSVTk9aCLDh6ZPwVlD/nVgvqXFt8EYcZpIeg+/u9ecHnSC51+mFTzK24jQw2
QRkU+X4l0tJhYALDD1FeYpHuHLjmVb41vP9vo6Ronkulf2uC6Ukhmkp34NCQP17n
VB/VNSvROARIKtz4dPW0YWazlJty9lnM+hmsLGHddvAoqikrac3irDKwEPvUfHfg
CrzkpgZaN2uSSw4kmJvli6hmMi4moi1Dggn6mCnl+a/ZCbD8sO8jzgdYxLCYRAxg
9zFV+xb3AuYxyQ8J85rLaJOwLuBHkikab/8R9ycTYciOpembJE/rdHRvMFccQmib
++S6E2n0frgCogMCoRW708em+i4cLH9Yfxao/1EgWYl0JAprmnwZfigLMcKU2Rzm
UrL/pPN5q+WOgBLC+qraywROP3ZtrE2I+ioQx68T5jbkR3VWeCgYAGl05XPYAfl4
zfb57fop1i/tPXrVXqpemMeajDi/9tyqtgyQthYMw87fWs1cNeDr9WCs+JVyVKJW
wOJOzH1UuJwGqH/SkeyRybQzwBvElFKk3j45SavLPKC0BQlyBQ9gk3JQMQMWJEPj
BBe0ZpW3d7dQtIGjrZmM6EN89ZPzr/Gf7KNKoEJKQV267svMEufFPFxITNmsP1pS
TOUBpCqTgSSOk5yVhKNUDsoyR6Sict7AKDRt8wjhnyr6X1xntqNwt0DunqSA9aAy
cGvRVxwGWawxvc7rFWJbFJbaDX1Gc/DfwrGHWhlPXtZyudhPeUcQrLgjMFFq+oWk
EVRUS1Xu1lGESfHJG/E1loZytEWjmig28xFL7HgrwXeJb8ha7pGNA08SamCsF9jO
EDJr21kSHf3PpZA2gcrhTkni2g67PUvVdSh4/yBNlUGQYAhNgXvEsXRsQzTn2Xh8
+5SxsDHJUxg9nIaI+MoFm/t3mlw7MeSN2N0Jnn+pXrFxUKx7wc30KW5FHw5JK/0x
4Z402Y7yKettqY6pitc8c9w9xZWs18UeuntNIMmmJWiVsorcJCYJxBUxF/6KLj4d
8eCe0SLh0azeU0voFNd8nDztNpgL56lcGkj9gxliHANa94SCsm7y/I4SVYdXIjAS
hI7f60gX5i6ChoMPVxie23PknSLEAaQUsEeTZS/HehBJRBKjB2MGiYJTf5gkK6Op
I9dV1fRE1aeNTC1b5LU+lRIF4LVWtRJ39yFtGfT63b6o3inWujCDxXPyz+pTQYND
p13Vgk/eh8UofuCm6KnjnE5Pnbjo82Xf67rC9sttEk99/DSXzZio6sedo7EW7OZ0
MOUrne4q3YL5X8mGFjuT1A781VqbLGEH4ttwvP2E+AIvCWSf+u8me3CG2EQNmO1O
fe2c0zPU1gYrW1uvjvT+7h5QggzBfLKTAxajirOJar2RGTtyAoikihV6yNh6PRtb
pH+CM8FDNPCFEJwo+wFb4OJ8/rU7aBjA+bY/pQ1rPS4vX/R6fc27DVqalu+dtGE5
8CeX7YRL1iYVCbWQBiREpRZKdFZGZWwo+IKpkUBp4L6hPWP02YbNWofNx/pH6LaQ
zE5lQNv2xHaLzOHwlvHXuB8s+fPobpo15IRgjfCO15JGTWgDQX80keOBzogFqnrS
Z/VdDM0OpIdg05v2hltwaoCpBJqq5lM+o6f6ecYG2qksIhbAZQ9keEsgcStzMm0d
ACm0L65i0uAjsv5RmghGlIXisrl9FmkkSlC84O/k/PyfdBo8Nbo08YxUoOLgQEsk
V8H2doV3ppzcWVdIZgsBuqGFiyjqggTwJt971Hw8dSRTbR2d2BEPf59g484wXI+L
iy5fdRaBr4J/+0FQAZPRnenE/fS/xDWtxNY+OMIlReDwTPnkLnUh9EeFsTUhzUGI
fEWwlUm+MU7aJMsPFTBU5zYcUSVGQ5Y2wdaoTFNUSghT6j/tUk7+vwG8AalLsLAr
Y5ZiYoObUyc8x3TAVK6rx6W7Gz5wpivXRDty7TXibVAa2EWutH6IQYL+LcIweN8e
PHhfkY4KjXsLFm64G+kXJYK1NSNjTpUPhrs/I/cIBGvZy85kAkh28A0fd84u4ka0
qR5TmR+ZhMAZvfkL4hQI00GzgYHCBsIbnWulX/ID9Srjx9xAv1YBEwiSCUVrR1zU
o89bzzeOaWLfjqB+RBHIVKWrYpz89TP85wC5O2eEvmCaOCJJSwb1+98+9nzNVnJ9
Woyn2kw5lPvyQR+zta3f7mh5zTW3UdOPoaJzLoQYaNqcaUnfYgbtMBaWT4CIpWZK
tzD3Q9pggV1zSAPa2sUDsmp5uXLZNWdqEKVpGpepmSAEDUTRygB0Yiuc45aVndtt
+Fw+ciGtgq3E0zIHJvYLSbmL/ewfOFi/V970wqwDTl84uBsnbFUgL2RBXwy+RdEu
EiXtceqgTX0Yh420GfKNuP9Q+ORD0BCVAZt9VGxbqvfgTaSKOL4sScJ/ZogYDPXE
rzmDUQx/t9gwk6ShOaQbTZsOd1Q53hMG4LJotmF3E2iK+/+cYYsodBhyd1ouGhW7
d4Pua0GWlAeUHzO4o7MC6f4SUL9bxM3a7g/Dr/1kncT27VDmDIBoPQm/nrFG/rKs
B5VCHL3cW4Y2tKwP+NwQ4C9TzzbQT7bfunqkJ4IaEueoezYPtdsCzMlBlOYmQ97V
4hyOgnbjD3H7JcLYioGbAPnJTbsVP24QDD/LL7QIefA3DeMNMtT5E6oDE91lX8xM
CEEaYHZ7GMhGIa6jbx0qKybyF/vnHh/UFaPgSt7AACs+QiRPr3lbxWZxpP6A6q4r
IE7YNwva5qVzUgEB+ALGYNJRH7MU6AUekuF80yV1Ip/FGqYZcIRV1A5RGBIzIJkE
85X4PIO1+iDcrlqr4S14kWaqWsWYzKFf4S0urDLa7/8GApQIlPl6Vym3NCdVa86/
AqeZuJ9ThZFjrGvlPhdp6Dc07EpO/eOABy+F4L9AYXiXC543JZHIVtaSlR2AoRoe
b6Irmo95vOD58lP9QIBoL0AF2JKkwSzwmTeMUiH6Tad7XNqydoAqGrDtcC6J8r8q
LWP2JlMs3mo1AcOKNu6OjYWC6XW+2dEb8O+0cqUF9UUp2sJrKE2Dzgn+JivjhxNW
C4vF90mj0M4nitmHalIC22CB5XEe/Q8Hop+oJsKsoAx/Kyi6khxYU1ez16pOuEoc
3VpMA9X42nCWBlezNFzO5wcm77COgEZETcNy2Q3tXEdT/xdh819N5wVi2DBa3rqT
Xvp/ihkLZspzPRMSGIoZqWB/kwvrzMmQrwiz0EyPKBzLEfqoF0gOwlSnCF48Fx6e
8Go/5Uy9oxA2uWCPB672mI2W2RS7hzBODwBHdzmOE09WVsspC48e2ueEHbF7RtfX
2o0GkD4EHXIqPKyHori6944DOBAo9ZQCZtcCoTmns5scERD0C2+ciMbrp2ApD5kx
ET6Bc1X5QgNPFNO8zONdHPEr4nwPQseck5lhUnMjuwrxJ5t0DlLoU3XJgs01Li4x
J9KiiliP8OtgP5H2kJDS7e34I4V41UYQa0lC45FpETXxVNt4bj0vzIuwQo4iMXUJ
RuP/lMEi1Tf140pHN+rQ1Ptx86k/RofpXGOSnJdlaWPjGM1GkKtxHDj6AHPJhK97
ZXd9hCpZsW6scePc425QT5vHljN5i6mJW2TSvv7f5NQ5FloH0f62KirPo/giseEZ
OjZIbOLqbHgNlVSdmuPxvIHJdbTogoQlLZ1Uq1DnYyVqD2Y6HNgT6/CSq8lTnucM
/2/Jp7Kmiuzk856HHHwHLOtM618V/vgpFBESVQBL1+XcsD9ijfy2SboUmilbo/38
o0qYtkcBYV6GKbLcb6KQk3nXgvOqKqAzQTl8ja4akZtzo/gBIEza8F3GdVwdgj1X
mEJtFpU3eyJdVe2cHAdB9EYFSAPD3l9lUcXlEYe2ywEEx8z7AzzWRv6iWuVXQcAD
0rG5wInuNQ/JUH6Gai3pZ8cdT+kmUt2opWZESivejHwYPZOL/EAEOAHrJnIfkaFD
A/I2MCikFE0enX+DiFOhUMYuNID/aw42rTOcjLd7NL2eTwMqQcMlXkQesAtw+un7
sbz662LWfFuznWgro2bfXk2jlxRqm9B+K0+n5odnvVH9Nmuyw1KpGZ2VKQuRPPrx
ln3xClfBv5Skch/j1m5czwYjcv3IL5LK4nzaWfRgsp8Upy9O6yq+mJeFoQCeecdX
SxEYP5NF6VxFG3l4hu+oog9fiPHF8ebnQIWHuIhQ3wvGpSsmm5vn6p596834RXF9
SyALRGIHEBQUiv1A3ZKH0xPOInTmzmFO2oGTPyMVUdlhBqTJFWdtWuGE6RCnL7Dk
AAsSaBh3c3bJaMUaM9jPu21QNRZHcTg2w+o53OU7TA8lswrWNleaK/AOAjYVuJEx
B6AuTRNc+uI2dGY2hnXvT0LY6/IJu9O1xN1/oln7G5+7h706hrcMvrejqh4p6tHd
ur2kaLcoBJf0oTbz6LynOW8KLhl/6C6gXNK5WebkXf82U22579K04a/i3QC9/1ss
w/adsSFe4Fo1MnteAEkLX+qw9vIb27EEog08YVcvky+/ayeRWvZ8WYka5+ipN6e5
QCqFsj0fjHZJeg0zXc5X+nELUdxfQmMvrlMoVX7n68qyk+F0rXXow0cEaX5M+KfR
/vBsxbQSFdTy9AKyIASu6hzWmNJyjMD1N2JT6v3DY/L/UYoQZ47FLPriqa3YaXps
6CDQPOAWyXbmmM4SGE0Wr9WiFKFUhGdZg6ZnUFUwXHxGZyyyVvi6nLp3QPyOsK4H
X5YgOlovpEvc4+ikgmEZgYYB6oRWXWqNyJEpgIPQesTq7Q+pH7S50yzli3gNazF3
af0lCNgJVCwjtbLWuUqT5lZsoTzro31yyPqPQZNZjLwGU/AhefI+pmnhvI8xusET
fscBWIFWsKAVUOyo16aRwmNlTeCLlm4wWrjiy2TqPBLSuBjQc8KFk7CrxEnLI+cK
gOQ4IOHqHVhGligemZXvjyI3eJ4+4/LFb0oQmUZHY+OGwZB1hMkTF5Kz/snY8UM8
wk5UpTyQMg6J/lPi0eGyNC/fiKIU3cIlz1FEik+p57iFnqrcMCq6l3xtYfpWmgam
xTf+6W4nEIzfZlBRMAEcPNg2dTp4q+0NcT1uDRvEiWa5UAqdUyKyjIrvj3qzhkrQ
gG8IYOxLv6XpezREvS/r9uql2VINUmuAUrr8lIvciK2TIGPHdOfL+L8GJPEeR+3L
mISVLc4aOuiBAbvX6tgSJrtsF5ZNMkZUlFbaBuj4dZ6UOLeRqhHRhw84ENxNPoQh
Ihd+AqFu4lQDCHdGOIeiZxlsWs2duu7PUBp4dpKsGehKiZdo4xfVGdhLVFkYw9g7
SvCZ79CjRvScsrCYYeLFuOCUPt0PtF+UwytenmtDJTo9n5Pw3bOPS3VZWhK3ApTW
FIdKRFRLKEEugjcpUCalxmo9czEYpHFKItlogFBDBoQ6LAZ3I9KVmp8Wpt8YpSSG
S8Gc0Rm9W9kisrQ8W7DZ7CojFBbqM1bcSfI2P/6g649rjXOgrK8P9C3TvxklHsR0
Mb54P/kN88TfTMDGiY4e4nShKvlV+lQGvgslrompBfyCHYQTHUWd51FQPRfd35Ky
xh5W2TVkxuDqNHvZ1tSL9g04/iqC9UCfKXocAgjlh1NO9eaoNbRdzJC+TNneCVl9
camH7iNXITTwLAVB6vwW5zn910jWCgAdVgNSKmP9cXHvepqgX8PzjN5MNwfABIoc
9X3ADChRHz5Wg4wOvRnt9nQC9a4p569zGzcY1RnNwGLkGO1nqAosVHEjYtC3jOlh
ph1XnvPe5mmUl0GZChqsyrP7+ISTs1vLeT0Eh6FPXZi5JQx2wGeF+snBNjZRUNIP
D4Nebbs1HvOQIX3Q7TlRLrTeNUqQUNZoybo3it2UFcpaCraebi+TRtO+ZYiYLq5Z
3lk3P9M7wdOxhyMdTmyuyM4PyHWsXkJi75RYViyDLpf8qy2x5FIYwiv4EnkUARWW
LijSW/gmgVhW4xTpTGOfcdLcNx+tGTVrpm4UeIYp/ErW46iybfRtRd6XtXdrLZrd
daspBDck5nv4RB9JmErBa1BnofWGRo73ifVXVtavOKfU5HYOyDz99/HMAN2U58DC
pCd9yfnrU0U9d9flkAOROm5FDTR4loB9AJv7/nTnFTqauPOl32gA2gA3D8xJJuuk
+YYL9a2vqRHvh6hbMbPk1CzlMqnN/+7hJHYracD95TK9LCKFcwP0Sih0YngUhsEk
22ut9VEbq53m8qJMYU0k5e/h2UhqHKudBNIWUvlddJPFobxWwK9KrdGPBoFt/pfX
5IszC5Z/7izGeFSLAiMFIFzTcu4Ej5iIskLsnlm2dQkpFbuwSjmuYRxgjomjtBy1
60400iIavs2jJulUilmzWv2VT1Df8tk/bTKW++w5zmYA4Ja7FLI2XmZAyCjI7S9J
fTPWJ+o6PCGgTZxDV2g49Kcy91A/srDyxZJtrTejojUD52hTV8NCJ57LFegGJztW
tSOqTlL7JoOl374NAobYAqftdowmYEaofLL2Uw+l+QKhChdIPTHET8Nzyki/iiun
W7ZXB/dhJqfcq5Z1vwEi1E8ODKLrkHuVgShehkZEmhNptuiyS96nPRv0rsKOhh8/
Pj4AEG8BABLB/fR6gin7x9OykpplN2WYnHkD6l1LlJ50BH88gYRN5TQIESLnNVxP
IvEUNarSOzew6r6FZf3q03ntmHkcpN10RbkbkRudZOAmvZu5eB+0/JLNm4qU3o83
MSB15tePNO3a3rf1WxMj6ii/73EGKg2yqcCMhWWNvHpKc86Jfc0kf2j71smdnlHF
TbpIZa2A9ICRKTMOy5HU9CFJ+eeUmxoim+jxjizcYF5YJK1AiJjGKSWqKSBnQ0NC
y+zdQFjKVOWATI+02a0Rzv8HnPJuzTpFd/p5P4AsqcyN9We2vgDC762A0d5Xl2Vi
ULsyxrX1UR+yCminvGMamZHL9906lzqZdroakaEK7MMAQ/nsbNyQkvczmiyrU5dc
l2eJDlGMjjyefZst9ZIDuktvOVdmvKykr/QaR0ozL0sMirIuUTNXQEYBHKK6R7mc
fbqE9z/dwYU2O2MwlI2fKJuCime7carkkYRgWMTpBjUMDPvFZ1M2fTXEBGhpbuxe
ZXH5H8Ku2mr++/c2Ma687In9jgWP2sdpC7W+vSsZ6daL+css1Tp/J4f9yBOrL1Lh
dV/WNWy24wLwAPcv3Bscyy51bJGjCZtFi78llpWlV+1/8uXKWmdnnE6vvgED2xuK
xaaqmJI0V4XGLoOAY6TzQeTU27nDq9vkAYw1jc3rdPuANMOlKG12yxOBxRN3rNBS
B8RFrUe8ZOksUEYr31u1fN8NqQA5W/I05PNmIh8xn412B2BC/wWGKTUUAox9Ypuz
hkJiHI7pFkW1ov4qIi5osb9wz6KEC4GVF5Z0OYDw5/IkiXx2QRjRNyv7d8ophI52
s3Tj37mYR1pEE8qKOZK8gtpiYbJF4fyu3EdTNnbrLPjyhBOqk5QVwqj/D3uGYe1K
EUpzq8m7HFw639UVui8crlBqN+wxlElty5y6FarI0rc+UJb0U0Tx8xBWzFymrm0T
VBTF0zs/d5EGoxSaHnTV5ZkIMPCc+OAClUBVqSTQF/gJbuemSE0oRO0cQbc/JJfi
Uxed4n/ijQrkBtfb4yZPxRMQOQJNAFcquPovyenD9n8IdnFzyGj6hds5eqwAuR7z
THXdsu+qbFIKI2JQkRochR18p1j2/7hq+T8feeT/bozzAOudew6o9Cw6D5zkF9i0
6CeUdl++Z++0Zb5JnkD2OkQHZvMQb9eBS6Uea7Twzn4C18/bfABsKlADE/eIBQgw
MVFG9pjWPYmJeDSvfBknhKc9BMtcTODe/+Zs9KyYmNx9bsB7B/JmAb/eIRGRmlit
tSIHNHHySUCmOY73FQQqQnK4hd4JVm89idwD57VtwfgqxedTpdEgzRsl+HyEAV8T
64ODYkkXIHCV9hLduEfVlMYUpwpcZvFNSNtJBqzxCKNcvjYdNSIXlc9tBm8oBHqF
0nsM5FuqWuTIOaN5xdZbnzWfWXsHPRgqcGZvq6sLJXSuxuBQ2CHzzfnsab6iz/W9
sb4HpSNkZWzBFUEsl26z3zbkH9h8tf+VX+ZQyRG40Zw/89o2qTJKExSX1SXAupAK
M+AD+GzLtl/97faNN9twAA==
//pragma protect end_data_block
//pragma protect digest_block
uqV70tuYl1zVaeSjsTvZG0ej1wg=
//pragma protect end_digest_block
//pragma protect end_protected
