`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
WCu2yux/bgzrx2Qo0jUPSOok/0GEe94nnTCIwbf19xk1uzapAy/8Nn3STnutDOwN
+oXq3NCyTJUrLUxDcekgVSzndY459G8lqjKMyPzo4TlAEiQMOVA9mhUtC4xPz6Ys
IiCZZcnfcPn4H85NrAEi092D+ZXx+uprNU6AT5+lW/s=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 7120), data_block
ErzW6ZPCYkApj+Vi3y+d4MPJi134EEpU0fWB2DnfeY8lPJn0epjYxDo1Yp3aQ90Q
9QoWHtLvDAE1z+aUrPWsJazH77CN5HWHpzW4w32siZuLJ2s3do2DNm2+HE7yuL/s
sULljBVT4FgfG4/Lwd07HSh9jNszPj4FgUYztWIVCMDX8Lv6afjHcitJtn+xab2D
AKTky4wWQYJExG8YIYTSxvMDIVKKOPk6NWdDcSFnyNi5lcqzVj5NFysZ0PZuOpcq
rsg4L/cPFN+Q88tIcwFptqCBEPUznXPTa2Pzs9RK3dGrqBbZ8cf23uh8sWZnRlX4
8rka63NiICBIsLauS5lGO3EMcUUjlMIBRgBDPUBes8lcPsaD8YqdVvT0ESK5FwKT
LXgKaD87MILwIVGqBqodKoBDb3Fg8nCrg5cUuP0YAMTljuvky8l4EdTLSh3WPy7Z
1XEHJ6ZGnWVv8ciuNn2ab+S5TgOKakeIGjnmLXHQ8+n8Z9MFqrx2EC01tRZFspHT
7HVwpu4tX9qEeNZfhhwZu6Hzi4wp37zNa1alxnMLyuSL1CbIpobQoyp3W2soYNdO
Dor9wr1Lfxj9U0UAsSMmH4QFgzNr8yDFE/i0gsxI8nKFyvVVq/JHxe1Xlz7vTQ4W
KMy6gGgSjewK9Kl3ul8N6jkuP58qVZn3vq51rJaKS+5k1/4SMHEKZQHn41CBiW3D
ceXj8Xo+//+aWJXpHQWB3qMYPlhmUPmlK9dnX4T5eRqD+1C5svpz1G+Dnm6PrIv/
cv986eobp2ZaUFHcGoP25Fzv7d5b8UuuiOcEdCXSLcX4ug/zz3CsV1vmkRamnF1c
OOsh9DJVgqgwWKOf5D3shrXGQP7aT5EM7/rDJL0xtsi/vwx90QxNH3NbwImZUIkf
z/0r70xVKlicP4O9IfHjG+nfLIVdl1yV8mR3n4PjMZD8dCUAwbbcDQPVtYGdYvh8
sYyrwuNLdae5McNV5QPfnltiK5T9EZ2/ixM4Lor7VYr83dqhwki8m/ky1PuUtEEa
qgvLnfBqjij3D+1jtQ0VORNcnilKT8rTF0uvrFRC0yy7y1DfoBLDbZ/d/kho5BTC
K+E/Rrs+sm3XB1Ij5JKG0syyTdd2tRe4BPhMM9s3uLo2K/UL+w55HFCN8yj3w85J
Fg+LvoCNu+fCLjIRb45f13412RbLLoOcuirVLzWbaB1WQAzKKUEWYzs65eAbzdXR
lF60Yq70JnMuN0cx7xPnZmyuiMEYpJHFO6ZjutHnihvk9VREYTJ0zrdzRbBpBsW0
HEywt/OgQkOzbHZRzPPXlKsKQfZf0RoMtLEkkUFqHxtnmXUgc36/KPThCSy+eP6H
WrekFnSEstIzr91+n/5WFlZzCC47sQ9OYN5qrd1UnPjKl8N3NfcJ1DHkv5pyv2pu
6KR6k5ez3UFnLvUw+32fM5Cy9Zg3S1qmWuwFmk+c/Is41+pANRCHMInb3vqTCoa5
YZFm7ocDEPVS9WZDM7hLuFKtooVEqwY41pMdghobUQDjHKofSqUtNJMRsxeGqK+U
1d59FiCcNIksIBONAtnSPvbgPzDqf/veR6V6z8jXu3pMOcGU5PDCjC1+E07tNx0o
ZNRT5OO3rMwq5X0HGDt/QdSRCjHUSgSItLcrAnWE7JqlCT+BNlGJHSUBXhdwfSdg
DeZ/UGmuJ/QwNCCoAjcjf1MwJ+CLXOTBZ502DnjlEWHXb3TbQf6VhWhYoXR1sbQM
bZlcCYq3fgL8jICPo10K4dyPqViXfCGUMZt1x07C6o1fY7k3NwAsfJ89JtNOupYI
gHflVb0gULz1Fh2y87NqdYOKe2/u1j6Yo4ySDcK7vOtMqAwmj2rZBwwITkzFmdQD
+Nz7S7sQu8Yk7BX2Fwqe53PbrNBIURSyj/Q/H4/CVBkzkHk52M9/o2ZPATm+Br/z
3Whutxq3spykWZWJs5B99OvzwCKs3BM4fc2wKYuXzSBnRIC+huDHOWSGoi3eBDm+
owotBK5Ux2/SeXjihlyyOhXA33BOA9b160B+vVt0j0G8hhnKandDaHm3sjHfRGKK
lsFvdeHS+l6OB/AS3IkeFu+DF4C6oHVFT26OY26e8OYrrZ/sDTcJtpHrx7zM9Q8r
M7W1snGoA2O6T9zBfGZyANcIW3KYWwB+zTXsc5Jbgsd4FJwF0tSS0+UTA9Jj7eZ5
VkkNPTuJNW/psF7rVRWQhA4iDjfI2ALwp7XD9xV4WFEVg4IO3kqCWqwxdlTb1cmt
n0ztb05p2r7/EfkLO/nONGuY4PaEiCnDqlGnZ6pA6LTwQXUGbvpTTYTksCCYAEdY
vzTwCOAZWM8N/HxXlRCRygJvkrgT5sF5hMGL/si56ZxqKz294x1HSL+XEl1GpkqL
JrjVxH1WRSA+1dItokR8VyrW/KYXs+BJnNC/Zps9SM2CZ+J3nrho3RetpYCk36Tz
ReVYa+JBd4+71KNf6h8QTiElS3po02wzew+eNfOfZZyphigeQ+rQm6h8LAv7NCMo
CZO8MCVW2iOZUkFP5EhkWCrZWjBkpLbPJthB4nFj2b2NU/HQQ5GpFInBp8fJH2HW
zZ4mSL0VmdwatLVOlrr4AehBstKsCtXHs564N62miYOkm65c8eSzgAlwYItZ6fR0
6GrRBrZZv4ZCKWpvXFYxwNhlvIzdJJ2koWoYW5exGwa8591NWZ4KlH0KX0xkiDGI
jkyZtbeLTzSXxzo6J5U1SjysuPE7dG/ZoIL45aGn/NuM/0Tuk0WfHCE/Mr2gU2+r
9eFt6Z2ueWJ5JvaRGGyMCqjYHPvQvEj12X0DoKBcu8NK6zeUAkhf9zOGE9efPoH6
X2A/uXmvYOcrfIWKbxGF08pd1Elgh7RwKoFmyYPhghj/PLkXJ5krgpxvKcM4ivLc
i7WaNwy4vktyQzU9Kyhx2Nb1RUU8UOiVkG5+In67LPKII8Kb789NYEXEnR9evIaY
+DlldPt/OFNbtvL8ta922opCOnb5IfyCK9Dj69aJRV0WQrXKU5X4/UM9t1dXLp1k
MFlFNLoXDFMatq8nAI15aGURY9cHp45XXXAf6JemOWoxb/OQXnfBxQrP1VGe8z1J
EUJpQcH205xjzld87BFSXedI3sI4GaXZoBUUQfiDl4ShcV/TYedLcA/v038T51VU
84Re1ZQm37MBEaRHdhl9y2SCVqWSDoXHBCRcV7oHG3AVu5SE6NmxNgVa9O+GpHYi
hf1G/t1FrXFrXoGQu4urAhy57KavU84qv7AzWOMcN3HUhaYgQnJxPgsiXb04etNV
aBwIBpOQnFHE5vNRBZH1hbzWxxGdPJR0+wAypofvjN77g9L6lGtDwBd0aPv4Ukae
0+CQdUrNCF3G0qy5NCKTRxqJ8PErkPyP71mBqib+634byQFBH/10KvovOpHR8kFv
971LRA4IUE2y3q+ZPuX/Jf2F9g5ohO3RFBv8ehhFqyebRopJ8DKcI9Z3attfWIc7
F9dBr+vaotE20uNK8d/ld1dV9EiawN/2BL0Ph6zPE+NkMNTFJ5PU+TGTrUY6W7+2
vKNNLwE83PwhN25sAlc1U1KMwnQhbug+Od/sp2A+U10ydAMdtk67IzVidY1NY1gD
1+DZqWY+KKu8N5FdvJbJVqIGHqXR32Ro9o8emmSo3tLpEc4/n/HDZxzo8Hhx2aG2
CjKvc0UVP5uoTZ9q2UJTlMtwic9SjJAG/p0OyhGCjmPLzxDfHYbK9onkZ/25yyb0
tQNaNDP4g4C73s35Dz5xhRaf+1wZdHTzoT3u5JiGFO+r7gkCIxM3L5vpo7mWK6Me
sw9G+dCu2HV9CT2DlngUIFrXGdMpzM6IKvsgjQA3QYo+u6f4FsRVDi0G79CIUVur
JZ4q3A6LfequmTsXVacHwPcvo9CpUA59DetHJJ++flpAc2ojlLIDOCp7KRLrEpnw
rRElfu4h1nRyX83C1+KTVYPHaAUFfZM+I4bGvrS2NQ8O/S/Tw305sNaQJkuz8/p6
XVgohSx2uPTl6dlcv/zqHsTgKhXrSyMUsyhYhKWlUS4U9dk5/mW6j7QYbWwLEggF
3Gzq46n1e1zwtbzi9w5PJwRPPQGOvOWamLiOcuA5TxEmAA3MHUGjQbN4xcQOemAL
0SwrGcy20K5hXn4OE7dTvvgHlJp7kqF5O6dK4/tL9UXTIUxnz/2Gox/Jy8Rr3DQ+
CZUfQ3Nxy25686wPTHNbFE29bXErF10/sAuRLMOPOLhnUSsTsENUw4HAswyQCUPt
3Y1BO76jEfTKRF5Q5X4YB3Sq3y7ALhp7u6Sc8wCptV4hgHf5Glu4CzmS7DLR5TD0
gfaKVhieooM9YQCP4kz+VYyVpriapfDXqNDTmpufBKnr7Gjtw3iAaZWb4P6KXTn5
5X8dKOxuUdmkhaoygRAAkhgu2vZxddIDC88rm1hBkVT/8AdkkLNg/jj2NrLBCcjo
8elojgzgOUkTQ1eVe4kqyzuTnKE0QUs/VG8DCylvhIc+gTskw+nsgTVsDRIcpwCN
J2GNd+f7Q+m1sIFhcAFF7vDrguZttp6lnbAedNz70AeW+ubdCoX4fFnLoNfCA2Br
oWxf99HvLwpWg0yx07dMQ1e+B3/fWIsx5KyunB91AVs7vUJLSXtEAmfjGirz130H
nuo/QahF8fYBi8k2B4nODn1F5loizESj6pvCzy+y7wPkpnkJlELg8K3ZD4i2nQTc
AE17SL9UDoC8oH4ie0BUmIPIeGXaSEhV8CTicenVWBC/UIUH2gPvSlbv/cEt49pe
TVBS4fhIdvfmPgwct0vZ0W0VciT1+9Wk4CVd4x7yqjKbVyITAV3+Y9/Oh5rVypet
nbAJK2qZ9T7qTnLzrNBkTvb0Z80UoVF2hf/ktXGUHKeJ+Cw7Rk1/OteMNpjFd5x2
FtAqGP25OgS6kTcdXRicEKI8SoI5fbe518Xd7kkcW7n3T58M/jBvzosbN+yWdEu2
OX4yC0GSciAXWF3ahTygqDA6pDo7LVVPICN3vx0WS7qPWAgPVtvrb8yLclqYWPju
imk7fct6cCBJvJjKseQ+6M5BzOslyjbLD0c3PJaThWcGWCGanHgt107F9S5diIDg
UsmE//b1dxJFaq5rylCxgl2+h/NtS/1mQzxvy0UDLuVgoCFzlDvNxwk0swwz4lQf
tYabaJ4OeYueA/HZl2TfS88kt8q8nDhG//vp82Rt2WIZl4+WaLmt743cjObHq48Q
TsAaWBLkxS7dGfpmIuJwXtbfhapyznJmilJGLN0Jc0a4+hIdkn7H/3JHbBzbeKu/
MmI8WECyue+ghlU+BEHCdgkggNHswIOY+PyMtJgy+FVijEFpCVk9eNAHk2zbaUx2
2R9RWXxFPCtWjHeP6muy8ExS4C3NPv6GSSpFqOjLKUz7YyhqGhdWaiB6Bq/BKgDL
NOQ32D90IojMrZPqN6W5OF6/EsSd7De8BH/SrLSvDow05IazRnKQ/sVgwTl3xV+q
qVr+K8Hy0g1bhSSPtGcph36azRq39amGRLigduxAM/wlzngaS/esb+P6iZq2OPOm
pQ/FZBY44H7wB4bzV9T6imbL7vQTjWCfk3qmyISqtALam3h6oiAB1pLpx3dbtyFC
1gnQC3Ck605RAf/K0pQuw4nQF69bwROGviFlpRd+mr8YWlO4vTscOFXzGk4lpiSR
zKRIbBr/3bI7TPOO2VMjK6T/9fUr6Ay31n4SYAChnd3DU7kIwUtcA16tf6GjFOO8
XCCKzVJ+FOGprhh2KrbkuBi75rYRGg5WPdVfPTC2JCzPpVeZTOktEtGdMrfGZWGM
faJwLDetOeXhRu4UAuXWhR247Wh5pF06gC70fOuRSNQuBmWEZ/RXCJP3oyJYkTSR
3s7jfA1SqBHH90OJL4Z68dKieo5boNT5A8zkjFYJFjgiRSwDETzKnGfKN0rJgvN+
ruHbLFeSkdh0gMGQe/OSFpZdFJggiMtR+CcZMtsDpTaO+HGNIKoJpRk1NVgKqlH+
Ydl5O3PpwGjPJtpiIMg/S27whY8CmJHKr64WxPxreki5/bIbj9Hcaj3yXLkHtRiQ
eleAsJoROR6tYvGDmYauVrWEWBY6VxkpnNib3uBWPtwFsfEXd09z95yXxedmhhcT
Jwo1FLpRpJkMi6BA2onsdI4Pq22wVQB27W+tiu9pP3tM0bxoy8lqT1lG5hbz/pOl
1VDN/JHHqSshIUeofHftxekNapmqMeHVYj4O6NXSmTQcJUIlN8DID6qIJeG5xiEQ
coKdodF5weSpMfsBqU6RP48Npb2iv4T+ccWIvbieOzUdouDM3HRfS+JghVsKdT9X
xG9sFU8jNQCWZZasnWGzRfrsZYEjAUPaEcFkAfh+4IfZUvLuSx27kJwNvlQtGagV
0f5CKl6ekUPJS24EWJhzBByE2tIypbvKtrG9MT3hY/WNmJ9s3RFlflSc6DB27Zms
Z1jdQTMDqWVHHbkVWWdmJoLp51kKpfynMMDpDWiTxXDIQnEFhBUVLlVyC80SWEjb
l983p3mfkzZuaVelaP0AFYckQIJkNdJ0MZjl/1Damdcnc7k0FZxbgRVHa+7fWI8k
IieY4LeWNO7zbK9nJgPV1okMVxoccFo9AscvtA/CbTmG5qX6Ha1vqpLvrVtWG5Qs
K/vK7aSzbXXowmEYK+SjKW6r7uH2aHUXjoZVYkcU+uTd06UAugBtriRjdPMSsBFt
C4WYB72oblYqGqEA/KpfFiwzkoz5ZApGjpIUWQQUnQbkSsN9miFGRuBDDM7nIRra
5ULg12OBDZg90t+azvlUF3FUSNrjrlYGtiPMXQkQai2GGp7Y/vfr/whDFGvL+AGR
HtuEwLHyfwmYXuACX5KA84xwwk70Z03Rk5Nc45+b8rP3UOIsalURZNFwhBamJW21
8sWaOokT/AHh56937c/cRr3nSLy6phqoTlKIWkMkk8i9dNEVumfvTdkt6tbAtiVH
Vg03Pj384uF2SADDCOpOPAMEdEQHW2MihcYcKUep8oYpfcXeo+F8/uX8a0Tn0s/t
UBj7W8oqGTOwWLi4TsP6usxJPvC86LY0ryD0uOqce9XqNBt/R9FTxd6q1j6RhwPe
crWL6g68+Jrce/HvWVIgugRMOYJeAHkbIX4w+ZCrjcryPFISh+CiNt6nj9BZ42wn
ysO/+vb7wi+sHGjDPlq5EvA50fKwbyjIjsQIBQSsvwUkyFwUdlvZlXhtPqYznV9x
2lV/wiT1AVkPd2h38g5JCJ2VAhhlE02wndodkKoQRxlp6B4706GenhQjZbpKe/g4
ophs1n2B9Tuh6tbA8/agSwkQvm0p/GtGi3qo9joGGa39EXTzLrD546h4kURt/hb5
3+RG7+8kJjvLfU0rZXzyrk4VF/6YmkYS35prr9lEFAFVEYJNC9qPybdXOXyPIkDi
EvJ0YBtmzLdJPKY6NpaY9hqDWEqsSSIB7FgLJ5tT6ckxQ+/PoKtxAdqplEmvD0Md
/CR7IG/c0oGmreiePXNBAJE55zyowoZN4ny9CW0S0CkLpu/ibSb1fC8CyPBpkzdK
LwkaBFBeXJ0FisbDTzf1d3jxvNaGQ2DZ8C9Z+Q7mda0YCGNAPKaTziuB0AMov53/
9hLD1Bsgwek4GlgQBPxdZskisJva3r6M3HdKGjJHXErRhJcPqHXpb+Hn5Y8jD6dM
8IjExDfJNn78Bx5M0H6O937qUM+Epse2ZIhUfSFLN1bTi40puPnOsAtMjjtVaqGr
WnNzCdeM+ycRIFFRp/GL1uUjubBLEB0av/pO+mNz/HhgiwynHNebfGU7jyhnoNKv
dd08SjBib8SDxlywTmcY52kSrDO7E02Egr9HS9hnZ9aUHMusB04iSKzMTMA4cld6
MV0gQmgFLM82UR6DWIOooobo85/5AfP6Bb3ScU3MbOhX2UjohqUBjTuEr57AfNF4
1jgWSq3HGSMgWfGPm0ziD/HjWqYvAF4z9nythdVdT1uddOwoiQWRxLa0N9+xPxSG
lv8PzEAtFjtL0i2XcGbjBPuWjhtXb8VvQabiWGxXfMZ2JO54m8yAbXemdARDrlge
TUsDhYQp5NdEKim1BWEcMp129cVZciSbmNptYW6KYX1Ib/urYLQPgF0PHptbxBcP
LS1Y9l4i7qhaQTXdGJE3vS/5aWV2ZgtwSWE6uGNUhoaO85WdhJAN9h6kob1jEnWV
lQs+RbCXWxBXY2hd9KtHCpO0/2Y45YVL+9inZ3BZy2bZDG30kfEWOarvcxvjbwBi
wDLfXVG2e1jtsNTxIdSyixSLRBDi6VKIQc6h/UzgeauMFZY4MNKIJ4zcM+9OGfzC
ssrwi+76s9ee1hfZRfk6ZNduyKRgPHSPjxHLGV60LOx7g33aiQttdH7ZqmFPubW+
Jlpt/uieA8Lr3+dWp+kEmhKoZG/fBYnOgDnUuti+7nYWsYSgk/AHX+7TVbtxVTrP
vK78Gk5QYI/kp5diqvGxpX9BKJt5ib1a5iFdfQel0az50QlnNLou+HzLPzoUbD0s
IHawJr38ru7Fb8mnb/OCNyorq6TiSA0Za9MZkaQnv65kmHOltwnorp0vRTcQy1Rn
avJcpExsFI92a438gi3u9jGQXVlcB/YgnEjaAkskiwdSK0IWiDKmSiDtlZ2wAnlx
sdCzMxRvZiHPgJ9t8bNZnJB9IS7yGXXIBT0SDncUAFRPQe5G50xfPOPY74VW4nuT
TzDvlzTqGoXZPrwe8V8pEX39dlgaZdj1wtsWFwxG5CTig0OoOhGQO043UyvozGAs
4LyzqWkCDa2PSN9p8Iwi2ONB0UO2Ozq1310ZYDVwpcUuIehAOGHTd4Pb0tWZK2Qg
hdJFv6qB6ezxzUBdnxSzeRsY1yZnJL5dx9Q2u44XAC8B42895tJ23Lbj+xPSLlRM
mB3HErY+xXxbZtuDuMw2tNbY7buaidas1DIOsD7/OJsvQJy9caNyKhyT2iWEXkJG
trsuITMs9JvLNXlSXM6uZrKt3iqY449DN26HShZ3BnzsTNpf8Ya1YrgddygHmhqV
U7qvac1xL0FZjjv3vWvS5J31lcT9ugI7Ngr5IuzpxYWRJ3If9s9gxRQoul/eo09E
uTVm9Y3tS2grgcn56g/aIX+U4gJiYi2zjr6xXqeLpJ4r21R0mdDvRZiC0WGd3788
DvxYq/0VAlQ+NrWxpUzE/HWM7WADK9t4FbNBKMrv9BvGHeMB1pbn+i7qmvTdpb/N
FsJ7rbJOY4WjB1QtvtGMLBAX/aEtYSm7kq4lP50jufrYv1giqjCMw/iY6cAQysRc
ILob+61J/Gemqzh4FinUwgh2hw3AEjNoC1hSvc7dGfb+gsgMO4JvD/AEXL+HBzhe
+Nwn/Nb9byDTLM5JUmQVdWXFsJn8L1AZAPas4K4m1eQn3nlKGnutXAzW1dFTM1P3
aQNg6dnZ+E0VeWUBAoDuUYpgpA+OOM8jnc1PhVqbMB66bjxraZi6qlGe/LQsPmDm
1hcITH31pf6TmP7LLoIXZ+I15Mi7Rs9c1nEWT1XkgIDiwjCgecTQ4vmNnoOhEbtW
q98qpizt3qeFk+xO8eLLNQ==
`pragma protect end_protected
