// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UmSlvw/Ko3SgPMj9GTaVCNb5SBZFULvgQm/ElYR3E8zOVzYCxKU2Wep5XOov
m/uqiZnWMFlddUDR7UexUKrZJ7yugL71t9OfMS9qPjPEsEnQgcRycVAWjgEy
dyT4fNbccmRzX2EWW0lG9mzTYp/lGy/Mt+qwY3zDuGBJSo6WhLjvaqXHk64T
JepoYvKbgeLuDOhjN1tp8bgKvDUTBef1bMLmFCnovJcJ/uG40c235rDH7HVP
eCKyOx2y2XsZlZIi/idoIucn8pPdOziCwCSgnEDiz7vNJ77n1DshdH2PsiBU
bfQptKbcXn9DC007IQpeDL9a5YrET3qvF73760RAUw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IpkxO7eOBaaZ47mbiZgRzfUPvyn2lVa+PAwkX0Vu33YC+xUrzgih44d8vhkr
uYEGcPPSLgQuTa6Escu+kCxxfTl/aFMwdaTMFKQbKGLw6hpTYM9WF9me2czD
nh2hTCraJxTD9tF3MjJ2v3PJ1c4QtcihmmjLbjHwoUSXoCPrm6huzkveFzSF
iO2jTNh0tecx8caN+kykMr4fjTEZYa8AbvbusvXCf66nV0Lclw9GAI8Vvnq0
zPe8SMWXup8U78pQKlc1uhPQMDticVggVUazDENos2zr6moyekVnpUIadgzX
22VrEsj6vu26fkTqfKp1KAzyeRmBXnslMGhZp5xW2w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S9fvBQjJ/6zBWC0bZy4Q5lRkEOtdOwrKcsafs/44J1mmv5/tPBD+AJn3egLX
3QJ48V0zNau0FkkRKW8d8F1F8kSrfTEKypdZ8sY4sljVUNaG5BonPrtwAKA8
gG6U5Ctlqyg5C4+PNhjfvGhvYXKDK5eszqIeIbSuaNh9PY3LoSUSvei+ywlH
9lHHcDE9HRv/aHLsLh4oHd12fB+Id33gSJ/CG36t9DHFo5rIF7YJ3OV3+UeD
XEin9zB2LLeMnBUVxvtfFJrWS+aAMmWGgGJRjk4/gfXuU8PTnqR6tKmaUKWQ
nnBWccP+Y/E56uT3p3QdywMkZ6E1ePHQQw1rAN7K0A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Cb8z+eSlecR0BEFWt3huKDS+Yk7R0YL9atA4TKySOQJUY2z+5QdXAxA+HsI1
RvCdntdu8Ob9kXLd+WOuP3snkznOtuYh27cSRIWQZOHdzj6kSvAdyQqiSfSk
qr4i6xFyxoe5EtwM5EcXgPqWGkrp3sxL+rV48EaWYVWs3pJQf2w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
BCPqCUN9GPEz39Jlw7YyPD+jQcD2PDH/HnaafJdytNAfTY9S8b1jsbynkMYo
jKBrNfOhCfhWUFbx0HZt7eW6g7lU1/dtWhaMR469oZLc+2IxRhONm7Sjwaiq
qqRQFi1ZqukKxmlEhTrDFPQ97IdweaBVoBpfAtbIyVcukkz4YX6VBDzmLeDi
c0/oyb+3cla6BNsAoXQmefu+XHNN+JLWjva4Rdi8Ngm7E3x0skp53/Wpwm0E
/w7sA36toukJ9e59snJCXWDoDEktl2mL+e9G+NbCYqba0M5Oxe6xD5+4VhGI
MGDPTIJeRT5b0UGDm59C7+/PUJsKy+QPvW9Pii1/GExnByQsKXhL8xywdFoY
FCcDAnnQ4JoXFEauwoDpBKqO5fBo6Dl4vMfkfB/g8hLcw3HGZT+szIixKLmy
6/qTR46iHF6GX2ZKS3d0UgTiYxJA/dYX8rJyusKIA45BvYMTJK6xEfBvinNc
RT9w1sbONKlaOEmwBqWbl9SFROv1MmbM


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KE6cTTgCxe4kGoDA+G2S946Pncnhl+6eyMT/r2FLg28//Go8xBnjGPO2fYxf
92truC0QclAoqXkdvizcucOhLrwEDVaLiYYQK/YXtp7xwt9PwMV/KfqDceOM
7d8//vghaxFvZ8thgfBS/maZFr+o/SBmPdHeIWDwAz8xiAXSqiA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rl9vpnJzwQhAI+gZtP4RuAVYAL9ESvA5dNoGG/RwpCSeJ704Rf3nj5v+onJL
E/Ed0DCdXriZ6+6Si7udjHALmGyCoBrisEsMlypOAe33rZLb7Uq2dIxrVV+H
J1AoSyu970UJzEW89t6DUHWY9QBjh74lozjhE2TcXjmvEtaIrDQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1184)
`pragma protect data_block
kVeYbEbE2aYao7YpDgDJBGrZiPWCpd6Jzeg4/6leNFaS23j7iU07ubmaOJ5C
j6AeWav7woSUsB0kpTjk2aHuc6ZWt3PkHe3DlrI2MD8bljtcDBFQssZMK8jM
jSggaVWqnoad9IVCEew/HWcPrFX2gamj6pwU9rjOP+uuPLRizAZ5ji2X21/x
Ssnz5naV8eavGn60ml4bEBqicAxqtkOq7K6RkDAIqf1OvYxNVcR+t22z2QaQ
e2LhtejGygQ8cL+6tubQuI9b8wUgmbzvUUxUHNv2FRCbD5xahixsi8pn0siD
tiBtBkjiVGpVI8Tty1HM2xrsnS9V0dNirOl6Kx1csrmc3p0fYZf2FIPF1JFK
E+iQ9k6KWJttBztMu9s0zPbFVuO+PgEiPAO5Vnvbsqlo/0QH+8L1hWtOcd2K
mtpS2huzFxLDgWy3QpA1yiFFcgJlwKU8UWwIAxAh5ytbgfnVJpUXFejBsK5C
cbq32m7H0HmD9NIrYTipiL9bflH5fKDowaRiUjptFr4+tWEuXIFrHbSRrhbj
XD9hIkPBpqir8H5nQEIPB+vAIGFwKWpYAoBlER2helQiFyej6+mcb8mqrSMZ
9B1KE2IPpfklSQbV8/XOYVQ7jrzMMXr6eBnzfr4X+YtaYFpOPIdTsB0P6Yzw
lBLahh0JSingtMHFDn2Wnxfrg75ZHxDpKDgu8KypTYM/vo1thasMBlrp/abI
rfjhTAO8qb5Hsf68Xvl0pTym/BHGHCqE00PWWJM5BGCnJ4GykfZr6olxFB9Y
r3qbPON/+Qz8AAZHjXB38bGciLr2/Dozunrh38QCCY7ULQNmJ/tUzttx3AGN
ivXv7THFMrKMgF7JBsgRlqsMBdqHdvHdXgrPx9N045AYWUKwn/W4LsTQl4W5
DhbjOQ9n//uVN6AEelYrcsUbw0wUmQWQUv6AmgqE5tNkVg8+Mh+HSuIW7ZoB
InFUIZAXwQh/XDbwLYI+UnsyyNZK80sSezpcZ/fz1eBb2aUsTHZtgnvUce/h
A87iz65YJ2LYcBjnp24xkLQaMCq3M8YVSoyCpY9tqp3MxTUJlpi6gn9bEyj9
i61g2/2TD9i3yxkodaj0gngE0ALyjjC/b3vRcdE50c2KZiMazrsyHnbaAKRm
/jHALrDaim5mmovKOK9OVdoF0T/+9+tdhRFOIbW8aOoLZmYcVb0p5RdcUQdF
gKQQg54F8a9VNYjJAtmNgMnd0A0CoBEiFJuJkO0L8G6WBidERjg9kV/npk6X
fJu+MZvPYIYIQDbPx7BbI3OBs5uiyrJq62YsmzzhcETjJ4YmMsqImI4EkoXM
OXcGJHqubs/ASvk60ENYzivsKdmPwybYfwykCZUaw63M/gl9FsP7uqFytBAY
nAsQOtkv4FqxkG1nN3grmS14u7beEEroJLQ62H04fW0Li/aKa1T22x1oeAYh
t4+dCIUmu3WZ8ttLukXNVzzdH4a0YYVldAXEPhBV0AwHcO5AfWGNinID3EvQ
32DQ7BwIWckA3Dedc5VjimAaSXbFao0a65/a1+VBNc9ho0CeKWJ9V3L71IgU
g8TifqiJLrQSnY5SXOg=

`pragma protect end_protected
