// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
cnAp4J5dB3joBRxSDDxnXYdpX7TpllUVJ0/834o9BGLTa5BHURC7YwWAkcCG80Cejjav/6UIZW3P
0ll8B324zW7Z6buwI+qjYDeMWwuykYwdPumfejOJTkgJ1Rr3hwqvP4/JXjZSx+qLUz03U/kNn01A
9ls2pN/jOjb1Bo/VNcg5PiSi7hg3kLBnRUVGUkJjIuiYISIvnJeu78zKXYpU2DkyElsTf4DJP+JH
BSa3A0xGxg2PwbF9hJWWW/O2eI33OsaCXlXupJvpgyLyDHKP4UcJWqPeXAsFPRA/pAOp9QH8ud6I
Z7IDNt1YQRnK5/hJAOYwyejfwAbOyfdaI22cwg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8768)
hHzWXPL74qT4Zl3j18vCNsFkKqXzwONZQYHJDb6UegTyXtCJbTEJv42jLbhyvOxmWNsO1+/sH1Od
NGjEDNiC18lsBg71COqKGML6/DzO07i4bxS8L/dGFEeUDmue9LJn9AfMKG87dV+Mk8Lz416FGxY5
30ge1T2+I5amu4od0U7cHKDyh8rYD4E3ZfPrIFF+EkCEp1D/itBbUjH9/kqQ+/JO/3yMNOn0ppmk
5Et8rky6JwEOuK4Nt8JOj7rI9xXvzfDeuV0Zov+peXF4FU1az2yb2Hb2H3OZxkhDtkfIviYEWvgu
Hc8hrOgVxeI/z4ar+YVTK0VfRbGxbqyC8yKkpP6yjDBCaENuuwItNwte9CfC6MT624IJgbb8b1rX
Z/MHEF+hJ+uDpkmzkIUQeutiWj0alLfG61s6rx8+Wdpe5RsVUec5/6BcpWJaO455LFXf+0ydfxdO
K8qFWK6Zad4TQh4Jdw8KZjvMiWcRaXIXgrK6KpyG4dm753Mo3rZ3jp/hn1q+82E44qcllfVYvAEG
OYyNg6DJwwT2vxFjiNm4Y73Mr0Ys4q5vmxgQ9ErTzdtc1v3gcbmiEqBMtYCeNeU0ZYgd3Ytp1gBh
qDu2BSkfwJG0OIBdrrd5DTof0cNloRiH2NuNsKFBaOyjb3nuejFSse4ieW9LyssorT2Tf2y0jxdR
Xj+E/ZHk2vuAb0XmiUip/MDgLJADQci3cIOUn6b6PjhIZxmxBQyLrRapOrzYNdOXhZEN9FI4sxTz
bSqAdhLwUzlRacpCjIXOnlDApAPfhtAJkhSzAqSw7opM4ee/a/TxcfSFosGCTZ8UFK4Fu8RyUZvi
cjQOWmalHKxg8M3vH8W5NXhzfOHDazE2VdptC1YZXodrnYIjEhKjOBq6Dy0ICLOrJiCHX3sbaLk8
QHZoY8itz19x6MD5+cIC/LvuM57zOPAbN5Z4aJOZcbMjxT6Z4gLYSIjUZiAcGywklA08Fx+ijw4B
JrzZJhGob1kFMzvnBouwdHh1duW1CksI/V+uEn2gFCbNzsmTHB5QtP1NqX3jzWrQJ0NdI32rdfyN
eS2OABCGpUEp2WNa4Vg+SNJE/BQrMw+GPQkKFCIRjZafpbmDEpMRFCzkBfomFMVJtjEyBWLF+3TI
3g73Pv/bd/Z+MvBLRtdKKtxz1oVvBSMOczJrWnLvBjw0oXV6Q2cnwdfnSEvAsGolVZQ+dd8m2jYS
YTblQ6CPi1HdvdMSmH3wLcf5kOWPWs1bMM2bfGlddslcIAi4HaCKLWIFlKjOGpbXqRosTvnsdJNt
HW+5d14qDZ4/iyGx6al46CkVA5vVPDFKOJ6xyI68gs3c4xe2W72EbJ67nrlZmmxtLSdUj5oDKlM1
jzOPv3MODXSj3CuVKTYfLqWK0q1tebBbtU8i91oDs/zVVoFOOu6LXf0JOtK66Ey8AaQmh7+Ncbaw
geAZc3gLZmrdb3Lkb5OncaREb40Z5NIBof/tDm1G/yK/yDkF0qjq1b0gGGeBEOKzfu9rr1HRm3DQ
7ejC7tQtpZCHx0NIM18tNEmqlogrni3o4nxD1qhPKcF6JRJF+zg+qwemUkTYV2AR43hvLNTuGb7S
D+j2Ywj15UO0riSSCbfiv6/K29ikYchiCG+pcFWGpve++amw38/eADvwuJVOnxjhH5SBSSoRRjzi
+FUjlqMaRvVcfbdwm/jvPqeZaaHFMZKcx9j40qOJz12WUJfJapkEzc2XZ9JbVJnL4RdaC66eHaL0
KzutEcpnINsPZPC9NCfH39+ePzAYR4w81R7qwSP/IXxw2HXe2cHWZNq7Zbe440S+eDOlYXdkQqfi
QV+pnYACL8iXvW5WfxO4JGvfJpKL1XrFkpynklj4b6uP+4rxshtTu2098tJrd82GvJy9GzhOqFYd
FBlWJyrwIi4t3BBasB4KC9pi0DlbinJAqfRK4IaBW20pHnLZX+4WJZPDyQmgVXNu7DsHwSg97Q8E
C2HfS9He9jiojD1aXDv4Dll7z4ykZGJtPAFM3J2scykkJXtCUaUcZXJNpxcgg+UMSc4gUUYMoiOG
SVNuzlpWoGFkESUjO4V6SCrusm+ewN03RZtYS5GcRYrskeSO5RnWuesHSd7A5d2fV1D0lmvsdaaL
pxB06Lha9ynCxxWx0m1sMbWSugN5F//ZB/YdgZrZ93Xh8EH2QJLHzGCpSak6ywhLX11I98OYzL07
8XJRiqqPPUeOkCx1b/yi8oVFcgiUjHtY6teux5b+0ZY8R0dX/7ILmP7I8/w4Apxlwjhf3idGyNfe
mSmwUIUeCyyTLPoe75Knf8F2KK7Aoi+dT4qCqaD/pj4/+hifs+Ye2QqAJMJlN29y3765J8STIpTF
AUV98byPQGygVjyeVCo6t3O89R+kYOi2KCe3KWAHcQMroeVU/63ouhmU1AmWkssUI9qk6zd2We+f
uICPy5IMv8CRy/C1ze1UiteeYTM7vR/Qe1Iw26/M01nUZb9vfmd5IuMcB7R14jo/Xmo8MZJSouE7
eFCxeGNorO8zYGzaSlZtsaWl/sSlshkkOegv50kHsenSoaU9ULwDHCDT9zuhEwfv2WxE7nRyPoXG
eBUs+AkVBgq0VlDXjvftxfeJsE7ZSzr7FrytdM6nkYKN6bUwen8NzckS2+nNmGekYSZqXI8PXf7R
1qxDMVm9SgMJu2a9ZdV8cHT1gRvY+adWqaUxEiJ7U0AlXXmYKlB742mhkTAuKaejjD5BEwQwIqT8
DL2HL/bw64Od05c60m7f44ddGTFJE4dHo4sLWQqJubk8pEa8jbgOjtQLcH4sLvm/8XggdAGrfTgK
3MXOdtN33cQ6YkZqvQQYyUUO7PnlNbrbrIRlva8I10oUluoIapjR0DUseI0rCNHe3ozeP2crEHEI
itgnKJHmC1iABhykty2TmgSSUFND5utaESOgTQ0BcafMceivMMtqr/oaJ0V0/oLELdCYEb1HSnqk
4AN64P7nh5TwcofzX09lKtx9yIHdmt+f2uhzLZMJdEYuptEzhGMpskQMlb52ZHjgA/CVgXL+ppIr
zDJKCs7qBZD1yxdRdqRv7XOx4Ro4aI5T7B4dqLbTWyvXbPbT2Ifea0H3zIOGYxeY1DtXWZn5kTkt
QSi/q1W2FL/LEPfiEu05VUB3/xI5FY2D/o3xESwGXMhUCA0WvuVFhNFFfJxRhmMhD2xxCPqFed6H
nWWv7Uva7uaq1760LvoEwqaT03/2kh7miRE8mJySqFcXWHUEIAbggOthXOONiz6kkjbQzj3AKzg+
h6lnWCoexJ8mmWfjY39UCseii/pajjyuFrOoQ8UgczXKT9iKPcrACTmyxCTHuI/0ilK+E758RELi
HFzn+uly5O/9d4R7X8GuJnPiYsF/nA9mT6CK+efVVrtb9oBQ8FY0qs8TOk879wKQWce1yKCDG/H+
hMrmfZw0dVmVMcfAlTPPlSu4XcIbpcXoYVTTC52z3ZV6EuvWwYfgxu4A71jbcksyh+falPb3emn9
XvGHUt5GHeQjgDqZGWXn7jJsdj7QW7D7xhmmX1Kg0tkCrXEnN0P0DQVFbFR0542/OK4meZqVjzE2
BwfDHVOd4kcUd5WEWG2mUwmn3NrAWiCAocUr3bliKNAH6vmCCmW/osAzd2G63F6IsXoWSAyzNLi5
FvyaWDPQq2wVoL8jW1BUF8+ItyrKSvbsKoG1RjkAZy0cyQz3XDx0kjiBt82aOTmJAfw9mU28qVWg
eQY1k6KRcHE34X4TrOM5tASUupGqiELOulKabC3EBFcaU/J+AKy37YhPt6wvXWpzdHnj2aSc5MF/
icRty4ZHU73F/lqNrSAOt5QtAvKD6KAlRq8pFEyI4espuhpcjbpT1GJNjfTcWdH9+hDsO5OzazuI
jen1tcA59fA4AvSvaJrLgji3nLAV9ZZK0B9oB1Ez8y8KlMHM+LDZm114Ux5fXKIh+oMSdNzfVZaV
/v6IrjLDAWZim1F4ERw61aecilOghaZP/fZORuO2baLU2jn7YC66kOW12/nKcOKJL8NQGl6QOVSF
FbkOGVJPWum7Vd4bufwYsNx+iPgp1DqYlgUZGlXNAW2nmZi0PRzObiK3EKwJ7QD2v2SVpvJvXxnm
TXrzZEHFkTpKBzlB03LJI/ULMf9fizdNmAAFI0Kb+4F3/jxfW+LM5oc8kmOYFG8UU7D+H4shHRWR
U6p9kI66MPDT+D4FKEkP8FS2gc6UuiufqC/FCriyT/d9idVQuuDkJ6od5Bu+doysnwD+Loil6QoW
+jAn+/eP4DKxr0fQp+ByccEXeKSYCW+uwH36kKWEIEhX50+iZsQOu1CDNdLMGXX7kgGUMRuqdmSo
LgyimJTD1ALclXHjVS1Lj+82ED52+f8A5sZNyn5suh03xBe1ZuVhMR3PBwVGQZsFBHAV0Rgkeksc
VbxHLw+W2iKHEoudkFtZjUCmzucuOWiFBU4TXCbJr8R9iJlqv/5juXZFv+b2P7TCH1HjTecYJxjf
JHMJ9sew1NMpksgPO70yrjxVUDOuUrs0bOB/qHXswXJ4IAXdJ3rzSk1gA+o+++31J9Oba9uUDdfW
c00lgSwy7QbLKJSR7ovYj9StqluZ/2WM8sA4aQSQX6M8pHCFEDqCwyjye+t7notADwTcuLaJqJa8
GXyE8LJWZXD9kPV75BX3tvGchzqkSYPNm1YrXefaVMeokSCka0HPxSsjznVa0Ki4C0hyuGz95qa4
bB5tVfHxqmodQYvvA/q8AwXMtooJX7MPi+MP4Nk8h5B3YEgOzuhrtyql88uPl9wuqURaahWAj26Z
/c+u6NHz+2pPZuYwkQpdj7rMmeyHnZ6t6LFEDLTZnbkLWX8yrZT+TGWYPdkDxmSC5R4XeZJfTDXp
v8miGP+HafLER0XrWR46c3cKJLrHhUbXtiC70D5RZBZ5LR1FnFLwpBz8v+3GOV+mkcGhdvA1Aj0E
YFlz8TOTPc7EoSzkC2iqSF0ajTVEUfo96ynszHb3HS0ms2JXJGopdMTKKUlHCmMQW0lTq+NI/i3A
NziQKnB1U21GBoYfwxKfq8wnOMcfU5rZNCnSkHfpAlgizFv3532p6sOQTdRU5OmQI1Lg0l+mlA2R
lSqUVPNDefgu9q3YDtaB4P88W2VcjLKBd9i7t0k9tfum4n66wzVqhQy5v7DD1gJCcCTzG0Ncjbce
kRyKj5oBvuo7t2tfZDpEgOYP/rYxDVErPWAlaWmzaqvHNG3O34NPpRnUwECE65il98+9QqVYxXHR
kEzObV5RLvBb9n/9cS0JIy6Ff4ZrIB7G1TvV3RmjjamdkZwDnjNIJd8wacXFXBtvJqplL7W7JKix
M1RmgFcretD9nihtxsOfcA/qptL2Eedkq5fslLneB/Pf5iUng13gM5LE7j9ysiF6TeY0T3kBR9NH
X/9NvyWeU3CILlW+dUV59W4v23zgIctKxqGhXNcqUegPhd8SUrRuoMBB3YCxo+DXBgqSjk0wKWHX
LjdXDCsXlA2F410jKi5yEr2mN3Jp2YKe3ebR90/w4NN9X78ajbq9MeSJJ4G8U8vm+SkXU1BD3i97
yL20PP8QnlHxx/ulTi7x5L51Tq06M/UVCXnn3vGXOn5Qrx68Wk33gy6NImIEIBm8cYIMWHmb/NCP
XtLssARP8KSPxEIywdEKwDGpj6AJ+jKhFg+iE74RiKyISEPKvm6bbLjyGWsRMnmiLSyW7Pj9oFJS
htxt0TKs87iX8YMsx7vJNarks3EJZBn8YKa9IWnTpfj05jHjdunp+yZjicLGoZwF8BXgJLbU97Lk
Df12w1HHHu05lHunGPyF+lOCEeEUn/V+mS2rIwt7X64y09xjxAwwTH7oymGZLOgJPGRPAaS0BWGP
4YstvwppiWWEYMwgPhl06nF5BQuCLsFuHc1oKFsIqk5aXB9WLNZY1jSrzLY+k7Z/KUg306XD9u4R
3gnanOh377NuvGnbf9Eiy21NtRH71U/kSSoxIY1uQ6OxezhIGpKY4Kk54JWsLnI8lE+dVfIRrjCe
z7IiFpiFzFlvLz1oq/FYB+ysDpTVTOEaYt4Il6o+mrVBuOINpIIxDRsFyRC7t1VkvTX4c/dfmNOA
cqbXc+fX9HGUT9l3c9NReY77kjPiuiYhwNjWJV9wl7Tv3LZjQnyMRRAIeryJNEWT2cTS0rhTjK+y
O77HkELddRcspQUO6YcO5S0oLTpSiwKUewHe9ICCz1BqiMNuDBj65wB98Smm05ZRVNthUUv/mpGJ
hNUE5G2MGrJ+FwZpx93ofwNZsQPt4Q1l4IN2KCC/9e0AvHwB9CHY688eJ0nYMlD21n49n3c6O3ri
QmBwnYe2jjJNklatfJ27CR6hIK7TjKGjocbxPAaeRNacV3L+nt9PDtIUto5a+493ZlkT2dK7w5KN
Yr6e0Hd9FxqI5h0m0toHogyQgH5AJ+a3rwdGkVBi3EdURQBDJfcff7jRUf2C3/3bKZM1vnlOsXPM
UkXQvpWBgoqsbTgM/WT3ive8cCW/TLv/A3mXwB9nusKmV/gjIAIjaipega5WrONbSW97Kg1dvJ8Q
a6IvSEuIeXNtmCCTDWTpp7b5buj5d8ME3Ifx2h9OCFf+3OaPBU51YKcUGzi3rX7lrFIaA+1M3nJX
TIGZOXOYT4Ftoc8J7YjsY7EHcHz80g+ExEGz+/F8kJogThp+689e2EG82ZIdv3PrGxBBoG6nYgFk
F8bJbLqWkp9e/G2DVF7DT+t7q7mkvD1DU0KAb+unT8l6pLMk9Jnwz1w9nAkxZY0m9Ky5t2AK+mQf
bitpCEFlNSY8zWtcH0gzRMCmTf8/zn+cuFkv7W0UamRgCx/Sef/S90umPoDiZIuglTEG8eFx5YCc
mt/+5mSmAk7TsrFvhVt7pZd9zm7XkrohQbMTaj5dIsPsRfHkxfvFew6dIqzHqaVrU7A+sD/QWuRi
ep7vNwWyzVWBFX4NF2rq4c7orcXBUl4sgOKCwgeuFP0DoBHj/Lt9JzkbUhxSPbg9WMD4vA8k28Lu
7gFv+0z/uFYvEezcZAVx57WoirBiaI/VDZulstFTZn2G+UXpLpP1VFvknBeKwk9ASGGLdFKaWSe+
IL2XpD/iB90KaxUQZ9KsuGU/2oYs+6JDmrGEQNfEd4qzUWZncC8hrtvc7KpW971yWgrDBQKO9hi4
X1QADE/WyymmBceQbHkx2NpwwMrDQzt8O4JEwTxXoLuIhTYc/3h0rHOrNvJstkMQCjQXVS6sGjfK
NhTJ5pPDR7UhYf+drbFWF3Yg1b1DHIA27+/aprCxFULnsipY5e3A1p9o8ZhXZdywB8eqyotvXaeD
Rf0KrcOqbeStPyJbsqbaverQ6YcEDRXi/d5H/7GsJlrR/VK4VwFwwH5TdVBt9x3ghppCyFLkpP9F
RTIyUNSxC7nONb1sl6i1XTMg1XPqDnWDnSaBIk/GrfvGWnBCgJIk77fjJZiS4SS7+/k1PkFVMsvM
qflRkBYMZIYIoEasvNQQwoWwyHyjb2S3tNaMPrKD4K+k35JY6WYRi8vIVheK1eM0+2RAedjgpsTG
DK51ehbxAFRT+5Fx2PbZ3PozM82EBycYldvn+GeD8UQnTALgY1FfOZKv3rwAJpeIJQTHfyOSqyyh
eSUh6DeXJaaMQYPEHz2ynXjaIr/D722pSff2hI+hqOFIjBwsNlJBywlPw4vwn/EV7OOqas6GcS8f
Cl90z78RHlNjvge1WF/wbl0/zIyGLQ15B4wAwG1JUShOfdAV+ezpbfMUXBJtawywmDTHujhG5XZT
S7SFnXKKM2bd/obDDeLpyp7xLPkY10G28gsPF/CDrw7AEhJ9KQ8eun1tJaxUQy4ZADOJaoMDc4vt
aJtbY1hC45aT5RWnezknyczCWAPg63eMdVU2zy+OIN3THm3j/fhikgKRIeUT0j3Ub9K7ptQYm6Zf
6IkeZc6kTDCHdTB3EV55yk0ktyL7lgR0PLT2na6zx4QU4qpMRvadXWgB4YtI95vZHiAVtTdlx5sK
NrG/lJcnfnJHN+EpvTColHSqqrDd6gaY0zX2VpjOZ+M1+UdncZrtV4oEq+6QVxfYXfLO7q+cjRkE
RjXZq3Y8DXMflmDjuiXpxrWx2O3Lxdo04eEnrbpPm8AV862njr89qcyLdNOgUXo+3RcuJege1z4i
s8WNSEnXkNtAgBxiTrU5I3DVLsNDtp0J5PgBuOgJD4+oOYrEN/chFqOHi4xTEkc2Tku3qTZgBYZJ
4a38fWtDor9fmwtEql+nzuY4ZUcu2APY1VwIKHdDbq+ojigmLfl5IcxPvD3Nl+NlirXFbTZJtw2f
dKNm1cPEVTkEEILB6MlVZFhRLls5lJ6P01e4ppGyodk1NJqyeGkrmna9kvfsAaiIwNqHi4QdrJYJ
I/QzGmEvjvFB0aAIL4nwNG3WIf21jA/ahzj9G6iicLyuBhb1y2zfSy7aapfhbRguIP+H4THNIZlp
k8c7SQNHR88RZ5zcj8nMi1ak6qxqCV7xTeDczQS72pfKB6PyPmnONdpdPpvlJj+L4EedKFFKgr0S
xPo4LkdqtWpp8Zq5SaMkMDxiLaQ2sfy4M7Db2QLly7Kxn+DfVuSFlPeEMYMJ+WVKWHBzguyT4F+L
yF2SF9y04pObAVa4eZ/xYhbpleRy/G6y2lC03IPChdh2T4Q1Zlraquq0sZqiL8tpQeqv0WjplWGY
h20lpJzXjPV+zfhTeN6B/EXmPm/QMXBF6qg+bLajzpnCIK86CCCUiBTr3cnFH5hZFYH+oQxTGLKu
OlOPKUmZiaqjWxEX9+rHoP8FBpZWUwyNP/PX0VKYf8Pow3NUTOlixBbX8hr4g6LnUTxpXEyUv9ee
NVsQfLgYmCVqjFr7U4Zo4wvjUr2IHsZfVe5xZon+57ej5q9GTSJn/5wK1+i3a/7fYlK1+SRTbEPJ
8xE19wpASese26nf0qnhBArSeZK0dvYP6YJhTUba2/FCPas1L8oOUG5PEPnDNnuyYN3GSE3UXC0S
IWV6FJaG0woHuxisMkhAwv1yTvLV0iSEV6+A01BXqXBXG6qMCzZrC8UEOWwXFi8XSyxJHSoRBfFb
gOH8kZjX/L5hAxf0FRg2RZif4HGEjQ7qwCDGFYt14mi0sbckA7lv/cEcs6SYJtLdqQ9GioBESaRJ
fPcz7hgiwC19d6+ThJU3D8vbLzRBeHaa7feJGs0yEm2S3UJvecX8Oln+kp+vl51vD8AmDayZXpov
f2yhvPV/YD5s/sW3fyifbk04i5PzRUqKUFJCKbtKcW16r+nbCJL0YbYXgfFl03lL2Sjo/0By8go3
k7NtvpEIf3jqC0lbxV+K5ZTYEt19qAr3MkyIrAi9D9OJD+f1vRntc+btHLtdBL2mXHUGZWeVBZ/e
+uLAtxI783ATaVllYBKWkuEZ+9AnMz34PE7T3Wr82mBvhDKdklVytAV+CGu5f97/COOu6GBaIdI9
uPz5iTdxRz9+gZeZaBCUQ23yKEGvevuTq0vOXgH2wdpCQohlApxGLTRUcEGUrybri6M3bopJKKSw
Nh05Gb57urT+fSj/v9FMnUfZ+atD3x+kUzeEdo+PAT7UK5S5BlVrCCgZVl7WN2K7TxpAv2E61aOM
pgDoIU1Lysf8ZesieYyw80hmoqlwodL0pZm5tT6AahlRH0O5BUG3oKgaPT+9yQrzDDaBLekmWfL5
FS6ZFMb2DtndxJNuvbvyyK8Lwg9tEMysvHWHRNHOXSwpMacJ/Z/FibNqcR6pY4Gz7U2FfcBvSXCQ
hrCxpSkWr99F7k8+tPiS1+S5C3JMnvNE6RmnGo/umSWQE4MbcY7wbZNCF1URG1cOULIO+5C8wwUN
LGCFcpgGKASI0o5b8VOai88XUMRKvNoXY8jwIaXFAIYykdJQaXVkqoJmUrjV7IHyW8vpt2qpqjCL
byEtLCxKe7e20Ye55Xu6/8m45J6ObXdYuUwRS/7wKIMwVK6oKjjIRDIMUgy2PM8GNu8hf71b4Ob9
J/bV5bjcQTc4VoAr4wz9yJlFJ4bJO2dxRVE1y13ptBlSd7Lrht8bMbY9ai7agxZKCnR89P3YtmYc
wth6FuHAs98tgAblrVrXpwzRW2KFYa9q3ATgl5CTtRf8j/SDtX5754/L6VWEmGJF76QUNvbPAoNc
NnSTWK/Ag86J+zGuXv9167pYXFLWOYhpir+BRiJux3HeVqwt/sp7HpZiudz4RPK0mJSgOF+TZ/Y0
unAMJtu0xEqxn1I0Xn/YsCkbVa2JZz18IXU1mYFGqoJO1q46/CxZ68HEWS8njZNXL8uhxObeBl+z
XNB7I9E+XilJTLdpQ9AyZw593Xys7yi4VFlfzk9TtSw61Ko3yR7fCYOt2VMuyUMeabD5xJI0nbG0
ZreJHB+egD0CQv/XS2XPkAE7Lj4r3oo2QhUKW5yh7jX6XEQhjoPtGrO+yAW9idyEJNO8DCGZEfpr
Q7aILe7YEQ6F+qv2et4XII4I7UOnz+NvBUE/CQztYxQy8KwN+FoDHbTj9DSj+A1P1zxSoL//Rlzd
wfgIPgmHmJWqsXuSA6Vo7x0s7W7bjW3zkoHQ3omYvy1muLqhyI4c74qC8TAMUnQ6FJ9q0vYp5nog
4yF4qIiRblFrjwd6J/xS5JjuYytEz/bK/9p7a8LvcxfHEY9IDPFMmgJqLSJk9moO467bMc+Oc9qR
P0t1SVux8Cd9XFygf84H4CGZyIl9qrSQCD08kNp+rgZbpS+t2YizJpWdSSgBmDZbjEBqvqejNMqa
v/QQEuFErmBQ4iZ3e+iAVhxNVcaO07vC82b4WsImVCCI3HC7sex661cjiyr9wWguxu/5d2CCQ4ra
2YZw7XlTbI0QaJKpcTC4X/IEaQN/Ruw+O8Y69JMr4KrP0tyVNMBXhfSf9/sCzSJ58lupM476dW5L
NFkzWIgPs5UFq1PTuVB+C8mt+mXd8GERVPx+o+kaZp+UhSOeMEBlpSxG6wZ49TUpDTEchC/fFj0M
UkznK0KMMNVF3JVQBAvOGIGKZEZpbxc6vQ4mThQyPatnwpsAO4a6XwSA2Jfg9ojg+lTvcTyo8wZ4
AzWVTEdyMpuXCh/6AX+hJgw6ePEXPeeAjnTXmMVe6zVnjPQbEJHmom2yAe6GQcFGmRXCq5pbZ8pA
+TfcXvfKru2vygL5VMOFchXt/nAcc3yhl/Ph5brsYMHIC8/EIwnPlcdUyQv82NdvXypEdZRf8Neo
Yrj5KbB+jTeSR1CtSwtg2TrV63UBNjgo0nfnqzMU8G/dGC58iiLjS3wAMudpBYhbBNNtZVai1HHV
6MJSYz6KyPKFPLoFCh0TsIf9LzVteCcRjC6AGhqSgHMKska9PH+LY0pGPtCiUp1UKIEuGxZdbaay
GgATCcdehripnSBFu60mh1ZG56yOiG1YNzJpSyTWZobtt4e13DY9IgbOX7zKrRKH90Sa0jRh7pt4
NFwPXnBvv2to3XYkfHduIju50F4tZFOVCnzBJMn0VQbEaaGBKIpipBdOEVoz62TJ2c8PULhVaXBS
7H4IOKkEQ//rLh9Zbr4oEkY91ihK23CJahs1BfEiiOXK7HRPUbehrHRPpKU6kuRFbdnSs5QW4Jwj
uIc5QFvbWd+JcrsrhFvUht95Uy+slCTEa/gtu+A3BGQKDeC6cv9e5bQZm6AyWawOP3VbYQG9OZcD
xCcSGslv2dxp9I+X++jpgiwDlH4GM03+VTTjoy6setKsIbEr67B0ERFIaDV78qE=
`pragma protect end_protected
