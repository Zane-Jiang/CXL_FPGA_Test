// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZnV/pzEMixNTN4EwWPIizf8PMjVIBUYkFUDSRd2kyTw5Mc2hct4ho+pPHWfI
OnOKlKKH3BroIWhTVTiFGPACD2vJNjKTAKlx2trU6l505t5VVlKpnlaSmPS2
u9fxn4uHcRWdy7blHRu3bZkL1ooLwXFChXb+bGL/UK3eLHzRi+0Px7n5dMnp
252kiQuguwYkC3+M0pW//yEk18UeCPVGM55YVq8XZDG5vL+cBEY7oyNAKxoW
fEKtZ/AyfcVO9GpE3NPH72uxGnyHyVQ89gO4NRoZFBacu9zDLXuL4YIKTUXl
dRYkM1XT0U2cnw1wZo86nozUYm6ZYGux/WkGiu77KQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TFehdaYB458nr4VPN3NrTdM7zsy1kekDNh5B16i6CekfkL6gtCHjtKYUKY0N
i6GoRr10OR6a0Nn2wZ+oKCzFfVWW7Fooh6D59JV6nK0BL/lByY5YbGr1g5LB
cLMSs5LeYe+0U+SiGbn8o/dt0QzUcskGWut+epOCUsy3UXyVs0fKM2aU4z6M
R+bvhrPqQK7r7C3B4OnamQIaIjM43XBiOjNg0HfLG/t0250wNBuEiqH/nyim
IkgBNouHyjH3+36B78BM3Jr5Qv+6wiXpQBStcNheAWaLjkmojPuWyGtg0Gki
/asp7VaMbXsmA9h7vWVFB42KQ9Wuy2CkuEcGVaB99A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pRUnHoDrC7t6F0WYgLBMNlFEJoBaG4Wm1LzkmgoBMl2NriiuyF7OtAjN2TkD
aDmJPZbx9P5hRrfgXO6/wM8SCsDbpAyFYF1gbiiLJjELF0cLR6NywQXhy8a3
S93/uxVM3+1c3XCwPOxrbt8wJK33/t7ybdlu0w68SiFgSCjCu6IA6XpVCM+a
ZdKxElUfW7gutDbfAbl6AnFT5PW/dZ3DYEl3gJdAjOyaGu6EF7IBUSvr+SEF
VmYyWY529iQJqlVBdjBwl/pL1WfFkEQ8+2xcar3CNExLBqiWTFqfE6Edg1oR
xzMpnPQ6+3gecZZzDcN+e84vuE0b2BmEL6nEKNgFTw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MsfQgqHBrARq4CHOjsBpOSC/A0DYssfbn+orbqE8KaiqkhVq+j8ISXSnxyto
k//4/mhH7TiyOVGMZJ/uWoAWqmMXf2RPpp6zQsbIiENlkN0JMahMK1cOPrx/
EWJG4IXXtaq1ftjfXa7EyN35jLOz2ET3WHkXoDoVEuE/bx65CKQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
l+/PE64m/7uoLewgDlrHjbfa01fyn/f+krNTk5vkb7K4A6MuV+3xBvN/Rbh9
ss9iWF+RH7OsdsyxQG1BiG2g7XBKdufdUabGawpKkpK+pIwxzWQ+LPsz6kZ/
W3tFo5uW9Pjv+5e3gZM7nyosAhlpFTXKhFaygp5msJqeOb1X5urwWCQ5TX6v
1qb2Bib/rDmTx0AgiddUTjjuqKnggjzaypdikcrDMiw8FtdY90cmM/p/N33x
DZ+35Bgy+Ar/jEiMpGrrO4lcEVgslRsaKthqksbDrtWtCyDOMNWkNuF3/F/O
YCQrc3LTQyY4FSAloUyHwB4jAEE0uYPfgMVUTyX6RAxi9kPtXTrwn+xQxylO
r4k7d253Tn/AMUnbbboo1VVeE9STMBcuVLx6nBp1QrSQAGevYCsNtSrVNNzJ
TRMLi97F/8528+on1tefRpxq7kPbVYMmHRmCWgn5mJQMNmYXqcMwR0YMTlPg
M3OxGtaUzLG445r2gsJCXKLvlIOnfADz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
un1JwatZ0TvJLJBp7LFc6Bhv9zG+IVcoCcfbZOcUC5PyJUchedjXJq0OUd/n
/BHnIJe0BZmPQwPR11+5xswVfQ9mqA9nDlef4JbXt/DlPoA+UENQVYxZA8IN
1SZvq2ovuEjEIfqp764O8lSGfwBOkoFEUuPtkTFLx+RjaMj5AOw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CbWr3AJBvRJxTGcS43u1ZCuzVZ+y/dWg4lIOh7ebEVDjOWQFPK5DDDquKA4e
PfO85zbE4wzysawj2ObMYNYvgetIu99xo1GXGzsS4aBjAJejYBdC3y3ps4FO
JMMnT4zgGkyvOKtaZXaKCMEgX0KtldvD/0hRJrBPLlys++HoWao=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12528)
`pragma protect data_block
gnHioLon+XrfWxR+Zr1Ap/x1J3DlDWFzglylvXTyqd37K39WlwG3kl1pSTA2
CwVxXyZdXcgURtLqGi4Fyf6TQEgDC30sbdmDHLOUBBJCL7X9xUX+ukfdKRbU
BkcvFOF8qMaLfRmJe3+mroY2ZmpdOOFSH6MyY2Yt4h9hPmGht7LEnj0oa2iw
lhpjlJhPgwfjcVN8LJ34ZgEcaxdOaKU9A3RBT8VkoIfhhIm87eo4hx0MisQu
m6BHe5XVjCjyYJU2MvN1Hc9XpuYuze6xmJPPZCmasVH+7HXh5KoIvr6+caKy
o8Oef5DE3mFbV/hLZQjAm6RwaWGqMXDfhN/tm6OmtURC/iibvWkcepE8SzfR
dsMEudOniEPHI580gb1rcj2NX/NzFMXJ0OQarBjvzzaITyvObDzlWhEWBpOX
8FFIWIz3oVMTdQyqyyU5G5Q+LiWLO0my4yOzRjwGU1s76jXsorwnpWO17oz5
ljk6x6AkGaK+g/MPBAV4JaAp2tQhkjWzvarOJz+fuuurM6JEV9DBgD5tFGgq
vLAoFrgPRl/3ea41YYK0HONFbh6O9GAqtJqiMZSe4MxtLKju4w+gi5pzcFGe
HB6ThcPcoZkakevQJUliH90jaimGyzRpkdIsYMsI3oQF9bkd/je9VNJoCaQn
a2kAY6PCNtTL6pQ5awuFc2jDp5f6SpVV8EDIlOSJRtugt1lGR4k7R1SuKJ3v
Yy0TNpLSN/RlNofUQwz0O1YRkLIhCYEo6KOzGmBBptJ9mlGVIj4vVh79+i0m
2uKUDgNzqSHgduCJ0vCXyo7SJv3X3jsExagbgfUUidp0XwVmam3ksJwKs/pP
D7/MMseVkS29yX2dWWP9xAvrzRzEV0/O26UDOiZOaqMKTsbW7OcBb0I8/L4J
X0SnAKc/N89PklFR5bSFVv6OwVIQoDUzbQpmpCe8SV/TPATnjWI5kkdwCLck
PHXXe9Ndd8dJ/e37EnG0dqLscTGff46RNsRjZpPPnAMBOyaEJTHl1s6eVF7H
0smMsJGl2eDRgiUNYEqlnH2zHDLZiiIiFzmpxggZPaTCKR9eLiL8fbCgFlXo
oO0M0MY/stKo9wIdLi/qUfwvGUBj7qqhQx70UrVfmuji/I35TWxm5qpeajSx
DIiEmzfx403A1MudYxmQs3J13XNYahI/OaSR0HI5Z8tcgCcx1Kqdqp4fDy5H
NOYIjH5KXTKJD1UdQOAQROf5ctJD0+Z9szAvFMG22p9eu3j938JxvlOWWfMn
gcklZvPh3Tu9waU0W0GDciPyWVlmTIpQSGnM+8htE6uFifIxwkyxZwowQxmJ
Ek3KK/aZ5TJAeZd7gI24WZ2ovmRQOJjpxpYnejodVyrp5fHLe6vahh93T81e
XxQqaMWe3BH5MvF2NKFlXwUNYtYASgcWLgXUFzCtWkdfDwmBZVjRRL1Pl1vt
SvEjHLexKwdqkRdfyphBcemGopbB7YjebAQLQVMNwQxvoKbqQtKV763Ztg1J
AFJD43Ak0pJDcxJNjobSOzFauNWZ0w5xtWH4gMUjB0QUgFsDrWanuLt3NRXB
LBQvVqWmzwx9F9rIcTgwItzBQ1NnTmfqj1mFkMCb66mJKCqy++sSkSO1diMY
W0yeAlG4vQNoqWST5J4xy7KNpkesZPWthYKDNpLY4FLDEVOT4j1dtJd8Cfj4
dTDAXXK/NDoZhyRMpx8T4hhLJpSrsWkSFu8IChL66Q6MDFU0dhrCKIeqRKHL
uWHjJWbK0wHHsTqpaYSR5Y3QmuG2BAmrR7PIAgm7XG9fvKtLZrqzkvl79My8
ymmB7jc1x2Oc7RZ0bdnTyXuB3LIndb+ps9Yjf7RN9P7fn0qSSFWzq1z9+q8E
p9YvdW3IUVXbZlNKBrk8LABGvoxU2la0irvDQCQyvQJyntSDFb55DClFdUVK
JSga44svFWOUCAu0X8i+pNjivUs7bLY8S0bEkgR/VaFJRRp5DRXBKTgRk3QY
XwDbAd5aeCeHJCD9se73mHc9fhSDMou36ztZiTKvLpeAdKr33XXRyNoQuzk2
IMNSJ9LaH5wOdt0KqBn4Bz1MNPallkxtfgmEg1DUZWbjLeWAPZ6q5EizhOc3
1qEXaxUTUckRrBCFDtL1ryROk3edYgQ+vv01ycGmQ2bnbIb3WECDv/PKU0kL
/QQR7i9zVwZgAUrL0Ax57YR5aQbRIaT3nzBmRtQdO46ZNNWy1cHautYPrepz
BtOeIjv4nmAFeVg4be6rasgj6MD9V6thCGlm+yD2uox+kzdOoDbJviey4/Jw
zmEgg4Nu0UbkI+ws7Sd4K/8m0VO2St3MRGiu7BPxAg3xoF6rqn8hmwyYasxP
tzuFzyFW9hpRy5n0qkn9Vs8IE7qpB8M8dSm3ioY3FI3me8Rwy0NdsHsbDKOp
C5t/Zl7xPsBx1ezIS2XMs93FafwHU1PP7UjtiF3yQzJ+iOpQn6jL+e+kTn5O
Lm3BsN5p9u/2pwxkT1ldt9kuwRR66yP4YfT/+GLL57URKn9kbkIFVq6sShfh
bEur961PI8piWSnWg7bBS1FwbbNBB4b6a/fjkUA3mEVZRbIYXLIESYqwKkFU
QD4U3+ocfXd1EVRahk6ckkJAbbhRka2acf74SW5e4VVBcJR0bE78Lf0KBgsC
n/V1UHmCmL8MRGYno2OMn7eDTm7p7uPFSGvCNWTJcstPU5Gwwxr4ldNS+Kdl
821gSYHCY6J/4NLIpwTy6UJ3I/K7u2UCd+RIydrh2zYX9rQaajS8eGPIbUrI
dJmSFmn14yw4nYYIaTJSSnNDKogfiaMAU5cZoCsit8QsXp4I9klmMCyJBATC
KbTc5NjEuNN2PCq6xZr17KayP3F2CRo4p8ZpC8BWFej0wxNGw5jgBnjoSkZn
m3pE70DoCEBjY9UentULHUPaHIIsJs0LkATAxrcaQQ2GnxwcdVI8tnTrABKX
tRmMmTmy7g91CL5wWKOR/V3XkmbhaADFqJ34KRCe8qyHIhgmYhVbbfCYHv8H
1jEgcbVMSlTZksK19TwmhLsfSOeJSEN1L20f6fT3i+qof8F85xN37E9g1Hv0
yQSA4V4Mrub7JdxJAzEWOKnczyUWRhcDduTX/h4q7zMAK2aE6d2ZgO8DTlEg
ItqroqmK+ZTmYS1PrKIVLh1SSfJtvZ97272FdE37bET7nnLGn2vtYMLXS+T6
akqyoYL2mFrJGA8EMgP49MV+Vgwz5ZKoe7LCxgoMjs9dJU2PyqdrDgQT3Wb3
0ptkUtvEaScpGJTHQxXkXeRayyRu3u+LTnpSH3K2R115WFIFRQfmyzGX+7cs
59NFgU2dpL5c5PJ6pXSRAfC5K7hcEBuk+VLH0twqCyoAsSnndCeGnHWoXpDL
HKlreH5VjyMUg5hD8hcRW1drIeV5KgHFuOjKedxaS/G9sQ2sobV62mDyomJi
VKMYykk5hDWpNao3p3bLFWj4x/1v18NuPRLzdtlkPUkhF0RJe7k00BSEuO7d
NlN9EQHnTiM4yikAeCY/By9yUFXf9bKs8ewAgFgN+y/oJBFHEE/AtWHFv6uv
cfw7r785G/G0NXXq2kZvms2SrOZ/Kwxa/dfxupuZt5eP//C4JC9g6XUsjFLr
VpOu6+yqoyrhvAfC+ST6RODOL16IjvoINIsbsoaXnK4q8/vuRVayOq/DxOdW
R/iQaw45kf7JN5xMlqUo6RfCqS5ZYOn6MfIV06eyR4HC4az6wyjsWDEOL7Zy
YkS8SzCGjV1quTGEUUFkRLm4FhP7FDMFL8AsOXjg3WfDIaKdQ1HXAaSDAwYj
Ax+LxRzn8ZwNZVpaAFM262X0hSz5x+bJV5SkcG/WK3G2Oxc85uPBs9HzuPm2
DbAp3VG8PMBsN5c77Sdq7pU6A0Hs4YQ1q8SW5QV71IsdEDRln0nCj19W/uou
o4u28N1ihPrn4pAsSjONSlsDQCnZ7ssQleMQ39cGdOZENWhTXX46g8wXNEC1
gEytPCaAPwfevwSdzhyYPVSIct1QjQ1Si2YvS4GJ5ZSOZOUVlPM2kXAM7ZIs
EXw9LYSuGqeeLxycShgtnP5V3SWES/ynlDpFoX5An6iiinjxAMurDA1nzVm2
SqkJDxJ8hWFsUML+aT7c/rYOLCc0be+wohvSQi/doZG0qxCo07Gqyb6weShV
TEE+VxrEAUqTtnP93uQSoTV3cJrXeYcwA606nOHGELygNl9UlgmDwEcKDXoa
nWIFO8q7hQ/g19Fn7EfxMOwraHVrat1gbeHedgTC2JEp2BkFX6Mb0LwymXKe
WDL9ujOSruCw1ufeiKw9jssLSBw6Gw+v4J8DSBc4VhGr0QQn3jDxmoQHLspL
GDuWcTmW3Xkq4Fnh9/rpjnSg5ibWFClRYRHPZi4gBSLHoA9+yb8sdoaTk4Y3
PxoLi29ThC8v3Fi5SvPSWdsxX1qdN+INHPwgqmxyhz1+qo7b6JtiDsmVIe7n
xngyvPzBKCNMJqRBnq8Utw+6skRyDxQ1FSXJmOyNoLHsx0zxYSVCqBuJQgxc
0gweSfg0PJhxeFenzo+Ms6EY/SW6caiAij/ZvekCax0Egy3kFAE+Qr4hZHlW
nQKAdUwvGdsXpVwa+6g8cVUcTqrbYhciiL5CSyZqnEwNdJyx2IPCJmfM6f73
Gc0ofCuODEkz9WeYfQEft0AgS5bjBgfv3FwHK923irXNcohGDbldU7DIw3vg
1MqN8lxF3UGHZPZXnfGRG8GIPoqATxjbhr54TLrwScxrQqO9KABprJ/Ap/23
R6T6zI8cmU+QvY4ysuZ15KdfK8rrmFOCFE90SFfMpNAid/dXtXl9ElDV+f5m
sRwhvmOi4QHGAGbl2KHU/0L4OTNECoHt2dX5aamFxrO0ggVTnCYehsXMWx4E
sBwOz6uLfbVs614jhQLfq6pAwXWT1PdSqkZ3h4/RO5/6URDlhrKLP+38y5Wu
laVlnNyWK1Owpp+JgJ6Yo9fa4vV+aLh8kvbN0BAZA/I1NEL03k09S58JXlT8
8RXI9f1/TRhp+pdkD0b9lJ2wfDD16g7UAUyGCxaSfoKuC4dCyIWWD7uGaiAY
Vis1BojKDV/NPIaSqq88iE7x/3iyws6iEMMG45AjuChnl28OXCtz8iP2f5LX
D0nmRQpzZCaKCI4YtmcQWC8Llm+vQpSms8wiVtigSnK7gT63b8sMEB0n7j2C
oUqU1GLIdg5tgZK+6PsLw2VebCj39xMHv8IA98SGd2mUKTJ+BXa0/dMMUv6p
irewOziYWAW9ZF+uO8gyb3ieU5p+2QpCYbkdM/YdPech4hK6P1Dd6mmuhDxy
r1hytZG+iXOTF3RlNVPvMX7iKc4yvMmD7+uxjYaWwyUk2E+FmuYFnqxTrv9w
jLwmfoA23FkTAZVYEyLPS04dG0/FIaJoWPdo/DU4tjmESIzSM4DqVcrkWJTW
WPvOcokcbBKEBAfpJIXCarH+upLo0ljr9TVZjXOvKJ9kSpeg+zFAdmWPd4Xr
uOi9ldnBps9r/J8DFYf9iwqlLFTa/4CvUb3Q76oaaN3Iiiw3zwLUsGP6etSD
xq8KFxLgQLjOhpM85PGIOUXK+0h2lK5JSK98OJ4IJU2HGIzTB05z2OTRB0SR
42B9nwPu/bAdP8OfN1MySvMyFfA55bUoHQ175DPZuTgBVPJeiHvXaN+gB1ye
5FcQFVjUS4OfsbtbhVsYo92SW/mb5Dy1uXTX77ZKt3r7p8RhaWW2kHaVb/i3
r2cb+POgYiu+OyKGGN5zw5QBVWzJL/FltOrL2m8yXe6oXkkFLC6GNRR+ocsq
+KePWzd2DnYD7nUwHnPCNDJF8ra/pu73OxLpi5Q+/8faGA12p/6CM9pHW3Nx
cnv7i+kmO+c+NTviYCEDasJ9BWUScGUtu0BImiL8PHoNpJE3eLup1L0sqDCR
6/U8R4AG+Th6umZ6iV2I0+dYuTRxfti6wa/whZ/s3/97BRu4ehqNbTfOPGCN
7oXRUr/7/DcQQNYI2tZcKOIxuA0Mc2t5BIsxeWjwVTPmzgL0Xdwu+gvnigan
BhkAwdL7ZhCuJqMMYgakfMciFfzJF5SlPMYsFpsugu0uS8LGeBJyqBOuNN7P
h5Fg8ZUpSQqrz6CnfprADLR2I01lVqtVrFax1FxogLcxwsTpO1Z+62zKdQy+
a6DHrQZALO03NPAw2Og4iyGu2r1uTbmLxibTjo4SaO4u5TUUWMhXbRmU4jkw
VQT7E5mmTjnZfnvSzSOlUaQpNnHB/Y7kqOtQNNHINNSv4ovCmKDUw7HoAg4K
KiFKicng3omzC02Y41XM1SGzGXJbfMamnCYZ2oz5xl9S1lmJVFLAk2Sbj/9c
MTSy217mmI7TJDp4fxojxBP4O5ZicQ+0k5UvaympN4vA9Y46yb5w8+uvvDBp
c6hxLf3cbjfSPTG+BIa5Ldez5accIN6mW4mDu+WEm/77oboJ6ZsOlFrrCAPM
mxR1PLQHkR5/GCVR0Z0LYfjQz10cc/HsSPKqWeVcv1DqvfJ24NS8JB9RHY8i
kFilpX2InvZWqZRfpikCQLXWeRYhZ3GHgQwk4+CgkAUMkMS/CrUk4qmJ8p9v
V+rduTaGDVq85YCHVGB7/2M6cYCQHj11D0gPK5dSqcl3BWFOSLTka81G9/dK
yGkOGB1npVXo/+t0M7jCDEumMrQ9eHtWc/rWMZlfHvRwYbztgjJVYWYx9aWk
oOY9CBy4nsTksw+zefHatCGjqkucMzCqe+NJwL3dzxc1jvi+BE4RwYwS/2ex
znW+fdt6zEJuouiEIND3hxFtZpgovtynUDOYgC6WVHU9iJUIhnUheYr76HVM
4jeXJXQun8jlG35Wh/rAFPn/rNahewuGXREbmVvzWysotfbQLZO7+Ym0Djyv
8V+Wv+ubf0eEOjDkupDew6LzGfXWRlLPJuQqm6dy1Bvta+MSUtHhTd7cxHUe
FW4cUqF7r4gNcfNbOOybDsendqZojes1VtWswXfk0bQTsixXi8wR+mYEp854
mQX6EdGFuR2UnGGHYsWyxFLWd29XcrL3eB6ssblFco/jOTzoGZEpOlW2N889
JwEs+RVuyrZ7vMxcoW84KNYGNmts1FQO4uN3n06D3N01wpAueOvdrDnOenmf
fteE5tCbz5QbUHNtUM5fT9IVxoM0kVkw8uq3QODB0xwwYsRJKp13cmq8H8iP
VS5Qyp4H+IDWYZb20DOPl9U0i2tsNLV0M1R4PCsUeIDcD0VhXq/XWakbUnwn
v0fe5n/ERn+FTuzRwCJihAAD7CWarUDcVSRuJlxHl73WiE+QHPrtEtd7X9Q5
hPuQ7bS4w8ybARZ6ooRxnLfAe39cAq2y43fP7QZ/OHFnMRsp7Xkybb37rte9
4m5XucDI+wnoSGbNHUaZumMJ1AjiZWZwmhpqwG3NGOhpbC0DB31tu7U1YjgE
mg0eA3pQ04yRGkQvcAwC7pE0gjk3/JHduvu3XMkM5EQkX7ilrreY7muLaRdt
fWzIJEAiSRvsoVP4R1BIOPF7SUKXs09z7l5PJ3J9wNq2qqKGCe/wGkNmyIUC
w2w46rn+Iu5+R9zH0bHj4Uqlg2xdm9Vzw2dB6r4GFosCKgq1oDS9DNh00jTI
kj2nPxhPH0zpOFbEGegFZjBqyuiMhwop0bYwIBYa5grSaC9lQdbDyZFXQUa1
7o+r8rsTBuGaKhDjygqrNYQUz0pShMf1wfJ12O6P3rIYcyJHVv452lBJl5CE
r4gbQH9R/ChSo+qxQ6CyfHTF8o4ZxqqURtuGB5a/OzlxLYHauOoNDDGovNOH
hCIsQE6znjbPClzYhfvCaIiFT5gdtkCcq1a8p4jl9Tv+OBWJ3F3FPjiLhPVS
9xnr50llF1wJJLE8XklgSgJqWX80rmCHKddR0keOK/1MA02IaCyOSUdkfYYi
ildhlJOsGWmjTG0pM3EqlaNyHgxiYH8l8bTrpUVNASshjT0NzR7q4Nd0jRjs
QaaRBMlwdx4q4Nka63g0HGvQOJqUd1a8/ueNL40y4QgetfJmRz/XJtgNGriR
JRwjkPCFbVm0/LDSjFHHF/IFEE77/f27/UpXHbZNN7DDvNSMUREfZVqjITuw
9gCEjOiRNUD2fMxO0SjO+qCZxn5v9ATROXuCWNiLo3MLHL19h9AfsUc+zJ8r
/kKsqBHsLGByedGuODy1L2EmNnOtj7oXLW3oAUhhkm1Cx9XWcSHrfyojV6zI
BWicp1HknKoQj9Ki2xiQ/sCJuMZTCytRQYG6uZEiM+9POQJrkVzzwbtcev2U
fwn/GtOZ08stZWjo4+3lx0TT/mkKVJ7fJIDeBLKvKVCamWa88BGOcq35zJSr
k8d02dWCNPZscrbtX0TCXrqv9+8EZJn5tQKyn4/LuO/eJW8ejYSU7dchjsyf
VdIEc4pf7+7KaOxKahK8u4Yf3CSIw25jvQ1M4lqmTH8Tsd8ezka39xn1P1Ga
5PSR1Z2nYueJ1juhN8CNv/sZzX4ez0657juzPH6uzIFilS0WtV0ao6pw5j34
sqVtTtQ1d8p2xzRMlOdn+GHgV89dHLa//wFINA3QzAGaoR+NpyNoE/Md5DnH
xsNWT1Shxv1kuwUCjEC1ToU1Y8N1x3ALzmGk/c3T5KwQnVlhmuP1qL98dwDh
+8I+sFlnTluQcfcBnfTlMrndeRFQbTfniUoGzrSa97BuwfySvrt6Mh913Aly
ZWrKJ1ZWBtx/Rs0h+fH+vLHXGq4HsBefu+lqXLqFvsYppoGN/1Lo63dY2n51
7bEu1VyEQl2FoVnNR+JvSWCo05C2ZlDyeUmjk7gQyyBiUgKd5Xal1l2pX4On
UWkprCEP0UUHC3R+aCO48G+opnApiwoDN4M9hcckwnNAxz9va4xgSMoYQruB
3bQpueCCgMNk2uHhuLgngTCzM72RpCHdfDcfPH0gJocA5jp6FL2GFHp8uNl4
KZvYIz3r0/4btD2Zyu2OZPxX5eYOgbzReBRERoOglY0xZssiyumKVL6TveY5
3HJXOiO5kNyRlXU+kf6MF0wuUxC5EA1BCsw+IgqyPipSM+25rujR/JeqrfIN
3NuR1OPDqmd8PN1jJWxi/49KUmZMQHjELfny+9ixv3LsAOoi5V5bqwcis0dE
ZM/33skkwaUTbWsJR4Eeb5RqxLtAWkOcYCejAz7fOobXsQPLXevdXq4iTgxm
5dMjLVTsqhy3RqYjnGtmS3Ksz8hw8QEBECFVTskP5tWccwoNLe3lvGoxMDV/
zKvcMdl0/EMiLmdw1YRdk/j0eQIbSrxdQiiUn9Hcfh2/DVX2S7MLRR+TE3l2
6tSmTm5ZetqrZ9/X8SpAyTrG2nF6G0zstNoMw1MsD/E0/qpwALsUGmfSDg0Z
ls0T1ug1vJs58jexapAgJaWoUjjYP8YZXt7Rq+BXAl5cln2QCIUNZ/3Y6bWH
N21U0tEV/u6eRZ2fnu/xzizN17OBILjw7rves1qbq0dzAYbwpXyuJXJF6GCJ
VMRVEa7ZUPQlSbVJ6ujWKZ5EkNvPwNiIxmjuFbWconMxZIeGGaOwdT9DU0LF
OKyFR0SXzbt+JczhnET3llt6zGAKTB2l38FALjUug5csfOROVlvHwBdEPjfT
/NKrtLyh8SM8gW9elPwnv5gv7ZjxtP8B7V7m8jREXtdd0kmt8DU0/7JskXpJ
ROnh56YBtUdt1Y5k9fUFdIKq96UUgaeNBNYzbx20uopZQ7jj+6Tj9yQN+Oeo
f8YKRUU41kXGUHzpY0Rirr9PxwfMwW8ZFOdqGZCO4nJ7bkCDR1AjUp9fEiWC
SL8XrK6T1fsqVqALNZsu0m5fURQC10hN7zMKOAAEY25Qqh/vXJelsZh4EBwi
Gpvw6ZhdFuDk6qZm1qAhdGDcFv9GNKZTB1uze0fLO7vfd40H4pTsMFw6ZBj+
+RJgpapS9HRl8H4oiDByE1SdQEFFIZXYTZ3JRjdnhiKPSjz1kUcFNvR8gK37
A2p7NQXmCYyq7R8lX/fpnCgwidGNADPO7Zi+FMEASKlI3Rlji/zpLKE/hZ5s
loG4hFCZrH6MOtaA3DJqnW7tqrxRRZnMx88y/oyGNq8PONmU46lIwj4BCDjL
URBB5kFAMV6zF9XN4i342KKvHSKpGsjLEVR6qWisuPLB7Qtg8tqwgwcGJ+q1
7RM6LN3JAofCchSgBCURembhRR7cNV6nOmOZo/X8lraSIVhsrPgVvRklLdiv
5V2klXTPWa7C0YMB00Y2Cn2pGeMMdZvlecWf4q6+c1OwY65VY7Uu/FeYAozQ
/5HeL1d/4aY6qnBAgRn5s77W7todKNcA5rzTh3DPMGGJKDA8t6yvve+ShFXT
ZtzwYZ5tGCEvwDfF4l/yHf/S4FykqWgxetSFbx47wdS8EF1zfKJBffCTdzka
Xh1srxQzTbPL0puPATItgSE1sNAFs6eXyyrCo4HJjrGW3MpMF5GnmJx3NsQP
jJXLwHY2tc9k6OdUTfdmUy7l5TwKQSFS/FgtMZkCltJsDi2xujh03NBNYtv7
9k4PRk3qK+U7tfAFHfr3I0TL2N8ioaKPDqi+1eYXlOjCGEHALr1FzFLiNDR4
WD7+BGZsGHkt21gdRHhRQu8mCQ0ux8wGxYVoJtiKw9lLH3AFVEzscneXZJaV
RGNw767ktGiuNi5uLuRoo7PIevYNVaBGgbgtWlUn4O3w3poVZ0hO3P2ueWjT
JrNjExj0hZJqjV0s3y3J5+SeLRVSCIyRq9ytUe3QXLZ4L6GguTv1tSyluLWU
AZKDWCcJhQmcj4iAlt7QpU6Dj5aXiJPoxAH/vPGAXXHowPUee2v2lJaZYV0t
iPQQjRpjhHLCTyXCj8tFA3VFpPTC1cIQY/JpvpxbhAxvTQH8C9DfSForl2tr
P3QQ6yuJuu46s+RxCbbMCc0MKZqsAz0EwIaoBmLRe0Kza3yGvszMdAK1sp7U
2DSdEq8+RPLfVvZHYJ2BJ+LJxDsbNNLh+yGtPqPANH9ngDR3zyAgfENiRzZj
e3V3rc3dWf8oEoi9qsXQtYOnJQB/ieKNyg2PAFmf6Zc/9OXEIfORxj7UqVCx
hAL+Bt+kCCovhHmiF/aUcgj9gg3luir7wBjlq5uGz/elSmfcxBOjwm3ulOzm
n3Y8PNVodCTA/1Pq4VvJViCkx48UEFD3Yv/oM+FloTrWQjTvyGkZJvkpghrr
/dxC3MckDZ89F+Pp1o5vMKOWc2DaQoA79c3bbm70JmGw8yYdTpcfDvFIBJG2
1Y2RQzh1SOOPeqthvYC/3bg1guPTmNCb6+WCW5o7IqFWwTBYwYcf32ss111w
RhjJNv8+s5bZA3zpODQoWEwAY0a1SGk4aUbWMeQwDeqD8818EFm3p5NAX3pe
RhyiscaAfMd5y/U4cchtef8r9r7VZ/YPaw/pnTV9nTpSNdw5iEgSIV+98BYS
B4rLTFkU3+d22Ma13v5Yr0D4dtLezkNR78ZO/zb0lNcFBBc928RdOJ8m9vHj
chzTazZoUWc1xodlDxk/CNGc0Zvb1vx6cWCTbDQSnrIn78KvwybCC5XlpPE7
DVkYcl20lKq81ciI9mncXjXXPRU/rPzia0XIarj+AcxAUritrb6xjmU0ZNtg
s6DdyfEMX6bfFevtZlbaFVCywj5IXN2GzqPfvvke4PQaTqCh0Ee7uEKYISzI
NUzSP8aZ5MWf1q+oyLzf/EpEAtLYspQvywXi8X8nGsE+fCectscYR7lN1AUb
5CX/u98AJb8YedXGxqZflMovsg3MN+n1PThcbw1d/TM1AzZYd6eEgLbYX4Qz
IU5XKNpL+wz27F77MVCdgRrvtkKd0Ali51ueAH3upb7bMP5fDWLz9mOyzTIZ
oVuWwPWueUQkJWENMr+J7NDthOukKndr37EmhLFqWR+RwzYyVNTKeyJWrurH
W7ErllRXMKXx7TkAFVObLRfnyrMHIu/6IdLKv/2NT6ynSKILc+FZDpa1163c
V4M7FLrl1VYDCurUed8dJt/9WKbRR4Gb9rIamZiFfqVOOefklonEbqNd/Kgc
j0oT49fsP9K2lIGTG8VnL+0m7dkOmqBQdKihch7nIEnpHW6xYhSJZhKpOH/H
tEb1XAYYiHGzeuY2ryQuBFomgJLdb4NSF0/1KgHvOeJygKGtWqTnEqeG+i5S
LQ1PsSMFztJN8Kkz7Hui+LI23hM5QveTqPcMh9GTNu5RKrXx4izawDZwOPIT
PDDzAbHb3LqXqmSTeFfsVi6jmYDB/Ht33v4Qsn0lOIrhgAnuZ9Ne7D8gdhid
OPBQhjAm1643mgmtipTVV5LrsqfSXyzLWIi+aQgdmqxZrYXMtDyQsdsp1hvJ
ReGKaPsrP2dOdW2gJEagJTW42LSLqsTzyxJWawIItu8348mbJ28j5uFzpFxH
VWVV2RuxFSH/w1kWNsVXnmACy4jOX3TAm/1OC81K8pCo/FzRQIzO8zvWbrkg
10r8EuXadfj8Dd8/8Cl1gH/gpgaX6EiGEwztZ+J/9IC7FsA48L44ERdwxwwc
CoKJxF/camlqOBkfGXNRFZ66k/BwkFz8zoRC4RtyHfX/9+Sj2/y3WAwMtg5i
NDMExBKn3W1oIcA/Q1Blx/SzcqjNVErhmdaAc23YNYW3nHn4AKIlQDrne7O/
939pfEjqW2swPfE/+t/i0x4J4OjoG+Ipd7PDvB+D+MvafIGu5v9xUHsGEiYf
cT9OpjSj39qY3Y8/2ZZ9HRnSNfOJ8QvKp1540b4J+WmwULy1Q+IAvsXWzIif
22lHRPfFmAP6bGHU7stKFq+bbZAnpeHu8z7nJ7SorkcZCQ1aHxeo6zADtTYp
kJhNl+JKEzjNraS5wzjATm+f/Jtt+nM8rtvIZGd5RXnr+Lh0X2osGLSjbIok
LTlRp8TCA0AAoCu3JtA90k0jmGzZYegrtCeaVjAcp5JQuwdyOfNQ0DRuHyxD
J6aQhY6tlsgfwr9ylG7wXWK3Rk4qzQtZ3fMopB3KVNOWWFJ8LwSYo+baFPjB
zJYTmh5ZSl+nt0WiWVhymArsI80u4L6BwZhjwnQRkHDM4/7J3j2r5JabuJnj
pwZoU3kbOIjbCMZSYbMvothJqDf64qJT8FxEjeyxFlOu0z3t/SVIJC7wmdBx
nYA2jZXnIQg5zSGtVIBPI33qabWA6mUO+ABguk4ODb4+jSsDlwXKYjJ1s0I+
Tr4c06hSE+UxK4Ls2YoAe1wmu4J5X3+Bz8pPJANO4PRsPn03MiRH2foVfuom
ALr2FehQ+zVJ5GeneHGn86XPr/gQjhLcpnQAH2X6E2OS+cVkyBntQYCvZwJy
2ZV/25cgXdIUW21g6U+HMuaeF8phFiDKUXNRo3eI2UKKXEoJQPdIbPkEvvq3
0jR6wotGAFjY+kll4ANY3PDhZkFFSfL4mBBAmwiQWSV8A5ugM28msroJM77W
Hz5SYiPH3+4kT8VNOa6qd2/VxYU9uwnRbEgjAKygedxSRqn1yFAMiXwW+fqz
Pbp0kcPhnSdjzuG4ljbBrNncIyvn595b+ftQjWtdHr4KZoP5KpAD6uj0x9Ho
0Za4N/8p9BGVVM4Uzi1WpVNy57v3aY99Th/9qiUOCbXV49K0nFF0ufKjWSYx
IRHnDTrylnWQscknKi4TvIILvthz/1bCM/LIRfRNmPSeXgO3Mz8rGVhi+cTK
Zz5QoUdBBIhQiXpWNZrI6PLyKg5a7P7ZEkxE5dn3iryzZevrUsLaISY3ZbB1
07oEwvDWdjoIjc/GqipF2bOCN7cvfe+c7ngKE5hN1Tj5X1TfG3Kc8M41L8Zu
8YTCOZ+4FAR9Ytor1y5O6yrlvQBBRQnHMAnXlaXvcPB6FQFYlt6kaJvRjZ6R
nXL18ih4JD0NUHOuQrNUVVa+E0IT8JhPDoyuyjK5BjtHdWqd+98ItPm6j8o1
F4LjBZ0ax4bugNt1n9tcaju6tcRtNgwD+trglMW9ASQm+5fskRSuv4b22I/M
oKzTOnOIC3BmkKTazQucCoZ+ra5sM1CQ7qkFOg50tjIgkQqZUJ5vyaT+41Oy
Jx6WY/+zOvYBJh8v+0SXIbdIOpZsIrFcyzgvycaTuBvBTuIp9F8Dc3VJp2Ah
RRFKX1RYd75m4HSVLiQJvMPEQMUH++pbQHD8RNJ/0AvazYLPtKGq6IwPakhe
dfZUWqdB61YBiDseOim+KYXJK/YuRk/Mtg/82LQeswfeVz+7pt+GJreSBg48
LR9zsP3oiX4igS6wXCX/b05Hv8exurVknT5kjml+wp3cBvvxeOYo5/4XwKka
BmIZONCKKWM6fiArrKlZPy92D0YjP4kL1Lb0aduGvcu2R163Qp73zf3baXeT
+c2fXo+L60J5TcdMpo36RoD2M8+x2uLIVACkQQOliQ2b2WrG1c8zVUp54626
EUQVmP3n87O9vBd9ldefM/fFW5xmTLLA2pmhT1OGZ2UWCn/sntaAkpsP5hkv
jyjjE5Vf7Km6+wlfc0GVx+LcHw/cd7Il6eAN1duhcTTeGA3wT+TbZeegjebs
AVGIKvIXPgkfc8G4XsrYqcAzK8BFZrsYKLI0uHnNvflvrVOGvD7hsseSEwSN
k29tiQE95Kxd+AAZcRlYTge4kCDnE+BvlBViV2CdePHn01cajAbacYN45LHx
TJ7mPba9rg63e3jZDQkUIDpcBZyuOh1Gfob9hdL2tWReWYqLlD9A02gvZS5l
AlWIG9vFeswmuYxKwSc0r61nMd+g+jm12to2asqRsxqyYaPXCwMcOBrzjwaZ
5OGXBFzcyhILWByUcqwbnzr5UuigUNbaRRoYAu3EpgTY8zkUzqAchbMeKTzs
uWuTlv56I5DsXjB+jL2PbogeEGHERrJUNjud44hVJyZpceYdL10Gd3+2z4d+
CIQCjd/7hg6Co2Q5BHRP7Qy0Vooq6W0/E1D92a1R7qI9WCX2BYy4z9SE+UuJ
qDSWLWFqNVLP+ry6Tg+s16TswkDc7K1SfuQBPYCJzqasNs53hHAVmxgZ2v0R
CapRfWF7IiePj1w3AvSsnU2D5C0QzxhAfOCxkEa6Iase08L9K4DCPw1Yzk7J
D6dH9NV+ZBPoQPyYyDT4iScSLa9u0ZYP/MTt9ObKBFeXX3EK2xbt1Pumxdri
gHAHgDnvx0OmvvwbA/VeTQKTTmHkZ584EQ+ICWc5EMvxHTVvHmwlXX8xKZFB
eJGDzZIejLoViPKkVD7Hyif/0Pv0JaR9GBVlf3/Vf4RmiVTeonrQUqJSXNvu
tEU53Ww+fOgBD2ENYWnJUr54XgjUook2eQ7Yz5VuzWGRltJ8qbaQ3J3zCWk5
cIGBjqD9LRc8SugLCbSIlydpHwXRQ5bfJJpXbxco+Z9Yq8qsDYpJ1mhFzLAf
qX/SLDgGzRx+AnInTjSUTopJtT2NqEwCvJrrOHO+BrpG4hck2795IpSW1FIh
rHelujli+RR4R+zdC5FoDfe/wV8GNsmrIa14NTRay1xXhpwzkovXjhCU6utv
mvPqR/44sszPsqhO3RzBvpBn/XCiMOM+fkKty5OJyu2hR5k9eyr1DvT7T1aU
csqH8RWErhYC4gZrB7kQ4KjQNTva3jp+J8yGMUmiiFrASFPu/qV16b6OR/jU
0FGiMuWbCGVgr/Lv5mJvFXw5Mdl5ql7CtvqmWB+RDnh7QEStxQy1xjtBZDuN
SraBTqc3iAaFnCJFEbRCK5DFdADDKRUiYajPwjFPhPQUINs3Js9rkzPx86S3
kZZRL3958gkQJgTQepyuwapLnm38owP7zru0bTG9P3enoQljW3mj3M32shua
G1WRy8F57+dErYwzmVG9Lj1IVwwPAgXFqhnlNBNnx3N1sURpmcZiukUlxg42
m6IGeSwFH9vpX6thhpWLOAhbiOvFCy2HI7e3HjLxd2QPn5K5F8Nv3Wpn6pfr
2TN1ybmN4v5YPmLE66JvcwTuDTXu0vuJLwtC14ucIsnR17YWU9hl2S1Geqyt
Xio22nAt7eoOili4voXT+GDTeaOJ6+SM7+dSm5eRZSgqZD17uT1bxCCntyj7
m45rnGvNL9g2QtUtZ+D435+MR/I0dx7EAT361q9igl1Wf1OCCu6lplYsq4Gi
8lzbagHOFB7Wn3PCP7LEuSE+0OVL/AVRk5GqxWWpyfcPInPf6uoqX/bx81Kf
hB8WJleHHfKlHPyYf0wGkqdviAKVGe0xaX7xBnIaXZx94CZiAFscooXiJfIs
J9ASE8EijzQr8vdoeML4/c+ELwO3nKDD2t9pcdREgHHD5nVy6dhSGDGHFzIV
Ne+seeQFga3y4lgYIjK7mJNg8Us2x5eipJDh9uwZ842hk73Vub2LlpSBA5eS
z9Rie3NwvdCTJv0gtr2Hfaramc8GQrtyINXTLpGkz4bk3oGxjBzz+7LdKsvf
2+j3nVSDFwoCy6CGaCEfdWg0oeA9sU/zz2/Yme76qJhHDsZLCErSYBRe1oCU
GoQFMBBjij4ooc+bvPwyNKMXu1V7YAnsKRvR0Btqhb6DrqzSvkfuTGJoMdMw
OO1gFFAEKSkPaI/c5TevjCW8yo8HRVcmxjzA95gz26k7TWNz2qlnys+7XbSM
JSrNm/9YG2NsZljAOLoebTy+1bXdDVn/WPP8WiMUveJ2ITV+L9bcV3lAuA/g
YhIRCBo0BSRxdLLQwVxq0CtTwxwgTWLTO6l3mhmnGP3lRSRdODVZQ8XJtiLP
QZYyVIOdijQWJOaQE+RhOO8uFVR/FlxMXkLeSlnRpe0z1k2v8ysMyAL6L3Uh
49wpU3J38yHSZOoY/lSmSWdaqpGg1QfhhucPYnYgJ5fYp2Qw0L7BGeWbjadM
6mU/QNXc/NOI0W9hqTsL63V0

`pragma protect end_protected
