// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wKp55ALtTYvYDUJev1EqX7W26FctEuo+SusP4I3llFw487RMFUhIB1K0p30n
wNejF91DmCrlr74FwAZ7ltwOrQb/MV3tV/j6+Ie9aG1XnQ8cesO1NxNt1861
TDL4dGoXJ3Qr5hdZY5L6JjAbudyBqzaYqoft7+i9o06R770VlGwXdcnLrOSf
SbW8o4J4hq7snFab5VL9caY7PTEBP/78HnoDUMQPC4I0Fn+6ZoKoR12u/3gU
CjHiJqzFke31TyOPTPQ9L56ZFrmL4D/oqmPFrx7xp7hsp/2/Esouy5n6tfzt
U4WNntTBnwraWbp/hgtW5SAqNFF4lxCIg0SK3aWunA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WWitvHZJcyOLJs74U9DoL7rfZbnnAK26FmWEZeifLxpjcCXXNTXptXTJXGuU
YT5L6hSlLaQuGlnc2G1WnOw2e+DaNDxTEivqGVcVSTsKnCjHYOVtH3a5VQlt
EC/5uHelGFbmHK70X4iurRnM/XFbuvyxtf3n1AXlYF1xxxIO0NhEE28kuGuO
R1tBii3OSNvbW8e8BJDf9CgLPSriVBVAesCQQ05bw668Ctw0nhhJloHhkfrF
ix4MtQ9YUTKWEAR4xJsjAgrhk12KwxpJ1pxtt5GOHi58L4zx/GUHUQrHuwYU
838u0ydLZqPMvw7/YjDwKycmMsp2l+nslp9hM/4Jgw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dak6RJ+WItENxOqemoxTq9K6IEC3HAbGEFDYiKW8VW6LRg0nHC58TMNpDnfl
el05smPs9pd+4W4oV0OR5HTySGhAgaMH/RRys0WcAZKhYhrgwYa4dT0DA4D/
78ZXiWSEWQDD6fiBWV6aKYKnbmzTnbfIxnyxsQJSVTVD7dGh5IQzfv4Q5NpW
t6z+1EU4ARGZLzxa19cHXGvPYE/EN9lqxykeXvjVVnx8hGX1siur+A1IZ0qa
NfpRWPDV0k7lezDu6EqxVc/OOte+ETZSKt6+KrV/+4nFbJs6We64qbaAcQ/p
CzYatRBnnFqcNAnG9XepU4gdWAMWrW8/VV55bQHPlQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IVrLwSon+UZ6uXSG7Pg4csRa00zZGMVVGxk2AQ4GjOnsCcVDKDeU9R7g2frK
OqMrKidE9eAdXSmIFYYfWzYC+sZORRbYc3PyB91k4V6LC2Mzly1pDCMJt4Ka
ttY/oOjZpbhLqfs79OsJqLLj5UV8D4Imv2IBT/Tx0iU9wGueogI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OhvNdyijogfYiq1GweeKp88YzJJiMW1e5nT9dNTS2HjRz7j/sqSfahniaEsb
/AhfLla04ZilDilvfy1ol+CzCuM4iuvKCFyqJKP44wnn5yANL0b+/ZmemTu2
L02s0BE7loxC/rYehcjqCxDC/ThatWJP9XvnOuY01LS+MRm7ZpH5t/72WsEA
ah3fPIX+3oPZjoziae0wgJP/1oP4PCkC+tQoxDgAQ5UJDvfl3xuiP9gGQGNs
/hJam9us8dlsKcoNVpfBwcDRy62r4GaLha65rniQHIvg5GWMYBxtgpFH6Pty
sEQ1HYGkCxGPyh4NH/M4m1HOwv0uvyuAp8A49LESSVMmF4njEcFm9FIo6s84
7LHZod3blI+J69yPM/+qkPSgR/ftW2qqiwE7EOyDTOIfeE6HsIVdSybBIboL
po0kCcj84Qj/TfhF18Kxxwe3UiCaV4zdBLh5ppe1EuLTahxu73EKsgUmzQrO
w6tYnVkIFcOOmBd0/dn49DbQw0m6FbcZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aqOTxO6Ft0ZUM9rjskJNHHfoZZ8bLo12x7YDi6lwyL0GQJuIYo1p8EnH4W60
BWhD9xcMlUtEw4cD40l4RLX8CWQ1mro9D/UOISCTzRicIH7FsoTso3k3tm4O
W+e05AaUMVZ+9jKyMP7pilct+PTDNcweySD6W4NTkk7hO4S97OE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R5GzaJz45fVunWsY0e8MJj6/rbcUKpmjtrxDT9wF2FBQlXXck8o2hFNby38p
2opTQJ1NymMdfoziBv2fmZQXJPjNHtXaag0meUOsJEVqExzp3cx/eNg5jh5b
hZX6ev9FXAWn0ZgajWNLJMR+J6lv31I46FIzkrEfjyfmF04XTZE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 992)
`pragma protect data_block
TVaHKcOF4L+5NF4bz3Qwvn7Bm84gK37nxsnH4ngHPwR6fBG2kJgoXKdJ4IIQ
0ymM1fXtv2OzH1dnBBksHQeoqYbzIhhttoXcPl0ED2TMpdR+ikECXV1ZOqp8
fICG+JXzIMDcklcH42eggkloMbRqP9jru8WuK2xQL+lJU+MGBu4zxQjLKihB
5dHx+r6g4IQoWOxkuBK3k1MAONzxIe4gFmW//ZNS1vtW1zCc2q7Ar8yNqcPN
jXi7eC70OXLFEZPWTXp9x8e6q3V3E4VHb20Ix2IOFhMPyx+fMQzbmr3l47Q2
AsZlo4YdCgz+T8gf6nKkkpflrzsorvavapqNS8FzHubPA3rL40OAlLexUnVp
6fAX2BSUTYWfNTPITBPYmS+Lb7UCVmjKPwEI2goQj9h1xg4lfcJGzSKkwTb0
ucw2gHEyHEHLmB5hC3Maevd71sOob/I5LgsjG5uOeYEjZABoAaRzC0//500O
0U4jZAqPKILM02wnzRbfbxqGrtKrp6xaaTEYdjcjhFdXknWwsXXQb5aOwf3b
5YnFNHqXpOLzCn+kL9HHSW6AsSWYBjpc7uBtVFpScMLlIOSGNt+zkPm5B3I0
yQOwAvDZLIfszsWRgL5pyeIBac2KRMp3cTgSXFeUlVeg6Syk2RqUnUuk7dNV
tdMWplYBCesLMaGwSlB947gM5JJjnSERVdgQyCilfaknSbdU4E5y5ui70hPP
mYBp9FCIO9I4TJEgD4oSQ3DMRgCEhzZMM9vgkz+n4kpTIl6c5jV/yikOdGF2
rPL91upyu7gxxtwh0A5tNz2ziXgiWgoNYAq3ZFDgu8fGauSN1C8os9K0NOfQ
kUOrrJ2iTJed6UeqAnRtm/puI3O+lrr+znmFURBZqaJmzGTpkOEvBGgBuvt6
sIaMdrPdvrydgeosNSKVAVkBEFxjSMt4BeScKwBT+EmkgG0BFJiLTwbQVhsc
d7guPfeXAq8eVlY5htIbbaDm7pDNkVpbSGCv2XVsA4cfh4V4pG5xHybcqWFi
4u9pjsSSUTeJr4X0vMNWXGCA+copQHpfjPnYRgwVKCttjfP6FT9ETTejTwsv
xcP2UyAwRbXhQlsAHGdsVTwytX+uSQoMF7hi0pzXynZOgTycsuMUo1ln1n5s
pnZzcef+TDWnZZlox4owHcuntNV5mHWT77/DYqUn7ZotUAv1wXRfi5Fl/zwE
wleDSu35CGt9948VHeW/vfIgk/lIcDLkIgG1UxS9VyYaxEEP3LpE4bbde33x
ttdMIgUNP8GYmx75RggDKfMRvUCQaC7iq8Z8JPGdgwaBjLcS3gX+uTrrjWXK
tSc=

`pragma protect end_protected
