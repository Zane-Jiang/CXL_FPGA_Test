// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EbTb0DdatU7Qhkd9DVkta0iIviuJ7SKBOd2IZIH9A9dwjnG8pHB6hnlSUAJ6
llx46/pjhDlIaFHIzXMb7UHv2Pr8FNP2AhpRusVIK/YyM6GAMjtUKp7pbCFg
I4CoAkUKTgOZFGBfM+VV25BjeFiJi+8bQZaQ3teG7LdUToMlXNGylF+BLVRW
D4w3nmOBMFv+4Z/p6RzRHEND4vL1ARJMI0t1jKSmrjzm97G6AxgRNmuNpizo
ncmFsj/ChLwsngBc4oPLuy8LEITRzJTerV66l8NzsFT/G8jgt4pGD8SV044L
vE6ttR4OZSgeVw4VPCiet2nMBq6Bb3r/pP9RaNUZ0w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kDd9LJpQbcZu5En3dZ6XkAusT3H6uHXbncNCFaeKVshMruy++hBEeoLTbtb3
V+XXZNs9oC6E2dPVMINFvhnDKNSTE+ZmvivIG/uEheffpMvvC+7PlaVYUg3+
C+Xe4cv+M/na1CMQfXNuyPhVCaaCqNW7f3WVaCM8SdMtT8WB1pBJ9L8MD32a
G3uzwRhNpYKDIBe23wRGpgkBiMtms3s4CBx5XWX9lGxyYWziQ+qUDYNsP79X
RL3olTXd7TlyUr4lqtmE6mcFnSLjlpfv/u+9z8AP3/3KUwd9fmd0XHnNrhM3
Z+N+Mv+GRScrboovFnsxaUg0yA7D5sOW9A6ePfS/1g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
B6xfy/BbiLfHFdOCELXVygxRusA7Y1MM/mG4M6JVMXs0BOK/N0iVfraluGfO
g3aDfnmlXPZVn+Gw927u9yBJTR8BKMq1hvGRoYzGeF1mYiyoZlnSWzo3wlqn
SW6EMQMzQgUP4VYIOHIaRiZhqgQWqhI9KaGx4LE8xPlDs5FLSB6BTEAoDAgy
5wfL3/RDoEy/TKh4pwYn82OIW1gMcC3xo3AjRvKz9NsGHYyFZ4bn4KbHJKt3
dl6hjdb56M3CqdavNsmMGYLohxnT2TTxhYgOMFJvfD7w/SBXABzzoKIZpcgy
8kEbX5eVwfoLKEP/4ysWyiu8V2GhwkaDtAkDYj1CfA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eo6SXPGQSPDRt+/kRN5boNyFsGkYsK/HF8Vfmmt45LbmJzJFRlPGQr69bo3V
IluP9wI/2oJ88EUzHFZ3rssV3uflEG+YbujZbp4QsB0i6zuYwAhHUY0Wcok1
2AOSae5DNgn/UGsByVzm3w7zHKub7POdU7bL2D9lBIUya2wwsM4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xoPmoQJt6TyS6dn5xshiKZzZcL97fdBUrV8ne9lGkvK+osWMrnSvG2/D1wcF
RGAw3LLvyexf6uWhIYW0NykdYbEEFnxTa4EZ1k5Qy0Bh763YQlCE+ULuu90D
1Jvtu9Fi0wHZR/tFG4MdmVcyquApOyd5mDVz681AWwRSxEp+vviuyQ9GsJ73
iH1SRRILjozWe43waFI0z+DY7bYLXzQtlKCJnY10bkyjDmF8I+VNnoG/n2+5
YZDvrThQ05FdGg3H7tvKgsUMQpVYw58c8aPwWjCpctHV7+niVGJMoI3mV8p+
4+Lxhrpo9MvZNJm5S2kuHTAWcDl3ji26kqwFC76UQS8S3i8BPkAUpzrVZXyj
+YDyYItMuvtxkyK/rxRfSVs+M4upg9z8ly35xZRWes00nae38TmRk4ZL5pMU
vywz37C81mbDDb6AVt1q4NM7/E3BygzKbYbAwK+F7ULLYwfUhRx2VpNoInXn
+vfOdY4gjbWsddN13N8rlDPcdpxfmU6D


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
F22NOXq8I4olaFBwsfs+AfPgpn2oqiS+Vf9M2TrVVvGRb2Uj2NftFKE3M2+y
Dd53PT1kU8M+80RNOStkBKbOLmDsJ0t3Ckq9m2tELliOF9G0VnjYy7JeYRDT
fC7jtJGLIM/zlD7lKMoRA+kBa4Tn3jqgJG6gNrwm4LLlYBb4PIU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pdRNBOJsJ6cYjWzbPwFKQEa+ZuiHU+AFzT1nUmcOz7T93wccz6w3uNjRiJbw
8/cIVCBxkE61eeph5pEwrMo5YRxwfLVPG8xURGODwPzoU76pgkKlmYoLff8f
/EvJ/+cdatfiLgP5of2Oq2a+uG8LtjmbdOJ0OzFQ0DmJPW4Idto=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6144)
`pragma protect data_block
uF/YmIYnEjUXKwABJSu98TK0SyD90SqGlnEzx5GKkM9GVBWdwXASRB/w3o9I
gBgWfmCo6F3UpjKUbfJLiE1gP/FB8HF65l6f9tvudkHUrlFfmKTPNEOGCoZ2
MLQXC2OXyLlbb+6W/MzDjlu7xZuxXkAm6EnFdB6XOENz+6xOIDI852Mpev28
25dyLzl2HhX5i/eMik+W3XJAm4tRv9TiMXhgTWsPdLRAUbwq9MUvlkN6QV51
nug/nkPwpy5uEgagcqZEtXiIr+Zh/w4rW9wXoLieKLBUnwzl4prtROyFIEXA
bvA8Z3zKnPJkqwvk6Tc2Sg23VdWFL6NMV++NpGrMrUtMvIa6ajlnfSQ3Yj+j
+qpWXHAQkN9lBofFoQ0xyjNdLvJTYzL9IuWC/uBhuJZhPyvtksnxfIejqHNg
y0rlUdsdHdOTfwpe4jpA3RUeYe4/CzaXvMD8W6ALJyo8+vGC03Z2rSgzCdI8
OREn2mL2+Gn/lrS7zlQ7NF5epNmgkOUCMQ6RE7pwneIyttxhpAyfBXWHQOtf
wOAoehSoRWSxB0AgZG8tC7cZzQjsxt48rECoNTLSPRVz4NiPsILtaai55K0V
MOUwPhTmZtf4R/Lp2uE9En/8GsDpJQCwTpFOnGSvAorguM2uQ41qwcRosYbq
YM7pcYeU9Knd+2vqgHq87wcszzEwQnTNxr4Ofvm+olJx6/lxGWbbe01JyprE
kMFDHHdHDnUqTKGYl0TrfZeWdKlbA13lHF3kHxAsckBJ0Xt/rQkkqHVq+pRe
crursENOj/jXcVCTeK5uCulY6cVdBTQEOVWPzWTeq7KI/Ys/7WtbZRTCGMqB
lqJsE78G33PB7B6C2cLYCWegcIKbuSy0oLzBKqoAWmZDtQ9QCykkAuPsW16I
o6XXvj63FCDYNtUwr7tCXr4wkm8swrwC6F+OhThVkmIr81HZgDhaQTCFK8NA
v04seDe4ZzODwnnTu1QIZ4Cp/G1nB0ISyCaq31gBkTsS6NCAO6zFC8kFdGqE
I5lbTM9XqMOEKd+RT3bWv8splm9ZpMYqvZFzLyVRqL4Wr6mmkbmp7dwTTa7m
0DwU/dBZ5YxbXeLRtPT9R02YMpYhzaGEwJeWfnyxVI/Z/3tZpMfJ2zW5k9Cl
NH5osvgaKYELcIYL4X6YAmpH/VmLrRxkx5LU/KFofhkAcg8+LHDCtM0tDsg0
PFllMI7WAwEull34bmrw3KqLPligflEpaklNuk3qPr8jpifb2lF90LQb5W8p
J4tKUnwM+4OR7tXBdOYPW0bc2sWs12AiTUWSiB1htYNZij4I+vBwaSai2410
BvLvI8fWqYnLdQYRky4+dZvdCFwP7L1d/FsEaNvAsCKMSy/6wxQe+J/kKktg
PHixSQ3ZTztr587b7cno5rQlpbFvSJoDgMXQqS444C32LqXbRWoY0HOQ7Ae8
ewhGG/E7HbJzhM5FAdnB/fVg5rSWK4IdBWYxr8clvwAzqeCyPi4g+sJyHnWH
UxRJak2q2KWkhwX96yTw2NN8gkyWhmHJKGmqLQWChhppCtGJ5gBR8EcDy90f
klCLqLPS3GPKoRq2PsEjugfs1m6mm9BEvyGZh87gtMci6XYs2Wob6vsSXp3g
geqQg8fL503c0lNY7B8AiV6LHcGVZTFNKm7dqwqcj3gBtRi8ftXucIZmIK10
i+p0ehEnjlgh3Arty/fgYhyk/wTQkj92VvQ7YV3QYTU7Mk8m8q152Vy9PpoV
rVfiRGW7RHZyW0wrcoDcKRE3tktmlRplqLm1dy58JWyDWX58aannYl0uW+XB
glRUkotzJXhSfGp3EMN1Kgi21KbzNCUDHIPTe5XA11Y2PmFScPZv5ZXNIwh3
GmPAvcpGa/HBHKy4ndYViQtq8ivHXIrKRSVBvhye1NH/Ydq7ClhYSpvS22kE
00BhgiVputt7ROxwtqI+nPncrXt3IR2yv6jOVag5MYgz5y73gebTNySkqyxc
O19mszav4vuZ1Xymj7YXKeuDmo6qigwZl5Q/THoiT1UzqS2cGlSHR29UAXcL
YFrwVZAZlg7jAzsGG4SvOHvKj2AxbWFlT0dEKQZivomQSuo+mxejDH4ubSZ7
gDG7eKfqbJ+LJIL1vO6HphQettoBrlVTAAmbLieb1QJ5qjslVyQYa+AMb35V
0aF+3jLNLcEZZIErCfimfTmpT3IQbmiUXPRtUVP6cGt9UYimN+BtNtscnci1
lGl2bcBgPkvXAqGJsD+IsU6IEK7bhNxtG0XP9GB6PPdu2WvkILe2ifNQptWn
dOP6BMHfyob+Q4hfSi1rquSZ0afI4cU1XRtp5RvN+16BjmN94RGsyaQl5Y5v
F5u9VQNpP6Gg1FdGERsUrMWdwbOKXqS05g5PHWIOLc9GgmQDJF6Yw0q3Bp+I
lvUoXyvfrJ1l83d9ly1N3wCEkQ7e4CC7ofLIOmgJw3A+mxQBmb9sGGTqXCX4
As1A6tOyUPyxRGkdlmnL9ZVjzG1w+sni3ozvnCtQDmJ0sFBFlrxOOWcDktMX
7UW/mbE4lL5kv47bepBGb0y8nELi8i9igCZ/xgxkcqDljntCmHAZ2wWlMQ0I
SU4NnNzzakC9JCSENXh8BUldENDcVEV5JEXzKiYqcgZciVAJtKR71FEYmXmk
gg53DOhioF+zrFoHL3oYufOr+rit5sWHhsdmLQyDQJZxGz4K/vKfhT1zcFH/
T0gIxoKOwcLZfQ/Pdw/M0mQF6QvxvO5SHm/DmfQOCGeey6o39WGc3yhJNzfz
rWZBlj2dPMuwb5qOsWLIHP0b87KyXO3MA7alWY2RSD257mgi0Fac4bD3z7GA
Dg15YUwrNwTygGFTduU66TwgSwHtIMXl32KQ8cMaJ2Jd16XJJloiGcAPjKnP
XqnWxsD5NUAaKWhfs/PdZagni6IxGGFK4m7kgixZyFCrMpz9wcCJTlyqrKJw
OmwEWeanDBxX1Z1Ucyal2X3UnqyjwcMEtH3MdzE1xmeoJjLDTQDgoJCOXV55
M9b53QnuA/sV/YveyUeYk0Ol/ZsOlK0FsTXxTZPl7biCUYygrPGYf3po7o9F
MDlPP+cJZXkklvkcL1LUrLq6B/du2Ofb7bM4+UzDwCw9Mq00P+EDz7l5Ayjj
GHzXeNH3sSt89KApx9oW8clifN32iZNqoMQwRkKLl+1XJ2x8zOqkmGB6forN
m4TzQ1WXq4vPZRoh5y3oEugBGQ3W2gN5MgzvwoTyJYaWKLbkuDPrKfm/hekG
Ehj0WDXXQnqLT8Arw9/jRjY3PypNxkO7/ryciNRNA4J+Jg8VRJJ6VZ2olTFl
HACTFOiLVbFBPH5gNqsvoikAHGygfCxUjgLbuUoYO9fajKXxfxrOjbngMV8v
nG9DquU8gfqXzCgmE2fDvHIM2DxiCxI1cCMLuiStbzE0ljhu/ZyjLOzbZz+x
ThJ+QR/LHobPps2w+0SSaj+X/+0Y8SweGu0m8A8CINesZvBUk/gwxBfyHcq3
nCnZQn0SfEr2DwiUwsFY8SzWulrRAaJHWZUX9bXFSNMpNkFZNt+CklOcFKfc
SZV5ZWHOVjbAnbB3zfxj1m7NWx09M/0CW/5bfRyBQQecF0d+itIlfou6SieA
UKfe9u1GEMnR2+WXxy8WdAPAnBJ80zdQp0nyf677P6uFfQ6i5MrjrB8xA9bN
33jnqepYjKi85dbjKNzY3Yk93W5dZk0tk+ozYeXxzYakkfioUSqwXA36pI6m
vo7A2Q9EilETIEKoF5Bp1kk2RAPuEVqjmv8SsrYrkkipEBo+Ez3mlXoE0BxU
S5FUbfnJGLmowUqPq6ShE4m9lju5GM6+5iI5sLPoWI/ayjTaky4mbgsbES+v
CkhBnhnKRWTASf7AG9CqLdupsiipfVePlRCwpMZr2O2+1EmR9yCg2fRGqUbM
mSzcfmlqieC3jkPOsYwDbuv14CYIlMQ+OOx8QtZH6zAz7yYdzIW63E6HOglu
Ct4QdV5TgeDV/5h964eHcaEr2A5T9ZEdg3ZS9FJ4lbE8ZlthZlqeq7pHFYE4
dHe74CTknVlMHQJCQa1xt1mni9I3t8zftdvic6Lm4Z1xHPpqmR6QShrBnEX8
V53V89Ux0WEH8dLRQ0ZaTbPfTqAJOGSaloZ6s5MQTX9VTOXk0B5xHTGlSnsq
gSw1M9/fVxuZ55x+9NcmRRyjyFRrlxdwfVZhlaK6KTdXzCz9rW57RnNpMa6+
gkL1bQy/eWYygCGUWHe6GRfAAWxzQDmG9bRRjAHXd6tvjWdCI1XUBUb10iVf
zqo+/d16Pu13mLA9UuaI9+lRWhSguOxmscu4WTebmwZn2ENLGeuEGEqBlLa+
ZEGzXBJB3U88/sWa5ur9Js7HWIn9vrvpCMdQOkMzv4YD7cn3cZZX3tQReu5G
BxS3RFE0D3/cx0LsMi0Tj7AnOW4TNPsV2jn0VOdtXjy4NQ8jjKf6Yc4L3KMz
l6dGaTppAPYhstYLQ2IURDy/w1ENjNAGAm8TDfFfLiWqgR+YCcyF1I87Rgiv
CqRCGMCaHi70/7dyXGUPTzLfxnH4oS25kUQrD8Cxdq297RNw+Li0MKSSurSA
HnBiZStVJjapkuo3wfsD/ti+eqZpLpLk04qu0zHdvs3qcHNw8RgMEfHJ/Cd8
tLQHguXcULouuDkFBpe9V97joo7vdJ5apwCQBZnphkHLjJ2NSyIjl40uXtbL
rRd1C6p4a7SpRvQzJh52XSbc+oMaSZbLhyV17huS6SbIxlokRdZJ2PJa+jDo
osX/U5GqN4vpsVSCxAJgZ6Lt6yItN2DUKmTym+Vn5KAOy6exOx7dfXM/KzlK
VdzKNJVnkXKF1QlLpuOSQbE4eGICMYD/9VTLrrCWlHqDFl0ut4zKz87KT5TE
p8RHa13Q/rhMR3DHIzkRB5No4nGd/U8gs+eFgwUuN5vnibdkgQO414vYpf2x
yNY9tNu4YhPaB4Bj8A0f7ORRBy0lLtXKqylYYJAcD2N9rx9nxbhCUvOEW7Tl
UFX7VAu5HT/6mblFcJxubLbAonwHQBk3ErLIBov23w0N/xY6pdAju7dMt3uz
ZJSLaOj9nWGC4M5HtEwbqi14n5c0xiqkGpg6rrJnOl65P5waafKPMnD8H/xq
LqAySxys8mCH/5kQUV04Wu7Ih3RWP0s6RTMmy7l/Za9WBieI94MSx/m2YRPx
8DAnU5IGnc8MiX2ojtiN2MNZmDXemv/MFFObvQpjUIcEmtMF0UepDzozpCB+
iXWkkINu8HJHg8B/3H+GRgF5UoCzJwA5TclH+a2FM0VEb81ADVAbVOr6Hf4j
Coa04lQVTKR9/rvwhP3dPL854HJpkl/lGHI+syytrqg4qiXybnKed1F2q4lf
3hldvBnZltaugWjo/tvg4kMBYmWTU75LMJ6kjSTMuXms903js/SdRD30ojS2
LSf2KQOvA97V0vIPpa/5u8iogGukpa7KQJBBYQES9WW56FYO+p01nApyxIl0
roqjG/oPvhIwfpMy4/q7Xq8tuX4eqVPagXqg14wXmRmLQFf301UOLp54RSxE
qZdTfHIJNvSLPsscicwFZRoQEZpO01vYcT3zB5Y7lN4QplVJ3ZXVwxRR39bD
OfeOUUNsrHDxZrFbmLg1weohZAPMe9IOUVF5fIrYbdhRlU9g7J9JPKbd3hyT
S+PHputp0ciDQgG91nGo/D9JuNXAIhKUiaP4bFtiSaVLu5mNya2BNIk6BikM
f31kwcJrGlaFGaZbgAD+7utBnKocoBpj0zvIaXQRQcXUKbQv5AqqXwY42uu3
ZPBkMPBFr28Af2/rS90Ka/ama6r6xSsLRec9JEGU/5sgKz381RcjrcTxdRV6
TMYHfE/SDB9FnbNoywujR5WPcJVaRt0Ge7uZaYbJuqN8Y11ZSzN175s9b9yK
BmpXCESF2K9/rOiBJN14tj+w6D9jgTn+6pcssOv4XLTk+CT3MjvRlSGBTKlj
qTJcF0U3HKQ7zKHJnp/DOFgqQ+bjSmM2vhan49IMto4L4uyOpo08osRW/nph
5LJLEsRfJIE46pO+mDaeHZVoP7kZXqpYZqobQ3CUVdqYAGrjLup+5BGjFVtM
Ex6lTRwmVqjJ0GS8iExNe8RvBua0kKww9R/CHnGDVAw5xGIIALPsua+s32x3
8+XseYV+KiA6ed7zbJL/hxrARdpkX1ol4jWiv8wzrq0jjMfWs372qYkAvhkp
lto26VCzsyAyKbxdKLYG85InSpWveYGC3O7Lh99m+ef6Hjz89EooJA4rcOJJ
YSTSMiFf3/iUzx8wkVlAKfwxUrckm5ll0KsBPm2/ygIorwxkUvLuBjpV8B8w
lsmyVgh/VIiG8Ooe08VWk3LKjUCdRcw5u16+yZ2nW/tyP9ov0VYZkKS+9xKs
tLv53dx52uQT9BDWkKJ81Ec1TVhaQbQwAn6tcXeTL9PP1T94UXkz5QegO6tS
8Gk+7wBQUMnc/kq1oMN2EaGbyuSpKCQvr3qUIX48c0hpSuYQdQbojLr2KKc7
CcZXLY8r+Oi88jq3G2d/PrIdXhJd/nn2u3rqDv/ZDGcvpghQbWCSTfCuXvJ5
zNNRGnZsAzwajWqM2oBJHMGmbe/rDU86sQ3A+HH8+c2OIk/NJWfpKkLcUQ5q
0fXIHGXm0NVPJiQES2ZrmPi7ATaGvQkIEnXeoZXg4MnTsCiouKJvEJfw8FSx
/9vPG/jgxi1D7DP0CUJ7/Hi585LZacHXao5ozCF6I7zR9yNxC5E34FTOZRh2
sp24tRpbhGcKI5fIYRSKuDde/VPZEbfkQuxSBYK1EbpTIEgay+pXG5QQl13s
A+eQo/Ngp03FiDq/S/0DkexbibXhYqT1OAYFVR8xTaCx25XNh13pK6Jj7B9u
zth6ilEev9bWOGQgerQaFWIsbN0dTne34YoMg7K3bNLoNggvEPueo7okEqV3
CTVra+0m1+WJy5hPtHwHYx+7C1LMUo383R0RPY0G5C3l5GmcxnRi98hc/F3L
GN1/fZ7F8buIJ2eJriNzaPNu4IfiolaQktHIEpNlV0Mcai82s+YC+dF2XNsL
dU35qPmcNjt/RC0JymKS8+XXOQLnuaOjaw0XZ6lhkRQ8UOnDNGnlz6ZQ1V85
DG3tVgGb562Lzjpu2sXxTjO0dWIBAqWnyZ7WvJzB5SSHOTMBZA42hKlnrI72
UFavum+KKQaoOBRn/BcV3qQAdSFkQUvj0PZkg04e3JlOoKE6L824x8W8p/Bz
b8WGY9W0qMzoaTwUO/kIih4oi1ZXOjuj6f8WLkzVs3DvZJTkHG5LAFPH3SEq
xzIUsUdD4pyKVXG9GTk7gaY+L5bGS9Vx65A+QDKsvm2PsWqNsIWRypDuvoOv
GsNePPtQab/QmCUCeAn3loVdIn07l3BTqFDKTz+HnOwCTcggr8Eb2FtyYyKu
SmIvM412XWVAOuUo+mFBIEMGRk2XCfScU3tJs2OZyMgpSKR8qXYWja+wG1qG
Y7cbHEe4nmBCTs9sn7F3Bqz2YoAvm5vbYdJlOotIpBFW2VypP0uS5GP3bKyX
t99QYmoI8rDyVP/nZL/fxnnwh8DJC+RZMY3dYsQku34bEIPqmtkBfCsTFXvY
7XFE4ybqdy2tMSfxKiOy8lYuwaBcGL5TfiND5WS5IBM7sAu7RwNeuI4JaZeV
BnUkVJK7OdGi++YKLyv9pXRsUclf/TENzm798PEgQWJRgGjO6mehg1Ik4sO+
sk8wQFAzE34yu3VOZKAd7mvlmVx+67cjncLJz8+QBBEOUfVY2W5xAofIEedR
VqskE1GXLnmn72DIX3BWyTJ5BoaWapyGVgmpeQ0UYdJ7P+MlL0lXA9r1eRtf
1hjlsiwBO+P1XoFDYOEXJOOi+UfX+xfvwDpM0AzfXsgRuXQm29K42cH5wAHD
Jf3JH6JmgXlEyiKdNfvqt9DKI61kFdfNM/Y5hLGAvg/7tDWNyNy9vJKVpN2f
/L2Z+HShBnKC1ef/xeWppUn+cwoKNgiZB0oCd+Zw1EcjOx5cssATfL5OiGet
FeknUcgLn4dgMM6xCRs/1eSaXjzyglOlHE69gXLHE60zmtbY8sfDWXIGFHvB
mNu2gaB9j+HrtZ8YyJqfLPMc3l5X9RE721msqe//K2qO8+duV7RZTgcUEmc/
2HMF1xJ6+Vdt+UJi6bE5F/Ib1GLG7MPiy7YxVP5bZYciuhP75RmysyNsEKrt
cfKaSCWM/K4UFcUmJm8txnY8ZrpsSMz7

`pragma protect end_protected
