// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
phfsQ7MPlAPjKjxDjg7fGEUvtLLbSeC4jJSxrzz/cqPp4rUCv31OunIACI87
DsPkf99Poq0tvQMb7uy80H1zkGzqVuq90JODfGzBnXj9B+55ZLOZNmp4d97O
xwrLW8U9qzJsHDCM5WBlwaX4uwH9Pviq+R3HmKXGdvNlayOUSnDCjqDcXljx
uQbnk73CtuMYmu4GySvfMYVvbCxQ48YW2BdyD5a3YeSBRMq3kwGtxFv8pZAy
JbHSSzU/jkps4EBhpZOOvy/3YqlU2W8HRkWVVJmK4zRf37hk7VUDh+62GqhG
agOFlN72BceJY/rK/5i5IrtYokvbRruQrUfn2xvf3g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JdOy1de/dPxO7AeSvUFur3apAGUr7/pEpjyy2YGQSr5p5ikIHUeJnibdQE7T
Ll3/OMaTavsbIBSAdN3gXWjS3BtrLL+Kxa0NxHQpY2nyFPKjpQZ/wAVKc72k
7oluxC+qOzsI8SE6W4E82nbEQarKdiXRpmLTJe1p286pG5CckIs6eU+wSoC/
rMODd+7+IhW+55FZFbQmEoF/BRRW6O3nt6vsXJJjnhR/xwMyUvyj1L07NiQZ
N8hiJjIeo+i4R+JTOfqOv7dhirRTkNyo4N6xExjtl8BtfZorAUApw7k0dLb5
nBg9J6ZZE/zwDVbhevvxfkYmKUThtFlbMKOFgWkgBg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y8Aoy0YloA89PXtnFDZoqjQxetI5mUChQe96QPMUV+0CKZz4yKcuyeODGVUl
fP8VZWrkuiW7pP5Fy4Svuxrt0v4vS7lf4iwsc69ulclBlWATOtw+s6Y/mmyL
RfEK4nOZnAJ1DQncVPlM0tN5l2yuc0K8hENw+hQy3Gzau6gBr7PyuocLCaOW
6ikeddRc8UKYOwLdvd3qhp8bHGYRvnUlOwOE72n9d0dypaYNE/oUK6zqpxVP
GUvwljA9/XZJ+TG+T6Pw38rt7xOtf4jxmYb234GI2fc7pUiw29oJpcpmXt1e
JxSUKmnUI++d/o0GaXMGDEifRWwDnYASeVFo3xmamQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QlPfkjUCO9Ceme8lCgFwv0zhzaT/ci+Bs81xscqQNCTau/bZyC+fsuqC1Uk+
u+o3Q6SBopNonUGfEUxLYUZE/dZo+VMOl+3wO/6NeNqC8mrqauO3Iwj/1H54
AmYNR26NfxOmd+OcV5NPHuMGCoKnK841NADwF8WOUwdK66RpHcM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
CulTskZ8+WHedeNZ+xQ0knl/uEitl2l48Jmpn+/EgvW+VX8YiTegtI6StblL
LpEodowKnhrWfdWeBM6WNaDQfS5NLb8N//uuGAHP1FSyHNW2FcWMzqkymt9J
2hSZpQOCg7k+rQVZ0m8DVtBv6FKHa0RRD0jh2XZlvP35gNQVvuDtSpsZMevk
/oQe4YCRgPCWyvdivfoAiKwOi8ukhCfi4pIfc7bM+lLoP8nfSM9mK7F2bjsC
e4YaOvJx/oM43+Kp+y88Leeb/YcsBNM9SoxbG2ouYzcPCWn/wCyMtGxf6GbR
yVcSITXFJ3g41dON16LRq/YyLzm855zOWkr8PcS3oFVo09dSyGlB6zwZoxMD
NnXKxeNmurzRBuy4M1ZAlsp8i3GtOx3cs9UlHG+ei9dHpposfcaDPy54ubUJ
OQRAWLekQxJ9r0Cgy4y8SjK/XJcH8CTihXxtzXVY+kcUBROcJCJECmoHiksL
+Zu8BMRbVFajpo/rFr8BezrtezkphXcF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AopO/4Gb2JzWP4iCMYoEjcYK45QuRCKUgVOVLIiaPj9TJzPYDebx8D5B37UU
Xeahu59/DeZ332lcHdRc1JQSEJxIMXt73lGlhnXCPUK7MRbgOwM8yIjEP9nS
ldtA+Tjq/DMMvUUoivfthO6bggnJz7fpoZgkOmzJFaDM1iHKaag=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dtZsSLCeE5+2Plvbo3itVV3yELRx4czz90Xezcj1/NK3yuu9Z7FCpMXrverz
WcDjXrXf5QBCmFOxn1z+cBFeVpwQ46Nn7e6MYzeqtk++J1bWXcm9Rj9/J29v
woLjEVIttRWJbQrPN/6f7jnbqW1pCndPxkLuzrdf6+XBmVdjdB8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6608)
`pragma protect data_block
A21i7NxYQ3lYvJaGXiVwuPBAOnWruL4RpvXYJPgMnHXxuYAYYjlBmI3duD6L
Def2e9LJAttaLJ73bs02nwyxEcYNYAcGdQgR5V0GQJnIYSRE37DTNIrdQC2z
6YlNqp8/G02n7/WOjWbsqLD6yoAGrMuzbjf2AZn1cOpcz/i+53YTlQZ7+i4E
W7GPEu1lyxdMcp1EhNKWta5ZlC8Yaj7Hi1E/sFrW6U/jQjWMM/tj7RIXqEUW
AIqRc6meLOmomvMgy+/vqlIbC3i1qaf2Mf085IwpU1W9/iKEjiu3d93igaJU
/lccJBy6Lav+za96+yYT5kbTnKqmX4A3e/uHoJ2YhUnZowKCJu1L29pw0Qby
vsna72QPJCeE3ab3JrKo/g85/A6VAR8JJ91cd9rmvyS0R4GNKwo5vEak30bO
Ij7DHcPYVHLyHvrnh30A/x2Km12JufJVcDRlJ4VXj6BhsHn7V57F22MXayB1
5NrPesFXBXHD3goFSGIy3nO5tYyZ8vesI097SrZ3DkkAlc57rEfP8KsLL9sz
vI/k8UwgpOL9dvOzn93uTatA+KgpTDBxZF+tm+m9WOdjelgFgQYttAjvC7A7
2jv1GLH7KNetfJ4elpm69Z3dznz9YabrSwr5gg5a7AIKWJVJ5MIs9Uguf3HJ
Q1WJrcXb9eUmjvUU3qVIWUe4iRFaOC1+NS1189kQ7thoHOISmMG/WRxRk9Fc
dC4Vfm1e3HN67+a+pY95PBlJtsrdxjivp3ALfC6ggclk2CoSlCSX/MOXHKFV
3YjfrFGjOfs/y7Hr6A4cELIVKB2lpJq6qmv/xG933XA9MdUfoHomIQ2G8Cq4
ZebzvySbTsBJs5PnTBqtxumogrbuqgHVF/tcI8QMZBrtX4PbNsbZSetGrBCn
TU963lbynoXh2Zksq34obxc9Y98bZGRNsKv/NqyYjxzWJ8rckbD40wAXJRJQ
hU/1fCRwX0ouI5t7XagfjB7qWhLbUZunyHgNykLIRw4SmskQtIibOC87C7g5
QEw3KG1SxNgU8UX//+I3b7s1VfWjikr+p+qmfNl67kYIkm2PNb+FtSh+mFzX
RNLZMcme7AG4XX8cvI4MC6LgTchK2sAYAoKdsqlfE3wiKv6r2wSrFxvi1zR4
gJ5nBqvu6A+vY9UMd/1VIzvyp5EgsP0dx74zOtc0jCMpMJEU/4HSHEh4eKYu
nbcp6zQRYbE8eGradVmn1YHfcJgY70+dCzCxMUDtZ3OCiu2+34GuwvuiO6OL
vUWQc37rvUAmTgxB/WfKnM3Z/G9+vZ4ocm3a076/QjK/xFncqvSgvXY9Uica
g2ZJe7lvsdmH5VWi9lQBK9oXoZvwbtFUNUQeLGQHvrSrPt6KaMtGCJK6/qoC
Byh0/MPaBiJd+OkXbboYR+qSnKnx4TmhJm2VG/OiFjC8MooXJcSYfYp0fOi5
HCBRrI6wG8t6jtMxLEB48+CpU2Ty9SczAfZNQtIWM8j7piyk2e2FxMOBuuqL
NxKvUOMiJ2CMsJUlUT/hxMn2NxXpR0hwHxqaOb2lBSxKQNOcGv0+iCS3o8IA
ebHvc6M8NVUM4LtT67++Y4IS9tPB0aDrqhplXNVsxbAOTqNJz/LT0cvNUzj1
2g8xbyHHyFAhOLPfYDSw8vki3Dx4wSejQUU1FajOJQ9HoCOPcMfujcj4WQLq
G7vzlDXAUXj2bKqagDJ4VpfizQtswmMfDN6g94zdR575EaKVeRPirg92Fxec
RFKCKCATTdHdyNLSHKPQh3qwbPaGrij3rzjgOqDB8Iq4iufQ4/sXObEeFe3/
jY9edY0PCcukq37+E92tUD4S1Jqkovh54adjDo5RPfrEjRdj+S5TVEXzG8xD
qP15VVqE25N0Bd7iZxTmEiGtUC8trMeB+VltW5Y5OPIVKxmXij5JorBsZvkX
Nn/Ua+WmZxt4AEJZkosVspG+GWLVBzDSkUQdhATCYmrLuc8VpDAJG2YfIepA
c4AuBSr1QNXi0uBl7XtOnr6Vjgjzv55PwMSepxjD4fK1RMpq8IouPITY+By0
IxkXVJVERhrDSt1Wswv1PO4gZT1z14XhWygDfNHIMMpbvRnobhIqbJIroxXn
Hqza/cM3y/rjFRQMM6rgBH1zq0m7ertTWm3br55uOoSlRs07N6z5oux8H89s
HTd6+oHFX0AtDnmWh8qZl0a4b1q4VkYDM0di6sEIipFa+0oYCarXUrJAN0K6
ok6A4xyoPaRDu3MAFHWyTJGw3ZhlOL8bsq6wq8PcvIqm8GyExBiiH3BrZaoS
vSbIJSL1XuskZijjhdZg065BMsCfKG0DODBrCwW+OFocwrfAg4Y3eKYMJ27v
sW9I91fFoNszXFpgNhLzzdUM8MWojFWG22uzChpVjV5/KtTeQMSX9eeEnjfR
kNq39n/4NYcXOJSqCbUxYu3GzxDFCZ/2w6FMFYMxmjqeRgvIKBRxgqJ3Qzh1
zlLd7hMXebn1hUp6vVKDJbV4eSOzBe3aoM1v7Txy3Fzo1b+06P04l6BCux8M
fxVLNcPDh7Xf5R6pNJ6mn6pz2R75NZzNaHtCfFUaIlu935U7jjQUVw4IKpw+
4ml1eG1FSXF+I2hkWQrqQ5VIk4siHQitaXFvUrPS0W/MQpdPPD5tEF5oXRqf
a6Ol+G4tdsr8J246/xf1Dg/EGw4eX1ZH2NAqhfUzefq6I3XznmZi/bLCeR05
lrBQUaZj7qKobbOnIM9nHGL1JuKXvWCQlLnhyvHHyMaIJMknFRNBf3nyHpZ9
bRKKmL2fuIOT7BN0kj7Ji3mHVcPrYQe8klqVjPI0mS+co2OQVXoufpE/tzfl
pzbon+aM5NYr5IauMUNppDMovI9HwJOurr4ckSQ0ymjwe+h+xWYlQfbjDIkk
mRcrMyumE4L5gdc/DkQfUL2XkysKsV8TapRIJDk46G1ypt4amxQYbKl2vbhM
FU6fl+PLx+l/xaq9WM4L6Y5/BsoIrdY6LD2a2+JrbaCdJmgAJ11/dBbAt5DR
qtykpE6Z3rxjoXpOWmPv9Od2KDm3+iRzMlmXLus3tJOdUhFpyThDQdnc/rgQ
Me5+dcfZ9KwOTZGxCzGmgXpLGcAaKEpYuGqLcXT0ousPWzETPoKx3Bi/yxq+
mqqD/gkUzuBLPuYfdqZpJgOgy3jyBQgR1kE9PYWieGpP8c9FhjRibycTK7Du
Vc5B5514H9rxCNWTr1zVR39t8khh95LkYtw09YB4p/w6OMHsoTvtjmd9Q2Ld
azQ/uqv0riJWIq1sD3Ecm/phqMm2Xlo+SVHfMicEwaiUhKdt2k+9I5Hvw9sU
lcxEmmfNvblLno6uoAvYhr5rzOR2+VXYsb1qMoa8H7yfUdHLhjlvPFCCG+Na
WaLo1D0iuCr2Gq1R+9Z4LwoCxvUjBX7TtA6xZbAgldEUCNbTUb+uXCezuCqA
kBsyXVRyy6HShKdKjBtJOOXTFxLJjC3kN+FGnnbGdODMcX5kB1tmXgIQoFSA
ASkHol3TzGPSsLVWijwX68Hgq62zyOzqaZR2pl5jlXavBNODloqwz48bZOIH
lGce/thKEfBVX7d0/7qkLKWVFdT+PwBBjHA+chcb0hmLP+e8hW5HOrQVNgwR
ORYUbdG3ADf3Q+Y4boqbD9JNRSimuElgPfl/kZJzByzTX4jhTIW/snwNwgo+
2BRrxtIRfbma7TTaxY3riso9WCi1SMX/eu0qVltaeeLVVtnHDK+Ui8zCDD/n
N/WbcwXR5qN9xkCCFEAMhFQyI0HvzAOzwup5gbJ1DExW71ROzeajYX2JDZAR
YEWOiGb9L05bSy6T5nJHIG94WXx9Z3lihsdxTAQXfR9aqlo4HhXQ9EKogyS0
VrvVa6J7Ois0fokE6O4Yepki7dXPbvnHL/R1rffetOzqtK8zTAKYEH9uwbim
KWvh85gYWpXLAyEJhpJsKT165m+4B5tGAXp+Ecb8KAK9nuDUly2HO8IJDU7T
3Eygwl1lNNnFxg3GZMSscZKvXQCvKL6OLTEHuOBb8nHMjgC0YR+f1riChUSd
eNKGRNfzATuBmNKYSkLzkfeNFhlpVu2lODXghdXYTeQCXlS4+itYilSTBdLI
syv3tZ52Lf1ExPXISYZSjWcPYKo/dT3tgO6q/DQYnFpF3Y1Nc8mp6Ki7EqlU
WD7xCInuIDOLXxtHiqEQDbJlHKqRDIWxKKbIU7eOizUt+w/ihBiTp7Hp8MVc
QG0Ft/hByEm8pWQU77DBSvabAjpnNzb4A+9fH4UX3228GqTPjwVvmwH59x6v
XZVMSd3Bublm4x/I54T8gb8trn8qjvR5pxTOy+wMQjPEH9TberWda5V7VojS
8efA1/393cBlpXU4/Kjm8oNcVj1nsHl7a9mpov/11QPK5HfX0z5DNtpsLoCr
I5rzAjdl1+uggZhJ5IQiRWWjAWMXAkmc5P6kwDChlfp2afOdTQC7YM8cpSyZ
Ugzm17zlP/PDbjsa4S2gHYpl312wE6LRjSYTsxPp0G7QVlEXFR5+Pox3HydS
tZktVK0BSLaam9aOXbgzzBaaS2nUCdG+Si+hLYkIXIUU42a80qt+SrDPvpfr
SbxT9PoRiKv2Tpz5kv0xJwP1naq9NCg6iWYNNmNqWMjAT/8h9YGduquuWIS7
o3exSkFC+pGkrKKpdpR0SH+Edrirg9Bgt4E4mVVkTBNTzihjmClwNzMsE6uf
NoGja4tKM0d2+Jk9KcVR60crZeetJ4t06rz12UBnwaqjO5odrSyGbb5hgU47
4HlwpBLftp6fk8fftD+xxio6scmYju6p2oMbz5zZwyVhzMcGsnyuiRfTMaIG
cZf5PXmW2SU2mfnnWHBIwJqT1dk0kzOliw8+I4w9LEQHsu2D7U+OtGEU96Ox
3/P43j4UTdWBanK07jwzaTnqhuV724pr8YPsECMMBp1+iFt88H4D1Z5gExe1
8Cq0cNauhJwGdd37DouPZ4xcES65LTDEI2xP+FCaKiC4TFiX6Kr7EMfwv7ql
oGk5kYTXeFPFp1A21Q9fn7VHSr1A8Sm43KJht9tieSdTXGP8C1/zw39k7pFu
1Pkq8Keu9FogBbT+tQoEPCUfyJUyh9Bo3cCJdRKNmVnU8CfgJcpJSpPt/Qf7
T0uXHKgqpIqt/DTs39PifS4mvnYj+ObjdPQ2wGqhDwCtONBWNwQjaeXX8EL+
CGW3F9Dr/8ht2uus4zc7Fltntq/eGHmzAjKXTTQBeA4v1G9du+GM6OKhu22Q
tIfiQmwZ2a+ZD3XtQZK3f/H/VbemvvuP+jbsg8UnxB9QsOltv5JiTUgdF6s2
t9an/VzRX9V5Zdk9cTJ9nV8t/AZ40pUCIUppMRJxzHNI0TPR9L9+fQB7zx7q
B8eGXZF582XYT9NejYCpeIItCvV1JFrkkTA/IK+cljJmWelb/F12HQSIutSC
ffMR4q83R6JvN6Fs3c2STCtG8nxMpMlreoUn4xCczPXXT1Y6xyoN24gGhq7R
FxSvkvtKE8Vi8Hqjp0v6CNJAM/MUzpI6qLFgXhOyS75hiwbiN7aonOupxVMV
QeCF6wUJv0xtj82UQfjgC0kzZzNjX/XGNDhnkOO77ojwmuh61vDnYFi/scva
Qu0TlUYGphBQ1yHb5i/4/Odf69CZxjWpXfQl+BadUlP25m5RyefuPTkLBVBv
6Ay4LypB1+v/RHtPHRc1+f55FHG1wslz4RGfiDHZYM5r5xval20iep+95Sa+
efwqvkLdzkCAhN7S5VzbcL4i/95jhUiYeQPRhiRhrU44oYSOAVbWvLr8rxMG
LH/IjlwvRBSP4OoYMPP+Lpfv/V2qJ+ErGsfIG8J9UtstbJckwPbPA57UnLKS
jfXCkipMMuPpBjX6wTxmXu/SjJWXssYazchbQQ02dBPXG4R7duC0op3dfj0M
t0EcPgb05y0gb71O+7JaKluYftiqzc0fWSyMthBFXHIvdxVU0hd67aftMXHT
D8+cKGvcdls0v35erwX7xn1kZCyqpFKXB4/yteEOUZnHpuOR99cxHt+Z5dYY
BKPbPVIP0Rmd5VhKRFJIJEogOYh4+CyfkzoXXBIgsLVkG33DP74GQvxwPccK
6RSNThk34GKD/rneFOin5Hg/Po22221zCvdk5nS4Re3lB7FoKqC1Nv9MD2jE
uZZOCsvEeKWS3y87ts38HN7dNWJuz0GLh8FBZosxMTfUkCuxU7baIizAdeAZ
HK0+BTrSeh0lGgE+6X+sD//Y88LOHop8LharBUPP7BsuPYNbGtz2e+P33E1y
E6CF2HU4Paak7vUciDJBuQ6GfDa56WhD2bzpRJeb7B8g5t5Tzpg1/qpwBr9d
S0L+567vpya4C1HDKfUWhEVGAEUvztN/i3fyZrWgFYWkjQwKIMP/n0uDjyG6
5zxj0T/pu5koYOQikKGKZY5wW1L0vwjVfIWt8QiWgTL4WotWHm41A/nBcCzX
Le6kzmlAGpWKLT6j/jubotJrcuKXxHB4F5VGzmONpMMfmzOA6OZlca94jdNT
QJKaIR7pVeKUZDI7aaX+W7NYEsNwbEetJLc8z6/HDSjagkHlpzLIdjcy/Wl4
p+AnRMDkRxz1ZjecXw/KUdkra5m1+p+0Y3/XB5tViXOtsMSbjPkI0Xsehys3
s0uFrVx8zW3OX7BH7d595tDlcV12gn/o2bzYd1+pxnGk9kAnS9nYJKAJWMpz
eDWsYUuvjEExCCFJTNXbz/OB2PVfAYvdXggsGkL2/UpRw718POZpFi1rIDdD
14bU50piWcW8RKD3QVepGqz23L6XwRZmEd4YppmO4fZrj7ws9MH2GL1+BANz
KMOLmyYYCz6Y8y8YwTsu+o1If9NubU8/cpSbRt+OS0JAj1tOYGDwN3L5B7p6
det02xzXAnQnn3TNWdNZ255GUKCqVdiRowKoO6DqUhV5p7q+wFh1gviQE5nQ
o0VLOrtWgN8ixnUqYcUio/HOYknZD5MdV/WA+jXprWzDjSZkH0+wy6LTosIO
SyzgWmJUIhRQWDwIS16iySlWVhbnUWqM8xbNZ3eNRkEgqCrQh21qbJTTBRCm
uHXhQ3UtUOmOpJZTA64mMH9W1nsLnl7D6wB0jq9Kx+HMlA4Lb30I4H3TCTZ1
OU9fZinw1Tih0hrmtw3kRX/M/0pgwZtWOJvOiQd71qVhmXov+7eLmrEScLLq
P52tnY4789woEBlU9FgDH0hhaMjgxV1pHYrcG/ZXps13/SvBqLT6vxguYEEi
nT142arV+aM1doTUnLjUYCxh7hsg+KCfthHYmQe5WVgd42tlUHLrHxJjviMm
JdvGN2yUV4Q8Q5dBwmHddWaO/SA9iB95IcZOb+cce9eHmvJ6vCzIjVorE9bG
Z8QRjhL+ELjRQATKSkNIZMkue92fR2B5eNFLpVtQ83yFk134uSURSiOdrmyQ
28wPPYdl2Z2gFaxll7SD6ZoI2kVWRXjWgbvsAOE0zWBTlk109junHAYHyllD
GAdQLFFpJc4KGntx2nHaoufXx2AUpvLU6XvURupKIy/wFQeuzmMAvKVycYCG
JiCNg8mdDgNYn0cFR9SRwN1aEGiVpTmOphIzz1fGeVWf3FkAwJpxD5/OHd+V
03EQkClGgDK/QSwpJPMUyinjuf96qW2WsABhVt8dwaFUBGtpDswPphP1LioW
2eOIp9XRT+tjURMYJBg9RzjG2m4rVYIhR64T3l/XPDzNqxvilj6H+lF54ChK
8c4uI1Cr4QzlHJx+3y/+MHIDjalzeY29iJNdtGqnXU1af+I2bSmUxJ7gZVMK
YpMjF9KodIc9px4+aRpv+KgIRte8ZRLb4X7IHMWIrvcJVmzkDsNI3d75+4V3
eH9hsmjueboBzx3UsIfZe5zLXVZJ+LcvS2T1JLVIsob/j2s2tDlVc0sreA4O
pxTjbs+Av5lE3gDhX7RzGQtLEvwl02xJo+Qe9Jlt9BaVOXT1CnQfeKz0gazh
Lqsw62uoZq6pry0lkNqVmyrQfEXyfKERqoDyw/7azwYqmpLh1TX0if2UDWrP
cj8GuMDF45MmHQU5yVP/VtubyR9Ocuoqv5LVTUjPS6YyOD4QH6z5ElNWHYNS
QZuqOovkYicxty2BWGx/TIjK4kE+bd3keWRtxVV3WGMU6pF4Lo+j+63r6oTb
pWdvaxEv0qtDcr28CY+eBJscSyDSI2sIpOEo3DwcKK+CnK76dW6Caq0trHcI
6VNxAb+baBkm+Ts1agmVKlMICsCPQrahlT9Us2U7x1AofWjq3NmMIfON46nE
8NN1tjiI3pk5A6HEwRas+f5YAP2mYox6u7f62U0wqfWk9SEcypJsQVW8Tsdd
1wRvmjBNYX6IEyAGZ3jOlKTiXxrcNPmfQ7eKnvaLH9NSNOi69+2+H9XZ59u5
RtRwtgPoCGBiaG9nG27AIEsXRxue7GynIa1TWcBiJfpFOuxMPcY1W99qaUgW
/zHvh94DxCmtk1f+tX4puMoTWPjJ01T2O0ubhqFy3jN7Kl+7ZGdZiMXMrEej
vh0Pq7xmNtc5wFa+Wnsv6CRps3xK0iieoX5q0eUt0UzcGM3YgYJD/yjA8XTl
wNFyQVIFH37PhGQO0CWnkuv04ZIuNu9gqgTE//9khdsJ0zdtINgidMYdMfJo
le4bF+jEhnbm2X8XrurlIhKFYyZy8egrerZhZZnvZ24yTlGYzCjWY6abvq2R
mk+zZE1KYbN/6YiM3aUw0+kvjgvN05Zrzi5AFwyS1I/d+qn592sW0ZY7FdRC
7hEIegk74u3StanUkLXrYJwAUub9waUsntHqRSznuO0iDBNoDeAlXBB2ymZS
JXCujtwwlqdUvrj1q6Jt7ps+VJCGtUGu5AEFcxmmR5Y8QLus0k8=

`pragma protect end_protected
