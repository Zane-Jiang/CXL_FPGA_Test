// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ES7uMd0qSD2BiTgCwmZfJykza79RDV76MpxOsrqp2Dn8YxlKZOCFEy7C45PE
0f/kHTUqzAgkRWMcDN5v7JyYIx1ZAuFSaEmAw7C2H195Ah5ES8vFXEWWqGPl
MieuiY/fnN/2si2NnlinCYujNDT78I3yycpV9tu0vNDdkCHGk9FPp+wNyREc
r77DgfxheLO9Hg1TthiTTj7SdYoH+Y6MCAt5N+MVSAfPj0NQV+KhwvpnHAca
ihT3idLeoDudWdvMnyQP0aZzo7VCIlacsUq/DR/rA3F2JwQ49+Y66hjNxt4l
vkJi2k4HIxCZxX47sUSfs26pqAT4Ia28TQ+8pInfqw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QwNltxoRl3Ra/tx9qdeoCrHo2xg3DDFdAcvkvJj9BCGeMffgg4CH+/qgcbZY
UXFQTcZLzQqlEMEaA0cXH+t5SCnd3vPtcmwpdWsSuZ943GB9NBOGIAHVRJAw
fhnrSwldRKS0zfmV4g03YzPlkQ260eOu4DaKtmpzuuF8dV4AotNAPpx+zsPO
5Qd5BIdzKEgMhfOFpv6fDZENMxIbt3wH0pSi+yBaHO8OG+UubBoPJ0j7gLDh
9WlGUh1vNEaWF+Ucy5guqjlR7jROzCUZb9crW3Pe1PUqdv1hHbxdqLPRPrOh
avJvMHal8IKM5oZuZohPYAVym/CeIgweMTVtkakWTw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
a1Egl2yJh808/BHRi+MWSAo+8AmbWfWCbGbjGZZjkqUyevw1anvaTdlxLLkP
YxYmSC9nC2e4Vaa5Lj/ovaQbxY7l0e+RnNOXx2XtKyaoG545EadTlGv5QvUq
sBPG++9QMyyMjb+30PC4iFlsrOziItHs/innPcETN9V59a85Yt7l2t5VMAQG
Mlv4+jARtkve/1t71HXabiwkWAN6F6f7GQOph6sSTV9szeY8hbqC6H2O73rP
tSdd4Ad+kGNVbLVldMa+AQUefm+eJqUG7s36J3WKXHmwgTXgu7kIwMxqE+cm
QR/et37osBsgs8gFNcLb4vQS59a6SOugvwzkEtBcFg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p86a3NAuLPWIw8wFyF4npLyk5VyyxEFAMIIKBuaUVvvfYPe+Yzn9zWjqzWaP
k2OJ89iat2znOeVz41MPsXJtXJWcFaoE+BnnDdjb2NYw2hgQmywmBzqWGPUO
Znj0OPveT3K+mNHihUirXv89jibll6O+XumsFPJnsUNhLSWhYgI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
TbAW4J2+1ejbg30OV6A49mQlqFk24yfH4OCBi8fnpK+snk/oSIxsrKivJvS8
YQcwvTMN46ybGX/a6ixPF2i/aUQvvRbkzpfcDFWjY5ScQ3yhHvkUbroTDsKu
ocnIwZYRJItjdFxXh/lUUTFzSv7dIC0EhX4oaia5KFw503HzkwgkqYThbzqD
BvZpeT6mGQ4+r+CVdh1onBmZsRb1BrhlQVxcvgVDB0b1FlPE0sKvHjVH2WmF
N/Oqhzv00zcHoE0NA+RURMJ59TDFXAnYpqkbIPF1LWW/5TF0WyWWez9ouBIf
RdCmdkagoutJovNwl9zFeuvpQB6q1P1ZFShbS61XL+krhifXTp//2ixhJeqT
dListM/b8q308tr2zWCvnruLXxxIYF5ed1AbuEfi8i+pLN9hPEmk/CvwaxEi
1XyYG7RngQFmhnx6ETer7TQ2+Nse+SO0C7hkLKvBlIad0dHdIkNWzDeZ8dRL
4DGla1gY6k5bVp9NQD4OmaY20rmb47Xy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cDlVsZ2t+28GY3mImmm4hOeolN/pxMRFH2Wm1H1uRB0T+RJvtBQ9gaNSJrL3
jFZyf9XYi9qMH0N9LfHskAxhRTHJJCSDELcuihmuSR/n+xHPeNkPwiWYI0ND
Oyloe5JKP7wtlqWKOnOPSvKyzd3lxtGES/VDHf4ZfQnCo0TwkbM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HQ795ssI5OJdQIys+saJDyp8TXYcF5hbJgxc4pYX5n26ByR8JDcBnIfEZR2M
oMnJGDrKLYiJNqf9vbwrgkdWOxmJUXSUIQv57VpaMiWaH4WNaXYfVa0o6uB8
OBY9z4If5hcOtZ9H59aHP4lUw1GCYtlUPycCVRfmjVaK1D1NFww=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1456)
`pragma protect data_block
0FW95Evw508A63MICYB/Gezn2ZKBtZgYmZHhX7zAY4H2nPL/OXil9MlN1oCj
k2ZJs6SIFLsriNCziAV9b6LVUcX1famUu2xc0mb43lp0pKWqXOyBVTh/z3Nm
TZBv8bPjp6cnGIR2EYxZjI5XOREKqHcR4spXMpIZAChsQPwgrfCIukGdEa2P
lA9y1gOFLxoeD8AfsqFn//Wv10JSm/xEy0jCOwgBfX9PQAI3qlcNZ4LmX3+A
11oKm0AsV5OPFpn2UDy5fpGJ8RQBCbpQksssS284kGww0V2IrrXno7N4QYNJ
8MwL7QiwHWeH1C5KMqvH9BPyPS437CoaIhtPVJDGDHtNqq+3Lr4Y9rfmVyGx
VS3A3Ki53nimD+QYRFHPj6KdlvLXeCJxgyWkIje1l8HMY/X+D7uSmnfeddyf
So04d2vYKuU8ECA1Cf88qoe9iHekR9Ezr1nIHVCCymtXeUsGqw+VkxHuYywu
OVMP6L82hOwdWIRYHPHt8b+mksxC2WdtfYZpVceXvPncLC1601FOZTYPSlCl
ShNNK+AXjuMulNUYBarF/d262ExMZ70jd9IUHYHHHy/kV7IEu2Hro6DMNqAE
htZYkUdXS/3GMMo9jo08joefxGwsVYc2j9I1UUroUzmKB3H2ayir5KVBeBMV
bkHzmYCWmYOCK2nlrzF8WQVWo1jztxfjXoapsihroHFRDOUU+spSX6sXps2m
0u8QSPNJS8UOa0WSxqRxmv6ADATS/ViYR/J3VTr5b4ZuvtY9uCuFmit6oyNG
Uhr5rqQ6yqkgaI3e0bA27L+oVSHprIjQhi9pSEdoUi6W6xwmMnByjUO93byc
gGhs4nSOvmeBDyTCfpfKJi6BK8RA+wK+IpYro6TirseSDiYQ8JHSM2BuHFbX
xJmJJPRk4KRGWByYPE50Rxs90tFxjPvQ16tgmR8e0Y8Z+ff1mEXMu09DMJVT
m+fFH3Ov05BFlY7hdNI+CZzzggv1YFQ1fOfIHAlBqX8AD9gOrxvN3ZODeHst
sN2ug+hMQz9HEBy+drWc6Sul4NxCT0f1xG96M6+zx44L4c4v0pUy19+Holo4
x5bYweFnV4u9bQ+E4p0I7MIEDbWJ0n5YIibW62U0tDdosDedNU6UXceol+zO
KFEBgSyDv/2A9Fg5EVOJx4suqJFnOwV8QpGXFkUz5V/iVFrnm9uxwak31aXU
c8Q7OB4odr0MDMHxmo7azhr1W9urXvu9wZVcksdNndFM+W7/3VGmo88Xy2/K
3LPfxcC+m9cVWBgAK7rN6ff1mac2rLUITfQCixMap7Vn4s5FbzEqEXgmR4Vr
ZZRr6tCJMrRrbeN8aQyZyj4CldS//6vxprzB/kFAFy/WNAbCsTJM7aNTIxdL
lnPmQNAjDR9tEaZQdWJipWF4UtOzAXfQjd6/pVcYXR74beXv2lCbQ05OhTi5
Na/WKLr0hKIb8msvAXQ7sXh7+I0fdtKiXwK07ZzSVC040/gexeOLOF0i2bmv
2QgAbGHZBMqUKY8zTr9NEHgoVE09wh+ZVjaD6UPKx5v0J2uah43Xa91nHbRf
8wdKkmrDscuQ1I6U1leuUdMniIodHAfg2woceX3ghvmhi7maBsuH7ISglygI
iDeWm24F5e0hRAfGnIbgG6YiTLSX6eQHF2MRmNn2HrcfbEFX+pgQHCHkyFOG
xTIxlVOaCnbNgUiHHD24pW4O2LzaIpann2loE1D2yE0ifUJcQ/JnHKiB+9Z/
v0K71GSCfg9xA4QOV12WqOFgX6lAFMqZbkVgMi16YssE3P15FSBu9RvcSbyP
KzuxRzwr0aiyLL/P9x4EHJ2G6P4YFadE5/sMXlLynKW45ETnJZugU2xXgmav
OjrgFN3iOzocUvRikFQk/N5fe8nhBdms3oDrfN7F3cADZOTO/wv6Dp9IDN2/
pb5Q1I7TeB/yQWWxXU7qFQ==

`pragma protect end_protected
