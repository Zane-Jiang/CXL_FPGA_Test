// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OjR+FTkLBJzQJVeTzZtYbMRRoSXRi8CHNWIU7wrbJ3jTm1xWgZfYfV114zU9
u8Kn/rPWxqNglUYRPOvOKaRz4WmeyA8dvJNDz1zmTswdw5SxemzlFOQUZtgi
2DZHNbr0qIsHX5ZtNi8l0u8r10u3hQUWF0Xs9yA9y110zk3r0hI+27HAco0L
OlWkfV0wQIu1aDiR9Uj/IsaeZAEAXwwYAdwpJEUZu0CLPXYFY2wTJS4RZ6jg
3GRvmVyFeNeZp4rPQ0oWd0RqMUpUx45uVY3zp204oZ9ggaEcV1+QZ5TbRWCP
7m3fQy7nDo5vngOw4Duw9TS47LP5wXscZZ/RfvT9Fg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
decsR4r1KH96s0KAFxQeenyBbKP60ok+sayzzorkadbRz8T8eSbIMpZQjFl8
PSDQ7BKDkXvI5enIkbxpmHGxZlApCTzKwesNTg+yXl/Se4Iz/0mCDDWHFjHp
ALW5D7TGD0WcGWoGYmlJuxoaEC5H/3JJwrogULI7pZ3peZsk495byX0FnhdV
LQufuMvh9fLdjqCRJ1SDawFVDQ2gWnQuT4z4taMG1Th+ORr1AzwBsIyJ29XH
zqWh+aYFbnFjaNWlNgXwu36k1cmi/774o0Vj8ZhgcRhKAByqnYNE67rraqe/
5r3GnwhVij7fc0BSL/4Vtlz4BVYywRcRklIlHqgY0A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KsWHsJN8fODJak7eNs2UOzHa7GFaPzFQEPsCupQvXJlnSaTs1ttjN9JrtiWv
6nxhl2hfQeHsliCCgjSozHGLm8aqq1twCTq4WHAy5aPLrsQg9OsqgOLNbRUC
xDv7rkoodQiTD5+QNk/K1dLFN9LxngroQhSD4j5GEVbhAEEERaNlHAuX+LA0
gu9mKdm8Cc0pkcgsvyD6+FHj54k0SqxDRqbuzibgD/c2BhvKz9UQg7yWpv4B
h3sXf+DppPswey/2VHzVeSYwKTF0HXJeZWniC4asGbClrmNF8dGyEoK3xFRz
YWs8J3MYNxaderf6KjThYmYxnJQq7MMo7wmMXpsKZg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Qtc0BQ4a7kszAE0MMXD5LGV3vJ7SEfylYaquahQu6CdJrryTm0+3AfRsdEj4
7QOginx/hHFNvXf9bTmorQMCs8kmzpxcn9kY6JuJc0peDUqPr6eiyGpYdFQ5
XRfzoR6mTm3mG9aymKodeeM+9T9z3J5nQRO/14d22RoTCt1PslQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nk56QFC1K1krEGu6yL2JU7M3qD8Q8s3NOubYfrOdu1VLfujHVKnkgP34b1NB
uq4rvGJZQZ601KydY6l7HHnbn0KB1oh+/vhM38+vuwRtgBT3iIbz2kNG4h5S
ois5uIHRT4/Gx1vvSseF9XLp7+NKUTh/cYv8N/obV1J8RDt8eQFhKcotAZfB
jjPo3n7zn77fnd4wX9f5Ph+fLe19cQ6FbihHAKet+3bSx4sgmP5YNebQ1aeP
cLPNcseLAfiGVglrRdVSsFpp5XxmUGaIpL2d9f7bkFC7xb+682re0+iGAaGi
e6eCoDPBBLRk6X0wMAYxTufZIprvjM9j76Mlbzh+1/FK7QoVa9jB+IpRI6VP
GLlwLAD4M76fDwgWVNxWaiZlTUkE1iwN/C7GawqAMFWWEG5QKo/5wsBWumCn
x7fHtSZX8/ybbIu9+YxTGSYM9AAFvEpfXMWXMl/kq7nNChj1h7Cse0Gq8QSB
45iVzY75IvPmsgYBlp6L77223q0vl/wM


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iQLnQs7nATo3A3RpYYGNHm4/vUqhRIDkWMY4q4sniiG5yTfD0U62VGwjzN2P
xw8YTyt0qvaF0cPk7dv0XUOmbS4sby1EKYxt9M40gTjpDrRtFl8wRjFFTdvO
/Wpl7fTVZj5fZDaJeq3Z88UzAtoXbDrHEtiMe9ImA14mmLX6oe0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hpXSDNxJopjvnaSIcKrzqzrrSWWfXVQ2FI3OcuH9MpaflJfFKY9gjaaJKJkt
H2pHk0qlDMTP1/6QmZibsGh2i0hBxn8/AgSgmdixWSDUMbzNGpj5JCvB6ryi
fa+cZvuszyHVldpY4DUqdRMjDRMnpBuXvAcv7SOCJJX2GxBF24s=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
91Nv9P/n8MQq/ry24jz+vOgXibHpI6tdPt7FchZrd0Kq2P657CcasjM0T/0M
CT6hXWTuduCqKiszlLFT8OhZ5ME5BbYAbgBl+jA+xo9XQDcAn+gEBLDUooLZ
ijxIyHc7ziuJLLSYFwAo2VtpbtbQ8LDfeOKHslY9zxwhC1DyFoLpGaEGtz8r
h72Gnd9bfc0gGoFTiNPT/2roeF2yLEOkpOxseI8+ee5BKT0cENiow2Go7Jun
Mz17xjItke+GxHHEcAtRRWE426bO9ftuT29aZSVeV0fkvcLI6tpgwzOC2Hdi
RYPn5uIZVwT/scF8Eiqbb6d+XsjMsTv9W+libxzwBVbzJoeP1BEYuwDMTUPB
ouEFRtNRh5g/w9yEVV1qD4WZID8dMj9pt3KngUkwIK0dhUR3036dM4dul6BD
Bb5QjhHC7KbrXjDsoCBozIF7em6y/j8Qy/uBbJ3QrirPcmObLKGJs6PLQXqP
VBc7tsHaTpHs1LtYcX+g8Pg4m3GL+h5Zo6+a2cLl50duASECS27YkqRm/Wrf
zjDMi78xVZMJ43eiOzugT2ymLptRZbVH530NL84r+7MHWTmdbJFm+f9jTJvE
JC5vlKV3DoesrWvS0MoTxnXc8yi+2xQmTQtNIx43y3Ki5ATkDlB51Ijv/k9C
CGHlWfpuAnUjytqfwDnfSMgBQ9CK9BBbun/jCaqGyNFMNzZMBXxTV58A4Ho/
j6U81/1ra/6KLDuF/j3B3i8oB/eNABpW2iDJMAeySw+Bui0NuWRg+RmyiGe1
aNbdf63UFo4kEWaXfGBFAveF8wAyZHMFx6Z1gRf9JtMKqzyfUtcLEibBML69
fRnzsl6DBGWZzUmx5ZN3XfuvCzN7KmQ2eTyIVc7TSJd11KpJLI9P0z10x4+I
rYydv0TXUJV4K8kY4KRtphk0gR7lEWQjw+k/6t/W/DLQ3QNTV+yo0ckwX6zI
i/4FKeRUT7hgEfp6Ax5CNVO14JEOTQnDeQBATNVcbWtsYw2i0cc/erTBgR77
mhhRjDoiA8fD4ehhOq946nslJudI6Jiwqt4t64p6Wdx+Tws5xPCxq4/583iX
7RJ7f2w8oTKvgH0L0cqCQp9olPpwVWHEVxWKZ+hjXpC0r4ZykT6qucd/hEZs
aLgwYoL3HtJE+ZEo1Wzey2mhgOBBrntSl2AiMC19SJ3LyAglyvcQASR55gif
picNxWuIQQTVGg9oQ3szRGS2g1TLhscqoowOIaoaDFimtjJeNRY+ZvZ2nW/v
cwKq+9vv8Dnnk9ZnNHZfk2crbdlLFkH+k0UhH8Gbiih/pVpC0wYS3wXvYwIb
zXidlraJswOKQ1nNhvDdfBHsqeij7rDpTsT9jOalkZhfFOlURAM3rsXgaPj2
0hCxw53Sb3hy/biLaI5rQQmM0T5A0v+MeFTY6OCs/vyB0z7ZG6BiZ/Kit+67
OyYJGKuUgdWhqBht7eFra4jm/txWo5eBAxXDuRkM4OhsRvrj8V5tAEmhH1rY
lQxy5YI/ZIlt5JRy01Fwxy886A4ewqsAq/Tu3tbQ7BRPpkbBGpf9FTmYdCqu
Z2gwIe7+gtnlSx7pBC7/BIfq4W2dRFB5i8jqK4n+5kzq5XGHsTLKclA/CL4a
hlr+S+P68yobqpCZlFEa2stiJBEyTWLObsz/ndjYpq1LdkfoP1RMYeo4WQmP
tZXrGnJrKuEHnYTLTAfQ0QrwJHg=

`pragma protect end_protected
