// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cFScMzZlhxwMHfzw9H5BltyTo+7NAJUVmlvnUTeyvlWEGyzk8ZKUS8/w4sln
WIEI7v4Hn+Ewa70JRJNGkgPTIM4cGsoMa0PQ+14AfnzKisdCEpPVpQzy+YXK
+fzrFCLz+FvBOXuXavsaTc2Ra++pJj5g6CPDq0J1FOJ3AJTaLh9BboQ0xacf
A2aDjIVoGjBLji62dERVgqlEDJFkNBmrWpKeIUDN34hSxs3b8qqi1jesTIby
jmMZ4GGbdIGkYAuoJetTjQh4cyUe61CJCdKA1DcODiGBozOAIYTebdqqN1f8
z7gtj+jNZqabC2GEJn+WZnWRtK9rTszOA3n1DiMpRQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EEuHQpdbiYfrw6RKeDexrW3PY/GAPA+k0qFBSOTdQTHBGVerQAIzNB+0DHt9
WEubCdAw0lWAx1haB7gbEV+5O3lKMzTCTM3jOr8+fdnGJ+TV9R8zcAtb/gLf
aiZ6QJOkZhtCfqmMj5QWlHY+ovqPkfbknScn6rbScht6NheQybPHsIe09eo/
RpwWR17ObA2+vFRm8sEx8JvwqTjPaNP5oew42mlLt1CnQr+ap4UlZMSyYetJ
mn1dVi9XQRxexbYHl86+/hMsvOq4LO2F12Eud+rK0ioHZs+exJrX9z4D7rRC
6GbU+D865IMQ9EqjlLkfG3hy32ORwPd56/BJLkKt0w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XqEruOCtbXUOiYzM0UGdRZBgSfZszWr5ZQIX066WYmX6AGUgpQKa+rDE2AS8
VN4oVlcNhjimAXv+QC3fnE2FPz72mDtcQGmWyYXZ20GUEYOWtIiRJqCWb5hx
OEuxzygNYqC/Llegq80JkHdTE4HlEE+U3xG4BKbUygmIYRV2SVP5/lCFxp0z
6P3E4muVNIG0WLr2FvEMVuSShgGiqlLAAnM2uZ0sIeMBFcwt8X1cILPAIXsp
ptxfsH+0G59W3yX4KovpEi1tFqao9Xy6zCLE68babR/1lNdZr/O2mQ/ueg9q
/lISzBuURF3Jy186gd/39jKITWe3PnMSkTK2SE4DWg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WYCdvnKl3hEkV7FZf4KzTXOJqAzgcXajLYhd2n8jF/qYHaw6YkK+M9F+KlJ1
F31kSqdV8KXurajoimcyFnMJlXaolmRjZLc+HyVySFScEckQemx2Rk1Di9hR
nejgpnra7mrrxnEbyD7acI9QgGcRvDfPfHVQ/kzJBm3RamA745I=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Si2ZaX1zgribmWd1bVT68OzRmtKrGMtpcugXgyzkgkYhn/Q5oIeeFsP3/9Lt
IifqKrfk4xYFf/mY8Imy+SAYQMC7oBxdh9QUOMu7YFeiTQmSpN+6Ilib/HDu
8ka19M/Cl++dbBLKZ7clOvA5J755nOvlUU0jsqh2WKAt24s9Z07UKDN/wABs
qKcIAwg7jfpLC9P/GiM04hpobeWcqo02fWuiPEMns/BpoHBAbqvDcrdryoaI
0QNo8pxVIq1lTPZrJcqS8PacHMLr3fVlP0b/fL9MWaNtbeIMOwEB6XJ5e+X6
Kb0Hf8FKm4x0qQIgvQuCvZZd08Wfchx+o4W4Y5THWrSu8jFt/sPMmDjjJR80
qsGaKDuYRf5rq9qFUQUlw4lOHJhJnAau7TvFdDa8iySfiRm+SFxCbpPnIoum
GT44r/umi60XOjNtV8FZfEIJ0E+slkeNkBzrjFEXJwrB3aGY6VrxgWYTxyp6
DqcnIb45CG9s7UK7ENbdm9axgm6PtY1q


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OZMKhKzyL0cGm8TnY6Zy8uUAbU8yR3RM4UMfoPokMSq6l5VFSkC8NZg+hMjx
tzwZIEZfqPWnWU61QypsAi1NqhwYY+LIfQ3JPGGEGsNzPmMkBNbP/vzujA03
8UHgFD0jY1RmNfArM4Mdih4xhJWk/U5mft3DpMuyhEHfwYXGYgk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HVAY/ZZa6hBLO7ppIpq0tGdGPdsipXJZgq+lY674xYcaxu3iH9xh9a/2jGZ0
W4yfmgdxomSwW0lz7T249PmBeMelyEum4NJzhl8vjKy9ZFm/ID1Hwrmit4yB
OFtbegX47NtL3REn8guUurpJXzfQuO6RZgv7Hs7xLEASgagmAo4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10128)
`pragma protect data_block
AskDQegkbSynPhQPKavC4rpMJWjsO0+5CNF6tySSfMmgwWswBeMhza+MQEzP
ZxcRNVXAVA/Ip0jXLgM/KYTUsyVK2+Ox1VG35kQ+BB2Vqud/29lmVJy1AlUK
UmPoNg1OYKp5eYqMz1Hc+eyvT003PLrsudxLMxDEnGWnrVZWY11y4TQJ2Cyo
LwMaHvS3xgnUfE8mx2jpgQGm/9R1zmmmBN5D51xZbigDhno68aax3TNpfRXn
clQtF4M/jEmEqA5qK76sYXbku5QqNB7JZ/6Uv/YTDZ/90Y1q0cU5GA9joJcM
jcbKx4NzTjvS6NWhyYRHWRDiilEZA4c/wG7TjZGYrh/RwzotV1MmrBNFu8rA
KjFTiJkUYyvAMPNBIA/IsW1d1V0eriqigDej2pUZnsjGX1k/X6ShgMfh9qTh
SthwFNuvG+rkBJpHyzSc1dwxFw+FV1hf0ZmhhYNbKLpx6N7kUx7wu0QDTthO
jBUj3nK8zfM4a9Ha8eaVoKrbZc2VXzuslTVSZFt3n4iR6niiYco8rS/fMpAR
uQTCVOiS77Vc81tMjATAzTlFSEwHC67OkN0GEp2UYXworwyar20yPg0s1lrc
C6ijTc0W4XUfi2ancyFyJ5zAkB890u7uODlmr15g+PaYp8dsu7auuo57uw6h
qjhBI+QvtEKNRqa+oyWTASkTvuJj2Mw5NJ2wg9t/Z6GlstdS0RokzRo3LbG2
2l/KGuYJPaSoKjnrL+1IH0P4qcE0ZjeMneb2rhWh/mgomU9MDJjfCQwcaY38
N86asyOqs0lOIdPgzATjLZh8qz6J0ZaASYuiATzykTx90oKAzbNjnDwamorw
qUUJO6Kq5Dew/PiI6TmwuQx6rlaIp4TagmjgUaPjvMSec8NccNaXIXdPRRWv
eCHVT/uEoBWoEUaxtB940g18ZiF2gQepwikh1uVlPAGiwy4VDqiEURFQcP/Y
RYQvbSg+UxqJ70b6Z+p0uecRgpy/ZfVyZgPnYpqv/Ycy50ThI2zg9sF7l7np
wnubWVZLaaVY3dyYHKdIfAeG7koe6KxVwxIWr/9ewwm2NBbBYIxUJh/G7oph
odQw2KfW/T2b0dyDW46SJuaNDJjWP0XKeNN836YRElrID5bHApZPX5JdG87E
VN/b8DRPe7YCReXAgfAgzyvXKSMbcxArU8ZeXT9wG6/1OkWq39Mxpz4mrTFS
OoTmTI+cdKqVE9o0cVE5nlC7BqHRW8aLQC+7NFleuczJboebWMl7Vy7QwxkW
l0eYRT9++nVYVjctWPvKhYqHUvAIfPpeEcmb8RleKu/AqguEyoa7Qpbz2CK2
qED2lr4SSYT0WZhB6QJd1yiZ1z9ckWwfpK3IleB7SwOAlglUqpc4LF/wotul
8QkFUZ6hF0ePWtnrmmj6cBGg4zOXaWs85gMqffKzFZRb67BueqdrK3nbggdV
vG5IF1qdHQ0J74yxvGGicpoyeVc0o+znEHYPKSKXi1vr68wjMifIfTGTRZZH
hicqubyR8ZqBjOYw1g2TK3o3edZvXjVCQOIpsihKnPpTfhqeKuvQlTx1ZZGy
0j7SiBQ75B1zc0n2M2QF2FFSH1OJgL3suPsFpyUmfWrzcOjA9Uw25IFHXK3i
Bj1ljr/5x4NnzXB/bItN9f7OCk5psPdVpbVgkGZEl+MIyYK9IlFN0YOQTp+B
8yrc39LDZH9gnrWYvYBiaHjK3B1we0MUtbiupydovs3QuWQ9rpO88Si9QpRx
AjJlxOsRf47LI/fYzXHxN8wgzALdqwUQwqIXSFtlDNe8NCpvTvJIvM1mDQ2s
KKMbj9GMatB0tPj7jPoBBS8AzauQfZBWXhMZMwOMApa0bRh4Kwf/Ov9bnDqL
LBKsRx6eF+N+8fQ6kokyrcpQTvsYfq6hmjYT5SuPn0Y3T5eVW+OPEeUeVYyV
/uM7JFGN4IJ/pJkrdPL3mlXevD9e0QvzWCD2BybgxXMFBe3uIKZUj/Rh06l6
w7NIPLxa2QbZwOSRyj8xq6XeXJ/9znnMk3q5y+2hQeLBErFoTNaByI5r1XtP
NtkqnQU00aO19Ij75//OrVU1MunZP0VtJSh90dYRMsxS+pyGL2zK0h+P7NaI
deek811vM3VgJ61UfLP3E5xwhf3qEteUAgfy7ufz4ck127xfHdcK2UUAwqYn
rFIBNSGtWAhbmibe+w4nW6ieslkIKdWaFB2WPcisM7QZPDe9DetrIyo0/mjP
L5ahCN5TM1GQsAJFzbLxh3CA4N9HCGIlKg22hO56wPHMDDu1cvbGF49gcf99
ZBR6HiXRdm86n9N6eeXIvu+Qdjrxq13AsraPLqjDfZppUEIkLegi801/csx4
8YaOft0d8X1pQys+8B/qS3kHk0hM3R73+cPcYo4t6xhDxyBqePa35s1Decqn
y2nHc7EkxGbU+tqFRf0jZb1gAmHlzRrqJTjGP/sfpuWLWDVchs01W5sCaavK
PM29BtELPzSdhienlSfcc8elKzc+SgMOuS7tC6/NiAEy0AqGCGG742Q1vHQI
X4Kw24I1wiysfLDySDot43B40K9wUwaVOVuwut5ZlEgTP3hWci98/CJpWuzy
W60gTN2CYXsgqkgE0A8ckTKbJilZ8l8Z+JKO0WtEh+26aQUimV8hxZ/NYDp9
stIh/ozgrKqg7r9BUTzQVR3U4EgxKHYBP0W0FRdaLiVoQFE/YRRJfRT3rbja
EAG9XQvEmCtn3G9yHMYpz0DCOL3fqMkW0c4BO4GmBJxakitCZYQ74FTzUgyu
CcuD03iCjigUPezQFXAH6k/cJY8D48BaFqFrQ1OZn3EkqbgNtOIygRVGf/lS
I/4XSZp2wCSG21kt5lccxmdS3DfikdDVl8WE64cIa1Aoda+h1pFNCR2+rb8Z
9ISTmktf2tgCVXWAzI9uMf8JiZWhTDhwy3b6KRBtzsWwBSIGxRceXdJw6/Yj
Pf9Ft7v4mr+MGVhcddXfFAYTlO2EkURQsyQcCsk+t4M/CWUVM9+eeFLLyW8K
2rymoDNWbq2ZKYPvKWAVC5vT8CrXGjTRJVqVLayVGpbUPm4uerP0IWlpigNr
ngaXhZw4wcj8qvCn9GACcBZp3GDUBnDOJ5AlCeWAlx1DO7eBTO2MYHyDii/m
WJb7d4YyN5L7dlIa4zvj8zL/WSJ/A67zWD4LtyqmPN5O9KdAsiWobd55iaRL
KRhymW9uDJ5UTCHaF8IE2DSeE5U+R61Gc5wl1m98poyfIkSbuW4r1gA5iJrr
YIvlLeIBQ1WYLlQYP/+TLw1b6kSMH7cEhAMiafztOeIKq2ligSu/hrT1HLEA
2ewnablQJiHX4gYgmb/VxofWpIXy7flvT2qeNZaQlgSUlG+EDCxfDhMW97BW
s2hCY3FOO8uZpDL5E0DrXKbAvwz1zHejDjXETWro1JoK61BdDnuzkk0eh1/m
VRJjm0B6bUz7p9d5uWII12IoRjKqB9PRYnLN+7zrNQjxMb2iTwr3KEfEjLEN
n6VtKGMH2yeQCtaUus0YFgsIU2cHWD4LuBChA3sab/vlf+nURaLCkIFM/gHT
Ra96Jf+zz1cmzSjDpQ9X42eaCQhm1anNCGLEd6glOpf+CbRGNLMoJ2oDJbAz
vmabKs2/iKEFGLhIA79ZUr0iynjeZefe8oqnwATgny7OE+9bpDCNR0tX0Wvl
YOkPnOR2+rVOLvNxe6R9f13KReIUsLwnVZsiRHvKpkhuygPbutgch4J0bMox
y1atzPIb4nsTsYZSASBJcWElvkTijLQek+8vUp0MWkqlFtBVixRSlkMSUenu
G2O8qUyQX5QYKVd6R7PX5FFQ5pbcuTewPJ3ejkX/rqydgKGr56lp5x5MqmYA
ApEPteVxeJtKWTlXEXfQh4dBTemadR9uuFiLOhR3oMEzc0zulgH71MrV1ROy
PqTrBtP+3fi1nTGNTxAW+I3EwRGEiLDo8iDajMpdJuDXHf5rfX6iByKS+G57
pnvKNFOyN/8QPOFWf2SziLMsime+ls6Fj5HBEwyP4YMbbIAPrD8EnzGUMuX6
1/dQK2HjzhCy9YE+tBJ9igoZJXPnn/Z2ASxt3cVM/6EMr2mUF80oUthVxJPv
amhozqE4YubivrTen4guzUSLZFVwGSAkpqNsl84PWrlX+nxVTrAeJ7+RtHeQ
Ti1y49i8QD7gF5uO7obhCOwqMJDFytWmNt2EmvP3o6UTd5l3MoeiUsvK/6I2
XpAtd1q2Lsma1D09MwMJhQloZyIFev33NG4YXuZyp4lxRUzK2FkSC11ua1Ul
G4rzi6HkfJ50NWHdfKL1KzwRWyeeKW6N8W5MWCTpHf6AIl62X0WsETQvXe3r
pY08yvoRruZlpBtJEB68jYAG484vwc4BC2sf0PQVZpG22w7a8nHGK2vxkeGO
CeOOjYLjJOymkrX4gQuY7EhAwlYSsnSnTxmQJFRJC1Tc/V3SVmos14+hroTI
I9LqNufvC8jQcHwdfdKTwNu8tPQBxy9qNh0SjvpkxNw1f5MylV1oSS41hLn8
9YqxXMDPSK0//qPUlBwqptWgSD8a/NbXyG/+svf+Urd0bfYhr0NpoqxdTFDC
k8lFxxtx5RyBiPCv3B6nfPLS8nWEjcuKRTb+66RoEe7iZAtTWjU3wYoY9Pso
2piD4sB10K6D/bl+IbtkI4M5TxV/U9SGgkaHIZOFm67unMPSW2cwDSP1ZfYj
SEGEha8KVdJrktJw9l8AJwWj0iwglbnnGwUFKwnPNc/z2YuDvLXRKfrs0ZkP
3ZPQExQBiH5Z31ku2CKHy4CwT23H2M6aw8rdBB2kHSrPVze8Fg4M5lbBvc2F
5KAqISlESLo2GWDDttWROnaZoir9rCDfqBlkQBBFGnM4dICidJ0vrqSN1RX8
zfnnO7KK3ysRjmBZExn9L3AxYAl27ST3DU0qJnOQNaX/ogBQp2C5ztRsaFBx
vqgWrdUM71nN4H1c62d9W8SSc7kwKSd6DRFFPPBz/gtDCz5T2H7o0LTMOy2N
nBnNhjqjW93Q1FT4sWfnwyNTEW96/m0neV7zTSQAREYA7rVOp7XmKioatzhX
lbD3T17iwKMLprA/qVMKaxYFmskkgmOk0TrW7ENkQoJVqBHLqY/rVEGMKDfW
uLnn4kVbmPpJ+Y7FC2WYlFq8LhCJ1BQrGNGGkw5ISF72B0p8pJYMmIdqyvhD
Ja7nnj3QA+BuLZdzUm+jXYoQdyVDNKMoVZYSTBlgzwePA/27Gvpujjv3ssbd
ENkew1VhYyr6Vqxrp0K96FrryCleaNrYU9VltuNt8cBBuE8lrfjGZoGWqqwO
NUzABeOiTZQm3HIYcr37zx2xY93CQKf8L3tIBH3pFkhpqvNHCtqNZzaXjwlg
3MGQWbGL4k8odqAOkRVy1culJAeL5KcjEKEYHyKIt3zLdj6/+kKzLuOMqnyc
md3ZQrn+eTGcvmXQ8nD2cy0zShKK87+5HjtIx1oPnzgPP/t5k21SSqBnAWtw
yoY1GW0ZK+1G9rKV6BcfzMgSNKIiElAUe4aydneNia9olQIUCfMzNYQPQnbP
o76+4Ctoi0SD52CH5mc6apFyngYlNGusJ3OskQCD0K6EdG9WyfwypEDk/Llb
cQJZhmNHNMEHkOV0dOmMFiWZ2DHZjxiTw/VZPpnJ9gc9O5PM3e+g88GRdBmG
vFSpIeFpmnV68B5nuycWKj4vcvm1qVjVISsOhHBzP1PEr6ObIZHJX5li5LvM
JfdEZIxiEMPk92bDKVv4VVQXrrG+IcXhCl2pgJfFws8Ij9pdxfiHQ44Q1OeP
DNGM8ZP9JpZhfLee7mXM1Vv8kGqE3MmQALiyH2pZyQKIfAxbK9LaAizpUsDZ
ox4vR2d4uOjDRHSgd63fVGSmZ8UV0WrMzzxYQ4iUE9PM1/fH6ad7lUp+SbSI
jkechMIhYbz/5nKlrytRPOKOhbSsrVYEdydUjAVnNt2BX/xjUBdC3SompHGM
Mv7GdgMuNrZnSUCTp9Gd9M9R5VOrUjc1vd+kbi+8yuRjnVD7UbH+8XXVkC2q
5EBCAXjPabfj6M3BuosJUy8iDgELtJxc0QiMsGnP/pdA4mmEbb7r77GRDMsy
Dw0lPwyb4HNqx7PMbOA68vNbiZWPGeFrYmfGYUB32EXtUmVz6nLzSkwjWiNL
J+T6pEs3UcOjHBpeA01p9NolI9Uqld2fBbAMhcEtlqEh81sJx0P2D/fwLZrc
j2iY1qKZsRD1Iw5EgJbeLV+7JKJ/DqWWQa486FU9i7gdwIZiVZbP0J6YzU2o
+Z1PtAaMiyhiYiHkSgoNrtEL11Fp92G0d8ZFoczvhZl+C+eFPmFW44NzkvZ0
WRP6mm7RY7xzmS7HI4jABhmw2pZWzD8zCDmso2YnjV7v4KwyG8A2fx5DAGmk
eDP9z/vbJTv4/9DaSpttHiVXe6Cbd2kFMy453H15IL9j6gCaljnd+7wSGPg1
EPFDg/em/K6UERc276kY7tKLr5g3LySTk6hdh1Vb/VtJNcoudOkLzQFAqo8Q
x2fpCHwgrEUVI80wz+W/IRsIW/ldtMEnmTgU++4Ievj6qOYCz3wgdIH6Dg59
ykuebnlR0BjLOulGJ+/SFc9gFz/pnRS+dZh6FXlmABn8OBZ86yDze3Y9/RFT
yAMkWTmDgNV1f0ZtyoJrdeq+AzqWTKYNHzloLbfT1RFWqVyIypnUyeI2ofy7
n+FWJV0JEoXHZSb5Smfj3RVyyQFFRGEmClb44PH1zTadbibFsXOd/soPRW4o
92jhEVrcosCzLgwSBAm6yuu1TuuDExVOXnWS1WPFkVnFsltTxTlgKl0wWJCX
ARrhf8j0CwsxQ/s9LED3KE8v2Tr4noDbCSzPGbQDCS+N1YDF4QV6kRftNImV
IgS2bM6jf48QlCXywPr5n/6uMLwn7gFBQ+i7P+6Mx2T8kkXb+5easuUvFaJa
HZnBwzj4/T2E+IUR21mei1PQnwk2LfZ1J4wnz4MQgxpr1tUgk4P1yWLxbWrL
pU8OPZbVMlR8ZGixsANbkUPHjATDjHUAFQ7H+veo2zGRCgAUw6VwOKmiFcvB
5OGI+5roBbv8rYEhcZ+NtLkU3UdUcDeMB/27SKF0AgWWwoJgeKYKP+92ukFl
fQQhdPlhGu0M+UvhVUcPrHgPsWefIzvG79yeia0JuO+WuZRTM5CphR6t9esd
exBPHN5fAD4DhDMACStbtn6VutSjXlcWT/fCyMAYnr0+NevVsDMtz0fTAzna
dwoTZ61vopPRZQ4mRYXJdU3ol0c1dkAYejDZq95dYCPFhX9VaK2A2vK9J46c
zOBZmzexyIbcOaTIyJRRPNN2xegJatfTA8DPMSL4Tzdy5fbk8pTh3+n5KiDb
Ms7VXEdzu+mNeyPVk7dv9lTzsH9ss5qTFwJlJ6DmOzjEIyuhiwQiB41Hdkjk
qtpdCC0L9yIasE4PcbEbKHHDwrUcIA9q0rMuKQ+y0KHZ9mhBaEq64V87zI7i
K/83ohBMp0aVM5qDehsIcjpO3DhPBzax8Beo4AxS9ofUcCqvh2+waNHFo7go
03d33DVk0gDlCjAXkVf3F70vrunAl5tNlMtiuzpfgBAEstxVxwjOZKmtfiw6
vG7xQ/C24qevIlM7L42vYTGlMivhcAJM9tzXTUoH3ixjhZF0MBZqOe14G0w8
NvUmYb0SGFSb/mGAeULjJpJMIKSbSsa6at+aa4Fvh1AbfAB2qCXT/CWnadoG
/voTmTyNIGNNklyJp2i1i7UApakF4U8xD97+Ea4NU3hfoFgYzazZf1TACZrm
Zhn6ELQ+RQuXq4qrRQ/54fxS2QCaEw+QHD7Cixk2Gnx+yOZiLx7qLw44PiVp
5NPprEzB0Jza/FjZ7Hb7HJbdpKyKnlM6LCvAPkK1AlPdz7aCdhL2WURmNerC
zLFtpm0Aiv4zLsVTKVBEdAWZ4/piAxCvMOlEKSl0oFSuxTsGXX1rXX6QjCBg
aZGiG3Ixa1UJzrR5Q3+TRX1b19qx/YaoBK2/1KNpyV8OtyeromF7I6xGy8PZ
73UPANtmZqg4ieiKS86+AEvyPHUEecNwm5XMLRAABUt3ke0T6NF794BLMHX8
aDc3VSeVZEa3++jAl0sLKxvsY5z8YW8Yql3WmpYb7UlaTMCLeS2B3l/T2yMH
857jrGJZAmTmJrZZI4VN6zHOf6mpYmReP1dcooO1MXAyuxsQTwAUTFU9I4s6
sxL0vCw8b7+GQxRL7xlEKzlSEq3zJxCOMscI7WhNzIyR4bLI6SN56UiOwH/Q
p+2OTlvCNDVrQfwmB9WLmQBXTsvXSoDjIPeolob54aZqbqNxUCE+EeCzXCPM
hqTOEG9/D+N/lcn+x6BaiR8BknxPVNghxJbsL5t7O9yqBqQbp663BYnyXUhf
xG78Vii6GT2JGdZxYVTDyV4xHIHrjvFAGkzqrz5bnMYrs+BrBozJAs34rZhX
Xo5AJ8H/ZAO3c0LrusshHqwJx4WFyg8obbE+KKb8Q1xpzxfzm0RUO8e4l0Ia
7k69vUGy6xZuij5X7cobFvm4H/anfHQefI+WGNBaP6SkRJ7e2jVmDpEwqHxy
6xW4pgKV7VXbk/gptlifh0jo7swb2XrdgG76efF47fXuP2QPZsiiclWVaELn
8w3ralisVDylezJzTgjaFig2JG82XY6+MtYNIgRaEZVeiGnDT3y36b1HD50d
ObKGYiE+gnUNJ7B4UxcFw9bUWFmLCldU7OlBQ/sSkSsyCYQJP/aa+33SQ5ne
KQP5SJbBeK9+4/YqHj8iw75nfn+R74SSU7GVInX3TNqU9x9FYIl5Fp6Pcatr
e0BnT3Mpo4bqK534wAb3/pYaavUfmlVscboJ0EfJJZmoFH0qj/3uyrECF9Xg
uWwmIYBuvuRICRMYLjkaDNSDzEb6gd3LtB6ccCo8qjftEK25Sl1GK/v7cmb9
V6/Mi1nd8JtOKzvLFiL0EDs+NEf3nWh9FX3b/BYajFm/yIf6ujUMEN+nfy8H
UV63A3RTDanWaOMMXy6Ta7+Q8CdGDBEyEdY/83IUxfCtg1FCbn1yIrJS4s6M
zPkgTZX9IMgLF7GQjU5zq2f84bhEZlIMXd3peGWAbHVKiunT0kQcklzt+hWW
4LFNcwOpSGrvqxM64cTY+u9MJoy0A0YU7jWfFWs6iX8IB/o1mH6JWnyh7xqA
RpGUFtS4thv93Y9o26vQoEWsf/s5bT2aGBIW5dyjTypIoi6q08qjudz7AXIs
jGq4AlXMYdHFBF2m0Mzvn4hYahwd8p1yvc4ftN2o2Dlubssq0+OpFErQS11d
bVCXV09atLfRgqxyESqNFDsJDl5KsG1oS8i9C9ZkWAOKl3Da3qBm6GjENPPw
GMccb8uGrfwzPLO8xiEhJINMVEY4ZgYIofXqfZLYPAtMGqv7EN1DmKOJXvGm
CJMMaUSSymtfRK0siArJJpjaIf+KhDTqvV2H/esRNvbxAMfWTCMAASnkohBK
IWaBiG2KckKHXaiJ4bNAXEKQ38sOXYQ81WnMvm3ssKXAfddEE4hYkhNGCsPq
xiUw0NPy9RbBMqP4O1UQ+G2eAhF9R1nmhRUp9OBaWIIP7Ewu+bk0ZlsT+aVA
jQsmbOnGP/QuvkXsdu+qew8mglic9Tyslhp7t1k6QGzDyq0yJyaRQHcF+qfL
bzuI0kj/hQTrci5xC6x1WaD8kb/x81ZfJ04TJw5Fr9QNRFhVdvg9n5ed3bec
QIVAAPSGYDxZ2o//21VxCZSJwKD4yoQkb068GmiH1Fx+wfpIxM6amGcXK4EG
FwdDd6+D5Ht90m9ZoLzXibfKsSRYiSG4FnCSaQGX+sgz3G74V4DldZSouiTi
KWI7JDmVL5dew2rkYvC4+ARhG6/j28A6NoxB9nY9TEBG0QFq5flW5Uu8DcKG
TmeTO3DLQ0wGXaIb5455rThUheNYWlIPGTFsWWkB+X0KR0hqcVl6hxfxA5Ab
t8be1jSVJJhDvYc/TolRz1g9jT/1HOywaGOmb65PL7Cc7yo0bgclJJHpYkRP
iwKqqRrwyF5+EVWJVWNedK5ES0iRRT9uWCxoPcgVCQroZFa3lBS/nkcWrahx
rQqxVVOxOyblYBdErM1MND/epFx3nDdW8odC85PWZ7RMzaHQDTMglfwmlpG+
trd0FKcsEoTv5J4hzeauK8UsX7FLABuSJPy/5KlKT6Ov9ASdFMO/ajV0mrvG
dVNRNVQFOVwDsb0OgUAsTajoW/3VQZ4y0VOD0fz/MoHJUV3CGZcjnJu3JlYR
cEXBKjUiIx8bHuPjWUMEWDsLQefLMoHxnemwN1x1xGkrOw8QU1joY6tfLr5B
KSqOCHlgB1MW8lsk1CDNDhgYqQBWPpO4qgF2NGCd+uKYpHAxJ17mEwZ7/yE8
Hy/RIMcgX7vityp6MWgXk0uJ5vX6QxJzUfdRHWLxCYKNMmkTtlHwk3PgTgp7
gWh02bBbAMTOcrmf6soNkHtlthd+xthnWh9MylOVarGUpRaJIKaIiWbMmY8/
TrcDcyUXrufBQntS38b5Uc20YRkWKMQLDktJr+h7Syk37gJC3YuTLYRUxxsT
+3Mx9z141QZI0/9WTiFk+eVW4WAcTEstCSVpecQXJRGwTATmqXhRrD7x227x
gpYoTHmyNyHZaaZZv9pI05wIiuqIrBp3hDHpexW59pPEonB2Z3uUp3so9QEB
jdRmUGb/2Ka6/3waINWYDV34TfqBC0spU8h6NadyasTSfuHCBaJ4yGmgHyY7
U1AQBvjl+AEjts5GjYzPO7jxLzvL5J4AU6KMbxLn88onKxxWdw+64eLdSSup
5oxFzlbyqTWyFTNeyhMiFMcgZC2NTNVayzrI01EBmTNRDq3U5cnEET78kf5A
ypBqNaPC+XB6BTNFr19ZVkITC21ouOBc1TDZ+3gsdVrzLP6npBZ6Y8VznA34
gya2dNtqZtAmKL3jKKZ3090Y8Hy1gxWsLy/g+6dBcxf9wkFzEY8jbDYZGgL4
oH/wBBBCv03DiJVlesMXhiKhJP9v73Aet4slFysNWJ+3lUK62ndc6lBE7SoR
Eh/2wdMLP1o0f8jDPD2NENrHni8ekpbkbND51mQ8F84auIqzJBsvS94qH+wF
87ulm+L0cUYQ1nKCD69CyF0T8AQ4Wwa4iZaBO25EjlWiL2Nc3doOZDvvZjtT
V4HNndlC/Hg9QLsybu2zUrVLxhgu0yhwlgb4awkNbHl3rOk/3ot5Rqx9VFxa
ipLRF88A90UkBklme7TDBT91UYAncnMUdVQrPEuW8+UQANszjvfnekjwf47p
vQLMfyVOoshJXERZ1g9xNRzTvohFtsF5SZzylphqZC+HUrlE4jrE2pw7HOSI
pdJKflpBkimYhAIOGXYaAYHCNd6/SMWIa7MUeJVZGegUzRr+9OPRJbnQ/H0g
nrWSYTNxq21Bp41VCOCWVMNUr4dF3CAjHu4aZV5jnRofO+fJrt7Sv3gB1Ez2
xsvZqrJSbGFvsLRUQrT+D1sZmXSiLUqa4SlUfvOohFe0ZO2zaH0+XbrpQ2Ua
ZFxqhuXDGzD0O4+eqsZR0lkuNufXxsKvh64Aw0i4puGuUZ2GfVmJwU3m5BRF
GazWmofI0QKckIbPYcbVyqN7DTpaYlW2vnYKuNgaCq262IKGv2U9/0zSZlD6
Vx+UGIeIw4bqgwzx7sVKsuwMcCdkP+d0AYJDLftyBFE7OoH5DcDa86zHOZxA
vwAUlYJRr+eSga6TysRG1sbh+LOdTSsDfy/lSergU16wlxvnUWF9M+9XKm3c
21x3y+KkF8HBqKk8MpkOWTROfT3plDP+L+1hcUcKQhCWLlKPIc2ZXkyAuvXi
INdxf+upbMuoqhmlBUEx/kFRuR1c677CISXacPX/0D6OjimUx6wXjkxCRztH
EmWduBgAxnpE9Q3rwC1bxXh1eCOg+4aiTnjWGe/RYO57/3OXrxoI5Xk5zuxh
qC9FD/45pk60VUHEONjz8NeNpsjh3Y94ZiR1OEaXyKgGOi698+Ht1bKa59Hi
UctxeRzYhscQGSqOn/xgqNbA7YCuNxLz8uidlEpA4vs1x0Fc3hzNs8+DiFfr
zccDZUTuUlqfp84o0NYmenOIOzfHKTRfyr8RtB4D2zf6ZA3HP9BGN53Op3ge
Pl3RF61L6yiiPKX/H1x4nwhhJeeFZTZkh0bYxi3eCi9dj+xjDo04XDfIc9rH
o7/BLmTPUSA4vZMARjrDhuTGhI9bA/skp4ZLoSlyre5aN3/ZIogh1z1G55nC
eoKZus5IimG5GgP9Q2gZt3ffwFizLj2HSyoAPYmiiKYZ5bm3QFqzrAo4ozNO
zGBngoXLlxn1I/Igtwgsebf+s63KSKs5PibP0UhznBd/zbEn5hIRXFBXQwOK
DkusSWxQc+q0tOeXMcjo1Cj8rJiGKEW5o1FH23eNOAb3r28AZY38uLpXZq8f
zGtQJ0YEoqJzyVFNQkxJVp2f77oR2YBnTIMP46vkkB+8LhF2Kb+B3bqoI/X+
6yTNtAgs7Rkjt05dGrkP4JWAAb5+mO3cKWKvjLsFr5lye7YESZXzXvSVsGAk
ihYT37BWsnDE0r01/WH3iKcHsvRuGgZ2gOoUXJhx/zdwi7SfGg6Xf7O//mb6
weCm+c5DWh529wFdyH/DgUxPDVX6UhgQ8IwTLi+OgU95iLoiGn1pjuYGXXdW
PEFpHwd+xjK3jAvGbux76MVW5gALQrQqHiCNYrEaoaDqSfZtQ0Stcu7GuoRv
jwrRk71n5cKN1yBnxaW7dRuca3KFA6mt8ut2oIvNUQRgKQEu8KlRYkWH/eCb
71bYh3+VC8r9iCSrmfvK9Qv75NMaLr7iHq6m8nECCnshfKzob30vSpW/Ap3T
b5TtBFDjSKKl2pZ/I4XDl0xCIXhNewb1NP0T4nN71HdsLSeYo0igdUR+Kohm
jTJZtfc1UDapHFwh8NqPrMDD/wX7viaDZXLmubK7C6pJ0U02ZOReEVDuOYvz
Q4MAP+W0vqwtXpxRzGVH+3ZR5LZ5YyUe0ybNrK0DgnfH6QTpq+IVuQOYro91
0gFig07K+u7732uqjPaAUDqDQtQBf9otHIjILRBWU4n6XsLcuEjMcFnawMTa
ZePHxCkHFT7Lt8rDO7UPdISvix0vyCkOl+Wdu9r5r911lJm/+jlA92Q6W9KR
QKRAy13SYbTvSthmdIYqZN1z6Ev/jFaUKVTw5uqxeI6ylLqcnb10AewqTNYE
Y/hCcQERxiplTM3zRzhzfq6EY9WYa61uMhAAtg1UDieVzMmifE14sjvoWTpE
rWFq6IcrC8lynPxwqh4gqfy5Tk2Hb3aaBXxsctAd3cS7/86GVPcZa171SSke
VCCRIe4lP1ooHD+HMqsrlOvP83TPOMV3gQpKzwAMPto5oUZq+P8GQVwmHaFe
Dr3JOZTwnJVJTLeqodhNB13WkzaGdnWiG18NZjqdb6ckudEqjy+5MUV6vAcR
1MLS4YoGvb3ShfvuClnAh2zxKgu4D+MzAQ7q2ckfjgzn8t3dviP3uFEoaFy8
PMjJuiapCKaRYLFJ4NbUahytxaqKH4YKgFQzDiZxI8d0e9AyC8U/cvqubPu0
wzvE

`pragma protect end_protected
