// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
iG9ksMdivO1d94PB4urD4A/lwc6kNRgqJVEaKCEvC5ub4YId9PeE5avZhkHme/31
T4Hcn2oRMJoZ5TKeBZh47kNOZo0MQcm2eNcdNX58e2DbILwzt3YZoOvmIyZUQLeR
7c0NerjSkuYzq3lw1sKhFOJ49TU0o6bnyrteHZPAW+k68j1CHDBRqw==
//pragma protect end_key_block
//pragma protect digest_block
zPKNxw00hCK+9GM3hwifeJV+4hc=
//pragma protect end_digest_block
//pragma protect data_block
t8qizigT4aMf6tAoeYSpbaeclqk0cQUVixptkaye9Vg96KVxFwD182kfZQBqfy+H
sb0qgIgnWAe67vZHnZ5IgZO9lkn2EECOKo6MrL5gXJUyd8S0CiP/8+0PAlsR5nUI
OHXo8AYleNoTgbdEBsJX2Kb1lNPZOLfLg91x5WYpjtIbKMh++o1Sih7TL1jS0wJA
UF/XwLdnCimkPMwxvAwTunIW2yVHdC4/SZfkJp7S2BBsDcH3Hp5iVLQJ1a3mhGqQ
hPnF2D+Sylf/yfeh7IUU4ZllhUDemKuHIxDubyeAZydl6B36tM2vFZaAbIdGqlGu
segihdGUiCc2CM/JXbaNji/q7jkhGhK/FpbLbjID9YrVjuYh++6lZ6p/nYk5GDaT
z793jsNLhWQSoWohoDJcRDZwZFMHyfygn8WRCNuIYHq8MY7a8cvza4mby4Inrzbj
Zr3zI2/7NYoHWKMl+gQmRklSGPKCRn1az94EyPyr2kztUhNcJ83CHmVZiDx6SVIn
N0yP5Vl3dDrIYnAuuSqHiViwSHpE1o+hX/WgdfNGSioyZCj6aQINhAXZ7xDGfNuu
zhfzndRzLhuTKqdOus7SNFvs/EkcaxSBsiO8NO8Mq9ezBXsNheCcrzaUwvqF0iuC
4D+F3aTw5RFi/cZSVClEH3+2L84X9BLLyIT2HYRaP7Q321cl2kJoSCvbJVib2r0w
2h8WuQ40RMBbJaXEXwWMirGKnilOeFT+dW7wlxKCv2defSOq1KTXUwTMdfQQZCib
6HvHW1ZZB8AFu33a+eziHfvV3vyfQXRRwb6r3ez5Bd8roXgzK36vDJfnUw5acZ2y
UCqQjeNxz1qO0utAUO77qfHNti9TyQovpltm31QJccZF6QiCdLsY+qeYQZP92MNi
+/MVY4N3BzEFplAd8YltlCXHCvzwBWqWi9jUztC/7RGjf5FV96KQElm0WuddC+u/
FyA1B6Nz7OMCcFMkNsaYmGOG/RnN+aIxJXD2HiMTaJ2WARuPm7Acnpq7G4Xq0/Wr
Iv79zoWmWCDAeZm3gxThIiD3GFOmmfOapeJUx7sJq+wqwsW6x5eaQY9v6DfiBCwJ
9dFZ8jrXWlrntQpiHuzCaEBwbP9qMVRUPkDFgqm1Ka6og5Hg0JzjPm6jIoV4CXf0
nw0PhwJgtOUjdrYKPVMd9JCQjH8ld64//gRJBJhpwKpy/TBSW36uXGgDax2G1eZa
GyQkoDSI12t8ntNft7outK/SdBoa1VrK/9PlzAyQU2jYVclX3zdY5vul/NTvwV31
hnudxtCShArH0OusGE921eG/bNFxzBL82vFkhEkDC978pU8ChYWzo2x/SE6uPtM+
AnD22P7OVnwwIQt/6f+fsoP2pUitHs9sMAtgiFU9mC9zR0BaHh24Cs6D76xLG/R+
YnvFbywnqVUQ4rMvSF2Y1Pxga6nYLGEboBOsFLdqrsPIjSM4V0hnCh6UoM52rX8W
/abDJJD/3ErRrepuTzWGeGL6Tmtpp7YXgdF0Qek885+zjJQYH6RyQsruU0+vyrpM
LGe1Plcle8J3bs0B/zqs7kKC6vdIsTWvJjwRWN0f4eqzULFbMHPbJoQdmwnUO/u2
u/VtsQuKLSl8OnwlOJy0Q71fzB92WUE2BxgNQ4RATfOgxCeqBKGUYi1+LARoOElj
wxmjGM4z9lriDILpz2yxhx/xQA7QPNSPkj3UopBq4nKDWRj9tPtT1AeEqPFgWhcX
TsV64PNI/921y5BMLfyxh4fQAG3SR7ttUR13Hg/WG9e2ouyyxQDPyif803MW1Rk7
Z7TYINpF3o0/3dMg2ea2LI+z2PXW2M/75QFSY3FBPDrSXAtoMwMNmr5QhDYdCrWl
qO9494UqGtZ3Nh8c8WOYJspLhhRcLz4+C8J7eL3atROU4b2pf7/uN6gKVCLvuSKC
dP/ANpA3RGBYCTRnAZAVef6fz8aCGP3RHcLb04uK1JZ58XrPGnhixMFcCpZe3P5U
yuxcq0u86VEw2uKeoyR1fEwwkTaBTkdI1XSy/itlqRZbE8bjuQ4KNsMCErSkaY1A
mB8hu1hTyV6EKKhvwNhNgaoiPXJwKSx4r79Xbd4aylLZzMb9BNzUJ62bTXTwYjZ/
m8qgV1AGZqxITki0WsP+bYyHgWQXBrFCrvx0mjJmuS3LYi1QjqVLsfkuqCnsw16K
8fX1wDWv/Wpk06QDbOT4KrJtLZNWVAzOGoiIsD1SlLKHb2gfMFn4+FRE5QlQmCFQ
fQ0im0CUCtpDEM2z/yDhUZkXoyCy60veS4pfeM3Wvq65sGcWVoJq6nr82oTGrD/b
5ihBXMwA0D4bjnWtlsGI/y/UfQcJewSkUdzTSsuyPNV38n4INgduJ2qKGkodE7XG
lUmdX5t1lVOxphXE0mN0Pm/BSti/rBQk+4+2XZKHySFEJh1Ott8L5IliSBBLS3AY
50OTfpGXXE603YLJXM7Z/2pR1M6qJL1ksZIIufbMdvxZkn106MmzjCxOvdBZLLgP
PlmDaPaTaL+Ex901kTW87L6rLDg412Zts07/OwDJ6pKqk3D/WLzSzwfG4X+JtcX6
7CEARO+dGEiZpcRXXovwG9w6TNVNqEmvBskt7r3BgNkpCJ1+H04PO4AJhIXg3deb
fxJQyKlINJ/R5iwxAouiM/gGdjVr7jXX6cbScV0OmRt6dUutJZQ0xGjo05uaZt5O
a+eoA0pdZS0xJVQ7rplNGXnsKGLt5QRSI3kDfq/pn/49q0DpL5gsXC+Ox6PXSi0y
xxskxGZnif00szaPCVxY5XT1DxtWErFokVNQJPVcolRsbARwAVDpbz+3AST1xc+D
R4FGAOqYnH82rJc7BMrsJ6aFJmuCASACokIRSA/dvZ7aGWHzkspU8QL/XJjxocrz
YaSrisxptBv3eyf/qhJqadzhRp5bbEodEbN0s6qDiwM0kF+PHUPHsOf4DuSjJISd
5mp0MquqntMfF9FPGmHTQCqmGilroHAa94JdMDpQPV70NHXB13eaQCagc71JdSGt
rX6OHqMZ2iv7p3YKKgn1hUU4Oc0UD42bv9VfqQ7csqvt0m/QEr+mr8QdCQPkUE+a
fsCFeSmmzcUr/tILb9oaj7tGoHqLw40TSLRi0X6KsikECwVSVjTQFAXSXicr4GOB
YHOnhR36UJ+gjBql5glFk/sXpN8ZqR3cf5/tgJz8XS0VQzlHX6XU1kAY03pV49z+
2z3Y/u0J0ZDLZoVtTvNIDlAsh6OewQN+XzuZYPluPCx2sahkqcd5sVbD/uFQ8M1H
rm9mLJV9+WhkMjfjLxrzOWJ4VrFQZhg15rr2qjMn8yapJyxdhHJIh04HWkVBdVi9
+G0XLm/fCPjWvSJsH24tRloJLe+/r7LFRrqtDEN6PQAK2qTgMD8wUof1hLkLLDu/
jAAbCouzpDz+lJqHe54Ms1f4GkpjrVFLem4h7/oZSnDFIKv/Zu+xWzZmNq0Aj3bB
hCd2iujw9k6mEg8KL7FIX6ATQ2Hc/OQWXOlnMixaXM0SnHCW3hW2BBzzNqqT3L08
OUDf8pn+BPsCxh7sWMRYvD1c4aWxgkWLIsD1viTWpESlzmnGJKFFZOQuq33eKSpE
Jorj46Z8+Nuu8jcZJic7wytVfStwJdJ0oRImWiDjlXPe707fXKGmL3m3iD3MXwWv
8YUFy6lLMMgAqkXjiKtJa2oZ/N/v/nopQyQMozxU/w2SHTuJdNsVH9giC0rFG6fb
Att+ksFhm/bev9M076Tub6MaKOoNLdhG99c3+d/6SrxHoh5nOjYEwXSRiiWyMr18
LBMhbnFTyPjLK5drvDOy6bbdFOym1vteadRkKcU52dTe4ejLjjgSnTXkmnrv/nZC
8awgmJkBr+/ZKdPBh6NiCNOOrrCgkD1SkaKx1HpmT89M/BWT8xdbLXB7bppfbV7B
MuYglTRBoipQke7INfcvxZlGDgWZ/n1svvbRew0gTBb0KcWVmafb1geR0lwiINOp
LeBuQjNTlNnp1AejG9aK5O+VXk9RezrY158WRvE734KfNHplkyhxHp762bOCK84/
JCyO3LI7uhMeZ4n4/xojySzw0nkQbNfKTUBz/xNg0yU/r0oYZIpevSlarbgTqXK4
vJJdFhvzzPG4La3+rsGCeN1kL79ad7R5dzb6b+cqs4GSr8ODIPzfyU8sE/EixMmP
SnsmLbCOoLdKjOkNL9NsRgVojA+APX64L4qkHt9TZixvTliX/x7MSHoap/4amOff
xm/EoXTq7NvQGN1YNj+ALMG+rYre1s9gfbP9dKRNcTjuN3r28Rm/yvWGzG7vEAqf
sP97hT5DCYIXOGn0AMvFwl19Qeaz9VA9CxAWxPFCrsbYNOIhL7SGFR636LFbq+YU
HJ073n53RnFtgmcLnVfn6UgLGPVFNgCckuSJUBQjEL21F2iRv9YBL5Ulv7m1Mzmc
esTOVxQmMtjxnee8OTj1tOVOmw23qT5uqxVPxZE+uyzP22Cg+mXxqs+hmCFuFtSg
I0NUxwhFVRy3x2GOonI+1EW0rAQBwhqfZJJamKjcwGpMEO8hARdRUIQghG0/i53d
JNp7OzDTXwboiGY8FIESe2aB+iDnLWlEmy2ZVceGaJ3H6cvGUn5rG8mYd8tERqyn
7/l9yCAe6A9baO2dhTOZ+zhuGsIOK56h9hkq/sTeXlacARQJMHcl/O7o3SykNBYP
0MzyNEphTONdRwjUR1wVcjul0I7dKwUyJSokWvwsYmS/WcScSCkpYPD/s4GxeuqN
rEMc5fUOyNJXHceu0FyF3ILHJk7rk/vdTwdsVuoeLtYZyyCLSnM9e9RgNK7o7J+q
N5tL1Kx9/S/fQ+KawBJRNxTpK8pw5QAo3Pt5iW+wrsSmhQLRohP7GxXbuL7wa0Ly
cJgIO33duUg0sBxitaqFTxZJY9PWrok/d+E+iyRRvu8e0YVkJAXXEDf5aSA5mGEa
+D2cwuYtnKN20e06NNputonXwC/ngrIx13QAZA/MxS+lulyOv+sBR/f45xFhYVQr
p90m3iUDmfK+mKta26WsLosI2u1kH/oQMDFoP9jnfgZp/FkfmSilEd6ZEiclzotQ
BN1KYH4xTsHi/ISUfv4lrLeQ6pG/2WrNWB9dPmKF6nf15CKuui6bH4/XUjWGkXD9
hx5q4aqpA/KAIxNP+7tQNum7G28Wp+mSwnq90sLM5ux0Wsblg921Fu3gDZG3UwlX
dzZN8147/dDCB5FGHQVTKsES2dTjhduKGhU+kTEETvG5WKK6Qd7tgPw/mwelEndo
Ft40oLyW4cDxJ6VQM9McVPkSr1ILlb8GTCNJogGCRU2zefkZriIJlaRONyAH5Egq
Z2FRZWm9qlBBqdSOJwsXvLdnch1E8gXt1KdLqRdmN+2HWT5hMaSiLq8j8TJYHTG1
VCp7FBT7YBfz55dh6avwKQO9NSYaOG5vbpRmg2LBZV0kPea2iGPUje8CtK8uvxkn
po2kJhct6xhBSC3zSSimiZea4rQwGhODsQJfQzciyg/Wat7sfSUBde0DsJe+UH5v
ygoA7UKGRtDIPK8tXidJajKPZYrMborxt9Jmid/ituTm5Oj8KaTQHZDzGdjKEBSY
OjhbUatXkeZKPwpjikqHoaB9Di01lnUyu+wd7DDOPXu80yQ/TId+Cz9oo1z7clwh
DKa0AhOE/0pMlqsd6cBhxbCEmUjzNHsFt0nvkcAwhAYlozdU4CavGYM8EfPwkpXV
Bd2oBdrqMTpjdbLiX72IOLhw1GnsuJSTSlMoXTtLs/1U9z7VlIQdF8R287lKpk9p
ZH7ATaw8jacXmue3ki3/or8gGtWXM7Ve/1kxcIitoL1iK1a/ajR9YOLmosfI63Dw
SOSvBYTVx6CZA1caVbu7wZljULUwQ+sCdGFWv4inOk3yEQSq1SlIpqXyRWJXAUXi
qu8ZO0xrHtZxnKns1LAubie/1UI7Zp9/7wpzk/Qagr2OheqbmzJAt5ZFJi0npPAM
auYvPw2EAsQirXwKWf7fKjiYg3TrZngwDxXJB5A2rnSp1ug1hRXIL94wBfvrQC+U
l11YeBkf7k0OSGkD+j2nB/9MHBjd1XxaCGDbCiis1hP+W4+jyAv9Mz9ARxRRoOiK
hxu9uHDXcUbaJgfLfp6+bvpz8yyol2Q6quliM9GClLHEMD7XosPTsHRqIPQaAKXj
sAsx4UbgPAFuIER1hE/QGQd+DcLCgJonvChFXCKaMxgdz+z0HY8CVkCFt1MPwn19
wJqhqG+wGoeCji/5/gjbP0zOGIQxZRGDdk8Wotom/9+JaWLpkDWkoWBBEM8GIHp+
teZfDNhL13ipaqgt1r9waAlcGSmuoRVE2ivv8DdMF9LJ46c6Ynt0VL4BCCDWVAsm
YKyAWwJlt/dKkPIq9s91w6iMh82tT0hRGlD74KQb+GSQjfcE15caK+FoMh4qkkHu
WJxJo+fCAJLBdVmLVM7PN07tYJBX77vCDqhyeCjQbWWlol/bI0trwNnAKAFSp+Ao
bDz7khKG3ZoDgTVqhqNqx8ZNuLWTQDLTge4gOnnsMBslNWaauhQmJJREZ7rYqUm4
aiaSTMxaucM0owwHWfrXiWpKkOCmENMcAjF8B0Q88JgObN3JF9vqJt+Klxl0A9G/
68ZztCluoC3JCdZKYvRl984/NxGnQaXQ0svnevrE7kJV6APDLS+3DnuX+fu3Ho1S
cO5WshQNXdpYLsCnnEcmtPhI6SIv0LhKyRSOtO3x9kJRrEa6Ee7cr54hBdhEciUy
c12kCPLOW1Uv125Od019jo2uAlTM5/5lBwMdY2AKmi9WyyXZcaKTMiYXMQQuveO8
+EUpDTE+VhL5etvCi94x35ZjUwOiUc3L95jys45ElFKapwQ4rLzuCmM8/2Z93dfl
aC8w6ZaU0PyaCy560Yk15/mL+ejks8Bobw72Y2zNOeyx5NHA+i0Eaqi34BD5xYtV
B+UoYnzmTCrILhpb/501Vgk3TRc4jDf7IOTjmIWW9S6eDgQpl6cttCE0hGkNIpgq
L/gQEMwQpQDJPkwHMnYBys4WXuNT8f+mB62NKo0cPepUB94vW1OOFo9GIR68R/+p
AA1AC4BfC5TQDGbxLcYp3bMPIrxV3B9ikqqU7Y4etOfCghtOT8mDPa2FaCkZNjZi
do36ZEvPFZoD7xmJqUyAA+cxEORc5ZplqVMjl7qEhTRRPvMpc6nLlzIobaYIi/g3
khz59nh6hMyl5/83v6iQ25AZIs9Yl8W+AI7AHHHvU9eMK8pDYwnbRiPidn5YjebL
wv75ON6ArkQV1HbVrGDJSal/JyVcjfkH+Frb2hqJGjpNQC2ooSF3Pcb9fs9l0C3b
HE7Qnszrdc3stZ+FYYkBb7Ypi0+CsRjQBNRnyGfqQkV2FfHrh1+8w1as2S5gWim4
J28bj361JgMjrQrRvJYWoROFxuCZm0MQ6RgdofHouWgr6HbfmuNsWqh7zvdulLuz
8VWKkvWcdryguYJV42KzLL+brbw/bl9flEZHmi9Bw2es6P9Rdr0vbCB+h0Akwn+w
YhjzY17mEJLWbqrkNXL/5Z9c8oO9BervAazrol5/F30sVubNAswgu+m3oZ1L3k8h
g4hommjicdj85gj+dIEN3DR0wP595kZs9dx7QM6HARUJ3L1lKHZZYTLXKKeZ5bav
ChgU/NwopJlpWoHRdeWz2Kd0LP5l41qPoWFlzUv2vPvSdU1M9YyruXKdXbUWPD23
+HYy3yMwL6UUML7FSH6THDas6/QY5w6jpiLLg4kpJG0e5ukRKaz0YCPEG+CWK5dp
EdJL3YreoNFyHn1PJ5FfaUNueeg41ZhWDx1BOcN0kiJwlcthJLDxwbno/Luxt0Ik
kzDPcyCVt2uW9x4/tlFDiwaw0kG+S4iTn1hGjw2/o794yqwYhds6ijTttddzS5lq
M4T812pth6neFXMNtxS4c7yzFUQibqR+MqZQmc9bbRG651g35o5vHeaMqS8BmrIR
M7ipQ9qGtm3o5+dlbIdXemqGMhKWeB1rQ6qKUjDOVMzyeCh+wVsjF+3uNQDLBT5C
DEgyiGb4ju4oALZprIVVAgr4IV6mTcx2TZJONuk9+goovW+SQhWQX4ZORRjstPJB
OlpikA6lcchVwZlBYltf/InVmA84VhPMKpSTdmH4iVDrUNzUJqRX23CCQrMq40MV
Wdj+f5X/CK3rpZvcU8khISa3DzTNJ1y2Q6W52yVADfwPLS0PB1PVRKSGD+n3zdHJ
GzVsZCXCQfahXQiAl0F4aULhQ12MyR4peD0Zclg7TMBsB2x+umrz5J1hsdtItGtX
+8SRb+vYT43EYQXl6GF9cl8o/9J295P1Ss7cdGLgisGeqDX2qBJT2UkWJQcLSIN3
UHcunooZ6LCRs++XhgiJQzNV7StQXr8jnDyvhLnjN2UzI3W6E6QbMeLdcliFNBaO
WurWmV72kj2eG7gWIvtfUTE4EYnTuNGTkgXcMqGsd9Psc5bs3rVaLJQc0zkc7hzF
a16l784ic9iabhqSLoTpquDZTLQZkXrZAmJqxvvxMF5QIfc1ES3RHydc5nVV6IEV
zDEbsQ8d8yDz22tqmE5Tnu02rCceNnS0sT0OHdG9z9BwtUszlYlUE8Gttk1I7nqg
mIpwkLcaIPehqCj9rFS6WHclWYoxJg/X89gPEkj49j8QG7CtmBebGyfWukwnzojb
2KBdtP0SbGoUe0TVnxm/9AS+uAfpDa7AImtqUvUgjxh+tG3e8FrbrQO4szYrnVJk
h88RzBLMqZRDNz1UTGYA3k9XdPo/8nQILuhP7CAVhR5SNYTLkm8cbuHksMDUocg2
V5LjzH7qG8HuOUrQlpRQBmPLLWZgAD/V0gZ72yDcVgyat8MHXZxxDkbQnPrKHeHs
H3sBUPIMKvJE9p2se36YBkb/CNv/WY7dZIqQm2jJxeXM/qEmmsK+xyTltCqZSkUA
u3WXmidT3N1WJLKMzgQpRD5BZOryYDEk35CKp34+4CWjFItg7iA4umHvhuNH3wGh
y8ARFsAw1/ejH8M6dnm4kTLxNWV0+SqHEKMLRK8sFjgEzXQlbXQN7PzS6e/87EWw
EFK8vuzrlKFI5AfXGlXY4LNZCCfvQ0J0PbkHa3wLk6t1ykwObx4IVPiLNXU537ID
BZ3/e+Ovs7aFrdwMzb5ZRckM5d0P3dFR1PL9XWr8sHJO/xx0Ty5hrOql9J8rqZ1P
GpH9aGbXwNjWXjB/gLzCjx0ZEndbaHqjskiB4Xw/JQ/vQ3R1XKsku0UrhPO1fRNb
9hZU44+jomLsFvwJCQT2NR5xWT6APmgSTE4LpzbfNz+VTfPsTEX3sOHZGXhkNA+0
wPA/lM2r0BvU5oQPdNCGWOpvzflvbM+at8etaT5emDaBQ3xzamVdQFAjrlbsduOJ
b91SI7GEljuCAuCDL9N2yxX+gckthhyzP//kjq2bReXAyRj6eRNAoU/rx55ruC6I
CNrQJBwutYJdoiNEVndJ5R6AjLiM68ejpwU/q7Gra9v4ScIGy1jh73yoPHCmFLye
dTa2mP0qM/MQU6eL/h8RZQ7j2GKdb6H4StnyY8TrBYLKlb/A2uMmuWS+lD6v3lJt
084gw5PREN+gkbjddu8NFp+gc3+DfZs7PJ6SS8NOkhXwpti8Hv4OPK1IDVbhhWuP
lP6wBTwbFr6jQLkENX1L4LiESvvRn0aOMWRoopU0/i/ivzxQk+fsX3wegomZeWRf
mZUEdOWcrrqPpiPDRVSe3V/HhqO2yYGMYpHh4tJYIujDs0GfWNlU5mwVM6VuD99Z
87HPXDhLvikMDvmCTWdfhb9TNrbIkcdxNFNxs1hx7fRvg6RLdwj27pwJcBSMmEiy
dgRz8JpsDh0yPeH+oE6fqh0pSTfYx6pMEQM8DUbIz3eqn+HkzogZ8W/t1AXtCW/q
kQL0I9U2eyc5VsFwKRjsD1PROF1dCKjjgNqLQJXeNUraebQHmzpZwEkx5VTmVW6i
sHUYYPuERdAxUM9CZY67hTeyblMghQQ4xUM/hJ0VHBZK0P3ogqRR+C8k3ieCShDs
ZA5w8nnHOZU+vlS0zqDArXQzuXwJUQNkIKECY1/0L80ooQU/s2A/cVsh67HExV4I
AmBxVt2D5rK6U897uzXWOfjXonKjIYmZ695an9F3+TxKCQP2h6aqJay7Sng7u/EJ
cWdxMAxIzsnBilvTsDrS3zbSACRRAV7s/VEXUsLKmdKQg0xY2wn9NMWDnHYPAuIG
1mfECWpqVzStwBRYkneQJIRajDV8uxGPT6jVQiGxRpirqzBuvVRKPBldEpTR1C+c
g8g2YFtnii0ZjMZmrRyQzQMn9gxtVJlc/e1RApLapHGhubkEXHmgHP9xx7z+JdJn
ZziU7nVbs6edx/s8sZq6UHVbsJkhXxOUZueyfGdkMUjW6EVJ2s0G9OYVuDkG5WcN
pBUW+K0ErydPA/FJzjMAOYFHrmq4ddTfpwXfmGRy5AKdDmFaFzWbtngddXmcE8Dz
jbuunH9pHKsY8CDrXOcVdEcZeKyqr0sxtZUazDOangWJ0S7biQ7d9RuAxIyQORpF
O2UGakB1cz2oaGaiAbjShidff1Zio6B9Y88RUwHiQJBO9JyfPl8f1Mpf/GFlvAiJ
HP1IiOL6CojTR5axj9oPRQprqr4pnXYiflcVR13SN73ybhmN8lZLTQ36xk/g/mIZ
W9zL6ACAH+YM5rMOnkLuvXwr9n1Dgh9GN3Jds1et5IyT8OxjHHCAlmPLF2Z1YMtu
rtkrZ8pJ1OJ9nPvDMu58BO9mHybltr6NbdW7B0ArDbJTqfZN4+FV3x5v3c6YWqCq
N24ZxgWcEJNUgVCagZQZMQh8Sk33UKa1nFzH7ziNLVTFzS9ifjJdtQln+lgSV1hX
hFby5XnjDpu4a35Sdqxvho8eF4vuSLeFhwegNGx2eXEjE9QKNHcOYFxdwj4ciM7F
BY3k3TUSOh0yNP8qcLAx6DS50hLCtzwGRMX9yI2h5UoXG8u6NgcM36CBcZVZEQk2
um4Wwsef+iP198i1kp9ScixqnJCOnD0u+U2uOaBvHf1anlJ/EfJCckrljXBcA2c6
3Xdlw+ZOziITceDL47uBx+CVTSgB+JBhzBuFGNXQ4aG3PhadNLcHAZKDzcMY9Mn1
BI17dm4pJfDwV5mkTttufIT8kLTrEmJfsAL8GpnbbK9kOgN2Z85xvdE/q11QX7QG
IxDjQdrtyBqR/IbaWt5mHhUYuSMtTh0jUw1OCPd9dLTYg1dCz7tlPmjgofa0si1B
ja+NM+ISpdZD5nYoJ+jcT4e2KwHLSUpFERxI0vBQqibqZmNdk9t4wXra2SVjkHKo
mWiyr2+bCUdn7t7Ba2yFBZWf32ysRV1aQTDsbGrH1b45Df5TDJUGPu+8lGzdsPL5
Y1BzXFc0Rh+21O4NHpS0OqO1itm4acO00ZsK14Y6BTG3+0m7e0gLi3jN2vqT8rsm
/a1I933aVTjKi0qL94wSpVlaH4YYlKzhf7yBbgSiaCK4NOSbvbqAhc263N4iufqe
Q3hGjMjPadWYq2jqjBek8F9oaPOs6ROVs/y//iBeO9QUiJmz5sbpyGTm+lQNuK3g
ilJzC2aUyB4+ihg9lgwKGQykLocB1j/1dTLu/nrPmN90VTJkxsYdvcrVvdzfurmS
mJoN6tBRxpUdLiG5LWzAnWcMp5l5SjbHKFAtroH86zyJyRpUEvc+Gu0DjdhzuFS6
OLsqvR5qT91sjecfbLBbI1Dxbk7cykFtXANaZm0BTm1Md71FbN/puoYtODr332bK
RVfLOUtVNieeG5IvLdcXTehmiu5MKxckkvl1/cnpCa6J2h5Wp7Nxdx4BkXHNXcHE
g0qjAZ9v+K9zkm6+SGH2uFVHmVss3S9FvPUC+a4wo2fZ+PA8f0AUg6kPHAhWNPnF
7XistuZIAKka4h9u0a8RaFjEEZQBFeeUa4JPdmO/NJcfnbPoEqvvxmCnBo6fXbDo
ac/vcVtnzHXd0xhRQn75EeDr2SffM4W1vgXx79oXqIfvndcC+Ld7yTUM46trLtHA
Lbv0B/DSY+JiFf2UnUBupIhrA3x3jLp3K3VqessAV5YFGf44hD/enLU9aZ7/+N/Q
68P1T/AU6gySckpbpUcqflhB3Jn9UJNJ+5XRLUtLGutuglFz0+0in+uiDvUdIgdE
qIVjiLBwH0m7WcXOg5a6tNCmDnJmJlW1Ui3QZi6dmCXUibzj5wj2si7Rv926elyQ
934jezj3d+cl1hVx6WdnVWOYAC5JLVu6+6nWM67Z3ybkE8lGyFQ8Ut3dAlGu+R3H
CsSE1FKdVPUDwYgxz92/mOqYX6jJSqyHi1ZAfOGqYVhUZZFU3m6OqWL/GJMrrkRD
mreSId3jKGqhiM//KZffQFSyj/kpNaD+IC7PmjE02nkuDnxvYqaEom1uGdbL6ouW
dnBzvFawyKRauypiMVOlTnvxPN3CuFqAnWTBTKWccbLP3NUU3Y17KhP4tea5FyuO
Rd0EiPkMJ/NhpB+6dBN7qB6nG54xA32mhMETA75vtk0MBGyFvP8GbAmfxXucZpPn
1Bxz40gUyhfkODqtfwG11fCft3vMkXt3fHq6UmKXuFJl8sm+bKDVKXpYdfuc44u/
ujR2RA30lFGctlzeKhjne4tqdQfgztcP2tEZwRuuoiVMWcDczEp5Ud1svLMQV9US
TU+Xj1+Wak0riBe7NH+qnc3dV3X/0sKsLl4JWsjMOHETTe8nITPIIg5/p/BgRfld
wWwb+y/MbWn1DqWGw4ANDQ1XUDbQtJltC5fjWomrMdnfaWCo3X4EuxbKRbFOyUFI
nki7UtR9gC1WZSjUB2Q6Or1bXAjKJndV86WtKlfOsH3KUPbDXao7DY87n0upNr87
50CXrN49/gBglVmsLIa7ZFHcC86dL3tRtRxrqUmLStI2GfG495bYpyqFJwqX+flN
t+eSgKAa/le+a8C4j4tgxYrSXbAeRuBD3HWnnPm9milMXWQiD6CztEVoGlrek+ZT
7ecpS/1QlY9Ukg7XgHD2VP+F7QzRUxywmIRi5W6SOEf06FBe+8kbri053fuw7Blb
PrCXIfJAxzhKEe7XjXccZQ+Si1Ifo8o0N3vdlu9D+urt7tM+DhUxEc0wN0bPrcKt
5OeURX+NECjZXCiRI71d6P/5JYcODULPQa3/niF52CBOLuCVVEkpZaLF7t81UaIT
6GWHtp//mwwR2ZQr2Spyl3ZxGg8/4LKtvFy2qNUOzkIS2LU8FbL+Mh+tWpXTrtiK
deejR9RJYxhwXquT+A2HCPquitFi/WvldPnpqXUKLPjdCAk/xbh5yHn0oDj0RbNW
xvcMGR6x4dURRMf8jbMKaOARcTtn6mPG04lIBdzJQJ+6nhyi1cqSJktBJomRvlYm
KcfYfC/o5NPGQ7kqvwetiDn+c0uFdUD3qzat2xhZJghI0LrgNRVW4Hg2Han13qHZ
0F6FUBR/b+LYxg3MBPBwJnrMjTssQkeLt/PmRUEj2tuB44yFqtlS5A0+jYQM5/XN
DyYnupfaZhwztPvwQ4ROugNv4elv3sMRUMuT1e0foaodMTrMPnXvBZ+XRiuuWfXQ
gsa4PklGNarTXTK1mdSpT6qsz4JvBTDL3L/jwI6lKOl/qk50h/DxtDHs6k1Kaz43
KjvPWSUJhGjeYlW6KJ7jSFweE5JNzdzHbk6bM4kR170dT0f0/kd8Z6tst3+4mwET
ozOoYXYSxwig+6vzITAVlrow57iYcVqK+OhwzGdW/9brT3TeEKd77UpRBf7SAG17
a5jV5D9hBt2iy6cLYMZu8GNRqOm0yD3uduMzRBV6p7H+N8xjyaQBGH8fW1e7clE+
oq2nZUOzld4E8twYCAvp+RvsgLKAF9MDZ57g8uUpPZy0tow3ehQPVBfcTNfafnsn
i0hHXY1OziJgZ8P3DzX6VZO4z70xHFHh/qN2AM16/iPxuSsLJiPYaZn8lkRzZm4b
3nq+qeMeT+IH1Xx4iUXgP1XEa6TVkLyUUiqrUd7nj89MFINJAnh/tJXuTx36eCkk
MNJC7P69z2rjfCTO8NI/cE2uaptAOz4bEUgcLRWw6QQRPevJaxFo2NSLtqWPh3XY
r2w1P1U5hdrov5AHdNi6OuoyoVSw+oTNGERz2HBH47aUiCRD0q/byidql1ap4nms
yb8Wwbs0l0Udd9f1ruh4d3JLAvivcc5OT2LiRESHAun2zQxPhyiSqZs8TRxF8nBH
YTjOY27nlCzKIGb03M2UWTTgbUE1+HwhMYWP7TVN8gX0ThcJlz8qMpa9lr88hab/
3KUXV29jzsImP757nkF00sj2vrOtfcv6RqbWHP6Suq7GH9r8zcaoQN+KfOlux/WC
yDp/kx+5jLD7xLlse0NXaP6AhOJgwI8Kr3ypvkpO4V71Rrbhc4pPYmMhGKp72R/8
pA1BbfRbk8Fsj1bu3uIKBk7ozqlA1HajkUHzQPpf8t+/r3tVxgRFZxmiO0MJvW3i
L6/n5xhYQmNMgfD0GPisw2Zw5E0Bw+2Ab1VWqE1pxcZ1hwgMwfyA9DU4+4DjhC8d
pXKCUObc9R/oSTKcmK7pI+Bgmo5QXO6ZVBme1AlptI7wmuNZzSKxeQBEpW7OvYVH
loH/RgWthuM2VNcMMJvoh1EwX2nTXyXVGAPEstzBzgtIzesKO/umg0nwfFhm912j
3gYTJxp3QBhrdSZ0yflLmZsVLsJIZLxCwLAlUXk+F7EEyLbTysPTMjAiHDoyvbCQ
zTwLZCw+lIeiC31VGdPJx0BuG69Ln15PNYpHFbtoPghRnDJj1tjx3zBiC9NriBba
lNv5gzaY79Uq/lnaNtpi5olvkoKHYLMyTeD5XNr1uqo=
//pragma protect end_data_block
//pragma protect digest_block
2aUaMgTF/PnthBS1oc/gTdVKLTM=
//pragma protect end_digest_block
//pragma protect end_protected
