`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
BZy2na6zG3CUrd8iavlAyCgutu53hwanpjX0nsMVuwm///7MAtCFP5cb9LX1GbLE
TtVeWx6iGOjoFxbuXRkCuVXVIVhZBEKp8QOxogpMLCm8wEM8ZlIu4sA3dfBsCnxC
+DoW49+iMMT/Bx7D0QT+q2sd+dSGEHgz+PZH8aB3/4c=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4816), data_block
P2v+r+LaRZEkhFQzuwDYUuALRcQ93ZPQXmu5Y78gg60Q1WFw6AUPYBFM01iTizQd
MQfku8HcuO44PHgJXn6DYNMOBfj0DOCqyHFfpt8PmZa/fcAGmW3ZFMo2VCvOeHO9
Dc+GZXv2FItOswGSEs+ZbQYuCqiqLSuL2q4+rEV9FaBsWVPZMjHhBoO8x8zuRUdT
a2d4OzSaUxAdHd36ZdZtv/fLwe5xSFzU8KQfXpfwJVoceuqFNbqSAf2rxtDEdFVf
kes1S8Tb5Txt23EFMDNkNKdK/QuSVvrfPZsyYmDRRYvZgNpSFRkWdqHA3cQ0v27n
bRRKjO2ENgFXWfCxT3iefSf2l2HrYSVVwoU5fzTHF64sWd3PP1fsPFWKh3LEWZ1B
GGc0LtEdA/2XaNQlGsul2vgORUjZ06CqJaK7okMlvVeSzU9M2LUvW+ipCdW4FViX
9KdItDxB1M3n77yqakNUxCb8WbE/p0Nt31KsBwuMqCY095sqQsXd3CyKmsDih67D
eIuMj3uoxNPUU7G0VONl+zauK40YNbGLyJEGgHnbx1M60kk9RAw0QozAQCxwhkSL
gVV1j3NzAKlhx33zgCwsL+SKQ2t25xt9BBRnDGVADYV7WBGa/3MYDfUN+x5K3Rlb
Rx1zLuRuiA7hBrN+x1FfKESeLlANgOvP5lLBt6K3NJgi0uLQfDgmvxbHksQDZxjE
hrhdpghEFE1ZDqpLiYHIGTw7oGEy3bnoIbfytyGBQ8kcjrxJtP/k2VGOrs6pOu56
bUGcXzlsW4i9TJBKMb3teBPQFpDc1s+04FaNKIewMCXy+tEnrbfvmgXRVnoiYxG5
ITL2AKACAqxcP3wI7Eb2uvrjMhvX0WLbdcylLKpHxvVKCjIFcKzJwxKSD3nglsSC
YahgZOB6V6DLBk4NWMix7+SswxYikXdQIXs4RaQBTp1371jd3xkx14FALX+HcFTj
ujZzuXrYlQkRbjIwfczEjCnKuK3esKl4uhPCPq72LZWIOn9iCxUf+CU9/wS2cH5k
1tygKnOd3LkXpUmajxQPamBQp3ULCijrHY23E7Mi3iewWOrMNaLAxSlJKJx+wUoK
lueuzJAeLKTb8OywBVPIq7YV3h9xMLwfXW1//Zfsqa5ZNSB227Wy0+Oc0VMCYkRp
Jvh1pGwAm/sexggQdBU0P6dT7lwUgjAaYaF59NLAbDYEIAax1ISUzrJ293NGRQ2G
WTmAN1Mv5Bxyplrm1W93ZnqkZbTjSllZqfzu+edXL90GT8gnP0wOUPDUH/0aBZhQ
9Cu1xDPVAInk7gVuVcbrPC2VjcbETQHxD0t4uKcnsBS0ifuHo5VP9TAR3iVfII5K
5+5NdlpgLq6BgT0AqmxeL1Cf312qh4PrIhvWLDcQ87wlNFUZpKC8g55QbGWLyTR+
Lxyf7Sjyev9uc5MDq6E8IyuTIeA4oR9VMm5pH1odvoctLL4YOXDUc3G/qLmBYmm4
LGFicJD8V7/KC05Is07ZTPTIXvtkiWC0BG/E/6Zrl4Q4RM5lwOLqD9i1NrCy8SCu
I5o0G5pryHsKf10y2bluMycS7iHHnZQUq82/sh4/Z9i+36j2UVcG4KZ6IyPe+5Xk
BBQ7L+Mv7IH2hS6zbPp0Nf8w945nwFqJeSVfv/FPMxfZeDNbkUWT26LjHCyfTOeK
GUlP6Jn+WEBdhaV+xqsHr5tn7o2zAhvZAuSGmTIjk/lHzHPMgUfE4Pg4XrF13we2
gnwFS5vfDly2oeXf7NnxJFuK8xpAV2mmy7Z5kfSEx6tbQfM4Qp2e1Wg9GWT2DADa
6XTxozMSY5UhT2yGrnDnhz5xsNEdz8+TUR/8R9p/+73EuPcdYdpXi1zZt8T2u329
1l2TNWxP7VyARTmBEu3paWnESd4+pr/4oa15mk0cB0ZjURQW8G95SBJ7sLva5NJJ
TzPo/mdmoc4iX+Xnuc59V85X3wTn5Vnx3EfBryZwZkks/aerFlQfhuz85TJZ/n6Z
QR0h4yeDnTHCxZoRo3H6EXh3E+wpvLP8S34l3nzJcvbTWXFC1fZ8wQg5jj8J2n+y
99plTMQ+GURstXj/nL088lRaz6j0YNcZP3yDrpOhj/7MVOXbk26Fe19QoJ0Iszs2
U4Pl0u6ozYlVUfbsSVLPqxtMBK3CUdq8DRoNuvH+fQVSfpvQDHxsAdeb0r7JH6nB
p2hYF3n94sfkpVJiNgdwFmHiNbbxujlOUXvEcGMx8gs64v5F9SMqK4a9Mnh2lPMt
Yk4qZ/7UuSPcJDGpYksqb1e6v6r8H9tyBv6viOahFJ3KIPOeXLCRt+beZZHl8Gw/
ictSrltfxkYjlUJuFSi4w7j6CtxqCP5IQ0a0dVzdkE+eZxFemLLMV+6p8cHiSM3t
Wu8ED2u+bohZEg0AWm/Vm3ZuFLUNuahSrj9pFy0UOi2EVZUmAB1nDt+FheEvf1U2
59uFvmg1lWNPqtORDgQBnTQZ8JeVPhPvhZWW7aiKvwyIMlW5Pp7sgcVUF+MBgltu
/o7mA4p3wH1v5/NK7OHAHwk5IMlU3n3c4oiMNJ0hOLXrQG72Qd6mRF+2OaYAyioN
1pSz7AAKzTeevJkwdUZpZ7xI8BiSCWivGnWbTE7Xt2L2LPkB0/cWCiisS59Loq2c
dlxn2FQdxii5YDt2PpNCT6xIJETAaAM1RBMDO0wTDUI844eMoSKMRuWXk5S0Omvr
xA+xNYb337ZfnhDE6zmnPgfroDtbWPJBhpD8370dPBUmZ4ZIAXitKYVYph4pirrc
047iGPM6NqWKdIabn0RAdbNeVOAWpv0nu/nRUkPkkF6Ts2yH5fFTbg+QE6oXaHgV
DxvDtVNP0+J3RMEu9691gV0BjWJ1cSKhW296cMt1jecjnpbLNL8TmvoJFcgvIpWG
lVmh7YaYJ1j6jjQQNzPzWNAGR6xIOqXwLoMDWa7emFXWQA6J6OWL1+4p91G6yUTp
8QTIAMCEUckzR0BdQgkzdJAd8uO8UauUzOFrHPFTGZSfRtQl8crh1hsQs0SquVCa
75JQV6vBSrhrouBBMPuHn/gEPtDQI7ZebKQp/4jGqNt7dX+oCVO+PFlblYIdiEJU
Di3XumLvYsgZjawk1ffE4ci5VBuwz50fxDwRSHeMSKYIwnXAr1YN4VYiF1WK6qh5
AeXBjWurcFZZHewEPvwJcVih8xRW94G8xVQDcMWHaS6iQtnOTa+BL5Ux3lk/SPWE
93X5Tgw3HegoLupgIUt0e/geJPX4bF4pCnlJXD/30j8BxQIUllGyER38TqK6kn3S
Egkn3AZEdijChvupboWofhP3gn8P5Xku3opU1hFMOlXsNPNQaG9/doA6TXeLcwH/
OYDi0/VobNq2yjwX9czy4uAFvlvWQXRNduYcWFXiA/cL0+py51CHapeWfsdAlvn3
vdtS0Jzz9VgAbe/ejdMpT3sf098Xd/TocPv/ZBEUyVwilrwiH4UbAVA2OgLf/BnE
w1JATyDTbMlffDEwE0UE49VA22YZz4Rp8Gqwe7HzwIZAxBlSJM/vz/aEonYdySYU
Re+W/sOvSbvlH4xwM+uMwMMDVkT2vMcAcHsiqDqJQXHhDO4PxgydCV9stUB4TFQ2
kT4itnAq6J9/Ctqddwg4ro6JrA04tFXVR5fiOrJI+CKCg+dRk74B7BcgKP4XwOPV
aXCpCpVyGMKT+NZPtqORRk1MT8s66tW6Zsi/w0PT7B6PdnPrAHsk0kxQhuxEXqii
y3oBpZM5oG/cVufiNtOYqjATiulb+ikeQfD4SR/lcNdFnNRriJx4700qgFoRlaCC
Yr7gvmmyrgmJAa/SSXr72ZyhssiQ6IIkxY8utDneMuPrt4I3hXBHbizD9U5Jgr1Y
en1FWYBiQWZ6Klt4Paw7+uxp3nzFXkVmwR0V7ICwhu/npoy0ShSJQF/AxsOaycco
YEkH/+tx2UpfNgVsb3qxs6AExd29GWzHtZVudAOVu6YD5HZUzu/vSYyCvS7Z1zIt
xW1BG1hVVGkECPE7EUwNcV+Fq2ktdIOJuJug8VZMZI4EvE3UKl5ZIAYSXRnmDnG7
YoTG95iA6QLyDxj/TjKZsWpd2oFICIzZeHPBC2kNFsgwyBnuPYQtHWo5jhY3y7Zn
lAJTbNyQ51xEgVhVfo61iYOLFdEhjaSYDRY22eu6MNQ6qob4OlUuAznU/ILm8PrV
QmoqvjSlr6Ed76yZOmNDG71wB/B2Yt3ufI2BZuJvGhpHd49KEQC5dYb8NtdMFSUe
CCSA7EDARcqYHMwgPq2EBYsFKXet0r3D8jSq7c0zLwCrMDsWfpb3u8kx0gTml7ru
i0X9YJng6QKBDLeukhP5X7J4pZdT8lILWB/A7/9Jyfi/qyHwuLGnOcHh7Oui7hc8
ZEB/hGeRTyqs7nUo+0M6X6K5m29ak0DnGD2nEwuS5hdJ/fjQlzgIwooTy3j3jbTt
yaDxiqUoJ4Yx1JOgOo9LxECEQ93XS4X9zvcKDPwswIoS5auDOVal8786U+FhsN7D
RLheZfmDqjZKrbRG256g8GKNNFoM1VhZMu13KdaJwtrsh/O3C1X6XzJ66NRd15x1
qZ1S5/NEPcJ5kqskCMrPNzkQC44pWm+a7lmTi8N1pBckgElH8R8n3RKHQitluXo6
JzFYpJ4i4pbNRnEpqt2ffijfddHhjm4B5l0Y4krSFophfMB3+ZNkegZX7a0rRZJH
/n4T7zXEVm1MbHrjSYeKkWjtrY0jCg51v6757DrtgSBFN4T3WKZF03TZQyolURAp
VaFqNcXMQR29QATLnCajMrRAQBFA0Dxi99kD5yLKup5mrUKK8cEcuwMxmupF7Dpw
lmltYs8MfdOOscX9SW1N2OWDht4L4EXshkbl1mUEKdgO+cswfv1mY+wzOdVE6w2l
gXHaEtsiX9JOxLeJSXlV/BYDgzaqF+RzRM2OUMl0APN1lF8QCsx8PWS1mpZ44wVB
CXU/0ImI/H8uvANEp20omGRdOPp/Cif2PNpk7YV2wzo4sM1yKFT7QgRLbwi9y9D5
QMYqdBJ5aOJKA1uCS/yXIGbDoep+KEJeJWSu1mPg71mDjRY+G6DQeORxWseopfhd
RiOeN2g9KCwn8E95z/g8fWI/WBgBIcyX9ycikw9GRBMvFN50hQMM9ux3KNKfgW2N
aEzLtyeWZFjbu2obN3elckPQFhw/nSlJilV5F/qzZ28n1QxUg45D/O9GULPti4ON
Ot+cMLdSVrN7MvatvEr6ZH8MbXLu9BLSa3CXIyoBGkyowPtAygenLbpdpfW/aL1X
3tNOMpKRwwqMnpIt53VgTS5BpRwaJzuMYRtQcYUq1pw6VEPlEfVFtNb+LN6Pzh4O
71Q4L2rfcRp5X53XhQtHkOJkNW50O0l00pKY5dM116WF69o+MunKQMGCJxmbTjQw
aPxDd7tj4irDOYNNzb+USrZChEuh1EpLjY8wKjMIj50kS9qjIpWMldIxoNdawSYB
+IfgcSMxY1EjAodNNsU9BLulFxoKiki9cnR/2JxfEozap+B8kKTQaouU32RtEcwK
WLIXutsjZxDrxh6VDvCoVmrCLDsQ5+Br/wnVx4Fy2waWASVZFcE1sfWfOuIA6dvu
W8R+yec6F5g6XDA5X/DJSjaHMXxTNx8jeBy01pXjuBWXm5lxnsmt2yjBk9usb8gu
AXyRKdtNXvePZKvFX/iEnbLWM53mt4/r4Yy4opITiWBqVzApE+/Is/f2Gw1TxyVU
jaAFZczhogvk0FKdGBAWq3OHurK4MwdAMm5O9JLhzLru+s1hDVx0OnchxVBptVqg
/dGWTwlQ0JaUReHr73HZYbC6V0bt8JfIb9xuEmLCnryQ7fGWgupwY+R2gSN0ay21
Sfyll4MPhs+dxmspVci3aPmk7Yvz8tgwHNPf4NMyhzO5zK28TlK7Hm2ychFDwBcO
Ft6L8nHa1yrt5zjowMweRmZPJ085lF2tw1qc5A7SnrMi2MK05X3mmp+3JHR0Gbr7
NZidj6Cu3+07Qu9k5SM2MdP1BG/s8TrCUS7sg8ljPUDMnISTV52OEJDlbTVc43wa
/D6hkR+Dcl5Jdz7bbZwT9B4tHv8qcil2jzNG57lr9Ab8Oej+GH9ZFBM8D9uuxPaw
m8xnJkZbBSMYr5R86fP9BlXzrXWV6EzHLaJwOG8ZygV9RlbWbR2ilGRuKhFkaITR
6VqaLVu1PYK722jkooualy9ARWF37+Vw8VzE9PIHLLebWnLjGkn/wJeudPQ8C3+f
jrYK7ymCtG4iym6CkQcm5w+sQhDvVmE3ing4k4/G8ud7AWHJhGJ00cjh5G1utIC7
7uNanVbGrUoH3avw0IldkMk6DZC64PTpAJt6O/lsTmMqGhMsYzLZxJrLj350Y8V5
huzQUCVgMPbNyFh7hNbl8Vnws/aVyL5/+scUUr0p3VemwFlnTbyaeyKTmxdfAt26
5QL4h5vvW/pX9CkQYkezAA==
`pragma protect end_protected
