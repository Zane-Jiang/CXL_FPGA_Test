// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Sxz+8RsQQd5fBMpAi44JKmz9MWEaS84S5jhDciMSa+w4+H+SGMRhRPsVtTgap1vWHiUOa04WmM/j
ByrC34X3aBRXBTmoL3BqsQUxrQm9pXyt4QYTQcYNqjQ6HOJ4X6M8p91g00dwC9aADmUrTnns1aNn
SAk8VUjsehxuAt9T79hNh/V/3Mz7c1yYshXCeQNqtoO9PpyTzcCRicV13Sdxc4BwX7pEnaLn0g9+
ukxc5OcCCtlfpOwiXMnIQWL7usYOPkzkQbp2xeAYa8WWbXuLfbf9+v43KiaZnHXv58u108f6u0GL
+g/sh4+qXqiy0cipswB4/Mv2N1H1cDNWWnNtQQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4016)
rirhdubQVNnp0GrSBOKSHlwS4CmhhMdNkBgWlbqVDrJcIPidh/W36h8cX1gxD17I3bd0yR4blipV
Yjeohn4mRI+D/bK3sX1yNvQOcinM3BVSsfbS1AA4QH9X6y7mj5uB8+E7HfMnld2WiSdUSWIkIQh8
aXscIKVdD+nc3s6LwsAJnh82A8cJ7DvJX2Vok8KObWjZj8PgBkuvr+KzoeH69w3QrTVb0Vio8uHR
wifi85tOX6TPQdcIcvRRZMb2DKpRK8nhE8VNAFaWwvfCjxiMD6F7PptUoT3FLPqTzxtNVF5dYEtI
Zo67qMu+33sqQ8Z5I5ZHLDyhBaTg/7AwyS4Y6mk2NpVoPmbE+9kN8IaZpkbJs/6Pof0443d3Zus4
UgYSO6uj4VHNF5zWvfGwBIGWHkrHKPv6QjmS9XvSgC4GjYCE8FK10vhr/DpOahSvh7ZDEnFOgpfN
p7E+lfa3Z55DNAMKf8rKraboe+C+V571Y90pmKnu/Lz187NsP21nDpFW9xfBqBoXAlu5oRyz2V3A
R94HQOPG85XR0N+6AWrX7hO6Jtq16vN1SMi6liWT/axqWW2wyIOAeQV0aqBaWgSIdcrqqcXgQFB9
vDougY+Geir3jxY4FjRoNdDFxwAqZq8688m88i83tfVyotEYiqF4W+/FFr7JcjJXvCALArEsLUgg
1t02P6cuC1ff/tmtILkhDH0l8vsgbIy8W52z7FNkelmjc6EO+xo2NwN55zcdRCIWxpk4i/YK0221
gFm1kJSKL+G5hwHyYWx3+x0pHMXQrjkxazsBKHyv4KL+AjL/O5OojhUJr6+FgYdC5vcjlWZ/MFT4
yqrxczeqqNMkf6B6sh+WKIEW2k7CI2xKLeIUJ1PX1KiJOR2Qa427ysPWqYiUzMdjwvQWjbSlq80y
BaI6Q/iT37BSaHLhMCt71+nq7tH8CLDJHmk9HfQEL+g2q4LHOkNE2rLLs2hWugS0U36D4nmtBgte
flYzhwAo9Qm+MFD91ZAjma3z40P8LxjLnhbsYKNIQDZe5SphHHEzGdQKiBDECCQJcdrGXUbyOevc
aVvtBBHqTFSntZZb/traP3JRbT4EBd4HMKo0jH5RJfOYgBAMBmSwlSocFgkwcMxhAIm8NLpDpoWJ
6eQXmr18710QxXC7aytA3/MktDPEgBm20NTOMEg/lxCOJBv/44vZyDt31rKUYnIrU/aQjH4o4UrO
4WYCmJVvj61z5/s6GH1LhbUYxDw7p6M/JmrH5Ev+kKWeHjNQ+XIOE4bt6iVOPSNcxVnCNVH7F3yz
mzVMkAJCka7DkY1oG+ex+qVmJiHRAf+TWF0eW3RRGOGF5GHwZjkxSakZyDc1Nygby1tA/J7DaUz9
qIxVmEgmuHrIumU4QaFH7YYzFu8rPbT/730pADWYg7doctXBqW2JwO9tMHMPbr7JJ315Ok9LNzhE
qABlrUgSqYPWC/JqSckuzbzg8oFmqp1GwWbJd4FzrM2rpomyQfE36gImP1n3ZonComR/O9DH4eHh
4dGOGHSZwh84Y1uuKeXDFHSW5cYkeH0bNFD5t2x7BLLr2Ym8vgfazP+fT8XxHyP6Ns5IrbRf93j/
bdDuddV46s46Elov/SVNxspmFhlh44YXOu1V7UZZJQioj/RFy1jaJk493X3cFPKRw90OKHPMAjDV
3XwKxr2N4c/yJ+FqzC6sSUf59fiKENtbDp8H5F/kizhUjMVpXGoKPx0B2i9tWx9ii/Xa/s0MotJP
1wVL9wGY0o1JF3kkw8kHwelR768o5KvSKHV5tT0j3gBxKiDdjswsXh6mMgJ1daPDH0HPctgJ91WM
anu+H7vDNq7npTSoyO51znWGcuEDCvXoZ86Wn5Ve/LMye0tpydv3uR8dKVFllyWBwbbBwQ+vTcC5
OQqmo4bhwHBB0BHeuq6sGf3fjTiu28PYkVeWDUts5Q2nn3HKA8kIRv2nemP2UTl+gFVfukP/DPsJ
1BdglzhwNlx1o+2POmCeBbOp4ciw4G42e+lYePytbiT8mSTdqi7SXqJAbllxv2HpAaZKN90smu+Y
WPu5F44R64Ru12Dpo3s+E6ZIX55AvXBsNZiVmPoqpWWBkFT+J4h2dn03D7TET3lOn9j0+fdkfzKJ
APMMfshhPLRi+A1F+xJGFMrd+zLTZdWqPVvXEAwkxaFQwzqxvncP0/N+E7BcSGxNGm7s6z1uU33y
aZRb74uWOUbEdZp1HLBf155gcpkhFBKcTEa5WJK0EFDAwwYl6WR26D21Db9rWHoNSQi9rBd+QXvK
oukpLJCiNWlv7hpK4vVaJ1YcXkP5GFqJSrV4WtF5xoqqTUSrhP6/gWtqrjyrrDStZSXOruyUqG3R
/cIa+4U0UjvObN/7F2lY7aSPBGjSk7CtJKLHWmzNXji/0npjO1BPDVfO/4jsYRc3wn4BlBBQ9heR
iJALbNr2sNDUB9EE8jXJ4heMSFpQHFnkKNgYFFXs7KtRtYtCfiKYYFqoYmNItAdA/rOd4SHlVeVC
dRb7QAInsIDiCMyWT+SOdo12GEIsVCvxsjYbc7UesdiIY6IEjDIKzfANMBscMcz0svkybCiEXprc
SIL1WC2IMawSd9NND+p9Rgym8X83v9eQD0aGZumh/0CL2VkB8QXiuxUGt/xbeZgkrwagT+Hk9hi2
5qpOVkQpB2OY1bZxugbKCAENkEhaZOiHgt1w/4PXO995T8CS43nfm/7kI09lnUIdl1m3EepKRzse
mucq7k7E+RNeQu+lGkFWaVYpaD6y36pVFzy4Zubs/McybDu30DgOlwmJ9NzI/mEr/urVx5OKOBmN
ajpY31GZrM7gi4fD7xx4p+lgpK0Lzn6nw/iaBFz6Ij+3iVcuXakgQuNmpfmhD0Bl/KRDWXp39gOx
7r95rbVOFx+7YpGRid+yieMAqA4ovkQUJOBZNghZIPYuTSdFN24sQ9210hehL9L6+ePVGPTs69sV
2mxWO+UxW3N+jFtyGWeofo6iI5OuqBauZlNc+zJfADfok77F5JYbwCeYiIcmFOvG+7/zIhy2bsK+
W7lY9Bdwgb5DdgFUN6MiULeTOnSFuLfcB1w/3py3Laz18kE7+5reeC6aPyOnzU0o0H7gn/UrrcUl
V0DP3v0zo+6VNg/tr4es1BY10akCVeq8hK+V4S9FrDQkw0OYMohFkvBBzET2CI2xsxptAGMNqKKI
2/SKWBzK6+FhFAM64x1jpQt/4v4jq82RaZSvyMK2/SjUqPm0ZKXUwuy164gyFYaEqpzqq7U46ItW
y1755vFcxqQ0cFZWvq07jx2wVuiAug4I+rq9ZqzkwTJCrN/GxYf/hUjE1Z6/XDIc2YEsBnZQemsp
TIckDAZlCp71XcxHTb2SCUQq1VDttBhTM59XmE4sGFYZ+t6ss18CLPPK8c94hwVtqFAiLbn/R1Qc
1gFbqa1v0NLapDMa/IGLoiUjWabyWZo8AcM2FEs1xVtsSZEa7eXkXa/drez7Zef2km5EaJ1czAdi
uWC7eytHz5FSE3WqSOK39FdfFqOS65BTefXOZNsXRkqRmBToWmkWu3VW1xK301etoIt8h4BLG9gx
XAQrGoU0ovdLihudNI19WDctNBDpadH9kF2UxXdRFbDck0p3EImOLmcFQETVk5MB3rrJkex4cgYH
PFwbvRa0uJeSRxcpM/Pk7142GX5nl+bLszDuHBCc1NycaUk+yjO/yrxGSXOGCuTT5N+vwe1yp4iR
KLfrdtFmWuqoZKQ1K8hX6gOG2ByFbbVSxHkeigTL0GQMv8zMfBG0KMMdk+3kkvWRbby26zpAu81W
1EBwlXGF2UsW7Mfpy1gr4FCeX25uOXKRv4tW/H+56ue8pv/CsdvBUG/JLpKgfT4RQnOZ6v0tuRjm
OCBAMIRjuUykOeu2Nwgq7bKkEpSliRH/gM6qmvwXAw0zojuRxbmnO/QQZvO6JtzAU2H9p5zBc7Vx
tJlKWrxwl4qi6q1vOQwjIqiWD3a+7HOwjRYJOd1EKY930rhTVn18AMDBKD9j4JSVs5SjC5bE3X7U
E9J0eiXFttjFBgdGfA1WOpNYswHTI9TR8e4Zd5SEj5rRH5sJNq01w8NfjvfX1P/D9bmKCVMvaNIZ
KIYJmifFe+gAYg3EQDM8mHplOlvPgfo+C9oCJqjhtmBHI8kvQ/+Dgaq9pfs9jbtzO6f19FjB35KX
R5XHwLAODobHMyPHuKyT8iE0HR8Z89903L2otJzjd1vPye338VDqoYW1vM82THLig9f0pRrGd9iQ
C9le2qBSJTqVEwx/XEvriwRH0jBW8ak4nqJARypdwXTz/Uhsi7fVrL653i+xg/R4POGDOWxACXJn
PpKLTXm+AX1eLxLvpIxts1EkJ3+xR6feoOcatsHNbnyyoH/1hHH4VFDeVXxU0B9NMfPlZBMdyhuI
Wp4i/j9P6io8roKd0Pq7yqmf6ZE3r1dRR2G9FlapESn5W69xjEtmC2C9cpl7vbc4J2+Rw0adnC30
hZtSGwDVJz/MEYS8UQrKTDZgZkbjKKgZYQ6hyXdEjbexR5RYMlEcIJaMfy3sUycWvl7XY4CS2Qri
uGBWtkYHF8tljbXKuSJo9r21UQbNjiAHa2VK4Lkamoy1pJqASLR8YhPXCKdMi9kmWI/EpAkKu7gk
oRe9S4/bXi6Q57XVjHS3++2BndstMX8T2guBKkuFNTWu+dLBfQyHBe9OpVtuYpCUSLvlVbgS8JbN
F6Krs6szBmfCEr6vitNuTP4Nt38BTFEnTYKIDyxa6BJWlb2lci9DO6PWmwXB2gVOgstorn9BilfR
tJVn6TtPkBLB1Ci9HNClYbzIY7E+k8dxoSV7GKZPLvKrdD3POHmZ+Zt8VqBeH8qI79gSbniH8Gr8
QCwQvZzBwL7mQ+jcHPWfFf0l+qQBMLxvdR660G+zuMRjKUleXP7YNgPLcBSDnA2Ckp5/dcbYE40V
plon4P7uvQVyiDF+WoofX0oykwzS25luk5qD42gRMoGLoWQPpa3JqdbccglvWPUdUCm3Ijok9gI+
VOl0X9nvEqlzqHHtTWH9HPZMQmpkwOrAyZDerLuQcLvR+nFJCL0DnRvvEdabDZWtQ+J9PyMlx2Ke
FBSVKAgTeCDppWOYdDri5DYi6q64n5amHecKeQQgL4BzauC6jv4BV90HoSx2XpOkVmOsA5BQH6jV
UaUv6L8aLw0Q33s+blc3OeRLIrzeVGHt5QBJpt66saScFmMIuIRTOs8BenQt1tdX0z5wfWHHW6B4
yM77XZyJMzB4kZ39xnbPfyctNb3Wc5RjxXk8V4oBJTkWjXS6Nst++/82riTQqFFeUvak8TXWd5u7
byKPczqmKLEPmegXnRmolzeKKWgn9plZGrw=
`pragma protect end_protected
