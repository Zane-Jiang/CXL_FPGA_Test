// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ELcpIPW87AFxcRila1EekbV3dgs6uGlGwRlPFAINCdSJI6vvV9KpECIeY+YO
DzKvuOLWZWYdtiTMZ9D3lczxRpxigOkK++p7MWy1Hx6ZqYJiHjXxp6i7ewD+
TOFcW7VcDEOVRBquqvTmAMscA5obgBEEkyr6zRC0Ih7G06FVsLD5ytMA3D10
4aNQWozC/kXdPLXpcIjI762443Dfi1ka1inVboamAHxUDJ8ZQdM+AqzzP0qk
n8d+KfOEHyafQpUbwsbfVaSOxLbonQviYBKuJwFkoOaYruWzjjX4/h4pQi2+
ybmdr+eWhKPdcNSCIGFE8l6tZQWesOI/zhf/8MsoHg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HAVyMELF7xWlLkDwwO17XMFw7Q2wisyrwnS08ulEiCMaL240BwiXq2DG8Oa8
3UVqus57YtlUxXBfpbzDAnD2fhkhvRMJvwsW6/ZLB5LCwFGbJtwOLqxPclqv
Jb24KhdLI5pG2txkMCr6YXLD1pJ8FfYj9LZMBCkeemGCvvA5tPu9qWE0fgC0
xOm6leiAUuOM7l/zS7BsqSp5nXW9A4vEu316Pyi9V5RSEbWabtFAL9dc7mLO
O8FR7s481+nWKne6q9n5UNo22jHWsN9wJUSfJmoIrrVYf4m/S38ogyxGfKKj
BXI93BRTTAGNnhknbgZabFSj8qMzVEVOpa6MHVFTDg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WWBbVWyZUccaxf1wQI08pvDjJ0n4/zGf89o0NIjmOwEPO4L+WLX5MhiadIJn
+3UrW+XEYioBVlznuXX9Oumh8iU88XRmAn3RyGOYSxmsnGDxWDu1HdmiB7+b
dO9I4tYXQmuU8HP8Agx6c0oBQIwVGvyC6/aOI6Y5ajDc3zh2DWIfUkl2c/mi
9qQs6FJWR0k24nWe5LsS5KPvqZV/gVXalZIloJJAuIZSUb56GouoCZ3YUdm3
MvSzjo/sjhhZEEN4FXtItzVZ5x+PsCtY/J9YkbnTrgBiYXSseCAfAVprLh3h
GQn5n2A5wpnjlBcNuA6RhBazNN4i7LuxRthoQM+P4A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JpRkPK6gHcKx3ZmGpq/Tj6bWcZc/C+6m4r8feK6teGbuAvzzDDYXEdUXzapT
UWobJJWvpa+hTArAVuvyPcDm6Ifd0QFTTuAJEZqt66VgfWRt37ZWGGQzRWSH
kSfoT2Mqsz+B3HkOhNjoGdQ2cM8AIguNWTDKXg84AH404Le2TAc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rZyLPB2ETSCmmIZJfEl6d5dL7KNdk1Bmjks5t5PRZqdKGpY0Wk09pPTUxYqN
wb/dYcqxV418mWfwoZvhf7JvcifHc/mxMJ0rfqyqlknTpZIDSSV+sXOQqxw8
cTJnwb97f6ZqrchBw8sLW//sbjV7Dfjwzi+UxhMoAyY99McbFLaIdBYNhyQ2
Bi2oCmbLNb8b6utYmdTvcJYPCFuZ6c0Bcr6hlnJZhnqt6KUxDtjrKHI/qP40
ePthfbGLj0/8wxbwLLCVcR5YKYYS07dSw3SIWzIF17RpBPFB/z9rx1d60hCh
1jPlJodX7rvgFoa3UqE6GP5lCrq2FDsyKRC36eyf0n7LWrkiZoSfA6XxFwjb
7KoFd9pcymb48ML9Tjvj2TDafO4Zcgq0Rm92dyirov17zwGFkbl4PocPgxzF
XhJNXAVxEgjifpDUBydgYDqLZYiGBqkIgGePMH+WYkgu0y3bltEGq2b2EzrI
FJWY8WP7H7BZKiQHyBKNKVXnchlBXsUQ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sCDHhbJiYSDP4pDrA4jxVqes0Y21JGDkRgGC1Fo2+Oz9nhT3dgjgKp/AjmTG
4xVmAYgC0Hk1ozegFJtUBFe6vAyLhYH7rNMeS6wI+I2DYqmKVc5lzeHeMxaQ
OTZKpN+IaicwG6Qz38thqJScC3DpTQShxpK7ninwERaolKe1iM0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GpOLmmOJesUFAMG3OhAyGKcSXtu2F8AUgnc2665+JdNvE/QJNYmBWya+Syep
REF+QuKvuFho6KjZxNnaDgfJgUT1T4caPZVCM2b0h1zG2G5ufOB5XOu1Ck02
Rwlx2MosrX3eCmyeO/8ofgdUGpd8E671Ys6ICBTbgFKZ6dChBzU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
pmV4ObkSZqiCacEfKJmZ7hfD80FgxWCUEDh4JxXnLNJFGo73NaNDTU+tmkZc
Z2IabQOkFYrL8JG2lCVbldyL1zCtFzPH9CTvjhnLkZdC3qqvIPXqnWfg7knm
XhJFfNmHgDa3WkA9jNTGoh4oeusVMn1rTGOVnp8BMfOxO9dEYQT32ISHdzb8
iT70fvaqb76bsoF4SATVFAoDw/wf+F1Qe9wvp081meXZc/kkw0+rKTIHtkr6
qNq8pV0BK/v41KgEqE6i7jXA/oqp8yg3qpNnZeS8/wr8smA/lOWiDd0MbmKP
4lI6N7/MPP3b+ZB+ugIX8zriSM1GXt6SR00uINJ6QZdCuvOgTWMfFQNQiCod
Qf9N+zZpscwAQ2skUpIa6+0BJe54+nqDRjx+gVYyws0FUKevC2x+lttpyffM
wLjtXEezlGhSdIac+ROTW7Q8cMIzZ5otv5yV7Whqrhutszl0HnXOrRaaz6AY
zxcueKwAyEMxJhGuxyMNBMsAscSNINqci3QkijQ8gMzmTIHUOnzJ5FTb7+Qh
1i87bVeizXQ8JKva/rXZJ75awtMykwXqbeHtMIyT0LF26A4cnfNTVfPNbQ5+
zehaVlGXIAeAD2UIbLSG+n3TT4ant5SL3QNYIOK4pprJp9/XU6J6wAjlvewp
tdGSA/QVzAJ39LcgVlzdNMv+UwRKo1cqFGvMqqyowS3zAK9f1EhDWZUM7DgS
mZ6vchqNDiMhRDcvO2ZSVoLQUx1ljlVgrfP5Bhjw3x+yUIXbPyY85pEBBv4N
m8qYWgp3f3CY31zBQ2juAjgG8M+Op/QsoIavXDKM2a7QlGFcAP4epwzF0UPS
iPTcmUlfrT5W/8qHOPFswXCFu+2I5O4k8nhqDuliv7ZkPR8BVl+RGsBBoOPL
tPutKkj2wojmHjhwe80Ct4Y+djITHmwHlHfIIX4pRBKNUo9HHXsdFdT4z5Oc
85Hvv4b2oJEfXYb7u+3suPZZOlKNYDL4PNyahynTzIFyDfR25JewZb///iKK
MtgJMhkzY/fjdbmIxDsX62LaDMkdnsZNlG4GpHZyD1FmLFfNEVZkMfSe96kZ
9Ki0syaDVoVPaiq5Vxuxt5jSpNVq0XDCsEj4I7RP9rUWBeJj8uetpFCY5fFT
yMgqs6twBw4tql6r3VOm/3wmMC8nlxlce4o6+vNtgE2sGFkk1Yez7Q61LYCF
mWKltzAOigigEarG7/vvFCZIx9/G7nPANk91BSgAe7I5bgxI/QsVp+v1MOsB
vKdlN+E/hJl2oZdyn2rbgjLQbEMSZ96ambEn+W5gGzWvuxo+p3lmrT8EDFO/
hi0UA3kB0qhrFYc/aHPpHpqBCjFk9XOXhjkqEZJklu8nUwoKJScGYDgQgT3I
gs6Rv0vFcOjF3akofyy9eR42MO/SCMs9gTw9n+Vn5WDKjTtiGYPFO7c27Izb
6LKtfCe4bEmSdGVBKq2Q39uZaOQSrRY2++pmzlZF+q8joXT+e/tqleGTY1q9
49icErchU0Wrlr2kM0Qw7wXXL+Fgr5mpoA8MqpMYflCQQUA8xF1VPsxo9VgJ
utQNmni5Nwp9qCb36dT+tSjo+iQ3DrzP1g2SHrlBzbZPQ8jyoEfUonowqRpR
sdcgma2E41LclGyLvjk1I/sv/Im2uAb5mDB1ezuVSzq08bDdjzpjTNIIpIm8
WB+jP5W7tffWy99O+PU0Qi7xFxM3Flnv3iBMPxACmLRafF6apOMOyA7B8nji
9jx97lsBPg==

`pragma protect end_protected
