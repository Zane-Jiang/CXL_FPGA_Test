// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
4dlO9C3XrQVbpCr8QevTUND/cEK7wWyYshu8X7GeJTEPlpq+iEXrti2Xq5f/d4tG
vBQLFm1deICHBhGZB4Yf0BsfTeqlw+9hvnylaoyatitSHJzqszuoVrqhYx8h7elY
B+zNaqoSrmwUnwRs7PkGWiVS3SmeGaUKs1NkfoRQg2g=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2160 )
`pragma protect data_block
6Gx0CHtOqo9n9kwUUFHF5KnlHPZT7F2kLou2WsBOuz7X/H97a84L5o34j1ge/aTc
HAN+UhGv6PxgYlTaTA4k8DhrdQIb5EvuB+gNYJ5mHEDPeKbKaFS/gu0b03c2ymAD
q304X86etMyNbUAASUPKveiEabufsykUBY3lvAQaa98MvungiTBIfqixexeWdfIG
QnO949gV99rGU9IvVQlcvGEQich4R8+xz/io2IlcL/W2BIGMeBMDj8BejzrcriuU
7p5roe/lFjJitYPxYicNmbSnHqkRu/2KyalwL+lCP5S0GtPH+GU2STQidZ6rfmxf
mdMZYADFzhW44K7XM4w953v0pjnsWYco9baYkl9783nFr9OjeolrJDXzfWrMTvqk
yp2BUnXN1bTijWTsTh99GoI+fYAZza2KmRy26uwqyWpQZ7JE03RJcDKZI1v6XL1x
kn9pOD53kwBMz4BJEMoPou2Vg4hh6XIIp9L60Je+ViDVtCG/vEiM1ueuivJ6+SnY
QHJf4LdP+gyqodDXc4oVRGU3xRW3bwMV2uKkNFwzIr+grtn5jf7M+GEAXCo6Ww6L
F/gV79B2BpCbH7duwyku+GrIYnuoXDZL6sMgiOD4aj+up5icVupIiKVQfIbpJi1T
2g3UPoPo1DMgbZlm6ZkTsSidsYEjvrv9NKelf02j0jvh5ODh3SI2NSkR7Uog5t3d
HlhOAJQRZfpAG9YntF0G+3kvSenKOdeh4zaWTeoUT7oOYHSsBmPggUKYExQO1HFR
ZWJ2kiIX+mi7dI7C02CT3NhkBRZG0LqLWXBXRskidqoEKZ20XEoNjQqVyNvq46Pv
5lNWvLA83IB28tbsA/5j4vHVl4Kyv1S1LM8AgqnkvA2RWAUk9vAz7/RZjxaKKhdp
EjqYzxo7LeGc8OGiJnhfkBX6eZIxNYxNcu8gEbv+X3SB2e0a8xEGrb4cl/rQNCL9
EDiRZMuJr98CuWpWIMNFBdcSITX6tfEVUUmzK1hEulQrZa5CPubcg1kS9RavCrl2
7B2BXMvLz6d2rAEK+NJveghYNMbqJ/PE9DJrXIOlP37nu6s/47djbQH0SNhoaSaY
QjiDFn76yOQ/nrxICuK0GzYsqBWkwJOPeLdju3GZfFA+LYoIDrhcBgK4dj+EAR2D
/y2ZOkIYaF3aClw4+ijlS5my11hhdFPi+Nlt74RTMyKg5kUUxih94qXDcUZcS6tu
moXerz2Lyr2f3R0h7KEmnnQJjyMc8E8vwfivxfLA116UXsXCf++CWJA/Vga97kUK
Ps6lIgejPKPBHwfDqrsUWk45lRy4fzSIv+/iGvyx/H+gp9xaUN4lBwgX5ael8I+Z
70OxAi//+NivXj8ZF6DOFvrYlukPi81wGvG1yoqYNwQR5uqd2xosAOZMIjbij5Jm
fbN/8krMAvGfXTp5Dt+EsKPytpEwsWamswoOy+WB3i4PUj3z+sbBkMyxwz49Xvjf
w7gyZtaYXBtCP3bvjpHCqoIzglvcAPjg2a/8BlLHxAuYarHCI/YweSdUQrQIfgLJ
zknRn8fl+TX8VuxaW08b8hPjXNMYvl0ube9AHRN2NhCYM9Ux9sse5bPlRsMnhhaI
ju7RZlgPMNxCtpehn3bPZ9qa0xRSiHI1DtDzpwPnMxLsBG5ScYBLl1zawpoDxcnT
lbf9yqk7JuF2cdRXG0XCXfqw6CT2p80J8IcT/cNlargOGKhKWfqy2Ply4LY6gvNR
lGZTncUMeJY8pDDrcE7nY9Vcl7bIBLTx6D5f5DC1MNqfaGOAEbp8Fb5z8UXsaGkk
OqKQWT9d3XZ7tRmffzCa/DrcEq1H780yv/ZtADp+FDOFAo4NuEhvMQksN1YlS2yJ
DduAJ9k1m+xrOF5CQcr7RBXx82u2jd0KKYgzyl7cAlSM6PBxNC1FmaTPwTEdb2Fu
+4/Xl5WJcGCIjM6NxL5LpKUY0PFwYqeJpCzijAvJy97X+LQ+1ZsbznzDIGOxL26c
IZWn057syHeUOhgJ5ZpvaG0Zq8akYA6QPe5V2r6D1qzBPJPImPUtYWJNmLoF8Bxa
ZNffgMtMNfTZgRAaxTaq6f2kfD21ORJ/nKfINkXakY6IwSv967Ixgv7wKWAgmwqp
dFO8PbpnAWtnMHAnm1nd1a33TKd/OCW6OszCKF9R6pxxE7mMAS06bsxc/Ipz86n1
gURKYNOQF9+owzVMX905/O1liQwTxo5965T5GY+CqLLEWAnFdIy5tpB8x2hKpl/x
ClQfzWMYp47aIOJmSJo8Chml7JlTdSX85hTXmcFLFos3WPd8OJfSCvttrH/aqYnt
4TY6f9lYFIcYd/PUvLQ+NEuuiOvT4qDoAt4YVacOvXxMw1mQH1Tx9BLDKQ/uDeer
hu70Np22k8Gt7VIu+sPG7mao55cdC1VXC9Lnidmr2YJT5UcZAqjHtvO22NwkxSPr
BVAW3ykFqxtgyKiyaP1rn5Xrh5VQ1kMSHIr9e09czMeElJUhXf4OsxEzvKnBTigI
WasTqqX/fdQgN9NfUpfVU7okEhLB5tArc/10Lchl2ANwTbfyD7qSjbnYRv4bLHTH
3hLsFJkFL+/n3QPt1EsV2k9UOca5qgoxspNhiyPCErwFIiiXKdcPk9Z45kivdfAU
RKEmmd9Ri0nwdMCHO0hOoZEvKaQVZgPSoqREZvnw0mNyEE7iVtlMdqTILqoLlHoB
5Qr0PJ2dP5TFFwm2BBq1ockkWzjTQC+95KAx6xiggFjOFDe+jMSsZsYZIG+SD48W
jl9TL0qQnFDHMlXiIqMi9U3UvaxqIIX8kokWAT6tKqMUDiIFJiylciWYrGdWhZ4p
1ENfcMX7ztsGlA46iEdYCa/PKNx0U7jaB4dxqwoTN5eQ0f5GnI9riEMJzEp9Ct+/

`pragma protect end_protected
