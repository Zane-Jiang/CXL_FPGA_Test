// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I/laY6n0PBBCdOACKfVMxGgigFMNjBtjir6ijhtvyWQtkwnJgh4ZZ0Gy5oY/
FaCZE0qiAVTXOt3OzskEfC2ak9jqf2rP6XOQhL24ChgoJ05SVHCoPLf9R5jU
Jt99tvGrZG44xmM9kLC17qUbqlM22gR7oI7WIgOmnUZlipNavEc+zKDYdGSO
XZLiUJ7o4um7VwPBFjRIgg6RFow0k2C9pPsY3NHaCXaGp5kvOIcbhifUg7vY
d9hHT8q1vdOWhn7iQ2/90khYlRO9cI7VHDI064tIiuaktANkHUBBqqpslGb0
pfmhLhfolyHfUxcbMJ8yOVDPHaXe11aa1oPdAjG3Kw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PiWAMvESZTMg1iNRswHO4OIN6zdc8yIFpFeU1y3r9QLdgcQaTac9UqK7cQng
mqt/Oj8QcznRKdacc1x57+tu2yoZLaB+vXTcrs8i09DBtXqESuMvymPQEo8F
WX2e7ceCg8T4edweLU5xqWN4DXfWWEurTAu8cifGLGsTO1vXMEVX4jY2SHqm
n8digdcxXdS7QdrYAA4d1sGEWvbfhU4Vb1SyFWUbb9y6t2COonaEHIo30DUL
PRtYyDODX3uYJ5OtvclExwb1eLTLDueIpjAUiF3VyXiJM1O1snaWNdF2rpS+
RVoJwQyWnTqkltCec5BxNdpNTPODySRnCoD2xtrOow==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n0uKNI/3gV8wBNWdV+QHp04WL8IdBN4xHErCawZV6oiMXK27c2sA9qCXfWD6
I92SpxL8iIETcLsn16SSoeAcIdOdwXyFgR7Km94I/oJ7uBEYR+MbuZmrnWaC
8YGmcpuQYk6+J8AN8vxe36U1swfBZOPS0lAp+RihlbxJNT/nxn6kbQZrwy2j
1aMvevv56JJCxXlOGjhJtYKd/FZZE8NLOLeZJpnZ8NF/sCc1WMqu7lfjdiz8
DWv3IXBc82PB/5npoexmEQn6cnn7xmTnpXFXGI5j2HLRyajDs+Tp3jpHxVpO
0N2JuLJb4lOB6UZqDLHSc7Pb5YpISAyZuXopGFTBvg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K9Db+yH/CdUUB4pVftEvtdy7X8SCJKeGc4zXf+aNJNnQ3kvyzZqrH4Udc2Fi
oZ14V+GdZyoqEKkANAwZtrIIUwLoJovZn36K1umL3QjQcBjFYMNW5pqer8to
aX/pzC/5375roF/ZBTKQOB03XUxFp0wi55oGZJ8KIeEzBe0mqgA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FNGV5hRSFf8aVhaFpTs5vq/12bPtj224NWaHyu0rCyIQwJygrnpdmLo/csaQ
T4HO2PsiLPpk2GXfgq9qKAspsO0E81xUzgEEz6RuHyf+gOorG1KYvgJEV0zY
2a4tWATYZ0KRorpHl6pCexgX8I023JM2X4pk9g4sJ5UD7bEk0+ij/dGraTKA
HjtSSxM0mS1PZa/TSlC0HfB9yERJ+UsNva81x71gzqOgrFn0zld9B+ctN4sU
JZE90cUNXbYMe+WUBmcxDzO0FV3cgV47CS6ry+dvGEqyf/B9vmfFIFCX8gHG
1xwx7RouthCnBgko0RruOLmEDZIMI1/ACeO34HQK3r0blHkRfrD/q63AzbX2
fR8xV6C96SKNqsBBJkH9zbpzxjy231YgnRX03Hs3YYu3N9x3rOyC0AbDEcNk
4ugzq6E9T1W/iRF58MNa+Mhrfmd2NIT0rKV8n1gn+MScu2diuiP69J7YaY3w
yVKat4+XUQ6PwUr4QkMWej9pUmOsRtLC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R2g8zlY0Ramy5sbZAG0lAgnoHZL7x1163kwEOg8SWEq2a1LYYNRDRjbULO3S
uaHX3v+ExuLW3lg7Uv9erEWUV6a0mXfZfu4bGvomx7XEHENUDYfZYPPwzFwW
tJDuvTA4Y15+L5aLZmvexhC4ZpTtO7GrQiBdqvIgbUsZjE4Gw74=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BQwiSnWFIt+/oPMSzsSnU5xV+mahEsrZG3xdtjgR8jWUt6Ldb2po5DtIDox0
wtoL7Ojekjw1LMgibK3uo/irpoHf1pz2ZfIFt5wOEP3HSepQ/Sc79p/MlkmE
Sl+HHoKi15MtZEPijj0hLbjKgQCvZEyy5qF2fBCZh2Yw2PdN9oE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46880)
`pragma protect data_block
c3k4VamNSphzr2DC11ndM/Sn4PX76Jaku/yloZl3UXDo5ewR63pgDGNcmpx7
eC6MF91ZEts8H03kGr9aUr6ag4HLUCHHCIPQsrd/c/ryLt4piL+xLe124FSi
m4X6juzCwe5hEQJhtjldKDsfeO8Rw7LLdmWkBRDdTSzsYT3Raggyc7zDKQfb
YBx6xEkCIYbCwzRFqQpF3skdlnmCZix+QYVergXg9qaG2ChwrSjGWPgubC6h
i3bjQKV+60nqLZ70moyl4jl/PIdrPCVcPSBfQ9Nw6McBwNTso6DQqMC5lrya
j4TrqN39IBUzocfcy0ArZTGaxLhZ9DHgo/BpQA1AjbxVJYg2E81O+un12F0h
oalIGwhWW16YViOvniBgxdGhjkSP37IX/3ASoxs65ST1susIzjVJqoRjVGuR
4J66jz/rsDB8kd/OUVfSI/kkDt2fy34Rk8ez9Z0S887ZKK15OKX0j4a/Fv3G
vSD1NzSYt1SBje+fXnaDnMHQoq1XOucWdzmJ1T9NbO8RS4Z0CaLsX+3YswhD
9y0xV+3N1poRzkSM/XoehRzPfvudmzbTLRESL8EwEH9/SKS7q8klQzgDV82n
v/jUMYm9h8c69t/pwnOmJZHaHuoxRomJrRUrpXfBWi2GhYSvWupKa8bZP9wA
iNSmkKJVXAnvQIWbHRHZr4MzhXKYgVu1eb+hrn4QR/4J9Xx/fjyk4hDqpZ+c
AyxgwDt+Cfkcs/d2chPy+2zsnayjBOg7iZQgfHbgazCNNg05S45PGovaWCwh
5y5p/zzxd9XwS9Tu1Sp3lPkDWUSrKRSuJPyIoroxhEPizXiI82R1o+xyw6ZV
qca3ySrO23T4o+1Q4n3550T8/foCeibecw1ywBWzOfCIgdcOh6Sue6CWiSAN
/LTXhOiT2xVwd5xSPrs04q648xLA6OmyySowQ4szwQx/Id5IC1RIsl9cS0FL
ltt7nedTWar+RH3n+JhJ01GCmRat2ewbcb4lxsytKgCiWKbhwb05+PMX4mzc
iAW0fSL8jQNos4sUaIXiNYiAW3Czfg7ULqToOfSAW7Z1kIlsLXGkFOGAdcih
D/qWXJ91Q2+3J+n4KRn99wjeJiXKRtuy8OlczTQtiH/pwAfK0kjqjDrl81m0
mbm31EfFZuovjmQzYDLlPVzc1qonITBWinYDZ5yTeceronOTcpJpQBrlvKfa
rqqevKaYah6rA6aACOYfU48mIRUVuBVzekWHob5zEwSzV+SlZgf1182aR20G
0uxJhlaOU9NnRiUxUKg0MNg+25TmCErwc1dRxxGsn+ttb0fM7UK50vVvqKY3
qmBNVFKotMiexdcdVpip7xWJmpC5nTjP4eUsdiikEgUaHytyIV10lRwRp4P3
fH+N8e7k409/aQi1IrsYpCNVu06IA5YBzlcAqU/ii+NzltiAPOEjk6n9NgCl
wEzjgjvyr+uBu0GjtNjaWcx1+Hll0NcWf3AaX9Qvf5PYq9+G6SOvYvfB4CnM
dwmyDnoRRuyiGNIRdHdjspZ0gH/NpBgTjVul2CtEir2Yr54yaDCATzdiUTQ0
T59bLe4IAwiG5aj36W+EbVfokp98tht/7SOZ7H0Vot2I8xBUnwBFEfjaX0HK
L5Psdp1dIBX132ZLlIyyHNLAGY9dQcGN5rIRVj3hEj5GvGrZDWVgZpRc7jBg
VWmEZOtKY0YfCuUc9JVjprcht1PT+zKiCT0PcqZCped5qjJTonCtHkZIhRT+
72ptGmI2GvXS+jas9BAvIpe/LLMvEwqyQf6L4mvbmFr2u6gRqAr2ihSkTBUG
9+n66Ew/F9rWUZwKK7Du6ic6NDEBQaVQ/HbL3c0dTmWunF0wp//hL9ET0i7w
VDai7bbR/1AzUe1tbULKu2KePijw6LxhvXsViqE/G6N2v3HNoBcEPbcXM7mO
aPjb6b+wnerMC+aDWoDFW3Call8dpOMKyh7K8RKbj5galde5KP6qSG8IES/8
B+3k0KDJVHkhVYdqz4BeOzXm/3QpxuP8TXTSJsgwUKVjMUFV8ew6AyYZcdmY
Sk80ZYogs9hx/apKI46JCQ6ks1l6ekFHnG6GYkYKUcRBDxtnpmMYTV8Y3aDc
hnjDDni4u9lOiguf5jWf7l0tf2BW4fTTUp107VSellv5vHqEK0ckFy14T3iP
uTM5urXMJz2Pm9U6Kx9MEiSf6AtdyZt2nkKQ98yjCUmqVF6lE00wlXyGKe1w
YYiFHbmSiAubGkZ8B5RPpYo7GjTLU3wk3TkmeyrwKC1d1nxfUF8sF+skAezz
eLO9/IFKZO8k+nfd6DiyXRm394KPKWN4IvCfnfecmJ+Sp2cZqAbAgtuTKen+
D12dwKj/oqAZr0Pw/eLYaAXlvsLkt3Y9QxXAJ1EPBk0qK1dEYXUlOz2exn7b
izwRouerzZWKkPJEqYAz+xLuhq8xov8M7QLGU3QPoYf+P1n9LGvy6PMoUxBK
Z/58Xc0F0hq2ytmq0G16TodtLimbbkDjRwN9iRRf/oF6xKPtZ2G/bQzKNew+
D8r/1zQpo7rxsvpIwZZ8a9b92mPEukRQtPsWFRn9qS/qrYO/R2HLlQ/zbLHz
31iU6KbnykNe65w0gG7aJXATWu/BaKtPaZYPiTurS3ntEY+DuKMlo7uj2NNg
fy6hTS/JDsN3zZeGeV3P97txY/l5GDRYC6u5Px+vtQD+vSSdtmdP74si3W3v
BJYyGopzhYKEJXep20NOuWbgDUYjX5g/KE37Y+xsoDPSUBaIWbj53US9Tw0b
WTuCmKz8HeJeGt9zspyyQCGO+mJldBdwWLn0jABJXuTl15mxJsvByDw4plNZ
LMsw5RidqoqS9EDJxVMmwd8aRFcAR5X20FLc7sMJCBbkceytWgY2HzA7mA0F
j2grfmSdjMoTuSIpESwAOL8dCFtj9xFLVJIDYSVGpTzOKFdftOaVGdaNC45P
6nXdGTkxBC2vzm681oSVyK8UE388uUqc7qIgSqmVm0wTdOAWfx+O+9cVxWgK
coVLEAIpKouTVxKYQ9vRHWjA1cUtpvzsgjRad+JRSK3biVQmlS8RgDo9H7A2
Uq2c/2ec6JJp7Vywz7TjcK9Ii/Nrdt4HaBBhvdTC24kXpWT5NzL2TrtCjytS
SI87AuMJPWJSB4yXb0FLHWPuMl84aMLCbFLF8e9rcUBMPNw6vCbKCR/IhevI
LuVOYWj0IXlSKmusHj7QQnZVYCnGqwmbug6fVwyzWw39KYwyeRJw+7mfsHAB
/C046uWL5DJLvkpoFf2RHhRwRFMS8A2PYcTyhSMSdE4kqLPElwWy1PCxcAcr
l5wjvOcGIOhZCpEWHx2lhQLFGG6oM4ecA+HQlCjeWuvRoC6JmX6WDJmappTc
dkkMTpxuKhW8jKRW0QG0jeLvd+YHzzMZXgN68L/AYs9rzFiNi2vY2OK5WRjn
UZNZdeH36nNwr/uOpwEnEyt3X4ZMQcU0Tr3LM/0FZfI09mjiwXr4pUG2RlyB
41xKeNFbdhZ9ZxuHDanP/Fyew0fBN06Ya5Hq1nXFRKhGomuZO8drCnWM7jeH
3OEUhGXh2t8dqejhYPqgWs558pFwDku912jDZwFXoDP3lMrZiDAwke5KW803
3MayEkfeM0nqzKRn8G19hVUv8Rob2xvebUThi3GChzDCwPf3dwzUqeWYuNlQ
Yjfex1Q35YVNPiluMfK6s1i4Qw9dhhhGkP54NumrfRQZvwdEg405nzuHFC6n
F4crOumF1qVsnIjM1pBoGXyz3eVZkn8TaymQaSP+xZFFf2BGqwQLUBaPizgP
fVt3zGRkgFdcAIbmqzyBHL6muk61Onbu3LgTtOix2MJJb/XA7Z2ggEemdVey
MlLijpC+lmTLa5MwEX+LYJm/I/Gyt7Q8LN2LXRtFo3C+n5pjsY1ase+GRlWz
98TyL0ePap+PELq74t9unCVr7YRxI3X7MJ9Aza1oEVkKkR0pyTwrIf9JsAzW
BCpNf9ua5P8AdN/8AsT2ZiRYPDbvFBaJAf0JsgAcJTX6w5RkFkFMuogZ3fJN
36rRXjqkVSFRdlQEFhrORUTFdEavTmUlReiQxOzRS/kY5Z5hRjkegKoKTZlq
AiBiznG+JRVrV5MBZaCSl7lcynetthr1fDtmjfSFrU7/dIBp0YG0Wox2J6LV
kpcjlBoMMDqVOWFNodlYS8VVqFnmV3WTQysSoUQYiQzaPeIcJT4ovlLNFp79
TwjoHAZ614zKeGLcGd7a9UsQd5vIlE2RR0+IWhHnp7EK3k+uX1V7tbATPerj
PjiIkEwK5AZ6hHH7RTbCdNGX4CaEVXRv+iSdPHO6dnSUNrQ/LTKD9/9T5HJT
kTXl5QFVbMIQFl4vIelyZVpAhaqpNdSvlaIW00QpG5whcMaCPxFyMdylVRsG
l62BfaeEbAyaoCchAoiLG69BMlcTIDfhsplr1NIRWsz80wF7CAFBqq7HZRHy
pFwjmztF0AUbw49rvr4RHL7Rg6cOUb9fZYaQXMpswaljqtnW7cdWsgmgKsjP
MCAM6qIOdNt0ounKJEC4pD0+pq9T5F4KjvK6HvliAMxuS3VmuxDihm22TBjF
rOJxyKsOPZcsw+iiQ4t1LShERUCPtD6SuZZwha6hN1eP0Qc381LIIrJMUnPU
aMkhNzTvs7QE7QFG/tcM/htXUH0EPsoRxH2dpu0g8BxDV1zSTCxqs0UaozSY
hsDPQ0GlugweU1o+mq9bTJKt/QqwvO/ZEmTcm36i7mpJ5obzEjnM7JlE7Et0
ntWK7Gq4vpCMLx5pRXD/Q05iUEJFYHp+eS6z1tTmarJxXCHOuzyE++YIhYMq
5CQALmITVlS5JwL2VvClzZpYZBxagip2YIL5pI2ykXBINWHulriWohjwcOlt
7F1nSYV34epBQg76F5nz2co7j7d0glwGMh+5hkNa4w7QGgdk9Et/HqSI7AP6
381gi9oxSI+W4kBzYBk0g6XrIkmCacaeHV5WOTofQ2/fiAGDQpKBfA5iKBA/
onrbU6afCeqAVG99H807Yqgow8vOAC5DUPtKzq3HluuhD9cGcVMGjwM4D9X7
yjmlDWc1XNGF83d4iPIfPE6XY5KmJAiBxILhKGnET/nH6M2GSxitRt5MQODr
sNYr/8SV8opsvLvhZ1dZIb80eRjMkcauSa1del3WZhPJSAR7rxpSLGq3Kf2g
CDzNeZRHqV9xWLMR2FdJ3/XsPEnpmxqCaRa/gOQs3DLz65ivi4xNQ4EGyGCp
+LHAF/sY2KMh0JLnoq0/pjT9dGR/CyVT4y2oXNkWGoWwtrAWar/ZtoTz0jO6
gp/HD6So3eJmyop7muc/UaiKhBSwQ7TDRuRT12p4Q4VEzh1LJmeZnvkq5S2U
I7HSbs2pyi8gq1edeAXGN4RNNor1f6G19WDlAIQ3eHxjrf56WqekzLcV7S5X
5rNrClN5J3EKxUqtQR+Isxr+TfA1SX0YnNLg4KhVU4dr7slReXmrggNAhfqg
6UXPKA1W8Xy32RVMVdC+do+cpTZdsDGbEwvHDe9KTaephzGu849467GTdMro
3thq68OoAcLq6Alc4mBMrOy3iK65FXOExYambALwhYly8Dxl0JrB4QxzBNL4
EgaPgri6AeAB9qLMDaWXqj6dKApwlfqjVyi3eEwUGX92M/x3tQWR0sjxK4kx
21qJ4l//tWrZBW+v6sQlCQYCWefhxje4GboiPTfgbtBAq23WCkq/MeXFp4H2
W2ky+xuf5oeMxunKrsq/sx9L7aruh2UENGRrrh3twmCyQt82ouoPgqzZb7PA
0ZErTsTLfICubIL4uyjv1ZUuqW2iKw6Xb8HqeR1+t1fQPqLWjF/I/8YQIq6f
Bh7mXjsvf8F05fOITWzMShuydifhWtvYd3CA3FNWXzEWJ486WQYnsczu2+D9
r7niJuJfFsuJU0GAwsN7PmABasPnKu8zt1UODo8ptLDtr/+u68yoaB9y6y4k
sj8t3aue8kMe4X517I8gPZH9VUcPX7Xar/2DN83DSZH2Qcqar+o0jL4xsq8+
tiBKnscHijGi2O1cVQOpg0f2UQ+hW6tFLTJXU2qqVt/YZTlmZim8CcYmd01y
ZodCW12CLA63g2G8D+8mbxW5ddjPrlqIEfGzDI0ix5OxIH1lK5zd6NICAEIK
nHxAmRdYLLAQyf+CBkqSHEhAfz3Fy9R+oOwOFhPX1ffcuoAe3lfNJokdotY0
X7pIdxPuQRGbjpiTpmAkZm+SBmeNtfzTr7weZaGCwBnzTty05scFWP8hJq4D
bQGK2TUr4gc518VjnU+2EuJ/Yncri30JHIP6kqMUpKXbOab1pLzL+PXu+HT9
rgnoGzbiLwaftATGBGvpzWRnxWfJmYjB94TabbSFUJ3Np/MYKzS6Easuh1QH
QhCzZRbHq78xUMlk1hILJY8R5n5i6ZkafozD43erjNmRMDmQyHeDBaDOpDsk
SseK4fWPdmTmuxw0SzVB5pIFQLVFVHEToUqut7WToG3TBH2q16GWDEN076Fw
ifQkS3wxJDiJd5OkqCGkkcxbu/gHNeeunBJtAx/LqtXGswDltPxUxp33t/ut
CcrEFeunsP8Q2mvHG6mBgnUiN4E9Dl+pGp/1nxvMxfkPGalddCSfcA9Qa/hc
uzb2F55fX55cNYRVOf6YWh0nHbcfrZvS7A9IePErWxnBbCYt7g4jvJDzdJBC
9KXAWYl9X4oq7SUf8/1jHv94z0nJpUUDwc900x7KfLNbbd6ecO1jPJUSl2j9
v2mtmourQmahJbrvcmJIRqbdEjHpjQeDuBaA0LAHW094BMjV/9JwghybbPFT
jmKoQ/nwXKSDQCYhR7qhOo0fN4+YLijLNuXn8cXqQqw8dlfMf7guiozCDYqk
bwCNfvZ5S67e4ezpHXlBC8J+hp9HzoA6sQ+BdGNzgU2yOuyo3WB62ZwLGusC
ZYU+Rn7pyR1c8G8ruEHlrxIf/wOdFQeHHmMW0jJ0bQuPMpcCT3ifZhuYFxPs
tRyw58WrVUr1wsoPb4i6zT83bkVrbNoLrUaE6COYgyz7HmNU7M6duy1zQXJg
vmdK359RJ2lQf0blmmHPN82VZtE+ehc2P/W9CePQiSMpg0kcl8JRyG5ay7GX
BzIuVHS6kLFWHR6BRSwmc8ebPpk5XhHYbCwioHqugH3DVNrtLukMuqGNDzU3
SBCNbnhokLa/bl5ULlydDbElY39h2VhFAlXwPmFzXi/lssQGCIPQ36SxI5kZ
i7lrqeNjMxndVl59ENy6IUj17OKLakeIA1RXOee108sAx4vY/TU0dFCI3KJX
PwYKyle8ofJZI1A1J1CTYXlLwbQ/8Ghm4csa5SPrm5dZ6BNu9zeFocz3aj5y
umOWRvcuZKt9XFxUsi1tSFafB3aFejbhiEo28tUiGUkDwS4GNIHEwS5rmBxX
5bn70OgoMa9RDJlV1QQZw59ZMkDQADaURI/doCQUQbfQQS2Jt5Ng0OGfLsq8
AB9Z4b9AUjj/T9BVT2GZ0eOqVxd1UwV+ZNWDm8q/WLrGcj0bp0H5SwdO34jP
MpWoK1cHeHHNul/k6iIIerdCTra9anTT4OLMgn0LrqjcNtVUOMYxfYHPZdr4
2XbhiN4V95TbbssYH2PGnTN/ENceJvDOfLUgFIReRoiG8f+zm9/NQGVD0O5K
C3JBZ9agnNuQKtiF3J8Pf0rJYVVctr8sJRrJV+ijEk2rEMgehtfVdI2N5mQ9
GOn9tTL7ki8/xGc4ovobALfC7vEhwoY0p+MdHbpyYWlMPMO/rrK6A/+d2yiU
8ncbsUGyOEbyFa4jJYEVRHICSW1RqLMrSjcNAu9RR3SGqCxjZ1FEyCuSQq8s
kMgZCuA1a34CSqDtW1DXXkZJMWB4uhQ/ykIb43sVc6pS/AtlLrLqdGZiSKH5
WMlgpSAhniQGURnC4rwZQiiN9lNqAy1+fRRvSuK/speXdC3OrAfb5lN+E+PN
uXFYJZSvht5JTiF/MwGWcft1fCqR3PaEfarMpcRMGPIM2XmLhu6yf1CDNnDD
tAygsCAdTZmHVGozwzBEMMtODXsE1hop1H8a2QuruKtitgi1JSMF38/li8oz
sDWQVbcpyDkLL72SfFw3lwUWVU2QVMQcT98bTt+6Q2g38qB8sIRk09lCKC+z
+re5IXEArMLFgOvd7sJXyGZYD2xGSSNAgiMz8SgWp+2qT4lHOJXzRxem2lat
t0QvWa0/yesWK0OvB2h8MlgrQb9POo5NhwMkEaXToOWpmL53h4LpWKdH98gf
FNUSXnc24TDjSbqNOq7r2+HW748NbPwIjgmbcLd+LyXYWJQFLFbPfOZXknDS
Z3qAyQy6FbGhQLwx6Kg0a9vOnc36vXiZ+j0z6BFGN20tmD0eCmEwDGefv9n/
ELEG0Imf+GRYkN25AIT3uuYfVmWmDYqtVVmOm0f3p7QN/+HdQN7MqbIHciBH
80tt1/QSH7OH5AnxJVVnhDtqOyZPD3KilKk9XFH4H+YO3GCm7wBYkKNMn3yG
4cX1zne8PqXAaPOs4lg/Dkr1LrQeq72JpwdL5ideIUFBJtG8xKyHAunmmqpN
bmc9tCkO6rIlGxxzsWu5cog4JEaFN21FGk5EX/8KMhJ8V4Y1WG961jqtOmJS
v/wi+o8KfoXMdp3NH9/HY3ED4WWK4DEEoPbn4aHvkYbaJIBpGkm4UFaq+Aec
klf/xttk4t2KExAuyJXOgOoAAjuz/aUv4My6R9wMj4fh66PcjOeFMgoeaaxG
wg69O+Ax7xIcfBEySnUHeqcQHec2SQM+A5kTppXp5PhC+Ayki2mfDVLdbO7o
KPXMRZnHOY+2pSKwTss1u5wdB1I4pIYe+jRXGx9XC39psWpJlY51wULkZy0p
TrQJZoOmsw+vs4xaPv3+JDm/9cXRMqMFnEo+fSkiJgAlLpS4wA3Uvx28HsVH
R4LqQTTd5/guav8LDn/84p1cNXF2QBsn2T/+JKD1We3XRALr86GXGLUZRF+c
9b5X0qmKm1cRd0lPbIPjsb1UjIcWaMvrMdFFuFqGVII7J1xOOTnctg4AeNHl
oJfpvzSyIyCtofkQZotHbd2ZyQzA9Xvq04agu3Rx8BKfvAVkPHQw/41pOvFA
dFM1r8Z+ZGjEdbIvIuBm8Kc5Ws1DNrvAJs9Y6cVxQAevdExCSadLajvCora5
G84DHnxKKHeYgCBg7piI9K0y5M7THtdJnF+9ozv2vb39RMo2CbXabQvE4JEG
syGby8y58GDa3W7ROm/+CDrWxXUTUl8MRw4V+HotJkYpf7YQmrWfkZdjZ7+9
BgQTrL7cPAiNAgnRzQKl5ESJ+dtRxLOBYyYbRtfMMlLKMn1mdgEtxoCEec1y
ENe0NdEHuCteykQ8ROzcDn13WAhsBySaarrsV3xis+YxK5onGED/7mu3zYYp
/IRmFLDMgnKZhDlIJM4W9mpnj/PObmF+ltDGy7sI/Bdbdm+XniQVdLtDVgrl
6H2ZUP7Lj+WSzH84ORSF6Fib4t1fINAYYMToX3knUAmHfyM4wNLtuc/3Cm5B
uRpJL81HESRYX4UHvKByX/5iqpoKqDOEtFGDWRSzmFpRqdyL/IN/ziRL8HKY
mcwW9Z5wBkR3SVAhA9HrbL6fK6gkhKMefxZTjn5ve1W1OW2LMbyc0h5S7Eva
ZsRd+EtS/kIyOI2WDsUSzrm64ebnMGimi1DvvJ5Ytni7NwHgKYOCPSz47lJm
5fAgJKVaMxdiMT5kMw8cRkNQVZtOmOsHmheRLNw2YLkuC0JKecuXeJw5jU1E
SbBQo8vnHUxCKSPZuf8LckbvEpY9FSTn2bFeeaIXIuzxFWsfb3i4OkWiCeki
tvmb3hpmW4O2OzPsyaUo7EUbXzuNjV4+0MdcBFePVzHx7SybEvLzV8YFnEDq
nM/wOmhfCDHx+CbWqadorsbAox4nH2X+2YdSY67NJzixlUd+XlWv+Zl3RBwM
Qt9XR1Bgg+xwgDAKBCEIPEcuLP9u67RgCdkK0DY7CCW8XKaIepBftccV18Bx
/1RdwNMO5IlQqh1yCQcctaqxmArouxqr30i037GhoX89iewSz9rjZDjI1AxE
4XAb/J+F8yhEYsMDJ6iKwtURP+3M2UaamfMjI/S4cxIK7iYyUNOmtuYZLII+
UgYOu4Wy8V8IZmv/Bbg/U5RTLxXO8pCGVDHIY8ms24YQkwTxCK1wBblrBUcg
LSZo5IxECNZmVvg6SalBol547zBxannL7y74Att9O1UiY85zVKS4eXWST9fw
OWRPefcNc1Ftdaa021ef40d2ozCa5qQuI+Uckv1ky1P0lCcupLAXOyB+JiL3
d65d9CDvK7Uhm94nT7ilXgkWBFlutE9HuByb1YuKEIz0YjYD+0rhc5hhmbhh
1LpdvRFz49ZkIx47nhOQX4I8TzbwfKuC24TL81CvmHEp/+bkwOzzubUp+YLW
1IExaz3fPC9jIeC2EOL72sazeaDDrAJRCytldjwCS6s9cDCmoqIs9IgeuKwH
W0OATJd/tQwQVCAG6VpN34b/m3IfZnnjqedySg0Vlpcfz7BvdjOaSH/m9ILJ
I0QgrjFs1qerlBEB/1vvaBteLzcun/vrL8qn7eJ4c6z7tDll8Xafp3dYz+kw
x0GF90A8Wd32skb5O1VWkqiOZogfL3f36g4KfIBfAZjwL/GwyJ35wxhSGhff
50MGJIeY37TWyZYgy4WLv6hqSXa06TEq73wGjO6g4fXlBH2QEhC27+RlsgVN
o4Wz1U0UM0g/35JXfg666rZc0yiAhIMN9nA6aadpJVED9UT7hP2GP11Vf8oW
9LaCOXcCjYk4WY8u1bMTSPTGe84wuzzlok4fvpnokLKg8F0/FXSuf9/8ynkb
IvKIyQjAm5suoqjVyy9czkD7J20V29TP9TzztPFv+sMlSHzWtHJ66wKz81Go
5Guonh9lxMd0BALO5JaiNHlWDAmO/c3KPpgmg2A52hcepwxBoIO0kyTmmNlS
wLX5T9i3RZXgeBeh/97pOighD+/g4Vr7MeQ4RRp0k9KZRziyASuW0q26iWuE
BSJxuTnYQqrGmdnySBAksVgD+sXDG+W5ta5lX+FNKgSWHEiSbWWYZtUD7R9j
CPpfRRaML/HXTG5FanwU9HZm1XZOZgXcjQztEGAZCdMvL7NE582yY653gZKb
SQu3CEWnTUu8K6E18c7Mv3eoumzek3auYDagVnpG3X+4REln7GZddzTGYjlU
xik+IvDJCLbjJRd/wnXksJ44VIF4HkV3p2WqFzzyNuHj6YRJCpKiYFhcELFG
vLEjUrpGi1FQOa1ZeU1ICegFBtHAQnYOCquypGlZNk8MjA1+V6d8h1V51tnJ
DtJtlF0vtq1ZZxVFHB1T++Z0eFJtmIq+w30TUNrQTQvATl13lnV/K46mpPUY
rg9w9EO313Z9ryGmt0zOFcu2ebBucSAD83jMUSiEUachHdUicMk6mi+rvZsm
xUOjfNjdlQ6ltvZRVVU85pnFLbsG/9U52pAlbL83E+vkZk+YYgz+AVLOWI/W
mnkc13HeEMmsAoiFoWYgp7EAQLre8IhO1UNsQbpxP6Kg0gDZRvpyCrh0PWjo
1G7fOksopzytNFVTJ+VD0ZpmhYCQQTDAkaJLvPeGMe5jYAQE3It6nRNUig3E
eu88rCOSQKuLDyGNKKpP+uis6L7bLNreSceOQvmtI7CtZvm+XsoUmrVUx760
csoQ6muZJe9M+/+xBmDscf/OFAtgAtwl92n8Vkx+w5MhULD/r5dePHLAXeNm
DVZkQJd8KTFov1KfgStk2JtNVRVCziE2oELkDpYTd2aKMMuxSBqLuy+Kp8Ck
XLh5xtD+vOxB/VqCFovWjKcoVbuQx57cXERpY8PZSpD0DwWdPA7oIR0OC/Fb
8JolOEcxnpv3mBnLYasdjjz7n1MpqhLaNd5MnVOBsJXqFC2omXGxac7y1fux
EPSxHgW0bhOIz+lsaruuSKGwDIBQlEh9Bv43wDSp7WF1REXcxIC3rN/49H9Z
je+wdqReeWRw6rtV4SpJnkJvOIkMJKeYzcPwornjTZ7k54K5FsWGZ6IRHaQH
vt+uucTIjq6Eh530O4FZEe/BVheuDEabagzDhOLtJtJYipE9pj6+jlqOjnYW
96obYm1h71MeVjLOhYDCziRqfjnvNV8HHIunGRDjOcA2CKAs/qeA3Y3V1i+O
kpvs56Q6mLNTpZjGrMDsYtrgQT4Idp3IzHG0Gz5HMkzq5rZt0k0ygdn5Oy5f
s8kMYazqRRIpMjlFWw4Grs9/DW8IMs/vhmYCeha6DUeAmnWZjMvV4eRzqbj0
2eFpWTBcj8NSTySpS87+24fVkZY/iyYRXae1BckQZWq6Esch+5ScAC3ndyw9
z4GvFFpW/q5LA3fNe3B9ftr4Mq38Hkjl0GDvhxQJG0hSrNNde62AB8NzLYUa
u0AxWmVEeLGkYWbU+B1iW7ZuoWcGcfRGbvy7wq+HsgfsCWONkufYyE1Wv6sU
yfZSPwfc/EjQbgS+xRCIlQcHGcNRel1c5MY8W37Bj7rBR+pAjSDqrBt6beE3
7VKzpS4Ctt++lurKcVIbw6uYAoE6XTSDnWHLThsEJX4sXjTad2Ua4UdCjoIg
5F8VPCuKTs/LFH93c8LuUevXTDNg1uCOCme/Arp+ih/ovU3dgrN6BDRbOq9d
dztZ4ROvmwstDGmqlH4AU3Sghlq2ZQBeYic5EJ9r6e+zoAZxl8Oo8haWYvpI
r8DIcKCpmd3cUci2ntzG+IVAHGa3HaitcNPeSGBLdINqWkGQeayer2AVeA6P
xwA149KYlKjOPGh2pckTRfqnE6yZhgbAuOlArDMisZPGPylRir+MIw1e6eeJ
37ZPLL4e0hCHlly6ztgkxJniA9wty6wVS3vfLvu6bFd1Zh1FTN7edk+oAw8E
N2IO10mF6EO3Bhu8rac9GeIDu66k+jjF+DngsZplXbU4MmZeFCYArrzcKwek
aSwwDJA5x2Yd5dyrP7fJSQc7b7zVJuyog6ftogohGW7EjlJpCnrko8xWZhpv
sLIBNJoOsrM40WlWnfcKVHgeT3qhEfPeYhrGCXw8+sMJoXpRYlGSeI79wi55
fe6dgKEWhzbBmyFj4zG0S5Qfnp7vJAIKcHnGK7Z6pagauIo5VdIODsPnM6bw
ZYmkJm0MgXsUZG6UK5SlrYbf9/WFYkk2C36xL6ATXJKMM9UGmDrBdeyqSkbw
Cw4nlcfF9xTkBX0OE4BRkljLg3lFvbXInoodMgyTZDidNvi5JYtC8xA4+qIB
ytAClostxuae1Ii3OawGvxqVZO3Bn7ty6dRH+OKKWgBPZtEchczHI0QxWdGe
nIMdaF0JzNTO0P2+iDch68EWoHEI9GxI3qwrQ7Cd73jNBu/EbNDtlzfgKxKi
YcJr4n2DH3Q+YP3I+rkXpXMpdrNh8tgoyhodgSflLrJvl6eIyzGAOAQpgjhG
R0g3dQc8qHml91aEqTDLHLre1mckZPQC/7vXTjoc+9TPXchyyfw3mAblMSPU
q9iKOYnRChRLpnMLTci2lOwkp02zu1e/DRCQqfn0Evc5tnnDd8dXXc++1i/n
ycoSKPVye1XemWTFkPfg078XFsnzfo+3WrZ94CFsfSsRwk/mrj2M9j3oztPq
8w47vnbOn3DYQ+GSpcjUZzNqGMKeo8jvldcU9O9+LtZbBwq9VjeeaKrA3p7+
6yhScRSGl2REJ3YoyHY/I1ztuxB3X1RhswSNPaZnm5qq7kT258WHUiO3a+1S
iAxzg0Y+tcCQvxDpu/8fMMpL5DxwIsWwc/zi+g5BPnj331pW5glx/iGgjYPq
EWHTECtWbU1VbL3ABe19MZnQqOzVAkE0AxhDLdxIm+UC91LJNX7rP2Y0Sdk3
e0L6+Dcbi6YSlKayBnToLMKlm3Uajnw3vsP4/O68GZlfcH9oMJArV+n35ofb
37wPgKFMXhmHY6fGN7k1N3wtvSN44rp+OnizygBYzIcmbC9dMg2+tx/5n79D
Ub7bAVjjpfvcuVQ/EBVi+e8eG3vZ21S1NlQO03jQxdM+659eMo7zKlPjrDJu
MOI9hfMCFQU9TgrkQP4jiv6Rvq8eZCwykh8k7h9N7yN791qmeU7BmRlJcO0q
bH2VR6oQPaYCeeiHJ8Mr2c4DFLClz4mh43TP8E8PhNEibJ2gRF4BXIYrsmQ/
gplFdqOxqAn8rmsUxb6WWxxnAcECX8ZDrLtJLA0AvY1hOriITY1ceQX/6SKh
cHac6OD1/+sJvMGZ6kxDj5Uv8i1zyjFOpk4qlOSxmxe5SUYtVZ4XPox8El7P
mpRKOMa55YP6VjBLgUGzYNmSAW3Dh4Yldeg1c1pyYypzVI/J1q5nM2zOLLG2
F+s6FfnoksWG3OpFAC4qdHdOw+mUdF8ChO2+7rQSZpnW2p4MAU8nm11o3wCi
ZjDBtbxnDuaMC6frDTeSTtsRvgY+vBIF571PJjlsmn4uBao/eqDZNxiuHdbx
0RJkuQADMnS4KwjpO+t8kzknsKBMGHhx6GurTd/ghLMPKdEDvjzHeHacWfLk
jXmZo9ftEPL8NSUZRo59AySuhbPeTIroYLcbuy2bZ+eybI2BnWWkwJ94KYnW
O9WXGcDEBAxXiiko0iuTAEOB0A8j83FvxpT3hRiOU+wcfIT3k16L9nz2voqE
atdRDM+ndt0dzOdrZVgc3/lQ2pN9IdwLRNefhAiodLBtkPII5u9J+BlCBnQD
JcBfltl0Dnnw1lu+DhqzIVKoiwZJMuOEC0ya/KI9yGFbQ2mFHAz5oaxMNUPl
bB0Tto9aZA0Spxp5LUfWELjmRjwpwMrSXVjjtwBfeaE1Ou1IxLgVwe0rh53s
QWy2SL8CMuuKcmmN2hCYzrbsXBk+LA8TXv9BNqDS/nMkZBMIXrsE/FmIU/dB
4fRvLd97NWMB2pOTo9SjEqwB7kvOp+N6Nfxuk+Whz9TxvREmbYSPGKiv+iKW
aqLCXaaXnVChauvGgDQV6dXbdQu35iCQWbJ0ZddAIaeKQeGxQPyJtYTEckl8
d2/eApQe8bXyCACxWK9Mbc6xsN+FT8Z8eBwGF3GYbqKRiSYbku15nP5j6ODh
UYkvO7XSj8MGSwTPno2ybfm4MpVT1DAlTPWU+ZHEsIFPNjDJRKyd+EVUxa7x
Rs5B9k3V8mX9yfpgUReXbX0Kp5sdBV67utnC0xPS0RrbAQ/YKjF6Rz/i/pAe
DnWGOqMKTSuVWp9+gj4ct+f93iiqWQhrZPKv3AYQtdHRnKlOmvKv4r03ZVjX
miHNrVmw6hauYUgNvEWNN1OHS9KH8P0EXTl91rox7d6iROh34gOR2EoC/61h
wqfCAm8plyUAprJ2zrjqmEMlYSMmvWKX7TxZs1CoZjig1riddvRpOVKvhj5J
ZiEP/WSsnHG8KxYw1jLvhLKMLOt0FmA+QNIiL/nlkggeRy2AKvowZjos1ZaP
GdOwwAKA0nxODluCJlynqcvYR2l1EN96+CUoZaJH6hLHmEzQneH0BDzkm7zh
x8GDY7PzNLH2ubEZT1RLwgSRhcbKx31TMgFk5LX+5xPwO/cdBqJAQiqptdAs
M+WAYcxurw9Lyb2tenrCSJb5Ukuq4dvUAvxh9Rs+zfcXFdbHnqtfuPLyI4oX
Q6i7STXmSMvsrOsTVMJQBVJhzhNW8PSIUeY1ajskUH7jO0JwN0cwzmqu2K8o
k4QvkSMqf6BKXVwy0O+QSqg14VgGCpqzUcfXooNgr4SZHkUq/GQhl2HK8aYu
VPMxNAXqN5ALhF+8sC8bU/VPwaZ1rW80PqAcb33sa+aw1f45uoh7So/Q/+kw
JFeJilRXTbGpJROmtEPLnhRZrFEwVBYkgAoOGxDMBEl0b3+ugGJfwg91AQ8V
UAoGAiU0wg94GfKbkhoMLOCOMQVGkB95S1iAvN0+Q/pQCPsetgHMsLaW4o+Y
RbEZNaK/CKFjqFos6MNZDQOz7QUO4IUcAxWRf9WCmDWQis91AD/RLXV+gO8n
BCB4S8v0/mDLvA09uJjHYMwvrpPnVrgNnOKje8Gvl//QO3unN6JbXCZBYjoD
OAc1WOaTv+DkuEQZENPeOkafVC6toSOPmIcwrfeLRtg/lH7fEbSA75eclHHP
LmAlsoBZHna2u5vlDbcZIDqGF5k12HR69zOF745JpMSfw/RmUYSxtNpZdinq
OVscxVyO3m+jGITD4bbqqSuoLjfl/GsPqW4S/YcfLuxSh2Sb5+G2EmqexyOI
JNMCT64Le5uyBkvcSqVDof9CyCpDpbfjjzyFEtRE1gl9Had0R/FZ1kC5pUk9
htdbxADYsY2h8XSusgPa2EO+tMdXba56QWlui1qZTS8uJJQFm+LQ9OT3IoV3
CMwtJiRZDnaXfusJuilbqHJN89v8TI6cQHXg3a1Vnqjcsi0gpKTOy18o/C67
IX6sa4PXuPuP1Lf6x2/9pcZyUEZ1GbZFKXbaWFsQNYGLKzxJejEa2PKuIfZ6
B820buO71ExMqUpjHHRdogbmHKx1NrsjUFF6uYMKTLISsxqRUEDZwUgX+zeM
yTcz6IFfmkH4C3vlu2GIrNn/6cP6HMalC7zHXHTDiJcbr5MSfdjVRZAnI/Po
QvPnjo76QeMy8JsTCE3iOu1uSzIV/VmjWRVuGNBRK2UERE4+hvLuwTU9KYOd
G0GyB7YNPe7+S7SZ+XEMmOM4EPpSEnMWAsdfY7pdSAGEg5H9PzTzAz0AR3Z6
DHPSIDn5pXsIrzFZ+DIXEoORNG464del7uK4FckURrmhWdQgQQg48e8pfh+E
YNxgeIdtlrVXI5nZGkmBE3cdSUZEBDe8VJLjkLV4XyrbPtRn1L0NLX82MHr1
jBgYBIqNm7BFVy5nH6UKSTyo6/ttyB3zYWFsu3U6SS+4VpnZP04KsPrLvANI
JrSmuLYyhHjA1GH6cxyOJRqicx2H8sSPIujKvMUdTc7FNSbzwPVEjqEpm9w5
wi+usFqRRauRaGDVec9BxMdKyaR+8ftFwI4qns0FvqaJZzeDnzB0oUmuc5di
EDwaZX2UjPAS3Y/O6iGN7UIUeaPp8T6PJhXrzEzdPT5172mt0EZ8du+ko8Jo
cQa+LSJ1kjZJexyXt7FkDEwdh+dMY6tzK6783npnDXRgQ5ZwbUzamDVg6WaT
VHWFql2Dw37VRPTmeGvzFA4qNbjvHtYWgRajOa9puCt0cLuBCE+t4Wxn6/ij
8eY1bkLTn+GfBm6m7ySMD/xep5qAzjx1nKJINICluxQafhrjt67Gt9wnwMi/
VMmGHtstsPMzhD91Vk/8tZsKTvoPDFWpNz9dl5foTKNsNBkpfvjoCxAjfWH6
v2SET3fzVk6wUp/dpOmIBQSWqzpodTFucI2u6+JyNi8lYCVXR46e1NsxRCPW
9Vx2H1adYzKmPPZz30kJNkQgUChbaqeo8nWkVKNxQa95g4k0lgXnPfiKzogT
LREvatZyhBMz/uwRymWmCsFuFs4rtF589Rs4807Ae4Rxonzpu6YKeSM2SSWW
sj1/31UonDyldnVf1JsT+NKDbU7bI/6hQO29t8+vMyLTGVacEZ/Mo4ad2x1W
vvxSl1Ya9B5/28/43hQhOkGrS7u2Q1L7JJEspj5R45pEZSm4ZIxCSsa4XZqK
R4DUrX7NnzQXqpOMiqVCbXoZB+BCwQuWxlvEXePhHMhimY0YY4NxK8iCrsIC
P8TNBwSIR55o9jcIDI29zZZGS2SBS9pmVaFtlgXq9dyT7CD9OB2WPVFZQ77b
XTCIsgrXr47Y7krAh2YcIsjyeclX+OOSW43AEG/h3bbrKDmVmDdcMRR8h/aI
zaIWYVWYVLvwR0r5h53Lr+9fVol7FQnsnNQtS8HRze3nTxaoLsP+afk/RzCc
VJ7HoONW10QGikZ6jRXJIX+u/XfwD3omagHjIIU0pRCoNv+Lzqbi7+pUwp+w
H5/WEwQwguxVD0Td26dB5vXVvG1IxV4lvkxl5qKcug8OmVdVo2T/SfDyMsYy
U6C9Yi8HFMh9wvlWrDNyZKCODnOEDCGPYLxQl/IYsVOGT8JU+DKXnGUT5I5X
9bqCo4UevjvIO2/PZduKcpUgeGbWPRiAx2Kfwpa3On6oYHY0DneCeo5MkAQK
cEY1Qi8ApMX6y4eqBdJPMRIKmYc2qdUCbShnYv/5+sZxymK3VcIZwDgqPwvm
HXRu6xJorJc+l9n+loOpQ9S58+2HB2GDUEH/zkP7cKPkAVHKEbhv3x5jnpko
3xPeefI8bR/JP+8ji/Y+hWjSHG9dxduES4FXvhtj3Qs/IJxgmmlKgl3YgO3z
0fUaKMOEWjaxtetPoMZKrtJZzaGlDd3S5Vdyct8ga0Macsf5Y/9IBNPWcG3Z
H58IAYvZpsyQ8l9oieJJr0HrgtCtypCkqPPMPOC+sq7rV1fm1WWfY6oSlcDS
wweFU1QL3/c3DSxhPI2GsDrZDJuTZ9IeNqbk04XZC5GC7h2j08fLuwEVSN1T
IyU07A6p6O6kCg6xa57h4qAn2SF/sj/FoGTnyotgEi/etC/Z/PrxlrMHgFX8
zvV4gkU8DYY0LOn6k5BWe+cnlw0zBR+F0pgeQRH9TfGdEJEe6NoFcu6ovbGE
2ccRToC5lDac3KOxUaY1n1fxpAeGlqdpatgf+CZ4KZls727WsxVJ+39f/s/3
cKz1LTQEHetAIieHhp7Hl5dJkHG5Cl4Pf6zM7I00wtLt27geAM5h0+ifzmgu
bKdeBUwPE428mWUyF92VGlXmyJtm5keC9kIRWyyy3FJW/7lMcjmna9tD+HKa
DcuVTadbUCuu0bcVpPl6OUdLhPoPATJ16jSpGDimPtfnNfCUQKmPrVru4dqR
eF6tguUDnebtseXhpApetcQSKyE6Fc0UuG7wCF4MZI5HVDw/Qg2q3WSq/zt4
11+J3KHUEnK6t2bg4MINlbpEKIvTBgb7At/8+RqA90yvWxUeYrhmEuMRs/WC
BOMd1gF7R7sZLppIrVs6IMPd3rhGQO+GAGT/N2zga2NO5An2K3qbYusTy6Uk
UVo5D/5erytvPYcR/xFtErjST2/61NR5tj/JG3I4Z6aIv0NDiaYrhaidFzYI
Q/0SZVlngyS6kaa5h1FKL6HiJvXYOpXUn8DcR28J3oOlpKfXy/DWUudDWzaJ
MRps3kT2sn6qhRLHCG+643p/u454dDbEoL7JC7QqQ0bXq5EhFdElIb0FpXax
Mu/YkS/mCdLYDF1CdSimt+SA+mO1o/MZNFAAvsDvmVteVPSBFP/OKTRbpy7C
0z1Nhb3oZturb8GfCuBhltYaO8eLumUJWZ5yz8GmB3mjESOd9b39BaNM4jhN
IBgVHKLr4H/su7I+CxCoFjM1CjVpeEmexdXJwVM0R3v9OJQHfiGTHmI06G6C
hkxX3Iz8hPAKInbcTxatlk0hs709mj2wf7OSInhIfi3W6EYvaNsY3WrJ5Vkt
wd37QV3Fs9j4/s3GNWajMfAVECLtMb6O1RuAmqQiW8gP3vYEZvmga3wJBZ7K
pQzEHL9u5uwv+jgZhh9XcepZ9iRiGV9MbUX0vDCNvXiyXPUoDgLKqXVlJRX5
v1+37BSoXo7eHjMvWWXT9zuEcuzuZOA4r7CmC4VmD+rrgTkCHXWgNyruqumv
kEHt3YL2xkEyYaD7vWQJ8Pt4KzftVBB9y3MHGMltRPyhQM7ZSrqbhDGNto53
2ON/lf906oIJU2IME35+w36AsW1MRwkNXAP1LPumQI00o4joq/qLbxoyeb2a
tgGHG9O3XhfTXiGE2K2Dlnpphfj6htlxOGt5B6+ZN75DCzg5l35XRXgQnfHN
fBJocOobMwaTwjimJFNQUyIDe/CoeV7dGwo2i0Goj8xgo1YvfIoMcP9bO+e4
+j8lkNI0PpovVJ4VAYqAWacYVKRsXx1NpO5S/Av3YVoLKTBrUgqJUzCNPQ91
fEcqFj+gPBnK0gei/NW8sEeXBPJYd2FVPOOjpxM0AbT1+TWxGwtOp9i6h4r1
BVCp4fJIFK1LabLVjRCf006yZLv7GbkhBt2/8tuGxSyb3DnOyIpPn/wSq25Z
Bvl7YYHl0YHviH5J/wVQiNYQLZHPep1vwtJXmpJoVx3l1JwpcUfuNXb4+phM
kidyoCVKOVuYD9lvWuvmWXUk/OA0nKzMXx+PFNaZLnkaxc6dZWW8W6x1LhYr
yrvmvMxX+MSF9E2OcDuj3k9fueiL52Snf4YLtmTY+2bW+o97QmgSLStOnjhS
lFnNSCCq/MZTGYyJdnKAv6GE8ggYp7ZV6vzhp8jrvR/ShxVpaE6mMvhuqWqC
VWMoY6qofWCmqctLb3vQPGZne0RsOhZe5ulwG0ioxaa8qaQSt0nhU51R66F2
tRUbgZ4PaWfnd+kGqSu1slSY2LPTLHUVTos74S6C8hxoVCnCyyuO/IbWzjeN
9yXgJRISKq256hv8iYi9RJsrkolKXcmFubXfL6WBrDkIKC5t+HJGeVZfxakq
SQxLX/iTV7Pc0cq2uperQLPRnRlOqTdwZLmG4JWMtR/FBB4eqm1AUDBGajZ1
ljKsD/v6x55+7QmA4ht/jSx6LkpjI1AhubKu3vIBbuxu9tpwuAJC4MlahYNq
uxXYakfUpSqrxc8gczkw/APbQNv65ww704Q3Oq3UeJpMUQHXh+yjssu8jiZv
lgtO3zEKDviw0olWnOznjGyaiuQythaKBqyva1FVYbR+ppxcTB8ahODM5ddV
o3G74lsV4p2232m1ETK2R/x5AaangXbCgigS8dhpLmUHP5CaGXcW1Aehg47U
7Xh2A0sBY8eMSriShRbzXxMA8EcZ3xGxuQr/qD5WxH0+I8mbJpNYNxE2HYE7
g++0Eo1eqksP+S9Vo5A1wTtznf2h7DLh2Pck43Jde7LsoeRgdIDOwzzVdr/1
XhSkky9Hv6pth1o3sJ1mCXJQfgHzPv8JaO8avHuEzlyIq+D7iXaabxswqBvh
CznMjbqdmOy8SEe+//S2Om0/rYxUZt3nrE9Y2cesrxVe3vLbQVr6ilPlHO61
8hAuB6cMLmaKMwTnZxO49i9j/sPNVXdR5Vai4nx8FRqY9PrIa47/WeMyENsU
nnBBncrgDLmFzqLGCdC8VphQQ183mc6P8/cwHZCxjAsl7LcFSWudhgOHhic9
VaNm8yfzHfgKlcEW06wXrbdghCTnYxUcuIhbLjcSmxGNWFY3iaY+Gw4VZ8af
a6ctFJ51JEQhigGbL/h70CLveA0+c0j8OuOE8gojS5UxatbbAgrAxr7MmwCH
O/T7e6NsM/PPYu/xGwGcoiNgTzB7077JRDS5PmGecSQMVxXHUi4bqvKwokuN
F224gKNlenpM1wONYn5Wcn2aF7sKv8n7b/mt7zDrLsMrACDaPsyFdSfVlcQ3
C+KWmguZxz53mvy5pCpSwF6ONls4dAK8jqrNNGEvGx4pdYNG+uvXdvEy2mWe
HHsUh6AcJwS06IrzEp8vQixYv0CBKkMQEjCNmp7gXIBLpvBgJEbhMR2z/Ffv
ivtJfOD90RidrrOCbgA25gmw4ThhPJGUtLSIRKZQGH5BCHNdOMR4L4Hlm64O
cUk+rIAnifHDJGPirgy9TB1DmhN3z/l2FT99eAtpxgGt63KXlbLRYbmFQjkp
2V9/LGasRa+9db+4oicNrXmiklK7f15V2QH2Ymmo9o8rFDaog4z2af0r342g
/XC4lcsv5gtFTdOX83JCXdynlJRx+/mjYxFJtaFshrlwtOtYG6rbO4MZqR9X
hDec+dbJZcIe5s93XWQYSowJKsAsSyKpXDlVjOGLQl+7QdSGyc9tvVr2ZhpZ
WbaTWNWfezbpU6lmhnpqtJAbZBuSSq51ERLbEi3Msf0fmwul4TA5U+D8Fv1/
ULEZrSyrxmISjhE1hosSEDY5Ov5R4G2keutIGWwLeL/VLjeHHL2oyeVcEngC
4nLT6h+YPhgcq3aqNDBZnuPLqOwiDjFBiKZocYfu+02RAIyg4Bz8nCYgaVze
bF/F5wq5cTHTEdTtm04pAXMde1UMj78q88sgAW3MkZGuQqzRmPMEo6SbDunn
hfVzALDEgrR/bNOA3+aDvKIq/jOVLQBZaZlgTcVZPOcgI6G4A4nZU1pV9wrF
BQKZrMzddMyz1Jrre9XNzsRcRIHlDlBixcHfLHEGAH8Mh9kxDYwfdiC+XOe+
00w/T4z5+3fRY18IvFK83ks5qESTifSHCdxAEQ8uPuNRd0NbTURleAKqqzXu
pHvIdCgNaIcKzpma+F7K2LsTj/BhR6C3jzylRUHW1u2fUAYRYLeTuG43s7Uo
PkZcN1fQcAb6QamnKhbTtSZfLYh9FF8h+8YaY8t/CySapi8tzvTt7z369i6T
BSZt1pz1GrnHDtalIRNOmEU8zVGkD2/GmvWTi6ItuT4oJFq5NfjyWf2PB+cP
4glKm5qWpaDynasbnnLzXknNvJ+c6KrO9tazFBBNRW4vkaxfTvSVMa3qR35n
X76HKwvYyfk5PeLqAUoF+zjm1ViE4V4wJTuilTEOP2dtk0XbBSNZ1CPVm+rU
/ow8k0bkxKgDcurLTr0/VgpI5vEhGUxBl+1mwaIo9Jm90ti6MJxD2V4Y/Qmy
W7rb8qDt+P18QAvZON9dh5vMFpVuTca7ULGthUZNJCaCEd7+CUEIfl2V+Wey
8R2W00s8f7fpUvw3ZGUCiFkFgagmgRKCIo7Sy7hYF3hpgf4Ka7nxD018U80F
tSXRJrrCPMF1U2TEaHqeHyrXgvpq7pH+BbpfrE0hzhP4ob6Hg9N5lQVs4j74
3oUlydYaeowb+a5SEEJNTmot+7il8GQ8vrs/HWl3DNeSEkF6Ax73Ww3vkmU2
ncr5115Hz6YtgjtLszxk3Nvufthh2qHc3thBvG4cugCG9jVpC3RtT709Y1Fg
PNbLgZb7lh5SSJnThx7h4iI4LEMajsS2GCWazUlr3WPuT+qh+A8rGyfrGSB7
iMv+iWWTTql/qnP2vX1GEMF1BvypEentTk8Zst/72YxKRKtbbMCFFdhdXZ0m
qp8E89i4FgzKREKlYzQlekwPhFB84xd6y1bL+y8QKw0ebX8hLO71Hgs4vzfe
C6uNGhmIGJIWSUYEsIXGNbTHIfQiZtsXeGLgAbpvVp5Bvy4PQHBo8qeZV+Wc
e/WbyQ1mlLx5pmBuhItpWSlfjrBZ2b0tCTrGNJftadoNae+TW+N48VhWyT0F
KjojjkT+lFGQ7PFdKQCHRW/uoYNnmVARpMg+L4Y8sbGS3zAIYm0nDL6nZW/d
ZoB/SN7skndk/Gt9kE8Uo99wSzEldMC9BVnUXUnvSsFABsfKmNuxF2FO3vRa
wIE8rCwwSFipE7ZF8J/B2tKXjX5wn9NsljlwIJ6u8e2de9e9RxIQBNOe9/vf
Ft0L/jyEVimccwKvJtH+ev/bhuI6ZtPfxBpQIAte3o4//BLb1QFEoxUk+hnj
JT0JgUQKtQFEkIUtML0nohVuo/WdZSIf+BcfnR3DBQKR4XigFlnE4vRG10gq
KbuYlRY49UTCILSeQEhYtkJSiytf8pkCmAz+Z/DnD2w3etR+NOXFoUKf/Nbn
jhv3PK0Jk14b1CXCcn6KP5YrF6JSouZBYh5kQJD4Vs0Ev/ZMJl0NZ3ZmbdqI
v1pH9Lrkl+vfadiubkHovFequvliaaMZhg39CaMZ8oYOWQDnt84KqkAPPEqA
Yb5BnxsgbVWCpHiYQ2rqwKCN5JL88oD8y3SbkTPzb1c9lIDURiygnVavGVHI
Rj4DpgCQsOsUR03wvna1iqghUYLPnTU6GM+6cKJEO6I2rg6enR4rJZhm+uJU
bT+jFCFSOIt8ZzkmkOERBGG8jApL0J8haaK82E/9IpqFPh3KPnSrezIR1ed0
A057IM1VC7p28Gc8Balt3eqUPVS0XuvSAjDdbC+NgkludFX9Xv9TRhO2mMXh
wF5CLAJsRGF95AXrXsb0xSkw5mBP8nIsMCWYO6mVPPXphHvQpefyP2ELlTFD
N3MrB0J9yKNQK/Y1kMyMP52HbQScnisDArSt4RwF3UvKmmtdkLFmLvL1/nWV
n9q8qzMTbfz+OTIcWqxl9wfjZMASyABDMJQ3srufUJFsT7kwpbFcs2SeESad
9znJJvV5FaSMUonn0I5qIjXj+jcL7KmukvIm6SINVv3DK15/j93haISORpp7
LuXj9b7pvOgXpSqOJvVSI9P3gE47xMDk1a2B2asp5IO3/kjtu9mFz8ibK4Pz
HK/uNKEN02TUGGDX+pOZ2MwiuwSZVhAhQ0NsBIjIL9Fo+T0We0xDvdUEFla9
piIoDsfwX4xBOL5Z9YWpVYZA6oB+QYHdMvVGwrmD6+fdfpdMP/wsE/xMzpfc
41Njxw06wyUhvH3yaW/Eu1y0n4AIijMKaoYDSrsVgxaV+L9/XRSIMU2DY+Om
kZkyiFAVwUU8KSS4+avZMkUnLV2KXJ57ZfAp5MjsXlwqHBOL4UhR7aoQnJID
ZAmPsXSzrehkEfILqhN80UpG9rJo1sbhtgBXGcpKCMpb4NEB0I4QWreo8D9Z
TRMV7bPft5LIXmL8s2LH4NQw/kySbtMKhdbBw49gNE2g+qbZ+7taCMiuwl/3
0FpJpUYtKfho5uvc9fYrBV+P3hIYVpyAmfchKuDudL4R2tCCRE+6/UliINYa
Xzummw+9148xmEsiUKeuxMLnJ6T603t5LIPU1Qv8Y5RYuFJkuE/rYip9/Rdr
a7FqPSVkSnVYvhpK6RV2ozKGCODDq70rxA5TC3N0X8yqkEbIRm487Oi5kVK5
Epof8SXkM6iXBfh3SZntfuluUtOETANFe+Spvs4vH6LCazxeWVZ4oZXbEENF
LJ1mtftIaoipmMVkYF2HOItJm69cI92mlQECU6bAvy1o9GaAfJYyg/q/cvLG
zuSP+QZti8t3cSqoPClMpdvz1Ey4dFKQAib3R+/kJkf174y32paP/Mir5uzP
9ZmoO4Tr+tpvd3jrL+ebReZOsdFCgbZjt2WOwqZR5DnsqGsHgu+SnP4ZWeZI
pKCh3YxOh+4f1unTUNle9JSrGacjHhe9Tgb4ckviMKFklDI9GnrerjR5OPZs
cSoM3OXS0G70VkCYTlWqEXUtGb7RD7Cpa8sC2jl+Q6EePFtMhvaUSTGHsAAF
B8gZqXQgQeRgZM8gIKPvqqvJbuvlFK8Jh1/I/Na4UAYmZAEGd21/9J7KrHy/
PuMCpQiYTz8qS62neQsE1wgOM+uQmGsridROiCFc9o4YkOVwc+EMew86+z5t
21eVy5/9cmxkL9vukT7lf8N5TfsG1dxqSK5cgNCdQ7ZH2lGDHQvBzwGGnqC7
PaEdzUbGRL02fxhBmXa5Vx0xNqz8IuXPnxikQcod4teKNyoZzcrih+NgGk9J
vmtry7R2kb3DrJIO6tUcjk0sxpFWJ4mxLZ7o7zKi6byv7P+0Krc9evol069H
Zc5jgDtQ+B0nHKaOez47lhFzlu42V0KjhjzY3Fna0hmV1bDUZeaaeS1gMPoG
C0ZY+XT82qgMHDKNOMYI5uJjaEW54LLeAjT4VGVHX6H/v3vfh+Nh/o9Z/glV
0ggQYySLtVW3RMNMf5L4ntWndNZ35HzhmjwJIWNU6DEQx5ow5kHbMH9jyijx
d9soNe5oCE3QQ7C9ahFfMywNeSKtX6bwpMR9kJ7T9lYY1Mm1eIdBo7AsvzKq
VQb0m2HghMn+BojQhFGCFONG9BAzwdDZiY6qF8gT9teKjaD4vHDJayaArfdb
pm01+GF+G6/cF+a2KgKkIhdEOfZ9xnZb4m4I1uxtbSTaRbM5dylrXYNbXqEm
VOY+urD2nXnWtPwUVGsepnjX2d6ag96t5BTlw7XQ1gjDezVO+LGWaM2EJZ71
zZRHrjCzQh3PEery9JNk9vCIm7cmHEHLRNtFnGi7pco1bjWW282kQrNMUEt6
Xk4a2xItYhsnWlBEJv/mlDsYH2dPeVq2n2N0MtWu8lUtSpYRPMyJU+7apdLN
o7D0cz9R79HdL3/hYmTEWcoo/fsEKTUb0QT116pLRB9Ee1tIZKfDf1Tyi82D
9wtk/bqqMQQV/eNxVzLNi4bem2i9hCtSha0JLTyh4xNxouJ1/rnGeWcAHZq9
GmV9KbIlV7UgJVw/8nP8nxclqxUf1wh4uE63H4n17iRnCzLoGNOE5CqDgX4W
35oIOxLpgFyB+KwUxERoAcP6DULahu+OGMmX3+6GM3BHg20P0jfORcgzNe2O
gwHMdO6K9oeg8qWpN8nGs891gYhj8o42xmcircpGGmvNITahY2PlmFgnQgEY
UQW9wEm5XgNhpRGyhCkprX87OoLTJh+hS9Y2sYiBFdmjcgEX35s7qydotd4i
iGjrzHR6GxuoH6d+zcwXROLEEDbT/qQRfwGQfygB82tIxHRRmHYz78ucaXj1
mksCYshKX3dRyQjxLrOZ+OOYLzhAfWL59smFJhpoQK4DBYRe0mesHoI3B2nU
vYsTTv1wHFS4VfbJeIsVsUwBLYuL72n9LbDvvgDTTr1AgGSR9Z5FRztA0ESy
2ARXusqzBpYJLnnfF+pkjb2iygdRuJDsqeMku/0Q1c0azq3k81MTdT9hhaKS
R5+G/Bo28+uxnCQPjbF9v0BKUQmy29ql9oWZ4MChICLtnX2/IBt+ASn5S4g0
92Unp4YYc2o/OBwzBUVBmYLbhb4axQSP2QuXrMvvy+pKEWprGcwsndQmo5JH
LwdTT19BMmMsA+Ri/g7j4I2vUEFD/djWzuNWV0YcXE5X4eR+Ec61O7H0B5R2
3OzD0JyUDYiU4zmNtsM4BX5N9L1YmulUFuEcxu35mBB2/9hxq1Lb9lNUZWb6
awvLk2T+9B3v/kQXfJXxf/ikhQkgn21yzKvg1lppDyHUdwFrzys+rMu4Dl4/
DNVewcUfFDNEB12NLRMCv8YzEcL13WVowJ/SvuSRi1fNwqoXoWxWFh75nuQ4
ldDnYJyFpS8H4TExGn9jGRhX0o8CUrZ82CrGgernS2QfDuvuY235UaOCfEqz
p8BP9gRSUXNh4d+87xWyqh3QGB3/ofiaY6c5LeruYyLUQoztGm9fZr0jpa+m
w2qTUpuBcyzHeU6oXe7AkGFqnxcCCNr7eWLtsr8ITY/HtDYzh9fu3xgb1LgG
uRXpIPG/ysXPaLpgImYkUc6pOaxGtY5R4YsmmHEcVtRtj1vXRHOKOd5sLGt+
n9UEPaUOwCy6bhL2MAQ+Hy2pitSshL2kSOc9UYnbHhVordjWyJI6slOl6i66
Zg/gY3JaclpMl2oMQwG/irpQ+QcY3/dk7ypKqGibX113vHuGzMToQNbYAPfV
gN5Lnst9A+2ha+AyubwwwJTY23e3PcwsyLtsbu0VnZPiZgoQxHMnv+K2uTTv
5kITx7h4SCX1GbcZH7OURBFFYOgWeohuXqZd1/YwckXp9AnwU2rY6HPc9Se/
lPC22A/wZN1tyKUMbpa8MhGM+wx5og56jjv2PYn2O3EOTTsN9h42b2FweSy9
bSm99uaviu/ti+pQUKoEaPbmtAZn7NJRBfu3PrRKk8SnZxK0NnPE6LRPADUr
IBjedufd8ZnrmaXCbAI4Y+sZLhUUkAOHxoOZSr9vuPH3cnkq1936p94mlS3N
fOVB5WH1LrmH8wkIE2SHXiXBAE/JOc/C2Q7ahaJqWj39S+otLBy/4w01tcSo
dj+t9Sv6n8JnZPMY6UdVveRRLJLJJECql7yAiXlfLu1NKGPAmUxXEj6zJ3sk
c3LMq0DpI6m5fLXqrSMahDA6oGQjCbBCTJhpNVrGSwZRTWQxS22v5f/H+g+1
2PHz2CTPiLml6OVkwLkCl9TUanQaYu5Xd0clYtP1xTCHk6mX783oViTCmtoT
ypJGHb1/+uTLo4ZivW9FKkEIft1tvKhw/Q1Y3NVTIBRme3hq2wxt12YokJVV
UXqqWKbZpKEBh61emZX3to/jLxjt7HytqCnWLSb8hS7xQdhO1QQTpioQC1Ux
lExtOoaRJyZowaFb6ILqBim4zcr0IpLx7VEnQ4bl0R/sd96wb98EBNkROwjX
TMaie1EcFrSKjr+53IyKap0tpBvFewNAx1rXj4y+PLuUP/qERUAR8gOhQAvr
GjqQz5Mo0KrmNT7MOV3gouw5VLOO3I5a6F3o+7+vo+1fu3kGnbMYOzsyWk8M
ln5OJ8VpnOL4giGMevZ/ztfgv3yqDm7kolbnazcZ7AmOL555NTglcumwJVau
iv8WhnCPOQ05Zs5JKsRoHoTvxZZk0DJZddD2gI8mWOZGKohLQKzHuxVz8QRs
nj5q1bxMDBITNHoIzzY/B9llLv8EIKehXkDT7BSP38nTdg6AnMXZTeXfi8vJ
M425HMVqdNla0nMqebsNSRqUYme5aQWB1DN6bwtg/w4O57sVeBSxcrhKSDA4
D/0VUsQMzrOFlr2ukvGaF0cZ4jid1cgOYkAnmxcjtP+fv+ktI2FpcfeARWQ+
Fywq7RZnkhNjQn2RGXYTgRLRLSY+2C/fKJpZ37uNqt2nNMBH1G2iY6o6O9XZ
3kCnCXD+zb9BUtD7WtpTNTFbEJLUejdaTjf0/S48tAHOsjwg06NUdhLSEp4r
K0vm7sq7lt+9Up6GLB8doYCYPFdQlBUtxkTu88uoRRVQ63NvtQXeqXvTmRsP
pe+vTMoen962STBZ1Phl7nFVLzUdHzkb6DlZGXbLGyjl22ZX/Af/u95YOLxb
/w7znZNQjg7O3yvtya7BXSwkw2fMNklT2AZTyOdNFHr6v7/hExIYXGG4Vc5j
zc+e0ZcNIRqcPn8XcG5+XBcVad+9Q+yUpOt3bSxcAbVsTALqndDbwTvStVcX
/6w1PTJejwE/MEF02hhiYqWYHS9oeC2Sv2bhBw1M498vYh/rUyPMGfpYBdEX
dEcP+7oCgENNogFhR+n8No8CyacynFJHR15Wu2DZEzv3LQcoRYC3ZBW3pgoF
rys5+NVLDAVcYzRJDM4FZ8qm8fAt3rhYVNQWtkEVpiXXQAYpOYdEfEs5J+QT
KkN3aAWH9PDxNA2hyN5YMF8J6kj7R4lU6uiFYrZ+d/8ts+Vb0Ov2e0grFhZR
GsVyCcHat7gs55mgArkHgGa2gF8/pcn92JnCPwy6aR3BkOT4H9/7TdksRgUQ
xMv7RFoKdHKDvnwmv3tk7gQ4Sp1hzlcxWnibfASze+cOqhab71R2MBi/ia8H
u7kwaPDPbr2sOmDG1bs2f+vYqbuRXFbOgEBa2Fq+xR7CGBU/rAlDpK53o8RF
NpJGZoMMwJX7Tq35f9bC8m1xst2gGOWxKBoEJsz9oeW1/HGzJWloz9LpiyH2
KAWE3lYZunPQsI0xPyJzmOV8IjEWsqh3lWQ0XBrFPJT/gqkYNOFhRhwe1AtK
A2PdOuH7Fssg2RdmWomUCdh26QpL9Xlu8VSkNomQAisVtSktuJvJ0wZ6wlyQ
pPXlzigvT1YjAzs1nocuG00R0g0cCQ/JMRRRcZnL5pcMrdxWYRq3gG82EE6y
9//VwelbXWUeP71lRST+0iD03UpSGJGR4/ch7xKKE+VV3LrdnpuAWpcHZ0M2
+15Ism/Fr5JWXNgqTziHbWE3FVp2DOg6KX6Bc6tj3PSK67WI2bDU1UbJxBdY
PqTZ1+Y0Hkade96/EUmYJU8i1UpPELERaxRZRRhpZybVxXrBdXUufv5BWY1Y
/PHxI9oRl/a/NwoiefrDWIvGZEq0zTD512PGxZ7HeH0gGoCgo4mPCYHClVUn
Ne5VdwQ/jOoJ4K6g8fJ+S7V/OKomDw8go+narfwUvrzPeXKpDXr0rB+Xm24c
czdFDo7QEhcntzEGUlovayU7ZxFouHWhUL0+1kGuo6AB1GA5cen0Car8MzuT
TD0SXC+V+PJi32/EPYWboa4sjWolcb1LQbQ/V1bsKc5ym02XfX+MB9cSICo6
WpIO5OgL+3dXkpNceGJNQJWfI1De4PI8rQ1dDaHgbECJ0bfwGx7PsMe15Dwy
h8/YjeupTwrDg/E5K9EqZw0i5vzsPK2O+A91gZKS8Is0YuuBe3c8dcqATdvO
C3iuWQDS5iJLkRM0w5IM0YTqTzzJG1p1+NUaS2quqpyfwXZ4lhCV1xJLICCc
5NDbBClz9T3YEYyZQJtQioXSwQm0FXZiYqPrx+oyNmgQvA7GiAQEEYQlyXm2
VSfF9YpWfL4WoCab85eOyXdkROreOnlGwpapxKlrcHyEt/2R+KD5tXhpoNvZ
chqjjPpX7QK0l1MKPIEMFYiXiWFXSmxNKw9jgiw5vSoa6tmnq5HSKccdOlLh
Ig0rzFHtTP0udrjYRcONg/T3+U2uChLIzg4x+Uhvl3LupY4CjyhPqtSVGuz9
OFK3DSwuOOxtrS60sEcTu+0Q6xJbVu2GlwAyDDb8N0j+DNQ84uYfu9SZJuaw
5WFZKP5B8p+tbaW9In0eT36vwRjAya0zKJFVqm8Cec0cIS6J71gbgoCS6nsS
4I3NZ8zkpldv+dd0xY9IumIrGWefONefjuNvu2GAv5UjBvkuWWqCgmGjfk91
mJnQ2YFKCU2UD2hRLODMpQ+E4Kv/5n4jFyR55jf8Uv33Cujk4NbkMcF5H1h6
mr5BsKXCWBjzQa1kS/m7OWODRJkXsdrButOE1QUvXjgoihOh8mk/9OY+2VTK
ojPa68iCQAFIkiJhobBdjRFhDRcmeslAumsJuMx6PtbJAWiyDqKxuoKero09
WELg2tlB/8RP2fzXLu4Q9GSD1KfNrVuU1hgpJbVAZ08yODLCMx0eIACZ7bbt
9kMz0LzkPDNZSIue1yVOPQ1GLvL7/9PLFJnRPbYsgqF3zbM1sUKi6C8cYpBY
sO6WH8KVxzK1QnlmrWPLR7UdERdA74Lpz7/epappHSrXD5+JuDdDakic2C2Q
a9r3WtmvA3I+Neohx/oXDRUT3iVVIXeO8FE7gugFf8Ccq0usarVS+4J75Suz
Kb6oTUcKsfVZWlgTjBNZz+DPyQWgJaZCUHKyYtnkR7GVAI7cBjwycXfa5XX5
6JN8jgIOd9IpMZA6Pf+Wv7ux/YZvX8GIIvBYNxEKK11ZkDer4MId9uWwvclj
sNXM3MXf6VtOLyUKx7skoYe/lMM6GGZ+XNJ1FQz9vJx9Nl4bE1+ieGXybg/v
CkCbokoBABAEfbFUNDJaoRD0WGfhyZnnnWzY99PDPCDP5kcZ9IG2HHfgVT6E
js7loT0NcxqQULOgnpSNo2aICLdo91ra+h9CwII/5HFeK5JsQ7Cf+aH7Qn0R
qbSOzroAuT8rueRINQ/5sj1gLBibxtmRz3WMXHrYtrLm3tApNzQLv863EGi1
cJztEHAkpgrP/heN2WfCAbN3Ifw6yvGxI3kSbVK5B0FK6uKFmfkfCYGBJ6pS
il3jxIyL0hqwwZ3U2h1vwesAv75XhV2K4sYSJxZpyVFKnbk5Kb3Sp+kg+OLf
tX58ilTd3mOQsbDdCmOyhgFq623KAsgZeyLnfH5/jJTZz+jyasozWaylNTyC
U+avQqMsPUsdROsSzZKH8Y4F5jN66wGgF3BtthwCGW6y8AErl/pEXFsEDnLo
fFxGW0nqCU0weRm4EuNVrTZi0yHRwUv3r5m9FHj1o7Pgnh860+5KLtpDKcVL
ICYj9yTorcTOV9sg6YOyv4hqNxXWByXhW35GYlPqLbDt/8dV48gxEZJN9ABS
YIpaQxo2M0AUJzEr8Rem1u8wsnwgcNrdlapuArEnLxp0Vx8CXBOHlKdwSwEx
9z3xz+q/8VWnR+oPq2UZrxT+i3ReyhoLvWoei3wrimolA1B+2sqZJqwFjmTl
tj8JIymCikhnRN1B61d1q56pP6oTI8UtovIN57yyXPPvqiVoRYE7u+sOPWyh
AhQXkDGT4fq2poT+LxnerNueTIzHwj9T4IhdCRGDR2QBHt0P+eBw4JP2n9Bl
SqnfSvWaB+XIDu0wgRr1+4LQBr/Kf8BZ9E9CuSVSdGA0TtvCCeg3oxfoif10
ok4BKdwBbjMtBH5dcoAqbhxb2RNTr8DpRLoxem+62TDfgXWS5Yu8ZPf8aW0e
bZ9PCCiP/xqo47ZcrnTvi7Mw0e4V5KNDbdc0ukS7lmxuJqmKKCO6Sst+HDV+
UaU4W/sIA5Wa1IUSt3cGQHF758S5wu260k3bUgyetkjiIEkT9oKai7Lfelpi
2aEaQD+6hU6ECRtjHt02jmCoq8cxlH2+oHHqPT6vESPcUApj/nycwco37F+x
Mw+zNl3yIlUfZbT6/emFEmKVTH5aJkEUqhrmMAUUjcSMQWCcvG8dJ/+wDhgZ
4fnnpaL4105RFDLhaseHgP8+cIjd3+FdobW5OjfRHNix5Z4D0/6hjmLpzBds
eMV5ilF8XADBusrogAya2I3abf3LSl/tFsqIFYSW6Nk0vcJ7zlZCpyvy7ndI
55GZc4Rz30S0LhuHKUy1nmneFJcnJh3s/Ad7EcPOI3ubn0Ad7oNQm1/LBY/p
CwdwvV/kldn0d1t+V/I/WQksvETgiYRg964HvaBH54TZ2Y9B96BoLXWbfEPL
BYBIEoBudt3d7wcmxUHcC/ALu6U5RkxKAYNM6e2GxdM2rcPoTw5ws3lnFSRN
OZyV/fFaojkosMkQJA5ROeF5A4bKrXD6tmM+UDRvwHF+JGTt5o5yJw1siPvC
PVySZZ/fFkP+rn4u30EtfOJ8t3mIccFqSDf7ICH5YKaLiiF7vT46srbSLgtU
BjyVbDO5NzWKJid46OLHcq8/mgud1zT9isVBE3b+WHeLiUOFCtIwXvTfopnC
XaNpir1YKS7RQLDvfC2U2EQzQnOOZGyYk9fpbInTUyhsGqaPyp7ahEkCYteQ
Wuq/tZHNkZuix0dm7JKQ8rrFnxLkB+TMHVx6RPUB9UzSogJhM0Tg5ze4nSSa
52d4xa5l+lqA8dW/6bemMdxCaOTgE2cLSo2iMVqs0yWiDlYk8rT1Hg/1jLiL
MHvsGQhYRdBM2Ku70fAV/wbJYa4bHEPGbil9ZUsx3oINsfFeQkeafNysHNm2
OduvavK7Y3SeW+I9Dkp7EdoOqAqfMoKE3e+LdeYzYsvEez+Qw0huFStjxenv
PBsI9U5foYrgGu3dp2I3/VgNL2AhaazN0n5eQzUeBGqcFZTUlaZCmgImcCLJ
d3mNi10xNRraa9OQcjRwCOO9zf2ZnBho+3AVGyBF2o1QFxbxe3JAMZeyjEi2
+R0HOEU3EuO4aOS3k7lNJ1Xyp1GGdUZAwE8lf9U7mliXExivhlEWX5WcOu29
+Q+fWHT0wVfAiPS1AXyg9UuMb2VJT+g7G7aWQhEXynFOZYTZE2/Aw9YCxRyc
hmj5cIl4UN7eGQspNVUQgylXXgva3MSfKdGUsz/l55+SAGs9bhdNBg8lG2U+
04pLH5WKcO6YweYlrMpHOUu9Qd54fYMrKiUDdpf+Qoahetipw1eGENiyrJbQ
oaqMdAGDVf2yWhgf6rOxXJitTykdqbeMAiYYVnJwOLVmlZ6/uLqCCH1qZ1Fk
vVwrXlJrhqlZehimwZTSjbauTF/ZCzyb+7B4Q+ufGSHWWyZk0Pg4v9v1G9hy
UeXWi8KdXZXshwmDTWeuF+ZZ+1FucvwpxJt8PbLCoEPknnXwBGl/KXMMvJz5
qEKeUndryJfVph9NuKMH/dMd2BuGefJbV/JgtNoLjpWDBD/9jEOjEUqz+kws
3kxpfyl3mima3LaOgtMyHxju/nYoASzmVhGAsDw4EwZXRqoUvUtE/32lezlu
NfodUemta9aLFvui7R+CzmF8jyIB+BtetxQj11MGGhHmvjx1Asg7kSmZTWcZ
MAtG3m9MjnwtNAtRt7LzkUsymx5N97A78Xw66DeUCxysJ90JyQxNwYBgNiap
fYFupQyrTF4ybvIciHCBI2spRuftYYk+pZ+5ymEzwGwX1wsKw+CWSCF3zWzf
Th9JqmIfEOxBKBK1CODWm96Su+z6eimbbhd1za/PnUZFVfzFQNpIQ8wAgq0g
vcVzq7J9E16Zm9bH37jPfaDjjLM4F17IQEYhGpuJm40MFI3KG46bZ423GE0F
KItEWV++FHdAsMeMXjrfoJGwDZ3xt/JbuV8wl4ru4t+XFDEHuRGc4p405lV2
yuKUyH17wVmmqKuPwtBMx5/3YF1Llre+H+EtSbjr0yXFFIBHhwOq9m/NWCYR
+ggJuG+nbQEu16K966xdR3t0hQzzaONLw01jhOMqD6le8SOJdnfR9ahmkmHZ
BYoJ47gROb1RDbxfJGYRSZBzjhgzgz8INN+KziztbBK1sR6BED4EQ0mmMqR/
bS128kXAJ+HEG9yNuDnWw119H8uhM/e8jN8AxSUZ/UPaOtM8Yx7w6nLg1XRK
GsM268eTge6IfJ4ozHI3q2S31p+GBYkugx5OUQ5ysUKaVRedArCMKOQWqk4o
e/dY4IQjwUwDfhLS4Q+omGm5TQRpmPI8VtOzMOdN4OSHhhWlNi8Hxvqwyo0M
KhyTKFelToGaUqjVTtf1B3ETyU7Vt19TF3lqU4ZXHjxMD3O/vpPqX3tC2mTM
UJJ8vj0oHIdI4FyC24rxDsxU1O154cA4aLomX1HdyJyQP/ctlLBZDP0A1agf
SN6chTnIPfvYRjKGCzRr1skbGG5yUg/FgFisIUi6eTeNojczmVSsn7WPBXO0
o+Nrm0JXRDxxlIVizEbDmopEObrM6zshKinhZ/ZOKS+1T6qyanpkWgB4y9SY
+NPboMeKi0k4e+kIoHq4pE7dnOiraRcJz2u54a9wZr622diW3clIKEfNhoca
+XUTLSQLe4xPP9dXUlQlqUbMQatgIGZ/CYtWhoJjInwluaVFBzVPvIYSVzdO
CnxYjPFvOq/hPdQ2bjn902EwAd0J2TMletTj6wx88qiwVkUvPmeGyjtLUo3b
0iPD7Q/YjZ/qSiK/X08VNyiW/dtuA1wD5+Wb5dct15lleRJ40yNhpUcVGeje
6gLCFcMEy/Iq7V+Dz6solF/XSRYqe4Uo0qF1Kzp/e2hKF10u3w5DUV2GrxcQ
SCBVbFeK/NdwETVh0wDv6gCsIVppJHkBsnOOaUtPsVZikoSOL3xnQee3S9B9
VI08qx4C5alhK/qs+A6NE10VfYuojUsSnTDYmQgW09xKCPkBwSzj4VdAcZCQ
D+UnF1QrOZ7AmlxgifukvJs14Qwkwf35rC/9UVsVG6QSYfGTbi7OmSChtZJE
PfQjbm8NNRjUdqPYzC8sYuT58Q5uXoOe8jUxanC0T1IaWXHpyoXLz97PFuV/
jgFzJhkCOYLhESjoe6ij75D3Cl5QOw9ENKv0/HBwxbAWekixKqsONS4vWVVE
8Tjmj/FInjND1esqeszkLPC+NeNvnvPQTvEcUWfYXpHTIPzzkRpmyPepA/uj
JRpJOqSqoM5bd/hKlluYOXlTfJmrYTrURSlg0GSl2cJ0F6JPtAaZU0fXIqDZ
kCKijqJXlgJwlsOLsf/XeDqsCa11Xiyvq0HPRVUDG65SFFO6tjXppDWykqIs
bFo2k782TwfcEejfHIKuGSeJfzALVDMiJkXc7TRmdlvkti0kPGciiqzTR59r
b3p0zrk5ypzhHGtyOK/+Phwiq7IguQ3edo/qZEdk5WY+EVyZBSeslBaOlOE8
bifuYddJHvHeF7Ic2lNh6FZRtBcmoi8LzLfTRhjteouo0Y14pDGVrNvIZj6f
NRFpTkrI7R8syo1Aw0wDIsoAbGMdDZWF/QqHRir7wTsVTXd0/iDrX0H4KxSN
1Aa5GfpPDG/Qy8llUvTNTGf9PETD73UrrsKKEufuz+Z2+KmGttI3UJL3XU1w
iwmhEoDxbPBI9WxFAYBZhJp7mUg9IxIZtOgQDesbplNHIFyF1kDPjYkReZ72
evP2BroLlEicbWu491g0AxXDsncdyM0eAZZxlYmAPzR8pTQJUG7nFsrbJrgR
mlL2BaXHmnvoH3mpNAKX4L8LHM9IfWjpyVHi1mrl+OEfPq4lqk+dESatItCJ
6PIvQ9QDzukhe40CwKigAShr5eJ8upf71Llt+U7bAbno2LEINF59n5q4mz6F
p252VJk2HVmf0zI9XXkNg2WR0CQl5znAC5XrwVPyQkL6BcpVkFAcOcZnZ0PN
68hmrTlocNf8HXye4D3RTRHqRf3tU4mRkKHys7kGE5kqSuCD418G+B7iTt2J
dV4KYYHHdGg+Q9XOnaET4IaZzBPle1xjOSdL4jUC+u7W/g0p0xf3bCwMSglG
kxifq48ArviJk6MibWjlhSJhCUreZVNDpIH8wZFd/LSENVACa64qI4I+CxPR
JSACnsdq1cDWV1slaYQQS7ARM8Q9bFh/oKQUo6wE9zZmxnPSvpZG7B7VETQd
c4AgM4jK/4qrOyn/tFiGBkAuRhfjVPTjQhAe0kUnXNmfNNS2XaWbwLvy8FKu
HLIn6am9Y6onpfa9BXtpUitvtDNaCT55UrHDI8/TWmoF/VQxhyjZ2RxoipoU
2e5IxgawvEaa76/g2alnqGoO4SyCNtFh71vQTSuiNUqVv/Ne3YFPRhgyN9CQ
h+aLoYhqKLVFtbg6A4DPqrLNgxqdNIC2ubqfVXaL98H8poN9qi9ExsMaQgEm
alu2XYNHjeDuERK7GjQlIw0l1QLPAoY9znsSoNKin6RLxTbAIZdbZwyad+Qj
KCTTuB+XdJNyz+9CF+C56o22t/5KIDQVh1xNFiSDcT82gIn6nMUdDZgVSytj
WP0eZqQDqYYszXJ/nFdnBal6zcP1W0tGZFJ3LmhfsbyiL3VyIZbr6B7iBVQG
Owt7CO+TpBflNB8SWfsOTbnpMZYjC0N8dr5kuwbNUMokQnjzKMJqYEV6h12z
Fdj3g5D9uMlSARJ4BqXZ5V2CiuW6yUqt/8V68JHAFLihLOo2v7K2k/x62t/k
b1cPSPt9az3HGeDVkJDKxzRdXBfDDManxaPzl1vb4vuJnNFpcBiBf68QKAvc
zWXknRKeEK+VaIqK75kfG0FHV43nkDGlXsR2K5xZV+tMImxL3PJpU3Vdc+/P
1I0xXpqsu+AMc1SYJvQUyMuzUnb3hlMAU/xVA8Q+lj6TuNKSXEjzccn5kzUB
p+TeIXV685F2anK16Lr2ulNki1c5zEuiRt6q+Yx1CfmU0dVCGO3TF6onUxwf
aDICRFBxpiQPcfwG64rNDy92sx4RkRK4mHqsR0v4+LJ8kh6Kxvs1AFiL/T43
zWNB22Spwfw0hG+2gVC94frM/5Rp2dFIQuvFB3HbhnzB9q7VATMjATwt8fum
h+k4ko1+v9H7e8VTeJFeq7Q4b4FlzBd7F07bNWSPKPFPL2/3s9+1fPh13Zoe
AayapYVsn3EafY5w1XSKC2f9y0PX5+0Y7eBDk8Ze+e8oYcuYR96Eq7v9zHWL
1SnzvHIqD9o/r7rjOmV9mz0SDu16CdQ+ULlkIJbicxgdPJ04I7k0clUHABtm
fsF9Krap1d2Hem8hCnJYL8sAi/jwyiR9UO9Mj/4IL1HHJwoI9NyrRtjwDubS
wMYZsLDFmtkqrgnQ5q6+nmnVlpSfknMJuLM4Zht73dRL8zcJnywOOj6UfDey
sZJLinl5FdyWq4Pf9dqhRQBY56ejmAkre29gtRDYQ0GVsb0nKW9VS4eV+hsN
L4pPL7YkEZV5U1KE2vMkmiV858GyUfePwLHBCdH4OzJEO5wYdtsedFjxw0P6
+oFZTwFOW07HfljXlhAAyPxEifY3VlN+fhNDI1XJ6xsrUqzGWXGRnngpQDMM
L7xgyXpg4ucruSyjQ3XO+aYqo1JP1sNdDhwC8V/hOt1g2K9QZT+MT2a5Y5e2
pQcB/4QVoYNoU93IO1iva9ReomEPv1acPHBHL4JPbWsl/S7q1oogn8NVOCZE
ilhvzYzafoqNoVZcD68VBDfniLz7a3z/t2YynSAOxEvQjDodieGC2N8gFsjU
TSP96GLnQ5bj05lAHWETkiaUuXCqHqAIwbPzn68rqfsHg2xuEMGM7MKyuSj2
/t83iHNYkdRjuI+XBsGOM+Th40RoLcIYYXW/IM5S2V7jm4iqlyMaehaVkHjy
LeBjEe0c0MuCkPGgJRgfbuGwBT4mlL7yvNxepDa7kAGnUk/ngzBW/dH4t/d6
G4M6e8EuQL6y9XKjX0YAgSnsg9fqU4kg+SXmzAd+gJ/Jpq3lZWfn36E4vhoR
XEmjZQ3n9Yzvt9TJV2xNyf31f67HXLEI696Swak+Pinmd+FnxiuQVT/cSBt6
zXyVcocsH9p8CZUtJ/WLGldN8tpY4z47stP9m4urtl1JrkqEen1S/qzPBuM/
0nnrh+hParDqxrXDJZk1Vz4oskMIvjW6jQLRjc/KtwuNkssukV6RaM4yr2+p
F4xbMpl7ORTJBE+YH/YWgx9iyv9liiLK3bldSgnSdCrR+pcty/ZAMsPV5tWU
hhVSH0gRlfPhGRLwYsZpjZ/wMepE1Uu1XilatEZyuK7unHyiU808ASgPbbr2
lFEQYvN/Ha+i07GlXUNcwm7TPIScFgWHIIdmhU+pHCD6CXQn3lABYzKp4cD7
IEJCY4D+lNJWF9NpFvHY1/VYWCB1LvszXXC2ZwySr0TUlil/ze75vdAgTRNf
OJ/9DWO2S3IteNnBKpa+r9N8IcZDp8qcWsWLdDpwsGR2dw6WmyCDTaOKKWFF
VHHdx88WVp2EJsJU0kjaXpn7MvjA9+obPwap0g4ONNpgd5FQ9B1tXrtLQPaU
IwCjGenzXklRQ01eV9tTFlcCV6nA+317rZmYMygdRp1rBc5mQQl3zdrdRapD
+7Mgj4PdngAaXoxcH21fDS9p1VILKtMwQa1rz336S3k8TQpfYioKPQ648XHH
sm5FQpOp9aS0tpi/z3ALiiG6AE5yOHz5iM1sEfxx1TqUvfYzNHoDayaew4Ti
v47C7pYp6KpilLHPVS4dPeQoRFhSalnyaOa9Bs02KacrckIVVXiXhEbh/iMR
U4TzTxFVu5m29wlrWpCxStubSdDyPcrvzUqz0nTJikeNIws662R55J5VC5gP
gHY6VUEQnboNiGbecPqN1PdONNVFXErR+oKeixcAgdL3OAMRdbV7klOUtnNH
eUo26G7uL6IHYwxdBtuuFdy1tltSTSIBeTWDeu1LNqe5icUXeN4sOz3xKtcP
zqJuDnv0CRAvHx5af4d0gITq4aBazB1yc/o34eo+8O1MmXOhK2l77kDmHIf4
wp6cnDRaTGkVZlrSZZ9n2AOImAw3mAI6dfXcT67KYk8rNTzqw3umaRbyY8UV
TX7H5DVyr0azRz8JX/F5ZlWZqH/HZH06+rcyrbbgBxLGyqkLLmaUg1yq/S5y
R96YRkTNOAEBjIFVqBx+9i6aCn0UwxhT3DJ8NSNRtVRGyWJRTG9aU6r6OLC2
n0b2QgjaBgBjKQw+kag4ROVOZCmCUsRpNCi9tyoMAqSWQaTDpgNT5mQ8N3E3
Q6DhTUNyF3/JLGssWtuvkZ/QlLP5ERB1ToLiljbv+CNsBsFfDlj+3W49ot40
CL0/mI3ucrPe2KQx9ibEx/vsGuW0uBDOwZoR4HfGKGWhiO3pke+vJfv75Q3C
bT3kYvpvJZ2A4RYwQ4ZD4ePzFlGjokwnoT29tbcf470wxqpmeHCIcvkS1L8x
7/LPABlLHgLKtfFaVRmL24WNc+ymo0/BLsweM0qVpyeU+z++X7MQq6WD+VeT
ciGdOFNTly0njkM5Z29K+Tj9hEMYVypEh5VGRb7WrcC7iXVU4nfVZiwIVOFI
l7F7QEJ8MZP9d7ahELFbVVR0XxzmkLFYuXMl5nYHgThMBaCyt7xBxwMVvvlf
gktBmeNRUpdTXr/3OEt9GXU7auG5TV+Tbh/EwTvg6tYd4bxthu/Y6jmpYnOV
TU4blhNsA09byR24Lm6PKZeWnMrUpbDuYlbgdC2ib5DlzfVP87VfYzkafONt
haa7Q+AsCNMekPgValGEThxuzvrarp3lUkXev79BX9H23tKVidmDiWbeVVOs
upsvJ3p3avhIEABsdi/lTqFt67VfNIlU3WVF4uHjjrBDbJbekKUMKQ4zsVMm
IQDPW5oDPHqXRh4t+AjIApRk2yT0ZSSJXs7AZDqovI987rxxGD7lEzNd21Oz
3iS+g5u2ONAib0Mv7oOWamQapy8O5Zj1VBkAT/LExCJ1PjhIA5kak/zHzFSj
2MFS8+5WI3XkX/OTujNbVwX+HsYr1TETnzNtNZYll3DxxbBzpJpfH8UvHxS9
HNRS3dPcG/5HYr9N+ezeJI8+tPn2nmjElZywNKBI3cpnJLrLI5Au2u69xDAt
mEo7Ji2XVQ+GaXayafYlLiL2euWF0mitN/kjX9oYgfumgeHI28FyngjqMm7Q
4ia+VSG3qkifS48dh8GrbMj1LKSto4rtiRO9LmJBVB9P9XmRV+Vjl9ItO7Eu
Ugil4J8G0E3ORMfYulv2Ep7GIFZzZdL35ycYQomvYSqVVNcWor3/tBo5OfEZ
MFwUx4RGFx2iJOzJbHUVmZxmBvXbk6AHopxwnR8FB8SOncRD43rgCV9oimED
29CB36Vd845AQ3yivDTqP1ZV9W8Th4PFmljYPLD+PHthHsgjHWH1PWdy2z89
cmef9j+lLkOyRMLcUKUbwY6Tch5hfe4UQWQl7svm8mlTWXxKPqhyREW0mjYl
H2vMWlsXV283l+UC8E6/yhPhKe56WicxtyU3PAYE2R76hXniHT2ThnzGqnc9
4CxPBCz8O6M6a+yYDh7pWjHpSZboQP2fDsBVQnYgaqX4oETWCjtuAUlPz7xA
Z3k381SVMCl/mtX+gFCF4cQytoJ39QBVn+3BFdG3tUU0LId5giYlzooFNqDS
eVMfcPjW3dCbNMsLqkPh91RlPmrKFWy8fbMzDP5s5BlC2JV6YPx8ZAxZjRnq
/VnxyZxaabgclc7A9rUUIPWnjJKQKmUMsArne/7wouiDSOFvp3RjpnOjXDcn
E8EG3zSehM2zhMgO2A3l58hAZuFSQ2TZSiRNJVdPN1q3PbrnJvaBZ31xIruz
MhCxnEIIENJ/TpprPd1F2o6pmAHzF0pNPfcTfzgIqJOIxpu+RjhONzkSm1WC
nzOHF8aMMjcSywMIpEzv4YyhaZHJlY86rP6PEtzBEB39Q9JzJ3nk7TDUtgRq
k4h8SAva+gYvWPJrWnyFQu5lXhxKpWkwg9vMTRrBISLuHx2xqJhnQQYguCBP
ujE0g5uuxx/hCcT9EtccCYIFAeBku7ivpdSwibqwfRK5p3gr8ZKsWI69RoAZ
pmISHuSXcqpV3d7//mWsk2d24icuNtgGDbhv80Z7gnBc5s4v9W8bF9h7idrH
sLTuBllo9HMNI5XTop/cVELfoI9lhufxBwoecNggjSfVeJ3p4Uve5camIpye
6eiSQsW46i6lsYq3MLYWe+uNCTg6TNHOtgaokBILDvIwMv7btvci56ZyUfEO
hnHEN0htEtOXfiG6fs8YqZN0X3kZSyMS7e+175Fpv7OhcJCAJSKj6TpeCej6
lL70puOW/SzmZUakhPuwhTjB6qFo9taXEMhkca+uu4l4g1BcpG9aamPwg4xl
fsc5UWifngKKZJrE9em94hdwr6+vOZSaVPeepdj8VJtB9dKao5S+hSf1ykxY
/pOr4a0jHmNsQyev4Z2RUpasUhPMakzZ4gpSJdaKEjI8ojJcSVbVC+M1c7Qv
PpWbLu9yPpkAlQeMTe/+xDAMuDlp9ns8O5eDciaLOKXmZMjHM1jU4/H1EOcD
BzjOGiq3VF/cMQt2f6QvZgPFShJ2sa3s66InhJp1QHNIfZ77thy36gXjb4sm
BKi3EAdXue9HId2rzXX+Gf7/BsSGjE3S21bpWZWEZvGKfjuaQRFPPdec8e9S
WRNbzqFT1430DY+Xiunvpq1UycXd2Gou/Xff6QtaGj+6T76zth+5g0T/Niz5
3phurqPn2UHhrGrpAAHAMURjNo/97RKwqNnjpN4GsdtgmWJxdeGxEJoqHzaT
tQQJBz/4elRdb25dfpBAKHBwsL2uW86QJ6r/SCrPlNaKjbgF9qs8jgvdCiT/
6rk5EMwsibcLwjl/CBVfpLFATtDrPMOnixYB3AvLXOHijU8v1HFHkC0pMHHm
Svpb2qtfMJQFEew/JChmHVF/Oh+6Mk2i8AOSZK+9WHgU5JiQEWhutHO9JinI
kdF9UhrrzDJ2QyVGTryDgrCg9qZmfmb4f2fJquhw+GD+/9cO/wfetO5YJHWN
64H1irfU7m9iAsj62h6XpZuWWP6iuefRLV72aeTwCvib8Zwj9WBnpiJ0IhuG
Kvel7AsmKNhvr5cytW//n9Eeq7aJRjx9NEiPmWOZ5iE7305g3cwWhxhfBuZK
jVc5BASmnkDOfeqeOstOZykD51o86y0nIuLCIYOszJP6Lu1Fb9Tp5KBK4+nT
XsWoAKEK++wou2OUvUk2O0nBG5zpjaS/5gFAzyX66cePYGNcZZEVkNok7xE7
b3eLGg8MhO9JyJ4vTj8v7E/xAER8uKM5QuPwxIxHUx/rQv3U+S4i36EhC30t
NpL7kBckiHEfl7zOjSQ+OGA+E3JbCuljPN9uXSMjhE7HPc3KWdjEx9QHPBiB
zyfUJbpwJoo+6NNwblBl3zXbxi+azYjUIKixdGqvqZwKRpSnmhPDXcbCD3K+
rtqNIakfWqqbHOOIFr8I4XHWokT8b1a+BogziBHtWbwatLmJK9CHR06hGaz2
IeRcMTUb9xafqHeUNdbiLS2qHONP4oi1BCxvTG/RVeFabR9lFQZlLjXtBLXq
L2Sw4isUHWtdJSoT1j3U8a4jphTGtiIdAg5t2KD6y7sgrtCBFW1GLOFdcphX
OLYLwJn+CrywFEJIw0o6GwPJ5RSqo1nsQ04YFZQ1cjDZguLO+8L4uQTx3TFg
RYmKBzgDSwFPF1y8bJdrEIofn48yS7GNvKUEVQdWKsFp0b/rck3ixcUgZB0T
MXqZcE31APxOqc+/xvEgSIWzwd9VULkXjRfkH1Xj7EEsPFns9yY4Gal7nPlX
E3A2A2MJgwFGMGH2Kq1qOLclftQomyQWi5k9K+hdjZQWW52VFC/b78gFXTJA
IOv8U+ysaYw/TR3UvwfV+xRmB2fPI+LxmRN93TU2zzSOCS0v2H2Rhr7XT/Oo
r0JTy5bMSxdIM1Rdxprlqf0wb7koIWlvs/E7VnDK3ofkyfmEys2t6oiljB2A
ayt1jBaIKxdSRFn7mqM+/x9UAdutiACMBwYf0hSlHk4RJXSFKuJciYaxqRHR
h1PbcG931hst5pLjHoa+5YYAJbldbEzxkS7LcomJk+bHBvaqd0vwEQe9Then
xptJA2y7WZROPobMo5G0zSYCWqQP9VMdAp7j5L6Hc+GdW1AR9636MQ51JpuL
tHpXgWdCeyoOyXKTH3iRDzLs+N2NIrBvL1T2pTDuuJGnEBmAWHmLb72no6jf
h9IXUxze/5wWLjDqhYgEt4+nOBYwTCWyRz3YE7CAkaYl5M7idYyF2a7szPMy
cIcqavSToNfAdWiXTivunT82B9kzKKS7yVzMQ0kPJJhxdbNfeNVkqpfSc20a
yD0A885w1n2CuXn+T/34kyArylhbjjAayHkmKYtWYy7DGHhUONt3tu/N0thT
+iPGZ7gt7XVPcCCrO1XJrOhjifBg4bJY0vTjgqRRETxHEvkcd2qW9pajCbRs
Mdw0Xc31ZKG0pE9RB8lB3Vul1bRNqdpoLydZz/H4UoSg+AnymAmIbO1Po0HW
pIsVOerI1M+lX16ofPFZRwlGHyzq28JlTiXifT1BX6bKdVZh0CCDHvlH1t6Q
AfbP1D7MWnw0nJhLcagh/z1iBRo6N+8ZzuVYU8vgjmTKxHA6ATB+TTwMQ18l
XYDJEGfi33jUEHLILzVsDSVLSucG4NGGQ6R5QoS2hve5bSaITVd8menlOlCy
twBSPP+Jyt6NHIIP+4l6elNRPR43h2oSy7tv0N88Ubd25r9/CeuyuC7esMY1
/47sM2McJYwJpP1XutQfzT9p05hTbAWysQJsmMdwhwKbp+wEZKZ3d/pQhpna
Rn9aW+sVsB8s3An+rebjgMMQIhl3w5TpKamzavfYOnpsCKmRSExvcRUEbHCw
Rf4UFT1w+R0jA2A48rdItGDp6a2qGo4rrMy4rBjhjfhz/T7qIdISc8P1wl/O
MfbdBdkdNODB2yWb38ejAPL5BWAhcSfmwrQw4n0mYjd/jMzOeV6GQJjBPBOw
07oL2B8PV7MMHC26Aa906/JaDxak07ecUVqFYp+F8Q8LkDt4+LBFWAO6itZL
lnPPCC45OUQnN4TR2+rOijljpXzwBqxfKuk+cwAdUO5L+z1weLRRHqoPQA/B
ac5uf/6p72Ds2oiU5mkFBC/x4U3ETiJRSmv9l7rRtV1b9xGVEvS3DHzoiMkW
h8AaQYp6gIq47vI+OKaNYSxFUhKQT5bumX0a5eAuQ0uS1t8Uuf2AShPolOWr
O9UyvIvt72AFrz7TMwc8aJ6OrwHh/cFIuLRfjATCaakEu0jbfV9diILZWPpu
yScwXTwuEMgNXKiDGhNdaXsoqgLvXXBrTAN2A1hibdmz25q4Y1+8+SxyZdKZ
EYEFSnjCnULLNxpXBbAdl8EjcRWFx2bP5UJXDT8phPF5iwkZjN5vFcZkR5YD
v93NU8ADutRZisyERy/olTkiRxiAmliyEo1s/SkOEWRDzUUAErxsNJPi1C/V
nhJ1HvmSNuzwwyv9DmewINnLHd210pWlp+DYPSKVRAQD7P07HQB3DxUHQVMp
2B+VxsAYjnjY7LP1lQquxhaVTF/ympSJTaiOzvRQe/dL1qSB4DMtD1srCycD
O1LX2ZXKHIIOc0Z/w79CR4+LnrwSstFHt5HOMJMrF/dfX6we/39nqg19F9YN
BKL45PaQqxhI0FmN47uvZ60kG2Mf5Qynbupq8agHRCgOx2XhbMAkm2brJT+R
t9/4SOekENIEV7HX34a6Ufgn4/iTpVBMLOD28uReSg68Ix9AmGIdV1DYn7TX
T9k2GjamiZO8hFePlrDtE6uGFZi7mf10GanVTuj74Xofaj9/Bkw459/wvTXn
zhm+p5mpFhvIcxTDi2JphekrDYdnve/W/kbMPIwmhMBjl0YNaLgZm5y1GYcj
FGB51J6UcfneqDCzwI1wTBmvniWTYhsAx3KJxAht5QoB1IFJOFvQ+/ZwG9rp
rC2YtLVf0brDQuxIuW5kp0BtvAp79UmdkutYOMfclrXBgfEwzrWhEglIxBwF
4P5hn6bX74cWeq75iNsKoOhzi7PvpisR0uSGwVyKgQnLmi+YBXcx6eggctpX
J0CiW6I8nOkaoBjaS37HLlOro/06myiVrzpi5YZzj7RmHhx9JwKow15yJIjf
X8zXHQA9PWERnkzS4FeVFkzhwiivut2mRm5aIaYpyOqpr9x93Sr4TgUEM1ca
8p38CQvsLk4BkjTpMzyGY1CGE3ga9XE6gUGE+hnVjyyOYVJO7TG0ansgFqIH
zNbzzSFQGbEp6muFAUjco8htsExbjI6+E5KWcRZA3PoXfjDxTLxhw+KTTAhz
3VOOoiCY6hX5SDokYENN6czeGYJwo2S+57EYgzwjhP+yDrZPAF6dIGVVkyPN
y5G8N2pISAirFQ0n5Jvfl3pHpM/PXe2ZSXSZ9UmoTu54xRP20p4eON+IHuY4
FgO098lC5I8av8JVT2mq4VN7n0Q9DOLGjvqQVZYYn0dneW4916pwWlnfDB6S
JWtXdnhu2h5lkAE3rMZYTMYzYDxksQzOutXcCLH7UBMeHlSlQHK/zF4s/MAu
5PHF+9v2YbGOVxD2sB7XzdcdqFevdO3O0wct5Sz5ARtxXcBpSYwhIhMrQb8S
G41I3oAFkrPmYWevUTtnW4s25kpWM2KQXiOu9psfqjv2Rgt+1YizAzL3LsR1
bdP1DCOkwrjsMnEwwVRAhBTBK6DyM2BAqm0dz7Z2ZqV/5oHt1lsVp60kk9bi
ty/GdHyEQw8U2YScdYqelQ3VnXjVWjKIxNerYb7Mq81z+vkzBZPDcf+my+LM
WfZKnddELdn1WDlbu+jKSjckrVB5wIJyA7vM6nh5B33k33e1qbZfjHLndvFL
Q/bmYwJw2X02k1KHKuRc3JSPoMyJV6xwbRtpYN1uf9OqLgJpteoKORnpWDu+
QcykRE+PPBvI1wRbf3/TyLvHrkAQ1tHgFI4ASxsqB06PDGIjdfQZOM7LI9Is
Adkmy31NmVnR4iYbtx3gLW6tpnEUBa99+9qzfcB0oHpwFCZl//5xu7C3qhzp
gSMg/G5CsIzDwOZKIPWzVH7yRImOOQAGdcN+Nd+/rj26QRYrve7RNi107JfE
KI4ZdITrnDqlGD4v2Dxh1IaUZs5XqyrkvCKcg7eugewSsJYAMHguEY2/gL3C
i9yAi2In1KKrT8Qx7fuGzlhcG/C5uZElIq0m93h7IwZgL/Un/CKn2rm2iyHr
cCPw9nj8qRVMCvZmaGhfzyk3KpNlou2heypT8JYtYALstTbwkrR+A+Rw5tbk
cJl3gTGbRR8vnPW5T92K5AZ1sllIiPclFWvz8He5dt0BCE60HYgCTarWbahY
Br6Uhsf8W7tNMMt/aqFSjUmfCoMBfQ9wZMollu/oOIFbYD0yQESdvr8q5CJa
Bkq2MrT0IUlF+Ob0RrJmoRLfSOwIrE6kDEXafXmzCKdUekZdHDfUbnVXuYBg
2OI2ZP3SrAzG8qxzgnxDziIiMjyi5Lk2qZefoWeWlMji6Vegt4go4MJm8t4t
lu632DzFfvxdjBkw7AvHtwucZUsfBh2V68TlhKDhjKxYNabIHwkVTjN9YLy8
5LWnFfo7faokSVmIAoZhIYvQtLJZIocesO32ORi2NX6I7SuO62D9Jd7vJ94y
pz5UGgmW82RYPf9ryUY+YQaSX6l52aaCxC0keSQtB5tb8GOMik02nfb/ZkL5
PIyR/j6Wiyemup0QB7Ra7CPuXJT5XLo6hblN76yE+a50l9rJKLAGZdgoclkc
RmBr0DkQ9RtsuBvQkFLAyAmerQOFMJgt0+eHdK36LKdNg8ZUmtFyBhJfdS5J
bmMM9r4nBLavEumIeRMmlB8gr7ccCTKjcROvgGleqWo+1PPAiEd27ajPVPg/
JqA5nqCx0smhUHSNSZ7yIxUhLtKF0IVIRfxJfIxdKLOesyClQ8sIRMYbatA7
ENKa5JP48gD+GL6ZBSXCVwBTeCv61cUgKnkiL3nq/Tjy5v6RXC5/5FLXfHNe
NgtDGV3d4LoHrfQWY1ftavZ5yqug2UfBjh97I6xwQXYWZ4IJ0B4gOknVjzlX
59Vmuvf7XFXTqvJY6Eq1VpfDem5hxLWN9TG8cZ0Fop/kOHhcto7MQ2OE0X/o
qT7zIK+CYuhQPBMcWPCZ0I6dCpmjTn6LO9r8Gbo1vNDUhOHATwsnXxKn/l3i
KDJJKIm9/QSb/DISB1tushrG5Tlp03VW9yvQ2hgdAHVJO/2LdHcmw9Hh+jF6
35fdI4LItV7pPsxnACZIB4qTuObz5acpE3x6msBLYcR6ASnOpDLGzreFEK6b
ykQpYFHuGe8dfqxdZCT7fjU8adW6r3aESHRROt1MGATvhFGYTqDVwWXDkoNm
5aFA9XXvjAR05pHYq5vUfA0SBhGt8J4H3UoDrAwJ5EeWk0WnM81huGfo7xPN
+WIf9sPIYTW+19/MAbzvbp0RMBgn1BK8w/njHVLvQwDZGjtOjisVV3iLat65
ByTpWWSw7uVi2pYrisrkFh4MnUz/fc3AHJgFfxXZr8sxosMo+Rnf2b3xc6hD
RoxcoeDirsJEmxvT8GNdPYvZgFvboXvRJk3RwaD8cqbw7pcAGtkYnWduLU5U
mtIXLsLTOepEhMcMQsSi1N2y22PXlo/wf5XfHSHCyiI51twKSdl//cO/+u1u
syaGcyWb5r9EcN8E0IFz81Une3bP7y7uDnLLtHYlNUuWOvKMMRFC/8YjGUJM
k/7rp9AXbOZJnDRvJXRcl+sfR2PGQmWKfVrwXl+/jetcl1cVuibQdYpMweun
jgTknOR3MkARxAoQPDpHrDJbpeqVqY2hwJKirI1aL8ZSIxz18fZHz0oDc0vi
VW9WiXug6NGl4QyTJSvgSzBGpAKBhqg6LqGVR/dtFD8NnfPRGF8MXtQiYwDA
QoqrH42pfbnS/gLk7UklLGOEPg2rG1Q9Jod8SPundD5bmeTeyBQmooHhcHir
J763aV4goYH6kRlKdejs2muaY9AD/rrlCela5DRsdL0hC0T1jcz76SBLWV5y
OhKm9RnU6B21yMBGodRfMh5gEReIvu8yWiC1QK22ktAxeLTQ8uSWIFHNw1hg
rOx0DIKIk5W75yGtyc+EMLKxFRFos+fxzr2hBHWNtpnAY/jra5ewCHdMj3FC
UE52/qdmorI1uhwBaf1VNCTyZNPtcnIvxBy1xkGdVnEsvQRDS/s1JO0T0UbW
N6jWr03C10K+TfrhwRdv7GA/tnaSe2xDTwXWXx9kOKHjnSoxZEOElaD5pILQ
LN4MfVjOwnkwDd/CIRFkQrI+1zWixLIlOAIxlyT7w+FXQaqljTgsSLv7azmL
6PawD+BheX5gTGMSlsCx/CtjfYbtzdqvUVfsNHNCB4xUSyBHFjcl3zjNvNvH
NoL7MykZPTTfIJANLmK520l4eR9ZF7UYQiPctCGQKgG43rsQVApZ89zvQTrc
1t1wux1RBV00fsQYcaLtU0QI67/kzu5mcdlO2UOBQuehuX1f68USSfjSpLsp
4k0shkrF9szwE58GWAUGhHhGGmbRnL3/F7HSjuDCjbuf5p/iaWluhXEr/ZJI
Aa7rVTjny1P7JT2a4z8+Cce9KKVhVGY81QSHParfJ5rcVU7W/n7TThduSZxL
1fGQNzDGBio0i97Yugpkc6sJj+3CDnu4EZDSPFkbrULliPj3IJd66DQPE8RP
T1mRHvu5I+JHb9eS+MQzPHjShWhS1kiC1+xMpZKOVzHg/iauec9cdHk4JX8j
1B3VeZ2k4cNq0kEYikYzNASenEECUSIJ4Mhq9d1a1RPMhnXJUmppVNzUWG6c
KJlJNmOCAOY+Ji6OLaO40857P0fnfJJWDyqUjZn1eqaYocGADscwXBe89JgX
dXp1/wWAsZl9iB2cClUTI5FjeWBBbjx4XjPjI0w71K4nOfhNojO43sg2V2sN
5sTxU+PLEYmHWQJZAVCixtxVUC3FUrLut3aROUMX/3zAiT76J3MQbXkuT5LF
ZIcbk5iP8vSSDefhvxQJAvTfHcr9x+R6y9614bSHs9FtEMKu8FN8boQuBc/n
pYFiZM686gxunSEzqbFsD/9j5d6MN7/A0oer9o9Y5mKe50FcU337sSN8fcju
n/ZG5By/GiQ5QZ/mpDdzMoqdufqjs2p2C4v7h7qlt3mHp6To6ZuNg0taQoaC
DvYLaAfv+tnOhzo4OGADZqMqJJLqg61s7RmPhxUJwmAwo3CuutjczuzwyPFy
uPrbGTG/Ne9Iois6mvf3P3xnCbrEC4KyX18/MU34mJEVYKvIb1PeKPFsgZIx
cCYQeVn278wRgsYHurPKhI/F83ikH63qsQ9hbX+iVqu9baFmjnwuIBdMApOP
d1J1DyOWGtoLnxBIAMpgzbwUO3Adb5pN5332lgPTdV6kNyNEULnOPGmFaXVE
YG1Stui5MxVgzW6gIyOTRXqaIaZM1hZ2GN3BMCm4cZIMytZPpBUtbjiFgdLN
V9iqEsxzuMhQ69UucI0bnKn/G2MAeMSz7+FG81VkwO+Ya9CErwceruVAu8gw
PKIOTOMZlPO2rNgET5kp9UMSc4CUQzcEjD0JoLB/xXR/poqc6wq5ReKb2Dcq
IIUV7RFLqRPM046aG6Y/ohtmX5i4NQ9KFx1xedh4E2tfRpzJ2fP9ENxKAEvM
1VwZY+Pd3TCwnGqW0YkY4fxPmlTWvZCluEGlkVjOeMxd/YvRi4EJBF8Bnwvc
fOEM0z+vUbEa0cGDv/MI/bZQJxCm7zu4Ap1L7bfxxrEN3As+OhRnOQ7vq1LQ
k8q89c0ivZOVxm/G8EVl8VYJ1TXcAQ4WJqusNLk/ACqgoTBTyn1xnAkSjQ1n
BAonuBETcL0J9ghsbwliwjTBhnPtLiAs+x70p3rLtq/32UbieOz9exUSDZUJ
UPWmqsUcdOkR4o2oM2yQt+/4wrqRVXyfXJS9YC/jSQGNOkw1/8NCTpztKEkO
bJsFe4itIa3xrmakryYSlioK2MB1Eu+n7kboqDR1dhIt8jZl+zwHzW/L982h
pJkHsN+cA1OKVh8+im/Kmz5jrEga8r1aAT1eQg9WuEvQXqD+0UJ352xmoW8D
B0puZYqB5liqsLCoE4RGjchKuMJrqrKs7R/JgIosflmPKupXeAmh01dK4JBm
n/NUomRCf5a7xyBVC9I2wOxlsY7xGWBZAIBqCL+cqAZvWphGEOgf9SOhknhD
/WLv4+aPKKD1R6nhF+FnecDLVf9FHo4SiPG4JPSCqBu6KdI6DdxW1EN+DUUC
371XBQ1ZWpyb4tDVbDgNjya+vTp6SwJRqVMSZ+sOvZtewjFNv9miWeeiJRA8
Maj2LFbScZuQtRcgRD0Y0GUc50TB20n+T7lVMVbf5h2BH0e/uYlIHf0+kMQ4
1dfi2AYrBNxZsBpCejrGVZQ5STFIA4ty9kBfTgn/UvRmpDBMfV7H2oMMV4ui
nWwyoLHZCsMyec119MUVEBhWfvNeJIsUbBMkwfAF5taCNm+k8hJWOKFuNKjt
XoqRDw0P4LYfjXuJ9sbkJtTCSHvIwW1LCgiW+s6ZMhiIdcaIumIezoCzQdBG
7H/wTYRr05D+FYTLK6M/aVs9GZn9gGjuUSy0iUrpV1GGXakPna5mR2VQC7rE
VXspkB/uaahhqDm04ILu9mK/lnPagVypoyV04O61PwNrwjxYu238QkfILATt
TEWaN7GBu+eBBcwN3vEuKQjp5ZB7lia3/bok2Lu3Ww/FH2M5FvmAZnDHPwi8
reiL4HImAdv68XwEDWvdfWDbILVI1cwtsEUeM+mgVvwa9Y9XbIr+7PzysYOB
gLq3HUb8A0YxhE8R72ReT1GSH23zV6R9n9k8MYGk4E/fQROAtC9Z87ZwwOhR
fZfsXhm+BB6Ezm8ABYvY2ygJk5adt9P9XomV7TAYfgv+9BL+nlsBeMQ7zUoL
oXNHqwHkOUOtRdxkDxV6RUCSLAaqZDogMnXj2+cOIG8tZYa2Cj9UUw7NnBWP
2Sg/1R2b6PfQyufaUt37bAULBkcsWHiWZP8IC77PaAH7kIAQObRKtr9yEXHD
zUS6JLbHB7t2pcTUQ/5BMW1Ws1Hd314JCISrrqMHj/tQPSVDRqxwHTw7h5OC
uoGvQJ4Ud0AyjSSS5SgmuNDiMpFMQdZOit/ehhI+cnk2OFucbGpRIxnmtllL
LevSsLfcc9Fy1sBRUyKiiNJcKfCKgmniWT8ERFW+Y3+3rtRFxXiqjqt8yrYh
zi4iLk0/zjvKsRzsQ/KyWDpJDAH4sdhX1xqTNXTvqi0lNLuxhkctmylZJXcv
4ci3DNaSDQOTdJ0btHFOv5eHjATmUQRDxUNhKSCyImjXgiBZ8xKpdItpKRCW
aPndVIUYSRs6IW4+5RUs4h+H4kmrrO5CyEM/O89oCgPr+uBcytPzReqn1la5
xJcQlATBURcQ/IQn8JZq1HzHwi+Vo+rlmtd3bICco+GbIlgrqItMVuv8Wzh/
K2GxMrp5OwtOMwlFCikMcRB5Aduy4IUMN2nizajZ4FE45vemZLLEGOzs9HGD
Qevo42QOtBIzXKO7ErZtg9Z+O4PjVxseuXjKnNfe4hO8AnYdy4IJZxl7cBH3
NogNN/cVk46pL92TBN5RNQZrGzsxf64Va8NHcxuKctmvgqS1poZbILXLHcqM
23xQSr673N/AeBAOISbBEMAuGwPWooRYzgzG2td+t15fiGpFAhYqIPX9dCNP
HDHT0Po6quLtQkhvsgEuIPg41J+VKkaBbPczzPA85Sk06o1hKVMqHExwVmfn
EhuU9BFodbTUfdeb+hVObO/DdfAX/Bj5MVH75kPLOjF07UO4wSD344LiWPTh
dZkPplXblAZco15sKLJiMji1L86hk0v/4C5orMC0PJmapvfuFkmfKpYiHFjT
/KUb8W59st/L7mNz1RYfG0XU/ECsAb4CV6khkGB2uDWwtCeBvA1ieA3O6YzE
/Q+NYT1kfbay9vv7vVw/EWXDsAAj5gljlgQ+OiBZUfgou2V+HNhbmxUnSrHJ
0F5m23cgyW1872v8N2GKJlOJFATUHKXZht+9jD786BBieS1huybL1Xz/VfBL
QbVUmA2CpSIWtgI/yEJX1Njxn8xFRCIEC97Mu4ljbfzxHsbEpWCu4xam59Zx
wcgCgBycspxDhsLvHDntY3TAS4WnmKhjvIsYXXEfpyCXCUz19DBcUmrKqvxO
hETeXym/H1uKR4q9ZNA9nxLBjd85kmBt7JNlzCje6SSp4CEA6+eIZgvazrWG
HmFf3xfMXff0km4tbOPxTLwk67O/74Pt+w7LY5Ye83xn1aAgknvZ5tlfLQcV
aSEPWK3fIp+c5NfhBORnumtYus/mUUKcLLdWd/bjj8yJCG1OrCe0LvWj4qbK
tswl8w2EnhcZ6TguATPUFCR39Su4DKpsCJzi5VkAg96fNcjT1cqRw3CFLiy3
62CEkJebzSqUlVwIt92SGz5aW7oIj9T1mx2z4vH+HBTcV2KwY9WVGARx1ZEw
kWGZpyNjeKseVdBiBHu8vgNOV0mntpArH+Ho0l7mgHHTGCNp2H+CPptVrvfy
hUovIkR9pYVj4+KaZymubpPC90XT/zBfhpYiQyIdU3D3HUpJPoWfkTt5yITe
w3AkVwxKDr0VEdhatlWCt0Xp2yrzDI8/NZlSfON7EJZtpC9Hln6QLceDXdMc
SSHkzjNCm+7rnDWwUFBqv9yZt0U/AGMICE1QsX0O0a4HbbKtE88CGo3ELjGX
icR1/6oTGj6hKRrDtV1MMT6cxRH2ycJOjPRWYGkZ0z7MLk8Rg+N1KelHcGm7
s4NPjihc74tBr2XL2MsPtqL1kcCMjVz7lTbJwwNStviiPFV6EAfxpHEY5Liw
84bg3ouNIrvhjV4TvP/Eez6Fd4gsGc/+YToxcii4wPYQohMs3AjvxsxzVSci
Y3T5uVXjPNk/LtuceTXHQO7feD6EZAaZYtVOEfDZq4RlW6T6q3jXqUIUmrOy
PnpAA+/4qs76HYSlKLSRMMCKuIS0c7Wghx9cI/TBph70j4lBezbtrKeCGZKZ
czkns2LTbGAeVsi0w3ePSiB9zsZOTSQthKq6XaVW3CnxQbFI66I3fc954dza
cKNWNPxOL+fGEAJCD2V5NOAFReLsqcugeaZF7X9KyWxOzd5CFmKE0SbHGKke
Q+aZYjWVKY1ejj24CG2eSaxhM4iv4uzfjTp6uj6TG3iPpogxm40etv4ZFOvi
xUZZg5wjMK/RV3vU1DS94d3vIlC+nbsyYS5tQlZCQvjv7J6AYPWTlh/1qWgj
Vdk/YR5h1kZtJjAnj/2ke3mn5s8c7FRO/jXEknQ85UimKqYitN6BgF/omRiZ
nD5Ce/orE28npoM2rGe4AcZlSh6ijngXaT3NRYlW5yJ7Tc6wDqlM0KtYjZlV
79M+lvjfz38XBIWeKAV6le8RYfq7+3wsKgmnsZfLF1oGcbg5CAUaJsMT7Byq
aan/+Fj24tGdSjs21vz7S3K12YC+eHEqrTnMys/2+IxDBIdGVRgPebF5eCj1
CGA4jCaXCyGlqcnMgFd9g416yVr8AUXsd7sqdDBW7OutV/XLouevJWyrCper
8IT+NlDDutJ5oJh+wf1Dh54u4N/5mbLKUhZDMVbyhB7sW8F+1gkQKKYr0iLN
Ax3x8qdClUAkN5vmA4wKJPcFLoC+ooUOqggThc/FPv/vyp5EFaKdN9zxc/dW
CwXoV2cwzDO2QaDHACKexbOpBuq4BlQ7FEDZU+RPoajPbiIFzgLzJwKnc0GW
wQcid62JF5YQbYfGwb4Ko5gh7shkbKKy5DgjOBUL1DJluIIzMcriP+EQ9CGL
gCvimxZFvonJQXrJOngSWHhkpspwRyLx+EHT8aoGb5mrnGaoBk0xJesoGRGy
7iZNOFm9LyUAlIj8fzsJPsn/u5XbwACW9cSziUJU2/86EiiS3RcDqmdnlzpS
KYH5l0aAB7NDVB0YP7DzZhwTiocD9WasiXSAO0m5hAXnknKPfho2HCMWXgKg
vkYJ9gyP4yWQIGAZ+wzcKmsjxqEWc/6wjopLC3Lf8AyA+V42bxU2GRO86EPt
yKtD2RpFMFO+Iu6HVKE9Rao/7rDn40UfWlq6lWvZE8kSZq6Sc0HTaYjwmwsY
p5DI+WOTVVvLUXIvtBQXYcJyj8tV/XVvKZjqOQG81BAkRt8OB+FmPs5laZyQ
Ez5BpFMHhxXG13I+yATAcfaZADaEn6XClUkIOfrgNHAe+8XnzQwRQB14GZ9M
82VhqiMprLc0bO0v2YoebFKZl4BlG39SSC3kJc0XK1ZNEuSO3VIfp8+sVw26
YufJ+83hjKD/6zOwQogu25CbUfClh/ClF+m1Ml7qX4t/Uk7/2EAL8Nz+D3ei
NjqKZz5hNkona4MYi1Ohabm0hM2h8D29xD6is+l5HgUjE/fpoyc6T+5KVxp0
6q6BkQAoW9IsyM7RinjPZwu3NeiHMC4S3TTOHGwBrF13X2ptLYJ/PgeTBlTl
TpbPYPxB3BMSZ90UdQ1MbqekhDhV5+IcrkDf4iTECSk/Og20g+plPj6ovQs4
fBI4YgDGEfM+DCJ+L+TITu95DGygPemxP/xoTo8soqS32KsgW3QRXWXk2ZbC
+fN+L/Px0X6EfiXTKRGk42usKXPUGjqnSbzjzGRdLfdw9McETBMoFu/0Sxq9
Zg6WL4pJcCk/i7zfn9cLhjpz/gVDVSp9botqPQS0EGvtYDovY1aaOzXF8oH/
qxi7cLg/o9tsIOm+AxhW97pAiTTmIoUcldqKlQFSQBp/xiN4cv13/MdLCzYA
HFPTR5vVkP4QFckB0WFVfJ+Xcwes8E+zx1IamSiunYbHdXCCYXbj6yOQQr5u
KH32k2LHGob9plYzg7ozuf4+ie45DRIWMuEEt8GlsHdksmEc2X+eJr9IsKGW
EzDt8XWNcZaJf55LPLvEVLjSDcqeypa7O1lY+7nNpl+kKO8NxEY91NolHVjb
yvDhl4o4V3v7NjMNFqO2U5XPHtNBGbGZJpxJsP/wqsGjreQ7Ur0BSxLGVpeO
+v0NA6LbnkCTc5kM4fV2Q4QA/o7tNkt4g/Wux2FI2u6HlWqxVwYY4eh6q+zx
Ja3c9yscu97pJadB6o0S2kt8FARAChOlytT+RYMhPldqT25wYBw1QY2MtI1Z
pioFoNo4DhYP0QjUTtuGYa7soynRm0XCm+goVkGoAcsFKCJVCCFBhzJDjD4u
LlbBxg27GZaU6b36iEqULc5IrWlKe94Hz41jw+uwEtscFwK3e6doVIKwdryv
X9WHzLAw1VOgYxQ1uu5/5WQLM5799womJyXENEWvPbe0xf4hxtCMHv2aJjlu
8Myqifr2KddlgYZ7xe2XwvoMqrlSrFndWcvc+VFnnHSUUCBuA4JTEhyeJfkf
Vb9qK4Wpfz6OeJdq05fT4WI9OMej01cDDMYY2Kj+EQOZyJ7QpaF5PmRhG4j/
U2knzo4NOTZRQDWmUVr9Q2SS2glQFiBAgDxIuJjSKcJ69Oab/uhy0DBJBgOn
tWnPocJYrTHncNUO+TQ4nXj7YhqOBe17DgjCoT/0fECW0X+BxtILej1xP/aG
ZFje8168Z4aDnVZa9Gl2Tq02b1jvmGmUmizn5UwGzJeM8Lwrd2/QtcE8/KHg
qM7P1PE7pE0bOHReiz7aibmr3zLZx72jdEy+SVID+/N85JsYvLBRWGNuvRss
siXHDva3U0Cff6xaDlDxJ7rI3VT9YI8O/GUhdYNyJil4W6S0Tb0mKtE3QmNQ
EIAxYCUPAxUcE6jlhB8gemB5lDyDYBuPPRE3620Cu3Ct4b5TQNI0YdnlpWYf
M0Cuyrjj80CMTpJKzaSNt9UFJH1x6nuVROGp6UgkQRKPT5ewTOSY+avZ6YAA
rundooO/gTsuXOTNgwvu11MPySpkjJQZpceKCmAP2WxGqPdlpEwZZhPcY04h
svNjljbmGCW7BNx5M1AHAdmofDIYZBm+Ro22zWrl+64WCTcjaWBpL1PXEb2E
sKLM9+6NZ9d7D5csyTcKy6e1r4o9NXOV15OQjlJr3HlNuiIbSaUPvCDsC0s5
buYVGGdvG7vYuZN1XjkeCDMWB43h89/jwq4t0vs30wClyxUg/yyPlZ/nYqge
fEIlFIQbSXdbaEjQoKrNLZTMCUdeicP9Mpn/MLBoZ/cqfkK8pmnHofWv7QE5
x+XD8UIJM4Q27BNCQV92GDb543JrPKtxZRGlOkMsF8zQL6+5GGOJYZu1ii+y
XmlO5tjiMGLDTSiYGYLsGdY0NFvESy+7w/mbv1nFWoncIrJz6/H4Bj+mawhB
BMIRddDl8P7X+g3J9aFOaBCumTffXRQeDPjjeixrTYyckfZnZ6eZQpcEZ2Fv
CvFfvX3U01fhwl3oVTYfD9Rmd+H57dE/kdGiLDBBLszRHJwzp3EwXdyMdb6B
81ue7V4Sk/Te/SshoKTo59CEysdE4DiRj+OPhNOvk2lXYWiuOcGOj9d6wpfi
8B6SUBx5t9jh9ZYOS3aiTt8GANruUmu5NgiAyob+tUvDTA8Jk06qK/CdExdR
2vbBeca/9iBmrj3ACeF66e674Ur6V9y0zEbFIejfofStjNg5VSonoLavJvV1
pw/dIi4mjSKAkIgrKkmloB1HObI5R1B7XqzGZGqmm0fJstK43HvNKqDQrh24
2rbSLimH0CB7riMyJjCHGNxEe0yFIEbPttUgXhvEkTv6NytXtEoSlz/ro5EZ
I6jRdBd3pW4+O9H500+kcYOhV+OWU2HBvfPRFp/uHaP7tqV4w2+BaYpRF4Ug
RQmvCtfD+R5cKGa04my/vTHDj/ukVNGk3+WIIStq5pbCXaW26r/o8434lXhC
HmhhqtV+aLHQJwKFBEru266HTXFsZuHmZ8j870qaqnsQVzEm3Hyc7X5Selrj
h84p1kpYc22YIRRzsiNuUOvmEiP8rPtU8BGRkekvHWW0PWhwOX4+zAmY1W0v
DYnGlIgxZDNVgQapZjUbslrg9He+/gKfO0JdWx0MwkDzJTFxqim8NoxwC0gz
qNtjiN6W2oDm7CXbpakfHuwaT9iEv+vs2+jkDLylyNcUgKFxoskdaX70QOnV
Axq8uTzUtFugNAO02k0Q3EweCt81maEzwbV6Coo/Hrnzii+ctRxOe487vp3v
FMPM6AF6fJMVsQIs8k7/y0NfCs4yd6wRe1iif7RmYZUbY7eBDk0oaKdw/KlF
oCqoA3gHbKbWPylW7J68fqBYGRAqvlIjDI0T/Aygvyqa6Y7fw5Vexr0yjpOP
TDpC3ncHGeKXVvcl6VUVVen3HjkZ+2YGq1epdozPb68+djUxBv07Ftm2KsDQ
ocrog6NUmA7i+Y8m0+BHvEcplbWAWQvWOpUu8WbgLWCYf0i8WEIjKCZOkeCg
SWsitKHT+jAG8Cozm8ZpzHfMCm/ylgfVb0jbfzsglMqpOiZ56jOKRUV9uFur
TJ5CoQ4ToC4vM84VIL5Q8ujoiWMHAvpnupOs9+XMJM6C7RqfRK8Se/d+IT2j
YRDYqtOKDxAVLZrCi+Uu1ZXcxOCC9i767UJkEgC2e+OAYVtVz9vBcKqc94Y+
fSqEq5Ra4PSVPVCbZEQYplO0dAPHKkzelfWmgInUFdeQugkhEh7+CxhVrzx1
QM+lwQ01jXAZN3fvNUgNjdRijqy7ZFWkYLei/W4fGc63iUDGhsuu02TJf8wI
xfb8zOvUgxMx3IZZWyDWK8/hLflSYA5BS9EJA3DV/loZCOQ5cMaFFi0BEvWz
KUrL5AAuMCnW+eqsnzdeanSuPKdTaAjZrWK5I75e4HhABJFMuCd29HBC7Sbg
HQUv7dYRpP1/aECSqevlptx5xJUgj52e14z1tRCGwfy+AspfTaYmm5BQcVG4
T1tmVKyJQbMa1B03SZxGEkZ1g3oPHj/boHRlrk1PR8mtXRsh3fQXHJIJf/Od
9d6eHpsgy2tSgP0nYiYeZ1CQXJ+24elFT7BH6ONKjAqZgRr38Vqg72PtqEIq
dF6q3Oc9eC3zqs44weoTx3bUsD2ULrXuetue1qWr3KcPHS2Ga8yVLySJaM5z
PjcMjg4itQd89ge5elvNVNkvno47LH9qoCOjH0fBFOBvnd2U1XNPY6aXUNyH
ADDuU59L0dySnxeF44Iviu9zBuBZAA0S7oy0VLZ+zUK7pfSDOuuG6jjqWI5M
lIsuZPByef3wC6JaZUaptE0hIekbt+l0lTssl0WZqJl6/CovmzrAWwrD+zKD
VGn4bdjHYAG0Od2Rauh0Nq05YGJU9IRwkbiUD4DQb01+RhtK6PKC6KktcmTf
R1ukcpTzz29m/co1FslnVfqM6eQs7o+yyfAjNtch4tFaGaQUWa2rX2yk9LTd
D6CQYk8NkIZ/sFn11Mic77S5gQnuGuwqB7wAUjoRFGZKmev0Whleu5asLeE2
9kS37o5xH4c8zGEiqqKef6qnKXhBAp8Dn8vigMx9hQwYfaV8Z0F8/sx1Cvq3
2+8n6kHRy07wyB0ZDgv0PtWBF8uEL5r6jJtXJxBnj25YPf5Lhdb8RBbnYZAb
a6xTQD6ymw71OQd8bGjcFzB4Gnn1FBKZIN9t6lirSg4GNzkqliUSQ7rMhGqy
w7v2u2fc4WIaWZPB/uRpbAl32lueGlRVihmAvZuLrez2kX1GxAVKutOgd01d
HIc2MSEMMPDMi8ASxCZhOd/jouPp9yFFkTqrToCZF8up1Quvfjkahkv34VYz
QksnyFCGd6qp1ZTEfHR9jeui3d18l+iIKPzQgBD4KdeoNHxfdtGQRnqChYbf
PSKKW3JpwjmVSjK/75m2G78Dyx1A9JkFm0fPyzaH+pZ0LMc9AGSwIGuMc9SA
nWXW702xkZvW05eyB3q4y2a7xZDRtKclTi6FLaGNpv7Bmi8gKWg/+y+ILoIq
JSFYmng77R1HdVEbkl31i6n6KUZXbIA9TpGywHWM/2cvEHcvCT19DP+lFr25
GcnQ6H9zy44ljN4+HbTRZYBANqxA0jLvFWF0iu1sresGY+8PKEDL9FO+4t5n
4x9q4N+MW0XJTw7s3HeBnUMzGLLK68nXl69eOxDHc29iQg1MXT+n93KTYyhQ
v0OQur+ysbMKtFqhm6KmBy9fT3C6pvQv4yE0XMMJwvG/+E47Xo5GywHhLmWw
tvJLN5D2ssGjbe2FMnO86ARjSaWbgm3xbxhz1SJYwmiOwQvB30zQtp9KdxQb
ObomYYs0bW0m5unfUdVKKkXBYp8iI9a7hVmB5ugDHlfKUkS6jAkQBRys9pLs
xD7D4uUQ2o9j13Wge/35GIPwMPqmvB2ep631dr+KX6W56lwzNlCribvDCrCh
GHBTRqc/+oXuuz4Z3JJFsXeGKVl+U7Sogb6Z3CdlF8Xbya21SxI0KurkFRYm
6XPGNG1oRKsnO2jEByjrYSVfKWR2NiPku78Y2MHBCshUaKSFnkHLKBevGMdi
HPXP3JyCf5r1JJd0WyHP8IoHTBwoAI34haJXsF5/C0HocWhlEVvU/wuya01V
YcqrZ8c3YwhgI9WVFBe3xrh3aY5jXlt0dNtr+ulYQQvZ8lpfdpAMS0rmEp2U
h6PQ9IxTe/UpDLXcriR2TqDUppsqnO42zSJ4WxoRpJ7J3OYYF05RfMqdeoQ5
OJF8AO3Bxb0FUKqinPRCdA52COwsXnhnz84325UBzKHVPkJj7rJ4nm70cgIi
359zaVK4iHNGnofK3bon1UIVKsdLYqm6s9GL2tO99gWWoO4OzvJbdAE3QJfd
VddoRr1zho+88Njv8LITmMsmt194llD8GJ7bJ8wwjFzWN5NJfnEKlp3Z7B9Y
n9fkBszncQVCLAB8gj6OTvz1n/CpxrSXrY3B2Wye2kNtxmf02ZpRyKJJHeQG
IsPir+X8iz6CkpENTgSiNq2uJ3ZoevmpsVnA4WeEVDfTB2HqSVc1KcuAkWNY
SzYsRj2s4L9axHM4Oj+21pB/G7u9fkISX9nEhERp+ngmM2EH/PuVdj7H3lyc
pCv6dHXZEFwJuqXbGvw0z+27UmnVhtM/uDCeGfUz5mFeaVxe9QoS4MoTrgj9
/9dVWOd4rwRqAC4q4AvAKagQ/rFreB5bckYEklPYoiUa3nbrPc6AbYicj1Pi
NDY/4uRXQ1jB4OAQ2uxnG21rx+AZsvlFScvVUY2RdugLHBoDWsxQueFMOCqp
AVKuv7wQ70DOp+BWgyf3DEvtsa/TxDeGTofOlDL8MhxwKeSsDjOI14argQuI
3reopiwC0FuyvZYJFUpXxk3rLJcfRgorUFy0CYfqdnujBOQEtESOsSb24bVP
xdNDiqGj8gF6t4Yn5g3Pxv69rGmyxh2Rx5Qvyl2Nazo1p3CL8TJBIJhTlj+l
ZVkm/P3mbywX82l7s67wkWcNbNAYzmbZP6GdzrK7ZKWHnXPduqMt2iHIsnRb
EDFD68Qm7C+V374vJWdWPB049t9MtjsBPzwrK6Y5fkImwrycv2oaxhr/2Vab
ArDp+P0RY2UYI+yRhpf2M7liU2maRviOpu4OvjJsMYTR6KGj53uk25Vm4lA+
fSkUND3dTM5Hv8uBr3e1rZRfSWj9ep33dtJ0K6e+W2WZEywqO1mKcMpyJmrt
gAuzV7rM9nNMmcDgLyodkLurJKK4EdnLPRblOTMBKqDDm6tGoVby7bi2Ebl8
Fz3M/G0UQTwLad/fMUKi4CVj/RuD82Ix0oWBkLZxnpS/CIU+H+sYE2F3i49t
eDlQ75snPNEm9f1q232HKPV/H4FQkiCQMSTD8NNua/Al3KThWLqZH18l/ger
ZKvaAB86ytnC6krlEZ8K+P5mc3WrDh25tFObJLwzgZ1xqvggp0RNMuN86Lf2
V2JOWICqnrkzRnbxX5U9a5IGXSgngWB7u0Wo83e8XGsdEjhtMdcOBMZHg6g8
t/eGs0i4Id4h768jOJ3wj0FUy3FubJL2tQtHanNVwE+cf28TkO+I5MvPtFxZ
qKBjEiPnhmkIPmrnrPmg8jnJaAYFNnQjNhKGC1rt4UBZHKfWm7QEKI5W0HUl
FpGb6OEC94619B7/ZJ+HJ8C9YQr793VUH/ezfDrXz50493lVrecvVd4cLw7O
9QQrcbfdj5hsA7eJo1Ii8/6LdsUcgp1TJn+xAZSb3cKGJKB8NyOAYK4992aw
PeHHfUw1q+DKA6YjzMssvC6iih6ftLVsG7CgHHbGNIS2juIEHC9qn66huIDV
cf09qI1JuOrxaQ30GZehwSawEKK5bT7hp+hMQDiR/4UO24gVERvdWG1XvIQx
i0kmtgkqKhU+fXGR0DGxUbl+Fqb/WLhEC29Awmj3ZTeGs2VWqBF0WYtxfWiW
hPrkWQdVU79m3iJmERmQzNj83WQ/uqvet/88WMAWiFyfuI+DeeyAAWJJuntO
hoMuyPh2tvH8odajgW5esP38p7WYjK2Hhz4Mnp5TT5rFbot45ksayEIWxdts
hGMt6Rfe/2k+R3tkvfWHdULZFgxVc+eEKokP+IKr7GQ8lZitJR7dVjVMCAqN
S6cDJkN9EHtM7BU99RvjgKf1QijUX+nwsYkJJ1XzFsnwewnPuFtDskSDTDrX
NzpKjFgHtDdrd+V508VZL+chW1SBAoWyuKwoMEWCKRhuzL5JUeTRbQueTYuK
sR5q7oBXW1Oqznk88S9uhcRwuazFpQgHMuK5sjnQyO2W110HtJ/RiORwTzet
zAzP96mqWfDeKoxBmMCINN+K778Ahh8SdkO01G3G+bvqKzHhX86qSAkB+PHr
ljqcpYFzAYzXcgWJEk9Su3rZKbBkcHsB1sZrhtM8bAwmZnBgykIMDjOZNFHv
netKhzug5y5ZmzBJdttNuJqbrW5ousPIJAaX+nwHEPF1CYSqPly/04Ea0+/k
Zj2IQm9C9r3ll69T9Lg2MJtc31RQGe2p7esj2aBZSpuGB2Ftp+JslT+cjTqI
Tp+upexoDQDex06fw2h+AfMGFn59vpBuqR/vQcnCtXuotzPCWs9dLoMNIH/x
eq6AQ4U0wmfUQTgLbxLuAlEZnlXDP+/QC48NB13/Aygladn5P8oNvSqwfB24
GuWQVSYFySA+CZNYa+leUEz1e/n1IGo/UIE7LtUV/MwRFp5vQpX7JO1P+Dgi
UPzu0JAYYXs6luLpydg1QL+yW/wpYjWYnySPhUO7P9UXV9kSVlS4w7sFCIRx
NwXmfY7xka1hl4F+vgutb2s/UjFMKM2YEG62LEg/xFo/SbLf3prRo5nzIPpF
WHNz+M3SSgpfVuHfEbymHLFLMRKOgXb7b1HSLCgFSZ4/zq+9cZkI0Z3S7cyh
/GLfqyAjl7HkLUWrLaKwF+AEFQbaVD/yMc79UD4ryT8/RB2w7dMPkdPzK8jM
4FQGK4esi3eGg37pV0v2ZiFk1qOfAlg0NtgaIF8okruUzb8G2bToB1xs29T5
T37MAtkyuvB/ofpD0ald6f09EmLOTreCIP4cZOs93eZQPuoF2FkhmCBpKo0B
hzXuhO6qY5yj6fsRoZ2bpZhESNO7bNbekrlwfs+I383OvcoYLVyO7D5zRo2h
Q+dA3EXPKGT5cnN1LbAVFeQSEgNtbHBbQJFbUdr4xVT7vbZX+V3q5Ifm3eda
nRgPvuQJTu3u+ErM2VLb09Y/XqRqKZdNW7ZlrgWswRTIlFuX1yVBhRXrWMv9
Fuy4uf8CeA3lPhMXCVhfh96tZlOpTEeD5hTVkhtHu6sDBd2w6sYvZQdoyvZb
aQsdoaTcNaRbcd6ygVuDvC4Myhv6pHtWGNfkl9dxTNbiw+k=

`pragma protect end_protected
