// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
0Ifpcf0pbOTnzgISCAdbqiyVH8bC3cFH0SQO+Dfh+cq/VmGIozhCUMf9j2uRUGNq
8ITKeh+vuVl2qED2aEBGJhlmQ3KedNe0Q62RKYNHd8B9KXZp/lguhHQs5nCCPYGE
1ccmVY/cyjSRKmFD/oRvo1aZSfsrKa1f5t7XdbP+rEU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 95872 )
`pragma protect data_block
iG/2mq29mcnpiJ0Il9CFGdvhbxEK6expc7T2rN6E4d4xRZ7SnDNx8Um4G/JsiPKW
iokgH90pLElO0TJlbsHp97Oxfk9a0xOTl8w0Lk87VPvD6GRmE4I4RoxO0cZdLofZ
5s8Gy9mC6huu+V/rSS+BB23/92d04lorjA+zCj3vtmvZbluIxMZedN4Jh2dfHMPe
QqU1Ec8uMTf8x9bzPzEhUYoF2t9P5cL9XT6Ht22p1MZrs9RYFiAdcNd+SP0LxHbj
RPe2hZPUBs1Od12HZrxSog6HubQ06akRbxsAl3tqNp7lmYrXuE9GhWUW8D0cvcGK
rja41PBJQYNQf4TB5W4Ua1qV0wljJfP6nh2Wu0KZOhr2MSEA11QQB76FnXXwt+2P
ZjwDIK29ON8vaI6TF/E3+cRp48cdQvA8JC0DmnEDjdTvKIoPBCUOkfkn35b/QxpR
xPndNMnl9DUDV4Z7si4s8Ta7wvBjRs/832240eKJvDuVH+N9TnyQdMoTmvQ8+ln/
9fTKKO0Gi11HeFWsmBhxUWgWwQMI/y24gc4lT4Mg7dubgQM2FP4+s5ypz771HGPr
mL2xi7AO3nDkEpDU0IrrcgEtkxFX0PCwZuNFLLTqfE1MvtJ/x9QDRTTsftIWs3Cw
gev9RaM+46RN7jbEq/6e25c75691CwiwpFzi1uocNleoWsIAezgQny/s8LISZSYN
KjpgoeJXftcyQjEOH+SYPt4M/DWw5vX9sPCZ+EA9f+qVG8H5TbJQ7HrLRsJK6QcP
3OunEDYPBTTIBqPvG7KsX4VAWAday0x8YxlHf5EuJB2A5VPA689MjWpSZmxOiUmD
blgZ7vBmu2VaAXdH1LpGmNcOcjGcJTQinfMg4gjL0Il2PcqUXWc74GZqsEi3lmbf
7HX1WLxcNZVDpEtG1+7f6essr7CMYxckoVF3SeRf4ygZ7jOfx00SZuRSooXhfPHi
YuukqUcGc218miE8KbxxibY1SHpwnu0M862etaIvBxIZHxFfwRa6YyJeHWPwJVVv
F4k64hOUmX1BgiIwMHXDJ4/BdtiiwKc788dhz9f9IanQglTkNxk3LIgRFZLm0R0I
hgTDHrkPcRLszSb3x5eZrskYLwJpmXS5dL3Buhs7FjI0SD+a0iiL7FnhGrcJ2IsB
CQaqf4/J+YusHNi/aK712FarKDVLwHEFE93zZbu9kKgxUCXleuO7nIgj+UVHMqTG
hMUb9tQDfoNh4ys9YlkCPXrD6nLZe9SRoSjYgaZJDxXYax2ChbBPYopbXwf8aNa5
/4wB+vjzvQgK5OQkxYY+j8wkp3mDmdq1lncOr5Tshs7387p6dTpSgrr0vX6rMYVR
cwysTHiNPvweoV4bqJ4V9uYHN6qiq6SHH/whawZbh0XBjvcBYxr4JM2Vx8f7/z1i
KLnYzp7DISKfkDxLNsmq//DIColSEVHtboLG3o2jaV3GVatMciz7RUIH7XZNLOWr
MRfOcGCaHbQHpykghzDUQ2oUFMCPPOs6FZYZZITzI5zcCQzqeju9gDlnIuGDwp7J
X6Knh6O+Rt4A8qliH0CHbOrXCkoB5jHGp5s1yFe+yiNy9VUcj/d2M82MSxiUnNYo
ii+33CzfB67kS5uHPiaytMwn5A9a39G0y0BbLP2z8EHWGzWlwj8YtyvM+nF5DE1V
vPwH0nZW9WznlS5inoOnps4+9F/wpf6MWKcJW/Z9darv2seZQp7hN2KYZojCaStI
h8MmNWogCktJ955j+VXN4qgoyPz6BoeY8nNQeM/u19D0pkTqbiCXk4QuXDkFhEXK
xhY9W7XKIHzZ0PaPAzfdTm1o6RyEhcxX6B/gvSMtZr+WinFujyLXXPyeugJnn9uM
LTtfKNRm7j2bOQdEoyvVNpXcmgNuvVsb+rm0qLST1EMFCLXmoa3AZJsT7FjQZbPr
n+4+CM6IjEJMADLK886SMTUQwGQDGrRVSLe7E+FU5FU1Hg1tV00PkZgkBxupZuRq
1kUfljnm673/HckPahhCnfOspmHohF57AYIwARTaeUgMxZBPu6h8+AvANy+a87BS
3Tv37m0Mxi8ABP7EGWo0rq/rO+xctRa8gjlO+bdwlcRDnapl5KwA2r1C6hDrFwmp
PdDJQ7SN+VgVnKu4bGFMnfpoUjscDA5yv9IhPFoDWahZVwdU3yqkQN9T6kTXos8W
QhvPP3Xxl/j8MHZFm6DZGtF6bcEycHDLVsI1ORy+n1AuVvekvt/pNOJOk4MLcede
5Oko1Sz6a+F0M2M/iYcGXv3Rr4/hYCbqmoJe8um65zjbd5B+jbz8qbT2SkTrxdhF
rVaCAVw5S4o9MsrnG6ph0n0/otIPTmBhICaChsSEnCcvrq6KQHoqdF+0DqAzOlFB
YP9/jY3fLdrncKafY6wnwjqBELIilwXA8aOTWzCfHTbqBbPgNQDcI9zvmWuelCN3
DmxU10xjrhha7iwroWPZtGVjCHr8L3ynXCygz2d1sclSzF+sKb0ZMObMAc9p+zKr
9qpfhyCPSxs+wKMI+SHb9wVfDtE9LgntOg8SO8LrM2RbFpTHglCiDfkLPRIeAlnQ
zwvYEXG99wWcnPDLdAZlVfySodCg50PByFNXlgwbqKxKFBUBpIhDHWkujAWGcJVX
nHnByfcOZgVIWeTMahNXLk6duXzwC4nuitIuGGjZjz+eOkaDZEVCzDZelmPu8TjM
Za23X5LFJe5ujHUYtGzSmkIuBv7xJd6o4YA0OmT58jg9zV8TLRsX6kyIkOJGQe/T
qQhOVjb1sZj0Rw7mL3UHHVPfHAosMavFtKhzp3Il7MMw+yoYsMqK7JwvVvtIVXsd
g53AW6is+sR4BksvyhoQFs7YAuUCm1M2QA0zhQ8EfDIc6fvAdJ9Jxaicn5D5Z5pe
slf7bM6D7L9RRe3XUFyI/Uo9poDy6nRpjAjJTAYZdkQJDF5vW3a3I0XbfWxqiNyR
16bvSMmCCWf4pjVU/MGJyFrw8S4PPj7XPVDxKagZq91HmicvysFu8NtXiExVuIXD
o6P5yGWYkq2gbVnZvRhm3Gwn3OACxLiueibxeZ917wf8y18YW0bZmtrTBEV59UWp
TdTiL52buKxqirUABRHZEFC6eTLRRmeBF99PWQS5PfFLrYtnnz4U2ZLZ9RAB9sLS
J4NjGr9vLcgPuFU9K2Yqq6okcSPWJ/HKViLyx4aRGuIpoGSk2Mvrmwg9pXMlBhk8
Z60dPEdeofj+/mpQm6ID14MQzzkoxnb8xkII+6x8TPiAA90XE2hJg24gK5krsRL5
ILRnhUb/EyP3j4sjKMODyBjBASTZO0xXk39tlJx8tQLyYocYzOE8C8m2U9QSWuOu
C5WbhZs3Eogdu36DP2yBWlYsZsjq8PV94Qp7cwmzCS/GJrozbNyvVex/kK+uL00v
JxUG4WGmU+Jq7nHAYRHK08BwUW6tawcdhiGVbXw9VCqgMD/wZc25McWTsKmSgtcz
33BTzItdL8wiDThLJRc9FmSArYrJdlutoPX4jMbV3t7S+IhsL2QOX3PEhZMbQ7YA
K5I6hAS4xTaUvvssqE1CsNRmh5WbQ+fRxBxn3aRdS/Tx6V21OcA49mhJ/niyrw7W
cdPbcDKPpjIAu2c6gxGUvdPA70SY8ppHJPR66bB0hzqFGFxfuefa6f3zlIspVEWC
51tUwAhibsiGFMIQhDPJbFqD4kBvTODPn92svRw+P6vwh7jKApDMMiDeaULkFOn9
Q8xYfxjrJ/DxSKodB98ce3JVSRHhhCsaZUSzQrJlSeoz03B2ZwZfTSf3JOv75z6b
Qqiqr28jSU+fzgOImyL1QGEBTnN7umE42myQOmKBeCCQ+C4OzeQnnTWB9BLL4Om0
GjWwfZu9gcbyiDayYKAEn8WzzZ+7dUxFw/Ja3OiasXd6gJo7HGK9piPEJXCIxS8s
IChIY7Y/IKZ7sZzlxVaCLsSkSZEOnBL6H4QNdwDoz3lBSGD86C/I8AgOIStrcYhb
i5sNF0+XjDjfN02d8KNAMEOQL/TorZ+OZ9AGsyTZwPTTb/amIMUuLJd1IPw5UYNQ
7URNIorr0ugwVCglcL4KVXR+gdzisr5eZny1tYM1yMkL0qox2eIMLQfoP+FBRdVZ
SSHHxXWAkrf5EJxjw61mXiWQrz0xhDqCBbAb+OMYmzMOZRDnTry+rOiwOJt+5+Qp
1OZ5G3Pgm2KJ0Mtt1MTFDWa9PCjl5Tt8BlyqcOXpFO/6dgyCnclcNYJG3Z1E52Ht
Cg06UOHmyG25kIFX4JQg1xZxpWLTJmJPTMrtF4BqnA133Ub4w9AspLahNiufSXww
19ayafi8uFnj25uoGfEExwG4EK0ms56yPt5cjkO5jRdRl91rtneJ60fnsvHcbq41
NveptPOXHOjDiAoatsMR4EouGdNbiniK9rGarf0h01IsKZ9b3y8YJ6utMCmAKVLC
9oinCMJ96vUbWjlB+xgExN+IcT97BLO/r+lCq1ewKR4AetSC6SkqCB2HYtqXKM9D
pK3m0DO96V1Q4Zfw01GGwWbngCMw11AGqPcfBkDlhiU+aulMnIcJzEf0bDRiDQmL
m+No4EaV6LtdbJ88DZSJsKVJWKRQ6/TnvYiou2ffOqfx76zaCttUp0iTckiwNqAY
ob7FZRpbqjIddhAS7jlddABdfwGdFLWbbj5UILR4e0BoGf5SxgYK7wfyUUkNoKK7
daoNIq/FKt0N89DLTSVBf+Oggei+ZdRk2Qw3mf/z2p59m2NG9msDJ8pKKYvLUeJ5
rG4yGz/2r7PtZoiu/oI4M9hp5UFnir2T2BFGN+gbsGAGiy9lE/X5Y6ajGm4Tu7j/
YCN3CAk0HMa74cM33PrWWBnPqAxfHpw/YihBY4WaPuneh4NByO6ltpQsV8iwmANm
Kv9bu4+KZmEHO1VnaCKPt6juB2yKYXgtqpxgkbBQYGfFb8DWDpa3n8On90oI9Om0
j9KDR0CqcwS7X0BVi1wVohzk9GoyEA9g6/Er1EhdHi21PMwKjQ7hKfzcoVPgGBkz
pyCByts4HmEcHiSMCcqJSwHFWQEf1fiJ1aTH2kPn5wPQylREL9zQtGYFXobqrCiO
DCsgdTT1uX7eg8f9/T25/PVbKKqAoJ9DpUMoK9r69QDxfjB9yTisGYN/iZsKg+Rb
QjpKt68Xlrh2bnaNU8646DNXia0+dTDXm2Kd4dIviB2KbcKyI4Mx+tCOnlomS4Ja
2pmaTfBSZAgF9b3l/qJ22s9IspzQmh5njjKRuGdt9Ld8IrFqubfzcKbYQQqr1My2
FKZbdiJUpVyPMsAoFet/DZDXX76KSfv0YZVgbi9ukQ1QaMpkI5sj2HB0XU8e0hHy
R92CDy2q9aJQpX2V7hlMGUX6bz/4GsdFd70CPLKxx8M3a+R6SiRxnqDSFUwvYe55
BfGiMM4L9wGdIzblIJocSOcERqgbQd18i68H2rnm5glmzA3Hz+vPnHE8heWaux22
PKmEG/agcZsZtXJADHRGUwkHGG74jsdKw1GSwAyC9ucWYgjDjRp/pm5euHL5GNEX
n9PLrqSxSRkn64rrDO+ZvNNhExDOU2oAR4MWb0jnhsM6CBdf1nz/zwtdPlFOfwY5
Wk0mJ+wRt5hqorfMZ0rtCO6fWCwceBUO9rX+KKH1sz4u4K7oJYlyqarLqwwrSrui
aiTJF0Y6h/U1HvUJsAmUsYaU6V0cLRXK12hQ2FCJ0QvZ2A8LJd5Uhms1uik3Viqx
XJDxp9SxGwqwwdD66mSjMhXT9nNkTL7aLSbfKVecVRPsqXkpZqsiCfA/ycQ1iApE
jnRG86Fbv3cAOJA+7AHEOxQTU9amEKepAl4qDunP1MfqisXWnsCAUnYEEFCpUIIn
o98vhlObz06YKUCyEeqk34OkGMQrplP/5IP7bRXmeHOhbdCdQExARawiDMVgTBJl
Jree9nzvASWOMQr5xCcAPQ3RdhDsvaz3Dl5+WVX8MBYfTxwpTQCUzBrps4DD5IMm
51Sun1QFHj+g+NyDIat8k93kp8UJpz7mQJEwW3lI02niCRl4rdPvc8ucyauweLxr
rmcLcpBXEmPXh0l3uazgzc+3V37ZTgzKAB4RdvTKOEnBj6VwuyQlx+c8gQrwcJZC
40Pl1RtNeTNT0VgXnGmzy2yqEVCPUo7bAhiO/jULB17Vp/gmli9LcYhmPQPrpKyo
QPLbg3ulh19m90ykmJrkZMVwQ0QkMelViOb/7WZp+fmGLLKQqiXrtOFNsjGuqc0W
NLIR4g9nwIuY2YTdFc40UcPYqeEEbkWmHUUmYTNZxiMhApQ161/i0vGcipFKfDge
1elBdhBMhB9rlEJJCeQrBovlD3e9P2DVrXiC6usyLRxPeM6//B7knzteJZSYAkW2
W49PPZOCHm9uxBIzkVGYwEU4l55ZKKiQKwpO8eUmyeXxrr7M5P6pA1ChsHHKpfiv
G841WveyEu4slIWty7bTkxoYk10+psbPyrvVEpnIn1JXL01KNL2bNjOkAWYozXsq
G4/a60qKgA8g5vyavaHa+m8UwUnxxuGXe+6xcSyumQT9NxJe/EaPbjDgRHgkyqtF
f2GE5LTtpc1JD9XT9gOzIfxbpFZEsNGZW0AH9c2jucalKC+ZzUYx8t3D+sUW8zi0
fEsP0oH5wFjkGunTMR4LZOlOfdCAp4XXZVMcraVb6c8h4Trs8PFnhWSnq2Kzb+cE
dgf0Cf1bMKB8i5Hdrfwi0hEVMdjixl/rqGh7YdIT+F86YSNwliA2BLbIbugIcZdN
08CNIlyzAht/kEgyyy0G4/8xjyj1bF6ftjWZLfjUHgF+DJ4dmf08/yqZ/8qoUT5Z
DqHkM1LsDMcd/MLpdf+wws1OrQgO76RMlDEwHuU9oeI1SYpuOhIYqvv2MpFYW0Jz
mlZV3kZGmXg78YCcHW4wh2SqLAhiUJyywy4e79OnYMHFb0MLXwwzYrIPN3zUjkMa
dHaBgrsxh57HwVgFQLB1LfElQSwF38S1mDcZ1JbA8eqdasFl92FtXwJifrxXgRF0
a3QI6JSTReWRL9aC4Ndw40c9/hMcBresi1sc4K6zamSVle6imZjvv26XREyk7anE
mdIz42H81jWz3S5XqhMDaM79ngLSopDqBBeN1vCpnjXY0pE8x+xoFQxDIenqIi1C
gE42QKU6UPBuNrRv1yBnq4qwxOnqVVe5W+eGjRPKDXdu1U5SaT+qM25C45ybfr+a
vlZkr0dzodtTwAH5YqrVeZwAOTaqPVSz9RJcwwxkDeQLkgrKb6ErE2BRxW0S8D4n
YdBwcUvJDZrXW2lZnMZol50OwAS+EOBaKnjH5cet6nLMs++LX+FUiBfV/FO0OOhz
zld6hZt9m9URhvQ4TsV87BtL3Ij/9E4lRge7V0gzgqzm67bpeJBQcL5kF+Modgy6
O6Ub4iXzf66BNYOsLmZ0hj+J6Smg/RbchNzIPZYm6/+XMmc5ebMF7JHcUJoijvpD
uhiFka7L9Qv6dSK5zPpX+u0Tos73l2ea3NKmu2AZfSKUZpiNmj1Zeqfyc8w2uDqx
MZGeiIZhFEuP5xNyFV4QOCWAeWv19+zKpKSffCFSw28yuBH4AkKluOmKOiIQoopL
1YI4gdMnI1lf2JvA5EbabX2j3j0XBSQPp9pm5KzhFznxiFnK7/9y4l+t7PsbDPYX
RNr5//di37JW6UNSA6l62JfXgb8PECfcM8ANGoYq8U+swasixNBI2WyjqUE26Ww2
GC2d/oAUNWWb0WxEBwa6fSsitmI75eaBN1/0UNkB7XgorG/B2wEfmCVexAUM1mKZ
x/cWyMMcNz4/ZwQ+gbNXvUfoQ+LxiBzGe6F71jlIaiN+i1r9Afd7xkEgO5fAKQIo
onOKAy5wyec9sGjSzqvf+fS+dD3BpwszbMa41l7d3OQTJ/EpfrtQ0VzFNfF+FaWQ
CWDF+2EnKjbn5hud8Rmd1KHJM1oHJ83ZvLh4JFa4tkx0o5hY/6xNCH/4KZGKT674
MaxyilqMzhN0mZXf1x39rNqP7IqqZZEOIsL9ErY0BokSbPEoPZ2T4P7XgBZO3Aa+
11C/SrWIl7eTAEQCNIr5kI1gauQQS0f2qSFfMilqVrG5ochkpOl6qaQPMnC6D5/L
45VAx7uIDj1PgIsArrxM4/FndtKtgdVeiY5609vEi1ly1Qd5ku/tYHTWY/zgQ9mP
xLIoKIuzVdzpDj+t/e+B3NRpSiEHM0NL/0C3MkWqrDRKMK4lTVO+/kVA6RMfF77A
U1CvzPCilKrc7qY2Tnwu56iPzEEq4dc2Avhc9dkve/sMMJo/oFQxejJLEd+HesnW
UBu6jnHB2OVZ8RUjcabHpl+RkPAKDD+S+2vXo9WuvShu4R/8IAe8Fm5iUyKy8Gm/
GgrGqEfzDfV5D6p+ohGMpgDPL8OJFZlqRpM4N8aPqJ7wvYHKHacbrp2GmzSbE0bi
iJryKcZg0AZcC3CrAkgLSqG9GgDMBQoMZZOX5kf801L+Ex57Xn4aBI1emV01skCh
CxbleHuRuZz0TfNg8VpFCPGYDEdlJUrmwiuIqIicVfF7+zr2CHTmHgcm/1fRjTJA
CiL4tWb+cKBf74hU+ywjkWLKUQ1ubXXBWrv5YDuEZF14evTuhGwYW+MooDXIrR7r
d9YbR6U1mHGyj0lRatrgnIIlrRn0L7yVAMcP138Ki/f2dKb8866i8g/LvGS7ETQg
kugH20Nbl9FwoazCj6+Nqq/P5bS9D9Fq5fdpLjVHmF7HgCPAiBROqGBTh/y5uUd/
iOIIYkkqcsvc/0WBTj90ieeL4FCebKeOXnpLbr/F1a/a95xqGfP6mHNmc9CkrfZq
zFrC9pgi2sFxVO48WmjGeNtmd4ST+eipVrxfj7cv0NyCch9qMVIYRsL8dpPHQhw+
/R1reyFTVBQCHBlHbLaO8TH3QG6ziv6wDTcEfVnsE1fxUDY/xdIpuimCj6RvCSa2
TIK0mWePAwL322uqrNaS0nwCXAf99L/iZTGvXN1PG4S+FskxtPU1Hs5A6voei+Qo
DrguqhajZI2Cp/z1QgWWW9SnubpDXoh6qFnOlxtbkiKjWzx9BXfmqeIniXEZ8SMU
hZSToKwA3EeNU+2M9S4iWYyfEbeMg096eRbnNbN/C67aVniXgcj5HarzNwuZa5ZZ
YvgfBFQO/LhLVp15KffqSpJVwSX2zN+9heBarMA4hSGLODIltpaHHVGHRePX+5cO
p/rT5a6SwrcfUCtGTk0zzssj649r03pUSxUYdGHF9CYiCT1o+W8eI0GPFDs9a1o0
itDlzCb+UkxlHtqI6yh8mT1/CiRIm5Ljqs0EEQhfHMjkgQkel6XcCQssM628DbPN
MMued35JeR4HqFVZp6MwWsk5ro+lIazIbcgPmYdoNZUYVciOhNn3p3pZwJQ+qTZF
NffYUtOF5u8Bqtqwrrc0Q/B2vcqDDX1Bkt7Fwf3q9mOypsQM6VROQhh0NjCIxs7k
dqZ8C6SXkgrRUVI3j50uRcwfUH6Ee5JJxCwZozx36kt/Q40hxrpweaqO21jDzWtp
gNax0PhZNHkURtU0TS2FbioZNDx99regB12td46N32wVZQ5XaaeZ6UttXvX9fRXX
u8do8kwTzShQIRXuOu62SX9zy9diaE6eNNJuHeYajmw+yFCayQklWEUz5cUjks4X
N7ToNn3Dvb/nz44nQ1eFUsOg8fp5PKHcu/cXgZpfHC2905PtbczeaRRu0UxYF0OW
CLSK+i8MOzk95vjxMFOQH5yiFeGktTlzWNSvDsrnk1gVqxQ4/a/raLuRu0P5puY3
UQI3fKU8HdiWvhhzKBfDzO4KSqxjqFZjrYDaRlh2gNe5rSHO4SG1ek6+O9DdGpMB
lQAoXm+2x8mVsFMk+aVbHh8Qva8wnPeEGLN1S0GZLqG58UesZXdLljeemZRREC2m
Q4WnD4CrtyOMwlTVZpprktmDLzTMhQV1u7leM0AECiWVG9bc0xoX2/o3cLjT2DQ9
lmJjftGqG96ZRL+VTm+yBsJ3nhC9w0ln1T1SThfscKOwTjYcwLGrFOkYKZIvTTKt
CJG1y+2xaA5tK5sIoknubBxaRGr2w2xxO41LCb6Z+v7FUzJZYHsdG1s1aMeak3ME
6V8pyLL24MM7C3HJCfevaNNCmzYpt7uADT51zdqNwVwbJ8t+a2FZ30yhCyNyBPO4
yl/4rACWkyrWkFC/B5YJD3+RjD4C27vl4LGfULWG4oEML+oxF/GiU3FWU92s73wU
lvVneVcC7ahZInM9i3u92IRW6nrPYJEZtvaM+ZuzwODP+H9p4VndPJhRXHAK/rc/
zwW+jYK83EH3zg5JMZrJo2eZgMsL7xop8tpTe9NFz4Rj3orl1FCdd7xwDtsrzEo8
7T8HqbEw2dwszqyZ4Qwf7Bz9Mdv3fOmJt++qavzDj+hiugHP/XhN82zcw1037zfA
lXra2a6nLsRuRsVxGpzPeMb/i54IQNCVfsid7qZRI70m6vJq19VCHCxUo09N1wCo
7JsGnBsT6owuduojvTacz8gdDUum3SRz8dM6wySkQBlC2gpHkv6xwyu0Z2aLNoqO
XbBm/eZJwNtgo7Jitz3oa10WqcjM7N2XIX+P/RvIMr8FmmViIatFbkCMOpowrhW8
a6/IdE4w0N8wevOKUpWs6KFyy2/1CTxaVwlvz+6sIKcRAyqOrOralY3hRD7F5HQW
NYjZJ0QMRcLl5fktgCsWTRWerIr7IR0JRP3Hp0igXRfZANoiMGOodExPzAdeOpvE
8Bmiw2tCj/6mxJJf7KTHntxggSEuhb3Ki539EPWhE+f3eH6kqGuK2jkJntZ562s8
/uPaDC2DzlSFXt67/eJIoNUwnl9zQTQbGSF8tKDCkLJU3mKlWGaKXvDVp0vOR4jB
MaiWPqSk1KuxBCyHwUnAb5+r/bCgQVuWnT5MILa2RDr/O5WMg5vGQzgelW3GZwWr
8muPg2XUS/E6N9saH56FTAkDojMJQkD5ab5ALAQ6g++if991bHGCno5NhnhWrWw4
FlzlfoxMGJwQ1+9FrjxYQdRtfj8uvzeE71uLITfDkEM60AMw+YSVNZXoQNep96CI
HSf/Qklh72ZdRPuoALM5fcFEhGg7gLuv1uTHcxwnfqvjNNFncZi5Hif6BHSAsTmL
tRJeRSsNQlz+GpaULC7TZYYWh3TaQ7WVtawLEdo3JwUrbF90J5Yb+3Luw8b1fset
o+4U+Pro1y0cHvLgi5eSNhE0RZbyic6oRpy5AHnHZuQHB3TgkVl0wgGSdn+HJ1eW
wKQRylhL2OnskVx4Lpv1NtJSrzKcIUQQva03qynn4GSo99F7huvGr+76uXHFDQjV
ykV1l+0+HYz0jmHuLbWe09gweWEY1h71XseE+OVL+kIb7QlYe4LQUlX4JaWNqrlH
1AVBC6XGj8Odsrrt8dNeRZDawjgAdknEGuGTiKUDNU2Zex5gUdsm//uYFd8RGsQn
UJesekld4MXnD5ohkiL2nebT/PSzbkHH0shICiwrMqdImPc28xkrB8bwEBxmyrQT
huBV+0X5tl/rt0XaCQc9juYAIBLFKRpiObzzq6bW3SOpFBsNWyRDIzNnFnGFhquu
iA+QBNOb9aYxFcwFwrs/vpR7HcWQw8zPH7q9ADTPndaeBpPtrV2n3udTR2cNvazn
wJn1LbRFpA4LYhccRCm4/qsoV5X6T8lZjLThpXFUiTyn9OvPFfH6frLKL+zXMQAK
lxzUtpmDWP1wBu4W2lAqXn0D2Uvu7aJxx3IoT9bbnJ6VlZnjBUaVX8F/jokyDGJc
lshF0PZgRBqt8mnBgF/RxH11py1yKDUUngOuIHdatXNMyZuKAL+VyuryME1F952+
CbmelnVUQqi0isuwFrtZS6/x18iD5WaY0R5Z9JTv/plBsCgVclWn5VlYoUf8GUWl
tUkKQ1LArzZXXthNHpzbERuybODGOx2h3EqvcftjkJASmBOAbpPYO1J7kQ8weRvP
DD6zdCgvFV/Kmc9D3/5R8bzTxGE3qXGNwy+Guyc3ndC75Evv2Kijid6XOJgZrDFm
iLK8SWNh10u0vSyJcOIERDu+Qkc6WBvEntcYwEqVaPuE0svKpTBCYvpD8UnTx9/4
6vGPUxVn0mhhl4moC3k8a/gHFZe8QLRhT8op/r1j1HwfKHclNNA2jjw3QQqRs1r2
g1B4ckW9eIWlxncHntL5ecMWdArgVOZF94b5yCEWnNwy2TR4XrPKgR5i5vV3jf7E
zVR1EKGiNJ3EaHNE7d5EOa10ycGCpfphZ0rdvH/ZZOQdafFtkgt6tQex0PpWrja2
Bw7iGx+ek69Znu+4SvnBjovuDqHLdymXrSzf3JqsjIHnmyLGDlCxVzAoLNtzypkF
P8e0fOslo6s2tkQLad7QeasBoMw3wvT/lq+iyMyMmaZ4GQMjukMAIaCh5G2Vd/oH
gmQv4j/4i8KIHMWow+un4JUkuTkJGpbDUVYFVJPeXlHghf7wnggpgsEIsOWn8/mY
kGQzwuzWK5dYpqKQ0z5n+yxzEUMv4DmRk3E7casZPElIFmgC+2y6dJXYxvaJbZkJ
2Ujb+ldXFPT6dbVZeeigmHSiYhfO5YUC59qsYgXPYL/arlE1P8MQrqdG82AMjCvH
kGMYgMnF2Y/kmshQAIvodV4WOM44Ky7EYH1eJjDF7OT47JDjcv52RCfCvZHv4q4m
Ex6eMmZu1yhQDF0GPNpuwzRqVOcyMNAe9aklvg73Q+jCbeU9f2q6CIUBBl1wwesj
zeSzOTqNn9+J/OlixmFHmkmW568U2vuqEvo/nDA/fHImfbax3q0Tl5rCho5Hgp48
hb6O4nZEPpa3+szp25H4Yq/0l0mo+IWtSZdUbOveSeeLdxMN9sJMG66Az1UENP+L
J7CHHvJG9hJbwE1o6bFHTDD/vJyxc6FLkQidUrCczey9SNRNjpV9LOLTspdvSyP1
X7YGNHbU35D31uvB1wXDkGasC1db7YLWQGfVlW/mxiuCjBCf0qPQ+OmIURATt6z/
Q6Mo0sL6p9Q6Ag4i/Ol652+JuCvlQ9PcfDldx3Q0rBswZwxKtdEAHaQtCeDLtdJt
+Uq6xPi9bRiY5l0URPzrZVIBhX5oXgaoJlNbWdFYtyZ8l0cpiHPA2qsJL6GI5hJm
1jwsj099vExGDtCQ/WaK5h/cQ8+HTKLOEv6RCP4AfNR3ftuC19JDgbGfXLtk1ulc
HQBBctpv9mQ22VbnvAY58Q1mdvte6X2/fbPQqPJUYvBX7jmTgBhKQQy2MUT2FQuW
8aO8fK+k5X6u0UsrST3/9yQIPgRwz1lDccwqCucu1PaeadtFW0ceWCAqtTQEdWbS
OBfegm4+QFtenIxg6IW3pYJ9sxyboW7QV+Mog5ZtJMl5g/RQ9GefQpuslAy5ksFC
HLaCeFmcunyUnwlvQqc934B5HHH0d1bVLHhkliq9ktnMvo/+kiK8LOLCTygrCqRV
dn1Uo0RFvMHKJulIjaVPNNbKpzwYrVFvorJ/QR8q0MSY3F/YBOyFGNV1BrgN2gK4
Cq9NFPyE/59vHsIIgVGmIorsum5rZkgkAv217OHCgk2PQda6MtfemVlbCpCN7eZe
RyZIL63VAA/EThENxZxFGPwlsO3LrYSN53dR/ApFeEU3M7vpFFOt9nhFB/5c+14c
8jiRJ1AoIjpYlO1unWwny5aqFRKjMUtnlSWemZEjpyIu4+PKm6nZC6QDJpm+4XRv
w4799NmXBdnsc0EMBdFznzt0cw3VBKeEExg5jO0QZ9gQwX+eZUQ35lMGCKKzjZRJ
Bf3cvLvB5e40HFghArtb1N0jciD6hjD6Dmf6zVPliFw62Xmno2KSugcHmMvXlNJx
6Z0aaBJNRDrYUZeoAnNnHaBwPmOFW9lM92poMQbZYQV5vfILrD3+qGOziZqc6Dyb
42WdJpRcKLICYhi0V85CC/kL/+bXeocILDYsNrgdBMGHmgLwJbqYTYY7gcgSUuCV
61dXFtYlrSRv0Ai13tnneLz0k1Z0F6CorbZ+PFSGsaKWAf68GRO6gNehPZhgh06/
zpUgPU6GBn41OpTMGXfdsAw/AMzMDdji7Tv2u7e4kwPja8JmQZsfB3eJynxUoOgL
fO26ZohT+vlbJMxYrrQtAFyEDNC9vG1y/9PiwtxIADi1/r8874r+NIONS/e8xV88
tcFAlD431wG9KxTLPbqOHqMw5w4afMTmNfOB3v7YxBN6WEw+PaQpJ3Qv2zWxedv3
Myg/7dLqmvHR7jlu5h1KhAJ3dtL67JsFMbLlCdYdanDcldhiE0HXaW43dur7U9uC
0VTDs9tvHjhCK4BaZY7e7JHsrhwiS26BVQRYG7Njout6NWN6b9DjE+3SbHj1Tn1F
FoJ+pqC+fqgL2bP83ipWWl99w6wWRJtzrijF3o1XQp8CDD7QGa+QBOzhVbFjTCf2
LkaiNoBIYOEN5hpJM4tz7QhBnWLDdSz+HjOHYvc9sE8z2IWlEhSUwr4fDtZDKbxc
NXxz2SKkvjpSdfzOkvO7i9e2GKfdBnIDxlGidDFMHZZj11gGMaNbD+AostWwCLwp
nUHpaa1CGfWRYuxGdleELa963lijnPhHia8Rmr1U977fE9XzLHk79bzgsQ1AtB9W
tE1jhKOx+Ywg/DzcjwqDlrkBh7mPSp3sy2m86WCVnIBGWqRPtJblbifgA7LA/5uN
riqEqnRx7gnXslvL8AbXHISa4qFBhG29K+1PRoJQnCeHYVmw6vKL1r82IiIVwFUB
9D8Elo76OMuQGvA8kkJjTpnPuK8frNdsZYImgBeWFkMXUW1mhuhrDX7w4SPFNhfq
CJPJ2w2Zb6meBBsgQoAg1K0STX7EDg1clpBdViqVYsAHS7eCIzzEWUKifcc9oP1L
dOrJP9s7jO9HV+z2GLft+DqLgXD9KWyJglYayk1ZlXg9UrUrO19+5/7VnPnwXV4D
/z+0AVaA5Rh0leluyYNAg2kks2U+qBD9h5Gi2BvYSySNMBbZxyfuYr3vdMZKUljr
QK5SJKPMenfta54+T3XagrwiK01K6m0v64dbzK3ZCLDq1204RjGoOyDGETpvxMyN
IZhHAv4FuRpceQaXUFqBZki2+aodz/mFcbTJzASpOEC+FQ6h34/reae8QRlm8YgX
6znECeWN6c6VidRQiwNUrRjnk16BoJtClwbKQeNL9/Lo0Do0RriTPFnngvT5hCal
wB5/e7Zeg212oAPIo5sAqloFvH8KeH13NQDdji4f5XkTh8csr4b1N+i/7GPIAWyB
EGs83hKBjoCFP41T9G+lbDs1lkIhFhoxs1O8bvZnl4YKii3nd/Q1uNJlUbkDYheU
aXeWPe/cVe39/jQ4zaAWCCHExmUMDYaQC6X1SBy0Tz9KXgHS1rdJqHi/MC5WQ9NQ
tSKHZxIYqX2FjaKH/sjuqRW7/F7+Lybmjn8UNu46cQnJfegQydZbkHqVMxXB+3PV
ES/WcHQ+EuTbP9zr68DZOACuHCOumL7Sx95qi08isji+VDk+Z/Pu6waMldbFTrJm
lnRiPwOXQpNKqDKVyzEGzeDreTp5mHAp8obXGF5/llkqQ0pC4FexBd4+0VqNdUne
wQbtD65apyN1wmp8h72l1zC8s3Kcxd7jE6OqBpdmIuYJsJ5YU5YsRlGMqxw2FSFI
sTTrQ9MjKOdOK+iXlhiWdQvAKK/9WsfeXBCM/wMyJqMRFaR2waLCo4jWHrup/dwI
RsMy/QY9orhafOCJXaHHzvB9hmSXI1EpmGNlfJpncJyKkwZaw5/QNqEXKfCfN7yc
V5XNCfodYeghWOI9Yc0sz9W9qdB6Dyxoj08NuXUHToOtq9F0DWya+KrQK/mFM0Mc
rT8nv74sUuxxMs2nIly1iW3gGQTjKHnWcKw44EB82dBmNCJnM8iT1axnNFMLfah9
ZcdZPYtpBBsd3JCRGwnLaP6CsrM6tIitaG+SM8trESu065FGmzECejW9VnX7dQs+
slGan4ad6TsrKkUY4RXNNwkOvH9jgwd5cor9YZ014+nyxJrYdyR+QFmuGTWfBO0e
zmB0K2NXGqCIGX5nalgM4TOXfVw96JMYh/jX09OKidvO1g/Lc9z2BK9l2/Dh5Vq6
qTe+8tQD3Mbb4FFmVopD5sgqu4FpcMdMzuF4R5kkVX4TFWAC+JHiXJOTXq/x40OX
vZ6o+0tn0Y+VOBcrnQIO4dYBHl1bNltpQ69RYRdAt4hbLYuua8WPFZb3AzTwNikR
8xWCpCNYOqeJDSQiUifexuRnohNjry+VZPTj+OEZfwbQCzSYYZ/M876UGnm6sd94
WKYOcLp5PkyCe9uNv3a1jUStudmP48Wv3BJ31WRze1YXfHXNTxh030IxC3rNMCAU
YBfKObGZlfwcJqk1IzIrCNpUwGbtiQQTHJyjeqY7OjpJUt9pAH2fkGu4xsuB1rhB
Df701g1V6KyJzVHPbaoNcQ2ThDKsdWQTHokeGKLLE41SsZrsvxKrOPNct1GNRmf5
mFDbUrfwh3G4h6SbFRH3LDTLxkPTwVesFLlCYlB0iUZKrpJ+1Hf2ooHRUpdKFf+Q
JfxoIxoEUgWy/fs2mB499rzdSkB5RvikeMS157JGTYkMHwCgcR2Dfu2+RsIwpKDv
rQYSZXm3A7MoehW3Kv1/cc627n1/anwRAS4W5sQjaid7xl3d1JUB00snmQbURHSh
WYQPkZlrnZTnrqrVJSdvlcYDBWoL9v+FIPYWQUF6QrhHfX2tBDsaB1EnhFm/vqfJ
CW1phL32ObSP9PJU0yLgtTDHuy/MdY/HixLQZfSGw21c6gIzwYRz4sIHLsGsNkYn
kt9KUcZ3AtG6Y/KhmIX8CBRm9//IdRjq2bQf1m3EVFsDWdb5tqAP1wpPJpMrgVQP
kPN71Fp9EwDTtF5eL4RUcRVuGGb2ZL/coOYwYkZA51HystIAy7Fc6Xyut2R3Tw6E
+5ngy1LL5B91H1TdwabG+HQuBbU22zm5yedlssTtTYqI/8cN3GAnlX+5hpEaE0Lp
7mNFkMDz4CsulEmaelelLWK+DOh8gyLQGZCF9liSbznOLlABRsEZHI3xAfUOP1Ji
9FnnvbyTAzolxGIKGo3E/YLONyDTnIIJG8PMU6a1Iku8U+zduHfIdfQbMBtg71Q1
AxtBaCVVOP+r46Bqzvf15wN6bdwjRtojSCAz6pGIkGApXwFtQodNgiBfGI0vnPA1
Xh9CmDwaYWM53CiraA22Go7LTEgyA/9vyjc5CiR2prdvD6sTBJMekHulalEXvmxm
xNrQu8kUtYDfjyQ8Jls7HJOvUGtL+CN8g2Xc4w66dvSiMsk5YqWmAZ2rTj0T/BTG
Ba6D8Q1FXZWqv0rllY/1yeOHFjToq1sfWcfIyPiMGxMkraARn1he1g8bluNTCTya
iqK697wLnHfkTF8xikCZu2m6Rt0dOyZerNo1ObLBO3A9X28UgAoNNJYYAbqJRjAL
HRJZjdtlir7xXEc8byrG8GEm4apSrgmigy3zFWvbgQVlZ7XrOxHAhC2YvzMiHbxh
2Qgtmlsnx1d3R99+HovRswxz15KAHwVZxR9kTJE0NrmZxzBU2IBpLuIUzA9FeXTI
VuQymSrBQuY/dYLIU5I5Allw9RHtgj3SZArjaIcEKzEbZSIF5Cr3XY51Gd9OdykI
FwHWcuosAvQILPoQrKQ1EFKxHUcUMehf/yRDGMUSXXq5qiud65v9wo4ANFSeu+PK
ZiPIkyZd3Tj/hqo2Cx5yMWFOHmyWdhxxq99eJ7i3rlBMAM2owWfcYMOxcgeOfn5s
lN5z0FBMVNdjjy1w13Ka9O+CQIMRZqzeVO4AD4g2WVpu79mLwmUdjuh/U2K07m3L
vNjfOgc9lYsmOIRcCcWzcY247Wt/v+SnrUq+jSBsSG6L0x8uG3vFSK1r5PJJ89g8
HmrgjV7JAKcTCTK9GFlZwlJ3XLdeOSmzkIv1ADDHM6f4bFYe7eEcRgGE00+oq2uv
FZhqlBJk00ymSyydP4f1SjumDteIYTpLlNJnPj9H1jK75Gytx2Nk2PjrmLYOxnEZ
tldM45t6gigQCzZlpH45zX2pSTDHnkAiry8/I0FV0N3yN3iJLV5DvM2d7wD0+lxs
G/aArdz8U/TkAuGbVlbFc8SSYnAkZOEPxflgz3DJQFUN47c8QybZZrpL4zKMW/Tt
AAyxmhgLy/iInNxH7m+zVGBVIEkCBuyDFi6zAghpd4oiV5rBzmIW+gRkvL/PIKob
m60CMyyjb28C7lZsKbIf8jAKD88F6HQUCdh5wZE/ZtT7K+GdwUurBOZxN4I3bKFp
heGRBXKyLHCefwC7Q5kWNyk4Mw+rSln65yxspncWNMkwcylDc+XUnMVZPEyNDAn+
ES2JE6HI7f3AQ/aygMSF1/1dVjYtS3dTXgxy6fpeiZ/pT3Cz1SV9IfY6R8GU0AE5
ZAeWR0+50/KPbFINpIOMFouTwUkNIjPkD2jDQbyaXIf14EmHTum9b9inIdPzeC/y
4+UdaAGLKzbkpmtbWXuABtJGioXZhFyJtdlQZTeksZZHGnjrN3JbhTxmfdpzb2pI
nN0vyGtCMNIou2LT7Xbt0F/ZqlT0OFUoqrWQ6BbW22wWK1eYIDDvdei8mXzxwsvs
Z82g6/PQUiaQSoIZWx2pI9ptSAHzHd0jUPOysLoPnw73AopK/+WoanXrHKPtc20Q
6DgdjxyD+uD0i+q/Ryrwc2U46fKEnLJ3EAY3qukbPVL14cZI/SmcEW6EpQLXy2t/
Tj+u69hYwPXtp1d/JeJyJcC5hl0RM3T/XQD+VssoePpcSwBo8Yjdqta0bnTp1Qb3
7yKN7AjbRsF9g/h1HpleFWO1BwKCY1Q2lwXiYZ4wK5TdRi8vukDzH202aUvBYtZh
Hbu4KgVlM3I3Ya9WJ7KKHQie493WGF5Xb281fRMNnTJ0bvihhCAKLIw2alSmUZPF
rwHZGynZYBomJhf35eWuli4OmLFzilKmWRCiveKU4uthGn9kK/1nwn2wr7SwyG9l
j+5uiMfGWVH4AO6trXwsmx7kgPXxT0Rubcd7jE/vBSUI0OmgxuZlfOJ/TdTHtZ63
8IfA7UeFLLiGO2tYRI45CRVhfU723MxxgOj2m7AgKvIcIjye60wKCjGZRg1lDfSS
gfH7Ichp+Ew46WpOzugQzpfd5xXAjHDhNkxVfGMubSGgPZSpyMpdHUiZGC9uZEhD
NqXnuVcBmpMLxqDScJ7YqhWnfY3MKqgX1R4e0AviXS+4vOvlPaH8uP/GSvAj9Xda
HjGylPnNTxpezzMujUScIQ+tmT5oV6k4d2pmwh1igBwZT3KtkuTrpPSu9qptERTh
xqUe5oc0tqu5JjrBra5y38S2OkZS9W6Mn+83t2OPnQkju5diRcnZf1s8Ngqhi8Xg
AJucBZHEZTDYno5zvZQxKLLNV8naBu71xn0r498KNB0Fq2CRnASOlEtxZW/IiKdH
+81y5PDCTe+WFlgxbU1u8jt8v744JS6mYeEkcJ4nDT8UUir9K45n4SDY6BE67MtN
uPeLyBloVvjiPWHlzejroMtgREOypeGjEt/hB/WmTOsqTsU9KmRP2h8NzRCUW2tx
Ub9M31AdXkbSxaH/yG8/73Yi6bURQFw+SUhjLbl5B3eR49+rZA9rf5AMquT65YUD
zezTylBRNPWRldvag8DSA17x/9erB9P3LYtOH+eW8ZHAAHNzmhZ9JjCX2EnPVLkK
WX4ks/L8JN3FPFDY5pcLI0YpkadYXMnmAwiXTeZx6MVWYelupnfTwJdQ1934b/IM
6AIOtV4UXWS8y6PodZYMeeGGt6PXiEvADauTGlbhUlpXyjVL7gB8+db0r4rnQLZ6
9lGOT51R+UdBguOBj3qn8vfK1Wm4u9MCaNhslgjo8ysW3etqZaBhnT0zp5Y5GTDl
3YtjvsEyxbDhknjba/cBbQB+WbXClKsfWe2C+IqnZTPFuvfYyJcWc77oat54Hy/S
mo7NJfShv6qDKECroKEFtvDinoRXh3+v4XJh0ECCiKrHzpga2Imphl0znlvpRELf
VGEec65KP5+fIQGuaCHz6TRRXcu+nHUtphZrgbai5fAXMDDJO4OG5YBRFweFtdim
Ti/5O/aleqpFzg4v6gX+BidqeXHxbfY35iORFAs12rDMeI7yhkhqS6twF/l7N2F2
+AyysFaKHkwpToUygKOMJP94NU9w99t2dnzQ5bxkLN8ahPFjZz/QXk4I6pci2Km3
l1LNtBGXPzWItACGwfuZeQsQmf6fb36JoojR3x+JephUJnuVisAUTzsJOJrtQXZv
vkqT6Hyyt3UswCh9sy5ocStpqhmn/L2n9Nbw1eYMVa3RUO0QWIa3/OI9R+57frJc
njr6hnN+zwUqY8DiGRSYdJycmfTr5NVrsVte54u1UH7++Zj1b2BRrLYiWEafRbsc
RdZQL/7yjgkB/4xRuxe2eg+pnICCLd6qxjMzadDCcOYOlxoxVMuH9XvomY3FHtab
3Ayfe590NuqrKNaoGpO9Njv+8acE2zRFUtdDGwX+E5u+Sw5S93+39/pRgpkwnSRF
fj/N0Laqr06JyKR3sxC0U0jz/50WOze8lyEQxELi8SIkXW1fza6auzQkKiebvBFG
IJUKDhCaGFr2T1ggncHrp4Kgl9Sx4YuD9XyZl4zlGIoyn02NrHXSxgzlCs2J17+y
SfZbXJ0K3c/SBrkIjUqihodlb/gTM8gn8jdyiSMhB+++py3oA1uQH7VumwG454M9
N/hLABbpjU5U+IjNg4zU5uFe2+9lNtsgJtkTPoIey3XIEUelLh5UlGabmX/pHtGZ
W9pJ3UL3q0gc5w9LtLPbTLXHqYH1tV3x+ZTEiKr7VANL01QWaxOGvZgxnoI3JvMu
Bv+OwybdtO0ZYPRgMhmWizdNseu/R02ExeZDyDn914b4hiEy09Q/5gfa6JPuDCC9
s/wAqMi4Gz4j8RHYVar3DCyXn7FSAFfc96TggxQp8ejT0iKRvLMe+HuuZTL9Sibp
qa2r6AxbGHNSuU9fDM2+FYU9u8EGHMekcOfxYpSTHYFlWlOunNgc7nIqiuWgSRqv
LPjG4VNoPeBJ2xxJ0DgHAM7coc/iopwG+M5Jh8S+gGxx6FmL7Tp2pvMtcVwY02Km
79Yh3/yvcD87duKBY70E7TJVpsGmc/WizR1vt0AltvYdPFVahBX7FbKzxLNnoTt5
QN/epCpTNUpNQbgRbElpyFvHgIdZLRecOvZRL4TeSO4aM3tZwrc0nI/QQIqz9wq6
s/ob807e8bRgzVPsRVsXRiDLx6zCHaEWVmlM2u35CAXc7/Xgits9p4N7tw+ifIa7
UDmkJIIeG5XKNqvoX2Iyz1wMxZQCb93BfZ3S5m8lNt9m1j6cLnyyphzq8kGfcWMO
iDa/uqHSy3BeNTwhRrsoc/Tt8WBTG8uTmRHXq0C0nAiMd2DMgAGeVWqw8VOP2v2I
6QZhf5wfvK3MhMJLmemc/S3tmJKtI7OCDzbLJT1POONnf7I0lXIi8iaPwfM6u76T
YlmhWIyn6csv0/yVN6ZxtCFq4xUZpaAFmdy0fEDC3/8d5YUoHgev2Xsr+YAwUoQ3
G4fTs5+ElFx5b/ErgsEcp7InK7xf5EEHuxGXt2QwE/b2uuODLWDFT8MrPg3Mr8Rt
qnZkkEuxwTd0BdAMV9bWyd/X7xJwos0pMPYU92Wy78da2YkbQEUUZ/y6JububNZh
b9fo6quLbmJ4A5xJ9XCZ8GIwuKLpEdWqHPOp63MamNCABFspGpluW3xOZ9v2b9H/
D/XaF4bvMcwD+qAc0JQ4ZsyhH81DOFJvCi+/vSdxnrDd3DQmmlIcHde8z0RuISQZ
LewD50226uYPIAoQuQZm4L2hBONPqZv9HVW+ZXL8ivYkVmhhdPx5FFrZqyTB7FFf
IMlIIrwm2nnRAjAFc9kTE+eMj94n6r6tnKjThU48tu36swRqwIYfLyEQ8pXJlnkL
gxdK1RQgNPnwxJ3GYmLfQGawy/OvQ2i0IW+03NQ29+zljiXDeiT+DPR280nf4t3k
OnCsFtzqqu/fvtgJ87EX7XuROCgjKy900epaam5yC0ufh0MdmVqiS/2cymL3LkZC
A3H3ila5glBibkjY+FrjVBNvHI15ypoHFPEW/OhyCbFpVzizFWJ8FVsBoQcNgqBx
hDcofQDFGEXiNfqpG5otclj9yfzHX2Ay2iuVrhXyNb10ZNlA0flAr3O7eCI7jpbp
7Gx0kcf6I9fvCW6wQVHkQ/gAZCn/LWisbt2avb2z+gZugW89Sbiz833OFlDjjQHM
fKl1EO1yOdaw513e00j8sdINEf5+w5ZxNRq9mJ1Viv2XAx6KvDDqUHS17U5RWWaF
X1Q+I2W9K89XCZmsO/GT8I7IV1ooGLqNSkA+nYtymYJvbvoVgJsuqhsjqdJT7Vr7
i2EjTrAXKlT/oM1jHl2HmBIKHqSpdDc+eZo1EvgJRJZrHmuf5mHHjlRSs5tkO025
CpIIpeZDeNo/KN/j+R0DeOvqZoYvSQrZUGJAzkEiCEhlrcaHQkUZcIFzYf2oQBek
rq/nfYPNrsVS+YhLFN2vI+VIUoGb3aNARYVYdcQvjlWHpR1JpXiJHY3noKQ0r9dK
bTt3E0pThzg0ALlGE/HOYMi2B8lRXcCzxxgq+kfDLYn0/n2/vpcUv6Kt+6seik3G
VyYKj5iQQe2zGeu4WyWNI+RgzLnYYHHdv/3gOGn4W59x/VX3+IEHXQm0oyF85f1P
G1Lu1YE4RaEIAxI0oS6OO/e2cKManMP5PWkfzUbkLTQeHbe1fEO+B8oG9yubL9Iw
1XPb/V6Xgm0pG0bkq+X7efHXKHG3bMEbTD7PXWx2a8ZnORR8pI6vHnw+S62E559X
jVizYvtOTy6egjXi7waAuQLaFAu9qNENuXcM4x30uGZfTAN0inm0X5GnPN/vUggA
0YxJH0j5QtoOqALLSkaejOyi/SZsiXgShutg5uUgVgQ7LP8cgX0n4m5TbS7G7lwO
//CxJjs0IbwxivlAnU6Fk1lun4wKEB0cGS+TRLp3K3VFMsuJz/oMK2Kq6T+OXhuz
MljDeNcAZk6/YmKpMS/6iF7gjU5DRwLW8wl0NmUUTget4TP3mB++5xqcdqwwoqIs
UDe9xc5jPBEbcPlt+Qf5wOgU723iIQQ1ma+zbKlnoIeyN1Br/eQuFHcwV9WZxM23
PosCHa/7egLOPgNjcosJF33+z0lymH4fuW4b5HidhzMkPaDLKY6MEPq2pUyzIcMg
ivmqa4Jxh9Y2Lsf6I1ufHd57/xWJgxZd7ceJaD+RJhqP7LnNz+vDyKSbYxgoF/eK
QSjjSJr3nHP2skPDafPrIRsbAt4j3REAw6lUMNltMe9anjhOcR2Xi4AyrFct418y
ZPZvw8nIr7gMw1q5K9zkjyt/QBf72O05+TvcdZX3QG208cj9lVvXglLLJsnl7Wyr
0UxyF27Nip3XotVgBm5oyPZ70yRVqiTH0XgkrtEBagGPauJ/zqx1HM/N4DrIdf71
QBxfzOrKG/iezCFxrMl5eTq7F4E+NCsrO4UzF+3/+2rCl12o9ZYqEssSwIOpTVOJ
uu9pZCY3oaifRJb7oz0dmPvCXZ2KYsIYFX1nOKB5zUXl8zESwbHEgXJR47MujMPw
EDqKGoZg/luF/aMMhLt35OTxiYq8Tn6y3thRqTufxhv1ImBh1b7CHAgzv1JR/1gm
5cF2OIb7kp1tFPuelg8UfFwB25OUmW+9w8Iz1bU3HY/5S6QeRl5g4AETU89QgW95
IId+sxZSb0lCkmN+HXDimZIkJ7ZrVjkI5Ss20vmZH4s45b1cIOLquKPsceocTcWn
vusc8CC1TOf3/fhtLz8i9NKFxa3VEH0vxntAQsPZrFTZytlmAdYu9jXxhd3GX/BZ
7o+CO1MAtXAHTgzbaKDJMSUql72rHQKdWmPORH0D27X8WQ95bVxY4jLbNBB9iGxf
qQzu7OFP2mcNXsaD84wVV4xIEJbLwkHCMlDquCaR9YO6mlMAUSFBk7r5KBzh22sZ
OceG+EWnNFmM/BeJzNwVnT4RFfxcMWa+qF9gmzD1U+mUgEj2pG6SxihtzZR7m7zq
pQ/s0NOKkG4RrOzp9OU5CG4k/PIisqFhI1Ur/XNRTj14r2ALOeE1wdo9p9i9ZPJI
cCs27dSkiFbX8YzwjRQspbK4ey8j3MydN/beud0n11NcfFTPknspM3uHAZHXd0fc
AzmAPvX7A4rDmuZM5CXPod4nKqwHhRKVrO83KH3iny7jL7DRe8s9nBMAiP9V3Ixs
3yThssZ4WUW0XMTJEAAYBfJkp+VkmvXQlRCKYAN3BAHbt74ke18DX9DHpkbwasIR
Sgzweq+UdqEBi7Xw7roEo+1ad3r1CRg02IKBmhn/QWsyXZbTlWV97Bye8KBBvJGQ
sx3RQ+IXkWXY/R9DVBxKoTqROPt4S+vk2YHOGp97H5Cto69lde5V3GNKfSzInj09
6Xuk48uVl+RpU9aE9QkKPQQK8weN6xxxu7oF6KovaelZnlduX2cpAZoI69hHOeXE
m3tJliuoFZXH2BOyFoKKzcJbNF1HWIYfSYVR1pSIeSRoUTT+AzbxbX945c54qC4S
aLrc2a1YRMVwhEJ3n3LWj0XqeSgJByCzEfrnQdWDU6T0QtBL9YRv1Ol4DAvFb2gE
Lq2clUUMFl8PS8tnUtS07Kjtjf0Czas9ako+osFsx0IyjM//aCGja7QMKEKXXmkh
Co/9vXBNtgpT7lOhq8JqPBVE5akr5B2gZPnv9sKjmj5+9+wNO6pofLOiTwAkgQiZ
IjipQZjkSx9wl7J6B/t81sTKWcCoX3ih67DKH+KmxlNDLSlU4mA8JCVrtghYARhW
FHENiW6Gnj3Nkh8S8pGaDqY66rztlDPAKt+pHP0Y7LbC07xKcrYQfenul6fYFBSo
cEnb55Fv6LQ112P6V4o4nNqwOVgnq98gMVvb9lU1I/8WwXsZKLmfBb2rhF7NzFUP
jggGNyxNXU9fJOCw/BbJE7iODaHpeGzmqxXzDEt1uT9Pa7anLCO5LGYtLLyOFEge
ljFgtzcWSb0E7HqowXUG6zuwzX4zLKpguBHYhTV0OF/13iYey3kUQFlczZ9S4n37
xYRBKquWc6X7ennvjdcWtB8X6FIyCa3a5HbtpYSZHdDu8eIeNsGJfoZj+P2C1Pc9
LU8dQfX+UeYZXL4qCxJQoEWz7+pAaGoqcqRdLPD4pmx6d59W5hBLv++kkS5qSUSx
Y89o9z5b8IeZkDG0e5qKvIE2/0x3S+tFGqyVVUz7ZEYt+skmLJJB+3sE0zgf/Q5D
PHlM13RFz7Qz/H5XaFCtGtI3259TEoBolFq17HzqBVjahM5VVQa4WSNBG2AG+9/9
EbGLkx4eX5T5iCqmfeUCsjuMPtPuMuT0Q6/jo0dCWPL7L2sm/SH9YFP/IHGCdyaE
82ckH3n17jHheyU69giWS4m2X5K4HO6IMd8Mii3vWHH1a8Ry0i0DCI46du00iRm3
QRncV1DpSxP53NvClijaSCPpcFjtEJMG214KJasDfOqJRMJKk9bHOxRHe1oDbu+u
wMcFZb8C9p74ajCjPeg3Ve9Mz0gvPmlc5vnvEkv/CKd06XdHFOsXgP2CH6DCxWO+
Buxct7UUCNPvc0RVrD/iSq2Trrcl9ZqFFZye8fUA0OIEnMiX6D6kn+K5z1KVkUMw
qou7K4QmvSnokXvHNPp/410IVJl769m5DlbKa3T2SCgM3SYpDjltcgu2h2mWWfg7
0K3dwSucVrbYLeJtgkN2J+ArxpIlEcyEYIQFeZF/UM4dAUiXs7lpNNEK4t4wzi1e
LAJHgsfVuFZcuO7g46ac4MgfVdKKM1hP3VEDQW7JOwWVGs2+E/FlxUQxphPfUdFP
KBx17/ZXl4gDNqdt91VYqtdXAV+LiKrIrnrwjwi1R49Msdv6mcNlRfVDRgl2S2lC
8orfwWp5qU502QwtddrDy2SHiddDCXDctcG8/HM9tUZ0rockfPDxZk9G+oizOv0+
Wpe2ioyjEnlzERvLOPEj7MOf66oXvNdYgvlLGJc0nD+v6ue7LjbmryIJWqmTeq5Y
8T+6BCp7eg21ylvIhwNwSy4ju2pb0ZVFwbfDWO+WuSzaA912FQ1/wqO/3R+rm7D+
yM1gsfKdgOjfRWIx8JGUeV0mW0f0Z/c1NeCoGJ0UnP3Uv3x/fp1LAJs0FZGvU5hj
VvD7X9VeHO34mh0jwix4pZrqTdHdoZCkWtxCtsZMNDs5UmJEodVRjv0bWLR9wfAp
R4uDWB07JYIpR0Uwtxqt3M8oJ36dv6ltMiF3cuxMdKsEHwBGQ7bXr6FA/JV9o5sq
w3VI62LfjtkIiSgdBBgEy6lGLHVUe+rKBm4sLaNcqnEBZpHzcxZRQKbOzen+sZ3a
RZCPYy7b6LJRz87FjxdpTDnAD8IXVjdgFtaafUw78536oQC3P+Kq1lur4lUBAV8l
zrneGyQx855E5S83mSlMA8RwvLeR3+ZKGYHhPh4FbmOgBMVIlHTF6B9IMyROqPkL
A4yh0aborLfRkfekZdg4MYgh8ZCc+ezLUUEDFWwzeGKntKNXzMctj+uvdOcPG6be
T5ETlkPfgVcHBQgPqhX1HkB78VdSCEKqp6aXcC1kLRb5LrKKux/thSDHS2KCFITR
Mwc/z2+eZoiqeDJBYJxz3G280z9h3Gt8JRyzFxaviz6izdGQIYjmKA1QkvOYmYwO
ruxHakpdwsOs4+QGX3bs86LN+JMsvz7QdDPdMcLXYZC2HKanwBzsn9DNj/i4uu+I
Q9YofjaZNH87c2Si2ntvFDVFK90O11lyTF+y2t0DKrA95kGNuXT9/WijKseK8aCy
A2BjWneikvOvn/w6UFtGs7MUqqcmZm9tUWek5gu1sXmVP91MM8DePkbJIedfpJbF
VqWLfWuUn5u8FqVrFnPvIcQt2pCkwfrzBxyksuq3c3i22lLdCt9sDG+J/o8gEre5
+8sKO9xB3bBCmmvbZP+k5YPnCtgeepXWYwExHh4AYuPEKWCi6txzLCm/WlZfHT3t
2UpyC0/Y9nEjKf+6gIos4gt/GaI3zZow198oBRstKRlpJCqjrbyFe90ZHIpqBPde
JDI4HpdzE4fIIFaxaEPNo1SG+vzpWCW3/0fX+Dfzs1qJTvRbsmvnsyG6J6vowyYO
jIspAMv8Hv2grx0sQEQ/8CeX1uCuPAwykkoRhAsu7H6+HxPlwQ5fLO7mBJ0DeOWL
pbrsuJ3bClH0OJaPWIbf2gVtn3R4y3JDnCWjrfCAOq1S4EnotRZMmSv672naHBCs
m6GQUOMqlHLVjfoPYUUhKk7Il7JMxOSr+uLvVRLVFUe7sDqc5JoQOGh/XNv5Wscj
QpEfHo8LgEuakg6sMFcDWoSNtf00BhywF/o+GaDDUb7uFtrOUON/Zu7uAWwVlLyd
uB0fXDTneiFCh/Hl4x0+oGFjd1aXTCwAQKZqDIent2PmX47P+vkPylLPFqZAkRxC
pHu0mxWOU8MrDjJ+aLxLze2N0UpbxC0U6LJO/9WkUkXMhE6wgoh5Ed7grbI/evwT
BkjFJQAYSypsbPaM110O7tyJebpgZFh/iAHJzsWhrZgosiA7QQy5aM6UFz28w++o
NVweXWVWX9HK/wM6TD6PrOEFkDfEypeWej+pGVaDxoLCv5SFkWO5S+iybpgJqAEt
IE/t5s+6q0+14LQs5Vs3fPMD5Od6lG4Z/9blbPNAwVxpBgT9YagItF6bjEmBLiLG
GuSAF+JDPYtztcLZR+2qn04TVYoGcAn+StS0FpDLbXRSGhSRFmJaqygILYgP9bbh
Er7m45OIy/cTAOecj2+ayuFAXVTvDxvZr382MOJk2M7IDwPUfEyPGalMiAYJb+0g
N0DtpUb9dt03EjiAGYZvHzAaS785m60zty3d3dUMP0Z1muKOnvHJjoePjqIdwSzQ
kp+hER+LbWA/MqjYaCNw4R0vss3up4YUoGMuWHKjiU9YOZAe0nItM4Mzu8CBqVuC
ltJz8nVnHN3+c4HUBybbxmQgmPDhTnmT1UxXYlZYzQ/t6IHXnQzSNfpIqsW0YwoA
Qv+cOmKH9asX5RUlv39g0YwlRLIKVte6mU88U4GM0x6znVbSkxjbbSy3Kp8837+m
akaR3yLnzvJcqm7ITF+1vqMEoEbm8HVKWHJSPVvN2ijP69f/pV2vkDrAmu9ZVuqR
11HpqNrHNZGowqukVExhhbsjM/45Vs8eVweq9cRwo8Z0E773m4GrzdC28ID+gBcw
IhMCxg9wZ3OpksFQ6zbvcVzhS/+T3vhrNyYqjsHV/5PYJt/ogmd3A4EaSAzfQ/Cw
708HGlF7nWnwAhq5opK1sAC3oXuUQAIBiPnyeszOy4tXM2acWPAJkCqTNF1JU9Vn
6Y5/AmNEcQtl1ufCZ8iolmhWxkHH1CMpSc9USPL8mJzd30eeH3FKsiS6CzyekoYL
Yc8xGrETXlyXbdcun+yk6roBGIJHZ2KkTWOwvfyWKY+jmoaOYYpTq/3wOgCcE09Z
m4fs7bIpxZ+L3vHDA8Hui0paXfqXnha5AWALjFMp0t1XbUVshgyO508wyXXsbQtJ
nvoUgsjgjJNtIimsvXldwV/XHUuYRTv8Ea3cJw+qABWpf2eWZfEc7JZcjuPCu0uS
l2u/Jubte33lYWo2Irxpg5E8COH1rR+ZAKwCpKLLLUVVOEcpucIFkjmGEhzgxUR/
Sl/r0iSxXfRBzYHNtWsj4Rukrux1c5+df0lvgKGRR/HTdP/dxjkqtdAwE87UdXdl
cL63DjBSzpapaat7MEwePWhUPYR9QEDJnTTF+qEMfScWAS+5c/a9kjyHeGjsIgI9
NC1m5cwhrvFBJWx1lS/KdM3oOyphaXh/ieZZOPFzeWVy0CWEnQICn0Mhd80X3Qhk
k8K4gh61XbTyfUPf6MVPiLsZQnB9MO/o5ILqQhyP1Sl8p/Junnyeq8xFmgX5A3IJ
kcqpjCn2xqJKudM0InMb4QbuRnvxf+QAPa0gKI4MrDlp6HLGks4RAZ+SNwMTFgTV
0WCZAX8GcxN85ze53MGE+Pt56QLAMuoBrx3vFGnMhSbn1guyxAQ+y/f+oykrsuZ9
XF9NkYEs9d8+AfVXcRRVCZbSihkGN+gtU8Fmc50Hi8NYYTooOYRRn7Cvbulimuon
wjbwGDk1e2LLmT4odgqIOkqyrkNN+xmlToBoSgZdr/mzltWC91gFGUPpiiyIezM5
/TwlPqmxW+Y7gZww+4lVNTkShruAe+a1hysV+cNjthrXHpzgVb0au5clEWAUSGHk
zgvFHd5kVrULHOLulgRlB37xo5F5Nnl3bX7TUx3oNEDAqiPOlXP96buO0lSShxSf
uWi0HaqSsJDSD3rgAE1pjVOh9KeiYI5uN04iEDgV2UXcdaud6hl1s0K/B3tHddIw
2rBQZbEamm1XfegyMu+1esF6dHhUkMEeiVtnVtAP9FDaVzEVEpbKHl1kA3dYqZbm
PTZ+VrZLm91PvsOQWXCIf05oWbfMU1Bi7jYm+hC7H4JUsd6nG1BqMk8OxCJaB38Z
+hVfOA02bsbT8SsDrEgw7o5bUD7KjS27owQcsjpaigt9elRwqjCDjr0QPJjH2Ei5
4SkUROFpevpJzH0ysXFYNY0c+eMTzZMRpzJgT+vNRJp5nWZCDbUTAqRW1kIsQg8l
7p35s+9wtnDaOsNX86Bo8JCUVEGPOTpNUg46K4LznDKon2fXEzAoHg5r8U6S2HXJ
3lLvp4cYWpxDHJgoo/yZ+Bgbg5fCtSxc4UrE+GwB7ZB5BH6P8dsBG4Q0mX/IE2XX
BLO2IaRRu3YbT/T0fHU4OoaUveiq9+vWFBqiDY0kVivvKNK4U30Uh6BNR71c7fJO
860xumBh3VcwwuKO90ubn00iDzNBMliWV9xA2bXFgRL7TkBMvT2BHH37TAP54+/Z
o5WHMoOD48ILUntfT2mfMOTXSSg9gnJOpO7ULaIsqDl2SYBV9FTHONrPzKSI6DxB
0dJMDAOPhqogw9K7pSHx5Lnn5vXlDO4AC9tskocorBFoVoCf5m8Jm1XLsx37Curn
3wg3dNGxcaI+rP3gh8RR/rH+odtkTKK/c7y/PeV4E/VR4Ny1iM13+shhvHp8ME4c
kCsbfOaVu+miLZ0RiqKdsXdjMQ8P35n5EHRagyTBDCt23ht0I2LSLdLk4DjlpBH+
lrXQzWLruGyBJ6GbjMNwuEnemAY+9ggWQ9My5y2cT+o89INeMBksUgxC4yOXI9wC
hrO+Nf+OYyMHMQ2BstAD4F0CPUKAggMNBvt9iJPgSjkYIgjMblBQQinpQTsJfsHD
oL9RsqAPiPAOgmT04q6oxbV+t1KRmM/fD+NZZS61UjpoN2Tn62sRL6Utq72TkExH
4M0dkdCS67CPcp2vB6s320v6ex6tAmYbAwl1huRaFD8k3PRdjmU4oZ/+YAeVrwXT
vtJWeacu2nzi8Q5TrjoEj/AlKQHaNoU+xRMUOpEDPPPfZmWfEzq9ONhudFJNJZ3L
ug4yeCNtLer75bRanjFOtA6IrZ6zONE44HPIyua1qzFK4iQQv6U4XjiLrs2z45cp
4/0VQuUOkbJM9sm9g35aLWH/7A0CbdV4a3sludeMZUrPTFJONp8hIriyWitknX55
g3Md58DRJrpVCYoLydImE3yWKIYI+6gFhUun9blq12RzxN+laus3sQ+T31o08QtJ
Qu0Xu2mBxcbG8vEmlUYo0uxwjlTAWQGsNwhY719sksYVO90nCiQ59ODFAlaAxm0r
7TWBVWH9zn7n8X9Wf6sRtpb1hr4uwEBLtB7pczWkAXQ/R9ocjzQOCjmtt9+uzXJt
Xb/HfjNjRrQjgIfnKiSgzzPjORufgw0zuIsovzl8TGVYc4l7Nooj+jKAc4a1y9Nw
yM1GzvIk+Glwoj4Ui1LxZpSU7HaHyYDMW/mGkMhL65UpiS2W/Be8cGrwgNcpK+Rt
EwjMpjHn31Ilpqi/RwXCoFFsXZzko1sUrvY+ypmvNr4n/kPYYubEFXw/MkTEJZYG
CUFCHOxqeFkq3q2dvaeGrBmuEW3P9h8gIa1/Csx2xS8gDq70wCxtexYWQ490HeLx
0KEmKBMFOB3p1i7m3BX0iQ01Jqk8IGo3L5qFrE/4szE4PuD0gT+huJJuSRtdd8E9
CuS8VGshwQfxnVemaTv8c3qKAyQuiBlponw047PKb8P40gV8W3j5/yw2Mfgt81D+
5Hhzb0AEarNaVpUUxlsT6GXyjnzeqckI2hugVINE5rasbLfkD5SiYFwpnAppbSkR
UTQCB8iL8G3FfZfF1AFD0fmbQQDmT9mdMoc3yY97xmu4hJNl12CxIScVsxjtCNlG
kZbuyPM1aUNJopLtTkxM1E5iEflxIHkV6CLzCaXRsvFpDlDnoDnBXpeVpbAaYdvj
RTP63uyDJtlZvpC8oI2VYAFObzeowz8qTX4kGlGOkS1O4lq/FipOyiQiYGwdYHX+
kjoTf7aepFE+HXWYC+Ndp27xAeaXIDfZp+bcS0e4srLqnP/yiX1XuZGw4tAJ0zMQ
3vRoSb1SuwqAzyDUwo88qCrenPknhpGh/5FrM8u+diNmLVbFI21sKHubRigXPBS6
zFcmhlcvjaWPrfXF9kUtrQNAvQuR1hLFqjb24O7Z3afLsqDRjWOqqlkW+ts/hqmK
xgEIC+zs2tJwlqQ6muiEfMhrsrGtlNVTQ2S7TRcsVdzwcG48xERP0djmS3og5F2J
2kbhKIbHo4WvTdgZYw/eFv21wMtd24k5/IW1INXkee7FHmn9stIfxzI2O2bTmhFB
R/JWPlgqPG/BUhue4fhQr51T0xkTlR4qTiD23djtwL0txEC5PkkoxFqobg/CIM88
OPqVkIixY2Wn7RkbUNxzMQ6qT904HmIFKugIKqBfyHH5cpdJ9rlGfJiO0YghCO/2
OwHxIyPu0CWpjgXVQC4Qzh1VikEdsWgIPACeAJeo/k5oBIoxEozPZeQWgGZnZ7ZS
58Im67ayCpAoXFQKG74pYqviLVRJ/EIqS2RPGEnKcckVfQW32m3kXTN6OFcGhLnK
ZI/Ue3LJZE0WIgceLIFDt58S42sZBFBKoCLCg2jPX+1nkHNi3P1JCtwLjftEPVeu
ZLUC0SQYQhQWk7AyoTV9j59OIhOOcXU6RKAbRd5BI5nTuErvWYEFVRsOo0UIKnu0
fhua00yMasggoV5fWx4X2hvYsqB+qnlNEmx8SD8NegVXz5REY0YCySvRO8Ykidzk
PaxYTcIP5P7HkgF7kMxBc+dUJCxUdV3u+erKLOenE3iC7wja2a1FtNbzfRuNUEDj
0Zrt5ZrgZhVJB3A2ZAXMy4yzLijsStcdXvLm6wuXYJb/JwCMEeFpnk1xoEnecJnJ
GDqOrXfivw7FTRLhNyTvBssxpvmfPGqA5kwrAjFn8WXYeq3lTl7M2zL3Nib4WAO4
s394ViceHwNsmwxyKJVVpSKcGq1ko7m278V50JwOOr0IQRd5+6n1dvgZGKiZtlXn
m+msA57L2faCoVebMfZSvB+oWy2718+hWHQZgsWwjKGQBV/xh+OYh9SITuPArfZO
QnlnXDDmDC4P+/GuKinKI9/uUuyGFHs9aQB9qzYHpYBMfUXlb13zdO+2+QHaMnPu
gyr065BzXIi3wRUJXYSJIq3TQx/9wEzihxwdkEVRHz5YOim2Uy5XVdA1tuKjROs4
TcF9A5Wag36J9vtF8fAI+Gavf8waUGDed7A7zBKTvi5VcVrstk7kX11C4hN3447n
AxchzNDToZ24uh0T3+3Ki1w/BFJ5jah5R+bxkdfmdzhlfAj1FKg5xHaRfaPt1yM9
Qsp3zZdy+hdLwT3dpU+HSsLYMIY2lZkfnZcbbx0hEna1rp3eV03VgiomWjzX41mE
7b8Ea2qMO+KAd/NmZDjCsku3Fq6HrSckba7kuaoKQoT5AmfCblZFyz35Jk4Ls2/C
5LJa+Y3QAU7KZOHy8FgAVZZoHhXM+oPzlWjIU3DPhbYADD8hp8G6A83GGXzBkF4N
9+fNMC/skr1sAjCY/skEdFXgu6cnnvFZLs6m38icLzRqhH0wm0rqiS2liTyitfTG
8+0sBei93IUAsNUUouUDqgvKSttNGjITdzdTykWLxfy5WZrAh6O4fGhpkhTveLMG
PqE1KRCDB9e3BkUHmBaq8TxJRVKlik5zrT89Hy5X8xP/UDTCBucw7yfW1IxhwRwS
yY4I7sOEvdXS5iflGX7uHhXByhUefLEL9NLSwRaDb9PyssPVvR4o2XL02pSgA1YK
gttao5Prtk98Xg9VqmJMsH07swm98EA2KWrOKv8lMTVK7kzVaWDpTf1wZ75vbW+s
+EcIIRw2O8UsGyhhz86bJbJbsJNtAo9iv2rZjSbFaMVT801MTZNJjxpzXe4xC7FM
Li4Ubd4f6JaLCyDA4PrktredqbdKAnbJvwcD/lzleTgvVgZ+UIcYRAo6tXXgnTWT
uEPUxQ5W3N8QcpuANd6ZkY3u8wKd1y1PIwrwFtoSh1GYE2rkmnd80/6Worjd0+2C
QDGyRH+1g5QKcIgTIurYqI6cGa7xMZGFZjbNYCQIZ/uiRTYVgwaCL18IM4VZPr0N
qd4fN0Peypo+VdCKgOUUGVxGd/A9fhUyAjFofWXOlZ7oGzs8FWamvPtRCWkXqGa5
VJAXU34Z13/jxXudDl0rqrnvxDf3YaR93txiwCcsXisD7G5GlaI9E7IZAiJHp5LL
3HMjzBRyxIzZJaZPRAEUpEHxUHeyIxB/mnaNfscYNA1NTwpdbzQN9uNt8w4kN8bo
ljZWepEFwi9aY7sUuwpSVp33grglZHw9cjjS+4guqz6Qz+3iUT5NS8PoEpKL0284
ILSqLWpkZL3d4dvZW/kaZb5pKzbdv2+qF8yozDElb7+3erxTLZmxvXRVeaq/lGxU
JIbfGVcCqbL3S8RoHFpFH4DC+semqZfgiV9zCwI2H/xfncR6Dq/oQzMVJLU3L1xl
VaXJEaIi+J38xqrMxvOFxwICILrgvd9Ws56fiRuL950WTDTXEbrMDZd3cL4mlV6C
GLKNOto4TDZoMwrcQ4qcC7oja6n22yw+LlV9W1A15h/3PD1IZbrg3WDr5yYnsMHv
xRZ9EBLlCiG8KP0JC+MvazktWqt8W3Fs5ovOLXVI+YzuprX0Bf3j3Cikemors/W7
lMKJSydPQy/7wtB1LiHMpmAC2Pg8YbecJh/wgQR+10wx8qCyFtQa0sfKHq7SCOKu
JIg1bnmMmk1Bqk2WfX4UIf7TAwEkCcYWSw7fpfQRpJ0uegHsqGQc3/D1+aEVlQnT
LQ4Avve6MGBmIYydLuDysaENggZ/2N/2i4ak9JbXwB39xbWaJaHsyn8uJ37m3/Sw
WeLY6GZm++8zGRirTvGeo33BMp/A20gqsed42qvYw+iXqGy66sta985PO9itL8v6
RNb6Uyb5oKIUITYUEdQ+9xeqZ1Frdn+Se8fk3KkK7ndBTRG0rfCPu7QgW8TQjwMg
KUlfTo+FrgLxE9BRQ0v0teubR+CB/Xqyn7GBmz0ZNracfZahKcCbnVUdOZRXcc4b
35feIvnVjxVu6bUxGalCvTXJP8aRrUW/ZeB6h0Wd/FpY5Ej7YaLBIbpsJMNfc6I/
TcI1CxwFWn+vXvu0t2hf7mvEUYkFNtiyr2362AHDq05AGyfAyANmfl6H3UwMNuiH
I6l93Q/rtfBEIO5heHrk4kAuP3e0qCUJTnYujoXj/J4KjhJ84M/4w2WzNyO6jIXz
XcAo+1jszUQ+nFimXto9pYqr+jCqjmR6X4+NrZRVilMjlGAzx7kojDiNWwr/UtMy
/gh7CRl2GiU6anMNuRMy75KrKl14M/7KNcdL2Ue++HkbpX//YF8Llr51Qayk/dQm
rTy5LKe+zxo4jZYJF9Oa1qOm/L+WC2rKE2rUoH0FOVmueJ4OuoiWvvdy4tX/uz9R
cfA6GIs4bBBwO2dJITVjtGayAda3LhQeCtfc4nQAqRTuc0tGJHAAZjfsrnt/w5hQ
qDxW/jq8zAyVlfs0Fsph/GPNldD78dvYuqHa73xnU4WED/+1asTZpeK49agG+7Z8
J+sQ7UmhXHKiG+Wae9x1YUWdVqpjg+IYlGNlij6gVtK+YXUaLnqxOmDWhQAgJuf0
muHzFeTogDm0o+TapqxU4d5OwBxLxnS0WVdxmno8S4LGogESzzuLdgX7BGcPpziK
aCzUkvqXg4r4G4qBtuDfxkOsOr7WTqQCmoaVN0pnxF7bxYRGahSf2V64Esj+83jc
WAUrqGD4DHcmsYWyqfpjSiMGibRh/e6gcYUBH/iZTy8jhoma8OzCarOamf7XKcXf
MldSvo2xuuXRSJivLmNQyp9354TVDd3HYJVczhNOqxsQf+3qoZEoE6ma/ofi2x0P
W7FdqTkllVKQW13hW1a3ZZyFh6XKkLSokCk7B6SNLcAXdmY3+koon3Fw5dFszBtj
jVx+qNL5KsjPaeCGKitDMCGVkzyaJmtWObfhXMWaIN4d9AM828PSM2On9r/SJ5//
qJrRjoC9H4xif9rrc6w8mEHnKI6RQXNzTxAKoEc2TFMciQz5VFoodoXXW2p//eSo
IaML7RjUyG9JZx/rHpVK5X5V8TticXtQWwiPrZ8MmtKkoBlgfQql6asCVlBzy0+M
BZG15SUM3hjaszYgq8IH8LZbQTg6nzG31ZvAej5fhgv28uTICNuh5RFW17+67GA6
W0AT2BnistB1XIgXjkF2N7srK/BIjTD4yfbr23OOoZj9fBrj1qCa0ILsSU2My9wo
cMyb24Hv11X2divojgQNJI72lYVY5+aacBAehAu6tmCoIqact5ATiiJI7Mwe1NAe
oviGBnk6bxFVFJ4bKWG4O+s29RmPmrG9t8S82U9LmOeDAl/Y5filLIGH6KI8dUDJ
Jn4FOJzgwV659jnluD9a/IaCraoSsJOeQrf8WwrYT6zNWD2u9sIOGL/F+BfTbGRA
toQKNgZQpahnKJMC3SONiGLULjYPwa1VJwqJ4jhVhkHfYej9qn8zVUWDjNuUtrht
XLKlmSchPcOQ8bfyeVMUd0XCwv854RW6qB1hLdUp8ur/sFsrkNuCGMEfiHeDDPDH
+nDJ8qb4+XU9H0ejXvrRLtRp4ybzO/rWOr6sRsgNMH7cDujyGKWhPzUSC3izt3tK
Kt3DlPksQY/VdcFAiyXZ7hR1xnZbbve1zKDSw0z1rA5udrwWdTKfu0odfOy1bEn5
qhFx3Jm6huIwh80sCMr1R+F5qenFxkz5/2S5gunYBMOpbYBr2xn+gha94jpHdKIB
bRO24qRLXwt+9E9mUF45CrYdZA8aLSuZo4dzuV0HEH8EK9AjxMgmyXZg+Q/7RVb1
BRmmC5BxNb5mH1wd+MVkFwbU8lh8a34wNIvSAPgL0k75LFDktlWgYT2+Uv+1Qp0Q
CVcZiu3DhNK/OGlJ4d/3h4tzQBXAc5k3nMGCjUzS6Mmue8Xv6KrL9A7ziScoVvr8
n5MBlQcPIVPxs57X003zNrCTNb7jlGKltDTP1Np+wlDSpxrTbVQ9JLLxArwi17ti
+aUlc4v9lDQKegSOm0ZcTNqiaTpiVmIt2qlxDYEExRMR+2Zeor20fiPSw4w/WvoR
K/OI0Rp7oWwBxck0++yQcL6Z0Z8IKrBCB0+JbSquCjJczcVYKCi4PCrEnHB5P/hY
HRYlQ+Vehtp7ktvL6Fyx8/0Ehl0tVHUmKJNfB53MFf+qQDVycgHhCJbYOJfpY92G
dK0hSGiatGIZKFYm0yTLi8qSTrz/1iMLUvDTOCJhrSR3E7XRno2Ku5a/Vzq4IjBK
rj0xjgI0LUf7UjG/IkId4uAXstsiPo0V4QlzMIwXKHweEC56tAt8BCpGeFN/HuJl
/gA2MQiVQHjTFBvBQOfM0NAQjyteqxzqOJwXXEgBL6W0spJ3Zlv7GLhKTop+fZxd
np5yPlHceshNQo13KI8fqFP2fdGCoH3vbfNgkpAkIM8FLBctvheooGxvBFJgRgsY
mupac5TZB6/cTZ5bs9QogwBc+pRSjJ/efsNZ+ew7Uy+0vvwdcMJHnMdJTazDYzfO
HSHwliow4XHaGD8Ed4ZpkYg+yeCemvTIASVYuE1hSAahaF5pcTJzREx9XlsmMZ98
PNr6kWimiqW4587IM2cd5Fn1jdA4oDSqernln1tH/FeLkLvCCYYiuc/plRZq+JsF
DXn4dWyiIe54stS5B9iHmcI2ry3grQmAsAETmnOkfQsyuRYt3vJRo1EPIl5/g+zV
Tbq69wQroJPOj5AgOJBbSI9AE/RepolhbTu1swU8Z5JH4xOhHZRfbrLy50cu65qy
JepCHQIPN3HUlqIiloNEghaxSSwnlyC48EXCuRgeNjN7ynX5Ep8iaqN8Yx4ZWJoz
m15dWPbldV55xBnOqUxO7OevIG8YmFsBXioDN2UugxiqCcd7p/GTxuY/W25WAtDW
bC4Brx9VDqSXuw0/p1cp+dDlSuFeHoGMOde/um9VWa1SAigwL1Ww+ntDu8mpFIBx
NZCFUxJRnn8FDTYzQ9aKzzjNxAY8sgH8tIEtsOmYgVVbeQzFyKOOPl0dPN5Uemd2
ECQvZRU3zsAxS36ZZ+tIZVwv/CJJBqnHKxFbWbxipMpuK+40TWFjZioS4wKU+aI5
Fu0cVHJP75ynd4ccszezp52PKD5IFcBHg1lQG9roDRPsCwxgegM2nex+h9HRectT
qym9Ul2eI3rI+fKGSm7fvpl5MmJIo/D06r1JTf68/Ubd/TLbvyO3xGR7obC/Ovj2
UGTr3WPRE6LqUyOY6Uys4RDCkQx8Zxl9l7cRBPH1VL+REP83H6alET70tVu3PGYI
7dggsmsnSQLeM/9LTc3N5iLsJ1OdQJv+sid+J/0o9B1olfTrb5N7SMABKRZbVA48
IIMfINa40CnQPYedqUEYnjyqDMN0F+aANGUrt3yGpiKVYJq0koDA4s27BeFmP7uM
+dZKPCAUpLHJJeb2pmB+bgIgEiXcbWGU7TyNLyasetxPbHSmpKMMX3S5lUdps7C9
U6fdj+hIKkQhwOcm55+BayjbTiMVYI4CiIX638qi+wMEYlrcBP7V2i2cREEEgYVm
P27E7GosJ0D8hz7p80Kksc1Smu0ELOy3SsGAYgSKRy70DPuaS1gx8xB+oshZ8iXM
yJ/mWlMuvecAyWU1TTWA/yBOl6rzpWGpSIdQs+cWFaxQhOdTtqQG3HLF+szUXvq+
78oN5Iut6hUf//eSCheEtrAzhZwLDqiABCzBY1AwDEPpSNVQMEY2700xKA6jxEld
bTDFK4p/0cByoQP7SvGz7qb7dnz3uuyEHBTNzJvwOmOrGmY1u068mIQyhycYyvgV
el8UOKsUg+Pvb26jel4uWb2B74tRvOJW4kg6pegE+vLwkhxJvMO0L3GuBG6E/rXn
UTzVu+tgEfcn9/eYSXuuDaUfMqwzRqOAoMDyFS9EBRJLnsDiGU32ahV8S0JNR5Oa
TTYovG5Rp9e4/X0OAz4qgPDo8VRBEEzQTVH+2fmCT2gwEE5x5tCsWOq3t4jkbxib
WLEwidjetAsJ2vAuyh3o09/Cn1qLAkmQh6wiByeBbI/iEzipGvsgEvvYAIB0C7kB
tKpAHbJHAatK2fAsQ0IiAh2Wi10Monn+z7LQzzoU5hFjv8ZaB2azldelvTEuefAb
be+oG8jc24NOg0+TGKKV+uBZpQEHWiezrt7dQk7IPBBYMr1Qh9NLyuox1O5kIIWm
l+Kz3qf854ZrpQJT88QnkNrjX6db1GrHMJcjejBbGe93/2yk54PZTttgaha/SfxZ
3zzfSXczrL0WHidGo0i1zNTFi6Ok5KmyEUNwDEX+JrAMlWlM3d9kBtcLpyPIvdlv
EBkKR5SGBdm4JuEUm5c+2dgbm4iI4R8NqpoazKtIiNIDCVtNaAg223hu+4L/WTFa
nE2Y1T3sUNbx+9qWhv30Z7h36MKeNyAd6cNqoy9spm6G9QAi9qiavT+Php1APTay
W8WcsDyGxKJrfnT7u6ZJ1SSYJXyc8jfzSMl2hUS0z4GBQdDXl3w5+WpOQZsT2NUA
NfEFjyvAt6TPGY811Cb2TSrSoQMOR77rGEsa7rMiRLqne68uIq8JGesdrE6TCPRe
zmTKJVHfNUKkGPx0zMvR0OtBag4pM8c4mUKl+qjWSIH8A961deg98yw0bpUKv5Y7
WjpkVeEf/nUwTXCwmo8U89VhQm1MAYkVyFHfRaXf462IrlgDgcixjrrUvVeIKUzu
uHVncKBwG1wFFmjyUSgiIq9GqDwlfiJcIQiDdNl1MAckPrTkQuRqGcWlDHhILZRG
JUCaoxzYfmZZQtlKOZ24nH/JcwdNy8Dr14aDds/Rp1357DlvECxDuJ4N9/J55DjN
dVvdS5GugvX1QF/1KJOiG1pldPFi8fDhbzDD4jddmGaZ7IHbHZYWS2JWDje7lreG
cN4Qunyddsv9w/Jj9G608T7BV3uPtPg+DE5aiK2Lx+k3Fe0/bnDT87HxZwZbcEtu
rM7f79Bxzik7UNCClG9AJ38Sv1BHu7aCDgUf4EKB//NMFIA9oUHXk8UFeCSKjBXz
jTHHQGJW+I3QK9Ks2Auh5m9RNWVrLyRbB7U+WHZdck+yjq3ji8qc1vn9TgXryZfv
a81SzEWFnoxlddZoa91Yq6CWvKGZoP2VOlIYENewnz3V6qbHlIcSvrtthtH79Gvp
C3HEURZVLgo2rKpjkU31H7OwnQpIaD0/jMlV5sEaxgtjngyOLaeEqmFp6pWBPeON
vhUbYq7uY4bqyerdAui6Jx+yjyVqG2tvrr7sPFJcGCjco2uOLsbNVqIulSOMWva6
7SiE3vkNaiJhpqaX0LVDIYYDP2hqhsgfmy7T+a/pXVBm1FJh2tLXBmYbVUYibxmb
bOTNOfrATgj4VT7F2d3AU4/zEIrwW4mz7sMKkHbDKJLbjjfV9sn4WV+NgrKqBUL3
W03NRa8p9sI0q6VRx591yaejS9a5BlIXzRB+msitInjmjioVFDv7jZ/cKUvCVLB7
NGi1yDduPzfuNO3Cr/MoC3SW/ikX3lexgyFNXqVneqnWp0kW5CYaHfJd92kaAIkK
xi7WQ/x5xFSD6v8h9hn6xMdX+CQQD0/77IzHHKYc0vT3JqZnfMHcJ4p75+19zh9A
rt4DGfQTnUWCI7Ge7T4P4HhYJZzs2TQQn6fsiCsAw2mGxWIwOySofdXrHp6DmSL1
X02KvFm/wPcL1VoUepousnTohsITIT9oEJhiiRF39ARibCMFCP2TFFnQ+jhD4bjp
KBhQxKytRcLw2zbzTr816yss5ny5a+UldiS1GFq8JV3nbHC950Z/UeAmjjJTUnga
fytBRCXZ2HGBejSlzqxap9Ej4CtvZTMyV4SGxFO6VcPatfd2PMyVqJjkavBLk2P8
F7sR47HTxxth1AtP91l6kKWnflePxEJKvQ9so320DgQi3etX9M38vrUQpeEJHE2o
ys0CSPoXOXJM+Wkj8HRkF1v3QP+dGELmIaFGqHmQ9P2docdMxaC1jQfBvfh6vvMt
yGAVYbjMeJcZZCmfNybY5kXJPv/viR2/a6sTV7VB1o9gPN+BbLE/UlK1uqOeQ9Df
LPBK1fySSbOOH6Co+wdBzU9MP0cBIObfZeC9TvWQxW7uerf9eXNZ3HnGMp7NRMSP
fhgL1QbvXkuducOOH/fx9zVAAOeO6YeCMEqyhaZMpdzkMaMPHbPup2LrWKFwugmf
7dO+f8DLcn+lY+c7+0x5yLWZIDJ9NVmmEluipxviudn2MmsNh+gA8xtCgvs831tF
iJ94SyBImHq2KKUm2EZAyw/qjV+4zsX1TnWxmIQ5u2XXQ8/Tp7yyjfNg+whs+2bA
n+mvwICYagv1Ulbvla83ltzyLnslBW6pnJLHg7r+BLtE2gkzyonsSZOVJlxdMQlD
DcG9MXz+K3fq+1bImcq3vJAu3EnHOYAiT7iLK/UFTuim90Fg2knyy0KCissQcdLS
UlL7DebQh/DoQcRtJO4eRpfRS0/qeJr5JOotp26bB+Su+7wlE6tFyaXczRAGb546
pmgK2doMywViTG3hMPgxPqL11Kfr2itawAg7t9bGq4fw/00QNr/pUhiN1lSSqZIl
Q3WpXZDUJe69OWJeTA53e7IWzhVLCqemtt0cGBF+jnbrVvO5/PSTH+BzXnL/8PMk
8uFtCC90n15CdOMY9bwExPUAB00A8ipedeRddKrQ771oJTePE96yVn6q7O9sydEo
xWF8+f+wVc9QKWMjmEJFvOB2xdYZq+rAuYe1Y+RJnlVuUPcaYPp4QGZjAzjPaH+j
PQCRFks1j8gqSLch5Pp1QEc+/Ia5ou1IRN7M2SwGFInf1UwLceug94I/O5/Va70e
tm7rJIIPK4VayseNoYyjoKCGojfpmDs4YInmWKWMocPdzQ1evRI+BcUsQfv12q3J
YzO9gbmjjyS4CX+f6Gw51wFFbp0LCxDmKJ3LnBUvf7H+kYhddEl3utq2STdkDYTH
PQDDBUBefHrzCSiPtxS+kXSktYoANknVWBUU/pP2PIU/CAss6G4heg6lP2VSSuok
bro73NWAvsXYuTLr0pwIeuL9yJYJ80xrnYQu9FtI3zcYce/W6Lz/gEj49SAExLC0
WpQqG04gBL7H58DgDc/tYKxmEYx/e2Ie9Vqk546L74WzV2A0kYfmigpqqq15pVKS
0pXdFZ05q3NZIPJK+v4sIly2mU7hW3mZsLW5aH2VksksBR6AEv+0Srcq2CQ6Ec7a
5jU5n4x/Y2O5d7wrfIESaeFpCU9ChFUskEbbp3woHfqx12vlHvfL0l7WG15swbzA
o1aCCA0X1BZCmMh80oYDCFCN17WKeeOot75ue74BcLdgbJWjQQlaiyjg7I/BYlLL
M24lzwQMhPbBgpD/cKhiAgu6aw3I7zQj4k3CKf5FERnXKIWy4hPz6sPc2lsdC5zx
IfzYGiUDtcawRHO0GHAIhFX6O1aJkWWu+buiinMMM7+FN68S0fxFjHT+3bj4+ypH
0ZOKA6m2sz4O8Kcz/njUZGzkrUDxY81u7a906FUiORzw3hcwiyZgRjupp0bKE2/a
DZZHfrjej3hObStD4UcMGOLYvHpBCKxpLQgNRY28Gg8MHPI8F48tbC/aFi56OJGi
MkZhUaqbyNvsOKAvm9fkfIyLyyDPZ9QqqTV5aTt/qLuwYKi83o+mt6wfIlaXxHIw
zlujRTIoKzOK5mwGwq+UfKUrTc0oFD5ZppqdOYqojO/uI8/tKM/nBD+eycDtLof0
W5cBBm97oR0gVqHsrBHdr2ZmUQoMCUzK+pJZ66fEtQ40BCHvCe8E3mdJYMgQs46M
qVkh6C0QCWdVEFQnPfybp9aazV6pBIzADpEusPeCH+Ir+nvrDJGz1vVek2BD5UQK
S9H7S87iEO7itCND7GipQRCU+T6MVEAdxjStgL/MLq/Qn/uoqOAaC5xGET42O5kf
BH0i8+F/rgj84UwGwh2WkEw5Rxv4r9ffCpIuf1rT6wUZrCYBg43MdWw3Ugi/Z2Ms
Or0xfbSuWhciL0syM2R5fbWHYN6gcaZlQ63rmtj4oJmhbXKSDlYVDsZp+MefOJ7m
ErMLxpMYtrwLAM9udeFu1QRJbq7DuZ623jv2e9APK+W5b6ce39YfV8JP+e/sozrN
CXBY6YEwEkdfumSFxS1yWYqzGjYdRU1WjOx6edq03G6WIfNWB2iIAQDP/ut1d4xc
wRnjmr86U9hG1sulsqW1nz3KMcOhClNYLYGcmQUS1t9cmz8kfC6jdjNic8Vp7X5Y
HCruipKOjuOkBWd1Z7aOnDouED6b9atixoodjcBwiRMsSQENsI+ogdmPQGQ8SVzI
T23vFtoY8oPEKmiHuiV0HZSH/Aw8wfym4dC4KGqWnIsoGKapumppInhTAjxWs8X7
714oNEyPjRb+2hxklJvJ2zq4uoVQ9rUFSx70bs0shqWulo2RM8MpKpSgP4dxOWdi
RKKUxW2WrKPzDkdFRGY1xEvw4gNLJ9DUrPzGQ4Fij2sGb7i1PDegb23UbvJG2V55
pNSD6Wf2trPfWs2BRc8xVDpb1xIi1YV1rKzZcQ1DnxBAKVyJYzp98RfvQLn1WC3u
CFYz1I6+YtiOlypnEcn6GMvflBIK2drE/quq5Qf6v5BOTAaACL02wFqs4m5+8LG8
HVfa1pAndCanP117SaEzrb1ocqI2TAb0bWbiRVFD7GMUfVYj/R3gJMFktG7fcbAZ
5A7qQIqTPFHpELN/pSqVhWaR7UHIktcz/7iWmApOrDy67nlseuIgAcsh1kKamTW5
6qRNlK/ZIG1DB2X0SRBqvLLnf/f97GCPU5Gaow4g90+RtwuHzh4+uObq6FpDxrAE
HRt+AnewOLhhW9BDUutt61Tnt3fFV7L8zE3MJJBBiqVnX5Kh8EPQ4COPjMARt5RH
OkXOo00iBaf+pZ1IZGAL8NqNNFSJ2pf3Xyj3TAvWW7wGJCOP8BLV8xbVOROVAxs3
L7TmFW35LxDlKEIu37jjqH8MJanRqEGmGSGyJqQoujRt/rBigS4QpCSZyIabO9v9
U99f3daL32PI/vmj+g5xzTItabuoZto8cUXxhaxc4eEoOxQkXQXVqBAwI32vOaaV
kKxugGNjMRv9nzm9dyLleWJ44El2UnGGXLkA6glAS9iz/VJ+6DNVlLonvAXBltOX
9ijkgxVBbeAgIVISdZNOdRLNFmAZ75NecgX7WrBF1JDHYWD64QOeMJrMquBp+zh0
m2uZ/D8pmSDpBGRqu4CYVDPMvX0PjlN3SfiMopBPPl+kiN8+rx5GCR3YDNtygx91
W5crnK66c9ihICJx796b5URR4/AqfsczYx1RKtm6KS3ozV4Sn4e5Pv6t7Ab2Uf88
c6a+UiUb0U7JBa/CtVu+2F7Iu+DkgOh7rJqjGC0CPpx0cLY+UHnO6N5RfVgD6Ylz
zEH8YR1k3qcefuXZm/XXvKR+mOaNTGGlGAVFJOo1mPugE5gkJJysD4Zvn4Jyqfix
9gs+P4cNAaHVK3O3YiY11ZbHx913c4Tfcbm8PTBQncg15abSejuvAq3pvc+d1Gyh
xgAz9hxYbcPjxd8ixhI7bp0Vr0M9tH+ii1ThO4VPj/Xm0ceV5mH8Tpnjmd3BGnwQ
31uhKaQcmmtEuA3V8hfSs3xgqhBdYmmP/qBKCJpsstRDyCzynbYa7PcwLVxdq3XV
Fd5ELUbaNlsrZagS9qrX9j5MntPC9qlIX7zAHMqQ0sNnl/zBOhN6+JKhmBDw6LMl
0PvzFxvoTVGlyh5AoAyvsWCneZGkigYRJdwU9F8rbnFan9FGzPhHFH4MFjF7sR0W
TprhJRgRbH92pC6SyOGh4+odIRx2lSE3bQhI7uYG9TSEO4G9dP4qykUR+0MdWaLd
GzqmHWw40hrf8dT2DpJgOp4HYQnLNszbEi0oPsh2FdTRWMVvZbq4smh3e6M6iJmx
US4MKvlxVCltYqqcYTPhGBCsT9HleBHd6G5h17w7r9Sx4Kcy8YDJHj2yWw2VhxvX
AdPLC4I/70L1+GoIQvAaDxKDyA9oMr13OsZwvNLbLRMIPTE+3F4+9JgPjqHpKF4x
1nATN9p+mrxRh1nbcJuOnLNf/jh84VmsJro0VqLd+oCJUTJAUp1DLYK41/mCSFt0
/YmBn6NNbmEdrCqZB8Hbf+s8C5uinUaaUimyDoYvMicd2ogI6ZJc+LKp9dFmXOg3
TG6MmR+tsgu2IX/pnQZbqG9M/y43Ih6o5UgVrqzmFANcDpcwE/1h2BENVSS0Ylti
Wqg7GzDKcPrRtZdMllF/MW6kTiWHQrVYLbTXeJLfa2FkEflg0EyR8pdLq/NgFzYH
lu+tGY4X5cOoWTEMwGk5H501EYrkNqMtxUkCA6Nq2nGz2wylCAnFsykeBMqKxqM5
xaLqfvfhULWc1UoiuLo4zV1eZbwsd6ttN6d7dULjfutYpasyPCOz1xkKiw7Bl53d
9rzU9ak86Tu2oZw0NQ9u6d5bBUGiRJa4mqeOsVD9kOfXbXm3iM5LyWTi9R3GZN7P
JIOUIRAESctUBO4CngzMj4LMfoYji0xdYzEG2K7p66TQsSdQErAmh/vKie2dOA/7
Km3rSyfzDcoJCug+VZ+hhaq06TEqnoF1EHIyNoVuFB3JfdIt7E2KLItDp961BxmI
2g4uJJ2z25m8hBB55nHbOUkyhY7tY/0RyqemdU3cgoKfOUj5XSL5o1czUk8re40/
gSz+HBAxWqC+44olEguttDXgu1R0K69dq8au+taZ5abIvLr7QWGTgdnpIcECfboo
X/faN5ZiKui6PGaoJneJtfKmOKpkDpdqWr2ecy90SCKeldlfKPw81Jzzbq9QguQs
mIcUE/TU/boTRsQBhEWPZH/iD8DTZCEjWSTHXF7xa9McSP6pCsQQVArwA6mRltWb
KUKPVSDHQy2q3EyrbbahMJjCecxQQwK51wN/2iWkOQx05gSa/hsMmYCvuABYKTyb
YbxaB3W/IBg0TQv/dt0kZ4b19NIDIE9XFyYHk/zrNYcesrUDBAkTxr1j8/oWTRj1
TuFuxTW/zbs9/qCzNOMR+vCf57sy5aKgQVBcoG+hJN7ERT2QCKkGGMXOfq2AsxH2
F1KCOIXrPqikfOtV2DoE114/8SIa+NLtGgmzMFrZLHLz2nL9lasQVrsKkXG3sjuZ
y1zDu+RwuuM2RNL6uMxSA1vRufHn4/BcwM1QJnmVajA4PcjL9zd1zfPAo/J3koXx
mWz7GH3L5f7UoWnXzLcb3TjZyKpZdJSzfpX7BtntiloBR0XkPWzvcxnqYr0aXDab
S89guYAxyw/hU4Eei2v4zmshxwYtEpvLFSM2853gwcng8pUyFLc5Y1fzQ0JFqAbl
tpbytxAlwVWbdeMAys8hyDN6dMEnE7NnKr5f5CyqWLYHSc9HeA9f6uqo6IvutwKx
LeSyX5KUei6iXdbYPEWBwWoKBH/OgFp6yguSILRP4+93Uz19aQEV8r9Iyq6x9KuY
2FNdNKfiyuABZnbruRCnL8Qnk5G11YI3cbvh2TfxLi9JVZIu4/hKQdPSzJ6Hl6HL
00MA8ywXQNagP8q45hqFogvbi1oTdZW1GOiNlGRHohQgVJ2Mn2PKWQByccdth0ns
HoH3dY+OuRXyCqOjt9M/O9a5v9QcBTcdP01AyE9QhlxScK3LvnkkQKw1mWDl5daB
zKbT/mPcZUMvDgU+XnHF6tF3wJzaTU+Vd1bJmbc9zTbs7DXPVFvvgKq/1OLy/io/
LiiEESnLJ+oJA7J4iNhYyL3YkvKYetwhzOKK660x8puDMvTVzhcjvGVcN0p6yF1S
IUFz5fbpWsfKy2en1FUCh03e/GnPV+Pz2Pou68C22J+eAwxqsZlicNG5B5oWnidp
c66KM/uuUoNbHb41pbkZZ+s/7yi/xgAiSW+JmhJt1tFLG62rTiwsUzcur7cP0u5V
1msmNT6NqnKKfIX6eWd4gkLuh4hk7rBxbvBimL0M3pFS2yw0aEET8eDU8D8c7o1y
aaji1HQR4CWPUNEXRILHqrGsIzQOJwW3xJeJ8h/GWj7SN3LV/sYMYTamFY6EkXHp
c5dQswFe3bmIpMw81eFk1GllXJCkr3c6hE1T2yJsKErc2BWxuJdWVeaQNI/t8K0u
3hg/HRL/oe/XYRXMekg8kIhjd1xPnmMu6sSnzcghOz3x+nrpEbsmd+NqMj086s4j
ywb9EgSiUq+T+7D3gIOeClI599GJ6hER/LK+hsFpkH+slOOAnyn4vERG737Q0Q/K
VMnk2UwTXGwZEbL11SHed/+Vwo3csJR44ZoSxSrgqv1IkfB41p5Hs6X1b7zaDnFg
uQm4ChTKQ6xL1OlXe/h4skrZjwijmJAJy75nccXLJXLUg1UKknyMXtFM7zvYnNd3
iu7gAIKbMTYusxwq6rK/3umXQRsRykvIQ9E/8pVnHQ/8CGMiwB/xrs5GXRXH9zR3
gwRZ5qsSRplorTwqY3gI4Sbb2SG443xIZ24CJTzszYPYHFKm3gILldMhr4EWaHJR
lHEJ6rFQv9CM+u/3g/bJPScfYD6+deV0zyOFoidt1xxm5aWx/w6+GgOIOH6XNoIR
AJi/gO8K7T7jjHFjxRhmTHjA0RPa8DhvHhG7pZzx+qMwUq5BphzEDAPLBrWmMsNL
hiYFHoxOgDQxt3TItXn2yPJc4SwrYVzHfNiH8j0V5Ek4aYmBX0oc81uGS8sCyer0
epxEydetsQixpf0Vv4nnVK1vjPBr/gMgvlM4oIpA1FvzkdaDHy8z5hNepPuOl78w
tUAVaSx35h+1j8OlbmQX5sx1PyU33Knw2LzPqUQAGjir6fGfCWEFu6yewvVtl99i
Z7Yj2v9GxTOmDZQEO3c5uoDNPk2KzWqg36tLpJuU27W5h31Phi8HkbHkEINkJNKh
+PNcIoTGtLZvUuHYOYrVvSclAcEADdHdy4V+G0pEm7nAwFO55m82iE+VaPwoU23a
ZcakYLZkyMmrrN6PM1QtVRmoFyCscrbba98On5Ce7emQSwLeIudoFTJ0jGu7AsXz
Rm/2mciQxuAE22ToT2oAJ4UzEdHh0pZbJ5Zs2b91r/5pMxci8sEqATxN1t8rZLKZ
mOksqzuVF6V1C2PxUXzZQy/ISoIeNeR+aqKFWu6hG79VVmLDB+Mg8t0/5bIc9p+Y
OQQwXo2WQdTDzg4ELw29nDyRKQvStm0Srw8cPAOM0v0D1JFLzLRRgcEryuWHiuUx
JmXQJi7q1hGL7xy8jgia/b9V9GP/LpbLZG7EFsw0dc5SFrIlzlORvJHmyU54LJpL
2LiklViZj7XXT5wRzw8we0ed5zt8Q/m7LBeTAz5vKET3vUmNgZeuK3QvMsh85n4b
bgNfMKwNQhWzOYWTnH0WweabrEh4U8Hf5jKiFWXzn0jCFBb6FXFtiJrnPfV1TZS4
/qYLqp+K7OE2IsdPirobzKVf8/3rnVcE82TkhViJj4ZspYcCI6+v9pOSvPQNWy8p
dIxFYA1JmzuRgA3UVrzJJTnzERC12bkYbETk0YaBcdii7wRTsvDUwAa6LRgg3Ots
byemvKHUwgOqdCfUkAm1wvGBohwg9pXeHCFNotl7qOolWhNJ/faboYs/fXcmjG3U
4yhhHERWsDe9pEYPnsAMTpCPSuac1XGuSZnyxxBPR8jenL+4vcMRaXiRsWYKTdiY
mQ22NOKWTi7A+4DglsJvfiZHSpPoTYcEpROBVLunQub2DKgVAa7+odM9bm4qsZx3
qed3YgSuyySQRHTmg65t/DKgWyNBp3UUxXbcwq0RbvPLYzoNmkXSRguPYb9tFyDL
KjEPev6O0ZAkqSFKwbbMZ1IjsXtpf0o0f+n+m7TzltmzM1XnVx7Efh8ghnRiQ+Cf
6COAlY3q24xef6s0TCRQtRXyYCkzpxFTnfyuoB1DXnVHvl9CYn+AC7nrx/e9MqYx
ggfXRe70t+5Q+E0VYwDSlJBwbvtV03uLEqq3AempF5WCtRjTVpNSdmh0QgPzISiB
Se3l+R2wrUiHA/YbMSTYYnGNPdQvCjHp9ZoJHgIftRqB1PMjmbn6G72n4akgr+fj
7XC7pcZAOmySs/DFsqHllng7zKHgzIhDgIaNOGxEWKCrRdHmLNsc+vgOnUL+T/JA
okxhjQ/oQKWkw36DlD9VipYiqACe2vwIzTOqijR5dqRjr9NVkGcKMmE29vwMSOf+
a1JGr8HDE2TiS1npSyqq7epEcS4gj9jjtRnY4jx7/3AVlS7aLjOoLfdivnJdnpUi
T1FqY4lJNqRi3IGRmHB5E5qx3+UmSxDah90vwAojx776YhD5oN94g07b8KVJQ/kB
v36Inyh4Jg1Xka8AlfBOmXO79crY1mI2xPxAZgJVwV8oF3oe0PP7wb5MFd1Ot0/5
R2pf5T+c2GA6B9PwkHeUFHsPEwr/3INKF6AH6JgTg+Jectgvuf1VtvRLqLdfFLVH
WvnMSYrPGE0Kt+s45U6YsDGV1tx6ORu/iEdjuuPyNQIzaCjzNs9iITnaUBz8FSUW
KdMknibv5t2dSLj/zqNim1jRqfT3akEAfhoWJwj7Mo5poQKgptC9e9Oqk7X0h07T
A2tGooU/m9ZKtif11ABJm3eKLH79JPbf4oCElO5wz4gGkCj4ln7pn/jjP1yIbyEW
cOaJuNbVuVrefh07e7xzfW9PPYjn4PIOdZek5uPmgh/JpWVBHiuJ0qCFxska0/5z
wOIUf/GnUj5rzwhIi7Xt3EgkXZ+ODhy/t+zRBWc/6HyABr5RpyqgB9UztJF+4raT
5v5IoZqf3S1ot3URFd32tkOmX7zWKvoc7CBjoZGZLHsVViWO2upWKrBZsG2eOfDk
APjJ8bT5LkYE612MswOEpqjW1ywHw28pLNQXB4eUZsUj6X8gMVbF5bSK9CHRmkdw
krvhffwv6For0qcgqvWD8AHUOFwa6hIo0Wll0pvEGAycXKBmWA4bqo4EjP+gTDbh
Q4f55+ph+wwsIwAEPpvdJFE1VgMtWr3xHpDf7yIe1uGSR5F1gbf9MWBVfMmDpx+D
wHKwjbQncKFWQztN7SIWXiYzaeKHbVmFXmYdPb5VY5V4Yo1Q+T2YWb0vVJeBDlpk
AHeFicgcRcjGLCW9fC8UbUaJRPpQ/1MGkodCD5ATYXMEdRjR6vIkyE6bieZjI4tN
5usRLbzEQZlYrWSAZaj8YAiTlhFkgTj+vyKKf6hIN3CI9OauzqajFkMNAvtRT1ja
JSAEmNAfX7C6GeMoBFX5q//HmlxPX99nFjWwporTEfTSWjRQc+7tvLyhygBl7qFq
lLLgWHP/gx6Vl+//Pa2wqRT0t8RNqIPZVJbVD22xGt2WZMBrQLxBr4MY/b9vFtnY
kAuDtTwWOc5zGxMzGOJQVquy30KB4f6MLmYPP5lyNFwAuxJsZFlafhlCjYrZCpuS
VZN35AB96j0jpjBvYA5HjrOc+Zyd2YAVzhFv7I7XXLXdMkz30OmO7UcheOfgTWH+
yVvzxGynogcWh20VS6U2INyT6YYJiLoFHw6bDhZSckyjNCten3wD3QmIi9T4A05p
8FwwtNuKupC4fZUwZLTiNMWrdCja2gUjJOnESIGzRz7iKPABvvHFCUPl9V6mhoxX
UCowXmnFYJ3rnp84GUXSonetyiLVv9nR4CED58VU6AcQxDnsSzxhIAJCpoN0vWIu
YsZDq4DEfGW1yfQowQem187NYEcGU+fg0EskPZ3SWs07nlriRajcqzNxAZvoHv0q
2QofzVIeb76Zwr2LcIirq/RmFb1TVe27Qr9K4LLaqaMgHtVvGal3SkqgIso7p3Z1
lbH3TEPFSIiDu+z6NudRBH8Fzw6Rgcr4G2RpnUuL3Eek1/O6NCcW2RttKQPHnTOk
0QzZcXUidBfhz80fKVcqgSMtx2fB7GDCnY18Umwjx29ag4nu3JUwNHg3MbUcstT/
z0EY+ixEpBy3TQZYAdeSKLQFz9woO+Fb93uhIv3D0z86aQJgTmlOA0QvoHcY15iZ
uG3KZ/m9w8TcTdgNcBUacy6tCoEEgRUTOsLLLNAKv/X6VR74CfeHtd+ix+0o2KJE
kSNqt63T+zLKvo/LPSz53ZPnFm0jzmf7qaflVF6CQHu75VwXvswXLXg8zKVFiw4m
l5bjrejY0yK7De29x2CVIEi34RUdhaZXQqVXt7aHl1PU8Yj2g7MOJJ3YHXJXrhyF
quT0nhIAS8x+On/Vm+vx6fAva+wevLgmvitc/3J9gK2sOpVdUHSqa7GSp9rwBJM0
oVqZ1kdYUK+shr/f3aOv1gQnSpmoQS/tlQ0sQEp7VVFyHS29JxOjhGDDdxGOItkI
WowHWCW0f4MJLCMZ3c+ILbJhlIzCF1/sGhbAvtUSWcQXkd1AOjc4lGeYVfElnSEZ
xvpO4tLQUa+5hshqfVo04W858ZJ9NIXmQmjtYzbgOkmm8sJi4CVkMqbQA4JYNn1E
fkMKLRORS5rE5htYs3+iNiVhWWnVMpqp3RQi0gHjaf540saX+XQbdRl2qceO80yn
awxM6SSqwXB0dv0LCuxYK6F1gzuCg+ce7zb/xNubHfVWnR9Ax4pPKqydDmsFVJmy
KwxJkZh7tAxrT381adLoWLj8oFXjgIuON/wGm1IpCM0iqeoVkFs8QC5d04l/nCq0
Fmsmxw+EPbJvoVKde3Xjl5bbgXL0RMmYOJIYh9O9v5G9dz2TfndqP3Oxr+weA9sb
XhCN0JqjNXwHgvbPzPSIMyMQuBDUCNcrYKKELdDfxvnoYgdLq0l19Qo0IrP2SfQf
ppXTUSF4oRPyjc1zRkvUqZRoV/TtnDyPijnd6S4StZHr6AsQv6bm2XPcadF31FM2
GJQzq7v7GJ0nLpC48S4O8osrSO6EIz4Du86ndRuXykL5NUf8vi3kxizb9xjRJIvJ
Az5ydCAtMNOrQX1aeUVT1sgOYQT5d1nf9XglwH93tHAGt++MJv5fKxptfps0v4HT
bBjPlA6gUTrweWNIuh2gU7w7Pm2e8iyS7gxFFPdFlRicWHzJv//rzNFv6OZzd1bd
GIc64ygqSMlFeNoRanBmpt+5IEjtTHZ8cK+2lpz7b7a/2uDoV2rv8r8z7mFFwv0w
cEf7kU4YJYncLqIaiEQ1dd+cic4SQRM99+ToGEy/HEBqfR+x9skOLJ68NHkYEde0
iQRsmXhsBqphQGsV/ntnoa9skgC4irYYt1THH9aSWry5gEvhUKFtIde+NeQRDOTr
eK1CUCS0wDI/QlQxyO7q0yFzTNQ1TCx5mTu0F8kLsab+JReZqqh4d77UYb1mIdYe
iHvXUShjfoYIuI9b8YoG8GjchdsLEPyE0DHC8zNcHUz8GtoBsZLPNIXriZTJ+Cja
uCxAElsCNuj/dCIC2q6f5njDXia54bM+BVOINuPFQVsig6JWUD/vOVDD6uo0O1LI
mrtuAqdr25fXaezMVgYpdK3/GaH3mh/NbnT6WStuFEf+l5T9X0CeU78fx8H5MrSz
mNCp2OO3pkJ0i5eBC8Cw12jFiB7U1qGFz1Fy8bVJF0hGRBtrVFBuV9gMJuQn7ok5
pZ0Nwq5KTr9zUgnisxKnSZRtumOjusX8oaesfNS9/08y2jXCOL2WwCRf4xhSe1SA
BACKexO1vYFupoJHDuBoLrvD73J7kmUAl7LQRDRYPGlVBX/nRhJ9+7/ALssvkcM1
7NxgkgaJ81W5zMssezNi27BS8fnl1QdzGvyCmzVE8g2uq1vy1//kGJQYSPlHjdeb
zk/IeTDLScPBpDqCKhZ/EbNKalVBx+OB0Uw29BQ3LvhgE5cPM02BtvpMKStF2iDT
C7UUX5e8t4NRJ4vUtxRHj1zFzKz5KFTYKJVB+Jh8fo9VzvFocbRF42kJHj+jCGhn
RK4Gr9b1fWLNsRm6FhDbRRafwztWAur+rmp1pwivt91iwydTwxjqWrgD35Jke0Ut
E3K0jraSn4VYrjZcFw4jwtdLYA7u+iqfExrNcpGagDtWTHI7qJA15WELGk02dBkM
vgYUcdgjv9KwRPBaScCiMtPhZQqTFROKIe5IvLbSXIK7xm0Yj3jBd8ddwflBx6Nq
xfOTheLW3px3ZQB5DszAAs+slfXgaA8EqpbYW/GgrumUZsWZHgeutmR8Ez21lQ35
0CwsSdCfbvZyv5+R+6iEqAwZIxlq7FHqk333kdcxUsDKDxgaxwOkY91HCX2anh1a
SQA1GS76Xahv+6Xa+v+sObHWkdGYh8jyGX3A+kBYIXHv+vpyxWhmtrZjxIdZ8p/h
uCcka3Ud17D7Zx7AP0bhsPD+/LvUsXUs7z95JzNHW5Zl8xEYvi7wQxHJ1df47bGB
Nl57vH03TSBtA2da3PqSymzCyO2xL1wA4sgDEsaO2hP2CQpclKBymKjhdxWYkdpD
3qAWZyXMgh/m1eUICCzauNuzV5EHkPDQBILbiyzcvkvjmMAY0g41UTdw+MFi+SFA
MxRHUaXor2OYvWAD++IGxzg8IOZxq2dMwj/n6U6jObZmpOuJjJQHhoqK5S22oFUT
iXF2hKXWc/Oih48rZGcm38p5MvIP7TYBKqAHULuDPLA2CdW2kbL2ErfLvAA6l2NY
rgdjWaIUA+3y8v3rKK9ctuwZoNeDSX3l9MNTqhGjAKAnWkm4nZmZaWGP0SVl8dUL
E1+jKZUB+0zgDf8Sn07jhycWOPwCdWA212qYHklWD52qGhxxBBpKUMiyk4vJKaWP
eJMqce41UnHKYES8Tl+YKXtp0Ninc25hMZKW2qDEiduYsGow4QDZP+VKN03kedHX
MjSDwei/CtxLbPrUE6fHovWwCzPhn6Xjk8veLqefPYjt3BBgwe9jEPo32f1pnq8l
dbPlPuBGQcE5sd/tojoGLvHr9Ubh6eIZ5zuELNvQ7PdVwZSx+iYiAQW5G07rHybt
7ZpM23iyxEsmUqkY3pa3+b50DFsZGpcBxZ9riQJYUTD+McZnJSBdLUTaAQYP2MeP
QGsybSb8BILC5Tkkbp+jTMOT3nZbqH6EgxIN34pqwMTeGpUitnS5AE6gomjpMQ8D
O+d2l2tbDcO40P22rCmx6kId/LNHxpqE9OpHOHWs+Xko9A8EYdLqkRn6eam622FV
ZUp2c+83IBuz650GhGxxnS91lTzH1r9HqmeTiQb2XUch7rgawmGdqWHqXmm951+L
qKH9zTZMjSXMuss3fTm9o2OEMJ49OJuabDZRyyvRD/sAinZjS1edmRqHMNi29Y0r
lyWFnnCkvYKJ3Qw5Zihm0ic/1EgFzJNXp7SHEfRv9xrg0xS3MPv+0efYehl2+cWv
6WfY4PV9Z7wNZU5m/4j64MYms2qqVsaJ5TVNeoC3x1Rfwy3Mg8+EKi4t+4bdM9cC
FsDD5iHrFwJCejytNu4N53GjC2W0UgtQNdEo4WXjOpZAByOmxcl6UGksSmyDA1Bf
RI0r1ypE4KGclFOwZA9STP/5OhVGb7ZAEtJx+lzhCFaHzCcH9O4HiNAji9iTVSsk
Dy3E81cSy02yZW05EuzITmhNRtS8RCjkpUxm3s6bQUIS3A32VkCSKj+Vd50LQQtu
gAs+2gSlznxtJMnVo+9VzNtOXD6Wmgrg9G4T09s0JBy6qpfk0fw7nr8hHol8960A
gSmsmcN/x2S0gtmwWfwzJyBmNd0BfFR2ozCr7vvKS0TdzI6cpBsg4ScIl5v8+s2l
tXqsn0l40pNVpnpRtOi88LTXH3ywn1hjmBnPQE1tRGsICwZGyh6f6NKYivrsOYy9
6ssysi3luKBL4u8zvcMeEiRTAH9IHzXs9io95QtpPRxz0fuh6gS3hHj2pFT0lslJ
NSVYuwR+SZ4nuLuJ5W4lWlOPCdEYU6V+ITfW3jdjt+Cpq7PYyWSQvKFXUUXyKqO6
aL56fWiq5x4yqtIW4FgQdYqA+hWLCOGXKeraGLOYDcRuzV9zBlZvF5JTp8/ObO9/
1P1+08RdFWImeRhMB7cTsYd24JPYt9mmC5FBmysEi8NJrBi7MaBnt1TNsmjQfWu5
jVqjEmGgobIaaQlIfMVTdAXENeFS/pCQVwzLklN+ZykBfGtQad3OK6D/ugwPmwXj
KQrvWQeyablHqMy0BJXPDVNbFHD9knbEOSbFSj4ebxvMwrMCPchDxnorxxUk4779
P+qeHSXmYBrE1Vzt9pSxavujeh1O2YLt/xfgmZ/zVlijMiWP0q5YWtE2iVFG6aD0
wjComj6jdIQBUP/l2waZlJ25zKZ5eOOerZHg9NuIG25TYoExa/qLrq+O6sKNzbuF
/VNqxsic0NjgFqNhwpB0MziMvOVoKDcKRumkVCR+jdP8vz9hWPDDF/e3JRK1/fFW
dAnxpZm7EwjwS1uh/fZ9yC8lkP2/nL8UtPwvwCpAYW4vv/GvXZy8OBSg+K6lRIIp
MECG+aob8hp0xEWQphvTidfUZ6LrQxOsTa3mz/Wcv7+ad1GMKEbHdoEt0rLi+IEy
ZCtVSUq6z17WV01+0F5EVqWvhJACPs6ZLkz+ReIw6r+d02Q9faGVBGwhCgMUuRAa
e8UN4+r0C6cpX1aPiMN6YraEavOK4MkTtsM9Y+uunVT2VLePUjrybFzNa91ALdBV
gLKWnUP2yTTQEGy02QGFDyiZvFy3uIFKw6fUwZSO6xdfZ1J+yRZxqP39cf0GzlBU
Joyqlg80sYHOKnFXCvbheaS2LNlajCvFznWv4S3/hy3Bld2rab9c9avSCUaeY052
PRHanOOk+RbCIzn96ehSiHCSxxI5WVROQvrpoobzF1bgNkxMA3zqoi9xrkzfXLRU
nbm1lt5erhPy7SSqB6mDuQnq19jCx8rxIpCmrd40zS50up+JDoWY1/aMSZ4cqGMU
a6EUf5TvGBll6KD93PdbGBseK7ZAlXybasSmAx5GG8h3ZjtJ5pAaFspLh9Oyie4q
xn7wqKT6iAptjLx7EjfmY936lfr6x896QDJKXVTvYAux3eGWmdwG9c1sCtot9yBR
Q2+VQXhBqxe9MWHizbJnNn2T0owzj+qKDPZG12sLL5neHoLOfcqqL6FE20WAesGk
Zbs2nwmLKvySFD10PwqxIfVdO61V2qtaW/ApL5Zr62PcFlUVoTiW+yMYzmXRuuyZ
MPe9Nb1Tr+45QCJQsqIzl3ICcr1RToTVynJlnPrLQj5yXczaR5znyrR0xkmrNZUC
SLxSUvgh5jJPCyyAuZ5sVYGtwyrlxcsZsNOsN+kkVAvhGhT21Ib5RJUv3Y//1ouK
wg35bEdrkheJ3CY01uqG9xLRopT8DV40mRvz48OQHsbkFVWbPw17uX0sih1E4oT2
ZLZ4r3lMndyEN653TgMG6WB3R6Exa9yF/TcGx6LzKJJOnZrO+zWvp+OMV1oQHz9j
U+/XlzSFNpAUyHswMZHuXAG3QMf9DWlvNhlw3TNWlB3ITgzaPpKkiTBQOMvcILTo
oE35OfADFO5RXVbbeunAGLEunk9PS+ud4y9pUjijNhFg1TRi3d42Q3t7J3GLjMyk
ZVNFYNYVETkRnNmdR4MAMMbwPxeGZzhRuJ7nqbgmIBV5OJmli4SVu811O0YNZ4ZO
5JMfMw/iK3r/gCceD8LHXEzjXlUdzOujAWzkx8smDLjWCcm2e/ToP6i/Yky0h6xq
nwpbkoVgGKX3s76ZenBEjNtXD2uu9DUn2DK9gnovUY/Oe03lQXFI8ogibmtlYG2U
BhSzdyf3Q7gOQYBp+0n0XhwezpRSD/N3aJvH5rhc8jpF73h6EsBExjg83M5jmCdl
cGRAUKgFV4g3VYUY/lHuMIfFearNP17mVxDfqAKDVBC812c9IRjdmhO4+8SUztD5
nvY12abOJgqh22tP9tr5LMBl2ReutHhCM8lNvVLXA0nP6YYW8p5YsZb5QpI9Kq7z
k70CS5xCscfypXuZr6FUoGBpRRuPXNVjGp9Uj3RCvZdsF4gdS4uXdZF3bQ3OWtXZ
R93Q+UwZx+FD4CtiIPGEJlsSVnQPeCVtLm2UFrbzfELWtN6bL5vZIH2hiiNhIR+x
gZPJbtWmigEjfqUh9lJedJqssXLIPsjzUr/p5BTQBb2xsX/ipPkR1+T3osXos97r
FVB4QXB6mjzXXTd0gchi927F6dV4SPFUdrjbUbfnRz0PhMLTR1wHdim7XYouSNH2
hmLqUXxdyAxuC3UzwlhSZOG+dUdGU9sy3fka5WFOA5JTDYc3f1M8ky2hAiHZfvtJ
g6vVccvW+DyNi49PB0MU+K9EVIkD3Z7pwbZ+1X+whhRtfTt4giwGnD7TQJUD9EIQ
52DjkaiHfB5Xlx2QMYOaA7TpbEcL1g/RYJ/WYvcyknhQCM7lc+AyhyrFmg25EyXX
wxPqFmpSJizGvIrp4sg+G8MZMRdzD48gWuiDvCSzNVPERg5qQMxPojNzpSJiZdXD
ahwan6JkUFt1esLG85vaRjoq1G46wqHM9CLe2q/6RHTwdJazPFcid6QcsTzt/af8
/CWWcJeB/1bnAm9LMw1DLIfVlrHTUucMQHZiAiS6xlQKV87GMYVPOsGcxChDEjW1
/3ThrL3Z8J15RUhjvtCr7OSmKcshyNQlLp2/l7cd3TeV9T/+Jrfd2k8oCItyXyj+
nP77Ir2rLUY5QD14YUziqPS6h9RjjUDuehc90QJ6HjHyRZIKkW31PU0A0dZs8T+K
QXOvcXrPSJWFGxR4qhMufV5a7sLJFlvqEYYBaBkTF7H+PEx28AogURVa7QL5UpJ6
ElK43XMH04a8A/gFCzWbwzx4J7L3Z0gaX8uwpCCbV+Ts5pOO9j1qxX2FnPbOeoy5
xqYIyOMXzpyJ7BqHiHGzLuar6UDy0xwOMGAiYgZp7ss6fKEyYY7ZYJHhubWXuhQ6
E7z3hPTRdtv2ZiKfSnFIQLhylJfWTbk9sRfNb018+rFeVy83pL+jY40nXzbwEaTA
S4lqcXKF70/Lv5FQ/DMMgTZqPUrt0fHt1YTF8fvBIKHZ7rAPLV+lM6MHg76btO9H
hYbtu4EM678cPUylPRLnMQTzFedi8AMAQc3HdufNF684x1JMLK7Pfi9jippvfGB6
eGfXiTWBA95ha9IdfTWOiT+aRDWyUVsHMwgJJ/dVbni/I+Jmg7ZoUAzYaXA0Klix
3hN50yV5pYfaLoyGyJz3PsZxFABkBydIM37W8YnS9ZzclEPVoQvy9UwNUtm2j8QZ
gifuDQpazHvsc5lpjpaG0Uq6V4MzsJb6dwS0gb8E5mUZ7YYKQEeKei6+Ap5PH9T8
aVc6twblMZU2QwcZou98b7HuKmOZuNzHf1btErPIrvsSPmtnwW4NDXEDK5ZrrnaO
jpSWArPs8fVw4ZMUoKeA5zvtSPMa5Xiec/bplOqtOOnNsy/DhFpcDaMB1gzPd90R
vMEuVDITuSFWcxgrp2OggmAijsnKK2OJ0vr5vtrgyy8wKgdmOiLrj3KF8lwrLA1z
eXgFnJjf0nnwnPJ0Iix/Vx/kyE3lL6SZUYoNISCA9OSD2OOwu3R9wxSBFqtC/IS0
C8YgMq4Kxmh2kG7jIoJKSRtTLM//Vt3UZoS8chfikf1Az5dfe4Q7H2aYnmlj58vS
4dzUE7M0GvE0UXRjT+a3aLGEwHoZJXr8/LmVJrvN5q++Zj6yC6t6lgm0QKitUSbZ
s7ix1PuKzMRYD1o3DZRjLdl3pkyXMilocsEl7gamIZY5v/wEyP7VkPFUPNnBfYWJ
jZVrxWuLlYnlGinQOaId6UfQvKH0P8vtUXpmWbDQ5uwEm6DZBrEP3OPyn5gjM2d8
ZD3xorqpO1GjzRGb7wH/w17uez42jBMe7D1tE/XoL0h7c39BmJQWm22B2QJxFG0f
8iTdPbYuaWfl7S9JHofWtg1FSE9uQxhhguG9M3j8/Okm+le43M50Kdm2u5QpH4wl
DrhbHb2UPWkzc169oqneGviPul3buFncnFHNwEw6yS0uzqKqgPFP5Gqp43Z9EQfX
KDOLMooQ+3rTwZUqDUMrWj6D6b0KdkVjFkKrtzQfvdwMa9hmqa+iNDl1tKsCwOi3
P47z9nSX6jq99+qmmINFyFsF9jY9ZnogU9hu1B4znxMDR3gP87/J4XrugeS0wm8p
aVP5EJvlnKotzPEHMDwherT+VoOnWChEeQKtaU0IRU425lBFM8+9dCtkNEXbJk5n
7F2QLG0w/+hBIDJRtZVsbRXXJAlHkrlEmcqv2oq1gQTknv+43fcWVwkSqLFSpUar
ojJRIdhr1ZDaH6Q91bfkl46/erjivGHHSUx8gHRZRCM7gejZRdXNojqYNj/WyHJS
f4yF1q/vldID3Cs1NOBpIZ4SqjXXOBpRVL9GnhTkU/VU5YIgPzZBRMGzEyzyfhBz
TQsjSzLi0KNNDWSMTOLIq4FQ0nF3bQHt4x9uVN1PCjEhqOVM+7H+zcFBn4vyG8vV
B2B1/bP31n65v2w5b/CNROZ/HOFah6GxH9nVtZNarYNGTfMbHEj/rLKqUgVnBRDl
V4BBqkVeBMriJ1CuZaGZz2fOBvBExUiewNsoV6BVTNMuiy4+HA1MG9hq5nt46HSb
aakmy580anHu5VEDxxYr1Q43T2bZfoH9snWMtAdz2UE9F0Puv2rguDrBaNM4c5NS
tw6FnYlwdn0U6k/KktKR8IvKdehgozdZEPCFwlftj2jxy/76SUHPKJmpcj/UmMql
iyxsnNP/cGppaUcGaDCoZt1XEwCvyj+l0hwx+Al661CD///4DrCxMlZuNVufaGpM
MhjqMgSGvEvwkcUikHtkKJQ1vrsLZ6BgOVP7aTx9LGT1/VUUgpujdJxgKNM3F1bX
dRoMR57h97IzB7bLUh7IAOiiHZD57xfBBBjQLmDIl2aYQqTec+LNHGgWs77zGDPV
BKeTBTqWdnLZ/pu2Aj0+l2geR69EUz7z4qb4gaBN2bApD4M+vgb3v6Xfo/mL4zBN
sWFNsPQ5MZt3ORTaLC/x41eTOxxRHmGG0ROnOuEPcoVlQM9OgcWMGzX4XVukZxFh
X7bpo4zHVk4Yqp/dSRT0nqOG1FrXrCARz6fbzZpLc3FKpmeVNQ/Y0U8tOTcKNZBS
Ox7VGTqHrsSiJ05zNCGL7N5TA1AnIsQQZS90kvmGtRXiCcFRMeEJToJIGhkM8M0N
Oqiyw85WXr3yVhBq6aFGcQkIF7pIbyG+25K3RamleYdiCIH/yPDZZCNuxrBqJbNW
Mjlq19DlLu/XOtyg6x3/mhqMqVhut6MJVmPca6HidJJ77d2Ywkb2GkeLIU/j7bBp
o5SDdgd02ORCR/XI7Cf2MU1/Zt3g/WOLJvO21sQxmj3Ii7tE59GgefgYnUYM8cTE
wakigaOF0i4TcM0A+ZOfkvG2HXZp2vxlLKbF13gIHK8XW3LDwaimT+jguYdMyNUi
uqbcuUc30Le4eWRjphxagXCulzq03CUNYo8Gai1qaxLUD6/kYh2N/5I4/JSCiKU1
BDSffMxq2FWs5h1PhrduymGxdnijSwiJQ3jHMIwkEgLPGhWE0aS5oUlE5CYeiqwU
0lWVwlI0jrPhf2D/ULzqa9Z27/mMEDhxfaBijfeW/uPmPHvEqhT2x2/qZNURsKc+
ssYf2u+Pa58LGrmt/UqgwZf1U0Hmgnx6yVk7AIyNrRU3wRMTdYZWMR1Ychs1wU8/
ZMuvLamwLlzFS5FLDOn7eUAljjjFLDlFdR9NRGGg9NqZbdWD8CsJhUPkYGVERSu/
OBS7/jNbTnSekKhy/u/O0OYRJGEZeO99XJg8J7rIDUNmUh9WqVSl69Z81px7IUy9
n6AvIL5o34UD9W2Vsx6basEF3lbh7ItCy+8LQGDsFeFR7HN4asIfCfA6p+EZw6Bb
WHL+4oF5EE1MAfkkvxWpcYfI72fsnq8f82FNIy+TWaXFRVPkwLzT84/P2RQxSjTK
QukRgp3pH2O38wrIsxAlRtEAmboPaMt5YvCaQ0KdNXbU9lfh/aX3nCnSb/JS55bN
n4N2w9Co6GvaOoNLBfN7vs/Xi5MtBc7OXKvJk2YGeQUYRp1qzYRUwdvirqMJt4W4
7OSzkqj5JkOaZi30+qT8FJlGa6Z2SiSeZhWbwuYe9K3fOa8fn8CIJ5m2QszBQ0dc
kDP4kHLfekKUZ1fVVjbeJ2evoFmvRDivviSKxjorY41KC5HrOW2jacH4KLAdsj8E
BiLHr26umtLKufhRsmFFyVbB3pOezzSUZWwJAJSCq+XmMrL6atg3KPotK09nIzok
lj6DifmwbCJ6FVf+RiRd2lCo7Z6FKzDGoDvlw+53vwPEJ6EOJCng8jS7HmC3LA5c
pHWKjfdT2BFEbEjcIVse/CL0LHIZ1TlS0QoUeFbWBJGo6I5KY7WKYhReM8RtOm24
Nt5HpWH6+XpIfWONsQux8WRrNf6GpzYKwiiY/Jwk8ZhdG0dQhGtX48tZk7bb+DUz
EAjrn2G2rftavZWSXNdY0wsDIdjtVc+CjlYRPTVuC0mIFfYq3lazIA+os8OgZUWt
z4mmRVH0bYQ+DzDmyVkuHj4P6FEHaxYHTqiv77ceK3l93rXR9qhLRXvwG1kyk8Et
kz2Y+QQYatKXhFWcMRbfE8FGaxCQkZRNg2CvKt4JC/c0q17L+XmfKHXP3YXH9hoA
gFqQoNUKi5KnL5Jb8uJ5jDqSa0pPIPoCYxnULKqxhU/448pyYtSltyWb9ZS9WLg4
xObeEOfhvb57KpeFtl5KL0DTfaWPZroRI6FuxoJfJjVMiSinVUcPAEOZP4AQbAao
NbOzIOea1ScBiZFtqPdGN1tTVfxb5QPqB7/mxwDw6ng7KqZjQXbkR+xZj6J7iLXM
htVbiIWchP7tDdpT1AM8DXNv7KYmZtGhPiNrZJ71145SoaKO/RT5UQoXKx59e8Uo
TaetjtzXtDSvkLocZepgLvQvne/J3HlDTh8nbAZn3CnqFXcLUZinvZ+Geo3/BbWY
2Z7e8WqJ/w0kGm2lFFPyLxpXzv61treV3M4HdINgsK0nJEi5uHArp9TWxFdksZZO
dsTkuHbzBvpQ3DNfk2aHxquLLekzenISYEcZnoa97vEdJXa995q2O1QaRSRqq44c
sR0lpMJYkWQJsuerZN5KwrHe/PnNqtw1TctDSHksUg+m0ju8G3T3cbtSo5sutE7f
3Y2y91tz03XASftQl0F/JSz0UJ+oQULrCSpQM5pfSstWTHmPJiMPUhcBJr/Sz45K
ekwiYXuyepPayfrtwDPuPbppMmK8p8rlH4vyfvfg7+AkZ2abW0xDNaakGhiZGKeS
JqdwuJCNazh3fau7UY3spwLLoNYz3mxCfKEGNKUaYZ7UisH0GoggW/3wJu6NuTD8
npWpo3KlSzFS/VqezT6jEPs3/svDNRqdPX8Gm1BSlb+RDQllTu87fW8IC4sQYJpH
FNAOfisPKtzSj9lSdkJpLEcLwScsMvZ0fxIuNoSTLDd3fukU6A3EABedKBEL3w8Q
yv7L5OVT3OUlzJ0X3sCvsCqiUPn+X7Ahjsow9ZoG70eML1MA6Nh1EkJHjO+MesDS
UEcF72cMR+bpso7a7MESVLDBSwknYI1v70DLmSDo+k5EU1l+vf50QiHI42Muz9aN
ZDY3tMaUfhlXtDWtpGNHKvlN3nMKtlG7Al0h6ndFXYLQROksxrrZq8eA/i+IIyNB
9c2yHXoEDG2Q/yO/5+bnalYjax102Z9KRPyusYbw4LV5+JjtTUabWOfjvfsM1CG3
PWxfoS/4bN0SPhIZ1jbCtobEarjFfPkBxC2D8tJvbrTLX2HsDOKBS9Kb2/xMbnd+
UfoTw9ZfrlQgEkUh4sLs4xtZFk9B3HcFbtbVF3Y+BcBr8bhZuxhJRrZkqy1Hk0fr
ku5e2sE5kgi6vbeWl1ZOOAL8B7oaIBPMsQZQSEnCABcdhy7E7IuqvsJpOk4fZ5KM
KeMozNUqUIv0WOa3beQWVdOpDaflVOrdlYJxfOWPYxK589ifo4PDIhRZFGMr8PFL
DIOhRjF4aHK+L9y+w6+uflRgf4+p8K9YsTVUnnMtrXD5kFIdJs+CeqWZXYqR3diV
pBaiX8FrolStmhgocaSLnt41RYUcNhUcuU1fuhm5XlXLr/uenbEADd7qE1avv1Ka
Mk+FkOAWDGwgr/zl7vfWmFS+e1V8dcZyDwVNf6/TCW0Ns9N5dxpKlMtKyhiRYAS3
RoGFlipm4z3GoELweNZq7/KHn4lwAAun0LUU9a/WJv0yehp87Bj9mylXcUXf/aIb
ojjoyaTi1ZTXVocF1M7dWwVdEfjiLUsq5BB0bmOFPzWvmQDYlrF1a49nIBekkzii
R5Zr0MO8PQBFRyh8uvK4HdLBMwDUPOCu+7UbETXDydj0T77kf4M6fV8LwG6HnMKa
NVwgavIt+jf9cwjSoCY3TrM+YVi/T2qjlCm2zmOr/1zTknF4quc/2kNhH2j4RqY2
Cm1dC4TREd5QpXVXn2ArYiCxVaLzQDwHqDR1wWh15VD4/gVwD/LTyJxSTA/fONsN
axA4HrlGF9VC6DjhM8U7RGxrYRAf1GBZiZD3TRAOjtHuTLNEGnp7azg56iYhzO34
iWg1LmFRWhy0ZYKr1QFSQm2i2k6YL2hbkawNAVWRAMpb5sI5GLmKljyf77Pinng6
DkrCntxip1cfhEpoGjhkcT4fzOYBCcO6KK72Dvr1rLQb4gx5Rqe7AGLiN+ivvMq2
Q3Imcll3FKDk9f1/p0zOVY+7FbArQzmK53mrk8nc6hbptTYpJj5Tj8nQl0JofdKo
LUqUM+0//sn+E9bTx185kze2uQ2opTtP5Tfd7IgkIX0cBJd1J80neJDwoHKbFiMf
mSSMq+43QHI/9ugn2zKRwl3f/4DTKFF2pZf7G6zQ90hcREHHCEYfoldatEEctRVi
MjlqjhsH9wLckKz9VlUuUfUe9ZfOdkfaBWK3ZaMCaAP82wx4FRNdY9f7msmPNQ/Z
iZoiEVN/YH+ItoiYuv5GpdspVpKAnyYD4PEyaTwQGKMlTH7ehhzK2G1CAOKS01cq
j/iAXXH+tLMFXOlqDIYccqvSYWnWcsw9iSZKSRPLY3+jIShUn/XLyn0hb+UqYRET
KQmGMHHXE+0UKy+6WwYXbu8cL7h2bHhDIyyiP5PE+rR9vULcAWUuGN61HkVhbCbI
7qe8zu5nvCCj/W8JB2AA+vi3a5QgpiVjWNQwBwHz9xsV8dErstL1Od2u0IKHMAGe
lGEDQuMSJA2QkgrzaP41AZ9/d9Z6bFJgVhyaR3itopCNuledr047MIZ4fcxVTZe0
FtcWhlod99Wq27udDy/qpxVpbCjCAhDTKgt68KeZLUeDNCKOBJyO/JhbZ8gNpUdS
+UHRHYSJl2PY/BWWFEoO8X/fRGEMrEYzZRmhtQbU15JRS+37ZltXveBglJ2wzr96
j7OJyG4go4TA/B/aUHM0f3scqfa8jDsbl3gyNcSmjhgNELY0dAbRWQqSPBk3Ddu/
j0ZUJW+50iC4/P24Af264T0AGrQD6k2UZTwtzethG0dr5HfIygdkGwqTRSTJTui4
Tfd2sDhUWpLLRdLa+H9ejOL1sCa9eXoI1DnYg5AZN7U/ZyYuvAfMfl4p/5xyOehl
xp4pmJbICB+0BoD2lmzxIBPQyERnlDPWhnUcElDw7MvaAM2TvUPQ38PBKP1JX/Fr
wqAchxdG1CBl+XrBqDnE2K2QWLjwnVrSk4QwhXkkfolURg9M3tpUXsU7WVd2aU+m
xXl3ow9Wdne5AF9kqcM7rMBQQYyoGDSSw9RG+Kt6+BgnRyDd5caI4Stm16rU7V15
M5Dt3K8BujLj/k+ewzu2k6rb3DS0keT8qGmhV6xm3WbQ7L4R/Oc2qkEqt4dmyMeu
QBZ9C3hjMwoQcQLebER1NyC4ExTrYhJpB0pXsc4uNyH7NwpQu7K03QysBKf9NjTB
CRGrMatTjMs6EKOxXP7ZevSvRCXiayL88tfG2DNCL/xBLKI99wjmJQ4tCSi7vlCJ
knqKmOj8M++zqitbOJguGCcNu0hkFxqnomoIrpIcvC77UN0JhYziGaFmdmasrAN9
ZP0+7UIWl1Zf4XR4e8oGZngMkzbx5M3xrtuERTdhVL0JcDtgB5I6oqOpUhpzfKsZ
Pw1yXYKZ7meg9AZAoT5RQvOdRzyGLQY0oddVpNk+oO9Zm7Uon8hbNu4pBQp9O3id
RBHdxU80tnQ4Y+QgZ0eJ+mQWg866nh2hQoCUzMiCXIjj8HfLMl06lZaf9rmvESz1
Lu+GE9Hy8UVszsEgwnZVBjQbN+eWnX8lZXvMweOc6UW/LHEvK4dUCTOYDmV8cst7
qObok+p7CYUOGb3AgdihYcSH+xHzY3fs2kbwuFIxFKLL1NJ07QVivR232h9C+Eor
3Hx7Y+sas/uOGrYZzbFnXpzr0Bpj0K1tCxQhsEd1kSo+fLULJMDoPK4QMqV4CMYM
Obi/ZKugGL3Tqn9xPx87Se5GR+boAF0IaxYV00cbiFwYq+fZc6GFg0JQmIOtLQ9l
is17kDA2soM+mdt0DohfJWR696PzsJ64KZeF56xRqWzEVRrZukqPpItINg+2oAvz
ZmMGaEacWvQe11RFgpITJpAp7U7SBS1smw828jN5n0N8XJyJ9OJI3CYUe7ZVr9UO
VgO1a8NgM3W0hyXzSXJY+lN4Nxn+ST9coeOacVyMZgFUrK2P5KA3ITs9K08d90kJ
YTau88wPjmayzKEbQ+SFspkDZLc7x1mfkmj/uV0yR9S4WFYiwBW8/c5wonh+wBg7
GkV8GfY+7CdaujinPZNM9cthb5cWFduwD+wbWkg24CAd1t13h5c4grxpP8rSFJSF
Gqx2WXMIKqbog3OfW5O4JulCYaX2r43xzt06Kyy9+tX7XLRzsjwo4a68RpDNxTyb
krMCQqXPQw2komfV1wJEIN1kP2RqL7PQAEg7VmHRxK4+k1g5kissuu+PRIVqFJ+H
PFPUpSSuqNM8IWRtSG0F/WvI38sXHiR69PqN0y2YdTB1IfmArPz7BdjwIqyPf2S/
axK/HxPE6XH+28lMrfjWqpBS0p8zIUad19XunSbfo9utA4zcnjbRXIoFQ1R+Awyt
fG0VaemH72OcE5cEE2lxduUXB+Aenh8fJYd0sei8WPLN+sn4fOQeYyzvBURXXtzR
pednJJ0Qn98zejcw4doM+xay4EnFbU370ajzi4Vit9CR8E7BLalpV8vCTqdny6YQ
YPd2MiYSJa77SZyINgu36B0J9e5mdzHfif9hRzuZuggEAE1tg+U+Xi7ak6JO8dtJ
T3T+rbCWGu/4GYHGozzK7R3YW/8gwtj+8Y4a5uiDBaw4vk2JvQWELAnwCpic/3Sk
EJmlhvIV7vQCXFwuJvMJa2H+NnywYkHz1Gw5K7j8Th0BSFteAqhSVfSEnrSFj4ml
cHe7VI7HMx2F5KhbayEWPFzl/1Xli77J6j1KF3q1wLXbN4+xj7QkSuRALs0LRP91
y2kwEqcba5uKWaW6OTx9OEMPd75IuDoGed5hcXlSnJ7feAGXyXAp9XsLnnPHupSo
M03nHROeID4R6E8ip32DFKz1yHrxUGI9JmQ+s/r5hLukDNPn38OJAaUuK5RXtopd
p2ZzJrrNbIsreG2/AwzMZI+325rUUx4s2x+3L/Mkg3stSi00CVOeZpRGW58T+WvS
iotiFxgm14vlTdxXP81ZxYQkGY/qyCrtnf4B/72R+ZldnCEKRTdJWLfABJSNnUPn
rO5iKWAJuaNcbRw0WYXB1QqCWp22QQ23yntYmmYwI/fMWSjW6ZD27i8JS+4Ba5xb
j6UyW/KRdhtkvK+vZLP4FwTNbk3sxSUvZaMa4FdoB/hXuzAE6MWSpKX3HjNk5vzB
LcxmicvtvAmqKJfu/BgDdbv2TSJ2LXT6FWUPbydmdt0Q2EAlGu5T5OtDAhpk28v3
fcqIFCwtndOU1nY5hef3BAYD+C76JtoShhog6dKgeZSTQCNFIqIkq2jORKSOm25M
uv+xcGISn8XtoomkDl5vr0ravHAMPEHaXEmQFGZkNipF2JUirdQr5N4j6QViB0fl
hKVb7JSPbZOycqea0vPKsOlOyOHg5kKF+1iNk5DqRczcv9zB53KIYFzka0jkpdiS
2anoMwXm1bIEumNfAt1W88IQX/msMV1eXjv/dKGnxTpVfigYF++AOuLAvSwnJKz2
bWR7GQZHfHtZ2e4URBysjecxRmuO/OKFKL1qIJU2SFkonDxLwOUhq618EzevGqCH
RB2PcKQYqpfffuflqGJo9vSnjTixCWZ6o9xuVecBOqdoVNN1OJVq+tKvLFATI6dm
nNwN129a1Bt57rcgouQ+K2QaX2ISv6o4Hhk3/oZp8aa/hCsJ3xU9J/d7QiN4MXHl
A9hGLC+cXs98ZFhUGsGs/8zzky7ey94YgnV/GZaqgTjWfgfEj5osiqw0NEaknXDN
lYJA/ZiQJrnvSd+ZdTOhGbktBVPCmhcvmqoeWD/pwM1DU34fMJo7vY8XHq+Q7Mxb
Pp/GiG800JQxPW/bh/2vnxW2jY3WfcuLJ+jlqUlSNb8lgYxcD7hWDteUvnGkQRWk
rWvX9b67FHSTmoBhSBMD+0v2/86oNGkni9aQYd2A8MmPMIhPl97mHYY092PZTBoZ
Jj7FS8gkaOnjVcF88ZLM8scKSgfr6hnUyM2EPixScTC05wkj0Pj0hwlXtNKurOJd
tTEK3xt/T7Iiiv/EFRk9IcM6L4AWsbOkYB66d3KuJ3CLLbuyLky+6EXCdkPGnMoM
m3rGbVm4rGGP8xbQGZ8gPBxZvqzdFDR5oxAmZYWLtuWRiLQKG57S6aji5HrVv6gT
sUSxbu6w/vaSq2GvT4AOXgz2tGsjQzzJcrjq78xqIybc7iWVYNbTdwhn3z3OWgzi
vDAdbD4BYbqQHZ1wZ/2SLgV1yH1ViPcyRlPHiqIFRmbBlRDcEW4KmbZqLTzfjvP2
ZvjE5LA5aydyCQ9vjO7i3uE7WLqYcsBW2Hd759yTGWZONoRFopIJE+yZojEwZ3aZ
2/CITJyGwsWde1I4zeJyKWu+Flsh6NveJF2nA8KSkg9SYq8y3HrjEIyP/lOIirQJ
OhyF8QbuhjhqXuqsJ+Q3PJcZYmSMBWAc5bMuaQ2A+YbTWWyqdplDlg5ZJRw69dY7
+VnV6VK9fjENhw33Ln/0OPvltQ1YM8mC9viiQUzCZA9Pk1vO/VRVAdX2YvaeVCvM
IZD7HENpxu+0jG+8aUUfp0gDi3xtD15ntfX6oGR89lPO4a/uamVRNilCdg48OHA9
+3BvRqoy7jc2KwkouyngJyoEqVvYO8VEMFqR7z/31vURfuJiDz3KWiKKkpRELrVk
pAHanosERxq3xpRd3191XVUAVzzQa58wpejBYRzVRo5epnBsczjtjqx5qETx9LzZ
whvftYl7xBcfBcvCn5y0RnjbUnoABpFQAFJZOq/O95GLEcqkSwxzBP0gxWp84vId
qpPgc4fOsy1EtuBdTEWtYSN6A17mvjB7FgOr1bcM8v8COkVwtQYjPyyszbGoHOZD
M0bxzGpZtW0QyC9Jv+RN/tTMs6ztxi6jcUOkNyYkrCbLdS+mJvynJLOJTnKkWLdX
6xzRRgqXbJ2l2j0S2EBdaKS36Vz7DbGHVMyt2yBe+D1X7teoGbv9JI6MW9qigwYr
VNeZWgXW/HO7TZNeJDrVDWYhhS//bN5qtYDUu7kyuCAIEo9LMICeD+p8LEYwkYQ1
7fnsqbP91MP8tDNwEo+0db2ejhburjdcgmd4PkbYcvFb+bViCJKrb806nYJ4wOXP
yBfCIshrpfTBixWa6lKMbNfgm1urClkqV0R6f/mqcPktwY8Lp84eRT29qA9bWWYu
DEexU3bQeJgBYTxJfnLsELTCnaZ/ZaSv1hzGvdOata01Y2ruf1ydqn74FJvuwwm0
aViPisFCMhK6qyG6ai21zPjv3xdGR+1byE8lObpaeiOuG6Um88+q7PB4/xW91o79
2sPWULMHDyVfNtCEsU4arDaKZV3gudPZkIaj7+zJjLs2EgTN46X8XdnQr6oj8evC
HO3foNHP6CHhwfDqXrQlxZbpCYGsnicfIRMgMvBfyYCipPwSE+WBJzGsJO5jpUPV
CwomS2XxADvgDqJE3RSkKEog2PaXoQ2hZK1ZGCXfMYQtqpxvZQLGm+1/Fyrpvfno
VFTFqMQ2lWmZh77mIV8aJgAkpEYwPBHCfpuol6LyRPc0h+8Kr/ce4X3UUqwZ4v1v
jeQhjYIa3DALKmDT9VclCEEZun97MNqQwTdnteYusQ77DHBlsJ7WAYwGEICUvIF3
azd+2MchX4VRLhCn5zfV/PQAB/P79bzashGxToOq97++M65pq4iDuKNOkgxVS76p
XFzbT4y5Nz2+ScbhDvnifXHHUoYgNlpltgUSWptVO81Ecl4H4F1pnW0IgZADRXsx
MLKl0bJdTHqwhTWfwgZCkqfxXn5kSRMJvlXa4DEsR1BUEJuEMTtH//oMd/5lS7HK
oEjoPRXLvv3D9O4/LBpzBC4knB9rXeQTxBc3t/azsJ6GXLRG6eLzjnNhvwY9t3uF
cDcFSUat9AyIC3G9rGfUhUUqqkngVsPcic+eOV+23zvWSPGKKWtA7tSSOsQPgV6B
Ncz3767/JGv3TZFIaNf/zMW8NoOTNYc/bhrTryVtIL4uoH3D9b1SS9c+H69rYD6j
JR2kIXDQbsSbM2TgMkWuOLOJZf8vJu4mny7mKtt3q8tMBMAK0Kl0MBSYkAq3VzKa
RAbIly0meznJ26UHszV9oJUzRdmNeU9P1wLdnNUJeDO8FoAQ/9wmKB8pqQUECcUm
qm1yCGR+Y1YL41NsnjwLbrZO4fAWEOM6vTZv6Iv3gRQPh982XfjfhiDv70/zOYMs
GbaL8+FyN8aJK7zVDkhUjahqX1sYt6sf0ni0gna0Rrvgf9KK+nb9EILMQmbPzqc8
8gUOCgaWqqx63DT6S9zreONzHKc5WNiFlVE/5pJMlDtcQSV2+FZSVltqGcR9tf6Q
jPLApOGP0K14ynCMuXlwS+/Ibq8tlSiG8iEBCGv2VHJhowIvqAGUKIbprljmsLBZ
mXSgbxik09k0uS/uwpCeAP+mWTGCSGOGnfnR22U186T/53RKHidxbRHcwUvSmIPX
dg+agZWwNtCQMox+LHEUvoSEE+tY4ND//QsEBw5NInltXeaGRrmhNIDR4SfEY4No
wy3/I7VfQ3eX7L9pq/+ve7kaU1IIyHPhPUAcQv3aHvNri6Hwj0Vt54/o+NDPkk/Z
qF+frKp6X/I/Nt+FNwdwsWuJD2zY6zrXKWk7TiUVaLgFd+mmUWP4aNPpwA9abcao
g1LrdWo595layQckxia4zGEaiq/psRAZdeHst0NzX5NB0VW9EC6TaktA4okWj9P4
jE/KfRBQE03ZO27P7JjKKvcA4A66NssUxO+upXaEshcrAVi9J8GErG4LS3tOKMxH
edxGZ5AbO2eQDV/g+5QSHjvPxpK7ky3R98Qtu6zhHgzUpRkoRC66XzzVtjsYW8Va
XfZ4H0iZTbzRqkGrX5b7jrDzaGcJrIj/awBKcgooy8A1z4vGoknfeO9Kpg6u9fbj
LgUns5qF7TTYfnPJA2OWxaa609uJGzVpdVD53b0YX6QGzHgZ8rr8ofxy/43aajZp
nBGWwGQbxvnQVYe823cx3fokN2QSkqDFY3VY0yj1QxhNQWbvxJjpzjetnQu4y8zJ
6UHDznEeMTECPdZzOprDqdEGJZpeL/Yn0YoyZaUSPCuf50s4UekvsKndO4zN48eZ
MdOf8cEo20veiKU5e92h9z15jFyTybh95qb1sSs7bdyiD3nON9JWVMS8MWmlI0RE
pEfj3kbY0xMwv7QiEH+5dytW3LvgDzgJLnoapo7cGjWAne2umNFoL29aws1QbXUB
FWhN8/avaEO5JRXIhGjn4qRc0a37IKqbHsYFZcxLUs9WWxM3uyv9dd0pKI91Z7LX
IqL9Zjpskxvt/ZuGrUpspOz3GdPf3NPXUyy3dLY3qa/xDwx5iiVTw9iOfMRz1zdr
JvZfF0m6yZYWNWLiKhkwLLyXKw5iWLtwgP/hmSUAhLIqNT8bxYp4+F1gmV5aargI
ozTtZiY4qsOM5taQ/H92vtLwSOyuCiPBExB+14b6udcFPotmTwp4muog+eDxnwEd
fU6+X45u5FUTCEWnkIjvOS9hgGIGABRlV+Eo1znlNGXHti6vfJnX7llyMDUByxkf
cKSjYpIFBrJxgild9ZAvwHqmCa6kzEyeDn6+ZMaIMfdbbZYe316biVryApS10Nr8
PlFwrGi+0JZxD3XiSdKM+M8BSf77m6FoXFmp8GsE7kUpp4k/sDsZxk4NWcgoMPfK
9bLte/F8avJhOfq7Db9/XW2s9LyggZKV2FYYNoq7dB45SK/8hOkqMH4HaUPN12bS
OVXDOKYOIVV27uApf2Fce8R6aQMMJabFvzns0ziDhdDUPTkDsjKxCDqVlpe9TmBR
i3gQJvmplTA7ISnmZThrKfy9ionm/0z30DlU8nAmq/EuwstTJOynwfDvIakrWp7Q
ISZ350iqUh49Sk/XeHwBM5FwjULSyEDcGCTrl/Y5HBa0DwCmoW970UBd2RYbjCbV
5iYBHduDI3ztII02U4HramRK5WdKfv+WbwQTSLFcSjDW7+Wajyo6rykxstpuraLx
MFVvScdMHHt2DJ6LuNKrZZnWPRPD81ubslGSzHKwnDsQziSsaZcoEFQl36oy1ceF
bu9B4JcfwY4JeNnBh4xj2AtordIS0gVZUyWI7PlskjqAB3xsKI7rGDn6n83rn4Us
sa/8H+nNIB6qQkwIsO122aLTT7K5yCsd6A1HvqTC+169Ktynuq0GotLVe/Nm4d0l
kC1iCQAbt4ZY3Oe0TJVu8WinLrX1P3/hxN1nI+2pBwkoupEQrt9HnMbPcWGVoaYq
x2u43N7yMFylIJqt5u9M6n5nPFFJwhCnFwuQzmAoTfQu0CIQnBQmC4lgxMM+17u5
jIrxbw3Usj2UUyaAafnh2HucR6D4wpei/PpBOzPYsEtPo+UoetD6ZJ8KaYPaW40n
HCGEEr0LMdNXu64ihvWBDWniMyW8mtePj3uSEvcUpnSAyyLtocC02XHGc6PBj6zd
D9t+c9PfPZ538oriV+yX3jv++EtGpQ62vt/ftze8DknynhJrMrvSwL2F/1YKL51m
lESTsUnbCtlzpSmWQ4T7yVJF7wqoxoi9wGN+LPMZL0ZYhG+/N/vVKLIt7qS/sKdo
u2lamibOKYCwW/4peRAdH82egV2fkN0OIkmpa6AJtfdaZfoDyj8HPO6GQG0XI24n
0LW/kZJNgzS8D+5HYURGlGAdEcEK38gHcML7wYbLI6eBQMsnv9960nZlCLstVgfw
p9IemG0kTEKP340/Y23d19wU+abvsYKDRjOMSBC/b/IAwZisYTq0wIUlNFashUuH
TVRb4v1sOnG/0+47c4mbHwSh2PWUR3/9x9xNUTvxKrQQDlJ3fRK1xPJ0Jm7K4R2t
Gc7fSjJ2g1kPXc2dqXZCNbuKLj9MOaPKt6jiqlOHvNjEmllSuE92P16nXv0FXT09
Mpu15ECUPCYYkXddGVCxqwec/iLJGbFSUZXjzSihGlm9Ub+NbxsHfVp2wSF0QlPH
wZ8OKyQbN3n39cJx+8Z5Ve2zIfPK5nCt7jPgUmQYncYjnlfz7yiYAvQXbFZyc9RD
R5WAZm44VdDpMKzKrimnw8HgGeZ9HKerjZmkDjxSEc1Wr/HnxEviTendnnqsC4Oo
GlZJcacVLxigPwGBuCKyRDqe6C3DDA1KXWFPkvSAj2o3Lks65e5AEOlKS7VyJmlS
T8lCjWgJeUYvYoBONXVhPgGei6wvg+4E9Y8JlQjJg2MJbmMfXqerF6WF1i/D6rzX
pYq9EDe3ORMoUPnAiEVXUmIO+xfIK9OuON5DsS+DZlPFXiu7+7IBMDoOfERwwcGG
zVbgp8eTZUxa3TuzLyWsBE3lMytxgJoHdvZsgX6pIZmAkzO80uK1k6ZkagSHjPHJ
Rlug0RR8j5pCMCRuyvHE/7rIXGuKZPZgwPZuS90OsRtzywMNR6szynqOnxGt/g2r
d/mX5sCcKokhckkKw1ob/zMYAWoVGoKM1K5UxZqp9RbSU0uu9J70/bO9wpdeOA/M
9kcBs851wMzTqTSeSoQnVlUPKVXnOqvm2qBEN7srWhcx2Ibrz7q5SeP/FDElfGV1
QiGbIy+QVXfydmfpZsCJQjw5vkWTAd+VL5jh/3LwbDp/6OioRrUdc3RBVhVH7J11
9+njwn5MzFFJ7xFECHx4bLT5SFRmRGiZUmasBOYrdr/2zmTxhu3a0jUJbpUDbrS/
K1yY8pzEay2k7q6qecq7z8UPPwN+iS14uUxG6lxoMi/4rrED+3pxhuUxrKo2tWij
EINebx4ViZSM8J8qyljRSuMtVHcSVaeZHOj6I8VaE9EO4WaouGVC3HhFtG6DktYK
0QG1U17yAnrgBRJ4XXZa8EUYtXmOZgzVR9DSEmGPYk2VlA9FcHADhHz91j+y/0fx
Y4ybvioYz9dk0sQqg7rn1Q5o7P3onVTivRx9Db/TdeYJu2IWqtV7nk1w8KLE4ox2
DZdaVgy5iR4+wKw7hRh1NEO8YFyp2e5XQHfkyYTPxZCN8hoRa8HEgGljyHOgEi0b
b1Kw3oyEXfeztDMqJOz0pZC1dcVDIrBuOyrT5TT60GVL4M73FseJ3aC0Sl/x4d0Y
nX2XA2GowfwrEMpu2dYBpPxN4V1yUu0v6m1O73UeggdPnmgr6dsXlSIM/JNMo9nb
kwzQT1NjvjqMBlfCVgV+ewxwCPO57kLS+5vSocqNGd2Yp9e/fINR3zX2TD33CLku
qvmxWH63b5xz8DT7Ozmaip9plZ4B11T75OioI1c9Uf/v8SS3Hv7EPlxIa2XXQdz+
pXdAChsecLnkffo5OKBzSnOuEcayuBC2K4RdWZyjOKH3IyYeUioTNzVSe5jtXSPM
Nd7XVUSMIEsZcIcUhcua7g0+FrtEpeLaxmLJfkoVL87cMGIlKKoF/xrpaFMMZ787
0S0KeSB4VwTz+rDmBuCRMJzT/hs+fsaeIOsTkkK9q8MlHs8w0s3HI5uM2u3luvGc
aU4Xt/MF+sECbAix7CFLhyk3F+o0pNi+wXN5347iPsVYK0USasEIh0rf0KLR8/rS
C4P+GVGJiWi0jPdJcm3rN7h4BLNInmpWj30avwp4WyP4tWaBbiT9BE06kfkjxGKO
wo+/HZI/MfKoCHb008Q6UzTWLpatodPxFDQd6CeHcl1fwSMgAbz13X2VFnK9YfxT
YjrwahQ9VzAFKyZIVG5lJ/SUFRUHHoufP5Tbgoyiew3DQ747UXq9zKxhIuwr1ooA
LbJfAqYTGib5Si6dYEjETzOW7TmUz5R2sH8/ggjCmXYJskGcza8wTo0MrNv3S9UB
U//3DRvKvbyKjiH/ia43Nh/LwWYGMWBb3SHDb4uCSOCCq3aXUBEib1+u6P7gNSar
EbUQGXkH5V3sj27ry77XArZcSyvmeSDrPRchB3rqYNbXxvo1AGJQeVLv9ks9zeum
HtlLco25UDFkMEIc5NM3VB1lr1uyAqhQ+swieXt87Owx54ngAw/WUzX5CR5KJ3tl
9SHyv34TwYGocD64oOpoytf2AVbvQzx1vO+fl8sarlVdOyC6z47m1xlKJESQhh0i
fxHqk+5tKwTFT2pFi640BSwkoGDpmFp7mPfd1t3zeKRCD3DGwWAYzodc06D7QndN
9HQ8b3bvtU8bp/4z0ZLGtZxNWcAY3e9kjxDXBXVwa+y5Z1dBJGsh4UzhstQOqI8M
8Nm2eBQsmL4vwft64lYDg5kSvBtY+xorukEIAH34hbL9IO07xvd4rj6XnqCD4PBL
0KrHf0BMeo/xCo+9jgBqYkMhfODJ9/2LsOXGZdLLC7qw6HkoxOSmOS8bkkX4l1Et
RgaMVzFOJVM03rs9KySs8L7tF2zh64FDnATpIkatUzt6v1OAbx0oOpF3H7O7ENdq
jzvDkE8JNB/8dyYJ5lIBI1EGngrBnY2vZ/yV/ggYA94GeeQNCSO1u9HQFbZVSbjl
qbw0SMbASPISiVNGglCF+ZMJ+hgtWmFPIG65RsScOzztlbm8GcDBmUegwZmdUggW
hxH850XURvzhYob0vI+Tn4uwCTToy8DBpN/1v6Meo4Wz+IuGFJJJHRdWyWFDO0Xm
nLDpzlvAkbhEeqbeHQvj9HPALFlnAjpWwSjssuFD7Kbdgaq9WG6jrl3EO8JH+VtG
riMfhvMFmBPJ7t6OKPErQ0CHPRpMgl3xy4RWi/rP+LXwWCZKRiuJGwJDfDIAPhtq
BuLfGO0n2vt3QqnASNe0WJEw7KuB7GWB9UgNPCi8+be8ojeAo/boycvePOT80WPP
6CIadhCJNCz0Q1CTrwXh5hvMnaFcBtStqztZtIxQo9mt8k53f24BECetoE2Vtj8h
Li+OM1p5698D6KNdU0KMT4Dz9vKELMcfh3l1Xa4RzsKo7oiHS2DtF18ptf+0mPa9
PYsIPOYd37vDSHpIMZaBTNLJrTHbPpXTbCM6uOsn6uoC7+wAdn6C1bhS7ohug0hv
lkKDMJKZ4a5l8NbEWooLzcOmomEXeST+qKDDQy0fDYgkHPOVzcXgQRruUdD9QoUY
5G66UA9W4Mx+C1hvg06d0nwTKgmpPN0xpRA28rp60J+Cij0ruYQA8BtZzypvI7gl
Oe2fLvHQKSBHJToITyekOccORZAp0gABnOpAwAkotfXEBuWUIzcTj49nN7saiW31
7mDBGGoRFkUzx9YFvB4bzh4cngqJAvMdglXIzzyUxiZFpU/ycosJ0GWAiARBH//2
PkJgOrf07fX8ic+Ir7/0avji2SSfvsr30kTJggn8ZTRwhtjI+4R7NRy/p52Nbs2p
Tz7ADySg0PHhWuQ4MrNGD3Vsh100Uz39TVp9SyGBwYjQd7Wl8GvSVuRVk5wH1eCy
d8VZFQD4CSaXdgChzhRfcgBMUt+aNxQz8KufssulH45yRPuJsdnSFTCAjkQ+hZAN
mhJO/Q1BmHoBdsAtMfwY81mzG6EOL8egJs2EqAbJbOPRgt9NlNA83PN+KHWp/b4a
o00HS7o/PCynqmWP0f+B7V36h7+48oHQToTP1ql65uDRP7C1Ug/fvgpRKu1N4FTw
UNznfTmjPc0miimRxmH+OwiJfLAsuVNtA/qUWUbB8ohkc2uHuv6qo8XTAcIT4JX5
mxw8ItQAFvT3WCvBRhvAjwx7zJOFjEUlWzR948ZfMZ0WVkJifEbAEEVoZLGE+/NF
yzQcWsORjlemSVKWeSWqeYXR4Qh4ow/860tfUGfpQyt8yO5HtieA3Hqu1ZMnWP9O
klB2A1J9tB95v7SYPvS1FpQ2j20d/a+2qF3AkPn5nSze7T2294XjXhL76M56n3Gg
b84drIKeMoJpguj7aY6pPS5VLKGRTyU3goz/ciyNXLzm/75UIVEh5o+0y4zWNLbx
LIGZhCu7vZc2ZF+3vdiWLhx7ptyhG9pXqWA/9rKnVi6Pn3oaGOed6ttUdQZQEh4A
WpIKUGW7WBHuB+GAasKIMMmBz/n/njwV/MzIcVY+JCH/z/lGSh/nrs1LiHg4ZMCO
7DzNTP0FRr72nFIz34MlBqRUdLGsZmbNUmYmh38XF2snE01e0YkfUPNaze0oR35z
Wkw1wQAYynIIL56sAgxTM6wPHSMkcbo9TSn58mcv/zbmxkTwSxz6gxF+nnuHja2o
7kl2dWw0RSR73EgFFc0D/ws42QqSf0oiFr2lFaV78vHcBMchiYQSCX++M1pVRPLo
BST6eP2jAo1jeOG4B56N7j5VjQPh+K3vEyFV6/ikJQSk/ipwFBE86DIhQswW+w9s
zVkl4rx3zqrSUYnhVyapZywCSb9uOS+Wm45CgJUJin9mg5vQBj98/N9jZ0oEv/Df
I7JDiwmrkz6VbUhXVLa+bZwwG6ud/eH81BWEAzi9eJwIGtkYo8PkQahlzS5hjtQp
BAP3SeplncJQEBEykpFF5K+c8Em+wEY9r/XqA6hQr7EUXckVT6eRkMwIfYnhOZac
+osddd/9plL0XHwLDW9sl65mYoCtUV0gFaCTg51u43RLYBkApZedS8izwcuZj1j0
3lzpmtpyaJXGl5W6wg/Dr/Ty2ZE9B5fiuQW6wm5cEB2NHB4ZSuFXMQEFJjhpcN2T
ij/u0LaASQmZLRPZaM+BzBdQ+g47JZsmOzjqKAitE9EELp8rQHvr0XDnRjBaHhTN
fxzL9KtW6d8cRpH/+aHwcQVxdgM+lAY1GS72ouIXBrtzV1J894zbhpAejAP7PpQN
LSBl2ai0NHLke9eyPs629b9URKzR76jq7dez6iljbrAiwnQKlUAgWnHflzVZVqcS
a7F9N2PXHrNoAoFSQfc+LoT3RT/DK5pmyr2dbfkYMAoQ83JsSRnzLpyzMYe0Mdth
+85MkZhnXAZsk0U57MXPfBhL66CjitiGTfcuGwVmxkY+q7nIhHTWH8YYJqREAUZU
0XE7w268RxKezBBqywc7db953+A2lqX+3OunGfCE+mglNBTy//+3xEF2+nFa38KU
EcJXHm1M1tMaWP1Q6TCnAZRjvJ/eEIw1Tp1gNEFS36pI+zvPvwX/tMTFAx1JVAME
v5dyZhrog0ohu5M5rWkbzbnWiVfA+YLwt5WFu0Hg//x1wHnyEoGjEvR+FHBl/G5K
dgQtMjzPSQXxZknkPS2rRPyN/ncrgFPbixKabQm/aoTs2aWk+HRaJD8bJO7NFK7I
Zjnx9UedURO/qkgSGlnljFLyl41TnTUXltTtfl0X8uwyMYkyL/fgGYcXtzLwTwCK
AV9TuqNjTZXMrYokCD9p/dqvQzMxk5uDw3mIprr8QlqvRkrsZZ7+pIULumndgKh8
we0j82hBm7C9/3b3nirY5opaouhLJc1FNGU+OrFobcKH/A8D9NgrI2el+b6sPFs6
V/XczR96x2++0tztnAFr69eznaCLUv8e2aB1jEj+f1jmLyxa5E2PYpqcFcuuGfxr
T+qXwUU3+PMreBsyzQ5LQLJfXaXexqyeoySrPHWR8k8Lh+yN2HZtetB23TWhl+B9
JXo1CNKwAaPPBPvekpPcoPzvUgOnNb1p80xHVLS2OwLMLPpTKZwjtrWFChmieJ26
UjPytwVCJtwh1+NHmOqE8ZhTWFFDvlmf4tipI9ZeTwFLBGIpEoyVptIF4k31R+Hz
+ee8Cc9ch2fUf5mBcU01fope38KTLNWbYszY4KfE3pE0d0J8DhAoSd7mjoalEyb/
rEd4u11YDIqNjysu95u6v1UpO2x13fsWSUK5RVNbqTC6aWEHZjUQB1mU9wGhLq5J
SxtPz8BzyzWI+uEFlbaavchyNWbV/DOpUKwadggheQS05gpxd1H9S7R0Hgs33zoo
i3Z7Ng4e3eosrtDjEVS8bT3ubKufq94cN7HiRWLZXYbu/WGWRNTX7qxR3sIKofgp
Zw41Lrqdv7z1thgsRiGMFCCqofhqanpiOrUoLUrVJ+Q2naYuHSKL67D8tjiF1OBc
mIDxUvptvhIQhhwFD6Z+DudCS7pciRpfZkKVFlHbwCijQP4HnZOGX75udqNTVMPi
gpGnWp2se7QRzhphphpiqZD6du8kgEdKXf/lqXHk+hBat0plHHUFWp9I3dx2UWXY
Qrb1nDC06d6jvekcNEa6WRXPtrWgnx6xxyJSNfz9Nr1w9sxSeq94kJRThsYBb7nD
n+43tHKKoabnDH52UpsDxVkBztuob7ogYxzQaHN/Q8WyxKxDCCUUb9Bf+LX07lab
dIpSM1DPQsa2gqqBT5lKvXPk4m0yS1x+aKU9y1HfYFYdKei9gXiXPlwqzj8B3Bdy
O3ZZEVBU5+9bygJW8qTa3shSyou9q31lFA6qzu4COXxqI7HMqJI/sCXVi2sgHBJH
hSXE3a86F3mTkZ3IUXf0yFeq76pM3OJlbJPm9jbONBOxMLclS7DhfjAeDibChhAJ
Y4EA8qzIXj8CjJFJwpwvkZ++jq0oes8w4+uMy0YQFCbrS2VGS9cZye9CWxsJGgQH
mywte2nJVJdEfffyorRwPv7wgXdo+KUbzpDjAIvHCDhmHQmS8rj0NgUy3n7wqG/8
avjEGHfirYEziB5dguN9btYH/6M5wiu5NFW9CztlUjtoidydoYo96CvURh7blNPq
RjODZd5xnNBG4qBZbf9BpXsVbs/MyyjHQNX/5yBszlggGeBrFQ+h1l9Fq6s4eihT
q3GLTaFghYIh/RzBcWDaHFyxlQBxfDiUg5gDaAhDB5bci5NCq4JuAbMHIFR6Tjyc
a5hz/BeXDbx+3Xec7f8N/iieait4E/mBEcVkSELMqEFAdTQSbNxUMnrh6sLV3ALg
rcK64esxAaNh8DZ3by1KbjXJBdHtBx8hD7YxoLyPUEa2q57lbBqc8gwzmOtjq1cv
zNPqujZ6tH0GHHYgU8stpFO9AkeXubZsV+EAuf9TvM/cpxMEIcsGZ7KmmFHMYisY
fp/UVBtUXexfqwYIWrjlIFnRB3A8oc9Koq0XZPXw/RRpB//fp2rZM1snnaSCdy6B
mYWoVHkerXLO0P2GgtOsJ1+UWhMUEy7HQn872LE3eYuWge7q1KNh1GNLBTAVbRnH
WdWb1glwqy6IkQwpFpmTL4NjYgkxdRXbMxQ0xuy5tqjkQIuS3tluUwcXrVjGO+uD
+0Ufi9Y7OfJn6JbDYixodTnDg36ESuEfMrbDNOHSU0EKIfetJhlZG5hOJh3WqAGH
fMdZtOlpTNVZ11ZH4RrqbGb6zPNU2DFKbrGwIy5EjXGKymuYoEeYTsydfVCr0690
hK9SlQ1aQB+pomRZ9AD+QqE7T3If+DWJPZdhJoG+RBAf4a9+LxYQaUmuq1TiVRH4
YpoebaKYl/TvVy74D21P5PQXLgguki0zD2Rd00+PNfU7K276aVvp4CDvf2Gvh5db
xyEIIKRnniqd4Dqm3dD+LPa2b/8MsNkvUzk5LMmYZNPo+1l/xYQkDjVVGTk6BpY2
Ho6qNzYNl55GzARY1hBpjo5SsBU6sdyvOswJsIdj9V5x2NMzq46daHIO3whOrAvE
Nzw/Kz4o6G7x1x+HYtRs4yUHD5xsrRXzJSTuCwXReQi963knzzLn0UYXWYGvK+TO
8r3gJab/t1bHhg54EkvhJ72M2jciO+1Aq0gvOzCrm9514GHgsjKLWphqWxKMGgIk
VSshoBzJT5sEKZFvr3mP6Qwo733lJFI1iJalA+1scDMg26ZV5XCpl2LQf80RnofF
DtBsg8RycjVgAZFbhmOR2nhA+vktls+E9rSJTbBQ3AFYfqxSLODz/6rHjEuxec5e
w5afJn5DdE2t49usBD7HVOCQNe+lWwMMyypjOVuFKFvddv+A3kaaR1uHVPviq1EX
9GoTw/WzpqN8GN5W0Fv63SVopNJRQg1nAyUUUodGKi9rZvf9jsfePA9CovECDKBZ
RMgHBDne7xFfunolf4dTgzCaGk9cDKCctINEu+AOqkXrf3AMZJPXHuJCG6ycRWcC
hO6Fh7ZU5b7sGtqXfdM8z/wfCboZxv1IKIoa7wgiKESx/ZDRrCX/KXSPcznSqvlc
sdofSNxyDgR+EvTE1AA4GXDwNg15FwG/7I/QPga67mLKH0CwOgf+iR4VOBIhcfez
kQOgF3sHKpwyAu0xiK8wai5lWUh6/YTHU6BWXGXgprIdWp8sucBHOmKTehm7W8qf
G7UqSaSbkg2muFrVuaocKmZQFIUwxqVfB1V5H3pbA2zu7cZX8GdSL/MM10vtDZIR
7nxe9SunSwxi1X0AAED1Ox1/MC7ws+Un2z3dE1vUAcuJpIcCTC8Q/4qr44iyBvUU
fE+IOUogmCj8MY68YoPuqCHxpnzOM6oVWcJLrQLr0KWJMlXTF2iV20cZGKSfwadk
VDv++fXt56hjvP13HJlRC+5kvF5PF3lLPOpLo7o4oBlJjaLItVQmjsXNIZc/4q1R
Vjlvnpqew5osjQO5Lb0wrhUWShRE/BcIROXSeeg/SZBWYQu58NRQOxyCO80Y0IjH
rSp+aa4Bd4/ZShTie3UKlzZKiJAMW5KUxjNj4YGpylw3c4pl72mkdyGCFgtQveEq
V09KPUkGgOA1ADQ0SNVmkaCxaAYMfQprh1UsaXZtS9EKPrirnsmucDmXzopJPaKM
jKl/E8VisYOwXU/8R9wJajRxo4VY1eHQtKUrnvfS6mMzt1MwZaC9SKTduJrbMUzl
vricaOf73TBl98Arg3ztSwAt/blSMZJeEzjL5/xV9Ss8HYUfxi83ehcLWWmMu8bs
Af5UNBbxDiOINxQtCZ4raMNNjISHYOgZCak6oWanLS0TN5EQkFy1k1T0MsBlhD8S
q735BfVcU4EplIXCRjRi4m+aOekCZiHgCJ46Bif0zka9sjweCgQMbuWGkzOVQS7X
jEq0ptjs3v9ZXGQcD1wJPX+rQFrYZ4ul+5NAjJYkZaBdxNXK5Tbk5Unuv17UUeoA
YbV+3ph5sgHQizGqPVmI/GeYrnFyqDg3Hcr0rFom6Y2y72IHfeXvjZU7WTIhiwnd
jPfSk3UzDnurKTTzArvisb/9hf6pBf9tt/hfjg9HgxiByR8k1rBO1qr5sFo06EA/
yhNBGsW/Ew9P/VC9VOl3EizRjk1mfyglW8yUktaaRfSOYLSVenUMN0z9KQXTvRS8
ZVn73EllCpHl3YrY0b+siPmHq5cq72Nqn5Am5okDd+hzZN7BlZae8filkf+x4Li5
Bs8adinMmFmBtAtqo/cpWZo19uyS7Ih0Igk1oC4n3Hhmrd8qHsUcwu273JplLX+6
RfyGSuC10zR3OwFdJgn4hWBvVDh5Fp6ejzYVLIzK4sUwU9ydYqQk+XGdgBy9/O8d
sOtL29TfwBjhSaF5lmeMm25/a3j0tXk5WPyR5xbIQFtGBZh6Yh89XYzpgW4QkVSI
lJXL2Z5FcI4qLbC8VISL6HEvveOposawgziR4k41DOVTZIZH6CzP0BJK6cygvESg
uTE/dgHGCOD2eBsSA7rYow/oJeiF9gszhxNRUjHSlmD+/kOTpcmL3dv+wcCLZhSC
e2UBSUOMWyouEasEvi7FF3BOwwBVCwhMBKV4DXwNTKtoGv2q61E5rFRmuNbR3V+X
cPjfUCtKUSTH5oYEbRrd0BV0+xW4wflIaV3/vdtCOWXxA6aQmRt9C4FtEZjTT6DK
OeoFikZsOT8E5yHhQwOq/3T9T27Oi6vpIdtpmyXY1/nh/yu5LNpc2pOLHZ3AuJOx
8T8TdJQZ93u6O89E+mfpuNWNpkCWZxZOYXNoOxxfBzav4eXhqPaEs/JNgEsvTv2s
7GfRy6i8G035BKkiBjWy+Czp4o04khb7XidXzNaY6gWrmi388Tuthf5Qh7WQMoWx
MGv5n9v1uE6sTiidYinfRA5zXjjpfQKqiYybmXiWJs7GQqvnrJPXCZc0mKQmQw/6
H98oCdHfXTNubTe937Q8ZIjGL5Eok1agdacxbyMmP+iCdehUiAG2eQdCSpjlaN2s
ouYbQ66t+029aUxvn44dp1E5+okXMwjiZ9h6NHYS7XBkdicG0GFJfoerd0B1GAaK
awcIo7PBOnGg8fvjmr2nx4HUKQ1gRJCPyUv5PB7WjZOwb0Q9eHz94kwU2tM9wPV4
JYT18BwN45Zc79vmD1Uib+cvcWNDi/RzTfxR5a3tWtjv8E6TaONrrhCUdeR4Ucpt
Em8ZPjEeza4dqJvjju3YTH7sCqg1iURxPM8WRjnNw57D3sE9nylwALRW4d4qd/jP
hEG2/4pVdVvG/G93F4WXkeCMEsVhc6InaZe+Qabqsi7R0MukbaSOXI5DeqeMCG32
OwfONY4vFW4+QtW/i/TtGf3fknsYe49BNG4hIAT/ZkkrnX20eZtNgyGpg86WjjOO
Vnc9JULh/vsVzAOEiTkgII+S8JmDgdi3wNjLmp6TfKhU760BMrBhP93f/KbN19QE
UBv0js0NamP7LKVb7I7fCneopUgbqfQ8oT9G1sm0JVH0yhSBkDDD/oCwPNFHoBrt
dnr/silIWzw2GOtVQkd7tBclZNfExhuFyuilzyufcs0Tr6AN+aKnSrLAGaX8Z5nK
oxXTEoLZ/oqazPNEeMJgZnujMj93EITlKa0oBv76YfZvuA/UV011wJBttTtXPRDS
Ojl6Oj+mBWjrwyRKVZdQiQ8GTlmz2tPA8Ld2RBbpFcdEoAb8EF0gt4ynpqASOusg
aWYguYhxDyfvlCY3VqHQVNFA/PgeqTkL3TnyKF2Y4TQWgq6YhCPMQGe+e//Ek/Xu
9fMKjVXECVQxgmp9FuqnBS63Nnof8/fKF4R9e3Rd2C8gf0PWda0mOaiuOaCawVKv
Q81+aI0VwBU8sKKt+PDC2q/z+DO0aD/KFuEy/NymmJJDB541AljgDsjHmYAsQ5t3
tdvntSudCTzOsa341g2a4xGmGrVMSDaXAYHTDcB/JqqgpYSQRGi1Mc9uqzsOG/yK
IbNihaamGmC8b+OYy6Lh+beGK576t71YVSdc0J+PmrsKZyyqqBcKgQcwE9wywKZs
VQrCUMUuTKTZcfdv1tQzltrFXkyucjoKlyKW+4T7+0gqJe54qlFMS8CnnPa8NzL9
5y8TzDPZ0Td6Op+C4IRNR73eDYlP5cML3dzaLIGOj0kBtdGRaaLqdduwjiUTwgnN
afL/Pt6y0F0Zk6iI8abUwEBWyfuccE0lP8PBMkbmbrttASrtcShlW8SrKUvCA5HU
Wv/duy4LcFZJxtH2cc1nbbQXSde0gZp8vsV2UWK8pvkSQtAeJyLsXUpWboG7VkGf
m76IpuwocfGsqSSbhEsNUkwnk5FIacr24xPDi+LtpRwdoA27yO8qu9gfCaGvDdBo
+te2wOUtAuTiZJMV5ujrbglKowPMdCJxFjBP1gTwp4fi1hNRz3R4Qi+E5b4rNCFP
pQ0KXtoXMvmUFQo5o0E9mM2dRQg14Q3ZfjPj+u+zSmPxCsNNofSl1Af3+0bVNr1L
N9rRUuaqs47Mr0pFRROSHjhuHkLvckO85hvsS9jm10LR9QgOOhSinARvIbRBJlWu
iyR4+51cc5N4FMbAl/zon0N6P3XWizfdy3OSwIP/ML9YyZ9yTXCHNTr5icZ59ajI
Z+WjI55Ns9b9MGkFRyGnF02D5txjYCUC+vFBNGqQ7Ye9P26QC/074JuKCeTvbtF0
qDKlTGEc8GiVRACa/jxaJn5TH+J4SLn5mYGyZTLiV8otjE6Bl7q32F7BIQv9DvwP
HESjjugsbdoYJrgBSFpBY+uRP295iIimRoH4oVCIMMSDnAHcQw1BN35khS0HNbBm
IP+tpbEE86IqRY/1ABDmsT/wrr+UjWHyN5elCctMsJgY1Y4wqOFIXpJehN//aF5G
/nP986/TvLt9K+hNu4N7yVg+CkmIDs4rdhepd+i+uNtLVb9PQtES/UBApyfVJbQc
2JLnuY8Dn7cJK4xwS1AW9mEOeqG8Nmct+xZL2OoQnUXEGkVmdOJq1Fp9FYne3M+T
SSCdu0RjiuOFxsv6nKTGtM1JASVhYYyLa+Iq17sZaW8Vyxto5OS6YbsWN/DA12lH
3WR0vBqrUcE0WuYRwAFz5tcyV0GGT8GUmhKb+VGZ4qRr/dn5zgYL7dZ0YHpuV32a
JIKgfrdniJSQokDtQoOxiT8dWnz82Z0gdEdkhqB21uMcUAyXvq4C9FCE8le323Th
S7Fbt+TpljeTICJf0knXU78DXMlLKv6uoQ4ZcpZnBOJTIpN8BreuBkODT7dm4esa
LvpqmoCUBcakohPxOShPD2UXrQw5NVAMhlaFTTVtY5u8FrPZK/8ndSHoynNahzS/
kH8Xao+4ZughDGtAI0iWiz/QsO8HBq/VCpi6RlkLLJYyENePc17rZDECE0HKpunx
AeB4oSqe+ybm68Ez6RUsHRAjPQO5j2xKiRCky3Sn4dkPdhujU4AbpQxyZqQVPDxV
U/ZBXOgqG+qfa75yYJjv1fkfUntfu5bKx1iFgxxYTw2hz8vgeOsFhNyxb5sz6RSS
BiuiLEeOrv9njQI2mMlgMWeNZkOXE7XE1Tzd/FSIGoEW77n09aVZC1aIKMkRm4zN
v+4zXXSL5tmB1ogb6h2dopNm93GynbBkAOEmKzr+dJLOuEoYju/XHSioFLP4sOhQ
yNvo207Sx0bD+CZU6XI+yvAxyPHX7WXULcvLw6V+jskO3XLZmk6PWn39hFxbXmqH
C+zseOrjLWKRHuZPlRhs0xP24tvOw06OLkRCm56fcJCVWjjKAMdWb2gbSXzQkkp1
kN0lJW7FYltcefn8dCxAHXIuulJdlQ/7wDbSZwhomOmkZqZ9f4tcc8wqpTGBVTvr
tZahj+FAuuqjditSFLXpvyUyMbzIO0Qooav8uBZ9i5Mp9GBNmVHbk/93R8Bmr3HP
m5X5ddePC0nbi8Jnsm4DcnqzvrVD9gWc6BiIwoi2sTDeDni7B916lhisiAqzYoQg
+Swd4h6lSTrKk7ow833p3virRxnaNHjrySD6X5joXIdIa0RqBW6wUdWbEjCWNm+6
cOYbLyfUqX9uW6Nr5DlxE+rUU8aNcmOL66ZylQZsbedG1Lgu7rX/fvT+UnmMuABE
5wueBvdG83Qumhrxnsq2yljoxFIMwQzmLUnsYMCzRkcVZsE6WveGBUBopT+xo72a
UERHaJYaThiun6ggMyGzEfKYTO/DFVLybzm85FejS6+BA5OiWlnczxwgCVp+KHJE
YSDKlUvEJIdFcTbnG/mGl2OoG1hTJitPnqsnT7NP55NlcjVKXpUkMA9S3vvKiEnc
Q1zx45HZIW3GC4oDi4tSCN6fH7ocYiu3/Cy/g0ckaP8b7ZL/B0aYXLNVN/VJzEw2
dtS+KyjmknPlrBlGoZ9x31Neqv/NkBajig4SORWBr09zhzYHTkOh95/1aIOvVQXN
Osq0kWqrokUyhRVFCXmt646n1AaxEisxhWHgqDMPh3vrKv0XPHJOStsmHUMmMGZs
u5YR0wpaMwmVp8EpXUlTrPonDsXK8mzEzCXTRdMpkXL/g5POVY8lAQFf0vlJTRTu
WPNCJeiTh6YwDfDR1GrgzuE7qGVe6+SVxKJXIwUCO/2TeF8qdWPsiTVHuoqLexnL
IwgEsvtM3ehqu6V7VR/+Q/qts8A+/WDmBsipEpMAXyLp+Dj/rNHAgtqgnBdoHua4
DZZV9/DOmjNg1MyQAqUTuCm8gKDupx1Exu3EhkXcfw3sRpUvwxFU/k+JTgUXyfOR
AMKfJWbD0snqi1ZLR5IiZGy3N0xJNJUhYfpuK050/WSSUL9M50Tv2UMhGibIlSGi
H0h+RBjtD9wuMFPlL8JzI6y4NL4R7Q22ewdS+1Bd4nm1lsMsh/qchisp4Epd/Thb
b428KSV3elMyVY1Yn36h2VwX4Kgxesg9+FeBHpf/IcylgDT6yZ3vqEGaEX/emKOG
Rhpb7JjhL87AhcUUxMqs3uFa2VmPiepXCCfTfJmT3J78oLLCeXacbzzCMIK8QI5g
FhYh9jwF+uGZbJTjZ+mnSfl6JdGn9wBOOthmCAlhvJzDO/QlvolqITl5uifq3OlG
5EZ0bwfoEt2F/c22pyG5Fjy7b7/QlLzx1XALlRcw+zGhJQPV/c2ogXdshIPH5Yy5
X7tc+/sKmZ2lvyxTC31Z01Kf0NWoTZN5wtVjgnjmNI6FZLUoi1MRnTJ8VqcpAm+d
qgLLAxS2Ul4911hmxCGqhVtCRab9lUuA3NkQugCxu9sgYr5AkN3c+0dqtIg4yP0l
nQHfPUi9IJhjT2Qm7B6wT5Dqp5fDsbEAXCSCScg1jEJWqUzORlDtx9Y2ETzYW/ES
krsGStFpkgLBa2ak6fxNBY5VSyf4UfwSZy1b1UW4Jhar5L28LdzdaxFXhfIUEgai
gHvHpvT0fQPL99cgu/scdKlyQ0T6HQE36tpvMBPtMfh9UJ+CR1cQyGxVYI4qrkIq
vo9kj+VSK+xw46d8ehLgLE28koo62eJuGA1T4rtc0I+hvMOFX4GqVb/xKZqz5VwY
Jbsc1+c1QCxBoM8OWqwQQRgKJpsT2WnR6zVFE3gKm2iMUcYdWVamhzKQtpI7tilk
3RUzr3gCUvhalGk1W6n/JPD2BAnsyWT6PErRRxtu6iVU8tAVT7TgWiLFKw2eXLrg
MUilRi6+zc0B+CimydMpwWJgIeGGQJwMZ5MdxOibZvesa/27w2THsPILLbMLZqe8
MU8D7r4lHU10vCaJQVUTK8X54UHUHsIMbGAUQmTrV02n3VIPeEuKCT8koEOIbE9B
ZPLRR15U/9yxGeakY3CQ3DWlM21EwK7C+eikhSXSpSgtRYPfXxijKUMklgioK/YB
yu0s7rEtFO98+jmeFRprKwIdLXRZC39dDPDvtYIW0k1A7f2LVBUFdRYQQP63z30e
++dkF4k0zyNUCx/DcFJTU1CW2TXt0+Cn6v5aZWNl0/LzzUnvRsLfBBT9JL1EDDWT
g/tdqELXUuSz2ddyto3TTEF2sFbKlOz6hhlfcE1jgrT9X4M9abG9gJwB1fvjPrlz
TVCZM0s/fa+MfsnWpi8uWyv5jvxvDcsXBs71+5vEyVXmw5lIzf0kpsCEKt5jh53u
Ndr+c5qwG4//U4vzoCJfwZwFKztV5oc6RWfPMtkEOMKt3BwMvcP5iPY65rw1SnJz
vMF5zJYPJKi0vKt0kEGett9fct5hwjkzIdqIIbKWgV0VkfO18AQ9JVIOURqVm071
QBVJDKA037WgE6oR00GcL5RlKXr1ng26ET1NSS8wrMBPXRcydwplgc6/7PsvKN6r
KdxSQxauFwDvB+yVneFcpUslEunxQeP5Ea1jvK3XL8VdeBPj8Vtffyj3iBTHqy9u
Vj+2K+6+3hwI6X4S8vALUMVFdyJex9ij506GmgLHOOmKbx1NWl/ZkR7upPk7LXxb
M5O5ofgZWwyF5L7qhek0khQ2s6gBeeq4aWCQGpNlBNI3A8+lV2dmFHSxppOCe0ev
ljCbX2WZm7IYD2KNnYCPJPiiv8CugPsMOqMJrVnZEh8iNVx4mSxxDu9Y/boFQ3jI
T0hPpWw9/7baNwh/x2YddeE+WWCC1TaxyZ0IK5RccowqZgOgH824QYU7PQgbbPcW
tFmh11+aSSqwjN7o7Ktytauc4erQRfStypWPb1h6UUKU9wi08oI+JK4G9MzQXKdT
0efexfRdB1AB00RCXwvEX5lAuXv3dXSmroyYCKCZml+cO3o2JdM/gyeGwLDNreCo
xl9urJFsxC0THqvtjkUKw9bb19JAyYt7dm406W5GMpQ/s/9kqY0J1/anxn/iG/1z
Zi32dQTiVKI4uzpcO/hRfksZpRvXJk3ijONCv9jSC4JPUcR/lEOZUfq9AQVUC7Sb
yiVbrGDsuS+I2GlNvyJOc+pZecsKj+uif4Kk5+jkytQrePZVOjeuIJ399VFerkCQ
+942x/0i8e/IY5pj5nekzV5KI9Ig+OczgToI0XvRCfyn+K3nRCMIXTi42r9XrP+q
90WIBoknwWY3y9Mj2Q7FAm4lO7gqaKVX34CUY+xkfDYiPo5HWL811wTDwmFOhK2L
ZGEZ73XePfetS6AyT2qQDO32GUkrFS9zzJL1oHqX3B+J9izvDVue/CUXKLFTPlp0
hxRK/DOojN35RAhheyq1yqCkQ8jFIqgUZl05xarKiflkjhjr/Bd8Vthh85RmZuhp
EY6hwq1AT/qEsPZnOcHbDdw9aOakK4+Id4yQuWk7VzKQaJ5Lymk8g+gSmoy4cXqP
ZtQAudkgN6qxP6qKt8e6h1XAJQuSRoE1+h5FSnvlIdo/XP5CPBlmyv/VgbXSBnmJ
9f+iLPxiH4gzq0gMJ3EzjdSB7FRBv5Kl6ViFJi1FVrhA0nfLo1wtrdzpTcE2t2Pm
Vu9uLvuW+0Bxa6ziczko1h5BGLzx1HRLnvrvmMdY7uRXPJy/1ndk2qILq0Ro0LWe
woEq0xJFcE1iQeYqXEPGOrP+ISnYEVF6P4gdn6225Vk5B1orcBECF541uPmnCb3O
j6Q93a5kwKHwlwKtAHTjXrGUHh/U8gPjl6+Nc6nV21eMSfPTNuNWEffntSdpgIeu
cIsmbQhy2UsvJIke/nrpd3BztP1jMSxSHNrYLZ6WgC2uRAD37pA3QgEq4ZzskSXX
543JNXKJo2z6F/fpFbkY7DYTRnc0YOyZPypYQvOnnERb+D4Xp7+d6ygDp4PRI/C2
VN7IExo0hJ96I+VEj8WVNDZfwJ4UI/xWL2NQSC9BMaH7moaL8ZF++PavIhVV3zRn
6FZJQKRp2DfrmStm/7e0qIxKXcc/Z7555kAG2wM49i5K0tv0yGQNzTJkl2flQwgO
FQ7X2gEtsoBLo4qGW/duee1zWnI59ecC82R7YMrc63VY9Oj/B4s0H39HBfyEkzn9
aDwCWsYIFC69+CqK2oNpV4Qnai0k5MBxUCZ6pLqtmdVXseeQa50obxlz1JORtsGy
RBL7tcspxLeeNE6a4c71MOPK3wDoJYd3gCOjYrX00ueZfCZGDckIJNmFV7dXm/OE
zvRumELbyTX8qYfoKTbU8MNXhpulpJaxRFE+56b4Gon/XTeXpg5X2Muu060Pv0kv
N/Lyy6wQVak5nT+xU5RtmD29wYFyd5DCXhX2HneZgEkPfeyB6tyB9C+vSqMmo8aG
D+PyA3vsIEq1p3jMHy5J5bj4AtQvKk+wI+KBP20gKqp4LjmuvXr/8r4+hignqGHr
1AuV00epr0f2B5fDtUSk/siZx8behoxRWE2Q4utay162O2TWVliExjCkenTLleKo
N3g7heDXoZ6f6+Q1Ap+t0PIhEhKEocBGgD2BBPGVP+JWmm3ZjTrMcL5TK7TpiUN7
jEKXv14LX+gO8hH9sXIg+QPFtMDgiaT1wO5ggNWGb7gtK0g13mCfc+hOyht4N6CE
nY+wtZ/yrrVdn65/Itj3UI3ctpxYdHVDUqYq3MvkeU7Wc4zf9lJTYqdxCx/+Jgxd
GJAOgdwmjCwlCNu6QnZBIk+FHZ4fZCWrwlmNoX5wWuIOg8h5AxDYcApXxQKPN+Uz
hsdrLDmWn8BugFY7B2SnA2IxO8ck4v9zV1HPlTLf9JhauNbhG18SVFKGSSHW2hKL
/WXwIx9DR0dBjFUj7fJfDjaIz0+LMyzUbcPdX9rY1SIoQTjHRTQASD3RpekRk88k
H5gI0OjGYgpnpGF9pOcUsaSjIgNX95qpOquHUATBBKoZWdekBRur2AZPC6opxTma
QW0P0xaj55EA/AUgiUtZarC0cMHIX6FBcOViW3SqWGIY8qqMl6L/6Yvjcfz8XYGy
99A9x3K0tzWYn4PVlnhHH37zIYuVU0yOkYVdl1PMqBIF42yBX5p9OWWygWEOGWPJ
g5NWUMgUf0Esy9KZ0j47OYJD+OaWsfT1UZ1/ljK4bLmcTqb53pPu6JnXAY81fsJd
ENEBlqxq2kIMm/OfevKbsLkr6BlJFkbKM76v/FMPXHyL3yWTZRe7CFG/TSF7Thn4
45QY5MGO9XhTINNYOhpg/0kMXaQjYDUD+ScQSCXgVWvPeIE628HAj9AudxtdKCTT
pHs4q2gFvhUdffd33Oc+zc8qyN1evVeg4Se3CSrJFkfhvyhZSlmfavJ9PQBkBIeZ
hV8JBDV0cFZvnpS3PAyZE/TcpoCfShtHcszu7C8X/lQueq1hraCEefLtJt4KsMPq
yiowOYdpmumNvWobJPHHDfOuHUc4njMXf6sXWwXb6eSTfoNfBntzvRzsFR91C+zJ
6cL8ewjHFc/tGPPe+gadXtM7Ef76hgZeC5FrwfzmMH+urMNA7iy//lFBjiLL6Nlg
bTbyJRjSfVReQazGwT1UAa/9dz9qpbS9Q9NcM7eDWIhiIWhm8L8RtFz3qyV/1Do3
fCU5DdtrX/7MAlyV+hIbQKdH27jmLqp0JKZJHjyS5vcDgGrKJf4Wka5QfFZZDPvY
bRXARYQ9KW5Cay8PK6K/Iu4psTM4b7zu8I5xZdWaz94Lp87ptghIEdtjxWzTD3UD
e8pelMeL7tMzXg1LGx4MKBCaoHLE+wDzJ7vGsCH2YrklmEEa/SYvqtsOwgDlJk1C
1yOI6eIzXrNFqI7RARrD8JGzMGatXFLDu0mJvC44rRNMZM+QNQeu8sEpplg5ASjs
SDUFD305PC3JvSLT62GpfJ05ZREVFdO9s3PS2pqtmNJ82IGh+vvgaLEhMF3QeouV
991zsCGTLhkuWJB3zAtGDWJy6F6He/5Iz6hlfClx4Wd0YbEdmGTRpbkhUWuSARxi
Je2FrPIfoVoMIm0XqIRtCA1PmS4NHnXJsYoyGPiDj1daSV81afHzzn18KaIKYeoM
9oE97pypcia6V0xQxFRlk7rQVW+2lTP3xBBpbg9yooTPUJzOYPd+Olx2Pl+P1Sam
Pb0iSr9rs2jtLTJCIefyzlcRErQbbiSdm4myu6/C3c0c1T9jqdBx66siFasJckl9
lse+zM0ggc2L3OSBxeuXvwcElGJVdmmzoHLx6LZJl0l9eIX+NDOxjtJCxn47NGZm
sPH4dQu4/sKF9RfpjckdXq5veGLYv9+CoSwo66PcNfJ+p1Nl7pnRCcRyVYf9avwT
I5QPhgLPsWSYbTwtH6sCrpSNLFSwjHo4RCi68I6C7gHCKjpIRL13RTfv4jb9Dyws
ky46GYEQYTRWmPIIAyrfl3Qi9HSH2Oha64BhXLcde/sgDPnsYFuOsftcgrKav//u
Aulh8/PzY8rXxtSkQdehbcn9HrnxzlT1gSmBWP7p2FrMlle7Wt8cV4ZQHhpkJgfy
CRb/ubGkI10cs61gRwEymU2Zgejupy6YaP8APMHHseSemTuKfEXVhSzDt2P51nGM
amVtvM9gt1xhMcwWxDjxE37bv8CIiXDlrDuPv2pvf9nMc/2BIaykwx8RJWPiuBmy
erIzd+4EBgyGMDx0nJoq4i0S3Poe81ktrWIHwqnQDCAidtljSj1zqitXSbJRDKy1
Hns9b7yCKViXVaT4mCxTWHkZUQ5bOxyCxRhaShTA47x6oRiXhL5k9X1bRx4C1hWw
f94Aa/uuw1qmLH74uPwz2wh5x/PkpzEwc4cQh/uK6piclE8OdT9aht3RRbf/bqwf
9//zbMPCNTgqt4U9KAS9XQiHTaSDnYvY1gHFxpEU5sXExWBjPYHabCYFDmZimLXj
m/tODRACJRuHk6vpEEDNyIjrkcEuIIch2Yk8baAtAtEtzH39MLQ5Z4hrFCUDago8
N39+L3BcCkq3/BLG2cEKZAJ5k6z9cF0N9BnG6dY1CVDsOHFrl1RuaLi3hhJM/Hkd
1siAa2tY9lerEi5vm2BRTGNZAhPO2trjW7kGV65t5CSH6h9luSwYJNyf7kEGYrZz
d3e3Q+HFnoR1j7tcSPnvQBZOtwMoTpC3mWl/ZaTTEXFQiNH3NDU+WSWScG+PsrJp
7RnZKxzXXSyzg/iRml3SnaD3MFt6Fb5yghgxlDmE1ZqYKe5U8jt01XpFaNw/F2Yx
g2+8A9Pk94+fUxiCYnw0RbyOAvx6F52VwGChDIEdejoLz5l7ZQij9GiJMFymbeZe
KT+hMrb0m+7mwz9PQl43lPALzqq6H1zayGkVWxssmgR19r2CFXlM59PnLKh0YT0o
4pvDIVm0VtgnaXuKOQg/fcNcYp92Q3qiXn4QtIyoaoIpKUNXFU6G7/1c4BwALfFv
i1y9eeN8lxEV77i+Kd+rl5pNsrPIMW38PykoR8QLOVsSZZy24Wsnl6kn7XyI6df3
DAn4f+zwGiMgpQbg/jtdUPZK9Ub1gQvBPH9SDPXuDmvZ/o+H9WcCn4ai44hcqkvf
RzrcUOjXitaFResREISg+Np3UjAc8qivL6DXtQqjtAKCHMx8yUBIrX5MKneS8Pyj
bBXZ6U9hcJGrRES4x5HFreMjA7G8pXs/E1D1RD61j6zZ2P2buf0dbTV6HFMnPsee
Dd+7lxdA3VJHiSEDJHmE05pjoxBCXqtqPG0p4GSQ1bKhb0lR3momVDepZtEAtqfX
51ozop+H+l4FeguF9f1IAQ5iCHQVuQMtGGMtYmotu74wREick2Hik+ec+QAq18TQ
7M1HLM3B771DEQkI+0WgB01mjxiu9qeVjC/nOTXmuh+DlKuSHqq4n2E49NzeBKQJ
VS9yVk/EDHDZdbJ5u/SGlbmc2sFDxbbDw+qnMfXRHeoz63tQr9cF/XCyJOcyf5Qv
v79wh1K6yR3OeVwKhZi/yK7zxW2xVpGnb/aCZ43dPYvQAaCitzbisjEafVuLFNSc
RALidwfUARf4jCsjTvycrNWU3l5UJsHzQleV5KHzjqAq/QIvy2uhmUjD48KNFEqE
ntIPCUmctabIhPEq4rk5ANeUzaxVJ+Ycc2QlOAExLeQ0ICgfV867VlLejuKvR7HU
42TM8iWzhQiOHdqxCHGGDwf+pY5nupJ5K/Z66KDEKKE36x8/r2xOYpjmsWWIAaJW
mrg676cLLQDopjJMk7m7bwI/hVFqkdlMBoGafcGFPP4+1qigXG41NBV8sxP192kB
yR/+m+3Sxrxn76hzcy+LNN4Jz1gbo6dpjM9cyQv0gC2u9paxGJgnUIr9sjM3+qqd
y7ADC3U5Tt6eD85woJBA8FbD0K4F43JKtswVCyB4G59TovSCtOWK5dwbk/BKkEJt
B/8V6rGwoe/rlUTMw6zv5Vxn90BdvC+zynYzJrR98GXjX3TqUbHnkLBZU+nVGENv
Pz2KO7koVBmM/UygqyQcZWuBQ3XQ3FAY8YlpyJRvNaP/gfdsL4a20KPvBR29JfX6
0QNh9p4YYnJQ1v2uWzEAD6gr7maeVRfC6VBH8cBoCttjbFWYgaYrhViHrPyPvrVD
lMF4dQtbakD5nz2BwmlCPGJvRvg/e4Ndnj0RnE3/MxDOpPLJ+3VdyHvCbMe1ViFs
kTU3IVyvOMpSvLoPSYfTMw8GA9284si03lY3WNO6PK3opx2bdosTTFTjTCt4rjoB
pCbu3mi3IlSVqcF7O6fTTA89bKdN5wCkZsY18Nac23hYwi8J/oSs2KWQ0ZixpnLx
fKp/Ify9f7pk2MjLkpUjY23CyuDSs0Jbr/M0cEfDBNEw/p5UVF2EkZrJ1a1VwnyA
V5YKCmS2wkNhjbJV/SbISPsBEyVS6Io7bZj0pPdHOrC884iaWexg1NfqtRyOAtbH
qDUTxEsztoCJOT5uIV6HLidN8SAg+LirewsNWIvnDhKXMR0f5WYBnf1eWR2gu8uC
if2yCP5fmuZn2v341VE7CbAKMsBzuNTj0M6qA00MtfHcSLghiRzk9zc9Sn2AGumM
KFnT7XhUUpdspYteM7MB/KeAZkx19YEot1zlVdHCag2JpDTApzz++e8g2sYRCVSy
lJ90+uXBhiYmBnHzvL1CzYGp9AqhpnBu/hNGFM+6SImy3K+fwUzQMh9AvtPqIuUQ
Y3GiiBmGqm3RWZtboE/N6ufvyul3fDwv+Mme2yKvemR+luv8FzVyESyPT/8562Hy
t/HIX0fujXuZUK8kqvYAuRKnBka7g6IEmBcptZEXAdqwIbrMDok/iQwo06xt+OFT
gG1U/J9ta4011FzGdhfa5CnciBSK0LLQO3IrdgsiSK4BIpY2oNWSs2n5sjWZ4cbi
LN85fgwtnfHkNgKmwV4Q4K1kFCEVZshECF4Rlw1nIwCXu6sMptOrUygwHcK6ChPW
q3nfUUGqC+asvHrCLXkpZeC+ZedIPlbyBQL7kHyLxkEySiNJUfOW5wh2Nt7l07MV
dj26iLuBGPtuCanv/1jpwVZtfNbBQdeocGeqgDTyWQWCNDzEKkiHtX1gC67Q/Mpi
1bCumu+E5wJHXtzloKaZi3uqBjuEWl5PPRP7T1DHwV2xzrcsXvbRd/f2D2Qeq8Tb
iKcZdR/VAVf3m+62gPXnHRWlwzKLc5tbfu1R86QSKl7pk7zYeVxU/Miw4MP/wnYg
6jMQjojIICrK34aVFazhiuKklTxt5R+6fwbfpO1+MJJ01ok+AX0HUWFNcXDrRxcC
ltJO6+5rm9WQLWtf/ofpIut96g84kJWlVymGL3O2/SimYBgv8BAE/nmce3pvBf5S
VMDit+UXjGkaaXoAHhsgNyxdqQGsLe6qm8lWF9pL1XSwi8h2Vhj64y6uhqUoinr4
srOVr6LsaJTYWa5yZ3tfBX8Pcl38TR6kMdDz/Bp4iMMF48eJaVALctMJmEwwS0Yk
qqnnGMfIdO4Z1AzOudSQ9gtPtPXvmqxsTBHB4A7J6IAPo7LdW8K+bEJaA+ER/TMf
Dsy5mhlb0L+jTby82njE7eKzHpKFFV26sxCUIOySrt5v9V+pKSPFvzJdettCxlaG
VdRahGfchHQtYpVVgLcjbPNrVYuvx4dJvxfY3C3wW+BbpXDLvjbdXNkP+zMgG0wd
LId0iHhCkS8DuaHgb8oRzRQWMbumNwTJ7WyMad0pc/7mws7cYOXmvREnv6e6WTw7
CVgsTXaA9UCRoE1H4qgu2LOFCqci8feicdhEvaPkNfR5gOai2u5W4HcxOCYnoJKS
an92NxmzNOG/HiXJCvcIbKgCFMi83mEUjvYX37zWyAqp0309Kvuld6owLx6/5wYV
MnwdE1/SnJ+YIiZCO5LOhAmSDUJp/aqh4kMYF++HyTc5fHKZmCBv3CxVvp3K8UYO
662Aj25DrmAXDQi9AUt2JSIgNFFunqXTQ31Blvu5A5c4SoSpWfF9ahbFSd4b14fX
xZI3l3W3cUQCBAISOpbXZHcBN6zdqIupCL7t9rS1N1utPbVTFX4F4btlCHyyOpaN
aBv1bOjjWgcMDF74Jx5/c8g43FYyQeBalioWliQaLqeoer5fnVce230T1qhEwnbN
91E9/gO6jDaziFRF1OeJ+D0goCgZ60Nqu5l37NXSijG4VqAQDT4GoOS2AkEOtBZ7
aFkNw/CIupDsycSsXH0MrNWRpGvwGeOcFN3J0ARPVmdc0JjFGjnoRE2upiYDv5LJ
P3fwRb0jT1viUKolKX4cBklQ8hUZmV32Ta2ZM7d9Hx7EogUOgtk5N1odqSheVPaq
3FSM/9HFe4Nwspeh79IX/TVQ0yEi5doB4cwjzBrdLrAO5f6wDHXKL4nQN3zKFYY3
2KAJ4gjrDK9v9JZjc4aJ2nm3wuvRT9tirkey8w60TNQ88IdXHgRi/ykngziv9a90
H7d0BYbVNSSgaTBJSsucfqDD5P0D0Mxj6lPz+qBo+68NH5Ss+FVLm1repAO6qIIQ
q46PCh4UnGLk2Xttawnv3eafC+0IViJlCDOfeSg5k1m0zTgcHXeytQBTGdvAFX3n
olj5QHkOQrz8hrZYXJFrgJbiiyTNmKV34J5mFDYNSxImvRLUsskU+hn/f7/8p0ej
ASxxk/BPaCkwyyUNWRLTUTdn+C3y7XU2l6e+buYslxghXTqB8bdjhUAmnG6dCbCA
L8DiDKHt6EizFtN/7MU+zpbwvr/efqQEuE6cnJp6sUHi8zQBQ98uiIy1kiiFCXy3
DJ63CYf9fynstsEKDzI1yyAEJAtuAfu1J9UGP2+8yh+MKR0enyKfyTWn072h6UIn
8gC8RyqwY2GyS2P7aFbgydWndAlGlAZSqGdeSxE6oDrl3vaVQYzrThpaI3p1n8zv
20l0FEXeEjGpeQYGLdzftH70+Hc5S8EKv3a/Jvfpl6ETBYaDz055tje4gLV27oVc
rEQe/+Akybpwb4ozKdnZfmxWEGkHMk7STHxM5e1qEgU2QkXJ4XDdEf8siAAGMcTU
tPUFjHtp0GYRr/th4plD87ogx+SXkU0HvSDNVvwfjJuNmSRbM3V5dBZb8nTQOZij
0pgt0PyFgckZ07ZTVAbX2BK0e3wMqp7ScGfqG95G0DUiZ43jF2fGDqln9QnhLSfv
OkXQn71k4WFdsFJP1twLxnZx84Rl3KOQJwYQ4oE3FSIRfRiuLy0zu85eSRN0rtrL
LhsPXV3ygDmGeW7Fb6sVDxiK9JmYKPeVYLCzgDB3dlrbadfS1KJIbSR/1w/9EuPu
5XzhIRYVHjH2ENa5wIC5EmRUW9Ubt1AvYf/ur0E2bAs0gn30m3j5r8JB8RLlAUu4
TqJfWD46vDHlff5oUcFnbw3r32iIhxnAfWY+wz3HzIk7kArSng3TrO4WlzvWbVy/
5e1ygxDLiJhCwgPwXoxMmI+/lNWFsHFnYiy1jc4OKE/jYBQzNHBoCpnx/Mb20O86
Hlp9o+RRjPj4X+wn1YNJ9/flg1nlM2cT+mNJXqQe75HQQbYJXRV+zj+6KnRIHYjE
fMl1WF1DgqxODnCM5x4WsAbloN4qGQY/Qlk2mb57Ha4AS/WK0YexK3DP/XQU2WzP
UANrjqOCGlL7p4l2FFXMQdLORJVv/8T4x8r5e2w8BzoUZKghnYAXIMbKQqNlYMqs
LmxczE0xRuiEGpuIj92pZ2yqnNVX3mLKtLYsPumWPtG2hnjaGmNg/xVdPDuVNhFe
0QWMgYJgdVJlVmvYWXZCdxZnnLg8GUaWUq7BwWA5TBQjGSM0og5XIvF5J3foTxo+
Hm8pwdi5znvHNS6ZUbePUTq1pxdUBKUI0qfGAHenkcj9RshSuBv2t3+tmbLTJFgS
DwBV6yYBgvNiu+p/kJptQTq9AmiYFX+WH0CCfqTqAoXgNneE3zWoWykYD05v63Bg
Gx0pQ00LPtqfvGYT+/Cc69CWtf20pOv1ho2ZypRQVvrTdluJU0aCpGyNZex2vkaK
/3UmYcnUOSw6F0MIJRptbkTQKl7ul7o4yo/m+fy+yG31rYZqLTDBWDHuRb8cHpFm
sNF9XiX3KpHorAuK3LPmxFu2BP3N7IWmpHDl+0HxJgnq7qQ1iXoPOkfv+CIdaTX7
V8rwNJvIqd9g1ezeqOqhEYDIuEGCnS9mv3NkbAqdZOfCwo6S7b5+qsQtbTAhGzKH
je+QdaTvzOOCx58VrxsM8Y29Yz/f+L28ac47wpAXdyh9WqJkUJdH9LLaKxGhSe4i
eBLtwkNV6StKPLmkSnLrRoL+j5eyegYOMoyb6zxR3WEogxy6jWRT57hO0adsEMBi
xPjxo5oHa+rGna6S5GGKYIULgY0ep15fd+0Vk7HmiOJxQ1eOA3dV5sVs3J8Oh/5r
pw7hdA/2xdEupSOVaG5JTkslGeu1HyGF63vYsyeoASgUGzHmSIyQ0OwCFJLagYnh
5Ia6RzsuRdHo8b0J+J1OtAYKHBvFleMTIJBfgVMJ2C6c7sAX4oG3KPAukm+jhlkz
sjo93sK1tnkvSLWoMaP0hTQogYMnMxqzslQJ6dZXXqgmL76E+g3jo7YkaIZUgpZl
9b3CGmXtKWPsqTRLj9c9jYrjTUHsvxOTwXC6Zf3SBZ1qGYyzstR7pML1UXQfWibf
aphNPQ8HakncIp/ABJSmZarwGryn2aWPlvNty+nuxSOEOsyOw10SzvTcuCscAJcb
vubodhb9hFsSmaf7xXn/TQO3YitKhi6jVtepxw8n1zS9LEsfSzuCM/qBEFXh/vax
mNfemP+Q6rtaMsKbj8afU/XTYRM0y0l+jsdGx1AtMUkgmebsctokkvdtA1pbEh4k
TQYaTArMpDcL/w+m+9vDGVSDav9/xgwDzv98OX/KnO7JN4nL9cVjmfQSi7HC4gdJ
OpAPhIR+OWZdq174Hqm1z0m00TCM9Bam1bV5TXA6V9pNbBqLtHtfj+rjckC81IUh
Hh1PufIo3Lnq0mUqC2iBEs06alm+/Y/KgLG871gNVURqpn6WYl+h7JCi1FhY7wZ1
THLJUKCqbDFPV7ybv3YDyreQRDwEayXCZ5rwmXduLhn2+b9PLHzR2fUMkqiYJ1bt
0I74nPmeW0AYgipNTlyT47iXk7UkBGDEN7eAfyMoA+EU7r/0shZieOBhF7110+A2
mz0eL4tEuBwsm7uXt/vvuT9Ja3p396AUGRZnTdw/9YZS5neF/EFLWHgxwDflPmZs
pfR857d6JCLD+JWpF4obJH06zYIpAKhDEteGn1X9Q3hQlLVHt2PTUlC1P1fPi40T
3im8c/0homsG7iB2LYBw1A0zE5qqc7QgLuNViPmcPjeGlOIQF61bnKFFch3q5L4s
Ts3hCHvOuG+SoRNseXLDV96CwEl6R7p+xdwmbOgT8Du0dxx5N1lsKtO+CgXjWMEo
l7Jjw+g3Wma+Xtpns2sCQpzMFRnmLdZYg8RQ0JAHgWOgxwLXgP8PYb43d44owHw2
LGjBwlQH8s3O/148QgVVj1nBVkfLVLY1R7SQspqtfrCV88QiOaZrgIN0nfdvSTJK
pj5251JlWRChy4ySchjErk9ovxzywIjeqJHk0aAIvJ/7Ou4Izm+K/41jUnGSixUZ
9qVc3yKjy73zWgSx4mY+LNUqRLPSWsGIteYvF9ax+3G4C6u+SnsfQ5wz1HUTLyhB
/EjG90ZvUgH0SOZGVpTKLItGmxGeH29V6VxO+ddnJtTXDyc5H3A4JqmWB6OQ8EbM
2ESQHYNzeTYNCb3tdxkMYggJhj7iUb7rB1ezO03UWjcb6pDd+dO45x95Zx89aKOC
NIVhEDko4VhkBKV8IUA2qkcitmkyqJ9ujvlO/cRVVMdaqB7JTwCyn/NcN6YcMpHw
kkhrViEpzA7uoSaw3ONZyLHo9KEyQ6mQa0JMhXiMIsARdINhUgn2TcKupQgZj0EU
UUiDbKAKtP2z0CPJ/qbpCkG/wKBC7fW89+j6q/9hECqdHFvjvhfn5IVQNmXFXPgG
C6LyAObgQhplkWkJq2fkHFPX40JFMpUvtQliH+psmASdFLlzsVQUl+g1AGgcq1vv
MtLgW/QWR75VMFqEvoGZBivhy1uThTR5Q9s84ag+zCp8k39LiAxlwWZIJdCGXRm5
fDUhe3+aVH0FTYOgkcm3boRvUNM2gpMgjwaZnQrgcJT4/DUhdxPhAD15sqamla+u
7B7ffSu3LVJI+KubXoxNBFIXY/Jlp6lcQGwFfEiPwKinyR3hJ08BGnTUkNoNaTal
47StWtDbWeHFB2X7BQKD7Ths9GDxfc3DZHu2hKpRHFLs5GpyCCLvSuSMneT4NQOv
uaeBzSIESuqc2Jv4tL/tjn/HXRrIm5Rv+MX1tuZSFSbD++y7YFgj4udBa9RX2rK0
c1m8Nn6u7FimK6Yi808C1y6IyZNnKnShnP8jVnl7b60AJk56TNYtXZMymehNhx5A
aZ6YDSRbwZEn5EVGSeuasI0oTGE+S1I1cfwesQhMknsSyk386zT5DhND/iiZGe8R
EdBMLDPEUOvaLYwBPoD2mRIPwqzJFdfwyvcIOUQCda3IOi8FVZPM1+mzaWWWCcrj
Jd9Yv+qkVW2o6yyk80yjNYlUZuiLddX97wh9WOp0WAeOVInv2Nie8ccmlwZH92tc
bAdv9wED6t8n20YpbUXv19HBb8zDXkk6SHtVEJ6qCnJIjLtHef2Sx8bXryYyyNPi
tIeirLJ41VJzIzswsIs1nV8gV+j9u5L/jqWAJzDS9vSLFQIE+1cWce5mqkEg51nI
ksssf3bmHsRpkRxbD/7zIe3EzPGlf22UzQ5aMhSQytxce3pu4yZs1WMu5jLUHxfC
fDtfXXcgPLsAJ+HxYfbVFt4z1PxPQ36bI/igPZqxHY0cw/qO82xfP56mkVKv7RHb
GJugV/SMu3c43Jrjjk2bhGH07T+BQHGRBcqyKOVX+siIzrARA00n2Cm23Pty8S/F
mD05Jmd4TNJyETil1PrdimYb4wgTec5utXfRW+3A+XRAdozyIH0+zc5g2kQt0W+I
mkQLlkBDchtVFThOrD+fcUxlPFHmaJxHNCnhJhBQmx1scUPbjSLSaBlgFJhJzen+
nqVsXFPvsv5ZM607jNQ/i2YRQVU9hkuvycYkANETnftzxwHi6pgk1UkC3zeM0rFT
edqcKydGA6+Um/iPRhAw/F3WDdZRlCPOSOswQmBbtK8Z8rBlmnc4I2cwdWySET/R
fyU2KDiqpntPKfF9gIPzhUKnYA4fRQgM4qX0eglp1tHNEzyBlx8gzo2wbpr8upvs
Nz5yYXSH8JT0j1qcfGguQpV18NpIaGBLOLdtIrRwPxcIyVHJUkVYmx9D0XX9+MzV
TBpsInQbKZsNbclbOQfujr3m1COs5HDjxlrzTp3j1Nv2zKEgHPUW8IZubTnDKFuo
canLofNfI5qNIQl7/xRgvqzstggOtggmOnpvhLt9BeGH3NUz6M9x/DZZxpED3b+A
nVp5uA3c0+HlLeTLARym6xznR6m7PimMTZhzNcRod2X74SWn27mg+zjkraqqRRsD
xV2WZGbBwyJSygMxmjfq1RmhbbTlaS9HCUSYneVnfBNM2uxvXNYxQkywuCf1xYOt
l8r3dePEOduJlh9e+A6k3Ub/2dayl82xXA/oFmQ24bqbz9k/0eGG3px0jswiY2hT
AZuQj3LDyoSjnDCIFrYtpi69EiJzq3Ui1D0RkuksoQhaQRakbdv8NzK2SUSyyIT1
zzvIrEz0HnI/KdYLaiDcbU7vov2g3WVnbZ6yORulAHI/M6g82quguoojXh3otNzA
YlB43o++nyb8Ts1a180fo1Alm8hBHxfKNCzYv9sanbvoXcwbnYt2UIgZfcoNl+ml
UDTSd92lqEglZFwHUYKwVSsWzx8GFwV3sEoKQdM+0sbpGVgEi/5/uuYNyXPlL1oC
4Lt3YJSw+dyJob8SfYpwKWYoph40dkIY2u5vu0mBy4i5lIlYeQq2bR3ojHpxUyGl
20gl+Flhjjdl0RBfdRqXH988C0FF4VqJomUu8z2PBSG+FI5FatUmki7aoeykx5x1
W4BakJwZItHOA4pKQAJ9h/qqMY4nB7wfNa7uHRKWNCoOUGByHkPPxN685a53WRPR
8QzD/I6OrStt/pA+0bz+rLWKSDzoQjjmIOsIeJiDzrpFpU9UAl0sOVZq+Rz6VH1n
3P6G5pyTwdPsRTXILCllflmJb1yjR085jWuzYhLnpNnEPNxUaEhMlTDM+vJFKvUW
fN9/tv/PvrXTvzU2nyJ33ycfjFzeCzkQp6wMnsPIiVJsHv5TY7H0bwaGgowH5ncH
EdoxUA2QbhPTvQYKdJyv2breZ3ZysgbC6U5kw1DXycEbFiDW7f0mlrj4bOz22ewc
8D93BUW5yQbioqVTtDxpXTHGupAaaCeFt50sXCZu2+AGZ3fB2sOQM4qY2nXPu8J3
Ip42CLS3/MXJkvfWwb+q+5J/bfI6kchvr7GH37ClQNtJ1B6qtxsZptpvxHNQpMU3
U+ZyNrwzmW5AvgjGs0A1TBZW3DjjdOKm+mwszN+Iks/ZHdhOPzFYZlXf9Kavno/z
sf2AUXFUvhM/l7OKrSa6CYe/QFKEAp4db2HSZdBrcGPS8WSgYD0z2h46EzwSFQc4
0oMqvb6qrUIo+nkMVHWVBFKX69NE0xDT7ZhSZSezxAs/O44JeM31dSMf/Ls95caT
QmUKW1Mlw803X+Xh11xYbUsPd+GAeptwc32oM1BfHY++amycnpn+q5wNZwnhsPBD
Gm2fOUElvXg8/M02usatHh3B64g/CZG9ymsyPIn2Z0bDmLKTQOiaMEDL5r7HpbcT
JwnLFw+ESS5n4M1ShfUBE+aDc8fSV8d4+ULjwi0cTLBL6V9DFIhoRdnReOw57ohg
VUObVhufnUmFybRH2xuk5V+YqMbv4Njl2eoa6EhHdobcEcmCMWXwgwfVuS/Dz/HI
WOY4DIjffvQU58ajAL681tlyXoikxhIFcT5tNadZsTd6k4ADuXfa7cmuwCB5eF7k
euRjsE9mQDiinKQkS5y3M8IGnoIekNtQdRZ33uy4viiPZGElU+mX0m0ZSwB+eNlQ
DdAPEkI/cvdT1zC55rUDXI7zi3d2tM5y02+LmLM55OziMVPyIBJbJBVNZ17se4yo
yZjPTfREJe7uF6/zn/ZMNF4SjhQZhTAwLMi1TLR5DPfeiEww62Npbjw6Hw3uxJ/I
ilE6JfoLWvpyhnzQJThQ2CXQIJUWd/adpHJ6HaiUcfk2yntaHG0mMO5cCPdIg3A5
cVlxl//HjWkGnl8PeVT50P0Pr5NZU9Oq6vSMF92mJ1HaKImGKmaJeUhvoBlThlIc
csc6jegDi+ndEItIGkcd721vHQl+mnJ9v3IXm00wxt2PT4Q2pUC66xKJ3KV0D3Ky
oxrmhK8a9L+Qh9up+OYuzJZgeB/cibRDpiG119eynCT87LmCyueskuGoiZxUiGH3
f51BMx2arEGakqIhV5BHUMoStxkQa4wK+8Fz1A5wTf3LlaX6OPMQgEQlvR5xj+PQ
cSSzVZfxOvcMNbpvK173ZSt7cfWicbPZCW9LJRHrfIP4ZdK7wRuYvl8Ucij+aWqs
JrUgNUyWKHISsCxcmacW8l07q70w9OUpf8tC0eMf2yVvGQGCoPMur2gAVSKTyXdI
8MZj5sBHdggcagJqxvB9IW7LMtOcmNL3zkblf0CNVLIlQXK5MKgDOzIUkifvLyJV
xxTD3pWZ51H+78dKDkpNqKV9xZuWqN5ppZgw5HtM/02VPF+RwyLNcA/AtCyEcSmE
fMlJzNqAVPCq2/YaQWoZzSgrv/CtQx7DpoLQRkuaRys1NkQoO5Lbkxe/4NftQzVt
7fv51oZlklIXO887y8xL1j0oP1313jdBZPOWIUUgzFSWBiRDjGTJZPVx2XxzfoBy
eJ1N0plUptaDa2A3McI1pLCPYXzNC3EUDemgT+ypIdVS9jYxSUq9O2tfdJ6qPvoX
xq+9MRnu/CtxswKfvoBejFiZvjrA2XMDOH/9e+iqMfWiw9d/L68DgxLMpOn4LcpZ
iA5snIs8HMVLJYT+eiwwNLMVhGQIzKvf6t9hIU1mApJKcYWrtlzs4MA4lDiCdBn5
WgeFiKFVhdMGRnE4bWG9nBxE5Gs+ztokcScPVUHdyXaK5+R1g1q1VWudXV1LJn+o
lox8x1XGaWXzfWjrgvA3EDezq4lr2FFx9CxXpLsefap9trClBFKYW3WRb15jEa1c
24Os7Regss552arFv/g4ulKuUa0RoRMzoOaAF0pvWDzU5BwAJqFK11Lbn6RRgzJk
+D1GF5/ltUp7jvg9jWmd3bnUPSfoj/8FKKZgVzWAXGmBTpAc3Dyxz0eZD3g2n4uA
4NW7a81ulsqB8HPfiC7rguGKPj/CchX4Z+3UZf7BVroxY4eYRoJrNlGp3kAb87/G
L6GHWkvJ8/Q3LQ3+6K10xZvkxRby2WdK3RuP0E7Kxp4RCLAIsga7ePogq8sGOVy9
bIGH10h/pw+8sWIn5kIkLG/T9xKvocuy4YebMwxqMoTUO2kGmCxPC4ODfeTwHKL8
1vyDO4aU0cj1kfgXMmy+WD2T7Gryc/r9Oc++ZrhXCbHMG8dIlUXkpfM9quAQ4PIY
NSm+izt+eH20MtzZ9C+SfdwUccUQoGcmiCfQnAXA3TZBH/c60IuVkpUkCQWy9mcE
iFpwklxmwil8tH5S8BRqSxWEZt8O2kWpA3/VhafrloqmDFf5k70WBoQwz2nNNSkf
nr+d/6Gu03FxWHzszbLrG48igTibx5CLxEwfoq8+OnuDsv265Br2bmrpG3vtpOBR
Ibmf7KIqBycUE8oqk34aDcoineqUMnQlp36WLeEAzz+wTIbqVG2gxpU/3pQuJ9+a
YPRXOBVhhoKRJcDm7P4W6lvrtQxFtNfNjaR4QxKXW+hTHWDXsyeYio/EHr2emig+
ABI5BB9yd7zn4KLv/QbeyiiSdIJFLfQBV3SgjjmJ8i4CgwfmF7smgxSB/5Rdcxtj
ZN5qfroxrKzrRzrInD0xXyMFMRMGDO3b1LX2fGUeU5gp66fBYUzYkN36RcW5bwqh
trCRrUaKT7niCc9KNQVag9mTKW7z/sTAlNBS3IQbu/upK+VbYSdmk6Qf+MQM4vHk
w4ndg71J4nrgSXfYBXW5tYTg37+m5bkYR5M0tsl/5VldEs+KSyCn40eMnRhenE/K
2Ree3L37xvB2O2BoMJfe1CAA3FHFm0txx+N4YA3A6TCsqr/nJ4sr4o0eFM5KeuWs
FoFkr7COZ/u/x71V/ACX4wR1x/KnrlSxtdO67vn1SAmdNd65agvEwCcXtApOHLif
vJWk6D2rbdUYv8l9wdI7tHGdqdvL9ZuphDAi06nu9OgLno9N1ThLHTDlAG9f9D4V
e+F3zPS0EIzZZp7RSEcGwIBM7LHdgg2g5l+UQ1Dqh4zHhkdEmVMv4Fv2Ib0adj8C
VQ7nKMmsirXOFm2WuOsWaB6alRkC5cIBavQACOEi5GQdENK7jyEndQrvVgrQ2f6n
goCqZz3hCw9Dy9Bd06NfTom1C5347rdg+Ec6s7cqfH7xDAld4j6TBTdVCyVBahlQ
wYmxsLKAZlLPHChyzkkloNBIqzJgXF0vJOZy/ujt+GhE6aq1Sj5uN6J6NLaQcSZC
+SFlJJM7y9w/Dx/YsbQngJf0hR3oD5HpldMFmO16t+8lKOjmb0qeZbSY0fPG48qD
/Uvcot6mD9pMbS5B+5fu8D44dT9zzULFhbY49pUNLaB9JHi5WCyd5ha5EeBS2aWc
zXWyEmiPILyog6cG6yk8lPYD9v/CDOxgUeMV+3qRSKfDfrCbmYKZmQfVXjIBxCuu
aDWiFupv6qkhGFkJUgygaeYbMoDBTCXI/dFeVKolFZvB+w/Os6LCYLHKuqziQGgz
l/Pvp2cqk0Lb4Nz8TDXDJGO8x4ZEEHLv/nHSqVdlfroUiQ+B5kAv25+Cm26nWV6W
h/nDcxvDQ55wAZ93NQ4ch7gzHUebNnSZJBLsL9T24C9PykYk9d2Sz6/dJi8Jup3A
KA7D6XFnM2YvrE+KeC00yKqhHlFNkkSAozQQlxaO2e9touku8c87/XSEwXkFL4lr
8bB53/MXwp6oP3ya/hb5ULk9i8L36PtdNGPf+HeQ0ikh5plNqWuZ6qnuE7LJ1aJg
zRYEtO2sR5dUE2FGaywoTUHlEn3LcelcfExfp4ZmGu27IdiDbVMzKwv6oyh0J5oI
++//WG3VdBmAR8X0CabMAk1i8bVAipZgCttAd408kaoynucLHs4LofuuMqFt9zaY
w5ca7jNvtegXBBAegAxHquR2jwTxPAaOgQLYYJFwWYyDjxxC1Ux15LsHHQdVXeKM
lCj2+KZtmlkRit91QS3s4U5CO2vzUVSAxVJMWJN5GvRJ9x0ll1sARH62+fDZ+kKc
JUqmqEo6NRQ9ftF1hNgTWF3t5SpTnOPka5PCd3s4VV0mFYjMF0nAKKqk3qjG9baH
9LNeDtvPrqWqR0VDJwg43rcLWG7vNHUqnpL0Qs+1O19fK1cx3Iwrc4q7JsxDhEqo
FCjuNasPUPNe8E2B5x74u6Mg0Jt2q5QXgOLLjHxjqS9fFH0R3VOFHWbRrF+kvu6n
1qsTArtS9+enyoyPOCsnhcxiJvm27tEIxL6tOvvtS7h9W+tBfhLG7FTDKoc4h0aQ
wVepZ82pjfCz9y48OdZ+bx7JWGxE8p48hv7cgZzflu8FHPEGPvl8TqbBJUBimx8m
noIhpQWfe40MVQHwIvG9ZCN3+P0rNnD/O69taJ1Jz4Z96oJ9kSIbsZoYMbYeaNLE
4Oqx8QSkGhACd2OFInp7rQRkv/skcrHiuLEYQ7/IHA2r9tmE87kvAG0hUkGB9Haz
kkrLR60oORlPJLCr+EdJGGmr8v8EE6MJLhnnIpeThV6Hm9eRoBMhW2dRygMG/jVe
g8/2++tby2DTevUfeTq7+8FzkVTCdGZOma374mzaCQFMmmJSCFFUBpAJfjYE0AHr
755NCYKGJKju7z0BO2RYdP4ENJvAlxmIpJdZsFgcpPeDweKahmEBbLx8kpCZ3jJn
+QrVGPY+b1/qeuRyDfPBrz2UYvFb1RyF2CWkr+6rzHWqMP4U0qCluhG8VM5OPK5X
mzt2JEMb7ACpqL4RwnwM5T2QyjByvcfft01S+qb2IL20osFvTf8Zw7dtryK6qdVV
2TGGPtfVbLxdppyftcHXwcRE7HdouhptOIO1CDKaqangEMRgOjvlu17zwEKUzOAE
0iZ+7bwFpx5mePAJUC7/QNd600cbmnyTDsp63b3lqw6jHA7AV9f3xj1seMeSMJfI
DW7gZqm0GczwdKskGcHJ7KHvOVlLqFyBC+3wz+SDQc/OqfYqfTkKzJb56oIGVCMs
KQn8MnJgrOnROloFyX2ydmmCBG7ETZvelHv2Slf9PSnFpDjCZaNiD9O0ihVs4aJB
87Tww/UKpBsQCfD65qq+EoWfVmLbKKSdL2Lt2w/shloQ+Yh15mzZ6g3WsJJxhY0E
ac99Dajd4K+/iwgPRZo3UohMt7EzbfzLwihpNdXBdUW3A2itv9qgx4cSKYIvQVhQ
1W8sdpEgMmo4NAp3zu2BRATbQOkrPO1YoIuCY4U/mtR7Af9nsjLxDrIw4y48WDnV
PHQhL1v67ry/fy/akh7S1awCS70DT/uc1HcPotqBju/ilB89HIFQrrGmD8Y8iTZZ
VP7N1BZrM7F25AuqtixQFEBVC8y9v1HJAKSxmi76c5oGaK4q9+um8qMxtdF3YGZk
oqgK+CLQlOWlLn47yMlgldNQo7THQVVrn1pdt5nQCX3rAymuYNprPA3Hiad7iRVO
YtMymXKtg3sw82nqNS4iaWKXyNOeUylclZ7Vko8/LbvxtUrE9EVScKaDNbcmB+4F
MQqrhIA79YekBtngsYzeNDBg8+CZ1W/CMs/hIUa5Rhim4wTCAos73KKPoxBZmZ1J
owY+YC5use5szlyjzVEZApRIfxOFUYI/+1Yv5HCSu+/+ZgPFY7VidbcoWIRG3GND
+khH+Id3cCww1MOu7JdGZko05D2+KZsD/1T66T9AQtBvRpihH6TWNXQhHAMPh9Ux
mZgGWrLddI0dz1tbawliWGXskMqL/4yxbtQp5/Fkiq9B5fNy+cP0qsbfh8Z09X+8
Tf4tJxJrJWnbqKwvm1S0i8p1ibYfKsuFiTMK4h4mptCeeisFJHOkFwMXxBWlvrrE
TZu6Ym7tc8Dz+Dr0hh+wHyqkqIhbDPkAqcWaKJi2s2n9UjFDBa16oKrPi0bh1qz7
AWIT6B8OTx2pPKVqNynNcA4HDy8rWlEWDkpBEKBO21mr7MF9A/LqDhDG9AO9SiHd
mitYGRLCtaQly011IN0kdBhM6K3auejgwnnERgKePY1K8LzKk+G4jDgRTxxf/m+P
MB1NkMvkLBLlkAPRzWBfKuW8Ifr6Ns85ZrGV6AnlQ38sT/Mg+i6QI3ul9V3Xlo6Y
sswnvWkV8I0NDyj4Q3QlH0GDlMay2chH3ksgJq7f4Y9HBhq2lt793KWIlQ3gqV2Y
QnF/p3YmSnLLOXECh+v3Dz8mDvIm87nhgT7NMzayUA6IvICdLaT795Fcq/tS81Sy
JNIpYxjhryfXZgIP3vGMfiDqaFKYY5ZBSlbmz+ByKsml7EiPZ2eGs07XOkk8ey89
AUMwv5hc1PdSBXObSnZtHTQJTgjKi+wJqdpZIAfTQMssA1t9vfwJsdvisUgAAhkl
mqEg9cg3fP3rrj+p8NsKS66A6nKv6DQglmB/v8qryRisOxx8tmGFVLTJNqxAXDCH
AfMMY65oWhajXrq10x93ktCyR2zSOftNcHcWXQEwZ0DOgpv3lXxRgQB61DLFuPIY
xm38k0bapi9o+G4q2uEMP6lUQMFgxKOFXfkBbce+RGBN0Yo6dNMZY4ikgpJzX5d1
tbewAFSHt9yh64ZxdxlxW9weZ+EwfMGhm45sjPI7euxqTO4jcIv5REmfG5TSTUnC
oQfZ9oTIOTUN6+AseBtaJN2A9Y1tKnxZdLr1h85NL/z9g8DMpI5oz+WVqmgJyWAX
UvRUML7hUKFn9yUEWzg572fXIgdtbBvNGFzaPit9XmToI48jxMWrmL2RL6ZYQNui
zO2CwUZk6Lxgh9dVwTweXevx0BwjM5rXoNc/zbWA7k3+1GNw+X3evRalKgsZ8pL9
jms/MuKJKUMwcAwsSOuDBdRjbtxFP8Htonf1P4UEdxtxx0Adv1zupVYJMyn5Wd9/
Z4PQiPSs5Eaf+7ljHLfpq8tXJfMnRyiv4oYQcJRNssSFwA7vUcG3U1Pk9G4RUAjl
5NakfrcChooeQiaXhdh4pZr9Vv9LS8iWSjqSshPjN5Jzoe9CvMhmI/KjSXrnVdAz
CULcWMH6Kg/F1eQrRpEYJo/i3p+qTgRYnCk3G0M3seF/B4DIOUzZeKX5EBb91aS9
zl+YSsaOye8bR48q+rTGvmipBRsMzmOcbQJFHtg70QNIfZSlGBUK9MYQyzKLipqR
/MAcwR6+DJ8TyFCHjOuHVbgxlC4ycOz45g2dsBrHtkPWPJci8fNBTA5UxPwdpuR6
gXa96LfMcJUkFMMBKGDDHTDeqaHK+o9SPkFOYIJkRp9zy3v28byHWJ3XOOJVylJT
v+B4QdIG6j6JWL3WENK1k297yhRwH77OqQ6GKZo/Mg5lpU7zSHtRojTl9yND3+m8
xVKfSyk7vEB0Xekx9oDCIfDhZk9FL/hlm8mulyB3TOze71gZ6scGDG5pTFMSBptj
vKfJ67NyvH7wxykhprv0PGDKV8frwmdO769fOn0MeXBOuPwo+FJVrnjLay46zAIg
ygxnd+Z5OalGaYiyo3TqwiuglVTZGVHApcqx64dKhbNwmNXR6iIiilNcxyrN6sNz
TtLTMjmiOJD+BFqsdGYZ89ymlxmSznneSOeooO4JysQWpCyAUQ/78Bpxtzo1Ej/V
TrSVzHIXGQiHTTGFWYT4WKgCB0PJAso6YRpA3fmMBZavwKIWEL6IFRdb/BgP/3CY
S7yylXqm2vLYsJrt1YxP/MW+VPqyM9s1olvAAU6aYqfrWchytscKUqaVRbqOYHXB
RRVxQDDCGN+gt+WAeBoC8Rowi/SRJ6DwxMVp9jOAMIHIzxC3mxCX3imf87pLNCjI
vgJPPMAY6ubiwO738Pl/NnD1S3NQdRowsWtVeLdpP+uv9LWsmV9lTFI8ENv5qPNU
Gd/dgJlGI8r4YbxlCBtNUIsLZiRtcBWC5dXwwWzdcokpyor0AMBIeaKW+Q9GVGt7
Cw8g+1P/Yn4s7mWFTFmSuHQOnlx9mwb4Gnyo9bK5lE2airkcXHxgur70mQqyavnn
ug6wIh4kflxKiFQ4Z2cgMV9i9t0SBt+sDvq+H/1K4Ev7OLeK77uwUhnP1gxH/o40
yJcXfG9nzr9SaGyfB1sJt7MS4r7/lKGEVGt3CpA+vzKPjrLYZv2yKAn5zp4rJgEt
PNbbnUR+SaGhIQxUX7UCfwuQMv65HfmPSq6DibNotqZC762IHZP6IQUGB2U9HMgE
nOjyJzDwVufWWdzULvn92aG8mU1ef+wq6DNAsGkWtCG08SbS2NaJfI7eb/YecXhl
eqzagamQMQFyCs+zn2lnmQrFb7zP0UbOhRfWWiEAcJ32Bl1yguwC0odeHAHdnwmp
I8tZRX8RuQGbmfpj+Id3EpzYXf2SQEcy7J/1ltABD3/r6IWSfmHxNkztABFMuOa3
FxQ4anczLGSScOyf2S+StrrIwn3T3hyyVbHAjxtr953U/Eh+uBM35AN4mDDH2hcm
Bw2lVoyd3XbkM5ycVzmomfjnVOvAqlv3Tn1PJRtJg+MyHTLQI2drniKPiwmOOLn/
/Ns8O0ZbSFlUZqV07++MlPD0Aq8TxpZl7Skg3Aq6bE02JleL1appv9+a6LlAjAV7
x/Qa14RFNrBNQsNr2wvEXYfq2KN8ofv5rrsJaIWhkqUfjlV7YlHepXITljp0/odV
F6XmuBLKh+r32op0DQoyt2J5F05FNQfFh+NdRLQTbN42j4VJZO/+GYx9vtvL6np/
rcS+7sp81pB3md+WvrHrZGnG4+wrA7DktoTXd5knc7//k9d87Zvima9UmWExHpdX
MZpt8bmOiJrt2VcAmP5ekJlp+sdvvoEvnCLsyOt12o7iyBLGdVMXpLdQ3EARlfaf
w3FxKkkut+nIDuz/He13B33sFF4s2yvJvUTUE8de0CxVe+gz07WFJQYZorzaS+eY
db1IzVotTkfw/9LopEVXy430YEeyEY/oAlGX7RzFGTXmNArtkoat5628Tbp6RcS0
hCxCjsfLWhqxJxXoVijGzk6BD495bKez7s3vxBpD0sGmu/SlwiWKF2OK49WQNftA
zwIel6RSzNDkQ6S95G0ROKshNGP0QxODeOF4R9lqWVJAEciDvDVmYhZKs1AhhHVR
nmlRrhXtghmyLBJEcsOwr3i0O987TpGdQBttb2xdUFs+zUwi4xf36cMZM8kI54XL
vXmQ4CrLltT7ojaWCL+Z1Nv7i+SDz1L6rEW7qSEYGYIakLQU3cq7Z5pD1eQ76ELn
yHu7dqUmDNoIFboR7MsNxJ6QGR3h3x9689IvtGjOzmEQ9WPWD9lFQ3dX3qeQw3nM
MfWWPTG2+Z+NL7GBjTlmKmMzD1ZcrVlPhQgT+t3I8hgcyR751mAP24TEdkrZ2e7T
aDHA/Bkl2nEVZMT01KtNQfl4/dAyBlWbHu7QGU5atzschZGUHu+nHg0K9qJ948lh
z5XB1p0BGH5q87Vlsc7c+BBjBlwoG6viVXuTAYjJmHAmNRhbnN1pFJnmcTquf/wI
z2piqgRfhIg14ZKSC6NNKUp/JhzkpIM4ZQW47AMZrxTBwOtWiZlLlY5fxvygi0g6
zDe4Ljho3hxc4cBM4PyazfDFLlj62Y/C5eaOHijRgMfJtOc+sbeA7SX+86NkEbfa
gkh2AMf0st98CJY4K0mqW61tqeY7TquQ84hGacCEbVtSUjkVndttxLFOhFbrOoMt
OaUxSPtQnVtLITewS3i13W57t6FP/iUPjH9TmtxsBAIglOHKnyf++ToCAMrq36tk
bTqztpI5RzXJ4CbC0OcSzdM/UZn83dZd5xOxWqUPMNekfcykqH5xBU8uabg+mFeS
sE9CevbmLly4PWxB9L5aN//Nae1WUOcBLUrvZhi74f3RvSktzVJRY7mBE4mWLZ+C
f3LTpfhxyopvVq/HPCJFUyeJm0x86Nccs3H8kdFGOcPpwiBFTVXpENrHYp/oS117
dOlNdhhSomuIFyh40Nuf5UGu7s/OCOYzwnPTqwd38nPyPcYyl6WpW2TYFReHY+Qa
ULAI2ORY7FAPBAKFaNhgtu50IlmsgpsOgoFywfZ95cOp2UO8tZBxbbApprlf8gLu
NsdFkw9zIiD8pSLpEoTRBHIddI4SDovBinwcylBWSwHodIw2SY3jg2PYi4mM72mC
n/QpgS5bOZ5dK55+l4WXX1b+yfPWDLeIn8s7QdaIxIx6Ju6ow3K5/KojXhh4dV8+
hcBU2wShAFExLJzm/Or1qTwjfeibLilGdMLYpnlppHfDme5+V50U09tNKoqOA+2U
7+dbdHedZxxgOKsd1KIwe52L1Dmv0BSIQTFX/Qn7P85sm5GGTG43KTWcL8urD6o4
uLydBgR2tRWcceAxX1qTIYbR/athZrVMey8wQAyfSRpj5WAB5/PXYVdhfajvx3Zs
AFfVQsKhfos00EGESkF2d/xVKzT7lFqfpShvzbGqP2/MqxGTRDVcOJd/7aFQxxKf
/wpZlZ/kGV0GNzKcvakJ4NzUTy9sfwcTWXX3EwukJzalZmzDdKRIdZIZyyKKN3wZ
UTlEjjMvqONAI9f2fbsUafUSsUtI9Zel5+8YHxRuIabVGqVKd0bmUUBspYYMbpSx
xmK2Jap64R6itumlSWvSiZOG0Oe95XTLaEWliBsse3A+nR8FPNRiSw4tW946Bgdg
gWtwXPpEuxRHJAFBaqimOzIL4wb0VPsRlRgFCzqfz83IvTVMKPNkuMKbkWkS7nHg
DB6zRlAt0Tga2DJ2pnE34F4ulfWkFYyJZ1Jw35cu+VV9HsBQvu8ZbRe98AeEqez7
zeVPoeeUqggQPkN0kfqug/TnGubn6rr3MZKmy1EevPmSXzPXigclb9ZNkWPr7rKg
+40J8I3Fs0/g5iPXgKjU64Fc3kvgNOpLDE7EIuvfGB8fvjtMZ/H4G9O42xZqs/sI
tx1a8E4LT4UlazrWYVdZjyDtrey3to5u+tkf0/KV2K6mNsgSI5XEsLrTbWJUb7f7
fHLqtbJk7LVxwwCTNdLom+L63GKVtBh8BizeGatKKVryQUgd54nOiNZ4lcek2ZuM
Q43Nnf4iYjIL/7twz0mbt4Gnl+hk4Y2NuLoolLHfFJPaCsBH8DNBpjM3OcfJXFYe
B6QtMXPTAU5kzr887FtCcksz+b/WYrmJMGdAuf38FehAPDRumL99v5VQhra+pJaZ
pp6xEmDSFQjmhEe12lVbE6s6l8XMIp1XBXifbo5ZeGvJhvx2BkXSfnZzObSldsNm
Jx5eWOE8wyvreALGdDdkE7QanzkQ/QTCWw4nnh8Rbhde+XJxsSzLsAndZJIX4YSw
INZ810jHvLpbg057a8PW1Xm4UaN65NHwKO8sfFrEI75NuGosinfz0aNM80yRnjCG
VNcbRwjHH7o1PRaMCTyF/QAQdyf40QjyZDvojRrBdp06IPExtB4WG6zhHZgKtrUr
Jd+cVg/X477gAeSa7eOsD/BjJQ/l1W2fyQlm8/vGHrQHzFG9H1kxsQunc7TD4qBx
M/Loy0+OcEzlNsHxJa/7UGaF+uGxidLBZxSVu2XDtOiHRXLb2yat9AoEKH504DTF
xehHawquFAOhHJqkP5nTnnNmAQMsMq304wterk3cVxm50Fd0DXTAQhdHiriLf+Xw
+SMfSg1J1CR+6+Ly7lgg0dEk4fb5+enBloKmmll1W7bxav0mRyUvDmyHL+C/zc4k
Kl5Iz2A+xv/sNJqy1kAqIw0ydTOZZ9jW0iycmwFfGphke2jnqdiLREqSwFlrFcNM
LmObnh4u2H8u2JQvmFBhDdzBGPKMTRwUGDElneNEXsdaoWErvuSo794xqy37gyyg
hok0t3NC2ndh3d/O/e8bh2uRNHmZLoxb5IksI5XMSWjNNiR7CDqDnXR22L+pywL5
/Dy5auSqI+RoEo7MEGhZY35sQphOG44Tg0oRCsc7fP6DKClRy3PNmWQ5Omd6P4Ay
LdCJICFM9YEE9md4cYxKtN72HR4iFEH63tieKCiVmrRZ8hl6x6QYPWobH+51YvcN
2LIlTpC++IDazQeLKLuO1sILy/YN6u/IHjunQ3Cv0lz09s8uHuLiCFW0qTseITUJ
cwG+yKjZQ0ORnmnahhKruW3a6JYHBFyA9oofeP/0L0AZ8FrMinENX49xKimid3qJ
NVo3nSMTSYJY/0OVoBlif63V7WL3ziVte9vFBuGJnA1g4RSiCn6sXIa2WtzPdzSL
1Pae6ustsbh5E8icc88cUMcl3XdKm5ZEWtYzH/mhqcwbKDdZ8B5OekPPZ3Sm03Tt
f9tqXluTgywrvIQDdGDqt660Y5lpumrOYC4TJBvaljVsnIh/Dqqgs4+Hjdbn3IwI
pEFNpji8f+l/l5S2wWyVVBRvTKMm/B/s63JDYqK0jjhcc92df3qI+H8Sf/Pe0i7Y
ohW74PMZNnyOxm9u1QK2FC/dRyrbZ9gu9WynZBnoJtNYzW1iYrMpizbYRGqKz2/S
vrfOGZ8uohBDmXHm7F1A4eqJ6id048NgBmDsbK/gI7TVHh3KoUgvbL9PwY7ak6mM
TNNBmTlCCRFaT2A/7+UhlbRi7Wath1IPkS+hxdFIGAjPT1JeRFrUPLFyyN/LE+bj
5BK/5WKE+ndwl7m8Jq7xk9Yrn8vb9bCqXMkAXoGPbMeD6rSft8lEF3fhZAw+DQAq
6ZBVuQfUcVDLzaeOU9g/7x7+K/0iKDusWxWpk7Y5S0FihlKtr73RiV4fewq6APPf
pQpXIeIU4+nS5hYOjLB7HZSbB7udLHh/avnPJ1ltVcMxYzMu9vtxTojvjOPFuQPN
bLHxmDrpmhL012EY2PPRCbasRVE27zKvFj6YbXLaLF+iQ2u9VsJScOoxwLifIukP
Q+T1inVhpStaKj/uCJ7tcfC0QFmayfABLSfJZPfnqXwuBtd4fDVSAPzQgFJ7ry4H
WUNerW/V6Y85dx0Wwz+VUZ2GrAPtHXZvdri3wongLl39saK4aHRlEC7u7rWGwhjm
iJlvRXw936+juVjw3bi8dlRBGj8aWh1k9dYVjclM/0JAm0DDV/fLC+UYtii7mdWC
obG713oKFmsbLTrxUAafrhhohiuyIaiu7pzr8nhDXRqMxJXD8DVlE1tzA4syGSI2
vUAZX3bE1mfciHDji2YaUtO9EYNwCdeZdmsssro8GIuR7Z4X9kFriNgpoygR5eVa
vot7rxxzvQIfTDaJdBxR/Atg0TTi4n1dNC8qOIvV1JflXiZNTCdSu5BqwnKJT6IJ
aZbMFaAa7OPrHuFi74dMO2XniqbZHO+1YRPjF4fx1RqueWyQL0OrFEAVIfA0nHre
Wf7yNBoP0TWTEv8hCvojz313aXBVBCwiy+Hek4hDkFwhe0PcPAWzJSmpgFHZQenU
xAJH9zVutJAkooSzIoqThDwGsoyQdww03xbE+Xhj7y3JaryzkksPiulCMB+SNgQA
TK5XJgg1CyMtzwTR6nCoL0s0eLcZU2rG2L7anS1qDtFZJy1ZOtWkrJQl0wDYWr3t
bQiVYWwzxb8gQ7LuqztBpLGVg8+AZtzXIx8NAoAqr4DKywnff6CXBlLj/KHA6SeP
a8mR5Kg6KjbKpRc0Cco+XIc/N08D9oX07l8XBNpl371o/hyKr+QL6nA6eX6+kAvJ
459Elz+x4Db3zjXb4qEU18dMo8okr7WxLwMZ0r9AV/6mQ2eMIOfNq+ZS4oqVklaT
f5wX6tkDq82IWBkSC4e9lRf27B54wGEv7BhQQd3raeqCRMslZYGCT5aQpTHtwOm6
x4ulSGL1BI59yxihe9h+3SajHhxxPH3gPx1fwu425xKMJj7mpbOqkzjZMmHzOGyb
kLb6ip2hAGLpdtZ0L08zqrez3VYTG9qngIKGCxbTXqyqf0mqNTAejb2FGLYpZTg1
7Er9CkLEsXbcvnkWSCj4WzEKtwecP7vr5JuPyA5oLw5nz+0QT2THpiqqg+mNDCeo
sRMTumMb0N15bseqgic3e/2X+U1cUgg3TY4i4zV/4JJeTDZkfn/LtXL6uxvxW2G+
gqFcvOGWc88L6JgzZucxFYh082GxKmHT5CdubyUW6BTxu4zM5neAD185w3Sh6yut
zy0aL3Q6KZj6u3U/oYVoq8i7h9CsEf7gwnfRIbG/Vgv3FvPSg3j6sEmmd43d+bWO
R59uGf4nD/ciAGnuqbzVygO9VxnVhpgO8Snsgh5/vkvR80XHlYMlK4lEok7Oi7vx
4OfAVyJgHCxFd7BF+1dBenYwYEcK4WHCHLrzvFbTdZsNle5dR3RvUGRme5vFsYoE
m65yke7xSgLxlFVdlmDF07zbpp58UpX6Nn+j5xznPfQEmzF/Oi3RXiTGK+yvXgxS
eIutHPa3kYpggk8I7idVaTunIjfS7SwVDlGQvp2Lg3YSGqEC6Mg7VYQdC12XGPvT
39IG+LMnRs82WQ/x2sS1XAQ0u0rzJRuQ4jICz0rnVGSagDN6FcvBI80NiS9I3cll
SunsvrEQ628bD2aBuoJf8gnjFW7MJmmh8QnCZTHL2lHo9SJcYmIzLTEgQ14KJB8D
WcKUmgfpix95ipZUbIUB82j2Hfd+nnJlUTYbSDA0T9FWKYfqfLfwxywWdGyI5LO7
/Z5hu55C/dVPK/5M3cyo/uwQlb8sE2S0dKJa4p4PPrEDabNrgiBI3cM1rvM05yrM
XU3WdvUY47WoA0ti9z7jhFbDJGfYvOfSUB785+155sruwmFTmaS0ORM8UWE5CW1s
BegpSTZFBW9Lbqy3LFRKvNB0+aAve1d+1LoRmuWcjwJbovzSNE793cUuog511wIm
oD6WCrIeEXw1QV0smtCaU0x6YVhw6E/DXCRlTkrMQPQgTTgHAl1FJjHMHpTpMa9K
LtShBMpWT762/6nwAwTXGXmJ08EQ+gJDu4ZbHdyoosfnZaB6hKh/ykJXATlZOHOI
mgSQCcoLKw+TPIxZcpw3PBgFNRXLcg4SVPpajV0w/hS1GsG1AoJuB/3qK/ZCRg+S
ThOxqF7q6nEmKmXAVrqGJpniiSOr/xqlpx009DQGLFlQW9dnkWac9EoMKPbhp0Hy
QNWCH4BVf0z9gjrAYZ+e10g5v1LPEEEzJM4+h+vV2xEZztQmEFmcpilXKVWHPjVV
lQWVLxmnFAaAkwgbT32yCdmU/DhLRuB/e0J9T3WzihBxa9aew0EWb1FfwsOX3QvL
oxRMzMzlfJYFd7ybNB5d9q3Akru6455lerPUZi8MBmI1QLn3JcoVVgK+bOIDP17J
jGWRrWxaTyEFe15bN2DopdIsC08HyT6H8YrUjap89zcn12ai2zLUAqVv38NO3tbw
afH3gm1pZNfEq4O3iOL/H7FglnqjJNAfyPekcpKaxNnHSpvDWHK1DQdzcAwRKCOT
yWw4C+MoFRzNlujGGYt9TAsmBpu9ud4wMlAGKyCCn+CYRAh5dlcy2Z4msMUyd+EW
Fx6PicryciKb4+cpV9AixJtw6ykDt+FJb/hdrdwmFdkOhtNbryou+VHfYDoOFpm/
qzqrsrDe6OF75OaFlhI9tHNSSuCdqjpLx0aPcQW1mgqjwMuSmgvTTQbO3s7HxyOZ
KgeJI3zTHWnArdFnukJDj+ch2dj+BhZPWQNThQL0ltMPWeQ2QI456xWsfs7eXzRz
3mTkllubc4jXNYmmN5uUGfLamAVT/Vg4nnX4HKyDXDHi5tKz/S0vf5q0mIiez/XV
mJHwr6DpIXx7BFZIrvv/LVbVvZ8ARqC3SI9JVTyGJWNgmmxRlV6kvKC2O2Ear32p
kgt0UTaQjbEyzb+PqqEgKfeffTjiwju7oHRGLJT70LAeG5xf0YeGBK1HfhUvpuha
DthuglVYjlXi/Bs1CjBfJVZ+VnfG00btgzfxPefh/F1OXL22ldcVCzIpWZShmoNe
oUTw+KjRrtv9WB5D7q+/3vj5myor651awOplJGF4ksy+K2JxdFoNV9J2RFJrkpqe
Zhh09zGPZujiYjKfhupAcDCqOYpIehir0liGKQl5ZvqYlyoPn3iWIEz0odSjFqUh
fP23AXX8eJ4n0whYX+om5VUr/t4VHfGvOq/bWwCzr1en/CmR/Z7EhxoAfrl0LJzc
XF22ZaW6dolktLv4TufcdmwWJRxrle6zlAQqYUEN/SFOmCCWUilUYmzCFZTkzuR/
Yjp3L55GB4+CILoo78lCgQHFEH1n8CqQznn6lPpGnLev1WMyIe1DEQdQM2JHe80v
SnMSueH4n+xMwK0jBGq2YwFCoXr9458u7eYwdkXU8wN9Ja0WzpVZHWYuD43Pttl5
Cyz6Uro52jEkgc1L2KTSrycVbbOJz5iBbiE1WgGGQkfu5moOA98nLoKRvICQgtCZ
Sa/H0p/Ycuh2hTVhlLt0aFPMdHYzKmIL1yivZ5nvl89xjahUPeQGN83PHyUP9LsT
4sL4IKKS/DSEOJakguAOnVpbyyb8SptYzo425U0nwTfSScCCrvBUuN78/1F57u1d
ca0+ky0JQNJs7ADVdqY8fT0I1Gf4mHgPsXcXGPUYSQ0ZLwrU8BC+6C6jst409HxD
Y0oRvhCn7PXwekhGA30nz7zjneGvQAsdGJ4k0b0LohRv8CBk5zu/DoopxCpoQovo
7S4QUN+C/xxAu4otATZhyUgVAeLeJvmvHU1zOM/6Ndjiy3t2rWYjKRL2GupF6u5E
SCbnFHPjF2gRqYtouas2k6tB1MHp1Qp4dVJ1SvyC8fQD6WvLpLv2/+K2FykyrhGD
G5HzKzZr03EhY2QEwmMq1JmA6T1GRawvF99S80N60RAKh3AAg0drRmYFvyyVPhf3
J5Ygt/CLR2W4WA3cKvWTnxzhzrg7f3kUHb44P52k2Rf6Ki1aUgtMaRj8a8E3cg5+
Tu8gJaNnfcfGrojZX767E1sKPmEr7NiYp2ZeZM+7nwVY7EJCEYSEc1bkmfDT9s+8
13TN1daMTZ2RGV/jIL0NKU6PQtvceipwz1f/Gb6YhVjIlgQJSACD/NIsy3v/03TB
hZL6LwllYcmebvOzmy7bE0Gu6SHSl66AWTI8RKMs+GpfXyq9hYalxo0sHg7oGH7I
uZRlhLvxJsyClTTS3h1KakpTM15jt7a0HwG64Ql2bGNDKyWXWq2x9DnvOYb6XlEI
nKgP7L5TqsbUx3rT7U0++UZy5uaYx6/OK62oXD7KqOFE07oLykGDpt59Aqawo9Cc
7AX8468wZpsTTUbESU9SalGYZCGk6BHlbaddA8smzP4VmcAchg/3rJFlCXZgvrxj
Yis0C1TSgiiUJHkjJIAkUMuiJ48USOxJb6pXC6d9KAkdhaCaheh8HeMYo2DZsJ2s
ICqZPlXmqwhXerc7w2coF6eIaE5YjQIZDg51+CUAh5VH+/2kfdtXnvj5tgHHPChT
24Sf5hq8A2pqCIYUmOKyrQbcGEjs83i8oQGM9702RhSquBTAcUoxMwfKaEg5HG8a
TEr6cdttJWKSbOMzpwPEFz4t2arbmSGHHyG6nBlGFKCmu0e2VVRq3JPvzg96bjKR
C10N6SaFVDmHR0PgRoXhiC0+pvhzzdk/JnjxGMdPVLMFQ3ILHVDG8B896o6PZqJA
UbhatpxktIT0trBsWILXKQy2DgSUhsFssXXxCMATDgqi7vTf2VwgXaAsR+BUc00e
P8MCIpd6l8a6nj7WnCdEkljXwMNP1RxX6EsfPghgkW8Vd859t8mxoQu7EsOovlId
LRx968CgC6YNsgU2fjrwJ5S6cvXrONZ4x7Qto6EA6wOheV8SRBDMfAC4V8ekTE3Q
tFN2Dq6bc4j8AMOXfqNGRodlATta056LDbXSLIKVWNQKNC6dG4wOBVh5J1FI3o8N
95Lo1ulucyDaQvVEkp6XzrUp186dyRPEgcEvU6Vx8uEechioxlThtCqpNA97M0nx
8JVsBCZsuD3mMSZ8cVJ4qYkVSR0zsy7EY0BvvB+SlBc4XEcsyd8Vph8A3gN5PWpc
RdxixOEYObxFN0h1OJc6iOQ34WMJwrpxuk/N211H7lAOFqh0ODExIAusYBJMIego
/oK/prHMP22kFiAlpABG2WMH2SSX32fnIoK+2B11sFlcLoXbkHa8h0ZiSjhzVFe5
99xahkY0KgFGs5avaBYM0CV7OVCvDw9Dve2MEww4Rbk9Qlx03NW7ifvBrCh2pom+
wGRX2QU6nOHAl9AN8a7N5AualciedMB/EIv/HbFhxUgRMmRlwPrGh9KNrAmr2o8f
GHKZQ/84UXgwXUhiuoQ6dxaSGDk9o5Ir2xVGnhLm24Oq0gNpp9mhBiAyT3By3I2z
MUV06BE5Cq9D+I8wTvLsY5dt8Sd95cf91wTs536b3/q7+NVGhO50I+xDvaTZrRDC
8zwvc/lEhTYLXbZNrCA81Y7F6JVdpd70nofzql0fYIa/B4jAZmMB14PkT94Tf27m
FLJUqOt+5UCmPAD+GRKycxZ8qPfwUxBCw8odIUrraYF6/UdB/UaKYty2ylv1l2bB
tEOklzK0V3TuSNosmGS+EauAs4z0UU9mAZmQ0gWScpTXFXWNtKa/X8VkRXt8rgGK
iPzWsjyRJ/BQKUnFFSKq3FkWP2wmxSoeT/DuDvAkkKRIxeKkatet9VMZPsRaCMKL
ZFH2lS3N9RnWmhHtpVvEX4oX7Bgc+16ZNDVy5IXXwmezBtu7hgkBt5hbgXLtxZSs
lQL3Prk3TgOmjWskWfrHvU2cRRdZ0HM3Azg7DUuAFaeW0VuNzKpZ9hbYWSOVCC0G
9EH0Vsxgi1e3RZamPa2G4q8+ZNnJGJm1Zoeueumd6gTmAq7cQh/P8cssuKpPGQK9
YsxBV/NS18Xp9FFkycM1X6v9X9XovT8pF/f/rsVZjWpIICIgxkzibIslE8qAjhMX
+3mpTmaUuWcY8AAKsMy/lgB+EuwAA1wAFgt9X7bmQ4vGjzIiwO1yL4pP0UDixLy1
GdyIF19qhwtWHQ2JXf2gB2wjKtXe7q0YvUWNeBV5jpzkF2r8sCx/sAqbQEJSe0bl
7bqTzDcPVkkWefJjuJ9pcxpZZNkC4iNwWzrWmiKh3MJZuv4GAVQAlISUMGZvOxlT
2hGbM+Hjk+D9bjQ6k3Tznm3lgQe8QM9JlCLSHI36S86FklfHI5GtHMfK5UI0GPk1
1qT0eBiLu/gS9/acDxEpeBnzgZO+iJ/9inTh6oVFyyAyFh+yU9QwgP+LopKStrGy
GlihnWnU/FqrYz/jKM63/gcsxpOvr4hsojo4PAGCoWf2wC6CcLH843uJour4NdEU
utEKQ6jCoUQGDDyYG8GaEKhf6Tlj375ad51Ek2C4sALFz5nMYRgPUlpKqCF+uyIR
c9SMPPwrySOjuXxTSjGtgsVHlyjZe2Ib9EbExauCC18TaqeNV/cluMKr0CJWUftJ
CUn5jzTMxwYBkhn9ZBenOIp5fN0Nbt4EL25X5QYPGIS+b6pNBCRyi/JRqXwYOBXG
dBT8XYc3Ng7Mrnlg0YGQ/uTet5gsO/w15nYLJiAkx15q6b+t+iOVU9jvlZAJss0+
CQ2EFqY7beS8TzJjBO1ENRQWzUF2C53dw7p/rpJp6xWE66HbbY+xD3eCeFA/4Id1
Vb+AUU4xxRPJi+pRL3KJQ6l1mLY0G1E98T3eRHyq7C1bOJBvdrVyY9CXz4k+BWni
YULxwm37WWoIYzFtWAusJQFjbrJs2M8uJuxyxOvnbhui4sZJi0Qz1w4Dy2n5CrpY
nRMvzuJWHYxNSgBDtGa56z0T90egPYdVlZgLdar9IR3PcihzjCh1aXrPe2EpQYhT
cmPIuMiGllYUfaSXMNr5b5MXZO2Y0d8Y3fQRYQIIFD2hP1tSoBTWFpXarTgRSwQI
zBUVLPLMvWv1qIdndRj2lu46Rwlx1fUcAPc9WNfvOe9vBlEPKzCis29zYHBfDTpS
wvBIi5TuHEgsfo1OUuU7GcQ+RQJV6zxc0Ogj3Itvp6fUj4HqYUQwEYdn7tGVcKRW
M8YiDEAs5IjENGQqrXO4eWgwadZ9oDNwe9FzJM5XilqzgX8Gr5KMMEoxOKB28CX6
cKCOA4Y9v8Wn7a+z/gcsPIILknMlxGKcAxe44rYCBhAoYkBL9NfJw/wawMggUNnD
lDPSU/99ocrZsmOq3LFR/D4qwfQuG4C8Ud3ryx067ONX4rgSeIkjrmVcA6eeks2c
wF1QO8+mPofn49F1UjmoTvmsYjwIdB9HS+80FOb+ROqTXSXQDz0+JyDzfNvFYu7u
RzctdTw0aqfNtx5WjrpKvbasjgjNff8tXVjRaZ9IiI1sLSpZgQbTr8ZlWut59Ue+
NMMNDUid7NxuynsqeSg1K/FQIXbWNJpJVbOxIBPgn4Rlm2f6tGP+xrKWIXG6PFK/
cOQKN/4iq9ZILatNBYmcYSKybBQQbo0Xzn5lHu8Uq98HHcz2DK2fx57AN6vr+RUu
J+HwVgTc9yjC0qkFNzOnB9XPeluCETIyi2b6AxuVSMm36K78RilSEOxxzZwYVJBd
cdspT0AznfoSG7FdO3BbTCpITkFHXRMyEOlT3NqMEMvE3N5PqNrNDI73B4BEO7gn
ZsjOxNLZ0suLVsBRMxwydbijkO4jvzfYc/Q3khLCOfJOA9bvcbZjld8c1jt/omOA
TNueMZ5R3QzqxFtVr5VkxT5GmRP8qZN2jFeBXaoydHMk53Y/6j53FT4G6JN3ZhlW
GpogPw5Nxe2Oj7b21YGLQpZHKX1W0zjpRKQ7m9YrDiMISRygmILqLSliByEzFuQ9
x5f/rCnFguXvD0Z4BrkHZ3fJ9V7NlCPCXdBepZ3sQA46cxBQIqXKNVQDdzAn5E/c
M4EjQPStOFknD0AqlLMXZNtcRBnUZe6e8e9On2ioE69cJNVtDF1Mf+4imGKZuGAz
wvdl438fepWBpJAJhAtPSuZJIEixp3UlSn6JfkvFiK1sWRgkLBkl9j8DNx2TVxke
0D79o623lybsu4w9Pd7tQ0opliePE6vi5a8g/YtpRfnnKewVc0DCKfj5H1NZkT0K
ky+7ytE5C98Xm1J9jPNTBR3HQB6p2BN0skhogc4pdChWpIFZ2dsaEjpHdAaUPjch
md+fD4whVuRHb/XifVtyTChMin3Uaf1Cpn8exP3NlDXSq5Pv+bvdA586WFsdNiqo
2Mys2nyN805lOvYOktWhn8Dbn4jFdPmF58dqnzOYq7Xf/G3LeEUNPWwoGDHYY9e3
HyvGIaUOMztK9Fj/KxRFBvfqI91B/PD8hnPqIsNNZ7GkvLpyFNvELYJd0ZCftR4q
uggoMTVkg1Nhtvxf6QuePN+hI/I1rJzmSluB+2LJPEUcEzYxQvJ/H3wjYXs0OyIP
5yhEL+Jm/SFf8yvFB3lVFSYSe0s9HOXrdIKa4hOoSq+GuezG2fukq0HqhEJ+s8w4
/TFVOI1LScM0XQBLleCx0jnFPEnlF/twUm0ChzI3Lx3BtsOc3NVqZtD9OE+4via9
sKR69hj9uopO+eoGRvxQX6J130AFXOuLTWHpRzCLx6OOeUkH2YiW0lTaaY2KVora
iGFiwyGcxhNuTfYTnktVOPqibDssApz7X9l5rQgmVLNOS8gqsO9ZCmajhGNel5Bk
9OhYlINjmTXC4DOiA6/ijBgAZ3Pnmn6Gh1oV0uWuqg6pwjQS4o2pD7cMbz5yS6yu
oflDiBlkfwuJ3oxnHrvlXiVFQAHqGAbfIqLgUmXmRmVyyPebPdc2pfxahHkH9CGV
1I1ik63eCbmoM1yKEqMIlX793nvN5tpbsFX+cHiGRsp4cIZsw26ZXnWSewmdO/gi
aTvmMqZwU5hBBTsm1BIwvRp+1bHMBM31MxgLKbp8xX6HXBOIjSWwLGir0+VFWsds
ewbxanqNMiYxaXLpg3zmVVzThyP7kJpJrZ0KPc2YfVwlsoofdstPO3O6FDN3hVB2
P5F9tPLpQFf/XUMQtVIU0BpmQ8rsZ2Y8k1vwIFutn09YtQ12g9oOF1nD86FgMatC
rJ2ITqOfKqbHH+eNlq5RQfX5oIXqdFbeUisGDsMVEIgXvQS3Srl5ppzSJd00W0CO
GhWDLcoNrkI2cRTHF0/RQXDqoOHH6Foaj6CtLrYZn57Ha/xPYp8SxLkY3qdSWXxb
qh4kg4gF4xZDzrjVR30E5ZRrw6w3TvKkEBbxVUBix2LP61P0WJNqftmHqWGawBBa
2X7o9WXogJhumJs6VLMgy5UsfltqJH0EuA6cc8KWWugjg2dt01KrBUQGWXH8upY6
a/Y996QSkv0Aq8CZ2EDGPlDK5XK5YQ4Vdsr6DV+NjlJFfsX7Cn3pYpEYz/pzQotf
lbcEJKTO7dkpDVeZqoXPUL4eZDF84GKYF2UNz7GaGj+bDozISuIKY69ME4HXQGiD
A9M3/7/tQuAnoKdPFtLcrxbnivESJFYN/GqjgFBkX8MZGAPUusmqY0cYZcjGp32N
u9FN0uqguhwXZoL92u+HhYZzTY+F9anUALn4tTOwkkLjsE3UzJ+pAw9ZRw1ti65h
TeGJpYsTqxKxU6HlgWcokbKcc5uwb4mZDPBHxdppLUDfLhnk5UxOb+WkL0ZCw1Pc
bO1Sq5q08RaPHoMTCKGdjPwATvFYoUGDpzSNL6sDrFqZ4uv6G/qoyWomjc1SV4e2
5XrAvKc5qJX4iXiW85y0JOA/FTeEzKoSwDxQGvFouw5QHBa9yLr1MeG1vVvsdA28
0+V+i48acZASM+cURDN1EK20ttMo/pccPZpX5p4ZIQ2Gk/1kwFQE7AmtpK5VEWdH
Tqa4gQRkj6T169PImI5jREZyEDTr+q+wcwVtQMoFqikExX+hWl1sFitbR3fMIr5G
YJace5mEAXueKhgs2CetLMrQKLp7PYxOMkTpsAMYogKMF5gj0rSVj6gpNcfpxf9H
YtNDc2LVR2PPGekyW9N9cCCi1YckTOogmAELsQ5s3Eh5NV9aSo4W6uhm9ASGEX5F
aYYA3VJBYiF2xD0YLyqj8kj+Yd1GwF5FmUOrKv7diYPwxOzdgUVTvlnLzrdKA8bw
awqYWBWXpaLx10j4AHYfQpT7k8aO3feEj/nu/yALDfIG5ip3AAvWWurjetv5assW
odpCgCwrkAc4e4IhqvwCXyaNIzx7q6cVjeAUrKZOvrF6Yfuox7lw6EM4fhzlu7yU
NnOUv+srZNczB1W08xdgBPGJMsWVNtqb98DUXOH0yifT4EpH4mWMYXCFCT3LfMYm
VZelkN3aeI/roFWVV6bXMROOZmuF2SUSIh+jD1qIRabtAWbLFNMT8LQDt/kKAdiA
7QNPfZLDguZ8hyOKQy868/eGlf408U4qrf3p0sPxe8JO8vr0YPY/VsMYRiV/teVx
IdOXeOwcb0T6c4elqNJpfQYfccOtlW2PzqgvIoxv4djaunggVEcAqDLqZJuDE6RG
l585H5oymp28OuDfLSTtK3WRc640QZUEPK4O08hkgQomPriDUvCuMFMCyFBbpZ5l
RReTibiFXdWp/XjCBldayrPFZIBm9B30/2oohj284/DEp3k4BmG3xCpCQSBxXq51
kM5jk8ZGsgHuIp3dKjD5IZJkT0L4scf0WrFDmvT+o1Kfbw5Z4BQYALxjW3bNoY23
kVp3NFr+OrqQduUgMOF5cZaUkH0+BAO7yG9OWuE4WT+LxISCYgj15+sJkIX/tKug
ZmpGMnlnaqTZj00Ba1sisZSSter0XVKjszp1Vm5x+Fkok1OcX6FkwD8AOsiwYRi8
IcuGF6j8oxXHA4Of6LBXWBfaR19dEqKHeho3+nObHgaG6tyabozKGIINfmsldREF
2MGet+AmApicC3+PSfjHFN9lHwR7ocAHzP2vJba20KifI0U4ZJHgOnm+6e+rWqPQ
4lB/0/R67rekeJZx9rcFcFNgGSC9h2U6OFqBf6ckkTepdHMfFafC7Cr8mYPk4Pru
p+GUTIfdIMviQAZiCka6X76DVY0Pm+c54GkUgfSgCWN18UxuTVxwVzut9O3etRl6
dr02Jnh0Lf7Yr5YD2dqOCTN2X5V3lvkx8QXNicMxLWIK8Xhnz7NKML736tC5jcoW
VxcxPz6fV135XRZt1wbUyCboEvDz8bHs6UFhITZNXdjRg/ejxaPpeugxG8SWHnSP
AxodvwleAk0sHTiviuh+PEiYn2lVyPAYwsqwr307YTTT45rzy0rUtjy+MiqAaob7
YNI+REOfT/IFDguV+UInxGB+wWKTarTCIcPWUeEWcjDo47PEvrvIg5Lt9AspEIH/
e1ndfjZ8NG5kevj3jLxGsUoicLcHfdWmtDpkquzszGApxGHXvAq9eBwPK842C9RY
/zcOMrLU6bRAQ2wmEmfXM6UwjaVZ/sHHI4JjVu/mZdC7oWEC9nF0NvCSgT65mgvs
xOataUHvy/rUDEH4niXphP1DmmqHU70C+LluVk44KnND4hXax7Fr2o0+8e8kItDp
gV14zuzLw/JMl/3XxdJzrLCXg77dvcEGhhGOTP8ygztgB/5oWO9Fja5RHMMelNY8
VRA7RaiaSAB73m6l6npPmM6+T8qRGyse/Cm2jqDGjL0WTQkOApRNO9mgW77jSRn/
hxyvb0afls0S1MdOyfmE1IrP7zYFE6nlxuO3P+535OX5WSHdHumq+r7J1XdRZyHO
sDTyC2jMyLelnpZ2Q6G10kaPLx1jDB9jFavTAyHo+P7UnNqjk6F/jb+ERNZcE6gi
wM1cGKjz0I+8Ny5w4lKzvueGAMvXHjBTkW5S9ov2dWXS/nAFUQOxZnh9D1vuisVz
717E11RnFz5B3i9PyzntYWBnujVaNn6dCm8ZO+mVIlBFXjfCO3eVuj9SCuzUJ90k
65DtYDUeH6f9541Nj2w2gEhQQ5DjSQciGA9hJR/2q3TEE+331M5DMrKsVyeePY2c
QmUo4go8li9/H2NTLEntmjSquk4qHmPWk6yC3Ujkvy2u0qEZkSjhjDZ2ZDDHYe0A
SEzuepY57sIqGQWL5WYZXXjeWvRil8QnTOufT+vGZS3FcZRCEGKUMOkq6m9NS1XG
MwikVpqfHWX4BWh0RTZGkBp4ByRDZk5Ku8DnM5s+9bgK76wo1hmtM0JmYeUIH/cO
kNvlYB7fBD9mLqBQT9yvFCbVQwkyG0EUiuqNygdKNyUdV3efGnGt+jmUm4I1E9Od
PBbkWKjKxsjouiZHE0XPpNF0HegoUNGnZbUL4NprfSzqVvYh1qVZKKsSXC9dMy9U
q39aYz3hTkiCrZ+/+kzMeKBm0nUMtEXTH88A3Pqf/9544DWo+56c/Hzy5Oef5y7I
K52kx0w4xU7Z+kgdsklDcdwCTXd1k+GnpjEMcbddsQMz5Cw+eQLyMflnoOsQEvHt
pshcZXrEhfgBpDUORt9elRDSpVpf1odRhwSYARHQyfSl/mU4Lw9A4yrEDeSBXIls
ycA/a+LwuuWcjl3u2j2LiBTiCCcvLV+muh+63z/yJZMAiHPthrljQ0wFg4EF24bT
aRsnCCoXHwU25PDfVS4Ay890Sue+PP3sp6Lbk7JfVuJunwK6dyzgQILuIZa3h4oA
2N12jNDSX0s4HUbkXwIYbfN0VLBrwiFC3K1oLW6y6oivSnOvCKJ+tnP3hOPZF1nt
GkUfoWXiO5lpi9FJpb2BaHdjmu63+3UWz6281orDCNHBtOiSuI10lJu36+U+xvQd
QJoDjSEnLsgaUI09dtmTLzCKi93zWZloWAzvPkk3PQ//duRnaelaHKwTg46K0JMO
B16YGiN86IndJ4W+OlAcE+WEwFVeeIIVEf2aO6DAAjNaYzPhzth0GhVMFJeKO3lu
2pMyPs/UmSSD3vjKbYyWP8xj2WfyFl8aRecwX6BrsB05icB/XWbvxhEcOoq/qmlI
c1SFzBHTz61VUuPFpf7aGY9d3PNUe4DlTK4YoydS6m0GvdXKyIPKHPnq4cewCOB4
/WLdMsbezi0vrj67S5kRralLNkGEMXQOghq/4wMDPI1DmCKHU0a2Pc616zsML6/1
S7yxr/h/bct0spz7sqrgTpEaiqxZWpRZCgJQ++sLmZ7U801E2/BFrAlocDppkvlf
uVU+EmaMoN54RAx5qIJv1Uxk09xgk/i8IhEn2zdJOblLl1cqJUHS/4YFoPE/QKSy
QwslMNe0FFDb9shF7jcefPykmfdgyEbD5tWR4LLppdI45o0W4fU7RecNq1ai5M4k
MbcV2tgQyaEDI6yjr9lqAZZDzxaCOxOZCG3M7zq2be63sPSIUYmM/u7vy0HVJxnU
q/o0DNzqitkhrn3NUVcoTw/8pf8vvk9cO42M2ayIY+4lhJ4Sp1iaGc68WWGTMZG3
VO2LCySAHc6xZkDVf9sCOsAgdu5uT4awQ0ZE0EAz9zrKBbG6xlFX102HyINSG7bW
Yab7jSv9IrNHW2HMwg7rqGhcutMb5FbyIh75mMDe8LSZAVkvyM8rHC5xQqzCGMCD
uukm+Qes66cYCUKFdRv36oTbTuNKQWjmB+Ty7Ee8tZ2hnibr8PfN0GrUG/E/hCcr
Zn10d0VG0dIGuCnwj4fyhDD2SP2IEliPpOZxqrhQD/2zyqjmdyoJSaekEfGxzC5o
JW2gIcWzZh/s+Q5sXQZ9J61o+mjuTUHL7nlKqb5bS7ZRM968Op+sOlWI7i5/SPGe
G08BjabUtCoqDB67YuHRCS48yJ3M1nbDqeuzYrSRRcMysvG8Hp4ugCsN96taSgXy
/ArqW/vQ99/PLRLjTvPg5t+Cu2ZzG0OKGF/V/Xb/BEAhSgBGNUNgk5ldn78wsrxj
7wZDLS9yRNQF8RnnBg61/mYZWbcO3z7JBlaBrAg52a44npqE7LsItzCQgax8ADDd
DHskX6SjBBK3L8vnYhhntn7Uj9MtIsXyAk54IbKiM5D09Q3+S9mQSsqNSVL7mJU/
NYfAe1OUxVIu4CIBmN2uCIJC7OKHABUFmeOEsH6vwLtTS5GCVtawbqB/vc3pCZlo
NmlI6Az6TYt7SudOKoDijlneqPkwElB1GRyl15k/8rIsMKMVheKN3f0ZbHkiAn6u
7em8/OVlUjzYe2gVDn0xzVBd7OQA6UauGp+G9bFss2yNRQial8+swuPaZvGH/l/U
q4reRyxfcoLlu7alZYnZbA==

`pragma protect end_protected
