// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KA9/f4AvnN+nVGeqWVDoe4I9VSOtIrpXdnuxVAGIIXjtr8BkFtpScErC+CTg
oQdjJPhPOliIul4ACHr848nr/nYbJXh1/AjlRfSFjzyKSmxqL5U6OhK32gUs
F7GhSGFRXTwvLR1gcq9RjHsKUUQ4QiaDlOVontD+FRO/QvaxdgHeHXsxaYBN
Uo5Bay8lTScEPzyX6ugnwVY2KVKfbFMBPmWtf8/ojZl9A3LjYe1UvGnGCklQ
3nMhjiCGPz2kA6m/TfX0S67zqp/6M66eCyuMQ7UzJo6NchPV098Eg9oNyY0o
b5h8uRssanjNxTNy/M7A+E2rjJIOPBPWrJYpmq2tIg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aI/AseYk6OYB9Rpu+/axDtryHbpQJpUvWZCK0JnVGuplVFYOBNgEE6awhmbF
cFoon8GsMKb2x07601Ysz5vDkqBEw7OvHwurBttOe5M7dSkFTuf/QvV3ILDJ
lsd2G7pSiqZOZqSgPk9Ddm8+7QcCg90x9FmzRs5cUL8xqSkJNtqIGVKojLZZ
ghqEVABK+to1RpBGzOqbGrUReKp6xwGWROG22tYL4EGRUTnkEU+Qh9602m9V
YvdzwJk5jp8A2zPD0f9TdHeic2dMW2oETA2/GSnCjV2MzMb18R5WH+JVBpNU
ElCp9U+T0pVeFrGUxhMGssetWQGhDaWFT65Cs8d3yg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Iq04CcBGE8SRokLycXULqctut2U7/ZDZxZgbAs6mghXzqz3o8Jd42lcJvQcQ
w8cfgBGoC6Pvbne2UowWAZItoM8gS2IhnLHVqWxvDhEsYnkT6bBllz+ldBTm
PcaJm4+kDkLDaiTOeU6p9aSMDmpk4qBvprnpIAHPPxnUJaRKzV0FWkTmd2Oa
OPVR/brLzR40Fnd17cWa7OL9e/Y0mv1eaXZKcceIEOndM9Qniw7XoeOTbaiA
TCV0pziG5s38E236byw2iY29VOIx1w9/BHApEk36ODUaMM+s9wcT+Sv7sgMs
8npuH4Py8DYh3yCHPdcv7ZO/BhDaxI6q4CZq1k2lVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MWJssqn5u1Ob67rNq2W6feCN5EpA/OCp1A+NPMWJBZb74XHqQ7hjQGd6+UG4
4CioK4GvfafTLbU2URnqlx3V+YMbjyLbQ4zRJPpRsNxmPIaNB4rwNcvF4/i+
JNkbqxc79k6Qd+5icXq5dhHMvuQgBKY869jiTRy+r6EWJx1+88s=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Hv5xMmwuAEa8qRsOQCVx0+DwPs7RRaP72lqQz9BiVjxxTw2pv49RG2owXxdp
gWPZjAUxH7SyGDYltqArFAERuN6J4Ju6twVYTI4Z8eFWgOtGrLVqSD1QyvJZ
6MQLNRZELuIvPVVImiuTuXeB5PYilKDjjIifcjKZMeEVyt/yihBjNbYWI2WY
tJ2SJlrNbVmcG1qI71QBf9h7hsIfaXXxWc0X/8GVrb7rmqbEWAKk6xNMnnmm
hLbezNhbNt050iQhHRGOnFos4ym/UQhQa6prJ7wcbz1cis0mofBGUfWhlNpZ
fGPlHlx4vtefsYcABNcqTrvcvI1GIj98loMNtsJgOAZP3g4zsVJu4uBttbwB
ndjDEFrAHaW1KedyCjE2Xb2hgWwqRC9cMwxh/OYYQj0ZreNoH3pxDJ7APmzW
YCsK9Sfc7tFHJbHO7D5HlLQD6f+5a3Kz/cwG3ufDM8IxT0gRCj/SfC4hdNxW
eYZXNuia44Ln5p2zyruu2bA0toM8Da20


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EXVUaPU2D4CZHmFXOx6Qe3OzqWLmlsivAfR/96nx6zN5HAx006wC4R1IqjpG
cPUNr4h5NGUGzf7oWtlAv192rR0j3tVl6sg2h60lP86igJxC53+x962KSzIt
VsyRKNzEddqFyj8FrRyKfPMOQWA1Ewjzc0cvuk0hRmrbedvZw9w=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bXIPGUf+e72elM6Ab57fvH9vmRtU2hlt/l2xgzdxxhcPZMdzifX70rfNV1r6
K8l3URa4pR/VYhu5Fy1Y7wsUoe02302dflsLCz9jVOZj+sMJsN+lndsYhr0/
6xFoWlnGPtst7Qv68slLpGQgBlyajzrZ4dl4IlScyMSViH4YDmU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1360)
`pragma protect data_block
PeMgT7VB4or8N2N85o/tk9JmFLBOMaqXZB8A0qw3oboXtZl+44q/VWuit8px
dl1bItx1PxNDr3+ziG3IH/rVcKjkvFXvrMsc98pmlvQv4kJbnruVKcpO9V4p
4Na5clnNUJgLCZytK3oKkGN2Oi5HzG7ggsoT1hwCs+l2WcyuHgDbSB7TEv7m
UN4n7aYKxAc9EFGSUcycmUKq0x6gY/oetDenWEQHH+jzAN3qxm6TM7rtkB4J
ibPtT+UK1CQV7hQM8mJndkszWppYYO6+/qvyFNo5GaVx5Hoyn3BH8yRlJnF1
ulShsUDkf33LV1PHW9lYjvmT1lYZAymYqtfkiEAaHZfLUYhQAtZws24Yd+OP
lXimDFe9e2jLcZYlr2oHw8KGpQ7woxWTXNayjp0Lku2tyV+LyLJ86E+6CPHx
BLdm8ioD0hoPdyHaBtoqRgA2s1OcRYBXuR6XpeUfKaBufROcvkyInYSXFryd
c9sUy+j7vSS0J8WdqfKhvwBeLtd7AdXfWWGz0SxlY5NYaXwGvrm6IPjLhHRc
WXI0aIwloWHUk52PPQJXGsP2jsLzsGrCzmx2aL/IyVBo1l2vmCp1yx+kHqE/
oorbOuOggDv8TMWRrscQ4rmNJQSfvn1MkrbPBAv4lvxQubyir8LoC+eONNfv
U5uXbEkT5yF5iyFGWJxh9ShvHkZ2U5wSPPQCNs2MFEiVcr0qf5kbmWXlrwuF
B6HUj5xHkRsyDh6kNdjn7X1IbUpP79/K8WCVO5Dr4jzQgDfXRuQcTSJcyzBC
Dj4+yKSmrLdy1aEKAlJgC0lQuG3S8UU4Zx65fSW0wACGi71Sv7WfY6p5hISn
9NYn3nTlglgDjOaQTK+f2eulhDFAC6w1BmcclFpI+wXiottZFEjccltj21X0
RQDlplenZFlxRkX025BVrGoV+UtZ3RLehnDIaoOi6u6DCk8PIBRnaTrIAyqF
FzUmIlFBVoS4hu5ZjWO+ftyzPy+2VxM63kX6Kyz6SE+E7JherLd67/R2Uxc2
3SAuKNOCNmzeM1oH73BPKGAKLELOGHSUqfVj5d7nRtNenuEry9wReKCp4s0z
t5gWjm+vwtOijsm+D1AqoVssj0a1DY7y3cv0BW2ylY4ur/s8p0KDZbZ/hrdH
mav/xNMkJxkT9gf3uxJC8P9NKxL4uav95Kb1pYN1yTlG1d5Cvqf/q61ib2V+
rqijKnoPNNsZqYw83nbksWwQ9i1gaarYb5lsgKPSQ6ucSDbOBRU/PC8BGZiW
jWMZbOnkT5zKwZkxK9gy3LYLACYrzul8jillxSW9xzBdvBmQY/Fp9EvRFWJZ
UfbtcgwMuJ7zprgSDQO9KWcxwiaRVeepbywc6Qdq2+8Ca/Y3d9n+657IDYC4
3VdcV3pnKKYz8Le1TvzYOGlIMpOrOpm3m6EtAM8fgieMIKSO5Ii9NVDgcV7r
3enw/8oLg8mGvNRsw0ZqDJJej3wWmYV56gXmcsL6BSqZVf4hYXRcCqcPM22P
EwPlZ3a+3MoO0mj/NmZtRUvTDLI7kzTlmFvqJVe2VpsXknZjMXeVvxrkNo+R
T5wzXJOoT5t097ZNYiLer1jMCz6rdi4+aX8ynGQkBTsBhmYlvQ5ZsjA9XC9O
V7ctYhcTy/WGsqDM57yQ93oeUXVKRKmLM9RyjjSS73PfxUTwLDh65DVeYlmy
ykahhOtslA+hoMNDNFNS63mIkqm1DsgU+1Wgot0xq+Nje3MN9s8dIYxNmGur
uyIf8/ubGP50H4/hL7EGR4gAmybI8k3eNlltuoCjmeyIBKxtqmhMnNMCEyYa
tU2vNxAHc3BFZw==

`pragma protect end_protected
