// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
KTj+OZxsbWF/Xq24zC9J9U2lhhCC224+WXKEc7EejgNzpikhwHO/OWo5ZKuBF9Ao
gkMDwPcFMciZEN6P2xohfmLcGj915608XPjb6W4jf/1+bA12hs7h5rHWhfc5k2HY
j84tUA+FbDNgh6J5xAaTutrIyUfJyDHF/6DG5vK5cCU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10560 )
`pragma protect data_block
A2ddJhXgK9w+i/ukI4yiz3npBmbLBG+yxLp1RUieDZu0hR99Pi+ucgFvLLXf5jhX
k0KZ7M6a4NWavk6VI4U2owOnMlOiyTyByT7q4NEUMuydnbqA8DsVcB9RxDwoU4HU
9Se9h0rWYNhd8XyP7eaaJds2duPuM3qDBkF1ooboMYWMEsOvNRP+NFWhkJ7CsPpm
eI1tlZz6aQqUs9b8zqsmcs13caG4ITEYBOpUx9m3qqnv9wJW/mv78UxtE0Whq/Qg
9s+MkCaRrFS6kSPVbgPEIovzGkGq7vkMYGPDtNufoiUeaKslzME4czXp99UnCcJU
v57Z/gSwu1UE7pKMAIunSOH52Negl7L7yyPppknQAYztQoJ9vwvNtYZvfuIunlWr
QKpljW8dRmf8sY+Zxl7Qgp/tPQuO2XZzo2599wBsE1e0Rg3teDPXQjSGwTxzLGYK
/X2EFUYlpw3n9y/XNqntHfKoBgjxhtsyFf8wr/M4p96DefBdFKrEzSyauIWNKZmJ
nkTqIi+PbkvmAjtvHI9BcPiaYbagmQEyTpcpGqWoKjw9H22iRkc3lmDwta+O2OP/
Xw/rTXzDsM8xzPQCXXzDONjcO2oKs9ojO6eGuHg5JGshu4EzRPSlIAX8RBxq4NFM
lcHcAacC/yS/5o6mZXIIZttHb0cMpbINC54OI/YAP8xq0dAAnUzxGJhbhlxFjUvK
lOfUEvr4995Tjr0WEYAwFUnOJjIRAXevFWtk2uVwGxW00uvcqwD23Fq6OS7xInwM
ZlN4vDGHjeBZvuUqtlg9BegGWUc1hi90BMkhrJk4YUK4X91J9WEI8k2qD16UJdtH
5qxCkCkk3miuIJDh1q6JJUBy7NHz0fiBPUQ0FAFUErwe9ECD4HqSDTP4BE8RpHNA
VrQZqyhMeP8QWYCEGcT5JbAHF172z74emQPsMgFn3DAwzUaIT0PhF/TWGoy8sv/V
iDmHqzrdj1L7IMFCKIWfg5fMCI1h0qD8gk5pON4AG2brckUInvffXA0Mppfpp0mQ
LSjWyh0/3cnIwMpmxVxoF6SQNuEYTFrkpNPwJU58wmm74WTAsXuxROYwjhlFJqPf
S2v1hN0XQ4mgtRxKRnw3IID9DuvmOJAjAIsO/CqAB6goNOAWeRmuC9nSSG+EsAs1
KZ9SfmZZgted/D+kbmVkeVpUZNUJJ4wkrFK2g43qZpAPCjXWUKcdsxBT7BIwCL7J
6Rz0s0JxU/rSTZQadxRA8VgunrMXJZRxF/Y9IFKl2qU7ggf2+ZGphIaQk8ETue+a
TE77ujYsT/czdurih6ERtJZ+FJJSWLXpOpd2S5lOTPd7vjw8/038ab864LecD51f
ybJbcTj5d5UQTCygdPXBMnamNV7lG5JARnxXbhUILzFDDiCdjPJnknhOxgDYG0sx
JUhyhOHbkAVS7sCl5L2XXsQKc0eGdY3s4J6IPbpqGZ9TwRRYiwaOtZq7ZEcnR1a2
+9YBGippoMw0ICesNgVbpTBO+nXa04wA9RLvI9iGGHNES271Aq905cH60AWBcbZH
7/VqqbS47pKYk+lgnbTvSavuJlxaY4eIbIt1ZIqCArYn4xC9YHvGRZLm42eqo8Br
cWrAc3nCXAwgSZZ5+oN+BkKm+tWxr9682BEGHOjtil+5/S9E1UrK3b4i+qQgbAjE
F4HwIlXrwLIlu8Rt1TUsuhvnnadHk5dLAV9Slo4xuLdcMnp+rcQTe3ALvbARYm3U
fionQffSrXbyuZ93bKX6ToqQiN9SlU1dS/fnfIhEB89KsgaevQEi2l679NpzoTEa
S37YGmStossTIC6qq+352g4jo0icnO8uetXN1vfJzKBlDtvjm1K/hgcA3lL9fSzq
Ms7Yqa7ZG5eIp1g4M0QOLNIJLzWWScyAQwnlNYR7GjmbLIvzoHv8lyqu9yOxqXFr
i/YtAMuy0A1WBi9Qrc66kq5t3Qq+EXNlxrRC25YZsHl0SuxQyAxTUTGlyRsZVwLn
6icQcJI4tlgLVxGCz4YY2+Q7eRPXQzCcg+RfmsTmay/VK+8uA9fvG/AVJ/lNFrVY
Fz8i7sUneOJV/ZiOanuuBRp+euiby5AwJsm4sL3Du4eaS6vCZIX0L9kd/+Wlyrjh
uD2WUKBbJF5kLYehmtoWsGcw92p/dJwoQmGfvWWhQosDAjhlw8lQHzvYr13tHw4U
TRIta87IB7jSpJFKUbUdOBfuZY87BA14obWmkc+EQM2Y3OpdM75rWJ6ugYzlmeJZ
dqPzpw1fIpL6f9iTk+Pjc67R365fpmw+sqq5+i/BYLTscOg1MjYZFZKeMn3r767I
yk/iALDI/U2pNkF2kg5Ru4Xi36wj1N5Q8yoQ99sY1rnX5xGELrTWHfmBKFkoqDyT
YpbXR1p6Y4oo8S2KV3Et6IwcgSmusHH8ZcppQbsizKd0qVg+Ll6s60v09WKuHrO/
mlFftJEgGoBIqyUBV2vBfsN2v9g+JhUCsAybsutCQw/kkoJBnA786LsQ+hqKNfp6
sbujzQQdPLMRB0DGn4orWDq9Av4QlO/SZuqebJFZMCbcsiodI+VeQo9jv0XMevqp
8RIj3DuHgG6Ti9bhewjoythY/HBRpSItJx8YLh+akh4KxZrZZjp1vPbYZcbG8WIt
Tz+8QepECP6fa2UpL5iorcSuRMJIpVt8xTNPTNNAOUFYdYSf0boUIveV3JhvAKZb
mqC+UizYAawadOvJvQShk06Jb2yLpro/jSenHSBBJODS2cLxvkyHNmdsRGWSxAHC
O7YF0Ea/zQnWt779hYS1Uv06q/vhrM03qSIWhFVHoICyvP10UiqJE4w7R9h5MZ5n
aMKdiBN3Zwfksh+cK2FV3fSCunJSwdv9dLttqxPIjniTeh4lJx+3e7fhL+q+2j4E
zvCrL6rPTl6AkclX/4r5CAFdu5riQ7TRFNYUJStoFtNdvD/2VykOYsuZOPp68tQ6
v+GqelrwaTwQZeOqmTn9b+SBXNhYK2go/tmX6MZZUtXM8La4zev75rlAOz/cv1rG
9Z6BbYhTjOQlQp6D4bL6fStYk9m1TozbZH8yBueaomz5HQepy1QvK2e+GTZG9xGf
KwpFgYN5Bw9R/+EQOEB8ARo0/cPne4k/2rWmS1GEu5siUjHGd96mxMRqMG8tE9tm
ysASfgEWg5kILKWLDdER4GIAn8L2EBLCXrXJbnNIb8xZxc9kOFE49v6/Thd49B2r
uVsiDNtbuw06WviwyCDA+j+l+/sj1MXy39HPDp/d31YoMLyZCNxMahyR1yoDQVVG
l6O4VJn5AqUrj5AFKuiuKhCbqtPQa27prEuXI8mmw5IbYacsEpuc0F4Vb8Ufga+k
gOz856kcicks80xFRxQXRJtONP/EDvXGQY7C2OyEFH6LBJY16TzHL4sh2ORyxi5m
Gwz4qqms4KbQTSqtJySOoazT0EBN6x1abZtUZ1dgJ90JH1Rxl8+9bjQEkraG9JXh
mdDxOCkuXbehB8PYEQ9cF2gZ4Mt2gcwLuOgDFgiydHmbIy1EoXYs0dH/Fho992qN
h/Ei8w5YVRA8GtyC7Di/A9t7cFktQlHek0wT0r7F+RwodV+usxUkWebvrhBnW10Q
M/t2HGlTSod8eqWv5wjny4PB3E0B7iW0Eo6oV6P4wV9hlz2tvRLfzPqnHvQP+60p
HAscLDp/f+gsjR+8wrL03DuEikIO8FMuGDiPLuz+w0sT0PRHKRjNLP57ADX4tOdb
y+hfBDpOj02dHKIOdp8ZMNLRjZuB0uFjmul3upUDZhnqSyaFxIw+Mj4/jV18To8v
reDfwfWfOxfnkovWq3l6lWGhbd3u2IrZeN39xVS1mSCObia1/CNqZNhF//2Snjc3
bXOA2jkb0NkUK2iL77CaczBuxTsldnkpCpnr4rBdrBKOGFZZQnIHEI/mK/u2shnH
ZGiPBlSVZEm+plBeDaaVbHp37Q1NScdi+CL+P4hdwop2wmudMLz82Kp2U2+QFpzV
XD657tUdW6Z9tOwhkUSQpjFiGytrHF8R3DBDqavEEp9poHl51bHZ1v4INGer5zt+
9J9/dSeOW3jRfux9ou4BaQxQ5h4Ztl4MYqGL4noXCUcI3yB6uBVpwPai/vKRO+PW
/3MXsfAKZxfhi+ewq7xd8t818SlbYcnKMUH45Cflkdgl+bljjYhEFqVCtyLQS6n2
+JRjghF4jqis4Ew3l2iodEnOQzz5D+OF71Kc9Mi1fQhIJefRMZoOb/PSKTSd4IVU
XrYV54KFr4HF/wI4FEKO7HtORVnvsghZT5vfhiM6/7285K3L88klRbpWS+jf2z9D
g/sdnovNoBzC3M6w2BCRR85LqU9AxcyQIhudu8rFf+QAYKqrCbkKROMOg6H6ROKK
ttpN0ZYT2aBBb0owFmVwr/IjHGoJLYvrvbD8zBHTAMa0D2IQLZW0LiyGmHtKB9jA
q5Z7SdhOS5R6IAfCVJhky+AP/v3SmlmMyM4ruvODMPE6wx957aDEuXXTn7pVBOvp
9YLrAuPtWx1sg+Fl2tHHZwF0niXIxJkrVxm2xd5dkbOfRAenBgaxSvsvKiMfqzsE
J4abLjULSJx13KnGasTKslw3oknNvezFz1xNDHeAlhLElDeEItveLSqeVB3gb/gw
uw/ppqFFqOvTnN6DPdhoR0hXPWNSaqahJIxrLYDpyjhIVc0cd36/c6uza6fHa0bF
tXCSCeQuvjbg538NNWH0WMVN504b9SfmK5a6WMwEGSz9OQ0DP6lhAUQGz5w5I7CM
l1fFrsZ1FhoqdEi2q1SKsusUVoChECrjHvQEIrbEzsANfxOHAziRgQn2G3JcgO2g
meaJ5tfN0nXyTXKCRGCBbBTmq988etF+i93GPYuXQyKb1jWP+MFnbzkHXz2Fy1aA
08sC1v6SYoAoJnV8AEF/Kx0P6RxcQQo2imZDJTUjW9CK39LmuFzIVSu5Sqwzw9k1
i07ijmgcFZsFtOhE4WHGCWeznJ1KyPoiGoYiRv7Kz5MQAZkQDKYbKNJbeiMk1ACG
7iieG2h3zGDTnJSZBQbhApObFDJA/BDWMvk4Mp8LXSWclItZ4yCQGzMXpFY0MIrW
kKQMCkXYJp59ktD53Is8v8tQ5xOrnrz5qg8NproyGkYSfS/BwARnLnFwW1x6Nmo1
uP79nIjtOhU+KbFBTvGJCtIP/t20WfAUIQfpoFrvvhxN+2WIbVE1eo7Huos8RBIW
gE4ojU5uPN0/NIW2CelJPcHr7X7FKY+QUwal/XEFFo34W7wSceEHpmqfImYHUAtu
KBy0KyI6ntYEZ9Ol0FwvMGYsBZH8alEG8AnMmbR+LEcOq1bSsnsSG7xrO9ZeuRTo
XHdSUe+fNSqVx4v8OwHozbdq2R2VyHUF5AXuA7Ng4mqnXU0199A56p1vTm2rPLqy
jCwnCtur/F/G5qW25XCH/AyZwjWDy3VKn9Pxb8UfJS5prMUm+lTB2m6p2CUnCbp8
L/Tv9hCMTHsKdK91pnlOLZOVrgbxO/okvCb69LokLAQ4Bp4N/nnQH+Z6azknT/VR
BN8bOHsG91JtgsdI/qwMxNqGoWD0IEjwXORbAoOBqI8cOl082g9UVUr9qzf1lgWt
7jzEz0tA1Hsj92XYB8DScu9OWDAhcY3vL5rr+MNenc2NWclKHG/ml12keA/eZEbK
TGtYEMcTnmwOSEDlN9VX4ihEJvb2pM7FckzahMxroGLxNIzk91xw7gVNQThEq2/+
6WDvQe4Z4hF7he7eVF2bKxWL4zfZzHqDovNgfNI/dPYfGPC3+VqdWMRc5cCM5GeK
aW/CJ1zEq55ka+iXTYjlmeRlGcTqyoanG04RahgjQ2ZoWLcAUA5w83vAxUXEIImK
sUVmqluKDSS/QeqlhoNzev9nzDecaZBGHRjkrh6wiJ8ASjzjaaSzHcnflZ6fy0OI
YzaLtVlu3Gf8Th7iik09F+7g+NfgWTbop08XJP/lpAlKStZVsmqfFTnFP4Uu6tS2
rkBEQfgo6WcO1n6Iexjcx1rquEUv+G0VVQ5IzpTc1unnepzD/67b64UkXYD2qtOa
4Z713oWaPoX05uhTjkKjJfFer84BZT+qzFq+QyJj6W6uslsT7uI9K+fMHa62ujLf
ujfIONFt8SV+OUQaowMhriEMBqlKgaAcpErsoc9pn5rSpcgv7P3L/yKkFltyXrZC
QiHFnIZSWZm0jLbYiPrMptGEQVdKzagRLoaNsUh8aTjtQORJKWyICZTEw04qArR9
nUMVhR586eOBrM9q774GSlur1Sf22gUZzLSMMgYIEX3Iym6wZGTvi6u3lEeYH0yP
aFEO+Gkwss4Iy6GgAvY3reQfvWwlf+B6ezF0rYxFbGrMtX1/a308uija66clDgnR
sdUa+p60Qh53qWsy7OMao8qneIzxLSEQOer5DMbocgMwH1wfEApx+M2JhdIoB7DY
raxEYG/gFiDeylGoU5BTx7o8+XBKXUGdcoXhNslfi0arlvULR+xFEKeQapDlosUu
QcqXu5esbr0049Mw9nlaxFYKwWNzb/HJmUGcUjwHKRL28YXmWKnk1eHERJBOKbhN
nQSTQ/OZwd/5XOeIvR898E6z+QSfAgcf1lG5szv2XmuYRKTclmSUWufPq5/7B5KL
5jRQUZ9MyxaXNtHPmXJL8dSdh7RmS4swip+sK65Vi3yf0L4tH/c/0AA36kP0RMPf
ODkXthRB3LmT92Yx2zduZTs26Wm1HnN7gp7vnwi8IMMWbU6QDrGXOFR4ySr/O2fI
GhUfFdX3dj8CCf4BUm9YREti9pqANAWpGm+P1NIFwlwbHsFXYuGXuVOcTOHqkSp5
M/nS5tkpPpGCl87jtaP0ivKvQb6V/be1j27nFt31BWsU/1ShaL9hZFLtPo/CQn0r
i3hVpwPOX2z8UnGPubUW2Qisou2z6FHODMwBJUje1G+NqYQ5ZqLMh6Z1v/xfhyT9
5472tvalUKkh2iR1EpK2A57pPgOguFI/VdkU0iqAJsUY9GzmGKtzTi383cFqMZZ9
V8Av9mv4Fj7jxi2DiU1jHUc4ltLlrOtl9UKJPsXu9YXBdXrd6M6QGWBjVcrGvucF
HqDKOg5+MEJQuXI0z3vybDr7VD8a3f5SNtH7cmyufE/qXyyKddu31nBMqAi/cnWu
xVvYcw2yv3lnM4YtS0otCCCpEoRg+Vee7BhkPY7Ep5kUJOIyyDxG1xOTqomFUofA
+iTOewINzUYKWozSfu75BkqHtB02+W2gQrBRmL3+AKhBwxiDWD51uRfe3gbGiap6
egiYdNVOvn0tfAtYQL9nD3lbvCgpJRVdVCnw4HAXQQ4gs7/eE/dzpTORegfLMuc5
VmPQdgwGRuaLiir7R7rTS7PEmfYTFHmWRc5to1WjeBPBLWnjACjHI7oZC27o8/mR
jEps0sJzPFSYHYXIsh8jD4YH/Cf/QG6LEu9ko+O1ZC7/KlZkieUaDnwezr381twv
KV3Ef/SMbeXP57HJaLDn8v/9nslnY70Jsskdqogq01ktOnZ2aP07j5S2xEbPhz0j
5OuAF0fujYZ/qrfjR6RNSQS10gv58QOkuI5F1GaLC7MgeMGSednjt6k4BwvFL1Lq
P+QGjAXcE4SD4KYodIiM5MK/DFq7bZdwCkwrJekUckdtMspbRPCPo9msFMJlYe9M
vNBgdZbhVQOJB51T2xBR9m7l45lHX/RsH08wL9oL4bH21VdHsuAe/o1UqrHMoNAF
cB5QFSMRQRhi5UJiX8Jlp7S45aS0gopW6kjjopUxNBcLBahFqZ1AoCxJZAWVTB0Z
yv1bHtRA0pZpglHy23RpPqO76axK7YcdhUlSc1sdlYB7jetj04EPx085odVgN1Fw
wf28GnHNbKcaMdHwC/19g5GdKh6T7+widZWJXCoP9j2EsiG72Fjiw4MDRtld0Vfu
gM+tu8sKKsI0RbBVT1CXzT1KIazqhDcdegLjJppwrIgIBBJhybvBBVx1SuzPn3Hj
TzXrwDp16pXLpJhs6jS2KoNFmSItfXfcr6KollMOuERQ9u1Pvnhgb/pfecdOgate
Mpd91Oba1dMSQQFa7z5SkmuT8XhG9/V8bx5oGHcpV2FoEMyDPs157/Ptj0Uw4qt1
uNFCn7MAUU3cVtsi3Fk3W2/unGsh63xK85W16NZ9981CWXhc38udPAZO+DnldaOP
XD2rmzwEA2Va5cFnp2DoI/4J3c0SiV7MqEUqQWeQZclF8waAVU/koK5jiTPSDWlo
1fOKf8CNvx/5SBq3+Zt6w+3Lt4X6LbDGe0s2jkwRI4+uWp8diWPVUYqa2KvAIuI0
YAcMXRTAH9CGyfj0Myi4KpkzYWUzn0Of91cc05g/3Z/8VfVN4soMGpU6SIiSfLbM
a/k+SotdJxm92XoPN1zLTAxofW+rZlPxfacEA/glJjAIrZsKN8pei6gdsHK8BHj4
u8u0zhxbNK7ePj8M7hUWiNT17vPja13LwfkWzbByYeTVh5pGN8lt3X90ipZtrCjd
NSWh5DwmknSOBA98KP+4GxSXpNdeTHhJfwBdgoMVTDhCNmEkvLoKUD4s7I+JTZU/
SMyxZy8XVFtg7lRygkXeR96rFH7iCpk2Gwf1nLiAsJxpTwXubYA8pJZsOePKioPy
NzNwCK0kRo9HEIqQH/qbDiW1noP3FsYOVqK1HZ3+Lg9Ey86Qz9sCeqjJ4wAx9Edm
2ZkRbi8BYH4+CSGxBnMlSnY+WHLjr3ER1jzuWe1c+GEceeW7CezaoWSsIrWhGO82
VQ6Bs+i2pExaZiFYeBjSsrWw3jZHXw9rz/B3n4GJ/fVm/2tBOjTqCvTu5bXD86bz
cYphgL9ca3/FH9jurC38ga1R5qkQzVOMUblAEyViRy5vBdwEq/M6JSk/zF3M56q+
slZDk4xalVXTdWjQAoz8xNYuBYsWVA09/MSgBzTU4kpiHCb1nS5qJlRJe1gPktHf
qa5+N+hb1hVgtHMSjB/qKX5//+9z0wqKgPkE80EpzIlUgqj0oP3ot/HTpUXwlNev
PdP7KNF6BVPg34sIIogAVNoshfRi3CZWA0wKYAKNAU8Z0U7xRZREcJ9EFV31RdeW
j5ulXbh33CUHxfnbqdgSwitMj7j8sG4rcSEZVVSpLYu5PKdnnOm3lp0vRCNFQVNO
rma7sE/oVCtGExsZs31ZYdoEVcHw1psNRkd8cCoidGgFDmxfasYiHTozrPEfVOPB
QWCF56E1Kuz36l/zEdjKw5ocIZhRq9C8UsEEybK6H1qXTnoZtL+yxJqi1MrbUsph
xlUxugZal+BxMZclQdewZF16NFrZnJ6eyjqr47f9J5LtSE+VcvP0Q84vVWab0wy7
UrJ5uqnXREIbfiGpARs7AsL4POXMUplUEckgeYf+tvwtbepO9/Bf4+huMQ+r+ruR
p5w8h3lQQdu+0ZSmeFqDQTz082e/WqaeRXmgsqCuY+qOQMMzMCx3ukdHUcr4CzNY
q2vDpOvKhw+NJ7ThVxcRwyK5GHbaKLaDioTN6FjYKdkuD71odWaXdcSlwuXbHKvi
GoEfT+CeJDlD/V0SLqQXE5jQmhnU3WFb1jALCKnT44bKKpnQpvwxnJQujDxQrDPU
+lunYUrT8fp+g4eM408vWLRHcKIbvkSFSaY9xQViY/6vacYmKbN/A1Xhu0I6K8KL
E+tCfzf4jjBT2eU9M9JrogaS24U8PvjfudW/yY6BGUQYkCyxcVxFkIFgOD68pN7Y
oCOrJbba00LpZEKEUiiqjmNV7wAGwIW9EMpQU6pbK/hOCBrjNSb+gKY+8uE030z0
214ZLYOIsKDXxpROXTClmi7ue1gaitO/jSo1vtgf3RlHl/7bn1N0Phs5x3YP8wdk
K9noFE4SIGbdGOtHwXZzPOMWuMw0MIlmB+uu6cPdfRBRaggN/ZCaW4a2Y0d3i9E5
uxtyQ85FkDS7vc6Hp1vALBHlplGYO58XKZZcPBDedjkM8CmeHWfPB0lbAR+TORKt
iTbn7YlmqOB1vDdTnACxKU4r7N2Wu84QjDSGVYBkKI9m0kVA29LRVF4D5h+oyzfM
5eEl3Nytydh6KCPbeUZ5sPl1Gzp9K6UUZhc9LZrtEjobTlG2EnaE154vDJLPc7O4
HlbY/cBhpK4ZbwuDMs8gsQCleA6KYHXSPaLOObVrQjuGQZhfAlN4Mnhbtx9vUTJ8
VIkKHJdewujzCELou9h3B2jpmkUnCYX6Hfv+3tBWj7ms9gHzFSFLHf5VOG5XsnUc
IPO8R0ifNsBzVTM4Fvf8G5/Ro2Ml1q81UcrogUjPi5zKgvzVFbD00ZyA4eIUL1aO
ZpCwgbOKAHud6h09docwxrl+nkLWCOSjXL7g50ZCjBudNG2kOiqxcSODRY9Mo1q5
scsYVBV4EOGpNqMGwT3vKJ+U4MMnef6Vnb9EdYjv/YOqPlUWDOXtb4giU6xmnd85
0IQdunYYOBGB/79cSmhiiKulJAQ9m3aiYvPdUBRUBpz0uvsy+yEcDNufKqT6+0lT
7olYtJl5FIvJAStCOWV5H/MjH5ki53yirsORfkec7+nY6ZIRC2qSpbbX2UAc2Yvn
w7e+vgYpi7I7ueTch5apMbisCszxDsbU+J80r81KERMvGbTITwlV+E/m9+JSHqUS
HMWPeXVs06oNeN+QMF1BOK8OmjOXak6S2bLBG20GyW3IMu9r9z027NgnlieysC5x
OtN9schnjtgViPA14GOfbmxOmwSe1bE/6FbD00Vzicwostxm3RcTlgs17kkMwmmr
ppKnzgZzN29d0ZvFTBQBQluq20/Kk6jAW6israadk5vCMc+qcwzSRXlkLXPhTQzp
DLU5IHtg29jlIfjK7lunNdgAHo3zsM1rMM5NTebXjDUNcMQuvqi0AcNm/fTTs5vs
uOOE/rQdoOwEjWQsXbh4VRdJZxkQhzV9RPzI4yRtQCJ7CXO3bXCqis9X5zsU5YbJ
SDjRR9IIB3J4CUsNFT/E3vbRMpGYJNSYfqWN1NbDJ+AqIiLpU54S1Cluw7q77XfC
5SwU/BPAlyghUAprHtTCJ+Q/4jxr7YFdvIFc8SZoa+ykfjhYFdlz3nKMWpZ/eV/M
8rKIwizZRt2dFUtYZWxLIxv0J3Dlepp+DMZKeDVsqamQHtLWw+ewUnGnfvIj9pOJ
Qsmsj4YcI2/BsHl7iZEhspYLgiNi+qC53MbP/3lQ8d+lwtGGar4iVgf+UffD1QyH
rhjmNLm7KL9oBkeGzeUPw3z7YC+TpgkvwRW+W4jBrRfiuh7WdeS4RmwAHwFt6B+U
VTsJB5rZWulRRlv18mj/1sF8CYaXAJR+fW4YOR/2tTO0i/4Ossb768DdgxYWnER1
aoNspo1fam1jR23RlMGJhrGMfjLBW7GlYUWE0SzBggmpJaanDG3ZiPbwLhYVAiIx
eU399FPrGZES1ha0Q32YuV21Ci0Ym3lAN8Yhi/GJNkt6gKK5CCiGf34PEi4pZ3S/
Qv3nJH3wPSCBQrafyDoh+ol4l2ewK0r/DqOcx6tL9VxxN8wN7yXPFPPt3U0OflHi
FjphlphqxeWSroZjaMcB5IB0MfuoFsWb+g74jYVJ3mggayqSgoWAymU8CPP4tZM4
iou1ziYxFGkDyKQ2W9Z2DkCVguxYINOrd3htP8SRWqeOREAY/RthERlK1iRJxXJf
Bke7nopZY/JyEsEjQwz+Rbbix5dSQvcUCf4VRooGfFCcB92caQGZfoDnZw9NHHnR
omZqLXbNyqpalW5S82EGVQ0J/At4QZPIJqO8gifmao897a3rDEoHIn0A7pUD4DVK
YXyCWKQ0Ze70FzScJyaM4YHO+OfCFS+9oWUkF1PoNoKfEqXqYRMSvseZNdXfpVtP
gn7UHY7ZR99zMm3+Z9O6nZKEUFQHKjK8kY94fmEp2lIWe0PJXrmTYvuavel6b3CG
BvVqG/ShuaIibj+RTQbK33AtdzF4fRagD3FRftk4uuHl+0S8WcQz8V8BMjG13kod
7AEqHDxGEqvVSuFaXqtzBeQbBvWIQbkGSZOZHEupGCztFgqTxdgDohSQKwQaUF3n
6HBqAWkHjU6ntU5mZ6RzQgJedS7k+8h53SIe9pdl1mOIz6YiZWr1VZq2HOb/ZITL
JOsqFgCszRncsZ1B3HfHyFf9RkF2iRIb09TSJ0tE+V1dKpPv+mm91mfx8EMszOez
4QBt2apgIP6UgIn9XJYcfm2kmMbZ4JcGONjf9nNnd62ybSHL2urJ9D0qY6sNNCHF
p40pqxvM6R2wfNsvjIbA31MyHK7d6/mytYcyvjfx78QirhqdNQ5YuIJQeGHmjZhE
RC/EKQfa4EcLjUI4xPK1aAlLWNN7bDrsSUAzRHruwb2z1acou2BZdCZB4C3SaGtm
XPl3UYnsNOMCHQSaVzEvJHyCieq2QNyGIU1MmSXODmjXSenkYo4oxKho0GfzKEMn
+0TCDQzD1PNqD6Sd4T4lCGfL0f/Xn/EJr23/OqIOBCA0s5eTd8E0agI0bk5OQy3p
1lqJQdgq7fgpJAg6BHFhcUj5fyu7CkQ07iuVUok3YA29sTvM+VVFgcSjbE0m2fU4
1EgbOVjBnPSvps7L2IcM96U3T2vqpdRaU9FCyOQulHFIRdX2d8N8XeE1WJ4J39eP
y9Tl+jlqM1+rSCH5tIlZV4XuWhVABrQirfjVKHFcNRd8d3SPkyqyqGdz/bVvS/Za
E6JILVsBQNxCdtFkZndrQywWa3PQEctF+6UtScgn5wc6Tdz0oRwCdsluz/GWpJ4R
HbiFpf2O8oqcv9M5SsVPZWt+JvqLgXSKVJm+176o3MILpl/Bz5mzDWKByLSmBKei
DIUlJyfdbSv8pHuI6WZdiRg/BXOmc8zm/q9UF/Ky9ADYt2ZdBJ8NJVZlEYAM6MEz
6UhMTMqoek1e+4MYJBOC1B0mK90fPAkq9w179xTCkP+rRC1seuSfbFx6ORvFVZFi
oY1sW9pAWrmCT769SqR85G3Dt+JSpIqlBQdui2GdR17MvN9rF/rLs/QueVJc5jWe
E4nsmN91kK/wtVF6ztCnqahFKsLa+sai+MRlAB5O+Ohhrx4g/fgn1BAfYHTHsLFc
WP2RvJeRTZSOr5+weyYghcHN1A2PZxVm6YxFJBNduhAwOMzcBnipEI5PTzEiyLuX
+kbfq6uI+OQ8WoEV/I58KUftFyk7ECMpboyU8wLY9bi2J/Mr1RRaGXCw7/7Owe1C
xR3IX2NludlKAbPDwiaU/FprdhUU2sO/03gCv7irWjZ4Z5TCn6bIVJPqMR3+j1ZK
s+zaCtI+fW7+6Pj9Ws6YgbYMeb4qM4cGfoKzFY5pUFwsiIy0juLJ8YyN37/WgGnr
ZBj1X62tFqbBh89+rZE1M8iOBaT7PvQBUt11t0HAEqXlXDdamzZsvOlyHhDKPjG4
UtzkMWrDor/FnOc3iOJfrTdO43aGWCkrIoZCDKlSLNz9AQbpVdvQZMBNhOmMGVoD
zOHnZX8u7AQyK5XNeCSlNYEUsP4UQjxcWgn4ULFyPEdScSbL9vz+YKkTBLoh4ID0
vgByFu4f7wUA44eSaxAH2d3KfJtfcQA5a5ZbokZNxtu0tm7OoPBTMAhfy8um75Xx
Q17kI/UQtTP0wIgyDopn+cpwhq7q+Tjg1tq58HJSz5EsLjVli5DbEa8B7pt+zYd2
dmpgU0PvkwJ++YVo9hh+MLUWeoc2ALqZ1qTUOMEhXljLmZxtTeySG/onIQKDZHr6
GDxl9rDv/wnMJR50kPfyLMRWiALVwSVMETIMaJBWqJReJj5LE8CoCLxJ0ibJw0Bn
RrdZENIYqlErG1JX38S4gyWfY91QXTnpV0pPOY11x7jPAAeEc6RkKmhro2TaBGDS
7BHd2yBdjmFki4KJHuTAP9EzJi9b449dUmGWMI6T7Z+iCTcrirJQ2aoPPn3Eh2T4
Ftns66IwymsqjZhyJ5Jq9FXtkB9raJDpzCQtPdcR+K1xgVvTr7hMJgLCoSFrthOP
vvGyOdwNQBvb9j0PLSkhD0krPRmvvWbHJ0AJrQsK13PErmioaKBrCTfjK5loglk2
NHU09SwBgB/Ll6GLMt3b9wyD6gEGBb7nqKNS76j3pULXOZo1ynh9ue38N7uw2qh/
dCAgqnUIPUWQ2INS/JWBUG+kDqwvqoBdGKvXYGCXuLSYl8T6pM8AXXTUtstH3mwL

`pragma protect end_protected
