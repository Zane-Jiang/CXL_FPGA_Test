// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
M+4cv4eIwkUMgv5QOPpNCKM7k6/DB7Ifp2LcJ0htTIFbfVeNaTCeci1+qRxt
j7HNyy8LDvb92ZTllGOhrumrkubFbl/gwwUa6JvsXZWlnkV0ftuwsglZWhyY
U9zoSU8WG18JP8rGr86pNOzsGZq9KAcFy5uxOLoG9JKCZHojBeqOgJ2T1387
yfUJvH14gPlLDZKuSJDPIGIlats4ii0uxCUB8jyF4LbTgWzcTnrPe8lIC9dN
/q5Zhw43OyZL94HFgPejDOy+GEBZF4bFyVEQq2Yn0293FfPpg5MbPAGBinmp
KvQp3z7NzV5z7i7vibXK/D07B5miWkFzJ1xTuiYkFg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EhyLyQG9CqNoQKszQoxsJIgTOlCu3f5WAPgxSIumaNeNGhzXFsNzxibJ2VD5
GckSxUCdcM0tpM0qsYesxdHL8Zb0j0JYBjC13uqu9qK5Jr1LLCSX5JYWprMX
3HgTssgCHco2kabWzdN2snGNNLc3very8nelWVYHPMdkmXmWudd7K13pPgrI
seNbZsue3yjyLnhjSHHPY5zgVBp1QSOVbTQav/mHf0DgjxlmNOXw+CiD06da
+IuHpRtnW2VodpdzeU4zE1u2najh87i57wYAe7b2HbgYDP29AgLFXMWkUQEg
lkx/KzDQCrIAbYa4s7oPdgGW7aRZO+xbbV+XfVSnuA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l5wD8DUT37f7MwcuL3fslyCnNNA114UftJYaOUH8zxBekQkLjJ3ihJMwAv7G
9MHFgu6gasrxLHjiCbswq4V6WLZ9s9Y6jesTwNC/GAwrkrT+aW/OtN2tet5r
sGC3ZSe/aLDaaAK4aLfBzug7bmTa9FutLRB5mYVSGIab/4uqqIE2zHk0/NvR
/5sh4hj61z9Ufe7JgWmhKcFz80he/nTlAGY+H/0oZeF6QzEuuMELHaOWuvjN
plhDy6fMXsWTOuqiUbarMDDuIbFdjgXXwhtWIk01ClU3DN9NkDbn6vkYu7oK
BlVFvqMoU58fWfDVTPvks3E/EcUYhm/CriQ8sIMtIQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fapQnrn1rfUG8RCcFXOhgFYfehlrLI/V5jYQS49i//YK7ScLc24QIFc9XKw3
IHDqRYCUBlWSnwClTi1zx/l457AhS18+tplbLxeA6EqH2RnhyUyNxHPbjeub
BCjQOi/XNeiDz3wZU57+JM8GGhSWP3/VGWTvWplkICE03L6LLNU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
j9hq70vtPipE4DElg0vrd/OwkBuIuTgTb5ElsUMNdpmH+z4sRMBZ/a7q+rgW
hqBcPFsZm1Qd0XVtuctVKGOcM1bHV8Jwf+zMz2wbqwpy4BH9C9+MYwqyQNpC
osiYMEh98FBwEJSG6SBE3N14T/60EPlyv/vlYtgq7YVIVLbK+h6gIe46NmUV
xEpKNeYEI/KRuAB6JWiW1VEpBR5hJFqh2WxkfXhcDH5jekZ6GpbX5hTKa3sG
Ua1qETvJG87aIXfGTixpgDHq3l046lVdkE5VR3pgggJmd39M9t60vSMKHNq6
O9sc7AT4V3fgvSp5B/P5MpUdUzlRbLK/cQRSUn9UE6v4BeTcLFKzYpO0boLD
ZZD+TmNoMt9SlHAAnn3EHmvnI6tv6Hu3aj5PdgVKKcRP7w2j/WQs3aMfmmKz
mWm06DRoesXiBkoiVzOyV37Zpk35cDWAoxlumtFjKvFkA38SQEUT5ZfPc7WB
qDFdCuLePVrGlTGub9gd9QJJ2AZFfc1w


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ffQJSPGvyVAT4toh1pzra1OTWDhWB5FytDzjTj3Ys1sCtVzG1XXwF19rzLLQ
VuXw9M1VJ1QbQ/vVqqQmXWqng4WDPQmsHjhSCM1JMjL2JveZMIytFG/mxNgj
Ko+NKfXNoV76iusUQO1NBG+io7ao6XKJO6jc2eMDnCcsgJlkG2E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qxdBPFIhoCGeFmKEEm2iJ2IsupNgofwENBugCuPaTWvHRNWLecF5CloltZWh
auZ5LDC/PPBPBTE69vjKhpXBOlH+ksmnVQJe9szV0yBc8EM/KEhFzTMynNA8
QLejE0RIfIFlR1W0BYtZWrfBkOOD26Nfw9iTz+GpCfD/aGXhEas=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 86240)
`pragma protect data_block
46nRDURNw/kGLSaFzUtXAiXZ3e4aJKThgicR2u2OEIUy2yula/ftP66K5HZT
d+h2d/JTPjSQ67tMsYQ+uXy31LLRBDZNVuVxedsHXLnJ7tE+9Gv6RUfticzm
w3rOdTBUzti+A6oTFELSnWSEe5fWYR/QkPBxdaeHPBbLdlLDmF4J0U7a53xU
PmDIHy4ENHEkSsPsdjDBaGu0xCnfWSwNZ15dClZVSeS3qKC2CRH38uzrjrLH
jwVyO5D5s/VQb0UDWAWouH02z5iNlNTUvL1Ll0utmlATjWXBkBTH3JQfC3ba
DZ8ZT6CgU/sEPVdSCtDsJtWehDVUppdgpQEGj2rQ28CoDkPiPeTqNGMu/Mq0
tj8C8W71UzBLFYWOxcDyESpNh3BhlgkUAnBCpytFJvAafKWNyA4ZZl2Jvfyf
5kmEnum9AOokIVXPnx4Vdj5mk8W4lyV8GHvHGiytxbkchD4MH9nkI+hPdHmp
YzrYCiY9dRAICEgUUhrLeztDbnPi1lYpgVa3Wnilf8XmHF1hHlTHELcnwRct
lJZVjdWUUF0sudnh+VAH7Tq5JcdE03jNiY1noB1Z6Rp/qOC1iXJtQaUt92Io
gRzRv4O+A+Eh1TpHx+Sjiww39C+5yvqlj1IfF7Jz2jVvzkyBNiiX0u53gts2
4pf1CuqXQOrOC0WtOsGGQuPhMTNNTC0CqDJVIGtzASmtN3dw+KJx1p4rD4Zz
0CyMERWSE09oBfMCBEhe3gQJd7B0BcDqg4Fm9/b1Z9WjixsnEXbEWMHXqJHN
VbjI1Djpg7NmqeiCBCcoS671x52d50aRaDmNc8es07g8x/BoLwseoZarcOsM
Km3ijilInR4Njm6PnZSdi98cuvNNBrmv7myimURE5oE6DQKJ61fXULYdJg4J
+v0rkUXCpLMBxHKdUNuQ0AWZTi/Wj1VJbcI9fEAeWGUaR4YkepkiNQBKAcY3
+33ZasUwbEfMQddaKm2ftzIEpll5u7Fy9/LxCCRTItuHCInOhGx3HJJ30OTi
PTEycy7JKg/LNnU+I5G2vxVlzOK4ekMBG5M0JjbV7TJFsdIdJTSzXU98D1fT
w9MRf80TkaDL75NBuhNnq5mi+riBhPyjfFksMsPc4oLReBFC5RuQ/qBoFdUP
kc7EYtNBELBO6eBXPyQsujuPVimWrZtVKRq+v4yiqCy7wjcqAg4gIlsKZZlb
CxLsIrPBKIOK1G6G6UvITj32qM4hKm5aoVpTJpPUkyToK4qN0TzFMs+pTfuy
ozUNSnoispwCqH1MWZPHstDW5UhUzDu4ypj6RxJeA1wDT36VIB5zargr82vp
7BYZ7wRHjZvoA9uHRn2C0xHcRGaCR11zXOuzIYnkaL4lJK1SE5YgTF10/VBi
3Lr1QdsuposLweycwa53KuJwWSxgOlharwYoNK2ZfI1uNvoKJClCtX1mgWza
aSLSTjC58USfYopgD6I8ptFNWpTwK/AKElnX3CVPYfwU+Zmca3IQKU1K+H7q
U/G5/fhRePcbonSZ18/PElVr2lxUwZcdhcr8cq2930w+3+cYtyAS15+7gPO3
RC5Mq6wxROJhlPbRn5akwvAZcB8t3IYCjRlsNz7aQfRIp03WDaUhvVdUD7cQ
QquFCmMKFH8CbCu0c4rdC9+2FsoJiR4DFyMFvxIz2bR3FTAobBBzwo8ya9mD
DYcTJRmBOJSD+hRocu1vnhYjMtXpNqhdPJlgu+2qIxkpL2iszv1nZecbJe3r
wAX31g7qaZfjBfzSMfnW7M272+uQS5SaaA3FihjhRIOaWK7aPgoUvSCLjzpb
Gu1ea9j/pwYgqDwzlNCGbT/FlMHCsw6tjyZvvF86Brw/+SxhcArVFPxnhAwG
Jtarigw5SAfxOhHEyJVKS3LSdQP3gZLLQBr8gwP8MN3XrnQ6z12kHQf2JH2I
RUmrQA+xDZLK0FV/k27oUhBgYfUCry92sVTcocKGYpUqvebaMp8CWjQQaRTH
DcwSp/nH7OpeMyn4xq8gUkuUWr8IEvMXXBY4N6B43w1ygrqSq5Fkq2VW1WyQ
0j1AV8tdv5yO1QeZAAsUMwhVcOT0l/v270o6KsP4PlvT1T9tWN4EW5K7N3zl
Tjf9TzxBHqbS+u321p+gBDnsVid6Bntbq9g+9cO5k5X8t6i5t3h6/UbiJeUH
q46CmrLxDdtZ5szDEhm2fDIoE9Q/6L0WBu2zp7OSWTfefBpm2Nc/VHmLTWSw
kVwUXtrwd8BknEHx07FJekEd/pXon0a4O4urBAttyeyRZDo5Fb6mILjn3EbV
EYzW+DisSWA5DuwxUd2b4CzGyO+ZV8pamQQW2ZSFDw3q5RLj1MNeDdQFAOcU
cRWQD145rpjv5eKYNY0pGe7sHJN5VNKfgEhRnS59q0d7RlDA38LayZ/RBOGf
KohPPtT/pqrJhZoPLPJjcWPcbn3hhsPvxkDwnL86oeigsNCSUN08V7uOsF/g
UVu94l0VKXNJTQje1Z7q1WRhvACcnLvut3kmCKo30IpKV+yJ99AF4vTaY93l
oUY/1YM3NLEuL1Db7UppLmmXgyL4E+eY4KCweM6NQXZEOw7vUfxxXSM8vhba
qRjw3n7kIwHn0qORnmoC3vhPLwkbRl2dup2Q3A/RlLRFM+voGsZV4pUOpV3k
U1jYjN3trMzgMObZQI9KCgYKEQbnwJAJ4ewy4Xbwio7prVpQyM0D2PwbaoZj
k3981xFz+jeRyZE1lxpIMHkqj8MzWNtRE5tRJZiiNgefvv2WQBOOH5M5omIH
nmG0TQ9qZH3QphjRhikGluKnEhq71giX1znDjBJSUCWxexiABdyZIBa8YNOJ
ZvnMvoNv7x9SyBBUyekDZ+GiEGm+U3IgMbxhEejcCF151CO49wPeN9lZHXLq
EskMQwleG79fXxNNKzXDVoulJQETy8FwjulkMwQfMn8lej7/Vo7ObdQV0AWQ
top5qztsyOCLoR5cuepL89G9B5Pt7ypzkd65ZBT3WgcgxYl/kubbkMhCkLYA
Ryc8mvI0YBHMx6VAjN7Fr9hYZ3SHsWQVeJtmLIYgAp+qgDnlv4Rzo1uyQayJ
Azc/AysgnZCVVwtBWZ/tae5645s5f0tNrbsfyrKeAnuUjYhRCwxJIXZcFXrj
d9kZ0nfMadlxq3b9sfmGYsbs8a/QIw3xR44YXpQP8h0MqEu9WyP6nzNEPSuh
wg3QEAmmtJjOl7cPdh3DUNNvRA/pon9tImsbl7ZuhduGEiLcaEcYH0Rc32+p
xgbAW2LJcaSW4lZzK+iDrfOzVxbuvgTF///uMIKEyBkRHKw8Hn6oxnJ2YilF
2jfGtP8PVwSUFIFD8c/aX75M2Z34ukIxzaed8Hu8tooqtHtFPyXuzNIetBMn
NQsIUA+b9mZH3GlOUzR9VSpTMK6GHOikx9vzhnzsmAFLKjnqkFtD0LcUVfFT
QOx6/a5rKfXkwXqsTZP2HjFsnkq5JX68mPd4md/ZrmfRq2twH7SHn1iqsQX7
pBG5OCgb4iCFTTaodfMRMFnx376tV+234F4tYxVLtznAAvFS3ssMUFEd5FAo
ryAgQ8YvQ0k2mQuTNJ8OblDFmImJosPq3tmDE6VUmJfM+TVIWT4LQJsNpOY2
QHEdMk0SO4g5ANcLfmtj0NMBWuAtgXx8Cu9vXiMhUule92VeUJ+NA2IaFP3p
VR2Vz/+I/e7ZlsI6YyGYsJ8hcnYrVuU5/jD62tXXhCnjnnFtLcUc/kyX4rxU
WkcLDlBPiduTbg5BdHDNevxcq01X5fw+uU0i1HurBQB+5lx4aeZz8CFKpOpY
Cgg7un5wwbfpy+4MJyv6jAZxv2zPyETJD5xZZYbTPhKurlwf2OQVQwBqvsRt
RfixKL49Vw1I+/M4mWwuLxpdAj87PwR921DddYfrPX22YdYTA0AygqMyfU54
SMNlKBXJ/aLpP8EXMnmV0OFWD3e+O5xjhDvZaMxBqZGu+fXhaYAPg/hRyc/Z
Cwo+YpCiyYCGSC+QWumEAE0TBoja27j8aYxC90Jz3wKqIRNpvhlbxSbtnCil
1Vfz0NTDiUIo2wf7B7+6MnpKtKVz4ntnlpzmtsuJcfCbNbf78WINVWgnveYM
waf6QhCjV7IWlAzyWEH91ZrPbx23jgs1t/ya/LjGG62qOCi13qx9gWhsBOKV
RwFbi9/Mof9RolzFH8rMTFFVQJjYiT47iztv/IRB8IWkwLHWLIOCG64puQHU
o+o23AcxY+ISSXaVYwTB7Gn8lLJ34LzPV6yDsbqGFNBun+YbZOSix/wQA+07
CVdMgrUY6wa4IXlRw+QxnKXOlK/EMhPckJIgX1dLkkwznyXDJKfKZZUHR2GT
ukNk1RA2/wJF1opkQHjjPkVCnv060g/G1PScfl9LAUCfh9Nle6j32oEFPJDe
us7L4iAIm5RmKgghRrwIUDhD7+dAgYFYuaQoK688pZYLQcURxzMAuKBU1xHW
kKm1ItY6cej2JD6n8gkcylCcf5rGa7+ge7YqIVo/GejOdzJVvZaqZdjgt2um
H/09ZMpLAuj/Z5PoQaitCKb1Vtja8SGxOMQexB9Xwwf8eFV15A/OVe9KwG0Q
4okrLmm/eW3ft0Onj9+Uyd59QcSRVE93WxR//OVeTUnhv0UqXbZ4K7KN2WoN
qkuag7SgA5QMmezZOI3gk4/f5kuT0VaVovmm8Im1AkIcvzzcYmFgccT08cpM
JJ2FAMaGE+gUH31CytjNB7X496ow+FS11LZ8IOXGVdjMcoqCdb1CQ27LIlkA
Q6GKiMwsUSTCtUAhajYvjZbMIuQhkVAXZ+u+uJIlnaAq+OFYDN4zdhA0jShX
pbM1Q1kBLMrHX6yqfZ4Tuzgvv41E7+Ul4i3BKHJogV236ThZK/Xyv5ldcHaj
xn/9v++p45o5lelncWQtHiU+3GUcbeMyLnzsK3ag0b2xCb6PTtFK2bAK+VwO
qTgyzmKFyciIHQiVGVkaH+byiGS31nQcfU2Le4fC7hxWVMhy00xu03DPSw2K
+1mHo4lnTt9LhNJOEgHIC2IMbCt3dOXczdhS1T+MfNwPqQIXfxyVk9bZ/vq8
VXr0Ba2oD2hWAaVWBOBqXhfNDllJ9NEwF/gVUIir3WL0wQ3kdLRhnFh0XNfg
IR8nTYUtrJKgFjbIW6pHk6ioKFPo/3GZh6JDT85Rx4QwjR7XKYm2glDAWq+c
1p1lLv4RmluPeCHKGkBUylubG3cN2HC0/tyRuNOE52qFz77oTvjuF8Utq+4b
BbUG0u4+NFrNB7tG73GpDXZTnY9D+px6bi1JcNvFwN2hMB6N/TQKsyCB/IEZ
LOXXA4zkfot97RREqo94oRAn/NULbwOwPkjgRG5Yqyr8k5z1H/cAUj4YGxAB
5WT2hmBa46V0O5Bl4RJ+zcX4DFspATZBOfqGMptvW3T0ev7jgY65/o44qwUz
GO298V6IeT32+31Q7UR6/MKYLvsC+1ix7krWXdPpUd4Y45L+cwqM2YBW2w9i
jmuefoVZNt29I+8/g9YvgWjBzoMe0pAOJiU+HoVHMPhHzWAouq9CRFAFIEuI
84j/6DZo5LXg2BnFLJqNVqzCNEmXIXMaHS2/lF/iAHiBHn9mjNVIQpCr6g1G
wuTlBP5jx12mp60c5Jt2u0DSlV+/sfrAXa2YIGGHz2k3GfvqVsMRnTojsVhR
Mwp4bb91eLZ80cOgb2vSjyuaeyy4pa+WvOsuUiVdUwmvm53VtDn4DC5SVszc
uUzKqtyssvot1Gn0DilCoAS0St8V5IaMjaEAOJcxeJ/cXkeGYuTZzHWw87m9
5eWcO9Pu3EEs3QosiiyUlcaPvGxNgj3m8TSK0DcZzbVB62OuDywAHFe8HMK9
bzDRE8K64w9w0FPpyeVsb5QVFS6BfTCpqBqu4UlXqC0bcbkHi0dcix5dWQCv
4DXAA3oGz71jMQRhoHGD8Kyc02kS7cNyyXR3oHkLZFeEr+21tUCszIgBxn29
W6IP090TsBy976ul3QO5rtBDg9144SvlCzWVt15OKiKX9hB2JPbOu9ta7RzG
+k839p4oiOOUIUKMULZmGUagDBbXwLRkGcuUpPHFFWcIXGwX2WkluBSqNnqM
THstUU6XKl2j9EzIp1ztzzlAqUR6kRtb2ZWQw8JUYmIqhRB+d713zRAe883R
dzAc4a4CwKj0ydHsO2lHHzorXlSsydetFDrGAvukeuH5+aySDQOOh0+8SmjS
VJjG8HoH/wuW7gboBerkqtEgEl6Ghn8X1do671a2+Yy9OXFFbZzOngnGNmQW
FvlAqC9Jhf+3ZXg6Q75sBjhrBl2EqzijzcQLGDDFHtZqu2qMeOLBjMxVHwUq
98GtAJJyI1HPonef0rOY2f9yzjdFvXRhiYwYkQEinnw6NXSKltX4ZCjPQsIT
tsH8o7gaXOTj9fecYhNQgN3FXd0W1fz+76wuPzbmrzj/rKQPT3QMBRGu8Aj/
7Y2NCAFMaTkyu3le3TfzhLa0mXG46/pClDbNlQNWJtH8RsMOnULRRQatcRYw
CieuQm1Y7HQEJaoRrfSNRWqkONl1tvBymNz1PMaki8PjiwNtEF1rcZ3xqu6T
gB3Udzl3D9Y4Mw3QgqodPEVMr5dB3PpMx750zHlpyJ55/Ov376T0GqFWG1/L
MyqNeSfKTUweoZ+Q3xY7sYCyyZKc0VA/O+ibTWHfZHU+YpmPWRz1djsvtDx9
U/e8nyTXD/KYQt+vzTiLCnZ3dq6xHnCjHPHXGPxFyMf+iJsYnDj3TIy2qgwC
elOC/oHkBglhmDcMJBrtEjbcBEOU0YncCSVzcGvlOlXiHmL2989YkMQRx8R4
NZbDq7Dc/JWCBnlrmgGKEZKploIrMLCsMnBhu92vuQJFrTTEn51F1ajBcZtG
Zyf2/gObWDu0Q39kXm8QtdZkLa0hjslHF8cGx986t4dH1lpjU6lbqsthxfd0
x4ZOGCkw85GyzW//nCzHp7MvIgKhUw6+ir7MCx7dJsgnJVB2dUWt7I+PRoFO
+bjl3lCGMOLTRdNW7XeGztbDacFw+UKfpb48d+P1h97gsUuYgJfaqTBYKpIK
UEptwkNINKb8y0UOZF/IADZtzJwFQ0+sJ0O5JtUrN22HDwgzjjX0NwonL/ny
YVTZQREDewgllbvZsW5+7g3sdC4dtwUcLjORq9AuaNEPn2hbqH3CYdAmBQus
OoC9A8Tx9J8mhs5n3dpBxsyIoWVJFkp6rC6QdBqnmRCSNY2ts4px5sL05vxI
2lPBB6/dNqeyIDHPDm3NiSNWWFIIt4ZT2ZSDFIkp+iNGH2LC2kluRyRmAKqx
v5ka1VxRH0MHUtWw9IqgaktA6ZPNQwju7uh8BBd50o9LtO4DgytsjouhSCMC
E+vbVzLD4Lf5O58NBsQOmzVlDAz1rlF1+rEuQMfiv+i8Vr35KwkpJ8blkKlQ
XrKeWo7JBsjYHCC4DmHNP98lkYi3LU4zaiMvkRYMYkJhJsQcd0aoXT9FZ8as
3yKXdVzc9cFgetGRz+9fHKvXydXg3oTsGMm8B5ucEo4jRIKV+fp5Kcfuxm1Q
OwiwW/+2mm8m1R4hl49aWhmQAab5jUKcuc3Pp7QewBjQkW9sSz+WN39HRY3B
UlY0wCvl2/jk2YnQc8cfB0wW8wPHiawFh4hCCqihwk0PExMLJGqZKakjW6wY
/2CtPWb63mf/d+jjYc46rNGcYD/i/ndWJtCQjedm3834DOxgTdd0IWfSh+Ao
yHABZ385HOYgmdGmkBd3r8bvh5MEInhMb2J6tKGMhSiW1aDVduwFB9W+sihu
PxXr+IzYHR6HUlkHTnD5k0cLyonT8p6PTOpcNS5Px8QAK6sIzBPBGubNpJ5C
zHTGjEilL7Y7jx47L1yExrieUHbm6/mo3CB7UqgtpwrKsbkBH52oD+KLB1Ok
e1+XG1twrQl82lBnJ3K0mokg1r+G0nKDShKOzXF6E+vn9OmUAmELqe+GJ9qm
RXaPiXMKh5JOXmeqQdm7UneBWRvqMQodLsZnjjyKXzu17PcWdhFbSGeD+7UC
a/GYYZDGy2NZNQaKteMCj0VrDfWdDd61FEMWKh0ZisJhLzCbfniu3DZJizi3
r6svbdGS4G9xwU4S3/AWv0/vm4mGuZBiXi9ah1wCvHsqq8eL2Z3PxZ+Er0fj
Rd0B6F+ICVECEpKcbPdh8UYn5EemcZj4wEBdZlC07NnaP0b6Pq4x8UEtRVki
nQZO75W0lgYlPMu1xIXoXtdpGC6sX/nTEJrePsWiLcOpCpc5UoJVAesiulCX
0/ZEWRzgtto3UMuACWBGVDh1Zd9DfQc6ihmm7xCT5mCOhL+S5bxHIjxJ9T6A
GHIty7oW65T0efJCZzV2t66bPhOvHPeC7UZhBhK8Beden39vqvGLwRA5t3ol
Cuzz8jsmJ4x88mVYnKLdPYFr7aR3fwAj0pdGfwE6hzDZ0+aWId6tnb5gPpe7
NEJl7XrZm3lwMyM4X+46eooXwC6agRpfeEv/szc1/NPphVJ5uBFgK0GmhX2J
Fbe2WtbWK25SOK/bxiUUAUzlEIw6jQR08XCV8/4U72TmiR8uuLC2qRz4cj9H
6BBNeGxt/5zDYqR64Ii7BP3Qa4N7JRStYfkSzc91hSn/rAuGqY6vWi63C9NJ
M4RzYTtV596nboIq6hO14hw04g7QY6JYFhWEYFkm5RbegBcQ+zJC9iQWfyAK
IG1TLpVs/dJ/nqZNSVguScSsjWQHsQCeI6cw0Dk5XlssZAlUm9xLE5qO/XlS
P2g0QMdzUT524fMRDnNQx2ixtqtl1z/Oi1uNGOwkkO+KkGENaIy8S4VPIZYx
ad6teO5Ngoe7T2GXcxQLJO57IaADoUrXFa0WKx+3xZ5P5a2jdxqDxnKeLRZn
4DwPlUPTo0fygoMdC96+6Wb9ajYZNpPXrV9b6MzBFYMYTQOGj2dE5OLYrA9l
ApXBCo3WKRMNFhOaz4KUoG+7m/aJ8kt4mmghZajRcYMj13BJPlcFKe4QzuHj
rcjnQFLF6np0enyiJGAuCu5BNmVPJlO8mwa+g+GlMiQCim7ie7GivXcVjS+m
ophzND+J2oDa08nW/QqmM3vh9uvFw3/EuBMoojkhCEOwawhyKNbccIW8hJ/8
muN0z/Ly9pL0R36KCkfQc1Mh+6+g6p1Bn6KHshHYpv19HIGEc61asOPpcsIy
xMEGG2Go1aZL6jOWDjt4HmK9yuXli3T3HkM+Fv6oTNJ0A+tQr9+TvOq9hjPT
Wv8PYfed8s8tGAVJV8OWE80154t/VZRWsHe1AYuEkr+D7uKG2lR843YmZNby
swn8hdBWIzrQCrLqIz4znE9KwzZc3P62sKBeEohhX4QXDQmpAoxnksbxG5Do
MkQ8n9TyFkIA8NY4jxjj/sf6qwNyOk7UKY+/b/jUp1CYvreHDf2TK/9X+IZD
jW6SDUtcVzc4AcbNf23dCMoBWxQj3ZuKf/nCbj811wJepP3fsCu1ofSGPKQt
aDvvSCxuYIiShUWQyD/Qzg9sFFci9dHFQ5TUG7r5a0bJ6uBKiE6rQt/GCZ5t
u0/clexwWPsSdHLMFzndDw2IommYKmApWE17HPRUHt1J9YJanv3OWfvK0p/k
0IiXVTskXmMbztBknOj27IzzleQXkJZCGuY4mMFX7VRgGAiUKXvumccBqy1w
d25E8zE0AszD4BSBZ2tlTsPIC+Vy1RN2y/l17gM0BDwVihNRdCnu91kvJ9M0
RWtHIPRYpFEEMqvtdr4KJGC8Ux4B/5/sXzd/nE2J+O7X4UC0aiiIZe9kF9MK
u3cWKBNDRCEsE1qjXPsAPLbEQ1t9uLp6Cydi5qFU2yvE+BB/BMeHn/6h0YGc
AVMmQGnPAZe1kDy1DcJs3tD4QIbgjcK8uzrhRkRTXK/l2x5GgVn3zYhme9nn
S6sgOD27Me9KTYb1gi5vSiqpHFHicFXD8I/mBkoFcjqr6jydthNsivVIKLOE
FjtIYYVr38hjsHhLQ9Kx7jNBINDeIA0n9wD6fSCwZo5JO8V+8IRmqI79p+ek
oO2prMjBuEW+Kx39pYg5XtdbJgD9PodirHzuPAlXGJL0bAWWgg/jqIbQo7Ld
92CGfgbYpUq8BPky1zPhG+JDPNOFPPf5UYeUyIPQsspX2lfvFdvQ1Pc86O46
CbDn4Oc1egv09g+mNE7OUppHBXCEAlg6hSfxsEC394pDPIxvmTAZl6UE4+Tb
0Ty8SCzFQbu7+scsbnNELAhkL5AlGX1QVUo+s34iwD+f3xSpdRsW++H02gun
xCBgaFrJCvNL0NyBkEj60gIxoovMi0/5NGfuZjaM2kdK22hI45L2EMV3htx+
/LCRHAlYt5N+/FOBSzpArmIiX3oC7GpJHP976cIki5HV7DO4fkc9ostJJsNT
QbxYHWNmX+/3nWQqyYoMHEgcoV44O9TpH83Zz46K2L2bTYhQQnNVe9GN6p7u
Ve+N/za/Qra4sTpza6neYIaxvRiwyeRWJcY0nkQlGwTP+TfDi2qQH9c8Cr0W
SHODOakzMc6/j09OESy4dZmwaQ8Ue9QVlOXs+9zgBbJb7rEy3WsQIUsvN7Xk
vaqOuiCKmums5SsYjlxJY6GQUdKXkMSuVgfQUaSpo4QfBeJK9claSeH9QuTs
3D/Wo1nQAdP/vnKukX6rKy0Qqr+JHDViZR2PBZ1FJN+MQYaTOXI+a345zSSq
l4R5D0B3JPW5slqzQj/CBIptqGw+vDFSauUqkPBSBnFQmEvMSETUN+80vPXN
9s4jm917t5upodd0BZlv6QIhO7ndshJ81cDESEnlPW1mziCJ4Qdy1BB+cRtl
6yWPzi1Tue/qnk2Di5HPgpiLDLS8SrtPx1tWBHeb4POYoPsO7K9b8eQwb43l
MBK1S8RVIX9ieAAGhfttVIWf+ElB2nZOUlh6pLXGbUD+58I1Pc8SnaxGJxtQ
xadCwvnEPwLiXFYSE4b0sqrrwgwd/TcsSUv6LaWFKO3z8fN0HltPs59g6UQr
jPfSjL4rqIJnuzZhRYYYZnogvjFGhaCAb7viEB50WANLM0FcA/cZ1ygghCw6
pRD9QjBBSWlq921ileP+8CVWn5IiedD+oxH0s0g/P7UXX8g8JyaUjnILK5Us
GwN8OTfhQ+cjXmqCRTsZxcKiNGo6alH1tDaFh4nRaXY1FhIgTgBfZjkiVuL/
YXLheo0bHruFGwji1TxNr8Bjm4Jj2uBOn8INx5xHZ1Qk3zUZRqu+5Faj4S4L
XlFW+08P05ABtGBow/2qO/tGMbgb9sjqVJf4WLuyevsRvbXRrbl9O+iHR4rp
f9xpHzt78W08xUw2ey5RxVXfahJX93BuM+RYLcyo3lR6Ts0XbTabuQDVDiJX
ey9MNlUYlHlLOQLQA2bjWagmpsLbY8Y/Qvq76qq7GhUYnxkWkLwt4g0zgiKL
n0m1JrHmPXjDdw5pInVoQhAdKsSnajtnb6oEVHYycm1FPbVSn6hwR2Ppz9u0
NCPG+Ccu4lumjp9liDTJAQ3PdGdmuzKv/G7UKxURXCIRvOm8t1Rh+imVBv/6
UyqzvcZ+Ym38F2/MkeLS75hrQietg6cXLMpd7WdGHfs5nsFr6RJqyE15+KQO
xiE/KZ06hTtRsyblHBE41Tg/6zmD8dCVB46b4i9e0ZAmJGZdShLPQDXa1DfT
VrOzwTmnlclWntquCSMNGTP6DU7HcUseXnOD5C44k/SdnFLckRCwt86oPVlt
IWjXEy36+4sHiQ7RYjULlS+RUM5vOnVfEYixLyJJm7ohq16/XUXemo/DZPwQ
MdT6SNcoNj9JL0TULb7Qj4FYqfb49vEI90kVIj4a0DHqqs0S1W3wzbwc5sKE
t9i0yj19MFGR/r6TT7g52TVLEL0DIr3MRizKIr36k5mFgJObCK9DQCxVuzY0
wH87kSEz46q7vmjddH/CjUw9ONotuwdQS9zaJtaZPkPtICAJGy0idrGr6Xlx
preppDqotMQheIulqu6cbClveIz99RQ4ekteczPwGcZ8zOCAVJ1gNNkgbnIL
fHhRbNGqq+sdT0oYX+aPCREo1qmlr3pvYVT02DuP52c7eNC1eg4wu3/X0l8a
QSa1IBxopE/t6D+xDP3FAXPfS5n4ue+SfEpOm19z0jgN/YEGBbrt8aNQeEJi
+WeWUgYa6hHojgw6Yolt+REjl6ZBfJbphJqMrQJYD8F8pUKqyVveXKTDw1vw
V9ZBh72gDCLaBKSVCxHGwKB2ke+uoc4plsgkqSoNA5SGorRll6ryj+v1r8R9
aKGCGWxyG/gcLlTOeaMO9+jO8WJ4CFP5zRELuqCsTQVYSPgkYLkYIemirL4f
r9GkER9Tx8Zx5aBMBKUc+gp/sOE5JBL8YyONCMC3klQqjXcntHW4ZaJMLfuc
JnCkJP9zM6Bil+bu87S5bhmqRdNhTt9wmpZ9tuWKJkmAP93ieLYRbZewkzPD
7tiQ2XmIyx7sZ9VyYwlTBtbwrv2PzzCW5CJfOwVQANVTHwWRvbVNhX0DiU4W
IcKC/P3r9kDH6H2PDaFfuDiXx+Ws3yWDlZ4RdFb50dv6TMYbPT5xi6thtK+8
wjF4GVvu9KwELJvx49AOFcx6cUAo+9Mlqdw8a+odnOHcsNxQSDl6w6K59A7i
SLAG/8WKTGX8Gxxx+8GEJDpMC/QYoGHEGaMvZv7uG1J8iVvy3JpeS3DqwBnW
3Tp+kkugamA4qs75QONWYSOwQaQTIcio1tZClmIiQhhLJbVGCsNQueXr2ddD
COSep7N+20krDBtkobpKYakw1ZXaIQ4fd7vJo+h4BNOhpwHonuSfLzw/Q5Lc
4f4pNGgpH+git6Bo9wXY4lvzLzwua430MIQbu1+oktDWNw/1P/Vr9KPx8rHC
Oy4JhLMIr75pXtqA4/Fl1wN9z0jEXFAkPQFyoGYkf9ifw3yknKYrO+ekVdZ2
/sC8vlco2r7recovGXCGZifzZ4oVE+7rajQWN9Z1qQDjCzvDNu9NN2bxYAwv
X+I9iRqGLJ9JJ8xWesdb+JsHHNwrXBimO8Bx5OmoBYJ/JWDO8eZzE8uq/zy2
t59/zNqy7Lj55MPNm8Fr7z+8sLG60U0ZchTwmW2HhhgPzzDEkwW13a0b5voh
6dYYv5IiuyYRcRu+kOUol/cd01AkNZQ+48E+m9HJDGI0QTTdAUikl+/MtEi4
Ivqv8Rj9w0ZX3wVA8Anc63tnYb2+SydkE2Q2gN4p22Pdw41krJ1QcAMg9DZo
VLtMlGvSnTogsXLkMVzZQkF2M0xwbiB4g7z3tbX8biaPnuEQBUiDYcOB0wDM
1Z0Y85UOT0Zw4QWT3wyfw6rlDeUzY2pmsF6JY9XFt64qEyUZ/7g1keJayvbd
K4oahVybnlxMhF2hwdSoNulhZooRHi3G2W1mLN361Cam8QBhJkL7eGm2ZWUL
Z0doYlacuYcfLDo7fzaDkGxAZa+rsTdnO7JPQ5Va0eVaBSF8GZfETZlOc+a7
rNz+SZrs2nsa2RKyR/URYiw8uQu35uTZWfeJcpb2Qb+bGOv3aJLQjwAJ/O6n
rSMxrvcnUIHDencVMPnUe7opqTqI+QXD5yKBWsCSjqE+bY1hjH7YKDsXGyJR
sjfw7KYFoaUZhG8xsFsfYVcVwc0ZrWvRLUHcZcEG0/lNVHNcR6inox++pgkm
q+JgtetZvBZX4pREZ8YjoRq5bjEYY8S7TRGjrw8ltyLAazeNnZrlyoFzJojo
2ZqYU8OEFsqnTH1OFRM4TzAfx5klbDwXdzSMm5DfMoDOwJJ2COauQtjopVo2
regRE9Dvf9BfvQtOCJy5TGKpFVqr5WmzGypKwATwW1DWP0mXioGAZgCANwSJ
sO92MWGTWaRxMiyzKz2PzFIy9urqpDmnl56aGSV3UaIC1sCP7brcKxBd24Kv
4OiYZ5oUgvn5wLGmGOMaG1KYIPtsmXwSBxWKaVguNEEro+F1M5SZYQs8NoHo
hv9h9kkqSVhwRye6x+Fz2n6p1XGXlsG/IaqTbrpNxHCW1dvtdvG8dm9202uc
dCkhiHsg9ep8e57uLhzZeNL1IRd2q9wtV5RlESW+mDvUBkadXwmP1PBoAu58
eFfu8aPn/e3sAdZ6H1nuo5RtF4kuvIwt1iAkG91Me6UtByqkg1qRPKL/J7Uh
bG6pofiXdiuBFFh9qvrztNKKbYgvnLpFsAuD/bgicKcf+5vAK2mV+Olqs71i
Fr88dvcuUWBo4NhZdfSZ8VVniFsUsAAachkgJaQhwu5JucR9f/pH1Kxx6cua
jcxUbsGhruHBdheuIj3eRHn/vfZwT8Y7jQMjzxcv/yz7B2G6AqOQ7ddYHr/1
/PbIA9G1urWn7o2aijbvyBaYGnqnLeZSFJEjNUkQM5GDdtZgsGMjYUzAUw2v
/BMINlqvvAIngncZQ5UrIIHfoia89yZ8J9PI1dodosixNtWNUdW4s1gtzjAf
OPQWdqvrjVIpIEMeXHxHzsLYvXUnT8K/hFUcJuHTfrY5gsM6v7rZgsfMzHlb
ZhnBBLqA1SmQI6z/qwAChDmUICOoo+2Cc91TCiZ532vS5KFajM4wbxGPuS0l
iD6ayjos3GaYWZ8qgZkMUMmhiFgZrgwV3AbVjYBd1fYHFEgWNIzbF7g9bxa4
LCLVJGSw91w7px0kl99md6wm9/ghVVureuTCSatDx/0WNl0BsQAxshqyuGoQ
uP35xzBSnaioNRqdzBsil7uHPVmWLZ8ovQC8ylXXUpCf6jbLD12NrjKR6cPt
GA7N+4F8/TpQId+8TzQCvexE7IGdz/FciVYrHZkjGFK8+zP3PZvDUrfNTBVq
WPxHBkEUl2aasCevkJTVttCiHZ6pl4rjAAwXf+uhighqH+wUNmc+fh+gs+jt
25Ss3QR/AxeDObiMOmqnMuQInqSwc+bnMOsy6paQz1We0z/PdS9sR/ZFnipY
mWz5C8wC2Mgq6bmoTsrPlnRNbSG2bjXOKudCYA7MMbOeHE0jHchfcUnzyqTP
YDnXVldWWz3zg7FLQcdofPWs98RrZprFJM2cfPqJYPV9YJAkBLDeFKuoTk8X
c+jRy4kDG4vhjZpxYsY/BKsefS9/RTLuzebzJMRbUA1kb0LLMy7jCfWHYfF3
UyDYVvakKUb/qtMiqBKVh9D1ZX5La9lWDTT7CZgwXxd8M5xKmoB7GDUuI66D
Func9g030phWzIvJomnRLdHMcdXNmwuY+2RVu412pS4i+AYSATxy5EYH7vTI
mBzumRgSjSe5YEmY/VN886HzmOzn6fFbfvvrYIx/2MoIPhwgr6CymxHgpt+x
j9cE33TM0934oCm5zX7FVxEkpNvcSbV7T30hfo/2qhAzJzGmx5yzaPyEmQXx
ucPQ3A5fdkhS/lK0379Txvlhb1MI8Svggwg9iIa7yj5CZmBCCDjaZYdYTsV1
O7wch9LwF5cf5YQGX7OSdtQLXfmPdUeFppn6bGJsNV7FBu/595xQscWpjdya
VN5+4d+fCenditwM2CsSyowTec4FGEhQmGjNiGmCO4ORWWEC9aQ+wCJxmbQb
J6dB9EqRhPTvnxvYvreUddoA/o1xeIzk8eiMc39JxL7y76F8b19MTOI1SDXX
liYKuXHHgxIym0As6eWOoiq0dzL0TuciLv2B5kgo65NGhTXb4HheNcWgDpB0
ZkMMFAWa4Ekb0gNViERii1XrlQXMks97akPSj54By9ybcAesa5IDST5ke1od
Q2gPUBOnYjFDmjxUjY90oL1oWIKPFzKLcLToo2ZyQDFTOJI9SgF1ICkbfOM1
v5iqKEPXHrg8/Bg/DdmcyDWArfTq/Y7GRjbaUJDZWbMt59AKV8agw/lJOQoQ
RC+PuRUdVkKsYYWoaqQgXxyrB87e6gSbZi62knsApprNyYSM4O6v3T6JtapD
lohhf42sMq6+HJ/Ah8IPpAfKjNsNM+x/zGnXlbQf0Hent4CTGCZyet1JS4An
Du/82SoV0EPkaej9fJ4hUqiKWGQvTE4I1vK3lry7XA1IisItOQJwaaf7H8Ze
SsxSPVM+kC3RNEy/s/cvhrq/ZTszJlKwVPO25HprMneNbCn/Ie+TqYLuaTIx
9leWCaUZMRedTrxF7pd0Ui5aJIFClldPV146EDQ59xN4i5dXsX2c3JxutmHa
3Epe9J8VkvxOH5ZIQJiwx+rVpGTtO5O1z9KVN45t/2r1/SnmJeM9nwr0eock
mHMcyfoNwiYNKApJc4iIsweE42V8OKTQMITHf17m1ry9eOZ6RLVkMXQo+SHS
sPXlDonEK5zE1/VaODidY93Xlhp1OxUTocCZskWCwEFbsxKRCEh48VrbGnUT
KgPBzLLX1dDS4gR1UPYJrMwPnnzpfm93YPWqLf9qZRW8LPftxLWZk0F7GyF3
9D+0CXHXHB5NGrJo1djbn6pIVwX9g/XtxAoquKw0M824y1RdfZVVtWVP8sgg
ncvpIo5ebzprb+UYkJV+8WIO2ZDmsrTlT7neeZmayHd/yjHxnHlQq++E5EH+
qeJD2/gFqqE4jGKZJQ+cLNhtcWupRKTX/OV42pCH/JkjQjxSttvGRHzaJ/72
gsKF9tkknzFBfgyogJ+flFiNF3CdkvcobGL6MVoQ7AcPDEBR9nGFtjtBpC7H
ZNJ+hl4mfyTsMhVwb2nbsulYA+0tOJS4JNihdJVtkCnw+psFruIwiMrkNdcD
fiQSLTX4Cttc2DW8QKspXvrO+gk/wBMKyu6bhTIB7kFnMGLTYAAWg0epmyCz
x9kQNWBijcarbNFknpEg7yaE53Sj3fYjfq7PH12tA1uloM3bPIpG1lJPO/50
QPEsphha9wA5UlRWgdsqnFoUFa77x4G9sx0x1OChUgpGtNJ3Vnzwt2XiyHRd
PWbxtOnNYv32KtySnYaoI6Ui6E4eZAZc2JmbxWdZLF1IVYj/JaTxonI5ShNw
GhZrWmxY8DH7w56rAHluCjdook0ll7+4/VeACqY34ASd98IUtJXwxoclmVxk
vPfcrRhYAZN15SB+3lGZNXKHWk/iwqleYgWQIAmm9r8HWxgv37HvxXUfMA8D
IVM4EuWUjD5tAU30Ow9QHp3mIRzseezIckTppAD91+8TuoMZUEGlmxMH1QXo
zODrMJ9S/KAu9a0XGCHzgldZ39tO6FLNSLEnsnxhX7Ezoq08wUYeBtCQSUtK
HO5tT4BTSxsANB2jIIL6JLOzmD0vhhipI1JMngzfMaSVOalI7D9qaezinYrs
NGOjI/l/gF9zPtS5I78UuwK/tEoiXxTkjgtyGw1lcfPMz2c8xAtZPTwVoTk6
aAs4c7BgLj+o7imjVEyfJBR9+haw0rZGjFxYM+0fbGdUYEiKLYHIqKnBboIh
8DYX8C3Wk53WnyZPHPve3Hfn/H+lAMgAaZKAEWrIpJ2HN0IDvC3nxEbtHjZK
gmdafdsU5aQYF/3Bl87J1LvfIUeOQ6SPbnCqqBWtQmUQ7jkgFV6y7SERIMFr
RC5JqfptDv1Xg4oP7qs9swC+hJN0tgJAYd4YNYPUksmglo86lixNRN6r+5oV
8s9c3q97p4LwWInWbIZUMPHNHBsiHKhyr4bEdAmYvSOcu8JjWSzla3hBajp2
yjwjC/vOXRtxhX0Py34SoYH5zsE/KGMpstVnEBm7DTP1Co/S7GSn7Bm2ZC81
qj1dEClRwXHw5ZUi8pIMPUBjTJf7Lv3Zh5xYzvz4D6wNzVbe5bwYAN13ZQHl
kuwXRbu1yJ1NLLZ6xoCGoWf7bU3E8DpbXnfe4UYTEpKP/IyXDTlucgFctAOo
xznnTBigHEypG+qSbEnBnHDrOapqKsHYCSDdqNdyoHpFhRgCTltyHGM71qAk
RyOcmZCp9PcHy/4Toi/4LdFZTv6wtzAJ/7tBKNeFo4AIL4HEZ256BTZr/Uwg
OCBRD/OpI4a1JQQliNEdbh1Ao/0pZEdFigIPgjRPiM+ykube9mqGfqD+9esZ
hOR8TfE7Db8r29qWS2nf4I1YypsPshHWjLebOPiPgQAXi/nP6/NKxnlg8lJU
PljH74NTtwyHLHOdL74qLMnIxIjWCsk019dygdIPiacl7T2iqOFVwWZ68CYb
axPhkK5J85EkqTjpyP942bQTi9Rfo0RKbIo7VrnMoVeviyjwyRoti7rDSRQ9
tKktc7sLruymyNOI8n9qS8wJtGYFajOq62IdysB12dvecJSXKEjW6XADVOqt
6mYRLTXmE00ZgAt8NADQTOQi15vZUO+N1fskQBarPiRDZpNGYxHJUF2ANwNf
1IDedKDI+S4gj3Sq7y7uqA62inyLri2/ZuUoybnHZSyCZ3lNOxpJZrVigewd
TbmQuDB9hxXOKcVB0dmsxbq5zMAI9fLUenQAP4gSPVXJPmESvMVzUZfuVxdg
BIFSecRAr0wIO1ZQbZ2pugHdqsDtYw2kuYWpCph3GFAd9AhYKDolJhwgumu/
En5faeyaK8uXUbuaEUvr4ZCj9TRKs3kVSReZ4O8kxO0mkuxq6LQAjRGQw9Vp
323Zxzg40O9ANvp3srtcn6LU9ihei8j5fW60idApz8st/KlKVlhXFqfs6VJ5
UrpqWSARcOxX5qtooCsEf34D/+O5yjyo0kSNu7bI7MDZ8OAffG0NVrqy82V1
pp+8nEHTU+NaN4KdEp/MR1/vZT/kcWdGUXj6l7KI0BFDTh6YR41c5O4SFR5c
b3U66O40OSQQi65qJoIfAtoay/A4+kLNS/FI/OjN6ZrVOFvipB/UUsrxvtY0
walnlaILvh4TdM1UzXyTQ0pXeAqgTSX/1TBPS7gabU1V4E4YtPKEPl+buam+
yLlHKvdSA+jcdQu6l3D3r7baNMvbDScaiBNxbz4q+apUnu5qtcGHZWLe9bOD
IqSeIh9E+9gcJlp378DB1mFkK2i3dqHtw//frJkQ6/2MEdp/Lj3Kqe6/jP5K
GX988/B6wuRqADrmCZNgcPNR694CxWZMRy7FbMtXR0JgWravEUpys6oCxJ0W
98XNN+htQpDn0g9nC7fj6dDhoh9JgWzI+Ig+3xmzstAd1zFQHcYyNKljh5dv
UzoxRd5eozckTU/ympu68Bi+yD9Y5mlRcaBIdPywiNP+BmwgIF9aSa8BcRqs
D5jPwWWhY6JbRMXG8tbratPM75hquoWI9zCrxvWlMbHTPhBNZu6PWUWFoMPW
2Tj5w19mbSjO2R+5xFRdhvhhRzAKt3UzEv1UAdNtmZTNuAkbuQIYMPrg5CGt
3CfnzU4sVbMb21P0nFXmegy0XW2l9Nc07WtQIjA2ShjLVEHpFC3upkXNnb4V
HE4vpKzAPeSknbU54XHtwR57bV1WUt/umZlpYPcM4cvE5l6QTVQU8aoqKoLA
JBzErrqAaqTIC15wfEtiM09GHeKMiIQ3p6QSWKstHquDnFs2Lmp7bhHT7bCX
tghldcOyczeu/AMKc5AkXAapDpHb41yc0ukeygIS0ae+zb4yn6NAiOl4w/8w
jAQgKAyfNulQwsr+a7JT0SIoB+s+cwedrJvL6gQpYO587nCyWWN2hwbpwc9W
3P+VU64E0HZYGjY9asMLEJ7qZzUvh40QRgwoDqZPc5xm2U5B2+R/cgqonyUd
mnsM1Yzed2KZF4jvAVPhUZZa0H2ehAvGiQq6Oz0p1hqrwspiXWeuT2MdoLow
4AvPdqRmeTDO5IjW5D6Cp4OMHJBNXTOlN9XSOlf9rFaZ6MBwwFWtVbp5lOc3
5IFPlO7DjJvrIoG8WhGHJJ3zRbTfkz0EegyCVZbsP/ywKmma4t66gE64AxHo
1eauLHTVUhzqBosNSUo5vmpY/D9VtRV1RFCmWa08Hfm38w5Yd8TBMYMSCMUE
xyKeNgyc5n7C+QJqhgPJP/IQQK1d1eXITT/Rb1dcZU4sXLSvAFYYORRtR7Ty
hvRZ/fo8lI8PE1GdQ6GXTxsNcxecZsTheo0M0Jm0v5tLwLIQvli1PrmHhXVe
cFElAGI5QrcEVeoMhWd2t9mnJzpscxuI93FVlqm6F+/i6Bbq1VpCfeiFH6jV
b1Br3M3mx+yTLCYnyRS7WG3a5CBNnBd4mbFTHSoWGsA3k2NoP/rK5i9RQF6a
AUpUr+syhBGQLsAfd4VKAg28GfzQhgTCwsG4e4H+oWYGWcLrf1x+jNYN9U4G
wdldAoeIBk0QNWwskracfvVkcX/FIWa3xL0xQQwelyensBP8FSZE6Q6uZl0/
a9pZxXrv1w1Rv1WlfXoK2VF+R3rkZ3jJ+cE2b8QHthXWLJbxs6MIMyKlrnf/
kRf+AxVVPKLd/Al4plWAxt57HUQ5r77lDyyiBxzZtXVMAbVM/p/ZKwG3lovX
PL8EWdlFMWppty9Wg8VBvj0vAv/R+fflNqJjh1yuHtOyMu7QehKE9eRPxUYi
4QnXIegnNEtooyPFdzyH4kN7MtVj5AbSdAMWRyQx3k0mo3wf/Xv4ur9XLXHF
rove4/Dlpe3a8UoTGyTSfeeqKmecwbkgi30c0G3XC9yzla0qmB1qmAJUN0D4
lkfgAU5+6YvJmcwTy30Qd09cu06oFwc9JQQzRJiwJlvz8rb2lZbyHwZKlZdS
tm0ccV9j7jhhdQTDxkahYcBwPCFHJ/Sqk8vumYrtrHM8MMrlvdo2AZYrBaqO
h9rQpI/rCYpJ9cDA1uBUnnHFLMm4iMwojn80i2aU/xuc+OP7BffRNB15n1uG
nZbTcxQPi4bKYHI8YoczpMVBrM+oOghhk8b0lsUfXTRPcyAQyBvvguLhyX1f
SZFqx3/8vTM8ck6KJfWd46RWr+PF7rdBV33ZPiGbv4Um7HFjVeyXSJWAwhR3
MWiXpUz1FmGTjboi/BMXMqQ6V86SgD3JoHl9mh0mCX0m2U0+iu2UHSVzm9x7
F0C4iKahGpp/GuTxDlAM58REg4A6Svh4mQlV3eQP2lSSVda7vNcNZIF3DZsy
DIkK2s4Iw7Ut8j14+bEs9Xy1XWnc7xujYHAA+MuL0SXaRL6D132qymUuN4Nl
W3wrJhD6h1V2belaFALqZiHFuwHEssS2W1sANiQvGZF6zmYd1iDUvmQ4dSIM
sey2jBMlw8IdRJp679P/tgFwAiVb/VVB/mAC0EspfN8m926YgB+Sw9lMqsRh
u+IS+hbX3uNUcnmpD+RsRFRFrVF+Tw92gFwpTBYARl9OEiwqSAPJmmv5YLd8
3E6dFBPvQKKfBB7bNLjLwT6cBKVmrGQpNFG52ipNs9IiNoBSV8qdlANQ2M/y
p7w0urPSiysA9/7EFpWBg2DuKN+fNECQpauKIXQ+8maDvFfAiXK8FnfCJ0ct
toNSFbKXB6UU9I9e2dwfY9Gwcba+9fSGOL/Fg2P0sK5QA/Tt+QYjYZqqWKAm
O1ygR6cMmI/Aheajg0inD39VPAsBWvve6BGuV1+YBHD7LrDk2TolnK0A80sc
r6vLAaLYdivUC/u/hSPWsMQov4P1JvMxzjEPhL1PK4TCZVD83XvcElvylyMi
YFqQ+VLzFA2w8jb7ebuyhq1Umo/iD4c/s7PXnFteAjGeqo1CTjXL5Rq3fXyN
ec2o1LOYCPJFGOryPcTeYmmAZmXAjRnqDnzsEC5WXac9efAg9FDFK6KUl3ZG
b5bQzRPk9QDCFlF6dRbhS4Ov1Kh2Mj2ZZjXzpPM0ApBvabQaUrY0SOH9uxmU
S0/Gk4Rrw5Qfa50uSObEGIXq26psRkHglN+VIRi2tLckWb4kedNXzI+Xr5IP
nHJJveegEAZKMgIkyxMa1WNN8Gyn2TSQf98FyA58gsKRmR8VuTUxLfLauqjz
zyn0r0f8JMgLXfNAlnU9t6gX3X3gHY9uiBchLj7xfJiy+xhYyHxTOWbWOKT3
CrHKpTHrhj43fl31LLOPcNxOsGSpxR4CFQ2yzBZmkX+dvAVJu3pck7KS9GqH
lIiQiU3frIIZAuUsRVSL0yQPW4P+iGfYk0/jGabQlCzOTpw1jnbEpWNaKRPC
8wxq9syfKDK3CYkzlZwvqQIQFNFollL4bMWItf6lDxKATbwP7rzOVW9JlgB/
8ZfncogfF0MDQTAoVKAOqZO/kSwxKi7KyjQchzTz1YW9I8JO2bAFb5OEbhDR
MzWRcf5kFu4vSxAZWpDl1FyxPTiZC+AGARB5UxoI1z7vUxUq5oQDMpDkBIq8
/TCovYBloD/biVoGJ/RW1BBR31fz2KUK02zo2t9J2kPCrLT4/9eVIccbJnpt
4yvQH3RyABD+RBh1Wm2YzwJhh5xp1ewgW/DK3XpkxTAkjotyahYjcWgPiLKa
A6tKPL01HNA+BB8PnMJBepKcxCLaCfryEKiyoVobwJCzmNxp4M5hHGpPEYJU
HRZUIzl8otl2Zt6CkkcUQ9LgTMuG9eT50bbUlU9gZcknuqGZu4TYtCJ3hsQQ
v9oWf1eKJkQnjp+jtZtlMfAPLEPRq2FxZUa23Cq5XyYjNZROEJZqr5ykdp6o
n3cprjuacPP0+pLo6J/h4eB5VC52RFs7QbomFcL54GijhiO0Iuv4U1Jt6oqY
FOhH5tnzrXSw24CCZe4uu3FmltmPgCG420QIi4TEw/3IUi1zR5taM/tR2s/6
GvU0u2/7QSWoRXWPxQ96sFwzzhyeYHHxbYM+p/eU77SFDrTQivBNyduvfCis
2H4eaIQFaUiAhYLxncvp0QCacCN1u5ZxQVDCzmbe8nwK9iYcguGmuC9VXJ7u
VP5JMaU97eGzlKuT+naTwsBSUwi6qf5YC4P54jQtF5mm8Y4zhsEeYVwBaQxO
gx4MUHAJ9x3BGOiMCbLkx92Aq3pgS+OG0D+/GF1LSiYPIBhAJHOQbYkKL45q
djg1zctjCd//oMseX/Ok+FwTH3GLpyykso37wqMCyHc2kpC9FUllZ0P92ePJ
wNwyBp31Bi6IhVYruwth697jJnaSvqkWereg0C1/M9NM07OPXbcIf8ss2WRd
jZsBzfj6XQxTEAYsp9bxsCUlmL2oK/TMLTgJEXkfayqowuT7DEGNx2Gjp/f5
kV4NpDrXuGbBTOYm656B1/W7j6lWwzrwhknMqXlB9J8XAjkNZjvdbfeQD8nO
F23ECrVzMssDw3ms3FRCUsINU9RUzF0+ajaHRcDtYKWnEm6Qd/tQn72tPxcs
dX9ymx7Za9rGuy+ustSm4FtB0noSomi2ZgGhj1c7vrZ1IxFQX4HWDKuksvBJ
VwcFFpeu/87Hq4Jzkz9KfWptNQJG2WB9v7FZQEIY1xXKf4w1qK665bZ4YMKV
PUtAJ+mV6NbdnTF2AQSXdVAV+JyleVjcCTzUi3jpiDGnZKwkpuWUox9vx8LB
pUIDmPBfVE6VYps6qqIs4QGG0Ar1cU3SjGgSJ8ESV3Bh9fumHSg9j5P5RMAL
6wZDQUpf+UZZjMK5XpVM0i3E8CWhkpfMbIU5WTlJ4l5d3u3J3yJTV5ZYYQjS
fbZpPEUEiNXOghT67uTxdmrJ6whonSWSkxgzbzxzwVgD9w8SsasT+vqiV1TX
CKJw+ZM/Jt39AinMXZQ4qNq0QdzmANKRURc78suVJFIQo+sVPimlE/+DgMFl
2/at4yrqxF8WhEip/RiGuhK5rPUt8Y69Cs7q/4AYpgzW3xtLEowfEIKVVm+l
8ZUdOf4rq1uWY04xLi6bekJ/uoPI9qKca0AU4fdypQH1SYTTNNWiOW73wgCg
PApPRblbs+xN77Mzj7cAC0XHy72yTcwEQgsOJzAMDK9agtk3yWrQdvzQoKtC
8FiNeczkBlvJu74ZEPCTBkNmiSsa3azGLa+U1jEVVgxOqooCVj0iTOcENmoL
JDCWR7+1TvWviNZIBzqTjErLecvnf6KIWDqH0oxTER8hREMExT/T0i4MifSd
xja910K4wqijD8CWYwNAFxIg6J6sz6kp25dBQ9RhM1hgULvYajwrhVhV9bzs
lUYEdfBjExKZ454yBomdOeaiQGPCjV+kvrD/qsa3bMsowmSG09nG0VB4x05d
cWxqjpdBxogpz4B9jPzO7PuFidkrP/iIvHCXNWlkreHKkAfxC0mXZriflFN0
m6p2HUtqq1HaZbK5Q3wWHlJgMToUXY8mEJYJIg+2TdNukfCNuBqWsScAGtSx
Nx54M497PzxxwmZFGiMnhR2f8LzgbGrdXgtkVULvU/0YCru2+h+rzWpi6xiY
F8KgZFXvClN+DETFLovZ8yLN10pdgJeT4ZIwyeGmSYZjTsHq14qmw5xUXWBD
g2P83Xp/z0zJoQsxGN4NEV6WsJe6cpsvf0P8ioTMougqW3PBx9mThDwLXo+W
wUBbaWQ6QiFeXIysjKt1Fd5dVA4S+9zIpN1fYH9RvPyPjULxy0jI9bDElq8C
2Uf3g6WfgQBQwGsmUikc0C9V3zbKX1gsUhcIXx29ouFNC6F2xJugHJG3bsYh
S2mMSTYGpguiZrmjQ6HjHIytvr/UJNzTkji5Y8vAFm1HjndPEOIRcU5hy8ji
aV+diHzfvGGwl1Y4BxGPH26sqHs0FwHeYeVucoqEXcTcKFrptBI6W/x618c0
epN0KyuOzZk01dknlHidSoxXGFhqH2I6kx+pGp2MiYORJcnj9PnXEgmTsJVE
N/1k4nSELCSKFAsSn03Km71R57xibjV9r+Ydi/jiRfFrAWg1wA3CLmJpkkNW
udIVeqZ8yIahLH70AH9dTovJ60fs9oKVbNUescdy5FA7hE4k0g21iUz7hqr/
XESByy9EfjBpj5kVEL3VtUOpgqMr0ccLKE1speRY/KQwM3fXCWaIVvCX800k
oWE/LfID0G8GoRLluMivXzWu1UeR8JgZSBWMaCnygFPsrjWAfP9OmX4n+03W
IUNN+Wvjq4smwjkHpYCAGmXrPxMK7QupqzgITbmnuRuynrAvj76BEGcEBNmS
I8Wl5vqaIicugPC+wDjptzbaEsXjhn0pEKxhbA3rl5b4j3/9aJBBFtZiZQiK
5RaN2bR8YbfYotNdBulJUl4B8Yass5B5SChIyyKDdmQbijcyOtgMVHosptR2
EOLMvoWHv/XhmUIYijdE+KMYsd7OiqN2qjIYojnZfz3ZvVjbaTzKOpbGEiR3
9H/f+XLmVN3dM9/3Q4HRDDHimxPu6RWdBRS9OgjZS9yDBN4eVGDNYzHiakAq
gnIVZs1ifQwWmsv1YXnFYAw7latfK6O48Y8HjJy+uaAW3d743gmTZmLLyQ85
eXQMwkLcVbXzANYwqUZ+Ben1RpFRJUW1K/MeucKKRpweedl4FnYL1xkUpQKZ
Yc5PkhBnMwIauBma+slSWM+UEQCmpbLfT1Svn4OVtG/cNeWL6Q1nx+IpTm0C
Z0+vqMKOekcXPHbyUfkR62jWCSJFvZZjjHEj5rp8cG0g+CSf+pajqe/UbDKh
b3hkREwlaf++wfOlxuV83OCamemx6Ht8T+cPx/xP1cl05T7r58mwPsj/I7R3
Biotk7aeaMvXjYjsUImyxsM3JR1nkquhna0k2qWAUw7NR6ixAruAiePwohDf
EqQma1PSKxba35aJkQEOPlryVEMYw8WK+vKZO2TBPpA0oxDCkufGwPSteazW
ViWrreRSUtNZ04VOQsnZ4OBjtqFszU1PHmuHaPNuwI0+cL/LTN2tkq8Rjwsg
Y2MBVXIAWAjY726z8DlnORS4ZpXbWG7BbjnoUQ9sy/PF4pd/48N2z7Ybmj3I
xRAw16bKVv6Ktsh8qYcAqF4XFqAG7M7wMz/txGV3J5ZLEBDWmPG15WHtY/z7
12x3/wA+OSZfIbO1WPje1zt/iAXvJb0dwYkWuLg5cQ8qqw7MZgJwpjkUjaeu
/16kXb+X1/GUyFbLpzL6Uk3HRBdWm2kvRUpypzJtx1Rk1gi+fO61pthbX0Ko
qnCfxg2Tn8evCwmvqsX3rXJP4gPKrLJ8sPAooCLkTW5vOPQuI6qMnftmV7ZE
MUISjZJ2WlZ7cUGUdMCh9RrIaw/jVcGu97buhxmicB9H/qHp0r/cKYYwdSEe
KdK0sBHq/Xb27Zc4s0HqdzWvas9oKiyOdKIukvVOXPT+Vl4xVwmaFG0h6Q9u
Y+ypvwhHI1YmcBtNyuqp/H1H5l6zqaxSEj3+lDBgRq/nAETaxOXSnhqd3r7S
Ws4+l5ghofv4JkEIHYxTpPgGudIGNFCA2aCeKDoCdWce1uo1xPljVckmPU+n
vIJOMzDbmV0dTq99f0CRd2cHSDddz8ATQEQA4F9sgZfSnRm97DWw/FSn5w8M
r/uy1O/0nFX+pWfXtV/5EtyxQ177qlmcg2PHDuDRpYKU9DUxp/dg+r2i6yrO
wYjBxoKdtoaw043L5RLN3dCjep7NkQCYwmBI/QFBypyfydiWBhhTZpiUHunY
wtLWuX5CzxduLdYnomOJ0nnxC8V5iyMaMbQYy9tslqgXkSauJmmyUSJ/vKSs
0JEzcs5eRGjJaWFvQc0IMjFguBcAM71gWAdIHFBzMp+W1905M80M8NXPVPoP
PJaPmfKpeLSXontFGYyayXmScqpcR0H5+4EnwTjYVkvampHVlXI4+nhmBhB9
oKZ5Ywb/LKhUjI7Q2chKEfKedDszuPaSNYO5y9sF/6hbci7FxvW3LdsMUPMv
a+LViRhiKsv5ydZnvFk8EAzD2QLKvyO6a/5K4DIhDT9O7mD/HMhrGs8Gt92p
F3CsdFuAL/tsNSsgs/+9t9Ap2RSYGNozQG3iukcww9Hwm1IpMTqsm+gUo9LA
1bDhzMTVFaLoDdufXEa1iQga+iPnCRUgm14bqzf/d2qXRe6SaF+DrVCkplpG
BPJcJZ/k+lpGoyiahfbEOX4ZIvN2t4InUCoIsCzq9dkMqtsc9l+rYuOkaz0s
dufEG1Ru9po1mnjgkky+D3aNhhvGrh1YjIN2ohz/lDO+XdztxpY/AaFTjDuj
lJSVwSqoYxmCdlPtOaE81MTahvAYH6qMKuPQ5oFmLBuGII/MrQiZgf0x0mvN
UKRxue4i5Mj6wDs8WFKDXaEQpU3fdzABigYoNTZA/1YevR6c2Z5e1nJpX9nA
sNpqzCe+ZUDVhu/MGQuHATqhsaOeCXuwnbOqqgSasTFgUSArjcVWDnX3AarH
prr4P38fJkVd/wjouw4JvDw2FcHXOvdsdOwioz6OKhM9jV4EpZUnmbAUtZQz
4Qma1+EHUEsa9nwcuXVQMcsm89ikAcS4TcE1al4SIPlB0O0zxvFNqolRQShy
GvBDDOfsXVAi5AkgrC/6JaDELKczUNMCdf9cF5qDDbr4fwRacwV9wYXbQf9j
H+7ta7JsSAw+juldM9gBfKQFld/PVwVlZUmakEmmlW9KM17+JTVT5v+5lkmQ
OOClNTpfTj96S6YvUK6Y1g1aDZwJ+Jm/KABaW0gM0Wnrh4lRxUrD7syhHN1Z
QZidmHyA1TAhk+YcU45rKvCxZSJ7dvJlv+O4/PB7+KeLTZBT2ZQb8yhOaKDI
Hr5nHhllJt1XPlEf78s+0ykXBIJ6p80cLPTq8+fxIxRe+NWkYWMKCv/mEEBm
NDIRj0q+u7HSBzjNk5BUHnQgqc80ioBCslmmDbXYxZwWGA59QzIWSPkviysE
gsunjT/JLXMJ6ZdOwTt++hQrUP49w1VAfc8ldFIFcwCAN0hX5jxcm2UZJM+4
wpB7U7h983AsuAmwXiOE96tqc+w5fx/bTY3mXcLR54UD67n9gtPCPhfnFUO3
xIymdLzU+sQjqNAl12Do9/6Anf5Mfn3sp+CA7O4Fs6NmV5eMCyb1KgAsb/Lz
iopZcwOTMZCzmoPdm3PU1bxyRLFLGjNm7vpu28u6S3BzU0y7071umfFCk4tH
AHuJhVShqhia+mPpVScvCrkkoKES8tjpm6GR4VRl8I3vvfw8OIhViGtadeWF
YJFzySunL1wccpPjHQOmQIY+gtcyOmcML1ee3eXu5lqXRKudxB94WaIrRGIz
30NrYDEOSnMze6oyOj0YzVJUGJfxeKPwC4JB6LKZmXTlh7YYngLCcmIjXefC
kXkudnUpPgYq9y6lubHV8VoQllg1V8OFuh/EmcejtCNjQOxCyN7GxrgRvrEY
w9ueXqeQewwhqNVgK5GwNSa8jItjS+O03797/riHwr7RBLANyjCvOyZ1gaWl
kc2RBJxFro3J3/mskznUbAvo9f9lFrwFYi6R+afCvfvmI20AvcQ/qnRF7N2X
J1OwtODlNsVq2GrY9vT+CYEiNR3/z7EnmJPtq7CRmaNcGZlr85l5ejs0hgxT
qu517uJPR1vWI9xiaAR9TZRJWNL13L3JPr8mksAwu8SdoQjmIcm9VmVa4WWB
RVj7uNu747lAUnKjRdXnEzDgeasXaZ2fRg9Jasm51iM5IFC4q0Qm/Ynt8fWU
qBOCB0wDWp6j9U7BvnR00OgAmDLAHTxH1bD6HO85Di8ZZ5e7cqrEaCEQpq8z
hrVX34VEEmRTiKvR13th++zRas00lkQyIFGaiNAHcO0VOVM0aYLEe5pc6ukl
7OfP3OnkOYv+xhCvRjOQZ8qQ9i62nPZnAoV96Mf5p9OLnSehpCY71hV4MRK1
0SW319SKZUF8hp61zxCRpflLn5SdFOpqH6cZmnv/WIVB0FI77hiOEvIQDiNa
oZrJG7mRbMqx9Ut7a/YADoVo2ffTxkpibm7lEBJL1KGlFV93nq9fBu7QIhqW
cyflI0V4yMLdjXfPkjz0IMltCphY3dJvUCvwOScaF18AlGTL18+A07ppDBmW
TvXnXEzAcDLSXXJDA0v9LCPtHTVorZ2y18bnMN3nYsu3s4GFcAHzDg5kDSIj
A72mTo/ZiWShB9aarRSrENqjG9P16NFIVJMrPHoxGyjkWBioo5drCCopFUor
PdMk4y8exU6uB/9OP/NiCcxWzq4bxzoultQP+M2wDiELUt+Mg6AENETXX7Gq
5bdUCO3u4Ni6z8cQYeEknthj2fpDxj/0SSud3xDJg8idzkC0jKf7/KzMCJJG
GFrx/v9H27RD1Yyycxn/gBJqhroJRdIUx2XYe39yo5ezxiJWUZI+r5F5lJPE
Jen8m/YbOUXy6/4XnBjYAl2L8tlh6xGjoKU4LUuFc7VBp5CMBfZcxaV1XZQ5
neBZVLoh7eOrEyvenO2Luvj00SrR2Ou7lTN0OS0QpOapFikyjglGRsY8vv6p
xFTB/htRUj1l3FUbyPmpKmUspUbpjXartDHq3lJEXjtL3r3FomkTDmxlf7vL
QPveCiDRUsonMM0SCO/87YgaezLfCA+4cdtTJPmCoXJdWByeZMPSXSQJitLA
suLQR8sTwqw9sHpkDXKnRMb4Rdt1amI0wVs1okgSDIDqxVcM8q+mkCDg4S/I
vOuLG8pASjJBawHUxxu98Dq5iDdD+lKKEBuFQY9oxsPhwEvDvf1bhuZyxDUd
NWjGPBwN0UjfNM1dOE8tQL8+NKe0qOCtyidF/vBTCpJWCEguKkTTJUvN6VSy
Z6RHs3JogREakzPWzEAEsG48D7cLucnR0qWlu8B20K0nWt2hs3L3ZzeKQ0Fy
9YuVmO3d0F/HzA7E7RePaVQVlFyWHjrhgR1EXULLosQHnOYdcGuDqWm8hz7J
QJfY/V7PvUIIBMH07IBS8oKvuoYu5bFjw2ppCTn1IGdEo7T30unJqpyDuWC2
R98Dmjh50udCTfLQrJpyH7Hk6olyFMdTM8O7MBYW3Mt1b3vQMUStzMwGRJL3
W8U0bp6Brq5uVFx9WjdQKHd8XhKIWQh4XUsrCGBSitPaik+qKXz63sJi7j4g
hVn0sA/9gAoe7dF1nHSPGr+winGgspEscGghJC8OUDJadjyaUfbOff7tLqo7
oEB7mC6noV92URLqvWIXX/DRuSndSlict2Vu2gKZsl0MtW0qxn6wPKgiH+M8
dkoi8V4kO+U68GKjcvRShtVcaeEFHGEyhZL6foy4g943YOqBqGPlUB/s5xjH
DBLbIRWFwWOo3ES7sqxuu5n2iSu/U3lDlXbJeeuegMagVBSKiuvTkoouspBm
/kFTvJsPZrDzpoPGSDPsTstYBxWqEppZyXLR8OkkJv8Wia+mN2k2LRpDsPy8
o7t35ZKM/kDA6jqDNcKAZq/BZ90sXnUrztaiws6FvgoncB234JlhLWwChXg5
U6D7Y/9tKTzFOf62dVkcAV2GXtisiY253aEN4w2a2QjifLHixpPRC4ht4bRY
foDXFwDktPauxvlAwXNaPPageFBzrwtvRo+wZrhwdDPF5FVdFBV3hZ4XoNMU
odomxAW8/ug2ayjIoCGv2Of5Q6PoAfZKHidwHpeOHJPgOA6MgyDErp3b0Jgm
xIKsIL3T606vVLmmR0scmlW3GcHNrAyubRuxvK6G6IhgigGQeyZI5ZrtjLxg
0VFs5evUMeaARp042lU5UiAjZQNZL/PxrZnVGlXhLKUW0Fh/NRO/CuOa8v1n
jTQznso/Qt8Gy+SI/WwKn45hr7PXWLvWbfh3s0W7JPrGQw/+/625lkAUYZB9
1Qv5DDVnrxMHXJgeTDjewuRdXxHJxgU2+NUPDdq5yKXUnwteh0Zbaj7IJxPA
6aVUY2RYKSBaLvJN/u7SRFlmQAgLRf1QJZi/VcjG5vMz9TtviQxBvpPeZei0
WwrU9coEYGzTmHwh5mGwCFqqOaJWZSl47Gy5XuTDWW7p04JwzR4yRqMtYYOv
RbjfBtnYRMMBu21eiVQwTAf6lt42aHLFme7fms3eW/Jk6CV5e1QoN+LoR4Sp
lLvAj2xAlGITZTLfLwNwwUjxGpJGSveJTwOIn9Y+sxzUVmCb0groOj6PsNqA
89cM7ucbd8TpmyUS6iOFUJGr9oJJZMYX98cJShqFwbXuPd38hkVOuj1cWIUU
ZFRn8W2fjX6mZaAgOfFuH2Od2poBiR/b4MHZ4BXPpgiRZ+zvCp8LDis+3ary
2i9yWSVP8GwJjn+yLl6mxRpGh9aMOLfIwXqm2X7ACxobAhZO21GFZn91eaA+
7daSYMP3cwF8dmooXW6laiRGni7mbk1e+uk/e8uHXwaoXc1o8LZjsB3mS7sV
bzV3h7YGwitdeA0lSLT0lP3GLixRGtzN8YTzA8qEmwLeKIGdM4iIsPp2iZR0
jqfU69XgJMS9nFZWuCq1t9zMZU+ams1oHUuvPblx3nJlxoJTpRguoZ1O/fuX
f5KIEmgdWrRCMoRjIpsRkbqAeRX8EZJtJ+DHeAhAPMoLD/dulSmaQZjHpHQg
AxSDWFreT/6q90HGFNpYMB2pccFJOrOlnzJqhtPSGjojiXvOdE5vLp2SCpna
uI+9cWeMvbm9gNZ0KJKEaMXVUaElQ61eSyoQu/IEMB8hKi12MHmrf3JKwFPk
IKkuNAUQkbOkIP5xGLkR5+eqB0mREJ4CDNihSLQWV3G/zh70O71rn2yvtLrV
UbGpXsiELI8G9lQlWBObuU5j1m/R1CHxi2LjsK/ByDeamt+N6JskReuL5rDZ
RVMEhIJz1Y6cvlIL7ZpZH6faDr7FeBMhcpXY7zjHYTGu6DYqM79JyOSlRKz1
L5mH8ui5zjW3EOV+AagoGXgc3avo6jaujzbzou3QBZ5bEXsQniPPpiweYQew
za7K3+e8mF3a6vGWqWEJCzWHQ1a8UzgozZv1MV7tP/dz3DnmTe2jQsfJ7SyE
eDO/jh1gpZwCEtW0OaHeYD/Vso8LPWuCZsUmG1XGAOnHHlIuHZzjZ0mqUnxp
O1OkNKTF+cN/MoGC0Zbltk5ppH4r9tM5iRTCnzHk+IET7+OWKNX2eJTWZZI8
97unePHQKeAwAqSX/JT7xiD2hfqz6OzwceD4VCqBxWgMZ6MVqP3siaBBzwhi
rv2A2boOvtNVbchgi6EoY4+AqlPzAotbwLZgAZdWN+AF0gtfLfs7DSVKpl49
1w0KZjSu0OFt/cLHDBT8ZmF3B4CYEteuQH4nhD+CZM6GeYolT013lE6kWVDA
VNo7k0yuz9kdEZiCQa/eTuzDhHI0CFBPXeeVVWhionVB4Yu5b6CQfSRIw5WV
zM2ttxI5MaagG+iIjtcFsXFoNg3Fpz7sOxnSyNmc3xFz5w0XXjcYdNsW7Z+a
BZX6Evl1sPCZb/199Kwe2SBZjpC9GuydTwu0//3DEwJ4y+IB4lN1yY079xdD
ePYl88GKTsqTTxT9PUwJK1tzSMaEDNPSl7Qs/iywyLdUHB+202rIhwCUh7zH
sg15vwvi7YNB3Cdy85LkFpxGfq+aNLuOt0lTmdIHtTHiBGoEHJEsUNPdD5PX
JACg83Oo7QzdFH4Rtp/m8c5G1SWI6crezyKWVmUa3TQKraRcJlK3RI24Q2k6
8O0PG0Pn+9ha3mC6/bsfjebnYHwBeJoxN+wqvdr+YL2Tbr/3XGmwPWa4TMnb
TPrUO4L+kuBZziYPRH7s5yQX0SrZpd+00jfnC8DkAk+hrfz3O9/RexD5q1jP
2S+FxtbRXYy+DZFvoweBZ4I+8kKROPkwr5rGp/1uf5icBnkYST7X+dcxp6Nc
qjyy+nK0JQ/sgs5pea2AEQKjJ/OCS7mXh/DKtoqSkekAuuHNvHKsj8F0KCEh
g+UJvdMGiuykgY9/TWW8OXu7Axx+4goaVDE7yUAz4/WhCY/XPzg/1ZzZbt6n
Ptprgg1tRBBm2KNlFgGKln5fewVAyKxix+cH2YJcpUN0ImOplGFKXVBwZqcQ
FSk0+CuajVUFZ57v9uLmrKphRN8mPWPopW6rG/hTI2SPlXg7hXH5KCRyXF9r
vB4hpX6VAJyn4XnMv+Cdku46Hwbq0wIe4h8tKBCE7VDYFBwuDaYQTI53461h
tBq53s+gjMUbG75Ko5fBwpz42tyhIwPcZHhdj+k01Ei3FeEEb7tJXadOelkN
yLzYu2QzIUfUZ8NyK58RvwpdIMCmV90mHwgYNs17hwOjK9WJcD6I4PqQvIud
1X3n9+g69fmCKjcXaA9Hzsr7hrxqBejTqk1PFmeruBfe3POS750Blu1FaI20
TXEF+Y4wNG/Q3iOc8zIZWD9f4EvRG+bl+kH+siHIRS/p5PldJs6hSQBpM8N+
G4nu3Ix+aj2PDq47q0mdLQDeLjGXQ/nB8WARk2PDYbZi+BTftmtfDpfHaKgG
vxS++dbnT6YkQG3u58ScxPFrR81RS2ckxeULq9ZsbDyTYCUnC50rsbOF3eaJ
s1EHBn+1aRTiH/XFgz2UCl0t50dJz4CepNgL1MTmATXjRLp1Bcue91NFa5Ad
iKgtzk59ZFvxgUgJKq59Nf7vj1ZsIjLkqE2mJSbz1lPiraExnIY6GyKBWzaz
m55mB+6C4thnY4Pe4Mer9us9AVwhCaZ05HlF03IDpGHCtkcnuBB8VHUTDyjq
uSkU7UjPN3SL7ZPJFmo8k0BJxxieqEoXmQHu+VWeFovc0UNi1D5f07i51BlG
ikn6IsIbWP1H550AWJbGBkrwwcJ6YBSsX+O39jOqLdBZUCClZtQahNgbDCsp
j9m/6zK+CggQ99kkjVvJ+aBqD1ZaECKuAn0jEVcsV2bEvReeWOFUt0c6ezsb
IcbokvFqb4tqxkoBRsoNzuZd24RiPPGOV9tE62fEQQbmKnzDmwzosgpag3d1
aur9WJZH7LsAqj9ClxYFU2MLgrgpF1hhbTaE26RHDe5I/stcjddteby5z/aH
FjYYuhKJWjmGX0gqTpxPvubcdhRyJDGwODkcXkznfo/xnrHQI15Bx6oq3Iox
vl6ZPisHd09dKxBtaV8sWGZZoRMND2DMIzjD2vlC8exS1TA66NTvcRZaoNhF
DeRqyKk0+x4mnswgim3Oz0f4nC3s+lE4EgvPx7F5SC2h6UY8nM1ktzpWnMcE
y/dSi/Pb+WMl4m8AbFvknjssM/J32hUNFbj67fF4C/O+i76ft5rI60mWWKFp
5Ywb/DArSpp5vKliB81NJPWNr9tozKV4ZS/E3kJ8U/Qp+XOPWE1S6Qw1+zYf
ujVa2e8/gfaiGIkQHoiqUcFUCGcxvXWtZLr0bST7GW8zKzZzgWJct02hqrp2
uLEkhzS4HzQTBKQduZUqiiAVCYvFh2QrGxkLxgakcEWLhd7IFMwbrXmDiSnr
foDrIyfF2Myvs5VZE+pEfd6AktyaCkVfGF47Z+VVC7tkqi9VpyUpPw7Lr5Z+
WWSXyxfQggM42/eIJ9yUS7unCkUe3dB9NC10bVl99IjfVztWvK24xzZyV09Z
WrUqhH4XicBRlu895Caz8KGalPx/oVIsre0Dz+wsPzGpWq2TpocH+N+uXZBD
0Wmo+N+jMiO9JYTm7+hpBiOkudB1x2ot6Fzg04QZIpsS351xlsYP0S7g/ubt
zExlMQj33ybvi8ahwvHrDZSUJkzLu92Ps6fORs2Y6Ul/ET5e2+UU7T6SGSdL
vLhno4lAKlbLEzS15DZGQXAnWns3AKtzVF4Ay2t8h0YMLIepn/fiFclMJLB9
BVVS0ptSCgQCJY/0/DZFLDQo+OvepnQUBjyWROfH5zC4N9EVPxFPdyS+eECw
qGgnP+XblaydepmKza9i0OgjZVPMZev1bYOm0Ma27hksH6AuyVn8Yilcnw2C
wDHGb4n4p42HFcbpbb7bonVpQ2qSvIuXa6IqbvJAtC0dM0krxk0GODHu/lNJ
Vy/K3zy2rcbu/JpbljWw57ssuviYAJK0mpObBlSB8LsAR8fWzaXRLJZPOce9
nO9CHshCC20M3mTUvbAzUcFC4xKQbvd3exk8P0DItnaEd9ChctbUpekXF1tl
LNwlzmaFqOPRIyEmfjAj/yKlnh7cwV9wvtcJPvQcvJlf16vAYKzNdT4tGJn8
gTUAnmvAJfZZyn1PEhesg1KGXm9+ImbhN0twuNj05tfLT4lKDP/Ljp/XXkZO
xCJnsCVqekhskf8WRM+qL2/7MRayydQ7uvkyORzBjwCrS7su5EbVXFDwK6e/
R9INZgc9DBtKoqkozBWI8EVtVxwhyD44fG2U+s/1LbFtupwo2gY1VlDjlknm
nncaR4cNkTlmHKW8Vjp2NvdGopLYcDkmoLmGpeDFvbxVNMLGtuK1b0ExlGI0
DRUr3CFOq6Az+ittuj4pDDAQS8QwaACMvs8a1Jy3kXHmGkHNqMIUUl7UXd7L
4gwOJxgoq4dPyoR2o8SR+sVWVzqdwGsaYEOhD7lLUqZ5CLufJCU9pw2HcGbe
3fAjvuTwUmxFx9Ss/Kh3YpYAqVW9VOZ/AeV/2aT7Lt+8JZYR/2X3lvG5fovl
qvqCWKZGOwQWcRroz2qDUyF/2yp1Tv+5vvmVb9xSLiB94hS3+H/0xXqnVm/B
rvr7E6ku5/er9Ah7aRRlQ1oY40dYi8f8kqzEwGPeQode88gKkYh2iWOzO0Fi
72Dztjp1JLecBEjEErhp3cqS1NcsUCFMcKrhZ6S1H3Rp0Sf6f6st5isopSxC
zerQm4HFVLk4BrmHGobHIDFeyXATxHhszzMO420+oWgJysG0JJWQ7UFXJHb0
N+zPbD7cm33y+gft/s742pyZL+ZX16VLeHBeO12yNcavyh3fhAdgGkzJD4Qf
wK4tns7YHtl92+XI1x+wNK6OYo/KTFqyXN/pDwEVgjdg9NEc0jA8XDOL0xo2
XLQal9XB8qw0cj2UPehur+japhoxxKKqOdfd7HT7IA43bkCUjgkVNEYAPCBT
20nRMa6ut3E+bZd5NcXsE9iAZTUYYM/243piryVgwmF8yH6FIKRSKfk9AKsw
Z+eGpLWp+3F6ZSPEYyjLNYQJhmW4dIN8QQ9h+0W73qWmuFVrGoq/148bSR87
9bfTi+4IyznAZt7svTyUs9BwDBzB2+sp4x2R2n8fts6xKMEBLYB5NQVk22te
CZFzEcgw5jWVWDX8GiCUD7KVyQTgm6gha+9qbbPoBPOq9MsRCmNByf83K13R
PldmKnV0MtgdbKIJi5kwZ632rw/JyJiB6N2/s9X0xGs1Et5bD2erHFmp1HAx
rQEur0dumB7lhzr9syqX1BwZF5Ou9+fJmLV6FbWJKJX1g+KkD8ocHruK+o+g
JQnygppQaPfUVyUpwhwxV7NiKAxj0imlq4rJVLZkUpydqXXd63uHf0d1TC6r
slVYZSP6i7ieDJUkDx2NCoCATy4q7ZHmPZxQTOxVQ56WgJY2xurzt0PyZnlS
RH90FONjktAgg/SuW+fMg0cxacYnW9xreWNxMCc1e8GzKYxEfQ9nT/bV31Kb
EVEPFP4q6KYSpoPsu4MOyK4/rBgVbsB+WQdb39MN4NJqENtPlMl7/+QZrEoR
0JMKyMEywCCZrXNnjHz6zXqldxSNMmvfHlEXwl0innuaek/5Y6fo4stNE+DI
WEuDXFISFQzXlqkvBKgBro0kG9XYU3kO1te8Mq1kRmh+pYr0KNznMyhkV9rN
zh7jHHGDylBIlZ3ohN8lOpYLjUR+bMJBRs39gwv5BAj0Tjx3OOmugVErDqiA
7KRSXQ4rsncyBKUUDdTv6eQ57zB0iFkzS8CWCJfGOcXxodyN5gYSQYC+mAii
nzIip/i/bEzcuSQslemC7LVepjQ7lgQMqUPXQk6Xxgz5f++AtLfGCIvUNEH9
eVw4h/UinzUjTORwdZJqNHal7YVg6R4vMrnMHu3+tJnO3GZoBgKQQbgvTlPz
e90287KqHnKgV5X5JSUU8Wwo6Z4SIz7Pj3LEtLSzEcC2nqSCyqsgqqybf+wn
gUcp66sF37NgGdyK7fkjEU6VDgEt82pspvxo80MYxfPRgpT6GD4T014PQTNO
9vku8nDS7R3rGctA5XDmt0y+HSO+hfjVDcswh6TCg3I2nm+5Xpp86hcCxaSc
mgi6e4RB7JjWwWw3fkTSNN0dCzyexp2X/2LahYom5sNLBMIn4/8fqPsSrCDQ
na0l8dOrioFocctF+X5wS5Kwab++q026kBtsDI2viGFo/IZE/RRRAVod7edi
7S5aF7QkecT2u8vupsyqflp77BHnI5sSVswlUphiQkpOPpbmPoJrCteAuGVP
h0b6uI8LecXg974wyaDP4zNOo6ZVBVJzqMxrHlVesBXitqSYB4LuFANPIh5S
PPaBqTmR8GMk8SCfslRDdzY4HKqCM5P89wQfSl8GMUqASN/D1XSoUznIYDWY
PNQipc0Vetb9SWF2DqfaVtXX1T6284Ocnu67uAh5vthbjWr3cP2qiwSfciAP
kH0iBfnRrjTUkXl8T9JWfaOyMY9rSMXDvc4L+MStmhDGYWyPfeWkg0zK5SgU
pSTLnaD6zkqpIia2bSeVVlG8wBGa5sIQ4XbBqPrAHvREOcKeoMT6UTvG7FI+
ZWRNqAFQSE3roFPhFhhj3XHd/V2rVTnf33nmUU+68nhvW0WpYNGsO+Q7SjEd
VtrAZU4gCu2KCxwg03+HoAwuFlUeG/Sqsq6SDlypIyElKgAeTFdh/HeIsMis
nWTLmjkH+Kh81VKxxvwiu5Ir8B19s2+rJGInL2Kpel3mLOZnZebgQK9vP9HA
RVIfDwJSadiB8Q/9YrokRaHNokrK4SEEUKPpvtcp/AYwEpdA9EZpFNxFPMhD
n9hM8UHmU4IMfnKoP+R+RzAZPD6lhpu4CeWo+TebkupERQ3C/QoJ9qQaD3lT
6IVCYByoNAQLaO8RsrEl1EL9ex5rjX+W5PU5TkSMLvpUZcomTrrAHagPPPuj
f+SLkbuGzmfb1pezAOqCBIy9XQk6867Me+7+TAlecxbxcaBwhA7+7az8Wh+o
lNWk8fcezboDYT4BcmWxGuMRcefTcWtGlJ28Pp+QqrlJrwUyazGWEwvwdA5C
K0IG2oUh36hduuMCOPWDPi1vx2u1PgDr0LVGmnUuJEmuo8ZjEJirbFdPmOYa
9g8gcC/ygEZcgrWkqpyM5neljKm/LonCQBSzV0wY5fUY4w0mSus/k9PDaP8k
2ux+72Op+VwhC003SSKQuuDWDg2FSP6O/qWx5RJfdw/dVJ5Yk8ibreMzOaQh
2psIz8LBOteS0+HtbpaepaFleffwAyoyXYjjnA/WFCBImJEMpLJaZgXVDSnr
MJgzsO2ERFoAyOb4XXH08jRKq+AVVFpjCdvQ8/UcK1nszt/HgXzRgzVK4VsK
mdGd7hyYPCKPs9558EWIeWc7/TrMwhMl3nKCt2Um8ss9FmsX0FJUs0iv+ccO
GJLwBPVUz39hDh7qo0vxMNClJr4M77BU85by59oHSOa80N3IyiDg2R1agdHt
j24oc6iTuNF/QQb8BYqZO3j9ajlOCpvSC/y7njTBCyYz6cQ3uuUrUuoSx17B
cTe/VvU870PGi7klc9Lbobipp9FSwr3FZW3gguIY4C2DQvWwt/NB91Ct7FnC
j0whHFjOZJfHDsVihwaRbE3LJaiOmL/9h644tvRYpfi69kt9j48ZapbEnNQ8
q8cHmfWZXDFP9JNzvoAd6QeRH49Em6uEFygZ9DtOeiwd9ya1Sg6AjwoZ4rav
KaY1qMvzwqL8IWvFHt1ahwpuwkpkJVF+cS6yXidYuOMK4KFQNIiT5iumbbw+
+efXrikBSq3kBrEOBRzmRnkqhaBGbEER9zq+WMTUqAVDgL0USGDQ8U3J0W6V
mwGFow4jcLLvW2stMGcAqOpbKw3CcTiIZNDgsKl4kkorbYYV5XO+8w+4dLGM
aGCOYKfQkP1RRQe6n9ehGCa/HsXFYXtUr6IqJBWYkHic+swKrb5PxKpxf7xx
vaNaUxuvruFfDbRqTiqWUnXKlE2/MpVVFctEvqNZCCHcl3PwDTq9kYJlHVWt
daSMHGzebTR9cpw/X+bE8qfXvaq+RYUR0h15QOvCt6fEmDm8cxW7t03geUPQ
L6asjlHCx/qPDd5L9Lr4pF/cFqKLECniR/RfN5FMFIuEUK8Mx1B47jneIwBb
0bPfr4H+PbBP8OYkooS2KMIAQabnIU6pBV5hrXwhO4BwdK1QAbmUeSiHvgTB
zqCHG4phg++XzuCSem8vO1o1GyUkeMICYKEIbEX+8HVaCqG/QfEnLArfpwPY
o6BspSlbn6IYGJkfqCxlRw23UiAjsShYJaV7BHpQ+evGJTJzVy82dr+qwP98
QnsG9WWhp6kqBeMYLNO8VVCq+lslW8ZiNSYLqEjhfp3O+lpmrteaQaWPzrub
T7++mibyTSplnvcbrMkC3tgQPdnVgJKWX2MCZ2/MCXGC2kFPSLQ9hm0Vgmqj
nuk5WG+umpyiTMCr/k3n8ei2J2iiTN5CSiVZZlybe1KmBAHlO0gc075GUjgd
AAgPlsfVYNdsZJBVmwlOamwMyDpQMWBKXnlNZJ2sTmtD5s077R9m22CU/LvW
Ro21QXe+Ne86N4tDp5Zhr1kClimvCFGce7JMQq/31lLAEcTLwvL5fxKbAVUy
vF9cyq8dVf4WDpoi5tr7j/Rcu7tJoxumpDd8HebWXTonzhkYIlOboeCFEsAw
DVS+eqI86UvnujelV1CaBGdOedsqOpLtUAvJGJ/OLr9KNhT4C5P5gTSYwf26
Js/kbbbhE0l/rTxdLjsrr1CtwaMAC+md5S4lc8OstQoGYawRoE/CxzcJjnGg
MJuEXiFca9w2DNdJgaSYTVVTh3jYvKWlEmZI/eJbGZh7dbutyAUwTsJOaw+q
0wzVfGlzOaJbrFs9QuuE6NB4aSnCf+2XzeavZpPMX4iVU9ePMqK7jVFtcSTY
ytxThOOTzyxm2sWo52Cmxt1AS9nfiPqKwcuSAOZqN9ph0zRrGr15LYEqD0i/
8U7V+DREuxHtwhCw7yavRefc7CYgtsCYeZNGfV0VfJYuVUJ3ixLbG6hc7GL0
9059jvhGMa1DUHnpBnZ1xN+OeteYWpOpv3MflBOAQ+6SLWlB264ztxb6w6OF
pS2+bWyqvkQxJpFJ34MdmQn4JW/nBtthM+1ebYvXfw0R9GgIMOYhxakUmNmR
YeltqSQvyFTd5eIKXEPGcXwU3pxaq13Pn55/aCaACXSBl776En6Bbyg1kclP
fRX9QM5d4lg19X115ZUA/v0kDuHsWreLsojyEzWvMbiqIpx/5He6FLq6xZ6+
hN+hJ6NVrQOGwc3YppigyvEZ8bHaf8MUKLj9V6jKRzNrv/9c/pdqomFdw1qR
6jXkzjMdP86jBrDYGMfdfr7EplmoTMri3RUXXpKlhqnKYKzyc1RFz11RPjTd
HIsB227M8gGGQZjqh17j3NIVu6QVq6B3tfxlUCU5JO4vXiQ9cTbasHA2yv/E
n/99DFTexDWszf0UJuH8QkxJkagSVMELzjjo4DuI0bNb1IeiHDD4wyWu97dn
FLBqGfwesC0i63nWebDUzU33JW6TTqnIrcYq8vgeAoZC1XycQMwpBgnukaoN
b73j6icQ5MZ0oPiohXQYpeblXMtIepc6gtrEKeGphqcnKTqgeSlXU6kfpMwu
kEOKyEOjJd5uQFVsI9IGOBHCH5Ny+qsle2RJo5qQo0+tjB3M50Em+sGb8pbt
vvMV7uWjzfh+uhR7V+dlnDw6qtt15ftsn/b9T1D1M1U8xztsjWMeqLo62dRx
2oyKhxy68UZ/HMI0NOqQ1A5nv+XudgfQAMN6MsA5qc7Z+p0ZXCMDkoIAJLpm
9I97R+HQtWRhpuVLDoiv/xcxJh+IGCNDIJ3rJ7WvKfX3BOoR0bGDuWkIukJK
VWDASlkPpKIkTfQDcqKu73sUTjZNMuyFhcZon7jp362kyUEAXHR2eJ8PrNAT
oM6IejCRTd3sIZuD4WZ5aUsRW0wABpttHcWqhdjrWknZQKObyUyZcqVMfOdq
PidBrH7gBqVgHsIsxswXb7TX3q8LMFsMjNISNAUp2sFVUZA14YJOupBFgt3C
nEDCK2V5+2XU7ahJUaN30a/veHzEhG2dinDtYBIlULOG9wmK6j5XC+bbLnWe
RJb1Olszycd4jkGhd30rNRvH356sC6ft4S8I5MPYVNPuZDnGpR64CM3qnuKh
+QKbEUuHFyyaU9CDAnVR172NCk6dmAB/TqsUyhH5FaOg4YdOreJ5eYtvHsUU
Eu5s+ETFlSChESXY2gRb4DAEiTz5euufiSIBrTihAvx6pbvStD/IO7DoHeBs
7z2qALVXKXZ6MFE4ysbID2QohvaO4yfVnNmZLnzhSg411RiqLjfIDlNlrKD9
+7SlV2ZE9w0azK+qaOK3qBa8QwwymYo4YDWMpneu8sixKLa43HmIxsuQcAb0
AHUNaCSQyR9xlsY/mVnGi0nsS+utJbvpY1m9b3iLPEuMWgwA57CnyBAKUJXD
d3uyKJJy9XBphY+/PBdOgkunQ0hiVCwUZ6bY6mhsC0FzX6PM8SjJOhDTg0e/
kWjaZDxuu+cq58smIlzuYzNjI+Zir3tg7Figqyujr0PA0J2vtCyXin2JJZip
R2Ol7S6KsTKFdbdg7m9n5Dn0Y+SUvnHbVRtwEvNx3eaImWDJrfTvs5gZkZKs
EVOSmg9VXwScaTkL8seulHyDwY7qLhelpU5PlOR/sdioV2POat/VMVDk9yum
YCP4s51D5JdfBrTG15IzJPj1Wppdbn1R0HrUtBwYdtaU2lz4MiMDk6bzulvi
Wojcygxt8LQTBt55RxxPNipnHOE17YFxlAp3WXfxtA0s90coDasZ4C/+Xkpd
9G7bEiyC9r9TDL2ozf4DTl05XRQ2fmiXIPk615h6yeUmVxO7nLhcCLDSBWPA
ppQ/22nh/ru6xHkaDOGtL7GcNFA1at9YBqd5vKGZcQq7Lt4rE6c1dYoNGKY6
iIrd9fqkN/iWJIpv/97iMqcAPJq/O4H36Rrr07lkafNQVa0Q1NdYRSqU+jKJ
Icwv65pXZF53T338LCTv9vR9vw1KaaPrsrEAesLsAV1Wevp7GebOlGaCZKxP
zXBNo48M34Aixa7bRH+y4KwlRR6r7lLuZ67qRa76NjdN9TlWXMdeARCFiIWX
mzcudyta6rSFRTaUq+vR3AUbLs9V22LSOzukFZdAXt77CTJkpVxf0ZdTiqwo
oCxK4cVkZ2iGu5qeyWXh0tBL2ra0By7dh4AK0duUuxKk0JDXZKptbAZrJBFr
wqIgHFAUF7r04iUkaB1o/LZlRtiQ3qPra6pE4Yea78i08zP6vdsN1pWpOou+
ejajBkXPdq10Li13cfFLMRYJNcxxzcpF3DBXQVwtvQGbXR/3Om6RIKd11f0E
+xfZtCWsyut0BJxCyvCfPGlObJqW7G6n+iDjVa+Dkjz9o2173hrCeBRtbuhk
oBIVgIoXRNCyv5pOjbijOdZUPsF0YDNn+pn7K8ajdNfcP4aACns+cnQx0KVk
TDybIs3u+dsCa9og9qFcY+On4JIB8tPPFRkPFfSsEiS+7knqzviMCNy7M87q
gszyVQakAGffA0KhlL67fv3InEe20tIsUB9kqWv1aA0yS5XiqMnK1Dyr2/b2
GucvYORUy2Nraa7fqUDQNOkybwNitT4nXwV4sNKLSw3lgIRiNsSfRhWa4B+S
VP81zyYemgB4NnlRopt+pPLLFiVfjVt5Jngz3i1ipUXn7Zu01/4JXyEReAyc
AfVBcWVTvnQfkK//RjefmfjGeE/fiRKaD0qWheDqHevCidKDgvpQpt+nATvs
U5QS2IupU4fdj2uU+cVqnarjwswlE5wYSRLoBPT4xIawfjge/aGlvf4+ThgT
9vOfIHlgB96Ss06Rw0X9YVqYHtig6yvLCSrEJJ6SV9Cn809Mid61zBwcM2BW
o/I5Jhk2YvXUFzC3Io90pwr6pHqrY6APdggPt4pffJNtz2GuxmKc6SIeTogz
a5F2FClzk2kgupNqDdLLWTzj1k5pqZXUZkj+5CgH+RmZ44a//pPceJkcl+eG
vGQVZsPjMi78evy12XIHb73fLvGtdSjwL6WRDwzTszkbughjGqzV64hraeVN
PN+3ifsO0nX5DKdYcLRa0Mt0UY5F9Ng4e3K22QraijWR6VZ202M7vsS2kOWq
E+P99vZeuTo9OBqUJUL+sBk4l3SkfYsgpSeUhaqQ0dfh95ZAqk9kszKvi6oU
lWYjW1e+kstz20ge6ijjk8zw67zt+RxMseRna7nDSiuIbhN5EcNChQJxhkAx
RPwiGtE7/Zc+ir9Wezd6MGDJzjsiIqR5m6VpngMi1VkDycpouuGk9ry11EGA
sYEDuxPt5dMaQEPJ7qCPnRZ3tlQjvKoLUcssTElFOgwQZj906ssCxBOjJ2LL
AkFEZrJKiPR6g/yJFm5XFWyGGMTB9Ky3s3RA66uL8fyrk+qK2RDJXX5BvKff
9hDzJ86x8GdffRX+c4qBqSDe9tGAxVBUprrZwelALHF8IKcbBoeuKYnSGjx1
IpnGGfjDAodXYns4P8qo0HLINk0jMrzVnLdicivaaL3XFZhNsmrIaTo2T1A+
3zeyHJCuZpD3WmcW9nsxsOrB/0Z+581wE/tK/FKYcQeOL3SxrURWqmmKj1hA
PKtYUujYxTd5D0WbuHdWJZSWNdogzxNl3hIz4kWcb019DtjFflxpltrRfdg6
YOZeb2YJ+bLXKM7SyoCd/iwIjJd5DzEgOtdwuTPM8jNoX2FqaZKjEZo7eba/
XR3VKuruBeNWeXK1m2RkWYp8xY9Sf6YvR/mY33ncV2e3nVQ8/8I5lH12VgAk
8W69GMkQ+5P8Cb8nZ8TIiR6IxLW/PZf7217tA/VkrUL96fExVvcB7TNAo7QJ
ZV9CHj5dIRGm12DXmINo5X2S48FQpwlkgwZNUi7zxF/xtl9vRhJfVHx587tj
9ZPpZqC4z7zmbvBNgAsT5zETVXxjBQBDQss+C7JKRQYP5iVSk4hVqf2WAe4h
IK7XQl+5PMeNy2j3OrUmFJTsWPkOsVYWxIixcZNKwAzuJldo3t8W+9JY4rFm
yJGqdXuR0IFnITFIrtg7xKblLb0P/a7vJzzAjvOp4IksQQmPyt1IzC3ppSG/
pyl06ll+yj1K2tW4kJxo5+YdAg1RpqEqZhOZNRgOGz3JZbyVRbYrIXTkrvJk
kK1msB73Hako7pIKopC2csFc7SyTTwfaHPE0hciBzy5xBOE0ADvxfoCyENpb
1e6UWRlrNwlR2/wSurnjkMu4bndLuIJXBYv/zoad1l1N5jVAcFAKTzRg0IDH
NL/fp88PIsqoyH4i291ND/i9ikd6y+FpzWqqbFpHmAVSRT97EgxjoogQOmRW
7RfChpMHYVNnMzo1sTEpR7tRmlv95bALleYjsPEod5g6z3OVt8tRWrOX4GVI
bxgaybZ2Eis0dO80e1T+60Ffybf3VBb5NOSVr3P94U077ePjk0TKaAxjrNJO
f1ur81Oa1HDKvQ8eNrTEYUtPX3RFpbO3Dchf09DNnjaYMOBcZwcWrhYxK91Y
d0ffryTfVbqyuDOkUHVoTAvlDHxhQewoRBOU6mzcvdmRe/7qIRL32dcfaod0
qVi+Om3aQKw2SEAdLIPWoarxhEE27Xl+ueo86HFmo6gqH0lRLcSIVjhxJ8kn
ZMVLEkAzQNgNM6m6bxTFFWE/OEcF3h50x7bOckF9/1A5WKLjaRJNIQfdy6Pn
GIXtRITkc3cmo0PdJ0N4hOWi+6iXjIX5QbfvICast2d/0mXx+Vpoelm/DHwS
wrqppgAIkknHbYeD+f/E4eKySX4Fo4YeneT9ZWZJ8FAPxNkabJLRS6lZYP9m
N4qDJses3NtpEgdgVTGggwteVvZbHGZa7iusTNZrMfaYVhJRYDJ63edX6zlm
hXaDKQpVPSSGqH5z+p7rpAY2EduSAshX9wffGf1JysYOEy2TPYF3vhhPY68O
yzPtOkVqWV8UpZBJOPrzp7Rj2rkTDvydNvHIAcrqR4Oc8TIo9KxrECGIn0qD
YodPwdM+ILdXcGMqF8V0ayUEDirjoP4YOS9FpWnbkTp1cKq7xXxPQUzbtSKi
TH/oToSIEHG/Zfe09IDh65MhLia5aFV9lcFXdcsORIwLEUWkMahmM8tu7W/P
oyg17at28OmlYZT/NYufQ6h8tKeAN7GvTpXWvx7m8Ou6l4TNH6aFHeKwfW0m
rFccagVbLPNQtxrwCfMNrqyDoMrpfGL9STZCOUbntEeU2ezTEfCHeKqwsoUX
iGjpzLTJscogQBaq7ap5hhyF/W4e7L+VTliZX4AExwmxb0HYid4QEyrPftHb
CE++HZLdgb77tQwG6OY/sBCp0B9LaAOHS5LXJi/GgtZ2LkPafgyR2cZO7ySQ
wwRi66gimKza9ZzZqWXaWbrtHtnWh/zAn1VVPo/RE1dQxCI3ES8CtaiIBW/E
exmwe5u9sl0uVnubjbRYxlj4a2wArkmw02na1es6fmCBllunvxI/XXwNXS5d
hz5rmDPbTtiDJPEk9Qxw1lDdO8SMHyLRJp3LS02J47XeCOwj0HxjCViHenYY
hdzk5Y/CjDqFEUmNVexwD4bbLRMsc+bonaVTRuSplRvA8YaUfnvb2wNpgpb9
Z1cYHFN+XiOAroN2R6iXy4bpIMTn2m9KtN7P170ioYPus91XlFFPnGbBooLS
VhMtHaZN0VZmpPX+BXTPcCANncxYwntgMxCce2AmpmIGeuPpqCyGaAOrm8Oa
XkDl8QKpKBYLfvBLOFwlSlRG5+/o1AyRJemwyxOg8mFI2F3j8eb1JMHkcYJ4
bURSm0KNOcUJSRY9SCxkvpMJ6c060VY36okfZHwBKcWvLq4mnOEpkdiIC7g7
rZYUiAd3XofU7B8s92vkhu23Ap2/PMoeZ15X+1GDhdeicVaSGJ/RTZAccOw6
u8PUm7A2Z7iFWmzVOu+PMhAd8XOaxKc63n/so8qVztyL4JGZJFU+s4JKZueD
KWzVMpuHTloSJ9wBYZx7aWw+2ymYcSgJUZv3ETnArTGFFZuIAegUS2GVy3rb
XRx4t9kFbU4awqpr1svrpEglWKBZ54YvKREG8eXLhSywAOsFPbkvroMc5efE
SimmT4FoUWO/QvSQTusGNYDlkh3Ilj3yrgcIZT37rpouXxqrOiFPrh1dfxol
4OllE7bwSFoc4RQdCYIR38Obu/zP4wDA3RUE5kjJjCzCN39XuQEr1kKz4kDv
Mx2Avz7z3j4vBxYCjfyOdgTTh7+gNPjGvqizYoF1sM0yoo0jq8BEnE3jaSiY
o1FVqecm0AO/vNJJu97LEkmoXHTocHYM88UcJRk03iHMywcuMuvxknv2SaC1
3G/0n5LDx8eZjw1nrFDsxtFlRrEeXzErv5r6pArttM2fTwEna02htg41V+hd
Ur+zxQdKHoJY8Z7+FcYij666NXSE3J3mZh2kQh2CyJfZOUYo+1R1J7BWEaIj
I11obC02ybmd+dpj4yR4VTABxNv60LlPeG+M4mxMJeL3PewdNviZy84GHZIi
gs5YCq2GswT0rq0NO/kgdj2lX9JNpj3qCSDbUELmqrVf//wMNo9QiZScdga+
C8h31lURF7ONTtig3S4+JWkvPHHz64nNzZdbJqkcOuhAk2LyDtjNH5HwLnfl
gDi0NoLdsL55DZlzWylpYoZetwruPG1BSp071P60MURX24Frff823IldSeo5
IFr2ocn5BplPW+SXm8r9kYQInq3pWTuRtixN28wURW2Dpx4KFCoR/Vcjw+PR
IEiycVqr5qzn8RBLkkXTbUcBED3FO3znoyCxszj9xSCRjsqo/AFGrALYbrv5
N7KyoqtkNBBE5hrP7c9p2jmxeZxSb7HxLt9dy7lNgpDhz9AEjKtp8WTgnQON
wYHnAi75AxRBnQsH/89HvSDezILkHhmyzQgCqKDUzhycayfQwFu7qq0UwcXJ
UerPP5XP9Nam9el9VYGzjZHFZpMTGTORwoQsW4NSULYFTrniAazsu0JJMAxb
fVp9EE1DzXFchSAr8XGHohHzbJFSK0s0BqfS9v3YlN63zhPW+gXQUapiXnIj
NOjLPK0sUnShksgLDnAD7hb4M+heRUtKQ/dda+piRYaaIEn8qDSFRl8xSvBi
vmzi0n+EvVI9os9ntxpr4M+PBXrU1rlqhOoJugG9iFgUdrxNaPwDk1iTXFa1
3kxBrL5v4pt5UwOe2onmZw8MSmw665Od2S87d9quaZ4s1IBZOv3CqtUQnh4M
058/lR5LOzrI74+PQ+CCs6kqUf2vyHjR6eDDrPue6IS/QsgbdlAP7djo7seQ
bJnFx9UxSYK6lYlWG3koyXkG4wo9dLx7otd9nwUP8YEHRim4BagVwvh6AFtH
3jknxrBpK+Nd9w+CL5vRqX+QElPrmva8A4s78/dg8GfettJSpxi7AUyFjEF6
5Zdq9HI79gkRnWU48L9EJIcwkP9AHVesk9zCuJjhb5417genw04EOLUokEpx
U/Na+SZL6IP/kT8NscP2HJNVV7rZWWuWDCeumArk1yfS64Jj8oWgBgyQFyh7
A2TqSJELI5r1cKxJlsniUILkO/j+mlEt5x8IPCRDr1DSqcP5rqiVxk+WFYW2
X8GSwj26a1vjp6oQNzRRTizMIkpZ9zbiJJVLE8hGh7UObZko38IKeDz0Sacw
Uj60sV7fhFLyTGxHD1meDNm+Ts/bRdmxoAkEaejc1pzOHDml0RxXFxILvavq
Gd81SQOexmwWVc4baMuYQfIf2H0ZPInAm6Mc1HLi4lqe9z+SBC/+qlEOXxlK
ckxRPHoWVXPIqbFPLomU2O1RjhRTwQAMRuXZS4zTag6YBTkS585hy4IK49NW
1EgPkFkimoEqRTIgOkkVdxJ3fkXXB95t12tzI8csxbXVKelpDbV0kXkEWBVe
SYl1xFMKsDddAA8F3rkUxIay8xrrsEft9bJdkvz8KoronPe8vds3YMHlko6u
60j4VvYnW+TluaR+MAGxVgaXPnZrUAKAYMGbqPmT3f/4HXEuo6ck4AdTf7/J
NS4VP4/uspajkCim/DWIRgU3ZcKYkJUQuXeWOc8CqANTlFRqlr3le5ntPg64
cdScLd7zTpgrHb0RY4mtKl+ePy/4h2Jaj3gu88eSLuCUsZcsfyc+9fglsj03
Q3VoXpCc7Q2LRKojKPZglnJNYZ0lkttdVphAVDXs4c0ontlJyBajP8c6IeE/
iqj0LsOtaYhqO+IF7I5rPXk3qVO0lmBHJFfj1wJjj5H26iLfSnd9SUYfE9rl
rQiiVzVYaPuhvrXS7HxwO5ItqmyUAhk84cjRHoCJYhrSUO71uiX/zQL59sxE
jwHLlZRwgLRuN9FK1UkXtUZS/sCxzJEveoidxcqTYCtjmdqcKK2ryvx8Co25
OenoQk7k07yz33DFnRciYhA3PrrL7hUmLPcWZL7BytUD8VrNKYKN2JvMDVqK
KcOa/PxuHXeX1yNaf3DhyxoyjZNhl9nNs46g9GUXIs80AXkMrIoS00BRzOE1
aE/iV38hlA0gYzP+yt2H4u/s+QFFdevpgDKAZa1t5YY7YaKhNaV4QbYf0A5Z
AckJR75sI/in9hAZg8whLbionS0NxotXHZttsqVqhtcOqx6r163+9BQP9m2h
Fqy1LFYD3G6PTxCA85/NdKTainT7hjlNwl2d3GRwRjtL/dAfPqMDQeKDHtbD
atOCrfxOlXgmDvWmGNldo1LBiNqT+n/QyEutu3f2z2Qtl7tSlw2Le1SjGehy
1DilJt4vb8kqAZWe+viWJAXCBuP1I4ubkE+V1dMWAI/D6YhduxM/5w407ICD
EATDTe+dUNFlLILABnxdbOogOc23gYksoEFoQrvtpZGVH04ZQH9MFkuq9Hbo
2HBhlZyT8dcvgtDjmCy0CcNSySftt/lUGObCx+Z5KXWpXmWOPEqlXGytsD4j
LUZaSZrwifftlcC9alE66JWX0wEkAvpZjxNyHb3b2dzmTqU25c8vzTv+7HoG
vmMIEcqoCZmzFTJNXUJ3nAivvsZmX3XgioqBGySNv/eS3/lDU6RsUVycrD0q
OowAxlvHjlKqwNTVmKkPsQY09TNwT9dScmemf2/KfQTRC4yQZt2MAdPnnUG2
WR7337DTEuHMmjvj3uqYKA7ORjoG6vtlJpITa1n31cD2w3bNTEA6NzNAsT/g
vGAlGzT3iM4cjlswpMEWQ7ljAX3U1y+Ds6bvU0RyY4lG2itJBGuhWo6ZO3XM
VxOy6788nt68hwfbOCL9Us0SbuhTBAnIVUkJqAID0EpPjCy7XNhVEH9NxfgC
gjFWsVakd+KHfZdH2B1fOlZZ2PKh2xHWMQJGRZc00mWCHI8qhYATxpMwBXKh
YRsgg6h6RiV+MUIJoQZD8RnsleqL/ngyXtbMwi6qL2UGIopjprkn3Cey6f2M
lZ1U2e44t7Rc381RFV4BxCqDKBlo4vRwHDR7CBKP2hl1G/aSyPvxbYrqUEWx
2vWjCTdIAQOPxLC4XQkJ/07jWjcaFHej4lotAo7Fo2uFPhWW7Jz3Ri00+alM
PeoByfHzvMXtv9s+OYDxLft5jUioir6aID5Gpcqhcf+0DJbk6SBSbmeOCJCl
fv9coTe1LXirWX3YRVituc0wJZdhVQEev6+0xWuHfxRj4IN/iHZsH8WGg97n
chiiB8DfaXu2TsEepOR9t0XteaKHs0SQdIDDFqpGY2op/pqqPAWRLEk1/YtE
axEwNmcbHjnETnnE6VrTdrU+iBL1HLZkNQorM3yOrz8smVtNrVeMvKrJWPJZ
Ap2/F5rc20LHe/juKTnlsLmQAI8GoslGHGKeBE4Avurtrn/qIqkAbEgGKQYw
/cuwRD83pKd7jf3lw2q819oWeAc65JBIzVlwjUAnCZMSqKZwPiRtRIFy4jn+
ND+7QRZtUFl0KTv+zxwiiHjqWK9zrh+s/AtYUNg47QE3wIS39mn6+B11Z/Ev
b6IqD4Fv6vcCq1wRNVsjJWtI4iQL+zrEwR9aKFsX49oPVdHP5AfyWsUW36Xt
LRaOx1S5WRe9BVbqoX4Jti/DBQIDcTM02m/+o0axaxzrwCtovqOpqglIybZb
TkmKdSpfCf71z+IHBQHDUAfP3jXlPK6w4l9b23XKoSpNcb1k3jsJ75eedzxs
fPrEa4N3FsAAZCScp7+daqE3Rg1pc/WwgA9IZZuc+GSW4MDMnQIiwxwJCiqI
mGRjY/u/iAxRe5wPPg1lN+weZ8rKMlZeMtPhA4EkdUTCGCppE8C91NrV36V/
og6HayrI49csQryI+PeHt7VC3i8KdcFRZA8aQkXiWnkKVwmO2uP3iAcgI9ym
X2GttCztfOAm+BMrKYEJTzEN3KgXk3z7SO81M16U/ODkSE3sMFp2A7ylmFhF
I2k4OVdd80RFnSr6qX7bneUUnJa1Ntt6c3tWGk4FuBONxoIBkaBqRhG79fb0
IAHnNYrpQarfxMSwSlhFjdHGAAzPVEhiuLH2mJOCUfQbQbHELNAOOCscJpzZ
Hh7rkfLaiiWmApum0RZIDd1N576DS+dYYv2i3XEGKJB7QmpPnLZH5Bpg6hl2
XdGeJkvJLe6m5rUuzyfM0Tdm8O/osQi75IMTFZxd8mbQvmK6nXDhKzqjUcd9
pCeW5SuG3vhGkPPAYaKwWukf6uXI+uAU3tXMQNO5T1o78dEcZ6endC84MqMX
AWMrIAagcP802Ks79/mCs5lmtvjenZprGi3r15RfZNGxPQD/fL493EAujCuQ
CYWS/LeCbRM44pNbx/VvcVqUNactbiyKebCgP9H9pWhFjLfYstVwCK2O/ria
q+6gfTYReVotRzoEoDk1hwXHGEzF0jRkDd26bInZQKF2V/cii1oMA2niOECS
wHxmV0lQBQ0+j+st6YU/nVVZlwWvDTpmqPeJURwpSLTrhsldIi7pNpRGem1M
5+SgsSz/NLStd1OjZPrMor14ACJXaJYehSzm6oM8MIxU9UmMDBbjunsKwgVH
+mPwHRzQ5LYnnk++EkPvm7MDegLP6oOun+3bZEV0eGmA+RPShBvCH95ZK6rS
0yYeWianHSD2v1hGapkzcMTuA1kBuEkyVbi08IhgDmm6dGxCREqX9yo7AQw5
kgWt4Qh5EUAmYFXLoUe8Za+r4yJNus46H2uOIHcTF1fkBK72yITZDh7nvWCA
gEGgIY5KnkBtZUyqTs+gG1hvGQ9hDLnfY89aWf9mdh0IPb8XM8EwJeufePQu
cfwPgiab6WFbh12wrqlyFphKd4M8ZTQOsUibUJELu/JyBF8r4rS55lts6Bxn
xWx1yU3Ikx9n4RYjJAje7ADEHU/V+1EyF80hvvEBeoE9mFXguf1OOy/WL9/z
ZosB3MQbv6UxmqNCkAvU/2Str4AR3Eyzm5gHLJADJt/1W0iBgACbKOEkpzz+
qFkRsOaTl7KQqVOAoEZUi2KjZjZN4HQVLWBSGSSUD0DZaSUifUfxY/zsjWIW
gZzzDQIU23aTiCKei3h70mIkmsUMeJnOL2ZzWAE0BhjASTQA+ZJ5NR24wi5g
CwjWXVnq64NRmxmfpdPCOJncRG/lCGjZULOOpPSw9UzULJqS7ZP2MfXJgwCg
N1x34IWeDvMHbZjyRmcDp/gVCP3iE2XtVJIkAzlPOgUnfmr2jJCU7Ea+vojQ
P2n+YCALjlWTVBzntlcjeiZg/yoUotImKX0KLTGJP+gP5OmKRxW8RDJDXijm
LgEuha6aReQm8lVtx4esV0pYAflgxRqH6EMQ4agp9WGsAUMonu+3mDx/Tx4q
6lLFKwzhO5tjZcG9CuX6E5pOUR+ocsl5hh0AHaLCz1h8YLPq/++tqvvXW9IS
EDthtBMaDWfGMDsptM0IxVtWtK8/BWdK3vQOUwcy00aRY/JOjbSNNSrepnnb
Wj/a+bQYkQpV5RTGoYMAcGrj+LUO2xY+05JNErkQHXFi4ym92tatIBtBMeUT
C8bOdR4IwlpAF/QCRZRMvq+r0ckxwq9dzjlWx+5seoudrtFHczgs7580+BNM
LXsG4qvTGEBEcqCbkAoNh8Pzn8Srj5/QH8ihGAGpKY+reizvS87VWvMoHyNx
c9vy4xHLwDDP9ADr3WX1wGJRygrMpaA9pywN0V2C/fdzyWalH+iFzHbMI7F2
B7G9wdW+K9vDhiYXAtm1ZfiwEBCWbjxkpCHeY06DuI2S51cLl028wlAdSOeU
oymavjEoVq/97oMP2yePX640SrWjG1+kcPiPpjGuK4Zpl14GKgQcm6VL6xdJ
P5SQrRl+oy+HP6fixG2ZL2u9fHAGuyYHbzfef+HCyJ8G5/Hml/qkFNPVpXcL
+2FCmJD/yA/Cd51Lc33aKFoCv1a3hBg9vSQR5o0gLVh42sH2jO5wQK8efmK8
+h1b7MdtI3cvJCZAJ8GWvpYxSTPvcPppSOoq9UtTr4xtlrjOWdJe1LIlmmZ2
eKQEP5u6naf+c7GuqheV3AuPBsEf6thCJNDj0thT9tKvSlDmDdvBAVpTICX5
VauZU/fngvVwuRwsJpt/smXhijk3J4STsjZeayVFj26pbM9x5J2NUXr2RLX5
mWGx4CLwkVlSrnnGsSmB3Gj8idzmUHY0pC/y6DcTw91IXG4/mZhVJQwLGG/8
779eDauM5LuXWdOmY7E6At0zeznZE7N2v/R8xTfVWMkrINDKL6qWWogTzJ3n
Uh2tNQn74uuzRoVhTRMFI0JkP8IM5IEINvkHXQgFs+IclTTQhcjWmBCA1pnE
zmkWGvP94CJBZBQB8H0xL/nWosbmN/PJJO1IEWSRF9P4yBZPp4GvUEDxHRcR
cVzoZXEH8EbuGuZmPHPwYW8BYs/bJ9xE2uRo1RoBrd0Cp2oSOr+3T3uhSxnU
4RuA3Z2MsaqoQICS068zR2p0M6jeGSIlNDaeVWxhC/mfhnjQL78n+IXfNZPj
rW5SgCi7JIwxBSIWPeGgUpPg1cPXkpFer7xvfmzx2K7DMkhM6A7A3HPcI4Gn
jU39adbQe20nY7ClmJPIZSYL4pjjjI7XjadZWfWLV/PckuIvQA8S44BAXid2
HlRJaH4G1DthM09umdpyEwmJ6nei8A+49AtDOCQRfI0tFsO2NqyBi3cJKb9M
T+XcfW5DCBP+0j/fS08Bh6kItxggsyAkhf0lrxFApBmaMrV15HAj5GyAxMqU
cSixZJpFiF+iEPuFLgEydCjVNV7C68Rq13hUh6nxvAG6gZw0iN+mtLo4eP9m
v9FXC9HD5emFhL5b5LLggRfXsvHB9Mk7tjuu6/yam7ap7cvIuOt7rbtWg8TI
4I6fWuQ1epGnRDHbgshsxUM+aqL2aSSkQSbN5Ig2VKemcigsbrr65aJV7xPk
TQr230IsrVzKI0w1elupR1qC8zUcFlZVs1FI8kPRQk2CAuCR+O7aQhOIp5/b
ecKCD25y0HO/+amJeD4tp5SYkJIMVHvtJWiy7BLXd6xHaDVOQSGNEkkWW6XE
IsW5xyn2zumGCl/3YNzGKGesrFA0J9hodpHUZEeydMTHkx+9YGvesFspfjmn
rXpm84JAsCtk+7SIvrwmEIpcPzltFZS/Ve/6rnVnrmTA28jIYuOn1VJjAYxS
KbpMzwf38BeRVCQjBIQ5e5nZ44t3bCNCZ23Z9Xc5UbW5FX1++ENw/YblY3Fe
VMrWZY1XVOP4jvMXFyLjBoRhMc69+PM9jK3ygc1W4binyDBKy1vGw5smOge1
VPkSvUXlHFsklXQOE1rF3aBUtQ+H9tzkXihTs9NLMvRVR0nCfOsDZJC4HGiC
ki3q27eeBRuyEszIZ7G+4Du0Zb4pXuOwR4TScfpBPwtM4gz6nA6Elpad4Gn/
yqTrMVgiMauwjlF3hsYMc3/GTnyBQh8wudI0UBBUfuP3XLnWl+FnaWC/SL5q
3x1ns0hS+yOk1q1tJTdmI7f0eWCq4COFW6aqGIn0azcX5mVumcNESAhyjpmS
HoxFwXpTNx0bzcmR8yVsfBNzJ9hpz/XekiuZ1Tx/6DDgK7NyquYBswLE3STE
aAJFc3irR3WpVfmDGbmrNWirPEYJ2+V/eB0kxFzhrcelompTpvHkK+BNzQ+8
UCa/EOjNjTHIPsozi8uWJl1kYgGaETJod9kCvVh4jmKWl8FGTRSq6oRFuUO+
IFiOb6bK8jnedpdlCJrwBtxdX1Q8jNhRZv+CQJzVgiM6F7yX06NeSlUoQOC8
xmXThW9E7iC/+t+h9WiqUyEnOPIJUAkkuH4foPt5ibLptKhgJwnLODu1TGCG
yRJVT2CJsdKOMtM4G2Ky/+iIiML6C6OmdOGUcDd2uGwZ4A+rXVzKnav9So3c
BL9RA914gn+ZjZuddTqOiMKluhllTvSHQMscj4ypJOou41Db8VaJ64ozRMoK
RlAqXOC5iT9cKAzBrfCH4TSpHNOiHzPyv3TeROVH4yiQR41w0JDi3JAQlbGu
TbJ0ExWGOu+Tp/jUAUfxZU3kluQ/jxp9BRT3aZ2T5JVd+QtjDv3/cv/A6PKz
BfawCsTv4PkZ+I8ycV2k5niRIegzLe+ltbdc9wRlDUoJWvmhWG0bVCVbOP8u
hmoGD5nCfr9Tntgxcngs3Kg/YHNUMVgKeEaFmPQxJlxUV6E199/uEWIEh8yO
C6tfPCcF8nEhnazJiOybfyOLP9WjlRTFtpBTl++ZzkKVBNw8c/e9MRXm7HCM
5XrLhIE7kbIhxhW37oZ2efj/Hyl7cWWQV4Guo58V30qXrcMHqVBhf0DpcCNm
sdrBZZUNz0i2KrlYVNW2iLamNHlzohBXBDnR2STjtYJaneaZGkfhRL5Nk9d2
WuE9+Kkb+hCAzIOc2OJ0umdu8uQ+9hVi3wkDR1yRKiinZ0GeWz5kpLvr4CNN
nbPrArQtazg5bDBPnHsruFSmHpL3PN+uRCwqGNNg7iFLSWg4guKOoCEOkKew
ZK8sF/nyME9Ksapegzsf9Tt/t2OPAYC+PfoEnDjEsskQ+MUUu+Y8UDzqmp7P
RuQHrQW+1jYgzezzagnL6ON0wuRj6ZRd+Ip4wjr+KYq4LSx/KnJRK2cxsJpw
eAchBuyw8Xd7VI6t2cmx0srrey+ODC2N+NnkpXT6oEItv/ngaWak76vulEgj
Sg9FCi3NdRsMbTYP7oF+bpuQJkd2ujHX9I1PJ+w5cIGUUC5k/6aw1rUSZak4
E7QOs3bSxgz+eVoS4wKJOWz23KGEVUZhefGgGd9jEeFhyJ0g8Er9nTuve0Tw
R0JSd1MoNfUF0pdgs02BlRCkgco9bS45P3DJmSD++l5HcO94gDA55KH0t+kA
uWaAecZNQnjPOab8EJlEGNcPiBhWNkHAPmRpjZaoXspGdrd2sEtQrmuqxSjt
xZCm81metROCBFxcnxu2aN7TFaxIJRjkqK1xDUIHlNJ1QP8J7ohvC1HP8YLv
uoPGYP5EVLGsSscdcj9SD5QilFyDAfOHmXGzDn1tLEqEMiYMhN1zIYphS03e
wnACNMfGSjMTw1pBRV+7ePGNpl43/ghzZm+qxDR52dbVlzqirPIh/6amFdyg
XGKNj5EDDvhC4EiZ1YoncyrHJ08P+4VWkfy9AfOL0QvGS9L5Kovx09t+ooLT
YBls52M4OszNpnRnecBNqwPi+w3cJ2JrqsDNh9m6nIBmnMMhGbRFmf/JejMS
cr4kEjmB/NhoiLkQnfDcoaP57PMJG96SdN+1ghU4GU1c0DcY0cq0H8sF8RXe
l3b5oJhIzgAB3vi81I70a6pqVSlt8GDNSeLizHP104Yo/07G4ggo8rZJD0vZ
YxWpOpSNa8U6joyO2R6AmJwfCK/MPw9jCBi82ndjulH9DhUcK6wko72Jwte2
x+QluM/Igsj+Sblf8UphVG1FTfq4MSG8P5YOqXEtIAx0USR65V/NlWce/9us
694p9LuXqbtJ8MmXivdwEXlSgwZB4eqYNmiw5mqnCjOOcq57Sw4Ztqkp7MRN
rwBsSKtRYWPC1RT3q9OOPsp65DiNihKQmxfOQ0LtRl5r+wENtI0TC3OhElOt
uTa+UyYZRLNkos5NRYOJ9Bo0UBYAei/ZArOrHRcsceFkU5TFVcTG8FK2N6iA
8mbh05ENfftU2HnfTa5hY7mcEMUxDQ4KLWqyosk32MkFn1d0+DvE24EXp6Ge
bvfPVmqcbBsj4z6AUv0un3/UR16TP9hi/Diz/2I3hSyTOcRf8W2G7i/tFjPI
HOxIO4M/y15ze4pvPjGY7aT0RRqbT+pW/wcsQwwG2ZMp7DZmbGHaFj42yq4e
jGRfChufSCW6TpSIecQPnyeA+7eDQrSYbTtCT/JVoke4Y6pAmdqRzrKifR19
Kh7ddQjKq/WWPawhRoLVUEjAWfNQ21EEbfRgonLEBBtJgMTr1ObfoKK0CQTz
nfSzDy2R7OKkPerFJTrZdv5DdvLNeYMEP6AjnVzMxvflWP1D6p85kL9/OSBU
lYu3rAezql93XdAlBOUUBMBOHI92QYVt3o+id9TuWwDvWn+5F6bXgsqM9ZMw
vRXGa25Ev0vDY/Dz77N34maaB+QFqae+EXkbIk22NRALZX917jM6v+EQdfI+
kx1BRm2sWzOKImwuhFlBLtGB/6+8NRnbkvNJ5W8R2sXE06PCUpJsjm60FiOP
D16amKx1BVorLuJN30WIH/v1bDILzcTgRLjoljDEU9DKymHQcByD6NZf1kc2
xES7LyT9GEYrob+DRVUTffgIgeL0PgVK7+KRMloAEcrCXnkmXKX3kCJGgq5V
aBO5KRcd9Pq23Kt4y6QPxAVCZBBAY4ODC9T3akgszCYswd6NjrUIvD+GkB6B
XWALmdkjmzL8oCgC/MMySMXssmxiCbU17zHylsgbB9UL/OHMsyFUtMa1/Zzx
WcXZgGNG4HpwX+DrLnZWK2zrEUXVCXbbpoKfOzrCxqCyiY3X+o5ISUYZInlZ
VGYiiPpYgBGqe/rRCD3MCT7X1x9Rv63N8KAIIFdXyEje9/B/fN2B3hy3vqbD
NiwsQKn7CEcQ8IIMBlzcYna6sKOTJWw7UE15QAe5wUb5PhQfHKeudvy0Qq3k
yNl6xTCnsDcT9M88XqGz5CFWh1tRJgF0M5X78r4KOQvnL66yRF6Qz6CeJU+J
orhJarwk3g5coHhM42+fsIPlpERRefEHzs9f2et8HDeSV+/OESlJp8O8hqnX
L2IHKLcPRFI4/3AW2aEla/FfMX3dxzkDp29xAvgF+cDm9V8CRSagFvmp/81h
NZFBBGGMpRI80TGnTUBJFETmlieFIEFf0j9c5ZVxfF5aj9TXcI107WlZ9B4c
T+WrZ4tTvHsLGkgdzJZ7jUpG+i41It/7l7l8DFujezlWEyl75tm7oyPvUyWf
1HXwz//cz9TKmFshOS8z7Atw8L8K6XVZZtYM4O4AFkVaAUIacceyUOLN1Vx/
shA51IMcHXSUm5tLc1+Abg6HQewB1rSzV2ioCSlhYE7IjPuEAqSUQ4WXkaNz
BSGplg/rjBlFJktZ/MXWOReG4Cl7dx1A5S4xUVaomJXntwkHv8QMZFS8zn/4
Bxs6UPChPXPIuCHPF+/G/6fuR+FkcbyYbMKE1VyW2Pu3ctE3HcOE8WyUeraF
dSNqp+xBgaf4ml5GLBsm6lefFlqcgqx39nQIpkPvJjzrs9vVjfZSpiPM/QGd
gQc+3cjjRc0fH8IMrkS37Sg3g6kkHWk638I+zYlV1id+fmAJ+DEKn6dDImtF
gLU3H2SUZpuclrzCCggWwkrjycydc6+7a59l39Pwc4U0uddjSh62FgfD0p5b
qTypxLegDNkLJUJlQLlrgUM7sHGx5mCf2Euf6yP4n3B8WU1wWc1+WBCzRZKh
r5W+juXOofMWR0vOeD4q30LRas3kq7iFtW0+S/ZQgxHeFSfuRXBnKPJd4tTA
c4apWzIDIs7FGVFsBRn75iYVGMYaTx3tMXPEMg+48txH70BhPVu3U/ATdCIm
TW45Fw3pS97kGsAZ1y//3mwqMj/bXP5FXvQX4uoycGpdg+OCvCbBZGXiCFzH
WPlJziJ2yjAJkjnEfuNS6P4e0o4vb/4KncY7OxgmTR71pJhp3G1gA80uV3e5
0fyJX2TUkeySieBFdS1QVEzOXEEmIpi8oYxHr0LKtyBOmHSj/XyI6jsEfMCN
BnqwVIapk+qS1hIQwbpfG/J8ZslYqIGBd/Kr0+eMvARfCnu6aMiIKaSkt3JW
/w8Cm/5W7aINigqKDfK1giWF0Qav9wF0nqaLrqtmza/pCoFLGOdMPbJCoSla
oDLoh2waPvjxpkp8/tV8m6/niTNKOPR4cTuieSupYwnqZd1TMUKrW5xvy3v3
Y3jb6ghMtNDMPjnZplEbTOzkSgL7LPox/G7yrnuTP3fVaIRaiEuZReuIukh3
oNeimT+kG4aV9s/fgklRMm4WXX9MYQ1hkxEmvT8oockpwKktnZsQzH1wZDQx
dZd9PdtAMvzqXvBA2NMrs1ze7gdJRupeTFTiuajG8mNV0ZtJO94ooLab1Vpi
nV27uxSkHcDKL7GheITVos3cSRhCH3ByL96IFWMUxeBKnt1AFv67GF+B3Nci
A/dBwR4TnJ8vfNZQHb97Uff0z/p0DfvVTp4GDdTC52zXa7e6NdLDEaZvI/lx
HebKbP6ZMh3asnKQW3KyisVqfI0+8BN7QBUJ4cR5O9eXRegJMO0mGVk6F/AL
5IeKMo3zprg+jqeFzCenljHVpiv3Qi6kaVPA+d7PtnyO+pKsbJjCoAamKpld
y/SoY1iVCq77CZ4f1+oXXj9vlyLI05fCHmgu7hCMGnSbc7g1K0fHQHqU/jhH
P144GihkrbNcQMAR2J6/CXnH3FurpeqOeNbfaJy/7d3x+Ms1GVYdHYxPyYt6
uUUwxEwvwraStSCQngqxDmivPHC+X8Jcv3AmkEudwfI2/Mpf5tdKuPH1xB8l
9UWyrXhfkHNRd0U71Lo2mwUeMvo0n1PDof4vvaXuqiisKiYL9MzKXuRHH3W4
fTYZ3mftrzXN6MrBMme6jtFigBhAs1uMewFQPwkwWCON/zctHK/nuWbPRBms
kuT+DW/h7EMJacCQS/SnGWJpqUiLN5pqVPgSefTwVcr0TanRwBtr6XT06pVf
MnKIwJcnDnd6j5YbZmZ3lYz9n8lGtFdvkTIYz3nzDMZYCIfgwmLaPk35Jbtn
4rH5pV3DFWnCEpX3cH4T7gYb1QiS2OExPRP2z9D9naoZFpdHdU+54Kna/C9Q
jWDmt+OnDBLJxB57yyPA2JeAjqRwK7E++fD6bAwhJrQhIhzJ1t55e8wO5IXH
FmMJX2u2fyVJ8Tf3cNWggAj9aZre6h6T3iSSgRlwtHMq5yhA3hS4YjniZqWp
/+TV3dUnGQ0mAbz9+03bqhJ7qKJZMy7butEj6drX+HCbXs3pN/USTuBqRgr+
iOczwfIeIhqXNJo70alCYqklnbC+czhL43bPmbho6QH70ZYiHWTyVMmcAkr8
hRVxGlo5T6ySkKlAuFYbko87oge4VID7AWWvf2pdYujYNLLD2SItqDXI7LJy
U6GFz10aRkGP68TWogQ6FhJ81uQTFhwWO6a5PzlOjTTMEZowrbdD14OfDrnY
JOjoYEtwEMvN9BTn0E0XTIOXyuQ8SAJyLgaGO1OCqueBtW4gBONEQ8qsWAkI
ay9wbCCjhSw2SuiI2qhcaHujQ9LeA+s44J2tHj1/Egnva7DYv00yIX/NBC7Q
QC4pBHN3VsIS02S1wA4mhANqXDdvRoHqH7zJNUJGInq8XlCR1zuKcJNT0fIr
gCkTmd+L7PtR/8YBOxbYcGBYBz1EOqf1x1a6CwwwQnLWdjZq34jLJ6pN3n9s
GH2w5AMKrf+Rm3ZE3Or37StDDCUMI1IGXGGhRWAV27UN8dV/jWDGNSiLYNBj
NQf2o9GhDMIRVE01ORaB+0MlU8kH2qLTHYSIJDMqM3fmwDrQaM8WEINTOwkq
PPXFP23/2jASLoz6w6ypnXOCJD3NhXCKcLhGhGfoFXp1Zqj5dC/bULHizq99
FRz7pltlmTcIcJ52+gKERSEg7g7ARBp2tNVCQwLbxE0PQz/qM1q4iQ6eXtm7
RzORqWaoE4l/dH4+yy89KDzVyP9uX/9XQ722ozbF459B4OSkkQkKjXo8RreK
Rjna59iQAhhIC0rAsjcPUCXB6zI8OSvmEDPv57ncsrcOn5szg6h76eemwgN3
xJWh7mvpbglqvP+BJUljSZdmjs9uooYkeCg8tSExPWCgsZPTEPjWjO3DykHv
fVcq1WJVqeCc9qMSW4/6UD4QO9ERIsOFifOQgPtQRq02qq2TRJ+/Fl3olhac
bFE1nKKaQV5iPf47Nbtsot3lKkvEI8b/bWviUc2X0/jgAjIBR8k/jLnuCvDG
9Ov1Wwbidgf5+egkJ9pcFcligFLYm2ZWz/GHF+al/xGZZaOh/mWOZQW5m6pu
zYZlESDLjeOqytXAG1YO2x0CUXSiIvUJz4WRu5cX2cAeC6nhcqHeL3VfNB1b
jXK6NEjIpei6uddEtkShAUIbbcEkJWkiHPXXs3FPkpCE8Zq0td90Gnrwjceb
h4xE/8v/IUlCtpLoYS8ShSNQ3Cv+p6Pxf2fRKRUdmp98/v+cMq4lAXbs8USm
Ckek4MQJ0vOz95ucgKfCuAYeLvT2AdwCZnpSj0pc/33o6AL19WBYuusx5LmB
/D941BIUYQJeCBOFiZmRViO65Ev4veI3wmPSgUV0tjSmi1UTCC5PulhiaDKm
eLq2oIKt57JQRPC+XpEO63U0Vlu0U63RsMmcsZ+6Ne18cGdr5YaPzFZfZUsX
hMqQ09dbJQc0vZPZbC2esf4s7NRa3DYrKJ/pVzctdHTtJ2GJrH0NCVX3wmup
4fqUniaB9xipgDX4mVb0QMqnFMUZ1+rtTBQ1rZ/I2Ze1fwUGusveu/KJuNiZ
oTkOilcvzJV8piJyFjNHCm8fXydgkKLZajxjA60DRhH0XsEFaHNAl1o2Ak0+
Vop81Om7ZpyvRyNfrzwlrLCpvWnBAwLl3OH6MgT+2Gi6Dlq9ETbEQ3L7NVU4
rNDyR7jAzY5ehU5DTfLKf7Qe4odMePvNpsUV+rsrK4IcSEnhof1G3UCQcsSF
yxqGXBIsoWdn8bRrRQv7XQFpmZrzN5SvZtMzOQJi1iteqCbRXRNowc5G131c
2UxE8y+k0+oeCmSNImjOXV1GY6fXBEj/7k+Je0pHhMl26lUFrdguf9v34tFg
4qTkdXV9v6c7W/Eh/76ZjV+RjkRYW58fXJrYA16UwJ1ZCjDgMN20W9EHLtPQ
Lkvn6CrJ7q7dU8XiEbFMVxxcZSnJePr1NHemf+nTjvSSWNzWVkZ7f0LSMmla
nMz2N+mY2+2hjTmNnwYJtjDiVW2dUppptlILzFhJG7yLKUhnAIysfTf9xv3p
5pA/xDdKZvYsNTOHQuoQGO2Z8uF2FK17SazxpUNfbHjMW2xMgVck+oyHvlI+
vzEYaTHR1Zy8mJ2ALbsJLRAcxOsfGdQ+y+FMYhevTzqE+r/cyJWXXNCcI7wj
mws7mzu1YmZWs9pPZkU6fQQwlVjiFE93RX8ZfMF+09tHoROgeRGF9yTqL++D
RP8oxyhLWYBhL7z/MGM15OUuO4hjK5A2ox8bnVy1iIYqKVaMl3MPTrifLRo/
IfpocakNvSxBD+F5eb2h/u0mpLj3j8Xvjd2osWh1+ApaYrIKmIRZNb9ksqMA
gnnGcrIwYxnmsr2LgBVkcPjq/OIoGdqOulQZ7aJbHGbpWR6c94CVAw5B28CG
F+2oiifYnw8Hlv6Z9UNCacjH06I8hKaTXA/yahcxr036jsHFqLBscbUq/Zn0
SRRAqWFhcZmOEJrM9YlR7kLXWLNtYP0Y356NWP35slsi9hQY3pLmj/08Bp9y
LLvdTsXV5AF4erXpyS+rwQ/MocwUyuMdSImBrkqshnkdsALREpfcGLU4md3H
wwwLCokl0DDTOUl4I62Euj4MmnKKAREKcahDiME7x+KmHiEgh+9G7WC3IlPi
BWXMAbRW1T+uGrFc5H2uGL26gjpSTQ7CXVnBqS2SlY3w97dOIObOXLjOsbmy
CSa0rAguTi8I9N40VGZWqFWzlCZ6PzTRnlKL/zXfBypJjX9QOloDyhre5/m6
PxjMKphMF76zO6gMhR4Qzkv0J9OwhIc19/NuortZ7lqLsBsttIGN8mePRLY9
wZzEe6MMVZsfndYnrKTUlWtljK1BdR9iAJdhBgQMZheVnNZeRHom6TufWFVn
orzr361PfTY95VxaozZ2H61gPKE2dTKeHCF4X+hfGK6mLh4wCcSIICDAnvX1
mG+xsoNh1kYbScw7i4H/+asOg2wVu2gECH5vpJzWAmL0aeST/FsEP4AnZQIC
sP06pDWqMGw0RemCt8gq63APIHsKhZB8eBzp/9A3nA6X1SqGbsQwHXnrLZKi
T7QLdSAq07Ka+6rjVJpNPPua1U1C1E54N/7jpmsg8L4cYXLVV+7pm8yP7/Ue
68x9aTBxTcfZ+6CijXE3QxeVPePF5khLBQrOPzBnyXdihdO940GYCZcwUfUK
jfoCYhshn5atlYF0uefisK351tMPOy/YT8TfBdAutKqmZI0OAH5ZjThHL71U
5ypE0jwST+GZwvDByWSBPcgbSgwySmxSXOdhnQPOxG8zjyKsuLIE/x5Jgw3V
505ePaykXOQr9bEISZAA53CtLvkzD0WfLrNZMIu2WW4Y+y8niLSy7Vhrh+xz
EOC6HFxlIIbRE/wEtMGhfiun+vSCSLemhjRrJD1DkD9A3aCwKo5L730n1lrT
aDoGf5EhvvspWH5d684T3zLUnWzNq3bL6xLcLvg33yVs+7rLbeTdsPbmu6+8
1AQLxWwY/bz4sGL3kiS6us5cdgUzi6haTZWImo/TUQ0JP31/tZwwhLS70FQT
yL0BFEOe5vHJTUWvhId6retOZ9xXEXbnU0GgTSZeMli2QdsCtNkDzruN/DNT
2nHjljAMZu/qnGlE8vauTxUKCCboeBctKuyjESMCLpUxakhIA8Vx6WdeKifq
qg45n/dXAVQE8fsaHLDXhsbFy6UfNG/BXmSYt1wM+swe+bQlJOTbfrg11DxL
61How6wKxWPVem9IgM9URIapoM+XMjU2VoVrF69riqMNwBENOXdhduFx/W79
pr1/Da2ipSbiORU2yoBopu44RQujmets7ucpb7pR9gQn2VeOQbccvrRMSjj1
kntdYZIpoiaO2wsfpuP4sTQavs6jES+RzMrOSaY4c80hZMD6RoEh61pAO5Tx
3t7KOadOKDsAxb8nW9YzNhYEg/gOYewxf6PWlw3heYcMxHxcFHVVE/eKQU1z
QGvd276ee8zWGWjOMB7EAU0LNQ2J0eipVb5RzNIE0+29JyFjPXFbNDJ/9ZrX
Rcd4/jlqb1FhrtraYh2U9YkyAhQhTwWpawOjogaHxMIGRUxGx8pGw2N8oXhz
Ps28QMnrgP539Ut2WtHsK236kJmGnUg94Cyo9KvdhBet3yavg2loG7POafzJ
1TxMzt9drwtCT3FGGD+2ir/fTdKs4df/j2gZyawtvkC+v+7xvZfP/II57HDA
ZFWN522Cl++JOY6v3D7LG3j4J75qP0btIaCtIAjpPwpsThiIPBINKPVx+p8f
7+wZZh809EPv2aU0Na259JLafHG4zyZVn04tFDqEWqhUPOHLxWZSUWVX7G8a
vGSSn2eoIWLYxyWavNagYbqlxcTKjfW+1d6M117jrrEYnELG/yUGAd0LHlcV
G5URgQOPpJlsyRp03eGUFs2lqLFHbtzSZWKn12SYB+TFsh0BcGsiD7V/xztM
rqWFPDYnKK7bGOXDw5aF54Agqf9b2NkDt5yQ6uGcLTKomOfk8WxVT8QSQxVb
Ffs0MZ54/w82gBjbqrO7eHZ66RimvMGSLWxQulru4BCuzFKP41vtOfFgXpOg
9o+NgPEBC0Asxy+4jAaced1KJHhvgLoGK9uf5dhXSMQb9fGWzzkYHhq79vNM
IRKtOrS91PN8gNrBfBup6tf5JgNK2klJ+pnObUptAPCuRXMGPgO7LU9Q2gtG
EEJRaRu+jkC7ufuYn/rE6e83sBWg53wGUgkms2Mk6enj6WlrOB63sigIoXnh
nUVe2avkLAkBfuWnbGN39hH/58v2zlGvc5QA4oByDtj3vHTlPhSfH2S7MQRK
x2wL4yc+dtzcAHZqJ4Dh5ruautR25JmPfszH1jbKlr1YfMhUYvV5KJXJ5ZQO
55gr1ceqk2FaABD+eaZGCg92eiWUd6+ot+H2+clbM8Md4xg7QFQgmZE0WtvS
++UEyteGVXkukPBNLXKWtoSop3yv347DG2JrrbfZTQpOctDfKWdUDeMAMX+7
KCNfdhtwn2gc2jwkPNq8NUIkyL1bl++h1iVoJl/h4UvdxukAGmBmF5sTGXnj
0wmvfmoL32JysmEYn5sXx6mOWZGcstjLDis3BA2WYeGJQ7U0L6dlewftwhij
Q6kiUGkfI7F5EFFg/szp4OTeCbbKhd8NbAeMZPRtErujabpdWMVM5gPREFhJ
HQTDiH4totL3JxTLoJg0EPPmiW51gbmZFlkLicb70UZEE9pgtQ3+/PUAhkVT
TufvBI9YCRYUfBFxX1QBBnRVNv0UaiJPLvXTIE85Dzg5osPD6bpcV/0AW2zH
n16j5tNIgLNGwoaSSquHDF3r5E1QLwZY7W2PdFO+tMZBFf1FrLbeXMrtjsMY
vggx1MU65Joktxu9pokOk2hRl8qEcHev/5mM8PnoMHbcxerju8tpxw03ONvy
aaH98kk3tZ4DVBBJ2YdTR5/83CLKkvWF9fFAJu5wV85OhGyKroPzDxdhXbZG
8g2R2RaHFor33rSS2iVZ57LnHODX0pOuL8vRvvK/qh4+Sq0AML+uTnzB9vpo
5HDp5k8RxXqTCCXp1H4yEUGNRci0tn6HTw4DVhTiz+0tYRBuXkHPnZLfmycr
1F8JwHCHpYiWISR//JgALH/pkqH9Tgk745f6VQFp8N61mfjz8CVRFHa3/06D
GjJHEi915I1d5bKOQiuEXGvkH5LgJ+x5kA3L30TzJQolLWoEAjXLCyynl/bE
XYLfU5ePSKssxU3DmSc6DJHypfYI7RkVAnz8S8b0o01THaJhM7x4NoJnxzLI
obPMLFNU3Jwc2iD0qIzgOZLeg8cQ/ohv5noDfT+mH0EDC5DWTGCCopSzCxEF
v8xTYSzDqsNE0aIpwCUFALFYO4l9b1iBValee6JguuqHF2F3LVwEhiNcIidl
Ys7UCr/lMoJIhV+2vTBbLIc50lFLeEUY30WjHYaGEe8PRtYxoLuwFrhMvuvn
hjICvDHh9ropuHwHfcJjWqznFwpI/heWMms0uNN704BT+Ypu3TfYAraTcgFe
FEZagSHK/IRLUUtepKGHIn1aQyTP55VYLEp5VvzQcX32Jv7zREmPIu9/731+
Zi0/yA9qEPRLXcgh/E6fFHPC/vxwb8HjMMuWdTPJjo37oUibATIHsh968+kE
qVNd9KOYdRzOrIxL+9LbxHWHTxNMD2Vf8bc4VthsEhQk/HnlL/AN9JMAEw/Q
Q3P0xZM14SEAeLEe8r9FkrLf51vfFBVXPFVACP8ofIvuRR1xUPX2SqegDJuy
Koo52BUWXweXNrxLdOnZFZjPrVQmCfZAxzaNNisx5I9yO3Emr3G4Z8WZUtmE
HrPKQpNwbpcRU0NGa3WkXnd2Kw6fTL5PmpVn2UYPmgh/sFS10xAEcHETx2ok
HuCzaArCRYXpYRQI5EyrB8H77XjZXTPukgbBmM0qtJh5Bcea+z6wysr2zEqW
dCl4+hq45EG/hHuNj8+4cDdmxLAXcZw6sVnrfUiyPOcFTCh4vP99pMGlkyMS
9u3fmfx+HpPToBN+ubWinGlU0xNA1XOzOWVH/LrxXfq0wW+3umQ0L+/U/4mH
IIdgtDyr0qAMJ+ZmShgYRwbcbsYKYdj5qPyKn5dSflm+XOCRYvTNeIWnFvG9
7UatbPHnOu/clGRRRYnemluVgycgw/SY1AnQWP00jrhlD4faSMJ39fOpd6g9
QYGoR8y0fM5rPMqi0wOuur+6t6iUM90mwhLwFXD6xwxmw9bXincqnM4pfhCA
AEo3ETQxhmJvCIoP4d8dJHXbgJY9ASBpYBJKRRTo4iMi1/nrbVrqd6Do+6CO
+DZr9WTeDiImmsO4nDA/0sBNhdI8QTNGRJ6EaVYhYZutL8AVUcpxl2/0IYys
UZiyIkQB4gvgl1SzH6Fn1WZEhs1vxqPAkQd7MlwlU6uIdyxuYiF50gVRbCFW
5d333mPmWCCOHrYrrZ4JPIYdgWSMo7o8QFPL4zxoQSoAUuTBuDukvKSPIKjx
GaJp8LQs8vnOZyReSmFRsQcLGjMQWp/GIbwf3RvqgNBnrXrf9R46Bl6b0SUU
LqSU9gA0CGT+4odb0UL7ntB3XDu8uo0NR4leIrB4zn1tRaF2ttrlW8gGEP54
+jEaZhn00S2HrrDO2ky3ZZD5o9XdNToEBi6X+usIhUCcIr2GigImOJz48xL+
UWe4uAb3UAPbUQ5+Pni11f+ZxFR7EPzHFEVwGi8GpRUSqkUzXoxfAgspVa6o
OhNuR57niO5PTQVQ9ngT2juLcX4BZc00XrH9iqLDtrl8RWvw9MfxYgx7uwcB
SdbhMkPRf+teNUCUyeieV7bGf4d3T11f/uHfXgImCBWsMwVDd+X1MfmAju4O
nNSKrEFbp+NewlSTFgFxRKbtDUks5H7vQwOxsCAVK9Notc9y5XINdZqa+en4
Rm55qDPTTaj/wKEeXCgPuPDuhbhYHRsmtOhhzDy6CR5R+VqBb8Gn4n8BiLVR
VS45CabMo+21AMNK0hRChBmYxyoTe4A12H2UHQ3Y512uc2uW8+22MAjl5ThZ
B+lrR3XBvt8gagH/tSAOnJOQnMZtJ4cWv+HOfO+airljFW3ovLDtZ1k2HXZ1
9mw1zf3SnLKlYHqUPraZVxjckAvPMkD/JtJzXiwZ77JnQ7bDiRnLK7O/ElhL
/gqXqSR6PhDRnZhRj+nT+em5rpzawHf/i/oxW2yno7Y+5YaRNAN3MYP8FVhu
qUk8yd7eLG/6XYmBMHmwPvCiU+5ArbQ0651NVuqfZsc7SYzRcupDj0OD7mYd
d4jy5b1yPI51b1peDq2autFdwbFKMJ3LdTeJLwS/F4ymECZeoR4LcuUC0qHj
S/LhcVDK3hFllX9Mc6ZUda3Y20uFJx+ISSbEhBbPuwjpnohrrxLeKLNT2VSB
dSfqakUw/UCIkOE1GjWEycvnQb+j9wqrgym90/g+vVy5e0D4hks5DMeNKUOR
+PLmpN3xc1KdMUnfmhmtZtrZulZs4caoNMMpnps8frim0BqqzQQbjo5habm4
NhC5XzNG2cO73Re4Punr3pd1iazsr5H5DDjFmtVrKcgupgKFTBVPJrridUNw
9PLTkBSqSiI8KjHre6og52BnCxKtAnb0LIj9fdVbi2u1ZFoCPEFRBB5ed6or
fsvfeHuuH15e2pxdK8S+kMCKj4CizZlVJykSR74oWDkqqjFjm+WnUkfdxA+d
l342uj5Maw2ooq9zxfU2js5o5LK3syftDfor66KvTLQ+N3IHRmXc0hFHQtoM
3zyr35d7erY9ol6TZnf6n1cMcOrBBMJn0zWsoy44H5GCw7RXHt8UM8a5WCCd
ghLMzkKHKgMY/nr8M/LC/kVW4vd6uwYygppnfqp0CHrlirkzzY+f/qyaE1S1
ZmyxAktiRRe7D5mkqXVmPirvyvnDyzuzhPGoT5D16ZWmvwizH2JZon9Hfz8G
AFrVPQEU15rPCfQt+atWcPf57kRTKtipN/WP4WqNqQBLdW/1HEi5exw/ItcW
Db2wIyDe6kqSi77Yzo8f2/5VA9G4gzWnqZUlipdRe2wMoiWdOnzH/bKeK8cL
/xXxDZJXFrXcU0VaiNu8eXWOC04SFvyTNikQk0t+MdXjhvtR5qsssfCzalZG
r4rONGlzJ9pM6gkhI1tdX1fXwL3Ov8BriwA67TFghcRgDSfru+Z187INxP2s
wbZQyhsRKvX0g2YgvM+TkSa1xxJLui6QBo1wFqhF2XAgTBVLhvNPlbCRLCz0
wirZ1V4JL2j5brWPFwrE14flfCPs8A3PaYGWeXTfE3al3WQDJ21RtLDSdIpO
ssVzgLm5p8ESmSHZ752yQC/QVLD2Qf00N8tGOf/kRKHl6gB68XEWzis+CP0U
ah9LHIXcVT7CWY6uQXb7Qz+wQMqCsfyH+ekNDmyMF1c3RbcRg6Ou+W5QuF8p
uvRcYU1Nj3jpHotTe1sCZGM3nQ4JfiD6CC/LdF2kafunC0BYuwf2jTlyo/tl
G68Z66SmTzgXgPN6EEvLrnTTbvWVZfcbsTewtzuv5EHKsjTs70vxhdk49rle
ANnv/bSRAQ3vXJWEY1lKdKAA5n8YwmOGMGj6hDO1vJIlwLJa5IK2MdnTclq/
EW1h3kuX+qxKBVkMjO+HtAwVMee3aNMNO3wkV0jhixDEVPI3n6s8xP58NwCS
PDiEe8w5hKOuU6cQbEBnfIxAJexeIBxQu8VCds6CrpjmDIYYAVpIB+yobofX
hQtLjstv3QwmnrKJnM5Wnxet6XG8mviO4neCs+sF0n0rk+AzPuz8UmnE4JXp
CWag/st7a3bZciUZx1ONrGZJ8uh1jY4lZ9QtRKXER1bE6K44mdCX7HJOTTeh
BjLt9KfghGV4i4gLYMnQUh6E6j23McaO18pot5LxnYo8tSBGuSzqvuOd7eiy
sm72AVSdwKwDLrde7vOmiAJkLIqJIyl4S1xhi6UwXJg1f2hj4n6e8/n4O8ej
L5fqt/ElzpSYoCRHuQwnY6pAK3AwkBXP9wF4N7giRqasFZFl+DX6ou7PE4hY
KzDpXUR4paBganD7qoBTvVZ3d8PdhtbLsLQca8WksRO6H+N7PeBfh5JmvXEc
d8LVuoKkXOok4L6Qpa5TlzXXAsS3peo6bLwii7+yYzl0nfpamBYLR/nUHtYs
P+PndX9JAzB77CCQsEvFesy8cA8lclP+1b1/be7Jz47MAu8sXsL17GyTkkNf
pDpDMw6+HhEV7I+wYuwStQfzt/RWD4QhMESvrrzK5JG3lo9ncyg3Dkh0vj2o
deSs5Gz82lDlp+YoP4nxGIerVBLDTDP+psP9Q0JDs4VJRoy5dAGmuMsZgG0x
dh0eKaiGCQOasNXNwE7VTC4tg6HxEsdrS2Ibcdw8xFzxVZx16joARvH7uWah
LTRKhkYpssMIV2Sg9/bXwIitENlUGTjbeIK6XywYFIHItBjFX+2e/GGopw32
//iT1tahsoqmz3kdi/GzvRFZ/FdsE1QuTygjys8hx+PAzZZAodENWrcgCWwQ
QPKEgz+MlJQZqput9+q1cvie9tPJ1qDifvYj+cydVJvyu2joLO7I86OFxUs/
YEZqx2T3H9Pg8eBWBSER/ILg60QnZ+gR11fWWBMTUDd3q343juHkYLgMOasI
9lAkFOeJcA1O+q+lt7YBPWdmAykYBNPuSomjFbDhbcBXixHnKtPCJGXMEGDi
lKqK7gcCrVD86F8kuyKZJEL9ZTkRoLY+fOuiNjCMJpk4RJhk7vVHYrUQLIFW
SqDJHkRF93p1VgnIfogombKEjae05t4D5gURjkdhZ4fSi0hXEQ+TVGMO15qc
ylDGbHdQk9IwYG+0ABtsH6mJmZ0o2Pgaoi18enIbieNa/jSA0QjgvYtlGogr
Vwl0gcYbsXir/i6UJQfi/Wuf/i8dQOBNae0iE2STS3ASYU2aSR+MLszXgE6W
JeUhAXFZx28KfHVouWRf7svfT1AnDBnEiYCgesQoSYYBJshMmt6oAg4us1Zp
u7E8XupPF/QGapXACy/YxvXqU0WJ8hy9cIikZCk+jlFblnu0mjxZPqKOLHhm
VDRnFa6KgT5W6tbtpO3t6jNIqVhCNWW13gw938dQgWULoOguLQdAK0NFvKB4
bRg6JCrwxHnOsnuSSQc0cU3MTxb+BABGYpgZWy5/W5lwqC1+6AWQ9v46DaDn
3XY3ioV3VJKkZCONnUKfAYSJgdtTQ5VtyBKLAtEJH5oXmC/FRBVhGKQb8RAp
jOGduC44AFeIGkLBUUjpci9bOmS73UZZxuBQRLmoDx4JPfWj0e13lJ1HKXgy
Io2d5r2584U0zQqwHil0FSb0nnygoPtUdpKETsrNE68bc1z3DIJ8t0jvuaxY
Cci5tuqlR2fU0rGeqsAur4/n1Upo3SzEknKIE1vdOHqb/QbxVBAjJs8d/p8R
U9ue47rTdKXzk0UdqNjW7o8CPcrRlck9tkphv0aJa8aPH0c8tinPCSFqFH7h
cC+pssajle4Chcsg2f/Wba9uCVE68Z3YmH6C0GHfAk8249Dxj4evNfGHNjFY
4PFCOVLcCbctWod3dD8l1+LKeeA244jzkCyYM5T01X0tSySBxoa2acnos22r
Wa9vHViSgp20WI6rA51hrbwN/pdDij7GD5KHkqdRHUlCIsaPrNAQn4KcDUAB
ouD8RgbQg15fNi9D7D/9BJ6AIfVmLpkruPfMN6JNrHcVah70WVpp/0ABoMcx
N31k86+cO0SckYmxDwBJfRiIoZB020PJifAWhex0ZYPnQhFZ5QJR5MVPw4Db
wFSvKHZFFJEkjYoQ93b3N5gSD+tkumxw/T4iD4cd6pCRaWejoJXzl3MtUqwQ
j5r6BRPnDzr11ks69N5qjIk7mWF/hn8hEL8YoYEUQ3A+tPRYo7hTN4V6DbGZ
MXailqqig6Tj2hVjwF9jYt2F9Rl1YWQyQC2DQdqkvI2gAkLoA+32ga98qecl
PR2SR2wAvIDQrCVN8q1Kk3VOfH5X4/uknmjCBR0c3cpyS0GzsTu2xUFJ+qnb
Zcs1WUFn+Uzo1mMjKMemNXD9sjdmzQJ1e6SzO5Mc0e9HGfBNXA6GQfhFP20n
a2zXgBCIWRT6dImChCxUgahLDs3Z1YMscadQODGH74nhoqBYjCu7fZBzIQfb
zImVpj6PcQXUM4C6CyEQI1u6IsIZqe5kxjaFYobrj1F/8N62FmlQpX/NNBlR
kYHyZR8qb9QZolQpZo7+WuoJSKrlX0EaM2nayrK2N89sUSpGU8ukPFNqLtWU
Amt4anVNaGAGFoJ7FFGGYLo20O9X51bAR5YuEw2Tigtg5oSt9NWYnmzUNuoB
W0+brXMf7u1LZ46QDRqyeWWCRFX6iNvlN5Y04ldTfRlyPYhbiQ2+h8mMIps1
/RtSw9bwE8vXwg7mNQn2km81Ej/yjYi7kJXPWVPiXqK/2eDt9ylcgzOZdGtF
yx2EqtxHs6KNy1eUFwmU9i4p2sKHWdHPy4hlXyPapxHEOvOXUMJJ+OmEGJ//
9ich5EUyResjqJ7o+W/G7fEFHY51lGuEo2UtH/ntTTSVq8gChdX2/HZKjwIx
Qem2z17fNiRP4zDEseF9Xhor5NtrwlI9AsLfcUYfoAiLGxkcO8gJ5p3C5FoN
nnYZi9u8LyDgVP93mO3of0kjEQxfNOOh1GI/rdBi2JgAzhyBIFWjPaN6Uc43
FZ9vpvuroVbPOWrGFV4frAKYqxDx81o3iyTrnVILk9ek2f2tZKUYBzM3qojA
0G5ZEVKJ+4FyO+gmYgi7bIBg2Ti2iimWSbj9l2Sc7vDZG0jlFSavKPEr4mrG
ZpyhYh5ULfyKF4b0tAFPr8/b8J6p54hH0D+orzepiQPM5h/4D2up/GEwzSwd
0BwtHlx0+FXki3ubvDfb9s/SBqZ9Bfrh556Z4BREofrQYmKS39MBUxMR6UR1
P6MHXo5pto+/GOWwSuorEl7G2mKuygNplmKacha9+yt91Z12PFdUe7TZGCmH
ZLi51L3yNpEkvVDPpaLc+3BkChcePOFr2HFXxNEi8NCy2GZim8eGYreFSHrV
7yzAJ4Hb1evSaCjrBsbLqGRNhaoE3+XHglmVtnijri1ZgebrE191IjD/d0+Y
AGKtf8njuB2MtLzcFgT8v+1V8P6eSzvBKDLDqBIK1dqIycgeK4uDkJk7Shri
3YZeSu/z5PBjTQukbqFpB1oM4g2cFzjnyaF4bMt8zPwWLqGFwrtKh4fBRYjt
lnX9rCE3EtXi2uzFTgDLBIS8stJ77RXJk2WkoX37nEqdnb1rCvn+4l4uDqJh
2e/kOUP8XEeh0Ix4chiW0LzdDzk+vk6AXdCwXd1/0t7ALnto6eCuLxE3Yh1Y
ogjyiZup8loHR2est5zGavWtOKZoHQNNg/h1aRNw7q52Nv3cdzSt2WiiQUrd
VDxzaG1o85sDflLeLyBWFnd7YV19wV5uIIq1eHlhEHFADO+OgW86fwsb4kR5
kaIJmPb5KQBJW7jCe1MeYU5HxUeZRTq4UgUdXg0xOxV+1Ba9XiB8zeI7Y0J0
nyQ4Y0+y8JuOy7KZb2a7QwNaBRL33AtGy7FUxFBE+TLFx8vs4lMF8cLPugBQ
OjLtqSlIa7V58dmXKkh/7MSNh0IWp3RfIgZHK/KTqVt90b/vUhUf57Cs3bN0
igiG8TmAf1GQhn0n/kFusDn7NnuvU5ULsasv80U2YSzVlAM0fv+zEd7te6lf
Ifl1+/ebcxEH+H6eJj2gDTgAWwTp8b2FRUhMKfkOmWAoEVif56ykuWiyNZ9f
D0Vb/r6PUUayazZiDPOCUyPR3jXacXTXYy4fFw92J7YrhhIYxIAIhI8NLFBe
mJ1eKgVYihr7MdnPHBxlb/QnY7e3ABIDv4dRXbDHdodyj95IBglC1nNxp3qz
EXsCNhIjul9l73PMo3gxmJo+92S2ddD/ACXDYYfgDk4zVQsxwcUZD+Zgvsdf
qQ0IwTImhALk5nGv21vGA0aef7BlsX0FeReFex7PwbQ8m+W3Vae4LbDMxRg6
xNSdLRCIonMQdFTvjOV5nuj+0xyaUnhqRmu6ILUJNM1v1WlSKea5S0lDMkEk
kyLeVGkA1bc875ZiWFw8niNMtkVZpgXmAobC73NsNEFBsivjgJUzuw0EiLr8
GnmQeHfIsI2HbU/FFWLUc0uSDvnwuAvaawl4x6AC/Zd0N0mO3MltEUf7BDnP
AimkvrhRSFw32lcS3Sj/b5AG1DZuuZ+F0dVv0Wgipa2pcHQ33PUUJBS4z+fg
h1brvFvCC/0GWwBPHTwJNoHFAaHAfAREJEZ5NeZUBhLNqMExnAJna2dm2ALY
Nur+nXgJTmnVhVP6nrSx0hRAztLOMQWx3t0l8zyAVfZuG9eqqxOKDVKT5cAN
WoEfaPRXSVBKMiun8w+PiuD7B4SHa2dPKNcbtdXHeHwtmn36hJaVnvhza4w1
xyBQcd9veLdEtICCfZFu0GX9Jl5MZZTJENlgJVPhqGyDXCcQ/Ja/Mtz/Jkjy
avTXKw8i2TLEkJriXZZ6QogDtQ1qA4YSCTk7tV9UqSMaBIjng8F7Jl+kYBQ8
xdWmuUP5RRVvB3DsFFqG0IvbwFSKemvZYSYVG9rqZUuqn7owWz3jQDVXSJ/u
sdhC9SWLf+HryThKxKzETEfvmxIt2+ENIYn56EG8iQptZPKALZscpQiieHCp
Tw50OrVJTdgmS6/N0g73NlnKcYtiSDyw+Y5nHYhDsmS1Y9D8tM16BobvixaF
ERjOp2OXDW53DjYzOFiAFp2HWPb+ofDLgOcUp/P1msjxUUATvVDW4vIvb1em
lvwc/EMS8xUXBGIdDc083LQpj8kc99fxw24pFUmFx9apNfxHg8yVOEvjtuOW
LSwRne7k1XHFoDU0S+xSArpnVsxkV0BCDX1XNI7AoFvwWEmmhprRBB1BcrDz
0yHDSv8AYyv5KaBzE4mdc4qQSODL0Q+CtOSOR5Vx7ktGNKCK6GQCPhARkKpt
59gMrbSkUxOXl+XwaUviyCaid+4vKxTdx2B1cDMDnWCJ0VDbAEXKiymg6R/7
wZqTAMqprgKX+hYLnq+CjeKqg827MIXzZr3TtiST+30gT422iXzNjN/KPMnK
NPYFbnDYfbqQ7NmGNA58ZkVUX53BwEbT8dOjpl2XxRrprtDE78WIOMijbMxJ
hfaQwpGqUICfiTpKu95LJdcu8SyZnNf+0NFTa+cZ8h+VsGClJe1OFOwvXolz
BwUT2pWlZ4exzNc7ub3leQdPECGm/zYI3sl5hm2tLMB4C1+7pIS+j/5IYtNM
sJl8QUAwXYTl/hSqSAnSxZ4O3tm9SPIL0RHh2bd84A6TXijWmb2TX8JEBS8o
JwFAyDcAF3fosuideZyNJD8k0tuA8kPhaAVmWM/+2Ta1X7HznCeQzQL4hcJc
g6Rs6P3QsYVrK5W7Hvw3+FatED1ayosgJGRdardu42FPyJKpbiHgtRW8ECPv
4L5otM9+Y5lQrWDjd/ztq0ndPZBRefKr3/goZ5TX2PioG3SzSZkKvwDDZg21
r702iExMByFHqV7HvtAS7p/sdXf8LaptKUizYVzmELqgkvMcN0Sc0uUFAkAr
6I2zOUiKPE6+LkNGK3il+DY6MUqQjOfE4HuuuIGc4o3z78EG8OWzuLTiX/b9
bH0z+dvtZAAA/xeVYdOtn4q7bGT0E0qVuV6zGP1ZM6ruUldbH7LotHrAzPyZ
cUT4HFbwiXDvflAqI4rpLMulDEV9ut1R4Er/F8A4td8C+a0ZNrweEEAF1ZUL
8wioMehPP+2ZlGQY6TfCmMcvYpGxewWWsNuo7EjBQt0WdiAZoqBaY0LHsnDp
GoWhhPizEA8c5hn6A+EeV5Kjau1NKbhzO3PrylXaeDYz7gayid4O9wC7kAam
6svLGqSbkXPycdMoqvZlCPgNnTqY3GG9SDAU+PMYLA2YIBluMBM4uCIJS1ki
uYgBbTjoWa737jjFJRE9KR5HPuW09qEagiRZ52p20o+uoNa0W7yAYI5zmQXW
oZ7aJCsW0D7vsM2gi1VYs+T7JNBkluvfl0YPior/xZJ8Kst/tgjQXKhtB3Tl
RUmgpvCpLUs2jtGyWQSW5IB3dLxsJHqVBmO0Srfpf+pf/pNamo44Jeb2qVcP
5j7ZcH+ONw/ng7ptpF909/MvPSoMv85FFnXxbSbFuIk/3sCxWdNd2VNFQXRi
mos8ayiUs/M+bC/xCzq1EChIdYjEA9fmD879anoW2I/9fjCbZVym7AmmUiFD
g/IlREhW+wi85PRzLzN4/xvfOtWQYkn5fQMBrvOceeaysv+Vmp0E7/om5rfp
jzuYSsbJ6kbRpMHJRke+9IU7VcO2+5mQCS/vVk5bGN5dV9HIJew+qnNroxha
v8ffUTuCa3xRDspbt3o52MyOB8R65CyV253g2v62gLQaBsTv8foPzJFPeBdy
KHttErAjObCxfg0tYPL8ItIvaEZqGrtm2ezdKRQ8xn05P4X34/SpSD0nD8Gm
52WHdzGuaB1dJyBVHHUjel4z6OPmEhCadNVl5cbfuZbjKJWgEl21w4Tx3wcR
r0VUcPj4aLHoZP13MVzDbzS5TmbhARsbFaMfqldNlIZTSkoKC+JJLRX13AL8
jsRmP2h0JmhmXSYIfp4uGGIZI29/Ga4s4x7M528jsGJrUfdIRAIIluQDdkYy
uqk1HL4P/s4vDA7p8c4KBDdIDz789vronRqSBdu9xIjY5T53Uh4/v1SvIJU2
GJXUlw0fgp8Yzk4/n3ByCW0ny6yAvPn5uv1cIMuRZl2Daf8Hn0qEr+MsBXq+
ml6xvvnq+4s/+USRKCpcjVKGeyRSTTCG5iCi4gWKCr40MN8FiZBYn93ktECX
fqkRjgZbg9v6C1qzKGjOlLoyqLJGL3TyrOqwwpFwlfLX/R5lLJhvzHWbtnnZ
hW1zkpP7Pkv0D8vJq51H2SW3TcKIy6Hpi4FY2diFb76AdVH3ZvGpN0kdkGlb
LMJBy9vcJvOlzJJYuiUuJ9bM8b+72Qipdd7PV02Hr2LwlvDHqqrtHIA1ydIK
mVvxAEqYCRmwS7B/NOoJyh8JjuHujsln+7HLWNqhb44oVQ61XH0W86XSDJCc
gHvqrEYXP6diy4rHm9g8OfX3HQd9N/59Sn0y8jxIvCNdNR40TX007PcI96MJ
q/UVtMIrAS6cKsBJFcmjn3feHzzt4hbfiMCCMWNl+Z5qhehws4qBW54SkJoz
pXvOxhqR0eappWDwBaqNAGyYY433apjbrNpmLumnWv5rH2VWptfFmMKBbOB3
2r3l6rNV4+wybJtm2Iot1sAIRrz+Rqio/1JUle4hnEcpZJmMSIMK3rkyOLFC
Gyuw+qgOac9ubTYbI2XBHEUT0HJ42s0yCaYsVOjPDzMD6M1ga1jEqWz/4sEB
H2RnHXuA1avdeNp9aF1OLys5jwS0u25xRekm+rl8/kzYBmFhBmYMQoTn5cCr
z/Qz/rriXwmRveZ5UPH8UWW2z0ZaTcIlutZJ8gqtqZ7HixKGMHfA/8gZYNiP
mwWSJspuSQZXCv+Dwwol+Dd4Dh8sta8vly2W5rr1iU/DG2qjygPky7mrBZu/
RBuBvwXjNvsSnnbLpxvPJfzVBtRq2VTsnJBA25EFKGE5RtzZz4Ow/fWQ2yyP
N+P4cYELsBgvmy6Q7mi/1eFcIgjbmBjzGAKG3op0akK4y7Y5uT8CcK030i4i
hVBVGpqSXaM11lJCJzyzi/Td4dUnqTlPUIX7MncUjXwGX9J4iknUOFh5chvw
BbCGj+R+k97gCDfFNYEmYiqf2gwZTneTF2PPyBSdMqP9HWs6XA+e6P6UGjt7
CJmzKNYXpPF27kMbpI67qPUrisCxThKXjxpWeany+9PuvIqfSfCtwR9Sq9mw
WabB73NwsAIFXMBG3KqGHlpwQnzed4hGx0wBkw759BL6m7QdSi8esD8qgUgz
eLdT6VOUGFZY5LNcrqCDEL9faqvxdDb8sFxSfaPwJvQxfSTjxUHcwjjceCC0
7ephZWHubve1GyTzgvDNadfshEA5oaIVGHh9Oqw9+SlxaqidXSY1yZuzU1Js
0Ydpixd4mUSNzFDQEWSl4gNlbFfDsJ2xGF3cL0CnZeOK08rpHV04jFVO0pS+
OpOjLWtRfU/KdEfHVDfXRTvfIpAj+5vygK0Mvkirx02NLZqwAy5T71xoI+iu
nuBb6xCxIziyNstU1xlkwL1sRcfUjOHt35WN8mLxNimMqynpj67kLKG9WeGn
ztcNFd/LOxv4cyJMyx2T/6tQGd+ZCzHbMRI9n3acqZrej20mPWctHkA4NAZ9
gTDfhgAUxu6Os4MkKfEiuUb/QQW36DLMQ+gFyZakqCFaHwjKhoWTwH3DIXPT
Mrvl6DfZcj3DIeJLFHN3dx7K/2QvtWi6Sk2udBeecLMNj6rgW+zZ1sCd11Ms
SrBFrRiNnPIje6tWpCOQpdXg+BqRwDjvxLaVVE+xpUB5zBtXvg17gZCynfoA
m7TRcspnP2lWlj9o536oPxeixQbpWsxG8mvQOhheX01dvN26Ce1RZmhfGYiP
Uci41MKMXq6FcDYLXM/YkuACvKM/1Ff70Ko2eeoqkqANcbYhPXh3iVQuol4+
TudExl2iH8Rd1g049jtqb/v/MUM8YbcgK4ngC53i17RYIBSFfe694UGy6v2O
+N/Qt0lFp2vq05RL0Ze5xRtonb3JVKjbrthsmjJPi/pW+B4QL6oVmcYlFf07
5ZMPiy4BYBc1vud7c6sdHmXnCUFhnxi107hp55H7RURRlLJPCWWV4QD+4Dx7
UkkMNeuHvPtWXyMJlMvWz4mjart/tl7ZwJvMHGkTCbdpb4t3MXlwERbdfGWX
Y/lAEMHbqpr2wWP5MFut7STTnsbdIU/LKI91WnyQDhR5nxvqRNUoHtuB5Zff
hligWwM6JjTXz9XyyJjkz1koW2i8AqvcegXlf81tjAB6RjymAeYUY+lfvDdB
r8S7INsDuBnVc1jrhmaRXaNTo7tKcipl8J0W9JbtomymJ0urIz6dKnbK8t3k
74u4HYChnE9wjvVqK9/hM8moGH5MNnhU153t7e/CZVTElAq2WmiWfckorPTW
zC7kxapQc4E63ncRlv9Stt0l9Yj+AfXzIoRq55o1hgs9jSuEyMhGicevG9x5
dE9GJdY8p70Isux9sGoUDT7Vtu1yNo6+DdEHLdQkjmlr0Jec1amn+arRHKzv
myaMPlE5RZWwDOGu0u5JBaGosXaEyfB+Vw20Wjw01QifCf9ckt1xH0OcJCNN
GjB1HOxaR7vlMztX2zV64KQXT+1nN619fdDN/61AIwLExFfJvgooC5fbyer7
ql2upbwlLe2Up14ILalowHUFfVIisw30hN+UQR1hClZll1EHZQXuPIStAtIX
x2y+f3WVEIJW/HcpUlv+5z0eUsqdIUoX/HFnsxHFkvIn2VOgY9v9jN3NmmMW
KTJ4ldiJYEjrXDzAMIxHFBb0BLEq631zhDBeLwXOXPHljw+u8/Wyu+hSasRK
Y2FV/5c9GLfHp8/WkIZWM06RfQ8h6DuoHA0Hu2VxPrVNXNc5n0/cpK2zpoFy
ZPz82gEen/PiNeeYSPEcPPb6GW4bRwIRf1+xepehPXFAtYh2B1COwq2V59AS
RpS2iFH958Nl/+PcI6xVpNXTXhwlhYQeYeWjY4KB3iRXlPV2zN1zqDsAZ1zy
1MlbqterZox4A2oJA9OaWNEfqMOUjH+3z4BtCyK+coSDWOT3Mk6/bNIByGAb
zReuYEKewZUqFlTfTIND9imTwYCuXHLqRMrlNGAadtBucnDmzY84q3s5k7NC
VUMYIxihUUUw1bRFoJX+ON76FLjsEgZjswKp6ZKQRVS4mj2PvONX+hJ96jVJ
S2vOUN6fSZOhOPcg4xvI3jzLNx57VJwlGXwpA4ptcpeDrjIrqFvyO+B/ayvy
Ky7+/MpYk2MPQA6F12MsU74KYbj3V7RMYPIm0rZBRXrfGjTEapx8TjBdhb5V
7QGpQscvbr5Jx1y/P4EQAV2m2v+FY6r2o/+Lp7Y18DkmTIp7gZ3ORoiiC8Vt
PWp4GAh77szIh9kB4/SIduSt/SA+ItvCvicAt0oYSxcigj1wj4W7gaLUeXsU
rIgb/C+gwqHExCFkmtbUrj6Ivu77m7mdEZiKrjfVJWMhX+o1g7HEl0GjcPhu
EWcxSVDNF/nI0UexxDcpJdy8oS22fLYWHXOW1O5dYMhXE5M19GlBDMJ9p4Y3
PaKMyXH3tQSHYKheZaf8IfufnkcX13zYOvrqCVKgGwIkGxqI/LEmbkX07bmz
nU8bBKyefU2X6yyG6JtcocDS9A0K9yyXHYL4moCPaRSg15KBHC6dxGGVJTAv
q1e+/JOdPXcnTnhmKybTV7aE0gxD+Cub5LvYdF35kXWNfynWzZy30ldKW2NO
ewGWhAPyhpDFXcIhMI8ehO+RpbuIDwj4BlJyVOkj8RK2WEzgDIhbNWMX0Dos
VJDJ6JWvP3mmi1JG5SWvPRo2hBaV9E+sW4dk9ioOV9MvEgXvMfDeS/LU2e8Q
OVH133+6/ent0KhG4QLDkVP6poKYN2WpeMqUf0iC9B0yA5RbA3ssMk84w0Bd
/bfwdMo2bS2PN1DpgpCXV/J3S9pAaeBLK4PwaiUiByplQJvkGeJXBWmGcjoz
79t2aAD/gRtKL/gCKffyF8LHMdPxD56CjBAveVZhy3hm75VEQzSCrkVH/jwZ
cR+humriIcUhkIV0WB7n7Fd7aJ+SJU1pEf4Xkq8JSi434x6RnLUBR8BW7eej
Ei6NcvtsW65d3c/ZlodRJubEll/nfWFf9O9nCTlhTB/tOl69Ak0xNajxdSWN
9krm0bBKkydhmauchjThL0bNyJBWp+vxV195fz/3Rk8gpcpYdoQvht6Qi5YB
XJkWWeZnT3OqZ0LBRbwOyOWe/Nc1K4fpolUHzyP75BzgSO+q2mecSFjM87rD
OU8gm5IdXDFA5vRcr5Yy7ZTzGf+HQEFfUFr5FaKO4x2h8ksy7kDPXxhIP6np
KnIhnZX1Dyn97N0N/wnOVfAOsQm7ALvFXa21z41d7OneDXpVVN1TSB3HQ8Hj
rRiW9Inz5OC5LR7EigeMiNMzckhFZCmMONSoYBY4LUaH6uopwj56qDHcVnxT
mv18nsEjeo+SXaI7vXytm1lJOT1y6G0iKdn9AXGz6iEpJVVe5fbypuegrna2
DxcKwD0BleeR+uwfuXZXjwRpYSYuxUfsVQxK5ch4NOAzO0P9Juv1Gpn73D3l
U8Bvwx/i7E4V8d9F/wOxbq9gUUiOnSOXjSH35i1pusEAmPbe6taowSEOXYBT
tObS4lkkpgz5WLuhcTlLFNU/h5ODy3WGVJz/GP08EU5AFFuAhefZ20iurwSc
A4x0pjixe/X95myDoDpoBrfrhQRnurmSzC0wBEo3z+8/AmECUY4HVXPpbLBR
P9+llKC/ETWWLM1sngqbYg11gkCU/J9Fti3A/s9yphvK4UwLisjcY9RWAKjV
BqkheqxQB+MihhFbw8Oc9Y25UamB+5IGdpL1d7OVHkldUT/WmQG0kyHQPUjX
ErwmGzM7nZ4Aq2pRfBeKMpzULvTVUHZua9Smojes2c5mPWyXtfFGzl1ck4ER
OIjh1zBZWUdIPMTCg5Tpyq++ec3+Gsj9HKiiGbgmnLj8Xk9wb0yEqphUMCoj
0FGmV6d0HeF7URA7m4zgO2Xi35bGp4zeI2cIfgLOI9ZZfyprBIzTidHNXCkT
3VNVsu2aH5335PvuBJ0mN1mehwu0wnOqgLbULy12Q6LWNMIVCOBrGS7AVszF
yWp0gQ0LpcqyLU3dTOz3uvgnhintyQiD+ImE7l9wVExL1R1znRMua5uwGcFI
bAG5m0rZUSp5biCDxkbAjifAUxCM7vxoovCco4kwHBJ6HKHieeHrZiZidurG
IKmawhces/croyQ7Fx0pGZwTLpo8mjcp/JyBMAdBHFRfPT8/9BmyvcDd/YNS
/07U/LPEQKhfmn8oHGGLp72Ng62c0C/eWbU0XIA+w1C3B7CROYaXSv9vJHVr
JiuCLQMZqLuRl3feNdnOdAT41m1U2C3OQPnnXYBQ8Vk2aQ5pVrAI0zZCx0/h
rLT1rX2Z1P18dx5BqbBDB6Kh4zYcJ9cr84RiL8/MOIWT8+rj76WWKT5N7Url
tcGxWU/IwYaYRd07/nBzF/O2LQym7dPXs/WuqOuRauHE6t/M4/N2GTF7kIQT
XLyT5riKbC4aQNba8Ae8syvj7fu4RArsK50+AYpU3xU0bdMD0mC/xWsgrku3
66MeN3/93oS0wgNK3+mX0m5OQFEOHOibi+8PjHn6m8HKdP5f1BmEInCwM+n6
ahr02B2aVrucSslg8F9u0ppRniyHFOcWW81dVfaB8aTcyp88f0koyj33HQ2L
SOWgDvdly00pHX+Z+sG0GBC/ntt7h7uTqnyBbmfVqxG01Si5Zr+NtpszD7rD
+vZbprz/O87gn909JOMyiOnl8AfHn8IGgEqXFXAhv0eItBwcnC4HfgjDxZvV
2SEqr7nHNsHYh9baVJyGyDgAh0WZ2qBWRNA9qOqMZSJXmKsvn7Zh4cU8Ey4w
/mhVuulxKY9phDbPJAGkBzNgHqgDN/WCJ+386W15yzt90a/QF8Bh1lFpQxZ4
ZKT3WioJ0wpzQ7M+dNzGmhHxwo7Lb/8nURtvr5z9mdcJzDGDPk0MGnw0GOUh
SweUbGy25uP5R+19PKTnPZr9h0ulu22iIaSOSGECUpka7Yy7Xxt8t1KN4nTr
E/Ytjg/QhStOXhBWs4C/gITxyIMx1Bgsq/zeiRMN8atIPaVOzutOng2xZZhs
9RclOVvTIIdiI89avgwaKVZ2YQ8q+jfB17NPKK50I1R8lIzMumWpVW+oyNgF
sr0ElSdR+0JTNNvhfy220W6BeAdfV3Vsja680+lbBwEOJGgNJsoLoUPWEMHQ
FiwORKe+SbEOhTA9ob34UViPDWsmbCFvxYuWbvtIpTRSNVu3Ez49P3m4dR1Y
zMlhkvrWUTkStTKDSZhYLegUZ1kJAxetlXN6puSprcEweBS5wUcd2FwpNdSC
nTACq1xuUhdIORW4dsvB2zx5Bg0diBiWT74sNWL/M+b1KCL6LE0zrb3WUTGD
Yaiv/03/EqKxJ09AI3CZVCv6v15lY9yjHnYTXoZQyMYNGuOG+GrYcKqrHDny
zoygNGAsrB/ZoA0nBZVkywRJH4tAfQsHjFod6EPL/P/wo4DBkK3064MMeDrt
TjqkcG5QygOKrQCdR4cX0r4q+OFCiMe+kwFuefFARzp/ms6KjmbCq6fPTeG9
EZWTu0s9V731ZX3Qn1nLcP/sXd9UgNzaYmxA4kabP/Y91S3CN49feygKUhRB
bpRjtPw4GTecxSffJZ41o8JkojWc8MF5fstbuv6rKrFXU2OdjfRHjCBWLUW9
RC36eC0iyX5izorAmSYXvwlM86lwG3vbnefPYllR3LfkmBaYpAKokjdBvNVS
rInQSsXy2wMvIDdS7d7+vFFIVFeQqn0vnoQeCLZfYrJD+EXjbDATE8dJttZB
Q5744HZvnkCUiSyuAC85ORba8vvvoVI3ndUk5bGv8KAvMzwlmcVf02K1FSbU
rXnY+QH54ISwE4gu1AlvAILFtVEu3++/ZAbt5ZwE5EWQRQS1iTWacA6oyci8
eweSPkL8kOT6mmU0YASNP9qHKAeHfEeqOR5+ApfaTKuSaK4b1UxvjyTZI+hV
8R+bb8hS/ph/LX59WWwWHd9tHyFpVMxkvqeIofi59S3NSFeFvAnOJebP8whd
C5BccMHX1z3d7qsgeBMoSKHlJNmktV4hj1o0SU7BWpU3FTWL3HSjzXEaVHbB
Z9Qz5Kb1u1DS9ILRo3smV9GlYWMAQc4H1tHTofrFx/YdYEWSqgXrhJJZ/3SP
egnjCnMIy+5Ij/jACi5oScjA0hcKoPmHYZK0BFeE3unH6rJIBmCzboH0t2QE
3JYj1VI0JiHhyTAMaWm9I03K3E8FkNANm+XrwVnVDaZ/+ie8x/hoTeOZ4jBz
fPztFz2HSrvVBIyPbw4w5i44SPhcd9jTspw4i4wvGGGwykzEtjFn9JBkx9lI
qhQrEOsjqrps8PVmj6/g2Qb8h2JdxGLYBHC7yX3/RKZivQ6fE6rWy5XFSMuc
fRM0sgKVF2Oaqn0Mya1n0YCDJ04jm0EGbkqmSvi181v2PEMOc5iOqWxl47n3
Y4Bfwbu8V+YPxEgtww0dhCE5gKdPtjmdKRfIY2TwIMVDZhYtGHdV2HhAwDWe
jCseO/xVn9EK6lY4YY6BTgW/yQx7MLC5hs5oI1LSCcVduxxFqQguudj5AGkb
a6leo/KRBTvFxZ7rM9FsTdawdLcctjxbyQfVd2VzLkIy0LFLuKBO3AdQMhYM
C022BOgb91+PmWqyCXmwDMRanjoLBgs2AZNAecQHhLzu402fX51mldzAf383
POJxjv7HW9fcMo1mUDtHFUhExaURXnzhSRdTn6BrjViKcANTKD+wYDcf2mAC
APCwcj1ng71w+mDQ/ZBvRuvFRh4suQQW+D51SCooVg8RR6m6VeAWWKYRHUGS
Vmo8mhOz4q1wYxLzNA70zUCQgkFjaZ1yI+KMT9KcQ0/V8KhZLX49QTbZ8Cnj
zhRbqaYp7NeWfbV01vMesIXmPacf5O4jUqf2VdcB4gnAGHx+35FbJDnoZvjQ
ddDdywudzaPOXFiGR1Y28yE3Qo6VARu8PUX0bh4VfWXObmAsnE39kEGrOJp1
PLUMTBadFtsAgU1Q2VMEJmTAvqXMmEfnH7LLGezmU9jfvxNgry4UkWDw5xim
VX5RL18KBITFiO6BP/4TFTCjMPw8qReK8m6dMe7/a4g2la1+DmOgzerw+Zw2
ioxtYiNBOMUmno3LfizwnN9FQToMUS4/eZ6ElPr9YdlmPxaogHkxxdFFGyI9
V0f2UGzZT7SDEP3pNhEZ8t13vuo8Q+RsjeY5GyxkXinUmZ7kBLpcjara7wUa
F2ZVKcNbDoGodKnGdIN/SMxaPFNMHLmoJbmkAmGMhkyEEbg4b5yySvS/ZBvt
AVJS6+wD7IjetnXPZZAAa8YE4Q532Ur2y4qSa3cXZVIuK08sbE5/z/bAw/+8
TyoXILGbubmQiZwZsqEUssSzJOjmj28eho9mtjCDQMpPpNhZZ1HAEMGnZRiE
2yPXTPzhVHrobMJyDPrkh6I+HVUNvHTRt0IUl3TYJjwfkTB+8WjM5dPjI31a
IHpPOU893P9KA1Wf5XH1brpCXdpdHRdUeqTiJmQ8JExmrBnn5/Joaki8KN/s
KG3LoTqCXdgELsDOgZyeDnqh1utbByEsiYLa0J6oOEp8metRw5xFbPjNNWcM
79S8VuCUIih+6Pa0eOvn7ONxPhIv2S++Go0DNe4e1B3HjZVNYB/pWgfcSgnU
Il6ju0uPyJ9RDLidbaUnyCbwuWXceGBaoKvtFgPvn9P8Xxe+krkzwg2ozOGd
ZCWj662xdid7h2fVJ1c/zsFwACcgt57cFGly+2VP6CS7i8wtDuCm2bqD9AIw
IKSGTI5C8oJtBkyUvHD8Cog5/0Wga7jXeEv3Fo92FD5YUbcJrImXPYxOTRCs
8fIKgUe7ztRpZg8XYKGiN7lbLxcY9JrtnBMjwfwxqEpRCSg6czLQ+MrQoozB
VdJYfBG0t6NDvKSwF2EQhvTUQZx8dNLf0QzOnnNUeoRnr54vVrg3He+Ncty5
qRUeAcdpdSCsRhpICeUokI6yAE6biHCM0rkEpKZWFoP8gD4gKlMivDZGBkVt
XyfCh98P/MPfV2gU8CAGk+weDPj0x6ScN2p4Psy244Qp5a95eL3oNKf5B488
yz9MeugzrAMfg6KAr0SObStui99wHl2JiCQE+czwx7u9a45RrRdUeZG7dU6x
iQOPr9o1W2+5lJgiuTuWdQixvw8rll+y1bxnjVZewJPlkO3X0f+2MpX8FCxN
FZbNzW+/U4K4vRtcVWTYw154NS9E09tUqCNxqGb9iKMAlA9SBLSvzTYCRsZP
D50/IR1FDZEzanvx+UdbQKbxgdgHgBw/jvm5WBHRgxKooSXGcjvc40JiZmgM
iH/zmZ9YVGuT9zSctUqnZ2uftTQRXO3/IY+Gb0x0AY7m5AgDbhGxIJW3oZOB
vgbAg2MtMtUlwZsSKDvNwDo6DhUwg175uuLfARAFJ9dJlqLF16+kopxm1Qtj
sd0XKRDteb/gNxwLuVYE83en35/7R6cJP0bBg/87v9LO4IML6Ytz77jIvNFh
R1FSvi/Mn819a/DOX3LHfH3/pa2dNTpTnntmc4l3DxOp4zpfnlUr8KSeDJhG
OqAx/ursMRaOMGpTtpgizWsU96oawH8wogS4+qiy9YX7bFMOOHz7yqr2FgnW
vicsdXqEK915IxwHZdxYr7YcUkdOxwYA0zxjrmjxELVz9PcLkBeWgps3UwTD
8uyQ7HtOaq4szvTeytZii8rayqFPpIUxumN/G7YPcNiaHPMxFI8UBLy3XI2m
MZki8Yv6mDC1FnTuElHAl8CcAx7D+WONuxf1ZkPLjARdn0PzK++ZuWv+xUlX
gye4cIdLkz6IsOY7QvVLlzaTik6VbTKafvrJG/hIectwFBYB0JsXmCM+uDnf
BiovwCl6ybg1MNR7nkhD1jvpaDceN9mJh8hBJo9hS0dCNaxkI0VyuR4SmWLj
CBIvlesmbWEBmS+raoHTmvqsM8lCG4vIZGtUflrjUwxeR1uRZO1BcsUCKnvK
y5k6KPwURoalkgobuZbzgXwUpyyT97T+DRW76uMPSjYCbbDACe746djEgLRC
rJnJktjEIPRKB8JRt+ZlNJBe/bFuJH6RQ1Qh7zqQ8rtLkVl7pZzzLSJLYLaD
7Vw9OjK01FHMuG4lqbFf8w/9cXvNvEEg4sYt3UxvUfUq4g8WYYMCsYCmd8Dr
vKYTuLIwvj+7BtqncwXeZkLaXhj+jbzvg6Ij02eNMSlp4QryHpOE1ZMcGKhI
Y6BO3NCa7Ak6RguzTnFyyDnOWUDWYMvzR5E9GF1+4Llbezlbtn2CAf/9BmJq
ACNs1O/autbfK4h47g64bSaCCOZSYRgxO4NWWREmQRNzc8gbQ7VMBYHW/YQl
+wUSRK3Wv6glCC9AeuAaXRU2wl61jbd69uMs3lNZCahNA58f9MwI3x7gSpOa
lnt3DPEJeznbH9PNrgAlchACJfq8Uyo+vCNlZS0AcniA0OEmltAI56WZTfwY
VMOGjxc99Z8JfEPHb1j8zaiQRkXNj4lwAUGwhPNrcnUmlTxX1g0LkxkX/OMf
EToSuBuksSJVMLaQ/tKtH8XuErcCu8WyH/ObRwRlkfH2c8jhy30sDmMP0+3B
lCw8aivZ2JK9iULJuNt2hPp6+/SOpHbGJzs2YGxHV28sBEr9757Y3FQHmn32
Aw8SeMd3jD19JZ0ehdsRqylvCo0DGmfxaNXmsz3XVMOOACAx6X8DlpRQpc5i
bGu0dMUHXN365mw4JSn1xIRwvN13EO0wp6JuXz+qBsQYI0Usd7FWG8ZUtFoo
1LIbzC074K73WOcOn+gtw8RPAc2UQNFlVAHP+Ht8W5ggfr5bhdgZQ/nmeUAx
/K4stDl6wvPMTi/CAQrKwj2VKvGKoCs2fF/cpAo5kAYrAGfHF/nZkNgX81rJ
jtNXXqlN/5Fvxk1VasRxojgp6pdWepSmL01WN3c08zMITeMyDBTT7X426l/3
0PZJSvG3OUmoivBTaXslLdP/ElPCNdrnV3uhXuIZcPceQk8dRCodZHD2E3Ki
/e8yhER/CFXl/nv3cQ8Wp7L5ZEXPjPhhTkhDbz7QEYUGXDEtzpHNEIV2P8Bz
HEA2AD/KZiHUhaDun0uJ5UEgVp1tUtXx2UGr1a/4D4CWIj+M0u0FOw6zh53j
+vlASWlNS4e9cry72ulOJg5t6aG3rbvqr/eViP3Bi6O0B8nTiUfrNN/54WqV
y7oOXinFH2PSgslhlxSbm/ZbqO7qmTeqY6AadkYrjBVT+KfU4xJs9FdFAbH/
sg2C/apPUTgdAv4id0eSvszgwtm3hli2XLV+8iFZk6VoZpEIJU0BXHNnbO32
5ipxLGnC924tJJ3ys1o1qwuAWhHytzSA4Zb78axtNSYVVe9QUJEgd9WL1FM9
4j1RgnHtiO+PaqVm4rqCT1EAUKEuU4WVSnWyT+6582my3Zf5B+DgvQAG+Uij
X6IRZQ9MIzzHa+WEXg+Yh97BUMTVcaKV8bTVKkuuQ57h5nEx3zsGRajM22by
NHsk8X9HW0NRR+V0WPOGSbA78UPdoov5e4Aj6RmkrOnk47tk3mOrMafC/Yju
mkLJ5taCWwOey0s3n3VYZ59WdKWIWIWX+mshsRfCQSNfp2u93Dq8pAN5pJXt
Pyc9Lts+1SbEpkqrZIzb/JbI2DsHv04BfTt0tb02kAoL4r6cmYWOhiXDVwM5
ZmOsNwtQAwaa+W5q6hv3mWrBHWglZvO+TcQzIj8MURXqPIe/0XHo3w1u9D9e
tBVBegy63XjVtcDt7I7oLSnCxG+Su+9FmGStBuyWdSZsz5h8ZgmTj8y133Hm
9tdIiTvq9j50ED60Tbimk6yQDUIiPQ90LYNemqVUupLnO4J+KuIxxWTE2Sew
bT2TLWUhnWf2P81EW9ZdfDc69adkg0yVTfcbHv2VqrDHvwnc7fds1hOvQgrV
o1lvd/NVhDNLJbvKGUflaoE+UnZ0gb2Ykc1ofUoDKrSiQFRBqaGwWcD6TvkQ
ag65ZX/iZ04eC4TfHtKWKnrMfrKp7J6SZLFrjL/eqE58ydIDMCtn0EKwyR+G
q0lnsF/rWZP0encptnERmJh6B3TmsmOAucawGSMpZNqPBlM3lNZ8HnuJNcQE
5MlJ5amflLw21WQlRDMwHcJNaJjpUuSKLiGj21voDzhb6POiPeAmhnfLrIbX
2Z3yKEkMZ9ItFLK2OGYeYfbR9IuC4N5BgG3fFAdYgZ+OQIvZxSibk5u50lXw
y/VKvATjpQuPXJhagB7uJFfzTUASLwS4AlpNyqCWxTQkE/HJYc10zWSE+IPS
5IXRB3/Fc9IQQPVhT4WAwvb2SkNGzRKTBSRoIBmqkwBTe87UB8G4j3LEvVeY
ECu8BKmNkNsof7na2niVgI/O1WNzZrxD4nnrYYcq+BqRVuQkewPgSLM7usrD
6c/TPJQgfnipJGC2cJd+tcKeAn5b1rx5vK1jY9VMSM7iO/NCxVtHZ8QncE7x
/PwU9GYKAggnHCYqjJka7MmeGPxoTbjDCpwYqPRaH6zGhoZn6ih/xxni4CN4
qfD1Ya8YikR06PVBkbRm5eDO9OKdcmApLj9P9XDyxQNak/qqW+FbO2fawNr8
gQ6/j+ECvjqjYh87MQfinaP8FNM7Dw/OwQvMLMrz4hCEFGj+rYYkY7iiA8tL
j3UV+f97wDIpKGO03PYnpOerUHfWEhcH12aRhDST239FKiVLa7kKDWszsFha
yhLSYzc6oL11EpkYoPnG3lQhXw3oaLGtXQ0QjiiMNrpJ/QRvztTInYCa1PQv
sjSNg8rk5Aah70okX/VWF8UR0NLxBr8AXzojs6stY5pi5llE3mnkU6us5fkn
QiVEuvm9q08RhS4o5wEODhidJHNDvQjPMDQBy5862sKt0j73SlkvigUN+C4c
fELH+so2Rq+hZxx27BEBagftsrJsLUZS++S4mlR3xh6H6La4Whg03dfQUwc4
5A6F1fd2J/SBYnGVaE0mZzIqhrC4RuA5M8Y+UbIMIK1uIwsYvRh3lmOqZDy4
ACGSnGVAN+rt/ia/z5yT2fioeUAncK7BvuIXc6Cjz3YiQFYhu4/qHgmE04+/
YvKGAkFfA6ci67pkN0PnBYDYiKrsgO8QjBN1KuKfwJAUYWBWjQ8Ubl1c2KQ6
9CEYD7Q5BtDnnfWoH+72jK5IzRUDzu4sl+DTrz+9zt3lAbZo+VnHUWa2rMJL
C5y/CHcNT/Iq8R0l2z4m+RvlagCuOW9o0UPSSi8BAZ8y/b/8Rs4X3lTFmOFE
Fw6hh6KgmVgNwaV3nywYX79AsE/NpgG09N5DEGsoFA0GTTtMu653KC3T5rsN
KIAfiJqx4M4eujSr8vSGponpigs9DmREYoJ/pwMCwIMIRSVINrLZSVdzvV8m
PSjCFRgn9sOiCQb3tNC3cnTyQIPJp7IZlCmkHAZtBH1qhEAc8myx1bU9EdH5
1dXty0J18tA9wQUTBbFmk20X5VRlWqeBqbx7O7uU8VyZqtiuKiS2q4uoa8Vp
eBmtURE/EAU4ZZL8v+uOBaKV+qOi0hroJ6H4a4asL07h6KZamkRV3SbTbV/B
bPsUSd5Ro7ziI6mqGv3HqtQiAJzOXblFnRYY9YEgyTM5UmqOxXVMiwrphxJ/
onmud+1gfQzHUxmCODXX7uwBcScq9J18CcFNNpsHoka3fwMWjIstmCYlMP/1
+auJL/qHMgAFcJxdi2TXI2AbFPMcyMXZ7SrSPloViiDeU2k+B27/tJCx5l99
CbzOfw2LdNTp2mgjNmM0mjXvg9NqzZagxHCNj6F2jvc9nxWGSC4jzWKEDYYZ
5YlMhswFgq9pRXW6N2UC4g2ZkSso1b3lmUeMRB954tzwjvfwfWWSqhitP9pY
/6/v8EZTEDqNf99fV4ARAT7ss1euOnnGSa73mCVg7cF59Q4uI75cLYbHD/Ue
TCxOgCgHNBDqcAdkkCAo/q2CwPnzEFIq60QNXMTiNBZvY0Pw5K6YGIOt7V14
EvemfUW9agfwpM3KPMW/oPd4oCJVt/jsYM+aNQWxvVsISiMLA5WsXXzlrBmo
GtQHGu/4Cfx0szmbMaSMi0wHKU2ba1BCIiU2dSUhbAi1yNqYfzaH5dSiw2VV
GV7QVFTa0N+CNQVdlDwADN7pSSHIhGAdULAMZ0+fXBhJb6/sXpslE/xshrVs
bHNUZjTb0jWf6aRjWoVHxAJQwqhB+JXQPSnn0lp0eUGfaBJz4aJV/pG7uUI9
MOEx2X1VC7DrykCdmUkGzMwSapO6Xsq96f2/SNk08oPSv6vK2DfJKfS3xCnd
4fb3s1om2nP/kJjwR1l9A6x0m+8qEitHdluKq1uPSlVemAVbOEyIjzax87Tx
p1TTHji9w1Mo0qOp6eoswr9pbZASIejvZpcE/vzDuKhlRE3GzNMlGFJgiXsD
KUZVGuOAhWCSoR5So5hPEGSsE1QJsoUsxCPzeka3Zln0sRcLC+hrsyghjEA/
aqQpb+LMa6729TPd9BHcvK9VaO/OUcPa9sU2YbyUCdgf4tZSIMHh0K98tdvp
YRTVEpl+RrtvdOJONRoc09Rs+W+DO45hzTZnxlgQcCKy/DovC+agX3T4lkLR
O3lInZRNUgXKkBnehfqn24CPUiBkRRU8rOntuXD9ylyMVCRXI4PJF1c+d5td
G1WZkyLQaZKMEiTcWwSqGSFmI5TtEeDu1KHUN7vJgxxbhxTau3n46qndKR0D
iX2IY/PrNCNBzaYKYcRe7vHmCVYoKICfwdNm+oSMvkTW4tb3b7vuf+z4hOg5
VnO3VEyabCJku19AT0fHArQS4m7asxMPlYuqsKReLKOMrlghL3e1C/Vm7v37
52g8B6qC+x8QR9xTA3RV1K4vQnTySlTLZc+yeQl5TpL8IEaTC66BY3/97jEo
D3emKQxIaoPGg7Jku0aLGIeZPGD+qzPduotiy0CKu4Zts6kCvK5LtTWJZ3WC
OjSZghj2GnPO42O6YYWz5Vuwjr6amlhtZEEtERiFzUJp5Rqo27UtsQyxs9Rf
fdx9KpvISgts4uVa28vr6WfaiGNATka4J4KBv8S5YSeKWCI97No8W9B94Re3
x5sHqvOzExMcagBJR5YVQqGlBYAjTVt4aE9+DI16+9d90jR8w6LklPLhOS0d
73Wb/xkMqI/fwK4lFZPXvtb0755tVNQJTLgIFBtOp1uBiv2v4TmbwYMdBvnk
JSElob46vBqLgraANbN5gwKZE0LBUQIPWD4+uP0pDAEjLlDJwLzCUGOKt68W
MHGbDf0JbH6b1/5X8g+kYejpO87TJX52woMguhjpBszJ5ettmHKRumAnUy5T
Ms9Phq08tWpkDUcXS9Hc/d6UPVUXVFdSkugx8n9bL9UhZkCuxFT/Orr21a/7
1CgV3HaNGf8QBveD/LzCUNgjk1vNu2DyIZ05C9d7RNnOuXfoKJwArZnJ4S3y
F48e9hSia7N0L4PhK4ffWj3R7Ra5RTkBB3ZP2wYXdzN5ueqHW51ll/XwTm1k
jmupk0NXbg/YZNQIgctm2ohy1aTGpGhK6cWfUgvIQrZ4/tb1JbhkyrqbDiTz
VoEakENxBZ155G3Jc5+DgDSSoFMva3GVGd4a2V+2HlqqtG8k7VDCX2Jsz28o
cHu3IDeZaxrg6c8x+PJXFw4vuKRXh2kWnR5COmip4CJ5Nuwdf/0T1rGgtvz8
mscN7qvFHVr4AOzAxu1eH+gLFf15vLSccS0Mrtoeg2jl4upFJNgYj5xqMjVV
icbQHQtNCJAv1gAXaJca1MhqX2m7yYj1z/XdCbsHw/CGaX9gPjxsR+9MYow5
cdBf4n2mzBkpjDcKDqdFCvQ8d5bL/awDhvhRBS33BTEegy5BGWno+Im6O3Lo
NCLBLt5o5y3tk6e/RkRYux2iwCpb6hXPB1kcfu/nJBG0hjbG5XnNFCct0WgQ
++LNCL/G6Bpx8or/QiyK3kqiXGhWMEr5XxbdngS+KA5qdsOOHNHzm9ig2rZp
X1qlmj69wonY171gWw3vzgJEv7SmMFXsB2jc1um9t0gmkHAx6gK6dOPamyTZ
4LHgszlOqSs5tcahwHCC0Plt2nWdJBHjwSXwAe/ceiXxcFX7zDFlMZxAwuGM
0SUBEbSmfF/4AUIh0JIx2RFyPZQ1qRwpXA9+Q8A/f/JOTE+bgj/bGUBdvoY4
fW/II68xckAXkZY6mXoNjdIQh2fdj/eNHkBesdz+Sv2KoX+opcVOqTo9D60A
kESIgIo3yU1XacuVbhGRO7dTEpw2q49DTLDT1g8CZX3gvQWIpGjjB7tPxhfR
KfYsrgZkCa+ToM6O+B4suvKg6xz4aI+KnYRXsH6m4iEeIp9V1sl2ZxitNW9U
2brT3F/EkWYqLp62uX3VFoeEoF2KIYQYRL2MpoD/pY2u3aE0GSDcuPPUXxXO
TKkuDveBtVMyQ+gIQz9/dLkAWU4Ba298G6YSyRdI5Hi4VqmlHgQFnH1TNjWB
CtyUBK4mJsTWneeqiGGnA/0EQFRWeAMo9MrGE4dkuK+MQOluOcXiQ4A5WZHK
BiQaKZIC+NB439qyWON1f65mwp8rQibcSinMK4YoHTc4sV0YM2WgiMU+y/S0
HQ3X2eOAzLVM1ko2aAAVRzpSMTCtCxSibAAxUhL03q6eZzrj0YMSu/CkkUwD
4qZiC5FmZCU8ZZRKtM7kPhUSEaeHwPovhSe2itq5VoHKTYNxLzq2n/7keOpN
QlEqNSoK63WUGgc4Lkto72JY6gukFh5ic0fm7azIU+fcjFwWNfwLgX1kNKrS
iFYsmVOkbBx1S48aMMzZcrEjg6k5oz0UFQ3l5QGeNprzWYVE6geFp2VmbdGu
jGlQB5e5cxMvzDAf6QGNMNzJuWFvXrVEXxFXesBg3svLw1d6mgwkoCuOMi95
NBTrHG3UJ6PjrIKr2eHySlQWKmLY3eAxQY96zLtWpu3UqCiYFKPXvI50Tnxw
fb7j4WiwsEs/aM+T3pHUat17Xa0+hWXFAYiE/UT4QgI2KY0wHekmjK9Hy+s/
5P3YzJm0JG0BR2E1aHdFqSgEeJ89rE90PaX4LiX8galVAiKwU18O+kTqKwzv
yG3tfClNdbv4vki1a1XHJQT/vuMOT8mu6UjrrT97QkdAB3R4Les37UJdAC5q
DrPBMDuRqrOykG168PoRMkj22JkZ7QpRaKy8mVMP1eUWIgjmRFQq8/E3r2iz
OO6LmZQX4snQ0XxqQ7BwvOgP+KbdEY8KcJmmpBVI8JDac69joOKkT31VGFNk
fZ7CPYkb154zJ3/7vstr14QCmVEwChD6aNIrFr+d86NCHMkHSGWsA1ogTCTT
4ARBTJBc/z5NxgzhytYFY/FuEmBZTIVK7TOx43zhC6s1THPQphPhx/r9ngNV
O5ihzRrNPFjlPoy/iU4btNnuo7E5GPrUVXJlom+Ctg784+IEfT5bDqFbZn8P
pWNq1ePYvIqWnnQ1CcgoRq2OgGGnyDLaUg7DqLjEUmUixEnAYJo3M0KHgYu/
JMKSrMU1TBKlQrE/Hmvxyg0VYUsit0ZvHivAiDjqBHZ1Iu5AVcLZbR8+9EIn
cFv3FKVmiTyyS3x0+3r2HZkN+fPKflMP7j0wF2fivNNSAv6pNbSToIatXem9
uEzsgN0Vxqu5k2uokb3Hymao7sUXqQz+etIx9dbnsR/KAaFrZw6ExXnKEFFu
dxD9b99DsRkHqlPXjVqrMGk4UnCdwGOKieuSd3VckI0XlxbzgE0wNZwcJSQ6
BHEUFkiNtb4pEvs3uKJooUA6vKnn1cASnfe309VvnPtzUAhZi2KQoYK5OLzn
dk/ZyzYzl1WxNTtqJrJykkd6e0qTLctAv0SQyG1LqajrEVEmCPk+pDFwGKE4
cJfstyN9YjsJiyN+FcAMJOqN3MOSH8oy33o+4Wlau6EmGo+c44EHAE3yCi92
vLsPO+GEOWt+nqg9zPqcokbF2AR6JrsBSGt9sOX8W2J3fuCCtf+NiGo/FPCO
DFkXD6qnlZ39H6sK5PV7avha4xdoLb8KfmEhKoLgRb0guWdsXDm7+YT7uYvJ
AIWVlrh51cGEoh3Yn0WmtAAB8kAAHIJ1xzLuauls1BQGnFm2MXk8t9GzMa5d
V773WWVYpGoOJpFw8V+tgbwjP8iL/x/5x3XP1X0DVdbgWGFM20bdUPbyCZKQ
3GdefVBAHe29vvWrKPDRtDdac1vMMf2GNBtVi42PYjwC9QtyC3pYb4/7dLlu
Ajw9aNWyQXHcejQZ2WbziBb1YWgugw08BiFzWeRQYdzgre9meEaC941YhTR2
xbgn939IXdnA3Ucm5id5/ZEPrbWwC6doHXZOMNEfRzDYlZW+HRT+FHSwv97U
3Z51iHNTeSJbsmhnR5nR4N8NPfrSfIRwsoS3mWKl7ey2nyh60jwJl8YRg6UW
DtxUgFekZRB+VyJR6oF/Kextiailm5FQzoqw9u6YdGsHU9BMOT0Bb7RbztIF
cwU+sEEwzijdkZF4+T0A+flYXDbvsEApiIR8EIgO2AbNUAVP3BlHg0tZpsV/
3iU4dbkazBPLJGhyHdEBEHPBVmkQtZdNS4Q+9fh1P3cxq6afFxUIqat52luC
c7UBEFwM/DewDf90qKcVwhFpGErbMp0GeIPaWuAuB3XS2Ef+hOvFBc8o4byl
4aikJBz3RI81hSBEDxOgm9eWO7XGJ7z8iuu9N1kzSxcMCkO8GaTKyn/UsygI
mpVdpgg4dsv9cWRZsQL6i6WAebokNjE4P8Td6PMSFB1AaN4llFttEIkmntJ3
FaSiWa5f8PjP4Wf7gZcDB9E1gjVvSY9nXN++uTVryuLzhxVuUG0PtX2tyYbB
dOmXVJ/W3gsWIVmBQ/HDSr5GkkVaXJwg2qEmB63MlRnZTqtguoPgJUCiS101
nh0Z52pcyS77LwMMkZxYyxrXv9oXIqWa3bvzAH6Drdd6SRZKlkHcdSk7nDz5
M2TWEuREk0ThWchy5DZe2KMwyFSmjN1YrT9lvwWdhNwkewNeTuUXia3su2Lv
DWUU0zRgwusWdIQfS8NSEmNoPVI0rH//Zla4d4wN/ZHfl2EinJrFNK9MfdKG
MgH8ZPTeG3HWtYOheG0N0ozrCs+MGSDZ9K087JpQKv2+p9rZ4Qspk32qZVrT
eGpffzrw2H3HA8+JxuSQUuuXU/vnkeapxPA+hN7gcTPWREKBpiOLCU/DGRpE
jwE/FgWeUsSnW9lwWgcPWsenfToR3ntngQx5EryO0v4NVxCssYVAld5QfWdG
loj2hHeKslVdq38Dhd/4juhJEEKMVhi6HzPN0QQ842Zba6sXU/ui/maQbjYA
fbpOgZRI+i87GXSBV0k6ysaqzulgwL3SMvKy4kER9FqwXbUaS9XlrqxLGyYx
qt7/093ptKApLjFQmn+o7B8eNmeRlPDLIXIVfcyXd04sUnps12olmTWjAafK
LN1O8Nj7bB9VGbVHKRT0pom5tDctjG+m8+yOsW2hODjaIaeHfxub1RxeoZ/u
wqKna9+8SM5Y4qBDXa4OFhlgmHzIDevyZQvrwr2+L4PF2OTkFVcXDmKkNdnK
9p6BNzQ4sPj7lI9OBG06fc2BQJdwI6j41AH92UNCLgNEaspgYRgFR6aBo0Dv
h5eDCn0NAtKzbS6cebCJ055MLwFpCk13x80hQWUG5nrMhRv8sde3Qq+3ElVV
Ftm4XJV2qtQuRW2lnKwXjqlJa0Q5mmnmYjLiVcjt88FqfH9Rk4Fcro1H3BfM
XGeolc5cIi89mVZdE+gVIQlx3AT8MuXjJ9UMdbt9NxeCdsMGllpp0KA+Nu5N
FaZYKqWzjsmoNIR4Jp25FF2XRrJZBuJfKeOuqG0GpAL051Xs7ymnwExbP8zO
mXiqOu69GeEAsNQAgTZXj9Baiw3Rdyv4V2ti5VD1nXPEt6KWn7j3Itq87rKB
0Of9dfd7bydqjINkOw77DM6R2D6ONxdSpGQlnJZI6Un8jt0yba5E8RV6Rde2
i9kyBkA8XRuIM2YVg1be1vt6dMF6ZbvHnHW8j8aiSmGq3r64YXLH2HPTZbT6
mk7SRU3pAO//KngjrpOoTuRvt9jwoBTnrPLO4NuMRUU/FNHGM7SnQU3MBarn
Iacpzg0Hr3cfrP+gQHucUnOT5BskYTAIQVp537rTMDgnjOIa7g9dR5KssAQH
4zta0BYO39uAfZJhzjGVgBnsfulgubvSHnWWzyZDTRjHjjAB6nkJJM3sT87k
di1Xdekhz4avxSV7MiU1VqFPKTbBv33FpGV1l5vbgIVQc4WkqRYi5QZ2mlBJ
A/2KYrt6/TV1S3nPu5irfvWK9ILAl6GRqwM+RDV5ISqzLv2LSNMAwyDoAJ6M
Iv/QB4ZYQBJdeTC13LaW4O2FdMeUhk+me5fyy229BSHg1CbhA6DKgJVItQR0
I/fXZdX6W04eusokNWG9gKZAFTmWwTwp4YyXkBJCrKShMurSR78HH0XlZk6Q
rRoOijYp2ERfyQugGBcL1j3MDn/gw6zt31eVEtEAqoyV6n8bh61pbuNpzFKA
6w36RFCPgohYZNuPXjsS0OTJfVjzaFM/5slnaDb4GWCQfjIdl71mvqW5p3oQ
jUdMBvZpscYVqOQdMJKwznxshs6MfpltDtCClbTNJNajmlfp+4q9JBpzM4q7
jSaK4e9X/+rWpvZVp90Uym2/bcOwyK3OW7sI/zMD2t1elZ+dhIqN2rz7zy+T
UyELeC78wMrOf9NUMwmDCTf3J2yf/grpSyZysXxo8ixX4Q1X57PQsXcj62xM
LVImoP8O93sRQM8XwDC+hf/E0wYqQH4hWBLww7jCNlSMO9kqeKnBK80kkLBj
mTII/5qVIqOiACZjiydcqek5xU2y925NRLLUaMclp3tf/3YAyD5e+EycxInA
C9hHWRMxGUf8r4ilHqowATYlyS6feZFe/QYAfcKXY2vr0597mfrnq05iDuZv
XqVwmbwNVdeb4xEII7gmmlzHaHx2qkOHPpyYfM3E3ILUSDHuGlegR/NQdgDb
DiEQv3MyMVATz/kcYSuazTv2H1D0JoUNDAWYBJsQZm/2Y6bO+7LjGGRWWJm8
EB45umI5oiEOV94sx3biKhuCyRHqVE9WzrnnL2/+9FxSC/FU5tqmw8ovT6qs
HhvO3fML7f8mqKXEN4oawJ2xrapIGRz+Tg5mlZ/vBOw+YTZE653DBrkCx1LW
6JCYOxz6qd/kiBcDyJGqHzGKBhkVKLCH7IarS2PY0Iq0PisOxbhV+fCPkrjm
32y31/14hbEZs41HNQKvxm8of2+HrJWtWbdvm/3UPLLEvkCZX+0+o3YbamXE
EbMyJN8tYhjIeXX5jfY3nwSYYOsnjX45zFfFAeoI0T3zAtoCFqw9UMw4NPho
uDgieTbCWmDOr9d/11vMssZVXDgJee6ltFzfRxHvtMUjVv1sht+jw8ceBSBs
X6+a/x5a5ERRxGEOBxGPEz93QISnZdPKt96b9Wg+7ThKRkO3eDqKTitVk/qP
38SBtrxc9buVGVvEoNLHOCw7bC8QnBvpOJYWPK/9IkDZ+4zlSv1BV9zy7bfk
UbmmhZKEj6mG4uOfn8EiLT6jrgGcsQdXCDfrwEBJR7c1FhetQxIv7MZHxaqH
Oei3ssTsykcnZBblZjgn9WyCWTPYv522JHBe/ammoE0Ys0q2COye+/ikB+Gm
U0/fUUq3DjcTrU1mfZrZreWO1gGfn+f5gpVgw4I6DQEHSiFlOiPQf1UV8OwE
a+p31Fp8Gu0Bl6gMMTXpu1ZQWGQae1ZCA7ro+5GKmNLmtTPad7P3x32QIc9r
nCSVJ1Bhen7RWgTxESLvpxmq0PaPlVDSX2KeLC6f7zGo5LeO1SWrzg6RW7rl
D8uRAVFfmcGWYW+/fNO+Fk0hxpiMpeyvU2/KhCkp+3+iKMgs/HpSEdFAfxUF
LbBtGlhkFrkrICjAxeS5K54bZo4FkLu7aGELMfGv+J9nMvsibZyF6bFC+Wwy
HnSXNCvHdhbRlVwDTAEzSWTbyBkHQ1O+RqH1nUEt1PnsPLUdnVsDJpBc7sxJ
Ziwf+cN5FOlk8l0eedVCvpj+iVtkDS/9JSUpmty9lJBMfTeotc+/jEUzMQ1H
pfSAB7u8se2lTo8fD+vzNeB2r7xocA3TeXUeWbC102MM27z8bZdrtIRkB5IF
tcpubtBBYMpwaq7StVB6BspXgC1W8P0rSFxl9Tqu0oq/EjlqtSn1TsjTIwiH
XPXqqn8VeBFYDurf9UCoudw7ff9Unr48CPHLQ+38U1lZIkLT8DFPYUYTjfeS
ZLcPlZZe/g7ucPbU8E2IV7+K/WsrXVVZC58hm0kvdx3IgzRx8bzYkVBMc3ly
c/SuAAYkfKWTQ+1ZiZblJuabE1OC9412uqs3hnQae8s850NTxzZ5puFxJsVm
xgTnrJaKRhHFN+xHV0sjwS6GmyU9dxeyXXx2MNtW31MrDnUeABkUIlwMUfK1
a+Sy+jOw69K+ROTvVcEwbRXVLpTYR7AudDcBhRxdsoFstresvVAmkHElhlXr
nRedp5KwmER9eWAdglhMILil1rJW+PJwivEqPYave25z3TyohdndnKrhraTI
+YhBaQydHWLYDt2nJKIefv7KvdEC/Oy6O0JDoHbuhZmL138dXBmdPlooTMwt
OkQfM920ycanhGgsRbfR+QeFcGwRvcTwa5Yg7JW2QAaoQuO4nfpblFb68p6A
3nzAxk7jXXdTT88Yjrfg8bRXHEqb8oWUyPK0igHE3LGA2WG6KkjbtpWpUJA2
0c13Y0VrRokuptEpQdUE41zsnrvdLZusKifN0CdHIonWteOKu4Ly6liCDO31
sMjDg4ObXrEbV9vLO7PEv2e9G5IEjBPYJSd1hOcQlPCp71kVYmplL/u3DCcN
fKlNZYuWExyJNbHb1bsSy/5FywE28hWHz/9xXkgkW1A/WSjEZiXz1fTLKcT5
T/e39upQipgg5n4zuzyqNS4ZZkiOT3b/G1rDlcK2SgWKF5pPX6ozxyf6Q0Le
RmHJgDrU0ca0RvBlTBRQjUGj0WlKXquEf8SsIqpkhA4y2HSrRwPRy0nvslO5
Czbe2DA2i8kewTho5uflIf0f95RYgyTtVkJ9zIU3ZJO/G8veO/OvRbps1ENR
n/EiDQtuSQhNegK/XoWIXdXvu4TtUBxOhsM3gPg8x61LnQVzl1cZNuPrXtjj
uyk5kva2odhVT4oZphfgi34rTHrqxv2Y6x2Pc4Jc5Um7PlqVHu7Jntlaiijo
CuM3AkRsP/ShmCL2f1jj0peBnfMRL2K4wV2AofhbVZZT9xeaE90D/1PXLX4R
U/XDUnn1ds109a8940i57nDLJ4xcUhZFi1DImTPrZ3TOlK0/OgjZqST2Bh1h
zPI1B1x7sqBm9iIPwR7/oJc+w/Y1VKVyDlTf0+2hIv38rT/d29jvHp3hZtKi
8jKPKoXy2APG1FP3w9vSiJG+tG7PryQEyQpc5NFXFfg+JUNN8yJbnMJNGyRR
t8x1Kd4X/FLOdrJEgr34hRVsZIHB2o+6cswt0x7s912q702zmUDqI0aGZGxg
ntfC06xhxJ+M06O+RJFzk6Tzf5eJLQVUrgFUk9Ewg8ZLP13eNScsGjhg/RpX
EwwFwNAs7YRXqlUw3TfNk/vJRz1mtvE27y6xqLliYHy2Y5tBlXLhjjqL/cvS
WCevkCQb0oXo3cOLMNfl6fQHzDWSIY3jVUUcM8FuCfoxJT8fHCHxMhNBfJff
05u8bqmFiL9zyChyT6DgppfNt3dhSnLzwoLHQKtUFG2hYDnixO73nOyepo9z
VynIBGUBbDIP/PYwKhCRGyjaHhdkCp2Yt0b/W1NIZqvCSvYHVZ33z7PelK3E
fzegX+9WFEnJdd4iMxBs/YAAc3VXmrRWtC0UhCBwnM3InxpaFS5jN9AQh71N
WKdtqt29t2fpZ7MpBZIQfG/KSOKWNtMAiEiT9H6d4i3LS1Xhlw2tsGKnwI56
EQ4h2XVYXcpC0Fxy2HJAdRmWZyIHpi9p6eZwf3gmEHQTsHXJqaUeakGT6+Bc
nGrd25h6y2Ql3yQcYPKgqd4Xo2yadF0DX4dwcSxEwOXjCiGHqhGPCCKtfaCw
Rkl1UzHZPirIs4Qrssswg/mUixkWjTYcGjC6nBBg8dIpd4fQoRcd1R1D6rOp
htEtLQlnF0mMgbr6y/Ep6hmaO3gYVKWzSWyEskRwGznsFYkVSbxGg1kBlWcJ
IonrtHzZVisbJhMFQzhwQ4hvWhItQSAOP3gpzMZ5PfGqxFYxTvizZ3K+BASK
yLC0FeCi25xT+uvrNErYgIFx+5Rfp9oYnY9XIQEPlYA2+OcKbhetl9RbkxN7
FOm/w5A2KfvzKM03BQWvdwrMeeWl3AyuWIxj1T/FCb0DlXWxmk0uLBFptswy
pW1WTlQCky8WT9/rSGN2Ri9mvjnxoNVa3IG7tcjqasgGbFf+Z2VhO4qZARPT
p8/0nsUtlz4k5ud0sgqEJEi8aZ/G0qSMgBzew2qHoTbQqDNvvGEZq1kRPLvs
aoWCRkSuwYJUc5+upCLn18XnIgHQ1YpUxrKSryUVXccPRusBqRlEThl3nOJx
41RJFJmB5UsYuFtt6BNQusr/9cQW9SpVxlSKGQLL1WcQz66M6s1cUHJSxPB+
l1GLPeBGR+FGh7fXsk9Y0h7Qnb9ub1sAMUU1ZyfGQIi0dLkNabqnHmBj9awO
H/skZ8NwKuDrATW3KUnLdHKKfr0h3+Iukl7ETmvSP1P+iVL6R4LzJCaJJp4/
jcLnSww9Nc1+LVLUra3Eeq+n9++4/4rLaXmzlMu+LxX5t2ywVIRq/6JDVpqw
vsgPW6c6bdJxbukL0Dg2XA02/7mqMbCSn901INU5tTgk9hyb7MRzRsHdn6f9
+Il6XcinyFTfTeCXQTx2tDP4rVH+qA2K3oES4Sz7g/jd88jtcB5F1zIZ9o2g
QZegCDemtZ4I2YGItFyUcXSzd+597c3vr/rYyUSXABYAzW7/kzgqBw1GStMc
zhPxNkqxEW/bc95dSGjrHiWjYvtEUSNJhZpJ+UI35Uy+7+4xCeH90HmNJw6M
2fBTXYy8naZV7Rr/9OyDRtNjdCe1exTNKyXfdDtTK9tnY5Pa+SuN/wHoXAtx
kk6Iv01SKATf6w74G6/nh5/vWxkgfAUW/20M9LTV3SpxP3ffhrygSty/MhRG
f/cStXlNZdzJrofq8cnD3C3Wwd8yNdY8OLykATS1K0+89IqJ+SvtDp/9NcQg
zKYlI3nHo66THAfzRHudJc+et7HZTL7NZreSp94N/Me7I3AUMk71lKo9H7S1
XkNfECWG1zuxkZo1gd3OGAcmJPkr9lNKpYV5nqbHF6386OhYbq2OLubL/Xed
noYf2S+fjDQQRqRyX2qKUk8WP6FWCYdPAxrOBnoUMPRtgMK3yOnpqS3dOJnQ
gnn9E+yJy0m8wXWafjOcM9KIUeuTAyS0PhNuvV+2ixJPUi412Vjzlqvf01WL
n/LQkgNJioEngQeBC/nf4fEUGvAHrT5XNCvZgaovSbFIrLCmQzyqk0lCDUdF
ATQsydjrvrrzw6CwvUaNFapAdzvQvKMUPJ+vtr5sInGbNY49EvflGlI6l0B9
kdgZIERcmnc3AqY5AyjqTGebCuMzLl0Rz1a5ycDUCmsjuf/+AgnFF4tE2J7p
3JiK5r4ze2byw31o4U3Fk7il9gA3eCoQuGjx1ApOymx9QS0yEJhdHT3eUMNB
MpSZ4g0ch4q+HeCDTNwJloL04PX2+JgnUgjnt42ubsCyKGChgYG8tk0vQI52
ZwzI8iiBXVSY9kfmARfGenncp7nseTnFfjUSa04rmmW46ah3k4W4l+KRWMAN
dfz3GiPcr0TW00Sof07koS+wVP+HanQUUWkTG0yZ0fpug5b/wTEwX8jg0BhG
/fDUPd60BmWMKG4AtjY4++pRg3715gWB/G1tWOfmtWjHjOvbmJwSaRenVhUY
oGhvZqphYE1xlL1Pe6KmBdIajFJ6P9b5IYZrb4/4Pxf/P+H74lSma68OKvg6
8jLnU7b+AEQrA0q66eocRfFwivNKL8XTsoeyr1kT3dv/10SxxZQzxAvLrk6w
YN5Rf+8eDWfADm2cVbhRxFRVoxeUooEP2tnd5YNBV8KkabPuLMcZHgaivpn4
R3SYeGZ4hiMCUG53HqSBSLcs8e7oKEGmdSG0Jq1R/VG7r9NRZpWf5FwuMblP
eieAa5E10jnglIFHchPPJol4aiKjv9LNjfCOr4YdxhJVxS+eMY64oQjEgvBg
KAZU7bEkXcL5dVhkRT8mK18zUaPtAVececlgZCmInZcewAMqMZqKjfPNgBHy
IdTp+/ynwGXXpd9ScQgfr7RsQGwEZnj3bVyscZSfZhRmOJ+eNPQEXEhAZu7W
yWnp0MRObrcX6GPSQzhe63sdg0jcZ6AAcXz47N/slFsDBIehroMBehs0A2iI
uJsHNXVem1DPofQxUkIdSvlR7myPZqWu1Bxx3iL/M/AQVVZdrUPIUxwg+rhV
65vcZDHqV9UyrP27TM7JUvkkOAVsKdP7FKT4wsTPkZ++3lBa1Tp9pGNWJNCI
HGesYvGywFl1btdk8R9UMaPTOoh5XaDQUmoaH2YYDbX6oCskrc/MOBeETnCd
r7x3WqS6Oix03MdXuzXZoR3ZGsKzU6F110zBZhxo1uCfuzs0YDAhVuQPWjq4
CxTCeJoeruBBBgp3+UNJL9RUgemT50DGxkcgk6gqehbHpO9R1rnCDK/RwVW/
oNJX1b3m8LoVqWxLTPqSNqzj4owEo8BrDvbKi2rsIaTWA3M2fzh4Z53jGkGO
jhu/hGG80u2SodfLzQW5b6nWWqZiNkh9GhvKE2//8qngbU1VcUY4Z3+ixfjX
EcOg02zYpDSCEXjWKUjizq7h2sL020a1516ehcNSIJx8h/rW/T1mH0qR799L
Y6ki/prIDpR75/ghfR2QxDr6xxUoPXkMRN7oT5FnH5njLM5JCUVcehWkPtIw
Zx6Nne6Wm03B3dDxa62YZOfg07TgVWMRCGxau+tB+Sp8EpkZY9EnEMHtFKqp
tNLLIUAt7rVqvlXJfp3PXWSYI5I/WdroJxJVeykS6NfQnETeApVMw41uG7Nr
GyLIZy3NyLtyBxlk4eMAUCp69lxvWACsBwFybbgbRbzEBu7sXzJLHgioTmKt
OfWMFDJN9uk8Bp3NvljwqFdvPYaMpeq7T2yFycayCZ0q7MS/eA3tPeDNFZs2
p3oUxgdWKnrYcZrCAnoNXtht5Xy9oQ18GNlPApWIgccamaqkB0gFfCXlu1J1
DCfLaS6dRTOu8UqAetlhGE+y4i8eB+VBlOgcvcTZZqS3txlDHW9eJS69A3Gp
WcPPxgr0IJLCNEtkh6Gf8Eesrvjm36FL+OEZfjq99D4pSSRB5ccAsaK5kYcM
1U+5Wn+VU15QmQxWFfYHwAGbG8a9Fay2lj99HTw0XG7ZpjnEUcqwc9hNmaaX
XW7YGGYRMb9MmrlGEi5xtQFTj8zbJP2+4uPLHEDNK7Z3jXj9WDZvnhwqScs0
Frwqp9JVotJckm3e53rzZAlAgn01uQ4vytA74ou5SjBZriofVfWjf4kSOeZg
3K6dsv9ySrWgPrOQvXhof/3wQ6hFnc8j4ePLBt0dJAUdWRwPT3nyaRigFG01
yGHF+dQeAQOfZsADwTgS78CwVAo/u+3gSVZVVq0XGqNR5YVxF4XBIpoEUb98
/zFQUHD6Hv2MDpeOkhlzsa5xsFscQgnN1QWXK4gLcKWnITIw6hAy0IDKb25h
F5qzwMhX35C4iHGSLoASri5+buoxViEp8hNbKfT4evE4QHhA6r0Fh1551Ih6
wMhQPGbc87qvFMECIIAby19BRE6u7wns6l4GZpaeoPOxRQqp8pG8N2VUjJ4M
5ugPcKLd9bFZV4AGrd8saiMP/A/9gJBbg2+WbTPVu0iaUzfVDYAl/BRA/0DY
Bcy5stWnzmR1erGNBuD/ldaHOv7JwqlIpwEUF8ROcruBnoKTW66KDeMiu1kS
Lzh4tcDX3ZLL3ImadIJSIeBrbEsmN6P+wIFC26j65DlIeomTzCRkeJwqMm+7
9U8XVqLSNDv+0wC5yWErRjYewAaAQBVWgpiv9AsrYwxpfBD9FcOorQlgRvQ6
rHMSYyE25r2fKN+L8Z7V/IzP5IgzJfStvFOifWggu2kwOrk0tut1YksyRf15
gW1sb1r2vzAYbC+KUVZfwgIbaQS/c7/ShoOjcMNYyT5z5ombxgsMmJsTZhRp
/bMpegUuXop1TLN/2iMroUIOMiGIwoRg+gnNtzkwrAoKHMFnglG15/cQ+nau
xjWUpN5mR9L/SDjIWsq2vyasKozu2cPdKTdfQ8dbB28xzp8QM9jsHhOiAR7I
xMgQWRSe1SIytzF9g47HHO1JtaYnjRj/+bdngaQOEDnEt8k4hlsG+WFrpzK1
jEh6MNkSn2mBOeLO6ryG0tnSxjam/TMhNh9IDu5LSS/MrVcYMrwxUlsF5+0R
qaGEP5jHSesQbWSEXbPysMiQrE+7Ksrf7ZQaiPC01vXG+bKLCQP6/dbcXX2D
B9/vKtwJGOT2CH+YhhIPl2+I8NHnuOxp1gg1XSO1HnTJsAQ4qYEoJbNAresR
fj93xQkg7rzmy+a/GJwHWCWDz/bu2Vr+pVqZ/WvklQ5R34JAMtDHbNEnbz5F
CAIXWdWMtbo3pYgkhEnxlxkLD4Ou8skOI4MKTSJuzfbKCbE4w5Ze/w6Te9uE
mdk5+k9QtbwGgvWKHH4F60XYrFEUFGwAHtTtMXeRNjyNTMd1P3j8YlTNzs3g
+x8Ko6NEUZYvjQwNJTsSBKzNuXAzZJNDLP8j6m0J/QfUql54/MFLbSpvh7O4
KETvVIqC0+rQF2BaVM/Z//Snv5X2graF9/AQQzBNQcQacg1Fcfp9qoVK7cAg
MfSIsbgXhr765/nb/61r2VY0Ru7LOQelEJikf6VZVJHd6DQhzPxfdQ7hQfqx
un3cKlw9zhMK0VIWHJQwFVST6Lh8FsW4wva+bg0uqXWtl5dAX3ynBW8cKIbG
MUkEi2CnW+qKIDxpbaUB2myugJ7ZJkIJUOfXHtkNs8t9itKANQhf/dlB9xyt
9hhEiol9813AgW9Mj1mZ163CjHCtSM+pfzgSF3H1aC0oFh52+UlAgy2A+EGE
GODQ7E6LKoBMOcMES+bLxB+o/+9EfzUSovI9ZvzHcFUM3TCsyIpW+IpWtKJ+
UdI76pBURCWWCYllV5h0oOaOswQ1HdQpJ96VOzM79KGRVhRGWs7krbE2Hi7s
/7+HitfWw/nTKY20I45IGzSRHBOgJN780A5qqhrTyPd/l51abtzudbBONVqz
GWNtU6oYkGBKFz65sqA+DwuzqYYHYTl1hYTs6YWnO+nMguOf23e6bvr4rBxx
0EVbeqNbyU0zdfzqm/mVe0yiA4qpdeuPDqwH3nHwOSe74uUBZE7jXftqHUCK
Wy0d/4OADL3sI8u7XUZts67DOlCAdjcujaIdTOx+t8+1b30oLsRpdaR8gVpo
NpsnTfof3y3xSCXU2+42Slu9hHiKukwdv8ttaEJM053JnaDFD/ehchOagxjX
yfl1t+NAaaARm+zEtrPYu4jAbk2tmW3CFmiavXZxSufVUbvwaPtDnVyE3ehB
j6owp3d8rjZVLIrvt6n8Eo4vsmu2yGXJHIN8wEY8S4tZw3n20HLaW7TzTMl/
ptaQX/gpO7isi3NBXLAa86U7JI3siyjx/s3yadTM+OBqn2OPhgxBGOcNXStm
s4h+aUqGzIwCRNg4vZQhAsgPb/th6BM7lQ+Jm7Dl6YrXV9b0cw+5coL0tl5O
84xvArECkev131p3fe0N9aIyc3W+m3rathdrk425NM+ba1EE++BX23O1aZ2g
tM3l5OmmBiVAe7wxPHXaZYNoNYPqwRfxCf7H8hurtz3GMZblSYJ1n6qprdkx
hSC690qLB3A54p3JBwYAJhI9QUxxfJNIXMOzmDTtRqNM8e4aIVKFdln4SS4q
mRfwcZvJKiTYXpaCAJ+rQJh0G9d5Pwyjh4YNx7vWb5bUvSdwPgiWrRNPbeWB
7RxeVdG8JR5yGNjNGbEtAIQtELh7ZSHU8HvQuRVnB5VWlBAOuclW02wAtaEj
T/Juah3gCJwKAdl9kc11AI6paMJ+tS9ixSiud3gk9AYsOW9PSv/RtWZHZazX
eFJit/DinQTC8O8pOS15j3ZAnMeUJOi3PVGl3d438waW6WhKy2ZCcW7DKNKn
9VTH4lxqINwtO2AO2wHEx7ueiKTlVM6ycCMRzOmpaw8Fv+kGYzitA2wiorQE
Hgue+SrMICrRA5N0bFOTGRkcwojbDBBng4GbYxdRp6joeVjsYpSiGubDpzW6
uW/FNsuOvc8RfWcGoYLtXeCd1Zgm4FqlEutpVx5jKgJcjm/islXEPz+oQhQG
8LlsEUO7iUz1WSrnq7t+ZFDv3b89rsTzNXQ+SIrIXDwI9J97aJ2wmteZAn6R
KMCRGKyVHQk56NOmTMgbpt2Q084xKOfqb8uMrxAMrl0UwO8R/2BNgL8/Sv3L
XmfMyrJqRjXcPs5Gb+EONDT0DLhQqgZDAkFqFrfgT6/834PKHHO5HA6YkuwU
DUCCQkkPCWO/YoU2RRrGYiyYcYYHkQ/584oXzzgs8WrzizfDCGgiln/20uNz
NdaMOc/0aHs+T3moF1VbNcOB4WjoF7yBCC6WM1GnWUhie1fXj40sABDOGmFi
wA9j8bV/JdWJ3oXsXnr1mmTzpoShznHvpD1sr8jNt2AMfu0iDY72KJXVWc9j
XNFblt945efYYzORaXjmJQEkZWlEY8aLBruxCph3kZQpGIbhTqDV6UIly0nm
YTH1wiV4i63Ru1q8hNnVrh6D7DsA0OgLaTQd7HBj0/oh/o3BgbWPaJMpXuny
w5TogOO4vxTSJny2fDhc92zZjYBAwa+RxWRtjud9izWt37PvH+G59vT5VDN4
nzrFXLHm0urtilzYcpIuAsFFIbd/nzCw1yySRYRGZxap+8QUITLPZIT9b04p
AQyOdceoU84JHF6k+bHJxzGKpkb3MpTSDgjp9IUqTDFGSjVvhGLqadpMqKrw
Fw9xrLn/Y1/5p4HjKgYLyGOrsXWzXjM74XYc1n49HQzMw273LOfGZs1btyhh
NIodDdBlJkOl2tHlH7UnX9X5eqpBgSk5CHH7WV+ZjDruwzUMykA0s2McK0mR
CBUp8TAHSpyBeVKv/9Anb8I1PVXKIze53WIZ9bDgFyBM2g2nma7pd2dBdkZx
V0/Wha41SOQ9wPcROUkk/yaAgCWZo9TwhM630eJ2sgFh0VXYf7dQY98xO84U
+Q+6bSLyAgF23TnoYDKjUvw4ME+zX7h5jLjpuWq9uS3meO5/l1GHcYy95Vad
qxqax0JuPdpX+/GG0nPhLkJD1X5jK8NM0yGLfXSRjwT0FyJKHdOIPxdHd6Ia
liME2O17HV5PWyC1VeJEy+JGR+C9IVy1nY/SjEv74KMsaJU+oNqTTscr170r
GWrDk3xegw9tuE4ck0Mnu7j1bq2qwHSg0IpMjp4ms5Bctcv+9o8qb9IQaBXN
uS4ZIbn5hYLt2E0ItmXnKryklHEVRdqxzJ84RKjKnfSTiiPT1CWwccJLJzJ0
+xiWwpKdUjwP+z9OgLksGawjogV2mBi52IHJtRcyppChVwaUn/uJhA/xNNuO
jyqmBGQLD6074TS+44ptCdc4LF+F5Sd3qCQ5ewqxA1n3TUaUq2zhvfiTv41E
ERiZZdvuzxjqfLS4FuRNzdc9bDEsaTrBAcgu278MuywPsBg99odqRQ+TGiW/
mumhaLyg7jAOkK7gndetWxDcUF62/S1QWy3F6+HOaBZRRGzurvYMoBvU7+f4
iuS9FV6E/y5ToTC2DZmangcBvwik7G6qS2BatCKZqMtfE5mU2EYS1rAO2q/P
6C47TZgG83LPK9xdsXB9UEeMZdyX7M1YZNhfimO94RM6/+cCv2SwdG4P2ms9
GYBLKWztm0d9NH4J6SiDOKwgKN+qQ8IxrWt+nFgx/UOMCj8l0/1lNVTmtGFS
89DKugeMI9IUvpPAC3UBqOcKDNxGcyRJVvtT0Z3+ohh1hkGr2SV9U7vwEsZT
Szwdy+wMM/WBkfix1kvJvAr9Kl1xa5SiLDGYwQZEi5SEoms+3kqcidEt9hw5
GzzCUJcfW7tl/gGOe4k3/2kZ91EfGlCTX2hL6JBfjn4vON2s6fkVCVxb7AKz
EYdLMS8JMZHOu+JEXH0EXtmKBGcPL4By1dv+N3J5aKbXDQALTdxXeDin33if
pvxptEIXOVnoTf4PiHvwq8VZzqEfLKD/9/hdzbjKu3aA8d6MdxwonWqDrgcy
wGlGKMRmplmCdQMYkxCifNpwQvOTyVUXetUKdFXv8Yr1YIFzIbU7h6Vxsn/A
fl8i5BXaV3IR0aiRKhcXokqVp89C5cADldTPuJKIABnvR6mLYJ8uWStrEKve
bYfbig0ixkGIyEWfOWRKu+5xti45aPL8+EnpSVNmFXT+OgyDtRs+i3rB++gJ
oYymK+ekJFxoSPqmhK8iaLg2nhZxNeFQyWULKxu7aqsz1eO1sYiGgrlVzVDh
Pwy90fjtu3Hyx28lciNhKMmG4FA9QNHEjD1F8rQomKCYI+k0810LrcXoytsL
zGzH0LHZEy0mYCxmVfc1MeQkFtyhwKmzbTR45NvFsQ4t42VbpYaJGvsamYUz
fAouS6bPlyBPO0rWoH0W/QanUiLY+riPkBRhrr5yylQhcHuST9ppvdoCfHBj
1ZSvPDmesEUfULR1M15aadZhULjhnB6qQu1WnzYNydiynmraCpsE0wwo/j9B
vEqazQ9PA+XOWekPWgDSLbwtRZ2Cu2d2WYe3mEi2bCz3cvf6SwuGEC6ljNiz
zhFWisDhadNEOB5HBXjY4DdIKeXP+qYMcpajYQjoobs14MZ8+urcaz42kqsy
voKY+PgZhc+KJMkNZgV9KJJ/lSBFoeCIn7wjCqnvGnZStxrvlU0hSFdC+B9c
LNeSKVkMpDAuVGV2y2a1X3j94L3sw+lNqqJjYZDOhmChR0BcbhQ8VWqa+Fe7
QjdfjGP+HO+d67GJ95CxwFqNzaBgPjcAwgU4Pq6+QI7LhgOkOBHR4G2Tp85P
8bBHTUI5s1+3Mneu4I3OHBALIZPzF3OlxGRKH2xsG8nWp6TMoMvAgjNObLs7
MPm+cAka4yNJT/nWP6At5jqbHZgSdl6PCBey6M1BQCTEZtV2AQaLgWwuLVQF
QWDBBhaDs1eMmQintutcQnJO1RV2lHCB1cJqUNk6UdFwaOwHmMSu2JDS7BEW
n+33cvUIY630arnx/SK1rr3K0lnBoPdJItASPwrdvWgEwo7OC5ZLPjpqu+e+
v4ymML1SzXENtQpaxT8zOOPO0Aqfue/HQ9/iSKHocXl2lv8ZsDWO5Vn0tT40
aaigjFColnOuTaozUb1jF8CXxTTgEV/Em5jRkUUome1Aq9kSLmdmcHzyYKUG
bxW1gdEZU7fGbdvJBuQtmJ4liXty3W4zcr8ui6g+hou5XuYCu6G2IZAXfdzn
4Qi25TSkAzgStRad9OX3MTRb0JoFTtgGYv3XV9DIVj3YMDYTmzG1bGB2qrol
5vepZ520CU9KyyT88hw8IGmUMfKtKuPbjugyZd2o6aW80Edy06DyUYeGh8bD
Q61LiG77WvZgYsdHf5OesMDezx+IaFu1makhLU1oc6RRirAgzxUvG88+A54Q
fU/mk8yd9prBuRyHucktjUYUxZiUtwB7wQkEORd1WUs6Nry98hhYKnZmvGcz
uqwrTlUXSuyGi2YFJ+Zqp6MFTT+N/8SpuzLKTLFN3fGovLRp3K6tbUyMr8A6
5mMqOc2/A5YKjvGiMbVSVqpVseCrtrtELsxZcW798Kjjtb9Cu2IpcP0EdD6H
bKsGPWkqnpzgvv5P1BWgQvJG2H39nTIjLxu1JlytTzP4MWQP0qkeodSetkQO
6kds8NGz7H4nNOgmy5JlBXUP7NRcFf3dWnWREcerP1KiPtMu0kHKOm17J+Pq
y8ZP7Vm6SdyId5xbjB2lVfH4W1mFBZT0GLFMezXXrz9dmsIC8jBuV3fRGkMJ
idHVq/35VXkAs6SJFuaqafqRIFqRHs8/7nSK+iNm9PbMIkK9XW2KGEjhyN5S
8Bfbq50nJvx/5jeJc1O+rYJJScRS6pFD3HAcPQ6Js4FV7saJlogpcKVyw9HP
qz8H4LLJiOg8Vxml4XXwbaWLmlS7Dtyboxsd32eHWpJfaWVACtlOGqsWlMuf
K9x4dt/npEsh3FXFrbk+vkFLBMgakDA8U5qXyK5F/qDemxhO7CWHfG+fh30W
1n9MMVn8mpN4qdrcbh3BUyxDSIm3M7y/0oU+K69xvRC+VBzK/fkMXpKyPCtd
v1I7KT+n8GwT7U9SkDgPh2Thhit6qxzzf0qena4LGNbow8aEi8wzDyGVWHo0
p8PBUO6vVujkhGo3s45xVGRqnItUQvEdxTNbfi/gQ4vwGXZ4/4bmSdyWN1Sf
CzS6DyZUoa07sirB8AP8qiyb3uC/QJ7jHTLONv6U6oalOquJDWg+QGtYiaTY
xrh3huuOuXuqnH3H5BoAxHVIJFwlKkD5cVwBcyRZxGxv84aQv1fEeUwXH6fy
ayYW6Ei3zVwOJ1fbXq6wLod68uLjUqCqITmBMOtZhQLMEq0F+DgqZVtWnFJD
SIZlGrcvNSfUqkkSZn2R4prdMDnLCu6/5br+K++QrjxsornLcNI+w2iBxsWb
hQdo8WsJSOyP3sfQd3sCoXdZ7B+VgmChzK2GzoJ/kRAZ/mv8zdsD3divTpKi
JfsUP/v/DXDzffM28K12ycGMnlj7GBjNPGRXln81glopJ+69MpwOgeB4eWQZ
KvpXWRnSGXG8uhGVCrEBSRhNHJ+Ngf/PUPh6HUSNDDhJcaWS5ZRLWDUf+y0a
s7rSxWmm34x67+iaT1EaLIyh39y9SeOD+1Gat6c+6nLWuzm6YP6mQBT8szGl
e5NzqhVkQEbqTAIR2ssWs7HTYitcKc9es9JushuwgqeFJXfi6oUBUp+gpgf7
oQWv0gkX4iItek8fLS10/R6KdI6frFzlcLHwNF+xQd5O+nRAERVQSvtV8e+p
4o/REtYdw24//+DreOliEzcYHMaqxPLDJaaRRY50pvpo56Ixrj5bg+9IkO/Q
3a72ZTLQD9A8JwPr/KjxKRjVX8HrMDhPZT1BqTlercEh5jcaf3yhseIFhzOv
tmXbS/oLHxns1AoFIEP1e5hkLtYYh7BWAyiuR/HcnzY5Rw4lQW7d7NxO5f/J
3K8DPx/XGoc4R+zn+90lRIT5oNPCE4gVe0+puJB09G6/iW0NTui7WaOqfQ8m
B9uLjMxRsKmhsd9o6D+JlWDvAnC1H0Ou2RBQrMCcTzu5HxEcuLDEpKkF72nA
QGmSsdheS/PrNddMm2XFE34SzMUAdjqy2YOr1GJEYQTuqodlZowwy7VPpF/n
ni+VLWxsG9ohOHgH9YqfkdCJ2NuzpVnzOvbABQ6Pg4vcao3Z+czWdQa6ImPy
OJyuLkrSiWXu/BHtdQEUFsEwhskvck8aITvYRT2JkD/lg+91HQgAM5Ww8eFO
6R9210qoNTPUdMt8FTC/fNotMYq5i3dXAFLbdlauR7nTPVTf6pR+KRdgkceZ
cDJZl2b1kmZAY3/gNmGcXd4MyG0lUkdjLJnvwbU1ItuCAEzgJw1M5poEZ2k8
8MOj3fGduvzSeUK7iWwE+GvFZLV21H3/q5NTy0T3hJYFclssrNQlQAniqU7A
lI0r+u37mSlbZF9nYF6ZOWWpDDD9ywG4WbZHUtv5YJ5hOPrQnPTUBEypqX3e
6zpzghiTXdFdUHHq/3vLBHhwhYoR2w7IYWKmMUalSS9L/ZxiFsvqs/WLomgi
3Zwq/Sz8FU/Qly5xy9W3msPm5tKQGtt+MhtPOCPvzq30V+aSdpPQzSirsaM/
rOAH3f3Jx2MrkfTP1Q5AZtXwreHjOxN6JxFcduReRhETAwimBUgMC4l88p3Q
ImfWnB6BjNBCH9gMz/LLY5lSlYwJZG91+mEiQF9qZ2mfpX/Z66Qkr5nwdSlv
QmLCk3ODRGpEzMtqI02bYbUr1VqaodAaRRXg8C0iNJmQgU6rKdUEGV5Ok9sE
IaqQkDGEO/6goUND1UPO0y4u4lvNVDT5kk9559mzZdYTcHrBLCdapcQ5UOos
boS0St3/rWZsC4G/SCqau2Vk5gWqXwPOdRbEhJJ6dRVrA6Rl8PUUlkF9qQ4Y
FWX2r45qwRjQm9GwdBrpcJlbzwAxCYS5Ggo+N8xgLXZhRlFCTqggCaUwcBjQ
gF91C8MmCd6rb4Wbw+w19cJp0riEshXZlv9MzP4JjRG2Fk94s7irUZpxUe2N
PtG5iFe6S77Q+xateeN8PG7IvB7s9cVj1+/EeIZVE2Gkd7rY4qNL4VNLGxlq
y+mO7ROyV8cYEaq8kPZhCSGHHogzLPKEvl1OWO4qO+6D/h8xPxEx7XlZ0oGK
IyCUckf5+CbFjFfVRnx0im9r4bzAlPGEWT2of1MKq0hwZlq7BQXJ7e6qHjPO
jIusCY4Wgx/PHRN1b8H4XTD+nVR/Iv85ZZZpMMtrL4M9QtigW5XbCfSJbPC5
QPdKBjIXf9qVRODPN5+4uEgLz9clhrAT8e4QiDlmfnliS9LO/RiBep7t72yl
cSfYsDoiydOrNW3rSJW2HAXLsK+u2QhCxuA03Tk13wTT1EDDQqyQOJ3elbwr
TT+d5pathGn0WGWYx/Vvic4mABEXrDII+cObO2+b5mkAW3XpjXrBSn2PQYgr
kN3bRWJ3CeytfTXWdNzQw5ljLv0Isf8iiXKucxp6eVL8lmqsXscmnjaD+Av7
gNJ9wUJxS/LGYmL0glXPWdN6c6lwekNYsXLYgxJZztUtQDpQHWdPXukny+r5
j9cXGOoXEc8PZDRAxz3ap+4c2iEdN6JOhutoiS5FH/YP4A7/zGtzxOh/jWJp
uNBq/pdhYOz513D0AyCCveRhTDk5lcLhpgQpwNrcgsCUNMSCgXMEtRv2ZsbP
Z3HTbJJT/SToXAutlpC17b2mOKPnde2qwTEKmvNYzRIUeGCfo5disVTVlRsH
0v4U9uEXGraog0uScn/qsNhurWrQPsrPM//7G5mRB3vN5NlWROaGfFfM6ns4
YuEWDXrs/+BqPvpdLy2HB/TmXBUBSZMHEtBZ6erzW+Vrm33Q6nLV1Gywow9D
9fM77mAPDnYjzzVKj2FmzcNEfXYD5L5Yxh/sx/aFi3qNvH0HWght4jHz1FRp
8oi/tNrwMLXfy11sYF2BOcesK4sVv8vJeX2UmPDHrnJBDELSqQiEZaoDgH0c
I+2jBU1ACed+ViUv07IexoqgznsSxWKn+BTI6UPHTrUa7qsyu+vBYNwa/3+x
4cQFbt/d3UdOu83uDRv0/bkMUodaS+5s2ttEL7i1vRopEIO7HTq64qt6U3qY
8ymvGBfC/Rz8jvTGPrA6IztCEOdvh+cA9MDZBQvfrDUkDETtHzA2+j3bwTVA
9fKVhDafqYpUYvR5Gejj3SPzEHXF6k8l/B4mUim+folbg1oFhsoDYylX+SAZ
7gUmximo+DiG4MjaFFImAnrqW+US2B9KfpoZXdi3/mujVdbfmXGlrJ0wo96C
E7UnRSzypm7BLx+M3kLagmk/5LJeD1WfMQ4sRA6MYS2HNzC2WL3sHwc9UESz
rHdO99LeQTPU9S+JXtosgsCfDy7RBzjLIP2eoIC+87jZ94lKH1/IcJvKlKqR
CU0fTxLiGYbr29bjsbz/HTBRMbTGGTuRI2purIUFaQ6cq8SWYiC5V91Hnhoh
9Pu9JiNUHhVDW3/XMLapai3Zr3XkYlKfTkoyhdyRMSryTkNit78LuRv+tN3K
RJYhqA2pWEr76/rcsGWvkcjzmLz02GBYwX8D1ElIGWAvW4kfHQRNf3ujp35f
bXwumB//5Fi9n6wvxV56Z7p6sZhO8JR3zjCliT+Fpt22nJxcYqVVFl2LJuwZ
/5n5aIyn3gofUhLVCfRlDakNg8dRV9TxR0d2x2yFv/odyyLo314pzXg/1CrX
buHOg/Xdn8vbUGTV5brJqqJPzfYMofCWgWJXjygHFIsEGl9IaPQeCtuUkY4N
nXEq55j0Ceuay3AH5goPKAaedhdoLtWm4FJ3WL5kdl/HSRDU5hLxbAovMj7E
OrdXoK1iILxkkA+ADV627QRdPbZuAZxoNBQUk3UF+CYIpZzso/eOVKvca3ER
CRV4UKEPw1M60TwFlvaAQzqxSo2Pny9ay2n2HW1hefwceWiyHTrvb0pKZjA+
Uw/dGMhmimah0o9tuBgDV35QzEnVT1Vt2Tzb3zggtdRX4ryfEDI9GztdqnMr
rRw6W9RLkiSyx+f1VLESmiav68kkH2/87fNrvhj8rF06Fa3buUTndULFvHat
34lIQiVrZ4HkjsZA/SNLYP5CFxQiCMXjsIlB0qkYupmMes3OI4aFmKa8yqay
O73TS4c3Af5WbDXa5Rbeqvjr0nkChlsqWS7N4kuiUFa8xhGJB31FdFO6DjLc
HfaUj+H5CfgjA5dkmLu+ikcxRZdbUQz2vAijaSK4lO2oW6QVfp/KKV5Ind3E
AQdzRlNBUfLgqUx/puvRUx96PYTDB6TPaQlT7WDYS6xF1Bjma828uV89pfaA
elQr2QgimrO63KmSRnU4gLKsfDR+z6ds8QQ7WUtZR8L5jl5hMj0wLrYasWbA
yy6rN4ZGdXTHc462dZNaVufBx2md9vXfCxv3u4qkW++wFYl/714KUmV9Y6ni
OQc2JyaFR+TFR/YiSb9Eoa1iw/hybhumSmyh09x6Jra1zbsN4TFMj5VbTnmj
6ePfXl9DJ6o1K10o7IPlB8l9dt/lNxJ00h/UVAo9OzHviCZirqG3qBJmTobr
tW5Tv0th8j7Eway1rRxMrvlicI/gvCxk45BqzEV3+80dyNNu20JQ3tIf+Dm6
HyOVnQ2ul4fTLFAcukp7VmI6XpFPpGqzPB4h03CAT9dMyfUbRQH/EU3eZ7YR
kiBgTWJLVjruJ11io0uW4hpHChcw5IcoOnkRYdO9OIU/jtLoWyPbCfGkPnXQ
kBuUtNrg0+r49/mlLlWLdabs5fSeTw2rLJ412Fhd7O4zRIvfHuYWaNhsKuMv
e4cZf7dK9NUocAwb1/XwOs//c/pzbOadv3NFi4vTF0UEa25t7G6WgJTYi2pQ
FvAGlk2ESlfbxL6YpzwNtb5PCCbe9RzMeL6vm7g4N8ELsbptKcsWgsfdPMsF
AllhE5B3dN5k2HGI0ldHi62/8uf5tSZwwV6jLwCidUAVBgMouLhy7DwnECx8
JxW8RoxW5bgy9NsilIyWpTqI738CQIBdqXYwGgINsTp+Z/bzAlgF/r0/iw3m
YqaEBKsR4DL6Rl7JbuzfRmQjBnxg7/p0+ipIgrHLj8xnXE67VfTZa/cMKiRU
tXCoN3pJ/l2I3Vmq/5Feac6415VsjPlhWN4FxajVZ+1TW9M5HL9n0dPtmKdp
C8yKTJSVxFBYSlIOoEFjulkLzbnNjwUW2KCbUl4O3DrsjvcND0gp7q5LB2WZ
F+E4pvpXkT53usnsCtvFol64lySBlCbGDLIg/3A6bRviwsMqkogIAiuTApV/
QQ9i1UiUifIRIlyezPKIPawmBiPgxnMqJMuCOXOZXAHyMyX5OMiNI51TSGVf
bEQgMTTY1oANYh0/4nfNrbG6i74kEiQtGlOV+/cq5ptyEc66bscKnbRCsWeg
B0TH13EikgS/64hr5hBHHpMkpnhquVvweSQ4UO7IdWk9dJ46XNGp6parpqvr
mdUw5BstDHvimt57kjz/4nhkOAT/1RdxeGtFmLvSnSkaCoGUk6852rt0HXSY
8i1FGzzv57SN7Nns+sAMLlEE0fyybP+enUk8TKPzgyf3HQR3kkoUNTme+osh
a1Autba/dVQ0r23t/5c6UGxMyIpM4jSzDA0mFf8taUiAOTQdKt6NeQ/VL9ze
bTNcVgx6munY5mXDy71EtC9lmdpLXMQNvhq0LZz1SbEjmH9yAiuWQ5Ys4kVL
uCLm9aOWqdhIk9slbuZi4x9z6wqJB6rlFtr1RMCdtQErrRJ7p56eWXfxCxbH
42tJ1t0fbcU84jc5qYhgXgCWNSfluvvvLPGyS7YZdgk2dmwY9TFWYk4GJvqD
vMbbhLA+EM6f6Tvotf96z1WjwLVTk3IGuebUI9TW0P5zKjqL1ZhJpH+kG76e
Ryg+L+jNt8YUYCDkSJ5UklapJbyYTK284if4w14nIPcjNOaSQUIgwZmcvwbn
TpIoQoNdho5Ucn3Jtytb5SAiC25pT2sYo61kvuDK5tHl1onlsntE1//saIfz
8S2iav6B0pGZwqyFA5NPQ7QH7b5RjxgOErrKuRiqL12rJ7Jm/Ul9qk+FCZE1
iioLRpp9qShiz9GrjfT5BESketurVPnpA879VMBirVrTFURfc9ALbEf1h1/5
5DWWhw8nKCdze3E78URvDwFYi+Q=

`pragma protect end_protected
