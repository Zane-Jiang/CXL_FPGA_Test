// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
r7QhBrYYeJN2y9YSxi7OxXiWEtVvDJxZhDBMWwW3rR7y3S4Xwa8YTvIqWV175Ofl0S7wITHpD17U
XvsrCJyHWplhyn7ZwOctMfFucnXRLPAi58vgTWjdR1PRkx0TnrrxCZMo2wcIIj+VNRZbWxsu/mky
xHIvloqoghxN4Um7zYm53RfU/A6n10jzX/GbwTazwkAhHKyMMhbe3SFys2Of/7A3YpY4QZe0XVzJ
1j/d6Fm4uo4cRcw7g15uSYYHQltvwmJpgFhsCjzQrbOOvZyZkJkRHyCCXxFXnltzsx+7qEV7yLN/
eiatLFYdicrATTpljetuRvrlkBSiiz1G19qO2Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 99808)
nU2w8hd73+qMcdsk6u3KqrkRvAA3ocTfZlqst4gBvd9kI1qluKjMLSL5xlmnDhAQtDwKKbzd+ce4
++vncBztcYums13LoDPIvW+Eb4dLSJewzkC2rfhpSkXSv8X2Px/moF6Y6YHuOPqPrbNe/f4xbD8h
oQwKCwJCrs90FlQQBKz4UHOfCfo8K1v1jFJ5tteOo3jIJGSOGYtVlCZUo0gN6Rb4oVELUfe8qKRi
ct17SnTgBpmRvLo0siij84nimP6O+PZ8vGF/WWExWR8ClVTmf6L3LZZ/+wRgPXOYNe8k6l5tasd4
vxfVlAZFMD2Qxy7XFsMUymh5Gs2V3yXKJC4yrZptRLNpVpFr26D1X0hK9mlMpHij4YEYvLs3ZsMY
H8pxmCUIRoKy9lsNw/zXp9hmlYKxsHEw4tyUDnhy7JKBs36M2st1oq+DFCJMOO95WN0kmQjojM30
VKGJ1Mvi4S9vvtRqWP0W6OOke07T+j4OKOYMn+dQwF5hGYaRpq5A9bUEjUonrjKKD3xw50Z6hLur
Kmve9AqDHJgUjvMUmAFLq44UFYLgnPg/DJAJMc2hc0uXUJaHDiz3BCyU8W53+HBwrMIwKxEOVRZV
f9S0DjQGrsI7EDDiTFeFoFQBLBgOeTY3WMCeNObf4UtFeES8bZXe1RybWmeVC9vFS66kp2FGEdKd
6FfkJnBSsPGjo3jq/tKOBojtTquw1N1u5O7/aX7spq/5AQfUVTcnzJDNE8MJ81S/z0Ku+/hGuKJz
bWLNL05h3Or5F1eTkf+Z6m+Att2gUwfkSbYk6+PBVRXr+L0OD64bYWAkpEMJ/CyfmcdYv7at3P+g
IWMIMbFZ528pHMNWrhzQ9JVAcY9xmy+wMpFFe+plmS/gFDL8pXtjbbZySwuY788CnRBb0/ZGgjdo
IramCMESMcxuIkbadkoPSg667SijScXLcyqBClQMPyAL5x/g5JSdwNBThR1JzqPrOYPXe2M3M92V
VebphYD9CVBcgU+/jCxdBGSxbGdfX/q+ML4Vo8d7vp7cTVjxNuA/rnD9hrt+Ab8YuKxstv0CSOHK
QGys5Bta+rFSb+pg/5CvDuEJJQDXW2ssFaAPUlGFgCwLVQtrUTPZN+SAb/kWcJA55Ww1jYNx2Opi
bSzzraNeyDsZosNDY1oeP1YEK0kqttSQgKXUi173NO6IiRBVKW0DfyY4Odz5EuwxL7O1PejyACr1
SISO/5X3GJ5ToFQozpPO7S8EBKuRjr+/8FpGZfa+u7/qYH2xev6gJRS2oEbpg2jF6O4q3QojD2hm
hsJhrzgndnD7MfYn0D5kAhX0WYWEzia4YxqnwpronfXb2esVTnW/5C9zwJi7HhJyPZOeBttXJIuu
uD2tCjFtxCBW+ocqltw7LzlUxcDu4DHAwYHsHyO14jAk+CSqvcsGL7X/Fr/NfPJvzE+7im8ohQvW
Z22gf6BKfQJ/Dl0JpDeEOkqwhI8N6L4PGH0df/bKL0CjEZyX6dBJqJKweMXVzlMQwprdtJZ068rc
TuKUevFFBrOLAJfDJQaAci+tl1VcYTXU9FYgYmi04azWPrZOs58l9tvSfWikYjrzJmsLqXZuXbTP
RdEa3n4u87Q6UnZo8BlMZbSW2mef8OewHLte/O0xZvIWe4bO6uBpbfTSHvL79nh1IXDBbrYJFuDs
HXOVRxw5qKtb/IRq/UobyXTfRSrqN2jMgJVKEAxZZJzNHf3uOW47ULBCsbvonqEXwCoP2d0goiNk
e3wiRaiTOcnolWdbz+OHex7LIj5JiavguV/3zx54UjLdBRoM617bpOs6YyA8Wf8h2bv3pZRMNxZI
PbIuoSYyk8Klx8WjxMzPN1z4Yx4ueVJWLx9E8jvSSbvk0tpQ82bEnaXtNmO2VoWcRWWADhK9GuEo
qTB/NOfHVl0TY9JbwQbf0WKjdVXym3yzELmG2PWY3P/KWNXoHQZVDqzPtiA1qpu3RK65kvUB9I94
/N0lXdayuiUIOPbMBDjtybKEM/MyB52PPii7Bxxo41rs6zTp4RP09qkI0QFWPYtwjrZNs6qAKs3X
B+29g1I7wDmOmf4/Oa4LmrAqWnHRXaDlz8Op9IQUqGYTkCOT8D5s1Jnp0MhwZCBC+P01v4ijZJpN
6pEXPa3xfqMl+nsDT86XCxobVqdfaPjzrrTeoicPD8vdticA6PAuOaeu28kY4irES94+FV6xFK5j
RCQKlCbstgBXXi2leWeT391I1rHfH4wvDvW9uTxGgFJP83EcGmCy8B/yUXILbdq6u/x1EIvSuDF4
X6rSmVeYqF0UUITzP5PiT7AbbFNJEIHwozBybeuPO10AjLEvagK4M8sxRySZiu+FpIIBSy2xzrii
/SNueYyfw4dkAN1qP8e3tSkDIVZ/r47n7rwJTaZGDf3RY4+kaAU2zBjP7p9XlJ5AhHnAaaJl8HJZ
e9G3CnbiMq0TlHhYCMI0YE/YKkOrjMi3S0+vhzTmivicVsjss7Q7pbPfXZbZFUUdtWubXctq+mH8
sh0Staj9GwKqrAZ4Dwk60jYcUxtxvERj+ikvDaEJLoDaRUw3OMWoXeUMJB5pY89wivb/a50hkg9q
bHWv+Mba+U5hSDmHH3oba2xah6Rfw4q7tHxcqTf7tcJhG6dAtkZIYa7PiceGthwLVET+kHDousc6
JEPFEEHQp5t95mmYDPuMSdJwPa/ddLC9H5fkvp4nu5kOGKW9qY4MG3YY9+cMJs0KqUqQUfCW/2I0
Jd7zgoaN0w3RzmtavMOfng200/078L0lL7IWdfUdR3yt4YdUYLKCJmV3PFDwNZ/rvwaBy52bH8Cp
O+06JQgMsVGgzEr381petSJ1EqY3lyrbFn/9MFXxkAneq4gXnzWZKOL5LBRtS790I2e42Qs53BhU
KSdq8uni5NgtqMMFeU/d613fB1vD/uMTqT28eluYQxmG7YYPNa8bD2J+9X4+kR4H3bX+CX5D8M+1
o2fAORv+HSJ+5lPn/Hj/GBY3XH74kVD0iqEO0oDPAhNChcnmfyiaYTD/BD/KRMF/rCfyGZtJXODC
MKj88OpZtPbiBBDqOvIdbGNxDdGfy8WHvFzItBRCGzZziqU/ZdYutqVVkTX3wIccQ0++gWRw3pAl
lRti/WtPHxgGBgMlp+7PPe8TauLtxUH+n0UZyrnDmmnDBw/OrE5WRNgFPW5p4yrOLXoQfHJfIWuB
qwCTNAvlQoC4SJlX5HQcZbO/a/Qjsy8/9kNIY7cMsAzGsBYnnTa0C35p6euQfsmXIeoXdjRnENt/
9gyMM04kK/5ycr9/vNP1UbHxib/EPL8aOS6LGXGJhzpRWEiT3nNHaaQXBaW8ZSkwHxJ2/dLHyw2M
kkIozor1eMGHEVrXAXqBBiWoZdxlgFQuLivheYGyciAigu+vpDm8DXGpmqqdoqLgUuEcXwDMTHTt
180b5a+FcF+Vwh9tMAMzR4tYd+tITXAt/+3+dGzJSXjk6k69YH46S8LNnq42uY+A+rjItenFKZ93
b6u1762CkhSN5Z16SyW1E5G+XbBeZAQm2DASMeie5hygFCY+HPCiVWEf37uvXLmUHbAOZMCHaB3a
ZCYx7bH3g5xCe3n1wXHQcFFyB182pwMXdK9jbSi4DRqis8x5og4j1x+LpaPYP4Fbrifxxem8SlJw
tQIS4kfrDiFgewxsTnVlWEcc8PgiYt3TkxrW2fTaHCla/DYy0/Oz872RI7FJZZ114I1BwrCOzD0b
wnXZNHekkxzFdX/cva4AGcVjdxU1CNOJ70Y/goCMvsAsOcAk+grJiJOY7TM96nhSAuWgy0jHGd9m
6DQPdamwt7K9EvHKtMDQs6tcdkeYcAa84lbC8KEyuGyhZezo+DMYsyocgXjd5H6rJape0876DJF3
1A9IQO5YkA6FBOdSHMHNihcwLzS0hTQNG1+z/SEZlRP4UfOTUSh+k4aDipbl1wIsihlHQBWjlwTE
hzvsUzed3D83ejIoASGoCj1KIjNVqkfwpAq00I+2lJcHBNspNYHEXwP8097wSb9KDpfb3vynK6Gj
vaQBsd1uXaRm+P4yYHbPwGqXSwd5EPm5R0CT4tBluyI3h0AQk4BTHiRpIvZIjPAdqHkSAuRQSiuL
QjH1tfedQUlNyCfjKtUpxB37swdE3x6DE87Ck0A2dUpLgGI+FahMlNH65pq3vIxaDm8YwRiils+i
cr8I7F/PHT5ud0OC4PG/pwWG1ZFmxHuFSrQbW2DBqEt8cnQcYVTaugN2f1ysW9uzawGJ9uhjV53M
ksT0yJMMXh8Tbk5oJybKTUywoV0pw10gBC6mrKlpOGvDDk5hieTtTruTBLzAuISlqYrZzvEHclBW
NMUgS5L3izjpvfzgFeDJCsyLBLkCAwvlIqvFdkb0+2yIdrhlucIlzbEH1uuVC/3B2trkRof4wTqg
rCs3NbKd58Es0YGuIMFgcqf80RgB7OgblxMVXPG0jOxjwomzRWKgrXXl1rFHt67nI3+3opR10QGh
y3ekHkCK0BUjsx6/DRjxaaq2PkZ/v76asImeSDi8Mety/n0bBOC3mZOl3ZXIGI/5n8+S56riiIzi
+VSadJjeSSqwe1MRooUKRUPeYaDCROKkBUFbkGdrxQxECYIV+d+Q13BFcV/xal2ysi3jmiqZawoN
fYCkt51YZ+eFZJ2TcK7imk/KYsAxiQckAU6+CTQ1JrnFU2OAc1dE7unCIGW7G3+QkJFxruXn0LSP
7SaVQL041svkt6oNoVf2z034/lnemGVcuMG4AGcmDNP/3CLzYInAuXMeGDooPeZIHyzCEAEvxs6D
+u0v8OhYYIspkV/VdAzgbH4LDVINJSmeOMCd1VkxNStVBPi4TJoxmDBLzcjDKg5RmZYUkF6Yxu0P
Mxh/gJoVWZ4U78CxYPm4pJ7JAY4Y+2nblOrp66qRc7/e8Lj6crc6Z6q9YW5c9u5tcUxBxdlShi/z
U0gXzpb07fwZU0oWhIcT9M7fCBcxj8rI/2czrobzcevYqJmKGmuRaX3wmQWBm4GujRavjCPBNH1l
n3EldNdeF3SPr00BRC4kL1JCWQTMb3spG7lj9kmmlAmh/M0IdeyppS3mHJCYYcT9mYc87MOuMGwX
q7BesW58BttkZkgKQqxxIGfJrpTl6wUPv4aZjcXUVt0Ph10u+hRKDm3CkDsO0wD5hiUfIpUwxMK+
TQLBm0Rg4duMMHt8RVa5FURf56RUCGBzVkn6py4UnnXOFXgDIAY3EBnvDlVLBYEpMZQwwv/nsbRb
HaOsZmFaJBYB2l6yMvWKmF7TxTJ25d6Z3+HkYds7ECPWdNlwpZtjYd2gjdfAS9/7IDucv7Fghy2D
nb1P2iZ6VEcHIL3N6XTEKzRA1WsIrOpcleT9RuSoeBJOoJA9akPOXLvvPE9/L7d+nts+ki+dEkc5
ZIarppOpGMuw3H7JJOpkXvsDqlRhvbr6Hw2dnFZBfR/7gYpMcq7RmRzyYF2avuHJvj5ZKjB6fk0j
J4r5FPVla1S4zqiFXtLYBnLuS3pQaUJZhxCNeW59RNcR9HX4dQHeaYBFfzDQwAfgiP75kMEPfyWp
Ay8Zxk8oQbtTKsfRvX9HEAiKBZHEkRdYbvLFw1FsLwxeTWCPXh9cYOJr0iM9waFmEDT17z4kW9WN
GCYEZbPF9K7V3wV0UvJsaIy1uuz01+1PeFfnTz0mg4PLjXGBPFbcNvpAfEua7tkNNU9WnPyGykoY
Xw8st1sK2xh/j32m7XVd0I7PpbZZmIYWF5uDiKs0Gm7ytzdrfNFzMnJXOlE9L5L7VbNPm3a2npE+
P7IpKgHGikchM5LTfKq/IrXuG40kr1vsHZQoLZIrZA+GKmoDh28JyWHhnHsCCINuReWV49/zA5ep
QiFL6TtLV5GpBP13+iOaD07mA1xEWHp9QVjoAqMk8hnmCVbmTXvyB/9KiMcV4Y2UxXpG540JBAnA
qiMVD5qR/BpWNAe9vEaTzaJGPDiXAV53kY7bK+sIa5mUD5LP0UJrjs8H7RY514ryAIuZZ9eQoJvA
JxgshpSKn0bXjyrq0pVOszJBhYzrOddBm+cKCFnYOiPP00PgUtjMcofUqc/4AKy3UIznUIpErDRn
SQYjNiEh7FyFBxm1MwEH0/yi12hAOmR1x/ryq7nqVvY2cK6HsFrvU4gJlFxt/fAApBi1QHUrQ0Ay
DB67CvWytFCx/IKwbwdtxCtH+UVcVNZWEchaVHmB9iJMsL+ewCoczsTS1zBMdj4Os7D77Y1JjBqZ
uXY7d4kvJYv15orYteuLNLAcdwVRGpK+wiiXXQF68RBwW9gR6/4ciHHGBcUbde1hPyQCvVv7bRgZ
/XnNhB/J8e9ZVMepfGbUtPsbdWzOQwO84hADyyB3aCDo5qjzkDzuxHuHwKZVykAk5D1K1yaqYudQ
hhISTYr6ceymPbZ8QY2wt8vkGDlU+CflVEg5sQwAXL6NhllrVkkkTm5HwJ8SA2Qs5fDwA/7glDSQ
i0MZfE15X14uSsiim8rKbKJ0ZdK7sOs2ih8y3z6ZiWanMypRIqWySKyijBev1GO+SBSsAUYX8ieP
XTfheHiKaQ+rKaWLQgE666Vx/nvWAFwS4BbyMGtGa1WGY0bBdPshjNZquZVlUrSJM1n5V3wg7vFT
1ngwZs7Lh/+YooLSwKmhFyVZ4007vyXcZtmpSgJAlJV2AEJE5lYNV/qZ12XWIU7oJSxhfodY005M
jtR5k2txFr4VaUGh+00iUjkVuBam+aybKP4o9i4Qy7MMww1GVCWXtdfIGmG4tt5AToXUGy3eR/nc
9Xk0bs9p5rYtLlL/xRrOqiTO7DTlwp3mZ4Ka5vue4kpXo1ZL/c1aD5d7TXby+B1oc9OaQFfSbGKK
CF7iW08syfDQNH5MrN7tEPGvRdUMClbIoH17NfeRX/FmOTzuh/wZ2euXKil3QS66p9lygT030EBp
evF8JKMU2KKDsifuEz+K/sqygQNSRukMfuKj26VW2TWdCeYE0WYhX7Nkyfoj5nU91m03B8NbqZzR
80aKM0J+i0w4UTLD05qkuKUbQ680A68lzDamxb0A0auokglM1TaoJFiqyaU3lo6RLDjnb+iSb8Ke
hiWkc2czKz3aeGD5n8hzBjZen60Y9xJdupDHg54YXXDoa5zBpK2CYrPzNVe0PQocUFdW6gjUFsz0
PzJJImjHxkOmVCFKjtGY4Gfdut76ghHXqAuDgPf0+PpBWwfwmMXHtsEI5vyRQrIufX+HeUkjw26h
6e4EainPsgi2+qE/dEe0M485UQJPdMolOXUfNvYLGGqE2l3k+/W+Gptg9jo5F1N3/M7bkL4LlVJr
tjZrSPnBGKsKoHf0xcNqCCijj9c+BKS/QhqTNyuXp5PrmyvlltxU44gpRVjMR/BOuwTM9kXwmWkP
ruwUgfryL+SJnQZieKzjeakOAE8sjsfirXotjrgYD1OkcBdGIANFzhXKMbbYxUgjP92Is6Lte0YM
RKLL4MVwLeCtC4iPc5dRgLc77N3zhRxL9FnSzG7UWGmTuSaQtgwXrfHqy6DmbcQu2+vmnydJ1Nh9
CL6GWuSb/uHvw/csG6b1528SYq+3Z25UnPy1LE3KAiBHtKi+7sUZvzxM/ek3TCHkFLJlcgggjKIG
5zaTy2rVFbjiN3JCfMuAi9wVwA4aejBqvdiEudnwiudO7HhTVs9qVX3DR/jYcNcXT/1b0yyBmSoZ
pmOnBN2n4WxHOsU4jy+scpoPP6oRrRjYftijxyj6pXZ6mr81jmjJRuEJvA9UuP/EbDW40bFPq7Cj
FohWeGRyC5rToJa8DsktOgXHLAHJkES4Qvc4nFf2bZC4Ehyf7tyJYszNNnnUVW22ZV0Y4aaQ9qlK
1QZO9ZozhHYvk61Lbv9RX+yumPh+T9+ZD3YJUKMwlOD/CTJpDETWa1i3FPgowJBDSHwhIAv1TFRZ
eZE1cIjFPkAa/KgAe10PsG65N0nD9bSMfG9+jD7dMOC8bPP7STufAfahwC3gdAPkVQb9SztoZawY
msnJP1mH+dEjzf95xFIcRrSaTHDW4/YqAwkTB2Y98y0NWLoA81OPvMt/tr3qne04CDd/PmReOJLa
V5h32A9vPYCZPAmhpulzwiA4aE88G1KB4DIWJTqUjob2J4YQ4ZSPZp+VipRNh0Ug95eicjXhO4zf
c4pcGBzz7sxbltJCCk7EI3yy3EcxD6cPBlVeMUU2fEYswp7AAu0ezGAVymkX2wmC/tPqjIVD/sDr
Ax0Ry+sJxWLMfQaclz89qtj63ELxYNzlaPwt0VWjKj0OItAoClB7MsAAIQlVXMBHE7lnboV6ttFi
McTmcyOjTW2babB4qDrYfZ4RcwT9V7/oeVpX7n3Ru3DW4vWu+kcD97WeXU2+KrolYv5jZWemJ5y1
2+oz07rB7ZMShlZqyjM1KZpXPxMqGRrpZjnUqblxmDsCdiEOOWCFxCB4xqq/ZzrAYt7LjA9OJhV8
6inhtYv51xNcWcUhqKYw++pGoqAkNxrKhoxkI0PAx0NLpDYEE75oZseaieOBsU7j2aGnn6CuKh5J
nqadeyiDK+3gcUCajsEzsCf40FMolJZtB4Ya0+rUzu4Vn3RSxlL1BS+ESkfHjxQVBKL2cp6t/dul
1YD51ke7KqeFCsQ1NodAzf5kMQUklAFMmB6rT0jxUlEO7fwBsiqhY8rHFJ+8uXkinhCTvrHJfy8U
y8XZM0tdMnZuxpSMxWpKWWUQwPCmEl82KwNiyTvFPZsRnrp8IdOY6Qk/zzkHmZAEGGXtoEe1RPbz
T50VE5JOUUau5qpvAjbwexgbaRdG7YWjZDmegvw6V1ZKkJnSSCZsQyszN+Zp/9klBG306kgVlZYb
v3//Q544dc8Q0hhWSx+xSGo6txllXIIvG+7l9gX5dfkgT7y1ud9kIEOQQAjVxFzFYxSuPqna3IBO
98VuEQdpLN3BpeUbx1fRMmLLonLf0lS+LaeZDCrRB3mxaY4P2t18p3wBWnfuf+ql3evt3LDaGQBf
Ob32BMrdZbozzGHBcvda33nLzoB3IXyuECesfFMuruP1Y5TbygfXsqQVuHdU7NV1tKE6Df095Guf
ik/gBysS+8OFKD+tvuFfFdliAZDn/BGsBFMTpyp/P62NyBYdjQa7TFMl4rhA+iKZ8clXpPgS75gL
vlUJc96pT1vx3i2tlW6QvcfN5FolJV3kT/O8E45ndpKqb/eI8/NbIcWdErVVrNNDB73Z5NFLn0IC
BEwgcFhxqgItb9/jln3uYE4M/SMjJ7GiNUmrcSdO6S8xlaH26ksuulvYn2ueP4H/Bs9tiTyjc/jy
nKWLwaCjC9YuUJDojTknxuPGegE6WgJ1eKWZVvZ8dK61JYjRuhSGMQB8TZsDH7GJdzTLvHt9qCIt
W41Swvi2dFRZ6MkXe1WrUvdCgH9B9rBHv0Q1VOFPETZKRdDj9GiUFG7Se0zTSeRpyo9pDyertKZo
7/e2/pMN/O1wbIYd0LX7gQ2E1wGPsyqM5Vj/CRn76FSU2/3SKSBoSdGl0EbSeCNFCZUjYhb47cMz
AAwpjfxKkuNevvN0nddfZzttg1oz28eylmFWiE7nN6EQz2s1glIgQeRElG4l3hYIVDOqXmMBiHe5
7XqmrfXZ9zCkjs2BJZN7YJwWrp9S+ES+a2+6PKUGfQN2sqaFRAcI9tf2W28qXuxftXuC0QAilMmm
SHtPviz5opMtpmmE/HbV+J4PlaBz8m0oEdCA+UaDRmvsD34ty440aF/EFCiWGbSUdWbUzWohpsX0
F/tbTAN8leFUR6nOkBJLqwdvK+xvOkFUbkslto2gBJAAtF9AwsV68gLzpG5UkBWwnhS95z4RogVc
5XI13fyHpYX1zB/AWTgGWhHngMPOPHhAUJ281OIlj779I1MFfGdZTK/3UssFEHOh53Tbp36i7ZxX
ZC60vA+TznGUkgYsFEH9BdSsnJz6Ec5WrvPnQd0aqIB8RDGBrfK21pmZC6mU+x3IJ8EYjoK8UfV6
hP38kR7el0pSBDOQ3eo3/HfEt3I8JFqX4kSbmSUmw/jHfXfi/3kbQU5UL3aucEgcFSAOcipZBFIp
4uaRkl/zYZ7cYJh68+MwbMWqBRL6LC/1UppbiY07DYlqd8ScayEVeH4ZHaxgYP7J2zr71JnMLMdp
LLWy5JN4FEnCKQ6OYFNtBsb643/Uq3ZhER/uq2IcNDwDwoJCAyudtS9a71HsxrGqqiCiEoFclrd/
ZG7rg6LtFnqsKwUMy2XKpILayTRKgVmBpz70gleRWf3sjU8SWaKf+Q3/qEzc/PsjqQLWbJaIsNpM
JFlwzK3Frtjisq8VLV3qOHGdhsbZhWXIplvrUnN6lCd1rKBMT4Pbgl18R4rB4BOOyh4nA57dsBJb
DwmwJtsHrk6X7YgN4IzoPL1OTV0J8OCLITkVpwuvpdlajddtGq8xZn/07AdhrgheSD6WLxEfd9L0
7ZDEM4x4HlqvM44JXQPa//Y2QhO9G0+IV7v0GzvwveHmzyvdFghxiuoZIQpBzklFm6t9yy5ce3lL
6IZE6baon4pkZ1aOKueWWoLV/P+4kELcGcYJcy1lt/3Lb34AQhISbRw8xd2Ls/Bokx7M5hc8dAdD
2WXDVmnSA2jX7t1RaoWIfksP3cy9mxm1XyFiZNnnQsp3GLqj5jtlVK0rU7AVfXfdGrw/ACn/ZUz2
WEE+W7otCs9/rgdOcW+BVcfa/bTC3uI/GYwDofZUraVCAqhDHhMnqdCQhiQjkdzc2v2rUpH++NA1
+MhfVjMKaZkPTedFOqjeLtN4kORXntL+kstrX0HJNiqvNYxZNgg0wd33plP9RH8Gwv2IUkTpdZBn
S9INpE6kPPi6+45SLLdWGFuGtzjC3v0RjomqtvGU8arhoa+Qrq7WPGxVvr+czaL12H15setD0noj
3ZG0K/su3EZjwS1OhKcnjkXZXgcGka6mb7I6KrfTwTr8SCOcL4zDqX1SsOlT60A+BoPjH5wvy43r
PPS3hZJB4LyL/p0xli/+Ex+rYxlJI+HsBc0w+yGGi/HK6JOUeugPHUGZb5Q2he2XLfOAaoVUlg17
PCe80enRsiM9O/ZCBnKXnXIXhG6hf0Oodmt5AVDfc8yYClmM3MfrakQWQ+y0eImiKrHIOxVnLCsD
/dj9kbEvJDGKnmBDoWrWWIUKGwwQwt1dA6Y0ylTIwpjfshjTlKh/V6Rwokdpm0gP/ezw3FUnKgth
G1CzgnyDoKPxs4/letdXCvn91b+JqoiqkdfvjBs0nqe+19jV4eqVEXvuzHjhBUolSuhgCqIc8/R9
9qViKXbWK/wPnYFEKCqs+d2q4MO8cO8rIVE0zoWsSmlCStvvrOXgNX6I/PX03lY+kDznrjUbZfF0
7RIBpatBbtk0B/yGBLEBdYmFWczrRoCYWHsqrIQfIeu5ruAl9W8nBJLNyGTNWlQrLFlMrfRgUHLo
WOoz40TJkU2BDdNcixCcEHbUH+DgpJEh4gx46wHNDSCg/4nES7iQv2Tz/3CvJZR2Hn4xmP1QI2Jb
AvxueR072kCf5UyIeUN2VEf45Q8aNHcfeeSGspAdrmC6LZPZAQ4TWETnQf/x1mqwrY9pfhvvtPAZ
y/me04tW67CymWVFFqSI7f568pcCAiiHgjGUtDgnpKD8oS1ezS4Pk6exN7F2In6E963dP63HG7La
TXWXygy3v4OBdP4YqTOJvjQhGo0/1KYK4saxQU8MrAFwmBPocwzzEnPBebLAeunFGI8Vo6z6wzTK
dOG0mFtgU5PT0xFzCkNkIHoI+6A/aativqNgkf0h3CXu3ezDn7iMc05Igq5hfuco9hqoO4fRlXpv
BR76R+Dm5rRiQuG8HlWBTRxsC3CNKzUvZrHnXheanFbGYPJrFgo19Gv2LU7LUag6t+/ybHgnvb2+
utaLzXLpTWE1W6lv1a2lFk1wX6QWhvELme4RV+uIJTfRTOyP8cSujIi1B8ACgVSpyjMhFWbIa6Ko
rkj3+xD2Sw5KkGeENVb9o8nqjGDCVu5q60DF4/Z0TidOS1AR2zenNbDrXC0eIr8LRdCAvGdVCKxX
gLCznzOoI0pkwWQScym+9cYibncZ6VRnAxUA52P1cGvpGYXQgKhJOKc4IuQyoVABWIKnIlgSnqzE
4XTb3jdrc8d6azrtO5jvEGA55KoB4BQ8ZF9aliymV1Y5kWFNNdr1bdmsoPTWhrUt8zg3VpS3d5If
VdBy3vbSQ6yGtDote9gslgr18lHl81L2fdU43eO1VYYtfsT6im6uHQ0zsNo245e8c+K72yXD9Hp6
4HKvtwSN61Y47f1eloLMwP1TJP1Ax8iOp215ZZ/D5nciw9byJnho1kFHYOVZgHKX83Ai/oue/suK
W4S86vu2MZGcMx3mOSpRdSDjq/4h/gIc3b2kScC7RuAtnV+wrhrPjMQnFS83y3nSfVGaALfBEO1J
D2fSUaEXJ4tFODWyk9135ITSCcHFSo2FCOcViOaZXK9LM7UOaCHsNdMzDWJd/FeGKc7qGluP+93H
jgHTjL33lKC9DWSbm7FIR+8P7FQt4Z1qi6T5YgHtovJlJOP7XkBxa+KETtW5rA9ir0ljjintbYnM
pQnuCDpW93Q6KYCSBzkMaEXR9msvhuHVNYxPxOXtelzzvVNuEHbmGkz2F8XYcPSDwO6Dhm3iHnEF
MpSqkvfnXLu0l+iLXjLdiuTMGjAZvcjz8LBaOIBU7ILLCXjc9WykOYllcvhMzKuY5NC7a/3PpAy0
y2Etk2HLAFibsNVPUTjqC3MEWgeAxnmzxCgyUX+DSsnzlTZOeJ3/5qYXRZLWjdbFsBJiaZQOEhME
wwmjJUf7nUqp8e3UOlNqsP3ucJNUS+O/bafmpuibfihNMiDdJROl+vRzcKwQGsTCz25KaPDRsCHI
vV7cdwlKp5Yxg9fwXqhPWW+cMlxMUiZHps3nIeY0a/jS5F2eWQh1ncDtQqB8y/X3xDtBcmG7N3yk
Cn3vSAUux1Gllpgce4uBHQiFX70RkJRtf6Xj/zKxiQulbTDpymo/oWiZLwnEmaJYCDtlx/D4ObN5
wcB7HnaCG/4BTLB2RvV6MplEvLCHU4KpySAXEEubYI/K1m7PQ/XWy1ZD6D8hEzEsYLXSrqROJC5R
ppUt2LFwa6WCl/7FVq18stHoO1z+JNbHw0oD6mk6EaoU6fWw6nElm8IxHlyHaHhxv8bjLq5RmC4E
xb5REBxkNe/sXjb+gJOSuUQHTCesIcOlOGicJSqwTyrjn0edw4Wou2TvVdPpSnzqrwBuWkNV5KVx
fHVuGcxjkRZOynBJJewnyRrg7K2Vx14metPfAIKIhZttVqWHrheEskKn+68E/Jq6phuxHXqE2P3+
5Y30oBGs2mZzAp19JCgDxJvL1udHrOSGkXyB++d27qaqlLxIkCsiAFpMzuKj9bVa7JdRIKpkwyhP
4sJQwWFr46hTE7vqKXRZG01ygtaWRuEyI2E8LqwAguxjbxadlzBE+uYpZMSBAa0Nd4ZqvxUD72bh
zUH4mm/4YcEXFEI/SD4vI1Kj4/AkiqMeRlrAw4iCyLT3gLYbMRVaR0JcXAxnw2VJ6//jo9r5uStj
3PObzJS7zCzaMdtGOE4EfYqhYQU4r2hH03M/AS0FiWgqfEn/2dTsvBbVB6aGk6tiTAFP2A4D/R4j
A+VjAiAa4FJa+gQBb/oEOg09sA2lwWAl4IGiAC4ZXoqMOSzQbQ2vSQlUpMe6fH1GQExP7cbgzXdk
9gE0zX7nePdj3zPuScZRQtDKF1Hy28a2d34bOLdYYA3UFv5GhmUQQ//UNiT19GlqNV9w+oTbg4W5
pZrbo4AAqRui5rjKGmTg9uX+Z/cJfTloHx7I8Q4h6qqFa4fCfXWeUCSNf8rrYJzxc+MLhy8HFhVe
pYJ1520GKOXAC0Vnbkfz50Qh/YLTk72C7xPTegFjMsYYCqiDHH3MB7H6TeoryRUtGVhAJmjoNk/7
8/lAmpEkO3d9qibyjl8Jrkaek+cRhS15PGLXyOjCyMTCBfaS4zo5PjuL1xaGS+wZ6lxasPmNrsER
kGj7FbD/Hnb3UYMj/d56jCtIhYP6qy3yNvMp5oi2bitU8f01Fi/I0BT0vxjrM5SAI6NTgZiQ26xc
QQX/y6Lyxf4t84hdAfGsNqZcydFRYIikfetvi8vuZ3pngI4IMylDVBqNJ4uUHDEhm1v+2oZZ/lGm
qDi86axu4RcceaPIO6X8yRiFtSpR+UqcFTwGtVW0sjqeNOfsUKJ3yIMHtbLSs4Xh3ySL5mltqBiy
z+Q9ids7DVE3oo7avv/SG5Csms8WBxxaKE5VToFWmgUcQb4c4z1USselywNjkjeYFmJnOIlX0S8n
iRwZiPItEEI2DaGBawDFpCnvP9grTiwWB4c01oH9gI9HthEEa48GiB/2D2hiNocwfbJttaXpHgiv
asEpEYJZRoQkP1Fm3W12gMXQd37eTvf5d76e7pmMbBs3Jzw+KbfLZZI5huImi3dbBzGmGbKEWcrC
NUBLMdcXoNcls+c1M/M1COf2rfQ19uuw0kiv105fm/iUc7OsqoNMJvULEY3AH09F3j2O7+Qe0Zp/
oG1xEkZzOEdtkMYUQI6dLpqvdegSdBsMgv8EuRE0vCaK97AJ+R9aP2FUNhQG0imToteRqAbbvMUx
UDkz7s7wKD7q1/AhQfx504e+u60y8lb/EewLbWV4PulQM3oguVwGo3hIL8uRuZgVMFZlnepVt61i
PsXF+YEXDVGvGZJMAABIlZGYTreCmqD2JDeyAwOIZHALtbA74QetryM+7nPjq9zAUQKEAJqyOKL2
SocOy4ELWcCXAppHs3MBCwT4GjuP0yyF+Zyt4yQKvGBKZ9HeDrfuQVRbKGgC+lfcbMKu2WtbAMtY
LR/GAb53HLnShSAc3K+sIiX53qPW4gYUf0d4wwS+bx6Ilwuf+cIVMc2TnPUeLA21dWv2vRhJmKQk
arBUpnYzqHG4nxC3N5hs/crJawdHsycOZF2oPoYuFz6Jxv2skTr6/lz++XjWj7u4MOu9cgEVvOd4
5qdRCJurm9RyfDR03JDc46dts351+b3MmNt1+TIrA9Pk3RBerYjD24yb8+otOJV6bel4r4zSkTVZ
Ix/Xab8CwEFmpk/8M6z9YJQmOrQfbGBNhlAUixAyd02gY5u3OIAiJBdtK50XE1WM05JVv1BI0vBi
ykgHZYUECnlwmStySfzFcAicetWvtB/BEW3Y4/QP6+I11/qCaslfS1540zauOR46LmfbeiyOa9Nx
iZC4mnVJZ8RS/1ItXfrEnKfbO6JviZn98NBfj7gCDrezc9rC0wlx2lOF5l8jE/Xq2miIzJJfXu5U
OqwSXCaJiPzfIE3FxdpODK7IAFGyfdWwjMZMSEmJZTpKUJA90ClLvz6RjIrVtwKTr2+4ZymAc1KC
C9aVFvm18HVfjkKhpzB2ipexc6AejXmpF7ORzEtIoR3F1An4G5rQdpXepT0TeWZRZuiFweOIzM4t
NFk3hzBlra0hB0E+0BSaLMH96rBpSxIYfQ+TRPrw3un8eRN5ylfZExwgJeffFKmHKnKJl7fbYUcj
wWODRA9gikTuyQcwiXUR9VCJM76FnPX7tBHHL8jpTMq2/Hcs0WIpz02G9DgMK0k3RtlD4yIFVdwl
lDpNJBkEPOQCsFdXvqmDiteSuV/0Poi1UPu1bMUfHGmMJmrVhdZY3xlnJvfJmyvnQala0xsxvVqB
fA8qq9nmMzzKdPyGMZPe6MAysvEQQzZAucrnJ7h8hJB/V5J41te6jEzJvJ6sbBW63MohpzAaZGwB
JFlZ80QPZCzPIWidjytU9xBg11wICfLJnpRjgZnXx4tUh6pJkkFSM+p6V430RHwe/2cJ9ysD1xNR
cbKUSD0SkNINc/XZM/B2Aal/1nd9psqaWEMKH7wsk1FGUDMk/iYnmVFLMUga2nNjKaZHFvt8OBwI
OPlz6p44ZSH6bkKNfoidunMRH/0s0CukPeRE+9mvOkTqIj4GYdhpBRSat1LH7thUnY0HERd6VoDk
plbqfVx1a+XLzyuYDdgbnQXvsmTMe0n8rgEBD6ts2UXXeKpuohCYKSLhyxPYP+t8uBPHEjybSwov
t837cgoaMfDXK8ObaVWiqO98XDPc5N3yY+ujGWXkLg7dwx0UkdKjCvilHvocdvqP0NgWgv22KJwh
0E+5coDrklQySZhc0zAB7xNwwplxCJDVYLS0M/oaeXzk7cF4w2I/WGABqyIYnr1y1V8Yu38TgaEN
lW9vdWV18u0YqFPsHyvnLFs9ee1V1+S54HOnbWXttwIsI8tbwfNhila8DN/zischb4R3LNip8WJV
JzFSQ+1LZnHbsJ7Rf944oZJ/7+S5Fn3yCS56rpzvsXyYS1eOAW2Zt4KvhOo+dlGdN0VRN/bOEVqx
/jAtEOyyL26FvoQaY3EHM6n8dqydfrtIdvhFGgLRekofV8hKmpPOQzb1dbFvRQUDmLRwwiGHdQQQ
7LSkFHymUdA+mnvSEN0zGCrR/P+wqVikp5jnGI1iSKhoDHwQtyG6qaA+p81Mx4Ay8Folb4PQW7va
yLZ+WrAsZWTM5p/QNMLs2aylBWRt+zTOTuxwaEvujGwWcocpD4NppkqxgWe0bLNNQGvN8L2JYV9j
+N/FA0K6S0lqKoIMQlwx30BXiN0PSfp+ybhCd/YxmjyC9eoHx1Gf6z5YelQvHoCgjXLgU5uLRY/b
t5p+hh0z600iyE/4rkjDWajid3aKuT0F9uR0pb5NMzaT4aCdfMCqqmSvVvBfxQZh4C3CxTg1MPVP
+KuTtbCT+FAj2l/UFt1hB03xPlnXA0iMDTaNzQTP6fWE96kANDWTizNpHha8iILaylof5qBzqhk1
fLm0oGERgkMwrL/MFiyoEzTLfOGPHlEhpwp68Jb8ltUFVQbjyZ5QtcK9UKyAnbERqhYbFtnRFbCy
YWfwcE3+DxkgnGAmZ6NmCLu1sLdzKe9+iE3bZzYYK/CuVRDQPmMCMmF5OhIfkLz9G6p3tNzabn/t
STdv9di/Sc/sJnVQJRth0ebAkZnDeicUPyCCnsAztziSXoUo+iw+d4qTXDrW2N1YR9oopiy6s4de
Q+pacSSZck5yMmUl8lz4Vm5b07mQC0SdjnAd+SAyaOy/HKLEy421z5tqVSlpFT84D14JV89hvE7x
+PmW4rgYmPZhXD+PK1uxfVtoRnVYGkwp6vP3VmcGdvURV/BfHXIjpgEnWxc9vUzMYM4hMaZAX3Uz
P2q/D6UwXRv75Smtci+XhPV6coGpphJx8++emzJ35wuOA8qpuSUmnoUmZta6WHKI5XQySOfT7gTY
1bLZxWRFVSt7FfBtWwEM9vWfjTqk5jI/ePxDrrEa4Hc3cvWYVK3wclakmw8KpV+Bghix/ZZEz+st
vCNNpqvmtNGJ5b79oBwVwKCrCGR2Px92si7vIGDn7CzBfW5suTDTPTNUAzw6LMTGN94C24vNEjsl
ORyVQZUettkWYuiUt2Lnm3O8kYLwrLSLmAaVdefggXxIgoCjkFRNtCVGkzPbaoTc2Wwd92ZacFC6
dwu7dhpGhxt9Y+xXozVkQQa6LRLfQNd0NfPMeci8exLcdOuUWQ/bu0yhBqw+/xmlC+rpEZNml+Io
xd7bYe7LwxDl89X2z53pUe9GlEaNyVT9HGo+ARZg0ePKpBsa6MYP1gDvMD/Dsg51kyPma+miJCGK
QkRhBu/Em6va9aJX0vp9iVWPo9WxbPUupYxQDLnrKPf4D/vVXncCCKA3CxmGDlTBytR4Nkg6wxD6
5J/I+iKB2wga+NPHi3PkI6Cj2G563f5sIowcpowvY+utPC8suDPMvM5pthoKxGO5MKfH6SEcV2sC
GHdki7RrTATgTpxIFjqanu0lOYLGznS0JOpH2ZT84AoRPcyd82d3m49FsYEz6keaZjypv9FpCrBT
k+PSsPlRorE+XmXxE8bo4EUSK/IEqxYTtHLI4I59LtWhRSAbaGJ3PogTKVncLEuqCEjgMmUSpb+3
Y0YmWpwc+fOpNeiNLFxHL1WNoIFynHYEfafbJHgLT8LN/6nhdzJ8j+0COOFF7Us9jmC3mk6QubjK
/adI551oJbDPnTeKimhuOkEAvGgtCvYEOlzcnsfLR8qr1/hrT/SizHVXVRtnTglHDl9R2iFefwcP
mZwUfomkP1EAN0IwVN7MBRtHDn4P9vCMRSMKVjLnHnHK8JCJJ5PBETuQ5wAryYAuOVp0C8Ns/AWa
QWFbYwZH24qP6MUWLG0cM061XuQ3ZWSTeZrFqY3RWIm76p4ZMABQvieO5A+uBOkU6k5UtcNUoHb5
Uql4VPM/OPamVJLBIkCHwyGPBF9D3iJ8J/S1udT4jYoEkP9Gll6M5y2sETgRHUxLJeVqCXnQKtg8
xErHu/xQ+dN09DYrhHzpEv4bJLSArbfG6fycFWwotVBUS7SGrTwD8jb8FO//OfwFYB3k5/7igshk
OkvrmjMle2xdLNjHWwtjPr/y/ct3qK/no1eyYeWOEoNYRrNH079HgKpO+5rmGCbUdtzIUGZO/PKa
DI0bAeLi8MavJCt0vM9K2RUyIS/Lkm+nv6P/flCT+bxSOwQ/8U3KZAG3frw1B9kqBbA1vE5/uH6z
pKH6nlDKhIZPq7x3wUP8BNqxi8z63uNurBv1AzD/IPveRgxFyuTXzsmhZ5duMaBMobP+8gHPeIN+
g3hvrkUb0a/cjKiO19WL8k79F8YDINCrf5XA8wmJwOwGXQCWBS50juZ4K+SeQxbB/Ocl9U1mOjjL
X/7l+Vy1HHGufjwBVDFHTKQN2cAN1etbs2F7RkMkFt8Bo81WJbJI90H2rSIED71U88XQ/KgrUQYc
690jxNKGiIqk0S5NYqmaBqdKw3uce9LeZGDUjYJasG/M2hNJkbJO+EuA43FGBq4cnKsBhn1kjHhC
c7ylzNq1DOk4rsmd9V5bjg9Qfe/ZFVFZN/Qe9FuGdeCGq2u4aVP9l1jO+8n55/fPYTh9twjjK0X8
+8eYNsBcPTatGDBSaoagOe6MGpfpoZkZewsH9uyii2Dvs3lCEm88zfYtkV0ZiXqNO7/rgruRpt4l
5mb60LWZepO7FL95Cn2HWWSLoaQLYgTpgUji6Ry8JVgEKi1WBxHz8+jhRDFGe4uA9oZ8Q3X+PVEf
IR3NksGoI4qZnQIn6KZIRtTyohScPggZ0o12OeB/mkns5hFQOfGtZMwQSR8RtPgi5k/mzKJ+d9ud
gSELX3BdyK4HugC10WHieYCw+N/YdokrXprMbeqIVGwxBOM7WAnIKKMsZy67IlQ1uXuP6I/gOZbu
2tboWXTn2LiwIKgr8Z/4UVM2rjQ559Xo2LmTHGDKkSzmZ1Tzj4ymV6t3JO7XXZVYDUcl5bO37C0G
OSe56ehf5kIUP/uj7FaiqjxL5AOh2UpCiMjfJS5KljJk/BXtHiqi0IDrYHQl3ArnDtQqbw9zJ12H
Ks7+eMwlUKTEpvs5hJIOzijJPku4vCJEinHxrp/S0+bm97Z8sOgp3vYM9ixkmLvAZLvQPOer+0Rl
8yTrtY5BKAbdlmJQvkv0BS3fNgdsuP/Dso49AvFYgIIEJglNXXc6aVTja4OlHWqBNGYsDOLFeuou
HA+JC2o3BNgyxohsWdLaAykti6IiQkGv66vUeboMAJnxQPZK1axmYRe6f777rBMP8swaFEa63VQ4
MNBbdnBhFfL4wO1AlqCMWT0wAZEDQGYRdGW/osMpC79+QLNPXo9uyf8wBM5iOrydt0M1SiBhy+5g
3apQIPATznKRkwduDcEgD7TrxwV7CeEl61phK45MrsjkfSK+GLwumzPxNISOzklCpvXozaeRdRdv
ULiFQYMOZA3Tz+JaCeLXfI2WBml+kHyvjW4fefWDPZOmuAsZ6IftkJiztiCPshg20PcBvHhv7J8h
liDMA9UIIvG4TpMpPtGLT5N6ITMg+7mJmqyK6t+rY+YHq8uGJpfVwsHca5VtO0rmf/wo7UL//KZs
fAeu9/XQMCVJn5CvXv+r6xrlLZDBNQcTL+tghhRK1g/pq6VSIx9hzxi4TD+Ly7E9J2QDumZoev65
3PKsEvHYFWu4ckIrjpM4jXz4IIKROh6YBJaoJ/gtYRPCVTY42CZdGnEHA0VM5LTYRldOryLhzc6F
Spuw2cQxR8tetNmVc+LVqM5VLQmkOAS9YVTX/npc1/XSjAU2U2Fa2N33nHKV70Pg64l3tCnCpVQO
IHwDPKpf5hfnrHdcvKyZ6leg4QXPfGl0VaDfx7JGfilT6rsFKIOkPdpGg9NxtXra3008zzU5qSP+
Rzj+J+tq4jjkNvTG3/BPRETY/XztFBXcL3kOj9wnW8mWkdofenmelldrGBmMWNOQMTpSGGOvb7jJ
p6kkgy8AE852X0eq8jaIYSTwq6vK0clp+OWrrLS82xIwXc7j5t9+rraR3Gh9hkoBxySP8XT/HEek
cNVfGx72Aa3W6ssd3JrlSC1w8w38jOyLxdlzjRgagHVWmFC6etJ3vILEhQEvQ6OerZAQDo/8G81+
n5y9VGMUjIBvOyn1xpAvOcJOSH9gs1hverxTsPQbENmh6lTvIXJRI3QCiWqTU1wdVomHMpOYM7Gb
rhB2VnUs9g0qRb+e5iVR9RJLVwTX8jYelu1TTfvWYXZGvxiylUFaYAzzAakc3APwEvB8iPUfaHBT
Fbh2RZbeLDXR64iUqComFb7562LFH8DamPf2gEREHD86Y/vYM59L3i5mCeav8/56y6pjpZ91dgAB
B3/L2k53HU5IuH3j8hE+hnQsv+JUzoxB4umjEskyb/BoSFpyw82rLQaoVKj45srMuf63J6C6FoNu
fX7tQ8Abs05jvtqypJIBGFq3+51SAp3crzu0//ksO8exniafC41EunTBLKYlCPLEIsMsC3Liq2pk
RHvQ6iIcxg4hj3JnyEcnMphoJcn+DZtC1Go5yvKEb6Y/nHsuJSvpkrKHW3jw6uKrZDmFe4pDf+2I
N2esYNHRQzMHzVGyrnagjBd0cS4nXsjjdPG7NojHv81K9efoCm6gtL5ata2kiHR1wLOp5F24ahbW
NYdnC0+SVaNgj6C7M3/k3aOxc4emDsUwveSGCdYV9VLRZ6J+dRa+CQBOfMJ9x4xniR7g6FI5FNIJ
4pIDlgEkUr/hXalG4T7cTqYPE/CWo0IWXSc9f+JlBaFGey4/mrL4fKdpFWsIWYn3u3cpAcdKFZoO
usqN3hdVywcGNBzRcctvEwzqnX9m7UvcIy2nSCgt7LE/weftagPhreZLqRjsZt5ukht5J36lHjWc
wuQ/cqnGhzJwWNM22TXzScPRFa9JKP4NzOWr24pRsqio+SsuMuim8D4jgs4zjZ2XzbSszomEXiPl
AWRbUomtS6Kprjlv/jhrU1sKWmPOw0hlsPEEgA5khc4zAQtgMHxo4JI2yc4lXaNXNGSEtAv5M0De
Cr4r3rk1fbWEH7tXEat7a5jKnixvMO9fzXtojGSjdAYpH+7Yzq//PA6dH7bcY0FKNaaSllk4m7YO
sSji0dgF4vcAfEUPVMlfz3qxJNAxQD81j10n+g9TgvUcHsB99XM563JOQx4e6xHJ3w1/nHRNhwVx
8gD4n3HYF8unEY9Y+rqO9kzigggPV2pme/d1bUH7zSQtnPQ9Tu4tN6aAFua5DvpuMZ6eQ9LyA+NR
amnuPjVy8uoqpbZ3mYGce13dIXHKcFeDjPgQWx3vTrn3b4N/WBo4od8WYRMlgiGzKSCCTROmcQ6I
/HS1JLKXf3bjlIMtfSR4oQQCDFrpMOus7v1FKySbME/tx3r2qmb4M6EFpG5/uHwJy8oNW3rsHGHQ
+IVv9ANm1Q2er+JaeqWMUTxapbXtpTKWHmOgr000fOaDAy9LCGqb2N5SFT29CWUmFj7Q8lf/kk3K
CbfmC/dZemKgziDYLNzOo6Ufg/dZBpggT8kbHsl9KYJSneHEBAvgCtFugbNyHp033TQuX11MCS+4
GfAuEWbTt+nvcFCOkNuXs+GfahbRZnOQwF5u2BmuixoDk4rYkxZcnJi7sCHVCXzIGeboykyeTk0J
GSF8ZzcSutAMWxm3K9swiiGwB2cchlD3Q7KA07rHXScZfMPgfjp0kqfJqarHIQhUKqisHsjYQEqC
qlnSGb2P43aHMIUQGGAJ2LL/H3CIRBldVz+16XN4jZubVytsWan3Ds8Dhi5TsK8pqNJoaBOX+NfE
7hgaI7IrnB8XDHIQ+xXOXRAPLai8HNBbsH1xRNBFkEBUZWVb+KyAXsyC6Tzy3jZV05HYN/OhbLPx
tSJqfCTyRiWtE44rBWTPtu13fRZGLoTa5ktOn6XE9AS8nWEI5P6p6hvcvYpB0WbgWNITJUY46I8a
yCIPTMb4LPxKwmGkVH9G9voGDzOcBrqHE3UHf1drrUKoZepqXwtiWwlF2bhb/C5T013xQDL5pHls
Pb3HNOzjoj7V+Aa2gnqz5zEfb/H0AnM+LGsOTQuYsV/IjMbVPfsO+4gwxkm/Kz5qAs2hVFqCU3uj
hTQpHg7sCxoS87OLFWLOJ0IwhDz5Yx6WxHGUEp6vhZsQIwm/aMja1vWcO4rrcFbuKuq09OCDWJGo
kqCFM++eUxnGmLHH4fJHIKcwA3cjbcGVyNx8NcUbnymcjNZmOY5ovGwegmDQuRFieNfy+w6TNZYU
pRltRIbtyHJay8yuAU1rX/UJElj7aQvUMq+1xs8j6QWT58AeMA48y+Bf09Iys6PtNNlCWpsL5V6p
5BB1kv59/HeBKSgKCukQp6urpzO3/ysDCpQEaW0fmlQVbGU1bQXeig6fYS1C8I3Txv9I4Ju7kZ0o
Eemy23i4hohnKGhlXA+M0cqFVyOzO+ljZk0/7ndAjkVtSUd9+5b8Ly0nE9AFKWbtDzm3nBvYzJ/T
exSVE1Dsi0bBpTNklTDO9FlLf0ljuiQrL0O7aKdJXhs3CIrxEU5cGvjxVFmLRD9ZDiKMe8BMcoF/
/hdt6gKJ6IvwPIOZa6KdXqlWVhJLJDH685VWMO5865IwM8o18WyJqcAzbWSlTHzkuTo4et4xL5rf
0F8cCSJLBbd5iqCCKLUC0OtIaDAjRpo2V/f+nu1coQwhPy3pVISpPN7pfuxjzDjLHaVv4npFRg70
JIVpZKk2fRx2cpg+c5HLY+zNc6APVXZGv/Lnz7xkoHSQXNnj/cO5APgaqXHo3dzsvF+Y6f2AbhCE
E24vE/T97ktj9/30soqtpg/66IoE5N8VpFF6MMvSIBw7tiWVCHoBfKZ6CThUKkaJMEHrj+td938p
qjvjLajjNYPBt/fLQr53MLkXAvrioXxwu4OztcGmJamqkTq72TUAEIYHDH/ClfL003uuQU09EGFS
Kgfy+q9n538pp+6G6ILH/nv2rRK1R69YyyfGo2GHQV7GxvbuM/hBIujzKSBbuDqRfHSvKngjjY0e
2xeTOfDvtBvNx6x/T8Q3Hl6wV8s9rut46SSQdQLycIXjkDFsAhvZo9ZrojRv+o1uYp5aIP1+suNR
fFOFeg9Lab3wedrUYTRAZhBVyARnMrm5MXqp5Sdq4KFAifNU3oi3ZSeQphSUECYbpSsm9N5t5WDF
FRM6r4dQLDJ6SjVq19/5dBFYPI11NQlZQ9Vo9TcsHJQHISJILrMkcgExfoa/fs696TPPKFwkO/VM
+Y387GZsyG1QXrD/VpR0JWx3mmLTuKhCDpxxli3uLJiw/vrvKZbGLgi6ZbT1LoV+Rc05MRvB6orm
czd5AVPRYlwsKoGFK545rpj1eZQMTkjFnIxsOrisUpHqQ4L5GwTqO/a12Ar1EbBHhv8Qy5wx9O17
d4qxoiUAWZ2xP+YDWtyjjwTZNXqY0Do7J+78Dz4K/9ltCbl4MjPwiwV3RVQoPYXsIrkyrS2v6z2B
Yl04S3U9XVQcJbwR7Dtt/AJI23byQof7cWjwnH3GLFeqBUnUQSV0MP3UaVRpncCT4dxgBXtOHKT5
l3VMVrKcn7lQQx3OPwwrHVdHw1TNkDaSdtyOjosBQQ5ogWlGAqC5kgD/r7CpT4b++/bCqFLth0ev
64/JY1rVbfsSjyJIx74Rp1j7TcVIQezWCNFp7Pv6afB9jT2iivFLNoXNNQkYQCFCG7eQWzx+vETW
TP2ywA6zSzYdimaazZFTGdiPs+HFvSS0j8jeUlK39AdM0heAGLY5yogh7BpZP6DDh4c94wQ9SIEC
2J73JkUcL0H3MAZrpa+o/9Jj0LQogYAr36/YOjoJNu/T7Nb6/M70ePa5fwKltCVuv9YZTDxMHbfS
/XOhXodGkiSj4Ko72iiX4R6LBdtx/M8IR+TXCnjOk/cAcZgu89h+PYtduIYMFZoC+N+lIhV5KvJ2
W9////6NetEV8/ZUYUm+p2sDTVCmTd6azUJNY9dZ7WBP9KVlQDG18wOqCosb2+fFZQghy3OSJaDg
AGAF3azHaBngoscKpMgVorTPEAENXx7mrLBrP4D+TbANh+IBQfeej1EaWXEjg8jKegEnpJBpC+Rp
IwZ/vwimEbbsMR1HITL3wForpRvR7/lmDywXoYuTGq3VZGVOVTPZIl8+dHw08xfJUbffAfYB9epO
RfYm/A8g3C/9KzwDMHsQJga2nqzyU83z+b6rhlc2QpCjTvqBBH5VjtEFkx7SM8e2CTRZCd+US03D
fcvW2/mXN+lFt4bH7BMVEZzH8enp4HGSVNmT8vghBVgyyuWZubOrTBly0+7JAHLanrsnwz5xc1Jo
VpOn3cnbqA7SrDJFunS4Yi7Jl1kxceS4ayEagNQgfq4YziZs3+zlQ2GZ6jed6GbnF3XO37GNBK/k
Bsa27aq/nEai/LcegBwv3XLvFz8W48tQ56YRpo7cy2dodtZShZLFl0rSa7x9EK50ZTwY8My83vnL
ub2YSGANbyfq8EDIzJM4jgcBoXXIfh7IUzYnIYJ4GuVqpgbE9DYAPbTrBZ9ps2fi23t1yF5WLlsz
xK/fjy1OprJ3kQhoxvCqgY6EzMlfY7WA9IRDwxnQ9B5D0UuLiiK4aRJTgeuQo7THK3KaxsdLmBAB
ZxdQh/WT0v51T0a+NYiCXp4u5eoZGQ4Wv90HO0dUr/+QCKgiLICLjGdc8ShiC4gUCv+s0Zx8KyAA
NLtQfuKrF/ww7PqJ0eV4oFF/qyiTNAT6PU4SKgkazB2M2amqB2LALLT7iXz4RSkdHV/v5m84MbTl
q58WUmffdRisu0gbgl8BCohEf3JhwGxIy9F9OHF7wn/3caH3GBdsCZRnTnpYYKBTO9BxSbhVfL4t
O2mNCCEVwb8Sn2pqltnZ5+4GCLk948aBSaHgzpFtMlYoFMwWXUtYHgmjCE1yCYS0iVhtcrGXyY/o
JmqbdVPx7p3SnWAjQJvukzUF0YWWhh6msxxZ1XPOZyLRHQh6hEPS/ng4ALgZcTyzaL79z8hge1Xe
u7gmgv8mzfbx96aG5cDp9sag++e1gf+U2LGYN5a09fZEyvUVm5vnxqkr6XV9/YgqIHqHcqHmtowv
s2mfEi0x9m9atlGvwjZaClXq3oKAPkeWId4yfObPHCqeDZ4WY6OBlfyMjQRGpy6OwyWksJn4PiJR
5qQjFUSCBB5p38CsnfDr8vgRLwj6mHc4/Yf+Ww5nnfW2ZO0Kn9GF+TXgy/l08c7BOX8RB9ieJ7KL
eSQDyBJyMKvwPnknDVHNMEUdiQsIk/mF4uKLOSB4ZWqnHQI9q7KO2pkuRIpI3yJuejFPuCfOzqGG
zXChqPWXKHucYG1GRgPr+FJivElKYkE7q8fNVeheTv0SdB4H2eplXWImhFTJoH66q+lX3/5hPjxG
089WsGaQerzWUq7zXEvqoKkYI0Q6Hi6aM9Y/y8BAyQn7N09Eb6EaPswBdUlE2UNcip7XoknWj2oa
EuEMct/N/69bW9iI9CZw2JN9SUqxXspWrvAthnEFq7ce4U+LRpk0/3vd9683HTeT8LqBlnme3H5q
qUGmMYtAMim0AqOj5HS9YnvZjftVuy+XqyW7lpzhC7ZO7Zw2TxVijWSEu9UePDLmdGP0kAjhrS1b
GwC46QWjIou4ZbUvuwcGEgShLOMb2xUM/jI3SS+/lhRH6uD4xpAdA1qGxJ5tS95R7h09P3vbfEST
8PiHXUP7BjfPottrQyQggxiuyvDLrrq5h0ig3xr99R5YmvgnBJ2NZgiqpEyU0zSDJNjfz9yQqn6Z
aGXodlTPhz60YuelaD9/VydltzgBf6qnozNw3x/qMGk8EfAFOxt7QaEUG4sPQIBFXuYVatns9LVM
VFGlZsOtEW1BFNVopMJi+G0dPLNXlCYLRkM4DLCkc7Ka0U11QSdn0g+Nykk2TY9+7gYIf4sNk6c2
BHUDHn+7e0/E0c8K/2mI/A5tQ6DJaAoZvB1qiqvQI/7bkvz6P7JpwOLKT39X7fg/wfdnSDzj/OXX
oBHBNDKrJ9CJPhSddFwK1WLpkb42H+N7PLiepyO3Se8s+Z22tL2DbkNfH0kgyd8S5xH2juhy44lE
y8RKlVt275lHPgm2QCZHy8XH0lSsN4W0RcnHijEVgkSg0cQP96KmxOsRnAXPC9f7h3B2CyW82eHg
07Mr/W7xsa5OctjdDKs8OXQ6Rnhb9qi6EgwoIDJ8Nju3XtvETSL39W6fPQWbtzVfV+HLle3ZfCb1
uE3jJy3cOuJ+fkzHp9g1OdJynLKjNC173p1r6fIA7wRijzOy1M4j/rsG99/ftmFRllfbAc9DyJ2Q
TNTzSty0czT8vBq+iTuedn9pFBjqTXXcnOrSJJfiHcrXCx/u9XpIcL3YA/NRbSuta7Ckbnlm3H0M
DO5QM8XcNxQy25lhnUYIXPjNA0+hgXMm8aWlRSMGb0HIPhmsB4I0TCuRlF4eHRFzPhodzh9viVoO
uHkU+sTHOyFXqZjT6su6XNKzh+MDMbCpBdQSwXH/JzxRWk6W8EIsxO9i1ssQp6K0frqu1M90htbH
m+N0cZvOtbtGrF8/72pMnLXSgUGdYVnnBb2T4kd0xyDZRwWrt8c/9cHBW5FBy2jmJDYo4UI1aRKl
KmKkQznQYLYKAO7zSuLq4r52dPAsVYULLqNGExJH5jVYMGDDs1ZHzl9ffOvdy95Rvqa4nJfbotQ4
r4qA0kfs0oX+/Uoj8jG3LEb1uumEaEVNDeU/wyNGas/ZfIu4Erqb7O7dJugFjRqtvfcLNRCHeloq
hWCup+2PbRuuyYiTBNVhsjAs1WHi1/k9aj1dCphUz981a1n0wWiSEzFFA+7epGOl7yj/2h4ibYMS
OT5hbPESiQZcSJP5sNEn8QSukqEN+MHzH02ed3r8pgQeIrPaJXLLH42n79d1yxo+bA0ZVsPnxC7g
8t2Fvcp6QyfoptRsSwAWU/EvgjIHvUZq9ullyMuwcF9loLnuYqfMs97PwYkYrRYlx3gpOWHXjZo4
v25h6Nl/jwc0O4lLIOAoaed87gfNkeiiwOqlKGJ1iH85QT7sVTWxUhkfRML1OJrdeYVxuddbrXkM
FkQOtmou92F10xw9EyKiqTpCtOqxPBOXH6IQKfnLaBmldblHHFUwMg/QxKbwItZwAPh2Q/tPfShJ
+JHt0x/FG+Bs/mLvDPRC+4qKBtet9/8EVivqoY8f6KM72RPDNM2GoDTXtEEXjfBqzODiEwOPtpa/
ofrgct3bkVkAF+dU9uCFHXw2iBG9rSMXY4W6xYe1YKhw6lmZ3QzEebWy/WWgFa3XEVoHvLHHD4Sa
vawOW4NZwvDKN/OvUK16UDJkxLhNHb93lXyxWfa461HiZ8mlDtOOWlhQ+q4H2IRYO2IYHxozFqez
BrnFG3OnsqpzWnaLqmdLZuTlSTaBThqOwcklzLj7k0PPa8XsFIQbkHsaAen3fu23bmupwSoKkf2J
LiUBzZjh9rcrQaI0Ob+EirWv3trp1EFRD0jlC6/NyfoQY+Q+WfkYSOaqLYIprGoBV7OiCx+e5woV
9D62inMFrfKJAYqiWvZNfI5UmUrzR4sH4CmlItx98awigA62GNTK03frKqkDGpoPqpizg7OeN8GY
Ylh6HB0qkYfXJ/VapXNd2GEusXbYmCxNG1DrDM3oph7xVmBIJSVmjIY6W9TP3t80gEm1Suq+80lc
la6e0owGVlcZSjz4CurdEzq84orS+qiy8CGiWww8nnfcZ+2oATVmThxuKBswHjSKK4pxt7K+Nil9
y2yhjBoiVjwzQxftZ5zGPjKiMfvp4tk2P/IGMVyXFTEANKFEtYszORLFB1dR1dZGRubD4vwItxnO
1Py1+LnGMS+OoggRzslmZ6UOmmJeNyHx+3/UJjN8dtCJPfCRTQCfWRVq8VuttzYsmSZac+ZgZQMR
SNnQ7Ai+zZYFW+KNJq+GWNRXL78q+2piup8awGPyc5OkevIj0c0b5phYwq6aFHaZ0Myo9HGF9j8c
WL0DbHWubnFjcjk5c5l+iKQODQFqu3I4oMrqR8m8qkhnAaw2Jps6UVPD7rfPM+Pu4z6zBJzEi/TU
Y074mD6yHgn1wYYrPfpLdW/QedszGVJ6Oe/cLVg6VyXIyLgpHZ2d+cYUTlkhHzcpn3Q0i4LsyO5V
C06R1Jtp+sS/wx6f5zTjIjE8fRzc4fpEuiA4ykQjfFSZ7Egv/keGUg6B6bVv14envFKdgP72/qCu
BxYEiA8FsVOrlA5h95khCfMpoCcsCUHhFw3YQ0H8XML5iHA+fYLhaWEdMCfD2j7dB5ProSrUohzw
ENsH+LULrL370Im/Jr4OqxZz9a4Wbi6ZO96AuYER6iKGFCEdcOuvsM7KdFxXUnwQEWF8Cpm8EUt4
qTmKBNnbqJn8lkfjoTD/rIDm11mKCFyBO2nsNxh8rHI05maEWZ64V2XiDJJyrrwUI2KY+oPAqu48
lLGYAloXGqdP0vYs8GTE37+x3MSWNygunTUEnQQMCr/BWCAkNa0jSch7Yh8RIRsQWCdFHglUin9z
RaqfGCQAin8eIO4TDdNG2IiqpUBbQPlYcOZG8EwZfo9eG9rP8lSymXrRle/vMtN2h3xUkxkm7hSO
5iGCTMIe6CPAzgX+lmzgvwH+u8pcOVs9K6Znw9cp4pn10O/hegZDFG14QPDfbAe4j6SWfGbRo/gU
FAo6EyrEK5MXTwV9nfjyhChAx0B4D8OfEkVE9XcFDZbu+TkqGQ45GGhKtzuBYiPGEUcodaFy/HhH
OB7XZlrWW/9s9HXWoCarmhR6/I3vM0rlCrKiEVqA0v4hu8j/+fzzYd9YLUhyoxsqPUnWgPMSBiFH
ceHFzQvbOq60gmxrFigS7cdes6f+2snEzFqHVLA33pp4TLirf+bR+Huk23M8SQsl0RcQ+pW1878z
IEQZhw+pMqBklnSuD4ED/4tf2NcC7I+dIBseappxBPRjZLedc4PMgYMwvdLYyY4t6UrXaepVitSO
iSAIqXx2Et8ykiNues/kz/fReH+cDGdtTrSrPJoMYJRrJd8S23w/WWjEZX25MybyNbFsfwPh6dJt
xn8XFQ4aiElv6niYiOd8rfK9nwqZWaeOG5+BjzyMPJjJsCNGU+wAgHjYFqIKYbBXbAzJNyAtf2BT
0ZY6OB35TC6dzJi/x9es+EA9TErBWJQQ9DHy/i7YYq1mKO1E2AnUUfYgwGdEafaGLmc9v9fHvJY0
5W+HoMJ5uX9GwPkrufGPF8WK9BK5z4zzHl9xtOFOecxVuNkadnlZc0ibk0jW8eKpTJaQya+prKJU
7FsDeFY63klx2eVGsrs3Y+xhTnaFvxWKIppsyo+vyGMMjm9RbcrlT2vyMnsCg0srfvLqU4ra8nuK
q33b3/EnivX7Ut2xEmhXDwJE9VcB+P7Ib47A5ctflGXFpNWmhuQrE7JfAuz+wKuNL0MXxLN0jXg0
AiDuHegPc676GfmjBA3SUqjI35wLhE7TEHvdUZsUaVmZKuXSLPXuFeTbRav7cAzp1tMC+M/jRcZ8
Tx+idHO4xUr5SAi1rOAlf41I7qPM6FG6NeXtIluNaAEr4JyYsCF0C0u9MyRP42JG7hrwdH92qY9W
lXQrfuUyxqMMiXejN8JRue0fCro9Jt6Uf1bLZiS0/+yMwgJP608eMzs+Lf4VDMSliyHDK/6RWste
tNnoC/YDAd+n33rd2zwonyeb/XsSY6EV0pataPqhEjN1Eex8JmHogcwGz5uBhVod5Fm1lT1KsVDi
sCWvL4rnWZzZjNvP6dJb1eYM/gts7JUEljnn7mIr0PrRSSaH/WoAjDkMJmLnwXwKSHX4rKvtvy6v
8QVcfDZeYAigbo9yNTVLvqr8wITB0+hFAprMFfUhDBrv7lVZVJRLZKARp2VUGkqKsGYvBtxKy9wK
J7JgxJRhkB9JP5ieJdlowRLNiQAXIifybZILQfk+HBLVpk0WT8x8sypXsCAIdijF2ux+RcTTFRL5
ikcbQw41fMg6KrpI/EP9al5WIbVEo08UFwNKBiPQEQ7oUylD8fEp3fYILONnCOTB4Te3kmDmt60M
OlTRtWZkvtrEEw4LIlkyGIN6jgPsc1CxjrdzqwqCRHY0YPnOQeHLIyzXhvkbQdUyFyDrwKG4IuBU
6Umu2xBvVFJf+T3PDJPJAFAZAmD0/t4G5Lo40+yZZx+ZIoJPb2BWTWPCMBEOb1Vrz1gQjf5q7CL6
/ozGCIr0rQ83feQzeyGWics/ln4N1Oj8XlZni6AAWCzIS0G+EMurNpGvzKOobWKbxswwgzU9FAbm
e4vXjQNTwvCIaMrJCrCZnNFFTCCcNdlhS6urE+zvmzNP3x+8xrNA+5kKBYDO1ZXrCJJUU3ydkk1/
YOJJMbowGFbAeYst9k2T6if7VEJS0KKnqiDzTOfNsQVwnsSn/Zoh0rRvld3nV56kFlVLLT4oMNMt
TrfHlhAe64UIfExUdj9kU0oGo7JGksi9iucBi4OZKUvvpYfMIwdVCRZapzm4lnVCBC+4qyy5FwTx
uWQ1oOtZ05ELmH9NcYpHsiWoaUecF4VnkaGG5TwcamUdBZkSv50gEWn519raDEjDVOWEdMiYjDcK
gjcDPnGJT8atn2uk9wVGvc5UOdwMOZW3rvq1VD0qglbIMNYehYtQ9GCUlA8WxPBL48rHCuQ6diK1
ZKA3jq1zgRAXN8G8O8rGDvHRQN/OBA8cMVq1FevwniYlyV1WFGvj/OkL9wvjbYiFrSR3uUJbOVCp
l6GeKVqdhXq8cFtylUGjupLK4wH4/zbrPXAOAYh9vzMAtU4sdcodRYacyzoFOmjYgHO4nZ+atXYE
OS0EjDHLuiZF9i/m8nUSqd/EUJZ0wOqAD08YnPl3cMRKZALLTK3PlY/ML/ge03XsIHnBoxDyN4iU
u/Y04MKC/Tq+dsNZAiFP6Z3twnZTHEdWFtSsc66diX2/6sp1URyd6nBhXYFCPbGCFDLfXPBlLdyw
tZmZbK1zBB4RZeMezkWjUGCMOcMotFRxBxAm9kD3Xtefc3awlL2cjnNkZAC0/PsXVeDhKvB4sfi7
hdllS0RgQjea8Qobf8FtJV1eB1HyDJf89A+LMVgH7o8CiOPaOWYM2JE8ORqH4L+dlbo0Qif7jDLj
PiGCYkvJcKX17JItcrpR/1+wGeUMrwYomyUMsOVHeacpNgfUPzkVcxx/m4FHUJOtBipDxEvCO6dh
KH+lgTaMCl1u4MfllT6WpQFTsRZzP3ObNEd2Kvqs+r2CKqwYSjoGr64pwUHF0bRnQQycm7zyFUwT
ZGZgfQtrMN0fYVJbA/4fYW9YzLfj9AR/qtbK7I0tTIQ6JMiYMGrhkra7Qo60jE1APoEtfdkOZdTs
y3usPHdU83BUFkUL0xH6Ks9+yrdnAx8nistrjcfEGQ+8vQU6dSpGRofEQ8Ppkrhs0NnT+NRQfdjO
mOGF1oBG9xWK17doaSy0Fr2VVNoNS+/QoltynanZf8yEuIdq/fXuYHARWLVjSjkW8GB27RBCL1az
A0eOwPNwiULrPctugQ5PZ5X4pG1xtA6KDyB9g9rClAKO6s/MZLI0QOy0GHtwIh6M0N3X7LdQTNXO
s+mxCnPYK7AsdY8Q2tJAhew38H8bf/MpKgDO5FNqeCWalO2s+wpZeg5uIF6CczZRUpH+GTvYsChd
00GH2MyttIu0JeWwDxgEnNCzWBSf2IKzj8/ww2i6odHfpcMwPRlhOBCM3oNA4AT/+ykVXPWLOMvB
dIit9CBzFLZKDxXczp21mQNC+GP6weD2ljOJiteRYo2fnKFQwx75z+NP+UY107O/FkyYMctP4fB5
5sVf7imGoSbG8nCKKSm1MsyoJJFrTJ3jQUy1634cgdzAq+owzpud6+z/M1PLBQaI+EmSd1touoDS
9dhWzAVk1+6ISWYjDnbPVZa4CL2H50OvrUycL9NdjghIrhVHGCp+t8P+vnUUeT7DbwwpZbnrtVW7
nYitg13DF+5fOxyMpgqmBmnsk44/I2gw7rn4cqRZzT0aMRHYaGahWszRy/haEAABxv1Us1yEBqG5
6HJEbqUG/zepbjiU//oMidj4aNUmfU0K3pfzOUW9FItSXSZrofeVPaetJ9xiYR167HIPk8wwo2wO
MM850/G3PzYd/5pmEB/A4DUgChI6pKw07EwCAl3U9dUAjrLTMr3szHgqslrhOx3TUEBNS0jtVPSO
oqnaEA5nRsnFaDi/1PgqLkehy9DOuQU9XhDHPoh4vWNt3I1/eV1qE6nwTM4FLN76ZbN4dEtsPpLX
A+Q8D568txoLpgaDUjddpyFqlQiXEBRG8jo7YHTqz90j9hY1ih1FN90U8m1mJ+4gYdzQkSr+P1IR
JAPymSOkcNXrJSu7uVqA27OV81hpDdNrF0vbFXiYO7zw8Pm/+fSvWmyCs237doPO25znK3kBFxXS
7Kyp+QlwsCm7CM76qzbSxYKTEPfyF50rCoCcgQserzzag1+gu9YoKLg4ppQFtWlflaLxGNxnGQy+
44OAhvQ+L2A9PJAGBhmPG1gIZPSDh92t1D50tmy+8JVxORDvrsHJmULW51CCsLYsSUcq5qIYM9YM
zTdunFNn5zKQg4ChzAv6RA6FOV53K9M7MzhM6U4ytSbbagmQK23rKTtMsFpU9TDOaZfDCfADzSsr
/asha5EfVSxfrtFrEtEA0r4ZCxr+OXNuyfDeIxEIzZL4Z/76+J3hoVZjG6rVeP9Tsp4+gUv+OT1g
Ey9BFymNropbc3QLxHMvahlkVQ9xPqhopJes6pzT8EpNGgPGGmkVOf04Gocl65j7Bzo2rgCpc48+
7nautuVGYZ00nTFLWgLIN5uMYLaXhnmiziHRWIvc3zEpTkEroXCF8qIiHCcaGenkT7C9Q1J60ADq
D15bcu3FH2EhjsU5ShfMBTw2H2zv6TtwUsJLGoxOhDbujCYsItnogSNnksTcL/S0YBlom/sYEFYo
ahpbWoR7bY5//+Ie+iemtd1Lb9ndDvk6kko1vz7swdSIFtyPWChmzcXbDNqFPjw3QAGU9jjv5jfi
S3+RZdmj03QtTFroyWenR7M9J1iKpP4KwH0+OrYuH0dBBNnQkn4nOZ/adLH2eJEBM5oqjy0x4Rs4
/KMqeUNY23JZWU5Bo/tkLx0kFfchCcideavlTO5n61tnRaCS1bIorhe6YZDQkiPSW67N2RpVe9ub
UBNyNt+WUc13HcWHloYIxoBRghZB/C4/InqnDvhOAAuzD9Y/mAixn1lHrR5acXLZmevu3Y2k+HcD
/eBFmgmS7hiUjrDOzdoCLKtsJ4tNcU7IcJUP0Q+6Zj/Jc3oQAZcOSKR7Kc50xTIEGiVTMLsalknc
h3s4DkX/Zbjr57h7j/dX5YLZUUEdRuB+cql+GB62A3k65ZFByxd/K2Ru93qHYniOaP8QmN+cEJuQ
0dNE87/qU4wZdS+Z0WHvcvTVfKN8spu0V4OK7xtwSN5PfWbBGD/U5TeSoOudrJDPA/HYXldpx8j5
TDXEK56zxjXleG2iSkTy05nWEWLSBujMC2zv21M0nYSP8JQdY8SLg7kPb1J51yuhmCFwFpDgibqu
MehWHG96lMUie0XBwb6Rug8XFpvdlCOLxDjqpvURTPwQcLevAhN9T0q66DVeGXVglfOs/+6CEszK
ctCTlroSx+94EyM8OinznftjjNlNdU5MlIg0UHgiVBQOjpplb3XXv1vceGfuF4STKx5zq4TCtbL7
LoQkFhVK68cXl99UTS/QDxMJr+l9YW5ISmc9zKUAGa/k4zq1J+5JXWIINbfe2dOXZMXFoKjDe3I/
sdq7bUiPm3RVcxaF4Wvc+jGhtJzyz8CYG62N19DO6/PstG7o/LbC6wWlyscHYtPbTd3N3TDHYY4M
M0NQr5vA7U0qREq7EuLDe9pHSKzDIXusjZWkmhF4mlxRQBIRIohUDXgOVrT8f+O9ObmrMByTlxyF
0JLbMyQ7Z3/FShLnM1KRnX+P3elCMaIWhtvfzsJbz8LN4E8KIkDV3eiVZuV6AVXaEVVe/7QjI2xC
v2D11v9W98WqDHZZTOOmz+uSfi+pnQal811eUxQX2TZSBGiEjHxtx1f3rdoNkxZSkpv4WpoW5Czs
YtpeL1ENgSmJIC3c+2a+zEGa35macxyDru2xi4Kh9Gx8vvFylTE99lylEoAx4HLjno4HHKc24vZ+
HS4yd5ZaNL4ebnDT90nPUp+PUR4EAJ83yu8E5Hc2Kja3xSIh9Nim6cc9x4WsU8lTlQAcWuoLS11Q
pkK5yGBXzBzTaw6RYm8LtUZTY0SoFhdZsa8MtXNkBhsFrAsNs6XD/Mc5Q6MSdbaw5Ah6VKmOlrs/
YFXYLHFpJlmRCqnQJk12Ckgx8fwJLBvryPZNmHXnVl+XII6FMGwe/6Q2FICr2W+zkd5gX7Kv/2sz
tUzVRFkEMxqvpjDQu+0CHlSh4/ITfN78hAjkE8K1neGmNgvtdJolq5qziuEMwdC9oEukDQVQHfEq
uXB1da2cCnXt0N46nC+kmDwRdx3FiBDZSEteN79Tim/gxKfscfJQtg3p2eNZx77IRmXisAW1N1Ia
XCHjmeqDCcBD92Ls5AyREjXx0Ox+pGDNptKKY8dFSrukS+lL7NznxxGDATV+Dgj7E8FTV5GmpqRE
jmixQLIbCqqt04QPLpT5wJEsqdrRsv6vzN5yUWbPT2Qb+7ri/iq9pJAJUP8iyX2/jc6y3hroQA2D
CrpgKuSigvOQHFZRWWn2JfIzPNIBPSo0+b2Dg8eWX8JLa1tvvs11noueP93zlvI6It7MY8cb3Yw5
xJdPMxx9oG6Fgyj3OB4IHMEpcZUhlSNLp0O+kuuelsHYdotFal3ffhf5QONc60dmH6PV6B9Ug7ON
pIv50+kcwuGNLw/ECKZ+AUwRRgiRoJk9wXfcmn9On0jEbTcsc8QOCdOkqf9pqvrlqK87M5iQqqHb
eRIwoId4SHQGLdldFNnlPaKfgT1cudKVukLdCa12RuCJIjxnpjL1f8AzdW2ts2VnpywE6pmeE1LS
lYe7GAbXdxqPM4gulLHlwdkI74bHDYumCcvJT0qTYiM44yc4FRz0kCVSu3wYAVF3IinhQ8vkDrwk
bD9IfwyH45HPYleqSamp/DVTzNxwsaw7ZV/EJeyYuh1+HEQN4wNIKmNIeCMyJ9O/yLLLC/w/VVDi
cLIIltJAx4lF5CxYsH9tiVG4FQ3Ji0WQevYcQyYIQcFilIxwj1pWRtHIARBWH0asq1/TrAJzjH+n
arPU99N9GuJDQrzivj8EklrXQzAWDISZJf3dUlDW1Exd8DHen8HYuDgnkTf5Vy+R6snv4Z49MqVU
HosZmbqFlkkcAfqEI+k3PPt1ayGWRl3ubJdZvrnaqaRtpqeTvncxPnvyZRKJgRt4gzPDXY5/uNpZ
5WuQN6OM9Ic97mCJxG9Tqv+tz5MAwJMTY7fY9Jw7xN3ihugLaLjTnPxuM8cRyJarZL/ZPTw17pJ0
Maj4BqO21EE6cnMfGNpfIOH6tF4/HbdE0UsXg1uCzc80mARIHVwj48Q3erToCCxa8X7M43+vB3yl
WeohB2+nd/ZdfFNoKK9N8o4R8DAg1zYs6jA8ytjqQTgKBtDYX+O880xDLCw11dxgChvvZtvov1so
UhiHw2B3L1udYD68NZzJ2ScuWoIto5WSKMnIMyPS3CMm0UMnOJ6NaJZqf5Vnw4xZ9J/0FeVmHbPh
NXA+zzTUExvmGBQGHS9e/bxRn1+TyVSJ5S/qFgB8qymskn2r15PFwmPg7JXrkb6hGauNQ+nIPcZc
m9yztFgDkD4QitMl/Gi1tBQ1jwV52/dup30C+UZiryrtIihlM5BmWlt1v/i3L9mV8RVUxaQzRyV0
tDxYC9zmGZ/fsRNMjDNi1xAcncR6ekZgiczqIh03G/VLvP/p0xj6E2J+Pjyr2qXRx9Y9uovfqR9p
LFf8yLrIswNsesP2f3TidnZqm40UAGYWlQXMBK2EDVcJtErzsKoogx13D2HD6FzUtmtDW+slt4AS
MiTTrCQYQCoRlNp7elL9lB8o+WVbqMObp5qe19VB7JLHaxAH/MYnAuE6iIUBrVKkt7PmfVY0GLxF
K4uoqHigTkJSscYtXVcmyOfhD13/Xl344CK/NFa29hd/ARPzWcK64SxZnIEDNmKINd9eWBY920qs
zeGRGo87ahDR3qnRK28DBAI/lGRZOmOxullM6Sw3BM16f4E6A0anXQI1aoVVxOGsFeDJvvFb+ZHP
6DY4PJJxTDfSU19EW27+loqSFFgYSm2588TbYlcGjt7K3pVE1MHRblkgYSk+JqimxA4Qg7//tRYW
h8glJhkqmJ76bZfTBMvkCOTWgD8BDz9xCSdm5YPKYwXY5O5a034ujjgKjlJdjM3fgDF+pU/O/DHo
ksT5fJJUaKeuKCgjfQsPCQL8QRHHLUdsQsJuVBA3CW7Z59UigBKtD0UqvRd2pEuZ51amSZyxHr/w
xh//A9AigSb1Ei6CCTuxNoKWJrCnw9XxoKsT+ITpEzAAw9UuNjX6bch4NC9ok/EpOFSdFxw2jRNo
J+Ztw0R/OEtNBCkDz5CA3BIQvRak9b4f1pr/TNG0JNvi3xRQez+vE1y0rLSxZrTqZSHub2gN03pq
/FgRWXmRZp4YL/kIcI9bPjvC+/BCHnE3qz2YEFay7ypCsbgmIIVWNevr140up+Uw2WfK/J11bTq/
lbsTqxO/LfPMPkx/tnJOX7N1wHJ7Dd2/r8cBLPqtyBqLIFQboutbbfBxXOIax+gdza00PfGbVw8h
7IuoaluDGtcLp4NMk1eV4qWDrq0WmkhRupWNNK5d43rtfpeLKlYBRtf6MHfQKyIithfPisysfL0k
3QDFXYj8YcpSV4dcIOxJnN0lVAR7eY1J9t+6/nsw+y03vGdZoB15prFqPrTiPvaoJfg6RuqvAO0g
t9RqAipliH1DaKJ3mxp1FvlAY5S55CbhpAQcaZaJuve+A2R6AymcSe+M4el4aY4e/D2fzxASZD75
XL0/Gut3ScJ8IQSpHEmqe+zQpUM1iQCLiwko2ZnhWTpbq7EvZrvyEpsn0TkzjZkl4Jl35pzWad9E
z6F+TZJ9vz92YhqqifTeAge3S+jsyur3Gs8lo7tvBOdVPeTGtuD9BhvDRIHagfS5rWlwiP9aHKm4
6XE1o1qIPnmMBIDjGHelajA5DRZlw6b+ykwUF8M+QU/UUUItOx6+ebJGF0huV+IuZcMzV5tpdP6n
iejqzI6Knj/FAyyY7GaKI+iSvnNq1i8RDhZO5CHMVcp2igcMc+VLRZEKGrl7Lk3exF5DYkLaOL8o
BxD9wiA/H9xczFYFuMkPfyy5tnDsHoisJiqzXw/ZoGbnf/UOBz0GqWcBVD6+SJvQ3oGQekXQo2Bk
+jRG9O0M6TNeRBVg80HRz83ujgB2eDpDUvb5Pq6JTzyeQaFdX2fsSNNmZv7CWWzFhgfqQfSzSB6d
Flsqomb0Y3GZTBCqAtoSvf7beK0emzxYE55rnt4J7G3fDtvRlajwqrJPNNBbBslVNxCnNSxLzv98
5q0csisT60hhDAxia6ngLAZEiOn+Z4qTDU4YreSFGZVQHS5xIg7Kz1YRbNFBbYGNFdJupAK16ox+
3EDD2WcZt11lT5zWUbjvQVeJcwOkl2Sr0HRS4g0wPlpBKaCPNNXmihwH90YxbjhhEHLisMMOzerC
SEg55ZtDnSAsfjic4Xh4rV7GAHo1nzT59FEDpbGuFlH3qZHdRkVAo6Jep3gSAXO2ijX1hPuXH7Je
6j+619CF1IWC96ytKd+wcsOYcM/e6brkFABAH+rhH3tcSa2+puwYVFk/ZfUw1ffDhNTL5PIAprQg
ITlMfHqkbQhkJJU0+pjbrIz+jofBpLprOYVbHTQzbABLTTA+TO5RIhb7tj63DJwPk613eRoDGjFH
hHI9ugmnth0Kr9wzhZbIgEOn6JW74BkTFuRjudVj12LYYZOZxtn0moFx6kfiI00+uUH1QGKfkF8o
yWoYbN3V8O4l9Mii7KKyJoramjrEIUX3EkqGtV1Ki4cXkm+28sQ7DxoZA+6LfdVAfiW172FNVZI4
L4cu65e4d3mHOw9Ys806VJAmrZ1cxLuC0pIue006EfVNXZygRy5P2Y+nArGvJjqq61dIfpwgqpmI
qua6CpLhNz1Mzqf8VhepobWMseBtmnnh8p47aTV3TcIbXlj8PBKKFG9tdokNUBOIslY2n7yO45qa
+PsjVCg2ci7yRoQQcB9D9unIAAzcC9lQRXL48oVDqhXDKZfcfysWcFGLolwFNwxoVBMjaohJSx1Y
a4SEmnTe4Jr5AV+tToXRG0ZPePgNUjqqlCezBswWC4EI9ZLnKye3SdHpZ31pNAfO4fQdE2WV5XWL
B6tKbB0Bn/UeTnwEkVLYyp6nmu0666sEAFDoBDCZHI0pM69M2khpOSeopx6MToFaw61L5nNIu6XH
69LWchuyTQD/adBPBeiHjA+xeET2hNYjtsJ3jdtaxirFuuSzK+PqzsL5FWx2MshETzgpWpZ5u7DG
6RrOK6qkg7u2I9BMMVACYnYMAIxFLYjFm24jc18l6ySOH7hTpiv3qKPbo85zHCBLhNqq4TjHXv6U
Z/KJpISBaYJ4PtXRN/oXPLVc/VX1X0cO2DYSX/dstE5979R1zJkr2/Vaa6VvR/kf2I6AD+/s6btB
zgIrdzimtJQlpIr3iahbGvXWjZK82lZ/S4UhvEypncL0HVJL7KEQqw3QMglHA9uZmPiVRiKf/ZWp
bSqU2E11uIPXFLTlid6h+tXzF3b9PqZiDD/7Ro+flg61SHVuWC9mn/Az0j06kFWSFJA81xTRYZFL
pXj9GC5zpQIvWndbQczv26QFAZ2ImRMyYgz26JvO0rYlfjRln5t1e8/OB6DMDKeqPCJkdjg1GnI7
n0bfOAzU+j+UDyquTLetBThq30drgk/jvVY9dSuJwWpwTg7z9/ob9NKPxb1WfykPvheynwc2E15p
WVn9Bgh0kpLqYRV3xlsod320ql01qNxwGgu2HvoIIpHRkxFj3GSLDb5IPcPq0O071lqZnrQM4hMT
pjN/fUqcLYkW1EI5+tNn+bnSsnn7wrHnH/Cf2+6ZUyxLxPijeqi8SAWInkgBkaFa5Ah/5U35ZuEx
YgbCzJAJconYfBYZjDPbldf/+kugcrA59ZH76K7PMl0xbRFNI9lXvf28PBTC8CvzrUJOY45XcvKk
wXX8mnvCaNksENT9ATFrga/X3Vr4swMquac+Ys0sYTzQ/F8IL/GddZI0Z/KZBs7mKEy343wZjqm1
P6V9e/+EE+R71kTT0RndFLdCe1dGohabM2c3FXCohgkehqhThKdDLIhlXN1OenzAtaMvdcaRVCN+
XtoR+W9QifFAG2Vp0JgclKVpqJWd7uTwDxqWa74H9iI4u5dp3NGEf+k91qd0sbm5MSzjpZg06151
FURVijd46p2SodRJvtoXSGJWiL8TACJ81/GtFS7uPGHY1ij0b/+sqFrmzVEXKvee/8mYLThxl0gp
lQL2E6/dOPzCn028sJYT8xTgmnFNc9cboR53sCA9pBasJqVqoOI2i+WWS3V5oEIc++89usyNpwqW
/s9Q+pPjJG2B/SG+UgPyuL7eSMwGpFsziNN28XGxnCzpJeFIwccTz9fW92fhJkPGlFNc84idpNob
+aOpCII8TSUC1kP5P16pXV8T3G1VuF7XUgYN9UeB1L+WI7gaFXvAz2YjVLZ43WhrpYkcOblj7EQW
jHmluKKC08M2IOYmazbptTF5ocktFmPlLZ8wCK5V6QfhXZwdEyaeKjoYAdZzqXddSQzZuPGvWWGQ
kqZMNqzRoxoU/XDZdqcbfBzi9JPnqVds4B8X22Y/CZLnFMvLlcqyGWjmnvbuX3/SD0B3NfctNAjp
iaa73ZwAhOAvw8SQwa1CsyprBZI1YGbaQuPqhOPvEiErI7jrZHa4+EXGXTU+kiwzcaqiD0cIbVOE
gRd0xgR0LL6oHu8xdoJQfaHcWveSCAQXnE4OvK0M1sxHEqWmwcLZ5EutxQ1UHjIoX+ip4UA6CfYR
QEIIwx1co7s7RZOJVQFfDJ/TUCl41owcV9uTz0w0qKtwV1fqA8icrzhMK7ElHk40BgX27thUGa4P
1LR+2Likqs5VTJ5X7KOmT5vVX3Fe7UUGGFmrIvxNELbpQ089MeZ2+x98hbly7V5tvCSpqW4uS6Qi
iEfFlKXyumdJCw3ytMGF0BrGDx1B5xbs/C54gSUxN1lBFyp5XqQYpym54z42BkiCaNK31O4ub8wW
xc05DMHWNyCyyVYv89meHJkNZdTKbIYO1i3Gt+TVTYuhhpZgwBWKbD39Yo2LoB8jGXEa15QFQURg
7kOfG+y348wmEqVVjYuTqvzcTTXl6bnvXmL/Jr5xpJksDvj6/B6WJm6kyKhfv5WILqSekc5bXS6O
4OfdtaWRVGtcn1I02vf6yr9due8B4mkf7+L1dWTuOyu7XAZMPpSrPIRESstzizI5QIu/iof6o7js
koZGIZrppqa0dNkuzlzEHAVnHJlW8Hn56nOEa/bFI6Pkb7YPRmPfluPuSniQHlGP4NKaqXU2UOzw
x72iJ+dTIFYwDihdftreIZWfmSgNtRxiuXIV1LUJ/l7U7QluARxdFULPkY3M/C8v8xVrBQDT4Hqp
2kk1r3Wn/C7czmrQ42Mym602c2DouesLN5jTn+1hvyeDagaI7vRoWowAsiRfkFh7wm9T7KiMbbjJ
WFDGqNldikIVIal7pGpSax5E8FVE8RO8R0fzDI7XYYi0w8W1uAkGYJpMJF+wjkf3xfiYzQlEkiHK
Tsh4xa5dGRHy9N5Y8JUqgl7Ct9yL57pxjn1/wTFh/+kK1DfqJGSPtI0V6ZJ4HaQYy/AfTBDeGwRD
P680PopAYV1HKh6Fa8rtCYe3v8Qq6KQSedcPdhGm7do8iOHouUaItxCPvP6trr2bn+y+Hael58xA
SN17+5VUqgkUOAivLFdZbFlojewTjvW9CrYWNJ8noe+BwMMvjgKV4K1fbfgOQ5BE0nRXoHjAHymW
By0il/bKLQeo7CxI4gHXXwd3RFqW96y/iQ96moglj09HB/aqBzjCDDG0u11+cZSw3dfm0+X/YYxU
i0su3J6yIZGto82IdTbsxTLHANuIbFrbU7zAPwzqk6Zni1hHOoN5fjPRB0MiVveShfX9PlJ8e1ec
eEufGpumWXZcJ7PS49wKnXWSdaIrGz667nW5x6wJWL6K3smsZL2osRAfqh4lXHX6zReuMMdER3Cg
m1A9hwiDn7VmyWuYRfGXf1E6xDNOgiR0dgbC5BZYxCUlqZKzegbmyJt6JyyqyG4vTs3iaFldAlVF
eN8R4M4hd31Sem5UwAJtukZtsH08kP+6f9+Q+EppoXJCZQEmzzZAng4S+FYcmbRKR5KUg8iOkW9q
1c1WC1ZB1NKergMhKjzXm8ZdOiEqQuEZjWNqiZ2a7ROUF1rfakEgz0bYK6Ntmicw0x/+l73vcPda
obh0JeHwrIAD0l6q/MFeIYzlR/ABjL/qTujW4eAXq9wyhLwtFwXzdDuJmKQUi6SovXZzqkKq5pWi
ysf4zhFPuT7lnUW7nbI/ITGAlnw6JITsVKahMNeQC003Tr9d4cWNHrlCUpyOvR0ftj+4xjIHjSYl
PIVq1G+162AYa7+Ii2utS8R2K4Gg6x7JVsp6mXLn6HvtC924Yz2qkX1DJ3OZ8QOWY7w6bMltrgtC
AilfNZoHIMBI1XwJwYy9grUA2zLR5c/gxKogjoegperHvwJAkzPXivZ6mgJ7Y5b3WTHgpfwLz0pF
4tYstraJC6DwHhchQftaqJEN/CedhZ98YkDXbE6U2lS+pUCvuxMPUpJH/ND2mL/p+jsiD9hlMY5Q
ppN60kX9Ry5f7rH13C7tdgyGaUnYlxDYAWltrT4wvd5rR/Ih3aFhkjEC38GB0Gm4VV7gLZdX7p9t
bKfT/C4OnGjsyCcHTQ9jofuzoFKWhA1f4jFpalTCEEkUrmvmt9Y0pJYxiYQM1l6xeSiSIOiQOGIE
CN7uelLaR6nEL9/ftDXshN6UQFkG2cgXgcEn8cUMmu7GDliYfIRBkj3xFTgB5HJlhlSjE4rX5rAf
s/s6SvIy9rfmi8fFTxMgwJE1JJN8JUg0MnV+/zxamUAvukoCsaxfNqTkqFKWSh7xN9ZfqAo6OKJY
OnbeeYrsLA9rnKTK4ait0Gxu3StKxnJc7v7peIBnPmSj1pITEQF6n7oes+OlQMVPyvLoHCOnVnM2
QWSUJ+pjUcqFLs9+B6v1g7dg00xW0/FL7u/2l4wSc63/jxboAcZud+L/8APMG/vUF7Ph82PkNcOm
TXvoP5iU1YQYL7jIvVrfO4I1+fVZ8jhoOVhZnRniQz8nQKbLCAcZIKg9bCfRviSlhnazIF9c+Eyr
J7BdFnsISapdswGmZKVdIH0RGXNH+TuaKFdXm9NWnrBzAOxJB6fIYiyaSVbekC724lYOZmj9FuJA
3Ac/OZsjwaAgMhEaAPIf8xmW0nO4cLuT0zORZ2mGmgluLKP4rP6kyWT5Y7yJrG5iq0dp4C2/sDwH
Sld8W7hMhIJaESfURxLpOv1Yxf/jLWoY7G2fEUeBC3VcRhdSEeljMeFPcytvxiqIIxITmrUPvFTB
MSVeBykhVZXh6yqK1v8g8ZFNnKiKr7nAllI/tU3hnAyiDaOhB/HiPMAuIitsAwyL/RZGblROtdHS
V8Wgg8/1d+7lClpyHXlKJxlNR7NQ7/JWQPmWIN0XwvLX5yERmUy4qZU7FLtP7Hktfdt8e0FPQe6i
4hY4kjGP3ANmMOn3BOtFQHq+w1cYGhNemf5oNTEXpDC1oV6szqvoLscIDN93gUefbnIjqtmUuHkw
XpUKj3NKWGci0TgLRFTSqUBlacaiIU8brlb4+RMs0aS8Ucpc/460jFaE1w3QfI5OP97xSEkyoRan
M2ZolwJc2CgykNzqZE78v57bkq/2/szslYVGzPVwAZS9bj4VTC9fV+KE+X3dJ3gWKE0z4JBW+UoJ
KAhfboD5hIHIE8/qqvxRkU082eNDuadxuukIZKDCFxwICIWfpSItPPoTLmv4zH2ZJ9mnITCli1gp
vGGb8QYOvBiGBe54ZEsz3Bk+HXdYhixKCXin1l5yatSAEUBmCqIfrrLnrLwdbb76I4gkZCfy7VeM
NgYhtjZnMk5SW5iRclJJI9+qnEi1cp0S2lp3VWeI1o79vOkc80AtnxgdSImO4yte9wmYoalydbSP
th2Lmj9X7PbgS+/J8WZPYYrbVV4bpqNWh97esbP1I/76zV6SKX9Tsb8c7AkaQLgnWYaR5GCB5Dnm
YJRFb2lm7EDLqqBoHSBXcuyOwdiN2/tzcmUVaXm+89fMwxKybU6cfVb/rNi38X8GMdih8UiQUYNu
4tTeo1JhpwIzGTwGV3cv3Dc/CmqX44ZyA2cqIYsT1iDslTcq5f1hmRMXQWc8Foo9DaoKeWlre4ZX
x8TYBPbLt19LUMJUwAPh0OOsKJIZMiGFB2jbbLHIB/IKGzZg+PT0K0bRXJZLZx9ZZxclSTe7cnb5
kNvqN0BTCZhTWv3CEp6M5HfZ9JQGiId35L7VppN/EcUTXCakDwOfsohW5KGBedd77HcXgdPN9gzl
+rSx0LQPeFY2Y4FlciuVgeFFuJaab9FVfoD5+Tqr9pX0yRQEMrI6q+ZvzEtKbYWFeHoAuSX1NnOX
iCmRUeWFWN4Cevlc2s/L4/9jArNBWKmobOesfWJFuGs/85iA7BevxWjqLItFsoFwvXzFQJY/7WKN
BarraRpNvDiaFupNxi73hIzOmFz8rjlPf62vNDjcL8qXibdDK/kGPxNvVsLfpVrmJ6fMLtMbKGi0
etxVuWzWPwQ/dknCDKXHwvXZykJohpzL3ywnyEwhwL5xPMNbh7dShlm2YzLXoq3JcAwrNPeanyr4
9vK1DiHARMTseVLVXHNscsypXcr/CLFGrlRKGZxnTg2V11K572MvhC3Fi3AiirRU5XCsFyzsvc81
MPBNEfROBa71etXhXjYSyH0IdsfZZKhEWu+GNW8FXULRBGtXShbb3G2CYuUcKPZ5MsewyefFXKyt
1jneNqGEIvcGh25jjtqkpu2LBES7o7xxj78/X/TgKKV+hIORWC1vWSVNhQyeIURzGBeO1SDAMBLW
TSszs8MJzSAeOuy6zJBPhDtdGr11Q5VFm07fEw4g57MZ/5uUqdkYgmyZ/+Ub1qNtq6WP1MYRNL21
Up/ZVni4nrKp2CaZ9XF0ml73OnzTMgEqolRGZbZI9lSc/QGOocPCbWH0bN1r4SOM6L0eJIEhQDrm
btONjycMLB0VHBWV/ealpesyorvYT7TFYRs75dmWjNeXOFOlwIlBkeL3KW4kAgIiJTEcU+K/Z+RG
Q+uu3k4lLmw2dHI4SMvSAyAiiSt925waBZxng/DFlzyhCBeUZaGllMXu5dOb3bXI9rpsFYWrwFTe
q472cOgx7qtlaO9HhxFZgirjvqLW7+wTdJLdLYgc9Nm4DdP1N7PUJH/gC4HQiIc3jZ9QLpYkbiFl
vFbJEJoyPufxMvGQSG2SzcKdDolMovQJZKBm9mUR16wFN8XtlKo4PDugy6+ZpNYxk2fsp+tYJewu
5A7r4dDVvOaHeO5tLAIzi1HQ2z0bGfnDIm3VfjxOfh/8eBvzy8gEis7gMjWlkizrWN2epbBf5mJb
BLS0FIQ1g4oaKrHgKdPPD3oHXFQzpaY+JHiUJinKf3oIMLoUM88DewgSwRjd1AyMiNc1f2EatcGX
ZkxIXa1xsJg2DKxI1OlVaterrsZRKWzrw0sNFIievSrOexjSKOukpfRvKtjNM+fYivX0Txlwr4S+
ow2ujdBXANCvbl6OOle8unxORJCi/SNSPUrdaXldV6KD4LDnvPa1VkRkuUAk+NivGOhU9yD2BSVE
lpwDMJbqXE5UADQYq9rDazGhyfin+faRtpO3KQRq/4giCbnGt1ty/FxAjTvrg0neG9+vEcUVxPkD
qDSwnkHZPC6qyuBDqUso29KPT6qlPzKCpzH/VoxmiceaZQLpVMVZvgCHc/EFwRBQeuI3v2QAGFoS
3D7/PVv+mw1MSCcUwWereGdk97L8eYetW+jjQDCLkV6aUr/V64j1P5D8+jxdB8gtFnrIXvTNSrp4
mY7eMmGQdLGASFIRH1330IgyWdN8VRx3cOOOUMBYvYsUXF/67LXCt8eRmQl9eRGKpGvqEqJY+I35
scBeWcQNm6XK5bFRuTujUtlGro7RHwpzKOidcXYBZ44k/+n+M/RnxTUnzj6idL/fl8Uh/d+Iig/V
qQq2NWgLUgqTHmdedJIzc/dLWsWdpDo9Yq49vzyukjFJZ8cM01BSpbxC1xzrY0sFk2bF5RASe995
VEfTbDkte2qOUw2N+TfTQdxjQfxa17jvJBNnY72kSr+8mRiHFAc/wn0K+fCkQOJkSyQYTEMyE4xJ
qYUYNDfWf8zS53pGeNP484tX0NHC9lQI4IQH9tn46ANCzNuJgtPikxhkx+/vQsR3TzxjxPh2rUo8
DJhyTKFlARAYO8byO/pHU4hDYFLS016Hu2SQFR9pNTkiP2a62ZIZcugp2u9aHtTdk1tVdg4zHGzV
YgKBM4Qjnv7ThM+7hGuAeQrR/uClHhIcNd/NdB6gyO9c8baXmSGxsH654noMCzgH4v8LdSyKt+fZ
SP5HtkLLtwocge4jJEFoog+Kx6b67HooNQSB1Z1Fei2ihrv+oC7JKKiVzIzxhd17L0yvanQWKvmV
z1A7NSgI+OoJIR5HsYqIZOuJsag930zHUAWegTziXDV1VeajkfOPJH+NoVN/0x7ouDsvgqNQv5Tc
ll+FHZpyZ0kcZlLIF8I88FkKnSphATd42KkO9dh+XZmcZbrPqv+r3cjbOz2pj0/Ek9dWWlYvCIIO
KhsWyayF0qZR7iASPPX3NnCek0sPMhnGNCaO7LIyCTT42tID2jNPmxcP2vD6EjqfraIMfB6LOspO
4vxqQC8py2DAMXmFmiewie5qbCzGqd8iQE4II700gfFqWkIkisHwKqmaeZznwsMaP3bZirkgeQ1K
QNYgz2Wts4jdmzObKiMzfIoOK1p0PwP/QcjMpfxhgXext4mum5rfSCnEPPNEYtD+WpVb1MQ68knD
Nd9KmKCX4ehQb63gkLyy1WjTGlKAPX0S/qyBFTy35QzQTeRjlev9NdQLl2MpY38RQlklJLBSlMQV
lFDfyp+yUbvXF6S7jLjcLTQMQAuDfR+Qr8pvgUcujdVocrsSHlCrbVbP6GBci6+VJFk2Tu0BP/IU
qvinc/+6Xf+Owt9y06be5kzIXcvIibJivxWkg/a4PleEKk8wP0YxHi1b76YMbf2IfiDcyD5WKmKk
L2tpv9rzWVxeH7EdOCX2EGSHTNSC856krNxKX8EHo7lAnTxNQDgqUevPO4wnGz8w+InFWcKPn1bY
emVQo9uyAMDssySIoVjCuSVfmWZlC+PXqUTpfxnJwR93dqlgfybh3GkXFYSl/a2tI8EX8cUg//Tu
640i4CmWh6WqdGbPUmgJc/wBv2FNxbhOAJv8Yir+UUjfeNVmzdvpBlGUTO1w73QGQs2zq7DLQSpa
kEu+vNKNAep0NuWVY9A2T2juEzmihVLsxuRCgG81HCGlDaRv2nO/KLlSSGZuptqCZVzhZH7ECfgM
ft0zuU2TKErUZMNKdOb4psJvfXx/Ul1yULuQby3Jxi5Q+GwkFsl0lvgAZ8Pw6ReE+tIRFZJIq2rp
7GRQgAAWILqgIDOmRuzlGsIaG7LBfWGSGJVZev4LdVMC4nwqRG85Jn9UoNQFMwUI4DnvYE2ZOyAJ
B31MjCUd/YMIt7PF5oQ7rPRT1Z4rIgTPgmyPCcAeBhYw3PYq20RzCmsHPKLPSZJm/+VITefORB+H
mEvYnADCm9Z3VWY7lX75z++3HttoSUoxrVi0P7ji8lRdN4FBvLQco48Qn8MVvW31uydfZgjJEuab
pDoGJLXdxR0SBFuJKoBTc7IMfCz9EYvf7LLVuz0pZ1ldfywO25dRhx137AT+sA2oAsqVnokeyTue
GeWDl/HgCN2f+LnMsmL67iS9rGr7KAqFoyO9pRfBS1M8GxGL/EQQAwiTXOnQ1I4gwAmgF7eLGupp
4S5b5dQTSA4XV08ANQfG/mBhSB+e1A1Gp6s7Uxrg0nr7PtuvSC45EUlytbn3ZbGeFzePnpEXpcmQ
LMTzVTh28F6vQSA6XQMr9aVJdDJb4SuclMTDdx6QWig69X2hK1VkJ8/fSkpTXqhoerQLd7GZ6fVT
8Hg552L5zO/7YMyCnLRrO63LlxAUhzAMXAR96++9b/CZSVggNeYbqEI4iaZuND7vkdcaDF8iX0bk
XsnzG4rKEFlI2kaBbk/Vo46G/97jg3pSE0M1YxEFXEkfeqp240P/ltv9rjuQ9MbfvDwvnApISF8j
4TzsPo1PvIWCrmQdhnhBWMrxCR70ThGddyT87t2FFsh17TCWmyw9eeHRrmDiP12yZRuG3/9TRkf6
cbGkT4EUjsdfTQfSyKCRP35ENKAiA5XokUPGqQKZcSjcdn+typLa/n2e2yjdbYAhTOq3m4RnslQa
kXvpAnwxLxA7DXk9lUuJJbdw/DaJRgCqs5fC8U9xPRnXDmeYZ+rQS+3iWuMXNqEFB9EYhexRqrpt
lsodF/mE5Sf2q57OKKbGjeRHTBJAPAaahXq45WyluB/wauccb71tkxoNe1jg+4a69pWKZ1VXAZms
rA56WUShpdsDPGvl4ihxRDyNq1ZCpxjJ5c/VadTUpYjqwzZDYK41cNaV19M/hItmbrRkmTtzYGFY
JACTy7sO1YtBFtXYYvPc+QCWxQ+EzNPbvSr90USXzJtzVDMb7armWhU3oWHqhhdkgidhQtKwXJho
yNPMX6Tin4VCQ+7Z2rCB3l0EUdTeRJnTHjA7lIz4RMsppp5jdOrtIPSIjwWjDFo8VJXQVn/UGTER
2dw9q6ADqGRo5gq6XXH2YgkHqzxhxl85IR8tJCmKaehUlTiwKHeEV/e9DpkldMfp0o+E8p+Plob0
c+hoNT2WDONIoB9HkTPs8nSBDcP14VjYfOkc2ZuxbHx1ZvskRFyZK85qpwJSBccm0gVMAk4oir9n
x3M8ephk7tlR98SY10jcHtUaTrEkTe87DFfE/d5g5spUcNwjCe8h9MFRD6YOiZwiOpDSgdm9e05K
LUo+2TbjV2BUyDr1E0YHZ1QTqVkB2c2GOwJNn+9wdCbNN/CdvMyoMb4TXQ/bH+OH8ZeamI4YP2MS
R8oS4yNHik2mZZpUlU2QEKyOWS+nl64aWNGo5AxXKWQPPhOiaXrqDKM0AycHP3xgvfEgjE2cyBma
SF297JWwaA1o7ga4IEPuOo4VBls1qttMNJlvoEMydSRPubNDMGu3Fp+7oRdh0WVGTt6ovaZeCpnz
X/iOdid41/tUhEAuqjPz5Fm4Shzm0AzeukPgrHyiRJfa6OhigHMLzbTVOt+VsfH9xraMJXqB2fL4
8qS73m4ge+ncbYN7R2Pjgj1BOmVPWvW9dljj6kxuvXUzhuZ38t3VMb3b+cqVRRsDrHpEXMfVT9RH
9QdYLeXNAyDY4AMwUqlOmyf6XbLqZuPv2BMc2UQzFGp5mGSKTXcof+rjTwJQN/U+qx6XHV/LfUF9
ob22447JSz7Zpf6ZQs5IkiJFQQPf+9vH9Il2qeDVKjV2x2U6C9sO9GDhahij9J/Ukw7XBWwdrIL/
ju5UlYks5EKsJMNhBGv0Ec+/+MRSETKpPAA76PlN5JsS6ifQElmAnQa5seR5cALfsu18dezCzM4T
+ELTaahMVXtvdqlJ8+6jyq9Nmh/eltjr2SjPVvusOfsrFK14RLv5NFXqYDQrsM5ep2EFuKuyQGh6
LP3fQcZjQbEhNqVVtzBP8U2Zhzbpyait8RGqkWsbLfuCMVMIBzCk9bDu34urqnbUjZjTXX83Moct
aML+EqIUQgMwkjWyVgfosx+ZrnZ2AmR/Yg58tST29TkF8xpR/Gmu8BNbWDCT1yIj1dZXlL2pWNTs
PquxjIJf9lMvPsEWhRspQp4WHXN4A5k94dCX3kXNE08kteawuzLG47jY+3f37iWQrMbyKM23RLdM
uRJi1m53Ezg8AEtN2hOBrs2PqigiGDOXaN7/bEovMeiMlWl+AOGv0cZ0dJ1Wz41Z+UbGRV6dfbTu
mZrteWR5wzaSW4gmIfESO2QDi5wp/EX8vKJxddoVWD0IfufYI++cfPTVhMBFxzSWH05j7dkP3bym
sZH30B/S6d5OJnRgP1pTalcb7QCIR5m3BKivvJPXgb8vcJ7cAvqY/uhYQESkaHgtwdMLelbAs8iy
1QrHRqBPjM8SOhw79i/ywBxlg0Jy9Ce+ToHNgpZrm6FxkgHK3gOW8j4xFj4h0GrgVe9mVWDIZaiX
lXTqVjVq5bJUdq2yJwSkYxVia27GCri2JcomW8AYQnxZMJF8fMV3q98z4N8iMCJv2vH1rdDxULMv
hcXJ0eRCUfrGtTRf5eadc9k9i9vZ27vpkoLjdQuZyukUuyMQaIoXf46Y9Yey66VXmaETfB3ADz4L
RSnbMgU50CMd0EhSmaYHd07zvO7kBq5Kj2EgnanKAvyZJPHbBROBDyY/nLhEbZZGuWDlPk1mD42s
aoobXNxuOFoniLO8DDhQrz9mLJCn8d4lDBt6USmg7Fq0fir/rkLPU+JulwIu+KlYrMSCpHUj8OKq
FLczfy/yDaPByyXPN0CN6Nv5WSN1zonUuaFSXkBu+gQ5gu9vQt6ITiV+/FYceCiRFZEYnzxEv9Yq
8FvUKCGrbStGlCggwVHieqwcSocDss7EhCpeCqk7IBs3aKcUrz773gJBcmYnyCfYittFN/fQmFvd
YUEKvBDuZheGDuSCx7VuhY96TLF83Lsj0Urf3rJKnVqanGyiBCjL11odzzyx5zZaY3Oiwt4hrI8r
WCWnnRonY2pW0jtmQEWVHAiPgGFSDFGhu+k8PUZH+OHeKuEPR++XdpNOmYmnJnmDWFH+TYh2RlyD
L+/W/Qe/9JAbR8398ixH2xPsXvi1HZCLWFwKN8rjucdR03Bn+tTEVI1yTAzpI7BzyQGMOswKEwSo
lbBwL2U/J9is9ZCAleB5ltNtDAWP/dpKRYmqPA3Np7zCqiIBJ4BJ2cq+YrDhZSvdhwNXobKzzZFy
1AsmWplHzD6s/4y4AcO8If4Qvdc6twzqHBeGgyjbEyVZcEcverVqvXmhmJ8ejWfK4tmD/KEGNb+x
8YqYYW5LCHIOlndo1aARk8e6gMEuyl4iIQwpoxaysSowKy3TYVHz2ph4siRFUJcmqo2oN7yI3BFH
6bRM/YuDl8RtESwJjqdgkS8ysH8KDMHruFwwcDa1I9ScOqmG+L28NWOCVnsVUHMJnBJamVjJs0BE
eWk6pVyDWx418tSSN05l3gBmDNJX6LGSUvThWQOqMUTNU2s9gymnnLAMDfxDGQucdhryc4wpFjsG
xhZDlrtXxEGaA2zJOaD5cS+NrT7V8iWIt8yiabWE1v5CnpHHsiUHJbvIODrhVr1eVoIwvjK6J9tY
XN5j/QYPNNJz0LhWKTYZRBOnkZsRQtdJpUMmkWwBcKDg5Gqktramovcez/plJmcndGDu1sddODqq
vaAUS9U1LRd8WCvpY2OWy8IPvyeE7VvIlsuNdz1W3gx5YCgZxlRLxOJao1NiFeOflg4NYYXxLmr4
R1Qy41cQjH920vfxF1pvetkr2TrQ0Gog4wHNjKFWS3CuFmj5FT/OoZ90mDTKznmjAZGoFdtkvh54
d6sMQHoDH329n/6+O5qq/afT/Q/dDSYJ4A1Q3uPotBuZoZdNbCMtwFYyXm1AQjriad/ByIOBIPE1
E8smXPNBrFIfx8f7wQn93FBJDUgWfgp84xo6VKh0S4GLfgzLab67olBOXCVqjaRjpRRXdApUGWhy
PSxwYdJsa+Dh7bPfAY+6byz9gSYlMyFabt2qj9Y6Oiav/CHEjbxdylTPWTByvhTqnMFQUTsswYIM
xk8x2wvQaAefMQq8fddcCdUB38qvrqNW0XyepqSFktOG3lTvgfCCBqV/tmmpYCNeuNyIRzFWcNH6
/QJg+YmFpBqPZYVFsVc5fs3thclOh7GMU0HJrvMuXPkqlm56oFM3ZAVlbUHNkJWenDdg7m3T7H3s
nBV7I3WxilwRVOuSJoQLAUuEN3a0hD6p8yn9yxGPiBxBnvpWi7iBMeT+3cPFxRuS7TMem7aZQkPA
UuTy6IW+tZiYAx42g8X9X0p0WeEH4hP1Lsuk5cIxkIYqPYSnDJj28X4GDzLQqt+15zZI+2InTYQ3
uAjTjNMlmQK7Y/VbxOjx59Y6c2kppnKyQGEVYPEbjHkMBt8WKCyCq66zszv9RBTmvykg+0fvd7Ix
vpOoy3h3TqTYfzh8uNoN7DwSUlx7AJ4n0HSCiLiQ7KnWRGZIfaZU5e61CRpDCZmwkkUeOgHtsiqM
/AW41TeXwYJj7QB56sjMZGEye1vUZqAX3c4b/vQap9tW2ReY7qs61RutIfpzgRrSYwuqqS1Wz9f8
hFQBuJURs4uZj6DWag6mzZdT6WTZBUvbEnUsv0ep0L3WRgxWls2+fXfY+alhbg6BBjmooyKKWjvs
0quMAHw7+o2fJs59DviTYqfwTDReM5xpG+jiASKTdHS87lokpD47cfoe6huKiAv9sbJJBSXkc5Oq
Rc4AcgLlSdrMygmT8nZvMVKfBF5BMMW5vkIfaPBJ78TVqGqTv2vXs/r0lXNFqcsuEzdTpD6+hEEB
M5twyTp6DtE/IQ2IYwLy54gHjO2hECLBR99IL2gMOHrMBYrXE/olo9KJRDkXNZfdzkvE0C1NRd6a
YJCTGwC30yWvwQofBXuw52EQbpjVNv3Kp5Om58p2gFsaYNjdRULnSsCXMbsm48kgbGbCTYBxaZi3
+otMj9wI0xPUcmtfLslMWZ22WfPIWDH0l1Xp3uqAXDTYk53ZzRJ/cIYPwqcMDej5WL5gtAwgh+gf
s4Gmo/GuFB3oDPtHDMwxPTGChFx967bzRro40zyaQWHiVjyLOsxSHN831PVcqDQDMmaSF6ADXMiO
MFzPOrmhqlA94p5L7WM/EmExqLGQl/RYKbXMAfBKmJ6lTob063aaJLK4ILZ6Pmlb2PZ6vRmRZlCZ
NowMsaL/gio3eVql9XGNq1k0XjMHYT2FNTJdfJpY2J9L7yuzmSr9crHOOY05A/mN4Iq8i76fKo4z
oB534stiBPG+SUlGCR8gYZ/aG267bTFUoP50knNhSfQMQ9WNICOenSBRytWLsYYo8reOE2612h5f
5wWtRb9Tit96kIdG/LeDKrhlI0Zfg4LemZCeTE7pTblh4FsEt9DOXhDzmXR0YSwBRE1/uZGHunAz
CN1ha9gPLSrSStSb6LN/yfuuRWZGe9gNTZS7kiKM8ivpblACAkmh+bhABGrvU6yM5iV1OKi5K4Wi
C7UkYVqoX+yErg5oG7IuLr5vQKgBfwWkGuugbjrFyo5wHCVOFtZmP3jUsIqYse/b32Dm4fGUsWNO
53aOyw26ZP14QjX1gDy8xWaPohzwgUTR+NDopBfZjhyqspuRedk6ZnwzRyf0hBdndK+Z8Fi2C6O0
2qNoKyigjwBcO1V3r7uarVTeeHcId3+z8Ub4TjPcFmKjIWlkvuY0IZCiPsVkqg9CXxIqShpt4oww
IGFvA3d8SrGCpUX23dNVJcWxQOm8jwDgLW6YyYMRsyRdMdzoNDdRFIG5RIGodvOZ70Y8aFZBF3O9
tBzsYZqOTQcXZlqZLplWrjtRqfTqg/bKWIdTaEb5ggxHBSrWWuP/s966Us+5NqhGKfodDs2VgzrA
g5CVcpnJzW9EkAGTbbCoOMjembg0gz/7pgzpC6ABW7l/dlr04FVIOGJbclrQnzaFMFw7j9lXYf3N
0w2/VqJz81t61gxueD3IpyZVokcnQW6SqctybKlPGBwmWZtGMThVAUMcj9QOm6NtvmpqybEQUoHr
Q/kx/DZ2dbs8UaMLBRITvD0VDdtCBR68gykfSXOXIHuiYlpodr7LQB07PMK2Mx0SULoDA/r7US5I
t5dBo35HWPU4Aop3wd6UDCRMtl/geQuDZEYe3IEWAiHoA3sa+AqxOaoUhIn7tuBDx1vG4ej/GyWx
+fjeh1ItreSL9jDTNGVIG+/Wk4PxEhC25nqAtO3aeLY6i5GpD/RQeKCoWFeui8jmqng6EKG1k7YJ
evMUL2VZ0QYxNPbtOaAke/7r2HZ1WsxIFq3T22qm+BJEvGu+eVPqlJX8YXFxkiWwmrPAEV8ftZIL
50L+0mMuQ2ynsTFkXaXLwqGb8KYgNZFx01IXE9uvoHnEljlhrbGNs9pPGZHpPCpi/+cX5qLGa+7j
xPWzuqQhHW9x3moCXRgQ27hg0n4A7UB8dPpzkv1Qt5zfx1CbX/d1rM5nkaWneqSIOjZEUqOznxyY
7h6ibrGStGCoAts3ypT0rDxit54+qd6UMhVVzPIyz7g5M3jhqxvXqHKR+1mRoMV0w6Gc8mlCY+6H
AMIccimsKRUkFYzIFQXzOjSTu6bt0yZZJWsA9+CciHscaMw6bhG0wmsoHC0wWKCxrxIsXzhcqVEq
6J3cmCwagU3D78Ymdfr4dv4aPEgDSm+qhspBygO16xDDRzl2J12dJvz4lWM23J3fbycf0+UfvvIT
StwocfhW9v2dMh5jDkKqdKis7OES/OosoJx1EZ5AkRlUXmTuVSnR9Poh2SYikkT3FWhw88GT0h+I
DEocU+mYUczg+tO0aiqCK8M6C/+Ni3l0vFBC45NQEj9rWWgFX3k1XDv+UfYju1cLMdE/bio3vdcb
IQ3DK+lljioOKES+5AZsgNHqC+K9RG1j5mrE0G8vjHw0Xs8kHmdCyIOz//xIyGQgBx3XZ87zdoYT
LQjgzRHzF4WBIcFwyuXf21Koe1PIHj3SS3FdCGARMjsPMo3LYU4trcYNggDXupMYyNM1mZXvq+3W
xJik8CSrPtSnfR9Bk9pwZP7h0DY4Ea9zv27oJGGBe519Ch7TrSVX4Jc5Lj93kM08PtHxZjDuLzS1
s5NGN+ygKLYgbP4xmhNZ+ToLJFZZvOyZMPOwvOtk8R4AXrVR0OHP8KhDx3o/lKjiCf5kXgjSHgV8
KGAcNKIPS8NGXYPHXZ3hYSzBQ0+Eh4glvUVWQUmOnbD7BYRQtpMNbGbpIxfeZP51b+B87CddD7nx
Z8Ty3zfSVplfzLQvrYtKZ8U8RKEEHPw7cFLlLQIpkzhvpP48ws/enhmCSJ3rrJhRcwuCR1iGlBNZ
5hidGC49/U36C7r7gr3oaEw4PNvNdS+L2DISVJwpgMCF19FwfLKkst5MiJW+1+p/c33oHEGwHCFA
mhXN3WC5mG5Tz9LQD6JTl/pRokZzxl3ynK63gUqT3JyEjWUy9RP1ivqXPs6mz2od0vUWdeBzZRMG
m2pZ8hpTIo1Fi0jXrUetzBGUPqLwX3LZXDVUMKVs5m23wwPxBYyQXNy1j5Nkf4BylnQ0WES/4q8g
bnQlq2jXDuaQ4LWVQuaelexCJAhhkBFMkmWyKCSwBG02yp128/RDqacn+FITUWDaZySVhNzFigtN
VUSRD8eGY7cSTyIKeNtZNWwQBYOmRyz2RfTTRQy93nKeYr5QUs5ecfsjGhxpucwivPtKZAkMvDic
RhKm/YtJ1qhNQ8uGGaV4Rbu2m1B4t9fUiFThhY+6r3YXLFlQH5Tmt8qNkxJ08bEgiBShafhqLb8K
BV4CylcvR4XiKCkypx+N2QevH+msSkCLlK6LHPbygqSxc50hh40YwV7L5oI8tJ7M4qBenBkQmvnh
89c2i/Hdxj/KhvpXLa8Qyyn/F/pOfgPBhLQbtKDqLCQyvT/Qi69c45mTpLd2+HJN813DAYCb17DG
jiPhrJ5OUE8XN4at4jW30U+yCw7RXPNcPgJxu+aQ2Eht5n3PSpdKChhKMEBZyVEspnFYjMjip5No
HhwR2mRRuP8796cKL+p0Wm0Nh/DBNMLecD+tV3MdE8BWQMpW6eEuIRxw6WjyAecW4qf5YdzDW+e1
j7uAMVE5Lvbl8Jq/5FbGGTw22363S7LG7GFh2NT9cICqhuFBCJqiVVLbSy/cWgoucHb4hwrD474/
JTlYUHJ2tNO1fUqp3y7PyRyQWAnzLfsJEO6r+GquOJ6vbNR5sPLdFnTMC6z6QuiZYtiz3G+L5FKx
ytIFKev3URkrYbYk5fEngRyFpm2ulC25PrqN+dYZLQz4ED7P4Vs5AE5epE7LqAcQWMzxNaW2OlTu
ya8aRy6M78HqXMVOHCTeXuUqy/A5o7cTxCBfurBbGq4563NxTWwQG4p2KVmYYY6awuIz13vJCjQy
uUS4VR9JutJ7mZOz84rHkisgeo8Jxy6VXiADg65vrsAIpXbsphGY3wUtv3xqScCqTCF1nxwSqzu2
OHCZDL8uylsa2Vx/qG+HT1crCeU6PRWDoXxjEvn62mNqWV2Zr4NTizpQEWfS655RecM2BFfQCsQd
b2q282F8/WW9xtDUUU8e38OVD+o6R9uVue667JSJKgQjafm4EaSm7tZhEinKNabWoOs77QV82tTG
OKmERWQkQ/wSNUVhYl+NPWk7DFqkGsc6i60s5IqFSVB/vDUShjoZAXn0zZkLgY7XBW7FV9g7zyNz
3uWQfZUe95bPHuEftvHXCUzqJ7CyHg7g7kK4mEz+UqORBIrf+LcuaHkLmULN2g1j3OYUykx0f068
7+OSIjMiqxDvFcSENQGXKPdhhA79vmHXU9amX5fKjM9kEaKK5uJEDaZBxwnl48o/3DHJ29K+oZu7
nypxgaz1/5j2sARE9qoE2rUd2cdE84zoy/I9rusP/QTIP8KGj2BJ/xa6sPXEqO9qWt6plA7w7Iad
W5i9JGB8E/VJlKxpXhtwq4FifaRe6deka1NSXle7N1otA8R4FAd8ppKvOsig/Rem5+Hw0qUsfRnI
vlMFUczdy6WCsdqc6pyM/5AAKdosBTTxLQJEhHtMiGajoyry4plwA0zlNeucT68QRg8nWxLF4pJ9
FymJhVlTyW9rHbidyIZluwMBDHYMeCL3RsysLgz/rdvAeYQQIedf+O69VGl2Vq1wrIcoHOtC/fW1
nHo2ckxmWF5CEThbNpPVYv9h9fe38jtuDd6oqxk2S5UP5lPGq4hNmEcCuW1MrkOO9flXPp71KipQ
UTv7ChX3BqrxRqO4SXqR8GDF1RR2VesqIURn0V0UBYwwoKHM1Kqprhhl91BuZ085NxTZWglgcYMs
OiW3KKMZW/WPFpJm3Tpi8Q5cTeZZOhdIxmMa53zhJe9DeRpJp0d2Vnh8cxiQdbcP57LSy90dMsuU
56gBk4mU26i+WFnYK26mbz/YoMu6n+QCxOd6NYJ/QaSDYU/qlTaexPs+CLPuGIWOMMpf3eEgM381
hcT85R0WzQ2aRrqSablmSEGD0Sd9qU7altRT3OFxwIydAuKJ174dBLczROxbT2yxb0grE3ZFYwQ7
yVfhN41fTvgcxHfp+wP7SAGAdhPcDN4yIY/eDbz9uNGmi/j1zk/tCBzlbmEiDEmkdFEpMtFPVNBs
mKsyXjrMdrGd8n+DIv/woPd8uWAaaOhvbt50OWpMRNSU1m2F44Ak8n5bjhDRjc4Sa1JC4ydiBoff
MRGIoW38tE6V1G0cX8YoEWYMjmAt7wL3+ZrDfvyUGMwZZMjcpxqvI9DFNjqMi+rxXCv/ouhM4YIM
LpsPVC9i9g+lLGfGDXXDPR1mb/lc+8aa+QffDvzJablF3uI8bB6g6sokDBauiKL28hph6H6B9Bji
mMGSxY+4kt2hlJIANjJQMaMZbJJNzBbYj7rBBVHe1Yf3pf8QucwTv2qgb+2NWfgcc2NJMosVSAFK
rt+CaXp3kRknMK0YXMjH9XgQydwzEgaa9naNX6I2a0toAKZaEm0epFRwwL3oXw/yESEJh+tRJoQB
OSJjMn/GyGGo3kHTt2bOQSIuvKg146eHJq/xNgtdX8Vw5iOd3mva7UL4yIT5ow8S9uD4XFVae5Tr
v/9SIMVM/P/v84qaWR/QHq/Fp93ZGQrXrM+KDjxvbSfuelBuHLwV+LiKLHhBjk92jTJQb9WTwRfc
sy7oPVytFzPqh3iQca+L3SbXKpjOok01geizCGSXMYCx+yjogjN8uQ/MzjiYYKQ+iAzT7gkYVtfY
WGOKoC76BRYg4ow88kx7QirHwDNYUwEtG1uXfB7mnIgrOWCZUk4ctDc0NE7CStMIujh5Vbu30y0B
NS0UxXM6GXraaRT44o9VcVHsDfMecdfSOn/FQCxmafTElBFb103gdNViZGt4A3rexb4Xkq4LJ+os
tERJUJF4YheIAJVvl+DGEjOqtKpvHpGgVhyhJEhEVOdoKyEt9icELj43NanuMFUXufuEC+0Ghgbs
DZCUZFTXHJI5bKZp5Axi6O80kVpl0Xv/RyowauqBTMckdtOWmTgxghSM+7qUaZI9Ikp8W4gdwHry
LG8MO+3WaGUZSVqxX/Shon8tk/pLsrOymslotF9jihJvAY1K8Nvy9qBtnOvCakYbeVT4lfsIgXaO
tMdZ043wLJOBMc2GJxaUwJC4ayktkShz3DK9hulyq65bwWtiKYpql8fliyCCuE8OdNDgieOYJt+c
So1POQbMlUHp/MfBJDKV22eSgu3FAzekDaoSo8izSK8sRyJBgG96m0JT3gpj0dW1pc8fqYHRim8o
lGIrRkWPRiswb56UQeQQwRt8w32tw96WVMR5BgNSVcMNVnq2fXu/qXsZFcDLFVZ40JtrmaWcypv1
k8Lwmu9RTiuuYCG2h/pKwb8uOyky3vK0nVuD6vu/jql14d4nzz1sBcaK7awrvwdQnZBQ8e3Fmwlf
kPqMEq53MJM262YNxBc+godv099pKgu0WImLdjHGlijla8WLMkJ6FzoAdSbx+8Er7sPpxvewHkcM
iDPXaquvGDUMHrcOD1SDj70tv6Ij2esApbLh8yyqxbJRoG3nssG0DtbsTLub+9PcPeK8d5rgmD8A
ogP76LVztb50qKfY7GndTLe1vM50wtntMC3Q0LDqMB1WGo/EdpdYdHo5RMJaGfNLYw+Exlhz9uxt
Z2pVLyKWxHh/MiMJcSItndIrwRlA4sC3GpcxXN3FdVNtv5c1vHYpfXy14uPIamaFlUGYMKUtQoR7
9Ghq4sBNmz24GxZ+CeKP28ezffnRgNo63Yd9ArYCnMEKZxNQdu4ryDuM9iN9xv2SUGWsagVDMXjD
Q7Op4gTgzWku0mQbdNIdzcKYeaxRfNRcMbgHrFEu7MLuQYqLYtWpEq7GVZH0KSul/SIwcZl7u7Pr
5XDtQ3UWRNiPZfaB0SkfzPukBsxPfoFIWjoDxfw1Glhzi3370qkShl6x35qCVQ5YPewZ2Ui3GPPN
T5sPtDa5MbxPJS1wtXp11NKWQ4oUKkKTvBpbjTjHx6OAw1oZWh8sTY9WaHUl39oc2bASG/nKAAmX
ublezaWmoPKXnb2MSp/7yz++xJ9X4a513IsiKbuzz/8QOvWJHjiWyB0aikxBijzl7b63DHuanCFD
0QGkPNXeYAwza221dOVPTITW/Fqb2C6i9LLEiZvyl9NIXXWN5xByCHiDa6egDmDCviweswRzq0DU
HjtgKNnMS5MTZR+wIvjFPsNYT/R4JriT8LV3oER7JJ2Xhiu8jw746inI3n/6m7BzSM9OcG7mII6M
7VVUP6nX+AqeNgmkJfFY7LrELrF7FMdX5p9sLc2HfE1cV5pNad7y2WX6c8dR7WEqIWIQCHSyO0Kv
wBIP6pUsxlnIDe34LIe/6ewTIbp3HTVNQfK7I0EFJRnGNUSMblIDcFYgdEghESgFPfD+3TnodrGt
nl/FjU10d6uHyt9ZUWFueeCL0WrV+LbhBuYvEt3clx1bkznyGbJs2eh80WO5CUKu25hw0a78ulG2
Irh/8OzwYY1sj3uHusXgBsJtu/+SsuT+1FOhBpIr7Xg9PfQGwGVZNWOLXJTqeVDhxOpXwwjlL4a4
NWaiFYJYkAuiNBeQAS45IKMig/cDxkvOm9sqxen0SNw1qXTNpgpW4BItiqCAPIvlAJT7/8xHd/sv
Wh2K0PCjg38Xr98CqOROkG3bInEVe3JM5Eo7MV0vE764No6vO0F7lNC1tWhpQg2z9AXgHIRQmhs/
rsetN/m6DhUWfGAcKu0nq/sv8/SFtMcWVu6xRyBrjU+D+j65/3ogEv9T+DIl36BXh840dFIVqNmj
DayuBe+NY9Aux1ztT5Iq5RiqkiOvlE1gXUq7S1pxUniMrFuCIs1+jlP4F9kL6KiEXyFGdaHEr+WD
lTqskDguWd+fu+Yq36KCOgRGmfanFdHtjYWXONeJlV23BztebJUrijRWj5/qOJVR+RO6ofoTcm6P
7YiQe7821/BdvweYxHm7Pb2L5q27Xy/3A5jZhmODag4k+166gYY/7EDDghRd5ib4vW44T4JYaB+C
knfS07dKto0hHGNkNAEE1he4Mrsn2zljCcGvwuI4U/bXE6/iytJLmt0QRbxUlFAKvv7ysBl8AkuR
fMXLzXfuy4cmo+5+BmlMhox3sUsxnP7Y14LFxplJ6y1BbnOkr1fnq8Xres5sMQwzlFO/kF8kljFs
RGNYZeN5uYFB3xVw81lLNXGMUy4rFxzVcFSyRZi77at/6E5onhw/rk6vj5yWj015wA5o4eU6eUwm
JPVOIfxXfJHZghNgAsQ4RdTDtMnNjtkge6YTRtFe++OhvWxY2avSjd95MNKjcXl+APpDzzUJcN2z
BfSuNo9iCKhXGH+4+xg0yKnp/l7zFPBkzrYGDEJFpwQRGb872Fz7h0wMk+dkUTSu2G3T7cfW/UYL
QIToLXQv5m4+PNsKaQ++Vzelyo4ViAFYUWBv/7H2AnipPuyeJi4jJ223uyIkOzogOvrKhj39Y0f7
LpCmjL0nYKQyMQy5WxS9v32zf0vb6cOKK1mDIfq82gcXPix24dQjxz6h31hD4JiDibE2PO2gJDQB
/kb6PSkcYOLw6UkpdYQ54w9q703RN1KH/cK2rE72x33/wFKfLqF+TvdkYo5QSgcqXmw/PFVKEOMG
PhRIKkQPnaz9b4wTsL08G5q7t6aFJ2khveXCqOW2CMgVXN1HiRa1qRK65IX0BvuutpEDzD6fTXsw
N07+plrTF6nuSRmEhkjEnQlmV45ZsHfOzcxdFBltrMinRkbWKgmWlSPih0ynZSSnG44AfjA5kYNb
Hv5F1ze/R3u4nRz+gk5LiKVjmmF7RN9XXBJ2JSciyHKO/Ck+XXe0jSTN/f56mbCAisWJ2j1k0Tp4
qhHM9/z/EFFbwhMuDhRmtsiek82mWbrRVxcTyD/RIxe6EenjZvVKHbKDiLJL8zegMJZqWnFcOJv3
gW0x2YfZGOBpKlNohyIVYWVdYEsFUF/UdS0oASD8trrGLpPuN0pPqDaw5lPAbKBcAfM7+2nGv8/y
n8vzH4cY38XrbKNLAd9i7u3AHXJ3yxzo2eBD1VkFxBaXEgQPilFKb42TLXgz5fgUrXu8bhtnVMY7
YVYDjUlFXgHUVE9IfxEnDE7DSdH8b9o9wbaZw1rcNI4e75PDrD1ulBAa9h8fL49CAG98Odq/qaLK
+bswsbMIHgc9P5MrRFxYuuHj3GmhNfjE4j4JoXYJi+Hduhb6bX265kwLQ7jhW2GInH4X/WEke/oq
tqzOYGaxi3zk64j6XAk0hLHZFtwgXiq/iOk4U49kL/YDiuesRvYduvgF7QQzuNtafI2zVpENTE76
aH/u63gPFoi1jACZY1lykFK8fxVw0YXLDAIm5SUDfRGgd1lMkRusJDul43y1kvkIvxVmPGsZchaw
brExUU2GTHHnZvg4umy4JwMudjHks4Mfz9IggOmqGGKMVN0kDEePaMdEX/FAjI7/4HpsvbfUJL7B
j/GOa1nwp1tVCbUAd1ziJEgcUmS0kfttoGpsv9mKSoeucbu81PiDUIlinBV3IgeDJsm38Nh2FjIE
vz4Z6rKScGfD5Ju0U5MgXZNz169qtgnMVKPo8VYx47xcq2QZGi+whAt5hyd21LD6OqUEoP7I76Wz
cPEDxBdfMLOQl8sa0b6v0vd3Zknie9MBvSrgk6bPJo9PoYMRxeWrl62ilH3N9Shw1gyF5cnc1lA6
IFogwNCTdP0/Nai7dU5RXtOADyqTAkxrnBvT5WW2S9jG9DgiZVs7IOicJFqjmF1U/MPsjxmiy07T
toymWj4ewK7zKeVmUlCiuFKpPziUGdyVFFRinM/8pC6q5MxqJ98W4vYCyjDxGYkTv7PdsBp/farW
YbRFEFLjuRH85bpOQNUKUV1fAmL9aXFmV+/28I8cNyqIOIPlIMqEuqPNNQX10Mwm1orWZD9mD/Mx
LEw+gFqLbva9TWZJuWRJs1QSY6HWRn+9lFRhVDRG/Em+2JAOK0J+9Jyu7uESTOnvUrptFoVoT3xC
6nxeRk2F6xM+qaE7si1th+4IQKoyhmrFwkG0eSDzxda/ROGg7tL+dff1n9lNrP+GMerR+PZg7lHb
O8IE8usHeTH6Tx8uLGy2Wb454DBpf0zshM3PgSgfBqiF1CxxUPd689PrA0kItc+lC2lOJ/Jcht8+
whjDO2ZzKtlgRmDC0u6G1uKM5QkFHrbuaKGpoVlvUnwuX3vdxGMB/BxJuRM03VZ70qb+PvatgWWh
r+lNPBvcpXBYi+msD/eXgyYhf701w7pjEqIfm9eHDZVMuZmUYrdds0HBij0Tqh6MBQaAChbkpy+v
yrfWVm1DqaWlCRphDRlM4lUc+H4bjPY7Nza1fifs+RuTkVhBsI/ldiVIY5+Uk2Hqvbw7pKZAXp2d
0BSrIjb+lQPz1oDVhsjliUN695AxZT8jfE/ZomCu1ZYYkK7NP58e4jV+T6+at3v+bsdxsFhD4g3q
85vaOAPiQByjVwhFR1TZ+uQzwXHwMuu1BJ9M1ID+Vefaxzvqw7EHw4KaPObFZr0MdyUMCTC149m+
0sSLroTVusYKowCPCWg0MWT3y4X43CFjZaMuoJftRYkQdBkQkyoHLwlByLGDThiAs6dTqDLhGeK8
2bH6WAshkhWY4aH+R1RZ8IxVPWJzbKfNlNLP5E6kPhNImuq00e2xcljUcREYh2cWbO7BpL6dPaAz
ikeiABM6da/2pf+TNmFjN1AakSZ2MgWzUhVyctTRRJFnN/KJFS6NyAxq/rP/+318fnqtb2K4BfJN
CvqjTjSLgQSi05UsHryR09mz56PYp47bg4CfmUJ5N+JCqBeB7Lpb/521xfzqKSUiBmhOUDBmMfXr
DoNb234Nd1gWQmvIo922FuFEJn2il1M1FtY0WRo0Zsu9J2LmhugPyMOjvqukC1LgAySwcKkap+Ny
4T9CzXyis5EucsDWPrjKQtDEZ2ZL5KSFbvXw5w1XV9W4lVzXrZ5CM11ZSKr0i5U0FrbaVStlwiaO
ONt62AjK4tstdpyHn2FcLpG7HlgRFBwBpU1F+Sb8efq7YSSI8sQ92JnC3Nmlm5sVJ0TC/gHVfcnK
7Rr13loAPh91eJHDUneEP1Yft1rukfVOPyYnqhahJ+g+N28rsi9Du6tqMhGWBic/rjg8I7xf+4rM
0wPxi2oZ6rUX0Eq9D7Uh/aqBvVA17rnbvc2n/pR1nl3lTKWnYFI4Uio/dTPCHTV+yCk+5XxdNYv0
IdK9n53NwFbtob7Ovop1JzYQThfcKNyGUnjtOJ4hqwNugcnv3SmNDv4lGFQwInXxGf5ejg8aKLvG
kZy5FdQEX6uk3EdX72M4EhN4Ru8MEYOq+wripoy/q6BUJAXa101FklpPCdjbUJh7OOhAr3hlnjdr
RNMCA7byu6N0QnQhIu6Wh3dHRnLkKLFa/yLKSRbIH7/X3W4wdBrb5dUpyBa/5XgwqHszUl+BIEd9
LsM6xgOKKYtBxBuxSRZmnqwc7l9m6Cjnea/QCdxJWhAtKncNiMaajW2N5xhY1n+JXmXKyDfoq/05
dgTvkkHnI/IwA+lc45Tw5sIwzL/NFbdjR9by+wNzft53g+nUFFA6YWuX1aAryvYejOnSBnUo+jLC
Zc2NYlu/ZgtjWLPVv+g7rFqxx00KHlVuWUNKzx13oBlBs63rzSTUvVPfQnO2fV5DR/DG/X7gZli0
J1g2S3PTPxTVSs6JUeF2pl/B1vLUHqlirh0D01gu1A5HkRkdpY78k9WvlK3E75AOfud2QaxPWDoW
vLx85Fo3B6PsP2os8mnG8UY2Li1i6i+yB4ws3BEOV8vybhDVQDxAuFO4J7aHCKwRjbfxGixQkegO
4m/UBnibmHs/N45a6DOjsrLCK34UKqDFWvhSt+znZ8tFS/lLk5p1RS316SMxFAcelrx7SqJtw1CK
oaev9bcB6nzyByq4AYYRdMeqtNIAETkE480lWEq3XVUrgIAHPVUQyinNOrLAcdNyHpeF2flgVHpt
U2wytLllQ9thMT4tgHC+Ch5XMuQB0jFs2P7m5Wg+dcFpakDWmf1+OPXEuUvviLYSUJF1mhioJovx
5zPUqipYta4z6jSCPuX3p5oEtLGZe2aq/IbKcBOca1glO1wKx9pw09MMrXme3yiwLb8IUBpilTXz
qrl3V5zMmu09RB+VeZ5Cgp8RWkGeOlL3IfkDIU2jeotdqr2ZWK77WlDroWdBky+CNfqKy4mV6kdT
wi5Ci+CaDp1sm4+hf+jGDj7L4D2txv9jt8rQToBJjF7PuLQAUTBLw707XD63/0uj42pIFYmUa6h2
j9Nb5NJv5Z0QkPob3jbwqt6d156u6swE9Ksa3spThInMz4PmQOMKxUXPcExxfBgj8h8SbjMRbr9G
W8x/l69mSmQxIk17NRcmulgDBavpTTo1x3mc9jQeab0bQwTS4aV1e7TrOzvA54NM2JZm/2bFxzYy
L90lbusjg2zxzPqgZlNzzyHKXD0I5QDDJxvrji+6mn6Po3QbopErhBFByvLq1M4E4dGzvy6cj1Xj
4IaG30ql9TVpeThOrqqeyp16A6awB+BCLrPmqDuzPAjkNvG2Xc1zO5lyxctR91pjuGJXRdo2q2vy
jFMuBwFNFK12i2NuJOFnl0LTXzTR8O6sr4z5bI6bb0JRbAbQltrWwFkRrWoqICcF8EdRDcOoxBFS
I67+UY45vXVMzpYGFRLnW1ikwhNspE72Bl3yI4hgMIPtQUOJNvfIkN5QxPj8oGrat9liY5HYXGbw
JDnXNE8Q2Y/LGZriONfs3x0bWtCSw1nEwP6unHjJXqlDfSK8U9eA4jh31N/O/lFbiG0Gz9nbDy/5
ZgPEGBOMMSrUsOBSdyIQNURVBXltTrRBFEEByIZbF/5TMI3DqYOIx01aY8gpYGzfD987EDlmN74a
ZIa7YRFDNXRokQsl3oJ8tTQambm2TCPqWVrvD4hGfkSnGyxB5RbnLXexHB9SwK5Drgg6aOrdHklE
5gLFO7HOOwr3QfOfi3qLWyJQ9ugjppNFanX0QEZrT/0yjIpE9/3lhLzQXKtWlKeddLJUHXvPAsvN
5Sx8dG/BKzdl2ynxFAcCKASMn8xuCkDbwAAGp4q3kz/NzOr7eVF+Ng1M7xhuycDAJtYPnX46MAtX
ACIyU4IXYMbDluqjaW4xKHmKGF7xoxpbTOiWxIhxh3ASNN/8HO8cjl5iHJaXpC66auIRYu8CKQa6
NkGJV0QxEcCxdEezR0HB5wVbx9UcrysMjr31bubEmcFGTp8TcPZGPhe9uc0kcszS+ssgle4uaikT
Psn+OTtvkNX+nTcr+cVidKAOYTH5fM1sJ2PB9ylas0oWkO8s7qWTRndwiqvEjgjUkIluH1Vng4rv
5H9UM0T9/xH5f8eohnW5IUt0SkD/WSMokVjRwAnfr1xxdwAm+HSyYRRyk5A+czixuWW3wpKxezaF
QlFE0jxjCxgnXIZY8aw/QyGaaGBn+U+bGFnffxnLaT9IGp66JvWoV+fnSbfvk/ooKMTA8+lEa/zR
Ev2Ji4uf4W0FBO1q5PN5oIsKKkZUO4QLhkv8H55rBZ5YS7PKfLR7StxEmoabrxptt6yO5HVQzb4N
Jov/n0v5CzyAE/GmAreGt7vgYaltK+YdRHu+B2nBGDsU8wwgS1BHKGS7UMcJer9juL4+9MRR/sd4
Tiau3RkkqT9I5kxWChPpTX+396gwXqk5dPJ/UR7J+eoDQvUUt4H7eNJKfvQ4cUlFSr1Bx7Iy/QK2
pCsskt4PeB4PlGROcxd7tSkeJUhRGPGEhVi7cx2Zy19BNNLb8Y63os/P2qufbf0MHyM0vDt65qHA
XPC1xDuZw9nLMUDIXWz8pK93TjVAYGarg5UdcbFSOhcjpen3elvbOBVHRA1F6N8x6nSUsDxWT214
9Vx66iFwMCHklX191HnRLOMFQ3FlDSj8ZNDNBfnkVPwpjtJkbLmzTUCMWytikmXl0XD+I08/+0cP
QgSLBed55uppR0A8lYpVY0fzCWvg+UTMWlbuXlTZP5OP6UgujKn9m9Y0mQhozYgHSs3LCzsZhPXr
w8v4MOUH4MjfLRcr6Ai9er5xx/15xvWmiro1zjYIB9LkhQmXnSltwj7SmJyrCLyTgta6g0DsrdVJ
h8Hsjvd7C4qYDDG4QII/X2KwE6jhBoJn4GtHIlJN1EJgk0dgG4bU6NzqVuJB1DDzN3kMMapYw9qz
Zshaqluvof3lpW59tIQ5ppDSLXp93/oC3OWdZTL8/ZqLJxyW9P/dnObfuZH+Uyt6HE1Ppz/7+JJK
lJXHm+Zl068HtEkVhzCFGGvF8/RfHpqT4R+mR5bVVa6IxoHzJouiAS1KdbpBSwfuAqr8Uwy2lfXt
mgzOPfjvhvWg9lwxbqjKMX+i8L+46AerdhZcVIa0zXAhhsCl3aOt2L6dbm7X0vJim72e6DnEEVM8
albM4Ei54RvpZiTd+zGqcvdWd81LO4KpZNw033uP2P8BWODxSQcOVW0AH8gKGnRKrhguJBoY2MDq
oZxnKdlaKY4q5uAFAlCgrBuZEgYMCVHOlMY5XqleSKvTgDjB3MJb0aUtLLwd11+4vgVWZAwm6KRi
YNHd6pRrwzY4Eg7aXNoJSTd18mBGlR8rH+ddIHBh22fG4f8qJcj6y6OTt7DhN1f9NFiLZhhvOvh1
FIGwYS10uCekQElYHyqLmjdfG0nU9/TZEFwgNkm6BR9xY6CAS9YK9QWzXvr60Bx+IG/O3cJZzbCq
BxeIiE/Sy+HNnuL95hKdhp3tNrkzCZL7C+wVVKsgA2sIxOPrY0wJD5xYw9kqNEj4lumqAqk92vhR
uMLCt4y+iAZmEoQdRN/uG+oXwJzXgUMfcatwc22BXVoDShAaOTgwm/oW2SMTWfk9NsfkAh/w8fbx
tsuGluoU0n4Hfd/rHWAFoqKxmhodAHojCm2dA6SHA/HQjeBXRNGYZ6BPsPGbEylDHQSF3pLpPVMS
SvL4/cGoS1osEs7erM0poxE3ZPHriFo0xXp5tgX6ie0fZ8fCLk78qK9QlRoCYmhoa7iKEV0WRsbc
+vJUAMBqLQWKZTaaqF9gcGpmJsPBLXBGlUDTYbBu+AhaX3uLuskaSH4ARgK6TlTN4/FHM8Ksmivp
cygZsKb+v5m7NuctIjophr3vF0dETu3wLfnAMF3NUJ99k1JJNuEqWacyhGRgw+FWs8CxYRwr7uJc
/FlMnZH9SuUA3Kzw2L9Zp/Tww/XUw5BDhshiE0QRUfR+oP6jeXiIvuD5y6AgBkac4oqJd44oTI3O
XU1NbBRrwzj/4vPDJnE07NjpLkpRiY90ns0Xh0MZgZv1FeWQOTNj8oi67Vz4ZwzJkaDHFyC1lrxt
8MSa1c1nfsdyW3Fpv9Tx3WWLEHOXAGsV6H/oU6agHKVRHf4cLwg711YAEaAu0C6X1g11KtE+VZbg
BrPy5ocHnFvz0W0uOyHszjwJccaxuTfdk2URJpHBbfnlCj7G3Itapj932SKi4OdIuq81oG2mz8mu
kKS+kuZsDjcruK206anvWb3B23HEvLwjtppREq9HJIDt9r4QU9g9VoJM5PNuOqMbmaeac2K3FNWl
nRp5jGK9BJ/CLGUHpg1wY4Qy9C/c+VsfYnqFKDUQggEW78ox6EY0TetTRlhQs/zBigJRhxVOlRaV
bjQlHaQMSYstiiUZwMsbdn3XpJg2q73gB35W54YxD3owHvvqa3g9Nmeu1ta/7Ko0dGgr6EpSw49P
fKK/073eb4EE+nFD7rgZYvZMvgmxfTpcuo7yZ8Be/VP7c/hEZplJ6WDrWTFq89u7ifkpFzAlpaSE
mkclscsRdkEW/39N8+O799vxWHdnDhWlMNoZuARo35/k1UbF5p12gJvLLWr/0S/T6XE3TXDQ9D3X
KvUoTvxCJN2M9OlbBSmIvyu8lZyO0u37f8MUdix3zoX383LMmXFmyfUTCl3/m4bwgN3KQcoQU74b
q1fnjngOuRwkKYjhNymL2oHhJWjHzobzNjNU5b24xl4Aq5AU+Pv+/1sFXar3sx4tU5Be8Qlz/d6Y
kIPRrBtHhJ5DecQebU/+dz0aYnLXuq36bYibcfe1gBEJRQizFEw06GYImEg3KnP8FDkLiqkS+y5n
j6GRVOxbqIWhAMamlMulUzyTO6yP1lyid2SeqAf5mAgNSVnV0zjRT3c3dQsSDpw5PYR1TOdNbCE3
TTHjzSlZWmCoLSPu2b7SMMH9qk1vPBVO0LiZDc9peHIjGIePu3GK6nZcnxgHIhPnoOtMaGHjoqfT
wexwhtiOIEUUd3tgZz2YBkykp1qM9iUzyqVpkDxDzSRQCZzDnIuwjcKHdaXhU+fAWEFOVjJlGFbd
yyB6IZjlqpIJBvstzzsTvO12+jtyy1Cce1LcOU6qe/VVHLatGa11LQGqKiwm2+iU7AHPzorp4hiQ
16ZfcaXrWPVB303FmYqJceWUns6NlI6rKWJH6UbDA2KSa+jbunw6pXeXGq2TO3Cx9hu4Y/JwhWtp
pnLC5r6Ebjk5O5WP6oxYtw4DkE2tRXf8Rw6pVKLTb7zXfjFhZQhxtS/nRjCGHbnP6M2z6Hozqnls
dbnhGsqlkdfKY28StUNjBuxdQlLtTrTBfCG0b+f2JsUczET8GEbsIVPHz/3WC5Oc7LiVnQAr4G1o
oxlpRRN0+RqZjXUd/955YsoGs6vP43fCPgChWCr4GzUCfW5xoBice4WaEamtdtZg36hVRX/SdUTA
1pOd6wT5jgUtL3DaSslXiABkJZoD31kmMxRIZXjbCHzs741x1KANtQV3yFJ1v6HT5Bts+XITIsMV
72SbmFsjOAu9mm8kgPvMw9URFEAWy1y3iX4g/k9IXj9HaQqXOP/HFL/EAb44tkbweSqAsH525Vll
3MeOxsrwNgSYkPpzMBaTqPlmtJnzMZ89qGyLvivkulWBT2+JDeb4b/COojVYknnkyvCBqn6DUArl
8UmyzL+KoD0h2C4+ziu/+nN6jaJi1skd5pzNiUo3NoiaYlPlVf9E+E2UiH+Oboqfw6ppiG3+6I2T
xiqR9YBL1Vww/jchfG98WnH2LQzQoYji3ZQq0H62NjjxQL5USyMhhUuzjOgzUHhHnhezyxH73ITP
bgM1ufhLL/7ouFYkDhkhv9YV/7wQ/Nyou+AaT3GlK+5bTPFx9kdgO3ODuIi7/4+NHyIuUVPRpI1N
94KqP7BRUF/HMiw18b86M+AnBq6dh6h5obp9AKG2B5NHsvrXITUm1gvvqufG6YWqRLJ0m32ZuTu/
YwdP1snFREft0ETAd9WQbc47QdnUjhsigyt0a3acTEna5hVSYsBRDe/0maf+NSx7YZ6sq+Aal9A6
iOynLIcDF5abc8hhpw2rJJOH7/3vpYqUroGlcVmM8BD8qp4g8ZlfG9vH/+Aq/iUvrSZyGSGVztt8
nGGfIZ6O5yAik30O0WSNUu4eKJQ6UiMThS7m/Mz4CK5tksiCqbdrg64KuXDKxQvXkpOhNzdtFKAd
jEPwIXBEBE/cR3xstw5EGofF81YZZD7KbF3HS61Ctsj8Soow4Y70/DM9eu+kbQx5iSpDrjXT2E0k
8YcjqP04J4zmtYQ/VPlhataMLZy0TeYAyuececa8pRoeRz2tBgd3sMIonSRK2U92KPzN4o/SOcre
aoFbEVKnM8hRV72BNhxHMxP0ZtwLuztzIBqYQIDGm5pLUiIVFCqF/eeWnPsytyoo/mvao42KDCeZ
5BQXK5aoXKMcN23jPGMiH4cKVEyQHlDDcQoRpu62nznXMcEmJy61yILg+w61h1yw86dlu6jcrJTk
/4/swTPJEI5rMXbcRdU23H8MK4iJu9gmJmU1a729un3I0fB9guKIjsGxRkay05r34qZ4fhrbFeR3
9bLd9MfFYCc9CL/FGh92igLseFtM4yU2RqsMdbXUQL+GF53WIWJNL4UWiW+wXA3clq2rYwJn9WBR
dOxMLdRUYDpxCkw8/F5EAh8DgLBiU8XF6qRt8qLKdqzHIPgSGVE5dsgrgzJCtWVDKWf1Ll/v8lJq
YV9coKKPprZ8Fx7Jhq2mIfOlQzwz+W4gohymtpsU5xicaVvdmW53TjTQRGynOslHWE9+wyoxsop2
UJtG1u5Uf5pz04q473xSI7iaDhqA71mc7YvoLhF+HDbMAi1BTAj0ReJadRprSkXfg1IGPVMfuS8u
qO9krcjLIB9KnnZengFjhaaLu3/T8aie3FWWeU/mbTUGra0TkOC6nhPbb8xa1ZG9Ls1ihQrSZlhc
8vYyHaV3nymBlUxJvO5m2FQLuwgEBnFA9wK+K6sO966KvX7393XjmkYUHsmCsifhhL06BQJyhq4J
b8jK+QsbbEJVExwPwgaUX2nnMWtFv5EQrdYbjfJsbVV1AxjOd7/3aK73wAS5J8XjSu9qN9KwD067
38t3aCGSSpBEhDE41OwgD1MuP5UBEVYPdm2WG3RiNmuoFImaMpgbpsmhUsM/4Q58JiVYd/0iXsKH
9zZWcM+lMVt8al2wJA63SfZxUnpc723jPg/hOFaqwqe2whRS343ynvEHeEhgrVOt3YRTOWrKod5J
SK7LVATK5LcOq6BEASorRSAAlDTzbDhO7NojlsEZ2lsBgMpAdON39/51peJzema7XEpJN0Wyf/8Y
FCYGctyz+G+NnbmHGYjwBfTqeA5RoIDGE4GyKDXAEUv9CaBX3qX+07U5lY+0AIUiWTX8UiH78Db5
iwM/mcKlSAeYqMdYkk47TkIemOJPMTl0//RSvRlp2R9zJaM1abPZwcpuIvcuNNDM2vcL/JStfgOG
1JrPqzc1TliixYXfkx7drnMHxjDeGBTc5LGnasoQdeoFDf/szr24p250ztfu3WlT8i6byJJIi+MT
ksQPFroug5PEOaAt6jwX42gmSGtxUG8NTj+JssYs5why3HOHYs9g+zYslFbY6hIQE/lfIPc30TkC
BVVbB2QdioQgAK+TPbaUtYXe/DhsF2kBloRvKiBWjut+fPHbXwwtIaDxxOH/v0dMn3Jw+kI/s5nw
M/r8pZ8/j33FuF1htsYZaiwGVDcl4wVg/JOUGgYz6q6E0tTdwi/QNqPVUKmYUcti+ymjZtlgAOiT
Q4DbSkwC59x1CsgAiOnREp/sKdPL8Ioh2Z+ZQfPi/vPZVGzeD9Mb9U6+1GGAgc8Q1vVi0z5GqOjn
JhQvfKiv7P7nRRVVGdpSjBKUejLAE1RjY8k3cJqe9Nx9mg7VpwkA7FjUwRFq0Wt+mjGCOiUaOcZR
0eOmHWoys15GiISg/+Ah+hKBOTa9wicik9+/eW9sWJ2PcuHs7kzE0DdxouxbRJiu8n1sL7entVyB
z607+ySXNXm/D/auOfKJB6cHB7JFPeI0gctNAbRIaZ0fAPBm+miKz9Vsa+KI/kXkMekVHnJnRLqm
m9zczYex357PjoHWO7nj5UyDMOZjDTCaWt2m1/KDmb4laNHK1+r49KCDGV/ko7T6GQz8GrsoDH9S
RYI+xapQepRNz0fDIRSoYrFrO2ZY/l3b1vn6uhZP7AISkZFTe2A1LLXCtrryysUyUwbKe2yZuWFk
4jxC5J3+2fREJ4zJJnfY7qxIid9Rq4Eig3BPXyOxZtPO56jWqN74Q6xDMw+u5gNU1ZmCzVBn9UHy
xT2tgLS549DPGtkc2oMUOIiruM9CLAVZnimlT1AuRUDusHMzIKZ2wfDy065/Y+z5Cp+DXK8s8/d9
iGYsdpNjj4BqcH5sGlDPFODUaKkefAXxxZ8NNyBOt64/q66LkZvHoYFNXgFoOzVcF1peH06oHAAw
Iqdb842SIZJjPPj8PJ49Xviw4DbViHv33MExYWpLDOCvjEP36MZKg1GyoMMYmye/Mq2rxzeZ8d0B
/UpxAYqN35OzvxtaBJ0vU8hble83mX21SyfBPb4ckTIS0Bmt+Pn8gVJIp8k73kR7/YzhTfiUSHYf
3meUsThdKq3sOYDvO8zpOfAP+PVekzLudotVJTzVt1aOGPcZUBQWg0Eyh2g8ii2FiWCYA0yZ5+J8
Mzfx4V4OZNZZ8G+3ypY34kUM9KNxXN+JHSijFiXHtzqMAQUfn1G9dO1QquQ55tmexNttkX4ghwtl
MVp9pgZQflRXMVkmZpEMiyMKjyYjwnt0ypbs1y1C3nuIb2SUsZBb64UTnUHfdfR/Eh+J6mtOAxRC
mtG2fXTCq0c8nhgMx4AeEmZAQZSdYcQiG91BNITNrr3U0vQmPEeB/tbd5YvT7KpCRQlXKdiKqA8b
RbrzoBnONFhL7KxHhl08tR7wCDdqp2ffE24hhHyHD3zZ66T6gWipWUlGuoZMhYrJhI+yo0ft7GaB
DaLjMxnvzv9jp2ovizxGIhzeclDBs96Uzozu0hT0cSj1NGWiKGI/fFZp8swsvL0L39zql06MIn9j
9cj4msT0pFBKD9FAIIORqcZeCWbesAbOlgMoxXMEOEFvqXYE0nOxvUY3YuoAZD7GG9wSlqJpVf0v
V+H86RLDsuHUTyfZUhdP3dCo93mB1+JGmXthQWHxhNroM93g/9KWKtnvdgedhqstCpwG10SH9roH
ZrIxTIqKBcgaFiiImt0ULisztY2vpCw+FEBfSz6t7BOXoh+XI1UTMw/MRXDyyCg/Sjdmp/nin/U7
2j3UdU1ZC2qPm2n0JwTDVHTQelMRPhPWslujj9FAGcAjmSzFQK1JCWKClnbLGSM2yLwW1Ak26/8Z
29hIVL+wirTyBpUh8/XemsIkhbDcOG2wBmXe2nVc/E3dYh9aCaVKxDtkRFkRi7wCF/2i5+B3ZfZw
WqjxlLuLqXvrguLwGL/+9f/u4kMMhPrfrX6Mz0rh3Qz6/R099tUhYmqrxV9r3AYpelciEUVRFrRH
bPYVDajtxq60c5H0WJfviQG2DcMaQ7wPkQz/RVUH26W4HRHSSc+yFvQdFDZxtsczCsh9rTqyEsf8
idfVJ5gcQEptvLGAKoWI4HIypbBOxphHKzcxlPSYPXTZbd2x77teVU5AeldJqUHU2Jk4juYi29ML
PG2cWjdAL4Jkv1EJPEZq6UZtiGTk97x6mGbIz1Z+/5TJFBH6cGdjzyRMnH3vRN7B55Zl53vPajOY
Tuy9rmpBexItnmmWoR8g/VkREoiXLTawD0Icy6/9z/piiYlG9zqwi3iOcgEA3PDu6d9W7BEf2GU3
q5LafMGl4Xrq5gypmQOzYuGx97yg5acIjgU2joDHxfjv9VeQag7tgrW97/vgXEUzmJTuQrjTO33r
By9ipSvYGIY2j1GOoVSXRAZV+5L+Lh+QAOZ58ZL5Sovd2IGLlF1olDXibjMa9sAmexWzy8SBzKqT
Pbm25MgNltmLGv/Hh2TNwGOsVXLf89kW6a+mjQRrxLF5AMwC6Kgke5wsW6a99WOwdzmVuKVtRbd/
ElsqM7/Dwk/RIXD0+Hr+OEFlEfGgnyf3h+dbLV24G6tOdecnio0r3rM8DxAZT8et+CktsLmXQYsh
AnhQrFJVIYgt6lmvmfAF+4N1K3TolMCxgQd/pRePEfAKpvmJJwLOXqJCWu43Z9WxAurrEtH6+LIy
/jc5K8xaBemNPaGuzacD1l7ZkFct7Op32nC9PaEPHqIsF0c8ZzIVUyz2MFxxxD2Ae5HoQMfjQAwr
pTiCLaXWnvsDlDDL2ZqJfA0o8Jtvkd43vDv/1cngskXq0v6FeSo1t+jRGAPCiOsD0lvgDu1IFEer
n45/DSr/iu7cXwbWrZrrK2vMgOVcO10hJUTy50gn+5pOpXkSFCm4jp8aV5jOIulXwx5N0BkDX+NJ
b/YvD3aKncVwTBmSJnoQKt/CmxLA5CyDm8Yi6B/EE4XpIVGt6OY7VloZV8cArOhwoZOEg+1qWXn/
H3xjA1j8vN2xGEVx/WPo67cluuL/m8OQXXl+jp4r7klnhFHevsK2QKyObggNui0Fu0wZvrafT59O
0D22QPDXZKua4DWM4IPOOcGzJunuy/g39VAmcl+qRaGkNu+77QggA5vMehSJe0M/EpqZdPzlzjDl
7FwyJmfhNJBjVze1Hl9Mck6otkApTfCHbKfuhxJg5HIePbQlllEdfR1PjLVjPYEkOYtIgY9kDTGV
+K2rDisVeqqGf4L3b6PfnOs+UXvhaQys8tJIW4p9DYZhL4CnBOngnL+q1nYRNbWPQ3CtcMuUL2qd
zicy46MSNxzadzRtaklwYwf5Bg9fpKXWPt+6pQy/+Vp+eEWUpMoTbvJzHmyMqD582OY6YVOGBHtO
L92Hx5alRgwijrTV54I8GA3OKUyhJLlbYOVFxVKDH7FhcRL7vCnfXR8m3WeOUW3/wqmPm3F/TIU/
xhc0lx7iONQB8fHSOcEyCw4oPiy7kHCh95L4mUDrEXlLFvGfnUW87XM3p0J6c8t1olrvcG9kxBys
353ScKr83Soepf8Mmdx0v5kZRBIPm3iPxO+Fb68LVrJGkQykJjKaELV670sI7yk0sf6yzhBJhAxn
2hwllQnoJVuBtoyr+4jMZsje2j78MkxslklxuZz32/5HU9B0JRlcl00aftMaQDNDUaUcRolFHms3
LoSbH4J61a13MWID9uI7Dc6AoYdStvjgqYoAWDW84i2cDrUly79LnI11KsQ+ZnjSHptcphhm4QZh
t6TOOiCvM36sjnflIu0C2nD9iaYl5YRh7t23YKmEuGWTLspApzZU0KvZf2335zxzPwEyntEP967v
6zQDx/e3yfLkEvAIzVDgkfv+3vs8AsqlwYzsAlKqdFyFI/agOPYLOmVzWsqtMBbwV+x3ehM3xh6P
Kw8YF0mtZDkEXz3JzszzLM0KEErkq0Svgfq/9FkOtlIwpUNCzdWi+G+MJZTIFzHxEZ9sOimiEKIZ
Bc4jmlLRxyzbjsVpLlyVR/GW4B34iYmaaEyhJWYUAsdecdbxl9xM2f+zV5kfc0xLo1zxJQLvNmlN
NlgHvagoUC3DKEMV7FXEYo6/YI7nbFZE/huM13Dm5bRGBE8/CzJ7eSv4TwxEsam+ZxlFdsGkYA1v
OphBWjGOk763uVLKrIx+aa0ebZzFeTGhqpZmL3CXW3BWg9WLJFc1d5Jd2FiNyuo+Pj8ZVpJR9HeP
kK3XEDGkfVXawHaMm6BSLcNm5dcPK3HB/uOolonlX7Yj/5CZKhLAfkmWQ0j6rggkKebwIQz/nIoc
Dz5glHYcPFM79JtJRQhzMNTBtWmUYDfvOkUAOiPjpRC4NuOVC6f8JQJkHfZge/gJJDcAhdSp0v9H
j9BSH5M0NZWsQLHO7Gp5fOO+9JSzz2gffTkwinZDMVYvta15ceN23DmMn+Lba3LW8Omw1BSpbVNI
CXhsWHqKz/PYsyTKGnk8w43WABSmFrTEM1PDQuUpi9PLfKtX54GJjWdA/J2MTIRGA12aiuMVMCPs
5/DnCI4pYUqlC2i2gEFgS5aGXEUqDnHbbH+bUoLtnRRKfKAYQf3bYPkoqkfXm2bgFCPlr0JQJCk7
JsFAR0hXMNBXBYxGHvIW0ew3UZzBFMkE27EIiq7EB472Ur55PFs+rA27HHOyhyjsN5k6lWQzWDwC
eOz6H95Gzip1+9HowLDKjO4C3ATSr5l2rCeD7y8pn7iWcLS3+4qfn9dSCZVaBvdsuJ4Tekg+Izi5
WlpvxMkiMJQocP+GkhYMrXPrBy49i2Mmd/Y5ehp9ZwkhgtSaqDgaZSo1/hRD6+mkngjKCNoFQEBA
5R7UzQaHc46nr5DGyezZAO4ivWUeQlhc4iidLMBDx/kdWIMHlZfvd5Eh9d4pk496Vr/8nY6l5NDd
CNCeqp4KXe989//HOmZ9h2uWOllXdWcsiD0Z/YVsHr0WzjU+dtuX1+srVp24PcFx5ccmY/5ialIL
jiurlsC3ytRzFsy27qZ9eMjj7LWYyoEY1N3jcwZ/LrGQxCfhQZSDtsKWNqdArx0GrZohnB0Eu8M9
lfcbxz/TIBNV6wfMOwEqSn/S8ciuXAiH7n7PGC638oWH5aG8BhIXtjxZwVlQ9AwyHiwu2ZWW3l/l
jcD5zi0/U05q6cgpgRoBcDkkNDR3DXzL8mAsaFlu+O7wrXYzKZPU08wMQnRcm+rVihe9OdoR3Y8r
G1Lzp0oeHT01TjobHUq2pquQPXIRAjW9tfhx0Uq2CfxSbfJjEJjUGrqOCgGpJpUY8LWzEMvPT4zZ
yBtRzSv/iYpuz6g3THlP06GkS9KOhUb1MoL52yTNVVk5vcM1whfT0auaRhxFTisQHBx/A29bYKFy
MOy7jWklF/Z/iPKhWrVHVk8DCoeKZ1LuYUDIZRkUdIZqFxDqLzafpUjEglhjp4/ZFanq6oDpy18V
iRFU+z/sJ/K4nsqkjjRYoVVxg+rrUK4wKjUzcbXM+Uu1T21AN7BY7Q96Ke2cQAbBZW0HcAc27CIT
sgX9R6EqS+NDZ7KfbPOGqp6XCH9HeNQqqGzo8v6lFHlHviu93+IQZybjqS33KrTHu72A360pgh+q
wvljhz8aGXjeiRzKSRZ1Z+uTAmVamwnurgMCaOCeBl1sJBUblb8l/Mbz3u+LkrDgtd2UpjXxzrn3
/D6zgTa1BrgRm4//zLO22LD1mHhdm1yXHruFW2DMaXYLnM9kSemzVxdGj726rzymYQZ+LF5hfb0J
fdCAlm7uqiGLhsPRvYCdy2qLf2I6UDtdB30guRwC+0f4JdX3oUW9lqFWhb00VrI5mTTzA2XImh9z
aeNsOlSvGXIgi4lMf1WRb/ALGFwh60lzWTWtKCL/vZJ5q6cakOqPIFJLzDl40Gy/sMRXhY8E2t7r
zxuJvpfWk6EQl5kxLbEbIDA1z2L4PzM5lG67EWV1xLD+phvebgEyUCYxZU0KzaAEq34M6CIoBLY9
BE5hx/CMAHGbCaMmXYRn/jwexNs+0t+HlKSHCGZKXEiYuffjwVkIwChK+ZJ43r2+vZEwaAypA8/J
Av5LQHO+CjuMJa9oxMWestLqwhGpzrXMzIQ/a4yWk+sQlKvwJ+jwNzU2E5wGKTPPqPnOkiRvTFre
zFXcztrJQaC/kfpPlxqnchrdOnaSM0672lV12g3TD06KcTErng7SzZve9wcQNwqWywK2gRmuVJkN
lWJK4vUCwrDKGFMxpfW1mVb09bwTt+UZIdptJPX2rEnhj51Id/MgAO9p2OGKPQpFAD+vPYDt3cOD
FTVgyPEENJGfyoLAv48+siqwuBDerxSpvGGbITXQyZ5x7SdXsxldVAnLDGc8gpwmBnPZzOwbiJld
AKvZ0h9u9/DhaEIKGESdy5G6f8LdK+QlOOLtJMaRJzAHllsvqcMInz5kST3poxMUEiKzFsFuecaf
iiUb7K9evuYQ3FmxdSJOomgme8pgjYduDNkT8hbx4IgIvllqa/VVYkaLTRsHMjSOuI7GtzZuaNM7
eoZMOhQuhlZSF9wDKLH90/nyU1iydshdvroN+ISgt20Xhz5NmhM2CzXz6+nPdE41NawhoDlvbHDO
ELH6fUd2piGKjRjS5BUXoOmFb0mY9pKA/5y2C/MV8YiwLdC8z+tk1w3EiYxfLqyq+GknSeJOzgNS
jcL3a7B5CRuMzEhBbd1lbfvFKLlIDkq9NdTGrpuNy98a4yqyc/m8YJgA+lAIGjr550i2bfQ/3uPa
fJJ2TGhh3fj11qyo7dD1GSlu9C11ckS7wfyXII2DgsD7GpSZyIIhS9CZYISCoQART+MU+O0q3O1C
bL0O4lK2VEo7bIFCIKCFwd1dn7KV4wSterHJtSFbUgt7fljJrv8DblFCDv+EAcgIY87DErXhCQWy
r/Gx2uz9BdDaH5VLk5Cllxdc0PL3ky8xPqWgTeHw0GDm/Bf4dj8vgj5bDG0oEaC+R5qnwOC01rA2
MBMbKRIOt57WeR3VSM5w6VpmFHzNiwesu+xkFFEndyUVbdPf1kDkYtU4Bdaj/3e8Vp4/Hi7ipFsU
OWdHqyaC4Fuw1rsCeOAAc5hBNioVfc2hIaBNCMh20bAv1H2OBtvv2pW5Fy3btWaNHRaWpbaP+zpr
bO4UD7ePpWqd9/3hNd2naDNC7WD3It5UknrIx1jcKHKxvA5mpSw+W4SE6aZGewaJDaeroZKK6FpA
UitY+c/neGkaYs09AjrbsUT4hsiOqgIk1lx6pwx1qCzqsu5qG5D9iaFuXpzpG2dXs1CdxbLAWj4Z
PwGGFDWbgoRWiADS5Do5AMkX+uZIXV3Ats/ZukG/zfvm/b531Bz7nxrr89KJip4d6cqRrW4BxUqD
3KnK/+oEETsN7ds7P+n5ajV+zC6sBIRk1yJ037SXAA0jqSfZizvVRkq8QcquE1RF89dWKE8/ga7o
hvYq6ffkV8/HHA4k6MRwXOZOizkAcwH6dBGW+AMmi1v4uI6oCTXcmDiISQowNoWUdzYT9qcGRVLD
zJ1tnqHh9v4Acw+YJXweb2vdgov+jKFEFQ+wOa3sjrtTt8nsLdAmV1xOWheFb2Jo+DTSeNHiYbG/
IB1CQ2VB6CHOdAxjng+xnlB1bmqt2PdO91aMAn6FzaJ1UnmYrvWnFZF4w7QXrxqUTRm1pSztpmmv
y80bzuKAJP67vLZ13A3QQaL+uyBywUS0vNP1/A920J/YXl9fj3bVgCYnwfhCa+6R71bODf3oToBq
7MxsWk0b2Q6u/d03dLPJ3A+CpE//9opTl/wBMH44P5k2AELmBzDReDjzRGVL0iAV45xxZta74UoU
hwvZsvnvcLASEHksGmgbc0OBXADMnTdX9CWBHxGghBycAE/xxhkazh/lpHoV8XzZYiTfCq24JCGm
3lJ7PPHxjtY/5q3xRuXAdjU72MFXkuLJhG/Demmb35W9StJtdFXukR+zBUWF7FI6CBZ9vTGJ35l/
iuXtuQPxWCbqXwhXCvhavjeoTfCgBM75gmpW6kEw1/oyOSADieuYEDmUGj2pnzTpblnP7cisbu+O
UTLRmo8tNf2CRBsC0eCzoKQ0sBSNJwp8LjU+Ns6ND7YtoGTfn59URtqPEx3b69V7lCspQDcL7BPM
0LUgL/8CWdHthab3JXTGDW1ovg4+BB4U/NZ5r+KVptn+8XkJClJQAVFdFAXVqghPniiEkqDRk8OA
oTc5tV4vs5dHUgFSzUGv2HGu/U3igMyy2HJCgaVl+SLxFdbKS4BA7ySJPwchssJcZIuuXIZxgqMb
CihA0GI1sQiForckkgjL2jeh384qMRwtd6imeev/hSHLCBqbBI/XHpuBtltdyYJFYz7PtHWVQRBU
YcqXTTwzjc9yvrkKMyOZHsggPF6A0TwzAO2g2F2cTjU5zXQbW11uxlgSw82w/wJeQdg1chlY8qBX
hzJ0yZXHn+CCUvJYCMFBEeis0so09U9H90gJ9joIzJiKlWX3RoPCgNiVaQ80OPjyJSQxWY8SWPMT
kB0gx+0vOZphcLw1qfszYenmQYP7C5JeeIJgcyjTnOgYphKULa79oZDL90rHhsKGRydGqOcXv8lw
UA+x3iM9qc7POa4YHc8qiYd3c5up+/4YzoHzcVzBsV0JQw5Yqfu5HuIEACr2+ZTtTz3o4zTr5bJz
T+lKHTwEHXuzStxvRfqCC+p0F1T0arwv0U/ovYORv3gY5t2M/e97gz6P32Z80tYGpim6ipQRxaVp
QhfPWykRJPtWz6hBZzX2E1BjcY2c4XTDnL6GAPjww4wYicLPBP6MLNCeYmeQSpXIzI7GSY8i5Zj2
bfaVtTgTWoNN2/etMpnANyzayqFWuWZ3taC4f3zLEweD3su0OX1ihWLY7D4HerPEO0uxzrTOscpl
4zrvwJUdcQ0xA9EGZsnEsBPfrtk9zEZrVJIlTMVwc4BFnJCfNiSCs9LMxnRALI557+QZJi1tl46a
jQqIByCbfBc/ZFHEBsER5JZyHC+o/l/kjS89oVFk95ri4SJYX9wYXGhRGb+jovcslrt/W1M7nPum
raqYT7CW5gPAczMM1QH+VadvxHGRw6pnKBEvyTQeeoaXPhUsXikYD6IpDfAgtNlR7uO3JVfRbFLb
hYjwH+lUN657o/lzfAwM+N57tEgIQ7+IIhrpioa971urvIqV8HR9CJzmqh3tQY294Ik2dLuBChky
UKJ/K5EAVmFoJx/knH7Uq28wsN0uqtvVPzJfcnaIoGXHjHhaMwYJqfBbuoL0J+e+TwRbtISbtM/I
mt1L+yQRjF+GdY2CP74YQD7/vVehifJZ3unpOYGIDALUJV8UePAo8rQcIqXOiGmsdO9S5hLS6Qln
jSgrKYTb45eh+G4yuJdrNZr8PS9dba/QYpmhaxju7SLaXRWB8YaBZVGpalXBMvgqy/k+rBjTOPrE
le+UpbjQb8eoDN21dWumFCxgoOsM0JgFjDrHnkyMNrPzEYl3oiZN+dMiBF2Gw2PJMOIlNRNWzM9E
enQCI3O+SmjuVWA0hf18XTXZKmOf3smRmzwqXrmEgJaiGh7zX9uQrFVgay0VYZx2Fd7Y9fVLlZ7D
LGQDIeBSg2Mhk2PgxA4dvVvp+b0lHGmv5UztkO4vc/LQNmcV8CmX9C/sO9Jeds9Wl0P7tnmmaT9U
cBR69ttebO3ebvCM0Kl+g2sHYU5xyUoknpVTFQSy+lu1OCYCAzpBjgD9/LO8t6RXy9nNpDWX/Deb
qTGUqWxqJVa/AdMJL5jiaYISsKQLhzy/aj3moJ43Y9ZefGacjJkclQp6hIgiYx5jExBw79GbSZ41
E1zDebVTN9ZcDOppsC4Hfm+hIDl/g41qmAxIeyb/5WikpdwwxLiPBBNLn63apwAbRgyY5/ZDpwTF
r1eMNlO7F6dhAXSpPnNNggEVMJKkDek6a81W6IuA7PhFe+oDcSlPMIjDlCWfhHF6SfYTGUpiOhs0
lw1NnS8BhqCj7oh9JUmHpImz/AQSht4c+EIcfeHvwtHsE0o2FQNP6uBLJaMRhhqlOCORceJj2hlq
bZ0K8vV7rhQ/AkEE6DTCzfmtScttl5pCesdngyLoKkxZTkWp4fC929QrMf0nlvjXLzHSwAWI+QHP
udD/Uwi0eL637NCabIq6+cnOsfpX0IYoAGOXpEuyTk2Ly1mTskOM6r3lbqAfziemprQCFM52P7or
umF4MJzK+6ZaEBxKnkcnr9fGBI8du1CWothnzaBiMpDfyDC6uVy/a/V6znJBdQx8DHgPjx6e302G
oSwNG+yYK0LDGnpwe1MoRDdwnxXls1FLFztRwaMvgrc9O1J8FPfaQ3qERMiiENA9c4AGr+2+pb3a
6GCxVGQUysi+e2ZUf12MEpRvjY8t22XvnBVCYZuOTQEMAgcBcDxXIYURAzLEdFV4tLS5fz1AxL9q
P+5zFTO/200wsyS8EtXl+mYRcV9l20KomrzTQCIrAiXExb7IAQRMDhta65MQDP34njCv0kBn8gd1
X1V2U0b6caF079uCCmqaQMIHhfauor7tMQMQ+gvmlDi3E/hlFXlMM5kZn3n6fJdzS4VZJpoYAT1Y
nLfzgn7zO0494kZ7Dd0euvx1oR7oSX9OCu0oHp+l/Bp2uOPyjVLeFNIeSObQHrfwhEzefNVpR12d
d6kVvkxr23LRO0yH07Ho7m24HRcIu9HJWl8q2vlkVw5NXYILrIzLirxHRm6ObxyxVQiXjMngGXxH
dHh7bb/IodWnacEa1U7SMhO39Df+FbymBWzX5J4OE186ViBjqvRzSAvLYyHP8D90n4AXYXc/+y4P
+wRRFPV1OFDvQDEwakOFF+d8x7fDlaMy2JVx6i/2SC9+h0X0eeC95xHgbfzVN3qXt15ffrRNWpk/
d6w/+NbURAeHSMPU1/2l2hXCHuZQ5iYenqbXh1qpjqvuZfg+Hc7lGcEu/WgcoVDAcXt90HdvY1tm
Q7S4X+cYeeukTlu0pJ8RBmq37NXd+6bkO4ReSZQTMKPHdgIlHIYg13VTktdHZWK4NIIwH42QP16D
ZAcSjX6fLvl4hwIpMjnLRyYg7ZOsWAce6Ktb36Ws5HJ9Jjhr1cSwE0z5TPq5gbnCPXwwq+kSv07Z
ksaDd2uNwCqM1GoN256x8I1bzfra1a2UWwB2gqtpEPsU3YgmeCrXuMGmXPLnr34gz9/Eqji4vUNh
rg+fE4Thd9cZW1xwGkPW+LpTKHZXFTncvUfYrEH6Xnzo1+ONTYjqJ3KmAxzUg6Fez3k4sgWv5E9n
HhmJRCZi6lhLTMuxYAC3FjggKDr7yP10YXWOo0P6eEQhfcuw1LXiMI02IFS4RHFio2dDw9n+GZ4q
UC6ES2i2CWBBC/plz0nElzDsRByni1Bi2MzXzbbEBAKOF2RkZzEeFTdzaeIoKLlUROYlk/N/inuh
VZykMkQvvMAKRvTyUie9OCsB7xanXu9AA46KQCWDom6CRspQdb8Gp+tNmm3cIVVm1QY1SJ85eVce
9vy8OQp2UOEPar9Oolut4e/LE3atyZFKwNZXirpWC6OWQAmgaKDKoUSnheIfIQyORi29k43CjY4l
cBfRhnKdZ+vOEhTOmcYHnQRQcnwZYv3NUc4wr/CMfTNA24V9UpaNVJqIRJVNJ/heCOtWk5TeD9sF
vlvg07U9iwy/tfzrn8UkkUtkSZ5TROuhL2Fg5yBzEiE8dDCniON3h5AN7J2DJp/d55+tjj+OLgcy
GgapMSWA7V8lwyzQUCg2XdWFax9cZqFMxzQCNNHGgMhQwXxYzv+L3blfdcQq5Q/LE+4v0px3bH4g
xkaiZBW/pqsHzombfE7pr80VutZZhG6PyblAFjX3LhpZiYa22C58rW5Rqy2au4/esLpUrcdVfRIa
uGg8YEr/K1U0xf10Vdv+20263ndL5yEFkD6WZySUg/iAxX4dPVz1mc+rusN6Wf++3+pB/Z3z0G+j
gBqj+xpjQ135OoYve6UVulJc7mbuZkU7+CxV1T2+7MQRMO8E3RJa+XvfD9m3fj9ogJr9T0R866cS
8I+JimKOOydOVaK+WmdFOkjwkGpEh7i03xjSNi5KWcqnWsqbjCj6N6f2Go4GhwkhFePwBGME2/QK
skWONKXGo+2f/tjVLj5jwcUL9xKA75vlDz7HbzQ4GdAHOpwG1O9+RdaK7usvd/K3cjcScmILeiRm
LEJLmg/5Kymq/+bFvHiHbdi2yV76HUqT1smRIS+A7JQqixBKSjlD+oP5KQMLoO2RUigD7pWSFtH9
H+0fNFEfle0GhXx4xd7pZpjGA/iiU2dsIFwdp9mMvyr4lIa6TNPDKB3jWC5PJq9Tuf0pEHSuzBF3
/qSMwvcfaM6Ta4w41Y0AWMqGyryIgvbR2jpvHlEDDEs07pRahCkTZ5aXmh+3Ggkqm54yaufLEZ0E
WSSkwP6BOcg4kzsdkA3ndzKypXwpzyoBZXnNqWePvgMvMArQtR1C2TNwFdqaEm5zSaezu9P9u43i
dsjmoVvVEXdLQheQhOm3CcIQfjKnvvUNHhgX13ah5ibk8oa40OCkGFE4+XP44uGMI6wD2VcESu1i
CdLHpyl/G9fThaA8yBHLDdrGtvirrqJNWDsey4b+xsLWWjgRF183hXQmVScOt5ysaQ7solnm341U
N9U0eiDbWHM5L5SIkRzSQhe7fZQjsutq0RfjRHF/95ryH0D3QxxZ3XsvHfcHq3yGEIE0/Wz+h9C1
Uu3gU2ouG1lLxNInWe91ldWF6ar/D5134w46WmZhsS77ifOdhqjMBPuOMZk4LJTi+hGSQYy48LQD
5t2UfHD2caN4xU2pAaHM58J/RHiiCP8oMfuYzN5c/pIrjHycKYHsfVlSZOFmAKxujgJzEF4fcfJk
8sdDwCbOzF/XtQgcchVWX12yjPgbW9RdNR0BJiTeVOw6MHxaMDvggJuKEdP9rU3rUL+r92BAmb9D
XaJNK6YvRTf8UnK1onbx2rDbo40VEq183YUCqeu7WKUnF2FhB300RZ7bhykQEsrfGrwlgxvXY9mP
gA74Xawk13/+sDD8zR1mNew20NP0DZDsKoOEGbOyErmteCHzmpfjLh8WH0qB2qUyJM+Br5GM6vqx
HgDVbnNDxmCkfVggAbqh1zi8jmkae8VUyppYVumYTrK5Sl+QV92E63E6XHsANCnfoVvdlhvrJ4Rc
0FcI1fdLWrh6Q42Tx4xG9fEpZ9XZ3/wFwupMADxB3+xA2uGzOSHpDa7Bg+xb+iuNy//gRc+SNzqy
EqfXH5OJr0BldSmMXKzDLkfWRjHA5/43FivHCeoII3XGcejOR6LXgZn2VNiAtcTvwyFjnupvFfUC
xi5jWBpJynslh6gaxa/GCRlTCfSOR0zRRealSttZe/ZBJQDYcnYGDA/hAWY7NQu180lL8EHiDegt
zX2bjXYUKfGPoXqXaHwSZZdf7VGswJmpsI0WjZGXz1+HvMlrgY1Oakk5BAJjXBH7czoCwO6XBTPu
Vak0Mkc/7LZ6ADd6JbX41fS23y1/pkp9BzcLtSTxu3Yglgh6TGAZwyZiHUVGz81GNyWzg7sogESo
fuV0lXOz2vQrkBDlGqZ5B9OIp2a7D0nl76NP3l3GxWa1kU6UrgqEZRBdtl2Jnpp0dY0kzTOl0xQ8
6x5oCYOCg/NJhzBCv/BmaL1ZH5EcbatRcHAkuMRW+fvnBJ6DErKcArATlRtwFwlHk7LqDRd/c6Aw
V4HIoib9dFgqy4/FuoaSKWDc/ftBCLcbdDnjk9tEpS4EhNqlWM8ZTxaXkU+56FRKQXa5C3H+BOyB
IxDFU1uwijvTXBOwvDLGj54DK8bG0fQZrK5dnj15mBCU0acNSzfpC0dbSzMLRPsioT1eM76Z4cck
jFTaje8Gc/7xSydzY+cmiVqM9PVOnnL1uE/kGAEM2yaQP+VoxcMbHDjULgHHlJCblb66fIxnDvJ6
Nr5Yd2GNLlgRPVlR7ADGXfm3erMACw9gCp8EOT9YIDj1qGGDup1zb5at77KuNLLTmY1LWuSfYpjY
XEniL3KfRPWTZ2cA6UawNVTisuUhtA/WGM3GiSSII5fZssxpvld/xnDx0hUKSXyY2ggqGHTVTH6W
DHabUe2skUdKDAHBAO7QONPOKgYh8c8md/yjdjUK041Zz1c9pfcBksnG/YtA0/e35n6SVU/kJ34s
EndAIWL1w9RD1UMT6/6zgGctQBsqerxUetPt2ftzMPhCtfVj9vVLoApFbv/W0p5q4eylWQxZd3bB
ayAHYkZvhQnRmNcT6eqUE1DTqFsOjj8ChCnId6B1iADhw9fLGFPLob+AWuHCpoHkvUdvGm9GsIoP
iXMrN/QRmtYqwLrFxTXpLzRSnlwliltPgVdVYf80BUv+UwfO3XzW5IN12OblHc0+yq/Qfh+OlN15
YiubIA+wnGwHj6ipx1AO8va47olU0rBhhXxg07q6gBvP3HyTDdrkr0/b7w2B637WUj4K++b4R0Rs
7BVvZzR0aw6qPBQT7ff1l9Rl5/5lxscNbIu+kH84mc1krBqW/9apX4eWXmPLKKgsCsytn2/6vm5v
EKkT4jcPlqVhvTCinfEKySMoi3szw/+QYe4syiPokWhkFbApExrpwlBQe98IzpCKE7Bdc3r2RwFR
l3Tejt67x8a6BBYRrAhaVEQKPn/qPkdIa/DUhTZTRsuqkT3ElxOXSlcmI8/Yt60aZ8ayXuGCLco8
yEYl1bG1EIKTWdhGq96fyULCw9xj1GyoB9unEJdwX/k8IQpWTJCZ0gmptTYWY+MYa0c/repLBG/P
O+8n3ItD6M6eFVhmNl+HXhYMWYPZUF/TlC6kUdMqYwDCM5jmcOaHdXaOn4efTy6w0e1AHTIM73Ks
P3lzM+NoSDBx7pjGPkZOBdkbFN89XkBR2HqMBDJAGbtOwqXntOEUvMaipLf3N9ELtgEsdcjswwE+
hX64bSb1AQ6qa8uOxQnI8d9L6H4hSwy1dErNIc/UWvI3eMLvPFYSGoJ8EuDbh+NTMUIDbsZR9Hfg
QwFKuDYZMmwBGMGS7d58Va8lpDcUk6RMIeD+4bOk9bE94O4ZmqUZDFCuy2EBQbpaXvkp+Joqy8CK
4MFdPBLnSiOg0uI+0zOaW3wxgmGDLlMcAxBV235LSy4DB8PI+2HuGA4yifpJ87lMBR5jpCXQaUCz
ZJJol1Xa50c52q6qWXnlYmpa7nSwTbJB8Z3pszgIeAhKpw5/Fa4zqNPAnSFC0HrsQj9MC1YVbEow
Nqd/PjAS7bWJMJRFLL2BS2+6sQYerufXGwc++sZ5z9EPTMlMcAFaI3coo2NUINSslg8fNKzGE+Hn
pyReei5uSL8ueo1pitH8uiacrwsYaREItlBXtT0nMMVkQWSRdJiMgDxDlTZMbP9pBtQvuuN7VrEW
vyYPEbypOx0sCU1btxdvdAi00te0i7M83JvzkfhxI6IUk/X1CMJaUQQQndaoCzS4Q5daEDC94V/h
tKwU01EiwnUpohIeEX8MS+VbgwzMVFiNO73Tsp33lr9KDEBGc7HmWNQPOXpX4cbpPQH8yA9kPa5h
20C9JB4xu919m6HHZOlSWylhzKaBILeJpgisvXGzklhWNurWaZrxNU8H9WKoSAWHEUe9bO38CyRH
+Bn4Rk2NpvCI9/VG+3KNAU9yp5XZVGJ+i5qIkKR6NxZNuUQDoOxQrckFJskJ37XDZA+YaVijFpMF
z/iXER+pkKlv67rALk8MbCfBFEFf2bCeUYXVue4uFewYr94nPBcrlxCiKSpmamwTmu9VqLq4G/Mm
7WN6Nk1OtEiGPjI1Pd/i9E3qXTe/nOYJJcheGE5rcLl95W74Vb5YkpE3/oXa2C1+qjxPoFmlSQNK
xdIaRnzlp6BaqAyDOOrIlroFHk6Il4ahg9hwHr8LN53ZVLsy2ldCMhTrUfieDtmP2TezcuRglVK0
wckx7BtJArxKzrYcwDMcEKFViS4AMkmMOEmkXUKf993CcpLtSc9XWLVAjNvhxn+g0mMR3lm4aMCq
QLf9K6ToXrb/HKdGxTRzDd/Fra+Tehto7aT+GXIYlm303CUzhznEvlJZ5vfaOq0Prt1+Zf1IOkZy
mbsDnKOfd8ndXEdT6KfqTYg2sLvQYv2c2jinslQwFTPSg+WA112LtU+Uh3CK9uzlli4rAVktEM4B
tFysFcPcilmZb+6qxoeyRWIqzM4oT5GySOuAd771FWtgBgdLf/wYAikI5V4YnmcAeDGbr5GPJ8Ai
6zO9lqrK5LTGNGts/IQ3MkVCOwiExiVo59kmuWsB6G4vlVbfnEwVOSQjigm5+s9y3BPe33asIWFj
C0o9AeZePDmTFlVAQp1oYrTfbSadDvdUvrYNs53k2x0n5r5U4Seqqo+Rl0vEMmAwH/c3cMu1D95B
L5we55fLNLGokKynEFxweMJ5GZMx0vwdEWFn2pd1vPypFRBPs2ah9pvKfiNNqytBxMy+ucX1+onp
BJexDVaoyRo3BsKU/7geLcQeSGINZ35dOfcBcl2CW1M/nNdV9B4xBs4E01Htmx64s6l3EVI5q6Dl
R4BNph5b4EBK0jJcNsIfFY9cMH+ZDC4ga5gI6UYJQe14VOGhuyQl9j9BRKm/ohoXivcMxD36Z6Mq
KiTcFN9A2sc6Z7Zh7CJTgxRhY5FDnXfDH4lCOnMhCsXyx6RiXDv23Wxz6RQc13pqo1GwMhtCjQ4f
2wevFlqbYOvVZpNAKTY3CVYGvDHItoPD3zNC8VaSfnfyrBUyMA5iozTp+7bEAisNr2SR/nH3kNa5
n1MrGkJnthrG2M9U+bGxHV7Y8wmKs0PVx/ksl7G2J2Hw8mv+8iJTIzqj4H/jIBL9krGU3okhiYe6
1SBciID8zkIHAa7QQXMRCXlE4Qj37VI39p46U7WolOWs0+BxRd+xbnSXDN9i34LextJ7ng0D6cg7
SIvYAsgYzPkoBuIsQw1S+OjdED/5aUlwRZP9v4j6vJ7mVlU95gX0fwzRcjDmOJdbS2b7fm9vSGRL
gWQWGw/Y/Ne5E4vi2LHj/dWeVjAuMiqJp+99LrcLRt7cAWdvDyocpsq7TKi/bTLmNkINNQMahkeM
QsnAXS662kWWsYdaqYlOmVCECzpd6PTYkm5KuEM2INl2VzvpJToanhSLdaZ5TlAiOmAXkfdWcxOd
sETFQqKparbJTiNeisUbj+We2DPqSPsTsVibXk8BkGSMZkULJO7x7fpNM40r4eHKPY6gQHNeM1YS
Ox2ANrnqtO4AJbCM2KcZ93kVSjS8aBQLQwx1yMFWdmfKjC1JcdNiwP5uPX1iCVgWwggkZCg+q1ut
3ICfdfvhUUbuIy/iLmwxZL2i0ioqciZ30Vu/vSGbysGZ6PlOnhyBJYP/w7zR4faXrHS/9cMKv2/5
05DKzosJNO1ASXh39feRl5KnQ8trzwze26yd5y/+oN3P8QAPfvh9YpGSsIAZ6i5t0k5XSJ6fGmT4
TdRilEOQ33eYQ75rEo+pTJ/IUpxwvSpdN0LlXEStelsdSRSm5cK5d235JQvxKn/HO1uFjk4e2LBP
ntDq9wfMORS7UDHcQhBqCBT9uVrrHY/tKiIOEKg99G1zzm3g/dlljwNLwn5TpFRnEZRmKx4rVA3t
g5t4HmduapKbMpB5K4wqCfG9D5bVWana5zR8qSybhCkpunIJd0U1WxUXRShZ4eVTrQvxHdI4RxoX
R8h59GefjwHPmNUvZcHYhR8bPaWajXlZ98vF85bT4RPV8LQTPS2+JARFry4+DKm0kCwlc1VCADLz
mor0XL7Hb+gp6YIlQkl+BUeHuF3ML30l6u10Ir5QLuFD68XOua4GRpLNmjQVCVuif8BfFChiJHfh
+4AwQ5xGnYC3JcblFYEclZn/OoD9f71bPIa8W9ERs0g6Kvz3uRdwr0YE71FnPCEZ4kIg92abNLpg
d0GhmArwPW/y55XOS0ocsFrDXyGh8aLcn15EHnOybEHpgQeERDZvveNKyA6jPAO2dwEz1Ia34eZe
7mKcQdvnse2uCVo+2psZCnjHphkmBBRu1Wbs52UwezWcY6pJuky6NnfOKtky7/RcxCGGJsC+7UsZ
Wrov6534NqueN0GtrQRzgrYhg9Hc0W4ks4FegwCvBtDNhZ1ZLfs+8Noa3YEwD7XO/g42WM6IjTss
+Pt/dXg5bcR+YUDAzmfTjClXeSq9t/R+K7cdsxvzvkSxHBm3RppiAZBB8VytrmxkuIAbdoz+gBQk
6a7G+o0ONtDTQiQe2yBNnwrZKeYzYdUU8Tsc1oRr5d/qXbRiZ/udWLJueSwlsPQIfSLSJDXuVahP
cUeLOeEK+jZebabnBG3GCEEFpIYxoCMJeeg+EBEopY4ynMJ8GpDHxkEcMX1U6pdcdcy3HlSvjxjc
Z+CTGnBNi1sWx1EDsv+gHjwMmlVxm6HOEy4GncuI3q2k75PQq8nm2Al27NlNcK7HIaUKMrhMn+vT
StZLPnh6hVqWj6/l9YyfnSbtBRXT8wQr8En2X9zaTm6ZbnnLEPKgvLocxdKG4uQGOnXq1ww6NJ0V
j/SUroBTgudZ4If26/SeISbcCbm7i9+rOZjlM3qFhit72n7bAxruWwN/eNmvbapGGZNAXGLeKp4Z
M2rj+eSMs1kKitTWJ/BwrXjd0UO0S5IxMeRy2jmBPVTXUim5jvG//EiwGZiRolqiBWL+4SCX3/fx
Sim0YVZGRY8KNdptQCch4/uhqZGmBKN7gvg57XjcWEJDSLnEoNcXn5RPnH6KZxcLbzWohSsf2fzZ
5gdynokR1T1XVKTteGuECuF+PkaIARzGa2qL6uKpvS/MsAMh/a73bpAUOqAaFak5ncoKgCQ3A74p
qUU6S8L+C1ssOV2/v3IbCiy0LyPQCbLFPS5ZdjM7GuV4lmMN/mJor+hG+ZY1kgmwjSUcinrya1r0
bn/zgJwoSrHRXpfOeXedYypZQ/SGAwAYdSrMYtMpMWoSEvajfRjCu52qlKHhk51oufcCzUzpQ6Zn
erhArBPVK1LNTmOcZRb6FHsA7dNcecOWfvtqUli+0Ay0L2S9YgC5RM0lf3CINfTc7KCZlRNzCSuR
sP4p1ooyb1bIfo5WgSgYDDX97YQPsfEYg//hVjQyMuJ3Rb6g/ZIlJwTcE4OgNRxguYr+o+xv7GSk
vH5klDptnTyyBvWHG2Syh6ZWJoGYxLcErhmiRh4/Tq0xn0k9iPujWI/dxJTGUrqH+IYxdbcOJeLQ
5sbvNgr+lWCjJAQzjBzuCyKHl9GoixZYBaP9jxh3E1fWV11YSs3F1rcZUOAEPpx6DwGlKbyLf/vv
J3MesPekoF3R951w614byUg16A1oWIRVNdqPM9NPIGW4+BbsBEQvoU0r7IIlHGNPbtIrbyF0zhUP
xJ1VKVsY0tERbywZ/OGEOTxofyjS4BbDtr83bxClwMvK3So2N+8+gMZ46lYIBpcCsax53R/d0e5Y
ir6CbKF02qt4W1plQMMiDmfXFLTgtcbK/6EWGSGV/CK10huqgAwNnW8dxkIf50VV3j7gdq1DEBsf
X37g/HsicvJ+w9QKLixuU29EKTnr+/MDT59DSJt8VTVwE70SDWDwY1PQ4wbiO0wZujn0soIKw4ka
+26TWNaDneer868kj52mO6LukNDGncI+DJsrXpa8OLcsofUHMve+XC7MdRsE4/5r57/AHKfR0fW5
pXdJKerc+tkSXYE33HQwuzE/o1045IiIOTWM+fXvNhEZroyfCreBYbU7tkESnXjUpbLyfQOmXZ9c
aRVbpPeCzyiGhpkAWPnn2Pu69QauzlvdAU9bMjFTpGSe62qxwAE0NG+3IyxhjgKZHW++K6QiC7vg
SvSCSuzJfkRN7j+n1GUR9F4nz+FgAz9Pz/s7JwUYy+VmJqKnwhnnxpSf/vwP/gbHW0J/ObLY029b
AOl8aIcbRxGhzQpGDj3vQyPPKZpGavYb6Jl38gvfrbzJ+bqQQUvkN4Y2r6+NValvAVibCeh5fMgO
L93rscD0MCxDzvaK/RE6RphT+WarJ/DKO/79kgsT6iw9lZq3LMoq1dlMRhzEdeRAf3zNm+y7tXbN
JrLVzrpK6dbp3Tw+3nZSjI3HITHA+3nkv6GSXHAnD/TfMxb64RUNv3n+SjuKzS0WnyqqKSFgfHz2
loFQaY8xouDlE+x6IbJAbIdPy4J7y8Sy/9garEJ3whgLziF48/LJf2tEqEW54WCO/bkc+jxhCdv3
bXKhMjFW6Wv5EoNsGzJJ5bPd+0z6tPgNTDcJoPc68iSGsma5VwoZMVleHnvrN0rG1fBSjX6TqytO
qlD3UaSIZzb4mCG8U84ToU1BRud0B9OKsTefkYaJ5GMNtiolCjlJfTeD84kVezeX2fLLfknsY1tb
PIG2MVW2przDpM6nTAYUmmlhJGWdoDoFE5N4XNV4LvR7Z3bOtFFUcsttj/MiC7xLmYLkP+Ux1R43
09eqz90Dr18rjhKuKMoIqW2wFUe8k2DjuIhFKzjEZTt3wYgl/V8gwgxUkZkiq94UAtbTHLOHNK6V
Oc9uEV3y145Bj2OorjJ1QOg7GqApe/pvPQmVhkKVAjp6LvSx2eVs3ecSwoGUrctCw+ArWASHb3Jj
vzqtXsiM2AnRehbmIf59RRPyBSUm9UE2f915YrZLjATkc3a1mKz/lFP/oVHCl2WvKiAYmoUJGKcB
p42giOfC7c9dwhn2CwUOupWu3C3TRi/edJKI0gjKUa22Ug6EhHS5VvSmm2H2xmi7SPgld3orFQcd
LpnXuHtisDR6ayY2qdkMTmZ50KOO2Q4bOmQX+c7Rgb2SuPT4Mg81xAkF+POYaFah86uEEYJnFhT6
GF9vZ04kHC+Tx4UQjvvrsF66R2/18jWV4/93LNr4xRNYbtxMlGaj7yBIAA0k9R92qqScotjypvIf
aiegrTsrpqvPhrmjZNN+pv6X9rn9OdlB70hE0/yKUY/RTBsKeFqxE7vWziFoZPN0WW1Lh/049Xpq
F3Tpj5SH6aIbKiCNWTbidMqPc2VfkS6aivz9KCMP6ZCWTdFugeY0HoEwVHM0lBVzkAyLTLImBZom
HLgDyz1T6Jx3FEMLZAYs9vXXKj5/ZGsmpRDGcOgTnWC8m/ZYcFIkVJD2iKqmH2u+9WsmtXQ2yDCm
4J/31wMnvAqw8eKV5cf0Mez6LjCnUdh8FUJ0PaXi7tMJsUcK1FPZeSr4FB0w9BdV5buZ6WhHrVXf
BydJ24p8PfFPDkZJCv7uQ0K4NO+Kdcll+B8JechgiFDmZAnYEHvkEsPzG/rgD4tm3C+bL1nROpbh
Y+9NOV2y1hPYwpK9J5Yw+utBhzJVjspDowIKGMa/W/lufIXtIcA3MR8COlMOJwnOUb3rQ8hZuLHV
Th18ZYm5BRCA+kODGTBEyzQ98gE4sdRmGgWOhyUvO3v6Sg9Mz4yShlVUwk1RkWOybrM/Deus8/tO
jcNT3vEhyHONrypkKOQZTwImCnXEMzFPSTYSJxZT2nKm+uUCUxXMoM+fw8pKa8nP8PeSHw89bpgd
MwjzlK0sxPZnLnPjbHsgtKK9LfjBR1LRQ3WL7Scv/MUG+bfTGDMjRQYaz8efupwtbcuh1ZJ1GcWS
hjHCDsK2fOAbpa7YhBVy3OezDjmMTTqaL9g0JHfZnREFgSvYbpIyUEqaoXanNet+Kxmv1evnHlAf
o74BZ+YxlP1QobWPpmQ6chGsZc6FNedCkXyeuvFR45xS52c9kb89TnAvGkW4Fzc7mNjKJXp+t/e6
kHDYLPh5GBGtdC4EbLuZ13rjl7wwgxzjxQz54zfqyKHJLm1GuKnSmUC54jq9sLZEqRkwQtmxzBnG
txvF0+LNTHNOj6czTMQw8Wo2wvtX/rA5v2Z06XWWBwy77clwUCsgwV1QnWYwgqE7FZEesthUzrEt
c6BU7orrNBHzV/LcEb5ztp5oNVunxxdX2xT/vuHUoVyAbrVlYcIby4QNIAytllzBVhrywDHEGZFW
6h05OFOj1fZXWM58pJkpADiS/cgL0UecCLiK28PZqc/Tv+FhYB+LMZ9y6sYuUJdhKrC44fGkV9Bq
V4cWMQ8hXSwQN7cRv/5Mn/YKFcSGDXMkrt+qakF7mICG847vpO/58B++F1m20uM/9/hh5B7gxU6y
Em8d7fEbvzy8wxOoU7wYC8N0c6ptg27Vl19D1+SxWUXZ5EbjwgoGiMtMAjs8ZoB7rM1Sq3oSilKR
haJRzdFFsRhkKwtlAP8NbPvoxoj0j6Lwow1KzQzk7rERdeFudUeHnEmtGrDsHmgmZ1F1cToZbOKx
Hwit5zUs90wLyay72TM+jWudLJQKz2fGG1R6cEeKJNww2Ukvs5MccFsQ24un6FB7HH1lus/rzSOE
z0KITPWwzG0ZIlN/irreQmSj+oLFv9At0UjDSjq4eRyDpTsvs+ZBSrtMXAbeNR0NllS9tNaWtbZq
Y+ES/pwykiu5AzyUKK32upQBmtuje8sVq9QNgFT0Vtxws1eGliu5OW6t2tX4ewCsKoUwn/lN2Hw1
j0jnWZ+mFBJvb8NePcJ6TRdASdI0jwXUm/i5XBCfapl62/PMulggPgSmCMeGmPlue/FxTlqpr04T
7WGZ+rQb4bZBfDRm1ZrgQcCzwwQ+dZIP8xnWtihXYFctiGgTXAJxFyiRyVB4PpR7uIdoHgKiItwI
AaHIcWf3QW2arh+cTH7tVwEWdRkKvnBn9HuBXxn7/xkF6AQXoigL65t0plrqgANYstnxXMbSpU4n
a7n6N1tWJDbtbxgVByAGiRkeJa2w8vyWHTAiO9TB8A2bXlvU7/jLWc4qBNgKj0J99gAIRj1bTGLr
tccFIsVVF+RMoUDqudA9rqxzak91f8k5GM1YblLwEEwOlsa9xXzPj57e+KYyF8rlqLvxRv6Kvno8
hjjy7pPEastKuMsTGsIcD3dP1+A7FSbzdYFLTzkX1IGFTcovnRFtdluxVi3iKJ8Eq5o5+XQJThNc
nc0qvP0UpX7VezZ/KSCTV/p/hjTGeIiV/B1wUl4JTjbydtXbQsMIDpVHF7teBbZE4YHj71pHTv7o
/nub3s1mwgdUJ8iXmD1Jd7mviBjsG4RLLJPDRX4yNPczO59qH5dqOO49rRKCP8WCXOsA2P6yNjzt
zuxEknq67nbYoPeGgzlxL1NGxxK0Y8tWk05ZaXEaZnKEEpf+7Urx/G08qeaQhELjNmlmJIIhDoYS
ozadmmJ6T9ytch9BE7YGz5x0O9CBsaktNMeWDD1F4qsfU6Dlv1pn5ekeda54PUvrQEGHD7V0727O
byzHKcrGGqCC2Zc5zL5+Emx7Wpyj5M+Xr8moFmmsD0t0Ln5ZPjUFHqozWFLTz3QMIPtvPR06n6+Y
+Taqxa6jN1vjys0ai/RMu7URR4eaVDtEDuRPptU0RQgepd6YKXnlLyC83nDQv3sQwmjOYurZuz4c
DKbIOYV0ttw6yjszyXyfckxlJLaaLzbFgjZ6ZAz3XCVgcvyjMQr5ajTIIodDEYO7zBOWTaLjnJuU
AUekmlEHxSkpNJjPqFQuNCTu8Fl40nuZLeJbCXjsLpWkoN3o/NailvXzi9SAd1htmHiIjGWtTptN
pPNXvsi3CCzVcSouXW6PA3d07zcwTYoqD7Q3h57p2JjaYJ/AnyTR5VFBamZlHk8Q2jQom3ds59yF
xCUKNnKbvIaAFW7fDCsgT7Bs34kjXlWteHyPEVhuujFqIOVVOedkizQsDVhMJtEUtWBEm0dscQh6
I7ImcVYWV5//xk28PyUwdjuiZUK4PyfVsVeFpjOeWENvce5z5SwOcRD6zkRCbfEWSsTO7MODbJfN
e8a+8RiihEdINfHZQtZKd61gbXko3u3Xid7PO7Y4/uGMCNaCh3I3oJ16zs0pbpxZNcm2vm/QiLYz
DqYRrweWVbRKedqlVHZlE6LX9xCrIoRbjvAzvgOTFhQhC9vqWG9DpI60r0dXJoUGt3RDMUT7oHJm
AwRpz70Yc84Y4iv6Tm66OxG3b0/sKcyFeqKCR98PjccH1fF+rUuw+t3Nlrek8ANnz9LjJWh805Oa
SY56REcNjTQi3q3g2L1vPDd4BkGbXfgD4UoDl8IiXuvqWU/6u0z3b4f0i/jQJ51wz6KV1Y7ABAew
Z31MkS+wx8VqWdlpUrzO1zwm47lgGJZthsbmKwwuyjZcSW36rN4TMwVr0ZQek6OsRmSo7N5732BU
Y8zlyrp0K8fgELIn/vDmbPnoas/gR9g+p5oGrB1KdGxEuElouxKDMsjsjGvNsrg0llqONlYrV0hc
AxCzOzEDoztzfbmSLbtJHZC7GU2vbZ6Tn6EIJtG01RpzLjNJYIc9I7JpbMHBzuy0qXfVbDDOwGL8
HmptrDR7yMbFsMRWZ810Q8YRHIdE0nRE/I+GhxSF/xLDBJLne8Jb1pioI7yxdR1dtBjvJWltE8H4
zq6xRlSUBWQ3ccXvSfeks0URlnYnsiZwKKDXWtVDmsn4gCvkPttTaesgmKfCL1T00HYiEtpCM9GF
WhTYfSeNrnMuTAIjcoTUNbAmtmZJzF/Qito09QTlbjuP+RqywixAAnVhvceBpLRw8+FDUrZoVGKP
Mf+rUBdXtJN2LFgg7VOeTMDoyokevpvasOF6Lzl71fhXul371BR7lCFU/G6TMaU79BVPPPQhfF9G
WOMHmp3QD75g2X3TcSKqecFLOem+Ye+utitYJWh+ZTH8KsP37sUuv8lb4ttxhmXcInYIwUmNGE42
djJwsYOkhc6en83nbOL316Q3YiopaaMVfiYxc99SIzIpdRdlGNq4YppSVdhVfCOx75Mln+t0IDQT
pnzXPN4xycBLCVdretcxsAHCrK8bIydxmWuVAM45Ji9yLIjss43l5ZPi5bjlSWUPXkupI8oWMEFQ
6T7BoHKOZNP6n5kVOV6GWJhg26YgS0KLz6OATTqTS/2GDXY8SbShBbZcchjWcsaU5Cc0/bNmXIFs
KMMqSvV0wiuDFtdbcYIgkb0TXebvKCQUpzHAFCIeedGD1C2Yk2Dt5FpuG184Q/sg6+K5SwQEdyuB
LHh1UtxkCu5j2QSMvuPiD2JY8Lt/GZt8ovvVBg66QqL1T1jn5Oz+7kJgdlF3fvHNk9Lifm1Fxs1F
agsQU0atuJc3k8lHxgqwj9FGlsMs/ldW/LrQdmhPSigbMB1DafdSR7NzyLzo4/wZQp92REEpR/HB
4QInlR7jKCC28kd9y4ct2rffeEGARFNmvBnDpOWI0aoJJUU9RcXpTeK94XVxhAwjAk+6EK7x5T2P
ALDMrWcZo0GieYI7Z7furU+rn1uageXt1KmcJyBe0nWSJg9KMF3l2N51TDamQQed7r6NygAqf+OU
vClWFCf6FDsx1DNUaH+EgCY7zu6j2+sGItuAQzW4UjeaD/gtPCX+b0rFFmOFed8MtQaYy6EyL9B4
Mazs+aCT8szIxdqCegNZX5Wnou1MqGzrPeBwYN5JQ61KNlnup7gzIKJMeuRYKaAUkp7G7VA6vjPA
aAvGiJS2YDvgWJ84FvJ+zQVAO4o2725/h6/34VqPPT/LSIXkfVikehfbZ6LkyG4Cp394W/ChyM6D
2CL3Ir99wsH1Q+H7AduIkYZ8GLRJcCq3izHhETC+BIQXVQbZ/cVeFALxuGtXPata5t6DE/CkRYQm
ZHG5YqjEFJOYQb1WUyM3hHQyNq0vO2T34eawk8Hp85M9T4XyqtkCt8TgoQICGZ7z3LomeTsX8w3E
QM47DjRZHlEP+P4+0CysG0iGyTTxUQO+CHxzN1eqTFjzMKk+rES+AbsEx7igj7eYMTAgINAqPju1
U2V9VjNSJykFdhQnVlzXpaWrRf6CWFuronyRjLZZbHu0dg01vnFnxymvkxCFwQsDXVAezrHVM/n8
1fB3ip3LSxp5ieXG1qzbI6WiCivwxcB5pKLgINHAX2V8D4uiNlWlbbBmwsbXUI3C8BmLNnGj/mW4
KZUWAdc6L2R/Vnz74cEMNUTjVycRfTzch7fKUCBOFn3D3zn/HcD9vDiCKTokfq8i/0d5C7vNbeE4
gCDxH2efwVNlCW+Z23HBMnJ1HHHJrwmdIHbdVkT2e9G2R/EanAUGfSg7u+p+BjYVK3DVaC/WlbIe
2gZ+7Ayv0RGbAVLx6HQwoTNaszHe0QLc6eAQir/Z1p35cruBYSPuNMbzBv5Ao9xXoVf6gQRoZt3Z
TohSBvGv4IYXgeBotRPdHawb9jc+vi96vQ8mqpqAsDV/4wJi5HdTPJNt+L9GUqsUzyLn8qf0Gtoh
Rz6vYsq6MTq6lEA9aJ9Kv2YL2x3rUdrpYfovXmeCHPeqSLxw74s88zaqs15zOu0veB2ipCMmq+zE
uefPGxtwOcFZeLHKr2u+4twER25HJ/y+T8CvOgyjDiaFGd6vS85iHvQz+pC9OJY5VbqXVn5+Lmwx
VGTauPrirvz7RGYsPc0T9rLgmmPmXSU3XBFN8lK52VIaVhOFC/jC+/MgL9wHGqyJLiN3YuRZGgwz
PKvP5GEAfbltggcfJFZ0obiZJOYxWVzDSmpYBDBgbRjEwhIZ3j+fzka40eb70z8qSrpRImnsJpRk
MuqgPR2sjocc9WXyug+MwZQygdhxvuzRyzZB2odB1UJtiHM6BkEFF7szmvk1Z1zFyLwyz3HtxNAU
1ZJu2nDtiph71XtIoMb+B+jsobOxp133jLMvHt65G4EI0cmJ30xd6ITBMNzwvX5taAr1P9jKS/1/
5le1nJ5Nb1i156o9Qkh0gL56m+EcvfRTBeYwJ4xYRn7UsAS7TyBXjJ100aFJOfieRt6WUEXZeq7b
SQEoxoTm5qzJXZ8UuDbBIrGZlmB2kKOcqb2+8GG+R+WecO/XZ3Rhxu3ZXlxhAvWSorzqaTnpu7KS
ROAKInT1PbiPfZCA/GB26sa0eMjoYULGrDF1D2vGq+hF9pxFc6ca7T4KSrXWtLcYZdXhIZn6+mEJ
lY/SbYdAbUZgRXJ8q++VSbuihtDy0QmKk70wuuB2yVkFUqZnpGLfRlI2BJu2QQWqjAQjLP5XfGDJ
AIKCcqNb/qoWtTzSJPpDgX8tJgWYICS8j2/VD4CvoMZoPkJmjh57VOpMojaQlkGax55FpKtlwRAH
m1xRvYmg4Dp35PoYRopweHYK28xlgwaqd6jTg1ww5My4uP5kYJ0BqstRU/W07wlLmir+HTjrO7WB
I7fnNJPX/e/u6OIkH0VuvLvo2wMlE2O4C1+LRaw+nrH+WtpsATHC+AsyTOBfdcsafBTQafMoDsuD
YxVLrqI+/QbnH3wAJb4L6W6+WX7yviNn/9yVikfD5at1r1QF6HuBticxBdxwJGc1uYwPREphKOpT
A05Cvr0N1MPREhtGEhKsp5cY+hoHAlsIbG0nag4MAx+PuWZ3gHs/M6+TR1paVHe0nmvWOmfACwvB
CLWby0HR+Hx5o+cWiVBul/tikmq03J+obCQgDGiLEjr/8cOP4g16bJEdHTeJjdu7ATlD18ukvCrI
oWrDBPVgKHM8EjkzGX+diZqhL0bWEfj9VCM1k4v8IaDqQwsDQr+VrcER39KckBVnoBFg7nzsR9ME
MsZwL5N/FvenFP1s2+Nep4dYrAzwda5XQoXmC1Tqpf7Ua4dFZCQg8lLPXkDynRV8bhviaGjqdFPr
um1ABLj7JY194usQBabG/FI/T3qgJLgd7m+BrLEcqxAxpB7uKhzM7NP0nCLJafsSSi/ankLKfOzR
NtT6f+f3+WmQQm0iqLDGa8e1ykvFFLYKxwEkO4mlTVVdc8DVzjKR8Z7e5iTcgLGn/d4X4R4sTD24
DOvE5zDbIpf4ncWgxhMNY9GFNoWCM5td5WFE1/WVX72h8FQ0Jp47aqnOztp12HdaJg/SSmXP7BIK
kVhUF9LjC5xbsw5uCQpnCg/klLoi0V+PZbpUBVnO2wosYjAgxFlz9izzqQhb+G8mzlMVbJT71sEc
cWSx4/dQ3OMNJ1zynclx+y3li/1a4c+sTb6lfxXcqTqLTv/TTWsdD+sIu/7hVfZVaG7tLNZHeb1U
QsIkBIGgzeAaBzO5yzfLCY/3sIOTZ4QZ7LlY1rVm7U9yOa5WMjVFSQCfDmd/7fKseDiOl02beeTW
M+bwihzXqVjhxjAG5+kz9ghTUeOZJ3ialss7pF7KOsE0Gp8ANhB6EyFPYD5i1hv9QsuU8qdTg4Tt
BVJEckiK8APM4b1iG9hBZmhwEOeHbEZxKL+Pdj/lfLwVhYtktW6grgdpzekK0aIwZ1cWwuM8ScPJ
dUuHbVtdXLPGLYEl0orU0W4QeN4c0LHmlMWf9stw7sUIWzM+bd1UktZMGjVDN+CjLjDS5yyoJ1Bu
69tZGzLfsKMU98eSzHLVwuva0SfndcgcTjmhWJLht/WVJPUeSMpl5fDIm1lgmvN+fTrsHyk3DOAZ
tJF4jkD7AN9ZjQpNopOqms1n4+JA221cjanEzYENQ+I8vwocfsDas3Kc/kIdOydfNscBLYB10FPT
tcxcBSPtlXnrsq4VVcuhDNp+nMkHI9HTMcfbHwaJ23sl1wQkIOqAhSzaM6dqLQEtfcImTIc9MH13
YiWhWuUUgMh0TP4Ip1p2wntEFpKfTDMkmW2RL5h9AGNAjK0vH3r2BAAaSpcw7HdHhBdntfNQJbId
Jck3kLzQAp/LamU7sarmQPG0Zv4HX7gVyqwJoiA7/6UceBNkqmcIkhHVcXwUu1kax19mOUSONVID
ZentdV5Hv5Dr9BHa8H7hlxcimUA2S60WJ0vNq/ul6iTSilcCLJ3eK9OVgR4mtLy/ACG/62m0krAA
mfTtGcohrkJ9h58lyMmMqfUD6CZqU6eV1WoMIG1K5JpDXybFPlKbiSH5mrtGszbKAjAarg1qs+4t
aTKiw5ykYfQjM1gAwpul3ov2EwTFLxCWCA39KA/b73ytf/w5XSDUqRQuTExhEXMKN6evrBzQYL02
Rzf513tkIrreb9bvC6BtrFXPkO+clIp8YvubXQaFSM+ryLR2d9cC7Fo4ksbOiyTeIt7GGUZa6kyE
1tyb0W3HKAPtyXDTNy6sFlcD2RMARIUItpSZYAO9IXbPVXuPb6uDuaBnrYqtM6hqX2KRCVGCK/yL
r1RM4xGbKlZr4oZvDeifdAFkwKjGq4NsSV8Pv/e0Gq8bJfaXVfW7VtrzasR+e7ulCunHyRdDZZUm
8dU+krLoRuke1HqeArhwt8+STIPkMFPODl/JC1mwexf8kZrYU1LkTG81t3d8QnWBR+hXrlgtbiD9
T3299gSot4I+Sc7IIexXvFUZZtp142oFQbs1SGtlhzVRAkDefSXV+isYzVWRKZEPupxV1CxfaiDx
HjxRd8HNXjymO18hSDi8X6pFeUa6oHukOr04BPMTp200GIM+nFjkZDBbOXDHeZQ93YWZwS7/I+3P
l1FckzAzcjLgUcHRi/nKB7DO0UzquFpSybiOJNMW/g0WgSPx0LKs1G38pC3L0JB8r8mDXpLHZd+G
uOjwOMeA4h23rzoHUXAmGGc41QoQUQ1xtHMA2xeqWMQCSKrudv53pT9VYdlRLgk7CMmEX5JBQmCj
PcKZpDHicWP1cwOJYPkMvFEV7VkuJoBvYaBjEiTDvCmphV4QEjEqxPhunvEZhbfRfnIDBzpb6xNF
zp6nZTG0zy3P5bc6k5amm+y8y9yKL214pkGJsnx6Dt21OKAEyxbZkMk7bbLL8hH+aG1bjSUg360X
jUewRB6M7KLCrCmva/OBw2ZOMWvC9W57npP4UqbjD2Fv4iVb+ov/V6KEw5QC+uwSLcuH9EW+E6Lr
8w6kuIB8Pg+Kyu5TAbIcEQWszqnTQsDQPp3dWWWCpTemCVAuPTXdmqUT4qXwDN26TalZSO2qyxrC
vrBZm0id4iCptkV7tOo2vwYCT2Tb9jEH3dUzHC4s8SCfNXHHp6HfB709YIxcF0m7tOPoIjWodES9
0TguxzhY9+ZkNRVOYhU/mO4oVny9H2LK0nb6y/t4c3GkI6dZnaZDcob+Gw1NAnPKIJPUi9uiCJnz
hMTass4qwdAGrbGAJgPKroY7lGe/QQ8G1Jonh+DYw1H6a6tvuE5Vuj2hXddoeDbeeA/uwcDO2q/F
qmwB4k8/HPLQ/Gd3fOv5j7vIivXNFuz14AZmpoXt9ZBIudUwu+sytJtKt//i37u2kGr4Nd5Jo06H
PbN8WqIpxddGXF4Iivk+/RvpS7f241aEN4kR9hzAcCdaSwSAKsMbceLNPQlA/fLZ7mF6vzQTtY3e
o0iYs5zFSg81l61SmfEzPBfYmiC/g+XWek6m6RZpBDSMqtHX+BIOqFJNSlqU7b+GkDH9H0lP7fzh
CwuFbwb6wZZ8TtwvZ0qPSjhk+JfLHQIS6rU1xH9ObOXOg+fFOl281ZWeVCxGYvW18XfN2Myl59dE
Ev5Z7/QSPHRs0+oYL5R9YKWqaIlF+NoAYl2Gp1fPLZq143cv+rvpJ1aHagiBbaCA9A7e52K9eBiH
euloZbu0rxILrGDCHb+PYEG8o2WIeRe95mGd5OIhX0PKK2oXeHyDAXmS0cqsmIlORe5R8RAYlBz8
WIKk3/wrW2v1epKqdI+cUj+kZEIcePn5k1TdfUyq2VCIsW05HFeSnVU/XFaOvMCA8DtSMEfOxZwl
nZ2YNDijEWIkrJyVwigNm+1MN3BaOtY6H/bGHNaaoS7sgsvngbZwOmtm6IYvL2kr/XzI3DTB7M7l
0SeJUdpH9v3xVpJt4L/TinD17XJMRdrcwFpPEO6K4/NzMBuMYxajG7TbvyZLvt/ZqY0/JEDWIsUX
Dv7ZHGrSYuWFed2159LO3GpX2cYrAJI1DAhPGmo2QBr1UK1/cHYU0CYqcn0UqFaK+JWEtmbsDnzN
GqXwal4xcSr9h3mDxQ4NfDb37oH0OTx7Rqezl5RI4XVK4kJDac0tIdKCZaPq2STLINg9HzrJeo05
w+olqt/BcEhbwd5rJQGTtXpq15QBlaNflgL1q8wkeUxzbrkD4YY/id5uCgTcWOsuCeyFn3fTLL+k
sGbvzJa6tJbFpRNvZWkUHxq7ACRspwLD7QkONl0FUgHE64WHpqW2UIsND4cT3CN8OMzFqc6UzzsM
R4H1cEpARYkFQitLWcrH0Uq4UN32w4jcHucxHu6LX/g2lm0TEH37Bl6brSJ29eKDrC4Klb7W3/l2
bmW5wUxAvdaZJh0ruJSbHenMhC4PyxhY94fO/JzhwRA21zn7HWvXLbVbLsj0nS28xDJuNCp+0tnn
VmoOfahOFcNBZu2VOqyQbycpZW1VCJU0FIQjeH6F6CUU+kz7Haz9VhHYCfRsQWkWfinS+jtAD6Sw
cIMv8tEAkI55z00/+cJHvtL+Nw/U4U8sMRKCg+dRHCCcYO3PGQow1tYPNuTYz8eJ7GONkBK9F2md
qRZt+kzAdrM5ROgVxkA0KPtbwaLw6QDvge2uJPHUShUxCddBni2l31q3wcP3XuY+g5tn+rwaxMWe
9Y2KmGOXg5EULh2ZogIggLg8JmgNeXinGzP4TVDTGN8yZ5NhAF0erDy+TG0IQCxiWBnkHNKkmPS6
Gg6KGagV/MZzxvkAuGNWe6F4T1xVqgth8+gw6x33Mrk3LPbkaGkB2lzptFm52Ubapsf7fAaccH6F
qWGCXoDYU3apu9RPdrOrH6QgFkILojsksvkVkvnePFPhZkpNwneBcvoje9jS4swyrpXOuQwgHcb8
DJtq7Z7LWENAhQ2qEH/QS/M0vo+sklRT67e7MBh2vms8LXfHcG5QRUh0QUiPg0h5066I7fIcIp3P
2CoB2PExjzBHu6rjDQkyOcvNH43kcFIwYrie5yxuJ/2dXi5/3GS0Wd1Vc2aI6QfRxatZRs4AhFCF
6p3RJN98l/XxaMg3AT7mnqRqdSqzs5wDmqgwAL05/UyLEkeF6q5k3UeZPrBf7kc28zuQAjjNrBPw
bOlt7P4voamhcP2xYjPSuMYlRRk66F+g6WN3XJyTsPCGZqNhvs3tezIC2eUhCCIUyAM2ZBRh8fXL
iTC7ZvBHZ5CdWJWBJRXz86DujcJjA2LeggKE6JpQbWxbkgHOieyPBhLtqqHmzbVvFzMvZoD+4EDE
LaMH6E3h0gPiJyz2h7qz1LWVq1LBubI5f7vKCO1I++exvkAfGcTOq9le/LCQq+tMDO0bBIUuTcrg
C5+Hs4lj5uAlPNUufwPkreYhU4NR3e/t5YqVu/Kik5tY46uYIc2J4YGLIsA7EwpuYljXRRRRSd+H
vjQ+GdY7EQwDv50QMzATFe3wjiYumJ6mznawwfxnItS18HK19uruzKWf++24kA4DVkRsgJBS61Eo
ZsR9tu16Op0jh+7KjpTldfSD917DoJ/3e1SRtxU5dd491SmcOWfUlA7GDAWUTz2qsgbTjJNOtLKd
4Q6g8xRne1UZwa4SNg6Ul7eA9rqBf7J3swkir7Ug8q8pazOBfPcUq3PrUmkutSgbIhjD0m7iq/Ht
sX5F478rGtitFl1U7AMEUwWOl8FCM1tcU/ZVddmKcaXWPeUJa+0w2iVdc08+ZYG0aXwcc1Zdcd/3
X+V604NxQYtbaonlA2TzkjDdiFDCKrIh6WTHm1rle1hpvR8J37nhUTkRRVZ7bPTh5c6B0ETM9U23
QuUQfimaN+nPlDQoXMZtSf+myi5AAFIZiB/v6hiMigqDobiQ2qTTw2224iR+vFNQRHMZt15hDh5d
n7Hh/KvTZYIgxS1+Iw60oFNt5kJMNnX/8hH5URhGvAtrO+4+oZTPKPu12ZKsSLBZZSlXwKGoRztN
NDuNTQ7HQtD38WlqsVfbEeyhOMsyqQ5/aoybirO4vIBOK2suFjCHR0bt1fhf91Lnoe/slj8Oe6IQ
ybsz5NWyCqjbgTOile2dfpV01NsttriIjd9/msS74S2QT4rsJRdYD/yq9yR+0HlCaJFTJnLOIuc9
leHIh8Ljvujgi01H77d1qYO2HLGzmSRxer1Xx1y9V+jagXTZk6iYYj4JuCLV/6BSfyQic1BqAP5H
i9w4j+8CybOtwVNtOSL8oDtE2nBpT3YvSB0iJg7yvRWX51kzcigdWZ7A1TRJg+WSvtfyujNV3zvx
OXkIjEkEdu/V1jSbbC1HjMoa/DdjD4R+bEoPbsH8fAO3p5xjl5X5pzCUHF5DycUbZAmR8qgWgyGM
XASPaPLzuwfLiDLYcSkuKyvcrIv4PTWA+BGm1c+PjhZI844xJMfztD9iYz5XOmd9M7vadiqsvt1r
P7s9TLWEWWsOSf5A2Joec8renaYHax/lEIazTLfID5TDK5i4xCE52JVN5xKSu9F1PmgxenwWZoju
1btx8XCdCO7XmurL/o3btgrSe5b38ScQCw9b306dWa4b0vuCCrtUZQbIqvFZTOHkB71aLjspBNAa
sY1QW0cPpXF+13tFY4m2VFUMHMxne720kBYmuebogf4OSqr1orICStmPLLznYOnqIjvAJoBbPSeJ
jwvmlAHZWH7lxRCYSUMFHnJJzlfVtYAV6FFN54Rzw8vtaD+GxUGkaRSCwyS6D7ZblAfRRx7eskdQ
3OiDqw93Nzx8Kj4kGHAfaWOun2s5aNR0j2R0/WUfHesAdLZKOk7lYAltZ9UoU40ATtBpwlEsQfWa
p8t+xmMbyw6YZnFidNBOgyhIxLRt3KXRCTfRFn0RtDC0/ibBXxTbuRLnxSJd8YgD7GmmB6Mf4YgG
cIhTPBxnUX52REVyrUbImPD1ZSvTpWHJIP1gVVCn9lA4U4G5Mk9fJftmO7GKgxZeqcw6zzrEtXde
iiIva1nvrk1+u9A7HWcTJwg3VBU8VKgBeWZkaHAxw8tA+B5a4DH58i9pSRyEqcM89zWFXUXhqlwq
tn9M5QuToJmgoyhjR0UC9m7uaoxy8A/V/+APWbr2i8gp5AXI7w6VqAL5F77pgkNZ61hpQJgGaS9q
sEhRmSzBeEdD5I4HL7pPSqNZ2vCTqC3wtHhxGJpJ+pOWTc/5/flEW/fZnvcMzoPc8Z1UOGsT/K4f
dbSLUWoTsyKsQrZGXfpnP5cHPcR4XBQV+1nTeYwKNX+VrZcTvJSG5Dsugq3P43YE0xhuC91RsV/d
rVAOppr6yawVwmEmpLXHwBjSG/lVDC6Q5l7/SM7VF9+8bkc9WhHSne5/BL3GowR6dfHvwLQMAWRl
OuB3CKOWO5lucH1VvH+OLpf1Mge2xAqT8q0zJsdBr/od+so5QEOtM02j1Eoje27AILX6B4/VPpqj
hA4T43z3KYumc83aZQHAqrU+bVioM+ysJGJaM2MB+zCXvgvZxo4FhJmKH/DDJFqp2Vg2kVb+p5g3
voIiMqCwojc3gRz2dXjYhiGwwvailL+ngzNpL7zHD+4NYXytTEToHZybbLH/jY2R/58MrW5X2Dod
rrWOZfCSAlxDEV8g2DKy1+715VTnGPnh8iCVBZn89tpRV1NuyDnmr2+hAYOP5l/SbEXlIhYxv77e
RWeOT8fNVS4lql02rttfp8Ugy2oC5E2OS8tmDieCIXeuSmBI90zfbqfjyhTxXpLCAoeVlOpjw0PL
vgSv9AFSkZS5NmvVny8edUXNH9KffgtRdJMflEhvy9qlJQPX5Udb7Rj0bwpStP+MosqiUThFijcP
A+YhL3PnzXkk1kTY1S8QuXhY3quQ2mdMA4k1lroBd0Py4bEfZPzluCkljLmawY2KlmSqCmWEcGBe
G/t0jDBRRm3V5UWrNyX/LbhbQohaFEQSWqKRnOn2Pcl3/qj4YEqdM+P6cR6jt8YVrMcnKhjudkjR
PHI1MvhSatmYYdw59eHYIccu6wwZ8yxmfVGiQVESPC1XZg1b5rO69Bnsr8g5SwfuzoveeGHzNEcX
Xjq/9+enQwsIz4uRFuO8BltS5+KTytP+QJvHycKXKjFyBSbqzhe9Dp6vcst5YbVnhOrEWyo2hi3r
eLEjjBpIdWlqpG8Spe+OVstX+NiuZKXpjqL0DHYv3Np4jM+yOEn7Xgs/zY47hMFxX/JZ1ethMLxr
miQ/PTZhQbYPTNN2SdS/EppW+4qQ89vjVTs082qFocbMQc/5bJD0OIuRCycT0WNLEXPDRrybhhXH
5OXHS8g3rmrdsrLAucoJKpETmnAqdZU1u1WH4flsCnJRPKIqpKKMbbyNtyR06zl+VtCTHxyuWxdv
ALMKHl/gC4j99vz7Ma2jnFGR81kKPb/Gi6HNIWq8JrpBgAq7t40HDop0DBlCorg3KktrGSXPqLbv
oER/8fU+/2UOQklHAnUIdYdh8DgyG4wRw2atiP8EjEDweS+B5R8tqqGzig42gebgd/NR3H7OYjEG
9OedeQpdPUGLNtoE4LpZ3BBeu3KqiDI+15SCOXj8YnAnrzStCIqhdqCgiRezoYAaI4OTskmDkQQ7
oqk+7HzgduVOGZTxYvRRlM3WXmt0gK4t8HZaUHbmDJh9+08CCRxeleJUSvvTnSSbB/KbZP3zO/fQ
eA/XUnUdF0vkZ8OYGjx54MssDtLmgek8KLZ1Pzy3EqZZuAajXazIF73ZQLl0p5tctAoXb7X9XLJd
RWf92c4k/3b0vzLs6U7X54GQagNqN8DGMVl/RttaCbOi4V1J/6IU3pGJmpn5SSc/g0V0mhoSuL8N
gPt3I0iqHoIC+tSrMR8rxO5cL9mKrwXF0bjpdIUFYpiDT6dlpY4dy8+6ni2fjDfrKPrrjKSbQWyI
3lkIeeAWU5Ppoym6k5unU7oVMrZxClvl2hfjWy5ISUFDfO3GWeVpWwZqyogI1tw9lsWwPgSqoVL4
EI55GmkErCvXdK6PIkBwtd/QloBZkWo10eLZrKKOTR/Ha1M29VDvgEmJYThJC67v1j8e1NOWPkh2
E43vdWlodLck7+7sQ43mAhJYO9zEj71Ag7kB9vlqegPBpaUjDdLHvJrroM6dZBVHF7xfNEVcHNhI
1N6hv5JuT08g/tRuc4pl7Z81JJTgziCG83BSfK/T38oVUCGp9odYARu6On5+hP+nTKeAjBClViIs
6vFesrwKpSg/OQ4Ka5buVW9nXb2vgpYJbsu2KkuMgLuIcIVE6iRhjwYYV3lzaQTVyMFpt7K5bq4+
J1p9Cgo/yDk9jEXL6YR7X8AqqqWZ5+jOeaEA5E/Ua+YsZ2jyP1uoSonezwdx1bAJ7A5hBnMfcAC2
8Gig9Rhdu3Trc1uzO+WCHSAnlPn/aQERbtSfKAwROahNVegFpedtkCjIocLk+HjUp66kYEtzFUt5
Z/CtChWMco/pQ1SJ8RodreE3ljcpmNay6YCDpd7jBY+Z5jsmEmSh3UwkqelfLA2dxEDtdapQYH9/
reLaWCJ298ftPBQP9Kdrp6O5OZFmWBT9q5pNIgCl7p6XqWadairHcqbOQBucy8cWI/hWxHJVjxLE
yj+8D4FnJI9adjbFOug2hicpo3QHaDMq2ZdqcT7z7qfMKwbhFwuDC9I7y25YLsg2aAD7Do8kPZIz
+mcKf4ZEMU4dYb4Fg4SXPTmTAff6EqZuRMKj8k8VLPhCMTe7en1vDZg9fUatX3tIcfhz2iHkB0zO
3Jzy963d1ln+mBKRBAiIkp2OdhclpAf5GbmgRBPMiHHvQ1Sphwt/Gfmc3Jmev36Aficeg5Ig7B8/
cAa9WH8tQfLyyKngvIRXpihi9ea3LwqncMIuO8WJ2DgdJFH7b6Y7Sa+AWwxs5Jqs+CxPt9M2DiEz
FbpU7rf9wXGw22px4ZpWMCckZP8NEaw0jazu/SJZkcTYqB9duBy35n4VWLMsb2rsLS4i2u7jQToq
P1hO0ByLO8lOvz43CIgc64u91G7vbTaFWd+HWf8CyFwuOlVBARN9uPSPMRMqtJR88bKNpFmaTZwL
N0P0syJxM7o9wWCcOGQzDgbDpMSc9oKaOCtlViAtkG97RtDXlA1aV9wJ+PWYMGIYeKWz+AHquoQ4
T70Rcj6Qj8a6Cf6BhrcfcErmhXLvajsRL9gtdMHzr4c8fb/utCvTg4tdmiJP0M5Mp2XcQ67o1TD1
t6/tAo+lufsi1cDUvGgB1FloIJcr9OM4P6dZ93owlqfwvcQKNm0NPuphCDM1HTREUH40MxM5aXDs
HxfMH6quoOAera2asvuanrlv1imCCTDYMpGqno/5ccuB+h7OYG3QRNj6wcghXvndZcl0a1TifJLo
x78J6QR0m/PmVaaUiJUJJrom379eWZjPUL4STICC7pFmva8sf4rslDk2Os8HjHpiqW3E+J1fDGp3
mVB9e4J6fsxObNqZYNHqSuLrzmhS6YFcEwXk10kav0IQZ2iCJ+fr/BEj/UdFOpwbMea8NpJmvyqu
VRsGIKX0MNV3fJdQF47e5Ato+/qvvud71k8is48tr0MkELX1lcNhaJyGx26tR4LIQA7ML8vpkvtP
RUGuR/CPS8TDajujJfs1JgYp0tz71fuk6/k80S0IWrP7KoB79pTYwAzHhPn2w4ptfHmkWPkbUnEn
ifsL3kAXexJe+h9XepwxkDWeYwOaTqbZNh4+sv2JhxcvhoNRsG5fjHFPQVX0fcfGLcMyQVTK7AVg
JwpwuGEhq2Gsotub2XD2Lw3voVRp6hDTK5rBn8RIUNtNwxi0Uv6oqab1HTa2i2uwT8maiSnCuseS
vlbQ+4Nms28oOtfTrltEP0emziStPlywsjgASPPNT1nVWsMJPLYci5tzV1ZOCCfqua/dWc7kSe4u
a4vlByuF2L0kTCVPz6BchGIPL1ldmi23reXSlkpaUimUaqK57BJxVzSvdLz7TWmcHxHrPsI9e+xe
3mMb6mWIFaRf2QISR7i6Um9Wgh15yqi0xwm2Z08j2I7sfftY3jc0Wtbilpn+L3o8IM8u4G0431GA
BKiK/v+SRcntYy7Umsq0jJQd99qCCA/Jf77yFYBOVWw+1XEB2UtoY5oAMMW4vZ1LMsUc+9w+hEAl
XFYgnl+ITNBhqXEbqdEqtTB0smAtALeBY69pqOeXjKoNM++XwxhJWNTW7OoLN1BeHQxgvAewsAeq
qRkiAZLiGjaa7iToIUiNRqRD1LlpBy3vb6A4bmK7ZXj4u18kgz8Kk4Cd1ayoy1vh6gbY6PTm5Hdx
kKexTJGbhG183QFp6okrRtoAvqS4D6OWrHX1nX+8FJ6XC8+ILmrqb80sTRKpzUgKs7sOK5fQQC45
8vEBS9AcidvNqwcrQ/eQkeerA5CXp+cZAPuGRXC4WUeFSEChrg2Vn394kUYeZUeldKjFfNpW9kdv
kwr414+DyIUOb/p7he9c31LR+KW1WYYzjgfXW8jJHHN6G5kWiKawpLLrrBVpRcsQGXQ1RdzEFc54
ozo0nsIr3810NJhSyzmBmbd1Pu5xiW2DptMUN07YceyAEdQ+DTW7l+PlT44vEs7pZUiLOYst65eo
PK/av4y6Y50jAbWE5UL3Eg73f9qhXZcYzirpYanTbT6khfHA3mWSoEavrv7TZt0VZCEIE7I5E3dG
uDWYXSXCEk+8JoNs/vOiv5Pp90/wrpOeqI2HIb3KJFIi5pJ+Tgoilp4Y4x/zLmABx/Y0JtS5MlQC
EKCrkgvnErZbPBHBZbMDegG2bIR22D7Q2ITRla9Xgq5tklKwiUtbe+uhC88O4KwO1Jb4jJcwdwfW
qFZaOSxCNc4CDXssXZDY/BJq7Hae8Qh01zEMJHrYABusHHZfNbxDzWgkKOmF7ZPakHzxd7dz55Ni
Zhj67/6hRbEWcwM4mRHQrPEwPTB8541nME8BniCw83HhD/CXwLftD1RBps30Wl0x5JB+D1wf2aP8
BjTpRohSsK+TrRVDcMQhZQMEzFNkPcas3CZHyJiDxjRzaotaSXi6DEdOO8eGukh/Cs3Hu8/ARmSi
lOmNJJ/QhefNc18YWH7Hp8DKJQqYccLXy+7gXhb/LzhqnKrZhkEqCihUEGZzHQLXsMfHwHvnXiLA
iG78i2PHAkAC9Skv0043wWK9rzkwwkfNKusifMlFHCjXihohcLSw+QBE32MPiTPgabahyu6A+5pa
pQlu+ItRJVpQmz5jMRqknCLq4bT+T/2GBu6HXmxvEPBjaZp9IBDe1l1aOq7VqJMeZg4cv3YlGkCa
PIxAeD7sFUuoN3gkhKD76MUPKIWtOW4qeYVjK86M1V0k8q1SbSwJjOE+lCvkey8TyUY+fdwpVDnH
JjAs1uBRoN0PSPkBvIkXvurPmSjQDt6+dVrCOXwv2MtRzesKv8V0oSHTUQS0Oia26E1bUAvy4Fzi
2vQ1ToOAJOJfccLP5iT0RMvgDUKOhmoJwqG6vVfrQsZjW1ZdEzOC0IHgwyZXYOOfXjNZX67rXPU6
5x4t2KpKXgHduuiAV5xITs5TUuw3wDC5L7dkFeyRlNvBrUUT7wVkPAE8itWO9G8ed3JbBKIVUyT2
+AbluP3/ruZW0Y/iKSyw0uvIBvVmtQi+N8cZ+hdyH2qa+4RpEEmJTdI/nLQZoWWJ7Sb3RqPMGqyg
1BiMZdm2n+7B6ALodwirVF8886Xt5QUnDUUP0dOyrI+m/ERneTrmttT7Z1QYeKICEISi8fGVEaKN
VGxHAPWk9jxlS4VfFQco+ZFjmGKa0fE6LNseGjuKIkFUNGYc0qTr2EgFvvuEnYfG0FkxIGPrCsnZ
jIut96eYs5lnXNDMhr6KMKl9gW30p9uqOrzK/V/gF35MJh/MvqyEg/qifBWWtgIzGYQjtsD4Wsvi
E1iBGCMRz9cLneBdKYMB104VCDKrEi76RZn165z3FMsMFqQ4D++0d6rJKpPNx+tM4yx36ivUojhf
JMLiejz9T1lQxlNQisVW1+mgRLnR1/ERDXE+WiXFSirtfJP0Lj2TAhml55xjZMLBTd8Zo3TCc+Nc
/18QOkDRMz42m6Bw5sxkj8qw6Htlp6RYiLemRLTU51F/qaikChqbpqVXLQwPYa0lH4HavKPoIrvz
GC59gtjv+bzht1ESNyBt0l6PaouRictt67x92xLyn9dGvIU0L6twXB2qTKNoH6ftPaKaXaMKpcXz
BbSq7xvF7wL23tws41kmb+0L3M+Ncj4dFi8i6P4LVmvaIVXHFBERIh7X/jZkGJJ2UsrV78Hto7CQ
kiWZzSfSrP6xC+ktYI0+BU9bmxd0eUNSz++xhwJ1QNNIcgNWdzZU+XYGbduZFfVUs/+FyB+Z0Pd5
Bz0GS1gp/6LuQ8ER0rD7306K6FG7u5rHznJl9PcGcu2ZHH9DnprSSC6AhI7DDWJS58ZpRYMp6myZ
5EKlk9Rh/9N0qtDg8fTJiPQQaJz0SVn0qVwWOawhY7qQ5eZG5gYP/QsCACDAqfg2xlOXP/6q+wAj
7z1CihzYxBwaKqU0zAzXER4x7CFixwDjUm11fHXKwQH9PLT4cMuakA0EdG/SCM6p3qaM+WF3ahml
W9eFEr1jVgjrGLNfdmiMMGJ8zuwMw1fkM8W4J/opy9I94Kns067mJAMvZE5U1xh9ZIH2SdVXZbH5
k2+458BdGhVubtk9TLzvRVQlM6we7Rzp77jC402f+3oTJNFX5GNlU6OR0Q+QFjuIRfMUWIAORJBJ
2bWD66UleWrzaIIHEdDhvnnHIUmFrJ6wqG7a+p4//MlatYJKDrw/hmsURj/GwUyCMgFIv7H6YSob
VeFGp3noynWDEPSJU4qStrk2GOf87qdd1HTmVR19f+mKpdKt/8jsmUmbmqn0u4SspPEWo9A55NS/
SJ9HiQ+FiJUXMyUEytODJJogMM95HXLvura2r4RcLXBz7+iY4jIHkG0zOWc8aB30SaeyRwpKrFBp
1hU0x1rNqTnwA1DEFGxssi8BuuqVNyyXdYqjUVbVyA2J54wHuKoModrUZ7US4YjBLBvLNKGme8Zu
UDsj6zdV5yn0WGB0fgT388D2Eazhoj9BFWVkBdDfWmoMg8SaU/ykRMRbKiwOkZ9RbKndlonev6r/
0yS0O5bU2cnIK+mTKMnJSqj+XC0CGsZexOTbXG+kUCY4DINuGMahl9nFhQHkrZGVWnyjZtuIgc2Y
/9qhFFU230+xmsjTqo11Ql8GaM2DOZfn7SJzq63hNmIDro8z+Pe/0OPf3g4DZ3XqHRhSBjG0AQUN
GVibkMTM/k3tKd2esGpeKw0JZV89R3xaWZAgy4EnvVHAh/M+sruLdCGtfKiF2NUbpTHi1ispkJK+
TxMpbQiyMD+sfKtWruS10ZFHjLD8Rgt7b45gd+8K+blbaOzPw+e+2E86auPhv8+Vrqp8TCsaBCcb
syihlJ1x1NA7Ev3FQ258gwOPmxz7kAXlez9XKaAPV3PCfwksHUqS9d+TNipwHlQ9eqedO1B9QkSD
ocaae/7jdhGpKa9ctGgSrh0aiMljpd+rZ/eBx3t70MPdHTiZIFgdjRRDQmLWc0z+W12CE3odpSFr
ZCeNMCb4f/pJftqYWMbac+IFSBdDrTYiUoeBtyddPi/jJF7SGYvXFQQdR9rbOicnfgY2ImrZG+U9
RzS5aYKAM+PdLgvblqg97c0DxibrubYD7wfF5JyTHyalSQemCogEDf0N7N9ZSLEzX4YtdAz0SkdN
HWd7QaQdA1lYLSaxA3feBrkt/2gMy3Q7r+d/8pfHSXmx2LKLoeHYurMa47ZaWxg+gsUg38RSOSJA
ryK9bK9oI79QITM7VbMvZUU6meFwzXPMY+0BHKVYghW6ZNj7nm1+599hJ4YtL3FsZaair0T02nF9
nOrM+XN3dI8wm6PnE/bmSywyBB/pvi+kFBINqFXGUO1Wig72wHEc0NwpstzDuMerqTY5RJxLZOiJ
UH8LG9rKNRLv+aPI9Jtf006rQ8anv3vWBTxtdD6uaOkyejY0T5CDZ1I2HeiDIhB5qBFRih4LYka3
dhde4hTeSV8ctQyC5a10e3Mw9Gr6LNNGNTNFyFI2F6LFC09P1ChbaaketvE2ziXb+vSpzmR9KpbI
+CZmfuml0AHeyP4VhcW6wTcDAgfye4GAhHVraA10Jwu545e7Rl9vr8WxSzhmYwdZRcjQ47lsWQPU
VCjdjRJbd8p2dlPO8tpU0jQHY9i6hf5nudm5BXjsXnMyu1lgN9kq+XaasMbVRpAkrvGg6sLO/9Sd
BO/ij4if9n05/wwggVmFMnuYxJtFoJDLmyXAmM1/qrChriMpIBa7u5yFaW6XndWHkd5JAcv0quHp
LsPgpfyqnErhkqk1l3IhJviSR4r6anv+8rje7dNkiSn9EAjBECkUiVYv/Dn8HLO8NaiVUwWTgS57
vE4rrrDb9s6T98n24nQzdDWYbw7AtQM7Whhdpy6DGUoraBAqihPuqv1PJltUXtUqgtcLe/LQcA7w
iNTAvmXXm6eiiQwAuMUCrtZpxurz6lO3DI0lyJhDy9yk9EAwXA9y4PgEGYeu0HutcgDoPMKPcGti
6rrvpnDHNPBxVNVTM0lVjvwdscGKXQFqcpMfzrrgsBkvlqy4pp9fbKnfeKpeK9TZS/1ohlJL1m5f
RKQbPsumvwyOrJOMXSYEyG199IQG5spXaXUc27e4V37I5RyhZXV6oT2Wbe1ASH/KI+Rij7S5JVvx
2T/nxhxGpkoSUKkRWnU9NH4rnXMiuPKQKbCipc7r72EFDvHmiuPW2Q+Atpg9eIwLxYJdkgLG7cGS
B/1buCzAjC58sVsFXz5L57Y63rubB9xAFS9EhDjZv6/G1qsL0koVC31TmEyHqSYabQV3Hb/cfrZh
U2XCHwPHnSU7WHYSpGSE5EBLLmtElD8fK0RjknyHpQp290AZR6IdSYUnPevM9vdf4e23raKaEprW
/Mz4q+XVlZm0Rn+ffbMINFErfUEzXsjJ3/68REwu7i4FgoZc1ZdKq635i62vofVRy55wy8BmcQMG
N3mh/4r62mcqq69+0CHWWII/RL51fSEJ9VWAErcKtW0vrk/Ik6pkzNbmkk1eQla+1GXuMZanmhb8
mwtBTMSng/RIbCosjybGjzs3Lky+sZLuT6UZ8W5sLRatQao5s5sccvj+c6A4RcC1uaf9r2cRfXXb
pc08doSWvWXOkF23OicR2vShwTZueg1RSSvKTTVY7beA2B/QITXV31nzkdzjdzuZID1xVInQokQW
5yFYxfVGTnewRMj7YZwKI1uHSZWBElatz8XgRXvNbFj1CQ4vphTCTJlUVIS2Ump8QFZMAFedxJ2P
7QRkhy/F45uvzFtRDJjJ5K3ZfUU8RdZkStwCrrDiMfULaSt229+EphkzztlYPO6JJ2u45wrhg5lI
GLp6pqM5GTuBjDD/Cuxy11VHiajG6ykV1QV0fT21xBDJtPaWYllYBLL0Om7Dalkvb7vcOxx5ietD
EpdiRRQsuPM4PIwTKZIxVnE4VcG24h0JMeRycCG7lUaCe9MFGivYJMH7RHMqyo8sdlLsPqkDerNl
jUME4To7ALz23QVe8B33+olM4bLZUEfdp4XIF5KYzIw0AABZni0JqGBtP5opTiEANeFs9TvAoTip
b2Kj+T4LldyJAzC/MZ/CaIcUdxqHjuWbCJWNi4H8HI/8m4C9zrDjssjgb/8AEX2aKdFLOc4eRCCE
9PWf7xLM3atIJQ4UZVkp78r1AX/+2GtZReUEf5mM99dZ4keNCyjsm4qms45BzxFc0NbCHSH694Nh
0AEWbTufX6CuL/o2j4PI6wc/hWwxb6FchrUNkYHPSqTMP4YCkY79l5JeS9Bx1uEGzrD52Tt9IbMN
sKFS+tlYk1oa2bloRKxqGoh5nu0qr819d9GypySnLDmugy6le80ttgJz9X5CRWvh7eRI/er1zUg2
Qgg/uYZF5Lcxt101PJI1SV4Wc2gt3ZBWCLKOaWEhSaXPegY/lzz4yjKUkd5UNZzdVogI0CLj29Xo
S+leZfD11KEhts3euoeylK0xC2MYV5QcMhRp3nCpTflHDNq4g58xSbtzV92lHJxs4sPWanctEbAn
P2JmibtK+dfwo3HhWGErKWUEWLNhSS920v6DsOQGJAYE+Ra/RW1ELdeBaCiUAgmzSs1XYDJgcBki
gUYeqo2tQyYMpv3a+fKrABYE2hfOOB1uw2tFwb4zjyVNoN8Ea3zre0/Ji2mG0ctHAFdZYk2q89fG
TI5GPcdeDMxo7cMi73rrobcs6Rxi6YjX9yCwG00cSlQsoguOV8lRaQ4nr/nNyZjTplyX5Ij/+DjY
1TXnD78YXLqYf7+fMcvft695byrhydvUEwcuubqrs+x2F02Ix1QJADT92Ayme9JA7zEnN+oYH2q9
TyNsnqflqXloy2D/c5Dg5tm/OfbjhdeFB6sa3+biNtY4QCdNFXfyBGqOKR/qhKPFtF7FWh3Gex5r
VM3+Eax6FM10Ll4GWqKIKSzlPgN3ZzsvDjMHErbnVar9i85gfUV2a2ArHl2dnX2GkeoR1D4+podl
dlq4m+/QtmnYtNIl1+W9EtOV4VQ/bJzKhdxVZGwpXEjSbg+3pDQ8bdanjftiyPZ1n9vTpXq7wQj1
iwcPkbkT/qyXQ9O4YEgrfI591dS17m3mNgnYLssAiZVcLr1pFMhgtZWKyXrxcZlv73CpHU7ZsSDi
U+IC63fEW4CPXgItCyzhs80ZqgYjb9OP7N/94a6oAMjZjiZ1slOWsSPYcGimKQ6nnfUIx38Q4cg+
sXGktbA8gnHrCzQLeNtCk6DfBbCALqToDRPYPsJTw4QpdyuK3xTCFlwW+9ya6OssGpzg+soSVH0D
kmf4tOUBynX777w+wiBqrQQSBMAtdJi//A5f1EbgqYQlSLzDo0xKxOM8M/q/28KiDMGUoz8+/ghr
xh3MC+SsdyrPfB5gCaWER6CZvHo3jdYXbzLzyr4WPDeoFMPmERIQEs6XiqFEsPOatgNoQrJ2+Z9E
y/yQywAw2KY5G/IXNYIrui7mVyzmIKyQS/8l0yfryMGuwVpwpF+N+V2MDuP8x2PZeimxbMeEKW5S
drtV18GE+NG/2W+bWafBCN/XMOwApzEeQ39PeUNHy55zXGSmvfBpHkiJGxseAWsKQNdrMaFK8KtO
Lh2IO1Zpe7mvoePnGeFYyreqvu2epauKLqZ27p6zIXoivBxP5hVWKo+9z9Tii6sK6qf8W+7a79D8
Q4xgKeUDIttHlONKO/wa30cgKtOzfPDUde7AHzeX2VyusjtfSD8VJPm1eAXbT+zQAm8Hrm5pngwO
1XPYxSBk9fqawh8wzsEOoj8N1vRFCCVIWb8QUL/Tnm8M550+72yJNmNL8GjEOxM/gdxNIZTkirF7
lhUzi71+P4sbPP9kGtpo/lt1Z5kEehdojw2BGjeX9Y26YBUJcDhQ/znnLU7FdNmIs1Pl5brPTTaq
hfeKg5ZzxOVgx6u+FRAI5zugPmqL1tvCSMEYwBppK3boFrg+dgyQSRkeKOCTdGwBLNfF25ODp6cp
lhqa+y72ctE++0iVYupA1AGKNjMUN4CAsc5r8nZFULb5Cmg0LKM1NYbGius6bdcppXQcNoymMFgd
vBf4p47tF6oLWJ7cTJ/Xf3wBmP/0DW/9bCu/7raSQNG2e9z3otncy+OQA8uQPy3bfmqBsA5JRBaQ
JhQE1mRVyhU4xpoAJyJ//imVGND5Qq1LecGMu0n3niPttjdyIjDQczQ99gy9UV5/1L78wLVMP+fc
ByFfzev7+EC3UIL4MPhtE2AAgUwg6aWqq6jg284WcQXvWaNQXkJ7z5JePkoLy+gxVuJKx14ers2D
dqy5I5BbalKwLfgiEyHuaWciTuA9porb1TX/ol6Z35dGSBg/w7PhxlYK0ElovmUSImJokD6qUrVn
8DYFVpM/tJuD3nsKBalho2/qxkWVCyTMLTmBTNKbC5yuefCj+rgG9VP9DoZggL8GDSO9Q1sOKuGZ
KRRMLAFSK7Mhhqcl8CdxxZVTmVkByoef8TAmbJcDUMwMNfmYeb5zOvx4tecXGlAqs/8MBmELbbM5
gJ37SVjtNYa305OjQuhoiH5OK+W2M0oaeSLQ6D74larq2b2a0439SXUkj4TQU28NHo+9sUnnUksH
LTDQ8eF+D5vy6yFXq9pdAOJ7fa3ufxLwn3TgGoyyEwLgUtPsoTCCxYFZZZSSYVlBrfRCy8D4JJUn
29BmNs9TFrM6IZAhRiWzEz/x+u6Xkqs8nG3wD5TxZzd/IqdJcSjIDZ0K4OEdFINkiFLGaMXe41Jk
a78dWcYRQ5JMNOuFxuZbLIgIkoibwi6fSJzVzTGdews2LrXzlPDO2kyMnVropUdSvfWU97H9sG8U
8t2cGfHIyw1YTJBqJhDEhFe8kVLcMFs74KnEu74hWWLywBWHwyqTQ/E60kooDsdJEAezswHHIndq
d2pe/GsSYv4KfMlmhLLHLT22ABbBgsgUSexA8BIPnwWPb1pn6swyKcFcvkz/ewGb4Kit8FA6i/zn
xftdFt/5SGdlxGd1wr2GWnd8FWbS0bvkwm5j5VsyUT+gWYse/EFHmDUIB/4aO19f09VxQrW9QiKE
AyFPFig8sNzW1OLj4vCSV2fkVd7v0HeBrhjhbRu3/bmKrQeAKuo1Aboyl3U2MWb8Dv1XRVHMGzKk
m+BDqK+kSgCv/sLYJBLimANASZsSgpILZ1SNK7GDGWFmdI1TSrRQWZW+4yYXkxSA2kx592ZsDOkM
e1YbU8+gOrgCnu78Za6VITXnVBvZQ08x7uvp71qISi1dwjimpHoRB0FtooB1xm+V4Q6xyhPcxlrV
s58k8rvFUIauiK6C854BoyPDwgV+gbur7Ac2H/0TY10KyhXmV+BrcpeI3hSP5Z/1osUZHiYcRJAW
+sEjsgpETXdKu2lyaChVxzrqQL4FIDpmBxaQwKwY0Zu8nZH5r+yGom8vwBVJppv0DC8lYc/h5zmQ
viaFJ55/aCha9aDZyxUUcF5d91RnjLSxBUXxEmjaBV4rP4e/iQvbRX3UZ6CE8r2+wKinqvReHTa1
aJa+0sR1P7Fhmkyl4E4TN2+9NzjcQo36zSLyfRWhS/NZv3zt+Zj4oItyen4rQXOe4poCH5oWYb/P
p9oAQDjBMeY/xIknJ1sP5BohkupTmHDyzO5r75Im6QLerlfgqrfYKzOkTUQyJFIMCJugmoIZE5uU
65TRG9AlArbG44RDcsrAZXOeynkTz4/HTE628ZIRWE6z4YoAAnRDbpJ4DejsB0fjDqW5T7YjLB1P
KgyCz2S7RJKvaEyNakegelSrzPPEAnPSj0tXwovfo4NLbDtb6Mp3MR6nL58Zot/wfEIIHqvWSLRU
LjKl5nwoH+Ebdi1wgE2ZXmlF9TKYvtpkQXAThxzDqL0nbepchPZmxHv36gTDdSoM7JBmOc6zULxd
pvXdhOGcQWnoXuaRaUvm8vkWIaeWPRIplxFXgjrjZChQu7fQPH4VNTexCnSRoPOsPs4JedDaue7k
IyJ3BZxWjpqmdds0VkyGMhW055yhMVYYmI2K2PSmihLjGC/yZE6xXo1iUAw9iwPxFazEqSyEYNth
+4C69zTPICO0g6LcCnVn6RhFUzymi3MWErNQtzCU05gCqnzucmtx+ngKVGZJEp2wAPCGvrDCqLOl
65QfvdUH/OjdjD74rebkjpWoY9POI5S9qQ8ct5BqzakbDHg1Uz3juEShlvoX+1zPITYeV/n/VqDW
jRONlkv0GGaa6FGLbTbMx/V/ILClqQQFHmVYdD4dI3nGoGpD02eoe018jbHaIcxjExeZ3+oUFb2O
4Smadw/aqE6nVMS5HlA3WLivGhu6QHfXMqFMX7H7/r7A49j9Bhvzim4oq6rJe4ZsOCYYY+Cw/FMJ
MN2weoULDqxqWtZutMO1QAHdC/aR2y3fJLjwyjoA0p/3p807eTsyFr5jqOi6tw2qAJbsDtBdQD/7
TStlLlbm6jCRFwNr9ATvFePG/HKJ/JISe8FXJtYUwd0dpaU4CH6OR1S6ejjUaaFXngDnN684R0CW
Rk8g6l1g2yBnjGgRnlFOXHxoKNEFmmHiha6j4glK+PC5eWLoX3wTb4Z6xdfe38GZA7gPDtfNxspn
6Dma++Qnay+kmVQBdDgslT76qrpWtWjKmUJ7w84z5XVqDn06BhbBGzqaXcSgDipJf/EDlSx4RYhu
XbCYlj5nMxKhBv6wrtimboBCoUAocZJnYfe9KboD3KzefJ3OLYXdfc9Rcma4MmxhbfcB+wChiMt0
bTUXuIZnQNR0oylbjXRBoBvw/vwN0ZRMgkJqRh124Qx2TOWAM51QF2Q1m5HTqPNe/VjJSn3fRFmw
KaxP1xqz1bYvA68vN6RdGGzFaFISkvng60GQRsbqE0Y1UF4fa8wUJb2A4g8lnJaGeRagDgYSfT5p
dr1MA/B5criFwQ0Yh2fkzvsXxnyqgoOr+r9FRyCiH0k+aXDSBhBZUlVoIWoKCe0q3QRA87ibuvbB
7T0uPdAL8xsPelo7uQEUnseK2hUZY4aN0S7wumCB02UnE+if/mJxIHb2aN/w4X7qk9pXpkpAOEuu
F6rh+3ahVsBl1YxuEYBkvT/TmPJJvi+Q68u1A1nBGPRvp4c5aHifK1OBLK8nHZZUWvyhJi2h2XQP
Uj09MXx/xBazxVuSI51onKCiBZWtJ35XbFZWThxTzceK2Mp0Q1pkEpI479O2I42DpA9Es/mYsg+D
j/q12pThhVegz8Bsq4JBATXoMea+htePLP8AdXNAX6AeWhAIwGtDbrZZYungdjaniDsvUe4jflm8
vsPDcg1ILPnQwZyEO6noUPB+Vjjs4dK/oaKEOjx2SSD2Cw2yYI0117M1Ouib06+Z/4LXLS31fmqu
F7qlbdleNFfG1BwmMtwQDAJfBNGgCAWELG4X+XAa6KhOAqxP1r6E3LjB3t2ek68P6yyQhGHNFN1u
qWFZsx+wcGJUxXGhFUlq+fiVpqDpY74fJsPbBiu61pmk4ouTecRY4ryzg9LgXCHG6cqfnaDT+e5/
xa3/HooZazRCAyiYqfBJ9WPKBcAea0hqyjexeyv5qVaKv7jAecGY5YsFmNTEqLdN5VANLxA9uOat
cDSW8YPSaybXd8z+w7X35bIZhTkYznZZqGlfeuGrMSTAW9rv8TQcYE4+e98PPZDOjrUeGrd3WdZ5
v2pRQbXOY+h+Ur2KB8PnGIq03samVaaSYlV4HbUkwDo61I11nTfDjVl5J+ba1nOZzX2an0obmssR
ExDMO/tIZgxW3mq4zlFskAsGORMvB/uVKw9nhqgcnzIZIt2wCm98LT/Qdxd6ACnlhej2crR2khjW
TfSREkgCRs+aF25N2J6lHhdUqJf89RXW5VUuhBUW2g9W1S/Udnrl6ngmDfU8itP4mneqGA0sMLOe
pNJCvpTiTjiE7UvH3RDf6OIKvuxlH/tao4AlOmuTFvkIswcZ0omFCqFIZV3ZYdOP2RsnnaAJkyBR
fpO1u/MQjDC/35hBIxpXX0o60GS5vy+iElgyfCRkZKcP1mqcSrqxxYEOVivXrZ/U0fRobqGlxYcX
+Ee0x0EPwbet2RAOehdGfeJQXqpyHcSQZU7JCVX5f/rZN7j0k5ks6XfAhcBIqFmSUlwKWgG0q7pg
xPtlbe0zO7lWfHTBmVvHjoXsphGVPUM9Bp+800kApAXlxnuyLVZSmZotY06erOXg319p3VEzPmUT
7cFd0pWYE4lhjvx4cdiEHasjeC1aTjWRhVIoguvle9ZRoV0Uap7zS8zFCJFldetIv45Q+CguvyOO
XXj6CsvBH/2j5Jt0eMMdM5u7V87wGdgwCMmAtffLoLfQD+PU/t2iG/1vNqLqjbemTBNLVHdRIZke
MjecXaHtuC253KLFIZ6F34uPlzpgcADbN50nK3FT+Zra7sKSaN7nm7GbpYG/6eo/9JGqsu6F2NUJ
pKBj+BJe3yzpVqj/PdWlvztOFKEShNzDh1uLPpH6jZOQb7CkMP1flV8cENUGkVJk65uAKoFseFy4
oCLRSAPA2BIsaKiV4vaBWu0ANiJP5FBmmLEa9cj7kiXTF0pkt3OOZjIXDCiND+GorTvZO98WOTJq
gC5ScD1rI2k7CA7t7TDa4wLMvu1C+Iqrm/+O5kGRmMjaNq9Rmv0FhHNn/Mg9cOLLKcrBHUkMlJuu
wy1qBLy804iELLJXHEesbU1LxE0eStf3YwcYmHefnyoZKGu6LufgZIBC/c+Hj7xAGUMV1F1IgJYf
A8oVNWi5H/QBYBAAgi4+4aMOnZsSXBAvO4ONAsFXDgfyzPu0fGOj18HFRVvkd6KUp1LjHk5YtE/a
iDwTqsFakW2rrWHa9sW8VAqmlDcpq35xtHaiwtAas+usD/HbMwpNvz7PAQv9MqfREVmTqdi31P+5
wPvCm/YvPG9/t8mFcZkQQt6CSwXrj18dGav4sh6B0K2/1HIDGYNWscxUJsz1zLq0ud9juWU420BD
Tm2hXmtdEt6Woh98r3reJEWJRGjI7csnpZ4WKbuUL+XPuIsOwChwUHB1V82+0dICeIDKV51G1TUt
FrWsL0bG0ko3AHL2HMb1xUpEvuwDQkV3Niy3Wh7XCKqgzD5q4kCzbPBsplW9nnaPSFDGQVONIdO6
zHdkzMt4GZ8c+eE39K27SDKIGCr5QVtYf1r51KliDNN0N3gCWmUSbG9FEt8M7Vb+rG4ohKsgvWAi
ldu2P8U93e/uwT9t/MHQLMnHaA+olh50j+Ygo0hm/OsYzDogBpmEikaPiYzNc/ZSgNCKjZRY/zMn
fmLV6of6jJI0/Dtpviv3GH8oYClQkqo8R7R4Fk42yk51CL4PjvpYu2yOuNM6S+t8Nvc/b0NM0AMb
jFq8AQXJ/3mL+/WZjhr9Zesvw1onP81EvadtIafRMIICW6H9tV1sFGyNiCCas9W6sRpJCoJX3kSS
t/u2YaITRYGDDV22BOZsC8J/IQrHP99opFw/OmHzACxqfo6+K2nDiRlnFd3bwWD8efhNb6zU2LUy
lE3ETw7aOZinRLprH9WWVhB7SlxBJP84VzcZEBdVl7i7VQE7DkqHNfXitPCN7RgjIEif16v9AJpn
bAJ7ldNqTZ/eGG5SxXMvBCRmxK/24tZ6dBqukOJeC8XYUslmPJ1dsuRDIRem194fjJ5uSrjvgFux
WXbaHzwzhpUQsLSvAnnTfumWZ8N+dj1iQHc2lvPsw59+hgt7WrX6BV53czOWx6mjdgSEb3MTwJTH
jJJNq1H6+QglsNXwe63egIt2sfcZUumRHLvS0tkNf7W4C/xgUmcNbPLmin2NEpeziQr925wxvGYp
3OPAALkS95v2qDF/iFrppsP972qvVPv2yB84nzJMSBc4D3G1jmZMOqVUhahiB4o0yE5WSLtq9X3V
G7HcbO4wn7Iq/gTOJWNCIiL+5wmoGi3vNbrvj2ydyiVWA21rJTLBl0PjJFveiESChkiNukoGFfdI
DzCgKEya1b5+kc58gZvtIRFH4Vr2ySQkMj80ygj29l04aI21ZopVS5zK/XvbIKQO8bF74x0I6nAI
GRFl8nRCESx/6oHk24YIoV1x8NzvVJQNbtW3Oi0Ae9f3Dnf7uaNPnXhtGPQmyO72tOTx0CGpqhR3
/S9DQJ5cl/kLyW1PYFHZtVXXmkWa1f1w7om5tEk6sGt0BrVbuml4qelYZoM53K153S0SLA5x+Lbw
psdvDokXr83KSPalGBo485qEtOnHiVHOCNJEQ1dYX50aMxyyrpLmvakncT89jIaGc1Tl5RMbq06T
HjK4ZR8IaOfz/srmXWoVC+XLZgVVVfrggSQZiWasVXCI6EvNi3qaDcusWQ0UxmfvpzMyt8m7irdn
bp2iNwPm4HlJa7vVpI+wytRRO5PVa8cxnjeVqDeo86nNuc03oU26Zt1dy5xnS+0TKoXDsiHXR2m5
P00cbNXdwYA5JCXL6sdK1cKfcgw3FbdbPQkKpCzb+YPPV1g3236elKqRxhLfUSu2IuAOzehIMspH
7HbJBgVrJ+6vgfRVX0B2n/pkHxqHZyAz9NuunP+byO/FS4PBxl0EJCFZi6QOnwbXzcE+9UeALiUt
6l8Aw4Me3y1DQm7FTqkQwbQTV/BpSTHaKzT3ceYdK+p+unDXDW8gXwJIlCGwrXZZBD/XWACZTogW
rGlLXT3Jw67RpUYfNNWpkRnapqX/cdWv0tB+TzJU8FirqjeXnnabVLs1AoIZqUDapwZFspZLVVrO
n7P1HO90PN1cz0vpFAs+TfFHbOXthHF+ur4rKP1HwaH0ESmwZmzYrtxavzYGRspJg464ryFrvPGm
f6W0rGnaJAg0C1AMe08NST+lW7wJCaGkgDFvVaK6ef+LJgPtoTnSWSIvcFQkbZGQFssDy3BuXthv
Cd/+wccJkJPqZmNxFm9L2XMR/h21F8U+24Pv6OP2Tc4pZkbeFZPfl+C73rmPQ02sT+YLcz2+1BIn
HNb1pLw2+0temZb9ReO3LCeiuehRN8jSeQSMVgt0EGKUDzWV9c+JT+U0svKVlIwkWLuoNuhzWq7e
eMGPGxrohRImEXTfglGl3H4KuYqvle7A+PveR+3mkM35wo0kOzYg4YY+gVznr9Y4aB0LuENOh5Rc
l+KPwmi66XZ++3ZmiYr8kw1pfkNd9332U6O4KkirkkpaUkYUCgzg4aCB4rtZ4oXLfwoTKUVe4zcP
ouudMrg92MdwQuGIj23Mi0mF4sB+AAhKDPsCj0b0lKcHkn+me6kEBW0ARqs870BLQl0PIiNUXRXY
W26Iik/O6GT6Q+AitDlnXGxStA/KrSExyI0yTm7puPsAfAf0P6/E7rC/mNUeEU9hqq9WasG+VFGL
pK76n5KFCwfLC8WLVKOgLWBy1ygZ3ZlnAwTX21vmD40Oj469spRjmFCh0c8HuBy2aIfF6FSDeUHV
0KvrpqBAX1euSJgDxEa7Sok51aMDMjAAa6TFUeDFz2BU/k5H/pirhy7UvB1AGFULNZpgt5iMHNsO
Ps/2LkxxDwdpx7Aj53yri48O0vglkP4MVS8Oe5o8uhlx2b2206iR7wQnaGQ+Zs6P5Uj6qOj20RNi
1MF7gLXfV7Df7aStNF1rSnoIrQO9qv/4QrTHJpSyIQirbaQs4BC4wjmbtSJmSUBqQlnYE4PDqxMh
2oypz2oh6QHC0S8RCjmlWZMBKj7yAgSfiX5PD1Y8myn+jwOBJAz4s+IDMI+7ZMgvWKdFlo9dvj7x
iv1QmvzsXbxGbv3ACokCQ182aSj0+LunrJHpXEPoUcorUPyDCQRm4MQkQWx9MD/CFbEm7csHaXVw
d3AefZMPP5HVhLsz9BcKQumNEyo8VPcnmHz0FO+ep1mAqT1KqTprKFDqeCBJFA3AMYEs1MpBuWfO
2AHmXY7CI4qd8yqrAcunBX+yR6w1h7kLtJ7/FosTnJboti3L7IIAGBeRfjZKnMHrQ18JweZAIaTb
p1B86Cp71Z1YL0zU+vGwmNZU5CMJNyoZIvr8xb1m5hwiqFJ91Fnjn5DvLI0FC9ZyUCLrRGC1QGdV
sia4wA263lQb56zfbbUkDIcFbPBcTJy7JtPkVODMgObLL9VWS9wjmU69lXpsdZBu5tAQxRYrIsEX
joN6AMMa9fFMBGQWJdBtcxl5PG8wyBuzZqIEQ85b/tDLU2vBzA7A95bR9KvGTl1y4EI0E8E4b9G8
Y3zetk8TInAtuKyHRpY7PPDvJKDuvil8PbD8v/l25u6Jz2/PqSTzVNYI64PqYVM78gN9HJFEpG3l
gD3huPQeW49ef9nMCkH1XlNuRJ+1FLDRpECmWb8htuCD2mfgRIiV+5ff0klhdtLeDLzra2vaKf4y
5Zilssb9+kRx0EGqqsIfzLg1tFSrD2T0XEk5/ouVOjasKFXy8SZ+ny9699kg2JOf7WT2fBpKcaMV
dKLy+Hyoggc75AKj4kBtgqeT4vfPIl/+7gHSjRxrFWUbCX4kO3z0t/O1GompoVF0/jcaeFI8f72H
+I4joJOvop2zpYxqbBaJ3uERlaMPEgyOpDhcrTBhutBOydDoVUChy5lhNGszCILeTELGdWzf9AXI
Pkl+4V81owaTu0bH9iz8KRSiWq+9z12X8haTtWS2wlGf5IC/O/VukQ9SssDwEmpSk2GHLpFh3Yf+
gC62+yaedrp5g2VtzSZ/BjQiBiiDifZpu024rknJ9szjslx/Nlli5UG1hKHagftU1TJBlxBgPtGD
82DFgH48rzT4fBE6YW0DXCXHd7S5PhdQb4vNjZYaHRNKlE0OZpuTKp7vWjXKwJtUZER/xVuuVz3m
luoFm2ZC3bn1sHjZ7TvTaMwHuo4723mQY5FcprT0zE8Kf+IvCXWBwCiSsmyTarFkrjam73SgtBdE
FMv4azoFEm1XLrodkKXUPZQMbMQ3phId22JIIu7IQuX4eR4ceKhlT3qCh/98LPcjXw32kboRZYEt
XVgFluFkx6M8blBgVyyVbALfKVMWVdrFZ0orxnkewiz9uZaRmLgy1ut8titbNgoEqeI31LbyDOX/
mXGxEKCN0ag2fuPoKKgwOm3CuQZeN7EtG4CC5AstiQ6U/Q6wH/EcwQqoO3ymI2b47jQAgYLl2cS5
UGFwADbJr+M07pPBknYzcfA5FdcjmWbwg7TI6zkeB8Nbs3Fr4aFsg4L8B88lyqXBWbCbvNetEmDZ
du7uYP5PS/4ufC8wm0CMsw6dD+Rb4LCJ86d7Zkh9DC64wh/6HVEOQfEC0zUs8UYu+fNBCi/oFqRH
BiUVYqltY+Va2I2bKZrqvEjw87frzCRY2aSty6k6+khQXK+EFkXzIm7yVXJiBsRa26w0lhgNVK/j
g2QPKQqjq3IBbEtKXqkqJoSpiJorSZGfU4FUMx2YLbqtwVX7WUBGe05SkOVDQP/OtighoZfr0YYd
fC79RCUiElw849gTZYoD9dRGGtuV3Uct4pvl2bZ3dt9i7Z4hJUKTqIbIHvmtvnNyvU496fdqE7O8
4KJtllcJrXL+ilMb+JNAZtrsRlnX3NLpoDu4dJp1A7j623ekHEwY2N2ndK/riBgkc8OyUONf3ZPT
pgCWdXODblRAEA0T9+O3OgJ6gq7xth+Bh3Utrgn043PTpIPcHJyil6n3lEFcuF1wxNlhbDz4QUTH
QCHI1D25TytnKrpHnnvkYHwpLh0Q1QV0dlIyF1qULSTk7DgFCBngZFzRdSDEl1O4t+Iw7HEUdRFS
YxSh8NrQ2AEQi/YQ3gdzwnxkxTdXe6h+eMQ0WOVYWPFy4uT1Y5klHBTMinU5hv2RFhqBScFfbtSM
EVcv047GsS+0/UxJRyPpB73ejYQMo9tju/hF4igdW4Sz0hDAruHBfDD4eVbEtkOUgOLU14Zuir6a
BOciqauJtrrKspt26Xwc45CwTR1wc62dNlCSPi1jWDVu6zBb6iEBZwNFRHqrYZPHH6QaLgUoeAOB
s29HSbUnoVzHHxjSlijFsAMZnEUmfp1B0nGwTBNOWEv/j1D9SoMwbjWGIe+WA3DHoovnDVlP8gFW
n36HURA1mu9VFQhwMOwamod/qWIPYbBdMUpfHTszcwVXJWhHr8Jy8iJPs94LBkcIObcCaG9PPeXM
4JsltXX15IgG60PP78baeKsszp4WKlOqtBDSeKzHizCGAd0GkMuA4gx8Kn4TxrwJw0QsIkVIecv2
gQ2p1lzTckrWD49oIFaivnnArE0f9O9qrp7OnJcBbE7f3Oha/QnDPXX6J2fZUGuoseZ3wi2xOSN6
GbIwRRfEoPOQ5ylCDsLrmm3CbQPlk2BMB0zfnYATS2DGCrDNUKSXI4Seh/SQ5+0EHYkmyJV+ckT8
L51XUDZpPQ9s1oEhG+GkbXG915pL6Fa+XZ49mIOOiksTzzf+HseTsjPDbMNFw+9BKU8bDb7tRVuO
8E6mZgmnwuOmxdAlKAPSZ5Mvg7rJsoh9RE+CE8PFB0cGQK2vrdmZPmJyPkmo2T7b/sdMtyoj/yXt
0esaxZgCIQfY+asuhZvefnDWX9br8Rg7gJZd6UwGIixj+QZIQ63TMbVfIWQElktdlb25RpuLjzQw
oDsanxAjfuZZCN0B1BTTjuG/x0hoOhKiy6rz5nGZaV0Y61mKqeLV08V6onc1tSSLVr+1dX/sb6G8
1uIrErlRVKF3Kv72n7nUZgim8mPa3OaTKVss5rTgkfzhuFGPTaAnGqjy3+NXhOB9R9KV15b6akN1
YzFbydm1GGgu5KXMx9/nP/5tturZIrW44lJ1M0RkH1p8cGkUl1HgoXkAHr+yr1TzKm3Z8QXQn21Q
HcyW3BcemZOPiFKwt0ZebyiLa5+SMe+1j0zwnklRowERAT5I1qKKLCG781ydsie/RUS9B8pcSMjh
ghfs7dSo7S5JvDBalTNzm1ZG581NP1dmp+lBI1EFIz0JhP96yMsjbBUv1cgH1UHYll7GU1MFwR49
a67bDnC0IzifUWH3B2K1LwDevuT6cYCkwgtJZO3hv5FuBpkdsD7WdMfi16WCZfUx7lNxT1jeMjNw
H57NuOoEgpmqebrjcUxPGnoSJY4tq+ErbWiUeMDS69QCS0uYiN3HkwkYEZIph3VGVZ1P44y6yzp2
SAo7lH9CvIY951rD8Uy8xlPcLWICuuxNSmw9hnqmyToZr0tpGxwpj6k2d8PuZxLzP0yyIp8xyV2p
+Uf91CsICLxXBYy6vVTI8OXPKpaul2huLywZwRFx4WxZfnVJU/pOkblGxBVHZNun21QPE1H7VYEG
uoyBpEyklCJSuABKxJz8wJjM3WU3NvW62yJ2VcVzBYYmV/9VfqT1oLiFXNGDID9+Zot8ETRfeNAN
BnAdgVxAG5VjeIzzmbR+iy+2x/bT4eOMOpgESsZXN+AzHnCVUwcpX8BXCXrVwdWq08MFTpLikVGn
LeFGu7l1XAgooKr817KZSVH2R7ZFKfmouATsvceQ3vPFPyakd8cE3h0ZflLaMkKzBU8zGvV6aDPO
366EONlKJx2mHdYjQpH3Dh0gddRUaJ91DPNywfqk0hf3n8pIIPCSyzfwvcsnQ1rqbyC+7tUJ/+Gz
EPzUMHm4B0VC9XAZZgI3sytHa9pnPFYQPm+71u537mDmqRIjMEFizwg8xobCZWKxwCX38SXTTRGo
CHhZjf/rLiJdNzQlqebJ9PqzBrjRMEg1mo5vgCZut7Hy/10Vvt/04gbtdMRdxOeMjHX4jIUP+SFX
IsaUQaGcJVKZUA6QRbFevfqVdelClF5DYKIWUNYMmtahbxLWAvLvWTa3jsctS/ac3VAoAtIA/j4/
eFqeTCKvO/qbibg+g3uhaSknGuemfR2pdDYG9dYf0tJIGnq+dq8unCUfcRK4Z+ry9l3/5XUGFRpj
Bo6+kldEPTjc6es6oc/T/URYgjYktzAqyPkJq2t6SB0eGXCpitCAPzbQRsJQOUP7wT8BT3nz0BQV
cMdL6uJJtPDzFQ8PwjOizIeQqOQyqLusCVFVAutmERlc1LxG8/6ShXwSHIhQxttEag2DdgYl5C4I
h1kq+KVAal4Ndc/Wy2vYKJjG3r5SUVMtRxxaPoZ+FpOlxQK+6ZDHr0rYaisf3TpnTJrYTiQDCD7F
6fl9kuUGfUjy7cm/mYpMHzqAHWsZqGbOVvq6QNKyhJp2/PfwGF+zUzUOg+j31QjA1An/VJ5sAlhc
8jA75TRWHL7Ldmqk06xCk9XMM9qnqvqF71jPoTTLUbrc6JxBapSuHi+TMypNVQB2rtTfcz7Jd41Z
fcFB756Q4xnw4wxLwzstTzggQPb8P71Nzgvprsf/VY4TxN7ia/84XhonQrnKbjIFKhjEyzbf3nXS
cOB4ZF7/nMYRFIqd44JVmGPql+JYuc0ilBCULN6VUSbeLD3/rUaVgmGNvSxcpnh2+bcawxOtmWEc
JCYaNNaUrW+GZGiSSipYX4fr+XkqmBG/5qQKXq9urfpEcdzQEAvJaFrhDqCUfSHKj5p5zMdH4YV0
wNdmqG5xuJrr9aRdsLbouFOECX1UxZ26HhoX80TryB5I2qlfyB8cfVVzGqcu+8rXkIxPWtOA2Edl
mJ+mEce9GCZixo/hFoCv26uNJ7rvf7ChsiXBjV2q+24Bbpkr9OY78pvMFP7qsXXa2wsxgoOiS4Q9
JqH+UxBMV+R/QTMc7reqHngyZm1eDtDRzt1Kq9p7SuWfi0Fb8oYVRJXl3/1NedAYZIi5/AU8xCOa
kasHNLS8CIgj6fvay6XGCITnC8JQFuUMwSJ2Lmlqp3WXD6cYDcR1Jh3jdt0VSu7q+S+HSTtkqEVp
d1OK8udfvW4uCUoy+8+Dp30DgtXXb8VMjROR53OtAeVXJdsD4m1AF/hMROHEmV1bLK1ChSfoKEpB
rQGlfmrf3ia1CroM4zZ5MCSl7LNKBFzWI1CmoW1kuzHmFIG1ZWjjQ4MBr4788BzF96CY+QTwyg7t
JjywpCVlYKgl9cJuZd278MBDwpAemQgoDc36mbdtY0qWC63HfknFchfADh1wL/YccQw2F5xYvBuo
rdPWWs4xPoOlpohi/kQNER/0wae/QGoRSO4gXLxc3sfu74IvP++aFNkU4CZ1xAXWyqIiWTGo+itS
66feJR9gMaGrbGU7YAIOJ00vYMG5gcdTU9ldRyeWxVDPPG281XrapujWAlhr4GRx1Y5/D3Y20Qoj
fcFOj8L7gnmohtu+vSKs995j+xCVnyRpM1f2H3uZCdg270RluLx1ng3u7kPQoEB0G4v8TfW2uGQ/
FtT4s/r6U23qqWj+peUBT5UgLcDeDqunMMxR1gNAuroBR5a7+FiStJLxQXF52QAUwiKZW98na0iU
WZ3kJ6BtVehcPP88lyG2V+PI89RPbqcMNeuwZqC7FKXraIAcpFl9Kmst6QsV2fl639dy9wTiUJg3
py3duPMSPXJUBXYtMqSm+lmt6GwumYEYzi6UljfOzsW0Bhvm095Mo4RA1YP0KVunEm6vs0SD8Udb
oqRy/aMKXRVA3kqwLK57XHK/+BHbiTI5xoT++myS+GjetsX4kBBukQEjZVF4/h64OrKQVOVzkZSS
b2U5FbBraJc/Vi+pkxFPsxoHsiAVkDx69SUeCFX/0oY6nRWGbvzCfMyKqLzPMLgMIijwWb6ZelWi
5ESTzekCEcUELo7KmbAL54E0T3G6joOsc7mR1icZSLGihb562KVJXIXgpJDx5Js3JBGWt9fsDgOv
n1DeQGBnRE7MjWRABPCfHOPA1RC2XAoPGLi15USMIU9YsHt9R/rmlq39pAcpImdrmciPfkxisPs6
OVYWFxOL/MuLwT8M19bCKC36wfAuUN2B1prZ+GW8TxdLw8ODmrKpVtAMThm3ikHjFhKCBCcXjbCX
wIWn9ecy3iFyzO/NXbYNfOL7vMgIahYAnkw0DMlVWuZ3HV7p1I8awUdJ3fCU/y/dmahDmhlt2PyY
YyW5j8AO2Zt3IyJ+9bIhOx8nBaG6uMzPM2hfJ/WEdenIhHYlL68TMxSIeN/2x6+pmq8VX0Udw74j
TYbcYjGt/8AspFdGuwLcmH0wO3yAWdXiLKw85j8NO3bFSLMntdTtS7JEccCQb5dqsc7k1Az71irp
0eTIkh1tPcOZDKO0ItqXG+dHa52DnJacIgOjhBPlEVf7D1dtET3PERD4g4xzFFnP4f4JEiEFLlOM
L0cpQyhQQWQSf19Y0UaQs84COWvh0VFTA5Eq+Gp1ZUZAqPQxgh5I2PGpl9kVOePEiEdO/hVKGajE
d/k/89mjUEKs+L8CVT6vKVJKukDUB6mDFg5pG1ly6fSFY/grz3twNYnET6q2Z/4VBLB5dB6knBF+
3F/+1nNC2UVeM/tOBQON4NqdMvNjIyViPu6OCnDekKqB9OCnQpDIHf6ECTTGbXfcSOZIOKOG+xGf
4Dn+gGJNQ/zP7+Fkmlkl2uE4Mt/VVevkM0N0wCiPPx/DhAqoXhg9TQQfS+vH9W57yZu5L9PiVF/+
4i1WWoDD2tCNDCEKsg/A3+ZJMBL+munEFPhxQSy1Sr+Z94Gio+BsTO3fpS0DJDezgqX16xxA4nLL
GjZl7F6JxHTijCw4P0a1yGRFBmMXZfVaRc1y1a5LBtQzYqHwLMv58DPAmvLWrPCoyxonKmBphrdH
ujppDZjN178eULxBPYQV+485EzZKslRPs7t81UXQUHKp2d18fyljbyVlnkokluQEu2SBDzxpEZ+o
9yyphg8Ak9NNztZUYikrxs2057uKcNSegM3G4Q/O/clIAPHXHCBNd+yZPoGqtExaE3MpQt4y3dms
+ApoI2BLGKq9U+8ia7gbIsP6B/DUTZz/7XO6FpVHEJM2+0jUMby14byFlQ5EeRW/1iz0XYncifHg
bn02/7d2s8olhpphwpzQ0DJhKSKWmhU4bzvyf3c+ZqpXy808Yy2EykE2qE6ZP3BwcZiHBwuBvD65
l7O6nTy8+GGfMXZhFBvE0wEfb8IDl8OFHSjSV6ldKjoQk3gfGP8DpsKGMYY1nF8uhgphXvKlk4Zp
Ui2ccAoHYKAkSM74i2rMB03BUMy8XfmDqtACQjVDFQ/BVWdcDtasr6fyBRtMTuNKnlIWY5YHPMWj
Wuphq85Iyq1goKH9BP8iHOZyGFfe3Bn8VhKvzs0l0c/wc0PCSVSVgE/WcomeJY+tpJQ9H5woDqi4
AjHPzqMWcr8XwAfyxKAihWXhIrcrnyl1NVXDK2Q3SH1QRtWUsJfMLNtI8cP2q1KkcO3hWoK9SKwS
z29c3uvVM7Mk8EXxg/2LDJUYbMAr7qKvySSggCXuqXxo1k1Nz9C/R4JIAftadROs5HC6LdXrCzuf
8GihJR8LBZsT2ie10h2eN1T3njBsKakA6RJUhKbrZDXcpiily9FG892vm68GRkMfDkLzazbLYmgl
jFgmtg0JUEaGEOzZ8Ju3H8NQd9uKlHmHuBpC+swE+ST58CjJgaI4MgztbXpIi/PCeriBs1SxtXv8
z/PWrQo/qRZ5l9cRVu4w1USWIichFspk1fvSxSGjB6uNPtp/A5RySB4nIHruDO1eSt6TipygnZ2x
DuPpk8WuleRQpL01QsvgaYoe3v0al4JXXcxeex281I9AGM3j8s+QKb4ozjCpj5hkbyTheVBBBWWe
TJ+Yf6UqemEqA0xioD7+t2YzfmW+dRtvm1hg3BsdmPtvqvEi7fe3Q7DV5Zt4nhbH0LYn38iPYDoG
5+m94J0E8WD061gwNRZnagjD42sCZ6aG1V/zDWmue7tlLydsNIIR9CPAz6F7A0Y3MTdfAkokwIlZ
7TbGXieaNg4gilBpVolODye92TDCTwUiK2HYlKmSBv5Bm3AVbH0xJYxwfDfJrzzz+WqUpmUEKubW
bndRh2Hv1DoREb+zL/wQ9m/DsCljoXj0QBm56xCEQzRC/rxaulwJGb9MOb8izt6+Krsa5Cy6ovpH
pjzYt2ldsMjlEk1ig0Bb7Mu7bTvXezFmf566YLlRU+oQOn75pgVF2ZCIwnXTj3aK3D4EKlJatnaN
8hQAv23AaK8T07+pWVqlmrifjgMBa1KS7OG8mT77LHadq9MOHIKZE4kZQobxpiL9wpqkMBJAy0Ov
rwg38+coWtEKAezoDlZVeugz56Yqzmk92br2baVO0eHO4zb9QdbKCsPTa2cSYUspXbvZhbXnVR8z
tAX8bPqqAioD3wEfJLUMixk9jw1OUpVTd0pZlSTo06gUqNjwrkOrzBvf2MZ23bTPTrnErlBSLGuq
6BnjUoy1pYMymP1CBS9IgAtnyPM2U9EQpzkEZWtjOO0Jxh1CC6WGL/IVNBD/tlZ3zxaVNyPXnxJN
O1YuWbQ2AV/bd2Ep+aR0l/2LfHvB6oGZjNClOdqbrLf38pre9gGebG+IVP+jISfJ7DV0qlZyZltB
Nuq33v3TsU1NPRnOdtHZCmuBbTYBMygixDWs5CADo/QaUkK/yARwa5d4jt5bYN5mHeRVcLuomqjy
Cs+0WuDXlebjOHqqO7KTm1t8kBXdhAXIIazRrG7y+yQNavcRKn2V1vAKZuM9dtcOZqISi4jfroeg
rdOP19u8mtEzetUSsJHztZUo6F5MibnlpqQTO6p9QHC80eRINJl+oO+VJU+nCCzDj8XAa97ZiB5f
kv+YTyvmbS4TWb/8oS5InyPdlisqll/dN+NG/k6XQeSpIa4Jss+KFRjQpNrpRosnlYfO25OLsO14
9KoMUgNSVIw8kHJF1Lh+uLYDqJ3B/Z8dtCheS62avxyHZpeTYt48lcaNnL2WzF2widAp0abu7VWX
0osLf/sEScJravCjHbyFRYv8Hp1S2dvtl3TZg01qneZU2z4KSsVkZ9MB3m9qUd+eW/Wy68y6p5M3
3EqZ15Rp0NOVVRYRZRwqUiuyOut6LTTTLtwKw6Vmzlxb/S+cUVeQHzW7lti/l198yHJWsvJt/t7G
TRUns2zAyJvdnezUy1l90vQzRk9ZLVSZkyPhihFBIFflnqmxQTKEtoRL7UPYxIbR5lYyjB3QuZkN
6kTUziQyafaLu2+YHtP08emWEgmJqWmmytrIIcd4NnV+tfOW6OLWmnY42fBBnReDKjOBeqADyn5h
0o8vYra7XbuF7PpB/t3r3H9wv2bAMIMQoEqFMxiDQcb2nyvtNOQ0H1A8p1A5C1zvhTwB9LiC4+9l
Ry0vx1fR+eyiM4XeV1ShS2K7oorxw5YTjGVQJypy9kemTnS9FBcvM1UQBXk2nBrn0GAtoqALgeEa
spLclcw/4comKRhInyF9HTfcgFwBHovMeiGHfVqwoJqBk4M9J5LSRXSOimBK+8vnGcQ+I7g50Hfg
FSRDQSwd6zRN0CMaE9wGauYmAKsiF1Ryv5Cml0DqPTil8U1Jpx7sck4xUSJSi8ZnOlDANnDe8jua
AAoxmblOH2sI7kc0xMG/UFOV/A+2U11vhccPky1o0ehnsSRHV8KSU4DZLDMcvL1IIeBRRdNg+PQs
OuEgBCNYEuQYWMCzBBHk0fDS5LxrCFgJOuTYf+YaDYchA/9qkF4ak7syvQ+sg0Aqq091uYSS0r8n
sqks/sndduKetHX9BLeEZX9fgTBAglJFzn6I92pF1lRJ866SyQ43BvAqBtxbwU9mLyfmIDNDLDSh
cPSwQyzxBN2hJbzSzVhtS7dYtnRVxGAr8MChUkKul7GzFTgtFf64oUcSaaX+j43VY1hsuPHbW0j7
1/XMJk/f4dU27lZkmY1CjMxDsXlyYc5EWLCu5UjXKjaxLShu/nV0Ps8hORM6C68fkRGhGEvI6rpN
Vw==
`pragma protect end_protected
