// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0LF1KWcf3LYezWv5syqvGAi0qE4WLBVANPK1cd7IlcepiewHq0o+bpfnnlz2
pC1PdQZUMukkTIBuvmwyoWRXWu3m9HqAIOeWBhIROuF77M2Fcwpsmg9cutbu
/gfMghV+54UZdK2NgGehNMvsWiopNmCC46WlQgQMGzArjtCff0SbaKJAi41T
7ALT/ATyrjNq8yk0WkDVmLR/E7UZclSh2NBViUAUd/73rcg7zpdOh9Ny+8xY
08bnzDjIiQFILw/JAc6UAwOngo2i2TC57DhGvSbd+HdtVvxbo6/PmclIrFG5
u932PHcmoDAzbaHh4WqEVvQqS5/rGv/jAAULDXfYgg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MrQv8qYlFxBavshQ8pUBx1PXNkB+kld3cpF8mWQi67fHrTLQUHe03r4eQ6WD
zm5XWAvK45evD1y+U0Bb3exkX2YmcsNz3rirLlR0DkfKX3dpCLvPdF0BW8iN
ogmqwr8TK5Y0OkMracO6DiV+g2uyNLY7jEsyKOcRdw8kMRvQwFpfnWZWg+vB
W2Ym9eUbpIdvAuB4QV6g3d+kSihostb0yzpJvr1JYLOocGzKBUak9am22ILD
re9C0JmGpK+7h2urIDSMqE+4WjE+87QFNsh5UpcQ+NQX1qqCS6g2EXRch20z
91IJqsaH0AhyAAjJmdTcAt0A6uCPxZzi+KZLuiAR2w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Sz0rZfdrMmyv7ICwuXHqne01Wyc759Bpm3EDKH7eVugHLuUtF5pp4TOzxUSt
iF6hM9EZv7a160+4iVD7u862HdklLUa6dJhM/WpMy1I0LdML0WB7Wt4ZtcjX
W87ml8u/oaHjFKwo4YWoUbWf2OzmWFr8SKznpvoI/TwwCNS9wJ5DsvtexuFL
kAWGRQF87C5RwKrW8FwnBBKWls4ey/n/NaGwad1kD46cQ5qTpuIj075glDcv
4FqVnaQJvXVDYJ82LISplduMhKtTBh135/QYd8vS0cagbNJd42aXxOEAhaA8
Gp2TJX4eMKAleYl0kd7et/dANDymkeJx5EiV87IeZQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jWYjB2Uj1IJ2U04pYkDrdQIGJdNY9G6ddHMmwE2r5wuJc5OWijijJJLdmK47
r6q7qZWDRu6LWtX0soVfa8BM0tOpaVtq82PHqC+5RFVXYgI5aSpzkbajJvXY
sCeiXsVOECwMwbzMs6A9jZMK5NsBv1Cejn89+V2t8JuedYKJXOU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
IF3egOA5tyBsotmYa9dffOISCY8vG7qwrGYwXz/soU19LljjHhA/p9tNecJH
AyHOIM/S5xjw7uehvAcOoRdhYwgwhjWeMN7bFZOtfGRV1FzcMeS66W4rX3gV
qFqlTtT1UQw97hfzEVexNsLDoyp4blDXYlGOz86bi83/k/NCDakLchcgdMQO
ank8HpRjXcfUGlt2EdkCMEgMR2SmFSisIujNFwN55upP+HdObXesGkZdalpQ
E5yn3z8gOP2CUpPHY1u+JeN0dxLpI1jcH2svm5uhdzFNPUUTqAZkYUiWhCyh
QZFF3eAY7l04rv0Ooo4MnxrwBB+v1DaE4p74USjzu3GEuLxHm4Yha9yv0nef
a5ZbRrNLr2HdpXjDWLZoKs+2G6Bi54W6tuANcFoNJa88SK8iY61NpSqbD+3A
GishmWCIYPtYO8elbnzqDF6rsgUntaezw9L1vlVXryCWz8jJyBs098S5SZVM
lfhXeHHWandpeQHs2/wtPLl9e67USCq+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LZbVXcDUtDcNNGGYtRGF4aTnrS44z06gWCUZes0EeysS3nA9I/E+bSC8zw7S
e3skp7feBhqX3nGxJtmfi9Bv9KSVDRHb7iNQWJmocsX0yOLlW3gzhMCB00UQ
47N8VDmfEt1NEJc152J/WS+PcM1oOvNkHal11uueO2xHhg/O3d8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d6W84pZeEjoVbYTR6j9f5cQn7FTM2R6YyWYvfhByvcd463uD+dAMwh6+oMgH
uLhn4LcdNG9+ilNahxXPkC0SVO0vtFs1K3d3/TLf49pDc6jtZLLQ+Oultvcq
93Koqxvs8UWI5NzUh1Z0GokXaDHFiGTrmkh086IfC3tVQBFc3U4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21072)
`pragma protect data_block
sZTq/Q9qqdDk8OZOaO+Ww4kdTyx6242I6oiJojYXHOgeCsL16JFE/aiAC7aN
+AlOef2vBDaCv4qXSYW4X0hHGSDeV/issZCC/dmiOZGeymh7MbKosvPFWQZi
RvqH4BGiOc/7M3p/rSyf/iTz6u1GcPcaibUd6YTYz2dNDe+68AQzvGAfTKvZ
9CP+wUj1TEnc2LTKZrDgZPikNVO5M7F2Wg88Z7beTZpdW6fZmEuANSiyNI2C
6V3E8JWafGU3LETxlrCEPMyFooOBUkKgIjuzmBb52Tt+0CtPns/di0jCyk/n
BIxjoiQmBfYjic8S2rw+imYjht6hkyKxHbSFAXeHFsuSV0PqrpT/Y6S3ZPHz
1Fn7/UGZqm4l7eVu6c6cMb7nLBnPrGsyNgBCP+yV5ZXsWhgKwCdltqt5kyvK
KszIzg5xyLJ64v3Vbjn2gvat9CRRWxQZg83s5G3vGEVAU2LeYHU4O0UFah5l
10JPsY8YVzfGuUkc07Nx3gYJIHMMzA2sLai6sc8IQO9RzkRCkGDZs2mY01FD
PMZJNd8QYvICTzy+AJuiG/H8dj9Vzp4drEjlabyIXRsqbOu+0zTZ8Is665LU
pz+5RiCMcszG4pqZtuKkMuX+zn6iAcUjjFy34IYj2ODqDyyg3NiJR4M0wn/l
0dEPFrnWnYGfQXSVToVm0gX0K9vOtf7FwaPOZGawen+BtlzkKa7HtyNEakpE
XZQQMDEokHhP1vCvbDTqVBcbG3knSHVu2qVbAA1RmPRxkZowMEc6OA6ZEqKk
0dmaPgi4BdL6UbTKUDJNxh99Z7FUlk+P28LXGDTPA6iddxHMGMBEerjR65lX
U5VP7Fe3/aALr8afKR9c2smbDq+g0hFMJYERXfPzGCwXVuMuk3YIYa4M4iV7
PFMf1rzX+aQVt2dIt0EiFZJXlzvQJBBiW6cnnAv3Pe5BzADx0hBjWBJPWkPO
xqNKQiookxc2p6jGNE6BJG13lTWsxpGSpVGIgqKD6BxaNtswIEnNuHEziALa
fo5ok4G9fW7pJ2JoKtxtU3F0qG+DD+chm+AGA5i9kRnJ5eMBLG5fl69BbLrL
pGGfXCzlNVab/7c8ZMzynWhezYj/pSsN7AUKKHZGrX808uIiVRpCRG/PElkD
jv0i0GkQQxA+XT2ILQZ5Y7wUDO7x9ej0V14Nnj3WIlupHUuzB6zUoD7NeNFE
y83OHJvGQtBX8S8RLduQLVWAfMmOwHy3kWTDp1cwrGMstuSi5DvqKQw86TUD
9VX0DwZj+ueIFlF7HAyD6xkoqjqPBR0fqPYEroN4WutJTPRTeDHIENdLJHiE
ny3zVo8omIV9UOex7y8/2WVD5laH71yRk20s/wcOnPFsUC4zQiuUqQlea+13
AYK2IzENOMiMEIqjlGCk7urxu5OkB858giQtdK5GyHX4A8kWRJ+R8Yc7gG6E
8pABn7K8ed+dhSj3Pq2YAXBgYrgEvTVya5LYi+1WxEvY94vSHF9jAKOphg4Z
GCla1Y2tQRU0edKR99LafAbUe/ujwD/NqsrkpGs3XdRxbqCaiyBAJMNxCV0a
bWPGPCJz89Nu+10qXqUk5w7SFrgABIOE6WBqO3aMwxdxbn2yYChzYYw8G/mi
Jd1ql9tC3SlZCtzrjx/g1T1C3fGQi+AydzXZG9j7RcHzTnNzhnjeoqi0Py/1
epAqrh4bQ56kpUcib31wX5HZ9u+uLrUkiF9gCrcPo/UJe8bXdJkb0wCdzZ3w
0b5OZw32jm8mMJkSu/ziCapBGdmOglkxT0TwJ+3wM8aOKtptQMj3nCHQCMMM
Jj5REbkBmJ426YG9JHwbz+dCFGz0D1RHHp2FRf5pGGdXWUPpGYzq0m31pPvz
u3qWMU9ZMpQBSYuuN41MWeByBml/5gLTLwkqk0UxVmG0lGvxK3B17xhxNBYZ
WtY+fLjqC0ncMyVwIQ5WGBY5W7SG8H9u/M968wiAKZSWgg8An2dgant5FKpE
6IUepB3S9ivIC8rFhxmDzJFLw9E472lThqprOvR9PLRCOn1ZnjtDaS7Lz4v+
9GChcqNTv+NB/VmZDFlThorKj4b4Tle/v4zkxCCvoSapGKRcndom0eGU1DA4
Yxh2JeHUpd8ANEnXhFarVOIMQcEk3eCajn9gAEUea5+ZfbdLm3ZkcqDVxaLo
zvHep3iiz/GeI8pRBWhG3VruaX3fQfdYpDnmYV5YGJSMjKmR2S1WCqDr8b1w
a1y0t6qFp8mIjQdORe8E+NkF6aUF4YMkCFaynt4JmJLTbu6OEFzmPZWtQ3WP
zniHwropR4uCRZTBUb5csydTN+5fx23WqnFO1ucKmfwaYljv047IkkVoOEvP
J3TwToDqGfAn1vYGs7uifMUTRKwp0Ioy2wYJBTfje15Di85bJxDjEcKClG8q
O8V/xISZjT4WpgWebxqfmohbWMfyh2BAtrt4VPseGXbAQTNeZ86d3gQkXBGa
5MDHU4NjcHr+uNCaARJ46VNrnuUPSQAFKHLPQo0lCUT/l52tpm/Twtp7c45B
J8vu0EihdLyqd1+MTodhbN28BDCuId7wOJZSeucY5zfcahFbdcdhqjdfmQcG
6V2hFJzwC88N7wcQaCgKov0jVAcpKEHnACZX3zA2RtYXejjAxinEIIjB6osv
ExDKCh+LvVYaSLeTtPli8yL8wqrRee02FosnT5T4EesVNTLqiLMSp24qESLr
JmYcK/Wr4s8/LTLzY7wshk0HI/QOQRdppiMZeao+I2RrWgSLDlSI0fciJrzv
h4FbpvzrnBwqzYG4aTgUgK35unvxb/Adx0ume+rk+g5dhoFzYanU3iToJPJC
iwi7dI1/sv8pVjNr9jaTHdV+u3fY0CYbLpd8DPk+iPNc4rkJgdYkibE1+y03
m03VODMoMV0RtAGV3zJOI1UP05XkYG2c0v3b538S/xaqGVa3eEh3TBNEgy1g
yDmGx8TbmJ3VGS/sIT/MySGjhhcQrXiyioAfL8FgAfE3I1bDoHiu+3LNvbH7
h+BxO1VxM5Nij1ScudiuE+a+nw9VwRSVJVfBJuBstV1oNFfln66A/S5/Tzgt
bCqvEqS1thF1VsmVqPeZqvfCxWD/bieFSwTROxvzFgYSaRRKfg4N7yOjvV4P
wGsdZMa2fIFbXcPIBbnQAjmQ+w3CYQa1iDRZw1pqPVeAwz0l70HGf8/C4h0e
yvjxCmDy5PyIIa52pqTU56p6KqTgX0bPeEXV66qRN/7wXQujQef0j5nSuRcH
dVAsz70McfLwElKn4CFfzTslpxqxSxlvwpLQC46EW0XmJYT1uMzen9e8c2Y/
hmbfXg5mT8YnDGTVEwZrGbX8y1z4pCgu4MkEsxXAAr91efTBrucJXf4dkRzf
fAaIemgO0Pt/Na4/YZy5BhO9mqEwrVXFSCV1lkgGmddO19rCCaqGnipUUTBi
TeKZuQz2t++AJQXkX6qU+mp6pmxpnUz8uxHvNV19PB7dwyolnw084AuS9Ge5
85EK8tDC1e3PaIOenxNB4Ufk3YVVk/qDeAeM1KFhhspWOcwi3eZq872iXRIV
J+rxgQA08u0mn/ia5YliDrYLSeXkh+2ULrRI36OPpl4ditEgu0gD/edgzzGV
rAH3UsFa4D9TivCaFnlR8bSJTDDVURAf2r4tjnC0ZP/CoRv6KxlFXxzQikkz
mIauj81l0fvf6E1ZERylVYiuv90xA3FDQ3uJNuMfEKheV0rGeTnEzJkwMbRE
FqZiMaTFNeD9r+b1Ulfsyooe+mkoU8A9qM5E+SS0yGXasa+RwlvZZK8LLdRW
EuFuduDvSkeLb2UiMLRi/x+kiw1At46HqZ+UBN5B+8sqVPnN3elSLCQZuAeR
YQ6+LzY0nT2IsrD7TsPwNoWzxk+uRW4RyisXDISltOW9DDD+zrACTvt3hyly
WZrCIboxl79JYlK/Y8tTymt+tcw2NT1cUyXAGWttPMLrJnonguk0Yizxbu3j
ZrbBjewNGWqROZOyqohXPeqdUMw5DOsPwVp88j/z7NUFQFpSwXmHmNkLBf0y
7fnW0nW/5UOVaOK43ZrNATYuETUynGWPYsmjmu/pcJU04SSg+LQSzoePGJMB
XqeiQ2Im3/7OD/S+d8EV42ReXsQAY5jYxFq0VXUCTQh2ZcBw7sbfjDE+0hX3
OpRELWvHopi7OYYrMMj9vku3CP5j1jXaQl5FaY/b62rJMGhTF9m4CdgtlG8c
nKPqJehhTJ1VTGwH/BB72RzLdv5EnLpTgzenC79l8QisOidNLn7jdvXz6fNK
o2i8hD3lmPuU+SCkK8w5Xjnqo437etABVoysnfJ8rI/ym8CQZBBhF8AJXIex
kRPrhGBWKFx5/QfY0E+x1ZwfpvEVnDrt93Jhu0jTD16qov629BwGiQbRVXu0
EyXNhB9WgWemSegzV6hmD5JYBGmn84JIA9OCFFqj35NWQCWIz35+KQdnOZNp
EPf8c1M3VuxEj2Go572NJXe7O+v0r0qj5zRgmUZLuGNi+epOEwHbTYRVCy4h
LXsS3LkuNETLrPiFeaBzm2jFHiyIDSLJm/dMuwKxO1H0ezCO2FXvG7UlqD+g
0v4/tDAv9nWhOTh8/23r58WV4y6wOJJLk8vKrQsMaHzM2L8JYtAOImQeLbtJ
rg+CXAF3t88xXfyp+iMlljDj4DxKi4BshqEMgfgJ+KZqreEqgkFADcFDlaNB
nFxCXwtDISijJ4RLeSk893PHk2PS30H9v7M3/daQIKzETexD2y2D7s28hutr
ak8kn5hfGGvV85Dq/7+dlLisW9lxIXQ9CrOv+kQeNm3PYP0EwIT0+uEvl72c
QQybY7tYTgsiFERIeUI/fUSuQphbQNWrDGQckz7w2k0giI7XnrbD9zEJByry
DjkNZms1d8GgJn4zwEWFKRKECKuxiqfreSYyyfaYprFTrnD4pEDAC/WYyAxC
MsK137dGDXI+6GE3xBKKe/TP7SR0fk9uJkkcBPcpG/t2Q2I06XH8SzhvUdPM
2Vda2M7x6MEEfka6r4IoV2HQFhHDfHvVMfMvV4GtMusO1oV4BGvtMrqABByR
yKosI8BQq7AOnWmoD82qptaL5PVK7L4cpFWbsA2diNlFVffN0JN6u+HTUKwC
OTTn7c6sib+SuqzVdDKQbocdfajJ/aNDhiYiZqLLz88X9mXDF3BZJSbiDBh5
sSwifIzep8Sf0YVK+oWbBiyjoApJnwy3R0CAFsuMcXyLOP0cH8/kZLHpLBKp
vu+euSsfzrRBoN+Hy1xZKcMWRIYJxglo3H8ycgYspoFuaRnxGLe94NeKjpHz
sH+ZuxdWVHinQccYWgVUCQs+03EfgRN2PcBd6NCgghkloRC4/rfxnodhpRep
HhNOjnjC75CrrXBDgWD3z0Mm3PlVx+e7EoyXSgBwcgq9rZUFaPRXCEFkGvwy
V/y7WwGpSLC/knRZaudMIGRqi9E9q6O0ZTDdp3fY8iLDBk1QBPUAsVPTokfi
bhpUjkDMusfGITqFD2QMYzrj6vSNtBe+VDDVoCQ8hEbi+q+/S8o57BpSovF8
eihz0/tjfcyJTGTxa+yAL6IR/b5eRCVuR3rpyBUuAP9GW4FKpO33/K5DWlfx
uV6P1bfeULqh9NMF8EFGKAnhtyjk5Mq/64gTqzNfroGculY5mN5v4aLV9zCR
Kq58nUfeEP/m4Jnib0tFDHqoNhFZ043Ef1Ob5SwOyIK5I5UFKtil2KtpRGbf
xI47Drl9dNSN554rIIu73E/eVYQRSpYP/PQWS4Qet9FC4T/a62BFv68DT7rM
X1+Hq1M9bDV3F3jgamqRDB+8jLrWTH63JKqEvfnt7IDKYuDw0r34PTYNi4Zt
PSZmwBNlDmFoMBNMsnXZHy/4LQiRq5BjlFjLyvSOi5ffJdRfbovEhg465lh9
tljoFy0sNbZH9w96f0ZQC5gtxj9H0QSYR5l/raqnjIlNT4vQJ30EqWf91xyw
EzUsR3bB8LL2fTifS+PYzPpGoRhj6PDchsZbB20wUzJzbWUEkYBNSt4dYqBn
G9Nsgbl4hQAEK/sYebkTe7bFNPnHI8y5CXDVOYqDavvpKaPpPkm14+fZnwbu
Y9h91lkV7eiJNTXbOzM5HqvA9UUOdztXaIjMVb1ikXHBz82zj9ZTP8U+HhR2
nQx1a/DrfugylpCb/0vZd9yqN8bqOGKQ3zx5ouFAI22I1VPieWTtw3NTlEs3
gJpgI6a34/Vmf6e/6M5YaBMAVWGADRWfmbCHYuhKoBkc10/m7kzxPwWjG/CY
72xrTywWI9uxe91i75aCRNTXIW5/jsqOJ/bltC9T9F+ymq37/yHkfdkUygKV
0hO/ZfrddsB25+AfgDlAqQDHyjvVbO0PcMArww26jn7CClkFrYFDxJgHObm/
LS06cBFnmUJYbyLZgobrvzNhnjfUatnYDL+08g35nAA5JRyUfVfIrPtwo3z6
X5Yf5ABaWNVJ4W7bcvb7xoIcy84hXN4ccva6VQSGK8snXzA9NHT87dKas/zh
NWfTPkz1AsIqMxb7DYaDQFxfZ5rzLhrc/gb+DUwEwTASOV2wU5dkkL0YvPM/
GZUC16FsAt23oX1hj//H8kdJIeP1cNgTYpkOR+5tbMTB9m8H80q8KgmS040M
ZxB9CW5lzMjNbn/4WQuuA7rI/RoGJg7XpFMgefuA/dctFB1GdYLge0wpAh2V
UgmVoEBB5Enj2cJCbeoqWRh8/4+7lARbfLHmCiWWIDj9W6GBJOuBydq3asCK
SevIo82Z6KkZq6Cs38IUOr07xBIFHy55sArUqelFUQMxWXZYYnBqAFSwNWiO
W/cFX48P8hUsRE/s78AMc3ciZpy9S93Jl4bgTGXQOUiSyxqovHr5j6uMP8Yu
OLrXThvNtSKMl/9ZSrYVddwDL3MhwaF4I3p7IuQQsRzPrkZUvw8cO/H6wyhJ
K3eSgAdFur5MCLUbPhe3UF1pYHR51I42ymR868/ginWPteYKQ/ECgohjMek3
kPLW1UsA5/wKXxPARdjEqzG6xzn8gtb/aonmGDO/i/IoNSzffKHirDM52rg/
vgOMf6byAqNgXBIPYMnsaK2jZGo02w5rymqItpzalNt12bPA2jTlJgLpgxe6
uwM1Y2G7MLLm4sDFK8QEQ0Pn3NGnCC7nsjUQ2UoPTDB/t9kGPfWMHzoLj6c4
ECBf04UmYUd/tzbjyKYbNIS7BFyQmbr59vgTkB475dylMxQ+XpC8sbxk+3bu
qizqTgVozJiFADFx/q4WZWbEmSD3r52ry4PD81v4cuKVNoHgWfI6yRsswmiw
9aa50cPz+S4WHl0JycAVrtlCsD5H7Vqt79UQjVggSDKeSEnl/RqBLYbtYMmn
HCjNPEhHlAQggWAr/+9vqOenukyeO9mETRTaxtHUg7zhduK7GwR4OsvS11ib
S0diAZT+4daJrOOrzzjhuAzBtMQRPB9QlxWGoJmjGHc8fPnOArkFX+dqCDen
OBLb2XLLwsxLqRDWYrxgHxrxAxArJSOS90/M6zKPd6vOFv2Oc2v90CBD6r62
+GpMBIQz1qeE/9wp0ZH6usNXVA8WQbdygqb4F5xHOXgeDPZ8P90/5YUdwf2i
0U0J1kTH3PHFkOQnmAioFTB+C3/zaUw9Jf6WNCYjjzvYlv5ndnXdgo8KZAOo
4p1VpkEd0h72P5rK/gYU8nPZvJP355A84LxpjCwHEin9CgY1WZbSMN/E7BpJ
ywraiqtLZn9fRHGegur/fzvM8hpx+u8fq+Pdf6EIqZjZPRkji4c/2z0GYpAo
7jEYdzX/J7fufp7VtM4yKrRaE13eBk1dG+b3fYaD9bZPGztMBxoejUrMXE0+
IA4dgmNk6n+c8VXtXLqLkce4bmlM6G6zlBvQ+HGT8GwaA7Yq5a5MmNtX66ow
FO0BsAxHVAaN4G/TWrfyRqqaPOL6XT0RyIq0BoLBWFWtdso6CdS+auMJ6Z80
9WkEgz2hVDIu6Yooqe26607nM2+mSx4mgYYV6iV86EFUJAyMt3IN/xkF5Hyw
zlR6iAmf4xWBZ0VprCjO/zEOLs3dw8/UgOTTv4nDoiPUfObpB8ZQl99Qk+Ck
rnVAa4ja0/MbMLl4WrSiY4t+CxvtUV+Zwtx3dFZE7JabA3ch36cEDtkJmYRs
L9T1HwvvvJ5jZ4/mfGudOuGnEt7hAqFYTkimFz6htgdPO4SnvmKCh0Wo7KXF
hDxmfT1IAzCwE2oE1XCJggCulgBLywOlQk+FuXX9D2VhKY9+Iw8baqNt6kKH
KPq/bRfbfHHyp43YFq4+RapA1Gkcq3qQZmvpTaSKKSP2fKT0ydLtJN1x0pdj
6l1p2R4Q6cpR2CSe7luZR8X5AI//LyBAc9gnvLnRst58GmRiVNcJmGc9Hagw
oSM/FWhltU0fraCAyfurL0O5r+DYvPoMp44Q6yD7FMPGnfEUYgy5hJ25ogsv
IyAUCvAH/XJx7oKz7wuPFYMZfuEeIwBqj4t5+b0/e+m0ReJp0zCjp5JbWJPY
msVnubmQ9/bBNXDIIw6x3HC2qePhVFrR9jIraIkgCDtFt1CN1t9fT5aXN/81
vOSq8F4S7JrzlAKMdKohOrZwZiir3/eG+Sgn087xxt/F9/oA+dn5UVMbdUCI
HjzrAEPgPQb+6PFv3plEqwkD6+jHcF6SUzWWB9ahq7idSPMxqhHAaXHT8XNQ
u0wV3MbDANT45bJn3Y7Ppu19+/9mpJ9iEhVxoSKXzQkeZdP/Teh4a1qdE+nX
REYHN3K4tAz29ik2Bk3RkVMUG8Tk0cNfwWI6pytLATalIE/BbChhp1z+vE0J
7nOHlOnqg60Yc16zVkCH5R/KDGC7BxfC2xNYxWyJZ4PgVHQV1jzztyQY3qGL
0x8iYU2VSMlMgDj/mVu4dUgJoa+PXDk8mwfXUbCS0zSQPnlfoyBbAIxhXkUD
u/blA9FzUGv6xEsT/3NJIJHXcdBG3SVnAHKxsCciHqOmtrrtqeoAZMEbhUD3
cjvu8QtjJG5e3yUgGR8qCcOTuIccsUxXgrH9iq0lfA36zYP/BZI7hBANyuY1
dvs5YUePBXxQigEtU83smYTa5nTJAjKV+y0LLLWSTdsbO8xUoGUIYNgCFNzf
ctL4k5R55mvCrcEjsn+RoGKzegUThPbTpx8cwybeErZVsiVi4lAFQwzFFuKE
T7d10s0toL3qccmeAJMB7IJKp201dsrhWX6dLi+J88X9i5qAYkK3KyIE/+wU
UWeVC40jCCwNSFvkcElNDAg2xZGQCa9cHKz62J3z6KnHvzkJIybmHRI2j6UI
Ltk/Sb4FXylo7zA/4wu8UPm/Imx/NJVXfMN42czxq4X35L5o+x37Ato0Hzl9
YDYF4SOG8QxSgf4cmrH9+QnsR5SgwsNHqcQejw8XNeH+cQyzm975JQJTHoIU
fGmIKwlso5VxvrLyYoBx3XHVN4XVgZo0/lB3uBN1KjpOMvtlzvucXdUw1L0n
dshmHoKFJD21bZjVuuUOpZQWGe2Iowz+GH4RWxlp4FHAcNYdLlcmAscIHehn
BCBzIoQXcGGsEdmpmlSsYBpMsCPVUjWi9MAiWNs59YPs8thQa69jLMu5WqQw
CJ9SkqQBWAq6+iXnp2MDfBrsBSc53oebCLpotAa6V/Ap1n46gaIX3JiufsRA
Li+on943Q60vMDZMxjPjm5GTKrbsynP26YWEHYkEJqjyDT6h7O9r/LM2iJts
C70pxtA0yzjUDVmmG0FdAJfXjoA+//pY9ImXCmfTy93C+jsox2VIdCgHOjRn
JvzmU1PBf6AKoFx5HiwViW1CqhCNIZyARUHJray6hdDRKzXWUDC0FyW0tJpV
O62qEY6pzzUlZ9RP52k9b6TnjhOGzEg2XiXDh+MLDI6ueol8Ah/Hsw/8C3ja
cZ8T7kU6z5MulHt9O3U3e6C4ZzqKFLbAJ3kYqhtr06FmezptsGvH+Pxjr27r
POCm6yP3WGlCjrXHRLFrZQcXFUoOPAiTMrlQRG13NEGZlBRAGwcXsxx55FIX
pNX3vTBioozdjizUBvKTlzdjiXKJrxHA6v9eOAn/7U0z9bbf/WQfu/eQBWaV
4qgRdG01sUNzYB7mi0LfhbMNJgrF5K9xTeZDJOeVHdbYJ/U1l2g6w33HVST+
rtuCRTnF/PjmKeRJ0jQCxwJ1uXiJmaQttH7MJJIMIS6PoY58El4l+3DbcQRe
j+oJMloo9UE2UWvIVy01KspmzMmvlG1gYmpsl8tlmJ3SpBfABTam5RfzRiPt
YqFD74vPufmjMsrjnhXQVvaIivKdrMs1+WN1ikrIYtPz7FFNqitNU/qKuwgo
QpOrwzQxTnE4UBZEr6f6tCSl3JNLO/8CNA93JA+TLEa85DQrDXndmDX6EpmO
68GxO1MnSSpqwhPAqfkJoeVJpDhrNxU4oXoB0TVMTbXECspG1tQU/BFKSJWH
FUCJT4Cp1sUXc5khJkLlUE5EQyYMgRLclbZyZ3vKCV1k+zh7BUY2Qu4fymAY
Kb80NobjCOk/wfRsnLlWHcQ2E/8V8ezZWjJkMQa41Bm1jlOGqin8sGp1FAAS
rgR6LXSxmwAPH6xjRWwWLCzo5iy5pEHT0VBuRnu+eoj0SQxTlJOVBItesLKi
fkuJ/QIyzp6iX6C33pnAnHKaSium8MSPb4SJGv+4QjLlvBrqLLwxi0uWEjo1
oAWy9c0Y3MNx6O+kSgXCKuhoQWMZU0nVS6cn+xQbzMZ0ds9vnQHWzOMT8g1U
n6i9/rg534oi2zqUiM+mDxr8veeCIs15dadOjen0l2Ma01esGD+V/K7I1Erv
b0PIHYlkGnf2//iIAdScVjjQQx1DrN43/6rd21OwshwBCPq12PNN/MRjn/wB
9didIBu7al8jaQDAAYZXGNMRnCbSob0SlR3+ldDqyzU84KNgLy66dNn594eN
eCp+wY+8m+HK0+rY4Sg9qMwHHAMs+rFIgO9ZSYTINbmLSPS8/yRTN6BVYBUx
X/tYRN4JVJ6nYc6IwqA8CU2nwjU0KJMoC8pknkgJx+nouooAY+to8kBJzH33
D6YGMnzsFx+mi3J/FW2JL5x5P5kF3dzgWa59RXU5rct+6MTvCKmjpHHcHqQR
Rr+lXIYJDRv/MrY7i3WphnPSQQ4uWK28XTwHxq9nkseygGfYXXKi1BYNAzbs
GP2Tzep4KDbZj/8un3eCnFrwNXd9KsmDW0Ih19fOzf+PgA1etRUS80y2RZT8
XCLtZxuzt4LKUP0viPZOCiHx31I8C0KKAg/UPmfTzth+I6w0MZI0ovdasvOV
WbztlDs+Ig4+x8TArkeJPdb8I2bJKuRzSGqzo/Fyv6YHWHHLALQI1SZ7/ExP
rlhoiDFL5IMG5b/bwqtFJT0HfQ3FaJiXGbZKvuTA4IqmnQR/bl0mhqfAtqSw
rfW9Rp67fJKrWxnqHuuqoFLtMA4qJ/bRWoTbfX5cBMcEK0HD9rrwV7JLm3Os
uSkf5tN+jLcfqzYHipvq+Susw7XC9AXrdq36/8lbVGQM0dPKFVsA1MnFxC+T
9qcp7212QkZwge9TnCMQbq6DY7SAXm+cFRAZJF+XPzF9PsPnb/OiQCpLYunf
dZPcuSzryv6gEP8nBRMg+VgUkB+wwT7HWe7Jzv80Guefc0RDmLDydOuVs2XQ
/VFQEA0VkBssyvk5/NemOhJjCYOstb6+yJqCduUwwdHJGE+hxksmz64a8Vh6
eqLlhHW6FqP3CYxMPCOcsd1cZcwvThnlw7Bv6JguwGz4rS6zc6H73FlbMBFx
1LK43+eiz8VksLHIXUI01jSnMYQRfk52OXknSGspfQbGhphva8ca/9ISgCBc
MfFTNM+Zpw5wT6BVmi8S93hSsIIZxJYPTogBebd4fDVFaD7ctwxMUFrBk6TR
6M2mVtC641yXeE48P55jlJE8U5g4EcXXaWqeYwIgwQ06nDDt2q3Rr7nB6ceN
t/6Qohfw/xefisgV3ZbOCXc6WQbLFPPdRZG+jLKkpgWUmr6z1tliiTAyRgo/
XskzSWCrKKeJbM4QA+9iYQ7h2txClKSd0QhGI68gUvklDzL/zN3FYAhLS/gx
oM3Pcw2BWZ7An9zLjFpZqWxCpU2bAeic4MNf0BBw7LhJKBubpDcaTc4Y5v6Y
LfMxYdt06ugFidgJ+tFAXJz9C13M1cLSVzgvym0zNgtORwCpNJ9Ta+49Uybj
sQRRpdpFKINZvNA6pRcEuYDEkUhSXtgYmg6ZeZfISCbI0rTF7toS1hU3167I
WjPTN4JyUZzp1RNnzqQ+VhH8pKF30Y3tqgx2Q1EAU/jjZsN9PgruYA2XHx15
mwOJ69DNHEM6nxu6e0m2WMn04Hi74MTE5O//4LjxmiGSskxaMVSAGIINNzr6
j/uaFxe1j5S8WfAvObBLGF9Qf2JuWauy/WlHguCzGb2573dClyzb5+KCdDNA
wExXCM3DBPbhMgYU/U3kvfqfFMYbW/qsAvm4an3Ro5qLrIqxFD1vXCpXpslL
G/GM0c2F5T1J6xmgA/Pu5xlC3sfwieDA+8CpUTTcSFdoftMaY+B+j6QTIQ8R
fWRJdNrN4MAJrJHVCowhKLgCuQ8sr5rQP/0IcU5vcOVnCocg/iNv5TiNVedZ
yzT2xs5rNMOgM8JFsuo41kKbdGDM+hEg2LD5q8l7vWfe02VdGfRboLxMvRYT
wEGz/APFRdsGrBcuGLvW2kZhqRVKJJrqu6Jou3nTOPz1hhqmDgUzxHgOXj49
Akg54Zlm1LEixHPn+iordEeTMVVwIs7UyCadMmoDYot4czjASZOqR0otM4jK
3wIrtAc5KbghfsNWkb8hZ3lNigq4aDsZBpvr88pbkAXfjpPgfYEoZ2viXOn0
wigA3SjZgZVMiz+wfVosJwo4++kqIVj7UhND+gKQTPI0l68aW8ptorxddx6l
CHhGQHZIyMOHLEp69ywIsszo0ozQMWXtEYdaWra86LodFTwvJTNLrzmi20LF
xzwGnnNQXNoKRIuk78sVwqCze3tg0O72qtEnexgzCpqzTxrhgE0OXc3gZKxB
rOLs+NTfswRAi5nJ2vR4fbsV3QzqzlQv3JBUbq/5gNit+TpjF7hd3HXGmX2t
S1KoUPpx627Bd/3j8hh/v6KnH//5h03aN/e0W6lgM5Ze91zlSdYwbTNXWNj8
0I/WB7hK6Wk46YIuv4Jz0jQ0wWfB8dOS6KuHrgRnIVVr6tL3zoALXV3atz1x
Na4ldWN/GSLG3UOv8oNBU8sTlYlQ3TcSed65A+4uQQP3w3WS0YEA1zz6HMqc
30oZ8UA9KzozQLGFdZTeOu8iUiH/0h8S/yK6VbtXpOf9T9Old8GJpDvgTYbz
L04Q0SGxNppbCzjHmWBnpS6r7VGduLDpC8Tr1Xn6MU/aRgTE3DaENVkBcwzN
GOBBzZcVAmkEjm8+/cOn5ATchRKLBgJI9BI0L0A1aBSbcCipem4Ma3aiCtiu
q4+LlP1/kBa8d1boHOgGrGrQb6r4/XYTixiJuaNWSddvw5s6Rgxov7YlviUp
tbzsN8mduTq6cioQ/bnlm1CTUUyWbf9VtqgSF6/V+RQFkjlYs2ebUFhe6/fU
c8ZDnPAHWQrubgktAhPCDCXLUHo8Cii476d3yDHtRL+lc87Uv8ctUfqLuhgg
zLKXp+tYSfXRkd2Ot01nmu2DGxdAEll9vRzFptpNLxmkkjHn+O4626bUGMpj
wjoTDhw7YL0BiiDkoxZ10qVm8lPhRjvMheXN6zStSFtoNXZEw4OYup6vXDVT
VEcIfjpb/S6gwvV5NxLx5SBkO/WBy0AJCIDGbQo1lPsy3x4kjyoLhEUe6Lkt
gJlf1TELTMJrDGywwM+yYxFJnutVC3VqiJM9z/l6btkPpozRpqV59JynHQvD
KFkRlLkDR8GquDmY3xmpgr846OMANpK9TFR470d5uUb3eM+iltaP4WZ1Y10n
WKLe55vHYsBUYMxD0ML0zxeXDU0gzOzvIEGs0H0nBTF7gZJhxY7l8637KbPS
WArbIPHBt9VZ6QyZcFVMcjl3eASHoxIAA2YV33NiPeC14FqMZt79XLjKrdEH
KrSxrR3fkF+odytYbs1TsKCaG6i2rKoE7Ztmh1EsFisJ4F1Bozv9VhJ2spYG
LYngAaj/QRIeoLjhD6AVhZLdsKrgcsYpob/cVemgJAM5mIJ0iwiV+h7Yp6jz
oLZxBoLitRGjzU9KScI6+tw4xp2LzN/joHU0RACL4O3BTaXnzDK4xflEIDlb
PzoPvwQhoZ9fJDheZDl35pgGJs9G4vXWVd0xSQbarrsncXMr0ixlfUP8BafM
DmmdrzLm0y1aDlUcyDx0UHld+CUmCw5bMXJz+KWXKR5ZUZkLdftjk41uXy1D
EFa3kbQwS4tyiUl0tLRXEecGkIMA0l/e5H39yYpYKBsaLVi7UrSnnqKlAkEs
FN+R5QzWjKB3dk0cAN4vHO06iaW8Uhys1qOdOjNpIi66Jf07oYw/PgxpkS43
+bSFE5PEdcyT+6Wu0UFWCPNtPQNX21b/olNgcvAz4WVeJNSs3pfVYMk2bea4
uV7PYtmz+X+K36bPmOVNlI748BZrFEgS7A27tZwHrNu+n/LMP1gnoCb6oza3
+1ZKEtD3Hxw3mMjCMdWa4nwHrEr1G+jXNa33HTDIxwrnuYyNPJDbY6qIf7Qj
WthwMc4SaIBUjn5FUIc48cTZiDzqhJb8AFF+DYY+WryCstYb+hcnP9Ekzfdq
UDv2ykbo5yY9bmcjdQ+iAKXUUALs3bTVAVSuZIUa4DMpLmbI80URpB4SWrpI
2mqDbIE1ufjVnzPP4MH77ghenXUGw/C3rlhDc529W3ZztGkuIjZI+84K+yfC
944PhBFyLHmgxd/IvMtx9jfar5/r3iCpGnzeNL8lkh7IaQEj9F/V8HB18/YR
U7U1jW+R+ydZz1Fb2XMCXPP+zC+R6zwZvaEjzIwf2ylL0c/zY7U/Cb6tutoL
7DwXtp4dWrSK2rqfizZOogPCEKbOEHdAQpgjNRZZ6d+GLUJCaoiljJ0I44aP
SYp83dD0kdMKGq6as31cl4vuVvIAXUqsoe0TT6vCql2aq7lWZ/QeDJ5tmh3E
3YTiyEJ7OL82T9nmq09SAVLl2a89Jpri6hQAnyNnA8YeIrzbN2BauBUkDR4l
73c98w/rIzq51DHf948uZikpMe3N+iVmxhTCEn2acAoJ6oUdOCtb7vPlIHLA
FKqgkJhE2Pb/+g7Zf/sXZEfF8PyMpA922d+t2Z7Kq+PweaHQ2YCssq1STEpF
47eVXPsqUj0AO1m42aEzy5MuHWQTBZSn5yLGYcgKfBbbjZlwK3JGCC973M0s
4AOxQNigtglSCXA9dEQCoHr9uQC4+bu8nvddmu2gjQfI3mZF+C8RH1EGvGpC
nEt6V5IUx2X0w3FJLCng7k3D51iawfg6jQwnZSliOGVh07naDkcfn8c8hZtv
RLYGO6dmWxjqfKTjBhpSXZjULj+QY1WT1zddMDMlfyQz8emdI6ryG3+TaixE
l4WLj7YgBYGTG0uuMGp5PZceT2NkDHQZJ1Ync2rRzGbN2fjkCjcoO4ODthlK
o9ddXkHz/zfTexvrfaoUXXV4s5HdMDZk11M5QTW7WknufJTh4rp76whk7963
c0X0oR6xthO0KUgRwPwu724h96OYZ1LJO3dodVf/SYJl103gW9ltO15O+GnP
L7M5+W6nkkkg2ml3R2S26it2Wt2/TQyYgFE5NG40jg2x26d5LWdwLt9+Q17r
LL/4mGYTKU8ueeJEtrYSgFEqJva1V49tGKQwMv1ECUvs1I4At6wvh/1vz7p+
CeUKW2Q5heeH3aPGszCyZrTT0rBUbbhgA1979AhIijtjxGg6vM38FbpYOYZT
nA1RUtodw7w+K4dzERlMmMg0uYHm6LkL9unpdZ8Q5hRzox4Lo3IK6ypXd1tW
TSGOMiYiMsHV5zlq+N9Zw/Q1aP1DaKR40YPbxGqMUApiWh6an1fLvlsfkgJn
Go4o3O1BGRRW+t9rRHnK8AzGyvwGkU0qQWdJeS7JZWoEFsm6UVzf6jJLXZcM
jOk5/TEWUOOpPJg4iU/OxKocSn4/FvgQ6p/hcAnyWos+GgOqrGWVZaN/JgAG
5M0BYzsIRST6+JdJtu8uU7Pv+f4tSK36A/wu71oVGwdJwO3gpAAYdcJCsg8L
/X3XICXSMPgJBEraeUy78gEbPbZcNkNclBzIylkBybUAi3YXMBIj4koWZjtt
9UM4JOvpDA32WGYpZSL+KjzB3XHxhRKU8lC3TyH7s7AHNmwJOD3tkC8IgdzH
cGJIBs1V35A8lBFIfFhhD4o3P/qb41vuoj8VgxA0LmlrBQbc1aLRhcTsNDgM
Ntgj9pt09c4rT8lRO2juM6IMTtkZ6z+JV7qej0PDrdeewxCrrY5V8sJtjN7N
B1WMFQCtbOMmXCJzymnngh4WhLHlkeyDfwrv3jp+pUV+NeCCsLddwYJX9guM
Xd2fb72apuNuzvKLRt9pkxjjG9QOYUoW+fd+QpFqtnGEYl4jYKb5okGJM7SV
yfh7QOdnG5rsft3qtS58ovt0/jrgWHGWiGB9kANMlZoCtM43qf9QeffZmgRy
CKGSqxfBorxJhwjjH6DYgsmrfs5dcJ9C/3gii6hC35N4l4bzbXC2So6RD7nn
Qd3JSwYmlGtcIQ+J0stWvCLn8GTiIpFVClBz67pU6c0BzIqGI0w3hOYNRUaS
oFLYshCYEEy/KvdUCxktOcwVUekL12ZzHpHWfxCqh2LgEDSwmBk8RaFwNKe4
gEr5bvEHpdnrvLFbSEmNI9w6bxeK/xxeDfulTSFAhwuRnVimIFsXMt6VDewd
cX7FwH7jCeSegDcQ6iszOazhh5aPDaXvS90QxhF40OjHD/ggXEDC9lj7wj4U
vOWXW1GyMbly5shyEL45Qq397dNL7N437ww4I0CZXRVrZQawTRnuethIygtl
BnWH2FXGnDODGZVQpxj0Wlw8UdEAM3My83LYtiXShit7X161FKBujF9A/mKL
XykUZWIY9H2fjvxtNO/oSDCbuQHtjSp5yylYLeFhmPJ35M4iLwdlPCgT6z/Y
FpRN6IGG7ffSNy7enScizchqRG7zd5pFjKQNcD7iili1Hku8WFPRFCgDy3xA
EdJZKt9e+/fhp6+a/DGZWShjrlkDM3aE5Wizn29Zo7c0jgilXefLY0XJ37ob
riMUmvG5VPUjJzmpfh/Uknc29oVY6/qvPJl5nFXnPVcJeldV3HjCEqJVs1hV
htTmfyXlrYY0dHRWOouKP4YgHqDT2ip2A3C+GLH8xL0GMuzgEBPwwvfbeKHP
wdE07+/xEoNMOOKAw6YG5trNh0M1AFSHdRLAHSzRVcwe1USTcydAGCJRr4EK
vpUgYenGId5a+PIShg0ZruySs/AS+gckvgOcbwOVFigXTEJXp4RGbc6/NKUi
EhP0yt7G1b8RNfGYM3l5uexP2Nk9yYuH+eVSlscDB0rp8t/2RLrpE3iDizs8
1K8Tvay9OHpTgLa4LU0Ak+r1DFMKJTsAyhbqQibEM+1e7auNbeu5BpUGCHVm
9yztj/av/1ALqbS88LbVuYHfBt9uAyHH8eLaPmfSQ6B02Yx4wBfS4OeLE285
GHFHiC6INOKd3UXz2GVTEIA7vH8vfYfD9ZASKwH8zn4K2AaXrZ6pS5fBJGpk
qEhubjOk+fyU+RZXQX8zA5D12SP7o0QPe7xYJ9jkspSD2GWQ45ZGf3nMNNox
ICWi9Zfikgw+u/V312PxLfYMlkP9srvKy8t6xEjOGN45WeophJKw5vXXJoeb
8hq4xF/S3/ZAfVSgDVCbesPu/S58ggpyPJGb/EP0jXh0HtUoenUywwTeeRF9
MkRJsxw5Q10+/ag/qyPTRFJtORK+EXSDIJ3k/fPBUmsRpGbPJUY0Jwqjnzu3
UGorNDuDzBUzToC4XLLQzfqIVKI17SLC+VYrRks6WJfgmNamo292HitNgttD
61yiJUHpBt+DXwZsl+7Mv+zMKSY3pnJQbJJxEpQdudula1bo6QS558+bR5+f
thwCHh/0aOP14+vlx+t8lxkRJjHCCh3n7Je2QlqsKrXFgwHuHbZ6Gtd76ENj
uLh+XjVx922xMUr4pDsqLoC43OvSfWcLqOva5bho1Biou8LJgYocquTi7ejn
NiSdfyzfqZGFmgq9oE0vbYBJNbnp6aTI+PDHU8C49yzKK5s7mbk4RIWaD3vf
fIx6S5vhxcyOqLbF2JGlSzKLDk4KgDdTIsyfpIDIuXC44KSiPXtlSsget1ul
aLgShZgzChwLJwk2857AkEZ+wnZdiGXPesabLBF8jm8Uae8IgqFcvGNP8avi
4hnztYYRHxhYI/1PleAka67NSXVnfTrhTdqPcZJGEwZoAEzSbCxyCXCFgsRJ
gXL4zw6k+CWHgNZBVEz/ToDFaTB9S/0bqMMrOaOKXbgB6CRwP+3RdKYguS/L
aUo6ZJqSB3827UgqL0AQqxwnJFKLwzGJjHYaFbMbLZobyMH+/znbh49vJsGg
2cVpWE3WckiOkk6RGTxnSwaj4hGLGqLYwpe0/T8Os94PbiL4TQ/7PB06C6R5
eMU5VSauBCYo3QfK4iobk9TovmSpvvnmAIjAzlXMaUWYe/a7XifynuGOmLEM
fftL/BBomC5tSgoN9r6RM9fwaP2BPSsn+yBSvUFvufhzGZ7KY3C/eR1/11e9
v3gg9UtMqf1zAfqbGpNawJVFnn921VV2FdyabrT2B65Owf7FSsi6WVM/RYdn
Q9LgvOxqVT1OgRMer1q4Eof0hPrlY+dC1OkwUyVV942yPMivvR9Cpl3OXY4h
wF+UOIm/HUeviCYThw3sNFe8LtppC8vA8MwzhEJX/TREwYbf97qnXKStkd7M
AiyQ63eja9gtKLShVJ4qieezgzsAOi12YbmsRyzGItgJwc3AYNf6p9MT7YiH
hYo44Fop8RV3C1dtQeMAH2Bl64krjUqwPLNz/i4Vfzl0rDUse7dFrvwY5joE
r4aw/fIt1DdD5byImFB0qijA/h+iC/2WOVXACGFlB6AGkO8hMdhAX+v1+rxq
r7SqlT4TZ/BhIPYzPsvsI2wgywX+O4abmxysw26Ctt59z4HUICYM4Ao50wjA
8Fy15miJ7hnnh4y7JG39gc4nNHbBqyYwoYWKawZ8uEwESzJzI9CBmSp1PW5O
teAEi4fIHIfiJvAhJFZobmbwDwg/2+d1IsZUheZ0eT0ZsECGpp1QA89GO5xZ
FPAhjUCI8TyAmKUYJY5LHtQBuczw3Kj3A9a5K2IK3P/fzEfDMvKQxHnONctR
AJpQ1kGpbfkZkgmW9XQirvF78ezQAIHGp/6hUnB4LDbAlrXp6VdxBp8HFk1P
RwOAAIOMzDKXWFOts4RlH+f6GU0Cudw/zYSmRc99CAT/F9gUvvar1/G0Nmmk
IEZq11OJBZp+PRiEahrAYFd1Vqkp8VYPu6x3qixN30bJVKUB/6K6IxNm8huL
9oJOislYBaCUR1PpwaurMSTF1qQovt0MYU4XnWehItaCU9ewje60hmNXieV+
4UhwW7yqlUu1GPm3BXUNlVrmBRx+CEdIhnNNYf7+JjjiUYShbyXD0d3C4WKd
Ty6MBJemqMM4UqUtK0Sl7MIZPsHArOEEd4BbtFkiuXSMYlmS3Y/ZaL3i/+FO
1diC/pMUkHpQZtG8U7EjsR+Wsr/lFrp80A4nNrp2aPJCRlvGOLPumk+VF4+r
Cjg8fK7rhnOCMOLG899mwbSNeoau9zaJYPGGWDRgAtJKpey5twrXtcCmhUdL
+I+SM2lu44516l2Ye5MlO8zEGY926N4IQYSZJZrP+KIZn/O0PjOZTcvzOMHb
ktCHD0bVnCdkZCHbcexaNDvc94NYEe5Q+UEgOou2OT/R6A6snK9W1RQRbNfn
yvbpPS3LcqqMOyk3DtAnM222T0AqnHppEsOATQH5IyhdEKuMUoVt6Bcbdo6G
VyO/KwzMqXJngrvqEzc5P252Z3xILufe15R7F6uR6iS0PrgQR3LEk0tCp5E4
fpvfP1OH9BgxwokBpdJJ8HA2gm/s6QkLmfpI/THoe0tdbRMXqpi3oerW/dmR
TNKqHgdBYx+Qov/KKZl3y60iXCpViHziv0sLftJaoyP22+sZfC/a6INWQEjh
l/jEZJ1CvuubmFStiyr8lCO6wHJEDjwmIwExRfa3KmkSDpyWcK2YhJW0VEVe
PxE2pQUVjAM9x9bkjeVP3F1RbYNqsjIrOQe8KGF0klAgTal5Tf7+yNclvmN4
BAY6WeWa9JThJjmjlkPks5OSj4l8+mrt26eBE0z/vFmG9knvLH4sxqj1zoyu
s1TRvi+HTofC12PkNQEY7L5XJTiT/y4rmybPvc58Uoe1J4tO0t//gBxYiAC2
LKS51WEqBx1Q0dokF9NMC5KEUxG8LYJnXd8/ujMKxt4M2IMP+qQGIHw4IdFv
9ISpErhwFLWN12SoZ9/OjIBnE377UtgQAuHHKPSR8PhFYGbngWdk1Apx/Uoa
/NxsF+Gg5CJuHjw3LGXztZmUm6AOCvXWiofaIaJciYmOioxfCqERsYLRIuoH
QHSTAEetjbes/cZih4ngnMPuupnHrhf6av1U+ZL60mxDn0FVTTmyLiFKwggL
8HXqnNwtN5JuWyfOt6WCbTv3+YLGzHRk09VfMTJ3H3DxE5aQG+F0elauOnLQ
+WELaDqxopr7vQf8MEr9fFoL9ZlEA2xvlWD4OMCIOorbJB53JX+9Htk+xmZ9
ioxU52OhIgI9dLPb3sj99nRrA+QCZe4T3EAuREcco4LhL0V0FaI3nAtD9Zkp
Y29b34tYWkks6Idg6M18iLJEFcHMZ3mGyQ3T24UgYq7JsknUwN4vWCYtjkzm
G9axt9VVXuUUCKNtDqbhunb4DEw3Rk63DAwad7iYZ9iWf4pmedCbkIBu5a5N
t4O/2eyP84jbh/wmCvfQFnwzeZdBRVRJE/IDIzcO5S7zAcpB1i9xNjt7PO/l
hHD0DAtRPXhSaDwNnELYMJe6rm6bgm8rQgs7BTyxdACirokDy5LNzDX6e7N0
3ayRiiFWbj9tUUy8Tx+YrMU/fxWb42PR/A1HSv1SGtOc2xJVQ38bHjtyaKYV
BSX9b3OMeqhrJ9ULt8ON1mE8Xy7CZda3wqVVl85gP0ea6LITqNbyy8uyu27/
ESXjFT7xkt3KSzSmpz0jaGR5Kdcwh4inyjjXFFeNoRgGGJT4Si9L+wPKZp6u
Vck7uSa7qHX1OyAaRGFORoBGNrZci3VqLCVQyu3JBh3YBq7TrQAkBiedM1vY
OclTZya50BkXYW1xvm3sbM1oIRFoIxHdke7gUH37fE2pBXGEosA4roeNbEWi
1HJTkJpn/4TKVFO2oi5dABgAxqDUORs8xc3caqCXkDRRBVRqXefVKnM5LG8q
u14cwwEFD+xoXHmL7Ee22CaruefpwB4ysx+HKbDkwQTyjxrPQXIbD2sP/3di
to5nyx23MMMun1RbiarVBNP8xYVCONZE90C/Jmt7ifsgV2hFndiGv9rXxCpW
e/A7zxUPOHTg60bQ7Z3wEylLrsw859m8UStXzb6GL+e0ouG7e9OnPYwQx8fe
RrVOX8/X5z2vhzkURqJfv6iBnYhXzgUMP+VpXZ+vbG+XNB9igTKvCMalJ0p5
iphqCvdli1w40a5eA9MG/Jl6GkQaX0lOQKl4AkAWvtXG/v62xBbp8aokGBBv
rKaaSpEkh42HHsgMQo/udU5K3n1+uJc7CYPyp3D4cUeArZdGifGzu0Ow9D5A
cm0KiT2tI/TpkgfkL5njUG/3s3s6cqDFMc6NYWbpi2nZ9HhJjfyZAYzBeY2B
pHR3Vy38JDzcm+OEbx+Ca68IOZxEWy4Z9LGLNt+TmJ5lu1e5bag+w2IWPLfE
2l64QwjtQelIVb6UL9RDY0+NBjGyBOLoh+tBdQsnuQqjxev8jNNNSteSTr5e
nZdSvOIKj0DaUUfMjhNubznwWdv2xPZOfDSKFC+srWMSFH1Hip63LkrhELsQ
OQ/bviaVXKXZYGIqJ7hypCEVYJ3mYPyBa3EN3QYuxfgnPgBKXrGKqs0sUtuw
YtlUbZiNyOfybRr5aq3UlV7tLFQTWKLDOAXve/k4r9kBV9jKvw0SE9REKQCY
O060EkP8p5I+xJyc46DfDVIltK9bk2DM2mJGcMpbpXVj0iAQWbopmwlFzhE4
oR4ocIfaRvn7TS63H4h4UliO8TMX1/Ov/n4Zz2olbW0/oLCWf93RBH6XNUlr
Yhi4YjlffZfQyJ2JnaPWW8ckvhusSG3mTo4aBp660V8FWUCT5J8orywUosh5
dFrzV+uvFa7ajxIHH2vovaloM1SvKUqz69SbPffPDny9v/mAixE1PTlsWHHF
RxvswfbHUO7906xothdcUUS4vwWB2zA85H5FN8URyl69MvHvrZnPk4WvNb6+
fPqpzsMD12qf4JtNkNxANfxoSXYpYN+ia2ImkF57az2oLUf0OjoF/ZB4aGb4
TGdWzKcdpu2xFg9m2L0tnQT9lYDncwwqn3V/GIvY+I+risXhGw+3sXtx4x7v
wFN9FMEBZ6u25WsvFbv07Q/FYW9rL7q9F07Hx00wVva55R0GsO2i3ynVIokW
cz2kk4PHpCBM0pGkq2oPmMGwdTC2pjkU3Dcl+pedFl/nwz4VyDrnu+DupHlL
4hic+/j+e0fPSqZg1Be6hluX9rf7h1wkXJMNyOD6YBUaV76Aa0twL/fKCyAW
/1aIG5qCKRXCmqMM+C5ymwDUBIE8K3HGg+FVvEQoHWHPqZ9brn8d7n4EB1pw
S/Ya3FBW560o0+VGtOYWa3wn01Zr+crC9EBSZ8/jNSkBAO6ASolQkC9s5K0u
rc0klVsXErn3MZK/+zokJv5VW1L2gI1KBgHBZR+SYjFZjmVVcHEgA0KJPxvy
owG3pVwSlMDDtqcupYI2ADOm5z8UJhNwgHoJMKZEVda8zmq/HL7a94vOeMnd
H/ppBKB5yHQZ3IU3DMgfprWDigZqKa0me/imodKpY1Vp/cJMLw18excwFrng
qNWdrhPxenDs8n+CjC1zEiB79fA5BWtLLz1nOKK0qU7EknWw+V2rkM9xUE8l
y6gy2/31Cqx0HRC90c5qzoCMZApR6bKBuHucdFpBmPPSvsOJp54aJ1syDD9D
hZjOsElFjwmvfytjdtomY41NZfxs5eNkraIvI+f9x/hZuCd4f4MP/BiZ/YOj
pqIxIIXLFO5wOjh1/yFZaFweFDCl9k+j1qKIxSQ5lzTSTYXCpZxasxTSKcQr
taq/Sydkie+CnKQRGZkdMAQGUs/XC/xwrfW5PMEqktCTHuSUdWcs5WrRRJJH
fZyr7VtjiGfXHlDunmPw7QOgCaSQ3RC7L6SBhRL16z5G80FsJglIeRrfLMFw
yNWZs5mDsEyXig7goiqS2GAhP5GwJMYQcTy7oulIj998pZy+BZm2szkAVMMT
kquP+uACgtN3tSttjCpwa0dygjYwN5LN+avmTxvvm10T1dpyVDcSjpTln0Ze
jM78Aj8cNiSnsSkMLa6U5zXsp7ivt3lseaxd+rspuJWnk+s2j3sKpcrvzC4d
zYE1PsJ4G0vogGzG6mEXN67Wj53FaKrKSqiA0FyVo9A1IYc30H9MM8JSW+1v
cm1ULjHMR0GX4PkRzh54VpmWoFtaxX4IhGatsGnCDJVy3vXSHCvHYwfVj0bC
p5JUsTz6viE5c2V3i+ZRxoLuCu6Q4NSz+qHITKPtV5z4o0nm+qcRz4V3nobE
Z6wAl6Q4E2aZDCJvlr2H0q4mJUQt1qKgnE8avPpIa1v7sDA6L88E7dI+Qyl6
pbVp4zkYYlnceA6fufdcvEPcWfLXtS9AwS22zqH9B69F8l9Y2WlkhitbLN1P
uuzTmjtu8ZlYBQKBykNoz0ozqYaWM2NNu25LqhhTCiGZ50FLHWZEYLiUllTH
XIiadulr2xRte3TIXMzwChxRzXYIzzLZVSoDSnDCdJb5U3D6KlOHREvOU3Zw
lHztyBHWJKlE3zBOuxfZV1B3U8bN9EDgVQM9Q0wA2y17BD6qgha31kBg12nE
2HH0J/590nDN1pvA0Nt7mjJjOG9vzPgHVCX34xkY8LybP4UQLtopn9FZK42y
Y8TWGE82Om1CpjedIz4p/TlfXpY9QVIoqXv6D4t68H2NSSNMP8HClcNCyzFi
OQ1OssxyLFuebBlvQyaUucBFWlXUVMWspzi8UKT0CA2bFiE78z97HvtBA20r
8goTpiiRsqTZytnacUTBONH/U7lJZbN+VJpcQAZU6BiCPNARc7NtW8bF/aV7
chFYJtijmtskSXz4AhLAckCnPwSSewS4gpMtoFNzoKSgJCWMiYHrmOH0ytRj
PFsHJHioD6yIO9EZFUekz2uYaLaBCMnFCQvsLG/IIC/bPHVTJhraiwjWiB8G
4CclDHwQbuYNQdRXBUE/3TgHuvstAg6HcyjNkFFDRInK5gm8OBjD04msE/sB
8caDtRQHtqjXwD/5xuh9H6ofDCs6aZ7fmQU1E+FfQyECy1vtu7iZw0Sv/jox
8YPM4bq7mgzU7MlMM2i2TTlvZtjMNqMjoNgQ7JFBTSqI1NnqxNuYkbs+Byis
TRoN6i1NeWE/ciQSUhuwnljbRCDQfG9tLzlPxkbg/4RhrafO2Y7T4AkENYjj
NfRuDnTFcVoFzUKXGQlrMp5yKQ30fBDb1RXe06Jlcn+k9crgPgKweafAo2NO
+RLColo1kXM1jgWyolJ+AUVauVnfpu7MNdZNXbFZnQiGq2hh0THlB6E4FxUy
KwYlcvKUKvxTIRxVKOwgfUSom4SA5wZjXDUMLSVZp9cHEhgAmHXo9f+xKBO5
qd+Sj7F9/y/2HaL3Co7Qz2Qtsl2ZEsPKCYT7/fBTNtA4zkNSea0d+Z4dK/Ea
YgvtRuNVslaTdMaBsIBZhTOu94o70FJ2/HSlQgiGf3Zil39CJStJ1ubptPby
AJ3Zx8JuYNsMTNz+0NEESLQeiGg2AFahh2jF31POtb+lUcnzNiF+xopgChMK
NRhNT7I2ScxxNRysxsMpj2BAZ/RnnbUK3wOw4v+63xINGg2GSCH21wqAZYhR
QkZMv1j7/BUN2pMIFPWXBINhbAR7TYs8WtQ1mDJYzzyft0dsS0QSz5YgNyCv
fkTyazWgltjv6lbSkuxq9NQFw6DAO6RRP0UskwleSD94wWeMRQPcRs00be8y
+c+zHSy09noUrPWU+DAkD76sjPXOIA7vtwtRvS+ZW4X8wFDs9GtRiBtl/bw7
SCtqQPOZDLNpy/DViIfLHToOg1ES+52jpusPziiTTI6jfe2rDZZimSQ58KCe
RKtZxnz10OV80anmeX2H2ugI+9PwF/K+RnfX2gJklFgzbhzlY4kpoZnirzYr
oa6dxhtg8vYQq0nFeM3YV50jraBJBXRPLFq9ZGyz/SGOVOARtZBvKUnPYCHI
GWINgHnW6TA9BsWNsLiIRb7kZ2ghk9K+rNam3Q4WpE0bDKzIiL6QFo4ptGFs
L9MUZVIao62UBZbIVNg3gcVpsrfJV6ek8fa6tdjkMUuFCB7xjegpFXqFeU4R
lqoep70f5/Gnr9oZ8yOPcrsgc3NSwU7X07JvhmeA9A0AbnKwor+7iqgnjdsU
4QLtATa65rNGNBfxiStcGmLE4cmt0TcBGZeDKMU/C07Uydcxww/gFakCNuHW
7O8LunfZNvGX7pAxw4/G+LMHn1rJ2AcjKFLO3o2MbSYSv57zNFBqpQPAquck
02F0o90msnG7U37Sz8FuFpb80RbOxq4h99BHUqOsOP8Ox0b2T1aSot9Pdwbh
eWTkmUs7Mi2d5/KdeJ4p4uqaDGtSfBUM7FVzeNzCQO5ZjgAZU/CNm593stFH
AkiwTy2rekRJngFyBh+0OSrf4tv13EVf5joA4YPF5/DAeSv7yDpmjAfY4/cA
n1xu4W0cFmp3HK9nGuV7/K9Tt31AAqKAfi27BP6bhbq8OI/Wn+zyLSti5dbF
Vs/ZgxZA0KeuJorCLZOiaOFu1UB3iX44p2RzBg5iYtvVi5iPv4DY+NbGdjSB
kUGv6jjkbsE8rycOQlhP7THLPuadMb7vlI4ZlZfCbGV63ns/+pkc/6F2bpNb
Qm0QNOp3DjRgjBgj16kDIKs9hkjUVjQMD8ka79jDpFpvIJICPaDwwPjCOdTI
tvChtMcaD5uq4zxgI/M7P9hf8kcXzmamVTt3w1wFe/iJyIs6PAlQ6fuoDwjP
6ZZ9XgFpe8WL6HkQapU7LAXJmygYQSK9gsBd+YzXempJJW6J4/5xIuv2uvMD
F5HxVgf2rX4ufeY7N3li/X1pbLatRd+yxlpX/kTJyZgAmYuaULfV4OuKSzGj
5R9WZWEEZU8LhS5nmO0/BRYQRkLh2s8B5UT5fY0+A0OAQ71LYFMReNVIHBOj
+yYA4WeYXtLj4LrAWzWCI6SBdCnzBLEOCiFl869jvyVYoS2m874uNJSq2FCy
CcQ73jc5HkEZw1EG7Vt5uM+DhVXfihwWrGurQghYXk6S/WaGrxtxtq/EieQ3
MJ1hb4AJKUKCXRoZ1mEWUdtwpTNNtBkjTuC0aN97N0Gux8rCiBO21uFFbDyE
Pl7/zcRS4wVI+HKrUdRZ3vRNHn3bvlQvpLdOpJHMmF6kgReUgPQlBjvPm8b8
brZQ+U9LSRkSa+67go7FsYoJeyZ0ysSf2USY5up5oxHVgWjfRyvv28u/MENj
0RH/up0zKPlaMUPyBZFIfEFE+6IdJIgc1Aab5w8hnjiwTydZT4DkSWhPYWCi
NmEj6ddZNYG/7KZDSgb/+WW6NrYVn9pDYi+OzqRiL3XLMa5kHYwUdnVkJEaZ
6kz6S9ETz6X0ywf5MRMb95ngkLZHQSi2gThhu4GP8CbrWVgr/KcZVlYjuBgj
izJkfxqFyQTHGJhGU/ajcNzukrSN1LPl7j2W/xxLTWw6uiOr7+yTH4W6opz0
TgUuwflIxGjhK7A1KAItAj95Lhhd2eJXKJb16LKWCMMf1vePzzoIk7AOr8aq
I80XdQfZhGP+qb3jpuHVzWetgfQKHnXTK1OOzMlJ4IWev+fsf/FOEOB7zQdA
SugmhAFOr8jNvmYGNBBkQEeblHDcL+zq9Zfx8iV7uK/y4ry2ShNvWxqswxkK
7jolDlSp9RvMbBy2zOJ+4WaXWYz8/HtDHP4zgogIL1/tpCs9bJ36TGlmQNp8
qIzGlzCEPygbQl+w40krcgk855ub1ViWszo7RkQwhOqiqQe3TBQWUs9MD7st
HWahEMgtk/sI5WV/UaUBdf5reWV2euWEwENrsWNtwilBSQDY78QH3Avm9usX
ZoqQmr8t04L/ceFe/f1hF3/jafsy1I7JbgglgX2ddzG9B11rEuGTuiyo9Myw
rxwcX8wWDCHIO8tzg92iskS0i4eEaHjPFCt+WosiWoFbA15N7fPT/W8XZAjW
7QI6CcaB7GWtMEOhhh6jlhdnxgm0CIA+JoUhrvwfgp6rn1o2fMN+9aP3pIbS
Tp9g8agEBclIuK8n6r/X8yFTQK44gAUYRfi8qhjj58+PU1zLF83fkGg/VPEW
aAwg5X6nZLug/QvUhkR5od4iQjlBxCmfArZvJZM+NcgBsqoW8Yv2Gg3ZPEwo
TwG1W2Ygq9UM+XYXJNPGOehH0KvB8SzxVG5AdEU0XI9sFgMctk/Sp0Jio/sC
PpfkAp/YvtoE+ejhHY8pAVM/+3SLSnA/7huxjDdlvohKDcYg3VhtMjEro7vX
8LtkoX0MqmOhAf1sEWIaQYEe3ovyLWlumsH5xcLIzUVEfIRmtkJGIrKmaAdO
ueZ8SNr48mOaR2QDX5cnMtl09vFbT+LsjkcD+vrkhS2zjzZvCMBW7l7pro7U
m8ozY5Ed84gKN0xPrASQ1bog6Wc78Woy0ar1oN+viFA+9iHF8chL+FksSEey
Lr0hiTtp1qgm6W98/4/cD60wbAOlBw1JEgaouhFn2BTn0Vho+Krwm0wK4/Mw
805xufgxki1YCxV/7OY9Jm7GFFKztSbTuxsSucG7xqbr1DmemV3Y3xaeG0rO
roqPWbwo6hLNoGzZkqVyqXxX20NmVVHG8Zu8KmoHhEEZ15hfRtCkzjRoaPjw
TI9aXfV99mGAOX5sL9tw28cvrohn8m7WbBV58yzvVZ8B64QIRZ4ujzZYPKML
HYN5XE5v1AuUJdpu5W4AzaEQiTEy3w6Q8N9bYIh3J49ThJvUh+FaKb4gunVI
RPTAMNIWicANiWgj

`pragma protect end_protected
