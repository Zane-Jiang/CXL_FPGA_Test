// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wsP8DuQ9CMd2Ug65j7G1GMYrse+JKxSccZHPf+P4Z5Mr5ahCXorD+3dXEUvN
prSa5LyuoGJpW50uFaLjP2wqJBOujeT4EJO0g8sz+CepWNpqZWt0WyIsUz3F
vrqZ2Ny0deKZMko0mrJhpYF0NapPHWs3ZU0BVJdvl4rdzkcHjAa5erkED1At
tOJpWVtPZsbyTJOuGRRpy3gz7LvH1bUHx5M2KgxYwlDByRstXkkQluCrwlIQ
Q1kNplja2pGEwPNqEpY7z3vvAJnwCubrXr3uFrIFxTsBDzYSs8nU55UirRkl
Xyzuzaa2hYm/XqkE1FghSM6v8fJ+Uqsz0TTS7B4Iog==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cQMcbsOEZkfIZVmIfGEapgVCHOqvayTKckEUSjKv2aMJJK/wFQ74yX9viSt1
Pz0xwf+aEHhtxse5aDILzZuaa63nzJjz+XVMC5aoT4wFGpC3jDUBZ1bAir5/
011la+x92a1mIW0CU+GWFGplYMDrK2ATL/hyxbbHiuAIsI1H9ZYlLBlueD2Q
MHw5Rydkr+2SCZJj5/bYEcMuR4zMNi44x9Pr9gmr6TQxjB256l9Z+PH4ySg5
d1vq7wmV+zdykLFWP3nE2sd11pCXZI3FhP/tTj2dnu9j035LmfDpQCk2LN02
XbQ4oUn0HXcje4KAXW2zxVdOjqxUHDhjwZ9Q1ZiWhA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J0VdKBTdYhag3g1/6ZcQAOrBHpOu5R/ioKJ6hNOOGxl/l22swTNI5rYwh7WK
8TeyLFO7jcj5PNtm+7qjxQuHRcKMD/0aeCMnjjK5fypb15IqYnlxywHnschm
aUXdL5HTQtudJ9eQ/ath71eFuBTSV05/sN3IO8K1EZN8pEP5mAOp4pJU0mUz
Zia4WzgnVkBwj0batTO/QEyBhyuf8ULRmlsEhqJzl2nXuIZhCatokS6lJGEJ
IBcErm0PP71XEFN/4yQSlvwtcoO/iSvFP5al7u7A2wqNsvI8V+2m7V6yhfeO
tFdAMXITFwO8k61D8HU6Xomf2DGAAWl6tqTS++dT2Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n9Vdl2NemQ9ZmC42BIe0TfsQ9dxjXxzZubZ9aB1gAIKueR5eOGZ1/GvOqpsa
O4aVdpEXAlVtVMOCWdTzSkxEy/NoA8st305FPb5+FzYOckrTS/vbA5xA7EeG
C9nS4I+uaep7Y4U5DvkjgLydaUiW5LzIQ+ZM0zu2bITtedkxfrU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hE5Jlwwp9nEn6gYmZNtFXRoU7wM9PlizllJq2VKGNDvH52ODjJm44NvJuth9
S2VSCi8AZgWpJQNBR2rH/Fcxxx7o6H45I6DvEPzLpGO4MgwWG5E+gCUKxwkW
UV7xxxffErvDUi6xMBDdKCTODXLDDPgmuqZBY7t/Vcf5+yWpebGOPqNyh9jN
AGg8NhfXBMdd7zgvziuiit00z436+rFzfHIxVBjtHUfMsVwEvWD6eC37JHA4
RIKpKuKIOLRElhwV7PAhBYUH5KrhoBVs7qa0S5XWSW/FmKgtCiovY9rZjLMt
+b6i0iArYuNHgsuGLGm6UJ3GOP4jEsyNvaHj13RFwYrz1WkMtheuK1FKdxo4
KlgLTP3enTQmU6Nv7xKYhp8xt+7UUJ8oSIy7W1wNnrkWXdD/F5bAUMZzymFb
Dd76Tyak3YOu25WRt7Ssa2Bj4T/PqYEH+LUs28oBr6LH4ZmLO1XuEnF50nRB
Snan88LVsbZRz82czOCZIe4UxQT5468q


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HLtc8oLM/NcXod67iEIdXXrO49q4yTL7BWkwzVm6xtFI+uMfEsHD0SV+r9wN
VIIac3p6kDyl6armvZkXR686s9GKQvjcrjqIbobfin63sDcTHejIFXipNue2
oAz/XIfXbtrM0zkMzehlIKE3yoneOo1qsAArVkUdwJIdPJ0iiog=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rHKHYp6vyXvRwjIwzFfSeYVLXnXGRSEgerYKFbpaJE2ooQGfLuljwVokVa3T
5FTnvp7iQNcWsfMWUaU3/aeAsBwQXRRYk0mBY+5gxt7yv+4jaBda/JG/+sPU
cFLshkDG7EHio6JJmxgb1H+9oCKPAS/VmRfSOQGWcdR9DSxdsnI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 214080)
`pragma protect data_block
bhpl1vZj8kxSEhSLdZVjCAd4veOye4w3BtpQYl2w+bj904IaAf94CkSRLia6
T6UWfTIxQEZHOnHaav6Pdqp2wQXnlPVgGKK0j9OZfGUZH3liZ4RyaZXuAzZk
EawbqHHd9Rg28sNpYehM5lLqutwGYglHczkYNU3c5phRcY2CzpZeWwBCcNYm
v01GyJ8FceiRpBk48uxkAdpp/9u55xBFK3eL0zCMycZW5esVXk0ghmX/m0Sp
+qAMS2iYjv/yAUNXy5ZCYg8JsR6mtwJvLGBiQKVIePEL/Kl9yO2VX/kDNJnA
bs7vKjjqzgVHWuAqwvUNkhEdxbRhLmCmVSauTHrbqq6NQx+ptYFEIqchz+SB
YDKcYM/iyQw+gohRaeA4Pds894KwfnPAiTK/8axfxNxnCkbzwq98Szmb2Ps9
uWIglkLoOCqUMOIVb9RIWEBwNsXDmptd5MXVu9P+9Pj5uDTD3hlqttxyIAoD
p1Vg//fmo7chaRyGjJTJYcwzzn+XAEcrFIDWpl8kWCjGVOhYVdvnsjlfygT/
P4/4lvzQwvJGnXDRQ3oQptrtgoBKwURuAUOEEilJMWSPcHQ+rtUFkom2y/Zx
XlcpCgj4shawu0p1vdC38Vywfk7j8ICgssyOxCrsgiLgrJxWqXL5Fn//0Lmp
fu2uG4Mdrqzg2ZWy7cEMBwMOY+D70k8J2dv3jjt5F4Dk3VHAUdbuDaqGDml9
kYx7L8a7mrVCUKkLzhU0kkz10ANLvXNlssC0BGpnM3XeCz4tnooZ3Vln2mWv
bKPIC1el5MNeKfzNUE9ye0FylQzkK8Z6ngV1cJzUzK9hpN1Llat6k5eVEB1S
nNNaHNMUZBmfv6IgalFRaNnPqaCNYRrm7nYHFllGjKTv2O0zUsK/c/LvtrCX
ZqF75HdrYaUeBw3Z46ULjdcKLFX11/DsAFfATv59AQ5hntICJzqXlIZ0AaPL
95VzYkk+LOV5WLvuvlpmljxoBB0J4xT2p0zNuQn+AD1X+JeTCAyf6eWxXAOJ
+vm44AQkeVXzOincexIRRuGeoOxbvfD04iPOqidBfflVcuuaZUjFUyNxzV+5
UJYg0yC0V5lPkzhymTzhOEDzSdc7M0sMroTTSkgjV42eXGJZXnCozgqQtP0S
sGmDFS7HL07XHWP6ngnqX37gIvDnUWsW3UnkiQvSpQIg6qi5DzV7kJY4toPu
zrY3krxBU7QLy9XnsXcVai8GO2TNQeDuXBljH5xOPtW3WM8c9gyl7TEEFzVe
FDU0CrNxXggnT/mVMuYb+N9FZMXh1DEE/EKeLgSVCyspBbg5ive0TLWyqPxt
revEgn8JQ8yr/rmgB+QVoXEl3gYkC87eYp+5+16QDdMJiiShf7oIhNXH0sUF
NJc6NnNVEXDSq+9CLEBvvAHpDA0OUpWnNW5quHg6co9DML4SgVEtq1wvrl0S
i3MdAMPBxr7kHC6oRB4ykiTzjQHdVQr3xSoqis3Oq5xCaykIC51zGCMFf7Tj
6+kOdB4Y83mMI9Cvr8wjXkid1KKGamxot1HRywoBSbrJ87YL9OeRYlrqy/zp
Ku20bDwP5rlUFaROEgkFLEEGZWgRCyrKIDVKqWU582wVtzJ/VZaBfHpshEsu
8HlQcyheTzmm55LE/NVfopoCgM399tzlmOYUG6viiF0uKSkxFJm7Yy5YBzGI
tv0z9qrRD92sLNABe/n2qmzZHvxNoeoP+ddpp4yGY9Yo+BRKlPJt1teL+EfN
2gZUPnpNFxLHmSuZa7PqGrbAMnVyTVlJCHMcCkunZBIzcpcO8Mf1i4JO/WA2
mYFl6vWFYKELy4rBIidaZ1pHefUkUUsyImWh6IepNZETsZz6K5v+c6/mzkL7
ogWX1nEyHKt1IU+HFHIP7p9IQzZ82CiklXIII1RsLJVZUMOHts/lnI3buoL5
8hkFkqOJaJa9j9iAMBweM2oq+g2nUQbXhep0Hvh9deViLfGHeReQ6UeHh+Bq
LjQbXteYpRoWy6a1kcukVYECyoWXaMWcvJ8ejxx1aB2PfVigmrJRtDnizlKB
lflPhzdTQ87EoOU4+8FhOBkw9LNts7vR7aiUoYBz5jkSFRASlBUNJehbPqyw
25KtKJOhirgHInc/duZFKw93UrCliqhLnD+mfzOr1GWAA03H4Y5jiKG1UvF9
DdB7ya5dit2KD4YQJIGRq9O9DuM/rvFQqHwOI/wE+1dGhNXNRqFjUhaD568T
+yjz9TnyXrnntheLiNAZr2YJSM+43KhVUZ8RMmgIf7u55IXh4sHONZCITkx8
UT5ikmcSjOVQOmaYQh3b2JnBXkoPIUyRBkrJN7kD2dvyfqRneTo0f/nsi5Pv
wFEAS/4bYcGlNgiJz6UJhzknJYHCxih3zNlnQ8rYzzum6jZHClB3JV0+yUAQ
RnETErrIGP/ubOhO82EZPuSdkZ/ncoGAdJSw3EnZ6p8Hq7j1DXlh28dv7hCR
FmYiwKT72w18R1LtIIy6aIgm4avaGzTEXvzqgN+F+CEquy1ZIUPjnLzfULyi
7SAPQpgYO1/n/7SfC60ng7mySS9Ofb9D97VgDkITDCeKpKeuwWm1hDzUFtzn
wYJBSpjlVaraMDcQD2VLcwxSBo9noOLPczSlt4e0RrMBo8BFzRd6NojxzwNR
G92VJ85pWZPA5uytiY2XbocnyBm30qQbwX07u0jMr0drkG+PNRtrlf1XYOV3
MK9J3qNbfdBR0BwhugvMuko92fwMiMLTW79KaZk4nmr9avOxNPuznQPNdlMt
VDY1AQbGcoA0u7CTk8+ATi3YxDVwsmGbEfKYGXD4asu9gtOWezHz/Pw+v0q0
oxyW9JmZMIqBfZHwem79lBUzYExV3WgbbIWm5V6GvOelpQkU9XM/CP2NryVr
vBwlvHGzY7cj6zfKUs3g87ZYjyMJxW2Pa+6KIAUDzm0eboD9mt53oCmYJa4c
g8BEUt19oRQleg8bn1iQYvlcJhuUc+HQYrToONQAWytoSE+8leQ1kGdjDHpd
j+7lBtV9c9C6jnJLlOTR/yiKIrM4F/152LgRThEyC1/aG6dxZa4Q7SSMYfdq
CZXpTUf/t3oxxCJYBbc9IgFElIv1hL0JhdjY2r8ndhq5ce2pBZEuC/lt2UY2
f1RYymevKkkqEEkCI3GFDOc/1WWr8yaeM4dn+Kb7uXTZNP6a4Y2PfHskutnI
8p0ncWYAXiMFLt6UNLxu7BvqruyWSxn7Eknann63dIn/ebX3bROrt41txKXd
QtCIrdZGb1g77iWo9amgaNjDY0dQxQBpaDwsdZIeifYT2CQsQRTVSYEJpQ7e
wa6yIyfjeu1JmvS4D7k6IssnsFgRcoP+RqMTkVvJ4fnjbfhd4lWZC4j4bo7L
6yh5InCbi7mSFiGE81zGE0iY9YB8s2+J3GQ68uxK/3fpxXVawdxWS4hJDjGv
RST3nwER+PjD43O1sgqLgfVqkiUi825dzVrkzmCZ4FA8wbIWQhvvfXibvqsT
Qrp5HacUa9qj7p+1sfhmmcid+JYHnwxbU8XZRNAEyTH7Z2BtN2QzuOy0dE0z
xyc1jGpwlLCttVhmcxdlMaaFK/MAum+kIKZSTNko3Rkv0PriDId/kkXeR6Ay
Wwi6NEVwbzhOCkGc0OXevC9Bjb3mN4XqvdqL4lwP8CtIAyHa/aC1fKpsobzt
V9BLHsTShEI5hNJHifIKipAkAtr1c6WjT49jsCk0G5YzWyq/ZhoLxeYCZUSa
besxYFe0jkQxkmdQgVD6yJTGykFwcNJaLBG3I+E6DMALJGLJAYS6qD94fiOD
16RttPk1c3oEKybRADCl/E8PZOz6mF/iA7VK3ix+NVaUfyI5osVxaeB91ryD
xVaQU5iI+rClB2d0Bv/b61G8ycr2+O4jp2WUdg/+mx1tc+hlj4tZ1qygk+9v
AWUHk5Plj90LW+HKVYFLmFYYqOoDYJb8awNDB5FT3QQ9o5LN/oiYnPO8mYCU
eD9cAmW5QKMQW6NT7rGFX1mGywpDUapaQuxZ/hyHOddisbuAdRce6ZYaAmaw
F1Tflxb7CKlEirDtat6YxdyG6xXCUeNFh8xLr4Hstin1pWKDQcUyutSE8eA2
3p0W0Wh95erO/9Xj9jhy0YlTKF7Y/xlyaZiLPOV97Fhq+gkYVx05zgxxe9f/
s7IrGh0c/RGPSDKQzARpd//QogswTZ8Z27bszZ6Ki/dc2Jf519MXzJhrX4WL
b3jXweI2vh/7yDPLozZxG7NqGO/AsgO8Ixb8dyv1bOOd1v27m4y7ra7Rlm4d
GLMHfX5/5nIKRh1PRLc3BzwiJv3CENOvuNHAY6Tv7BBMXQFC/dbXF8kzltS1
eAf6B5KhtrfB7lP8p8KjwgEQ32lQ/R+tGJcIszkUwllW6X7dbCmmSDbcog8Y
o4xxdKH8rWi9bS7JkbTJdS4ST1uHrxY4xjXsz2ESoocLxpLr7GndN0tTcgGB
qeS4viKkSdzl/RvqVlALVhF7W2KYyZx7Mh8urqZCqyQayPDOMqCmwl63Amzq
+OyQ/iqMmo6HBA77+Q3IyiJna4NlEZ6vprVjPwRq3vMxEzQ/+ytP0TTv1zR7
9kzL5/A2p8ov2hlE3WYOCyaqEaqSIZkSsa9l58qLatorcFAmZycjJBGnBxh8
CZ3ex4yFRQxdQYuQ54NERWyPs849Hf08JrXTFV+pn1vvcEd+XPyYq1yFWc+3
41iDaK0Q8XwrwCYdlesnGOkaaFoc9SHfet+afKHnY3rRJz09ftTauKPTD+eN
KvVj2TQLxRP4XnP79vy6xsTap/msRx2AYuTFTu0Dc//s/onQ4N8gUoLTW58l
lH24QItj0JuuoSLjCXm87SINmbbD6F4YGFnIV8/U12KPnTglV+bJcCE582nB
0YVKdYrwUzn0NYw3BPdF61MtWnHcmiQYKt+NNOUqmFv9jdIg42OOTmpBCev5
baMTaY6vm7sI14Idnv+suFXFzhOoqFqFdM6Ye2rcRpyQy7NyP7loIfdT3gSb
o3LcVRhdcMvg2osNtYT5BS3qiBmfDHFKKFy+QEB/yVn8mXaKjw23fGg/BmUR
6aBc2Cu+aSVBeBZ3EChp0JAKmj3yWNV8wou4mjrbrVkym1nIXA7edjDpXPVA
LdJ/nm2tAgkpXK32jhwSAMvFaesoQR78CLqTjFsPeG8xEDYqn/eXVvBd3SPP
0+8jQ+A8AcCA8dr37cqdN6Gh1BOBAC4SFIJRq5sRGaxOG4RkCI+bXoqR/faM
Fd0P48dMBrKumwyu8gppyO/uyY+oT3TfZ6IYj4ep6fo/lRZ1MRfWLj/85fZl
ij5TUOP1g5eRcHNQZXCyTGrFTUUbVMkjakY1E9X2757qNjruMeWT7SGNxD9s
WGRR9zDxwg6Dl7eVriyHo9b6fHol3lSwADipNe5+rBSBjfVer4X/ErgE+fh0
pGl1G3kaVJz5nMsILsstBVfDrjBtyUb4c8aAoTsGNSmw29XHIqyyWBrnkgPs
oppidbT1arl1mzsY62N8Stowff1+Xt9NjatHsrqtuvbz9k6UZsFaXuIy4zZd
r89qYe2g4SroQOlF3+Oyk6ikxnPnf6TYG+Lbt2d7JPeMEVGUSbDimMdZX2vT
r3VtBsOwryQYIK/96irUIwYeYjwAaEKwMNe7pz3BY6l12ZHvZ+C/KQBJyTKL
Eqfo1PLk7mf57MNo80Ixm9+evBbqAktXd8YCRjU+WbYQtktfOjvgWAuRNVen
Nqy6QM5hpAaQbZzabX7dUKlgtL+aeVCylQdRPI3Pdee5RcVrVMNb/zRuKfcC
sq1TDo8H1+kTTLmOUDY4LHssOI1QiYqtMzzpkBy3BqqrmzCUx6DXAsNV9kCF
/kMZ0HCp+LA42wsYOmGXnJMJ1CvbUwry7m9C+J8eebEacv+5kc2LC3fpqMRi
1pvr8fGnSysYZi1p7jrd46LVFYrFhZH7ObDIeW7KtaZIGffn0ON0XuX/Kd71
+6HETRLZZB3QsMycA/eu4stYVdFqZmSnp8ngk7yMG/J1P+FoW9GmqiMiI5/7
+jwBfZmQ4rABAyVzIBgqUqGyXJpzxcPbqa45ZNm+6RrZujHg5GnvecqbOF5b
43qbMixrmqTBfARyRi2el8HgTjgnhwhcC80tAs533/xJHxRPu4LWHQImPbRe
b5X2pF9FNkGRfsZTHbO7peT5VP6/cXyEdsJRF4tUBblWT+SbEnMnFhlknp1D
mrGzp3Vu1nPaZjb87z1koGnP/MNlERJ87mOra72/IWVCtdssp97xhedHNTFb
Ga0qfyw4hV2WFEUEjL48UIXSrK383lGvlKwGVB2hCNbgf1AqdRBuKuhfziUN
tR/PZ+HLZzND31E4Ve5ub9K9G9E0jvjzUkFNf9KRx/AuDLJWX3mArBdO8rYk
hA08sDhGNHJRBpZNGeW7QJUu5UUS2gN95VMz/nRkOM7tYQM/w5CM+CdovX7l
gK6b0Sv4CeiGOHA0nF8lBSJnWjN60n+ohIzAzg/NXC1jTPOsMKvBEefzC4/P
pFm9P4RJqK/T1jryEWgnqlX0WXwhJwSY+bcLcm3aElTM1EtGGhIscm9p6H1B
1xuvyBJnuNG9239GHKRT6FdKxSx6TxjaGOt50JZclBmskpAmWzmhNHEsdx/z
gQI/z7uYp4RCo3gI2MZQXX9SxVWWZ82QK1QppwlxwPma9wRmYDOsNUJ45Sk6
BdbRsQUDPkjwXNB95SHd1bg+4JZNdJFm6yMVM8Cm+E594+BOz+dbolHlccKd
670WRrYTmDv3P4BhxG6wVRfnEfpwzJe0eq/uh5uW8nbHog0/Yuw7yQTEHAqC
3GZEHA/laFaKWMgfPoJ/xzK/nyTPGbwDSjHqGudSsVm76VUAARBe8rKLzHUS
GjHX5ySSmgmflIDnHKHBEZrgWyw9IP8thwrrR+VpMq3fJo5dOo/aWCuzIVZU
tOIBM04PZSUmb+x/9M9DDxnY87i1GNt2K0rStEBQjLPgcp/Arxzlzp6MSbRo
uyGe+zNI7Yk85Y3U3bOPuFfnoabup3+RxaPJeMAZVFa2a1/Mtldnsdcwx7b7
W+hYUTf37xVi2MVZ+2gy8Zfj+2NtL0SkG5dU6gxT5ObWB1nJftpaq4f84Pmc
iU6xyg4bR5s09Gk7QTURifFwCrihXfAYxHYNWwfNygse3ZBUC5g7TghHfDs5
3t41ynW3lE4U9+2EsDKoFweP63vOsGHgeCK/Ex4Ltn+hIwV65Bv/Bo1vGkSk
d75ZxXY7rD3Xb1l4hgzXHaWfBPZhGkgmSAb1g88lV/Yu/vcw2C5zSGrLZ2MU
T6HoEXTtVSsUOveYyXvT3ukBN3veaJle/FOzsdr5/nFAIwuqnYHLyzUYb+2F
nl9eURInHSwY7scNZRBvtlFSM5eJcJ+4YeX7QJeKitml/bTg5RZut38JqWw5
8N8iIcUQqNQudRfvuMJe5IQjIjugAWG6sLRuHs1kk26LeFPAWAE4NtqoVMrZ
jrcelngkv8gdYVwfZYVX8rdH30LohSojwmurXIEXmN1/Kl6C79qUqBlMsCXR
cTN662DAdpHtOI5B51AIQXkpCUDz7bxzfk05r2x7HNTusArrtiBB17Kuivz3
P7tLAWaMZ2XVLwGdxDeDMI2efeiGdcWpr5SS1/YTFMnfoIgAgJSzLOjQhH7P
im5tUe8cJHtBYH4mAa+FYmIUQ4cecqAJFmFiTrR2oMP5NcjaqSO7/8+Ddc/J
nIwzyJCnAsqx9QjzcBHvaTBU2wo9Zbp2uFHuiCATLpaG5Lau1EsymLxPWVxA
0S9NVc05R2m84ZYcSxPXahyEfjWf5hivIr78MinAXRGdh4p/r7Tzm7q3XZAI
exiv78UNJFE1+uYAYMY22LUmoRvXtyBqo0h7x3HbWO3St9GS/RcQOqgGl4+O
muyf3iQlvVbAJ+VWaPD3232Bdn4OldUc+mPPWbQjm1rUj0PAJdk9knvXtsU7
nJe6jdjHJ39sw5pWL4LFoKtkijnHQX05MlzxQEoArqpGsnHTM8K8aH3v/QSm
w8zD2RrNj/fLR19QF43Md/ZRcXuofqf3IdoTu1SvrtzYGoZG9Mg8/buaAlnT
ZPSpenVF3ZyjmLjMgdDH0zFmgpAIodfP9IbR4TiHkdCpHxEnap6wTDCVRHgH
nhTW9EWMNORhd8sYTrMQvdbidJonEy4s65rIdrxgJFTDWPWG6yezfWQf1dts
YYuk0IRu6AnXA5yGHiDtwLj4em/d0m8k+Tt956C9hM+luBdGU5U0JkDIUni3
EvCMzQqr8pbtPBh6CZsxUNeZex4i7xXMBkivH3ce4G2uASM02aSxIOoKQNuQ
8+dXScUg3rHiBO6VqvJUZLiencHsCBFoWzbvDxxMyCqFiUFZEBXAD1MFIeD7
CW1zq41+yJKU06a5VXbLJ+GHCGliNVseuLIXae+wRQlxx/h2WTPhEcX/Qp/h
+olaE4WHGu+JBRLmE4doADPkic/Ix4OVEiEsIomDt6u3eztWBKYbvxeNK9yg
KoBGO76xSaTrVwijgqIbL3WXcpYICRDipOl+Uw+R8mMcU4IXCi/eaEg3TqI5
vqfYXmTMF5wQUnUrAxHme/jJCJ7gSCDlkPqtVDq2qFzpzeGnDLXlaFpZ/J/7
ahxGKccPB/82xAne42sPrRBRTZSJdA5gRDmlg7RgrN77V/xx5pHgOqkofn/r
Mm1W7HUfbA0e7HY6ou3imw7UzX4VoAjkw8vv1YXEnhTvhv/OE5tY/VhnO1Pv
XkROKYYOs3hTCz8hhwyyZVJVyysjTydt2Ngs4Ex8guFGZPom+Yjo+9TiZzBo
mvBbNWooDGLK6IzEgwvDx9TEdDuNiPL5ICRxHY7TrzQ39NGu8yrGgSo8P/zV
sqE4JjLBNT7IJrcEM1rVlsi5Np4iKgux7nnRTxCpcyyL+dWi253PxvjC24GY
Hl9bbO0sf+1w4VrdNnMTRF2qKjvYhXzYy5MX+oTj46GlERwGpPtZvnF8NMAg
fXFGRScMwPMAO9awgd7eV/v8xgC+txjFmBpTBUZMiwN32GEz9r4IMxNzynKR
oJyepNqlBJbkR/2OUJu0j2byRSRVGXzKGyrTOerj0vI3tREBNGG2col8M9kd
QUfCBUlOfsMbsOprpo8+LL4eR4WRxHoX9u/HjpCwn9Fo3C20drcsTNWHC3DM
ruW2mqogmQbXdNbUb4p9ZylYO7pHRpjuh3zxGhHslwga7fZ9mkdZmxfPeCcf
LfYpxvE5ekbtLuqNfcn+xdrsYT1QfyshZKpfpw7+TDxILDgsVTaP6vdZc6ek
EJfL/nUXCOHU5IlPK7coK7NpkdPBDDPVSP6qpCO2HuINOUCyo1ZKIRj5VBZB
ZNRUKk/5CTcIi6GathNGVJssnYT2FqN+hfZJjpmvMqanwmMe1Lx+W/KVfcL2
aZtfDadSzy2i5ENASzzIm/11JcpVFgs8Si8C4wS0ZDUcAXLnSPofABM9oujB
AjRb0lKnH4g1bMI+itYp/N8BDo3RIRh8b7k7vZgn5LcFZxbJuKwKfPEFJktV
6GgCFVri0/8AOEKr8DtEiI8Tm/0BdjNSHIeSnc5pFpYJhsDf1Q4PqX1d/Z/t
QxtYAe7PeYW/amfFgeIOq8qZ/10YpjV7NbuNLPJ8z8hSH4cEqZqXgz/0+0uK
48GW8n3Kk5G75gEfQ36h7kTFNxu/yF4M6MUhQOaABIIyWn1YNPmLx3I9Zgdb
dMW1tQjuOTbL9Rp1xdUSh23hz2lw/ckwMdyuwK3Q3s4qp5Z3bzkK2vtZfzAs
wot37OoDT+87jde4jW1DwRTA1tP3anXy/UWNrFFNSrC5xNV5WIclfgvOfmgZ
5ab4U3FcCWj6SyNdsrHy7DfZZvQ4BkVis+td/Rikh5Dwy+eBYDEp323F2kb9
yvFwH8Y4c2UVyE4r4xuAUbIeXEBV58vO5c0tmqJT/zpuFZ1PCNyBjiTG1TQA
RFZY7cYgERVzzNOzvTAGMafuJtPF9v0q1cJR8fZETEOiBfG2xjEsvt7eDZ7g
CaiUuxPTW8QNlD1B7C/9Z4YCZ3aLV/Au+7+DmRZ26JU6AdvKKiHK+We93xpv
H1+LCEmgkgnKSi+VPnblWBDmdiwyK4uXn85oByl0tMbzGdCpUHI3rtDCl9Wo
Kl7C+QW5T57MJyoIrL1fxDqOcdLClBcvZNHFtkBE2LKE61O5TN6hN7Xwo6uf
h0vjjEkJzyzVmA1yk1UJQS4SPXUKzpmCEKkYACljrtAaUXbUBHs7H93Igt67
/BmM8qqfJXklQShbkyb4KJI8DZ4t0Nm7F0VkZMH/xqvv7ncstky3zc3evitc
wtkTm2fqY1rQpghFBIXYyxK1KqguNdQKUL2pVoIoDgqzh+GUH8CWnxgRupAI
RT+h1c2vqSQYvX51PN85FCrlDHqEbaHTZHAKOSsPf/Ddm257tGQ2yhQ7V/Zn
pd9ifDvuVab0sR6HQPSuvK6o20CdMkB27nDtvVXQ3Tx8DYOHnEGiSXVZE3Tr
pckBqZL1az2K5QpTXD87og2hbeKxf26s7E7gaf+RnBj3zshbOinmHlugUvvL
yXCg7QKF+Ju8FI/6vVlFEK1plIFj0tcACAOiLvH1JrqscUMAZ4m4mTiN/vrn
+UGnDX8ySUrcDb5+UFS24REuY3eA9xuqmcOqiJPLDn461+4j+g8uW2DK4iuF
eE7U7W6DGktaKon2MTWmRI1aT/3agQ6izDyRQmezNC27jxWt/Pef7tuhubN+
grfC1XFyrQb02TOH0c0G6aYllJMm7D2u0IxkhkfocMrFY4sFG7dr65BAx+FG
LHkTnH88IMyPWfYItrP3cKnJ7779rSb7od3K9ofB3001aon+QFZETuBe16+O
S7xg1CPlxeC9NbAYZpFYOc6+SckuwL/BNrfjaQs/H6gyrycfvwGsMDpNGEZs
xLe1hlSP1LGr1AKnYgjEcMw1gZd/rlkkABI6P63t6B1jad0rhVzT3d5i1AvY
TdE7OJppLaPJUvZw0N86FP0e97QujmttzrrMXVaYIKs8r+L8Tl9kHVNmqqnW
929yCZJ8UZb9esyrTYICRBXkF0a2HtqeO4EtL+mnKGDVzrZ4ckL0hU1NUWkA
4SiNW2iGEl1YOwq/DH3aLejU1Gc3Ud/14zJcVithLRhmGOc8n8kV9GPopQMn
wPM/Qelyos0YojX8rFECUdUBlkxyk64TwXjJZlEj3Gq39lKGLfe1xHSeOq+E
PesD+RthIvB3cuymXTZK2fbB9i3P6Y/R1mULPb0uuxd7VX+CyVIDGpfNW7ld
1NQOMse8uKhCXRo/dehaHlFai46P3G4v9IotnGybOHXbb5BjTji1FwqAaUDn
TRFXHlJv3dTD5BhUW1+HICPmfWfleJvtzSv/UNpikx9sVDHFJZyoF504B/Wr
3T8fsY7wAmq50GtlSSceL3Kb04n6lqo/v8/mqCkOn2EelaXN42/RKEjoAR8Y
+cLVmi6gJIFkYW7ahems1QbYa+QM2qKORQ9m4E5U6/dAnMjN+koXQq0f+I6t
yRkzgwtLDj2euOFaG0OYVSMbNi+rrgan5agkE0Jn1CflAOySMbeI4YEe/Akw
n/U4nt/eLxtzAOJ3EXv2VMTlahd5CO6ykMsrvOwh4S2vP8gpkfcp/VgPoUCY
iod1sOXRtw/nqiW2vJtikvmqhMegWOEtF+E+3VWxBwMsO0PYbIeyq3mPUZBA
2OTk7C+Q/dQvcGOinvk8KPb1ww4cahrKjD5eFaHMfFhzrsuJ7vjb8+y9/fG4
Uz8i90THvLtHoLv994hsIO4Mq/k4lLXsQ+mki24Py7T39Oc13iNaCT2x5Vxf
qp9dRvFnBM89zu5yjk5wDJVuSXPsGUvO3s1lc4qGYwBuCAvonMYYhHbFcBnN
DGAEm8c8DeMjyq2qcVnlJuqu+dKfAzP6nxsFhpPhU3B43j2wqIeTVtTq3STk
8eAwBmuzcYkfBAMUne7q5ixISi4xeLcKs1/6sV7SBwCAQoddiKOBRmmoglUl
JabhrUHol5cW0Ss+BFxj4j++/lPEjlZVrQDxOERb/N14ZiX8VQrWP1nX5spq
q4Kl8EOdkawRGcpbPu8YeHqChuwUe9Iq5vvk//e4HQtxl9+aqfGA7Q7y1iwy
/PQ5Gcg2mHHrzMcozU1YMuLuHKfrm3wup87SEcPPmafRyu77wgPjQKkAxgKb
fpilvzP5mg/FIBqVPm6GgTtOnXEMLp9AG4wxoB7bkMk73JQUfZ4Y2LcDn+v4
KysU8xoNg+uA6EcMbmk9eV9p+lAjODBI2RrOSz/80ND9lAX4eR9WHcxYrki5
WQmYa7QN7FsXwCUPiPY+IGRWGlAD1SrK1dMe9OEM0rnFbSYZQDS8/i34WuUA
YTkdxsqbbD7jtkAQ1hbyll+iawGi8Qs7E1WBLoR8mjgPJFRRPAo2IHLQZejh
N+riENFNqSa0HP8LJTwgZdlB7AQOjYCITGKGL0jE2ejE4xZskV0buUPBH2xa
NL1krriOtbMPprLd9gaPrpovHO/8XkxPZAWsP0zZIjzWnSIanHa7G7lM754o
TNAmjmsu/ZHXzDpnbBZeN7O0Q7F6WF3iMWR4Cn+UqZxtRz0m+u5by7qXYfNJ
OyE2xfoQj4sYs9qtDT47jW+Gz/SQnH3RjbY7IcByvBJOQll5An4XQ2brkPOp
WaJAjMO1jqMsg2oWSlUTcADbEgfnyh1JywAaXgR7OhcKWTg3uDcYfWGD+InI
+HmI2qR8yB1mQbmpoehXBbNtlPSEZGsL9iRate1gRgBbT0ZTSF8s5xQf88hQ
jBaShkPxJlDtoyyRgx1+qBDsJ210UqZ6nIAOzzP4zxjkhvrFfTLaKGU2QsTb
qm02Ou2jsDy7gDU94E7j5oBmmXS/c10LxE0fBOG5jSOGyx+hjrHBwbXngTR+
FIBlYvb9dC1jbxSDSoyYrrjMEB+wfG6bWLOq5zhefRozDOAFBBZKGgnwd+Xt
/3Kfy2wrG7V7m9Hu6d1jjzXzwOT2C9UiH+V1f7EY3/66cFI6YCvNvj/mKURz
ZB5jQIhsPKsR1Kzex8+nhbh9DrsmZbF91QpOamCh6cOuEETGG5DI/f70RtGC
WSB1qDZ5EWYyziyC9zvmf3bPgQ76wvDUvY64+KFXn8/yCKj/TghET2T3NL7p
k/TO/Qasy9buDziwxNoFOKtJLYSSwKww6cpgBvtw7yEeDWEJQvzIPe6r8IEU
fMmVmb0BH/CySeJo7qPIP5IfHGl0ASIzqRmqEinWP0uvy0h2gIewWtc5SpCq
3/q39GYsMb/LfzR6VLCkP27VhnyQamfbOV5p65CkXYPyG/Nlh24mgLmOJ7gu
/UJf4KI/67PlGOYp8q0pHiB2seuDrN5lrMegcmQRKzXIpGGYJPBjj3z65C/H
wtp23yrkLKuubLeCulqM3RYdZzZgCJENz44lfZbbR5g72sBX3xwFpf3Uug1e
Mq1OFvkpqi4a/7BqKeSIEnKK3/HQgDcGtuOtb8AXuOYC49se1IXlzpraTPX0
GYBxc/fMmgOS1LdSdLuji/t1jVEdVGKI/QuYXckFxjc8PsB1709A6/ie3nDs
3ZNULy7Xf5J0oMxraolTdXxYX+gM153xFTuyjXIwmANpminEYl7NqQT1WlRD
vNaOmcHPvJY9DbWAMxPLTsBRBDxOral7L57AUFfxBfMSMlWntBOCCjjzsciJ
c8+lxyguWTle95PEWjZ7TacBivum2Ema5w4GiUrdxCqkl9LteuP/qUut+zaT
NXMk2e8YqczffKFVkY596ZIHDDiXtfWCT9IBEdYAjieshWh80lYazGcTZfj2
pXJCUg8Dz4+i+Pe7/v5wNvNYj9QzsNhBr7/5ww4e5v0QF4Dqtx47aAWrdLah
PGNlM8dxtXCQ3Bdb9ijH0KD477mjHPsvWzyM2jvSEvavrrVgiI5dfqI8If29
P98llOKq1p2seXC6NJHLN5dTzQbXUNTgaqkhNyGb0o1kBw/Ha2DW69Bk4Iv3
kRcLQPnI2hVHL5+m+kHC1XtXQ4Ucp8NiOmF/dotlRpCfCU9yAR/hHUXExotX
OAjK+P+rwfwq/yGGqoHWzM0E10I6oEjTR6BCSBfE5yzrsixhzq6nds3/cY2r
Q/gUv6BaOtqB7xqTUr/hNkCBGMPCewA3WP+uhOTIXtzBye2cGL56WrdqAP83
VpWLPLOCBazqAt9uRltN2wZxnQWsxAKdRF+O97/lZYchUewLvdJNZ5h2RHS6
Ln5ubX2fej7QRTD++PfhrBnEtdowWF+fvvijbOkhBQnd/kf2ooVQPvO1Dqxt
eDqfCVSUL7q2/D5S3YrhOG7Q1xhYp2/wiACYE3qZ4bd/V+/zjpqZvz9Tbl+9
+uhnbZWcsqCENdibaW0Sha2W46di/PUNZcDGuNG0yA5Ix01fqkd7XgYVqXGC
1HU8zj5sKUyp3nQDmJqO7IZ54gtQuDHFI4tCgCnLb6lUbjJrAkq2dreqmI8D
U6k6qS9s6l+EzNvsQ8rjElcgab+9yoH2i1oQEHBEDurm0P1KXFpYfIYI8h2G
7kgfw2RYtDsEDbyaYDrkRAdFth73ahJwH0jwZMKLJ1dOZTg773nRprs1H86j
cd42aMgsHGg4caCgEqZpoe8g+o/8KYWJ9aV9TKYUN2dKGmAG6D/eI3ibNi50
V2WmFftSUuwHkfdtlZsu5SmvSuZbW92z8Yoz+C2K89/6a3VYd3aH1/HlXPlw
/CJ6l/umTaPtb7kP0DoLTlT5Znb+76/3dME5sdxcc1fzVj+6rbwucNv0qdrD
y+f6AXv8jdnQJgrtZgNmQBSNIPpFBDMViVAvW08lKyuzme4WgjWhv4Qc+ByZ
9k2kIFHxFK5KgiuaWDlBD9orYJBMR9t9OGi78SJfAexhvOWPE+5hln09zKHw
O3vqyjFx2hlW6LDcO1LHOu2KzNj8/qUN49H+UALzquCseYGDgnhQOOyIxKAD
QSw5Anw6MRFEKHgOYNwFFOqmfPGLXZQjR8hNf7AJCww03/GjTYOIPI+WN08D
TFKWhv5ecEYptj5n8Q1uLedA0fpmEgNqTiEuD9kTlExTH1m4ITLSuTKt/EON
IoWJYlppgmLUtBU7zdK4hV5Na7ZN1Z6RPDtfV7adgN8KCLFWaJPoI6p9wj0m
RrYKw3DaBJnSoWSu11yWD4AYayE4HBE+RZd0uAVXOWk5fkzNtvV4k4RDqCsu
1boaEMe0guHszX1o4LyNYKkw+rzNGsa7cGFW3J0ujw2H2bXW8YPuM9vuPefJ
3T0ti+Z8/nxcKo7oOsE84QJ6NgasMfucwBafrw+mzY/35I8LHQvUCWggD8+I
AfCywUdvGsV9w+yoa837UT8YJBfz3MpJmcn2Z0b7S4cyf313sPSqPEQlDPK+
4ZWmzcLnvyMdmiZOj9yE1Z7t4S3vTG4S2qPdLZ3BK3edMr8z6ZJjRlcIWUBE
7d1LninzotDrhUyX6t4HOPo3O7xTJZEjyr4avt87kly8CQKa8TZ66k2RSUo6
L8R48kZfAHbaaQqFZAaso4hpQy5/MqtyN8p9143XfwXi1vnDyo/NPE/ZyP1b
Dzc62GelmDvzqJjbYTpaIKwDNalGzFUq49VdvHe3FkuSVUHntS62xRVznj/m
NTXdmN0xE/lRU2PqD0Y+ibT+Zd/t5a7nQP91PQj5EXIJXPR7KZGh8BYKK+TW
MrZV2M7OSjsV7aJYnX2OlmMCupLsQzMPJ9BRS/0nkvSazGy+2T8ciSp673hk
T398MexYQL+EEzKy+fRdrUrs2+mE76DeckEBieuV8doOfFelvgEB9uCFRpy3
A0/FPziAxWppIwP4Y8wZGqFVRbGeXV28uuGBXKJ46ytPxRe7YgyVPz6RsD04
hpHRjvamJ4E1ueOz7pGTgge9iHsCJoNPCgp0yLl4AwTgF8DaMFUoelFhSUso
pLC1lFLSOBdQFxFnKHDvRg17Fa+YZkE4D9BWDbJFDrMD2KkMR9U49hJeoTl3
BFFmUTJ+dMt8h7LHhkBwMyJ9VT5y7Xc8oCOe4Onjxzn0nbriRpPg7A6j35oP
r62myB0XPACuwFclkuEwmpGNHLURNMyrG6vOQVWhB+zagoDoBuDYO2ISZYNm
aSIHCTosGaG9qndGSX8NqfTTATHIhFuqBZjdJN5PKV3cpqLrraT4Jmd4qGQY
I8xgxU48+Dhb3GwvP2c0FLtU/geYFw2f9B3Wvisklx2PZQ1faLLoHCm6GZ4R
xhMr14MW50w1adKSkRaLbrXVh8gBGucZyedvQsWEq+LU+ParJSbUeI558LdN
oh5/6lja4ALFVo9lbI3qCSPZNvtCLQXMl3g0WSq4fPLAsBPmGTQPL4lgMBzm
7XjLAoQH5CdAQmkeYRtRBVm6mIvF1LCZ2LDsHXLoOxgLbJAlz+A3LwdA5XED
npAqZ3Vs9OBPZ4ca/d8wD7IHqQTTu7vGRxF4mjexwb1+nE21sdvwjAYRbxrR
7jv55Rpq3BD5Jm224Sd87y95BRZy2XA8RJhBbGUcDSEPIPHI95bjphZvIWV3
4J+X2BcFA9PKH2alaa3Di/KVK2/77DJU7jIHjEzN+d38y5YTNhJ05+ZU7c2s
vmYuymVkxNHxYaB2Gfp6eNx3TH70kmOuXTs5wwrq+F4A1sovg5HB/OTgD5At
bquaaiYhEzPISFF+hBvfUqj62wLgKW4Y1yQmLqJGVDUnKpU+TL6gVgkN/rXC
KwUSYuZxuk3Z78h5vblbRv/6TJ2L05AJ8WCdHslxEgGl6teTTdb3lNoXheRW
Rqq2Wc4rf7gFtKMIX0FDpxUVqcBipm0vE4T/tvRJKEbvFgWz57RnW09DxPzX
XA2gL2JjAsUNRLsMGog2lA5/qeXJSMUY5J9qGbA5tHfiK6Y/8Otrmhg7L2Cn
z3XgJvPnBrJM9F9muXC+T2fHn1EqMJo1sgK0eKt8JGLUcJ3Esu87N0YioPmh
f9v8id5eDTUrnt6hNs+Zu5BBH99v0XPVh0FhAo7yTvj4N4o+RmHL5+CjTEct
hGVB0LzdwupxKyM/gGT40jPfSShF06VRLSlmTld2h0SIlXoLwYDABpVzJLBB
0BNgBUAc02UFulPUG4vR/l2QQ/3UADrC0TfpfuGOWMbBqKTWhWPizC+8uA1x
l06EuLoQJXGLzDnqO1kqr5cJ2boOvPQEGB/5iRGKS6xZND/DGJFykxoFvOlq
e8FnPWgfQBemGYOUqImeqgczrr26vgne481PzJbC2Ikncks723wWRjExHfTy
slMVeMFOmhk9HN3h8+8IJfRWZeyBxuDDNvntNvbUswcrQAhoUEi3RmkaKWSt
+hHSwlm1KqzyZ0VZCIYb4dCRh1vNyo+ihXG3JLJIHPJRO7hJcmh5tfzqbQSH
td38ZChmBxMTr7fbdgS+q1iQjyERZcoz9nz3qSthfKYKx/K6Tll+tKk7OduI
B4zHMJvpPhIOaW1BQM0nR10r+4ERF9EewrDwJ5lFRLMpdovRk60qRy1Vyxub
dwE0xfu/wmJxLqYXKT3Vm63vzuCQKaAMtNNiHhnaf5vh37UuIm4krMkic4rf
zlVAduMaXY91D0EkxliizY8X9+QGStJOJjW2x/J7DW0l8WZYLJN9GJ5PR105
tDkSMfZwl5W0yIb3xp1t+yVZhqbPqaqMxefC88ChoNkM44JxHFhPDVmr3TJz
x+ZhLfga74hB+TArGWHTvrepe6axULGJw1Rz7nZJ2T/GGROxbynFKD47YE67
bS1MiTyiSefm3yCAB6M8kSzretOOQeqSXC6uxxovp780gWkuE2FX2tkI2knx
RWv8zRnUsZuFy9zNESuz/gf/5vS8ax5LmVkAv8VtTOgah3ISVi5Ee07oD/Wi
EYCQLIXQ7FXpVsR5XXY09OkY81g8P4zsBYJ+ej1Uw1sFPbuaibsBg2Ea8jDY
YloaSLGVvSIokZNr7xIeYuwDYaXMZfCqvCKwM46XSdVUN9mt9QyxU6QiUJpz
e2yGaTmyMwjh8jFShdxdHEfZUsohEs0yjIEqNNkjUQSeCH2Pp/EDaKYMozmM
YLj4rEeNTs/zQnK8U9Wrd3TH4+dcAOAzRJ0kg3L6vTuv+qVInDkeNsN3nwrd
BtMT9pjx3OuZ+tYiWPVnDAmJ6Y+ISwHZv3N1yPEDoyNGJzNMImSzcUO9JWfZ
eTTUk3jLAe2Dwsgb/Bc2gKw32yCKkZe1vGOLEIIsisEjJg0QoOPQebna/oWI
QKukRhiNguetpEa2pIPb2Ewkyu6xzaq95o6oYSBgCc+2FtHGhmeXcjO/Gukn
0pPGDmimiBphQNHuR3RuFA5PxVb51/PANkaoOkveFZm+KpNwjWh4y+sLOBLT
35mNcOVh9ogcKO2NbNPLtejXlmxDrROp6ld0G5zu9YBajo95QdYDmJQm0oVx
kkw3mdkq4S36o94nox/w43WKsTHdCK8f8hbW7iDPLhevpaVIV6MuRebDF3Nk
vgDiwmbRcqYTqnBqgQmhDXveEgNNQTSzZQ/IHxJxR+Tk4pgLsZSM7K7vgsWC
rrX5TztIa7tnt7iIMTIGZGIrrNUUkuBJ2iuECe/XtdfeRzKQ3gQrwu+axh5T
asKEUneETj0j2WE3hLw0a/VeUD0cWF4/hAtUPM75+0Uh6NE0dk+17i1mZ9cI
frZT0cMcbQWR/zB2Nl9Rld2Kxkym+VBfubYfoCHfDLBkFXc1gKyTDVMcqcAr
zzR9Y0ylNpP1CdsReV1NN6JbLD2iSq97S8KenUi7AgyuybytbEeWyrxV6KzJ
VVWIcwS4Vnx208skYdgs+1++VoaJOlfe2EWn9n+IrO9Fsw/N9FAxUMSjEy7o
2z3wCKzIKfV5o/SyD91AUKct+QjfMFEJ3+hsJLVi1yqgOUyWyhp5JzTNUw7k
OAnOFV6LLNj4oCYaf2b6Ierjt7GYkWtZ6bOL0SR2hqC/6Qb6/1i2XkWcZTcH
YRIFraUzHJze2HpM7eBPasDzw6mub/DJy8DJkenv8KyLXoZw/dDGfyNzQEu4
O1IfVUfItRBlaPw4/qgkP4sF1NYyxFy1r6e7gjORSOE3aA7b8a/Ps3Ni/xiY
LfKeK+VJdKD9vOs6mfpqH6qDELGuMdUSD8FmzsBPDPDH+nFAiJ8744olBkb6
+t67pJHl6mLyZK+8sGI/bHxDajCcfOUPA32FUbdFkNwUfPXAP40sv2o3zz/1
3fV7ivMk9FSJEa0F7s5JYoVHQF/7g8dLv5lxG2Hl4nsF9RBW0z/VmL/ZWsDz
BT1yOXysHXZh62rMTiO4WD9OPcXK24NJXU/dHTajcWX7vfKnHivolhvKd/0f
Otxj64M8Ti74Ha4EMcrCYYXC1OLGv3RD5uirPa2yYQq9V1PByp9kjaxt/VfX
iM1KgCo34C//OmiPg30E1lKFe7ah/0zGAFKx8sEa4Q39oOMnha84ih/MGNF8
Uje1BIUZMxq8X34yYAGbLEzZd45+uOMUOKj7Z1tmaJ/5h8EZpGJ6HdLp2RQ0
dn5BfJ3QPXD6YoUPRUlgnNHX+NEF+t8U6i2iQTM9n7dS2TKkgp+rv50cav62
Z44QpUczQebHew9/Xwc95y7FwYo9b27+2WvygKv73bzIdDrISVnbGhf1jxhC
Nzh0awYwH0HughM9zqmJq4S5DU7JIHg/sbPqBFZgbS66RWHrf0nNo9SkvGDe
gxxkK+UwzPoOQ0Uecmj9DPv+Qij8cD1vNNDT+dM3wLbB9dXeQzGQUN7OO6mr
AIZ/EdySJ8W2WpjbXv4nnahIv+jzQo13sPweLCSY/orrqfwW0mnNMh3cCUat
+qC76drfM7+T0MCulL0d22IPKPAazFN71I2AeJ3JQ6l4Q8fGblerR/s+agd9
auavq4TFRDizK60yXDZWcbs3tsa9TTzqB8gllDa4zmfpK/GLw7EjoE58DFo0
QDwuawHlYMXoXOIuOH/K6ZmDQrPrRGf0mTIIR4aXvL1lwjXZk/Qhy0kQQHkW
ENB/jBpOPKtH5w891mPEkFMUzoK7yjaQGjhX3bWuBrLMmPNh0siF4DiFvv5S
hlhJn7iOuPFolb+rI/EaacKYmXR29WvSmnihUAAU560wQhmoHVzpyUksDy1f
aOYjBRsJT+sMMkuwYaQ8TOVq9pUZvIAe0L44slJaCEXFc6UmqRXEgVvTUCc2
WQEE6E9eVJOvOvp7HqOTT/B6Zd/tR/odHkb4CKtmiX55E/ZdxnAEmW+dLMMc
OQWWvoUrn9rlheLBAof+babe8AexZqdMPA4CNl5uKytUY+X2BgTi/6sguR/2
JWSycLFKhxk6/ml0wpnbw+LOc/Lfzw5m9o05q94EUggp1zRMbnVGKsXt4wcL
91GWBchMUIoWt2yQL4j0JJkzgoM2rDtiUBgGS0+Q+/ZyVw3ASGb/IUCtYlZu
MaYYkVhKZR4oGi3pxtXfb/7rWG6FAtvWcFAKOSZvQ5P4r0YWLBwP0tfBeMlK
chkieL4vUFsMGlLOGGGgF4ZGHzwqzruYtoDnBsLAw3YohbrLExMXR3vVDfib
6ECbQD4Im5jlXvVXTDePUmQqDCn46+Td/uIfLxYCU/xkMEis1CchPmpK2O4w
0Ph9GpoNS6Bhy/S/sJB4XJTMEcENCjTRv/df/HIgY5l+O8sIWsZz9oEuFYCc
yIk3ejp0wgoF2wH1ylXB0GL/CQL1i0sZlzjgibDyrsNRPod3aQ/Og9YuvvzA
l/ZZ3OlW06a0BZagd1P9DapggFEeRnu2wRJ6ECKDF/2GJoVYgtKg7Z230htH
nXubcg/Yo+Pux4UZ+ESCXorIfKrEm3M9//T37gGOrR3o00gpT0INEPRTPG+r
v9MCF/TijPHZ0M5APEpPFTUVmnqoBNaTh83BQug5cBaIRlTESZBlaWv/sw3T
FtCFJDQTNABjp7m+gmpHYLi+6F4RHeRar8x6q9YfxooFVCPKNi+5wYAW1s+c
Q0eJsmyTv5FGkhKHHIiM+wWKBkt+pU9zusytwYv5twPcppbBrGCfUjRTvi4k
9+k5IT3V5N8hvegeHQDgY+j8XfNIp3X8yZyd1IvBqHQ1Omy0woWCAp2MtCt4
VbqcIAZDXhaxTF2tvY1WTwyyjRpoNqMiF8wyInFSlVHqvUAd4kz0/XWL6rdm
T398GzJHoreJvjtW4O3ftC0TA4OKetXsx7ZejmIL7v+s0koKkJsxeqGyAryN
02mhXYcOf4VSgaZhBT43KzzLnTd8N79iDW1PJI/GxyIS4c/s3r7upeWd+hr3
VUYVzN3Bz09LDGpXqtcnUIdaED/4t0wjWmaFjfllKlpHXFY9KnNawTtFQGNo
qFbf1cxtQHVYhgcEOysLdTOWyhm0ON8BbzXLo7z6UMDzCSUZdxpQF/fmr9Ux
aWsVqXs91B9039vS1uNphHwPjOKk8mBGMvZoe9KW0HOBW6wWuIzNUG/dIHZf
i757codfUp/Er97qtpOynpCJBXQjMKHIR7NoAT/utfg8KL7Z8U/3M9KZMFFI
USYsRj6Khke7zDs93rt9o62N92rlgjve7t2suIqjhIAHFIDgeqfTXIVjIBFO
4QktpNYE6Ll/RmXz5Mx9bFsddQ1p/zD0c0kWhC+LukZkdNRyupjKT03aHCYf
eTI1FXHcF495aNz6Qxh/c+Cok/4eSHsdTbgtypmKCqeLEaTw7LVSPV8fJVIX
d5vJmqGsXWEHfYdFTcw794cJxHPJLGFAKm56VY3kjZr+ZfptlrCsX+PHVwyq
hYUD6dV9veQ4SQCu97xNoJ/cIGsZt+/SEtLU7goBQE/iwE7eVfr73Pv7r1Fd
+TzTdqmztTf/S7bpKiX2gx6LF+9Ktr8Npc5B07SlekXb0Lx6PR/I/AjQiOA/
IvE8o78Km89jk6xjVkoWMA96yBxXgL9bTjEMOUsXV5FhsYaDCdqamLBMiGgX
XGIHGC6QSD6Ga1IU0f6/DDPPpi77OCb3GD5rJMimkl7RzCc8uKISxzV0BM4H
2UV6HFmeOQ+vIJNM1A4n1FmdjUowYafU0LQCo4h7ARTd5xaHOibz5mNPCWF7
GuBheBi8dW3v9FHWFhGzXAnq7RR6HWSRkbPZ2sAEVtxK3QEr6Z3wSUU/IHOv
jLcPqGEUHR8IlrD+IYFmdkIPeJ48YK5FcAneDj8ZDn8YK1SxpS/w4VYkXIGh
VMo7i0P4oJDzBBDNcb2r0G2JQprdFlZGHPzEFx+V6DLJ9lpu+7Pu6h0yec7s
P/Dko3aVYkCigCAPBfCx9+jSJVzQhKGr2ZTUK6UU8xuG/DamienrJv8T2JQt
6sfJBOiuhXkpEz4M1fuZEEHcgJ0JJ5Il6FUtRKalHpDGOUMpQxONUZ4yBU5l
lx1KoSDIqVdrF9r+o3Exr4W38CZC/HUp44t9ZTlnq38aVUpM0gL/6M7Yzwa8
OzlgY7bayekGHYiEkhGui9D824OaAKOHAnBBfwP7aIteyWZ7fNpULhI+sIGc
kqcz78dPIiVEahR4zcuDi497bRC1kODexiXIw0fkUitlo9ae0GpbJJ9QhKvg
KjFCkxeLh7O3eJ4/8+WAN1lkZ7oCg1zKybRP89gE3Gmi7UBFTCTtk+IC2J5l
2mvNo93tnNTGoLYzsIJpwyI9ljOTi/mJdbPNWJBSb5lhTfYbpVD7G3EMGJWn
D+Hbs4OVzmVsy+CcLqX5788H+/iHajFwFC+haQXogwHwvlWgQYnNujDeqO6q
JVIHcjcMZYa7DoVqA/5ddqVhPKD51zScmRjXnvvCZqSq4q9fbUDRJrazoXq+
Y4Udx6eS4OYL/UjKjWc6AMD9AICtd1xBVwY64DYMRNXiMj7vMThK6xC4lFvG
bVZPPMF3qPr0icQwX2LjetM6AqGHXQW0sANtykcSth8dtbnBnuPHyLrFZqJN
U3JHzVY+VJrARG+bk7OcV+NA2w6Wus1znn0GfsCn7InWsCAEDIhhGOA+UWkd
1I1JfKb2rZiBpJK7u7K74gU8AYBCwiDVrwNZSTBawFJMQ3mZZiq+wVKjPu3v
C9CXRUS+TbY3X2q3iXqi0HokBCATT7pt+gkFVb7vdJ/o9sRkRw2ODmfnXPVV
H8Bz/Jrai6/5Me9+Za8jTwOVLbLyuAXB8j0WVnujcL3ovS/hgxpKH/WFDUZe
0ZLwPTH/qWaJ9ZIjwyziVH3yCqVXdBSCko2d6qDK6m3b0wBblTG0wHeegbsK
H0BJNFVZKigC7vRBJh+Fwut5gTb7Rl2wA7RkIBLScN0K6TzUESNEP0BNOZSE
JFs2Ku6WnkkFxVrocrYfVaUC83ziaEDg87oVrKEA+OgLI9g8tInQ7x1mlE6g
lVWQpnWXbyqPSNoJylEk+9OZVRXRLoZQAPiH17HrG+i4UvnhhUCD93MoQg9B
dvFMA8ZFX1z6s9K0akuotSgM5uzFDEX7MKGwHn1tIYoHNwTmDkol7pQIfQ5g
GLvRdA2YhQ2EjFsHdPIfAZK49SyZ9h6qYykDE3gPR+6RosmpJkxMSxsNsYVL
xSX6rlS9EYwj3gQu9tfGYokMms+jKX9AU6N1HrpCZV+az/+ytZWlV/K492Pv
gbpheXx4XmrpAQVwDfkDv5QkpIkrhxT+ZzPsfbZrFLX2S6qiqgpSOaN8xEPv
W+q7lHxNNVjjAGBCPSCTrODF8vonKLXxPW5vIwrzjG74qKI0F7+ote99bUPv
yIrSkuGhN3KEEEVQHjZaejP68NkXAhzZtjgeuVPe50UBVzFrLmSbZ1jNG8KB
KJiZNRvcseaTkWkpuRcy7e4Bs9bnF1xLFHjNZBMo/44WKcNB43m8XpO1c+3e
0vpOtHlNLy/meHy2wytjgQhHBzM/mfSlmSdedekbLnBhEzxSC+fxAf+/K+Y5
z5QfOKXcZc6f5jQUx9cl3VLeD/Cu/ZuDiGUmOasgJFOuJFcyAF1g+4kkWXLH
b8Og1ROGOZjwBaPqsz4T+9xmuDIkoq7N1F94SPoKKXOMWFaP1AY1vMK+rf9R
D9S0y2ZSoKBtF5WeUF7NyiLEQrpc+qqE4SuXtvLjJrkqyqZCU1ava8sISI3q
bl+ciI4wyuOkRKm3c5bWKKS1gJy/XJ7Xw10vGzCa+8OMFZhOXSLUwhjTq0sz
IKtX8L/P234BqEOpAMm5+HjjdVydxBx/8O3RstsxU3J8AA0931dU7DVp3T8b
itlUK9ETQW4ricBmdkIdIJB1sURG3N2tUz3Q/ov41pFscwn17dBjoXdMHzLn
EIkoR19u+5qR3BpLeSZSQfEF1kDPLJoTwvqrK3HAetrcogWSDZSj8+u02V4P
bOjMEXVahcfJdI7oygveZ9xHWqEITN7CGF9QHtK9MDsAaosUjz3dv+nxSPgV
GvRMigrCNEaOtiEQMzdMfSDX4J8N/d/RuubuPl1J+D4oxgqtk8oySct0Oy12
RFpS0YVjM+ucQ4Wu1pXnyjnXmltIXpHT9aGfxOVxAj7TDZyskoKYaqVPgO4o
Ak6dPfUDyuiYER2Ot0/Up8kvUgFb5b/vP/znZETO2m08nFXTuhvAM+cF6HUf
CGX70gGYfo315g0UavJ5wqi9GW7mqY9BuHs18a0Rg9WjGn/HVfd6PSx+oc/c
ZPbXo+B7NtijZ0EYBL8SE9pWzqEDB8BFwJ1UhbqA8n1O7rG0837PCD85w+Us
glyA2sfUFcBC4AOTRr9CYQBaTBRHTGDsTODFWDmzJrFZ9T1efg9bb5cM20vw
lqlN/Vh4S24ATDwfOVSyq7jkYpQqA8RC14IkhgGd+r5jE/45FKKDoTRyyuc0
/QKbVLofUHHPX5AF9ncDnYXBheC8Dt9VBYIaWqGGEBfay0IYfQp8UpbJ8zJ+
fal2Ol5Ft2BaxgFAtzI1Dc3LSB1GKJNlRoD2dq2nfwVVwXGOwL9dyjYMRd3z
y8KN98aTslfHJDv92PxIrWJWKu3lEeN2bQgH1e7jj2hm0ETDy/Rk5lscotTy
VNp3KU6G+X20zkO5x3CnsuoRC3nHoL3SOEVX8gXbDG4cFaeyJQNsAQusDzQN
GHOTkcNmuzDERAq3eC0+TKdNjRVlU5W6TV6chfirBTj7/5PFoQsSUAuNjaHl
FmpDtKdoNG2ZZD3onXMFyIR4tXbPXGjrXGZdRLNW+xjxF7GkS7P2HGOETsPn
LCgd40+YgJEBOaM6VzayD+iq6TO+5SoQ4BSRCyiP5LnaifuHG6QUCjAu3Z53
DR9BHVqE7/zIvCyuX1xkf1t4jSW53x6aVsKyowQRvizNiqs/dME14wEY1ycN
BJ9honUg5Cl9SZdKSCAAu2hkJVNJ/NPeRkedBsTuSjNfgDHDlzuZ53KyCvV8
zSj6SE6g5Ak4S8SULzjpDU0gSJVOlZ+bbUf4qw3rmmdVYDbCqtduiAafacd5
KPBkln/fbuUzWgtQGwiyCQiUh5S6Qcs/Bd99fGH8CEWTRQu9kG3PLqrk72do
27xgBxjB+WhKSseOniI9bKKwyZrDsz5lk7U4tALJIq6A6ep3rDeIYmRV9Hwr
wNNGBCcPcusUqvHEi+wvcWcDw9ALbexdNQ/Gp5JKmKfcsjjfDZrL4AgZcY8a
a7UlS9ggGTCca6cBZV2i9X21P+bdHrCO63xw61lToxa7Uc1teWw7jCbAKIFd
jNM8qTzF6DCdaB82XIiYK/tflhUpK21J2VQhUFi4Z5VaVEYPg8OhrkaN7ctF
rErme3v/Daaftx0hU5rID2gAP44D3aRLWHFuS35K3gQKCthpDQIG4cg3goEA
pcGN2ubgYUuvsAJf5ifXRqtprThBH8CmSHfMopzjC9ckD9Z7Cv/qM13S0Vu8
/lbmyDyNWVBzKwXSGeLnKPuF7cYnnXSRGCwSfyPEdniCFGryDyPoP+v6wzND
sHkNVkhqdRbc29bYSslg07jsDvi4Q4X583DKh0wNm6Kfh/SEAmIcYZOYsYQE
evfP4D2ipo8KNXK3zJcT9nmhIXcvdahLQmjjugoLq7KpugbHcUadSay72PwE
JwPkR2KRvfE1ZoV0qKLsbBrmXyDXvJjCaq5ZXAJJyq4nB94ecJoq43cryonL
BDl3TNrYn2BI6rvIMl4DBq7rAfk0Z0SVpO7VcJD/Flai0uErg7etnlGSeozD
Qv5Vqcp8miTqN4/Xp3UfedRExS85GYn4GvZAMvjEc6IDY6FKXdNQnO0MhMmJ
dVFwBL6FHc9yrXIcDb0PHoFSiaQ5M+IGsCnJpien+QvIygurMTzEjDuQuAkF
KejBZuDAWphIL+jroLid0aUlsaBbpIOBNLVGVg/940olc7Z9qdqGUQhpdtja
o6+bnvNhZPMqdSJKlFZruDWhVhUg2BIGaRAZ7F71LvGmMr3Ezbb7t1rJWDC8
55/LayZkkjsNW3HTmuWNX/REhB3Suj2fqz1kD33r12qpGvPluADbR8+ALEhy
wm6DvqStacq1Z6OsMp5U0WsQ7L1Ou/8lipYnV4P5WBiyDRgUN+UoVmaJ6smg
EIoOICmTEnHIrF/4yPtNvKeDIYPPJorgU3W9HexpoJc/i0YaBEutcywtC1h5
1thOStq5Sof+dSho9bCp3dogFStf2o0nStbsqqw6vrsZsqFU1rF+r8Mo8SiJ
VHV+gIlheruFrqBzBPgpKzuReUg5LO5scNKOx0PbBcA1cmUzzV9YyeyiFoB0
l2RqDC1OL0fSEZDPnhq7ZiXf3MU4EXu4rpgqiyETHClvB6gopbRPCMtLGRBR
2YNoOx0JhEK7XO9+umFrU/Q3v6r6lTGnyfLD7/S3kNpq59aV6+wAYENup5Az
d9w9YQ/wxxb2KsVQqSEsGgkC9V9yfTuoYnQdWh3ppcd6iyYAryqqEuLd5UAW
ADKd0GLLsbm3k/2xfYRDVOdoA6U5JaEuBcUGpLjJ3SF5QJuuu5kvKAMxYlJr
9smM6S61A45UpXZ7v2mqYbVuVxsZJyXQaTYsuRVOzKhrfp1rW+xo8Add86Q2
4obvsSahetKYGtV6zqXXYNuhqJZAGquisc5665h4BFbDsfx02uun2s9FGK7w
0NvXkSG2r7vWzM8vrV0UDYqHfQScY5RiQxM+TrrbXjdB7U4abKUbb3JjlO4F
dP+26PfRSG5Utg+Dir101FuwrT+k9g+rvgb3hlhiQvpQRlPFIJYT/qI3m2ho
z0CGEZ4ktqjfWs+P6q+SV6/vDKiydu3G4odUu6SdlZYV3tdWSmeux7ok4f5y
R+vE+a/NfFptv2qvHShWdvtsQLGysAYZzDDo3Q1hnVsgnaZ+M67S4zkw3gES
Za1X3UN54oGTDnNuNKz0qFrtaftIxUs+apDY6leF8rL7aUEg315E5/ifQOOY
kWF/rYafxoeTX+NYNX1FjAiNheyL2rIBGBFuSZcdXgLngfpECO4NQ1JZUhOD
iCdsd2QJ0+/E4BCogK3UbXV4qh/VLI7KRTcAdAe1IQvEqIjgU2X6UDwaaKCq
sjuCN4uwtkabk8YcGUTKgdRg++u1p2qLltbNiOU34Pfi/IGzqx+zfDYBnejt
nBP70Mtot0PL8ZomIX9dqlFBCvDkd/lv+VsoWZiovb8xSieco4jKZUKztWLC
+lcHrVu76eH/Ys0QxMbvIm3eEa08K16gGmsUoFJ+LTuDLSH1xy68XoTKOQvZ
QBBgJWtnoIvO3AtamVdeQ5lW6fCTmzqH+iol71G6L4NKOet/uB2dHWnfo7Ib
v8HuobFyTr3iCKpGyXgW9He4MwXZnBaLPZWWWvyrMgFRA6zO6hXOriGRtMKt
nDQOXDi97yLkHkzK/d8z2yMHBJbCdc8YL/42yNl8/XH4ixPJ0qSoClozld3s
G6SHZJ7lI0EoN4GbH8MtfIT99McKvL6cpTfzW1E1l11LlpfrMlBnZPX2KCM8
KpcCrOPijk88KNOsW4+vPVStFNgwTqS2FapqQDXY80AlZO4gAZoO6M4BhzgJ
nbmZGaDb5Lf4+ry+eWY2mBxl1V50y0eQfYAG8tlQ5Br9J7/e0kT85hkZ6SZl
XQwtTZDvSQEhLUgWx9kdesZ7nCyo5Sqm6w4cEgDEn26oP8fjQVbocYWuFvaZ
QRNR+80YMCl/msIUQD7ZNA4skAvo0/X2vk+KrXaySuxIfV8vjGlS15GSs7x7
KDIj0yHPhQq5J1BoJ+PrlS3/n2TDteLguJ4LJJMk0I5PT2w1CeL5qV1ai8pU
/WUt5k1IWWCZe1krCyz5s7f6MLHrBPf4kHk8mmUrP+vUpqUjsIlxhgclpLn1
JI5ED3HrgyGA7+G7wWdiJGx2Jx+qeg9E+4fWsCblEp2gXY7SFLx8ddwYVSOP
pPXK/CBZKpn7UG0vBx4a/7do4i+Hylt0H8h+Sm9k9Y7MQWO1yLYlFT78Rrdm
oo6SeOKJdgQwQtvNgnvrzxNaQ8ZwPsrHVJU3DDfOKgheX4pmpEc58D91yQ3M
HHS/yjMUBHBdPHWTR3i/tP2DXGKU3hXYih66itRhyoTTn7iURWmCoRJrxpCf
mkNROo26XyhV2cEVl578zV0Gi08UWf1521lwNrdveqbdJ+6JRuJz1UAThlVn
8tRwKDgEJjRD0VXVfuUHQRQS8oDKvzApv5szNSxED7zk6XlULNYtFiCMKYDM
6PxqRUPvwR1UHRJDuTV766Ghlo0daIPz/9NOrq2rJJWeyOkw8QJj/uOZQWFx
v0t7Bn37cFowACJ9ehUcgP3aiAptD887EfjYdFgP1Bsv0h+l+zI4IT84Mh0Y
lAaL35sRhcElxFX40Wk6Xn28+G85qNmcsu2WGDkgb96THQ2oQtKT1lw7k29n
ZxehCPJR+G9awLZyapHKneTTYyGDnIjcvblfmrv8HEW8StqDyRQtoyeLjJZS
v4xn9lcqlTO5O5m9rxsdlRBCeOYgirim2cAYs/fs5ecnbRTQ+jPZ3wPiK8LD
xr4+l4jCkd+/KXTrISSssv7yq0Z1mtNcE621PXn6JjHIJ7tByvfCkCVcNJSl
I+VNpjaTS4UHVePzE19P1pGYyuCU2vGvB0v8zHed5IlbZhZ3clapvxiz9c6o
zFebgmQu15O3PNNGfOx1oJ+ODfUqVx0KE+p3Z003q2RvGRvWt8hjGCMehROc
AwQ5psDO9168CYQi1Fr2pH8NuArCm/k/qj4zLd84vCiQt3gRoN1tWf057gjd
+xfZWQDfrAEf9reJSfHWo+G1VuXT8/QMoYETkQHUZqg9iTBedcvMcn1d5DVV
Ii3L4qCHNiZ1WsiTYF4sdRFv/ThGYFtvFCu8befSwIUX78+Bs15ILJ9Hy/wW
5dEYgIcnjfKBhXzSuTykBLa0JRnoFl76cpn7tr3/KkkTWFv1goBhDRWqRU5V
l3H9lAKNl6y2bbYWCimMYwhzaqwErbAHepTqOCOXaKdaVEnDPTvHlX/nAC2Q
SAkd5oRIo4Zr/qz/Yg0YTn4UlZRVp6rNh4ycgrIbcx8+qXsAGQrNr/vJ6u4z
G1mCPn0cYgnYRpAabk7d+VnUd43qDmtC3wMrWN923V170quDNWUXFYVSG3ZP
oSlFD31Q1outDKQ33nSJxC0RcNbost1pOlAb8ru+I/F4omLwbmTMhR3dUoA8
dhlIn94rhaqlPwbwTrk4BYhrmz+DRvvoAy1wmEYcsNKL2zMK6iE2jzBRi9FV
+l53HoCCZu2r3/ToRDMw2uIqJjrNhup2vwMyxRzX/VzkbI7T+k1WYWY0oK9K
SDXz6OG8OU0euO6yBE1TXpSRlGBe5ZQIPNUfsTNmfEW9mZrZcq24y44G8vUn
Jr0gaNHN4ATPR1WN+EsWhfo1YysoNfFsxlF1b5NMA6iymBD2vAia1BfPfNTH
Xsa28a5YzttJ7AyOy2RoLeiu4WHj4tH0V8noQPvwWO7gTkO7vV6Fl5hyJtjN
8wCYr1P4WfmHHgHeHE3iNdWGooDNICAK4nkFqg6Nj7TFI/Ho80uHkyAbJPGE
dYfyCwp6sPNtfa4wHrUFZn6eK93xBYSqDm4w+VyIt8HqffMEhpRSw+3H95iM
kychE7ZOYLqjZOSIOjv6Ud6h6GweJ7fptBSqUh6TLeSG+pTEd1Fog7fDaT71
LU+iKVdlhqVCrQahmrjaBvb7Hl1dY67bMoQAmNmlvFRmcEW2irc2BW3Q+DLj
JLjvTpoNGhIRbXU1g7GIBw7TlqT1O97NIkPgZAWF2YgBoRBesOHdTjQJ6hpc
aoyj8grg55x3j4eM4rfitKCCEcKMSqCRS6vBdbu9yC8zzUMbZ0wsaIPOeuPr
aXGmYwaAjsUWlGi5s+ErtDe/rfF0UyQCZb35qTCvQWfI2uJIMj51WnfCXkm4
5FDOwkYiHl3UdEdZGO27ZIKU6bCPYVzsSMkvcgM4PPBERK41zKDJBEHYupx0
bLM1H9I9ZuSaqSEAIXLBO+e3GNLG+dPoUoUtoZ+M/6+1z14ARUrmJuexrzHX
R0z0QmDmi+qctoHMPaDZnu2g0paWHDrBpmknhuCY6xsMzbcDu4AxbapuJH0c
0YahgqbTvxNVqnpaC10nArbwBAPM5n4NzTI0QZrFrrkZ4XMWvrck17a5gE8Q
CE/eLr1FCgIioR1r45iJCpvpMrQM4RxecUNbQYIq4IEixl7h03pmXHsNJm12
kS2ep5kMsukE8P72nd04zcOjUqyXyQuSJ1kCyJXP8agnQaAGJqWkoa39kg93
OfEPeabLWRVId/w1NqVPblxhE+ih9Tuv8nuHVuoP6vSjjhiDCfiE7OBZ05JN
8+Jd4MyKQ98j0xTv27oI9VICh/Xo1KlP7hKyMFbGucy+RZKQ6SnvwP7h+/In
A+sHhjl1eg0rPMUfkUq+FLf6NpCf79jX/y/0mIFWJpeGX+koefNBcPucMrAB
fyOyT29PixxMJWtoNC1sWfb2GadEDn70exPOHEzRo/5PAxNzS+0iMVaP+xIe
C12/f5G6GUNqAbRUz+jd56wk/Z4wNUtrdDrDNuar4mWmtuCY8o2k9mBX7fH0
sQQXssBQ4Ee+byp8DkmN97TWFndjrQavIesOKpOA4KKDwdXoqVZzWgaIM8BZ
VNUuYzyjFwppaPZ5tkKOqO47NXom1S4/DnBSZ9vqdWumul1TQayDQWJwDxa6
5cW7BQgXN6NSLmz+tFKnMfG4xONf1r96dnZ12thDpQXQjPRbzgVJD4dUrOgl
DPntkinUe5g6RGAeEJxElQ3r5F/0gUKlL7/8lDS+VNea+1eSdkRpOhDFuswz
1Q0OblbDWPUhGyc7HZUrfupLLmLMZikbVySdOyGnyW7ZIVE3OOEYEewUv0WT
v3t5DOeL9kh/iS5n00UY6AKo6g/noYlu5B/W/1Lzg05jFIqJR8vqQxnU7T40
cUN4mMzqJWs3GG1VBCprg4PoE0HCTYGI2gDIOx2IHREbi/HhNeREif35jynh
rXIrak5o0E1IeHCuIT5EHpf0rjBynL0iaiZ9KBU5Wrod0saHoC8zb4cSwXQ2
gIfj2ZxZ+Q3C+hbswrAMnmkD4nta7q8vGn4uQAUjVi484vvBdsRr1MbrCBc3
jrU0MoeR2FxmtcpkQfMhS5KlVMYM9Cz2G7g7UM1YVPaZcIdSfdrgDY3bISp/
ZTVVB1XAy7ot9QnCu7hDy1zmYuDsiKs99c2vuksEdBEad1n+biiW3vNVde/I
k7/KNcBohrJrT5IS8Y10vypFjx62c+VoSPMhk0QQpgtD7rIts/auZPbRfMRe
hGfIDFPNirvKYW4zXlqESsQLetIfHtNzY2LO/LkXgI8gIF3ADEcheYZnNaYX
J1mXkg3rLt5lZyncAs8HJlcNdFMxs3U8d0sT4NHhOUj7NIILjzWkGlpwBYda
0KmR6MC1V/G28f0JwJ9Mx79gKt2zmxMm30qq3DM2n2TLZvEud64Sh96m/uY7
KTa6ZEdvuQLlv6fPuSnXTn/4nKb+O+m1jXgqpUARLpjgPXw2oiM7FzP9JBod
Q9fSrtZ+iN0ZIySnlsfjpnzMDUCVmdD8SagmkrxrcAiPtnJD+KQ9bEq2K5NA
u0+uvlhdRMjFsSQBms4N9oFDq6O0hhFqJiOOQFKm6ssobPoBh3dKtcCKKygb
EFvWvIBVOdpqX7cM2bH4q/yW0InwbsQPxpg5/VW2YGMLYa5dW74jGWFF9Z1H
qS8wRi9jyqh6wXTEkqJAMVZ19d6utWBki1E5rJfxxH/5R8/L3iGlGokKBzad
jNyNduEQqHizovXsDmIdU5TDLmLIsu1cmsDK5/Ui4dGPEjeMMR49Du+rQED2
mR+8ebMKcXattuPgdyNgjAeYcuSYuVI3qXL0C3jhdTVCjnVGmtNk9EoigxlB
RebykOEnGdxf3lH552lZJdd7NGucfPNm6yKVsO9kZxiER1BqWRE8jV7OlC7I
BsWj+QjGsZsv0E+GQBntcYY9hm3c9TRbn/a13uzmy5po1H3DIgg6P1vsPUFI
mMCdrKW2ct0HA9Mwy/9JuzHYvOqbzs99LP+x21cUWhWVIlCpsz14+JoOXFxl
Yc8TAiNyqBnWoLL0rqFCDPQhpIV+AsCc7sPUgu/Oiy+LJMKuZDneEtWlkZef
RT8QEh2wrSbnIR4uDDyb5sjsAo69X38DW+CBNoc3m6it2A0IahhxM5FiCjPI
Ykl4hZ0I4lEQTGBBh/OAR/KYSxjenCqWK2SAfieyL1vvWJtgmHB0IKSPGSxx
5/iIpKeNxCuNfLxXrhaiwxh2YRCgBTPIGgtcZNvob0dfnkvqOSNSIfIxvVj8
ndim/9Q1BxssAatpNHV8fo+5J+EdBnBaekNoip7QRtXxRmvQnlKuHL7whl1+
ueaAWqN68q5qDqc0KOgy+l1GpuoRtx1Nywhw3DKVAbdy+z5IK9ANT4aPhO+q
imRAXh2p3s7qFvZMivwM0vxWIr1WrMT7NYQpBnvpi22RTqjieoE/JU8cXOUP
3x8CWebmbFLptfJkgJl0xzpVZuDF7152YGSi63vMsUTDRYAcHA2m7ZbRqUeM
k+Rgz8nVw/flfXq2Q+fDGoIr/rDidlBXhhYbNJtKzzpZyTg+fw5nU816BnED
3WSUMWFmARzP2ru5nD0PYkKEokaAJ+ZVXtNXndkAZhkWmlZlwVb+wnOJiJP3
hRPsw7UVXqqoDE9VWFLk11EOtAygdqgamWZKbFHDU3GxRNCXz7p6HTVJyePJ
WLvzpMDxRgdwNZlWwFLF8J/howfYQT1srLAsvFfQnHYgINeSShtT+UBB69yA
EhIKw22UKYc4WFd7WBt235MHIm4FLUEZD0ITVOM5wuctuGsh4O+1V09BfSLW
o+mIJeR/rsJV9zPPwK/Jq5rzgzNhgyPI7Btrv/3eENMJNd+CyjvbSQSUu/xj
GL37uZsLbeUedVzQJMfN2KBHDpRvHO47MdJbeeXgXxn0PaMCpjucV6KloVzu
FTJHcmSVBoImIA874YTasJrp/J09/wNHFpmhWwJ+Vsxb6Y5kfoQYVZzExe6Y
pOXZA8kVr2ImIjOMxlPYjwTICKQr3WIW6D0CKszoK6F29eIfzjiADPhshc9Q
jQaaxLiIx5YqITALM/Ge5YxilrGkAc3OrsmNU0OwjnyIGgH9HiYjxp6enVJv
iG2f3ItOMrXEC6bb2tPD5aElWiuFw9hxhQsErFR2AQv16wCN0X2ujBea2fpm
e41ymhlW/cDQWLQBLJI/Bjgt0DmAvlABhLbX2LwzvTulIPdAQzLQi0BaJWsm
WlCsLqOPdawQw/8ZP0UvfmMmTnFEdGlfJvhjFYE69lAKFsMQQ+gZKlbdAi6A
iuOZ7uOzJh36w+aXPCV4ROlJgMlWwq065RF8tUuFvg/9M7MOG3KLGjxs9kEu
iqCLjyKYglaAQDElu0sG4MSk25gMgRTNIGh6q/h3dxfDvJ14kfntnWLtQdPf
JRO/sjzSGdP/kB0Y0E/qyUJ0twvQZEDeD7OImv9V4A0Ld0iwd9Zc0FEd8l6x
EyK/3ZUllFTIKvx/5Fdq2BCZBCFniAZHohuggaSlgyLXn7C+aTlwouNqXmfj
Nhu2n8SkrensXsxPBqukCKumLz8WzAL3Tq+XAOcLN4udXtMjK1nlrXXjuV3N
rzsaH9sVw27gsji3qQnXJF9yScs/LwbY2d713xOBVrPXaZH8+pPz8djaB48p
51F+JuqNNBpV81rYvQE5E/+RTf0tivrj++hxUs+jM5rC/aKUBoC6sA0R+oO1
Xqf93Gn6HHyvMErILdHDQsPY//rDPxwZDIMpajAVLTajFxb5pC8KqCJz9GEj
riv+02lhOoAsYgkOGQ+600Kn2iLA7uzb5msExu4hI5M7znLG4qGZorgffYWQ
/4vegrMTV4MKI6Q5I7WiloLWbNVuagqF/mcWb3fYg00FbqfdG+gKLtKi+sKD
j8mFUhCYACVc0OOyYzkN4EB8TwoO/h42oQWh624qHNZQByXwHm8Wwxo2Rq24
ck34zO6Fu00LO8Xr3Ls/zybb4F2ipHgwiCVJVXmuJf9qtM9Lhhzm8TKPS1P8
3EpP90mS1ryzoSVKWWBy5TMeKBSxNDR74n8rytrifiCFdQ+LeFEO+t5djdIJ
lCm7cnWZJKEJBvdq3GMq9Im1by3Xxzm6dshfVyx9VlyBQZx2G2rJhzhpzztD
vvSSK0wXUy3v/c0JCDBJnMEb0+oTiQnBIaYM98XvjlKVSdfZ2irPWI7tII0H
xUI1tqIBvg1ujxJc517/abZG0hw6PRRNmpKato8eaXGHwcwHQMW8t47R47CM
xCaUl0Y3i+eT5mOjZGGo/ZeIgOO3hc0lJ9G2P1NbLs+UtA2OZM7U8r+S2Lxr
aGFe8uXIrKA2w45WeYqI3g3YxMZs5fqnIv2vru4y+/YNukigdDPy2pO4dgca
5xeqqJJ3+oSnkFMXTcVM67Dagy2IK1SFPwKqM3lWfZZfy5NmGugW6JTFWOox
3Fzh2a2iW4Us14Vb1fvJfL4jZJYyFkEc2cVl5tDRZwHcp1w04UM9nrFjpgsY
8NGcNEktwupdurHy2fh+IrKEwCjUj2H2zkRcLUNl7bxdllmybRFHMFoUYjtp
xwbMFe+6MI2RTVnneT+wdzijszQ0hZ/w25Q3BsFLJmGigqGmsmnQgsFn9w31
6OUPQ9QDSf8mMZ/qbGaLZJilOg9QO0cHiq2x70vRKCaFMPnws8rvkVegLYcO
2QCTP1U3byq/6Oi5Ro2HCgOdCgjwHABYoRmfjujWxibNkqlP4KqEWli0eY5p
jiZO4fcMeeu3dDDUjzl15B7F7NUwW3XfYD0wng/CDZDy+Qb8Db0m4nHisqHf
0dApaX9+gk0wQgrhZWFRjx6DEcuxtb8JVpI1RjBl4KWueVX4Sb0PxOIN5ueS
ZzjrzVfd4O34r5k5RONKfrPo2QobhpR7w1OF/dPbzITmhTxHGR1hHQfHz116
MgU3Cnawsf9aR/FT1SlNPTdGboyxR36cY7h/S4i+COHwT4YElprBY1VXoDWY
Xy8F9kMZn8zOWu/EXKYiv4LAkTgRfMqd29s0E5N/dG+kSQSPwJM69Mq12+YM
fTEe5sQn8a8AJEVoaWSmTiBwaATWpFjdMYN1uqf/B3vWiX6f7mr/AxKx37WU
aICFy1NEPLdvWvQQyO6SkmiIljqY2i55amWLW+IwBAhawdFjcDEAKrrUuYJK
iGQLEMNG88HutO298Fu0JRLosiD07ORLax3EEZF+xp4AgVcjC8LtpHxuxe3F
v+LS0AXzhsGLNbesFcDsN/shRCTdB6Dor33X8MSKEDqOaOJ7apP629/ItQu2
i9DJoWw9MKxVNYA3eg4N0vzXAzi+x0OL35EWXY6njZhsntHAFPO/29frFRf/
WBXx81cXbsJ6Fa/6762RB0KRyBqbZPr1HHxpU0YTGRXifl0SEuvlZEXAgbgP
cPtNQoWsMFgr5OUvZewNuG5Dd6SfVmywr157aDP2xY+4jtizj2RVuSaNI+ph
tnqR/Ox2Gpre5cqBlh08U5pocE8s7QSbvaFQQkMNowrZhs/XaLeFzQi6zN3r
Eg1kgfbIErfp7boLDTJJOJq8ZXj4Gta/HW7hMBuA5DsrFSfadKbCerozW+Y6
8alhRzDyB+9n+1XntWKyqdBXENte3e/EgHGqveq1n4v1Xae/Zo9e5su5moMI
igZh5667UZ5WyLypwjnijEJpObs06o1hF+n4o4kce0VYloq4mQrgxsDRpHnN
1/o06xpkz/9iTl1T0r7Rx8ef6rzYtGAkuWobapP/S7pBhV+3/H0fFfAvEJWY
FblK1s3YmMPcrioxCy3l+/iEgfK952MM3MnAb1i8E9UF+5zrqPIIxJR+jN8u
tvxBrktriIZJJibmWUallmBwCTXNfiKSZk71nRWOletHUNe44r7R6QR+q5lk
udt39CvMQZi6ryNmPXAG3kCmE7Tf3eZlncfUGqFNARczJaoabzIzDWLtpIIX
D90+NFAqLBLyc1wgQdJaP7a6652si0YusgZUIz/AjY9z03ctPVPDR7Zg31Kp
GR77QNK7TU2q0wFBFs87ktHLQaOtyXQ4cHfSf1nKGcxyQIFLyVBh1dneas/6
WexvE2OZ9BLMI5AcV+xQWsmER59jrxLrZ1iLjRddWn7svJpHxOa3QKI0H6gR
+89pNfq2Mbx6priOUv6PVK5I5gvUfjYDFHD8DhxJcMD1N6f4VDfn/B6xnPWT
Aff7IHsCsV3vgdnpvl4nH+Q4e+aa9u6WH2xqxvG/bWPxDDsAmZmp27dQa6vD
6ezvlJvFpBat2Zrnymc7ot4XsRS6J7pn2V1jb3r8y/FDlqbt53sw6kk4osVN
G0jQoXD3MJ2JuBOLMo/0XWLar+9LFFpdS9VNYGHaiLHzF+CYuGQh4h+b0Kcf
ZZfWPfEIfzdZYdqujT1CfWYRDJOm0L4GFLE3h6EWjLC3+YpGBDU7ap/3NnOU
HAVz7lY5N81ngu+iOIDl0c8YSrpDH9iWXiLjQaapOXvLcX6+B5AnvHUsQy07
hruQCI/KjwiQP3yu/RxYTgRUuppzf3aehqUNM31Ta3Hy2XiyCBxKu95ulYo0
qgLVUDdzEsbMEfMERGOV5s+po8XmfSu2PIJhLqukSsggX8qQX8CYWsbeLOA7
uLtkjiZFwD5aTVb2c/75yku1n0b3Kyslrc10O/ECYHngfS9dvtsh41txMzF2
hcUoBPuXwkZnZKQbeyDO1jKadTdLWc/UlYc2l0/KPQ1XL0ziNr/dgLoIoQDK
hV/gXX1ugGYSuj4vlCmmbh2cxvxs+n3x4QPutz4AMkziegw7uP4lA43M3qDE
o9AxD9x9bSel1FIrIQ8C7xQ1K54b7ktfiTNydi4pXOTOYHzsySRK7EYIVb4N
gvHPo3DExMXAMzgYmtY9y4uG2fFJbDvFAZ+NjpivrHSJETtQTFynbyipdMQj
eXu4k+GHN51BcfOBXiGgBWUVzK7M6BhUIZ9tMfOmIiGsjVtmQ9FfdTG3W9Z1
V1PCjBWTILAKQNfqGuu4JQN7FPR+sJTc1399azkx+GKqqrap63nKz8Lx7wPo
oocu+4GCAuxNlKq2bqn3Ywpo4TI1ekN/UQRIcwj10VC9fWBHMZedc/fwRM7r
RdQoiu0R/0MKxmXqRCf82fqfK2AUHBf5lcZnP4IYUpL/4dIK/IxCPO9PlOAl
2NqHVjWJd1+2vmff7kdyQz5GipzWPovQR1GAn4596PgaTNehAOWROaSCdnZp
geOGiCRyA6VKWITYFb6RTxJJRnKzv/MVzNfm5YsIfErprFGd1kx1HwGm6tbK
a/kgzXAdBppzv7MQwqUzTzOW1BNja/vzdpsJYm1k9ypjxcOspQPqLMHlw/86
dJLF8SyUzfj7bquMkH6+hXz8hxQ6bFUnisSWUNpZfdCni6+NBZmwneQp++Tk
rPnVlJTnazU0hcpXvsNJXaU2RFmzqWa7AOuFLP02z9BWBV41bF96xvassB90
qvmi6+XO0LGLLaQV6aJ5bBhVbM+QRirqSYgI5/BVWPa4HAIxKs2b3PCpT8tY
zl7/tez607jNXXq/tEv1ZKStdGg/GFXkt3dCVUjVW34R3CcGddiQR+UsfDTC
p0kooG6qwG2aP7PFQF7qs3ITjGNW3/DLJSZX4umWSbNHxE/85SrQSh0tJSy3
plEF6ERFozABCEt1lqscyPAH/r9vJcKOP84ZQqV0cWoCH+n4zMkM+8gD/GCA
5EXEN/M3y46GBMrCRheu4qO0AtdN8tDXLd4pWZlzKvckp+hV+yfySzYn5Lv8
/kPL1YvX4IRDRujZm1tRcaMCcD7behU4YvmjlNXevZByZ1/jixFo6vlh5RSc
UmBb72v7kGqTyV4OOHzmgGXPWuIGsdgF5EMoIFZDDXjuL3N4c1YUDn7XdTDV
QXIB3Sz22AIGwyywPK8faQvJcPPeF7o90NOieHKMTeLV9UQq0eur/Emp49D9
96Rju40a5VBJiJT2ZbYVjqDbS4XdcWQrxM39smkyAtwCWbo3ZSFCtCTwWLEJ
rb0lefZxRdOcntBn0aRpc3RX398hhJLqkCIIpZnrFhW5RjoKeIDD5b8P4AM4
zyy1nfWmenBhC0nIm2DNun58DWq1kvxM0Y/0WUKoXeiq2Yfts9JjPH3MFNUA
BrlCJDYQRfR9rxd+5V6XuA5IVDnBRCto9ikW6L9vONMtQ4mpHMXfGP9M38NL
BKXW+Z7ZJjLRQ1ABbvD5BaJeiIBXbtHNnGeJE0UXOIuf5NOqjgiPU+eRctEc
KqVnWcF1XT6WeDSXRC/FW0lUvlBpsQO4tg7r9SaKqoFrYUmOBJYgJTpgYtAe
kCphkmdSxBYpEr+3zwSAkHTxbSF8HhXqio/3d7TaDcoj+Y7bn0btKYWcKUuG
vIRMNo9eE/S7fQv1PkcTPpUc+R7XRQgGr8rjyr7qmmI1ebmNIOQx6+2jxjb8
3u+WwVJ4b+LJrVP7F5x41Zt6RRxYlfRBv6+b7ZGDcw1ETZJ5dhbVssG9i1v4
xweH2htPShLuvkWs2OjhVZ895OdbRmIkwA8PLIJrh7/VmY9GdsMmb06eIBCM
mdwYgsr6JV29eeNWmwN0E8XnWT1ucO8vBOhdzD8zXqtxQh47dyN7Aeai7WQQ
xWWpVfFphBsycxBJ/z9hGATc2ZjAKKU+pm8hN0/ozysqsFgx6imC0ID2xqAu
ZdtBoxm0P48al0gqhAarJGAP0+EKBroQaoV/sJkooD6Kr7ikUwDd/39N4i4j
Pg0dXkvKNoP1SL+l/4xo7gzIHAtaON+RSlRPL3nTVyQtCOtCklwsZkRFi3Dj
Z1QVvuJ2ojuo3alkXAIzuuauaWjtE06M/JVRm2OkADxcaNdfbcuNTCuLBLlo
nup0TCHRmMyyTUIU/vx+5vaef8Jv4ZBBKjy+XpiuXWibOGPLVZdhOcafI2Nd
mmbA2bNNJxBgloTm4AN2m/s9WxZQyM0BvngUEjfuEseEO0lF07EbMJXqYfxI
6AgcxYHi/r+Swomvo1znkOnCkE4fi4/M3ZeZiZETqXr/t/71eMVFzmdeDjqX
uY3ab4Vc5rIEgzEEgrSHR6fxgD6OTZF95hX9A0jnOdXBC6wfSFP6OyqcOr4f
5AjDexdXUiYZTo0iOBiFqceooFqDKCc+oROe5OU4JiQXzHaIA90Oe19Fda1r
d4OJqKWSQ/zDF5U4DyBExl9TutTj1RPjgoenF7HU5cJExCU91BI5oS9q10BA
1XGcqJJfJy/9lsYi9Bhb0Y8jy8bbnsngMlh7DBez3jNY+mY28vxQFXdZg9P8
xYI9Y8RoK6Uy625qiuJKCQyUWCRqoXplwC4mwunnCTO7jK9q3rEdnMjv4vek
6+noqiz916g+EeQP33DW+gIaoa0cLBIHv/oMEoqquElxPVMPs3sQ4+3GpV0h
wI2PtsCdAwVdcXf9hf3g5XHzSjGaWGr4eFiGHsRx4Vt/kUOAXYoZFpqdplpF
Tci0sj3YCD/LNPWrxXJWw0SJc7AHEEwnRY5cA8B5To9O2IfEkcuM2v/pzc07
F93Wah7nEdR/YwPt0u7C1N2kiqH8YvdWhh/MDal02p1046xMW4pDS7sXUFA1
VubhJwA06dR37SQYIcMalG5BdVvx3+6lNd4Wbq8kAbVBJrhQ82ltBF4euuMv
DkUUJO7UfAM4fGR8Xh2XYpVmDG/a3kP0AxnX1M5STlUdEecaRQLIDqS5c3Iz
P4RjFK/cmO5mOcjlddDYKbUVVKRlbZSIZYpNb8Leh0qFFDKJCXbZj8Yypoy/
NsWUl8ySS6ZiyGPn4myLGW466zyDwJwNLz1KE7ureG9LZmyIKTj5shtrL++u
DZg27Ow+QKEUyU5JV/I8tLm7/4ajDG0BYM/EqLW5JGJLZCpMD8VGnBSpEnjW
lbUKAgPISCVSlaobC8R4hzsGq09jWko28kc358otwMyvI3JJAyCJ0fLTe667
KYidnbK8rdy6qmqkWDg5sZ/mny8KVDFdeZV11Dca/PLtqj6HqbM4OZwV8X9C
78dNmG0U2tTb3CYDWe55nZ10WAjJcw3nrPZQ7IX5MrCOFK+9X5vV1e/VcQDz
sGCjHWBEPj/hQ5hRpl6Y17VyMmgGGrfPBQMdA4Xn4M79/zVmWBt6jc3Fhyw3
dp3mwGxrmNjCmudr4aU31ZYKWfWc+bTbJjOTKz1v9JhiWVhvtG5CMnHVEkzG
mg/sm0uvfg6kQcXS0TKbftvU9DO6i0gZ20KHng3IRNVtN3SF1uCmhm1qlQvv
k3U52it5MlXyxsM+54FhE5nMBg5caCi5pNNMd6/6kp5eTB82RGzZ+W0Cdelm
7hbCTsKBP2Xzg4DfAMCISqpXMbsAMZ0EpaGMUqf+21LuCdwp5syQ/FyXsyFL
uxESkF6mOX5sPShsdF7Z422sHbd+m1DgsWicw/2J7Kmo6L1OzcwXsBj5v3oN
6eWLvz9G3XEb3QAmtZxdZZWjmevC/4DOY0ZUYoJ6j0ZtHU2X2lJ14YNXenqI
0WECL4m4QkyJJTlLTc1QbkkyhzrHgyeFtXzuhTAT8LxWYJq1V1bWIsTy+6RI
iCn2E7XfGf3dcx1c3G6qzvHJczwDZMsH0GC50r25Q6A75Xw9dLCOqCPPA4M3
1id7ieuXjy3nyOaugnUygzlMYQipbF59RNOiO7Gp0vNJxFbrPFp7Yz+21Nde
/iV4nuWdzP7y+ozXnS7NHP7KFEJSXEgxrTZVV70tjL31HD6tn5CFGAxBBkHo
wwTZvbt1YB9xGUp2BAYagsowp5C1kp5eui3gFBZybmXdyP3mOZVXDC1TUwLI
i/tCFC/eYLbe9x+vVa1cvzCPsvBZ1EPzFHAyLs5Ccy/U20G5hiEhIcS/ay62
VhkQFc28hGBYbjYQ1BEAZpQcZA2VLas2Ga0o0s7toFTYFWuDTDLPm4bgQ7mP
yi337P4BJTDbQmFikYZwZ40O5nlFMGAe7u/t0EZMjrmOMAoeavPN/TiMRkAA
UsME2fTB8gyj9IyRAxLNcoXl6V76LpuERLX67vZ+uEMOskyvTmwbP0dQcHJr
D67zx8dS7A+ApjP132F3tOOKhjG8r98cCDpAuLR9RNC4Ql3zcqgzaF9XdjCh
hDT/FQVcqBS3Xu6ftBGprhi/hMZYiOxosvRpFMVNss1XYhiZ8jR7HpjIqzBn
0bLnIUpzQeEUnF7EjwGx1qH1hg0QLjSwjl1fZBTAstl/vw4sZUK3v1Sgzroj
4pkV3KbMsDFlHMkWDJKmWa8mF9Y+0Oi08nPBMtT1Qbnb3vhiG5FcRc+ojDGQ
r3wd9Od7zbSuXsr3VQBVLhNapOm2UjHJTu86muAap9aAy9m68Vk1tAQ7IQjf
YExagSKZV53t8YxbMbQqnAw1ZrmFjKdyBSO12GMKS+tKwUjL875YJ9jeJkwy
9g1rqShEf54QkBgtcakCsuPDVRB/NP99iBXh/1dK62ZB14Wv7cOMo/6zTMS4
6BSP3fpQXfL8MA++qoE1DkDLEys9INOjI4LA+Ulgkh6loYzkL0AzmrhrVcgP
g0xW3rLHykf90ohX+1w8YMiICoiKEa/vAXFUG2/uUqMZfWoKeeBzkCnNprvH
j7ZUmAyadLfq2PJ8Q0CPo0YVcd2cFIWlNxeWRt4kEzpcZ3HuWjrIWMVTFZ83
jv6JxXuk1sOWb2YncfhRHzHgqcXOXJ/p79l/Pj3pOz3g3+72KY62r6JuOxQJ
8TblEQ/8LMy65JlqdXMqxbhKpEDiFOI3j6RdQNjRrUXo252Px5AqOWKCfhm5
+gVw5ipJNA+1TT2+iJtYO8Y0KGii4UfLvsTjzPLgB+fSosInvqJO67CcPX2p
UlUVVdvh02msvSpy7oL1Hj3Wsac7hMiuUbPxc/zpBcs/177JST/Xtrlowg8w
i9EhmNEJMXIKRlMBpxk4GlUm1KwzbdzV8YF2gbcn08TzzIn1WH0kzW+6WaBR
67dNVJcfginLUPZ/yKX//QfZbnnLe/L9YFFetCn15Pdd0t+etEAmLzUHEoMZ
bmPF8zhlXrlhM8zXqHT8iYkrtUG8DoTaUaUvwgN1lHko6e+bfdyOYgod0sMv
gkPWLDkNBDcR8NvD1gh60HjgWSwAqzs4NGsZlFxPzjPr9mzM328Ozm7Q1JRV
lb8XD+JlfqWNxGEJYbjGqXQbkMJ1vC14aK5sNqADHaevXNKMsKm4CaB5ll3T
j1+0/EdpZLMh/t/4jm1Rh77uWwTzn7SI1qNx2csYhF4PvJmxNn6Mf2/pp7xN
L0lyr4UwpPINlm14NrNs4qeOiP4iK+geXKxeOztaX+9YmV5wq2c4edppTSLX
a0DlbdWvsYE7WuHJNDDTjtkNWEh9Evh5yrxTNadsQw3/quvcWUNKrFNnM+j4
jxQ/uPh9AbGh0LgL1sN8FG6vMKE2CxPkc+fjqxtpfgdqxfavR7bsR+wevtvS
bDNzOIC3YT1cztjnoijrOJ7Iq2i2qtWNGXm1Xh+fxGKhqZ5YTh/NgCjEvavA
/7CH8xqThi3sGIWS2+j3M7P2IXPIdFMcB2mduFG7+mA2TstaDJDz9Iov0ZNV
6Wug5vKELqv5VUS8TCLVG3ktEX3HFkVL5u5cD/j+I8G+ipO1pyoi6eFErlWu
YGutoi+WEQofEO1fKmQwN/isTdzCjS9HStVb4r3fFhAwlvbwfinORp4VRtOy
kdOI0MyQQfV4/TMccU+a5mjG3Wsnzqb1nvX2MJPoXqlFlHCtjYb5eswxhnT4
leqwW0s6NBJ4hJWmNGLi85LPotrzU3yKfSuUfzlskJ28/7i9UH82BxmIRVYf
WyhLXMBW3dWFiOwz0NzYbj+5vFTL2VkOE/cA3v+XVRhOSOzyvyb80/RndAVH
+zMj35GkERQhb9XJRLTxjFPL8Sop1Y/MCiWRJQIAiNvMLXht4bQq/4BA6f+i
HNcTIzp+VMzaLjHzx28L/GWsGQMwYczwiq0AL86cK6Is+80HrlTqX31svl4I
I3anUacHpeWnMkn377VC/uPqF6P6yStI2Ph4D1rFRVWngURCt4o7ZGsipSjj
wYInkDeSq7l5YDISN8zHMm4RTlst7FWWUTTUkZ0KZyFtDSidOv2jFUc8QcJW
KXZe6En5oSVjJ0Bh6ofvH633VF3DQK9bH0VZiEsMP5ROGaie7/Nsn50rTS47
Did2WvFS5BvVmPN/peYC2UXWQnOr82VwzhEHc4ap/6H5mR8nbRmR6lMRg+Z+
e7QD+CFCQ6HA8VBlWjx3H6Tykjs7yRYdKshb7pcnksT8l0Uvd3/qR7xOX5Xw
XAIMPv9QVTtf/XiFFRV6pVxUk/jmrUHpN4uSHhTitSJWNZhThvmTqhIKiC9k
rYgKJNZWM87yBtksVVZ7qw7mGcXPzHpjdxSOc9LrmsUvnjgi+jlkOogTkKX3
AOWiwldPti9udEC5g7DxwVDSWSFhoouhqyWSQU0P1p/OxBPg6flD5QzWVXt6
GAwEY+EHvol72h60czpyRJ1KN9YkFHm3KIIaTiEtNsk2Wt/q0LHqYKA5NJpM
6eqPSVoOXfgqSjrpmVsISlPx0FLwzPpPpmSiw0B1Okx96Vmc5y6RSeIEiTSk
3qM3xClGY6168bwy52FPhEFPu9+b/12r2GQ7G2eoKtvYy3316zLvOU/2BfIl
Hh8tgVajuzI9ZnG89yNz+6vFibvlug7KaeytPsEsV2mVRXzzo5BwtLP3/+Bt
X8HXWYMtwGkmXZQyEAsDQwBrwsDxP6KBRhpgZEXAyOKUcRG1CvPnb4n85FWh
7IM2Yp0i3pPiZGxoU/KEj7T+69jzl9KK7PvoHaWqP+4/oL4yxXrmJyuovnWi
mR8CgxUJTRBeMhjZkmts22Affgl4nFuq17bu0Iy5SL7kfdJ1PE458ICTE8JT
/G3slJlH3IXQIggCArEDKgpGKTICi2aiExrr9Iom/vE5vQ6FMrYVkW57iXPA
O51j7X+EEmIYPpTtRFfNilbhfS/SvI2UA7UKztR6K/QSgWqoooiYqodAjnKn
YSB623VgAw5143Mev9u/vyw3E3ze/Jxpil5+1R/GpDDlReMViKhc84V6xV6L
OqSHYKtQoQIMNojrMfmOc/+CjOs20QXjlN6AnCr3CO85Q+t2C0SlRPC1sg1P
9p44W5e8Jz9DQKY9hQ6KVj/pVhbPRPd381WeFbXcrbOG3rVBRMpFfpZIRrkW
ov5vJ2blJKVjrLy3Qzcn8X08fzBM4qMhAKKfpPB8ujc4wbxBVKIP+abqrvsr
jVVeXmQ+/axTt+WSfrncaEdxmdSSMnjgdenPhqnnBqA4oVbFRlPpiKFAN4qk
3uRuL/36L+c0B/51WzFdBdt3N7S+LRMDI7FDMtGn+b9/rwCUCqkdieZptUsf
WUVcSfeKIi6TBPSiIW5Meh8CGXuVXxv0KXrGi5rmars6SmnEVB+yKwXBkN8V
xxCgtzcRYmUKeit8nN/zlsAiiWKKkaNz23Km+dQMgsLhlfUHynRahKLuDMLj
J8QoSAfPJmtUOjgKd1uVFVJqjwV92tEPmvOenbrMu/Ea+rk0LOeGwL5nU6o3
4mhoqnciBUmBbceBz7sQFtbwTHE8ToIG4SK0aK7vUdXwWIMF6wn344PhD/Ux
e4473krOQ9SO6hm6ppvSXIT+5ZcOhJ1rKY3V97L+V9DHTTCivGnwtnm+4y3t
BlruLuqqzbwL/7xSRkUu3ORmv9hefAI0MLGfsWbPtMI+D65YWPW44b75DnMy
rXUXNFtIRFMbF++jmtgHT6bc4JlOZwEG5N6uTRnN8OxwADEo8mGORbGFrvKG
Pp6KKKkrVmAa4RLH3+J412wgV/7O1wk3QxbqxUAzvHiWTpAzJAAwQv97a3kE
lF0nqKNLbhkAxsX3zg13KtEn2M3NMXYT1VOkK9wH/KaMeYy5xRLXuaZI7xmD
B/MXOmK4kUKG4Q6LW6l9YWry0ujE9oA8ydRrWKGpEmVzinF4uJULU3IThaUc
LX8DR38vNDvzZJQl4nvHvfunud1rMju3b/mnft2vZZ6jKQ2D2cl8+Fn66szS
ARNdpNfbhMrtPp7r/poN9SP6xmXGQ//2qG9gqyuP6RAh5XQU+5UBEi8BqDOp
zlAqGB55t8sgixEkd6Xm0xM8O19E7IE1RhgCsmR/Ht6bettP3yL/N0r2oXt1
v0E21DuzBtNfqrVNUOKUIkWuWJre8K7XZizwr7NrhFZzJC2yUMR5BPw0bwqX
iBLccO8C6SBCF18oXKTgpfgzU+yllUT1SLjop62liTb81vOTkv4Xkhh8Embl
itdPpKbchYJnb9HjSbVr4ODGeqD6FFGJ6pUDQFrlN+7Yin4UCCQJV7WFVTWz
q1/G1KSES8krv/sx5QpOC2c8ujAnfrOOdtaRMv1QF/7E/8x+44Ze++2RvKzq
4f00zRv0VRuXU8kDpp4wokV9B9aJwv1Tw7t8hV2vkPmu+RQvne+/A/7YD4uQ
hPX8zQFe8gdSG3zJdC77bZ3LaXJhU89xO0E3tXL7mzUfaLw67hDjjHlSkUsW
GRQE2D5dOligmhJM70v9/lNrjl5pwFE9YQXIliiU+/wqH5riWxiA2SVowIOJ
FrXYAYz18R1jLAfJSa+9I2PlftHl7UQouWMTO24d1YxqcU9qK/+W9ODnZZwj
q7bl+SB06BDotUIw2whqWYR2Cjs4w7ahV55got2VeaEfeMeWkqqtrmELn8RY
lSv3C8EYERs46zITaaFFHFLBUplWTBZE9XP84DQX3tUSuu6DHhdCO+t51cwQ
2ZMs1VpU0S8hZGzQ0PsAxBuXKxAZqd8ncS6nlH99FuWYqF2Q0amlZTAGfHVS
mSNW0BNsCF9fRbCJoBRTJKEX5e+xjF8MfS5l5YndTZEygG2su0LcM/JRjQEw
XmRrsrdtpfPsYW8sIKB6B8C9ngXZWni7PpDUJogVCGbQJfwocBCXAXCSWjzj
Sd+8DRrzbMAasYc67uYr1QTIBlxFmDoSyxriWbnnBe65MCNCaS750NyqXC5g
XKvy1/CHTYSGHRt1FAkaJf25wyWZEfmpgeP6hmxsC4+m6vS2cLsqM2Uz/gR3
Pp2dXWEg+YENIMhRAfxL/VHev5TE5oNHPHMa49mQzZVABR4Ly/rgSCzc4lg3
WYvLm448nfwojLdRtLB/2kUDlPvgJxfLXWDS1+ZL3CxA6ZcY4H4gdFJlG3pt
TdU2I+AxlgaRhTZdy8SOnuvBHc0zmAnNEQZS9NFG6nhpybAhBRGib9orDQzI
tJwsp0pcxwiqD7yOjdHwKHg5LdKf2sXv94N/aCb5BvzDM00ZGTzcx1d2TkGP
qtihrjGpCoXb1P4upvB6ZYqfimSvtftmUDm8O1H3cMCcccnsJn/ofmZwSWKd
zURWXq+xP7mZcjLhskxBWin7wnMHJVigaCuT3xa7OKDRUGnFW9r6pwyTPIM0
gki5J6GVImg/Eja3FthEVlwvn8DLL7R6X6yQ1ilV5/GmloyAjkx34wtQVpzh
BtpBT8cIjfjS5L4QwC1yGhVlX7he+B8poaRHt9z+oy+32zlE/M8WREDKhTZE
17DUNpTMMl3EKPpi1ygg59IJgXeVJhvNt9jLrSsVxYe2ov8GSpXyLUYNNiSl
MCyXyo6d9QXUdE7IAPzGeBmToI7g3GQKa3yKON8jf6y9WelA3Rac8FL6zxou
uET+vBnCyD1Ui24oSgztzqEkyuR6iz7f6tE/R6AONgHLmI4GUsNbaCaxwGFN
OpT9+01e6bHPNDsefeZ2MRp+UI7LeY63NZchAm4KhGq5FLXzrp/q5OUqvuOg
+B7TM2w0OVAg4OnWEyAY2PeiTQhr/XTHHjQ4+iIIwFcumK2s1+ilOpVFjXvo
kFd73O62E7eqfHdn2YXAxLOKFtHUrsJQ7aEgfYWUZoeJRCrGkWoZrxo559yB
h68eJMFYHW44Ry+TL87YJS0htbWmPIUgRPaSVY2aFC4wGEkghJjbWtonRLLC
2WYnpil4JGTxf3jyjWY1gaUlozIq89GRodZIjneJTqoi9gjsEdKcXrL+76cr
K1cS1Een6W4o2v+OATYtUtA0WjZ+TdToMr4hlBM4gnAvLelhruxJZSblsbNy
Dh1OAqcivqJ/AKJvCSMmrjSf05On4ZqrP0nHnZJ3aPwVkESfHpoplPRnOhrT
UNMfwoPKYDIL+wh4YF3PHCCWuiWBoLAHh0XaRa2gXwgrUGeaSjEtuZXc1wJw
Yml6CzL7NEITShg5QvgYHwO98MoE+bI5pj9T0N0rBzn+mQFrU48FW5jzN0eg
zbMLr7DSndRYlIKREGsnokjAt9G7xcbYXdyurvwGMgsPV5S2p79n3/qJ/vB+
fptAmd/swhVplIlxeziAT2eVvh3o02YH73Oqd6tHCGxlg+CEjKB8apV5htVv
4ic2uDc1VJlBxOnVJxFgZai058/L6OMLnE0FgqQMd6JIBlni19210fqYhn0X
1J/2mpaEXHfNYZHQA3E6djBQpKlJISzQqrXGP5XQ4Ue9Oy9Fq03AZeK/xtgh
inAkYCA+wDh0v+EWReohessGLQZCyLHNfqrDcirss71PxPtpYo7BSas2ayUu
Qs2+wvHO1BIZhsn+UMwuQJ0Gy/xTPz66QylnEmXww+9cUpVeeio5et1jEpya
SBFCbkuuiVpgSpiHqNEJ27SKx17crolQxuYUJGxa6jXM0VS4W4p/iHzJaoNj
qUJ0pXm+coleovR7QFiq7yQLwfKaTykOJpWzMEbaLI0DYqHd03mA3DZ8O9eG
Su+R379XAHvOTnwq/AlTUTvj8RyTPXKahAzxdzjvAJjeY+Azp0Nq5aOXrBYL
nhgG5bJJ/HQGWncn7bpjfB50NHw5jQStOWxxGyFC9V0EBxbjCtJTjxgxg3EP
GGeKJnlhA2xHs6W6bgYI+f9LYKLr1rJgZnI+vHqTU/lIDuSHR3zHhTJaVcRx
jFRGyyXV0emjGw4NqclHRmDfqjqQaXrAOgt3G39fUbeOkpM8/zcs8sNojJA/
kWT95Dc7S4//IMU4h+vGkBGQLEa/g4pTuYqkhcZALODgiOngZ7K4sm8P1vli
fhKTj5/cfIZPtDtqnA+DlXzErutTQFp84/nC1WkxL9FeFgK0qf3DEFpSR+aW
Xul6jYEJIp44YE3kAGJ+v4ofr45w5tacXNxpwJNuaSm4hvQp7TI6fGfLuRE2
Pxy9vJBDiCuMyc6JQ2mmPnWhTt+1zOiV6qDXMRMiJ6nSAs70VXV2Kab7x4yZ
SaDCskjX5/Cv5UOa5nww5eMwePOIaXnxkMjoA327gBmd1nmbL7gOzsCe/EwG
hE+y9Ns/0QVg/wDjG7vYwOqYF7q+LmQroNNnY7recLnqtFYy9JR/Us99Rvch
Ie4vrCgbWBr0jEoNz8dtD4NqSqlSm/jDpZbG1w6tzO8ekQTDug24pvR7cbHl
1NL+k/Qngh26HDxD5hhXaoKBRI1+zKF7dEMCna9l8lwWErF1ogXTw9QdrHC+
oXGAXNTDW+yQCOdEHoPvProIvdGAOImEwTSWo0W8bDgP2AEkE+vXter3nYAJ
0i0RWFEJa0NtksvosafMUwLBVYre/7koA8CXSPJV9pWTJPMU1EDcVGM452b3
Nx8S9FBd/QUo0zXsRgUKiC36LQcm7KUhSmtCgeLpg9Cjb73ZoptInnw2VwkF
jcJfotJyrQCOXX2+KFygWIxWXx+oaPFzJX6NvaPGeyc0W/LfrcPJShsP3cnS
j+8au90+uE2A7sSNKRljqH0Vkh5VcXC84DkiUK/9sfDBbcHR8t7pAR04z4Gn
13mU0j/Ezd9JRaUJOQkAC/a+23Djsn3CzT3XzpGTposdVSLl5fKpKGg1NQoc
rfOLXIlIyeDhAZWgtwmQ07wAqpnG+dCjwOy+ZNdRSNkWYwfWNiY0UiRk8KsP
yrg2WdnAoEg89iIjy05OJEOoioAAdimXVFgJykXTRZl0vzpqcXyZOccg/eUm
o7SvoXyB3O+H3zUFAB7x5H0/Ls6q1CPfihMs2/lSNPezTX/RCnRN8V7jyHIo
H2mf88UGQeyKLrnMt8zjFl5FrRstA2N1lQmwewGfzfGk3vZyLzsNuUwjH4Ew
/5R+/kTLDjYTbTzeo7TbZh/1Cj5so0kFdftMbucEHPywr36wxMAfjAthNHSH
aUrysAFlmLJ+K1C6LlhvqTnPvKmu6AmT5v+6hYDjgdLNbYzGj5K+8IKdCEWa
TRE0YG0FQIRFXSDxVq1d3U5yu/BJ0dLBv7iR1jV1OtbbjXJdTfwzvBO+1E4l
bHoc267D5A1+RRlbaKNQEKHzrxfh7rvI3zb8WWqqZA+Y8VYG027Pm4VXoCFz
Y7/u0jpfkb2YvDHNEjIEuiR2zxCRoBT8QKth8gGgpVJSeuipVW1OTkJ/ne45
FzswjyQc+5SQdwOEogKCPJeVEmDG/22+juPW4aX+Vh7g+6q45T5BAHRAYXRn
0ibudngejp5tkzGWVE3+Oyur7YniYcaKDtU8891ElQ60ApDxejQzf6/bV8j5
HvuJsRsbc1N3rD4MT0bSWsmou0oIwAohu0UWcZWZNp439GffkprA7hAPTkFp
hlCsJKR4D2jkoe5lqZ2Qtj7o6lXxbmIRsWivPzgd1N8Km0AIMZ8k45mLa9mL
vwovnsU3mUjNUYeg8QatnZq8h7sHxPpMt6brDIEc05lupmC72DmTg4MoLurj
GVwJUYiWlu4PtSpi7p9LH0o+cJ5ncFi0Qnu5tQThng3o2u2vANVDnRe/Gr19
Nu8zy/RX+XpPfOECX90JFv2d/t6XEBgmLa170C3CNJqqtnmuUMhytU+g7cQm
rp8U82npbzFuM3ZK1gPitbBkqiisifKQRcZpM13wGCBIBgQK3CWM9co2vl5n
Mc+Pm+ju/+fGSUkUHuuu6Iq+sUbQ0Q99rzLHrW2DHWxwcWGjcAinwKgDZRPS
Rzd3XN7PXTgD3b1A9XQgoJFJayAuB4T5r1YOV8U0CL9c/tNUFrPC/+Cxzvqq
4f/aQPP53TbFIr/v0k0FPSR3S3Z+IoPcPyIUtr9HQdJmg1yY6EvgPmGfDP/k
RsX7bdvdEadjtV9K1FoagtKGt5syE49QtOf4A4l9ij/oKA92ZNCKb95sOQlx
keu+t7YrNhOXxBV+lPJHBH5EKX6Nh7FegSbyJdaFhHRWUpUEBb4bqClbn8tP
PnJMemK8RG0tyVFadHvD0We2F5M1oVvOuH9XSVYvwT4BX7RgUheLhCUXZXYB
e5VRpxspf3VlRAxkjFy5JcALl5QqlP37L96fWrkZ2+ykdGyi9dgJnXUbi/sY
A9ZBWZh9+HUyHDfwQV91ortZEb7iJcvtumPeeFz/2h3lxbEjiOMcGEc26XmN
1D0j5ibFkqeJLl2uB9ve3RmCfgXi8bFSq3P8eOtxXGZCkPurbut6+D1hLtog
wSElTKKR6Pmk1ZOM5X3furbdEpDCoQoqNrivAweRLt64dePf2PI0HGODHQUh
5ErUvqbYdfegfWUKrGVx9bjGN6d1izq6DrdGwauWTzFbsP3pDah2CTkU2ns9
AgBw42DQjbDgERxWgS62ALOSooKnQClqLFwAlvXxl0tKdaXN0ocj5IlURkEP
zY+U45Lr/swL/o6Nj99VUeY2n6Wu5Wx6QmCzmWtCktVFGSoQX030NFOiW6iz
1sNe5ul51eQBwPiZKq9Ncuf3EF7mqAnKXlD4t3OVZ22yPFXxZHhZnjXFTLX/
lzK8GEm9oVIq/ckA47bjtY8jUI8TG9Y2XHnROF98kBkPGe/F2+HFGc6Nh0jg
iLU25cc5KaeAZtS5x0OPMwQ3DHFQQpHzDb59j2uAnbzBZ5TDf+suW8RHRBtC
e1GaOLDKlYMsJ8aXLvkCcKQTqE6J/FQ7WZCsqt27YGEhG6eF82u/layaj9Xe
Pe3GNwJLTh1m1gxBLqsyiRikkLfPqYbeXAHKBNH1YtQGL6eDkn8jrYL7XhrZ
MkLfYU70vumJiczFHfOWQRjKAJeuXA4jQ5cvv0nOKmdR+G6cgZVlZZNQcCYG
F6iNbCZV8UUKvYgB01h11k0Fl+uKREQuwzbJTf5q9QFw3TWX2rl6tR0m8cpk
kXJ0jamOP3n68PbOHPIbkV3xTREvqaYzeBrkSCaJBGtnDIoV1p10mc4JG4EQ
l+kE3jIBZkFSOy6mGVGzvyDYFs1cl1av4jDqjwqbzEKCw1FdJcfy8A9h1QdN
+VSYDbjNNx0/cVD37SyBDJO5J+Mp8zPrqvjQbJ1tbSG7BBaMZ154E2XCyzha
Rj1Crb8HRjI+BSIbDB3mo+Xj0Se5yymrMnkXYrMrkgXFHQ0zrpYORTKXBaNI
eKy9MPSRmPgSefWktcy8irCWXoQ2Lr1DkvNzLeBnFGyP8RIwtgUZBV+BAepp
O9hQqoiA04ae/o8e4K9L24wD206gJRxZz/NO9QbW/MeisLQgoMy8Ymj4FvY1
LCQQIID3309pNptvRyIV/HCNKw64XpgiM0XjLeaCsKWN20URI2hUiX5F2vnu
LNQyjhsni/PO1+/+JTztMcK2UA7sJXjjanFc0lAZ/1R8Ju+JUab0HLdyBGi5
/JxRv7sLMvltEix2j6zIF3fyokDZVCIUrVcUFIeEF+JnGdr+ph4ebOxNLS4B
whIhvKBaEnfu3dl0GLQYR6ciVIOWT9BoHe382d2iGZkmjvOYAvANhqt5v4Mr
Ml0YC5KIOUs3OFX9Mt0QziJZ+BLYFCAZOlGaMpDgkvteR6IMTyjPaGvxtys6
6zPGa+6JLfAjJxT/V57EA0MvJPKhIvGUZ6+dK5y6vGFZ0dXIRIGxomUIuWWJ
CAbj5R3iNs/PSzRgtbzWMlkYjyvGYBfr4JM6D1C89I2ejgEV6ASAbZuCpDZB
EvJWzVfGm8GEwvKRN/520sUY1lxdRm4xfZWKW1ewCrWroEvvJk985vY+ROHL
M5mqnJIWVUrfHprxGWHdmP7tnaBi+ms5j4ZGc4ZyP3sWmZeaN5a6swDzuoqZ
m7C556L4zGjMTJQyK57djDjc80rzLgzD9k72v0mBjIKlMf8cAJZvPUqsp3wP
Ruz8A1hBnrBqUbNxrAHLt7t8IS2UcJCMJqSAA+DZ19aNYvGMan0QjiLZ9Ivc
tpJVdshDppb8eqCdrCrlqn2h+lpdK2Wzgt+vlSPoY/5ucgVsMury/ZJU8rlR
6vGiRkW4F7yQVwkSQk7bvlGXCp164wCpZMFVf9YZnFgQwgW1g5qwWNlsX4v+
qLMZPDfeAL2Ly1EPZBzswc/ZqVjdhj8h2ifsMgMT8OiV2kfyxYHlDmPX08QJ
BUUwEGIBMjbmNTqGQB/TWab4x5HqC7McnawAsc0u1KUPCJFiUZem7Z3+7OcL
Ajt9KDc4g9VKzwfzTEx+pmv2t1t67ZqR8J+7PeqlHXRT+OvlRcwY/5DNTUW3
WTSHt+gXYYVTqnSlLEho27kUHvAXhc6MQGW8UgZkrF9lc+QHsaOPnJ3f5yRx
c4u18RdUnRc3vDnDHE974nv2D7lYhJ/70QJ/qRobn1zgiVK5aBH4tR621AuV
3/HeKlSCkYlBAu+iO16u29ljEpHLkbWA9hYrI3TWzkN/en+vRdwib2d7o0g6
bAis8zAaFHeAwfy8AUqRb3wVHlFMBZN7l9lmwZWsZWnujJgAdZhzXfR/BN7w
aU9oBEAtm/Jmlfd0Dm4C7UOIMDIkmsw1lPrKB3RQIwSuv/uyDb6tjC/UjgWr
seM7vh5GJ68CVfzfBQ3AVM0tjJ9A8N798nL0Pn3mLfLauMg+WhY24naQbr65
Lnbevd8Y8A/pCm4zE1682h+MTGtnbUBj+IYWfJZXYGqKqnl3QNFtba7qo2aT
mZpMDm/MZLSr0wIto4Uu1m1Ktthctt7N1oZZLIDw5YFNHTDOz1gvw5YxHt1t
ah+WWfC6DjivcOtqG6NwrAIj64B6vL/lz1MJz/BfsuF0zbQ39sOkeq5u/hZp
5Q9eh44tSNrWm+rM3brS3mFsyNbnBrknYsll8W1HxqgH1eKtO07qqBgJqdhs
367kmnRU9VY9lyX2jMcJ88W9OQT7IwiaXea9EIIs9vD2+G6WkbNTQ8MFWra1
qUE8KU9TnInDeW3lVAUehqnMPF27ry297COzJ/NWwCyDuQxt3LmB2y4gFHGq
GjqFQg7IDy0swvQ8L5E2akxpL/42L3kqbaMZZstkb67m2rsEXiKW0nY92+7X
jZ5kIzTo8q6VT+Iva/vFb5T4PyvmWj70FD5GjD3gZvbRYqRuA3VXfbG8oYdv
9zEwagJkQwlUnDVpTXvyXoXzq0jNQhW5DSLqY47YWb3gLjet7OcR3gxeAo0/
wb0PM3X/nLFiLRofhWPwPFxgfcv6qysQ7yg5qv4/bWoPZ61Ws2uBo/XSoMWB
Mofh4JptS1WW+cCKcUy55gCSxaYNghrJPzJKXtJqfQrJHUvdWTYKOfyCK0up
atKmthcYkrdSqS07JEZ0bGgrHQK+viCggtvyArFCQVRAo0dMyezeltD62m8r
RCkvAbYt0h0aPi1Slz1lge5xZ1PuGaggJx6BS0c6WCDwTRKEtfjIrTYgeRgf
WdOXzLxTk36cz77Tg7pY9ka3Y09tB6+GfWY3B0wjqCRqhOXlCF0iiICpzMDR
81Ql6BjxhqCU8aIk5FB6j8DIOomkPToRAil6d3W2fGGCAMAMjXLv8w4/mfY9
wN3dOZ31CvaWJPoJs15P96MOqVX4PnlvPUYU+98qSvKvHZgZJyh38UVnk5x2
i4CuzTbKIP6EiP/eG4yy5cx7/QFNOE5KyRXhuOdxxZF0+741DBM79rYLZ+Gz
/w3U7mWDx/A92wuHU4kYoWqvTfQVh4g/1nNVp+eIKFwiwDJyBsL7JZeY8XIP
9QBj+ok//lHY7qMeCsnhkQbumiUqTIYFZJNSkq6tPywL/iYIoqpEyzZ0HF3t
n5JTTMczdA9iuienXtDehkAlKCpb9+4esVP7vNpjIvv7qqYJBtwVjM1D81Uo
7x29SDjWXzPqCJXUQsb9tO954oH0GhVU+wc2zaOXfAQx8jnHv7J56GXGqTWQ
gPf5mAYW8X3gexqLaP5kXdu0yck0WoYf/lmHYNwkh1wWOHJB47Epfe0huXaU
HjVaCWFVjmdDPYFmyXMmCSZVw4O/NxveoyczAxBTj+DqWiJpRdIHp0zE9194
RbsyDktLWTwsokjaT0EX7aQjLx+GBG4e4wFXpb6qZM/IPadm0cobmn3dORQ6
zGof/qqAIBRoPvlGOfPfES4w/Wyez6KiQM/2kIUtTNS473vC2mTurt5kyy/v
1pvgvvBGDEkKnE3nEEZoMfCW4XOSn1Zj4nGTXGLfcu+HNmg5K9vlTaVpBw4K
2ZS3oTfLj0OLeYiDWYz5ABrpMjdngQEJA0pDq2KCG//Kk/gg2XDFNDc6/HAY
TsWPuy1Rg2bFLGt53qmsIlbpv+pn66NMDo39U5qXs2UooVsr4S2F2fcrqvwq
RMMdx/cQRP9dBl5NENbqncIPerqWEz4WTMSs2ZnfdpTM9a84MThv0OemA9g+
jDve/FSkgtVcF3tHVQ8N5sTKJAB9+66cquaRX0F66HO+OPSMJoU6OQrnxsnW
hEQy8WzEEolQiDHGvm3ZlXOjYsVHJwM1zhauCrzNNDryJkVRa0GFuI7t1uft
v5/Isdb/dZpfP8aEwOXV1ShREVd2yuzfrEssiJjUaKxztZXu3KcZwPQ+HR/V
c1uyPUHO9YL8C9wKmeIPGcb5677tbbqCSXi5XQtWe+4BpsHRoU1DmuC5tFJ6
o5b+cZfKoKUJ4wTC+6yqXz+juYtlsnE5pq5Ykik55GjwRfzZM4hzc57gNgoc
9BOdCVpW8VCjYLHhUhagM8wNAcDTyhDYQwzHXx7OIgFXWUaZRXwhJboFK0LJ
k6SksbkOh81wKlwrlZh0Gkhkc6UMOdqDctYobL1wZ2daDWhePBOzYJeVWjWx
L/C2XYigXSo/n0XcnRcJDEK3tSIj+Nd60XYdlp6ADaPJbZuLoTxEjCxUNBJD
sQ7CbFPk1zLhjRFUH/F1Kx7tYzNH/jHew/QMkz3tt2rHaiHfq+zznyeeh+WU
JV/YMYFhxQba4teJ0XUrt6bhnbEmdgx2oPVKYxDbOCSP/AnEB7UvuopRKWHJ
ik28zzJcAG5USc00jp+2e1Qx8v1NPpBVKBTHeLvPeIbkRkjCaSqsYNJEr4Gn
bFBrhEjOuA8r71HR0VzV4tPeixNC8LHj37m7i4eAlQHdhh5U7nyNEhzrt5sr
7bEfjICpu0MX/2Vu2wJAusCZBTZ5g7BDLfGW2+hV3xxEY5rzjTO1XyUkRVHx
rmNDp4SEZ54oemgwNwH5MXjbgRdvHO+nHcP9kMF22w+P6LuyKgDcsvqvjj2y
S+nu07JNeYXpv14g9hRm6O4cZPFo7vcDDQb6Zn+6mE+8p4QKWbEkMc6+7b2l
LNFHAR5wOsydkLbKHOUtw1r0bc8jiODilh68cqciQKevxcTgOQqHkYfdBpd5
PYed2FKkF5GlWTt6qSpvQ/5bqb4Dcno2Yr4+sWTMnMve/IFx7pOiz/9LuSpu
w6FMJ+M+9qR1kEtEIzQ5bJFwtIJrJYHaI8GU6wx93Th67OrdpvsatJQ681Sa
RGWD2Yy94Bb7UsnSEJCxbMxKZdkmQjE+RvIU6+6Wq1omC7Gpwem2+AikE4RX
xkD7N+vdJhzR5iLfuwT4zekoNV6uq5J0DLGTPG8+HwHylhEJFu6KTRhoxR4B
XTa6M9btnPEC4CJnzBfj6cCrwjnd23dh+x9Qqh8oIyFSZAuYA3vQYKEu3+N6
BO/pRPoV/nfSc2X2TO340LBl0jY9ZeHhaLWDZXNDIsd75KoUFM48f4nmTdPe
PdN6agdBCr+sr9BSnJh8IqZYbYV3I1IL9s/DoGIoaXkq+fsuS1Ixd1NiOACy
ekwH8Z/qYpRnDMpIeeA67y8es/ufvE+ZQYHVc2RbArjezzqp1rEYG2KXv/K2
SxqDz9RsKaxtToR+hhEnqm8XH7DV6cCSfBWhrZd8QkSemk4DIUvLHmbEHaX0
8gzd64ggRx0tMJvdOU4/xsUwNZwdp3+D8foM65yO2wsau66S/RIfBMmvp3LH
LPUwC+vrOauNTzUVj4Jxnrt7h+/l9uRxLh68jeeKxNoqmvPBjZK4lIk7sceM
vZ8tnbu9h0moHIMy5T4486d7WYg6RP8fqaiWjpjXZn/g3wk1C+eo7+fcBI8u
61BIacckaPpaF8+oLCv5C0vqAwKncvSreMKiOIQaaQGKYO6AefS+cl5mwLuG
J3lLhABGMvHRhJ1fx2PJBND8C5Z+TnADyG3/8KBmyEIqzGC3gTTrsVzH+FGH
NXGh5bLpu1LDeduys60nlSqCWUgnpic6odgbS8FqJ35s9CjCqkCWMs6f7WKN
aMLYrMH83XWaCUQHNmbGH6rZZN54zlvTRFrw8ceX9Y2Zr8SRoWLzZ4wPfHC8
LHau+XnQfMuSS8XCMmRX8vOtDkOe08SF/a+8Lt6mVKpQyIvqvXyvTLThGaxC
KRlmo0JC6NkWLVdsQ2xrpxoQf1pb/C31Tq1WVLpwX23RYkQOlO3qqSar2b0R
7w6iLcGZeYCVtREjmzqjxDUMTR6LEUO+VaGJ6yPOGFx2eIZ0Hnznn2V7ZOTs
GofGEPHt+zL2cFSATl9UmIC+CgMO/UGL1VmpvQlJ0b/s0p2PU+CsXR6YezUq
egV07YC4U6bXYdiqPRioNi0iOzom4ZS0cPYiIvhKf8WWMgMo5NUzbWGfdS7a
0TPIYQXL2qqNbcu4J2qqF1eC3zV9RrrE4N82D1vq9936blDsnx4DErOVDCBy
GL1/Wokzbfz/W+hXXXAZRhIDpRkQDo1V1TLDEWlZoj6tyBMQycElCNiU3sDC
21y9xCukx1kdgvyun9UzeBlEFWwqiszZ3xw5nb3UE4Km+P9WuHLJg3uSdEeu
F5BmnsIr0tUIvFiMKhl4HZbECu1SbtjLumkEJ89OpwZWOE7P/qL1R9M1lvMe
Hpl/lUa6zs/6Iv8BbTuD/zOKQ+8y/twu4KoTdI2XCJCCrpPgKux9lvUclWhn
LczrubZQB2yU1XOGZxVZuTNkN5cuGKFTRvCAhWDvXsIVP75PjfgZ7RFSPxAh
hndoMvH7KI8Y947W3Y72b9e/Wf4BGmL542l+aVjjTKr9q0e2UGWaZoLFO06c
iIbfuvCT5RV50ipVM2COwH2d1DhGyKmM6gP7+a0WMa8q+p2SUVCWF5VWWNMd
PVX4ljQKb7o5JzW7AFJ3hbv13DSKXKkzNJehF0EEcPrhMcnjziRKjb6EBe2a
rDHtIgG7PYtaYxmJq5rTKQDx0Ktz4Zi6K7NOT6Nlr1wMMh/YsE5v841sc2jv
JgvXnIZVybLP79zXp01OO3S9Szy0uZav2VCssFbVA9dD1iTC87YbAoagCauV
/R683yfe8N7IDqrikHDvCEn1NE1v0UoNXpoPYMrOMZ/DrlcKyu2wAkvv4Ep9
QdfxY9UH8I2BIyunHbL9PXaE6lnE/pLyX7J0x28WycwxMdGMPO/U6/GVXwuv
3KHgm5cs5p42yUJ0SEiERR54o/9FLBqGyLm0nzcJf8IB3lxRRcE09AgiRp02
JUYu/5vannqpaPyj//nAOeStJ43Jmgi/MMltzxQY+PfITMc1pY6bLZd3/8AV
HOpfQvM4aNGcik+u+UKVLJJfD87PV2Tb65AwhfaJPE+67i+/PBOH+NNPP+5K
uDYG7/5tBdsU/4g++TKSvcrYYVbMITmFBhudqWB75t9cHEled+Yp4+WkyOnd
vB5f61WMBJmjmHGWeO09Vz/h+smaFBa5pg9qHRSntvuM1G2Gfj4ZhF6EYced
5GXKyODrMNjTPekXjlVcAqHqVEbLn0UDrwWa4BN9C97A15DoxbxV640XKuZH
fJwp0e0jh98/4w1PGoXu53IDpRu5rKoekwuHzXsxge7rKXUAU0A9VNz8nmNO
zVUZSxlUcZJouQHm84VPncMv789FARzZbc1dO5fLi/hxhsDUs4Q16kAlSlLC
bJQOL8h3OQDQ+9i+D465AWZswHyxu98yoLkAfTrBjDBe6O4SnZHxrEBZWfEh
5cY7uwwzWO6HfJWKuBUgwlo/QKi+n0v7l/W+Asq2G917Sagb2aL53KNm2txZ
jRLxTtZtT3FwTQRgJW1TDHi9TKDlS6tOggTw3qR4TJ/b7yA1hN+RE5ErV6Xq
yK1nqlCXyxryi0YRrlWBgDWH90PumcLwnhAojGKhLF+XfBInkyo9jOuu28IA
H8uoRYMek4jtD6Dc3vRJPUlXgYUCOSHKk4UYaYi2rjE621PhriwG/fokVbWa
x51YOR6poybqXy0yOM8FhpVNnJTPOor0khwjU6ihe72492w5zdl55xC+HJXV
OSFVzJVAEQDs5C108+kKUHpAgn2UdIxSOl2TOwFwimt0hHX0veDTn1mrtltu
kl66RXVS8Ihly59aWoLOsjF55hzV27vK7ORQEPtsduSgMzYo8+QkLR3FplS5
Z6vk/+SZKMOuQYq7pZojuGQRKgp96Ngd23AAtphjE3v0jDI+QkGPJuXZaLiG
72A0Q8zt57ybkwV+S/fXk9ASl18f2tYZCKVp1n9PalWqEskc3joD6LM63TLu
tjeUVjEbjoK6S+/8DI1RmWiNfAQ3AgazsQvI0hcJQ0mSU+X1VX2IM+FfS9fv
TYfAGW8a4yQ5t+fzvAnjvBQKl4pWhho7P5PKa0zNwVL6ayPC9r7oVZo3m1/f
OMlwadqfcyS4uc3EO16cMDtTvnimvqAbhwise5myL+9nAYmUz16VQAotvVR9
h1jSNvZKTCa2DQcM+cMe645mEzl5SYNgx6rRoFttGeU0lbzIHg8LmdL05v5b
aFSp93LuLrRH5hr2pLhI1/MdacyXB9NvJBHMfEQlUfcfbxAAxMb6sp3QOjba
l75o7JxFfkGOPwojJXwmlf999lk0Eb1y1wvkPc59eXQF5xUO3yi4VR65wi/y
cJM7gyaKc01EMRA852o0QabTBZwsuYKlx0+RFJEsWr9qlOiSqWiSg4JqXYaB
qYFOI1TstZfzEDDOvzubQLWEY2vDLL1fxt4S/CpK7+ZCaMDsCY/nZjeteOoc
jiELsEKT5q76/x7/6Beo/jxSTcPV9K3OP+qYMhvHE3TKNC/Tltc1Ewysvz9a
R6TVNzgyytiuEwuOj+h9MXU1ToqJWJZhx+IIpj/7j0B///201CVMXbSc+zoG
9fsFGTHF6fj+ALZZ5AqBrep6cSnODrmKgTqa4zgaeL+hwq4Um9ciJv8zYDI9
sSwvyLYV2cbrv6qXmlKB1y1k4BP/fHq88Au1FhEFsvNNRP/oavmhxJ4Af/UT
xncAFadWt+N/utNkkY9n2eDMCxdBbo6g1Jb1c96p6gOhPWFFP7a9+qFZ9TrB
jB0ArBbayBPwdf39xzewA/PJvfnrOaI2weiN6T17f8E/IIE4/LhOxko+wPm6
3lBecsU4OV9/YOsGWm0uvHmPH6dH1QZw5wUGUjbg4BsR4zXO5M8q0KAsbOla
lWnPc4HHnAZTlMMD185iTMI/i6Z+ea1FgTWV5ohQl4jsRFX9PUIF5X/7ttQu
or+Agl9Ts7otujD1KNIdIRBV28PidHVXJ8+TeIMgAF/kud2mgUNG9qBD9LvF
il36JQFvWfhwtorcL0gI8kpJsJWsYj+ESJXpOG2y68RePEMIvr7hw4ww7o3B
2AeVlFBhlbS/FVZhzi1gj3+0xuCg5yxsR9jWJ+FwydgBNmSCtLFlzMVFMQM+
AJ0uV9tXMza1gqscf7xFFbVxKC6/veiPXAJEssMRo4xm1G+rxCBQwJ5JzvGu
F/W4yz7Do/pW7yJSNdl1104E0OpB7b0olXPZVE0TBcfiEmvafknJfPBr16lO
yLw4YWNGnl2FF6FoOIOXLAKsw4ClYLQshKhuqdwT7LxRfnToRnVXjrP8U6ji
YX/NsyvvorU599sXJmmgQvpjo5vTUmaJT//vNlvF8Kne039kagtHpGHSC+w4
28tVDJ0NcX1XK4RiU+GbfoG3e7aAPWaJehlxqA34XEltwH2ZEO6vaO7RBLEn
zBe0LUlgWP4YKDleARrF32Z1qzvnvTkvDvqWUdzxvhuUFQg1jIYyQeezovMv
d4mAvsuCVwFD1drztsC9JEXwhgC05i4iBEqprwHC2B1eNoEe+iKhaJSZn1aY
oaLMVAPze3XHX8FbZ3Wb96NDZkBSn1KMaBOH5X4nQXx3+R2B+WW29i9DfosX
GFNZh9WwBYWlSEgMI+McQt5on8pgIbtaZ8SLs8GfgPmNAT6qMK5aV/+6zd2A
Z6xsgbdafkzbT52aSvauS0Ln23rvsFTdb9wmW3mRJvkMPFY2xr1uWC3yr/xw
6gpUo4VzuJVP+935mIh51djirThoK0S2QVvfrXz2XIPznEXy8ZqQMV/lHpEX
swP7hqnyNagm9BqpTy+LZ0cBwtSldUqXDoHX9ecf1gB+2xAc2jLn6kKLAiGZ
zUHigSZUYJj0k2MmSNGy0Cc8+eQeIfT21YtUqRfHjZxVUFZWLdZfiT67wivm
PaXJmShjIL/A3y/wzyz/QBJyGfXaPpvkZKJpKqkdnzQFAhHNaHwMNoxsswZn
EyTf5muK87KjUq07CS/678ts0DM+J4wBDFFLVbMsrD73QlaHhcWfElMUyPhy
XvF+UPPyXDXgMmF7h6EUuY6P+KdW4zCaB+1xcJ7aLTvzVUDtfWT2g8g+oEmb
+5j3dC4cyZy+G/vdN1t6hrGf8sK8xphUrZUsv5GgRoAbaGREAnaXRdC8TFxL
U73OsbkFlszHXsSrs3Fe8oX8Jpr5MQlWB1nf0RMTT53Pn9Exf5FpnsduZvx8
WlwvHNryqGz7XWzn3zP1Uvqf3IAeOZq3T3H8atSw8mXcK7yYt+O23U98yO2m
4RJ4x2UhTEnuBL1TWsg/tjGeKmng35PSO71WzYrT0Pu3mhVyNd7DqlSuUymd
CSBP9ayPFM6HaiXkJP6s3WYPXh2gWXLNRe4tT5PJsA7zVzy1AOzRdNnxhZTB
dJ1O8dzYuM5oghoyYTZz60BQbV2sAoM7Xe2bvHBHXUIwmmKDMNKsO1yQ5PAP
RcRVwsN0gfPJBLyADePLH9lb2wGHzyTfjDEZNPndezhnxrpEoQ50ySUfZb1s
prVQnRAxJvqnDJGTXLNE87H5zNgrRLg2MuDj4+HccT5qiX1ePo0KynKa92AG
qdfuurHBr5ZX3D3T5WWugM6FHV7/qRS0yY7PbIOUo8+ys2YwJy3Toe7R6MlS
UzyCl8t2U4O+u+H9vO+eaOPh60Dop7pJBL1abAuQYwSv0PL9QwHxtXsv1KMX
di7wi8vpLdC9epwuoXAIu9W2ttLYho+ti6uv2PKc5QN2DhL7DWvBCqfIKE5x
mXNscCdE5T7M+bXohIp04IejCqJazeFVA0SW560DctMqHJl6QXFODqqHXbPH
gnuvmoST84ocrvr4uS09UkcWdkiRefA9336OK+7DrdkxUTgAhwOCyxG1OU4C
/yJ4nQdVcNnu4QkOcHnUBIMRWOIUEUuPYq5PQgHUsDta1j1lXiZWMj/wj0Jt
wgKLgQIrJ8n12dIT4QdKeb0gSEwrfa0JNBdUAHMBHCxo9462x8Do2b5z/UP3
Sk9NCgXx2p3w4VKSBC6//d+ZnBstFYA5x5ldwSIKDSe5gAb377fmZ15BToOZ
/DqMuMVxl2wTTZA3BByV9BoaoLCn6wYKUWywFOT+lDsOrRDC6BfhYuAMwEOI
F8SYKcZhb+/e0vh8i6xhrMAlUVvXg793oXB08s9Ic3fJ+enChIqN4jHOXXWB
FWK4/Qoe0a3c8fOpoWyclwpfoiCNPWOui7lfXnqM6ZIOyuEsiOc/woTA63df
5n+6gOHreoXGiztCVVDaAi49Hr685/Ak0hEwLilyZQeua7lkqxlZ0QP2N1eE
gQdo8WAh403Rz294DK50djwqPfBeTKEyiOOHxxqtrbXY23B3O4G2ndA2um9O
DVR0t829BXiR/dj204rQM3bY1R9FQ9ZYcJhijwOJ736mbUYA52t5khp2s7/o
sj1LoPG5Xho93RpWAlsy/EyAgkzEeHp7dSV+IUTHavEh4G5Tj26bxbZsxYRo
WQB8Xm6i1vEoeY7LXxq1RrsMJiIMT4w4vDBxXae9RdJHWw3BOLLArJ2Al996
PiKixpqEpbTS4nPnxh99iS4UBPOIeJnCs6EJb5ddAbx4S5uDYNLbb6SR+tsW
SuB6GOohHA/0m8KnYLj1bvY3l5VezkHWgkAbCfE4K7PNjfzE+BK2xaE9hZEt
klsuEc0xNyhkzB4zYQyOAWE3SJnlxYexxoZXnGDJNLiAFJS+MlSeNx8jI9JI
8OpYg+njNtcuuq9ICI0RuzhmlFlg2xAXpo67Uv4Gje1BQ0ZfcghmCPPXUVdU
GpeK7NC2N00iZBe7hLoME/FiQou1dsA2PzhDoDVWTDnAYHJ2VJXv2USqkHkD
j/ABkKs0r3JHb6gfFg9Uy8RU2N6gWFSq5C2wrVrwJwj43aoCOGFQZIPshZKS
S1dQ8u1j94Z8jD1rKKSQFkfrmlzEvD1UfQpDlx8dWdokPZ7Bjcow7w8FqJiY
LKsP2B5uk4cjXEkH3ATIDNW6MviO4DlJppxUJZBQo80uUxvFIluf7gYCqdgl
LA/PscbImU4voasgn1cUocrn6UNbHDZ7dXbrrzP77j0mmzM8ATM/k8NnYEL1
BYamVpfi+n8ns23SFKxUnhbS6NHE/EBzNj/Tw5CkRpQsC9cg4w4QXpAn2Q4b
XbM+aJ33EKwvYX80OiRN4x65OjVinkfVvQUC/bsMjNM2EMxM1z8T48NlZGRU
R/opOxbnM0VTZqfX7hqjK3D6ZeSXGhnvV1d9OmCtB8p1Z481OTy01GUH435r
IK70k7v2P8zPu+8O7r2t2d7olBk0v8W6FE/p4CxUxHUDKClIDyBRVoUxNLg4
ztaWUtypyBA3LPDcPQPk8ehsAWCluHScCHzMvKIYwnP9gb3iWe+0uiAtJ4du
tVmjOMDCRRZU+N0xXBCTNS+sxFjrCJhoRFKTI+wZT13FFxUX949qxNgko+zc
5cz4cp0Z+RkCHGw26t0bo6lTewi+Y6mcU0rEz1YF7Pse4rFbxwj6xVf0rl+2
J3CKLc+lzBXylD74B/DywcpC4SpADykSuefKmpqI0vXYiWxPhjo4omp7qZte
DmIRVcBAtPcFG6mGqLu9not5pGi4jgZvX6WRm8hr8k+wsmDWOt2rYWmJ0i3B
lXgoN5ZLMpArIwUyudXMm8GivbDrLn8mgfTMNGT82JXlId7GmK3rTmst0xd3
1hj9fM3UGCSlOtE7HLnqvULTcV6BK6b/S08KVp6OSTAtku02Bsa8iByzeqoy
QtJGOoeiLAXXqZyKVYmzVRtdtskV99TtgloNLWNyRK0+WG62/pUm169xC6xB
k5ejW6R04Z9QsnyQnyJ20hR6NfehyKYcRCPXBjSvtXxQ86RhL51eoceak+Tk
HeyA2X5kMB/Iur5IkCaVgWxuE/Nt+I0rZ6sRRFyu0jLN4Y+TaMw9TLTtKbvW
ngnWPwHm56UuRZirYTf836Mc7AFj5dbH6PBym0WChKxaKVgjZR0HA/dT9JZR
os1nauybzXpVPfd/WXP4SyFpF2Hh8HAJrHj6GZd9/w7Sa3oGOqExyY/x9fET
OBnlV4jvxS/rZRL3CHZaPQfs63Rq+S7dB5bn1dmol8ojvJOR+OQxKD82aH6G
ZbWwGgouZBunclE5f/KkbwZmaI6QwHwzEdBlKRemn9tRAp6AMhWCBLfF8JFD
xQ5dT/Sr7Ulwx/by5LzWEJyp9YoU4GtlUEZqQGMdNxUvcIRSor4NK/9ZAfgn
cusTphIg9WQG9yTW4XVRvxRAAd+4PgueEzNZ7UossCmct41IqVhSTWi5RMQw
ufXMZ9fhq5iI8itJMWuja6jtEIInIfIAabhTdcGuWEG8jsmZd2NcT+Q0IBL9
H0gtWgNwCLT2xUIQYbLxx7BjxA+4tjygvNGCcFNhy1MgvfScVcZ5oWvrNZhq
NLnNGnxg26jeezExlr1bThIHqWR+0l+QA/y2yOIryFlegRSux+49fML+A/VP
za38UKtMP94tEXWQkHWx4AjpEZlOmv71uP49ldg1RRJAhVZSjt5fd8s/GGFB
Oy459m8vJjUUIbyOdtILiRv/FY9egWS57S2d/41X3V3QkBnxABRvqXro5UTB
qfF8WGxT2Rh/PrU1B/j6RaUWnfLi3JyKOBNYxQfEB7UBE8mmd1ylmZE+kSnr
hhOHtdIJfO352nv+Hhks44D8g04Ct/6TFW7Os4Migtd6VWj9Bb/LNDUi6Xt2
Nl/FAB7JrpadLzcPq/ayYd5rORYN1khrjJ3IfHzqVvY3iwcmp2/iv1gY3sGK
gEOTWGziFHffOYdjFddzos/lyjXgOWVYRtmjIATGy08eG/cBsafJbyiqLh43
OcKvmcxQ7GrPH41Vo0u3eAv4ohaAemNAWxgn2Jxhax2Myp92V1HIW66HqULG
bTJLhqDlaQ8sFX6G9hgrZn8b1ADcKDcrC5qKBgPfQTxfTT6oYP3fSbDnU3fs
C0t3WI+dHa5DPpyCFKctV/Bm0bnx5wcJwRkGp1s6y5pPYe1KbEWmc/iNDeOM
HgG68VKHGVjAOAiXjIp0ahv0XyV/zcb8fEixz4m1dZE5xNU8eo2vgIyywSaD
KkzaFU+EG+SfJOrhdgaxDbt5vjXUAZ8mfoATN7prAOprF01RZDuPBMFLZmUY
pxLwWnHtRqe1nMduzcbpSCPn1nekGezIXc5rTVl8Nh4dOEGrfGsYS1wNU2M6
tC6fFPydtunhtzShlxB9fZK4cqpScI45E9rbPWG2tcaNs+KT8y10MeAWs9iw
p3qAHQEHNKuKoNHxlJDFNmUCE6HZo+f+5lZf9f3dkoE4H98CNQG7Ff1zzgTE
s3mlVj3UkRHk+HMRrtiMtZzSg4MgYESHlgYQmaIVGulbUP06EQ06SaeIzXNo
Ct47rcteWawX6dggYrvgUQ4A3GxpFUN5vEe7eg4mrRm80vf36jfx48utAFFi
2oqj+RIc7aBWLYP+AlA6Wh3rj8qgIKY22ztaB+X3biIgShAKk+yhjpmfVcOD
CMLF3rphdfGsjtpF/2WSTvrEzeOOR5DyP9a1I7fnmJYax41JvQQenMXOqFVw
YB9ycfBP4kJupRp/LpXO2TiD8QCMspueXBg0VxQI9JlIa/ycCaFbsLHpyjAr
gd8BtNxXOV6V9XdKgj4kXfB3C14GJWcUaMnl2DoKyHefjwmrwOy3Wdopvntc
1JHX7l9EsLysmy2gbePHyed8FwwDkyT2Ksv8o51A134BCF38t88P5raItZxO
U5TSScnyLEsEALOK9uMgWp8kzInRwDBYRkT0lAtWainamUpIbmqo1E6DgSDD
IL1F1MwKb9xWJr1x2gdtvXnhZjnmxeJj1JIsHECH9q75JoK6du80+vugvUUp
3q5r0N+2Xm9Ayisw59ny99BjSh2CakBAcVj6IIBBUPAIvJ7VGl5ZUEex9gQO
0LVnzB2zvi29/gNTFvVPzxYOSyILxFT8YM5MiWwTZswO3H8U4zB47/RtVGUa
P6mu4XHl32RcRVW041sE11iCAdDdLHfEH+d/Q8PzwjUWjXy6N4MtZln0JA+a
9bWDLzrNADAbVEuImZbNziwV4uVsViUE4PAP0OMgfT85lPccbmcCI56UkrBJ
hcG2hbLODNEkibTKJp7BM5NVmINWXUtxovBHVglAKQtx9yj2TyisconzWJzn
pL8mpL5D+8ZirOXVg3+jSv0OJLZU/JGtylWib0NvZn/s07drSmUY94hL/+UR
t/9BQ18OHYCSJzJdBwx7T+vlUUXvAXk+a2sggpnh++iaXdA7L14Zq9Xil1z+
Z5sARrUV/XFnjEhWMINebLdNCSa2BKNxc9HCF2IxSFgqI25oZr9SODve/US3
Vp2YLBvNCiEE5S17pLy8+II4TXqgFUDNdusYnY0W42sPyNDhKYgxq/FgOnWF
kdvfumXfd2PHsQK2gRxrmlnZe0pDBywQ3wvSIA5Pj7Rf8gKu0I95UAkQpm7T
8FLTdq6dDdCFUepa4XdnE3Ea34dpSwaGkZW39mnCKeuMy6J6kUtQiPdxHWl/
K/Ztw+FNDwN6tJjh5/5QJwnbxxvXQFZ1P7crb8vS6cWd1R2Jlhitaj9aYXn2
fwqu0aOy8HOJY/iR9jlfyLRqxmL6EBPQkBF2wAp/hrV+GZT5Dxo0pk5Za9Iv
vGPIhJVX+HQAh781BeVw5nUxHCVct/BKc7VxCaA4w1AyO+ocqQdoxJaHAchy
zbSQZ+C2vtf3fByFmrH8rhQZ7+QQ0sb2DIsUdP/jVs0lVJ0fKpNDCAeDnNzM
ZGB0KAZ8jk9/zruMSf0yJFOINYySkRTk3ehVzodd6CcgPefHl1Hi6TXrhFVO
NB8UTvpfMk9hhGiGSFdo8II0xOQezqqQuAT/i+KCsCwovRy0Fz5dDWTtEZbj
HOytyw3hX5pdUp7Qd1cnDqSy+L+uD3YkbF1phIcJvjBMtVGwX9s0V+Ync+lL
CM7QdH82d+rNBZ4i7T6PbpFQYrPiOtMJ3QgtFr2Ymwm60zIMN7+K210MgeB4
fRiQd8exPW3qOTdvFotRK0Pqv7nXz0aTR2tOcmtIdUq6TzJqalfh3A1F1QQp
U0A8bEZMyJoc2OnFJdf+2AcoN6nGDSfzdXThqacw0eCsq+1D45TuZxomRSMV
dR33bCyjao/xz2gAYA5WuxpuVDbFnTKuR43eri5Ih1VQcUuP/XFT4o4vplwk
Aj3oi645RjNyrIV4YtY1fx74WG3GtfAWBYD/ND65FIsWz+0JMPDiroXDtENw
vbWnmbim4anhq1FZNM2B00tMxoLNkNWYuy3IQ6jo8T8P5GVDaYTM3eLELVcZ
//xMfMmhYY/JGXDghR8xVU4Gc1inKILD6jf8D7y6DAfrjzqajwqEqNJrXgLQ
vA3VHICK+rG+mAbPqD6dbcWAmbOltxwEbdueyFTa96j5IBsw5KMqnnkv52nd
tWH3Ou6OBOl0HJMGHuxaP/6WPk2vmWD9IHMTrVkdITZueQfVf0XLfXD2/UpA
PjT8OeiQYh6N0cBza9SQKGsS9nPFaZLGBXtUcZ5Vjez9t9YMFccVrGKg1GXL
NO9jAESrL1yWR+fwuPTKbPwQCdAAwzpsdt0xocr1/Lr5f5kykMi68lnXYcjE
IRKn38sK5yymtjbrSCruY1lUTxRKs10raWAmh8HbqHWTWkVMzrXLl+1SM2QP
TJTkcIznuFyfzhEoFt4DM8zzEyzIlwLVoty3xMTMLoi2rBYSHroA/Ev6f9B5
rj1RCUe5HMUJLdoiNiPCuM9ZjBNgHx8ds+yoeQ3Ls1JCq/Sd/7wh/v2o0YJ1
MhuDjkVEr5kbcOV72Yd6Sf6xT5vhdQptcmdRGg+SEyTZ0NqwuTsKnJYjRcXN
ZK8KoP0KTosVxr0dm5W0EucUV9jl8m/7bNOI1w7ow6hOIurP1vHU+tiwKQ7z
yW1OX9fE7+aNgLMOHLrOndqg/UsHJnDaSkm0RzyY9min2iqWALyy6oxmKqo1
odh71n3DouMtHIFxTrkbVZ9vfE2mhOzlc+C4gyJTqDrJa5CBiqWm+zj8kJhR
dM5/xkJ+6Ml7sI6I3ScwupqOZlD1cPIDLIqr3hd2YS+sx+ioaqbQdOvKogT5
V1CyOFbvsLCpJVOY7KwK2XC0Y4ZIVitv2Zlc5g/10HMuCiE5Rvdnzqu8kksn
Q7KoaQOnqIl1L6MtIhrw28zHsuaxOF4Mnql6oP1cXBkVG4AAI/J7cx0aZDxq
LWmBcoltwmahSdHC0i+56eAyK5ESANL5fCHWIWJOLlmej3mow33NkyYn+9Wl
nZ+tpcWO0kSSU+U4tzAOeK3aOsD2Ey2wSsMlCK+WVWnIJYmNsiayFwOZOecs
H0alc9J1QDcm+OJ1pFLi/U5TrK2wDfHqlzEPKp9sa53wvK4JAgC4STa6qLsB
nNausaIsl8kAbQi9Ul0ghbyiBd8xqGNJMazNIFbeA5IMI5qszIL9N108wZYs
gMKYslM0s8Ry2QskLW7p9B6WMjPeRh8NX2TvGsSQFcibGwzRS8jrvr9FC76K
aFfBHSS5UiqdtkAnSXJB0TksknaLu9V+5Y3VxPGXx0qN+fV55eGhBa1SncI9
bFATPkBBKobMBxx6ovxaaMp4r+Zb3cArehVWTxuNziJ27dA9F29hSnjBzmvA
Xz9025eG43F/LCvGn9LDYkS699TRmAUdII2GAEOB/TCSPO+PfEtOTc/DVA9h
M4FseteD8nLbkJEZ04jmhdHBnD1w5GdqxsgFxGdIX7HtzwSkIUhfT2VHEICJ
asTWtRKnwT+/WM1Va0Ov4GQkumyKksSg02vDg2qn8agH3d2SOMTLKnxy9ZNO
SsSf0XV2PbiL5SwyQo9GXdLBrXp3p11Q4aivDNNNuVQ1oDdZQs8yr1j8d4Ol
VNDsAY4oiocAwLUufq7Ci1a8iun5e25F2srpxfPvGRbDCj/RyK57hQD4Ylb1
Zzhh9pnVYTctktdJNaRvL5Z9T7mHeziTx2Out4ANQCPkFycx2LtWYqJZ8g1Q
ojuMgGvoKq9eNy8iN0m8vygMbZ9WNiBaKr+IzKdDhzLQAdCr/V8DRc4PgJlw
+p3pepFcVG6Y0cnogZ/qXmbIuePbenH7Cae3kEMVB5+w1VubnIlKk8NdYj7L
2o8hG7rmJSe8Uxk9yVBqaMHUSEVAOTN3tD9aYQ7i7GpiKU34pFiDj9K5jHF0
hglCdD465pRbyBCM0Cf1JnLw62CtRUxpAu5FVwGo8nBkrU8/B4ZuoC90Y4Mp
VzalPOSa0HkTtBzJp2aLfx1HCKYtTFpoquLdjaBF0FpKvwLmKuIPxAWGR5nt
tbZIQkKZADfZziKfzg3boqhVKDiKYo1Y+p4UoGwC7kjT/1whQVLGfrNVbNdl
K/VlUS3do3RjKw0XKNh+qR7kw5cg79k4XD3zPpuRcN07stfVNVzKWa+Y/3qZ
hzBbRBWJTGYc4kOZ2r74xxVt5KTyIgTeUGU0UTA8DhX6y/5eUguZeUgvk3FS
8F/TNrZ3Dex5cgaCrDBdjcEnf29FkPvoCsv4JxaQD4Fv0pQIUc8LtPNhN5bJ
DnMcuiu8gSpB6qa56EuzyUd+Zgm/wEKSmO7Tb4maD5Zt4gNdkZ0WUAKphIFI
p1iEfpPPK8QrVGHlOxk+paaq5a+5/VRzZd2ZF/cK8O+3+pVRBDZnbZxbAGFI
sCkkkDB6/NZt7djQWYB7jwIDhWFR3OflzBvM5v5d37KfnPYIb6fxQgcnScae
mrWQk/+rd3ZDVBTBcGqe56LTeq1NZnlwSpqAO8bs4Lsjhgxj6ktOeZjs/QSg
5HWOgsyrZpha8IRsIg6+REOHKOHoSdv3k9LjP/HvS+vUOOuZCPGCxXyjrwt5
eJLKU6p5pLMH/edLvspi2cHTTwBQThRTLJy/LdopUiF44KKl+4Pkvvn724OX
aQMJuPQTs9TtelB8HTWlq0AjCTZJpMp9nmrIttrRrf/qEOHK2oksqTmycIwm
RBQpd4HmCoSjwJETvuLlySQzHuRjzI2hJfTxKfqObSCuZBxVJpjR8bKKHoOw
KQrA9P25iTcKCsmWbyCTkHcFWr/ug56zsccmY7dew0/mTUSEVjtLIeOhZzsK
YygrI3SwGk8dLDzA0VOYnw/RY0GYZkNvwB4EzBC2zLvN2X1uljNdRQQJQOyH
1ao2Z0YtbscwLbqduQmnoPRYT4QLBJ97HAMCWKyPcEU+JclrTGQ8l3k+vzZM
vC5W8u4g9WV0BEGjmEze6H9AtKFWA41AMVXlejqQbUOIZ0J87SuhWBPjypXo
MtGxGliuMSnETqXju9WZ1YMYuHMPoUXRcZsSZl3bYnd16GnSzdhJQoREeUza
sGGVMFM0YakbrglnONeFM1MBRTfkxSMrH/0KK1zCaZ02xP8veoGYeM0DpgXl
AC7Y9RHmknSSmHXGpyw0OEbC5nXluS0+QCioJyN8/hQIl0CbxtoofnMcKeVZ
jZVrSBNm3LTj2C8Y2UgJ/oWxotkPMpiIH7ly0fIcmtl3eBdj6m7Iv3wF0YD2
BkVqlLUkUoMIxGy0BBLm7VApLxeVVFM/Jpet6QoOu3D2C1kZR3S9Mr2GviRN
JKXeG0RKaxvevAGUNJLvB/rjASxgfx6fO9ChPCIAxUhJmC02cETI65cRyCok
TMy4anssLGk2PeiALTlqlnoI9KjkUqa/MXwBTv+MDybjevXz0nRkZtrgnLen
M1Qr+P/BNaqjPLLpnr2ub+iOJSPuCh63c55F3Ed5bOquxFB24fRVBhDSnMoR
uUnL5J2pllcgpl9Oap8KOrK9KlbRuM4a0ifD7SbKkIQ19unyIn4BdMjGE5Mf
QdklT1sI/rb9Kd/Rr4N3ttzpqTxrGtaIBe2pjhkgR751pJ6ug9/WnfzMEMjO
4dEPNdDH+uRKJoq9dKg+nHQpnk5k5+fQ7wi9QtRsPwz5rtxgwNAYqVCFmHRX
55H0Xp5CDIo7qZVPAMNFP1/FPZsG+BzLXHFVua5B3X4mYykGG5eJm9zXZJBQ
jmCnqgsxbmbxmVn/kpwetyl0Qw3KJ2FB9Y8yxylqfLOvIOTZhRnedsaMhWas
vojkINsBdxYE9gFLxQULpZHNaauaxNANKQ1GLy2RedKOFSYEimoc/WtPZUK6
HU5ZIfMOa6AyetiJcQ01bRL4EwP4eYEvvc/cbZnwaabXC5U76qpijPHlfafB
IcxV9MMKOcKDEiamVqSHdPj6t8lQg0Q9Bm431ED62FEkUZWJCb3Ux8sI+5UQ
0W0nbXF/P4/VetLoWAr5DdpXoEvkGLx1mePBGZPnYB8E+cI3YSGGNoif9gxB
aW2coocv9xgtgH2XDVVqAKUR8aZHHBPNsM0ooF7dLjrlS5MAK7juQFZQWzWr
vc9LBeoPz9VhhB43K/qZNjKi2xYdKr3D691Z0eOE4W7iAH0oLjp2tRwLm7Wy
SQ6cS9+pvOaW9ECeW/4Tb5QzTKDqbVWC86efotDXEU+deB/UpAqn6kh9hmDK
n7Pkx7JZuzykQgOlE38b6feyZUt1oEgYIpe1MlypOBoKfWZjXKm6yWiXg5OP
wxge70LaHct9eGbHpT7EyRSn/+RXdY6X20M4Oq6a/1+seyaJCsP4fyMt5woa
YdXR8qXlRHS8jF6nzBtElZr+TWnRWtWn2Jp9v3sCCULDtKwtKRIiyaXq2mWr
qLixHPblvVAoadjpHG2izjni4i+Fkls3vcEIy+mltoSMq7HcS/TETiaflV4w
sx/11EUEwwhetKm9td/Vrg+74uEDbjvBTXoh7I715afkTiLl38jS8cHyLlu8
ZgipgqWxgvgKYG/ywio2RXF7fvn2voZJJT/BVEYNXz9Tk2s+1Jl4qgZhSJ7N
3vViQjtXGbkMhXgERuzpiUDjGGPy8AKl2qME/HctO95lH594es3FAn0DoR2w
BKmRQXs6G1/9niFN/FSYX9qrutID/oDyglT+zfP0hZLp1NkdKcTRSkOSpbgc
749HTS3cr6kJfmlszdSz330J5ehTqF7y5cchK//4WtaZyu0zTWe3lm29pD50
2eZJ9RYZyrRAVR1bQR9tNl5F8mkt2rdb3TikCiHk/Zgv1lL0kJsa3QhPb1k3
jhtaqEPAC2azAKa1hhZgWD+63bN9nhSoacozyVfi6jj6pm2B7nlIgBDGO6Gk
xTzEsmCQ37Y+XG8D++eSX+8VHedK1W2ogNtS8fKto6o+h/Ng7+QtBRksLL5j
HFkVORU/+V1FNkP5PakqEn4fcgcIR2e25Q75GbqxotPGxyZgvUCqsNfY3y3m
uyUk0ILwdO2P2BDKtnkwstp9N4qHQ06EpISmbbIHubM9N1o8JGdwRm+HC2Gf
t/YdQ6TqW/yn0fq06MCb0aDK9onKfkDLKzisOZ/LMx6oqv5d9t0xfk3mcZnw
Xbe4+Y8CDz/SUESvpwf0kP9dUx+yri0Z3quAVKeccp3oqpLrzXeGlzWYiWD2
DVc1vO5sf+tlmBFgiHP7xdkzPhgixCRlsDFy95g1FZTh3cxBFCXcBFEIM0uP
M5CY5ZMXeWiPpnrNPZCiJrpOirg4R8Wyza2XbLTCaxEoGyl34WMC7CR25kOt
5SQ52Vc/CTKqIF3tWE5ynw/b+STsKXRqIJTF2SIBIcfysc6u7UObv4kjMoMx
Hg4Pm5WoYng0R7v2KLZxQEBRkG8cJQUpEIwFzsQwdeMUmGp0TKgxwX1CJKPl
/x68a0x54VR0medrhK7yPhLq6StkysnNwr0a+c5hODQ1WSaTzjQzO1vgVVNC
xxUminyxgrdMTRnVOzEjoTd+B7Vw0waaU3L6oEt9DQ7OPJRY1exBuqbztp3Z
D4FqMOZ4QdbdNlSig5WpDEwSTHrvcPJCzVg0NgJ8fMjCQ7X/X+wp7jHEl9j+
nLZ/USNyXh3jokUmimUmpGSqQWdy0KKHB1tgootM/blh5USQAwqpJRM7W+Ql
7R+l+EdbLtL1VRkMfCHzNVYpr2bdxTGeEDHyfPr+EQbavEnt+FViet6zIKTR
aMbrlL4XXHKxIZZ0LUxcoMk9VlyflAk5AQ76rvpdnU5RjzhxPRcujCwO/aib
7NtJfB2+cIdbRPIZAlabLugkK+MdaxZAtV+v458TMS9bFYa/LB9WOZ7SKOn4
Rn9znLpDF9UvcF7IxfA3VJ46YcCsEADj6YIVXwaq3dFUe7NaHHm4kK2Utdk2
3xOjJOv2Y/9GvYDks8knCJjr2/2Q70r9rVPu8sxIdE3wTzzTbSu3idUZPuw8
02NEy/1/gSyX3Xmd20eU7vFcLd2r5bN2YIZP5PpOLFwaPH1CJcLyskqdJ9pg
+/WCDp4Czp2l/8vLFe2NxMSjQ5b3SDM6dNIDmtulAHQwovzvKemPRbRhQqQE
HWRwhlxHASAD1EhIuh7Fq1xORC0tqHuCfBIHXwgOEjQCl1LZBSn+FpUO6BMG
ptwcB8Yi9j/hi/rHgJsCYrTORkpccswUyuCbWxpoz2s1FWC0Pod0bR5LRpIP
0n5a9mgUB52fCr8rIPrnheTRbc0jbQPmJIiwkQVjsIJAa1Mflb7vKK/9xF4j
3EBkU/YNhatzeloqWm8BQariADMNsdhiDiElh1RdxqS2t3g7ki1C7dMNgoli
XTsSZBbFq9Y42DboJ6U1DzSS3G9eW4M7Y62smqH5K9vwveowaYBjzLVRbwfj
lxxoDUgVUhBK9jiHUzLTcqbPpX7/MKQ46L/gHwv0JeJ93dGIaqfP1lzetfdB
Dqkw1YfwBXF/lLNiVEtW4wzfpjUR/0hsb6+zP90ima8vsbeyJeS31qsySNaI
NRBXxtCwni8IMkYB41re3DGGEGn07mGyxLRMHakXbiYYqYNgvTUjD0BEIA1K
DqrhbFdn+QFT35sFfRKjtf79/xO2dAVHN+WfwggDmCiHSh+8KtXmTD9ip1/2
8qYBRjwDSCXBr+aC4mhdEiwIG6D/VvYKdxCcIjC24lZpjTUw8qViLPxRKW4s
PN/13FAPLVJFIn+ZBfYkJlvhMotzu+i9gHQBEV1Z/NqF1abq8VfxliV1vDH5
HRsqYGBUdLSzxZLsQK3kadlbd3osJdkxtGKWpwF9X0kx+n53vjxlJz6yZrnh
PUdhb1fNY8/0w/dydAVXhu/Qz++vUUO5nFJ2QpPwV8HzGHNMhqT/ylDixvuw
WaNQeqF1IEbxbRP/DFWcbIcoXRC2eXKaZ+cWO7Jp8uf/3Qy58Y6Dvqd3o3A3
2lEtekIinH2qq2W/sYcK9cH16AobKaoU4JUVJLGPPdKi85CKP6a96S0zHcrq
BZE1Aw+/qTMe69YBYtoiKftihqtrRSYocYogzskrf76s1IRMhnM11bscbqNW
U9M0fMDt1S9pzFjT2lbE/7o9pWhnJMiAZw7wDNfrYeiymV6LZOHdA3d1VkBD
8gdmJ0gQc59G42fYJe06n36+P3KqhXrTdXfX1bOqgNLXIi6CSR5hfJ8unsmm
pB94NOFBbYdG4VJB836x8RdvaQn6W1IxhnuWMsbDjRIR9pJjRAc/NwURop6m
j183iekJCav7f5+xPLOWkzZ8BTPP5GMINfsnqFw8HYOFRIlXgRUHAFTf365d
q8bRJmxSK0dg8cHLJEh/y8fv1cmDEzlOD9rIol4JiAhPh+qJJS99X5QCQvaY
aeX2B63VEcZbRXcrgtaXD95vwX2RnXj7JgR5StzMaXGiF6ejXGXvyBHh991E
OkUdw9y30cosqisfxXssb+AbbDbgwEAv2YE6j3S2VBp8mkOpL/j6Xs2JhRTp
JBAgF5nYwxaHi4FGTFu5K/fxkROaQqZFZv3Q1AN97uhqlS7oVLluWYArr3yu
EyPdNuDvNZAx/YX3xWujlEUayA4CGRFso8Nr0PzvxklalckNwYK/1bcS2RBY
o6FR1RhRhw1DY/bdUusETrZvChEgHp5Y78VjF+YG+JyeLY2i45MV/lrxuV1Z
lXe4plMeUiQb2keCdUGgz2rX7JfU4MFGAcNt4ZUcfuSaswwjVKfdEktaUt2o
lI4zUh8yNlXfCA17T4qTbb1UXL3Di75cPV5k8XDf3NJ4fln8ZZpiHhsKyKKm
ELdMo0knpGYXSDGev+JYFc7GWqrKgQp8kdOANbkf/cskGdqoz6xWxrl4p3v0
u0Eukb2XcUzZIFKYcJQkiN0Nxc0khGSCzuUNEi22V/lepOhU/Pvc3lfTj/BS
WrzH5K11gYQGe7gI9KLv7SKL5Sn1AvjCQP945/6PnUf5z+wMHsolYRlMlqvc
jXg6NwoII0n+JmGznI7Jtqis1M8mayJM1AaWacaszh+qgBST6BSKUM+NUkIf
recCCh3P29jHhCOhYU4NqOGL8t3mon2r3w4hLtNjBIb3EVtNFdSfoF6zXW1w
4knIa3x8iGEte5gkr3tl0BRx4JYXYmv1GR+7KOZHfmoXWr2VqeGqiyfjOfkz
gmFnld+Km/szXyWAOTYjNPlWco7ZoSDLqj7U79kk0ceNziayqaOwamt9VC09
1mUZ3X91M5i57TRsWWRaqQy9YOyu3DNw82pvIB7MgrIk42QxgYAeJ1eWDgQY
k4iLgfqjmLrbsLUVYXKJGH5NhBlj7TxwKB3r/1wWl5enAtPNs5GoUlPiT3N5
Xa40cBTk6U6y/MoTAa0gza7+tnVxNQdUZLCUZmAMhnLiFrrFZIIyjvRuCov+
2rHoMOQOmcoG5N0zmcxep3kgFMqz6bS3txeuFzm0kW4xCNc8935ijcngMLgU
zJRMMrokB3cGIQjhILRuaGaAPGwp8uUKVnxScpcLWWABbwy6sIhhoepRuDqI
wMC8AfSvOow1+tsRaWGwTRx3Gx7gkMAUsobMjKl0DZGq8skFeSs6i86PhWP8
I+LKjM6mz5TESlX1OhWn++YCIFM7axiU1RUXG2y7FjrZal6550Cu3j02vJHP
nx6U4ZHXiHsBwaZX1jpY4pcGoQ52Cf1ga5o9jUx/RHYMW/iK+0Mpq/1p/PeS
7nC9fZTOozUM/oykSw43dBsSrls3JAFRpAe9vavdiKO5jOQ7hYvR0dQWiRML
4CQxOdblW5VRtawtPz2g1lL6F4ImuZL9TnGNEwHo1pUJpmoROhp8cfZdbhZM
A8/Huji+YiBQb6X+2UmeiBpJXlgwFHZbiln9sb8H0uET7Kv1MqTRzqn4jV7R
FZRQjy0svqwjfOYk8Ix0L1BoJEvCAuv/srrtHE30fWLtFx/cdOpZC7GLf5kK
TdI840Goq6bRmbv152YDKNrmrubQIIWa5lAPOW687BFAcIT9fXWhUsk9jeHw
boY7dCc6nfLURMwV89blkZdYpBp98xly3KQqIqKMGOSDnlBSUKSrXax/4jjm
6x1cXL6NjF1mEKq7AeabFNqU9hN0L9AGexY5D4wlEEM4N2gtYOWpHNrWzU1J
NGbyuKIph2i4vivBdZGJ48PWa6u8HU1wjT0ZXW+hNIhEgq8yglntHszqr0Sq
X7+ZIJa4kAmR0vWpgR5FlYpebHDBy2JnyfadGKtNvHhHL1xF3HVb933hH/cB
/tPcAZb4HaUGbABeD/v5p/nGvsEy3putJ7IN3YU/hNwgJgr9fS3NxB2VO0Di
PMkBDUAeSbk537Ymm60r0oySnv118RI1f6i+OixHJBfzZFjeoJ89+Zka8T9w
clbY0xeZQlBeGCQrSrdWjVW7b43afYyIawqhmBNf56VDHqv8gZ0zPv4rHik8
AO4enS0NYyt9aEW2aXnP55xzU9Azt04aKFTSZLIFoMMzuKL9hqw+/LUfxz1R
K/h89yPvrWAE3axTMM3uwAXSlzaS3bKkQseMksCpvbjPOb8w6vfLiUS4umyR
wzGs+iqxki9eD6QEPBMo6xymhtJ+FnzjTEIxw8XhXzBIqwZYhBxngyT2pX5O
AHfsNFPVKPBJ183gbCftRn0x0MXkhnWxiQ29+ub4T2OSuEDEKf9b8u+p3Kcn
KjBmJv7mVnPCoItd5RZEh2AB6d70CscW7SOpcWOfjX9a5KVKkqEwjY/pwnMf
Mv1xfuqQwdOnMxIHvcBuIdbA9J7IYGI0ZcroPsrN8fQaWu2ymxkuefJ2/bHS
qE2s34Cq3AM4XcMnVBNpGd/iluHdgcT5HeDPZhL01VhzXnYno+ZG5lnD5syC
9VxAu/gslp82Hz2o/hcu5QVqjqa/yPnBWNMEwk1agBGg9sv3CR8FZHwrhBLy
Ttm6sinJSbq5MLmKsI3vwiGLzMtt1Lwu7Vb92Gh6h46y1zP1peWQQ3LE1C1e
WuJ/Q3tuecr8E+qVumH76CZY0/npQ6CW6M4+AoChuQGqwbOQMZFeautXeclk
LFH2ar5uCr6/EOmvWh32GrN20peqsq08GhW6T/UouiNR652VXGyUycvXXYbM
xUuHbJGxr2Ux+gFOaEsataSl99r2HxZsOsmTf2fOxuZ6X0sYF6yH4ZzE80D4
orfPBbcc9SmEKdqFoG7b7oMcr9e9HfEZR4ms5XWaZ4lxPnDUjUxUdNNsVh3Q
vOh/CEvW95Fnph6n5xS2/gNTYRrPcVinkHa708EEv4D7FbcgEBd0iMS474LQ
fv1lGAum3QXWC654x2gJdqbr0Q5HifhdR+AijkdA5DR2sZRB7geRl2G5fMTt
B4QLI5pZ6N9v7tOGBrxb4GezUu5bi8K5DJDIomTTdHpoiBJ7H26P6QTTj079
hsEQ6nqlMlwZDHGW7MDHuWNsXqKOHLgM7su6ayZseaIYaa2jOdEbi1J7SVG9
SdvWaMun+8UI6HDSnukyc4JdwWXJFtgLu3juROzg1UTIAXsbXnS3vy/0Qv8U
tQdzMmVqLOiwM3dg8y1Jb62dtn653RQIvG5tA196QLJD8GuEi1KHsrsGgK17
SNoGayDlQ42SxJPTeldi4wRGRt1vKTkJzeqzFXqURzp1xeOOjUrW8STIoMvq
ahwt0zmFsgNWIv4UntDyfgAjfeCpX6IYhnN6JxGMGsTa1+zqvQ/0nvektsVn
um27KsyajC5n1pH+iEAhChuU4diXxJF5Raf9rXRHOkf3wKgnEIn1gdYkMT09
Jv1sODWRznHKv/lZl30+Y/Fck/E5qsLahRNMvw7CsOKiJWnCpkrVxG1dvfyd
OivWntFAob3YGqyy5mUp196hdaKY2PlMt/4wT/TTgyoxAiivNPUdqo+2uIkC
Xy2S+5JjUFeilo2GYdmyaawNLVj1Fns7C8SIpqMCPpkCtZUhQpjCRTgBYyFm
acj0i1mIofGQNQyNzYuK7odMIcHCGAMS3l2iVfdTSh0d6oTuUD2sI8JEBQQP
YVCoREBhVm0S95+WgFFMteVQthvUPBRVpNZH3AtYRzkwGGZLC/EYi1Siy4gI
m2XzUzjeG5RQBcigMQzNZ+Z9YqR22VWk6NzdDqR4IlWz/DFIbSzT2P9RCbUv
bE1DB951rteIYSZcKMJw0hziDQVppvW5+RO89+8AlUqlCuWqLqQpgDz7JoPa
BzMyVSEM2H8j7dOVJqQhU0X3hyx11Ikho9pLesWTKbfbaiZrnDx5Dx0AinCR
eNO+M/yXl2hchLc7U0y4ndyi/in5oYFzBwuhfUTze9Ib5+7CV0LYPmBprnAy
uWG48MZXlqFIMGtf/E7wXRLLx1YxD9s1lNDceXHCH0FmJZ3KfejbK2hPbegr
TRWVd5fV10fm9pfqHpLiNUkQXmB6Dzf7uByeFFp6QbUIQzPnKjt1Q35C6z26
6zw5b1lwDu9D2RJQQDpGZ1pi4kfzLREd75n6atXOLpJdKSqdsd3HxRjv9U+o
4StcuPVdUDidib3y0Rm44MiqdIrI1AxvjzO7P+ybGcQOqjbpxL2sUPkl/UrO
xn6R5Y7IDq5Bo+2VgrGtg5rQNWjhij9Lne3MOV/xuNVaYpks1BoWgpnDLU+w
78US05W1RtZbXJfK31lFPDrPLUui3OrHuJDyasq/pCVqcDSXyUKYAcQYD7xL
PfJUlCuH92DIQtacLW+CnwGxuUmtD6EjAReEytlLKFlp4+CvQx14RZgsXFT7
zROVQm7lXCeo4tAC+/AiNCfQN7lIXwIyJ9Pbj6Q1G0Rat9Pf+XmIVxGg35Le
0Gek6uTO+Y+wDs2By5/bPjwPEdcK/DjIcX/RYcA/QklbYcBl+J71N5yU0Jw7
UstzVaLsuRNG6UKojY+6A/cRq7jDCMv5XYpu2MoZuM5XqC6Cvv/j5ghynLJM
T4rU1MhN6qRXc/IzY7GxRyZVTZvUul9qfRqZq/6TzewzQUUblPigWO7Xp/8e
xBeaWu0N0dnFCuEewE4MUIwQcHEm11G6p4yypozePsDSt+Zth5aFaSGaQdxC
PE6X3OyIKPhAY9b0ruZ2zLogJH1yuBzvwZTeXck/r7uYucriO4CWkGFUpNum
9bgYuPDuecodwbmtvDzzObdXJaTSJpSSRbXy51d/Geeyy1PjZmtfIo1CEyf6
jht2M2Eyx2TyFJDrnoQ1pRiE/5nfVt6WpHC6yQyQ9QsMCHQENL0ecTblFQCs
qyiB3sHLpljfXPNzj5ubxEM3NWFES4iB3ve9M0IAq1PTKtlO5F/JubXzej3V
LVReegPfhfW+3XOe43cac2n1rDjLaYxzw+H+ZCoSvr12sYkVVAmQQzDl66oF
n3CHDLmjfMncOY+j7bnFnQoxvCTr5kcYm0szFpbGCETbvaWSrz0t/GL3Jj+/
tZauTbbJZM1/0L6ZILQQIPaX/RrNGBAwghiFYXZ5Le29rhrVRQUNtmbRqfyx
I/KMa++Y9Y+l+z1JmfJVev2J+3Rp2Rs8V8DsahV9pJQYzAcc7XSbelR61PWe
/H6X+l2S61V7UVIZ8yWs2LQAFlTTztLaTNmwC/Wcrahya1VVNerM3KzFOrDG
MTJad5GoRWdmK/A+PEWcsvFwqz1ZoKhKXAhzJxQN5vYo+il5TchM0Tz0AbLM
LI3VUsjM64RJtKmc6esqrYYq4dmW2rzStgYI91w4E8FxaTLYtCgn4YbZNx2C
uUKSHk86mRZ9tawyZw8hbAoPymj+t98E72sDz1Qsde9GgAtqR3ly0/bLicct
vg+PqDtWXfaeAcdXyUOYqqzdOERgbxuYz0m2sUSXqWlbSgp9YaR8PJw4xOJa
0jYid4WIPDF6zGzmwcQcjEohoQix7CbKlBCPCIykhKVMJVozIjSYckKmYy2X
E1tiR/xUvKlM4raZutP38vn9oQORLagg5h5L6Qni5BlbnDR8wG+w9OZHJKTO
snf2gE7ayMWJ+2qsLMeo1jbPu24vJ2FenWnqx5ni1CzaiaiTUyXwo066M0p9
sYLShZQ6z+lAqc1Txb8BtuvbJ8JdMPgrzK82k/z2z70q23lDrRi/+8X0Fgo5
EEGfD9AJJb7DNq4Nc0p6B6ZPAF4xZ5xdnvtECK1B695Zv1A5Wku7FP/azYCj
hu8/gTHHpubnhyUMaEBaFLoRv7EpF/EPtMLb4eIV9ZyRWHIU+Zr7Aa0b10bw
lq+C1As4X5gluEQRH7brE+QmEpacpNdUSiP4f/rD3UIlNvyOulI90E6D+3eP
2/jZ2wIODFGNHYFfTI71zgXLNCzxF1lh+R609V3ZBphSA5g3uvzReqduiw+X
Xu3hkl8jhyUg0byB96wgfHR3UpXAmhGNOd8aNpnwQIXp1i4YjEyllZVAO6uy
TfRcYt/Mrtawl4eKiUvtTFj7Wg9GFoWPeiErBHL+MOBZwxxVuUm5UbxKpaMm
5D/tUB/j0ZLK8V2IR20zmYle3aE5dUudOtTKNeZhwu9myw6B0PnWhgvhw0pH
8N6F45fN2+vZZdpPgEhMVPvLOvrfZO6sjZiNjsU2yqZzaYmN2H51ziBlm3Z1
ehyyrpbodAkQK8xafGudZwfiYCb2/Q+Pb7KXUENd/zHSDxz/+Ia0b5DWoTHU
um23rRuVHh/1gimr4yTdPXSPzoYUNNiera56uhUMQf0G8EiYNtTO7TRqG5O7
lFh3wk637uw8AUSTyIlcQwrgZk6xRRu7hQnREfBml728zV+tgfwT95znauJf
JW4V0o1vmmt6hHTVPEJj5YZcSN2xHxomFowJJWzAQJzK3sPwHopM7jHNns4t
5LgIVGqdHI+C3adu4EPYblZB69uK8czDblBXVI7geqA/wOnBjJlTVAnJfoPB
uZgKtBVYwmutDpZo5cp3N0wBMIFUuQy0YpvaT4M0x6LG4mP4HvXTS+djV5pi
ly4g7BWPO2KLibvZ5M5Ilb9ppaRkv4HJjpgEF5A1OJVzdmsYgGdhZxWm5vtB
iptkmqZfoMLJZOi0NVsuqh7SyZe8dEEzs07A6u1NeRPcBpoocoL2sufCsTrT
+ORChp8/flU3Vl4TDLHY/PY6XCWv805S0AZRDL0srkuk/sBWEHMTszfm3OxL
WSTLlRzdJ+7bkyF7B4o9U7Ysd2FHXV2C1qowAOVwDxsEifCWCqEuuw9IAC65
sxtBi0H5DsjNJNKb7cOhcbHYHKuLp+UuIZUO0EqW8xVjL0oW0HPtwsAE0Q2U
iUv6L/kSC1PF5cGmxTg1GvkWyXAHSHa8XUWM1u13AZxIwT/bSRpN+5AxKqxz
je9dQi0iueeb4XrUks82hZZTaeqVsir5uteYpSy8pFSsRsUTz5Tkiy0gi9eB
RsxbfjT5xSZsRI/m1oZp4Hzx6iKneLE6TCdJudU4UvqciTPGmgI2w0NXUr+0
7XAXU4ltU41Q93881izS58T6znJ3GvDnDB5r9N8d9EFqvEmXPp3EHnvcnNfz
3U0WGZmql0o7NJbpB7eYu32uwmP7qt8t1DG/NIH3sEsd1xAMXjbN2B21VjTX
PPfpm1pMaI5ogSHDy/Fhn2sfmgaQ0Czz1DCKLFgNTp6KIQ7Gfn8dVampW2Uw
pcNkRda6IKQgI4ByrQEBuJ7xM87sjI1tXNfRjchnWgOQy/UEGIR1Frr2axaV
ZcoCI7Wbo0vsCZ8f04/MdlUHR+gvUCvN3+XwbdRDtvsuVr+Mz1+A2ekaXnXV
Sm4ioKkE95DKXIsBJhqDbzZUXFYNofYOmeq7A+myOGkR7qMkpBbGWLgjbqdW
Qh1/f0fepjXVzTLYHD0bZEM4cEunHaZWsCRvlUgdhvTT4CINztyqoOm2UcK6
z0JRPcmtlciLqdvsGLx9RsUt/8DNj7elMxDkHNShN9PyZqwEkzFXQPZVbPZ1
GfS4VKpt7qej+0YoS7b6blAEsOTqhlM/hhcojEWi/PGYfHmT/JPA0iqLilmv
sV3EG9BHIGs4UkKTH5NE/3flG0jZinXwWNJnvzbGkn9CInkjjgE7tREOhWFS
zjogyN9NuatZZVam7lYLJVygx+TQT6d/LLuBWPUkBHInwsWhhRJ5t198pfHM
SdjruVB+vKZxfMQREu5WecRjJPTNvz+vqCziKY8oxb19mPSfDeQapv5Q1Sd9
88DllIfQvwHT6ggtyK0Nc42lZhXkpLf6jSFlxZIaFT7aShw52bemMEDATOcy
wlQdgcyM1ldSxS59bQ67ZeDYHHOa/j4/vWJ4n9kuc63yo+nkvQEU20d2AqY5
ENV3zenk6E+BUGyXiY2oolD4/nUe8gE5MKOq/Bo2lEGOm8ExzTl5eQk97wME
Hjvdh01DNElIVBP0a+H3m3PeU/TaNXDBs1VPAm5T6cZhndWFLofxY6dShJ5B
UlOyNWcYJCYNGF2ta7xfaC8N1z0d3dWqvW3VDcIaRAPva5UKGHmijR/VwEPF
nPQj6Usap9p7NvQjoSPrhd341BEXqjXVYJN0vNqkMZfwakDKcNz9wtNa82rL
Fbr24RTOp8zxYB9e1IRbmonGMMAOQo8jKa827qMO83YQ0asLmS14mhI+zNYn
0ZAfK4QoLm9cc+xKoCwe8gIJiaEPIbSdWQTX+adRvcqGVi/oc3i5YjTzZd63
1JACDsWdIDe06cpiJP1oVOewbGLGudzhv2vKH53A1/4XC0VfyJX8ZVB1oeSl
+jL97RxRlodnSLW0RQS1dbLpxV01Z4wSOi+3BvAYTLbfW1L88EXVrn9HyaMe
Miwkqd2AuGWvwpmaASwhwHla7YDITpdt8JwaldCjzib0jSPYvqoi2RwvhrOj
Z7htERgagQ1pdobM0o8sFZm+W9WAXIjJfdcGQQGPxeMvaK6+23Y4wq4HugEJ
19z+adePCYpnHjrjvu2MAsXKAjyshf5f/8sUsM0U/K400jF8st3VcH9jBhod
okI57PEODPimGGMPKqd5YUpZAQTBH7e10uxZWpiFvNWIWR2988e+u4h8S3EC
on1lXcT88AKo3eMuQyIse320T8/2EXh/IAjJxaaPzKI8gzzq0pfpRPRYm+ue
Y+mhGHQey+07BhqsVXBgNhVq1TUkGzLgg2JXwt+Gx1bh6/sisc4xkxooPkqq
ZpmT5LH4ei40I+FNDG8gnsoXc+Of2b1AHOyJXeyPOj3dbWU3lldy2lIRQwSY
K+eepxQQ89UZL0gsz6sv4aYnWLQmFZGhaa3MCFxn4ApmwSt6hFXO0ia3IGgU
XoN2USaCTONPAoZ3yYET2nVA2YzrXLv4xU/yJvvt1gAZHfoX55Tmjbi2rzs+
mwOu/626kvJwEe9WMDkS1NJNgm1tf9p75i/NyY8esyThUCZg/P/sAQk1vaRo
vwAevi4CSpiGNpcvCAsyIiEfn1kqJd5gYILWlwVRSaJb7Kf8XgHhsvB8JGaV
sDmjQLkBV1RAtCCXcfiZ+RufOIIXf5HgDfHX1PHrRfjIjSCpFkQPd65Jo1Hn
j7rug/fxPxpk0RcDsqam0uAx29gtG+VYwuN4nko/JSD+WNuuPIhH2tidc/c4
T7EDcWZi8oHIH6G0aVLbUJa3MHCU1jE8hkt+jcibJWlyK1qjB9Z/Dq4jUzvI
D/fVOke4QU4C4o0plu3ULFJn0CaJCcI0TpPZJW4McYtUo15YTW8vCPnuXaGV
YEnIXS3mUyM4OnhUSqpwHzbX1TyzQvzW++YoAJvYm7QrDmxptON2qcFl5vkK
dEeNbZtM5eXrdTI752q7UQWB/GnyYgtjSuYc/BwGv7zGLWAznRDSrsFqsoFV
o5I7aUGXXlGTk5DgiWgeNNUBBNjewZkvjzUb7PcmwSj5LhXe6vGAUFK0U4RB
Uq2YXeMvTCYIBOn1YKZzGRV4hREhcFrCM0Mzne8F7YRM0P0o5lpnSMybuLj/
f1w6l0+EisjHzXp+meh7piQdZ2iiu0kkoigLlivo+yHQGTXUxaYOor+lpNHE
eh+d4YkTpqwZ5u8zu/sG2oJSlMCIBu3UD+52uMN3Z78qQ477NeIl7TNGF3lf
lUIgl0zEYAtp4bi5JoUmO/zTmAWMteIEDTpKE5eCEzzw8RY82fBulhEhPtQG
P5ng0Hy254Efww552bYSlYAqYxFepo3mkUZ+n4/0FjZZZPfRgCQnGWAya7D4
m51dh0Q8DN7UT+WjEpazIu7BSeh/bMJYWq0sMTv+er2+nFXTo061MX00K5Rw
o7qADg6szItEZq9sSdyPIrG9tXNh+k8sDggWRGFSqvhvVwFsSt7+r5xhvTGt
1zFRZ4Qi2yP9PqRVS47BARiccgicWUCC/2ssN1y/AAg2NfeEK9OF2ntAYyZ1
HpBK+RO0Tu6qZTfq+jPd2hswYHbFLxpjh5cIUYCiGTkr+B3wo+BudjnfROmy
mD47tp8RpXmqFkDHCBRzcJd2hXwgFoSQRboSJM99duy92ieQiikB582lJ346
sqf+Xy4pWtP0MxBiDkjyOuDReMtSCiy5XoktZvhVwUqIjEqoE4ZrDjulCeUV
sUDLs/Q4waOiZYXJzZavM24w0pqQVhib6tE89hGPUPOd+eDwz08Yn3r16KVB
Wq2u0s1mSdPZ2Z2JaAnMJS7uFnpZFW5eRMoeH2Dib8j4pANrfc6wSaKMqaqY
pRx6EJc9SDdCW+cFVXqv5Y1NiRqXLqmhBz+tCEQQCxXfgD9PUjkazPycFkNE
W2BMiYlZ2M1Bp+/Zim0/IvfcqKT1DcXEkEH9rb+OKQemzhHmfECJ9ferBG1r
2r8i0KpJSvrxSn4dunwHIQWfBGoEn4NA5JEXY99bDhvjXe+9SKg1X1ti9XKA
auj8uKmqvXNx3iqC2VBfpvscB1U3iVk+lBLNMgNIBozbyyM5dQmT0GDzU23K
3C0gdnURYfwiblzYNBECpbfVI6KB+3l8mAHFnUv7j/CcYki1XyjDIA2fDPn8
PHajnotFdS4MKN5DrCznC7Txfub5rVcLiajgiHUQM9M+mN+j8vaGbtBykxlx
tgJfJzUXA7PCWzVNK7zr9iE999A032kfFffYlPnqGYkDur7gKd0iCrvbNeYX
2FhurnI84Ro95glSTvrS0zAI7rEWPIOidCZ307AFHR+pFxGnxFGTPKDww4yT
HgMt4KybqTT/WoxEAbHzjwJh8otvlGXGJ8XlZOFG/xeSLYvfu0b0wI9DF20C
6MZozrU7SCQfbHgWUQhfx6R+lqqIdwZNQ0JpF7mO+BtQCVBXi+pgoCFXJZBD
039ZVi1thdpaBElJyBFFxivSj8WwqD7i2WnXr65iqkOscQHLsf038ZFR0fKq
jUgF0jXZ7qirG/YksQZJBWFPClFPxo9WigF9bMSPnvMdHhaO7NH7nA5z61Pt
sg/SCmmoodFFtlzpTpdGitMQufPI2DwmyecUgTiVedwrhOx0BGdS4aBvzo/u
fj2YXeRpyKkL7Pnx9GMdj9RXd35ROBA+UxSNp6TMnUkDlPDU3owmirf6fsd2
KYw8dvbYwVAJVKKn0dVXCfQp85OW63UKQk6Og+optp+YwQDNP5KOD+Ir1Vty
9i6SPshBTD1OJg4Qwl5yBeH2O/vc6miUQFUuf8PUdaf58wKMWGzvxuuO54PF
FWRuLe53kzHZIfTZNfIYH/YJ4KhItxq+uv3m2E5aQ1UiNilDvau4LOlANUjj
8SoyipMuBg5dFyqA9FTJgVIUTFn89EpfH5JPK3KBbPi+qukmeLBZbsFDN8cV
EiyNv9CZJUP/vZrI/sKRBSoQbKhfPbTQQjtnTXFheICcDHxIjrnaWAGmOqAB
z7DrKHgk6NjxAHKKRulwc8zytstngPCA9veGKaT0zhvMDBajVxjlk7VAiTTZ
nmN9/F6tbg3+FMuKG6zJgdlnZYOQjlq2FYvdfNddobtCmdtsboIZTB0V2Yfv
WPNP9rlywwilIji16K8d54+mrIq+Ea+UuknMlG/PJ3m8IR2CuU0WoKC0L3BJ
nK4GbfJAWqOFuhOyLoAucwSE7NIZjsYvBbu/AIys4WWW+MXoJHG4lbi0AkAB
C+f6OB6PP4GVBPLgLPpw42ISHfFHDWQPSqpkdh0boN6YaVubrerYA/6YMITc
EuuUrQGL/PH8kYZcb80G2XAE7MVYB+4uRjGRjEaiO1HlGp2ppOd2vTivAI2U
xdHT9/PCG/0Y+3pz9OkAkYDuR7T/GJQ6n7+zOKmnYOrKPck3frfpzd5j+5Tt
UweX9pfWDpH5tbFdQkRoAg02N14AlOuvMn1Cqx1/h+h3sjQlV9iWIwz0gRbA
x0DxQ2qSv/xnNHRqqgA9sl3FVm+rn/J1GDWX7EGhd7d2xYxY59goT3t4uzVq
bJNwTFFpfJ/QeLQekLri/FUXCEvoHqz5z7IHfU9Apxo54txjOc8M6FM8iyDS
fu8946TPGvMkUGohnclewxowxw0bQQlppnpyGpwhPjB0om5aa8IckpmWXB+O
H4YXd21CMwVLAOCOhxFtsr4kf1ngFNxZDrkvNHKalfxwlsAhMM7dwgPlOMMl
88rM/H6l6eEXjAxG+ZP+DYCTvk0GR3WhlYyHI+VEaBktPL0aAPHEeA1lry7u
Ab9O2pzthrdqGFxY6R5usBU8k7w1ksEvcBhIyg6807RL1oEReqtcqFsvfpzL
3Rp6VYj7O2nhb7kaXp06dAa2ICTttvoeyKOYEqkPmTzl+9wfRZSTKgif/QRl
kzylXYql2r7ZKKf2ZSM4gz2ZE1z8JvWNDyErq8wL/u0eX3xDfgqZIdGaVL37
AOfS8e1EANuQTvMqtCVQjVQxWlQvN8jSrLC5kDSWiWVVQOAOz6no5Xhglp77
4I01Ek0zKKdAMRUv1MY7UAm7CCduO/zpjDE6A8B9UpDHcrbFBtZ51Re+1EMN
U+U1F7K9eI/OXC86XRBYNYtfM9Qb+4VgF+ejDnoOvbFx8AruFOiBASkGxt8H
4XbxXhlyXFYDvT4KMHwuH0Hq5T3T23mQo0T+IgK69QbS5x26GuGhHRurFb1A
h8Ips0vY14X5C5BVQV4VioI2z3lMt+1I/bilRWCNPAi3zgc+VMMmPWkTd2VF
HMMmkMcepCscNnLFS87LJ22WeUnxGggMRxFWNnSvDzkDydV3dtxSFO6EQhDk
TW6gSCtLz/+uCpXD8wcti+gQOXVh9KBwOIkFaY2dxjG0gJ4BDwgiMWmIaehD
gtFbykE9kT729WniyqK9dT3MpQ9IfFIOUYNhyeGezepNMtOimRxZDorEc2k6
02VEmt6CDV01DxetqIlL53P137ujB2WJUll0mNp1eYiVNj2ItHHSsLj8wtE3
4YofS/TVQ5f2lGitiBCZY3uryZBt1bbkS+8ZLfpPNh8GKAFP0gvjpT760IZ5
tPPLj0Uo2Pi1uT1B3KMC9ogq3nRcl/05GQlUjUZ8AP1OPKn89TMgzRgMh0Mt
FzePT/aLcJ+VhXEdpcbe7wknKfJBbo60dnc6oopLR7YR1aBJv9KI12OKdlpw
zQZS+/fTl7HUfSgQYT4LI77fRkeeX8rzYFFOjncrakkjshaFW3bau0DHRnyf
K8J5KhVYP/tsS6u6Fz46imzh5NtYypbqcTvvp/fvPJ+W0gu2vCLcRWSvOtC/
J1VI05zOZMR7+ID0hjrtfTHBQb+F/mPHkw5yrhOXKGat6jmeJjPKMViSWgJS
6xS+XHCSZWQtKxe1ZNYHqx4/V+9sLU1oG1Gq78dVA86uN3DNwWK47dcDKDqv
C3OzOau8lQH64Jw0qrxd3grtnsgsuy9zxmze2XpNlVfpINzibB60npEB7irO
bHrwoU/Pbho3Akd5Ov03NEHjIUH0/snD06gEr5OJbmdFw58e/VliQUC0hGJH
tFD0aMcy8D3PKL8+bT201/A6XnFuK3Ijupm16iM9joSd8w/4kYYklitC50Dt
AQCq5xCSIj4VA6AnpoxzUTaDppkPKdlj9gtAZzHGhUyb3gizRJZSdSb1exZn
IDH0GZdAgK9yWpozMBDRl/IRKAfOZKf96H1dsya2UMUNk+CnxaPBOTcCNJke
QclTlmxYgiAoAQg/2rCL+0lVJarGb9iKVx0uFXocmLm66EBtVJXDyM7Wph4G
dOeN4Jaa8/NlOrqCrp7Yw5L2mu3eET4qsl3wnkHMuQ05DcfOReyq8iBu9Emt
YPzgKR50HsBJ1M/YPJDcugZXHDC50pPRmmDeTW2rx5yNu4nUAIqDZbJyBDjt
8s8nDicoJ5rpBT/jFP1in3fJMyMIEl5YE7P0CVJ8LD65Wc91BYJ4fLPOKpl5
EnSoZ5DqsfWYq8LSgxAscrGhHD2Ax9xHiUpQBE4QaKJZRfRwoME78jcxLVvR
KhQNkTlHsGNxFgINMpLGrYK4CWdAjAe7nTx2PHcecyNxEiOy1Qv8a7y1Ljq6
qIbffCiodP/Plim4TL1AhqCBJuzgzHZ7oeE2m2ofCkFmJ178+o6hYwdfmSdp
SN+4W2Qz1nSt8dirR8U0Ui//9Qo1IMfBEF4QtKXSkTuZ/ImXzl523lNyFeiR
Bax+kDopHPWdK3YruGhqx6PSA8ToQwIq2K+OKBcTB4L7H2aBpkcZ9P7nwnh3
AvtFNiLiZXxMMPmRMGwHOkVxHlgCiH/f818jSJExgtiBuC74vey7UlgjkRmg
Dw3w5PTKS3t3acsdaO/kroWAhNuOFexqT6igolWWPQPQzEfz8VgxGCHMsnoU
xclAFT54FWw4aSkDirYtiVbVkvXE3suQVYcUWbkBkfJ0j1ZYhqbHhoxd11eV
c6ecSmsaWzsDEj71DHwF2Z07MqBfeiMs4R1iiLfBQ0FQdtVhKZB+T8RszgVZ
qFvNEc1RJrW7gzlkxOyQJOF0DjbXztG91XHMEvi6/Pgz7wsMPpNstdN77fSt
ax6Xju0C227/L9xFX71xAcagA5ErJ7Qy1nQIE9KO/p49hKcF8YN3fok9H4mf
LBrlFQV8IxVmmrI7C2R1TShli6uDmHOq6CcoiX2NKoGzG3zkJPqRDNAaDVtT
N9KKkHORSGTsjctgAgGVPijIWnzGEXMYnEAEA6OZIVQbrzCjDdwGr3Uih1xN
MkHAxyPBZsmWVn0rLL0ew5UN4TyHsvqPlRv5T9QFqMBnDHO24t6dLuJ6D4Pz
FPNj7k4eARWHFrD74/EXk5Dw7CwKqJMkni+Nfa9r+cfIRGT2B5lwGcrHh/hS
a4OhCHJOlntBhiwDGNWyvKaDDUoMEJFhNJv15x1HnpTsLA5KhPnB3+G4INFJ
0HrbNR2um7SvaINLpJeQU8xr3dENV+28Dj2Z4J274kRgG9lIQX//gOmoXheX
0x9MIOp6wl//JsRhvRs54GCTuI41qaTUWqb5eRY9U866wwOrEWkbqfmjPGaR
APSFyizb7sjfHAtyUt95IzGjzrxqZu/IWcC9Cuw7uYKEFpfkvQpe7436vdUe
TDE08tJBI5g7SAqhemefuNgixAz8Jg0G+6BQZ9uBxn/QXtg+j1+m0QDOMT2b
ZwEvjOA1OKh7rk7ztsWPYoCGyDqaJJqCgxTUwy5SM0lavwz+9b5W2fFNy1Qu
Kr2ugh9tMImpXyIa2fQVeKXxiHfbef76SmjSOWAl8DEuIrji6Nekd6zBPowx
5DF9MeyhYhqPNf4vsoenqaOFps6iQOFr7gxrC/uITInqiXRQtuXLwPCxYdJ5
dMbbQaiDPpBOsnwj1/ATAFUPvsoGkIJg0Tzl2Vn5gj++boUaUB2mD5OwsKyB
CTdKEDmlPmrgTuR161oy/tZ+7SJJEDqwqbFgdnc8IxTip3aoY4VPqqq9Pork
MLx7RakwQ4xtW2zBiydLZeDRHtXdiGlWPtjMwcqBKUapMzs51JCTt0D8tgNM
drozB1BcP93uih0Uo6fTpcM/4DTjvVveIrh/xHMsMUnWb70M3+fO3ZYcMBUB
OXlEG9WSzKl0JdwYwMSGWc3GrkLpMRJAGEI8gAV/4SLza94utDghjWnwWZ/c
++80P+mcoZMFcIj/s8/zDmijkyxQ7zKdMT45hswssBvkkhMXs3DWqP7xu587
nM58AH9/H/3Z72Qqh19AdUAZMXp5tuj2CMilNYp2aCeDHPxo8qRL+i7PpQ7U
77JUUPz1ONC31frVvZM6kZrLNywgAJg/ZccEYwPtTK+NVIvirN6i5MgXkkeM
OT2aacjhnjEctDEIKr+abtS+0o+l9HAqanw0HQw0ktw1EtI/dqcyNAfVyn7g
ZCC7KVnfCVSIu+sF+bjN2dn9PVVWlazSozWomf6IAFH57/sB/dV2/sjU7ake
QmgcaXHULixPECzirlgE2377UNzdScFm2MyrraK+vzUd1BTsTzk8k9XpJLWG
qoTjxv1b679Fi3D6/xf25VwNQAoTfTgqGvb4vGWc7OaF3mFVNr1WgwGHQCdx
ug+CsqDNwIawPZqaWgHb2LhA2i1kLANC4W1k23pOr3EVrHPjjfxZUWygM6gs
6FZlLBFG+s06j+J8GzzVyrMO69PIyBv2x4afCFToG5+h1g9UnM87/Nd8+kVg
oJ1Vv5L50dGN5xHJqSOTB3IHj/X9enGW7nZnsRMmgW/e8zu4h0JdRRohWL4d
rD6N7DmHBen9P+tTOadNM5bMs33klxkn0RJDDsLbZ42XFQYFPkhdT68KSDud
tJyVFitkotJoNEMEGneuqygaCkTfkKw0ceOvdLz+p9gfTjPVVor64H+I8jaS
nBf60UaXbt43PCa4nb98bLpacAc/qCuinipjb6PGi7sbIf+yqzqxzqxLTZGy
o8THu2GkJ0LGjuu+3MNErjrlWoZjS8sbdbAvXUIiNB+9fqG4WVk4eBW3oeBe
20hO3LmEOAyxLUJWFAsNrv7WsqRddys96GMWNJqK121yrbV9+AGauMqOOU67
3Iib37VkS0e5PKLJg+7KNmVOvYPPV7qVvXGARc7qUaKJh5Afhv7EN5wobQcM
JQV6OwKNRM6akUgycskVijRh3/e4IRZSeQZjKw4qOdPT5NNz6xoEyhPZ8YUA
A0noSVS75qhRjC1xw1BzioXw2SMvbyaNrO/cbpykZ7XCVlq+jKCWSmHzRoCi
+MTVRAC3LHPKtF03lahmElnhm0YmWWLNwIoVw6AG3GBob8Gfy7kvfDutkIgz
gI4YNggfPkebBsv6JZEpnB9JntJ8fxy2C1fh4U2l2SRvEFl49G/mx+pQOsN/
kbH6EpxMlfX3mHwqr40COsLZ6dbxZSCH5P47goxsBBFNJxvx94xySbHhW4G4
fD9vxqezPlrfX+tiFSMmq3lePJK0oE11yNGo+pP6ZA8Bhs3GlxXANcaBxiy0
5P0WvdpPzFO10GYUcXB0IkUdsE3i6oEHuAQvlvubE1h1Nav1NzD0O3jWuFoY
dcf2swh3UA5GLcXJ9IhPT1VAVVyhJnE4Vf6MzM3lsTCn994Lq1XYevwaGmtD
aZoTsXGuT+2ouySSQUaglxCJjMnMKlk0iX8gKjg3wJv7zwaOG2BQbvUgEIqb
lKJhD70kZq0C3hvGDIDyGdeH+9wpxhxKcmVlkyhSngiXsZ48MZCILl6Enr0P
3bAwDN3KgxDu+QL3+dMa/B6URuEPMOAPX1+JSFswft0qmJSPzf1J/omNFI7Q
ahrVeTSCVbxkYENiR1lZsbJSri77szVEYFO8KNKnpC7AYjOdjQ5xnn/drbVf
GOHgsCMY6MuxCwvToyVXNhaZkbY245n08Nn04wEOazwcI6aCgirJ5JZeT0Vu
y5LbryXp1EYspM8FI18azgMA7C6mqJ/9p21EOvx0LgC5+fl1tWjQGmo+hzJc
zUMkjsIIYwidBiL9xe0tJBd5TccGil4/+/vmm+9d7gsYkHOyqwZOzd+bOaSE
JQsudUVRIXHph5vGaIzYvmrMNE4V8Q3hCVdQP2x4KEuntPbyIk04qrKgR20i
CFU99A5YXclBItrhFvLT5sDJ/N+vsrf1QpPOQwSDkBC3uQh4ePSI314n1M61
p7pCztBoFLnjnXqNnkuR11ia/7TYshxNF9ZkAMOV6hrELp+COoRGW2t3q7bd
SwYTFpxDlphHpfcq74yS+u8FqUieORR39qu7HrLJCYY8bSf0TeftOcwY01HX
vcqkf78XAM0Pu9NVfL385fI10/u4z34LTI2wNFGXpttudrc0lgnM4/zeojJD
tOKgOZ8dXQVx/iMqeLVo4HST6tadsFkOMLaB6k6Mq4X0Ee+ralNGf2nXGL13
tfSJ2Px9umRV2oDEDGW08dDSIFv2CAzTrAT6ZjR9OOzaX4+envZ+TngBed0s
I6jZuU7JnVChDfoDvH1NZcAREzixTzMILsFilDdsIJ0UVlhIPZzQHQpr6ixP
V9YvfNP1lqcH3qnphe3dzNW6H4dzYxfWf8UYIqcNiHilHnuUvE5xJcVy/eIm
t3Wf0lSbF96ycmcMbU+xO0UqyXM3j2ghdbFe6q2Ajl2ZI9R1aq2FqOPtjSth
bIZXmKXU50U5qm49UtwIfndr/+8zxAN8GLUAHz6UJ8maIQG4EVfV8wC0jswn
rLdadGlpth2KLyASzpyN5S0uIuwRoUFjc0Hqu1jK3ymtO6Lex80ghZrQx0p3
k4onIiVO2ZcwoGo7TUDCath/d5GeqMaTV3PWnzyzyn8r5oHxtkVIW1dSupi2
A/TRo6cXQmGneO4z0bLM56GluYtWYK35k7NnLAKxLYfSbdGAlIXEPFYsbyyF
WumrqcL6lXbEKnvlYAv5XcEfgIrTglFDovIgyJHlpHFu/hFDVUQlTz6lQ1eS
mmMYPzHfV3kxPKRIYrDwdeGMbMeOL6jBoQKRtPzeeM4QMauV8MwqZBkh78h+
QmUtEbplm1BACq4JkQfbyDYFKq+ggo+ljb0piXVYsjgvL7iJ8uKKQrJqs4PT
pSjauHP/He012ps4FhWP2Z29dnHZpony6dcg6dFmNFxE729MWJkgp1W82D/+
zYmwWvtngCJK1nDyt25dpiHBZvQ9Xkgg0PHgRSyCwgJffLv5VwQTFy4pBQZr
I6I6wrkUxyOTYVMLEOkrkZfIFVRfRFivxWdknd5J/Nu+qjMk7KkvKSjgxpke
FM+cwJHXl1OpTLirDtHovGRAZpBf7DkyY0f/vvqir7IRy6hIgODwDA12vxO+
hBkj5CAYWBwi0CM2r6js1IQjJ+3MiQVSschPI2M2zXIMfXmjR/b9XQT5s3j2
I294V+Z1qys0eQbQpjKT/9SHofT44THsJFIf9Wny8N6ukuqpDMSxaIYJ9rZ/
b/uK+1kHtIV19sAcF1QrPf1zG1OElsC892cE5fCIFQgY8NLzkxhseVwYeK8V
AOrz5w8mkVbckE5dehLZBloagx5YHpB7shgGXUazSWP9cYQTTbv07LgMMSOg
RxGh9odxYowm9Jxh8qAhLyW7HisW6v7ULCW0L0Gp0M9PGhpFtGeqjkveBIOw
ka1p3X4nH6PBeTEtmZYimtSxOO7GvEvTdZ6qju62eWW+mPvLTsRZOroXpBUY
CQ/swKQrgvqrEl9M4ni7oGJpSXAsc3n74EOA/Eh8/6hI6FR6Td+s0QxEEDnl
BkVljn/srzac2Og6cZs8JGCQKewVM3exoLyA8cqPDGvkEdJI4GiZ4+MEXnJG
hRFcwPbwRpI0OCfJD7YIgg6F8+G7ozkXSYM4CDhfsZzU8o02HhT/tNcUqRsE
GRQHWVstF2NpKgcuv652pFjd2y/a+CVOv/+kEeGxz7i8psJt//7H11RI5t5O
iRvFu5/q85WYLPp/YmxeG3+ieBo+ZhKQna4mIX/7i1mH/SG+RAE607wtdKuE
yvF+9jsOfDEHZkuT7LElj5baws9hDWD+AIlu333C4nxdttxYtJWAo+5X4KtJ
2jah4znUqcSO928Otb8DZRuC3a7eozVijeHdDo7cCN436kHTLmlNZMiy28i3
gJiwT9Tol8lUhBfVuFdOoaFnb4mNiWtMe6rQyoe2GRD5MLyYYLDiaessP7+m
6Whnv2WG9zJdTB3zSn4q9KV5/+7Vlqo844ob9QNZuA8fds4nYA2/nevMW8l1
Y4603/lrcg31xGN96T7f+bYfyEci4nxZhO8qI8ScdS96XqCBrwjRF8fKc/Ee
rua+buiy0pSu0ty088ztaZpvsXD0Y7Exh6u7urTfzKX/lXLlZU0VK5WuMhfB
wja04IRGjdyqloKRCvL1eEdpuf+qb8+EKx3Oi8tnv1Dl5n09JZwpq3WStFzB
KoxkLKabPJowXS19rebyiRbS+nbJwLNu1JMvlO87YTovbo4ozslzOFf3eZ7h
glKwcSFKVANhxRYh02fgnuZ3VOMmfpiMK/EoD/GqJvkDAklFnRedFH1ScPnq
yfJGqUa8sM6w5je5SinToTfecFiSsEapz1d1OkLuKJnQHBoc+BwamGeTjj0g
K2m5i5DUML4DHEZcjaR1ExOxrX/7TFrS/b/AMChY0LPD+0+/5aGtTJzsqZyW
1qTxCrm/FvWc3UDnxtDRNeWc/epO5GY3gFfL+k5GyZNywfbKntbDpesMGbw9
9Or03PoHeEF31RY23/xGLRCfNlp7ZdkTpBKG87orlemORsuvp3XDwr4OAqSO
fJc3xIOk1qgktB+vIoMuy7NnTNdCKv8GmXUe6QlPcIJ+r2KmWRWIqum51uAE
5sgPITk1mQ8xGeuc3dnXy+M2Fr/baOpT5fNEaRmFN+BIZ6IrJ2ZaoaUCYmyN
sXGrCEhYBAjBhIeRvFvlNE8eA7jBmY+EaPIQSZVcgERLbpAHyHcrzg1UujLa
n97KqFwiVHK4iTxYqWSLAv0gtXFtuk689apH12LtGJAzEsoxn+TNnprhVdn7
2p+7q171mDP0C/L5h+7acXd9y6hTQQVoenMs5/X07E4gql0u9kvMuk6J98Be
5TCCHJMHRTEceIeuXoBpH4Tg+LOvHsC7nOO2iwYQjCy1R08XAkkPUCWIMTxN
n8/T4DdgmzKhKERIBeuqeQc14NuTZMbKHWrbY0X7lw4+4PACRyeX9AEx/hzV
/id7Je1Vp+ORJL55C8ztx5A2brHQ4SyCSDkntAlTDh2+NELcTMdE1acGIwOc
sPQZL92baL8SQhGM36FzfQWJa23If63rXNpZ9qSdE7ROp1hsoZHWZfycYLYm
iLOuCyYyHeaODjlEYMmqvuB0tL8xsUDJ/fZeusWPbpDLYohuj3WGxq0oXU0E
1FiujWGPCjOOq19xvRX0XA1aOQL3LgbRj57xw8aRYz8Nxwt+4VkV9PQ4+PSj
iYXHynsqBM4U9qadE3L8IJ9xnsiftVLBSrTa2HQ+gQaeABHCTsm+6jQbiOii
iKJkyEvtSVWmHAFA5DMUCg7Ix/dFBWf7wUmc2P9HZhHn3mOCBKTXdyzUC/yI
HIGJwO1azXRl0+hRZJXiLDdRFxfAmUwXI8oYSmNrFCMcS1JNvFdekeJHHRD9
8ked6LIHiC0KXeyL5ARCg3BiA5PdiTWl1YvnIqvH3ElKWe59u6+9Z14eXVGF
N/MF/hAKRO2pKJMpGFMWAyEfDluQPNwWXjs20IkZ5WrrKjk4rFQypdInFUZB
HWNaKnMVjd3n3Blzwj3oAZmW1Lzh4OjMLo8WdAVKeCrLfWU6gdArnwASTCmm
74gm3iSByKGq/y2PUkLEe+0Eu7fObBxhfxnzyPP0jEirdb5Ar93Naf117nvg
90waCgzTIHDwDUznJD1+jkcWKnNtLGOFHuyI6MKCan4Eb767JO7HhGxeBear
aFSUbGjAK88Kitev2cS6JXS9Y4xBHysy4u2NlwnVE6woNju3zXgG7on9HjYW
J1YGS5cSXrrrOMxpr43/TjynQOyRQvLSs9Est1PpuCgYCpvBPa/bpxSHSO84
MtOw8X/PR12fi+aATdATtjvevXNRQekuzPbC0fVsVuPJ3r0Nuk5Ii8frvoOT
cKkPeZDYa0+YWV0hU4Tknf/eDE0nEQChJe5w3o0azi6BBOFgGFb/Ws4j/AVq
+tuuhf/WfWfso2z+2DFyymnZwGJBcUqpVmMAGjmH5UW0HC8qsrGwL7zJJbfm
y4dNmIV2bPmqSrnbCpYBh56wqPI1nK7a+0pEAmlq3SzqeL4tyzLc6ZabS0S5
J4I+6EIRJMbrqC1ytxpFQ3067bIH7vTyn3YtiQvxLgKvw2PqXsJdLn73Yu6C
hBMFXkZn7bYDFswlDVGrkodF+opCug9qL5pIyBsmtOcqm4tDQoG1TiaoKT5g
On/XNFP93GtgU251wyQsirTCri273GilGJb3p5K2L4lHH4bTa4gCzJKtTNai
Wm3rLE9QjK7Vy7UChCTM0kdik0sYAl0defQcVLIbSun0S/yP3NemJz8orVPW
ufbqPVucvnzoMcTLk8Qhne9X3D63Xx+pEmKNNnn8hg2j/QcLHbf+6zNYlEzP
DxXwOmk0/sPhGA0uU8FNuUQdG3926P3kzNdoS39twG9qSkQK/1brwkHxP1zM
0pm4dIGT2vfoC9mcklw0TN58Bk64IJSft8xvtRF1taxzL55zzSWZNV0bWB9z
GGsafLxrc2eKnB7NUGu646oCPG9zb0FqISX3G3PT6BfF2zzB7ZIMyHSXJJen
6XVkCJ8+1b7mG61+bs49qUZf+KEp8Bh6zCnUlwBKbE6wKAwijouwMQM5NZPs
heVPKtl+U7nd8xbiPzUDZXeuiv/rkm/R8VCPRnig6HbmSC8cnkXb4/Q3BZm+
ghDuPnwJcPVLtPDGtA3aMUIKbii85bo3jWDAtRcwbsehLi50PcJj5LZD1ZWj
4tsSI3+3SpG/nK1R1AUCdb5ru1cF+SSnSUzZnc3cq/2jVzqaMuxqKtPkEE0x
GtrtmaXfN+afdaV2AtxfGuLMwwKW69TcLBRlVMQvB/PqpSGyJ1J9VUPNTop6
lcY0bsWCKEw4nQCOThy766c2xPVgyMEBM0zyAE45cYdk5Gh2+Cb7ISnncgMz
5c4FSyiVDQkrJdCaPMwUpLncH8/XIit79tpBTZnp1jYWYxA+6R43OtEFJCWs
hjQBFdS/EyVB+ltWZ4uZjpvg8J4aFIaJ4mbFr6xLeUcXQU934l8mJTrlTmej
rukwSbiHDQY92F3K9Qq2e+t8tMMif8vOC/Mi1IfS0BmdqTCrCsVWC07nwCGj
BzmyMsrVKD/c0CaDgYWIAPzLNDNLAgaS21sKs7SWzJpOe1TRm5LUmuLxdjXV
a/VPNqACqUZ+75JxO5n/orN3KNYUedpNe+JaPyjQJM1h3fuCCrnP/GxnR5oP
n1UGgoe5uGBnS92Ro44j0bxUKG6QxCHUlnUiShWFbNP205+ZQ9WrGX00KWMw
iamkp8aZ0WxW36V1AEmA1qGcU+caRXxlB48ypSPcTZZcRhNqGxYNh0RXxjVu
9fd07m5SByGIavfeEBbSSITBNz+KUXOt20cKmrwWZFEskGmudQJg4u+ZZYHs
nJReaZzcBsM44hzfgtG71+AYQU0BgD607jNEpjZto3K98tkudyHBKoUXF9gz
m8c0f4j9mrkvgqhpdWhMAkduvxHpto1ZJL24wq0NKHTuDclyv9evexCFtGTJ
uTDALKSVi4SJSFDofFzG7/ubVpOhOLjJBvz9PD+bWMl3xMLHzS16oKVYeI1t
ozywqFqr0GZvfcjqy0csqRTU2Q19bWo7ZG08nx5heUq/pwMk+jam5dBceSzX
jZf+VEVdpEMoEs8/h/b2JzmpRRClj96/tU7RrmJmFjkBJAdZLMKgIz05rrlu
KkS4kIn6+/dK7QNkdKG8q1LwYVxHGePcMQ1l6cyH7Qeo08QnV3uN2nsbuIIG
MPC3RxxpQOlWgD/Xr00Ebf4s61eYTCaRTI4YAmqJGLqq1BaeEvkF0zh/HHfV
e57CIHtVYyJLEqWQphuvqmvHI/7eZ4WAmZ5H1XA8Fot6H3bXUqPyDpnIq7H4
51FOLxuGEtn5UcN+yNYvYthbSUDC0fcQkT7DEyQKP7Crnix4VVNQLwAvRjV6
JERu1WjNrQjLVBh9fMylb8AvvIMNkn5DJTzGzDaDTwqBIVzDNasIsZCmWFnp
ld3uc3sFjXf2DMnAxBICkWztxj0YcRM4jH8s7qa9aJozTS5w8g4vLyxgNDx2
Kg6Mrb0G4K4BT/kaNVAxyoxXcFA0coWo5SpXqzzYm5n5OIxBDHQufqElOnfN
JxOfy7vPjD5MNfL7zeQ2tgB/t0TP22qPdRiFRiQ6CmNTV9HtkdKwCbecBixo
5gNgvswcsrGVJrywZ8479YxemazNvy+vRErFcCoNGgU+vQlJk3pIHSA/igVt
NddLw8Bql/akw2ci9fSJ9zb4WxYRGBXJESeTQZDr5vqWlYRg5HvpFszeJHpp
PAkIuPO2CjbGI+p6FaVifQpdA93Q47aX89ADwosbq31uQbwsntMrLsUusGW7
Sw3EAXvmqau8koHgMvdqDrsWJ56ehjt/Peb9ueLbeQHm2HAszpaKTMEYkem3
Ik4i/GaxmgnJ+7VCzm4x9tYjxQyIaxon0p0JQO7jg5ouu45wSXXzmmGj0JVL
5R96tphcNWt5/3OFHUywWbmIeJwANEhEsKhmu8nrO9PwnTRPIvhgGZ8leDI5
JG+ESSfo5Ty+WF3IC8E3/rqCTeqa/s01uatwW0bqs8gsTUdiiZw08xk/VOir
Zj+iAKbHlKL8kl42olM+pUHS/Aij3GmoThcSs2ds2OOxNQcKGZwoC+BzIoQg
w42394eYkbPmL7XCBiByXbGI0KATnOrYOGjZ/thAm+kec+MkPjwcSLvYnaEc
IHRQetyU6ztW3axCsNRnmGRogjMb37h3pGXz5wHfkm0Hdk3Kz+iiv1SO5ILh
GJcNK9R4v9g9zDmPMXKge5rWFcdQQmC07K1VAPvZMl8Mgd89TglubaXy8dt7
pbCFQn4fhoV8/X3AFAtK+swyFUt3YkeGwZ2cKAUYyUqSeR6TI4IS3LrKguSe
qT4mQHIObbrD4ASvAwwMlw3G3iAS4pTdU9toiTZuiRkJy3GtMFieMVk2Rp2/
QXsznycuue+/AXDwSaDj0vWvuKLvn1rv4wks4si0l1a2LhMav1Ojm15hr5LG
epcTqxwUttuE1ucbgyhv3aNkAlVw3M7naDrkyghD2uYtl2dT75nHtcEQIQTA
sHpR/XBkv2SkbZqUF7iRMg6sgHXc94CrCPT3A+k8Mea8KKYfxoZjGcEufCaT
y/B56UzVNjAPd0B0WgNE89Ok6hMy+Uo7+4HHr+weTMVXrcdwKf5KwadXe6M2
25FFTTT58I6JJpmy4ajOhykQhR0OlhzwN18z1MpoPMNUHuZdp7cUpOAvm5NS
by0MB8OkDI9A1qIotuEcMxM1o2/QChtuv6ZIKXz4zaN0RtGBrroQ5Jg6S0xJ
g9uvrKn4eaRTWv2imbQQH22OYefVTAGPGhfmE8Sevw+T1mSCkQRHadfmd8Wm
yFJvTVDqjcCQ54Ebo3xR0kVM5nlo7NFO3EADm6SMv65z3xNSsDHX4rwKhkqx
BZdvR4APMv/KpkKVZraZf66S70TNkB/LsHnHQJ61L7wP9aMIArNd4SUOQ/KO
pUXCbYlYxS5uWdsoN7KtdnFTHVk3qIDbEVp5pSg0Gt3eB+PKB0g+sYLx1Hk6
lrhTjNNK6azcxcK78IQLstiBdz7TaWSE9I8l9ydXM1bH3y7znD37GbsPcZro
6elbcqvS/pjMBh+J1YPwRHm0rwWwpm4qYlg3qyAmtub/KprE4nKfdSsYU6PH
CPOhuT4Tmuwq3W6/qCLXLeDl6qkspbtlHXbopbS1OK0vHRGcpI3l1uq2QYLe
BBdes+vY4F13hLM2J91t6vpd7XjJXW8yv7PbbnoWhFW7DGgVFwzN5nA+JPvw
793+gUwaqZGNrJMaR4TK41MlFF2fVdWB3jYOy30gHjNNoXzlY434AlxTbAqm
AsQ0KHqdr/VmeKU5TSeTjwXxkpQQAcPR1mPoBNbbyFEpG1YjWVFGo1c01pc5
NFZ76LxbFowY17XragprlccTVO8AjzVQkYkAUlF1KTqV0nRIvG9pP2p92EAz
/d13nq3XUhCmqBXUmn29X6z+Kk/4H1zKCP9gVYRrItZrylUea0L4u1il3xWO
nLwKwbO/cgsn2t7zcyJMSDQe3aWazbxIfZB6K20mFvZRjTuKecV8fMQqw8EK
u8BhItNgd/iwkGBIH77g0UThXs55W7Gyb1aJ94nLOOZ3vrLBA2urrdJnc0mX
El3vbqiY7Eud78Et9OEGQm/9gDsEt8uBBLIpKh33A2TUVUN3p/FsoBpHf7zi
Fnj59ERc09kwXYFMwy1Qt//G20DlDhJ5UvUitoJz9lMLu5smoL+5U2E80DU+
mGXmLQhdLvDQ4tFlhMbVUNDMz6xeiX0rhwoFDJ+jlX3f10cv5e7TCydY97og
0AO8iH7vtOwGqVqtSaxEn5ylJwI8PStBBL9oqtHkFjeHtfjsRPl23MtnzRMv
9M9XXEqJEdh84V8cGuCIyjUfcgYmV5M0JMVG7cIb9bjsfudbWYj/U8Si4QOW
OKy45mQbwTpITbTO5p/0Dkm6uX4IBt7T6M+8X8hAZq19M38TwOkj7DezqQAj
M00CKh6pX9lF75c142QoGYjQPoZwFXebhXBDY9g6g3/jFQK/Ai26xPXe31ZO
5rbIwr7EErVdf1X5Ac9FSg09uB2Kh1zsYVxbPga5z5hsaRqdlzxs+F/j/9RI
8/Mupx0EJyc/TiUFRpxTT+4JGZLO6oVYDjTQVCM+Ey8cID7dIbiNqt47oJbC
aEdFXXyCRL9H8hTFh8Iv+bgV/koJT6mW439sHSM50QmntP553a4O+hmDiu+y
87B830JwfTo7FGNFoGxmg/Ku01hwGrVIs53jE7IBzIz0GmkxL9uuQH1ln+/r
kAMk5+3IVzwWEzTt8AnkhDOoTMUcfYhNRW11bKpPfhV2nq2CdcFlbvawdZwm
iKEdNzy+pCNuLlkJTNXOIjwYd8kY9/YqW9g6thevXSE6lYO+tPOdDECvHGfI
P8HvPz3ykZyh0ra+vlwCbIV8A4cnRkqqB6a0VAkzXsQx12/rfgeXy89X9CAg
tXEPraG2mqx3wfxmksUa7AFsr3Gb67Gljsq9ES/RWbASuIc3TAMduYR5aoes
efUAg9VzEaowoiiCgZXZL9R8tvO50q7IaLofybigmPOeCk9o7ajai9qXaYfg
bbGWgYTB07NenKBRceqD9zLLQ6J6vcAfH9sxwHmRll/9qb6MOShuXyl90mbj
OXryv9c28Fabs4beViMc5PnYTjzdzKd2cMi3eNa01Yy+zBporb1g9omtdXab
i+PeBhFCewHOinhFhwPHZBTMTU7rfmaDzDS7SYGXBhCQ5jXu8Z78jeOqQpos
a9mlMvprqPw1UkZT7teILqY7MTeeY/g+1YPszdswnCwTza4jc1tNw5dzRCe9
XcyBl6/YP9Ru6d4pVvsOdZjrHutSxNZmUa8jo3mQVojQIMp3xkBc+o4fQZxL
u8HKWtbkNTu6AT368/JeDUTqsy3+OEhnMVY1BQu9i0CGcijQxajgrUb6WJ+l
/frFz+C5wdYqdac9P+qwp3w+13hzQn2A7jOKVq7yCCchPSiGSCP+nYKvebvV
MTGZKz5xGSTxrgOmZUtPJ4vEAsikn8EXbkfLj+hcjyLUkaL8DfpBM1vfUc0y
gSewmmaI0xEy9X09Ur8RGAe86lN9q5lhoTy/spcoq6Ng9YqCUmE6qBFczH75
EJo7DxrMVU3aQ2kXlOP2An1ywY6QjPx5xc6UwBdiTljkbXhRc8XKjLoM8rPg
cbkdTT0cibOh3OI78IrSkdIoplBcBpme/Z4leC45JpAkzZum57+G8wlN60wc
tsyqu4ah5BirI121c57cKxdnRs31e+axeATF4RHEYyufdG2kBAg2hp6AAqJg
CWneXbxIRC133vRy9DJlIOh6PfNFYGCcpkqBDWdDlNDSJAzYSnAJROwnCjK6
eczlLM/mkbiWAXP1p1ZAXtvum54fvFgj0Ntv8noXDlqSntSRdJ3aT595DAf7
ZJnItlwWJJrdqy6ljBCmxCRmlm2cTjbWXLayq2/ZGrNjnr1H5AjLrEVXGC2R
eLbQ+h4U/ECEgkfUYacixFVN7iBf3U/rh2VxKB3CXNW3c0+jEaPH2zB5Abmy
a/ifjFKA1NG7ITL5bAelfHRsN3tf9CqET/3bu/3YOpLC3myl9PYub0BBQuGE
tSZ9N/Tppr8uv2qZw33VBjeIhlNP7ul2MZGsPy/zVeObWP1z2ux2Met5hFxL
6Z3ZYFNdR7Bptahu9cffLYqETumf/Q/SCdxXDp4lVey4zjk7MjhQHrrlrJlO
oIAK9kcU/GumAG5wzaVZyXFOXSZQf2DUYeTWlMbEliYx/0PUih0COeUb5OX4
k8J4dVkYLR4a9LO5BQQDMCoonAxq8nOP+Yy+urRoifMiGSbt3Gg2uozDOJ+B
+EEpRb9hzJ0ideWova5JZgBg7GzkYa+wDCg9fDu1qjU8TBgSWneB3HnL/bWl
xvhMPgoR0l0q5prV5RrsH5xFxmDWXuJ9mBs13MnJu6Gl4bllcyMw3uiayZUP
3L2gw4Xy1QW/DMfOVNjoFCIZ0iM6sPUIrK2VH2W/0dZL7wqaPw/o3o/dTPfl
ZeoFcFzajHzBmb0vnY7dnHIfWXPUrx94HynHCoAs6YNrbvYKR+tisiAgg04O
XRYV2eu0tYJL5plqJO2Yyb7iBEPE/X194VfO2g6IpdOZ57ZbJaiIlVmZOFuD
0aWDNHs4s8nY3tY85KEGwg89sImXBjdUAXNLpKE1+CeOV9YfXHhgLebRLhfh
N+fiGIALWequj+1Fcxx5q3/fJQvvYLzMs3aM9Cu/jkjeuwuvWEsMXhK3D6Jw
EP2HkJH5X1wJ8dGchhPlCRYYKkpLa0loc5a1bJH1XwovNpYU0WfGRLozU5wD
ZCSgRNBQAk0BmdN+XxDrobyjRB1tPkGZcZ32gsaYD7cbXYNsqgiDt9lQe34h
sXqzE3lsU8G5rmuxCYGq/AOCKmIvBDvbaDrejGHNa57sAPu+vvrzscYwj4IK
J4Rkh5U8rDpTmXIL6jjIsCbgrqXOi2kM/k90Mp9iXZz3McLngSqjDhoVU956
YdlW8fzMr6iHW6m+kSssIwKSq1jmaoSkWuZOKOSn0esD9ZQnxf9Dy05jjD9e
5TeVa5KOCLffZ50YRGSozop1mUgTo1e5tJ9mRulDSLCorn471B5H4Q1TN0mW
u9MmZLn30ncGdv7O+X0uAdH95/1PiSsaoP02eznOMqMoEIfgROySIKgvNAns
YyumUjqa4vtpfTlbpw6ZZGGHpMnsb4Fp6iKxwNZqeGhI+JTn2Vt6fJWSt45Q
GWOHVECut/wsWkWpHqlm+5E5ta8zcqXYliqDTS5O2jdCPj4WqjYe73ug8WdX
toHUuqhVEhEMPC6sh3sUN7nw+lRgy4lkdMrCeg6nFFE2PyIJvVytR/br1iZ1
dCsSBAa+4aNQ66jA8enX7lv2BEzumja7PcF9WyrxgcNs/khCZlhXh8tbKbFg
cW73lXYG0CEXGW9MI+wYFqA9VUEiyfifMTklEE78unQgGoR4TO1UIrwipQEd
SWp8UYlX0LhUweVFq2+t6zywC+lgMHZTqjO0ysfW/p+PuryKi/4X8HvFsQ4+
B2TK96lYBU6Qte18j+U01iFEnZdI+42uBzCpSD17YFkp8bVsA1Zq0ZHj07hm
039UeP+VSyNhYhT5Ap3sRmbz6ZDYY9Cq1vhiNTH/0bsV1hXZ/+tN8IR9I4Zv
4wNjGKia1VW5o0OQVa1LdHQ9f6uJ07MLFEt4xtnBBnIXRniKfPI8mlPA1NKi
ksHDNF+REKoHuHv8kdHSKJcpUpiFHt91s2YKrMfS81EFNVXQ/038uT6rq3jI
KN1kJ2khY2Hwts3JK9awaCyKzd8752I3oBZIYitAwjcW0X4eu7tc4QC3Upwh
gOGpwwZ9Pucx2RlPKLBw1haF5wjVcntZFLF5Mr1DYtYlmgn9pe+owGZhke+S
CGsWKUWdwMkVBhJJzafVYE+wyciuAhLjhud+it9i2KIjw9bi/pJQH+XGLc/f
blf56uCv3ya5edCS42wGlpQFddCd+OhUYUutNBZO770KRVaVDDLTqBIZypLz
nxYakntgBX7IDIgzQReAsaaXY0RIiBLJ72bSD4BhWeNRKC3aCr/jVO/y9Ah/
7J3ADEn6oV4+FiiDRju/ef0adZmEm/pQrvVjJNMFBY4ueO7smCFkm41O9bef
ef3m2ILpYte6Jwqkno7jTE8Q/Ltb5UGRqnjOYy5BKVI1XMuQxST2Da2hg1mZ
eccWAWsGTZEiRbVRENPk0ixRQGYx4/lLuTA0ISD9TMJZnKK6JRn6IR7HQKBt
OsTNsHjx6dCxQ3U6M+funcmF4TqYpiS5JesprTeMQ4OZnt9t8tuIUNLbE/mg
7DrPJWF31qEehTVfz0k5Jd6ehKgOm3+E4zGr7ZOWzapU3efK7HtDMwtjiffM
ebQ21hLLj9Ws7wqb8MjkDmXghGB5x0FjbeckzF+tpZp/euxjvfX1TNm5MD77
Gf9WMCLf9GaNGZEmY3GjaH7oviTRhZblkuEFzYjiXAHeQrSZGeU2YuqOcw0z
5Kl4vz3SzlSAelCVT0UKQoK9yd+/jKPRVNtlzTm/w3GVILl8sAStWbTROInn
UgToJqZelvemaovHXQK640E0WjUaf8f6y1fJLjPOJtUfd1T/HRIOrkc8anDa
FO7btKA/Rr5wQjDPnZFZwbjuZmIO66KFxB5dtSKByTm7VgZ29P/CiLU9Fj/c
bfFCC3ikxdwbBt7+a3Ya2gy5pAAS/lw5jLQgArFYP6TXK5IAE4tScDHW/tJH
JEsuFShcSQyucerhLEokueqWWExhePKJErzvYHG7locstq7MJkvKkxvt1jAA
5T2V1okH9ibtMNcFr43nbrwrz1+mFeqt2QB7kh9QVMRB+DYk08u6wbufybR5
k2JCEVU5+3yiaH4wLEsXX2D6F96Zz9j0D39y0bZjh+L8pKYS6akzOY8Z9Z5X
VE705/Bz9lI0HTf9YH16CxSzjQx+fFRr8CgVr/CZXPJt+u7USmnBTmf+EGcv
/p0nEK3c0+LMVafP/ocbs+o3C/jDmDnMTOx6HlTscnAjVjFRpovH/YndtwV3
vuWnsMKgDRZqdfn2HjdLHKDDCvxXpw/43qWCM+HD8hmssIKkl9CoOhyKO0E2
tP4Y9maQ4chrqJcVviPcu3V5ZaQeorzSBdl0YU1kgQZT37atkIGr/LV5rtQd
p8w/sR06zOdfs0gzCMluYLn6YCj2bqhtCNn6nNIOkl44YWkp/BpAjw+hlDFO
qQ3+ogjzienhCzVbSfocnuyzREWG/29xOKl0Uh9DwIaqblq9TM02vDvtxsij
WHGGCT3J+9K1kx4nZYcnwb3ZY7H8xKnQA+BHLPmO8yrGIS3LHhpowJjutaiF
UZwS8AhUtI+jTobIfdsSdK3QvLcuNKXU4X4lotFLOomzSAfWlaw+B/TIMklx
V7SOjJ8xR/zE4RR0l83mu4UAcK6z+BuT+3pvguSneLfQC8yRTBR2Ws5eOTHd
naC5e848V5UuUfhj9sHcxoCDMANo7AnHCqdojIFFSNwKzQcEF19RWiqOX0hs
hQFNmDZLJCXc1vyS1ERivk5a8wTdJ/8I1y+oY3Xuvgz7J36JQyH9BonQHRe3
ZOvmt2N8+uiRkdTHctYimILCfN+MRLqNQuU/yp13K4AH5Yl1dL7XDxHW527R
kdKGszzGt/uezRkakYS8u6ns8KIjdBmYDgn0Gs8EAkxgLsGoH5ZjOFtRgSX6
VI5tpljir3el/SBJzoyY/NNmxgcIRcKZr2wqbgMQfJDFgVICNOVDLzLktbMW
ORZUlAeQq6rhDe+oIzTDeo0Md7nBINKj+hnA17i6WWhvGeirfMTjyLNMtFgA
T5Q3bgdoC4SphOTpL0Nf9BxUmMzXyFCNc8JAU/rDVHsKYRQxDuj9Fq5RdxfN
HhHGgppaIIxQ60jYg3JJFJHPmSljtzNKIoxWu+ZSbF2NxXOu09SjLNPyG1u2
T5zbD8OqmH9DELWdhYWFJ/0SY+4BfIFK6A4MJ90NTFIq5kqUA/SrM2W6Y29s
1fTK04SSR6G38uOtOP7gUNsBFVImzlA4pzoRNhtmDoipUn9lOhca0soHdrTI
Fr9qjX5i82qDYH4ILGzTmlItfKABHD6BorSwTUkxnWxykdOD6TZdpEGnwMdV
czEnW4gmFS5F11hLHNN5XwyvEIjAuSBk8VP9rOI+Vn/M1pvBRhZIQP2f7j3M
ptc8K04dAnS4vtaBEEij+iVCx5dO0fR/IETjmFp7EsWFal5fYr/csNBf7Ey4
Cv/dX2A+hr2GMa6NtFYeu3zysiIIffguvgDYMtgeWwAa+LrLHyqK3M7oyIxu
AoSPL+F/J0WpF3fXpNJ3PvlmMWE8w6bZTfp1wY4D3mwxd+Foz6tewOz74e8N
t/kXhOpeuU7HPueXjgQgUApIJ8YYlXXUxmdavuITLSuCJUZEWfonIss/WPJa
uv9pDSKIeW3UWmZa6hhX3XBwXYl/VkiFVoMh0DkX+WrjOlbTz7vSUF4Y19SI
6TF8SECGL16fpxFjhWwnRRa6dVk9bGlaU39PhvlYygchKfQANFRYQKFVCIjH
b43MDUaRZSvJdV2I11AJ1kSrmZxiPY5IxjPrfJoedj8i5rtvpz3XMPeWA1hy
hW/R2h+Igy4xM1MBwr5SOXjEvjF4OwAOMCng9L7vHXnwXYL2bG7ZweI5KaOI
uPnEwOw8J7QG9tZjLvIZd5evQpnFUH32a4U1H+2ZprZqhqWZTnMLqD8tjVsq
DgYWkqm8TN7JISmgnCJ56l8T9KcI9BZn94/jrfmOEafa3FG5G1ca5xkd2JGm
vDYsWG6G/qQp14s+75lUZf2DG867GVmWFS9mRX+6KPy2oPpXHy4+bvn+rUTP
WxjYq67RUdq8n+gpW2Y+TdMaXO91T1WXj2/u3XqdRcjLyEE78e54nWmI/qD4
doDdxf7W5JL7dSdi7+duxB0O65YKm0p9c/ZG6PQEpMAk4NLUCc7NteDUci69
Q1/X2jntAwV6icIWGaUYLbuLrfRGDWG8CZlp9J1h2afP0wnQkg9dgQ2zcFin
CT/k8oBy9NiZeuSQhzWQqVSMiWLM0V/suh4D27O6neJjeVdci4k6rAEnarAW
UDqnLOnj/7qs5hFEozgdFDjBuBIwAJZ5ooY69sQk7vm3xylgdYwqV/CiWdfL
1qA22y52b1z5D3xGlC92QRXdFTNDPoxNCMipOG1B/QbLhlKGXQ7RCgsi0qx/
3+y43qFnNGLUlDOTiMpYu7UE99mVYYbhrFr0qSa1IpISZDZ8EmWPFid0f4Cu
Js1RKuhC4IYAWci4tDfwv6WYSvhtnu/2J2mE8dCFrK14OCGxngPYyZBvYlFb
eAThezdNU9NlY9a0T4NAEXgmVRxIkOsCRYZCCiBPzTRtt6KdN7XOUtn/wCBP
dn78HcduwJnhGXxTDAtkGA/s+eW69LPTVYkfAgd+E+AHLHKnkag8tEnXHkit
G77af2E2C2odj10Z4y+TxulMhawenCDRMUcocAk1aOWdL4vv5pwjaZnJjvVk
h9Syde9KW8+IJoyJ0PzaZorqXsHE96mGUWXLqMrwgnrEvWVF9AICLnVs0fya
04eyUTyDpVbb1h+GkRR/ehYJtwPpB0XnEt6H3cY3+SxQKVgUNBslDUFe67OF
o9jQP95EK+GJ5GWnNiObWsh9MAIaoBD9ET7XkK455P++G6KNnAYV00/nr2eM
KgPlqyv/0fsRlJRFTQmRlCsNfHJSdx5JRxkwPQYth7oeTFABqKiZ30qXRa8Y
WhnoZTJuBb1c3xqmAoAnK33Lgo4SgURBMA0PiuF+1Fb0Tufu0NAEYq/gflmd
79TrNqgdMxhMW7i2nR191yVD91xJB0S9h6m6NM/uW/xOgcO0Zi8mZIEzk80p
knfJPyIrdYuuJqbAIx/MpJBl46cojT3ZBk+4Cau+9L67DPK96lqBcJGmVXOF
ZpBFocnm+4UDnTg+x67mDwKGGfPRCWx2yx09BnAKK0B59Sur9myeQgQXrTfe
XZg03lZ65BMEZN2WGPGUBlg8tI1Io2oUwlMhEshoHfM4HDyxjgfUco6iIeWP
1v6ml4+nDHxYc3nm1Hl1i3JQTCSlqQRiSeipa/C43TE62pGhiqaBebJwgU4J
WkUoxZ4v/McreqFDreDyWwZYtQLkMsaln2NC/U9sq+ytat5tfNMk01hyj7/9
fLS5Mpydg/1bpJDr7QVGoP2B0y8h6ItM4zaRZ4tCNPti7EaPWNhh8626uaH3
UAKg7YbGg5Ez929XwMDNDnGIh75+v1QuQ1w4iKx536doUSKNMJv4DbgzW3Z/
sjeth5c1HVPJSmlZPirVshH7D0IkqnpT2IGrIVgOGAxR7AeM8w+rDITibIdf
8HBY3cgAfFWZz8tmEy9LgdPm1HJPE5rRDqat3qpScYm/0HbDNI1hVh669tBm
BC1cAnBgeD9foEdqlruyH53aDYAwm4xv4y64EMo+u4gdTazXhGf56kj0dn8v
1W+T/Dcz33ZJipxVNbuQy6lDjBUCZ+kk6WpZOgiqOYnhw+JujsBIomZb40uk
07GM2dG53A9Dfw/7wmqUuUjU1R053MgzR457BG3nrLH1Vy6yKjIGjPYw2dQb
48dxIFEbGKci4Hlr295O9fAClcWHqm7U7xLDOmKSFZld37G0o09dJQy6X5TG
pSIYw6q3jvbQLIFMdDnjLU49HdGRT9b3/z4FU3s+jaHrsGurDM1RJMxpv5+x
nojZl0TZag332ukzr7/T4QCTg6OLvMLCffnW9v5IWyfo+yW9pH/nt4utiazT
DKpXoyulOO3un6nXxTB2e6GrscznwRO6YDgGm8anvw3vu1VE6CEUMUirLNgP
x0Pb1sEapA3tnu8Q6pT910Rs9WchMCTBRVrFJzC0ARAthJ+3K4mmLtbMUu19
4+YC3wiCI+5fdKSgqvn55zxcVERIhYcHAB8BP2jyCSRKazIvqQJc3gUvjzaA
xZUX4HTi4MKBCPZBm4MQef8lVcV2K03z+G8sIdmQDBGLgQA4W0GOISp9rLoe
ZLn4PB+9oP84jS941g8nitVuYdgiDrWrDbAjg2iS3ts8Oj4RB1HSiWmcKl9X
XJTs8OIXJePBEkZ0cWA7uwrFW6Cp6GypzlSnp2TGl9t2gYudVnTnOAxNxkFe
VwUkI/6nkmpvOM81x0s0U4LEJO93k1vpAIs1RMrlLiQs9nxIUhP763+IooVl
etui17M2Typ6xcbKxKgT3FyI/55TGx59YtJ1P6M9IHZZqj09OHOpJoW2cfTG
QBcS7PfMVP5shhaXa+JaD/4yctHMCEgo/kwmgrPQDldOQQDRI3Dr0QAL9NTb
REL7T5YnEsNVRseBaMSHjJ7MCQns5eGV17lIzf9XI6DvPgzhL3OxM4UChqOv
rkitRmtsnSJFpAoqJPSngqIiHHKe7SuG1X9ERxtEjkZVxytkHoGAdW8MRaKL
mzfOYpvwZW4nmw6TU4kglFqOfJFpOu/wOmGmse7lgEYapn/CTcGK0NGxB5jE
f4SMBOUYhEHMbqNh7U/xgE65L0AMbJR16ww1PVbHTbDokhJXtRSlW69w0FaO
iKfDwAH/CJPb3G74hQSzhpy+fRHz6MnOhsVBrXRHYuPXoFipeK7lM09s7Uiu
5GygGIDoIM834tLQm4O5Pp/Yfwsn3cMhL/l4I1ZC6WYBIy8cOK3CJ9JWcVx/
yhCXyGDv2slIpfZ+PbPK9TpdHTykDDEtHhry4XIt5QUFDoXBLIEYPWPO1VKh
WsFv0EEzKU3ONUpVLzf7b2yKQHlASgukqw6EuuWsVVZtl7hvDjvpxJie9Qhu
iAtDWjVCbvTwfMm/EYVgXp21bK0tpO7Ki4Iu422Bxz1q9orMd2aqeCK1SQIH
owe23xOB5B6v4mMiUays8fy68U4TLPXXmA58diYnUK8dfSU1ZKfftsVPtq7w
PMbA/XLj1zeI7LX+RNqRgUX+qjDqQs0e3YBOSoxx3pj7hGQaGm4ymBPdGOjM
OBfbDV6onta1s4pG0XsuzrkiTjmEORj3MuQIRrUiw3+MFTUE/BIcmOrJZC5t
5CcE6tQ1U/jIqok3BPwTMfw3bk0RRTeK0wNk4Eua9BLxjgV0J99IWrkum3jw
hkRIIl8voZ/piT9nsPw2afp8ZIubb3UT0k25HoMU7T0byTVvcXea5naNHjoo
Q0MkuouqQt12fxTHf/+/dBVj4CL90Ec6q1v/GVC4TiLg7782+iP7zzYTHK6t
YE0x3eO45c9RAhuOwbziOJVWFZul/40o9B0SeTlYdS+xrCs3uD1cuF75xiXv
Ra5mC18mDiuk6kqA5feFKcvQmIwAdQ3awoqT+/cRS4nd3q50I2SJUQUEIzNc
oQHANroXrSuMuFz6MFWXp9F3VVaW5vjMoL2i2oAS+zCDfkbTL0rVv/aAumMl
zuxUw/+VrBl7FH3AXUUzJQlkTWvg6pM1utXsPU7rBBfIyqr/Q2ZKcnHHGOYd
zRM5xFTI1PStVhADANOTXUHJgrTZmLuo3jjMbE1x704dJNzCBEjEm+DFChyp
AlYHm1FanhD3lbjpnjgcjBw+G+vckWNI9swib3E7v/zHjXnQuQfe/Vs16d5N
J/D84qTGR/qemtpYX8qUWw00+uEyFijVNXljg1IqnuxBPB5GKJKWN50zRz7u
OG9SeaGOFRihAvKLFTGKbS/xFNa5EgtrrrKa3470cAm06qLKbiBxSctYkb4z
5aRqIHht0hSeynhE6zAT9CCzcK8h6+vg7cq5IdVi/i/yqqZXtJiukX2BXTsg
E/Y39g9QGuBBHec6emIl7ENQ7qdmEp5V5eih+7Bw2eFY87JGL++o6Lbrq5JA
p0Ge5n2A3fVA21x94ETDitigjSzPycSuelUHW6gKmO2/DW6qmQtWf2zIDSvJ
pQMgrMDXIfredtjwIxy740peJdsaeDulxGgv462najaUQptNQLWh+pA+ZUmS
veSGXazTZ3JJXQR5FEjNVPHWUJ6LcxlXlUy0asmsGptWQzLK3A2q9ahYaSD+
vFTxnax3ttX3IfPGX/Rue/Dlb4+A0ICva02Oi0uOk7H1VfR/km+yVf7W7Qs5
QgNdAqGw+Xkr2bustW1IpgVq1EpsqiDNx4U6VL9Y+3nu54/7j7p8+JDQWQyv
4nR8hOCwXlVpfmHqnpMWXqb4qdw2BA3G36qKa9VRCYcDapRNOPjqwY1lRiaZ
OedYIQGkb4477sOxpqdDAUIzNWheFNVKM2CtB9yX9aaYDtVqBqIrznW9lnhW
fQRrw1w7KbpVHC8m5E3b7tLUDguDjVEtklEkK56/MvanY8bj/w8qIw9Ol3ai
Mh1M1meJMcfaakrpuXZ8O0HZvJeAMfAsrtWyuJMw1o4VHTqbPwJ+0zJVsMGg
7hNdnStl84ievtkKUDXCA7DCU8m/hXODdErI8tdIoq9+rDHQWpaGONgZehRm
9j5o/4M7TGPrZ7vfwODVf52vwgtRCoFOu1nBbCbD91ZYvmGDVLwz8GVcwage
ahXX1o9hbeXFJ1ZZn65TehYb2D8fFrX1zoyLG3fQZ2rtB1VmMwqrJZlKqrrS
Y057FDqadWyclR2TcHgIPJ7E6rdy2/5HlyUbHP0x7afmJeL5y5+8QhYA88CX
COKIU4mRZ39gT+AHv7cBOWF4VP5AvVKXGrCZHu5v5aBPHx6cayyfAnNSR/Ld
bial4Qwd7XgZ/LiLe22+oRQRgClULcyajZ6njUM5FBbjlDO1ltdU3/luLwKR
kMMsnB+gn2bPih2Vck8Tcmz0MEFE7FOtRp0bofimvq9SEZE4UpKdHvgDfpzD
SKDnSyGOYxvSt+Gd1D3/QqOFsq03hnTv1w8oo1z3HmQY4RvakX3xFyoTUgIw
ZXd8aGZPHwdSzUkK+WaLvl5qLyNW6nqRnjzMk1osbSkOhU2tysj1AxXneFhL
/HKFGVkTXe16DtJBuCb4tybXCpH3GHBDimr0fqo4/8g1s7mB22ZEFNT+otds
a8Uii0qvK7wLbFabXbwcodUjT5X1ncUs16XresJAPv7xJUs4q0aaC2Ppr+mE
gyDl1JUhXH9b35pd+3Rn3kX5jqG7Sh2dewkBrhEzVbegkEEBWaUSBJdzcYpb
2cRTSzyTXIpFvQQjI2qD1J/XdlCNjtFQUkVUbvXFeFQlsVkLv3f8LzbFnucu
6PzC8Jr6aoDmjo2bajke1R3ckM9lMe3sqfgGSCn5d2p0qZoJyXUuLBiPFhk3
sr6oR4F6OfdMuggCokYoUJOrg9MTqhOZb3J3iNGA3C3yWBcB3NApj/xKnlKW
WuhwC65AaVBZX9J54MgCOg2MqhRDHYzRJvPpm/i9VJmwMAYzHckBk9q9lptZ
Ku4JH01WQb9JCm0OdNLTNOhqFNvrFsa48RwrGxzAAMnipq6cnahgQ91ful8A
/rLX+JIC9EufYQdTPXhjNJFwxj3KnW2mVev1SFfhN55hj/YlrcFqXChaQvCW
LXmiArAOvofymkZHPaStsX+SWQlSoxUl6q/h/e4QSkMRI7vtaI3ZsTOG0Z3U
jojBefYpqcBdcfJZj5w3KmNLr7TcJWq9387QaCB6IMxn7CZ2MAw855RUcAFm
QCuywaM9WSYF7gevkmEN7/DdQeaGxlrM2tYzLLOssO+V4+5dYcVRAlE8NiW8
qd7Gtgbra8FS+nSoDxXj5bPVEM9vcVjfIa3MbAbNGveGNYoTwSqzYsyNGbq+
jq1Ajr7eD0x4DfKjOSZYe6LcK6KZz3ccY5dvMwe99I5N+JrsfabZF0yLHMa9
F47uHKQoCAEbE5A0EEMRq1YEWKzMbkREv0haiiDaHbOqdfNyZucg88pS0Uhq
A49tbytiZyUFKboc8sdQOr1e8ne2fFgIzGopnjX6ZjE8cz9CL0BIqyziPrPY
Ae9apAwSI8uACxfjLzDEDTkh4RQ3DsLLnuRBE1EgYvt+xo8Eg/GmlAkYDIln
FvbBV6osL0NsaMgJ1/dWMvvGzrt4zkva7WicZ0v6Qcfj2OCeghxGan/STD7d
bQtQqZyWuPbDr+h9Steidq2OMh6QM39EV3e186rYZFmeihLlNiKRjvMzXcO8
HEBHjO+1Ki9CikKmd9c22ekH+ilNKarYdwXG3EJAOeJBJiP/CIpxGZf6Yke3
O4I/16oLJZ2W6/3hI7W4pOoV3YijmAWWyJYWD8Fbx55eOGGiDl5mEUVPSZgI
c8+UvL/3IFR1bLwFRK4EQgH6LwXu8UbbxjVIyyvLnPNP9b80kAG9CGbnRIW7
DtfzvfrtP4fzmBs8rrd4WezMunp/GS6mLCfmq2xCEgDzdL7hLB0ozUZwKKa3
1sIOTmjVmqxe3MeysaG4y9v5TZjR3n54ijYakIdCGJlJ4okNBI7GI4dOoJFe
jjMMlhtGqN58QbaFcAsf+j2sHQr/SsFloiornFUuaoGmAS8HwtJ1PlubpWS8
EVI+ocrzY6o1SdAPia2EqvBhFRPt2PzK+428DA4HiJNquUINrVHC223LAzab
GJAIybi9tUD2FC3SKLMdlPspXVFKk7Zfo6CVvhG9ZyovzyvqYTbsq8sxxw0i
ey80vWtaTNjVSNnzCCKX53k8etXfr9xGnqEbGs8eSYFUZBkIOV5JqTsPgT/H
FXvdY0N8q14TGOrQW3KaXT06I5umeke1J8YtZqIOIRSbRjov2gqi6ZQUL2AN
wtlQT9DRJ5b+0GL9jiBhINo3nkvXnT32v5BPaatBVCjSoLGBhVL1q/h3vPHc
j3TmB8tSGdy3Y8/1PCo7JWwFrj8HOjz5GpPpFIowMHMrzQd1HgXrbq5f6Sm4
5ozmNdg0YH43me06tF9B40PJRli6rf6s0xITVeVWgdqj24hjLgdrJ1NXmzfL
FRpWwJz6UeB7yyMG+cMZhL4flwUuOFfKXK8bxKTDA14n2xmfTWXmfPjgcj53
VihJ4H5VuJzinz/jA9b549k/sf7NCioPHwGLGd7+XRbPI/DnmqaylNSWwOl4
SxN18wgXriSNlCJFHVupAbBuP4rXt32VIwpGH549/K8rMgM3cHpT9+LJwUPP
ODKy+/Ts8ivRpWqG4X+L9dfzzFFtOzAibqhSFQk0PLnwcwC4p0l4UazHILo0
EJm1q2JwY3VADFDmpbO/3rydDCzjvuzfH8gTi8E86D7kmGJHKC1FjOwokFQK
nsfDarJSerDZko2WZLHAkDt9+tHanNRrVrvR6F6d/yEVWiEjV7zVT4C7JJ2s
GBWceErnC/k9e4q8CbOiLbYs5LG/2zp+JqX1P9G6i0CsaU78jEK+is/PjH8f
68vNiSgV+FFOYm2tUG8wYUGwXi1dsrE2urotyhUgX3Vl6kSp0wM+gcVvFhyh
BVKWcl+BCj2vnhJUR8jfw1r3KFARdxoCO/jF1cCsKuhvWYZQpLvwQXWDQ5iq
N+QtAtXlSb85C+CaTd9V2TBfQKNHxcvw8WQ1rDhNM7wKgn4mtPV5yYeizXNE
QeKFLcg5JaS4VwPObfxogacz0PLkNIX9pzYD58b8TtVBsFDq9Mk5csyim0Vh
MUwACtxcHzgmgZu4VvKkssWdoib6aL7HKULOTZpkurMP6NZDW0xXn0O1beSc
dkK3HSYVpaADxhHUXQCm7kytfAa3pbMGbr2H18QrZAcCylXQV3tmqTlw+VSx
g99APekxvSFVqzflQsMpyL+5LkGKPWJ5efgbA/N6pfFqDdCsEZU+kYoB+LcV
3+8QCevi7fMjd648/UdkB1scjNff/r+yObuWfUaQPypqJn29nX11hrOrYipc
CBPS6PkP9OTv1jnZ3nzvBcD6N5YgkO8EqkddOtAm01W1tUKMxilwJldlBiin
fdhE8SmAoUl5BvMQtjHBo40AkJzt3OwuKTp/SfLp797rBVNcI3VQLyTUMRal
vnqSR3riEwJqgdo0Gjobm9AIqsCHyVhbyucA0P5RhrCf1lzgqEGf2mXDzQAb
mSG2Bw0qdJwodc9qpow2dKl7dyWPMcUcRUZao7B2eTPYqVpj5fW3n5PXTaAb
A2WVwnMk9HwWaujqnb3E/iPLLZtsg7FwO0yjuOR/EnymHmkcBJzNYbRADeiq
AXYsHW7sYfoQvB/mtlvI4e1gDKv9Oclx4O3Baq1QkDc97wEN3W53xSKYHicY
qFc5DGjSdMelClUsCx0Zvu7nIDFKwz0xRQFlofW29EzdTvRajS3eWcxB9VDA
Wtjv47rr3hFNjqvbI2s9WXopPkzquTeNQqXDW5Y+vbjUUSlBMM4VsytXDFPV
hQLqiUUC3N6yvutUmiDPutdR9LM5p3bui+V1SrWcLhYiZWweTEDCHxzJ87kt
hBWh9oP9tfXvgxfQLKSzEHqH1lcJUPGy4O0eO25yKyiSTeeR3WqOCjbGrm9v
hG3RVUNO4iSw/kfik7OCY4KiMvynQijS63dUDoD06QsjlZHWz66gtOUcl+CO
gaKVQk7/xHxUWUstRDeT2oi6t/PEU+dlP38KIp8Z0cCvUqQMv9TmmbeHkZiT
HNrXXkz90I0hhxW1BW/G0WKgO+cF9jj2n/5uy+TS1UkFVBP+7J20ORjOe44b
WEjWghtcIL8fu/qlFrc1CWPbQRfFvb27cnlNnqwNZLD8fSaFA4+HkxKPxN6y
2u2UkYGEn9jCkXqarAd+pIxCQ9xpWv1FaX/uIcSeh0GvffDncTJ5cQsC2JPQ
ucU6JHJRWoTpdrIuE4o0XpT9ThKz7Og48gGTjlzIzHZJjC+LX1czCDV3ptHx
gF2yQ7jsM4gqteu6YNC6NEYyA5A7FNeuOztPSGQQjOGJ7uHg85SfWAGjpzvk
IyR1J/8o8j0kFjBjUEmjXR+Gxab4Q5j9EDaWzCnqeiRUpvsiUS662pDa4fOc
PtHtvX0rhGt8AmRFtBeV1XuQZE//Qswlqzl4pJ/C2Ef0WEgD8J9j9YqvS8s6
nhEKXQUYp8lO5ljEDf0PbU41NTjgMI5jCe6RiS6tU9Yv480w+4RtQovmOhyt
eEKLXh1fADGCTeD6103pOZxH2DsjGurosyFRTunVoybty1eHZIlHIE3SU8Dh
S7kMApNPfHorU9+Sw7LBpAgzJA57m2tMH410zkVYpReH3HrRIIDPGJAzc/cg
kbJ70D0nRCme5ZRFGNq6HZfYoLUEyU9Ph8UnE+5+Rvb6DLbAnYYU7tOkoPkU
XbTajK2ks6IUQax23zroToTgYR0wYwhXRJuRz+I1fwuZxCeOYRZfZRAu5MTH
e6C5srkXAaO/kPJLrNtGpxXWGJLTi9LLrAS8zhElO/MfVzK8XuSdQSFCpFfo
UuSZK9I7t3KSU8pGDT8ytjLgPZRkpsnZsJQKk3/5tUMqvbTYGOW4cSLKpbu+
KaDx/nirSeoBwkDlyilulZwcSIro5Nr3zkaBmvrH9RVB6qj2RIbXaln2Ucrc
DH4SAtIiYU8uoHFhKa/loRkQsqrNGvcbGiwKruCWsbCDK8prnTiXbVNzWnjO
O1qAxmEtDSVm7wEZYcb6r/1+uZFy4P6nQHY6GMApYjW9geYwgq37rgMcWA0F
L2+4JvPOcf+Z8hl2iuJFO1oDOvGjJoR3tRxrO/LtJcPMEeGmuEzzqT1rmBt1
jqeN4PJ1EvLlyG4ydFjs8Jxs+JuJbkbVAqJqfx2nPMHwl0NMG4rnchD45d27
1E5NvFqqojr24Uyfnnj7Pt8e1orz9TsaOwiIWeQ0mCsD66RcMBnei/+bfEsX
tUguO+goDvMss4kqAjEZcA9vk83GJi4DhBpyA4RFhOoIfHdYKTnVziyeayIo
Kc+TmHzkdlvf8SryTLelPfpbuq96DID+5e9PIW+DB7L9LcFLC5W8sl7yq52A
iDRzyQMt7oYK2ib9fhArOiamYi/3RrzYwmn1t8m9E7YYQCry4pIMLrK8Z+P/
6sN7jlTy9v8OHbFr70FAqWDeiB0Wob48yPjywnU80rdKhB9a9Q2pdQhNAseC
l0NeO+y3Y9QJSZcs1RaQrhOROnO3/xTTKb2ytdMVJnLWwCHwFyTD2TMmpUYX
L4KqlEcW2bKH928jinSLshachZlLNdaiA0VoHII8SutvXOs5JHtV54CqbgIr
gBbtI9e0rwmSgQNXytntyPQabyJUi24DdjATUStho6w18r3mFNQnyT1s+sHv
vxZ2m8hzmDi+XJNpUXrcwSzH9cWPFOWX9vxhthceswtHPZ+yAQkRWBinL60Y
TNW28KZtDsDmUqV59qOh2UTPzqftnWadSXOCSXTjB+ROmtBWOjIZrRMuS3nZ
qJhEy27Dfko0e8fQa3vP40Ajzmg1CRJXLUkS8cs6EcuJ4iMgfup3LlNUAybQ
lNpsYoqw2cYdhe+xhct4jhcdhQnPdyZPfAF2B7ohkgILf8+qmtF546nqpJfG
oUBgB0KTsEUOhuGJ8zSaAqq/u6nev26JtKY0qyucBmFmhDxMERTt50gx/vyq
NCIyoPXVPDLBZYDvdmlLJcDIVekoHv5+RiKtsaXuvFPkEO+Q+P5ZmWMvuuuD
LJ3zs5mtKVxLN/ZlLGBL0mIXZCw3L/pUf1ku7rXYYVLtHIRY9zHv2JVeHjQP
7DrOJR4SGjtzHBZJvrEwMKfYywFkFJc+dIUtGENkmyUz3ZSuQlQH/jJIetCu
6wg+hSFivbZHSQUxsOCLmdQ9PiomdknxAT6G28m/WCCnn59JnU4tBxes5IrD
YJec9KRkxNt6wBB6DNK07m9uM6a87/za8WuMLo6sf8h36VjqpEw9JvfE/gjl
JjR/zlMiBYJ9QTuFXg26GPWynwOtdEDmkg9F1vJSJlKhKEssbOxIaaPon56/
/m4wgYmuajjvEwzjJ8KmoBe1yKaeoSqJDpkvXZeq0aGT9AaLs3TEN0/0/h0X
YuvgEIK0zDHrvWs2NQUIJXlgIe03TfVQ1YRAu4bJ5ILCGNoyqJSdgYHQ436F
S8L/LdiRQhQqUZXtKe3qQMfnuGaBW6Arg4YAyXVTLHOrEpc/LX5EXLHuzha9
DlzlYcOsxJd9v3im7UPf4vCrMBT/LRTw+U3zToNjdY+TXr1YFmvwqSIWO+S4
FY66V1RZmuAfOsq4IbhZWCaKqm7G15nfmhrKx2hqs7Mx7+TTjITd+7B4M+Fd
KjXCuoD/bBVsWz1AO96TZW4CGx6VfRR89dQXYViGUH3rG4erYw0dX08zRYLe
xnqrrZQkVPXTNnhw5TFzz8pExw4R3eSY94HMYseh5yh31PQoaWG0z2w+wqAE
PVZNpxZAH08lyPi0BAqO6womlJHeU/STsHqX83G5qdlyxkORhA8w3vz2Phpm
a0R2Oh21092M6uS6tWTCiI9+hKXA0ALrKl+QMa5uPZs5+nnx+vtPAOhLQWB8
PYaz2w6iRPH4D5PH8EpsXROFhOn6C+JDqmmSSlXdJhjGtB1ZuS+qhb06RM/1
xbB5EkW8ZX2t7kpUzB7sFCFwVWeRB2PMSLc6qOY0D4+k5XSECB8bm7f1FI23
JqGq7tl66DZzofbPaygh9c7m/DJZeo+k2sZ0ZXEfTDVXUkcjE37V/zm5fed9
nDVN6bEO+5h9AGkoo0ImwfwS4HBeFRamlrJ9gX1vuPQz8IibxFMY6o0bphJP
5guh7p4XfRL5h3rTEvOW6W6wtQUEluX0RZvlTQbCYA6cPxplCgcB7Vx8zfXp
rqHN21rB1SyaTh7FrfnSSmYg6g2krGUU/ViWTSbzNNFIY618RQfSmFw5V+b/
QU7H96cAznZgAW5V9/xrU9MB5rvukchL690SlrwQl1bb1J9cq3uOMt4GZkMK
idcl1LIR42bdT3pmjqH0YByCECf8KhWMZr2A5l4n0o7M4iMp9pFWXL9pH4YV
BaCqLZHr9TNOKWXBznHLxJo/eQMKu2qIdvs44TIjj6d9B1bHAf2WHWwxWkEN
LIHlLznZe8sjwQ42c5vsGc+Ygo/fwsyS2yVIvNRwk90/42VHfQi4NxfE1gDn
HKgjLzzZpYPi0AMrzTklqXHq6KZPdNxpRyweDvWfZk40EngrJtBfH2kWvIyG
BSpwjhA3PRlJd0nqmrelXcM2dwJ856HIKCToXUUicgIj6pjVifeCDNir/1If
m1obsIZ9tWozwPrvUmpJosXV+ubaDKybZiUMiqJcmZYvgxqqMcK4E02mZ/jd
uIbu+GM82GGhpL1uuY2F1+zkAvzNJcB1sXF512C2cvrkmJ4u3VCx2oJILdY2
oPD2nGVpl40IiPVa6eMfoh++XUhCHq1nIPigcJpQsTjxH98IGhyhisiexY2c
Aa44J92YEwHTdo6nznueytfquV0CEWhIJRWZ3xN46MVHOBAMVz2D4XII/+zu
Wy/SKxQ8wjEIzfAOwT4b66Meh4UE8S/lsrpqSVtFoR5yIrwYMNqFi0XITtoA
Q+kUaWoi0arUhdVl1RTYpWH3GZ6e39J7ZH+P9ccyKVWJxPWFm3s3Ob3l8OMx
bTrZs+Pb26LaliuBIzVbuu6BSMzbFlHDtcpm4zS2nFlfB0BUI+a3eH6bmqjJ
Bb5qPqTZfd4H5NcNbQiDLvoBV+a+VZG7cFA0j77QWdHB0LciPupDIbUeXMWo
lyXEzPQuTp35pbvuxm1pmY8tnwmHnrUfIG4fcgsoZYMwv+0//DPGL7P8R8Ry
rjKS63oYTgJXTueBV6nWJZ+7I+MnLZ9jESk2ZwcwrUePlJy13mrIlnSga6SW
VvGZ6+eSjiLgzlV4lcxcwmFZJZwD/psGJ8C+YP3alzSIDJvqNhPzS4IOlZkX
ys0q7epA9J0iESunPpej2wGnwVGgmxpx66USbmUzHER9XpW6L5YrH+e+w4ha
7N8BoeKc57fy9pTub08EgGpgtwcB9hGpBFUWMaAjERN4x38tpwH/gUm7F7Ch
ulgG3+l+KxRCFWfvE+mgIQhgnCgUR1Y9Mw1ApS7zT9+JAey2ABCWeMsIzBYS
bX5LE9+9leLNjemy8M9m8i9q59bW5v8btj4qIZQNClBgopf2OuFHTy9vAO5Y
5bQlnI8zAIjEyu1kATLLzwHaLufYhKqM9C98htq/bZXeW4K0KR1AOiEM6flP
KoNsvGWUkmhcpeVpa4POTYI9zfvafwwk5pEASfrAmHA+Y6lIRfvYTErIcsgV
zhafIJLsNEkicneqPmGVhsmFUaHOa7YnD8xXxFj4qpHWtCcquiULtOQRqGmB
jGgnsWcuHOEY5IWg47uGewluKOjH1d//rvtbgwsX9FJswakQmx+7ugaW92ZL
CR/SKSnFTCUXWLc4RVvHJyhmsE8weQ6QLhM9MyTfHT5ivmcvlYTxkl9uqzHH
9zUdpghK/00NU4voFnyCG3nc4WoJjVVvjQ1kGIZmv1Gkc2B0uX0Q6E/gVQk8
2smtGn+By+9ZR/fPuGpvBVxet0wHwk5xuMpY6vta1Awfq3ErHO00752cL/zb
qo5OTXlW9VWRuukxAzvYcQr7Pl7KACXwIcENyUTptmwMVWwVSxe3dVVesXkZ
kn4qjllj4RRhpExd9vtHfFQNXdtGHfEQtPHdqMtUhbLfKQ3V0pt7I6IqIRui
2u/ZOv8Bya5oJNanbE/O3ZlLZTUj4rHMoYQ6lt5GIpipUDBSipmT2Be4TBAE
5Ng7hk0JBM9uH7UJ1OL40PIIJasEtBCmUBZpDIR8NN4MAuY3a+F44de1GLzR
LuCpckEeYu3wTcR70zzfAU9ohosYO40c+oLnWThKnGU6nHgnkaBumNi+iHXM
SSJ77pY4Zkhh4tIiAj+Et+LDPGoVFmruPt97PG99Ko6sYkDYSNgcx81IrVWB
nFnoCJUNcczRWnT+9cASLIIBAMW7Xd7Qqt6C45v/72n2rPUkGmQ563QEXF2j
iGu2T74hAlU4nyWsVd8Tx+nmIfVv9t4kquyRHgx69/Q+I+dOqzl/nZv1Y8G6
sTsV5zIrcz7C1slO+WqwGzxYTH1j5nxOlNWcZNUBTWqGFpS2MSxHRMSjQxGQ
7eQmT7sqfQ8m1o3pJEYyfvUsFCdxC/g5MJgwotpA6X2SfxBNZWxalLzv/r5z
9Np/0koASQl/udeA9H77Lb8g4TkWm6SjZtFxkS9XcHiXPxCw4EVFkz4eMvQ8
4vjs3i2MBMm89jCTigqaRwzd7YW5wf9uxssfN+joOjBPXQxvleQ3X8ZJMu7t
D1uISaFl7fNDSYeQmhnGKRx66he6cIrrOrVCSqd0x/kBAUHCJ88ghpdP1eqo
kbFsIK277/uSVzHpQdLS7Em+n7bQHb5ctZ3hmPBvEa30quREh3x0i7gul4R2
I9/8iUsa5+G027ZrqMQ/TY9VWrC23ggFySpzRBoLmTg6d2o/zqzRq6q61rrJ
ggbx5XcjLax+OnulhSosKO+UhwuafLirUmL1TRx6DiUPyXnY/lMYBqGQnDi1
8/XhVbSF4tbyFtC2NXXPT+bDSuu7mWtKJqmUKuPhS/Y4b2hh6WnAnZHGV50J
uqUbs2VZlovRj0xdXquCh9TgtpO0uLVzs/sj9lB+NfopM5hucVYMrASZVDTq
tspzXhSjpmoa31ZA9RIf5hsJSgHrSLw7KLb38lektov5E9l65mC7LD7CgB1+
li8QAe7G/j92JbQxN+/njMW7h/x/QKkuKNeb6i/cQP0lq9Ct+EAd4nAyDFvp
BDatoe9AVA2Xh0T5mwuDvDGlxGWWiZmXhd71sSh8NnAZWLKgqG+LeNhKiKj0
C10Ej7KKcopQkU3mOVuMC8kt1qGymlOijlRqLL5IFH9oiX5G0RUg117CoTgr
ixaAWY4HQZSIid97vpUI2lPVLpcFD5NBURIT7ST7rf0oXQGWD/epzUEUZ58m
tsqbZyqbCFk5tROYdZfbRmn0W1PhemcXtmwyk2jK+oYYX5F+hdxix+49D8ca
GH+j54bLcS+TBdN4pdsert6wQ8285PYTr2HKApGHr+3XTRBVqRi8cHjuM06S
lA4zLlHUMVv4mbzfM30K8ROdtdi6r76VFJyRDNxLgM7XR2fXKbd4LbOpj9Ow
t+ZsbHRh2viN55xJYbsMe1PwwWikWRlj1hHTQ4Rthij/SPodUuZFH6qXn2NQ
sVCfz1u5fEzlEjuzKSJq0k1aDQ7mkyEdV19TRWNlHFH82NgCWJtCo/HzUkA4
fDUvjDhPA1wfRtqlAi0rxvoosxtupuSUxg79SL2v1xikdzl1VI62mcCOETpd
WUBQ9MeKd4j+j+Ju3IvRPlCg+aXPelAcA31ZCNI5XRkvGibkxq2l0HTI/Rf0
RnVkU42+swdXTFjeRCE3bMc7BjPVPWPTKWIERJsQX9BwxOkx6W38Wi4gqhUM
PPDGeRtVhNIwJTn1leVkmEVT1I+LLRMQEUrNCLb3kPNjpFkvhjG4iGj1R1i8
MMJxDHUkWjjw5fW2L2vEMt6zySEIxo7aORBfWjd3ZF/NLv2PyfhTKCNWvjI3
IzMUH5EfrnSm/3hpsLlJOnW+uK/+OBtZhEMXBPvpFrApswEwIv0OiVK4m5ET
bGa+Jr44TeBy9ZLr3Xi1fgDDki5kapKbrfs5H/z+9TeqSyR6I2qGyMpwnm7u
VdnjlFO8N31zOzc9gi/7pdmJgjp1z6FL6PvSWO69PJYYKuYlcZoEOZ4q/M1k
DuS7pGxTCqVWc/2sq5xrcQB7ig4/nOc5njSkUl87P5QVIG2kzkuWZXKr/QB0
PhVxEMN6rAbIJQ85Pu4UymK6rK0ro5NiUJrlVgdN99dGuywvn2f1KPeSToeP
Sv8r78K/xGaZH4STSS8ZjtcdywtlFX1DZdK+7muB+tnAudnC9GKxxFqdKd1Z
DeIjwJQyODVMKpabSkgh8HIvoHc2v+1U2+BwHcD4O1uOMQ+E1UzMYx3P4WFG
kOBqfhqsbLC3urxU3ljkQuTFDKMrB8wtp/jqT1IBCUMMyxluL/Ma+1EQbxsn
Z3qMon3H8C698pXeLT1V/CcTmQhGVvSkt/2+MmeN4kmVP74TMjowbhe4zNsj
Ttj4FxDrmGyxm67tpclfez/JMxZFPNhMRtmLduGrnLQa5P+nDAP9abfaKb52
hH2tv1Py/Jf482PmPKi11NwXOHU4DfrlZxemK/z0yQvSQtqdB3lqM7KDTeGY
Y2hs3njc8/FoqvqvpymlkZv6mJKNqwCaqZW8tedFedJibKrTC6OuTg/3q5Hn
H8217xl5C3RAb2zV6WW3XJg9BRCDy3R0GtPzBzWXusIHhXwFEj34ENHEJNAf
RUIk4bnThCZTgZuA1bjhn5G3zfXBzIDZwkN0t8+LdBA5XuuA/KCOOdctY/um
BkwFqPIR2LoLyR2JclOSOp0grJX1tXe1N5iCMZG5Tl2o1VkwQEFr27EsTztE
uSZVs+W/08FALEN2EHWoBOwoaZZfg2M8k+1j5sV2W1+k5fFKorLiaOSbZAOF
9QpU7NTSKiA3RPzEBQaZlbGxZLv3piKUtR0maOOBcDoScxVQlrPHQ+/c2NiV
AsrUlLp6ZNODZpEjvLjzEUkrVXFz7Oa6VYj2wxnCp6atgZWZc6dyUTOHfWkD
c1TZ+SOvow8tJ11ppuzWItjrMnw7TVk2BejZjQMgLg6ugW7XjRgUXwlKiTEb
NBrRf+M7RcLYhciIrMtUCMa2hx3x/hgtV89TYchZ6GjH8BdbVuTikdbdTSjP
3YvI1C22Vxj4zeFmS0SuKRWu1SKI0DtEghTudPnDR9xSAKzF2wcNfXZ+Hwbi
kvEt4HFFyXuz2HDFvHeWe2noMFQFLHpKKBN5z598/dzPLNgE2hM1JetEbkZ4
b7gaKRDAwzfH1stGRZDNHj8PK7s+SAsulzdiyvjf46+UIAKMBTnIgAxl6E+p
sydZGhARqkyXlTAHCRS/0jUjPdF9J9Y4ppvZu6P0Ajwb6Lql2Rjpz4lD48BE
lQSW0LvJBp9nhB10ST30i+wlW32LPfxyoeQ73pIYPagdaQGxzULMUJ2NGFCe
LlG3x9hSxuz0/3tVXa3wIAptvFegNNC8qHEroTpeslXZ5Kq7j7hYVIz3eS8Q
RpbbjVKLdMGWUgQ1bCj/GWqN0PzFLd9UjXWmi9zYs/81r3OUeeVhSTuiui3R
g89znO8fJBAFYQNWUaoEWcNX9mr/MViEEponxR4HwJ+eiYgkGz+WAXEpSgX3
jrnNdrbL8RQtXULN7bP+Dr3AwjkBeYUFOmH7ggr7LFSqQGqsY/ZzAcfXwWZh
ejLP/q3q5gKtc996CNWHfPGoUIAulZcqZJ7EGBNpse5zPDI2+dtPqtBYiPUR
RbFqI+ZUrOPLeJe6IlkWGb1XPMPwZP9KxiA181RFAq0oQ6Zuc+T58s3/z8m2
CmRiFRMOlWvlXx1OAgtAR0yoR+/xEPhPRgjBs7tlm/cLmwHIgunHUGGuhhf4
viWFTSm577Llv/UpNQfwshyrY4abRCd0cguhiVulVkaWy27KTssjZeayj+FQ
Ap2MoDPIf75jcNOSpICIusUbFtWpJ1Cyf/BEBnt/YDdxa7p2LmuyBEp/Q9dU
gB4jGR+bf2G6uC2nGL1avJ6p3kKDc/erVrsd+yxiGHf9Ebt4mGqIuI5aAF6S
f5floSCqRzKQR3dnuGCMGkhSYRql+JfZFHgi9iJf6fbNFyKn5/C6ifL1aXY7
casFF14aTJh+DwGLmzlU2JK33BjbT6KqMka9k+fNFYpkRWxW5o4R6MeXcKb8
AaPsZnRrBztNJ+RX66sn0ydIAij1nNcv9ZlagBbLVx/nhuLENFMqE1ZeVdem
zGs79c8BO0E3zqxb06TCK/DYaUkrfe5eJlggGnV+hYyAsxX0Epu88itQJIr0
iaywn5rCTH/t3ghQV/J8l8pO9VMNPYBMIEQULvGZbYLtUCqYlwcEKFl3YJcy
bsZtJHur3IeRxoEhUpQAThypglbsp0IdfaGEeyOKiFDHBu+cQeB149jZCRct
5MNmGEX2aPKLy58pjvvZ1GzJRh9Ej60tsgftuyQUIys8lWuKrOYTUISJ9mwl
LvrmzcxjZ9zwlmqFoYNpwNLrC5ABkG6srq4tK4DM6WCEq3I8JrL3KJxbo77w
CgWodSFLL2gZc/uUto50KcGE3cLGjKqJHDtdE8EeIshIdGOHPqP+S98o3OMz
BwF5qZ6AE6XRmpNTeCNZbrs/yQbZwPIi5aiHYhasvNt2sqZ4Dtw8ksDp5ibL
htNrr5nfH+VRuEuxuVUOPhUkkMnUxSx6a+yjbTsYf+hidY0fWikWCZVWHzWw
e0PSpKf1mScUFmiFQzablncLQFoJm9I9psZNCdfBcdWrwT+u2bVEKiOdyFdA
4uOIP2iwUUJUD8cxvizPa10uNbDk/BDEwwcoGiaQRbVj+oBuOv1fNrlXzYZY
yHbiHWyQ9pyr68sTXctYVZHU4xgLP1CfoqPyvmaQvbdxdG9PoNPljbJALZR9
ifY5cc4RaTXbiYQWvEJuEUYQoxbzUODU9rH7ufhoG2wC4gvABN33WZK7pC2B
ghyFN1azOi2ehdeXxX1thM7vpVjBCX4Fd8uAsxv900B5Q1AQz+pDpkQDbdon
PAU2/i9BUXeK3aHIGnHJBsuoQh98sfWdnXnxdDsSSXy2sIhXZDoGzwnUgPr/
C2iksMDaD3FEXEhAe1YdCMh6I081I8Uu787r82Bb7RP9PPI71hMQSRChpqR7
V9/WBnsTL9JLdK5uJWdVASOv2dweVGLbF3cbfgowB3q+0awFJQ6NRtgXeXol
nhZ/yvuWeO+o+pDDgt1FOokJKRjd8nIfzjsEdF6lwnaMMWIf6sCexmVR5iKl
2efXo27fbMH4PA5MOXmVDOJjUrNqPQEPcMSU2s2JhG2VX13xuG3uiKWPVI49
0p5AYqtGaF0FiLrgs9M2wvoKIAu6WLZ6P4qCBUIwqARhEUpWMHdPhnaFHXEh
d9VolgnZuS7i1yqf/rh5C4vqyx+Z0PTwu30i/efU7CIPHoKpV0ydxc0iDNgc
RfMEHaAMbWuCq3pywV26znwDaihRRrbpO/Jmvexo63DoK6FnqR22cVYA48U/
tyOb2uPyKLaxKLwDxugu9X5DDobECyKAEjo7vgny28WCPJplUgnm4iiZco8z
PwPJy8wZy/92JyX/o8FqCm/sbrBAv3p0RT/Ebwh5ZV91pTcOeZd5KybfLIDe
+SoZTdvionD02fso6wmaAHt+/jITS5SYFgnnlAJn/2tEq4gO2IVYKf2O6Qgj
zs+DqBS2nG0RvFsthU4iEcIuwf2ylKf3iXxHLV/PKtMjfkcx7agD1GJNGPRj
HWYFG/xF/6++GcJoPmHm1dW5KO2hf3GNOVyrGDqPwrqf9TWiMYspRLNBQAnl
iyyKuCYN289RCVqMOZJNBL9GREtyGmBLm8oSNWyioPd7Mrng0+Yc09FVrkWc
kotsOR5mi7PA7ONIMGQsEIF0yhLCLa2+tZd0CF3DF3R63LQnAlaF7uV3ttBR
/lJqQtBR8fuj5suUC16yHfi3KrbO0BfrYxNhIikAg/mHEJjN5QhaLg7C5+Do
C1Uc0YlhDtHdAXAVgEu1PujO8urg+iA2OLWV/a5pPXpo3nIgxRAdKtaoNl2u
UgXVxaF8bpAywxmGnQqlWGtSAvellyWK3JYOFXB83ZKsaQJP06XFYkg1/8FT
DiourhuxN045K1ItiA9quTuHQHClyt9Eoou8Yiuqd6ATlcFaxUaQdETnOJZe
bS/0/ROsumq8DraLaoZPeJmrfWcVG+AC658Kl9SiqaBpUDE4voZc+ZkayMY/
sv+ylrXiG5TE7mBXPlbKB1SQvbnzaphEsLFiqf6w5ZKt9SSHeAXIU0RyQwYt
oUWkPiZLjTqkr9VlA1ZF2avvTwcFGaA7/sZP/wHQIuRdsl2jj97gHipLQHIG
bkGE4iINPF6WYMHdMPOGZDIybwmnfMc8O0AFuMYEY/OICJZo+iSREnjRA5Wd
NHj2uYyN3PDz17YOG12H7bRZHRLD7c+3YXP67md9zEPVX3BybqmodbNyQAjo
T+cIYoPhVB48ilI/zLsZYEuJEEKW57YijWdiHR+2a49XVAmVywBu2gm28wVn
EOISLpKMYMGc3vIxhdLnJcO2Bvh+wAmXdTdDHahF/pQCeJv1fb810Y3h0MzS
y7zHTlIaisu4ldIklGfqmdALk8ildAWjXaKbwuEnajaz4D/LxCwPG398WiEA
EddFWj/6DVhDH9z/zFivyPDaiO5cF76pSEQ7Oq+beGI4H3S4Zh75KItPzW9f
q/8Ns8qkXS1tI6JOEIWUedbnkQeBzLosQFAJf/k8VdrqPLbb4vw27gcvSOqX
0F/sj8EPlXOk6kGbIBwKMdnLQyezzVSJOA4LrptBG1jtWwJhq60QQwKIK0vW
BuPbL/jioINulBplIsWjJixchQi3DLfyz9pmec9ucNl8NamFzINtZWIsEvbw
6auM6rvfZph6Uoz1HOkQkii8nljUNqGtZax2bXIZGeJydUH4u6a/Qeu8eEXL
nYxUlThv9JZ7bCc9mz+6oyqE4fuk1bZ/gQyF2QHIdvQPRMJXULeRwfHJM17F
I7TpIERTAIcrmYgGeTwQkI85/CvSdQMwmOIFYhaK6La4UA/N7Q4e2auirAcE
FpnY9rB3VgTWO0eaT5OgSaffk2RjEEWZ01ZWMC1q+C3j2qayUS1+ubRXOF68
BP2Rmqdb57tGu7+u+Ts6JqX836SUdeiwVVDfPr/Fx4I/UkjpbvY0z+hSYPKL
Z7hjmm+qOhG9cIuuEMFnLDsn87sXS/SOrjAuN4MnTLW+C5GAAVSgIQsy3e41
KODaTaSNZTHvipccaXTE0+HIe9rjMbGRsIPiNPEpYfO9hPfgH+Yg2t9tedYO
Ld8+P6CXdNRfIH0nKSWaG8WfVuIwXUTsJCa1cpiePmaafWtreM8npi9Uc6QT
s3crmghRz0rKJwt5LjroqocHbl7UgylxBQGOtXGwTphZoyCJkSpEl92ocDAH
KswHj62b9Dwf3EQbARaXnvIjWz+HsarnT4fcxS+XYUAz+H+MhPWuAKx4ZlSd
1/XXW/bF7snJYTe78a6qc5mEdPyBNevAPoBKIm1O9ckKmpVzIeXnxYkr2IS8
7e7bWAGygWrob/N4cD/i6ZwVCo+5r/hvyOPfgVIDpBBTuWzMxiAWAZaKKQMU
Nku+ztDkWEOT3PbksVFWEk8YD26aSDFWqJeENLHaDqUvCJ9/iEQO1/Oi0rT5
qIIGMFQs8rNgp1E+edutv8IJ9CyyGvf+RN/+JgYbSI0yeUEuelMaSaP3XdiD
DP1iuD/KmrKY9Iz3wKBQRhJEAheJ+mhxkS+5O0reV3AfWHK/o2zz8ctMLGGo
4VQgcDFChVdVA7gSvXnvBZrFb+wF6VFzZWInfg3c1zayqTGAvqBFFLC6RWCS
dya4mAwwrhFzGBeL4/jV0tJktVrV/PddLjfQpeLc8/7+iAxgFjZ5XgtKfQbm
38K2TK+r/+8AipDIBVTaPYqnQ3Fxl4gvUIZ0oqEY/fvHUhjphNoyk0Z6dJL6
hL5kAIWp7r2e15ym97tChUXsMvcBY+GUDnqVzImoXMYPChjDfTbtFbrxa7Eg
CFC9VmzfXcVGaw59bblO/ZAJMiBSAgwAR/ViRDAeKFu83/+5qQPhkOhukkVB
qMW80WkaMDzxXOAOy4WCU80s3XKeIWt+hABw3j+lshL3CBVIQNyvuYer9PKE
AbpOXqqRNbq+SOfA9lZTIHVsNGBZvJOo1JTBT4jdpWjZ9ERUUaZVoxufn49k
e2P92c1Kz/OHS9wtNYIk9o6G73k/BMZBjFlh446wwx4IZq0jZDlWqySwyVz1
wwSioGziI0UwkkTXlcqe+ceZU3NPZhOJoJQ09d2nM/aQ0mu+N8EwzjufErtG
l3FqBhGYJ/KmWjr28p/r1qdWq3IOpUll/PyGwM6iwtkUlVrYCXlfOScv7Bcc
8XLASi/rns+bzlXmuFdlqNncwUkd9Tz1Ss5E85llK3mf1cVk07FrCwdJ8DdO
8pERUo2o1UfAReXrSjvt09Jr4/x00P/RSjnXabJbvMGprKKYveP5ym4TUwoW
e83GvS197f6zrZr8vw5BKXyxdXD3PIG4sNOV0FyZciQEEHHo3hEGKVO7LNMD
fbmP25QvKYagC/r3PmeJSDhRqcsQsi+/LuO8nIC377cid7nTzUJ86UGqq1mH
fRP131htW+WC6+npqOggxiUkVD2+kjyP0h2Fz95YbaG0HsrozRma5ZDhXqQI
vpvOHYgBRGDvpHZ8cGLqBQ6VqrashSeu0kNAOp8V0fWfxErpgKJsQx++c1CH
UALSWY6rQzdQgHMWCtRKuQm6dD2FwlsS+x+KXwyisf9hg/l/kOQkGJYTt7Nl
lhqGbDDgrlYQaNh3dKojgyECXuIPtmTX7ZmVkr74NlKghwPq7p1KVwbRrU/+
xNlZx9lLcggS4boNgWNWI36zVHfKmPk8V5co0AbhMqmiOwoaNZmI/WQ0CiXq
PmFhSWGVOXnDVR+r3vMHwC1Q/m7XWZDK9IZP6mdNcW92yVlMcu//ubUW4yEG
I989mU81xhFHMG774+GvXNZs1hq1CGcN5eTPhF7hROn7RSy29WLvWlRbZXvU
GDa/k/7KmWKtAd9zQZSgXFCtcQ6x1LhDun8jlizQDAx6cHUmelfj3Yi6QDkO
QHB4GDoEcqVX7pcOkGTjM/OZAlhkodiFAcVnWumCvL9Zmjb+CRoyBPqbMzDR
Tn2p1qG8R6jCAzwi5wjzbfShlcmfDZqxbE964XeuGSUY2LO4jDpjUd26AFtQ
o4EaMgjuk0NHaYFHkwlRe/ti0A1yMquw2BLEeRVUnsFY9G3CfNWLnuYxv/H1
hvqXtn5UtwPb3nz7ZtDZygpU0xUlN5RJsStuPEQ09qWRzFOH5Px8ykDB56to
52a0Cns1sbXuQdRj+j+y+Z+UVeFdyQNfCnluXbDNlIbsngakPrXeNlxrnLNS
JShX/BJjLPkmTQbZ8ym6UHoDxFcHTRdT2dvXUpy80SQrjGnYsJDZqbF4e0/D
0K32Eq4gtD+uQss/kZZGhV6521k8wuHWfEC1Mwi7CScOqaQUoNhNsAxSiYhC
IQDiTqaE7WZUR9Jxbf+BcaHJZ+99bOATuCgS3l06b1mt3npWCaDZ6Exog1MO
bOjkBCyoZrvRaQPu0z0C4YHTKcTRvl+yRocH1ro510S233yDzWSSXRILCMa7
uvO6BzIpkXWiP4wa16Mhgwt4jfGE8Nz+JK8A3fAuA71LcGF0XsUcb3+LqaA2
b4OhsihUmn1gWEtkk2i9jVQ2/QB/Ru7lBZTii9KZwcbupe7Cqu/XmfC3A2bI
3PRMYuapKayOWc6iY8fWIcACeWc4zG0KBVBLVyXNqni24mkgCjSoHpcbU5qK
5X4C22b2cJU1EGDTPcY6lQ8HVBqailu3sinRa/37o6XOGfpJQK1lIG5e0VUj
hrk7ja/Xp7aws77O5ozvmc+sbKNFIyug0bso/pznRnTF90UVlmj6Q/AQ2Agf
Q31FrS9Wzg1rYeGB15vcP3haR5NjhDYgAeIpPef64umczdglS8ctMZwiGH3+
UXl903bFtx14OLhrg3aCtr3Bl94aX0WvPffhl2y50Rr5g1yizjy57A8l+gpk
KNGPVTvd3P9JRQpcRktNkCnP2+mndEpTOH9hJ2JXd7GYpwfZBTYLB/bYMUF7
mY3ajZbX69Vcvf4NZ2YauiSwmWk+GRzZR+b2UrlwBN4YtpQSEZByIQ7sW5/b
vdmrbMJwEwE5VC9AMn3LqpDQIOaj4vAJ9w8j7I3T0/g+5iOnS8dzwY0cb2jg
f5GgAwhVigVZ0VKmhAAsptHA1AyHCV6Mjm9DltRKoQexYQyDMRgzHBkl+b+S
qtLEULvtNuALQyWyLQog8IYsKUJDqFM9Vk999KX8uo8Wufxe+cldDNm7d3zV
DyYsiXuaXT/eNoj3SFudJBfMpJPC6HrRVJ2dQqFgDTJVHOSilOHdgwCkM7Re
G8WPB92oGmMlM2g3d7+cQSVcW7bAw+cCwv0gvWb6ACnL1qmBA04vwAGkt+dl
eO8IHomuodTFnheFWg25Q9tqbYhI+qpsGhQSRHazP9hkc+eF6Wwpz6vEslvy
9qNvlp/hS/ygf5NiDrHF3xuTrfKaSRP4TxpIYZqlsek47KHZO9F6f8WQvU9o
B9UW3zCvQkRLKStm+JPjCLHK31EMY1w24NvmOK9D97Tj7H21Ow8z6yISBniN
PJ2YK1+H3ztl+CFaDM+oTzAIP3be+f1Pudvh0esYA8icr588vw8bX1wNbuHM
lRzS0LlfCzZajOUSlLR7q/2R+3kLgERrZWg1QLglR3A1uU1N1rttClEmvJ7c
rcoibZxjnj2yHxBkkwAI9gCga0u6CpL+OHb3xb1gdBBSel/KZ8L3GKuqhco0
b8OWyVoBjaVIKr2tIpdj1o53hDfMY9iNSurX8PA/2jBeQ+tiWHew81cZBgab
lb4ih4vUcU9KGpxmcVqB0QECryHFbnNGH5BKr654TL60Lj1D43MNVuiZTZM5
xdT5tQqIAhnAsKiyd9BA4qFlyLBMGnDTxbh7hOKhzstqsRGmrL6CN6i6wpl6
7YaWvtplyuD2vBWB/azntGaeI+Y8Y+3MipBNqN9FqNIO0xLiHSLvGhKUlvrj
HCosJh/Y9tV8KBzgpnSfZwvskTDVm0cFfM8HYnmuobnzCVjfcEKu2pKfWA3s
IKFkqT1fnwphm8HQEK9NxD/cB7Pk5X3IbR4nyuk/Sxl9njFvfPQ6nABzSHUw
19Z2Lz90DRarqjr7ErYKa3DGrHr2uXlj+3Ub7v/au+IzXB4//GSLDqgoZMrJ
cGE4k6zXk+fjFwBn1Cps8wZBJwz9UFmc7C8rDmkGkDfQCwNc6TLnkS/niKPa
6oApXcF1goFbTGi6r1TN5lk1JacbX24+WJGPeSPt9VgCzxJTTG99yNnMWdam
1fEYu7cIFztcQnfFhhbOlS2fb8P/nlf8O002tebIh4EQ4L3rqxnnMGcs2Cc7
mgWp45lvr+4v/m0P1WhXnFf8dU0XhDNuBYXQT4BmxefMAvKun1EozlmxGe5c
5Ky5LaKG9NplIw2O8f0PWTzje7rMBXRVeLTmpXpfkaYQFES2KGBneC4jpwMg
wod734ObJnEQdoPcrAGRmXM8hGyAuYx6D0TXvXyzvcjnx+uevVQQY/jb9NoF
ZnzfVigLHk68g60qwDbwbTrhsyIg7oSOLphFFey1zxlBtUr96rM/zRNM3h8E
d0UmzwAJpS0YfjkrSbDZ6+klfGlG7w8oZGekVDmh2xZuA2fguWQU7CehAciR
hhUmmz636uyvN4ewmeZioSNn/ljz9U4YlJL5c6ZrUdkZX9Vn9oi9ErqiNyjO
SWF7RhAcHPVEM/hihdjYcDE3D8F1ZN+PdFpIuVfvGgJiE/KFQBJjEtJszvPE
sRePO87rlf/GEA8gMqCv3YHGAEyGp1qbP+UEq+lStjMyM9PmEADg6nLi1AW9
zayuMreB+z2aRNSj5sfFTlKb8Ba8bHVbQJYmWGXYKq6Gut97Uu2lZtC3PzUe
iS1pU7RsL13pQbqOx4jDiAdRMOoKIPAPEGc37k9jDcg2vyGmx5Dr0HuRHlaa
1M08vDYLSne1Gb6yfN9k90DxCYoVcwGppobPQXd02QTUhf7VIIQGmeP3kvHC
OGayinoTW9oRkd8TxKF8MG1tWVLNb4ma6gi8LtNahqeqi6tcMtBhL9RuVjI7
heguUbrc5tqq6g0HwN7Na4qNcku4oiBhEFphf70fbEFSmQ80ysK84doQkgmD
0oL48BVttyWANTko+1fzqaUWam82Z1ln5GxAscPFLniQH+lpx4L6MmjrYVbR
Eff4psWXptHxk5Kht3NnfKtAFQNAXPqwD6OkD908hfJrJ6FFyOl6K/f2Tua4
6yf8GQ424XEo8LHcbi34FEodNH2eChIlpGw1iAOqMKqrCBWTC65/dZYb7Hxg
vWuk3Pmx7sPu924NmnGdW0YVAzbS/lTEsWFGaMsFEoHAGnaslbSyNShzQ6jX
ANWLSxpLg/HlYBO6c1MmkC6UIyUowr/1NQynSCbE0bH8DuTz+7nFiNnxFNws
1NKrFwT0RYw/LrqwUliin4bhw6GpHMxj/A57d7voK5gahgKc7C9OQiy8oYjz
xnlKXHrKZtbgP8i1OSRmTiTvQm5VIli62Q/MhqUaKBjoyIJG1bO1kRivxPOE
FOrJYWXxddp2xFCF/phnM8w15n0beALz1mq0cL/AgWA1U1OTs512R/Fj7IkK
SvWGz3rjwW1a1z0A4BM9HRrgMsBYMyBpuC+YuVsk8ZsoBhBHEUci9PcfmbX1
dBxX43GUatP0blxeHvzWJt2g4JhQe3NclqkSwnbiM6JHDWaVBks3rrPM6+2S
CxearURQyMQOsGirT1ZPMaUSzKxM4FNPhbZc7Lw7q405AOzzjafnifONoHMh
/dIeqHv1te/yxw/67j5uvpo9UK5WsQOjgQLozw4BDGNMaXSINEx4ZDFbdlwY
3CJL82/RAxYVjaULgp98C7Go7vUHzB+HIFGtkLmVzp5qKi3NpuNjopN4jXn4
JK8XAAul6u7W0MeOzBUvZrTvTGIauK1SjipKto4/eF4Po9UzdhCpFWZjvG2+
0evuTJbfxBKQ/sufo224chZRqtsQRefwWsGxUaONFuhjF2pxliSCecoxtYAQ
tT6fwuZBjRaXfh9hT2GnAKItdshKsHHbyY79i7hmbeTFimV1gNqOgTgNvK9R
XEbihXowk1K8rdXO78vvX+8Tmw5mDhCUlgIeTJ+vyKfMA2z4YC+VBh06A/KL
9/90vHlyv9i+SUyGtK71TexQmkAlliHR4b0fSf3xqL5WqRfRwH6LWpLFmtaA
eLeklUdpu1UCcj5c57um2dPYAkBJg1BPsmc+9cqfArvv1C2bXryyX9FVYz6q
I4ejwESp4myxGHnycnv4pyRRyseYI5h9yR9BJDmLyAQmMHE8yIysoXp5yxNE
MynuArdIaNfZVJsY1bfXq4ApotxuyIeC+ZLqiDVXPOgvC68JTL6cMPFj5PrE
vgD/6rv8+bDh078ZjZVCkToYajpIMAFf91Ymd2+66diYyAGO8as2sOj61wTR
u31Gw2uUUIxpX+IPE7KDVUltmhRlEfwE9Tz9ZX3+gw8esNds1ULyr4a/qKFu
Q39670+GqoAWZro6g9BYbjlMn5uZ0u4xYRGdp8RErXUIOdjKDXV38GLp0rqM
Bpy1/mR80WCR0zsLXzc4skcW6vyMlcUPEjQ1WUV15TgI31Imd+PInJjzLQf0
kkhfSSryndb5YvOtykMt7ihfscWkqqHwaQblRWSt9t8y1PTWp8LUmNVUq2CV
GOf9FyE+mgwmjVq67tIohVZtHlNPuflsfBl0ilTeJ6thuJmV95RWUd7Xpib1
db9rOdtfgem0N6wpkFwn2gIkowHbl+CHEvI8XEt9wZcSatL5Ws2hoXgfUGYM
SPscdX5bEWf471C9/qbv4l0qU9B97ZwzXsc/B5b5UC1dUA/iShrzRzKzZEJu
bBmeY38Sm2dv/uOGwAQoyIDVjo3XGHr4rKkZ8CihoLcCgQJnslFaToa2M8zm
0AYFdoTL2mAg6K7h536Ko3BnDI+lpKVzjzXzOkEEFfRbYHHfYMyOxpNY9Yol
LdUtdUi2EdPZWnShhQhKiY/89WtlPZPS2ncDWUE6qizluYGh8nEBrpk2wsiJ
9zrajIht48DhpzcC/Vubb9lsdnv0B3Zhv3/PQKFtIq3iaUeLW+08ItGUlJfT
Gw87fnNGEmyXQHKd1Q0wzXaboN9Bx/bN5/HHmdJdFxMFhwpcm8qTe3wU9Nt2
pGLV3KtV2FVc0J2y9N8PlNlDd3M1EtBoLrvlOmUFOXLX3Ry+lKVDC/oYqPYV
mja/6v/kBuI7We8lNVvYWTsi691LW9vLxidKnAAUPKzNAWA2HZqCYFtUV4Kw
aKfAs6nmvPpqiLUb0rAJY3hWIVvF5HqOGLlWfOIHFh1ONkYGP42MGvnLRFir
N/E6CQikGUufzASIe4SL2ZiyQEqFbYpd+NoSktllUzEUzxcFRG/IHXKoXZLt
sazzPlf0XoL6eFy4jU9t7sHwF/pJwaj2ThJL4UzG/2OJ/8Q/BRAW2UrK0E7N
dyD69IcfgEAsWCqYmw9OEdWz1SGceBtCwh8R2yMAy91MllsCvC184qybRlDY
xNqjxOlhBPvpnNaf/wXZwGVeoKPc0HeSEV6OJ0WG3l8E+INSR3yNHTc0QBra
SJ9pKheUTNuLAVSk4eCMlrzkFT2g5D2GDIo2RyygCjy/wcC3i1WeI8EjPNEi
TPCbV/57/sYpNhhXsGuncHfoiw/8rvUc1IrAfKenrd8d/TKVQF0X05Nrg4qW
8oJAgD56pI9KxrdcnERcR2X0ZE/BR22HEyXOewaw6jvgBPNv7kovPQXhk1Yr
rx/dH142AsxVyAsvMfKZl/GGae2Tnt8Oie7Yt2YnXrydZyXddr1J/Eh2ZPe1
WzakantNaocFWteMzfBFGdchNAUFti7+3UYnKUxzh7Wrrt+FPJDbuEIKOp4/
AHCoD3DCOcYI1tiB4uBNocVX6XVmJkGwA0dBvdg9CE7/M34U8y1B/px++A7A
x9OoKQGsFfRsUzRHuNuquokWhiLkOUEx/byvkDI/B2ACHmYEnfkOxzxLc37j
s41Go0XK2szp2Nou9DJAyxAPo5HtbibutyxiEeT0Aev9Y/Vt1/rLWy5RSDW9
aNY9vdQeuI+PZbgIhIkLPJiwYMCQUuddkxlNxZkXkK/ksfNy6W+fuzi7yX6Z
g2yqxt/NINySQGlEllEURiGvh6fQOK9TmQ8qjDtRh6WFC3X0q0lwKgGITUOk
vHPjGaq2v6lAfvk8HT9MaD3uy6Hj7eLVFAIjlEtLAzA18gIthNr62t2WbV4O
FhkuPQy5f6MVBEkF+ewyJbCkplHu5DdATGXjfNO8n1pDiDX+0+pK4GAv5KKp
++IklwRjJr3wH7ONzAA4fkqoxaQX8MZ53DknBgQC9BCIobPAYpAcTY3y4tbL
qmwDccZuuw3AkOrYURhHLOStB/3FnQ2R5bnuWHswBwJN76X8Wwy+60/LZB2U
3AGOW6WRB0jAEeQgNfDvPM+CNzWarx7d+oSt60z4MkR3UA/ItRqr7wh5XGIa
2xv8cFgGWWXuox3SU24CsCT/dcMwid3EcMURcLCW9MG1v4wa36mlH3//j6Rc
la42IfQowf0HFa4Wrf5nCk5rmf+xO1Bwqyfkr8+mOJ4/5LNok4brBWvKumuu
jR1HRSO3wtaG6j4o2vwOzgeo5WXJ983BAXpGifBVIWDYlyjwv9J77IhyyKmU
epz33akSZOnmxJQEeFYxk90qLkr2JzuGEi+ntpxKHgDiUBzXpLeF5diFgiF6
iM+h3DbWH4JlxBnzFOSkNZoeF61fHLNNpGf0+mTbsOWuJHGgmh8uXlPzTmxC
KVaMoacR/VTvBZmg5mSyhStKAPFeCAW5NhINVwKdy2py3+pe0h/yTzVpqQnY
GmCLF4HP/xKEsMvkuXaRZdmvpbu4pv2nlSAEq7dpO1mUrESuh0VjYYinMKUJ
PHAUHpnSdm8Nu+3n9NUftTcRi5tR3X4r9naMr8alIIbRXNrcp8j9wMR7GgEf
EEUUgR7A+jFXq9szcmJnDU9GoUhLE+mtuW03nzDdZ5AqbljnWMLvnkyC1Pgf
iL1IFmGpszv05cVnRRDlnSXyO+qOFIXxJh42urH5G5QBWoMyPtG1L7ca+v6d
hyY2+rbTG9HoqFZtyBiFJBfbGNBuexscVWQ45KN+4Oaf5v2i2+6Z2CJVFjD2
gWKSrKXEeg2y6dJn20FNoZ5hLfeVU+CYTJ8nD4J4a/F6W9Ul67xIotUAKNNN
adPdvq6468KcYMH6KfWSb+2N5AoLwMZKubly6JVRqglz1QPmJGUBPKW33US/
svMu+lL89PFJ3z4jWxu9eEbd3m4uEI87EOVbyYTTNtO7gdqW4k3WnF0WUUyh
0PdVXB98mJtcFVj+IPq0Sgl3y4N6qvbMHjUb81ZZYwRiIY7ukkkPk25qjw+i
Kpt9cW92uPNnki2LilfRWbkBPdUNyhY94VwdUVwnAzcEfNiHLB0ZQaJbLclv
/MkWp1+ijBv+65+lABnI1UWTjI4EU/oiJkFakml51zsoV7vaMaySV/0CbHF5
oIGUMOil1BtYU56Ab5JNFGnJt2/aeGDSVeomSLHJn1sqf5rWoPHQOcLcrL6b
Dkaf+2+3ZSza5q5+e25nIoZEFDpZoYWhwjVxFmoM7pgZcOCYAvDrRzRG8Y/p
BqW9y3o+prgbaNJedOqSrj4thv0eGfc76kYf8GLE5a5dqziYxm+msSMPCc6t
1QxsUpyhAspK2Km1PbbneHCoWgqP38lxDsWOz3CerpORyUpn7zRieT+isZk5
NUBDCIgRJbrzGc8dOzajiciQ7LWOj92h/lxF9uO86uVxmSUfkaEOfzMY42y7
73ZpbHybg+rItoyZeS0B7ysCIU+7s2i60j6KZkQZwWpzeOEfurZwQWCPuqod
+gJdoJZj3KTbeqbvjITtd593NusJRc9RLRGZ5mfgUPzscZyFBU9PO5J2/9Q2
Yu0ADk7WymoA7h9HrT6Rtk/G9gImJKvgihRd6gssBsQr8UmNLQu1T+Nh1tn5
MhpHst/Q302GDPJ1khrBGxY2QjqhMAat2s5eEoFDfaZxT6fJIlfFSmChhApE
t1EzqxtraNYBiPN779jeHU7BowjmVFjoKU8V/QFbr4UxQE+CQXcJOeqvrGD7
M65Kq4fhtvKidS0VG6AGSlA/jyCdpNNsS65Ye6ZWdA0qYeDi6dDTg57qSDjd
eNHOEI+i54v5XTaRyqtmcPfWd4v/14cg6qtswIdJVThvmnTJXo89Cm8LyFHr
N/93kLEGa+7f2xWj/Z9I9kQ5HqPycK048YV9iLyNLWIe2y17TFMdAfcJXBiV
sLhJBWt1LCysNUQo5xBETpYidx8pqLuAhVIYZZhUXNI5PC0afjyKZtzmVL8F
K9EQwylfc50sLeIuHJ9AO+ZwQ0sTc3GZ0a331xmzE2dz2HFgeeUSN3ctTZUV
gd5Fd6rVeI2Yszjh8x/QplZ6ElqwREIjrQ9RUzaP652u/AIBZZgNV33DeVJA
gf7qoWuXFVqOubfWSSB2e9vbyfncZK5i4+eC7TtGQlHMxP7dUz0v1nPvqg/j
iMFU2wgUXQSSf59vhgg+AazWyFSWv5voCIGlM8atiQhmNmgKIhfwLMz4piac
ydscjWLzkQo9Cxtj0GBeIVuoialom8iYLiQ0DDLzxNWQe5u/APw9V5UhyNyq
x/ephwDhoxQf+fwiKEsSS3qFtBN0anZict7P0O5P6KfohS8JzpsMSnhQbKDf
BEZPANcbtIczoTdGxcdSuUF3+Z2DDNpntY9aia4wsGCXDxd994vqcVky6R8s
f+yaSUWvcAnBXKFdQTZe/3LSKt6ls+j3lK+sxO8bMJ8qs7ZEsZoSsJw70lwF
7LVo4uJ3ZCzRdIJHOxicIkTw+fh/TCrJiq2ufIFQQ+P1quIP6QgdUuhSXmw8
1/H9m0OmsA4cVV5p/4mClrwLwV525Dcp4oWu3FXd+MtK7jRWSgndTxdvHhky
KiYRGUdw060k8climV52YgKRruLJyzWbIqEY6kjpTCgh1fxKPtDY5TnCNyBL
DHiQPN/sQB3ad0rHM/rdPRLteKUmkH/l3Bax7PWyZqkJRAIV6VTJjkVTPc08
UsEETWZJ9Vo5gkrxRFXx7DGmxeXfNkTbt6KF3WjJ/BSuvKyb+sU8uYQv2dGl
h/R+Tv1QlfH6n1FUXhnmv2bXAommkXrbkvyAPswefX9SQ5it9yVLN9Y/EnJ6
cJema5JtaAOiq3Rm5dfFpcjNbDd5keagp/rXMdX798FzIK1yCqVHl7E0IGo4
1OS1cqjgcQz9xfZp0Ui76HhJegvEmpfT5cVAYEG6XIRSSXtTYpDrcNvuvJyv
y2k/Pq9CeKT674Je9iIR0DGBeCUAPpFPoZYk1YkK/HdYAaQHSzwfSdkskdWb
f8osqbBQMbPfskiTMKwpks4n3Kw5ng/Zjy6xigZnuV+mUYfqoAStSo0Ckyjp
vW1fr+BnD7HWvIkvLxNsdDZbzcRyvSAmUvHQQ5yIOfA46+QKMSHE5IpCwfvk
MAYec4OsOedoIxOIM+XPU3R1FnGTflkvDn7A+Rsb4X4m52nWCkRaDaJYSbCl
5uY3kqgPFF/yt0M8pUSLxTFkag/Twk+7noO+aEwdDPzIaZdD4oXp+9PhNSYy
hpoIHGyX8si4D6AtrXWVTD8AoCTj2yePwcRgTAFxkLPAuniwdkVAHbiuTsER
/RNlCTamyJITrLB1NzmCt8yOXHd1mZuAIJVwkTv+Rq4/K3JFtySJRQIw+Yyw
PnbNqaJxaP7uSXvjI4zHN/h1hK7o0gSsa8knfZ+AQPXTN66HN7FBjjYLE1hg
dSbzXXuqJliL6pMyJ/Armu8BtoRRjwQMLaeYEVoGSUSMVR2hGIPCPNfiw/eN
h/u8yONuRvLXcpqn6SIuEVFJzlYJvLpY39qqV+6/c4hNidb71r+vfh6VtaY+
1x2GbVvZ7wEelSiMNwhtrYNrUcgfqJNcQ6irqSBGkAJTn2YerOfX4Q6DTATn
42TA6q7Ciz834pLR+YjJTpyAWZ/GuBUIawZ3qZCiBQZxEBYvByEXP9sdbOlz
PrL/Odm32yUYB9bkr6fKYVNhj1jbANdD7qCeR1oOPjHMPZltmF8PgueLwELs
QS/u80Ye2p9FvB3Bnc+nSo1D1LhqxNS0YUd/XAYfajHaGymw0BES72EltZyq
QrS9maV8sDYDFeuwqGu9hicCgtEVN0E8HM9Mw79/4UzA4x619gBSE/A9+62j
ZD5x2/McU351qa1UDbIlR0/BEE6PG7hzwxbPZlw/OBu8z6rl/AFseVRh6fYL
zP71LmB4A4JX2WGxPGjTgWdZ6rP7rZ++NP0HZiRTLu1i0X22QQG/9fD6pEGy
97Ai1sXVXAbSfikD86QzL5yivTTRnW6pyWk0V+g8+Wx76lUnvFyo9ofuru2j
wAcPz+eQ2GvPUTlGWRwTtglxqilsil6oks/Q/NffH9bw4lJA0kYTw91yFOxt
Zli5vB175A7tllX3fzEm8kYGMe+cYg6D9pxHcPZHWfG8k/wpuDy1srYe1QA0
4Jm21VwkJyGftO5W4A7csFkMWENGJqiznF3u49ZPSbGZRMsiGQSSQQgeeE79
e8RPZpyGzgFsQcAskH/Xo96+ld30QrigA2CvVXp3ZVZwkeK2SKbzLDLVbNxG
CSSriRcVB+oaXz3Gu6LlpF+NTCv3LlnE4gOQ6YZEFhGV6G5qQllIez9EGk2X
P/7i01CpNQ9XiUP/R89t6UrcdTCv3+cfHjfaKcgF23LFj+hz8DGqb46OpsE0
LA4pgFNQ34LarbdpABP3xQrs6UgMKUP/EdC/6qoHosSRjA0oLWXfOLiHZ+yi
qmiM3T9bONeuWiDg0ohONvK577jUAb6mOb8IJR8EY9QUxUUaR2oKXazTdQVv
6r5H5zBc9xPVJLGvLoiSWHnVG+1iGz6WcP+5qeACmlLJT5aD9vg5BXrqGGnG
+kPgVHdPUcvAg5+tMGnM5Lghv1fpGGO9I6cF+OFsL3B1Q5jmphV7KsiY0BzQ
pM/o6ZftzFcNkfgoWVv6CWjU0LPWUmg3wFrsdjX2ByS/mtbnNKlGaLBNFaOz
qJRvp0uuvhG2NmNNqLEneMT1fLQ+vWXVQiFnOdc04i4fRAmShoSqeBBJCYGY
ouxMyd7HOs5d96bO8IYBxdq6YzPbHb7Lt42eRvwqO1l/hn+xYawEr4ouYfuA
aoEPTCvuBPv9A/LHwYos9hW5DK9As0JhWG4iYwnPeV1u+0kiflLem3baeYby
byKGwjkdJ9miLgPy1ItGn7XHzwzTgIWTOZ+lplwWiOHWxedr2xJivoo/jPHZ
8Vp9hOBSuos2kXeS+ZwZQZ4DAoa+7Jf91IllSkHr8ICRXw5r0WqqWj0jxxnz
Gfmz2Up1Ul9WRRsVPxi9wGrV2t1xrNH70koFgVmJLYL5wJ1noqVdunD4ShTP
8RoqY/+7/lWnlw+uJlk9W1ljY1B8LlDrTnC9zI7Ur6yjs1jyDtJxxktMDp9k
IKiEWmqjXF+6+aB1xK2FM9cvYDIsFsaBWsxM7lieru+JzMp1Tgih99lDYRWZ
66j8doXw/49nUtU2nGBlv+/btS8eJ3+802bP04wklvCWgWnYHVsAse0M68CY
FMAAbh3HAr6vu44bLzAVkv99Atz3o8yQTTrkJ6EIkfqkC+ZpPW2b4dJRZ/zh
kxgyaL4UfyAICoXm5rOb2c/z/d8prC6poS2oyJpLvxUg+1PTNRDv5H0HPbxT
VbectURUlWAkRw2hXMpBSLsrI++ntp09Ys3uVddpeNIvk1Q4glDHsofCiMhp
rYpNJWc1upBQuC0DIAg959SdmHfrB2BLNZK8OouZXj9LDBUsZUMrkDRv7fRE
mr5p++CH/ZwVPuhzxaCY8gfmDM+RiKl7PrwdEWPVInrlYf6JkXBL3WCFEGlY
P+r/deLS6hFHo+g0lbVYKZ4AW03IortoNDpQUfd8iYNvJEvOd0eMDgA5nsZD
Aop3282XfJVjgyOcMg6nKW9WwB+hD7HKE+vRCgtfkH0w86+pkOR4xDmo6dgA
GsQfiH72Mj9cHspCiFC16oAMhNzfUY6io3xjNzZ/e1yCuVnN3LKRncO2XP7C
IuUeRZM4ZyyeSsdkDpk2ARJHBn4/SsnWJjB8mYJkBwS3Tl1tB2FlBh+b/dmL
J3nzQbgj+PGOLfEkU2H3OQ29USrSaXA3PMlqHWkdCMriB4PgKYWiRjV7F7+O
/GiSx3wsePWf5HgTeE+TZpqrD1zms28Pgk61r7kOg/52TE8uw0wPhmRt0ksw
+YbFkEdjVkyW8Pv4bRdiMX/jNDTISBk4FPi4L0zj8FTJ8Kwe7TLXma3zpXjg
pBJz0BNDH+IF4xgSNOD+MPXbgatAPBOCcEl0QKcWPvWyk3Adz1i4ewhM1Pmw
e6TC0z47bbECOyTzfPa8TTgTA7beREupk+lgOFqYsHdH2Z8OVmB0T98LyF+n
KrBweV0GTeC7irFEU3fmChXlin07hgef8dPwqDeaAHq5YauJlgVS4/MEnBme
u2susuLNFkCmLqN0e5en9ulPKDslcwAAhAVeSuBO2He0gk3f2MgOXNJUYu8N
GIL0LOyIIVdF4nbSTDmpxpqtOhlbORNHhJ3kFTYDW+twjxS+b0o57kxtpB2R
1hMFIgCVb3+huUwEKrI8mDo06ajYr3aJiCzNmq7Zud8rzzEaHgCcf0wgiEdK
OeU0e3gsoLCmUAPHwEjRwv4FWtlLj/bNqWE/5HQWO6TxvaFKEoFi8FchAMH6
tsTM3ZzE/59tJAzkoZpCle0qfTj6Y87S6N6fYQpQOORURlJ4jZ4MzT5EZaaq
sNQg3aFbbo+BRgpgMTMgM7x6l/AFKuTZNZnmsvSUy04/cucVLMNXLUWp8lhb
o8Jqx0+XFgee9nsJKsJz8qVeMiiWw9r1EDzMjDtEWVbNI61QmiDwFqoQcsRe
ThcDZiGWxPdTJl4KdLPUcGvVOIaxwUTyN59nsf3y7hckQca60HF9QIv1Q8Uv
u702Zia/nA90dfaEu0Dl9OLlqq33KUYtRVMA2kyckDDCpACpKr/9xr9XSd3b
0D+XQPHm2Zf4oN+PT7GdeniBrzJyQ86AYlOE3dvI75m99e6edW5Jm9jFmAC8
8YLQuc7ziVmeLJqOJb2WlfeqkunRaYRB80xvfdthnQ3LCrF31T0kMdMv6jT7
E7FG7FB3AZQBO8mrFFetLO3J6c8GtxZnTXphR0UT71j+mYIdKjhNftw36PbN
u7BgB210gVgMb71pUBKbECJTEHCXlc6cXuKBW9UireiU8JfcSTAJO9qljOHx
1cLEvDcduDp/QNHibUK5YlDf+dj57lvrKMphXfJnZKNxbGv/aJap/KhlZpKC
f+kF2OYSnXrPAoopZrzKgdwaHMO836PC+omPLL1tjuvzWowfX6moKhRwriPE
smFoDM1Xx1Tr8JKyr3uXjCYtxZJzvvQUn87BSkFeOPWIKZm9Fg7s0ErPOBPc
9CMQTBSjT8mqPqY/YzD37A9aBdJvj+qEKD3nFm6fbodydkVFD5JZvqjD8bFG
tjsGToHU7XJogYMrWLTiiYXUaf2PEX2nHenwpV0zjuGnA6jvT0oqAduqlrmc
QFICl26EVzmr3XHoD8aClrjr9lUXACH8Zn7VAt+1PEVZOjeGFV+1kV8nRPPM
PCmu5LDOI5Op4QULmBgLB5/gYyyVeazBhKDeCI9Xb8pq4HvtpnHL2izKUquw
C8bcwMBZ+kLqrtiBYL2R559xXypeYTM9XGSoFKh9ui/FZphkVQTcxFOV8Ris
e8q7ZbhUi1vKhGT+Xqy9w4ypZ1cTFkStp7LZL2jHeSzf/7q+88tAWFiOwbJe
xn7jDFKXs4HmrQ8Si61zpQVXLoI9Qovl9R1SizC9tNyyLfU/c3KPhxnJNg6r
10W5vtnLEgVXeYILijA9/fBKw54Iw9bg6yEv5ssLW23FIdoH0QQnCZxYiAsU
DMSbBofxIuwliLQPN3LVVh5/tTk1lnZWIohv2IP3YReyENlzhdAoUC4pRS+b
GRVv7NDnKqiW/R6PMbVWTsHIMJDKmylaGzDjVnIk6jgoQzKZTKxwaTfyNva9
emFJC2hcvtjE+QZnblL6gnIVhzwCLxmRkBeMrOFah9VZGsE511I1aowuzsOe
E0maooy6Sl4rk8sc7X78d5Cr9xkw5km+CXcUJuw/Wxsgg75VyJdJtNQtkH04
umGKMFGwnJJACRTFAN5Fs2KWdnvr85Egl2yAF0O/TDqu9z6+H84evlKKRJQw
tk3CFTrzaPqHcGRzbNSCM98cLjmhRpNJAP45yXysXJpe1YX693VZqqwjeNoQ
0hEg2FDNLFxfE19JdpjN4NnEqLY5LhAreCe8yOITgdMKosEJg1nR31EvaI55
joMfrSjBnShIUhJbzPacHJzEb3J3WAn/+TzMWF5HTq0n0AD/bgqfx+vbFOBJ
Bg3QiLvWO6CcMipDstYQ06tL4LTHJJeObE+aNX74VMREkPWasQpGDWDH4cSs
2Fss28Vg5uuNyALuJj4z43LTafHVwd9e/hRQdPtKzMSa8AeXudcGuTmR5U1G
aNg+hzuvDvx2Y9auuLKgTTK5ObclliYgxRQsAglpCz47eEu2Jjx0IVSl9d4X
5w4CXjtO89XiSp8sYPlFfpccnUBMTUTf4nARu7RiyAcSjq5IKcsT72RbnEnG
u9vHV7RgFKy7+PWDa62rLzVUwxZc1d1lPsxGIc9aee3qRM7rNyzDMC8QkWF7
GTfZWm+zDh9POMBZdPwt+nfHj7oiwnWV5X+RJdU3IbXyCWLH92xd38EvyR98
XBfcCYuKqIkzdDuugmrskCFiR+v8NXt4dPBQMRr+kYhwTbA4H2CdewNwVZ6I
eg6tE2fCghVSAzTqaZF6+jVZ6r31IQmPXZUUJdO0gRnlhzJ1qGiCaAiWFVmr
pUW0l9D6CuAFBTYS9GRpr0IZs5UmJMzZZrnuIjv24o3B3mXeFaxTZQ+yhUp1
DtHFrh3lh+y1xOGjjiLn7jeAO8dg0pLoy25+b5L/y2/CQgl3RXC38u/Gm9V5
DlbGUNWDHdEJL6VtfgYOm72i84A/X7TjPJZ4kwziU/P3OkT3h0V7IrmvMHkU
cn7uOHGPgncbgt5fGBMSncWFP2yT6pOmtJImM/jMG2+N2aTTTOvxsOVQWx6/
+zCAwiKVz17Xwc/1AyS0eFItT1WEx9d4DLEP38pKYe+1paISpC7qMeejvJt5
R0VCetGHZGPkM0sMH2qceObypCVyX3pNuXdVrm2XMBWIj8gSQxfyQ7DIiM2y
GslXUMjF5t0b7Sd1Z4R1DTD3Iyt/z7zyfMIc+HwCCQw4mwRoPqM9qo5ulxGZ
TPqPdzXaQWrArNSXJ86lLAAmvZtlw5OVZflL/GT4+dRxWa0+PxnaGWsGcocK
Nw89hJMXQmAd8wsRk0i3z8X528gmQaeJL1cD+qOi7XHZ4s+xh715Jv505yKn
vxPZ0EkfrhNidxVWf6CJBu9xC31gvY00sB1GpU/lqzmXJc2pCJ7KISy0HAtl
5H4mEntzufLcZy60qxfgvWz1pVBl2bPDbDZiu7b5I47bgkxDcP6HCWAtSyAC
vI7KqARYQJnsQaJaO6g+3Fxw3UUGnPy5CdXbMjGD03JxwJFT9ukdzYIVZGhi
m7C6KFQQVcVEDD4iJ/Ntj1ZoLK+knqeHQt7wmyA9/hnp+xuNPzYM7Nxt11GG
nBY+j+2VxjpFOv3M5vYfqBSPH0FSHvyfolzKZYU245K39ixw8uk/oPg7LECH
G5Mh2//cuqTjltAZ7QFU0pLgJpYTUmnbUJhak129U4QAHPr/HU4NFwqhPcY4
iJeO+5pVu+P7IX9W46l0kCeOdDGRfaBs3/c88o/oXmcCbYwMG6gKoWLUAIhQ
RZIVNAWy2BFh4RnReby0PlOaHGj4qyxletFMvTyHWABtF9xAi2V7pyuuKrZt
WEW1VknKfGN4b1ZnGnlwolSHrdTFDpPKv19J5iyoX4np1PIRKlUhrp//j4h7
T/x2i2tCDf+vvGsKxM+I2kp2gszsMCt5biNUrH8hZZAAekjrsB1hLBlWX/FG
Pwx0POkMDRzasNaN9PsBtoTWBNKCY8GqyhgTPJoKi2gmDPx5A+DfaiWA9IrC
km5kwxegWCm3Sl8pjQDuWSu7/bdnL62rrZqOGSvgIqgoiF4/mpkHBjITDCW1
GVfuALn87JzKO9OM+SMiYDHrx8HUftlp75L2HapGJUmXJNLZciplIDywhMbx
I2i/jQcg/i/FKaUB/qjJfjaZJQfrzgzth2Nz+7AKnYAoEA+Fc20dkWewtZDC
ul2BjcFUp/3sqcIzdfPFNlqqPJuqk4otHnjivuMyHWEAnmdRn8TwuC2TFEtf
6pwMxuH2ujbWPqxUpvymezBRiBbZRpLgBPypPaDhVfF3OPmX9kd5BnnwCPjc
MukyygRfDYy6/ghRe5vE+PW6raaPPuGYmwVp2EAB9UB3PIsE/YJDxuzYpMb/
vWrIsRHqnf5lqhzvj9icUyK/qUlpLTY8sk5o+U+xFvempkqjrXTNiVR3lGuA
5y5zuP/LOBsEo2Vc/xvVp88dIOBK1W3Ji1V2aLl+Zv16gGaQcz0yPBXampI1
up7EyZ6Mg8tTBEi0y9Lrq9sNDRUGwU/T1g4fbBpbwWyirFhNFxQ054uQjO2P
GHTjTJaXUCiSXaUHYRftETZYnlhHAKNUZUDStJKLJNXDKlvTWVq1JCE3k0t4
sez4zFzkmMWxzBXXVevnzxXi5YTWXSgAALiruRZ/qarEp9oR4+uGx/NORMZU
iUBkoLDdyyk6l+mZ3ucBuukWq0I63RoKMM4z0peEOD6hWI2rZrYVPsunBn5x
7rXqL9uBJsxxpLfjPdbpSXg9CF8wFtV9LsqFzBM8UGlRKybjATDbT6Vb0FJB
Zo5Itodik4RM2qG2xoqHk67ORpeRQwx+Yt1aSDdKweJpBcTbCoZ30PMclV3c
56wX9B2/utDlid5nm/RsF5DM2cmLYCu/cgMqc3qzVhJRcovrxJMC4w0Pa8kE
Talm7x+U4ZYdancPLtp4nNz8dQ1wFFXyyj2UnYgBF8XdaETM9W4h6hz6pBEf
58VboOllHClZ3HKUCE9ZLcarIjI7wjTRmLLq+GsGW1JpuAK0m4rTSbm4jDRz
5fIOGBkczN8S3sD/BR/UjfXR2QKWm9JlqcMDd4WCryMNKsT2PDBvznqGINr+
GCwZ4Za1CPxzNwEPDJqD2k/Gdu+hmh34PT1zZfAV5QIc7gXYEAjOpCN3wun3
c3ApsC3lZLbAHj1ug4fWQ8xVdLLYF/16iqgNJOVHZGIXpJTewV3av/AVs14N
y/31TTnP81nFUyTuhtxJGTIiC022652mKZMrsE08T4VQs5rmMwg9Tj1UmkxA
Cov2anS3TYnHeoSxm/M1GCfzxJHhzGmvl6h6Fd3e5Bn+JVjBXfTjHRRq8XDD
vdMkukQbOAAFJi6b8/m80lL+FEKrJc+f4+dyry6Gt3WqLCiZWkssOYjeyW34
0UeasDSh+iw2YKmm2WTkViy3jAh4dOtRd6bi1l8ACw95AehhHrC/qeEu1ORd
4UcGRWv/mrNdeui1vtKrO3mpsj2/sw1CSWRsTGugZOhOU7du12EfSWDOfHuQ
F02PZG2c6O+cM8cCiVY6ZNMouedKnT8gnkj7c+EXNVkx9Q8/RKJxbObsvFVX
L4ifRpAU4h/VQsDfigRiU2I4vha6D3qR7SlktAVUPKLsnBu6LUXFSHwzXzFR
ccLDHhFKS7xtkXANwjsbaQqc4t1Zc5kNXynORsD3yk2t1wCjRKmPVOo9cPA6
G6o+TqAZyUdov5gpUP1ufSO61b7vuKeKdYT+OwMqTVWHoXTcfEhP3LpHrDNj
hRkzEvtUBSocdbCNs41//oKiDu9VrjLpfOq2YNUsLEyKsXN5Pcgvs3OX91aX
W5P/1AWdJ1qBLpCVumHBJ2CzhWv86h7J2MRjt7bsylvoPs2lbMbOyKXdp+5x
UxygUC86LpnR/mfmviLBNPP3ni3mwZVx3y8BwS0qzcD1Bha0XMpK5UMv0DJh
i2hiyQSsqR2KL0gWPK1t7I3TiOnMgstOBY83UvvTFzMWTu2dlztbhIWlxZDF
FHIKLnzMv+w/BEMclHhda9flPyJU4cwnFSkp5Q/srvomL8Qb76FpxXWT6CMn
9sHY5/fp3vFZXoEje7jn/bmFazdaXyAVQMjW+YRMp1E1NtJwKWESde/yFfvn
JfWTvK66MQBmSbR18B9/iTBKhmWWdTspx4ZZ1MDdxwMlzKzOiP3akXuIA13Q
/L76b7btX9ol/D9TD7nLLsprzptPLQ8MgRn6Vsm/aySy5VCbrNCb0kGo3YWA
mTqAgYfJak0Imb89nuOzCwLD7NVlvo6fxQwJKmYJRAhcVF0R0GtclLp2/Yt+
QH0ataQ7pc915o/paQ5ExefPG7pI0X/w+mXZ1A0uD7QDLr4njQfNtQhmKGnf
GVfQoPiHxfNRmLqlZhmqyEUjcTViy2L5JE9AlPLsuaTJxSYWFe88+Cq9kVcc
A5q3OD9UZfOOE1x05HnU9c/mVQNkw+KQFmsqSRMTxc5FlvN5gAtWgPBF5hrv
hV34zA2TCuwrHebAVBxqnkp7S9zk5iwVrw8yu7kpDAKV/8PZkkzkkSxaUBqr
ociw61w7MNgvs2HuguxtR0LjWk0MfCxNUavAqUjd3Yso4JIn2rXHnxyVuWVe
qf7NXLNXPqFE71uJ+GMv8+Uan2l6Z6BipITshZHqXE8j3eyGGE2eGUr5LScG
EfmS2ckpOl+kOZ82m8sOPX8fSjaJVJZ28OtkvS77HQDRgdteGdEjS4xeyvmE
3KmdIoW1hQgoPBE4w9i4P/mWnBJEvHadcd8nQliXnyR5yA1j9y/k36a+vvUw
x/ul//h2sOYWSAhubiDxYWPqHPY4E0q4Tc6bZJBKkO7/IpauK+ZOY67zHo/Z
u18Zc9N9NEIb/0eexoRdGlieA1V7cOQTBVQbsRWnD5eRaJA4jzcymsjveKrd
PSDV7yM+TRILq4mIkrTmbSKCKrdaXSH5fmu4OgPjQ7fj8s3s4TsWcx1+gX2L
YbrTDyRvyH+1L53klCKsN7B+RKih9rkKznJzRTqZWw1VoLwfpwCwUvXkrSMQ
KL9qzgiAMLlMDYIgkt2v5JWzeVhPQkWcyIgehjlLmqf1Wb/SScANFpT/8rvM
J06SyPdwLnMJr8zFKC1e0S1EjHk4buLA+UGzdL/kOfBQOPO+oSNJeaxxjQsK
z8uKeZz2PCpUu6J8oLqEm/RhZenYsfKU6GBjKqDtC2tRoruBTxd0BkKNSe8b
Lw7TXL8yT4G0SS9fkhh6h4e9iQ4bWyYxEX+C16QrgwE93IzD46pJ83FJV1nx
aM+8mqM1K9BNRY+AjxnlnoZDGz3cUt+46IQpAWFPlvxOgj0LiD7KRxxSm1EV
ZHYCNlh3Ygg3BDFj0SNs2QQMUQPXPD+d2S6F3p6TkTtL/o5wBzM1h3e/W+d9
mIUoEkmjBE+L6j80MDBngj81DqI/Yo7LB+Dzijlf+tMZbgFPBmYmYH1DLjM0
NgxM1b/Page3IdnL3Qa7SShf2E+RiVPt9gUMjwROvEYAkGBmtMsxbI6VYPCm
AZiVeyyUAptFx21eNANimvLPF+D8h6wOqTIYl6nxZ9sSrTeBoW7G5kklDobo
s25V2XxodFLlcTIVyoPKcg2dAZc5R0EeP7TaU1xJQD3K8zzwu3xtBDf+3cjd
awk2np+zj3S5H97rXvUA+3gHXkWS/I5v3hfIY87t3uTKprqv4JTCh8lmg4g4
5TtM5Si5YVfEn3GDlf4k3MUrBZsBjMqyQm15UK+LvJZcem4OMtNVdUT8A76C
YAVjRxMzf/ZogiUiteTHswSivVriBMz3uyRInhMI0DD9cFyyc4brVIMaqFI6
hXIRIoKPCrG7mOZLm2kakukGqXi0S4OMUEnel25+jD/cwyy0O7EmUfOLzqXO
b4bgOBdWnhBtVLyHHtYkX4vK/uHXoNJjXhB6bGx+IzSNpA8zkq/ne/NcFLp7
B9qCzk7L6suZeEHyE9ulKdaw7T7cDScCHhFySVKAfUDqteEzq+qP9Ipqq/1C
I9ZOALwoRH2Lov4k9tkNyteVP03NoCr4CUrLDrc0H2ztODVpoAttzuzeRhOT
AXB9Q7pl+qXjA7QaguSGWl+at8QQ9qz4bsC38wVUvDXnEWDOMl8/Yno2+khK
Q0LlpuETxPW+KnpvVs2iUWDqdxlotEzRIb60xnaH6bVteC4JXLTuWiytBUkX
TPGuGh318oVLrxLl+XSq4ZzSTy6JljCjm9kJTZ+yy9aVCx2d2wTiJyRWAhWT
0+p+rFdhwkb6kppYVIfJlQec+cZjrtRWF5SjwFEcTW2J1SdmmszPBStJ8jQJ
0NhTyIEmnzUFJ6TJADnd2spLcu/RYQevG6LOoVIcgQzf2WK//dlWkRpulhSe
9gXLQBGpMFSk1ZaAmWZV7RX/9k4x2fLb06445ubFrsEXuSnC/VcKBXC7giZX
AlxPcf2tQKzdAJXJCyAethwFwM0rW/XdMjLfRKVPcVXlWFw5fBZGOwj7J+G0
y69hIQtS3DdeoEADOAxYZP2hrdqAt7zqB2w/1Guvz4Wo6tSH0tNyWFRAp/w1
EdR25JJscM1RXmCWEA5a9+ZdaqHm40Jz3hsp1BPgULKOjxl4qxyvmaPUda2w
67OiMC8rmWBRujZeyRoTmGKpIc/bTC5yOLHG+R/Ze8nwgBPRQ5eBbpS8MYtt
WzuePhKm077MHAQRQiEsPNVEmO9cOenN5Te1RS6edNl6o1jk5+7SujBqN3aN
sLouPmNiWb/krwXfWC6wF7T7s+/P0hG/ZwObzT4Wflg9iC+tHbHzc5gde2+e
LI49nUl1B/djrPz9hqXXsbEFBXmx+9BUPIDXoVAGPNFVOcQmrh+TLLV+9gyG
/0NcStTvWybB4mCeAeGQ0uBXgdoyFRiTG/Lq6emIwGL33svqNgENlYnxFMr+
5ejzGYXP8+upwXl443/JybZj210w5kMV6lSMpl36dOQ9nX1hzXWV+WlxuLGu
3KgJe80nD9ivRzguFLyPwbrY8qfBpsY6tDhS4zs14GDjfeOK81emxXMn6Lro
YSz3BasCvxzWl35773oC4T7MygLGdXqk8Vjz3fcP/IZVen+Q71cGqqmnDSYe
QZATrSrYimPvWMab/A6uWOCs/XfCSVea+0ag9nBkTdqUArYEMIs5SjfLZ0Rg
AtBNl8JpisZr7JoZFPyMxNLs5UwCfnQb2xetY/vR3XCxwrVF/HpFoSI7txoF
VzmqD/jU49wnBctkmBtqD6TyPvUaZOVpIpMFJJosT4q86vW7HoOABlXYuqAA
93PyRKovOwpoO+z42w5eaUNKn03a9h6zwLgnjcPfp1naQWgTnHA1w8ito+Cy
EkVirP07wl9/VWzHumCUICbvnqCW1kOdqkboAH5QmRI+JBTqbE6pWyKLVh3S
MXX0c6fWpjqP1g5Pcm7cRhu5VoxO2k3Dj3Vv4wuJ27tSrR2gTkE/wu2XQxKr
RY5qjHDtmSji+/NVldIzpbu7taWherntsZ20Y2MYdkYTj4QvSQkS1QIwnRYN
9BnwpB+rVhgcGsS/9PajRlLRHph2uPeqwsWxXr1h1NJWvhvx6M6RjMC3r62c
ve+J5/ZSj0qGja4DdWNPkp/K1OMeLYcgl5mZAb83ZcoCurgOPsxUTnyP+hs3
iT+B/Yv8vry4GwreGsN9Nw7svaSN/k1FxCYdLBdy53+Pq1m4PkyTyeM1pbFp
/0+y/yut5OCYLF5ME3hQBKK+HqMaIld+Bt8fsWcYND1v3oceD0Sh2JYRhadl
BhWCigSBU7V4RdyNuyNEgrEDcU15X5njdAGcx/Xtq7Km/MW+bRgT+dismCoN
QBGfNa7VF70Mk/4S/m/gMR2XdlcfY9lfX8vW+KSYTNexiCvUbW0TggqHYMb9
fk+32YioD3OMFoyTiTtfSrFc8eNsjSQ7RSlG/83KQH7BIUIVlVNHbQknZhUg
eHp1zivtbWXS/NH9r1KObE66uma2q9Qp0syRQ7ZSPdRQy/TowMLZq4fnwxS8
q7zrfciOoVVfZP6iLy8PoSxUofmuj8Xrf1nNCSOZ5tRQaHr47VJW8ZMYthBs
Pe5KRfvaNTqFHAYQCjdeRFCwUvoDve4DOYZFnImrlxDSu4ElH1EITo38X7tf
NeDt+XsQufZdYik54Z8pfh/nIkh10LR3Jj5KzJEOU+OlijxF97WLSQdjJNzo
ExJ6nROFzZfRwjiB/CYOu1z6feEwNhOc546zLV8qWcc8txRTV1mfYn0kTXVo
9fGc1dCLOoOpgC8i9WgJc4wVcRwcVyPttl3RRBUCQ/j+98ipnq6UuwotEoFb
PlCcxSuVX4nwVA5MTWqa+4btJv3CyukUCIZru/La/p94OHlPAYtxS7zlArFi
uNV6pUmR966X2Sulu0bfb4kHTcbn5AS6p1Q8qh1x9g/Rf3eHVMRCwfiGt5GZ
CeatYO43m6wqAOrXhXsaYJhN9XZ5pY7m6ydWOJQL5u1YIkJobVq5+iEfpK9Q
nujTLlgeuXMlAnhKTXIxHOKCuEID6nwO+qg1PT3+mS3op6qn3P9+P3QFd32t
6ozwvuxXvyT1KsCISl9atHGzHkAoFeHTqg2r7d6CWI9Gge+fCy4Bt8rGoOrF
ftXT8Z6d8aRfzdReuIHBO+JmgXcU13fDsRiuwbq/NQf2psb1w7rKwQ0dVPPq
OsaQU8X9iuWC+7z30cvbAljETepFmUHeD2eKY+asCRGKlp4go6ID8odrywJo
E2EThDsh4YV1o8PSU+dmHSV5/3CMWqmZx6Hil17v4RFeVGjj+qAo/syUZmuD
79MyWiIc3aj7NEvHrvz9Cib48GNPz60RMU02FE7JayR47JqBo2DTRnJ8K/0V
hZnUSOCg8LkLlbNaRBfhTX7gX8AHwS8TRo8AjqQ1T+OabjrVRcUl/PdAIMmL
QAVt8dQczHWOaw3sGWXruJvu8RKmsF6FwAz/ZiQTtHv7/sz0cJYAQI4encwO
x/x06PeAYp3XbSP00Kb2G5Kb0L7d6M/coiIz7B85bXiSSimeIPvrxhD8iVSh
1Dz8aBn6lCIXsgFh+y72WaAjLlefvWfL+olOtWhCil1HMLo6eoCI/BF+GN91
VaJvG5qUIfKB5O1BuPIJ7eSnrGMTYGHmTAXFKMXgKNHmCzVB5I4TXa7TNXMP
79uxgnToTxj49fbbbb6dJFew884gFPHSq9kNEzvk88vhq9Jo0AJ6RwdBEjb9
nr/WXiQ4yvaCWN9IaidlicA/dq8X6ktxihsL8H2HRn6KiTlj0LYgAOYAEmZ6
MIDBqZP52L7KL0yCP6ex5K99uFGGiROS/Up7H1aNiGb/+mwOib0yYM+y9vwR
WC4ScJkJ06ejtDeF+MDTJfX5hVzjzEDx12/7wSQnV5YkabJNZmYCYavldIen
b9CX6jeB9uCJvTZIF23LIAVLCsrQ0nJQbF4eBBr/h+N1YiMyuwOzroeag1kU
xAkwtpFTUZNC+iP9Z7/fz6d/8o2Yo0MHbMxt5VijJGLTMXNBkFFXIIvOi/cs
mBjtBA1TCDjhMb4RW1Z+yVfveCVkIhrH5qQ8GTqEHp/3StrUvwe0dXEQXnzI
mp6MUCErslcdOnB6Cn+L/DXGLWdYokhHhYqNZ+l6Ywdc0FWeFeKvMRiFIyno
xib4gwBavBWoMMIc9BQXP7N8MCMHmQE5SAXHOLBMZ/0aXUWgzZG5uwL0Tklf
HZvBrfSBJdor7noEQGgb6p1CJ6HR9fawMYMUYDds7SO63DLBumUjoukK0gAB
cTNqdAVAp8V4khUVq5wlE5TFBlqmlMVwBMQctxZiLHT6G4CoeCzC8trOg/dY
jEKnUWequT6vA62qhja2W4zH/6nJoTscy03XZvoxNoklvkQZxnvkfRyTGykA
1ihr+Cr1sWDSrcsVccW16jmtj/ETdRaq7lQm/5uD4Piu7QZcmhT8qn3YSQpY
OuN8fQKQBfmt9vuHbq5ddSYRrVXQHcY+SfPR1heGaoTYt4PiDBiFBCl/DuHd
mu+Jykb9kNfVH7XpBBSuSnfgAP48xiGd2438IitGDetQz6MGXR9yHfCcyxE3
mhBTcl3qnDuBJJ/M6sNOrzM3qf7XVHrlPkuhGENXFbaGwfoWtmubOC/4aSNT
o6AzTSA/hPmP2b3ycBC7qjHQ7/t0dwKHmUQ8sTglz5Ektua25YEUg6iW5qPj
Xw0xQ5l/CBurI5N5fVlsxqP4FCBJvJSWJEMw/Ehe1s9Li+XDm3zJM9f/6I6d
NYkLJOmVFpY6KtKeFxX+jWMYO50Skrw0IeOXP/56A7zD1WSW6cXZM6fFQLYB
QfPv+0z+YDKHpWflP+A/DpH1cb4jE2DvPu8OaQHgZ1isJd/VWH2mVh19l2rw
fOz15aTHm2PR0ABHRtzaj5ivlVZWEljncbtgJPxthij/xEk55aT7w3ZEnAX3
tG6YvJ6SECey0iqneBvP2P2fvgXaKxaQKbbvFcBt7VVWhnGGerzV+DO+Cj1F
dnZDA8NTXhdQBfDw8DRLHRwiMA5RZy2bWa9fqEgyZG436ul7PLMEun83xjP7
fYiqlV+TxnYv8Gxy+8Ri98ultQu2lzG1O+0duH6KAQAextC+ndH9OHCf3s8o
12yzFhPlT2BoFiTC0lSCfM/y/ibHLdPM8k5bHitqhzvilhadHVFjPcSymSiQ
R6n/YX4zwJrXLHbHnAhXQr0tzH8mRz5eD92LHYySDa2yMmItZMZYydaUUL4M
1JrSlgq7PsNF4ipQpvtNE4VhP5DeArrwaZxwnldapEDqwmY9u1IMjavbnE6M
ClafTq2uqwa/GANWCQbslhkovMBvVcZAd8+I/WHMYXZFmxvvm/jKiqLRHTKI
Ql+qAsVF7oc7OON2DMLz+JP8OWTNTdRQUzxgdQ5nXEXuei3+dmI722a86Vw4
Kie0lkUq7fUM8LIvUD+K3wAkDorNeCbTxuiBmPyYkoW2j6p7rY7mgo/sE/sC
CIZns50MVxJutJHANEcZ8NDi2g5jVhjYs+us5su9+RK1Rch7mpShXST3smsP
y3oc8fP6r7UnFh/EfHgR/WBAEQWCsv4wC2fDN7/TPyfv/gsiVclb5kVpKhuW
tT5gl4b/+0AAmRX+MVnZKKvdg4pdhbr/pjfdfzQ5HrDmMnKzTjuHh3scmymR
ltWHcw7bxr0qa9RW7fuiLXPyRHTMaH08ENWP5URqqUjKHlB5qsZvz+N0YrQA
a9MAuqCb4hic4T9O6l+K24UrjMvzO+ThnmmBi8slsBOsF+VRmnZBV+ZCLmY4
ydP7aAgFa6XhSi+0xb0d/tlebzki+dZuqaDSQNZTVgj7pnNmXRGTm8ofphTq
YYmA5FLtBjeZdtv5Du0j39F+yVXxOP6ADqMo7JvgRAgvRwTowklqR9jtleN/
WLN7jyCjnOscMfyi1QhxIKCSrmRHjNZEbMTAiydXW4TSvOiDEm1eY4ynFC42
4YiylkZWqT5JJ5Nbr/NKvpg47RC2So0h7DDmJqYhYSuRYQoyy34o0jHonuo7
zVVosDLF4GoQONB8x50hRTdlOtYUDXfL9+h1l8QnkXjVQ4ES8JSYwgD3xB2O
B3zdiY5xVx2xal1kOD28QzyqqiMMcmovWw/sl2H8PBBUECFJVHSAsyGPyKI5
4Iuh6o2I+WOmcocC7JnCjD+FSZ9KGVzsbx++ckdo/ptVInSwWueGcShliYfP
Du22+SZY24jedQHyYT8zuSSVoAFCPlXOEHRz7pOTwczijqsKPRrjLrBf5y1P
0IeYaI0wYUOgVVfqhgr+5TAEj0xcdirk+KS/sJXxaKK6CNHVbY8QUMWJQMKB
jo3Jv+fOIMqbMC7WFj8cFw+SWIKb16CIjHOxQ9sU97ICZKvpL8f4vWI6iFGG
Pe/IOeEkgJNClxgGk+1FGEZNbnA17tnI3TgG08Vivdf1uiE9XtQBkPTdh97B
AM7BRgJlYRxtfnHmzyJpcPd5P0LXCE9K3UkyjkrTRfNZozH38ol+klpW7Ii3
M/LYHDd14Cokca7USDZQmLbJ4afJW6af17dcDmWKXZhwJ78/ftmtmbhiEmn2
plLG5R2bbwb2yqGwjJ+b5O7cv8g78yxq79JFnicOdwbN2rxMhPrG4FhZNwFe
D9TuT/AiDuhMBlN/bj6kV6DH5PCanHUyW9Saj2XjiYA9ss0dOFrg97NaBVb2
6Pn+er79UEKX6M8kerKzse/fh0mezLZJJEqmRTMORLL4Fg6ERN+3R81GWCm7
W7qlT/jRGfMNPYuu7nNyTEzOPGwFSq5xS/LrzJRjtjzQqRYEJjz1UWwhYOur
iRRnT08SCgZuOi5rxFCLX4nioRnUT7WLgy4QFQ57zCAhof8e8P+voTMKKgWB
/tcyNzAruGT5BnFOKMnJCXF1Lg/xsH/ObB1gqGqXI9G1mx6GBBQ8FzFq0Gnk
DeAMTg3I1IfRpSAtCivmE+FO4JWuTvJdIVaLGVdW7AjRb0cNiD4/LA2T3Y6b
lza0+2Gqta+1SXuCkDEI4MwbT45kkNwXtfQUv3SCdTrapPwyeA/qKP34qv3H
HTZ1xTkPKrGwKoR73G4OBlNCFUqVS9qQbDIAVMWDCMDO5Uth/UT9exqn/gtX
XFx4O83DtbbEVuE6kjIX9bOZd1ffnuahrUzCjhqFOrzfNdLoScpLBZ2iVUwb
FIxA8c4kPmPy4ITdrElR/oZgWHuSAncawi32UBsCRYNsms5eUqhYEraEE9uo
DhrcvJSu2TqTqKy9/RoR9Txpwa4kBV/LhlVerLuiW3+YfAkojQ+fE+kGMCYQ
u69dUdb3c9a+BC335HlQfC8jh+ftRfXem5Ky53u+nI8hPVuFQJ7nI3f5IykV
r/8fpkSw7sdQyc3/40XgOP9yFutoCeL+S1wmTr97n7yTmjBK84SGOzJx9x5K
nypiHs6d8FBCoKLF1Cdo4Wdlvjy/gzWhfOrgKo6df+eV2mfxHPXOsHHSMCqk
/5C+64YtQA/pYYWr8Rq6V2T145vMN17cqaxQU/jCDYqFgM0mCPC3ROyulOF5
kbHtJPvkDLmP1d85wqdyNkV9pvbes8Z77hgtCX6D/Tfmt6iQWxkh3C7VXUQp
OhiiQJzvuDzvWBF9Ycblfa/Qb2T/oucE7a0nC0gY/t8IFPmS/g2inVUMDiFn
8Fvhv4fBnAg02ZonPXCb/tkXBILVTYbeocpgGYiOkC9bMY3uX+uT47uiGfDb
1gxOxGN4bCR3JKFYTEvI8LACGWvrbIVM5ZpCsteFRWQpgh2Q9hePuNykAPRb
B49dLCLuf1m9DZROach3KL4lmYE6P3Jc07icSR4GYStAmyYA7TdYLjnW7Sej
sWOul+9LkXTgVF0X3Vx1Oy5hE5q7u61ydMWgJ7uwQKBBTlPrxCkAXWsFbItH
J0bGkpuyd7UxQeudQT8pwJwWK9jVXUsKmCBpG0ZGGzEpbKuWqZMa7AYZgkIJ
A8Ezb+prcHPwaw0N3lQp3wnfA/S6A3b7qSGaXTEr8bEHJoiCHeQOwSO2SBtm
Qa3sfkBf2dEx5Diieo+fSIYMT9PjgY9UOHrP4Gq34UrOxKiJhlGqW/go6oO+
9Pj5e8F+t3jArrRdpvHQPBK8R6XW51Ygub0HCzVyefr/m3RN8oNJioF7oGJO
7F5FCTta8UIA8xs3JCrp9hf50Nk758hrkrtA9oxOhgsa560Pv4/7cN3kPELC
L3XaLCZswZxULRpxUY//6BAuz4NjxekYJYxfHrBw5nI/wxlq5jr2GaAZ8rBm
p9gFLRnAAPzNwI4XLq7vNgQIqe6GB3UQHJDcQ8qU6Q0+dqQlt31J9Is+myNb
/xyh4g3jj/8nmhHzHDDBDkoEyD06jOGF9jbSipeo8wlYJQElSz5iQYakms8W
/ydkJ6JiGDQ0bqK12sSDubhYd8OHEIy9Yf/2ed8zybVR8Y9sie7FpMBIiLzG
S0L6loX5B0+TyDsXyHSGNVVp+VcThzTd0ZMuBPWZU2odZdRyywdaQdNLdS8Q
vEe3hxZCiXntFnHRB+GWdyisJK+N+aEydJy2YlEqMKvQ8kvE7NsAldm8HfBe
5QvrqtvdAo2MiZ6vvZH2t1mgf8hFY2H8iwJPV44ZNoTIn41KI0j+bE41TwG1
BAbQwFWaUAqv4goxbZy4fSa2B7OYuRJFX4T02gy7Jw73dfiL8BeCItnToM/G
nvGgcoV7AwQSLXIhGzKeg7RXRoekPWGXYibOcsABfwtuV4Y2FRWj1EbM/53B
LdpDdJFLgbLMiqIj6FD18ObylDcUzRyBlxWZoHzMFU80DgqdLy2e85FxjRkg
aaGz0U1Ow2W4ptN+wT4CJLH12RMZsJRDqx47Vuf9WqGm4NalF4PRxtTeDSxS
tsO64QQzuscuPG8ndet0+97Mvrwxwik0ZYQ+uxqW4Xu3VuzRofgUzpzM+rTT
qGG2O7O0HKrIMDIyfHTeF1/ikh0+rTMSRZXBCMaZohprizeKcqOVDca7PsVx
/VczJhGGMQKLsdjo7mOTxgT3cULX/fyrc4ESlw0iWJr9OmPRQyNt5zbTJSI5
1jKMgm2BS1IuxkuKR+ZQZ/jfOqXFlE0G7pVXni2X2RFs53RvdsaaERIW8qNa
kxdwSa+1GZyY8ALeOB9zUca3TDJqPtmYm59bpOYW8GKzZktONd0XhJjjUZ59
atWO8IWxNFIHptkfmHzZ8SW7XQeOa/JzyibCmrgQdCzasEcZRNNUA2e4Xrpr
uMO265BjFG3cojy9q5/uH8cjnk2O7Uv5m0rAU9iWxkbu9aEjJEaIOuZgUQvu
maE9Vt9Q7cA/CD+wuoswD2fDtTS14BvIDPtnIT/PmXsQ4WiolJIvTKrgsb2h
4qFtF+srCnVUHgtIpiWnPEFo0fnH2Ky6DwPLRBL1tsIrM/ls4rR9wn8iDFcl
fqvCmBKkHSfC2DknhMJf9hwXV6VdbW1M3Gjp/yuXagOrOkdLjM1lkhd7789w
wSQE6PkW3o7506pitspjQZM2QTzBGt3C5Kph1IoD5dKAAPsUnXHQtTeHohSw
62dBNa0N106C/RV3j1LF5rRWKUarPjeq6qcFBCS36XUtVAswk48IKRMu1oxR
WdL3MiZlnX5Lq21sled882cuiDJftncCqrhN2LHoKViK9chGLd2DA/KTB5Jz
/kqonIsMz+HpNZIdlai14DpUECf162w8w7ubbZryioMAyvKW8ZMvbCalL8yS
RmebvXym4EjqoF4XPk7hKS3BFW2/S5rHgwBObO82MKnxEL2gszJ+c7BX4cOi
8+adRkOSki7MKKOAz7GJ1uXx7bPgwNgigOUOQHTiArPJQQdfR+ryVRcFsLo6
JYoNe7d2stb1WKtA7R0RxK3QqLahhLZppYlFrpz85qTXAgmMiX7ISty3+Hy1
8rpp0vO2eM59o8IP7E1DyivsKPJWkvbDnwZYXQ9JgxaZqgOwed/cspQFOHZA
ZM1jUX/dOm4Jl1zhsS0dyIpLVH9WdOuTa18jCZM9Jq2bHLvr+VqJx5PHXjP5
6ALqwuZ/lCNdtho0iSihMMHLwPCzSx2yLgYUIhTRimA1E/2G1Q+LmYErWpBv
B2l/JZlGE9Q4XuSm7X9ma5BEQX+BwlKa0S2A4acMGjhckJLbRjo8Y5eRwidd
JLBG3Avvkpew/KMI8ipXjTE4EF53cw9p3v2o/T1Llkf1vXWDswb7nGe94J/1
8Q+C1MZKZMGqWaR1HXaVmK/cX1fxPzg9bjjlsSTQtFwt3+8McuFvKk6ojgqF
jIeypzi+WNV4zcSYYGh9m5TQ2BDm/Svvs8oKYyXyCHBaKD+JUJyE8hL/hTGZ
grQCYqT0Rlj4+r10kqrCp41fJqSxoSz6zw2udsT6dlxdWeECiyZtwZlYj4DE
Vjw0AApLe6b1SOOud3rL6USiy2YdirezM76XzIMqFqdUhrUwf/iObJbjccXP
M/EX+Pf35UF/MSzBKuMoqG7FVx1v/pphfd8SkWUQPtvhf4feNNc8axf9o04A
o0n7gScZIU7/TmLdhYwPvG8CDo0zzHgS5EmNky3OOhHg/fIYcU3NVovAQtBM
BVnU0ERrcKUET0/HqHEEEJfY+mr20ZjctLsXCIlFCBM6m35TdZ3mqzH1+q1+
Cu5uznAFaWHDs9qU7UxpYFLGp3HTUHM0U37ZF5IBaeh7nZtgqyzb1r4bbbJT
+g1LmZsZJA0chQ3bz4oHF2vpPoO1aipQ4K87HILbSHk+nihQTLnWqfJtaXRj
Vt24QhQY4S9pMhCI8RXdI/Up3j+1xRI1E1aObbzTwr6EQNleKNimetEsfXuP
RLLpbDk43biAfDJ1zVzhQlaTb6DHegThSw0D8wCleGmYKmc6a3dvSkkCXdsH
ztaQuGkYnU7XjUzunOBi7TnqvY0POkJCt5BUcSus2kgh5L18n45jiinYNx1D
1WsqtW/p28GUQaJDlVo9ntf71Eq8QnUTt0Ed7cTOhGfGwMxmIrOhY6gTM/qn
dAEru11rTMSfF5VpduYf3+g6GNkm4Fz2yOw0tcBtETquAlQjNHgFUa0Aft1c
LVb5nGxnOCT+kWG81lcI8buYUHJnmkf3WAN6umPtb6FE83HilWX5RePPxPaS
qaCXvAwIVNmLvUbnGXZBJIdNkzhP4MJoCkCD3/C11ODvX6sTYAwbbRTOcmrp
9XLTLOQC0SjTq66zKA7sf0C9LHKIeStkc0/LzXmVpQ8ar284TiI9kCRQVQY8
Fafzx1ZMEirG38as9n1/r8t5iCIljwdXPxWwqD3chfJNzr7pmsyUWYaG2b96
JrzhDB27zXT0+BPiAcl9oXtfv0TLBbK4h+qNAZszgDfhP8I4ev25tLYCm+BH
uWbKNkny93ZaE9ScFuMN0eNh1ZEL/HEFG6JdbubzTm42i0iiCfu7eDfneb1i
LOkVxoxcbWjS2eFFGaLPF1Q4B2RiB/U6Gho6PQxepHbA1vHHYO9SB6Z7WW33
+Qr15+SFEK9uDEv4SN5mX7AGsuQzbrFUEgXtQnX6i6x30Xr+MUSwgB0Lvnvl
IAfG2iEEuRORe7YfvCBHwGcveiFhCPVHRdRwyoblAOeKEWUXvRzd7fzp5OAW
bC5dsAGwLrXTa9jeoWYqNae+22Hh7HhKB4WZhkmAfTtqEg/OJ/xVm51IeQu8
2fRG1YlXu0kM3+mnDrYIxUBXCmpXE7KkCri3VxrklGJ5SowW03tE4PKjp3xL
FxZ88q7fLsiugxDSeUYETBiHX4wvUVlZB37LIIBUogyW+5aFRE/DQwTMuGbb
qJpeF5Qull+wzr1ndyFlBxb+jK2bp0Ph/BQHIlOlg09IFXweSgVX2NSghZ7B
Tkdb86WT9viNH9Q62CReiZwCpjFeadD2X4vr3i5Fpl+9uxf1zw+h9hAS5XN6
DtY93QheFkOYP6NksMHPPPIpoB5VOjvDQg6IPs4wc9LQmcpPKkGnXo2vbakD
yncqRpbNk97mdfgwLlMkFUlHe3ca5Mq1Y1HNykTpMpSupdDAmZFc3TatOKoN
rvoFjUvj48PynVkanxDRaBVwt3jqsSutaydzYueQtIXhMDB7/VzrkqCRikvR
zco78OAgm2aK9rcE3RX79CaoeDHRgwrhgg8gZPXVcyewbeqlxKvs/0yNvotb
JN913AI1gjhS4/SnrwZ08BjClTiGnbT9idxrjPDLCSvwaxaKCB6+qmHNxnqp
mP0Sh5i1umWXifaSNqm6aEY4PJ0BrQ1X6Kz8R5SP+aeouq1AWnsgl1ssQL3K
z51o3tEUS0WNAqY9o8tUaldNCxM3myYYS0Ds+EFfN1Sy6gVal01nGLIWkb3g
LfQdmbsdkxGy2rRIMwMCqbibQw+3ObxGoCqQhBiHUUTB1zX+/M7Y2gRUvrxH
8QyTw8AfwLVvcwZN8enXlBtYT3i/dK3m6IXIg7qPQIIgsNvslCnaeJFTuKsa
yYhixXV0n8y3VYv2phJ5v8Iib3QuOS5sbMDX9Up5xF39FBqLbbeOjNrlEijN
RUEsEhRzelVpRjn/Mwl+DMKbV/7oPdvxN+Drd36Hy4Qk2HHGiLH8Id201krl
PmIA9brapWgS3r0XAH1JDPFXzIhqFLy4oSbqD2c/TwwFLeZyUYEnpi4CyTHh
cGX/j85qIwb2AgfR0iUVHjncQgvX3+wU7yffPlGSLAM4kTKkycjzCR8yG3nS
vFK03WQ4vlnckkcbXJZJ8QGcTItDXyJbmH5e3zf81lnwgEhCDeoEkUXMAi/U
bailzXEna3fDbnQcDv6NXYJNOtiR9n5NZImZUgAQw3AMchwdP9S5nZjQLqiz
+ASAT7z9aB6lpFEXjoGR7S/+qwz6X6BBgMMuVZdWcWay+AMuQKDHiFqKOiGG
7nrWoZ9SpM6PR9NI1vEGjWyM9zq3fGSkcEvBDOL6sdi5OGkW5VyVJHZJ2s5X
ZRMxZC7TxksNc9mN9o7vQQIVrrWSutImSxWwcvQzlt8lHCw/pee4REZfHHPR
YqK0LIDzOFOOBwYj67WvvvtyzIEly86tl/HPgjTIzys2+WYn9CKaFbI/kpOd
WOnJG7/hFW5jBTbWpSTVl9Vsv2mSB8wrzFjDFxkIfcEcE2kqFfkX20LCqkY2
RTQ54gab+Fb6IneUVbPk271YrEtkYAUW3WNJfj9KTMzjWwqXu7Isrf3FD9nr
Kr1FzkvnnjLVtxHDW19JWOLVZ+4MwUqbebMmyD7t6oASqPxezZVHB94mG3bM
nLvQESXS5APYjMQskQ0UNgdT+XH25iwxtt83bWBirRPzc8vSnmQK9MVElaWE
aEenoYJEZ6xMYv95kCgSgIkv3jvCsPjoDFRKRsPePu2T1YoUCeMfPUc3R24h
KnBy6c8aLqFdeGHAWIbbl8rJgDQYC7ONlpQj7c32RnQbpUfKs7xkr2tRU9HF
BPuKSHKcZ5to+C+K9rNWznQ0OG7lRig6xhd98gYNVVZqLyPkDiWV6gfY3rcT
oaCrvwxHFtjiaVnvVJFsm78W7p/UTcYlSJL7GA5tyZ5AtBHhYGpB6vNIQXfX
DcGd8NCixJz94xsxn8KrIMMjbLoPb48XWaJupF7BeCE+9oxNb4oXTXHYr3V6
2lPW6UbhYK5YvIqxRqU8vEZPhC9Z9ZzXCXtyaP2rGUs4hxNDiiyn4XuksYQN
1NB0m8Gf1rlcut1P2g02VkOIWj7YDnFp35bucwsxFr3W3cAl9vOFX1eI3eWd
MwNbRo+l9c3XZRQUbNBqOffoPMK+9cbxOn5fnIAoIatNOsnOTK6mf/wNqGt6
oCaIVDsMj3hzjUDH3Nt83Hw/RVeEM46jPZrcTMZdtbpuLeDKjVxomQC0V7qp
vAocDmQvszwJk8EBVuI3loyLmgA8eLzHhNQZbF3l+itySy51gQFK2zlyjcTj
71G+tsTuMpfP51aauoI2O3ATBbNRKfV1LdRG7iOs+TyDTyJtvmHZ+jP7NHg+
Tepj5/R0qgRv2IySPJG4FPKWk/C9j0D+gPcfz2vHOt98tLXKrDUkHIK1sPcA
HrWzq77orrRLqfGn8dIanZxQI1gSV1rH/GYSQJ7TscQh0pDo5wMtCgdrrN5Z
9CMyEpvdrwkeLxnThcjiz6APlIN/arp6CG1jzwbJWZekMdPRpiYRJmURC2Dw
Ag7b6Ee51wQ0V3mzoq/fn+UZykcVqkwoUF3NksR8rx8GgVjOEr094TMuv53A
DhRWhKzMEuyXR3HtUWGQqdupHWtkTOOiU1VLCuH6e9omx9Zv3AQ/g+MuLK8u
9r30Grnzc3WVmN2ER9D+RlEz09yvZX3sl9Q5u8OU69qzIPjoJyjF7I4CyaNW
3kRSd7itb+QBgsh1TAM8eqIFA3I5W+ahT83Q7UK4nDZna0yaxCWY8YgpLDYL
9RgDYMJRswhCgGo4rz1EVJn2bx1p7VDMWDTqxx59OHXOxDda7tp2xlkD70qr
/tM4GhOA/dZSFD73OlgmW3R/yMe538hAhJXpIOhFBYOAu67MU1/+cd1TMipp
vpRVcnrtDGFBcIrHa8fF5xCx/uqIuNzsdwESlk3dVlTRnrcEczCiyDKWQfCf
xnvMyX5sDsE9u4+I302wMUYiw/uL25qf79cAq73LoQUcP2LSbEvWrORbxnnC
Qt7XQ2/1I81l4YvdTLX6alzXSKxs5pIMPnzB7tWxssxq5WsDhloE9L0H4rgX
HmeMOz04/UF88S026TcKLKqYPLbISOnHp7MRUs4aNumdwSmTBdbE0Fb3CCpH
p2dPwlCu8p+2P3JwUFCYnljUTFjn9Hb3/vuTNcx43oOwpICGiCluEn6y6eWR
ZTpDmc9pswW0BYaWG83394mub1GURTPtAQI0Y8mVfMML1vP4XOKJXzUIJjVs
unQ3bnOp40N1pmIcmdNkZePh0gTj8CbHEqpZfRyBxe2BDndw2iPs57CbSPb2
/KZ5uO45gb+9viyIOdm42v2s4Re3Fsb+SoiISc9k4+6ZwEB9gjFkFfzgOTp/
XFf8Ch+o/Vf9HwH1KClzk0pMjryDHXnV+fIKjqcCxl/QCf98z4S8wzJFQYwn
UPMB91/9UfagT8zABGmIObI0StlH72uU9qLfmkhDsEGQNr0p3G/8SG1PeZLP
4yVWpnQ2rDThvjT/8bl97VPl5G8F8hi9JbOuO33Jyj+CFEi4pu5RgQmrjOlJ
UF6w+JNIoKgW217Ciotm0SQuAj/RG1E+J6J/l37rQaV+A+p5VqdnU+PwJoSr
yGDd49BW5R3JE3KGQSCjxGG+eOVo/DegNoMGaxpkSvs36xogITpnw4ouKMjr
oFj4dRdVC008MaBUJq35uCtX+hfMeVV5+LFVQ8pEl5cA9vq0dZ8Jb1N0OSEn
UMBwrwwkeILscwb4ebZahhg7RISefLlbdHMpCWLUparNOlwZpOjT4RqfA6Fp
zscOOwBxxHsx7uPMYzXQrd5X8hNvw1AK6Z1RRUQ936yz4Cd5zrP7hAfrK4eN
DMahsxiq4KguOxcnRPqJST2zahMKq+/cfhdnVbjOmlEmeCniMcvUdYVDKtrE
yxjZQkD6gAeNeMVDJvdwTsbop6T+al9ODKk4EpSVzUzqmbPyLJkCvqdzVPxo
vwUNL+wfQpmQNEiXeC5JNYNqYOqIbrYTmAYTCXQXt+znHzzd0JYmxhn7CVdy
Z5DDGHK+pbO24UcB65f+wiwulenqLYoGSALXmvpuWYvTpXRsWVc3ufiFDhp4
gu3IAw0kpGZSMxWG0f+U11V7PFv3RDNAIVIYmnwmKdIThGgQV6m+o3jYAPWh
RD5yOHV/K1RyBxjKROIVaM70v/lp0DdW3S9InWIcVU8f4eZYL5Wb1OsHmKRd
wK2o7NefaY5XnL5UjFH6s7ZzVyjnQspTOMeBwxBZwJFGXkohaqTLEuZlulgT
gLqS3FwMwrcIskvYL8IIB0KJDXMoymxQWjhDuU2EBKAlK5sqsUL9NEKRykp2
Xb/o5wZVbuYi/4rifXgHQkGpzpqNkDsCPVOcz/gDXTiZ+0zJQfTTYKlh6BmE
LODooHlY1p47y6CWLzAy2B4K8XI6TFtPrS2Bn2pETz3PHELt8R/KDTH00iit
MErfgaQkVocwjjsARk5miP1kQxaCdb6HJPemuJpg1rnABe/MheNlC/wGU7q7
EwHYUMRZDF0BDG1sNTtA5nm9hpRT8F+XkitnfA4lrecrsmDQsI9Qj6FThySq
3x3nLRcrSldjcpEXalnCpHYAz2E9BZkRaScqD7ffwLFAlbnE609fAbcMm1mH
uk9MNktMUKIcOG4SYSu1ATgJ0DkphsGS7m/2zEi/WEESq9Sdr0/+dQXkLEDV
qkUekOv/Gmvb9V2OLWr44FjB7tv/cH69JywJVGgrTpBKbgh0sL0jtyNr8D4w
LHZN83pdmwyqipF4DYeoScKnIgHm+R4Qq3KnQnHlR3jQ1d23DZoMEEbYIpDi
ja2iObG6YhIG9ro4Jdra5YuxLo4aScNVHCIhKMhCMjqrigsqNVi1mZv8bhrs
GmcD77D+qt/vKlfpxk5ulk1vJ+/pi7dL/3iussU04FitPl93YQi6XAeEVbxA
FOPDCsXG2bi3jOySzuO4yUOQC2HiirOAHKha9m98ZvQRAle9ydjuycSOVXFZ
DPeLAyBJEle6pE9L7oSkhWtQmxwHY5ihjb8gWSSxCnsYQdsC0Sz+7rKfIIe6
AQsc8a3tPChzzQixIVZLnfZ68LuIGl8cvWqr1pO0UK+JXj7wCm6WCXXdNA15
NG27GNeVwXhNxkfVoYiWfAC+aZE53Lv09sDe5vOeLMe+pbdWopGqlmUOEmWZ
FpnnQxn/Km5jaBF2VP2e2UZomDyh6WXuOMY7147gVzx8RtufJggSj98FWvhg
gg8eWOF5ftQXSYvRFU0n3nR+ZjyDoK8VKeMp6Tl3xiPZse/h1h4evmp8ZHrn
KOl1xtmsbq3+8rKkMxK3ap6y9Z+xo+EpQTtg/oXQvWs6veJ0230SSy0QB1pP
Jwv5G57BkM9vObdXfBdnhm1ftSqzDsUnjNnfYI5dz5MCeJz7an4Hx5dqhT1w
27DCPD17jXa83BOTCVAOjUYZhmT1v5kK8wvs4ZMip1gIcTLKFRjY4oXMB/NA
JHTPyE3X19+m7jo38NbKAIKSWVvAKl1Cjm7ROu7FDqaY5JyD1pAYesAPCJNl
QTqq8xeBDd5dNCw6ueE7V7+MSNzkwagbF3x+B21nxjGuQW1wSbVchmYjXgpS
DqRSDVtwiXV0w+pFfYZ8HEHGt9cAo+0T1Mo49RGTYZ9ecIa/1of4ZvLcU7Fx
6dK2ZjgdHzEHk3B0L4YsMVayZ8n8gQZkrawBQQCVTgv9VH8MgoQVVBZW8Fb/
JXTeWULQC2Xq7k2UiKN4nDwMx/AQDQA+q/CFHYUGwASKx0EbE4jBiCauFSw1
PJ4Q8fx5b5OQAaabUrtaxbQtYqzREV1m7kdg1q6PUfvIfgBsGJvLK4qICp7D
vLUoMjUia8yGipYUlbZIb8RrrbAh7AxmUAlYppqmqlS7hx6CPEnjwehowBrB
Cfh4b1u1v46ljXzb/RUpwRHTH7QXhHdMC72OnFfy4kEHMcgpBbnWvMA3dPCs
MAj3UjRURBa433hNdOeVVA4fG7h7VQPVziimknj7VxDtWJjdqb85TsOjdQDn
JLKTEPq0HpWYnsGWjCiW1w0+GE9RWS3ht2UQ343TJuMU4yZIqBcHqIGUSf3N
xsRESsbgROldb5MA8UruNtnUkokdjOxTA75YQBF7+8XzCgyP9Ra1lg/0fuxR
NMVopT5mzka1On/89dBn3GIGWduGfE/ODp26edqBHRJ6X4HaJ6smeKW2GgFG
pneA+IbG69zTdjsChtEHitkTxqhlLTYX7WzM9fo+sFb38M3A/OaVLBPez3ad
QZicUCWwCyIsmeFIlHnNjMeFk/vTBK6pgO8TgfKMXheT4SNBDoZupJ+Mez8c
OnyVDZkaaVTrOy6/fiiFIBlaDPs1uzvWVgDzk+SrYtio7GjhSwLZl/5oH3bX
n/k5WRE3bWd/+TuAkPRT7sHSX6O5jSVvn5EAi3OHL2VHYLLE6r0ODPVjjn0l
fwlXfn3Ba6JDCAS2disQbwYC+kFkBSxxyssy8lzd5fzezFZ9zOj1QulidbSu
uhwPb/CPvK+Zq4wnK6cW7nuhX/OLf7SbAcGne7ULh/R1QPmrOu/iwsClJ2Gw
vlZGHgrp6sdI35LHAn7Z+ofd6vSqZ1Wur3A8thPgh4ptpZn/i8Kk0OcosD/l
IMUBloFZbox2l7ZcuNB+vLX2BvtCJa09Ei7bRRbkjLVGjYH2ql5KPxutM+p8
cIM9C85/RZigAa0w9+zUJxtrM0rMwlvMUauCYAhY1pun5VW3qkf+PuafSMMw
gnFPZnp0fS5XQjqUlkSIovqXzcbwfP5sF18qrqGgntKCS5JwQWSYZlNqsmjO
fKPZzSchV9l5MusZ5pt6WUo5r79SSG8I04zgj6GH5gZj9zDr1ScqWZN4JAex
cvcslnAOUrfT4rZCj4tgsuV6gYfib3YOnDibdA37gXfi8/r1CILXob53J9s6
rL2mux5OA5lEJE0sg9GsE0/y+Qvtv4pRXn7jDltTez6BCqbKhBup47CmwqzL
vdVEAw7mpPriE8nvyIBghVXQ9aZm34LE5S3oIGKaNW7msmGxjg9YL2usIcpu
d/6ctYm7XE+k2Ni4ikFMXyw3N2R+miv1tzWx8hWj+aBRc73cAKJJE+Ugh1TU
Eg3tGeifnom3Xvx+Zze8Tt+bHhgJ7jRvdWoiYYtW7A6/hq+UuOKzTlD8aCDO
G+tH6MrQI5SiN94erqW+CRmt62u/uixv3i+/OUyzawOZg0Dwy8p0R7pHyIWF
cNIYkpEAKUqrRBaGsmbcTW+8/Ph1WUAaI98NZ56BB4/0H7AEnzyUoxDK0u79
h0C3a+54SdYTkNJdDzVUkxoW2Tqlv+KEZMDvrKvoyGqpmlXKfz+EGLDcIn3X
YWH6ZCRhX3dDUZHB73J0R8kAOQcRpgg8/BTF/gKjGIUzLGwlHPuQHa4zqt01
sO81GAeHv2QR2OVck1YGXOOP7SZI1U+h86CvWLSVTIKgceGXTCAf+EZvElxF
g8nWREYElaUlmLc1Rbybi0W8mvVMdLWdbwu1eA/mFmFMShUXary4ln7Q7cdQ
YWBboamoHMVZXgSOuJ/EzKZyaUdWGDOILKQ6NRBIZhR7wayOB6o82cXQwgmF
Bqu5/6EdGTkanuK26B3cFthmQ7tcvz0KY9QIs9wdSR8a5dpUXYOODvHyzcbf
TkkCowZMzqU26VcGJJVzx2neXvbom5fLTo0J7ip38mVnPF0QJvJcg9ogLK8T
ugEfJKiXKqXk+yXQMTyYpKY/FC8vi5AeLOa5rFWM0XwQERQUFrkZHix4yyz3
i7V0SgM4Sz6tvStQc4Oq4zv6ZARnet/teFaIhD7ZqluinAam4KQvJKECb6kD
SqOzVistHXjWFlsXBGaB6leb/kTcWYyPlqIkQWGgu95qmKFHaMk5L25qlYKt
jGDxhmO/4i954tHV2BPlXPoUpOwus/Xt1ql7QIANEb9hHrzD3b9Lv97QxPvQ
6xvIoHp2uZxQlZFqD1n8Ubb5Ce3bbkzSQEQs9Ps6ozrT4glEu39AtxPyx3GG
S8Tu2BovihiaZWcuYBqXck0eUvapn8UuSxLcM3SWHU4fQAzr2z+B8F3mHd9V
8EysrzoWgO3SAVvgYDvuff3m9lc/gpUnppFWKslec1zkTVkH3Ddkhvhj6CuO
O89DJeq3ml4kH3Wtk/MHMdIUWqwGLqZIgECa3FD0a+0ARfqaI+JigQCnkKrz
5qU7yIU6Yzn+Mqk/MI5eddfbHCEqr6k54GyI0LqM7DQwW4oJQ01+hWwQw/z0
54sXD/ZP7SUa9QlmPkRxX8jmkAYiWfgVru4VhWdYjPLxO0dysZsmD2RQcpHE
Tw0E+Ba8C7ifjDYKC9xkafjaavv8x3Ab0JIo11xNRKntA34vRgNUY6jKgLIw
wMdwNF6HTUOwcfmotxwqrEnVp3rlK5wkp+BF7jzm4Tg5FniX7Dzln6Ze7wgs
+ERSdbjwIotHvAwJTxWBHnxBpM9zwswIlA9eMRNHTtoznnvG5LTHj23qoPTG
+8D3VDtaW1gz+kVTHivTM9MyzdyL4RDGHEPkeS89tA/NMkpSlAN+ZVkkhgqA
gZMn9dC36qUOIQb34iUFh6qxLWxPZF/7z4k6v2IlLKJHsSpTPT7pV3iCRO+t
YSK2WTG+1v5pWzrjmBnUKkQ3mMfFjaJTBay31mUzYauaFwapDEgTN0tdVfNM
RkTF6nC7FTG5bTwxGny3yi3bh77yABJjJYm9UYmqYrJR2/wIfOCc3Vkf35K5
ZbpFiwcaEyEBoGxOIhJfn0fyIboOveCwchmVZ6XLxO8hdl4kUEIYOphBTWBK
eJdN7XS+DfGjWFIUFDXdrHXnEkov6o9PWVtAI0pRUTbC8Qoyo4FnhR8XWCIg
zSkw1jt6Vguet2N87t19j/ib2b7csjuidacbNyKZIMDbvqsipbzmHr7Ls9Eh
yL/Yre8nlwmXdirigCRhcrv5rWruNyBY1P++LNKdKRnZz8YXpDsmGTzVVC33
ezqKdku6+pPwaAw8kvwpMe4G/+bgY8hD/KQNZA3eOlrCAFD/AUkPtXmC4Um0
j+DE/xg34nKHn7zh9e3RXP+fRgoRlKyT0ALrbTA+/fzb9jtMgtVa3AE0XVnO
d6A1f/sgxhEONtxOkuvYBTnMNbXZIVRP4QZibi9V3gClPvBTTfJvwYRSpC4+
4JEG3fGx3b9otp/QQaKxoxq+JN87KIwQ8iE37NEYOLmt2G8o2u+NV+EcLDcx
XK0wnp2TVcxtr6oKTfdpPhttoPDZnM2DYloYPC1DMYZCTs1nnMd/PPVAWbiF
vD8Cw6K9En4FVzwyfoXDeJo9eLHge+T1v74KBqilbvzUwNTttFjpl8xY+E7h
XRa/JxBnh1dEzdq/W3/mbP55wNO2uLX+2mZUUbuP3Ltp5RdhGx4YZl0dUBf8
cZQhY+cWtLsiP/tGWO75CqWs63PQ5la0zPXCSLoRsfzwwE+ZsMZs8zNiIUdr
XY0c+94npgD/10TyJ9kAG/1uFcgANCAsES3TqWyw9VRCpRB+00ujpS5s1TFP
skNDTKTfJ9t+fG2XYBOcxyfC7a0kcMYOtM9vpsRev9DNKXATfQrrEJNCnuul
hOH58eQ9qVUUiOvuyiPE6cWB5v6KyQL9ScrLbcgBIX+V8hLVFc4CQS+qyrbp
oj7mDY2PZr4uPw0Y0Ac6GqQW/DALwaAaQVqtA5hfMuP8p+yLio5rpsp1d4P/
7JZO9Jzyj2HXt+yfPS8+rzxucmjJKZh+P45FVu2x2HU2FdGgmY+CqG4O26X9
eE4Z3kglmxq1mg6TL0nxFifykFn5ExXbw8INyO/g+Z6walca3jQtfcOQVuKU
zjJbdc5lH1CL8atUi73t8Fmjpnr4D1ue5yQWVbM5l45K7TlWQFWzGMKbiXsd
jtnRn7ZKSqHvl4JEBKPaebdB5btNCtKsk7XNcWbOiJNHxMKD6+EV76tZ/El8
V47b1fIEEywWNGXxqPYjyVTwZ558aNGsg6E8LmqxRALg8EhWf1qBQeoOqD59
iK1D05KSD+4PDaD5TahAeCrO6Ilsf8XWmjuJaMSIKPLKbxM1Poe8blarFG3i
9xnHhQSFsm3vEv5IpcSDSdYmd2V3hsAnvycCqgaRLNoAuFxEoZh6NyeCCdA5
zKmDqQtQXIJ+9NyD3px7pHrm67MGSq+sqVd1cjYl9E2T5cUTEqhqw1BG275k
jZndkY7DJICq9nRYjdijA8iCd0QppadgVlRqm6XDNrJgfGGz65BnlH9edD5z
dpMJfDI/fc+okIQhM0G+dj00WyHE9RYUZNvoFqeFlvukIjiSbtWkLDZAozfy
6Q6T51+zHz5mM+TGdPUj8BGtTL0RFUaELaYj0UOhwNO5AktpjNhbDli3fpk6
SEQUKJfXAICFndRJ0KnmQKWrqiLM1snRDfuyhIhzv0ArBLFVVVw9OIEuFXkt
JmC0ERLLCE9ezPMNVjzQQKKNn7vSi8m0b+ksTWhr+7oBpX5rpVWL15emOnsg
xikQva1rl39Zi0ARhdWtASs10v28y1Fc9QXuIzHMWd56f8LUujZAnZqKQXos
tfukht50wK7jA5njLTvIDNm97QrwPs4KndoC2d7odiSMXU0dvqRYaT5LCx/l
coTGGI0WmZzBr5DVfHXlysJcaNMkiHZJFKQhCzCXwnoiTgNZvCfLpjAIHPW/
M++tl/nxzBRFuZIhMpL5i5zcfx5v2wBkh6yTnW3ut7zfinW3uYVZ8jrGGY6k
yyyzb6nJxPDIiQIogjtk0DBXRIN4IqrBMOrWIyw1x1390fvNHGrMj+hzVlXM
8YjUgTpGXncHZdVuyT9IplGgN5cWfPKjm/p/P4wJNPFTwaKVTkhDTWAmcRWJ
zNUu0jcJ0cQQo2IZhVsgKdzEvOEVp8hO+J3cARkr1v0Twqs5V1E5bUgV/NnK
FaiX/O/hZA+PcjO5WK6YQlJ21wZh+Na8IHyPpQ1TZsHBqjnkYRy78xMaGeXH
L96EE7DGQX6GUCEsfeE5uI0Pl+dGUS+1JQY9stF/Quwmgmkz3m3ymMJUGchX
KCO0/1151jaYcGVrydzI8C3N4rRA30kjVP51PADRE3eVj60MZteJLwXUb0I/
Fjo56NdltbMPs1FVZHHEKa8oEzzBlha2pqZMU3NNfNVvkJSkS1i883I8nGhC
f47CUp622iPkjxbhnWNK6QDLJOzt8onhv4NGSaEIv4ruYBYZcTXNN0/MDrlR
le0kzQmpvJ1wObZXPqJQoMKGNHm3xqYSMkhfOba+10bzvO7DAF4YM0TJylMk
EnQFLnWTImip9apX8rgkTLjk8X03udgG1LRvzzxNikSgmvUPxDdS1Zx3HkAq
60vvOm/9Afh4UK4i9MHYziLtWZAnIzQ3ZsUQbwEO16cpq20ptvUwtyMbC0cv
m/SwPm0Kyc4uuZi1wk3+YIUFfp/4pJbEYcZU9ldb0jUqBicb7IzESFTc3uH/
xq07xMkBM9sMHfYJyRG5XdCF0Zp1O/MWuXWUAMSa8T4ANryYrycuf406Hx4J
RgGgEQ5NVIF8HxOQxz7qzoJJLiCU3mG0X5rfU8UZyvM5ns427AAI/FOXvpt/
DHePrXDNEDIBeXH1lgywM285LleeXznlkG1RBQXB0FahDeDCLRRIA0xhW4AE
VHdZsU0W1VA5ulyDhbec/h+w2dKOMLaGP9Weu++gxSpQOoBSClM+HUvluSHq
vqmZmhrmaHH1bBL8pKu1pcEpnny4iP5vlYo/N1Yw5i5M5oNKDAi7uyIpS8pg
rxizERNAIAy2wt1BCRTD31pqr7Twe7mShTRJunPDONMe43olYRRjSI/AM8pB
4GspXz1oIDQ4rk3JSbkKvxRyJLHKJwUE/WJjEAqYx5ZISM7pIxxQvTBPFXZn
DTUeX8OeorE4A2af+PwklvDF7SSkJCh7Hz0o8HGkqIYiG0zPgpAMqcP5sZCt
aw7LdnItJaJGrfBjV6u2ewgMTfh8mQWwF23CQnMuXnWi1e2NiOhtw9aygR/L
W/hnewlvnistoColQ2FObR0FhUFfazykEc4NJL3yYhu12ckp5/84pSkS6ri7
2JIs/RC4ASBbP7aZ9ICjsasYZ/eaFhsw5gEfrzvBND0a+iFqVFZoOajz/QgE
EQyHYJekCZkkNrHqKH2oduU5bYrRv9rZVe1TXYKj3R3P9MCy3Cw5X5RHwCbR
UFctbiHzsWc74r7vomA+gWgttVLycd01difP2+4tRNwVlDYgk7rcwVXJ7EzA
9M//qpBD1/fE9he3/36s1G3XXRQEXELH1SgQO2UNmz1oV29i9Gq76qkAiL0Z
d/fR3riuFWV/XCSodWveVld/V0TH2lpflpbkxWhT8wMcprIpgWIE1vm+xi+U
tCxAK84iDGzYRZNLr8D0yJM42wsaH1yt+qXN041VGfNLNa6IcWYUqPPhC3hD
RqiaY2EXds0yHq0nGZhDNlvY36FbLrl5jG6ELz48imBlnpKsHSkmVekJx7ef
XlGftbtkogLvku/nSw+1+5MPvAQbD2kuQNaKe6CCeaHN2I3p/Ugth+PCH3Ho
2RL3TfDF6/dQ1w39S+x4r9rybO7uororyIWww1QunCJMBddOmaAtmVxWtWHQ
3hTDg4Gd8+kkwUBpAsgLynCo5+Vi64+bgPQ3eXrIZ74Hcw2s0Xnmzx/3oq6F
KeTqohjOu69L67HNVa2Fp2rhoscgR+ckoctLiNgZf3fl+abOvz/6NC8FcQ2k
UXLOCNrCDW5EQJgN7TgurpRzWUWLgnLaqn2SCrNNljkoa0d+hYgUbauB+nci
Bzfy0IQr4DvOQLBlT1nJhlLQpFVBy4u6sIAOMh15qPlH+QgU2cOxWCIeTcBI
m5pmTfTvKqVjD5DCMoPVrPAuR43HgXJAzoWD+OQbQkUj84IlQ/eqMeKnSO8I
HgwP3SrXQCZ6LW6jc0k7gJz5uxFmpl8D9lcY4SDlv37kZTQy4ah3gT3ioUX2
8ZLUYRgKDfl2mwngyeHpx+jRwITE6XLbKaXf0B4lWC2UKotPzXIz15RSFzUY
mCiZWUVXYq0dSXFQEF4oGwq88nrNKCoGFzt2Vi/J+/erekaaf8iKDtX7donF
aOzMzYYccOaxpo8ELJbBvqfHEWgyMo2uxTxe8wUmM2D2dsbrXPyUdF4EK00y
Nlodw87BOy/FTKqE0QXZo9xxMVxqJAejXkOenqlytOXBIAf6RmmA8S/8qCLx
DX/mQc2CABsmpeXWCY6z5XwABI9NEBtQhs4A5vXyl259M9wuUtOv6lzXRtVQ
/s2ve23Ec++hZ8h3NNTGJI0+b8PDvzcXJxBGbWUpfibJ3pq3iedNwyI/zuZo
VEq0DCEvsAtzCL0/DtLagp6xEvJL9lyVUA9EauYJar5Fm5QiFp5T0pPWT6gZ
87EXylcAFem+oLi8+aPt4XB8Atv9BSxUXhpUikqNAISAYZ52dP87P9W7FgH5
qIQC6DGWNfDD70MabfpugPbpCqN+BoNSWCJOXI9rGPNMQ4pXxw3lUmtqXgk8
VTndKmEBNLsdLXqVFJSyVokeid14yYgegjelRdrnfbEYHCvXYA2DFrOIVkMP
Irnz8ml6qW8bSK3ZH/n33LhMcageEd1c8YHowVJocCWo0OYJzXKtYfdqvTu0
D1kc7xttRDqvPuEcWD3xQZtGNWh/wLSRD54/rQl427yts6zd37lYIB5TBWWd
JiGU0f0kv6GoG8B6uH1BYg5xdQg8u1gBIns5FpmkRJymbMf4QS+S6vsOHdN3
Yc8/p1CxV6BqqRymdXstyHTo6BL4uMDVKgmyFue0eZ6WS5GK+GZ88oPElclR
kVF1cayvTfDrMFxi0NpqXgcEZlGJhH6VjiAaqXHzXtlutZa7I9lGbx7Ec7I4
J4Gwr4QY6J82RdTsKbEv3jORDiHQmt76qPQyZ+KfDiPkbZ+lMloIgfYSs8+9
FrYUFeV+VZee9JeQ2QL2lgfuuLgsVjphEUdMNVGn8plIX2H7DWvmnuQtYvcH
PI2gh5ReLdONire5kMev1ln5n4stnBx1t31LcDZDT9cf3UZFxKztx4Hw19E7
1e+LDfGwd4CnPKVVsKbwyOXs3wWuJAEd1TeETwDXMHGTsUYL/GfGWDeOaOtT
sHWlZzF7IGsH8f6adWJbIsXhzhRVPK1Wo1WEojSFIGohTovhb+FFyIC/Gk9Q
9tY5G4pgGRnZYWT7ekiNG4Xd0OVow/jQHWXpRugxBRx3to65mNjZgSjDFsW5
S2MFPoq7y7q4h+ss/Ur8DlAJVexJ3L4/lTKOy372j1RNgMSeAOoDmrYamuKk
8y1gHphnKZ4n+65MaHmGHq3SJeCAwZm6SdId5gNeHrUUOxX4hI1gxaTDjbie
vlntxctkyeRxsEBV5I5BXHlFCXj/xekINMvnQ5OEJzleWNcDN4fS7U4GxAJv
2gNr01Fu6cvWQa9SOBUVMGCg6f3F7KdoqJfWfN2bosusNMb5b+xZdiyYh53K
Uv9naZ5f8ySKxE5vtMDDRkE/XPZfr/adT5TEjGrRPgYxxz+4RZLKPoS8k3eS
EW2eqxspARp59z/TGiHqCLfhWvC+3q8iyIx1jpPu9McBJq69rL0L8Q74RuQa
mYKixaaZRsigvwqaSbVcU/kysgldyA8hmm7w1+8ftxGgBVeA7KcxxyhlDNg4
h0AMNY772Stazq2dN//PwVya4rUlZtWGXEq1MMiiWb6oggt94LxR9kwr3fAh
g0QJzKhEmkQsWUgiweucTjFzYt2R9ZFxEMyHJ/QVPylA+7HWTL3Fb+IK3BWI
jlcae7qzevjLtMvTBDf9OdyinTZbCcUWqaeMi6YawT6SzU//6nsv8+Eb8tJF
Qv+CPD6yoKJJ+HMTj68BQMB8LWr9vpKudeMK5AUhD/PHsbj2JV9Wy+1Nq233
V2dAMvv/KROPEwwKjLoXItrZJfvh0VUmV6L909w/y/qyFznqkCAbs/V/4n/1
jdvrIMkHmZbFn277D2rimSWemQLyikNUIWnvFq2CsuxmKNTTwjArziPacQQa
J0MJyH4TCHKmbF/FpqTDp1c5wjBYYn7tI/wfUsEnPiBfQu+LvGQSCOdkuAsm
QG3SaE7IsCvEdYlsGIhMGG+Vv1G5q6eG+TjO5BpYUHV9FQ2mFX5f1Uf9Hl90
O9SDrmITLfxY0LSoAziBVNvr3t2NcbA0vOGGzXLfTchV35TLwOgSZABmMIs4
BxzmtrMR431OYrdRPxPQAY1XP+dO0+Mv0gk+hAKh4T8469bvg96mU5Jm7G+6
xNfORxlMx/34Wu1Sa9hwWomWKZm6ndnXlMkePlwdO75+Q0o+87RFjeMYp10f
EDSXwhHAeqcD0zFT2DFrMBFj+MmEbW/FPmPH2c2Gj+jjTMaBK54FdNb/vAEY
aa6B1FatdmrDmHCV3NiebjKAEDeTEl/FuBH/CQoWj+uMFHwMvr7LLXZNToD0
uqEbEHcJYgCwiirBrrK5lD0Yi1ZgJNxqI7XwPdj8AxhNS76T2NhxPMD0ZWMC
jU/LJqiR25MzT0YqBp1cmceRei6ljNNbXeAzgl8+R9TwyDs3NX4IZxQuYniT
6h3iDMTYIV06f1w7eb+Ua1t0N4UR3/jM/3atuTEV38S7CkOsDkjyx1tUmsD/
dzQ+D52kVJnkaRl6bhOHUrLMlHYjUKo+zcTdnuhvUxbkqTK/34svX5NauN6A
l98DfU5+W3zUeDX6ZcqO76cQtdPkMLlq8Si4ZbavejwTzIcKIU7n2+pqCK2O
CyXLc0hUQqLTG7eGGdWyzLY89nnz4a2oaToQWd8sa9zZPPwolyOTk8PUe3sQ
2FiCKBDNBiyqeZUGAykR1hIPdugg9a7FQaBWDKnyxsBfLfAA6hDZVQujb5Rl
H4DoyBiF4nvzbasxpqddzAirfoSBPO0pcoEWK4RgUQ/t3uTJK9OuNHcQWDcT
H4kpcEtHluZEhuS8CiUh/WbzXoSB8gLy3Ez1d5ZpWT90jH52OjY4d6c4Cjk5
EKjgS7mThNs/bnxvLz+14Yg/JU+taJ+x0kWP/2PYyeKO8Z8Em/0T3xMn2uvi
x3mr1pWqjK7I+tEpTiqKdIyIHnhLtJq7KrPFMNCoW99AwTPqNHo0qIbi0MKI
gDO/1w4XY5pp/3NYNOJV3S45Mxx/cZ+FAEe05z9r8KAtAQDg4lHePA27NWQ7
RzyngS9pg7L9pEqFt+2jdOd9wuxg+ieDLsZpf2bbD3y9ZqnkN4veTqmaCHZk
7FKIZq/jOpkXWIA1hq2UYjXQ6pypLi2fQ6Gft+NHlw11DvI1Gg6dJijFf3U5
aC1QjfkUjZMOMF35pKlVnJNVu57Y9CV5ar3bdb8CIFCvla+dismOk2Mkd9PV
ufgFd9XKyFeRdoERNiO8umDS9y3vJFjtZ1Ui3JSIqguR91/Jun68F+6nu+kr
D3fTWF/z5jOYx0aMmk0i3Gbqa5D0Od0NXO4KM6WuewSoidEMYkJNnLqpVULO
MasvENGe+ynDO1aRBKk9Ll1zsclULqAPurdsNANLNLjV+nsU5Q/Nv+7XwVoe
Om89yX/2gcnFmR/b3zdKxVvrKtzNSJ1DC9rKG+aLUDjxhp3k3pMvke6fuaE4
oSUyHGMAEsCPHSb/ltk56H4ydFHo+nmDm2V1JeU25nASf2A9P+wUySIupgAO
c/LvgyJFQSR2654/+dCU9d/IXKIERK0SrPQMIbzxsPMrLi6dDkxcImhnM+no
K7gGiUUpV0BPec1aYtQlglpWZwK5/zRVEvdnuEwH/LK1gX9idlrrCqcN5t4f
1p5hdGI3L7KKMJ5qZZ1mZTPQJdF41v/Td7k1B0DOHPYPyaj4u59sF4bTVxzN
D7nDTvAE6XtCbkOajb6U5s+3yePlmzsKfZSKs50J2eyV6l+MLQpGuWiwR1vk
v6Qkp7uMy+p2bRMNNb9zHqA0dReWC+0KQik6SrJS6ZE7GwwSEOoLe+qhcS10
CkzuciZeGN5+XUDl7LTcIeKUxzkRRasp2jRVQFOTmmMo/6FNLBBzKbZUzfSC
VRV+AuCsTUH4qbQafYOoOOl4YYyRKbiqDC99KQwDBzJR3IFanQpJEvrnrB25
qvik8y+H/MuijfAvlEmXB0fQ87KJL6N8ugGR0hxxjTGT9jn4b4Pmn0FrIjxD
RRYN4sIUqb0WI55sMoH/zsnkOHZ8VH/NGskTQSPElNTQ0X46XVuQ6xkqaP+u
3nV/Va0TWL4rd3VTXlaKWzZcqnsJSNxd9959Wkc7pQsTV6TutD487G+z6jVK
4iSB8bYhme5FXDe0H9YakWqDzj1ysewKAOI3P5fkRzusEuCOr8jxRkpHm1rP
EvpELL5QbisRxMRzAlykEeWGU1SH0EdQylzFQEQdYenYWsr2hrSwlCLm9lG5
tAFRQQkBxXavUfiQfcX5F4YXdo9+sFv2XqF0GLs0L+zyU73qG+s+swMQ6hKn
MHZNYG1iBQSMj9M3FfosLbmtNx7T61uxtgeO2EY6/VbB4KD69Xpbpz9enmmH
kt0IxPMFhaFRhZp4YUCZLdnh/fCJx8CJJ7GFuHe/HYtxo1/0MIcwZgaOQgIO
Us1MH8SV+XGMm+dhKM8FcCwXrKFboounIeWvnNFQD6ksrYZvc7dZDmP2qC6M
SWugj+YnCKc9eHhoKdbfhUBQYPBBNIIWea9g7q1k5rkP6/5uATbNbIm62HT3
Kj8l3BT/M2Ok1nrBavMHbcWGe81lvZJwuKBEXN8EDPQBP2Kz8r6ynjr9FQu7
IpsmckSHGDC/F4lmblfdEf2vuG1abdqGJqDscqWh3UjWj/X0cTI24FdfBeEx
eMe8Hi2iMJmR/ievcUpuF6cU/MRJf+MnC1204zJoxi0iqlw56K+FTDZrY9e6
k9u6JdzpHZpdjU8q+/+dMHI2qkmsBMduuspcTzh2RST1PlOJUff/9lZxDays
3YRrF5mg5aPx/XxvUxAl7w+B7RqJ5eZsuWD+JvWIEFHEIw8mXEipsSIte2YP
ICGrzofgaSC2HIqyV13LUMkTdwEMiHYVWjK3lpCp/lwr8I9FFOhhJ1xhWGO5
9I8dRWdqYxrR6Sf/FfjnbRy0BgiK4EVaIOspJqL7VCevsMsaG+2pFfl4wGsm
C862N5v15fNbcAal/8hlHF7mICLb8ie5S6xzc4tM+OWv/XD1e81W0+UXf9Ot
0Aq76vDs+i2lIbFJgr/KqgxSF04tQY0P4qgB6UAMQW3vhVP+4i1uYEg2SwRQ
RkxHNXu/r/OMsItzBbEfYiDxyTN6O1Lrh50a7ZjStMWbf83O/effZyzeu0Hk
oc6C8ADW+JhHZkTjCkWvNVtgAzKOJ76MPuHGkvP0uyhihl5YiHjopMwkC8gg
miSrH4L61dsnYwJ8VvxT68VIj+6W4nUfEIdJL5yQ1Z0anLnfrHpR8R542/9F
r0R9f8jqcvV0vtK0MublmzARcVjvPholXaVO0NnBV3rsFyVzoh+uyc5OH8vt
aQkQY8Vt0WtCvsLpKiOk1q/Vip66P90I3EA6VjkKMTofjzMZL4Ufmq/9eTRs
0gFGF2GiCy2ew8Qy4F5XPg7KHLbSHUv9ohRmm1D//1kDE7ZbMAZcXxt6bDMR
nxDzydwTgjdsqpzJ8G8v5GNew4B14c1P6z1V9RRerX5IC2O5hXRGRVOF+xrR
7HotBiAEnOoG6buXFVu2PvPK4NNFJ1i8exgKAsW77He4trofoxkvr9NHZGsw
ZhOAU4bFbkk4wamsvZwpPYDTaxN1mpj5FfuBU/WoNvYa6ldWkublXcu4zG25
+QtJo6bq5Cd20fdlTJlQaW5BUaaj3ZcCYGxZgFFFnwBlysDKLleTmQNI7dkn
i+vpdYAX2WQvjqpiTFYC80kYoRD3X+Uw9Vnsafu9F/23YKDpn+a58R5LYERf
VxKYQprkaJRAaAIO+A53Q8w+Co5Lbb6A4k0k+8LzH2SgWrfrEchLtVyXtEIG
uynm549C9MsJvSBtNrckCRRdvjmfyNSjmTRRUcgx8bnU1QYx1Qm8qH3wHTwT
QZquRQz4v3i6EbF2Zfc2tSjn9ZB6LibNL/EJpAKeZh1RFeXCn/d1XSKOnX16
AERIPn45AC+UhTrmA3q/3NoLjd+phLtDI3m/xiqTmdUoX3ub327oNrAaCJyK
4zwNjSAS+XCWKjeMnhTUfH+088nZw+3TlrZ0JtIaDoPfHqQyiE3p+3k3ZZJs
tG8Z+cIAUm7DwX1TiUoX3IlieGViYMJg00k2/OumQ8wXXw0mFFvmFl9p2IgI
vlPIjU+sLYHykm8tnQ2AWsXzz9kcvtrDgM5MeTFqJ3AA8nOGYE/LASK/6iaF
lswxLHnfPhApZQEDOAX7F9aCZ/l3Taue/E5cRrALIHkS9ft2F/NNPq7UckMw
oTmfDo4wKJ2mQc8VkoINmAK6W8xjmwEfVozbZwCnqsW6TrmCKV+cRGNp0o9B
kI6JUwfSKFChDwKw2r0+662Q+fUU2+kgtLNtxkEux7+/byOlS8qZegoMDwDx
iZTDLGIGCKoZ/0C2gYOHuDPi0A4LBek/J3VN6Y41WrwKMAPWcJfGj4PjKIBX
WZ72cKM3PYgI5VNupWAJdK+0C+fRENNOkPI/n4DB7q5dOJ87BaKpS2QV097K
3cG/DNTI42M757lQfJXSB1Baa7TGUSueqwSroB6cIbXYNd3O+ToRBTXLygUd
Wc/Ngrme0rng/b5hjixDkDr6XQGpln3kJ/zJ3fLUN3Zd88BxSaOsYK0Djk/I
dSD5AaOp1w7Az2r0gItsWLLH7bbsbWJkvO1TdImj+lQTNBIelpr78z8JOLOG
TAmSUFYwWX9Y18W8WONTH2ls1bsegMzeMnGyDgs1makj+V+k8wjNtbc1UtkB
4brFSYtI94FaJ+uLa+AnldixcWMYjzEwZZheymuVRW1mmgzZnM5qp/ekRLgc
cunLlMzT+cC2cx0a9TkBmVthMFniXigwnXudtmEnDocQQE7BxSugCgWC8Aw3
8Y8Of0n17gYvL6pNuS9UJUW/rZJjBUwftKGrqC1zgdgNaL7uaJqxvy9dGu5e
uAHAiYmxfd94BgpPwWhkvW353zhoca34pBGokG9/S7O6Uk6xbusrPKvrDE+p
Sf01Fh/oM0MqCrD1hDlUoXrEpbXNApVoZ23pX7GJiiEmqAquD8DmeKXAR4Om
7Hf0niZhO7qXwjplRJD6lLS4jqrG/n65Gt79QyEehIorWfrNAJPs8rs1rMSN
SrrE6NsQyam6iHeED2DI6bqP3TyGOreCUKAnq/zXq+PtIpZDLCWJigfwXhCH
g7V9ET+ObE0pnsP3h6Omqm0YJYu314tGiiHodAEFfptTkH7LC21DYSSi5y3K
1FqtZA+6AnpIN/cFj5FbPN8wwRqqAQjp1jBH9HTkPks60CbS5KP7KkPWCaxZ
J5WVDfw6qDbDpPDgFjuC1gU77XAD99Z06XGa+pckjyDdUNv/kyXPO/GXRl3e
Ci7xk3MRdk/f82mZGpIjOCNHZYRlLWnnFFZdbGM80pfGXCjyn+0wiaf+39Xa
2ayIj0+WJ4WAuDE4eISTjDkvTQ/DT94gzzfKjbwMNNi5ojbu+Cqsfu3p0V5N
Ii0ADVPMjRIRYlkXSKVnm7UTege9dMoPg055KIqkMk1ob4JXHpzNcGH5bZNy
sm6aOV3KdFmRSQvthG5L9YNJginYHdZ0hA8R4VaBltA6OMy0P8FgELSFbflc
tVEj9y40/wGaWt933RmEt3y4/nG1ucLPx4uruIl1oiQymD7ZBbJNTmXgC9PW
O7HyjIVKrOUGMehGI9dFu0WLDgu7kfeHsMiqAM6SAtfhvbLo1rBpJuPcmHvR
61PEgW48Z/5ahlDcPrOX2UOA7lFBjeCpLJCWpvUksaWjm2EFgpOZi3whI3YZ
y+Vt924xTu0NwW5JXP7CULbW7ytNQ5YH3UqgZU/JZl1MacMWSyHXaUy+d7uV
EUHnJvE2rO2wJjYTvblAhJgQF6racqaANtKiQ2nu055QlaaUndn4bXhVEw09
Rp+02eI2hp3WWywMZhiYHI4lAszNs1vkqLrxhRPY1sLCOsHTkU+taiboAzhI
w2ikfjNkuLip4nHTfmrdJyt27BVCslXp7YTpvxw76125kw8PYLIaTLIvodBW
FU9vGycd+4zskATLXtCebz4TqNJj5uSA+HSQ9vnOZKg/VfzVULuU3JNqnRQ9
2RXekPiKzgSoXzxs8ibQ/gJ9/dNjxFLOmhR9u5v9TotfqpP268fIn9N8FL2q
KfXQzRSqZo4qffOOmrGM8ZARKI2zWoikLnTSz8QCrnaOWVUtce4Qi4kFxY6l
g97DlIvl89I3KAz661qZnors8+n5nMfZxlgSnk+z7HlTW7Up3bhL0k6sZOzx
xbmqAGUBkaxjQ3YFbTuiwNdD/K/KXemgTbmvSWU0rgqSTKDSFKsUS8xY4136
JAcKiG/pQoAvzsgYJFRlk5pj21Y0M1FGx0JqCwUSlpwDMczkZXCzCLXk621M
zZ8ovmqM2vaiO7oCsyCovk+9YAH2Y2bpyIRBJFaO2JrIe0mNEACd4Xw9HgxY
+7Zu7iFJWGho4KIyybKExUn3J3Sr5xQMiVchkaZpgKgT2POTqOR2+hHuobma
4mnNkGzHBllekoybr5zPRvhObhqiu4YBc+/2SoIn9Cow5+YG+WixVyUJTDfG
k5qc6q8iiFlt6dw6wgmDvSFxB8o7i8irMJLge/ZOz/JTnFCW4QTZGyGm4fjl
2uqONCIKgYwvD/gwav7VaxMMXYZLMUA6+D4TGo4Ps5waYjW4Nmmrjg/scJYg
oJl7QoL2t8++MK8W9G54d3gED6AtR59QJLr5xQQbtOpp/VPeLDOFlVrDHOsc
rMsfJxRLuByA7+/BwtH+/iaIRmTX9O/c5NObyuJwmHEclDhy217AxoJbpvRW
Dyw9fQ7cxu7nlJL8NCVFz8nb0co+ESHI4ti2WTac7WgLIt0/qaGsyo1Ct5s3
wqQSB5PhNRsLJw/98LRYhNOC9Ur4YqmwLaTWI6RmMGuP8XKpjFsrGbB2baHH
NTDwcHzkzRXx5csDwnZo1wonltyvrv537G49hpv5Ft28YlgVg8X3zvFU4IL5
IRrJ6VRa3xugZ1H5XXCH1GIeZlixWUQYwtKb2jajwd1CoZXb2qziRd2yRvj3
tLoroDbkxMfV9xdovEOfvslstRJP3An3LRXO2Vx6liHDHzoUFAjwNmIYdbj4
mOmGBbNjPXmXwJuU5aclDcUK6xv8Ap4IutNCIaZQUTKQeWft9HSF+HPqpQmo
AYkgkyxhlYc3fzWjUaleTY7UqUltLK18YbwOOYDBVvo0FyVGc7OwGXcQzPsN
rrWI78Wj9E7jgTLy+8MQoXya6Tx6talQFHsTQ3jzfQkfkYh/OMlojZWIBokf
/CICCQeS49YIFC3/4Mt2UWsoV7GqBt72i//KdQskQdIa48px+311334Y3MXK
mfw4el/RLWmDBANQNOMOfzJ648Pqvd/248RxUFp5b07nJAO6t8ZZ5QpVxRmh
GI3twPVvWkY74s1L8UiszAVvxuPmmoxeVmwmbHvbnfTM8T1dd9cmF4Wkj/aH
WZdeUY9ua3E/mPKKYpvLOzqGNfMY4D8FwK8/omXvOBaErIaNGYnQd5aTW2Jv
9IU2YKJQm2AyBxaQDdAtxsWIovW1CWlpPPgM6w42M+aZ9a0epxMy8dUn7qtk
RJXRb1RBiu+5jlvAbVNB35fBGrxXKtHEc8574WBtmK+BY6oydI1lDKMH38DI
0udhjzZf9w0JqE7mnkrzocLe6Xw1anfdbnLcOWoKXNzUwpiMd6/mQXdVCUfC
SeD1OYkKsj5pe0ri4WCmIVr8jJZFkLkNEikWpEBayDLkBPMNKST+wPQ05opW
+rEueFmqq12VB+h9BGG211v9YKyFUoLTI0bhd9c/cuW+d77ktyJUPaNYBIpo
dNtNv6Xsv26IHeaLBZobh3TAtejeZo81zJql3gl4OKU4d5eQzwUG8SQef6go
P7P1mljTJDKOfJcelN/XH+qeWq1SWd8GeWOp9H+kEZGf0LSRYTzFjaipLT/z
+447+ZkKAXBp/jd9hFpop28PsNPalTIP6ZeGuvLZHd6CDyqpR1Mz1/O6/uKe
CckYeVLL+WQ2uOc1BAsdvFxcj8QLiKxXGp1ld2PkOwRCT8sXKJdWdaQkPmw2
2fB8hka3iKhm60/zcC8Q+CJ26aSoZK/OPwFTKXV2rCkeC0XBmPo/TM+qoHud
04BnNh2/qT2lI9xCujE5aWtTirrZqCpxboOLCmBdBiRatfpLle720liBxKxK
KNNrsXv8yJoT4BW95GHnswwZqZXAAQCTiNr37bdKyzGDZaJUzUb6IzssYMV5
VDprZBrkwLLUWAohz98H190HTf6yp/yhrSQXyvuAIVyZzrnuSCSz2/QVJww3
sDXCpEbQ6jaUvFZHFDefk9RbIUFaasOv4cUzmMBL3fH7+Gp9l7aRCXbt1Owt
Xhm+gR5ofaERAyApbon2NcHFNrNutHBELuzxGaqwQ9//vW3CJSOMpHn2YwyW
/AXfOlDbNhUPhQK4nx+uOHhwc2rvdQtUToylpEF5hoBl0tM7UbSzk7nwGjWX
s52BMm1FrcjzvNHezI5xOjB4VhsI31mdGWWeGlhGD3PJlASXpo56eg0qMM1H
3ct0uYpymSx6n+cEG9ax2P3ClguDO5k0wJat03I96M2oMn4hOeDLlVDDkawy
jvQ2gun034tWhK9PWq3AgcuH+YWDtm95qttsDSoROJ22yBjEweNv6zrhQCXZ
CLilkvtIV8D6+dw/mXmmxwSS2dkzatvlS1EoNmIv+/vQOH83rK2bm0gCVV0E
a1gnN6EeLbcjD2/HvkkM244Oc1FoxgJEPTiasDUeeHreOwroVULhFJIhiPq1
N2TT8ACuGQ7dIr1kybNu/gr0ZCtdfiRrWTDwDGJjDHpneI9Gp97wxzV8Op3d
bFDeU4rgtJZdPUXMnPluUy1tB99vybpL0tkx3CtfhVy6Nu+noZWK5hUNMHoG
hMwfANE5dBSssArNqRqlk2bdl4YpcYZGabqApzxZKXlc7FCLqSxtwX85CMDv
4THF0UpKrt8mzqyekQogo2c4fdoDb9n49D+LmXxMBCo81uSMjSqKY9zsl2Ds
1Wqyftrxx6sV/Fusg0vz5cHsfRDBNBAa6kml/0HYCzuWCqtSLkC29MdZNay8
O49chrOlKKyj8mreRrKHvH1CvV2VJgkIm6kllb/kg/xM3pqxqGE5I0arVa0B
lMWTb0gR6rI4TrLDzsdYQUngXg218dtJIhQvEJj7Nvlky+ojN8FnUnSo30SQ
QEayrj8j6Bx1yn2l1OAgbySp0s0Elr9w8ozMwTZEL1OkwseMAUscSpRYGjf0
RwfU4ENz6e1BmMiBLiJ+qWI7nO3skrg18jTzBmBu8xi1Ye9iYqJ04vkOgCEn
c8awffL83paCf97ssOuacJSLqgbjiqyDTdD13XwcKVySn1HC090nS1Zmj0Xk
q+Aa9BBHYhc9PVc+DCGpaS454SlubitVVUNOUPPWCXPDmCVRFCm4adOjyhwL
jJG/yn2VLLmnKWGCw2PLXJVcvturnRhbwHul8hUXPRzrM3O2N6v5YwMnqNCP
ktl8ScG4xDYCurUKQZ64+3LdAbXvgUoK9Zs9hdwisiKnIVMDMj9gb31UKZyK
484khn6xlJ0uCANstCPQI1Z38lxghJ+P/NGh3+JTX1nmT6NJ4BioOBWxRAjv
OJ4fMljzIamWETUa2GEQ2/2EXSoAX+6MtfO21N9QoffXLMUJxWsMGKPVYJ9j
+HFwdMO9GAAMsMOdv325TjPgaJmmsgQ2/TG7dFV6HktWmsioe2F58sjV1P6K
iJqbXKEASfZ8iMOr+haPi4Bq6HWoIZThmUjnnC4ddwLWel9RpwO2DRP6ZcJp
eFwzIISh0NLorXdyOlCHJm2GPYMl6GRAMzM8ECd0cO9D7u49G9x158wsjDDG
gw076qS/hE1cGxIBJuxIv7Hxd3XPpNCWIslg8rymKJK+S9DgfHtuzRHEBf97
DRyseZC0xcQWd/UhQwxeg3cG2t6pRz/WrDQT8rEPogqf4ww0tGt+fj0pwZ11
VWTKkcc8oCOHi25hMnpPYK56Nwv7mJ4EZQSl4t8fPtnZrUObYojhEIxxAVcr
woR0SxwsA/AtgGImxxvpHC8hmTDsDmC/oalSmfQk2gVtut/B5nLW5AB39ZLc
hR/7cu0L7z/2v6tqGKmfeHuR+EwEWYhQu/pZ/MflWkw7SE3mHCfKnshh/D8n
iMQVvEdPeBCd11WfCdUpm7u9OWIk5W6Gba3luK5izmhA8OcGc1JOd9z6iGGI
X08Zo0B/UGX597byV15ibimSWJ87eBlMJ19QoL3ZKr9LnC7JHFaD9vH81ZP6
lk4xDvjBeTal/X94I9jP+UQ6bV0KbksWZvzDXh+BZSrzvhFjRw/Fpb4V2veQ
Oyq90iHKpGULSr8Ba2EfFGTI7Jbt8Ub/qA4JKnt+ZygY/CvZKO1ZTu317wzl
ovXvubIV53PcJFd+zVYmFvOrW38WScTPzjI00ZMXWWje1D/BpUkQGsHq+IMG
R+nb5OZPjSdt11v4HjK3Hs28S8AMVer5Jn47hGJax5NBMznRcnoaJGIABNGI
QRFCsn/x1HmddzuLKIH7uTVVq4qFU9swxFfu3x2d8+Ibsq+n5/lvuW5qpu5w
GMXHMQ6dcYp34cofoCZGIVotUBhm6SiujBe8RZKUpt+T4/5NZ+c9Vw4VBcfB
W8WmH176SMaQ5DZPT/CjHRfxcHU7gPGFKyA9co9zKRmyS1R58OX3IW0Tu6lj
2Vu7VRjJ2oBNSAl7HvJc0o8/49/KVVvhpp/IrD7z/8S4mU6yx5/c5MtPPet/
ZBEWREqHRHgCkw6ZiAVhQkVKrd/uPreCQ95SxshLFXpoESpMKHWZ+LhnoLII
LFFAMzRGCCHkq/UA/4C0HL4kqDAJ9AQfQV825/WQ6KsLHlCDTSgs4tPNNgg+
bZCqnvArly/vLPwepYxqW2RS0z+6cxIDkxD/yfeQzAQ/BcrYDvdhfsP8OE2t
0oN3k2Kml/XxLY41laK1NjI3lUbPM3pH3D8ex8U5M38TzXLeBt+SJr+WDvv3
ijKK+nAgndwEeL1gbnTMISue1ebqH2h+Dc7UfMGDskNWR0Rgo56ovw53Mb9/
2E+JkIFUA7XKS+dqJPv8aRPEy8/tCTj2eHEAOmzpd7kLYSCHKBWvQXI9Ixje
IPzVt60f7UPG3u4VaEHT1ofBsFc9WPLbCKN2zR2pjxRzBN33sNiW4FFhenNO
jK/eTsZ9lbCe82xi10UTMkcxgipEfxpkYrk7Dh//QoY7pDcFKGPz5tTRd2gX
zJE5FUXx6VzrxXKHWXUtE1Ezar6QyCYAjWIjfHAbsXV1E0qPQ0sQNPJgoS8w
3RZX5EyFh5QL2Xqj5LB3HSiqHnBfT+3g/+bpKp+uoKyaw3Q+Y5KVCQ0R3Wb9
fN0Op7dj2oLHTFDZymbP2cGDKFJtbU63B2gRUbhlib2m+vLdOGmbntV6cCaE
zbYYnV52eL9yjXUxgKvyuf6fXRBV2HIOuTt0VWwsHtsd2Ww9xo3k/kuWzOYj
6K2MxNgWJzhXIh0MrncE7yHzd4cqRXw7YYo8WJtlgL8Qn1+oubRVQfDVYflt
b1VOeOG4xFNYK56yw0S8vlcJUR1/C39afUlS/kw1kBTDu4aQMkoWomJI/Ult
8xH211ir6IfotJEmCutKsmBGdPST7N01VYvsQEYdr912VQHwHArfuTUOt8n1
+ImCwX7KoXqIJ79RVWdmgI8a4Bq7r5KXjoyy0m7O7/q30Q+m0hnIvZWUChpl
T5QgiTWT6iLgUpr7u43qdTN/8lZuXhsDtX51kfEzX44z4QacnTuB1LFCyORD
XPtCBibyTTXN1PhEwtTQ2d2viArYKEV5+LDoohmH6XAu5vmG9RNqtzYGYOGZ
4xmWSFzgtel2jsmtQbpWKRtDH5PSwrPNA+J9RHf6QgoweLV1cJq8VcrUeDY2
4cYNtkliuI1tGIMYkAffTQfYQaiT8nT/2Kv9VwKjE3icGjETm4XtFOUNdRAd
ieZ/79heYiogEiIbFeQ81KW149LCDO4BMNkjIKhDELA3EneD4Fqu56SNT0TE
IOtNydcoXip6bFnUkWzfBUEJG7tJ8F1yzpuBzYS2KBVcWt/SxgwhBZcmtmgG
MuW8yLx6cwPlf07mW7dZTpc4Oym3V2UgMldlE2dVAHIi2lvJ1wvI62BzKOt2
lBaIvBG6VFwodnPEpOk8zYPC3LfH2S404ufObIMAt2sCe7vCCel5omk6Io8q
521cexMuwCzyY/B7bNEG0OjoTSpUxGVKBOT+IB/lmeykkqokioBlMuTLW3xi
Al0S02kkmRhuVa3tYvBpB79shdSzRvuKyJzq31f3cIeWvCY95PiJubkzq+aH
Nav0lJttgIMHnzLTrELr31MH5oJKypJk1hXERWgzJj5C3rndp9AZHJoT8PS0
YhQ0ILI7Jg9Vak2kV1Fxff/ZN6NMssMhssLMgPdr1ZRmeLpyCljcsG6lBm7Q
QE4sGYDa+EXGtbOFRUz4WUAjD1ZK5gJfrBhXD4KeJcUE0O+9fiDnM4WTla51
SiXmWFVxfS3p3MmI6RB4fx0Lwwon9KtUczBxppRvuidGw9+CpLaxg70HrAlj
lumjGOX+TuS3TuM+i0+3ky3kVaKsHj9RYTbQZSgeJ5C7Br6DbkF+xOeSNcS8
VJlam8Rl1tRr/PjgpPUlRBt2JtllddwAapJE79DMlT0dscB1/o6sx8at9gqq
av1dzOIvsWjdWnIUrWhS73GOejXLSWcUqfyobh3iTE5gmsZYy919mXK1Oqhr
i5g6A5FTzqy8KvnQVP0+8WfXiWVtHrsu3oMH34BUASqbjzqAJdXDfLtN9RgO
tiMh+2QIZlJPgsmTAn4L1oopD75mSPsTxeIiGeib5uaqaJ6cRV7m0e/5iVMg
iHBahQcBtUTxG/f3QXjiQ4hPsTAg16wWEPaIh2FsWibmJRTDN0moavuLnIPT
NC6fT8oXUI/my7fHskbtCGVFkrEbVN083mYCI4GKHkFVbR0WH+2gl9KmxdH/
jZLrJLzJ5XLIAu8zi6GpkEau+LZyWhzoXe+leQ5Cat995M9eD599JW90JnfI
Bf1evsgmTnNBv2SbqOXfDtaCQB/3bnjk1uLj3MKDOAiPHDGd2fTIyuy9Bn7A
BOZdbhHcn7Hz0esXx3IlXtFWoJKdDB8X99C8eJ6ha3tpJ+jk1UInhcbnsxNx
7UxFXvIgkZ1Qpl/oNsu8q1Zg4We+LJndomfWtKW2i0fQS/zgEymykodaQWZg
dLHUUUGrX80/5kNsfnRZUxtxY+NASLj4w1Bwgfz9IwwKGlM8Gm1/jK9Jb51j
xnG5UqUWVw+JQ4twvFKbwk3PNbs8G/u18b3TCoCsEn4ZEShBSRWcsTVXRUZR
7Heof1l4n24db0cr3tlRW4CAh+nB7me7+st3EcRJwnf6shvCAhvmZyRoezNr
wtoeybAt5V5l4gl7RKan77wjlSQW+6UCfk6EjpPff3bfKvVBr0bjuy34mVV0
C2fh7IPvvINFQDcyQQ77nUCvX+9hix10I1csKhujyrMXfsfPegKjXMZLX8IP
nk0cbCCYImVtYiAWWh5KUsFuSGHLrsRC/olePorlXL9UoqFNIfxrJpC43PKC
iCt872LmneQVeSzGYQYUESOMh6qS0tff6FMlzs4HVQBtl6/xwtsV0exwu00Z
I0UrfWyUByNr/vFyGYF7Plhpr4qa4fC32nE/FEzfb5pWFxvCjsMzYa5z8coB
GVWxUi4S9eZ1/yvJGVmCW9bEeVFoGWDDe1ZgiG1EzJrrx+3n5piPZ3PlBBJe
pmXxQSpYnCezQtbWSVRg8IF4UqPmzBtK75adg95Rzfl+UHF1REn83Zb0sE1T
fXiwuhOHtRGuh10ucl/QiKcWFmoXQg9AukF9OqDOQyWn81f0FpRCyTaOd+lJ
CayR5+wQSErMJs6/L3LxKQSirmLQ3ZHR26ZR2XosLOOTcdy1Gvc+nZzC2Iw/
RYvy9NSvoL6rywNrJ/iqswPEE7jGWM9g8yFjDQQgY7tyTDEL+UQVijJ5+kr0
o1ai5Y3TQp+ilzxbIQjghw5kzIOdBbZ/gxvTWO2piJHumUoVFYP4Cv6dy5ml
VXutUYswjqJd/TWrD77ri38HdrZWRyGOf0QSMT6K+dRKRPUAVkoBk/0i2RcX
/xxzUK5jtPwnlJOHucZUtHqYfluOi5kGd3ipvWxZiEHdnK4UJavizAelyJZK
tbC3ohZ17wk2UR2ZpGas3uRP4hHZ5RkYqOcIBw90veMBxrr6C4Oad9jqCR/d
hTlLpaGOcoyBx/6Iu1tOTbh3YFiLgMtFfL1+REum6rZdLB3WbSyFeEMaM6x4
+rA052hQOnSrfB10A3IKQcNmqigB5tFK8CBSo09jKdOEy20wlS+X6oYHpR2o
y5gO53osAt8hKfI7maUmJI7aIHeYqiwK4sBKblHuavrNgVXiYt0xU7d5URz1
WxPyOtpoYxIQVvMwZzLO5/7i08liNQX9C3JJ5F9Dj9me8mAUqRnyuabRVrGy
fk3FSMKE/WLILrOKZgMUglJWHc5GZYH5C2J1TR8Bd+YlN6zbLzTz9IXjQgUi
fkFuR4fdh/I1ofEd8tDVfqOD4e/mUInjrp6ME4F0rMs4vqJUjpOw4LVeqUtQ
w02S4gbVZ4jIBjET6Sxj1gsnSj7X3nHry5jKMAdi4wsiNvFnzE7yMpvSpxBa
NPS5wuL3eTw6rfbUdJCNQ4lWO9/8EfjdHYsnqzwznzUOMsl/3CNUAdsK9apb
g3iM1l/FEUbPn7oJLb10NEGjrUr3ZKwS4fd5GQMNMqnOnk+UKVxl7ZQ+YLl8
Tsfjj96isqustIpwhL7411de130eLa+t3UwIStkXL4XMHoim7MHqVYF4R6kW
F7WKf2GElLbe3Oct/8cu5QuFQYF3ifdwJ8790PcexR700EW6GVLSAwQxHPVl
QB5xy6c2HIPV07kYP72W7Ep2l97TlpzKJM51TqvQXcuaFdPuqwdTGNcKS85M
egKUoD8dDg9/oyUqOEfDGloeGdZVdkWOmWPTyrQ7UaEY9YINxcfcfIvHViQd
aU6BaARDUNObfuwx/O8o/BGDAdahHLUDVhwd5IF09ttjtmhXC9EnCmirafGZ
1U2cJeiv3pr0oRXXREJq95Zq4q9syWB8ReP4a0TAdqjUFuViTWarUVdLqCi/
N817qncFFmYLVxs5R7lQ6BAJDXscbC0GzfUJRGMftcd5+/bH4oKS7dDR6GOg
oEGeZtc3Nh2BTsbdrY5RFtYq2QC/fKHBbRaCBwIqNzR4Y0rwRm33zFzgZGDA
4HEbhgmA5xAkfOTCj709J9/r+COniEUIVp6sjmJqUCqcmEnqpSA/5XCAFiwQ
9UIRb10Zpe2MOmUYveKYeSfPPkm+rg4dyTBuWY7IG97i81Fnw1A4PHrskrX0
f6Qtuf8XwUx/VxWahVmI1jgcDDS1+sTmeiWpb8VHAvyTpaz99LtY+cx9FNff
nEqWUvEO1HJ8z33PEN3A+AnAvsmQ/pE/5eTHubcISJuEJmEd4E/eK4W0V8aV
Oa/xNntxmcR1J5Mjicnss4wFG47z8iQ0LSQXXpGlPOlLd5gx3a0u8XMEi7Qm
B0StqwHH40qczdPrh4b4++4or8+2NEy9tUW666neluxQR2vmiUJYWh6hd4sX
CIxWjs134z8ZcBEVIpdd3HcoUJZkMX0DklG7X29509zdtP5C+IG3AXfymhZR
RZNZ62XMxQ1lMrNiziee4vLJ3EY3kZKoBTMFkloFUaZNL8vMxgGxuOaGthX+
edqTRz859nj9X9e3dOgB25UcGUuYfU0sEptTo59NKfi3tFCAq9HbhWT+Qdo6
HoOUmOVHg12UUnfQ3nd1L4jpC8Rdq2Kiyo4faZUJybEmUTCVsBoXAa2TKyzN
hlRrxrfJO1EjKxzZtPdQN++8pkNIPcaprxbZRstX/qviVqFMrRxGNJHeITxn
U2mRJoRdu58BmUx3laY/NAeo74RK6ubynruM/sm36BTY+WyPk+7D6gH+PVt7
BrAbtz+x0EujGVpof5c1HS91dU8ArztKo2Y0agquswDpNKAQx1ngDwZYgWBQ
iQC0X3f01gEyVBnf+6R8D0/x898TCU9emAMwZPyrkPnmw7WV0237Xl2gdweX
vEZyKA72hMrcD8gMvPisx2BdbHODqhsEbyYaIwm56qaDTBTwjAL0T2gaTkZU
dZW02O6qZdflwDdfuIQlTZD//i3vmRQKm0LFC/amPAn1k11q/FdxWE/Ju70k
/677Oc5tqswXL8hbKku6XreCoc7JOjW2rmAfIuMom/XIZdEtcT7Y5IggZMvG
kZr7+aI0SF46zJdcUDeAxbw/AEyJ1kGA/KejoGH851X+ub3xoaLR3Z3HlkGK
Ql46OkbA6BrUSAwGdhb1zquCuKUxdZveYppkiY/I5qbtfzdxPhbTXrWciu02
aZ8DXAuhL8tDiVnE7ZvXxSr2WngSt0NVUYCNevie8qAgZqT75KeQsaovGkXP
0IChn5GXbQvXr6yhqaIRr3tjFmzX7bZTDLpC217Yj9VuMHanxeuoWR/7aK6x
LjBcd23ybBKXYNnEwH1vzDVAwxiKqW3m5icgGWtCqMp40PWhooKRse0Gr8ge
zbPfwKyqwgh5zFwddumTY5PJ34eswoYKmiBVf1eaG+M5/6RBM3NxTZHFj4Jh
4dI469aN5Vz1XFHpMZgVF2JoD28gWie/yE2xMk8H22CjKwjvhDuQx/Mbus28
gTA+e2zh+UNF1EKTfi8ivFPiy2ez3/u0EdIU3aiRL+zHsV7dc4kml3l3gcYk
0UnJiagNQXS1AvLCfe59v0eqozoQOrO0NOTKr6+3RS1fWe4er8sT6mGDrshm
WyORBBrJmmnw2I5iBeq7jwodqVAVBhHSJ+qtHtqFb50AxdK0TquyYIGS/A6N
JM1TpTBKLXSYNu1ZBYV2AdzjWZBqbMvK0meHf8PpdVOv0BR7sJ95PTfNcHf7
m+oOi8VXTNY7eH5VjNcT0uY/Z5JV6LPxzF037qjRGVVLSYXNqKjJfAqLmIgr
5h7gA7EXWJFzuPjEFVXB3hLcpqEkUMqowW4SpcrIWQHAnMz1D3v8uksfZRIm
6Lh4TcOaE2bzvehdS8GHeUaANFkS4dwIDw0ATR0qDwBzv31JgdmfKn/C0fmc
qRSD7c8jczAXj7bNXPoARL94YnOhzeiPLPyfBms/zHphFursyswa5NBfVMSb
R3Mq4PX3cBwTntrqNXva2uZRPpXVt3iz+kZ9m+J/BzL3g35LbIda/Yi55Lpf
k9qOKC2lAspksb6G3YgFd8LDzD0p3wI+xD7vKDybGsjzA+ucsBk+On4qTJQ9
rgipapeLs80MzyWowGRX7lPWc8HxUzoEOiVKFlH1KP9xFy/9YXuFk+lFFUFx
Vv9GgrVCglLf9RuzQemWfITvSkVZScJQIHife/nY2eiOMPTOeGqAkRbRq5GP
VCVYjU6mcyATGMk+m8bd4+iChDi4sH5TpW3n7+2wIsT4tfDW7owVGSeweof1
2FLK7cg84mGF8fGaLyOYOXaFnJHUcl0q/Hl1NnfF7+Ie3O6H+Liy6NCOTmCz
z8xCYzndQ8SkAxggzD8a004qeytD86TDeeDYresFWN8cVjAsXQdINS3hWyq5
6Xb/oEbft3+fJJI86ek7sLxTKmZr85M7szZOhftL1YsU6bm2H8SZD+hztGbr
Sgrmn5vJ6qYTSrN6nM1OGBzNtDDERBg9LZKB62/J+FOK1E4Y8w+BpvlNDpFB
qpik5XJzbLZNHFSUR6ckhkkwZEm0NJUHJf7aEZHdK2kf5j+r9ewPALQoZpU8
wiY8ZM98gdoAFUdhyAyFk2bWIzCbQEpMk2k/dcY1aBmDbVpZYr+UMFg1Putf
Q9/9NdAwWhKG3pXrY0mPzMChp8q0bebxHy2I0uNIDNwd7wwc3cHkedwcC+PT
f7fYlU7zyiQVFYlBfwSRE/RrjRoRSB2k/mL0SDqemk6BnmiALa3UKngxD8xT
sXTQ9aiVRWjh/417EV3ZrMFubmH/H6rvfVt2dFU0Iw0IblGlsatuef2Met23
HCGynGnpuJUiz6nB718Jno8JPqjA/C4tSMklxwbp6V1aRWkzGqiEDZ3rXs1Q
qccd5zULehPZj2mTjSLB9MD+c7T7w761A6jSuNh6eaOJyI4wwKNtKujGj+6V
XjZLtFBPYanNK3i9JcjGahQj9xu3wTFewS8LBGRkhWwX7tEASfFLB7cbiYLx
taaFLd0fTl0D2jjbH2FrKDlcrgeZ0TiPAfrvUtFpH84XDufb761Ha5uLV+PU
P7B4z7IessSwKbGjKeij1FzXio743yVYBZT0pVe00r5digaSPIn6lx3yQy52
5sH+tMTw3C8uC4V1qmQlMNF1XRvF6T4spwEm/e++RWkOFc7Oms2GlZlpOykV
/TYRWuY+CcEMEr/4h/qcV7pbi9y2bqMRGCLqZLyKzCLAhQP8U/iGqV6bTD1p
XGKn6xehbJcF3SmgSlyBJT/smy1Bp639ByyJ+sGrpuy1Myb8VhKuI2KMdmJS
Q/YH30uUwwUAVd7fRVqaEZYXZRelxdijI88wXncCeTvyA51mAMfhZQmguwjg
0qqUVKQIcWfDzHxdmVvO4dNPR+akc4xvZpJ+AN9kj/ooo9wiEGVbkyylKXd9
sR7IkuVmwZMxmf7X0p/TMavdzOYtlmNQrourq4Ku7I0aJg7rxCRbrTOw/yfr
AbNUJnkElwWif2ngDtQzStyeCQUEUJlXdHELq5gzKiB9786pdu7VeNcoULbW
Vyc2M7LZmgVqrpBK7bQA255bVTmZYbDenXa0IAeCPW3IotbjTEz4J6dJrJPk
kPHPjVmctZ/fXWgctNyikvOGwtyFADhDAKah5N5PBXMo0KY/Pw0xJ/AnoUsd
vRGqrIqzUtsgRg+yzWANIDuP2sqVQ6x9bGOxrQkJ8ltPAY9IonFMJDGP8jNd
FMv4Z+9YcX/VMmxnMHBfACgF1HCeLdh/mJxq2LGG6GsArINjrRoZYJFaqIJQ
R6jJYlkoZj0wVhMaiNkuIPHLvknI6+PwvYsXAR9l2Onz5ZZlqILAVR03uqBh
skc0d39tUSe3iX+xZN3zkSNlNBX6Uuoot/B2wUWgzep6xLeEDci6tGGIZbJf
m6vMMkubcm4mG2z8DKqYQuDDroz6xFM6jBExBH6AO+yvUpErr/0xBByqPxoX
9Sc7d4RJA4r1JQXv1lQ6l6ZSZOYxdmzQxMLGCDHe4j8n0cRL/hHbmSm3w9lc
FljmDjh1PhZqJsSsQ0JCLSxBFLXk7RFehol8NdWzZ7IfXypdjVXdwFTywcqd
ICqFl9otqZbjEXCR19QqB2d6ULOkwggSUSFVh6a+7v9Lreg6sR7duYnkvU/U
HFivqhO11i/EtEc006spTvOj4ocXSCMRPhma1nObaZkw3Uwoqewqnft/Fdah
D0KU/68AnuBJNHfGMUphgJvM0CJJ8KUmk1GhBP6S7Eg7uQe+by8JvQFSQ3+D
TkDWnjgxX9bcuhCipiIYPR6BTF/0NMjYMCJjL5lyUKkdJj4riQyjXX4xdYl1
r8diday+SkFUA76KduImmu2OmmfsfwYerSPWn58pz1LxVZZrX4u+I8GiOukD
bYhQa3j6O2CWOVKN+ROB5ObirBfnuRIspfLTiLOUTrbilu3EjuJcPDlM6ADf
PxPmxxZtdHALQ58Pokql+J7tZs7yW+/Q/9JlhzhBQaDajon2UCkWWihEuGYq
GBZAXol9VAVD/06piOSDuL/E6JB3dqi4d+TDKMi4oRglPrKYhSWeeIfC5zF/
zVLrqgM5moRQCWVIu2y/DkX/JmeYMGovfiz+Uskh5wy7xf7L/P6PZSyTKHo4
W5RUmGFuoSXzCB1ZhmKoX8jCX2R4u8cjKnc8WiCq7H+NYI0PghO5L0D8LBpN
cW1S4s3xiakqPVVrDpSTqjU8cB+p5GIkeF9kHalMjn3aYIx/FGIiYWsSaG0/
b5SBcn00yIYxK+iqsl4zV/rdbRB6yppP3mV+EA9UYRmhlyRxD4UzkmD8KOn5
xRFgSmfM4IemP1VgyeqLJxBWGyUJuUgmJvhgck0eEnlUu94rjdTMi0W6jtI7
AVozZ7t69jX+dwUUd38O5voU8+CNEc7I2zxmZemdxOLQysvYX5LnN/UHEdfg
QVwj5Xm5gbJTy93SPLFK/N5i/PhsMMpUSM/wPE+2f++DnsG2eu4Kdzc5Ve8j
1SUtxT9NzzvsglUusUsk5Lvt3+n5lWr4XJLiQrm+g2ag4EK3AijnqzWHg2Zo
+tT9U4Dn0E4Bl2O+hLdeLtlULOt8bEVwI8WmLZqqcBJbrDDEw3aXD9jBIIRc
eVTpC84ujilFZGQSb+kwv+rknHDdIjssq9RWnYmAdX6giA5H4VFzpzhG/57c
0VQyjrkzjOW/cTwZkV1+GVOj4WkiNzeepFzRExhNKaSWwshyHFwplJIqm94f
AOkd3DMJt3pzDqkY7lcAG6JrO+4WCNiQuwIpPFBQp+VrxuBJ4dhwNGkzDeCg
CIcaZkDnKaa0OryYraz4ibZ1VEXkIAESGf+fGuyqvkyljGL6tqj2EfxYrFfq
Ye4dnNh39S44QK3VSGhuRYhB2Can4C92mffqtzon+3ixIPx8udxFdxreF5pt
ppSXucCG/W2S80jN5zOfprlROWOtI0E6wjskKj5wj8Jg9Hh1Grg4u13fR004
UAjND7TUHJO5AfnSM7Xe8iQQcAO/igNuh+fSxZOs0985kcgb/K2M6OZCNxqR
Fnt1VsV96vqGkY2tBvhlScWcPl1Gqrq+IHyJUIvsGXVPGnhYvR2Pl3KbSrhc
xidCrBVS6sGYQivDCGngZs5V57GixbT38Jkp8rNCTNpRgKDSdI8pUTjt/DLh
7czJNq81vWusUmx1lTxqHKUEtNAxPx6UqO9cDmcn7TV31PDdt5TMleUS1TuW
4To0SgheOkFD83oayl+xApjUbREOsoYs+XI1VRAmp+IjoWZfrhb+VJ39Y1pG
QKQYN+JL2J7J6UYC6ocq7nyaL53n3C8mwxBjvHgqHh3tC5YvV2g246SVT75L
cgRjMcxCg9tZKkx11w7gqSB/WhznJwtmuW+z6OniB30sA7imhhjPRzvu0Z+s
cgOADLm9MTi1vguD1SAjrOwrAzFDAsrGAHGt2M4llCKRYx/YBE1cJEU7ciC+
rq2u3YY6ZjLX4iJBNwKIr6CfFWJ4tCIQSeVDjTo9hymljWj3axP2fT7SOELU
htNTrD1kkbuHPQX08S6mQs2mJCpz66ELuM+qVeu1h8DJrB611wUxm9kvxYXw
navmLJG3Ke4ZOF+R4cU3u3zNyifRQ/jClw3urALm2oDTrabWKM7MFMSxmPfZ
nZ/HJEbwKszBVQigGfY9xoJHZ1Uf0kedUCIScbeiHbfSr91c+w2Q3UEohK9a
yIXn8+5nKL+AsaJQM+1Mk8FdP/7qp/+sjJQCy1gReXlVkngrzDMPWBchYlRE
qrImeAVwa958FlC8uIcxW2GiA4+DeFqcxpwoG8hZjS8eon0jnBsBqVKnT1k3
hlr5uR2i89eAIeYWMl1m8+jJH7rs4fw6wiK22WpwEJiGaKslmOfEQl1K+Ni5
f/yNylYeMCO4EEXxz4gA6N3wrj5aaA4TW2PdJEGHTOViZBKiXUIlnlfIEATk
D10OreKp1WryQsMXO3vbaVikvwaGgQf1oiADPvWimxWCevI+ispN4KvyfDag
LrhemXpjeTjuFaXKmsTUGyRgbmIS/sgQbnstTWhTHUM3FyIZTXgztqT5QLed
ihtoZyutQ01H2evSLYTz71UaIphtKRQSvt7tByJ6VXX5/qXOdz3d7mgkDN7H
U3/6cbRODS6LTMMOmztOuw0kMdzB4dd13vNjjE6oL1HjhDJkbMiOp0OMrqUT
O037E4Bryn7ZbJcuKCKqUgpajEYrCgm7eNkZocQSPERUQGc7cCOmrmYinyHV
tfpNbecsD37szlbqD5kTBWX9+rd9GRygeQvg5wmi7pEC+hD6q64D2D+FhMxO
14e61GxWKE9itOxQ7R+IW4gkzgHFMJ5TAlMOP/MzXvnNMFYmkXIM5Tp4xLVw
+PYTJzj2v6cYACD+l0NE3PozCzCZ4u5lCZFgMkv6KFCKG4yzqqQSZbcJSiRy
v3qGJ5KIDaiMPFOYvii11xBUWcO0mcCMdYIgegm8sb6cIpX38WufoQyw+FDH
mnoA6fdvYNKZDy7Z+P6zJIBmInM2oBeSswY/ViqAqI9KjzcqsrsnNLAdZW2q
QRAaWLEKaa1u/W/YvyMiqMMLWa20IITURL1EZXioavj29KyXFgPPBdlpAkUe
6VurRyUGI37hxhmZKiO5ddDr2fSYPgFrJysBFIse8LV/7F9Lz7vlMud1Pl2c
qQDylrRR3w39FAQLwiMGQMWY3v7QrMsojVhyRyPgkvDO7J+8GSqGf0xg69yO
/D4CHzvWzSi6un1tGqUMsvBLbcoXGEXhUxUT8ES4L42pqWvZvDAqmix5LFsO
QXXnL0k3y6mOLHuC0ERxTHpTFOjHBhHSllU8PpAyeQtmtANOqvvlOL2I77qu
fWBC/mjHDQ+3fCL5GMr7FZddrmyRssa4PCD9OFO9F7N5QVc5MHGQAf/UaPw0
LK7fGIgbkiwU/Erpv7EBscoFMmB1hChpdr520TgKrhkrJP5DIR5XE/9vDUhr
exlwYrP/CNsd/dd45fmS0QCcBCz6T40zrLQgchuI14Gp40Zj+IHS4HiXWurS
8Tt+D6Vi1dTZI7cNFD2S0oLYucjihQk9ms90zfCXRJkEZzhaRGrsw6NSXjw5
crqZzxIebwsGWlBzMxUeletTBoG1QhsTxo70vArmfmYFJroprW+PorCqnHga
rsWbmeGdCfPUydprrSjg6kqqGuiDVJzkU8aqEJEiE7+S7RDNXHu0ZcB/mhCc
aGHBpcevgSaEh+EaVr8P4Ywx2BL5nn1mEoPj4dML+aHXQg+8eP2wxR35s/Mo
Ib7ZELImp66NL0MEYnPVkDzyjCd2SyX1UEbVRaPngy3J0eMdkk4KU45nN5qR
TVpxZXYCsi120E3m3SM6bPksfQYk0MkPqMcIqmKkoaCdsVICGvLr9SRqdaVT
6afQ6ycaFzMGjiECqHq/7NwCbxLoMv5wL9iIua7aGhOQ6BEw0Cla+p+AD0/O
GfyQvVDB0suhP4xAaMwBeGozLlC2h5Bzxb+PCfK0DFO+D6UYeqQFM9jrsL2Q
dxO5kpXMkrvyTSfZFghM8IFKCIOBPGZWNbqaTnUenRluto/UPeI3ZnCbQz/J
Pp4JQGAcWp14e8KJYSefNtA33XjSyod+frcqp+ZhcVoNHuOuZCdFcqnHgEFf
YZTyRS6aF7qpuC0O4eU3UwW5UqMc//gLsFSHLJzl6KsFqvj39fpTTiPpnjew
AKaB47SOEnJt0NxKO3C//Q0I2OOeKACf1zP0d7Av2x7rHk+eKHP78L74LX7H
O18so0cdIOc/19k9uqiF1jfrPYwTJ7NJrXfntqEKuaMlkU/TJouIGV6gV9WO
0lUxZnqnLUNdUk8t73MYEqpIPyP/0ehbWvwnIl6t4nGGpLFh/dNsmEcasuic
mZLM2/oyr3EBGQaQrWbwMgx+vX46z5By9aV8y1esnEXk0n31+Maw/fCDt74X
qkicZtRzDB7e9uZLTccZvtwym3kprAln3lbaDztKYmH72jSfy8317AkDlj9W
JNoSkzr8aEzOUzFsiimFMdMxBlF8CVUxxZg6DaEyl8R7zQwXJYhlJn4pq+1c
IwICsxZcx++6wU+wKPa2n78Ly5V5jiAcmYkIRJPQF7WD2mpyTjbNSduFJOHj
1BeqOVL0MkEMRjdvpl2UuxUtJQwHHAPVfMYKki+pgZRhLVj1QGzWekGawOQM
E3JOsEHq+7CueAgJr1pjWqWrhPeYvp9QButN5T7cJsq+nTtk8db1182R8ums
wJsSMvVWVV3V4Gjsw2ZzDT50+eXLMhj0X/93CruJvHmuMq1WHXr1Zjw+r+IJ
AKYQ1mMMUlZb9LxjcXG6mUICYAw3IrBKH4x4JBOvWKD55LApQjAIjigtzaoW
fEySn9w4/yyCN2JVAwNn+7qpcemcEB3nKuoEW+kV53REIGG1e1QQlgneUHir
GxSIoVSU/berIuqMoZL5+0KXn0WxWx0E9OlLN/ZaRcO1w+EPrbaVhnayAlE+
VXvrwMRVFqJ/nfPhOEOZcxAFWVK7L+Gchbx6GkJljoB6jcRVCkec5J5r1mIs
o+1QI9gG6jz5/Uq+nxCuVBM8Bw3/180Re1LUno3FNS3Bmy3BsBjKOF0Ku2YG
6UvW/Qft1LqWMTJOUvUvafVbYdK5kKyBU/eGqA4TgPgHZuNiIEWfcoo9N6cr
L69Jjwhobz6h30rfdFgNzTl8bg/H3c0uM9Xs4lWHT7eSAKfAhrKzjMT97HPN
FR4gKDCGcvAfiQK4zURgs71K7S5EFjjScPW696ZfK+mYQ2RwaGMj5yJzgCnE
AuURSVF03m+csUyj7D4Q3uE5qWd95YWqCA0cBzsVgF7QSkv4OM+jxbS2/C7l
JCOEaTVivgq8wc238nGJn4RoRhZDm08emgIzNgciZm5iK5Cf3a/RDGt5Zd6z
ZQdEOYayBNZlJMYlbDnsuicRWXFd8KSTK+wo3Nv5vK9G8oLv7zqc6gzdx6D3
mJ71oVqzriFSN9Ta+udgL+98IEqHsjhEUpPJXpOCWljV4aEmy2Fp4nGQ5yCv
WX+qJQ73OCeX1l1Da6xg5r04FBQp62PaubFeiWWUcW5/z0S7OT0oRgC5KeXK
BdapVzboD2t+nNOqWlgin3lxsLBQCSWILuHyFbcxvqLKVQq+ep2EWGwxqZqL
2mP5AKmn3gKGZeP5jhoFSqIIDp7TsHY3SoLKlNGGjb/8gsgD7fnsJEguR/5O
GSgn040R4ecSWcX5/qVeP6GWDSpq4EtdHpspP/TzZXX7eojVUeYbJcr0EZaE
KAmjnosyS4gA2BUQXvKsBoXU9K/kvuRlJjQY9XCTW3YBu5OVQgAqKhSu6ZgO
ig1quwAONZJEjRcJaqqL+rTrgRgUcpH7GS5dadzCjvFPt75/jPfML9yf+9hz
WCIfISwPPa2paPHc7SPR3E6X+4Y/oZH6Fquuz9G/vq6i285PSY980H9I4C+C
WvZF05cR483Af/tWYGfmQuTz1a46Wt6iNZnS0O6t0gYjKtgZDrBjAA1RpPds
x33pSpRHhriOJokYO4eHLxzNVbFSGOFaTUbXONmqQys6YY3QCf5KyI/mMXpP
pR7PJKAMcl3NIxLGYI1eUPq9Zr/o7wNhtTEW31xWENdfeCUPSju52qolxd9Y
LBwm2RujlWO8CPoFXSWWuqZNZjSlDKg/7p1hPUmWREtPY0wbV+NPsLn0jjxC
y/1EJfewnfPaoInK6ZYDStoqKuMkz/jjh3gWOmBGv6K/6TFsw8BrTkXF7g/V
itoaqIhalKpA7Yu1YmyKwnF3L/vpOor8PLEJJqdLpDc6g3GrWMCcJQ+CBL5W
Vdjd6J80g+E/Hl0P1UpGMkPAPSwjAng8kvuvF1YoXPtAVAokhnAMQHXNzBp5
KTpccy/r/EBU8lmWDNhOCnZdW5SBe4m7TbnaCeEex1wsWqqP4SrF3ApPsfkp
dkRCXmSK6t/psjsG2sz6h1I5hmupTyo2hMxGBeV7reTQOO3k4/LnLyI3Vg4S
ZpR/4avWrAKJs65qhiCQwemBA+uryRg11rWGvqWZcl0SGSklARPv98hRhBT2
gqBJ6BMp4fYrFOQ8ui4t7hSoUyjYOKIk08TCqWKf8DC0UD4gYnWGI73SQgyA
bzWGTnpnkYm0M/hgr7HyRfU6bc5fFDedVm2XwUVRDlkaefOaSh/9NUb+Ckb3
+wKlpFRLu2bkGgjRdzzcLfzmeNkyIO++JW4v0iUJ/m07P1dB8crzATbff2+N
HG/tAXyRQkZBW1wA55t5POAxN9XOxLscACkWI/mOSWtFNYo4uhkfWntg6kbA
th5yEU1rUXvhUE0iu/erImrJbHwEyxL4+17goRw5NJLsVeASde48u774yQV6
vt6gwkWZV8/T29XRE3D/TpHSslVvJxDytByABdVyhxq2Fi/x9ih/kiYW7sOv
Tpw1Ktek3Bqal9m8/UPQrf8wk1OhSSNngsit0UbB7+Jp0nPGi3RUYWYZUa69
RNz8ztQF9u22UiYe0lYJ2Gx/bbSJEK0iSBxVHU9WfqvRUfdua+3Th4dCU1s3
7H2o5aD4Hy757kfgoTy24L0jo0ZnkLshf80vf2bn5g7xrRr11Ciw4n7u93/H
h3BoHM9T+YqOCJaRpOycQHacHcbK3GBFB6u2SuncXz65yyitzei0FGvZ84lV
IhOfVPLfLS915el6K/q2ObQWoVTFsYvj60BN51xHURC52d95mgM+nPDcQcda
4LSERtIx+z0ks0+9erVWTfbZojmk1aaaVvwCNqM6Shpavkf9L02T011nL77R
MH5V3uSmei0Ncu8Ams7a40addheqfNlTYnPcd+n1ivr525Zju63l426kfYGA
y7pUhhr63p8MVlMKmoftuEeWPbu4DszVK6cskr0TQ55NMtFrHy2Jdfv2Vl5/
if4lj5YAQ7I7aWtYAuoqGlo+if2MQ9Py6jbBdR+BdL271pezfZQkY4NskLb6
CB9nIXeii7hR2MM819fIeJtWbV0N3hbAXA4T1DwIn1PAqXNiNBud3yZb4JQs
GpeBdZgA3/qLm7ehgN7FBogVkk7HqgLac94NR9vT8NZbJzREAD19K5j0SCNk
issa+mVHj1IgrBdFvhotUCg2hxYjha3wcIJsUQSF7IMX7oqdraEPQBPo8YpE
+SmTEcp0eZiF4LqNMs5lx28nHnVU/3+VITOzFuY7QaGs56V3XbYQKxFw8VoG
WH2J3ZWsSBWTyp0lJANjDUW6njWZ1JGz8p+xboClPeEg5eDn/tOORHnX1Q0o
ZbYM+L0k1MJ10qIu9+bNCy4KjrN95oRMYOxCJKnyBbHqN1RyNOjChRGa9UJc
5dELU+on7Mv+yxOjpl1Nx27Y6HOPwGRXySNJhK6vOSMuDHtgOyiLCZB6Y4wn
1QWdrYb2EpsJUzib7rKCw40Zwyg18MoTpEGSLfYhwHz5A0Yxw/1C4xQO7rLw
4eGxqOUeysUuUcTxHaqx1M1to/qAcyRePzIJ6RdLx6La6SrtvH/YqPBsCi1G
YUkFV/djp8V3vNtEP6U04uo44QJiL/lljT6d7kIuaxzkKxwLgU7xFoaP+/Zc
6XVMr8u2eMrgHREH1juK4SsNBIc/ORgmJKYR8hDwe9XPtOlo8uvxXX8c/zU7
WiMhTw1zunvHOLOz/M0gOqtZ5rhdwsomilHh80rxzweskJ8qwjkh2UDdOThQ
vuJrDBun6FDQpg0E8PKTKmN9YFMhdpBuu2UwDH18OgsaYjGI7l+DmWAfRdcy
FVZOq3ihofaD2Z+kSzIXVCgrJcvVHBqnhH035KrIORS1N/8VKWgGRyEShFU4
KYXCHA81WgUO+ibDOIATr2IE6xn1RCfcoe54ERW4yZnP32QC9B2+h37tf5SQ
MYPYGGyVg6P/Pf9rQg42nTBSlunteSbNS6jeTczP6K6a6zSMVNk2l5XhbKA1
57MeYn/+zdKG7RWPQenrwnqcaZHGmFB7dCocgwuoe10QEVNjF8jfmWU5mdz3
sbXuS8yC5R6vTfoP7w34YpdccRCKMvehYW9xZqyPHV+UtGHXXO3R12TFysGi
j65tgFHclvurUAYYmJ/8CtKUoAwj17W3YxdEcSxfsOoPaA9sVZfWtDd9Kjol
5AgPOj7KFxPMAvmBUmTcs0iZR0C525HNC6YmTsSZpefvE2dafzPGpVI+EL9P
XargD7B+qCg4RGPDnLQ9nI8vT1M5dN8SGEBwHZTkcb0Oj7m4eWTAfzKV1+3i
yV+YDIDRUF1C4IgbgsXpYGQwBkr9Q9W5yVBsXzsi4qkWrv8asaYvdeRR6tkH
8EDQN8jn1UqmOPGUSBk8dJl0SU1+PUNH0E0h28kZ6GSTL7Ul3QsbTkBKGl+f
tsWTHDwL7fBA+iI6yNxPwlgGx3C7XIPurAp9G1LRzuGxrxsFF0YbnEbzdG3k
r1xucOT4BsevHHShVonKPyNkNVTQbf2J0CdLO1pOxDmo+YuFSUIe7nLn8AOe
9ctikbuLvn6Y9DlwlmGvdUkZ6+wBo4nmBfyg7iqz2yikt1JExFJsi45nN17G
qlTCKtlEXkldFwHMqnWv6LP7touJFqnkAf+1QaP3rT6+2lhcLl3fJ08NyJUI
hskej+L8dRGq/fJ/33w6DQVgK8WfaIa6cEI6pRPGLOpl0v92UVfEPv4be0Tl
9esiYvbP02wghNBD4lz6LC076H0Q3/dVytW7MzdyqvgreawuP9LJdk/bxukt
vx8PF0g/Fi5OwvvUFIleFQafB6FaENstO+fVxEMhS84UzyiuYIbqCTb4tpjn
okXoN+fZTH4SXUdVmhLUvSYe6d0EgG3/0ujSGsP62v/kSY7NxBuIubSVczRj
ePiEQ+kizI6ogA3kuQDt0O0J963srro0THZH6LtuYkGSubepMKRwrCKkkLsb
YdFX/O65dRkxrePUuwvH+Ozi7IFPLr3H57u6TDw1g7faC/bB7o3JzoeMhnkz
c8lKSiAR01NKPFZ5BDdCBxvJ11uIBzW8zsP44Scnyx7MWLkdZesyik1XNJPS
5UcAcu8pLFvPQC/i2UBo3vxV7LeupYgIQf7t8n/RNqjlelwpdjdBY+pYyi6I
P1NQddMeY5LrdJuK+f8UIsnAecbP6BEN3JJVlpyfcmi1kbz0Cdcgf1Npb30k
pVkmnSHDjuGr8xuU5GbBlGyoM5OgV5nj8R9PCcXhiWiGipXSWPWvwvlGARS6
0odHVOXN0aD5ysJKwp7H4pUedvUmo2sZZwBFzxhdc3lfC6JZBxQjRzeFb2iq
GJFoIdPmoicqDFwpBdwYhZ2KZynWgJJL7yxmrPiPYT1fTywHcJ0McMOsNeqI
WxgUy5S2Jft0vpfGumFN2eU/jTec+3rgW2BDJ0JkBIV4zSmtw0IJHT+dMxHi
kJkJSB341iBtwSfztX5P17eVWjHJAyKrKtJi4qxwtWepZ30D+jhFfpr6cZfD
/yXkmRp1Pp4Hiduo2EPFf1eBDS0+PoDzKDq1zkGYRkmGYLQLnNnRalmMwYAf
DNQCgV4p/AIFRAge03C+u4+AI8plcZ8f34PvvYMllDd5FmxhQu0t2pD4rTnw
FDt3KUg+t1Sf2FsMaN7L4wkrUOcfC0KxAGRPP704jOSZhURGFyGPp0G9VEys
/1pdXcO/E6jqKp2qyxZgvPx93y8blpskgX0LJ+qdcVEVVXa+nTK3IOuUPDaw
TqBV2PS4KL6CTNdMHKDSxoq79QIwcjIGTXh56QEJOIyTO282Qh2L4AvUPHE+
KXedhl/1qewBL7kPuc+3xF7RSCDxlDJcwooEWrq5EhWeGo9Q/k0EFI/0ks6l
ZStIJiAo34lWLNWf7cgZavSRiNPRINXUDngqpBjRRkA4TdkR4PWxeYGO80ky
yc7PkmxlCTf7y+cmKhwB+FnZMDYJkYFf44TuVTgSxopnDywsjAdvm5E+gn1l
SUYxJ4eIKBDCZxQi1eDK8r5SXFboUVOf2525t+OBh/V47XnM0MLiS8vPXndR
xxCV1BguWHMaMhyOuPz9pSOktmTxJHnxLFkP08WCwANdtTUcOce473h1l5ln
SLf/V/dxksAFUWUhI0aT1wLDuBNsTSzweg1ne/uorWgzgWh7XIy0OH0Bxjo/
BqElSgzqHp4H2vyTpQ0EhQzYIb7U5ThBQCs0z9IjPFfWjGxI0d+xri2yGiFT
YARFfZjyeh/5xFfpcyx9KnUF6LdLYKEVbwbmQEQslEdqgBSg2FLcT5aHduIm
LSg08w8zPg36men8+HxtGz3jMT+8zHEbGtYiWXQfk0r1CO8/y1tPtD7/ok5j
G6PfD/pyS76vdX+Y017i4T6Wrs+tqxQClH8bQp1nzTRNh1fNzK0lbgfxUEj8
3VOB/UWjo6Wr0/a/hf4Ex6ECVZRBarFF7Bvwd4DkSnsnW3CHcZSlfLuZuckR
Q7EfHDZhGO53Rha/MMmh2fGMNxythEyocT/9MsWi+UiV8lXJDVy8P2N+Ps5Q
F5Gq5MpePv40iWSkro6D6M+gDMstALSjZWXdJtowCxlgUT2ax8WUAcHe1689
AkTfEL3tdb0BXiG5U/gXmm+nDqXo/uJhq6/SbJjsevqnMpnqCif4HZokIEkX
VnSRUvT+b1oTAZW8iZa2LM8kvl3OC1/VPZeFf+ETqMUPQYQVW66m4lmOm7Nt
tvp3QnjkZeE9b2g7GwVDf/9d2aaL2E5O0y8NU+5ai9SJ2cAxorOd544C+MtQ
zRtu5m9dZLGPBKmIyCKjBlS4oqZx473SaSXTHwg6LI/ZDp1WuBwRF9TV4Mi2
EFs84DrugAinjjr0TX3znrtiEcJz/br1RmGk0um14ER+9XuqsuO9Xf05aMip
XyFhHLtQUwrzQK4MAeoZIHOicyPQLnuCEc9PG1EoyWH5Gwig7dlHSmDYKzUV
neVxdQXfGwi4xtqhB1QfqhFdQ4Iq2QbV73Hj2ClFCf3bTeIh4jTyP32sJo6S
LKZtCn3lKO0P3ZHFjUApr+iwrP29o/dCJB/RkkxHMLDMtNWDoboUHRgWKmYt
CziHdlvAxG/7Zg6PzKBQSuoN9qU+rle92SGf7bohKBydoJ8AMgMRSFUN7Qr+
grJbhQTD4XnHZDmZ+tNNS4teqsQO3rHVfcQS9XHPQFs1T7dgbdk+Lu8CghMd
bRq1ZuMHl7MLS7zgjDD4fz/0PdGw0UL1TdU+/DcM9vZkB9OXFsZgGKqpJe+n
6IHBxnmoQ6ioAH2EbQ42kBrVLjFYMWDQQR3Xl6HeHKYlTddaPnDJOB/jI7YA
fI+O+X6KJTt1txm5zqc3reswdS7XMBOxE0zEZc6Ii8+Hkb0xexG+1PmXo9GZ
apqKA+BV8dBr4IBeqJPLAFKwLI5yMpGNyvdqx47xjiGZHNdAiiRSyfUpSA/z
ymylTEgo/PQSkumHEplY7R+E4Jr89TrJ3w+LaAR7OE2jknCojGDjBD2PvGx+
IcLTZTE9nG1bozc1UJTihqfAKuRn9a9cptq7oPpAOdQniNGhWW/MtJd2KM13
D+rMztPZWivGOxTdh/7QJ+oJ17He3N4SoGHRRDlGzwiteRmaGfXLxMqmt+aA
lwx/+wE34y1f8z1ZPpPoqKOrARDvttLyZqc+VcwcnQT4FHQRvJc02SYh1xpB
aFJSCHkz6Kod9Pm7avP4oMdsYdX+uSalvT/s31EEz7QHxmmO+zlY1BEs9Kqb
ZB0NEgsmOvxVWoqpO+O+fjhMXLjk3sFfORzYSuSWPnSWdCGKE0eivEmPPTtz
FbBVO9fqDrhH4qRQ4Mt9geweETTxN3H/hNwtgScejWI358hV84s1HfjnZ5H8
8fvSBKv31o9O+PdaZ4TJEQEYyUmI05NfKeANcB/pzKez3GspmAn8wl/xQYeU
zkeO2oe9z1vhI7Ax/8x+S4Y8W3vHaJo+bSXBl9TqOSIqA3l24RshOq2ml+5+
2kWnACOi2h4W7t5rK83WJgkHEL0oHod9qOjniiFUAVsmtA0PgTjMLSfPO+EL
h7AESblBQzo1+6Ax7uhQTR+OKzDy3yAZpuxO5Mtf54mJRRshLHuG6vTHkL/m
tflqXNQT2SzXxnG5i6eEn8TtUT2pNGnJmDmM5Cj2KllnlapH3xWwLbccVIYO
046SuOf5335pIRABq01Vo5jJieo3oirt4D1h/7fW99V263+Tx2ShmNqrvxIn
ZWYqD8q9jRFmRh6wJOIKnZjIy9BoMD4tknJ/+zRl1RHnpTS4/kGxhl1cxZWY
EZf80yMoy/xqaLznBwFxM4kTxY1tZKhv9txGJpPMOTTAjLiSja6T+evzn3hc
VY9nQ6enplK9tvfnDD2w1Zk2n8U1HzzAyVZ668+85qLw+TvHaV7JovfqaGbk
eYAlTqHLtJCHsg/vTkmYbQgzIxYIsTo/I6oAn2iuFJ3aG26M70EL5eqHIJ5h
k8huXvCk3BywBr51kavTSewkvWFIO9M075LZ48E5dbDk8Js7ebHB/tkvbD4I
wo5lgEcNKp6GRZo4Od27VaB4xurm7Ug6NeoPOD+Pv7IMEm7yK6tcDSKdhgFh
uQr1OVRRgZ6nlYKfxH9RbggnB2gVMfpfYmymghFONzR7TJYLEEn6LHr3mRii
urIkSI9z6bR0Njeu/nWcNiObcqcG1T2rCYhDSlAjQiXlFoYzi68eAwOtmq0V
fOaAhK9QkPumd2ACqvUNDitrVZA3et8jrwDJn5XItAD4Xnp4mpt8emVPHWLb
NYy9BvisANN476SKVj/h2+ch70o45eJxLCnBI/aNaof5NvsQ/xusnrNkIzrR
5NmqYa3qSUPv3wisajnER46epAA3iiMT3EKjcTPJFlt4J4XMqDfCUlPmeuDy
DUM/Pl8ZchgCT807WegNyMfAETgt4L3kXfEV0fqlDtVhfXRYDR3ORUxoUDkb
60ws59vUl5joHIBx6EsEmW7EHsehOYyx8LcGU+8kJk4PTYKtvcN78Jxf5ccA
OoaYFcLLDd2Yd1dFNPqDT9HBkIdgADSXnCmt/n5EeBGHKy/KnUslacNYfHdn
2quHoX8nNu5Yqvek2iy/pfqeJ1ZAykJjyDViC/rjzoScmNt810J448ubq0uM
tCl22XK8pjohdIVGzoenwjjINqil7AlMVn1OT/Vr8ek8l7tIavW5IGDUvNyG
j9E/UCwfdczMezyloRWpWEbYQKaFPwYyCMghPkcdNt/n3jL7z1U3hmGooz0L
gVBRTcCbW42EcytmTp7NE1ugwFkqh+XoioXdmgzEbItIq8MABk3BgDbztgnk
Mdo/8Rmf/cUgG84ZeObRBiTOsYHi8o+UTEyImdCiNYuPdujU2yzoaIVrRnAc
GriDx1ryNTVpiIISUACmacxOrLwjWnvM8PUjqoAkBA0A/CoadxlPJkBhfbBo
AWtseStOY4yq/3SdScDwpQl0pb1i5V8By8oxnOlfaO6uTZQUl2VkjydUm8an
31iXVl0VNH/tV7kr9JzsLSqNZdp4P7fhefEC4MZXENIgAkqzGbGfdZj8bojN
tU32cEXM1lmWxsW1KZPq6A53qYgYPUXnb8wKKloPXemO+hHnmwJX6Lkb/EVp
Hw0j4dDMKEzL66OiNYkCo+jWx5gMXrvqsxfs3gbEMp3OIk0Ht5LRIxBSvCBK
INcfRh1d7wGIeaC1Rh5c8ERTakhTO4l6MbtRPU36wYmxFVu6l8WXOJRWTNST
Z0zIneQwWIQoXmfm/u57Uz+iEUo3hzTzdJaJWzq23c8xdHv2loa4ZCQipfqk
5eseR9TRncUEnQkDM41XIVF/tgWX0sDoTaph3ApISPOiSDvbrBjaOXImZsYx
RbnlJIIQrRdwqiC2TrOsqYwsklSgDYj60thb4SBOa0QjWFOA/nR4niKuU/v9
Nm/+ZRWN76zOBfdwxX/ZfKMtxU8SnmZ1tnRgNkRPk43r03ZaJNmmYXZoYpDm
QyAk/6w1hML0YrwspX0idSTRgephBW8/VwYbHPwQvDbyEt7fLyAh8eMmgRKO
x6RRp6rx4jF++phQLb87TsGBF4Y1jsB9UzSd9fvBtpGoU4ELNW4Iom/ykFu+
yRSAEqMPH7/u67ntrCrMD47iMgFoYUbIruc6Bs+ovrJqQj6c3bkRByAGoN2M
koS5Nd188anmEnupryAilljH9cyfXj6lBSE3zMVa5EzNfTnKdPTEct3bNJag
vjNJYtrTTZ+BH74jF5QH0eALzk2jPNSArwJcbXBVESL99QjDfTy5sku3L6Pi
KLixX2oiN+FhtOU2psGfmX3lP2iljifD0CqRRUCdnwg3lfUsRc5hvgTV7ExT
lrwsMypsNdP9Hr29Pe7aS60HbFHdVALwUfZ46x1iMUuNce7rKkwWuN6tisGJ
C3Qed3Y4oa/kxEAF7XlogQSJrG/zoR/+y/kgHGEqDt4wX9U0MoYhBkh5GOLE
EauZV2QcWcyqiTwNHY9G5upeXTlvniH3nyvnGfiQKxF5CHvLXgsdnucSxYei
HNVOn6nK0NCDMgc+q8K3Thdzk+2dQzGb7uF5wrDQ8OrrkMDOkBvFJvpNTBVd
wXVCquy0FbXYGWkhIuycF5k48yIZIZj9m6UVcVMIVDSXZzHVk7HSn/YFpxun
NXn0hMsttQrewLsVZhQW0qO/aCKyTGWYB5xZoHeqkoOH/rQ8qm2PdS+6xsnd
fnBTi308/34b/rTTzdTe1XiJv+pehJ+LnvE3Ej5yZdu0cuEPQHvlvea/je+j
8KUzGZ/Hzn/7CNMcIVJvRiuLwrInlVlPhvsdgu4Iaz/nmAPj5RmAWFio6brQ
GiGSkC9zvalMTGX7WrV5/o8/Agllb0Fum9HYhx9qlMLNmLp+lec4nQELHVRR
oY+qqxej8LbUfAwnw2xeFLhsKTYaTE/ZemrK4l4pkq5dCHw5jeHwTiZ9vpX3
P/fo98l1WXVA0s5mwCC3uZ6GinljRzJjgPV3hHoX5tI0MbqocwUCfudDNOA4
O15Gsfz4KhWsHRf7sF8vjrN+8zGn9ocq3CAofUNbO+N1EEkrbNFWZtuiv3cm
VzrP2jx8MpJve9P1fCXfXvKUUOkSqFg2j8qWOpu5eXVtZp3Nd0nPL8hLTe4R
rt5JdKq0DxqLKuUNMeZtQZlgMp8ap9XaI2OxQW4pPBh9JkCLHlUfkMePy+FP
FZtnmf1C1BBP8dEylQISgrKeu1W1IMVWjKaRIJe/jS7N5/3L+ogXcw9Wexr9
xdCNG1CGZT9QeYY++uC8qpbg+tzhy5Ns07NAg8DFFhDYIvwTATpohoNbj2FG
gy/MBmK1ZmBLX9USZcav0VM0D7+P4hz6gISgCxzLd0XZaDWQSGcygCxmJIP+
QHL84dEncetsi8x5aoempfM2Z+drBKeKjz3y0dYh8kqhsbRp+PE8Q2xNmuHR
XjCqy/mSclSBE2dNIYn9BPVq/kMpTj8svYSUnqwi15E7xb8aj/2Ji2MlOM8p
x51dpxEwdk9DarwEnsdgbJw4R6xSJd1sNIhVNjvF++dKlPx7kykT4BmEBz83
Gh5dBrMwsDM59KaCRgNmjoSlVCwZx9+a5TzqRAYmsopX072JxrZJzEzMcv+F
U9w88TGFebQtaWPP36TSK+48DE410qx3xbvZ05zSi+gAol9ZmYe2kr9EMN3h
JM9/5tf1Uaz6+lDREgHlficljR6kQTxKAwmhJSBoKu4W1bpFw5nAssZQCX8Z
RF7wyjuYiQCSS8g9HODS8i9vXDAzXYw/2lEZzOgiQQ3/CrlR37iAL+0EQVQu
FqSTouXouet7S0axSWz5CwtipgAU/CNTFxTpGTngcAOMaH/0YDbxg21V1oIy
1WTGKMtY7ESPUIvf8vlr8+CH1LaejXpSj/Q9RcBhU16gm+rvScQoM3Zss8md
Mq4jx5a29uox+Ft/vpcI3lIqFcd1ZKouSk8r/nQcKlNnukFTMu5uTQEMsqRb
zK9KkarLocWOLH/sx7W33z8EIWeHEdon0edlnKpI7JdKINnwnMzz3bfIw9Vq
DrWETE28n9FWwKIXNvNz7yD2fqzKe6+WAqOhl2ysnyAU2e0Q+t9m9b+zwfqn
QCKg0HaRbKMab9iDiCxCnCqwUifjrTxug8oJt+kxuhPZEzPT5GmZKJ5Z2FTa
SK6OaGytBRQBcqh7h/YAjqVg+JGjmZsR1SpF3KlgIEs/c0FyVV2dCjkE0y+g
3q+p2KEdgyexBScV7dhQJ+uNQgMXG63hOmkyeEPl9jmAnmYwKc/0xlar+w7V
kI9W/8OiTRcqf6hrcC5zde+bqaperG7R/85CMQPIoubR+YigqRvubHRQ9aXN
uCNhvmaltwtFLWbSsRaV8eaf8aVeQMGzzpqXUrmAED5p5rO2Fxwh4Nv5zs+/
YYk/TB29W/o8j5+BVGcRwvEsq9HvGEBwZH4InBV8YuLE8jb5ziaTY7NF/eBa
cW581Ox0FlUOx5HFKa6a9gHDcw6u87a2Ws/vKyTWgEGYMMByIXRdRyIXJnuU
9QxmX1fEpFIQ0mn0t9ZTHqnvIEVSWDmw/bpzc3uBPuSp8K6trwMYV5nc66N+
zm/Ow/5YJhPpq4Ku0Hb2lJgNm75x8zCnfySC0Tt1iY6ie0i3h7XNApaNqEmd
wdfW+ixza6V5a2wOdI9xDkLxu+YqqoYOYGm7I9ZvX8kRjsDOJBtDujdt7QLd
fo/hiKJ5oOIm7aULRLfaBjidR1SgoTBqmB2E9Hw8eas0cX3PDnrZaPSNQwFI
ujrhwRD/0VwVV87TOXoPA0Ct0UUco32KR2/lTknULuDO0Z2HShohyJAM+ZlA
3i5Npp3fsW1dxapP8HQwk6CTyjc3IKxDMkuRy/btwfywoOEVndzfMuN7HZri
9I4uaDMuq0exwrsLEAcC7LqPn2dfQbHJWU3ggc/abGZuwOefPISh4kb5vGlc
jCP6wN0o7R10l11V7+nvgkHeE816Nj/0w74Y/tyrzsWNSM8vvqYRnayanD7s
cGjBorF+mqKYHQzS/VSdYOVvop3uohS863VejbrdkjYgi3NneGIOC2jVDgfz
D7R1cxx4wwxnedkrPGduQcRGV0AO3hXqXGe/jXRmBtfzRCCJ2tMxe5YQkrIN
zmW6XNfexxCS2x3hsWA1CQ9A/wMhiSYL6g5wUcmWbKu1DBFnluR9F71l0zsj
XaOSdTTRTbrOGZ0z5veWmsrqEql07TwemMDNsEm6Dj265R0rax/HBJnYle1Q
qT7gMiVSbJERH7DoSX0zVgZFDITkqwRfXKeIClPgigpF+O3GQs8yu0jHV+Wg
GqHVoht39UBfMlRsDpyJpJc7Z82RL+oOXMZ2WdZSGwQXI5n4TtRB/XtcP0uA
bQglezr1Vq+n3UM5DiAL/4kCnOW6OiJCbgHhIr1ltVqtJoDGVKzlXLKQmDix
1WfBNmiHZKPkx1nAQx4StGxdca2UYXe036VD8j99PqSPWYx49xCql4vsEp4w
Eq4dclXQbgZXlUS3hnMRxx09QZqrrjyNP4dYLhwYdwrHHGGHRraeWJYwnEjk
3p/einI05iFB6KzPuPeflXpmYwG4GB7WMZzlAZ4zH1w3oa21EdO7W/Q+3JvO
Zh/GBlMQ84bfSySzPW8QXcSiIhUNifqhbuhSCYxy86oJGjZRIQzcaLdFfu4e
fqnBOO9Wxo1shAc1izMOEvcL68usx4fvCsSU/Go2Fi/FK8wHUZDxcpK1SZDD
Tho+++AXH2aNx1/OawImTmlGQAeDeLMH09EQChCyR8UW9QZdD/dv7ICJVuWn
7MgVBwp9IqYfdkgv49JFxP/iror0rDi6th3C1bYA15WRXybwclHWdtYIjPU8
qphPcWD6nG35WL6VWqO1St346QPsiMTU/XCxwaZtuCZIfyCvIDmULlFFoXnV
L9vEFQtF2Y85QHB+44QVnCCJlsz1vvfqcBOqz0iZ61AQQN8THA8jJDxYarAd
fRh89r1lftIrGqsf8hDwkvOfvPBC/+RWwmKSGTqGuBenbcoXNxmXtpeqJj0Q
GWISOi9482HoxiGQfICLkRHJ5hhQ6WWa0NYL8gWyyrGsIwi90a0KkP/AIN58
70Rkp5gvULspiDZS/NtCoBcXhn3gm1bErf1jN3+cVieH4BYqUDTbRVM5bnHd
UrFKyY2SBcx6oecTK12jF1lammKi5efiFM1mcZiHG2hMMq2cxChRps+BMI1O
RkEDcme/TMFuDppn6Vj3Y9UCt3s0LpWVbfwB73+M3qRGPz+Q2qayfg5ec3hD
4OM/LJ4mTZZdUkcxNKOFBo90V1guoh7BI7vpNLpXlP8Z3k5XabdxoT3GcT8w
jAZYmVzJPcnpkhgwFdyH35rbY8tD+DpOuIBbXYK2ao40MN+LcNX9Tg86B4hp
GJ+zZCBmkBxQ2uE2uXPpAPa4tSTckTRlByBHxV91bGxQuUelTJheMh5XgI76
RnycPRgqHHrsIeOatEq91YeI58m/aeBW7/SSI4/CxTPdrvkzbObmXdir4i0N
TbOCwRA3/xH21cYS06q4G/59m6W+JZZ0rDjSiUqCOEUE3hsMQZgiQ9VxGFC1
Ik5oLGXQp/F96Gdtl8bwgnRP3ZBUOz/+GrKaGtg+YhqK0LHatExgmY0st6Wq
cNF3dRMZ2GeqAvxmCZyiuV/R25fs2SeczgF7+5YDceA9UTHI+U/Th2KJIore
blMjHHLE5nC2lmnlXm+fSetN1xzdTVeWzXoa4asAC8uu/eTZKd4i0dP4Xrn2
+dr5bYXRC2/ats7ClQyw5e0afCeiDXK7fLsgU/STOTeCz0JuaiEiFYd8K0nF
f8CzRyP6F+baMnH9Ry/HACHUWew5j18uMQgI1Oh3QWnCgRFpDAireP+qZITT
EpGt4JnlYpFyJUUfjEPK/qmrcYOeXqm5NMtOnymq+b20qYddWHFHuhF9q7Od
vY8u+H3LcVmLOoQ458WVD/zQZ7bFA3Y5tLypfydPZafZOsK15dFz5+VPm/nd
dl9rypVcZqthx/h1F4Y8xGOicH7kvbSyvGe6POHVoHft/aee4HzwW4Y8z84F
rIrkImpc0H64+zUaHLlicJGeW1TzApk+u7nBiy9Bd+EOEDwR8W0qY/TtN6aR
U5WlkDQ+P3RipIIOeZQkmdKiqAj980hs59IpFAhCJvBFOwgNOI2nIgQ9wdiP
CdmpjEmZeKs7UwZkxY0waTdgifW1wWolwPBSdxs0SOWIWTGNgyLEHENO+ih6
41/VpUo/pqUKNPqPT4KVs5HhBJXKLq/8ZRQhVhNfMCLn9zUFt2ICF9ngkJDQ
l6TwGkZKJxS37MPJokjUwtOoROZ9Wol3357njidC+8Sq6iQU5iTszeJrtNzO
ddayYFBdxlPxBgp/LlNTszTCu/wI5PC/svt61Uz2eY1q/W5d7AqoVDVLJPhW
myc0PfdhWU8dLNwDdCiLQ9Itybba6A5T9JrqAfwB3wiNH87n2gAOr2nBu7sj
UxQz7Em00qWAMr+HvkIJQL7VrN4kliusgDUwHUxajpMlYAVpkIbVjnrzKN9A
Uo4z+LE8kjTLQ3B2v0t90s97Vl+C9r6Gti469Q0JOqChw82dG5kyciiEC+LU
pcKxYpEcxq4bP2SvAsoGN+eg4t7gXCzk8T76NZDmR3UkoxR6eCUH5dthwvq8
WY6fDDQIBsQcKzzjJkbgWZu7VWyxT5Xrz55e+oR2rc4nP11xEtPk8XvSlCSq
gfswtAg1Ho8PQuVxjwBDrmAPpDqCTeCxGEKfKQJgf1NAf9maPprLN7IaGF5d
KmNCRoZrxFmBVU/Y4ZCpRRZ4nojy1rwAwuIlHvsMXWCvGpXIAA5KyX9O0enL
PfUwdVe4bfehzWt+SNHg8AVP/lL0bKuNOx8DsxDuVB2Af0TgM+TsWCkJfwlk
M1fLoHRKt33MJ5RkCa8su1j2VOO6ue4zfabNgeCR/AiC+TVZoAiXCbnoUDPB
ADeLg8m1TzuXzFsnHo3bXP+PEwXhNfjZbFev25YzrOeYYhSc80LSJUkdm/6L
gW21JTrf2o5nBzAxxgNOME9O8qBbVZUU654ufOjTjaYbylcV5meixT+QijLY
qub/Qzhfp99J7ObaZB/GXZDoJVmSOabID2Difwx/ZRWgUSKZ9IN8Ar/U29ic
vBWHBtLB4RGiaepaCVjC217dUUOtwv6xBkc5OvpBRJFkMDOoCvSwScij/E//
srRUaMlArUVRbVDhn7knO03kGL+89od8woDdnPSB2LbzBItt6NUzUQVu5Qvg
poXmUlB4nQBFVEYqoYvC+h9regzhMuzzKqM9Qgau39J0RUvp8e80hqbv+e8A
aDRPFKEPPrYjxmVRX2gBONDlphE4mKsawzmMxXB8iisS4UZOb1/xPjpkZ04C
9kIettOs2t6Dv04MjKzvw1SW3l64a9fCLIfNdb9DjUwYin2MHO0IHLv7Ps0s
KpL7dPGZbmoxHgu0JTxRjb0WNcjMaL+UcsbEo6Bs9CpH5OCaTPnd3Xa1zwWB
rRhbNo1cBKLhL+qNqIgyVKSjeuIyt1UJrwXa/48NBqPIUClMeCX3wMPe8fcu
3PQ2Vgr5N5nyj7haDPyBf8srl0J8/AWo5Cd+DHHPgA6/ZQ+q1Z5lm+7QO+H6
+Q3J+v9apT7PRduaBhqhHbJIq02AMIx/tda2n6/7VGEwzlF1G/db9HSMEo32
2QYVDOqqtXQgDx3WwCZtwZLts0W1gwNZl2jA6ipkcm+ZlDcvWju4t8YEPeos
OzLAB0QXsUynjm5VAjmSXKBzvQqbjFCqnHXEraQJVdck5nnZ6ysUeqOmkWnv
IAyphdn42a3+jbvs+MZHuA72fAfngdZEk95EA8kis98StHdtvMa8nawgiH0D
KAdp43EgfNRn8iQSoHj8oviTMqN4BmhCLq1pdg7RGZkNQQqtaLCZ+SOrO3Y4
WYT58YTIL0ZYCHaINY2var0/tz52wtGLj3rmBYo7vYgIIiAftX94VrRDjqcL
nX67Tp69pTAhoUlpUf9bQUeIBEMTFbewHHTCn3pYQXDb67wfuDTg2Pw7VgHS
UzyOQTpwXKJwi3lLCK2Fdflo88qoR9UoCz2Dzcgfyav1j+P0WyUKYshu/T4z
gOx7pYDSEpuZCUdiPBIfz14dM/aIwFOsRYXyxZgdHjVSYdEfxU20xz/IzSP6
qhvFaZKOF0UlKw5iUh8fU6v9AU4g07Qn8rwfOlljOiffvvYIVByYW5QFL/51
XGE+gffGcQYfcOJscT2SD/OcMCqBY0oVUX7oyyegaXEaVg0VUAVXWh07ug2a
BpvWyXb1SAHRZFqa8CBOY3KTzvhd7CQ5rdfICfcTAsg+4Z+CydgKXLsZzvAu
VLt1qe7pdELiq0oWFeAzzSCgeZQC8FB9NtVn4H9N35wXuhXeEI+ztlu779D3
H3i2ss+jpzDawGv9uHb91kRQrJV6E41U68xJ5xZMMgb+Vs3zT/FqM8GrFLK4
XELs2M37ZVk2EAwEvx55X5fFe/LqYW+c2XKcATtxNQmXyNCjv5QGONPUeSLl
XnzJNp4vJKMyOeYKvDRZll3tN0JnbMtegsbVy89eoby+2fa+dxXlf/jybyuu
vWyFghvH93qp04t5oV13dG2e7qCJT91VFZnb9lWjMmf0kNYoxkP33Rr7DeSq
O9VfGWAi1+LA44Cr54g1usJwnoHZ8rqrQRBowRwkqgpAgsena3M2L0vnS9Wf
1PPUp8tCqcIU8AodHog+rEy4kc/iZIpJatASrRoQyqYaq8h16GfJlCZLdV1Q
MEaw9qGBk22kgeL4wSAo/yxwUzuqjOxkJBr3+Pk470V+ZY+3/15E/ywo9gka
DlM8Bviw3hVHWteMCBgOt0Asm+lTRqH7uAWZrjUlr51Xyr5E3vT0SLFGN2Zk
gir6n5MTV49PEPHNUBQ+jAow5XrM8Ks1elECJugjPm96IdfLfyNv9svCkUk7
gQUpEDAVGy++u7ySONkVtM7f1emDXoqxSl3XPcGgwEhhkQ48VX/WD72sNckI
871Qzdw+sb9mToiC9rX6+F6Tf7HY1c46lhkfVcYpcxCEtrzxZyYdVq2kLVjT
xaOKty2lFqkgemd5x8/gATwgAAiRebzcTDgTMDxYw6qYTlPx4qWBvBxosMjz
nIbI3TOnvX1pzouNV+/6ybxFy3S+lgkKyBWrVrHpQhi2Pz1fKwJO0dwlNDjt
pKjF1wnP1mP1xGDuo1OULiA9mszHd2GBtinS3ypSCL/auyCslcM7TIT/GFKo
au5JsFhetBVvuQ3LvCr/rNM39SeQrxPCxnEGYxrDn74pLCgxyDNVDneLGxwQ
EcTNyBw/PruZghfvBr3YfyudhbGkFLdrHybjlC2S1jU6FKgCccfv4y5zG0Tb
EbHZ9Vgd2VoGf0BmhoIZBXuKg+xiD0d6dJ9+R14hixR8RZ+MD/rfZxxVh+IZ
Lnp+Xs3HzqNvcLkXn7yIGaDgDnLcHL7Yhs22bUq0gBvMzw4ThexPcuGQ+RCU
uXiS7iSd2tq1r0l5tTU1anmbvnc6iqZxqW9jAwq7Bh2gZV7z1juFYw0I7Gvx
4mZsyWUYR1c9JY+UgtJ8cJ7ye0KPU/80hi+q1BiDnmefe1+wxQguQnhDkZU9
RdLp4E3sBD3PfTT8i63siNq0aQJj/FgO5Vhm9sBzPOaIiP63MIGPaGsm/GDQ
yNLwPM5HrSnyJ5eROAXS1a9+3E06gJttyQ+gQOR6gnBbBnUqULK7RY31mnpv
tpDAdjsD7dAidimo2QMhu15keqmhbhaVfPX0/zk3k8liS1gdOM7LjtO6sxdL
k7sr7mh88BtSs7PsBIYm7fdnGIPGmoF1UWnIGSd124R2A4bgr6lXjIXUQjQ+
WJMnanIcl/O//6TDIUnJO1Hg+xvyAU2s4VsVG1g+yJAjoHqN7EvY3Lwy1+WU
GL7cPp6Jrq1Dx5eQOLIQY7+IqFjZjZMnY0Y1eCQqBL3Jqg/I+x6sO54mltYx
4MkENOEzSQjsFye5EVcHqE1fDo3/p7wxHNNZku1NMnkIgE4TczBvR1n2KFbp
WGgS2dw7X4f8thsQU3vKK4P6n7fqZJG6DgJRQSrxU0p/yR6eTNZbx3nJTjhG
J8MoROkFKHxcYKBfAt7XRt7EDtpQFhx5wclSG0GLg51ol62tt7LchjFaljJH
n5+hmNpiiC1TjM5WRUY2I5yqU05KMZgqrWngQk2iriq97cpWCskVfk1xHiBW
hUIuciEET6EjiwSCPwo7W0AvsHzPT2Xa9l+wo7e4D1Ygfw8HBZKIqiJ71AgW
QRG7l27bjdsRGXojrR8NhtwDo14F1IXhYGldmV5EDM5qI/d3wtp77XymgkhT
28kprhfb4dNAm5Ag+4GUiGlhlmbkW/NrTHbfGh6ouxkj0mSrrqpd3Nz/OUj3
s74ZPg550ndXzJh+zHvi9KFE6UjeptsyDFF8j2hgjaAed7+LAMGpq5r5RNag
ODvSPzgbCSo8sKzTzsI0EvZWZ+dFbNGDs73B7x1lSfz3Z8NveXNwbzmcOSIb
1ZawPG7UlvtzU6c61ZmHCwpObWZa2P/Q5vD4LZxf9ViQNr2YBmmP1A0J+HlX
7B+BiZnaCIqavBviVEfNo71FWCMW5DfheN84o/CTEVLCEXuYtW9J8pP12dNY
q9w+SgjaYPiPV1AdHLzQBY77hlfD409M2fNkuursDhU5z3ukODbzkYUb+Mhc
Cvzg4eU0QNAOcnDJkkPqklqcUwzP/A1aM6TBFK8wYZL6mM+gVVgllQnY9arq
pp0+KunMOIxu8GO68VAp5fM1DORJzevAZNomUbv65muU4gp0FJT/4WyLXGjZ
gkgciTdYbxhn8AKEFMAeb7Cw/WQd5IcCnN7MQzUOG5Z0dG9m4kGul+fQ9uN0
qfUbkn7k9w/FDl2WrQ37Ymd2ERKrsHqgqLoQEIqCmCphmRrmgv9ILKGRHhoB
QcJhMLG94clubFZZ2tQllM6eMs7555UyVyYz+o0MWp//uw+KlPr3HhrB3OjW
aL8FbX4Uon3krjpkqy8bw3qobFlUuQ9+bp+qBk5VGidcygo+cO2GrSxwjwi/
tHSmipbdrgFgTh/8RXgBz3SfdB5N/LriKJiTaW5v02vzV98kmmLoQEEygZ6o
3hjb3LTxFdJ6Enexazlv/+CiGzs1vvZ/sakwVvl20CMRLvahLzoqoz9DOMG+
LWZrnd72DJ8kHqMTYH7amKRV3ZJ5F8Z+8p9a/Ji2EtsBO0V1lUH7hawDGPkP
cr9zivgzRFw9/KKNwSmKDvKHy1bb8rrC+BXGCccqaBvSvbI/8a0vEuiHe3VN
nsTk5ORwMd8JTUlbOOnFCwoXIkAHRTASTEFKP/DH6nLaSqs2U0EzNHfDuQAP
ipbHowUTLwhoxvz2FgsdxH38Ox8p4EYcSAQ5T7ec0JoF7Zzio2fvEOCq7KtV
T4dQMPYk2H20W0qaMe5kmTlFOCHhDtYhxrDLsunemXlCmNtBT185OJWa8oHu
eWvU/B4J1U0wPDG4tI7n2ghinGmD1pPxMc+8eOolIiCYkd/Gm7H5WzvBlr8B
myg7tWwkNm0MgThG3GoTwMHhAeWKgrzshfXCdB61m7Z8yjUp3LVrYBxEY0LO
QbFv2EseiQPQkx+2vqZucANdr1UaSJ8q3bcKE2vmKdBtPEGwkGLMUuTxwIde
tyoyp1vjRrw2+blFTi2B50rEWeys8lhxOzrBrpjOsrCrSxwWuBARsnfWjKty
J3vWxmC04KwOZmd/GNeoGywxA4rZx9uv9TScdkoLDJOGBnWi09c2DiONyN8K
V93/PZ6WKmpZRubhdGpCQYcgs9p91ta0MwG4QXxEKJVxPhSxEhM9M+hQAEZJ
gCwMiy8UQPae4wO1rxANkWc+yMiPWkxEv50cm69d9ZZLBxxOwoT8v0f+oeFa
s6bfjWLPWmgZH+fcihGPybGi9FLA6fWyAhjwACYa2nqtn/VwdhcXsr9UTI2e
gBI/JU85Fz+pajSBMML4lnCcgDiROfx4A9IzOh5mLeIR/a5xGKu7L12AR+gj
RD7JOi5WCB/MH3k93P0wwzpERw++ylDWICvdfjEF+ryc6XTA3Q6n0OHHysy1
DFaKvcffj4LOVYjsqb3wLFWAJc50G9EjCU1/WDy31RfV4XRdVVB0UMQkpMOc
NTGTxGMTEFtftfSQGyVzCotGTb69V2x6d0kWuSruNSPbPqrOZjAlErnleCB8
gVqG30yZEmLbZpQ50pE09PafhYz9yv/SkTej+OvJaCgMawT/+V3EZ20f1JZ5
T1fJxm4TVHz4K7UR2+UlTLBP2O/IXspoPPiRO22XPtksbv/7+oM5q9ENeLU9
lUHUXOXsrKGMXmmKR/lEfkTThmH9CmW0WbamY/KIC6XQodouzVyLTU/iFbU5
EDYWyOAYJVzdasD6/f9vz6ZzNANgpeSHb3kANaW6I/f04+BxBBb2qqLSiUSg
JAX+0Ikiwyif3jhvKkYh0A3BK/hGMKkOBlrxICrY6yZ3Cqympg1i8zM91flg
zUqm3uCNdgU078jl9AhEvYLKwkkNnf56+Cppgq5GatHsHFy7BjqfM3XlGQLM
CZucdfULZWLFozW0HBBHppMmOnS1lpdXO5bbzv9w65UTG5bFNpCNyIqVn9ZD
s9v2RLWPM33m8SpUZvRLRVnavxitfgV8g7umstT0kwblKd0MTuvCcJFwk/f7
MolDu2FYiI+KwWWtIW6KYshhHobbrHCQmpRTkf1gBRnbP6va64gnTMjIGux/
3owDfmxbWdekvQD545zap+udUT+vXNrGzKENz69IACVYMryLA6Zcsm0IETzX
NYSUFVQowrwoJo1HLEU9CWgryNnjL8ChIB5LwWJXVJqTi+oEAE5eW8Hw6dlv
599n+TiUNDYWaNpRsbCCZLYtPKSno7R8BeIHrVfm+WjdDuG9Dc9LCdaAcdRY
9VaqX5LNOPrCblz/7XYGJRaCS1RHJxfnMbB696X/hSQn0UwhDl7P5W1QnQmN
KuUATZ67JxJ41JNS016F/IJdH3HfP6X/u6itWf4SLjMs9iPrRwHa2LSO94Gc
5efZNGIBVFPxzKLgL7KFpZfEczS0weuI6M6J5d2OBAlufDArAcSA20DW+KyD
LINSDCj87vnQP5dhrd2fquOV9ThcTSUDo+Yd2lh7vpC8PqETIiusRIQQK1h6
3gaMNeKWsbs7FpEWQBx4dLl9pqMsHIBVqmvcyY3oKlo7+h7gCXgg4UedaElt
/PSFQlu+Gy52wvrhuQcRteQ0MidV6M6HA7huGBECPatj1aGg6n5n0PoBrNGk
L0LGL5Dpp3SdzPjFV8BeCzOwLzgJU6GA9nVWskht+3ah38Q4QKMBim0ZGWPh
dS3MtnKhFywKIIF8RI+wHs2DuE9XsAV3XpMfaVZnzbzEQFXuCWXjaOFmZRqJ
CvxlaMytZStTIEOei/QxZmiugoEpTCz7A/MIsFQEpgq/4oHaIXjxW5cPiH2A
ip/5YkDtrkzXCpiiI2ANdkOs8/DoLqOwClcoZFYgkQDS7xbBbU+5fobtjT0c
40Yvuz4qW2neYUR4g6iLYAkofqbudJqKUXtr/Gr5RTlAUFhkScW2DkoAymuI
t/yuirCz4f+/owpHr+keZ0eYqyv16U709+1biRM7tX3/4eAVvCZ1MQWaZ7zr
VBulfII0OZ8JPbYVWz7Zgs3SXr5HOLrrfavxMtr2121TQRt9cRPiQiyaKVgo
24qtuhep8MhUf5b8M62CrmI2WdaKtXT/4M3XDujpVDJY4txVkl4c0DcZGP/W
d1lu+Ns4a2/WbyP+Uo6KjX64QEQsSsmHLEOdedCWTvn8AjG6uQQNCMF8SAxK
s/35JT5x3X7VJ9O7G1KnIhQtPy5v1/b4/KZenb8p1pl9znt+0KlpydSi3qmn
NWA9iljyQ0Gt4VsZqYc8tJdjXNLFGt9R1koz3yRvs914vqtFZJDk/wwivGu1
wC8QvrG4gvjBMllCkZ8qSrlWJpja1Yh0nvOXHUa8u6yljfRnkKJEMVWRGF/M
OardAh8Vzq4dL/41nWNU1mGfBtau9LshoJjtY4qE6yDqiif8wTAj/2R526Os
9Km5HSMIADppy9sw91VOy2zaXgQFIm3BKQtorc6fIi6fz8GerZlvysx158wh
Py5nZcn6JtxQbCWAJPojDSe5nvKEfFcllcA33vTXSkqv0Hkv6u4KW3GjAbV8
VeS+0wnqpMvCDwvncDI/gYat7Fx20O9UiUlb4f/MilmAKxIEANXdF3VRw1Vt
OWleYhZX+XApwZuD5o5Lm2uV5IYPMCZmraDfxemurGIPg+2eypM5AUkWkYvC
H8gxy36xgnncI4qPIyXRnN/6asnrTTyHgRzxqLyIiCofgEmwY9cLSqIOEZew
hMWAuZ5Hsqey4PivC5K0G881SSOUBiUwNY+3LgpqLAvEkTZEdUsp/vQv/J9f
bcpSyE1iyXrtaJHII9r1GwTEF+DvJq9gE6Zv1WGYq3xJYI8YcD6+nKcsosW7
HqNikPqXPUq9P2/L4Up2zIoG7+Hn4OUSGRN80FGZaA1Z+5mcGmqAbstnzbMW
o2TWtClvspvxV1bktoD4KDtT6C6ldrItjtsmz+zbMh8yCL+PISC8H0ubajQo
qZfuCdm6nqoC+4KzAXpirA+SCaszSWSfSDa59AtxDL/2Jte70QhQHL6aIB9Q
qGP3+kte87p2+upmCeiTazfUnysl/ailzcPV9VTlClGzKukg0SOxKV+74kdv
yyJWUpU8tZVSmlnn+lg3yWu2oiaSRnwQpjlWzZS/esvZmo2Ynv/8FZjRkqqG
+c3pYlrfF5dz25lzxiEZTpyPZ/RiFdSABmWtDlWwD5Oo3I5LmTmZ1hyAcnmo
neRyDatnuyB3reoo5PXfTM1yVXJOl6VXmZSLHNtj0nYM/j0cOK4MAhd3OQr5
CCyYmB15rQjlkrstj0gjjbF9zI2Vh8ie+yb38OV5Gpgme5UAvz90OL4+i2tK
WlTIbX138mtYlYtbfNwXX7EB7oCHa182s52vC0nnhN+/71mCWN4OqT2j854o
/BbcRzDAEVb3UCKsNeRhYuxUS0PRwTZhM+Z3me747/XiavF/bJUjQFmplpRL
qh4CIfRqE8/nUDQRJSDunxB0bk/xCPxmg68CG8fYIyGkB+SBxCHWec7rlRnL
mhbj2Ax5E5fHhXR8+kxuEI4NnPsE72tXorw0b2+Cr3UuJIVa7LK1VbwUUl2Q
k2/PoCRo4W/270v9/n9j1oRifelvsutHzrccME4JDJz2Cgfcp8T0J9KXBYLg
bcq8paqWlcs13n8sstX1v8Y5SDEPCEIyoXhfUaTdIkMXR1RA98u++F0xRmm6
BAnWqZehWqhKL9j5M1JxD3nEprmqQquPEVMTnCIHTsogA8qHus75+7TElEyE
Yp9986MAn6MU3+ceVW3pZ+bDIonhC2z8o7N2K1kS/3+9shkoZuruYbmWhdZv
geznLPwv6CMovB6yXKVJzltqWXjG5WrfBC+3ETANlL3Vuj0AIu4n12yZV7xD
DiD3B/i/G3poXnvyatmBs9XHH7dRhewb0Wwm/JQeEXHMUqJsbBWjlfp4zBzt
Px5x/4jjvoTqSapDCAoUrJWCC0llncMScTpMtacJWRJ3Yi2pkjNo679sVrXv
Kt1QnCwFOtZgJ7E4k2rlpwWFmBasR2tPTCUx3nKkDNZryyptx7NvSgZ0d3cN
cpVwWX9CeYfG1ntpZvcj0skYOMJY28E+gnxkcbhyzDClM6MKA1ych3ag2Dcz
RBR6/+/8v+mCZM1dzvziv2vu4H781gGaz5XK8cWiMeySFtmkKM/HArLvSudR
fnPMpmfWc/tfGVcz84LIeEtEyLzOq4FRTm/2Cw28bUO5m/dxCzUEteJ160hR
ApVJTLSthWc3vMN0WbPhhwGkfzDHx5mDpa/6IFw1tpEP0ZsKblgpwn57e3Fl
oVXrQjEPsMR+H+WcNZiDHqL+L6Ila65uOpSF9WHHhJtqQZTrCQyH5HL0q0oK
409y1Yq12EAPquuWaR8SL9qAmCsslH+r78Am6uyX/FNJeBX7kabH/bMuSplG
UL7YYmCcwqrshmIg/G97+7ilSZ2jfk+u2lOQeDCXDfziIc/fOzYdrw5htWFR
9hHEJX7K5dTPqFN8544wiCNj0Y6utkxlv1Y8QYVPSKtnUx9c0ab5K2Eroo86
5EzTDs+Ml8X5co8W0gfjIfcqjUmScp01E3KGF61krVWNS0xJBKRk5cOxS06R
G+tcgULn3F9LIzF7ZzRohLQ12ACqKhwko0Ubn06qjmjIkSUDHcPmUU6uEJie
8u5VA8iODkVvgGGqyWPkqyBl1W20STeRBe1fhdz3OvSGPz/cPiGWDMutugwc
bBP+6PwNFZr3RX1qchuZchlZl7+pGipr2YvdbwZ3hcjfHoCDKSb4NmF9SZ/d
1eNgP8fI9fGu6y/rRbuflaErkSZq9NxPo96gjPYN5rcFH1kHHs1talK40IT7
3amXpblBNXpd++glbYDItgHCxB+9mmcHjpenK5XNtKTicKQRdbgEhK7Bhnbx
nj5B/0wfBigWkoN3hmFp44V7sLxDhtLgU6etChWK651dgf1qdgFaByZFNiXM
SmWHpMKe+hhtww8b1G5fmfXI6CE3QiaaywG+OBSNWNAjnW6c1V2Bu7Xa6/qZ
dfr66QHNCqa0jMRNBdnqtMFDG/YocOixCKh190Xh446TXyaMFJCokXTajNC5
tRUCq7BNYZ1NPh/AYlZV6KkKDw1I3g2z/ge25cif0VLC8mC1/J1gBGDSA0/u
isc6d3u+SrvoKwtLkhY8ch5O4bxEmIt4Hfa4kVQwXqt66+2NnLu+N8HF/0/s
CTMu00t3n5V5/pVGDWATKOQ9uXkGUm3Ql8EFJXjg0Ey7n5XeF8OfrtgIcYZq
O7FpNEN4tc8p1hcKrJFKNSINtRKRdFVBKZLL1dxLZmQyAKwSvfSJ6M4QxIXX
Y+Un8vuHkU6RBmVE3aCHCOukO+NxGfrXC8LEOrWBUvgGNaHLGcRzPBYPCBCv
nuJaKb+8wZVmmrp4ica/Yuxmtqb11ENFBZ9jPIYMjMdBj6gUj+g5vdgN/Q9+
8M6J+lpC1MTrCGiuRZSYHVnuwVHQ/URB9oGALk2w8hCimU5R3SBqRnQ68pZa
hCFR7momdpBgXq1t0HFG47kfKTAWE2HDYAv+1MOs7MfaS69p4phbxmIhzuNK
8uER4W9IPmIMQG/KsYHTfkLBwT2Kw+R661CTh+qDgWGUhltCfnad5GwinuaH
vHuRys3AzHRsPQSzd15zmi6nSZ2V9Qb8mD/Cagd2r4c2gHI3t3n0FfFGLb1b
0T98elWTX2oDkVD6/9BVUtUHKOQBjivKpVt6MgFaCij3SmHq8fCUAzc/O3O0
m9iJ/UmiBxM7N0wsSbTNe3vtm2LX2zRHGaS0tCYpVhVf9D7wsrbXkZ07M6Z5
LlNr2+wIgxcW6JMAvDcOR2xAkgquTiFHsnKZASALCX4feS38FRev3cvba8Nk
Z8+hAQPkSc60uAKU9IBYO1ajaua3ySMPm0A5oZQLyY0YEyDmXEI559E+8oe7
9CrzbnFXfqje0V7p6LzMJcsWlfYVfA9pqhfii2lNVmygfSNz0ZfYCXaAxwBI
kk1hm5jx0tjPyxbG4qT7lILMhplodCk1LzKfVYQmzw+5Pqi0x8R51ca0ZUwz
4kueRvoEVFxEfnj12Q0UbSZFws+UpST0E+kgzb+OUn5jzdji8hTDmmpJuTZY
yGOGUBYBRzzYMxSWZhtJZIc2ByMKW9hONhxkuidpMc4XTSNQFx3QMqfRKQGb
EBSwkWxNayFEKaZgD7lUl+4KPzB0GQmD5qxECbJabVqC4s512/dDpc3pkUrS
a42HAs40YD9UocTFWY8t+cXrI1FkXE8CvYKflFSqzMizNHz+9xDZjh8tSJ4d
wg2s+9GCSNBzg4/+O+/WDUy5Tue28gMTcjkV5w+Sqf1K4HMTwQ0Sa9quZJ0N
6+GhwgkkyJJbR5wujg2Q3fxe4pVVQ5dHjQKfHV2fmxRcNSERwwtMixGjJDAn
dVcWiFo7F9Br5IKIRdaA+pkM+/7iT/4OvfqnlY49yyw6GG3SLHJff6W3Mzea
uq8qrBdoZ344QxcNvbMUNBxx+1c4QLKhVymZmasT48abI5IOlJeDAvOP/bXj
gviOOAGUtNMt99hK00WFoZS8pGrCjvfGrZv1QknwZKVPbUkp4ODmycyIoMnr
70wSrtgBkj04mQP7cZpyvfdFW0314W2FCzJr7NdxtL/9+rv0HbAH9M7QjBEX
JazEsdlwxCMVUEuPjUWUHV2m8PcmeG5xHOnDULEKzkcK2WwbtixelVaPmXYM
fkX1JSXna/86ThA0QnKq+zibRecUxOCA/o+fyNcnywuvV7VlIozJLsZiwvhj
WixKMY8NaXAjeo5pGvtWxrZTZdmGcpVHCZiE4rVUc2DJx1QfleyeeXJ73qaL
gclp5PcZIxu59c2vESgLFOLT1c58pcA1GdyKpqMibyrUv4sP9YwRlWpIZJaf
kMbBd2R6bXHjcDVQJVyrfzoWMu9X5Og1EmYqyG+KGeVIYOyXo5PDuhIMl/UC
OKrMzvUCMoaZu7/NrbIw+QDQ1aB/rEPiNrJ9WUB6kVuXhQY4fTCHqxtuyTr/
oerwloxXoSEhdTl1SjKdiEiQetrw1plAbInJ80AosffyR4CnvTsxd6WYLd3P
/W2rGlVHXfmrxsPN/WNQy+QtQwWC1V+DR3tkJxKypzlRgfPi+jpvybBf3BAQ
M9G1MaVEd9sHp8l+Suymhc7eYFpii67eheuyhLuXXHs40W8ZKvwK2ljt3PVm
rpM8umT39h53hZ4IH8n7yH3+ezBbP8e17hTMSQPPeK1Sk2rgtLRDbPXMcrpx
RLjdXuhggnRe9KVK9TjxLKy84eC1arg0tW3Lkz0HIBkWFcMf025J2LxEozWv
JrFujwgMxI80FNkoMED2gUGQFRsmBDY2tdpH1syeGMktsqj6KpfvrTTpeHHu
ZRyKjJWDKDpNwur5JvPho5deZ2CM6UgaW7t8NsaSMagwClx9YPGgQFV/vux/
VOZoVh15xns7Lu77tjAJnien8GGHg6VMiT9H2wDWXqSxF/oWTVXaXyp3VcGa
OWuTag8dqa2cknpJipwQsV0CF0k6Y9ZigQAnGude3jl7N5JlC6geE/XLUnL0
t+pGOJJ29h8FrxHkuYR2zafuDmyiV1LQ1F+U+4U+WgVs3QBa674inaubDSB/
o4pVyFbOTXUJPPSGAkw/zqDIZI7dycgDW9fPJJHFVy6kKefr1Y4kg1HzgT94
pukYina5/dXb9Pki8Q6d5tOpPJxdIm9HHOnyEuDM2LgYehDBNjLZAQQqIRft
Yhgnh5Tgk/UeJI3MCMahlouSvkR0tGEWmugc7ZAukVGPMxYoWnRRKWZPaZao
M4Tv1HrkiEElDmXby0IhBnPoIJBXPFA5dQ2ME9HHgR2+Mb5E+83muYcPa4pP
taxNQz2cGIQCTDWwrL0BDY5x56Os18IjrZifz1to1Z7Pf4WB0MnTkpWRhm/0
9gXeXYRcH044iySYWP7KljU5EtaBF0nroHeK8nEcQGlEfcQhxcfIjrS3jXl7
sFaEQBq6TxeYKhg2ncBE6Tbp8VOM397Pp43B92nNfXN1GnJV2J9Cg13JC/Jj
gvKd8A1mNoao6OGdMPzJAuXC2vZ57lxVmwlkFhymriuhGvWDYcLUFR59dd3u
WKNyt675BXfqNQJ4y8Y/1GHJdtZOuLz0hCpok7HsH9fZyEU1IKNIzq9EyEbh
8+T0Zw/PErsuI3PedmRq0TwXCZT8GiK4Y4uZjHb8zlQSDI9XutXaHp9nnOh7
8iHGpQ/qhs6YGfKImPvz7mQBJzgEm9amIxOTpAe95VQeHq3iRGmzwh9W/jXe
b/b4I+P7kJ2QqKdGuuAMZf4KM4Aj7gaaOoEFd1VITBf4LNPXAEGZ+tjghDip
4KGuv5vtREUN5iqIb6uWh9ccrJKr06ALHxuTxD7hqMKki/ck1mNYlXGXD5oL
AjJru1bNpjZG9eTXLcuCyaYlGqoreBt+SRZmPaQIpAGWANwEOSnOfG/2ewO8
VvmrhUZerMKFLMJkDXAbwvOF+ccm/jE7cfm900ZISmW/4Gx9vCtzKIpzspIm
w+lnxEWpaNLB1B4SDOys5jILx6RtS94iaB6PgEi2Cf9toBMgG5rs53bdZyba
r8L5yOED8Wq/a+sl2FE8H2Yy4LcZIWvxF2KHk7haLeFi5MQ+GNMZreusozPS
61mpALmui5xeSJaF2W3bTQk4nkpD35UCNpqOa+TGKsSk1EH2k3ka8FHLmowO
g+MZR3wQ8S/BBeIGQWXht7jeEQXdWtw5t5Z16AGvNfiRHAz9CWbknCJCDDVy
rDQjrbkJfx9tvlUPOtwrR5UuoP55BP+2SjpppblvyQHIko8RTELJbw4tnIwE
XqiOOLUHL0AR9kraEpzvS51q1RKsbnQSCnLNNhozFwkQP7HpzCKBvFX9YJk1
AZ+Sbz+AgSWNSoKiHnSJKRMRLtfnDN9cPwiaeBQV19GDDMLomlyHgS0wfZoi
YqbQ3dTuq/rXNDK3p6jznH9+0Rnt7pEI2tS94uGFB8k6RAspaTV1lVjMzfuj
6dOpdUdO5cWDy5kzonKabr49+LXklaTKiHhGKpCD2e2/YaBPS5NfH3jQbG/W
cyBzEAMY5kNSGu+KoOR/Js5gQl0hk5L9m3yTd8wN2e03bB2glMGCUbhgZgNr
zja8lV/id3cp2UsQr7Eeb3VKPPl5MEAsHkI4ewBHKSVhXO/HCU/vXiSiX04I
/JMzkkriOA435cth3AYjpusim6kTUwBBvz+7RNfHVoPRkLOYWtM4s9WowiWk
DF0Mpry1TtN5LHYWl6Kujv+2wX4bQWUFPfzVk74pG7Ocpk7H8Vn7AaYg27DE
a1Cg6ZiFe/DX72pLImBWmTg74evteBAUWJ4BwiYRWD9XmX7K4dFbOhAviPD2
04JDpOK6n0OypfqLeWKxtXtnOYHXBJpRwHNJCGCgAL5Oo1kd9R2z4J/BDex7
sXTNOxf/t9SGi1J583/Y/EKdSGXDCYs1KyvhxvJitzFmTOOjabw7Tv7g9+p7
z2dPoPUVBXmkbbmlQTcM5JPfRaYZWQRph6dhfvvwIOgr/+AnFWZi8rvxm9rs
5zypCf2bqEFmgN+7g0gM5JuDI/86dJDGRF7s9fO1XJyDeiBTuA7lXBCYIDT4
d0XDgfG2T2Sb/kZBoN7yM171aG05oNXoYwCjsDEkhYd/b+NJFgr0JO6aeRUy
2sBZK3n/UIe+nrPlcwEFmBe+QHmTc351agUAi30prUaBlTPYCo6psKNNcg+4
+5A54sCODpTiG07osqkF7PwTC7lIVoQ3T9oALw26/OBX4wbaEis5ufgicKIq
+mxJbCtAfrrNy/DgwM9+fwHHyr7dhEYlLSpj3qgHavzAs4zNQEOeZn5glmUy
KZoQCu/vzzyXOdwlyjJpvPhVighumRfrPHZXnfwg89jJkvQ6F7v0XNhZjuOR
2bAdOBsux3ef9a9V1uDb3f+G/TduQMd4+Eh0+07yHUUcnVTjelNl3vkeV3/c
NClPCWwYBxUvZ94BbgaZ67FwDvYAuJhlWmx3cdMd5x3tbcn+wAss2jfpe813
5wfjJzfNR3zJV4WSThkHjJGL3ImFc2xXzb7dVXwMSsaicECXRP1NU7LNc5un
dCvLa0Nsh5a54rrRDlPiQzLHOZ+9g028VhwUkvoO9JBVRmZYGFjBfreR4eUf
NYUIYBOgo8SvlOggrJmrP6vdkrnvZT/uizHV/GsnS7l7USvMYLKONh0nTWmx
wHk060sSKkdKNh0VePyPdUxUbB45sQFsGmwtM1Xakagorv9d5Ia31F512/4U
gsIuIKFD3mOE0wD1V3gCh8nF5e1JieXFSVY+U9/CFTnpjgTOIgynL5G2hmeF
tphbh4hI2ObGlLQsmHXR9gJwLmhd0qBBHaKcv9q/6iBpPZbSMZY3l3b2h2RA
oShx08+0PWCjxfSgC2aJ2kbks19q1qi+d4jdhx2IAzMKB9W+Rh8BoTz6qDBI
RwiMbLXPCBPoN0Ye1J2PmhWwB9aG0qKWBH6vj4MeWtN8M7jLRVqWUk03bgxX
6/1fGVkph6zsFdSvf4cXIgbXV7wA3BPHqFE+16Wq6+qLzAaScC0VuZw3oSL5
E82IqKtY305UGCmjpqQQoJAchSf5b4C3j08gLvNGPKMMNrHi+I7jtncsDUIj
F0JHLp+iH1u4j1wOF6xbbpJ+TIngZlHrZ8O4stm/NDrZ34xPnpuZfAV5LoRs
C0suX2ATGrzd+KStUV8SvAse2hIVL1Zu5m1KotW4kQZ7X2xMQuFTmAL0zGUl
PZvOG8SnPDtluPR2J/ru/2FNclVbfhp+xjQib6Z5OJ6rDONk8iL6CdwPprWL
4q9rgw+OvDRq+3BVr8mjQBBYUEY08Y6C0Camos61onV2gEDkueZjXdTHrm01
C2Qii8PNKWF0Ua62DBNufKSb+H7SV1xPKb2ATbK30PIHKLfiyuDM+KU/ukyf
d+BN4o7V3Or2H7jZpmPlOonIKiXqLPpsUFbt0Q9qu65tRZ2YTjQx8H233eDE
pdq4ktm63dNouS5zAvf+lutf89y1CiSb0oylE45kXqig28OoeGTnSavQ0SJh
0o926kaGxK6A2MMzHGRS4xLpIdaMaN6rSIukPxqvWTlg4DNmDMxrd7ARm9mV
TejkTuR5/DX8DKBPZJ0U30nNBzi8RTeyST/z4ML1rjf5Iqhg9B2eoIn4WW/0
ZaaZhTjD7AH/zrvdVKt+1Bj4HTgtqvnERO4rmNlrOYnhDtk++j0U3Xa5OnLQ
Lvr2g6I7TFS7RvR4eG/MyGaIwVHNKzn40wQKWI6ur7zBxt+6EbEsUK0TvdLT
o32qwe2OwW8xt2V975oEN6i220H/By159uViZ07sYxy3dLZ2HQ4LtpAvkgJ0
0QXU0mS2Dd2p7kIpDMbBi3DdLfxN4uzJoKxPV2NwbbqwNkXu3dVrUBlG5nzu
W0Prkliu/hlQP+WgM8hob+aDEi41/vDbDyTX4c0R47k8mIe9+FKupedxMf5G
Gqmf9flhgIxoVX5wqy5L6dX2JVmAiz1CdqItZuBTmAUAU45cPUdMKnvxc8J9
+Tm/W6wQzW+erRyS/4q56j+K+id0Jwrn0RixV2S2lv3J2yqZNPedeMQE20KR
J8GBZ8+waFmsWewDb2bECu4WLUL3IJXo4iild+KOzx1FLmR7TCbdg99fgl/f
SAYvmAIQ5BV4I2d3ZzsmstvooAcMGZJD3nruXWMw+3q1BCaAS2davbfWHahR
HPoCzNcnZDp8FZ9sH3kBoYmAcW5zUx7cV+PoDLLsRKGisod0vrd8np38P2tr
x0KtHb+eGnCozcx+Z0bJ9X5YkFGY0Mbti2jQyx/DTiapNg5+8KJQzsn7m2mh
7k/f4saUe6W08ZbZQooVzkjUhUxGZReP43ytvEgWaLUDCE2MOf7iF+i1NATy
QKWfzWcQBtE17Ipx9DJXhwjDbvf9kIfFNoobUWnW8TAzU1LYiaCLzfi/kiy1
tBfaqCqLQRr5DAqk01xzPS0rXNj29E9gFDzxygVrdqnT6EAwvdOsEq4my5N5
Efi9KhRRzgbpCA2UVQ6s+t1HbO69iNBw/g4GHsB6vnHFg5UlzZnASHTMmsjp
fZzBiCENcWcobJFUIjnve1lJZcnjhBIlAo06ETFxJkriRPohsKO3LTB2OQtT
9FbkjPAjrEBV1s5buPJ07XxomRfE6fGoFrgG9yyLq1h2vAj/3jUB8aScu+r/
dNmAey9ROCN9XOVwDlngsJGnGJwN31qnlgGDO/G8tSaxrti/EBrHc/oZ6pI/
sPtcpNYVT2slLsAZyFhm1vfanIC+EdS7W9s9V7zEteJ//Ak5AJcMbPY7CAER
aaTd4c0eK3O4ke3T82UBmYmIeD3imh03CLL7vdb2M2hH6iIi9ERIdi4RKGRE
rkHMD5DBtU0GbK6fWZvBmuGU0LOu4IxGbJxrrY+MnIKmDATvdrO/xaMALqYI
bh4bggypcI1CN6AiDn4lfpUQBxDiQQ0hU+/kkUvg7Nt5okHJw1ijvT5mb5OJ
e282uPmRqs8z82ljStaE4j5ZYR7vs5If33bhx667ErC+j+sQz+NUvI3QRC20
ogxw4ZbQKF4TXyS2PPlnDq8I1VljJf3BacJFszFTep8s363XOIcbz5FFPDHs
BYu4aoYblYi8IKFKUL9d1JvSZD4nE8VLQvmFcApMqNM4gyDzNNZL2tm3n3AR
TI56YQRywkncaAClaHKe5BH3bij6rDFf7MiJWpfbodTnv+GGS2b+BYRXrOVR
BRbbqeYlOHzpzljOkh9xJ5VwCUd9m6JTs6ga+30m0J8nOLnjFskEcgdJtuEw
rrMSoRF7WqqITnq+5+tnAFrBUu5K0Slk7E7s3bLVD0o4rlRxsIyY9Oie92qN
QgFrCP2RhIRlTrKOBLuMjWiLCMp6o8qgZUD3QuAAneSGkOpDdcMKtMw6AHHx
k4cW00DLxl0Eit1XuD+z9Of2+Yz/i08+hVSEnEbnpRoAnWn3NaQwbD8cB+w9
MXPZU8Kf9HDi5So7SoKbLUw2GpC1FqBi9PmpltKRu4OlHXphY3+CJrxo3/yT
wAEGRkNZi4rZGpZsSdu1O0N54Mx4wt/qbbLz0tGdsalaPZ5oDmtabIMtt1lO
QiG9hz6tm0fRy7YhY5+JEbBj6Ww+cotQkyqsTPR5k799i+3ZG+4xHuTswsLt
+yHfQVUjPEpeADKI0xWDobloj9l3Rd0sVcK4WUdmt3d9xzb+cKVqm9fKDBNl
QU0dA4ifX25u+TWNVU0kji/4V232yJhXUChvm3iF/BXj6x19NQXlv9OCL8wO
5EeQait3yXCRMjE1/XumurUPpOEcpatJIHdzty9WQx+DVocyGIBHWWAz4xuK
NJtlV4S74rTVMoluulnumIwvvtw/2xhWjamUDVZMvrwFgIyCAQAYbqe1dz+V
BcWFQJlvoo7SRlTbml4DcP1LSW1+/cUDgaG0SAXuz8sRiUQT3sE5LOnwzGBz
3Z2/RkBVHm0GdjO36mPI8gJbYpSIQIunrGX607tw8sxvliCGuppIjezp91W3
4plEqs7k11cngRaJZ9NW9X+Aqh2b7bbpxOYSewSXngLgoM5PnYwQV7kyI8MK
tGSsi9jzrobLp1ljR4joOp+88CJWcy2T1riyo7fiyFx7HTMNBxswehVQ99fT
4VZ2g/nFthwTlqUJpUETBznfIkW3lo394w92Jo5x+24Sjc+0Vvob9iuw67Wu
zEWx0h2m3Ojp27clX7a8E4TfqHj53/da3k/HeHbKltj2ROVqEG/iaXrpI7tg
BFV2G8G9yXX+tl6z3N5nI59XWpX4ctOp7NCmiv4oz9+kRMCr1YeFvacKohFM
enY4CyDhrVuKJleH7yVnQmB0z+w61VnSUn56r7qTjjKCwosrS23LTxkYERCx
b6EU+nrpDrztu0POt3kueo5tSYanrPWK2Uz66mWnM900yKNc0HfQdBSOqnXv
3CMBBlhrYLR6Ii2DgVC99CocgZiViM44PsEAXl1gxuIIGsQhgXm5CIZnLbyz
dDwVjDS+Z6S6TfU6FJMk9BqDx/TqfZ6FFZA2+QxfAewEc/yGQydRFV0mKEps
SahwRZgGWT4bLvlyizmR/z/BRCqwVlEYpl1JImTxQFkiM9rSc2fY5y+8NX79
GhiiT4Hu0dnASGkS7cURhtYwDhmcNOXnKkhCDDPd6+GGhVabAawgka4OLp9+
WewiB3XvsvHOUMX/8wVDg/yLhN62KwrELDE+pmNFfS/cJQG6fNnXgjO8RTKM
V46BFBOyrZ04AFcXBHotayDALen9iRkS6+nh3V7UQypXk/TdkxgvPCMmjjSh
4j0pBwLqH71BsJawetljdCcScb7M2gnpm3GQs57TdvBKiBjHAD3Uoeq5K8BV
YD7AZAce5e73aTcr2mYNl3Wr0OxX2WbRPmXCnKj7PI+7cLVD0cJPXyoX3msv
JO40TUX/4DXkuQIIR0tiKxcIF6bcUHRdpqQzxI2jenMnlLdFe+AWegfvoicI
04QOwNnaihrQ9FWlHsSa8yFFEypxKQEGlDFrhGb09nFk0PHOXipBvUOF6MH7
kEkZF+h2KcOf9eiSxMW8afZIxnvJAo2JeEdknbPPRCgyRJCbvOk32MFXqNzp
UWU+vqatxxJuuXISxBNulNAwbNJkb02uOk2o0EvSOk6wG1o85/+HSw1DNYPz
8Rt8apiXMvnORjBdJrSp2niR3bNHKrloLNtoIKQTco3K9AHkfmDSYPpC4nLI
4UboRNNIlJvm6dbMdea5h+STJY2f7hsuVA84vTEEO65DSX/vs5bcan/MOqzt
bg12RBU4Uxb+piVj4Wn/uXKB5KC+o0Pc5zvRMjybLiFHeBoH4G2KnBp/kzVz
F0so4KAhlUDDDb71Qt8I9R8BafMXSC3i0Czlq2xaMqgO1Varsggb4tnVVsjG
zG9QQ2eZs5gH3wbhZecTAqMayK82kzlYz/O+X/aRh8VPtucqCWMpYAwH9L4f
mHSFqHC/LIDzAcAWlfxDrtjcV4ObzTPL89Dd3GbIGyRf722Rr9CAdqjXGTd8
aWEmcz2ftqqQHozYzmJwzIdgraOxYA2AK4ufDnTiV2UgZD3fPsCmZoUaiEVn
f1dNPLMVltvF9N2cpOXA3R3490/xW4WK9q0iYOb+4BWi7n5EIxORsmmPS3eQ
Z9eaZKy+sRcBDuDhXR6glnlg98G1qHH1zUkLARoQZuOxnrHw2hr54jWULM8J
ruBx1gUB6Bb7uiHASJXKnipK2FZ4dxOfKTwJOdjhDS0CFSmkGK8bD0PlS05N
EJuNUATZZrk1z9ZtKEEctYOcuIDoZOUvxIs5Qva6ztKaC/PdrbzCb7gze3Nw
4SEfcpXlCGGs2IvrL1h+edBu18Mx9s06d76tOztQTkqv8q1L79BWk6kGTIdB
KR+a2CyFhXYlb+cmQlyMglXG/zviKocEgSWPVmb58zLL5RmbNrhOzYqBORcC
lNVeK/vXlX/oknko9F3OxSHevJX14ra0ZAe6aJ0VwlWrPJhaZwJnmxqnM/e6
wSSoDf/B43f7DF1p9vvci7o1k9hiZYdwt3sTNFHwJ53HBfOAIeNqlS7tI0xq
+LRuPLhekkRsBYelVL8h2PWlO9MxpGxeU+V2lrnvB8ZHOwsj8kx3Kda0iP3v
NoI+0Za2HGgmGDqN+pYFGCmiIZ5Bn35YGlcmhYgiqQDMNSZIQxXgpdUGQjS4
AbnTGsdw+K0qcXmKtpXVv7hR+LP5mfnFHD4lDgREY/KjK3jKhVJ84Xs4AxmJ
416U2CFGjyUe9UuyH73GU12hxAUmGEL0QtcaK/wnO1bBVMotm1P70l4PIO/K
2NDTTf1cox89bmCrrU3VyzEYL19ekNogb7DtwRic88Z7rKeKqHK996bKkHVC
5OgsEMc/G4Ain2HOP+5vrU/Do6mzFHOMA2kJGVrUoKoC+Uu7njQhriCUJan2
uYy36Iyo5vhtTGIW8CRLlnZCPH0P95lo6VRrmG9qr0csgrfl8JKrIwZIRrTZ
qtLKljBS5AIR/SRIv1ODcfXq5Z05hc4UsYayTrZ1x3G/uT52hbsTUH82a027
2jxezb5pYSniObGn7D3H4sCQMY7JVnD0gCS6CK6fmKg/+C1TH2Ozxu0jdtON
iBatvmqyV/KCoCW6h+b2GtSYjaZ3JZh6XyGYwR0MMaPaIx8mvpcKzPvcdHRv
PHWcarb3WfVVWkIdnRqTxgZmqjW2XHf2CLykRnljeHH5+i6i+JKCqgRYHg6r
oGhD5wnGPcr35ajvb28aYcpQBk9Tdk1jTEDQXo2ROA/dTGkiDv25Ni3v0hwd
lO0oqI4chuNhGGSrsGrKXpeJxiesDt7rvtDJkxUBedtQ0nr95RtjnqNqaJRw
60KFm/rpJ7nkKvBuRm0bR330IFOSdLVCDFQC4QYuudYZX+glArCKj7yORRzU
QyGmjyvUcsUVIAk+qeDM7GIDfUYNxtLF9tVzorHFN5xGa1VfjomOF9zpWH1p
GEJ+o6qncwJm43iVxxJS+jXvKdv7HEnWFfEDXkSZVFByaC8SmI88tKCd4rL0
csiaFrM0rHql2qFojrsgEV0wAoxzrZbn+TwJue+nZFYa6a+GF67n6zH2sYZm
O67aJC0yMAaJg4FmkLndnMIdwn2HTVE9qwpPYf5o6nGjGTFeT0s3UWUcAa3g
7frXMY32bdSwOgzIFDsI5g8DSyNSYGckWGBJNXmueSDDX5OivrH1yurpxzDX
0HxXhRmXF9Z3sQ+K3EBDZ+zXClos3eQmBtIScdQ2lZr0HI5T5o75Otq3hMhY
0rXxHxdXPkbucua0DbyMRpPsn8eWgjh8OYgKUaYMDpbhGbOb0uvHF5jbaTB3
LEXbjGTP/bzsDzaSMkxSNtwFBAXwGmv3FFGEj/sXj73ySB2Z4X3zWkO2JG7w
wavokbZUAj+3UEa/Hgf7WoxMrn/3NHIwYHA/Die+3kGLwHW1g/a10KY9rsKY
CzWqS6emAMqag3UEknje/j8xFVbiWWoyu5CDlHKGKRJKA5iiPzYawq0IB4bE
4meALYHFFH5K3Y7G6q/lGI/ogK2Ig3KYPyCeun/Vy4ru1BQzIWFdg9Jerice
U+ykfyOkwGMAkIwOovsuwVjIzCsD0jSQipsMhuQkefBUA7g8VD3Lm6fLQ6Ju
PMP7HSQJICMkpZTMn/PmioqlXaM5rLrREhPJDt0QL+s6xODIj/nYct0MsEvJ
hWWX+6EZadx5LSrYzToUJBiEHBj2d8hCl3fzF7FrPfRaVWtQET/hO5Aawy3a
BDIynX1KtUzMMqLclw6m/oOcv7PYfjx2h1eDPRzuLbOldZgBLtKA92+wxgWa
R/c26hLZ+P2C6/TDxasFyML/XrIbWJgfTX2IlAk7a0tn0tF/6nGbcHU1k6QD
DAN2o4Wv81GwWi6J0AAAmFuj7ZnZbpwpboTUBHsDTh8Og5SxGswLxJkhHkHt
qC4K06aujO/A3jhNMhaVNLph4BIZQvwLfgkdXuNimBfilGtsLzvKFvV21EJT
YQWYhJIO3XH/yGJcC0MSfboIG1/cmuBAU2OAhUvd4dbb/b8p9PQm2VQNDlHW
5GhR2EC7XP9qZUyEk2gaWobx6fYAILZ21EGFr1uUirL5qKeXOlbm3PUu3aip
7qT2hi+uxIqrAaqlvM4+FAmmZEyUWQxDRsAM7VkcRaIasg6Kpz3vxcAZt4sw
gKLNmNaS/zeUViHEpB0ritXYIvc4PxlYaHBUc8fTdxtXiFDF1KX/nlrwYFNC
hX9v+csNveRHLmxghT3h29jFEN1WRAg0Cl8LDLoH+PZ2DLIr3kq3kn24znTc
5OI9lN9ahQ2j3Ax9CWxCnAkG8YOzK9LmD9GC11fTnoSUThV3kN0uMPxl37dk
2EsJ44AEMqVFPipS/IEq6qO6WCaB8pMk7yxTgIK45XXV16gNbFCNPmFHbBag
e9X0bhz8YWqrcmCQqDr1dE0MCOYrN8fbgcbQ2LXX9w/9akotwErtzW7kKD0A
2Ekn1P76oMmvu5TO4kDK+Y5x+zcibB58GiaG/Os0az8iitAAaXsQAHzsSxtd
bdQuphTFjPqJdluaSNuZq+nLHuygJpDZHN3eC+Rft+o8BhcBv/vLrWcCifEG
zEFNB8va3BM3/s1KGeErwALekXbMZvoziAnJrWjZSssUeYEo2N1qazWAcdKz
tVOyW6MpyoNygXkWirDB/gVX3aMptvVqdwnxNzrxJO5Hm5bORrT1/7UZlTqg
yEK72EqgDhzrIW6yjJsGMds0fCWYYEClZMSDekDvqgbBs7omGIZuXluHYMYE
degIvkCw/gSN/24JwCKaUbR73lGYx8IXSWxrTfmWywbaZMohgQLhcGBBcZn2
Z9JntgH3LdK1BBd0a7hO2b2maEkVYnDDjQxI8ClCtCs+QzGgA2Xx0oN/qriI
G4rxmwQe1SzlHXGOtG9pZzE1PCdn2sVrEjCP5tfdlmVFLg/EYGWykQw+OdX5
EuQq9CM6nvle9ExbyO6of3wCpXETDa9uZcYkzNJDIhl7hwzvlHTGv7KthLbg
ADIMRsOQBJsB229Ri2QdDwTLcP3heA71VFoOfVqEhdYNotdy064gZtMWsnoQ
C33Pne1a7UNxKjcITfral3KmByd8Hag87hiVIOG8Lb0v6/Qx+eDE6jM7n9EW
B1FD9T9EU/rAIPEwlakXPu+NUvd6+Q1ID/LtzhkKP0i0/Cx+bamxDl5NdiPn
5MLecupa0/xxuNoq7g4Sr9psUeQKnhtU3O5QIk3AEyOo6u1yBLkLRdUulhzU
hdS25p1UUOv+wsd07kT3AahaMcywBP8PD4SG3useUHPlhFdFEh7dtRXFLgD8
KyrzTYBXmdvBOq+wQhcVsjDOgqgkbLv63T3zHahDfossC9cNd6bUGpPpgH9T
p/VumzvfS/owqgJ0BHp2G0jD7JpLBaSTotNNLU0S7/9Zgme0Ufb1g9quGsMt
T5YRcWGuNiw/5Ox3OEote3wXlN1Onhcf41mBSZEEv0or9KkLnFrZ/lGUfvHt
ZwrANRpemamNFQEPCZiMKlqnMpQfgo+q+X1TWnPIiRzva+WWdWFuBz6iCHrA
49VLvwr77wvH2OIJzsya9G18/iGRHfydfqo6lqaJu0wOsY5kVXjxOb/lhqX9
Jm2/bXsgM06Hqjd0OpTRmUc/RVB4yPHPqQNgMC5oEtRkU+FOrQqzL+dNIkEH
SrW6EVrCxnAbxB6rOJR45EcWZe64AcoqD8uPlR8taa17faH+fzqgn8RlX9qo
A5ZBFOIl6/W86FbsTLYpUE4BvCj5BPITkv5IjxAcXJHeVli4UEhGEJMmZ8Hx
+GCS6opzV1IrAf8Mt2YEcPxqAos4BaPfzIfEbGOS0Qn3zTKJdXmb3Mbf08jh
3SDgK1LvBYWR2pZccRewV2bcv7Q1Arj/KD9WpGe+xkRDSABxf5CAFXyUs5xk
fiFGttQ7+IGD3SO82DwjqGffJe/XmnvfhiafXVr7k78tC8uBe9Wp4X81dScA
dqLorZVncjGpi3wlJTRIwULYdP2htHX88GIsjpcW8Hydb3vHoqiJ+54QObAg
mVufmy6T8tIwENADoM8qI2vrQzMkLSshiy5hGzCZEDWBRwc78BnL+MLBULqE
m7gSjnbSy9lOZrkRfJojw33dvsnnlYvA902s4bzoRGiwtRWT43epNcvCZt4q
5AlObQtjMAAE1W8KXfmrE/SPwqe9BuBrwZGSyzefHLRtdxxdrEYNN1SDFLIK
F1SHZsnnfoy4ePFNcnHh+HmWn91ZxjSVRvsQlqkH8b8q4TO3S03rh6Gxx1mD
0TK5ytNRi1FLYM+lLyXEIWnbNT37e3zUQMajE+KXm5dSOIT8WlnsUqKTDT3K
s9Bhs4GW/ZM810dcdrrB2hh5M/4uPuVqL/5oigoIXSWFRrrBMqSOHcw/JCzO
o/Z/YdBk0Va1nPMvb1vV4uRHDd+QPLqGrltC7MKbJGxSzYNR3dIWBg1DRh0w
MJDsHH13MxMWy9+zDZdavDrMPhgCzXgQRoRnVihP4PlCAsenYKrnXmtOlZYS
heq+icLjXay29qvWOhyi3uGpYke2oQg5wQ1HJP9xDahoWM5cNezKXaX75EsW
89HX1hgWZGA+vj4tuW8XOCoC61/UmJFc2TK4BVc1Lk1M0b4rmX3ggkQB52Yc
Ej5iTgf1+drWRcj9+oN4jmubllnB6/lZ8mnoTKHQVUexW3ZFDdborCo5zciK
cpDl7mykLqaKzqo33FPNcFKAwvlXUl6sfnltLnbXIFfcXx9c9kMNmX/huEpL
gzFoyCDCGrv7cVnJ5C/s5Gppj/myZYvv2uUq2xjW8JkaPoodyR8ufSBs8Fqz
jfRiAGAv0fA3vN4IGV8qyAJ5rLHMUTFM+JA91sWEj9YSUZegBFXcYKdQlwJK
YMLUy+mEZPGJK1ZyfZ5WjCoI+6Y+mhJ4f1xEedgeBLYHQ7EorCiIOJmWv3xr
/aYeseFlB7g1MRw/jKrvutxmlfMc7afn+poWDRD3gaNVVpfTYf1aV6mg/ol3
O2+BGNzr4I6AXs8xIk3j0ciCsmoQmKCBm3MwKeT5IubW1y5Ezs5KM5FouRSk
SXrfmCoD9tIHpHDDVeJCk6wQd+EBUJO/r+Atfim+D+vQZcnLRtGxMQdAJUTn
if77jsNc5zpGSiRAGzhAQAIwMW5Zsb2w1xsXo1vsmzMzRQDQbsOw+upcdwOO
D+y7CQ+epVpCGZBA5zbynm8I5WvvnkAz4oykXaftih9hAeV8YwSBQ6PaOc4C
DU5nfb/QsHXzvmLDgeKfVbm8Sn15px/D4vYVwqZ5WkmsnQ4hnKKIrlg7L6uR
U+P3+pZOysjG4UVNYyB9dNDclHcinHsyqILsevd+m5dC7QsVegqAzXygDwUC
79p+xJXjTLvHhMIhcl7CBrzABoH8EtBUxkIGHCi+fbt4R7bhhSlBrIuCAOeR
QjYo564QSrb9RSlGS/WFCED81s8bloSct2uNMIjctGJ+8fpX6pLlOt8hXNNT
z9joFOCXKspI+JKG1+LDhiysGs0pMdugUCkgWTnXyW4bCEQt/wL2z3IMehgc
iQC4wQ1JcMXDu7791sGQRJVQEYcQ5MZsFRuh3lCzpgPuvxkmq/bYHzW76xz7
spxOR8yVnwP1ymsX9M2mhpwwTht/PiKe5a4WslhrA4fGect90ZCfDY6wFu9r
KM0eqR6Ku7WeApP3URrx5ZARK9xmcnuk2oTXcgiI1C0Ukn3ogoiQY3BPqgXZ
UkRHENMQxZXsJaVaX4Rk/IXuFM6lVqVY2AWVpiYIFaEdsEZZu219PGcvfo4d
gbE4VPPCU5xnnwc1Q96aMmkfh7nUFemkTUexaoXXRcAT6Kb56IFh4MWVZo/5
IPghHbGQW4vng3OnUYk8IpwEipatrzC4Y7F2uVlAOr40Q2TXzlGUMnSlrypk
VWMWlHhCjthLDYwHnvwufZZjMc3BLXsZ0XB5yo6Q9BpFqSu74G7W4wVj/miS
l1RRi0x6LYn1iXXKgZKH9VVVRU3yilFZh0cPSGWTnXLyMtBvAYFH1k0Uy40Q
Vg9MyfqTqg4PamxUePClfZ7x8KI0LTOAftHQLZ0O+nhG+mTtM/EPucskLOU3
yjZJLR0KGvaw9O67jLG+Pwxc3ujsUJpcgYaM1MSCZjy8yFaysfUVX/hKBj0r
QdQHZ3HUimaZTN9f3Z8tuz/w2JlaY46iAQnoU9buhJtetDyD7NNHV3BiUmfO
sWE9MCronCFDoywmX1N5dzmhPhYQ4JHfJ6KDVIKfcQ6aNtyhEfLBNN3MnONj
1EYDqmgkIRMMsvxvUhFkBTRlBGj7fDk5+Dz8bx5uswlS6m3qvgpDQTHKIJqP
GZN8qBcsKieM3bi2cjLhWtmL9hgafleJ0u0ykRKqXSpNUELYdVcPK0tXS+J/
8dKYINLYIKJ/QcxJ9zt59zbuMwwIC6HimlpD6FRe0Bd+C48X7ZumJkRL0pOU
j6o1/LpHp18l5fHFEPSfV9in/1WD3CywnfTNFK2PIad+vfs9MsQXlIkahaxn
DexFRoq/xsRPzNdW4UAX1eWGjZzHyEfj5JkUbxzDqCcRGYUKbkjWsfthN4Vk
TV0ovW0YbPDJ57SrZHhm8jWAwlG9cloyaGHdBZiITxnYlzOt3CIbFsjif9n4
dOkNIFdI6Tf4j8RCnwlIPwpQCxLKYK7l+QYx28Jn4ZwMY+DkfDkqoV8nXyHw
lflGg9rNb46j0XOW5dxTCN98rS0dOkq01yt6em1Cg68f/QFU39KQMPY3YLIe
LlCRSeJ0rxxS2qpMu4XBJAEFHXyU6Ir8hJ5LRjG7FWRORHxoVgb02eK11JeI
Kd4PIv9Rr0lkBSnwm6w8ClScqJOQA9mfPN+rjHRLqLslsP7c/IftROFAJE8C
vTsd65ZlGBGyLykYYUpophSqW61JJNZCuloh6FARCfQWk+yWhm6g9vjhaDp5
HcDQ9A+2hPte8iBX2/T/e3UKMq4jozz8W0a0euHWTX94EzHJxgyIaw79dFAR
hLWh5/CnhaBw1An+kcvvN8o5F2X9P0GqA7BznXao0fxcjfglSw2lEJDCF4OL
qgQykZ4Vw6LXTrEb81VKwwHutbFK6jf11A839TpMTgYBFj2eps2BBzQdYwEk
VIvu2u5ESj6K2ab0fJuyYoBduBeoUfjn5T2ml/xoiTq4H8Ks1/CngEHqViEF
IhUwoLW1tv/dPta/EpvgM8zeFbMEHOZdPpz5ix9ABxepR+VOtRWuS3G3YP/7
q+nglCUee3YOZ1Ip+A76VdlSB0jEEAcaZcp2rUrfGT9yAUp+FWrmVZAAUTg1
ne+7XqrJ8L9beavy1A7dAHc9rbev5IHn3iflkRqN63+GzQclWcE8TpKzG7cU
RnPKEOD4l3REuAMy1gpiPgiqovN8kbuKVUvol/xoeYMlLG2xvAgX8wXoXjjx
ghsqaXa1L8EkrIrO8/76IKDfqLbkhfodcFEKRMQGI9XygIacBn0XZC4tSJox
lA5pOTv23VMDSqTKkI6587r9TjQ5cnV7sEI2d92G/uRczuqJX5apjRdczDOE
CLkyBNcSI21wbQ9Yvd/PGSTnyNkNymqaQUkU3h5Oabgloudv114K2oU+Mdvh
uJFTI6/ZO/l8KPw+PmpATDRJFra4dlJnMBrZQqKItr2Kx7Os/Q45/XZ4NHbt
s1ijV1iafv96Ntt8aDNApWgQ9dr3mVTnb+jxt+hfijm7RXVfXmL9B86vAWND
LpRciRYeT0WfXdeRppamBYhzPsSP4a5c7fhKo2wEjvi1thuigximvTRJFnQ1
GfHsuJEIIwuE/2R3iXD4BYeiCYHx9B/HKnPRlw6IMZyG89+zPeOCOjVDafSe
6/xMpmMnYVG7fc0OTr0ozvusTnNZqssM+YQfeKHobxbFN9QCS9qsMk4peVa1
g9FDrH54sPbPZurrC2wIsTKD4GjLWZWgiT59svDYssuPVO3OvwGh8NlrwVgE
8icYPgt5ngISZrVd+9lKLMBf6hf66X9MjXXJLNbuwSsC+3SEw6Il40QOn/Qu
IFVivSJ/kWYAjy2HVOpk9k0OSeKGhx7XWbKrFmCj+mHTjPZGP9biLzcbGPnd
ZT795G3yFqq8zliA8Pb6ZnbzE4IxfJdGFHWog3LI9fKJZa+a+iJwDr1R7Ly1
CebjnIM63s/Ghf55kcgPgs2R9PW0uuxk6HMVXGNihnayb042r2QKUsXPQfLK
Wg+Sj7/WkTYhHJBFMtoVM+goaWXMg19WuYiS1pfuX4Q6YfXjLeVJK61kP0cX
xkuWfJIPpG6pJIbe7ZdpZrBd3a2bcvj23/V7P8DN/KWQ7ozVbz34F2nFMyEQ
zvt1Fh2dqLLYs3BKGdLK29IjY/XjiI6jxjYs7hdw0YT3rZbpuWgwl8fhEqoi
FA+lkFvm2jv7CwBWzplxoo+pJGZy/AGRUgd9IxGtEFVMw0sqdHV/2nV2lTWV
lWCGV1Fcvtso7EolNv1gISJm7s5KKZ8SW7NWI2uPxSgpLLgtf5MSGsSf+mYs
ISyB8mFG/0a2ReTUgdVXH65Mncwov6vgbch+1eEn8nQLESnOkVJ6ewLuW21M
tvr7i/rwV2BA6/sBR+Lp67m4GNL0uYA9w9MRtITrNbaMPO7dWpBl9Du0XUdp
RiZZZA/0lr3Nvc5LG1iELVTUKZF010skxJohpORvmonAXQV5U3hkB8/9S3Hq
goUPcjOpA+AI1v2ZoId3YxQhH4kbfn1KOt9h1JwSIOwuLe7WRALnBhLQEu1s
+cgScDoYxbzbSEVCYkRRXikLYOFvTspQt5/Ms+q/W9m5nJVOcoYv74VD2cEF
cHvoXtyhSMe+A1oLfx/aIpnulmTEq3OeVscro5v5WcsrajLpGZUMKcqSr34w
HXP8HahnjU0ktb6VSPNzhJ5FlYZzmneNGsaEatnoRzPV5fiQ7/AIWm7Tm0F6
bFQYN1x2+60Iojrjspv5j+Uq3nGUfSZVyknYFkqZFmH4IbLuuHc4gWiihB+l
iW5f2CsU/9rW4+usHQ42oDnNTfAziibj1R3rAPTpXJvqGbJ478KYVZgV0aPs
nMwvUGFj+K+iEwC4RYxziyyA8C1FP3fINj4ZrHu2jmcSzimKhhLhiNq9UX9c
3oB92f4MOPCWqnf7bmY8eI9dcPNwzEGGOgY1HCo8bDcWTm7rju0jeyrxRT9r
BLDu4LZ9AGizu4nKxYByJcqkAAfSjVtTyWcov1I0wNu1NQIsTjqmpt+Zdb95
8cf59K4xr4Jq6mWDSXpoDwIhJNnaQW1AVyi7wlwmen9tb/Dsc0l/ijS6cqbb
BUJRxFJnvPewMwAuoziJIzhD4l0OYaeWtlUP2W5X7Oouilxg4Nc12UINYoxo
kfxdRTzv8Lkg6BCdw7A+q8iZLZQ/TZl1M+LcFCGhTcH8KIEOQCu7FI0ZL6C8
8AiN8leKBauJYV5ZOKtlPIxKIZBg21zJRWG3hDIFsEnqWZgakY+QpQ00m0j5
TOz8ou0Twk7loMnWww5ZRo5StO0wXyNTlPXKJIgFJHlGRMvPaxLDkF68UK1p
Gm5v2EJFwEnxtSvrqx+Yv0TD1nuMZmru+uuHebFPjCgCDaqZ1lv6Ay+S+IrY
rtupbN9PtiqgS3ExCJo4RXnnQXI9gcASITCN5fDFiadCRfHylA4XRciRlw6E
pDwuFq2l8MZeZt/zlUJxA9l7eRStonQ/5/5WmXICzlsOfwCiWNRLwiOhunhu
qzBQ/k3syy7f3grNrWazebXRkS4Q6l1lTR62cbmDg8i7aJpMXtw6i5aMfFCv
Lk+pqVoEAYToDxu7HmJYQzLZL4jUD+77V2WkX0eBSuE6JMTynIeJ08vSug0N
ROVdLaT3Crld+Qk8umsD09omNYOxXcKrly8v4qd4lgZZMYVL/CzSPdvQOGXL
Wl7RRa9fhZ291EvutzEyyqV1zBACb6pDXKJ9JOzm7bzpXEk2q+YgRvnpeGeW
kcVacjyFoJ1j37eqOL4WK9L2WzLIjE1WtT6fxHiAJz0eOHWbwokgHLGW0INu
PZTpvTEC6bu11l6QrP5boirUJaITDA5HzrY4eZyo5csMdZDA7LzKTqiBgoOC
EVv5H6bGt8a+jsNqyEQRwBC2615DPhVF87Vz429pwnda2BtIxDKgmcKmNmlz
cyGN5dl6cbQK3149I0lTbqJvlHb7l7T81xDuKB9+5I8X/w0cLNbnZLuLLVKk
uVclIHN0LkrxiZFyRVgzILnUsXzZLTt76lXLjG6PCJdBMUm4uLuTQ3J3aH5Q
uZSJcjx0abn90DtUcGkxCQrj2qeHj/NeYgcZDpoJJgFOHTkE/m+vy2Amlf61
XQmm3tftyUGNNOA+WMlI8Y/qVgZ8SAq0xpKN/pv7Tqqd+PsgcYM8H8nb3Ms7
CaQ5wSXDShomxmpoxK7sn6WC2fY99EueKtTdlnqK2EVZyjxTikzWLDQL3NEy
I+ZrCg2dTUwbrlgypuWL2mjklKPMDz+9Xtlx6MMRfWEXaWe9QuT9KjogH5NH
lnrBpqh4xUKFKKlG4EjUNeONkch0l/9cm6FCi6Aoqv/F6h8hqhfHyapJd9Yj
xmMEpc8BwaQ+7aZOPIio03rI8gQbWJG5Wo5h14gSkZ7ExS4uRva85EgmcHlU
ICz3Wh4i7vpHZX4OoPRcBIJmLZUdbw32YoG9Qn2Hblmd93nw/jiRaZGCBtwh
FFn3mxthFfqc0QIKw4POs0DMktGiXrUPcS67yxOYCv/w+JjEK45JhuziIDBp
M+6fshYKxRdxEZTdHBdnzB2ZxIbv5WcblrIZoH4IfJjabHtmVexjONJGBJV6
m1eJlN1wpIvRKpG0/gizigxtGQbNzMJ8CeX/03gVgAQroz1kRtkDreKWTW4c
KRIBLE2ef47DgmwWQ/ECDI2rX+ALxBc3DnUZszBXxTMFv2iG2Tnhm93n548W
F1M0Yuk28IpJCuF1Up2S4bETBTmr/SDmTPb7uG9LfK6/jBsthY8mYMAqhiOy
8qYo13zvOD8LzNFEesUW/Q45ADckc5zgaw2Bx6LEhmcnbxd14j+U9xUbLpSf
3UqwgLeRAcP/zDZJBxYZW/u6LwncpeLIa0AEJfuL+O1XX6lzlj3e/9UJoU8K
VG/lfDEjuo81lE5sYRlDjp+1REa0UiaU525hc9jOAw275XdNuKWzfeEUKZwW
sgB6OqLTFORZlHlYhOzhq9oZ61fvcybFUJgX03eLbtahh/mGmE/Mah2qBiu2
sSS5+ayH8Iwoenez4ye+DcUiH55X0DEUO1ij146VnkyG8bKxkBRMAebGb7t0
nzhXxpBZIwq/tNhLBHztz8iuI6rmsklapQXTlMRnu6Xh/lDMYHTu3giPrqky
vuHYzqCjgm1hH9xWQwyZEsWGKm6DkLcmDft1t84AZ/d1Q+n0bm00MIYvnTF6
el/BEQlgZ2F52DFHp4Nu50QjFPQgugNw71SptfymjSj2nnjjM3heGCDj6xFB
gljAE+HWqQyY729VRh6zTzXqfjZVAhqijBUz+Bzzrt0IJ/0pYhvO9EO+ZW7s
QxsqH/z4ex9BnczHviEbFAyokkns9DqK+nnrJwN6GC95eqmHdvxNwOMkFCx9
L60ly9OW0PfwrSXZcNmMJIIG36dFKJJHRhTcXTfrFECeLNyxsy20rsq8KA/Y
z6wBuu7kF5VIBS/GRA1wIITkwat4qOAyxEXA/zfc8tj+NRLw/6+GhtHw01AN
weTDXd5M9EsKtcAV5JUsr0ZWc1zAg54Wno27b/KE5oWKPo56iGLeTBCxAaq8
2XHzQHPorj3uQBX/fKIJI1whWuBS91HJ2TP7HHpDnV4knWQwT7+y/60D2/eh
96XBt/yJUJ0dnnq1i1P4IMZqMfffNgLfUMSlCCewdDZ0vJB8wLX2BrHJeG7V
Jbus1dUgpTHJkeuDb1Zlcaouhbs+z4KfEM9ksmb1kf/TKShlQKvMEiaN4Q2a
L+1MftTJ3268yCfJlAtCH1bMN/xe3qz1qwiAkPV4IGm3YWMUxvqgp3kOpbVJ
Mf3AD/L3YmyPxpdso8m+ovoHt8qz8QjWEdEtSLyYgsMcxqhZs8tQI+Iza951
39tR8vY19bvQITNa5NqylGGn/dcEvtWn162A/dsGNeUcNuulpKPHEBriP/Pl
dza32KRoWEt1nHvCkYbpWOyHjEC7DB86x6freUFcNvieBZqgFBCB1SbUEQzI
WskeF0fNqrNpbdPdmqMEjLRCHKMYMzPZyqbDytgTvn8REhBaj3n6xH4w4Kiv
a3uFxr16fewHC4pz8u6zFitLXp8eg6sAl6L/BFZwVbpeMVx3NvQ1bJlPvh6P
bYumqC0AnWVFdgOjeHk1aGFSFI3aHijuBnQY/MSNogHOrUILQR3u7elLxZ7u
UCfHF5DntWtfeSm7+ovvXk3IumGlvkSd2dwx4halTcsj4HKUghNptS9PAEfU
HqT2bSigHT04HpR5e6r1a3sAbFLc64uTkGfB5ti4PON5Mul3qchMXppAoPpo
0fSbrHLpCa92GxB+4vZZlGrMQXDCYeuliKHCsnnuTcD1YIqRuwMI5KFse+cn
6cdvpQizQ4yb7vrh/SJ1tbvbmbmWOvQ1ol0It/dPXRUnOkDzNyrJoFlncJMz
1j3jUyb7Mw1fJNiY4VzCMASuhSKGLbVB3wwRdH7aIbkwM9ysvyJEbEGNzvER
m/Wop5WuzjNHBspvShmF/fjw87AfornVlFiNcVCQbFcv7jU5SppN7v1F+0ZK
Afj8X1mVRl3LinphS7oU2ncV1JFd3BQEHueEvUqyGXI//3W13+6f8nORJDip
3hCyU12MHOoI7cHmeIyqmxFwi0y3RziwVFu3h6x96tdm81+xLMjKGUxY/uWO
3Y4tv2qtRWqYqjX+WJQWBMg8sYfl5dZTg44mcntUB1D8J2RAw0Y4Cwwi6u3C
DH9cOxka2TD0FP9PERaso1I2f+NQc3G2JxXpHmu01tOXw9jS6tO26jWAYDZ8
WFjgGDnb9TTJA4MTtqzuj+6MjeVE6xlGrPLp7KHmsw93t5C6wqmLiocbp8/9
Tt4Km01ddqQFc9nHck9AqMi1gPr4cn01YzlxUMqGUm4Wk1J8O6iN2c8Iabxh
iNdLZigJtNeS/7yUhyJZO3TCn9aEEFpJL+GgdLXg8f9/PUIXMIVAmLJxfOw+
1SVk638WgrR4rGWqCWgTJPosoO7WUUSUyxqnA6/hU2gYrSwSt626RPSpEm0w
7NFLr5kgJ92t41K4ANAfs0dGSGT+GtDEYvoQ477oDni3kT/P8QnhYG0XeQNY
hJYym+mQYxZSW3yyrwSl/PmyGOj2J6B8mCXExexEY1+eh82ZxGvN5oOKGIZX
i226GPEBA9Cz3aphJcvwJcSTz9X9hltBdLVsOUdafx8A43zstPI17pac1deH
eyQhoUdcquRxmghEK7mXwCEBfacf/Zv29QN5/240dt2nCbeWkYA46LptDXN0
SuLJu9kR7c66Gp/kjfd543yP81JWBgS+fKei1RkvaqqXX58rRHb5W8Tj3VMD
WPmSmDXVLTJb2k9D918+OTG/cDHxlYGawjOKsWUj0Gu087R+KBJUeUvrkHr/
p8GOkNOizzwET3lqr3O9MoZaJRURlS11S4xeSaQa9JCbpozPxPfYuvK9A6J+
Hh0iHkpcgZ8Xn17NwxIfxjWI2OlA3Nuai4eA1LFbkSAlvX2D9NbNYIJ3vDuf
H710Q9c7rl07ZanFEx7QgWHQOlLeU0KbXw+lrIjhVEL7CnPUeMEtA3vrA6IP
pFkLHX7n0OpkJ9Z+rgcey+Xj08rH44zJ8EXWTx4DFKjXA5ksw3ZRWUnTfUI5
sKEsNYOo9vfLKFM542dWugGZiKfrKj1BFezzSt1Pvoy/fzxAy2Z5E+QopOCu
UK+UjGnlNnwc9sKQLRmN9cLkd+lVFcFIVME/HsE3+eAYaoGTm1sXeEhZeLhD
gH/eaXv9MCTDG5lFSdNUw89UM+AdKxR5UXBijPE7/702Vf55roRZkfFccJRZ
iAfzY7NPkDZ0CadQwkiW1zgCeHkW0SutDR4vWRoSdlzLWSjIyjB4qGRbuSNx
zcU6okmbNA3fqJbwbsp1m22chZg24FaxPjP2QUequCMwBT4u7QXDfBssbNCd
lzuUNNpEccpFBGpLFTyOkHeFWRChrDNPmmFpxZ+RbGjn/YXZufkaFdg+Ifgt
JQn5ASAOJG6m27GZE62QHQCZCYWZVrlN3TOX2deNwme7i4S15ccMCMfa7hXj
vImXVXdw+y1EYisyjvzBz1MQvy0/TRtK2v9Sez89b2Esw5+Yw6ykd8AJ8ZID
y99O8iiOJbwKAt6d+LwBNx3M1yUmTgSiloGK0vE04I0E89DEZ2rV77SbyNcb
c74ObX1bYAxYig4+ne67GJ+uaEh7p9f0ffqaNKRDh50UHY+5AcIxtxPfIWK9
yf5kR26okE4Gl1xs0fO5tucmVTpbPj58/QbMpSXsQRx9i/EB1OoiPTx/AIw7
uUXMumfsGvMj/4Y2Pfw+FDWYoIujipqvScEqt+37neaqC4HGCJ/rPXrBLCz9
cdNFFqg5yY+xUZiU74hXeTOMPalwC9c6VKIzQndIstKBhW1ognn38N2d2Sze
J88xDx6fwLQZX1Fi+bwROvLfoKl1YwSLaZcUWnbTPJqJOoSGJLq5l/esDbJk
kVSWtwuoXF1MhaCMWI0gUPqseKTK/eMaF3ESCbuxN8+MCRjUegy7Js0f+Ftw
z7SymiyxEAp1HJ2cCvKugfWXfvL1VIkRcJ6J1s4ts6fIQpGPbFnAH/i/jAIU
/ND9XXlfjjkvDLBBQo8xmRK4tNUTSeSWCgOhHhzseKYDDwSO4q7vVaCq9Q0i
xEgtgNdUjJ0tGojYP8xQbhL9JONwKbml3wjMWRqv18b5nvG0Sw7C9JmHMKGw
dniGCdmxxDghZOvjH8ZJOoPeBC3Y6n8Xnk/rJkE5SgH8q7dH07vAjsTNLJIt
lgy6B2iV+JtXLuXAfPgsBVvYcaYgC5iApFX0esdBjn8mFBwGrcOtd3R7IHs9
XkiOMtS03HEBcAxgIdETRCanKeoL4IbAYSXsZk+tnvBhGpmzVh2Flf5ncADD
b5VKSDpVHIFYqt9V3+cnlmHlgDLN8afrmqNyMQni2Hazye4GbigQXi1YRWJ8
zv64N7mdkTku+eEd/Jn6QbtC/ZlCVcASfHDAoQfzfYHna8qLWSHslpRS/u3B
gEXOo837EIvAVL5TJhx6geayHvuuBlq2lk6XvOFlE1srf5iqh7s9/V5qawA1
Ap7a/0KdY6+G8X8XWRcaHPmhKl6vEICkxexxFOhNh3SkyWMESAMaMb5CiFR/
PpLZCRcUlKSKdrYd016D8pPGe/3NrTaYYbqpbV/8BHxkJIYrttMt7o3AHVPm
KQAzTofUDkR6SdlBjcZg04sz3c7GAC7dnwUhXODauCOhJ4LqUsSYYnGHJQAt
jTw2CJu50TDi0RlPApAV/SX1bw9O62JmKDrW+pvcrDvbHtwXKBVSozQ/HGiN
KnLhTM5V+nsMEvflY28O0KM9foscC3yPlsX/3qqshVGENz7WKoEeqH1xs7n/
AqN1DbDF065ZYEXeglRsK26q/HSN6k/5qQBB4gj6vrL7nDluKBTLQFlqTxRQ
CDzA+35PmUSh1VTM14I0AjNrnMjCMUoTHbbdyM+8iIWKmTpk5g5kzEF0nFDK
PJqypUQLiIdavD6D0zovrWSJjFL5FYOkAdTcm8Cs2NxTKc/w+TNUDbVYURo7
dSm36Ur/Dj9n+2oBnA99k26sJKV25PkcJMBQ0q/AcFNfWPl5FwWm7ercvvP7
Wr5HLaklH06QPAtnl+9whWf6qQgIvn9IfPUY61+8pxSdPFWWIyHmpjokCxBB
A71ZGKZII/HRDZrW95Dn10jhjcschmaww9SkUvt2cX4O9qHZZLyaTc6Cqq5U
uvSA7Rga8wG38O8w3/6N8bmbRdGnGNDk9O884nJWPK3fcygO245ejolKU84I
GFKPLAOkFToB1GB9wqp2iOsA/2UGn5efunYoxrogdFTM4G3o7Az42fESe4wS
cKYZZpGKlXmCJ404mvq3GT/6k1d+Qs9XMwpATbkf87GEJfx5/FboRNQgI2MN
HM3FwIUHOgz1XADkOHnI6yTseNzg233w7faO82cFLL8TuG7z9k5811eF4kSD
1kwMxEVpCXaRsq38l9R7CAgy0BdFjVNSFn09Vi306bZ7n3LTZkHJLE97rfdN
blsTOozmnhEYK03VMGbSKPals/CZqyMvohsL27dDUNPjkRxYYHdnXoJSgerk
yH+9TqiWR/c5mq9ZON08VqlpN37yhoLLtp+Trgdk0bkjT44Ew2pFjNgJiYNM
LLPuiu8W0BVoJld163SEtdT+rPhC5IEizaL9DXD7Eb16xXyupKd/Tj5GE5qf
OheqmukPcMV4wnnR7S8z9j6UD2RyKzVr0rZ9F3vPc4ceBoaT+Oenh/fjOUKj
LyXOTSwA8kdm97coxuC2i4Tw2MQwASooic33WIj8Dbg1m0FQzjdq0tGX3i6D
K/iazwmE2GvfbKFoGaqccQh6fKsW2KtZ11fSHu2VU3J0hBtzQt0dX20CcmGD
HF1owziivX8UzZLl2zddTkKRStfBQcRhaAdJi18cztwydY1k9bF2MMZT/fjS
SB6BNkeYqNct1K7WPEjPDNKCUav308Z5lB69hUOPzsY+UrX6h8C6ryCqkZr9
bqjDR54/5O0NzrDZifbpr6NYpAtJFv3VzXsRh5EIIMg+y4iFN3f06fwhGaCQ
kRD4FcjPTXsHU9VXi/OutFsJq+GkYGPHXx3qLl1GhBExqWxnx/TvlkNP9PUF
DnhWolmZuLM0n9HJresGRs8NmbYSzaHC87EoUV2SJU4VQbyK0cUspCY1rSl3
PJAA/+nIHQfr0ZoMutK/qsPhfCZqWh7t4R4MKKKw6GxG6Xz+UPbRLPtFzcfI
HaUn6JlAbk5jcu3tJaL/KvX+254LHJ/eHMg98XdQCOm1LmkWOWRbkluSIWon
+/gRza6yKFpOv99uYWJG5HvIEkfXiVnDAhCkAj9Hut04I2aBRbK1bI5u0FMJ
IMX5oaC+EFbBP8JSA9huFw0wjeBax77H4sYTpaQtEkbHjCcVbKaNHukVGPor
/bgCYKaLR3V214zD/Rz1YaUOLeP7/G3ttnc6vw+dhzU5W00RkNNIGgjQO9s0
iS7EzQVKkx7Jy+AcTFwba2GYRyxXYotOwevbNtwFq+mm49SUemQocW8OVwWX
bll/EUBi2b9WFCFdcljxEeZYD994mvP/xkMM1GrtJTeQmv06GNbsUEWwxR2/
5qvVxsA22DQzybq6V+iDde7n46h+I/5kUktXhfckuJX8MEBs0+TlZYrKJHsz
K0GgtVvwsPPMYWkkqZfAJxaogS2EHJ3JwzXtFcgI8iiD5NPDk5aJ5xJ1ppSE
sZcn2jDDAGg3wT8bg3o52ICq2Ld3N+EddONEa9tTcho316pwxNMxFxOcTmdb
T4Qv1MmoubpDYTRZzTiB/6CkyylEaq+ImgA4WMZSDBWXYFPaBcBGvBYVByzb
HIx/UpcUJVoosY5tCJ5dNy49Phkvwjr3ssvFP/3uVXfDhP/Aro0UGEpL2h1F
28L8MRqpRK23Na9KQS/g2rm+tctSMIx4ZYZFAOJM1jS3/n5AffccaPVkQYG7
+ss44vqGWOoPvQRtQbDPbmyzT+oAK1zvlRTpGBm4xL7iIYzqYWR/+cXfhqh7
K451W+R20xq3iocRGmvwVJLzQa+LDBMY/3ioEE1NSgaZzjvMavDzsxdeUjmU
wHYi5PCAOj/G3xqeBk9b1d2n9MwQRHJMTnEhG1x5sGXE8gY+NazXOQnhUkRL
zIVDyrv3zpWmPGkXe0saRlQsL1bTXGFNn7m4jjIQYj/xC/PqPI8zrddjzx6F
Bm4LcfagN9G9hJpRNuJfjojpwL3FGacRrKj/gsiA2RGx08T6d3hxuRv/C4bc
bpWKqZaPNKFWKSvEWtxlU1dbaE1NjsjkGisPau9CPa+0JkWM9JJ8CYk8+KLq
TzLMiBbT5nRHNvXZHloogiwdOuy6TCv6GV+bdZEzQ2b5/VEt94R1+5TGWDJh
sRdEWMCQb0y7L3aJzEpwJhx/8aKrjZ8eReJdkG85N7Yj69OaFBH000xGtaeD
ezoUApJTWvuSQH4NDfgex/vj/Fn0gmTaE02zgt/3KSXy5fu3KsckBnIfvChg
7nZvANZriXQ7TecxcJfevRmnOoMqAm4/XSHGZ+64OUzl5fE49pP4fsVtclpe
0cB2o8/Yu6PVrXAE+PC50VN5Fj6eQjXa+wbPecxDGrlgNFW6NJGX8HYShCVD
2HJGrHQ7NJLifYsCb/eKmLM9azzupKCogd+7P4AaT16JBlQlACfwthk6MLag
ohRZkTs0OiL3rIC+L/zAnasaazohemqKPRgkFm2FxeIceGHQsxRCFG1rxH1s
p1vTP+9DNEL66kIHAX7lJ/bXFrTTrHFT7jUFypey0j4sipO1rwkov1RdDIpo
FJTGtJfspDnk4H0y3IVcC10YdCsXCM3OhllRnLo4gxvO8v3TAO/oN+AwPdTw
Xz52uVR2t4RM2JeN1w/M0zXqk+J2/Nnbm+Hh6KtMFncQn3y8LBueEecggPdW
R7t4lpDGP9/FBBjSBN4aiPxZtxkk54/IjYJ1HE8AuUXyUBrkr/RuG303OU1P
PP4Gr2TMMwCUkGs/yEPlx/iiFx6qb0wo3/NVslvhLsiGz5ipq5/PgaKTg+mL
XfI9Mx/EzxHNgmW/gjRXyCCxbJIMF+2Xbb+/+nYsBbhQ6aJ5k/6+aGCdVSx4
GT97g2zbXyXXT+QLKE5IikwcXicCAewrEWe+TB4uLhpl3VuMPRVZlBEy9dRs
J2/OC+lRjWFFhVZJGCeliqQl/nQ19bS1uW05v4lI0kGViZAhYUOpiN15u/01
gDzPiX/knvTmWdR8bG4rz9nPwbopYq82UYQjHtJr8HAnKv3eO6fBPHa2Jz3O
laAVXAL7iFAzRxdTyk8ZU0x5Hqs8wVEV+NfPjSdiADzKJFAqat1Tk3zvGlcf
V6Ox+VMx96ZeTCrbe9kVq1v/KLk6WdM0HBQXk0vWa5W3wMx8piACfknx1BGK
seNLXzq1uId1C8gMJBTwmVxfFnT9+xoUxnm/uuk4wvMnEtxtImVuaMFXVYCz
drZqi8wUnooOHZxxRAQheWp/mv2GG8SGBChCgBufrmxLl8fj0EkvVXMXR9D+
uiZGIU/F9slv8a5BA5abtUDqFUlyNlQuCppmrYWT02EIZZ22oGYPHIGr7o9n
c4RqIoE/OS/u2qc4pHh8R4EXkDQisXZK4WTWvBeIRU/AJ2O7TMVN3k3mvGN6
uyrPAKi0RMUCnCXsQXptx3k9XoU8h80pvEu8NiNw4eQ77Ih0tbSx7B+z/71t
1ZgoqmQMHeHyjmVwK5+pXrQ2EIXvLZYym7HD44kT5aKxpCSr3gJZjEJE+fq7
OuWQ18iUnkjirb99g/h/vk5XcpiMhqr3gSC40LIsksTswD+2dmGcPc7KZKQ0
trZ+AA6J/oDTPepnFozy+t/wd13ZZhtMbdWdd8pHrBmWScz/pGZA7cp7/CwR
oVMsXphMIh5J4/AHswgvkdc0dRZFMXnzHUHgl57IcE5WKZXuvhROLxpW21bU
ppnCED6q/twwhJ+zbQMDbpUCcCB761nfRbtNTt5omCfdaJE5l1i3Ri+u1jOP
aIX51QUv4A7sz91x3Nc+UJ2QHaJ58JcVD2ovtrY34gLvbV6Cd+diNc3NwpBs
HpzSjiEk9gu1N9aPYJ2ctXp3FIfZ1kqajqqgGr0EvH/q9sf2JVkwxDoXljwG
N0Vs1hcKxFJ6OYgUcFGrTrdvHELFgJtcHAxo9jsPgmGYmAePHSK8uuhDXh2e
LM+6qGDKJ7UfwP7vKsapBCQlD9v+IIF2MrALkpW2G+J/hbCU77QdWF+kv2Cf
cHUYMgB+MuwP8oFDz1NDnvw4xomgK3a5oC/kbfyNFMxHDC3D49EqvFWGaMnd
qahsgvKM0EKOl1lFZpflmqrdInhUkWIk+NH3w8r4Q0W0KylyaQez119CFFJC
FDH3S3PT9RV1nkzkzKcE7qYFOGYvBEPxqRRIPldo+uT6hNjvBesfMKtdG7ru
SQ3xbAynxOG+eUQIzLcRhdqYBvLc+vuOfdSTFKWpW8vvyBdKHoyOSmFMV8iB
AFMItUqi7ZCDvN+4p5WlHMC2Qee8kGDempUdhrmExyKxsQMkMiDJEYZfHC17
aLdQpr+sU2jEYcslb6q+InOrT90JTcThhjCnKdSptPdXwJM3QomfLjlYdv38
S1qeKlkqbtiqpsf8HSPxaMttbENObv7ON5/Wen3/MftJ1jjB12gOd+DHmvrn
VRuKsZJ+n+jF9tQyU0kCa6ZXGxHn4iE2v6/EMJi4uG8IO2wK8Py4/rXo67Do
hTHeshl6fdanAl13Jrj/DH1Y7+vUsfQ0qdLq5LIlwhDulhqSzIajepb2DYN6
UoLln01lYHHjW6shHsXz7G9uxuJ/i/CbNa87ABfnLjDv0dkmXvaaoQ2u+IQG
FS+Dza7zchK5eG4IOcJJXmVEP4xhbHRq+F/9uMFHO1QjU0SMvm2NtKPkOvVh
g7ArE58q1od0sQbTFClndgUr270yvI+9woa39QG+oaplznV65dASz3q87iB7
qefZy4jHJjiynInK68PLr6tdSbsJ47TwVY+iCWq8h+MREyeuEm+nYxOGCm1P
BwDAQiYODybOmMkFtqOETjuDQuBVtBn5n0lKluevVihn9VyuivticxhmdrXS
JMRDzu5MMhytXW+IQIEktz5ghfrSUJq/IDiIJe6ZkoN8qXe7HP2P+RHOVXZe
1N0Zfo+/kz0ABz+HD+gF9Mg3cQ5SnzO/g5eGf0BazwJ6+uHT6mLEZTE+RKAn
xPM8tlOpEKosdRjPZSf7Di13K2Vhn7aENtmr2faq1GDTsNR+UqGa/HwXCkIx
gjHzSthxgO1/bGczqdU6FkV32ITaC9NZSuUBm3iZqfx9l3D7haQF6DUgHwF6
F/5rosnLaqcSeoGMp/d2W186SYzPqsEbBzUG4RdkimJfyb3syy56/gRdibfy
3Nw7I9nrHmkOFZ6p+67WvMukHcO61i8bny27CFWjbH3+XjvIDDCwE9v5Ckj+
c1bkW7nSMgvp2mfJAKOVo6DXZm8KJRqHQPG1Wx86d3d9b8b7EBdd85osmFgk
zYthfPBrEB/Xy/+yR3fbeSaWDoU8G8QZXZ59DohaPzCu9m8gK/mZhBkSdgRV
rNIv+zYJ1xOwPDhb2d63LhgUogliwN33vxs0EEljRA8WGR+Y1y0xL24+hcBy
WDMarNseQl/GkNL8XhStswXU88YBa+Ld5uD3ZPK/W+wLFuHzU0UcmlLkVZ7I
qqwbZaoptIfOH7WB+ixQBwCPnU6U1gn6Ye/XspbI17dtPwb+9/dsn7F0cCqX
De6+qVAffynofnX4fZrh5fQKzeSgXBy7ep4Dm6UomT2zAFeZxawsau3hVy0/
jInvL0ANtqYvqbqpZd2UIHDQGzJkibf2feKao8N7u7a6SuiZNV7ddAuoNdaK
j3AYiNhSmehmwi4fS4HiMPfvyLSh3LxRDy7CItwM6/RqwNIKFqFHe3+8JfCr
MI5S4wj5cz/+DJNQ+QnxcaRfuXJANjprf5kFpBo/6YmOf7K4oIp3r+WVgXfv
6Ny4GMMXX3uHl144kVMkO60WTiXku8jD5zLdjFwI5TiWvqY5VL8yo4UXQkkn
hUuWRIsO5DX9IliCFn+0kQC6H+wJjzGkh5a0RonSdNcgcVF7CWP18xLOjpja
pa63AU381iZ9Rem2XmbTChItMNELz5hel6DWqL1zfjF3bUZtx+JsqijMauET
viu5geJEOKPwbRga2ar//6cw8/cMB6nZVNbqhE0EKSXCMW6DcxLl9Wc1PFQX
Ru93JAUMuPMjO4TPS8LitpCH7rrKCB4K/z6NrxXh4yuvOtlZN/fQ70hw2Pct
lnu201cM66JVhy1gl3qiIdqc0Ch96jyCBn9lTjVbKrW1pwrU5lvI0JrQdoA4
TV7LATCdos6Az4gHIWfW63GQ6L+VZDLQFKSKfaXnCpZFrUtx1AchTWoVHyz8
QasWkwS5CrRr9MycczZRc9UaiIh9/284j8Rms4B78Lk2OMGgU4emxdkNtSvw
BlwjVxpTQayEJ6wuH8tAngfDqTwRXk9g7wCTBWKE6ZmphW/QOSAFaF1dTDqy
UQ+Ur+a+Wun4bMWCJOmjbrnxZzCbUJ9CXP1OJ6aExabL99ZHLRY4svVJKA+U
foV/C8D3mugsvmg2J3dmZXLQkGiblDJ3FoXTcTUy+Nboulk6RBIA0Peehy+/
0m0ZAzv2gBMX1kNwWhD/pGPRNHiEdooiWfyWqDkxg+Ah1qGAabcpf40OA9aK
GLfgMzB/MRQ98UaU81scw/dcm1Ta6KdQuP4fVpeGMFc+yVY2rhu/AkMIt22P
N2isIzz/qB99+OGubypALgpu+XH4lJH1Fr0fWtpTYp+e8O8+jsu0IsfTCmWu
XQi8UaHn/AN58PO86dttm8/hvaxjFQAnAWaSIb0Jf8TKkxr+2gdVKXwTN1NC
feQEHmiJwXZYyEprIzbWbt/LwXjuOme06Bkzti8xjfCviU3itZQHz+RMMSrW
qxASGGYr2ulz0qBwy/bSUjQBakKcN4WbpcZLHz6rOM2aptvqztKWOfNe+BiS
b/96f+CObPmRv+7HZWFQNIkV7hBVELNYimge6DVH7VlMvNGylyuEu3hinW+6
D7QCOoZ4447LPN40xopG9vgUoE7lDp0IVskrM3+i5g2SzIcniBmxtYU0dsmv
pE/bp8QdH+3rNF5XcDVnW+5Ir8YS+n/Z/waqBlmBdxHTJlHzFs1U4I1aLgd3
embjIGMtTs2xdDKvdnVk6Rcof/aUR2SVG47fRCOFYgPyqDqFtzqjppAfJP87
ikyoAWqH+yqgHYH7pMPJVBuCGj/UGiCIzBVJXfDsknXB53iXpt9G/hzfTBz7
9hHzP/q6rMm0cf+jABxpx8HUJtbJCiso7G/+Ojp9j+nDhHx+kQCA27LRfApe
VC4gUIn0FbaJoG0dO1G+oO3tsOHQuM6hTGBd4Xx8P2LRZ12jb54iC2MbpJ4M
Hv3QYyjHJePMrKDpn+0LMzGWPmV0ASDIfCCQa85pZm1kEZlmqCtriGff5iCI
IzFglJxL9OA7YA1mfJCOvrTcTu5XvMn4CwMq0hK/NzKoCIqZ0L/Vl0w8enFf
oIYgAS5yS6GpjR+WFDayEpxy/4BxrdX0CIydufFt05nVoYD6uBs+WM7m7Zk0
/aJne2iVfg1zkQsJUSgKBWIEhFp07hRHFmuN6atM5mee79DuJpCqbY7tyWgo
fapYNiPFLPHuOGZ2J+c6SJWDgUW7d1EsbWS044Hqbjzl2KkLz4LoKsFimjwH
hrvIb0HM90fMnpxLo7ojhB1GaVygf/vjT9OLzXaht5TkynxhBGKgeAKtZQvf
M36f0IrVQ/6EtsviDB+vS/lhrXcYuybz89u0wx97pYJag/hE9KO+zx1mTT6P
VsLV+QFYxxx3nNb0ThI7Nz2ALcequpa1kgnPbksQoOks14OUcZmLbIVZgGwM
F2BZdCs9SGhBtoLs+NU5k5LvVWUot+sR6tDdilIJDg+5rle/+5X2QenbA664
1kbqhMpbUsEg8BLHz2LnnGzJqnKYDHCubCpKhLUvAZZUEhhVGmsThVngzu+x
XzRy25tNGbEYxAigjcTbvoB3H3+AI5Ke3JSyqyJh+6OkjBWPp0+45c0ZJN4p
YaWmyV//Bt/nhUg1NKbFjghH3lviMzw0N1RDBc3Ype3r2UuE208Sq1olZH9Y
nAnIXV2XTGcUd1QoxsdpdQkdNyWpLnfUGtQN0g8LQXHXs9K0WKCdXsG818dE
qyxMe9325vIv8FKiAUjsU9PniqgezzTqZ+bH69AHnSnlGauObOBVGSKqZQLu
rlyyM5Q0TbpVjena+BdiomSyL2u7oftjxigvxDAWogcLQ6Npc0a1xAHmw0CB
bMG9UOTldssQoMza3MUszjNW/tKOzygKE4AThwjMbzPxAu+s1YqDB2DLD68B
7EKfYerVJCmCIlfbuNFg3uD1rqlapOzdiCZnphLNkbXwfKNm4+73pBNqRBdO
i+P2OnaEsKAXnx+CXBSlMloJcXMmFinSO4zFTqHNi2O2OcM/2NCwLRQpqoy1
b9+1wlBWX7XDYuyVzLiaVzIFkfgJ7X91ff/qkWy9dssJnh/o54BI7HeighFB
FXLoFz8lenq/0IqdP47UvQlY27czFObNUUPk/QSAYfyAwGCE9Jl+czW1gMHa
sQSoTFygpT/6RipFSz4aScxxK23O56aaW+Ec8JejjJqmg4r3u4900mFMf7y8
jSTikjlktwMjMPZqX5IXwwJmpbMkaIqv51R62GDH036kKkjBQ8+QVh+NoOuw
ShtSD1CGFdFBbV1ZBo4FQB0oL3ZxXE0t8znBdayN/0TmZmQlM4B7UJznqBK1
acjmm6UA0DicicOWbX8s/GMqgQdT/S4kT7QKwLzkYJ/ucUBjLMIIbATshNV4
qYyV4YFUtlWkwlpa2qfDaeHNEv2f8+Uz947zXmg82s44wxOlzRzq3nLok2qe
HM3dkCze0jEc0GpMySlsJy1OQSwJ20I+/HToLamCxDgnEekxElFjIgGG35hs
NyW66Gw/apmpVmVKLnqyDCMMaiAo+2pkD5hAZd0Qtn0rXuNbbaDyH7xkYpsK
A5X4ppEWMdixg1LjOCMpLX8OwpsKGiItF+NUohRYW+XaUnqQP6W8K5N+aoBx
Qrs6L7qUKqVRUEDq2VTcwRjfjS8J6Hox99jwCheeHCFMFzMYv6wv4OZr7yqU
X3TFg8w1uEva5RtikInzp9vHz34EXUESsbsr8G5HH9+TsIuCQpKdtq1EtG/D
p49shpgTeCocY6CjiwaT34hJQJaGn7y/fyPGIUL1bk0Ju3cdpgWaJhNiWlDO
16WwjBubePobP9K673Joa1n+2eEy/oQ7qpWRNT1dW5g1M4vZGPnAyCGKFlLM
t8aHNmXzmZSr/3AOtD3RoLnTkP5pc+a2YxsBYo41HLReYdmJ2TJPNkOtLpTr
DFEdqJAkmsFZ1rTT4E/Uy+TaKooZGfjaxM49RUQlcaJPi7zMSNew2G2vm4zn
jC1wZksovzMr2OGZI8K40ifGmpWzwoZvx+uI2yo3cpM875BoqSb/mn66Dzju
vJZFTMGFUdl9dbE5hGmjzKtFhFNOcQLmltCr8pCxFBjPkCfmzvk+PDINPTiM
kRTZghqJKiwcugCtVNAh7dJie6r7b1qJC7wrFJ/sDHWVvkkg6p4ovMtr0lzl
xV5B41HhYuYnLLtnyKbXTET8F3qhif8De7wcxAEYWou0TUOEeleVP5idivPp
Ko0rKZA8qY/42K9e+IwRC7/xMlDaHv+v0cBHK/DV4iCctZUhnAcQxnNsSvHn
H7phV5bv5w9suyBhQpg2AipxcQyMTn/4N4IiqCl+1yat62dMMFRYkHOLLdo8
tQxp454zrPZpMkeVAl8KC7/XWtkex/4hU897ERBJMJ3XOIjdLtYg5UtfVr9H
CHPAVwqtsjhWS3N+IhWM4d8J1wC41DHlPS1UIIhSEq1v/YWAKr/VnovCDWIa
bgPMrMH/CrDg85uhk5GIfInluLyV+S0myR6lg1zOyRh//1Lt+SgABX0oE1an
4f6lMrHEY1TmVHsuFke8NNEpfUsNuOOXYMIXnS8WnSwZisdjYDEY73svZUGg
lMrrqqWzZxuY0Bn5sPRFNWYyc36W/NPcOGTiC4CUeoOjC7HhISB2EVWq6FpQ
+WzCPRI3o0eArM+MkDu6NZlkQZsiseA7RrVbTFli3dwTLkEOCIU7JVtdajS+
dQC32MBs9FbqzgRT3Sj9QoZ7qCgWyluBsMdScZzaNXIlCdcTsCdI1WtXjgs+
zLQyF1G/eKu3rkUb2gnp9Q15tu0be/525RWEFe00ITD/wVV7O/o5KzO4EzpN
u8YH/LVdpomtHMuje8xbZdGi61DH6Ip0jspPuoGSukrHNX9wqn1UQoemTRA6
PsCALiWSMWZbaIMQWtJoksKKHi0G9nNevLJGdehHpupM65knRASdAZuOGSLj
7v/idxVLqzguFuLDcS5hEh5EiC0IkXti6QdKOQ4AUpmhOWa2bvihRwQ+pp2V
/qWFzfLW7uPvGVFT/BoBJrUz9e5/978sS1F8SoCVJBcuf89jqLepGICzacP/
QejqlarLGxOL0Rg/ofF+L/10Tf1KPwniVDAGo04D2HPfcAp3Lh1o6GgYnRn9
i+GA9tHovq2UYJ8TrT7vUayOuDb9zFmDZkGt7vJgw8AJ8OnegSbq0l3dhluQ
EqxlKjiNOhYFeDVWsWQaHy/7A31sLzI6P7Wi8zgL7aNIKK2zI3VR2Ewenwvo
lETzVp0nTUD6GvbffemblzWBrRRp1iXeRQptjrb6G/WgJgkhpZGoTj0WxCVu
aiyHS/R2zgqfdkaQEIouNYxZYZ6xK0FPU4Zl9apnUKffvOyVLrGybpQSH+H9
ucr7jUhWHhApCkJ7SvrdJEZ/6n17Cp4Liih1sNbpZ0UvZcAq39Gvyr0JN0rS
PuOEbBJlDPeCbbOZZVjW2mfgMu06IqLA197jabsbXF5vfzKdrCiuj3VkyTIS
qS5EzvG0Jn4HSqXf/DaQU9+NnAS0qNE7YHfD1iilpBKDhrXK+GP2kBuEi5ei
I2i9TTWl+gMj8OJuFXEssy9sr7hK/hPWo/bL4WrkqeRiwyLPl7ROV8+2xKLC
/+s3JaBXDv0isHlBWancQbq70XJE/gcB6lpU/NZshpIdN8uadKvh79s5FSVb
77gMGV7A8AVV/lLQZ73My8GXbLBmaOlcezZzr2UbQ/BNm1GNv0rlQU1kVmwr
9KxFYGdexeqkSE+4OBNOH166l+sIGpcpARmjeJHrSlSXhZ/EkZ+618LXWWSB
BKqD3oTG77Hn5NQZmi23CU2Uwai9+qweEZOzynz2+nU+66Rh/cMytfkAgk5m
22O581+wW5tyGMCty/uYE/M4klMMLThVaKg1re0FlVTcw+tWFNPn2WDqs0SR
WH1MrxKWpj4UcoHWF0kAd971ojXDnk9BOGcKvD8jAzS37MQdM2FoqeFzVKUa
QhqPgnN75jGpogW2/XFGL528MMThDoHO3usajlm+n/se5UKpi9o/XGFj0Yf3
ha6O+1KF5VJWMy6CcDYdqkxnYZnflZ1iEQW/TfPPCkNAPd8KfhkcsLjNQkER
gsbQ7Rx/oT6IxYsYSx+U83S0RHBsBXGJI03iz+2fbdEzfnZUPRGfCN+4+3dk
4iAiGXm8qjeh4HmbuAx8sQk/+cUgiAeYRRpGAFN07guXzPzm5PQt8Ar+IB5a
q98u0cFsO/FhmFhtoMBkTJFvB6my8+u/9SkRp9GTBCgBFLwB0sAC5SJL++CG
LDz4SdJk5INkMMLOII3nhLr8rSE9PzqxFy020rx6YzGOLIM7xzKhjUkIQouE
UzwgWDFUwbaBsXLI1RjfrRlV5LdZIsS8TO1VklzsZOyY1uiAfTduMDXFaMHE
dk59a4ZnBy9qu5W6aeFQGRecoOmlcH43ZUFEFX9wADK0nihxw4P2zctSExGE
V3ynRH+iDqy0fX4N9/qCjjDR0sIyujEPkAshWbXDSkoOyZ7s9zRkPCc5koht
I7WE3zjYe9Exh3EwxmhoAMj3LvNWWWlIGx7bo4xtBgyVvS2IBzsLvR4gz81p
CnsDKFvKcaeZkgaA0y7wzNeAPProJrnVtfkxvN2Dw7K5nq5vvw57rg2/Qp+b
Og/f8yHOYbzIKqvP0puu/z8NtswTH7ZH73A4XHtzQa12AsL+fk59UPyZB87j
vReNr4SsYaUenPPsv5YnP5skLqk6YD8oc8AvLm0foststKuUyxQ0k08bNgGO
QN+/n2H+r54MfJdwm83MYiOORWG+3NqeqFZdhlX3V6l7YvXAE8qqTvM09tVl
aILo5UKqWhL27NZ9u91/NOniA27Tand5KeULS88thAK/apknQtJvRYqQhGOT
d4h8nj4gdDiW2WClNJf5smuHSw8YlVXO+x83eR8hgqqLOW8mDpwg+rDRS7rl
VdLfxT7pqTkpHAM9iO9NwaHTDuGakRcCXf0tnT50hLhnVDsYEShppFW4pOcO
Efj13qiBkuhMUT6jF4fXEp+f30JXa+9Vyzl0GKuaHOb6QXqDPAA4rc19KW2S
/WGxR8P0DPoZ22Jk+R0qNTyy1DEHP18iNuqhfxqLxtPVS16nU79P2wc+H1Dm
aiEo96IOowwhFdUshAzsa9nFyb2IVLiyzYP/BIWE7c1oy8idbbnChZbmVnrb
BFFznssvKfwK1obiLWF6875w4ZyVz/lvU+sS9rnMEfiYL71ThFF0yCT7h36o
GOVKrHcqIa5FbEkl8q/o0nzL1lQYBG1JwpzZtnklKGfk3SKOkGHWCP8U3mII
ccvbtbUvLsTRNHt6achzK4Xr1xq7IL/U9z3ceC5UoRtQo/mjkRqA6CCBvtFZ
cdUNWHP4WhNr24CHbzWxH0mFEJ3TiU1PeoTmvGrTPtCK44jhcuBiHBy6QX0u
1uarwW2YPtqXmqM/EHqDCTJvNFLuu4H1M/bF+C2l4fHZULz/yabi9nSRdHBV
PT1QL2pL1OCx3BgbO3cg1M8ZhjK2VrXsA5MJFvb2QNI4fE/xiwC/JlL6RhX7
pYbLexGJyJvIx2wbJbT9Cq2k7lOODJe2oJDSAEYRElKQSUVdqwOFqXLgOX8+
3zx73BktQL0HQm8vZuDTaPw9b6ViEZa3JQIei9VNywreMEzevI34WRxJ9JDF
Ko9EoQKCA0zIUSzkzBY/lSIH4M3I5njjwboA2SX7NW5ceS3s7gilOuH2Rdna
uNu4Peo0uS0MkyTzV64Ly0GNq5/QnPNEREUNL4J8k+bhqoc9ZL4PA4oj0fKk
YeMolMTRdXWkgSascEeb6Znsz+IrTFfETZpFZD95jPIY0av8sEweVaUz6sfv
1lZ4CsYXt3DuEcJ9AFjijy59n6qAG4zsKeVL/BFUhKYFQMw0/btok3xNaWuS
iSeDF8LGWsJjEeWfNQgHyKeuFjmN1oN8Of0CMureAWKvmHGPoNPbA8jZW2d2
KBp6MwYzyNNXmBd/AprhlERPrAxR9jh28QJTyEXh5JL7cfe7hDpbZdZUV6qd
lpWFdvzAOw9eRgN6MUOePAQ8AdgGnj6NpWuvbO3dQgPXJOlhDPfX/LnlVJCz
DYumuNEy36s2Uq8RW6EhaqCti2udDxoEvjPihR6vG/aFL50XTCmOo11hLiQQ
YF1TuClXsuYTJfMitKqeX8y/XHgBEqVV3kUz1+3g1kIcA8bawFG2G3u0Ydqa
lDCPgF1+T4PGX3a7WDrDhh9zrbGpnQt2Vr2K1k0tJ5T+XDgpOSbgUWRhrjtl
TDAA9sMv+f4MKiWlj3nEG8eYYoFl9Pl7+pPz0Zd4/m7tDW5aSt5UOMRTnGSM
IuZjAm+CE9D5+rV659Vx9LUPcMaaXBueN9VyNkQKM5KEVt8SCPoWc4xE10l0
ZXbugjUwHWiY8c/uecY1BLlDIYndPzb4+Yg81Bkr0Nj5Y5IzVHDH5wLuUMoW
a3uuk/S24XUYGtjO1o9S6sGsbfeOt0X+UkONrUwHGrryrPFAcKH6FQZ1nZbf
Dwwpt+GTPEXSBR5qQwYE4Y55tjGv8DxzPFgbi8isoUeajmP20jlsooA8jWuq
nDtcL0afOvSeo+62wulUnw7koTop0oh6Cy/KdfihXJtdOuJG1CVTlP7AuYDK
Q76OTygKc01UR1Amda4X9tnGmjIjgHveQNmAnKZZ78+WUIM5nSCeUkF8sQGH
Szftc0XZTmggTyLf/TP3Th8KxHkI8NsQLfO60uUg7SzQ/bQsNOHJmspzoOHP
cYzl//dy5jl9Bfl1RlpTsbFprvW0FILWHulZ2UvmCLxQ4xRae3w4rwEeUPUk
k7pu1tpSqkBTNyaCd7Z9RCE5ZRFdA/vtTOc35wJtoNV03xol+h9rI67kKOIx
m2QAwE0zMoPw9a1LmSOz4t8wBaQbpRrOqlcfgnv8OnkaQljzkV1/A4lo8cYQ
4CN2lP86ttQ47W4Y0NxL4zvEvbGKLgds+OHqTQ39WuaQFhd1O0zjeHi9xjN3
aPBZCN7BROSEye/P4nsau7ogdITI7TX4v8yl6r0trSQx2z6VpYy+UgoN8yVI
+fc51D36O0X3P4STi4EcU4H+gZEbbxIAFjSBABRVYLGbvV0CI9cu9j6actvA
cOo/6XbAJD4MhbCChjwtT8rt6k5x/1cAdA20Vtm5LoBa9kfn4Zcj/X3rTp54
bGR3SBN2h6EAXskzNaCZUj+dTfmANIaB+OLQ2Vtls/PZPvtkm6Up2VJYnRZn
50OEVVgDTAWTIsd1e16SzerW3pPiQNDGcKlj22ozepUqZyGonCuDqwkK5oI5
YdV7bVx5TAtlTEVBR5V8Fgo2xBzydLMuGKapztOPsTj5SkkhSDmc4/ADL9Yq
aOxTKomeIRQcFDPSOeOehAZ2cBQd9tSk+85Ulk4L7TksAed0rKrg9r5WcToe
R62hellvwYAVLrYrX5gEciu+U/vrYMNY5Xd/ogVT4fMYu6nh6jgFtS2GBUmN
E4EmadOwO18h+BuvXj/aTqN5xj+loUb/WjPEYFU3YFC0ZvlJbFrBWAp7nzOt
4S3iteONiUyl/pxvXRw2VK53bZdMsmNovac8Q2SXd9lVcJ83W7fUEkVgo0r+
z+Ls9T9aHvnV+HFZglsqIwxD0TzmFLuRonYS9tr4zyh2KRmeajg1uiALqJFB
F6pWnHFGRR/ldrTSnbWJ4BmZbVfZC0lfLkIY3bxykdEs/vBvZduWXXyohuX7
a35uXQp9JLhU05qvI0zv9zSF5AqjNw4OH7z6e2adJwXeLDq1luNJKSLOAui6
o649MnuFclUd15X1daGgCw03yuHV1yhRclM6EHRsgNoypHhmwxM/+zNpmR0Q
RBtKx5M62GokzLQyX6odIeJfaYVjuy6V/lOqh78hGmkoEpWDZsatJ2xRaOfJ
QsKb5hdIeltJ7K14vjU9NlAIISirECJnCsumWjy29cQl+T5iqDJzOpaDVrW4
QEKFwUCOTjhSqWqCoFWHccxXw/ou1FqJy1shk/O41d9huVUWws7tXeh73db6
Tf1W46o9o6hEzylJx7zzguGxJ5wWJT8lMtGbrzR/6iCZVdfwXFUvorsKEId6
r9mgoryroIl4FyrV3K+ySmzsKyJbg+QAx9H2Mu0U/1RxK0S/ef910HLGVZ1H
AvQu4Dpo+WL+HO6J6ii176FDkXrEL7OYwiuLquvVy8JYJBZcBp3w2mDdrck6
SLVIx11gnDM8i19tbwNh8w9O30rZ9SMeWW2Oz2SVZUuqr9lMJKrzw3dxKvps
nYOJeZzU4hpEtCvqt5O0HErrJNQTgxw0D9+JfSElzgrzdgfkjG1DMmod12Bq
eETIbYqZWdTGSXBejKSeTF1wwK6MbE0Na3ecjghMHURVCzXsyTvXzCP0dUcY
+L24qCdzqbnw4xaElJ+APfA1MPDsmvgW/1xjYDOn8HzREZ4Q6q0zFAT7pzJO
43gIuwMdTW9dKY3HW8DCPbGPQHC+lZSP90UrANu86G5Ug/DMyC7PwDXVskHW
vPR6vH2Lt82KL/AaHwGlPQz8MYathNY+z/XTzx0OShbdomMAlwiJ8zrAN0ES
IUrgTxZFPdkvbJRiKmmUUyl89jcyOIIcF4o45wkEhGtrEpXZeO7zYsvwYbyS
zAIGawma7ZVrfI1mlafQN1cm4l5451B9Igh1i+OiFIT80cvzQ4735YS1KyXz
yplFAz1ebA3YHlYKsvLzIWuknrjrgHpGTQPQrUNnVl1i3gQyTk6xvAr0K5WN
KQVCDYdkw1J+A9GPmTsFMQJXCP2pBvLk0GTimaAXAaPpnd+ikqPI2gF8as34
0/yhq8tkIpAgs5S2pkeh1yaPF4CEeCxWbL4efkW/OPHZBUWQKE7WST/BcC+C
jJq+TCG0xJwdoGcHU/URW/TQkftHMB87bM4UxSjJ97/binaJ43j3RGq6BtWi
Q+hk6BXut+4XXOCZojxtZjh6D7EQPmvStQ2At1sAwRn4e/M3HVkOGX7/MD5e
0fsNNPQVoKpRPK0asTYLP2eHbKkt/AwzNS4DgY0+WYCscmfXwFkUso5VPPc+
KdlzJITZ7fF/BkIudG0urtCggx5bRNUrTUuQYfEdEHgSuPttLtPpKLA4faSp
ACUn9Fm5TEJIehxb6PjuQeky0326sWqDsEGWT9ndZzK3+g4wp707ZTpfYgxV
z4Bz5/olXNTHocFgv3Gb858SHecwIZabaaLJCjHdwE5n5wm3y4jOZkQEx4T0
WdRrg9skUnZiTjVThUG8hoNSxWNm991GauJL6LF9cS23bK978JNbxHgobL9d
RL79yL68W7jPI/prMoI7TmGYGFF73diw6p9tKNuEngM/xDxZxzduZix+WPfw
z7wIPpZT+GS6i/epOifHRW9ui+ZRKL5FM6db+Ioenfv8kknXRkLFwKVnfUNy
pE3YijJGFHI1hExyxXuuFi+m8WJupXh1BtKLsyVBOXBGY3fNGnP6M0gasjiZ
1BwlhDdH/MyKToqcZCISJzPCjOuONLFI8kfoQX7hkMNnkN0eZoy6vhrkP/g5
LVY04jEInIfT3iid7+/pGmI6NlCEEQNk/Ax0gNdpeJq812xsPGFAb0w+b2Vn
sptQaO+ZQ4XwPELtQj9q2cWcJ47diej34hZ/jnRfXeVHMH2Cozxfk65shKCi
xjACbU6UQCHmIWub3i0ccupDy/ceMa98dflOSFvJNvvaTEjfiDlwJ7zKe12T
ot+SAmaGuTrb9bVOdQo4K83OPj38YfxgQp/7KYzCg1rCzzCQXn6gl2lCNFn7
uFrpKaadA52UrWQdVlsk9TBzBhQmcczo3V0DN15sLGhFJ89GQ107NcqCAnLQ
AonbQYJlZIiuX4825iW5MxbfrO4NXR5YxzzX7yvcbKvAekieF5mCrLjg8TjJ
5BrhheMjdlaKRJdn1NNne7wH8BjpKNdUS1rucqNxElcMScvZk3/0VooIMxV9
q6v0MYnbNSmUVK4JYJXn9UXN1Tqh3n3wyt6YWFo8yOCDTPCgXkW59i0kgijJ
vVJdAWKdr+mjcUb50/d7EL9uVpF5UtP+uyAqPaZxjSkREp3oOOx12y0ezTq8
/cOacWq9AWtUzN9+T9ZIU8pwzagNagwwI+MMUBR0whbajOGNdfz6YBIQBiga
3IF8+zEF31J9t1ps8O1p2jbLDrMsz4fbBjPCSG28efTi1TOEfWr3KeOViLt/
RryyHQcNXZsgckBSr0vmzOdJzoSaIOOsSwmeigbMkghv9EYQRU1bWyh7XOpo
XEtlAEhRX7TUWJjRTTmbxpNu7NFqmvqWG+ELoOhB9ybUi+NX4XFzePMtBK+R
4Gdthg8dDrHOUkhN9WA6fIeXFo68DwgzJRoKiNUvKNL22p308ohXz8COaB+F
yUMvFy6Yr1GQ2OP5ixdiKOKG2W2AcJDWvZ7/eboiU0ZCOmzITK986/GkiYeG
g8LkFgCvGPmbh0ECgmNZ67/oOxj7lT7JoJJyXBeUJHBLvyTnE9Lls75YJxIK
JzAzbcTqE3qh5+Rs3dgXLIj8LHKh4BYQG1gXr1hCy9tKRsed4Ni1WS9NUpkN
mhxB+chayAKQBqmiWVfOEkwXAgOaVv7IK33JEvJh/2maXP8Vt7+2ONE9jSET
OU6CY4yeFL1mLF13NKph+BaJEbULlz/z0TUt4LO2b3dnIk1wlTrIWEG7xXxt
TbCIrUXqJXVUVyeq0SNMpjLweYXvZ9MZRkXTJAjyR0HDnw5XMnS9JJXPs3Ca
U6oxqVru2CL7kfdK/BxST1PT5UAA4bFW8WFEusZF9aWdO9wOeSxfx2cUSDXH
iQnxaGBf+2Nllid7e5uz+2CegTA2mejoWiJf4stIm2VdOlG3/WMaBrtvJ+ny
+dDUD1G2oD78AgNWfSmbE3mVEGvZyqpcAFm7myDjGUgHEKMI8aPy/vWPTpGD
zzhD9s1dHifNWem4ct7nowNL0mhVsfwXHPM7DZHX9h9XpBaTl1H9Sr+rA+QZ
wnGRX6RwFwlX0lwCC0ugQi5PXpyV5b5Y4B5W8WVD2foPlLvWcbdhVumrLVSx
mJ02XWJOz/LqIolM6NU3+NlR9cSdyf8R3u6iWNQv2ONogTXlK6UVGZ+G9OeO
/Vig5jJ3N9by+2HnwIpi/O7G/Q1czIssdm3DIaFt9MLOFxqp8wZqdtkJLQre
cdMXW+7p6ycF+W7aPbv5UdOYAQrxYTn6HHlWZJ/8STk8RLXkj1dmveAkZCIv
jbPDWVXnTXO1GtcuJRWPV7Oms+DSPjNHNWDDMqZSbZCNTs0Vkp83vblKMY9F
QXueVQHtKtOjkxGgnOn5FDyajwqlXbnYp5YrlhLm4ZOc67o/2oS0O09XytQJ
m4o6W/5S9hq0QOK5W6JOq+XssmME37pRme28WCNJkoUqWpH505i9Wa9MnPHe
SXleNnUkpqky0/F13hf0f9FxcxR8CLqgNxhHNeY0pH2U7mcnyq56m745/EVJ
zPlxWgJNLCPEK80bfQbvJGF+mDIYXbvYQRU4KFYyB6h3KdBEpYSAW8qavns+
Hb6exIcjnxNKlRd5YOm2jftOB8OFi15kx3y/MB1jFJu8G4OrcfD5upepceGC
BcjiJFeb6hWUEHYqJgnSemR+eg4M3JtGJTAA0ZAdQ7zWmGJW4fEbabTpcRgR
JBdP5UUMD41/Bwf6eYJE4mujv0DAE+YmEyzVbQNniyPFoCAx7pp9IYM6sjuY
Tx90Xekic2EifdKz0DKcvpIaBBFxD0Nz2RXrzCEhbrPxr4nuCj59M4bkAKJ+
UK3Wxjh+6ZiEVm+v40NvLK9f6t70waD4U5JWD4q3Ze6H82kr/wIpux0clBxJ
BAvmsqVgNOuPjDSHXXuSNFafeDKXrivZ28EHV6r/eZZ0pav2LxNbeTHXVS3L
n32TwcPjlB+f4v4ln+44iD11HJlVF+//qhbUSSR1RJOLktpXX4RmnrIIi6YV
h0ENm6vNzDyQRHOWiTgu+iQY47NBYl4lob3ubqBol/tvx0gYS0hRv+zDvS2G
SmhSOb4v/DlUVcO+1HD/AaTw6rokloHJuUEphhLihGrvO4dbWndmsPElmkaM
Pq8sm1tXDgpAb8m1AmE8dqIhabaenlfYIPqQz19YiZ2NDBkFFiQLyqbJhlO8
v4UDFhnFDZ/lcEsifE3QuboTlwXNFheM4ykUqNQXZUo33l3d82/SzeXmBAJv
9+Wj1qnNtFjsvnE3m1oeSFwOa0L/hx3uzAHrD7BL3Otckh69V8uRVgRtNHlR
7QKhwkGZUP/a+vYpDhQ0XdjR4zkn9GzglGF2Rw0s4WUYqIN9eIzow91ZU4rd
ciNmZJfVBjhp9uLq660qgYrHKvcBIvfhnVZEMa5VE/J+u2JI95F2gf1InFUu
xTCDJl7D1NyPfWJt0v4IxGOGYRqqvtzf4ib0A5PyNHNtHBoBYQR7xnnIvbE5
bnNXsuh5tnwz1KM2Mz5JgKars6XIBoNJX3PczFmsdj163kpFi213nGAL0eH+
KlLu0iXVacEtVJJpT2juEGgpCAgwr001ujVjHItBp2Ik1s+edfLN3rTNjm2z
iws4Saz+D+YYBctQKDCKlkDCr51WE2P16KgzOosLDp2yaEj5aiegsuMDLtZI
F7XXk02ZyuXt5XxMXmTYCft/AAkt4d7zP8DMH0mLEd/UEyRnNByVjXCTAQkg
H9603VFfIvRplq+juj17FLK2n9PgSjtrie7fohJeut9x2+3AVbKb1MbDi3xO
LgIdNY5hXw2ZBouqjW1eUfDUJrHNPDPFrJ2hXCGJdYjo7wfWwqUVk7bCdRgK
OOTWbGi7MF283rqjFBPs8WRY25uasLPcmdp+e8bkmhKS3Z0vuRKBewvK280u
Fw8MfCXB3Pgk68IupVAtGE69YifcsdlSG6IQ3N6IUhQ5Xf0Fk6Jk7Snzw5VY
lE9fSJbOa98m/NqSeMEhwd7LBg/0m1KZI6exxJpo11VFTozp0hCHzKsD3cnS
bDZNdKRsOEyv6XergeIKS+e+AXpm79AY3GjOI0NcFK3aHj93a4YY9RO2mFso
1hZBL3dxizKbxOIUj3c47uWyUoGM6hlragMJEJoz9k9mjtbHOxFPeSJDd2B0
f0e6JUHdSQdCDqQGIWOj3WbevTqGtiA4M/cEgjClN0dNz8zdwj9CykgFO65Z
f+prq0v5pfN7M1s5htUX5cniNqoUjorVFeorGAM32hbgYVVpKpWH1ssrOIzK
XlCspvo8+OYDkuQotRbh4weOaOwe4rjZPUyqtBoTu+niUkNzKjUHIWV0MHk9
3jhckxfIsatDDOzI+7tIGV5R4c3iacfcr6BUBexzPsNeSal9GhXJtJtHc6P5
zKWe6qVmaUuBsSaAEV3BTotngWrDYfOVKOVons+zdFeOX8pHlvvYkWKkqqy+
t80yHD7WxaySJ/lBWsaw2VP7RTVXBrqcE1q7/SunQlNCzYWUZH1BjO3RCcfD
W6UwJkbR9PmmMh6f5bBBsgV/I812eefPULSnqob7W4FhWERh4Q5P1uRsw0Hj
Jr9ZUN9zucxtQUFECf2VJ6F1FFGzkEprETvw2ni0QxdnHV+n12Yja4ujThJv
zxo4y6SeAjDF4i/tVg3Li5BQjwcN4Vz+39kduST5C1esZipUQhqwfo4/FNRe
YbfPHA7t7H89Ir6lF0KVF/LWZlglD/eibztNiahoRxvSFubrlLB1ajkbU4XP
pleRx5fOlhXNZnOCVGGo+bsffYwvzyJ/xdzEXRvqCqgSJRczcbyeovr0WgKQ
/HSWltlmQIKmjF/xxPzNnVarhxouuVpwOASXEral7IPdz4zgXO4frs8LrqP1
gNE0aC/6EZFLXOvCX1q6/lsG8ly6fstvpmiHgxZqLlaTrG4XyWmoxTfCthiG
Jltc2oLe6BYair1LV6hbkL/820/if4Bn9YFZ7BmtSk4m+bIH8kEI+wezatox
ff1xSPSFPaYL/7mNE/jtvPNGPuO2h0RdX0N6whUHgVFGlOspNm3Bj+FdfMTN
11KIcsuLGMU8Bwl4P05F7WUbHnepAnW1KzPs9lSezX4YMeBnTaU1RgzkfXwZ
PsyC1RLkrG2BVPuFrvrfXfK/UI8GVHw12zM9MDdZbKSai29kkLduPvc5dV07
H+R7je2cn2MfGCfsyhZI4UnVfp2I5Xqowlnj8A1SH+344WarCHsZ9OnFUnzf
NO9wWaytLr4rOJjDzzuNpgHHiBuwLBhwo4DuG21S4p/WiKYvElxynmz9OqEH
Cdrky2NeFAfKATbtWogqz3AgfqoGn5Bl9aaoAv5TCR1Ajzc1275vlPQK2Ssu
pWYAxqK04lkM3OkOwkBLDjP5YdUQzf5i2o5LBMFxG2hFnqCmsTya9lzJn0d0
AFpVvsg7nD5FYTKS1pWPS+yCxc3DlINe48dxDDJ3sGhvl494gasKKgafgmsC
gRGM46SLr3NDNJ9TkmuISyZaxabia2OVDRlbPbcZ9GtWp37F7BQSLIWFvZkp
UwclcsO5OszfPF3n/3/KgWBRvEFUKkoF+opk/5C1iffqtKRC9j77DLZzAb+1
bE8CTOJJe/zje2T2t4fdoe5Pi2LPWy3l17xhd1N/0Ob4PdLtUeoXtkcYRrop
KEMKzNASS4xNV3CxtU+68dzLUR9ytpPyQ1XdT1IGcpP/C7Z00DKYZvt6s/Up
3EXCK97YXfD0YfkVsfCggt3Dz4KRq94UIk8E+vxH8GrXoHpnqe4LJIz9RE72
VXxws6Xp6WcOAmCQDN+02vbcvzzcTAyeoUBXRYI50zuRsdhH2fRqjBFgeVsK
JCgQqg+uUYsuubTaDeNcblVNIxNQglKILMLvAswDLErAstByj1awMTJ4LCnh
l7DAzpCEd/NGb6BfDKQtvAcaMYIoPqQb/jQ2lrkkI8AoavSs+49rVx9yqHqK
A2wjelep77BREsoXvbgLKALZ6clY8xMT86il8EwT+Y0hzEnAv5fKsxrvYHdm
0JDd30zPNBjDwiax/8JqsGnXEUCYpHZl+1GKl8s3eADyokwWrCrci/yw3GJH
pZr+1KAlX1Jv20cgcs9x/B7vxx1yYJtslyt84+S4iwPx6JoA9m43BB93FWCv
Nh7hqJKmwBh95Y8zDYJqC7E6T7CJTNzPbfW85I917gD9EO0wgM6SWglsp5u3
FUGxmpQ4kR7W18B65iqeUWuVZmR6P3rFgBs11CUcrbS9CU95qmx3ZNBCoNaJ
rq98YQitYlzGgHLrppfLdJl3kYuGlgHPpispIOJx31yDc9YicfRxkpGc6VAW
u2ea7tUPSgdivirX562JLogIkCgljHlB8XdnbjCmjm/xnkEwMqxxxTQBbVNh
3Pr2jVoCT7SWGSVDA5IAd8WoqngwDvFAcH+i4PTbQNr47GSV7MVONOZLvdzv
KKH4+e0rPi9kaFBYoqBNNMW+zWG7qmeTEObgbbsQNpJNhwORJCPD/lLxHgVQ
rVw9qzTsPsWsdOQ3URMTWZLnlX6JT/XB9/f9otogUYEGFL8IuBacBQjLeY4T
CcTOeb9w9L5uxDXruX0MEsJkSnu+j0wPaGif6B0o/UKbHuRFMONpXMwnnqIc
iU1A3Dnq42U4cy8Q7KZh4NjVWB6tg9R4Mg7mTGz/1hfbhq8+QXK2OBTiWuLa
Ttsaur7/oKhV3MEiLaTC0Q4sF7Qdx+i/AMBtdHdX2tK6nmhhzOo9P6t0dmup
71AH6LbvKzk/DtfFjy2MxZ7FCVGhDd0UpihJp5JUWSRKKo0QMzlYEM3+mxzd
0a0deNxnKEHvHQPQbD5ZPr6ghI1Hz+sMnJciAPTOmG0iLz4iU8kMLcDnI2IZ
5ALxBdFdcTaF2QY0n2OoQ2Ef2yfKkdcsE8D6lGdkKjDckedIq2zkEkEMqNVG
ERFVaVwGnJownLmdY2pvimruIEE4r7jC7NvmGMU/M97TWh1HrvnSKLd8w2K8
9Yc6aqCKv/m7gD2RdM2xtUWAtu4hxopyrKLQmHLraaX8Jf9pvgrbQFOzNkoz
BxumIFskFO3sd4PBLmFpbBatVp7OA6+WtzGO8EcFbyR3RiAalcSrbkts9bCL
A2iqkmnXI0jd2ozY1a8/tGtuLtR5gcp7HYCcqIjtBpv5EWvEJlujCt4Zwmxr
5hRQ60f1ZiqT7yD+Y77l57S8LFTTG2FWU26V5ClDVo9ag5gEMidnJ43AjLg6
v4tCIPlQ9wueuH2+VHL4wN9EwQ6YsCxkaBedfsLJKiuJlOkXwY7JN7E1ePgx
yhGEjZDhvZooeGTTcJPzNwQXx2Bs7e4jOSkhrx2+nDmCCR4pYayVogt+eUR8
GDrl4aCjgIbZ6NmYwuecs7sTRuzeII9MemhXfGcSX1gylgKET5cclQrSzSbR
ZGBMWq2q8FhQ838ntXmPAMjJG0pOXspxwr8nMeTE3Rx6RzKq+lbTPELPqE0T
S1LzYIRj/surIQ0SLSmg/IxQ8PVbZP/ZrL865kPT7Kx1rSnDHIai/DyuFbZ0
fTpoFYdmLg1KHlb+r92ZnhfX0UaYnuUjN6HY2loAHpr/VoBcK1e9QvKRagHh
tG8KkZGO5jdxZ0mMEu56v1JYNu9adqAToJQwY2jn2I7jrYYHMsNayigPLsts
3WSAm73wEz26zP83Y+9UJzObDew/NY4DCUEHJ551PaL/VdwDQ48uC1NQwkWR
dOv879j8fVXVIHuxgjj4Kb4zqI+q4+duNrsMWIhDEVIwxLHBAdGKh9ZXlSvA
zV2UoOZOxgDDKeLerGSIxI3bM3QA+2NdE+f5drQ5SnaEQYg4qWYcJ4QM/z4x
vk28CnYnytDN1DoD0ME9Wuw1zLwR2ksXPTVCOQQ46jdjcGVYUl5wN3EUTfLY
BxMK32KigrTo7yu8DngRnW32aDrffKgnQoIIgRGTPNsIsh0h7Cg+BlYTQhwD
CuvwqWMlirecu+3KhYQoAWY4XqQYKY4wm5X2X8yZuYFtTV4CgP6QfiQUiSvO
O9QXmLFeJPcdguCUZ/MTBZx/tt/CPFLbjlMUjzYKaJ65W12ixsPtBMZnbJFe
ICQchCw+LVfeXaEYYRNubUkNKAm9p/RpI1L6Kfp2xsnk/F6JgU3NV7jnUAAM
avZ6EZTY8VAhLUiXoidDOAKX5nOF79QiyH0A0fMlcQzgmzQADcfHhtOpqE0s
ahfohi75YDHEh9hpK/w6fHT/Cx2LC7kd5dmZNwP8ZR99XC0Xke1OqGJSKOD4
4GlkrgjH+VJKg0muHpSel9uvCzQZQvtMbG1P6nAkttwTEovawWMJ88UO0JS/
W6rFQUr5KJZzXv4lmx/PfNklyHieAKXS8jKu/Pp5BNPgnj/LPP80rbZHFtMO
sLPZ0/BXfNXdcNQWRbVlCTjGhi1UTbBzGIZ04JKhfwu7rsLbkY4A5z4wyqoZ
WZRv7JjAlz+UxAKM7aGO3h59AwiVRxvbhlg3fTnMNECSDeGE7wq719dGPFZW
wKK3NGlzPXJn+h4slY3McOFa+MF+h17XuLBYBrawvelRoJIO/PLOgd38e6ww
XtoykSO8cnsFNgU6fsLgjoyQHBlt4W2gKm3tKaM2R16EbHHNxA0WQrTHTPdp
0hktoccOvpEmdz3Z44IPY6Bwbl2eN27F3WZYp+GsFXs1leFcKdcK8evFjFFr
3cp00lNd9GAVllQHNXg4T5ZUs392VaKIKQ5oBHCcyA/KYaKkx4/K6GS4phFT
8Ca0r/ekhsOYDueDlHf+AzYCr0LIIBtgf4I4551bzSx5lP3+oPBdeCYnP80C
M/nIy4zNT3Pchb0oerGoJ2NwrG3EggzIW14SAfF3qfnPTx9IjXGEVk1MXLbY
4z6Z4CC3CPdONcXUvXLFTfVVk3F+KbAhQKuPIAGL6iZvcdpJ8+9lh6j1p+VS
RvAJ6MT+Z2zBeK6IpIq8ipgvMlpbWkBrux8XvAmzi/NMYA7e9As2OldV4Dji
ebiPEdfot8qDKn08b6pOOjP3cOmJDphl4xj0DdFpjSx3I4O4lExsAAkLlk1M
0yxzPkCblksyv7C1hsWL46ZbllzpV5nFft9qx4/R91zExFa8MRJVovvG/nLG
Ds1QSwm2DcRtmfrSj0JaIJrtQMR2HmOre8lhE6Oy3QHhvCanwIOjd7Y5glEe
YT8G1nBAgH0gBcXYpE9N/uJDIwwMxa4a83Vr+bWQ/X4xUieoK6Mpemsa4x0+
++d+2gVortBho4bsiTi/qDnrS1SlR6T4Psu1mt46K/qhEZz65Zuo9vPI7kVX
Ybv/Go9iukyauqRVUAK7uyviRLOtn2JQn0XI1QedrHSOUlen5Xe3Zkfl7nRD
bEwtFqvJzqUbGr6QXs/WE6VW0NBtFwOcCZn3aaF1AZkDTS+nTjey5cHNkOvE
jzLGU2XrUksepScYxsjs4o0ghpz/YgP74eNoOC4J6TVrlPkDfY/RwvEgKyZ0
1uw2uIl55eL7nDlQiUMENkif/fmCsYoMg/yoZrSncR6oJI9Ka3c1Wz2HGZk5
KDwnkaWq3BezRrbyl37AGr7IsjqZloLjDUAhDrbhjz44t7gQ2bQemKTFtR26
Ch1SZVuwXUhuCGPvuk8LEcYFG1/UnOYO2xg2CZULuQ9eqRGAEyHpNatq3ts+
16uzNjaM3bCwqvDZT7Apx0L+XPoAjCW1Tb6zS5YgNkFMJqXwNt8innsIAZ5z
vfd+puVVLuou+16QWEUx79XMXsRH3Sp5vQC4vUGAozkQy8/KR09OrcbJqIkZ
4T/voUlMfN9MNMAkhFlgry0I0zg9tV3QSgirRrS+1AFaKVA3AanrKg+WAMnD
/bQajIOXbK+DuY5tSjwGJjq89fosD1Y6Z7Mz0t2saZsZ7+7tFnazxcUf/AfX
8dBxUYDsLupPZAgJiYjHAkXZtblGg59bXKRneApwbgxM0guPoEpuDsGpcSxu
h9dkyGiPmcQIUeLGKh1WY4CCLlb/2k0TB+/aPYBDYmrMTcLC5MA1gzh8Xcy9
kPVlh2zheB2aHlCDmcDbo9fEwLrO9fnPBygeC/XgjQjJBVLBGybhv18ScaY8
lQ7LDuXefWazVqVQriTOLnbWl3O9DiZa1jB6g9B3U/2JH5xT+8Hnt5ziA44M
9xQ+ZVfKmq2QwGykxQkCRuh+84uETwF+UGBrgqMFS6xGtALiYzuFN+X1PBxP
KPELo0LTGx1zmpd7on9RLMTE57rju3mjffRRCx9FZhFmbVavp0E17S9XeRjJ
/u6zjrqErBdLFTT7wWTBUeVjAB6JdRi9Xei1vr9hhdSh1R3nBVKcIrrHyV9a
/q9FBmgBFeFv4nGKb99uDw3jNr7H0vFwYEgAlGXBudhV7YkwlUM89QIynLHO
W/Il0lbyWTfkK7sheX5jsYe0gnqU/3P4PnMwIO/YmLujIlHuVc7X9MeMEofu
is5fBKsKFtPrqspR6MrA2/mG9wGozQo6fPt4ynKGMhDGD+NTT3+QZzlzwZH+
STk2GAmYjO/i/jAu/Oxke+u5/A9FnE6Vq7D2RTog4V9hGsfFWQJeH2fSSE68
m9qjMjFbJkaK96jm5JnoCsr+UmB6Qv+iPXk470PRPmxLeblMCwoTgVFBauHg
PMhS+SUHl9wYZuxxeJhH04BHefXEha+ac6oc9unJS1bAg8MUHuVj3pRz7a9f
eWDysMFJumhJHT9BW1ZycdoDhUIycVqYaTWViLnYLkrUesncVTgGWKSDPzLh
EtjcA18MpoJbKB5s6ofqH376/vHprHc6oxq4OZXxfYcWT0LZQiuvYMl28ucS
6rj9HXf5ax42c4AIYqFbWSlBjfc3hZ5zFlkNdRazjkhMgKaXxsRwMikzj7tB
Eem/tGjjPPlOb6TpLMBlGBdMDSioUUNwAOOH6yKmeEdWM+8umABHwNDZF4XC
w2RoF5oykCbL4KWnrbYap3QCyFsSaUxMpzwP3OjnKlS9fLcvVQDKOlqYR3rF
RvmSaD88lClX6KgjuU4m3Vp7mUSFKJucG92Ee8/vMNRXJBqXytxdi1Vc0h+y
HEHyKt6AJX/5rmwKxrEvIk4kp0BUXuSv36ANDrJbeY35TzOipspcvufcvL1N
q4ocW7cA96FS6gZd6uY/SySXfBP3zY9mWJS92jkIa234RNbKkAxikV0co+Zk
TcioFnWCo922PYUNixK6SNM7W1tQEdFyxauVrXWnFI4dITboRH2vQMonQ1qy
6jDA99+XI9Y/iG9dY9G2PabZ3L8M1li0Xytc9PmqwMlbx4Iao2o3TKrKBubv
x8t4XQW/vrsLYoENDCqAddIXwLCLe/NUgOoLi6ed66wYYC84d7eNuEnfHW19
MywxL79Lc8eS+bWRXIRgW0+TyeX7DVXw5prJNwxpDZEm4JQYL1nL0dCd02S4
PC18F7Ph6h48qGDRRQQbV4umctO1WzWexfguDCEkv34vnORBaoXjM4IHMrSe
o6f0XHLhqP6v4tPGkd5QXBWa1FHc2TYTR4ez7zrAVKAXEaMUlDY+LxDQ2dIY
hFSv411BqPr/wsh7SVV8EKYx5HvY03xsMdM/4dkfRtkER75wCSeXKsbwW+ga
GjOalb1ORnpA4PfPzOfkNAxnqzo99Hka6rOFkb+O0GbePNHEn1htRdyNWJaC
saQX8JApLFlKTsQttw6GhmMbvtTUD4dFDlYJVwDuRpHAix07XH2JuuntfaiK
ewUf/f2MzPB7clgUacemaHlkgFRJI24WrmIeg3anXge05iY3+A175YeJvhuj
Be+w829Uj39NVIixUBDYfgjdp12O74uEYvtZ8tPnJDY5eMQ/oq1NFbjtGUmZ
mJ8R5eJz4lM0q6GWSbChws0gekfvxLUFlCeUdK0IejgAJ0d1iA7/giPRnNih
5abZoz4u1QrasojHtf0IEU6RMaAh/kcMXfcZylnPN8l+qsUYJdewtubh6fCk
rv9xhdHRggi/y7FyN17pOk9gyg213wQ0rJx7gGH33UzEMreCQmjIqDFylucV
4YEJUUSM5iidkupS4tBTb12QW/sdrgZMzS1cdGTVu0AT1l3nDOvq1ycdevd7
M8awZZKnymcrJO8bS3vWD1kJ8XmC/o08GgsVNXLC27mlP9UPmByn5lj5+w1z
yc+tH5umyh5Lf/lDBlMK8Tx7i1k6AQcC4663UfTypPVgzpCLH5S4biiFTPJb
5f2TP3qRjjJUtP54es6M5igubXPYrjEhgdduKw4x4zhDnm6HmXCnB12hPkXv
iHfQ7PXa9wrz8vt5WXWzYj0EdxWycWxmDnX6DmJKbea4RQqP8LqLfyTd/11B
+V4P4dc5fE9bdFgid9NkpMGsqUjJMf/OgDIEPtwGFDIjgxZGU1Cw16qasmJ6
H9POYH6Y3N61gQXAziGlVBEN/tM4oVP5d7qYt1TBuNFNLEKoTdsPw5QNg2ZR
Y/sGRSr4kFySgUUYJiQKpTGrQGi/OqJ8DbmBlEdm2epURc4kt6kWcL1x9IZH
iuIRXf85qBhRPcKEtIXXPux4rvArsBJqffp4CXjp8Uvasr/vDt5kwI4jZ7uh
9ajbGN1h0CXiJLtOmj6BSgSb7mQraPHfkslwrgNhrL3X4U1zPK1pFT15IpvL
8KQpgjOVweD+VsMHMuzSdeKfZD/+zJTFqjlBkVnBVZsDu8EkOwHRFotr0dLa
wt+XDRJyHNJUtp+3PKm24QJEmsEg26QRTEd1s6JE1RSmdhMoLf24O/+THoHS
dq2yrO+r96PFoxkLLBppPCcq+yTZgZCfBc00vIGmVqNLF1JPF53e043E/xMn
lASdkrKiNf5ZcA7NXItyVw8dj+xlrh4kb1yM6l7qCcldi0ha6ozwRnjkOFc/
TP8jac/yajtOs6oqez0Dyf4fpoTUFZdSk8oSvxQwsZVC0ay4sb9UzT1NHlcl
1Gx51hiDIlvz4CgNZKmUphWOHd/Kl20p6B2Xwdgp+Wu//JCRz1KMO4pnuc9M
PNLWUUm0yXnYux+nQSDfLzvhl9LS1vnnrMHLssc2iDbrO/ZMUE5pkaePLbkj
kG1dxjnGJSRAp/BXZajEWgUgbguuCm5PwA6vWf+2qvXm8W8ocuzEr37Mlrva
inWKeRrLq6xhNI7pISM+jB2CTyq0Xc2CnsN7sin6VdxD9j22vRTGy+XelyXS
gTPslgPzLl7jJZ1mHuCGMyTy37nLeUb6QfgO9zMTzinJs3nu/dZDolP16LYo
CSnt4EkKcoacVLibz7oBikFBf85h9W1pg7osja5NzjGlVZex4OEGSO7PQJuZ
H8Lf+grjMt2H8+6tvMsrtnEwphAT6fYm4MNhT5ISveEWiXfCzzcYyyIjBTWh
v2cvzrFsriQ5cYvUUJw593vn0upGDUJViwtxyAoiULNREZEQVUK4Q3CrDusv
63Tb+Gy6i3GQqBq3enTN3YLqr9losrDPnx3gRNv4e1H76Z1OHaLbOHL4dAH7
1vc+CpvqqiWtqeuO13BlWa99L6decRVpSvJHlvDvTReRwItXOY4X7NnDe1Tt
xILQ/RGAf0D9aAsKTidKtjAM0YoXmm7zhgwgH4YJ9ovv+aLQ5DQgIxXkd6HX
j+HTrdJqXIfEB5S1mmqlAgkLelb54uuRjN/FUJgK/wn8KZGm61f6IezF3BIv
+zdT8LtQEfl6d65tgm6NLbwuThRxqMJLY8ZM0QEYAycASnoFseV2NM1xhGDW
7SBG4DSD23F0x8FjEgMVMrr6VruyWVzDqg7sQ16wzwDMm0tCC3Fd3s7v5zZ6
ebmAXX4g9A2b+A7iaRYrD1M6+R4M+GD86co+B80cRFtTbsIqYktFv2F8LQws
PBY9I/ozv00kq/zvPqGAM4HE088ukhCx3GCkmwDX3XnJpgPn2ISOoVTdke9G
Y1kKsl7CK0HgHvWNIFmU3dOjcC5HLraWwC2w3vSwZYkxeKJ26x3hCxKjQ1Hl
vdNwj9Rr9YkG4C3dxu99gKvq/jtOLebZ0/0NC891vf/A4fxd8jB/7H3f5esd
gbtEvY3FEOhk0GQoQxID85jW8DkVUxVCZMwxZBMNjdjbhR/RK7BnHCCnV1/q
CId27dH7RNTza2nLd+runkRYE6/QnVxrqTAn1rQQdURhCYB6ct/umNw9knzB
KcJf+lJcvVtcbL0FRaBao+tLWZywk4NZgSzcy44otEAXuW/MYzVOOQwYMsPM
cBClZbKzd4QqRftqBgTp47QzdhDYDq8b2bMEX7A9EZMUxdXIwOXgjWHEqDFg
mQzaVXMJlGINoM6XZOj19AXOD5Fm1XkZhB6VILjWXMpeRJSB3jzj0wxOzGgX
gKGwWeCvS+s2oXnHgt0Cet0ahE7u02flLEwFF6RCnIRf62QosylBzWEZKTGQ
S+dotxbwG/KFf1ZCPR3lI6FeeK0iY22YrEbpGMZsv6TwGZdnshKOsyf7Qj/q
bs7Q1Y75B9jTcb/k6MhmLtlzXcUn7IuKg2M8JHbR7FEt4CrKuEE4e7p3WeLc
c6oYLCyx+R6Xd2BwRSaETFTVDuf6LreLqrxYYljjs/NAR3opPT+W0BqChbPG
zaWvKSyDpsXSJPWhLWimICdWftvxtymch/vj4XMjjJhTqDUWoec5mn3d+eme
jNee3uDQMsTWgmqmzNPvtOGCEXsoImlZjtD9fHYlBifi+fcr2WKjC233a6Gc
uKLfaUIvbHsA1ylE2/+7IIFDkcBt/fSGrzhsnF05sdPTgakvQZN6EPijRAj9
u+w0KqI4YXjmMPccG73F3pg/4j/FNBxLO1gQyDst6/LIzngr2/qxkv26JWrX
DB5D31nVYbe++wRFqdR8K+y6VZubjMnSarKo9SSVvfKAcgbzJO/5+XJzoB9F
CFjPmLOrdEyvTjSy84gRB4TgA2f7JeZlaK/tIiwwgNH551EDZkh7rVkaqfKI
86w8Tb4HiakkNepGBMA7SD68yLu7Na522/FvVrcIgaCSqcK/MtdyUj6qKC44
8COopnsGEl1mL653WMqad1Ngq9oJhQNJzRpY6DF9Wl9qG+P+0shFdH0d2WWI
kCCtjSLdwMyOmsGaNTwX2qtIPatzS3ozjJkAw5kUsHDppYo8JAR4Sa3Xt6Bu
MeI1OF7GJjTXuq4LeqSvdAIztACukB9sXaQejdy23zR+DBoyNpTWPbPXiThV
2ritWzRtstvVW9gzyLevWs3H0D39Ewxrozb3OdprwUX9zQoaI7ZuxC3mxJrG
YpjmZa6tiF3t2PNJNLtBwsIt2jdKlIyLAbkfuSFPhrAux5mTiDcjopmixyYr
i6WU4ChPutyG/BgjwkXZYKKB4iFc3Tit3jx34OgSqYwVRpSsRGg9eFAQQG2b
SsMfmGyw2YOFIS3w7BWSs8s+S63xVH/Us9PadmyxbskEiMNnRTVBmyEclPeW
yLIKWMIgeMkHonbhiJplmNdgysJX/LCMr55PQ8DyYfC0Om1XA0t85x19EUbe
Crf7BLt6j3z3CeBWQ16JpUuFZRmZk78rS7yM1gTD9hykFR1dRY4vLQJDjin+
1DnyV6uEZimNuMyoWKpvOx8dMy0a1NMT/k8nlwMsQGekKS48Pnndf1yWHOn+
lUevnavHxxjBp4vIMWSruOjYqTRL94vwLXlUUv7QTnzyGTzZlIspEJCCi+wA
iBvK0YFszvMVVFGcbI76PWMYR5iQMbuDkuQPv+hO+Jo5dS8emF6kMjs717TV
HVlrUQ0qTXWPA2rdqX+Y0NrTwQp5CiS7rpA/SAtaopuhla1XDH9V29zISVOp
3SzV3ENJTEt91FOhS7l290DuNjUOytiBcgspBVG70+eYzLU9FHJZieSZIlgN
WBFGjPoEBw/Ix0KLJ9kJRM0jrko2750z6AsEbJmOQPH1RW2C4SaIIiZw0nuu
ePgcYbEy/atmlUHs1pHRmbEI/D5wE3D52GABiHY0OQ+MBNDTuABXsbu5KyNs
bhIDwPGbbJc90qZw5c9OwnXZuSdhex0e/RIAOkNF/UxU1W9MsExqGgKIYwEy
bndNqIqWjrr3bvy5+Q/v9m9gkxxtpjEdfCIn7wDAEvAe51jR2tvRQFI9k+TI
dkKRgJffcqmwdBybDYwohpaKvUMo4vxr9GVtoBx+Gqvjt0AGzuZl1iFEusjc
6YVZiXOZEG9Mabz5orM154IJfJdpPQruZsPJfgXzU5UiJ6HhJQE+X3cbVS9j
CIk30hpMiXX5ij/Z5LRALoPzSzZFj6gJJHUQuP/FJYsEg3R9XKjRR/nMj7L3
SS++nBJvzgvNk8myAdXgccUXuJkwi8GGLqCux5SVTpFl9CQ6tJqQaQPtBGgH
pmbdcFoXRIAWguya5/80W2RFCkDf71aW2xBGr6xraEu9yJlea9n+BwxYPA56
UtqPXlVUx9ru8u/V6tpFo4RHFAwxgtX1a6A9pDR9HKp76rsuoRZW2jRMlCw1
OPfnhoZ0cAsPSGtfJH7olxLnyZoNdwsW3t6JRon+q4FctckjrUG9NXZAcfVL
CUWvTnjmyT+nu0h8zirZhyjtiCXDejD5nKUX/JdgDsZBfPx1pj4zmuyKkc4K
pV64XjnnoMwsLFWzBM8Y7YEE+D4iY4orOg+i4Nco6BEh76dRuUltzLU3TxbX
I2r26RRUQ3lamVBzP8Hui7/XhKTd523BSja0G3kCwodLoO5lXYFWZZ1DehVu
LPX+W4lPj44uoFwO6o3KVX50Hx08FGD1Mlh+KwLqg3qH9bEJ01NYWCUXPMJC
5M/HRtcsxQGTvKFzWW5euKch7D5CGAr3KYGhA/i9NR3+OIAodxVXI5kb1hux
ViQAFQRY8v9NVG+wMHcChFzarY4DSstb8Ex9yI9y+9jLJYg1jDJHCyGpyqJY
6on2ZQl+kn5AU8u0uuEuLT5r2nJdIV5gdC8nCTbIAayTxqnB6/ZPEyCzlspf
NBljJgrt9j5/ThlIJy4D8LSkZC6uN/0Y03tI3ICHYE/I9FssdmNYVzCDeYOJ
4hjLhPzL8b5ONMwmVTDfuozE4HHPxHgecqy1dNwEVbO/IumhViK6hndaH4jQ
tHUcrwzFmen9rjh5IJ+ZqlJZMB827jqCcL+bi07MSCMBNorqh8RHZu1L5xfc
CMvoxL9zXozfhgaKW1ALavlEAjtuMQwObKJn9ucgjIPDpxmZP86WZfOUVyCO
ERT8IzMMwm8jb+E1V2QIgFQnMAqvLEJ7y1MD5rP1GlA99b4PXETSd2WSZtvS
v3kOU6l4uSFiUyxt61Fu/QG8YKDGtu/NxsmZ07yCSLBK5/oj3juRAdB7ZC4F
D9AmlyZ6K99mDo9Go62b0R3aVXXS+zN3vseVHAisKHg01oxcuae4wJT3gBnH
Em/svQ5c86p2Q6cU2A7v5LdeO8uL1lBRm/Aq7gc9DZA0SzyW5H11VQOEd39n
+//nMTqe09v0bTAG7wW9mHUu45cdTuOnSjwhPHj2WAMa2kKs8cmN0FEaYOba
S5jmDaHinrLk3u0mmgJpo4S/1UEINTRp9Kh12To/ZUNfQn8dDUDIW14wFj+J
DXwtO+adP6g90LIebHyW38cKC1k3tr+esm2e8RlxnldtsKpsTSJxZYpsOwXM
E9RRUlBWDzs22vX3kHUpqTiv6To9hNzd8CrJwzw0M16dGsBzmDc/7gVZvZDp
9rj8RpbV0l77EsffNhILfzaPvV5Rxw6leSfP0lrq87yvRrYON/ozTGjd8iv9
UGr7AEyOfq4Zbv3tP/xRcn4obkfQqIDw0TG80aj7RZA4lLyiwurXESky2LET
T9Y99iE+PHd2XbYWlAjoiOSwzo+cwfeqo5uiPrFxh3vnzaQIc/yLBtDJBqAX
IeDpnK9sov8Vm49GsMxq+YMYrRfzxKfGCcJDw5Qty49Rei6YuY6rdWAi+PZe
If+sM9KcLbfU4/6nqFtR79zzjN6oNhm6j/HKv1RIuYbaGpqBg+cZOlmtIFBm
VclaIZx6QjxaF6qUh2j3XgpyXy7M3vgYCWyPTGUAVaKJ7MK1Lyly6ko1UpZp
Dipg3c8+Z2KZUElPxhVDK4R38+bNJ1S5CRzjjYgh0w5sMlmkMEckp0+ZTBCt
2XFgj6HyRU6H2rbRM76194PL3msOmuafLHFJtpYoGruNCl0j61x3uMQf6YWz
lOdLTsgB4Wou8jTat1iQxbHDtiypMWOuSInvHvlWPxHzSSjIF/RbqLwb6vZ2
DchwSSn+X90l6jsuQbZ8YJNqZqZMTWmgAUZXvYxD4M4Kf6KS/DM7RpFAg78l
W5WNzbU6MP0pObAHdyOOigaeb+s8wMM7LyTi4f0QLu9DdZshZqE8clnmHE47
e+SBYjkIuh+ZPvBaTuLyK2lHnqM505GXqsernygP34u19X4xGEex6WvWtb8h
oBwwMD7+UT2xsCSUvAczxQuykvJVUgx6G5i6uN6geEQaR0YJxhA+ZwzdZTji
Y7Dx5hyE4P0uTTriXq1aYwNEdaSFZFLMmHGu+Ij1z/txhgi6Fv1OTzT88Obi
5eUPzOrfZZNc/6CJTKPsO85U05UjrwQg5DXse4ODTRpsU+ea0fBpMH8Th9cr
hzYwOXHq+lCfpjK+7QzfkgSVEy8jZqyC4CbUH4CEW4szMg/EsavqTjHwoQZL
4ZTupC80cvjB17I4YUGyIlKEwRvNsBu8Wk2EYXJ/SEnxFqZMhUE8piN5n1Mv
UBMq6S3YfRCziSBtLvcF+sOeQK2t3+D3Fg9VNyiTiHK7en29yv1qMXoTZjZ6
gK547UotoglRxefP1kVQMnczvc76+24E4X6AhUCKL4wZkyFkuy/YlP2lQ8Oa
OsXdVkpd2F0Eyari3QZ6Xb9OR6G+btlqb/B0hLNFGnGdAGXq7ATg2ZMJCk2q
17FQq3QA+NfpcE1w/myIHUv557uh26G6JFpaEKVkayUVShGCB+2YFkCE06eQ
IH1InNM5hMYXr/OyjV/45DvtkOFfwaEwDKdyCIXinyrMxgvZt1ATUa5+W8u/
fV6nEK4X87UcEBnxr78R01lBaEfjiQ7iab7AlfidW3cFOxtUu4JCHyoHNR7r
aukTzLSu/jthMk303mUj

`pragma protect end_protected
