// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
yry2K0XnaNsRuXiG5tmT8Epzbp9ILRVfcvSxexgrh78a6v/HQWRLKVpfcxE8
g0766lIS6PuDIPwcFWl7bvQamG3RuUlw75QsrbcW8dQl5+EyUgTJwAL1im0n
kyhd3U7RukbPHwu2577G7xJEMliqiy8o+FNgzEnxavTs0Vsn+jM0ZP8B7ija
HvoL4W/1BKjUqwiKw3sOmCG4G+bFc4RsZQs1YNNOr+DT5M4la9I7GI/Wq1B1
7sn5Wdj9Cbdlxcey9bQcof+ly+OZKrKGHFPdjstIZTzA3BkC1Ck8ZqaHS9re
hf4ASoz54Pzw5Y67ylr2PG+BNd58YAYaAUqtqfo+GQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KCaFzMBSpJ6UdMnm1c1s+wBV2hzd/kuBzEAhp73bZgMFSf++kVijnBUlo3Ob
kXenM5naMEEJL7iz4B2S1uZDDjmsEAAa9YJ4+Y5IerYF1Sb6evlvVs8XQpDe
IVQl67mKocHpgYG4e6QZski5dPm3OuNWvVRI3lmJt/bfUoeGL7gfPjwr7qLn
76mSMYvfwRYCSkXhJ9kRrkdS7MVu7IiXKahv2FRjkIfPyt224Z7H10wAFgVk
S4GtW6M5Mjc+Xeoyhg2JD9mVWBIe1gCFnEVBj93cp7uVkeycOWOnReTCph39
aWd7DzMsja4hl2W0clRjIVx8YM93doqJZW/UircycA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HQ9kQbwXsKtBcR05mNpV9LGaeZpUZ3ddMD6MgxwnXydHbRUqNEbkGs1xCe+I
rOIyF6jB9pejfChdMu9Gioorvw/j3xWN+WEaksfU+XsqTK/9GMgg5gV/J9k5
rt+pUxPBT7pPdwnagugz+NnkcrcBJCVx+OTL10nqZeVo5c4QPL0XbweQ+4nI
KSWfHdRmX9wb385At3IMkAFrf30M16+sJgGW5nb9IJFXwb3Hy2FPxAZG6F6N
SIc96Hsy3H3mI38ci6uu0Py2KLyerZFw3M94xIZavRF5vPa4zpiArfuxA4h9
UDEjn3VOh22lV5p7dQJugkFtM9eAbqmtQq2YoBlK9w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
S9y3xqZ+OpQATh6mRPowFR6L2tJk9ywBmRaXX4Y8LrQPgMFDcTYbOd2gpfZM
aXlCUsK5VzBhlDWK2dq4XfUrGdFtRTcZ37pSCjGGr1SJN8M398fhbL/nn9WP
YzOuP+g+caCTzHZP864CnvV6iL4EtDWH62G+xM+qJxgaQQOjNcM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
S01ZeY7cl4zUq4UBz3pKomk842dzvUD8tZQAk/8XdY3YmwZalc2ObdiHqipW
tmqsQOvGoIOE+mJOe2BpY2h39vj2h93f3rByk1U7TemAqb/KWWxu12ICbjnv
4Y+T0uUy24XelsyZ/R2cABOcg21swR5uzhH61fpkLkEyA0gdac7mbcQAfOUo
3gufWR7P5scvfF3zLNmjOmoHtV2PbLMp7r2G8xXmMVBruwjlvyFkZAfmfdE9
tDTFAbHyuX8YN34a8YSfmBPt8bKMsLgngprEVePFk5Eaa3pVnEK9rkDNrTme
6AvFlYsfn+ZqW8sT/wNKVpVA66QRYCiB87Xv7L0K5UnKx/3JlyBlcdb51teN
2Hv0cI0gLIwHcFtMncXG39PvDqcBnzoyuHEzpjeJU91uGnAjwTvjFlj1vbxQ
IJ9ONQ87AFz4ZGGZQ1nUAMBR0pxFBV2Cig0J7BHKZ2QcFo3GZyEPlV3/m02h
qfy5NO/8DWiHAPDjK+SbUfiObs3WB4Bs


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PFND4vrh8DMSGc4S4PKhfylr7ogjTv9vgsGFHWS46G9SFOkS+Yx1LFs3R6uD
75/sRQ/bHZNsFFKGlaewlDlnjV/HFA3tacE0CVN//SfreeURdFrOZfB2JxQz
RB1JrfHkaPqfN8FZkafBbfilCWoyIxnZ9NTzgEipF61zoA9YufI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jQVZC1TMjTYvMpQmad1cVAvDE9HNZFJqe8e5ouThzPXRiZnVMDh6uVQlPAsd
2+lYsUOu3YVNQiCj2nEMvUmXvhFeLWKNd+8+GTQqmUXIuw+zwKFWDusvd3R6
eA3VmntaVQBvpDaT3u5TopAzMmJ0albXj+gZ7r10vabAgAfB1fA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 25760)
`pragma protect data_block
CTO8Nogloskz9hbYKmbe1FhFglJHndwaJZvs77EmNUtwsAD9qdcMYHUY1a8a
TaWEM5VjgKJ1+lo4YGueG7obUgVIQJgT9CTm62bGDsEEi5Ca64BK0y9+8wS1
8BJva6geZMo5MOBnokbkZB5FCzwgb8ec9FC80gFrxLNBYkYsgpCkD0p8fxmR
ppVnJ4ZFW3pRIHrBATd9Pi7oCiNsnZgUypszGygzDdW4JwhF5FZxNeube1cF
edog3beI9xiKMEQ7Owl0g/21tB4++uPDCHAi3jn0+7Fon47HKdxKD+ZNfu7d
g6sOFRbnH1Ags+zTDGOlWkhpO3PKKu2OXs6jYp6psbZjrspHFtUUvsLp24ao
a00tMQMIGJFLW0xkENrx9Puo7ylUuuD8m1CMeXYq4+FZ3zGK9n15sfRs6S+J
Hrk9jQH3ESeSGwISkqQW6D06nWUOzGNP8AbiWpFWWD0vMdz5NSgLaKY1GNa2
MyG7a7N4RYmKUFG8ORJClAfGMDT7I/bxpjIytzFewSVdgvYph5srTBfvuIMx
qRjdcRGrRSIHgvagPU2j92mnyXuL0ojMEopNxicQEn13cbAZwLvDSpRNZmBB
6kQ5d521pjqMT/48Y2GppezQ9FNrr8tbPQnOCnMCApr6A90OnHzZAIwbEBG9
+Zw6MHmAJd817+2dJ7ix3YOTfKUJgc1GDwbQCLuWyXAUUa7MsD6/7H0pnEKo
a6FAY5vB3Q6EF510dsP+KD8UMfwvEkTRPdDOfbNbgIWBjsV/eVP9FYBfoAYI
r3U2/ZJ1Ej6rOJhazWUMkuMuojpew/HyDokNi+JyLRz0EC2NYU4SI2dfzz5m
RbvksTHea6ADaCduWZdUYavoHQfvHPXIiV0PNLs/sMutIryReBAw9dk157/F
lpz2z8I/5n8nwMxbG9bc6VSeSd300HIvDGlOeKkV6vrzYdQmDcEETnvupl6K
nlEqgdxfIN8nHFR0CGV5ihwJZLbg7crAT0cCHhFR3mm2Obvgb7vtq+PaMc4N
TZuXI1RHRX3tGg3ZmD3UOLuSDEjJPf0qAfuB0RngYza3KFu2sntXnKnAJqcq
a1rQjVyI6LWgjIs8KVz3mfhIYfqUPyfiALqugd28Pd8yq7adsUUfGkauZfWq
S4so1bKtQqzQmBx8XdoxENAXbK8tsMbxHyXg/P0+hruUxWWkrFR8kvvNlU8S
gR9w650dgq4+ty1PsaiQGiJ+HBYRFa9409k1YNkp1kddL09c4tzmaBdzrrwD
SVf0AKCoSVpz1HHWlOCwPI4n2dFTArDgDJAF0vvjTI6XZdf3FAeqGPXEsG7u
AxVWYZyNWt3cn/+jNVtWUoB2uPBJaK31ncZSTucRyr+A1rYEuIIgd3tVgslM
HM+w0LQQc4l9CnfzKB8r0QdxVOFFLwQBPjMUR1pO3F+gqt7oWLCTQX1iG0mI
MGvRbTjxYO9h475JljD8ZP01fRAf8AqhrSq16q/qzbsjKIiU17IdY3UaI+0J
MotZ7Om9PixXvOib3be1OtfEz6yicFRs4UFdwsVhqJKZ/cqw1vv1i6uvl8lo
4DgBKZZSt6Jzy5m3DavILxGY47RJCoszW1ta+01BGbWBjrWk/OVQPab5UXNk
Gr7ettXFAHWjTLmA/TnCiEWgqDxPnfQAYXaYtoMxT4Fr7/MlRXsYW0VriPgi
xCcF/V6EZ1bm8vnf3GekG1we3eDEidaVsyIhXRPUgCNjvkSyN7VJQvaWYUvv
2Stom6Xq0faEMHLc35XVdukWUaCLeFmUD/QR+pVKon8LIWR46Zgi0vKVciWW
sX8M9Zc9AVwsSlJTMszzXVijReX13+1+EJ6FJMN3KE7VPLcc9kQCVooWHwYt
z2KSVWPtsjwVWzxCVwhIznqISIUawmRCKRlc1AaOWYDEt7UMHCoJNQbULT61
vK65FTvXcvE0cO0HNveWRT7xs+jOhMf0iVtICP/uXq+54M9/utPDb9vDXwhK
jVTJ3oDMrf/Mum/VikxeS2/yQCB+NDdCzN6CFmO403HB/s/4PZQ/aiLITBB6
suRyOXuX2T7TD3I/VYoAhJA2Fphk9Ld5w4iavZuo1MrXoSAomAHRNJbbN8Zk
AtU0Zy55/JGakfu/L4NhQY6Iik2dLN9KjnLpt6MQrAMKEDu3PwDORBFfZrJa
9l6Xny/O484g0hdI7qa4jcidT7V+ydx1Fn3ii9e8he8JgDDWt6A751/kaS2i
k9X8dIFyQeWGhANBJpidv8Ghc4YZZxUY88zfKwj3lnE1co2Y0wNtndQXtMnZ
heLWgygVBBI00cN4J+fetTS428+UPDyX166Rj5gs4LHpajSTs11W3vyoH5Gq
w9iTOH9ftVmX/W1wLvBCYzxd5wvly7ej6BiMcMmVpGiNq9qfrNFawEWdMwkn
5xZ8JJ7OmHbLljb9P05rrisAsOKbjm7NlhezWIrol815UO3aUzmjv5GiXpC9
LazNzT8faKg6O+Wp35r3A33GU6zIX1jLuzhRM7nyOgbiaG1bxL/elZizgUjy
40XApFI9gxMRVeQ++l6ldZ+TInvw1cs9sk4ke0xYnqZKw2EZ7WRP1EAGzMtY
ADBQwIM3PxZBzTt3vuYwvuzIM8bIIHdU3OnjrdPt/sSOQkN+Uva5Ze/pUesC
HnijvWIbdtfo0kjzXhw9M1h8NBLBTzVmiHeP98d9L0HJjTmYoMHmnbBGIX5Y
aPvgTc0gFL+4OKKtURlSro3ise0/30MzJUtYqS+hdG+prASzNGLEfeK5qU/Y
q9r3uBZ4oYrFCbqH9kBuTeNvTDk4Z2i9uZlxsFKteiaE51vk9GpPN4EnsCfi
DVid/4qKITb3zmn5efVj9nhTMNzJcUs/WOH3kHucZHf334GpST/gTuDpRG6X
QZKYo0bSNKUqXSqDBfEGkAhBnstaJGNaFDzscd5kHvitaDTKXzEnNrWd2bKk
3f3Cz7qDNf53v+uKqfPN7zIBKoZVTh/9NTacIGFsd3wC1YdBNsz9PpCveps6
NUkfIuOP9FazcAdH66AIcnn4+ClrZ9x7buC8ZEHpzFb7HdmCHvcQ6Vxf+Uhf
rQwBJi1hwDBc31srqX40sOcKYHrTwmTVuk6y9DuVLtCJFcpqszUFRyYYy3Uj
A2tAs+wmf4nckWfATFpeXYOLMkTAqkd4gdNOwSRZeHgY3ojczcb4KJFJrz5m
lLjDvAREfnHHZ4KoGs6zx0MUm0LpVhF91kYV+/QCA7wJyhXT7IgZzQeVPIOz
tW2oxR84jmdESeapDqgLyIjLCE2yM0+Sif/YHN1sk4S8zJf1uF0ajDB7oV+H
BBtLil3i5DbQc2TML0QC350A9DpwcwdVBfyukz8ZKS2Dns6f9/YZ+FBxsaJ8
M2Q3MmCC9re75W4HZpJGhep/3TSx710DTGc9+MuVLgy/aBw5+uRnEwQc6gle
NE6dHvB3r+WUiYh06rylFh4rloBXjjiRjOoHPHPLG0nk+FV0vHkrCSF3Vrmx
//KiGZxu2u8cq3LE4trZgiGhrLGOSovRv0bi0Cqj/gXdNwoH3xgx2j4AkmXc
07BIwTh+teC77unf3VXr255oY8keEVIFcRpRsAZRz3s0mzptjo1WnQva2OpN
6FqLQ1S3i4ho8LBwpun8vG/5p5uq51qCoEUBGgotsrHMSucJVxsXMzlpwTTk
gjtYa2sEgDJC2Ml1OLh9DfIeQXzM1yg0V4ZQypGqfw7vGn7JJUtfw7DWsxsw
1Olrh07Gl1mckiT+oWjB7LZbThGfscfzNee3vhMUvErhgmvU6EBcpa0KcYsc
JQqUeMenHnGR4+hL6xhs1jtHWEePp8aD2PKv9rh1IRohEoG6gzvo8z9XRNhx
FWm5ZuRjkAAyfqB7oKFXtMrTrV2nzTzfRUk2gNX6E+LK1IKkB7GbR6hXT4y4
fclbPkXZ9aqvFEMqKtXZUEOXEhhTyFVgoliwkljcYpD1sCcR79HSv52UuL9z
nq265dzTmEZpJYc0ER66WDy06qLXu/bNSdXFC672Cp76McrZSfhvps840ogN
WkQXH9SGjhqLa3kmJnI5RNzqJJ3VHgGeSZg4exay5Y5jpUdXO3fuWxazwfgu
DS5+Kw5V4amRdpWGvuk2B7X9RuOwLaVI6pm9JJOxO45MWjOD98t5u02qZMvM
9k+4r0B7rBf2XEHRbkr5XMTtLiVD+/k7YV4eZvpJrzf6oMXdVcGqF0WVbPjc
lZUFAzn1lZPwzEzdC6OuimiRUe2ff62OH+yB31n0cu9sDcHr/TLIyArTzXRU
pO+0y7+p7X8nhA/1IWqWmoFdx6O+eXIOABPDs1cG4a+zJHdmnURE7jzN/XIm
QPg96V2LeYygvytC+YouV4dPgTuovlAOln4zmnlkGy9DHml/kMHWDT0rIJi4
YgNF6ud+pit2Qu/+qTWUllEevdDOtCkcR4nluRq4vPQWudfnf7VUXa4XBqsn
Hwf6lP71cOsYZOphqUIs+5IULu7UudLecmvP1++jPBX2frSkDAhlFRIR9Yle
vtC0fvOfeCzS24LqXyKZLQRF1glug6nApBZx0HgxzPFlOykOE6sqzf4rdFuf
NKJH5j1mpjTQXQVB3k+Q7+1h4LKqfASPtOJR867xyDGHcmGw+6jf/y8kkZzp
Mi0EKHb9jfC0hsk1Skt43MgZpLicngvyP5WmjLxBX2T4WlbAXVocm7YJgAxH
96yUIH1X0s3XR+T66jcUkZLv1P6ZUUUDsNnTNxwJAKS5u3nMgoEPZqNmxloS
d5xokMpRaxem2RD2bpEYFmcD8it5nFNfJ5TGpHtlJ6rtmLx1izp0P4iKQRjm
19FDo+4mWqLW+h371HJr5T+viYQFd1e7j4S4B5FPcNa04Uq2ZMmYz1PVPrLQ
hyzC9UXVk/ayXcPOHIWDddtGqB5dqrqitZB7Xuk4s9c3hniw//bKMpbtSYLq
xLkzmvnLAAaILy4aMHUh+xE8ZU3wWN1V68ssOFOYLeIknue4zKbn7pV+EUfz
daz5iFbm0uscR9oTLeZAXByPpyxMkBnpWfS7ZWXgUci1KHKmg1jR/iLq9Lan
+H2ns/Xmlcgg1tddgrVpK/NYAvdN4mhp+szC/0ctvfjegDYHTeinTPbjGshG
/5yYUiOzxRVQqUNKY8w7XCFnsRpf0vJ4pxTTJ+MP9AY+57aOoSqVIbgr/HEj
MYg44vZWAJ4tDXYr8efE2UXqiQzNy1w53o9PYegJ/UQenwmovWqkr/A1Amt4
s74aTli5ma3vC45e43pBPLSNnu6DmcshiMN7tGFjn+btA39u4847d6EPgkFW
M7oFV6pMVIUKrYzQBXtIs/X/Gq9StJ2waTHDjXt7q+tXSFvYBunzcjkOdzm9
glzGFuQ0AcEQRptwBHSsr3lkVTG0kNUXsUPFYiPaUuRGXduA+1jYITcwKeO+
VR2ZNyLEkuu0ASKqYT8Pinpam2hb8Hhq9olarjfzzJ9oDWVNgq/n7CSUhjn1
ngePWMF/sT44la7WR0Ayw19W7KHSialybrjD+gCXxDstos66H/A8n21XIDLy
wg2nWezCABeRm+zOQTALQlQoPMyQxSErpj2u2kSnyz+J04aexKpc5OPZkUMP
iSFSA3W8muFuNOaX/K3uBBxtemipb7U4id9UgGOFWNgize8wXZIYKTnyQ98X
gfTzal0uViJi4SggG72DMtHnzzbc9yaGWgSWnU1aVlBu4DQYTqfMgcHHH1YE
47Eeh5PoLJzV2pd650n3pavEGjkvvQVWqp9u6S6Si6/0k+khOzHmOnW66w2L
XDTmFQFi7jKUZWZmQUXEienhZFP5lQvZitFPh4yIREc5j0/9x6elHmRz1E5o
YcvOYkZTx1FbKZr5tfh5LPfviKgOzYiuNTJJf6ZEHN9nillJicB6J1pcdzP6
2CFJhz3CE+sigXd8Gmr2Z0GyJjiSBfgGPuTo0ODJmZP4CBFMA8beLbvDy7vl
J2r+R576seNFRH18ZfA7l1DkzrCYg0zXG8eJ7WQgZ9OPyKqOKNIcmkR3sIbb
Cskf+QlzxWdOcA49DkytLXgwsAXd78ofstJ+JEb67vHzjlOL7vOCOAdg/4cP
sgrV5NDYOzjTucu4ffkZH5CprAB03k24quGb9a1XnN7jygTgPpIQ5FQ2ZTwb
VMPaKNOkFa/+C2Rd6At289QmjRMFivl6O5luYWKn5v/88ngUSAN2z6xAIMns
lKTUrvwacwU/mD46CHOzqbVDi0KE/lvEOKfVOIsARr5pvpFeZZT3nFITVg3e
xGT8SAd3R/69j40UH3/OTMi5tLxWJPmeWQAa65+DMOub6z0bdeLq861k53g9
7T6kb4RqK77TgDX/O9CuUAQF7lm3o2mBr02ccrS9F9E9FmU3WxkdXuZn397X
xMcWq/lToUrq5ipANPiykHq827DYq0DhxMWLLcZZnX5kZBaFoq6yuDDIbK0E
tWj/1rZG8w+G8w7h8KH7LOkqm2t4WgZOZTsaTbrpsWRXyuxfkaaeQuVA8zGB
Hrb0mFbqrC5ASEKyw9rYbMubohf35Xc8p54APBL7i1vG3gKxhmTlyUIGBqmD
fmdMCY7m3VIBmJUYJEvk+wgNEp0Zlp1rdWy9C8h48tEAyT70/tEbRuwtlRvG
lKJR1nWsJFcz6TEFoK3ODWgT3XOL8VC66O4lgtnMHItxX4WCzuShnHo1Vu7m
CE3JDdLuHjW/dbsW/S2DJOx5hgfBmv9Fllmy64qqaZ6pUGBGkMu/sNNJ/EYG
urL2fQ0e+4W5XB5XSG0J0n0CLZi3W91nczrdla1AEKpiybmNAiJQ82XWlRWL
GnT/FoOs9+vyianEWyAVOmMeVIzDBpD9hag/9MnwbC3/88DXRSuIi3Ur75g5
RJWBXM2LKomRvbx3+Vr3bY8+vK1KXzHJU9kWbxUVdkfUrPDVVItKIvOT1PPx
taylcCDlNpahQ9ImgUbPxbpNhS1bLfel3hW5ff9iN2P6p3RrNpGCxrxneE+m
yQIoLx5k5LcLdzNjxTr+Zgczel1uhWKDKHudsroTD+nOdyQEQaAqxqVxcodS
KtWaSKkao/Ndq0D5jrH6R0yUNRWUCEg9LkSnR9blBJqs4dOFvGjc695LtHpd
lKQWpTM9MorgDw3fVt0r7QOHgqFIfjZPeHT8a93zNZWNMOExQfmHqreirJs2
YjjxvxTviJd2QTHjE4Nbd3nb/MiS8I64KasGsl0caSUTul1l1HNMLWP069AI
mIQph1DQRGFrsel9rCr3GmQjDYBxW45qmBH3F7o+fGMeSuYYU0yWX7ERh8sQ
iWoMrBkpXZs6VObM7pANM/VQIhk+4yVoAVQekl7j3yvwyBU315uNhCVHVSk+
elr4BgS6UuluG3ccwGnC6J0Jw9Dysw3VzNqoA/rshl2RSCz18Iy82sA14zC4
yJ9QLsjHWf5hfnEx0oYOisHa0qNFGIya8p2shAC9/LsGLU0i5NOpNqwR9B3v
nO1ewLo449yL2+Zlabei6NeTbiIJZs2fqF8Pisn0Ak/b0/fg+xLmedR9PePb
+oDiP+uOjsVIzTCR6HBFrprHXoGTLU9NMae+BXClVRhYFKcLs0xE0T1Ggp9x
zQ/Q9IWNbJBSL0NGNMrdFPeBb2o9QR7vOLr0xtBGXZCoqj0UB3AApngwr2zU
4r44IdRrBdP7BdkAx9/VObqGN962m40kvzShPDxYT1PVdhsF/SBOjKXuaTnq
HPQwL0D2lE/CJBIDuX/o6vk7dRVRpnw8tfRaIkNpGVhZMfIpY0zQQ+Dq00Sa
70OCSZ2N3m9LEVNUqxZV9cnu8f5fPf2GTUqvzYSpQMlAX+H+0QJeO+JvBb5y
2Vp3HYR/n1deOKvjpuJ+j3aeJauou4qDEzYOXA65uoudbzKaqYQaqhZdsw7P
haullszXCat87navHyPxCgTZn0dLjop1AhBaUKvKx6QguM6OrS8TKWi8vmVL
XUPENLUWXCA/Brjg+M+L+NbGwJA5bGbL58I2myzvhF3ppJ4QLC7IXijgaN4m
UUORZF8lLnqY92JOHX6w0COcxjygCrRQmnanwWP+2PwuOv1f2DdHP2ccwVXD
yCCFH48zczSYHEkc025mjDzhz/hmIuUahmaDBj9EfGm7pefVgY+zj+WwnjNc
sio+bGI2N/55o+vgxSxaQyGdOuvhIAaNU3rFd/wqAWoV5w5VuvqiVZt3PEuq
vT/UQe0Y+CmWwXiZN18uHFNJNE06/EN6wTVCnvUGdjzpOg4iMFAwsaJHG1P6
n2jV/Xpj84RdQ/oNw84wnFnT5jwTBZ3KKo733pmJHFeOOoEh8FNVFGFSzCyj
MmZUKFwO6x7KqtL8gKBh8vIo8ffBagD+wCAhUgqe+yxzgRn8fCxr7ygG9pnA
k8kQRbO5CG2SKK7X5nl1MbtSY926/MKBoNC02CLM+KAflAZdaTcPLks+ZcyC
fTF1CVsrB7FiZyZXXZMz3CJyuzBQMOY4oUgfKwBulddmHmbwmVp3P6CFVqqv
xqJsL7CJYp8SVbzeEXaZw8IJOC35+4AtxQAR994g8r8czLKKb01b8JClBkMj
SsEo0Z9JgISiFnZdWdZarcGxZiovDYFw8l3uJ6rHLh7WwDyLaOib8LrcHm16
PlbrmrpPhDJ6BmNxmGR/R4Su41SMvHlyzW3xr2tKxwh72KU74nPOElj1pmDe
sJ4qMlYzgr8e3FhLxyCGEIO6wI82wp2B/dJSeBHVEMQGMyJ7y7swtdhcy+rk
3fuMylFlXo1jfDwaocOlUvJNI1rtlxUQg+twYaYrf6xB692/Qj7wzYUgsPkp
lfre9E5fwCczYmzVchlcTTPa3cARegxfObdIpH5vq8glCDj+C/gRvg8b7Ojp
amOlW7+5+5bZ0QVS3PcP9g1o6s79x0HbD34k/Bbk1BFNE+pE8ljyNZ3lXLgz
kYQnZf5rdSAtZzhN59cLgBBJhL6/C9dR7SNJ2GhuiFTacr0dbmJcNm2V02et
CkcQYNAnInQ4dc1JoXLezGU0V7DrxXIpb1XaeKufowzLWfJRTWY/8v91LFcU
6Ogugo9CuwlcdJEIp1/YLTtFeK1Co+N3SYX3ueQwD1g9czSVOH/DlYyTp5RF
kweSSzAUSxYHe15lju0vnEFNKjT5h+KAQeVolT5/i5ovwZpx/P+nUf1KYE1W
5e8/uWMf5B2BSx5yVDarjO9t6tpOjBWZi10QvIJpQviw3LCxTr8okXF/lfGC
CjNxHIONfnyzj3Tmn9DsnP16h7Quh2XlqVDv1YotZthaKrz6vV5ww/NwK3ey
9j3S9RF8BKKXUIazz9jppdwuIToSuUgrW0JEonbJacKDGTfdLjcQ7wJ7k8+G
LiOiJbWXKrryhAmnc2mXKa56RupSap6fXrkqfUoZ+kO9nAto4tc9D7ctA0Gv
FHrHdTctBqQoA/fpD2q5I5wt24Dfn4JjB9lCxe2WcvOe+owPMEzWfvQGFSOq
wNvcOnJScbLp0/clL/s/7tMM26gRhqeB/bTyD19iiKFoMifV9k2Qm4FGmEZ9
fDutZQEs3cgLXfSjDP75w/TCAtESMrBCsScW4p26TGwoIAHe5c2A/uXiE099
4ZfTy46lLjsyQwWpxW8VIaxyBqkKYzvJePLItG52ltUns+pJLxNkacBJRnZ4
KLlaNaRVgS3kyCWokZT7QEUHGxyuud99W6J3dtjvaqMmN3jxBAjk+vWnE2ro
LdAk1b64YfDoUfFfh9AxGbbg/cU5Vx/wYF6JM6ASdzEbIdQm9UtIBkjaYtbG
EesmSY9bqzSv0n04bOvCmhscfYZnxfLW8yLomVguZBiKXyeYgXy+P4XDYMT+
3A+/xPK9jBQZyQx7cA7YcXWhu4X7XfINaXqoQWJoHBbTFMSTgiqf0ImMHlhr
2nxORCLa2oErAx0gLsp1Dw/Gacs9Vcg6xYaVLFSZ5kpuj6BAsTLl2+n+OOQr
d7g4khWCJB417vPV+48nK7GEKC0F33duy4F3wjAE+drYkmMeKI4MmwEGFxBP
LPN3tr0v3nb6cNtTiRf+vZhsaq18GADjl9z5+P6vQDeuABVXOMTUPMbBQ4g8
BDg26MGWtjqqwOSQX4XeqYIPJkmzSOPa0x94LGK/8m/HjgXlAbkrogeAWwaH
+/tHC4P7JqZ4RdAstjJ4QdHrnrdM0FU3Y429X7qwY05L9o0p9sVKdClqXiFu
KeBDL7NtbRqF/PzRFU3SYoaOw+6yBJ942WlwE/FRESVKQRuf91DUYsxXRYNz
sxdmpo7kmEEqxqt+YdwexZIWEEOihznUK8kDr73x/lhasXB/UH6iAwKPp926
2JOvjIAGO1R3tX1bcNV6vD4MqDnqzGAcvA0v7OG9GLSvOiCoab4DFIlJIDOF
uq/4TIgG2ARK7up9v2FSTwAxh+cyylBUf5Avw4TC3KMW1NnG6/BA446mi+PZ
jWQlioIN+aeM1H/8LEV8tmSZ0y8sgs6fK1034I7n2Xv2XkrOrB3tf9wnwaiF
XVM3WHgnNoaHv1mZYQdH4BAuDieMUkScTjhckq6B981f9yL7RvbXVMMYVy5y
eefe0IR4tdKNfn4qlzUmRkrHXcLSeNvcGCrd2U/UC5suL2/w+qu/fK3iKdIe
qg2j95LC5TM/MkHFC3v3TMsqIwSEHdYD7siUQguiH/ZASQYRSfpD5pFQLnM5
uTSOu+4D6ipVGd4DLgqbObC8kaf6/yqFoFm7bhiG6+RvY2DUCE7QlQ8OxfXF
f6zpUHgi0pQJUMyxSq+m6ZgKe1rruEoHPCzEuvDpW0Duc9H8wSX8XgOmEAgl
o9Xjhk/ZfM5pck9stQSLJIXAhtX/ohqkKRZnl/id4xD5oQp3wczi2K/6C/6B
YZ7w1q9jzgQ6hWAM/WtyM+gAgbNO2bf3sV2w0EFEFM3GJxF/Y0V93xTywa9r
0/B8vyBYDpb16zWNt/ZSHo5qPoPPNTONxziAbEKkwyFYOkRUkpu2jxJPitOJ
FZBchujxswoO3d6qczAGbJaxtVH4oWd9RJq/x1nDHhgRtOuuSuejBBSqw/da
unqf0ijzTTijqSEF8NGQk6ZkK9pPwMyEyNWCkqHPtkqWw0P74aKXncGWGq1E
AUdg5SvCb5OYG8EoZRStyRloIXQ/9G4oRO1SNrWWptdErr7ZZNMfcQ2Afh/x
9SCs9axM2Qj29Ks6MMGMv+iB/g+0Kmo1IF0fB/Vsgn6QOpqW6C+8aAu4/wwi
ye8Z0QAGK5WSfg7O0tzZGmQgw1AY45WoHNe+d1WjwBrI2+rVLnLR2HkYrWHp
SCeLGJeD1D9BiN/T+oRZdTlAzuzC3fiDSdYepWw2P5pwsvot9xK4oN0OZKm8
xpnVDmko+qn35wzfIwxw7JWSxjsKSu4zf8x/YVeWF75ozBKmPrcNqJbIkYh/
v1MlHorDJDTAc+xT7uuzGk0qCpw0SdcVJSz1smBTKMeZpYOb4fWnEy4IMxEy
FThVuEKWwZz2ysKXlVF4FmrasyrKNU8RuCj1u/bU2XmfvCY4B0l5qrkSp+XW
+H6g7VZ5ekrrZx2hB6RtM6lVBu5bRiFtwK53v61cV17bJXisv6NKvXKRu6hb
Hbj4ZyBICejbUO+AAvzFhpZ65MZ0tVvo/Y/X/iGOUqZYuOVeH2ENNaC1UrWu
p1oWqNgN7fUD0TBBUV3cepoQBvjsJRHY11LY+Qr0yQyJU5xkK21D5pnCRyfA
96pFn3P1kAeq09HB7O1kgt0S8gsx4RacaHJMSbdA1/dedPVfx6AdzZIVqwH2
Mp0ZaHqWOl9xx7owmjQBmqHrbtiwbygJZ0f4wy+XljsXguM6IoOiTttavsHo
26ZsKLNZsNGpZwSyEKuiuNOiQUZay8OTJDo3C+oqLU3MyzeD2KcwLunWcA2X
dl5XDjNE2osgzxhygVomnEXMAQfgmZEV5n8pmC50V5dj4m+MEreNc0gTCWss
T0DJgRZAuwVHuXzXuTJCAo65ZxLlDMJ8MTe3EgXhxI/U1TWlW8D690mHWygy
hLwUNmT+sJRCAE5ypJuEhMz8ZuBlwZtTWEUzNAiNN28xYIQEmRva0zEOg3vF
mx2Z8FuhRLuwyCcH7OKujB7D1AotE3Of4K6abM2HGBmwDOdlrCKLzHqGYcBk
DQdjnHFlGpiZpK5ci2MYJNrcVtcfQ+jpgZXT7PYEqDA2hVff7XoF8RM+jye3
EwtnmSpugJ7WS8yw6vio5AaEPuzaUH4gcOH8oYCApa7Yxoy1ySqWfjfRB94k
+FbEaoq0u47DEAlJl/xZUHGF/SYXOcYSUXFNpnZKqjqO5ICq1+BtbWM0qIcv
oHcLc/QjT+o4AanzKNM/FFGVi/PGNRLJX9bjvmlaSKzJKy27ZWVimabtDkju
H/GARkk6gwnK52Abif1ANmpLpIroyusNa7wwig2k//jta4BKFrEQ0BXwH1nK
N/seUEoNIOuw/qAOgwtwSLXUZG/VuvtoGKE71ptFRSzzj1vPSSqCmnYLqZXn
GfHrrnznfKVZAo6BBFJNSwoX3vSzfDBqobSxJFtLp4I4A94QP2XDmuSSmLPt
d9G9vZlqGKLK6ybNrGK6Nre7qzSif7cTn7Mc3rzdJheJ6D5xYFmqzyBpYyOD
ozrVqpXEM6eXaG80K8Udq9iQGjrOhvEA3sJ3/+cOXaN2oMHLYdsKWKwP3MDa
njn60DaPFmdBSqJdgUZDL2mcYQsXjyot339U4WtAMPhsRfXUYqvpcJhisGvb
9Lync2CoieA1cRM+nuT2z7jZAttl4EOci2SNjrHh9iSQpqWNkpnWeJamoUtO
FfijG/HqeAgaBTF+/zT7OJTxNzFZVRAqzCwBBDNn7xAVo8s0TnAglP/wlse9
6oU5m7O3UgBwG31p4osurAcXKqDWLH/617mj7NYxIDrWShYUDW9w3hPcuo6r
eUBbyC7sGZcTw8vc8HYcyQoWCESWw7MJqohgo8Vn+fhUBWryNB6lL3wEMhQj
Cu9mRM9dEalMjaFzzSiBHxUZWTQocq+un5pcv0xNqZJ9pNiER5V5VeKNuKJS
CRibQn2cLRIuGUpT3Qw7y/dvK5yLVsX+4LeJIULSIFMOx6NFnnVPP1dRtorD
iMTvdgHOJM/ig2DsibKfC/N1xDuZbyGXZJRtr8OOeZYyThKx3opfyIbB55qE
n38iPNpGNvtQF7bfW5fQPYo+rcKY4EQD0EZbUvVz8Bk5VgWmB+p99opEhbyR
i6YI1N0sO9Nq/n8PCt/gg0i3m/Bgu9V10ejRlqap3/PGaaa/ggbpkp2T9RbP
fXo1/ywl5u5AFrL4cY9JAQOPrNYbzt5oMJSk73FKReLwzpWzCIaXSiVEHMG/
0hxJRb6mAaZLixafWgRc3uqICW6qJYAoQvNn9ycQxZE1nD0ROkHAAonaQwy9
lyx1CJCi7iFWnXJxzpRzmM1W6h/vV77en1J4plbgHlPRJ/zrOvX7mox+iaMb
feETa2H7XEw05lCCP66VhOFkV3el56iMGlXg7cxZLTqOImr4RmhOs9loH0Xs
t0DGCZdzLgSpeTnKACsoor2N3SlPHFAKctfVWnoylFwyJ7zngZPOu4jSzUY3
1y7Key7TRR3tNTDjEJ1yYBYZMDpDFZ3ZUMoP8vAnjljBFOPNlZS2VVuktxQW
KhdXaOtraTU3+y02dMkFi2axOybsMC+08C6cxWdUwTNv2Od4FulKypKhhUUc
OM92mqitDrMrufQsWFTJWYYgG/hoTtcaIB5GwVIh07Tvar4K9hfgDYfD2uv+
ZfdkMfZjWKhK11VYJaFSQo3iB8hB8ECT3iFqKScZlSMFBvfIEbIjSP253BS+
2/pcLEUpgacHfwZ2jkr3l5aLCezqJQnOef3MTePGdQrqlZa6Fx8XLPv8z5rt
gFOtLWHaMzDsD55+kS3viIrAdarYC3kEs1ajw3reZdAA4qoTEmv07rL713hP
V+9Ex9d7oZetGvELVuPDs+Sn38FmdJaz4iJF77WTTsLYaNi5cjYh1z2N5t/r
Iku0RZeQNtA/bbvq02zUuJGyAPP3MIFx34E8ey38x9JGq1Vq7w4r4FZKj1zz
Nj1pxEjRDs0gpEU/TUwInjDlqfsOhhFbARq5mhDMGxuBAZPtfWum/b+BvEt0
G/Ni3FnmzR4eMjgSQTDzC+g8/pRHAjYbKI+g3VxpjP2fa2N001rbXDsQZpQT
XFot3noZU5LZH9Nws14S+ZOYFgd5HF8AtvLoSsOfp8yS8akWyJLKEXqi9Z3t
ZTgzcR5oXPfoeKLeTF3A2kOAoTunQQeB+CwzGHub3fZXxGqelnubTF8I5gC4
7fdKFpKuZuwyHN7HW2zTmu5Z6GzRPInU40qO4ufEu+abtRWQa7hvyrcDfgB5
Iy1rOIemoP8deHEaRJ7Q/osB8C8Gf9bWY3vhVB+px/QjKV1v2b1l8GUzR6nF
xJ9bFLzMTx0vhJGYHDX3+i8uFbJsQDNilKo5LUvjdmKrBQLslljyWMLv0pVN
WXNc1jNdbDdzGSkdDSUr/O0J1ybQTLktLxMpd1t3JfiZZszgtduOcYuvcacc
TAi1cVJBDlDL6vr4y1T739Mb7zPOCWRaJQHf4sgpYfMeVszQFf7FHrrWZzUr
QzAkvV6OZyHKp5pqbOBfqequBofAT+QatMkZXn7A0SKlTwJhmAsIYzXM3+yB
zo6qO2W/1tm+YGhC2zh453s5Wm7ATF6vtULbRV8HzwC/oCyLVlo3Jizvje+I
rumRxH6uaSLpzcreM0MNeaIKB1XgBo6RPokHLtDbL+0foU+S7s1jaEirC1ys
qguwUzx0h/sGETztiAXj1j1DrCZZtqq9NmKbfwuXA/bBVOMMQAr3a6R1JoeW
cSc3mWVAgFt3YMJVxTymEoTqO3dTrFEtpR8BzCsuf6EfyYmSSst+g3x0jb3/
4h0McX6KJ32In8GlKWnIv3pm13U98BQichTtGDCBa5C/DFrjA3zgy2KucTrq
G60M/emwrfe2ehQoHWRytIgctURbGGnGOi3KY3vR3qJ9MFK/M1R9BufwFZ5c
H0JvNomD01cEe3VKbdVbybMag0Q4/doM/8elzGAh6Nr17SUs9ecqD++ZyF0L
o6IQ1yrPt4kkdooXr9J0+9mEigPaJWC/0yHHWstHLTmGLG1SniyryJIZZ+7e
WLpEiMuzNjVJwSpziqpGbeJ0WQFlS2BIJdf+8A2zzIZgG6ic+DFwK7t+4+HT
aKkEFKtECn/oZMj/vEr0d/BMK/09VzA4j4TOWr2Fc2sSmEjCWkDFGBpI/8hY
P6dTflAlPSMWgiwDIA1WruWYN1Zj/4FXIdMwuUX7OE6g2TSSRq8XK6NDKJ8u
CxSey7VpEdpVJjhqPAipxIzUmsA9Z0aee8ifxRbrt+Emu4eTbks5GL+1Aqi7
yvImcNlzCO9YPhITSs+wmYTe4Hq2RShI9WWpaClvFSXGifL+UEE3KmI5NRJI
qVrDI8YGbOtLIjnAk46MbRWOekszHo5PMV9vMTAZJPq5gouWSCrDwbTkdkRH
+H1rp//33a+4UxXl+E/nTASVQHk7rUHnBMkkgMhgr2NMW/6j0+gwc0BJDISN
puf5XeJ5kyeMHbl2u2dkHC9mNCWnf+r+dpFlXJ9lu4OrsatdM99O21dFi2IY
2+ti9SCzd5/MthewVhpW6rj8Na1iHW5Ef+BjrTMcpOdWPFaX+IhV9xPkNLO7
KDQ4iYvzkCUkQpUj67oVhIfO7hABrNcxAdFPFmxxqTJP/RDdhE/lwN8gMRW8
/sACBgGtqB8LrQfT9533wDjJ09ErAMuI5Kl9R6e+5c1LSDIJy03HaQ7A6DmU
4cePheEMtKvXVrCPkJlM5V//+gpQlMmCugup+i+ZLJFrvBEsmYnOLxTn/H1p
4RYqQMvgXOiWtOMGC6RNttNrrc6n9gMLS8lmEV/7S3lKA/Avh/Eop/YqLI2V
9XEECqVoiW44keykJ2i7f3kwC+9lL+8gQZKUFKoVdipm5F+d6Q5Z1YskrpU8
nmHI+lyN/Tisl7tnVcCkWrpMaRexlMI1exYYP7p48oeq/lmGmHELLbSEPGBq
bznLBSR3jk1y+ncyWWdWfFtOyU8BIJyo/zFSpCWLi+gOvmXTHJLD+R2FlLWk
KzreVsRKmiIyCMfBarcSrFasTQkmqKd4wk7yR90XxLPPvQzU+DP1/chn/r5M
OSWFzqohX5CDANPcG8pz0/7BBoSTNQ27InswmRQ32GMRaTzdrzo/vaPAGD2n
MoutGDU2Td/A94BoxZX4JNmoenJMbFv0/C/2JOseEy/PDyOlvUxoCXQ4UZB5
WqXxYdniAfEiaGWv28WUfrFfTurBwKU3DTSIhDeth3WqDtrs6vFogTKEESYN
vc4lpDwfwXUN76Qg/ZA7CEPR1i8BSI8yxQa/o/dV+VKGOpUrVmUWtPfbWKyg
SOtZ8D1HTI+0BxPKCiNmz1VYuGHeNJ5e+coNMSYcLaB0qd5OLK2O3S+BGZhX
bpbX2qOrcMRBeGvkbaShMrxBhHa3j5fnckPjFR5J7JKQRXkCy7JjO5HAlEeh
cpahwzInadBnZPzo373EBEw6OyNvUDG+A/drrt9P7SBOS40GNo5hFMfS0TTp
Q7bt5amy1lfwW437bii9+RdT93ykW5PShF1Cvy6KCgof3ae3ZGD0DkTDz9x5
JkuIv8mIGQ3RNye3TXYA/oq/rRi+VEOZofKI26Lgr/rdFFO1ovzIpW6k5D2L
RYULCwAXyAEXME6wrJHINAZYZ/3styVCiAMknbBk7vpWH7s6BNeonqzSePVN
ii1MB2RNqIEGUUGwymIRhKVw3K9O6CvMLvlDOrBkgwHP1kJgv5hKHJc1SDg2
sbdAwEzHR0wxBwj4JRwmJ6yBk3z9W++Wxgi00Pf+aVWyQagxQquLS+h+TN5o
W/4VO1M9TL3MAuNZThsdjlsyKQ93PVeTnl9CuuvOs3soIC43R9dFCQMOqHvs
cZt+vOsXSbTJbbekk0fIl45NuUOJDiXuivJ9QVuLi7HY6QoiIZ4oGJs5WSVe
pfyGlTeV8Vyso03Wh0sYJfztaP1vjt492xuFcE5HG/7W9o4AQV7+a/d6yMeU
1otFAHsB65vwBm8zihsqnaCb8YsBBmZVuPexb3fkOWaRq8nuypFSXJwdDrjj
nFHlge7eYZFXzFldhBHtppJUNNocZzyUc5GwgZFTMAzi16xGlMjwRGSFtYVS
dbj4QHCSaaHpVCNTB3e+3P+vTWzKaj1vndk/H/5Y+pRBgFCu9ZPIRYR/NW1C
wtWsJLU03+smEpXheqq9zO7UdbELPge8wr/d9AjXjgh1oJFaBFMfZZBO4vDc
/ma5WxpF9P36NYPdfigR3kAnRvgvzRusrKADPQJkGeDQaQbtVC5Bxv4FDzi5
d2gG2m/Gw7Yra20krpQL+O2UEFPU+mxLmSWmh4oWuH7Ry5zlPKNgEs/rOJwE
oTUC6qBj2J7hjT/94C2RbOqapuzVL8jesMDqpHEQec4c80++KTP7DzmbM4t5
PTVI0sAoMWRMJuu5bMi0OrY2d52Lo3Ikwyui2lKALSaoRTC30cyk6FPZg2oY
vzo+F/Pl6/XqCQtOoekiMvEidZapXMCau5a3A1pHT1Cxhoscy8kRrSLlF4Ol
5X/7ARamZyX8qLlbxaLXHdi5z7EFT9qGVIYipwkEI4oxBDo6ZZM+nPBJbi3O
kktYkyDTrepejiZ5F9XZR4BSloAd/KOWzOc9HPUHwE9ZH0chEPrY1HTt9ait
oWSVvM5HSozIWvyt/ljBWbGzZVRV5Ft0vwEsfLmTQ8PZTkhK8U6PMi/nMKuL
BvwB3R7JS25zgiNrziS6AgilLWitagATocdvLIhsPHnSA8QtcDRnypGuKVXH
Y6LYRKmBuTWwv/GriwVhsKrAGxDC/us4CMpSjPz7c+agcVNZYnESnz6VRPsw
DSwRT6TJa8cA133R0FEIT0ibY5rkwLnEc8SewddeYr3kVpyB4dJnyk0unp4p
obAkYnR38oCrQ4fAhpJLsGZT/MhrTJ6DhCCZbuMncHY4RxRjp8BjCznsrzpa
UjmK2q5sWj9dbLaUZ9ZYa/ufWgwE7YevCCUm/Z5bgDEiU1n5TdddRlZ/ZihU
B9xQwPkgOIpD7Yx0JR6zAbKK6keLXPK31ZVE157cBMXVR8amC4bO2JFZ13kM
9L7CuMdU39dx9iWySsdGT8kBYLmCPgFXSG3XzA/aSz+QlYypO0Wgah+QJfKF
QtKS1Rh66J1C+bXC/XS7Hsp0F6jjoe/0fq9ctxvE3TYQmZjOh+h9u8sUdHec
XfG0N91ngDb8sGkOSdKnoDP7qjRS/aGIVRAfbF1JPqC3sm3I9hVHudAZXR49
CZCzoz7C6PbrYGKvinAY3SdWGEplq++faKEw2SkbpHKJKJM4u2VTFmZjRnRZ
Xe5+UtO0CtUOGUJZGoq48DMEzRO5vOCEDL05bP42GN+eCoYC/KKNUXM5CYlq
qqE5+/RiZRSwbQr3FCmBFOYDYZzz3yr36ChOuN9tTloSYQ7cTAUkB0LHLtyO
7xlg9nfFIXKnL3S/2KupX1/+tI+p2pkZiiTm2eOO1EN+AlSr5ul3WrPiBn9b
ReJzrE1bZnJD6IcHfG3GTt5lMJyJxo8c2sa086bnZwVKlBSb8nAzVeSrT7hF
imi+zCXRwtE4WExPZIZ9pKViArW81xwoAUWYHjIDrU3JPZqfEGtIXMsdVG/y
luw91OsRD8Mbfm3+0fcRo2CDdDWLRwZf5uyPzJP98zxKPNiEkeG+tgv/Py1b
TNyc3B0VTNwIhIabE0MFTa1e7GMTMRBtzAVW/K6KaTUnW1y5hZ11kNgWyt6O
bAjim1rW1UzEEX7oWgUOtKRDT29QKy4h5yoOcyrtjQR/q6W2QnxSZsBURPog
a1MJsJqdqYAJskg/ZMzxXsD2nJRrnx51lRXylq04PkDhoDZ5YwPiIC7jXh6J
+6dxA05IjUDC8HtIxJPI6N9kjNBICKOM58k5jdNV99/cSmMywm7ytX++7D9y
5rSpIckQa1eQqIciYit4+oYuDvPWFR1ZR7J0FBaVdgNelYruehxuIrxC4sJx
tOiuxBrLkZrBsL6xoZn84h+kHLnuBAMr5RItF+XzpRMXfJnfsjPDdAgJtBUu
XSN+nSCd00DtXmnhFjFNTTShp7qOc8tAI4A8cq0c1wUGuffXT1AsXhuodjhE
Ua9I8Gu7DACrwA+9Nhm5hTHuV3GXfq45iI8iy4auBNCbFnlSw7opP2dF8hq1
t3ICE4m9s50KkTsP5u1fUYyxKTHFn06eI0HEMqdBkGT25bZVReu42Ki9SkMo
odjZp8I6hjITuEguU5450GTBqvDo6vbPL4JcGGoREAXxMPyeqE04iQuFy5IZ
mN4ss92DpcFZ0baMaj+4OVrkuYztCmFR0GYdlheWttsoAXDDn6r6UdJAwOPp
vjKDCWuSUrpnMRJIpmx4n7VMKl0ap63i/FUEcCYcztkgtaZ4gXRjwetB6rv5
c80CeAXowGFovL2SWCiJiA43f/akvlqmMJhZPSLUJYXHpsIt6lo0Y8ezu7Ou
r6bhglYzIuEBD174pZ9Uvt/3XEIGg76EJpfAQogELTIpYlXL7b+VZCbd4Wmv
je2dSiuUN1nM5tbhmOl6BZy5WKbSozg34WqZQCOFTjITqKtpW9XOtCWV/vov
tlhvz+f/cpmzEqAnAn020gSCfTpQV/0qxXGovfzmjrYb2HCNWBIecneLls4h
XU/Rw80e1p0vpBfVKvwtJZdkH0HQsJuQzAKQAWBWem6eykAb8hgYyPZRXpFS
Wo+tWIpWC1sw3m3JbpRE/f6hal4f3zv78PCd3Cem5wLnoow8SnLJ5YcB3oV7
aLHidtVe6zqRpOS2uHU8xgpJSr0CPm8RjjYxDhW/drUHv40jZAaP97Stcu50
Xao7Fqog09cLRa2QOrVXnO7f/5SZmGVkUDw2Cc2uyxbjFNym3Optnh1w9Cpa
mrE+25bpjr8zpgbZYPRwGJx+S0YyQXHGczjn3yaSnNxQZwcRe6T6Ejp/o4WB
3j5LifYeJataul0Fn0qOonEVknry3d0/uWqHQZxzCwT6C8hPW43Boq85+okj
PXCvG4Dj50N8DyWK6o1UCmJP62PSBIJDUkDq3iwagPgVobU3YOGDdfYOpDEy
lhE3i4yma4EKLNaniXCndbQHMYMvpZ00eMVw2WnQtVD+S90Kft2yypFdUcEr
nkMUTQ/EJMXDKCqUfs+vJJYKSgK54ZXW8EiwSI3jXnqO3++JLXVCMzx09D/i
7yqRo6go03D5p7OiurKA6Y7Y+hAbY3nbFt26tdHSTw3GS1DNDgJczNfylchh
ujhT0SMzCLwNlLEOZmOIbC+9AobTns1jQK6lt9MmbWnyBz/rhNZPqtZjikrP
DsCRSG7rMt7EBCigCZppuWwWOvecrba43mHFg7r5ixCMrVAsFoNcI2mxjcAo
vDDY5ybRYPdGiHOPuQx6UGYEsRva/PJUqOcG2M2Z3OJPweQ6ETRZpo/9MZu3
pTz8FUixJoDk2/5yv9C5YoGRe00M/Lw3qoNjmH9uUEjwB2EO2TzubBuPKcqw
sz+YNhlhasU63zvPdHB/O7pLAb8Y/wlK43mxKnWn+9MOuXanR/Jbe7tQAyC6
5TGV6pArhmVB6RCh4SA2y5m2tMp9LAVty4LeW+Gd4Og2OxVkCtNoYNqIec0U
uyIeroQbwsL1v+KMfN7bVu+EwD5cggE0fy8ZKw5zguQSXdzyMYKu7eWfXr2Q
9FeI9ozCr3MLqP/BNZFVsmgU868UtgseFsMijF/znUlS/xk8hJXYQvPcPTub
SQkgpjnio0qsuxR/PS7OXbs2BEAp53XlQh23T6j7pGt2xTWC/OuonUg23GIi
LyAjXrFteIn2tl2CGTlKGcvgCHjQOt/E9xyoyW2jZLJOpWTkzjZ3z4r/9lFV
MsalOyjrfUks0WGmplKpn0wzRJmpiwDiixxl/eglGU1CY9rihDIXuwiBxNUD
TQaKUTOctEYDq2nXvMNXvVQGPei6cJq+y8hD2ggl21REfbUWjg/jSpFD0xoj
61rrAX1V7h7XlVuDgG2SO0KT6z8ZOyY7MBiIC4LMYEjD08IyMUo65QuNjfsb
TN4x44iWNpUg+TJGcYA9+B5GPIyuN1fYttDizaKaJZRIvV0Wb5r8ateTklre
gUZqXLOy5KFI4eRHe+zt6fbOSh0UAkrsIFvWgDCQIElZ7Sc9pTU+q43RtyDw
QYNUa8tvHrYH1+VWM38ngY0hMvgF+tV7N5huzd5LixIKohsR2BR7l3dsCNRj
3xBJSoRBunwWpoRYVBj9pv0boIwoLDZh7JuLY18X3cft3sJHHmNjMI13uVkz
OgMpTZr5vd6zpfwzJUnBqqJqVuLucZz2kg8K+Kox9HVHsmhrWU3akDP6Pt0x
o3rXEw2556eeUKnF5RbsCubu6RLyLt3knkkbNJuDgS3hSA0F0bYW14g4H7EH
6sjq7ZJmls8bZbO4R0uFB+RL2TAHQ+lUIYmWN8oFlBBBe+EWruavLkabJOnr
mopBQBQtQkkw2BMP1J5nYNZDZzzuCv3qujfktR/C1hJyzCNE1ntIfpbnsswl
u9JYTV+k2PccLaNve7ENIOSH3OrJT6l5kZhDcw3pkA/DeI/vSNFfiVJ3Xtoa
7qpWG9lK3NJhCJOfAb1lhaRGKJkRSuuN28i8I8YH05ZZ6/AN+uKJt96IS+L0
DDzAutE9E9bH+S6XCf+wje1+MTNiV2uVkZ2r6C/mpKb5pWz5uRmUOoHtyBEl
Czvl+BCyK1+F+qzAKe0P/V/unM9lDOc2Mlzpmd77bjaNl7EBG4gKlVvmRN4Q
6ptyIXFqFFrvSLpNy5cqegV8gaiwHh983mUhTcjpqLFg5wu9dC8G2Vja0I+M
KctYNp2PtVZUkc/UgBDYdcLamM7ecwFynx3zlnJpjJd4olxdRftedpEJHLX7
6UVLKMbB7HA40g8e1us2Jgq0zzyt3eRO/PmQXW90PW3RDT03TAmwrCnxadoX
3n1EViykCBwXEyXVmM7vTryhMyf58Zk08aoPh9SPzCuPTwlAdKmSXhbseHJP
Jqu7FDV8A7tl6exO7J2+Z17UaINaNhsZJ1rQg6P3Q26KfDXYOry/HNARw3KR
wabffBkdeKv+capyAuEAYWgCJ8YLSi35pGMattQ4RCtclvn/QGtka24k7Upu
hTvyzB8cnRpw5wLAUi5camKJ8jfBMyICXqYhZIXEhsUpoe+X1j5tT8NxduSb
SMESEeLIkk6hohwOXcgBIfJ+B99/dnLzsrxDYnIBxlBzwMMiURzlISTmYBxN
UzbsGg/PUBgIPhGEV4uwNOj7+fbJQkd9C0ocbmFlsDDks63CMdr74+UosqoQ
RAJL927UpTmKLxbz/bF8eDOJGIR2A6NsuWq9n1DaoYPvNZmunZ12eqvzhRZD
a0MZP9gsouFXjfyhqpZUCtzK8lkkMjbq1wUw2hvABdKh21wo7PloSWvGMC4o
EIAB25xGVfLfAAC7CwoJgAEPsyx87i1wa4ZunNoKabMMsaKSeLGVR6j9BpDm
wVkICNU7Oo/BrHzV0K59Nm5iKETBvWp+wxaS9Og0MzZkCyxHWKO/mZvbIcBC
clmMUsyJTc2iNKTFT+b5XAfgyZ4VqHERH9RkCmLmJBZt1YV2b2p/6pbaqe1z
w3ESO5aTtwQvuRQuQb2lIdZH1vsoscFW6Gx2imsmYMV6XlahrJffYbSElmuP
3bL9PrE1z3bTjEaPxbi02jw45RsUI/lsoTxecH8F5Ln6yqoTETW4KGx6hQae
juElQkJlqwvQ3q8DvVVq4BH0R+1807z1y6uwGnbSFE7BpGr+zEOLK8DmJ81b
S6vNTyNd+SgBJTEZw4VKPNnM0tkvAFVPWnyTqfNd9Lnkp2ahl0gdXauOoHNM
S2VFLbWuzFTCQMVH/SGeBclzkn/IPj8KugUhwSLeLBwO8rRGzBdZ7UyUsVQX
iY+UJFo7sw8VHoJ/wA8DVAnJstfyzoVMHZKW1wfTDdKwEe1MTfi7q67z9aX+
WIqPN72tZ4Vv5MkBst3OAB9MWvu59W64ea18DyKqJnPsFbD54F582dayva73
cNEIJFCGIQfk3t41WTOy6h47FFyppFmTOXc+zeTfcItZnE42YsidDaMn7wBS
A+5jhGayjg3vp0oquNJpBdFG0MfTJy03cOhGheZ6xoIEoHX9jLTLPi/ZhgfM
GZYlfYXr4A+nvmr4xJUdpJb5x/4C5ZJbT6m49IvQ7VndZcZcSl3z1EFlNGuA
TDHos3XTF2YUTjeKR9O76XzgxJmgcNI9lBx1fV00mfy9nKfXCUGIhzj0jyDk
itT85xVrw74EEOXjJueKl4626cHfsds+MbiepjXk/iOj40GFXVGTDqd+teJU
jMYgQbN0gvYJ/tEKEbnZtugqTYDVoSpuLwoY6qffyLJrK0NfQM9GGrDfuLKu
B5IjunafK4eolYfgCAN38+HUBtUVTU5xbmKVTSBid3U9DD0zLYsUX7t1Apcm
lZTpgc7B3PL6vGDLE61x/RpGqeJFilXh8qnC10kSyBmxIwjPJaoiH7kxg13m
HWRrrLaXHOdnNwDHzT1+UfJqltlqdrKshYqOerWk6dmR6+W9cCkdAG6PLJKm
NHFlxDncKecqW4vMstWD9OFivqD3waiMgW9rM0/N9jrVWWGPIIr8zUnC3J6g
xjGE7WiL9zGnK3h1OH3Rc0IyTaWRMHoANqnMCYkRRX9H5Yj37hNrXK95nMNE
FMyEsGJjYpG1k3W/piBRMEjbIpL/mqLwV9MmMazpkuUmms3dUjlNElbITawn
WYGJRqfJ9kEDC4i9tilqEsoxAmOQ15+B0T/NZgDh8riuuG3eJYQu0ykqz2NV
s3DqmZobvkzQjx0n0FcaW6zUv6rJGe+I2QhVEkoDIMmHOGm7oMf3AOMsAemw
Mg5OozSdWNEOJU4Un5se1ghMpVzpYkyxYvd8CrCYIl+PipdPB74+kgRVfd9g
923/7wEi2imFKHe5Ia6Dm7zie5UjL0VBJylkZI1/7ERzFq3Kq+MltycTxMGv
ljHLiC7ZMxyUcxbX/HJefa0sQuGuz7qcDg7W8zKhP+0gk8WjRCQcdqGo6LlT
MnoLIzXVUbOkw7jIbqYCkepc8p/i+8lvTmyzxkgy9tpOESMXNQ9CIurYKxtY
ZKnTD0IhNWjFdellJlOimkXUgETDnmSHvMUry/geTnf9CNLQGIUG4gWUv/B4
Q+ud5cpPa9uBwfUnlF7VD73+vR3TZXJoqW4YC6ESldtuHbSJrqm5TGZ3wLtZ
9+GLCkbYGhpKwB13qAbqZFZUrPVDy/IHDQZMJzdg0WszpUWUUe8Iq9+SQeqj
/SgUdyCfexFns/QtAKwGrGOvja8uc0OG03xGOvBpep1/JBwWLXaJxjuwBP1o
b6ZV0WTuXDeHJTVM0G0kMeSvee6iEkMlkZrLvzpGlrAAdq3IDtXacxYN16ri
lYGZW49GP5DxC6R8QeTECUAGjxyTD8J8eM3ElDhxPdiM11Q+9hh21k2RFACC
A1OTAqhEQ4Bk8S7MvwQ/Hspb6dYcGQJ2lI0JIPGnN5IKvjn5OA2yBovlzVwk
XFCipTVoJpS3B05K0teibCgmOczRddazbTTIZkYg6pVBziZtMleRE3MW5/o+
JL6bLbZXO9xrz2OBP3Glo9wvU+aYoaM+XSXlglg0Vn7MM9Vh+ShtmksMmgIy
XiI9GGFUOAYulTKrXpY06t1okZB0KXgvew8Sv7SH0dzTngUPRCM2dNrcdqLr
5Q6TqDx/LxVSWMYzuiLvtUEirs2yMYMO+S52G//3zsKjU2fSzfi3FSCLTv8a
ZGQaf4whtHMQCRV8LPlA+FA+qYXbvHz2QTqz9sCbeK6YEo+79BBTDLVM9o37
hEj0ljGjz10420Nf/EVxF+aX4fJZ8QfLNn5tQNdiJMwffnDBZ2TM9EkMUeP0
uCt5i3itx8DTj/YCBvbf2K7ybiXQWBhyzSTYZLwb2c7s9RCo/y4JCo/imC4I
Fr3rNlHTCNFgfGEeW6M8Vn2yTKyvtq8p3UbSW200bOiJExtpxb9bI39Geu7n
4E9XKoP5MlFmPJUphrXi7oroUdwGBVMFajDz2RfmMFnkl3m09quElMD13L3Q
3DKy3aPSKwQCLib/EdkeVz1a3AyluWGW9ymo917mGJyxcWAjosp5FH2ZAdTQ
xRG7U27DV6fDv0j+0TxqWQxkkTagwhJglMShZyAvua/6UQIKEKE+a2IWBW3i
5nKFT/tsj+4/78EVE6m5yv4bMIJSD+dL7CJZQTiHBl9jOWKZ9tAbLBpyzBWm
65V3l9RkuVjPSf48d11GdkIWNMtSwMjrkHpMkHICTiCNJR+2ZiXvQb7bugCl
2OJ0vtUUeTGiNMoeq9vnoAbnW1ki7YjXSF85/OkQxFs8b1YEJMzVGtz6aiRg
g/VQVAKaPvyxpFiuz2ANeCJzsTw9cN8aoJ3HsPmk4V7DAQ7RrECFJVltn870
wPYhpNZ2V4Q4PnsxjKXbJJXIgPtZtGSjUI927YbXSI8glFkysNB2IAOA3V2k
1OF+Tb3Wta6NX7W+gAJo9oIBQkFSxy74rrbLYeNvZ32wYmHhD+RQ2ZrL85mx
wB+Zkohb3klqHoTJ5Qbhhy7FwQ8Bs/UhshqM1jxh/q5oW1avur5ikc4UjTwc
jzgDasODjb3XwSBeGL9KJBcEE3IXpJdqyBD0cZ6WUoxKMOAYdKnmcuycSS6Z
G0Y089ZA+sGquNOLlgUcd47OyxpBN5WY1njwGRgLpDw+M8b81jhXMueDtI6M
okJZoYHkDVrOSrTay3IvV/jU8dbLxapsgsy6QSEJ5wCtVE+YRQdZgbdnBWP7
kkXc7anz4UmGjiljFeUiFaqLek94yQklJrIEHbWkUyExmFYW6Dc+/rI8bACr
LucX1glHejf5Eaws69V4TrQOKtbQ1b7cNqOhTYzbrtjhyxCmceUQjY6pu1fH
7JmBn5oHLyyXPSJkv/gxCACxtc4a1sOHsHczk8jOh6eWfeTnY1pxL5lfJzuU
QZPlmNRz388cA32iKhDDngq/Gu0un/wNCE1z9SjzsjBAC59ewGL5T9Ixqoln
F5AhCIqw6wARIRGeN/+2NX7wdlVIET+D/6ZS1L4ywGKaiz4SdvxAr4/fkvEx
funWOK5XEOJQ3oP/WgW62njDhDsCSRoA4p28D9RfUR1mKa5z3qT6RDnlvQo2
6fnTl2aK2UKfTDniPm3u35M256kQ8tExM7FVlDR+pi1eDgdPv6lDqrndhjkH
uuGQ/xQFemFjJUMnvSqLzKp1xE7g2/QaeWyjHH8B3bcZ3xzTlyDyaZV1339+
q2BuMQv0TtqxGkZEGR3NTUWvL/QXQqi1NpmPZ6vGF7xV5gX6Y89H7fIgbadT
K3poZVM2h4zRDqGpd9tAQEpdt1oZ9G/oxSgLOZE0MldBAEXqLvLZ23hNIOVy
zXcXXa8PXUpsPHO+7IQC0byFwMDWlguSTquCNWy7820QlzwIDZu2gAEEAz8q
iuvrL7XPHmRGaNGPKGdkIBiD4EjXGG9CmVQg+96RER8A0zZSnk1nwGfMQiHy
ZAIl/MYgCkM6FJfXVAl4aH+U6iFqx9vpo/qrUaTtqu3wqtYf6CFAMwxRoHgM
GU6FvUQgNHYz3CkI0jt9PtAhuYbvwXIV7fRacM3sQga07L7Sr3aQlTcrh1Sq
eKBqiatUyiggWAwuGSQ59FIhUaibxFIHaJkNeoMk7zXjx8/IhrPIoVOq+25j
jkIHpB2wKKHqEzdOljHvxceaRUuTqDqeMkOEZSnrDKa/yL/n/biSO6ijOFes
WJonnCakgnzLdMvJ78sXqJNvN60cPMtTeY6FSuA3JCWlBs6DFYbuPCPo17NZ
D+1WsVl2J0lzqYKj/Xx/v83cZr5QLtDmdnwPBEnr7ExT3b7+EHOh93mpCs1D
GBnB1MK2LyIFx6m3FjrbuiuQR6O86veTEjnN8WvPnAD5DhtnmLNyaq9Xl+9V
EVgwwoKxeLD8oOwlduyMqc+S0MhjfztsWkBFL96ZNgwTj9yTIYIwrNdHHKj3
DbrllfCwYCFQL18fBgZ5i87b1D/CToiCERanizFkKAPtVLShJ6pSvLDkCl4L
nvOhPRR9sjS10HtsPNCk67PuAMKoYa3aBkB0r5RV+Agan7RyaXTvIkw4mP/J
7sNgKLqHSTT8nVLL66Dar561j2o+j4og0ZGmJjUeuCNqYAub+2U6MYz53yeK
+Yju4hVwvApS1SwmLGXjZoeCSCLK43PM5jx1FbQPShek6qt+HiWUGj3bRywM
E8U8876nbT1CFt/h4qwAk2zQDCRYy+O2QLSA/K1rBiZgk9mQqx8zBigg0yE2
WGHOUpKWQLDNMIr45lnAklpDve5PT8pG/L4VIFX5d+vSr4rR8PVLJTzo5hct
MbcGReRmdAH1SnKyMxri5ZU3yzTmmkyhn3p6quuneMbzHqp+d1XTRI5JLcD5
MpEXEBQ659E8exv/O63PHvzl+N744oku6DBrM22OuIU0UPtDfFRxMkiYHHQC
O4+Jm79X1sKR0y1EjxA+Ml18XGINFm9vF8VXD0IoWhalf3wwW3hKYj6Xy1O1
qFkKe3KmhoZF4Qxb+NQtVAn8DGP0OqTooI2/pIovM28LOeshtDrEn1/0FGr3
xnHpCgVsu9fhhV3uxiYPKygvDNkkZjmbq1GJ6ovjRIin9i1JhyHIHmQkIqB/
62rdc4VWTliPW1vVqYWp017MsKmdqsvzBYjE0Wu2Z/6tgQUtZ7vVdhOh3J3n
XkAcMdtRFS8BC6x4IcRxWzI4SRoqZUkXDjCdG0QWkn6yoIL3JHuxJbXm0TP9
d1hSZNXetGBMcbWtNZHSTnRdyL1EXWqTlwBCokvq9X82MX0YIPJv2PxiS0zQ
7MDeUwcX1c8gy9YkmTgUvHmR6ETsQu1lDSjWTlPvEFkmtvDZ5li8GHg6vYCe
MiCvfkylcnW1aF9ia3oZKEdlZUBvQtsvmr+3zMNVpxy3oOVL8jvUv6sbyGD9
YIvlOZIreCL00TVk70aNDYhammoTYBsShup40VXGTfTPTDYgEWhiv/Q5mu15
9cc789Sxh0cKQpnIum5yoghQFzxsf943oiFXI0MG/Jl/EyB0pQqOjK04LWUw
GV6FKuqMx8wbs+uVJfVX42jkyWCSlh/VRRhrrbsSKl7c/VlpZGpATs9LpWI0
bCthcPbu2qkCaWohFgl9dqSK/tuwZXBfSOFN7VDiC2PWD+0h7qHaVAL2rBLJ
2d+GehqJplmR+cMUyxk6YJcZLE8nJpp8RfBPL2Qy3jWd6tmG1AoEB/uJamcA
XziEyWaZSJjySLQYTNKppVrcqKaBolw4bxfUtuatiUcobpE9aKpttf6pzzQz
x3wVovu7lxxZhZTIqT0dOWL8GhCIPXDkhg8arx9Tpi1AL56/ItlXpljLlyIx
ERsvmqTHICINaZZ2d3FU7h7epyQ1k2IUeM9RLdPt1T7+95yZvvbah4ZqzuPx
F1hXV0XZwayvhK7KX3uB7T+YGWIuluYTRrYLRYrNX3zhStjCnmpuZRCU+UhH
GG+7wHiUG/5BZARrSDpBzUf29A3sPkbEgumeThOBBqt2eXOeUx8bFYnj9bkC
9NzwlHB7J0Kso0edv6wi+FE1wDXYUpqTBUfLDRIxFtJQVHkrUJ+kEVALg53t
q2EMlSo3Qzsly0jYSbbsjuVwlTLYGpTCJghsnd+XdvHIBM2lTccUIGb8+4AG
kzlIr0mPqQTUyLsC5UkI+y2P83FNTaGFvJ7MIlapH3Josj7S6dkqzWEuKnGz
qp20kxTWyXhcXR+8EpvorT3rlgLmEjIYhi1BHAj5sNMdtaDlsPEcyGh/ivsf
Y1ZB9RbcqS4PLbVK8VklYYO/iPB/lMEeLDDkJGG5MpUzdjVhAJfOb/29I9lC
V2oLisSZyQ9HIyrnnporUEM4WVTm0/+jsh2DnhAJzS9L5mwwfME250Vo9m7J
kPOr0d1ngQGbdy/F8+UB/ffDgPhxefka408JQp0RQdvK895PMzgfW8hERMxs
cUk09MbBlWKfRAiGzjBqrmAuC5y2O9xqjML1TqbhfCiwXXJtV90z/9kSL/Mn
UNdad9rxfSIsqB0tHyPpO5Qdc0dp8BuMCrI1LzDJtO0uR9w0ZYxGi7IBTLXQ
h6OF9WJKMsut8bbtVb7sMwwkdUhZGkP/w3dUU94GIMVrnirTnmW1pCtH4LZQ
G98cTH2Ivp2VPqjWm6RaEWtnXzFCERus0ByCqraERytaUyOX+4wfgJG4fZWR
IAhWgowfBKi+wAO2/IMU6WQJ+y+FL7ECrSI/Bu72UG2anQ2Nxa4+BTeA1Z5J
zHbJHCMSQ3HjSyY/AD+vgcver59HueDHRo1BQww/AFFFe1njO1YSlve6bGlf
vKp8C1l8h6IipRdlQsWo0A3K7qymJ0KRoEy8XvNnduRBRmuWTRjYPHeIUFS6
p4oCohqhSYTHpDmZo6Oig7fOrtOxViMSxxEypEArOOdG4aZfKc9OFseJwGle
TD1Jr0aLwXGxdZbl+13Eli6hiSCmmZHR/PZ8b0V4lZHWB2gGCwX5uoQG4osp
xdoits8Q4c/1ToFAqZ4Upmk4uT2Pc7pHLWWgPAQEY1UJS77jkVLoR9C7qzwC
X3zqbqkLRA9CdkhYn0zqr3EMp0ocEV1i+AvveW2qh0+KIMEKK6o5NqHRd+zG
aQSxB0qzuPqLncAsFXZYibHprRuE/dknmnFGWjbPz34V7veP+Dmdwt3SGUcq
MqPY4bx3dOZFUB2+XwDL8dTgLa9HADSM8Po6z0zGoL7Ak/8mwxd8XxzGv8HS
fV/8dEJNv9XhrnsqqhAgHt9WwCP09YHDbT9yZnuLqp2yz2xQ4AM4zEZj+EaK
+MIGIMEIaVuVxtm2spOrgLwSqyBH8qvtQGA6w+6Y3/ZnV5XK0C0btW87r82G
W4tPy7kBWh2JKLmEXVqaLVN/u/mYNCjFjenZXeAI/S9nZr8PPeOHF1nsQztZ
ubuoTGmoO6rSj2x/cDpaDJRCfNUzAkHjm4nxbB4V5KZwfcKapLaezJjIl723
2h2ZYXkJc6d0+jveIC+PfQnfx2+9k/BAgLq5J3PAFQwzpg7Ta1qfFjeFlXXf
OEUHJQEOabizOEBCMkJ7AyNsd8ST+Qbxybxs91CFca//7kVuuyBHe48N11/0
LF+gpUIdHJZ1ZtNTvJ/FLtcq+c9Y0Lagk5U4JtIiy8nJG+m7s1goifI7fDab
yrwnie27pLFyiI43KWwaldeB2AVe4os9G6QQuYfs+DAb/7QXBnMfuN457pHj
cr+W319fxk8SrT4tj83oiFbt00NZ4aFJcay066UnQaNiVNarW8rvx/DE3DlV
sY7xwVR21cQX9uviLbbhBxT7ySNH1o8ZGzXiCxO0PBK9Sbj+0K1gm4dzy/Wp
FYl6lqUKMcjNBgSwsQUeubarmlOR+G+HtjkYqasHYBxC1/6yRADhIcj/tRCd
pGfI8tlP5Ui4nYpOJfcVLPvpUXo5Q/7xU7N7JGJsXei0HYxquOuNTUFfwue6
djCOUlsGnbInbCfGAcw/acQgJGzFz9HsVDiaHbH/PDKrghu3L4ICUcBj4B2y
DR+xBpuU9+F++Rp2Eq/D8ECcMJIs+Y86gHkCaT0CZSSP6RnTyWfVeqGunBar
XAIWYrxrXWPJ+G9a6gwfjIZxR0sG68amyy9yXAtxhFx46gvLmmlf+aasDFNu
RGPcVuCXiBcQNme2qjPOg51XLMSkheet6cCny0OXsZp1JJm4yJOiHwkclBvC
MHEZ7oWsKmRE+0/oO5Z+LZNsc/9zAaqWWmov0UMy5Krhlm1a5/j0kuepzYZr
o1HGBaIyjs6/TaqBu5NN5akfO4wDlZmem+gCBbfVjFNQls/mhSDfZiI+TSf7
XqJYg6Z+YghDDpDNwBM7UFYEIq3TOrodbmb26xnsWMiHwSDV/U9RYtHBpWuZ
Fg45pHg53XCRDpBR4WdZgUnvOZlJtYU7LxZZBQXifLqRpwAAv6ReAltx+/JI
Lk5SEXwl0UKllY33aZazXt2xuTLu+v7jb2UbAMS3if+eiWL01NxwqDP/uMPq
2csWmAswPoQdDQSpRsEI5I/GYw+Gy5qH0NYW/1NeuuU+nIH1Wxu7+LQjFmd3
Ui39cZwofL4Fqs6S5PDO/LSJiRmmGspKG6WnM+VMtq2HbjFoyquafcEpnheh
jY2QtkGMpz7turGlfnoLY8Eo1Fuohh9vkogRzKYZU4v+5+PoO4EagN6KiKOC
JuSkf/yzcjELPwVo0hez6zYlKkXscSQpkiZrWZHAbsE3GqscnQqc9Abi2uP9
NUNEgROObHvwrnp2T4CyM6Zkes29JFiNILykWhGlPE5IcCr0JK/RN2qpB/fg
dnkMr2+8LJh6CdTM9xQjKhZd+Q7UaRx/q8ipADim42eG47DUMZuQx03TF0Nu
yJk2NRFftcHslRVERPJ3+wRPwJkgbOkAFCpPnUUNhnNf2lj9H8EDzlhbLJwG
4erx0+QwshV5SYA4QA059Yxnk5DuVtu6ncnWlxX+EpgCUMVKcdOGGAvrhMGe
TSQyak2fXtRDeLvcUxytYIJfolDkj09fzOETkr/wBKBkejqblOJWqcyXjrlY
FT0t0SMGHd3Muavg2UTaIlNWHpAe9onmqfJDtPHqi8zFC2zZD/cHRKcsBnbs
pIGTg9nGnwuHBqbsiPOz0cR32xATAx7EbfiZ1PQ+VUPd8233sxbp45e+aSFt
2IVqBWFKujb//gmKktV+jHgTVVpftvJ47OA8BpoiQnWZdzsMXCnb8tRM6rbR
646ZvA9WnrxQAtL4H9sYEAlArrUzeLZIV2ra85T7RqlVCyURVno/xvX5lQks
DWt0JAoMeBcZJbh2yP6DajR/i9QIYyJgxMlvj8DAVh/eU96LzQV/jTz4Ztf+
e/oX68DXo6hJf0MD1sBxjY/VrX1vctQByHTNEDmhCLvv6CqvB+YdLv81CgKV
JoZOAAKWwo5v7mv0CJWiSLQsxHs+jYkES/ea/e5SdyawQ/TGdBEX1GrSesOQ
vMqnAHwHT8wzjbsVi87plP5dWX1jbYP9oCKFKFx1LPE4EWJq2C2vn4Kx8Kng
yi/9BLCKneriZunK7dzmArU3UVEVBqHyKkNtyEXIXTmKkvivxtVlH7hHBcm5
xUI28h0qVcQ9X8zOA/H/WeNtLLRqbOk4vCr4ELQNMXsgkxgP4nRxd7wT3Hmj
OAfMYCHwm3Lpr3TGSCHnntxDQ1A8fJE2ieexRvKCGNfqQ3xSFez3FKu4djVh
EPL3U92xKJCvdhLIdD6IcMBXDmv3EebFCjqpI9e0psGMv/3yqZjF3H434nt/
WPkhvxd6ojIB9NwBfOjlaDnUY0w2/bPSpzfOLFyUTmesDxho5uFtxBR436x/
lwgbf8rcF1CoVvJFDyRxrfojQapVKEC7fxEGGXSd4fGPrRhU6RPzye3tb2rl
XxY8FzzsAOZ3ann7o+4IaUBQg1Pj5FbZX0f0iGK8YUHJzgogAnQvPzKBBCXH
j63L+0H5Ens19KNCLZro+0gUJFTvoATPWY9YCh6k8fdNncmJqEcPrn9a1N7/
zO0cgkl4PDo5s/i9XVSCts+i7Q0v94jXK/ugiq/zib8NMNq2D4dMz9MgEAl6
+gATGu9k/Klsrj8Jqnmmp5fqRBlllsWhAeZkf32QIaeq8E3LIrhWhCev/Mlr
kgKOyJCFCGDoXIl4XFLKHXQDwGa+xPqxouebwYNPhL8Go1JRIjp/ZOv8gAD1
xHHG9TuIeExqpRVQjerv2D1ZqxRj+lXpDm0xJURjmdEgKKVRLyeL6Ok64neB
GKRU0u5gLwntZrL1EFUokH+aKfITaH4DDMwCmKAX98QeMmbqcvA9nAfEbm+U
uMmOv/U2bs6u3Y+jMlkQ9nWqzKBgHgUr7ZiccYshCkyzWe5iE7CF5z6N7YOc
K75jWmIF99Tz6wEN17kZscDLFv2Z2UdMiQWJP5yXaRlilziEH/sIFAaMZOWx
cB0u9KDUDi8GZTePUkE5L4wo3ROpVHOik1/Cs9lb5cinYa+sDvCmuWKZqusk
SAuf+vc8aqTiExPyyfVKl6AVni985XUliOsfrogQgCJNl0gb32SYzTEytBXr
gbhvjL8uUh6wBf/n73XFeWY28jD7r48YdC8pn53h8Du3HOryDuC/Xhd3ZwSH
Vt0WTB8vO/B6XLtcc6LYX+WO96oVKGxA9m/R6mKFae5luThv4L7HivSh7uVl
c7HDwrHllhV9FbO60kSpfypMrJpTzwggOWJr7MbZcyp6wfv0pc5UUbgZPnrA
3kg7rotG5vIvvbQieF0T7w1g06JIx8aF5vhvffWEnb3lk00vbBKJtxIY2r9+
sq4UK+u+/QmozeVHLm6j52a3oc77z4WzAd70RyJ3HgWSlGo7Jru4ToTxTBkW
erFyAGpO7CtzPuYgNHatJHtfF3uFOGMmdUHFN7EuIP5dWHW77i/30+cIo5X7
c7JKjngehvnlKJTukc4J64b44lcCd83HvNf53a3jJ9D8/i47QA86s0UR2O4j
GdFSZP4N0CjM0vsCuJlHSdTzgJtVm9BPyEQ1t6YnbWxKQ4cx6sD9RWDy+8Pl
ZmCa9LdTLQhwpzSdVIhKFn0qCsd+MrQO4qUMouOQY966Z4g+Xdxano547rU4
ZvPwMLojb+tZZ1C+74M7/2IOkQBL96avpwQh4hH7MYExXtZk8g/6I5mmmrgR
h2pwlmEFmY+6kcWp2g/ej+9DUxynclhwDcI6PWNb1hlzpvd6xFYBzeIZ9e7N
FPUAkuCpVU0Qp2enwIeDThZ6O5x3czQB9LQ56nGDvTotjen1j1ndJLP6le/5
aUXJhE6xQHNTjFnI+jPCc/cO/GPftvAfqp+3q18nrxGoBOLAFol2zDE90pSj
WtjoAEhGNcoazjCOLLK1eL5pTlBSRqcweTcqZ+3OTDgcq0HbicVePP1k8fkc
+SCVKa0OUYvJkYNEn9TQPS9sS6G3CAZuZfbWWfwH6wT7GfXk1qOz48qTFW1O
L7RfHqfPi6uuRfCO9h+1YtzqRAkYAT4vasS3mMurZzhUmTWsJWQ5T0oycEeL
HNh2896UKg9iKGEhSb6OxHErBqe6shhlvfw9j7BQPnGylw5V8J4UvnsgSzkR
SonxQEY8/SWVZU9m36H0FlqxwqrEc6JuDk1lqapLMO0XnQAfcA5rEYsUqp3a
6RV2+JpTf97hqz3N5Xe6uwTLskelJ+IclK/btoSTY0dy9Svwo7XX6W96KygG
2APcvfmB+j3zisb17zz1nW0kWJtemJnqu4Nfms0DCdoBPVH/3yWqGk6VU6Dp
KhsIoGQ4J282qjqq5S/YTJZgpL4yUgTH448B1VJa9fems6xbev5dXiMYieYV
KWo3JKpQ9Xrm5KOXJpPu9OuoHYYYQSr2oVAubGk7whkfGebtUIPd+5XzBB2W
utAAKam3raHlo3HvxKEtoIHeDRc=

`pragma protect end_protected
