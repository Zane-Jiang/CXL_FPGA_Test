`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
gAw9yNGZolce1ZNUZLCPJQ7fxtjwaQvvdXL5CGNhnEhdsHF7qlCKKkOahOGkr0Ck
KtaZlmG72ab3g/hPv+meBnPD4j2zxKeuGJS6OygNlgWLXtU0oAbSpE9K3Pj9DVt+
eJj6wl3TusRfGNQ2nHqGFuoZBN+lHPJbyeHLCGyAZAA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6768), data_block
XiFlO+hBnVwWTPiRBgET8j5JSVg6Txzhrwq6GRp9yaiuPfYAqwaBXU4Yy0OOhSk/
thIFluZPlIu7tjIZ2dxVcoxdKkxV0wujZkNBY7F27NIf/nBIlzaPBb7KhvDFBwtf
vaugxTMED0qLH7dftQHmgZuzG9zkT7cjQZNLbtBqpr7E5VROM4sAeYWIjcuHkTWX
/68eJWHx9HOajNRPW7QhEhmGxfak3Qoe3u7gPXnEQJRHnqkdzIRJcqvcstNAqI/J
KUD9favaRbgrAAgjQegbUOIgeBR6ymONjwRmiGW6Tss1m5ivXjDmcVUJbsTnwFlQ
qw37HAX+cJWAATOBM+i5cIoczBzfHp3+Im9yUTW62I+Wfncf/GedVL3HqUbj45ee
8WC7b3aTw0OoMzwlAqGedfgiX4nhZuUaDjklBdWaKhtYSiHDRa6ndnvhB9xy2Ksj
Muu8QIFfyorZdVVxH6ihDZ+wLDVhmoSJIah6yFsNpOX8TWpLvp/eDUfzGUmda9NM
Yrt3LTzfp/YPpQ/0Hxnp1NJWasBxRWvGw9atyq96zAkdpuGpc0LPNR6A2NIC8MdL
IvEv0Lf5uWJO7M3LeQk5Exc4sblQU7x3XwzTVmaNedZ1np2j9Zwr6/PzGm1aiKIp
9KIm8VIm9uZawrxFXiZoBX09iITexXYr6hZgYul7GxHqrfseGI/65j1Avle1GgAB
WHPUDV1hOmflE3XGq7O8OOB9pFA+g4n8E5KCTYcEItIoptTMqCeXZvG+2+ZEpdAs
dBpNH4LCe8iW375p9zpVHZEBMaAIb3mJVOCxmf0JdMDQ2LIqmU6kHZsL2X0Chd1v
PZcnGZMyUmg0L6udBdzPAwABcKGyEIpi00RUr3HULorb5MQTfCpW5zaiaag751ZN
+8YdlnKkA3G8QC9zr6BW5YL+O+n4QSAg+4O3V99SUHG4NmUo0UjDnqW5NtQqq+Qb
FzQ+5HmLAyQfNQpAEGYWQ3VrXi04Rz9pSSTK2RhRzn/2wd9PrrvQgCLnw1QYkzhb
bLK0rQh8GYDh9wiAM9k1c9gbmKws0DC6k3uOd7RDoIaZ/kfLCBEfgK2HF9gNS57N
5qCwf8e0Lsj05+ckguoyfqImECl4XDs2Lk18tdQmmKj4KnFt5vht8RWKozWcmnk2
2+eqJgHSuvN/NXl0jZDZP50wAG0iZnVZ9KeKuzpcD8DPbIqwMnIDQ+53OxzhCHMg
qAs9oByLD3BeNibWgMEj4OmBFtYcX6p5RQijZKLwqu4d/o/L1mzD6Q0ciD2xIv8a
0I75lIbjf3f+QEtP1mxMbXHB0KwfRtHkNoq7Rg/C3V4ftoLigtJ2SjdVYmlA5Rue
Ri7MA6QHHCHnR7eD9K7PH4ROSaclbvr0AOyez1S/21XpW0LnB04J3iFWqVbuey41
g/XZLraTE12XjRQttJenODcBpZygmiWLibzqUe7marp5JMVhSurpZuOMVSObtNtn
S1lsvM0VElMWYmuAYNhGwmx1J2esLU7QSjqw85I3NaZMJT7H0JSeK1PNcoH36dxn
vvhoEjtM13OPnpRzcTeI6zkcJB1yzckNn9LRpBkVKMkvSxX9eqeObICr3U1Z+cDJ
nDeyhzyfyPXeWLit0x1fGpWVlBVBQnNTiwQjeif1hCpPpzG0YSOk5Cr+tK1tfYl5
FqNUUZYp/vlt5PdodRhtLmGpXgKGqNlDeaQ2aarEKuBg0SFUrWLAOW1nnLWY3zzc
7n+DqtkfQB+DXbXtFv9fGUQr2qZ/zFLYf/diV4Hh6WA4/yc3ueNX/h/VrKL/Ke5d
/9rm9ACF+RZB3Z6ZXjl3sBCyOn+uEiwaQNXfcdPB/GKg4Fx2agEXfog85/nSMcEv
7vlJSesQfMAE3or+nrt7qD8APqs/ife/EoOWnicTivdXTVSvbqBEm/opJHZeV2LA
d4yRM1ET4RufinwUWAF7yjCEsOvBdNIVU3iKr1Lln1Wj6BNQsNHzxlf9eNCS8UZD
O/IbUjGcvDODrHwnFqp9vGE1CXwrsByosM3JLtcCfqimuRLKL8Mw34uDPfcndB+y
Emq2/J51IIs3H2VylE6/mneWqWKrFTh7RIcGXCxS1wLkCb7Ax+heSXcgOEboHOXC
eEBA9sLN7Qq9sqJAiPEJoT2wVToNk4wkrGJBu6V1a13u6etTKh+sDPYd1jJJJ2R+
eAjBuqOmMxqBEhiBuSORKV0VpPtulnHBVPI4LUkJ8kZSNO84uwYVkUQHoFQH7JmX
UKt0D2Z6mAnvQl39U05dEo3uhFjDpqTwEfNk02UX7ZWsMF8PZ2CtjNU4KKV0pGam
1Me1kM5Mcu5zn6Rtuy+A+dOL2jM3lG8ExOIAXCRPla4ZINuHGh/Xu2qOL4qVRNdY
qq86t4l0xC+UWYCii5xMXyJPdFHpbBgtdMoyzj+RqusHJ5x0vzZRalXup5zoWR02
Ge8B5rFQWaiviLDEjrdPkfGmAoidWFnWvBMZZYaW9FJ1afBQF43u2NyX4NyPHgAI
HZx5sCC7y/wPrBZWRot9BSprBFcg35+KpthxZ2BiLPvk3CWRS/XBfBxsNSZYbqxf
sUVcRabbYObvu3KORNm3rfFpAsxq2S81q1/TMdb4+FsRB4lR46buV2R4BZi/hPcp
yvrOkSP6LSrE9bCHM2eItQRc6RJVxSF9RTe03zyvHFe5lT9sZxljxSTm2SXAm67F
aVRQ87zyrB7VtIHT9KPRKOyu2G6nKFGKZ3P3P6j1wn79Gs2EmlkrqrA7gzIv1/N9
r5zz7sK9GXuf//4T06JxrtSPRwSrdVVjdLMrAVImuFCjM6EU7sg/Q/wXcN7FZIZ2
Es/kieNfqcM7r3afdD8P50A3AdrMHQc9A6b8RReXa5DjEMiqxyZn/zIGDHSppUmE
pcLCUWEGiMIOB8RFRaMBnQPeYMyyspR+lOU1I+qBd1avaWraV275YxTCkDjJGtrD
uGPanuff1w54QJtk08rOxQpzQSdv3Pj4JHD8UfFsUmKJCHs/ywnQl8fmA0JGsIsf
p7DtgTN4VHj2UxtII7b5pOvh++7nkLsY200eSJoHcWx+N+WNkhitprfmf1BZvbbq
ykl6naQLVJbUmk3hVFL/YMyZqtvqmPg6uAs4TGtzOUEgg7TK9yUGgbNJmjiWQkqg
BsPaSr1iDQl13mE3hzl2b23gZjSPwbVNbNx9KJquIsqFrdQ2llVFhYWAMCz2yLlQ
7lStQSHOZezKVfggI0EX/7Rup5XP0BVvNH221wMB8Vl1ypQIcKYyYjB98UjgMs89
xlsrsJKTcGpPDjRzzRhEjV7mPif5J0dq4UI0a9MrIopEXCXC6U+MYajtwssJOtpc
WmnTtUW9uBZgkvdJaq/brVOcgfw8QjTcpnZ58AItWQ4H2bnHM9zRKLB27nvM2/9N
PpHpaNklZP0uT6ngy4XDwoV/Y2oT6lS9GmutULnM7XL9WMdknwkfK6HXiw+mAU+1
rXFjm1kOIP6ro64N7XDjnqOVrk71D31SV8BgKlIVdfo+o5v5ECxLZAJJI4kvdIrG
j4Js1VuS4+HQkU3X42cCQ0phDrdWdpqCkRMFWxvd93TIdsVhq5f803NvzH2hGx2F
2L50lyT0LNRqQ3BI7SQ+0HSvqGzNHu73jEKY2M8wJlTlVnBkfRa3Mk3+4RrC/1Db
DgGjIip3aw/LfH0wqg55owKipAnlqYxi5NDWvT79RBbtay+Zb858tfgH7DpnrhoO
uStzGjM0WJ4DHEeg4anD4YtNGi1czdRn7mwZGGfAfGkp2VvhnEu178bhLTUOU5pl
cWaFhgY5c1sinWCH3Fdj1DRyFELsJGPfMWGS+WAOAxG0Fw3fWrAcYZhvhxAXyI44
pMQbQp8G01mYHuWr3ea3WaaN1Pou1RhVF69eqUDY+r2lOsV5lraEuDUngwf1k249
oYRUx0bMwH0u0ln9ntv+kUWflNJMRbUd7I4J3ao7ITElYXbNfsZ3cnB5nCgRnhm+
1Ih4jFmnzsyFpXCkXFzEjkRa0vyjuaor7/Rs6isUiz9SQYrnMJbv3AdZhZlDPlMd
sd3wReN2SxGAtum5FCj6QBkmIs0R/0ZbDygQXHu9S8JzbJGsxCzFEo/djTZg3oJD
Kq2Wb7kqNzbpsPE7Chq31R2Ng+rq3cN09kba/1mTsKyrHfB245DQm26zEhnlR89B
qKrYVsrRmPNIUm3ah84CaZ2HGJumyuWTfPNfp7QxFV9HWHtHsYCtbfExeQRkHuOR
nbbsIzzgj8bUje/a2vB82oQxkW55N8t0IicksTShFFXy+NLojDoRPi77n4/sqYrm
a7sGHHL0OEuli7z2G6JG7aAZ7FpquB4ZUmuMtAcKuhVwSuDnz4mqfb/bTBfCUrx0
smjCE0W3wayhX/mnEEgzhDjOxbuS4WOxfc/H+EgRifE0iw/SKRBi2BkOWd0YXrWA
rtmh940mv8ce3rk2OWZK1n9hoisWBbHZ9C2J0AqNT7jZLyGDjIiA5O2uVukrrIig
L6MzBJhis0PYOl13qA4S8kKmP2iPHTTONoxGp3KbG/9lX+fRahN6suQiNHzYDRHV
9TY64vg4leQQHk3vBuVS+oCFBJXpwoUZAqkhnU7hrYe2OKgATXKNpnr8FZoEA69G
akEgjqnMs0Ysupvo1JPHq9UlUU9AMsnQbkS4ZTvzSh7YfzDtITcOvLLQhyyROkul
9nP02lLDFAHexXioi1edIWVpWNBOva7FfXj6cOFdiROczGICS2FA80IdJV5gG0KT
ogOkNsYT2TPI9W+42R2z+cQadB50xrgIQtRSRy0+q2UVeoeO+wq2idKL7O445kZl
xXT/h9Q58mbOzzJWcruIz16y1mZEiNy+WKQ0xjmGE2dW40D4RoOECabEUCnbj79x
k9q2ydFZsx/kz9DXknJs6Lt7WRhn25etfsTCv9sjsgo3e4kcqVNJWkp/4obywt2I
LYi0gb+jS2CCbPIFZ5ebPqi0hQPK3oY9PkLLIkcVy6f1VMykEYA9CqAyswtglm4Z
Y2fg+x4zLFaXhjyjY28UNtunkVQOzqJonczKOsiCvjhE+uovxPn+yXvTHI4m5i/D
Pcas5tEaZhdA11tKag5NLzocRtT8MC/jyU3S4UUo4ijQjhX8/eGrLmThvzORYtrP
MGynRG+C5zzKOK0G9omAqEfCEvu2PDXn6yx1x45I+7EQG8BTkF4NixMD8OThnLSE
WXuiWNTWyljTEC83BtxLGcAqD8h9ZzNRvg2Sg70/0FiNNZFZ6X2CGNeuwPMpL90w
Y80iI+fDxdWd3DsiJuAFHkvlEXEtVdU3OzbeZMD1SHN952qsaJimiafDzvHf1pgP
Fq8nScv+xojYA8trrkz9ka4B/vGr3wWgRqzfkIUTnU1uNK2BICiUIAlhHe70qJ3P
zWSsuM9JP5Cwn+cUriU+CniGpv4fNuq3DMDv+DaO86wYXebEyJnfLxQhct7IFtTE
2rirXtP/eBREj/Doim3iqTl4VowhNN80DGqnPOv2+O4mAQwTeK1/WE0XYGR2SZe/
Cnu48rPhzCIrUGKmuxdMaeAQrw8iW+CVE0N2fP1tg/h7NGTVpz5ZTPLfuuHgyxcs
zwEqIPXgt6s69m8YDpSiGEH9+c+CCUALQSZFow55gPgsHpFSbWrTy/g3U92lncm7
HLZL2om4KoF7k5/kX/TtQ9ZFemLWq4ShMjwuUsBM8imD3LaEgs5BybNk8dqPgAKS
SAN3lqw1ykspKLomXAHQQZVlmERDnroDuEqLglkqylGeV9RmMTi5RfodC1qsvreu
FEwsf2J+FOpIC3FKzU2x9cvwHk0k+joDPaWsXkmlne74jsZVkQGl+Nr+LTxdLgoM
66+Puh+ohBYcjl5CwTXUvp2HKF4YhiWmc+op/GtxDgq2nbNl6K/dt8FcgS0t8u7+
0c1ZRvY09HLebjM07PodRyvR/cUxR7acLOhgt8Jl+NKvDhS66/KVC1d/65ubauIE
aeOlK7uvqmsuh9xvr3/8Cslkvj9DXtcEF08Ardd53vLKrRNSNow2ZR9BG7KxWluu
N78xWOQHJk28+N6vpy150LxLvvpXjwyFQRVlzNaE/7JSKkZ3trxOHMiHKsWC46Sx
lzQ/u83lMQQ4kblJWwbA2tNpC3gXbDJzBZ/rXnj5aQ/XbyQZkO8suxrgphcKGlsV
5YQ03zmd1ShydjPp2KuyfmlbN79gz3sI59TBQCcstmy993Tl5ww3QfloFSm3lQ3z
906DwlrOg+GNazMyRLLtN+YC7Tp/qZvqF0R9VL8rVLGOcDUsUUryfZ8xP9SwN+6P
JMuUn+R5IjukonMmXG0+tByphRYM2AdqmYCw/Rl3ww9/gC19CMpMI3v9rrDbW0VH
/F7Ewu98zmVw5FlG8qDV57jQpbicgfTiTwGHBuWv1KVrIMvCGsf9gXFDG7rY2Rm+
J2xX9SNmOFm/lV3yC2JoDtsjCxCf+l0jEGvGrS/W6CmrosHFzhFKP8bv6fZA579t
yFqgQwkLNFxF77JRQ5VlwiCvodqRjQinfRfFVg1lPfiJqdconriFPMFp0T42Ua0e
kGUEsw046L/GCayKiQ51vbkrg9E8pMeoyFQMz8KgXGOXH5iX6oS+uc6LGczpvG0P
5Zp1kcs5P7qAyqzIc1GaDr+dOrKuhsrFT4PzEGg9/VT+BFz98xgavnCvv4X4mf0m
9FFKuN44QCfzrsrqCRKUZL5c4GmQzLgVW4osjmbkBMHHL5eBYRJ18KDmacbGXdsR
bocIbGh2HcXF37orY7rey72IDjfjXtYOfQaZ90rvj/nx8mWVsLTUUHiEqj8JnjVy
pkoYj5DKf4G6q8oI9nclxiI5W7XeMlqSDMyKS4dUHejLM7JuBq/WCasfYb2PY9Bt
DUkszsTL2QOfTQVPUUjXmJR32GUZQIx9i9QIXZ0nHY2WDloZlsSWL8qCSh5uP364
ls4AFE+dv+3IjgP8iGKFP3udSGpbVYZUm3mEz/oXUUi9nrVdgHk/XpCLEX6ayuei
xfz+BFQHCIKW00yDqyaEF6HfWKOZ9plZToKBnwoa9oIfPe2eEeBWsIbjvKmF5diQ
0gf6kU4x7SfHQlPh05cwZKC2v2CMJsodW6XjPU21M39GYv3qQcQjsXip0jvV2wuo
jPzlz6lLWAUxa5hK2J5Pz3ZSxS+OxP5RB8Tw97yVxe3BKGNR3UktaA37JVGRV/NT
AB8Clifj4U5UFg3Fu2F/mD13IXOv6nh17sUShN8T6cQVllXC7H8Twurnsiw1Wwyq
4TRYFdVojDI7aq/SJiVkn0DjRxw9qfU2e8+ygDdpSsgdfe3P9TKkHBgXUUPAVYmN
dL7bLnNsZaeGdpV+4MoIElXQ1hTIu1OQHBAt+cE8ZkK/GsoBJ1PEVXpBRQohWZMS
e6r9jNUF0BeiR60TFJ7Mu/E7Sd7ynv9d1IZ9Bcc/8isqBvBWY8xMUH/Byhvn6jC7
/wFmQsW+t0BRc60xLedxiiq5qNcwU5JCfwT5URRBAQf1I9q8yPAaPD4p2XeZLUDo
UBPR2YgzyOGSWBTqqcuFpv2fmLZI9K7GjIowPsTCaY5uo68Qrz1GFKfxjA0KOtUf
FVyZyVCF2BnFvXtSUEvE9s+bA5TDTHhtQh7YAoml7Z2J647XwdOpnhGcWDbFyOct
tUmSbLpDtViBptlKM+o16RPpSbia0ZQt69jlgmBwXKO3qDfVGWyUc72kq+xX8309
L2IdfZ3Zl/uscn1Gcg76bgIi2DyR3+F4l9CumfaAJ5P3TYYU4GAjynCO0wuFc8A8
6vgQ1gqfvaiSPWbv0VRLyifovc6PQQkD1ZKw+xnXlth0E55Jm1rUn6XKIjTRzMV9
TYfHBcQ8QLOPSf1T6jj5x+924SQhy4HrhYzFed3BJSDApoKJgdgsbhCI8wI7KGtz
Pi6j3nEyzdgVFQFtlwOVYjxh06kpAD+A6cd/CdT79aQdw4+bvgel0wWOwmpHFwJO
URv04619qz8gTmJVr3IyzSTgRNdYjYV3TZVsstNdGYLWDQELJKxBaHjd8KEY9MTf
6AhhQFeiQXw+eQJB38xBdbut/tsUcjSMINjzIUobkDuiLuTxBlsDTS3l92yVcTqS
O3OPCVw113lIiwpAEWLpWPf5tlHKm0HVSgwl57ev4lshpJbk+RMVO1D059tgsXNV
dBSnvzcabMAps2nduvGbc5DjdCY3htlSgJtAad8qZVYxc/AeifV9StJ1Ygz7n4xp
SEnXqVBeFCMF6wDnCBpTS3T/RFygQs1+8FNB5g9ZMOhWB7/p0d3ME8X9IZoPRyWZ
8EiZud8iB/hLi4Fw7JELmiuJ/PKO9g23NCjLhbFJqo87qgTtuS+jEGJJVIn/Twct
dH+woL7k+avmyU3X29fT7o1ZLTQsrJpMSUcjq+EyQJ1T9Nbx6EUWdaiWgadhhtAP
6KOQpGd2FpZ/YND75EBdlHiFsBycD8DRgwInPx2mUzbGTaDHL5N6CwYj7ZJ2WtM8
xS8hKwRyVaKPnCoqvz+hiKj5naHAghcK2sE/QygoQC9sCXlWIhVxA454HYcM0uv3
7IS5PRr/7ly+nAzG4c/Wgv5Su36jsdYAkeSMCbg6i93YFdFaIAagMlXqr9cv6nag
uRVVagJSbOrUNMaj1oHHtSnLxnf7VvwtejoHng6Bl/5UuRczxOQuKb8QMj0vBZGV
eznc5NAfNzxJNrx6hkfX4B7yr0hm3fOYVqCZc7oqPO3VX52FL9qeDecpUIDtHPAD
YdBcuYbi8vhH48JFVMrFa4Gkz2cCIIzpiNOa6dBOdv07JXOiy6vBOVWavAL/cRlk
PdB/MRL2whX0nCVNp+J4QcHnAWU7OrBmY/imyJ+xNpASH1LPckPiziNZ2yxkcwsF
JZ42moSulQ1OiOAyRsmK2r4bsHErEWrpwsg1y6SCgkgLAbpvid7DV0yuozfRCOa0
aIAgEL5O+UZHF2Gcq1k79VMauLz1ywCoPX9HM5zv686MQ23wqiFo8fF9Nu+T+/SL
wdSYzUg7WDOGFvp3Gtlyvw8uFIPIh3Jbv0MmyYal+sy9BOM4+qOHMI/vWSdFMqpa
`pragma protect end_protected
