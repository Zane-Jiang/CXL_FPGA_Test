// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
AIvZO6bR/MEOr03uM2K4OScsM2QUcTOe/sZsvm2AERV6UFSZKlxqucgoQ03TNGCL
Y21uTI4zUiDaYVJyoo4oSml25vchLdCJHRTc63MrAOefRIRmnEOs2P9p5ji63pbL
i99sJ4s3d7F0wHUvt+iHWOdzn+le7kTCSc2Bz08GuEQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1328 )
`pragma protect data_block
89exJ2uwU9xM9sL7AKoXV36ASZ7m/HHsI8S9wpXTZJZcSGvFsv0dIJ8JXpkC5ILO
szSyOFImZZXftAj25PiUC0lP1Y4HjGeXv7CkAVpDnIL+FFlOoSm60kZEdppmmbnE
/9COFKYnTPqZ3fdFZT99+nVmNfwPnK7Fz+Qr98doNhMUpa2YWPDilurmi8zo/jc5
wfzvdLx3VPlZE3BDTOZ94DZwHNv7VEkX6hOp8/Z+ZVgFD3dSSl2w2o+MNVX2ym78
NPq3P2h84cGpm8N2Itxeul+kOqTic8ykivja7IGhYHPOcYlx8M35tZu42hDa5fQf
ra6MQrWYdfgiuM62ha/C9YC4jikHKT0/BUmyoeQxsBWVxmYCfxyZRAJvjMr1Aujb
K2Hi1AvJqpL4mAlIsGRtALxgujsdJIfG9crrMEHpalMEmyT1BxEo24QzTKsZ4Rqv
fcYUaMIESVJlZvlEFGfDj4g451GBhsctbZjTUhcvVGEtOlk7fPQ4+bonXV9X/6zi
IW8o/c9NSYGzSPxL1BBK64gC8vmNbGE0V8yTyHFnPBFaardZKb0JeEysnJz9L/30
x/4SPHE7lJBVwWsdlmWGQcQBH+oli3OgKo2g7aply9Qqe14l+J+E+ZKsaRp80OEk
LL7tOYspjKarMnl/4j7qfLNEf+HEEEMNt7zJt3fdrY9mAoe8qRlNTF2LOZZUF05r
kPZJZ7C4cDTDRlHz9All/Yq5R9kpAdXEJVStO1f5eBsvoXVQDEHcnB4Kwm6vMBdI
rMZdA1OPv1XIWnB/7dbFBv/OVdRtrMsN1fHEYg52m1k+Zr1OuCbYCF7M+sJcwmtC
vco46Xi/3ZnWlY0CN+wQRtiqXUwOPoXzEmwa3muVcmekGQ8E/83LBoWO5eXjQUvp
cp8B/9yeQRkJXl+pJJkTz6ulPDmCaesq10SFh+EAR0LaEw8Wc9l+qgG6e5os9C68
+IoxClRQd96xGtM8nqXJEfpzXeCOGO7M6mR6WYd3z3jWskLPZfAR515RH/7pdhxc
r/+PhwAMmliIVeRx9VhZhZQx2v29Q+ZPJgh5c+FXiFyqUx/bfL4DEbQou+6PB5Np
1T1NNanIboyHNvojDPcESVU62qqTIT1tOMexWhEz1hQOwQrKujhGlRjiBLd5uD6S
wbZByQ+l9AgV5MhH6V9s8tNqDTTbQSQrZjlX7aTvqimenbLMfiaqWXBfcK27/fmG
AJKVcoLNihCh0JvkJNSHqVPBzUCZ46qo54wPtrJPUUIwq66ot8soTZeLeZP3fDNP
WpYr2FVSU9DSCVVa7ovhI1v9SY+XgVACuY1LMYh42PsODbpK7jDQLiJyLEIc0ROt
B4fSqHYWyX2TOUZ+J5hr+ZMxaBqCjxk0CvfVmgZubACX9TA4rP1F4UR7g4uuYT3p
cQ0QChHCuGiWpS6diTkta4eM9JXWD6Z0de9jaxTI9kNrkcgcp6zeP9EeHdBkv7Bl
kVBkFd7hoedxNRQebBCINjNmLNwi/7ee6ffnTddGxS0b/iH+Z/DruCVZghHtUh0T
wKcTwoYSFbLhqb1fU4f66v7sA9p1Dm1fgXMvmm38ONAg/Mh7UpVL4ju0qsw66h63
UT4M6OhKfVDU/p3n1uEAhJk9wQdeDUY51SjqALjhh+21VXiacUFEARQjphZGlgSz
lfxlPcAH1ei6VnZKJXgVHvk9DDR0p5/R3wz2vmdgixp1pTdMeqTY/1BBv9fd5TIs
k8UaBUKwoRoLdF5LlgF7i2la60Ylhcjjh5RHmlQc0uw=

`pragma protect end_protected
