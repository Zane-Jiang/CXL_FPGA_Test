// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
02KLSKQkj7n71VjJpaXV2YPdHzkWrXuyHlj8ON2RH9huB/cXtU4b0fACm7UJ
WNMAyfhAhTsfZAi3uynr9aL0ARUWzOuYjGdM1HGQ/Xffu0JU2OqiwPX+Ee5/
YMr0pKdpucbQJHivdeHZ0AyoADJ0znM4BUvfXLQi+xmXAO2enesUc4ELjnnV
1DuAw2eisq4gECgJHkdVSkal8JEGl5ZAplnpLmHmXmrRAxDI2KJSXKcCAlQ5
XReiE7IEtGpvIIy/pAOPIdO8cAWL17IKOfAbQrsLisyg7qSBYLYe21Clfs2L
4X47kkdTbk5smBD8uFa3saD2D+LgxjL3MROUZubLNg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IcRcn+bTkzx+Sq+KsgebeusUKywjooaP8r6/OAuMf0fwCXWp9JQKbgyMPvfJ
/xOzf2E9X0olQ6yxRheRqV4pRKO/rGwSNhUSioNJbShkBhYopu62BhbcgELG
Y+ggq4lP3Tklg2GWgf0p7PUFuPA94vxvPbJ4ARoHMP/lE/pE0VbmTKpYgJDJ
ljqQ+Emre6csmuAVwA7BxJGZOMoVMW77YrElMXRdT8zHnYJgeqFFN3eM4l2c
+pwk4avFcVKSuJbB6BJmBgUjMsMjTcXaNSBvtHzAmsDaZEkgfcyGM9a6759g
VWvP3NTcLJmpzFqWMIAZhUXLkj2fH5A6+O9tPrXeJg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C8M7WSt5fuF3p7rZqknBZ6o5kneUZ1U9AD5c38dMX9wCJjJEmOch/oZql1fv
VRsBQcOVSBM6j0FsNd1/3R18egNmpS6yoOEB+FC18n7JtGR2rrJMJnKM5gUK
E6xeHfw137XtYIXD/i76hFzBWt2uGYQ/BfHJgNzEq0gaxVOqwe8AGajmxc6K
WuKISjnpq/uqveZkfMYi6YO4MU7MOFZui1nWo5VmGoRTqP/0K37Huhlw+PcL
O2ZJPKK2ph7Pyn8JDf5JrSdmOCj97e8e24feQ/0rEcA86uidEhNvYzucBKq0
paSnh2xpke/Rb2cp2s5tMWfac+kvruXp6eVuPqDcWQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gcBaSSgQh+XdYaCXp321iVYn0vxxeVOkBSm9xH4figM71g4ibJdhjTwMgMuB
fcTDSJtQkARRPnTxBegYlWuHwmt7svCCxdk0FuiKqb2KbZ8H5Exs5JHYSi42
JlYW5j6AhzrrHerEt78aOitmWm1sTBbazE5t2Mn93U7s6/yKLCk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ncKlDAEgTx2lBBiriIVz3dtlgFvToFrNVWK4PkjJfoO4CKBne8oFMQlRI09G
gU/fzvEITbKR6yHZAk9j4V21RIEybNwMUPP28zPPzQGsmczLtTAdQCICy7mM
moiHBMDXojuev8PcGtjlVqnOWdwfQu0v/hPrrLxXeFBq5bUhcI43vXXyjoiX
jYfgRCIsEeogrvzSLTcJpGUbv5JnXjWv50Prbb7RKM8k16hanRjZN6eSEeNa
H0oW/2eM2W2VreIz5IbKcLC0QSV45Z3XL+XFd+0VwTvWcHKee5d2OTS0qL7A
Sug+rmu/KqTHdPdoHs3VYnZwvHeOodTr1F8cCD2/hPs2P7qp4uEM707sulSM
/uF6ba0LQX4B0to3U0MXwMB2mOCPJRUaxRX9oMCF8bhkfkqKVp83QEt7pq6G
DUm2Wqc7R7r0lz1+R5+ukhT5hcYuG9+WG5rb2zmIBXdh++U3eN2jzJIooNMo
Gqs09D+fR2OVj/UAlj4Fuf6l36vvgdwh


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ht56T5POQZNaLxdImsKcPG/XT3P6oAeD6utisBsL8ElDY/dQmMrPWqkjjBpx
P2j9zdasoqaqqsdgBh2FPapmtqUrA1ewm2RDT6Mou+URXh8LoqwmBVp96xKJ
gdD+j4ggDUwEifYCqLnfMEBYDP/mWgmSpMJXyWIGWbZIzlwxzy8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uxkSNVpi8NMQgSU5DwdbpRsv8U+XkwHS9nY1oMaEqVdkxW708ncc3o9f+032
A1kxBbQOymuhM7bRZx5sj1Hr5W+/Tgipu4qiOIRFM0/pL3sm//hJb3HY+jXV
lcT1QwltOBIISVx+SdbnHG29vIIw0i2bbffgM2Pzx6q7B0Ickv4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1216)
`pragma protect data_block
X8rSiJK/8DrUe+hHMstRhQLTdS9kAhvm0IsuZFYnqPsWzI4zxDoAGF3bxwpr
SQaY+CNgyjqA0i16pwkBfDN3UV1aqtcki+h6g8CXcPU7i0hWm0jqbh99zmEZ
i0IfE4slD7LnANI6oo5xcghm7DaEjGPkBTIG5KzaHddMyxp0NMq/iE5Ta83C
jdd/FNzxEqJrJMmFEM5B+k14ibqXe1jmifqTYLBE9vS2kjyuqvZ06KSiZs+N
GT0jDn7DT2QmKPJB+hgqt4OYs57MnzJzGuIzq6pXrogboTmW5ahp4I/ZA5ds
/3hdVGzAo+12s+ArmjMOrcksy4jqxBF1AdqSq68eTXZyqDgwyQ7pkoMjL4tE
zvTm4kyaqbchCnCQ/UNkktSnXbWlXVzKxx6GXGkRy2jMdNQTEh0MTEmH08ff
+2A5rA+/rdQAk3y1DYw2VA6ujlreDy4G7fooEInrcU5QlPpqneAEGhbekR4T
4yHj41+Gk81r3SJmg9lnSpI+jLIG4PDwRJOT1Z9jesAZ9rlwEQBxYGVl8cWY
o5DioMBsLnYMN+2lS0cY5+AloLkphSZvdRgnk6GqTcgfE7ukm48hL35yhqnt
iNDHyKyFluAMOb54U9BEdR9MHlm1IStRJwA7xYdyVYt1QeAbZX8ydIsd9Dox
AHdXGQ75WI/onar9Fp1D77phI6By6Cf2uVZIaF/jFIP1+U/K22Pv5t1aDeO/
d/SyOsIJXiDp/dcQVEdtvBNIJYDF9a2k2mOsr6aW0xecaoAGMZzmD9LgaS1t
8/HJSrX6sxfLHSacxns+kLvOfT5CyhRr/o7U8xF527eZZfsPhnGS5psEj5sB
+yBwRl4D4M2X3iKOfKlJAT7OBaaU4HzmBwvjZ0GeijvY/D+Q7VPOrmoqRhfF
04jGyA5bqvBYmZjbOiptQwzzwjxys203I4FLKwHOqurEhwNBj3D688G83ULl
vOYCbmW/jHgft8TrqL+AL+84PlUtFdOcfdzWq3ZFf7sOwvkohzm8bGRQNfCv
DOyzJAy2VNDx0TR3JE5LShRDn/gGdMefTeMN/a4oCX8LvN7uaFxWebCcSwPm
SQkQQDvkGdpxrd65hURp81OEPqPJDDpBbuPqeghnhomdInqS0JYVbn14Z9qV
E0S+Wi+pPnEkF/+289VFgupQQMyVEdlqrlpNUBMoSung2779SMd1467kZaxu
XGbTPcY2P+WgL+OMB7d89dVTG36bl+5aD09IMbqi4qXkg7bfY3DIWA1ZTb4T
uhBZFz7Sk/yaAmqhOKEQaNE60s+FzeHYa/SMumbDfW7iJJ8md5gAHlj1lW8D
2kp0/A/Uvhsf1vwHPBiNH0ew7f5uutjf8HEXZWIkFBo7HfP5OG/KG4nJco5+
Ft/9Lpmzf9zgGaly3PY3zMAVUioc4cUvwnYUXd0dOsZvR9AVXwOasAUmzAAR
WBI2d7k8+zv1KcVvsfT4o85dwAkhDaQGFF3waFjpA/rK+HLtrNrdO2kJqXYb
WKHhKx31WGmtEnUXL2yp9Lz/3+9D/EZ3m/oJFflrkPILNC2M7T680E90hcls
DSRqHRYQZ3FONPSdbXulIu2Eor+bnZisyM6xspN5ii7vkgA4HhFKRRCnEaEX
VQ==

`pragma protect end_protected
