// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
uUEqXscGIsFxryBwrS0d0NZHjlgC7rpIfq+MqXdQMfmRT3FZRcwAK1qQ//G1g9Zp
oqEb3f4DL3n6LNaJFxZn8k2qc0n0nAYtNHE19UE600H+SiN0TGJwwuOUIT1/FztG
TT+TktHtVKoZ3mYu5EoYI4K0QVoSJM1KGyRmQS4jXv4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 38896 )
`pragma protect data_block
CYTK7ap/+NPGT9MwIwnd/ypLiHJu4+SeUsNJKeIeI6lZ6lbcshU4aqwMZDmf/nFJ
UhiwAjFplnP5U5ke+h8GvZLTIWbbC6/znjZCp8EqV5HBkXUgvsBoNp8cT3HP+sgD
YhDqy4la9HHkF3XMqKxSKZRDSql5BIEM08eWrdVbX4QjYomt5yRuCdlaXSTVMbQe
AmGGNpqJq8FHwZ1lHyH+kmBchhJ2++vuwNFNGJa3+k9p2lGoSu8XgYVjwncZdn/o
+06HelSjskGxtNRA1PBSdpZV9+AQpIpQtEkTQ51TnKqDwBemBdh+4CzReM7v/UDV
itvA8HJkajOSLfV8qA5zFTJ00i0ltfNcCwS6GdwNVawb6IKy43w7IzuStTZH+93d
8fNTNEmsv9HJfPPHgSdC5qPpGiHl6kUzeabiPFbh6OkFFRHuMHX/l9TKY+ZaXttN
Kb8YYg7tTasf326UE0hJVhglSegc9mrS1KU0w8Jjd8ZqOIp8GAM8zJDvFVS8Hcz5
nVcRyHDzmQO3dHpT3pzjov8naS4EOpPOIINlrXmEJ9P+pdTWZL7kixX0nSGA8F9A
E5kRnMlcC9t+b2Q7GQB1THlLnskfP0ZKeuV5e8N3Dt9Tnzv/gQC2Ek3eGDSrchrm
5bngkg9E813j8ZXtOSph+sY9PAh3zfFxizDhu+eq7t6AYL4Lwb915uQdoPESOEU0
AcrtSgcWqfYU8FXe/P/jrLU4RZIbSpPENU+WW2voTTG2PpIXB+PDh4o+5VtWF6v6
yX6uTDBdM+rzfxXyYITj932YL4h+XVQT8k26+0KfXXfGJqD1xw8dhkAwgRInGRJM
/ZZDMifekcwCJq1jt5rCVbBxZFDPrP88MXK4Y+MFAVRhb2LQBr+z7pz6XHKKTq5g
E71KsxMUPP7Ez1ytdy/BHbTNI4xAjVnkT8bPW0+30Feu0mg+PNs2XnBXipTawpgk
HfIvxXlEjytWH/5YuZ+Qi2Al97lvimNY3EdvR1ThGvzz1h1pEP1G5h8OPW7vxgtb
kb1++hS/IGEHYdu9pT23DxxHbLL+BqmIji6MVww4MJ2wEPv9aNoi/3qW6IXwaU5X
BWgbEEGQLtsu4aT6pCG1V1CIECFkvVqDsFMNI3llSej2f138UuciimJqPthpvcMF
PFRAxSyoofCucwmxCKhN4sZA0PtpDF2rACVlU+b7/NKW3iyVH1ES5NKaRhdLq04V
bNSEThuev2lRF+nkperN4DvC63/YkX2bBi+qF8Epl7pNcfAKuXWKsZsHhNAW/eaK
57fMJ6tRbJ4gtrMmYqQ/tD12eORgom4hRoWr6AdEJIT5xm7PotxbK5QLT9dDJKPI
SeSuKcPtej7io//7Ecciib10OaHi7dVCZQK5DQhj2raSQsrCQPraN9jt3WtVYAj6
PFXQlEPVl7lUNKlWEOVsgI1c2F785Diij8KHBac8q0OfYPfXFOojQ9bG/IvAGSpr
h0qjZ0uWYRLIC6HjOryPf8/TGJPQNJ1OX/tGBVD/FR16tf5xLqiis28rEPtIdzdh
7fap0SZ0S2CzpXw1FOVLks76Z7PlhcusoV5EsJHS4bClV+SdZXP4/ODIjKZz+0bD
AYVcBEVY9wQRLAcgq3I0cAW/XLFBTtgbsJoEeh4SWDlk+bBmKvNSYyLyaBZkIxkG
05pkfAEwiui1rmzOt/NCoaEOTQXJUoPK/xCtcxI9TA6BOCM/4of9j8BGXXX/P6cF
1+cWN2yeLkWGmJmSc2feH178jVMwflrz+H/FEZa2+us0VvbfoDGBvzGYp75U665p
EJOtn13T+qxKgQa23hKMfrFw8DcaESjKPOwcvpsbohFpck0v7QasbePQyif/vgzx
50hi6bgx6+XzB3vcJ9XGa0LtkWEJJjm8kynhdMD5banEQUlC1Djc5hPpOo1F+2/M
pHsUiExKFAIQmdTy1y+WftASP4b2kj9jIhMKYw9ZcLuFBQ/e8UgVdf/GH5UnP8S5
R/GspjZppUzjSDraZ9d9J7bZXxnt71SEKmwBRg/HL9EaKttTxwyqwXDFzCovfe4V
4NffRcZWXOeWkf6RDv6xNgh4GqgDbYN/NJNmm7Cj7qw7lXe5gF7K9NT2tlnHGHUh
EQgZ4+/jlJu4U8XUnLB08Hx5db6ATbMIYPUOIKzUBpHG2Chc8o7wrbrsRgCOAW41
v4V/p6lXmwVVMW+mpIaxuxncsk2uedJuRpDADQtI3hQpD8qjU7kDgQzh8GmxZN94
bmotD4REQBbZYYQmpgROrV5AW492ZkZDzQkKDLeHx1I1KkoeZfKMkWRgfbt+8ovH
OCuCQyTJ0HBwlYvOfyviHK10W6kGNEpAk8sdUwIL1ddG4Nk9deOsV7EyZyytHl0z
q1F4IPOHsCg0xn+XyeiALaoo/xQsP0hC397CkB3eRn9l+j7Qmc13w4VLhiKWE1Pe
FkJwjaLFxMb5tqdbAXsJ1/QcuspnO1N8Z9Q22LznbYraVfG2f2xEHcAVUIO58zX0
aYofk/vKiubduQ6C76GfQPkKBTkTmch5AbDWV/kGXCEzzUoGcMl/knvvcWyNfu5p
X3ZuYaNIPNQBpyFKIvJ9l6oXVnVOwEJxq/9WCU9FHH3KQOu1LiWw/qbjvMT2RwDp
4WCj3Gkz7OwWTdTD9sPxu/0LB1d77K6g6gn1qFNqK/G2SByHXZYOzlCsXULejOwg
GZH07xY3AopVRZpoS3WAO62QUjIyEc4Eu1DqWxfbUm7xexhsZsb67ccxBqv49Vnu
h0Fd0J4bEn0fxRaFzIaWi0f7gX9IzYw0mFoiXpzGzUcI94wrq3m9gZn3M6LW+M79
FaOmByP9WhjCt7ubHCyckxAd8hSp1Kw+4/5/MouqX6ssMvEu8U/k1d5m+qlO9Sgq
wCXHzK+KWjVetZCVvkciWhAdv48JTwm1X/+GKG/taZIgqUYsTdVIzzJvWNimr/eA
AGkQ9lU9fn9TBt7Xpu6P9peWYnPyjbz6UtocX2kL03Czp/lZy7d2RgTW6/neRB0S
hfjgaoMkXF9LpoSUJmjxxvnufxCyE1ze8gH7b4avuKsHX93AQfAO5ldVqV+Hqxjw
9KDlw1hllDpC42GjATtUCRjAvzPDvKi+K+H5CdpR9Jvf0Nr8DO5alTgGVWTVsD2J
NQwU4CatQYYouoD+Z9gMG83CAgKLLkm9JO9nUjP/4hFQ1Rwl4FDhW14sR/IBJlkC
Bo1taFABXkiV7ndLS00nD/BKgvqZWZvFvLdLi9Zlb5xphx851Vgiq2XfiCNTxlNA
9FQFP26Jh4GaoJCWMVqSEh7Pl3tMil4oPIpAwbyekm13LGdNgXHh35VmjGdfIkaU
gzXr0+Br5tnNgj8reEo23nafvk2s30NzBxfA7QCkgpXSd4Z6xFy6d1zLduCYtgJS
kVMlrS4keSNmRg+mqUgbgggYDnqMTWFerb6K7aTuQQN8X5/RSHkH09FN7KQdVlv1
cBXL5cXCOjzPHtB7fotT45WS2hAd5byJoKdozZMqqg07HGuMNAkJayWWSypoJ25W
EU0btMbbT55lVDzSATYJf6EMEueEjK/LNRfEwBeKXF0rPgbTmmDtXifwaORe2XmX
kH3hm0e8cUlwljEky1ddt/8LEAVV0/Bm982BLVDwBVL0EiLiuNNxV9P2XUO+3yPU
EP0r1RX/DKX9l1BxZPsjBUXI5E/w8onTP0lsx4YR8PB1ETM3IkRgvo9WeR2/Y+88
hKg0XZ5ku3xNjnc+ILZ0w2xGXvnJ9k979Mc9HGpDrTchqhO7k/OX2oV2YmeshkWU
G1j0QFyi6rs3mfkNE8Pi4TWYvAWY55UTKW20rdV0TDFSrW16Z3/fKrc97/GFyQMh
LLkMIFBEQdJgX47p9OUDLXb0q5uYUrRjZFywOLXKxVhTx0ICyYhT/3WhI4rkb8u+
QHK/n68OTaOc3fCcuX91emoLPkQYA1D51uSPoZBnHXOxD2x9ABzt3c1UmSciy3rv
4+ghRf8SW0i33MgVJimzM4L/IciB49Wnm+45gX3XPqndqz1NMkX5i/FZ2/ffeCI9
pOrTN670HqfAszjIGcacUZ+SJ2lrxrAj12GUC+E6uDICoJSSUWkxq6aE8g+cMsXO
Ht5Cc1yCPYkudbhS108CQ4R/N53U1ovzvRktN5Nxl7GU4fXkdYtVZapJgqGyl7+V
q0zrVoiqgXnVrgMoe+wRIYaXGi51+S7C90lq9imX3ZsI7uSuUUfOFqNs2gVodpmi
0heg3fhPMJS1q6bXLhkDJHGMPCt4hmvostoqW5Z5NPlFP8IdkzUVTcSd12w0/mZL
M7rRhFyp/OkipBf5KmzOKBO1T+6uxD/ClUCeEh6GflOf2zAnuRRvKoBFYmMxVrwQ
bhikS5UdKuZX7k4djAg58IMbxuNfIUH9fGQlPiqadmA0k00HIMuRBskvzmGoObUs
wf3SWtXxgiPsQo3iQx3glbpXmrK8/ccVtIt60S68qYLdsczk4gXR42HgEjKgye16
sQKzEzTSKAiooDEtvLFwaijylSoqdcWCDbrUdTMDLYX2Af37x/ZBOcoBi4VsKAP7
rFtEGZjYanQYQcBQpYegQ4aImLGHUyambOmtHZgIxHFNw0nPEuvpfmoz5ftAHEr+
UVOpcEN/pfzA3AR1Az4oaZLGJVyErvhdI1EQSmKAg87F23lWE2sYIRZeJRba1w1Q
lHoi1hT21O/rLgxH2ow+Aya2tGH9ywWcO92kWCBOMr5daLa78vHZ0XK7Gl/kzqDX
CifREoF27LmERtHPYW2f1APx1bGBAJN1vzXICV9EQjZC3RwJZoUVr6MYWgqQ7ktR
OEC+tu7Q4EDIdYytr4hcM1VTnKHpxbjTGs2suu6dPJCSJv0ikW4hmLt/DDXiC9rb
36w+GIfQ4hPylfeKgPCN1lZjTssd4YZTozkrZsYMxeLG5g/gGzVszWDGVuvsDigd
Tvz9FuaQWKQOTEHcZm3wAJRnknK3Ts8oZEA+mDSQHDhNZ9EXrlj1o/yLl33l8M0e
Lsko2RZHd/T6eYwIStX1Iio/ebuw5SQveFT0zKqDtlULG1e/sU/57+NNbr6/aNGq
JiW/f/hk6ddft9oWlFMv6OOtz1IIPvE5qavZNgL9ZKpuIxmKFPN1Xa9cLlswJ57U
x0u1BFy/Lq6RethcYRZ5bTI7GGJSYXxEImKx8pwMXODB+/F9xx3TYgBuTJyuYHmB
ghrecGX0A8LJzFa1+VU2UP5BjIZq6IdaTnh037z2iz7qW8glMT9USz2xQjvLijiX
20Qr3eQdL022ByO5KqGr3K15aGH95kzL7xyBAR/Eo17L+84CYtGkrGoliKAScF8J
63CRVSW3NiTYHHIbCIBjKKIpUQhT4/uLT3NadqX4UHm5clsag4HNQe0caaKHX5kb
E3ozKF5dr+cHGLmi7nAixim1tL0pqjT7UP8KaozA+R4UEE4++9btRquOv1TVLA/x
Li2ST9kjw4+OBlieSck4OL5bfopGpjWFUXuf8Frl3k6iK/aeQvO6HO8knke4XH3O
RJYBVlWuZm+tGwLXxqm/sJxsZmut82vXSn++Ra4VnyRi9j+WDsD1ME7UHpRqKhhE
k3VyilZOF5NVCOwxjqZH1CxMSUtQAk6tKl32IoBji916JMVlvOXi+yBW43xKqyx/
Fl18o7opTGp4l93fZe0MHnBs4Mz+p85y7qYSlagPB74xTucZkss1NDRxE+R71Kte
oLZsGFqGCaK5D10x4oeZe2nO36jbXIbzKtLsTvsax/S7HeQHxrPywHPy9Lu+vIBA
Rb1aBckY0/05TH5FYg219oH+qzgL9vDkncM2eFS8PEkjcF+bSc3Ayazevn7XcJNO
NZpE17hv+4tl+qhSeyLvA7Io7S3BvpgJsKfBVORJ67WwlcahixsnNRlrtJqtbf7y
okinVEepbv7HZR+Zhb1eSR62srarFeMFwHYFhkQA59KkqCr+1PPaEhZfDk4V20kI
FZYYwn2XvlgomnDbEq4W05tnRZowcMXVvPGIPDrcYXIVxL28bL/iAi+AfdVk8l8a
RMKz5S33gLCi9TMDwf/rl99KkJaaiZDgWYN2L7Cf5S6lHpzxo6EzmSRRnKrPKpnq
78HGzZ8hlzHdon6Swlr7ifq3uCYIQvoUsXhx4dz4VYJaVRaXReHZlHREHU4elMp2
t1sxNnLcX3ievmY+g5uH56cydNLWvxMv2QkwjTkvf480wSz7ash+jL+FIX0BYO7t
2juqMMDWr2uR7BjbDHlX3X7kB8EwKogzsgJQC6WcpX/n76PL5BCM87YAzeZP0aQK
grrqeTeRn5Qpz8Y7vnJtjeP2RrfhlILd59I9pZiIEoxIlPkKvbPali9UIlvUFY7t
p83BtIPnsOrxelvs9EWMo0TqvFl6/7a96B/uvPWZlW4FycWy6QQpCoetx/q2Llgl
As6Lms0IR/328rSJ0QVTk1FHmQms9vutweEZNaANhGxjJOIbILso1ffzM9nM5zgj
ZsgS+8a6lSns4P3Rz3m7JP5Ul5D4lKh7LnsiVv+WA2uZpTQ83opPgEG8ZC5EmAEk
az/W8Uz8DevxH9QCTSPHjIzH9k1je+mjtrwNtXn/nIr1/vYbx09fJaa4Lcklxdi2
eWJEHWlwkJ3zomBaLw0LunQ8wb4lddrkzySQ1dS9UEPZ25Wp8XLyUPRBPEhIW96D
1a1GD1IoOw4fW/jyOoGwYMCQhMY/5tWT5rQWgtYzx5kxxb1Z97KriZ8KLSWpoRCr
txHwRpE2JeH5BMwFbN2Rh5rUdpR+UIP3v5Lj5BIAo/J81q+6ZgppveKzJTMCw0aF
Llyk/kP+jHcr2Nyn6noyf9pcFdeiBBnrAY4k7S0IJI9M6WsEGE+Yxfww8xjpiXHT
K7Gy3+19SPp4+WtrXLdlHNCxxByF20FMYVnEcsbMYjLY9dgNHgPfkispp+rnfjov
qOoQXwHQbAv+LAmZN5fRDSXakRLkaE7G9rHRHE0qia8Ue1WnG2YvbO4/qFS1u2fW
0vaho4Z9miSHVwpPP/p9QgI8toG5Kivnkd/Cmr/3PB5ZjW5TkYo4dwSKjm5rFo/f
CbLLzUv1flDnnLvna1VU3QhnFrUNe5LvTVz/cSnc6XWMmgKwfdMk1dp9YRJSmj3U
1syjnli3BuZbxeVXgZWMGWy092ASOqdKsEs07VzlgIy8ny0FOR0XCCI0Xx7d0Ux6
uphFGhERtDFObySgFO+/Y3qEQ/3kGpQviRynbL833e5Se7BxhiC+FCqLCPzZ+aw2
AFEVCeRRr24Ky1QQCRCkPeFNlk3R98KwR4Gb1sOxOHn4mQ0pN6wxePY9FfBiN+V5
7oPDHSTk/ltDUuOKZtPt13x0/oBiA5wWZT8XAmM/w6k7qNBsSkEK6PS7v/l6LBI2
vDgvF011YinprFO6ITDCVcO+KjjbPPUsU8gq9uU8Rvsq3fvOhz6IWQBB6kEn4bKs
o+BZNdxt4/OgqdP6c/zL5ykTJedkp8Dlsak6766WevyApBm6mIyJ/THLg3osmjtG
PSV5GBz8o7Ke0Q7XMna+nKSG9mg+yw2AOkIn3aCjTGFrfcheR4AxTZvn8GiJFJwi
LRhzo6CPXMIyuREDiAQ+V6cABaPDD4JrsPNSspeMz8WmpmAwOOwMWqQpWvDTde3t
455hhA5nHHY5m+66Z1UeNMA9xMnupz44f7RoeZjWZYSjbIOld5G3x3pZxui6QKqv
EM1qxhgOuTlZjFAaSHV5iFQoVoX9NKRyP8a7hh1MTgJ4yGnPsVJsoSMCN/CNWInn
goWA8nmslLkLqtNnI1GpYk5nuO8vdbFWbuL3ERBVtLwDedtiGZ2qeR79idz0o482
oeHyGXz04sU/XkIIvaj0G/6amQ0Yl5DYLG8lBykeb3d62gYNclFO+AJBZ8TPMdPH
8qyvs4Avn2BekMtkVWrcJMHqo8urTBvhP6kzO7PLdVFE2BQatTrHpuMEj7Yne7So
UsW1uBtpxrvhHDIzwCtOPb6O+B6KOXlu5C8TGl/+VvgjiXjWqpzh5YKtZjD3McUo
g3PwQFUMsduzJ+C7MbSHgSnkSQJ1b3r9kEKz2CjbonIt0rTCxDFpMQbccyVG30YF
IHtM8d0gukq5eGRZi9/+PRIY5xtSfYftudVq9+5Hu8DSdhQ7YJ1CN/GqTL35CY6N
ngjcT5TgqGiFOoF4z0Dwy5/JAO3py4svp4m+1ty/OE8KxdvaaraPV2ZtJi1Hq97F
Gxj/Nns86N91dIJh2kt69GmR4OTIYyL5gU8wr0GfhJfUhrsD+GmNJST1JiVx/VP6
V8jQIAhMCcNPHO4mcTndgAjQswqURgJ5FvnrSgLRgSBtkY7maFR0W/rsiCmjt+TT
7P0+ao8WEbkgGEsIl1tb8vo5mSBeERnLsZ5pYByQCI3BSzUignclXx8cmVQPxBv0
fKVybXy2Fv5k8NjU80ZSxIB6tw6lMTFf6bDs4l0IpeKX3aECp7giW0fQ4NdFsuLu
wpupEiqzWdDtnRiW5uNrRSB4+96K/GlRmikFZyEltsgH5wqrKHP+Vw9VYtI/jAYj
5J7PTJQLA9tbiTicvxkw3bgXOh9ngEIbC6A3xAC0I8HZqEGxN7wTHsXBSQIkNBgQ
81hPpw4PjRHoYB403WKgAvtNDTGsSyAFP8GbV1xpoZKN1MuUAMHUwobSuk1wDyFP
EOomqyfztsihYsq5oo6mW1z56K70bL47pbx1HmJ6zQUcL0wTX4LONxIWF94yHHJC
2AQr1bbeLz3g/834z6N8Ogl+I5r5OEru7pNYdrzUIaO+2jAQmt1Jq024Lx75HHis
wJiYElX1Dg0QxdiqDL4xX1YmwIAdP/o9+G7YDsefCk4rKdHgqZs9Mi9CUSiSzl+u
aHWVgFIHMUuB7E9gPnqskcAUvrcvtI6y96ICjfyZoaXOsXT5X+xqq6C+/GnG6S5L
EHIEirpdW9vMKs5QxsTggrPUViyGBW/4tohPWB+SyVMv9//FiGwm7ix4z1ndBx08
Wed+OdI9f/dlRylm+QHgDlsNrzPiOFvaGcgmxYUqJFY6/Nmrzys4mffeTDBM/EcB
Fly2x0gfL4mR+TZOSGK6i2Q8CSe/O1Kh7kMnSpfrpjYBySqZ1ytldxVX+0HfXH2n
vQDC4LKXUO90iKgqPH8gscFeBDHeHGKXX+3eOKgW//fEP46irzWCN+X3pC+Csngf
d8a9GklSqikXyS3ZHbqPki78IVDzTGSTtu5ZR/LppSOwuGCcfVP8dacTiRgusLc4
KrUN1O07DTUJWJlGrzlQTfsELvhHmUE6W7FPkDHeVfCwIGcii+dRxFdbKS5cY2Vq
kHkpF2mjqn0SoyzGs+BNwDdQ8wApNynl/HH1KIY/eLvtzgVMZWU9ewW2bDeVX5Dt
keBKD6C+HYcuuu1NPuKlbusrnlq1vaY++ys3Hy+WLgLVvV9kRz5KBwqqNLEolb1J
ory4rNEs2qGzLW7ksBJHcVUAA2cMT3WIPQ/QJatwv1DJ9Sv2UcRWxx998dwajdm3
9mv+J9hn0z3LyZXSxBUaxx/NEmELoiyPDG/jgUxcmyCh/ei2I8H1U2tTB/XGb6w7
/JnF2FEQz1m4VveXKF2qg4lXN24IEWUTIxv4AOLyha/fJwIhLLVlql6EGsHlfwUj
IhhDoIfbSgn8GJflBpFUVSKfg4xRsgwKyeTwqTAXJig+KXr0nn4KI3Rk5gdJUeic
X3A2IK8Tq5N7TTjZFHK26RhOcO9G65/pKQP32Ao6yolngaknoDtTeiQMxQiSkJDp
jIbGJbG5K5beFzbv/dwbjq1hmoonJRuRabxbFdGuMsX6uKHvzRVhiL20FGv/OYlk
VsC5Q7dKBIX+ZS93y0ArN4+BvgJRdcn4HpzmHJR9CjckRP5CNnB8fDj12ynG+7Ui
xPWIzvc7XZiy96V8DX7DCsylirGiVABDtfINcOYPNqA5/oMtZC1fkaEUNogAQgiy
U8kzqBeBv7QKwYHa8Y3pv7SQujKJuTsUTdNPUB9uLb1ZHQOmmzEEJwticE4akaKK
kt3i8BXmRGfLrSrjI2u5nZxUSMpS+XNdYwuO6wYz88S5z/C4lml3kerfrhJPJJ3s
im5NHLHgRZR99KzhXYiYlly2vMUJDnW+ZCNdkjOqv0QFC7Zm5q578yT9NSKXQaDl
nQsaKVmmAewEA8pVCgICza+lx8mKSwfQ8npPRW6v4h64nQELQrDrt/W7SB/iO5+d
8vO04pqZu9MDr3Hsq7JX0hyiYhWZkWRwe0i55FxtJkbbc7Sv7QJWOQ6UmQkQdHKr
GaglncLAkXSf7hubT82he5BQsOPDcosyM+e/o+0spkXVXpCHCIev+w0egxsriY2E
U+WglcFjcXQ7/P/fWiWcG0wisRjjFgrtwz5eywIJJGaUgj7005+o+IFGTObjOgkt
Q12ud4SYKw1/zKjC++VrsgLJzHLbJXLcYHlnaqyK2lmayEjOS9yxKkz5U2+5Gr2I
zTKKwL7TLTZP75DP2iz+flv/5CUsyGi0cJQYK0d9SPGge+yQPUvocvhT5iW2WG2g
CO8Yljq8ihhIofdDWbrOTfXfktj4grueo328Pz2kqC9kN56da3fp/jvLaXTQcF1u
aRT4Hmf1pc3PU+BQpUDAjh5OFQNqZHLV+T52lRxaGI1YPRdgLXy7j/QoR3tZNMuo
L3+sTmBM5xVbDFUWdOu6mv2LLq6ci6Au4QrtYs/1v9jx+Jp86vz9a/cqQ3XL/KcW
7jnbFFHdHzGMhjxTKP/8WBpnLJtI8rsWnyO8aibrvBgErSA27eRpIAawEaBkgcQr
EpSTC7xDt0knhS91OT+KerzxgZ3vT8XAOqyShPS6O6httxzo80LEUcdaRLUfjF+F
TjVChvcOHqRg81ZLkY5yP6AdeCPC9cYBlQc48eCQwIkRiOEs0/6BA6QV49sUizHC
DJIm2D9I5nMslYX7Ik+2/1S0MI8wCJWbhtHxMVV7ASt7kQgdfrnJtep5pr9X1VCo
5jHcW8DCBAw41IpJuCpxIMQUL83S1UsVlyDMVvWFi0OS4gPjnnr8Wh6J1hMAOSd1
Wr0Q0s3QHj1jb5K5cVRi74DVnhkcw4GaQuj8kOBIU/7Av+v/Ya2r1RnnlD3z/eyI
+lc0w7wN+39J+1PTCWlgEPXFt0kQHUZQg30pi9rNgobnABRs0NS4tmmy6A00Tjoj
kDMoQn+FzE9gwJ+IkIH6s94k4M66tfjNIcOMqjOm5gUt32129/fib+q76nrKmYcS
O1HarpD0VfgFKso/qCSdw9xSYcd0IVnQA/rf5QhqPP8Kp1wqEVBOamxDTOQDpgDz
JYxntLua9XK6+0hL11xZ/Zn406wXorppnEXLjLseUZ+3cuWWWNo1cbMzQvn4V56d
Ef8Yv/6hxIovZXgZSjSuYwa7KnvtapABz8nM8jpzusfBWEudte7uHb1/fgIOcT7l
dEf7hsvoA/hVXGNLJkvCLkMiMJW1OCtPcDOb5TojGEz/jNNGxwVAxh/qSBR4a6f3
cPguP4YvaHC0iI/Lb87IA3h4uf21voh47JI3hhn9uexV2FR18X+J/GW95e1Ba09S
gjJ9FF8tNZg0BWNny3ELIawM/KI1RIvYtICTaqKx21Jl6Z+WTC9iqNHJAwBQ62KC
x8lVDPCuOzkY9sMHl2JOMFyT7TMZ6eYGuVzKT2QhAS2KL06YPw5/q7dVXj2+/s/4
o2GABWAVoENSXgi8I1K2PV5Rb21iOotRZ8MlsRQa84NBDOBDUzxZDH4dEn3EQUbG
UgH5FlPq44zKbt/OKNdWPhKZ4L3YcHm4dWnK8TgRfN3jettcOv7MyRgnsYx7PBJ8
k0YQ5iWnLXy3bCBSZNr7IHM9wQfWAbHXnSC0gk6yp9EO6LNMCJ/GedCz4efx+1lZ
Lrjap4DLKtm0R8IhFX8heigwghRrHC17Dtjn5dE6cQGz3sO+iGWPK6P0z9JQjLep
97MsMw3mgPGGtzIkw6AqI0MAnO3UGyECVT/q4QtX2PrqaXGQgEITZfmejzVHvMHo
1EUVu5nvKmm12NcOZBsncdeow/5t9Ub7d5ZMdqDpdqvZq0VtjQ6Ky9nReNxa7hie
+053KH5Izww9LPB7xsZ+uD1WCJoRg0n2dVQLqHz8S/h1GC+SGQ8xd+Rkkbgzq104
y8wK1uL2kM2Ary6YX0zDhcQ4k74NP4oQZRGYUVGoceTMH7jka0dvA4p4DwY5HVan
F+OUU0BdQ5bANP9NLsC81rhZewTqmtvAcc/nNjKWHGF3qBqMQkInUVPqIvv6m54H
naYx0mY39zRuCoXVemOR8OaU18xhNgldSS5IOXtiMAtOMgv8XE+hvx/U2HCC/DwX
qU4wOYTf7rSmhA/JcLguONECoEeLEdRp0xHzW/TMZhPkc89HRqTWWGv58cF6cvDW
S06gl82DFqcSy6LqMHs9YX1VZXWx5qWX+fP4dnY0dEEhEIpItM2/eVFcXkulit9t
6nBokgyFmKcKE9SsB5f0w+uUdDgCnZhgyxUyr4kwLXCQRgeRaEoTZnLUwnBBDnVJ
TQFLpYUx+DsKCqnEGdhqBOTR9cYfQ85ars8aiTB82AmY/fXC1zbZsnPH5lMEKQGU
qh438luWtUpjn23Iyc02tNDyj3t32dfvgBYaaYjSthrnIeUDSFXujvdkmrJMk10u
D/e9SQ1ISVMSB/NGZg8zUONVf/MjSnpLl37ACGrCHHMWVkAfk6VghW4FFWxCQz1b
j3oPQHOJ8AZWtoVHE+zEOiaycZpO9g+KSHaO6v8AMMjDv4MNix/qho3D1VjKWBu4
otapasm/5nZTUEyZRkCly0TzzA1BESfiBZ6YumG1VY2tWl72NRidoUxShYE+Mgui
nqvSFwxCzys4QqnUBtZJiXbPO4cx4NZtfJf2lJfKA7p2nmtIjeLisLSUMS1V0jVL
iIBFaGbnjuY822C0SbCJmMNrGhMgCm8Vxja8gX5Hj21b9vLsxJI7VHwI5KYntMLL
O2pZ1zS1JfM2Ugmr4P2vTihiST/y5mc/mWTKAOYjtB0GlLwwR2mSOJTLYluWTzBZ
xFt0m/Pi5FZ++46YaPEargrZoJH7NSkag9lXl5ct6EQwGtPddcj6/wLsGelHB2fr
WnYP9uryQTOVQnInUxUZmxPnTfHHrIs2k11kNRU5mFbX2Kdyhob5SxDzMhuL5nMk
U+04UVehP+e/aA970v6zdJtVXnY5mc9rrU54kJ4pmq8YC0Y0s17u2IBR+rMxVDj5
bv4XFeGu8DCSRbPn/gsIZq+NoahEQCiwJTkCmPbQl36Fi8ueXS3sFCS4j6dlXKRP
yDe01FyFtPl4js9SJ35fq06dsoyNXzwEHh2azNAdV9Y+w3xLmsXNtJx7r3/i7lQq
XxadEJTl4ULR+tHoDmaGN8jKs2n7KrZICLm2b2/VQxYtkIwCK1mz0fEzDUhC9p/i
bKclWgQXW6zgG6/BlBnQja1811ILA5YY3Djv/1g7eX/DZRCGLs7+c85jOPieDhrW
UU9stYXWpJ+mP1aBIOBpx9uf71WFAOTNFCScm5hxFoFy2VybHTEXs1BayIysReX0
TB005lgASKv2pyVMfToEMSuDKvFa6RGw4C8lS4LqTqrjZWvvYYm0iZ81/sWvqOBb
dVos+BduJ2QNdKMKr9xdv1d3MmryNGhMRq9OY1LQzWpP54t7EPbmCeZLdT3jlc3Z
R4kz4L+zBApjNz2qFA5Vgj4ZuSvNjgjZmTKUjgjvWGoeCpEYZibN8IWgLQj8D5on
1RNnipUSrzPdJG6dLeK8XDjrjAz4IfeLA43WCsgihhdwKMTQl7ummWIcAE+Lnvpz
Kdvk8hl5/zTXAlFY4Eu/a9DB/pRDknFWr428XNTYRChKE7GflAtRxBFpCZd7jrCO
TzHekDsFkTZeDVhTrQBETzDtprqwj9qsBCTe3jPbF3TiKIoCC4+DvMYhLitC+v/M
pCfWYw7Rzd/m9VhsB7061pVptRsbpzApHlLe0OvtMFybEG3B55Jna4ljXJFTQoD8
Pwav0HN6/HCVaBdt5zpeNLDG3txoAeTXkX6WECyYSrIc1KBgcmyiS6l9M4kkFCEp
oNXXgPC2rngkJNhYc2g8b28vZ9Lk3RRvbKVpWIOA1cb1pCV8IFAVo/RbHGi1F9+M
+BuPrhXE9a5p3a5Zb5gJCY+xcJyRlw5JwGgUI0S5d0fLDrQMHaXlTjFncnvbCVZl
q9VtG9Wivkm4S5JsfgktmTxVubvBROo7hmurlVOldwtN/KMEWQTzDcaybBwIsmEe
5MoW0xz/B/RzLLg0ulwYjxFbhZZSUjFsP4DzRD1HtCbawKWVRK+8dKkeqyUW/Bdl
TtgfPDwwt0d8MWMSrBIUaOdpN8oAuCpmoWF5VM90Ai2uGGFMUTvRPhrLU6PpNmsE
FOPdvH02Q7CTCC76idThm5bzdO2AJz5Ap6HahbiUpCOEUUJHyE/f+kTkZGzL+Aw9
xcU/KVknuloYp/Ar2ecGxE9tkgOvT2D7IlOd1w+vFZ5WVc3LnpWpgaVHj5TbJxVI
/W5B3RBd4os+3Sdgr8+ezsVyMfzWoPO0JRqwUYjQOPtdIFDeiP3Va+HTu4hJEcoC
YkHnsW5ZW7c3KBcFju6CqPbxQ8FA0x4SY6+hDhu+U2ZQ8TuxLR9ufO6AkkNt+1uy
ZCstH6Dwrlc+UQoqeancO4LwmbN4hfJh1BvqnwWBTcXTpepFZFEy5Yl1JC9jpMz1
wREe3vSSoCYhiWwl7BoOAW+aX2GAfUlJFB2uydDpIHHVTZeNTDV4DNjt7d4N9K1n
B5inmS2OmmmNtb0hICMrxBDamMDsS1gEON3kALIfnxNlVgU32JwvxDX4nqSUlfYO
siPr3xIAJ5yowbX0G5vzZEJ38NRQnfcj0Jb93mv8rzR0iNbAv34SzZWwhAAknKui
dayhhiZgIybMU0U0C9joCNZnD9SHEnBHWE2ZMjqgQLW7zhXDDrT/bE9JL7Mc3gch
0k0vfGDVG/aYE2YYXOT83A4Eokv3bZ+iXqpR0qgtGkD1Q2xnpl2Bb+DsaY94HDp3
8u72EXafT+2XJ4wFbo2BeRs94EAWGhBBy4eXvE+8HlR64IEykZsNQPHZxmQDp60F
Qj8yfafT6d2zqZ6ij0E5PLqqrAWppG1KCYYMNsMKwqnu9xzT9P51PyK59211+DBO
fxAbQ3mDUt+xpoxSpxIm5eNzWFxGrVsF8yJ+nmYn18bFZ5dXT1NXrdF/R4meENl4
hKHaTdjpYtS8ri1DUGe6qyO0px1X/LuMOWbMZbJffkcnCPbw43uk01qR2wsgRFXM
KTdzliffKGFiA83yOuZuDCz1rAqu50ro6qmvl21cjy0uXRqDedtm3LVBmK7aw+ya
faIX2cIhsnOaRDlOFT5Plv630jS1ibqOv0uDpZ6pzcZEauhHef5yRd2VGLxu5h5i
111KLpMITL8EZFS8bh8FUOx6d6DBP12i6MV5m6mBxMGsCusFAbEaONgiwtU2wcts
IH7tBwgmBDQ6yuQnifKQNaq6jZ+PlhVzQq/Mlbn/u92GX7PQz+h67vu3W1AkoCBK
F+qrA2MHY28rlk1Mr3Jjl/+FFb6UP7wETSr/YJEluWfIWCu0Od4prnVzxiAlDjhp
y/nARNtDawl/EWiuiQOsWt+3xOT1adpqTeZlLqBVOOMX8jEWV3PUpG0NicMWqj21
lrGolfrhXqbHGjX0hrdvCnsiKxBRGVB/k5xJR3EZ1vNiyZ/B2H6rIFeyFZ7O7lZO
cCOiUpjDFZZPwSUWf+s4mjWEGjJqg/vL1HvfKbF2HzI/+rCjBGu6kNWW3C3WtNlH
tx6l/mX+5KhXEWoC0zQQDOe7E6rkYV6tKXViRoArL+IElnBd9NEJrz6AqViI1vRE
dM5P3zJcjsEkgBZ9YAMu1XaFJy6Rzhu5R01Z+FEDli7YZMifCJdLJ5cUhCOMNUNN
w0BxXivuE2KeNRxIdRN05i0zOy1dPP3pnGIv0Jv619GoeV9KJObcybZ4a6jeG+2i
PTDYVofwLEP307jP+EW1nSVxL8mZKIODxNuGXSGkKK2+B/gJT11aJJohhQ2a/yl3
9CTyj2D0dwLrrzYsYAQzp2ajQIfJSdSQUxu0BK4ZpPASuUsXjYF1nHPkKLL3h+jY
48bIABpFN352iWUp69V++jNkL/6mFhVtxqzVvqy7t2Jy93r0cVhN9xumhjg5BOMu
O5ixjTL+PKbrl7S9qmO30gDcA5Ne0cPfUkgsCGKO1+jnRlXch1nX1hnWEwZMLa+F
/jBFkNmEAZfKedbzdYoCETjLGfh/A/ojWhkSDoll9C+zhjYYlZbwC5ayshNhh7fb
Jh0GvrrV56a7zjbBsQG31czbkgH4OCsCmeuRficQb4m7Q3nRBVTtbwLZIvxLCwkI
ggDjpllT+EdyvObPsAu8JWmtAMlHfL/4NAIkTNxf/VuzGiqvB9dBDpSzmqYAPv1J
YHvPwDfMz0XAm3J5afSChIBlgUWgELUXFoY28tva1IjUws8m+K0NV0bVd5uhtgDN
dKuSqfpsm+8ddag7NGACZ7WxUi3UclJ3Gji4iKB/91QDn0cYMZKyZiuuqeWM4Cdk
lLOT1wYiKUVjkNUaNfEUj7cDHV0t2jSQltd2uyERYZZIXwLZhgcIfy9X7ASNvKdS
v2ALborXhCPb6T5xB6FXptZTMLQTFvQjkN2IP1M+lnFfPjJE2BvWEyEsE3vDx0Z9
HEaMEWyDjYQojWYA4QlcdvH7mAsBMbKNqSJQgDMiSeUNBnLy2NDHZ4NW5trvjVyD
MASoRKWs9oCkGw3q0g9eKBZ8Wx/KF97aDoLq5eiUsEOa1wXV1dtQwqahpuOEU+ur
F+DT3gWglorkwtBXJPrcbYZ47lmsxRggwvsC0eta/9JZ7ttD/DSpxTZ7/gvhGXR9
bCr+UhYhKIJl32B+U82h3fT/CXCpMoWef9YXSGzE12YSbIYAFUtq8i7il1XZDzbX
7r/yX3aIr8U53qzKgFkGNoTOdQlIU9bsAdB3uWhQ4ZboKY/QEskgE0xJs664mAQg
OrPi0ky+k5+8RNQqSpU6AJiK9HpS3znsXDM7trIuwqrz6aDKI2Oa6uFIZnuIOeQw
SNozFDjhmGGb0limJXH+jr0YsmZPx3+OSlKv67ZK3ODufMCza+KnlBWPcm47S30l
Wr+vp9Sv4RHCyfNUIvBTqYeMYqcbtJ3idQ8BNJ2NoC7LEHIhN9tz3XlqRSS8cb2z
8J3xqEZ2sJ5pDgyfUFEf9ix+HTQ1uOb1e0lMc2kC0cwUBuzI4+w1VwiVPzjNYpVE
mz9lLKcZXzPZfHknYYX10HYlA++JpDwfJqXEDRrQdc+J/2CKP2pIdmft8/i+5Lch
vjayVdub0IVyOeoAv/z0bQP/gu7XZB2LejwadhH7Xfb/Jp8LyZu2nHrHKOYOMLMD
vipjm1NfHENv9iScNwZyykrNqUoVNIgkoqQ0wEzxK8pcld9eKRa/bo+2EZ9d+FBy
oJDYFbt24/0CAKAbmITjbPf1fIeYQNr+/MouZd5h4zqbsU5ADa0bdcfTvIBfVsPC
3qkj5JL96zReR6mxbyjyN7DGIMugo6pef1Esbke3vE30oYolgmicMAONDIabg4uK
2qLblT0fjHf/lOIhbNtEARtMIuxMeiqGtDq1xkhSe7J/Ahjb5EMOO3DJWcL6uRCU
B23TQO4ICK6+1xYqjlaPwv91+yFpqErv2P5zHnhPeJYcTch12q40TiISFNC2KiTM
2E2uEX23whoK2yr+9QW0HG1U3KCNAarpAKA3WBfmpo/0Q7R/lLsq7uRSmxriv0Ni
5EsnKSSMQh5s/piuulFqhxFV8MU7GeJxKHBzd35uVFDzBbV2htsRwKkb0KmCdYY1
pDiuxul5nshSnXVZi/94p1Kxy0UuaMjAf7S7chQfylBv2oXUvjYcNulcf8jXi+a3
zp6eShM6rJcOrFRCDeTCzTV7MtzDjXPcf1oupN5HoEHr3hbZ1ZakCM/5xI/Jlbd1
FeoDo+s+0HEvDmyjOoO0GF+thf0nnnzIAeUOoTzoI9jUzocxF61g2byntyOprPBz
3D/POfBhIRFUIyX5axCHXMI1o3hzPf5jeXQfvaQt3pPOc+H+lPNzdNhfKyKDOXoJ
zym5Av4QxaB54YgzkPQVHHLPor5GPt5G2LNANRdzm+nMiiFJBlYxecFt7gaXyDH4
RmL6VbO5bW3IKdd6J1QAzIDLVPxf970hx1btAUyzIqZoqNwXqE1721eENA8m7OVu
aVN4aUuUk6MvXSI6dTCB7c/tunDRozM2qadOZ/UfBbgalwvSpUjlq6YXVxSGCB2O
CmNxHAnq0vEB6jgw/SM+aAO8jn6yz/hG5KGk7rni9VHt29Qur/EUbeeea0zpRynM
ddk9vD9Hs+sfVvRbwVZHjZtcDExJ2m3KOklK1jTLfCyR3Q6jQdUUNxfjXGq++yJ+
1bpSXqZKRHwd81bivSCZ+yJElb0QSLiQ7d5siV3y/neJK7IBvyh7APsVwgaSH9bn
Umw+g05v8s0YMHoVKiUdcMYFp7uR8cBlpwtgHOfpZZGPmC3N260kmZ17fTPgxNvw
MiT7CUb/XWBuJMC2a9/0cziD3+7GLR2jBV0GjP1WgaUfmkeVzUqbcCkDygX6UMAY
w4GTDI7xg1gjqwdHdFBKUrJWj0ZsbutLhNKKMbL+wEGQPh/Vg9wnh7DkWMKG/zdk
kpvnNYzG0jx0IKubmZ2GQQCkaEdwsc5gYDV6kWOYApdCS8r6qc/szESCibh/hldv
uL6nqZqEzBO4TkoFF1N38CFkRKUnICkDbav/uXSHUtwfpNHzWFTjPm0+8a3w2vii
bS1eTwngAAGSWYByMXSDEO9xuKIQRBaMOnU9RGEj8ZFPabGAYjRvIxHZsXQrs+1X
2OY10Jzvhopd6kYjkTu/7ozp2UQtmJ5UCqG2IuuP7j3/ykYuApDQA2G1tCsgH3O+
G5wVT33dcTUL3ZQWp0UuQP2yfPtsgHOlXJ96y/oVIYteKngKEgLa7SJop3Bba4HS
LeuGR5sbuWI58h04LA0bISjNmMPaifFgryTuQ21gjk/PJY0WDx8+uxpWWhHhJkY7
3dRZnAZQuMc5BTjGUe1KG6xUVcYUykngMdJ3eEoMFWqJz7TYnmMjyqO2+DKVTY+2
Kmw7zn6o3hitEYhA7/MiU32X2cveMG34vTwsWJOBZM+UsZsEf7YqXHwl4jYKZeYg
32voz4WXyOVR9s/JFlLnf520rXi2CPLFdQwOCJkFMacKITZBBvJsUnUgIoS0iPRg
n9CrgU/CkQBEEUs9NDvV7Tl7dDU3QXggCiWYA7Kn3wY4tt58Pq8zYX5vB3YxFWdN
NMD0Gr9Sf8u7ZSGCXiSr/r0fMkCgGpGwpxytC8gAMsvh6kqknzeMmxDPk0NaHrgB
4aO0ngPZpqsIj6PcJfKzpVtN/G0ZE+LnTW4UTEPObMrFgnTXOygTdEWwmVHh217l
bLy+Vt5v+O8YynJr7W3fe3B6nrr+TxLbQE2b7DJ/q/Supjr5TxkOxtZSocDYaSbF
K9gSENN2z7GXXF0K0Y+PIkhBTsi87V2neRZn0EQHwZn8cGwzR+PlICpF9EpIRMSG
JEVwJbpkM9SqXI23tzaaf2MBmGALpE8SQiRZzBfIMhdGL1UtLAd8L4tLaC6ds53S
7H+9ioxk/B04FbWBBQQl74Z6LS4Sm/d5H4Cqf1zZQp/75InjS+gCvJkpYNuuMR1L
K6cjkACNxA6Vyki2ya89I1MHiVAD3va6ZTjrwvPxCPocoijz0yRusGUyNXl8VoZU
81ivf2zLzHQ22wA9WdqQLqwdrJhq1A1X39B6zvo62upr87aHLHaQ84PShiDqibp0
Q304SQD5Nwoxh7uXOTPQP9tRTR7qBrwCCeB/UuzkBRUaNfQ7qRhEj9nNSLiE7Gmn
dhRA4WrtXlt/XqJiLGsjWBXkW3w23xfr3dXMGTiFMKmQPVsLnRygkBvuj0zWYwTP
1q9jUMUZWWMmrJY+StXfdf0RoS2RdenDjDwN01MxYB9GJDPkBvz6WDF6hsyBlwdf
8/uYUz/Mni2mCtThaAVwg6ZIM4noDA1sNTFfvXdqV4VwNaG2ZGaK5l3rdHsz/9Mt
cJEVQKOYFiFQ8Oo8yrQ2xmmSaASZV5rtbJ+yf/qoMHrvStQvWL7K1Q4eBCja1MZs
0fNYMget5tvAZ1BCC+IFKf1nK8F0mNoOYI8XeJslFfu3p2jO5xEtoGCx+o0DnGjN
aBonyUTgbI4+nnTpIzPRg52floEUT0l8rhmTfftGB6LFas4nO4eiDePtZ1nKr2wb
J4mbgoLLOxpiBKLsM8tTh1D20kvemXbNZZRIdFiZqRsYnhdCeCKHm9JtnGqvfOCg
kVze0F9CqtuMo7D1JXEdFWHl26OLTpWqT1vD2EhS93zz90iJ1zP7bjpb7vNDsjWv
TI7ysrvzfXGMwuvERVnqNARhbQ+8/ngG67svLDBajUxSukzWV9CN7ah+CM/ldDP0
A9B7ZTUHn4cM+KrX6AkWHW0i0wW43GndNHSxh6rM0bu+aHxxvT4KXYx88b1B+f63
yqK/xftU6cyoxDmEi1Y7iCXv19IoKD2XT5M5tQS2u6EHZZb5rKSzBQS9BMJxfm50
8RCDrnxNViYkP3JdiDcqKbxoCSC5D7tZsmIXc+jmH1za1h2gcr352ALW97Nw9jID
Lk3yv1uPOH26P5Hg78wL+Kl3NBq51V6Fuv167K9aS3ca33Mf+G3IGuNuLsMlrmdr
w/nqziFRKGVaBbzGeUxNd0d9x4SCPre/Do6n20rdiAqxHHRHn52LcM7CTKFRQO1f
58tTPo1lEgQ/Ca4ooxAcHsGyTg9/XkFvsyOoJz/u9gV+D2FhLD7n4MzzrwYu8Ord
TrXWuKkCIKCnyZF2EVnGQnOUe66x0EgTa5QgmaIIs58hVPpDFbdBVW9nYcK92nP/
vyNWGyJzYnU+Sd2fp8/3wT3EysHR3ZI1sWYsIcrvw/5BZUwrICli7l52bmvfjDA9
3opGVbs5Ef/8evkPFaQDojnRw6WG4Sy1I3mOj/x7O5hYIdL1SEQ6Aw/DnpFVihRy
NvBgqUOfeL4YPebP7jNDT7R2/666QliWXYVpLaRXMGR+Kv2hsDhKooTr7jRB5LLZ
mv3eaWUFfk3/OZdv3mHEU67vEBV7Lt81YCyOtNvSiybXplnFNCo3ttnfjrWCslUa
OWl1WgY3/o17JiFyBBMij3ZNIfJr+YuiIkPY9dD9/F1Ay/UcL3av2xVrf3DfBajE
B5YtK6CV97mrl812rHLRqWW0cjTvAOB7/31yLBN7s+iNA3gXBvQjKvjaxXkBbRGY
4s1SRz7zkHgxFia047zBv8grhxm72IK+jR0Owr/4WaFpKZTT7eb8yaDbo5M0ta28
1jN9zx9oXYAJkkHKfj3NTCpmCDZgJHsZ8TQDTVCFWM4NjgCr0HeoLoxnJ7stgwSE
yRTnLaTyqzxYTIBNi2LQLy188Dw0FgqPXv6fyXQPj40M9Hf0iNA6uwnodjSqW5R+
HG6rvPFKerniIVexvmLDSuDixD16YMRi9+Wqa3gPCKLWxKiGZf+oENem/BzEmBAR
F5T7YDH362cjH8nIv0iQI9t/FQ6AKeHkVtCIoJq5uqRmKVzBM1FQ0IzWuQ5Up+Ny
+uOpGZDM1pCmJExf8Eps35bzquVsEPa/JEMVY285fZKz1ni2q2Y4o16vfsePuTyb
K72575zCRKU50I4BWz7YYkN41f5W0is6rDKA0e8847JB37eIsLqcx4IyJtz7Nq+r
1zuCCQIjl21hdKkIYVlMdQDx852RzuT4REgnhgfer7zF+cfL/3zG/OIBd4OjmHs0
5/xCL+DiGWlCj0UzhGCr8B8+q4ClUUEJ90YI1j5UYuzD2JvXtvJhyOu2+TiRn4pr
XmQ5+15+QK26WsfnaWN2aZagJ/VYV8YFRoEd+f4O9jzC3UsBqhstK52/zwDo4nLo
63eDTcCcrrA0ZX4VKgQwyaeluV06scdYsJphaUCuT6x7CiwjMCel+9K5irMYvNWs
+ZYQvtVzcAwluKKRJCah2tJLK5cUKZr8wi/sZCFXQM+0NHkw9gmgZZTnmKS52L1T
ZIJ1WI91mFVdeS/FdWnEgVpsYQDNFUsL7+4B7ET172H5yAwT43s4PofqjAVvdXZ+
Tj1dPgN4i5q3oREfVPRE6SEeie1wHQO7tpt1EaOvcEp8NzVcxKuSwfedO1+85SV0
/IPFOKNmdpC8YFGY4dfdxvWwFzUsCVGMXntT4vYAxOSLHfRk+35TvDOmqP8ttgu5
jxpPdmYcI6fvgvm21Bah57MCDOA0vjVwXLxmeNVldqSk/SRB7mr+EAgunKMye4B6
xHcxBcWi25vRkr+uQCJqOy+4SiRR5R4WYM420dSPPurGqH3/x8nx7+YPACaZzQQ9
Qes5LkAWzv6PN0PACJNFAsM4AttZlmSCj216V3nJAIUg7zEFvfD9YXqUn9Co4JU6
6ho52PPvIthDTJy3iGpDxI/ANSgCfTeyEBLn2nalaJgE1ky+DYMjf5rfPRILZpIR
pYNKwGDmEs6uQcTWBqrdNWrwkuf6HOp2JV2N796oPje/aIHh6ImwbxR+nzhOyU12
6V3fBITNZosQkOIhDCr1pknhXwjVqvSoxNOD3PsTYet4pjfkmHlWKI4aKbzBj1Cq
vdq528TixRf9RCPGcHOF4gGS0E5yFEdyTkNngKqNlcJW46dQ23R3c6Vjvbww1716
J06DYxWddMVy3MCrx3TTVGLD34rjJF7e2Kldc4UWdEwd1YQx+JQGZ6BJvTVPMAT0
uZxiC3fIxRG+bFBgeoe2fzmZY6b5nTlnfGoRQF1mGeLW+uNHHBWji7VqgrvQXRWp
b+BN4OqlTqNQGX9SSjX1BSZUVMK0rKYVH9QL/HjcvG+Yn/a079NzdQcItmRoebp1
0izKWJzhhv8eIq6YSMwXvvKYKJ4QRgvdpycae5ScoXCTpsFhpsx1o7omTjEpHIYU
WmGn1ZBG75yF+UvKPDiqQITeC0aQcgeIh1LR6//g1N7rtjdEohAVNk2LWu/5+3wj
AUDzd4sK58EdrrxNkeTlba1Eakd4H1xrUwaLozVvcDmtvHM3l7JmQu5jH8P0nbHV
T1F8BxoFI07tCOq+x3DaHlkaTO/ngXLHnYHnJmoSGfuREWCFd46dN+Oje8cQ/N3V
BIX8gAjuQrd2DIT7xP3c8B36aXW+hld5e5giTGKcl68i0IJLPi5xdCiF0nBXmR32
clMYqucKnG8FIJBXM2Tat+VJWxtBKprZ5AQlowT0CKzToacVXAqzg324kUTtfjRF
2AJRl5F/FCuRXJkibhE0R0yuqyPjPokteL6Yusof5GsE1EMopm7tvSbVxkq/opzu
9m3vZOB0R0G8tvmFc/uUSzQe+I0ovAHsqMFOMn7/2UUCrr1xnPOlMQQVzqjCBaub
p1M/7WwRoUBsQ3lTaaxpSVwuUY4btBf9f/5CHVOR5A8fIEZn4OA5UYRuji37GLSB
vwf7l8dMNmZXZHNK8G6SnmKx1SOGhf2Q2Rhd2O9H0jDgLvQLV09o5+fonr+iVZQf
faP/t2I0mzVBrnjgZXx9ySxroj6qB8OExQzrdGtSujDlnDffXOniHiwf6IRcRLZM
I2EJr22DNE5CEtm97eZf04MGpHWcXT2PVO4DMPtwx2S33bQ9c3OHmxmEcKeqmC78
m23D2i54c7OSyhhTuWTIPywjV5AXELbCJCxuHBzkJ2ZpJelOeHDHGwwf7IYW+xTi
bSbDZd3QqFQ+pC3f6A8p7K1zGCMDcstWdtAGwIevKtpIuQoGldxXCt8XNIEM2aWn
ZwGvtXG1D8J6UD1OrA/GqL5t6cvGjUiuZyT6AyBEj4NZMHYsQzbTc0guHFJ+Qrau
YRixX1+i7zxgl6zZxRisR3YhfE1aWXifFSLL3pbt55zrXzANYVLHjtBX442RuV4f
LeH2JFWCwrevKUNYgjY+fNsejkGqdFAm9jQanMrxEQiKd5ZopgHXle9mO2gS5Nup
eZVP/qK9JGg+95ELOcFpDpx8UWtJPuWBoUhbh4Dt6E6jGG55LqSQrDB3zNGP5o3z
svFrVtYdaiG/nOMiWekINgJzCO7u2YY5PTKXML9qw1ezVScx7eGSRkP6jqosxY3y
W/n8EKfNO0JWQZrTGw9uJLD6pQKu/eyF34xu251mbRosWtG9SnEw+Snlpy9m0hvQ
lC4Czl15z4X8tgkiO32FL186g5ynM5Oe/6bvIJAPbVOtjoo4Gh1g3YC3R8tK5ZAG
+QsDeb9G0QNL8pkBR/0ghC53gL9FC2dA5+6mwNS/0jdB7j80oKoL9yGwE3pR8WOC
3r6k7JKvDpoRfIpq/fXE+e4OUj7031y+2LqAljfVwazuAH5YdL0qFKZdCrzWiBB4
63YBr/hRM4BeC0gCYMBYBhwIqKLp3th1ljauC4+zfahYlEjJWqCYa/5BF+aiiXjV
YWY4yz3Ryww0PorJ5am6eroRNC/wekt0bLWWZpAJ8pOnkudnY+nZNo+2bUd6XCNq
R97P0lAOsupZLwxDINKW67kr0Tdrcz9rKCEYGCrx2xzNLvnaEtfCVfss39cwCwGO
kaDMEiVdOdgWGd82wn9kjYHwHRLjRnHPSA62kueUbNXCGWoWcMQfpHoQYCV1QMu7
Yvv6dScAFvuNFo0gKnnkGIDIOUwwZIBKXR8DKSCR/MMDCYVjhE3ScZIe2MOI0eMZ
j5PptGe5aqfrd/PhJtEiqVkryT2Y3P3nzKv+gjW+tw/HFD6YFpuNalA6wJ6Nb2iH
og+OcjrkyJvm1g+PU4Xa5XZ9hxERuTYU0SxmtSRwJEBeS405PwfuH7wtyY/Swo6y
LPPcRW3qxkl2YpAPgAIGp5x+iEtAJOfgRmwkzc0s/5bUFBbuFjeEOK6+JOXhbjlA
gUqak7JdLyxX+XziSq3VpCSzgx3DoCQCAxRT/JBAIu4GURT6cnyN8uoq9umQLkq0
OKc+aWlnFzsZ7N8Rl8F3RTze6208E/fbmB4y/nKAJb5WLMFnYeR3mnNVcKJcEEPl
TbNTF5wqMuMlN7F+LlXFnmhqCa9fCmYGNzDbgvKxEqzrnrkRMEKljSGZ1mSWSXkv
E/gizzMYT/Dx6ipXxj3jwJrtzW6M8nysgffhXLC4AxTsc4qWsop+nZRiFXR7PyR3
9HkjMqD/1DfRazBPfEqGfwZdYMLcvmJs69wHKhSaqjQzgYq95DbIxTwnaScZCo9b
h9fAAFmyyxnk/6vWUrz52IwMDZbHgIeapWou4/VSziulb3s7UGCrHjl4qv1UgXRh
1iE7xdyK/YX+90bTUKk5ds75gBuEtT+x5atxN7C/J/lvjO3pAQGRtQ6HXmf5IffQ
NGPG/UI8+Lyc8YL+sW42idde2ogLH/SZS8WW9FgdZ/JTObdh5Y/lrNkCHuUE6OKp
I/NM3aNcy7ujuXk/4HrHmR9EkEnGHeaZH/EWcCCO2JmXA6TpmH6ZDEjfDqUkQ/7h
2Q2gXPCmF67PnrRFcfV1dVfYi1LfcP+c/GCa6WR/vugZvaLX8lH11xd4mB3oijuf
hL72btERXTr4M1Lnwq3Nh9xg0KBKoVjJSdkk/vR/wy5195pzgN5PubAh0g62ygdI
dJ0w4c/jzA3BLorx7n3Ie+CiPVGf6lr3RKlRHUhZzuZhfi3u3wKumbdn1SpHZrtZ
kqyydQVpwiG/p7ZiwJKkCYSX/U3DvS5lQLMHSDsACzuJxmOg5syJIQwX+5m7uMcH
6oeTHJGOCO7cxuBk2GQrJVYsxSIs77764JlsgJz0uf5GDjkN8OucboEagC1S9WX+
/xnNTKY4lz9WQDe7Va143Je9QZER6J9dsWV5uSHHw8LF37MoWDJ+YhXN8sfHgZ1S
qQkP8xt9QCkOpbHJ8QcrijDZIbFZPmt5eynFnYEg58n1YUuE1IT+HUE1HjfomArl
nDN6CJ3txx4czwlkXHP5/jC3qtyTicBkRwzxwGBetpXfOsAcErrzXhvqX56IDm/9
SIZxgCNErq4zeibiY2ymDmfMOvVNKg8IOHfuEKoTTarhJ8f4bLdHBih9Qat1hqJr
UOehucTgZs5N8gfQOsw9ceNMfWK5uhM/dW3fbRfhR2VGvNJVlgulmwvgPgVTiUoe
JqNCTG2nbVwRM688+xXOVYVolx2nKftkg+1RAbJXZbB7yndELODUgEO9du7A35Gq
zX+d6kzD8LqUVs53pqMmqKJnr4NU1Lr3NdZU2cxWwlGAyKlECYyVxROJ6d1l/wb5
637VWTzxponUpneTuR+F/BMJzi3KouLiCrR2ho+HtvFebYoEgr3EqbRLXBURQQGP
W8+gkHs1qssr+TjOTLNNll/6dm10oRWVVD3OZsY+PKTvpXjswIQLLk1fMnozYeHc
qaav4C+Puuzyla+tIVy8RW+jgvliB6YwQZhwgj0bTyytTLgh0aSTZeuXkAlbWMkT
mbjx1OjWT8KhcGXOh1TC/p0Ycxw0MOBGiADJTEPL/6zXkZjp4BR9KItotmBHpwl/
LbaZNC9Eo6lKRZQQV1cpBdP7QSmEvz0/03O+wf7vOMyUcb+0MWOOzthFF8yoUiIq
3a6hMj28FcvFGNiit5EDHZo9vlZ+aufZwZD8DYieR2Fb6N/8gFjNEiQGHULNaYbg
TfwN16izgxxhOrxQgzzM7yXnuoSGidpDdB/s2tX3DV2R/DSyg1YAaMienSc97wfC
NuYXidZLsdqFVl2TJeJZcPRi9kHcAaS2zOtj0GCOciazXRVs5tkuNHdqIuGrVV75
NXL80UkBjBuXRZJmiT+tWYPazwgj+F/tg59ypEt/Q9+kOXQedHWsIoSnSfx41MLg
4tEpWIXzNxMGrjyXQ0WCzQXYMTE6lxYl5u1RZgOtYhpHbQxTTYbg9z7P/MCNA5WT
IpXUkiIkywajVPgEv3GM37duLFScbooj54IhNklkEly1RcDhFJRvwKZY3kisFSPO
XTKuUVTkZCb0f5tIjSEkfr2ZPshQZtC2PgITXLjtNltwUkfMA3igUy+SEFNBXfqJ
VYSPNQ9w+yJ+TeETZ5WCV+o1cTLTKBMPOWq5pqAx4rvvBx1rp8Nza3pDRY4/OcXy
2C5WSD6LhdlzA3Gt6x+bOSTvNUu9Jo7KgLtmMZwFtSmztYNBzh7GiEw6yW8o4dqy
sQO6xohrX6eqeI1pC44AjXUY01N/YcKhHYuebryHlWjKVv3LoYL9ZteckbJ2oE0n
+25jETY652k7HFpygLH0vz5//O7vPbwO0Ect6iS4QnrfC7dMBH2XAL4U6Ql6bkPU
Gk9dAEtGBkRU0/8rDCK265KJl5E6Vlns3+zMhQ5I//YYUIAMtN42C1htdx0VF7/z
ONpeRQzCmjTLNqiOo5azOmx39vYYql0Ky8shlkKK3DCNkUVym19T3Y0y/5yIXrDV
BSY7LpG1mwiLQi3vVHiLw330ByBPQ6ch1vilQDOwUMLgiE7qf82CE07jmz9gSzdc
G+Vu0J/IQ/CRIT/ApGLaBJn6y14d6WHwEyJgreCopQDkMBuL+1TfBIMDxtCQm7YP
0CcIa6+7vL3MMAeFGNtifsKvsQqdAa2HNJxvOtPxmwDJomwJtMNUaAmsHYBzQ7mF
aZzhycEVC0UaEyU8JJgs0w25EqIunxh5ullr9t9v7qNoGu0DLMMuTqvD910z46J1
ckkhi61ceyTM4QkvuU9I+8mKImTDkRyUF5RTH9JIwrjpgTcdfVtQdJzsEqKI56N8
3OmNQH2ZGHqn1XRPvzqIje0uTiMqRix0c552iIksr0SWw0irmLkJgiYZFmrzRJiM
qW6ogwRIsbG8AkLjwJ/eY5dpOBf3Q0SldWtg+2P1Y6D6aWhDY0oZMR9pcj6Kw4R5
FQA7G9X4QQyshE8IZcNjtiCM14xwW3pWJiZ8pkotjChE0rimHyTK9j4GU3wdTXr7
B37MDU7IPdDUJj94YxezQG6LpSXkS6lK6rLCGlG6kxl7rhK60Ry8SDhp0Mr7aHgk
mcnL6CO3QT5PtjH71zJqaIEKNjPb5rxhbe3Nj6uwUOBkzVNrTlnUAoabaXZQ3lhn
f01DauMVBo5QvHfuQh7HxmORgwyrkDqXkc9Igc429TLjdBAE7jdqgCoHRtsTJq8O
wKw3x34fIph9IykrNPYnLPciaULm2RPO/3X2fPbvi8mYlTEVWc78Fp/IkwZFf8r2
etweKqp+YAjILaAjRjL1xFd09+a1oTR2VenXLNLPAljsS7EptGmjbUHSA+WuleBb
rWnCDR1W2b8Qu+VmsUTf7MHJHDa+crn4lm8cQmvnLuvhvyBOEMvtQYnZJcbLfJke
F+pRQR3/hDgOEEyU2IHqx6DrSeEB9pwerjKYUOWasSfg81mhrFjr2tr1QNqMDcIG
0aY83v7Qi060Fq5re77CTE6T2MDPdDiX8AHUgl2dIQwphyUI+7gYlMkT3DOzTwA5
Wl2dKTds6/f09BrFucudg/bEV7JTuAtD1snM0i7DNZcccYwS+QUDvE6tONX/16cy
Xw5ekxKoH9dG9NgAoilSt9ZIBHwzy8eYSJazfUm24y+9FWkLMvkcq4rPzwZTPn53
C9xkcJhzLrFygz6/byTpZ14/NL9fB4crs1Vd42IBlGA8yVG69WHnhtrDxttVvUmc
pdt1aMrBpdcfOw2ycuOhpJVK4w1SENlRI/p8D+u4tJjh+ZkH1QMAr6mvGYw62a+T
LT7mX5/0vHKTZHz3GDZZAdArk0KhVyXD8oOnLcojCM61GaHOodyZ3CsTSpaDq/uQ
3/nXYMeeIk9epOe2Ja+zNsM7R4jMIOFv6AXd0WArmpOVO71A7WdwiazTv0fCNcno
7bNkbhwrxZQ0fC5tldv+ClnOFqgDDWYIzgfThX3Hv9jbfS2l+/Z1oF3szXWwZlEA
W8TbP0yQWGspM0qe0C33G7an3p84Q16xgVZh91RsBeu3VwbA7FcaLxyxf57Imk/m
kpI5+j2WTUWgd3QssZw8bA9rzK4ja6aMFe15omEk2PIANW/sj452mt23NHIb2ZmP
iCRKVVTKX4booNctW4bQfPmoan66kG4ucAOgoQUxabkY6dwrnpWntV332bmB7Krb
AOCGIpMbITFtkoyVxlFzy9e9uDaCt2F99M9rKralIFF+mRU4Jbh1oLWfKY+sobtl
VgK3UDoI0OqX2aLUU8DMrKV0v5bnLFFvLxw3eqW1xJnggyzv9ne7JB+b6DlG5KHG
U+Ta7hK4N7+gjXKTHMy1t/q8xjVYPDFv0gZ+YMmM+TWfOfiHiBgb0kAiXTaq+Q+g
oitxiWTpmvXeINISVphFwcd3TZ750T7KShdkoWIPTktCw3hc9VAh0zMqipWJ1Be8
JLHuHLxxEDdoJhx6eL9IgMwzmFlLO3bXCVCvonW5Bz52O2UKXRt7wFbKoojQA1BH
ipXERQREk4Bu18kAn5rKjEycOQm6MfZgulGbL9lZNZ4DZNlTpjZK6adSUJo4QO5Y
uf8VT/g7AY/2okO3ppdVMcktYRKo5GR1qjAMRn77jT1sgp0ZLLGxYVH63aXg0TgV
F2R71It451tNMOruoAPNvP3R5xizjGFNRwcDqQxWvIL8JbuVUHvFU+6LX9wJKvcH
YaDLUlfhcatQ2scTsEHApDtS9FS46X5Fn1tlTYdsaPaiV7co4tUJrWuRQNASSriZ
zQaRy5wZ9gmq41IlxoLlHvkCFDEi5cfwd/KG3T+eDOPB8lkI0Fpn9n6qem+kA7Q/
vFcGhy1pJubY2RHmJQrfB9Em9JyxOtU0TSv+d2uRnm76WSVb2wLFQuzYLpMnuTLF
bix+Med+Z5Aun5vY3kz3BkJIwdGYOzZkcSl+IUW6pmD/TGFTZYUDJTzX0jq51Ld5
3WNRdWqTsGM6IXx9ySgWF+wVWnBpfbN07ABAnm0Ve9T7zjvEhGmS6T9JdolahCdG
YghQnobR3e0tTgKtHSiFliGTP2NGtc7Ayg2uZTdQumd6aLGk8Z4cd2t9qhnYFCzm
/1960KVMgiFuCYKucxtH2FotHXkm4nQGy6SVllpJ6jUFJ+7ky87xHnTLUBzxn79/
fUBfdeWZGqZ761MwcRcKWGOmR2DjWyoy83UT7B/LbwEshFXPPgaJbk59x2GI506i
di6XJ94mRN75IbVE6/ooJAuqtaRsEyTu3I3qiv1r61rNPP7Oo55ITwAW7VO9aukH
xQM9d7Vxb2k9f8m1ttV4yVi3EkosVqHMM+meetVlWJJFIKt72T8vfP47QmDrgyxh
M99bBe/hV31+47pJpASYFViRUxoolgfD9GbWd0I2DVg2OklYRoicH2cCVgsIZy5T
HWgoYEENp35F0UdlxfIKVg7AVDfJ7z0NCxEKECnalX6s4QnW1gjoLtEis53hTb0G
awPILWIcGgYdEtHCq1mXPNHy9IYHBDF9PgBePxsZQHlh/jywxYlfiB3kRqxqMzur
iFfwwydSLAVQoFyLqNjWEoxNhdewVAaZ7Uthp4curNSPMfhv5npqempp4+XVQfsy
9JxAhPs8Eo6Qqipx4gn0MUYTDyrCax8772ilIV+ofGWcAhkD8TozX7DW7gTUJXE6
WB8lop1jhxAKSKiKEg2x21OGaxopNasP//iGb+jJljB+DLClWQtnGio82oua1pZ4
FNwX+zKi1liNduCzQZcC365F+boe1R0hGJPgl6zfHSgBr558+XbQu2tWSu8i9j84
fWNLGUpXmnAGjX26Cwx8GvIbqYZaOHKuB1D4f32Q5nVuQsW735elA1svO19ScdpM
GrjF//qtMi3wTZ3SyQAsUvBOwPHB1j4iyYK6TaKvsr5SXZb7iJtZzdfiKU9DxqKL
gEaZl0UoA2EQmbWhkDxv4bVIK9X2YdKMV5HXkexla6J2r3xbjRfGUw1ixrqEbz7c
p88iKGo40qene6ZsSVpONt18tNH0OurT0euaD7Z3ynO7IklfjZKChPMp27UUkqro
dz13B9skT21fBc4h48+tXlYo8Vmn1qxWD8BEh4i+VA3YoVOOjizMNM4wMHjgNhyZ
gaTe9zNMJpONotekSF1wR8IoxhyosWYZMcyO1iLLrjvHozbL4XLu/HDb02kqpVq6
ao3ES1RyPjW4LVSqtDwC8TCgcJL/rPYvhmQZ1hj2u0w+aiGLjHG7Vub5WPUFFIQo
UlOSjtcvPJEvf8ye06UmZzzhdW8nFdcYAlPUVLlZWSTNl31LGcvIqfw5Jd3o0gK3
NtSTfC8pnYb6yNndIYP6Oa3GbEgot0Frf/FrRG+x0qJOgOGoEF5VWP9+5gl6IPed
Ey2qmmXRUg6bn0CiUv6eAtXXtbHp1/Uv/Rp50cKQhde64R+p5u+qfHcd1NvVl07S
+Abu1jbVo1nlwzPQLMw48f2NdhqpNDgU+so/VuhBQcBYPzXE7NlbzObmKWano7sg
qJ2HSnXQ1D7hRM7Nbod6d6bnkDHxcSPqrZtQ4b7rqDvhESP9Ji0584pNaLCtASyi
ImopO6oy5sOsqJI8+WxViVS5ThbXQlBIoaDBmZwrHk2Ub5vcn9CtlDkKAWfV9KoV
177Ah5mI9ffPXi8ZpfcYtXQgboEqvTgWERUPwh7BF5R/JociyievtjpjwfZKbel3
fJD2zIBf1ojXPw2r46qRikTFO2UQ/tbkXtT4aIdf8ih33Vh2rtw6bMld15u1eVMd
ilgtAML4kpRvA4OFwmutUSGEU/O+0AQ7R6flFA/uQf41dNm4Lb9twNggKZpN2lu7
nidFf1tuMvdFMiPq4nhbulW0wB9XYyOsdxT3ROqPeS6ObEQzbJDlJHLtt1m2Vr9d
3pBHDNNDnA81+6eBg0Z+Wdq2kG12nBGz8jcyDhyFNdUozjuIiDB/0VS0R5HV+9ZF
8P7a6AQozZd5+JHb/SQAp9VZhaOUsjLQaDn0VfHLz0hQg5MEwhVcW9CItn+/e5CY
csHeG1/QW+k6PXFHXy4BjkFUnv/JInTHuJuayHKe4h2/b9akoW7k5P+4QE9qyiRe
tNxEGhT764iMVAHTyw1i2ZyimAJQHVNugM47oleHXcQ9De41LsP8Q+3oVnwyH3d1
ycMxb0H0QNrbSoQvsHwOSfntUbjs6oBOyan/2TblFXQEY2kFShBzRPjGDm2jW92Z
YhD5r+prCQafugbpAqm5aGYIRffQ0jq2QR5s+2lyIRxOihTDwzKQ0456MQtvGKVu
O/gmatU7/iIkSJDQd5xK5ixrLxe81dMN0Sno8xtyDuNsIqh2pwovXknKbPm2jwWd
iORNv2HFrVQtb85emP74KZvRD1WKZCOQsjoAU8h/jTnLrYxuwfTALizIeGndtyHW
ycpmp+XHIrEkpccS1I3YjTtfkCI7VUYnhOEsbyAxa/M7kiuui8O3f422g13iQnRs
SwwKb8nSbAp2bF8hstMVkpM+Bl10V5LZzBW6mAo12lo/0yhZazIASfjy66a/Ll6X
aO9jjdRQKODtCRRW0GONP8Ep5O1Vt3nsDjuDC3OzY80nD/IT3ilxR0EbcVKq+FZg
28ZPIsjFEAaZ3jkcqSfJoaQku5IY8pDCt5o9tZ1zpQqwRnySb8jcvWRGYWNKDhYt
N7/yk5zRrjZrix17CRrIvE2nj/1mIoY+ibl77qqr4XhVBGTiWD72J33DZSNWQrte
M1Y3OrjMRce8Ne/Wu035sERvz+qr/hIhBfy22oG33vbxCs+mBL3SMcbf+q0CPBZt
S6PZydA9VkjQiU6zae0hX/RUF0BLcdITw0jMDiTYlP3Uu4b3Op46gbc3QU260iDq
3r93YpMrn/yYzexDuVNICs2Ge5KVTCwObj3/gMBnTnamnZxdxpdhl8k/oLNgsjlb
dl0mnpNfEi3z9osvwEVYPXyHuThow9AlZDuUqgFWD64vCczwtenS/VbSPH15H8Pd
A9XXLAXO7FzUxmy5izX8xAqNYJd+mW3DNg00SrLgyLL0DPaiWiMYCEp1aS4AO0H6
I3Xn0ikcM1PoHAZyOYrdYN9B/LjU3CavFcEAWRegviBcTOf0PUCUxg29RsmzDdMA
zh3vEicPSjUhPvCVuxjBZ0NUmVwT3SF6K/MF8iNvmpybvhkjGB6ToxihgXsfApiK
gXySNUsZCk5CIXDFf8599T8TY+Ekw/HecL1/3JyZlJJetCDQFrNWfVvgvxXEcJAk
LQnvMszprDkAGv0VYLxjbymJwc0ZOb/6k7zMLhkI7oFthbrpmAkgBV9XFlcOuMRU
b2lx05RGefrKtoHuR/V6fD43qgUJRzdUyrJqXzOoqzHeB07gOZco4f6oTTuz5xFG
vscDZgCd6rYXGrRfL7Ix3CAbPbp/zPbhbqI6QogVZk1xziriBKOuGZJiPRq7NIEz
EPIub2zPEXrPAMFWfcL52DhbRNjQNfIIPcLdnUZMta2NrNC29XFPKytmGX1DNbHE
b9pdgUkFsTLGvMTdOChjHpTZ2yyrIgs6CbvZlCuvZbedKjBGMP0LD58TVSOWV5AL
B/wL2fQpJ9GCnApEu3GgTaotiEk9uV68U2UmT1NwVrNhftbvGhOvqvj3aPO7dsXW
FC0qWvT8ojOUlC3OuNR0AXBGNDLtPbshE1MJHPbcvESNjmJ6fIpU0F1LqCMojdmG
MmtKej7E6+DqVC3wcttGXPswdxOVzdkMlilRXtPatvfEVsTeRQR8kcdnnyW9iNz7
VoO4b4BHYu+UmlRZ1MIW11LzpIn4QA1mEe5cbTyIslknQwdRaLsuNqBpX+Q8+d4V
AbsFCNxgtdX0XXxWfkMXNM3el+avkamKhaPE7hbgb1IpOPu3FX52jSfklDIE+2kj
5cB+gE1z7vWt3jK9L3dahyfCgx/Ni7CpuHVd2ItNtiHW8iH+678tAESP2LA6/J9A
jzgvNj2keDmdJ8FLDsm9qz2N/NM8cijyRkIh/iavdPiocZQy7D39fd7g3Fo4sLye
fkf1OIUHkkjtXQUsBq48ECSuZ77lFc+JI42gbtRX9BbyQy3L7vtOhwvrAuCFDSaE
KXcail+aI+w3O1lUZj7Pe4Eqelt5n68+A92Zh7G8j+YhImoy9QrMIWmhgl3CtBze
4/QtXyNSOZU1aF1nQ6xjRdGv6axd3GnJOPrg6Tt5jZx+6c3IT8PJ++uSPMTMBvah
dy73TokwKdiw6KS25HSMna3Efe8XKQwPx6ICsWrV1vtdo2k5xHLwwU4Hig8IyXhh
zhyN6yrTI6+QJ55UdjcJ+1ovzHnpKGLw+XK6Ww5yKWX4PsUUdcKm2H7rzYN+2kvC
v4xRsjp1uk1wsn+JP9btKAm3CHLOwBE8XN1Ong7s+tHKD5KaavZMgGCSM8b+kANo
0y4/lQH/fJvj7oMLY3Slp1Ufku/uL0O27hj9r0kqOuq8x39GWESL6BkvxpKyMAoT
3UuWAyPkdT+rLpv/2Cl5iZPMbtB6HeoJPAsrkr6CISZlk21B7xRYQHoNj9IHV7cY
U/RbdO5Cy6CyI5+/V9k0Uil67Tno5wsE0vQiEJbhzE7KfdMqkkZpgV5e/BaTDeEk
Ox3mcyd8z3IWl/3AZ7Zz9zjujis6zHZnTwrnja7PiEEJDs8XLa8Y+cFQx7aGw7hs
1zLJVWFacYDTOZCD/2WOoicTX48ynBnOrq/6ASm0qnkQXMtndk5Oy8ls1kGtJdtd
xSCovYF1Tjmm5Dz1fAoMwVFGaL/RXxTV0TUijGdN8nIYeesw/w1r7lH21J+zl+jU
rQR1ytdemTqSp3BssGKj0V0rH5uxmoj8TsQ8y566bfVrkTZlCo3R5lzSMKjF7ACh
VmWH9zyRCvED0scFZx8U/M4/gY3EcWARmjWiWGxh4F4neT+Z5axmSC7gG80YrgTz
wLdskC9cDm8urL8SiSyBmh8u49WnKrQnlH+DYzp6vxIDVQpfoU8GnZ4YIE1B36Jb
EssQPtLEj09FLHLWwfQ9WSr5d811XCKK9MdJ9juDsaH3NMfs0ATCtES4VTjPdAfF
HlyH69JY9XPOs/Nxdirc1GJgDhEQ0iJtUSfp30ZkwP/0AjUvReLIP8YI/7LeGukh
CHYEk5tRuZtyKYh3h89sHR85PT204F7Nx9RGztT+QDGVNhSlWXpjpBbphQhEBrJ9
FKDibUEhS5f4MHSRJ52aiYVsHUCfLQvS73kkBq09imBQ4O59Qbe6la3Hyt9Tzy/w
hlSdAgCFcv9EiF23i7j4YC/tnkrdiJdrImxAvct8L7wj+C/zcjBJty4C21gQTS75
/HYDNWWPe6jH+5vd5l3GMZ7SM/6sSWOBc5HTkrLcfNp/keCRx8gbqrGlxQYrO09x
8D4LRukSnuhVLgu8+kvMPDi0eXD2+m7E7UNImDnftgrT4Y6Mi+PM8LM/kgMUA1G8
2DmDyo77OA66RAX6RmEXHc/VPw1AKTSv0gKTnzEOm/vrgvQcNrwv/FAADF92nSlr
Wc2zOt59ma8rHNaINy/WP7CUlSbZrG/rG2boRKWAQE/6JMy8XZTeDAroUha/MoPV
YfXZDnXijoe0SHA4SR0osgkkdFXXmo0hapZuDBMzKYdmYOsRUUyMHkxntAnuCKos
H0tMyj97/Lctgzctdf5kXQexgPG5w43HVLAMuxj3vddCtGHS+77lIkf6sR23o09s
WimZMnP0/1tFgwIfYZhaZZIhJ8GjKYxSwEJ4qQKzK66Kdp8rp89759wbt7mHbNX0
pkp/KFV5PY8yzXJmJgDMuuG92hbgykg56uFSba1D45o2faa7t1o1HDhnuzhov+RP
w3aOzVDFREDfMoOD+DYK0mgB1WKvzr+uxTKHLhtUgZiG9vHZGQ5jq88+O8yz/YVt
E56dsWlgSa4JugAAjGetwZFCI2s9lKAUKQInFujZxtNziVsJzXjUnI9k/a7OGieO
EXzi+Gv1RVosOPxGPrjbwEHuU8FD6cKQDfZG6Nrr7XTynzw1GTNtZt/qRuIhPWrY
+hQWmWksZ8eB3KZR3DPGSiFRvuwOqh+PZ2q81ACCd8K6kF2xAQcYxtq4bjXxGjUg
+XLBDMjW0IWdaDmsPTZntH9nXPpMswy2bobqEFh54S6GU03UqwRUw1/liwbWGtVq
TZL5u0FPgMjJM2zeIucpnFS/mGLB5DpPzwDLopxL9UFCMB9cYUVEVjoezr8lKDad
HC5MM/feWUsTDxVurMXFYEWVn7DaMwmMR5pOhOT3tWl36K6c8nXiBOMw7twa1FO3
N7BB5IYRMTHDesye8nZgjz9D0cukVvnNDTJPCB4fT9rmw0feD2VWACyF5ZJL6SNm
GiTvK9TNP01Lf2jHCgUi1tmOfUfysi8C/WKiZSoRkeRbhNwIXjmPq6DTzB+ZZFhi
6gSxzBoLaAV5dEebLaqRcbF5BBB5qrNZ7A0EHPPI10wZrRDm8zpgLDeXpReFRKL/
m1/yfv1o/qCho/zt7K+ddoMTDGxif6GnVDrjaP5kJ60w8fxwJk9XPO6T7j/mVjLq
WvlMPHvMczIRqUOZEa9i7X1u0H6OXB3CEjF10ZJ6XC38MkoqDS4GznPjwXXG+I9I
NyLkfkGrG1EdYiXGnTWYjEtpxAeueAI0Gslc0Iuqhha871CcHwQzxNp/nabBDTBm
USbB99cji/fAs05D7UCsWb3fKJzlXfyoJxCyly0jrTqU/zcHkkTf/sPi4FrAs0h8
RF52gWcZ7CxGucNYhsOpjTMz5bV6/4kBk7EPDCBE5qWzX7cf1iQP/RxZAM7b2fca
BC1Uk/pASrU+h1d73dTEstnrKOZmjeu8PCyQmcEnO0e06nrz1hNTc0ae7/MgiBtX
RQoNztMxMWClS3QcGlLh5gIymvG/rHCn6MTUzOUV7B6aZchx/vqxiEBo1RuO0hDe
xEi4pSoKkVEuS986cURSPujfgA02gxjbJEeGO4Bajao0ist2LvIzbr6elv6e/iYr
IaLTy3Ipl5d+LJEnqNG4OkyrqR9OD8PY0Dv/ouKPM6phlCo0IUOhEBt9+UNzxLl/
WE8dYQsc3oQPQZjw6C/I8QK5VYDqG1DobaZAzMmu+THLwI3K0+TPrHh85Z989TCw
ryHJzs5DaFeNl8iH3vwJEpoFBJm8gdBS9zT4t1n3lBShtKDE8lWCfLglErCmr+n/
cMqPLx5EqGnpJjepTS9NSJ3+d9ARH/TqE8UJZ4B4r7eJnVWuLDSG+mI8tIEBUI8Q
SitZSqvn2ragAPFRxJTN3oJxPMTxrgO25+uh/zN02Nq9LzHNZwUHh6EeDk0EhFPq
HKT/VcIBd1/y+MtUxqNzUG5lkLlNT2b1ZjrJ/Doun3GLP45epgXRAvGe/QQ1tRSt
y/kpfUvzabOlDf6hHB0hPXGO+dfDycX35BSZEd1IIG+R0yaFdYpuiymrJNZb+MW9
r6BajoCFRlUEe+8Utu4uoEyxMylxJmuJrpfml/7jpKvUOTMgvSvHeS0DKppHhqcl
hs9/KjiNVjbd1OXdY4Ugh9fM4waWPpdiXnSQvkkJkLOIWMSOYgRK8qgEIKRTy9XK
Rn1cSzEkX89ojUJXoygUPT25ohNamaK1DiLH/YG5E1ijTIRUm2QH+PI6fgMAfroK
YMu8qYt6pnesJ1oQ03tW/CQQHT8nBEVu0j+meyAcM78FkkVXkodjv2rmeY+y0cBX
G91znJchrocM+nKgjnC/Tm/rRN3immR0VsWhjUBUN7oMy2jjNrTrgXK78JY9mlwl
e4BiLNos4tp6DraG3S8rBY0esjWwXbfcUNZ2ZA9Hr1v4tnNdDL1CthO86vNaLEnF
Wqls0pst9WcXNSbLx4mPT9A9lC7ukbQotyYiDo+ZWhFj/FtI4BjvJbZQY/gQu1Fb
1k83tyY/iBYc0O2dodHiBFjTltUlyihPQmmxDawY00DNuvW9YIDPqqCY+0FBF+0N
jK8hqChayF9ePqh4V4VVNwEPaigFn90UCIbwT4r2iIpVzOar9mff3kuZFfIQBKnz
n6lAz8Ado94kHhIcXZl8CZywyDBeCSiNYkbsefhqL589vKRCnX1uW1VbsKEKnLzI
POny4PmLKKm9CvDpFtCpxm52Lrm5moMRL9lS8YaKf4Y/iInQH7tdP14fuoWbpAJt
5sfbKvV7/xvsOHfqkFot4oI/s23sVpNPCXrwoLu3seDV8oCV8LnH9CUW66L694Dc
B8AOxqMd0y2JWh6mzH277zMbEZnLqhkp+nShRmDpvgiB07GdJi3jBRkh3a2rIkBe
xuaeh0hbTPQlTleKYWQEVa+ZaJNt/4poJo/7YX8JPvQAjSpjeKoDs4FJxGVsjhMa
ef4Rzl0lITX1ic/7ybICo5LnPVsUl4TbQLdyBHJCNL00jgqD9NeG7JLZ+IvmTX+u
akKZc3UMwqJC6PX/OwFPmOzqbnCwdp/Eu6/XC9R7Cz414w4JdHyfYhZsORMKdPzK
ib9nzEYoUde1hLhAlXM/26KIdOhpE8MqvDL8mFZaawXcofkrg5XoSJ6Mkzm1+Dvy
UdU7g/N/DQzOFk2PHE54CrvGbsFzqrrq8mfZTvHGqr0rCN4lqBqvHyfaryy9odJx
N2k9hRNowrDCmtduWwy8jjDFgOmWge+i50GL4qXeqBxX8cmQRLIccdAKg4UuSNWw
wB2+y/yrVXPu8djgoiaGSgTkN9qWJPnWi0hfxvDJTS274lFxryaSBkvAocvWnVJZ
r3akB3jOY0eM7qq8Y0YiI3cbCUIoYywer3D+kXJkV2ZK+6RvKEivaXI++mXJXn0R
4Xp3UNVe6dZaF3ynRNggFCBGmaPCJ4cS0X1rQk3R8g9i02RKJiaN0wgB9md4ZhYh
UaqTkyEAvlSk4MfVKm4oO5RwMvShinAED5SdZrebR6h+zNrxPaWEMP9TRFeOyAUp
8oS1jaWIvyiIxUWtXf5tuoYnDXsxOD1P9b4sqXt4BUDQVnwU4Eoc7sC8aM30Wyyt
3QBtx0+gNzosjdJYnn4Sedxhto0zCOeNdcc1t313nlfNreCb1V5A8KIYMhUtyvNN
XOcwikzgHNRQQjWLjO39EPz76GsojAc/0bLn8KqXbE7k0nXj1jEYZkToRdNeso+I
HfIBlsA6/ehJjf6VXx4iKpLQzBEX3sDE6y6aQEvuI51aGKebkZ+oH+w6KsSGHKsO
Bhq3kG4SpcTvRiYFjT0rBUZKF0FXKnmLjcOE8r+abRHo2JJooIqLxvce4SUk8MpU
IYa0Xgf085zy29wywk8MngZ6GNFJw8ADYoJB6IAeg7hWu4RCYCUJQiwHRtRKuvMV
MEB3/QBwdC4yam9wvhWWiy1orlVkE2Q6z0K+N3gnDAR0Pqx4BUHdQvvjtxt81oU5
6KnSvT2bI47TFIaHMu28L6Kk0vA7zPg4rbm8syIxE9ol/bnHwxfDZzWYsE9xYa0G
2VmxqPEer9FlNVxR2MwPXxTtJnhGfCKxXuUjVdhqZMhViXVs+c0Txj7jMVHfnczw
DdT6651J+eoPpHnujQLF00ZIlk6AMriOFBEAPoUKNRxNliY1htlwmV/vfVul+d7w
Vj5OdcbFesOu5aGP3BQEQJWLaMvAwUXSv1hXi1aLGNLrwANdTV/aUp38fZHxa+kF
IeebPGVcv2IdglwgDDgf5+yjwwps7kJHf5cAWHNJAe/cSnOTdYA3gVH3FIO8xIDq
iQ41MubZz/a0pL/9LxgCSBb8WAje/vINgbsnM5w7kSZ/asmgoyA86yl+hGKm83M6
VhBGcPOMoV/Xe32Wj7xIKJW8IyZsr/TjTT33aMCY96s1xP2BQNi4p0a+5eW3zPDZ
POSBosTU0nJt20fyLXpP+jqK1AzCcuhktGgi0DFBKb8cSAD8AmzI5IBaLP3sh5G4
7FlmRfKYGwOXHukSWPlLVfOjcxuSrOsPjAStymVLNRUAVHJIYintyIQshn17VJSw
7t4QdrUBh88YuS/l0KTSsRuOb8OY18wzvSfltwL5mxV+2vfNO+4v6Lka3YXbrjF5
SMPdAxY8kUjcdcjZXi5j4pN9txdXfs7A7+KNDGQch8sn8r4lzcZ1Kn2t+4Uw6zDD
GOPEINf61sTkhKbBfUPKS/Jlqi6t7T6qDv9+5QatLs7hRyHukxyCOnzJORkluE7i
QJR7kA+D4OG8Wg+2Cq6a6420hRWHRqeFaoyBmVrQ+qTWUHvqwb4nz60A4q352Wul
iTv72M6lyxnXfon+4WORpaiFjbxoeft2Sn7TAhO9mZ2VAizHZT3MpDjp/9SzuhpW
TwPiflpH2s8JXk1WLmZbAx9KlXnhGxQ884hMBrQOSFDqS3g4/W7gt6jTVgFPk08N
GttLQnqcWHovwRLLBMp3EODdbBbQ4WJlvfNHEisAbZb+rdSmMs/HgKU18xZUtStx
lKVAPcDKLx9Th0mrLEpztuaj3yTNOA9CKGjPmB4aBGJueySa2IoQDjJJnzd/4cTv
E8fxNmiPexqi/FomHobmgy9SnWohbq0q8KgMf+Vj2DreS+fdgkrVN0ChBMMEuRL3
CeBc5mICFd+St6IYDD+agy/ST5b1QYPd6+cye/qotuArdI4/Zi6PSGPdLqwzrBf7
YkliocddpYvRnKEMe3SnsocfiJtCCyjbnbiobEjFU/1qtvzDGlQynMnC/hnFjKqo
yJHNtmc1BVXN4tQdQcRmmLrdXj7rCKbjFpPYgw65jiiWU9ed+3aE+zPpn3qL0AY9
bQd7nWymnBdxnCZkPFj0LvCWhtZ1NIhsnOEWN9+ZO7WTYzjdlszgYBtSbAmNUhj6
fbRIPWARQ9yYnXmH4UFoMHqCNpNB/7D8X0qFXuqG+5bXo2ryqWG9Z7LC5wCFGnc1
j0Stuv8EQwpWQDrbFOuYkApyL1cn5eNwDI20gjhQGIlL06AT9mK4da7TIw/0WSKo
AzXYqPS32YwOi0o36pdKUOzk8ZQiTWYNdl2KUoE44hTzDL+HryU3V8CNQns4UZfq
/GqXm7u7Be8RX0ilLyuLUBUaLWvRO+vArClV4UX1QnCbLo9pkHHRhPyfTFlKkF5F
DHL6EkJg9xQhjNqnq+zxcS+sLt+dHB1MQOohdvKxUsMUAFWT4q3BGPSCLW9YnzWv
f/cKs+GLpVJLJB6wNwWHPZdejiIZJwz+BfbPmhVh5cRw5zyF1gWZ2/OrdcBSqBMK
Flnwzh0o+UkYULi4dMB93Kj5syvpQgmhdY4SzMhxX5c2/7dvjrzPKQYiMzIR3JQt
AZUrI/uUTH/IdnJGLkVC2Udky4mUgMOyzugPJ6BtkWBD+x7YcOLVa+a3USwmrkbY
R2KvIndk/IMwHpDa9LlvnzbSgGYJ122+J3NDFg+gxvJDPQqfAn6QYyuWLfbWjgGp
YuIv/2LcjIwGyQketl8IAa0y7WD87c8ZnBPfTma2xxVLEY0NOMOu9+lGo661Tu2v
XPPe6/MgBBBgEBE9WXaVmjTb6NATMMHeVd1HcID262qq7j8JVVuVunlonxRi7nvh
WGUxWbeqqiRV5s8Z7Q6RCgIWLzwhMSphW2+PfIrFxWKBv11gm5JwRngjgX2edL6W
0CUQqucT9pOQpFPoIwgrxroZOF/+j/XLAzjPp/MJWdcQGl+llBg+E3vnrlpGWZbJ
P753bz0hk7PEh0O3yLjKRa5Rnn8QzTv27PpIAhree+k4NVkqwjgS9xHQcZqfA2+H
U3AtKsISHKmU0j1Tc2XAF9oPv3n/iMp1GzaDWbDjHyDIAQ4NGcgAtuMtx/Kwlyio
mD0UzOEPDTEi2FJIAwBIefqIzOZ3nG6i8PJhM3c9lVDlTe1On1PQW6rMU/Gg0Lx4
Yey+SRl4zL5uv8XyISz2k7VaKe7tJvZzbuEzncfc/cJpDJFq0XkcgJ66289YfTBN
KmHcD+0tOK/8S6fbmLrreZDhO2q2qYCcktTfWq2hiKrlb/jxLtR6SYtg6o+pgEcu
SaNradBFNzjImYejmQppPPd7hk5fD4BVQJRmuZrTUp3/E5JESRUm9CyKcpwhxRM3
GcvDOeEnH4ZcNYmJW2YYMCjjWfBUpEH3Fb5dgofvhuWvxzCwanAhG6FvPjePCCSe
ivTNdmqt6wdOukLmFkIDimpSckOJdWpLGA6RoyZnJx8T6SlLFL8xgndPWnM9kqM6
ae0nMa+rgpgpDDB/CvclijKWANGer32WKeaZU9UoPHy55Se2UghlQyJJTK7WqCzk
6mcatrrWYx9oYl70wHo1ZNLmHgmYo6WZtNJfnjqMD8czZIJhJVunbsyKyx7RE4F0
hnA24b6u6tpHbSMBt03Xs315vXP68EBFBsB55VhPwo2DVVu9VNjo4pOYk2MVFXv6
GFAlQzatAxD8HhRuvOnPq4bCe8WrDPtm/hWMMlhRH7Zk6x3R0CGxa3h5/KidgpT1
9gowL6ru2As3vdw2V0uswbhBIIZqCuP8Kc7vRzSH6bekwcLU7uCZkg496pQS7Mpu
tv8BIMRSpLtuHwoncttNzvkYJ/WaQ6Ixcpx7wKqsIXpEFYQDJMizXClutw0VkS6v
Sfql9j9t6tBCCJGNLdehT6LIaqEmLWvK7hXVOORlIjgcmcdGvdMBwDLaH4942VOQ
DLoRhnPzBZE1NOP9E2OC8OpCRPil1sbTyHpUejhfziTlk6IhX56wMJ9gVnX4Pow4
XX1H+A+A6ZQh+kv3zrf7TlXfiKZX3m3DG9blQb23GYvJ49oAlfPdKs51FESJ+FcK
NRvSiD1JsjRQsAwvOXgz/Cgq1t9xQJpysjGiJxLGGfClamr9Kb7ezQcNsiqiuQsL
1nHyJHYeYmRpY2cVlddU9PmdEghhvX5RxEtYXldObjEh9AnOMlpi+VIfjboHu0Uu
jOZGyBAv85VDRptQIdUkEhg1cy/dM8ZsALRJvwYM2x8pnJ9/n2SkdXchFGtmaTPx
Bk9H8QFB2mwV4wJXAMM32XwL7gVRVE0vA7+WLKiok8nvviVSYZFrKHwn58TSHHM0
QL7yxPXhaKUx65zFOL+MgOJ9jaU0jjmddBvdHlIuK9/Ys9fCFvxgxT63W+qDr3Yi
yRWxPttE1CBOPAxEUEu4MJLBgng8u/6oOzRCyK8KdNdaNqIzQTdnlO70j5Q0y7ll
UcDk76Pe6gEw8N1DLO12gjRTdfNHh5dbnp+jUFX3b0Zhfu1U9K9bmAu4oXrquuRQ
ss5tBhn6yJMdOCOwYlcoVrzSLWDmOzIe/+7n5yuLE/ou3pDdMgJiMfIlraKQ/HmJ
wqafIhvvj0HZCA3/yRkSK1OINOsf3K9tB487jW/uLXhdaucviWuC2nEgQqHEImZo
OLWhV1IwNf1+6zIndcEAhs1+Xi9TpVK448qMlNsxPqsGFay9SQrX1sJ24BuNJTXv
ruWfwFKSGkJha1xt6lBlz5iOwOwobEXJuLmtPfq6m2BP49YDVLA0mTpN804vsuHu
/jCqEiaw1DBCaKz90vYms4RFzikU4mw4oT5lokUGvGlXgNu36y03m+PUOV2s6lk3
p1YxhJpnA9aXF880RRCWQXNfIoM6B5xmrbhiaK+MCyXXXYcyjj+zOqhKvpQApK8A
MoTuDJQDnz6CgUsI3DNFUL8ya/DEE8l5jyMSn0kS+cHRsZcW5a3moTiZzghxsKGt
/f4BJ/0LGq6KntlIAu7PGTXeXqwPP4/oG5GA8ZqypdQVyA3nsdXdMkV/rWxOaoJQ
QQzlagb0pgBddNNOrWUmVjUXm6CSOzJpeOFXqedjz5gWcIjsBSxGjKMK5J+/IrfO
+Yq4c5j36rgR5Pi9r6hN/xu3WzTGC7suFfKH4z/BUZNhL4jW8cGIYwzxeqjyNmIK
ykaseyDcjLzsgr3Bd4WEKuKmR42IS2996gEZOPqzqBGe0Q/RzSqTLA5edLu1VeCf
fYbuoQSHFyxRMa1T8qQdNlwyUyL7SWknf7605nWuzh/ut29HAmBZhLC81ud8jU+5
HzhsDbU72W5lAvmqzRSbKpU3ImTxihWxF4IcJ8LVYzwc+RXbVDVIzro20gaT4HRt
R/izhjPdVspsno+8ZrZ2IEYD458yj8VOgf+49iBw/09LeyndFeo81gbDCcsnWEUY
qzSY4D3Y5qox0sTJw6rn7QLvXE0zKnynffzIHFRbQGasmMXldbu+dUSqY+5H/3Qm
7eDtKNWNt16ArBD4fFzOERi2gIbt3O3dzm+K9BAEKc815TgL3gY1ZFPiyV5wKoq3
MxPjQrST7YTC9IRoRtvVYCNVhsft9RapSgOIoV63IqMb+UueIR/+HjpnIgZIr3JV
KgLr0OpUqd9XiXuah6qO0zzlDkFntXFDRbK6mc+FawLqib8m6A5rlZpD9XMB9Tur
QQTdQ1y7kTvT7H9zIifm3dizN3c7ssVPcUH39MzUuTb6bTJashfM6jfFNK01kTrS
Agqr0B2au+K8wb23Ugxe4WKTtLuv1Liq5LhfNUe/Fuh4/hbLjjvTnTfXTkb84LxI
UOmWPzoCZoquzqsEvNUJu2HCA/dmTQK9vd/aJuwpfk1Q2NCLZqvSxjxYLiidBXPe
xLWTErjj+CBXzP/Kse0R+/21JGEy/DCy/BCMqMP4Vm/o8HIN3YPgWKAQFRTC2AM/
IDwWaqi7wOy7OLXHX9+DV2CjQXkMaXYFHbFz/7nQjRI0/E7ZxxuysRSScjf/8emW
7i0ls1BJc9s+PBg/+t4pWmAZoUinUBwukSlaUzUL4o2da4y5xzVnaPhLeoqSgrEb
IZK2C5wwu2Q7MQoAT2PRvmXRHCxEGPxmzePCWRPCI6EwA+t+QfmvWKEEGgKvFp6T
2SoTr00dIx5FqZ9+q8mUDV2kdQFq3fhYrQBzhGShlr70j7D6PbF6DWU7gCuNmwlx
5OCcio43h+2snaVzFGwmk81fkRMzI3w/n/sDhUIpCkZ6K6FmIgGPUUc7LarMEhBY
7BhsveT1/0zPfWBEcysZzdvsln/1QvZxj3B+UzhA1fkDZoybCfwvz1X6MtEeVPTS
AORH2rFyQvTTXe3sGw5h5xS64l12zkQ1cOb9LDj6yEMdj3CUmSCOINaMD2KsdbQs
iiBzqt02ldduhgttGdOjRxotuiHJ8l5Q/xaoEG81FgMyXKtnXRKaFNrt0Q74IFeh
9rXAwwXyNS4IR68Zx3k0K3dU2zD0QmesQCx3sPexh44HpnlR6rqc/SKOefjyZIdy
IFQKXe+piRhAZ6lE25rUJtDgdcjTlKPSB6zTJHnWMzW1+uSDDBzP1XCyUrErFruQ
s1DaDvQtLCor3lpUtGF0nz9ACP/6FGaJ46JJ2Br0O88id8yp0GVgBCNzuLZYLjJt
hpu7ujaNd/bcYXGTHszLNwKzUrL4V+pn/1B8jCdjlI48wjbXrWbOXhMwfXfpvDAD
mxPx40K1bJsm3YYB4JT2BOYPlIlmSR8RblOFX+R4fJHNpBxI1Pbz3YsMvO1RVo/Q
6Xz6oGnY6taq/5ldJhaDUrAviXz0ghefJywtKsyligjNJ5EAcR899Y84/w+ra0i/
fZBaHyCqGGwvpSjhT9UVHWc8a0ryX4GT4s8bD1ei+NdIuKFY3rufMugPhXXQka3Y
L6LGMfItmQ6drQcG23vQBguXwslBzsPTj68ZqqB3JHZMj+NTi79wPt2T9XDCn+5/
q9G2uSQxXk3IJwt1pvQb8RtcU55mD8fLojDUpf8Abi5Z+x3SBROmrWj35LfrWiCd
PwURqUvZrbmI4AOo/gu0PkaegCN2dh6LfPV4tgvn2HNk+bNQxKIOtj5yas4qbRvX
m+z1hXDJ8SNNQowD4+6eNbeTPRI7SXGq5z+k5Tmqq/VkTJR7iWOOsN1hsa+Z7dW4
so1YbE1uR/sYOr8RYmRrGYU/H9DMEsTUk/PLlGCHCtoj8QNssEgCnkhqggywgFC0
19jkMSnmS7ngXJLqlERz/pd+7pciDt56j2oF3QHTSqwp3IW9vy1l+/85EQIlkw/2
hSDBR5Z0iOloiqQyLgmJhzR+zUpN0EsY9A9w0fCWHslaSUPyZnYAKx2dFdiLLfQX
5s5cAjrxyJotFsmAmQgFeNFUVrUxNxVbKZHeoFmb989LPeKL1yb5o7m3qUkF+R4Z
D+deMili5fV23mYSN07XcSeVvxgfpiFIWLq/3vaU2xBrHnRjeSbz837RN7EAtUMh
Yo/teOwYi4YLcEgNvZkGG2ZAcp+TDLGd+6H1o/v6gL2haNtleyomeC/KuI4NVDYq
zvEITUXAGThiq2HlgxfmJGmj79VNidZ/qNm6fd+06lt2vM6JQJ1iuCLAkv5QubMW
rGnAvWKoeha3HjSvi/WoYcCoEk2nWoTs3gc9Lr3Xz5wjEqN/MdgpRww59s6rdvCV
cJpp46ShAMWEgrHbzI6YOk1fx9B2YgquoQjO0F+5wVwPDcdTjlgJFDSo/m+UkOtB
i1R6/NEXtf0F6W/cEAMJezpMWS7309aJaDMMZwV3IZmP4lDA1JbbVDrhG/8gytCP
mGP7uf67M9oL78R8X77mNO6c3x5itytPBR5KYIXQ45uhAG8vzsgD39ypLIjQV/wJ
KtRg9NXcKPXo6TuHLnA+0vWDBTh064dE6vDezL9YX5aeVwzkiFtW1hO3rBwXhJOp
K8A1IjZk19rH8SCc0TPRe08+UzOPfAedKGlhaRXGlB2vA4gBKLRDp9g9Niex+1Av
zYld5rjDgh1fls2dT4Lo16IcBY+EkCE3OJUg/KUOzvmTeMTYovYhJjiA/Ps2KWa6
Ko2OIjCHshbcq9hznccH2Fo3vx9TUZJJS6EMo2uP7J2SmgZ3QX5idxtsyTuwB38d
jD/pTI0w33jF2bEZRIM/q6sxlIW9/3wCt0aX6QijTBCBCKF7CJuQK13Q6qZObdaL
UYoSGTqy2QY46iBAZZidUNkMYoIf7HTaIzF0KKT+6zTUdxZNbdxvPYfY8BuHgCvj
rKRgAqnGcJi8BD1UJyq3mGP2L9oJFHHLn3Zr/yBoC3I6Bqzp9Iry0lh88l/OqV6h
/XleriBcaiVMNSah6KSA3+4KrQo51D2ums6UMulczUerjI/wTzc28/yuhRfZAwtO
3si+INZUkZkQCIapXEJNfvzXq0X0cadnjk9zqMJdQx9pE0KIau60IboM78FULltZ
lEtPsJpMU7etNZ5YaqmEFd0cq1rNW5I+/V7ivPFJHAt5SHET2HFrrusSADdn9mmv
aSIS37sYtWrtxL9QR5Y+CYP3tUCwGCmcUcIWhvycrKVzwrvP5dyjGwUbGM1SEY9V
iAn4kOgycXoYB/ssZp70JGRrpW3SN9OzX2JlnUmlKZgboOr9DQJ1trNBpjQXYTit
5o3kgyjOtv+ZTYLCUY2zcF3V5ciKAHQjoZDL3D3WaRc8Au//dWpnZ/DgNZqzaII4
khO9ORImDvf037ggSsZKfAvqNzJk2idpJFL8vUsuhYjxDB61oh8YQAUCBkwLMhqi
NnVGdmC7AmValjB6wFa4ZdzcVq9A+woGjt93d5Uqdb/TxV96OFx/UtmOtwrgXORU
3oRtTo+Fh/n22f728IirVxUCJbOiHcCMOf8A/UWiFxG+RTUYv98phxyYOPOnmmqr
HjWNfLnsmn4cSaClGDQXEY51pYFx7ZO3dfQS97+4pBJEFuaKLwznB+uvjUtd0pdM
jgFEonLh15PeBd7SEZayMHWxqi1IR8FeEH++rALoKb1ACQNdlGX7q/wgdWGu2X1c
UD29ct3IFaE9wwYi26/VoHbsOqgkpsgAFSMbd0BAbHg5snoSnXHxWbyqRB6jfGyl
9/v0spakbSBw5felvJurA1eXKoLXTqNNqU9UQh2CHTUEJ1Qf/huzIt/UAhUqh/Vg
zEJTDnpS+YYPn+XZdEjYsaARJEcP78GT2QNdSMtFUwiCf+Q0DDUi3XK9nfFoOFWp
RpUEV+0LZrMYb0Vzk+zEBraH8sjKi0CJRPvZJaJ8oFsxQPcb5c5zvAfVEvo78a56
3BhyAi85imWX7cEUd1i5BamP2p0hg5m3qLLYMw5CF4sW79WkmPiineTmB1f+zGPy
i+gIAz3tt8nDG57x5SiR+pn67WIfcA/4U4O1joFFkS3MlMc0vpNFBmwHbMia56Dy
YN5/AXYm5ZYwGsqRPPAPhq+wEjO1E0uVrC1kIgfhctZ2aV6HCmFEOxpvRVj+iQaF
df3fZ4DCw/0kagjaWNfGMTBp388T51k548KrVbT3Ab4r5DLT4kv462y/Ehco0FFN
R6RPwglkQHgD9+h6p27yuZfEGx2pNJ/IBToKpHfEXICmo8ES0Qg/R8vvKyZMiiA8
A9BfrLXSyGbVdLY1/SjBDe+HNB4q1dfpL5xG9rRRYjXAsorm0JjRHX0vd7wD2Rsc
dTDUhGJi7N6khreTKAmuq33/l7QqON39tVRJerj3EM6mN8DrqzhZa2/OazD7Iw1+
mauIZ5Z3uXMlnD+iKC52P0eUf+Wn0ivrbFtBUmWaJE0tnGCjKC1Tc63rVWAwGCU1
tb0jCse0PJM8hyOwWd+4oqmptCW0XOv4ePK2K/zF5M+WiyjG5ZyQYzJMnRjKr159
rh4srJLxJlaMhaV57E4TpQ400X8mmTGt2Up5NjfSo6waOg1iGAa5uZyVFxokXUdD
w4NnSBT/beNATBbeQ5Bty2rDrF6LEwwoAIpv+B7Fz//42hdd6XO4TDtu7T+Is03c
7Rguba9yQH+yekGpzFVTHk8IBFbk2xOCYaeQ1SkzFMzZdx/9RqoBEWdRUiZh769Y
MYS0zctksaU++WjnjDGnxW8C76AhxXsUl6wmOiwKGK6Ck3dflIhe+bZg6BtgjhJV
H0M/Yejc3nHsrD4nPhG+cPTDAWIrqy9TwBsXpdbo/4Mc54oY88uiYf38/zcUNsMF
Jd4ZwCIUlvLmiis+nzC8SJGW9dsUmfuQ5DdlGirwsI8lEJd2gIZdFvFlGUbSfArr
TJE/GySBHFYu+Syq0DM0nVxMQCQ98fOxhz+m/G38O81xLBsY38iHe6eyUSBn/k3H
912HiM/XvW4VUsRhBO34HDt3aWSrd1fL1OYCYiJeR6ELf8+K1CV9paMQOLJIzbAl
dlIqmlSPMZwWTTGn7DYJ54CSNSK92Vi9uXR7vnO/V9V1T1Ly5uHJgiXWMfxbbXjm
CLRaqGQ7KppSqf+5fFse+msz0mzmLJgJVaqsSS+qxp4U84WE9zV/vRCApaCHe0S7
pVgyiDq8xQ+P7qKwDYa1lou/3hyEUbYGQI+/xJ43nqn69MagwtJEWsDHM+HnzEup
0/tpf1V06C2ZMcR/ii20joq0zF+fjGddWnUpA0ZOxHjRgk8V9b90PNAt9ZfkXFrs
Rm3pJZzJoRQowpumYWVaAQp1f8XzCY4EKqCC9VhTteKydDkVx6UXJXMQH98IyYp/
0xTNgAS9bVHlgfqNoJQJuLDnx98qgTst66omVkVYeICOEraMlKHmzmNTd5bIw38R
kPC7Vqa5dUPoq442R2pjSss9EYfKUBa+L5E9sNi0gOeGqP1aV+OBMsc+NuoEpoHN
rk3tz++7T5WuiJz/YmyN7GCS17QGCNmPiPPifHiIvxEixd8TT3Z3D0rSdoytnErD
f6q7AZdyeOWN+pS/PLL901xdRHjUdsfT3d5lhDenZkuUtDArjEBgaWvCaKGWfBxb
OWKSwQ6WzCfJrsqzoliOGaBOmFHbfIvwff00ZZCPLKveY18licl+yW20ZvfPdrT7
Fs0cb0d3dhNEUJavr0v2ltDW+ym7lfN10JcpUT4hdN6Zmj63QwatGwBf+Aem57+k
ZZTQkABqml8/ax2uzU18xqvk4q58P0JKrhSC+F1AziQoYgfoRiJa/Q2YltzsPu53
M1oRS/eO6tkYL/UTdkdknZLAy3RvZvRGbWrs5tWlssyzKF+YbQGidKUxs3TzArzW
HnVn/yp2IxGfxJdoDDCt2aF7u3BQdJHzJYtAjKhcfm7to2NuhAzapPA938kd+8gO
R+sB3jOlINM0t1k3PFWM1kEKOPPx3chlbkGyE9Eo30SLqA9AIoVXfaQc1VmM2t1y
TM4Wkm1FHQdXT46+87CjrYlRrlllUFH9ZcwDIeN6Q366W95pgFpXXNWWtlCXxBwc
e8bOuYBUgO7l6chYi3/mfEDNEL7B9ivgeNBwTIMbWY+S7D4HL9zya+3QM+RIU/oy
fSGXn+/Et48W4xc1f0EbV+gE+Z6JauKnmsxMNhIWlst4Yw9xsSjiLAnPaZQaaayi
9OwAJtUoYLcSJlUQEgLpO0s0dzNOykAZLZlgqb2NjgvRK2nKVl/LZotvQOcI822m
wGTzwKlg1PbIJ2mjtiO2+g1vwivRoWLDatPjb2axEkOGlxuOeNKC7k3/ROzqWO86
kNt1qMjV23YsZA55+CjPiMbGDvlJVLv+8Z+EB8NTKnswrvkN4czIELfFHgcugiQ6
TB50M/AVNjHBQq4oaQHkzvhsAYOtmQFuQdIV7YIpNpHtC6wji6keLCIWC8TVsgS4
qSkHOg3IfRL8uQYMRZ1KN+U+B9Gve1DeulGnZJK+340ZHFf7acEXRP/ZSSPn0B3u
i+3oOvMbqIpsu3GS05Ck0AfDDBiVaTEqoJLS6KyuBRVYmOE58feVIurmAwAJ9BZ4
7SlLGB5N0HO1TAOV76moz7E6cjQyAHXIEt4Wcv0NwXUzV0QgAGtP90gWvfleMEEu
i+85JG/r1yLgGAx+6uS/Ydk6dFUk7rGhPXTpBocGrv/K+xq0Xlk/ZUHAGCcsz4pm
b4QL5m3u/YxSf7/tvO6ID/xwv9IBgPL6Pib7cMMGF3EczmB9Al9mm1M4rAfrS9Vf
aKEN+a5TM5mJWbTbWwBh3MhSocsP8E8xxV95bg0ZF7a4HCixJ7jzxdumQqK0HkjV
KPZLP+Tqy1IP//beaVdhxO/e3GRyIV1otOGkgEsGcZcT0I7SYMxg3LhkMNp23oL0
GOJKNWN8vy2SNKwu39c2AsQOBhZ4fYLUJDp5bIuL9IEuFp+c3PYAbvtmXx0ZX7S7
/e3sFpcUWql/1mvq6nqJPcnOPIt0xRru+0pYi5REVrWXRC9DRgcbT9bFPzdjxBDp
g4O4ae0DNsu8rxBlUV5265LG9UUcJX9hFEG55D70stseCApNj1Qwt1+mSie6+aDm
Q7hnG5xOCVqD/XiOA+RnoyFdzZFoWp1f5INYg/3pW+rhL+/wcR6PR+8ivx4BEtdP
RVJJVGDMzTbuNFnfndJ2Ud85Z5ROKJNrMQRiCi1pD4zvDrP9e06SWTkPeyLDVSRq
z958ALZHm83HW85EpAgxD4cksA5Of1C4N2s+/zXvW+OS7mxdpPw+kXFnsxnj01f1
b8e9HDzip9PDdrENMiKOLhVSrEPj29h8+nFiHfsSWWSpso7rytvrqW4eBZXiKTwb
PK8cvdfjs7vR/b8nY0SKnI0LL7sA7rjpXXWt+Y2b5Uz3WqHVjl+kUScReOvVGGL2
/1C6D8mHoR+t0sUy/XFAHxIGEow7SvW82Xihezcah91AvX/bLwQqtKKLmu9O2kWj
wQroJr7za+ZU5+0kUxDJEHWu5VFUJugTqbdWfkfuRKbSyz6Va0o8KD2MuXK2+rmW
3jdLw/OAqEAcGRPqVM1/NmB0rD1pg52bhPET9vbSIiPSSPhGjoGGz25Q/G0n3CFQ
28AfbFzDbk8RpUHM+Acxv1pDKxXyAmcg7hxytY9cqZxvxEPGBcIuFu6cf/QYINza
KDrbaHYh2bs36CHlANdVSfaGsSjGpV8t1sgd+9bPY7tJCLThkNBENh6LFPzqnk0P
fJItVbrZj+C3/oTefNuzc/ljo2oou+QUBbdgkorM5NLFpAKbMH/NHwjE/Hqk8WgY
BJHCQzq9W3mlydn4DVGN6kaiHslZUwIA/vNQh2wq6+kCIGXoLsxG30VT9Qq0xv+o
codGLpTFkYcULIeJsLwHhuMjGk0alNTikeNQjdwdxElLd4VjT9Y9oiaDBlYMBH4H
buXiLUYdSTeOlmpg8WcQh9YFY5hyt0n/KKPLtteVABsiPku37oEzetoVro1/VjV6
spP5N30rMOz8HBpzGiaOWIB2amcGXwqJUW4oP5fALyNiyWHjkMuSO7PZKrDIydYY
iDREeT7KnSGzGiNoffcz4cG6p3f9suFZntR5YMDA5ZxAxaezFSV9uUfm0IRZXh6B
/gXcL7JXZ0bSPSqiAj21EvH3RkbdwEvBggq1klGS+dxDLD8aJW1cT9v6nDJ6orcm
kMM89JtT2DEchcKzDMlZPw==

`pragma protect end_protected
