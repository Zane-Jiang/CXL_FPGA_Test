// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OPIQpe8wSlZMCsiPG7tYIQd1vx3/VajKMBCNQYcypVl1Dlj8pQcFQl3Jq9y0
8gGE8mb7ixZeKj3Me532KQlQlfAD+gB58PFaKhGFiZzm2K3qaSDTIUHkD2Bf
DRLOzHkaRQBKKtyOtGwVuiVjn7mUWNpRMiw2/ZfKsERyuQfoovBZO+tRm+WV
OC9z4LGcyJVBHIq5SUSJ7qdHn53XXSxYdaJRC/7M4XjMZ1sXrMzs1WleBG0X
Qto67lw/PxGtfo1vqMP8wrhd42eBEmgEzhYSaN3Va5DwlcHP3kuWMPRNtxb5
WQ6W+cefaoXtfLGcJs430mlS1KMkx/8iAhOACq7RVA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oQwnVBVKYvlmuQYx4twWXg9YF1rf79iA7QxUx8bksONQzq4Rlh29pyd0KNt2
PhKF5w5H2wl7VuLq9Hkavcuab3zJDiXbsl78g9FYYw3IfYmihgkODkb2hqV0
neHJj3qZ2H8RPtszobXmCisGjT7VykerImx8Vn6tq2vGrtpYijdDeguqJGtT
KEDuq1srwdDBlelxtGeqqeYZrC4d8odyag31RMDThZXi5bpYg81gJ9QAIosh
LXGeeLle9Iszi9QSiumYJtTdRcOAu/QWjFdp0hiOxgEPzKE9bfN1a7IorVYT
/zmp5hGwAd3Noj4rvBfGEVgALhS7TtJUh81at8wUHA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b6n9kXzoV2I+DSvGyfY3/M0LP/4XkYHzWbrvXMiuhPtXVMBu73oRu/AcAkPx
byX6iNQ87Q11OB2/nG2RgP4OBqwN60Hczdymqhu/nUJgvvC5G2BgMTEwYF+B
7QteNX+bAGzplFMJVV4t2bRqoonozUqkMEUjyobFNe2p5rUhjM5gmCHFBfMD
JveLcvFnNl6wS18BedBJNkDDXVZ7m+emNM+ET4gI9ALlE6+CgVB3kVhOPrG6
m7tvjlS5TdV5CR8lBiwrpplnv9rEeX/hiB0GX0hv91dByuvxZZCBjqZYWWDM
46ezKD4lYMYrdtCosVwARV7sLG4NnOu/Xxh91cDqWg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m4+mMcMALdgaerB1uzUtfl5F5b+en2IT/M307LlGdvdzcldM9BIkCzmsn+b+
+bA8KiouPN4MU7ZbzGrgkFXia1ZUWdjMm2L9e9yuD4XmlLCnuyPEHaTRAWXP
fqgopVwefrCJaLL6coMyv5kOcJT/HyTKRJTaH/PMxVcir4+JzWA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FdyX1lbpw8SoyCvBBDAX50j1n+f4nxgVDCG3tZuRHS9TeSprf97VywRWACpM
F+h/hcsWcEYN2dTt9QPqWvfoLs6LzhBpFtTgXN6jpiycYxsloBZnNe9l1Mrf
6n16z0cClYAixTMUEUH+EXNWSc3OdHNGDqO2SNK37lJBXR84aoGpVxpZPTSV
0BpLVFX2KHjLc2nsdMFnvNwB+dCEaomDhQGHEnIbxICSJ7D8RtXLjjGDfRhL
FN1U7KUvu2ciI3HaZzmyaOk6nxjhN0+mUBebnLWj3omFMwRQ61kuLGrHZ5bm
uk44+dBW9f9pN79A2bejSMp8sq+SWd1UEUY1ooTTxgX/8uKcNJvP9/7twG7W
h51SiW1QadDLf5JsOExemFKzUphJZ1r9mDzIlxVQVD8X11iu1Dk+Mq+6rZ/n
2VTy34asyqeiHjt6zlXKsM1i4gB2EGCKcb3iQ8rK8wnwVVwC7oerwdw+5QGF
/MNGhODOUUnYKw3w+kHR/VRqmcrBUJM+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kV7UBJy9Csm6MFDW4XY9juA5+JWzpflVTod9ZvEBqU/NjxkFBghU0fsTBwrx
nmNlMwjqgxyq70Juxn+I7xso6EpOEpVsSqqI6hxO6u3/9AOQEPaM15QwBKZr
uzqhLRjSj9znydBTTn9x5UQ3D7em2DDcpjMR7AMqi/Oz291AYGo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mznu4ZKxagp/xAPvF15j4kR/YaNyKgEOwzeUSfNq6YMCYh5E/Rzejf+k8Wco
rSklMMBmxyIahc21IaGux9qpnfSLGLCRgVd/VzmzfHfIV29pC1NXdgEj7JAw
SmonDJmombbzTQO3nioqswdtNFMAZo+ScDo8TJj9KyPwzKQsW+8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9856)
`pragma protect data_block
LD3rhTEfTMPSaoumWvOiV4US5YYEkRLptGNVi8943fxmxsdsi6rTHNb9NHnV
yCR5FEiycEgK9H9jcZ2bHXqZId6ca1M8xkdlg1hDngzNOvdRgo+z6AGpfUi1
sVPUrU9G+eyfDzHcU9BB/QrKXXlcSkUVuKGvNv9/XxqV6wlCTasiMEjZCYrV
77ygsmRpzcFvJxEGuaDPneWafA/h15GIFz70nVg8HdRp7cbybd3CVNyyGAe2
GtY+1ry02ujYNF2nB6CgkP83gsvBJ7u04Zzy3AN/JBSYakV+8D3plvlYQGb+
qS3qLsVnLvJVDN1LyLTigcbHwkvtkVzBXm0vVV3We5qdov3EH2+bu3Wm0ZAr
tp3vjb1+hw3e5qevb4LKsnp1uS/9pCrYb6rzfYkjKt/CvN33FyGilwQMfgYz
pj3YELUNTE1vj18dp+r7GfjV6cYvM1pYDwrCAm4wgrdsUAdEaS3L1ubtAbQd
6yHnWUL0dlfCd3NCK0psPa+wXof2Qis3rBAUQUpWv0kI3X7qVWur8QbQr7j5
R+BMSsXq0l/yfANGZom4a22TAgXtzK0QDJa0R6vEi0OqetC1TkAXsUEYJUJ/
7lNxGPhSPI65vMAgKUvl9hmhUsjDWrWPFqod0nPfMpfIh7X+jt2bEWqTwLMq
53Bipsjl7JtsPOjP5kbld3CdinZgCy7D0bTnz3bkWwSY0EKzt4v7CNmlkLPR
RGntl1TQKN4ngiBq4i3fnj6yDIqkRN7MCmlWcsGWezCTBYE9YyKQYjyObrOX
TkNNs0FTw/WcnOKJGwRPPfuEhIYQwyM3RSlwXe7e/G5zaEclJNHHWt5RIWkA
CpOoFvVqaYhHfQYgjeEfS8NvrE5jMjdul5J4ZXxMeZU2r8cJ04E6eA1/h0nw
fkr9ThNp9SqnZbj/rtiyUNmZ4ZuI+sbm4qvJFqc16yRsflvr6dlbKJ9fArLI
B/1gHyqisRIg0JBl7zDuELl9FJ/6c5HN0RurDrfLBICPXoSoNscxnErcctH8
UU/EHpvBR2lLVajFoF67l6d7LMYdj6YhKHkLohfrcs1e983/YrDXQnXsbgGh
d3HyjaHbHJYeb8D74gRH6B5EZ2KnCHpoGEK7SiVPT0RrUCHaj+Up5xXeLXAr
sj1fDBim+xp206KIB686y1qYdMzRB3ss5rwqE9mFstyEIuvuIMSvOlCovLOb
WqcPX2ET8Lra3w0T3hnxGfw4ZvJj6mYkezSrGsbf1hAVSEfj1umxDH1Ay6e+
W9GKXAlADR35kyE5aEKPykZ0bqBr3/+4ZRg3vNJaLBmemtLDZyNHeXdGAHuO
poD+4X2ZhCpyJbryhHsFeD63qxGaOO4Pc4aRkR1L+9idYEML4QdCtVbmF3dv
C4+a6EvHL93BRp8qpbkgaDKzojdI+P9DxPIU5Iww5kmpSuWRLIft0+42GGYB
mlk1qJe5rYsSJW2jZlRM5KSV0hbBL+foqJ6HaEntJS5NkNIpIAtMaCfYCAgY
CaYQvCZSbrNbYqj/Q9w7WTDn8fxAdjdzrqiekn9s00/WB83KpDY1lL7k/l+c
BDwaYjTgw2JlXfj9TUIH2PDryFNYcNAMEatsZVH7lgPxR4KOd762w10PEesQ
dtwehGYZRblMGR1txqiiqzRsXshflOBJYYOAh2BO27RLnR9l4EFsVcXdizzo
+mdeJcayZ0XqQ4u2p3Ya22MeTVhmnvLYHM8603JK2sAXVCfztPTJ1+lAzVsF
q9JU59ryROxWDvOyyyfNzOcxDKfNMGTyyHxZn0zuUdVOpinhUCuU3+zDhrXZ
rixgvYqiXvtwzKYfEHhrG/KdRIlE9pDRhuauVn5NxdcQyKyzqvRMTltRU37C
01NGZSrJT+uNHleCO4AoCeJJaeIZyd40K27u9hikIX5t7aYC55TpFF8KnpfX
IUSf6kKnDQgBAM2EueMb87ZoVaLnWirfZQhiZqVPnLF5PUtWZBOHjpg9xJs3
oY1pP9JVLeGMNbeL9ZfrMsVl3AiRxVsC1IukMZutoT9Wx7OQhhEEkOcB/gUb
jAn7GV/VLHXNsyCjGNnOvn7LF3tdHKMmxMHMuWD5AyF019XRPFPhFDrdqKiF
QEn74GvTGD/f+scPxZJuvO9qR/blC7l3WOkiSlHtNCE4Fml9b/lqYozS9US/
Wgo/a5cUqVd1VuB6NGo++lJSPQidbu/siWHGNl0e77GyyTw6pWU+eoDiAAtR
XEb0eybYPzX0dRFiSH3VQEfJgF4qB7JVNOQuLKCB58OfYNLxP6WBcn7XD8Jh
pSeFXXG6AVPYHfQv/GXqEXM81MHd46w0rrrJZnMv9bbHNdrBC4RJRqVgu/IW
dzYKtjxtBn2HyBEQPMJV5PwPbrGGOJ/9uK1YMhNwgzlK6KOFr8grFz3dLw17
NxeijDo/ip5N22CGPSTlvz8wfMhFjc9urnW7FJvbb1WR8/sYreqlv8C1wG34
lW7F0Er+8Zx4S0xIEgt1tjA7kq9htU0+x/MCN6N1hG2AV1IwiQPfrct9+HVI
EIXJn8PvOIJAiUM0Lku4iwIxda7gO29BRy7cUXilV2K81UvvT8m3SsGwUyAy
py7vYk3o1/vt/enEeDnKe0H1zmFnZjq3Qk3KFTorkwwtJ9enOvoW159Ah3TZ
SlKkIHpCNIPDnwA84rkCm+6FPwnMtnzutEXg6xY7llHvOrvoh7La91xVVeZy
2AY6GJY/oYX9+D3AsrD773NemR2XCuuStrWyQ0GV915Tv0/UPRyl9hH+aXfb
gJcdSTN6496ptiu5cbeaKmn++GWLTPCVaIdCPJIVeTA+9/BtpcYj8Jnl/kw4
bPVe4NkBMGojoaDww+lN44yI0TxXONqhsV2xZrmoy8DmtgvuCa0712GPF1dm
rtMiD2XiJ32Eui3GsV4I4ENeiMR0lrRoXbUCpIvAf6nU3HxuiZHtrHTn1ciL
BBcSmu32Jes9mzddoYpNt8gXs+rxZNNqwf0B2idLxxVVzw4Kd/XpKm1irhSC
d/CGijKLMgmNkIelioKjpRoebSVAS0c15I5Nv0nWLRt28Yaft7mUhUR3PXjk
kjgvDKQX5Xp3kDscpIG1gD5z8JP3Evle609+Z7RiBtZcw+0eV0M5ZF5Y4tFY
dmi8MznmED65nmlJXA5RS5G4XgroIf6WF2ypwyo/54rom3BNhoJSeBRpYkDc
R+qlc7PzC/FIuNYBV3aMj9GbauLDeQ/aa3KRXrJVEermXLEGdsf51xU/67dT
l06pzDCqleUYj503wvS3ZTnnwOOairWkZXpOBREIY5JeqN4jRlc8np2qc72D
3tkxXCqvAbMA2XmWz3X+FX6aOVFSiYDuoH+BfeudBKa1e3/PLETGez0f/+pQ
jy4IHh5rjcWnIBjPd25GroMeJnKTGbiGFJPQcON3QljpSm534FTJ/JepYqJl
OaaT51E6Mnkr0IoXaN2Qq7MX2LDAMRQLoBzmSjFCjvY/+WU8EallqXiC4ait
6x0lW5zo86uBGDMZ/LKey/upiVHvetNg4te0iPNMn4bnqiXna2jb3HA34eP/
S3TZeaJIS9a1FtP5Bt8BTP1Lr5y3g/sR+qq3DJg9/a6OgNi3nJWnYrVBaamd
oXODPwel4JZCsSljdkPzTuB4UuFrr0wSmhgEx5YsIpvRBUw2zt3CQXwHmuRe
6/yb3Fds/BDmTnBQcHdnXY2z1zE1kNvN9w3FZS7LXxYw8P/sKE/JSd2ktPBa
AmtXqc+fJtMYKYeF83nke2o7JR1KavICAPhX8AEob8CHClkzn41LiKDv8GCc
oUvzd8yo7DdwSX2g+iGsm7tkj075tr1H5YXHqa8QTu/k6I4SekjWEQ8ih8Y/
ahuB0I3iAI9aFbXk/vgCNddomx63ZZQCgum4Ofs3Z8PDLdDxjMlD3q4V6Vss
r5KsiKK3eHpSgIXcTCMDp8RZUKuos8g+gYNsCuPR9RGzEm6gSgKrdJssPHLp
OsZUNuKoZiwiJRd8ZIMaoFTl8ZQ2Wudu4iq83pricA9glYOL8zijL80glfN1
ha1AZ/XtTu0Xxg+lMWA1mx+9Pp+roAcFxo3Wxq30cAL1fbYRnCt2voeP7X87
YNfu1P7Pept+nsBuuNtiEYVRebT4q6d9YJeQyh8DtdDMXsKRIcvRdhSzvJty
4oz4C+HMbzCiKpkcLyuAMEaYq/owl0HIOdoy+gOgvU0cjuvk63xAV/6oBsAK
2HBwmf1gVUxv5VkFsCqH7i7IwoxHwvFKM7bUPwwGjPdik/gw7Opr0mO7xuvF
43spH62x9NG406M/BedISCLzQjUAmbIlFRsGGQMdAydfUPDvNIWlNheqeNrg
Q8cLlruUKxbQEi9pKiURN+aPSaZvuWKGUGgDNznU3cFs1TPOAhTrjrRVC9Dj
tfAGl8l7BJqxqRcfjmNVTrHZDts3n9DyUUXM+QNZRAN9TdMr16kOnrqyIE67
+TowX7RbfjYBR/fQsl0Djd2WSjSF0Wq30gUjEVxTY1WFg8EL2MPx8XBgmLt5
SKYDQZ8eSccMDL9pBm9EKUvKzvanb5VdPT0iKPbhNLetQ9ILIMjDpOiUpY5k
EDHPvmLuoTCfiVSF2c5Ebm1lvMIKdbtxx3GQFRMRIIgoVZxZIKPZdzWN6vIH
GazsRHMYhUs1KiIgD9aZ0v08et0zXlb2n63ZOoZgn7eIYuNYGH2YtDzbXqj9
FidNdqWyDM7mtbp8riNHUzi8svHYdA7fp8OlpyJofvzgqxLQlEbtHkjRm26u
iY7AVUDVyWIdqE8BOrKByYaCaT0LbLX/80DDdawtvw8ido9nsrPY0ZVIpdG+
jo3v9wa8izbj8aPKONQCleCk/VZ5R/FP+M1/easSwClx5IkW61E2DKzfxHpV
egDzXheJEmFgRlNSIfkHGgTqNDEkiQPk9hGdLxsAG00G/BDjeaSal0bm7LzZ
Yw1zH+345UFfF2uxHI/Htzt8tiGSm6s2SltDU91FCn3iXrnq0S3CNQ3Z2fEE
VY+AOMnL89z0GNwa46trrznNdgZXIklltLucrsIpFIqdl41J8qXygJx6JlE5
qBL38lAbFl3Y9Eo0s0l6SHKHY3ZWmC8Eh/qBy6UeSDTtEVbNtQeFJ/1svSgd
euTTeXJq9fXN8gcFZYBWS6xuxhVDvE3zPCgj84ZQtW9HzGTFHcy2/shxSTKJ
hEe+aX7OWwhA0o8wxwVFL5bziOS5WPf82l+2TLZ2+lojyamIrEndrcaJOagg
Ptc9ya4tDwah/cgES7Lch73vlowPMO0yyTsXELl3pe2PmtWQ/IzNnH5qGjWz
f0ipbbkhghnXQCq5HwCFkJuvKNhQv/BO8q6GAK2zCnYxUnRpe5R/4Q0/QeEV
8fk41JLvnsddOn+QCNmcmISdCtr9ZaBHnbiTGZQ9oghNLYIzTR5zXS1RN1nk
4V3Ybwr772wVVsc5YFqcEwL772jaitN/F+640vuGL4iUwvubrxxQS/uTJaZg
d5wbBkAMve0vXbknsWaQhdZ+Q0dI/KghvvNeKrwy+5Y59LzkovC7zHKyWqMx
8+gs+K0K4WmoJiqretGRQbAe/xCZ62udjND/HlPQhoEob/BApslQU4VqLSdx
kG54a8E1xje+JALiR7+UunKVndNLv6lEUqWKMghkYPpCEH0YZF97uNW7jpa7
ks7+lekpH367QimcRAkXbbhUfVQXEjnHTJnTJkVQi9IStgbfT7xd2M4yxEN4
dgdYgfsBMH7W/Xe+gighq5TaeKd6UwncpgTbB28Pkbo/X2DRz6MEvbCt2pTw
e+pzc+ngNC7XYG+9WJu2ilkrxaEamQdodlJwgF0jA4IfSKW7zJskJ/YsChpJ
5UKtSixKV6euZc172oLKhftS4AtiZTN4gaZr6Uf2rXKjiXqe9Js3pAoyXF/Z
m/QvpxzFgn5g3PjiW+Pv7tAUnuJuxQcYSzFtAg+7oksb88+GOEyGVihPYXjk
EFNBaK3pbc2IV0taC9uTzaeS2LhupvNeXNsU3pkj6o8hi5Nf9WVUueY87LoP
bVr9yBYU6F4s+9kuw2rV55N2wZ2YXF78QohjAvdvWQAWcYfqu9wLyzkspLPH
MHtmHO+LKAaIOkwS2WFM9/50NogzKzHF8NjOu377XK/xvkD4pQS19XvA5Wo0
92qgNPEfBPdkKAU/k8vL43zeA3LUo1FGquQHv1sZ8lS/X0xcy1JrEMIlx3pH
h9t7Ex7dD9KoNiRGtCVlI6OuRgKK9axr1VmYkqpP8mX+IOwipwjoS7IAatOs
4L3p/g9iJI9gUI7gGwOB5WcYpiEOk2aBw8ua8SZkK60TLFg7/rWyeIFMQusM
KmoDA2dEyy6ZUsU8aKnL5MRQFtn/CbZFelnE/+t/DCFAWz3ifJDjIguLMTKw
tl/oanHkm8GtG3tpn103KSLZ18EwP5gTiQXllKTeus9+qE1WMUCTDyTBDMKD
8xR+0bLiJmIjz828Xhb4MMMHCjdh865ZDQv9VrJramqOZQsN3qT0rE8wkec6
9JNoNVuAADX35ucWrZlNFpJZIPfZLJBWmbsRQsZDfT4jMs+L4LnLP5MS4HOQ
hJGrijBSLSpI2HGiPQV9q2TSLU8VHC607VS4xhZnGxmXRaTQT9a203ntz5XS
6AQhPcl4qVU+Qpk82a7J/pFgm4Vw4TkO8KL2ZmsNm1FHjQtxuT3ogasVXHzz
DdQxDhpjXsav4d8aptBMbSuGL1/wiaFRoWCoRcTZvK5PyVBm6fkApcuVA49m
6XpUjQHUZW0fBj3xFv3i2PncOucNyXdnbHB4S72bcCmaoPN336JcFapu0bdp
iUAVTq3xqHpwME7hDUOx+i0c23Sg4Hqj/Zq7CwkMHz2JaH7+RkiuVsmB8KWv
1KsBr+zQRH9vaGjWmXuMLa8ypdkbNF0PW9EBReGz/F8KWTE+YRd8AsFtLYKs
BGhIfPTLMDXq00twRH8PAH65OG9hzG2Pg+ZOmnm7J/Dveo90XT1yMy61vR3n
4fGXu6gOqyk1TSyWg4rHXr3v4cX/bhBPawwqQ8aDhRRZi+76wCdIdQS5SH6u
MKT9BW4tg15fG6k9+zgJQQEXf8ERRHiuJDo0FUsfv7emSDIQZS4Dc4+ZnMGw
u5s1Bjw08XGQVhsi3v6R+oja9qjWw22tVHdAKSjxx7+yLbdlVGI6gSVz306Z
oQc6u5GjbIl40H+819UltaCr8V9jtyENmWopjp8ZSI1LB7bLZjIsFpeyHNQU
hgWSOUQW+Sei/Dk9SwrFlwhq8deE3ldgvX9T6PkRPiQXONNeghemSi2HGCGA
Nzg/Crrq6wAuHR622AXDLF55xFnPD6zrXOuRXAuO8BnsGlBgajCUpekzGU2k
R0czyVvF64uJh7QZnTzJXa9YvJ/bd28vkG8WtI1BcaRyT1fjVHKkICGckG7l
la4aS6WAH8IlkwZt/laMpvM6CVTcjU+mirlHUpcnMSxs13dPicY1ow3mwJXy
zML3IvC5Cia+fR5S0sVWrnYOvE/dlRTXWC/iWBydIO+MREG+QqevCCvGKXbF
m3ACJiLqPUIMKMP8ScIJMBnZn24Eu+fmt0+ncEvF4yXpY2EjMyhr0lTvXitq
UYJ6TCLvsb3Agxhd2jgOcJXK8DH8VCleVvq6JKxoL4BZcGloGIPbIUds+V3+
0SWdQSksoH4wdHU9/6sefdM6EJaXltLqO2dfPByTbOdGUwBnE9iL5c7pcSnd
2kmNvnXRJqWrV+nNlD1c3CzyhjGEum5/GJoKTQSmdss/E2Q0PmQLMICrSizc
6AaPbv/jCaqlxH6PRf5SH5xsixpaME2fZsKKfSoiFl3GWNZgTJXb2HK0gJ+A
FCQfEyKom+xyEORPMU3UnpbcYGcXBY0F19XKu0wN/StnDsrZnEC/O8RjOmMJ
kv4EHsV5f69Rqx2wyiGH6XEas7hVjGgZFu72DROnRXb9JfkugjpbO7TfIcBW
QrSKxkTJiZ7B93q6Ag6d7nJOvvTx3AAXUxY739Yi5KXfJ3ljFMnnk7KSh4Hh
BJ19/XOwJoUb0Oc4c7yZ4v6cjL3XTV6xWy6HAxUHUPn9Gf2OLlsNwV6N2rwk
plYOebAaIO/1TiQ7Xk1mKRZOkchLpNLengV1lT+CDT65XlVwNyRu+6wLqA+L
OQfq8Hjm1ourU7cRuOLOkmF4J2Vc/wTCJpDfEG/UOinHbGaGoScKjqXmubFR
va2nUYM8LZIgx2v6WkJI6Mg+weTghtcBjITHS6/CJd129Jwt/+uGOVnIGeQe
5R/y1qdzNtltFab8WdTtRCNegonAfiMFoL8fZEiJp+AGH/4grFbhcVhtS7Xb
yTiD3Dfh5hnsQh0F+evHXHLZxuZhm1fzK1VuYFZIgmZMkuRsoGHxjUZs36b2
6WgZFt8yXSqU5k03cOviAubLC1TOT23KSKg0ezLzv80emhMRx3AwFvjNswYA
Of9o4jHSzjG07FczyUeu+kAI+Zfcdc39e+JL4Ps0DiUGFy4XAh/CvWCEK4PC
G/IzNDmTV6JXuLaiSPEJQ9Ondra2n4V3UUPBCscKhxidRi4OM0bKHKBlKRq5
laOlI4KKHSPdd8GmE46Rwv2qaks5oyeehgkwIfDG0/U/9e6Mx/Y6sOkzTHyU
hSvAPrDtXdCmVjT9AhqIMQAHIuGgTwP3YOrSQhhSoCAekLbk5R0zvWaVcnkv
R2PUbkcqwWxrvf/dcYwAr/LyB0BKF3qwUiAS5VWYnBpxAjhwZfBGhcPM8/EG
1WBDhcVV3v3I/JzUHALxWvFKkjiYM7GOtHJefVbSKWZXU/1HpWvPfI+lfuah
dRxltbc9etPyalqTVNeNdSDax1O8/i9lN6uXZ+7J1UsF5St34YHMN77JvPtS
PenCSP6wHuXyBcLp1TXq/VwMxhdMJOjn/Df/abqpqZN4/CuYbBzvs10upLtT
H9B6doViewp6lJEdfIeWXn89uxngieYEpi0PnEwaFggV6FDGUiUrCjp0RgyH
kG8Do+I52ZVybJ0AwXcgQC0K+wjMSLpj14GTStI6BDeDdxgkewBJU7YclHe4
cUYalRy7yjyNGHUFi1lIjIVb2wnm9CDlQzmyzdHPl2zGt6Fzr8wli9Bk1NuJ
jtUJFMcwOnU9CIIPgSZhBdrR/qSNHrABtvNSHy3y5MPtTGvQ75ic7kzRc/yE
5cYUV9bRJIktQ6xCiKepnDoeN0ajyu4ztRWturqCM3CZWNSPVd+DHr0zB/8y
32VrTWjZKgsUGmnPFDaCgtviML/K5M8pZ1sFI0yfn9/S3L2e2csz2zuwXSEF
Oi5pBtWxHQ2eQI1sJIKlcRRt5zMThPK3JHlQIh09Th7NBFG8x81ioejjffhS
3w9Ibxb4w+NtPu8HFqO9WZwvnYLKgSj+xca/wCszwq1Ak6hQjg/OxZEx5lI/
G5v8JKudH+zNIzuIh2Qj3/26B6k1FkKxUKojgStkIHfI7xjDltBA19n8dRpw
CpALohXc4KqRNmgBoXfnfi3wnLbq8cQN7cLfZqYUmHtIu+6mbzE+tx+TBnr0
7zlCAWCfegd0GbQp9bt6PMT1AGVgbcKDEh23iPMz0VFMvXbY4RQqlJeFA1gs
8BiWBSWHdbAuOwY76cBWXNL5thmYNhMtIR4gYlrpAYd2m45FwV0IHhvDtXqN
K2I0yJQ993KbLC+hA0y8uvYL9ab/AZlZ0QwFcYhLalnH/dqvuVHNbDHS79Pi
pDbGRJLeJe9WZ0MUqhIJDr4niPdafLFNWvgHpkJwRLnQ/Fl0YNMyaLngZAse
D5dXpc1AxVhtNLTAEj93dsYqZ3PFEi//86e1AjNMwMoHxd6AgYsyAbB+s0Yn
+0f20jiBSV468RRwju5oc7joeMrP8uA5aOtWXWDnyUHI/Q2Sx8fysvFQ9x66
rwfG+M5CQJEQeFh9wTAaoNTAiaLdXGwAKJxtoRPhhrkUAoGD+M34815LvKTT
SVNhhzfSeRi7gusTUCMK32XppPHDPstVEGNzJJrS+U5GbxZzhS2gz0BYMszI
t61naSH7UegtynfpLUKKHY4QDu6tCVcXuLgXGkolWH2U7MjM4TgVo7nAyTSV
H3e1g+4kdR/+56CQ3PbRAtH8T/lJ+dTpFs3IH1H5VgQLT4OJZwkhfvEmtXX3
U1dcXzzi9cMfHrs4RTYCtUWh6jL3oO+7WD41/0yhdLpLXL6/Q54NeeoDzpEs
JRiM6bZUnk0UUzxdHOB0xvBvM1IcvLIAbqJuzqcDNMEqYnIDkIie0hyzif1L
qo5/2TG36vcTA2epSnGXG/LCvZacZcSpEhB+IssoVf/kv4lUNm1lCa/tyWO8
9vpPT+/tqA9chTY2b3NB9xuIHJzpqlvgEIqiYovGTuT+bqbq+XZq1QYJ+GFv
yl557SxQlOs86Kp752qG4R0kmNwDtsTOMCkRpaLJGFgeW8iEfsG7UW1itufa
pASNCqU2EVWyj5sr007WqhO0zC8xe/FDrzIul1aXtChjI48qgdgwuWjT7RNp
vcvgXDRXJiheKk9nnbu8uXKFDgveP7iJEDeCdfxQYRwMQ/PXk1taw2EgAFlQ
67niWZjm7FpOMnG8JkyFdaFi9HVqxcvQ+AyiVg5qwx5xc0yhSpgnco6907z4
Ma4MSx87naAUiPeGRGZdq8DR1apYsi30X3JAol7ApqOud1kPNmwe7B9zRD/0
o8SBfo2ZMG9lkanLwDqISnK29lIi/lpXaB9xK0ry37sdq894YR5ASmS0OCUj
nartjCq+gKIAqesE0J00H9gkJP2+rbWNlOgx1/y6S++vPhpG4JRhjns4/oLR
XD5HrAOSklesH+KEaWXHRlgvWYpEPBWW1S2xzzPQAtcziGyPiz9AfjEvAB54
2P+00JyDD4DnFl9QqNf+WT8TZRkrKoxcn/GTV6kEjASWACFdG4kcKsuG8mpi
vKphSJrQKOtg65qq5DEBRJ1q4nWl6yhsPgCyyLkq6ZzVc1wJUFnSBiawJZIb
++tZnuAWGR3Y8AteInIg7XPUe5wdkgSAeLdSAmsm/MYsQ5o17tZsfF4Q5P1p
pbW4+EC4ikOwbl3nIb91k5dRFNOQBns05jRyzW5/CeWoPCSmyNbJqOc4yVC6
C3FaNtdevXKGnbB6KXO52FgnlQkTSZ2VyE2VUiOfw6UalWxBzhO8XHoMYDgd
yNSDUMUiWT/Q/QeuOVLHI0XQ+tNPGTGq1eba9Wzin3Om5DoiGvlcyhkTCF1L
e4/Ub0pQE7cXkjOLxLe89Gbctl8XrEgWlEjp3qCEQHwzQ3kR6Oe6CjB498wn
ZJnr35N8KhLfxkP+xJ79Z23YNhXZMMa/TPVW2sbdfWct8coAeYlmvmZdOHPs
gdO7CBn08R98CZZrkq922oY5+Aa9Ia0AFnHAYJxOCPM59rfciAtbaZ70xPsk
+HSCmmq6NqJHrSJ/0QnngFlvQVwrwGkDMsOLuVKNf7km+YBTViI0C2i3qKbY
ZIIr5a01BoDm0VqOAs9e/G+NvEDWREn+y1qbMfuq8ww6MGnnjM1cottkOCDj
T6qYYFzpHZeEfhx1hAY3TABX+AyPwq/oOiVUIYYuDRUhC3eMVpLQmOuqoOPA
fAyepusEOJCEU5yUyA5zmka6uQL+7xlUcc8I3onU0h3Bb9SOed4hPhil2eQH
ngJbGvpnAf4fFn3ztXt6NIM5rn4ldd7Va3VBpAiyGTftttsZxRf86HbAOuAY
4busPuxPA9NHtC9ppnHpqoqR4W+6auJLOgPLs4+MumioWYkBG2DbigK8i+Hd
XL/ZggR7zVPa/903dphiRMKGzWrlDENmCv6M6zsVZ6+jnVGWLJ6+fn8OMmFC
F1lXCk+Oi1kH3DCsCHZmDEh//DVRjRO/UHXGmD2pS0XedEqXMDX6PPXuLXFU
a16tuRc7i6mreen5IM+FgUhYO26BQKhpAug9zq9TTTIsrlgAqEPl7JSaCfHd
H2JNE48pN9EnCpWya+jMrcPCYczGKvAsceKYHVKsW0/bde/+DYF8uZxWxObl
7miEiH2XHhACiQtuULF0C+g8PWjpg07MexL7WzgS6TmekwkF9JZvlVZjK0zo
XbWrd2Y4noBquj3+o3M+rD+463fTY5G+bv1MPSeR5tj6NvAYEs36OqK4kBTd
5hX1joRZcu/2W0PFGbYr5xVUiYUpJBsOP8TA5UZBRBFISu7vkIpVG5KophP+
EG6grd6vfau0erg2H9QEulVNjN/x9hmnizgstVWbv3VbS5LiKqggx0sQfXX5
odzFvBc84jrhSV5Voj6B8MQ+fo1U3EmgFnfiOYVpE9/i5dHirhNxK+pRnyxa
SuAVOPzw63BHy7RnZFCGZBSJHudokN6dMlR21A4y0ipl6TtImEPldf2c1B1w
U06dt50qrsn4AkISgHT/DOFO1mRgADxULhy6E9pZ4wUTnW9Wi0QCy15zMUSL
s7VMNHzhdcUkOjGy5zXzX7yjulgHDmP2+hrC1gRtZAGRmSVHH1lWlCw4Jzrg
1CF2FXA1huhH0wphFzKXNbe4yvqtGPjsLf2d849Pc9XkQ/YqK1uWz/C8jitY
Ia63JGLAFX90yNUUFOdHGHPQODlWsyfezGHZXiAmd+gGNbOTQ4JS7vOOTHt8
cEPC4QM6EBflbTSiRFb7n86glNLRlyIpf7b6wYODwToghdvYhbRCZkgnAKTe
9L4Q14u24IWA3j2Z7fxwt4zcpntCt5OJCVyxIKvEqaTg9HnQvTsLiDrhVXHu
++XDtOQqBrWlA3L6DYCWHPl77Yq+onK2H3MYikzzsuAYbzTG//V4vIltrKLF
qG3CY9IiKSPUwpwV2yX5o1kKB0J+vsV/MJ55qg4rztA1Cc3miMb+9UPH/AE+
c3VIA/j2Giv4zgFBcyguAKjHHyhBU38tTQhZy9O7GTYXaQJny6BQ/sCmI50w
n9bIVc0albPVNZFIOtAUrqRwRNiM+1W4DTKqKhscvrH33wjjMqgIIT/r+uDX
h58pD7GbC6a1DFEJiS5UPHUjot1NOc9hhiUPFDadPmM4denXU0JL3O9GspBI
FMiaIjrNxjMI25yRojix4p/hLMcT7TCmJyVE1tEIaUFRoFZrkXOCqyfksicQ
p1PiljFtwrSbIlPaXJyPoHR1lTPxU2YJPkJ6GIK1TYa2ExawdbvEvq6fQH5q
z7VjJssw6KM5J88UyT1cf9x2DvsbkmOV0NuczLwwfqoQTpDIwcp/FVjPNLDy
NQ==

`pragma protect end_protected
