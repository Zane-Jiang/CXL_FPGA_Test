// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DqvOuSMaKhST1E/5bEIw7Y6SuMzVVhxP+C6OzzxSBtMlAmce4/+4v1yA40NP
jY+UbONZ7nBQeMKQgAECgn25X+l3ALxiPKNCXl1D3SilYqU4tRwZCGxVrV5X
W0PW5NkJovIRx+P2J/3yV8ZnkBNyfEuedM62eqgRmH0smg804FZJjwgaL06O
SIvAzfU9BFNsEeh95zk3Mz4re4ppqnOGc/lNQdj7dlpskBHKLMXEAsHsOiM9
x+tQYeaQsRXQsujiP04Gf5003QuWILNVn4XeDNCQdcRKTE9pLvqVffPY9eYp
UMaCpV8uLWJc0hW37yRqWb+j4gANnXvyc0ZF1SwHDA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RuN5KY8CAiYRxo5ffnKx2TzP1D++CeHUJkH9ofvK0qTub5qXcakBw7AmfY8H
M39TWt99I5CDtO0FDzWLJbv6+LA4olvvizGll/FNju3d7A6Pxiud2Z7GZPu4
lNL68s2bMgJn66fX2YPlwcMlqcIAhj6NUMmKwjCwkEf0xHqz4+PdBBvgudPi
ytAaGv9/1bDVudvWwfU0B2EOXBvK9ykHmvcIaGfLPQd0euBP9poIBHC9zGLq
gJNRfjEo9mhsTXfoQCJpmymLd3eMn4gpKou0cILhZMKLKlABZkt14zZnhdCa
QqFYgXdzgXvy7BHVsETss7+kRKUy65ApwcQKVXX4zA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DlDxuIfxkuRc/XEcc0iXtjEkGb9o0n8P9wzmfc9e2nXpg1j2ZTJbmJycQBEX
XH2CF8MC5lqNeJrCa8UHfWWbo3zpOB4zDEn+pMqca0rjkVcdWz6PiWFZUWva
0YgYH+a8xGEv5mcOw+2xeMAKN0InXXTC+VDOZZ15Im+M8izHI5owX9NJ8Uoa
LYeXf5/ij1oC6bwN8SZWeinOot3lFiReXPVvoIwO0/UDafMjftGiF/2LNyeA
Wk3a2pgQKmLBCe4zBFyVuFuXemaUbY9rHzxgMkbI64qFow+uUR+rTfGsX9wK
s+4b7UQ+5+gp3lxw8GJArFcnthkQJR1/C15vC6cjNA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IH4FbMVGEtJsE7hI5yrL5RGbFXNw46jk6m/XJwYltzoEaF+ds9duwZ++reN6
sz7j4qEBtumkwWKpngh52CzvI37PYxinPDHir0wkayZu0IvN21TF8hFb/5ea
FzjglvrcNE1YaZPDPKnqldY+EFpnAiXr1vP/3fh/1j4hLcfYgx8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
YjBt6rDe81v0bZB1D+PTa7qsJLadRGhk4Ey9RDNaoy07dq/h/8KOQTGIp8rl
4LCSd6uWUBbAIcA85VbQ1ObjLZnA3amgCUmxs9JyHwEourbCAK0Zpfztk4xD
Ep9taHS5BsWhpxb5MTXPAVShw0Uqvq5x/6NIP8AADEiIxY1HazeGc0OljoP/
U0IqYd93zNfh210my1TYS/bYUd8+IP8pbC8eJJ9A30Pp2jJ6U+UdAHp8nnK9
IkbQX6EmjUurT5VOvXW7jrQiU3ymU5cimUVaJuQS4knVhutWUqg1A53BrNgF
Lme4f2TELkch/N8U8xR0+K5Vtt2nzT7wYYFKM1kA8Q3buPL5k9mQhg8L3hFi
MBalic+vTW0Nfyf3qha734JEShDE1vuRcUe+VtrsGgnegnpHqCFgEKxCdI8+
2xpY4/ZU8/4Gn/O4WyFzLPIAko8rBW4YgF7fvoVBZqIgfM5ETDny4cskM/68
nO13AqcmmJEc2VnHDUN9JkIZbEjsPMbX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BiMFhcthNoW/n4+z/+wRhcmm5Pbroga/Y5WZU7+4Q1JGmJioDFwmE/P2tXU8
bRM2NnsSmOSIBgwr7lxuSPKufMPMWlYu8NJGv/UrV0h9G14oKG3p84NzvUfZ
AddlwVIai7dMbrBVfDJa43fRxium9Sc1H75bjn/X23y3VNYt0XA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hU2OytJSmH1ei+Of0TOz0Eo8N4FccvS2/B1wZIiHwZ3ERq4LRSaMGwRMfM+q
bW0IYvF3KDoUeV3ICQH4RhQPGPkZZXXAqKHkTmijvVf44OyjKs4K2tltoCnS
GRcILvr+vDGRnIJhvkLSmFn/FyQxqTt5xspFftJyZqlm6ytjzF8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 64128)
`pragma protect data_block
Bby5KeMxjuR09bhcv9kPxoiaRXyMwqPlv5VodXhFDrWBuxhxWU/TMXe8IVgf
uWrfO9MSduJAJ593NoS6qmZnbYIU8tOcUYlOd1kNtP+2jKcJ8JHpzXYrUEfx
Z4hfmspGg3GltjE0x0g3vMllbyjmNrxm2HCT1kaGCaKTXwUFkt1J5qZJLZW/
32CsTU1v3NN/93B1pm1kREvh+sNJpsFB6Nn/amhx1mDRBeUzUhD/7SaFZQaC
dl8swoF1e6K9D7bbLJpWi0tgiq0ETlYE81O0oCle8CGl9h1J8MUP1dCpEeIP
qtS6+I9llh6dzfuN/nWnCbQpRdVMU/KcpBr7Pz/jFXBxrliq4EczlkrP1Lnn
Ua6vVgNyO2ZhovwM38nBXkmYwu3cpV+6Ejqh+Wq2fZ8yorT0xex4scrcdsqd
aI+4K+DBJcMd13pT2v+5tqfqES813G7beZZmu7b/3CE3HGF9p/hUFAw/V4Lw
3foqyuDGEPqFcFCNoGRkv2MQdd4ILBf4o+oyFPuDnolkx7CPLOT1zdXa0G5s
1rzhsk2fihAk98/0tFvfVqH7gHPu6eFml+yg9P6g0QuoC47x7y48euZ2msAC
FQ83FrP5UyJcz6za0v4DKuKCHHqb9WgaXuR+xFuWb/xVImYV96LbwGtmjpTa
R/yl2mN0XrxQkKIOwfH8wAr7IQpS+j2RqEKkTTHFJkmrTJtG6jiZ6ubdY/UW
RNh1yMrOcSV4arblWer8i0FsJgvBZOFLBgEnvogvX6dD4IvJnEFT26KiyT1o
1B62BjQ41KVviWtxwXP90UsmgVU0GNIdpvC3SC7p7lb35VJWaLvvTTgeK6MV
CdY/VU2iB8Xo2sFbGezbM9jubIWE3HREiGoHY4rSESwyFnD2t+/efHJAR94H
vypjQsHTuViihqq5RPlgybPWB87xL8R0EA+HPCX8EWHf2LksNrku9eK2AdYR
ws4dy34n0GlHFHcbHF3VFa8chZo5CkPNii5cMl06Ta8z4E78dbZ5IYdlpczh
mrqZm6dpHpkZZuTjhB4VBIWxr+pG3JE0Zh6AlXk/c0afsk+z7bIpPzTceHjU
dtWb+eEIcrA5LTmQc2uWr5AMiEtFduFgYVF07+PKHW1d6bytq4dJjLgQ/UKB
K90ef2b0fz5zgOFKJjxb0I/bG6DMUuXM9caxGW2pPegc3U2R5SIQV8+ITNyI
BB/8Z2XY4dK9OYs/nIatnK7tM7cf0ZneFVtq0siZFi+1ev23nM+EFvubYTq+
v0N8AccxNAaAmvp9t3OPl/kYNYz646Q+ElHbEMoPQ9VCf+jvADk4Ye6JZS5n
d2vkZredNtG8mJ+4HkaOu6cNVPmQfxw5VXyMWFng/3o4cZGMTdIF1t0VrKGs
hYGLZhFxab8L18C0ZAt4nXJaN4+pLUjLtztQt+eyP3m8araLNrBohFBmAb6V
nweNoaBep3B2Vk2a6m5qzVA3C3lgRqFTyW2wp3toGrXLFhljtc8+nAmUufY9
zUbljmxFReUP69vxLg3+B/Age0ihSGci014GPtAd4jEvFIrymvp988mxoNL3
IXwD08FRRgxvgLygbymokSasp48OIpyTmSPCYz68JO1Ex+jhkayK8Q/jQCtl
GFBegdsBccPo7x8bDmvHGwDLs7RpeO7b8/9DcfgLXkC8sZGOLs2DW4tsQ2v0
bKHXyGluKdGbFRVg2fAQ9/RJls1xvjjNcGJEoePqLek78KkLop0JCYHxG7mU
0+tzwdVRMqFJtwMirrarVyw5liLbcJQ8yCsdkxRAsaCjoQeI1uMri6+F8eG0
Mbl6dFCTvgbt/ixocmqlnoUrTbZ01i6nJxQPsVKKIrxAnMcqBb6QIYBASuHF
1CHnv9LBCkbqWmkGIvkRIt2/WsOjj5JsCUBHmog58TmeaRnWAfoDKbFGV3cO
prg5ZS6xa8sHThtsFPoQtYr0fHJpdBhS8JYyUnwGOxpWxHd2W+IJktBoMZDy
X3bgB1GWnTTNpeJQicnaxxEjDzzXX26UBSPg78EPxmFVyQusocRRAi5WV/73
R7g9ltmpNTynJV1FZi7X2fUDfOn30hk+xcHqQ1srwnDM7whQhN/sKUD62Hpf
zlneJpCWNiNL61iZSQd5IRKDA8AoASNYiOSk/zQEpy+hz7MtigSfs/g5i3eR
ZMsnc66jvOr21Dgb4G9Cyk6IebMGQMTmhlAVhHUpjTmRv+ZXV/XslmfsDj7C
qonYlO4f5c3MZaYDUysH/fa4D9+r+jSRjf6IGB5J6e3dWiN/RfFlF7HaNfDe
albGnV23xO3+dNHlkv8VlxPJh775qGl6+lLB42dYkiM+vFnuu9gNwQVQtiA6
bcb5Hwaitj6oLdeNCDswu/rBpxkvnARCN+MzdI3TNZr6J0cWt9VU5Q26G5no
68tk9MhTz/kkZ6848B0lCgMkaR4wKGBGoCKZeMRA3AlA/+nreEv3zQhQjei4
dRBaVNyqgY4f2atH6MIvjGZXy4lgruq/pxF+vYk7KiFAqx5TLPsLe8gzQzyh
p0yX6c+DmFOGeh3sfS4SpUFcAoQyomhgtgZmCalwH9QylHVywUxjyObyl36m
ieLgcxq6ga9F/X65QHh8U1FoNHjvP1k90QGeQBbOZYnhK1cD6dJ5UskTdjhc
3GES3APpW3/7poThlGjuZoAX0eX7+vS6pkACVxhNJ95cLeLfgb2S6sWYRGzz
hdTsN5/F9KyAy/tyyDnST1pfkS1oEBM0ZK9AtmqxaSWOYLGfahJwPqua26uf
4xuIEcF6QMZMA4J6KfX/d/JVr3nMRrcMKtCKB5dMdt/O5E4MEw5uLXpEOQ+o
nQaFSNf0fGsWaJWStykv28Oy/ja1nmIyftFa1fYbmMryviyVI2jiWrhQUkml
XIcA/MpogxpED7PTAQ792nladaCmLPLuT71EsSK1hqukzocEFW1Qx76poZEf
huAde7gR/RDMCx96VmOAp294IFClBAA+D4x2xGYwMIB1/aZTXTpU7wZ7ta+h
svQ1K9scM2XE6vru9LzFfnMIf/0uGvpmot9uc0xlWpZ7tTvDra6ziUfIlldp
qYIit54dVt8pdBPgfSHqbue8cjZw8Dy9a3EdLx3GhY0T3s4Fm/tT1HsuoBHa
xn0jxB7QRj9S4IJ1eY8yDZq+AETPNW04ZrK8uJtkj3KkZgE+YnF+27Ef/ocq
2NP9u7yjvUqXK0QEB6iJkQn5kl+Z0kxS5ElD1xodE3aih7x1r6LYClKLQpV2
d+nUpVS7cT/G891gUz81un+ognZfnhOR+LT8U+ZV5prziq0sNn240mBQV8l+
0q6YEYxUQ01NzI55YzD2TvESftn+vd4OUk3D1xvzDOlf5Jq1lltNgs1e1kTK
e3uijsmeHwALrBNQ0ZSA1VEhHd3m3/5tLc1HGZkgVJY9Djx9R/eyV694g1Iu
uN+jocyYmzUjSBOaIA7qCZ8qeIKAqB7lt9hJKxYXv46pc/8dKjtCo3HLvW7W
6A0tEHh669eU2a0ifmC26CqyFiFI6r2JY+e27npBxvGTQkLu++4kKSKQY8qz
KiB8GDeWRKfL8OhZ/i6b7th0hT1qDAdQCkG15EVi/oFIEM/IX/LLTaXqmsXM
7XUh0uKH+uwlkMSNFB2QHijJHzN+rm69MYmEYWNfcHyujocD5S9uJ+QKE/zF
q0fYhK+FGy+/eSXoaugnwlMAUKJe++0ghI8eoYwkihqF2slP44rXiTgldRui
RVViRdoddWhMDXdJ/rnIBuW86bAA1KNTH9E9K0NriGdwgxlyAW96wH+jzcZU
wJNf1lv8gvrSSN3RZFajK1DICQ545Pt4cdAf/hXCK0KN/p4UCiiEAj1M/hmT
OXak/at/VVW73mNa+TVLWiPcikJzf5oEr9JhosHRtm1XbD9U0+iaE01JwacT
Kpk7n//ruf72pA/wVY5izz314o63AOyParaYzBd1QTeEkIj6XGClaEe4ibXQ
XgAjPsjVbkjIzUJv5cffxRTq2GXY3NpWTGeJGWeyRI3W88clhP1L0VGkJaWJ
zSVMGg14UhJmgjfrYvE868eK/16Yp0HuSmYZZDIYzT6IBnqfT22ljnARGFIV
vLM+y9kqZ5T6fVp4BRrxS7MVxdfgDUkTXCuCFq0VFrY//75bHGK9MizfhXh+
V/13LFmnXMwCkDHGBeMDq1eGknFdDFZKPiSxwmJ9yMU0bMznBAs+DFbuSrJo
phqTZqTF+V7E5vtTsznYNF4LuWBNxbtEGGtAQUdTjy5IEV8YfmhWu/hCro6g
Clw7txCbuGr/S617jIBmwVRT7bNqhe3nYyA0bAi16895N9oYtKvXZGWfJePj
9Q+0YDmrZ2erNKypY+LeuolTlQHl2bme+pJj54VHQzhpUG98uFeytpijk5jr
sHfqZTvl6XKcVPx9iIbKA1p298Y0VX1hilNPk6nt8R81Mjb2SIRdi/3oJLce
gueMepmKztIxgAGQ4vcVCXk5JEjw2gVLwWJtwBAojc9c6eXFc0uk+OrMW6ik
dDBUpxjfphZkXsSO5NoF7JfWurZfe8agUtXwTcllItxRDrg8zIHCBjfuc7GW
a+OpxzOgC4pVkwt2FnnSEk2IMqo40bgar95/CQXGIcDtx078G7hN45PLsQXm
2JcuP8rn6EaI5iFRj8eMQINX7H4418x1fbq+ApNOKE8kNCfd4XYKD++I08Ai
Bbidg0A0upRz6ISfoiTUDAdyLSumDjG6cRJjJom6eApekiYJtc6483tOk5Xz
ADm2GaWqo/VagxjUBwtcbdQuqcdFHZmdtnjq6aN1DmiEcOa/TGlkkwGCzzi2
vMMvfebvImg1mc1XNDXZU5fljz8h8UqZSkePhv+MF/JHbGk3qxwIVhQeS+Eq
pap/XM6nGSrDgRx5FEm9zmXEFvTzAsvXpX09IOl6fClTKX6xQvPELWZYkmgD
V3z4kgI0Xo2M+c8QJtR9gPsrj4p/qHjOLlvMoDbBlgQ4qbaicaxDPs2ueYXf
0UAx+Jiv5k750rxYkDBgMydr0xWGmm2TVduQrwvK1ahVT9kT16ckg20r9R0w
jc+PVC6lngMqxvJKgFRqeP1Bl0NNBGbpf3ae8NZ8KpsIqF1cfubNw2qVuoBz
xiIOPzj0HHZAuwc9rjAkM3vAqY3QK1qHjZqKriKF/U1DEehIjQwA/uqA/d0Q
MBlM5miq0nQh7NhkgwMTbQ3x7nyeGKCb7pvAoVIVzDECbt18nIVotaYTC0Vq
7IdqznFzkxQcPRNEv3LcQvlWCxak3Wn2FZX7u44E77hvAmxPL3+ghBmWllDH
iQgO0t/FoRnHBomESaCmqEFZglqiK13+dnMCiH90XgQwZQS24MjvAeC792e4
SJ8jQlNXPe6xHgV/Mb4LXR/70NeuzhkSSZHqNe6m5vxofuVenCsim1/yoF+7
W+kytpM5n+2ap5kAGM7zTieRJVn3SSHdFPG+GVBAeHdtISNnqraPSxOyONdE
esK6mRXYQ44++8mfMhBlNNVk9v5YnSdXjpnjoQEdw8fMwME+vg0nG6xYtM2N
WTxDLmM8Nwi+l8oj8UyDyfBwrZMmFy5/K7BCf2R2hGWIlUVRXtY4wi1AMl69
YO/AhwjChfNT1a/atIrTX1O43Qm96Vhl0DlA0E9G9D7D40Fp9sM0snbzt/ZI
ppE+9kpuWiQirXTA6FGbxgk3wXxJqC+fyPX0MOzweLaXtg0pUwhk4t8rDeb6
blqTd9Z49z0i350I9blY6V63v1IkqudfMgzO6FCbAhb/NvxqiWghPPV/qOZs
oYEJlW2Bd07KUxF2ZpGIt/x67WR1NEwb4QUqGXz7VWA1v+yP5LEIYNeeS3to
NomB+6lYlm2iMV3o1ZpUENqQfDX508e3eih0W2Adejn5pADhVNpdCnEQzy1N
7ltZf1GsiKcvYNGujj9PNrEb5/isZ9pHJX0Ux8AoiiSJE29paV8T/DdmQXbJ
X7wQlHqYNxIjrT2M8khlxrvsaLziFTNf2/d6vbboRB5xc5w1fJBwVzUnTkj+
yW1ajCdT3Lu24DD8KmasHuiWUKOdfHQThRkrEbv2/B4L22PSaoI+8escg5RR
/ldultNGjwfFapLv9ZGSaYsRVB1OvXFivRMQvsjWcGRHRWdTsvZeSBKt3Nex
7BR8Bwf5R45oB4dUeY8G0j4+tPeCbxb4f9bWNhI98vdmNBeRaxhKm+qA7k9t
Rbz1pujSpSqXD3B5/DXPhtw59lVtVMDVTRO4mlp2StEwmXdnQOVJZKX0hpuT
SbvW3pnkJA0EBVN6gw+liMEppZv+yg2L5GqBL7rLpYcay9+VTsQcy/ZBs4YT
ZX4oT3d623I+odNPjZlzlDDdC2J8RQIefNLXNyaL8wnfZFKeXWGmLg39ptC+
BaCK+r5POypM+k1EddER+xv0PvLvTyOUQB+G4tEUNr0PLwVb4Gp1yg4zI/ls
MIgxjp2roDdY5BY3aV35Y3oxzSMgWp0FqpmgvL7sCYWvTTnSyWyAQ1ZeMCtb
6dX9v66spPuRTaCMW0qd7gtw4jyfnQPMldiT5fJIUvULW4jsW4WoxjwjP1ZC
ybffFgRrd+KbGoGW5zoaHvh8eLu5tOro3K/usHC3G1UzZ++PfTkzrN22GkuV
Y8k6fX+luarHBmdmxZ9tGj374DMIfWfFZIFUOLxCNGN9tamUSVwP2muMzxL+
dlbIHeQkccbR9SEuF0x6WHFj1UTMfY8lJXcRdNGz0U9t44dgkDKMOWr7EJH5
9VZHJ9CXimPjcANltVmrHq3Z9zdC98VrxjVBZhM6p4x48OsFMOqPwJms062i
4Y7wtIJu7cuGNhi4M80Jh8rNoJNow5jbSks3LrFK3ejL+998NWtbe7+Ecrhi
TySM4O9ocy2SmJiVlyrhBhHho5Xvr6+VfoIiOGQfbbVM/unD18LzuoQodBmB
jaEwnYeziq68eiuZIclu14dzyeVjtNrWdpIi7F0rVfyOGnuzNLE1iJus83j4
qAtDiuJRCY2vDPbzwLE10LZ9k0Rf60irQgH8VhuLVNZPAy5GJIPLpECpCRRf
hTyyrsCHVbjw0KHVyXkDNykv+tn8rJjl2RVES6IqCFu2R99dtAT4Kbyg3daq
4Q/GK8C28XhI7gbCiH1PNJ2l45F1sXOrGo7MURETd12EadDAU7jMjwg1m+0N
z8wnJTqlIBsDPolBfHu/U27aMXsJM1x3UTUtF2yvRcKvWSpTxspnm5ps3t4t
4ofuC1uHJDwkkxgHm4BI5Kbur450qNKVS4NWMVGt83delsjukMxzjhlsv3p6
SmzMe0/HYDrd9FyPGsVOmSO7FCJzVH7Y/44iMKZ25APRpkJ5my9jtA08rUHU
+oGU2YAcQWgUZ1mLq/bcYF1lJ2SZk42MRjJO0pWjhalHBmRmRkO13MK+TXAI
EM5rZ+HwircRbnAleSfBTVlbGvh01A5tLyEMwxJIzMbLJJm/P0v/e4DFfNWA
UostBcNM30fNMJFXIa5UAXw0snHoomCNSvuKY5Sp/VUk2fF18c78Q3ZuMAZB
4MMYJcP0qLj+DjNgXXv+ptAO21ssPRVBssCkxovQKZOMxeHK99yL8DFuylFL
KpOdum9YAmFfSFnaRb6CfeGzJga3tZ3RSV+hfJX4JwP1GmQSbXCNzaKxdKvE
7ICDh3R7Ukdxl9Ftx2pq0k3KktkwzUACBrJhKLp3NrASqkFaGBekL1pRn2OD
fxlnXg1yXxUIgGXlB8ovoXd2QJMuiNkc6fP22G0B4Uy5S7Ma5wFURkGAhngi
MInckZNTQ3rWeOFkXKKz3IWKPZKjY4MubSkDN7gQo+WyCcW2XKhIpS2L/NqY
xSJjC1EWEToWv62By5wI0jrhC8yoE9YV3QTBmyW5dykuuenGcHAj490CebjT
5PGIQQeApVtqxpcyUPqFUSSw6ZPzQf4UpCOXqxrvL950WqUU8v6SEUeBXAiS
OCn/KuSlAS5EXS2brdaV5zpVhvUMwi0uXUV0dn2hab2I0P67IJSrdOwuu6Kj
mL8/bPpVk8RkOqcoN+4WJ3azxxnoTCTZK/kXVkjxO3ejHZzri3RtEeYQk6Pb
qxCwl2kHvy8q0my0lVUMq6KkZ2JdRH46M40tg2HmjUXI9FT1zmxTxW2My6ae
1ApVEEA8NtUtTtHTvU9Yhtn955AUysF7sYPo0tve8qQq9//o1wsJ8h/RMvtd
hVDokzzVFCeRbAdiRIL6TXx4U6oeV/KeM5BHshQ44TAnLA48qgkNV2H9ptwQ
1zpp6m4OngoM8Xx+EJUSDPaTAqaRX1h2JdoMGkCFAprxi4y9HZcc+JEP98QV
2v09zy46oX6UibzBeDLTe2AC5dUH8Ufj7NnaqZElm0rrA3d8GV0hzlX82Foj
iQBbng3KIFwYfDgxyPGP4/7ZsCh+JrCsMIgUTYh8wrEExqwzGgaL2jVs6PnR
/S/Ac1QytNlfYvHJ0QrDb6rkTRrLeb3SLnuTU20mZ6j5apM6EuJVdd0SeOqs
JQS5lZ8mQoGrlbcXR+9DfaZ95B9tHvedpEMFwpZR82v3zaIvP+CXjgAlavRK
RmSqf0/yxQl/OOVObChRYZP7nnVDc7EaQPrLDmqiRddv/E/VqLYhPL7KXIPf
DOAFiYUZo/krjnzu8dmA3A2BVzGi9pkqdHu5I6dpBvJsJSQ1PnHqvykEIWrV
3bMO8zNZ6HbsKq9O5GHc26k1HPuWMsmT2nlr2IdKJNhX5ntF8bJobShk4l0T
wctOumUvHSeir/vOypd7zhS9dvcCf7/+1ZNSSHixqH0KnDcTYrzPSH2V0sOW
YWhiUQ81KZmK4USJH/kJ0i04ner6jOrn4h9lqTJ2EYmJW3R/xlPo7c8Tybdm
9I2fMwXf/6WJfK5wjqVJ2s4Q9daVTMI475Z7JXZMaM1mTjP++/4yXnJcnu5X
9gJ688bqvLAT2tuD0fJ9DIrye4vLPofyfi0JYFLFAs/w/MDH4BLk6bo11JLh
pdR6+Vv9vLaBzuqRcLVyKvWAviAA4dBjx4R7CQEXs0nxeIALyogDI7FJCEqu
8fAPKGYP1asjvHW8PG8YbuI3drBy36PsG5xI2yr6GVQ86q1XwIDR56xEUVt1
di4gj7IB32n24YE7W4XUuam98SDFoNJF98abM/k/T9iiKgNWvsrMbbY+Vt+G
XhyuIG3Bl2XjXcJKpAJErxq2hZj3We0wgV899pk56DKgeU4shejNRTeVBSHZ
Vc80gCE+D7tZUghHf6m5M5CoBXesvOjq2iEuSzH9vVARYEaVEpPcsz1/axAz
6wkYN0gsHzcjYnUBDvyDeE/Q5IfRue+mtt1uUx67mUyglRurOeiyMTzmLIOt
5HnAAYw14lcTorAkEwls8Ikh0SNo58ma/qTwWPbtU+ywJUqVCfu1e1xammUZ
+oxu3+aS5OFKMjNAxXJoqCd+lC/EnmpVYeQ436AErdT4B3xc9VHYODMIXG0l
vLf/xZva8NY+FaVOFZGJvfPxtKf132lFJAAC7w/kMZKiQb+Fwbjpkd5M/eKp
bJOsIk67qx6KaRs3412MDPC5HhL0Ji8muon0z9xws3PWNApVaUkXsbq3f+vv
a12liRvsX2EMJ94mWfy6PG0mVT3OTtDd+qaGzWFhOLc2urHcO2Cs+7MkUIm5
yNebKFcc2cabuPzxfWK2uuv5l6vW2GG08OAY8aHhXPLJd9gtG3IB1ATI0OD0
Tua1hnP2VZsxS/2u6Zr2offffPVgcoVDLaGFdzG4eZG+yaMDiO8daXXt/KvY
AfumrPtm1mD91zq7ik2NLErrGBHiLbeEbAvxfAj8mUl3EfDQzvC5tAbtTD5N
yeVtqJliifAw7SgY+CaqNlZPFx1dxnKmRuXRdybwRmmIf8KrZJJXSSxgDmZt
elQzeIAQvyIWx+6SSL8+RWZWNh2AI49PnWqCR37b0CfOsrOeyHcuLEQwivjA
i3fLt4HAG8+RvUHeCMD8rPCH83Fe9QkiINDhKG33rndibgDmBhYdn3tZEPnW
JOaBUBul1/Krg6yLGGRSRvwTjdmOLvey+zw1EJVQWwAk8rG+lpu97xqzfDWz
mR4j00ZrXGxGNA7npuQgRsybCit1onXvrdVOx7a1wcfFMjl9IJTorcA4JXCP
+aH1DX4b7lgdsxePgrdn3VFtmPPDap3KR8JZUwZdJZwwdpWknzyd2Hn79W+u
HyF0oMFX5WIp7+glXCqtwOtr2DBHfJNbWVlDkkRVyw5nMVlYDVbdseTUGsDK
u9Y1iNupqGOzYX9tkXMhEE/fZniiyILKz4Mkg3SLG1JjtdKYTmOA119btv3l
lK8IxjONDkb2oMmtWsmFQ5JJta4u0aed5+6Y2ExzkadYJq42yaVVURa+Nq0A
q10CWj7ArwnbogooKyvEBF4K3Ee75QIxjr/bxXeagNCT8I9sO8yGvyAKXA4S
YNFlvFusZkfoI9+RsoF/OgTtt8X/U7n1J2qtKYQouMotHuDTOQeawmiz2ojR
A2h11D4u7BAsUzdws2EhjuUvKBFWsZhid0m4yE7UYaf3yJWlkjzDfbBjQP6v
0wRf4JjFzF5YDo2mUrgL5yI+wk0V6O+XcPekeWa/bu/zIPAKZXnQJYEV5Zr2
kOEnADWtvUchN2+GkF8lUq0CFtY1hy+oRxG63yzJb9dOVmOX3GJKxb6H6vwW
Fb82tnWR5fswoCO8jtMT6sU/vFS1TH50PB4w3NmLYg7WYsmiz4GCq9XTLk0q
M45ntc8/o3NAqN2XU6CRUDaLeSEgiz6lGPwWX9dp6ny2wmklfYoB9ZTpfp/U
pzoA9knXZzCrr7IneW07/f5w5pFd8ho8QJG8Fjz81Klcy0ObeQpaIbznRAjZ
RM4JOnyFP6RAzmZLV57i5C+z3vhTh2Xwq89qqv97njLlORj5hHFu52uE0cPQ
+bovmL9a/W3Qfza6H5Gv+5z49uknASN1C4rqeRg/IR7saJOMnOEFQS8C2Rxz
OGlR09gqB2pA4J1nm2HtsfqqsAYlSpfP/0eFbehk2QY7jf/sPfZb/8/zElSJ
CsDCxsDygGmzV7yUxnrFc80fGmgszmTNgkJgFWT6UJB8oUChZrLqVGkmXzQ/
0q1RzxujTAmIMYe55vngqPmiXPQSaE2G8ov35d/Qj1MNTy9KmC9VZVzcJcXu
pFOqv/aOQvE0nmNZwZ8uHA5bKpZnAwEGja0M5+q0e4BINhkNNsZ1wFvld1B2
bzbz8cL5a5zXaWuUQEdi/1ioFGDfWtrFeNsSyUnpFf2hRYGTCVHoWUMbGfvg
3igLuRkkq4BsSPw7q3oHl3we+IAmWZyhq/5fwVSyHNt/zTQrcdIUsNVHyyKD
Y5i9TUFn4POafwpY8R53sDDDQ6iojuentRhbaoEJGYIq3pVMAr9mHhVjg0FA
rmVXpwzoN8L1oe5nqHamnJBuPgbXmF1knMc3l0WmAJXV6GAWoZSXHYl1q8pY
2b/4PxJ4fGfzy49OXcWxw4eQfFBsaHfmWcOqvmRLKIDDsCJsmwcgAYD1VTPK
ASvHopuh2E+83Z0IPLglM8b9j8FooEUI29/TzjQir6Zi7ahX0lCCspS5oBFS
VSvovbPveqwYqGyEtapO7RIMZbYXh/X+5PygFHEWfYLbkd3VqUt12xcxpTqy
V3E/XsJbBO/Qk3AGzN4OP/eWfFllh26sslcxg2hUzHrCL608EQ06/BdQejCT
mPb+AXed9wNJJiN/Ps+9/jMj6vlD0hQy+7AqNwmmFSBMLxkSAZoKUSsxV6sW
0f6t3HNlEjS3ZnBuI8qcoGV5w/r4clxyjwbI8z1r2QfgwEKoA7p73i8OVund
1pnfcUng2hrRne58omgZYAgmfTAFu5Qt8uq+HDOR34yBUbEuYqCymJQYmaUB
MsdXtNBIV/HZ4tZH6yI/pNvTjRaFW5RqKDLOeurqhTebdOJKCDFqZI6/w7WZ
5a1uTslbdrelj585ULgV9Ap1fxESPRSmNobbhxoqPJrfMHIV0Oy8rws5z8HN
uNIKkF/VsfP6tkVerGfUXompRVNrNnhxw1zVaEy28r2ckGoqCY4B1tHVqdyu
Gwol4Ekjdn+vIHegXfbXfrBLLtABOD0dkiGp1zReVHriPtP8EsvFlTbrMV7z
vmpM5TRYODO/T1uZWQzG0FOoTNuoPWW7xRJBTIjQI9Rg40A+Tflbm/zZu0Zc
O0LlrY7YWayOw6qg0QOuhr3NIg52/WxXJtr4GAwzkgdTUMTK0AI2j4YTcdWW
wey6h1qBhAswDYwbUKt4R1cNtRms9lnj9SD1aTMnRkLTpS5QN5LUOlNA4fTl
v4MWulSdxvF6LZ8oy3Sd0CvivW52TjzzUszKrfooPbcSIj+7JHMRFwiJmWhr
sayPbM2iYUZa8XfTvv03ihi3mPYIV7JEwUxbRwV16gDL/ga9PqQ1l+26alST
rsCGCPFpIM0mvm6k7MsP+zI2ctsQt24qanYpNWVrpKrL8/o9f46PhIjurXMb
gcSsWxDulGjLujbtCAVA3qNeVUBkVg3kjnwuouacYtI/Y8f670nwVwZhj4xD
9+TSryqzug73nL76BJNXTFc1ClCtdZj7q4GVgaTvzbIc1b/lfdqOAv1LSDqB
cV/jHh3d2smv7svuYERZQ0v4qc0WatsyQ2g5/jV0Az7nK94bxRDRGQ4nDR11
tFUrjW5FV7KP49kMlXUeGnXbIvNLQnRNY04D0hMt1dCNFCHsV+LhzPlhJgib
ySkx3Y/fghTL0I/cck8t2Gddcf5C7m/X3Cxo/1m+PDRcnmKjw0bqqJXpjlyg
JtrQ/m9JDqo+JtiNhDTG9y+2iq546iZzC8UquzsMpQPdoeZsy6VJXi6R+V5Z
GznSU78BY7BCg0ew2L8NxDsKJaTNWu17dLdkyxSb3A0GUImk6iby8uPkIClb
9a6FAWZY5x/l09CfNjofrfgnmCe19lh0WqLi2ivC3etosUPU1XTNmX9a4Pc9
qvL5oC4egiA/VescYXwUwJO96+cLYg5fDOLhGAkwQYtdNC5m/++fh2fA0oHS
4K4hSeBS6XYYVgPym5Q9X87hyfNXpu4MLU7EGqYnFWYrjwdkoSPFkAw8kU9g
TVRCWuLa1iAHOHRoV0BbdfpiUdlix/kG7vVTyEo4szR49+NIdP2N7Pf8E70w
e4k53gkV44Zqp0ecma6ghmAaju/t09EYKj1dcWwOME8dNc3hrX6Zf7HJP3GU
bsm6DtT8RisQ9cBT4GA8hRELZByHLRAcG+gGNXQ8CUk7pmr2wU2xcAV4gJCK
DOTfUtjCJjDH7LcUbMdXdJR6vwWxM5+gJvrqx//ax1Re6wkXu2O0BqDSLqbq
8EeZ3EcPJVZE+39j6fatqYv4Iut4RNnOJc8iu6ifBz70RLcZnW82RWW9Zrs/
p2boG7hK9fZbsCP4XEGRY6mYwU0ik4WpjASf2Fqpu6B0Eug5UKmXemSmzzwN
mcUvZJu6wPsrKaZrP/kuu1nON0HKYK9Aq4wyWzdRcmYdyAP4spJiTMp63E1N
vgFhfNHpZLx3YcQkL+Ey+tlbuv9N2N/i9cK1ZLTkzPyu/ns3F41d21mFKWh4
bIcsukTZUU5MXu4wirVgnM/VNu7La2fXafBA+kmLvk836nqJyTa0cJg2wMfz
d160pAf6udlr2juJZx7bZ7EruZQN0PR/jnM0CH4nJiVzbwxiPRYLt0ktGQyg
1n7OvCufP5wlpHFeQiczz7/ihBx+hYoNhMWSyONSiu7Z0xIaYSJ8gnM0xNGm
J+JiXLhCbC5R5CHbFW+1T5Art/4aum8RCw69tGBGhaKN9F1dXRqNGCD6CCIX
c+3GO2NFrtqnlYEPvI/RZdTw0ywpvcrHuOKJES7qJRQaTe2dyRTFxjXxL3AY
HCm3DF2X/YGuvFzngAaoJooneyQ2mq7jioS+sL1cRIRYZEaRb6ULKmD+3sWM
PUwl25JA9lSnAS2n1MrGHWa6RHaQzvQ8obxtaU2Xv+yRLAdKUbjQthYb2Cn1
tQ0a+LletPSNswhAyrmIaHSUAJijDiYsBoSwCgy8u+txob2mu8MWc5NXs6/7
MHCIE/WVwfha5BrF0FDKsLXw4LvYqGGsxGv+/l7RF/3BicHbn1sUidG6nSKL
P8/qZcn+sQO7ei5EAkHcwAMhasGA2j0p0Vc4p+uW4wNjzrHA02yANR78bC+J
fzZfIqODtr2TYNAIGQI7zshdGt9bE/ABQiIw4uoojdBxRtqonPc3mSpEgW4m
qGz92/sc2xjW8BtXXnXqwl2vP3sHB9mP5woD1wSklC/8BBJZHO2QM4K239kM
Np0NY+iO7u6DvFMUIxHoIlwlXLLeZrwkEvGuL3NTJE5w0YRQHV7GxJhNgJk9
gNQ/lxUtD4bo7+tfJnhMhVTP7lk4YHten2oRdGYL3LcNyikxE7bXwSA7txI4
9b4xq6g8S6GBddRLsmYeiSKXLWbqquIaqdtoqT9MVBTkOLTMbs2OnQG3Ddq/
gqLYKBzHiP89NoLxts598lykCjFvf93QuUJPIwgYxWFB3wIONxiy2nE0MBrJ
QPGz4EItgVH4AXARZFc/2qBNRTTH5oyniBGb+GneO53QGXjQUU1CkihNd+gb
w+X+xAqLumzwTza/aquRIEprMuu12jWCjUCdnNJxNBiEr6nYJ/Xne4uZz2JY
QN6SnqvDAyrt3lDpRgPO2tK4VATbyZQIplkOJOmb8GOOke3CxUfc0OQu2336
NlcWTLn/xFz7HLpcGCfc9V1NjSnPvX2GJUVm8+PV2RUOeNbSa7qWckEw8inj
8rVNDqwqciCFi2E7oMUcil4yfm/vzC4xf0BMKb+Z9K3/3v4bplvhF4L8adAF
IdcqYYGhpfbUkND3uMiOsHNISBxTL+E86IhjXjc7gACujOdjdrbQhqNlDDFr
uzWpNZks55iEfzowKSwFvoSeOAtWD9e0SNxvaFalBKAJWLZgcxzAYSZDH3eg
ViRB6EkbCqv5IzjbEF5N1G+P54ZEl1P+Sco2J87N6+66ZmFrzvLCktwXmkz+
Cc97947Ce6AzCU0/AUgiyEhFoWQlGKWNVgwHlkCCJOdzbOd7ewRiyvg0UZdj
NU2imrfNRlS4QaeyoISAmFqjUNxR+8kDLsrHdDmhIGDHkoddC7jlXAqwERC+
ekPwctlW5GV8q/88xLKeWa3KaOuHn9whzINwrSwJ2iKEisTsVGOSrzFWxPPn
icnhi3RjF3M533g4JFvz+vcV7E7jQIEseUqmBhvSDGHweKxan+7wVEZCGY35
uGDf3AZBpsLBmUYis8AIp3jFiws0kitS9i/EzvnTyaUhEZkA6ubNObRjtwAS
NugXYYO38Q5+7Xpi6QyvXKEq1/jrjnXXpXc7JgCbFUdIHDnsHTPcBh8f4HnX
SMDKusoZF5w+ePtqdMhHX0EGqQw3vMTKHtsYiIknZ8OrrMw8hAspt1oG9dXe
wBs+mJRNbxoxUTFhoqt0pjgrNBPu+KNbqHwSNTqU4PPfk7gEzSuRlhp7W7hx
3OH24BAIorC6j0n4MXlHgSDWhYw1Dkn29cJ4P0D+HoT4YBvY6GKIiwigEL5O
yVd8db2m5DrHd3h3bECpCef6BwiTjGFZhH1rA7eXft/ujD9J2KDLmyge7tMO
F+gGWGXPnj3U0sPbnuJBeqPtWV77jns8tM/vtL01NMJIuRg27PbUh4sGKIAN
0k9bNVO6cTsr+mWf+Y9+ZE7/F+jPF/KIq66hIy3YmyZeauZfpThbbuFtuvSf
4EU3ElOpBPR4z5CHM/AeAsomxPd0ohKtobULA1uRmXh/kpJ/iE9uYs0at7vS
1acxyTAWbj4Nt9xZ6+vPOg1rH10bgfXdVrFPPbcl4Eq6W9cWwkw6PGOwbJu9
zH70bNjyE0jtvd4trYWADiLK20LrZmAlyjI0BPbi5TTP7YcnJ3c2MbKVLQsO
xE61swzX/GCC+7EAsB426g1ZbNs19H7Dmh1u9+QLk9PMxTiSBUjbdONnAYeh
yNYfWcijPfvdnjRETn5C9iWSYHLc2dgua+6ehrG/76wmV6f/IZWszFA4rvtY
zbyN/KWaUvzpXyNfT1NcsRfmVtp2mznek3h9OVJIHDNuY84dq37pbn1ZQDf9
k0T8IafCH+ASB1LEQkMbtDMqFLNRSlJ2sddnv3bXl8cnJZ2VPJmLYPdpCaOX
LXtT8TohR2o/KPU0oX+5DjXum4oA+ktvXUhXRKqF5YnRUtFDX1PPaqypzb/z
Ebbqa5hwBmewmXtf08JDJtc/bVturW2Tz0HNb5oveO2HO3sI3/mBCWzeKmQN
Bm377UFEiu/zHIzXqp2kGz0SaRl+cL8maIlK1dCvv8SdcXl42Fji3RR18DcS
sjnWyHKPVOBWNrhU37RbMa+4pU3/MqzEsiG1U/6tdhgqTjl2gwV3Ogi7BD4+
rJYN6vfqUkliCr+HHrb2ao8bcpLTA7pk9N9I1aAqoMm68vESCwBstzSu5Ex6
KusnNxrjV8695DXK34d3kwRl12njsEuB7KRF+SmN8xJVq1xjXS7p2Cvhka9v
kdzkDW+wO+yQgEp10tgn9nWIhsHzDx+lTbebFiRqkSTxqQWBrzw3aFeEkl9n
kIT4pCSGpHX+KLWrcrx6GVG0tErCwAUD2Gr2fZW0F5IvP9PHqZ60TzdZYTtl
A/M3W56WlI2rDQijH41SVLhqG0xqvjM+TTPGAm0Tn+DQQCYljlgVaDWfbUqy
Ms1ZigHLzHoFTfivu+cxvEfR6zBcn+pcK8IUWCoUFwBMezDH9YoOmgsoAz5g
gzre/dgQ9Ex1dWE8BeNvSh0ceV/VjkE4tv3o75pbM984BfMacEI0PedfrOdt
nMUQhqzEazshcAFwpF5NtIb49QzCvT+q2w5E/vG5icJt4Q/tWzE7mT+4yYQy
5oSi2PBfvcQC+z9T4vhnUQM8y1TFIpymC6nlDBgMiWIQEcSEgwT2SMBLUMMv
Gf55WDljtaRhr12ojmTM6+9h5EG3rIWXqAs87grEOvoYyKgk4Px6LW955MUW
4Hr1UDBzkZy4xWRKNaITIQ5C+SrbEfQa1Ab8ol9EV1nwjeH+eaEfaiHaQU93
q6rWuA50B7F64xLjIPzTT5JivDYs1lozgmQwyemsb2WDeaDISIgBGnONpCv4
7QqfcZfFd7qG56Jl97lOwE+O2Jo7JTe5lsuxTOXN7FM405U3nRwjQhTFP/OX
WALm5UAZqwMftNAwwt3B8wcRT17JULBdQvz1Qdyh9/BX6no61o/A8uqq+heo
mw3iIfc03hoRrVRU1uXlmYGhGUJ+G1YThDI6Xw0VNKYsrl6ikrMwQS5jmZOj
KfXWGc2KTpMBlj5DxdiupdFWe6KO18dIqSwzZ8CmpBNRp8R7/WoNpj13PGNX
nU6irX+vUKsllGogXJXQ8WB2uPcaGN0fk8yMkUeofHsKQBeckt3zdQetG3JC
/XI0njpAedeUYmdAzhHvWVz6nSRSslmJOQfVorRidU7GN0MHYhAojoTKNLwF
8BBxpXunrXdqPGCFsM07+EwTzfPbR6tRHUuRNU5PCwglGnSMzRHhE6KLCcjd
GzPQRS9NAmAXjrhX7GBO4rhvCKqQtbP4vAo8zBRN+xnQsTlXaXUpIrg4lc8D
X+7WAy/Re0gjhyv0w3Z4eOkEPdeYTCblJ005ckd/wXMZ4gtkwKORGgQPnyhI
7fCTR9owp8AIso5VG64eAT+wboNidCgj2BD1tKvy9NibtJovvnuhWpRClW9U
q5elkwuqUGMFLKBXG8YDbRF5144TpQShnzcFgUL7ynV6WxO3yaoDbipTx86o
YdJI9Eijf+xDR+YsamVFlLJ5XconTN0CP1+9Z9EV3wZwq6YGJn1zhmAGDPZA
r3w7AWow4T3tEnpyRITxLuQOqyjOW7L9NK5RxLwxKMTpmB2KtIH3HS6EfIy8
OcQ4+zSX4TVIJIhXMOEARJPTjjYKuj++GbNGqbqdQb4N9uJ6iwO84wBS/006
pi9UdGimzVEcgYmrAoOX/9E6JVjuvzhaeaqo7Q0jRy5UVUo7MBTmeArDeCLk
mpNwkUi+BeyIi13y9kofuT4/5hXsnZQxrH5o77CoCVzpD9kIDF/X6roPFdC5
rYN9n/qFJlSr0v833Po4N7xhykszXhjxD+wsH3dlJv/QNscdleXo2YCyaDra
56UQ/JiatYqav+Tcoxjse+tO01txIkSVg5bnpqJNpF2I3G/GprDS9BvQPE7a
q+ZLfXjVzSejo3ccpXFsD28cTiBTnpHtLpB1rv+wGmaOYU7vPCsLfjM0aJgv
bwQXBFh37JGdPqxoqKOUfNa8ULjMJ7UKIS3SXqb43bHxIfJxVRX9MB/4v9Ze
uiFnw7/ftgAm0/m6LMNKupWDFdTfnp2EI1QeGw3/QOu5jiTX6N03D4FtL1ts
FsnqyeJHb5H/VpTGInRo4o9GUFoS+DpuFIbJ8cYNeDBgqM7ws2evcpo3qrKs
3aRbwasQ6KsVyzGKnZ1QX6oPhOWu1qf4bBmRrZUT7lncVO+0qOl93+JVgp0E
h0ghdAudS+89F7jtMUnWySsLW+CZBwowIqewJHrod98vGMBueHeZRvp+9JBs
OTZ7T66dR9G84eOoeM7BNj/yUt6ou0TOghah2jYXEOlKPa5fkgaIebMfkwX+
1rfapPKVN3LHipmec781bqntrWNPE/+KrQZWMTnvMJ5umCG2sOvU9VnOsxnD
bbd5Z6+EgzFbvPBHkrl4WxSxQB8CQr1iDKNv43YoRkNMtfWxTojDLsxZb6r3
rwd5YoP8tM3q3l4DvBL2Lgzwn6jmjb4V3T4bk4vcz/vnOUeYw3CcwyJMtqLU
W4sTYvAd74gh5Ikmp5H1H5Gx8POI46IDgQ6dFqUfLRUcGHuqE1k9+Rvy93pV
jfW5u1fVlXdUGtKmi2TcCY3dNzs2nubdzD0O2I9R8tiQAD6DIlXhiqrg1pEQ
h1EYenpS4IeMy8/HhsQP1EvO3b/vwJ9NE1ahztVw8xM1+SirXQ1+nN9SyCbq
P3sFnt5uCSqO6WEDez687lcYUAsIILmgFS/hH8Vlt8a8Z5DNBJThhxZxP7ST
SrM+2mKDbCWNTQatvnhhOWBpv3xvI5R0ZsQ8LTAmvn2WzKA1DddU/PURJ0t7
dgoGvkcpeVNDwRVkJh35sHTxOMpvCK7abnwsETSngoqgcyekobd7qFggkYfS
BXWEOTMUTij+YMD6Nel7oy0YkZQPyv6UccbFNcdAvGj1Qf3MjoEsA4NbdFpS
n1lQPWdRSJSUhDI6yGG26AqKXSYG9P5W7H0nxKF7xNqPfL9JPlJOk7vpiGbY
8k15vntk8pK1uoEbybOJUEv4RC1wJd7n6KLbzDgg7l2HQblEtlPRVPsxfbLK
7snuPe6VwxwqR1+JXStM+MHStCkOnt/2312uAbH/ik+rAwFUexexYa3Vjj26
tS4M9DXaQ/UzGOlobNhVa40LaRDNiBIGD3t6iwdIiiuGKt7zAmk7JIVroFHw
NTcDVvP/+02RCTDcJ9FqOH7IvuHNXx53lTAhkw0eNDdE0xF2dSCDVhdpBG2g
U66CfDW3eukTRMg5T8AhangZlkKYTQjaMH/SNQk3xi5mwwKasWjlUhQ5j1kf
ATqqy/MqjqmmF/qKwIrLYW0y1epPRVWdErI6vtmw5bbZbZn5vhjZ56/dssbx
nrRhnrOgNU0aDCm/8gZ8m1P50wTB01G52n5conRaCc3XBCkqao3OA/ORKyg7
+xUEOu/uZsF7xwzkXcwRvqBd0B98qhl1INNpY57ayuTLwBPNY9CuYblH1wQC
Dde9XE9qu7qeEgHA00M71UnS1JFaI46hCPIMbRwJ1YQ1hHnGHplWKOyn9d/Z
ep8XgwjXcrP8ggsjfAUbMZm+qgt1ah6+l2RQrcBIg1P4tTH11Eu8z4FW0Kj/
0QoIr4++bEzDw0thRYVX1yH1UgT1PUurDPhoqE73DfN0WUUdgs4M4O9Hd0Tb
XBjTGlIFV0UhiojGPHzoocjAOrMbox7rgihahibRv/etEmxq+xBWjX/ZVdke
F7H4VHaOztJ+mA2MNVhVFnKtZCdE/XfKDEp946KyaeFGwwELlaJP9DOd977z
i2Yc48sLoR5zg+FKCKUUTKXtzCbU6eztfoEqMCg4C6DYvfnjhdFGVoY3jVSw
9fYCL09S7f7A1+ggYU7PyQfjSpCHl2NbSP7mWjhmYb2qXtGssbzGiFd2AWjH
YMZzjS5e55of4qPjNV/FalWPjStPwAAKs9YBfe04t3z3suWrOTcaWHtYxHU+
5zdlVODUk1lTm3A9wO8x/+SQ3/WL1KGrRpito3M8RsZSVhTWA/u2TZ6Z93d3
GvPgYdp7fw4EFfDG2yLwZuAFVsCy95rATBt6KUoYeeQjATqS/6DftQLiDc9W
bsByodcosGU01Mdrt2WsnlFrBxo7SkEcU4J2LEFU0d6VVytsql+onBIJ3GZO
t2sfVwiXfRFsobmKN6+BUHf3TnVyuyYSnwno0y90jlMvj1lT9yfE4GvgaDsf
HKVY+LLt33sE3YyYQzmP4az8TPlotzlqtvaxSf0MPu5qmIu63gIarvCszsu4
QFJt62P9LAn4Ads0IO2+DpzMHFa9Xddx+ASfdKPrUgRUxD+s1DZrG0VJtDsA
oPnCsWrNaSHeXgQOVJdVz1isgbbmX+k7NKMvUwqUqIEIVO8TQ4Kk8TRFZAkZ
ubpKKe0aUbFaMRI5FY8+JlRXooYaTTrskLHcEV2HK1V+4ITrKeItMsAl8qlR
y/SfRe8pjb20dXiD6U0mjq2FwZ2Jifgkr/gszg1kxX1amz1GniPLSsModBkK
+EuiiHQHMVe+sYFqWZs0Z/CtE7XKhAaFNkfrEZN1gVfezXnn3D+sSU3//tWk
O7/eA/602Fj4wlTWnwiZ/DEnx9DAJhoVUTWgvPTP0AakH3TXGd/lG/7M8EN+
xJIZqOXXTX3mcaPV4z3FjAUAn22Rjs/F4/xfL7pTqJmef6D809AoavYavj2n
iSma2rEOPBC7oil9ckxs58Jplq2vCMaXH48bOLiJZmywk/fNf6nXXQHUCCe/
M6OD2lbflrxVyLewykAFsFGdRdhgUQ8IIXFrgGs72v3tzWEKVxphS384LDfc
Daqfylfrl0RzTgTxn/hSJORkPy0CzejZ/+gy6PHjrrBPFRoaTGuF3RfHsrVb
AgQNg535SzhyjV5UZ4Ezknk6uotmWjlGxJqXv5vwKYuzLKRLyyJAe4BkrMFc
aalGhWZEE4IMakmEOvjc7+lJeKIZdwrY8HFVLMTP9kE5tEJpsjsZIADOSGIP
Z+3oWWXSepJ/IOhx90+x6QD7kASkUViEtiKQLvzhA2t3x3cBB53gRlY5k3Oj
Fvf/qOAygCNMCQeu7GoxnQgesEfzrm/LPuBKkG+4WlBsXUj9p1TVjmBmtV49
eeEDADaTVgBlRy/uNm4VCL8Z2s9NlsdgbHg4NBEOPgb85HCky7kPwqb7rb1F
sCz9Zmvok9F6cPBxS+cthflLQB8iDM/PURJW5pyfs/8S5hFjgLp3JY1XyZu8
qm8mnBvx2ICzsUQTdnzyvKA872b/Ai2cWLIKw5320ueEk8nfmVRTS1QkVpYF
h8nnIEr2tZK9zju6uzxUU32u6+QqKvtO8x/+2I5TX3IbkNPgzAt9lbDNZbZZ
73YfNXplLOxBfB63nLC1DW481tRGn7SYaoGBaI0cvuynCmeZMyKssMxFE5Bf
Yf2UkEtZPWLbq3vVq2QzmEEOEJFQbD4BwCa9WzSyen1nAj+BdziLFaZzSGVr
zBFBuEzG69KWIuzUEFogQLAA3NCST+Qe/I5265+WYdBNVSpW9ODiSv1lzjHZ
fhGQ7LVWibcsJjnJFvjg5UAxhGiIGIaKjaZGKhko48b8DTJEewPGCCPCJRmU
AWc5i0YazObBsd+iPtVH+LTtzXDPVjG4QkkR+7IhWu1dliOXRtb5QhpyXPao
R1Ac3pxQ9qlaezFGV5L0N0OrAw8ClGwCkKkSWXU9K492kzLPTyUwFuRpHdJU
QwZofMJpnGt1k+y5Qg06aUQds6cDBCGHeZhs1RPDzYn72gm9ph+hxo54iLyv
bIiMfjUmaYorSbNe52b0InOmHDz+9dSjUmAcZ7sU/6/G8biIhTzJsslkfxh6
ncIj4Vq1swHD7v7LZRsTcT+nQsrcLxdkGSLXypPeF8NrtIkHScrvDzpkB+Hp
82VThUKDKEiBBxUuqv1YLDkDf1ITo4FAaxqU/qBQBuKj6gSR787brmanZEEx
NO3uodCtIdCfeVDI3Vtb+us0dZADxSk9kina0BRLUlVisMCDIv6YpPRdQTBf
YX2QqR4L4pMV4cjbukPx0SpBDa6eje7u2+/Ds7F/6CEclnOqzw5pN7DiWIHz
HaUxACcJu4GFXijpwwqNgHe2QDIPZRpg+BlNRbd3jGzyTAYz+TULkYduuX2Q
WhVgHXRBrgnYVOActfrpTv7kF3acIjUqpnrfaPGkL7OImfku++/IF/Vg8C4s
hivI613dmTZLbCI1nthAoZgZdH1XDhRmV/X/lugaMvfXU/LDAG2ScVYsoGId
XPLC9q3S18rRMG07B1sR7cwk5J61jFqYv8j3vhUDzYMnKrgW7epJLeduB4Bg
UuhTTJqmBPem3loEDffxCXuN9lYs/jdnhGeQcNiShX9wVkWkUmrPRgKTI6ai
CchSXZumiabHzFmwHsLgDCDG6fRyRXdgTjonRdBditH5kMP7rpStU2S34fOs
G8JJUWj9HA8dVsitvfUyzYlC9Vppt7vV/ACVzPlIaPUnGJQenQ5xtUAAWgLq
I8DlOQH4nJ0cYcAqxMcCCqWDyPFP5+4f7MVhDUwULx2p1teaGlLH1VnrJYDP
KzXDf/LyQWqTp0J9KpqIwDZi7FG4F9gKtz54ElvQmDEDVfYcNSSP9VdtziXu
b2QwtuVEegU/dTOwmagWI5SO/YvbdikpI+qIOtYSVnfBmhPtSFQcJy1zkE9v
nu66cZwfjRnoICe0br4MbgyIZj0amt90+FyThzWYz8qIiNCHYdlj4t18xu2X
1zCfKz1URY/ZlI3LsteRlMyFxo0TX57zJF3il0pf70+XIEq+mBahlKqSSP/o
rjZHh+5NDnvcXGkvFg1g9cVDhxVSF60RJxmpfJQUyz6XOWOcvKfcIvKC2y24
D14BV46kYzVMzthbVuC675tZ23FzXsfmkH9hzq/7HpBXEbyWUNn/4P98ze8T
xdW+YLuzRrKBebCS+xb08AcDbA0O8z20uwAX0r1J2bnJvsNDF1vGOJKTPCnm
3wMeoZCxkkoy5PkBo6PEs15ZbmmOegblaG1+f3H/yeqFHYzfuouaAScOKDjT
xkATIZh2/PaKuGYNf/B5S2ztRMaQmkXbxQttfMudMXmchBmMG/bneiHtmiRO
RXOdwhUGDT3uSgCmQzgyrCIKVEuERL+Q6MCCTyNrOcPvZDuQ1AODZzvPYHRw
yJchElNEgTegiak0ZUTppY5y9ZGPY2nr6P1C0+k0E7JrvjapInL1nxfZBEwQ
Ycunwjhv3x+DUK+KYZs4mdGmfcJiyhn1PTHmgZXgjlhRXS3dp2u9RCOkENJt
1m/18SyVDNRzeKndo+m2pPt/x8aNWQvMqRcO/uK6akMmHc4P15K8zLS1flBt
P4MBoUOgKcv+hC5RYmlvKbPP9HpErEN4Dh2/UVp5xt8lFgRdwXu60Dn7OZwe
Hj/3om/M6OfXqTZb43ApvbvAbWjeMiYlSE79fNwN6aFoB+URcugnxy/OpkxM
92MuDE6l7gt7cJ/aLXkVX6aIBdsShoMPvoqV5X9QjhacS1OgMJiOgiSutDCh
qPFMsYPq58J4IZEPv0mhcca+ZTBjMZ6JclL1l+lPU3WRj//+q2+TQlB82LrI
47xbTBAkl+BT4GdUIqjHOupWDtaRgx0DpM/Pd9JtS3lwIO7iJOWzzQvW1kbA
Dv4596f8T5W/l33WGRV1OfBFyHdv9rtrCem4bF7TbWzLD36RSWxA8aL4Phil
EFFw/NpMpWxJuzs3LHQ7trZpZer9RIK+e/qO0e49NiK87r1BapyRJpOvy0M9
26Fwwytrei2na3lDslOB+pr/npOr8Z4Z3GsNRehVtuqA/k5zEAv9k0tnKXCP
TAsx+Cb2PFMYqNvrFa+X1vctns1NvvQq7z4/HyS82evC5HIgnsRuCvq30RDF
1lHk1L0E2f/2lW84roseBpJZqrJwHwRhAfyqqvsDg18+4+lgTIhmkdawgJK/
riC+1DsCtCfoaCmdv/iuMzUq6D7E2RYGx/cWKOeooJMsJy0d5ip8ZXZzqeEQ
dxEMJLP3resqgVYWxPrKU14RZftdvgMkcXrMA+pVKdsfpoUGie3FNZH9BdT7
QRP3YJ4UDL4kI3Gzm+pWwfQyAuGKEpEOHtCJ/k+t5RzexzTSVNk0QX04fmRP
ehBp1U2SACqdchqkRItF7bL6au+4yJzwOWWB0oFDDQV4TKjyDcx+d2KPaSx7
9x/j39oIMHTT1mtKYuQQMwV0vgtb8KQqjQxnQnztpCFXw2TNYNWBp9zCWWaa
vOQUbmOOMwc7V2uBq3sEcQhLF8zXmQgGvT4sDDuJFLbwRVYk7DZHj9A9vMdX
1h3zqPwoxF3eX5LVPkqFFxmaIZcqx6m5nEUYZAONE1KaVXw2Aq1Oz/rT++zn
IumQcRWTTJllPuq7CETaXGRFusYbiWo4qXRsbhCTnOit4pyegIaqCmFqCobv
EWwoYAY5swKnx0D54zUPHvTOS+I9DvSybW7hjExI0/qivYgUFBY3DEiEpq+2
G39k1/TorQEZddspGCAXYc5T4T/UPJCF7El/mxxwCSOP2/59LFX1U4sT+q5Y
kTPaCWrxjY50VW0P3vePLqo+DH2d6Z3Bfy1KrlWa5LuOPoSoIB+llYvjROL0
c6t9cTQ+nKczNy2onkMe6GTTQH67+LtOj7+ey8tsEQ0EW2FWBKctGGyMz7hV
3wMNd+46ZVQ4McjJTYIk5fd2Bmr2EwSNndzcKin/aKS5hrByonwny31YtQCa
Xr24eytfIMdIZvhqSHoBRKpgEPmZpVP11gyYbyPiKNCTLoTxanVkyH1zq5n/
LrHlv/lZUWOjpXpGnA1ApdY8oiuP0VaSZIIbJOZ29amA0jEVeud2ccqkGJL5
LQlCrntMfJJD3lA48LW8HE5aKXZopRlkpwBgRMMmidttczH7EIVCQbxARgQW
c6I1gypXygPOQ3k59p1alV0K9d9dicQgwP/5r5PhL2LlaldnhUiFsmxjrYH/
+u0K/d9ajZQQ7GLbtle4JwlAreUZMsEveJSUegNiUAep7esAp2i5Wzc6t+gd
ZH5S3rxyVsB6VcSXIjq85BatH7Rb+69J3qGHCdrjAQ5JJw/1rpLE+rEEC4wX
FBVoPRK8qmZtur6Py6b8zbXUqmh+GFXtHfnk4pCMhgED4SqMaPYfARQZAAvV
QCerzRxtbDqaPrBcqVuJ/7W+W7bwyGIfmUT1zbFea8kOM317lvWRq3Goitif
cOu9VYHid2+bFUmc6eLfnbzVTFIUZXoacZ0wyFdUk7+97+vNG2/WuFOtrzmQ
me/P4gwgo2j8u0ZKGvOau6W2maZvfP6h4p9eekN28oWmFcbWEI0SNJOE0w7w
+lqhFAW6bsUbvpSqTPkE82X7AWW6mw+lw1FGsfl4pDZoP6/SeE8XgsOvG9pr
orvQ+FthkXuOaMLNzLdhyOcsf9LoyfIW/CuVFDxb9t3KJqD5yJsyN82WTu86
2FYYuKY5/xQa+xvlsuQKnWwQ1mPs7r1UNXJmMSTf4xx/fl6Al1DX+pbXb6ur
r0a7eavFi/Umz6259W/BlyC7g6o0VPHnEzAof0oDeqiMqRGvdHBxrPCsIVcL
kx64lceVgw+CD6WNxSagssf2JUIBBJ841tsJUuwd5iX4fdKM28DF10e79KNm
+Hr1pu3xS3VbgijMMPxv4z7ddNI8eu8hC/Xtnba5H1kA7QppgeLw6Z+LcsAi
PmK2RFSuWv9VPX8x+Gu87GO97dTZSECUmMurJPvx1WRvAghfMCNOLpdafTX3
Q9Gdouqwzezx1QroRaSAMSBYZzwTfLM7kAkW6IvsjLQUJztukNCVaAUl8FgT
bN31b7td0YfdjAwnGxUrnoKrYVhOvL/web0E2eDoIwNE8tKFHdlafMESHuZg
EcxuprGG1Y0Dk2Yav3p1Tif16UpmSDUYrrjNWdUaAF+atjjXXhUJpbAgXJib
JpZe6PmJl6r2nPUSp17F9V/Yfvtp4qa+lRTyGZ914zMBgmG8PBeRnm/5uo8x
QpAk0wekErvXzVC2UQhJd1zysDiBLFTWUu5tRFMeKlmuELUp69jfo+PlD9Qt
+LSP0O3gZW0/0Xd2AV1pojVmbUGJSCq1BYuxjHHoI17qvWuXI/w/LhNAjTMs
CzdebwTYBcfOCZeVtjFcFawDU5B5HGcng2sH00Tbzoe3LU+YgGzw1VVnpWyX
/TXcEXk+Lpt39K9mdhzYQ9xTgk5KRekrRhHvEfH+uvylt2iHtHx0RGT9jnrZ
Cb3cz/xJEqXrbmwA+6lI1Zz3ExbLSRpcUp8+cyjtD1g+EKdNThE9akmERDqQ
VeQr2nEwwPJDaNDjMO8JXJ5lsy5HxPkitiwdxYjA6swgiTH2927BlOORWJ7W
rKvH1BNd198Yx3zK+Sh4PDe5NrIKUd+FNeAvUZvZ0OxvgIX9clwQ14VvDloN
zW9XXxrs7elxomFfNGzgQu4nYE9YWj4cJ/ruK1FyPREpddx5tyzNIjPfhTN+
AtfEJcAziIo9NuuZr+DkzKg6sNxp48ewwLtfGj+eoAdZDLrxXF/JJia+WS0o
XE4wRC3uc6E2hB88HI9C76X4IchLtbHGA3hxl/DWUt/QSI9yH6bVfvWfvIs0
Ye96GWWZ2of3BM/3jAduR1kLtOIk0CCgf3htzG3hRes5/dOV4h6SwmQjUAfn
VMEbUJlHbVgeyMzqs/5CyGgsHxEVDfUYk+XMok/n1sqkx5KYxtYgdoLmx3ma
zopmQcrOBngN46UVnrXG88OKE7k3F2j2rdLvClUyMHdGuvxlnrbMu3PdyqPz
btjPLSabY/puShPB6v8xUXvm/w3VtyRaXSJkV509TK59D8jYGWhDK8IFdffR
rTYcgiv+Hf+kLiYpwyEbTy7m8kAFHuRQ8xwmjOlgxqIz/fUaQaXOAB0Xbr4Y
bqgOlS7lfeHOt/YE78EeiFeA6nRuQvq3X2bmzh4mCG3WbuSI+kUXnvnjoIeh
MnFXFZLpFRmXNmBoHXgEALkWpW141/nTy4LZlTU1Na1ik/9lRTwozQeUTyKG
fRcAKPWwQ7Wjin2Es7QZqcbP/StrluZ3rEG0ZJzT+1GrNEacKFXe3NdXeMAh
Y8D2+gs6as3PgW27tXgZeTjgd2VBesLlrMzpPtIm7cKtAAVZQR4+26NdYRu5
nlhxet7ICXh++bUt9rssxU5+Z9R9b9Mg4Ej7Z9Cpbm0h4pTOEBDKFHD1as/3
RDX4C0qruCtjsdZxtHhU1OK5z1/gFoCxP2U+vhkINRLFOu8z+oIPmmDrjum/
GH6zWVrr0bHliRLAyHnvniXkD0D44oj8TMtDobl96qVXtHaBROpgjau9NsHZ
55pGN9Po6Hm+lJeE0CkkxK1/n9bPgHyerxZzVMkjPeLwxmfncHPF0QHTEwEf
hTmk2NXcpajewr9ESsTzD7m/KOZLWwFzWcTlHElsKyMO4YH/XVqNW6Tyrx44
k+gkn+oJ/vmZVvqgoVTaK/K4ikikRNSNz7uY+k7REkMzvwDvopYPHWuSpXcx
+M+t9Sv9Er+8fOykpUS3CJN9P+lOLJrbsZ6wn6yj4/UxZjXTcXvBNAGmSYOJ
NKoUwo/RH0mMtEYd9klp8V5Nnm9fT0zKe/WnzZErpmjDhyutYjZX1NoE+TRw
LmzlSH8rS57qM1E5ILoZGFFyMUZFnAdUgqXJ8LY9hwVNtCsvElHh8eQDto8r
KrbZmdz3e++bwpBxKS7Al0AY/agPe2dFMIvm009zhLFL9y3XI7A0foQPi0bw
uarCT9d0Gj/DTr6tvzbRJ0csQ6700SL7i8g7XluSIPV/1n8HwjFQEZPdB8Vg
lcQIlYFUtajXN5MemS/apC5W4gsoZ+2RlplDUoIUytAUM0CqYIkJCx5VtBk/
P4SiFa1QoSfkGxcsJ4hsXW70DXlKUpOtsoqmaOdUR0g7uHF9JDUIAJanqw3V
afNtJcwFLVQGSqwitPTbNcXwXSryk34DFyXKCl28iS1/q0PbE/ON4WP0U/Wa
28LPt8MW6f0aEKDwpiWm4ij0KYnO+yGJK5KMzFfl1dhI1EICDr+7KsDsIhmU
2Vdw7NmggExBRfMWgf4p1MOlhinN7rMebIdjqmPdNUt+3SWmJbQe3DCuS6to
5UqVo+g8qFuvBWGjvaZdGE2bIywX7HMHa+UOMt6O0rO+1ThwxanJGgHM5B4n
pA2DLDl25plOAEBaGezc0mg9/0QAp4bmmBqR3vg0a3RfftdmJIw9kCGRM7ZD
BrCFRFEOub3Byry1eNpddyrdkQpSwTtlL0ayrFWfjuUhCOCW4ptNuYpt1zqW
toGce8PRMZxgnZOx538CK/IdzwIgl2gEqJEDSm4FkiDSdJoDxMN4IqzAr9qC
Fe8SBx8tnZXubreagErvDdbEo7T5kzjE3e2DjDKTMEoMjjH7SOem5I8zQCTH
ASsaLdzUvVaLPTJSy/rWE6K9cYEYeevhoW7ZXUJqegyF4lv9HQ2tJfh37RHf
HgMCp3OQvh3SyQaYBlwEiSX4s+gQ92JNT4AEinwT1McUQOee3OSjWZs5VWBr
jS0fDBErWbWK0uVJhhrC8J0SqrJdjA8OUs9yB6CDSj2/mGL/fRyWBZQ5FVuI
dn1RJNjBz65AmvvkCPLeuxmnm/NOFuk3I3Nd1lUMj4i7MlqXY6BdZ4ScEFQz
Y/z8K78jw7MKPQ2zv/qyLdEb1OeLFJgc90ioYmlCVH60B9Hh9z1uVqt1gH2H
iILTzmiAJvuO+BMKp2cqDKmC5nLuFil4jNms89RpvyZvj/Q1uYBo2hPI8MnU
iIy7bdN5euYaq4y7KrhzokRCiNxrJIKybyi2HXpJ8c/IGa3beWG0/u/KBogp
9JzRA01VjQywKWlsi6p6Gw5oAxbhobp5ZkmF5aIa0NG3fVoLgy1EOnh50xkw
vTa5f1U9431LR4gpnieiE6wpxbMILffen2ioEAVZSzz/TosyH3IROtopOPL4
PaV3u+7KLMN7HkYIdIepPQmSZLsAFSYRZYSz2IU7Ndrue7PZu5KWEkRGs/Y+
4efCEVj8fg+sla11hiE81tXuAvc1XVSu1TK42kRNSxB/XJqCCbzpt+1JbD+N
fXbE4yvtp8nYnkBzVbR/Oi17QYWb0BboR0zRBtlrbKiYgZXQzgQPfi1zA3I2
jBd1Sg1CY83TtSX4YVihPYsj+pmL8Nr0G/LO+D6CE0VzLNuyezLbSVZb5zl4
4RdB8dt7JwiUJunAnIl2QZ63zX1w0xjxran5EuxJRxF11OPYKyXWOf90eyEs
BEI2C8jMjj30KNY5p5xNlyiaXOJfuYncGa1bCTn/m8pWz2yvSKK3FamWFCLU
yYPzBvGr16LjqTeQsmR2OpF3pKrkeEmbw/kbG60QQ1xIHACMD7WT4QmXgamG
EXGLc/SS1wDXoT8yDL3SXR/dBBHVq4oMMAFvDjo6seI+nuIHY3SPKtxI76WB
Lm+TFrpn33ATm4KP9soQvVzQKPaNM3KiMolafCfWbzrBjmMcwIaDWJ6qkhlg
nUVnBAI/ritIycUxaGzJlSOLKYIAE7bg1GQivdkrWQmOoPL7CZGCOHP5Iy/6
bcruTDQHwPQtTabHnLul4i5ciD+gzDBsVqkDKpzDbyeogwxn78sVbrdVXoWG
O0Lh/8E84JeoBS3ZM53eaLoV7FulNPF0/PwMpNrB1Y/VnDOHpH8dLgFzI7yt
Tr13gJ1DuBurGQk1G6ZF5GjC1QJxsNEdsvhOkeha9jwQOk8o1cMbbXprr3Eo
bGktnvax1Bx4mW05qzPYFTqQ3F4Z2SrDUEtXUoswj2FkH9cfNKYXexHMozb0
dT4LupDJ9kfi+uCnv8e8y2P+cxvJdeKRWs45A7vS9FeNOV85FJwT1SVLaqsr
uFJ2UNxxpc0nsk5TcvEb6FwbjqUzB85RTIgfrKmMPS25oWFjy4DGU4vjal6U
oXfcubBvDEWm10QEqKn6pHftz3epHc2oOoIfdp9q1I6cC6Vme2Q8caj0d6no
0nm6TneENFFPjcikk8DKJl3T0fapc+LuqGiieh6Yuxb5Bd3MI9/IvU3pCiCZ
1q5yKblLaBOmq8Gg9LdNxXhhJhPXwc6s2xIB2iTQhSDbFUP1bCtgOny+lTjY
zTrnmqkzH/9nhnaiJK3WBn7cbynd8D2VwJ3av6JjsFdHml8htciFUmCIWkZL
Ok+3XoNFxFtgo1bi2zhGGC/EJjCmSvPashV4ERArAZr2U0SbBKZES5BUKpsy
2huj2ppJJRAeIOrb5VjcOcFky6zUdAkaJaxzqxfJA+sJJKunhmqYROmPlk8z
GjoCzJyzSkDo5/iY+tew5VQPnelhLyi8RGHq6RMLHqJDajUTVQpbKgfTMRVr
S9cvgmQ91wKyIRx9grZfKgumRRDhWHif0UTfCKynD/uXdpWgGbhsALrE68cs
/jgDJfS9L9YldX+jwEEOXlWb/6JoPvXyqkceKiQbQQ9HLdCmeBD0ld36tfWs
NHyxldcx32SK5/HxxYCQM3daX3JI9qCdNcuqmTEDmpOrl6pco1qwWmdW0Uzd
sWw4HkzE8YPGzXEDrWxGehU6ruKdbeOdcqPLgKpzHAakEVHgOAMUI2a4WrQJ
rCa8osV0q4zWEjM1hY4dHzj4M2XDacLIZKCjKcNX9gbCJP7uAsHVGq8z+XBl
tcEysIfUdhXmJN1BdJ65pre5VmJFIHwcPSetLV8d7HzHJASsbXkcMR8lTl0v
6tKbjSBWnGugyI7m1s6LhByTIa1lDShxQ3C3+bN4RF0NLyjy7zkJOQtjQQ/P
H2seQLDWdIgRbSp55ZAFQ9aahwNf43nQW0G+wbsg8rxaZTmQ2NqO8k3GFvAg
rRRQxOwOHg3LU6vbWtfRqqUkIcg87OknsZohoCi6eaU2Ti/Gnq/55DbKauA8
wBh5Y1CBX8I2NFKplVqAwAnoU1YRqavYOWo8AGgyNWDspQauwgg5aM05j6N3
EgjqEmLfhWYrlp5llTfJRl4fIvTLdP0VfXkcG+61MhBLRcCjs26K999Yz+7Z
WTySGL4T8VtV7A6M3YkatpEdDA6gfpP2AMeEYNfIaz2UR0xKnEX0pOUX2wh3
hbTH7RsNv4im7UE3fB7TrebedJrpxASXgk9T14TCfTFQ11L6435JKBDurm7O
hTHePnseQshCNpxSDPbCjBqm+uLkiCM73qy+DUgwqWs+GQzincz3IqNiJJ2h
PTpFucJF8PHuWR3jsMUrihy4PMrKe4XSn/7tZFHrDr9lTxMMnlqE4exYGtZA
LpU9aNOfL9zJhxpxGa6p/qnJKORnF33QGSz2+fOXA/WW2qwljlTKelkotuTK
IZKkvFCopYddG4PFaUvjEMo0hGYt1K5Rvj8Vh4gYARIO+xnOt1Rws4qKVLRI
+Z77rEJ5UcEdFZFY3SEwKHEszY39vx1KZjLORD5+Vcfaw6+J5ljKpoOXSML6
scyy7bHBrpel4ic45375edO/myvhnX1YdLitLsRIkCWs7p6dJh4JFFfTpJGT
az5x8G1ZE7SoOPcs1nUVZlt/kap0XLCHAFpEPw5MDD5ECHSjzF/43gNCHrR9
1UuL2+7Qjohh/bVGCVylDbY4dVVBxNlhROwqoR+0YXiSUeNnfG/HA83dm5RU
xuHhF3VEZQIEkFDNFQW7GaugYG4kkHsdWUApUNplY2DO6EpoXwMQJyhWRJBQ
tfVYDJceKHb63hYsZqozy808NhlJue1/HXxjUOIYdY4TdCSlvikWJK7HplAi
RYDOT6RtutbmPp2mgRdas/CowO4sz1GUC5NHDemjaxmtSrfXvUTm1kLgedue
EpwlhP4/ZV0fI1qKPp1gZzYQAWd/tgMkJvQKp1gt5Qi/PWOVzzlM3+iY6pbv
mWM0O9VNKs4SXKEEeHlt3sPuFqmFbaPO2CtyjRKTK/7Oe31yU0af5qSjgR6P
ML31ormo0VU0LrAvXsz6ICiMVbZke3dZpHTBP8QUITBgJ7KTYsssytyXj7w6
gGHt5p4Atvko5njW5pL2KYdbrGsMLIxSHO0lIeGxOpaV8NZTHSOF3Ha1+658
CdocxspbLDkkWcKsdm9aqKqyqCqAQV1ZACoIN/okfPN5/tW/HiNZF6wKbcIF
jER54RW3unb7I421RBY/22oYln+nuiiYLDwVV2ih6a9pYmQfeJZxtMYrNIXy
b/FMRzwtMvvJLj7Mts/YrhQr4ttu+jnIZyhpE/IjyqV5L8Fpp+MzkxuHgdRR
Odl0jg3dm0gKyDelVRjspTqMMfSlF7YAB027nvk3GcHhJkdh8lzM0D/PaOC3
zSKZIAZ7cC2doApnRbHWzSRyiGhXDtn9+dl6qzleVIOt/+4SzsFCaRp5iCjU
ecTJUY9pRTsqp4gMbaHn+9AKduXoi3UTpvUy5dgdvyLBSac5MrP1hybgvUwH
xeNtflh/anyvlh5832j+f7+vKrjeBqndzTlpjBg8zXK8CVfdduIrQEWeHkgL
sNzBdg+Tbo72X7cTvTT/zrtMH6A6+wRRyyhGoOUSJktu/tfszJkR5q2X1uYR
3zd6+F9W4c/T4WDpbStJ9G1miAxxfmGo/B3YtlWOP+1t7a7wKyCyOGO8ojlT
MLHd005VFBukEeXnfgZWz+kAFruVAp+NiZKN1y4+1qG5DDFiDUtECu2MxGqi
PhaqWQKaSprkROgeDd/X3DC6GvV8IAmt7AuarGCzJUGpdSP9IUGwBa4nAMMz
kw/sA9k+gtoc72nC8MYTWXwBe4MSXXIiS8qGnSU2I4bzo9BJ0A/YHXjT3B3B
G/mhhqIWA81mi+5nNwijCNeOcD1lvOQCvJvKFrhz4RLWZSxiG96gOsTloqpA
WusHV3mj8cHbExsEOT8B5N3rvVxy6N/3wsiEt0woi8Ol8vi/KtOHmy21SiLH
S64ge/+ManW0ehDmyCxbJo5iWYmwX7B5bHGuLUmdkbF/K+JxbpchtWKtRtSY
Igmoouqgu8vIK/ikWJq8txLrLTGF8MlPDUWB2cQGEBvaGDubXBJI6ePqPMvd
mohREqavh1DUKtpF+QvJSJTG0qzfU6wq9+zKxaPw0P1tLn4Ymj0AyYoV6csk
CVzR7/W5g3YuzpqVs9deAA2oRFhRybJV8qNF2tsRl+yOMKpOUSm1UjGBQvjZ
EEW6DJL46NDfQGj8nxoQRwugNdDCGLpAJEGHsP66MIU6hSb/NvJpMC2zTSfA
tIt0c3cp7McHmRpvm5FNKvBEP++ZoQsTWO/1W0yAsHad25lxfkrWyExa+c/K
HCltVk83Xy27lEiXjxqNjk8wGOro0P4FigoWMNHHne5ek6QQzF/z8xrkWS4c
nj1bICfxh46bALNHMtfsQXHqYAzXDMo8yqcWKqQPoryrzmLcbcGqiB8seHYx
UGvuSdDWaiyklnE6WIUwAvL+VlKRP29sQylW+M1H8Bmx2lHMbJmKZ/aNMkAF
hJXzT05kNmdOkAL5RLdga1ZugYmYYEdG50DZfZgU4YsD18SsHklPr7puEEB8
WUenWoBfga5IyNYzyEwn2ACd2bi6IuY9I3YCmbrP4qSwzDqhFkyp8+a1F9d6
uJtbbq3jbO3B0xTblGR3L9JlRkUdeFPBfkDo+9/9K6BpJacEtHddtrOxNNv/
IJfMQcy+thVrSPkBOC6wr8zqzdCnexIATT6drszo95tO5rMohzgm6cicvrua
qosYinpa8VG3W8JNtrIq+nrgh4n6qG0PkwLY0/wI5miFD+TPXc0yGpNIPYdc
9L1CNctFm0ejD0o3+pp3f8z9n+mr+sU51QrevmcRrquC19xiVOe3Kj1IHC9V
x8fZvtFDnHO5AwZc9kozHuE75+YZp/lmLiGFKQ88l02ts+MRYkz6E6zeps7E
oqoEcjCn5FAiZPzKIHfmNJrehMeFImKlqMWNIYy0lOlRfsS2vLFPBmV4qdr3
6CiOe3e2mhdenSWuS8GN2OUMG4Oa9vdLRK3sD07G69VBg53C1R2WjeJtbtDR
2+xTRjCPzWlamwE2z62TZEjpbPWlCjg37+mJQjrKqYM2xR0uzKsTxcDDT70o
A2UkxCnGGdlg2b3s9LGqm5XV583gZf9vusyAzABB8j0E1HIWQINXV3plIuiM
uPofDV0UoIWPePr3YZc0O4DMTyW9QB6pnKy6J1yaxoFIN/kwGSUIEELQn2b9
hQYiYvS3lVKVC1ayotOhpeQqYW9rzzQWgNt5uitknU/G1rtA5dwP69oHPAuE
Rmgk1p/wIxNvZ7vc3c1MsQRHeNKTafXASm347V/JlnUy1ADhkcRXdGbd5SAw
5cr1lqeIGv8PVoAoBWI/Z/n44pL6x4GSHN9KV/weNh1BBKv/lVHbFFYgHhWl
Q5BXeqoiIVnXJwYY+TOij93TKGb3t06RVcYnwhNo7K+oZPBcUqsuuBbgdomN
sfX9+QEbHk7WZ33Wds/nCYzx962eqTvx4ptOhVGprMAyt0g5m4GHqXJSy7cZ
m0XDY6V2HnSuV4NTP6bYgUpOO1Q1Ie98hUXgNrMiDjwUatjmpX0xhUCGKA/4
G8sZFbGhvh4q9TRQSBNlAd5mqqXfS7GUHxqTH2/zo4BgQpXEYWqwYlXKyRwF
Zh2ESUpx3COptDgRMkI28SCeK4cPkfqRuUV72Ay99glSU2RhLH+zAFBEiSsA
jSmpYHrHSbj+y0m/ZXLv0TUQZoxU1n3vKF3s5c5D1iCGmypaIqXVOsRp3HNh
Q6XhlxKcvmEATgc+zCAZmHbPiYnDv6/dj5X2KZAOSFZSknFKoouRk7hwjyQN
W6X7pMrKqIolyePHRTmeSLcehUmFCSvQsCa/+7NKn5lYkfLVaRlOVb4YWsZy
JNjn/rtiegvy2RrE484mi6LAGvFe0Jv/QjSm+J/wNE5/JeauuZ1coAxHoHWm
zyUINtqW50xdYGo9g5AdRX8PropWLxv5ZXd/lydMpvlEDbNJvsmQluE2TwjE
dgyZhv0hdcNl2cMGuNadJNGwI2V5ES5MIjFuorz+V3qw6qn1KYC6C021VPQW
5uIOtaJOSdUW2vYlWmBP005h0RbK/BtSX3PcjnXxvj9y5bOasZPTPI0CfwOH
9PC6EFunQ5+T4xH20+bd5Cr2qFXBepLefxFhrMqSV2/z1Pjjwdo6AEb5UGLe
kXpmVRaAOqhBHGLTYLS7ZP1SdZp45XqUrlgaxXTPrYwksydy9GhhIYhGA6op
wmXhcyYna++cS3L4rFImeRzs0IkdeJkby/3B9xp6Yq/VjBKP4r5RRCowDZ/e
b17txx0MRo6nFWTOQi+A5QtdF/gkh+h/aGN6q5QxNEz/yHKGi6rVOrEYAHQq
TZXBzZ1Fg4Z4T8vWMd/Rh/O4F453VzQLVIogpIGW113UMevN7k/KNh5lu+Wo
GTMRPN4Dg4IRIuWMpXGZY4c/+Qyn8Qlz+eYstZ0IwmzsbEmSkL6ZeCqHLj8S
nGexL0sDEdJ0R/gyyPa5fZsNrNQQNAHbUvSbkVFjNlSoymVes1a7t2y3ajtE
fcJXw7PIZjcb9oDHiiKhZCCDlspHwjBK1ah3ya+j3T/TtXp5/eZzmO1DeEuv
+GbXdJyG02I6qeIIot+IXqsjz4QTT+Rx/ydTeaCwH4R6wK+uauZyJbWo/s59
1w0SiJjF+9Cq+uVNeXUqxc58yvKEZoIPArUNFg6e1x1suXmEgc377hOXR5mb
T7+C8WvKIvAG9VyusSwkh4PdYed4yWQ1L/6wP/CWK8y3wg+XthOZnCQkEgZd
MH6w0SQtY/QHmvOGzYGs6ahLT2R4itkfQPsYK0qqtVNKfw/ZbOML//zb+fAB
NLN3Wsdq4f6KMKQDx9fZHq51IF3JK4tDFlFxsLihOegtjy9tCdyyRAj3U4yJ
TId5GzJ21AthULD+8dHetcC8o+8dwnj6Zo9Mf3G+JKiLSosUqOx0+v/u3Icn
ztnJk1uj7OkkUJBR9t+udjtCoxNR+Ui9k+qNnw+xKzBLbS50ZHNdh71yLtRd
YsCye8nsDnNOZhJZ0I1qBDLobYDx0RpBhi6q4FPO+tMSOjXWq2W5OudYoxHu
o50ECfPYXCPX3NfNl0oSXORQMZLH+/P/XVXeUvrn1Ojs8dKprh73cTMDYkQJ
z8Rg1JWWF4d7wAmRdGLD1gyCl0DcUJdPt8kygyA8TBY37rS/ZJdqTdMMWnsu
naJWOr7dkhv/f4iYC80iPJXzz6PqrHJ16mY1a3CKZmKsFlJFy8nXtfbXNpup
wFnsk6bDgzQTd/Z5NXz+krJnpAdX4pvDu6M8x25vv32XXRZtAsZSQStpj2r1
0Q/SSEQCoOY0xI9jywRvDJymdCZvixZioidztnS5nz6lkX14nLUYnNpLlIlv
8ZParALg7a2d7nzfmFWbIPw0YD7rjzf9EcZmYCGQn6dqPorUWGgg+sq9Tymy
E9kezGG9FuMU+qKlBezgdRUF58zzGeBoKRvCtNfwZyzDx/2SxCXU2EWHcw24
yyps5w7+MK6q4b1CDUOCmC/FTKJDU+IAnElqVzdfr5TMFH1BGpbBVale7xdM
ZYO91FTXMg8CyX40cDav7aGXFmZ42sjcW7Hh7u1aoXmW81rGSC7UBYIiHHRI
PFAd6OEqcN0JGINuuFKqcCI5d2lvUoSOCyGf/jajRCnOlvthDc+rOFk+Apbm
ki1p5+ilLpCoTmEHKGaU+JPX4iusapaZMy0VXP3OGDx5hxXFZq5JiaFQwRoQ
R/xwV3K0DYENFGYk0h0HEOXbc56qnG7OJ3zB0VLsOBbhn0oiujHGAFOx/1Xa
QzQhiOLzisDm5ZHxRR0z2A5eYiAKTj3gz8oxMsehEj+w+UNPo8GQn6TbG/qg
XG6Qp7QGYoZYwBkQ1Pw/Lf4xb0Idt+IafC1TaQRolXjVEt/R6e2zCDZBUiPD
kfeHUkVrie+lgofkPlQJ4iVpC1fhujBgi0da/ZVWJHR8ci7A28GQC2Xv50C8
UO6jzoYuwNJlQHmAswDecrKBhKmj0ljbkjmr0PN/JjMEJ7iG95crKTiRNgrO
f8USjkxOw8R6UcaUETQ/HhtvMGOc6pXzMqKzJCfzcnBQYD3iXmNwbOgiTpwR
4FxNNRKO6WqlmM2HFQNMkcOBiini42xKqE7IlljnWA+1Jl5EhTW3i916NxeH
RjmODNe7Zt/MeCQT7QLl+xqRFrL8pj3kL5h9OLE7kf3xXOwpgLGwkiSWsIEn
weVeQMgm9oWvzvBIti0wIsfqoUIZlm8QTO2PRoeAXHFxQwImGDhUTvFoMmI2
J1X+KHtk9G4DF68aL8cASBoS4xGEeOxjJps0fjtpKzo8ipUfK6Fg2j9wXSBR
VbXKAlrlAn/Ff2wu20hRWNj6VnEPR1tm1c97VK0rlZAXCaIfUc/XvrOGbp/j
tOFaF2qhJnePSwQpLigK7SLNYV+hFrFeRvJlAjBjVrQBTVb6fJfL3hYvGCC6
oYglE/B5pXEEiVl4z34hkPI3GvXXjEyuiBWY12ngVKhchMnFjrGyGfplTYw+
d6lsjUWWb/3hcsV2RYhFZF2NqR8DVwClGckHWq/WZxrlmTSX/kT+W2yJFZgY
6OAlARMJQFJUeuYDYquNEYvHrlM4FuV4H0n+7BpfHl6uzP1IUeyhoczfhD1u
sSCY8Sii37AvyzTcYXNZfHFyc0U20/i1SALvN1KFzE71AQcFkJC1GTRez+9P
u4JPbOsZWr6qhN2QcPO8pqPKMgFOQTWyFBBNosWO/thsbNHlpOqnGhFKclu7
pC+lVx3af24pI4ptmFz08j1Jd0AMPOzOwWZWjTkVvPaXCE2+wJRvbCIAO9Au
5QYI6skLdlrFzXi74alkLGKBMK8X+DMxezrAt0GLcft9rk/nimY82U7YpYrt
36oBsRw87LO04qvHy1bJyha5q+wwvZJ3uaESVUtWfSpeeWP1YPgjfUhsyr8m
pOIv084CP2eexO8eDhTtsqA4ObRZUazRSZuB+13JXGUn/32epkf8V1M4gUiy
6l7Usn1D6lvFHWUgFo0kk2oTNrX/YABF+0XvDavLbzLTiTv3b3Is2onrxCFf
E0CYj/A1SULylsNjjEX/hVn1mucezX88qIMWknbnJ3Tj/KsAfKj+euvw7BQr
Lbou3uUd0wuFZpVclgeC6IrIBRwDUVoBLaUdbaryux1MNYEk4ziELeUSAuva
HGthpRozwQQHIWHT2uvsc4ofmOQQ4wUlMM9PYRv+yPVfXy76PR31plJ/2LKQ
U+5r147/M/mqawrE+M0J2VjO8+26YWUmdA5+BEvaBA8ceXFPOcRJ7XO/iguF
7XL85b0ptbU8l6Fsta8xf0w9U9INDcReWgVH28YUiqdMfKxr/SyLCvtVC2D3
jJEUD/1Ff5W31AlGXm2Dza51WdRSNE4On1ohy25uyRlg2rPEMsxTTK97WbeM
bmmCeHO8rvz6zLd7W3SHVr+SUf+bFwqRXWiijFRiH36tY9v2qLcRswHSbcWW
mm6y/C4o0MVvCVR9CymJ9brXVD09i0kVEXwGuyyAkoIvFKaHaL6hTt2dVmj8
IKiEKJT/AjrQDnZo9BtcU6JEbd/VJU725QRktJKvXsLC0Dc2q6prVnVBJsoI
fxQlJB7Kzz8q49mXTaaxiLBH4CGHbArFK7KpChnnL7WtKeN57k5F7MWZvKQs
U7uWBCb7aV3a2jK6OSAEjlIox9xJQ+hT9LqX6dI+0tNRQqDBZlTNUQ1wHBNo
MfuvGSkcH1VmabSLzjw495ahfx1npkGY/E4rSdj6U2vrUDWuHHlWY98eHddK
UI3o8lxhWtwkwOWE3WGzqKkgkcobrb1sQADBaEEx4K3OUbQzPr/f5VnA9i+v
SeGnuwsEA7LA8ZzdahlE5UVpT71nP3cI60uicZAby2H4iRhhCTOVlrVb5AoC
nK3u93F/W8tO1g9x2dY5WLPuG1F9Qr4LcHwE+e5BTzerfJwtQQJ/Y0qHR5+K
6brDeolhOKG1pHfPNs5MmAwtLMFJXLSgIg17HWxel/3lG1U9XZf6N9JuC4my
SOkYsHV0ngx8CqxlqqhODhyAG1LIG0v6o5G65q9MIn6daiMhezGw9iGn+7Ss
xj5f5/xe/9MCwuPBrBMgsXyUfJpgKbzeHdZQUgWqYH+psv6nXjvRK3WYz5Y+
BYr9w4YJXgLxV9shSBf0lg7ieS3Vylcz2Uhb3Pk42wQQoniuxcSnwdlfo7fg
a5YzcNpPs7uSgSS7XjnujxUmbCGebKlW43uPkfiQAPgm4SlNgwL2xBtev3+J
1R/JhEd1E/fVkSOjfIuSdPUdEAtYe7883XTaw/88K7cvflCvq6nCMjO506lB
gEdR61wCE18ODmzJRoU0a4EpBIsV5wu9QA6GIfgjMUxtqH0qDmLR+JA5/jaz
5pn5xyj/w+v8ZSxIH5IRA1E5WQCI6yzGTU9Cnlzo4s7YF6PP2qtl2fXvfkar
5MG7z5Y3/yIFDFrGxaIRCWh5XTNhYGUJuTC/AlC+lSjLr4idxSfRnF98QTgY
S55lCVinnv+rCXGZTS6Eb1VzgGkwxFmqZ7vl/ori5UWhswZCydZx5R4wIZ+d
54Di5myvCS68wY/3GjqhwQmCl8ZfLxCQT4vBu3GlfSOCcrn+2Rpln5JYUB6k
AQBP60rLRgKsXfMykYi1pBHBajYuT0SWE6D+d/VlmuNuIA9xnxbYnn4lp0JP
A1f2trzR1qZi6BC3kS8vvv0HHbCUwsa8Csb1TEgBp3tlhzhnpEnqtE3sqMQL
OsCStR43HEFG1DPFdlFuxDSIyYFmBVjqQqTjufufRsVlIJXWjHBztvSIub7v
zH4zeLJeU5TOFNg/HyGOUDcGcxVCIs5wxiybt2yMZKDPzE9mZBwO5aPxvIOT
TtvwhcMIEErOGWZe+EIRrK8+eQVPhcS8MVtBqvKCkm7A8QGcvawS3amrfZSB
1vO5OA0UApOnWy2O0ndMd6bGteSueXv7cc2RYdFO57k61G72B8cMMU1ZIpcK
xTmYe2YDoBNctzYmPQcrhfhCfcAxD3E+DsDT4fWIAV4gDqHbV5Cxt+by8ABH
oZQHzDdZpq6njfk5T4JB9XL1lzyIKRkp5neibLLiEDtsLKKKymfJdgBPrvMx
eGDV8RFr5yMr9NpH3isSvH1uUdz675RI8fZZYSCKSp1MdvTmXwOY9eNZbh/W
Th34w6QDE/0D1rlRraEg5hfzqnEHH3YSjsmK3JjtfZTDK8eSt80Fbqxv9fFi
a2ciDvL5judJmw3iTMseQtAdIPum9HxtfUfAlGA2Y3sV5bQnZQs5Sa305k2i
VPLS23lo8E3tm0AJO+8xdmqDhwwnboUupjKA9LD9Zh4AQ9A+V8ebzaR3WsX1
Y5skuKkeMeLEWomCqrWs/Ehd8L1eYTVg+g+EMkRCeOvFtwXQO8NY5a974tw5
10YZOI+8LH/kfLeTamxPdL55Y6+RuuTN4H3Uz9lwbHdizOevrL/RELeHDyXm
dSIcg9aoIc238Fa7g9JUL5iJzGos3y8KnhclyKc+QYDUyxTO9ecYzEgm7ce1
7iXMCS/0saeKZ4VFxQXi3MEi+faB75HlhdK98lj5geIzIHtuLHo3urxGa/UO
WXHdUkbfgYpGQ7u0tpySl+zjrkzmuDFzfIeik/XpGXTnGdTj2wgxZqDwiJAu
iUZVIujFP2/7rynq9B0h5eDRL/of+SHN6clMMzMU3yCdi6cwrnwKsVGgxa6k
U78K7leZVgoxzYXyzmnLqhLI+LsNsPGL+c8ege2mfmR1F8BVRerZ61iNdW/B
5qszYemRfDjOTuGpgakTRlncFqfgpOmnOeA+UDccK9N//46/bcVtBqSeAjKr
5NhSVSpj19AWfCxhBlckumbwRtw27t+oWy+NlhSWvFOet66vmjk12KSG3/89
0oC4q8TJLZDVk0kTI0qbvQs7DCMIxtbA8bMnSg46g38PXvl0TEOn10KLa1I4
zcPctbBR/wdO95M7r94xRmPxv9SucBpjp6BKbCAIk3mz10bPaCIXK8ZZwkTW
Au1YT0niDQwb7NW04OGogYPF4ClPHbxP+919pLj+cOm+y0ULbohynkxJG01e
Qb6Yd5DILefJoBwDY11UIx3Mf9vRgbg8tGNRXUCELp9oCjzrKCa52EZdEWS+
FaoxrAkDPECAbZXLteD6YjVcO9diOjdC4/TgNS30PtXQhHQidHF6LmuOH+OS
SMyDHPqHhfkGhgyFZbAfSjskdPCtPKGVqSXdHTNn871z236Cdb0Bcr2UjpN0
xttMtWFJH5fDkN+ssz+e7vNXm4RFcKyaezcFqeGwjjZwikiX69r2v+2nfvND
VRuH1eKBfERSMTmWP2EP4BEnKSjsrr9HBMJtCJSeuGtYXeZADwsH9Ie8dVwy
i3AzatGa33XFNbKhj91DvsunN7+4aEqzFLgT5qf+7iBdTJYfQ420xYDePKhD
Y8ltbWV18Nr/YjUd2c/RDSow/hkwMdGgbT3b6px9iDOg+VL770MXXxRspMZ3
nrkkbzLBgkBieGX1iBLVpWOjYKcJOeubLHoWbLIVd8VC31e0nENx54qFq4fe
AU0zKeDnEa9f8Bt1Fwel+X2sQvN/rGiiyqFa8ec/B+3FEJGq1agJsmht9ymX
BoDwY37QZGIIstIMg3XbrbPh2viGxIV38IX2hhzdvFo6MYBkG+968PSbX+mM
rtj56OrQUMTmPY8rYbYyeWQuWKtlHR89xDJAy2Ts96El81QEVpTQ5nYfnE6N
NvN6V2TetPXqjyeKkQp6nN5F0l7L53D0at+an3Z2dFvQ7uE8FIpUIwDI7iwh
zA0pzkT0lsgCyaUGMb+aNpxAu6T7nPvFsZ/45K0t1y8MGDC6xapT6wGvd1+k
qrYhjM/p6xMaPBsTV0MIDe1tU82IfiLDSNX6CL8L3b2ehJoFE3XGJZH8wMjG
YXZZcJosarGvISzYpEFSq822IdjxjNkeVTmPBQmfOKRKzHuyxsL8zgIAW5PT
BFiK8g7wGj4mo0+sc8g1VWvxw73RXJbRxWgKfHQh70A8eiFMp16hopQ7vuy8
BfMse9taVxoXEf5qc8VX17QGV3OY5j0sKZB4mB/pM5u91V/BMLLHCpPm2lDI
jfefLC4EPK7ObGGLUAp2W3K7oxhLEgANIDbZINKa4c7wXwNl3MnhYFQ9fs0/
CabfBBM4oo2kppx2jfncWO6JnNsj2APMWLajUyi+mskSt0VVuHqzhVBgOc/G
q206qjhuPTRHEnEHjXWgXxgKK0p10AzoXiKPIqfJ4z0uxIC5HV1ejQLui2vC
kR7kgiROWVO4jV1tXQ20CPAGYEA25eIBrukN9ezgIVWtA0cPDe+HQuEREKmS
plu+I6aMfL2KxeFVnKhWK5Ms4rVNbXvj21MnrhOcNNFkv7WP0W5nIKzXlsMD
EsECMjgMHZBfU+OwPaOIHYKQP6pSu9wsCh88Z+CAwAU8nPSIghvZIv4GTddR
7x8Ipf2sdFZoBlYo6Za6m6Vj/lw4Sm6N6IS4PbtRJD99viNOSI3vnRlynAGJ
00RpE9gaLnOKWyKOOAfCE4dYkU5PWTx8T+INrIqtYVO+CwtwA39mZ95rntej
yl8im8hxv2SMxRLbsfarNZsPINojepeifctBaD62HNEHUy97bVgsrVl4r0TY
2PfXOe/9mRlzJmXbDzCmRm1dW1fvu8GiercH2R1WZu+jXwoJ3ZC1b6vAZko4
QB1gDhibuFsIdknvcrDhWB0rIceYXuDfXrDvrGYgobpcA74ersny/6z2Qd3h
nRUX1wdSKv5CniQsGTdQ5QVkWvEHRzDLMHkPgnej6Grz/CfDppDBixQGsv5i
IbVFrkGGkvjwBQJB0n02/xvR6WJj1+W2DKTpZW7qi1ASlplv6nsmYVpIUoiS
IIBWQfOGTMwU73JvZjCs84FksdskTrowRh2+WcQ889KtrHdNzSN4b7gEpQAV
HEpCX+SQD/vTDSTBgj0iiFJObPj/EpNuFtSX5D65EDGMVLZI+WtCZ672BR6h
C/SNM/VpHnDqr2l44SBvSXb9dYAmlhh1ryoqMf/HowRthSb2wwFS9SCuCBxd
M2brk45yJzFngLeED7RObQE53XRH54GHcVyRP1oAnfZieQTHguXVAW6slbOf
wsftM1jokdTdDBuIX0noVESvaJcF9UD3H46v3l+McRzRf229oNQVseCPPSw8
4KpIDas9EOS9gC1f61XlCOGO8J5bgR1DKXXc3nqjEPfDKs/klRHbsiwhlhKl
Wf8BdTEHzkU7F19n8vhqXsFNpzVKP/gHSTLeK3/2eveYu9kPQbQ+x0NLWyHH
o0LnpuEM19b5zqluJj6euXzq1pFFSwL/oU2WveQh248x6Hm6bjvekMnEJcrZ
BvABUqXH4OyBNQFhWyz+yWBW1e5zwblD5LtYcoGBGvH5JQ39K3kfVRnIMZIu
BiHN6Gbw2NkvhrrMW3KTHveM8+04+cT0Q6fgnjA9+Gm7s4tRXq2qnIYvjkAD
R9D+OBshnHSJcrx6aoRwot9vQMHa8Do+my5eg95l1w0jOj02IN39lt1mUMm6
VYhMI43UL8ieVO4qmR2KYBSjkgbf6TsskrIcyi1P21bWQKl1x13mez+M9v5D
7OgRGkBvwJbuIKrcR9v6I+JaGAAwayrYXJmAy1nRdm9R3Usm1VhUy7wfQyoi
54K4+S8CJZlrnnCjKB73LHqTZ1XKSnpJepl6IrkfXu3y5W0dqjdTfqXVX+Zv
rIsNJdzOXIBHPMfL2R+PzyrFcVoMj4+FSEPhE+qcW/A1nUNNVKtLkqa9Z7eX
x4prkfCHWqHIjDci1JL3Nugfdwrc5DQKXiOMNN40I3Pa9YcButX5KmoPOwdC
neUx1+5Dz/SIWPBdPwrq5RcGr+J4Oo2ekK8JGiCvZJvu+sWcQqtpOY4U+erj
S5MWGhwykVQ/aCcGvuBBEIfr0qf8uVa8XsfAG96P4aZZoRFf+UEV+uVtgPlg
4UYNI4LIlL5VNwmpjWnyiMUrgq5Rha+YTJrYa+wppPalVwv8BonsDBGK2XAX
xTUS6RnOrwmKAGmaywn9l7+RB9mvqpOfGqnf8reiZEyOV+EYUlFXKXh78Lx7
30aNNaXc5F1laeOd7NsCwbJTd5MlOQVyXi3xu05ZXhcpqgqnreDJFh/PyC6Q
V0dmS+gMMn81oigWug6eQiWdagZKMG/tpO9wy/DcWOpiV7uP1RztNA8cgt0s
HXuSrvjPoGn/U7wZd8FGJeQ2/Bcy8Uihrf7v6S61mh2WURANcmTOJM246GeJ
74mFoKNyqBkl89KXegIEKcVBBf3aSifPjgkUExxurbllvbw1jXnBuIQUPPFZ
dpvkzsAKi3aQzoAp1BmJGJsvrZ4L84v6svVrTUV2zBcs8gGWKWux2S8lsVX6
EJiii8ogIuwAR1WSS1zR5GGbNPv873eXW9dh/3w38kH/G7ASjnJ98tbKx9gR
jiKrTz+dIC2dSVWUstNSEL89LhiEJ2wfmzhWDgmj+PJY0ZjynCGqOVZdj+Os
tNxyp5Z5Wmo1xDhVEqrTCz4ynQkYaZd6/Of3kB4n5cxZq6Kgs6Blcv8aKSFr
6557WBpKrrU/I03RfcqF0iGq2tmwQsxoxAGD8lEYZGPUXOY7ZTor4v0Nrqzf
+9JUoAP8QPLjd0SnZG83MIub6h4tfkdwbuXrDGcxNVB9izF/l+Iuvp4mVKV8
oQXEsBtSeiGSfzDjtBgACAiIDTW/rsiP2LOF6XQ901cZed1vH7NUNX5IdXy1
cXrW1Bpn/PIOKEcc+ruQpddyXKcjGZtOh6rsRIAyda3H7dzgviWFDXWxEMm3
vEk6bfPe0YBAPk2dHhJym+BNUeYhBzTFRRWl/ZE/9J/olMgjo6V6LJ3wo/vj
xE2wNRhjJn1OtYsSrWncmQysY6tKjyG7mL+3TicN0U66jcI2eg+DriiInHZi
goR8P2+0d4LkruGjrawSXCB7cMR2pXyq234gV5VnpvKtgJ9FcrSLOsgwdlMX
JeW52ytj+dfQAzUvz6O2SoaAZ6EYZmAL8UnatP1+BjoPYV/8Li5WLfA6hMAr
cYbXFu1riO0MR4nqnGe6rzGi7xlwO/JLHGb4YeJqhHfILvdOhOMMgBsblmt2
Fj1Jod/w8DrSbXqWrFmu+2ZC/uezvvYd7KJjejxBz0OMAz4XJBRu4CsM2i/P
s83HTMQK4fCz9YSWmQbZI7OuGSaXEqq1X9IB/r+eJwJbxMdIL96DTb5HVTjy
V1VT7I1LvPsNhnNxB2zyI6ntshoczBjC2wLtKllcSJOmjO0WF11aC374dm4v
BsrwXzb3nn+DkcAdv9NM+JlKYN7t+vHuAm556U36bDgV+0+VTERBtnZqFSFu
qP0hMvpYdd1SUdWTAZG/Jud/mZX85EftHkI5Hq/NMKRFDctGsF7J/0ePG58v
US9e1Hy1dXUEvBazs+PXqx8eFtnAxS7eE0OqZFFVItrP/ESrgl/0W/qvIieI
4mWyiZ4T5YSGZb6FteciAE1QTXq7EXj5VN/obOOIOO42/DIJYGYGKkSA9guR
pgC6VwkrdNg5bAffw2RJ8//EEHLHgk+5zfD1KoDYo+Dg8G2dy4Jwfqu2vKdQ
Ww3wiZ0is5rTMqz+wIkPmObIZkMtaSMskhNi3HmRZsS9glKk3IkY9ZfIOwwe
+xdvlLDNpDj9ju0J69+tib49iICVCr9bDKf5w9tR/hmtZ4EdL/g2qwAOclpc
uadnsWKr9agGjhEyU01hVGq3rxxnZyq1Fgb60Hs8M/kzAExoo0oVHj0uho3I
bSH3c+sFCW0CP23iMAPR0CSIghoEeMDK8rEWaKpHY/MKu/JZ4aR3l0+Dvip6
xazhpznCNE1MKqxzzRLlNbtFpHnAgnz9fRYZPE5BeTRJAuJvhVY4pq8OG/P9
jWkPMbB0KVor/3nzX3YtV6HUtOMyR8GtshZImqlqbtVnAY9wT/JLmNn/pzFt
9I9ZlqdWygEX84+pViIzoRkvLj91Sf5OHaPElLE+vb0u1AlNgduonb4U8gdr
gpdS6SrPLg6WB7j+dg9w4fSgF1qtg+6b3ETv69Skkj5d7WTcec0eEi4iYhUq
nLxkiVHKGaWX0nSvToOf05hokdEJsIHYLQtuSuTUS7xLt7uxj/XpD6VvkQNw
RIER9ZZ4emOFkUo2fS2urkpfBoTOqf3pwvpZhVHAINT8cEdSVZUC9PmFUuDl
hzDnENwK4rLU1/iXsQzReMFLxIuSXZQBzNh3TgjsL0px8mz9x9woDvwcGptT
moyAQlQfhaAfqZIWtf3gefngr7ifC8B0RhXYyaB+EE7Y2DKRXv6+SG1ltFEg
kt48xteH8P4pewGm7Xg7l8wdZgwH1XdZfLTbyNnZRMTv/denbuY7H4sQtWCF
Bgvoa0FtZgZ5tb+nTIKpGtXg7MFzSVst8QDXM95loD1OteCZi8qApVypA23D
9xcnF5Aq1jhiv0qxMhpFN6V3YB9PJSQvplpF5GGKTI0w1VojCWCWdIfjykBE
Ie5B1cpvtsCokN3UI95RdNk7XO89houQ+uKF12rh3Vte21YjkXWdO+FLa2Nf
29XDOGURx4SIioZUkk3VaG7kVBrGzfLMGR/3vjcDmzory1d8w1V10Wn+dgga
mfxxmtf2RORstoouTDKUn2DUzyPWhaZLMR5iaEiM+4zuCBU7PN/W8lGy1Xbc
QtmqXf0Xb/XlXB+FERozrUsNOfPgbS9n6OCMHbLwCJ7cjKJD6yf3jZ0oTFg0
3QBHZXtXRY08UyuO+O3fLuQgd/0hOAuCjhAdYYbtOLmOW34BHyG5jufsIuPg
VJDP2biM3LCcbXzkwIn7yit4ahEWSwhCSRywj5yA8uUNGyLXbOhtywR+MZvj
39dG+M7Ff4Dlj0/pJwTzvZwHT5h+eeAjhE1VZAYq+vY4GUs1LAup7EWZBLTG
91JMlBZ983Aoe5prLXt1CSSF+0kJmxUDOBn9wImUroDWt6AcH0h7LL1+ESSL
uL2A2gNuwHStdMX/4O1u+E7mm2T0qXE+JGwbRbc6R0GCLXc38swSLmoOcn79
CVz2NiHdfQrPsChy9sKkZCx8IBmKZz1VbScNazeBJKjWL7JkpF41fiziauNj
7/AG+f0VTbjJ+hP/eOE8zyDlB/V6ls5U0zZI0Uk/5fe9vYNnQVkXxPza1xZG
DpbWMGXUlYl8hLswxNosRgz5tdztnGojMNmCqR0P4ZpJAsmMgQGZlMjjXJCw
inSAUKrct0mjvmnblWAGph/uBV2XeIWbIOaYR/1JpnQwEOrWr4NEqRGhNkMp
PDqtxz53S1jkkT3XkQDgj1yX607dkVq2k7aGROgGdyKyvGpKeIcQkQwgKq4d
rA5dQ6ARRpQ3m0m6MLEpCzMHB5DyyztAwZMCzvLGECufG5srcRdC0KBSt8md
BsuSq7ul9Sz9OcBmfBs9Hbamd93zZcdeeNNPXbirqacoL+uAlCeia3LfhBq/
lRF4Tu2lDb5cg5iwdX/Ok1CLjl4wgh/ZYQmc632EW0LYZYzbq/6dYjhtwUrC
GnNKM4ccXoVftYXtLWiMqNVXIziT/B90ulo/hEL87sPRHcEtuFZQlhMSWWfc
rvlmhvNhdB85trg8v+5lMoGhuLQi4eYTJh8RnckJL5IvSPDhaqdrsh3sXdgv
Mraw2M8rHDlm3EXYl7Ic0kJ2DrDZRUL4vA7Zln16s9woC43uOwsdl6N2kEqa
gfYIq3ILr7EAK8DrJoPi8tGKem+pkllLdWEFfe+4IF3Xki94dWv8t0aX70I3
x1Wgd9Jn7VZr/DzRFXapbgbKa2t9bGc9c9/CQqZDXuymNiSm7y+JM+FnEkdb
Xtf7Lnmhnm4K5B8TwB9q7T+WOaRdcqh3+mL7t4aRawU6U2PgOeF1HhX8OmU2
7MEzadBcrVrUOueZl7/FbR5g/1CPXfFKn9cFok7vCmM67btx6hBEs3wnsAts
5q1xdTiDpBnUqbi4BOkCLd5QWkaERFFJVWnMsCaH7Oc2udOa0Db16Kth22qU
2EOV9Ms/54PZ+HkQ0G1A+QzOZEWDkUItySeH5I1OCtKBuF3qgrrtCLknQMcM
tr5GaCdR4EgV9cKCOCuudr38olfbw/WBOtm/3cnzXlv8biz9x/qWHkSusfKd
6lUUxe+DSurjchzzczvu8GwPAnDtuoPzyyjZFas4ukLQu9UyeUbDBhROLfRC
QMhOuEEtDeNTC6I6EXmNsYDYsN9wmR6yaEPeRSJyxeZg3v/1Xgpm+s29W/wl
OfXRP3/Zxgw4t0BadxZ+3eJgdaw2F+l9ybh5I7PoY7HjsGK3lC5E6hgXKSO/
HjTQ9l6fqjZ/XOeAg/frq9Tsp8MbRpk4r5hmJqoABXZL0v78nQzB3/gd1H0w
TM3Oy5HKVXqRvdjRJOHskZh1C9jk8EeOlvDaumybgAfcN6jQVScr7vyAstNC
+jJ6L2pmNWQEFB6qNoFvUiAhBo7uBjvM7QYVS+U0QY9n3HjRt53wQe5GrOHL
J9rjIx9tgsSLJiB5vqcJV8hFtVSjrqtXfGj0l4bLSn2BiqpLaRiOOgqDKx4n
4kxaQzK89qNFBnYYoWPa3R4hAFYsuP+4AB1gOOcbBGcUkwp8EGBuTOUnc3MG
MParptxLaCanwcUjtEDlJ53CAXerT3DTU5F1+YpGk+d4/piXVXMU42fV1hAI
YkmdoTyoOIOIp3cBldpb9N22nRTVRinPnc0nInp0zX2Oqjy4hrfz6cfeLzD8
9POu4ZRTd3iQUcydnmsBWcg8/K1Ek4XvVbVhjKPFYT+4CuN1aWcKLEE+ms3w
e3OFXmjt97nqt6dr+hNgjJg9PmgK8E7Xo9V9UQkb7Ryb/Ndf2hgPTRo+G7Gm
CukLwhh/YbxOA0UkIoL6zDc6Ohuots33wN7DEd88if90L+OC6koXYLgw5urJ
1FRbnVIbLdPC1gl478GI+UYScOiUVec66XhfepQ/Mf9noSJnxkP23hCHToEo
Sl7Tz4o7uGEuxXujxRegP8nLZO8cJc+j8OxfvAr9yYaqgK0myRiqA010GqC1
f2y9RMoPV/zyIB2StSDjNeco9xzAXmYdmzHH0YDLbZwUKY0DLka56pLozCFD
WJxu8uxq+6tHA4lJvk1RzbXQ2m1KnFJDzLjNKP4/T7XqW2BevDMflnilgk+7
0pyXBmA7/cpbH7zdZ4rpkDgD68JUMmIO8lCf4KMo+gdnUSJCQMAGSt6Q7I0m
FDEWUbqATNbs7wsj5xIAdny6sszrMbN8k3Sq1wRHXsYIQb2mai1mUdLucdxM
NmEQiSC2SCo4rcjdjFfJBvvKzzXtfkirevVRwMbPQS/vOOG//cQAupM9w8b8
UM329v41tc1RCvv6wwZqjkN87vxu/K/tP6tiC2FIZZvl13AXyHhuKKlweVig
rhjJiBizTmPmv/+L5cjFXjmtFVz5haVqB8kDS+e87Skjz2CJTQg+pVJGZqrq
Zm+rA5jqcpxi65D0noZJFEvnXSTdx5V66JR4a3BtPLdgqOPsxkvNErDLlYNY
Gn4KWjT2k7t+eB3U3l3ap5TJjXLBcAD1vZxtDZlmIgbtekoBiW+LgSapRUbK
PeNwGq57peth++1OnXD4q1Ll/svuLaHzcP2O0vECobtD2zEtiL9QPzEudAk3
8cYbmlWyG4u0iCT4PX8lgasN8/OCUle4q/+de58xfrsyWRs3dNfiwBI4VmKV
NzjhwJJ8d2tpXRuorfHmy1lqZlqaKNblSxFPS3eHWq3x3JSC5xlSkZHR7PWv
D6xyjbd+77q8TZCwSzQm1Ri/wkHiOJO8AzVGZxmkvXPW+mpIHMTV1sCP5xN0
56YgUyygjfugE38+y5w2VPdH5UJqGK8Epp2gaEMSL5J9lJW/Wb1LWXbDe+Rj
dgiJzjuBM+c5veTVvJbFTr0TGy00O+OTZm+kQxe9VpPTntoE3Cw/FcsO9hzW
LbaiTSJQeyVFLHRfBh2z3k0VtJ7LCRgd/ZKMfisot9wrv3Sxa+jAy5maDNUd
73jMEWNqTWUNOxQ6SPY7MfbDhU4D5YBxdaf3D4fSwsq4BwRJqCynRlWE93pF
hEaa5ev5JdJLVWOYitlML0/RlD1Poc9IFZaVLzmCV4hzniqqFhvtGpVB/O3f
b2kInO63VAe/wr0ajYi0VfV5RsX5HiMO+rsH4zGXnTchuVPyuCwMBKT34NTn
oJgQGpl0tEP2XrwDcJhNh+tvk0Szu6NkOF/sV1Nyp/QnaRzOrAX6ZyRBEf17
IXoqk0VwrN3qJnqw5lkM21LKbm/eHaJMpZhquCM42H+J+zd3Pl/eFgXBE454
buATCkaJ3iLsxZOpvNMAhJ/q4/4jdSwOTBvMwRjrOFD+vgRmJtHKNjA0FVvs
rTVAbGaAcAbWcGjcPLdm6fx+59UYu/LWyL7/PYTqdjL29lqEZHWGF/gKyiY+
5PCYLiFI6haxJYlzklExRo5fjn1WRNhZyaNuQiHkzKiOHpZ01Y2NSl3HCFnk
4JYCfgkat5V56s99Ki1JhCw9iy3BiGFwBYaJRMevgXbP2TevSKLpbpuOWqyO
ldujpJ6AXuUN3M4DL9JOAEiBnDhKIg/NQfVlXrQDh+xBmPmX50YjYYblOTpU
2WxPPaTRZJQpy6QPMiyuagyqvlWXsThZLHPmsc7zs8mOzxdFuPIaanP6yZqX
Yn5JYfPmCCqZ6exaHbjND3Ylrdh9/ng6/VvrFjwCW03QvEzm28RKw5DORp5C
m9Y1+9oECl2kS9SSN1ql7BiuUxK62qsHE07BrYJAYzIC5XeLgF+q8hgfxLdT
tf2WHYnLXVyQeNc4CGovzAS1Ce0lrUM/wrwFv56sRwY8y6/pC4FCMO8fQ8vN
Y5XQY3bchKc+Nigag1TG6vMfDxdRFXipte3LqGiBUbVqEE2H7ARRRK2OK256
ue1dWFigLgUkZ+QSI1Fc4dwgVrqFqSNNdBZIjvbMz2tlRQlKLToiF5uQtS/K
UDLf5cQd7bHNgUyIhejdVM2zGk9exoJYl0hZIX1iABfmkVMpOR3ZJ3s+/sf0
xRNM6/0MCHucztnF3rhedqp8RTEAH7WElLuCDJShd4w+9NbOXCDPPe5QL0mG
jzonm8jSjbWlNnZHUaTUIO8ya9W+xSDbEe+FP9M1Wh28ub6JDzOfAQ/kaqtO
5Ou4YiF1jOOgE2blspH+uajmnJot55Kv8VxnM/KM0rvjERazx5UMtjfEz9es
hA4zVX19q5DMYchGYjBfXmW6poBxOMzZ/a3nYyyKhipz04WdtwxMyLaRqFFd
4v+Rs+EzjUZX5dfZ0Pdlu2z056tQXr7qqRAzEC6RFFAGPvyELACvEFURxNA3
yPCNUtFbWEBtVjydqiBGT44q7N0OB1pU0Kf83wJ70E9H3sdGYRQd92yVWNnj
SP7K4z7JLgAiWce39qfZjpt5hAz7r5uXGYMA1ePyYvtXyjwyGgPDk9jiiwkw
e7N7aTrm18vU1IF4DKsrJKdIedwP6z6i7rvki1WRQgEI+OiL5/STmvsBQkat
dyQqKvvEXOMU8NaGepBrGvP9dQYleQOd/l3RADTvcvpiz/R/S0CNkQq3qIEy
yJsFqx09NvXWCP/xVjO2jBiMHVB9Xe7pOd100rLc7567YKjPzuIFl7oj0hVP
ueXUABGiuesmW0LppJUd3WautjAj/syfrkN23zPbnxX/bIsw7D8latMU397b
YZOwh0r5P7U/DVU0BVMvPqY43Tp0z1gQoXZdGvW0c25/HhsivDrq4QFpl/PU
IJsphOs2/E/RGTOoPKjjfb0eByy+q/iyClMQ7XAdnsNASc7w6hV8aK01dVFf
y07TvcJ96/BUKtHxQeoRzQzZKytAFK6m/IWnwrJaspAqruZzcHDNsYojeGob
Vru3YhHf1of1H95e4P5PNf78of0Zv5HhupuN+7eYXw0Smun6JBPNi+0kYrb0
x4OJvYxoHcIbgOLpcKFJTKOiuBUkP8y1fvgQzQB7J+zND6LYDXXrmL+SVj0i
CaNO/Meus++q2ISfmhFKEw9gUiURnGKqpPb35lGS/AxMS4gF9baaYcb4a4hj
L9i69Kokru7bhKVRsvPrFvWcAUEdr2DlAN79kJBgWPQLty9pPtmLuOtm2Vrt
t/7Kib/mcyhXknzcqiv0/3sZIJcWP8EbsBT/4ncdBOLV3ergNz1422JrZ5wB
PmyemJCuBvJ8PTnSjn+QgVejmVktqzROD7amK9pvOoysSScR3EyWfq+xUhFg
/p5YVzDWRa3oOULPqYkrxmUnPiOei9cDMCqQlOsEd9idtGcLZKA3rtvmTx3g
3WZrrfYp7jtDmRM+lo/+YCfsPnDY06hfr2k7yTYPDPra/oAI0mu2FMQmKxAu
pYP+Fzio8XiPOFIKZKhqh/fgYZuJaO7EHvkbgF7WMAYSa4zZTEG3/l3b3olu
AxInGlBZJYCpSROFhVQJVhaMzjfopsM/DO1wx+r+WIEJ0VVMtrlHwY6nsIu3
+AXTVHpwFoeEWpbACvD8WpddT4+Ru3WrcPqpyR2Ew89CT8w06fCbopUfAIay
7LKqP6ITafsUKj7p+pN/1eoLSGbhy7uusmPCXlBHAQfbKbacom1gBeM6iQ4P
VRTEvPrhcKP9iEdiOGSqPMzvKTOkH+jdxdISydbvqZuSDg/ZELb5Uo1ZhSMF
EySQW6KBakbk9Rv6z5t5P9wDFNLOpebikzn1ilpPEtMBQBiyCM/FBbYBnXN4
EwJUJ9iCXHuJWm2XqvA9motV3+BjBeaauuNXXaoF28OpeGVQ78xwRZcYPm9U
y8BDkLqbQllM7JZj0/rn5Xx988D4+5q2O69Cwx1aRAYH/IQuUtL2cba4J40S
ENCj0neKiHTFYbrHQSafdKxuYWCKN/bVe4ICLfSs2Je6tOIfN0eDRjJQULp8
8aBOBlPuBi/e0IpaF3PG/IPbWubPYnt+6hu9fzgHkO0c+6S2TzFDpzEf57c8
V5ieeHhnOnZBirTCJVgvuTEJs5laFNt7OO2LYkcg1iAQmnBMzwlGoX0DT5fR
GVd4gsL0GuwMpUBjo5KSLD0xpnsOELOWvxoWQ8FTD+3EFG87xJrjx+TpQaas
QZJYzUQjAMrwuCQnHG0x7fi9c1nUFHcoY9bu1u6hwdSNyznCz479E3IHnuZm
6SUS9UbNefGbOSwpFqsXL4I3ZS3nXE5a9Wizcr4FZiVjA/CIN0pz8MP78W0X
CykOiyv75K/elXxxnni0b07mtGaJN8ZDNvxKyziv+NPz2SnSg880pWfYup2D
Qabl0v6fPa2gFT4BPpmVnrCydM63bG3U3fjO3y9ndTAdQzNY5SxjOd/5QQpL
EPWxvfezFPhxts48NF8b76hm4X60F/TlcmO4FVlhiSlGZ+51QmsnsOT1ZhNd
kA75Gake1T0HagLED8Hfwg1MxRMFMU/oGvqmC0JW+wwCWM4Bao67s2ojbVRs
5cHgBfrwP5EileMpxSnffmm5lS+eL293MP5VvB3FqUUVYj6rpuhPJzZSfy8H
9W/XjPnwx7uJyd3iBnXWF2dyuqvrQDlUO1CVUFG2zQYaYQwNfcEMcPJitYa4
eZT96ABqhfHaW5PH87dYDWgRRXF5M8foJdZhrHs4sqnkFSbiA8T+C+iJSLQm
v0XjoWzy+E9EC0PLO90sQnu9oKnS33bikDgUSJWGBcS4BATfJViIhleDRXay
4mHLVbEoIp+XpVSW6Svvjqd6bQj/NueS37Vz1N/7mk7jf1wDv4U1l8KT00b+
kqHXs2m6yKco+RnWpLAIsZIJS9Ozs/Wsrdapsh3s+s7EZ4Qv1O3HFcRkTcua
RkBsy9tYuYQIqg4422vUZIXO6MuTm8pyME2WkYorzZr652byAMSWMvPhQTdq
TbHSG5UdVAopZx3/3Kt18G8629JrpGXDEmfUjtTI0Tp8NVeqnm8UcAdpX0UH
B6afRk+EVPmmqPnL3u7XkoPXTHFL/FZWad7pZyOjDHRxniGFBY0BIoZFTenU
lQOwoVntiYahb/uQ3g4Pugnx8btsAnv8sgiwz+mFfevUlYwJ3uZOOvzMbRgL
KQkHSI10H3L+ITRa67U1Woy2/EblAuRXP31MiBSOCzo69KbQ8Pdte7L/4qAX
QO2ufa6jWU36J7BJhxe8GdeKCvlMxpvAL5Wc4kkFEBDyzERSagOPk/Hg7ys0
DVmiZCGXeKnI9z3f6MyU0ddPfwVDYzRWR/7oqtDqxOkggllwcHhprBO47RZe
nZEBR6psfl2KaGot2U2oKRqr769yYMvnUVEf7D0yEo14MEmfmkSDuha04FeI
KGl4rvg7wuWJ+jQoWsMlp3kqbbOYMTy8jjRhZMLlZUbDgNe2B7c9XWsBs/Xo
CtwAZyn/BEcIiSxS8/tqmBSrIWVtLGrHXV5I3ZpvL9BfF3rKSbaJCiJzgm8J
xzLw0qChdkFLNEgvhGj0qrgzsfCZ/2U87orP4K7uSP/INOS/iAWVOFrul0LN
+JVh6Vb5qJpBWezXnIfrc3xM0WzqsYwl9quXA+K1+VPZ1ZBfpS6VEzIkkEO0
72qsOnAmkwVCPYVnCfoAR55laSeAZnGJVFFXtjcdeDtxXNT0nVIz3z5I/l5c
xwL3BWc6tGTtbOOHo06U8DKPP71+s9YYrbhI68/pcGtD070Fc7lU55TeIJlp
NqC73XVMJBHude0T2k4DydSXGNhmqzHW7uTwDwgCqklSlcNjL43lbOBPjbZt
HLadQRVajCBOF1fSZa/4HREjGqV5Gg1j/P22SyMuQchHVZwR6VzauFR4Zkyp
GnYDSoa9ZRegi9UxPc1HHBuEJkTHxNBPKV0po52YVnwV7VMuBilxYjzGKxuO
ha1hMuUeEE4I4Aef/fqRAPGaddXGB7jfmqxID2tRjRgME+tcSvSNOHLCSv8v
YAoR+TTe5Jw1EktwUv41vVPJAvxprHEF03aaA/SmZaur3kTKZdofBb13dmmu
nkiJCII84Hug2qPbAPsvl08nKzaFzxmCLqTO99DkhkALM1BneZgu/2srDciY
kpUf1JbZyHKmYeqrQqC8rEqqK8BEqVxEZ9edpMy3HQQYKjWzZDgrLfQNvd91
GeJf1dudevqRsvvR9iqz3sD9E7iJyqI1VoSZUZZCfJ7U9Cfy4veiRgkEKOXZ
FDuPVggs337259jcedYLMzPbnjgV9XVIK0bUNjDEqbwLkWJpxp7Md+OszWGF
DMVdpCN990DZXfa6ewtT48cDm5kPSQkgXj8csDpmcZz19bMKhpfjfWVgKzJZ
7ABM+8M4uD3b+igE8+Z/K7XC5Gt3eM4m6vqClQ+NeOROry9Vz0+xPQbBuJJy
qgRZ+58jYUt24FP5et/xSujKpJnqGLlEJ/5a0MpOzhGfrRBFYfd/iHi3rp3C
VGQllAn9xyV1XP7hX03YoWw7kF/xMbfFtUdtc3q4pD2yR/otoFTo/Lfbu0SC
KrPEY+8BmlvzpYIL0Czs5YoJw1vG5jFN92b+RvksQH1ot0QS9eDVi86yMYE1
CE8jyWyoa3NhWnOm1JG5YD+ojse9K4QKpaY3G6aJOph1a09OuZis3Z1YjbyC
BpMAtpaeifc++P8C9eBcWTa6r3LMEf9nrxM+OtqXVvB7uAUnHRJPa8x6MKvo
hEVIvKFpRbKSPqYFEx1RsZJmbdK+mZG5ZJ7/PeU4o8wmPejBJwZWWp0kmV7/
lXPBxUrSapqA2JsJ2c9OpJDUT3vQvJb6ElHFAY294Co1gCp6zKhtit/AJjDS
xD6e5Jrz5JzaiVgBO3xjHOafK6eR41tIqDZ0VA62bNol2dEfvoVnTblrLwnP
kze3YulWQ1xD1/zcJNUDzcIcClLeJ7yNQ/1Kvxn8DepsHCgvRPqUqtDI8Y8o
Md/UxK+RljoSewGWaExUZjnVu3LKg//XBNHOQGQrGhKewZON2bwb1Dx6qqWJ
SMDQbDjqpz37vAzQ12cX/VEukUm87YNQDVNsQi5LaI0CFdN6pwrWum7LeRnF
ujv/Qz7qmh0FdGWSKahT1NoIPFH8I1EYeQHxQyVh8SkJRgMNy6JygPsEZlzF
cfQdvyz9cWYvl2zqvvA9TOW/Q8++i9T5MZ4R8WkIGaN/J5yRkhv1ifEqkRAI
4Sbwl0PFncynriUHSfMzVjNgGxGyuFQS3L24KL3xcYm1OjRmC5zwSISyM30V
duek/2ObSkJHUcbjKEPWasMTxkjS1bAteCRwvaXtQGt0ukUxsmZPuTdI0lZ/
Ocw21OuPFSSIgkN70axF8Djosait/CmrkyEsrcuzlCFrPAFgN/d9wa+X4HA9
7OnjixvsYWnHPL0e/Bfgwz5+bLMUEfevhfOqldLx8QHqdXfdsCeoDVxbrqCm
8t/Qweg+6uYltMCMouZq977kF114JWTAQXDUCchdm8QDaCgI+2kNCYyh6EaR
QrlU238elAd22+RJJfbc/0rrR9HXTklu8D6c3/sTHPnLhagp9ir7jS2bveJZ
uZLWDXLM5Goxsa1dUi9vo9zp7BdjNrOvWYeY64WgTGYe8Mnv8VaeLX7MPe5D
3XIUvBoFXRvZU85nj+YsUEEnxX27IiGHHtUB3jmoL6X+LmglkvJO0q/pdpXM
MeOAT4hFS0nEZzkOPgufZm7KoaTXQek6AeheK3OmXIbYFJAZoVGJpB/fDV3W
x/mI4x0aBi1gh/iMSgShMOr/UheQwRKWbl8QPy1/nt5Q2N4QOPYvHCYjYnJC
oB2vQ8Ukp/HjqTPo4FbWjfecCiExASr2V+BqXyo0wVWeAuAcWpcj3yl9NJVA
Aln/s8H1fJh6yZzLpJ9Ybwvg4ZuHLfQGZaIg+jNFekitB6vTaQZjb0DIXyxA
4lb8xGBhr4Rdr3ZJyYethNYXYUt0i7IzFi5I2VbZuTr15RHK0Jhby9KuTCWk
kUA0tprM6ZhF+mis1UaKFN77OXfZ1hp+ebWnedWshmSZEgsYqVKKCjQDAqwJ
2lyD3j4UcAJcoHMrhsqtB1yd+53IM8Cl35frewENGOzJ/e1DHLmev3Lfaaz5
75wArlLdoVuRGvQGeBPqIMpk7vAyijBy6reOLNgQug6Tg5AewwweFwvKmrsJ
NL8vYDGnwU3+LaaOXZh6yTOsosH99+vOkNl3DdU6kIfd+g/X0fHE2Zz4KVig
yRzUTksPW12OSIZSWwGFIkcfy8x8wycJH6CH9IIFS5qoyVe1AHhZGjBaa1iK
yDqkh5MAU1snW+zrIgjQKLd4V6oMnTIcZbtcmUqcNWSw6NvoC/Zc8eLFc3E7
W9IwfQ05gh4vr8nzSeG+9PAt1bB9iY/mys/ke9bmOIKsYqRaY2IXX6cEi3K/
myOLL1MYmTPyGPp3esMH/ZmR+WlnrBIlGwfhgreLKnVhhBoDHqvwMYAYx8+J
hta35dtP9GQDywR75yHXVw/w4J13jTLa9GeJEnPkyAdIWzfucB56px0hiNe5
WJlE7uSPNy+ZHelmr1xtIu6WY45bU+fhlfzAwfAKoMnS8MAmTcQZJA9nVfeC
6kHcwhAlg01z6Ra68A7URYjubQo8mFPJVCOVY+0Yu4mhdntU3rCcuZxecMAb
hCwoPbRmw+MLoqJ+l/+vSXis5n0WnuHh174u9s3u9w153URJD0Cxr53AtCh+
+ClIbBvYw+4szAlJrPkxPMs9LRxhDw/i6iqnQGx+spr8g871JfDrZVjNgXAp
8hPVHeCmoDG53l6V8+UqnpcAoXryLWPbIWb9e4nQ/26DMpNxI+p2JH9NnzGl
ILReq/SDebgVjwjclju9kqS1zpCH2I+vvcWfEkzWY/r+aGOauYrSO4BYEd6o
ZfqGmSJG17K8dVvciQ/rBMbsT2YvwZ5HlL/EhqBJK97e0ZdYU0ZrYGoMAe+X
JwqLJUZ+I91906prjEJOnW0Yfb/s2aEum5WtP6jikgLgcXcBPYR6puaj9u2u
0EDEf43OONt7ez+5JoXx+N24c1edihKZvNNsZL2oE5RnLEPhNiu1lrvde5QH
BOamiSqmhlmIX6rwQ7do7R+SMlAA+d4NXVzdH6jtAggb+Janl7fMfJ0UeLbP
Qqxov/fUcRgkbRk6tWVV4mR/z89K6yoXbKaf8o9rV6UdYNy0UDyOUixVmUnE
qTrwb6p1KAlaMvY8PzgymUD3Q1O+xziNE2jswYF2xkcV7zx+o74OmNeLVfpP
KPMeB1kLXM4b00Qgiqnu3HtiNeErbqMVoHzsjtbWp3/Xg7AS492u7ejDNS98
Cbwj3W4vjBnNHC8kMmVuZ86p746Grulv309ORvMrLNQ7Q9F85WxKFR302um9
RDuMKUw9i1m6Kf6T2c3TCz68KcLgMpfAISQi/w0Aqt0b7Ser6zjCn+Va3HbT
Lefs70Gxaydq6WVEvFcmmAVcIfBCE0qN4ejKm3G+Ts9GU2+3V3+EztkLR3jJ
snhUB1Qc6MmNweaoEmA2lUr8Va0M4vc/eg0KjCfRIoX7Xld2GvXXWdd5jaP+
y1Fwz6coAuylhnpIeIBY194zd4wj21YeQZq0SPYHhXBsfDMB6tPbTvmCcsV8
0JplYJzs+gO2YIqMiYYNOsocqna75hBFexNI32KqnFLhDoKEXAkZPB8y3Viz
QtsSvE0UighJLUAse8yQUrIAuZi0TG41bssUe+YraaWTGuTpdKRhDMxKAgGs
6LcJAWtv+h61AfvFpLyUgeJA2hkbBr1WSeDcSi19BMwzM2Vh+byveQQbYtxK
ToYItLFTwexoeOGROu7LEE+HDL7bZsoVrX7nHyhYVY03zG6M630qE+GBRiHu
Kad6q0JbE0cyi3ZtpWllpJPth2y540wgGkGmip13Wqrr2IHF9rze2xNejt//
FnIhEcrOu8XKyWCpqXD6bsy9vRrFqoGZmFGkiR+LUbdD0fzHY7jdKwmQQliV
I3pK5eIM+9HZJnYEFPicPRCQFa8zq1cYFbYOukAEngmBF/5hbHvRLxKFfQf+
kOvlyh8EaKE7iSTKEoun5Ss4Qju+fHUe4n5wkdqIKIZQLttWlWeng2quyRfz
3PGdtI8mOWGKJ/JKwkJVMBhNsl/kCdpYng/jLRalC/DCNgIBgFsBkulr3LAH
FVvGTC6cKH9ACjS9mnyWUJKY2hm8NHlDJhZ1wNtlBxGELp12B1bqbrI5kiBy
SFkAVeVTOhlpqNVq9YzIzq/9kFCPIbzCafbaZaDeIgQ/koQedf+kn9sDkICQ
vaoLeRHgsYSm1h+5UitHNZ/nQBScF54R/QijJU+61tJ7BSCRE6E8PgFSQr6Z
II8u5wcts11zfMY3B878zDNOa/YyS+QKgzlXPgn45ftRyslQxk8LQnjrwQuX
eu5hehVog1Rub/6PsQryzGTGzGhCbhBt3sUxFNwgibgenwmg4DNLfXGseBBE
9cZ5LUYLuBKAaFiWpQG4hLmSThahRpIbvRmbhdlwG0GRJEqntw1r8PPRETUO
tF4/PkO0HjKFh3V0SkVqKKiHJPkoFqoMJwYmKnI3WBRUq753HgFm2a7IN10b
bIqcU7a8AoVGV9HluiKxrVQvIYZv3l4N5MmZxE65V9vf2ErzzO7C0j47xBc9
6+nxunixHYhPaTwDNWuV3GR0AXhRUwPqbmBljdslYY1K8qsQwzsy88TjG4Ay
3eQMZ7PR3kjpIH278p2lnR/cwicW9SEB/wsW0gcSWGmTmvXjkUIw+/6JT2JW
KqjGkgeb5TM2TW3LFQL4zIjUM6GlDyXQjbpmgSVP9PVO3bbCwMTEAlGhIWcj
f8f61+wsDEnneQDaJeCrrb3FwhbR2vLPPRAQZ6EM634uAb6WUwzPHi8g7A0o
HZU6fmvPg0OxQ5zHovGtB/vJPG2tz8TSNHJRAZ25Ied9c953NURtD1nlKQEq
W+TtBe6KE+RBTGB5iGG4e7nPcycXeocKViaLwy1cjWG17mffAxty7UnUzLoH
GBW+BZpfGg8/yGB8LuDm3FQ6zgL5cfob1LGx5gh7cGHnJUnbjeYYuGVASKtx
MaEGEcPPlhV7uXG4RI/FjjZt//F7SCiFt1LTZdL0LpSl5j33VTfR0bv8tDm2
9IYBq91H/MVJSvMAoQawDWXgXfnPUJx4oJje956g/iHQtYxc/pu4/Z0fwKM9
C2FYq7sXpv80xBuvuvacoIOW5BEx7e1sSX24CQqEkX7Nx+1+b2RIqGowOr4w
921ZlswXPYh/s/3z8192yWcB5hezImAg9Wzzj0LHAXaD5tkqPbpv0rRQosK8
DAtSIAxfLC86n5sAlpy0mHIUjxpoMmc87OXdltTHMF8pXgTjEOUERf96S+5S
BtEsoPanORauAMIR5b6rFq9XEmWtFkY6GSqG4Z1kp3/l7iuMMT4ahvAS4uMD
9zeyfbbkT6PYfCPAGXyqOv510sH0Ad3lwkC0jITxBV4gnk7YNMRctReRyljT
aynO4WGHGLjR5KYS8pLG6q7oMc/5fI9xJ1MMQgH2a2czrKlHDMnKNRPdm3cA
Y1HHO2UMkr1Y6Fqz99aN965SjMfzdPSxuG8j/z2lFxH4jxp7DtJl67MP9hQG
TZ9VtJzSFzfuLXzeBr8DASCJVrcSlwcKVHCgw+Xmmt86bx60m1NTEuXwzScB
yFEWwfc5WMDlMpZyAVZRmnKnk1gmRiiA3fGLl2CsxVnBg07c/8wPq2jyynyx
PF01fY8nBZqGmzDRMC0HWSnQNGJmJvcS/iVzYApIttW1t2tXnJxnXPvdPPp5
aZfePh7ofGAm0TAHjj5BTdnXNdvBCwim8xBKEhdXC9NTZn8y09U4yItjZLSv
2q8T5s9maXB9jfHFnWFkHxkdsF7/T+DK7e2mPOSesatOueHAVXQQnTpxssZD
oTh0UNrXsBFycx7zTH72fUU23E45AUEm5NSohUmyGHOkgO7+mXJFXP4PT8JW
mVAPafidAlqNyNlMufTEFq88q+9bXGengfxaHtnlGGn5RUhtpB5/Ai9iV+se
IpaXwDZ+U85mAV+USKXUTNwWkGlVNnEONqNO1dOuPrU8XfnORuRvufPklDwx
OhdyHy6DPyofCGmGUqmzqO+QmUa2rM7Tu5Ydq/OLQjC+xaC8WLj7xK4E1Nj3
KGkIQSkCkXEXkKyMVd+WadkQgUyDEBT8J8A5iXkbNnnJtNU2uWoXwxaSWj/F
rnEKIuns5tlL2pJx+kfftqPvKD1NtIjM6HidrOxRuNbmdUuj8aUVxECK7vBU
K5vXXnc4uVEV0O2n0OIEUWIdPvBSDYO4rQ4ArI7Uzn93jPf3YLlHNzoeGFRv
0yVXenMol72jeebfFxKP5ClVQy5UVJuur0QQpsFNs0TFGu5S/mXkXP0AzPbH
LVQ/YuD740tbsBo0jW9vfdwRKUMTXFIbAyGbXVQCQIZGsdxT8tzirij5R2KP
QBR5CLm3TlxBjNbe0TH38csqaiDs3Kl1FFbsNUD15+khtWMnV2oREXhOAF5J
9lkQ4p1D8VNW3KB5Iz6UMln3kLRxuNfYxHX56Q3NxhHcWuzot6A90vcMskNz
squPX7KoCIVfYlPKUEHVeciWkredkz4Fc3TDQvlq0rG/y2GiSKHOKq5dAlUu
hyJlbloOrg59A8lm5F5lHQ+mq4WodS3zkzwmnBu+XANJ2QxSyVQGOYIkUr2J
VB6K8lgZz/1uk7MnIBb9kv81wCPCsWvHmJ8kUqiAvVrp7zotl2A5tnaDSSgc
DpnhcSwYhd7gNP2fZYNILpl0b34Am6RS6ZJuFtvee5bY5Ez0WIN0VS4n4zHo
+XdfrJWw4NWIleMX1zxCTQcXvoErvMAK4fNrz5JdYTKBce73bhdyQYKuNBPY
Owze5UDWhalQHXd/jsDF73EdlLn4rU/0rh/8np2BFZaAMvkbVdkxGiHC7Kny
qzzd1k3HenUBbkKkGujfIBF6ZWVAjzJT58+Hp/NqNrCgyN6hGbJOZoyx5m6d
Z2alJqi+024CwoxyrlffjPvJx8MBDmhZEPvwH2mNdghGcissnao5GYw3eNRv
gvEDS72nItdp/DG8iGZoKM+U0r0NNxdUKlpMCeZX0rMnHekIG7HMfuaZt9Sp
RIfLbx11rlY+eV+xP2zxqiQuzJzmM3bFre1Y11PC4QM94O8HyWUIyaGSvJIJ
xWZleuJw9S6EHw3L8fuFjKrGq0Z6ZSICTNXd8IQMKqhO8jWo9R2NulYuvHMe
jLiYe544G47bYZYIdsFy93ko97NG/GQD4W3MYprEJFu1N78QZGFUsmtVBG1u
3dX0ucdww2dUh77Pe+ImdDHL6dfNsZqP4MS8P6cjMbxi+8MHlzlSAIIo9e2I
jc/8N+vGtKqzbuPC/JsXSDp9gRh76zyf/aEyCI2lZyGOR7qRSoE3fLgs6cq+
yWBZyYg+JAmjrAoYvwni/e6kFmxHa3lHVljUEdRl1/DeOHUNI1I+mjK5OWL6
NDEniveg0SqVvPJn0bw4nC1Pqj9NftOk2onlmLSoVL/0YW2XRPCBnw7GUfgh
V2/aNMWCw3VUBaRceoGxW0TdlqOVazXm91L575I2LOr2aSuXMjmcLHMR1r3X
/3/msWXFUyQ3E7G4PShAcUkPiXuu3qQ32WqmrR1ROK74m9NPfmu4tPtihFL5
0n0IYnBd/sckASsrwdexOLzwlzsRXuIM+bsIseGv0kfkHtx7rT0pLKTJOsAZ
6o4M5BdFL3xY95vYXN1oHz23n0rk23rUA1eWJH33sApFxFMyn56KYuBXgMa0
p5hqYofi3vihTFgU4MjRxs9TDGFWqztlJ5OCdf5UnPz00mecXahR1RqLNjDJ
zhW4I6ed04tU3f7BuGSSzEF4mu+ILiyV2ye1du4jxbwZf4/31Chfu4aLAN0B
CvkfZGC+JUL18HP0ujLL29xP9UTIEFFYfOyBfxesaqeqebFDL1FDie7ibksc
VGjNSKg2qAlMNnCFUo4wkZFl85+KqpYbmqiS7nsujUcepUTDN2e42/0Dmt42
J9foioBuKJ/s+3AxCg2jPXZFPJ18Q262kVHROGg5GC0PRlUirdUUiyZiA+Ug
wPC2klFq+p8veVTao4Oq6p2SyJSPQ4zUCw0rh99DmHOdpLRZ5Q1p8DKx9uib
Gbe/dlsravrCiqNbejbsO6XwvnIFP9aFcG91dpHShSj7U2WwFtFFzaKlC+/A
4b486uuKuM99NiXnBn7myowrEH1blEX8WQPUVH8hLxjK7LC848CSClQHOpK9
VCYCoSc8NdCYVeHfegi65vIv8diIZVLN3262Y0XsqLYd1oRWnjZS5wbWkwg1
R/1MLdTspPcPNDtRaMs2I2X2qPstGsY4v14/xWEkSBaCZkmT4P3iKnRz7/Mg
VJSgaYWCAJT+WtGqxljLuaxLf4DGebHK+tZ1AG8GkzcE3LEk9ZsE9D6/Expb
VIJBvB+EAis9WJgigdyrT1x7AAfp/8bPTvxHHbhIBwMGOEYz5U23d+8F4hwH
KkM/lDhfLcq8JEwdrtdIlZTLFfFd7ADxjcdrWBYr5BiR28aqGC4uqOIniqIC
CQwOJ3UoCBNp0As27A92ZVN5IDoURXHRtGxZGeuPbcTv4k8+44kB94LaDF6e
9earUxRWqm0zz2ADLFUqTgcWJL//jPXBH8UoLFu7W1234cXUc8IYcZSHNrtl
W8HPWBrNaTyr5AYg9sfqdCqTJsbUY++aPoOvHTa7ViRoUPwxZIOspa5TkHdE
GQjUGlm7e1Wnl8oANosvGS2mp0uj0DcvFIMUGzdG6GB7BNH5jcqDYxnWa+ys
bxLRzhD+ReXRR9sKBnILn6T3EtybHtMF3EHuLzExrQi5/nHCXX/3Yotv17zE
HkKgVukeA7cVdMRwJ5cnHJoyKRZBcjW/PUiSjnRbgz426TsLhQlIOGZexiwi
v7MG+8NubAz5QAfC1Q9+qFwuSeL3bEkYjH2ntpTS2Z6/xVTSZc3CCg4ak/9n
LdzevStyFfIlTSR1jWEo1Y6CXeoAioPMjI5ab/fbcoHmPAXXljH+1PKUZmw6
BqU3lhn/xTtWzrqcJAqPPRDFqFXAq49Ji0XAVqI413jYU8Ma1UqGJGkFfhRz
jek+NSb8l+dTRjd+a6FRnnYqgWqEFXa4OsTAKbMZPkRNAvFJtpaxjOrXp45L
7vGoP1KU+Aw0GVY5VebIbq6aYvQ2SRlC/Ma2EFda7Uq8HTKKxQVqafWYeXDK
1qZBXiMJNqj2xQNEOjBq69o+4cWAguqUcvL4iBvbOlidgLDodCU65hfzQndh
cKqRO4TaTT+99nj4aTtiLBdnKblQJwGTvZoSdGBw1yTn88Prd8a5DYsKzK2d
FKeNECAkUT6BBNbY+jEkdvctBTSe07li72SB8S//kA9XXApZyZ1woUf1rZR4
itxTisFmOnIYwhrozsdtDoRqo1vKSvOS1DfwwETbYXhSlouSfk3lBaxooWLM
BJ3KUfaFS6n69QdWKT29Gs4GHCw47U8xOd8onf/m+jz7/kf7pSeKpRgoiaOT
QNlV2PveZLIbkG/Ug5uEJubNc+mnxCxQu3bxoHiuiofpwYa63NwHO/twyHA6
WTWs+kqC9na9QpJgjpBk2UgAqlGv/Z2pYk3zt6EpNaPoN+IMAvLUHZ97RT3s
5e3TNjRmWhT5Zl9a9r4gPG9/08GSL14re985T6Du57XuH20Cnm/lCH/4kTkZ
ZiIX7355jt6wpN41nDyGGUeO4JFVrsKPC3XpNMgR5ptfva0i2JuM2s9IEhTK
Zl8B0eXOVBE+NPn6b3vDn6QTCrkbEQTp4z0NQl0w9CzGA2tfkba0kKzrvGFz
aS/QhwgfSj4MvfF9ZLuONuTHJ60/UfPEl76Gd8GqAQJu++n6ijEtJ+PG1u7/
Rx3Qpc58tA8Bs8gthnrG+5nVqhzqApT+e3JtrRsHBDV4i/pAEgsvSVwGFuTV
gsYK5Jc+/jU0SfNipsbsGb7H7atBB3asCWa2iej2g68LuLuUUYmMP3gGMoug
h1oGTwKT35p3/s2ldQl8+kk9Fto22f8OHbD3F1+FsKgg5yCBaqdDCcZthJUf
YZlrGo8//o+eyli1uEQQBmBwcITDOhrIZDoAtK0JV3dfeEZOnJSQ7mIdGMQc
FmfQFEM8LGIV0hY1GBFypUCSLRKrEd4l6ivuPJSiHotZGXRhnydKg/Kxs4vf
NNNPqGIa1by/8t+EWD83KYoU4wsu4i6Qa6Yy1zEzV1NuAtLVXm4m5uJaFpnJ
Ho+9xEmIioXnYONarwafDfPwTYmBJ+5i/AbZe/ktgY+PWCvNeCUxZiGn8qbK
Kpo+X5/t/P1T2OOphONQjDUL07G7Uk0wCHAflWAhFUWPQOM8MRgRo8ampf5V
62KdqesmxcBL3I6r9RQwz2D5QMZs2/mBzMkYRUZtR1EQiNFduHcwwZLS/nFq
VPpZe36l96ZRF8xrsDPXtDjmdn/8BqmVjptwOYGeLQZku/b8sR6E4aeLOj1l
KwzndI5GWZUJO5Fuu2s0dpEKaQRuPuiwby7PUaJCSzJ37R/1IPNGFYE7p3Gi
FGRXv/qJCbiF4VHkCgL5/T8N0biEY3CaT3OEdg+thx9iY3r6dqOcZ67tna4h
USMZV8jIo962hOutQC0Od9alrliBqCKgBVpzgkfbGAtfmTDK6/H99SknZrmr
Th/waI2nbQDLytopqVslJr7Qb/30TBQhHHm3LrRfvwDbimK9kPHZgibUlBdB
egFdchCbpiH6xg3GU7QBXNn6iad4UH9IB55dbDdc9oEo6Rd4Cyr0c9Kw3mFe
Pn0FZhYiJ4riP0NR5VmphwqIhmKkhBP7V1til/BdeyJEpKYsr1c47zyJNv6J
AMankaGX114a4EI4WYEK8PN2vZw0o7AQjWOrPWPxwioSReGpID+hiIwo482B
Ayls2fIKkdOppmdaHiVtn/NAucy15WZ63kkHjKJOo0eXkqU0aFhItjhlaiqu
1apF4ERtWt1fpfATpUGePeOS+qRLOx6t3Sm3HKwlR4dDjkIuHKwnbBIiYQjX
9sfhw2D4g/ZkIHBzDRNtNDyZ3Fk+IPhNRfOi3svZDj1ckwiJbjLUD9x+bcc1
FzSiTEkZQgb2j4SFZukDH4L97K/zAu0pVsJ2CCQZSBMEjbrM6J1UtSjHR3Q2
bpnserJsp91bhj4BmTIrYh5rqKHPeTWjjFcG/tXSLDwr+i+9dIlrGMo5D27l
HGvNz0KC+0a+OWiwDJIkW0I7LXt51N9MV68F3UOsB1GWEkPpBLU0i0ZPlphg
q2UHw+z0/550s5sHr36de+5wh8lc6RWJD/Liq6ttAlcnhkoGOpRW2WbS6KpV
UjXB7qVRjcRW8iWEyv+5qL5O5ljYLhIRQ92i4EPtr4+VQ0+AD9hb6SEWzyfQ
WqDEU2w31+1HR3n9cDV7WxtlbIieBB3yJHneqYI0waZztJ7GBRyPc5sMbuTp
uUFGW/Pd1IhZFM6zDITYJYsB2ORSPC8vOUIpNnyvBvw5l7X6RLhJHpl2Y3YM
piN4U3KKELTxv9moehCES2vCFSFfDZdGR/IucGi4Vmegekl/ZAhMmcZHBQCe
qJ0kZxCgZIUiwC16Yaagk4E+UmEMaBOTgHaKIYlLSS3JFdFYg0L67x3+q3D5
H1JL+m/+1OCQpxXkBgQGzWtAzXcMjuNSqXk5Sq+VIRfX3R4Pqdi7YImzuUcX
dsNJFpMT0Jo9RuP/X77beRM7zoZ3nMLns2cu+ZzF9KTXdLdYdhEiezno3Oy3
miA/iSIYZK76PPZ2UtDCMwq59cfbVesbrJwx//aqM94eS0x9gJ1zhRpcOZ4R
ahwLoKqoSPxgYhniDHZC+Bp/nl4vwqeQSQkxshjc8ja4sQr7vdxzWzmLpaLG
XPVD+PsNKsYn+gYphTeqIls+lMJ77TuY3CCQ7ejdqd9lX7Nryn+h2X5YJ9VW
cghZZDzkpY/zabhweyNMkbA7jvCkaQOxw0+NfzpWgBmfzsS7ZbZ+UHBb6TSk
w18xF4CI8EWvwuWLPqVw6qmuleT8y1Y4aIiTRoPSWH9aDLBRi2di8DcrkFfd
WzaF+wMs7vSoUClUn8wW8EM6R+1fAN8EW0Liz9DY/KqLTOctP7r8VHQ31G4F
Vs9HxJPMYwbUmxVp8mSI8wAYNwRZ4iNGCs085JPSfNBQ9uQ2GuJE3eLdKhh4
nEdWB28kZCECCpZrN0/PhXytA4eCV1Q/zW1WGVm1l5C7ObcHxJMarr+0D0rp
srn+5jfgI28RXVl/d8m5/NNyq0Tu5jxHad2sDasw9HgUhvXH/wcwdCJAfNls
pUbXy2Zq4Bc1ZSbIUYqUS1c+4Qe8NUFhHe336E6UBsvoWP/G0H4OONLo3eaU
G2pLf/n0gS8haHq0nnaZp1V7nt8QzVc53nK6z0FHP96dUHH9M2kyESZhy19K
nDUohCO4MD3l+PCenktZSCDZ6e85DOQSA5ZJsldtRLaxeopdOA7ms9EyTIye
rpqLlGw554B5Qa9bOGA8M8Ltb70DMvyQBX+RRaYKvj20UTixni4C4x5ptBTn
ZLktbxd5dWT5efwDA9CwI3+r6UUefhmoS9i2NoU7eODIv3Ez/+4UCf3/sGEi
6q0EJZXcP/20o7FLOq4ZOfB2IQ0Bl3ovpkn67RtzGXXWHoLv+0vu8i8+/ZOm
noVUOB10jg5zdiygqJef2RdykbVVw2NRLKM9Oq3QuqSiK1LHySZqceOgCnGy
uBObR5b0nJq3yh7vbJZS2hu5Xx0oBx1Xn4X9ti51mTIrB/oIIOxeST2va9Dm
3JkLO/iORah1RIP4Y8rnAiBbQZVWYF4LOkQpI0OyK0UMnhDzE+s+aIp8bZHH
muF+c2o+6IhP4LO/aQVxetyEZQvslkemZb/EiD8lDlkIqgOI5R9yxcxSMizj
PmraD47yxBxZXLHGiL9x3gPFPEs7/NfpRk6kNlE6Sd8ZRYtbSrWOCIoaWhd8
ZQm1MXCJ1OP/gEYAqKfYVLqUcbrJZtNf0o6KDQ6PH9aZYWszushBEu0SS+y+
YaRXQmkqKLM70fpZsISFjfzWK/+I9FUgyOjvZs43/R8mGvycGK6JOFuoKuKe
R/xMxnqxjTBX++Z5RnzOeeUdmXGhj5YA4Hx0HEDKk5hHApDFEhRNlDWd7McE
ftDQMnsL35hMjBx2/YBng/0K5tdpBG1RN4z86ohORvKwGJBrVbOARZ052FxS
cSRL49wzGrB3GKJ5pkL09+eMnPfbUqVuVuK57+ES32lWn8yz4cLuco5SHrit
LnndlWpEBx7wfOK9b9SICwX3bFM5OPKAtLuRF9CkWxaAV8q1LuHGomh16ir4
LWnpV3o8PhIURq4isqDKo+EniBBLLZrVn67sOxHe2nZNT9WWkbCvERA5rkJo
BSeCK/egwJWq7AA+qYKMunLQDb4J3ACLk1i/U+kP41OO8TOXwl80dX+D+UMs
ZTO/j3TlOJJ6JEI+whh8oDazWvYdH3vklLGYfSNK/DqfX/ERX9R69DE79qNJ
IhTTi9sgP38ZeK1uo5bldjYIzr2szhqLfmKu3gsBTJJUf9yJRLDRf0AGrd7b
+0MN0PtmUEQ+VAEW8XdaM7s6xULOVn0GApjSADpTaf89N9XDECppET1si5gA
nwP3Q3CrsrcK+2oGQs20Aj9W2mWCM3rvtfLZwb8On2ftLVBvY/L67Ew4a53+
e+GoC5Oi7t5iOPUK/HZauxtCGd07HQ10eT73VmblEsmebPyxHv0qgEDJ7xW/
J1iSfKyhEf0Q1+RUVeYuo4av4zHFPLJwvf/kXkA+rGQxd/k3OtcC7AwctoUn
dd+/ZcmZbqZ3autENCa/ts91AQlFUIrUt5hDENUmBTYdBlOvOqM7nSTX2iw2
8Lxc9W+VbRgC2iExVlr5Wmz2vNsMIqLN5Ao/82T9CV0oY/xgrpMcCQ7zWdKt
/zOeoq/oURbdE26pNOGhDxC6zd2OSCkH5BdnFl7u48PQXFsrMNCBlbxuARCq
j8VXQoKyAS7ROJArBUKfH5zFKuP3lucWdwgC5kdBDXxDp644vYhypqdIvJyc
72N+/BFhPKe4d+l+zbVj0RYcdKnLJ6tLuT/srAADBJseduH5p8J0Q7tfuw26
noQFaDi/AsU2D5ts9Ocn1PMnZCV1UBIivPy2jSzaUADL94Dkw7nLARBLy1DP
MMbQAqWjBR/qsCo555cOEyjbJZvOQrhcnREewIOMo8PO6HtthW4+ycHYvvN/
vv8nDmSqcUxHCOyIM1pRkupZQo41+ZsXfuw41FDT8OpOJCvxlnNbi9arsLOv
7gPgsGRlhwjeTVqkd2Co10/g0WylIIyvo9yzLdutapKACbwZDoUzqgNWbw7W
1AcQ8Sq29r9BPrHzDwCSlxqn8SMnPMhEXrUQ4uMqQQb4CUzF3ssVx4uGWWrx
AVnwTTVLBYLpfVNI6++ce+uzwkoZb4nHDUNTxopolFhOSyz8e9gMUoX4c4k8
pxUqjuRpUzAlTF3udUTfYb+7YCpw4tD6ywPS8HLXNs6iWjLyp8cOGay0Pvu1
/W53ruoYZvJbYzLWyR87W/Yk8L3XSaAwaTFTSyE7v6pJ62giVDFLMzdxcuG4
pQvPiRetCNhQkc/5KEV0dW8MAppSScJnrkQ4ZttwGFlJIPhQtvVAYmQZ28qn
NqgITmyyi+kPZnp5kjke+K4REYu0+r/sFxdMwhAkVQV6HAzXX/LjHRwzjXSc
mlG99tm17OpixDZVxY3j7SOTjz9F7x2SPCymiFNU86QTdpJKw6EYAWfcfHGX
GH5Ci73qQC2JmaAqhG1c4+ICSy7oiuG7KhWKQ9kHk6inW88TkmkxAhH87GqX
rBn+tfKd/Iqwjbc0hLLrNrhG6UIYyP+9GszFla8gnxgCU4eo8TIy3Xq+O6VY
5jQNEhR+C57gIV+0zJqBkhLvdgkh3K1Q+JrRsvIPCX38XMDCEG1RakwuW2Sy
Rxmpyh1W1kQ3ovFMm8WKgG5fYoq06U6NxlXegm8wc9RuWtfcj4pDtfKB0Csd
BPXPnSsLYhq6/H9uPiuRVz0P36Mbsci9INwat2RroOnSZWfnO8e/QgJHBEW1
Dfm+FsSV631teqgOYgqgbRW/NgQp1MPYsmanuoOEc44dwFLSmmtu+jhowrsH
B78kJ3erkCujFk6AJC27GX7Vxzzw+iIjNC/FPyFb9YPzUym+5XBaqzCqd4E/
RLLsa9DjBBAZRZwqwmsHDKaCC3WkpO4OMBoKD1EHS0K5BQwajp+Yon7yOVLP
vmW4pmM/9buHAOQye+/kPKeSdQoCTSCnKvUGzHF+i0PVNj+f01VqLgczLsWw
NjC6vvWf70oal7Ju9FCNMolyw5fRyniJYC+2t+BQPSZhpNrcaPoJh9eJXsuh
shefRXKaYb7wzhW0D5cV84qqHl9NYIJuariSNw0YrCE9sBOEfgHVOFbvOu31
aGjD5pFApRQY62yedaGaqrCPuVUWK8WveENodnJCd+SpArXBBMr3ULLFiUSb
YP3U0PPD9yTpT0LH7XYhrKgnXztDZOHEZXepoilUB2P4VD8AvvuQ9F2KTTye
DDeYe7oV+JB9KCm61QMiSaMEqVZm6T92tPBZWpbJIwC4QWCTlKXoRKt7KzBA
jXYEYxw+oI0NT1D79oSzlGdXDbE55raOJl09yx/kif0ouS+lfg7ZRZklpHY4
5A6Yj/kJZpHE2PS6LUQzObM/KuuFtVa5d/iogGr+JptTRbFIIzsIh1CXc//a
WADKWtZJJl61agQQqP8NWJYxIBd8shGB2bk0RN7sNEsCNQKaHqHvV01dxRZG
liGG8zX8GX9f8V1J7RviZRMp1iLlmxGHC/Hr5zTdMMpoC9cff7A2C9Govfz3
K+uOQJd/B7+SlxhB0E0lrIUe4dlRHwhiWBdkIYGl5cQqKuLoSF3mJdbpjHbN
GSUevMr+FXv5vmLY4dbo4sqaaE1UrLuU45jEaujMjrwj4nJz93z/0HNurNwF
5RHnBSqYlfX5t2B8IX+kI9+kZzycfX5itVv9bxh2/hs+O9DtUl3T0+Dejm9u
zzgAMC/Pqvz4HCYjgXFdi62gVxW52PcjGcBsWc+qdxwYtzr4+0UTbi9kahYW
ICBYyP0rpl99+VrEE61G+wDzn9pqgBBmxvQTcQN+akHpPO8iAtWpIsc9eM7V
uiLnBx/t5Ms1lWu7RwB48SGbsR5w29X1IRmnuk0EFCsbl2bAeJVxusHNVePy
d1bNtKMZyDGF3MY/JMQRJVY58BMm0O4YNJB2vdkx6AAziBAfko0mYVuT8CDv
/jcvkdIlys0HJM87AIZp1Xq1ZdoTr6Z2H56/yYNlPg8NrORK/mHZDeuSpibU
U9XF4PNrtRO8A0PyUESBRTpgLILsTEk1nUKJHNL9X1peRsc2BB+0nODMRFXj
1SNRV9C+jBYUTuZS0QF6g3IZQGv6GMvmhjpEHa8RXx6MyBZ9LEDBdxlInBkX
fDDbIXZebBso2dziCR9JqezZ08FqkXdOW6goLFRNmQua2JFaNHIJ+AfyI8R4
IG+bSMuE6JpMj4tChwM4TWO/Dm+c3IQN4YQqx1nI8Fa1iUW87DsSZonMZBKA
VEBUhpJJTBt95YlnnzjciRbak9Se0CuV336Cfe77uqy3rwu0OEQVPuKSbD8+
ppafTh9TLfzJtJ8tPpK6HXb4E6osGerwf+rt6mqOFY/uSqH2scQIB9NxQ6vF
0ZLfIlmeqvEewrxCui4XU3xQaubnmLj1v4Bo5mqhsoAsNTCJKbC0agf4Ff3Y
NoX1LzPkZsCwvxRMLhqdKVCU5mBhloekll7glin2TXJjIUnv7xJy5iABUGeT
+1L1kEIQlPLwh83ht/10Bu2ge90EYe0YXVQLPBwGR3X14y+vzhv6vZujvU7P
1ihDkH9ReKuy5sW+5IA2vn2B8NF2dmHuVxTsMeSuOBzgzelvH9ylf67igxDG
9jk78YkUAVHeFPG5DAK2kQSSjkfWI+7x5txqz5xm2+r2l/bzTw38Eb8v+8dT
pntI8bwc9Y5WVLdnDgXwS8nAh9d/D6mEMzkivCUr60eEpwi+yVuY1yjsjAIy
6U/BbudS5sAhsS4SGw4ZS/602B4Qi5w0FASzDH0MvfpUXptx2Eba0jrKoOi8
ZM33kfDLdDZZ458J6pnpKvEFV+Oczvff4wtqCWV9vFtrxd2OvPCKJ8g0vr9P
cLszK2sGA63VJXwiPn0g4r8XyVxnF2Zss1pCvlxoXcLhQ2amq2UxCp6dZe18
qbLGFch6AEeCfd6YfoMwQbfXKMZoe8PdFmptg7KXSUBjeGaWjS+qpJWj71nT
GgWei/1vUCJNIYBP4eHVVuu+pSuQc78vjrkkymTCpaRhd08WpkqiV98VbKiQ
HEzQ3zZw2LKJfQKw4GSHieVQCp9EfEzwlhSSmyKVk8THjwruc/41C+IOj1xC
SPRHedZzekIk1WfU+txGd8RDHSYc0L/4aEdTRJuSl8vz6R7nZph82pHwT6XJ
ezveIKcGBDqSWrzWRWFzXTsw/xV5f86XmJPmYYA0+uNd4ReFKjqzAkgpJQLP
V/ZmdONPCoeVsYm9+IHhHCxTKDt0uLZ5/Eu3rCNAZZsPSnlWiHhujOdBBWy7
tQNbRzBCh9XRxnfvC5V8pE0XTbKrQgpo9d6IvLP+HRlHYrecwvP2w07sucg6
AF1kF9B0y8PZ3lKpuB7MxtYdHd1UqD4c8z59eBnTfGyfGG3pK/J9nF6s5ZFa
cU8cTHNIhJ21jMbes7vq9e7k9w6BfH0P9YBaZCec/Qz12uYqy3OPd/nyiXB+
+Jq+ghuE4OmmxpGP5U3hkPDlWp5B0FMJ2ZCDWKIp7LWQePxvEMIVUP9lWyLA
Ph2mVgiORqMWDS0vyZumbAujDUGTP2GRdgnWrRs5O/RMjqCbE/V71apd4li+
xSBSFImlmkXhOzRh8qt9AiZp48MRRpYLnDEIcRvTnTpOpB3Skh5YOpEkMx/5
qcp7NKjH+0dePoLmZRAh7f6ICtqqfSBKVXLhiRjRWiY1TOMVg6og1ZP8Akbx
2BROgGv90Qy69uRKJ7zwKvriNHFu7cW2GnSV8fyPDR+Wkt84oMw8x4ZJF61i
eCBJDDO57ZI/Yxk88xLkjl2pTuukFgjEcC2hLse0KWKOTQTe2lEW58jpIQE+
FtvibAqfORf6EZWotUNadmrMK6GFRwlAB4pYXHoVhc32H0ifXB2x1SmJyF51
s8LIVfW3BLOqWcI+5D3hTgXrihJodT6n1nSD7cZ2iNKh0OwDBLW4druxPxrS
YJAsHvlI5UlU0ecoH5odHu9vzR0svLtTdDoR5wrpSS0pC/jqd+zSTpmddVrE
JhfAM97Nzm7ZHnWTRBGRKeqm4qV1nz75sNNQ+IjZO4+LCL9WEAJYs/opAQa9
xiyoerudwYsqAv3GLONl7aGH2aAJ1AYSefxFoU8QGth2+nVwvq+yZ69LKVgD
nY4HlikNQ+GT1+EGbr8wtdXPgNufKyuSoui5NStCoN2HI5uLXIDuL1NWZ3u8
D1Xyth925vaMvjOSncfbVxC5jHDje+2GYJ/ybSqB815ybKrZ2z0R+LxGWfwk
c1FP8q0+L37GRwa/i2Vk/CJwk3yicnCIXcqt7UfyeRcE54g0DkEDIP23OcPN
pL8/CJlJOyZvu/5Pl3DUavZsw5kACqw8IJUuXddIvbSMpQujkio41oPLm5xZ
t7mZSpgf0j42i3+N5VUdU/o7+mytv+MsvOoJ2Moh7QKKx1VKal+z3isxhagM
hbiNWVSCkIpr6vVCX6T2ABei23sfEAbrFU/twSC5mpeUMg2uK6HbunZqKISH
f6pcVhw2Ty0wVSy4xGBJC/JMss81eL9rCCIv92XeCwo7nzvga+cZuEZMS2PK
pZ0NWy3snsroHVXuigS6bazkZ3S62KK66Usxx5iUisvY+StwnbuxF3C4fepW
9SnnzRxn26C8gBTV+7uECEeAaHu5GRGpU5iFPoRmsyYR8XU9iiGYKrhbis3N
Gb72J4x82PvNV7nRsz8eSNlHOG80y5xtiwInJCpQv82OD8ys6ZGscZwh2Hb9
yl/AL74pv+oCc18S5MXzVmKEajOdHI87w/oSUTl6IIA8ON7skbzD8Ilg7gja
AY5NUc2J6S4JgiJkeMffJAnprWIuhZ7O40AgUY7NdJ7SEt2RX3J5Igul1ill
HCDv6pf5SWmbxqVFuxcmr5QwaVxuINo6KGSQhfJSvXHfbkXrYLf/rUjG+kzp
5gSYh0STxzJoKx+8/B6mJhmCyKbItZ/R25veJVutJIBgQE6fFaMUgFgx4Efq
eBsuL8jBpUS+vDmB7XeTmDSeCD00e7tD6QQkIV5WccF+M4bv/sX0zke0DO+U
5In9eBGtUtkRXkGzLHdJ6pwGUyzcuFOgmB/owYI6Kyp6UC9KUTANeViGlhtX
Kn3+ckvAlQC8mz8nExztyx21CXNceUy8QNbN5khxyjvbsLIZDYmo6BFunSfK
AiydAvX2peO51tiUtGJrrcAF1VQDxa+VovnQ/kZ8ukpQN/LqYfReGUKJSjNc
hcNRJ73JEWE3CP9qxFIawqdolrz1OsUaU3V+H1w/x5Zm+P+yCNducvL8IpsZ
1X63BQxBI+FdMFZHuk1qulwsbALUFdSumVlj3dkeuoesKWLOavmZIXFrpyjn
1ZhSjwjAY/MtnTnvCcZRRyrjiRXU17LBIRPkkvtjaBevInfhvBc5cvGl4dr9
Xb38PzO1rG6BVGszj1j/rJMZEZAWmHxpod5l7ds7pb+lzl/vZWmZ2JhvNZwD
C2vs1gBINp9qyMsBtcHj9GjGSVdHWXmUyAkPEpBsIYUdDjjYtecbDFgCrDD/
ou4SKauZwgM2Rvqe526gouxv4kDRHnsLIxV+D6x53L1Pl8VSceBF+ixLLTjW
rmhRwz4NcGjV/xDhAbuCrGrObAHIOj6igPQwCaO20m5kKs/+cTEzcxHH7cAO
M0FfazCdcyXvApD4fNCG190Dpkc7tRJi85ccL8Q8gBpaFjb00RymPeZzauQH
tz8udJyEeXPh3FOCEDxQLvRETr7K0l1Rt/Ql17Yp8pJdopPuGNAAHshfCbCX
kHN/wMvNdCBmbYNO1hylGJHEpmfAuFZOo1aOThOXootDANVXcNeusxJNqhrQ
+ku/MRBiFfDoqP3xiIr3zRrK8vlu9AvNEYzt9koG2/wTPn4Oo8Jl9tJHXiN4
GiCz4IZ99M13z82D/nnex1o3O8waHAmvRDcO1t3WpD4/1uxNNw8y2uZrRpoC
6AV6NeL4NfR5cOA1K8d0kO1MyXeESYmWx/M3FlWnlxY7mDBykTtz954ipeQn
9SLkKZNNMXuQk+a7CaMLCc2uWW/0vNm8BtMPYKDaO5iGjUH32sjcbCVAimVQ
wSwVIKELr5vLtcywHn7jBZN2A4FrBpI20iqzoUgxX0zy57X01gF0j/xAs2Ms
BgU3UKt0oZfKhMcVg6aQEvzgqIsp22lYOtJrlhlIFH2kLdMMlKyPB/J1ZtLk
UA3xPMFi+8SmZKDBh0aK/tuwnK7+CG24LeX8ldG1mvVXWUhGy6+VOPxmDaHE
XR6m8zVsmelJ9EC0Fm31Is9QRz/y502QZCQlZKQgOBogOf645A+oOeSppntW
WOjno9oDU1mM4Ek9/hApdvckWWeGi0I6Wa1AqDS66PodSSofB3BrX+kVasDz
5JM3IwxvWi2wNOI8KctUg+l9E5vEl2qAyucjiOid4NOGhK8g2v1Jvcz1I3lr
CHe/OqExTFesVi9++3XU747X9bJQeZqqLqEiIxfe0Ykk8lOU2C2Ez36+rmPD
n48WKAgz4ZL783t7n/3KuhI5Jj1ywe9u9a80Z5K5uExEAx52BnqGcjZl/Tfi
VWAh6tTB3eMHpPKi5nsPQI+h5LhrVfam5k4rfNnSxTbF0MswqXJ/DAR8X+KX
4OxuKf+rQBhQnqmOkJOMOL19KIUlR9nf46q/WCoYKz6WO3a+nVY0xnbxxPB2
0Xho/s6JOFDK8D6v02l4aJTC1xqosJ2T1Fvw3+hnXgE0aBhavPg5KzoyPEdy
HCtHlfUtNedj6id3Naq7Ll6vd30UXsJyb55WgcnV2xTcbodflo2Gs5gRmP6g
AgkWMYVuzs84m5fQRKZnQrAZj0yA3mTafq2m2OoX6HAW8CRwWnPGLRi/iC2F
kVIh7XiAgyN3KwjhuqC6U9lCNoesdir9V2ieK5GpMDtqOWZ1F/CZ91y5A4q/
V8lpvoJCV/RK4BIpsNvnhyNJJcmAqAXtMKPJV9SXO8lueY6LoZcN+z5JELtF
WlIlz2x9xg5nxKMdyrY9VJr+I3lamPAnT2gF1NVVM+PYKFvRnPU0OCH10C0u
GzvRPCtL2wpIqCxM+wR6os00x2FgJTzTe88fUn4UVcUCDJgo9lpVFsQ4EcaM
JjZNCd0G7/hAYaK1x8rgTUK8C4dkjDx5whWwCR4QJem7KcGYXaBdrDD9Q5Zj
crYrVYL5cjp/T0QquC0yq5fHVrlZb8YMOgtIOrpo2wAvn5IMwou/YIdsTLQC
tLOsRN/m/DofDJ7GeUb4xjhmcm18cfzj7FWeXU+j7c1bKZcpKKs68PPCpZXF
0dMRk/baZOU7uBSffiIuMMhfmslsH8UkpfwN8VKgd1v9bbOR3tbaedHmhRyi
WU0eAh+HEjymKIkCu1q5YZcBKPsaDHqhgbda548Vs2IU+8OtAIJdQ6DKyr3U
9TxAmI8U0aUvAi/G8tn2dBB9bqkNTi6bUVTlscek8Vl9BMzA28ee/HVIy3f4
YEBRfq06wzd3t+MzgDYu98ODJH/wcERaj+Cpr5RYGBiZzX1UKD8x8g1QvNOr
DA5VC6OLbx0TZdgOVGnMdwGS0SduEffkzqPoQSQg9ULwaGqAeo3w65C0rkEG
LysXP7NzWzveIXh/gXvKyReIF69DQiGxX7TveBWKR1ymvn7mKplIYbpQ8OjK
sJdn36lTpCEfRPEpprpltLGhQwgK8t1WB5/YI1xpbXPYyE0fBDTcAtPbGuYe
gbHbthxiuQ5M/pJyhvyfqkrlW3TvLrGGhnFdh0GdA8ZLU8KSbDf37VOGEw/y
lbj18BBKnWjA8TjH1YuO+894G2hy58JuyvSSeK6zNo8ImVyC0rI2NGXW0+rS
NdhSH/HApEVQ7jrd3dd8lYlYBlPfZvPrvODvLOtLVnEqvvqZkyVlTVWqnJgq
vkk0vMqLCFr3duURw003FjEVwaIUqW29QcKSB4p7d5EMwE1fHZ/h8ziKRImB
HKqCxiBaytuzzALXdCdO5rlqyOY413+bwIdcdzCqknyF/SKBHj/CPe/TzjTs
pc/aXwGoenVC8FRwhviwjC80nZzM7rLGq4LAhhgYQxi2eKGIHUxQi8ZS7crx
G23hka9ChzwBSmZk2dogckJ24KiU7ssXXuqp2Cu+Y52vYQS0vG6uDW2FxWGP
IoSCHEwYOQk4IGLuT8c9O+txr4ASJ6YQDqOfLEr7sHTkfHIzR4OXS9fisydB
mekIyZ76nCINV+cUdXfRIzUalYqCNrp68zkiHvbTUPAVQ3qXP6/1X2HtCSNc
2E1fjRCp95hx5gmhzqVmuWDXq4vIL3s3vbEO/x/vxuhLTnjZAp99vl9UA5d0
QDDfakTCd1pXjne3iSBwy2mJ8OzmQVqT+HCXXSPVGJNI+8iWr8HghwEnrdXL
5KdqmMpwXF3Ey7hCBxu3fZjVzY227DSc+KFOhLfoOclYzkG2hOIHD3n0wgpH
nHS3KjLavMOO9+VAmpyx4mt3+ONsvbGCu3l0AWCv553YSuT6xTmGmYemrRIR
MUFoE1Z9tYCHmn0e97owGCCt62s/Oxf2zhoYiNWDbSAuIC6pRqMhfsNQe6FV
hx7XRthW1gClgYCk7iUwvlGPpUsMIq9rYpL/3C3X4q7VsxTwlmzGIGqPSai8
3FaX8ukfTxVap7nLiOwYxtACi2oU6KjhMtr/OV8P4HRpTFj0zGIyxrLX+ZIp
bWreJA6NJYQcSuwm2ri6LruFvYZMul/DQSrJcFod+u+EA5V+j1HqUs72we4i
Tgr6svIsHahklhqL4DpiMAbniPFOJLpBnYUzyQOzbbUT1eswFPew3nnEpYGv
IL5zKHcT1W1I2j3VO8f0W0Zwf3HdaVGjDE4vyQHtAo94mRixWEYqLDj98dSd
/4p9Ufp+VAcZvpxZqxxoPK9DfcRf6uGUZj9MALNdvABMvWEVzKSG4iLBQ+ns
ik9pVcHy+7M2yXZMAaoUkr66pk6iyhbYAwjrlc4n1XTUprBZ6XRaHBPTLlYa
hcfBa5vAih2EAWBcVlpmyJxjwRkrFGvDtGHPw2//MZAlmgRpcPo4NRwYFuDO
XJSrG/CN35oAFUY4dKqbrjBmKPSdCnV+faSL+YULUPrwlSom9D7YkkCZwtYF
b3QxGIIz2bM3669qlqJiaICXD5A9zG7usEJF/aID7wJj+o+oI29iMfGIKuWC
21p23zvHA2XNyngCqAcMTYzsthi8tWjNreanDuVManvshpZxmGXSduOZcN0p
oI5TtvOakRN3O0fl3H0pHtCIzLwy6uKuFPFAO30gwrM98N3wQlUSaEEBbjAs
W0M8pkPUzKqhj4FEkgfZgxWYbBUoSwMkGEAreQtLMsRxEqBtyzA3ZcH+I7QE
qeEtbntvPmKG8vHfZjTrlqh+1tJBomnz9sQgXlXA0O967HzaAT79RcL+JFON
BL3+UW41cCuDEv8rQvubuEcCHXOp9w+y2+Pklk2ckeelL1B0VJpPEnscKL+T
LaiMgw+kNUJgI/2ucmEBs0RLwa5q8xwc1YVQHclAjYoHg15lKXK9nbBUnyBD
X5erIZkcnfRy8lAFg08sUqsSBWa34KsCGL94er8kWWdgZ285PxXIoNqTQksu
ctM1RVSeh5YKn38Iab78BY6v/VuyjwRisz6z25yFMExJ1K/3lwuabqjgvvvR
/fAPLS5KXbL2mX8RVlLi07/upj2ubqD/0o+lcT0rFtE8CBmXgSQwgJuLm+BC
lP1CXWNR/o8wnY2i6c3EO7JCBLtapOwfEvpMGlrSacsV6LD06pk+9B4kFEgo
8ZU/OxYRkFbZ8pKAjeHRkDQq+5FaeSnw8RbVYKGSmw+QfhXw/FZ1VLyPGIQD
VNHxnxm1WoGrokBHQg7spf0Lf1S2JSc3zittVhCPWudqwqvBgqlXe8EyLuUe
X7P8/gF3ynuqqNTT6QqJo/UpecFHLnjCx4SUKRpXxE6cKwFJTyiXIjCGDOkx
Vbs+Qr49eZV15tChZCmkuthpCf9qB8VAjMOKmRm93vxiXSs3ov44xk0LbQ4y
PbLjxlbhoHBwv/Qka+Im1i/ELLUuB1s0enrweGs0lcMq9Ji1N2Zi+x3wE/rU
8yYWm/9k4pbR3g7drHqj+lIxfZDlq6H2gFU44YsfCRrxmP1kndN86AEfYyqA
SCaoYX7AcyP00UmLmrT3vNjmPVT7f1JffkaDYjq+jfCwXx2/qPGmLbALryqh
WI2ny0zGd7ol5z7Rdm/6t7NBYQ/CXLR6t7I/SuBzPkTF8o7EzZgylBwaLt2L
prmk0rRaUCodR+PevQJmlc+i1uvamRKdYzT4V8o2K76Nkp166igAtB8RckcZ
LWo7I/z9HJDZ6Fw4bHoTcTxGywNEtIpghRCCvVrvK6vmD0kFV5F9bhHH32Tn
UxHyzownB8xQhZvNtbV0N2aXwzJ2dz8i2O4eU+F0yGGzbU6QbKsNxR+00WIX
jrYlcv9bcmoAeN9dnyQuq5R5AM18lZIGIDSJwGNXeQ+rLYAToBxfcE4dArU9
q9TCobLBoPMgtoDmfwb2DTdWqeo5yqMBuQ3a8SezETvxdzytsYHkl6xx5MCQ
mOuN1nRpAFZ10Nl3pmwYavfMrtTK+gEvqIqKvm/HtfshGlaxEUmGZtlRPL6F
X08j8p1LvnzMHPxknUDQS5nrluYtIsE1UFT6xWk8K/gRfmZWPrUWXXAGybXs
IxTwzqd+6SZy56qa1YpAIfS7+0dfC4yhDYMjcMS451cFSAQXTwATPu2SaRe4
kKE2SER3eYhaSUNZqTb7wG503MsFiJnLRGrE7FJ/rmi8OtuJR5MxUZOrrf3r
1dHgSgQQLq/PJCMlUAPe2ssGSH26+39+V7/rwMmkt8hkhu+jvi3DzZvKKaMV
4aIDWJ4TQpUwe3aYoSXZf7OTJXNgaJbDUQ7AqfQmraw+boqVEbM43d3yaQaS
6zYzT6dOCGSa+fnU91PSZfLleg0lvJLoTlihbLWwsE0ouoRsxjs2nr8Tv9qB
RdAfYdRT+hHFrLS4/QnZhraLeDjTBTtdDcM/h8rFK0VKdFS7QAydfPUR7JI8
Se2AjAA2DIKLsDCVIsRQ0OdzU2tI02szG5zW6fzCDN4QTOUUp/YxYunR81v6
Zc4BWV7GjD2RjBTB0idB1HAHcbzPI0Dhvp197R2NRKoKb86r+CeP5djFeL1C
JXxDAjI6enhw3mQ+n8js2qbZNKYH/56ytL+UfX6s86R5MKlKruPOvFetRFY/
SwcTm5IB0HgYMxIn+63ZX6syGsfvNCmWnJ59bYZCcM4pPLxjsMs3lSt8ueZJ
gWa12ZZ0TnCQ2Lr6LjdkMH3pp8C9KXD5Nmkqm3LADYDFqAS8jrNeuqU+/7Li
YI7wGkqY7ewkd6N7did1hfhV3AgmabkVhw6MuaD0yDkpm1fMsv1HuLyq9Ncg
EwTaPMNGeRnk8q7KF5zZexleLdWdA/EQqKiwVkkQIRR70JrccFV0HsHyEA/G
1sHqGzPgpo8JkefPDT4Ol0KsOHqCvBUXyuexxHpL5SBeZzNCEqKbCiQL0sVS
ZqU/x+pu4PZN6CQVtj3il5O+Nh8fkX8c2Te6N7v/AJYBIxkqw6JRVOw3vlYQ
NdiExXHTlGJ2iNK7vIoFsQpt+EIK7PqMWBzwLlXHlkzd59kqkKiKxm8VOUDt
UHZ29znIJW51ArEXdf4W76tdsbWwQznnGsrE50CbUX8txjMgpnWvqVWZl9oc
EROmVCLVyOo+rkJBa8stICCPsMXHWT1+BfB9dMEzhLRVpAr3yUbcLnYUkZJl
D2BEBC1SeDW0oAjUhJUdZgetwoPqEVb2cNaAChTvNdTqabQZR4631blZ+sMr
OB0jNI+388qj2WcK9uHqACHuerLdWCVTEsOFvYqYP4c63eQ4sb1TM4QUilZR
ZbWbBQK/GjHuYGhd5wW1Yl91c1mN6VVP7WzSWPy6Mfl8vuxn7f4Uha4cFd2U
0ca1CtYL6EBKu7z4+HpU/8r2cw1pTFOTrofyVv2aAOlebaQbZjLZLqT2+TC7
WxDfSimikX6aA+LKnmlDhXtJaxiLJUsDnbIl6EnTn82kxl2GRRmjBFBDVGRW
DPZoVU+Nj2JRIlwlLyhmY9kOvGmefgizGBAFk1enYtCH5OYvYbc+3EKBSIAJ
WOMyRk5LrgG/mOPooKiF9ZQPOx2RLabxzsUGBvKIjIEH8lu7OYc7bCV6NjB5
1csTAT5wTTgthrguN+6Dj1irc2WrPghGrRX1UsYx6Fh+3Xp/XMLfKb/f4sO6
+3j5nbtVDU4C3f4lCTI8E837948ZcAA0qZVdbJk6IBr/HRW8UBMCqvKMKVGH
/uonccTwkS7rOvYv5in13y1U3fkBwb+Q3ARN5Stu7FlK6oXp7cUNMXr1bmT+
VTgultM603v6FvG8NxMhjdMtEbjySz5N5+VAxpPsOi/gCtNuVw5fhTFRpT8Y
vO6y/Jn7yaoyLfsw56E2CA/3/e/R7lkcDvaIstnqHF764kKIPOgpoWA2yBri
F/4oniWdRqQrP+JD5rFKXrrrAf6JJi/lu1FU2soJ/bJ+wg4ttppdPqb66Jt8
3GMhC6kgEnJHR7wO3B40CpCW9UTvWza6xO60jTtg81AC1mGcBGsKS8avm85s
qEbaeo6Ofij9EtiAGM9Ek/Adk2BAx82PTPvWtzn8RADKgQqmWZ33FYvKXw8g
j8psRxdbpU4haz0uvP+IHzUB044EPb/52O7/ce1K8RvAlSSjO+VtA0gXmZJZ
8Xw6608A+zxoSunWOaxB/3X8PRN4Ul6dpQbw9PxRkHG0mBE483+2QhjDQWUu
zLAHavFeezg6A+zUxWIxenbsyV0kLxzL5ZmL+mpITYawHP8GxDP6/Cwnuu8i
xWHdOy7ynH55D+8AsrzQ6iS79TzTquIF+vcsJ+Ugrpr2s6g+vFS0jHcT3sA0
1AqWkb1EaT+3NzM/SArlVCg8AfLaNMz56Bl+3YsJSO8zoT7v1I9pSPNuopvo
qo7lAv4ETPNUFo9K83ThMCM/eYcsjScqR4ATwF2wREVN0uRkKLxCOCv7Mef3
IlWZNSxDxOzKJDcmahlCqS8g7L37Wza17heDWSL9YQWuur70qA8sl02t50yi
NZsBU+g3FUzi+tp5Xv4P9g0QhQCIKVTkA/h3wo/g+NfRafkEWYXyVfOe5jFB
jFLzSOzlicK5mI1pUyjkbEkefxX4gygFjthCXQISIvhcCbC7/mcn6R8RPNei
c2x9kCrqSefRwR9tNDTDCRNvwwPZ8ioivw/iKseFzEjRWIant/jb+NCYVSAU
vNymh9mKCS39URdkS6Lg5Mifr+RoMqRihCeGerXhTX8twExuaMJUKzu5lys0
mz+beKN5GDjxwFY9IypfGBehfR1mV+ILYT9KimpeCwTap88AtcU/DBY7uMhb
9sDR6ZgelLspG3+dyp0DYEpyUTzepf/+zLP6Xr+b04Onr92p6D4WkaPuMEFf
Rxf/tqmhPKj9T++nyxjvMkW3d6RgN05KLPK4VpLGqtiYuTkX8P9pdPYhuMwT
+c66kbZq96bnofiij7sGC/DPNWHAq+0X1EchybmbF+lCxUfPY5StLzf3LH2I
adZc7HCWwYlHMObPKfX3H+RC9gSRR/XRH2dnWyoyX6hKIkZd1F+bYa08OylM
rpFcFcneOyACXM+t0ZBUebAbO1ibuOxEhEuY/14eUMJUInUsbiECe54s8huS
OvBd9CjJ4a8ERINxgWM0NS4UU5CK5rodOFk40h5ebVnND/YF10Ex9mLXF4Nz
lc86QSmdpbIjWkBcpg4HIfgg0irJsfxJUqDNK7w9CZavkKX7H3Zz0lzshzBH
LkVvgKuDevFoXce2TTmppLE4ggnbGbmXI0+oX4ic1efC/4mVdrSzhGShA1Km
zRuaVwm9onZdNRN64EgrQ9SA9J4QH4IRZ+AIr7n1vq7iTkcoPBClzOubpte/
vLYQrMBYDUn9UQ4OKlT+ANNWFekp+qU8d30Mvb2dWA9QHekviXD+F2rNBC9u
whkOIr3QpcqfLVEAfhEpl1At6DCWCgQjR3iO67hVMQATO2zi0V7265qsM//z
9XAp2mlExAtgScgvlUyckiKqBsILab+uZHVj4FOPbVsY5VSc9vKlYSJcB5Yc
kN4K1no9ZyCwd6ttiCmXsSHFO3TnHD09+wRsTWRp4WC0VEN+RBHchQLf90IR
TK9vwGnzz+HWemXC2y1upX26B4cRm+LijlVkCNdebAzYJeAHmEHlLP8ujJbT
/S2XKRgsyTK5emM/BonoX3eO1yecj344JPZQ5jvDlrS8IPHhorPqozReEAfY
FSG4qBXQNwHfN7LdbUFVxfl1IH2UlOHJXq8VVbGd+91OrOPZl9pDfIx4WBHn
3NRJ8h8UtMv1EDSzhguwSQwa1DwKO2rM6Wdh3qGuB6RPj5n7TWQbc3opfs+7
k2XryM+9FOrjL1w5YFYI0a20K4UCvHHurtvOhrJs2Uzg3Udh6BUgNXixHXJv
FqZPjmMrn31CEbnLzFo31M369K3Ppf9/9H2j4xfEulIgWjRa3Wb53xbGXumJ
roaDJnxEHo3TRcQIJ0G/VoZzb3FCVggQDX5KKWQ75DiLQRAcM3aLeV0oEHL7
C7/PptGk07zQPWV/ns093EW8IhrdGFZqTM+1hejBB73UK00F/ylKXHbfElpL
pZS/sRN1j1baiQgJiWwmzk2JbVu2HpWhlwxkBmDtfls+XMD+jgtF9LWpLSZ3
+5xfvoPwhZnFlOriuyM811DYs5/aIXBX1yaBdIMSYaYqlNla5vbx0DRCKJ0e
Bx0Ln0REuT8JxS5GirJyiR9OKGH9NJtLRZVBmY735D6VNv0iI7hzP3MxMRrp
QBlQr82aH8hZfGmj7S+LfT5pAyWK3I1SXAeBUkjwbA082HT+EO3ptOXzuhvq
TtlzGPtDddZ/ZWuokQ7BFfqbRzoakTqN1XwyTosddDTjK3ovhfbOF9fJnAb6
4HPiI3AAV5FYWjpws4JbImu+KSew5RnzsF+N3I7zQ+o8LHpPtegwXv5HUbV9
+qURPZQZCslOAdLybH2d+9CNo6+P4cuXLHmhFbbPKuA554gHu/jMVRzCvs33
41e6pbiHySpUcaaDyrF6oPwMuYxd1+j+vZt9ce6mT9hRcul9nzZe7kYd0wkV
Jxryiy8n+6ZADDfscWdZLTje3p5pRKvIIA7beB3H5V7y1Ibw4xNY2JThoJSL
j9DsBkJqz31/uZf95arM9wTmAGLghns3q6id79eL2bVAjQuI6cVHTX/a61bN
2iBQVJpHjcEiazzLlgr57E5cfL7ZCjgqoPlQs14Vsrn5gNV4KepDgl/0ACd/
0VlSnymfFZD4R8/UirFqDyd9q3EB0LcRXJN7pJS5N1aT9hjR1aPWArwolrWs
XAg7A8wJZqght0ntfwVDz7xTKwT4nSRNzpOTNjtj2fAUmKOEctlNT1VXuUYj
ofxWm77iSwbmJu+GQOXTNc1G42V6r+ssxLmJyKKPnyNhgPHUszA4VO+uOykC
/41xqLHb9cCMd0F+RjYYAVA0Oo3itbwlmgTpOwpoLuYXXgXVQaewtbcvFI+2
Unjd5Kmn4X26wnFn9xhcVa+Hv5unYFwLagnj8Et8T+v8xpjWhvDMeLPaZAAU
pfth4eDaleQlRs3+bxwEA64pQd5ZBOq6LdU0627uKMc5caUDaTh8TOK87S66
hpz6+vcZpTrQ2/JW5VmUHsOMVmb6/OKLcREITK5BNaN2aceulq76395GigKv
CqMQS26CrE//CkIlaMd650/67nxkzrtDSCFn349tQqYR9Gves41YWtysP8Hs
sPg54VEwv+suG+qckwblUaRcK3QXCXgUGJln5hqFBU26oZccgc2Z1hNIY+rh
8v1MMVDhGCyZubJzqK0DFqJEJajEorcLZsnuSey2tCRR4LlApII+fOLwytY6
RXIl8Ku+veZ1WS7MqxLcukJblJ0ZdbI5rxdO7KFDUdIfQ3G1geGR2gly5ik0
rpfw7BTYCWx0qcdBpr5BtwvP/pW+IBKt8iAldnAENCUZUG2egS7U+hQNcppq
KTipx5JRM/yJxNrUvlH+ASAU9X610vSwBORQ+YYH/9V969jJPxiLlbZUZHxu
wc4VABgLDe11pBLIcVXwzwO59rWH7t33wmsr5df1p+yvQX5OzS5EjPNeoV0T
5/1yv2U8LvpcJ/8jj1dqA3RG6aEixzwntSlwnhUZB5TXnXq6Y1GCAqSw8T63
7Wpj7bzmX/KQTRaBy/jVnKNBcsevM3MHsolSNRhrn/9X72EFnr60roRFupj2
H1FGMeBPgNpRYLUne51HDq1Mh3cmLHnXbH18m0qBWXoq1tvjwPpFjSXlOpu0
Np45/yBs6JgAtu5YVJp9D6plZ7D+2tIhRk8BJ48E/9DyreItAVhSS9u2XaMv
ktvJ1GZkcM/+vJuh+3cNZP+3bo4+u3EgLrl1z595QWLzus0qTko5doeqzcYs
khXo+yj4LLvFiGk2sCu/XVzMsRJSbU3dX/3UlRhYWE9F3R32Eq2D3dp0+Aox
hk6p

`pragma protect end_protected
