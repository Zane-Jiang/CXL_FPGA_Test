// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aJXVL9VjlSf3eZgIboQQp/hJNbSUd6sjyZ/IVYX+BD2pQIO4HETUdfEq4jX1
9W0d3nvhL5gPvt/gxd0alyFPc+zrf6OLY+Nrrs/i2Mm/ZYD9l0p5P/fKuHlh
mEDDOTOaYYtqqZnIEjLXo65ZNKPv8CND3UoHYvzgwtkdvjnevsTU2GQzgR0e
dY/yBRvssfbdRt2eelHDnwsguNnm9rc2HItcLoGCmPnktyN3itSGHD4cKrPW
D9y0dRb8eHGs7zPR4QIBsQ+WcrRvzmt1ZQUjLJhxjoimiWakMsFB5AZX6NqE
UJNVbTolbHShFgZQm5f4t6zqa2NzAwz/Ty+bBJDNQg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kvZQ/23ptmLQ29kn1Wd7oD/a51Gq+yuMQ7uPdGyig8zp2EfV6xtydH8Zu4hD
v6vz5X8PloEeYJ2ZsLUW8R42g1Lst/0lR8gEjA4YZ71R2r60EKieLcne5vh4
D1ZT5kHAsrnQo4+5i8cj1s2Z8an8TWc65LqY5N0xLd5v580YvfzcirJTN3sn
PX6wkHoHNup2oBSq2t8m/F7dxNag3gXfTgvzba0oTn2UxOfvNr1NkYAOmDFz
HLr7k1StjVROe6IaK0kZihsDx6osu2vmD7UKS6gSN73k/8bSi7RPnu1HNOHJ
7JGIlXzeogBepq1orAxKZCJHdKHeZ9sE19qHjKpAzw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d2+oWjF7XH0o35uyyX8XBA0I0P1JWj4oZ4QG0DCRbXp0XGhsCmU16nx2LBN1
y8rmWt/amk1jZ7sQsh03ekU8XIx/k/7QvdxDOaBRKsKiSG038K3cN5K9/CBL
9HAMQBBArzuAz60A/ZZpd3vx4NwuRUoN0HG2yKoP3+myUcRZ8KRr4SrA1iD3
XrzliOoTKS3NoIxgmoY0BGjd+g4SbuolOFxdDLOCd17thNHdl5lOXphYtgmX
aTisxZwpBMpgdfIuqwLFj6VOOy11jPWoQnwuSP+Fca4ZnZpOz+uRnIlMCbgC
Z953nsYx4rx7VrEH8ip69esX7Q7qVivImThNLVMJbQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
drPdvT9YRN9IeJuJnp8KzkruVYZc8BSZ6oWYFT6aCm9wHJPL43OA1Xvqwq7O
+eFX18PV4OrxhWo/y8D00F8hR6fCXF7pTxTZZkAg8QmJYDOp7bGFTO7BTeDD
1ClbPo6hd/rn1n/nAorZNyZ1csVdNVj6jdXShj/FM1E8iy/60vA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Z6DtYB0RX/yawJl3qNtyqSrHFUujrgqVhAbFRmC+z6E7FPtgFAz7XGp4SCpV
pi/uslupDx2Z5x9UPDzZIGLQRDLALg2RKUQ4AeCMmSt2yVaFetK8punxAm5P
5At+u/Tyvf1kNIhMZ6tTL/SA5jF/QRsLyXwNo1/tt3v73jzxKvbPqaNtXw/r
hunkPTvgA9M4VELfu3pjGHhqfqki/RvTv54tqKazA0U6m/Hx3tEVDbCbk1G2
sHqxNNDgNnQmo01ZbodnsYxfoRMEhaJMiopaKUQt1kjJIxWQw47jTNe6b+TZ
S4WgnZcwp/R5t1cAl8NADIkrCAfnhH3lAC3xeXCH/PidADJDKwqHHyTCqwal
j5iUEr5t/UUH1TanI1Ycr4EqBxNZtuSZ+PIxaf8+9mmEzuZCrI64wxq4wQ+M
QMwwDstrN78PYAsXj8yy6/M1ojUEYg2vA4rdpI9xWPylzaofI0qp+ukoaxjg
SibaevTHVzXpcojnz0A/1iUVjdwsavDd


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ok18vO3V1rhlb4abKORQYLRhLgnBOcMrwB+kbHuJoo5pU5S/RZ69hqRf2LSc
6sHm5bIqXDuI2tZaApXdMnmTP7jnjkwUlpT9x90TAyvRkJePrXO3WO0ySMwV
tWGo+dPmFBClfMWFNOl6iuGFD9mP/YXD/6Nosjtl/WYvJy0dhi8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MQTi0rhRvnOGJxSkmcukQH2GlvvDoCeepPdZlMaZ7FV2fDTzmMgwWHtGda2e
WuhA6Ym+4t0w6B3/4L55juTCzBMCW6sNWlRw+4mY6CB9gu64ljOa4fs3MiLn
S0gwO6RQG2xd0pmjjw++B/mYBt4y8MyahofvuKAEJn3YG2jAluY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9008)
`pragma protect data_block
stQyke0w8V5Ppgbf97L1FiyXTpZrw1PQxv9g4EzIHnyfo6PVDvyC+/KbHN6d
2FyhgqUTjXt9D0Z1v9cKGnoCeLKnNq4fVSIz6fW36nuWHRBLWDb+3BaDgYVs
Y8xH4k26UEngSMMFOAM7US0pd0KzVcPzvtudxt9vnIpmooKGYOW9LRxUKqHt
A7aQqcS2zkXVgMcPJAdy5y4nY1SaM16JBaefalqp7gCLMpon/QkX+vnlU33r
xFdE0HWnt7cSLbWd19yzhPz7uVYYoYa14sDtDLR9TFTULEPaFZFmT+zcrvTk
hQynL0j3+Higj/paNL4nwUyxpEx7ubdmY2UE/3s0gLJo/Cs9IPDkCpl4k1vw
sza+Wffjh3iouZimHAJ1XuovVuYJUvxUArFOBofbuzCAw5VD1jdJYRprLNRZ
h9ta+SWNlq0+IVZjcuUfYP7ZeOeuF0SOeYC2R99xMeHl9jfSAU114OU/nA7x
OnWvCtltziT6pPSMIPm96u1D6j+CmptKSfI58nBXWRdtU/1Ks186G+Om4jL9
xtTKX2lv+8LdY+Roz2iDCR6PmXZ8sTe6l8ZESOHkBSojezethmQsY3VJc3bi
afm20JZWGIdx+EHui4C+iVh7EAiIZY0jIFcxicFXxnUFHXfJjIZhjUhjOJWt
Z7NVSV8ZmZScpi6v/0SXZ4I8RBqqXd+ONcXhgvJ7bYjuee/ugdKhY16pxz/I
h7ZVc0Kfcaox1o99TuGYp8sFYanxUiD5kIHe+IyzfxzLanrEse1cN9bGmKW9
YADycMPKHKAG8XJTJs893Q7VP9yhOPvmeb51/1B40ojvikHCAaYaMtoGjaUq
NvIV6a+EfNZvqed06aPV6ozl6WsZxtV/9Le2SLlWWVOS+i9fMHgqZgqYoicw
un7DNnfOjV49Hm5lOYgrD0LJzosABbpOONX5wubXMSKQF93IUjK2WxFeeqUr
c0Prp5QG1j3TqYKbpGyth96ITW7VnoEZmwHoycFq6cqPNZLPDgHzRAiMX4Ag
sMAid5qnsDkB5InZ+29EqQHLICxsc6PNgpXEt77h4p3OCpUCocTnbCTBHYe0
/cVMT4AQFSk1sTT0GwJxl+g7QDAZtqWlPfozYs8WFn741L2wTySfNe+aULan
XJ5Vvp1HG/LYYk19PHAykNyONVMBLcKsBBPEELuPTIuchsJeuTNM8LYSF7ux
4/83a0eN8WSLncDFMG8rZ+i4Xr5jlCXJ/ynE8kpXTeNURBj5PobYOKmcsumb
2Cxq2iesy1p9DbCuGytqMCHpYsicnMIn+/MTVd/MZglk4I3YhqOHfeEi5VKi
ZtT6GrwZ1Ol8FZqoF8L6U9dLkZ4kDqI8pNNHwz2Co4b6tWyGsx5S9ob5cXW2
4Qn2QUfysZi8GzA4TZzBHW6ZnM/X/tX+iGOIBPlzWw5lxPJ0ndrdFxcOlLIm
Ve3tMegSw82rr9Pgb0OksIu8zMUL6I5lJAFpbT5iTXIAJdqTUKbxKBRsf+BE
qoSz5CEj6uPe9YY3NI6p/ar7EEiWcAjtLEgwXAkDq9ASv2+EP9Ysl6yLd12i
I3lZSPfm7ZaJ4StivarieRfa5I6YvGvVQQ0ycxKLNrU5cCicXl7HZNY/01lz
EVZbaWUVInpdZmw5od+80IXN2A1mBiFLemzo3ZDgJk81lF6ckGp3elsGJHsF
Xzkqnun3pTP6eZYJ9sn7WKPGPG0Ha46eDlujdPIlwmyQq8WP/zKPpxi1amMM
7vvINSjspEQFFGRhYuvW+ez3lxzHMn4HJbi8idfW18Hdkar386lF1cTmR7sg
QlSXNKiEyFaGwRtdLDUb/kXz3hM1C4EO+IFhcRQZUVoIC/5VraT+xLJ9iZjG
yIsIDL4q2ErG7D3GRLp3B4rO0euf+ggCmpqbVWBSGop1UkRy75fVWSnayPlU
ii7aAlCSK1SFujp30EeuLA7SYjaWF0ihNjK3sgso5uTMPiZ5G1mwEEZRs+GY
0OHMEEsb77JRrWDB7Ljg8u0UOmW3JxRMvd5A/VM7Js6kIO1L0TtNtykUKi7l
1O4kWFhL3bmAAFRp64iHlj8cLGBlsDIW9HK0sj58dsnFNLtCDvMQaSdDiDDL
DiPhvWGya+AQ/ETHBx0SQFdXS9SKDSDtVlMLrH8qTJfKl68A7rGEnQ2LHRx8
868NvrCLf3lc322X6zMBFuawm8KZePvb3S0Q77zLTtU7cZ9lj4oG7PFx20KA
/+FstCHt3C24POS2Mnu+Kf9hN7MVr0oNX8CpOI9hXT5QoyjGYiGxl7uVGiu3
OY5PaxCRoc0jG3ZwCw+l0xli/SibqbiGKLboPDAm2TftYucdHd3mVf+OSdF6
B1TLL6xHSOqawIqrv32kuEstvwMdAqXncjmUVb/qxshtc+H066bwLlTSphdf
3XiNLWoZkoAuv/hduDaHp6bsl5f2dQhOeV7Zs+LXyIlDraP1XeQZcZEfS9GW
23FT1ui2YekW3wgKpBxTzjEp4Gcd+YPGHYyy2Qd0p+abX4zbUbz9zgucqsXp
/N9elZLQCy6CZ9GGFS/LjmCfayb8a8iu8GH+kPOmGFo0Vums8LsYi6tHsyIu
vjwtJj9JTQVCDJTFY05y2GsVxeny0eq3EyqFR136xSGVDKPhwuiRkMziNLcb
hjyJTVr5bCjbXPUrIX6R+gHXYJj28ZyMx2Z9aHLMGvMD+WJG/thrFTH70gl9
666jyTP2symOsPkvcqU9XwYdrhjYFB5iiKRHYd1lRafZvGpJMMtioJjNHmeM
6i6rfjkA6mA2aG2kaE8BsdYLzYcPy+hkdLuez9aelInFCOKO9zchnp/Ahope
Far9m6yR3rFkl3aPb3nh0QwGnVdfpm5Gz20p2qkb7loNKPaRxXOYxB0pqtJ8
I/GVe5A8rAjYcJvaUm+BKaRufWozMDNBawjSSWk/T8Sethb1VrsxCSyAXFSH
Wow9HdenU2jK5Naa0G+NOfUpNTFZmviQ4LMDZRV/3E/SISR+Oz/eanO7A2Yt
RhqFjwByB7tI+BwUnzq/bXO6YXDnWS7lUT95ooF3SLsEBI3WWQfOIUWJmE4t
tDoZaO8jX7+hQTzjJJ3FZY1VyKRSTuKqygGIEgOc01tRlQqHmlmq2y9+g3ej
l9/+B1qyrcA/bfy4X9iKbs971idzJeOIgAtcKLGvy5kxc0jgYfqNV4fvhRRd
weg/y0tagVl6JfM1xJG/1jh2AxWAc0Cv1AqeQAPVxhXMRAqEBp+O4aKRQugQ
Kd1cgvZ+SW2opfOJ0QGnBEVXaJfKAj4UcLvW374ONDbf9AOcXPFXW3Oc2Wqo
PctemHxzNHOibG3I74oo9V/PKsBzCFaiq/UZqMDkXDUtDGq3ttWO0UhP2xHA
v1V32WUbmmPCly2U70pcBM/z7tPtg/AHSElWnW5fnNZqxq+lggXifc24klvv
Q/c/Zc8WfriY9GPFdxjMsh01B6t11QnfE0X/EeAEbZY3JL1QzoGozdjB8GiN
cPQU1hvQywkrZ36cZw97iulKNTJzx+Q7iUi2+/Cc+k3Kv0Qz/xwKVmu+pXPv
P17sDWNcc2xIaMgA0flzA+xnhtuHixCS/shJH7dxjxUODaMhUXfq4VxUjVru
aiaZjaMbD4ifNu3NeuFjQs2cPTU8IE12Xtk7BSvzQQ4qvesg7gQ0NYq5SJNH
y4hOzHTj2sWx2tVnrxIUi2tA8qs8essxuj2aVXG0H9/o/Kfv8wVgevzgZWpW
gqh3WXFD6hK2hFDfJeqIilv7kIx3Ki3hZzvo1Vnwjz+GRPKDHoqyz3QcLfSR
Uj8pM5w8Vw/eWzz4p+Sdq6XGtaafud2ePMUI1qR0SynM9BokuqL/aI/wFg7+
i+p8QeH1mkDLZZCC8Xy7tA0mBE3usQGK/PUUuw0VsdlXqixqY0he29JPfjIG
9NC9IK3dV9ktZW+qtWgczKzbk7Br/EBJN7+wqf0M4WubBcr443WAnkvmMQI4
WxIIhbi3lzyf4xLboT6meercVxBH4BcJcTNGwhf7XknX7zVEktFuVvjmHDLT
rJJVFrouOh1Qm/yJHPYzHz8rwauYua0S0zyvXW/BhHvp7kp7sp4k3XVUU2d7
FODM3s7hs0Miu5qrKiqeNMbS7jcxnFLxyO8k3sFAmXaIWLvTQPEbrHfe8bPr
on0bgLeLm4MoqU61nKjUNkJfj3I7SYPcV9pkZktJUPIXWigqprRSaIbUWtpo
Du8kG9hQKL9AKavZMcRioCA/LliJPuYshm+sL2GK4VXo1bNqcUN7mYXUDeDs
oBxmaundXoq4ZCmJqxw9SkBA0EMBVnp2jPp9AmSev6RKOpX38WGFolQ5nceh
sVtpW+o8ohB7TNNdTbRJYLnXxukmmlm8/AnfcIUcKDIMcZLGDIlAPp7tAeJ+
ikhcjvATanagP10Dv46YyMOEB+DRFr/HxNrEA821ebUMQdHyDC+0QPHkcvn0
gAwsBfRuP/ay811mJUx0SmoKvE3fGawffAhsJKkZK/Y7kHSqmwG6j1vraZ5D
Hfm+Po3pBzWx+tWpiykHa8GkotmdB2UXdcmCdQ9dFl0l95BAetH596/lTK2M
nOFhZXPYf7CRfyl+KZZLVLgUUV/unMfOSYd0F2IGcjHrhQSRJTSq7mX2ge4B
5LDKavM/nP+zB9PvJV/JNwhBgrYDlwv2ATSTdi3s2VD9O26SK4yqmgM7PVwA
PYz345GyldVXWjSAvgFAygCyzl60awz8NJA4NRGkDehKjYavgD+4B8K6E9VS
qryBd5j4YPm/x4rYpPZ1mDymyShAd7E9PfCHExbzI/q7FKSLGXR+KkNmR4pA
od24GLlAqaSvqAdLCiprLnQzbrr7yi7Q+S6oXB+t5Yki9efI3NW9fST0W0q/
zoLqozgwAg8D/XL6pBB6fJLcv6q9KVBElYcLKeFMZccF2/HtBNRHl+FjmS5v
MkARaepc1lLQDKSbOhgPsxBHqocO2oWdnedHZSbr6Hht1xN/sA53nsWYU3YS
wO+DzqWbxG+oaPuJrOgvXVx2g8nVgsl6My89L9zMSONyH22JrYRodlYhAA+B
3NziF/xcTD9fmFk/aKZDObnsfDyoUaN5Hi5fKM0ccZa82kIL9VODXjGXnBQJ
RASkw3LeF5/5WIWmD0QmU0Ex2BgYt7YQ+y4eW4bku/BQBP1KW2HUL1q9dd9v
jcbGvVBzvZ9txHr2qXlUjEzEDMDxfdt83dpT+/906I/Pi3E639UzHQY5qgmF
3f1jrjn9AfpnAakrdbZdNg83JKnl4NYDFLiIRG2ikCiYbzM91IgAO9Ny9F2r
8jGHbID7UCqWOKrcmvZ1LxZTudTTbR8IBRlHjrTAdvD6W9J5b6gYOetR0da5
4zLN8gEkmbyffPu8CHALCsZ2pMyOElG7E+y9UcNqr94cLVzoPUY4I/0b6lpt
lKu6kXQZEI4kDhr2DT3tjcqbteENoWbegpQOfNI+qSAAeW0+sbVirE/tDrJe
8tDylhrVgBv/+3AID24ZRRX3AmpQoCpeEVZKuXCOuWlmjueqWbZsHm3ybSjr
vIa/w2mTcfWDHDlsSFHSxU0dg29L3rMZ9wpKbwSQB4i3Y44KRy5Oi1k7NMoV
NFTHIWapJAdIaPKYO/UXYU/JzJEIY6jyP5tk0VRBYADoKWAoe4XKVNfOO8u0
w2SPPbhQWpkV/9kLlSa4gkuZpDknGJLPLRQDpZ2I8q4HoEJeQQpX3iD8QijT
JDh4/23pDSsdRr/R8gZgC40YSMjQmItM65ktjHHf6yvlcXHSXql3jHuTrs4R
c/D/CxrebW/pu2AY4A/SkVOaMojXMUarmF0VWf0HR4c6MahHcrx4q30grFve
ilm5wEe4nrLZaZhQOpRqrxuwbMTBm9jWLaK/Yas6lRjgaLSHStoIakVlVujx
lSVDydjm5OGB+vCQj7AdSPEUA402R3Spg4doz/QgbM6pQe3gTItuwjThxDYh
VWlA1pXVVy/WMARjYpjD1URoC9GEJco2GmR9Pfnb7ZFTIqmz/CJGnbBp1a5A
0bZ+hmsVLkWw7qvXnzklVgOkgdyTycWWYfh5Sg289elYLS0zSVb0mQlDFfgu
nFo7+wX4ZUyUhA89/4r97Vu+tSQJx6PDKIUFx0mlGuDxNDwrpizlbVTL6Xtv
4Yhr5NWt6E9aI03frUfPq1soqbkWuthT+IROa9gBGbOXQcusGTzO0loGmdFf
xcAiNmUe/CJMNiDuem2/INsfy7Aqr9tu5jfNLAnGEAUTJ2OHex2Buo3CbKxh
USx78wwltFIxUk3qdjrcuxRoria/hOaVtIj3cHhYcHZkS/EayuZVrn2hmz2/
fsyRY9xFQlZNncEYTviQlKDstPI/ecfXtthaEdy7hjR/GEQ2xG4XnCJSVubn
Fd8TuPpBcjp3mZIcW6Yn4fxoKke16yvbvcZNiwE8CQwGNpY6G+Op7QQIRjR3
OVp1LgfPpKFuDjNnzH1nCFgd6P3FkfYfvnz9fAqYVuTwzhUKocOkxTMshPMV
O14ZlpZscYoh9hxaYaZ5cxhuWTamt37Vo8au6hEJ6ipp8abNu4+jRVEwNhNL
eLT/Z7Uq1o/X6sDccTCytVgUEr34Dx3K2prKKanmUdYXQ2diVUT8oEmYxfyv
K+TvvH3MZ/Lr/H9VbWfvDHjjfdbWiW4cB2FCQNJtzjwAlJoGjhFms0cKiC6K
6zNFIq/s+ztX5c2we9/bEKHVAoQ2CnIfUmR6ptJBxH1ihI5otuxBllr0mnZ3
vD0ADx3eXuPXOeIGBRlvbVdqP22J7A3GAEZy9C3vvoOc0O4VUSZoaSjcG+M7
icu3Q3Nqs41fdUEyGox96neXvV86fWb6+UHfbEFc2pwbbFZlqQGq7TfH+EEI
E/jSyuv5n0io2zLkFg43LV6k6p2+xcxIGqFF64zdKWp9jJB0aY9nBko3Gz4B
eFjpp26mYApPUBxTSh+1zLj1tqBebkqe25Y67HWxvtjwZxLpyhm7w8tOCrty
xk6cTZcvQvvMEWKAUh3BAmr+ekF/sWd1vcqijt3WDzRZErq1hTIN/kaG4y7z
nGGUo4iKDOMyE9YI3rfGEMed86K3NrqCAEt97KrFe/QS1m0+PtZ8iGPoHgfb
s5imrN12LFIAG6pbKDVRRQ0g/20eB/jcDmHSiw0S3UOdJ8mMuw9SMU4FVvco
XmuF0HReetgk+hNcEs3tXXSoKNhhhL4NgB4WUtTtnUEZFYtSZB02CEZ4E2CU
e+MJLnuEqhRnYmYhx4uNMKf/hiFh44H1VAYV8AsN4K/Ni9UEfu36WCskdO+l
0FXZcmbF3GTjewUGXIxOxns7fdrS6V82Kn/pWmD5dnc4QHyhYLwCEDT//DId
d4/w49sbykRU/feW9INKhq80i+YGe/wiRbqHaC3tWXtDzlPww2f5etx40lM9
ROTaOuTyzFLI/bfd42by3TOXuUwu18joQH9CNgI6tSJtRx7eZXVyUcQR/Ug7
k5YyLT3buEAMHc1Th23Ib1AkuIu9Ri8uhgYZ7ntsG5sjS/vlJMHHCAyWHZZX
weHmEaO23AFx/+L0TaLmR91OmVb2W8vnZrrKQmZ2tjJi1tpmGomkwMlk1Zsq
1ApgHYHl8uvZuX1VozpyKQ5DaxVvxFb5mPdl7sAECkJlXs9u1E3e8HSxKI0r
bZ0O3CACLSSrlWHFJyUTeu/o/RgC+UAEW82mXE3aRHRZIrCJj4DGEBK/L5L/
XJ6iYrtukEEwedi2lsRoKdF8dDhUatwiMIA1+ddKdCXLaZl54TfoMzWgEhQW
dlMjhyIE30I+TFse86HHlRM7FNmIyG7zqT7hpDZRLhtYa5Pw1KhdNgXw/Jhy
S4Al3ANwdqQ+UG5p/LEKhYHkRmWCGPbh+qrSR62YWf8A6LZGmwvsi26kBKWs
nwRJ8L8RkIwwXdZiBGzkUzM9+wOQtS+k1FoIhpkrAgO47Niwkdr6tA1R8xLR
hSKwVxUJ37Mz4V0acwg229uWnUWo0+zTA9iL1bu1SO1ghcTwpJIwlXDtSJVA
pQLU2mKVwntLMy60YOQOUCwuVAq3hn5gI76OGsMwowUjrTeQTNycil9lSUZ+
onwxabNd/jTQUaXxflmQAggq4sBAQnnviHr6tJ3EPCZBa+lqvMUZgK6oxMid
01E6x0/evrpfx73qEUp1c0LLt0GPS/wJ0WwNfpnLLwf9tvcl0zZOd/uoeMhm
hd5MR7YQUpCP1QV48PdsNOU7F83Fr+hnw4LLslKT4npxzCBsu4YUkWQ/Te5k
1w5bx8th8Oow83BTbvXhJKUK8tly3yqHfPs0MiU+nJoFl8yP9CvaQbbfEElC
ZMdm4cqhXfLLc5xb13vNc3M9SMTeWl9PHRtKwdGQ7iIhvEXoBPvF/nszXRD5
RLVtTziO/dqi9OqTP5eqGdeWI2DatS8/9X7k4wOJAZ5yzkCV4rSUebDi7MUT
rHu+MS9S7I/boNyzf0wGRMzU3wcs5HeKWYZvZjR2qmjyBPrRy7CTcMBWCBuD
963Sw9qkS7dBZ9dbNPPZJbNMsmxZ6cb+8rGL4UspjGtVY8UXPriFVBgPbpIf
NTt19YrYEYGkGd3tiYEL35OhdELsGWJ4Lu0pNB0WB84W0i18Kw8+eh67oKIF
6dkqGHP35xQ9WVpZue+XiOS7nFEFAWQ/Mk04/RRHEM6eeQP483d17ycsfCC2
6kgPOkCJDX4q337JAlKGP3ikQHFzPrKfjkeet2VMamofKCIQq8NZwwlhqowF
TIvJfdp7RBdWi4VGeSLPJx2YW1ghtFQVufSEE4V9+00ZBGHOJypBRojJeRYp
54AoTRHHHMsp1DqwJ66IcTd/duywztdAP2xLVVst9N92M/8IeisM4CvTMtzW
DoSjwBHNZ5behcCZ9O6yTi22iXJKtwOi7FTx/uEBzfR+xm5y+GGzMdMf+vvp
nbJB4vU/YseyEph+YwCBgQEJgMaKgfb67ZCkER/dckp/tXdLVJ110WPAzpSf
2gk/guOXWEimLZUhtJNibbStZtczv2OGWHoejgIwxExG7WGVf8VeGVZ8xL0I
b5Vnn+rclNHJWIUXVfsd3qZ1z0OUddTG8mz0zFnfPt1vb+SMqvy7D7KVzIzm
787elVxwFYR+TjOZ0LJuHFIH1quWbh2mdGDpTUPaacH3q7fMZW5ZXninx/0K
S2B7a3flKYUVKon5CvWqNzd9wEeDakFqCLA2medHLm3ft/KnGH8OXAsHfVAK
1G6Rgh35IowMJpqZjW9eTql578EubXW1pPfTPwsaS2MpgmP1afe6dBjElRjH
VLNYOMygyAc7w4/7EoCVeEGcyLv0DAkCYDwFEMWaUMBe9pKAze8xMGWPhul3
ORJDs5yE9XG940kDnmVM8/ksdKFfeGink5XqnvK+i7H6ZsR7CJ2raoNUv3RW
IcK1Dxm0LbhpdU1Pnw7zgae/r0FjrSWg3g1eF2+67tuaDEXbATPy4U4kEBOM
IrXZynqwYG9j7wEQjpS5xgQuuOzQVpTibu7+RKexKxf1Ar+pTP9d+eAIOn59
t0PDK9IkkuNfRrU1TrM/aRjPcqX/+L05dV6ENFAbDDil5Mc/0R8ogqVaF1FW
blQ1gox4Y/37X1qt0T89LLCBIdL88YjHX31JGMfrE1oG8Ba5s/zWxD0t6a9U
iXmAVUq1ATykarvf1GD15RSuwFklwLgNxEYysN7FhLeM3Xn+DAeBSjhMguZd
zmZk774XLrfABkJHQczXGzgw+tDFv2QyRZtaNRYn/QYjHaqvirhHnnl/gk4u
f1ht8grpC+/EtaS+LN5XleoIt63rMP5B6QRH8Iar99yKl6EvHJ5GWcPUPJAl
XxHLIigMa8d3MQOxNX2RxCRFiHt6LlfgJenhfd/2EPL/OJKDr8BI7Mh8WoCU
MowhlHAub6NUCqlnywzWCORIXWyWoZZtJKQ2hG7gm6V7QjGtZoUszkAVrUkd
mpcsS2ABjAWpgTlpaIWsb+odGuY7FnXXCqluaQfLyGIwGnCR2GKJgHxpZ9HA
Hr/dd7vcF4gfe1dlVSiTKUuWeOGBYmV5edhvAfWdIbMRtjDaMJd1ZTeXMIIe
Q8pKqoq4kxu+YL+BXpJ3B921VUHMgB9RXp1kcX2FeQWB01crf44UjqK/chXr
lm0JepFLS7xzxKYF1fGayNOTe7ANDucAWyHhD8OEmX92aAdkUR+G8Oo/VmfJ
QJIgW3Gu+8l7vbD1xdcrnEhy6TMisETDVHsH4DqOldtbXuW8UvKgUERoHJNL
n4Rei4RpMSIYn29T+p4at7zJ89fGF7tfJo+RpkOIZ9Sbv9BRQvb6L98dC2aE
h+57Z8+EZ7EmCEECP66Ug8EoWMqQNQ7r3Bd6Pql3B+WXaozRCEh+GnosArYs
l4JGONWLk2PxtYYhvBjzFwyFy8R4hgv8f9GO/6y+zLwO6ACwbCVbMUNgg4g9
0nHQB0itNFqZA5kS79dFICgW5WVY5G9fyDLpLEmMYiJjo9jyzrohMlB0CZGy
DgKsJ1Vl81K+f6XZv/6KdErruvzLg7kFhcWKaSYQ5mWIpzc2kmQtt6QwsAvE
YBn5Bwy+yuY03yg1OnWevsm9G93W5zSGnyQ9KMvvI/5CMqHtjpvY6hYatY7c
X/oGSe34edCZfhPNUWV7jdFAIyhGSV9oyDUlCdTp2fvOtu2jMs0cVadwAe2j
Ve+A1+cGe7ZnhKizqHSQpwvm2zND7/MoeX2aFG5KapxvCErlGd4FldLljOOH
hmXy08icdqvIsSTt00yNeXMhOerU8UIm09CarHqLCF+YiAZjJB0MogEEvN2v
wXnkkA+YVywE1ipz2PXdNyLaUwDeM2K2fOv1o46puGmN3GnacAekwgDti6oL
4lRSjZa5xUDocHhVETCx/xD9hBl1G5P8Eizgfd5to0pit828Ag9kI9B7mAaV
3Ya4UAmlOzFBT0G2J8Nd8bfNoxQoAC+cEv3Ql5gl39fD9YMyByHCLfbJKl2j
jb/2UXFkPSKOE0SZ2u6G7zRbZwTmKOlRNLnqqNV7maRH+DKPcSQnF094gtZ8
F4ApKdspyAnqPeDuWeDDbT0JHA6d7pP1G5DQ6wqI0ubdPzPUtpxsmr6EPNOV
Y4g1bmOFrZKs47T47HyIpvXdl8D+OyZ5IQvJzNpj6ilZUCDnwmeB7M32K38E
jsXF/jtTd8MW0kge3JsCOcFhb1NsffUKheTaPThRO0xrZhGouL3ELjCwUjXL
kLJ+Z5Hsi4gwsBPNOB/f9pfw3uwQmzSKWrVte1m6P1QEI1d7zVk2pgB4mN72
x90QgI58HWwyNwVBp8F9PW9vsL6fkNmpnrNi/HN99wxE/3+zz+u6ky6VCRnm
Ghl9q/rlz+N4h7+qBpVXFTXnDcFMf/f1SGdQJy6v4hV1C9J9Q9JVJCoW1U5Y
+j+un5xetQL07BON2Hv9qo0vaJLHIN1vcqSeDGh3HUoUGQ90yx4eNggUVgIL
dG4TGC1nMjZeLxxEX4xrWysw51SjR8WC26+34uDUnGdBM6jNorILq6jiOJ21
xwWaDeLcvW6i4ak0Ct9Nv0FuFLximh80Wlc5c/XVZ2Jcw+NN+fDJMX79W5q6
5BqlEMqOJ1fW2pf7Zqe2FIvONBYCD+uPmIsYJqXm+sJmNmmFoj0TDgjyrIMD
ubRg+XorV/vovnmBuIW1y3Y+L3CKjj9Vd01uk3QsPG/3p9pgZ59OKCiZedP/
s02cs93hVKjbBV2lZvAFWgC+K2sCQTyqtbRO4awo4LVblLtV2nLMpL6BLJq0
9uiilDnCtaRVaXboIYQDSL+ZdLrMLXlzEJBNgy+1vLQ2rV0wA0mrlTIe78BS
g+L0BG1nihJAFKHfi5QnP7e8q97QEPCDvghaq0bxKuS0U2OYYwz7eZ+egC3X
mY+72o0td3eLdK/PYOjNQC80vbLzntME21SN9+pGZ13xTTT/YDobe6OYR2tn
jzkgSBYcfwLzn2/PU5PfI0cRvVePHOOifxKzFc1m1jUf3eica1nQyq+BDuOT
FYQG/e2Q8XNLmbgKUvNLpDlfgnvGZXk5XICaehuL2tPT75LfIglJ9XU8be9d
xSMuRfgqHB8=

`pragma protect end_protected
