// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ShDs0n/14TG1XfHXppNUPS/sAYDrIjYf8tCYTUFNjl4q4xD838Dh/PZFA00pVJC+
21Z0G7OB9BZoHrPvi2D8q8LWrvEioWV+axC0ZsvQUgq1tHIdi6vvRf856ZxxpQ29
LuwMWHRLPXQiomxrS/j64frHz+zHre88ZQEWe3f0QgpZcq7Z5Mj5lw==
//pragma protect end_key_block
//pragma protect digest_block
2iWiU1kyW6od6LWQSAFwJJs5/g4=
//pragma protect end_digest_block
//pragma protect data_block
tlI64g5/4EpV0R0nvKWfRtIeTkLong1V8BoVPFE8AyuegPausMf+txz7/RujiX3i
zc9s2Fx8ljg2W36yoCZrpnap1MgEkkuojMxxqjwHJgw7ibr23bban6k8V9m6yZis
rjNoeHJLTCLZDHCOo6ya/Fk+adjpVc5RO3LzYMkBm+Y24PGIqwbgItCezxBZWsOv
7+yx6oE1vF42PfLDxvwE51Q2fn9vxAbFWgN4y77h15A1kMNPwzK4gjga41nGAhX9
uyOeuqRzLvez7LTe0YDFZxzZ8u9pCqofYlRnahiCFaBi1oMl96j2PVS+ZQ8be9/0
JDGztF/EIBvcU2bdM3JtXLapXfnwl9shk/vrFswPKU35FJi42o1PBTbYsi+rdLGT
9PUGoUXk2zfJPRek3ThzCOWZZRsMxaOc6Hg6ApbBX9Tgi7LooUb/vPgW45crHDYW
+2HSjQJ5sMlCpUlvDrapJyosStHyuIF2zuFdK0XJq5BZ/wqoSTFYrH2yPvAXlL6t
yiXcGbGJw2d8cICYKijE8CnEkGbA+jcUh9BREeY3uhFOHyiDkGZD2ZcALO86Dwz+
VmQSEDqWJDMIvfokjriJR7rZbPlVHz2mEaXoi0BapqIkWRdTz5RCuXQJl2NzDPef
4PmM1IalD2gg6Y71mQCsng2OC6Mxu5WCcf83rqlh/4RIouMi0rvrUwSNINZi9O6n
GQbqIcvtiU6VOQd5rHtw5qk5q0rHdVFJyZBNVVVo1orhJpOkghW9sgbMq6oODX02
IcIYtpLs5du+bODLsoDzccTWXFb0+MZRTbqrupzQV9hY8ktO2hKz7/iN1ywfObuF
48QSPy5yWpsFZUjet2871YgN9nGo43KOJMACvKxiwH7/BbXG42h0jDiAxFKAC9HS
h1mfzB8dkuR9fy9d+ARy9j2caSxiGaUqr2COUHJ1/sUYJbnCiiN2IpyyWDgVNMza
fNFG5Mt7x8blJXhnKSleu6KKYOvyxjtAXAQqamFeWR/b77yy5Ejy/hjJBm1rgVxI
0xTCT5jR6uVnERESgqpv262oAEj+a+RC+6jSL868YdsRcNlRS0CwtNux18MkzOkA
gT6grZ6DHYLAm0MX2MW56x57ZyjiUxKWorV/muHoHMbaBo7uVBqU3yftQ2b0nD9j
O+B3cgWaZMkoXnglSdvdpDr9MUqVRCVnv85MJ4gtDGBfBR9Zfo3FtVmAcp+NPnnW
tsNI3WuVWzUgZ/r9+Job2nT59sR6f3EzMAveKxJ2Yzt3WeWGySKzdsbS3qbZkzq/
xo4JNBVEKx3bV5dZ3XkwnAWA4+HMTnQ13Sbk3t1txKrb6FwOfV/S1rSe6lMhajQo
ubj1eroqgEkPebi0orZgzUfe2AAqSmKFhlZeAsxJkldkvSP5dK+owTYbveDPq9yy
uT230Z0GCH5QbtDXz26Gx6XIirAqPwL5uXakHQt8Fgp2fJXsu4lJbUCNJnOhJSzJ
4Q+We1RrVa3USExjZPBpSx2LXQXvXnMnPK+6y1XkzGPZUFqzh+K5v+fmCSHGOKBO
golhm3DVklIso5dNkJU1YgbTRv/jxGFEkRgPeMOHwbux1umHk+sZfER2KdnALHkE
lr9H112nn1+cTrjhzrXmNLhH74SBZH7oGqJjOqLx+aanxrpL5sXY1xKE1+QwUB+U
RO4R7GGfQyyb5iyznMFvvwo3kNLOxKmQDEWXKY4mrGyPAB2NPoKlr2AOTfsp+NUm
75XAUNiyEP13mylklirFCAXKBx2gKMn5Vtgm3kJbah8McRQ7IvsJMnVz6CCpgwC7
7CMzHuUx4EhdkSYwvJjwiHgFVpIKPBWtiOUy1gOMxfhDf8XvUj257PvI1wAyWDp2
MepgToqjF6o5N2RN854dlgSdl2SFLZUCg1tzyXq/FHtVNKm4H6gWLmzimn63fCQe
sca4vFJrQD1qbW/adIDiZ/d8JMHzDM7zrhq/7sdaku7LZQqt9+ng+nwoNaKDcea3
RZAcHcA30E7QrqRSonu2GdjLxYwe+1cMwhzytqOhGaSimrb/glc30k575cme1HTF
qWuVqkA6AVipmVOWC0MwsaaV+2DeyNRrkwyOf941uMXCL+nTnXkYhzWzouln5hwG
3Dr9MlLntv+lJHOq08qcpqQAQp8jlc6F89MpYF89IcH+xIdmxosw5DTJcEn+KSCZ
Plj9qU3gfE6haGoLX2YG7kGuGAXadrI/02/xxZcMRMp9EAiOmoiV8vQPludeFvSM
nP4spaxIPI4V9u5sn060YI72VqVTynjOaP7Jm7QYxl6dilwaqqX2WZMdXLB5aucq
bUZyXSQ7I90vT9JvMbMXTWmHLqETXRTO8i0fY+UzVLHDpMzuR3G8MuhmVKtjoaml
Wjq341jmHXns2Tw1YxGrIIx/T/VeTNSDlOr57QxUbfIyqoYcnMSNYawT+jRAT+0e
Kc0kIolc8G0UiPEv9GZGPZfp8j61ttRlKumbOXEAQZYDOylFLhOLNYrAaaOLzBeb
jMUWUqR9O2xFxY9LEHhjTEnQsVpdO7CeoXNqkLfEoGCuiZyWKItHOKPm3xGABM7v
ypL2cZps6rd+LDdknWR34slDJCJiT8RXb4hfvK4L/JR/zmxJ9HuWkcriuDqh7mN0
BcgsGAJOo1aIVFChPt8SkVAITF6+HB+vFYVvwVUANvpHYr9B9joeMbp84K6YuDNO
U5gdSrRui1NgYbINT0naspmg2A35sH8EgAxKQmdREjigL4AV6MTQlz7v/aUGg546
AVtCBBokJe/mMFNFN09amTAUjqD04p5j/brUvkbPejnqY+/GBhL/8qOZ/CD9buKH
dCT6miN8ltIGgaBJPfPn/ygoSolgg83AFWZltoT0+mAnZVDl3k8X9QGxA+oY4LTw
SPTvbeYqfRfLqggDlJONJYMqrBiPVemJ2CMaCNXfXe6mH2avEcu/HwyVwFslRT19
MR+d3216jaE5ZHbcKhfGyIm2Zf9QgN7WUbwrw4E2T+rqQxbozTgmoH3Ydl0TaE33
gdQGHzd1ywabErgkRzOuk2XzpuaMMM6kseAmEZCYBEmTQnT6R3GmItqvRXyJiKYa
7qYzpvWvZhQEuUgHGGfKXnxxCL+2mPhWO+FwcdbT0rsNPCo0FxmzIi6HrkV7a1c0
uQnO29LPaVjSVaUsL5PNH8JfE2FoR/9YUzc1azye4VdzU/F3t+FNitDRSv4LcfL+
vs/XP7dRNrD1mbnj7OEHLUN2CGh8q0ryVy7Ep8FwQwgPKEJxg2sqiVYRnnH0KTxy
tZp+0gFNu7vcBBqG9F/4GSSZRartHbbFiIk3hWYRKFY9f56oLaigt5kge5xlb0iH
Ip+vr+DmdYHM35PQ2wxgLgu191/Bb2inHy8FoSHUtDV6mZrKgvVec7pdljF5yuVB
FtDQC46kLLM0q3Nr5/UBcm6t4Nilt57IDdyCXlYEn/uyuVCcNtTzffdBV0UZHJ7b
acWDsXZ/0tMVSurRQoDht4YUK3W6HkchQrTWEyBmKMTRhXxvNWSrTqSqEdHtGTZw
JeJwxuIAVduswjORT/DrJqYHfJhhytRmkxe/q/0w/Ab+3mVZfGvQTU2FmCGreQVR
GQdUVLKhCTFYPK/NXGNWhcJ3Xs1Nc3KwYv73hAmcBtDiqFAEf2Ean1oZaNnvKA73
F3A5Ys/JiEqkFei2/yTKQ+qrNJMj/WZDMMxgtPfK1qtutGgnNw8XLJvCjLuSUlwb
10pIDu8R+6hOHwYVIBokxNwJhP4z/355gImdo+ODkbzPliL4olqRyHGfMMJCQkwX
kpE4be4A3R61q/bu71txsmZ/2iRAIN/5e4xeaLg6nXzy55nEnFT7E8JzRH8GMxkT
VP4euxH0jPhqwP48PbFohug8ts8uwn2JBDuWFQ4exl6R+eXnVDJxVwF6f3f5nCrN
HIAroc+hXNIaIpS6hGgj3oxJyYB1Ht+CejkTnBQU4HhnlixoIpTH6noJ73hL/dIW
tBzcak8A7xUNCeP4f6tMp4sT3Ue7Dl2LDSNXgCISAkJuuzJZtJkvplSFzyDsoUi3
e0U6BIvTl56GOMHEMwlZyDH5AI03UYlTka4T+Ei/FL91o1xkddUYhEQLl4dem9hC
KwdzPLC0+393xUApnqGvMtT4jejIYXstmaLWY3fhZpC6VijfA5XmIaNMyjcglWvU
NlO3iSw/nIPpkvFVsqBwl/smCu+Wu9hrTjfWQ2KchEhyIQGJLhyJPa9v+VQyqXCK
0uFh6OSXkw1+L9E3WhWsO1Nn4KSIq6i9dwTvWK9IRoDyx+rBO4SONQcdgFHUBcYn
FCfciXKcHZGwUyObn5MvwJOtFcu0vnbD1tGiEcU33lLL8uj3FF06eR+Rwgpg3qhi
DLiM/sZegIB34bOINcOUX68vRCJckVJ5e/a/4Tm/4mVC2vRqD72v0vGcQMRYraRL
nf8HmzaFqrdj0j6ntksIWi35Hzl0ZIxJKnVC3zBH22QW2Vpo3Sn87YWstNsvSPXC
71CzxERNm+QT8kB9pw6ByvSpotzAuwMzacBoowx0rbroqgABAjiYHD4YPHLnrdyp
J/3/8jiS/+celHib0oLd5NZjg5XLweUG+Q3ZksFjI2SDjAfZr6YLBsdGl+aCpbTK
B3xTOQy2FDstx/eJb8VLCqDIC0ByN4uAb040RbV1+X6kMbMwIcdcqq9eixnQlzOc
mc58Wpn7c+rfnkJhBfJLZ8ZzMY4vWcF96mexpW8EpDlszkf1xzhSgnGwp7jb8NxQ
NXpPud1Y/a0Z9QIqt3NMSH/NeL5/nWDQ4q6tgGQWye9r3yFkRFzIwEyo17QkEj5H
Pzzm3OAcNZ96cgplngjx0I2gbiCXzb3JH3Y2J4PuPR30Z4NzJVLOWSwDdwjkKg90
ku6vlsnIpr5XemXRWuzJZmAsBxlABAGKfCoj/+RWJspy5YaUMG2Wfq7kiyfmydnj
MqRaLabjHaLRq+YY5PYoo64L5FmN92Feec1GHCZbQVUGEqC9xBl/1/NmxVHuXj1a
TKXB5N3BtX+KjNcX7687W8ptCbjDbm6Yi0MEBc1XhtreF63qv9ME2d4O4Gf3IS5u
Q56ieAbH81gZ3tla+rw0J00w1wMshWs0NlRV0RpUq8e5cYy9R4/DRzcznCmHU5cY
W2atICEopPuHEEZM3dJ9wVaeRlLi1Bq1a6SuS2P+Mvp7r90dCSK5/ZqEKUjoGkZZ
KwNwarxXWSOAF5F1CV7MyfH1PtjywrxQoVSY93vJpbcEX2DXuNjwK9rCzc6M9cIA
Z9HLpjdxoKjmY6Ep/zAbTXP+wnUmiurqkGakMl048ohj/5LrDSwcOdn9sNEXes2D
g/VNMjKZgvdQZ2WlmBHw09pVQZqIyv3uzGbp06LFDgQ9XB434DGfUJduakdPOXuD
TFQaWCoLAe21aNk5+/NYpJRCYXp7EqWcRjNLXv/C676PtJezaI4+hRfPA3OkyC2t
+cvJ9VBN1nbRWBE/6GWo1L21nNWM2eHth5+Qdkq5nzhSLI32SkfuFRRLm1HLA3Ly
u1/Ko4lzEuROrkAt6iAZTr4NccybVDXTuMSSSWXAUg9kNZBjz2jpGi90uq3AVcMd
UVQT7eV/o4QlIJFQ62iX3x4jfA0qi6F6DTJb9dtO8FGsHQBL+zZ9VZHSdU/RRFD6
Dp/ciG0N1oFxF0S5IVHdBMM0mdAFcuFFWbVYs2Lo12sX8f0QYq6zopXP3+Ew9y2A
LRk0HvwBY3XimPzJhJEsrxIGsZ0TDrF6dqr2bS9i5y9ZZqNm15WVjigX2NroyPym
koZGPpuc76xyH8jjWb3DPcMM/twrYqZX9QgoODdEoq3xbivNHUj8Mh995qph3dX9
BNgZ2gVk+WQYX83XFMG8e66Umt83TbrFZV0z2ZhjaDMMZHcEx2en9Igy4i0jXrVB
aga3JTv7WzN0pTrbop97rlv1tC+btQyPFpok+L2NtWsKm1nR45NgO02EEVNfpp1A
eKkJRRtG124yKu+r9+Bz+Ok1CZwQK2K9k4spKVrG4+GRMKaSMcidXTEKmUhPUBsy
XF7gSpWA7631gZXhcswgvNGzPzJb+w630JRJ11P7w1K/9J8v+0ozRu2nsHOIe1Xi
9iHVYDYUWlUyWh0Teuac9x9A385OyCKuyCwd9TMS9b8JDCm6hkP522ItpMnPZ3aS
LqIB9lt48gltcCY2EX+VtqeNG3jXRqm3Ht2oUhBjxbYF+Rh2DBDFgo+yQ3rdbHA0
/LNiH6DLtzT+EEP7mpNdo2gONi9Q6uZbttpx0j0vFXwd1tWPfOxDNyaLhLKowosF
xqsPhQO4R1c0qYsJKx2X0ZjZjRB2e4B3L2dasUiqwGiQYLx5o3HEuhZnggPm+Zkn
CoZZ2iUF+l/TuzZGN9cRtfa06+u8UZ69TPEdxmKkPHkwLo1H6FL96kb4x1OF7oiL
SHESjQiIQui+bn+L/TVKMgZkcMNQwRmxxMSbSmAYYhDWW9FyP3ggSaZ5Gyl4N4E8
WvOKDNfy0g8j2v8rwi65q/kD1qvdigdzyq1CqLlRw/HIKbUKnf7xhqDk+pXwgQ4k
rdkRiLim8yvlKr0lhORndsoY/okqfBGts/l+hPiaScXCehJP6qOpMGeudToT4OAN
qTKbg6jvdwwuGqWapa8m1YwiiL71TLFYjhf9rl564i+Jg2x/7VmXoJYRAHw6BjgR
Bkr1rT4nJeWQ1xA68phPvSod0dpK/wG8Jf880dYxkvCx9Pk+iKwXVgpI1FoW6HzO
KRyMpZW5KytbAl5BqxMGQfvisiNVnvWckLCHBuiMqAyOJ/uu/cS5uRMTbrc3eEt3
Z2LT9OwJcEu1efc1mJMIgtwUMhsP/Rdd9hS49KULJ4GxaqTEuY0jy5MXMq5LbCz6
6r/fNZBlhJktBhSmoU88+AL7SlLaMKC80Mi1jIOySY2EDKBQNnMDl95cFxI8GhWn
UCVTSxkNYllFrCvpbqJLJpqF5C6Zvhed/1CArQs38hp+uD1dHNtNASuupTkG3T3d
QgzpJUgO0B9ieK/g5TMdfqaYppdyb/ZlvID8RE4niM4pRY2mlZItYy0YZ1DTsB12
55rGaqfxC3v7khowSA0STGAcBBMRDCpoaQSywZbjizlquYbQDv2YkmDhhJou75GH
xjz7Hb1GQzseC8SyTUeT0C8Ku3GBUvTC8ZQ3ESXTAp0FyQ2yaSchUDzsizQT/cXT
XGUmBc71FsOkwtrO2+2c19iQIuwuYhXZP2uw62xsWVUzzQfR6uXiJF9rDMDoSrWY
8qaTfu3Xtg8Nb9NABbsvDm/zsFFnk49WGVEAtBIHzYixAnrNmu2tclUrJPMJTjas
gt7UshklmHIjAILRo+0l3hIImtSwGRjQejBDI6cXdRI417/+xfhNTwSQte16rVYI
1y8xavU+a41vN/Dc+89g7dsCJ+S6e8Ch5fO/cXb1wBZDnZWIx/aYV+YmcTmmDpfu
EjzdhfPlejbULldhe6fFKYuvHIaSKeFxT9mw3fQXzIyL0lGIO+9TI3fKgU/Guf4x
HbyrV1NXBvGidQB0nEDpNDhKC5R8TYKLtaUTtAFC4GlOXU7JGDORJ+6F0QZzt8LS
0cTyRaRiSs84zzzmVIsZZIYxbfdj6fH7aSrZmAVrUvOIDeWry7QCX5sY7rW3mjIQ
+EvfT98KaRawpV32/NH/3AGlyj6fNTtyyUIxOVKLoFPPDccfHFg78UmZf6BHxuHJ
SZ2pcdrcdRsdxQLJrvcee0afbVo+kuvI2XdafQLRyYnToIENrpI0TmOGEELJNgrb
rINpBNLfKr73zOLTTlLezrWtUEnedcKUrf2iWcc0anImOOcnFhgwc9Ktw18QdZrE
IVL7O/hnMkR5FTSCrS/cmRo/8FgSxNlleN3bdkU0/yrTND6O9ocF4sT0m/Ab/QxN
cj6yd6255lN7rt3fYm1ErfTctIfMjadqm1EFlm1qNGK99qB+Y3hyc0MLDsoHrOGB
xYuLu66rA5fncDZ9NZqQSuApLuWHAY9a2NMVQRVYUc9ppHiYImjmLKEo7OhT0FvL
+o4enZ6MV237c199yqZJN3Pbm4sUsCtpxYmg4XSj6YZiP3de34djRinZO+Ak6rNY
DoK1SZPgnraSDnDtJrJyzunW3h/EykQMLPxwGK0VtchfBh0fgPKvkETbHsRNZB3J
I/yXJtlwCyfj7OwIv6KsIWduZwbNcJWWKUvDk4qugk78LTQcoqTy3pGST24Ta8oj
maheVr5CXix4iPSgtNH90iDvnmO44KU5wYUDXjLMjw8xyUY7QNxlXsO9llkSu/Ne
EFkrMeoElKO/donKBwvySKKJ5HsfU6qXPZr0ZeHhptntYUKiDHyYsB2392ahaLZk
CKlHTfl2e0Q3knlcQDhrCHtVE+Vipl2A5tM/y7tP4kSwHuAT5qPjGDm9wLKLGfK7
WJUXEnaakt1NOjrdyGYMreuhL6lmsrk+FcCIfGGDwMpyf/13SAEHCulfpe+FCUiG
6TTYiZpA/T0zw9NtMsr5csDdTcmdehkGToKys7yDR5VCo5kwkwsGskaA4+zWvK+E
dIsAKeQo3LcXDHR6bvoHG0y9sDR1USZSeJNsWDiL8CVQBGtFrohwfGIcUecdE345
qodJan/OnRpHp28zzVyZSUTyuCzLGg2QnCrVq0RNYcBDjnHOEbCkhBI1yn6keTli
jvOWXUROV3TcDLl/NUqNQemfMlZx6an9kE/6IlpWklgQDHRfzyfMLo2SbAz1FftT
JHWjM5XWVeLJi/Au5IYYbOGHJrLJgNcDEn3RZ9bgqJmIqDeO/WW8PUT1CYRUI1Ve
kXrI/Xc5jmWZxnqQvirokfr3r6DJ9KlNKwggvG5uiTQCkpB0zyJad1mpktMDkSuW
enhg4mocfui7wP0GtDoizrhE0g1yTq9UJ3nzp+/v66+++C6yZbmAn249bQsaKHlW
TAnhBjmjPRijhkDb9XlYrnpifhjpTTpt5+FocgIZXL3DFG6yIYUKwcgoEmXMU88e
X63ardWhF6OSmbw8HOwrv2k4P2tNxzoep8Ir1VF1Wx56SVU2o5MRKWJrnVqRrpoI
Vx2s/dsrxZUxua0s0LmYEtbr5Z991zjLZUFkxrxW8+ER1uJHg6rB2yqDk9OnrFSM
dEhoFHq8pvFZVQNLbFZXETq230Wan7KJCjui1Ut5r3LDTawGQrY1L+L5/xl5O2g1
Gsb0HYpB/6EuPZbNMukgAy05KJFie0Lzzq0hGLX3sycTltOkaK0/cZYF4C/rkHUs
5FtRYwpFEhppjKJ9hYv7F91aI4wLDRUFrTmB2tdsLL9NxKbMBtjfWdiIfLfTAQg2
OHH21HTo+i8eCkfV0Kldbsjl5/dxjI87yI1Nk5WupUhZnE9K4Gunferh64O2BKhY
Rc29c9n+vF0g9Ayg+VM96MW3V1Tj6ET0nmArBrw5tuGuX7uM4qNyOpib4UJlgRMm
LVda3oxQkZwvrVZXOm5AlgOXMNbCPsdUvZMsmeMaIINx2czg/FrSoJzm73C93Oi6
/uXJaSqTuSGjejWOlHpjpHCpNowhZUYUja/E4tEV5HIG3rZvvyzmw/ulKSpAfluG
wzNaI7VQenQBbQDpz95z4F0fizr2KMD36HnCI1sfxYSbxyaO2hDLt+P2NPEtF1a8
1RfyyLMKdXom6iaeH8RzHOZptijYIR0wmdUO3M7ID5mAYHnTNwR3fOX3LllRJhgV
9FmXD7hTCL99YOLlJ8gXwRI+MTPqjZT43/dYx3RUrgzjhVNeG9jXPyoV1I3UWTkK
bQd3flG8WZxspaxBHqjo5oqBh3zSIR3QDruUPFWplgemqYAW1Vvi+zqrEsrDSAaz
TJpRusCLoreCUHActFTNdEj03mqC+rKyyTuY4tYPSTViOf3Y2o+W9nmJrT61H9pr
QftTd2Q/qoibjY0qpID0tLo6I94TKUzJLLe+/M37KWjo2l16tUyCpVQhY+iGf8Aj
3/mLVZfQfb7cpzkp+37T97vO+/Qz8oQ5bETG+qXEMn1TYpnhj70ojm1jTh8ky9y/
sDyWVnqB9P96tktPILT3ZQWCdB9PX6JhLprJwP0HMYSW0oYk73JI1uAvo6Ht3LUd
BvOIzkiHpyUheoDoum3mi7WDosg7YZsdFZ/ZfIBIXkQjeY9pdrVnqYimaOEOTAhc
oj+LJoQYzgmAWAyDr4EGF2Q6ODt1xbgTEfP7dBoSZkttkaLmZ9GVOxt3XEETZZPV
WBQzEMVoCr6FtTeilLIEj4/duN9DvOUNaBbpIKXUXU0ObzR/5NsSIMvSCqGozndG
/9H4jX3Xj0vM/CebRZnRtSRU/fDkC4r4B1XoVVpZSiNKHp9aJbHWW/Qm2DfY7WSZ
Pqnm7Kt98aZrsQTa3X3Q7wjNRgt26zfsC9o5ulS1hHhactE9wVErqKH0My9YCyLa
EUq29LCIld0/JvnPUAG3iDXDlnNxOBy1809TjRPB3bE50m42Pg2lSMW8YHgBsp4m
UopJu2HZX75Y377xx8c/sdIz4/6vCeEOd47LcjgXhWGnvbqWc9y9sXrPIh6b7mqW
zn+bwDbt1DeAXgANj2B/OUVKQuy+xYSXXe/ZtA7ffL5YTVQzhQtSwTaEDbNmhbiC
2hHaVwXlknD4BXX2frCjaTQq4BGSIk3Z9UF7jB/8oE4SpAyV5PlVY21epdrqWNJN
JpAHcTYlE1Dc92ZbZMarAKUImEZMnEQRkGaqn4Qme9u2aL6MSrF491DeLmPSeRqy
J+IizsvnpfbVPXyBXDeHzsKE9drVZ9GVJ01kCwyZ+TpA+kEvgDUADj0vyiebsLv/
2rfLT3FIFZ0IXGSsin369aTsJt5VFhtwZoCS5gwZNTWa3swTesCQzJgfbB9IUsMg
72hsLgv2BfznJqyCUoPDmeW3UnT2Y1yafJl0KNeFTX09reCQ44I8iQ7PhmH00GPL
N3MdIgqxVurWsQCUjZRjyzf0T3aePtsgx396z3NPTCKAgKZzEKAhlWj/saaMiK9p
a8Pv3H51AsV/EWW8r4mwBsAnCES1uTHeQMCb434xJ0ZrrHoEbfNkqvUZ+t/IQ55m
Xcbqxp3gtD/uYEMbHK8/Zju6gQyJhbKdx0yX4cgBobR2qtSxX9I3GESo7BGDTVlI
MrMYIfZs9WvzULyHqkQpmiDqaKYQN3q4IvWEljhrP7UqeDqeZ3wQpx02iLGQ2Snt
Z6rykqtfE+enHJF29wzzFKh2vIydVt1A+lBN6SyzI5LH8OFeVCzVc6l+XDPIEIws
9XF38aG0jVF1rlMqZ02vOtS3NdOsC+nlRLhOAVD1K3NKD5jOC8rjq+9Uba1MZfEd
wk+9XpBaYrxn0XyqDAgS/KBuWH8RFRRWlvqIDJYTdYvnPBt1UxZdAEUabfzJlo2z
/t+lQ21277zPd3kI1N5KM0zuVZ2+6F7VVB/FXX/A4RSw2k0ACvV7GrEfTppPx8uz
ujIdkef6GTHqoLXFG/1EWrtjGs4JI8nHRurA4I92NukY4D13LJnIXDSR7VXW6RUu
WGIgLuax9bdP2P3yj8RtQb/Fk1g+zMjl9aQjRUx9ZtoB/RXiXdCqEp70xe7EWoME
i5AxegT9ueUBVB2oO3mMIdVfUfQ+xcwD4koWNysXwGdLCCQeiCrZ5lljYz/+jyQJ
dQ6F2WYF6v24TaXygK6Oj80l8f1MGuTC/U262MeFMHficw0QvxgUNYZM5JvLaZSQ

//pragma protect end_data_block
//pragma protect digest_block
QBbsZwXnab9s8sD9B9jM+qwRHOM=
//pragma protect end_digest_block
//pragma protect end_protected
