// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2hAeRyhpE36h4eyRcG6fRX9VZahazIJZZGQjhRSabo9WiiVyr38KPGVTprprCF1l
QeoXpOUFbkH+/INzrzeWvKuR97DMYX0w2a/N4LV0OZG6krpN3StzJnoaeUBXfJOG
MxUSDGe9333LwGO7op/rL+MkgosSo+8E8mmGWS1JoQIWJR7OTsZNRQ==
//pragma protect end_key_block
//pragma protect digest_block
r1sJ6ogq64QlJczyLyXyVHBMyxI=
//pragma protect end_digest_block
//pragma protect data_block
NmdR4FG5XSLKxi2luVyz0TSQdN6RrN5BbTTkDbN3KlFsMh/bTlllfyIhwEqfzghk
/VHFlzeVrt+s/aEb3BH+6FqQbCrHkPkTD2lMysmLDyYfQHrNWFxOc2CAcO+mBqB0
pUlQQ8tkKjdDU7w3GE4QtwLTJplydPoE/Mt3ksmAgGcKV8SGBlB5vY0Vr4uiOLqY
xHwkCzv+VjWUY7PqID+jQE8iPPUGW7IhM4yUvKMI5QudQFnY/ZBiFuqsNdj+70Aw
dhwPyoY5K8xUWS4M38mc5l8M4xtDZ1jktRvBscc4IArUuSrQeq6oRAuMMqgB/nJF
M1K0ILAMcZW+NwI+1lrExaY49cDQWXvr7x0yc5ZKDlCkY6Kqhr8AGXANCt2PO700
lYvjRyOsexqqeZVAS/fxjXAuIxf8zUgeJBm8CLF6P//R7vAgY8iVA6yVPr1N6rxf
T3vhwxmLpZjuLcTDJdCLxycUwVzDznn4pd8oTi/t1wZwriZibVgu9+dWdd6LJLnX
dYug4wezSv4hAH/1LcYFeAtxyHUlyRgiKr9Z5/nHsgXv+zEPqtlBVsOFQV57YFuz
kklbwtG23Y+eLcr591smfrcwq3T1Fz6yL6e1k5MZDuNefz8fG16oIQFasSQzKoTa
X0FJo9sk4SKZGCLpbm0SjO6lq3UF7TYimE8omDW9IUDyE6hM/R3qmh01uO79x7rg
KXdb5qp+pZSWhYfvNEMZsDRwSbe8JUt9gy7QBn8fytW8a2dJT1/HlEbXSdNp2CpB
wjfvFMrNBzA7+MKVh41dK3CIHbit2zzinU/39+F2Sb5OZoAUHqymimP+0X2XNV0Y
mcLU5N77zHJF/otU20gHdT6+0Xf82uHMZpQ5ULPfJ6aA1d2WIrl0HkkUXNA35gND
xVwVvAMrD8HRxvWHnombQP2++R4+kByqHtV8XZ6HKOEuOMjly52orpx3sjofm9zJ
U5x19+/qpEq2IvZyPx/TRQW/EHq0dsi2He9oqNIHuUm4YyDTqVtbBug6oscOtGEY
VRKuBwnOjqdGFsEIMjj1S6yEjM3Q2t5z8dSMfFf71ha9K2Vsm2/hk6da1nUDo0yM
Rf0K/2Al70To7M2MhnIQXGbDs4fUDbdAo2oBdSAIRrccKIePDx6YPK/SkcbwPYau
rcleTQVSQtMuQw1nF3fBU7VKiM9QFEdF0WCPPRrcWuFdp67DhIW76ZTRHaY3DkJU
EOP0Z0NiRi39/Xt4gtk1ZiBZPIYq9BcPIg1KELy4XlLnD5y2BIp0oqj1anAAMCty
er876+ei8EOf1wDGqvjE58Rjkis1MfvmKtPB60vzIYKZK1ipehn2OmgeIT0CuDvI
F/EwdfMXxGEQFONYvsWs3qrJjl8ebVtjR6Dhxa1/FxBLnokkLARr6bQ5IZ/dEj18
GBJAFCnvTotyA82F1QHGzL2TFW1r9ou42J7HnwzhYZlb4MZm5RGLF7PSahXBnhCY
JHq62ltiVWyZONJ8guiH08nvUIm2tjSiA6e1bBtPW1OJeCc9h5CSOtJ07E5bDted
B0iqq0IfeZcXn7P9IjSICCoZ/KV5xuhd/eThbdFSM/EdJPtyvopYfMUHeEbK2yRl
LxmwdjMkY/c6XaUf2cW55C61JyX8w5s8gWOtbmulvvmLZ4HdxMpt0f2gavw9faog
TznmBq4+8XqwTObey3fYCnxXlb2rOXUHktaJyI93YcdSi6V27P7cxL/gUzYcdrY6
wSkuyZHuY+XogjXo3K0KHWbreLJM4EjAyAuxGULUHiotCerU3M8LjX/68900ozIA
WWLnlncSurfgDcCTVD0AE5xk3wY7FDJjcCkK9emCXAnk+bqdiI/7HHo4wdtKx2oi
ievnH3Ds8guT1XL0UyrIiBdj4MRXyw4/lx9DDLThMpAyq157R+RPD3zSsXNrWD4l
qx8wIZa7VQ8Scl4NSyEgBIJXZ5bHIStO7RLNX3AsehZ+CQ0h53G3tbrDx48AdDy6
IYgkmVEXz5TCF8Sv1t8qIdZOomAwbZ5WBTvnQezZk1TPV02kVfu0qSdt8dIWUsoC
R8wBUQBUEnUOOAXP9yx8Px8MHD7CxENhk9eNGnwvJmYKADKWGCAgWjvNDP20flD0
T4LZkdEepkfOVlzOIsmdoR4gKzrBiMcQo8vTjCK9kY5w8cl0PL55vTofHqWDiFIF
QPgCKS6jG2jdzup5eUgK+w1Z42PYw5l/7EkkMjADXCUflrDMBVB53HrJpC4s/c2l
14b4BBu23nnDMSOWtNOHjNKvoXxB1m2sIMkoapCqsyISl9UtwjstweAmUJqeiQU1
pNRavyUC0PTW2pmXMKOgyvwZZ+DB02QYPhEjXLhgtvX30xzcSQTIqqZUFqfBsbjL
2cjOpJZbkA5b7BTEwCIoxDfAP/fhTR53Xsg4d/x+oMQ2d54rdoz2uvt0I4D7bx+b
6TZ/go809Mmf1CmHqkROfYtvF5M0ZPb8n8TlRG5To5/T0ckt4IC1yrhiyDHhMKRx
8Dc5m9q2mi9cSHvQRsLjHe0+Gl9AnoJZ8RH7RHHfjwReo5Y2FyC/oOgiob6MgEyx
1pgAo963e4//G0RLS6GGA3W0gz1+oElruWyi385IUM7YCXLBdSbzk9MIdYOnvxx3
/JVSBGqVneXOkP4BM8ICF4CfEbpxfJmmfh5JPWK/tD+I2SJhvx1CVvnDXh+uMn/1
FmI4+nLJwVT1o+DmMbV5vbxi4Yq/VMkwNoDdQgoQ94mlcRz14x8uj3S5VzWHeH6/
jm6BX6QsmkPxEEY5Vny+oIy/rNpopRfsetGBCsR17jcdfeKonQ3CpeLspKAGVo4Z
Te1vC/klTMFwhCOSJNhYsutD15t3H3LavpSKWSWGqVGGeUD+gf05/VdeDY/Wiub2
pMQZcrdtzpEzcuduIGMq3/dRRHDcHK2iR1AE7nju26DSIByLbm9ezGQkY/HYk7xc
+beNbZUFx/Fj+8Txo26LZDaEul6gSIuJrW+y3JUu30Yttw6b2cHhPqXoj3+EqYGW
5oImVYoP3/hPZNDWxTZJzl3Eh97CITzjg02loikoEVinLfhtkrQxvmpNjBIG5IMU
fpd4qySeN2kb1979DerYgm/ey8McOVCcOzQSth6s2XOKD5RrT2uD4er8QmbI4RpW
FcDbXTWzpNsd8wmXgSxFT732lP1pXeyxhux+IDdZOrMFSzlHy3VSzPZOX/lMPlO2
2awCBA5qZPPFOP4u7nmexvVjhlsbeg8tjyXWkOiaP7na05kqM4Q5WmmwVO3pOybZ
GOFJI4AB5STRPOBHWbrmcMxqa0WdaZ7vBGuuyOReTjluNbVWETfvUcy/TXyIWnuI
BY31S/D2sthyV4UTHHRwb9g+bxxKjMUIOjZ6FEmmJL54xIQNpeWbDTNpwr1aDLwh
1Eeqwh0mTuQGQO6pQzCN5Xx3z7rw7ZeM4Zs3SRLL9DnnXgKTMxbUo7qdJ6f1TjG2
tsNdSKaip11sSEGLQQxQFMiYQJThq/G2KgW2/y9zxOvt6iGtkpi6zSlT1BBfTL2B
WPvlKsI1CYNnOXv24TlUXNYw7E3YjYXHdWi4WSXbqtBqp+NdTmy7P/u3ILZ8NVmU
R3wXnO0T0To/9lIg7hYWNCVfodv1KrZFh1ed+QG8xcK82AMkyUBIAVEKxxs9X3b5
cJRtnZDB0iy/zdHN+ZayB5Y6rl2CUwJCOJU8Og26H2g059VUgpia47lKKqJu7eAZ
9naEbq5wr6uYdYbpVvstYqp93YMscRTucX4tmObyd4AknmYlmhlLQohleL+LsiKA
H4UBXwNHo9G0hSTxByM+yDye6VYJSDwpRMoQn9FbpWnUQTaN4egE54IxCjLOILeU
KxDENm7ZdJwCDgdcMIgjpEdhpTspSexk4nPlVWCf/hECCgK6qsQhi7akfhnhWyaX
6ClF1SHj3j5XEEZEc3tdrrQKepOgL7+QxT8q7UzrTefJk/EsxgitXD7GpbZ5v+Vt
Mbin3ph07HT1pE5/V6Sqh6JdOzn1HwSiIMWuuM+UGYmLCV9yQkjz0qw6J2XcHOCh
xIa3X2g5nWThH2lePO38HsTJYRl8bQ026ii3u38CrTBnn3J6qFWFzNy3kCmpb8Vz
lNCFOS++zq+al7afYtMzAKDAB9EuASXfLFNIZvk3f9ePQcdTCehTHPZ/QF7ujry+
f8r56M4KKzGCg9wsGPqow5M2YX1vbd5vPG1GUchh8smndcAY/CcycYp2pKMaMUMV
ExKyRpBFVRWEU4g4yHhNCuj4BLZlYz+D04N8Uvl/+JdbGnN1PUsoBRM4kl0UGdTi
1enht4xrTayACGk3IVIo80q8P4ss3BSmoIyIgKUH6X9P3OCgKa4pncE4XHoLa2es
+cTgaYTHxZH9IvhCtlVml9bl4riSWzXbNra3k85nNFdWuRL93WC5FjBIpwmZl1tG
ZxqXf32qbpIeoCmlUZuloNB9IiyXj51hQPpqhIPeZ1mWkcH6zIRhcNwMaW1j2k6q
95LKJ9Pt4EZ5g8VQvmjMhM5HBZx2VN7eSMrv+YO4RHN0JvTTDDnLJWAjKpZTiQU4
qiuAtl5EdhrMwC08p9uMyC8N7rge91LPGkRdP5aw4mRf7jvpTSxRFSRGP1PHa6hD
MDxE6JSUhNaQ2NwQhjFXiAUJbV2Y+HboagAHt+O9kcCVyGl2XS/lBeYOmLatQWd6
8HM59d4vXZb+Nhv076wPA/oC+/8dywjQUSTJFRAZLUOfggZ89UrZL0GvUf6YCYQP
RMZK1r3x3HIqAV5k82MklQp6c87AgQN5yiXm3AQEZAufNsYl8YZBP76YtHWPXxS4
dLqecVyGatURBlcg2xTP4ixitkGq6Pi9HTnyoHg21hDXQtqiU9fitpk0+PGyhQ/R
Mq+2OU/Ev6+EJqCIr811wmaQbetimfdWnq2MZdmA1BsfyuKF3HtpAGpXl00pBZw1
G4rpd3ntJ+/CzpqahnpbIwIinQKzin+0K5BxwVtpDkjY6VmxYodlpW1Eui3pW35n
MgSzhinaap7DC0m31fBbgJpvQvwpx1fWl5OygZOekM3efJc3cpTzJxQChH3/BwlY
Gl0Ni77QddpWNkkyzmj9kegQk+6Md4ZEC1qtFz6iWn0LStbcltzd2z0N12u8L9Aj
+xmac1HeaVkOi1ZuWDtRyOp5brZwcNTtHGglQCiZMfdkLgFgU0gikouMuAph4V/0
Kq3SiBtkGNr4rP1k9PUQnHPzxwjGY0EJNYc1jA3gzBU9VQfum4wbVxvP/IQLR4gx
8C/85vYU3kJdWjQRFyvygYMiwSJyWVcMyV3RVCZzsYyeqnaLpxirI95/KAwBailm
g0hEEZWYvf7df8kd/uKq5B+aZN0wZxbyf11sauE14mKctdt1mhpg4mdrb5+RZU25
8wdGw3Cay6HZdkqHekdCpyeOaMqvC5dqiHu+tviQ5oBuKC3q86pbjjknlHMwYMNA
ye497epMND6ODCPFkn7ziKWrJAb3E/3OKfo3p30kFQ+9adnMtIgiGgMRjtRmVcnM
BrexbQifbxXhFj57ulLTmAfvtTdRrhpO1bB8Lehkc5UBIkjDXtEs599khIvMEvgr
WWPP2oRKkNIyC5N/2atZLx7bSbQXNkdSkVA7F/4crltJNj+k2BJvPAN7oK7ppwyV
U2hHv0aAdvdTW5uOKxg7OxEk1Pmn5rePzE3kWanlksUSrMeV4cUpZLbIn/s1Y0xA
FC0awV8UaxkVwH1rDv0TJGKL9gVH3br/6C9KqH1PNZeZnG6HpYnI1xBH5a9lHDZt
TMshNvTBiCQvcYsUFy/MDe8R1fLA8QTN8+4/H+YO3f/wg7PbwcqoGjPh6pTQwCYw
obGCxhEq4s/aYb1caTS7MInxgC4SuQpd7iZrxp1tUv6U9iQOwPuKf7k9ljyPdHDC
P4g+5PD/ZS17Yj8rR6pztrg4RGpDNaypqSbaV1gOAjbqfbkcdA0v6mZnEog57+gt
ed0i96mU7n1/Nr3YH4Xct1WTlhxHQ+IIEaWk1pduo2AVVSwOH2+Uq2+/NhLXvdLm
hXLjaNb3pODXM3UtYAmdV5bS+kMYJZggvJTKWEGLNug1MkDarJkxpOHgx8hJcVc9
mTp68Q+fc6aYBNLk4u6N/grHTcjBFxK4m35+9OEC6O1bvH+CEaReUvnMIAJydPX+
nw5ZQdnlLD0eV5g0EEmgw54UtbktJeeg8Tybpa4z75BaI6Z66qXilOs6qkc835pP
wGsKoWD9+SRZBhIVc8eb4vwIjMtV+4J+GnEPjSsrTJWXSNM3zwqvLVDf1ozbT8aC
ksOmstXRQU1oMtQN0uBZxnrqf8W1qI3DbV1PW9s8pXEbznhXprebmIP1gMXpYIuh
DkHzapi8RLd5B9JjWzVcn1H3cNaYFzkG4olhj3ssUUYzD447LkBbh3xQlUswHOoY
IhrknBYOx1LsuGTzjymq2C3O9yWBc3WwRqVr0RIgObLvHooLmMd19Ja3DH8uJuTf
mgPazMlSqnzuL97ZW8ljT/80Syi2A56ZcTrsN/OHdJKlsLjIzWOP+/0EleYwsLXT
vy9Soe83da4dyznahuE8YZHGWu7njzhBF52rmdKbYSm5IO/iKjvN0BHbDTsN4NJG
aDzZPTNXVXpnmgdii+NVvho75Z+6hnkf5w5mONZo32mwuCEsOwUjAZ3CQAivM7II
IWqWjtZszFAR1/tk0XkCwoUMur4E2abMA4l6JBZjNtNASL5P+vIUI5tTNodpQqni
hb66qUIMXRcl13zZuueoM5xNyUIHen3g77uq2JrboGh/TZ2HwTchKMqeuuPH9bf5
gFgyjl7hUhwSRzZBlWeBuBXj6kmVbRSDkULMSPTbTl1dFj6LRFuQogxt6jXbYP8A
B9+tFYddpZqCy/zKmwOhYzh3QI3IXJy0usyQuTpaFg72+ZK69AoK92j8adwiP6OG
ldROn6xDosteh1Ks3e3Vi4pZTqqXDDfPNBi/h6PfPABvq+jdfNcyX3MrnC60LQtm
3r5kaHb7v1bgh+O9QgyVS7N/BGffedJGbFNcGhLBghVIeFEj+DSXFokjoWiLw7fF
qU9yXBg8RykjA4vE48MMQOdQ43zLq877fUFQtNd1yEA4QXyOjkgLOeHnms2Vc8jz
UUFhVRMnvn2pbsgpKM1jvhQL4WMzP9QNvgolb7cWJtXEyl4Tl5yRYCjo1UXNbS/Y
LbOo9TFrgcWhfzZlPYfTdKWjaMki6hYQO41oWnpBkDNRY5cI7lw07bvybew5vArQ
+1ZA0MON4LTSPOVexuHQ9jxViFZZAjYRAGKtb4YxEgCGTPrE5801wkJco60N9hVS
0n0U59ZzqaA2CZ+KK8TsBB2QEFhaprUeFV0OHyR54gnbZ8HJPaLenBhKaSpEOT5J
2vGmDT22LNtzj0yz65omnfGh8o0eLN7OgWTQjnAbVu2Yuh+JefAnVLJy00eyVFHM
0nM1bup+0Y9OyKulzkfyRbLPwfF+pn2qnjzpKSVKIyxzZn799zJ1fK8CQJNd0+Zc
g4Js90pfFSwLsMJxa6K9NeklsZzYAj1t4jx5VzWVXm5cfAjF/CJKQCMGt2o8Odqj
BBqxeF+pZzYXfE7m8D2Dg6ZC/+WThelVQ/kesgw/S4sPjF7/mil1QN7QiwVSSmZR
9iDtqhqOahEyd45cOCTdM8dMVhz9ES4JgAkTHcveKvEQ20IzNh2eP5HxwfbeW1Vp
xoHuXCErL5UoTV+rlViJ0RTCn+GpdYiAjGNxxxYyj82+xEsF8TB4skcGg6fnAbZR
+kZ4AN49N74o0OsmwYM7e6qaEmqU42FZXIUBx1TPv3/kknYf7NbL2CINjECy2vh+
pMPguXRfw3edWLjbJQL92B1VR+/iqpigbHXb5mAIFUiDypeWAt0texSYK2a+npaa
qQI5nWmEDHZ96OvgValsgZ7NHvYpNGD4MQCn4PQ6lXiJ7Ch883XWHdIxM8SGpUVz
bJ6M4vyNU6N5tVKFIEGj87AaPZ/EEXtDc30Q1a0iXOEbVmGCmLozIMNVx3m5fyiS
8X5yjN9FI+xdb518FBkVRLBIEnYR72/bhtbjl8prDNG1NbN+Mc5kLFp7Ae1jnttD
rwVvtTpMATwauYbpPn+V208ICJZC8QKHufeP+1B51EU5CUB7zsOJALo2JniJObIR
sZD/x7bgRy409/IUFszV0z1aRwFSWEEPqtXSs8Orb3LTPdF2oh3aCATnKMHzB3LW
tmRA6xi8S13EeXYC2//fcYhfEzc/TkJII5Jc2E4F9QsgWNqRZX4ZX076yXJ0fMzO
pH+xb6BEwilbzvSbBZNLqUahJmdmHF7r5cJBUh+fppNXZwJ7YiyPLqQpBD+u8KGm
uOheSwQKt361c1uVNUXAchDY6TlybPdiJGqgMWIpdseHl0eSVmkzaWy7KLQAcdet
DfsY3xRPdoycz3NUcvO92oiLc93E3CWbhht4V+ugWzIeBkMSmZQv8xA4EplvWgAu
SiOEqf+IoIBZ5qpTm9EdCJFiDdPuclf/r4aWp2URMn37ViZIKM+C/evPIOAEVDjG
Etz9JvjqMoZn7G6VA42EkgjSeFL+6qyh9E1lQTkcyvyZZp0Q33ZzXsjPo8gHKjps
llLU0YNW92T/4SxW5jAjaNeBdjPxCCuTMXnlykGnp5ho0ESHK6D4PCGc4snXvyFO
NheZI/ZlMoW7dhk2Q8NAAXjYSw9ihhmv/fdEFMF8LHacAGqwMNYyzj2K5oeVMhdI
kX/s0hPCwoeozShcfj8JalArdKlypjRYXxBle95NYiUoflQUkkSQIE1V9zkyQJ5Q
tKt819D4jHdSvC7JD0z8ZcqxyIKuj6b5zw3307J8WcpqeJj/PGN4aUL2Ijqv3Yga
tbYUpQSlb4zQ4bOSUGsWKCYbCwyKxxLlCP5HEnRJFSPykTublAfNWyiYCSqEO6Hd
MPL2cnlPBGqSWaZBt6fHca9PW0AdPCnqbaUl1xbDodwHSLBo6a0CGU6KgqxwHdhb
aY9hBb4XXUF90uUH9CV3xAi7NCMXFTrR8vUWN/fwjcWx2t4pfBpzfmeJfRPeh32B
9G8iNa7ted63iyuUAfmgPgJiyDw2BrdbF1WZgTLJda3wgWTuK0gPigFB6GZrdXS5
+JVcnlg4gNBUj9WGNqJGOXmsaIte6u6hiUuL2CDhhBdSh4fzHsvZq6BoTq2W5E5f
Z7uWyxKA+8GA7GDEzXVNsVHYq1+LyUmm56Zf6bfdNSklvUZ2MdIiiYJY5Jg80vOq
gHuI3HzaMA6aDGBDF1IXiMvMfZVrEO80uOMBzU/pTBuV8huxmFQ5XUvF+ICl+321
u/zIpF17wjSaMhcAmEoM06uZn4yQdni+rvpNL/Va/4QVa+OfINWJ7FLmyEgEi0+l
qHJ3jbhiI+iva3omtO2/hquDKEYA0ePSpmu6K5FF0YqKfiVsnMHL41gqTnG0GiqD
3KdXzJqC6yX61pJis+kIs6xWHOH2UsIL0ImtDBdL+u/mJnqiQDBuCRqWwBeMcsZe
DCcnbhSvbtR9AIEuUylZHuDp1nsAu5eSaKHdlW1Rs/sCxkdpX6+JBh8axJYPdnqw
utO4hHoLPZkNaHcrtiXWl5RhV0i/bir42Tm56DpdtmlpTMbjOIxk7bBlDKK+ovy7
KQs9oFzb8CjG4SH2M4Vuqe6ROUB4k3EyYAHO0hbi8aOABLVE6UXlEvBSbny7zRmJ
XZ+SMca2znm21aYIvMlCu/32NmhLX0MkInu1dBQamGMAK3j+Tzm1oMvCKAUcdTzQ
hQ+baXtmoQdoM0QHcO2LVrr74vixV1MCj8q1M5WP+aFnYXEPa7XNpWs53JSmF0fJ
fTYwpXxI+MsUCEtDYCvlArxx2bhujXRebbkVtbeVkH9ybBm9waqR2XkPyLtJbMIt
xWjcL2j2tqh90syZgFmSXLHsIe4XZCIgSlBuKrEK1DrJFyBv1vskzDLssIiy5E9H
ZvWtAC28iNfjs0/pyfwm4gXk+vWKcz9fkaDkad1o91qh64ZFTeKa66rrufL9qXfP
kA9isi36oqWQwbWCDstI3ox/jrZfe9Z8ab8Omvqkh5UOtJE9OCDpzo4MDN3gogcZ
qHKiYJcex5FuhFR31FFyLBU36RLZegujDOU/tLa+QbMtfgzO6PimCAf8XriwfhGZ
/gm8t7UiuaVYBTMkD/7lQzxvZQo9Gbb1mFjX/AuQFll4FBufEJlyMBSVRULNdNWi
R7WT8LzHVMmq1QYDSmBH2rw8rpZZVMmpgDMbSoCUXxVRfP1Uh1yzoDtkg/OclJWQ
YUMFFS33mxWVKGu4mnHgq6FYx5ZmECcaMV27yV0hJ2NY3c0snIjbZ3QZC6e4b/I1
FTaonIv42CJTGsYAFf3uYETC1I45469hDLLp0KBNFNDF4zJSQ8x7GaOnnLqf9c/l
dFw0Ut3w2gf/BUgPg4TdVvLj3zFW3+tMEsCfAulUIlICUVeFbiDVGh+fBK5lq40C
JSHLhRFRCn4f9txHhFRSLzkZ3l8INpKFhZA1QaCuDfWx9LgiENzvBFgnRQBKbcdY
ZSDSxA16bK0kjy9cKDYEnre3OiL79JklQ3e7DqyrahOolcbYWpr1P4AFJ0kawGJk
yMu4p5HYsEmzknmRnTjaQ3n0hY/deSlbClNROEJClyBvYbKCakwHdzK3nXbsZdnv
qGSMJi5CrxlhGkGr5wTvNOYo34IuEvfUjCBYzxS8MSIMs8GZYOEyCmDt+v+1nzv/
DRnwZQEKK9RRxLBqyH7KeMAGvaay4/YpfVlykGXyBuSfM3j7BGy1cLOk4O8f2Psz
6dR4eqfRCVWJlA9KYnOofKZUbjffVHgjx1mW2dgfURY3E+Py0bw83jFgEODyCrQ5
9QFn9gvqVFHr0jFhaAvHb4d+lKpD/ieZpHMHcKzcpdAMYYVkupu4Xo+lsrvx0KXb
pGp/5byJvT8gWOtGQoJMCdJaVYEvRFWkKjXTFMjG+ym9y7KinOrFG1Fp4e0e3IP4
WFhHEqwUJDYFM+SwZ02mNIAYaKrAVVbSJFMXia5VgPO+jxg0gTF5BcIGPMy+x7r5
T8QQoj7TQG3IcWB0KxiCJjDJn2IUj5zrG4I1qFotVQ5m52mvGbfiMm/9VhKxbeOm
eexWEIJoKiSlKI16JkGbpllJT8DgrvPMQPinU4jSve3DpgWMm97mNPjkngtuXjIY
i5Q8tYr3IET4TUAVNVW8zlc5jaR9+a25I/FtM4WNWjiV3jxcX3d78g28rVAPagkL
xX6oIlrcXhqmuP1FJ/WUMMH8WxnNs62E5amtLOSbz2Lki2h/AIsiHr+P6S1OE8NX
aRO20esI6yZCaSUVyMpnt+017amXd41sfvTkD7zZNKsKcxQscYMRs+15qdnIjowP
05fGQcW+eK+iebJ29Es+N+uGJeQQMAY9Ge/tRWlmXfbIpBkYlENFfQY+ULF0zp4V
Yglt2W0bX4FpahRCN0Gdq/SRD+1d2iTH8QD7xDO/ThwEfaRYtcBfr7RRyRtkUA33
SX2TNMlim0UrfrmvlX9PdSeNEpdKaOCeleY9fMVzu+ntZcGy5xSlb1zVGbN4jHR1
MJH/sCxKdnt9G9asoD53vfwMxRHxftteLW18CE6H3mBSyanRO2HVM/S7dM9xRmpJ
I9q36zSUVg0v+3V0IcOv6GYK1QGyQRpeB1lq/5doK8cPUd8O0VhAv02q3OrJTKe4
Ko2mJlVsCS6HETnNZ+I187RDKV4aAA+CQ7Olq3dmrvMqr1A3JZplhiUetgutyUzr
xmkU3G7pcHPl8DQ7poLKvv3zOuaR1iMh3WRcJ9TFf+1BLYyCKqRyEMSsJ7btIFbl
X9JqiTYc4nt9Nfsz6vGGF8FeEKH3xxzI1S1P8+LQDGF0ZVuI+aVBASOXSNirgKzJ
uuRqcXHC5V07sjURkNO6yl3JgV5dpugO1vPyc6xF9KshgSbZkz4p1IlbDIA5cv1l
XKkuQeJu/v+0EfSsenX0HdB7StvvgVndvoG63SK/053eRJvXWsn+xrbN2Ieg3lGo
o7SG1sVWA7feelEAxJONC/cMLZjd1wmQT7kvR0imhzYzVs0gbzwM5ons9FHQgS8l
FgKSHTQQ+7weHx5Qeyb5wSj6ZBCDvjGbmc7HN8SqDX+pL3iRb9TZw7m8riDuo+GR
YOGhGjP8CwDmuoqjILzstdumMNQrwXLgi88Rpo1CyUAfeeG9l75yyl7RiKHeTMfv
qfSdVxkbVMUj4/uOwxwLzagDAM9lF55WVNrUGNfGTad35Iy7DDUVXyKyOseAIVHF
2JseSgyyZOnvxAysk3qzpYfckyjOs4xuOlDRsAWM6fYWpgZFCaNWDcXMWaoJfhEk
hBUIOiSEI4zeEcrGxdpO3Jlu8UM9Lg2u3/NIX3tgIxTQZT4D/3P8ClLw4KgPXI4C
jfFVqKtMYgwoc5+j4kFij8n8ocwxlDK38Mot2CxfktKrXavd1e49WLINR9yrhF8p
fMDY4XD0ldWTRtpu9H3DeMU6hCkAsaBIqQjdaHJc4wUuf5qxWG37GTv+QAnx04yN
PBGn+EbPB4Lhhyuk0RkKmtD+rvgle+PLGCtQseH62G3XTcnYr89eoI+IKMCekNYV
5AliZemuTtQDbRk6kpRnSu+FtUJBBf6UkPD0CL5cSYnh7y/v4MVhlWXdYf2d7GTk
JP2IDg8pnWNbaDFCTbMdQnFHUiB+4JAroSv5M45TX7KhJAkIurKCk5YeyH9jytE1
voNeLCKbZepeXkJ6XJoxgwlNvgrFeBjh0OrOfA8JHoY4VJhcvUixp/fSvdjfvRnH
3AlIuvrtAjvN6aQ7nev4XmjdDn8EFEq5cu+hwgl7nTWl3wysurPkPZL3fsQq+b/S
/2YJvbuaq2LI6q/5ey3b/uGmKQO5MceSCGHvbainAp+M506KBnBYl57jTlCQxI+A
6DL+MkuczCoAU5C9W1k/JcWsmWP2jhEXDlNEVZP8ZoJULPmtzkoLlmS9lRWhDBtu
ybBgczkzAlbIaPeFK3JElcCJseJCKlRvMvzyQ4TH8/dx0za4WdFnTiO0EBYnJh95
FWO3A6qqlRDbA3/V9heOPUKfMCeHtpI/RfaXSNRrsBMh2GoOBBgRvGOYhLAmarOj
zPwu/bWrVS1pN0f3hN2yhf7nBmcj1Op3rz7TDIuB+Wu0iJ7jQV762A8Rf0mBDXub
6PitHGIW09X7dJhIU9arb26OBdDz2DSqHionlZ5vVM3gyGFsvlRD/Rz54Yl5OzFQ
VD7dpJeJqROcSco9NUlpcCzbrwfju9gA+vosKZLUICsyLc3/jYC9W8TEUwCYC0WN
Xf+GmJbkJUDabO/0PL6FdUJBi/N/ld/fa/eSA4Ab/2ARRAfqziLN90pFWZNZhVZa
sadfEl5pAEMqpEi+978JtitgmvrAX0wfMHu4wzdUzg/1OPUBvMIS0lalgzMBqsyl
2ZfXwpFDYzugli3PyjGrUabO80GTlsuG5W5FQurVn+3cKTZVzXxf888vpH8kLpeb
GN1a019UGSmjXuYjZmMy5E5Y4MERipdcrJHPG4vwbIe8q/p9pbPfbEX0Zso6KqEr
cChoc2akbga+4mX04OFeDIxLsRgA7a+7jmo4QgQrQAXfQbW9+JMYOrZsfTQOaI10
8fhYwlkxutGbg3yPEpQiuUQgjHeC5vJYRA9m84SSd1ykCTzGVOZW4pNQkWJwowbl
s2fUvspuWekfOW9nr/D96AdWxblvxdb3QHB72J1YfIe6uNWJSU14GQvF8DwcZIaf
b+8rvY/reOzPvgWQ2CzwQekUcFvuUNfXTc4RAYQWEqwTsue0qgKlJyzvUUhzJ98Z
iAXsrP8d4UwOd4Lf8vkpoUABiLp53xbE4t7TxUOT3xK/RwhAhFTuLHhpwStmGHz6
7dXvEF0a+Ri890jS1zOZbmKmS+HrZP5o5/gukiZfbT+kX+bc9xGUCja3AU3/EjYA
KdEEKCU62GrNWu0JP+AZib2/IEt8uop29MSW33M60btoJE1LT+5x0F1WWyyMft+I
AXTkeA8YN+ElW89FbTfahpfaleKTAXRadQ3y1qge6JYFa5dxmpsHpUG/O3A5dMdc
VN3aBrfR/PKhwdPoRjIFP4tGgwF0RIVU1A1xhtYdB5oyptbt2XBzeRcjzFsoOEXv
ekPmlQf+2j965OM5PNj0+RDoDu1Z85lMdEnHekkec9MrozpkgPh1znpC8xGzZOWD
iZfqOBUbceebH6O3F30U1w9FRYfA//9nBDa5vF+RHhPcgeLx6UrxeCM0oZktxLEX
HmJc3bRhsg3EBkyQreZQ9kpYpBwMTaK+xJc8ZwD/4ZM1Tbyg9DDsJ8m9WEcvXttg
f/JS7+UNfnQBtZMG49NkGc7mDl7sO6kuLi88qyeqGpaNhbzE/0/pg8WvCxz1pS8d
ucLGLezgoH3+KYpFHYXcEWpwFmRbIk+YWusNKMoIu/VSsXDEVoX4gGpj0fAMmn5E
TdOAs6kDyYxnN3aCBPqzDyFZcXDKtfyaA3rrozD5aeJIiajKO7t/6LchynWzpVul
aBs9V+HT4t7XNDqR4FJJZBn9ozaVIVDo7xL6ccTgYakKtuNQQPBANUxcQp4BxK+d
rcyW+CNgAg/8f1Z6ATvWaR535/H0jWiQ7TsmoR0I9Wqkrn0frZn5F5DT3k2vrp8j
A2EAMQfbbUXevcu80sINhHNfBhWs0zHzIDJheswjPHM8xv+M/zEM7BJKo+ye088W
7QLn0N8IU1Q08XPla5h7jd/wLJDmAD6rnwSfH0iN58NrkRaAkJI4e/AgExy1oEQQ
s1lqboDdSpU2zbYBNBl1OtnziGr94QHkw5m874KP4o9r6vYtm/ZKBmJHLc+tC/4T
coSLl8lUUmLVSHOSofi5chANZ4k7RcAMtRp3YTHI/+AmwilKfwfxD6lKsa6ESnL1
/P0Z4kb5uRSjUKMzNCkaHBU8OpEc5FgMPFmfA4lk7TLe99M+2ZAmMZrl9/PJZFdH
+uE8IkKn+fu5QBBFp8NLoP7/9s+5ZHGwG37tDDtziQfk0Wc37vCMBVjZpI8AVvAw
RNR/NeoQy2C6jWS7vf5LFzhawo7rOmiIUUT3gKWTm3/Rh+ApmqinNfoiVJ425Mjt
OpM5wjQVjncAwcQTxz5GnZbFt4PAmV5toKx64kziYN3zy4PelPG1L0LM6oZmuepT
v/K8iEdeGcaqH7T6xS9cZlk4wvfgDug7nuKp9y3VtTpmPTDB1UrOLrjY4NrC33MO
t20WbRSPSS/7WmWO1/xBdQQoaLER/A2yyL1slPcXwBLkcJ39bEtQysw4Irm8/EeH
PrpGwLBn3uYrYVZHtrSY5UjnwZ0jALPX44zYttwyah2cCPfWB5d4Me5wX2mlVIbF
mPiNTtioLXIH169Q6Uh30UICFo2c7vIP4aDKoK+V3p7za4AiX7KDku5DwXwNjByN
DLb6FxFi5IgFWWWuzUwt1KuVfg5Bt1aghIR1SPLdo/gr2JS+YwaZokPVNRQuym4b
c5786cIDOIjINQH13aQmC8k6NGniwf1jlq6adsfr4CnEzPAdXSj6/CwgolZH18u6
CbXG0KAs5HbkSTYwXBh2b0lAq/mlAlk8IC5A43Ih7IQxBF5JV1wJwlXwGggMnavz
cbFS+FqMSRcpV5RtekL4yjzz9JIkMGBMuwoNcrBYJAYzcfYZ6FdafAKI9/2LHIlM
FM29stam6BLxqEUfW2+ZZvHWZ3RwZ/+fPP6/HbPUWAu4YNQn/9r2S6YpyiJ2h7Od
vot/48dzVgfZi3OmgUdTAAQHw/GWEJ1HfmX5hbjyNFBxmScDcQpw+sCBUtWbyflJ
gligiGPGNQmhgoYMjUld2OytshlHGs1ODNSpLoYqvoiQzHqwbG3Op8VIk/6Mhf/z
1cyU0oqafXY7LCMZWN2t6FfcvQqHVdF94RDPK/YVRDr1TLbTQ71g5U/zogH/kR73
9XD4YOrZMj47E7EcgBlOmvd8JPjc+dclM8FkLPTXGUfeWyAeORPogQowENWXYZfZ
zviXORO4/uDw4tKoe/AIXXnDfssDoP9Zo+tKkV2AhLvR9LEMKXF7UJ/MRy+D/hxy
95WV2IPx9XcVvtRbcfoOI3MxEcjtXLoNnxjyThqymYfKAoRjgp1RkMiNZ9lt5vDP
DB0nEVxF1iwugYeld80uiOVvJFxq1WPqAKlFp20E/bVPfO17Hb7DLDPzuj2S0l1i
K3+Kdn+teZJNCGzBF2vMeSzzK5VmwIdLrznjul+ywWg6VKk8/mxLfLtKiVZgdOw+
TkeFkCxIRhkL7diHgp/gGMKWoIgvLVnZUXKlSPN+a3PTR26UJJ8n+P0Fss5PU+/W
OLZblXPFwh69pma1fDWoniUlm9TLlF5GROaee5P8Hwj49i8QpFSue0T1u0yaUbbF
lFnRsSjK8q6I5Rt3z5Q7WhzQzRGcjS2nLa92hCYBYFp478LOGWGD8div8Alotn6K
jLId060OuUu9hLYk0cSEsup6NJ22lcvCZVQiAmL2UoWXt1nYy/xQIJUMfJhAzh1p
0wrPo2N8T8oLsjQ74Ga5GKDIzA0k+CVlkgD2tpfrLJYingGZ6H4xv9nIUR5BLgXP
YFqVqDS5INLTXc8DuvOoblOwF9RMVCW2UPIAy5YD54OuV3URN6RVEzIN8dP76Pmw
ZRY5rlikHPYn3hbQAtehBATRUfNHzHscgo02r84r5ww9F0D+ATwAIP6xQCGEx1EV
5co2ZH0bLrU8hF9II43M1n0GkwvQ3py51WpJh9kbMvlaEUCmd2+UROX+vy0eNnEF
J9E3pxMbK29Z/yZCjA/94FtQ/ivtniQcsMjt4+j+6o/Fde0OwiWeAG4mE4ryAoAf
EbhG3vlw+JQYX3ez+5RN0UmxCpXMOXMLqqb0hgquPViHyTGfwRw+V0HDld5SNhvV
SLzGC4n9ES4adK+ETxJhexVnvjT1UjWyiQaJb7kl9hIhc/Yb6AWycU7NM8QB5fm/
d/7cbz+eBPA6lTykPFOZ9h9QK1T7wpYCQRSVpFKmeZzMr6+e/1/mVJj0voBESw4l
EQb8ezTyXP5ls/WKPDsKvJjxuIdpYrXyXqdYbZiLcHMWuRWXlPo86eXrVEXshB2W
w9Ac0a8Tuu9XebLOEDWSmj7ySz8kqgqrOgdxiekXx3uFoc1K29FuBLoHTrN2JY0v
BvxA5b3jLMYvmaiaqbe7o1qYomh+4+Ux7x2+ui1olaHkT5LqDb1FnGZlgZJcdM6n
QmjSVV1ZYeRhiQ/io9SqSbp5mvJ6rHjvcIGBHycu7kXooRUH79DQ5X4LLwVzBYis
/7Zqn76iaM9YorGejLfHkz19qjgsbN2NwAFslkr/1yhli/eqB54BbzW3trJ0B0xT
X0m9I3ALQRZ8VCbdrNTX7BbAUjWHFIKkboVfh7p2hG8V+7Fg3SXTi4A6qyAvFN3j
+oVZD4WRyjXkcHJ6JCaV6PQbcLi6RvT2VjDKT0yt22VnOgx9PQ/N6K/uyEcI8oZs
vS53+PJHGhPoeambHa4D5dxZSdeROABGrUgHd583WK42hzNNaUzEhnzR/P3G1lzC
ovhSlto6EHzJwXnJMZN0DzaSTgBb2dCD5dprWKG4iTXu+3l5KDZNrzrmU/XUTQEd
YLQ8/5DVymFeOMNSRCfd8gVBUqB3y9BJG7yzzRkNTp4yEoaWkTezVOwMlt5LnGL1
lEXytfXL62+qiMcV7p1sViGsvXusygKKeS+wv5K4IlIXtuEVtDRTFgjSKpm1zYOK
iu3O95zvZPr26xsy0ZgX7160GHgRQwZaPpnsG1gVu5DfNtxYmWBMK5eikdq6hPIh
uYKtJIwem0RUPazEGnZnibZzj2a1lXcI7JzGyOXkILeE27u7XFOnJg4Etiwu8yUi
e9lDIAJPLhKLDNq9r4M5rIAibaFVE0hDO2TVj0NDugXBaC6nfkx7TVFWLrvPXYlJ
SeO0fNeUNWb+8Q33n3INw0tV+ixp9MEbXX5QlX4kuxq8BmvpR1NKK+ifG4TP9K/W
yv+TiJT6P4Qe044zsiedB0wFYwTs6dZ6lG+YaDPEClsccvTap0z906HDVvqRYgjd
Bmi4VWd/KCQZqfZ4yosUpu05DsKf+6RDz3OPfs0VuVOcma/xK7f4VMYKPfmFvCVW
wrLxnzLNufIB87ZNB3VLHzf7mu2+nw6wR5Wu8twFC3pWjlXevcPNWPpSjZEY14bM
8EKRnMAvPXz7jhiZlSBhsmOyW43+gneybxFcoxfWkj0kNMvrTARlmDpxwBMElQLD
VGQlthZPtEuM8lpOLDcJgbeuuRV4ScPg7DwgEPHplNctoJcE7E5k1r1WfNXx/URC
4+fU95X9xUmCz+dJ647JwxaZ/M431YXCSjWfUDJA2wmtekqY9A2NC1IJcfJJc5cs
2ukprqROF7Tnb5GuM9XddbYpRkeE223J1rNwDpzzvPVsBQIZNmz7FCuB4fD0CGQX
JQD5Ile5hVSGYxlk8QLZeMjj1yzi8jmxRiC6Nb0ukj8rMcF8CKkWZ9fpaFPBgE+4
YgZgN+eEpTgqmDGBvUwx2qTRaBwI6z0zAtq1MdGqvo6dBeTecMHU+0nwkvTpb6oC
Tmz9VnhjiHVodO+wTMceLaKl/mqrCWvj9gXmidJlP3F/zFO/vKRiu1DQJ6KM2knG
mKTunako/2sTXwB2MrJIaplaa6mt9MqZ89mN6i5ubNN3iiQyBL8zFX2O3OK+Agnr
tZvHFBFZtk9os8sRt3Z40RWcvwSZti0/QKxL5Urfmxi/2IMyWv0rroB00pDD9Iwo
cMfH4aJ5yaZ/IGsVjKpIgJEKIFaNsyZJe8sItL7KO1OytmH+H3O2GbhqwnI1Z7Zw
vj2ToNtU90eNrYrAZ3fL05ef6cJ33q7fgb/4Pe6hgsIs/Puto8Zle/4A23FBZn2E
fegulrGWsksVPk0CsQL8C3j1r6XXUNe06+AJ4bfHPMRY9KSg8HI3RbGZYC+roLd4
pXc2S6FWDYZIc5aRdBeG0HFV/CVqyBGUd0efURYI9Htz8XHWl7OqgwbbLarSnF2f
meGaAyVxnMuuM+PkuWZj4kQIv6AQRvwvtDn0cRNxJPI/BdS8d1+H1w48sSif5hgz
QGexra//SkKKwYzHOA5kGi3x9eqwxZEabMRtkyM9ZfJye93zu4DtQ8aYfslf40K0
CkHJEDWYVgUmBqTKhuf9QKwb+9Jf28qr+FqOc84ZmL/YxGgBjkMUEZ10gTzAcLdO
Un/wYKD+Y0wPbYr6uSeTwNUnhY+Vt0pC8z8bI42bGJUUfYp/PPYhDQ+9sls4REAm
y1JWtaunHLXTcQrCvTlovL7fdSmN4ZdTOo46Cp1HO6M6Bj78gB+lkztnw/Tm9XhL
wda/LciYrMi6uOtm1bT/vZGAv7b01KBr6aR/uKYHacsgAK/NatSWhiBAJ3CFFrst
gB50fETL91+JrwupJ1hzV5zB9LxZllvtFKYURyRi9PNlmeaNSt3gsvFi/CBiAjIu
4bFsjCGWSdDjEH3pPJ5IwPKDTWfAPPDiwMAbYeiljc7J1/iZA38StLUcnry6IJXe
EEAxufRG3l9w+VVIJm+66E/CdQBcyZqKfOB/HuVQ8LrojWwaZHd+mKcPiy9M6zcg
adHc84WmhYdqD6F89nMCRMgGNtRCXPRfOeG4oMVRX/qMtRAWFfPzvHtds+mXroU2
bJGW7N+rWiroTrf+u7YkHyenpjZuRYGXMcTCMXuGi/gROF2mvQs8yXpjWg3Gyvg4
zg5J7imYx8ZdlEfQNv+VqALhEmANOX9lvJAUez70X4HAFl4ziZPv5Dw19Z5syxlu
dibtbw4nq1n5dZL9JCaQyFwPTZVjimukjQCls74wSbKuDMTv96H/ZuDrlDRED5hY
Qc9Y4SZvZsM3/A4DDdqVh9HVrVgCXDaZlDi5JXDjYqhM6j0fSTTDlRWitGRe6062
JXUTh6X2bUENMbh6oCfVNjE8deM1THI3Wfx6XZFPd3fr139p/+QHdNL6qs/CDFsF
fNoBSbDWnNoNZvb08dLkFAoj+MjM9tfiD9aOEE7jzuhUg+bHGB1bXze3UMYkzvoL
+ehY+47H2bzwxIIg2BrkUgiw9evB08PehH18oHWY2in8115YIG81dCkNF3ejA/AX
o9tSqNfEM59ix08ah/UTOg2R4xCOIYfwXm5CPEJkeZYV9NsqH5HT7UpMbAz/j+28
GnVveSTzggJdjcYlCQg9JuHPHPUI6cJuveNeqI1n+0Mys4gpO60LJL5vDBoAPVzX
8EF6n0AkWdwiDVJ1+qJv2qdUnENt41Ir5f6SlpZhpfLl1NhlAwxNsJx9o4NFptsA
5CZJ4smWxWdQZRn0LZXlXWzTxoZtGvWSQFP82Sn8bOXog9AooIvduXBsHV6YXpmF
kWVRK1yu/l38VkxOrATjkBG830a4YS4HlmT6DRxEoBMyJjwcDrDDDta0VMna3FyH
GqISMvDdjv6UJNXVsaqRElvQ2jVztTWiDg/nmcWWkc/dqL80uAjmNbGtTx8wBf8W
+5mjUuZRcDGFRAr3L87xBxxcrK+L4tp30R5s9anKZJ5PwPWiqI37MIfR1vQJE7p3
ahky0RRe9asrXad7di9c10bPBUZdTqfS9gyX+Lfu/9Wk+vByAGOBXSdY+99zXDe0
OR1h7QLNfjloGW6+Yu5ZTpeeb+qVDxep4CZxu35d21atSM/CV8zcYcLaIB2g2q3d
oBV1v5nk7xZFo+uGUSdC/uYtYUGX6leeUKBX45haaPSFyb6eRJDefPu1AOVvkoe4
K6+mT9Rhqq15ZyZ0mcek4VVKNZ0ZZYUccd8d4tyBlaYsmGvt51kWutEwRkauqE6y
JRt+HVW1qkU9hXW5t4zzG+ofU6wx4HFJ0V4+pFxyXyiueO98yPlisfKXojHoNU0C
3Vtlla/Gvzb797Qmc3NC68w785IfqS6e2YL7FRxeKKgRtGRMPITb5GoAydX57Q9f
NviiIOp9jJIO/rrWUp7ykkktVfGAPkKxoSkPL/yDHj/PVvVmwZLxDzsP+iRCf3dp
dGwdkj0Rk5B2UMm6J0yAge3WtMHazHT4JrL/cyrfcZPPY7o1JlxF8SF1ww/DdKGm
q+BPV2wylOaMyvCEQnuip/UkP6fae+mzQ9QIUU4O/B10IwVKBFo5qsIg/3ELfmFm
7dPuISU4K9y/SCynXBwfIeENozC4tFbww3gHyh5gdK76z6bJnVSSx22HwLfw571x
WCEl/HdXB2gxijKuCWcmwV5GfdmOVmu3JqKiHxOsQDxOR755M9VkCZyjDXJaS3LF
ciPUU3zt7yQBVyB3tMACb08Nrm2XySrSaBZ6yo6Znqwob4LMrxbZFgZajBGuVmK2
VDVVi75VWdYmajiS9+s5Ajh0ugxxLv/FSEqecbz52fvj90omU//VeCxwk3QSBlf8
//34u/NmFFEOvyezwxIG7RA2b2YVfB2AA6HGhEalMg9aocfSaXkE1UYlwtw950rB
OF0nAwJaOpAmnZBGtFqqZnjVPup70vsGYqOoKg2nHFNgnTz64qHdYZhHP56COv4q
KCmbzhArVNECDCIWV6fRWhQ54YDIbz0ZAU4c76z8qn4z4FZfvALhC/A+kkmb1H0b
//l+VIQ8L+IPQ+UJtwY0wHqt691IEtgQziOZeRZklpugAOVjE1nZZq8zqVBJW+RL
AsB2yYTVHfmkGTqS/8JOeQ+qAHLsZtSMRI3//mjH/E4Ngulo3VU2ZYUFoZGCoKt1
ZL0/CsAXzCG7Gc2f90aeQKzP5BzmTd4nNo9Uke2R639WCsS+hl8K8M7zanNnRt8i
56HvbmU++gR27Dv65EzNK6f0yGFI+0dTeUOn2FqnUrgMDZUOa5L3G3yfa7XP1j8S
ofzr2Obvft4efa15PyU86oIBJroPWpI9ikTPh2g1ErWQ46I0e0xUw8uvfPmjPeaN
BcaokN6FbzLscd+SYMMhIICeXMlyP1kz+a9f7o+GoKhiHiUNpPvb6nUvLUntAMtg
+cBXaAnLejhfC/mqbTSQAPQVExW+Y6lgUlCRCPGsk3F40ndUM8M5Qsx02M3KU/PS
SVwc7Pl3n56qHJKM/t7FDYYKfOhsyxOLA3jy23FGt/nPcwGKN2E++6AHnJcU7t0w
8RUvWuRt+leTf2wxnwI8bMq1tBZbrw6e/jiL4JXRZn34s58Zg51zjucz2QohSJV5
E0W67WHUuetm9upL6LDp1h3rEsOntZw1jgPcLnFDzdo/68GtuW8maAZVa/NHsD21
2a2CxjxrX1xp2wF5of8VT60gKNyBMo4pJU1ELTU+wuT1BeTaMaON5JlugsglOx30
MllE9NPmp1rAt2yt/m/+4KoURsislNtlx6ZQGgY2v1iz84BeOo5xOWBf6aoq/tVc
Cuji+fUY15eK/WiMTsBm1QzreRLPTqLEN3W3sn6ROsqk+9xGStwjX0UfwhssDAcH
weZrYXVdF0zzsxmx7A9tDVQho/T8NfQjkKdabcuTQOGuoXUed/tQmTOiR9yLSQDb
lTZva3q2sK3FEYK8c2c+TLJAxdTH33A9nh2IyxFVOhehAOHSDbt+JDWE6hUTFFdL
z5libqdKNN9T6IwMhmT3ZX21qPRCAW6OAQhOwFcaTLDiMrsyFfpZxYHwGQkK07tr
VcTONVe7mtVl2YZPw10sEIA56E5lfognzkmnJ6tdDBYYFxJcbSr+oLXWseZlgRp5
T/DjqjOB4jD0Sa2UKtxAnfV+cSAqW2oSL9jHxLK92Ooy5XQl/6bMQ2kAuIugNHoY
vWeut28vKGRDSv48/B7ANxTbO84HqpR2qaBAe74AMP0T1F57on1KIuFrsCldCOzF
GIAjIVFH5Tx13bl9wVdIkqQvDN1xottxBwkHQnIS4gF2+hu6gNTNxCHGh/5pBicR
3MiLqmpKegrY53T71pYvwezxrlhv6DWoi+om5Mkll+qCIOJ5G0vjOKQZ7DdBFiqw
dcm8JCmxofiJmLTHc0p51Ds2qRYMOfi6NdcmeDsucfGFQCigMEFvSmy1oFLTXdP6
OBd3qvxm6/aYGmgrMzEzkQJqR8fqOzvDnOIBDz8+leQ90y5CfMiavhpBh49yiFpR
6OVXmX1p/4D6tErzXZAwJJpXXxeMSK8k1VB5nCGhYdeaAj1rNDA/EV5LO0UXFaHK
pYfhrs02sbvarAA4XY+hJS0vqcwU8w3pSdLBP/0ETFh40OQ+Rc2h9TmguiSf26UM
3NAXAfXJN0y3OyO01yZWKbGsE/3o7D/VgXoGIHYuVL+g7jpAPoia02iKb1tbxhG0
Pur2GmpUGZ2CjZRgBQPZY4gKVav6qwJYVSs3Xk4E042VwLYgmzJ2cbzX2uNoXWDI
uF/cQ5Jbr4Ed8Hb285ULAZ2u0XHenWqcXJYeDSZhvYqk83I4nivznZL1xJr4saD2
+p5t6Hq19igxfXIEyiAXC+MWOnO5gvtTCWTqn7WsSCs2dMPVROV4GOUT/nZv7l/I
88QFb7Kzim8aLxGvHwra01WUz6LXrcxYez/k39BaP27BR9bo/IaUrrX0Pnm4Vnwc
ohnAEyClJS8YYuRIxjRxICsnqko+UKQVjyjH34YH51J1OU5yQt90eUxay1GktAzo
tlOgXbOxut+cWEvAsknP6bPD0UVxaaubwZGuC1ZCueye71J5cfHiOylDC/faPJMu
Fwuu+Yc8RoXEeISKAxQb4Va75veHGKkMtgDGNTJVl9nXEt4I4xGyK3mY/SgLmdFA
J2CkYq3/PtCLRR9GuTgoJ7Q/oNCaFnJfOgAfB+j65fuopgaHmG1EQPbcVp9R/vWg
43/PYQJdocjdRnC4tqvWgVFUiA17WzNnoJCUFj73FilBa94h10A01P+mpL3WRunu
8J6QO5y1hr9oRvmr2y74wLaBOagmQAipA7i94xWmAZtBgeX2tHPMTjM/dlIMM1pq
TnYivD+8kJKDLWXmjhi5JDriNL4fgNF+PmPLFnNyWM3rK7AxG/GM9NZ6ecITXbQD
3cH72hhSm9zgo/F0yNmeHp3RXvVspEgJWplnAaWptdnSrRLkXxsYUupY5pgX0b+A
GKM2vRiYam9kIgpgXOrqX2a4jgdzuP0CtMmfJttn1dF0yp4il/fDgjd39bEVRPW2
fpus8yAyOD9UTzG4DY/x94vSjMXvf07E+2dy89rI9WixrPdH3KcBqEyt3W2zLjL/
1CSFBGXAsCY+N6O95OPK/t0gPwSnJlqQr3tIbk+V/kcAugT7hXSdzHqcWLuHJidm
ISe0XgaWcjdQSpoOaUzUQ/hw+rWUKHXRhIG/hKdrBQfxVEySbidfYkR0Gu/DlAeE
Vmsb7iG6DjQm+d+I67ojWABn0qxIGVhM8F65gB0TzBGh2fIFG1si8jP4/LQfVEpl
whLVzLryyn0Y9UBGYW7NnYZ73mHho8lL0i63ZaTyTRWfxluYrGPxDWa8FMFj0r91
3y0ydkihJeN4d74Uck0xLq5/zuyEIJ6Cct/bSUhDJM4dL3QQcUZi0Gd3fjc2LEqS
F3ccEqYo/XvxayhrfTi1ovzMyOs/lnHZ8IONjMojPhvNvio7yoJewBkrMDZxVB/M
GRFJxiT/O89XIxzHgNnHNsp9fbbcfiAg0mSvqmEGt/Wcx1O1Eu0SHOIVdi1v6SaZ
CUvELFrn98oEzFGfQODA5RHcptGCW0gHvScVR+AQqI3vTcuJMa/Mdg9R+nz9RmyK
45edxRNDk/KT+vk/FnkFVMBdB2Yj9OqayGajS3whrpgTNkupT648vBJzUaQdPOxk
O90rZTLMkm6i78sYPOKldPf4TCI399KElJuUigXSz5XBgQNzQ3B62aR3bZhmkD9w
LOXil/DKNJj0M9Gvmvs03OAsTvdXT0eJWb0ET8b0IAZKXYD7uba/KnVrP6rLnrNI
nfv5YRtTEzLS2vDkYTaOiH0rj85tgqfRkR8j2jL4JfQvT+Vvj9iyNwUoPV6wxZol
+lJT4MrSZVKyAVReZVS2XAHIvrVx3n+guFzeZAWz8m+PNv/kh0xupaieYmhEFEB7
ObXinnqY5ssO8+SadszhF+Cy+ZFFkGXimIYfP40bjI1clfcUQbT0Q9rvzcH5VOpw
W723aISuqmNJVGJpZndI0PkpJVIviCHhDJA2uCtMlXX9xVzvfr9xdjzV2bP0bWjK
5ecn2PZ8zdvIvnx5FqE+LzAA6nUBQoOaN8QWELpRxiNPcrRTud3TFWWZ/QkJfA6Z
+SukvVnjgNJruUAdrByTnKqBehC22vOwKwSS1ibjVzv8MKL1UX1My/5L0LIyR2Ds
2GdqHURhEoRKQ6iFw2GwIUSw75ie+HCmPvKKIip63QlDmDgYsnKPjYETVjybauGs
ttJvu7jkuvkuoZqJ6jKnyQBg21r/Xe5a5ts9jnpS5QAxOZzhSVpxjWHabg4GE4c3
Xz9vrbxvsv0gnIoIsG12Irgx7rUjg+vj9VTfX8IziBThJwhjCy49LQXYOfP/XgiD
QYzp7UQlVNfyWr+Fhw4UFEFY0uOnSP5mgBoiH3EggDzASSAdqVgACBSdvRfypQid
MLJCR4/ny6SA/31VTEh54UZTbDnqR8tiU16ocsx8rsDIOfZKMHxsMlrLyXhhu7m/
dKTZxXAoEy943jgSLAf7CXDqespkvjli4zgf+wXosfPpP4RA/7bFxaBdmHkm2/Od
M5FADsADex0vH18Ww5RVKwNVKpC6C7VqCDP1BgJGt1ZMPTlaMqf6j10QD2RLTzmk
oCwhPYFZdlPutEHY8d9TnrbAW0/SvuOKEkvfJ+y9rgWZLSM6DO7xpUsdwdCdVsyI
3d1G43s5/A3WD/5tt5rx2nKpGyYRYDfIHRGKQcfCjklXZH0uSCaPMy+LrmF1GZNU
8YcCKFFaxm89t2rumyW/cDG9baut4Kaymqw7ALBZBcUiQrn5DUqxav1JnrwLJwJv
ywT9BRtsS9MgsCKENA/EIDQkx/PEbX4sn+VXyfmHzwqAGe8TPKbqhn9HafzIfC3V
t4lPlaHzL+QMYJBBt8gesaa1NznzTRRFRofjjiFsedWYnqgMdeEv0XCFYGYfPgdc
hmXfhgKvJ8U5wBZ85rpv3QhYvgOudvbAZwzx8plGpSh1GyqfzYklEh182Y0MoNCw
cn1vE+LU2y1d0wzuZl/y1Xq2nZS848HpVvfbC2yjWk3SFSOe0PyaR54zbk6SYBHK
Aj8Mk9IUcdLlVbDNcEErcrDbZ09XiTdO3GnIp+AxkfPrzpSEad8fFGxBvoBlfAMS
NEk7B+8pRXriWxKBx3LXLc8/tNB0s524ZP/EMim51KJc925LWqLU/LGu//MQCeF9
7i7gZtyrssKS275Im6IR1COgz3755yTLf+Z8ksbrNjoqJ6eHNhrjRhSqbH44KLP0
DJ4h8yGxyvaBle21LDjpWZh1GFcyoMG6PrHuC4uoYB4PqNQMkyywVP7EC646qMVc
xX/GgacWYjaSKMOYji+dMgUdFiIAYWPzt3oaDed90GYW7z6XHTabihjv79dfboqH
wZFJhfoIyDRoEC1EW8AbGdxZoEAHuWeuxxZoHgWnEHhqFxhlugmRYIA8Q7DjuaW8
9clJ8lga7jtfh9+zqfkdkutGxjRUY6FdiGCd8MwHuaYz53R6hT4MfzfGrIst8leR
AGJDFSkIg4xg+Xce7gkEbLNRlJ0+rO/gHMTv7ad9PLZsSX1+uAuLzgJsG4GJlour
JKqqu7qejIWqwXdL/eDah6pfta5obZiAqfw1CePnerY8hkoJhz5+srUaS4FeFcO1
lD7zcKck3DkLaoRcyQ9CCZ9tNwG7BLggbTpFzZ/p0EmLSBkiIUl4yqJcB/sjuMw4
ceKBHI5sTWafgLCnAvSEzbBpMtduVx6CWsFuDwu1QE6ZryUGE49GAaKPpiR7/7hU
8zPAMApROv0SVwMRqxGUyWh2rpIx9fYYtCutz3HhJ/OYESuFWcTMXiqqvY3g1Pt1
zi8pgB4MZUj8VX7nwtj6io8sCfXxHGEAEqFf+Y7wgqaGngk3zEbQdLV9xNGLFPeC
XDM16Ch45UexhxWso/WTuwRTqh3Pis0tTZw/wlkEJn90f5AYq0WteqmrcQutqykg
G+LrbIV9r4cD27rRTOhmGODYfDHcbE209jv00vE5yBoivIkJXXJxnlYpjthUxoSv
cGysplesiUmBoxqKb4JNUCB+UvkpAd7uaZvEsmQoRT6vVHnexbdCqtAFfeVNdcZ0
odubFLGScls5Pzot8sDDmvBHi7zPBReVyXU1gVTvVXmGf6Wzz9mL8gXFdbHSCIoR
VD155YMKAITFBl9mmSjPdJmYTdUBBhiRG3B1zVyfgagWmulqGMKyppazO6PtUh8m
EXHkuzBkGwzbxR06kMk9drYYmjAKS4EYn1j5hBqux35DilwqiLAJmON80Yymjqdc
W7KbWJr1dXUAJD+g3KWAVpY2PA1RhVh+JnzaJWnpJd1CLrUoDV/nyoDus51soyTn
tKtogS1+eowx0q9a2qXhTZiSleapygTIoRJrJYHdlIHGQ1nHxvx/FjTUqL/dJZrw
/+ezdy2QqFoSlfNDfuEO20KK/D+ZP/IHCnfKhphUIHaGrQ0O7oGQm58EikPuhAAS
ZQmaYiF0RtdHoUZFtvk1PXGSd9wsXN7KxBbqxjL/xVgNaOuZK0wJABmllLSJJSH0
+QAtBOPla49IruR4trKbeQ3rWoyhcpFthfT+WynDFFv+Z3+jZeyODaJadsXE9LwV
OZNj+rzTulB585924nFdtsHmB8DJiZ4ytBH1JSQDVekWFvkojxKdwXvymoE8xUQY
CyNpCCi1AOnuBPaGBf9GsvE8D6cENsKNhdP8KNcdqgJe3t31BvUbuqI86Dh9yV88
EyEU5f0afa0ePxTY7ErQbVlkix2Fh8Os23ulFIhaBEVGascl1FxKjEs1zCsdRC+5
ZYnJVkYSG6RtJ0XLChEFRVrKdVPWnI8T37Xrc5H85YTeb+l1KRunZQTxsyPK5xhr
oG7mUiFSiJvmxe/ybcsWItL2xQ6lJrWDSWC5X8vt2iCEKiDnLiXPR6+2VtF0wSVt
7MgRn7WYrKwrhgRuogE4whm9fVhtXMJgMTmKik492RimOWlELusAcEI/6pcpB1zc
qtioK2LNpxpcLrmiYBjrnbLiGh5vp6geSlk0eZq7a0CgCbaCrtsizal7hZ3+7Y0i
koxQilTFVLzM1ZMh1EmlfwfWNRvaTeNgSvQaBxIZamPiNE8nrOrD5671TtLPmktx
nTzhNagRKxg4MXkniqJmVwZwq6wyUL6DPqLS4b7ALyXfzQb8WRVtcoSD8Pmrf042
n1gAz4Mk7xtT+py8E6O3roN6wbfumsY5u/bwChaesTNYdbzFSA22LeMlyQsLr2ay
JYN05CxxjLmqA+9daWmZIuUv+sXRPZdPtHZBlKZDlZbENVEg+tFjB/NRjZBdx7sy
PbfT3gGGJF2UUZxzBc4KXKa0g8023TCpi01eqrbMmGGuA1aw4jgEfbyqQwHZ/58s
dLA10AGt0k8dZJY4bFbUfuiDMLsX5CCBMwFj560j8LkPPTHBpWAzVAtQ1p+I2ekN
mD9QkSOQrdBMMqsIFSwBoHOkiDZHzhWtDa7MOkVBvDJKKAmoN6FuM5NqMW/8dse3
xSZk5P9CqL0SNT9mu8ioXeL/kOA3iDGCLAhtm4EbEhvrQMlMvvOc7XswyA6ZlnCr
6s5ZOvJUd5F+tAMYUw2cJPrdrgt/CQutYHZ3lc2qo2CLkaInRp45OtaHzgZENH7j
ktF8gE4gfh6Vic2EpsmdCmNIaAPJC5NLIVvdp/RmFE+WPsbZ2FHmP/xMipSMlvK7
txTP5Xk7LRHKFlUM398oiV7N2a08Au2xrCzhtJOrDkWj/7KcnW5fQF9lTdQRoC4Y
PV9Gp5PXOBwOsLjgKaC5lhYN3NdE2yE6jiXEOQUg2nle1gOS8A+bfZ8LqAcsG+Jm
G7ytc3ZOPp4IuwNUvV+OjhHo7mpo9K/fyubBI3NdAz5JJiVRT3Bs0Iqp2oGDiiz+
UCP1dOQvtTG5uASCQVKe9hwltypPd3jIwP2QRvJ9I+Zljy4WFNgf60WkzSsHi+R3
HCHIemw1B0AkfripMw68bm8Tm0wPyrV2P243j5BtJasA0hrb3e7ihgS4IDuHWgTV
91qNsL7SfPLHHAkGVCkuZcdcbI40QBQmXrA9nTs3TO4FcisjBKiNfjTLM/MUPGX/
dOj56Z8Xqjlvlko3c8pOpt52c9AMr1U5WlJXCDvwvwcjWF74iskNVOjW1Iz4Y1Hz
C6FgSm3kVIkF0FOC+CEFYfyFGO5bmpd6y+nftnu0Qf4q6ymDTQaEW6FuZa26UOT7
73vQhGYJ/Xl/P+ddUnJQDWlFydes2yNZoNOAfIggBKvMELqA2rV63/o8vBDzD/1I
Bc+FMKKfz1/H8U/wmcb4iPkWPFeklgRjYnxmhHzBlv9pLgdeS++FXj1Zc9OrSyiu
uVLTLRWETW9mwpe0cuwL+xQFnoJ0yutHz9rfvYuD+0XBIorNswHHhR8ND0Ltr/Ol
MUmWhiCPCb3lMHZWrtBl94LlkNIVWNflebbdbe4ZbsmV+9rdjRorggcu4bV9nxLQ
44JsrNrFupmXj/hCyOVo3GV/g3x2ms+r5r4sbEqCBCOLFPUUWiw7O3HpQfG7HQfx
SEF4cIxfneTB//qX5j1InwORZB6tuRZEGAYfrUn6g3v0QCKOie1l+3W4hH0cd5J2
XNLsIZdUMXalQRQVDMOqORgzeW+6hI+/igJ4bdMeTD+PW/QtyISG7qZFnPVe6eVb
9FotWKVJivm9pYUYFzujVN+lqGwXzb+I4lIszGZv6ADdF9a85GB9ba9x7w0Cx1p0
US8xIUsnTtbIIdaM6gJFuSwaO8ndhs7t7FPNCV63fj8SX/qHvKukKrG7uWFma1T4
oYFWfQre22hb24fYjCpwN6o1FMUpstrpS/Qm5RDdT2NZlHa4Ss/UyZdbJGWFY4NJ
1Fo7319u7F7TudS6begXBOMqUG4X1F4ibh0jhRaOcNXkqUDJCJZ8LSO7fLhBAFEh
FoyIRFpGxjUbip8GQWjPm9bVVq+XTUpF+wjZcQGN9iowHzIPcaF7U4KoYWCNP+v1
Qpdql2/Md9OmcKdiWx7N+G93nmnqz52Tr3uqutM/ndL3Ui1B97JwmPIn+3v1fGYv
R/h3ZUIACHMkAsaUb69BxiU7hoqFI8ZZyol8/h4/J5WvlX96mo+MpVNEwu0S+h94
Jnfag8Gdo15BPFqAxb4zpZ3aL3xTa8tES1gRD6if1IGJ5ehmZFkp5WETWSSrrPpC
rpiUjZPXU95+sW84eqUApPbGrxDaCFLJ90zgmyoAiNXW9mCQCKC50o/K2e6cMERV
yoBKOe6MZ3osFAyHQx16TyPjaGlE7y+pfEFLmjlk5vZYGEDWUT1AGKcpFhZDS+x+
yPP5sCy/B73QZbYVZ2+3rpwFDaJ7fs1TvL45Lh3pyhVjHR4CqEYXoy5Vc3GqaikO
UKQyJjbrGRlGKhGkqcnXBQCPO1gLUtq/JWunDoMToAfwtuT+uzA02W4X2i4TFa/P
cPf7HgS/NR6cvDKKY0ZkpE5tSEjuPCODPTfz7z0lzGNcRMC3Ly14gE/k8k90An0o
F9N5RpCURXlFh1Rm8P+75kKt8cZMRPwt+Bq4+2W+/Rrwz9/xi6cB4Z9s9dBZGgj/
5FdoX1+qaY/cpDVKM7eqc216GDKiZlp8umbCQL+/acRjDjQy5AJzS6u7WOf9R5GI
4TxpsgM/gPJpZIE/UNvRic+JaJBJXDjlCedYoPIvp7REICeu+3Qv/UcXjQky/slZ
xmEkbJBPNgEFJaw5Fyu181kva9dt/LAR7/f4LX/pX6diF5GhCXfjeQPke7YboBXo
l79AFt8eL+FWM0WRdZO/HFKaoCdSkt8JsRID3pyKTmOVFohB5CWTrTAjc/W43qIW
LFGCs7Iaf9WNibuHlTF7Yo5MRzdp8xTJDdV10DU8hLkyXqO8u8MZROKbEU8epn8R
ofRwpqLHGoYDWBDNvYdyYSIILtEylGsKiDlMrCf3niwOsw2JeNzLsv78ePki5+pE
sysy05ACBL9HtfDvjc9L7M6gGchsY7fPnvvltZT3NNX3tCOC7mmV1hji4LoxYIhA
xa7Ue9kPj+c/EHCi65nSoxnXl2Na/JqYPYkWN7LJYXreOOVw/E2pmIu9sUFs1kgd
Na97VN0QJ0qD4j2JncfnB3G9oGNwlLBgqMSxL0Bcn2ETXBMY1Sw5/YvvG0yy2vOX
+qXD/6lpCqSCropO5dBKFUGomos+U5DeSbWfIBZxhW42dntWgoWYa1PjppmaV9gC
2mBoh3DKWpDYn1LJMYTx2N5GwHbP0PvyFJHEx6k58SpqkQ/9yq/iJDx1RsEG/AoV
9shc0LdiJsOC/87YlsWzryqOJm4oPPMsnd8awmKj6XbfM8IDIXHuGIvUyCXfC1eF
VBziN9LT8V8rcX5S2CEqh59DTJ30b8rcHSooe7EYsPWqVY9hUOiY0zgdyHyRZkjD
31zeLaJrhnGShFElaR+24BNp6br5fuiXZUP5vg202aMp/uoW1mCAU3DdDpKGQXV5
tmlpkfl//lauI11HSX8T4WidjAitiSgnA4qYJdX605p7r5SFObE8rBHa93O6b62i
T8D5WLaUNoQn4qbpljY42tpqUxkGqpjwtNZymISGC/utEMRj9IUV7341BDcC5gwU
YDobnxWeusV1t7qORNLsqBPuurqIq3f1jTy2kyJjGGmsDkNZOFjTSMz3GZvqdFGF
0Go06jI+e2PL+p9qt6sR7XCGRCohGY2vDAsdKW/19P57YgyKxywY6Mq08a3lcNLY
vng/tV1tzW/ejA+FdWFBFUTdj0bb18GhE62eg6K6LLc/NJrcocnQg0mGncE0nBew
H55MC855Lnvo5K03EmHr8WVDq+dFDckQGdFQnPBnL7m+kW+/qLkGIQZOj6scRYqU
/ywDeRdPyCn5WbuoridPu6cnjibAvkcUX/ny9ZVumdFGOsUkZiGRLAou5EZOyT0M
4sr3juZ0Elp8/opSRAmioyK12u4uAyBP0aMvXI/IngqmBS/6pD34uT+K7TD+XAaU
RBhZKdMPDhrZD4bOX8pgV6TfRkaBd8frVhWPNhsyYvTuZG4T3+nUIGQEbIRQ5B+e
J9W1kgfWrxx8PshpkjfqNPtvZhRiBy1MLAkHM96YSTmoCkMHkGBOlZE4IVyq3MB3
bnQnsLz9Q9Rnuiv8PRfjG17v9yqVc2/4BfFEUlRqtZ5xJxwez8UFD+bZA6Pd/f1B
lpQJgCUwyFRnaQAlewSGrNSbY7XgjDHpEgC2D3rNACUloa6un7dbNrWgozl0aVeL
pd81Ho6/3YMiFpx6TpyyYEncIpvIuRtnuJ2QPS5StZWrVJTXMIS+aBkf3YQgEjGL
iRiIZVZVVI/4NoDq4Gb8upIJZPwC98VGLAinvTdQMhRDybxJiTGQGzzlmZ57brNT
eUdKMIAINQyBeEuA8Xs8DkUta9SG27ajd+jnci6TOA7ev9ApcvUM5v5YzXqbM81s
tnU9SQMlSUAtn2UYjhzP8sqcqiDBF7ReDsAlViLzHFGtILZ3aQsiMkzexE7au0bN
Qlt4djgWrVAOauekpchetoDxzs7Y6V9d1bnTPHP2KYQz65fnDAulZtLW6+cG/IT+
7dBT7W/Gk2TB9GCKfJ1kJNhO446X0iJDp+x1fnhGRw+3L4FSiPq8EsYSkUQw9oJ1
t9YIJ4Xts70LZnZFxzgEnZhxS4NwslXT2LkWdY7/0tK3gX1VN4+pXDYWpJdJ1Opq
6MQBMtTy+aIE0wiEBZ0PzaxTDd9CExJXhAIyDE6rks4MNuhcylpVPPScLz196dK0
4Z4hRx8EPZ0yXtBVGXYY/5+s2ZhN7mDAHoySaDodLL8pElqfdezvovNaIQStnRYs
LEWYc0DgxNuCUv5d7O3W134PT9eU2+aABnBh5Ca5y1zKtnALDaQOczIuCm/csorZ
MkhuE9w/LWk18k/lRsmLVPnJt5Ua38IfikTrK30JrRFfsijwrG3w60SvJKufkfg0
+J/WXu0FAxUA0CyEI2sbKknXLyhyvfQWThCUzSQUPoTPxy3izGc2DYw+Rn68zt0I
znbKYWb3xmTA7Bzp8UN88OxI6Avx221yD32w5NllICKBJ54vlaGMbGOolocXL378
C4VUF0oKSIRzqLdzrCirKKXEeA4pAABaEJI/LPkRwr7lrR0J9MFVVfvWd/nLymuK
Qib2hliSjSvQG4QbxjDhmQUzjCspcopjeVvzqmSMiJ+duqEJ3Hz2STNTResGancx
rdzI7Gxup2vy8ERdb95psVqup8HFAHC9IEaOfEybR1uQm5xw+pJIKpJDyjZEInOa
TV+B+j70ROShyvpmYQMDbruL7I1hJCqWpMErgikKtpxVfB4lXEtEuu0smz1oLreL
qToJOXNtPB1BLI7OeZJfrxjlfGRvk5pOCicl5D41ar5xri5Ylw0SNA0a/Cri79ja
sVNYLbgKC6H3npZiOWCSjDIbLC+wsLh5ibranRczi/GxOIaW2GZ0t+nWPdlS8s+r
zydJiUuPhiRJ96j+EzobBc/K8/M+pZmwgbfURbNYUd4qazOut91LwMxuD7pDeDRq
p0BxqX1T1y2jw7ixiZn5sbAjSHtKUuEZ50qyQWB+EgqQVk8+0X2d8CNQO8EbEa8N
V1wDYapSd0J49FY3G7r6m1p3icfmDRpVMN1qM8Hae4ep+t/ZSCozBdy9C7XTYdHD
1Yv+Xh0oVKoY4nv32honKovz3zJMasbEHLerXfuHNYNRs0JvAalVu2GVA5K2RnKD
H51xJU6jP50j8aDjpS/jO2P1wFk2Mm3Mfq/nymdrLdMNubN4OQAwAyPH/TvoFbEN
DA5aNpGlD0YwOQsKGop9JLM7SjdRuW3/tmxq1g4fzo9g7E49waCV0YHQ2t8UJZuZ
FPY4aPG4j2bP/8I830Bmc8MYYPU+dgIrTZGwuOO583xbynhrgy3zCmKc3PTe3Rsu
jNNiGGRQIVN8XfvDn7WwzX30WyQgbA9eeyzLJz2cT9bpEwLaSHYZfHaKjDvignOa
bjsNBToP/jxoQY2akcaQ5W/uCc8hDbsF96+Hh0jU+owVtgKUQ3mRfUM+qxQ0HWep
i1OxJJiotywBCElYAmFMi7TVbCrvvjFkq5Ukz1cs2dLaGpvrbl6BOUtx3KKMmWk5
wwSpIqgW6RR9aADm1Gtys50uAHiW1AD1kJMxxx+7V8TZRJteNs5p6lSc25RbqBna
2ErMzY/8sa53POKS80IFB7zNCix//DxUasoS8Iajvs1b/eHI9uxBjT6RlfHDuhqU
LDInOC3Hedjua6Dh+adPmGPpnivWEXTw56LSkTLOPQjFoElo9Zi6rPh2bvFtN+tJ
wIaF2GKwoFnTYZdpt4CS4vTJ2XsFmpcmd9Hx5B7rU4f2ulN6K80C5v5b7LuWmMps
61uL05FRAvRs4HPM8F7TCxNa/rVBa+9CCNEnIsoXsSDCjww7cvRXF/IcavTZxM5q
f7ckvBfsbPzYVcIpYc9IHZN9SNX6pgjtjmdT/JedDGAswPM/9YH3cEN4RxUjs761
t7V8hR9ROmxf8/Jvav2TW9Cd+DH3LZww+/UjzLGKolOvE4pqwqCjmR42Gyc7sMn6
cRtqhD7k8z02L1RdZCFNUKaz7ue+oeiGoXTBsuo0uV22THMgjnJwyB+2QQEngkUu
rRwbO9Utc7cDkcsClOlq3C9jYgCIYsaQO9GDIL9xAddXHUcc8TekZnQNsUinq8x/
prusHJXzpLqFRchblaJysER3XaHuubOECDSBcogMehFf/hbcorjjpBJRlbqA591/
FCIh1AyMtOe+JYQs5m8Wcxi+BHKU0F5gTHPxSiHHZnVDxHfWciorSJNCHjh/mPW+
/15ycqVmslT3nMs0hm00SNrZ9/ZVmPBB4fapHJy3hlBoV7/tzL/1bMg/2Mi5m1aG
+O0ZToSOBGRKPGD0ChmRHQCbS26RVhkIAMIuviyVzJZPor44KCPiP9OS6TJrq/pD
TgBFA4hNbz2xr+c7aSBYakEuh3WLXRw8JpNNyVD3vYbXkO+em4/UwWay9cGk1khQ
oLheyuwvzod3NEfJwZBI0VDxdzIEJBuwuLE74EPhkLoq+S7M+ftMfzMeoGzHDp1/
4MggtuSHgBXt8pfDzlTGBmgJJlc5eYNXrcQL0V8yFAOS006N/D4PtUf5pWq7cHmq
DdnowX1YJQV0gIYNP+mEbPQJOqvMSg9OMq1fkAMQ7ZuDAHpgmk6MQKc+O27e2ij4
60nOXz3xHK1sM11/tIm4whpqEKYanWxXwvnUVXIgzLfwNu15lmgXrDjP9JprZ+Ei
Jy3SL9dH2aI2UR29XZMRSC/k1BhlYPi6IRVR+Ri08cSImT4kaHondKb1eq8edWnM
IFMGaFTBcRGNj9wZXUecTPY91MbPI7kbcZTOS10Hb7m10ymKiN5zVX6qWZn/rFuj
pmooZ5BxVll5B0UgoT/+o3EGgCu6BLwHQOZcKKG+Rp6efO7FFV4Ha7BkGSZJsPnu
mltZ2fFX+vKMjv4rK6DG5Ngvct2Zo+gBPl7sx1Nc8BOvHT+qK1E+nC60myer8nbe
2hclvrUPcIG+Ofm6lxpy6oKncaoEcwnnb7jIlK00iee/KoXo5fThTFxtLftNuZWR
yhNzQdjFPT1VLCH9pcVLs3J0BFVtukdmLbUGzp3VgjAwj9BciTSfiNHap4CYwgLW
d5bHC1TMkfvRB/XX1RUjbPChFpnKDgvmU3R+7+qgvK7cJHHDVKiOmJ79v+O/8XJz
oi+q91YGHN3VIOhpa5JArfHqfZmeDbKUXCP03sF1tTS4pgkOv9c4j5+fdusRlK+R
ZaoCsCVywrkF8vajpjuStt0Y+IbVXwRTw758/b4oqFHfzeo0ANfvsx+vmr6ZC6Pv
HW6DYYGSDLqCGf5MYGDiW0aGhSKV/jltaWZkjNMBA9hiN7npOejjEwHLValztH0g
ywvW5j1PxkmQauXwSHKVUhcFaEMl7fJOxDXJmWGIQj7AzX/07yilsPhIYVOZZNzq
qOgg1c03A89K42AMM9PPsPUWQ6WdsHL/eUwfLwbSOQGlj6dAreY5JE7liKJfM2My
uXoeanB5xAbSvOqukuOSGtpoYU28QR1Q/gVQN0LWrolNtHzvGWtbYmW3eJZnxFWs
lZmYZHPKhYCzigS/rQ9lu50IGah4GzSVNVnjhXlYrqpcPdue0GeYNfzMC22cgEh/
4KYp1TehDnpkcywdtxCzt6NgoBMOHjHHXJqqZbw211L2G6njloNPyrQr6x1ytDtf
nwCLTUyeLD3iiWZNlx0l2Fg2dusibuNV6hxw1LM14i0ctmlAtDm5be6fuPdL3YN3
VdzYz980TcdmZsvXQ099sYMEhzp+3YhCeEQqzT1fHLDXX8wTtIlRowfDcBEaJ76+
tBKiznTJjdnAhn3nwmDUr490YehOYNMTLnJP5FmLAKADNecBl/yJSr5ROxvcQ9a1
Wgd/MAkPBHXnOjL86ETZMOHQnESlT91v2baqW3vY+Ju7QNFaoc6kESOfbakn9927
FuhlbLv4RJQ73Dr1nlkRTXIv/y/9mMFyiJsYz+GAns6DSkZoklCeQKtI/lRp3K0d
MtHEiJ3skQejBRrTbHYlqET6KrP++woM3OqtPCTrz1d8IfVnHFJtkT8ZEIU1m1G5
mlfgJzj+RPeziCMToYGIxrKw/4drZq6koxToDzydULe0I8ulHYpoELO/82y72oVN
r8PNYfgG6NKEnx9pTjL6ADsGcCbXIUUy6lAyw+P3fkxSQiRCC8hn1Sc1fM/hmz/W
YBU+JlGimJK8ywYqKyG7EBGqQxrzzkJ7gk9Xt25P9aZLU7yoYvnEle+nQUvo+Rct
i7rYxkvxbtVo9YLgWbzL4Zq455YjZ66A35x/PolBh79lHPOfVmPz7suk/hQyoNs9
D4uoVt7NIuyWugpvnHORuAMg0RFFypBInxLCndvh2uqWYvnnMs5kG37zmM8Lumjy
Z0kSJyEgeLDxXqoczwJxIUB+kEDVbNoDgsWFkepVcvnu8hCykOia4i9vp98/nI4D
z7v7HcFGJcZPBJNpcgiFJx0iAFrD4fcTgDF/VZ7XDEHVN8e36urtxWoIM62PwF3w
9CAYtUdf6bxtVdjMm1gCn+4dpV4Lsd8iq+rZQKc2Man64oNC2ApCtHyrhS1PTVw7
TmnWSGjxlESqCaHlYQ3EETI8eLLBF6R+qelR4HUnqyUs2jyxPkgorwFmY/AarXqq
PXzp51D3fbQtmJDUuj/UldlhO9GK+PYg2YaI4EIL5vi6O0tdc4aM1lj41qFuk0MK
KPAVEQxonxJihYaKJD5FrAi07xgPNaRY6fzB3lxR40UVjx0MFYxQgDSzQcgpgko0
F1krlUb3QqGXvhMGTphwbhrl1VWp/62WpeICmhIKc6L2nafLge9OoZsUBWBxn8mV
DwZ8ZRgn8ERjx2OLhbmTBVAG1NGPpa4lwEBXhvTXUpkrryLwJBNm8srimIq+cC7i
U8Jb4OHXXDkMad7/vdp7+HXPqrUEbU7n0OsF/vxqwdoQF9pn9nDeG2EWtNmqT9tE
aGP7JQIubXNl8IQ82Nwdw4Xu9P08k3fqmQMfMuIbd6sOecHHdOZDMAdMYfyWtv4e
GEXzKlsqW89OQi8eWMmk0WkuIf+pO1DLQCIxxRDesJHPMnMPfiHvJElILGPI2MI2
wJsOkIDNziDHS/omy6jksGmv7/ye1JHo4D3fpMDesu115pfdNaX8PcagUGXkH8LR
MdfbRRdnVFrdrMnQSP9ENmDvozIdN4Sh3XO1LpU5Exbz4bX4E8yxe2ZFdJF674QY
xTOyUQTZQ+oSaFfmSKO/u6I3zCXRPdB9/SF8krPzReAFkYaisPWUDyIIFcmnT1n9
DXcG+CTpSQ030+jbVyOd9pM1Ql2f++aPoswrTgI76IQhNtIhpir+VER3tre+viIS
hq26/QbLCjQp/fX+QJxDLHJ362qk9HoxbE1e841SQhJ8vNvUZFSeFFfBmXo+sBuw
83GSsG8iB6G5X+MSD69rKkDoUnZbwFxybxKhNDS+nAwynDu9D1k0bX/iuXXAp7iJ
92sTWe1D3hSQfNQHZZhmQzeN83czN8k30DvUST/cY+36GqGLCIzr/Mwl+j6hNANl
CuMTO9kGTjTJHUQdmtnqYKAdgTHkaa/pTf2+KJKW0u92iqfefHg2wpKblAEX+vLx
RkA0TRqh8uqPzE3UONxtZ0Fn8OiQISm+6bp4MtT9tuGP3G9O/Z1+kfrsLXgc/4bL
9L04y+qgoueR8kBhL+XClGAYvgELeiHJDeMysHK8DwwQLoZElDtNH7SIDmnXNfiL
LST2uQoX0hqjibMOrN/faArlLr2kaAwdRn78rK+oKGPvCT954W3Olq7OKIhT8Ts6
MBsECavySNhqdR1UJf4qD4qhOeuohywF9dLSx6L8xV5siTTzK6hvJntEgCyfe0/9
7vb7JojPqTjxjGCLX7KD9dsq8SZ1Cxl+kz7qLvb9Q4sRidafdvB67/at8Ds2KHl5
P1cmRWZX/4qkKeluJSHkcn+Ns6OR6pdGqvVsC5OSxPu585H5bB4slmMLq5o1zjJU
a+iOLGGHLRZewoSbuPe/SgdGpdZDa/MJptDYMSxl1vw=
//pragma protect end_data_block
//pragma protect digest_block
uOWxWuAxDEGPCFbDRu3HfZp4Czo=
//pragma protect end_digest_block
//pragma protect end_protected
