// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oR9/ne50lR8WexBaWmV4UM/s3QurgcsyS51dOV3PtQa00jI3rYUzXcTrRgqh
aKceKvLRxsuN4JWbme/gC79CuW5snNSgUwQx9NmVOZzD9/UY48/fyGPM29G1
bkT6WtYz01l7WmSrwLdmGmnlmuoGcOkXuunuyDo/KkHi0f5TawfBNxBgKCIQ
zrnhYVEOqWfHBBQyCVXVPvOp4Jg9zWjAyMdfyGlG7+7eZYbro6knNji5suKI
CVooKdk283V6D24+/66GyQErfmSB/uZG/H74ZhV0Geh5rlIfQypEt6qvFSgN
Gggj8UNjstaz5JoDZphmxSh/lzZ0or9ZjHTO0QFKSg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iVK2sSNrPSzsBtrieSeKKW8xs8dUYqLpnfzPm5OU8OCCJdysbzQof0tUT+zq
dcziNchv681womftPDj4sa4hSaeMu0ckwSm8GJIAgKhTxzi/I053YPqGjM9K
kfAHnHHtCE8tEDo0Z6dczzVtj0xmK1gCYVQ9Oc+RQtz1OmfExRh1Ltz2fgMs
Jim37we0wGck1gHGY2yObXBtpJzdBDqma/lv+Af/IEbeOUjxaPBd4ZmtTnd3
oXEeqa50e5JlU6y3W1qBxL3Qv5bRB/NqjPgvnvIv0Mx9DQMhLi82mcSUHQXX
zekL8iqY9EnpAPxFUAesEYg+h3q/1rovPT/esMjCIA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WhzrhIi10mE9ZMSRQTEXy4QSbn2bqpOr30gkNTlduuT/HTMVJPVEiJzRHOrT
6Kvt4iXFD77oOUZivdEkHAyxuGiXAbPv1uAeahhz7fr9hTK5OVdnSYQYlfie
nxWKQd3kIPdVkEC2rGjIRA6X3V+RHj1ZOKwKOoPuUS1D6cTcZ+SCvsTfmRoY
vrQ+mAvSuhFrSrkK+vMwIxnDbqldJzp6/PePg/t4bHHgsV5ssCDm210nCHXK
SZPdL01KLvw5IZoR7lt+Fphwu2toxGmMiv953K1/32/tV0GfErJjbcsdo63z
XV2WtrRSypAwxODFY1vsZx4EGzJYe6/uhzrqwFcvxQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pV1iD1R18vO05PHyuYlInd9iqO3JsDfkfNa7Wjmt8OM3LzPK7nuCw79PNQ55
p9iSZdUvUAUfDeFpCfN48P7HjsZtppqQub+l8sVYUfNeIMiQhH98xUpR4i3M
LktgrJRDfXdHx+mmUMTZEFQQEVQZnggVeLnJYCnTUa180W3awXw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
p5pip7cF+LZu+l3EvZO5XEcsmRWUbQe215yfGDYk4KT2Gg1J8W2ITGVKvO8V
Uf+k429eS8DkMl+bySt8O6gdAWfJZSGndj/CtR69g5pW2BpSbfOh9cgFhuxl
kk0O7LokBVG+agD3QIdUDTpeqZldWkeR8XmqC7ouU471fqYMIuo1uOi+PnvA
Drzh5Qovs2qJ8uaKp2htSl7I8ea5mGKFmS37WRmqspAUuN3aiaTeE1xVTi7I
Jghx5MFKQmPMHeQ1QrT+kqsgtWbwFOQ8x1KFAhEnxgSOcxFYTO9Sw5SqXIlS
iwnGAdOVOGqsQSO8DVGWgwVe+33DXMyRumYz5bu/z9Zh3sw0CCBtymqQOH9G
rmM44CeZ6wn7jyUq75WSkjen36y4OeaTDdVNFQ86kksQ2sXeC6DhqM6tvZwV
v3NwS5KRCdkgtUzpS4FYoPt1i4dIUg4xss0F3lYkHEthrJMPXXZa/5UOj0WG
Br6YCh14dsygI6Bhe/jbHPo3/BWkZlg9


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cUrpRpXFQ4SQxPgY2rpNQwHNxOaM/f3BDCrsUXRNOGlxZcOgiK0N0PWVJCDw
HRIXa3b5oj8K0hK/K7IWeH+/JAmT62C5pw6p2+yKiVTZiBSMv2fSwtVENt/W
NlnJbu3tOyoCv+ZlXvHdCXPRmMh9NozQ28unYoBNY7sMlubTCB8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZGarBz7AQOfXVYmRrQP+clsC4KhM0sZ3DhVTx60DLVdhjppLHntbAz1xqLK0
6xzAODXkyL4iMKlpt28ltdp2IGpHEjio5iGQO3UujeUwB7oLtEsDeT9jdCGP
Msj2DeDP0kFj0tkdRLI6Lwj7yrp6dWfZ5E8wL5gwN7oLPHSYQn4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
nFbv0Lb0QI8dF72dpl03/OzjKzLJzsShuNsPbpkTOsh1HeHIxYNO8LJkAOaK
ckOIwUW07XItBde4H/OzfRQ+swh6X2yOgVXCzhKPHLBfBKTuETPUsCn4tG3+
f7sVR3xzXwOCl0RkX7FwkpMSJRiFi/Pj2fbJvpQV4Jsv/Z09qkAxyur5jSQO
a1wFAPEs61lllUTZivwQHCiELGTrRXkJnBTWqUZ3ACcBEXHOtOYmtaLDybe6
I17Fn6qr/lNevanMAnPeetJG0QrrlYBz/HNOIys6CenZ2+sfHhYg5TyATJDq
uc1BkrHrUXHzIEmjBlfyAzE+sGg+R0J8xc3e9ILLoRk6gm9fFBhR3ywkmJX0
OPILxeJGVFtwv9F4ioQRJZFtj/cDIeu6/ltV2VVvQAYEJHNLZKNlU1IpXX2T
rkziOoyqiz+2nnGwFcojgU06MKDYZLt5h2hAoEyEpmaJ/CKtY0bCdqu8VpQT
R62bhBm+plqcmvcOoordu3h9AWYuoXTpllR2ZgnwwS8JCNKUupBt8tJMJY9a
CP9fi669act34YaHya4sYUul/FvBO/JeH86yu1QEmjLwXduR/5uR6uhPUyBE
kBQ5XxOUanKL6/82zXxIjWT3x74Pi2ROynhutroy7v91rCulRvpPrhDjnRKS
eFPQAU/d7dFm7A6/bEcvMG65dhn+z3WzKrRXwNPSwgGMOCmbhiZt1hWnEaXu
fXGKcmKwlrTW1QjoctPwLYaLeLMjgTNO8JvSIK1n04dzYFqRdbOjejsQGwxp
k28f42SfLw78FTuWDX5XNn7i3dEpLx3SQ0myDJK2wkw/f+6efIUB4aST9G/k
0GaPCOeXoMOYGZ4CGoygx9+sArCuKNyZfjrn0scgZhLwH629oLFc3VV7l2VH
3JG3Uv6QG8Mfg61bMyuA+Uds9fFZ/wuN9ggGya4+A/RwcUBu/u6+f1SjXv/y
NkaHm5My2Q0/jqw8uPXwbvNFrJES8BSVU6qb9TIGcBznQQhWjcxqosDAtVjt
+PoruFOMZHetMLNKyvFYiM3bl1KgvbMxGjk/KIoJFtxrBr1uQrb6+5PCY64x
kQnAEMXSx4aA1TWBElMOEitmFO5OWOp0mwE3uZREwhTKftIgW0kb0Bn++twp
9M1aE1Z0wxBlrM+WFKE5OkAS/J+VHcfYfU4GFPdwFuG2VLXj8JI0lUcKDpH9
E/tzBFQYPYI94rIU9vxHczAPap2k61N4VXGTbmqRp4qPODD4yO6hRU8x3Hvw
BAUapjKaj3AQvQRO54q1AwwkXVLHnrrnXpGsp7+ZUAlVDmugVeiOxK0sRSX+
dlQgi4bOf/EUh2Q04cUWuj3MSX5BC0BUm/PoyET2caB+a0toqqWgI0rmMpmA
YciVKTR8YEzLkq+m8697m7GAiWzRKnS3/7jkzk0UTt0Y8yf0mXHGHcNPyYhb
82bNSMlqfhYoljJpcotSzroxagjl1k/AqP3BVjr1FqBjMqQ/S6fM5iMPGJCq
IbfA6JwYGTJuzAxlD8SIcYXPVSsKkBndJlBkMOF2DbKLkt6IZ5qjhaDZk6hu
rbuOv6e7w7XNx/C6jW0FjgrZP2C9utPWCVcbyaOWazJiihXcyteivWVZRSl9
vipKn/AIKPPEEz9AL5E7hRFYbhjNKNHYtMC1hw5QGwotM8JZLAjvFJOi2bfB
PwQgjkn8015srVlENg3b4sBETHDofYHtzhNbY3hKAnBOu7YU+DZp/WwTbjHT
8YszuUpZ/A==

`pragma protect end_protected
