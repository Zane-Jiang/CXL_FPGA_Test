// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0rfVvz2HqYsTf80bEBeLy/ioaPi9xGy1zG5tDXyh3VVbiPEAcO/UllUBTuQ6
YdskFZaYp4ucZ57Y1Iyu7AE6DHRxQ+65AyXQaxVjfGzgtDdOjji52ipn538+
MHJ0L+b6iGTMwmjdNLdwcogwgCi5BbCe28O5ZZE3n1B4zWVojMoS3f5ZX468
1IqyYqaHHS3URfO3TWRRqZSXuDyxYaZEsgUXwIzVfRnpEBBAfqf8yZhA84fq
0473tQcE4U/kPZBxIvOnIMLOQZBrsB7ZiBM03i/D4n6lweUas4kyLCwQx5Ox
bsddb3jKaC19WcyxWGwziDEDGsCYNxF3oO+qwPlGkw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ROJRqdsPBIgP40ixtFbIjMp+t7ICpc/RCQPUCoolIa+Wv7Kv7A9+46zAJvcP
2yixNEdrg85+1lgHKcAtn3X7+L4dr3NjV9574nvO2UyxUj+TfmI8OI7knRZG
aanjsrcE/10tyxXg6Sdwjr1puGn3KGgaHshszmxyK1n6JhjL/8orLlum0WPJ
s/yeOm3fMXdMuyp2vatsBSHlvAE/CoFcfbpxGbDJrEq2irQR5EZ3lGVZLovc
YFEXcBB2vFpXsJxkuA4UnrXlgoPPg/cki2EJVgwMm82xgNjtLeCTwrIKkMdh
n6nnj1KnbJF9Ef2poerFZ2zbmh6kAFe23kL8xg8BuQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oxne6bm01Bq/k4+HtPMIROWfCYsH8p1dJFyUL1H85Rftma6zwYNfuirxlRVw
d/yYzzycy6RDoS7B10oc1v7S0b74X6zDq6+ctXrn6+GFvZPpDcI8EXnl3xtN
5rffQ1FnN7DaKo0DlE0eitNpvzR1qkOEEpYqLAKmCMSUl/EENbFHI5ZavHhB
z1nySj9H7J7d/Q8F3zKQqdvntgOSfL6EZjfonrr1b2GVWvmrG+PpXaZgbeDr
B0ALEat9zkIyowmo00XUw5PY53wAIDqvUpO5lORxI9xTsO2YLhuNbzqDYqPU
N2d6syFjxvuSpB13ee61wAIjuFJBwwZ7K8YD/P8unw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KmXbb88p6mdDZNHfEFPGc97erDvX2jejWcyxI7a9TxWH1J0xdwBVBbvXrhdC
6F0mLE1Ufn7FC/Q9/KxjLzNz+teHDe0Y/XOjk2j/w2RASFcmQWlrlTA5dbT4
YExq7qXL8HBCajgA8pOCfB6FqCV/ggBMIar8RW4TBsrGEkeqn1c=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
h3abKYSwH1R+hilKvPwZxW7lcbDk5vSqOlliQ8C1ua2jR3pQiHFBN/5PC6Xc
5WKXdIQQRic8t6yh4NXnDELd1zhGBJeXh1KBzFloGtcAQBc2KGDcOuIeuRvg
6WGXtzPa8CjF75mM9MvnVvjDDEr3T9ArRphAsdk9oM90zqW95TclUZNP8w6d
F6maDnyCog5IOv1qvTpyYw4DWiaFI570b80DaEjrTC1VmeWee4u5S9lNW2Oh
DCN9tCmOBPsw5PSxDVS4GS1igqttMgvAt0d3CXAyG/r6b8Cctudz3EAUu16U
gZ48UMgj0KLdEW08oI5T+yLC30YN+p6bUr/Y7D6uFMDJ7D9Ukqsm466l7rXT
kObzjguVmIqzIo3xW44RtdsiLNcG+v79X0mxhUS+8Q+4DpoaZ86kBlsOoKk8
LRhwPlnOxpYTM0UtgzvlFYwNOZYazXa0uWj4hO2G9YY04uLGb7d8q/f/zclV
BK3n13J6zw5mNw8ZLhyja5v0oB2ehU2O


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dIY2u1JRLSACm/iDu53lXQS4p7qFDicQmX9Vcb/LrbWCcuo5hRad2kljjkK6
dt6JZHn0HFYeQthem28OioetTRftr41NNJTxZI7zfDX9mfdiXz3t2B7bIpnf
+1C7S5j5Zlojf2HYzvlvKL23C4RF22VeXWx4B+0lDSjkJieD9WY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R/FRsnCSf2Nn2fPSKYFI2wT8oc3aQE/I4gClpk/IWmexWW9YMdP3vbsYjkCb
UoOe8rhWiJs7SKohMQdUwM7C7yz0lEJdCXg8AKRB3dSGTUGaWP/JLnGeJU+G
VnZVBFTlJMw90CJ4fBuyRHVs9EN5qiT5jvgiU2gO9AHjg5CpaQg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2064)
`pragma protect data_block
akvnrXBPYkn7fRuelVHyZeVpuvthpHKA3Vrqk0pr5A3ewSRR2y8ZaMWkmnKK
CPy0c1r1Lcsa35C4pQOeY3OVyqbt4/wQUhvj8ELm3jogqZ8Ps5bM2e/yenp+
LZv+nPKzKAtq55+KMBjx1DcRwud+wNTENoTPIxOcXPsyuvUtm3WT1DyiNc3c
D2mMdz1dLMCugEhkYR5mT1AcD9LIHnTNHYa29FA3pLlQ7GeGH6CLdnpgf2Q9
jpkzm0GWFP62B1shZgtkJU5n60oPMuR+SD7r02sFgUOEHprh+hOGbS3yTDq0
OKc1BRQD3ciVw6+SX81lhG+cBeXSTtYMNyKVFO+dBLdapF+LnRG4nNMtAYjN
vK5xbjNkmcLgEDob1LX+9970mo6pdELEg3OS+n1os51YqNzfOsbGi4NEh0DY
MRSXi8oJDbfKBCuI3k55GwnEcpoXouuFew5DPuF1czUKTmlNyepm7zQ8s8Zm
i12YPFDhAIAo6G9wTmV5eVDg0UvfG51mtLgfLZ4p4zPrXiDeLo0K9zJibJ3J
2xsgwVCK6Mir8p3TEBz50yL3td5VOY/BjSbhj1HKyQgl3kFjm6S9a/WPPtvZ
JjOCpTuIF2VWZvimz0D6zzbcYkzTIdZPmxu2sWoYJsNdR1d7BFUWk/LebjNw
P/RO1opT3PTclOSwBqqBfFtzdpIPELlUhbLo5FGXJ9orJGxUZgMPbU4zKX7C
P3/EUt7eOOEB2i1mn9H9/9bel14HZFsOwb8LcqrUdT6yYO1rbOkw0DFPB9ms
ahi4s0a7KvyNHrccPCa3hBLNjMMQnjSEda4kKhrWqO8cE7/0tzaLwVbSa15+
fkXKxWnTbyfTLjhsOughdtu54z9NIHsAPpo/tyvM1lGRNGrOovogkhjTkRPs
HlJIFvRz7V0z20iEjQ8nwRFNYY9eq3LWY/u5YD2SzTqmQp4qMh5f1YDHSkif
kP4OyaMqpxXLd3zb1VOqDIm+Og1do8btclJZmUjNcRHZaXs41PzQQYnt8W0i
1AQ+InTYEpV8UNtvQk8CIcQBbF/1OvlMcLq+Pnn5D1b18vQJ55/qf3KGZGMO
E+h9iwdJILKhMtIKsmUz5LoPO35QAm4mGCZ64QPoLbO3if8mZyulq6pIeYtm
vOqBUGEeShV8sE+EH6xCYbpUcvDLj28Y4NcAX5E3HnnMbpQgpJ6Wp9qJ4dKj
plSl4/sAHpGfK6gjo+OFLpA+rZIEFnS06EqMAO4G6uUfBxtFUDUP9m7NyOID
Kw4lRRk36NAbyqxfFKAzXtDs8il3f4A3XB1dHZ1aaooW5gpP566unmux+4wt
dM9Vhc0T9WTQNJ6RduJILpNxkGxEdR3zCsNvbkjNogRD72q8i3ag1Lle4GvL
ms7QB0mse8MwJWyWCdJT3WgCRTwVuGJ0ACIqFnYxfgoAxvAm0e64U0SGy4zz
irvt5LKXZI/NIKZ/jJqEYybT6x5mEOCoJWTQ7F5PY+Xpu1t2I0Pk65aUbxyq
TAPZq97ptNIWFRUibkmv+zXFjjUJ271Yu7fDNtX96wiZbP3nMbWFPw845BQW
pJYppgNN65QOd8SIop7Xl73fSXNKCe+804NQP6K2ch4b6UqfawPTxosUOht5
Tq3aBYduqTKZh+HQxwSATcQ5op4zpr9p7Zp+hoaEIZfrGQwUL4qwmfzGoagv
S1vUQSJdCc0qeSybxQE/d+7b0TEYEQO0mB/nLjJC6IVW7nWJJV6r5x0r5PHE
PUUcQSo7auQIavXzmDX8aMKCpYs5U4LKd21r8y6vF1AXqZGET+fvXiNZrUlc
w+W01qT3t4gdkcJ1s8HleBRuL/Hx5pbxPf0Fad2OUohmPui434h4eb8kbTSn
oW1I4J8gcD9FQKyN1p9bkiZg3VtqDamOkBTU3KcjoQvTrPtohl06U2nLR+Ln
Y/VYiyztIDN7m7o6ygv+myKiSgX4go4Unc/rSBLzFM8/1RQh1vGrgtHkxl9a
2NSlqXe8Z1O24vNp2wNOS19s+QxcMlohgshlYA+F/C2gQENvV2zYe1+7ImIC
Ct/2ZOiT3UVl6KUhkbALJjaRHmOluLlMjZ6nBZEzxk881As4rw2aidxPwkHK
VrMvQPwESHQ8nxsERwL0totYpjesqBmO171aT66H0fjsmp/JXf9Z2ZIH9Ail
/d3zTKiU5F3L+4nV2r5+3nXWDy8qPRJ6k4xTDpV7qpqFKW7JxkW0nVmpg/5p
4PMpQV86n7CqRSXZikdyxigr+mESM3/50JA60T3rxwB8BLf560bX6YERFWb9
1UfBweB/lqHWNSxhwJ7xTezCL2WA0Z6S2ZV0Xk2/glVs0bdgNBAORzWw3Wo2
yTbOPPdEmgyzve0wNgMPuyZb+RF1PIS95u9QgFbYJYDxqiwVbJMpsjWCzr7w
NB/mB5A7ekgIA7/2cpQ8OZr+qJSaZ2r2Mr63h5cgtZ0tj7ol3/++23FokHmd
4bDKJj4b6OK+MLBoZmj9qwAfl8D/W2LGN3RA7rFDig5h2IV7KP0MYH69M0De
wiihE0o63GBDS/xCRC3ColU6EZblLyPsnDXxCjYDJFAZc7TJ04utlODlMugt
SbMQG4J/inRB/Xw3GkZ4a5nR3JdnWvLBpqk+9sUM8QWO0apd2r6qB+35XghN
Jfz+DB423mD/sAgQJDPARwFesFEHn5lqf9dikV8G3hjLTEaFKtgglQu0vaHY
kOAeDnWti878s4G7g0O8YlM9V5csEQoa/8pqB1wwxgrUgvLcQh8X

`pragma protect end_protected
