// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
H1SCCWtBPcSE4Jg7FXz00slF5njqIiK6cOZU683m8Tbwec96tzYT9rIAZp8JZr3d
ogchIS8kVxTuppqX9jOqbUmxb1ECMRG/yppkCUWiZwIm1S0/PnoxOmCAjGWHGzdN
2Ui2VwmxH2iQO7ruq1tPYceHi21CCf0ZxbZiy3ZLwV0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10272 )
`pragma protect data_block
/sJXph0wTpUPHYdO1Uzl63DyDxpuEx6RXbL67Q9si/XNvAqyn8FdG+4nrM7TOn9V
niPZSsaapPbywVIDArrgYulDEgiE3qc2iWcdJOApqQh4GYw8QSPLprhahrTsEArA
4jtQJvcv4W4saxF5d29HgiVh+sK5LhIvOtAiLGS/4DaWXEFmFivjRHy4ZfL2DLwY
AKRMKwXBmE3uF5Gc+k2Xoegli6ItlN2qQdLiWkoxwEJ/Rw1erLwj1Boj/JaC4PWt
T8lHqKFWnxUVmMN3K5N1c4V3k1YXQlnBxF2KD+s08LrNXQha8zqgOHHhBbtmO/Gl
TSCcnysDAq3F2kSvlb8oCE8wXPmGylVCvLaBVWE3LBzhUtHK5Q7UBrPfTHVHMMSI
22MDpmCMUdcVU+Mwv+l+S2YEkpHBqEq6s+9FDgJpKYgZsjlzKaE2/Kk/t0CQxjZx
aMYyj9I8d7FWas5NTJ3uLk9gR5TXgvl4Z7rpsly7v0p6TUHUvgDkSTAtQvldw9b/
S6uIcnqDJkDq8NcjZXHVNkh+T+/ntI7XrnGLw2py8WxS16h2pxsoqExkEOcER7pr
t+lspUYugLxYLC5E5gcLROJtTPPIwNrShxUguOuhWN0ocpQjBSqqgt0GLmYEH/i0
BNs9YL40qkaqu84CCWZuZmo+uNbZl8QLQ1AyFwGSCJDeaAkjH+I96FOnIViPdk3K
z3p7X0BkxkTjcSw3BCZsQajH90FJKJrZD7p+P+LY+Cuqge335o7Vu/xKmyiyJgxI
805kARumJBqTcXJoGQ505D5d2z8hNeXoED9sOQyaoKEhfDzIXJCGAm4ijU07WNMU
kRT0HZ+X/dmMUWPklhBuj3g3eXNabgZmYldvBvVGKHGnPVEfbyBqzis+A38hMZ6a
KFyoJ26vGHUUaz5xAd8vo2v7Dq+H4P+RBE+XjiCxjpqwlZ+Tg8VGSpuUEQ/faPE7
K9P82+fMonGl527PqWJu+AfXpDW8vAGVA1cr4GdDdWUvMdMZXl68B51twbWDc6NV
fC+9IT5HPhBMk7Lv3WHmpixVNfFmYGFC0vuGsl/rsakJqhHUt/YEO+EnMaxNDbll
D5sIIwLj3EljequgwIfA+QPYc04WNKFmjleuqmdFAm3hg1g8vlvwTosuaXKwET51
NicEnBohHguzWm227Wl2uFqzp0L/1gMHwvQDgIt1+h8bPUSWYh44nBlTyTlx765j
LsiPEF1EwE/qkFaPK1r2XrCR0sZBHAxqZPT3dJkslro/zViVxm2oYXFVWBEPGj9c
sSH9ULXny3Z0g3PzFAj41ke9WXiMm9R1jSbaEzEApOsjZz5t0R8bRmJwh8bMs5b6
UHnqgcgoz5IeZ80ESFEyZOaFXLfjnhc+2U/I9uHgppuGjP2ar3630/6g0xV6+Qbz
EF98RAlzU+zSZKwFffYlbh1BfTV5xo0ByfNThyS9LqL5WrlVGZoKDveohgjAm8Qb
zARC5OA/omn5gbo2OeMWEipt9LvRH7hwzBWDviLZ1wHu08APzZ+/SyeExLad7PXN
H9JhYuQqZZW59SV8T3KlNBm0aZDwU7Y9gHq1DfPr5IJRTdcc39uhfmfdl9hnE7qq
YYCHos2tsjLt4ugnRIeNuX6ZF/AAjoWpob2avlqgs+8zl7vfGVaWeEBWvwXDNHez
G49aSL77eW7rzBlWDggqRx26XVEB+R9ppNftSCLDXBhcQb9hxbB101nBn1Y75a5Q
/wboe4DFBv2Rryjj863cutZZ9+Dxa83kaktwaFdfDvPZ2HQbP4TiTyvIYd/2ut0T
w0ojD0n9ZEPWEHx1pc+sGI5WLXPoUH4tT7o2X4KG0ReL+8wfW40ZOUHPQxsVyQYA
MdZJn+hDIgyUYrG49uA9LqXgxto/K1JkKn/kvq1I+YS2m/lHxDOgV8FSx0eAd4ON
EV3QoHbKgjonr7XqsbuirFB4MV/Y5LDSzqDqw5J67bylSfkLslBQBhtwIbPGLOMw
A+xEKpCfwh/uJH9IQezjjfegdt6cmHZM67C0LL7qbvMQzhhTqFi579pDQJq2LfSd
jli1MGxB3LaL5FLnadrG6wcGfgpOvbHB0v9Z1GbeolE2il+2pfMEbq09vtnUI5TO
hTpG4GkRDFBYMb051Bn2N39d83inyFm13GRvhjJpkIgSZHHrj3Ff5SceqIRgh+n9
+9L+WYZGavU8M5a+rZY5kU9cO+il6WRUUxr0paG4uNk6IRNIVl/b85wrRFugLcO8
tozba0r5kr8BL/skDKZlxANkuOzE1K6T0CzQRzZXCtyO6Gp2luRabLMd90/Vhcx9
I4q1ZC3PBY7lL8K/6n0cuP3zx7cOJ+KzGVMkhgaoAA8trq3xkt+0EwiJ5Tmq2JzH
tLKacZu0tRKxftaPA8CihoU9+J1apV54IT/y0S4oO0NDiB6uXvKKi4Q44Z7PFJsk
643gFhpZjVEgMwS8DJIlifdyOsi/Y05BFfK/aL3v5Eqi3RvrIXSteZ0V2UvtEI6a
86sxv6so7GmDH3oP++DHP+VxR7QFAuPf+6n/1qI+han9OnVf2GnzQygvo7ZYIep8
JPtQRmxY19JGIQrSfswvC+uYuqY38franUzaZRWWyEG5NTeQoBfdTUC452yfxb0F
Z33nI0FUU0Ptcqj0NYVE4KgEQfMos6HDtliSA7Kgi2dz7vXtrHFBxaWTybgbf+Fh
3YWdJxPlhsSFoVJHGWKlS+vt0G0dyAYQIqvbPM14I0dj9GUoPc/DXd8zIlqaMM5e
cKJ1RGpcz6/CIHbuRP2Uh9uTKlqi2xAa8ELIQmzL+lA0vbBsgB2jR/BMzVRHp4by
P8/txgtHzgWs3iMmmNq4MU0IWBAYo8NVfGiWhkD+JQwevaCCqiiAUNZc4a+Vs6mO
FAXunhLYTALAY9nKRRKqZenems9qv6DxnITAxag7pOnMElY7UJIV3m3yqrSKajNy
lA0I9I5KzULW3skJEkBkT0XE2T9vzSDVfR8OYSF+4IECbJ9rntssH6CApZ0jr/5R
Dcqc4WoGmLKmK3/x82guPyZp7kIMrRY3M+0ZIERU1yOgFu6UR/1ATZTvpxm65YfD
VSdVgzIrqFa/QZuNEDsX9v1uRQk1vaLk71hSHYOdOGXgg2mwTci6fp5vGISRjogw
mJfrWrJPiuXLIp4JL8q6n1s4/1aEIJP85AkzEA5NdFl1/1s1ONHSJdhxaut1l/ty
niiACp34BeWtefV0yCBQ5QxQ19yI/ZCipj58WYk35KgT/JcZWjHrXYbhGGr8R74E
73S206MBvoxSN8XWEOrjTIZ1+5JkUuTR6uSXxR7FI11+9E0ZdhUCdrXsaxYbGiZL
LB/3Jz+Zu/Rig8Pavqy3kRSUH10sGvmTiOaOynlVH3lzu+qXGTl34Ozzfj3l7N9S
PSZV419Yz21rMAYnho6NDXKEtKFfXlOwDrW2tIa0iDETTfSThKKxrH+LPdNiEENe
ao+bkM/YIGG9KVvmXEBuN7HcQMAtJVmhiD9km8R6ydX5EHq3ONXivIxzKZklPsDu
ehaRwEWNxnNFDTAHLDnGnYvuFJgpkOqstQU4OB9g/n8Z5OfCnZpByyRQU4VCn1WK
WdAxAqLkwGlwhkRyRfrOqCEAEQIvFskkLpi/iZ4HBakWXDtVaNzoDIWBtyI+3WyO
cnDtEteGiaJ5hj2QI4w4Z9O7RQSoM8jHtHYRK0qqIwZc6gkZI2QREeagjFN8FmQJ
a3dEl+d6Q1WsLwoW77fIeWxLiKmVnuB5IgYhwikql4nF+afGXBn3XLMJ7BPIBSv6
kHZBCrdzAFjxhIo+FMZ12OatCMmiDE05u7sWFFAhMhlVmJagkusI8IHSwmDZmnyC
zYKbMJqAZVqLM7u48fVzDFKJ4IO9g9ouGBRYR6X8YZ6lUgnVbZVmGsAjYQivdt+n
2udh3XvV1ThMjoT2bs7Ok7/XVh7KS8apxS3/2GlxHGyLluZahBv8aTStRBGqELiC
SzpERq4g8UclEhpDBMX5h3c+EBZExWxJ53kWrwCUcl2CmGtLfTrqVTOLMdJljIZF
wI8QvtGUhP9iHIiEV9LCtDredsOFKnxfEdE1M35M84pWaDbtxGs6kV1Ls4nxTtn+
YfzBco/g0YPrs25kkdolYaxKmqmBSCQoKWqOXLQrCx4cxfmXR2ruPp/w5Y1hRZ1m
4HY4iBqoyGnX2vlAjs/2ignByxoQbW8luUuQba0/TuQtyGjNl36NllYSl6c5Owve
juDMZp1DTwwsVgohvYLbk2IiGXEU70BOQS6dhgSPTc4DJK+e4+ewKhi0B6McQ8ur
GBnF+4z5CbpAQ7JyIcvZ7+SeH9WlEwfsyJHjCTbSivjJOzBN7Tf909HxaGEmjiia
1FuPTo6HMljU835RMbm1QF7FNp1Y2aNrzWCpdYPQgK0bKe0zwjdgLGzpAL8qH9AC
F3dqA+KSluHJc/5C/11vcj4AT5+1UFnnEY8G9s0a3hqYBtWdJup0ld36KMkBHWii
dg9v9ALrKyqfNS6j4QjlRkjINT9lWzh39Wkt7HhwAknQQ4PmvS85BvLaVm3PJvU+
Lta+dh2q47CBPWMxJXwX9FkLy/J7Bl2lBYyfVzZ+9jd6iFyGsBow2VgySSRiUlCX
fsvTBabPWWKBD16o4gNvhlqmvgb2jzz7EGaClfgwh2eGh7Wg1CiEMfOn/FNjlvrc
EsZbhuMYVdsBB3bP/3L7gJOE9e1HOCCglVCu4GCiS6cpuUyRTcbOAIGOVjBKHpl7
Xk+vUEkO1c9zLSEz6YUSn3s2FPz+rsvYsVTMuV2a3bTOTgaYD8oDFMzHI4K2YT72
CrKC4oQG81bYcGT4QnwteLv2tM396uDP8C2zULXbKQedMXe+h7OzQjBcV0TVJ1PF
duJ22ybl4MBrp9wrjhMgH2c6RfBgHtwC4Tok6m0LZJQEL8Tbyf6ZWmB33dK4pvFf
KBOoEeKQZD0e2uALiTEuCwzqPBJdU7U5AiZUbN8d9+0AczkManQmsTpok7ln5uKi
rB4v3VrssJSigo9BlyLgNOmkR7tIYb8pgQfL3UStiAq73o9khHWYbHHIXZkGvr6i
St3rSGjjVmLBZHqepII7q4Ag85WIse9z3De/9F0QC0gW1XHjTH8Fl0mLp9g618Oo
PzIsFHY10f8wzFPDpTyc31f4aBMSfiFdKBTye4j1LyU572HnXwX8xrIUs33mqC9m
12xMQAA9hvT0QzrhUjyxJRHw9dJNUO0/CvXKZLn+UqWWqpbCKHgWJH2/yYtUGEIq
GF5wggZuoeU0RUzP5kBc0wvaQn7nFEOGGLV8i46okL+dB6u+yvDLjyy08Xx2ms+z
D9VOjDaX3YJkgbPjNiwPEB9U2NZVDmnFDX96UkCmvfn9GJKTi6xg/+ESGGse/wTD
xadYeKwUAkc/aokT3GY0Z5bi1iwUbkrAE9LiWiTbih3kqzD2enco4i9r2xRmWgvM
x9LcnrxQPghiCLPhTgm4/fSNWatJHFGds4bCOnjWkWBOHn+rHgVLGWgSwEuTHMN+
JN1OwB9ymlnPVJNc7XdpnlMxZV95Sd2ZPfVUmf7P750ljlEASsV+ufbv8Dz08rwK
ZaRl42q4qPogZwjVrLBmJTCqs7Ogq9oJKvuhFTez9m0kNGWQGKO9fK/iiCJjwlUG
Gn0S5WuyGQ2R+2AvhxQ1DbBBHiL5CmnFDfKRSQBEY++zdrsHC+6lkc86OY6KXQ66
TZj4ctv+IsF4j0kb4QWiQ/yhZAXLr8W8gjw+kF5UnT0gIqiPLVJaOpAkdpipRqGW
SVOIArKkdn1PyUoSHQZtgPudqkGp8J8afHJqYHR/Xz/HW4XCrJE4adilkUrT9osI
MsTz713hdFovCjMO/iQ8PZF4HRQT9kZ0Kce9ICZNUNxqkibn3l4ZEaB2VANTrDAj
egmSl1J+ciwyeuCpp95+h5A9GW48vIHgZO2iZAoxTZzzXEsgSOTlWxgwk36g8BqS
sbEy9YUDzVdSm3s9DEAu8U3QAHPnQ9cXHVANFENaeR8H5GGkt00KqeZRWt+TFPsl
xaW08XC1jG7ztu/5mcgG1yowqKD3JLxagPEMeqY+pvkzEthqX4zEdXw5D2k3cyO6
cnEe+6Ya3BX66ISaaf+4MmLZnerT7wIeoWjkWqmWGSNinbBd3DVeV9RQgDXitwwl
+3af1T7tURk7KltuyvWK5cOCs5bfOOIqkaSMLGrMFoobiUFfx6GIBDHE4d49eLuI
kOD8/7jYgkLgGiQaoyb89nV8ssdPUQIYNfjaGnVgB+6MGXQCn09IABQeCekte4AN
hplovAZ83z0zOT5e9CgkXeyk0rytv7VQ8/NbvgztbHN/ehPZCx4Okq7qcTiAi3sE
+0wXjY/N+3NhJSFcoJh1Pp3GjVOoZF+2w7QPOJorIHQVRxqDK4drweq5UH64kUZM
qNpJs75genTILkBKa/5flnDRJkRp71101p+d/qPIzjkUA+zbIkjKhcgNtKg+pkQQ
kd8PTbfdtYzvTpGntC61Aj0AFE2wsw9f+/R6+yZg/o5kwDtNHJboa0kDoZQuiPgq
nB/wsxS5tBVlxmmswtKSNj9Grnt8k4lpz0cYs3yvkv+WKS8N2rROg5QK8SOLsWXv
L9Xc9f/JXgv6dSSBmuR56uQaZ55wJ6cmuzUUp9j3noDJp4qMC/QLSRhJb/LD+gYq
T1sQB+lwKckyXtAgD2hWNvqs0gYUMAiFLl9qUJzQDhzs9jDtBjl7Rn9sE+KmuvYU
b1Hncn20qhVsCVeFsWkhFmKveC+oXRCov4jsCVuY6Vv8T6KGs7TKLyt1zJfPG809
JkvY9ims8pXxSNBrBuRdFJF6xH9wRFobg0cmZ4knjosNz0fyEO6J4De66LAVJqu9
QleYLR1zRJIi9mpfOtIgn3ZEDasY01IvwCn3A8UBNQg7+F2Mg719FglYkRQnv0MH
X6zDuGInejt53BbLU8LysW18RVkYy3FHW4zC9SdBcUrsrECC7pGh79bS4dO2iv4Z
zWFJJ1f8hBrzj2SaYGidHGHYwM04QHql8mtaz8bdhMCUfCyI6WaoWemDYSmuUdHE
M212YPOtngcOdGythJspVuQ7Np6Qull3Q6kBDE2IJa2W6bTOmaWxvw2RQwCny7BO
eMNS5/rme2cD7uJNmYopTziilK6p++yqiUzI4LnU/i9gzY9Fg3nK12b9xpXZwA1i
sX5E8oikHOraubT3IbNfdX2AXlPhQ+ZeVGkuUVs4H9uFm3ah0OSx7s7alKX03pCK
CrwEIUMfXWQJmU+s7untccgbQPB8BqnVSMBRIr3vyqq4VmL23Qw4g1YF57866A4i
GcQ5otLG1XuBrRz+rMu8vmAbVUJ2LtNv10Fe+Q0MQd8qWpvTqqa1/lIhAnt9AdZ1
/oMkLDQiWemS8AypOLvUqQlag664yfe8gZtPy0UHyEv8cCaQG1foJlu0cc8xZhEO
rFpnKhB3sm6UnSpVB+ZVrN1o+BiKEM4+bTxS6aCjEv51PVj3xiRC+ptzi1DHoBml
KBKA20n7lP2Pt1kAMiOgVW6ZeY/xNoEMN4rPJ0mK5jx1l0vzkCwTn9x78lyNIVgJ
A2273J+zz0rrJKR72YLeSDA8OBKhLwiaNDNl4S0k2qy1/e+n4hU9eHqLPQClXMHZ
3GY46ooYtzPppeVPREAYzU1JaKkr9dvD6xAzEwXEEZXUWztFYOuq+5HaM4+8t3Rw
7w4fLiC0grrkvN/QoYIimf6JPz+0BbfFHXG6m3b1K8sKaMhIYiC2ukPUebhg8mLQ
jPyDVTUuoAS35NbcHR/NceTAuVwnDmqyDTMIWzxEKIcBNTLW18aO2VxeHcecQXUe
Pw3cw3TOtbPpNiDU1IXo7qn5W38XFZD522pqLQFSAwQCSvFpZ0RQdnwUubjrBMXN
o0Hl/8myICho8UIMvKOU3znBpOLJISHCL4hIpit9DjPRevdbLACmAxfZlwMMHbk9
T+waJWTkTsw2mAOnymcWoIPSZGi1+Sxxjo1cWS90SBgwoVp3HeMOWUfJX9cM8sY2
m0sxp/bePjHUocKlGBMr3hDTx6tW5xfy8wqgC8slN73Ol597ZuWcLgZ0aqL4NzPE
Iu723Gc+qX3WL7VB0ggD7ppH4Wm+i1dFfqBz8o2pHNdEEZVpw3KNVxFRBB34TPHE
GW7k957q9zh/EPQHfoT65t9lv7OimvxVKCQ++Yzm5hrdpY9Y3Qxp3E199VCa4Zsp
1s953dyI6i9Ao5HqICK7tCVWNSIXf7mABRvJGK78gLiAyxgfHvtL+OrXkfkvzDmi
zlL3U444rjnAf76Cj02DrXi9aLlCojcjtNmLB7crnuMVxNJi1XGOs99uVZuxOltu
raOKR7qRnOxVm91gZIVyzNSJ/CZrOdy7GrzV51/6J2NHqD1uTPtBYu5nC00f6N+F
bCr7RABIobUFlhgyFvnvxxBS3yG8eLfmok4FsJj6iWlRv39dPZp0K20UNyrAk5hN
555lFRaqHW8JyWOib6dufxCC1n+YDlzh0bXBbSKXwAuCdaDGUfPDxp0UXc8/J+GR
3FYNlrCqmatFenKWvRRLSwk0uJFF5ChqMzAOmWdYZD9ckhAEBJr11JeXVKuk61b8
gCv8sbRsH2nvWBe4DN2kD1sv1b7Yb/CK1zBIY37I8FUpz43a+ZVFeyKtuzXmlb4F
ezb5y9vAISsl9uulbz+Kz8ip1/mK/HjL1gHCv9fVdl1Dr//zAhaviR5Zeu4Rsis2
qw/PN7wJ8BRbuPecDEcNSY44tDBnuTwoft+dulFLAwA1RFXDOf5YneTPkx75PBPE
9RcIj6oFEdfWyDw8AALamY4fzrfyiGUKHpVrQaWW/1lRmnW+mVE9+Hb0UvWnQ3tT
IAfpyWo/Jis8siOxykRepWNCVp9wT83Ft4Qpssnx0AU2tavFoVMQd9roTexQw1Pt
9wXxyt12AQ3DmhQq5qgpLz85h8oR/Guma7MhzFpsU7ATfDx96u2eqGO13Kx2rQLc
tjGJjgP3z8fqTnGLSY1FX8/RWXMumUfFWLsUcvIHulU7J/IZrPF1Y0Qp+ZhorwYk
eIxKAhMgs+xowzcvc75RlLCnw4xCUx+2UUbAcIfDn6SN2aJuqCqxHHzIL7L/Ik8l
08rOds1GwkxVQ42UAci8uynt/iugeak6quiaShkOEcmmE/fH9IH0BSEV1I99SBZO
G+Rq5fE+ARM/nyDdbEfd2NYcJMDCur+/g3pL2/x+Js8GZu2/378BCIvdm9zRX9Tw
buLCLSrcT/K2qLyYAOUN23Sfd6/EtaT8CxQYUSZdKBDJKA7zLAkKiw49m+0JeuaI
aupCJEG7M6uPb+wOpCkrv3nA0NGylQfe8yitCXZOqffrM231FRaxsI720fnUTZHB
3AtAwQNUL/Zfdo7LEt1IuEp94/q2en2PY91vzvLDZ2Kyf3GpwUG3GwMbuYKsCqHO
Wpdz2nAPpTqIiCA10w0A61i9ButF+zBdCXA7biVtY41OkpMZyg0Phz+GGS/meGdl
A5kswXcBRAAvNmL74RZQrO0pgIWgVJXhyyb7chi/myT256pR2Ax/XxG7U4Ery1j7
LK60cd5hvJb6af8peEczye3t1PgZRRHAfYy3BWR8PvBckRV35+Gl6Dg+5jllVWDD
gQVUTJmPg9PhdWU2ANuPZTPOF2zux5szlOBKp8VF0G+Aj0X9umYfKcnDXNvD+jy/
WJKSfjlnCznW4Aa2m4MXy7AuHoAEioV7UDxLkGzmm9mENjss8lTd4zqJtwwIP880
yWfXv2Oxf3WfpPCZrhI7zG0xgBbFdbN0KdOiUug3KRLrOekgeBtaHDIUAB6IbLiS
dIJL1PJyZvfcPaz/WfY7LcDDIaqFlSMgbitUFainJelTSKn8A3cGhPcLJNY0kJze
OFAC3AhY6Vnho9pcr53E+sygNAlf/AzOYno7PJFlvvITMNKGYZlncgcN75izHzSJ
w8jg1ShJcQuNNWRpx1iyHRDkzIYgs9I8i6e+Q6jSqoQqlv96D9oHof6vDVCQ/nOs
UYzIlWiKLftn1zFTL1FveXSGCNrBRZwE49bT8BEbv2ZCz6WT9GeUHeeK4Q6ZVL9q
FCeiC5Hs64pBHcWRw+7BUXz8qU8Flg7q0BIog1WaMN5YC2/oHgPLYUULFN07df2o
A4KZvZMjeJvFby9a0ysBG1DMUEuQDNGsPGZ8SuPMopGaMH8XoGBD52BWSvdCizWG
HqrS3Els9qpjGW6lBZWd12OBvivUVnPSJxpX2pfETi2XdaVxTRsuN2fyVB71kHe1
ZZcno+OCGED2TjhIbr9QaVHLc3By/gJtGy5Vww6iJ9LpRcK77oMCwneizO5fT10o
tiA/0AnhxC6y359v9Xzm88xeMiaT3EFyy4ds8ff2oaZ3qiG9d9GtTiaMu3wRXk//
bhpAF2g7CY3Jmw9Oi/HLVd8rxvsZ8WXflhqLKA13W+h9EdwkgXkDt6xzPC6EEq4i
wffVCdJEi93aELhuD5TOyBb0bzcKO9vNSFgdU9iWvGFEgdtlq54Ue9sMjFONvrDd
jwOi3QznUZbJGHO1UN+xFPSif7L7XQ1geJVfndQzRsUD+y/p2B5W3rl71t6cGeZL
e0B45uekmZ7qieUfN0LxS+BGZ/sCcEEbzKKXMo0YrerVq/ufR29y3TOsK7fmgK1q
deK81O2ahDxXUgoowakFbZ8XkMB4FUaVbFx+tolMCXOjG+l8QP4TwI38kRPZiGJS
sEewt9ielniSO3fXjoC2tdG90on7Ew078Cb4OZwhE7zmabFLzj9EYndBPctH3a3S
jUPB+d4nwml3iELbt4MKbtIzOE1dMxY3nUkV6YhxLkTkOTJGzL2goqcdsl1sBQCa
e3qVa+aKyiQOqhyoAy3QysH06fYhGZcCt1Ef2l7uISdEqFtjirDuIISUcUhlI5yU
AEM8fgsgUZK8w2aK7a50a4C1a1xtVBLkZZMiuRWqugTji9vnLaJMkhgn6Ma5nskE
k9g0JTkPI5Nfjx8/CaQAVtgXMF4cFyNVr6TvdwDexl5N7lFjDQM/i1SJgVYuT71C
aa8K/DZb/TXr0DFhr2OPl6JgciLSGxiFCXbvARi+W4WVanO6RzyvmH/BmiBTeYsI
tTmsQHKSbnT5RVyzBCkAMThlissa+ux/I90Y+QwCkSMnOJ3VklBdMV4GDFu1jJ9S
gJ1a+lWQkQEMOv9BMR2CBtv3O3OPjJapWFrOOl2qPnfBVyKtmFJTHuz1HVPlAQl8
S2mB0KdzQHooMUbzCX564ZeqGLRFk5MmZ48V0v9tJET4cllMeLeDgomy4KFojus9
aQf581zfREMinWmn14OGkDQnT2o4/SWHSzqlFEWdn9Wht+bNY8LSQ5OOnurot/uD
8rfTtVCsepxiEBKjau0dVM2oLqmRzZWwoNTVZ7J3kShPu4SEDG8/KZw6BB9P7Cdo
SP0yPxUxlFN8dPFNcE1Df9Jmrmped7oiJnS1Sx37hyk11NDHWQxlW47D/T6UcPgY
9oA3rzmNi8roHgRZCXbiX3O/Qb30yrCWFB7xV8l5RTUbXhbV1lME5GZ5mOYrFsis
kiZODqZVjw+QG0pUUjaCPuwfVxKY0p91E1XERaBOi4CloTs0vIL8NSnTiqksKh3Q
82OqVzk3aFUeB0FdYCNTa+T2F1swugHnf1yc8v6KR0M7BF4TaOb5weqrB7cnJYGe
8Wy8g3GSLQxasM2tK1FAl6tr13ACxOnhhWuMgRvHf/rQcs2jVZx3OFY/SB6iLdBO
Qchb2QLP83mkJEk5xB6huQnp2eycNP4CHxyir0TO5HihizaD0sN4J7VHF3/LZ1d1
yzwoItTfjQato3/mCFf52LLsqQT11UWKjPVokL6IM0HCSnfXdgFWhTQPD3gt4DBA
ekTzvDdJnO8U8I0ui6QxVMjtYLfV9nmphPqWhZFP9BsfnO7nkxJ1qovc61BOQ+Zc
NuBQqidQjCkwWFctF+TiGTGEC08PP+PslnG+FtFGxUCF+VJujtdYBsmbf2ISYDM3
vSfS5KRT2AXLoyiOWOqflcSZENcqUE3qF4E2LPNHzPAubAJc19rtAnU/GBQpjB89
E93toc7YkkB/T438tx+lVDObV3XIhsAcIorgT+q7K/y+gaJsz4r0HrkrHvdUfyZ5
cT5uUxM6IqiuIEtIRF5gyHs+bBUNBj/2Qck3iKNlLs76CEv1704I2O2KQfFMnrzW
EkKZGBxtkfeCiCrcYot18xlr+pRr+/Ph+gP6h0gyFzvvbZLP05rY694dAqT4KLW6
b2fFJCCCM7KvLV/u8j9aBrjn8aQGpynKD4slO2jUNV6YJfaF/Zf5kl4cYEOHHh1g
cM+cyTr9nLlAjW5yMFTdK22r7MeZVeEK9G9F2XUkqxq83uuWTrcx2htWVvdTxNyu
hPqtnmApen8IDjqowBa3atGkJJ/+UD78Q9429iZ6nIE7ASrp0bZW/TwcG5IYMpeb
ub95/Q1Y3gVMey+p0SkuRZnotHKrQ/Xl00+YpGe1PKPzikx2QSZ6P8V0cZcu1Vac
tmXO+07AjebjdvKRYZf33kBLl4P7Q2dRz+DuepqOc7lLY3igqSmJVEI1ZLxNkmEP
sbdGAw0/ALTq2Yhkpg9PIf6da4LEJBcXJyX6ZDrFuP6c7iDG92HxybWhHFfiruW6
bQkKEibb+OY69VR9dBnF+wwvwGN63pZrquprz6pOmESvUQhcwE0SK5eHx1Tra9B9
lYAyW9V6tYiQUBfnUe6Hn5tNq3S5gD8hO4xOsX6GFzW6Cr1Z2YFrFGEJloZY4Id5
1aJD2H0vTFuZz88wTNV3TmWPfdHSCuFeVPAUi3gNEnFlZCT8HWUPVxrEBSr38lA/
dWzX0lTKnxBRugC1nbgbCYLKDuL8tYbIPmpUJIs7T+SJDTdZfHzvBVpaZJdawOIC
VND/cTgVP01wbVkEKUZPArBi3/FxigLlFXHf2gu04jBzNCHlKfIw3dik7+un43x3
+uE8LS6rt7cTedZrvGIPPeF8G+9RHy5H0DDYKF1D/yPgHbmID4uZNZc3js+N3HUh
qNR72oHl4QWXtvd/w4qgPTp5ELtDGUPPou3r1cchI3DQ4TXQfKsJbVcNo5m1Yz30
iwphaJ2hAQNMtdcrNn74IgqfYTQXHiVE9AndvJOcnaYvvwgybc19xWUAA8+MsTft
w+Z1zgigFupyMT7NZgSIw9CYMN1pCwRwHheE4Gk/FdMbLYYkNetMSjqAvVOShaJ6
9kaBB184WDJTLtaYJnGcoId21WKR18I8N6gOfSpBwExhITCdl5n6XzbR87tyV+bC
iSU7hJv2+0c/2REWwQ0wMOmoSHvk1lyCcEYiCgsF8LNfNcCY4uD3VlT3Kih6J1jK
JWSzONMMSunL96qI62bt4Cp+N11Z8bqne9D6pB4CYFqf9/PNl1ScVffsQsjcVWGO
vWxaA76aOcv5DT2vctXWOhBMnOupHEX/DKT0/SkM+AU6y2Ys3fs8uoH02fRCByo9
GLXPAWWE3sR+Vq1BzxTcrlRrKAP3FRcUoPq3beNUVrSQj3QSB8YvbUx4H7vwvoS2
oNYnffbuJqOWiHub3nA+0CMj8OQfYa8AFcbaA7BESlblVDZ10IJouSHYgvG42g44
oDwrU4QRIj0RO+eOarJEvMWejdh5rn27ztLn6fhhJ8TLCPIrk+Lv2sIg3z3rTA0t
iAbK5rxpv+PHQFIruA2KoF1DOv95C39aAVwmbnvoueIB2nksMR3Mk9+X/MsPzE1D

`pragma protect end_protected
