`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
YwlxuNXjkGJwj9GUDos9Il41awTvLEKky4zv1Hsfehy7MOT+4whkimJn0O3AXnpf
gXD5nlLiWZlW0pXmof4gRelSkY32e4d1MLmO9Ml/GMdkk9YuH7Hb/Q1oyIfybhl3
1FVUUXa4l4YA6IIR3eQTSZto/XyW58JFzgmbKyYloTY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 7472), data_block
1ARrx6M/GmIhP6NaOCBxM4C/Vd3Em64iZljDwKvRL2cGEY/OYBHAmMaDCNYRaGol
uM36VVkoP4hkT6/AcVw5s1LwqWGFGL8qxRpt9ViLfG3LkY9nG0YOYpbPY8KYFQ8M
ozJXVNMJrGBSRg5LlsvvAOsBWi3eWx75l5rADdeeR+q4C4FOowxMj7UrGWfzr0wk
2FI30oiJoiEKS4jD+7iBbSGLHgIT8S3eZvp6iYBxNh+YFtUjMZmzW33urqY/i4ti
kBmk3cig/5RXtKwETBw1IAWCDJ7fOHAHuWVJfmBNGpNe06SL2gyZkhzzh1hjGHYN
MViMWVMuYn7kkcn59T7Yd4OXXikw5P0zLW8SaIhD7yKY8LN6zE9yV7NT0ZnDp8o3
b97M0e/2hES/oj7aw4IrMOn+tldVHN/Ekmy7rys8CC/8eT2nSVT8QpdkFVP15cix
zcpDN74B18JpBIlXol7OrkYUhzeaitVV14dB9R7BF5SRz2EozTAmlS9WOo8YVrre
zEMZsr0a1llgiQWpCUj1yaibID2Qe4HPEYOi5xo0HMfgE6Jzrs6L3uRSydixKwD3
xYYIRo0spcv5VnRU4C/vaYgTc7z/6zpvDza9bBoy64EzLjEI7EojAKajhsRuDB0j
6oH6TSQYH9FmQt2JdVyvprdHZ2qYvYMv1Okx4JL136NS5u3eIae4uo0HzUtpiYnf
YlJSi1UK7a7Fn5e8Z7z0f1OKGU6Hy0chR6CpR1SYsqfI6HYMTWHp7LiDxDZ5aXT9
PQV3z+1CpkIUBULXveJZdp4fWZmB2Z77Fi4MGrnZbkOJ4E3+cMSvqnecsDxr65BE
t+Wk3AZV1aDkqJYQ/cEFri1noHhQ1nGiQFXnD5bFh6RtAckiXR5QP4W1l2ws8MOr
s37daG7m04AMNdxaemIY1k3ltfIBXpWaJKa6Rt7vTtwZ90s1QKV2Gdn7LFRIxVnk
te8KWTuvZKybodgvS0qiJHhmScmCwdAKfj71so3BwmRuLM920Mp8N01GO2W/OUMB
izjfSzQuwoVtJQwciEOu6xc499mQbi7xA0OTV+UDaV28WXuw7FosDRblUc4sid2B
JKXZfKpyBq6zg1quYPTgw1U2hH93W1COcO5dU7YOJVcJ80t3Ndqx3XDBhs86GKWj
PAItJNrDQ0VbBn9TIWVkCz8MGH2jhnaGBkLu623JjOATZOAM5/9/hfdl3Mq+L8zq
pOJavvk/dzkOXYrYGJgCG3OCWlkEp0Dh8sd71FiS99S/q4EwmGUes4LnriVulxAs
Zb8XeGEjkofhQoO8RqBqPMT14VOvBmprBWAmfdHTS6g2yFMmaaMsxtV3vMc2y3GT
GePi+D6ouPenmP3FJSt6aXnMt1qiBvA/WKZninvynnHRNqgeYaUMkTHheQjAso05
1pOAwANEgWDW2WWdKQ6+z7XjdB60wJgJNy8C5zpO8XdocYos7uQxWkBnWNsV5/Qs
FRe1cUeW3jMja/Ovw4HViw6RwXhX9G/dwVHF7PCo0FS9qcz/POybzYc2JNqGGHRK
AAgl6q0eM/pDPzHpM4ONQNFSg5le0idzB//uXmXcboIODW5j9zyNLfnyH9/CBQvg
gwr+YQcnTikg0Fj8RZHi86NF7G50edg3hp/oo9NEvUsozNJFODJUfKcB/950c4Ap
f5OgrmUmr8eXNbWlI+sszrLJDUIQqumuhaV0ITRUGjpK01z3PtXZhTA7bifUfBED
NeHVCPIBcQc4PAJiwvzMi8fveiN00NhQjVVf4HGuinVSTOxbQBS6JNEiucL8dO94
SlrYH1F04mIBkRpRGwhngWRYNYvVyADc13vHmFZXR/ZnaEbKuBVGlCcjrXP/Nu5i
TeH+HPzroKeIcvxTB4C72Ju5GuNP8N5QzHFLw3MJKLTRyaMJIPpcFqgKeSypGB+L
BjXtD/2SLW6KMIpX7czuY6qEIW8xR/BtNHeIeyTGA/ItcWeFKtQ4wUvkKuIxOUId
u/eVJEpxoX/l+HHA4E7fxoHYd4kUg0083Lqmfaqd+mG3CDTIE3ZVv/YkdWY8m5uy
FLH/TsfJhVNnL7UWxxQ6TdqpZxEfQqhT78QhPLYFkmq53FBCxDadCtR7ig5BdcL2
f0ZFRkWefKFGCA5HORDP4H8jNndDDrznpBspo135BdFdvDHhgOdOH0fWA9Bd59i9
65by04hMs3ZtVGtupD439NoUOx45RKmkFMTxJx2argFCoezbbZo6yLLux49c7YZR
+6K+hLWsFTEyq2s/fsiUvhSl3mU9yjQQxgt1Ucq6koAq9BAoEILIlQx41We2l1yF
e+6nS8Ti9XEDdQkOok186Jz2YWqvCSvqnaKdUYBZdNXvsURu1188LcMHUL0rUIed
e3ayb6e2GXGXg9NI8Z/zahwy0S1KkfxY5FVCevGR2Fw7yyE8TYQSZHE+SZGuCqgO
x4ITZia+/P3ZXuZo+UK+YBGwt0gDItozcvQUptEgHMWXSuQziWDQz1hC6Hyk+Eda
Q/HnrOjx0FAozZoFKsUPNcmccxGsDR9Y8WQ/J08gMAIKz9/cDAZfgwlg3Xfsc7OX
FJydydlNz411tuOBAn6gfQ7c11iYvdNxU2w1uSAD3+L9ZDlDHDjCH8AkigtWMvUo
7f9zjH0Hg9hcMK7OQ64fKpgyiIQBE/joeyiW0s2vVwv6TrWMG8WKfiYNPGtr83S3
f4r9zEYN0En6vcaF6l1OXdrmYxYKNNyB4G5cqrSf/M9LTgafnjDrPRzD5Op4Y5YJ
ONBAEIrZh84SLBDRLWchGpZaBQzBSn6j3xX0TAVqM1R1p2o77aq//uTs41bGNC5g
lnjlboUOE/HI2J4bRvq7Pi0ufznPRcJtJdSU2RK2Yf8xu38IELZ+w0lOJSmHIfp0
cFuec2U4NQIAwgyuijNYL3OqNTzHtGR7JwAsL4fjc0BrFkFKfRq1dF7RleABdJFn
zpSLmBroyMVFwllRwy3A35N/bv6YWi5kL+UCjYDZn7jGB1mfiSvsoF61z7nref6n
+Giwl4/4ixCkZmCiTQPN5cilU7GsGm2Kk3Puci49GYwa1B9SWkzxeqh+FsvYOKrD
s5ZG77Pd2V4gDwY/LSRxAoJq+qXCQ0jXpiP4vBvA9IH8G71N4LpPPWlcvLlPwyzd
D5MLo2yY/s0dryeSe1E4At4vdX1UjFWN0znvsMkryQu6bQgAlld1zW1GB8zpFDAw
bpcp+yzwAIUr6fY8UWLnODdTD3js50gXnztIMi4Z0u8YMJj9jW5BA6/sceCj+BWa
a5Wqe4FdtBmDYovPgqrvBNPRita+0uxOJsxSdH8TvmiD5NSkMcLpZR1GlI4FoiA2
BkEKkQkDtHKIhB8aywiUoQ9vaje3yM7xggw2wBe1qZkfxXTNq8nSOBea8NLIk16Y
VwNu9HPO8bM3rj2clf2EQtA7Qf3qSVleF0yAPBFPmFr/fQnBBEhfBwmUFiGKhdTm
1TlNn3M7hZp2YYpERmHJO1obFaZfWJw2utyxN8sqEbLb05YPf9JWvgTC6ztM/DQN
XjeLPI0e2C5xNDYN4NvrDx07F/9djl1V2VHjAjgwjU90Lji3lfWJhuR0oQEsdEAJ
AlrT21g2Tx9KMj3uATSczUceDtdyumA6TCUlOHM63pCSFGFEickDpJsJJQj5XlZ1
OwG7cQhghJC8VdyWYIfqaIoPbk4DG+Em+DA1bYWlHbofhQwYprKZEUFh8ObkDE7l
jUTnGF+pDAfZ2jxIEN5y+G1becMbXhMtLr/z3DK1CBN8Fo0soorHx9S6NkTBG5W4
os3jmjciLH/TzQY/YDNn7gn5tQShEr6mZWK5TmqAt5AnxhuxK2WGHN31+1fZqc6Z
O0kSfxAbu2Av8T7B1oob0KreptIG7NfBN1gZff7mFOJqCa4+Lbk2PhVI3NN5uzNh
1g5ojgNeEnByW+126S/Fj65d2OSvXq5478n6+Nb/lfQ7hmhAVNVeaP+2/5VeWC51
JyUSpSH9jX4N0D28zjZKHj9gD5l4ZSgPkmHa3zA1Drmtbh7qsSrsnYkS2kQztscr
kAK2UOHokTPFbZz32ASx3dpkp1OGFhupoUSX+cKvQEtO2XAplUIUdgGa2QYAzvtL
k8JwhNUzP64HwBQcfkVq7RlKV1I4AvImSnkhaQqMHTqRdq/NvKJuJgyYf80DPDF8
JS7ToQl/+hsExhu+xt/aiuMfCFYmA119TzBKcoXdjyp/DYgmOuc8L8b6jDkGeFyC
8Q4Y2BrndG63SBGKcyvvjDYUL9v54nNkkz4LwmctUd1q9lM+Z1+iCwzbbJiLZ7+P
+g/dXfYNKc+ajBMtNP+BFrxrsPtML7WyInTriday8Tb0+SCn8EQIBIHHa3S+EpwY
0TxhpU5JacEJ4c3FrtDN2K+JO0iZAMnQHrvBO8jMPcDMI0jC+E5/cq80fEgV9/Xl
Hs/9UlxuhRmgQXlcgHFSV/KgH0gB6lxycmyAY+fBdTaKFNeCcB2EGleArQhai2XI
Q7AFbafdZ1GpfhoPg03JujomJHArsvA/0yLky+CsdiGC65JdpQ9Z2VCTKrTPkQbK
V6z7DNjlfz4jFyNWB3KOGy/WcZo9J489c0sVISAP17HyjTvTfNaD8ugNJ7nsySRz
bWYzi8+Iamqpn+RxQlSVZQHFFeHbUZ9tPRtnK+fiuDX9C0Q1L0IuyI/4MFiIcWLR
USYGK+TC3dz5Ceo2WWUavXFWRP+GJ7s3DZpVWBK3vfV1DL+yV19zzcD1Kvj2u2Ns
8LT7oAResSUkYoMuOLm1CrVoDc5Fyan3miXiVKT475rsv1Xje7L++LFYFO85alq+
S8iBhIx1oj5K7xfC4udtokIhztBhoGx+/xNaCZ5e1Nl6XgXbBgGAQYTPf+E9RcZq
vOOJgBZca+hENtcAX1b39OUT1g+Pzims/0IFsn5DXhdIIuGVyhnxPXlrrFVFEGQX
cqU9idj+sVl83Vx2LKBHzU1ADAk3ZTSH5VBiQPUDbtFmeojAX/Kqc2ON4Du30G6T
FSrGDIrE7L5yB+1xPtRYbDTOmPYFI+SAiqjVXDfVyRTfWM+pX7GdHVf8QFw0jJzp
r6lkydzm70io7TzIXNr3lVdlm6svPbYM1sHmDYCCiCdBdO0iXBWmhA9Jnu5ew9ec
imdXu4o9rOkTqZzra6LqghDf7DxjaQEpSq/C3znsfD/JRaCDJ8r7iqYxVomhPUaw
Z/SUdit9ifaDv+V5IIt78nf6J9x3R/TRzZcxgjyrHBChBmEg7JVWmJIfVw6gYyDE
fN5gl3HIQY6cuj1P/FOb8dDHUbk/5cn6a9PTHa5MudI1L12zy0J9mjAqqa93qx9C
9zYlvWQqpqJed/Loybx5eJBHDUw4FBEVfl1GUEptOutqZq4aycxLU/yUb985XLWy
klPYXSymG/WLbjfgoTJHD02dryPyyLeCDGYC0M9lBoTyujd4bF1O1vbh06K5h9Nx
B25VJQrTROcwNnOpuWM+KGyER6eI1UpdHjw06Q+qbNIGPPYiFZeiGT9JhL4mVkrW
87+QjUudjqwdLGG4fsPtB6bdrQLh7Ub6Ikbsl4/OCqQejUajKpx/X4CUKfWxUIi1
2EFY80zNHc5DZIsxVovIsLbw/W9Llh+e1Z4K7qeoJWI6EPrzPPCn9P06jEWmHZXF
2yIq1NgTbCHzdoYSePrD9tVKjEF0jSp+fKsTRyY16QsLYMKp7QHpdQN/mUzYk6Y/
oKLNG7hUjtANcCbPEiZo6NE6uVWuguybyOEFV+g5yQQHNgeuMtFsR8Mf7kuPMOdp
fBIK5dubjsPMJNGXZZ1JuFxlNsNv/IaO0W+yb07fObm+NJknxcYpxcwSXoKgE/Ob
cYMctSKhQ/2PmSsC5yEPhXlXjGyOGVdmXzrXrgo8ul2SZkdN/MJm+2w/o0x5cR0s
DxLd/iMwGfUiCSPguF4/yHZfuzAXJ5a+QmBMsUtGpki0ON+XnlUgRE7VAOdN+/S0
E1U7DFikMPqZfo+TghtU53CimyOD6WvWH+OPNAOa/WF8XzvXyPGDE4WuqU+YY6GH
nZz9Lxt6JFBnFvaHzmt4uH+MKdzi6AwDvfpCJ/hPlaJqV31tGcUyEbMySM2U25nG
IsS1xjH43/heOTjuJnKgBuR0O0sauJf6DNQHPgAHJnG71HbABxupTsmXOBtl5uI9
lNNnXAL0PHeHq4pIIt53eDpgtXccYj9E7iTkrYDKIP/MlQrTCCfloCqQQB3cyee2
CjCq6PSqEmEyWvgBX2pbpRvJHsrC5ZOiGlWvNpOaO8aJOE4W/vPhJDjTCC/CCpa5
C76A6/0w7emma+QS4gC1kIv8lYLOZRihJhdu66lf03J0wpQ9vPI+eKQUo8KdbJqq
LYABL4HE71ravKAroFm/DoHuZD2NPRuodnJ9+vTBTaeKnQD7QIZqBBFglBOohOwr
stl6QrJ7CXPzabiAGAfUVB678Idru/d4VPGBXKtbKss4eKpkkVmIXeM7s7Bdp+6D
CRSnVXU988dEoR6Bjoaap+Np0v81mtMQkgIFy0uywL2BOLG4uPnnz7ViKITpVcew
n1t7fSaZTPO38/bOhaPJiCYDK78IEjdvgkgkqcuuNKECTpBgB41kEKsVao0cd0x8
eI74IgJnXM/lAMYqaGz0UwTYh6Cn/fTrvBZWuarsg6dJfphHHb2rtFfJB8H7n+X6
FZa5Jfzy4SQeHbCjxhNqlobBwbN0uWrd5hSi7Ecv9X9OKv79+Jo7HQLRlB/tE3g5
T9ftg8rakxDwip9t/iqBBegj106rfIHyQgWDBOGZWCOrMBWwJXjrxn3YjeRB3JLT
nUvvzC8z2oT8OzGqtX8ayRnIwct7hUhvv0NERx57ymOgw4a2iZKAx9ccQAJhW5ny
zpAvHTu+GTZrD/HO4kNXiGhXNfg+ryUQSxcOOX0y0eznxDWM2ZEcB/CcbUIgfhTe
q8CWZL2iHq46IHf2ZccNxYaoyN3uTWhVYPJy4zmxt1U+l3GYE7PTH3stzYJFf9KQ
hnVD51XNeHz0wGKnyqlUr4DzQ3nOBHpOtW1Zr/SmhvdTy+dtjv1/t1w2UQP/xqOH
iRUMnIG6nb9mxjjpElX1G8g/AbRwtU+oYKOYE37Dx4dF6a90ZvKyfC/nVeAQuk6B
sFiLoEETSEKlNqH4Cf0QuQg/SSjHsYMsE/Xa+6KhNvLyLSCCnnIZRxQWRxyXMDoD
NS3iNogWQl4rfr27biXnUeD5AG6TW3JsIeVADzSDM7AYIQcLwld4BFm7fONJIeAC
xeEVeV9d96LjrAoxZzeNH0BFap85np+Jddq0s4d88bAHN3Hpm564XExGWUaQKi8g
rzcmN1AHLg17cEwV2kHfCmE2sLJugjaq6nC1UNV3/gvny7AkaT9iLHz2giwah1Ik
2hbSvKkQR5duzTWuCKH7Pf37fRsu3HOgeaEGB5as0YzeVKoNsJRXJqh4FSKnXhlQ
YbX5tMpxXzV67DnfsrDu7GAQAYX26LQqEQZ0SuX0rX5Ib8dvMZQJszLDgPo/mN5v
XN5if475HlFvMhOFjLKL4lOkR4YTm+/RT9eIIlLfBjnPfWsoqURJ4vsxwCxzq9zI
unzjlzBpn42FWi+RvRigQj6ap1QoexHndVHSm1QNj6sNba5xlC6mpLXgssq7nlJj
2Xvhjgt+4JrbJTIzaCpuBZ7hTEokNL0SoQeKzdQBqWZDAi5jH2GVS2X3gYss55Xi
+3UPhCbGMD2h4aU5M5ZJAHaElUsEuCDGegxHNjawMaHDFOlb4frsXcFZG7TBpfUp
+Q2FDEyTflgbikJYpOv1qL1JUkVb0loKLs8mV19hUrOcunOUnG5odqeUpOu5/MPt
6NsyGWytCQmJY34yYgroDGHIo+PNXKUIdQHewgobcq1op34/4Ec7GPehl2htIJUc
2t5WRB50amosX8aBuJUkP7L4eeJnPvk5Dwju8QdD3bKFPSsj/9ap9JttEO8z6sqv
j/dgMN80RRT2WywoMkPsXZjqUIdSQC9kF7LpD+FS2YgBPeOZSzh6Zrf/6OJE0obe
8WK6weVvesHK98NyyNlPaHc2KJsuyPxdmGOLJSbVB+gqtsdVSPt6mdwBoMADFTx+
pIV6NUieLIx/Vq0Mqzpqnlap2QVNU2sHELMOHOyj4PKkAdmVjYJbfEOTB8n7S9Gp
+s2qbwDtjJQ2XShIY+PyMo/xZX2GmapBzbNVXT8Ggnh7yaAOjMKsHdUUb8Us29G1
VPV0mv1kkR2x5OUMejrxdIA7ukm2XlfgftQBbkAlLVoJI0MHUeRscOdr5L9j3s5F
juCVFnL5lvRgP0Ed7LnEZ225VrpWFoLvQL2jJDPM6I74bDBKz1d/w3Kj+UxWHRJs
9+naR3fbJ+zZHxBju2+QHS/99HIJRbLN791CFgaByeFu6u71DWYDlkVJpyIeTpmJ
A1+6nNBEr7U1zHYSqmq1RNUupVRuDqovlSPCUgrdW9kWyvFG3duyPlKMgISuNro+
atuhqvlNDsRjo9vY0SRug6WpK4a+cVNZ5hTif2nDf8Xzz6QpMJjzrM60WA2bAgaE
QK9W5iLa0SfD4EnFJaC3wQyELUjdvdrPXn6aIImbyzTUWrm4lxpy1ilLAene622k
+zOwkTnUq0BGH6iV5782qV/3Ofjsn8PSiNOay85WPISKyZqI7VIzepd+j9OWO28K
Js0/xzzH7pqhB+zbA0noSyxVyyB2Na7cI94Cscz46EGU9IZ+T3fuRdTGvB8O5B+E
h1q+E+A/MXb+kutO95FMSd2ICUaQiBWuUvHDOkdQ8kgWBcvuk6iGyELy1t73CGI7
9s1II+V9OjGEZ6SnWvimvUCHy0Qfw3T+JFFITk9GkPB6yDeIHzNugIZMzBHXPmvx
F/9ziYqRCt5G8SiHvDsWpyd/ycwKDJVY+ifmcpxi9G1mNYZJEA2Ii7KOUwwF1uK3
tTvRzlvQ58rED2Zk+2GHmUH7Wt+T+Kmlg2RVG7dOtPJGti0zcHUqVVxR8iFGvfWe
LSVah/7/HdZBM6xAOIs7cv4s3jJlFVZyfjiwMrIaW2sJFI7XDI9q8wAVMV0XfJQO
5KHdiYMSAbLb2oF9WT+480MbSvr9nOgEqGMPczkgMB04AwaZfNzGjVNFHU0hXnBI
NeAy8aNmQFlzalKCyyJJ5YoI2qpzFXnPJnyMP9Q9DNGs8IewWSGwB2TyS/MKDlxx
EMFk2xcn/74EL/eTZuYLkI/pdReJt46RW6z0lk++ei5om+HeY6rKukRcnb5yO9G2
TkVZITZXbYQB99xeBv18Rp8I85aK+FCQnlicYcbVU4RM9af/GZBUX1r2Jnbxx9GA
EwvAHnIKUB7y7dOlEXNewLfVhN4a2bgmNi+mOCdjfY9xkjc509mY0UXPq1DQjsMA
TbSJQv3MQ2Fr/cGMiPqAdhFBLDNXFvZMpHqG9W2D80tF9PxuI83gBsvuIoiBnayo
vGZ9bY/PjTzkko+IfTX90W0qN4gXk3MKFRHQW+mz1m9UzE/+Y2PCDkDSWZYB9poQ
dwQXylSwW5xZ8V80INGlpLSMcTC6WWV5PkBju1rDdqBT92fbRAISjId9tF5Vb4Xv
PJACC/DzfSamCpI0Bu/TEUoDrDbRJReZXMJYFq1EcriYScYX6UBJBal9xDHT010w
Z2iS7mbpsC0WdJFA/ctY0PEtx5XV0l71+WiUKXN9Xl8DUuUEQMqNdIGy3sxi5a6A
vY7IAr6B8RfxMJ6CN+VL+LmWfexsSw6XiqdIy0mpZDSYsvQHKdsTOf49PIQNfAOL
rMiP2Pbh6lOMMl/kbeG96OxcQ5omwWdLw6czOnMveJwgqSxbZXn51REFQkyB4RU6
D2oHh95wk3CNwZ2wpl6m+zgxeDSUHuIT/hvKfBDwn8yrpSV3bqH+NA9qC6G/JE1u
Yty9l0e8Hi1XWL6Q7leyxLoeAZ4jTk9hm9qaBcycpjUMICJlDm+WZsg5WFlO1w5O
U/2z09UmP1Y/dK1bBahaHO35TIs3M1RC0WBj5Cv0hg0=
`pragma protect end_protected
