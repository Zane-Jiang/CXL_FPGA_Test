// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gEMePxXbasrbIcV4B1CJwE/cyzkCitsLTOYUXQBb09vUMGFWUYNtEgvNrOk2
M33zp7MRU81WGWZhbR9efq1YwiQsKM9LUupxXkl++Ss4jOcpyn9fcQ3p/FEG
KR0TCRu1O+nJ5EPrjlznUxcvLB8w/cMJKpWuN0YpiV674nkJ4xmOWg8/p6yD
W/+1W5ufPK+8rBmfA1vr3dV53fFifuvrTSOoZNLIlO1WqikMsjeGVomSDMKv
rpAkAXPYfFw+P1wR/LMNT/fqYcQgPhgRuWcxVO4ijgbAau4xTzzLwsb8kBQx
DZhv47tDuU3hRDpDUp6CLDMws9Jz8VaOcm3y0fvxgQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
byk0GfpK3yUbOCuk7ay5Oo1On3Wn2c3auggeQDcriI6ccmXYQ62O4UO2V4Gy
9lKuYa79z/E7ssXoneeTO9jkL70KyOwFSHVlry0ccm7bAwnhu3UN5U2p3SjC
zGHbKbYaeyIFo/w+a+mElVmp7/nthQ71O958wd0TBznLzEp+nLJ7rMlu6y6L
7+LL2Z3/yRs3soyrqLkvaQy10Y4Y9VRctGk/kDPOFSpbMl/eSojistwowiNs
GsMMY8IHkU9mDhKqV6S/s7zFmsCOUbhDYix9wlrDJWmK7uDNKO9dBEENBEGd
Rf57W296XCKL+fdh0WJfqTDL8JJ0Vd3cDByyFMpQAA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HL8C0nVyXqxjKCa8f4CSRf6W6IC7w+Zp95tz+Wtopb/ZDNZTroWxzE02vhqq
ejgWB+maN8+/R0aX6+G/uqbXiflWlisF5bUeyHUAvg2QeKum4xhwycmXlzrW
44UcvWm7pTF/RcEfIwTJjdEo31H5fvacciGcAmh0bO8zjqk0pXIv8E+AKf5X
5WwXV1lFTWALc5vj/SGtg9dTo7nAZeZwGMnMmpqJKVCJb0Ize4P+xc4BY1Mv
u/TCCFMPT/OiCG+iF+gGOASvQT9XttG9iyzD+MNP+uVvibdev/A7XhUW7J1e
rVSNZvhziip7dh9A96R1CEJuiuJGGnC8h9DWcLBwjg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cp9YmviaQxASy1mtvgBo98Edui/z+ggXEBhqAR19s15glpMQ5mUENbWdjiiU
LJF4A3y7u5aS3IxErBBgnDkq16xpjUl0KXXqEVgYhwYGZJ54xj7MHLpl8vsJ
huk3TFFT+XwJKqamix1L/ivdQqJnvTpjnY7OW9IqinZJpRnfFHc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ms6ftChb0LuBEZTeJPsf/Dm1CtSvnXxsE2ms9+E4p/gh54xhOP7/KmxXoCDk
F1vonEVnWA/KGEORdosC6FjzGlctTmbKlt/+InMZOpceADVBLFuih4w1R4D4
PKBjszWynv24Qhm1sX7kJBDQuWRm64acBCAkoqpx+KyWP4A3PfZPg51img67
XTT8lxEppncArPAECSpXkQGY30W445kSMX2j7Ivoit+LnFRHzPqgDMMwAGTz
JRnvESjqGgWHjuKLsTeTTbdfdda2aVz7WCE36aIxCqv63/pwmgaffimhqgXB
GT8aJkmCiCnGCb7kIKvW5OEIJcHO2xAupNKkdTMPkkIEkojOvi6DU4Rq/MNN
3Fnvjv1JtX8rDXxka3iIScAcor/8TjsB8pBOCrBhczGfcPI2LA3YQzViih0C
/fLsE8hkHm5QYNR83Y48M4+tpZ2BfVRYksC45Dh6Ai49tFoGb/YIyrSUEoA0
IxKRDHNIgm8Afu2me7j3bP/UX7tCgpsD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FPkiV/b5LingQTmdXq0MzO8IRAGcpqdiurb6WCxRpozcRSgV4DaUhHMJK3J1
fOBnqlnEXppoFnC5TmTirfXFyClClxOgmWAD+JbPTNv1ve1v1696OwcpvNjM
PN7ztdWyzd9/h4xeUO6bL3c3gZDcC26NjtM+Wq2B1XF6WbfwgUQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JWCVV6knDGTlGFcekfVYiyvjcoAgaz0TbdS2c5AHrhaVOdpW91revfn6a0Rb
6PT3s/6CtpJN/DgHjIVQt5Gy4NnX6AgifjgxXZVoOFIJERsjIF5IvmsnXy5b
ZWqzhaXUBDZTDDhi8hgtgeIbvB4VfmDIQwLxybJtvL2LIGwAP/A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 37072)
`pragma protect data_block
G4QRv5U8MKGA4TMDpOpymGTSh02CVHHu4OjEWrCK9vwgB9eaWsqty0/faTPk
tI5XjIBoznugKYMLVNFln9CHVuhm4cgO0k5CpYjDKD3ufIi/fuXE/758DxKJ
Fq7n/7gztGLCA0Vl5XSboR6m7NoASGWVRXGLyfOUxfVfBe+neN/oxRxBwR1N
JOYKZJhgdAXP2PhsDpFyhA6DijrnBaFCd2t6QMwmnqkdBzf7MF6C5yi+IteB
RiklSvrq3IoP3TRGm/uXxBNiA9iuxOGMNSCRj2Lef9uVwER/l6AWnn/BPsoq
vJ4zWaETpoBHz/Cx7whQlYJr5XoWm72IY6q7uRju8yzFSW0Its7I+XxXr0VP
ONJG0VtpcHxDfTlZNye+2XVKmhGXYX+qgZjoBYT+Cu21/12DoGIdItfW4Q/g
XEDAIJpZ+rKL1NS7kYPx4cgh6ewcdeGtGzJ78QhsvrFbLXaDQbBCkoBh2B2I
jpqfjaATeJOWG0PGS4QPQ+cnBYvcrmaLmXFAryh66xRmVVKF+1NPdPkDV9V/
K+N6kmmFUJTBhVFL8RsWSv6WnJOx/BMziQZAmT18YZZlrMkeUl0BxgfK+hQ9
3RfOcyU2YXo323ecDZRzxd8hyEAaxBwzztAyz4qwqFw9INwD8DX0NBpFqh0i
1qkzbGDuGjdU9ntZPYUOBAdhQbx+jlOPRb/LbKHa7P1EAwNexfIvKorj1FMF
WrSpHCnD+V9U7G5MarPWqqPVg38ssKUMAJAXcHli+1B1xbUy0VJw9c/+ehZV
NdZDAt/6LpqeNL0Uir4ayddDtrPBWuEEgwLRV/Ez10mkwlLAWQeqS74Mth4Z
LgynvNJb135jGyOjJ7c+2QpTiyb8ZzVr9GmUAnaGozpxfh0pOVQ53e7oO+b/
XMH5jwIgxPO9chqnTo1hfacw2JOdJ5bL14jki7OpKqQQYADoNc2NS3WSq8GI
V7Ne2WokS5pG9ug6NMIWBgliYeexab8ZNE3cXXtvfHNQfBj25OL21VYJXxwn
QL6jo5OQeCl7B/7O+beW9n23XJ047AYjO0Xa4FzpNr2abSt0aJPofZQ01OaN
guPahbJXBmP+VnLCMijurXEUug0fuCNIH7oeBZomVIOUthpOt7Mp8yGWZMss
SnvGX34NR3NutFhQsEd6uX/gCYxWqTgxabVTRXtbjzmNno0ljsSux2YRok5v
zfmUyO/941qU+IYLkEPueSy2ZQXPwwyz8a4Oc4WUyGtusMAu4y9crMPOniPs
p4OcKWlflI7qxcfhPoM1NQRl/zbye33c+pMGyJKsqdR91kSIAFSlMl/7dCp2
y9QIpZ9oItdbAxsdEqUFg6B1nmqcwpLV3Kp7uvnEVXJfyIDYOsS6CVGMCe1L
8mbfuoEKhLAoQy9cdGCpplFe5g3qi1cvjF9GroLxMqOQanP2Eaj9svficRPJ
2L4I/yGLtrHKL7uJbxdstTc7Pcwhlx/AAsJi+mcMH7hwH/rEHadsGqAjnzuT
Vr9dbPPcHLnejTrGZ5phwXf8Rqc9NOtRL1i4Sv+wyxGW63jBYxC6sv3yQrFl
OVNS9Tl7jsbae5IS6S4tNbkPFo/0Ck7vW6cQZ30yAkRidF0WPbg0uaxtMiNr
ZUoQW2qAAbHl81QZ3kZ34pLdrU4SMMt5szCrF6k3m7Yknc562RMQjKlpU1pO
iv3Etzz4sFrc/0XZXKvX1oN5fu5i8jzJI/68Nea5ZYJvR6cDFdHk1TFCDFWt
irmYxbKK8uTHsC2F9Na9Ye4pufZEuHxjbXF2/hvy1eUuERuBZymqiC3NKohJ
Yu2r7DuO8XcLZ6hxk0/bqeWiaDgcaLhX8M4kMJgAaeRAOhFjWWmJHhj3oak3
yYPva08vInigzq6d7R5Wxu/T3NVXRVN+9meaMZ1LtX+yvISFptqMNd1DPEHE
9u4LIj1dibQKrHpwadzLy/xp98zTuiEG20kkSQVs5Jvxc2szJT+3xYMJ2mGj
sPHSdizAralPVxkm9laZwdiEIaFGu15Cj84fJRbajKX9FClHexcL6Om1DIUe
iJ9nYbMupeWtnsqqRNUJAFceFFsDAdKNs5k3o/CR+4my97JCg9y4v3jauG0u
8GsMSnZ14INthQ2SqOVTNrsdJXsroW1YMcleJeeE6X+NlSXi4Mv/Pn+irYeK
ysBeFhxG8A+i+9/yY+ATDrRhn2tcSA+E0gFJAZodA516pkiKNaEL74EXLpnu
O6R7wTjcvPIJfeSxU4+I3+J0FonIh7TF9wCaz1ZKZWuUG05+CsFXIli1xAmD
+nQPXY3yZepy+jrBRGSK4ky/mRK05UoQDZ0QvJ0F8cM6UT4P+RMman7ennbX
gXq3JiEEyAarlqk7rSgJwQfWcKb5qEklqQxQ7USu3fuE874sk/2hxaFlVLCy
mmbgGVsOc2ModSt24IJDmUAs59nTnuqTrOA4tDZ/OBNB4kzj6kqUmR1MWcx1
OhS73kSmRkaZC/KCICn732kpzSgB6nRCaO+Dtjfez8LgDOk2n3+ZG5IwoIpG
dTITA89a09HpdYqO49m8HijjzTUuTrEWKnSpymucLqRA0rI3hNgTdZfIooLT
yX5hIAJ2iMNnBA4S4xjOcqrtp6SlrWus5I99jozXPrrPwEoPnEKPyUwQL6kT
gOKryWD3h/RZ0V1C0WKlIfMcjzmXzMNM22IqZDkRooksdGlJSPeLlna0lL5X
I00xLM2OkR3bFuzZWmdGB/vtOS/blvzQdArwsGr//i1butPC8NQ3H/A3YimZ
1lL7HxCqK6EZ5Iv9E/ojCdqYcIuIb7Kf1Lgs6DS5rxM7VhreRZreYeTDNsRF
gUHNX3ZTX6V7ZEWvfm6QHNSQBoPqGlEkvxF764lcq1EKR11+In9NSrO/reBA
Z+Gghg3zdNg3vQV5iTbgINU7oCCEdWg9bmughghSRVmPPzC22GCLRZEEK08Q
aHA8h1s02oN7ou/54W0v4D7M5Gh7+7Ak44HJ0IADQbqGplTco6hjJT2P82Qt
Fz6PLys7zYDTyK8b4L/1Pe1wyQdJDflz5Su5f3nNpRTktZ0uIG4vA7W8KP+i
KajO6IXqoM/TFHJBVdHRjfshVaaMxCEcAjxAEkSe0apxVNwwqmjOR5VaeeEW
wSuLKPu7NfIzRsy3gLQ5Q93BlJbAa8Eoj34Mtl9VjF/4bML7uq8De5ZvjEGQ
g7jkM6aOgkWZJrBn+xNQrlGk2oS8mSu4SmVTH6VlnF9Ou/HSvtHFqOXVceAt
K2FMbmmw9ToIrhEgChj34Ocqq4xENF+EJaS/NgpQ1mD2OuI941Ii8l+D5dZ5
Tq75Zymg0q0gJANDfZk5hglbIecYhLi+Hhz7qCq/JeNEnrmxywWkxGDWX44X
OLdCamWOaM0EXzJ6oSo7RkVrpFoRSgnX5IJ5NA+dUeGS5LIj9di+UYT4E7Wi
/PdswRScBhDfqah+fie5ZrkkCoEFSlGkZy4sSSAVsrVHLD/YeXsEoxnnwZuf
dX5VhcMI9EVLbXjmG1Ye1fCKbFBa/IfkZ1CL/g7EY9rhRBcUF6eAaEwpT0cw
idb+U2DoAZ1uPNOZPrXoXlcLhrQ6Sf9kF6VeliqtJFfgsP+lRwUz4Vwflsew
pysIGTwoQRrm/RoGtWVwHyg5hDfk8CYXNlODfEErV+VptDJRXihx+Ba7Ex1l
genXRvATq8GFEXcSNoiGB2ZYrJnvxM5YwzqwNHteA4Q/U3tjOolhL/nMw2KQ
+gHkJdKIdmpzwtgmsJeIROhhdrUj+GAo9D60TUanK3arZiLvs8ArgYIyYr/Q
sQzJ9fgUiHFXkpZW9pDKOhPHNe2vLAvA2yQi/oQ86+byVx3IsDfoEOru56yh
B0+hUdG0+eqzEFQLHzkl/Z4UVOKS5EXsGwYPNhKOVl/yR8kWHDe4QT8OyW6J
Eyr5hTNmZu6hTflt8voQplm3/RRszl5rIBVs29gGUU5BdtqBpidoH487McVt
aT+HF9kpqp11s91mj4ZnvnVqlkEkQ73c3jYaqv/1jIShigRxaIha/mQu4U7S
CLqtIOwdWm1d38bjfluuZA3stPY2fUldalSZuZ3VsCMDezxTLFb0644TV2sT
kjbe5/9/3OKVo2xkdhuAYUa/vebzYzVhnnCoM3I7cQlFdi7buIg2j+1BfgGQ
OsaFhF2qtqL/nfnKdvv7VEgzklaGf3o2cdWZYL4M1JbalRSIq27w+lKlGWXs
r4BiWOH59d3hl0MUitA3Dc+mG7HNoWCmt1yp7j468WOAY6MqFUWAnY95DZiT
Z8ld7ge0HCz3jmMhMuM5cKZ46RF4vf0K1bNnfwk/7RQZ/+Ipcy4lgGWuWtWU
ixj/RngRxgAB9eLT+RlFbNF0qhEq/HVwsIgblcfK2Dv3dAyatfCigzFyfxxR
hQ7GSb6W6wSk4Xawgm7F9I9zg6QGA2iMYdjlSkc4E/JK6KKwfJvnCPKcuRiG
36lyg2q7XCw+Se3O7FXQ8Z/+VxVcNfaFepR5JEw+QqTeTo3yHi5I0UDt1ujw
6AsfMCPoGHqipgmfy8VOsEFqiB6mNO4HbvLGDcTbJKDDLsInKGuSRLPzYfE1
aOfQvHWSMfn2aXs9nXTimwJZ/k8Ufo482mOhQWIDaxLWJVTD+W6SzUMzSZYe
0iMkdDrVLexKkhbJNBd6r+kDha/0Egb2PMJFioy3YBonjo6u+14RdgaYdv3e
tFtcUoOlxBU6JPEBA0vW3NyTsiu6TaY4hChzZWTHC1WVG6rq99ePSd8Kv17A
qGCvI5nSS1KvW1bmp9cMhLZnlLiK3A0fr8pb64+Tm6PCpekcaoWCl38EffnY
21trTk2ST8jpWzGDMJF8FWuXYEXn/xyTY3hChe9MEjv7aHyHeyKvfll1esRX
ZLPrSoPB3bBc6UYQO8WWyXdMNrNqCE88kB4s3yFC/QdWOmG7gcCrxzXWTR0F
wR+ZfeXEx//WY3CKwHg3hx5s9rj6hlEKNd/WtvYjhzvNd9l7MjVhKI77yssp
I97I/tV2zqsvebwgwXyJWitm8ux//L+vAvHj7KvuhAowZfatyEkDqTQh6lhf
8IO1c4MuyyIYfTwVvWOjY+V9yu/yCu21c/U3jsybzkua2091FByKbiitExN/
t1FSPVInk9n9M/y73MqqlkSMoVqaV5/KNGODr9VkwD+sTxnqGOzacUPn7YfE
dUiV1+WmY+Xg0hNIYreurTlAGKag68MjK/NCbotb1rROeJWyp4UwDWnVBF9Q
792uUv7HAWDgRQsm7mp9ZOrGaaZ+2Lf5B9u/Ygjwhbd7dTk4IFc0qf/5Pcys
HlfPU7dZ5z66QRpqwlHA5L8fbqEmcbI0DuELZmvMeFLi5JHvE16ELqsqzMWK
SSLXbf8ITytZ36JsmqOLwVKtphxec6dh9OtLXztn73sMXc5bv3OfvEBeYosG
ZiHyQ61Xiomkr2WCUy2dfOyTgw1ddPllxuxl016GKbru8Yr3+0DagzbThNYC
JM5dimF+caF+wKY+xIbEhTPEJRgAbXVTErvGCRgwIMjDwvWNl5O2EiZh+GZ3
N5zCKnZzX+yWeOKhEttWxbaOv3RqXt5GQgrtKtV6CoPOHOT8arlnVLOXeEs+
Kw2ucN3XdlSlmpitbs2mepbdcdLo0LFFdGmA4cOmy+tH+9OXKijVeWmg5SRF
VrOXzTjAqr75wR0URco8war2c8jnO2JkyoAkEcec1FhxJMK7W3VjDHAxWwnF
5L9xd8YgFKdvlL48atrMNDmj/rf+XfOW7SKdUKBDfKLC5My6WII87WiU+RtS
vxJzifV2uhFjT/Ccn666sOQ6BvmTnq2lFts72Yhr85rEnrfSThhwf63yjXhL
PwoH1wfn3ztPTFCo/cb2UtTasC8DDYRx5nUkL7UvtT5dUSFAaAyU1W8DZIkv
Kghdw2splFGHkx5IHEFfAjzZKFIn9vySKfzM2zbn5BfneGyDRqyA2XCVXUSB
dbz7CTO5xN7hr+OrZL6QTc/aA1eiZ170ts6PLeO1OO0q3QcnGmKaMMMZd0i6
HjtxprpNxTO3R7BweV/+Ziag2+Xyo4l727EHc14ogqZQtlRUf6jm52jpK1sI
ARmmEeWUEKPwTqVWae5rffUh0tnmsTPYr8Qlzw36xs02v/ZplAAmE7Ma37TQ
gw4nnm4TaHSyYBps/zxaM04u1DR+Meve3a1jb9j4NNIuz6RDrE+/C7mmZFdM
ISHFqHDjD4qRb1d9jzZ+iIwpW7MRhTsSHQweeQxBc4pGak33wy0Jk3U0H0qY
ZHC9LzlSiEjHw6XmvxAKXYbHx14ZK3bLaan/JEyN4/4OorBppq/2uJIv8D6q
7GPFkQOe9frB240KHUDKxrB9hnrZQ7c5TlUdwTCeTHs6aDIXw/hIXET9alRV
sG3NIrok57CSdrEdAG4ptMYE2NWNtCsTflalEwL8dxHmR27G/C5w1vnsr4hO
8OYg9bBGNtDf1H+IlQAQIppGuuIp76T9kvrse66JgjVqt5EyC7k5b13iqEKB
sx1hEJJLHQQh6mVCPogjXCL2fW3JK3IaMDdkr+4fvjYX35SyXvdbO+auoEaA
TCO5vAvjFlopKR1FZ8OavuKuVfOIJtRH23aM2oxBwK08wk/T4KE1tVECwGmG
ej/NG8t6QQpY1URHeVWHqWHnqKFE+7eLWvLy0DPxJGFWycAGquy76/Fe7qPa
vIzM+gBUq53pWc8mpW0gd9vwkKM75Yl1RD0Nr6StEbMdMFFsGRDt+mipGQzO
uRzR4gAylGHgLrqSGKeVMcNHfQoiEgcMby5QQVMxSnjBGZDmR/CE5dJwixGQ
sp8gHPKRlBO3CK8OoTqDLwip8PMR8XKU3yWQEoys1IlAfgP7Qkd9wPVDU2se
tVYuSayJgjRRUVJzclRAO4aw6JnTq65eZE32Uc7auZwSpsGzEN4wX9E/1DZf
TKkO7CUM5INundfEReEUA1/vW6gF9h6ACqgKateIsHdxGh5f2c3213MTFz8S
YHmlZwaAsmQejXsAs8EVL7S6xLWmDcjsseT/69kHU1Og5e4+biCFSmQfV6R5
Sr4yCj4UdVqdg1bDmjDoA8Z4GrmAx0EwXPHktuIx6+pMzVF6PhJSL7b5S3Up
B7m1A3LYDnXWF7DeCYOLnc7CsZSH7j/Oj+fJX4gGHZmwSPWnK2b7XQ6WC9hX
K9NR4eLDthZ858FaE0pJ7kfTPB2p9malo07+SnL1mOH6rBAzD/AJiJtzcyn4
0HEbQ4tqywqFxcyoM/hgRA3m0FGzbkr3aRzcamLRJrSE4Vqkk46YLNuOu1jS
dZ0dyyDa2Lu4PGTYHNdFVgLczECMnrx2fTVzlXs3l3zZXIuwpVXaPHhFZe99
0EX23F3kwaN/MlHluhQQUTTAuNVSPbx3WKz5QMyysQ+VPRX/FB778M1HwGxU
QSDdKSH86RL9orzE9yiXT8GS36DMcHxyGAz254bCa0jmnlDc32RLe5iEoPVv
kFMXOx2HhcxxHbU9DhvdbgNfOkkol72YVF+uIs9tuKxAZsecfW42acH79D7+
SRDSDPS1xe8YijSAh2VBWMaCNrj2foWm/H8ldtGx0QPa3M1EndcJNAUi0rWt
YkLZMt1xU72mt7JZswX71HalzR2vDOGznTcCrsbORm6vXaHiPbK1wDbG2rGc
ArNziaoid2ThI8YgPw8YvVuzm7yTHBOt/TpFk0Ao/ovK3cUaN9QgE2gjQ3JD
xT56IROugHupeoLGYxnU6IPQqarcZChGWthYkk47ITq20vuWUcXhMeTeetrM
fwl0W+M0imyjMfy7I1MqULtWSRb1gPD+42nXhvMLnWqU18I4TZGA4Tiiyump
iMg6fOkYJEBfEZWXERzalcnbngHbN1a7IrVuf76JTcxNGnnjU8+Bk0KjHXDF
lIOHLKFSwa47cR+whzb0655O9++WPgivQAsuTxIjBGnb6Kc58h8FgeN8ZE8P
p9uaNBYSAEv2BhO+Fr3AuYqiRl0kA2pYuEalMLF/sGx6spgCGe7opHSaS9pd
+OOY7SdP3dtJL6dA4hp/yptvplB+p2nwwpefeP8C7MquG3Y9RShtWHsD6DkJ
8V/jbmQe/9ttRXx6HBPCRno7hdiJitYNYOY0dEV4CjvdXJCTnM9uuuw/ir+h
e1qzTkRrSw85ypOQ6zEmbOEUL1tvdNMYBwqoQUc7JbuCx/VNTKD7SYH4D44q
YttCrp2EZdp4NRUZvt1e+26b6oWPvSHiCTQKe6qmQdkxLkCI4fjPrBCb3P9c
HWHE0ffMQV7goC4asS+26R9LYsLCL1NfB/YDPAn3WbvSRMGzZmmB/Wt1e/nM
l9+hucQPerkzDaxn6hL5dFZm8EZ6VEjzDqkcCp9YGYuzBEtIsGbIHFl9pZoV
xYo7S8fZbrRu2xf72bzQRvS3xVTGi0LVtJBK9HmhsLXiuMJbv59t4bCaczuw
WvDVN4UztJt0lqEGflDPqgKKpylGqVLBGXQU2GFWXWLS1ljonJQPhTwd0oHm
mnhjQ+Yg++fur6OdKE4+QoQvhGS52p1YGIZfO1Nl1WTcFzkPikNgCWtO6v8R
158p/Axijrhz1PTbGxiz4QEZCaq9qp0dmzniSl7f5/tk/A0gyX2DBVdiC+VM
v9DCYvDIqXtyxKlUs57wiROLZCTmmCRSy72K1YaIaUE5Qv8yAEbCbi6Ptv/p
w+2hn/TdifNd+lLrklglhss81cVmrxkCJXZ0/27KcklrbSwuo31ezukTbBYF
9w+z5g73znzF5eHWzL0+9ZMtr9FaEvlcbOSwZlE0fp+du5orpLVAac9N0qAw
pTJeyeNJBf0vkcZQFB1fJK6VFc21Pg71yoEzgKApcCC+Z3jLr0Ms22qbTJlM
qyVP+vZTxb45ie1TTusAlB1jhnpp/ddvcgMhoBQfenYtx2AlNYEbXMN3JWNz
Tu6qQstgvtVU8bzeohou+syiRQWg8pcnBAaLkXCmRBsoiZF/hoBkx62BcGjN
fCzdlinmkbsuJ8Z/abNEh1j+bA5YIYIc4rSAzhIUMoW9FJn/yLGPoQpQ26Hy
i+3ExYFOF+w71GYnAS3GV5+IknTc21BfXuJKzX1/8lZP8iqIdOvsv5jnPcv2
PiRrmTQR20udjTM4UFPlfi5fQy7K/IcI/HWt5DtREl0LSgFOkweTAFNHkpkf
w7GmWePQfRK4bRbIMj5c3CA+CAefBeHAeZHXCFS89iC4so/xixBTY93ewtut
dilYcxBBQFYu/YmAJ7CJ5v2RPMKq7jBKD0XtkfFxP/xkbnRu3u4J48RWkdaa
DZTcJ74U6Pym/qgfOeW09y0eaUSe8mgu/aMj1h5rKzHJKv4Je6SJc1KPr+xn
HdPS+tYqaxIwQ/hjMORq1ixtqd2Sute7P5cuFk+Il6UNYQt+6jP2D2r6VSQN
BnI+0Z4towHY/IGRRBtRmASKEAo303iAdDeYXnxx44O6N1BQRpHhj9PWgimI
mBgqw6bTHKaCVqRY+tDhqUIA7jS7rMIXjl5XqXbV73JzhcpcTlvqhFDHPd9i
xbpvPGjDENnbyfnyv8YF9EFE0/Tdo+HAgr/1b6YfQP+lhbn4ZZSgN4M2ANIk
pxsysH2tHme+uuidpFQqHsT7beef+f9PnvtH25/3d7VOWN9njIO0j24KdhAq
akeOxz2hapRfKRsE/qi8GNFMuvcQ9J3VbTHLVhr4M2jtfmLKqO39lpd8p8Lm
ucj6xm8mobDt79ZRsOmphZiRkUa8WV9/pO+Oh3ybGcMEg2hvYVzQ2xfS76fg
XE4BwwxXUZhfank0X1EUf3CTaSHLAGIXGv75OjrwKmg5jaQrUbyDFsHN+eQ7
MWDbzHaIQts2tUfJSFhhyHJpEMaeJOlMhdxS93TD21F5cVieQCjzs854dYrj
28xxH91I7UjDhAaYLI80X1K1sr+cU1UZ+5lezDHlV33y2ZArD2tlPVD2nlZA
NzKWM6dCUEXdwc5WuihPhiyewqZoKvQuk9muyHPzc6mYbiBDO8kLjRaKTrOs
83iY8hP8E9oAIBdbj/Pp55O5nGhLMjm+xRun6nHDg0tPn9TcXE92wSp16Z+N
bbRd/PUNpUq1H3pfDeLW8+hG+XH6g//Ry0ywn8VczwwgXbpDhyNbHfL6MX5C
/UtEFF/zxe0iZoZrSHFDuJFIgEEs+SxGboAsUisJajUMMjjR6JVEpzRRCXjk
uE2dGFWZ2RLgR5k7LjI8Edw87BNRP/xvS+1oqTH3CEkLAQvlUAj23qE1p+TE
9AX11srfGKsxCD9AZP42qK++nKyCvu67MJeI9mt1OOdmPTRpP1OsTEQdORHl
KFn/cXuQ9g1GP5TA54ECSzCqgAqqQ1vhjHQyNe5lO5LBbT8btPjKOVfYtqoT
98Qf5TVngBLfffYAAv/HK3zVmREiCTV4xnv7EqOZ5wwk8+BHsF0hHkkDQqVk
uQzyug3QqERecX/Ge1KN75+l4xWpUZxjdrOZ1WDeXL21MLgBjlxQRJcYZOkU
Tc4T5ff1N16cHsyBFpyB0ECM8MshV37hTF4tbygHgR289iDLOUiMGkfqT6RK
bxUYLgQxqrgBVxAwLkiK9IusT67kapA0Xt6AOzjfHZFJdTzFlBLDYjYPm96g
rYdr478V0AO4rKxDM+ddm4zFbqG8RKmY2gjf9OsQsG2gJJks6+ZNBpdL9yGb
YwmPXttHEQOppkyBN6KOHpb8HNY+1x4kiZb7gAbug2AlExraYBVwxW8YaCIZ
lHITikwLEROPoUMTbSHz0O6uhHOgacr1VK0rXa8vJ4BA7NaCJch5tXl08Fzi
hQx4Yk6BgzcxifNRl8bYGotOcR8FBmcxxHvz3lWtZAtL+jmqZiFDBJR7zqnB
FZblJo2L5Ez3GW5C0kxqAJ4YpXBq3futay42fwvE7NqBSelHVYZJvnxHmaES
vdidlMrTsZ/NRmT4VVrqdjAg6QwasQFvOkLR8oQ14DJqU44DSIFB2pwsdFjE
QZbD4yLPkA8BHnkvaQHdLlDW4Bu3p9NVf2e6BUgH8VkpY5lq4M8P0om5qhkb
5NvasTivVw5i75dTASd9SIgwmpJWvZbeMeWe3TYISlDvnbSDUonazkHWJplH
mfmA5bFcSL7cNDkgbyWfKUJY01tsYrJNpF3JYgKFDSSwkawYGBciGJ5+qvfB
8XcmDaoGlKOgBQR8DNETn4JQnEGcVk4PzCaQvQzWWqM8TvPUVB5zQSXCOzgA
RBe56P26zJinuEluPHaxtO0Vb9EX4idNdgEO/6OZDHVjxbkQz7K/LY+MsBuI
Awl/5L536N1ECdlGLzGxVizXzzTczktF4hg5rg1pd5JZFjoq7DH0cYD+CFgN
lNGoAjFi3mAuMo1kGZvnuUHsarPHjcFD1Zb5YHEOyRntAZ5XHDoAceO3ADux
I0jeUn1tCeSmoCfUpYmjlrSaLapT/sYbEKqnxBUmJ2m2iFHoAUNepdtPrEB8
jOjBOpUiMFqUfuGrX1P463+OW39MpScaBmNhDqrSyk3cE+Io4wrCUhxbjLU7
c295ckwbdsrkesV89VIfpJfDixFKWWgdlpN2/OYfHf8AOqBvtNvrqZFp9+uU
p9c1UDHWbBRdzDw2oOIBvKLtdu3UnvzF3iBDu/YkmrKh+CVmvkFizpAkT3Yc
A+BScJ+NlkaE5ipbRqqGvx0jB+db9gRDX8fORlSFmd67yjdn2CNVf41cPKzj
aUUJtgmkrho+0qaiZaaIINnh4DpqENh331AWjBqAD1UbfkdaHcP4pUIomN6O
Mm1sOJwtlIRNG2HkKpW77HKEuPyKXPZ8DhOGNWG8sc/z9Di5oEPAe+RuRjXl
2sICBEByH4C/Ntmzev1zX1x9V0AdVPzNDivzUY0ZBVOURtDfZZQAqk7kJwNZ
oWVCj+a6VK1CrlLBH1hASqX0FnGl9W/CQLRyNpOrcundSughRERZnlQ5tQty
3/yzahZTfQ8tV2yGveaINIHgusIYSqxXT2m97DgpfZ22PHF+HXA1Pwv/+U6B
5os+dK+EwMXDIHe7WEwcNZSWw3N47P/KiS7/NW7XuZjs+qy2xJGmdHEEtiG4
WCAmjd4QPoQePATx+s5E0AVDl47i1VsanUrgvp0ozj6SDjZfyu8CrDr9EzAp
jxek1hw7SqRw9VF75i5Hykv3YjMF6jm9tpPKzcwxnxX9bAtCAe87YRjyZuGG
c5UXKGrWUIPj/OuotH33HJ20gRegVmYa9McJ2xRyuNo0MPOS+1kvGAxDa8rW
8A5IL515yKmWXij/l9hpfQJRYVgKXQUCjFvyhHCQhviDG/+c3O4emuCY1xEG
P1dhfzCJfD+UU6+dRISih7APDlBCMNfVPqwWuzPhLzVkBDORkHmyAuep8iwe
C8M/aynkEFwS/1j0iDXq3vd9JUntLHYcV5Kd0wKf2MyWT8qQ7gIQ0SR5fN5N
b7wcoz59yywqFiHI6Yr6cSsHNA/WjXvqHw2i3qVStyXxIgrS076w4Rrc3wUF
BfQZ2GTQHVV7cbtpYlnXFsEfQZU65bz+RVnYaPU1jNcgVVNBVLfTOJRN1B/v
VJgMbLqn2lp8WDlgZdhLCREi4nUrmFypQzAudWIt1GDLTLgkhPpTf7gl8Van
nsfeEnFi5QXmRonYMjc2hl3KDGvMY4rMv+yywaVzKCzc9BwYBBXHEN/82sEG
26lcq5lJZvsW6zZK1NH2MxhhaJWuhJiz5mCEsEkSBENXv9SbtMdvFAeka/xt
TsFHsp946W60rKjTvyit1N3g+U++eGCOkAn1hq8if9QUNbTX+2Sx1C23pOnC
7vnhgw41CVQfDnthCc7ZTHXylW6Ytbm6vCeeUviw9UPrT2om8e0UmeKBigMA
ELCV4nhE3S81GZUEqiZR9OZIONL6nBbKnKhWcvT/9hbUH+kXpngC8O/rHzud
vS9IW7vuA+woY9h1g6sJGXwSdOySAeUbqi36tQtlUgS1Xv0dglhwKNOllz8K
6N4MX4sHuSFiEOO2xlhPwQkFpr48nW1CjDpOB3QY/gpMdYbgrHPjB9NP3tmH
JjvjSGkU3J4xb9fIBJHXGjW926JqB7Kj4sdx07SNFJnzq4kdPkjeGz3oeGb5
sPTLcrs6TfX7LcsaULoHJriV3cS7uinGpr2Jfag/XEcE/Jcli2+C1LQNrPXz
U/JqwN8wE0XbOE78zdMfOfwBn9YtyD3ezfODcnXdYZHkiazw3hu8HI7FtEj7
XIWXcMzv206Cq6dQ/+V8F8bLnFHU4cwwyHJMCvIt8qt2aiv9s2rDzxlA6il/
WGEZmpTSBT88rtCaoRglU8bahBQ6s9xOd9lKCf8BFpY0bI3QZx8IKyo1NF5J
5CpuPEvecJIIJgLN8Ag0kxbJUk/e6kv4qV+adLjFwBZM+NwalGpicXAr03FR
6OFFhrgAF7Iw5MUnBjQ0KiNzVEie7lneEnJ+m7aAGo3HONAH3Z1wslpxbzV9
r3ArFEX7vPPAKjfGrVe2cWCRpLyN7gVDNoJ1DRS+c33onRkDc0GBotr8RFyx
bL1OObnHu0PuWiKQUxAKqJQGNac31p+xqyBiJoF69snHyM7RhxB9taFNquxq
guy8YTZbf4FmSaa49cz5D11X4mW8/c/A2F6AW8axewVpyGq4ZVcVP+AvUFPU
1knCeK0DYu+MhwZ1vuLxq8SsvoJ4Ge6m1qRqD1Oss+QNd87UZozZgyamZB7Q
iqdBMtHU2GHQCTAkm0nRCLRlci7LyL6TgW/mZB+UwxjMSX5Z3qOidkrlj2eR
ueUhfQIPKYSALy8NS5yVFpnogBlgUn9k1YYk5eLr3ECj0+c41PoOB4K6IfdB
zSvWYpJz5x5FYLfefzaTLzEgCZ8o8kGXZ2qe0Z+s3rdKDkteHlL+rsu+QR/l
870KOLAzCFEQTb5c26ypYp3nbSu4wV7T5wckzVx+LFYxiCV8K8k9UgIK2+8E
2h+sO2hS107AazU/g7MXDbWTVrWnnG0H6PToKi4PncCbprcz158tY2KnhqZh
qo5g+gQnMHupHEackIvy3E5nKXWV0DPrmMdIhCkOk5aXR/BKMJKUrWyun07F
txqumtZKlpHOaMBsyVZebhcStpL8rEEgnp7wCvaBMJLQh0Lq5zGNy+ny9oqj
YZ7x+QFD7Iu+OkShMk/bU60JPwh4wxtqSSwYxAsUXg1TtEkC1qvdSxY5qCVr
tF0Vogyuf6DgHe+YbT0kH2IDRSLx7+qiJko6ccFrABxBdUICKlNndkc1S2j4
y5I1sBohSn+kxHEjFHaOlRpywFEbHmpzvKTrOhSrhe8hyoYsQTWu+PcBWWVM
srS/f1T9ecpPEQRWo4wHMeF0+rDAB/JdUmhoswgC4wRQ3h38gPnoHQLfaFZW
hcdFTfFzO1XWqEe0kCXnThDsdrP8WzW8Kl8f4gMIxY75+b8ijZ4EB8bd8SlI
jlEe6SKYBfHTzg/xZvqJfszIbYM0YYOhQOqZYf7nmtcjhWXjsuf9BnCwuWGf
vCqR2dWlg4Edeb+8WGpapCfrJfTm6Ic5AZNJ57DIF3CoXpnMJsmMjWZeTo3L
RwX/HM/IIbgFf0aTCv+InG6e09W6a9NuT6h9AmKZQ6zb7I4m6fkHICoZZXCg
7JcECH/CkVTg1LAOleUv2rNExisEaZ1AelIRHNHwwXlzy1S6D3fwE5q6VevX
yqkGtJmytmKFOwtaKUcc+jSJe8lEA4LI0h0UFdVlO/1ez3w0MsomCSiZhkYU
Goy3jR6RCmvH1ZX/gYnphO2XFqDL5Fe/MUden+Ji1qYpIvJ3kxXsparPVPm/
nvQqa2XKuogDOww5vnXhuzM/d3SZGjjzxSnFJI/jj024OJ3H0tbs4OHDtmk1
TmUrv9xBYZjtdVRyo1KtLDpviMw07+iiVtGgD61axkAMJ+olYW8OBVf4aK+C
Jjelp7O3l55wUZnKiBzjTR+oOoxuNbZiqP4nOhBpIDpGyvm6LbZAcEJqGkfo
tW5uDVcIarW9nTLVVORnBf1WnaoExhf70xrgjFQ7J1QKkN8AWSsK+u1WoaI5
Fs4lalZxx0QEDiDnZHsUqXtEYSgNf9Bi+azM6RxSj8jihOBGN9sg05LPSYwZ
MZVOIQtUh2lVWW5PwpxuXBUZoooAxGZ+UPyxiZ4tzAncgDUFVgIGlz/J7RXV
p38gJePeFctP3YkLJgl8S3BpQw+xAVd8PYfl4xGIZ2CcFfIN3wO1IaDITs94
mgJq9HyrDmQiIFB5CktSZOAlK1NKEUgqfNk93VVwlWY0Wx+Wi9UNZjYGPEIO
FAK5WhN4vFLr5wQTl+U6GPwzhxAQhz8SHAG4ismaeEBA6ve9FN6wWx8odN7+
xNSQn6mCnHQC8tfLO6cg/AvuJV0kJKAgd+Vz1sU7mdI1JD3DXBP81H/aSqng
HI34SuKyis+bAz5MefaVRKxCHnij22rvYcLwo0kqUpYVgSe97N2uLOkk/8xl
OLWJMQMXeb/TA4CNuSghozHGaN8YnoQa8z9Zosor62REmoO06UAkWkaN8Kb8
oHJ92LHOrHBtqEmUm2f/ccRDnRpoZjFI9hHOy3nIytEsV5Nv3pXyodBTMl2S
G8vK0eSYTGBj265Pq9k0gRRhU2oiK2wtFOas1PumITD4J/ypHNsSir8MlgRW
HI3ouzUOPxzPgHlnNFhwiYKDBilSjF4PEA/HevgRLjGvj8A8p57feeCSCohe
h+7uporWJhuR4i+fjouwrGnGCVoiVGvnyBY8LU6FKhgXCWCPamCk0FH8DHoh
2aW4wPdbB6adXuLchLz8Y3U9tyzdzS+j8VFVAEE29WmT4JGTx2kXwZl1xwDr
vcixGQ1l1Y3r81CUGJ1Hto6KiRUdtHBTXucYyxEVwBIpJAZKRW0wEnIe2tz6
m8fOugluaL44mx48T1x6t2FVNpCa+uQgpo8qfVsUv87yLd3Y5my2BLaiTy0z
CM7Aq33+zQzkqymLR2cw1mlfHVDVqztaaVA6kdyN6bcCE7pvGaMpwF4tJd5Y
5jxTY9xYKGn6wPdrk0vKPFPFd7jZEl6xQk401ozgon+gdBFIdB5QVbeGg0jo
8AUCEDCEIJuhTnQcANGrCvS90QVq6prGZPSQUUlByogiJrqzmXx4wmvpFDlF
6MG+KTXrusO1ODOfNyjEJZMjswno5yB6b0IDZgS38MGrOyDco5TvEX9urTPy
cQJiS11dee2qOkWtU80jkf+05MtF94ZMQVoJ6LZ9kVoM+1Pjq76tuyxCuc44
HoTO2msZuJPi1sre58bhcL5xq/0/xjq4ehxNsZPemESZTFQ0qRHsG3n5Wytw
nwtWrRk+CStTfTSdl8R8QgD41pdnc67NswhaZ8WXkut/OowxKclapLf8e7oZ
xYMnff2c8jOMlTV4xv1LZi7CKneinlpNxGjysBvdW9Nqns10DtXHYGHT7SI3
omuqEiSfktkXMSqTGncoRmKjq9yNL0fPTbPkhDOR98fcPjWGswefHKN8GJk6
XYNtLrD3oqH0xadH55r3XZgZm1WIJZqOG0SaUn4OsMYtwzaH0TqgwOlulEP8
s+aYGRelRGH6K07fXZaAFD9+oY79snBVopn+cGyGNc7rp0XQhcJa+DEXevta
mb+Ou7qy/TMmWxZTZWI4g+EXmeJuCeMg6lQcp4ra/aAWIPd6rrRjvHWIBIBP
RncGMGd3BkicveDfeHhqQIVcwYJEFxE+tLjDpYcfmW0lpyU4iTZ7AsAbonGg
HzPGHaSkqM4GPP24lN/kzVvX+c0/cMUkOrrzsaMV9pxKl35ORIuuj6GK6D4G
nOQ2bhCzqaKH8dXanFM2Sa9z2Z/ohZQh8ZFGDeob/ffZ84CnbwnvkuPWohYy
96eTprKZtsKa/Gl1g5N5CkMwgEMQYcG0NObNoFp7v8rSR5QHnJgSp768920m
8fE8G+6hagQz5QsmBNuG+1kHr8XGo7NqLOsAi4fg2zhu7gyQM/8yAVnXzjUP
1ZMmTmw81H7C2grRRksojrPuw4mGkg7Z9ElURP1lQyTEUT3DxRQqf7QX9GmR
JWBRjylx+szOLfST91C6BrN3zG8mgdyzujNRgw0tGivshYKokyOxsUDV74en
6DWY9/Rhvi+b+WRqZXemoY1B+tHvrgzavz6Z5aoZ1lhnvmJ3rtKiW30qtY6H
XlVY/pg7RSKK9sdZ20nksmIRRISQes4vbcDKJ6s0VLlPdrSHAXCYqalmt7Yi
HQT35vinRnyE7gKXtoSb+oQ1tm+KaHiY2/VewGBD92LramLu1/W+Ej4VkpxJ
qaKlILOnMNmYKB9wEqgfMvqt9I+MXU1cva8DiFmYV+9dfSF5NBOwnkHnkSOp
fn5zx6AIHosJyBpmwSNCXHlRhwnWN9iWm/61Qclw/TkEvg6564iBct6oy+6a
3+QcvrHbu5s2VPjNzK2XlOtT+Vbm623DWIZN+AnzTUg2D1x05C7jCbgGZC6H
PusRteM2u2rJ3l6kQf0AncRT32XCirFIwEgElT7w7MjNKRP3o0KE/zgASyHG
Tl7hkd8tg6ewpQEpS771/b+VI+dOdmo8VEzZtWHR8WzDP9RZ+QIMnOp8IVEG
uqReJO2QRSV4aQ5IQrWblS4wDZ9lTh0FwSyWCY3rWgGCTKs4B3HK7DJF0mEp
9ecvnYiTydD8PMXSzY8k4B9348XiC1qteQAXRxeJQy9XDQK6Bha6Ej6PXtUk
cCIRRSE7NNs5XnFZLWRuLYax7E9QRXme3DY1k67Vjpq+rxQ469WJaN1ABHA8
BQpKvDHQWHmG6olScZxOISe9DqDaUq29mRnsPgfLHBSDCk3jWxLTJoPANH+3
r1QPZ5wFzx/iUmIGd05hqoe+n3+beEHvvOx23rvVBuyLyZhAWl8uk8yaAh85
OwRCT7Ti4CYuDyEdjk9uLB9kO5EjhHSnqqM4Re2VHcm7KrVF8i03GQmFsx8P
g4DeC/kktuvy7nTtPYfJkCcaq9bRr2TDk28ha/b3cOD88QMcrou4HBXZK4/C
b7pBibpmQ2jUIvohSAtR9khjTUOKm3rXRrtVL+HyYzRmvWMjjvlE6thZm+XJ
m5zDz2/dNyU/dkVCVAGLND4EpGYRgXFIchIyK+XR+X0/N4eLiqlZDnRw9OSM
WxCAn/WfV3g1TkkM7n7sUI5LdJZHmYdGRp6t8MahxKI6HVSTGL79KvPkN9Ua
2I/oHIbMSdPB6EAWOL0mO1gQoy0A258o7OnVgwwO4Grc0tPctfNq0Us5916x
6K5zBgy5G/0bwt9SkeNwI25xdBSdIl23t5X9AtsDEQ+P+YHlpppiNcaeDxbG
OzumdjlicRlH02i9pRuQ3bb3EkCs9TQVAZsaUc32HHfKtJDMVTD8GR/uqhnL
K/JdNaBpLAj4oledQFASe928LMk64/K7B+pd3wxFOYmqOBjYPK2BPdXTTSuu
Xw3V/Y2hyKs6ft2ilXwGz2N+JFLZDTOazYc/yAYTnKz7/BUUFgQ92+sMNpKG
5ZkowOgtCjt/DT8+iDF+aQDKnyxjAxajokgh+JYJo9ksV5nM7ChHIGeeRrc9
Aw1santrSl5Sho38ZGiC338sZkOoDT8PmPYOCrL4+F1Nq+vA71Lsc5/yk/S3
v5tAp3iPtY0Re1AgP345vbOqSeOeiNzQlFOZmFAs/0ZogLrDnZsRQSxmWBEC
Fm74dgZ9ChqPBC+qy6S00xDvMr3NJc1rz+DEkG/2+OsXe9/guHpipAV6tDPf
l7gCKXA8fz1lGmaaFVnDQfXaA0sqqO+n+M6UA9Zr8FnK4mVxd2tqvus/0gz8
1MBwc8BEY+unZvEFW4k85qx9Nxb4s55E2EeRpaLh1eL7TZrGfcMXk6CIpMzs
dFSiiGQWyhSrMJRKiTSuH05oBRse/FXovmIQIZ7TJ8DE+p6tfqmfyS5n1U5X
k1qqh4ZRi4yTR9lVCc2jIxOfITpMJfuUFk5unlieiU/BOFxHNKgOUK92Ofki
f6VSX8RwXWTm3vUvjE5LYajbD6Xli07u9C3j6L4Pe6lMgfNKzVvt9mBCsLmk
dq3ALOUqMcun4Dfxoy8s6OllU2rI6Ec+NE0R2AxqRJI4yD3cjlxXEjCfZmIO
atmfLuEujG5n+yBs1bqiKluDEN2UHkM2hLs+HyGgpWZKIlR74NdB/9Sk0nPs
I8ZG4SIPMC02+8SkEOL9YS0I3vS9S/BVWxBtg/XXbyrjtCtjBkTOI7wx4AzV
HuiqzANei8fWaT67k9HnjjUbcSrXn6Nnu8p+BHfFkX5pGQUdPRLdfwiDs4Rf
z6AhfrpWu7kTrtspwswE/iPprmx9C4TfN3xeDJ4gcGFEM6tTjZdIzItEuEHD
/UFw9AtSAaY/GjlnqJ3Bl9lIv1DeyDPcvsanrQYnCwXbZ/SjvVZwoi1EfWhV
HqMavYrHGgqJ0xkO0UXC0IAiAmhZh+2Q4DrDZ7O+2gruTFIHnXEBnjscsuB2
cE+cjoaB18WxzrysnT866fLL9wTW5jIB+qg9pDzmrGnk+qQ8YqUo9ZyyQ64W
FzBEQIWdZNZEYSAp4qwHbijwAJV2XM7/nRr3XlRUHZmu46LSaWbCDl2dXgWn
95o5QEpPlwJAc8dmxbX8fICdJgywG2UBx8wu0h4/RBN63ermoo+0Jb/zbdzs
IZIdrTf/N9BR2pscgRJ9Ima3hf7bmCRL7+m4z5c06gAZ0XcmTu+4ak2Fj1lB
FDtNewJsB/EdKnsPefkVV35FeoFmrNbmGlUlFrbMz1TsujeCA5G+fygxf3j3
zSC5KlsxETnNSMZfa8cLOBAlALtsGoR1rbdPQG2zVxRz+0IAk/8Ja7m6REWu
AC0xX/dv/3MHCu4gYIojt/2dFSqaOhFlIs8hr7TtfEYRL3XAjKHDtX7CGlxC
kiAkHW0fYOpL0Jr9NRtHq4Cbcc/PjyJN9zHkew0kZdIsAT1X9Hhqkpv7UduN
eBwJ8VawR1ACN6MgSS5gZAGWXqNg/BgHLeuMR2MH5TrCCAyvMOJRyHFplnl4
4KCqFz6JtRTZ7Rla/+mJu0Su0U7oagYeFPn6+zzFu8N2YrYvL4ioQba8vVIR
u3ooKwRCL73umNhjeBDbx6//MAMVNRtwlHMN/yK9ubIBkYa/Am1+CLFA6w1O
qiXYBRc8LEf3nsosLnJzyzhv25sSRLv4belpYD2e3La1NU1rj3MuZdi8qg43
AHs4s3nl/I3xf5dJ+P3zw+smOjrvYohCbODs032kMC4QoYr4TZW/Tw8Rf7Z/
hEJZmq5HpO0nxwWln5p4qltlndmWlbsVxB7hpXQNOkuBOPO/9P8kDDRGkony
YDK+rePEm7VmUI87c4UQ6qQe+PfcPSsR94Qbsrxq/MsVQ1eiDW83rvzxaqmT
qQmxpoa2urtlF3RibQ7K0VXyt6Ixozkv0prUz0Ny7oDGA5B1GePsK/0NMn/c
vvRv26DHIoHUdD1G5ngAmSPWpvgSLQ8eLjGBAZTkClN+c9PIyUGU5PLV5faz
FtmLR6Dww2oqC77X2O7BFwly9D8wTTBk3B+hvcbX1cgStfyUVqIUDpirRkGh
CEuux+1azLxj4dBnpBWWtTha6b8KNQgLvKWDOY1anhTk4N0hbfDouSAF55fk
T/pDigeZDDxkA6tWW80QSOsXZRd7icQ6E9L2PB7DJVnwSKFn6/B2iqef7fA4
KoJB8MaxLkNC3FKE5X/3XgQxWBz5iPadT7H7lrf/rw2H+98ImgVy2GdOegoF
GX3pJBzOy4/LPhTDZGgvVdj5DVfCrAhdLy+Ezt3y+ICJT/ubO2gw/P5kiZSB
o4yToDHc1cDyliwx0F3VmRAnDF4sC9BB8LnUFPLsdc0sRdSptAF11mIfDVSc
7Em/bJEOhzbJ9Iq38wvfU1VVQkM8qk8aWT5Bh7Hh3qPyCEKLSNUs28zXpiYI
oih/T8F3ihmQbUyPz+Eh3q8PkRF4w3mOFjnPTHkC3TReGGL4+KjnKnd9LSvp
XR6GqjlA5X0MO3ItMY9MyFLUCCMd4cXEhNo7qNMrX0Uyw3IKVGdAK6sonMjd
B+d6E/OHMgrRVGuKH5JW7hgJi7q4EaZsU0spFNorK/vJQCqWr7iBqGJxeDWC
Q8ZgFigLgqAvLa7WDHNAN21DvUtb3ZKih/O68P4mOv5hOrd413xtG/SRUdOk
PozFi8czKJkRwDv73EQ6ng3UZP/MsZ6bjToMy0ahckXZ+SWpGZvuN9jMOaG7
FLdv4dseslTz76aotHgIR3JHuxgtM/7Oi5sCK5NOZsKrfYqVeR+7ntA7ryeD
FlPoRpwTfAVKzZuGRM3rGrhPQN+MmwSd+E3k89FS0fgf/Wix6zxtTQKePeew
5TLYCI+hFkKuFj7yJZrStYZveflyazuAFTmVuui26W5ywCuLqkkDludJhixN
y4tcTciN/HfrkQ8e5TVD/Evc+1+5GZgCMzDSqEJr6gNSQdU7AMzUdNxNk2WX
nZtyeL4ztSzMoAlyXicEJal05KGwPmF4Dkbvmp6uB8h4PSdsu3a73ogbbnA2
V9/PpD84sCCtARTnE7B9jTCscTOZYBB7pn985CztQX6OulFTumv+36uVHu3p
+0x5QL58qmQ5cl+hSn5ZtHgZzqtAbna7wUGzRAXjrBs0fsufYLbOygw4M/1B
wc7a+xM9rRSMgOQbeUStMkC5heuzNtcdliWlghbqzoCruFFvofxaueH62FDM
oZuCkHb6c1UgUrLN56/+5Z+VeXnYsp5zb3C+w3rBgN2B7rISnTwgx0FO8K5E
yrKsDarxMS03NKG0dcuK19rGZg9sWo5wupfXzqANfFTLPYYJPvI6OAo+6kY5
2wDFsmi6hEXGVU2Yhiffe5Eq5P3WUiUbhZ9gzOrR0DGIzT2bMz4X10xeOaKh
6D5nRxXRY8HsC7bELw+fv+/gKYqZDGnD65UswVAcYbNuoctKBSrm0vHOgaWN
evGy4WMy5sSOkPT8riN0uCqfKmSsilxq8H7VEjlnFHApzJSykxlWXpS1IHD3
kKuOFM1vJXXhB208n1FSTnzjIIWVqIbeUHr3AYTuT7m4xnZVb4JDgriV3bL/
q1Uyw6YPzszgbST/pJ1ph2BLm8W3NS5nBdpRn5QIcI/4etqLmbG8hVAqHNvR
gvV6MhJTmI13gt4KqTkQGnCWwy+wLY2aR/cn4bHglS76jFsYChAxabaa33/p
Exv+5hzWBPTr238VGmWDcocV1AGxOQ4w18K6YSchQTSrt9mYY5Veesqws04G
aKaZ426H9G34QMiwumyGoeXrGUQ1yoo/iNQt5lwSRMCnuKBeJANwTEM3LCia
jOX45OlVR05cmPyFpB6waTIgDc5uVLnxsN6mkEN3Ug3E1sGeOv9xaIw4/tVP
3qnrYOn8MCxkFl7E/bYvwQlFpoIdm3KbBSFD+cjDjEhyNLrsFsMgOGAMBjb7
KEGhvV+jRlGH7YsUa9riNreu3nWTQ4fA/Edu2F/qiS1YnyxZNu8pxXNJdVYC
PVfWJAf4QRtQUqd3HVV5ZPt+0noH8rCKNT2pYYvkUNYF+Bc0aWhnxkwZZMPm
LgxyhTlyBKCzCZjd1CEyqxC2L1C1JERK3nRZcI2+T+DH2cdg2SUImfRgV4bx
6w9NHuMecBkoPtkWWEQjDVHQF1csawAP3C4ChoB+b8aIPzf/bP3B4u5/oMOR
Fk0hxE+Jfl/dcdMW1hBWF2w3hjZGfzBXihXG3cf18kRuqrPv5u2lVjlCZksg
9k7MVEsjA/86E/ZKZGS2DM/uD/1smr8u/YrE6GNslFjoa/jGcSY3DyIsErhS
0GEHTW5QCfJ5seNn+a5LOMXO3P9eZwgVnE9IsSmN1CzTp/J7em4dXJM504Ey
mrLPm3H88vK5wxfWldEa7KS95cFmnDBmTQFz8gqcupd65e4BH8l/RT1f5J8y
FrEBYhHef4XNtrhzjBRqu9B1iFTD30SDxCiIsWs4mHJAFuiFkjl4gSJ+qEb8
IrszRaGDcjbtmrHuHJP0OnYwYqg/P2DjT0dTbrvneXolJYOkxWXovDjGGKFd
nHc0x515+1QM40ykC3rljiY/D8XgyaLfI1Rz3ZnnckluWn8Tr7ppwWhcW5Ed
I2NbJS1hcondxgMEXMqZC2+tzGVmd1spWEVH9WTbA3c6v5RQ3BXKHY8OdnAG
wQ0XJiZyC1t3TKnjRhKmpsARGLhFI3VnCUhzqzA/LMs5tVgKgIyU2x3ajb25
5T+DAl766jFZ96AJjY+xrdkdgZjZ4TXfnMdp1sRhnzDuwtiPT40wOgO34Ant
2Z4qWjnOAzNNV1m3sYJ9VW3+yQ15W2xSPtu/8rdAfKXW7cXUn5HkgfJ3Nil7
c0Vos1ZKgpA6rVaFSBAE9ZbDipdSuFXGTDDIumTWVjalgWxvs0yUGdNaeFgF
dlXnFfNwZ6/He8woj2m20+T7SDp6F/CwyozD4I27FI8aWFY4prHaPBNmj2mz
TYY3tiMR9i4Fczw+nVS0474NeKIawGWV3ZEWB4iJRdqCj6Unf1rYwuKJ8MMy
EJ+j//euRE5mLvXRdEhd3P3vAr+WgdtK6Xgkk0xNjVPhnzHERoU/QpiRXUtV
s4ixLxv4lI+MI3S7B584hMbunC/Bnfl/ycAkufPPCQbX6l5hwXslThX+B1pp
B9oOkDOtrx62ivpODxx39Tm8mamEgEtoSO2DB7URjgg8dVOp7HnocDCDHiK+
xYPRsQK5XdlmdvRR8PTyqj5l5Ca874SfLVND0djpbbAcAinyzNV+rPldCuO0
7alHHaj/heA8CgHzEnKsRLqqx7R0BFVsL+MKkig5xLCeM545pesa6nPrAo0/
Ov8JfJLP5XPePddnLUh6XRiT6Hda39wn3gxOw2GNZmgSxN42At25c14c3NvO
fM9ANnH3nRCteNc06AW0isxok+ujJX/IPp6k135lkMjXpWfLbYCdQ+wV9gFE
WAdchHkRzAyHdKUKbw6JnbE2FJ3Q3D9yrcysXEmv/Kkz1OrJ1WGbFFgPMLux
Vu8ZETatEbj/8AMpVEM97CpGnm2Y22PJkUDX8rru7dz5pnhVGT5u3yEjtxzV
gBZaVkcb6yyzZJcwEtismE6e3Hpn9+Edyl4XAXG4ZDTxSe6vEdmxNopbcsMx
SQAe4ZDzBo691c/FCxusbUAKGsvo36oFSNSyJWz0PG+aQat3FdQKB3w+AB0N
8eOv4nEe3k08ql8ZHA8zXALciaa3klbsOg/TIVwwVFLddd28uoxtAliVzmh6
1H+13p4LsI8tCnqKww9EEHPkOpDqlDO5sFNLB9HNFEDNKb6jwiAdPKyrzPgt
JLGIjfJpnSeTGQ134anNVO9NBwHXrYyzFDbktgkD81W89d5adeZkvbNbtNTI
zzBAa502nCfczaHAbio8M/ZHXYy9PtBLSvwb0JAXEw91LGAFU/ezfuo7qRZJ
97brdKKNPh8lXiiKs9imXdXWPzx3lHgdWFmqlRzEo5OMeTKZG0SogVMyj7uK
4nc4iQXC2OFY8uC/+KMOZ5ss5hSGRbCwYEhxgqczN4YfDAkLuKlDF7DhMuQD
DGXCrFmdl0ZYsgyn755Lr0H+tYeP6Y8T80RdG8juzLYLUJ8kuF+ntK5a/7UM
Ky6N3VxKfpkN67N5dyASsOcQtiIN4x6JRsv2YUAAZYUzBOaVSSiHxwdxf8wU
UE7aGnhxDXIg9hiU+b5nT/FsBmnCQlJPnWWL/hNp0t5ibfSVYL1/nJHFB+AX
1Qd+TGLTMHa1HFZk7WXN1wprKQjqfz4mSAiaPXU/PfDicHgkz1XfcQumwu/F
TZRKdCndL9nvtLlun8obrhCr4sqDqNrZgEF6Ri49AofqkRUdEbfiabJyboZQ
6j+0OgQXOl7fPlmO0JdYVooESf+00x1iWzbdqSoX50u1RnWNix/JDuiLuEQx
2QMPqZpQz0HGjTy2fFOn3ZugSUFQ9t16XfdnnUNj2p9rM1DonGSnSkVnazpw
8xYMeqKGsCqJX+4mbCOu/ZX8x0DxOpakfMiAscHGlal2zr2aTcN8DEIa7SAY
7oGoLnUUgJezz1Mg5knn6P3tXbm2bQcSB9Hgo1bc/O/x7yGUtC+Cr7JXkfb/
Z/22IlMNp09udMKUcFc+QOfvVr+W05OBMBZMab3bfpHJPrV6MHokikx2gvjn
S7wpOO7QA8WB85hE/fJItKplGpB/YN4LcxSnFypZ9014IQTt2uVd0FXqYQs4
aTt+AC6POf6moohXfwmHsjaeTU8vvlwcvj00vF5K3ecuGWiQ9oaE5NYNV2ct
wq6AcMqRJF9fAk3MUMcrbLlk4Rlm/Z042koUWeFSVv+adesNbEx1P6GU4r+v
US0TqUDNkbSiwp02QsR4+DIUvx0YfE2TNuVhDUNdKcR5EWUoF67lq95V1Neg
WuaQzzSismgLiJBy/1JbPCtN1AOSmxrRkV1FIHKdqRE07XL/5HcReS+B8mDR
+8VZmP7HM2jVRp13A7NDTDjgSC2DS6LOEJnQIsywsdz2wh3zSz8QFJLC4K0/
m7px6kGWqCN6aF5poHMuwMT7vLAh6BXBGziqWddhJ3hnic2y2h3LJStFA5U2
d75o+8Ck/0vzMKbDLaAJud85RK8KzxVfVi6CiZ/tXYbz3WchaHDNhLH/HX9o
vTxNdD3BpotwegYUTMTO7kITd4iUC25xRT4fVJ8nbEIQQ1UJ4DK3L+UJXUi6
3wcTXTJmLlvzZrIN6wiHFj2OThdrA8huRGaR2BzndrKoLSW/oQJLQdcW34sE
J3tJv0BwcJOVx5FYs/pq8GDUXI9WOo5/+6WA6m3kznJglatyDh1jtSdcpHu1
zmbnjRGpkjBN+gKLTBUdAGEIkPA88EhQxESqYsORf4D/NKa/90FNa7wO7v0n
xP7mo8f4nh+dGc8Eo0PDkgRuQqQNaKjNslqhVS5dFJOT0lwEO8cifAZpPjsz
rbOSzfUxEfIoRRtxBXpb0UWHeFdmwrBlQ2PPn57gfTvLIO/Qsr4RSu1q0QCU
tYSsFYHcI5T+8b//aepsT4oltgQ6EnkuqLJwvcD0/pU/CuaOrIhTGBnopcPG
CgDed1uMBKZVKSv6Jlu4G+rhhesa6jb2BHvdvBy/mmiz13iR7WA8NawCXtTd
MXRKSXsBkW2Av94JsGQwEV9m1tjWDUzDDWH32lHM5muFUNkafDzKXsqXWa1Q
w/nYEbl0IZlyog06+3sV/akWe5EBubqa3zh7ArNt5I2Ni0Ik5ljFy+AxCyIn
g4tWmjkmOZm5b7KxLq+xGob0kxiUAeFP47qMkIhTA7j4E96SsgsVOQISvk0Z
wm0vtbrc4dvtnmemYZ+OWsjOnFNrjnPeWKm8Z1dhQqyucilyiWz/m06WiJBM
v6xv4jyewy4q8bfcOgu2bF7GQdeEZMAvT8D9Mug5H/6kWN2SfJg7VBGXcFZs
dFprUJgANiTEdrgSlWM9AyvUBGFfj7i2EFUaeffgNlCprSOWXoXtOSwFJME5
sOC/ypv8P8BcW3ekdiDHJT1t2mjplIDO87ZFcPViFOUJp+RrTinp13gGS7yD
X3l/RNd8cxUFqNaEOcUZkxmhnlol/mKXv1m/yfHdVWjJ0j09irb1yAU2AFJZ
1oPPPXUjZ/cVl/bGuzmdaVxgiQ5t1ThQsG9ppW/PIUWsuez77oDq/tg8iy/w
R30mfsNcnNqwrIvjmk+W4RJw6ZNzwIQZ+7LzdmcH55VezU+vqOfXzvtuXYXd
ORdg1+WQe9qwknDWOL/bFzlAb7A0drd58pMpXjo8LD+W0iz/8ZaFtMLm7pHy
FGDps0AxVlx08NUG9TLVL2Tr6RuTNVXpoJQpJBxG9J1WKIlUHpMkuu1DvXnQ
VlKYmXDGeyiqjw56Gdrqzyxp2xiDCJZKyvqPimaMI0a1q3PF4ydg/eeK4V18
9g1p+02FlNpIiQTW4oIPsITKOJSlVnpu/ezzwRCpGnj4LTUzcGXtRMQCwrsB
HqUQL4JUutQNlLyfXMfOfxHcSXoPrrnjXoDqRS0xCeMPzjdV8jC+1hO3+LRO
A5D/kkhCPKnhoZRPo5twCwZNSGlSErICJsfjckQPKwr732PMUYN0qOzzhXb+
B6MXMK8aakoP1aawbfpJqlx1jvDyiioENjPWiC61ePfq+HRD67R3bmonTyQj
6uiv9YNyhAoN8iftpnr9ZEDlffN3cm16x5vXIQg3rwkXq12YvqiH4kiisZtK
5n7LGgsaHOOT1zog8z8WDuN7DnXcWQoyBAu/GMobuuMCqrjQvuZEv/+SVj4j
efsshksEO1a4dUkKGaXGBLsRT6ZtkyH2Zt73pcRUhWPrwRbMYP+XHMfMpfTL
xobJ8sLWLsDBBk2X/izOGWmubUhelebNUW8wp38jU7YZAd2qER3yXkhIhOKn
yrxPQ56623UWigEAh91UupPaOTFss/gJC4ZjTvPAwj6fX5zatt35DuJ8/y6p
lM0VisGDfudHLcKMIq99bU5sSnvsdzJQQ5zy6yoCwgvrsgmQDct1/ZS1BASJ
h8kgMDgP3UMYnq8qML5grEHOlK995UfMuAfSDB8z+NbOM4LB8abno1DQWECS
WW/72hw5xGyMYR/mHJYeoNBMKDBPPbBQGugsL+ZzpbW5chKxa7gS7W/cHLA+
vM89vZ0F4eriI8+jfMYnA3zjT7/Q/GpwvXyV7uNCjTVHaJqjkGiJXok7HF6u
ljlq9VerutZkfQqqyG5f/b3y+XZ3UYf1XBDGJg9svfDS+bAhdCmlGEGZEDV9
nbVwY2k5nKvPXrpewzKjuuHv3BWB84LIarPTovGm7d5vH2/VyVgRmQovzwkI
D8zl834wUhE2EXdcKh3eMmzY0GjK3TOleTUaiPt41Ee7AIzAkSYr0SRn6nt8
iFouwo3iOoh35SkneeQ59qeCqFFieS7iRP9icFl8690RPOQBpDzSvFyFupQd
6YFKQi/zGLCSVZ5hdXeDeHGo2JE7fOcCd2b6mNSWBpLamSFs7KcCC9JduT8W
mZ4IT4a0ZpIZ56bbhjDD/7Fc0svBv7eCJH9xZhKHVw0MWDE/KbvTls3DzTw8
/c2zu2vNCKlhCqyCe+zx3nQ7QYv60kfBtYrogL2iaDLpRZX3w1VedyQt7Ix5
SzddiPKK0g6UEd/ikw3VmnnWN68eu2sGz9VD3/AGEi+QpMywcoUUVfLZNPfz
rNiIx4RkVLyZfoz6jcGKlHTEKHStkSRCpOK5zvS+ULhdjKJuvYti8ui4x3Bu
/qhSbRnrCWv5mrVQRsZvgIFSj4DDy2u4Loskd3C9zjQKQqH+o+IhMillxCw7
irAspLuxOjCDBm0LXm4+BMLbBshVxm+GtP7ld0pFyVfw9VgVmfpC4+V6JFSC
kD4cEDq67WGcotLv+lo0xQG3WksuXEWELdUHo1j53GZ1D/zP8yh9K3mo/mEi
In1hFDRK/5Xlxb4/GRjaZ1uoeIP4CcmTFCXGX1luosv66f26JwILPws7fzPC
SqOGuyhPNLJTVPCaKZa+9f7yBz1PHzei61dsb19WG9xfwyboiOC6PTneJZQD
Yl2gzlCInBC6XodOFBf+c6qBFygBPSDIHYJL39bBjX4Ayk4XGLA+/w8XF1en
2AdGpzrR53SfjaGHk0v0vt+161uzKWK0TtSDSP678Z8n+358vNsV02QbHomj
Q0kOmwWaI+WctSHuD3XjoUwA88oORSADYLvE2sZPicwGjRPdL5tVveYPnn3Q
+6As5M0njJs5oEKfoxmFuIwmsDOoFjKxaxjveTKzoEwioP+e0UxeStGhFLMi
zDCTtvICqK19RELbcgdg9p9unkPJycwjxePkMPMsczyoNJx1rCAcDKAwodc7
OP480+RKhqORt9KXCzDf2PdsZWyVvTA3EmugLMOra770rnInLyLs4fohzNvL
l9WGlErZVwn5VKQWk+tclQcyzpAkLLhlMz1QHXdOSl/deJUEh1/hglHQoYQe
TW1dKfBZLY3FJCEtmrzmkBZMOd1ihrrNT7Yufrr85aLVLrUjBP9iwzVrhN7m
MyFjX7t5IPN/0lEUiNOZOZ14WArX7u++AEYfBalcJHv2pavNBSmSGWTqVijY
V/THEyTmhCZcvNbKsTTGdNQhQ2JyKU5DR1LLuCiVrgJxzCD5nEAhKioAwRoG
fIkOhOO3hrRQY43Ju+E/nvPIAgkhFeVrOBpHRBT+KZmU75H0uEVGHsmT+Dd0
u1plTHUT0M6TZnP7oDLzuK4OwWeONqFqbpcDjT2pReORrzLRcSPkC2tAQYCb
aCG47DfDwl9ox2Oc0JzZWxuBvCsag9StdLJ2zYw1kJMJLGoYX5Y57JA9XUUh
EyTWU1V4toMb1o1zsT2D25ZLr57J4pkqllJ5LAyKjQy72I6N4TSOQ6qL2fF0
nNToASWTaC+h7x1V/b6WbXUDhQRfhvjk3i4rTvueQEtjucw8EoXA5Mmibmsw
JwItuocMAejeSn0bMuVaRQjnsfO6LTjCBNj0hCZ7Wz5myM56/LrjI5rYG/az
Th0mjPETuye79wH1nuQhxwQQAAKgeG5GxSvrpMjdL1ynhTIooo1VXo15mShC
+wcvIRjQX1fUIhTpTspTGVZ+IR/jf0W2ky5J4W4yNkOxbD3VXp/uKcDG7ULg
tnhanxQCO4tIDDmrh9TiXLrCA+0naXMXtP+s9dqKtOUkyzJtDnhSFlE9E/XD
ffUXIPTpvhtB8vBN94Z+CUXXIH1+5lv0SBl461C/7tiPEBOWM+rY/5PZ69IM
V/nPIrGCkjvCitk3o7qsN1axWBbzrZ8bx7+z1OaesLnO9YOi+HIYVJQ9fFrp
ro8cSqZZaeSiojbSmEKRYKrF9wgUMZ2YzjkncYqQ3ATLxZ+evU2bXmzhG0ZW
PhEEwQLc1TcMzjBmwrdGn2VpmiLVrQh9Cr+rtK1QhOd71SS1unANdtaRW+tA
h+sE6BkY3fF+y9lw3kDcL3iPpyibXIYTxMv7Spa8j5qDiowqY4xqxyrmCtU2
fxcW+CRts3nsR44lZoJB0JOiBCSaLID1MqNBrDWou54k20mqUar2vIQ9VOGS
/MFhqYHeyDInsjHRF6jR6/xIeR0XFlozL4/UqA76TGEFs1k777LF7ENaLUWE
eRCyzliWFof9tfepohEku8Cph5vS0NriAVOcJvvIBUDaSjwErvfIJC4wnfbp
ZlXhWWyJOdTrmll/39I9SU/YxTWDne0RkUE37IQRAaSx56iWxDWU57xpokX0
3vc8uIeWGO2WwgM65jMw8adYNCjqMtW2l0eiXCXRBdCJ0LcUwyp4uEuCof+t
qTLyexjPSUQiNvaPgI6xgQuSHInb6CVZGl9cyWQ7eNvXjOOF8MM+moM0ikBc
n0BAqdzFCvlZ02jM0XlQv1fREBBraYWqQW/oG1AOcqiCKuRcQhhFKCuYoite
MY60YvtV8txsFdQL3BbV/km4kCMmKtiVvp4vgtO9karKmVTxuBSJfz4/eWI0
DjuDfQcqS727G4zrSak5qgpMhGSshqepWVB2Gk6tbZrgoROpY4YWgvJo65xg
exwqFcM8hx4bUrBixYXLp6Masr5j4KeJPJox4YQ6snm73xrKF6vnBf0EVUKT
inaYNQwHifwifzxcZ2Nh3pSjS8VOHcnBDNXqCQmkNhAu5/ILbJYoYFPfqf3x
WiJEqMMDgWLlD9ew7L8uaWvLc5mSWeBcwAyxVHjCZA+RH72GetxRcvMG60z3
SL/YKW18/gT88zXFDN/b9gmx/d7eBvf9xYP30kiLPcb3BIvFqC0WFGoGUnht
CcpXUHuAs5g2rTHkFagujYyN/axlm1hRNvo7kx990lKtLN6ao5DJDzvfXU6q
GoNsAXg7PC+6R1qSfjIEGOCvyVMG6VrcBAI5gqfKBHLVxlYGV4NvO9OW2eDY
v8+CnB8im40pn4PcanWdu4A8ac7zZ8NLfd9gI0tPBqsU8Jo2Obcce3sSisKl
9mIbcuSvNIrMbVpsyAGWH8Fdrkpyc+TnlZZedxyfRYUEsQvjtAxEFruAAkPt
X9MaAnV6S00D8GUheTFp94Ziy6txwzi+3DkrQrrDSIZNM9Fhhv469U1XGu/1
UdGXW4A/qYHK7bCvy7R/+imCXANviAWiBhr/0WlRTrwN2wT4LbLRusMYe+De
lyc8Ta1CEMwtU9cDymi1qlidqDSypCd26dKNMMBRwK0o8z5Q3L4bugsvSxvs
QL/eOho8+ATYCpnyhzRIPBtunp1JnbF4PaQe76kpGOBKyTj6wJ1gnH16YCwV
s/uWmWVubI+mx0cW+/FssaZOA2F6tf2Pn9Y6tMCWzEkbzE6Gb1WBrMq7xs7v
yKZ7GVbRdgITbH3NS84fmANQ3iSx+KXSyJ/tTk4Ao4WtvBz9/vIFFmrurMKj
759ViK2Rh0k6qfyFrL1OaAmDL9sx84GFCOIJNagcnzEh9AYsgwSfAxpbvmce
6gm05H8xYYSHXY+2hQHQwtIQiNTNLjXHc+AqX3mQNJdZfTjFGqdpDP9XA+9v
A0MG0ndJT883uHN15HmzZ9ljcSXkS1Ct6saWK0POuAQWZ9uybyitVR2uqMM/
qpihlLiIf/VrU1CNH1QoYAH2S7rqnggDwyWtx0GMkOxYyf6UqRsmb8GgwX6F
bI/0QINRGpGS2mKd4aQ+zfizwmp5iQsiu1dc1t0iFys6bVgMWQ6oz74R7NVf
W6PwKXfWC6Uvffe9ZnvyKGzbsXd4ZMu/Vb5LpO5qkfbylQibt0mXCTXrbxJP
vLOdNcTAPRVJ0WY5Q+vXpYy04reuQUMTpeyZqUDPTUn96oMtUt/x86yFZCnw
zHYpN9j7DN21OdQsaN6yK61zqX6dPLJ52b721bzSqu4f2lCs6agI5I6rp8aV
O37cV/MRWFK/7TBe/YiaiLGmXKnIEHmsLcuWFueNwgC/Qqk+ER56t6a1kNDD
FKTBtkeazWahV3nXahZHWaKDR2LQGwqxlthBN13nSAAinSwUsMoInv/wIGe+
/NBKG7ul/U/ASw1RtCdVm/cj86pIhtGBwn8uWNe9855hZM/utNd6ZtRmB5Rb
zYh1tuL031VpKIQHjL70f6KABNFqOCloA5Fu9YhQwTLSpzPkF8H0c3aR8IgS
mZ5uPeDK/Qa/qFzhH158/4rpTqwledYP3BYsSE65A400TzIwiv6D2Nj4AhX1
X+cyKKKdHEOdmJD0a9+zkiGr0HMnrj/Od8/3BBDJ6aIhaXKSWK3cBqKsj5/y
r23YV+foWT1JhAKtGnLAgfdh8MHJx0vYz5SK7So/gfu5fIQEXMgZXtPAd5Ze
pv5rMo42I90kTNkEpFrjweLXZCAcYktwMD5TjjtyA3uWC0OIiu79WGW/OYXr
D1/pZm6ZgQS1zpIAUIJMdstKH0wvbfcG+z9BVBhqwLDh6Vci+JNroTUz3qnk
Q597ufOJx4uH6RfjKhz4ijBNiD8+dFWm7ciWtSNn1TsbInZe/kFb7S9aAGRc
CUqa3qR9rmEi9kMDEx6Arv8czoJFliuWyddmQWnm3tXXVNKotIz7Ub/bGRUz
mNh67bm6WX/Dir3n/OJ/QSaRErbspB9WTLmYuKQLfrcv7uXv0x8gAxKKDQ4y
fkfOI+lFMStRx4La5ipxfDLP/p4hxy3kOcVDzpkVbc3TfaBpntZ3mSRcLPTn
foxiZftVpGRIIoYfyvNZoEW5S7n0knoknyeJDot0ztIZabCltBB7e5VB5jE/
Ptqx7fXYOgvkMctjvtQxmPI2rk0lJS2i09G9UQlII1WaIL+sAgqzUzkh4kjW
Pz87yEJRFqPaAwLZwJFu/bS77BQ6wSNGxvQNSEAHuG4BjC8lIB75CO98f3Q2
/p8i7wYJ094fq5lvdvqmEn19Qb1NsD6rgwTfFuaQ8hkDWL3ezMbAT2HypAeJ
o14ngFJP5rmafqiMwFmsNVTHmljjMRD2BqnToadCKjSES3bX4sxuOCuBhTi7
gxZuln3q43DaHAawVlRWK46FB7iEOHUwp5hKTFr5T+9oiR1MFgVlaqWv3u2y
hoSA3k1QiDMvEF4vzPVAaI5AKZjCEcNhd5gAuKhw/A269Nis+6RTtY+Y1Hrn
FcctlnwCE8Z5l6kT5n4pfDcKu5S+vrpOwxyK0sXr+2iakhZWatMQolNM/l8R
oYCgmPrhOeA758rcPnRVtrvrGb2hc3GDvWltbSfbLZjmFmnazjYomKaBtPW/
6yFMH3jD0CQ1zz9wLPIR2i4uVATz1BbEifPxiLf2MMbMbiRg5y3C/1ogqybu
uVaAktzT5a74m/XhHrlW5VMCQmUP+M+vmXF0TE4Jh4IsAcUfW8H8SwmGbPT5
bT3ppBdjdZA+2RUbn08CbclQEo1TjNwai1HnYd6jKcS9rj6PGEHtCi2F5vs+
ue66X8qRUPwjzXTOdu5inr5aPa5VwSt68CaShdeLQ9GGOczhJQps4kdhcbmM
glSiEZgmbCq/Oq0/FqPi/UllKm23mP8eF3uqGGtZl9FllMDFsiQLc7nHmXj/
evMDsrQIPmYpT2hgx/Ra5Ju7BM6S5zKQG9l8T7c0fEV+92CyA04p5nxgPnpm
fnYd/MP35Avkg16qYDJKnoizAhcKJo26okohEtOWg6QrxQ8EvnvXUWpgbVcm
VRdgkiVJp3SmsLWpGjvctTWSjImhlSgohxzSKTEhnIonOpQjY2ajip1IH1Le
vVG77btcJGUb4VJHJlch0eKhyFaUDvrJjT02xEFVOXngFl78gd23s1fvQo3F
ELFzgyqGKFApZ/iHac0fRwmMFtKG7TkchQXU5l9/p4zXgBRQ+SKA5vIRpVj0
ImHwcF0HQ8xRUR+iqKiBC1xPJryeSX4GKEEIIrsKhUJB6K/E7Cg2wOjb+p1+
cmPFw8Cjkhe6/XzDuWtlJ1eOvNUL15SPLRlTWObk3NCHzC65lwqTgTHVNlGa
yBsq5GpyS0yY4Av+ZothLH7SPwapg/8ziywiVVKXbGpCp7DIgXFAWS/WUnBA
LwMUSt35l8m26iQ3goxJ99pduUu5mMYmN0l79SbPCHPGBdqV14ycAQd1IdPd
cfDgBSMXZT98+5oUjMmdWrBrch594dJrdyn926SD1a6YE1R03yWMDf82eD9B
qHUHcUi4u+ZSALubS6EPszpFNWf+5vSrdl4jwd0t883cmeVAm2r5GDUxQeMW
qzucUANK8E2WUsJ+9rpAWa0UyrZCrAjUP1I//lpsLyi8tFGOzV3yiythrG00
Z1jmXylO+jCDHwpSveLprt5fJ4wUKbFhzbhUQ9mVL1m41wE34gUH38+v3xTu
DgimXt8Ewnu0id9VGJcMBxRvVL3kplfyKsNRd2pF15Rayu74ulnKCHsfJnRp
0lFggAtnph5eg+r5oxHCP5HKQP1O/EFX95FzQtm3++T2e2IcJhpSQWpH4hNv
dAoLzuzCXS2DRyOVYKXiMEFUGC6FcFJJqWFntr07jao4sIl1YR959ryyIYF+
EfO7qqIFBY1P2P63iM7JLDUlh4N8b8d4eMhvPTMHaN63Th7qUI7XXGUfYtki
WccVb+Hpw02dZS8t2+E0CWWOFGmalbSGtVB/e0uif6TGReFlKo+PNMaUMuWj
T9xGqymvSTtsae0GuCuw5PYRdzpSlif/+vlFqZ/c/Rf4SUKDkjQ2kZ75f+xo
8OJunZUDT1YX4T0MDv/dx7ssr+GMtoCOOqWjdFA/90+OnLkeEcuEtUjNGVXY
2k0FSqF9mMmDRdxolfNggNTzpaPCUI/7kfc8xmp4BkuEnrm5fu1jg2RaSb4N
feQW7hiZKAJXZ64G0d1ifFoiH4N+lqgHwF7/IxaJpMqSJJm0isKJ5I05EMBq
jH4af8nML68xkxjvJsf2JzTHybSX0Dwr+qAk4Xuh71hSCDXp2ehfQHM21lNT
vgyE6CfIEPtl1Vqs7kxOEKCNMN6eJws6DR6MZ2XGdKrT9wqJAwE8YtKh0bhg
jJoUNe9LdxaSgX5k72H1j0Que5wiUPiWXie9D5NGFVZjs+f2ElBQmxNpludm
hC6JOhkMn9FMlT/z5JuP1tjxP/qIKkATVIsdiJZjxFpymjOlaBoRfR8I9AU3
ml7o+S6hl694mfSl5JK/f942KUg0tAnGtxaesdjPLBDaq+odtSPAA0TTw4HO
cCfO0j+r8tjQJEeFD8p5FqmirY0nUhK3FKL8XQz7HQjxbmkO+mAA3bMJE12d
+iig+2klmDZxD7I3gilWZ+1Z8R44/u1V+kf+sSzxZ/2A1eDBRb503qHcyQa4
/n+jCphek3qVGIVsXP5WsHYgDj8d9yOp7yrdtEeTQ8n1OvPoQhFA3Zvqppva
NAXXL9q2U2na6jjvcR+Ia0Gs1bsPrABk0Y6mqgvlgZd4c8w6FyTOOqPofXtH
xeC7AcT/lJ0XYGCKolRcjB+gLHGH7Z85noxziaMPmTnW5HZVBVPsvAKm29Si
oc9c6dDJhHRIHfMPb1Api+gJ/1KKu3vkcekENkEBcHWjf7uGEAjFuS2+N3Zw
lx+waZcoWkQhfJvUV6frPNl/FLJd3EFXa4WWl2vyU+xOOihuvYZ1/K5rQ3mM
Vph3M/0U74dLtCDAuzVd8hXzG96t1I6hrcrGt4c8DsOoWgwB6dHL6VoZyt+7
icmTdXzL7fYo/qYko3gyevsoHwDyTON4wlMxf2W9/ZvxmVWI1LFnPYdHoJw3
IIidrtLrUe790KBhnbECTdA5R2kQFsjy0dNVsLns2Souus5M6fcNvvCkQuKH
HwfIRW8gpQEi8b0EyuBYiDvS4JeCXxDWE10Lhh0CgbhXOM0NOA+rzS4jXVKM
b/sqPemltPi4tzgRLP+yszVu2hHzt9XZm0d4Wfkrrq7YhqMbl3qRUrGXHGsV
J5b1IQgJCJC0toZNygEsrFC+DaEPwz5vjcH4coDgViw6SLVhID1tZT1vX3Wd
IRlI5MXF1652owY+TLqG74bTv5Y5pvk+d/tz/m1liUdic+bSaE1wA9HR/17w
qQuyJScdP/Ip2O0beI4Ifw03bvicw0ELO0VNkEoSBYqf189az1ibT5zx5h5f
QlWJQeWBwdx/5iuWtmA8F7t0bAm4XDZNcUHzYs/OvSwDS1r36Y5VMNpx4mUq
C2dZ7k0UEsgHGXMX4rc9GtpW9cVWo1l1IuTi51rEmuBa64km0BkgvOz9g49R
LPWb4ioK2wWIdITpjM2cqP+YfAJ6qkMwy7iB3EuJMeHdPRqClbdlUBtrBBxH
vM3BdUzWg0oB6GqUuy9w2h5fIumhJC+Mkb6uuJW6HS+o3fE2xspKLNT2g/H0
c96TkxYwcJppoUg9o/mqSrREH77oZyfTX1+RAja7GXzotNf5RuJQZkSc57+Y
JQ9tIDQt2yk309cySiBZtqSU5Z15w0viQnglE/uCRIvZGAGsSqkxjEvxaoLI
petTLrsl1noZHjnKNQr1HgsBLz1N7pXltT1flmGycW0OohyM2sWqhf9Hj0Q+
rkCOtn1J7GGVkF+5+xJ0kOyTjEVn6rA8A3c1IBrITXNP/pMgFZd6bhd3wPxa
uq3JhrgLqFGP4qyWhg2sjrB48yX8+N9iD2iWtBPkD45p9pWm5WGFM0qieLzL
wuhiWGkBCOaCacYBGtI+4wvKujIYwuysBkfzey1fN+B+af3HOLmfamtgsttd
siQpUZvsMeEnLo/ZKP1awbgNnno5JZPHafGdM5gcRFio79zOp9BdUgOx9gpe
5i4XRgilOmqqGa/9Hr5Og/5KZrjkP3A/djPnwrpDsk5KSQsqPD8iVt9ItUsA
eHAsv7/uIph+bDoHJWe3G5Vs4hfrgIxbF6BbZTwFkgQUvg+AqPmU5YHjoepA
mOLOqfuI2EFOv0z8jUe5cQ/4BYRwKYXjD/wjTpr5tIslstwNtic6LM32JqO5
/WVKtQp2PLzcT9J0qaTy1gD+M/eTDo6DAR8aVp+P87q6hwE9ZD7dMoKwnD6Z
0HCE/jnwa+utoklymcL6JDb+DuTOG3YK/86s0g+/vL7zEVXXkjgGnyOSwxyI
BcGd00y3axcyNw5TIzOWYizKXa0BFO+XI3r2oWW21oXGpMB070ymhHLUhp/d
lvvHu7v8XL91XmNbTsxajBNe0NOQo++vtPpE3/FbHjnpF5hLJvh2HwfHx1pv
UcVtLHuYqbNJUDMjN77U81Xn/1qNf7CR1uqmrsH1hF3mHAEiYlh1zmZsneOy
8XUPCr8qUF3pk+C+OflVfmOsgoL89x8gAln6Eu9iGSTLKFBa4duPiHFXmhxr
e51MzJhQNrCuhiHipMoMB43HaVYc+b+Xk8HRijsLpItrvxK7bcFbf5KVJxg+
8yL2en2ieyEnRdk2B51k6ipGEW5VErx1Yww5fMrQHHjaDB4Sr2mrwoFqu/gY
o8GWWiUmmcqFIC/eEa33ekLeaNYDs17EPc/Ij/pursS1PtD8qhpEPdq77qYd
Zc6npmqrKN25iK2xhuxqo6sHA8t+jaPqX9Ows7wezBvMzJ8NXjuH2nsU/VgP
BIG/yj86npiT/h5OXIjf8+pvMK0KKOB5fS406vRbMAa+ZQsVMl2DZBshqrde
xTbM0Wh3VcdltTYd2OkLUuzn304ll1gopCCsSCwgvyiS+rymCsM9c664Qz0t
u7nJssmPBVaOLAaYkWie5xjQ9M2FVb6r3x3EVH2Eha1OqiyAJcojxJ+e7Oa6
i4KZgrt2UsVmZ6kkhm8ekJeXu6ma1ppHc+i8ZuWMrsYYiPaOk2XtvpFbPuT+
WRdn5LdqG+VdqUCSvPka9SdnWr8Vwy2SRh5NfMoQU3p9b4GHnhq78QfSjvC9
CsCtlxgzLKkaZPTrTbRFIvky1cSWereHRM8Udzs3TCrh9QD6ErnR0PLZv0u/
EPRDj90aDvnsGs7sccssT7OCzEv1smzsbCzBR4+dak8MwvdtjngaMVbqOtyS
jv19tOQ69Qxrt1OgNI1Czy17zKP1IYUmf7qVoDubjNKAG8DWc+FL8IQMt+EF
tfs27puGeEa7y4i7PileMSjEX6JcR2VcQfm8bi3J7Oa1ljzEGVkt0clPPVRC
iR0VDBq+Y8Vv8sKgt083dSP6E1D54MY0l2ZZ3GiiuscR23zrt3lVFek9qmvN
Pt2W1HWrppqvuzie26vainKQzP/FpJO6DHoPcrf0xqNo8J/3anYvjlNRKCCr
ttghNy22RFCn/UgOvakRJCwWFmozNFkURUfd2FFw0eASbhPgzAKm+hBQh9mF
Ivn715WW+eh2/BguMI7Von6mvO+4VymC814CSOLvd2jivxbLzNmjz2cgTJgU
dIDb0k3HZtqtvyB/YGa7p6nlSbp6glFi/TxTrCbhTTzjNNkJlY+iTDbPLaXB
0cESqZRYp1tQAvI+UPTeC+fMYIkoesAajrx4DQTmmrxJeY2RK12yJ6qW/wmP
5wf+dgMXu0Vl1LIrEzTRm57CPwbZvfS5oYb78OhRsNp7Vcw+Oz5p9ZIOAJc7
3jdOV+NpKSO2JSArX9H62qV2+85intWTIO5C+6O8UEhkFlT57tGMb3nJfG5t
HTXAYvqakCu1x+p6dTUgG2U25YqWc9rZ3esK1C8YL9NZnE1PPYWrLmJIUvem
kZCiDY4jhwBZBCdJChX+P82nGRoQuL1RjMveVjm26jxzc5OG+STdm4y9ISoT
pXr3zGhh2qyTf9W0Cm6lEZpaypB4HouIHKO93/eX+fVO0MMyvlhM/0cvoTDU
fR6tJnG/mJliSmOdLiRCra57RM2Lk2SCzfgnUXqthBImata4VTOko8qKIuV4
mCrgaMvrMIZCtJPLJtxpUync+UUkMq8V6HGN4NEQI1QK9c/KWc12mLS1kaYv
wZzbJ8BQlz7Xgb+OgZ/SzPtD5JKnJfxkbI+WmB3P2RDQcQGz7dDGB1/czf5N
2xFn5SMWbwITv5N9Bb+u7sA1ciQH65kBqvpVHyKO3UYHb+UMBkTq5mjIzFwL
oyENZRQUSgOnb+9IhMpGuZ3ODd5CP0JgTAQ1xK9hi7IgWMSbE0+HumdVmN3q
Iw1nlBey7EFzYyD7ObLzQQpnWAYCrcxFBa8DtwLwQc8kdyGwak0MlcXXWkrv
rgZ3ej4KN7qgG0EwRp2i25sTIwciaagh9dNZsTQLevt6ypJXMIZCI+7S1xp8
ztVwe6+8TXs3gjlp/Ex7uK22Od+eKCSFTTF2FzeGqfEyAEqqwQD+YmXwyuU/
Su+56xy7aLfbn6TyG4fJIT5+M4ZPb4qBUGJyPXTbbMkCBv9CVhw6eukHZhIb
G9RmV+TEndh2MovpRTCJiT0coBGp4MdkMEpxgQh8iRGnI6uKbijWzboRQeaP
o3zkM5AQI/Yc1YwkT3Q0S085HPCXBNpBvN11x67nbYm2f9wWANBBzkaYLL0d
cPx+JYHGAE81/CcqpA8lYfVvw0MdfkwB/hulclZ/xCZw/i3zmLXcnWnEBMbk
aJPQEUI3gB/LAjABzQi8BjXwBDJf1PbmrbqrTEjYPkp0QsOg4df5qIooiYGi
bVCHsKzJGQyz58JHV9v+uL/jp5ZXKM00zSSsKFNbnpmdM0pk7PGexVcJS7AQ
Vwr1vddYDS0JtXH8Llm1KijIL0Vu+o+E4TaRCdsS10DUAWtixvlMcBKwwTwz
Urgx508MbH4iGoFDCu4Wu4R8dIHnXU4wxDn/SZWK5dqZND14qPoZLnZT6LJf
KOI5dn9icZGJhnU/jCMo0/8QvuFnxsjSwKoRTIcLnKP5Bkbd3WtWTegoDJ2x
lI2Zu810np2GuXPJfRiASRRwitUC48kOJnPvOFUpvxKgY/IMWfRhRxt/c0pZ
R6g7mQp4uUbRMfY6y5/seZHWIuQie371q0uwduy3fo+TIOZiUqyGpHjq7K5E
npnIpQoh5ZrhZ8iqKicPWMqA1SLPIRilozOAdt0Wbyt8USls0KTbRO9OJTTW
3H8TbCNOOtRexjqsQpXpR4JyJzG5PCBT28mPWBh7vk2kOhW1xuDxCcPn/kQ8
Pk3rZUHhVtwnQ5XuHSB5AD8iUD0IPhc7JZ48YYRTlLQdebpRK5CZ3eXjIaDW
ouzjbSq8mmJupjZvIY8AkhINUAltTguQCUzheLB/Tpja9AnClYRy8wTVVuHy
cHgoUD38TuxUkvBubuxuxgZ4S1MOSzXp3YV9wM1yjRRaZnXPAa0NMZc8efka
Sv2HrkfdTrYZMzh81jTdS8AihjlwphW7nk4YG8fOGMEK7snwGAHQWJ3CDlJT
qEvJtDSAN42L91c8LLw2JTcBp0/KxG4gX5LZ3cajUatlyVxXtuLmWNqquzpt
pQRIMVlpe6AYltcXdrXswPebyNaMzGe0B0TaH8PZD3MbrZqtQjLZi1kJZSMd
WlgUj2WtuALpGFuuncmlnVj70FqtDYVoRqIlFRpo/GCzWz6Z6DvWq1lRJnl/
eNng+GYLiBgK1clz/1+6ehD/0wLO3PmMs+jpNlTbfFOkngrQYzSTwUYRf5Gn
cMNiSayBc6Uff/mZLKd4d2AXxX6F8RQY2H6+LfPwieVqErpsvYmcKJR5GlC3
N8POk7PUm+lk6zG+25v+i5iNfYhHOqQ2iVTIv+p6mvlpDqY60yCVG9BPDLfQ
b4oZZciuSZUNz0c6Uqn2BDFY3Duw2tezFKjO331gXiU8X4og0FpbI3KkaGF8
jKzVe0r9ImGPnmOnhN/EVdt+Bz5HnTXq+vENfkYp6sJupBh265P+I0iypuk0
wo3HBv6AG9QnSD+7eM+C9Rm+pG2lCd8QiMKVbGqD4jFwixwcnjFMVwmsp2s5
rQnhLCQz7ORnwOfvNtMvN/PsO/SskgY/ZUPvQOwmSZzdlkB+Wa3+7GpIQaee
4hmcC9YzHF4/GcSnK5IrH7Piej9oB+O0BLhi8Yy/lHyFPkPs0zLrSuzk5t1T
Xct7KbAQFvX6zPsqBn7QMch4IuachQj/EOfYILoexuKMe6408XwCXr5dCRAJ
JR0J3yCENRaSlAftNCqqXwvWpa07cPHdcXeT7bcqbe6eWGX7VhvVXJWtX0bx
AQePeDGAKJjcdGLP0IoEdRAeB9YahCGLESYnoi0q/gn4opIY64/+Bg1QTRFY
sHE/kwg71N7TKmzBuxAlIeA67XBs1lZGknQaAXjMZwQYPkYGYsOxCXKsv4ww
4B4Tcr5pF8jR1a6/zyYHAOL3bI4+FAkaj3sTbiAw9muGdmAIfrXvRDmgSs41
eKXXSVK2WtkPRWD67gSUrlsPqziMXsBK62tSAyAdnztV1F0BXdkGmTieilye
oDGG5EzQoBOwiKObjHAwsm4bkJVC+CojRhCCOduOwu76I0fNrmAAeWf0Bh4r
ewGBEIpEA5J07Gk+KKp6OIl666ypCv4aidFqb66TqKHVhz4/j1FYwZwlYfjS
/cJdGrQJLKnNC0/Uq8Do6Ii4L27IWkPvCROGlgiZmMx5ay/RNmmacRdN8qqp
QJ8uscjwf+D9h0vtmN9xFsjDpruKoY8500hfURl/wv1hB1hd6vTCGYkkhgjB
Kah08JS7R+fSC/NGtV2PWT2fJ9k4gCKuX1oKL43CqYTyBxRD5225r2d7HtPT
xjDX7nn9gGhODfmgoQ+uo8AZ5QGxaL9ihj873ItdhXpoiJBca9JqXHdFdb+D
PPBIeGt7smNvsuLawL8aSueto2CbPvwatAKPNHSLWeVntpice+U6/ecHagkH
zHFGFfdN3Y42bBu6u/uAqYc5MvzoLuQMuhsNnTE0doUxJSWq8C3UomzGRURP
CejhDuMAt795ohxajmQQTm8PWRLrafPijcXweYBiLgewIKJXfoiRAyVVPjve
X87+m3g1Hg9u1yLAANRJli/fpKEy0kMVtTCossr9lj40FuR9b+9cZv7ofYJi
PBGnqwytaaEiwukNy4sN/CrDPLVRGJQSutYUOU28XBufdxgSKJ4OGyVy8MX/
V72yJmi2wrT/RV9wYo7Or6vP3VQUjP2/HQlmTA1hxZoMVrER3YhYPw2hTpg8
2YqprhxmWB2HiMbjR48LhhVmcRaKzaWRBJu+RLNVDEZ2Wt/Gds6kbLxEm8cK
opBQHRRzXo8DP5uMMFVUQZsiCyK/6/fkvgPETAS7IEn8kg2i7HgKo+TMgs6F
zxgKHvWZgcfiG77wUCs8e9+OU3JxaBJmWnx/5e2AcIuujr19gjdIXpWnBdrB
jxH6NpAqXewiKyjab3O49SaJXnYHD3wBie+AaJQ27OKDJuR7cLBg4covipIu
YS1XOGGs8DwAe29ZUs9e5Z9fNYbEE/uTILbUaBE0FDAGfbGmHoqP7hJBjvb4
gAVfN0capIu0gcA40/SZo5StTG9kaxSYuaIj/eXw9oNLi76cLSgX3HM9cfLL
18tXyuUhUa6DpoJY0CF+c98UrrhNr/zAnOyDuHLMhZJ9rHO5mmZOtWzRdJdN
M4eRnKd/tVUmrzQdwTRji+26rWXLe9/fKvzRr7enG7VQ7lxOyzX5ejzyNnHE
xQXjXtLmKVSPfgq2+BXZhUTFdGP8ezbVulU3KNpJCaexS8hNSIrSXb9VIra7
quZup53F38DCVsbwIxce+NMsoj4ug+oKnF0httowjsXvRpJi+OdtIrsc0VAb
qHVimvuTNjiNbq+f109C2/S8H7FftwuxUz/WyYJKTPxVM3SBcc2cEFjU8TA/
yrLPrtRJLLjHzCXFU+pZ3013SMj93oHCY8vCLzyjoOgVQBXpylechA464K6l
k+/qVyQc1stC+CcDC6xKdQqtU3sKPdMEy8NNk+4y+o5QKgfbidmIOqF3lhzS
BUtU6aQEQZ/ZgNTCDi7h99nxiKY9MDVAGFMVaQc+WwvMrIIPROK+pEkvtngW
1Ln7k/RceUq17ncQHjQ6/8YnpQjkG0BBlJKePB2Ilfnmb71W7db23Xm3yaHv
99Ilj8HA7edbfpFtQXxPT99xDr4aOQ/DrVFLcyipdW/NCJUiD4H7Mo1A/W8U
m6iqFIwp4iYUtoQt3Lt4KdNzqNGbiQ/iaNN+84k8pZjDGgeYx3RJTdLqssc/
DPSpyis5C5ofOakEtpqrtolyFSsoaMJp+cAzGSYWaB1jp3qaaAhJ7a+HaBCg
YdxYiyuE33Whiajo1NyffvDSymcMndEsmcTnBh4XPZTOwUNOyLGKwhUiJ22o
TmpRhkac5kvQmNVfKCA0csj4pH3cyxlB6TP8PZRyAXMnuEB8gQ235pd7ELUv
Yji9Lly9ZSzp/swkjEe2D13ckZO3KNB8uzH2Vk4mNHtNBMr6KXVY/4PBOKWv
/6SKb0uFd62/ZC8KwxOo3/FvDNe1HqsWUkEnMf8iVz1e/QJ6Sr7QYIzyL9DY
UmPcBStCcgF7scfbB0Wi9A/jRiyMEOkjGxnzstRXnw5Ya4Srl1LFgu6FcoE9
hnjvNV3kNzq0dol1DpwlHffO0LqxACdjr54JamA8zhHmbF+/5C1m1OHuP4Gh
yDr4VCsBaGPexAnFbL4uznwM4t+k/6jajo22VUhCA3q+8HBdrrYflZ3IYs4a
hM/4SbkP9NBxGf52JmrEOb20P5GQoBcNKgiWvwAlHXDZDjLcFhcLBPr8p2/b
ZFbPSyE5Xg8TKl3yAdFN9eZ8AfBi24uHOEZqzSS3+rPKLWahYHcVkZ91K5x7
HiJNscn14Djw9xbu2oYjbiQawgzfJu9znnvFatL+0/BCSpScVKZ1SQJ6Nshz
lg7qw4cCsvWMPp8CVEje/MyN6/3ivTBpvA8s2Z4csGAYHLGgRBFHorEyU4rF
ofZxZuWfB9oWbJJQeZTIiKt1pQnkvAH/MYuruAZixnjxfv6ruw6L5BwWTOd6
TLIHWLDRA4gufhaN4riYvZtT9Q1XnyHNLvU3E/KRx+16d27gugs+YUtZFbHJ
mE2vNuGr2kXCE4K1JrZ4GjlDyoAAypIlW7mUCijch1dTHpIstiyRHoQoG+FD
N7oNg64Tm2hXXDwDEiZjM0j3JhFVibxr3JvZ6tHfbB/WexxTnTCyrKR8lWPq
n180FcYLkMX1PHY/E8biGm7xD5ltsTNnUs7gxHXKZWCBDaxp8l5siBvxRvKP
XNQm8d4rr5DAXYB/x6waWtCEvEeM6jtjPTtxbgetA4Wz2u2Wn2gApqQ2YBN9
fyRbbSP8bWjraPc70lt6hUY/rqBw3QcSxs60ALXNeA1hvoYq2gKtQ5kgOJlP
KrjyKCwc/JEm/5JT8HaWaOII8BWTgft2um+m8+OgqKFiBFu8lqluqkxKmBVt
JSoNXIYRRIRW9fh8GS5G4fYl2TXDLiX3UbvS07q5DhQtQfHS/kbGV9Lc6yO/
E6yfLHPKRasz99U8h88wgzEXzVClvxALWAtEMoFyv898A/PRS7OgDITVBHog
L15WaYJcu3yA4P9+q3IwZl6JPw6pVG9XZfo5ETu9fas+R2s2aFYxydN/yOKd
7STTHPX9tpg9YeySG/hOOIeSNkYPag11soXNMdqz9crx7pd9LNVYM6cherME
OSbTS6T0TH0DVX/GhrdU3FzSirHbVUiwf5lpnXASKlNbYsh3rca5I8NZEbQY
FHzHYn8SAhiaxSGuo6STfckvBO0CA67Ffdzx/7+lbzBAesaYulw2ShB30dKL
KaJPFGIFaoWbmmZhFFtF+nkIl9UiZI1GZxfYcwEjHz7xDlvqf1cco9ydvPJ9
VFiFFyzJLs/xmqhqv9KhVtU+Y2DRYnmM5y8o8ze83Qlc+1fTrgZVLS3L1buI
pVBxd/mLh5SCmm5NN6ZllleprsJC7iy5303bKogB/bZvBEws1ftJYL6jSYhO
HO1QTqkSdHN/NB0J00w425unP4fnIEHVci9YT3R77m5NIoZUcuRUl+35COln
83ymrszEcfiD5yPfmpJHfBs5XHg9jbnfhomxyF472uQ6ecr3tT3hauF80W2s
lLwac4I8AFFywVhYy1zBjBuNbN+CUzS1wz1x2lEWLBmmYvdFavOPfRRWMPq2
0M1SnxWZHHhLJe7CEq9B8gKY3C2FThXmtJmlapzDTgJTrtnJwH7I4oJQ3vX6
DTnamKY4xD2GZoJ4bC7ycLJi2eSzYxPsadISEzaH6iP8R+3lPR20T2oEh1wP
uWRYYy1sqdsQvuERjZVvZvkMV21DoueUOLeFHAFMv1bYXrQusL/6Wh43N800
Cu3i/PAqf8rPtaPOriW+zX5F0sDonzZ895avIeqBLvewmdk9kPVxPZDsQjpe
4GpFxwL/ul9IuUN96aoGfvLXsKLz7aJ9qEU43wj9DjdEFPFSgg7gFqkuBq0B
K+Tq5CHBytLwR9sS/zxgERL1teThXewQEPwqx1lh8nDsJlPAT6nR0UkXgX+X
j4DRYPlvOnd2y8HwmP/23gvlD30oCDbLXqA10utcPa5qWqv7pQVWI/cP1oBU
sn3OUiqSV/pXMjh2XVskAcQyJYW/OukABnuurwxlFSahZn72FiPVZPviFYfW
/gSm3XQLccO74bL/vPuj3NH6O1M8HyttLP3iv49prm65e20UBrb8wZ3dHJsS
jsu+L7vpRuO8Zhb9oQqbIAxQNct++LbkygrQBxYATWY76rL/M8YVvqyPT2s9
0pkF4vHItD2dcG75ttuYkdNpJeUDuKyhjcbrE6ddiMaxT0DNpWjj5LqQP3T6
xjqZsdoD75TCsnKIgQCPcjooE1a+BoiDKwW3OvuBRS4nwrd59RfL7OcVZnSR
0BRh1rrOLn8Q4AO1FLnt6Li+TdXvAT7HcPFjOXY4hgI6kjsYSUxG6Xx+Oyzw
UaSw8jKlMgJnCzYx02ICMRPFSHzJhmNvHXm99ka88ZvFJbtyfENscsPnSYOc
jiRgubMe1U+gyx5w8/OvJhUFn+d5MQHtogEeNHZ5YRc4S3HmwyB8AG2c8im7
684y/4PEP0EeE8yg4egkACaCSvfih8QpcNGBEIyinlyzxaZ7EwDWj0PonqWF
aG6/ienb2gnf3ZEltdYkjKngdXQLbLjKoV/s1IZhfx8hxJ10SRcsGTNox42r
eh5Em5pTOjmsdO5cbsA88S6ardT2+ZSI2V8xr3KQSVtjXH13dV+b4yeAds0J
qWSBJKkp30F+PNxbyN9m+s7Uq6A0om4lKsP/SCraAwAfhDDP1Q5BaxPSYMfj
udwTg+Ne7p7JQNeIIhdx05KDPbLHfC1H+UUQnp3ekmjadeQhejKD466yi/XM
lNTcph4kmpyn3GRi2PYEmhbx4a9M4knb8RfbthUyFT5/U+H/OYd0zRBHtXlq
595FQrgreKN2mzRI4XpWBTUogpNiCojNkilolCrjRhD69RPsW0qJP7MQY+jz
ct4Q7YJtdpFnVQM0kismiMV/vyNZkeSFIKtKt+de5BQSYiw2YggNuq2MqcOH
ycEQansv3BOLAibmfcywYqsloXRyff6kSnopCsP0rd+jIjNEMjhknT/hpVVQ
VXUs4MDDldy5iFFZkF02wYKDX6pzS0iEqajZ7RLUEUaVFXlnIn6Z2nRgrMxa
/hXRSxpJ7SqppUqbEtp5xdSozkxJP35rUSbN8ZBFw76n6J94KQqOeGWeg2/I
BcfpABwPuTJiOhKs+dEXXBwJ0MP1tVyjrqPgC+ZUz5tDk1+vW6cBU7fmUHlr
kkaNOV3QMNcD1xDvNmMeNXAivjEy6/yV22Bce3Nif10SOpJ+b7ViXWwI/o5n
0vVZsHpqy+29k6rmYFD9xsmPtbUhPQcEhK2LUOZHNG1f84uZ8sxfR+dzMHBV
dFEa/Xi4Mnx6TtWhqhcizqCnhhxLjN4tcBi7i/6L67fEBAADyp3RnGRNdMUO
37rTyuvObKMet82OJr9l/T4rTy8v+Qq1m1fztZdIaVGh7sAQPbIuqWZTwT7Y
i243IxAmwqrRGYtHbI6vnctz69ksXmVFqanH78SmJx5lq+giKMuhlPFwCwOX
8ao7MLl5P/eXLd79Ls7v5A8TJ60VJXwsMW7TIuh+MjBeNkr182Ri2o2Vdk2N
BR2u3YnNp9YwRtCknsH76OU63NKuoCcwzPJZay5fHe4dMsNrkLMaES0jMj9x
vSvOSGdx35+WYuxjN4LNoWfjrXhqRKjeMdkrJO09p7zNPz+4IROEZ3+AJk74
Ogq+D9nBUJP0cscFwdGGm8KV3bbohR0nWEmffi01zy6vbnzRmeRBg6syVwAP
XipUQ7HhbipXVfkegUtNeiDMo17AJE/KmNG7iMzkH8N+GKyi9oL3bMWVPEyh
hThb0zwsvw2WnNftDU6l2swoyNBllPWguiRXUM3oyaqPZanvbwZrOevrtOPG
5vvgjRXEly8J5qGWTsNzC59Ahqf5KI/Ydy2aRW+rKibi/HEgv/v5AI/8O3Pm
yNpr24TYDGxmOU65Hi/+M15H73IIk3Awua1ShOWmkq6ZGb+0KLrXfQNOV05w
OLqWWk77AUdL8v7NWcERI2zRd62y1SLPlRFQMB9GSv09AbCvty04MkGrC1CW
TD3Nl+lkBKhs2kCh8W7WI2Hc+Zcn+V6Je1P8pcya1qXfMorwOe+30BQxwmPl
N0BmuGcOFEhvg89CxB91ikr5Whgxa18AtgSKSp1ukpq4UfEA5TdcqGO9dAB9
FTSUzj8Ko2sS/6cFc21daMnjFXmSnHdgzadFPdST1Bv9a7syuzqZ5N74Cubi
UItmFh47tkai2RpbLY+8UUObuSaJhOLnosws4R0q7YUr2wmDlJavmxazG5MK
Ntnjbv6el3yI4YArejhgtLUR6MgUJ66Jo9W+xY+N59tx0QTmi3p/ofGwj5mv
bEc3F6bWp4LvuKr8HjZI+uk5xrJAEvYOfQLZofJkcZCo4fVPFJ4AzHC+2Ek/
f8GksN7twU3VzK3Ue32r3vCkT5XZ5P0kDp7TPhbihNYs/ZNKJnATv5CTVF5v
s7PQPAjz9kYIO6gJaIj3V2bqlWHc3pBOugSNCYb4J2DzPGL57sqK53pJ3+Pq
L84TZBT3qFoj3gP0dQDvkCD3w/7+r/x7AEZur0R7ui5DMjbAsHlqX2yWgcHf
h2++PpBbOd99ABNhgNw3OLBPRwpcTny4KUYh+wGLX51Xt/wH7dQ9J4/Q0VYR
/41B+DzLcOgb+YYhCGA1QgWz7k5m4arkLRQHpos9HMIWQWDbW1RJaG7hueQc
82tEpZOqKXBYW/esdzSM1i05yl1rfX4YAtJ1BzczaKgB/WEzm2uHrp2AzGU4
VMxQyFm51QG36txs/tseWGGEh4RmMQDZxep/hDJyieJoifcLP87a413CCMLp
h5LyoRL+tgfoY8YtiopMrMlfLXh8cdm6vRva0cCuLxRHr0qcBPqR/TFGwib1
IPrPXYhUO64vAep8oizvjeHZNA5YrqyXx2ML2ukAlUWTSnK8sZM3O10hi+6x
hqgm8RlS6urj3E6sEOjzWA6NHjBinGg8X6VKcTn98ErZPqhrr5GIGvSLnOWe
CU+6XmCJGFi6VqBRUdjWPh105zOXL99GH4YZVHfydCC9v7BG5BtzL2hV4tl+
I34ympIE4xjdqSO8MbTxkfPSrbl3eILNKETis9HCRcp5thwV5VOx9E/Kb9Od
N8/RY17KOLgheR891u/w0DFA9feBQ+28hPCVzvuTVVwj+le+kUPhWcdW+dCL
F5ubut6cgm+KOVpqIuereVuN0iB5JLf8P+oK7h8NcYgtpxKyTPnDizC3tcMn
ITUiATlja0JE9X7Ttnt+pTXDlPitRKwXbflUfyIffa2LMnguEK8c6wHi7qyM
OpaaU3tIVY7NWjuAeyuRWNehCibXPYDG7qvsdl/Om8V10hKZ9DN/m1ZPhSLt
e4d9cY0Jk1STeZJv9R82hogtUYHWBrycls5kx5Zx2cRv3PEY6htFgUVBnAyo
6nGMUNyJGdfvfQuHBoynRI7JRytz2RsfqvAmyUDA+3LKj+TPLvWoLMnQZWMM
6Wo8OucFUfjbiyMSzklU0p1nrC0uOqelwRyDWh3Mt5UPNr7FE/Yxbq8/GRM+
/P+JYpeCjsuRTL9M7v5iNw3NvbTqepFKBKRFX07cFkqpOvkupvnNtNA6XI8w
loG4JE9rIAjyqI5e2Ofbov4C5YeBYF3cMGKIrQxvNbuGk7DdWKR1MVgvXKm2
VGfsr4ZsDamyq8c9te5p3YEoC4O9k9QJJTxbHn/MJD8/mvyAh2IJFXjk9EH+
Ci7DZwRre6juXM+cT8LECqD+yzIgTVy9Sl7Y2CBZHOXw2AkeZ4cRHuszB3e5
9OKM5EJYOIK2VEscjC0I/+K2AeekQgeaN9WJ3+gPPbZzRsewW2TdMu6POlp1
9CpxupOgE2aEkkbId3nAeE4O+SmyuA6x5KR/wHZRT2VLd6MJKM6iXZy5GyoC
HMnYmHYXSa98t+mspLtDxOnkrCPfgY833AUKlq7JNtDvsfXRetQSq73Azsl/
qDSleWXtPNuWrlZZ9NjQzfIaQZrMoLWR/spTKkrM3w/FpQKtTCtcgeK/PlIn
of1tUxWzXvHeiSbcWp96keS6o/UInSDzpfQL2K+qOR6i809p1ENnM5ZpCA5I
XxLZ1tckeSiiHUYEbQoLAxxIZvuzqEjRW86wMkvJf8RLxKhBPdRtuHpupIJG
rdRIIWouXgS3fI3vG6eGdfD4gEss8FUVHk2LwtNgK1qn8bVxy/VQ+Y75AyL9
4kjJMw2yjaotSmi7hsuCrP/MmhZpTwiydGXbJzt6DRIn7m2HpNV8TmeRCuOd
eARAsF63l1sdrdUnutVxTpPnVl9jD5cUgpz7Iy2/38KLen1LdX5VmkT3vSBO
osDNPhzKL1kyeOQyUH7lOb13zGuOtULbJn8ebUW+jDZnP7OFzP70LLfNPElc
a/ukEucXQ/Yhzket69Sq7SgZQu7DWASUDFa7md4viOV2OsO6XQ==

`pragma protect end_protected
