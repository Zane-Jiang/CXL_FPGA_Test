`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
sSQLH7OWK2skeCPOxAddK4hxpUoWfvP6RF70QsXNu5NP/IBlSId75YlrsAgEjRV/
QMUf2VTV1GtjZqln+BdvrPUpW8wXoWvy1v4kBxUvydxXZnGOk1WRGEKcbJbdOvq6
JkjU6hkmg5qv/D+DZDTUAdUS+B2O+r9ZbreCQaEODRI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4096), data_block
71Y3Hvsk1jm59o1AdTklAdD6IEFVVFDLHGkMtmv8wibAXiXDOXJEbYIv/hGfmZ+X
wiz5pPwiwA34oNjfE2uUsU4hbqwTt+keLjaYUE3UC03n/6/8WiLYDFoi6+0ye6BY
00pURT9i+fteauc8qghsUWeQEDBMgeNRvuaKGmUz778ZPXZ0NwHKZlMdiYDY7Kf1
7OjZJ/N4JK86WwsOm4i7AJayI5wcmcAPD+yE69S1Ro7rYAtdLnnVMvd61U82LNDB
SddMB9wcutshrIHVcsMy1gnNfLyIWFDG23h2HitkoVc/nQDL6NotIpwL3WaPd5U7
quMoXMb8d4VDlRndggtrIeU1bAceTQ7CHZOAtNKJS/fdt6wGDm1H6bSwjtA3s+2w
EdW/qurfzcyIujFMtS9c88mgggD7s9ZsKCAfIQWVVGFZ+qHJDo1X829sSe1hUsod
tHsKi1wr6aCIt+QBgkyCEX3zJwufJIlYm+E00QIXwz8k78XkV1H3jmn82G/BaBl1
UMFiLGjVoPt4W5OVfH/9QKdJNeNlSwzbLCPXQ+Sh0p5H5h2fcDxZxpwalrIjFW9Y
1wK2yNiZtSG9wRcPVYAwBf4GuiPhU1tp042/Z8iujliTk96tOjpJBXMEfIPdZC4v
a8jSSvh7IsKWadZusDTgIhqgyGsA8yJaNc3YRrKsh6Mce3U85KzqR8/TlnNcQqkU
dHqGaEihq1QIhrWTvdTb7TPcsy+gO5rUw4tbnmE/bLspxfnNmllZkVPc0px8yJTM
Bnw4LJR9w0qDjp8dISXnB56h0MwFF7VIccq8+hv6cCJGEYaRSLUD8V+1laDSyaRF
6tLveDe/UNnKyvaPRZmKFkzdeFLupx0XLCxKyxmJMcVF2UZVcrhe0kKdbowvkUmU
uXwf2JM70t27LOi/SiF20ll2LqJ0e1emxBA+XgP1zN8HiQDbylgUdIdykUvOzknw
S3LjUkJ9eNONIaPFjtPm1xgUvVlmQjB3Dv+vIgFOPPLTjt+7rFq4nwZgC3TsokdG
1RxefM0tfg/SGrWI9wQlSlEiRX4/Htf/xCluritnhBoPiEAiQhgu8nu9W/McV5dz
jwmJubQPLw97U/ISa8weR1bXVnEcnx6sHipHSiIYBzbJMVP/KNhAhJs9AFrSPd44
qY6tHtZK4dVlbrhTBCDIRS2XkTmFDamk6v7dMaXmAoNZ1daqhY0RVkzGA4Yj//eM
eXkj7cAS3x2+HO56PYQ+EodkfzIjDvEZEg2I7TNlCkDuJBbzrtGXbhPsCRwirrAG
ICE1isBHAdDUBhxyG+MW4BotMuuza6h0qJLd1y+d/bhEESfouRhT/4MUafs26vZL
6h4bmKka0aD1KCc7uff3CERcwCQw45siPNPSZmzw4feqa4x+x+C06BkvfAeWaeXH
ikaiRIeI0S51YisLauU87CA3FZp0D9/2YQVEj5sKMwnRA0DKXJx0G2Dpokkf/yqb
ghYvLKdvsFOFF229dSMD3ah7NsKWlx9TPf6haZaGVrB3sRj8z4aegK4VJYp6gMK7
5sUv+Um0Yk2Ip9Qg9+7Pcxm4Mk8h7116EOePJ2Sr7IJbRPWAHgY5iPZmRCu2KTK7
4rbU4AG/NBE6zQWhCJNPLkmbRFkbfpcqjxJFr/JM22Jh4qGWjGiHb7wsvdObRt+0
+wbB03j5f/rXGLr3Hn7jENxQflPszq7tjWqKWrWkrvWgpfghWjmPf0sdiF2kX8hw
HbHWpopYQSJg8X6IJxD3f0aOV4IYUKKqDlXXHrNjzXl7QzIX+ebEmkJsPtjB9N+y
IwLyh8lzk72QOg7LlAELCNDrAhUTj5Ti53vVOulpSHz17w0Y+61nZHshmF1zmopj
R8IFc3PTc5YwCK4k+2mjuaew1+ZCGqxT96eLOulDbFUEa79ct7ZriLIueMv90JRm
GxxAPZTxY5tb+IlEEe60W0X/c5tGTEihoOhku79SKqc0VtN0UahoIA2E2rleMR/R
eBxh17L6bmoAHqAhndXWnY3Z0WZGD0q5GBnSdDZ83r/8woD7rnS/ShzDs6MRftOH
7oujtywLOQoDAam+H9BuQtGdMbu0fZzp/Fiz6/h6E/GICicIrGHggaBY2Lsn4ieh
RzWnYTQJkbLM241cDGqJM5Wh9ZqXSe0NdVGXwebzCaH5mllTNPUaAG+nJH83IIVf
n3E5Ua/UTqz0rYARU3IQcuZnFLP7RxBDoOpJpF1RYByk9Zj7SRWqV/L6NiSHaO6u
+GA6l6Ln8NITGLNX8WPPzfLW34o6b/BLVij0EG7XUuvOO1sgFBfyFSpP97d2//Hl
vG2hTHik5u6pwcw7lMg8ZBQjSmDxzzYR8+hWhiVOY9nNBC/VRJkAwbSuKfbyd1F/
hMGhJ6ZpBLTToSC40XVmCpBTOpfptKZmEdX2HfxECUdSEh9FldIF0A+MY4qA13UJ
Ay1cN+6/suihaOX3ThZ70HRbbxeYUu0seNUXzjOxYWoYDUihWzbgbQp0aGp9In8u
EFYHU3Hzl4p294KogHL/uNAtEXLwkoYzHEBuM/sO4dY6E2iZHwgEAVW8vWoIguNv
cznXu7mY7vRvaTleC24b40oK/4kCXylYXHhFIzjk7jPw5S2GjD2bT+rzZOxo5syN
hgiel+9vhlDgu81Sawk7HTOVfwTw4lRQYxp/Y8CciQVb3j6zuXVqGyi0onIKbGoR
YPpUyHVZHZb5p60lhlI78yuScliUSpktqWRh1c9KXmtV3UADcato/szH7A88ibQd
xOjmRDYt3YPGO2qOk2vfg206YvSgFQsWK2kAxbG7owQaca/ZWNaL4mFTG6tb982q
fmQ0qrjoqN7zwHe2TOp2I4adKpaDHVhqXACM22ptkXpixhsGnQ02/AWHq+9b7g89
c4aasqNflqjLbHKj4gFYU8xVUaJCalshaxSWNTNisYOKYTT40Dzz2FqSEA9hn/Jz
0O23oByYfTnioPVEfmV0N1/E5XX+1oZRrR+O21geiLFhGe/9NofHYQeVU9StCzCb
l1rtkjizFSJytVzqhVIMhQlT5uh3316NyADzrepFHZ7hwsA3mZLWTDCwIYkgZO2b
gU/n/VTL/VtJkDGEJjwHGX0Cc73Ek/vBi9LMFEIEJ1caFfdsqoEoQUNRZ0630Otb
YCj7OwHRAImNdGTMKqwhU81IoM2x/HIKi2Iv/NQsvfDJDJS/bufeD3Vj6M4h3rrx
crXEeLIduSS1e38em9xYTPPRnLb0aB/IyM9gdZPh2+KzmxA9kqoMNcs1I/KbXOwL
xALdiZEuuEAn4SYc4mqVs84LffLLfezBZuBL7Jh9vxhtm8xhyPVV6UkyQZjQESqQ
70eiAIewUvxTUTm0jNWpuZqtDSOG6h5r4PPQqooZ9QL2QXNtIrKZu9ZKqiZ20Ori
Ei0yov9Dktym4m9IOZK+UVwehkVlOhBaQ2M3TRdxUhoB8G4yQYRwkDXbwO2we8UI
BclqPB1ruHCMpucqSToY7Gl0lW8Bo9mUK0jcSgx5ksYrxm/uxdUcUlJ4VntZCHPO
gOoFGyPAPZ/sm4xEkKiYz8uqGyBKN+WAkymYpj93kp45G+sgfxLj5R+9SQfIa2tI
K2Cro/snR7Z652t2KSukAkHfEzIQJ/XkKpVkYcy8mPM7FwqnqiTgGXQ8F4Y1uSRk
748lgw39b4++RGGYeF7cu1g4gVqlGsQTuvRsdyMnFdfZM/PJ1jMc7SWj8WPyhnP1
FLeqe51g+GsjNUHOO1+39d2fyq+/IZaLL7ReH++Jx6+IGVar7QVFk4p6nTtrq7Sl
3f9lXehC0x/skpC7MWhY6gnzpMdhgcnJEYkTw1tJ63cwtYuYJgPZF4yWcryHlt3r
D31Fl94vDtzOWkO41iWz0DKVbUPh87U1dJZZ1D62RHoEXaTNUg8FfgblfwR1KkM6
JdIWTLBtjlh6IyCz1X6l0dxwUGSv0ZQ+J4wEIjKwnKN8NgryKVOfaR/XV8+zSeZZ
U+94sgIBpDSmlpIZl3bx37bj2OVAOrhJdKAtCHsa0n2Ed9r72dhwZu54Qw/NbRqf
6pP4zL00wbyvk3qqUKX/0cuRUFZsKF8dM5VUmrzBUaBavTO3S1JIfIZSzVPNny6x
v3Tpno9l5o7Bi/OfU4/HTeDdpZ/hCtkS9TmWkH5dxT2t/e2b8OHS64SQGx366/Zz
CHgmjf3cTxjrHIomgY/GAOQq0XeyRTQM2Hv6vtWFn1nnxafJ3hbqaxJyL922QJQR
4p3t/8R1D+eNNbBan6kOHCF3+lX2/MKI+GDQEueQOu/gSQz92GYn9u6ICGHmkSnT
CoJmOWI9pIBO+5Psn+N8TPp1RgSHhX7hTp2OLnNWPOQEUx5PDHb8O6goKyjBDKPQ
seyW/Adl1850/inBIJAc82rQhMQdTCMfF+OXNOm+2RbUS7Hlw9jfBnWqubWo3Mnd
8A6IJL+qOWq36vmvX1KcdMzh/OaxPOduAvABp/GMgeuVORJwA6MXlSSOJysmBOiI
RAXr+ruZdw9qx23aC8QWXAQRWoA1pM/z+oo+VtgKF1NxJR9uXed8jCjZN+D8207T
CkLvn4OVDvUb6+RKWWd7+p0Xz40zdOiKN6xPNmVTFR7rOsVV9PCg1m6GwH8z6qd7
MigwB68tZfHtp+tM0ehmX3K/kOSCjjxcLO1nYDccDA22Xau6vHcKMl7Ft9Tfwr+I
n8EvcoOkdCwr3gZ5u7WiApjb30wj3vSubgKj49vlkCUfmRe6SWqHM3/fKPT0yfqe
1s2YlBTnBHG4ad7rp9lsDnmaPxQTjrzBsSycx0GpNC1Qqj6x4dLajTOdSfyRjWsS
CfVTox7Ey2hZKbJtMWHBq/DmiIVUKUP3JOP+07EYr586dwalxSCNizXP5uIIVH4k
YZqfvmqElwI/w906k/JW3enU4+rd+hB3zAauf+UHZA6iURyiphTC6o5HNPf17s5Y
KjH7Zm4guMbAipWq7SWAKjjFNEl+Rf1VzJs1k1tr7gZWEX5Qg192ARW2d4pfWK9X
jRhmpQelw1cHlSIvm98GekPL/+lDN/HrBGtZMRXjY9cN0t4UGTI7IqQjvKhgtAP4
aHQpuhG88crM82v3ojIlpioz8mU6SIC9xJAse9nWmOwM8QPUvqy6NQVjLNCW6jQl
959DCE+UCxJWoMyOmScws5pgcwFplBH2+BVaQq+JFK5HDhkKL2Hg+ntAOcHD2Pni
+k00JBXGW/fVox96hIWmRvmjKW+dYLkplNZgibjMTPpSEoqyC6Xwwf7C3olGEv4E
T7SWIQBOqmvzXWv8nZ1vQrfP7PF/gInLhPBKKKnL9TD1rF0i8OS5Oy0kD0H8fNOo
EuVpfcBMnFDIn/WIeZ5kWVH+ETeze019BLfmk5CXb3XIB/3CTHQrKnTnwlENNnYo
8mpVCqAp+b8xtcIUP0sf8JtrTgR7wJ0ejpgmzent/bl67P/9T0aj0W+MD0T468MR
MAc5eNsYfs9OQISY5haxvQ==
`pragma protect end_protected
