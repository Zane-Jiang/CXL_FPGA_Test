// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OE7p/vm2Kx+WSLfzzJYGlnQu7hI2jdZ7rVVs1tzcbDxAQJGSGDsrFMXOhm5C
GD2eYlnVi/W2V6mxY6gpWfL7DtmW0wGV1qgdsVA6hi8ALuJX2+eWkTCHYCWK
TIAerl1bf0AllFvYK89Lzn9RoqRN9XQYFewRvarU/K0WNOhYKh2YJvJWEsEH
7n7016eVnUoY+2Aa8tL3pzG8WLJOvNvsZenkeogFm3IsBWBT0soGCbqK7pAF
hM5XOHMRF/Mi5Jc3hRWMobqW+V1Wu0ABKfUMAyl8UvmsKe+2fxej/0eypqMY
GogQcSu2YyEER2HYI7ZU+UflEr88C0TmA3etR6gC3Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y2burWwIYYolJEgSaoeTui4Dvy2/2T0qtXwjBdWNQFhkXvsRRrS4OEeDQscR
HXxpIH2HDZbBMwlOyXJE4CGXDWIrp84ulZ9egBotaEW62kxAprM42DysZZZS
Xl/nBAvvnZRHcZW000iLqnANDECkel/o0IO/sNg9GigXQiwPlWIlbuXJhD+F
55G179go4Ur1fDUdQusOCzb6HLUVBi/977yObfQ+p1bR2GpvdrP32CDZZZMr
lC+94dc5NaW6DbPCp8rT5uFQy7q+Ey3dpzjTvzhfEsdUmW901ImwR22eZoTK
xMzrahj1Pk7UKZbQFAWek9ycaxR5+2qZHy0QwU3lmA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A4VAZDzYEcQjNFbmnUTmUO2oY4122UjmiMa+GFzPIUnSN8OCWe9aESFb6Dxn
2VObjHv8ftQaJQ3KFzH6C7XHEvQb2gGpRIL72p9X5bCff8zjCi16y/ep0zmz
IdfWeFzEAO3Nq/xbXiOYVfLWJl8xPf4G5pd71xGvFTLDK80ExR0Uzvy6h0RG
f+y+OmTBIr/MZ4QOu2Fx0bXmeJaA0Dslh259JdYagapKb5k8LvW8aqJVmHTq
/9uiz9d2k3wJcZFmnWPlBW+YswHHFpD3glAL4ZVZ+bk+gZXjSREbjwFpKzPv
pi/oJwMZGyJ4mZouLYh2nM5Y++g9ZQiwTsvZ3TElRw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Qo8dM4vmbnF7tfcS2shkJoOPPGnW0KGQuWXa4msAyvecCgw7gE8HUelz9gfg
yGUo+KkR5tzZr51frGNtsaLHHAV/99yXmClHXVwokmFAoIq+sSOxAOTghtC9
eH52g0y/ChtOMalb5NoeNXnCSnK0A5xU67bj9W6SoXqkmmhZuGE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pJmQ0DDK7H+qm7Sd5snjkavrAzqY2v7JG/A7SHDxVyeYI4UW5zJp/vjye2bI
Il4zcs2VHS9DfPvi8wrKy/qAq/gM4rTr0WZtIDUBtm8nVDvMsYUczAgH0OJl
AQcD+PJNfsjylkHBbnUG00VMbFDpcStNa7ACNQ3Os9BPaSeow4DU50i+viqF
zauG7fEmeZYrlzXftsZb+COiynn8qFK2vgchA2XiKNL1slZt9o3VAuPP1sbK
KECKMVGn9dOXO6GZ6ygQbpQTgSqqeMPaRcUN2J3qNyzetExUZRQJP1lz0ifE
0jij8/1GD6dOh1P6PG+iqG59TpY1b9MeOztWqp4bUkEdXcz4tImVEfw+JsDj
e7r//jz043fJSAVtJAlZFkokx3MQBEvx5dJnGQ5Jj1syO0p5hhQOshjSg49/
j94UEwzzicuRP5kqmLMjMKTKenQpJq1radA+LlaftRFePy/+mBzXyNvYogwl
zAY7AJvmGHnkKOweiXSnHMGzc5utHHQt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IVzXOuw6rRP/xXegDgbYm5+1SMXuX+QMTmgj/zMbQnYAcps//g90DhDAG6CY
4SiCALjDIfEil71sCFPGGbjWqS9xuRa67GZQfoIvPdIy4ooj9c7w8hLmCtLu
gieBFX3c/PRNqCt1uu+u39IQ3dINezwZot9vWGz/M6C7gaiIO08=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aUtlcWLOmdRnhARxrN9nVgBpGjkvHDVkPB4Zf//mB9fukoHR6jW6fkOeSWfP
Ac/4PgkAVQj5SSpuYZ8+eDXj/6l8oVlKcOzYJBfB2/QiKq7qylOYRA/mHuwj
sbSTNcVaWQGKRr0MZB53osX/pz/sffoe6uhDRxqi6jvQhoAJMWE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 37152)
`pragma protect data_block
JUKC3JL7W4ofc0IcLhN33JUUgxdQifAQaqym/MQhhgBnw/XxB330Fd8MdeBb
tMtYvhA5XPu8Yb1s/jgocjrg02JT5fCHlN3cxS4eQBVnmDdkJDW78h5kccn4
gCDKSFdyAcznbJLJIvDI3fZqFFgQOaefd6LPe97VVilVmEpg+AoozNq6YdE+
6bYggaKJWFgpVnUfJH/Xqrmr5khhmzah7CR4bdKA9T/AIIWQrJAFJRuEodVx
I2KoeJgmruaNjIVO0CMTAVKeefiQNf62x7/dF//pnA47BSg82wRbJfoJIEvb
R9HkCN2kZGTYWjcsC9KBTFOYY17Ww0at9wurrV7PMeYADpy1iOLAVXJpaRrq
+1SDY7xJYy/nAZDdzriRuAVaZRKARtZrrdC1wB7mff2tgtxf/hPsuxUPL5NC
Hmyl8ZAlWL6VPekr0uYVNFmWNv16hQgQx34xVyU3y9PdrOGhQamUuD1c3sin
h9Fdhjna4X5ebQwsANiaIz9Uz3RPpELVfRaKfkAR3ya1iO1u6nqpbF+C8hdA
cZnycK8zAu3+HPl4psditSeu2gBDvHZDdeo7CF8ho/hHM0kE9tlu2Og+dG9o
uTiQCDh2yDEj1cLkEERmGX5kUvI8+DTir0jROGF2SY4ieUPRMkEuxXE8V6M0
eevuPR3r4W50rcEvYVmCvaj5Q9eRO9cCAUDMhQA+TUcdhvnLOiMZoOVTIKi3
NNidoQgQ/N0Lv+NrfYAjF3zk57bbczPHIbpao0hRa5MyfPrlZcr17Hia1AXM
s7s4X8z7+dBge4m3MxPHBEK0+psFtKiAq/52CUsGcM6FhYYBK6xCK/HE6dvR
6ytJpR1V9XXikY9jYvOZ2zs8bVIywIvvwBr4WDcy5LBcNHBm6ETwB3qCq2T6
OPLopxTONBGZg8gjs98+muAjYIRV7kwqLzhbEJ2DGsqoCZ+p2Dea/r0nc9f0
mt9M4z7runjOjrf4pDI7TQXj6OXyxJHtaEfOLQpdZp+Ma1r/NR4FMOTkR42J
njnnl/RPJRw2Q2Ex1RP8DFkhsLCgApg/hQp/8EkkJrBtWq4BFf55SWh2WR0H
aJ7p9jGP47wvjmU5dTSCX/Wf67zuSjQ4w0iCBnOrX3AZ7dZKEWiQN/MZ/iTq
/u3Vrlze49+t+tT0Hn8rxDQ+L92zgxp3GgIcZSEzdtiUkwsiCKzaJbD+emJ4
G8AIT1acq4eACy2QfLwOg1W0opUmYnS90lz06QMT2600NVxm1pfZhSOuTmfX
q7q8uqp7QcU1uCnlKgreZetf9/8/2Ld88fEqQqbDAxJS4U9I/gQ6nxItI+nS
AUeWuqMTSCmxhiQQHVRQ/OMvVUJfjtw6hKk40iw4gERYK/YRjxIoYIMGviAR
Egw8mpp0KeqCGdt31ltZ705WHAcF4QA5Q5qpV5GZDQD8yw8lLdYJ9ikWt/hS
vphwBCIMNIjz9vkMTdqrznDyc3nOotApI99GMrkPlNsTw8L4nYLKAyVGxpSB
fMYq10Lr5Bfy0pqm83xYKpUpKDJ8LPzU/VH17qiGGvBlss2/WZDHOGlIrX8u
ptLCZiQIDuINmMqzXEB1mBmNgf36FO/558qLlaPgFOxEqZkjXejyTfbZRUQh
yMeG8mf8wTadKwTxDEcj2buQXm0iB3tryGHVny1D7Sto/Nvlg4AMpP8QNUIK
CU1krZpQGAGbe7nTuFaJxPPjxNG/I1c/qgD/rJGQ9f6k0NLwL3/wHFd+KMag
FpvhtB8axI4Ce5URGtq/slnKDEIxX60/P8kxtkQbHZM9+UtYxQkJcr5FIxrc
vh21pBNV7LhGon5kVjFRSn10wIBX61jNpm1AlQJFaglRwA+Nq9Ydy5Wr7KCz
+afhDRmHoK9QRY4CesoVf5q+Nx1ytMlj7QzmLvWVXNKLW+1Il6BlNRSsRfVp
QGZA2B0Ny0zUqk/eXShIQdGL8eUTtM8n7/CAAeGzRS+wjL9QdqHwf4t+xKB6
H81aqiBSGIodlFCPDgr2CK0otgqpiN2SzZHYpYcssdtSy2NT+Bwb7pEWOTkJ
NsyrCTbyGznMgNnEylmECKlBZ/VfoXd7+pctLvlDncMbK5r2FaGgFqvtSXSo
6wYpHa6Lqg61GZw5vsTlAoz391VwqfrPZTmELC4+fIShKz0/FRW0o77wJl5k
X1+9iWs9jVg8L2L4OvcygjsHWjuYXfsS9+pX3BtEubnGDni/6wY8Ou7ncUcf
gnnN3bDy7EUQVLtlNgCUVWhOBtifklRIKNJ75OdDjn5jVgtIbb/Q0M5yzEIM
QcviF903HnYS2IMPlwxlSiXWOEoM8iFx4qvVhOstXTS32d6iu3MPHKXysxB8
FXHhUeb6qFWXMJfA7lDcwB93eQ1eigiOka1bcKdUr3ojQcBL30qabswP1tiK
r1XJP7XD/nLOdIiJ9AF7lG0Ce3PMwfFb7tzKpItQk9FyZHPFgpz1FXqLObCt
1JpDitenolAUnh4iHLMjC94ayrJ7Hl9dXHQrEpJNAgolpBGKxb2SMOKkw2Vo
PJYVxJCMXq3+pag57+X8yOXjumFMd9Z4ncOAhNhZ4g+/KWMVGBTUmAfZytbk
zEuCLkliUEDXNJ4NLO7Rxq2c0p5SKwLwLfqsoUUdP+yiYrXZSU9Z7jo2JP6g
2rmQml1J6oaH0JGV1PPt1sSD3SOK7gLkNLV19K9ah0PRVGpMNSSVTVxkP6zX
Ftm7fdPyyhzJSfvyBBDG7VkMnj5IsMNrpiM9IEF2UbHjiNNFB+Bvhh5BlSrE
LYFj29CB11lqerLN1NhSwXqbDptnrR+/p8jXQ94z5ElA7sc/1Kr/PtNQjefN
w+nFRWXU9pWstCADE7+1mZwWVC0+Eb6Ek2o9Ql1hKx3GXyxNLCaKe/m85DUb
yzJSiN7LA909k/KQJ6C90DVeyQyIe+6D5ch//WN6E2163NJzibAnaFAIS/qk
1wNCKAn9fGHdBf+SfKiT4nLmUruG7yAQujlfMGa50xf2YTg2iazmeYZ2N1CE
p+HWk8kqqb28nUtxOyulCFqX35Pw6gYYJbuJsUY6t9Zs2b8UH82k8RAqyK9B
yGSWXzdePGfhmibskXkdbczjplBtqEkEfBVevz9lt87V7WrEbyGB8ei5ljVa
4oi04Nx1JlKLQ359pibdlhJX4VPboZquySuxEP51ULi3g+TrntTi1E8qQ5un
pcTl8OAN3SGiYRDKm6xQWZh0aDmRm8Osp8OH29p1mSPtnHX+9/1hJs63xpu2
CXW+2Vwa4h0WmQEJWdiDkTm9FWw/U+pSDrNZ9H3m1aDHvlTP8NW94Z/52suR
0Cp3qBFldPjthP8R66wYaiCCeQzgBHRo0KJxgA2scb7qJ/DBxdPuaRdJSHAQ
cmLE7Zej8Brs/022wls7UlsYt7n9IdFC+YUavYVdj0RH/Uib4vYT2CF0rCCF
G1Fhxop9rvTPubZWFU55Yx16d7RwY8PIkfoKx7mXIkkPPomxpurwahmYACSf
DttWyiFSR9zAFp2TFqU4cDlYhinuIljptx4RBaOfT3XS4YcjQp+LhKH4HreF
4/X/AkTzgaeYZWLFMhWKtUf7H2SP0oHR8DK86OzZJhVSysWyOBFAy819BWQW
NzviXh4ZrNmdSaIHfy/kmwId8wmx1VTxjCKD9Oek27ttHz1x9UK5V0Sal9iF
BoaCQpDaKduorLox/iSbVX5lQ9gCSdLm6TZPAwFNxPmLeY26zOcdjBkrWuf+
uoUBhi1JE2i/Ny79v2aLQ/CAMUC9+7PkOl6noC8r4IwkyzwQ4QbhVrY4zD2b
FUB6mDi4mzZwkRcMu2DsxQpLwYr2XH8whOd7V1EAP6rDr+hGfmaCgfRpD3md
Lv7ppx15hOezFbixQMF8MyK9FN+1WccrE5Sx1YnXwS7y0GUbPjF8DDs1Ybq9
KLKquLIVHu5gggs8NkrRj8NNYHPzfcSmG0UuveknlKcj+3A7JY/ljT2cegYg
YIaOZzajPuxPNie1/fvK3usDLY7SC26dKreCQkhjofQSN4AEa8O/uCsyNLF1
4izrMX/Gdx0eDY76iy8Lqax7eD3ak60aC4xoctWrVnqbQAMxZaZqakie/0T+
ch8sljU6kLPFOpZJcEqbo0iQvgmnBj0mS5XP3Hy9kZWNqijPhEd2bisfFYP9
aXj2/KMIaMmVByv+NnPIl0Eh25vEVv1568g+wuYHk07w+ZIt/6Hcr8D6yBDW
vqY4owaiyDwxk5gXQIQEjuD/pbvGGKxIUTuFeTZvXvSnsBjKy6uV4R10f5l1
wAU0vN8rMo2MVWBT9qMna824/iAujcTtiP2lu4DMS0SRtRWnXPoE2AzgerqT
3n1wYY9k6Pn6JJQue+w4AiQJHSYija3axkmoWimir5RhzcMnz5S1FVN0LHUE
pqV+B5wdKynD+XMuBcRtmkLXdRNvIH3xbnxbjxbhInIrF5DPiyVznkPJj28j
UgE2aPL3gbW9kOtFFjjoy6KBZzKg9Dle5lqRRtB3OGHdckFFhFEegpfreHUD
UQu/fw2sVV59uHbhMUMDazU5rRObs4aexcCmxfhcWTqgMRm2bYeQlomnyM+T
SCyaQ52IiTE+RPzZMI6bE2SMhwhRauED6244cC+tlfHR2drP69ZQxaxmaCKy
XzTTuVJH3qTMbxMCNhsduattWuCetpToAC9H3EMr+TSH1MeP1iN0kQOAWyWk
H5Mbc7K71G+Ebv3eeQgqPBPz90V4Xe57iAiQGgQaF0JHTXG0Mr6AEnvGjK/M
XiM6dpMjK7kbNDI4jBhTNrJAruy+YiWXluAkNjQAQ5CnEl5/lgPoUsvUyb8M
3NSmeZ8xE68vqipN06KDVO87tAgqUV77PN1sY+GrMCISyiSNMLAs0PUnAjWg
DTm4Xj1iDOw2AcCK7kB46Tw1yMDLdl7L4NUN1TTiMLiG2WLPuNZdC/liRmdJ
0Iw8fku1JQZVb0Y7cioUm3L4tC9zhuGj6Qsj56iFJyB7J5FqckxqVv7/S49A
itgZmRN8rVM8bI+MmKal48MdqenUIfdM3FOpZWckazmiCOvNo/s8UEh5Ij82
4U9dPVxyQWbGwwsmUWGF8BfmG4gvYUOYrz6K7Z69psEc6sUjFRAk6KdAwzgf
xIuf4o4KysrkqsvkRkgl05WiF5mKatSeEhhZg5KJl4QpB1XUxYzFp+8TlI4F
mNq5FcpjURQ+uG9CPaONiv3e9z0o1pwJCfutG4mDw0XgYjDougq4do1MVIDd
K1NzAFfWrM2fsB+ERMQLN9Vj24WoChxpra24TE4D57lDyh48MkJGmhcq7J29
1LJBPEkN9eeMiwYSKp+lZReqXCQTVbxj9p4+p37HRaNLZ20dZcc9UAXua8Mk
nHo3ZGp1MtoaWALEkuXJ4afQHZe3XkTu3yESltApw5H9XyoUjKigkGFDFCkB
B9BUxDnwGoD8jZNPlXB0K8Q92NXXOcML0BhzjE3sRu0hqXZ/g/nVXDP7xdaN
cUMqjoJfe1XHvBAWRgU3VEaIJA4mOC6fK3XIO9OCvZIW1Zpod/qvqg9VnPYD
VH+88/4cHa/YB4dfqrTgafCUyYZCW6v0g6Fm792Jfd6Q8JW759hJf/xRIOQx
smqFdWX24YWPqI2t4ggtv+I3Z41/SpDcJkjT3IMEBrcoWnFDqMf3uhDK3YTo
fIUL23qkPiweBt20mDgF1ch2aTVZUnu9Tg2Se0817MniklHwtiXHwLjZdAOJ
QonzH3V6iEauRsKwtgrItK206zhlxdCrhYYhMvlNASg7dGK1/Cza8LK1PXAh
Gin8oQdqplt1DmhTDtwmjmYgc7WeEtFJfUDd6Cyyzks5CtfRwGrstXb5vu7K
MTd9Zs/k6WnFZKpWkweCOB6BgGRT9ISHNhHf/gZZ2+X4PLV1p9XlOZVpXO+/
s86p3FJooibBSuLoEecNmKc2350MLmM7EHbnkyIzEoZBFUSu6t2wvfwW9jYi
dNFNjuEWLZ8ycck/h26C0RmJ86i9LKxSs4oeabO97ZNWXa9fXm/YTVIbFmBi
UAEyw2gpqwogTRqUoygIC7UaA0vS2IBUTRs7dRk3VouuSDQOKmNsd4Og7reB
fEes0+QVnqFKhyfKhNGrjg0crU+IZz/ExPXW7TIw61qF3tc20YcZe6zi3D2A
2gMu131hYIiXkXtg3LoAzakTJ3FuB443Bx0EB3g0VuIwJj0GKEO9I5diduZA
GeA7U4up4jqfySLdoQhzmZkwCxMsOogvKSIGEOynqRADHZCeWvDeBMp+IVu8
2a3CDDrB0tE2YSjqpKcgAHE36JP4Rgj/fUMQUZEeOtZm5fDqOW7CeKRf9MDQ
MyKofsD4eO3mIkDaRFlAx45nCMiNYgACbleXC1WMdXcwmefxLUGhBQE5itCb
IEZSOTB8RXHBN8KH6pGUVb2Nsli1ueC9aXafDfDcfSSbf9AAmaPQWfJWSt5P
taCTe8Yh38FgWANN1+NqAt9DHW8XFKkoPRfN7cGiMi6QVK3B/ZkMe91MZH6s
HjbXzUKKjRSdUwS9WljlBcqFtsZvxcQjywrvgTqAfQSA4pwMBnKlJeclAx0S
wiR5anGdSpJHGtsLPkgIGRayAVY6QtH9SzOKua2o/84yODwLoRCN1RrfdLwF
Ub3hmWk6R3thj+w9zBgt5+auDwSh/hbT9OaaR5/JwXBwvXR7yUlMbxFlQT4c
4VwtjWD8782WlLHDQgUi01KJyTQ47OKepDCUfpyEpFvmwfsNnBXmxaSN0s1x
IbkylMHb74pVGmfLVW2TCaqYaHlBd9AAMQSuC5l/6hcRCXrRRN9MZ0SNqpiW
MPUPt4JxPRoEZf+70GsnZ4ff6URO2z9aW42EdL8hYYJNDz35WvrfiGvXDRSG
p/9g7F3GxZ+sLjzksDCJe5Ko5WJwhYfWyLwlYYkNm3inw6WqeSjl39BW1Ny1
TWOPgebt3m+8elWy9NL4/DaR8G6dO5OAnhcX/r+g+hMTb8sGlCGXWsUhU+Dl
oEOTAo0QlmTqKYycx2YqaUnnR0xwQdO8xet5CZcyYhh96TYwV9T2Ha6T4QVF
Ylu5DZ5LMRgDW4phZI7F2h1ErZIViEm+XpqUgswKMgD8jd2Ur/Fnn7QApUtx
rYLSLaZPxDsGKk/dZrvoJuHgrgKRBVNdyaNjzVp/+wtESFahga4sIuwjOBJ1
AIrb+/qfCxsnO+MKsK5U9DFQisfBoe4rTpuOnolk0Wdq17BBtvOUNVsboIaP
J/npqDNOGxmNJ52YCZa1ksqb2F6P5zm6Szfxo8dOYPPGbOhN4sRYw/bXKoOT
CN3uGqfCaO6TKkAm2k9fnjz6jmD6CaDWD8jdh+1nu3EQuyK0oFbZrObRpb25
/4N3KBKsLKHjl0IdZhfYCFqrKN0TVN4OTMg0rXtJNFjYiVuEQ/OubgapViJx
0aUBqnyXuKj+pukzLzZtoxxnQfMS1Tb+cE5Akg4Si6sJ7lIImlAxPSsdaOfq
uBBMbh+XykmNJnInBcITZf41DFA1L6NFuDv15g7K5aZajh4fXma3wXy4vubj
Kg+cXM24n3sjSlsRrphE+sgRceUy2oqzQ3hqQ4iVEf640xXRtRjacvwV+fLa
eWkbPiuCAFl4q3ditjcplBQXqnMRgHsGVzY8AHlXviySidywggFKadIUXa/e
jweYamB5U0s3Z/xSdVOnUsQYkYarm0ztdgaeNsbyQE1tSizSU3RLWPS3J/yn
RFsBj17jPhAL6V6mg31CCN2U4A2gLZkpXlK21x+KRYIWXIfuD5ijBCZSB4F3
HFb1VoFKQ0WbtoN85Jm8KhGOSphF1sScKyISrfHPcTx8gukBKQYQnoSnYqbE
suCh4gWj/+VZLiYrJQsbw+X/cE3gTM95xpwLc15fp+pN00sUtpbwTeuYHaea
zT8sMefvVo5GgCN7lsWHoxu01fxZ/Q9YEYReQefjO6oaCx5rI3sjTLT8vWIV
YQGNjIJ+QKUSPJLXDMaqHAmjNdHmc2tVFwlvu6Z3u71KpBO3tKPkmxUtFtE+
f0DaG6M73lCCaH5/wac+nLaGtrx8VINRgARw7hQYGokgRqWRjlbNIA2/TGgA
wQa0oRGnVELGp8Fg8PWfJBLzYIsqzgZiTFE2jXQD8zX8Jb7cPH/dHNxATOxf
Kgt4FN1rC5fkOz2UErofUcjtTmXW41yRH2aC38OoBrvGEExG967/l3aMbULn
hpLXg1FSEQH2TSPgel/IHU8Ghfrfsp1Yu26pa3Jw9pUWsibx9cBGMloHJPKY
dfdnXQ543NYXK0wf0AH4gpHdg7jpES+dOcGNj4CA/2NrPHhDF+H9fJ8ZFL7M
+9QyMyeKd/8pqWqHSk4B/on5w6TI6LnfPLjolaSBTH//o92QJUf6XjZ1gSjb
sDVk4kPfio3OO1sAsvJPuIb5PUsLWlQSl993DrW6SpQgAS3RkEMLfJRaQdWS
WJPY5+SaX3ELVFZH4uTQ7RvvZTKzkPbDMikfJnhCXdHGE45edg6tOmXSU9og
VkRcoBqr3/FvMWscEkEIay9wLmzvafOmQ2YcQu2ReT5lA1femJEQ7MJB5Ba9
/TG8o4MFT/bpeK9lhKE/pMjjqFco0RI58QH4ltgycs2AV+aBnrd7M73kmuHu
cP9x6Y63HsHmOS0IxNBNf3EPa4tt85Fr+y4xinuwnWm/90h5xWfh1QuyINLG
9RDrMcBEs371/abmW783YRCsX9t0DvH3bOWj6NIUsOSqHvo3RSZD93ceGGt6
WP+dpCHtwmEqbtcKhq00rAFXQCXGJQ2F5deDBBPJ5IXB3UGZZXTH6Bohl6NP
SRSON4HCEIHOm/ky2IHAByCwxpFzjyjlMSE/uFYCQporxZEdxDlKr9dY+LnM
OBzRWYh8GkUf8vHYxS65s2lWgu9UetEvRc7SLYl24M3tV7rcdgmrSBgad9VP
syob/wOlA6fCYULp3IRT2PoR0DvQVsvIciKSnynIl/pYiXgK+CV1XF4v0Pp5
dNt7QgPh/dJSuvgRYzHJx6xLwBbnyUF3afnrIK6sss7Gh2gLuFxbOG9Zmaft
k9e/49/Ux+1S3FgXmtBsFJhjHvmT4M7EdoEOadRXhkr/A//eR2earetNvVwr
l+UvwSk/9huI2omAjx8e2IpQNDbYMEuSKHGPCclrqfQ1/aKstFXI8J8Qk5LU
AlWHIDuvS/6MSaCbCm71mMdaiw3KVkP4rYitrGlmOIw2cRNmLqqsRJ8vv3Sp
47sLg79HtkVZKZW/JXiL3Lm0P4lFKkjImsSJEpGDo04v45pzbNnRp9A1S4Hj
2HexJSBVwyaEXi8xx1X7yaSaqsaeNs+gi2hrVfIhT30pzzz39C5OCsnCguXi
kBm3tVaWKriD7PZpBIMOnXCCJ9sEpyKYb25pQSdVHBkr/SKzlvL4YS8kDWI3
ir38bPhWZYri2CaJWM7yAVilsLriUsjCU29lLF6+0pu4z6Rzewk9PzI6+DRT
SdvL1TzvHQgjE4nKoVThALmNmvqCVArYgkpZxHjRJWbEKbYkVYy/FLjrZx1O
2LsoReEMYRFedhnTJkXxVuz2we4LI49ilohgyA68i8psLNAE6G/SRKKajjyH
+uMKoiPAZsT+X0YR3EYwYi7WzoLCcJJPaZ8ZofDv8zAy4dsfiMB+TXaFgGdm
9LLFYt1LAFLsot7ZoY/AiJiYrdxzY/BMOlXMyysO6SaXVTYcqiY0GEpAwibS
e8RWb+CpI5+r8RZ4Ln0amKoo2N6hlXOveFK9YOWIR2v07jYxpbX3ShVjNl6b
mOVRPREX0Uims58ktuuGbJYTWofRr7sf5MohxKSQEE0QDCiSjDPYkYLE6WoU
9EZ494NjrLHMzw4zSL4rdJal4TGvF5z82nMlt3PfUHOnPSBiO0UhBGeJUkob
oo5SQJ4qyVMVcpRhqPW34OKEqu48Uc1a0o4H2yMmQJ8dPVuv+N69Hh/vSSmT
/VMeE3JhdfvJwVTpBLL/m+zpZrA8jpsSD7WnBjYM9J2wd8yMbyl7pzXRZUwJ
QB49noU2qiOiCru0nS6G2w0AAMLEWv3Hhh0LRCGLrp+cE47feHHsPS1zygud
Cmbd3nJV9SWYSBBdBBWtbUEQ0ZtsGuSh//tvGqaen+1BZJtel17PCRGKOBSj
+1TwUUQk+FepTmhyGBIaFi9qZtgNMLfwC2/PsR3xPVrkoTeZNJNuJilLTOmI
/ydzUvrEvWDjocZeaoEnCZh9CrDHyaUtm52a2OQgFC6NIZOOJuV6YOdWbz6E
W6Izcim4Y6kNamHE0NJZtEY8xJAwimGQzyr+Et8UxXt92nlXB7KqjHuwBgzK
y18PWSwXmISywJSowxF6X4I8LD4PpuKQNPUspVFPJjS/Mi2ZEMWRuICo6+TW
vvebFV7py8dEsptYciZA5aBwgLz/KRKQDcV1BXo3HdwJUXN7ksoZ+u2WhcGA
iBL9T2gVoKeGzLfE/ayTVTurqXE41DJKvWGRaB61fO6fsM2diz4Ych05pLmZ
Hp126K4LaUJuIoMS/7Mil7cu1mhHKD4wtHfPz0LyIIQgP1aeYG90io5LwQYd
rt2AYiON1en7P+oHOdDzgPS7PMkD+Jfx4oWlHYLOZEAlEb3KmyB2yA6DhOpC
o7tyEe3UAE8r567OReKEBuyJMn2po4EzpA6IhNeH7rzc3NnHjK9Y4AHVIQGI
FGvIItuWk0IgEK6PqFs2ExBnFE2s3AbrWCdazkexALXw0K1paiIjM0TYALtq
ThGEheSs45eYfQeHaHsJByseNemai/G+Ewe6cla60QFxgEjoWZq0HSh8UKOL
5mrSElThjbPZ3++ZTWX/aPgGENoXztvTp8noIcg83CioUd/D6ws5nrgh2ofx
KmgdlFf77Y9Si566Uw4ix4jc3JHhwvhUb9RIrhDg3I3MU2IkbxGr/kLD4u0i
Y6sS/dyA7bNvnY4ZjDoBH+d5M9UGKG1DDbbhviKLAxSzzc+m05jTUVYNWYvg
nQVeneio/Z26Qo3L98B+7LoH5bim3kDtxgJCtRyRWB3BKIFbGHPvVthq8Vjr
DqoJmgHCBW4Q2I4CCMuK5LYuWxdwYeloNBFS1L2bzuTg/c42Vb5Hef1Gz84m
YKmqpohOZrgJojuCnUQtelF6PVgjVb3regchJkok75HJzH6UY5cSQ83zC94Z
eJyodqp8Mb8gUbfQiFTHrTTiqlIPXqio+rHLPK1Txyp5KbsC2W0VnI67pzwP
YnV8cHtw//oO5rspvkTkAUI+OGajB/FvPSxEKGC1B/BwuQhDkDaI4d6mKjmT
GRxnXT4+bKxk0Qb/3BFxQ1nv/+gZicWSZQyIc2h/tc/bUIYxhJJkRhmgvLTp
iewjqrQq3i6NYLUta0ZhFGtPfz/0KzA0mexXzhnGwijHIe1JIu07ApBMFuV0
WWVr84KN4YCzLHL5uHd9iaeDuXcWN4PhtxLj55E/D6YewUz3Io+rFkd8J9ja
ioCR5rSpWhFVL14mFFFkFT/eE79VauDjnGcRNjFalhAZrxn3VxAVXLesFJE+
hBxzLMhTiDD+q9BDmyz/SAtwHs5qbMRrfgtJ91zc0TeQ7eBRI530M8NuImDk
iehttdmPMBieQ36zJkCrrY1xngQVzIqHWbB5NjF6jpB8/xQWDuwVoykypfNm
HtdgDuB9+cfxNFuaMK9k01/DuBkuWTziAWUuQw0jSD8CKyjMoXoq9rcyniIy
d1Sn4zPk/M7tGyN/5ZEB517sEhQDSysj1t/x0mD7kXZDijS0m2+X57eR7iF5
1zkF7sDtmsF6miQ6dzJ13TVnn2jnE09W6WKzLOb6GFhKWGyAEYKu5nbDJ8xt
7JvUdpVikBQkjEXBdx4/XPyF1rPUKLMGCU7Ho7ZltZeb8QZFdNLin8g3B7o2
47ML5tKK71HuiLsDQm65Oqrk9xhiyHdayzo7vicQ9P5eJ/4JOpQIYWXF4bn6
rrID8+A8yPSY0Hm8AejCKpsJUrVJxasitfP50f+MzZzMTqiGaA5GaNMYFvtn
CPEeNRO+WkyUI6xl9kTb+nCrjEYF1YpLRuPMHxxxcANBnLSaOzpxM5SBtnOg
KUKRY/u/Sop8TzccWMJ9RWd7l8UYrtH7T+A53b4A9gNvblNrwm3EZB/9U9pN
XBw3Eb/RFQoLJVXWRCbY7lxQWQRjutJtQpmW98hu6GTYkz+Ulvk4nZHVuvmu
aFDDjMQC3yk0qgnDzHIrk6yLyfWxDMWRr6l27PwSeoM/g82FDNau/QcmbHzK
BFJvKcZLj7p6/rDag1VTv3o5RegcbDivvfoAfMQ4Ah0tbWLhFm3T5quIL5n+
kFNKHDrhUc1eYfrn9GkHWBJLd33Zi776g6sUYLGEU4pRyOyFrHmgD9l4H/qD
HVCFH8iXmzDo3OaIqmzdAPNzGjXfokEKhWYd8L0vocEqhrJ0y/5bTQ0DGKtU
6z3imhbVjaJ77DHMMa4Vh1PppWtY47Ezu6lDd9w5B06kJpptgctbgWroVydK
E5UwGr0/JEu6QRE6Fj6krc/i38ESr/nntdAWrTRxq3ZKgnftlp8qhogy3amZ
dUWtz7jVWwZS/jOuCnkqbQpAOoIHd2IlTVhc4MR7VkQWsvhgK+NCfHS1fHiU
teFgjSL7bNdUMmtFCl98ZRlIXL6HxIh8dpm/DkR2JwE+lWXasKr6jAA+KfH1
aohQfx8Lq+U2YpX29pc/phrthI5N3sSOHlaffFVjg6cqkAsKtkgLHSAhmBD5
gUcfc8CUuZlLgrce2BE5rhzBdL4E8+YG50BAE5KtpeHDHkuaIfhw4oLFwPTQ
KQEAWzE6Ck6LI+FjPRckvy1KrzHCmuXmQqm7ZIhosGUrECyCZPG8WYk81Umc
uXFH7Xqfy+RyR5X0e8XobaSEeS9NEQLdqSZrJ6JBRsgMxHborr8+sCoOGw8/
j3qTArsQrYva1Bs9gjpf3k2OedcmJVkBNEv8GLi6jFpNtg9B+JA5MfqlONbn
RzqU6c8f5PJuAaVDYBqL742kRnq6+ofBrej4ZAIA/lH6/a/0M/Y1AIV0j1N3
IVqTjErIhn8/jVH0NB7rgvIXvuMkSVxndRKQ5WC4gjELsdBXGi3LRZ8poPZd
DqEOvpln5+I+L+dX5PemiOYto7HaxdlUhIV3bUfoRgEvwY9rLygbH58Bw51U
JblKbJ65qYuV+46IRF/GnqsdOoRxrvoqT2SSBbhuuqp/ohd8B9tOhegD2R3v
ebCTgHIZ90qP3ND/lutd06s6OScbXVCpzisMmTx4hq8xAhMtb4ZcFLgqWDk8
YLu+/7KJTMI1nr/ND4MziLXOrOfRH/9P2FjxQACNCtQeUjdCqiK0Licb5Lg0
3pHVDc1nXorojOt8uJKbWZ01GvfrrSjfxUt/n/hiuvgYBWtGYT05ujpfjl25
2D1PSP3+pXqFpQqsaI/jnyvX+q38o+dSgNNUXkgNrkc8HONrmwmunPwNEvHk
k0X8JDzy32ICYexuNxdmbj/w0TynC7E9TGtGyBWyx+DMsirQaKgnQgLOuBzh
v7QhG+oxOP+rdtYD5Ucy7P11ImzZdeuftXtoai6OvTzHaoepTnKK9ULVpzGV
66/dSaa0Jcdhl7yUIFpQa9AeXdlVP/OkB17rIGgcqWxl1QN+2gtFIzXPGuBH
sqeMQgWu/cKokE3peP/5z4Ew23uCKwVcPyG4QtEUheGUowA/qmN5L1JUQKen
U4W/AdYlu10pVyfFrb52BuvkxkwQd525gCwfYyBFHqgR0f38POiT7yDtR0Ta
fuhWwvmQKY1SixCW73FvvRrWtlS4J+ne8c90L/KJt6RDrxmhFYM+12dQAUb1
y+dPP9Q8J8rt69n+c7KJa3pQkH/rcvYrCCDs7xDPUMq9k8oJHX2GO0lONYfN
pAdA+MP0fvmQgYG6DWIVt7BuEHqCfEtsmsNAVVIil0fqhZk7Ph5ZIyx4Inif
uPbbjJbFJrzCy8acGI1iT+25tAdVlOVHRRgzQYXiHCF/lMh9w4+4eX8qzZDu
W5QlnNYML0FeY2uoNFrDSpK5wYB8wC/yVDdh5v0wnc4z0bDQaCc5kxSlMRVC
teoBcUMDt3p6nmPYsp0AxVwzDKt8cHrSbjitTduPRaOXBSstmlPHgkeMtrGu
f25LFl5JNhG46Ngby0VEG9qvWxohCb3khifCRKM+Eaco32nK30b0kTLopvk7
ApgLZEmGdjXNSxdJ/+r/0O9sBr0pybqLF9WemjzWD0cQHfVQkiO26hAwowMU
dmiNtr0XtqfxPz1VH57+JG0tfO4f1ONV8e9RhRAJy5hY3cIP3EiueZaikGEH
yAxLVYc16jV40w3VUxeR/FzkE6bFbEA47BuaV6NrD4+eNLAYDXf6FSTx+2oE
awp3+VJdu1ZDFgOamkEgyvhd3JlXuO3wQ1YdnYucYc+rF717OST/p4sxF7b1
8FXtzhBGfu0VLUF+smR9pDoQv4z/psipmI7+YyhyN222Hf9M7rMHTLHPi7jd
Di2hUA3YwMtURG9d0LRPp43Glz/P4OJd8HPRqDIIgsQkHDQdlrdDhj+g9Es1
KjrUxCsXocajYnnDrNpcEk8q0ecm7DF8K0eHC1uAZN1RMwIh78qb92zqfi7q
YgzfJ+gzY4weMUHeGEmr2uQkGE3pSiYI6TdFS4nM9UsQnT7BWOn7ER5UxDeH
F1XwBeFN1Vk3cpxHTmkV0zAcjT/vo9jtPihytG4hZgoQCYk+E9tdv/tWwuL2
jJLOOcPh2j9VDFCsrAQcFRHaP5kQBs/W93zUI0wdr+xz+hwtOGQl64zaSxy3
TN3evMJQoBqSDz5xm+5fGZTOcrd+YQm//c+V92Wa+ND0WbHfjjrOqIsPg+r4
KgzGlANMUgKbqF/LBZB2bk54Aik4mnhks+CT7VqE7nHvHNHIyEH8w2DkZpz6
xUf0d3nh1MWvmO5ckNYkYWu1ywsVxjeRPfUtkNbvd9LrEgmFmPNaGWgtjhFU
0TR6B9CgBSpBdnMuAsgq4M6GmNdURUsum8ddAPx7GDOjCrrWYlpr+6znFj7+
MKbODGKOgi4dLsoWy9yCm/PDprk61Ly8w4+Hn/Q5rUEmSvtj462ZSFZTF9ud
ra0uT6GO/LgwF+ZbeKehtVpiopW0zF3j4gERq+KnkBKCdYy2HU7V8GQf+u4T
7C+NTe4ey69U6UyZRnozAt71FBUpD4WGLQhVn9RBSmOpLUCJ+OBx0/agZ+uX
4osi9sFPZ8+NFkXNkBmyYXm/QgXrbcujF6SzHym2QGPT/VSCaLm16yLQPERd
rIH0UbvsFHVV0dBg1gLuk6M+Vxc2Ff7aT3NM5ajV6gKZKVkTgZhw0EJ3LtkS
zewrRpdVyB8mw56bJPEtj52ONU6P1qTyDeSuXcLkg2gcJNnu2lB39FThU+Sx
jO76lLaVI9SfqzC1Cr/A7BOTXGMOhdsUP2ZJDXFuHazJb/fe6s86u/GLr957
Fwb5AJJkakHFBuxufHq14VwCCp7R181HMgAw6KQMeAEY5CBj3fwg/1jiOruR
Q6Mm6lr4XtbOC3MXn7+9bLiSs+TEEdrExomgYGfIPt0UxaObBCu6LQ58TFFO
EAgN3dJtakvTbeUF8vXKgmbPG+//EQXRbHgnL0pWXcIMO2/YrMZDxZMG8+LB
zE3M5d8kfW+cA8njH6yRdw7CuiScJTC5pK2kvzeRWT3GG3ZFpu5fvI8rNQt4
cKDueD5lhBYcx5S3ROBGyqPA0CDMYEvuVPRP6p9DBqN6n/HEvuhlJKAdXJRS
4nGSr7OxFmtdsuWym9QEHteiNJzjDyOdWyrNEOKQEY9FOJybwt8QaCRiap2k
NLYqmyT6ejSD77EWgqMgiwZ/8rczoP3R2D7ql7gRsTnZxePuJ7jY8aTBOM+S
Fx/aHqQaZhCGleyWtvcKfeG3ko3hLw6Nugm7+MnEotnCw1Axg1SsgswFA8aC
eTl+8VvuntsDD1oaxiJZgQr7SGjenu9xgPkn/2aYTv/GZmUFAg8ch66koepZ
PwuzxQ6mXn3NUR2OvaKZemVGWkoSw+nEAB6Bc9G+VgN6Gi5kIpcsJwFWTiNN
5ZIiEHonQJAQTyYyQEOPK00eJXlMTD9hnEZuOk+RffrcNbxotTCVnambrTA3
9l+aal+sdP1qdLrYhPEaJruT/fQwpHU/fCxRXbCiTb+X3+VunTyvbW3N31Mj
a57rsDZEFfhPJJxeb36qaKe+g8YByVKz5GVhNJjwdf7hgu5TK0RPLAeMkzIW
eg4aNEmJz+BDFi1AH2rJkIUUcT9a8+4wd18OHQkclht7F7/r2zR5Xp7Zx7/o
0gBfEy8BXLKDpg13SJ77EIpCgjWh36wwXIH06rKwcEvcJAuzO1yvNyZTN5ac
d8rY5wbDnYTIN8B2aAvRRS79ggl9h3NLDj9QCX83HYsjW4OM70Zbs39/d/zz
D3y5AiiXk+eKMBVCnUxybEGhoOVT5W9IiZamOH4+4eqj0+OIMSmSXUjBTyrn
9oc9BqkkJS3fJ8ojn+GAL3sGFYWjj4A3zvAm80HTtKeGA8d+1uMbQt7s6f5l
19yklIhtlo9W6BJIh2/9RpKtD6TjFgyGeepSeVQA4XCVVCesh+ldfhzF+bcs
XFkuer0Qf/XIZQgoA3ejyiXpFFqqGEC+6U8/sTLWLOzM3BKmW1O2Gl2hRRe1
HgkQkyDTGOReGTGN+naHYa5kONWz1SmprDdv8rGVpODd9ihcHByvrm01Fa2p
ALuAOFGAslsBSz5bbgtmN/VFB2WybJtNHw50Gt2vx//noH4GVzAaDul/v3GT
I7rE3NgqbcGfJpgKGF7Z0tueYzFbsUmgQb9zLEFdXiahs6M9jjy/hGkPzUVL
7mmPoKr4RrWhrEs7TJziaq0PsSnAMAJDEH+mz6FzSJAEZcHq4jeOTvMDhCoY
gKyOZa7OYcTYfR+pBzkj99D74GsQBMTsenbATTW0DNHpVtiq9yeO1i2et+VO
L6WTsqTqSVJaSMAzAexzklKv1lHr39zyXD8A1hqP6ZbSawHO742w+54md/dD
4TO4TxcOGJM3vAp+qT71lYEF7A0+jwe143zjVmsknRHpKbD18VgW+QO9ew+Y
B9+HJuD2zb5MRpWgPgBlf4DbV3P01Y1d0857R6CRWDO3FK2oPe3+pKG170F4
arot+dUyb+5gtzfIQUBWvY2SLTT43xrweL+dRx4O31lN0kiob5zFXfqBotTl
A4UA2nqh6OUuEvcf7+63MOI7d7Pim8OhbPck0AR+t/qzsSrLK3pj/s1B4xKc
ar++HXGo3R40bQVg0/p09dlzFkt/W0bwosewkey9fk0Yj9d+YbrhHbGFHSEc
WBPC9GtIbTYxlaCtRYltm6wjcJ1BYRaAJzuq4cJMlpW8DHRAVJUQ8pZkbLvL
gbsSxjBu52PsLkhWLS19fXCXscz/NHuoOKylTdVFU+w69YX2as7YVvMWSk0r
HWQlJOpK1uutax4fw3L8yKzxTsms5dL8s+88Sj7OTheNqVHrW52ldSEiChcY
tY1Fhzg84Z4HHhRIKHMnQdtp72A9Lu2Og4gFTcL1+u+7Duin7qjeGCH1Wkmy
DFvUs4z9Lr+XChcPq5Z8V6ECZ5dVs9L+PlDno1Ofsz7MwjlXFntmGEaUmMjk
VrE5uS90wz9JhyNeo5psM5ev4aARsumQXf3mJBEjmSEe0ghQ7Q3HSAaXGdgY
Cg/cyf6dSXNeQHQHc9qGbk7NvBOkLlEwsG6oszqnkeZq8BDE/vtyVKMB7iVf
iHE1vUDNbyrA4jmAzc68dFC7spQmPuVOmj0U9j0ZvKcoONlGgimLE6qq11y2
TpFx0LUcnr5R/KcvmNLEDGzLruLXc71MCtq2BEH7nHsJb6lV+a9RTeDLj7NY
yl+EC25dXUtkvG0wjh0YzdHL2H7KTtKrXYCxjkJV+N905JjtPY0R04OVJxGt
tERDkiHmBaxebUFTjyATcjHprbl0R1pqbQkiwoiFJZF96CJy171Noju1N4AG
1CR/lSyiR/2ui0j9tE/IXZZPWabbTDwmz4iGN/AineMkGNu5rqbNf1Zex3b8
Az7LNxVgp9Q8IJVkVmTDDivg6fzJQk8gmD/AB7Y/D7QKnN3A8kJaADgOgB15
U6tPYk6ibLiqUFiTcMNm5TKoTDiXAp96OurWmMUmykrnRs3zk9wYUTNarHzj
n0FLqihWVxXEKzNH7r4PKBe32QFLRB5S1+cLzTk0Sl8DMZ8R4HMs3b9pbRTR
F6tA5Bi6IirrGoOjchoGq78tv2z8vRSHovFzvGRaKIkNvoc6WMQvTtQgyJF4
rRh8qr1G3ZF5rV+pN+zX7LW692P92LXzF1glJcxyZktiN60jqtNNecwWfE0e
aPxpeEGL4fbw7PX+SOPnoREvt0TlrH+Cc8XV/jkppgMhp99bjlVoHpF7SvHF
V9wJcTWWJ1092G9B5eO/uH5OqUWs+opuN5SQ2MhCsyOYbpxhCfb6Ir3TWAYq
Rpy90gF5g3tpkgOxOqKDQXS0ZDbb5ihObNgMbQIP4k6HQshTeeH9MMlfQIzn
j3L2HnxUyG4mX+3OCdDsCUD7nuTbC/61JEAI+iaBjW45IuMkDdvuyt7It5/o
3sSKVsrLyKo+HRmb/pFe1QQAn4o55rSYJr2Mu55Mj10A+1zF+hSUJIHgzpQe
iB1SWirVMIepnf5520+72P2Ri9LrgcipuEoOVNY95KoX2GayANjpGfSvyYD3
Lt5UqTLGfolZAxrbQmUxX1kcVxg/zZO88ubpBclBiFgem4+1KGL0wWehLSpj
j0Xg7ogIs2Hr0EXsB46m/jAWozkVKVE2w4+uNfMygBP7FUxnnmacf/iZG4Hj
2W4/NPEHXgSLOe0OEaOipf460lX70E5HqYQcQE+y+ydXvWALbQVCJHQDKvy/
lh3Gzg2cRdX/uJYBMhjsDV8Ub0ELscbWTD7hXwEyspDjP7dZ84KMct6+RuL6
Q4LhyMsiQw8F+NPBdfIblQhPCfe0/msftLb6dyLnSL0/Hrq8qVYdERcbUTG4
gd/RPbTfMdBIEtnMmGO4I+8vacx/X00N7JzrK+pE9P/hLe2OX92A9ppxdQ/Z
VPf29+byF80pul+v5ETeswW3cjJK0LycZuEDSw7jJFB3pFzSC28zpNcZoKCo
6oMLkuA4Gn5RYhnOaQiWeoyW9x13M9Ki+jJM6aTfNFoLTaENnNGkKiCTkjzt
a5+5frscnNYrjaEXwiOExtxlU3oGYhbeUkas2buM2Ppp13IzsZYOkxYX4/BO
hYPP43pfW5Y5ttyPOcCIg2D+95EMld6YUwZLqVsSRLwNrCcXSOWuNd+JQRoW
V3UHzsLVZthAr77FBZbynaD+vi22yrb5N6iWOISzIjmEVNCfwJvWjdrlONJ3
MGpRRx91btD6hlTiEjQXFt0sCP/vK1uy89mKPgLWQu9wSDJPZscYa+NqxUc6
XQvVElf2q5cSK1xIXe5eJYlCI2N2aWOHcFVf97XsXeaaWMKJVwwpjnVDuIyc
W3gcrpWKmQ4Fxo8j95gOgh8npv7MdGQ3yqBb0Rol4R8U+EXDhwbjUOmZXWo2
ymvuRkWA1/zDGBcKet92zulakfq+ZDNCgIkUUWpGJh/W74utVq93uBizC/BH
bQEqKxs8O4jX5lZ/jawYJhZNEsmjLew8OKOlq+aUlzEaDYqKKkAHKGNHetfn
AsAuh2HQMDga3xIZI7Qt9RcBHJz4ZNekDPmJTauTr/XxQAcpC5LYlvOovGgh
aEHPK5B2En12ND4KZvGH0cP5tFZ1mi7jjxQMV3vXAZz20E6Krbqjwf8q0l4Q
/gdZ0TEhI4uY6ioJRfmxpkFtZXzTD1GUKqNFWyQM0/uQMgEjVOnSiq4Dg1W+
8zExtDSanok/PmGJZ3oOfTW/7F2l555VQuU9Z5gyGbO2HsI6avyvB7YdJNjT
oMpQg0EKlU+wYIrqnowi0N+RIAdHAytjMHMkI77TaJU2Y6HtpIvepp+tSn4P
VDS/jkAyiYuR+mOQG7agNKe5DMlB95o5HZVu2xBwiNWqmFGQvHIAlQi7JmvC
NyyoBfL58yl/4H5o8PhzmRpV2gWWqSmOHevmY2uTWaMQcWoTRFtCaSlViH6V
mSm5ro3gVURi+SpaZc7NpXE46Oq747UApqoWHi7ILPreeidi05NaxjlvAMtP
YBk9EooNYFdXW3EPyNmhecMIyJcUlyvR69CMjrOgjUqPX4XjvjBIAsuFVxyv
EcVvSgFt1TcQSe7cc76gEzLNSP+eVzljrcxK468hGp1TAgokEtCDvj6Vg0p4
TBdCi26jnPMtSghUcmp3K+DvvDW3Qw1TUrx0+sydN9nEd3B1HDhAqMvlkQLc
xYLZ9CbN8hwJx7UzcRfnZVJkoPv5AU1Gun8ZIsKmvJiErnx/Fo9x1HAXamo5
seHheHeSURwmByfm2z3LhQ117FhRGCAVvEDMXMpcf2cc9MR0v6+BzPuLjcnO
Xa1YKn3A8wpvQH2fQylps7BwnjRj66h6Kg7V8U8X/aYRvivx+mCjyYBRS2el
o9jAK7sqh9db0Lz+rUf3zMNRd565U+CPFr0BApMh0HM+qLNZDzpMQJt+pkM4
/LXr6NK0G6XD6FPXEWcreAfsB2YQtfnXZCp2ZB5FM2PBSpJa7tDGwm5kEq4E
wO8EjBP6bnorxl94k92vgdxaM8lBkQScPgUfCxINsTJnhRT8GUVSjPyV06qu
Ug5NksKxStHraPBXQSmxkM7bPi2eSwqnLL0VitEJDWsqBMjSbW/m85KUkZJl
oMvklGJmFLtI+sjGwxzAhGGleaNLU6jad0lXWFWJajhagIIiR8pmynTxTERv
1EeSwWMKXZyK48YafUOvF0YT8HznDKn+onvQ8HxqDJpptXSYBvhzWlyRzsEH
HJ3i8V439HIn56oU0sLGYwWNCgvDjDR2FvBazMg3va5tjlHfHukCT044XtW7
dzkX++G91nFgpYsnxXjHRmA8B8VY4YaoAeA50XZwuThFpniJVhgNISQvu2KQ
JkaCiiy+a/T/FTCu/y2Vde23QKClT+4d9Y2IjjqMaEnia4+/cGZv2o8RkLs6
O0w6NFkYrn8GCUbCF71/SlLmpOBhj5ThAYAXqvOGA4GQGtS/yvvGf2PMAlM6
1UeJJBzDka8WsNNb2khwBEPf4EkhnopumLVPor1jg5LPZqQsZDuslZqRvMb/
56MWJwLSe+5zo8uCtUBz1aM4XyurgQUYNMqH6kuJ+/G3GzyPih58PtmV25ZZ
z096U1vqttF6GlghB3xIuRPkVlbF9IseriH9V20SnT7FqWvReYi8Zu4QRudy
33VbThITlkFkXcZqhBeHJcaFrNOP49TkUKTt5ywu7iY+3sKjMi8AkMZmDxoR
bju+foCZKhkVp13xXR7Pg77m7zIEsByn5PEPOtwpH3gDWSI0Br6Ps+8gVnUG
Z38ds4TcrSzQ2ofFzVcG5M5nCpqA734m138EpAHseNPELIPhxZMtXl9Rqic6
IRnXOaiePw/yB8kjgZlXowqWv/mYaC8k0NXPtEGPlwjST89+g0wMEQl6+k/o
XgCqpaGzI5l+Yk7+8bqhWcdIkCGIX4YhxaGXXITS8luZxj/oOjtieV2h6ZGj
2MjUEExVL94Hf5HkYnUK0ncHgpuFkYQi1q/0redACVo9pMmzOhKXBxhfC/1G
QqxTuJVUIRm/6prtLbLbN8AIEV3/vsQH59ZpszVbzDBwrQI766BRGU7N2QSl
uMCfRGfqYQfeKqtqY1gisjt1mcX/saeIyZ5f1J4hTaZjKkyhkJD92kAG0m0T
ZaKl9g0a6pkzKOL2J+oGdaq6voGU1bXNiyPZDDP+LnSH1D7C5aaG+abMVRTI
zzsBChvQzOQDn9tPpe9kY9c8QSe+nrpSx6+vk0kP/8EuY632jYiACks+4hzn
pVUZnP8/0L4SsvjGGg31PAOfBUkTNAiNYB6kKzaNh0ooXq5valxCwuvGG9NN
FxBN/TtZgKCtU4m3QR1qG3m5X4Oypyw/h0wfIbyW0CZoQCz0dB+O8rRbWzBg
lAmd2vjPaVrZ9EhahKm15bIqldATJ1AMWDCBr2iUYhovTBLJRsYDOVWZc56Y
5tMMhU0h3mSt8+6xGmRb8ixlMWyATRl18ErVVzLChC9iNoxMaoHUdM+iN8HL
0EYCngK0UBO2waLq293DLWh9DM7d8q0w9ZhJDXkxKLFK9+HaDFV8JHpWCkmH
fS2VE2BLvV2bZ4vGEqptbc4X68kc5Hl4poQC2WsXNwXTJh79XpeBtHTzmHmQ
QABV5/BHr8pGFQkyhE/J7UGWwpWTVdWi+6Q/KKTLseEbaqQStQbj2qind1le
5+rSsjH8rpIPo2peK2PI3wFYVDbLMidvAdt8qEjveuBYaMeTavmnKE3OgbTY
JEnlsZj+Nw5/mz8/pYmB9ymevrJSnmnimr+n71fZWqh938aWiqYp+1eiKuve
HMz51XMiqM51inZ2wydX1Myv46A+yqc5HqkTZIfjrDxI0N+TCbvPyGVNp/vb
xZJF9gr88I+iT62Rx4mWXJnOfCTNvuLOcEgwcjYxV75Z0vSYDpWYCLrO0QHr
122nEZfQoCGPJWzc2RvNurB3xduoqPslo37guLXOSKCN86QY5lExhB+xuou2
6bswWx2LiJ9COPAkGY406XrCVChQCL0yHgbXasrG7nczx1daX+pnVZ2nIjpJ
L6PeJgVZ9rk/Owo+7zlrwu4WRuBtecrJkw8iwj+35YregJyeOxStAdXtjlPL
V1sK7yU9mL6Y0d220J8QOoOgE/WU08eS5zXHxllD/QWfS/2RaIeM2QVmmWjH
65Kyc+ca/iICEg50rqNlEc1tg8Mgx9ZamA+Dm8HCWALEyCDhd1rOSpAkTPs1
sQ++ZIk2NjF63zk12+WjOY90k6NxgShhn75BTUiuC2s7UoLAusI1YUupcVVH
VXmyjPqUEK9I16d4rsA/mp0TbigO2ZA8X9JcpxZDRPs1oBliCxKoFCng7qan
SvKXVS9XE6eWXWkoyiFDwB8y1X13XVtfCwnTu1sUlBOQmsTSE0HuYofm9WG7
KnhOXylthknHbLpvtlBmJ1ck3aRDmj/otYiyNYHWVb9VOBbpz6c4F0wtJqHv
MRWW2KJAeEICHH1mq9+ZTOXrBIBexKLpuFLHTC1P8ZoPrYQb3l9HzOZ3aDQN
U53Zb3KwktbG4FXZ2GX4LBP/TwoiIua8VglsVfIePowdSAuV3nJYjnhvwtD1
Z6aeE/UB/OjjliJnei06ujT6WzNcCOezR0VLmAnWjcIMTtRBsv4wEKh+PcEF
RybAYDAClWOIsT4zo/1hwk8uBCwVH2jrh+aj6YPAFtB38ap5ieyxdlO8heLZ
QVAbYSu+Mb1KUybAkWXTcbKb0tF1a4mv90rD2sntf/xKxfJBZBmoZa1by1f+
EvWBl457RP701ZfDsKz/hokgZGPvNYrr6gVBUUJzkmDwh46Fm7sMcpohI9rq
5zn0PQ2X4HhI6GvMMKQJO14eeW6m/wi2zOvM1s4cL8mLGF5cbzZ5yLiacPpk
yXdD6B7qG/NES7caRzGpGNtf8R9BBN7qGl6hH4/jg//hrPrsaE+06pe8y/3X
6yaz8sMena0khK8eyO0GFle0ShNNhEhjSVwIckF3ScKk3k6GmTUjYWrt7uRj
8ymhvkGEhzcYlngZFuQuslSHY6vdjEOqHT0RlYWX4JBIMkNeVjiqyLbYhAM9
rpHRLGmmcW372vmjfYVCCV8+ccIX0kX2D5ctKFNuZYg7AzaLgkmRwaz7BIlC
qfupj6wzxgYyiVQBdic7GD1inwipCUK68vP7j5UrPuvOy9uxpIQYCivtapVi
rnhkrFJ0JLAhkeXA15Rr0BTQL6YHihDszFq0tLAoBEhoNsn+Nx/hY+eRA2UJ
gQZyoc9xr2+GrrzRS4i+EGBfKu+qHz62rtA2J20XZ18UIjcFLHq7vJv2RboZ
FpTeqJ7CSpxYa0ZS/X09iLBGkhkIawHTjIpKmMI6b97JUAFHPppqncp0ovQq
c55PpMgs2SkjhbDuDB9fhMwkS/ld+bqglWiAo3L8bTlVmtatJiRZntjDP0+H
K2iP42XUSWpIRwbv9f3ioXD0bnqMfYgHgGGVxuP661TpiAX3jeq6dSgI+Hyt
ZNqm6l1kRtU84pRPjd3QfS3twy+yT9mRfIoexJtmAEFtifpfzPFszx+mSETM
wRlugpPJO1SBl72JkPgeBVM7Z6LatgY2Ov5huLgsNudTVln/IaViUBNseqTH
s8jLSo/3AOIKrZ1nXaatg7i6oU/QHNzcu/QMoMS815wuIQnst4h8OmyBjXCR
t/PahdEMwnK4BuJQ2nqVMBC0FfeC0Ci5NnYnbULBKPRvPbqPO5s8PZoruEcu
CXTvyIkxceyq8MUrVGhr9k1zyVZvKdqlZxyg7TuOrWsZbQ9yW/wmkKcsf7OE
0bYWc88gnyBxsQPBzva5KlW8muPV6c1KvK43/m5JEnS2jOrt4gD60IRN3zb1
ugoDHR3qBvRgLWXqzz0+KkNGiT5yckyWbYce71vZCBcCGTYGavU/iw6YNKWt
U8IJyG2S8w6ayFAkTO7rQKkVDDFy8ywU4t3c6nPk/1qzVafMkQ7sKziFJjuI
KrMOA3ycfHTCmGHEyVv9eGg/X6PBmOGVlgt8Gjnog795Ngw0KKnhAwH66gfc
lPXkgHU2RDQxdtSrng7sdWVPSUp3xs7yPU29Nv3KIRnuh8/oxf9dsJXlmAvI
3WzjEE1T5y+R35EZlvSK43SfmM0K7KRBqGRdWe8f5s0TyYjBRN1gN8oJKxkj
0VyvBVrQ9WJCJzP64hU7aLPqlVnHb+Itk3sozKv3fmXUpVwcsaQ6G9L9EpbV
IC2iYrdezGWNBTVYr4XGaAFltHaGGhuoeiuReW+WV03M0DAZY5uWi3hg0vXL
jlQQpLbIUq0wsXBeBYVodCvO5/fwEuSK50AQKVvA4qVPIg5ciZwH0MP9n1Kt
OQ87FieKN4IGlMuMl1YrlklUaZl1bwHBzU9vh/9EGK8aSoUN4jLjcM5FkKsb
QrkpLO2EbygkGlvdoTf0Ew8hmchN8/6y2+2n9ihVTZvESGAzUp8yBjmJDY95
OnJyqSpzjkkFICx6F6dpP+TPxfqCC8kJOVUChOzQ7quNT5gZjATlx8iusJ0B
xgf0S1nny+uqq3FbXgNBRMlnb1CasNb/+x3aolbbVXOmOg565Ma5RGXtz2nZ
fl8ajyA7fuevDNFZsVP1Ohb78bRVxO2c915RIdrieFH9F0+4HQkyP/p06be6
hSgIQbSp+iJJICeFzhJxbJayucdud6tYqNt1mMuBm9pdGaG/BMHtHsdFfB4P
hHnEE9fxTXyOL6ES/UnMyze2BJNSltiig9cNQ/aqHQve07ahznEHik5qmN4S
jY0RVRAtKPiCJWV9dhGLm4asdEJVnWe+B6tE7eQbf9zy6uGk9BN0kC85uHTR
gcxcxt8hvzEbF1gJzPBub2IDVqjeoBLnI6VskwM3riM9GgSPqEAO/J0xSw1Y
9YUmAewSC1GKaz4DSXdYm84KA9J25uyHzNFf5AeZOyACZP3lKEcHkoMkq//A
T2wfi2o9qPgoT2ypaeWy8QJlxmVcpgvIxaNAbOKVHTViAOF95ZYLz40svrEI
pxKmXzd8/zJUrVJowLLn7+i4tK3sk2kpMxanoiN2RWghZm02pdn4DvhFh4N2
YpBTq/tfAdWe/7NtSGtI6rcdyZFf6sOGNSXhVJxdTQJfCxxFthR7nyflNh4d
365HO5YOq2dmh8ILXbxiUzNvsXWHpeHQtoUonGGcZLUQtHKQrERidXI3c8vo
xCZonmz+oGRHsxHqvMunfO283YuSa9taORBtqnyraBpaj7jKI6CWY75Y7Ahe
dwjfOh7briCVe7YJvEE0U/LzUq4qicwA5lmzZW+2g5xYh8bQ6Hb3DqDodVV/
LTsGqISTK0QZziPvFicOodjXElOuBnhpQoIGJu9WSVEG7MmfAdW0mglk7cJ9
RuKFsBPvuA54RhSVEMip646FPwn35DCE6QzB9D2vJOOzcY0bkCouGbBSXHPy
K4ovjsObjpoE50xMcSOvi8pitJ1MooI7pRuZfAOhFybeHjoFmxFaNTj3LJmq
0vXzEr93La2Gh9MwWRYMUyyD3NFjXAzQ68xLHc1I5Qs6/+SOz+VXI4tOI2Of
iZ093bZHYuCyzfVM73ffHM4LP0PJngKV3uQsxU9oNIb4KJRAu++EmgF+DYP+
7PXQAZb1EHwLlkg6z2HXSRdW392ndTI2iwgiXs7WE4pEkb59Jvrqk7TJvzxd
R287ERTPJOrE1ruFvHq8WmYx7M/iDltGEz4yndpOq+ZYu7SNwyJIaqnoS9tu
DYaEd40dQjnZfHUj+TurlO36UhUNrUeFlUn9DbaBErIS4oDakZUDsqd4EKkF
5pLIuRd86D8cKTf4JFVtLzJES0Is0CLQhr43PpFz6KtK3nK/41xPARrzEbly
pP8DYbqDmSwYG8fTKJw5AcOqEFOsCr1U5JmCKJnQ0T1kvGv2Vm2axmrjJCvv
tffBUiFqIuHqb9XtPlU2IPTYmYkX0+zkJGYDcB5aEZNZIRjeKcxQd6FD3uAz
oV9/DIkh43wr7TLJpMGo4vX73giZOZtzRK8/DLYnSsIlbS/FgaPkVliLqP9z
m3WjhN2LOiKM8hoosZkRaWKjcVVD6y4uK/7Y2pZ2doK8g4W62PNyAVJdL7AG
YV4wbEqGr77ab4CfevWvW2X7bgq5eu3wSZ0a0akUzUGrxhVd6JVEJp0Prtny
g82+JEk/F+N1mPLm6Tzkxj8H/sSmjnOv9uaSyl6Py2GHLkAZ6ud3ifFyYD9q
7fpNIy7MgwwzlXsZStfh+mWnqwQzsK+AfMqv/CTJr8faz4AIXV4mRFo+XIMt
lvhkmkoTyg65jT41lsZb0HcBgj80Tl1E7nlSmeo/LwZDCDZNzvLGuhCCJzII
+MeqLNXGV/Vq1XEITcAZd6AV4wN5wsDnmb/i/120R+2LLslopbRgau/aYp8L
+SeR0ycVKraPLx7SDNamRGRPAvYjrR5MRIlTRFzXPqsGQqyZTzRZCVgMmFgJ
hauVsoNVeg6C+/oizXU61rCkBLPcAGe/5GBkjSp3dRtshPYayUbDhmU83TS4
ztm3U2KkryMpZGjFRgxQ6gBhT47wdmgxtuFv1vPY94AtdzjxbaM6T2SRn4sw
8A/EJ5Omv8Cb/+zpoe0d8TvSkSnKSdWDwZm3ND1Yd+pjtS8u323A9MWkKqOH
yUUo9ZuuqV31xGtexBximPLFuRVD7fJBx88ZovhvSZL3DpU+au9QVvbLjRoN
WEKMz5zBYT26N2hi+dMgWmVVe+pH5vA67cKX7HHkFB5cD0LuFmEQ3T7EXa9e
0ShYm+Gfh4uuGin0vMTnC/RddxPS9kYPbkht3w4yW8wIbM/Zia1P01f+9HR3
+tO0YCpCTRVnijFirvlhWYPEUoF+t07gsy3jdji25+93hKnazkceO4Ytvj4T
kGJHHt+QanA6Nkih7LVo4qdbaTDtKOrFhwc1YqCbUh6PENYwbEkULVH4hZ8d
fpoPznNR8EU58IYo/2ynuNocwXlDVr4s6ef1UTVK5yiUu5s/tlj2VXZjqGUe
OxVS51VbUf3dSkSRqwpjOYexXp0xsUzG9o4wzx0ttc2F35eOJA+2ErOnkqP5
se6HV3v1A81/7qITOmVFiNW0xnrlB/R08rsgsikwhkGe1JdqxWySzLqwXA9O
q5ZN0wUlHQeUuqSebaDCIJCqDpcU/HKkUSU9KP2vZBZR1RkjT9pYvtP3STrJ
LAII+Fs2DQWDPJg26vXig4KR34KtAUYAuOZYCEd23XRUKTtXCgYzn6pDDVG3
69/gi9EgMNl/9S+YU4vOrtLSVyMnKVq9LaI7P7+Wv4VZ9eKfy82kHgJQwiPl
niadjlJqbsK1DvgfxY3ZCaA6Uaxbnn7L3bm/SPCCRye6JKVLTPdcLdabcWdf
fQ0ixMOODOYv2NL6aHi4VK6sg171HLD4tm8Mc5ccddigBjRur8vr1XfVWSXH
vI2CvH9NtoM8k66VJ71pcD50epsucnN5w85PV64ofisT8m7ufNWwk2sTmjAv
WWwe3RSQiMuRRj1YV+tw5IroLn+/v8Hz7QZMNRfilM6SXet3Xx+I1nSgkQm7
JGkN9bpnPERTfKeyHa4ZKNd/yuGpfjtGmdjlb3DWKEbbZPNnYzK6JKODaUcl
JYOefNAcpLb6EtM+VFYmGAHfVIUNPcQL7Hnqzek+0RKG+ZFmEAkpyOQch10v
oTXnOlZXEQ8UpQ3DStrkks+ZoXVFqYPPHqPDu0nH4p6VueDIimD6Otgpj4Pe
L4Q3cNBuP9RzcQ5TDqmIpG0i/GL5QUcmyhjoqv+YHLclAZT4TEFngEeClwQQ
OG79NwpPROrgr89Wl8kmHxINTulzw/6XK1iBamvuHMDhefIuFLsd5Vmu1KfS
CwWW8LXT4uUr37GX6XT7MJBOYo6o8UCDaYnc8kKhjziL8BoBkhYFo34EPP8B
KJFRxOGTsUmupE25QbLSzfFcRQTYtQFMoUxqsT6KCx3OMqkrznSd56KuHJj1
NnQbXub6e3saTCO/hTzB00jXzRntH+ez/mYrkL02rhQvPwA6KXHYVr+6aAap
LFgykgPye1/DFALdQaW1uTYooCaY3xl1GmEISVS3CxdifjSEDrKMK70FSJWn
mXoPqrgs8LBakZo4Q3g8zl+0jKm1fOrr6FQXJCTTy0keOjnFanoVrrDbtGDp
7B4NjqB2Dx+2wL8+JD21J+Vna4UX2OCVQFeIMzvgK6pGXL2YTEicpkrZJ8Ir
UQ4CCVKLqa8knU8eO7r/OFWgLixguHz0seSQ4y3TwJmGDMakYtpXiuGSBPK2
wyRudpbZQ2+bs8RrNg5DdmPr+1kH25PEY/w3vPiKC3lPoV95N4Hv7xqBDXoL
L7H6RABskrvihZOGET0ca20PdnkC2hYEEcOQEzLPnwtRoDsrs02uD45JKc/2
zhAFaY4TnrvtUFnlwT/loTU/BMIGXJ3rqiHNxzzN9JZPAMHnIYAjtKmxEOoL
z1sZKNCQLYB0D8gIOAPX+AV6DGcZwZb6b569+mt4xu/evt/wmWZ0qShxFQBe
xMEzCAroftzMNhwqhHJJzvPOlZqVXXBte4AtCGhHzc7di0F33B+ARIb8pHob
SoDWyTQD3x9Zr8rpSomGPWL8Ep4bx53C6oJB9oGvScoe9OU5pMurstY5YC/V
qQ8a0LfblxO+mbUimFMQK+eQ1fJOhqR+9oukqbPY7lJclDUR3k3MYzAkVfdg
0/0NLpNZ7cBhAzkZ4XqVeNvle3AK3q944ejR7A1UxqIKbZGN0qTYaFDaEgev
ws6r04+eL067l03pd0mTMmQBQFbGJfR2hJoVxfL/c5Msq59FHzcybuA0spmB
fjoD2VHZwoo+ni0JQaZPEoGTAlqMHHbjDeO0JZnZLDdYSNjaxUmbQh9PMfBk
od2w5TsEDo37S6/oo4kv22mDfVT+tMKRWiAwK33M37d+z+/rqveA0USE8GBD
OOiPy0dG5YJT9CXg6GOHJGQPBhd7j1ZVNoPsCUtTzUpp3YvIa1CWFZlDFyW5
KpGXW7FoMEfAmkknCSEFzgMj3M0cArUJ89Lu5E6NT+hZLrARweQcaxNbahoD
HUrDQ93nKaoyqA7r94P+y++K7FR34QtCSr51NFrzwuEYWBrpFvtix2V+hLi/
cEVlgedVvnYFc7XRfvBI9XNh9T63yvyoe8DwCwyE3Ez5xOM0gwL+Thn5KCSo
avb1RxmzoLTnZvYuRPUkNAD1XbiZAnt7OxFeEKhtbgY2jNexO3lEtnUZJpwl
jrvsP/bAEprko9zIk6sWu6tv8GuVYnDyml2xVH4vRNF8dXXxXVe/9yasGU/8
Ut0WK7eRZB4NCDwnP7ijNZnQTanJ4aJQAJAw/RHVXEJDtXBjbRNZHIXsPAE5
90WHbzs2AdiUR8aLvFBH/Yl0uHNXATcmHZiI2ay7oHB5vGHtHJu7TLmUW+yg
/PiDgRG7LnI1lvsUkAKDfAeJ+7IummPp2QfrhOqoTcAW1mHVp2zlI8zM4pdp
s0lg32IHPHR/ng7sE/8+2cGn7IWBquHnxw69Zx8VsnDBZ+5wXsSxSIklOXTd
5e2KMoM2HSViPmv8gPyQ23iFs2WNE8UUjIJ7Gqj2Rfspq/7+RiLUEHAIoUy/
Jg16dBRrphbxZ4c8PbyRdaByHLCgRQDRzwB1GM2nPt4tiQ8DqScGJrHV5pN9
LY/hrjH77ZnwUbwMjEZYa/BElmDCf46L2Uhs6AiJ7nllsNq9SKDPLg22lhX/
ibY/ng7cxfdGE/v4S52Tq/lNO85Vb8kMNh84+bQDSJY+Pt+vVCqxMKQ29cZ0
rP/aDAKoZfLI1zjcz7gRLSIrSYavwgJGRaOf+KAIBiDeDLZpuVNqoTnhdmlA
aW1dMFd4A9ewsjZcoBKwADn5AaljlUbw7/U/8FS4kH8z5Er8IbwPXvFISgdx
cIpaQIqynG13MNAkTy/fVDX96Zk5bgsdALKjgPcM3nBToRK5SoNGjpMl33/G
Y2VTl5gpBVuwJNY6VlelJN8nHzOq4Ph/c3lXkWtddARjyE9/lHgYy+MyT04z
F8RkHZZog3wjMSf6OloGKdemB0gaLtvJspBaXQpYVzHgfNygautOnBfci2Tc
ag151lS4x4ptFfRdRZ5aBgPMkHh1rH6342b7UQXJyn09JkNOQWfZPLUWuV01
elUzzgqoagXSAk8Wko4ByR8s5WU+ZAtmsfp6jbFA8mBr2tm3VwKfpBDCYF4R
KdUSIU7TSX0p+wMnChFTl4EiOZtsWpKqZ8YKiv9RESoqEPW8ZVgIHpVGj991
T1sEyl72rk8EjHvBeKEaGl9GTh4Z8JInTkx5PDPpQ/vpcR9wuNgotJsOfmEU
2AQBbmZ6xrpxJOiRAav4WMM2svG+kgbLnfi1OuWixtpOe8hfhX+5X6VNGxL5
8zYU7mbk18DeCN3FWrlLtAHPe2ZzCqfjFwvYocw9eaMvuWtFGuWRTCJWyREg
m7wPIaDVyASoryq/nJNtYRy88DG+UmDs8QdmcHglAQ4Q3Q5BLVA9Ci4v1eW/
YiFUnm7GZlG0k5clXpesizmiuEJsGESumByrUIBVZvugczv1BrTR347PXusc
MiSEIy0CpDkXyVnCpUfcMv7c5muO5hiokzCqjV7h6F6+plGqCRy54U7Ry2kx
1K4+Bakm8ik/HcfaD8LXzIcR1PaSTndDkCFYAA9A/pRuNc/UYbfUOIfL8gHc
pcU2vdL2un4RAbUbMA0LP/Jan2JVtvjZeHpFsvwsU4lvvFHaXDgK50LFauHQ
DyaRXrXa1vLJt/izX38fOIqid3Sig4KxoQFIX3k0IiLQTnM2a/jwCAY0hN+k
tsCn2Vqvo7TLrtPPTLWpPnMflU+T6zT5paBnKKGK9qOEUjg7bjyKKUVcP1Nv
HlxY5lRFFl+5xA177BVbVrQKMiokw7m4LtwYLw15gb1n1gs9ZrQaxs0B14/q
xxjwRxvcgj26+UH/M8Ku4YfIwWbm4g4pYkmUMRsNwoM86ZCFgdwCXwoFK+AD
vfxmXO/r/c2VyIQPtL/Frf2mF2/Fn+iP/yOcp3CuTfk3xs/pWqqJ/lNj5C8+
zx40KiBp9Ko7LTfEi9WlWUvh3AWsEmp47RJlDe0xp47EP312EJ+37t82HXFh
sSaiFd2BwLw4o61+RHJ8TVQ5wGRtpaMWY5qbBVRhtQm0KfOJHDYARGXpzJMb
tqBEauTaRsaniVCJkQe8mawv7Cxct+Hg0u896ZnPMySpV1c2OQTRjdmwbZCm
N69ZJdufBTNt/bVB6SPuIT+QULOxdwm1Fx/GL+CP/dqyqQNRMxGR1617JYx2
cCopx7Q9glAdeZ8CgzG/LOMKnq7V/vziBB83T/5vjWoSRgHrI0XfG/XrLjKt
nL+7jxWGE9il8+UgDfnX8JNpCoNNc1CAcXB674bifJxWialE0/ezn5dZJ64Z
Zfe6xt8rYv/WKStWPtJezBB/xKc5Q9JiMLXiPJzGYAmOsUNSrWkR2eTsplZv
m1nLRZj4zlL69d8bm5X427AmW+sQ1u8uUuYRn9jEoQpP7gmAGBVaNLTkAoMx
iRxLwdlZWtlE8/M+sUVd/N0iykF2GLcCxJCmwUXr4ymBS91nmthTwjJfzN59
prXlfqdGMt8QvPRTFxLnDB6mhQ/YOhN4vpUcxULJRcYvp3ShFzrsIW0LKwAT
edQeC2uPyEVc0IA/iN2d6pECrOx8tKj/B6O6KYRcKsU1h0C+Xh9S/C/WbL4Q
xuR6TrDGUdT/w/mJYX7+cRch9miR509GvayZPuQJ/bo1xHynZgsO0R17JF2E
dqy8+ONB1kd/eOZLdWXTRB8Vh4RsP86rU632EEWX+oKo5rxG2d+mZ/pdXm9a
jB5VOYNRKT0dWTTl6UK+W6cGjixFtviV6RDdu7fULqSX7ZHc27QaeevVqcvX
+1Iq734LWqvi7ys3iiE+zRKOakzkbf4so6Jo09To4ZfLVnt2Fdftyh6TvKzo
kbxp/TjTNepqWa1Gbdg01/CLxIKZt0N2NZ55RmZIOkTguEPFL01bv2VWTAo3
KBCRcA5e9Wl25AvP+hBOqQEsLYDUPwbxZBllKgmw5sMr2wBtvTVcU/TNnM8O
yBXseqq3TiIgbfpRIuMLqdtfsvtzepkk7CPWt7+MsHIuJqD/ntos9pIn33Vd
n/kae5DEQxZ/flH5ENZGqEu6xR18o1PqCypsvGdLKSHGrd3LVijRIaGkpD+5
lNmqO0lNVN7Sa9PDjrOjFgxAY9VHzep5C6fHXuYRkYZdCK0yY1RPmEwD5HBU
SJb30I3oCdFGKSxTuXleTPMBlrhtEWKQarZM6qOd4qqtlHsfR0AWqcvn/eoY
7/gE8I1mZAfRzgnqA1tzE5XjiRc6Yxp7iMShbjFoxWG8zXJTFLMNOFTn9uOP
gjoX2dLxhWTJhQahUWIG4KvoIpXIZ0UHQZU6JBxzXIJYylhtznYsawQ1Kp77
7+C53G/wepN0YkbhvYg3KXLHi55XhMjiB3xz+GlTbOnh7ypqUI7K8EN+sQSM
enNGGPT6kiBhNIsGnrTqpEIBWUDwmknqeoTZ3YafSVRFarkbjf1z5q5bNJTk
9/hOHr+0d/V/MyAMoNe6X5O804tjOojee5e3Rmb7/kW3gkJoV5FPgJYW2xmL
5EM0SByIWB4Am+qRorRAILM3zZlcJ871fmvIAh3piSaGmK9uQAwkAip5JsHP
8fWRlKKB0SmaifuMnBzjVS8B3m2GrcUqVOIvcJpmsxuV64Z8DMsFgHgF1a+l
yVvCdIZlupsu73yL3HCvAH1KacuMCXNY0XXIcpxPbrQvm5yWYariL7cXfc1l
8XfErAFNiJuTXYQiRY9ZMgK8UEGAXS7h09jvKmwheJmw7ri7iBcCIF0cfROG
Spmp39sTlO2yYLyQ0fKpe89xHz0m+k2fM4EbhztXM8v59hHcyfkMIj7DK0sE
7Ioaq//Ja0R6YC+Pah24KqOfrS05cme0MgJ6Q1fprsPgsLszimgauUKjAMlf
VEcNy02+2kL3nJgNAD6vkjmrBoJltqUeSQHIybah8JOTTRUal+04QYF9NVCH
xU0Wjck75oaH1zOu3FnJSv/IItZO6TtvHhMhX2bXdQ1bWyUGyB3/1R785DCO
vFD6Yq0Hcg8nCSEO9AB9IWP2WbGr7nk0XXq4zju1udJOpbdh0qVuMrjbWyv+
aMUC8RWRprGghCD9BDHtK3IogGCVCFWT6rO5cfpI9RfCid3JJ4q/caxmbrfd
p9DVu6XEIoJc0KMe22ydC6PgBq+UIwiqDgkD09K7xrvaALQ9N0PwmgCsOguF
lGBuYNFyTfW46AYBxjEwB4VVYUIjeprceug3BDer3DS4JSIf5R20cfjfdLh5
BVlyOS2H0hEEurdbgY7uNEfFvucBPe98sOfMtQAU9szPm0Cb6+kGCcRrDrlm
ykDhBCOKdfBHXdNuAGzFyKaCko+bB1jWYVPenrE2afw61mlWB4YOoxzN2qbY
st2mtt4MlxS9ya//U3UCi68xZnaqD+RfMtcXH3S8oFRo17btcdsDMeJsTpnG
RoE/nOOEIE0aUMMpvpsSueix9zfJtwcpsCITLofAuB4uv30lW57r6R8DH8Mm
2W4Ah23xqg/17BSsoQFjrOWGg4N+57yP17BHBe38R0ASn5vxBBZrzQ1uWYRB
EdN82G67tk4g6f10X8C32mdg7UxVZLX8pT4zBkCowQ5qVW3WEVX/SOGiVew8
AGjmSrQgMbTn04U1WLLvA8nqs1aE3g4A8tMG54Pg/B0+v8kjpUknQpd0SQg5
zSB41odWw+7ZZuUqxnzqJ4IEwgLpWPp2061lOF2le6fKZGKs27QAYmJ7gxVj
9DN48Km6z0ck0hgDH7mhYX3OPQUrxR8YCFT3wq3gHmFBnry0ex7P/5k0e1fz
sw0ba27m8svDGZljshSpWoMyKE4bKhiTIjrWLJ+0Xk/FMo6YWYElJ02MEwI3
B2rklsOkEfKBi3I8pehfMzNmzUHbW5YTvi29iNKLbBHXrVjWvxxImeRH8sqJ
7+zn7R9zobUhuU4BjScnAnmbC7lUBNBTgX/TMfhuEScmRplhznJ/Rd67K/lG
3nHSm9pY6hUetL/eisjKmnTJwIfcSOUxfa2b46fx9X3N8Vf5fLxGVL1EK/Nz
RhSifG4ndLKbMOf0JO3YBsFJRVulkNP9CjE7zt83vI0w4Ayl8x1fyx/O7sJo
tzqvd4FFbOp9k4cY7hhaIyks/bjQoKuqutsEEOubMOTxWSb+lSTBfU/r7Jcy
VD/8bJBZGnhglvKcI9hPplgn58A000f43BJ32nWYXAE5JkrdPaUdhtib/dZk
o6tWBbnOK9cSUk0NaoSviU6Nm75rlJ3Cy7enEKtXRaNVjl3J89jfK6KEK9g/
WvzTHQODRbQw9vAHKbapVvV0y4dDNmR8jlF+fmtXXuY2ypZ4ljUV/oOKv88Y
D4GlrQxPzT0g+u9Jq4Iyb/gvt/fk1+wnN8gTnsUkovBK9dfee5ch4mipQYjF
AXfD1iqDq85ITL+fxqo/Aac1E7Thrf8ym1n8ReqvNHGVw+Wzy+KC2i5vzrcP
Yt07g9/3BGCfz5bc42rijOYlH3+bZbxXhx+D/+LRlh3C8qisBeE3YLa4fdl1
aWH3RF8R253QrjyqxCSaL7JjVNh6243QawaC54LFf3rxMP0qMvrcWdWIxNTb
dvm1SllyFNLvvERIrWqmvEOn5EjwiSkEajhRCKOTvkeZbOLZZ5/QNbGSbr5R
O+7a/ONtxdQJWd9tswZ1f4q8RjNPFccQuw+ujQ4WkEwZSduaotMQL8pFXKsJ
NjdXqnDdQ15loWYv6sH/KYtw0Sf/DUh421JxMGdE0BSvSRkpxjIWqKuwTsmn
hlYUGvke3dD/2HDDESYie6MMULrBHwvpIBnBWmvcrDXozxxvw31l7YGpeFSp
VlOwFX7Le8b+f7BcUppkh+mgQiDDyp4pip3fjHJmAsS/R4gGD2H2PjULi21k
8JKOXeG6hWqAK9lomtCFV6ypEWPTq6yCyRce1WgQcPRdhW58fS5bkRKrteRB
NLwnXQhskNxbW5SbBwdZoKUWBQrfG+RiulGu57PpCM8Y8XHZB7n2xH4uqR6V
Wp6Lcbo56cJ7Zip5KMDtXt5RWNMfWbf1bFX8jdub9/5pEjlGQElJcZV8JrpI
7nhHKb41uLYHpyB6ou9EDTkM5SczBabRJpHscLlXgbAGy3bbtF9tnQMC8VnD
6bOgoRUaCE3xBw4rQkp2JomePUTcVfX7/NeqNDPsjxD3SxKYtS6L0R2b2BpZ
ZSQDCAhHAk+6YTugDycMWi1jHddTydKjMqsRT6LgEo+Ja0JTiXJEBuf9ul1x
qm9WhbQ9ZCd0tgEzzrObNxLWCedKxZ95oJm048c7Acld8Kxq1BXsTspGEOrf
y1wpjjOMGF0k5V1FLx2NSRZaIjR9/VVfkTJug8sre/VNVwVFrLtbHqkiP6DT
gBdxDBgNwgSTmUuvjM/4OL3VWKOb5QwKOJAb+o97+XlHFePA7Z7zbwwLNdIU
JKNuwlZbyHGJ4RY3rfL4JlSzMD9w6NSLvDyNKsT8n/VsYuFR2LZjHJ73I6Qq
IYMuIaxvkoCYABO9Gv5aUoJS0hBioQN13CjLUcPsuaFzzxqax0yYQ9vBDqwp
VA4mtnK2TnrKRsnefRBwrmiNi2GN4KZ6BRuE8TAqr4PWk34SYwYb2JKii860
S7hctyQ+nH2f+GBxOg0PdtaTJ9GMR9/BEn8mU6pS2OL3RI93ivDfSRgch+MR
VzGcCvHkw+XOIHYjImKvGCmfrq8i4qu1oFAA1QzodFBDm2DxAteKDPfHgYMG
biXT2HlAdFZnJl2MkQpexHrtu3DmFDURlfco2WUKCO8eQed3n5WPCT8UfTjN
qLWTlhbBe60FYSfp7kwaG2trfv9nHO2SWT3MItN7NooGEiCPt3xjDKtN3u7g
ZOLCBmwfr2fvOyBtGQ7qsSXqenjBPiSv9yQ9pWz+AmgjkomQ7V3Wc0tls3Gk
yEJI1c2SaZzth79QNAbEfB89OPajWbcWkERPFQ+Mt32fpePh1GcHu2ouN28p
hsAK8CIreoEPS8VoU0pm5JMgR41ka5uUw51lutDiUthZ8SiuvtQHvoDpv49/
S8i3qdyq7NV9l63B2nSJhOMLB84sfHeSd8e0zOj/r+f68YkMeqJ5GWYhBMiB
4vvxK8HcXUgjlCRuuWCNvf75V+gE+kHKscFy8TfCvAujdDDj3HDXuFuRFfac
qqetLDdQrkr6P9obUBl6TJYzrPKjfZ9mgwJwKZCxCNxXMMrJhAJssGFwbq3k
O2mdZMXYtQAWH+6S76y6sLtkf9bfF5X9YD4TSOgNiE1RmoUndAamUXaIR/zu
VspQ5FwDa9WiTaLVrNVhXDCyR1mY8vaIjtcDNxAgzewVKpnsD5DGgHbAXHzJ
mayg62udU5/dITkccDtyd90/NoPa089CMtUyF7tNouXDiy7Cxhs02YBg3lf7
clOBLlQyD2UxeWC0u37RD5rTrnj/O+uz9AZi7VFT9UmduyWCFWlkPyw11PFB
WDsSYu4qbcT3M17cxryfZ05q4GcE4UncCC2smyzzN4cJA5oZbmieJcL1Blv4
LJFqJQUNTHpHMlEhX+p1atHvzRbDvIz3OVMQngun8mr4v1JABQeSfIruWqSC
zQCqDlg2/frojAgcffox8JnqMaTZhpShHniYYqxWJeqTSKQC8ByMqonET4Ha
l4j1cvszRcWFfLaINQ3q7ml9Q48ts1NeH+u8mgr3KQ3hEcRQ0tj9KBlQ1pgD
i7+hVOC+v1ArWBVFeOV5+RosJIzhzEof7adGRf0tGfMHx6oIA2TE+7SSHpfK
IokUla7Fjp62e9Y/ISG5GyW4jCfW1XmMlzsCCjloZSXuGbvSmccTbTr8HK+o
sf3zl9fBG9inOXrNSlENLndLAlaNcBbUSKj64zqARXDp/nm8JgA03CV4h9r9
lNubHYWg+49OoM8Fh0BbThGn3UOWcGYYRQvpalfBadsEKGFMjL9xYvkmIofu
efDgYYsbECpopPGt1Pu/404tIkVvXAXVEYK4kgg1F20/bx2yrKO/Vfj4lpga
UmInzcdzJD7V20jCBfdMYATadWQQrCoRSPeF06iAd6VHbdUTj2QmFQ9arcib
rkUrMkQNCjbOBhBhOJv/KBPioYbRZGQKfsQp+YQW/rafMx6mrhXdyZ5sUT6c
+Flq+E+xsiIaG4JdsZJtFExc0nFE4eVgfbi3AgboG13mKICDPTKj2SpzXX9Z
K1IlvLxjvnE0TvaIjy1pe+XA4bLw2JCbgcEm+mkFgENJEsutQLDMHKZhBrgC
bQYKD5V1UiFEFio1CVk27XB7zO1k214Q2kgSkFiQTsxJAkak+3DlkslDKYUN
WVoE6/75RzOuNf395Xo+U61H9iaDdB92v/f1+N12jOokQ8qp4y+eQsbSXqt1
dkSJszOm5j8UobyKgsWU4ycVJzNJnHAHO03Go71vWCCMx2YOPCaj77uzRLhQ
YhY1BFsAGxKZV9TUGo9zbPsb2sBepmRGTANnwCDBKNgsL9suUnmEY3j2yS/m
ELn0JONtwbyhUTc0vABN9Ub0p4pTw+eLfLYwUEcBDzmfpCftJzM3S0LXnBqj
9BwMGRQAhbwUjDVdAXGBRYXGw/WME6AfBYDPDL4BWSDuJbIX1aoZcu3QDyc1
4XQ+4q7FMK5tGTb+Q9qVsmrHpuA93fz9CdMJLtLz8oBiaBG2rVNr6nHSFylH
MKvkEBfM1bAZhk0UHMsu4nXbCtQqp8tJ9ESOwiXtuY9ASZaDTye3c7ZOPmOM
X3p04dLQ7+g9P4YMPt8sQrUQmO5jRShkEN1NG2lI8iaohDlXRpD5LQdVCPjN
juKjFg6iqUtzITnqMsu08eZRbMXFMuU+4Nozr6Lxwz+mGpWJNCwYM6bt8yb/
oDc9AcauekWK1QBJuiBGLlYFuct6xd4jsKBz8AdwW5spZR92Q4kxRFxqNhN3
A/iNn4p216RaemJhjh1VwzNLUc7sKhZ4g9lpmNuAwSmfl54GcNq+xzBIzt5R
lfjBnR+F3bLFly/25JuE8EGm8VQ0s14QPj81ApF73CKr+2ySykBb0t6k24MS
eNDj8Kti1w9foDhFsGHv38Zn1/EjN6+5Ru/Zmv5pjtZ5GibAXXojAhRfnp6h
F7QYw653Gcb/c3ekwL9M8pkpMaypHz0JFLJuXoL7+AVSZFxhLr3UgvAmuE03
5FollQgQh/ST935IJRG3kaB2p3P9OrqWuBB3ZOjN2hIriZ+YU40D/9cRuU/7
GfzDwZ0EpUFTdLM95xa2VmCN03Q2tyC2hcpT5/g8jKEWqyZOWiuVXwMHDZf0
p/KfWGQhLR0w9XArRzOEefeAIf55bP8XWxmyV9x1MIzptEesixKEIN6/rzlF
LNDPIDpxUz37u+vImDMivY7P4Z3lEBCg4woPtRtSqRTGhpdJ9T4asPTu+4D9
DYvqHjtg2iEloc4HYCGF2iHRcSGPqAH28sADQUZXaaMX5tctVd+phFwkCnDI
66vcta/CgRBQ5DdLT4SqAJOoU2Q+qyympLXaIcDu5P8XzSsHcjvKf5a3toJE
4jcS9ZWPG9AcNIoJd/W7Q1AZvfoNIgP1zCeULqsJLIX9t8G2xfsZiaLJPwrB
sKNtDKPHrQTjU2KYspQ4FhV/NMilVIPPh5lg9Hm3mC+hCAgVkW3K7+ZS8CFJ
Xtf5Te2cV5bx6jDbg6dJXeJn4cLpVkM51Vl1EYD34R/EEegh3ka6l4fHpjWt
BYwsSczo1up6GIN7EbawBwSSGWXTVrV2C3HQ0jQmh3gdeZmwUy1noXHWuU70
JW+qzzb1IkTortpitHX+AK3v0OJRjTtk4LU75tFJsxkYHcMIRDiSq8atoBLO
opda/+qb6G2ckP9c2G3Eij6cluMasFT8XKrh++5AfxUo96MX/0LnzSR1MXwq
WnkUgioQzYtpPm+izI5XJPFJGrdbcU4ZpDnWXYPxVvS1Y/po5m2ITeWit2/0
zkrEXc/CEo9XQh5XQGil8+VyQ/ruBb82PYcb/k07BFQzCGygxSjJqamn1Mjq
hk9aIl6/wzC1K4xp9w6/K9jhaiyM2KaVG8jJauCLspnqOVyi2KcvDc7B6GUt
istwyHIJq138y1KIyGpne8VpLWKegdlUu75hurkD8i3j0XjyJPbAtjDMXruA
mywQRXpRHaeHjLY+GGFGXVMfpQ4of1hnXNYgOJEPQZ2L3Vxt3aJhBQkYzOaS
LPOMi+dSUaoqdf72RKNsbsEjR1dX4hBy/RpWDdsdpeWLSqDk+5uz8jdaaylH
DXEVEZ9Rf7HIpi/fH6HppWiWn6m9HTORfUSNf/hl2+eSJBLlH+OFZmqTq9I4
y/OrZj53VEizk/Mc+ATESrik+Eudo8foDJiqdJdhPsDwZG0G/QbfNeTSRZ1g
E7dOf0HCfgXQmONqCAfpNxw2BoGmrp2OvzGOoDKhdWSuGHHdANMZZzBoTMNY
rlxMY/jKy/pPEw2JWmig1xgvFZY/Qg6BVvMZEzmMvn0DszSCk6XPDIqpul+Q
EUe1j60UES0Y9VR2hFDl2Ql8YdX6c0dsQmOSuOYYz0RLHd7DGcmr8SI3CglR
rxWMJyyzXgn7sf2WbsgiIFyJwTi4c+j/MrMMZVPRxhDqlOWELf9+J6HLTnXe
dH79wQyY6tRuLKUmP4A1NvcTsgLcE1ATO9FgEo9IU9o7WXPdlCAsD2Y0XaWR
lHTGK3k2ssdiR7YovAwXrl74X0dawIBVENznegKF0XEmL/f2/jc7q2sXr0on
Yjjm5tHsAo5hJ/ZRIoW0ncIePcD3V2MtpFzzNMY+jmCIlK/yWbTnAxZv95Kc
QlaZqbFw6f2Ljs1szMpy9M16TctC/hxqu+Miy8nUcRV+2Izgr0Um0dz61bCV
IiZD4QGIdnHKZayOAMVSc/A2fwBQ3Qv/rkdSKb/SguHtjWnlPYV9yoF7DfKr
wzyxJ6IxlxIm3zcC14gaK67ebnHUkDaHodJ7rVBL4tk8kzQRBR0dZiA6jXg8
eOwvKmzTfhNPvs4WkfCn6V53IrXrb8fMAjqNrsCtkwfAJpp4sVzR/HMAhDmL
gZhweNSSuiFVq112wJzqowFWo/PNOWisgFnTUeIHV/zVJbj6gbWF4EqIDS3s
SHb08VyntiEN5lg6WpKQq0mQ+BiKTpnd9PxXQoo4DmX1LazRfdFluPOtHddX
Y0GtaodKpsFCPmk0/j1zYK9cSHgXTIBwD+p4JCSoLoiN2SUZB+NzJTKESSnZ
9jwje5h2ySp65yhgxeJOh9WZ4PpGWPW9xuQCdLTv1MeFzCt4/AF19294yAfr
EGcou4jT5AuXvtGM9hlT0g8JO1CNSodvFCyuUJiYaupf4ouC3nRW7gbovfDy
jy8vIKdVhftsaeV3wetGQ6BZGCZdPJqZWO79pI4vNe+ZU7Jb7R4QNoNVmrlC
Z3MLZMcg0pQRRQ/jX4zzFTN7IYfSXXDy7o6+aMH1rP6Z4Q5h9TS6mBEBiafi
AfJFg28eADaMIiYs93HTDmRtn/Qb5Uhox+0dvYu/xEYAM9kN6gxFeApLlbem
iwAjg8PNxp/+d1ESk4iB8T90zzVCfg69DQspQ7rRXKx/uEjE+OkREcJ/0xiZ
sj1Op1na5li33+gx3nBx2/2wG+99cpN59tvLAer/GxvBwN4s1HpfKdyw5Bhz
MpaE+UC9bV8CDmkwc7lj2FTuJGh2WUoFG/XpZKsg6lULXvvaNeRgr81fuKJR
gwwX53UBfqNrXN1F3A2FFmnpHek1S837sDVzHp36PvBq/Smk2T8TRtv5yPpR
xrojrezxG+5ZDIIWJwmDzITp6CgfV6pbFaxxEw7XPZ/OliPJEYxlaKOvcPTx
OQO0VUJz0IXcDKs2/Qd1a9rTXvBDqCAI2pWBGeGEGjVQ/qkdaPHEvcGh1pu2
xjoSsxNDbbgkCIEDma1Utg+t2xyTSjfrAYLRK/8rRAhP9PUkRfauSnK4HSBT
yAQcMwP8hu6HilPvQKKANzV3fs1x77L1GEj3HVTOr6XFnP/9Q8HQtehopIZJ
r56FS1BYq0SmNA2B36we14CaJc62/SPSiiGYGnGbWxL5YfEl/9nndeRWFESR
BiuKUBdIm4uMHObd7qKhRC4uBhx4yI3Ftnov38xRAg518CluizV86m1eKP/t
F6rxwi8YOpvtWnXxB0/OBCJhDx6lFDli2x40llgnxlhbvigBg/9d2sovyGoP
bXHYXgwK4GYV/bfYwDs/RdWRmu8aoaeyb+1uwqDscqeNyIZsRuCM8r4KOG2T
IufqeKdrEDo5Bh/1ylz90Oo/5JBW0nzqL3uC7d/7kXvTwomIZ3b70zduLihx
hnDQ9xOKiIDgPyoNT21b04GoPoQzo5QOgHrFwybnPjpXWkkU7O6da3oYqQhP
g2f+nDJSe79g0L6r+gK/TZHxsQTdhhDvtDoSYEJ83RIcYN0a29oypeVM+/P3
d7Fo3W3ufWck+uYKj5drDIyYkXvjglh6bPDTOBYpkc/MIIsLdYJ4EDRrwFz2
erJkb2QOmgC+jmXHCww71OUCwn6+YWQGi10L0kIYc6Ay0Ffr7qYAkLBUGX35
XfldtXWTuZC8d43Y0CbmY/4GBjRqMZjvX6GIw4mmJ3RA/0s2DB87oJjEYBRz
XSFDeMN3vsIzHDHBbrJB8f+diFnuzVS/06dVDy7JWJb08hjnQSHYSbAS+ifC
MUwcibTvn4CB92zOOtVfFHF8dxBmVenx2XGrI6ucqhNVo9mLdexJFEegjqMG
QFPiKwpdJpMptWHeS9KuqGUGksDcunlQq2sS6YhxnzUkc3juL7CIDeKIUV00
jVDWrbK547tmbx+zHAiQKug3W6ImZX0NVMgUO/eRt+D+QFm4ezZTxGbbj4eq
XWPKpm/XlBFrAyg0mYnVtxjodauCajST0lhUrT7juzYochXZwItCO/OGBJ+z
4v655LJVchREtsLLYWhjxDXmi90ZaWJweyeBfJWEWZAMULgrO/b9MiSL6bC2
3pylK1y7OGVRVMRqtFLKvEO+VUrswnJHdCe5TeWWtb1R56YryoOieebHOCu3
CWSdOgbEc7Uqk/gjKzz5QTKmHzeYH2krFam+xv5hYr1JQVHn1+5Da30QI+zl
MaXrfQ+oCP1x2g/lE7NYyxMks2PYuHyZlA0n8RSi5dt3m5QEX0uwuE0WpIq6
i4EUHKbjcjwAqXmyjbzjf3m7neMW97JCNza+z+Jyz6NzPRdLj4gW1plVasCH
9ToX1docTJrCkcsyruB2s/kZWQxhh6AaCu6qWIxoTUjCMyAXdaoKn+mGVpL3
nVpOiqpmIsGaCVtHefnDlQtpuMdNnt3e1GAHHG8uP4W+U+N+j1GzIeLw2TLu
OzOL9BF2DTXpk4Y2YsVfuVrwcMqEwqDrVyDwMCE3lybVpPmJ/6xmXqB8Cvz5
iuADw/9ImwMUZS0seuwTyJH57r3e6x8I4c/qVGk4cmOvk4QceK/VWLh3I7zj
K9s4BB4/lf7ljxmULXhcFTvpCpxDXJvZ73gyEzSJDOndm22VZJj5IK7MEbXT
Wi77u3MHd0Inc6+qP3Y7ftCyEu75JkybiGHEiWG4tCATmJCdpsRU7SxRvy7N
5Guq0/N7dE0MDQ8Cwjp8IBNbNai3kl4ibriNL4+v24zxCn4HkJaniTvXu+rG
RNNI+/PTtM1sJD+VQb5LSZDcaVX5k/4NTHocAUqVw+ns88He3d91KfPJnnCl
iNw5A4JCp65JB3jfo6GF8pUc/Fvx1d8FEuW5q5nz17CrqRJg6qsb6sse5bzw
JpWVV5CbklVRd4D0xfwrvFvw43kLUiXJGBOdgVbkU4k6ETEm+nruVoPysPBe
kXxDQFifjCWq/PtfpSsbjTRIztZioO7YKLOiYb3fbBQFfnG+/N5hEPak2D3L
0yb/64TnTy0gz/rnhDuPG0EDj0aM8sfDg6asOD2JI+boD1tVLtxbrqT1b0AP
jsZW53PuStmW7pKXRnGsJXuyR63/XsMoNGp4V4mDlyW8qJGB37Et1+6sfW17
iwZPXS7C5pAaUDZf+OhfVk5REWXzEYHyaMvqId7ySUNKE4dqpdX9D9YQleT0
WXzwOuxuyOuK6bu6gvS377nC8rRxsVJWh2e0VMuI3vUBjMY211IZqHpzZNip
Z5+sYWRMh0+ahTxC/Uum/ltrqJI9PY2+RmCL+OL9M0bFqiyEqjCHhPKYtGPR
/q1NaKTQprN0ymcya4mbJlK1vlv/wOMoDa4/S8kxxf4vIZv+JjT6x1z0J0dL
Mq7fmp5Ql7QEsxioEL9xl55Kibrc8xMGBy1suEHxdxvJxPRukro9h/UhyFdH
zK+sS0bLX8/j4w8mkrQojuJA2TNGUhRyVrIoJJc0CBt2SGUsBUkqju1QAKqv
wlNvSN6fivFrkwWVvrJIS8eIZlmXW0BYvLlk1xT0tlSLdcWnFDNeBkhk+ZvM
a2DFa+tozdF58k88dHMEqYfoYOvmcE/wHTcw3Tnkt1fPouHetXKbfVhI44zL
r9g+s5tXlm1MuequtwMR80QD3+sz7KF2dgpTJm49g3UnslNWBN0whsXeQK2c
FYRTopryUMRIDtj6OkWym3pITALsEsV1tOXKeXZdhwMlmMpM75gvc6MZQ6gH
T9BTX7Ff0Mf1QdVweJz6qiqDDihqMB0lBgtE7Ya8GIfGgfM0fUynVoeqveqg
lCKigF2WCq/aYddF7yWY6dSrwUlvyS7Q5SMVoXa5j5UFp7o6WxM5dU++Lcs5
YuSuf+OkliLLrGcO7awptsRBJJAZc+KXGvVChZEd1bkF0WvnV2T042a9W2zD
V+K14XiB1HDIeL+dtxNUQgX8s8/NMZDDR2UBRyqLBENrLFZuurEiZjeQSbSi
1HNo8icU09DjKTDworcLKj5rvKutWHFgRMN5pvLOIO9mzxNV64LuNcXJO2kJ
DvZlDiYBsOikapZl+nL+tUViQyCJNzo1DLZzT1FnVElpV/wvWIE8KtbPWW/b
JUSKG40DXT0Sg5cmpj1CFVRUN3hbvh1JymiwsohS5TJhzoOtuL5AXIeK4uR0
sQWfmfoij9NabFOSlVsnubZm3EAdBAYPNgxcOQ5cSMsEgC8ggxRUbahPt8qZ
TEmjmNF5jznOiwDa+vy/R/BdT37xByi87X25nyVcKTZUC0Kduj4EI/AZeQd5
PU/BrKq84rNyQOPgEDepyRgLE9CeBoAac3KwhkJP/c+PZYEEH3UKUvXUjDyX
hIwACP0FPFn9Kikxp7K+YZGm/6p2yD/Y9pf+vMyKny6OIvjDuKGDijvxIvM9
Ls9IQN7qC8/rXyOcHfm33cUpph3Ujk53iQDejJ65bPFhgv9ly2Ya4eHV776a
xSPF16b8J3ahVNk5NIml+Cvp8q8sv+CEHfVjw8iyVOc5suK02/y+0XH9HGe/
bVoPvU0AC4XfuckFclVEH3k2tO+afDiB6loNeW31JmQYKXA6hECThJCUg5hs
tU3XMzbFZGALRgT0Dxa0h7H1IZRTmXnM/Je8k20M1vtNTom00WtFZe8gHXG1
pKFZHIjeAWjx2kHkoEztJo3ftwNJW0o8fx85sbiu0iKnuItPCE/ydmytPehR
hpIfEgfvQRc/xR92FXZUoFlYyxa3p8WgQx/lRDaYZfZXb3lIqNrrS07KGDcp
0Ye4XvfHVaPYlwQrzBEPNCf5UZSyaxzktSlf0GP+DlbkFJqgyHD0eNTFD1TZ
YaolnetXHoc8LsfXT/VVDWSsLlpperDXa6hbXcxGuFx3wfWlW7s5vHHc0uYq
zJNpRc+a99g6p8tNAYk0NDn6TDW4hubIT4Oqmsxpj3B7t8lz3zPyAtZ5x9/9
8FqrjmHfJbElG0KYGz0+JXubUGbyLXIoiRg+hwY+TvPT3vWAtfLT+Tkfq83X
lP8vK16vwSjzE3h9LfU8UryD3h3QLNTd76oVX3jXpGAvEISmHrFXK67qW9bz
ngGpVgZ4DTIMw343RHBMP0Gisr756FVJgCqxcKbrUceZQjx5s3tlUwB6yiGi
Ps9NmUIyr/OAVtd8bqihMSuLA1fy9zrDJqPVW1dX6b8FZAwcvXZr04mG34e8
8y7tQHNz/rm6X9kR4x+E9mYk4wkylkqmNxLRAHzJl74KomyVf4c5udCKRV8w
b1tEv8H3yB/kmL3LQT4RZ2tMKw4HmCtdoCj696Y08xWo8KaQ2m4cffMtYvcO
F0m9izCjEoxV9rHNbRgbBAJ09bfrbG5DNtO7DFF76cZl1/JAppZBDeSuBQB9
qsKN9Iaw+hb+D1I94bUzY79RbRnhd0KUFSNZM0iXLt7cOLKdg3Mo/xrY0c0m
oX+7J3QJiwHuoeFTGm2tlxOs7Sae1P/Ac0Kwyvcj1NE4yryrBzAm1+/WRNBy
oLpUOt0GCQaTnxDEXp8jUpEiHf2Q3Zf57ni/tOGfQ9j7rdYql8101FCuHoGa
dulOPxVL3hdM+KtpkM/3bAXQX+TEEdn4WnrEImJAdmAWcPdisIR2cR7uS0aR
hcTkrnJ4MmJYL5/mFegdkfI1OPugMpe6vY6LjTYthInFWpm9Rj/+espJcwSH
pLjOMPyBRMlFrasPem9trJ7icWoWjpZ3O7Io3/WTedh5sTBGS5d2NIxIdWVM
sd9pzU6aKpmZyHEXcg/N8R2coLX7XTAlmcAt92MOLvcCs4GbIxcDo6I3HdJQ
Y4w8R3hOIlTi0aw+9Y8jltkl2yT31nCXW2trvVhLKdn7mL+6cTWqX5IoS4Sb
Zxh75gF+o2qaxS6wq6tDuAF145MxoODGgMvGXUbsEl6yTlF/o8h06rbXBMwm
EafBPUjm+QQQGoVWBKFXEnTSifURMsxmV41RAaxa2M471UWGU4IATDIWVZBl
aBxTF2aDjLYPscuic3V4ucugYSkAvaznT+Mjm/l4uKTHZi1BkFjLPNTM5+hu
F61y0rwqmStpCfLz3yhvqAJ1vcomK9XJMe2JRjHs9Ja2ikXv/Tmi3NXtw8V0
SPHKUoyJNET1iknZg6PPCTkPZ/H3LXMDVxyakH49rY07RtBld5UiqO0KM5TK
nVEtjQn7n7TidOcHwUupO4iCFdcKIIBOGkwSToIAe5RsxMTpKJI7ZHCLx+j4
shdpBvOqrfTnAxhXngfhKE5HW8EU+i1epIgvSw4plqJjcl6VvJoIxXsSxWWq
uqxEQ/2fBbKreGw1u7FOmN5ZirP/xXyHLhnULvi0IcINNzV/gqux1SxQqPUm
D79RCLjHnWoyQ1OUT4DkvKY9MpFc5ShuS0oY78HflLdK+222oNObtQH81igR
nbmoSmBBJl2stcuWghQ26CA3VZKbVM3JA6jTze8oUvX+AzjxvNbj2QnFEpxi
DRjtjoW9iQMOR/7iTE0pr1Joa5oHV+51wq3V1h13mg/yjeI/LEmWX0g7k4KT
/9nj8rHlBHtujzA39mJzMoONfDHhYj3Yh2GY8XaEuM2qKa1VFHE634+Mnj8t
4riVckoZ7yZq/uaSIsipGTRS3K160BpTz0n40pVWsjkGjz6ZD9R3Mlw62vg3
Fegv2fW0D5Jn/GgdfYr1ZwzZb3l2wxz/AdlaGXirOsu8r18ta576yNs7cq5P
HbLqxOZup+3tzSeR+OMsVrNF7zfDw8nk5Fr8Acc5gVikj4T9RSxBnT8dAnSx
8Ric270VVEYUD1cNm9Fhc7HAtSxyBxoo3vznE20RhLZ7GJitBP/CdSqtxU/z
zEVJbdiCJC9KA/0DK6wWEMxueZoUOFAaEJyFDRc9+qLmhY4gFGymo74I8Uij
/zMAt4IwJo8bOcO+A+hMFTemCte0OB/ZtR/WFQh8bwdQwul7CWygjg8VOEbt
egPm2DCcr0YLqmxxg2dF4gYYq8iEpBvR581X3oC+b35jQSI1bpuPM/T2vUu3
uoAqVEbtvbLiaGrO0ZlBTkuhmUozAK/qYpKldAvMGW+6AJnaroP9UI+dnDzS
h9Ei0VasiuVuqXnAVaBY4obk5Tppxbs2uftbsvAUHmAHWJMKJHDULh0OI0Rm
rkeRXYRinYfk7vUmF0YxdG4IjlpdtfINdFZw72F03XfOXyMs6m+Ya+R8ZjXT
GR3epk7vriTyKoy2tccyzIePzLSGl9+OtdbeP7L7FxI469KKOSAfw+D8U8fw
4mnRsfhtA23czl3UypShVAf2zS/KzRp0XeOWJZrGnAy1LTmYZdAbyDsxtEXP
fsPpVKwIcQIPQExI5OkBOo4ITrenqioKcczavHmTEO2vcnwHBo8opZooM4lg
aPyBM8PDjHYMGZuNi4yjIpFNiwt3vhwis2o7mi3CPSa+LWktezCCRtHmftF+
taZ7lx71Ts2QEiqqHfwRtGxqHd482InrCUIZRld2ZXdKld79h/g2ZAPnXIN+
HDJ/JfLpgr1zLG/fJiMb1AUspr1fLxm6pgn4OEVAJ5IMiqC6wFRd/VlEquVF
vBG/0tyER13kqkYeSp+EPB6YaqE8ByeuSkHaxaP/jihvk8QIhIHaG6oC5iL4
0Tdg3GQtMo6SXsO66XdAIWZtyv05tFDagl1mIe3Uo9z0Qs820J//kqAqXs4V
ZJREUD/BCsdNARdR+e71VHiqcXDc7vAhDMDgvR+c/6saCjDL7IhZ/Y7PbLCB
a3cTzrKIz1IliW7rWwGvkw8kw76Iqz6HQol1CQSduM5VHj3SY/nu8Th29J7l
w8qhVp3Wy/MSm/9KRteCnn/GgWrIU4dn0BXF1czXgaXg7yefsIYDqwSnD2k5
puJy2C2MdzLXN9Hfc92PDJmgL4Z7jRnbt42C21GRJNWTxzmwqkZRWaDGDpoP
BUJ5g565KhxfdMKn3tfzHNWqaOTaK9DLCItD6O/4cdAY50nUXKdCYMSChwSu
AarqU3xBCViM1hlDfEvOaICq0vVF/h2+Ji5OuP19K0xCZVqw61PRYP4YQq0s
sDDuRbV9TIDoRfr0B3VzwCWtx/zKTQkpqeNEGs/VhBQA4Yq1DmErIBTIGVGM
qc21PFQ3sxCpYAF0lnqFyqkrVSKJi5Px02KZTFZQ9sIncerfmPj2ysWD9E+5
zSGsxns3mR3QDnGykLcehzqTBGdHUoJj8GMwzeJCjFO5dBwJHZixZ/QfvNjv
tkwmP7At9xI9+4Vhsn1AmsVXY940edqG0n7iYNU6RX5o5G4DoHWWI2eu/TxH
Js97ZKymczvd5/2iIIGwrhnnL/OKK1M0A+SOtQ/Fy3W+Ae43d3x0T8+2hIfm
MCw3zyETROVYKfyetfGYkFBQI1bVKiIahuELA3UoEPA2T2ea7IMIYtVoO+nj
id5tCz6mhTUutGTXaCX0mKp+YD4KsHlFxl8x0dIas3rwCUbWrj6Ef5ODTeyN
xGru2jJAounq+hn1boKrRa/b7hy4N/TdC9MAPhLj9M5VBpzp6NePfGkdNMBo
NXbn/OemrrTh3iCbfczWG7in078LMQfow3Uh2PRTqcIXtWZIrivhQK9pyWJw
RWBtOExwwNb4jecQ8MDR3SjryrXORYAM+LWLgtgv/H7p1ariO4BIOp2cCtrK
GkyZ4DKxNzBoNjGavMSHPr+ZQ72mLO67RK5ZZH2Gf5xFcBIEVvxcx0PR0oP7
xoRqGfCPVUCENfFGyjcos5SyugUAWfeTFXIgrA6Cab+3/p2hXWyrAlJ8glwy
sdVdlzomJwuPMM65xZP3hCarWtuNFxPf0ZI58AJy10PNbRFTg+Zw6GXohhss
/rolGYYCp4spJ8dsrchmmFsvHvnlWjSJQK/+GNl53hCli9FpeATF0LWo2n/t
5bFdSXAMfBQdRXQNrz7JHX7gr1eOFuDKuKEem1kv5cSg4MxLPX/1sMKICGZU
23Xq93jVtKVA6in/3b4QC/6VUt4OONsxcFWsJmLUM0lOoInB/iCpRPNnhmQ7
wnILx/8de/phn7XIM8PYIqT4ke+ER42LjnUiVoWP751OzTP72R9M7FnEI/GX
c9XG/kHLsqhbjgOnIf4r+xpolcfTQu+LbhXib76KyyTMXATlCY720a/vx5VH
0MKZa7wcdcmzBM+O47IHQ63CuP0ze5E67P+ZmmvAAz+Q6bsd2WtoBuQQ8Ntf
A/VgvQQDJcIlCqhWwyv9U6id0631ijRxM3IhCSco9AjJd8+SPp6ZXCZetFUS
U3uIRWuGvxo7cEUD+gENpYXkoR7ruD3TN6FD

`pragma protect end_protected
