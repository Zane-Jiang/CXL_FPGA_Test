// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
jZ7OQGg6qwtGxz8KG519ENp7P4E1mC69sdxxZp1IIFz+Rz5FswiOat5RfIawRIEK
euZ5jqZy6KdmD2P74h747asuDCr/pIDIDq8u9vXQD4ws0tY5kbvKZxHIieFdkewR
jrnXqkl0hLASFM4iO8o+4ysjk1UCOpEMlfqMdRYgp6XSBjACst+VIg==
//pragma protect end_key_block
//pragma protect digest_block
DioZ8wMaVn7X9dif5qcPiRcWQF0=
//pragma protect end_digest_block
//pragma protect data_block
DaSNU/+35cWj/dV6r5607dt37kBsFPQYGw2jh2Gt5c2h8z6RhgrZfBpBPZNM7CjN
jwbNUS9Fgnzc0iS0YFhUIAmRczNPCG4YgP7zcCYboFMOOixqV/6CqQ5J7Q2rXHNE
TqJTWbYWAqurG76tfvs1vMvgoW8G1yP8Deu8ZnCISI+YAAor/Ws/I2EtCORyvMIL
aA/VxSfTpgR+v0wxT7o21VfaBl0rHzgJ5lk59P9UdveUku++KnjjmDrBc3LEKQwZ
4cLm62SudYMaOGrHSouiOOO8Y2BcgMcQoZ6be4X8xjjpBWW0zrRzxBpLe5Bcy+6n
2KW1Msmmu0IeKtPwK2CpdsTFHyHXnwkomt2MpRIkRUEBAjCD/7U5nFOVCuh4TB4K
msU7L+LH4AioWEahD5LI65NRNoR5pWkJT9J9sg7+W0o4Elo1l008Xg2/camTKGOu
Xs7RWL/S++UQnGBrJJpzEjsYCC0ZdrjihJr0NOd17evEWGBN7wP4fZQWkkWDdHGb
TgLhuiYhxJXrkXzM1YJ025jfBduY/bqnrt+nLc/A3di8Ka6exe6AcUin76JWeg96
yGtWecjNDyHW8QAEkI1zgYaZ/ADKK0naUxvCEb21PCkSczdAHipk5wGdYfE70g7M
4mQ+zB13aFSlNNCU+MrjdsljAgsXJOH8xioevWZsbwpvCpTDfVqieaHTb7pQ7iGB
YiXt0vE51myiCxElc35cSLEt0NhmzA3x6gR7PzlFbKMS/bs/+LFmTWP5DxLbZGk+
u2npC1fDdLUoMZNUfiacCQjEOB7Ez6iD5QM8k/8IQNn0ExalSS6u2hrpuz+rMvaj
WlgJnvCCMWxavryxolDVvTu6LHL5hOqDHow6FKf8AtROtBOyRPymfl8aoZ9uIZCb
DEwmHorb1OfMZT302VqmPYyU66iGcHNhcx9ZZemV8p9gokCAyAXYoIPfnlafg0hJ
c/sAIDsgyFEUOclu1Bmjl1a3eAwvVRaDFsFUj9C+PO8BMyab50h0Mi4v3PkQTwLH
7nFmpSwqHf+7Bu134XTxEcpU484jmjQuIs3YJJzkcbYpSyQjmaveuX94zRtI38h4
oPjzP6R48na13/zy/Npw7CvP6TcDMq+mVi5mEHpLIEdOPaz8THPLECzmfxvEgJpK
1Zu1RMyArDSxIBHBjt6VWpySgr//EDF+20dDTvEu5AcRp//nNBG9Z1UYAnwq4pyS
1vesEdOEHN3mEw38p0czkHQVkZ3ttM4uuYmKdepbrRVntxIlHfsc011KfQnC5MSk
YpdjYoLFoXyXWjdJK1mpAF+GVCm69BwGLL+jD9qWrK+qtQ6BhHrfH+SkiFrDkzjH
qXNX5rhiUvA501kiRH4lMRSWUO0MI4vJh2nZy240zHN8oI4+F9+fvku7QDwUJ/KQ
YFSozgrOWDM64fwQtV2OGYMRTi18QWEFgk8aNlx02YlGLpy18NU/f3awCP1otG1S
pE6iblsZvr2K1iOutTeYFxM72fiHLRmNrgxXhsFmT+Bp3pwvKNBshp2Dig/O56rS
CHsXGJajkMTy8dy9/seT8zL0gdTt/H+D3FI5FHbuqNoDDtsnnEAtrP8NB8pnqnmH
z9+FrUOB1lbezRVavuq7ah2A/k66D7Ipfj5ZzoAWRUTYdfb/9tqbPI+QRifD0nRM
EdEp0pasakX2tVMm5uHbFgx+Z283u8Aw5f8X3e+m3eCMkbYFH9Feaxn6iuAPJKav
1bsUfXJOZI65G/Xs32Z0loqV7va3MtN9/M8A3cBaIIVHhIHg3xqDiodLaiWn/rrU
6Du+micuxW8a1LtdPbyWmOo855Pk4w0bwRygqv3QJ95xGvRQdBMAslfdSen4pMdt
OCxwEeXdUX4VN+qqWfPVx0sXUuF7oREOfWSyRFwbAAGC2XXH3fEeHJf7YB8lmQ3+
p3TqirCVl2cubYlIqoHcYIMl9A+dJXOyE2t303prxaGYdMTQyOzmfo+jJ3mDwtxd
BbP1dVxQc6Ws8QSc4e/wi7PnLpSenqB3dL1RyF7Ztf4VU2XiEcW4hSMS1lR8u161
PSLu3c/hLlgJ85eE1vBO0gu1FKiz+iQvmkRJ/sTR3/u51J5SGn2NmRT3BC+3AiyT
XDCAwli0HcfYrKrdpr648HYtrvnI96js8PfAmWBEyvlEAVUnxj8DIpwdv598w6Ci
h+k7ZWMnWD0eNr/f2V5d9EkIYOaG/Iuy9nOcM/IycBVbn5dzZaKvKspLupSnRWc/
7T4UB/TO2Z0IVBD/cqCZAXl49RdCYSOf4tZrr1b3Uz7151NRxnlAZqFwdE+HlHgx
QQkidtVEylqhP9GBnwyQX2a3NTugmpcNApRn/wWkohGt2OuBOoHZros/9sN8zY5U
s8krlpfxXIWcdrLjLcCbi+ObkI3L1U5bKF0syrE9LXvqiMSPBpqhLGTFMiBWcFnI
mRhEme1zQDFbKn4AiD2OQXH/DLxOTGPCNosQy1CeB/8ryx45BM9KMEiX5PjPl5Un
x+YblUz9iNkBXBnYCms/Uon+cBLyeMS9vkw8Rwqw+uJqAfxZe0lchz6MOIiKKkAs
YnIWXdLXTbMN/flRyVLPapwQNF9u0urkYK5NfxwJkL01cs49mFSVReKJd96YFp+K
ZjSVePKFHd6p4oU/fwcLIpDX5Tdut0Pr/ipQj1xZO/M3OnOeNEyoINHC2/1AxRpu
wDAjpCj7rNxnjxhKezEql/C74xbGAdSCB1GW7H1eAK4KpiWhoL4DnQixCWxG0JTn
Y1udgFhS8UMvQDp0aZ/y6P7LDusdptU/OxZO0AcIE/qptrdHUPrfxtIrUsE6AAkF
mouxkTzdoBdBLpgAxNJ4XDWcT+30i4OxAxp6okWT/vNReFEnKw0TPDMJQPFq+8SO
WO4K7rXWzkR1D9cj+9SRTphtGSyxJq6p91REp7eshvh/xqhq/U9FeORB1r+/X4iW
hEIQuWCUxr6nLklMrIDx7fRbaREgpLLJXHWWoKsiZIap0CQQGCq42lSFSozK++kM
k/u6TsCb2Pvew10ICoJYbzkPisW4gR8p+UOrK4m//ytb1O8deSI+m3UtcwyQF4+k
Jy4QyfKyxDKUyFv5+g9Q8lT4uL/8Jm3velaXmMuJuG3MirOvUJjLcjCBvKowk2BV
1jtuEsEEvFK/LhqGC/N2w//sI/47uN9uT6nEGkDBbarjXN4v7/5mCbnvqCEs+uIg
BI81tmnoEFzCfRuAlpS905whAY+yUVm74SUBBO8/3VNzgSpWnXTc/Af1xUhL458C
bq1yy8y6xEXZ5MsUdu0ZNL+6vsgAOyxi+z8B/qnvHsKHPgAwfFWYew6HlKbdzWtt
ojirrFPIt+B07S2ZfpMcPOzlCL3lDmtXQu/yscX69SZkirNV+KI0WiO6/b0P965b
C43DVl/k7H3T3FSNpRm3kH04ChOQP5YP9pa+zCzLXgVcNy75MbFz1X4WTjpsjKeT
imUvxDROF+mlARSR9JtqfwlioxbCSD23i9jfN/TjWVhDRwtPSOVzk9upWw7tbJR4
Q5LSaGzfvuYSDR27DoFOSUA9faPH59riDXIRnXQP7CCTlbq4lhvCspStSl5mP1Qw
qhZv8rpU5qR3Q8vmkKVQoQBN9IPelUdmJi5E2/ME+0u/fjRn9BQeP25Irzmz04jw
/mE3IJNREdW7wFaLN39Z68IqrpCvewjIJrJuTgwzASWanua0XAuDBPFTAHb3lCH+
pcxM+iC7NQ927u93oMs9EgE/9wRfwdiN41q6PHPIjhhezamAvHSe68Fk4qNdVD0O
JN8ZOdkfs41AUJ2YH+ijLpcrvT9b2gCQWToKW+7ZI9wmN0pZPSPsjDNnfkzTsdnW
YzKvXl9rCpVgHJ/8B4CMxPhl2ey+UZODwNFRoQgSEwfY/8iLl22jrprlp5sbaE0D
cPjkhcPdSAFcB4elxTKt/x98gTEUQIRqRcSmxFv1FD/sG545mamkP5KBONHGtDas
ypXxdIIDPdcdz+7pZdSk1E7YCbCeSAfYk9rSUPTiLWI/9wCoYKOQxHfMSnIRgOIy
tSEdSkF3H/gQrfh/064nrpyiMESW1QvUboHBpauZH3dZBlnmYjO8AqWV8EgH0Ia1
p1h8ny0Yd1Ps9sKiRCRC6z8ZQELHRUg+CFH9gCjkUIfowmd+S50+xMM5RfCLxEml
ALNSt6wVL8pp6GP/bAGoUD/9OEhGk5dRupGU55mxjecR/tpXWrGUS3j0snkBWsN5
RzWH5e7kNtl2T0gEW0F9NsYmasiz6iIg4JvxnloETqdHRc48oWSBSdtTEmjncizC
Kn8MYLmQC4wTd7md/mj4X46+MKJ/CFsxl++mLYy6Zo6efwWN+6+pq2mX6lS7y3oR
9uBzBNZYoFUd3mz9xrH+b39aSUabGcgW+tx/hMawO2sUq8cAzhKUjgwfp4FX5Mdu
AfzionmngVQYh3+pJsJ6K0h7clWXhqEl8SYDVk1wg4In7L1o4L0KtrFCiy6i75KC
Y8uW3swbJx0i6mI7hmWh7jGa3r0SGucYwFbnub2UolhJg58MKFhA+rRSvNiS0zPC
EhNS8CkqobvvCTrUef6qg/rDUrr1/ozLYiuZWZYbtu6grjDq9QeEJERb2l2Gl4os
UBjNbbSW307CWbpBw/X89qNv+cgIJWqPECZdkrNSpA8wXLJ2f3tLyuUPD/biJE9L
bCWG44ewRjrI1LvVstwdxR3pYURQdjiEgTaufquxA/ePOy42vm7f+dlTLhcBDN2L
xarZ+benGA3oMilM46YfPELfgu0shyMsA5UUP0jtlcS6xnbGXsCK6IxzAq88n7ux
Tul5S+hRN9rpd3WRhQcINpv7JS+osIKvDh1RDHkjmRBPq4O4Y5N94kFJv5UhSCfn
ft21/cNOhyAk5FAACPQv4xZHDHiQYL5b4z/Yrm5P2nz/rckjB2O/Si/oMlVofWbN
wGk4r9lvHSml/qQtk8ErTwN61QloQ8ATzjUQJFv4O3468kXkxQuzCA5fs34L9Spw
8Gb/IbWaPqG4/nGrnWM6yh70o3pxr8gbDs95Hb3/+TvCw3ju2VaiJMBlMXw2ww8o
AITEEA0SJ+1yFwFEAWkkQ1GW3LO4gN0WdafjBeDfsvQZqMcOBNFPN5GDk0S+k9cg
aRYptwBitssnhxniVQ9icDUH2NoDBCy1QKgNhN6j94X41vr7TOE61/I+gOzOPyP5
n17TFmdjGhqPnq/Xntzp1aUv3Y+DIG/eQpqhy3Cr4VKZpdtvXwQWMO/lBUyFK4nS
138wQwqpplf1XvD3a18Q32UdWgcyZj96S6m21kEhDW5U/WEFenHG0R5k791U4bhz
S1kZLGjOzOYS01C2jmu6NxK0DtGCPzHutCvWhv+mV6o2DS5P2WMXxWS2rnQkOdXV
5WgpvddPate3KbvefcA2ucS6oSYobbZDXsynXY30wZ19SkWRBZvtb+DenibmcOy9
UGIYmA+9nyijWIzUZuzWOlqqgCRD2oNC5zhoGpAFdFAepwjSFiUFZx4WPxTDLnZf
44h+61za8oUKtDfshJcBt3nAosQHiCuVGWDJrUhBS8Onc1T5PwJ005hmK6HYjS0z
L3qcXaMuy39dbuohboqrr1JKyX2p+fkvJgM3fX90/NSr0FQOXsfAYrbfzrXPNraY
Xa1opqeogaa0AjAXYryBBFiRU2AzDj0N0jD0udvjrXoOrY7T4NVXaM4eFIXfEAm7
u6Gnw9xFx2geC7JJ/KWLMCvquXyqlfiDaOU2l7K8716B1esfZixBU5buTsnyQPpV
aG6lWf7pr80wonCAAa4rzzuLxG3uDECQEf6lB2ktpofyelRok5PZj/YlSviXctsd
QLbrWvgV3oetLZiPnBp/eyzOvc1HMiEz4NgFxy64d7Mxmsq/owsdPg/VxZTa+VuX
WoC2pk0b7NdfTBlNTssOOHdV+/ouDbvo7mzdRY+5lwd39+fsMw7HAIgBP7svdzm0
+zg22znAblPyYZKDbhytWBwKMNyLO14Q1NgiOs7izGNsPdl98o8+XZOBX+R+r/6Y
h41DFcK8L/ZCc73MJn19y7/RZU3H/nxY+WBBbWZGTgpH4WSY1vLIWGdzWEoxckji
cDqWuJltYhHC/sr0ixVJdiDV7JxpTiMI+h30PLHipYYA32Jpmrb5DB1Rzy3vFKar
UDiSQq1HddSVOxsNgH9+QqCcTXQl2O/nXR1ktBdPjac5jFOFvPBLcywZ03GSaVtr
mvAP3NqyMHlweMckttX0C7G0hUMUcx/9T5TdxB6mzhwbm8vXqNFu2ZLc7wwCmkN1
4T8Cm9/i8LiKMq6zMRhDipkPHccy1Vwg99Mj4A/WSEQqOLAzVb7EdsHqgVRO6ezR
84cibcd/420eySaZ2c4hgu8EcVt0M7sptpjEegPCNqAGKPZMPXYtbGEDl7RWgKck
4H85J53f3jyZtVrK9Y4MmBe+OXSRBmYwVVMI807oviIZJqQHZV2SYplMb+ZcfPnt
1hvy9+2vt4fvyJ8r/mA338FvN4aoQ/3EzkteiT9KrwD746pUnKdyY5sM8c80uKT2
63q0pPT1NJzuCPEVWvuO9x1SYTQouz2JgCiMiq2Aj51hMlPKxuDOFIrPrfopBk0C
3UkSaEHivSUc9yXFq21HUDo1Dx4M20Ag9ZuMeGWK14ZoR5XXtjrVUweVe5ESyCRW
KAz1+YugZgBn747+wIeiZOQrPlh7lZ8WZPyYUrOVZ9t6Kqp920OboGHuVzg36Sb+
Ev5cjxulwUlxxlK5KWrqzK7yRR6iAKOCRxR5EObIBt7LV9YoDs6rEq9QDF7VsuxJ
lxIoWA3Vhz9jXTrzXH/+layiNVvIQz2+32+W5UWSfQ/mviGxCyp5MUY+q7Tf5dkN
zRc7mc/Ns6lyAJyodRMzzQEKaaJuemYrKBDvZnfNv1/S4Whj5Lun9//fYUZ2ggJH
S0B5tlfwkIe2zSQNJwJtjn8AUkp0CfJC+c85VoyKIj1wrag5jiClhg9cHIhxrj5k
Gk6JXCSGum4IbIBBZUhBIAjDa5QMlnUe2q0+Ph/fyfmvYJ08S6p2eVNMOEK9PuQh
50SjJ6d97UoZhhtNzhOKJkBeq1M+64SLdjIjTRqvNXeEaQMtub3408oCWrpH0v37
P9gg+4e8DM5MlZ/I92qSMiv8MEnEkx1AGXEPKRnN7croL8XA4jnUkMceYJOAHI1K
ejtScI69uzPh717cpPnreeS6/oLw8q0+jbl6RJra5cN6y1ihkbfn/z7YmE0Ahr/J
OiafUkDwFQklgXTDd5zNSA59UttWs97S2IrKLd6FZ4TCMCEIVKf57sDzk3M2qJ0P
GU6qrSXVpvnBDcS3KKjZNiaGkbKbAZm9NgLT6EiiJijjLy6Zc1eDUaVK0QJzNaAZ
evZ93PBAu8455yyIZ7CISNcVQ165dW2vdz14JJX7LifYAF2EIE/MR9bNfQ27MIFN
ro2q/vleU8pIslxyUFfcITN1Vn6LMWr5ncR34K0A8obmNmiQ0RYQGZcRCT5p6odP
XSA/IrIbRSD8kk1iW939k5nfnl+6g1sqegpQpElyNHGSsRrEtRRuR9xmMQDPVajX
y+X3eap3T34v4P+vGpfOoevIJII9niNtc/BFyk0EAtsVjOVvEddVjJV8eCzfRP2P
WEMhgirg0wSgdsPborZoX9tbmaMKZu/FWOemeufGPj2rg7GRQOWfRTea2QpWXkX/
OVa9q9QGQyGqTaNJhhHyG9woSykuHPIm/RY5PZ8tIm4NAot0JF5KqB66TrD8vO/x
LHDIpE8yO3JCJBmxjE/g+8hXop1oKEVqdHlcWIKGRRaKL34fkNqVY9iHiwuyhI/I
6gV5qn0f8/U4Wx/wyOM5nXC3TD+XXOFZfXppCj0sm2ts9WzIz22dmuRixDIDR3Ra
AlB7xLnSCA17YvqHGBoebKajnQi6PmjFM+ZcA/GrwWTU+tnljiBIsGPlnsi9wbkP
lWe13tDinkfyZaqnGbk/pyDsoCi5yUYN4pCL870oHC6b9oI4+TKHqcspVy9slXr5
SCRWbhBYOQiDIrgk6YJoqFRy8K5k5PBQE7IYgEJcEqJAjjFJriUmAIUA8U7h4E7p
eibWMP/epHWkIO76VmDLmFndzxrB2NyRe4L2Ctm37WCvG4+y+3FeqbDJpd3sBAAM
77yOQRsS/rm3RtwYDsVre6YgRTzvrS6lTDATERqEFrW/C5x4TaYotnlsUzgSDzGi
FdhKkRq126DX6148RyXCBxdw4AhsUgtQZfLN7UXQ1NOiK+vwNxJojlQwIcez/3wI
8zs1dfsd3FXiGsnQDsrG2NxFGJJcZeUqLirDnSREHPRkf3M8KDU8ypt8sbsCZeZ7
t05HFqOi+SzDyK8sobC+qRZEf80cj/3lETwBmse1q8Vcr/MfiXt3kLTUdb1yRT2R
yRF/XTWmrC9L7/R4e3VYdRo7eRoAiEfup/3ln/KHG0ZrKRsgDhcV42hYxy2G+WjY
2cstG3EKoqpDb/W9gaZE66zB0XUUcqbHvMmjmeXZwbjCFaT92uQOItwjwFjcTUVi
LLb0XqtIdE0tEaarnnogdiTDQs5lglqlyCN73zlgXJ1M9jg3wnIiY/Z4T4p2f/c2
rmPzmdTAXKFjgkfdnH1LgeruP1r90Z/EXpMew3iWjTswAJMi35VWv15d3OAnsIdH
Xny3OO0eJ0VA+T0UxoUNVJADVpb2jasPEwwEd2dQnfkFmc6oBQalMO3QbZ0q9AX+
N5Js/yBj1yURQnSOy7tofKZCO2fmfFWOJ9XSpwpg0s+axVveNtTDdiNTf+ccnniN
KLsP1qpoTy1Dttzd3IZBoXLJUq/1uJa4xq1SbFEkkyICkYan45/SDxV/4y19wOXz
VJsLJh8Pf5nf6SnJ6o633wr6N4k7n5LEENVjTZ9DOV7hVDArPZpLCNx3XyLYP9Jr
95YPF5iDYDDinBkdfiogvdAfwNIcozNRsNan+nPSauzA2W4QK6J0MURC8OynFI2N
SXEFAscTMrUQx5bQ7m9UtymgZ+ysXBsjpSljqQ0yW2jmrSbm4bOo0ZDg7sQZfOjp
PS+aNCsE5awkw8L8cozVX2jnDPlpP5SPwbxGzLy1b1h37g8hUjLaMJdfZF+k3RWa
l7PLrMzdDi0yhKBDaO44whyUJj4IIRoi42kF4cOLs7XhRBlMl2vt5y4XD2B0EqTM
9ZTXMI4fNSfZyrFHHBDzHnMUcxN9gCiZf4mqi3odljDZsHP0SbgJxxygjW9nKlA1
JfisMyaPZ03Nwuv4o/37/KyHtC+I/fZJ6NVWvhDqMIJGZJjdfYVmca6MXmjzb0O9
PGYPz3uHsMfYvXNLghhAEqhlGJZgvVS6cxm6m5YpaCRxSwyBLijCdmVYmSoHkx8d
ezK3wF8XW1TGCEdzyHukiRqUsNnbKPxURMRX6sD8E8xG2Wa6ZYJKQNCWN5IC8rDP
tEwK9AYdKEuGHKRMgugDqfwZFJftWxtIPdwYi4GQa8A+Kq8idnu0Wem8hW4dpR3u
wrt3/bnrhGGsCoOMMPZzKW82BM7Z4Y7KTTAzvMxpr3pBtBDBofuEOo7tqUrGUmXq
v9GXxbjK+N1K9sGluubk8ylMxLKDbQHlII+V6PbZuFZoAaaEOrllU3dfEVozi3Tu
k4qjT/LCaZOXgRdPnCQFstndEtVD0km66R1XbA1Kz0SpECrZtMNcxiKMImXAIVFd
qG43JuOxTILlyIeERDf1gEDowTaIgU/RB532jWUqLoIS4CYftGudCv/ntg4jQx0E
cFDbVwxZWK5pjJ+2BNlTB+Vqn087euhlFn1VLs1AKlm5cO2KoAJXhMKOYs6Y4gh6
1YlSZLUwPGOfIHcl/jVZCyZwXbpe1L9G+LWvuycmV6Ani/vhWcZdSNrGV0stwNVS
drB5uTh5hXOH3jIGLVTCXaAJNfvax35L3DM4Lqgqqn4GGwxXAztI7hh3+/miRzS0
CgP6Yk6bviO/9NCXzGMgCM1LMjA/YDzYTziW/U60CYclWdG/6rBkX6OAZ1DbkmTG
jag+QF9f3u3170XPKDXU9pxUZOwGOyxTdp0a1IyzM3PfipTVwE96pBbZnFWTysOT
TwlMj1lTAEX6vCtFpjRnIj9oyzro/XGeJmZwzMyFDd0XXAQZzgXfEoT2zyTVM5Vk
FNsMjRm3TIP8e7FeLzIhfm368vL7xF9x3QkaRCGcgRFhHVTrAgZ98QWw1BlWBPF3
dlP2o5Jx13lgsRc4Gwe5c/xvEF6GHSFmQyob9r1O/Lsz0mlvYf1b7IIup2pcpeQ8
rArpaEdFnv/8QDie3Gcur6pBD9XV0W8WK0B5uajcl4l1J/8orpe2D2qNl/yO/imH
blX04YaHg+i9t9+QaN/Bn46MvD+MrherRlrirtX9yyC+Y823hgZ7ruFHBJk+xWoW
6brkYsf7lNhKnot2C/8U419Hp37dYJXHQ3gyvD946HnbWM8KnLK+0tLawaRB1mMk
8I41fribv2tIqJW+6VZV1MIVDx+SVRpnvsVVdA4uKeraWZPjNLPOORsmSZH9ocsF
1VpP28JGi5lE4o7ioxwozkL9AQn/hXEaZDrT/MMsAJo9MiBioiZOvTQX50MhxUCN
A3Eid9AHEez09HfrwujgTNasxIVnBe76lITAPrsl/JbgIUs/I679UsOSzEN60F6c
CsfMvWUoo8ykVZvJfESaXm5Gt2yJK0wCO1tB2KTwJn7dEpczNKXalFem/ETGGVdu
V7e0z31Vwpvi7A2zQh5DMuQPKBZhy1UAd4364a8NM6fhkHhxfm4CzHfiVWAsDKsz
CUttFcJtSQEcUEo/GeYlItuB49yNcdekKsbTPFFy0cYCxZNbY9dmx9cPhihnlO+v
NZi1FuW9FicEPIC2IOTH1N/pGhaeSrLTlG0gsRkLJmRRf0yuXevCIaXYCiC5pfI9
YPWa8Xg3a9nqFSLyzWsUwDtuVdNYWfoamV80knp3jWTNc3M9RiH5oxAbCGUy8QFH
ekElJcZDo/bVELWGHzd1PraM2GlEaKv2mKJ4mm3Gw3C56VCRXMLab6qSRNccWOpW
YiOKF6LpUa6gtkbcV0Y4K6R4A7TMOrlYnskAxNP/ZD79Z8DqPtepMrB9DsbNvvww
eI/ASp2Y+lYWexXUO5M1f+PQFBLoWkYxLM47BfcY1kF+eb2Hh/kiuyDfSSo47RUU
PlnRLqEc84OYkm2IpzGhvz5NadlwFHtwu3OVr6LMLXdQ28lNaBH2pxbIO7pagqOE
p/ziOHdjHIt8acVCtcg3Z6XGJ8oGxqR3VA4yQNMfXC5KyO3bmVqDGutv8dOAOZhc
1Wss0kOEF7CJzWslwcTke+zF2mPEH14a9lcMAbIyB50PxvKrhYqPLjSKiKULLqA+
GT01QUDc96tRCwOhSmULrZy/xLGBk5+aVuSMtr+v+vQbRhSZl1Y6WC4+1jU8e8G0
fqdLPQ/LtgdE2WoODrNa7ogWBxup7rCC1jiMWXcEqLu40qff2mSoD2Z4r1Zxm/IM
BpDCdSLapaX6TxZVkzdMhJ6TOudEQtZ9wGw2rtLYqCaK7jWI0E5EBukB6P1QDMSW
sQRN3D9A6JPtszSv66/XKlS2288LYG18/k4tHx15kD4sZAKywz6Mi5pq5zzoxEH/
00XAV7MhaokROXRS1PFYzyRSep/tp5yIu3ft16vCGxlt+8pbd5nmCVKN3oxX5ptu
0GKgOcgTEOceTJgC9DJx0UnXT7caNePXSDIPMtK1LDqmRUxgnJPdfGGgbxJQwq5V
aB5FYg4iMrXlVgR3b8L5C34FCQLLnj/tc+DP7Pa0dIw/hZi/G8O3/bmF6Rh2stZk
DOkLIlgfUcRWIj9m4dmjJssWRe9WQdpiUxK6UDpyH+VRxW7Z0i/DS/AGnXJj4CP0
uehsu8AXgNGsbIyNckOi7P91M3lMxBeJfYGtoqW1fCDHOF5g0wKmqBJ+78U8tYRy
F9eqMeh64JVrZ1Kag4ugSuSSVXArdZa8xCUwA2EgGGvnGYfuFxhrInRVZuMAedQJ
YN2KrkI6jFX2NeC8ITuUW50AUuLnqbyjacD/sm0Jbt8RgykpXbaNDXRR70FZFYrq
Qpb6FirhJjFnrJkX7196tr5zudJIxY6IYQKfLC2TjnsO6xJ/KEa1HH9Ug7s97tIH
5u1Sy35eSYqTL/fzuEaiVoq3mO5VXAyVMPZnlcb7tnGlUEQ1wVPeNZR4FdxJSt/w
/U6Iujq1bbqRzLWDfZEpI2dvlLIdQo4gaZnIkORZQCw9xdHEI0rFvW2rFTY8lUwo
FaOPXowxBn3RzsjvP65czCKL8oIlrHwpJsQp7zQTaA1dVTQO0BvzHF1CUw3lNVDA
enTg651Ufcjk2bLCVsE/caM9tISP+qr2/OLKbEDwoZmzETqoGiq5RTDCZX83DeMQ
ilfaLb7Z1yswG8AA28VYT+cjIGl98ISjUmC6CKMi75RlC6Q0fKs+MCqU9ZRRWloO
bJhepz7sDdW+vKyFCzONvX316/2v9b79QyTiCenw21dIW7PZaVig0iCv+G1GdDBb
XJC76sXsfPtNH7GD+C2vBWM0HIXXfXfzeui23dl0RhDhv+mN4RJ1feMUu4yIPj/D
3i/QtMAiEhK7EB7RZfoT8n1cl6i7IHq0gR0m1rKoOVvDrudEetHFIKo72Jj3Ijji
ZR7e0Why8+sbXdYGj3HoCm7/VUPwnqEOTXWW42GvPBXPjQCK7fHA3rRN6clQlc/q
7EudbfO1d7swaOsjnIq2d8IFN/ZgQ2chSpiRFr5M5vvBwXGwtOy/Y9yUPtR61OC7
coXmtpFgHmkP9LtqVdUEFePsjIGdMGhYX2c7HWZXvWkyPsShw3EztHpg6w6nQttz
RPA2eRxUTKhocvttLkrijHj4gi0Tn2LGOKCsY74XPRwsxdllpmKCNBqybIyXZw2P
AWUrLDkcnlAmvcfwfhn9elJlEAaCDh2uVruBFDko4D2zKNc+YTNLY8apGt801ws4
qYLZHGtJ3ThKjHfzWZh18c5xdJ4rBU0vUor8cPVNl/6XNqw8PHtwSy91cItnFu1g
hVr6oaGWR2qv0V2neOnp6tfPlEI9gII75ftc7tn1SuChkjjx5NQkrkj4qTsSERyx
MZTkttx6jRd+QVqw40F6H74UaLy30RAm5uE6YEAB4RaFxM1ilctg2Bngz9Mwce1O
sEK1lNrkQKMbWhz/lbbXc6NK8ki4RSbP3XrssPtZ5Rqnrq5hmnXx1JP+Bg0kHWiH
5yngbdN00ZaMFekuHWFxWxuuTEefMxaqKtaQhnJkDy3spvb/QDRdXjYRYc3k46ED
/jkC14npcxmlrqF3RYjv6oL70Uky75soSBQBEoFsEumkEVQV86LWy+IZyB8wMQnC
rQS3zDOsnSg9M0R8d4r8jE8ncByl1PFETfD9+8KY41wyTOdEKkFkyDMIgiDWpv3a
4fmlkaMn/jhRgyhTUr51Ej8Yv4X8UoEON0i5VjHU5FLkpyClNYAmn0sWsAn82x7j
ZRTHh1pEGoOk5sD2QclGOdPg1gyNzQhMDdh/wUZoLpzEC31kg4XrYw/+X3nuirta
92hc/fd0RZ9nRvalVzggoonUUfZT63aGnF1JzFRnIwxOt8mAFsGzpf/p0pw4pzUg
Ka2Z7IFjwC1STKUd0CPVbub/Nc/Y2S/usdbIQPQx6CyCqObx7yFSKMvm1m+DMniK
qKYDoOsNtsCiTcKpoKIzJoHqUTa1sE6uVKPLHovTazrkFPzv9E2PI9P/Mplz7yFX
2F5iTam2leK7wvc4YlSxQqJW8FMwIhSUGKbf4UOxJ/Xq4eE9nYK1rAsRITLOHX+I
qWV7Oc4phmoL11wgPpNvYN9A3pmuOXyr/0Jf4i+yeNYLmS43FzRL1h2j7mL0A+ck
r3msmvIpw0kBzSAA+VJXgNQ/YcXmQbZeSrfPJjyyFBqmd+Za/BHNkbrbR/o/iMGU
r2PmD1J/pWBVSe3yxj5W+DLp0x1fe6ecbKzP/v8UR7VMcgzSmiBZNtDY5wE408Z6
/zp3/ztcoUJ/llfKHf2ZAfVmPPku4y7Vw4O9bb5WLcemgnkirrE0iY27DgY+20KU
VEelvCR5IRxYW+4UmqEO+L0aMH3k0IwjW4HH2stJZ3KOooo1Rv9LakIR8ZGhMHs2
kLT7MdnFXiNRIF+ETCzR2kK+j35ly7Odone5v11tgcLPA3A5JpsmqxQkd6Q3phk3
PHzoI0uMOUPY+n3wwYYhfagTMXM+QUlaMrXCR+FJNb4pgpqoCKRw9JKj3nkZ4yjJ
eSJjJ0v+6oMTkElgDGqpT4rvTqA6qM1N5x9WMFAtGE7PPLINmOZ1hojEYJ9RTfHn
qkWruhLWXEZ/iZqTmS2mzrgPyMeFCSbaEDE0ezAE9XfK2TeL+u4oYgiKfOmKVH7K
ycvwzE7o0VlZvIcUCFggicQhWNXBlGRfDjhqMHlAtxDs7v4itVwjRWufRQLTo3io
cBgJMvJj9l54OxAxGEyXLXlIlYqhSKhJLzdrcRZxyFqbbccVFL71050vJKZTfKwc
xt5Mu8W6kFmjttKvFQWiWXbCzaj/icI3MQILH3ENQdscrF1zKmzCFrnNjH9EZMQq
hx/AIWviVE9GSKeuhLX3RSC424FqUclytp6tyEqsIwtT1RjQVEHuT3r1XXIsYfhJ
VhoDoRh2SyVoz+dgxDwbd4XqRSZsPUQNygwCUASnY0xFIALegJVgLEzh5I152u/L
y+1HwBUCnw4krRvrkzQoR+oU1eV6Tj2Uyixqw3XxT6vjZJMzZ/MXS5v11fQW6bb9
O68EtjyEogiSaAmVEosHIBqVFDXhYfuSPikaixvHLpk5qax4CsLs/ROXaNPep0Sp
wkimwgk23zrWJdjLwlva9ALFcdidpxUfmcKOuI2k7IZoxx+77FPv9DvjV/A8IUzv
gXS7w/7LWvHhhPcFER9gJ8BrTXSOPk0upWZ60B6FvZw067hN6yi2I/gpD9FSNGnv
pk5CjW4rjrIaumJfUbfejaoxyOTOlpIeNz0n/dLOh5xBOLenaBJGUu9aR56XOlzJ
Ou3s2wDqvNresdnC7EWjwtksAJ/vZPWN3DiHKXrKXDgBZdVP6n/Z4NZx3JMpgOxa
DiLD7V+WL2tGBBhMwk0UvgmdpcSX23HnRuK7mRWW1VxsPp7YH+W1Rn+5meno6JNH
vTb9fPifdTewpGJXhVM5124IriiQDRUzRcRsENBiplK+tVuGnsVwNLOSfZyI7ecl
DBrXs8DIZ/3VXGElYMqPjvkVUan+tBBOQ93LYqdB0OSBcZZ9kWRXAp8E98SMm3o7
vR/N/0nhjL6ZuFUvX/xb/ONUHsVTQ9V9w7v9mK2B6dTy2jRfQcwt3JzvtyHO++Gk
uT9pWSeIU9Oj4Z0cIOjxsjrq+kG2B2iQQ8dl2esURisSqMdiaMY6L+psAmKY6XqH
ppexd1WffK2X/Fu/ePHFzfhvgRuvuqoMNyWRvVCVF+k4CqMlFMwZiRzUX2bHriWV
vkU0CR1zRZ8iH3oqWQOw4wjvIHky0gjbCprrI75AwQmU1qVbep9gcn7D3aFYs21Z
puiWzDjFXrxXqqbG720rDpvzc81VuueM2IEsy+QS0l7p7i7xny9V823j0B3FN9U8
kFZrJuC/60faR05pk8P8K10BJgI0TywfY/WYJtQGH+CSNPM1L9PSrScO6Z+uh+RD
RqwO/QBg+gzIYBbj9FoZw2pNfle2nlt0iqQ/4UZcOs6K+k0NXbjaWkqUxKJUbp4s
+0u3FrNtJ60x50gqMaKHtBDTXfalBVobCI1f2KQzRcj1KeBbZTrHTPBAHLsW5a+N
TAKIWfI8wHgyrtYZcO7CZ0sbgv2jqDRxj4AYqdMyUvo5PtLHTUpZX6FqZvOJMHVo
RCzp0mf6Tdv4X9C6neSjF+2lAswmfSlggg7gYX55bLNCU7qYOmUM4ruLuqU3644B
6CECmWn/3YfYVbNn1dtYkv9qW8hAUhnSW3cgdmfMEZVZMLQYwBUzTgfv4s4nTjs4
vKcXC05SdLH/tVW6z12DCHZCFVH3Xj6b83hYdvDT8BZkrbeMxzSIS/iYW0tZK36j
n/dpP8satp3ETbsbH9Re5mU8JcT/S6o4E8yCAAVnFnVOIWeRJI7l0Z28LUcG+E2V
nW4NwcNhjw44z8+xMghA8+h+TNBw3I4zwvsBPaaGpXUR5IdUCddXNkl0H/286CDz
3ef1Zpp9LHo2llkkO8PsMezS4d1jGnbq68wAG8J+MB7rJ3DauTY5Q8I9OTWlvCxt
4GhG8JnNs5AuLip0Fbmv0QB1rCiowx+YZa239fBdHkuR2QiZFrvTcRoMu5OTopGH
l+f5znqtyXbrTxIgHbEEnw6xokQaP6N6lJe86hzHrS64kG2dVciyah3GMAUOLhND
omRZRi8g+fY75pQbSWE/JoQhqwpC3g3Ry0ZjtLisE6wSG6NLRkY4OEXpwujM2k/X
LlqM65lan8NfG1HyOKMQsQhYckMDCenneFA/RBWcEIfvxjjpXRFE+F66Mb6vkubn
PJIpy98K/AABX51xQdOFM03/lDmnfPzDSCKVbmb54VSsyT45+e/tUGYAFSiHIKqQ
TzjGUU1Z+9n9eXbiZIJnpkcPwdcaUi0UCj7WD0d8C7e3g8mPz67+BxzjLYQZgWLr
O++wC/v34WG+lFZbagRtvB3h487xyRmGisMCMxsV+x714BMGHNoVoJ5YNYdbzM8w
Wb/1uuWhkpJwWPUkRIoKdKOxifI//AjBMCN0zpUKz2A9z1FUSeGMVwWujoKru/fN
BKHKDqavdsxITo/XU0YxK7xpzkk9ua0wN4csA4e6UgS48NTXO2A+C3+bjXOwYQ7y
D2AOkJSgvA4+iQMRrw5sdwW6BMFpC8zhxxiCNoar3WOa0fek2xtQNCaZA755SsNW
9cQKME6qqkmPRxvC9znOW2OnSMmysT/0ygnYE9gl4iD9+TDQfB+ndMZQYFEkrTgQ
N9aKqKCEFhbXNt/r84g/0J9SsDCv0/pnZkQmJ98w3WiC+F83UuueCk3998ZSqjaB
naBHjxJzssDvVtwrnjLcNPGgqyKu6aBrAE2Dby+cKa4gLd35/b7ajuftREopkvbF
y0oKdoD6/oVaX6JFN511OFx5LtcNNnR1iKNW7t4MIIqkO3FDbycHvddMY/SrM/5l
l71mTYNug32zyay87VkpAfH05531nS/vV41mE2GJ9in8RRVPsZchRnMyz3zFr3H1
5rp1lDTI8Voj+8G2dujVgtaZCHDN4tbY3MOHZsanwfWRqdl+Ve8US0qjvplCAZHI
Cl0w4i1SeINQm26oSgyb8mqzr5QQKjDp7GSejG5H2egt1+8qhdBI6ccntQ8F8fKC
LIkODILBPt89NMquWEQVTu0PDCbD3ItGd+BgQ5bfrEjzZNLxq4i8vl2yjScALQSv
kPIyLgcNwABpFOwLzYqOuwrd2YyIQsE86ksgTE+mGKXbPFV0w5tZaroeHjBxQTtm
10eu32IrAj4v9qLtb6uDPcXR9/mFJGMLhA79JVxMdkCoV6yuWdPTuwvCNqsRfLq8
BQ3UDlAoJ0wPQTgtenc+pP8+UgTuQT2TOtyQVH+5I0dn9EIyj2fxuwAMcu0/KHW1
pY/jS7zB7bOjRwe0gN1meSJYMy1mjy7KUHfFnuptpJilpEDlDu9ToQJLaXo1gIhP
MwpyA6JrZfyyD4Cxan9anOft+rp/BAhghFQCb4vmKqyWV2sD4KVwwfHTugzX6aMH
vRh7z0ZZ/oRRtCNMRdFBb+uqyZhHGOIF3sXoagcpzFgxvUKpHNy7eyFTaAf/BFP+
6b6Lr5Kza3eAEoe99s+eu3dajEsMNjH6qHZf1oJNnJokdE3qM7uBS4mzoK3wrivE
raAg2ctWgQ/2WnDLGMzwj0tr1puZ5vXCchzQmV2gL5RJ3/W2yu8GaUfJODYqhTe5
RsASzEqMuo6gSFIJd80EuuZQKLpEfQtdlM8EUYFLv/VG9nI0MqTT5Wy2ozChgaen
86q6uzrVdv3+ML1Wf0NQ7aAF+8mgk2mYy8WWn+UqbQ2FLNGUR6L6qKOelHe5ZOUd
0ajtf4v23WP6Q9XNxiyW/jv+5BcIqQlpcRAq4SCWe/EWDY4d8tZgkDBS5K0z1E7r
1ZBm8aXUEHok0Zq8DTYymbALD+N5M08eDu2Aoh756vlI3pcwxDKERwFexMtNXG0D
GZsNnoESlgau+paHWKnzxugzBs0DN7cjtY+ESL4rCdRKdaAvtDUqbKxTrEdNc3li
ANlU8/iTpPjlQsk9vS29EBAX/sxuMvtq73IXR+UT7o0GLmFacws/0xK4U82YKQhp
qW0HYUtyMUV6HQWVLY45QZ+1CSOmZF8CYtjMycqDYVMHdV/L3lsIEFkaYQHk0Ub3
vJ/QSQg7qvvz+J7ufdSL/vNVZ3GsdnhH4oOCk484qPX/HpFp5/t1LdV/ozroDOqT
beR2+PffkvQhYzSEPvl3jkJOYqbrkMv2W27IAx7KYEZJ2A2vPK9ArpCxIjpKATul
55CY593CRsI+5JRJg21AAsu7bAlnlK5opmW55ZMON+rN6c9PxwddjG07DcoR7BU8
NFqKsAr4t8BBn3pa7q1wWXCdtEE/jIAPnHZJXS2zX4LtoqWD9zTiHCIFhROQ9tJb
DmudEZVUSD6uspN+/Iy2rU5oOPn1Q/Q5wBfg8IpdPFzEH8flp99lXP2UUH0qYEI7
F/lg6cSy889mMYaA9UKqwDnvP1ONizUytDbP5mEcHf5rkMXkYbKr+Fs6FzYXc6T+
enZ5DnEZGkmU6tEgA26ZQjV2Mkq3bcO30r9UUcsSxLLvijez84Vx9H1wu3Vx/k4k
vreOdqLOKi4FHk4GDnNYts2MGSq7dWM+0z4Ws8EBke95qzDwVdfRtAaGUigxC2cG
noqo7nDMPbeJBhKlQkyaG4X8zNrz9QAGcUxWynQv5Z+Q+cPoR6fsVnWSTNRpP0H7
W11uH26DqSMzCav6zE/NPqow1Vn/FmTk5FpRKaH32vqnUmOveKSPSKPl1pFWeUXv
YfC9/F17UMHryctYsWpcBTlQs31PMVE1HoN03fZxOTFytZ7wStifIM0pvsvhVD6X
iOQBzDCm/OPQJ4j+HgUAeT20a2LaDMDqxHm8udvHKOs5AbD8hhm756WIxfpQGNsQ
Aom2QJK8f4MfnlP7ulseeLF68LYs/aV7ZqaGm6xYZBkOnxOIqxJ+SxsW4ixH2VRD
4Z7XdTXkapMUKR20239Bg5XIDiK3PgabkieV5mnVtzzt9BRUd8UnOEpwJAJHra8o
clvA0f++MOlwyWrJvA8zPw/meaQeOp9+I4Pb4VHHBHLon+b04ZHDp5USQGNmcLLx
Nh0hzO8XC0QkivW6VY1Ym3kwE3xf7qDgGIl71EBW1GWnlFGLKBPeu3/LRcvGLzyK
8jG60pevqFg5eqAxnSydAvD0dMgirUbCMw7DgVesT8GKAF3U5tHArGC51J8QzNeb
PDTjL2g2gXq5u2j9nD+UomfGECsIbyLeIt4fePXRFO+aXUVmqQ6Qac//GQiZ0ecF
I7SFjm7oUavaCGy7B9BkBCkKBGOktkmAzqxGIjQbvSkh4sqHXaQLSBwrZqx6IYVG
qWljoqntTw64xIuBho+2uMcxWTjAwtIctAxJ4I+M3l87pBBN/3VPAka6cIxB9i8y
Ct4DvnVVuAlJGTsqMp5/Q/4CfSD8mIE1kHbFgZ8dB3OZdpaZRTbtWBehJ82p72Ft
3vQLQD+a+laa4JN4ipCw9CzNlGbMoYvM3sD1rGIJawcsg3zKaJlswW9pwapa+9d1
RUyWoolHDQQq9cn5/ncKnChYD++illb+lBzSJB3tsi8iSAOMTE0KeWIOZ0ujEl21
YSLswJcjfParfSm1hwQWTcE89mpZ5mxxkIy2Ne5N6957nKCTgBQNbIfxRvB7jr76
c4Bd4rjKxeY7rktAkqgGBFsYmi5IfPxLY5+tsH4baKIiV8w7jvfbtW3TvtMwkSUR
GfRuYdfMWhkDpujY+kVsV0i1mIc+xLEUMO663HA0MIoo/sqlHQt2ATArE7oCUxun
UllzT/4ZAnPFQ4pKWQsdyUiydu9V7uWoM/UUxdKnKLwJb55OxUvsQqHeZamx1pXn
KhNbLav8KAlYIPt7Y+Mh6+ACGTf3SaAhVs4Iu8rOVy9psTzLoHRRNBtis38OXu7O
PCpaslPo8L/saTgAyT4TtSLvSSD3CQ6bEXvafIvoj2yO0wOrrUuD47/ypA+92hvQ
vJImCVNrktt0ZjNEUpNT/tyrKv/ba4kwiPbzdridD+op3PahdsRCHfX2HzEJ/kVn
37h0kIeVe+/4GGi9G2ykW4ewH5u4+XajMfLGRtfi0qEbYSBYxkzeFmMVzE++2eVs
aeRhqyuTH/5G+vr3mDKltZu8LTQcHzzMTnyLsRFyCSoxwYWGIVtCaufUAsSLROdi
wAa0KnZ945smB4YTo4fkW/1Z+jPmh6fLzf1esjnroct57D+SaGBo9ekGyPUmmeYv
7NwSs1YAtBW871IIY+LrUuS/55LNu3+fQUbIus6kH2Aq78RtvxkV69XLDOtOs8AT
t5Bo0pFwVm6XnoLNL983NxVUgyHOyjZ2TJ9DneP9WHhJugJl1L2vKqz9zi/p2W9I
efipscEi618rLt+BaaxHINSb6Dkr7Ml9GtILwuWsGesCS2o+C4lc+X2ERf5eLIqN
+R7yQI1x7/iW+P/3wpXErZzF1OrNAEhsiC95BauZF4XUlAAaoFm3ZCUpMNEsM8MB
m/nAu+gLCimC67vsSIjpRFzyeZT5uCjSCE2lEaPwYv8i1K9Vd1uKayNIBsrpRMij
izke6GstvDvzhCA0JA1D4jYFIBa3HUlCDSrUxRp5u40GR2l02PaKjXwJCAnXIj+x
9irhAsHCCccs4y5baoKQQ5fEC8DV1v8WM4lke5EfoQv5Wz/kPYr5TIFG9jUhqbl3
p+NZ4VQECHEU1ve/yugyvM7EkyOCoqM++lEHnn6Kq+Duofqvr5PETwooVVZYtzDn
OJf44t380QGstAmeWb6NbBL/lRmw1QhIE6oSkDOVwD0bOBEUxSClGZAXzwMp6BDK
HZ1QywL/LW4RoE2mP4uKAAffb6GqpobV1T1TgQNnyR2D0buhMFDm4z7nh30yd0T6
gblTJmSH3gqjnQ/4oys6hLjx9BB8u0xk41ZSeEdU15q7TwgoKLZB7VYNTeNMhmgp
fyKUinOYQs+Ne/KMvT0ow2unR7Mz5xjRg3pkQvSblE0diXQzt0qJ47iqrlpJQ8fa
bCaOFlUqwl/4WkTlTvkjPS83uBDyglQanLY0EXbi5UFKQfXGxerPSWuqcYSDCpjM
vhDkNKTOXtqx4Zc3Cuuz2ig1kE3lBCs71t+IPC9Z8JnH5FRbiriwTpnNItXw7FPg
wkmUwl5PcIDHT7d0bEIHSrGedXhzkmbMnciLSR/MevYfwOnZOaBUqDJ9IvCtdRt1
w1XQc6vT4eCdZcliPR2lbRl/taafr4ZPaKs/cHKUllj3C+PESa/PW/2EHTs1wKRC
Xs5xExPc2yj5rqhUDbdZogsIDXMHqfz4i/jG+BqOg0JF4pg+VsesMkoeeBgwQ2in
8+6Hh3ayId/+7ybV4yI8lJIPUCO7rDEjxwXn9gLDkG0L9I7yKgpluaTn9FqzXpqn
hh9P7X/mq7UebdSzn7UUFBwXyNjK8FlyI0LFSaRbKg71kMI8wWGcztcfc/XvUl3z
dMS8CVkmuEaFenQRHymgM6siA60o6ps//LhaHZsvh/5HLbdtMoe0HhwVdMtiwtiG
n0gkMwHRnptQARLCPDPoohCoLOhTOe3En42zx6AnF8oWKrlvPbPmdIuNDRDGOxap
Ga0l2u4iHppcnckYRJYsLjxazeBtU31/QkOEBm2rEyQ/1d4fye9JbDrjW0E8ozXj
wpEVnx8FL0bjdxgaNEspCSbiSTnZbrU/FyX1rVlEiiavrRBql9pAqR7ajwrTJBdB
nqTY2ajKnQ8acb0ISqcFCJq0Rpy2NY/TJWBOFnLvrU1admi5TmD2J94hCqfogMnX
Y3Vw46sxuxo6to4VhQVx4rrl4ORw1nxvntyJpC3L17SblTsSFx4PzypQz4FFLVt/
vM0wT2sV0ygxSR/+83gtajb/ukYcldgRgZInNjiuY7WSMbRYaki9Bylatc4G4trg
6NuLNuAkBmPsGYaMqS2M9hJJtQAyx2FUehTKM+WHnuwdkLh4DMPhcP8xXHbXfAbK
5S5nNcVgNYz94g5o0MKTcgUku9vdSjIKLcpCRgEPYzOxBF1RpzPvHks+g+1sNWP/
kdUeJ8AB4eyhZYyCdtYTG8dETiyc/yX7jJiMRnI9Cl5n78NuLnTy86zK0AUwSXt5
W37u8TB+ewdNQoO5UZ9ZCw03mt8khsCQVZbKtIk7M1DNzhvxlOlmEfYICF3KEvXS
tacUbmeV3C3f4iFu8yxNCjcd3gLw0Zk6CejjijMGFUQCaQsFyS1jk+FTs9zuy4bY
z/p83RRfDC9pmmsExeltLSHVZgyNIXfYDIccT1CyLV0+mqemu1w62wBEOePPZzPx
SsGEk1YR5Xk+8Bi4g3dX0aKVZeidUOIRqolnyOUjAJosudLLVlFjqhPUWbKd+Sz5
Mi27aKa1edoRgtMwQRtzfqqMbsSagx/AsxvjZtw6Y+B8gexFYNseajpHNQse9KLn
MXpn6MpRkwLmbIYsYF13yEHQXpFb5CD9ykVitoKZKCG2NMRDcEF3OPI0Fko8zsej
IP0/6/w/y1EGsgNQkN0DxaQlFavTPnFIohwk2FwBynE5sh1N4KY0IE0ZKGkkY0FM
aVfqjDRuzaN4W3XIh246c67U9Itwp/kSmB0pQcbr3KSK0c6DP2TE6xgv9Ao5SNDm
PRjvpzXcpa8x0zXkcAwFcSEA6sgnY9yxxQ1waI4jmITNWaN5QJwp2nX1jRThRKK2
k2nypv/G8AsOSomWrOIkr50+B+NA/Kg8KRD6fsIgHDgagaeP5nPjJNDkFgxUoxYI
anch407ZPeOew/NuF330GD9aHXcGjqnzV+OqFof96ehD9ReYLcTFxQf2NIpkdWQw
SpIyvSYA9SXs+pdNLPuwYKyiXT3XC7fjQrzuJx2X8MuT06gy0zjuTh6Gdx7SoDUl
PGsQ9Yter80f0//KRHqzLvTifxs+SBMfY4JuG+I0GscOZ9eLUPUeOxQz0dV8OSMO
Te3a0nTtTslp9s7dZXuRukhrpwFkJbPOxnnElsmAC1EAgCKzOYj7AlmmJpKUpFW2
VvK8+wk4AWCelggn/tUA0FtECQBZH7yrZKAlndL/lPtUDcqz7JVwcUHXo4zSgUBJ
AQbZeuccxUNNB5UVArzDEfwaB66NYYoYEdkHOj0Jucio0vFqU5fp4W8IhpE03WKS
peCnIpU6qTekEldtWxBD7P0ypVDVxM8WsUxWnIAM31ZnvE7JOF/5QvvjY/eNlKN9
+Ijht+9PjhwMh3ak8p0RbmwHV+QpqAeWx4/6kabf6f+VmOZl8bw15SHtnj3HGrnz
ECF3ON3bMFyj5bydeLx1yKEOF5YabpVl2tUVr5JSL/bdxRy6qqJIhZMzj3gvytCi
vPfECyrYAmAI2timyy3bOri9X/Hsi3QLux/4h6e7RR9qdUJfTGDlO5NnUv5IJfY4
d2EMzaScOEXiabnAwDWSjXEyHU8k88N4VHOqZ2xGEbkxzm5RdUXWUmQYX02JkTPn
RjK45Lr8wQMl8t6ii699q5I5Bsg4ud2wLVoOjlRZ0+r5S8XoN4yH76/wFU4dyW2i
a4QOGeF6To1uxYFjshPqgnztAuxcz1CDQgYbyj25nN79Om56DcHXHX82PJ83JKl7
7IQf4hCHiwviATk/TN6nsYb8Weg+bBkkSToVVX+9NWz6iOtRdVWkz1zR1gptsNI+
5S3HvMq51DLz+KpKgptvYjCiz5pVGOAP9ZD+PxRC2jGhi4ki6Diq3RMspVDlHaWO
UozbF8X83aCt5EqGRj1QYlgi4yUmCLneg57jAd4QHQmAFQX5yetcxW3OGLSc62Fh
IHHbAshwbE9c9Tug8jg6C0AKjHJ6UKb4iVjreRrHwAa/45rGMq/9tHr4DJWNIJqo
P4044TUnZ75y4W9BV0jWdz3mMJAAiYIb2W1pcLj/dIckBDqOWEex4pWFEdIli/Um
7nhwsovvGGbPjeeVLnCHXZn1kd0L5zLWZlmfM+IgvLtPIKjR8iRNBSIddYfXao1i
GNfu9PtJm1O9LaMXRj7t2HrUF6JmDpwbH2hP4yP8AI6dDcqjqls7dB95XSdYpf5W
TA8svRGMRfs5hzSmgzm7Ytklxn++r8Ozn3TxjEbsDPkBpwDU0XU1M9vRJrhYiFGO
hp5TBnIazLreKrKJ8B5dyNwT1XuW1UDNAnN4lnM986BRQuzW6TpsMskiZIDsBFm2
WIsqxAHVBOLA7dPfnFu/otOuRkUIki4tAm1r6FtEmIqvH+DJJTBn668GS3Ko2CdY
BKzMxx85Q/A911foJ+SuCrAEQsV6E5+nbfFwB8xZV3uSu548A8gYRkRXqDktq+vH
WTp/iyTBt4j921SIAPxyM86mU6fj3YX8ey7/Rh9jjKC4bppgdF2i4jY9rSTnmdso
Clb6u6PR84JyCOTi+d2pYDRJQbctQPDJIfW1CE2IkqsYtrHpUJP5fma3cFx6rymm
06UwZ1uJjyAoG7D0pVVQOCrMHK1asHIgtxq8Fnl8NzNjwwkGMCnzXOwemb5Y4cT0
xpHlft9nQsAf7mrK+kH35wLd69XHDW5yFPQTByXeHfddpZsXB2QaMBDH9g+Pz/lV
rQcLXULEFrAo5nWPBOE9hHfSj6os7ELZb9FfBDSMzrwrCAj4vbOyHIc/QQ7d4NuX
ZeVqdqAC59IRjqeb5JpGZK8yaJJUby5rZmftrDA+qV/Y5OPzmm/BE3lFu/6NhhOn
vh3Wx+fs2AfemOxSvKSNqBOugjmoMoC7Q/iCi7fKyMvpxckWWd+/pVAHzudKlZBq
LaNi4TtgSGawq80WFcuHCo07FT7DBOefUFuhjCpAa7FoFXu0SdAeERosEDKqa6Zi
D9bx4xHCKa6HBGQM/fTzknccsv1D4P8zTBjk36T0aLVAizX4sw+QKD97JNfqiGcA
Zh0YyzmEcZhmJhhH14ZajFVSL4c2nUqGrqAnIH2VQZq30BYDHnmQmR6w7O2N+XGK
OSXElzDd5xHCh1PN8pfgB+IJEAG+vTjwRa7mPET8rGdT1Nm/MtuhsH/vNaeu+iLe
cKtNi9tvrt3H6D5c2oiiy6m4oEll/WEEU07lMty/awUMSiNmTRrxMrfsjPCO4cBn
rc6CXEML6S3fbwUkgZ0P2k7nPC/OFSmjeXUfa+jtkJ5EQMHZb3FVUtQP+7GMIQYy
Wa/O4BvhAAB1cYwqVT18ojVYXfq8BaYsu0fgM8Gz2VaD2lmarym6EYHxsATpMGWR
DbMwO2bl2l0HRPb2KXPtJPQTnsIe/2VdNpXt1vj2InnxLwdDwUoflNua0OngMPi3
1PDPmRd+zPeMZhZdGkj8poX3qmz0U7wxWPB/1SnXzMzrvSLyIMSMJvdTKDCxgS+t
UVc99U95AIdh1M8stFIaUgPZaofheV0TFX8lPjmxOiooTNQn+2YpWoMnNeDhTZ/d
EG6TtaTM0k8bFwe1mfXvW1/AOi0N7NT0DFj3pEZhE8/DR+miNeiTJMKXBMKw4xTJ
bXJRmCKH4FxUxwI2ZJpYHcGbc+dl6yMvLqd/G4Dhfbazp5HporEPpMrvPlawWJSg
D+2LHtZJ+kg0fgoZaYMM4/tqIuEZ8L5mZ8PUQFIOEQ1MX5h1CjiJTr46oBZqnxgY
433enVHtuooDqg0WPGkSHe2hF3RTqElhszZ/xRsj/1c6F7ddLuDxhXYE9YG6GcOT
B+wpecTohi8KnmtIKk1gZ1ITHIAoCUWNdkyb7Q2aQLPfH80gSAa7zV77S06SSbIJ
nZvuPm8Twva4gtVcSonYGX5kz7nQ9pBrZ2q9kuiwbiTtMqzenlkegCYgJU1FXi9C
RNUVjawlPO2ag5zGpbxxKR9eepW9XvM7q8jBcPDJ6Kd9YmsbTveQ5Be70vx8Jym1
5EgKrFiNanzR1aiPbV4mHbV68AUCNqMizNoFE8MMkYN7k3LRGJMuJ71lUL/4cgDO
9S2Q0QoRwKNNj/bZr7PmXhGvrOcM7Q3wWshpJ2cWwnNJa9W6ch4aAhKbNs1R7tj9
3l6+l1hM8+nD6c3wxuZd26dqgcYMDxpILqPF5NYRB/q3MpIfFs2bIwojT9I0CQ/m
fwkkkzSOaFo/JZnKJNy1DpQvpdlkr0O1OVF+yWbIgwbWPK1tbyK/v1NosNgKI/XV
QhMsbjB9exA3jM70I/u19enQiEHeLW8QNy/o0jDKSG1nc75zegDfMY+hqNx/AG0a
NgmGksi4FJCKRluXIg6PCKh9UTfXGgeqPrqNoZdIK1IOUVm/bbZpZ/B9KWT+9Ke0
ajBie3QDFg+YH+NqsskHHo8/k3Zb0ZA9nGTGRj5ufaviNkAeVtOVQlkT7SDSkQlS
AcUDpH8i0kx+TDUFNtzc4P/T+/m0KQ1BOyWPf4j237a4l2/FhxWa5VyEIy+671Wf
m+l4Klli2VK085VQGdRZIsxXjgFdotsBTsquOuFwrR4RK9+CjMa/N5Q/bjsjF/4w
7/2cRcW1qM77Pv1SXYF9FozUQA/A6ZV7scv376VqbqReZHcJocNEFPHXuxMchWR6
5v5I3XvWHxoF3V4BwrbT8PbRbVHS9npoHlopFrnUoa4FWBUm+4nyzSfFjuMaADf1
nFOajzOlEjeufsMHYqK/73KGKE+hfcD+tJMzfoU72QusdB7OR3RRd6khfgn/VkTX
IKBIVDpPtVobaMMpLiTkFAi0IjAksBSj4x2kb1b0DmIiZ4AqPjYcHpG1I4VOaVRb
VnKCVGdnTwWrYOHsbpOphzLwbDTPD3N2gl7NtsVR/ulinD+VpIw0PW9gGFWG+EaF
cas8dchOTKK6DfmStuItzslM08EWNNUIpkZhVEUB6eXx+EgQ+lGydJbJsZJl5zou
PdAiJTxj4+F6Nd9Y3I3046nJh0182RUxLo7aQL/AKu7868IhB62SNrw69J8qY1Rj
XcXCZTanYTOXp8L0tt1yqRkuTsw7elPsJvhCzwqwCpZRj5yzsj9GZpvkmVHn3zbu
vczKg1kC7y01KZcrGHbbC4XFWbYD0QIvjItzT+fQmqBiteMyXxmbS8Zt0QGRPJKB
WTcBlGo17LiZQZAsygt8D8+aF7EEYbXvFCug4qLSTMopzoh30I2L6SzfYmW617zV
kmZM1jmFtbytQk0F0tag51OxhSBiM5Wo8Y9audDEBbaFe+LnEEAa8O6TnpILHh0J
g72ITSx8WYzcvNClskkBDh5ftMKI9mmG6Mjn0pfLqGzzqGKhm46huFBGEyDnNn0h
RuZWchidT/4t5b6MPUSLlFP03mrOeiMhZDUl9kJHHdu7Z9I33hhg/tMe0D79mg8u
ZutcSVx/vpFayFHzI74JF0d80cOj1Twk11yF0TR6NguETsyTJBs5xQEpfFoAPFev
tctdYdiTBC/GOTwFYAKP96C+/qp00Ysv+5kcgVUbhZ6EVVx8uagwyijgxHG7wDSs
3/9o4hS4LSPNQock9/BchiZbehk0Js8NUzArYwfM5Od2cC6oc2fEayyaRUBI7B52
xJxe3QSP8NzrbUIAs0oIYU2fWu8Q9EwFBj1R7LGj3H0VEJTrXgj+J6BCxdCewXl1
qz7b+vjVXvydlg1eltWA2tcVF01aMsd3oGEq8CEyMCoa3uBSm3nPZ4g51ZraaX66
AQcirxiuzIe/btgkSg/DHeAvyCht/okANvmJCeQAmjJuCURIYI0nUdKt/hxg3COA
mQMMURRlY+7P/mgIfeHWnfn0qS//fEUHZ5182by0lQ4zJXkC4RBVgAYIgMJBRRCY
s8rr9qmq4hl9eGF9fdJnH7Ii89Sc4HMzqsJ/jOnO9/lVEVnwy7IRDxHMEscqSZPG
mEntxxNkpNRtjKh8rcho97Otxl8iSWXP608n6EXaOw7JbJi6uB8DSa3t2T4+ZzFn
J8XT6VP12Gnfd578e+ya0sbFJH8gtcMy9+cYoCQbK7Hgww5JbnLcHC9VkeRSXfU5
PkAc7TtLXoCIK2ULkiekXGRpuXQO7r/C40+T29Ia6mPnY0gV5bM00q6topchLekO
KOAe47YQPUVR+4SLrlqIzChCQLTjDEhdcctgj3dBDiq7zs/Cqm6Yfg4u/ZyMOIsg
WNRKP1oN2msr3aqG0R2X4DeP0SIhl1FIvPmv3K5CmgvrQhusPdIbabTMT5xQkVmi
m8vgDqRE3EtywOPXCi1mFyDnspzT1HYut2D0748WxNWxtPM5sJzKT8h+WbXJ5RHV
kZSu340LUPeb//Xy5neV4Jsi8KrAWbtF0TUIyVLxeMKQ1gw5xJJqPM5O7WqRNiMc
vxhbIdCKeTWF1F8GaXS1MVh2EuUX+2IFDYIhvumiARFH/AwGhca5CynA5TmcJNys
j0MbDY0zf/ZoZRkEmhtis/sgDQ0WKMoDtxJmcoioF0e/ic89bKLOBg+7VSF0WXcn
tWWSd0/9feUpiaAjO56D+clgFC9k3DuebK6MDaAZSoMSpVEpZ8ZF9SxA11qIZucc
W0L7kX2HOEkZfIw4jjgA9X75G9F8CF4FcEmyc7wYcrmQFdkVzUi3rAXSbxdUt36E
qkA9OK5M977r+dz9MyCXJt4VkrOolAr9/68t6KJLIV6be1SVqLneWSsdx3YONJO/
f4LbIQmfNhk/QrGT3Q0w1+YT3EFOVbltdzsVybixYrpY4saCvIneLDwNG1vIOcP3
0ctssoqns+c8UklcJn+26+sL9Y0Tiitc70pgyTSDDIrmWivDbhb+i6Y476idert7
5Sk9ShQ7smkxFkyp5MeWKn194VWEGoCpNZDiwggiFdAKbE/0OKqc51n/G4KMId+v
2hdA155ugYzjGdOUkf6V5rQ0ELP4hqy5VtgxV+vMqT2y2k//HpCHhgltrILOKFSh
nClBU4e9NAjMMHbzYDMqcESeYNXMzCLKFk+pFNy4XB4XIGG2jxHlzMnolMgAUBTX
dgEp91iYm8+xqy+QGEp1pJqvRsDE6tD8Ev3RmPkVw8+/HfeLLAfahmlHc0n49FRo
xUyk6omOKi5YYGmnlhaIEqRzH49JcvEW7foGnFyMsysHLVd42ZsERxh++6nV6hXE
dtLHeVBmyH3WDpg/gopEY9sWz4UoJQE9KPYM8JViin7X3Vbw6L8b6Q0htjAeWInw
zHrpJe1UY83nP01A1Cp9U/DZRTCT7ytKA4FN2uQUOa+ogAUZBkDXMeMG5s0XOZsH
HSZeMgKIrSZs6pGmIeH8uZau4ORW4WVjecKOp6tPg780vnMPCPTUJCoJeShSpJQH
pwS80bNexy1ZLHZwGCWvT34VSlRdpHLvLL7s/5sQr4Bpwi5mSUb1V1sGGZJYVP9h
ki0A+UPY/e/svhV/cZt1+mPxkWZJbKsqsSDfdsf6EAKCmeATtBLTkdUHKi5Yi5iD
wNatE7JoQtRQecrda58SMV1T0M9OPZ08VzTBhgtEBGuskcPm+cOjKx/7iC3VCe07
lUO5QBJOP4io9RxYCh4MNZwfhxvzBQcmQ7Ht9MNkMeeDaCVaG+y9XH4eZwsGjayh
JUBUOcb50gSVwMatzR31GeX5h4nbJN3KDR0EDx2rg8gtIGeGa27TEm3fafPpgujc
79n3GDbujPyEx8IYDtbFnoruyAWuEtcF9a6K2z6uySA4Aa4dhWKnjQjTMDgM5tlh
wOAb6lwUm2eoUpwPFzZ0YOaDlM4urUtuK9OTMJQkECUx3zr7xUF1HjKx6iL1vqd3
XN0+/XPEDebAJ5wjDKxXEKLfRqSVgR5q+Fj2E4qrpHKhAVmUZ262Jb8EoN2PyVgC
+dLfzm8x6RCmLqCYhjBTkIV8oIjwAGrjled3Hga1T/xQetSptVIeDzqcop/UoQi1
QnIFWq3WQ8fATOTv79K4naFaTWIbvkdGe8DfcrbEInzwhDzGW7Xx9NEyi6Ffu7eQ
wkHXL1LWssN3covVAOr1nDvlLlT450ZXbfrxWl0jnv/dzmSNILJrQpwejX4VT7MP
RFhsVlPrf/S8vbxl4a4XMSzn3s/xPPMDzmmJZJnMvvVBDYNbG/k8zki40Gub/kp0
LD3VcyWgllVNdp1ARCSE6lEPHOe+u3yhBQdXgaHCWxTgGm0vsJ7P4e6t3qLY7YoL
NMJXOBifP2/stjgF7596mLTxSHotSgBlzzeyeDjViDt6h/siwVQG3bD7xp4xfDdg
CdSE5PGFcfYDCb/AobrfKlveyUnWVPTJvTGeVrXMHZ5qlHqmNZkmmUpRJvzBDoXz
arRaDfjT+z3dLyvWJOVIhq37NxlpJW3jlsE/sgJzkgrSCI7LP1PFdEKH9bAzNCEb
sr5AlacxGhrTuO1BGRxBJz4K6pPFIh/RAjM7ivZG9HmdNbvA8aw3Pb7uhAfcBxuJ
nig1dFynawUo6wtlnwKVYNFkMjKSOwKGEn71Cgu6SdP/dn0r+QsTGqe4c7mvMRfd
GZDKNTXEAyVZGfE42BnwNb260hcXm+jRwIjp5kLWrGuSUSr+N06+kblRID0rxvdR
IFkV6eePV2FenJzAaiWi5EbJroWJCNvv5+Ir4bcz3t4PRD4/UN9n/TIFiMr9StLa
mP9NMqpoa86TqV2yqcuMz+veHA/JBlrBlFluQSzZwUMT8/Y7NzheDxxdA4Ib4v1x
PG4/ll/IpJpP28du/O/AxzBbN9e6bskNxBMpHqaD5NNpJGbW+5tbiOth9rt5HpSv
cf0ky19rjrFER5dW0QCNs0qjC7YVERwpc/HuB6Zlm4S1FhEdbbqT/uUTwHCIp8AV
XKhsFfa4OYz6Ucz77NGEeAV8w/WzV5scyyd/LtY+ZiUyX7ZDPHQlOafGwK96pMYl
Pb0NZj9zWG/KnbtQ4dYw/Sr85rR569E5BEeYKwJMX7vN/zVDOJnuCyrCeZsRZLP7
l9nBIZ4vI2IfVs2F6CucmspgJIXnObNRK7KAKYWf9vD+xF0zRv3S8/xTBsAZXPZG
faHOF1iGMDYXr4FBTQHU+ebL/whnFVkpA8fwtpbPn2v2IJxt1iXbsjeL7mv+ldwC
Sw4O1+k5eU3kl2wmqji6YucstpbHcV6BVOxK+aGEiGbQfvizM+vHfOhpyoOlMMmW
53RPAQ8wkkTZk3D7Hfe9lAICvM+kDZ2amfHI8LtwnqH64wsXMN8QTqSfY00feEYY
qIWZW7y5/5yTdWDFNAMaVMJE7nZjwpVXtk8QCr3cNSZRRaeN0CILOtZPCFFreJ93
n6lmbIZX7Ps3ERkpSVsyxI//1TATny3evDkZ4hGA8/k7vmIHTFJJZroW9Ab7n6gf
adLMZ9Lty8nokDpy/ujdEnwOgGfkXdsuTWeLbAJEoAaGgUsysYpjz7a0Su28fRI9
8GhfR+9Vcrd2/PzrnsHAZNT/AFAp9wU3azKVkbge726+77EsQ+KW+7u+LlqTg59t
9T4Ora3mtlmoQyC42lpR0q1siRJs3uC8hE31Uyc8HCr92Hh3Kck0eXjuybRzDJ+5
Q/AsO9X817va6+bYxZ0U93YJ1/S/ktbe/tATIHFvp4KSsmH1z05s3EAb8ba4HKXd
QH3GQVc+O6AXU9INP2RPbPmpdt5x8UW9hvPgkF/IaVYeDI5GQqvTAsfYy4MmLYFE
JVUgZVNhSIwDyiDSBu+cwZuxXfmZzOyYgfCJdHfyAzqo2S7p0H2xbPDSLYtR24Lk
nUrUvG/7DdqM2lIw3RvEPeIT6rsbBfCAFbi2jiykz6UGJ5JUriiyzSG6YiW+x2u9
VYVIzDm7Qb/UG+F4HnnGy6zIMKRXhK+1nnkxKYqHjdv/r1HiaQbauiNSzHwcUkLh
SiDS+5VwJuspk/AEGOWa9aDjSUvKigADjkIWeNNaa0sqoOFpi7FXromrgZjhmHX8
R8WJDvYpuXcIMzNCxLXGLxk8I1wpqA8JpnLnahTEgV8fY3Bfn7ynTqiPvWqSEfKq
h3iOcRO3L+qsmvipgx5Pb2KYtqJ1dulxj2Mbcy9Hh5z0Qt2eEtq2hQ1plrvn/71t
5qX1rad5xkULFsDvN45Oah5Np4czUcLft8qakUnq0qkA0cm0NOoZ6ASRD3B478rD
GDeW6oGMnlkyIozOpPraHp/uNCbOsk/U4WK940lTYMBB68GTc2YYdDhnifOhjn8D
1+rOTno5G3xpNJcPlQRZsBNYG63d2WQTsi9HQUnRUHwc1jId7+9py2VvQidtBbT9
AMzWtqYnbo8I3QkQRKm4T8bCn4gsUoY7Ob3ZHJU98yhiCT/zOGHzSa5OrbXeXI/F
g2x9Mdy4SVFgfY+GEGncFKRwyNKWb4I3JpNWdD7T4abzxU9bm9Dj77Ey6GUuBjj+
Lb9kRXFduThIXwE2wONPD8ZoJe72ZoSIsQn/rZ/DVJen44RPO2PwigfbdyWVacDV
ATqYDQjg/t4vzrGCUs8cinJ1TPrtkiDhXVkwlaT02I29OeCz2d/Rfyt0ogvY1g0b
/6awQW7oVh9s7kavb2o+Rz7V7X5pkcs2ssf5O8+1UlolMJU2r80c4cbw5vmZ2TwB
eKEH/DdiDJDG8ykctEzsrddh8m6fQ74mDgVL7NDAiJzFzpYVoplpAqKmlR4PqG/X
MgSnk4D2pFLk7Njqoq0G3FLQI6xVpBQ4Bb1T/xS1lgtvgPp5kCiwOUnQVD6flDXz
PpGzFJM3dXMtVQ3c/otnBy02gViQCDpInwg5ycRJmR+4OWGyZPY0RsoiPDOYf1st
fH+BhDeNNQIuxIrDOG1FCWaE9YGgcVtSXmU82kfVro2R5lTZNb48UCB5JrKhlK2F
21EJmU41/BilxUT5+UEgoAEYJD8eg+80mysLeyxoiIE3MCxyoHLw+Uyz8L33OQz1
CgRR0Z99sCEh+MCQH+pDUBiqmS/bqnY1fZ8BzLgnKwI0SQ5pjhnzQsCodHd+VCrp
M4L4I8EXCv9dYdTMd6sRffxbPk7RJxrh+7q8cgWfkhVVj3+1dG4pFGIH6teM5AR+
4rfX3ct7XgqyUjxZUqfcGPLkx1v2OrTUutZY440kf9wiSCn+zX5AQ91K/6N+Vn6D
mX5t5fP2i90AbfcFWmuqUT9WIPGji1jXSzQxWmeYIJ5ly95z5qEYRG5AiRgnuYe5
ITULGAhQn8OCKBCvwOaf9FctlTKPnIBect/IvKlx/nf5ansmW7+ss4Vhqt9jE5vO
18tLQxiqK1btUIwlryvbWoiTikR1pVIC80WsTeAWtm1zsZ3cYSswpLjSSlHpu4Om
CR9SAP+guR7nnLc/O/jXjc89ku6SHpYduEFD35rAHQFl6yXO6kqkpjWN4lSgFZbf
a2uqQUeAu4+8m5ot/rJeDk2a7znz+CAtq5xKoMmUtu/t410BZC41VuPLaQKI41Ts
2xzYVUpCk19FvThAmvAQD03ghjmEhM5Gye4ejR1qrTL1g5cxfIZwILTv10pFxsgh
H1g72SzkihY6lWy5hnYDRKbNKkHBvOuJNvCJQD2v49/PDd+rA3UX0mqmnNUx/Kri
OUhYxdPlOHHDi+geuJYzkOv7mMtsITVYOsl/0u5zgc0yKmoQ0uLZAMWpWHrgisb9
ooqSR7EAGDjCbBed1BbxoIy4QlY3mXW8SMGnO3bMEAP8abt9aAC+bWmWbvSRyBkE
M2m0NMirDlMzgaiO+IRRXJDwPfiiEZV846Wm446T3qlAEXS7uBkDkcelaWaRIc5K
DCcSTFRat2N4TZFFKws7YYG3j3OW5tm0Mi0MwQh6+RHz8aQyH/3UZkdBOHi7z/zP
ie6K7yqHv9omK/SeS9UJo4TPlsswCmT8KbIzByjirZXgLyewB4XGYRKzrI2NZ/ZK
FQHW0YQWHDH8N0NPIMici6wEclbzM0AGzOF+RVBSiaQU1psehSJmjiYl0ky4GFSn
BokTDcmOuHFotUtFMUkZgIcMIHCTren/ViNdDBcWKQZEb7BU5B5BRegD1KMFx83T
jRZO5YCF+b/ydCi0oVY0xe+lpbrp6dDV6QQQNBR8l6rm9CYi0ETDpY+SFXSHbrUX
0F+YVTgoHq0vo6msBgxOaTTyK6xPczx6yFZDbglhMji46nICR4tCEc7Rtz6OmcFY
GPPIKdkTsnCyGwuTvGuJ8/QN8rTiJK1z1y0jN83ZV8FlGX83SlIW5X41QeYt8uu4
jdOmJzN5t2hWA/SmtPQdqruxV74150BbBfl/x3X3o5DVXigWbsviI8O00fC/laAi
jVSoOK8DtmL+zDUijnM+Wd6D6KinPiA+WYux2H3lL+wzS/4j7pIOZ21SmOgsOU23
WGQpmvWlzwNgwMlCzDLrnryuCX/1/wuCT9bUi0ESsuGVbqAbjdRw5sGaGCr5Hzp5
/mjkjORmmP7ivwUCiurzblW5raHNtejWwZw44zM4XyIjQ28NM/qHfz2DbZEI5K4P
iLndynZ0EIYMzR4/OX/6o40UAvT0ae4nruYTcLcf0u5kJ7iIQaMcQpA72XNG7aUv
mTgXwjLa/nxP4AX6lDL7UQIoIOUNDb5URmFxJA32cJqrBZMHpXemHoKWztj2JAWT
Lk2B8FdNVkXb/xJTdARH0AbWNrJmcT0E5KYZsrOSiFXftjgcbWQWPWBYnPV4fETZ
mALUb3uHNgoORvJWhumeY5vwjhSuMHOi1GRvtlv9wHRWprN1nQEH6JsN258zfYvb
1wGDRgfMSEcBayqOBcwT2q8zo/nGz4G9kpC2mb6K67xh8pcQN+Dxd6caaxK6yENk
uh70Wni8Aejluaax0QIErmMVFXQYD/3iheMHXNFmE1r37B98ZqxxTz0dNvzwgeiU
yTOQBpU+lO93kGgtO9Qq3LiP9m79pKH5EcU4sBhH+3VSFhNkKH1gGxVI1yfdCEgc
5YRanMlLnxN53/GV6MyICGEUAthRDFXFCqJZzY4EYCdS4afna1AGggQTpSz35LaT
m/n3x8njTKv35yTqip0SGdkx56gvDMkIY9W3H+/uuJIGLPVRsd53EA8XKTABbauN
6KccK1wE0epQfTfY/X4jZ64sA1yMqC2+wV7vwUh7RuuEpl6AFxfyerp2ckObp9tP
SzV0haY8fan1gjktzg6s6mzKUUjS6ML1sHWWOOlgIiP/84Kij50m8tE82yXo7JMo
B5rJxza/6EfvKdRwcCNYxjhfBnwUVmG3QYHIXHEQCYcb0LWJp+tZ4WzrGeZWHHJR
cC1AyfRVEio+Ngv0OKsT0IVNFldVXkd3g0A6i5BHpe/20Ltce5nonMDR5/T5YRuL
Vz39kEfU4pyEWVisXqkFIYYALwZuFYhFs9h3AoZHBlKmeBqmQRf4PhdFdP33JFAd
X+xALJW8+xo1jjzptSDm8ByypxDY6ReoQobRgLxQV9mzURaEAlWhz1QwzFIsDDRU
zrM8ciEH0jiNzg9UgdVOvmA2l6LAe1s4L5cVevXz7NWt0lHG/rliu61IM0sX0Cat
jX3BN9yrBDuOaSem+I7KHJ4Yhu2gNpg++LE60HCMLMYWGrWfn0gz8iJj0rEpdWmT
5s/9VRHpVzbqmfC9rcqKEl0PGZblwPAo44ZVybyMpKbSmP5MfTJ7FqzqDMLxgLUN
kKai+u9Vk2AQNH0XMd94dY5Xi6V56cEFU2qbp5pOTGJd1Gg3QnwB0oiNmV8zvmqH
H+7b+6x02aAMSxlncosetz+ybl6wUIbR8wiKhYgvJNiZPq4OdN0x5JFuhf7aywqS
7U5Th0XDGTMWTbbfr1LUov6nxjvH6Lxp5PCnKFBi1sOKED1ZaEGTuZ6a6tdyEkyB
ojGHKA0RLQ9gh0kuTRnGHok7yAkBMJIbe7iOHGhddw/Zy3Jr9C5F/qZ9F5dL6J37
qe2Qo3BXRMcf7QaZYWYO6ibZ9gPsK77JbrNoTfPfQ4VwSPuedk5qvcn6WMe6mx38
IATvIQs46W3OD8G8IQWfejUZEfoNDj82DBJ6HJmPLTPHjBn79sLTCCcxafWAZ7tN
NwhvxxGwJcwsv23TFmaOvzaZbf/yaAmVePs65oX98jIV4lHZ3GrYAUY9D4Fc6KTA
zjOvoZ23WKGx3HdEtQjswUc3HBuX7reVFoHgqgnanj7vf6jmjyAIeHpU3D9kHbxR
4AbH8PUL6zGo/3Nnhu1v85ED6q5Or6CZeHJV0mJeVec/snboTwu4PRnoxoTqLhSp
y/5k6YGZ7Md12+EhSC4AGllASfPUomgPPVDAZY/IAkZHrDsD6Ui/4nIPkGbkPjHA
m/akUNEmvELVdDZi+5k9+uSbrFK6B/2yIKTlyjMGsw6bobm3y+sID+TW8629al24
wDgFDmha3YoPyyPXn04iQXLb04ZxZ8E7ClMsjxLRx2RahCLzIAsR9JelNGE+LWQB
6Mb2K4LvRTEghXGzuj4RiEhEIkLrxH9Xj/mIQpmuBbD0F8VElwlKMemGMmNiV4Yu
n/Yv3/DEf9PFCZAISw7MpVM+hnJ5aqjV7tUrdVjCYac7Hh0EzppmpmCo5pIGINXI
/psjyyDs5tBWCLoyVzYoVAA4NVlpOHkmpxOgYpRoB7/7z4qwrw8Z96o8u3viLJg0
keUXFPuhJD2xGuw2j2eedYPRVRL48K7yF8LC5En0GgDXw8M7m/e+POI543rDFvLE
l1BS7xVXGfsWjufiPsLdXkArCKm666qO7tNnESvr5qCVhFzB7QUnm7IQucakLGOU
ObvGZqGp6iRs/bDClID+VM/KmqloZe+Nfz+wS4DwmjHg7XGiGm0x/mulkHcxAsFI
Q/TxySVMM37JVfqAvCPpb/X3TJMzCbp+ZZqqPWjbArKUJ9hX6R4NrS/EapzHPpjv
tUfP7qE740EVMQUeSs7zq8e2HALlNyKo3n1t42CgTp81q2uBdwiUQIM8o4NySNaW
JU7WGqX2cmelqm3vGbxHo1xhl5R8l0z2siuWDmQWnD9ODR/cIUBi/zeG/MeFoCoE
GCyrjl3MKWpB3I+GzrVfMbujbBQd5rI7TNzxVHLsk7oO5spgvZfZa1r98rwc2dWV
SmWK0hsRK55ToeUphCu56yuvUTeIFs8gLHFTXmmypuVFKgbPVZlv9KMvbHR/2ah6
1teus+9HQxxpMxuXPtvwji/TqQYzcbCuJy3ZZHeaWdy/Szc0WvZc5WtkXsEcuOtf
ee3D/V5p9wUlpB5fhA+zik4tyQqK1klNd7sLbw01TonRjm3pbUwa/Vk0vpJlNvRD
gc7kYa2W1zXFgs3BbGrhqt0307EOc9RWEaLk0bwt1Qe4dm9QQgkS1hATej2a3KYg
VpR8QOAgNfQVrpSqa6p/IZuqMV7Y8d4FM6k6QC5OJqKMvz6bvTvCHNo1A9wWM/jA
bUfI2B6S64cQH4e5DWmcN5+B4v/a+dzMSp1eXGYPiF/T1WP4sVsMqo1ZVqUvDqwm
2MZmnAiKnY8dhxW1DTGjRBZDpl5NB4XIolfE3LIqioYKpsOG1F1xhq6gXCA+ASDP
cRvfvf7oezS6UGuonEwIFbeyUSaQYUCle4wvk0uwU42HIbNSlDs3HRI+M5b92CNm
ME6aez+8WVgP7oUx/4ltKGTVOHQkWuaZTAVdFABOfk1nFYB3felxjaPtxX10O3/B
DfGVPZvcj6slUZN8tvtSAMNaQYsPD3l1HFugAIuUVFcHFKF8QeOKREohEgGP68M1
lrjKKOsDmhPy2vHtXE3lGyJspaS+2IfgZdrXrES+X8X0FBXCdjh8xEYZhAcsEzw8
nrN316NjdiPAk5/RjInrwqPmTbY/KMGAE+uWAsoVwQzBjwfjSoGQK/IksQEh75L3
UCKo4Uky/bUxeXuad6Hz4NTQTitV3Y4cDqb8hDxTvDMD/7KrDdYNvdBkEPQe4077
qyUEPsn2Q8XvqoEluYnRJGjzrGGM7Qk4a2L4TCAUUZyAqc1bsKpSiEsG6CydOUYD
yN64tP4mdvVD7WQz1K/JnqhMYJuU+BVgPwJ3727sDZ12o52gtZ9v8pDv7JkeYm7Y
Ls0tJwmdonuPO1Cjm5LBpTnKMGUibpchm2lZR+GGTp36X8gPtM31Js7XZ/9LwJRA
fsGL16CnJeh2RoACHRfcBQ9b8NCbXogH4ACREFw0N5Y5oNp01xprB0DHUeQj6/SR
fJ5PMNbrqaRxiih7s7pGZZtSTvuvj31JkclN7OEM8O9/NULCTENdG6IkWORgQCgU
qEJqNng4NYWa61SdXz3+0EN21gRIQQTVwHuqbAByALmClVw3Vrz1I6MdTDD0DNyj
8ogf2RaVFojH9LSsmTkqoBW/5xBlLvAHPhXLdlXrqaJjnl4NIn12PQMiabR/NE8D
BYYH9WNwkf+qyG67DkiAfToIdpPq1tT/01rsHV7Hfxg52exdCFhLCnRIzZJ2uMa4
x0I+xUVjsLufyrz72Gmvi8k5qXMa0dBiFG1R3mZg06z/EjbOAYdXu8tuaHtJq0Tc
LDHF9Lnst6okkNod1HvXwElwq0VtSJ5cAjKbPBDWssPN8kkb5AoLAyTuVzsnwN97
1B/1DFrXK0kPdd1SgFkotOyq2LsByVwsBDPli4nQxYtrUhLt3sCK1MbsN2UjKcm1
fHTQBM5f2aN34GYb639kkGAykgTvuZvoPr2Uxuo05fyOQDzNlkqv65hWGtC9tVFf
7cH+3FY9hJYQFHXny22xxF/0yn7lx141U+sTn1yuQiJTe2aM/cttXfH8ylkCz06k
rXB63iPJfjVFPMsw87mMKBmIGMD3vBTiF24/9w3va2pQpP1A7HhpI6J0sMUbCi/X
qJjoFcrbDHkLuKiLjDIp6HEJ/g63O+2lAadkNkZ4p83Or0f6jtgG4jSj9hSe/bQg
/ndIk9Ljphf8iUxYqjjgVfA4Hp5ruUfzvuYtgyL/In+NPY0i7RlITD9evXiD38VP
XGmpXb77BajlP9O6m7xHl/9Gh2tVa+AJ7Y9vv1Bm8oFIqKPuJScVHe65NrHoeKOT
o9JLfqF/RU8iLL1tW+Lpz2K4oNsTnJIZTp00GEjxgewp9rOQPBi6QfkPI7rpYVR1
sqaBcFbSos+Om+8c2nAQhx7793/OWqAjuZ9tDVCpr2sNRFHfwuyDFdlm1yqwOrMF
2ESdXkCnrzCbjmAn4/XltA7bzpWaHDRT2Mn/lXOcwyifzfFn72ibcQzHSgfO0cz5
Fbw1PuwqaYyOKU5O5CYeAMfpHvjb+eW+iFa92F+EuAC+1g7LD7n4K/KQcK4lxTQF
LKjgP/f9ecUuo1XtNBPihRg12QzSpZ3EFt4tE7y3H9fyNtBa5+FsUN4k/fNdxulw
dXAcQsxa2yb21k0UEsKcfsEuRkhwVfSYkMO/dsVV5DpqzBAQUqkfD7BjE46W5xDf
mOkNEo0Vkhu8OKFzKR7IoXwED/RafkhmOwIQFITyxGD9xs4qDMA3FsK8Ps6EwXFf
qYHrrJzyeb6QkuJgCDw4s2BSx/Jfc8rLSpnWyLDrG8GR7982x9QZHjGhcXuvU/Ky
DqsmOfXZL5mMlA+rT4jvOE2ROjlbW8xMAGIm3W429yz4zS1bBazLwqg8cCKZX7CC
9fAqeInSs18LCOhikdQrTSrKujx5yJ/fqMv2kRjLNEWOnPKla0pWiS9bmURFGKoh
hRp3az5RWJxfHi/rFz1gpdtpk1zMiDKhZ1ZRq0UB7RD+WlHQ7o8pLyxt8KjT+WLu
Ff5O3bC3Sl8SXdkic7Un7mULGeYrAU6ZXkoA34DdCB+3tg2Sf6CkP/Rve78kwwoR
Uf9BaS6pp3U6hal2IMhTsnB7xouIwrJJmcbUoMJ8cZVUwOxSViALWiaS6k6a7RPO
z6HRAYE45l1sr2hwna+Ub8OEAUge1SRXK2GDqx0bqf2oiusgxKsSmv8A3fV8eWQw
W3mDydUCxF8q9zmh1PqLFQw1365uktmOZhndvvSAFnzR8Qe4jV6XZLUXzp9qUgbB
ponj6Kd0Vp/dZI9cv3t7nMQlRKOJOkvF5cRIGkm93ptSTe3Hw+s8U1PQ30TVBft3
bgIJqF3BdisNuh490auSUKNoWyBuTW9Y72mkg8M8eVFHI6b6U3Spp4fDnW1jklLA
7zGszjSfG/Muc+1Q94Tt02eMW4HDQt0/g6wl2bxZ5ap2vCCWOWTcw+7QVyoj6Upu
HNBH0kl4wnnNZIT3Ry4zdbDr5Phua5zTCcjZWn46i86vrWX1wAZ7HglDKRrDGQLY
7paq4s/VFyv129B/YMrwEHf40h5SDtZnHtA9jbbzO2D17Qf2yZ1QEaQTj+0riTpD
dTJtfVzR5lB1L68g/9tjojetPGx7uLHieVGwbJKDAAQBTiiSjMDKx1fzRxU3cj1v
wB5SM/peLhp8dHyChMu2zIAEZSLj24ttHXvfEl/ctAE6UPuoAnF2lM9ocloHtSL5
MozgcQtxkgYtS9FOA/dG10RqiRgFt4hGaYrClw3ZVeCjb5dZYKCaDWMosFGuoNLf
dC/5JcHc9NCuccjNGIx/z3gtiewr0+JPUERbUrJKTOhp6P0t2/6licSH7EJjxBoX
hKjWZ+ZZvrr6oq+HCql4uieG/pb7wFPNM+uYq+1m33+aZhnxc7Oqj4HgWxRYsp17
+WNbQCBlWenqhl8U5n0fGRchs5bUbznwkfxP7ze7tTmUzqIlLI8W4KniO5729q8w
PgOqd8Ou5c94CPvrFbyCCVYf6g8cziW2lfhOd/aVw90aYQdaakab4zqB26rkKFRj
CKNG3MzmXUxMFR409+9oLICJUNhH1aLAtlk1ohz82kEwbz0sy43EEXnYgCDytD4J
HUizaVF+VU7R0E7u70z5/CRxlnxUSJnXh41JVwlp8oM/RBv0M9OLzy7kg71XYhlw
Sl5R/AU0fxSbAFFqdon+im0fAcnxbHfE4fU2MMNGgxY6xUU7l0m8CQVAWyNwgeVS
KgMcyofMVCOwdhFaM+gHBRAEoiuqik16sTPIW5c3irgh5yRM6A3+4K+nLgsa8dSe
oy7y1uoueTYc35GNLPv2LITvZvIKYMGga/deEqf5zsrRmtNADoKu12RIkFPBa1eY
fCJn5F8CF49+2UbLjZrsPlF9TyaTOFGfREfBk+FxvJlnJfhRDCp3W4BBKWbyd/Th
OlJuOVP8AplNXgr+SX3l93TlDiWK8qSg+cXJghKTpc3Y3qr7RAQl3EgpwLTphqpw
PtPw1PYeDw6QYivOoJWuMdeKkcun0NT5Lfg7Z6gFFYnvLuytLG9FhuF0R+EPEnVm
HIfYcbjr2fPKwngUCWGj8/n3X8qWDjWmRve7MZMqPsxnhvgZIankHVQ5/0uNxBq4
DK4BeqGtRvWocnlOr140TSgL+25J4qXvvcJjz8tPGsNVjEwDMNS94Rf1/Lb3Ua5b
gF/u9k63JtZGZqNOKNbmcXVyWtd6qI9z0TStNCmJz2K9uPqDKIKrmm1yKhui7d8V
cN8GaEiSInJpFsPant4coxAFPWn9y1du3R7NmTNYXvaKyzLK+H8qHtosT868AkAP
ELZwW3+kfJeU9FKuM8yQ6+bFtbJCougNHeC587B3VxA9dd9DxOwv5iVvstIueUFc
ImKQl9N88EqFQ13fs220ubdtoSta1DX/p7HlzwS5ZU05B8T1FQVN465q+pLV388h
2cLzVu2Z9bHTjqvzlpWgFFgNrcIMC+TWFyRhdE/PNBXOSJ3LmOOCMREeqeT/DOZW
dIkeu+OYYmkNYcOWdOq7lNj+DxnhQWCIeqbltnh0Yy7mrU44XCy3ztoMS35KurgO
a9bhjOhk13273JzCJLdZs/ZiNYamQeHq2qKgE9CJjDhsdLDXuQHC1wuO9qXNsLVX
o3t8WRBCffgN3Mic+mU5pdUgk76/tnws0GcPAbAWTX+8W9z0HmGqwMim5lENqHwj
WsrQs+NhWpmxRVej+eol+gOZ96VZ4GQ8UudvyWerJKsfLQ9Q10XFgRHV7NuvwJ+V
3JNeQl6ApEMUTfiLcpPaiBe5pqPz3FBCmB9NiM7u6jkXVoSREIfWsS71x0zm7FQ9
OpFhkJT2d1mkPNqI+h7iP9ZvN4yMmCXl/q60wSS0ULIuHZUfOnIvGeGoD/O1AyNt
9w0FntapEDvFzKut4GI53S3++SKw/8q77Tgaghd/nRZqGr49T67Zn5mKfyuR9AqY
NPqFgrpBQZAiva7CAUwMEiwHXpAQRUJTHmGjuqHRXPx+ZdAUieJMPkPiTQHwFJoB
E54GD8i8jsyGOwDxdJHFBte31dD0WR6oT2k9agQ+a1suPmtUU9dFDhd/goBGuWv/
ySbwYTe52AvpMGKt03MiRRAT+MZI9wgn8DD4p9nntrl3uh9c4WGnIilcx8bsl5io
wLdMYuUhSRwtp2360Gv7IHXpbEPjrbS5s27GDcu1jQU9OtDlZzVq1Z7OqMnnUVWw
Qn5+nZjkdbC26G/ZFbCWPqvXS1D8rvrD8xKmE8qCsSnMP0yNTpf8c+b8dL60j3kU
3xqMSGP6XvW2+G8abm9UwYu0ArjsV7/R1elpLu90a2K5K1DKRvSobNZ9yCY6MYYN
gqYgVgDw4fi4SelF9U8vdT0hSS78gRVs4WI4rR9BGon699GNVrGR91bdDNk+OUSB
5JPfZVHroUUDfPFR6RxStI9QbWzXesszLvm4RmnYC2qYJuwFAdvLgkQ9yuujUIu7
Vm7jxmudMrLVm5XdFeecNy1kTweG5Vt1byXzFRxiFgyaS0hRMG9ylsoT916P1jS+
621RFaL1EDKJ/MXJQRYZ8/Q5cHNswhoiGCvL3Vtjz61eh9i/lK3zADfCS86SjSei
4MlYnRjhdvoZ8UEJn7na6ZCiyeo7VKm40LhSWFIc7j07MUGoq4k+KPaX+w+cwmL4
L7pLeqOv4G1A/+HO7rHq1RLZ3OqrGZQRseO/8ZrNY/PbbxpcSsYhdfu40TAaF9v7
/6YOuk/VHOEDuCKv5L8d2etJyQJ71AbF6gtzi/AjRhNbYgN1Ca7pQcv8qN+MYC75
UgGDeKK+0yvKIsZcV9m4uxY+SUGdhNl+t/8r6GUbiWXUS4gJmaPZx7D1qE364Y7R
nbIvcWs2cCj0k1jcDV2vOYC8dHfdlmTCf8d2LuxwRA/MywPnZ74Hme/p/N3cnAqQ
4FteDtyVLOcGWEzdW3qrHg8oT/06tDR4X/m1vlhl93hiKUQgDubstRJ3IS2b+oeh
pLvJX/B6YjCtakF7IO/pNbVSVp5seZb4HIgZY27ZFvmTRoh+fSZBa0UgnzrZDuMl
svGyyR2FkwGr/Nm3sI+g5I2k9TMtzkCsVDNNQH4ag8H3BbW+KYIu1XxUBWnymEV7
HBglVDcFm8MIO3LWi1K+QubsDShSXtYOP9fkbLKu3CSjXHGAhAK59+YRfst68EeV
wqKri/WkHNGY7pPD2f5OEqCF3IseTJCBEqePgM9jcA2THmkPiGen14IbinR36lfb
KwN6+fKlriuiaV3ZGI6WTIfA0oZxYz+x/5iy0SsGFUa6D3xtim18S8vpeGq6smxq
u7hUrZ+gv5dEDK647V3sngXWUjstEq7p8wlld24y0DUTY26bbrDd1EiWfI9g2lQN
CeZ6WM0dlkFK36OTxUnuh2+EJDIYTL9LKXVPPjAnehSU3W/bTfXNM1C1NrJ5PdlO
3V3J5mBXlkJlmFkjJiwYuqWuVzGI3vAleWy3V4/DpB+bsL/owHESLIN4sJ5y0k3W
xlT6ifTrSXU6uAbYkaYCsu1ofqrS1CyoB2c/w9mGe99wj1afQ26wgUG86dvTcvJa
Ty1e0QeQZclmYnTVGTuKur4A8V6GIl76DMM0j7a9QQMEOSrOBQe5cdS7ZKE2RATJ
abfiCkpZtClk072GoxluKb7TuR2ho+R7J7cIkNEeuo/7xSpr1wSWgOKmLxe9jCCT
K4yJGp3P1R2ixtbAPTYKwnt89ocFNbao/CFwJO7wMR6uDlvP1kN7SpW4mZAjNn+A
a3hgT+S0i0npQzgKf0KGfjje3NAw57Vgkd7VicJj6blh3pSpziOK53xLGG4ayrvV
1HD/hEFLPyH1N/ZwyE4KBxNiABHJs9qKptpLqDlhuM3DzOagFD6ByXaXXJTsE9l0
KI8I4tdiLahuVj83AraDMTrUVoaJsvF3YZRLIK8ij3MK9EHwLMk6xqCHkxM0kwNH
bLXQkyRD1jzmink0ZCWqx4kYXxbzR2XznadE+WuKdtkhLrfBG99RqgwMG17G9WYf
vBisBzx48ir1kKKA/creiYUaTl2ZP5I3CuBcgiEvBXUr4o4mN8LOa3dpXKvVl++5
/rj0PgdHXmeBR3BoLTczilhF7OxuqoycohIWRCVKX0+1MUaB1mPUdgwXh2OphR20
AMhZwXlrxnhcmtAlvZ8CEliAvCNrV1isyBk0x2VygNbigbLZPI4vbQ4uFzDn6LhD
0YjtoA2qsX/7buJk4ehZAeIyyD/ontaO/fzsmxcbjVvWIQFzV5hyQNoHNo/Od3Oo
4De0aiYTqRVw/LFuhO65xniqbBq3smicSZ6EQOb0koHicZwEeh0eSjhyklOiMmqu
PNLLRIoXRh5ezSFM2gUs5HOsYNkWkp1T481ebg/WrPA3KZLGeFof+1978z79lPM6
LAD77nZmaZNmGKOSCEWMYYEUUJcl3MWJrNIegh4sX1V7Me8g6qUshS3+E4WsNAnq
izydpxm+PM9tdM1pcK7TYMS0wQsXmoPcvB4sp+Ai0iMaWHBYSFyD6DE5w/SuXLqM
cG1OpmXlMMeXHCa1euu9D+GfH1OShnUirLC95CaO+/ZXMWM9VuXseK5kHMBOdFrC
aCDTi0pvapTtFvECZMwil37aFMcUR6fW95PwyzVScqFGk+F/CX2rK1QzkJccQK3f
SiIgSfyoTYhzdfOQbbtIG9A/7ps0bZsGoSgsDug5I0Mrr5GBbqo7Yp9hqTo8/uIZ
JXitmcwSGXUSpyKkQfHZi2UPfuhpWBVs3jpXfceeeXkkIPnvtvGkc7Vqcze8DaKt
pNHiDozWeZ60yE4Uuzy6d8yvkP6VwRBwUKds9ryIoLfedBWNdPci8nHF+BMqGkUj
cziLfeBNuidO2zxY/zRDKR/uv4T/DBup7ypgwaqNhCOiM1mQzVG5MK6WRDr9s+Tp
M/yi8ciNTp4llMS0vHWQhG7UgPiBpIwh9jpyq5ZRnubG7/RGM7FIfnKFNexbB4oC
rLr23EJR7yxxwVZNi731WpJC20LeAKhcFmU8yW8fL+e/Tjg606vSgoO8aT71HRP+
AJ0vPM3Xpn47LSFDxMmIaiEVWdpCK8lnOrxM7r3yKbb2919UCxmpilrOEJ7bev6T
1kKn/ZBy6ZXR8wkZ/mpPYkJleh6kiXL5bnLpd6eK/+wKp9KrL1anhseXX9ORMzJ8
p8oQmg4C4eTjmyhBJc/4ACiuZdlYrTz+p5viP4fVBbMlVDXF96bv+wVe4Ee2kddy
4SHrm0SP83ZIxuhaGkKvXLbj3aqE7rdnAFhEw/7QpTpfUuYU/NqYTZqEHF7BVjG2
0hPB2OA+1akYOJQ6b8W7DpYWHQVI6PKPY6X2UNqFSl5ZY6IaY3axFeySOXjWb4xO
OWY7ONUbjph+2ojXpsFs2Co8NxI4nwENcuyaTomXw1FZPyr5GYt07MmHFKF3mWUd
Tyr0OfYu1rlYAqxed/DPQbwDcgQX612yAzJ3yBbFFn4E/xll20Sx7XAG/+srQonx
LoHeIWctRALUluPEJ1aEuhF+nOArVVh2U5mJmstwpg4zP1qzZXO51jUS49YlYB/9
xDPGK/toiAM+8XVbuyQbpX/X2L7i6+UtOcxlyZNR68F6X3V8IRXrMzR2aphykRdT
x+XGsrYfkTV8GU7goBkVvwjPhoEsC1jLRfGSdhfeoialxHzUEme9bDqK2WtxuvMR
enDH5FV7jtO7m+KPh8z1d47cbO5r1oY5hvqq8VnbJ09Y6wdqMVhFNdmG6jiF/iHW
OmQ4CMfra2bYz5fQTWn1cDIGzHf+miNowtBZMt9ejwAcEU4TeZ15p6XV84l9OqE2
gWXBcuTfqs6M6O8uD3BOZJDfwdo0MB0WwgXKGixeZLdxfgD+pIU6TlFlMQdMn87o
Gf4ZKAMZFZVQGB2+f5RSkZPWwTXrdmWAuIsisYTrfYdLTeLzyBp9c0zcqyNhKZMx
fB96pgQJLyMmHdwTqV9EEtlA27XXfWJBTyz6thtqHLi3pNeY8rFd96PA1yi7TgDL
6prvNYE/xRF/YvJiNNAxwn9PVAAeP9bBWGAWIWSrJxx2o3JsBmsuW+4aSHyUuxq8
ugOn7MeBnVPsTonVPV0mlRb05k65MEMemzp1VAKarbsOrny1hQBUVYQLQ87cyts0
PlSFScpphlc03u/gKzzD/G0xHgNrRzTbUzbuEmHKjDecpSWU+qp9rF26/PMuUS8B
jpZ18Z9aMtEwO6RZ1wsr1iu9koq/M8Vj2L5ZRodbru6MxI3/7qWqF5d9aqznV6Sw
n/VNG6yQ/0zvF/E5hxrnsFljWC3rHhUsqGfPLrmEkmvlwX6Y4ERV3++d7Vj+P1gH
c8t7OOgYKkFg9ItEg/f4Hqz+ego0KTi4FkomzKqE8yEpouvv+6hV3Pq8DEjYAYV0
TwxC69V5vDqUBssIvaN7KoERk2IptLUgHaTZ3vnbJeeiRPPKY7/b2TaXcghl7k70
5+DaICViuglX0ZkAFK+NLqZjQ3jGBQ5p1I0O2W096g5Eke99h4HIgsLguqGmwFBN
SDJbILafiWDAK6zt9CyGbSqevtQ+ADLRmYAOCQpUmayXubpkg13XAP5Q1AOSo09o
JkNDt2XH9JLfFsesLHp/hu6tyvtmySlmSIV+TWl2qwJXVat2pz4La6HDlCsGWL+Q
lxpM/oyp6Z27dSB6HCEPgIJfT40/YJ3ve5kT9zixK5BFRAH+1XqY6NbDOp86bpcr
aH42BhD3fvbzX2GSInAloU+ZAZVK3/mzUy2+C20isF8sUsTB0jf0CngpK56HW/4f
Jwmz/c0tCB92TZuaWwyxBR/Qa7lPTdQ6l0Z6L0Izf0YMibGxkFMZBM7xrEot+9ie
c3rTWU5eY5aB8Qze13YHQkqQujmFWYHTcU4yOc9I1WZN92Kv/5+gN6ayeVlAIj27
/m3Exd0SfFB3RjJbzlx3cjQL/ozeYvIyGliAi9HvPf6yJALakxDF48o6M3lVHCTy
lE7lBVpHOiOdHRq9Aip0WmruZ0R/xQDMWKdmVmYv2Pk9JBrbXe6hZaoUP5+mvi16
hkzYQvRkQkcA1hr3w402I2y88CqiXD+ZQHr8Stt9utkA/93D9KSBT59RBid+T1Y7
0a+c/SalNQQ06j5mAZKMyUDcb9Kjp9zFI3egAWwgsPte6aFC5Q1nTh4DuUNAyMN1
fE5UFWeRTxrlFR+3Givwt3eZd/OqBqLg8bZo8LJeVM+O6ImuTLglIo55A60x3Lty
fQD/fubvGm8v1QTiq6q5jX+cCPuEbUFROgSG1Xsnr97mRKTPfbs9RFFiDlALEc9L
ehLd/0EJVEccXRhvsncdfi54gNEsA9ksICCR3yOaQUtZLJvIDGI08/qCeDO1Ia+F
1TtOIY7SKKlWjGk5xmah81XThfjLj9GjpoyyLFWI8vB0AHCkvMWXYFdFaqIKowNe
1jUk1zLJeKQy6CUH3lKBH8waYOTKGqryNoH0GOSVbO9AMWzQ2+Sfviz1ouwdstLi
WSN7QrVEFPRfP77o2ze6fa5RBVk9WjQgDAHCKjvQBYh81Ov1+CxO1qXOx5q7FWHC
fRPQ9KnxzijhT3JhThGPvUkdlnIXi8IpuO7/xTTlY5/tPdJHuMgCQeH+aAQeXApE
55Gvk88P6kmncj4gf67ksuFjA6lOS+J05wVxeYNtwoGsKzM6LaFATJOtbwyw8yJz
Zl1CeJlDoKFOh2T53hzS1by2E7j8nF2NnVgpILEDn9HgwQmknRR4OU2TILpQqouJ
idNGnAR1UXArqvoc9esw4uieISmGv37Gwlmw32tnJZNeZRjRaXRW1fkDb/kzGNMk
UZWxcZVsNTwxy3Nq0gQZvz5QsGrBukePAo0ioTc9Y9DGbRBISSOk10xn3Wp2l65i
LE3F938Qs/Kh9XVqp84C2bcz+XWUc094zEy+Oas/aE+dFH5Xl/980R0CYXbuu43e
ozR9Ch6WfDST//GIvAvP+Gxah8KeiAeq5JUOrgTF7jLVqc6NHgruQWse0Svjg4vf
4SLqoF/reFqE/HsOzUDJjFcJpERfZCdSHs9jzdSqs0Pi2RHvVqCND5uWg1j0tfxx
OiGkEglKUpYheAySGsUWWspPBUC+bLMtyIczQ58g/PPNKN3SNvUlwQvW42h5vUDA
3y6T8QOftFttnYATGCoVuhGke7+WtQko9Hg9nTLl04TNJhTeV377OiWeesUVMWjT
X2lTochFyjfrXiR3X0XoNcxrSjofTtKIgiHPpR4YECDLQE6Q0w9DVUokft98HgzR
HlrRMj8qoMNrR3fb60RGd1iwIWHnq8yKipeP1TmquDghRfp1hUWtJACnZJbqlFiM
EZ2QoF6TgBMdeUepk7LV+zGW3/QX9e78gBiiJq05W/8WpNZwmr+hSG+egFcPhgdN
Jado7wWvNUfRDwHdi1e1RNpudp6dM5xiUe1HrBAZeDJsnjDBUawxtbH9q46h9gZf
myzFU003gWgGIJDQUtfN37RVSTpjyKwX9FhvFTboO/iAnkSDblFct4Pnq6x6kb5+
gZUR9NjFEC7tpJDowm2iT50sLZgwsGzugEkny3j41BX5e+e5m9CJh9jqYhEgN8Sl
+Z1VWa8FP5ZphRGuEXCOSy7iGlKiKESE2Dlt/+mipTR31W1jTGJQgPR9HeIhMJU8
Wv1YvmQU8bIiqgUQNJ0to4plNmpghtxOyMjF2v/MhO0iqemdzo8a+hOTGfrZE5uA
d6u95B3TBqpr2kFWWnM031JzmMoNZXzwEipI+hYSRQoSaTCJaMZUL8M4xSA1zxjJ
UhViTX1liVrE/adKMR712JYF0+THrTxk4K5SRj1dOlzANdA/FnqoK+yQ/SekQnyv
ZMLAMKbbPoun1hNdh+rFlfueQGhSMjK5izIi0OX6aOFjxeDWNcVX8S5vQhL7t4zO
1rw5n1iMUbaNOBGb89Eik8KXI4vSVY5rslX85vTp8twqk2XSn9aaY6BvOJ2nBR77
kP+6jCvrrqnElhl8lIBcji5ygBJuAsybil1EGyF3v56Sfz+WvOPZIg1MHPbSW6Qi
paLO+kYIcGyoi5SUQmwFRqzLaww410nzUaWSflTainuyH+R2LPNNuxwleij0o79J
zLg7gJpu2fVhwuc4l5NrCaCCwSbnADewxYq2LhrFI1BwXPo2prk+VLhkYH/0h0u7
4S8zPaQ30dojk7/9vg+5JwLMVpF7gOkZnHLGpFv7fDYjZmbCRVPDI9pwuEH1oA+0
EsQD+GDbDP4lkHByx6zcAfOfLqN3YsuR89WTMu84U0EUMkEHXDI1nIIYqQmFPf0N
3cEXPHYYCYTRXpEj69Ftdp9PbleaTKh5bnePbkADdEkBWuUEGHQ/q37EyRG+RsOX
SHpqxWTOBTBHw8JK5cwEzRaYlqkFwF3nqsT8h+cX+P1chkcNKU/1ieGEiXZdo2HB
wxj89L7dX5B1OPm1bXzWit8xRHCAyAS0eDn6cm+xk0n6H76zwj/8aRtPqZMVEimz
gYcBP1zM+Bw3Iey8gD9JnQ3+bxGdB8/zv9FbkivYMdBYFlD0lq/r8Ua6jSO7vTNj
1IHD9zHLicrXDLiJJaDlxXCNNpp95bLDom7TcUfv7mBoWvaxXJEjiMJgbcaWFzag
U74w23MW/pjwVEw7HMC4WAVL6iJIn4lB/gbzlzA44PSlUwjrzaYyDpFhpAlGrNcS
pUQyCN56hwFkb+spt6T71BhTdaUiA/RhiMs8g69/RSwyZ4dvBLYZJjQNL9lfBlCX
GLPz480QxtklcR1aMOmaYTL8TafuBvM2NA2LfFOV83I=
//pragma protect end_data_block
//pragma protect digest_block
ViZT99hydlPJFBIYjKNvHEIhHM0=
//pragma protect end_digest_block
//pragma protect end_protected
