// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GxjxbhKg9rPT++heJAoDjybcEmIqbWw6VZcrsOhezVCCqT3sOzXQQhOFwsvm
Ij+lygmxBpOio4rcyXubiwhKRqwhz77XlIPlKfWaVDLE9XFCAVCdk/GLW4pU
OOX9gQ20/CQUvHO6l8u3t8eFjW6OpsxehcidxnmqNR4vUw9Q4D6hwvXZgWI5
9GSuZaVe0Q3arIqxmYHL4se+v/SFZIybldSWJ7rvXuBu/e2gV6qXQ7LYny2R
mSz7A5CmoXSiaTVZlkH/hTmTGLakw03FGoODs9eeL4hIrVN+yieeRNRrxfdL
0eL6HMH/CV32LfbbCDvNPkeKE/EgHmDTSv8KTJWU6w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VwxsRERZmO23hRnmdjhFvnQkkzDAnK4CgtWQYVmgElLD48zL0haMWoKIkSIl
H81pswtHzUNj3dW2C7Gpsw9vZ0VLvIbnSbe/eNv3IoTKUyT+LK2lT4gT41Y7
l4Rcs7PH84oxYvD5Cm4cpcSOOEo0R6DJ5i/3zi++6u2y86bia0uriYlzxnbr
ZvYpRUYF/u+R5o4MMyHg9eH5+IrMs37/91UUH1kt3r4N+teAxz+O2+OtJvu5
K0aKihaozljYz6K5pc59kUYsz2R3qzxENDarVomMs0hu6WhGYlfbhFayF/zs
rxmCBtt5zG90HwLCGWLFRESixk4MjhVb3WycFmIdlg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
G6C74GRquLYZFu4GoBxUF6XVBAJ1vTfll9+nDNPVnLh4qx91D0bqR8yHXU0m
0xcZ3v0vCZ6KBwX8cBmzvrDLK3sgY7H7nFKCpOAtBWnn8BKHLrDFHS8GqD6/
Ueu1lf+F+l0keNYpvxHe/6nbnfoPPeE5h2gpyaaCHPtEj6WzlSL8HV8voglP
MF0xQY6JHkaOaTakHKXlouvyJbfLRgy1IJbCAGdM19D0f3OcT4fmEyh2V0Bz
7wbbikLhThlCwL9rdVKNt1XIqz5NGHUNxeRk4KhC+27GDleaImivHTndu6Kn
LDgSFasnlyi5yyVB7CKn451XmarFTq0ZHUqnqI/z6g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pfaDELyxSpQok4z7tK4sZHhUMBKuIll3Wg4LFaUtNiNSJUEenMJTPo7Ux0XM
+a5/KBu3VJ0t8AFxxSf57GlWshP0aTl1yfOMvEa2QyMWHY3nx6YU+Gjq4m0h
OPlnhtzgpkfbY9en4feIlHyDzZeiSxiYU+/1LtTt/VYPwOr8kYI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dHkA17YIPFn/YU6oHTOB7/+Y8A0HICeyCfBHKMj/Kt7Bdty6tXdBPclivs68
B2I+qP0sIduRzSwGsWaKL1xt2yvj7NwnYNApN5Ss6t2YzrTJ+4JYXMXQSUJv
/AN0D7SFF8n9oS7CW7zWIsfRLRyW165Zh/TmcwJ1U/SIKeHrMefBOxTJbZWx
ns7P01XjJxUFwTVQIQ0XQcioQHbVjwfOF9LGvCbgDvIbGtFosLu+Z1q7bweQ
0CSdTtRx/pAKbJBcqirxJdlAy07CvkHYCnxIk8A/JVYSxxFfEj6pOo2bRk4t
vz3+ouoTJJ38wS2Z6D91fyprtjA6O1DbJX/Ut6qT17fOSlCQEi4/lOioXs8A
4CxabJS4gWiJmFQPiImSfBgqbS19LGpXz1vE7U9omNxzQpUUKuOi29soU2eG
Ws2OEeagVpQjkLr6GxG5WgVgeeUMGO39F7D+bvQrIy4iRK99d6FSeYXg2xdF
usyl5fUl9VTcBs/eT0iFNc5zKj6yjyrB


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Sn43piosbdB40fHz95/d8YV1+3UhWQlIoMFpGAnW0m1eEshraVNctrajfEWv
nI3z9IIl4gqkswzFUM+7CiOQkkKQG1oFGORxUWo7ylVyTaKTFM2bC0u3AqQe
4rGf0BnDGp475dWPG9o6Gs/EB+LzxRz5Uo29B4cAwp/NqGGTTfM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ue3jEBfkZmgt9AZAbnMuHP7fqUcwjHtNCk3AaUXBvsx9XRFMrxCmVpanY6+q
pxmg2T0lCOIM1C7SMlAZ9IM42QoDH9sWUGPw1ylvoMOsna0F9kzRxkRxzdR3
KmMpsda5rwgJ5M71sWSx/yk9nLvlfpCX1GwITgD0ryJrPXSz5dg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 75232)
`pragma protect data_block
CuFm18kXHCWMJwqTgDCAAwBOcWFcArqWQJEyf60Y2ha8FKsqEAVFMCdzGMaY
Q0ZXQ4fxtXVwCmn9+aH2jwky0ep/X12m4tqAqKUqNOk/AozARTZqbHfdLQ9Q
2pDe0BodMTM0LjZ/i8wC6RSjOcJ3MnKeCNYvO5h84VUsKbC/yP2VwC2qEBFG
EjN8KspaBP4137BnXASggW3n0l7ZW+aFpQvGQbqkEuOw+T+D/cTETHrJZMUQ
75Oe9bvDmIwPbcWUM1UB4wHN3dIRN/IRABK32zHC2h58lVrs/KCuqNCfv7J5
ioElITOSDTPmgKBWROeZkDAnJGOeVoAUN19vDAdKE3kXqD/gXr4jvwkj3tYB
ASDojCfzaZGNJcaXVABRs7tw9b613in+Al5vC5c1KWRyhfOWaHhAUn1X9y/M
fKWUH9ri2FLOXUFzW+UMGGmOtCcyGmm33nVZbADj9foTrKN3x/TZcKWnOfEj
NdARbHnKHXDC+VHYfRuXIgLnB5q8vlrG1Rfcn3XJ/kO/0uwVDcL+vf5wDWJG
HHLX/2Wgnx9remdPineiqdmQw/qyZNkrTmW1tLOHPoAEFOt1kL1tiH1PqEH2
MOnmdlNVaJBGAiw0Bdcqag/FKXtLUDd7GKC8T9Hg8MzM72myWul+jZYGsokA
0sq4odpaWAObkZ2EHyn8WGX32LXvJMsvzpyQI9CYLtf/ZVoWJAkKWbcVwJSk
RzMn6w3JVrVPEjd/AncCBX7EcBuqyH+QYEOCC7HoNL13aSHVnrdvesPnb/+1
dwbObwQkoVHsdMOPedM7IZetXF6uBH0zObmL17j0Ye1EzuE8f8P6YEwvt5eR
rZ3pj18WYMYrsVRYKF2659IJd+yUpsw4ZKfwb1XJNVOvIS/vSNMvg5aEjoBJ
igdL7I1oGEtSBjI8rfnRRGsxEwkjRP6FkmFXg2LyNGwTMW5YY8+5jCD2iC7V
MdAb9FHAXE2sBlKHmvEfESlRLHWcmHsUSaVp8hDE8JKIGlsYs8KKcUqODCqg
hhjAg8qwMoH+DZEEjeBMQfOlGquh7VFXjkmR2P0wgi81H1Ikj3QL0Lg8M7M7
R4AYdHyivv4ZnIsLyJiCth0VhKBLlBcR1KxF7k3FLqC2ga2Rd47hlbcWHQy0
zsdSuTY3+xy7CsIS7LptKks5N3nqWuZbzu6kg3ASSS7eIUC+mDIybEC7/JyY
tcDXI1XAyFfN5Q+giwESt5x5BiQVFN/FfDoe4CIYhdUk3JrgeNaSHFA0Ge/q
uLOvCDdjQHIIOmEG3Xd0RGeMu1umKhyLOMa741HnfNYXBiy4FuzfCJ1+F8Gr
zpi5xeQFoUUkGtXugz6gQBB6OtWqB3Qe3TJbDOFIei5v4snTGUMjC6nWwH08
IzVpjCSlieP3Pp0X1vulJv51C1sywnzwn7LmvlDZaPE1CR0A+vetngINPa9l
w42D9YBs71jWT1BXnbNR6VRDIBut/4pQLLWSZYlrbwI+tTB4Q0rBiUZmO6am
twT57PfIAl1QyMv18e8VQMVw/iMjBYTxDl/v2BN5kKSl2qK0ul4fXCQIpYGD
B0yag8HT8d9+BJRd4bmPH4ImNpTJ4S6Lm+qs4P7Y5+3tYtA8PMoIBY+yU9pI
owsLPy4td7rSG13wdy7KEtyWGDkpGrlIlTao3CIqfdrqfc7I4hJc8FObQzmy
rA7vle7qg4sx6PiXROWxEQjkCyBnCGCrSChcvI5+gFtpWZM2wQn63bqwjC6+
l4eZo7BTJiI4YiIagMTd0PnHtJo4D8VGoHK5kZvNoGQc32OCH513s1XB/OOG
G3T+UKzwyjT0l0fBQVAyye6S3hEIPO7I/0+KC+djpOBk6tq2djwDSUGfGsY2
jCXTOINN9FNN2lNCD9uNp7suujBsRURdKMT96mN2pCu11sT9BTMoJvJaXE/q
oOw6Ji6DUw9ewO1bzWvS1ZclxVxD2vLBoykVCCtjK6J0BHjGzja4LbEcwQK8
tSkvx4Zg8kzc2oIABEZ84O36VflMKn/eYEa87NZIb0vKKO858I90V9MHsg4X
eQyxxCy2iJ1Tv5nJD5q8X93hJ6x5t4blFYeql/LILpKymqgk8/5gIQmBMOEL
ZObHClOLL0Ekb6zMGxiSENWttbom/0el9nklwIx0ItaeEZF4Iu78t1N9wdTB
XFcA9sLQ3bgnfTi7ve0cfSP/ezwC+Ye/HNp/sj2SCMMtsJUKM4Z3XBSDRu7Z
dwJxEncazsb6w4edS/T9T2GvXYyeXzCyr4xOQCW03zz1wfJ7BNkhKzJUTYR7
/M07O/+YWYTAh+8u0irBHCR8eahxvcOeWyW8kc9VfEj5FFgO8/MlBFnZVuZb
uDMev2oJS3edxNtTo3O3gGef6OWwtD6WvKMU5SPZWIB8Xyu+s6OXATBfmyNU
N+reAuru9d7xOqJ9VXYMInQq8rJMo0aFfTrIP/3tzee4VkLMZ2D0KzhIvcrk
XYdhYw2BJF2e5ihGt5+/bHhdFG9GCDoZ73X0sCK5wkgG37CAfR1Lp9A7WqH9
bre83WwNP9/262IFLrNNsXmAT5UYZHuBrN6flnrCOtMVwrtNJOtp/+/Mb0X7
NbSTKvODDVhVZ4NdqU+2DselJZuzb0yORFniPpXju1Ro/vjYABVyXeD+VcbI
x2pKzGbrJqvgYyThauoYCHIoe1/z1RSjhhA+BFy9wNavFVToZzoSMO/pQbbc
t3XNFUYCvg585ATa+kPb/eLeLoYcfoPF0twQmK4BHetNDLyB2ZPrgSNjUah5
oRsaqYi/GVONHGvzaknm/WMf4TkA59YnxUTXuLrPmhsMqSyuT64wbneQdkG7
apF6n1ded+muLFLvon3araVMIr4+tv9yVMvu9gpaC5n1OojVtzkB9A5MkNwa
FGl3s0LHEbjXqtSN1LvLW3ArVWIzZpknyOVu4DawFlkQtcjv3dZibsYS5oTz
3b5X2G6xKdudrUP1lXqDf/6weyay+QiMUCwCEp+zmdwdwBIphA34k8WTgkhl
2DK+9Ga6NWzSCuvtHZdF/ToZqCYyieje1sTynwUgipaNVs21flPZ2xvtNQqw
4K+JZRNVFms589A7oXhDFtSwnre/aGJTjJXulkH40bQmInastVxQCFXTN6eS
kmm7McDGU3VYOdMRwxS62siJCWZTr+WgQ9lNBnnSeJ8PEXMDcgE6nNWb43Hr
RPZm9QgJqvF3mYsfyMqU8SHaVbixoy9l6THbUZq/AjONODn5pdKEOpAUMITz
1ljEuoIzKKgnPVDw8b44T2Vi0pVAoZXR21oyT0Eea6Pjo3gp+My+VahNg2u8
T/XKzm1jMWtWmrfJ7yS4s8GZqVXqmXWAD7zMDo3/J2vGnR/zb64pWmsb6vLV
OKRPoQa43+h+AlJRcK67VOZZo4Gd4VXBoUfgSrbw7QLFf85IiQzMMsQEbYQv
iCFEnWcP6EMgKshK/WGc6CY5jwMci+m4A9XBUncxiBizNXqJjo8XV5/CS5/0
R95+J7+cijDJ+hHO5Nb5AQ7QjjK27PkEFfwaSd2fsfeD6MCC/kiOMols9gFg
5SFDQIdd1eYsaP0d3vbvm9NbzpjSkfUvhKImTNNtamaWLCF3IULeS2/aEdd5
e0v2olieObpXsGkKwkXIPv1QuKjeBvNkWs0Unz0wNOsbh558Zh1zvO06dNfj
r6cjqesktqS3ZNAJLMb+23S4RK9Jp6oWQH8qIS6ghC12o8hprDxFQKbi7NqZ
usmcWD24TuqmIMOK08jLCSm7QIpODkQqec359ipaKsoJfrD7g+8blUNi/fA/
4F2xJHYPuie1lc2vfQkzdH68DWezoKHAQaWvNX3yXGdUAIIgz/EvJuLrG3cx
wjpmmjmnvUSZkcdOT76xL12A2+gKsf+z7Cu60TvUXyOgx18k6wrX9jhu1Ayx
F3zwUJrlnCwV+WJn1F2xZAYQ1zrfnxo1qaP6ZZS6bZWMGu1nipOT2QAoIEjd
8y4x+Y+hrReI9XLyrlEBg3CZOtSdwzr0uBwaKXOu4KrBA5DSysFXyFuoBE/r
y6oTgU+I1oKk8JIQgZDwiURfPfEi//8fnepySA9c8K2DGXYZuj8FIS4wdDVT
jtVRMrxIq+cBIa8oF41NLzWW4xHpZkQ8G8mH1KDakvMWt9fuBwhUEwD725WA
Qk7RvmjVNXZydhre7x1CD8Q87w+LuJONFgKG9mTjDIKkYooMQd6v1LZIT3z5
X3/3px9vFEUyilpI5n2t2i0ehzu+5Tr3AkY+isfUUO7bpidWwHX7EvxdUIWS
nS/s/NBm8FlxnrDtvdygTpKXH0/yubAMdkO6txsvBJ44LFqigr4rJNECV4TM
cAmMkx7oo3or2LFUkc19j5mrVni1c6i8iSyIvxADAwZNhApFFX4Xh3VmuIN3
gdvJIYYSptCA5kM4YcQldlpGkQ0YkN24s9FlHFy/5d1aXc/j9iKu2/S+c5z9
HOiV4LtCb78bRVJpITvKxLqiC9sY5fE/qtzbMVABrpmVQR8lyhybHxeg70dU
eOd2DWE+VhVodKoMfKFqJxYlaiTp96vFg6+3+hYtwVguVrsX9/JRZaMXE/mx
vS8QMvRh3CwwgwZzr/ioDAKVp294kf1jIH+vo96hVTyfLUUhr9AzFd67kiFV
M/fmNy6czoNiRZpbEKM4oOpyXp6cYhxSlq+Toj//qUD1hqrggv63GE/+rtba
MhDv4/y+t/SSxl71xfamHOCIkk2aJDN4eJm+lWhT53WE34gUQb7p0yq1atzy
N5f/+cfwDqlzwwgI5vuPRcXaGOMSiRVpXg1OwwLH6oSnjkpsxsCPcewROc7S
u/onSjaDBegOJz+yVOJgdNObAbtCQcwya02oif3iyfBbjPKhwXcOeNkBnY3/
UOJQ6TVe7nTIVSIWqowyKLhbGdiZ9S/teHBgH0EceXPCO8nkDBHERYUcmfcV
aQHrZwPP4LYvXmSvHF5vJAFnH03Hkl3XaAiTgI9hdpYAI0ccXGFLMvPAl5mT
CxfPD/BbVy6dE8hit2BfdE0JoU7Ff1S6GceiphIKStNx+IILt732T5maggD8
vmuoqkzwsc6HCVbCxRnwKWKCmB0aR1NRDbh63Gnsd1GH7ECCNaxXBq3PEcoh
go0Z46ZJeVcsYhukc24rIWxMCXFs5fklkMPf7aa8obhl7OeA0GQQ+TYUJrN6
JdTbObJ5/82LFftwVB0wgROcq60Qc2B0ix8AlmpmDlibGxM7VWtp2z8VrY0t
kmIgZcwZAMiAn3dYaXxl2O4FI+T2Ym84UyjQN/FuXKuQ4g7LZZV8n29kY4OA
GZq4ddmqF3UlKKByatNm9YVKCCON+Lth5+Kj18/vCxoAlFl5gqQj0CN0ffbx
rGbB8hO+jleNDjNgXwRVgQFkpNK48quNVtOHUXrfIKwRgZLCVKSEIZik5LNT
gFhhwZAcZEPYUs6YsQH1ZtmGP1yz2TGfYCvg+ZOQI9F7uAabulQcwDSB8cGJ
XNOTkk8y0Np9usYrxkfANbzaYvC6y4dMr2E5iua5BxN8E6V525cueLeIoOlZ
ZCRrK/UF5HkJaAKICgWcQABpBwoHeVBbKRiXmZ5nnHmNRJyw83f2I/MM00nM
fbv1tYk43h5yVrgW8BI4Qq1j54uGDOAwqTgh3cJBAIrbJ2BXj6FrsM2XyBZY
7Ts2/KBlDSKZc1PHkJimcfHViU9cfMGDLyQZZ++KgjOG2G4rbQn4WRgjnL3g
sytJQotusi17oHk+P4cSz24ztiF9lPAYBdqWPzp+iv+Y7TIThjRT1lBnkXHW
OMI4AE25O13gyieJk/iz1+VmS4vnXMhETjjMcjifbzFuBXq3gF+S7djGNB0T
Eu+w/yyiD8q3INxhMakicBDZhpMm26DeXZyrrkqVEX85BtIz9UGFrqclknrQ
8shtR1SucCSvMshvvG84B3QoISk9hbCg5bmjCX9mIKqGD1QzDyb0pGOi46yP
XhsodaoEk4aJi0G92M4s4jsw6sEBuHvoximT3vmGpa/RSA21ktiJbcbpSvD0
plsC5z3/iYajbDv4SeETF5wCnuZXju/u5wwECJp9k4CJ7iyeaQaR19ghNl3u
mMDpowg5JGt5we2PIx6y1OxwtyEZmfxBh33B1JgH6hN7D77NlwGKVANF/z57
sx4W1sH5ubq2zfMvLq9VuUymS5EcrICgWOKIj0D69AcF5eVINtMuMCKoct2s
BkkIVYnxz6sYTwwxCerS63sEZuEpeKkuXYq+zOb8nyjq0dIMTwKvGtncgUjT
UYCgltsUTKVo4SW+h0LkFb4e9Oxlo+wdDgMTQcY5b3Ui+IzQrZzb5c+3JwLN
D9ss6hBTVAgiQnlns/S4nhFcuCJPVoJb5mIzox+kr/qfZWgmRYUBnsRmQctH
w2PWsRWMlQvyJ18lFSaq5VjhNpoJdWLhRBddl9uS0WCeM+ataMAQaqL558d6
YgcHC19l4w+URwtGEEnJWc1afyuGbntf838rqBtqehk5VxA65KeUyDwBnBUb
rdVVOv8TdklMdrRRDaINPRNVb3VBtPH6F5QREOQQSduLWM7XqYUDSYzCzobB
HT55ZaGfCQTmw/ECdO14yUFKaBOkJQtro391XQFVrnhNqVQt9uN9Uu+c1Mi5
qAhc4KYpuRBhJbGnFuAuGQyqoQz74C9JomDYH/m8dqN5Y64Q2d8PUWrkRd76
D+CgbyWHjmMptkFxym/hJIvW03pen+zC6KKAj/mZCjrMH7z0+KjcKDfbNDVc
tiEHXng9GJWJ4cxCZsNlOz/1NrIY1E+VqzPXDTpD7mCLSooHAewVgYodDHRp
0z02fqeS1eSo3LGpq2u33hHD19rXTy8N0Yt5I50o+R6tXfRiEZiwQjoQJrDi
yxNniuuWZe3KZHoqrTHknjT83SutCCrcVkwX2IYh6ybG799q+Xhr1AH53d+X
M4lqwCrWlcu/3Fqph9F0MXACZypAmbs7qMenV+aSscWMGxU5q1Mh0D/OrNta
SE3c9pSDgGGJkrNUmQ4ijiAdmG/BMxRSfew4QMnrvaPhmVo89piAOMmm0CZH
KsxKMfDzfQCpEMc6wqGdpLtBGzFlOVg5HLQRpsDMpDpBDLQ/20Iq6VYEb74O
PFyukp0+r5jsh1RkPy9aSJEs4S9AO+uAbzR1mq+VmbAdyJD8WU+RXBkjnrmC
MPF2WtHDWbu03ey/JC/Pd8rSLpOwvezm9yAG9pWRhQ9OWDj2R3KvJybKbrcs
ZjRE9Ta7xPEF8JIlNR2XvE1rszC4EYXcNGsKnndnd+G+xqjm9VPMgzBQZKhH
a6PK9oplsFWb7gYp+JidBBFiOTCYffqcS4bz7iDqzqFewC8ealGLMOQKEXuY
/yNcTK5sGidhQ8Sxb/OJCXIZUhF4IfnMvwmT706gy4aTT5YKQUXhrUCz7JB+
j3XH9DbqakVcgtMjMh9zAh6dxPPI+yxFTH7zU/SneJ2rcwvEJpYquMVeg8Tz
w50tJDaecAC0XJGFJGZ13X2TlyncEj4ZckJ6KmmCUI06M3kVnaBPZYiMCmX5
P0xtfyFzXLNc/UH+t0+eG3p41zkOCp+dhAbbhj2+uaNlOZf3EfDk+hady4Az
Q0qp8cZDIasfm8v8PoSMvHzEVlzVmjGzscAxk4AGI+RscbsQQn3AuvySgDO/
+IwWHx+UXVyD9+bYvR0rT/vYt55p66WY/lfjw8y0IjwXOSuSsu+fR6JnqBi4
RK1CTHEtRwJr1ifygGV9r0Apd0+baYdrNw2IN5/StilPuxBL3qpRfU/hfsvh
t8R5m+kSgCcVYJPOd/ax5ROekzbEkv6tflqoJuLGzwghnFCGpKdkYZpys7QD
l7wMwGq3gIfI1nq4YPDySoPXFHJTJknNcWCIURN6AP8fBwVOggsph4NkxWi1
Jwotm9nqm9HRCZZPSDWXT2pk4BAde7bYE/GT5JvTkx5sIJw/qcbgg5KeFBKT
rTpFeRVlFaUpWs6N40HkmalLOHTvLyteX2oWpV5xwH9zdU/5VY3aL1wyIzHX
NIeJ/4khcigCRmjsHYo/9zUU+vswbxLunJIVP6GrVkgZYQWuzPjHVigHp/kS
iEykDb9SgBRzQrEhz+rJgEfxAzekLayfo7cAHxoiiR+gzM+JW0/qkKX5QC5P
6iRuFOmCWn01ZYV+r8TqSapr03QEXR3iQ4rrtX2wiwi5LhVouyC0KJI0+NqU
tXAlefxN2PHV4hbzl0XWCXbq77D4qM+Bs4oCQm308oi70djrTNgklFcL8wq8
DiAkff1oITqke/PWGwYxHSk/kx4SFgrmcltpNiVGDPep5QDrOGwskcBXkmrl
oJE8yt4mZ2f3ovPvLvdilh1YAQqdaUsrxyUwc7sp5sDS7FU5opQaMS5STLNT
MUWAMzxHgPwUmLIgmZzN5PWoWDVPAZ+8DMOUdfpGVUJfvrYtNhp0l4xiqcUB
XRWa9TsNrYhwsRCeKemzWqV0ZnjCSEhTgiray49Qqxy833GchsP7NZi9niB2
oWA/Pw10W72rYV1fCzsNHH+JwfzU267IKh/9jX8P2kKax6YBJJ7LexnxmIDQ
8VLLHY3nObdm1L02U2QJJzawvOt9i0EBbcWcLgq4kssc5BGdtiBiS3EypPrC
aRt7WG7WYBihc9I4Jegn3vtrmffHKKKk9BcuqXUgPMIkJgN9JesliAPG994S
Dx4uJIkidhMZCXNv1btBa8NeR55HeM1Vlv9XmZkSFZcTmelegfRvkFoCeWfS
iqTMD//WI2/LK+3+SXHhaiM2O7oB1jPHtmItWJeiI7FEsKZTCz+mEVv8QZU+
y3Zi4cvrIt1m4wnZXo70aB0L98LBaaLYzDUEGKR41utizMcaOwBuY3YlkeDT
cQXVtei6iwl9NSEpX5qzZVgG4rCvOsRgStlqDc2Xvn5X7h77r2lQMtQPWyKa
Mdle3rt1JZOGGlhmoZwIrVdivj+sea+4cnrH1yLUJaBARwcJdaojtwqdueGn
7dCr4l15/zXCoGvDMCeyl6IjmePuIHX8RpyqylGci6TveHT8xdluyW2dHll+
3dcSLlxORNCHtEX7FnUtKSOW364JUZEJ+niybICTSQuhBpwx+mHoMF63SxnF
I5GH1kmGRIK06WRsvCYbCLO3GbG54cWQke+SdSYRZtjCfonCOzODW190noMr
zypwd3L6B3OwtryU5wuTnueL6q52wvjgTSdRpYH7ZtPBueBGGCQwQ2dspDrN
FbXtG6xRBI9RFu8Y9syFBITb3TcSuIY7TmPPUcNMvagT49SObu9l7QRfvSxu
J9OF/OdbsVWS5tpRUmWIeO8PYZcO9kYLXzQyT/QRGWyDv9kk6aHNdQZ3YBpc
ipcDTFvwKSes0ARPErfv8y/68eCw85Um/7kwZpMuBPsuDVoo+Mw18h7COPi0
LDziq8O2NVY+0NuTJU2uUcS33EqfwSeWI7cBV8Bfv5geZ6duM/QnOD5pT9s1
fBb200cfTI6LQBG36FtZxgCreUtG7sKxrKuGbtOIO5exvPFG8SehWEvkU2if
rX+m97sVtcCpuTFkkfG4MyEif5rGmSjYTfPYWD7hDG5++mQvxs4brxVBJmug
hEHPv847GCPe5M33OnmXBAsgKZM+/l9sYBwvcR+gjKKbKbF/f3fFY5UXpTMn
HvKXfZZpqZ/607upZuvIIwlYSkpcEoi5snW6+vNlAt77IfIKlgGprxHAZbwI
t4r/scukJMzLy3OZ9jY8zQKQe6cCaUP53W9mMXPDi8drsV+7RhwkIqmE3WIM
42tSgTvM6l87d0y47cMc5xlvybNrcUIVTsz+t/YrsCwByYzXMq0xYTQU1QrT
RbGQbon8NORQP8/QcCuJKUIsecIPgmiYq56gRcQnMKNqgw1dW3sEbL9egHE7
I+ri8D/B0fxIVrUUQP6XTX6eKSLGqX2OnnAPSf+yMEFjbG+VsJQk95i/ywxF
NGgeDRiOBe3NBDg5x5hcoNHVafpZMulXgnHTOjkuqTyJpGhsezy793i4V1S+
oocjy4c2m7C6Kn/n/xy7dHWgCqQ2z5XshMS1uh6tMQFVBkWPmtvLD4NqXokU
PcNO1tOti83dnRuBnFgOofaB1WSmsqGFmoN2x9E7zYKfsR75RHQRmJ2ULi7r
Rj+YdXkRFnOTL1Jaf9uAvhT1rZiILzrBkvoVDS1AEAXHRuL0/THVZMgaBm0Q
DSPwROGOsnmWmqdrkUc8ZsOqLr07v0Je63aV44ZQrl0MAVRNV18WWAITC6Ym
b8mYUHoOENNGK4VeaVka8sNYMSw22XCOIP9KvclevkG+EdQt+Qlp4Qu5+SgZ
mkBrKiYgWWyAnrbjl1SvkbInGJ7momIvG7iizzE+r5EgLMBhQ00/mFMqtLZc
r0gUlVzz/zYNFbhe/uUX+vbm63lYu9BjA9464oJB8dHcQ9q9Lv0CaeKQpz2o
LQYnkr211XVLr9fzCkeJ02wBdaw4HSqqeZCuTNCVdthFP/nMFaRHUk5Bf0v1
UC9zXDpb3auZ8LxOCN50tYOf4Gh8hXujJ0fHTtviVzgwS6VJDogldm1Mr5Dk
nPqoLZr47lXBkLSVEnfOi2GRwO6IstkY0tAj/BfhNdv9zSmefnDM+mUEosrU
bhYhH8niNZqHLbekn5PTJO2ZPBUmLyrJ8k6Gyb45MAFBvu4TWi82zDj4RZYY
nQN57ASiqIKF7Dm8VPLqqSNspYUY2w1yotOmuwkROKf3H7YvF72R/FiKwBuO
9aHbp9p09rsFxTVgO/Q/OvMdtQQImhhuMLxHMWhQ7T/rPJIuuWsNAw/HPQe0
JztYuFLp+JGcgWRtbMgJt4P2aoHd2r8QO6dGqwAOyJHQSzVYupotvFhSE1xf
yQTlZOwaagu5oG74VtcTjgTiIuLwf8Q7uNiA6HTxc9Tk0VPHayi+Wg31SZp6
eXp0LYSAqLFrzlcagOgKBtmUYpWhdKnzVpprLIfAgeHD15J14RBQgyS1yX2X
teqHN0nby2grzKNh4cmNUraBVI2m36PVFwLOfRtqfX/jYDnvMaX6OneMEqDb
K837nIV1KaXoyyDtecL6MKqT10TShVli2CLsDCstvspZILt6iEkCUaNmurT5
NvQcTpIdBczA2qQmiddWq4Y3WusNhzWUL0J/tcYB3bMg4UpiwCcqwYtDVvG6
M92TWxYq+Bj/o//jEeR6icswyA5uTaoRIwFwTRPT+qhk1q7u1AI0nCm4HiIJ
Eax5q7QFSOpT6G0HUWj7R1Em7PmPZIXKGbAsUYU65Z+FbFJbr7sv+XFiBhs1
+sapr852DHNKXJn4mIVnc2S+oHjmU43ARJORLAcqi5lALa13qAgdj/HtdyBP
Euoxvvlk9RwbuFnucFznjWhSuriF0v8wrITt1Pa2p+8CWHTHjarXe97hOA5x
f0/ANIsrfxHABnUUF0duI/Mstzt/xrebK0FSvLJ2NpTq9CcoN9eFJkGKMWIM
iXu7uEnlP0JwjZ0VnOxX99SX/GsJfKc+AH2VDFyOLrq06lql0GFiChv+oTpw
jwK+JyfADYf3LRf++oar6IF5dgvHdV3yYG9/5uvBF41x+EFts9K/e+xJ/sM0
TPpyoIlLcmdVzH7+7cj47KOT88LdgdCm1H6+evxoctIvbi2Zbp90frw80DlU
ICVRx6BaGrp+Z4FowTLbaI49XDVAbmjAFzWxi+Q3mhlWVoY+bsN0indSrl3v
HN0UCfqukqOTeD/FHjygAIZf23o8ahZRLP1dficK69ivzFqkh2qjvZ9NLkJg
jeXiLCTyNdPFSX6xSv/tWriWTgo7YiSTeSesNO601xWLKWToOdctvrj9FxBL
W4k8sNQFlbXdGtgR0P0CY+wVmiDUK66f01lFpS4k3woJvXmzaTFe3RHS2y7N
lYfx+QLFdexxYIuTZbvazGwOIpGgmSAvrDrLEpO7+uD9/3L33t05Ex2Op6bN
VZ/OUiu/TnwKPTX367dv/p6zreWtoBjlYQPGhWzeFiRPSagkRLVtytnP3VEP
wZZXXzyeKGd5TyBjOLM92ZemM7FGh/jQ9YeIUXmKQFU7MiYec6CJj7UUqlrp
FxkuhFBm4Kw1tHeGQO/6drAMY5vb7zScBTzotbldKMUnV41PQ6x99g1xEy8f
3VECYWqkIXu//Qit14Wry99qj9Eu+IA2L+evCtPmiI6YQVfuBdRAOmEnxm7d
M+0zeNl36TKhdfwJlJFIIRWSyH5jfZZwBUyhL3vveEDoNJBzZegyyWshp7L7
DPgc5sXDHTr2tZmKgD06Pkj8+NEXG2YgH2IB8n1Box0qrmwnqa/5QpkojZk+
nEsl87cjzesue7RTqArWuBepMF67PGAid2Ga8E8iBesmz3X7ZbWc9HYRh/6T
c5JosMHDO3FDUg/rlYlp/epHQgC2xsOY5BuyhmIpd/zWgQZDowqskCjloKpo
/y2KeS9GFmq5mUIPCainPiEWNz7p2yBZA46hzQl66aXZBqw7QUeMMCcfUdRH
DQoJDzrhFfBI+WNbeVELgG7JnVgez5HcvvfIEq47DjcUsOCsTdYSwY4555qk
9gR/0T6fXsW913IUMkMIz0tfxySEgMb5p9NL/d800rqb0zN9v0lB3JbGQZia
3JiG/2vjipSUCtrWQtkn6Cx1nU5ARs5onperT1I9lw55hfc8xY5sAxrHy0g1
dtNciEgzRV5o+VZTLaO30AMbM3XKhPDrFZPPvJjddMaud9SM7aTMsXGYf25A
V6w0i9zbrT7FrEgf0JTW6gL/PdlcAN531sJHsBbHn76SwQsfXeRKfj7eWu5c
mdZMIfBnhI68qdeUWcEiTqKb1Bkh/VcKeLmQQJ099c6cwF+ZzgLsEISZ/GS7
N6rneZE8x8FqPDElm5DtbRBOOic0sIDV+e+WpGP4SzdIjbbnR9TlwsFbXW16
oQJUGPpw64fM0xHGwyJgdRKXOt7WgP+LCUMboWuqfOFEIFYw1z0hqfiYdLHw
DpwhNgrOp36dA9uk9nTOcam0r/O1k52YJPh84FL7Pi3IgZLmo157a/DR5UIt
pBICHpzfc18uVPqaQbicwXW1sJ1jwu6hAj7TU7r/9rE36VZ94+db0D9GF1YD
KEdM3z4jPbs4uUrnnmeedK3l779BN9RDR+e0HmGTNQu/63wL3Rzhi1UpOvtz
ocnL6rLmXksX8dVEnaVUzQvHq68X8YHrIqgVvc8FJWG2kxysJPVwHSl6ds0H
2R0247dNzgfuzgbqJoaNAF0zdc5QdFfbqJVpSgahtqXpDDPSOJJXAdYr6dEv
NhApVc7aRO+vyBHcCvKZBearPnuBHS2Br9Ug0mbW13zbytQ7y0QNP9NfFazb
I3rljAFM8DNivNlrXGdtVQGtn5DAJ9cyZHWp6slA5Pq30fhPjGaCKusnDZsh
TJfXzV5T/fM6x06IWurx1vygqFpLdqQHprWGqmFM+rwulCJtb6N1vd7mkkg3
o51skd1r4SDABtxhgve8yIjasiuJXBJT36JMuP4rHi6zQz9UTTDJK67lihFH
GVrSmpZnTH++3W7bCvJy7Vmjill5MvvUqUe83MSZl+XSNrBlJKzXalZNVNlr
7bY/GTfoeZ4yz1nytEx8mA5ZvUEnnvjLKvEu/Ov/D7QcAoc9XSG96G6BjrwX
pcxQI4vYER22y2aNq64RLm7r0GLw5dRCT49h86+wBlGIUVDzOOKAhq9M4846
x5vM7zSLDOBzWjEmQY8GvxKcxBo/GIc/gQ4FWRr/180/v4kAX+ARu1YHiqgp
if5EBhwLU07zPC23ryzpIRBkqjM6c7gqJucvOQ59z2h9u/YMxogS2qQpV+gO
/Y5++6gzsJvOYtFzZtU4xPfV7tl/dOac9lXuyVLRCcsC/ChHHs2WZUB+apVX
fQdVgy9/DXMuDqPtpKCDMUU0EPaO/AloEwX2ncKqLs2LgzwJyBsAjs2K3sCE
Hm02w9N8ROi3SjMo6F/AOXaU18CKO62jDHZTCTqSVfY3kb7ZWiWyD3whhOKO
wlajknuVrgZdXGd9NUMVeYYzs4+geTg+f8augGgBpI5U6HRcY6R6t3MgIW2p
XsK4xYyIdNxIFICI0P+GjYOxkrcdXxBenzV3yWbMswBZsidR/dquhVjv3EyK
AUWFlV6m5qynXMK+892aGlooYyhu8X9ZrigSfduIdB3gm7in48/y9U1k+bS5
yTQUSbnBnOhYtXEqX+soaQp7s6xGgiNNJQpKdXxstEebIMP2/pvoA+rFuuLz
lX5fYeZ9VR6y/vOYRh3AGny7M/yJfDUUCHQNUaJk1TGDAghaN70aG3615Jar
hrPF9IKxo6K70uS3/9a7zG/tZ8rjZ4wDFbdyCzId4ooGRU+FyG6gWC9pp/bQ
U/jgZ0RRJu4K2SMKm/ydGcNGTuRrt0PQf+cUEZjB40SC3B9q4H7pnXGIc/aT
SCNihTyphBR/PCsozYs7EgOUghXUZXbdEaTbZecuTXkJuXEpU38MACBlHn3i
m/C8iQHiJ4dv5nKo5wafymYJSg/FN1HebXAxJfQtE8FzsZB1JBlxk5A4LpEe
h1HEZb9howVG6O8LjKdfiebg5zczmMieCZV0TjGLmJa2OF7E8mzPIc/hSaeM
rN0HvyCnAK2XlVkkqaST6PmNfSqEp00M7MWr4OnfOeoR6GlEmTnQNxYRCJ2d
g35sMv5hhFPA8RiqP6CXXe1htCohXQnDCKtv3xNco6B7ufoNqeUp04ZS5ir3
B4Pbpv4CpCY4TbrBzgvxmeOXCPGg7fUcTEKt38Fqc31Wejlb7TJAbmVuTZwT
d1DUE1T0BmqoXIS0nu70lNVGwHk65ry+5hUp+lV/5RKewJvqu527yYUAFXkS
NyNW1IHkNCNLHa0oS2aZlX5aAZ8KG51W4wDJNtlnYm2FwAkj7YXdGm6R2mH5
WJld1+CEYnGdDk1yAX5PD6SiOzkE/sYg/xrYp1mPZPAPhDAAi7SUlNcHUWb/
TReP9Smx741CwWqL+R1YrnBkUqTK+hRlb1SmJZDCdDeJzi+S6g3MpmWEZHxp
iq0mLG9FB0Zl6IqBzT4t1A9XfKZIL9BP7eb7dZRDDJC9e8GYpzv9VsJOGcN7
/l06q5W5QmcJ7xpep7XqL2HgRuhzISmCrk8MAC3hbjN8XJefJe8Pyth3RYeC
dAmf7OitSwpHVOom7OJqpgG7NamDAqIopjGMpWV4unrBMtQCg+XovnUOFvFk
SIDxDfOuUG24D1GLluqyRwkE1pQCmJJC96dvmOO2utL70hNIruy6Eu6MMiG0
IZNKnKe36zNYgM283ubVPcjFi6+xb7aOBObtBLpL9Ctv5hLTRfHVCH+Nl8+b
KcMdWyp5UDALuJ5yL+VB2cgZAeI5vm/6wxVLLI5C5FISt5XKt1mnjvb2QmDQ
7sx0dulK4Ew5vNCjZWI6jyABM9PC+uTQnCdQ/Tz6IR7eAvx/jmWIVa6gDC8f
wCczyPH23jjKCOywYX/Usw5sSh83j4tNf+2cGfmKmy0b2z53qDcjSw8rk+Pg
CH9cjNLuD1LwJ4W4jN6zFnZa+udIIfbPxAlycU2uSX3Y+dxSmQL5NbAk+7Yg
Pho6rW8BkH16GSbsXp8igaiUxpGea2Kw1nIkoauLhbaGTbIl/Ho7t8oArQSw
78YppERm0sDH5xyPUZbsd+K1/du7r4RT6ELOwGTHTr5VaDzVPpCuDx3+Wcrv
EW4URXFujPQ5nTYHLrIeiEa9TaxWLC42GGCGltkqpbc8RbatApix8iaGKhfV
kjWPenf7n5eMS+kkXpLTKH4yPowZXoaQnXX7rglWVzOhLdjQyCHLmHY9Udnm
qq5liC4NPRCqSwcHkjuruMDLN+zjkhsl02PbMyvSdtJ9n4H7E2lHASKD1Yo9
NeUgbYDpIGQ+Q5IIr4DNJaZzG0lBGy3r9xQ8ATiCr2Sm+5XpqFtsppfhINIB
mNRabRgYOksEF16BdRodwIh36oBHEMPgkiVgLbhzHGoLSVDo7qmRY+3Uz1rS
MzaA5giTrQ0Id8V2hHFBCY4cCde4/gMHGx8b9X+hPj7NDzCfJhsBm1c9CxLI
x3fJK6SbdNzSMlTOTD1bCVHvBXsn/+q4NEOJ1Vpg0APaY6MzuzPqaH90eiFL
rs0dm084EGDEkBxISORUO6sXptEocCBWht9KSKPBqObxcr4SqLLMFMrCVL3Z
o8Afo8HTUZTNQehVOxwkdjmSImBuZHfczJuFYbDxLzAu1RmlhuOBeqM17ANy
h9XuIGmLYUtw+ZSV7jc10EAPSMOmHdSG3dYf7V8azv15VMT/r0k1oNDx/n4f
qtjSxX/IFPDvdZa3U0IF/YS6JmSCCOIPFivbERc2FAu5emfPfB+w3w5UeHEg
9LLXsMJad9hwgPkT0ct6+uLjq9kLKqHDTQjDMq68uoFSCy3RLUvT/qaCxpSy
65CzOSAPHyPzJKDPEOnJm3EgK45hD35rk0yt52zMyKRBdRRsUwHEEhaL8Bv8
CYr/7mk4MJJnv2KeRvBtdCs5q6GyM+ZzZLij+GztVgo78ONJ2SHYV+SZN7Dy
p+LZdH/ttpTgNMxoaav1vSUVRI8k61gekdDZBhZ+Ep/kK7rrlvkUDIsZTzzV
cKNCUM6zAk1BDkwogbpgEv8NJZYcM8MbInnhCpVG/BShtzBtE8R8RfCqnIFW
tc9cvxYJ2fKTbdvFocEK5BzcSZaeochjz/UCwz8AF+6oc7RDmem92E2nlTLe
R1NrYuzbMpWH5eoj3985jaTXyZ7N1Rtq8G98a8sTXIvBmuypBQYMIcY5HV/w
fDyASa63AoNg2Usu3F2EIGZzzlKSOX6MbYSMpsU3p7Z8sLKAi/BL0lEG/2m8
+WM7qNC0echord3K95K+upN4TMh8WAUWURYNqs3eVm3R0ao2v7ZvApycbsZ1
/yhH3JuUfEEuPnqC4oIYNdXtDd4DmFHEjF5sR35ahRUBsfwShUjtkQBj4X3b
ouSUMxtVTATZhxCXRuRTuGBj6oRThKIjjx6LIkFnprMfLHqXWUkycnzsAKui
8j4Ko+YNEAyFSknNsXEVRzzhQ9/pRCOg/b5LUVVJke9mFsVl+b/nEXkAYUQy
t0pvX/GLIQw83rJ8kA/A9QTIUtL2ku29quaYW4C7i8nR6Ugoh0+ww1cI/q0Q
fslUWviG4emyDO0R4ZxTzpQcwR/030TJ6GO6gbwcnJGT/bCH8uJX53ZBcEEH
figXgfYy53A9dFOWBFQmUZypcCZg7Mf93gqC+lbNMEOFzEXa+TxlmpLQM2U2
HmDSrjOW5qXcpH48w4E6ozfJxkPAdGcqrse4Ef6G1j3EfHGpl6igXS+7HDUD
YvQiPwppo0Y9N9i5gQaqAAHuKE3Kldaq1omNauWFKVDWXosEy6fh1l8qQeZc
/ayjIUMvanSe2mZ1AiELFcEXh7J9XTb8lmcOVp0yj2B5SNNBHlIFNb/DmlcG
BPGle4HCjeflqOJKT43lSo9h3ivZz4iMR6UpxB3MavqDGmHi74EYqxpS++1w
ZHdA7H2Wk2kOXd/oEcstg4fxb9n4EjjNnZKDVNqIrROpl+X9kzaswE+vvXVA
zQqr3oLLP3USQBS6IyKAgI7HOUu2Yvwpzu0Vs7XQx9Fm44+OY5ca1A24nvB7
REd9ztCKuCApIWoN+XHgkEpV9S+V8kowzJ7stV3CrLk9H2eSVg10oVkU2Czd
CqhcaTGz2A911hr53r+jzxuT65BUpFWw+eorXy0cvU5HtW+QYgiIH29OpYJB
dLL8mWFKZZBsdRTaSbw3Jt3teLpsjdUFDzWPscvqmIB05g1rnThm1AWlv6KY
vA029+cMwCHHbbxadEpjal5SLsQtYu0d3gGlJFUuD6prVhsIHaGNTHFwQiZj
b2VX/0jHrNnWxIgiUi9bpeh1Pukw6MgqMLLV9msXD0R1rV8d8h7reZ4yVN+g
RxhbZc1fFtnbomrkP6AQGNENqv3lcbO2XZQ+Q2v6AyGALsB6/ZNKiPFGc/ek
pnbVLwYYPI79xiOsfXnes2cQIHK5ruS+wRIn4X8vC9ENLxqcCr8l5zPWr3pf
pvmr//rfRZRvJaykaplXXFNtycUM+EBR9HMdmeqhjqesyje/OUuFiJnzY1vu
+AUpCl3eK/ZpniiRvTtgq7B+e65qeKu4IKXmPxs1uqp0qYUeV7JLb2SurXmW
RwjsrQA+WvQTkvA3iNTekQQNtrJeAp6UdW1+Ln0FLi0ieHq5xPrVu8tSeDly
ccWIBKdXlL0HwzPubpoyjfv7ZJ75Qzyd330AaBlQLVrfpNhsYxY32lbIkUgq
T4V2aBm4OB6bt4NvtVDSP3+R8KFh09WnzqIO0dHUjfEbLFzLixdN8eYSKbXC
rkuprZgt9NJr8SA1rrkWAgHUNmirWQcmS9JspR9jkWiQAidh+sSsOpO6rYvX
0NpuHfYzuanB3RyT6xLaGKd0Q6W5c3vTy11PM0t7T0W6WfNc0Rjeddqlxnnn
tqM+XBtUjrWxIMpFwJqlO3l51utrwBlRKj9Itm8wl8ug/dOuLql6m6ZRAiiE
89DXI4lCMpwUxXW96NO/sHWaK58+P1g6uRiwOkHj1h7NJBMMxl8cshizun/J
VuxQNNRlbb9+A2mTcZ2TjD5ZC8j99yARIwKTIjeFSkQ/K4dkYFFFrS3U0KXK
88+ZqSPXQw/rr3G60Sg0mdD11wZv1FhvEAScPHd8o5BV5d2TqTD8np98EgCc
fIGYm60zDDshWHepOk4daAjQg4NL5Mup63ldcD9pisvNGgx30vOcIAMyDKul
xHGUSBQeIBHlqYavrFeR1QEi1SOSkA7FHSnxv1ciaAecUhpmRXMZqmEoF/q7
+wyY4F6TTfXkMKynTmaJrbnnv5N8lPlbf8W3UfHZqOoyH+ndcJ21NBn8OjCF
/CWEr5g+WmVvQwjvN83hFMVzA8XrUstiKsPeTnUHsV9naB1/fqgbRpgsTzbT
QLhVSo4GwkKXjr0eiUPIU8S/7IP9ZskLSzR8QFoHs2gMkQQF/b1J70VNAHZF
jD5jnWSzt2z3RcnGh9eWZhFtJ9xn/VS/ao3QPC2jcLo4QW59oAQ43Nr8qsN9
jVJdDOEXXnJI4MKtRgZ3JHPM6GL50uREkpbRd3Wi8foj2SvBoEMYfk08e5wO
naRKsCjInj68jJns21UAZPC8D5xGovY8bbsAimx8TSSh/JKw53FtpxEu7NCf
3Ys74MvIH01EkY4wKpYro3UykQ/DS7Wd7wKNA+bDMhZyGf3JXwDpUbsv+RAe
2BTehQ6uMxG1YI6NfO11sRdUBHt8ZpBzufjF0cicFsIy35YcUqkEDhoSftrP
cHLebzbvLiqccNg+KwayBnNMr16VoCWGjVo8jAjFoKTkCBWOBcTOa3j+AtlV
6EspFkvNVzZZ9ZvNsYQ/ELKGxhLxWjOh2WUEXA68sGsNPjHseXHq4nN/u2gt
UQcDihzJLYzudIEy0xQhgR44OepuzHR+YelUZJ9AVBgZ2ShAZbH7kZ5P7QSX
g7ndrYkP7hLBAtNGLmhyShe3b5xzIVJ9GK5LgOfsB7PpCXGiAVRrzXmHzUDP
aklUeT58DCMYKD1V2ny9Z4KkNheQHY179BP7yUclmksuXfAajCw8Tec9aJLW
3mY9oedWrcS9z5tjGlNBVybmmodpJq1ckVR2fKIkyOjFJ40AAxbAkWo+EWuK
eKm3AtpTykSMbcDUntnp9Hf5UNNDDy1YcN0s8MitewhEU8MmLrTsXPnFu4wO
yPDixQ6Hu6x6HYt1CAmegryQEx0NdwJ5eKSr0EdVrLrFXK5BINwRSvr9Fwb0
rjSXlAfpEQEASU+y+28i2a0xFbvGc9voU4wQgTjBNZVHBFXh6mdxO0RJis9L
xIwfNsH1xcztdx4Pps51K9hITIxKMSLnj6kfV9JBslytnUnS+U2zEQOLC1nx
lUS83710e2ZlzGYWnxs8SrNaXdUPbUBugmYpWxkb60GwJIs45IHZwOFLKKTr
Lf7iZCSkvx/khe4SmIL0vbfiMuA1wH76P5q6r4R0LtquYT03szL9ZMVfjC13
yh/IebV1/Hyc4vt5VvC1AO3Ttte2vtSQVCTZLTAteD/nqWFlAQlqRNlFttXZ
7qJJNbwNPipc18kACH+Mk7pfskemMC89tcRaz+UNQU1bgmJhaoTmYnPcHI3p
5g7OpfZTgVaNnPE0gnudMKw3GViizoZ2pz1Z8kHCN9CzXTGvg8LtwPOVgi4j
wHtCIntHoodFIoZzoQx6vTs8/eaBm2wUZXxTadyhhNJOj8ci1f2rwjnvLuGA
ADD5mXcVEwlQ/e7hz9atx56pFtXJonNYYxlrSHyhYF8L9/Kc+DQzaupAZnom
P0DdOizSDOYEdsE5DAFu5TnTYdihI9b08Sn1u1f/u52q8O60TOIKy6ypfn6V
G0QNYUvZFq2FBxIO69NnmGf0wxM7wD6f2udXBdgxf5Hdgavay53t3gpq4uih
NQEAP67vxo6wje0IgLV3+x4FgRgLlur+kEPBZuQ7+VyhGeSzFM+jE/8k2qwt
9yDwZL4U3ip+QkCek71RsYGnjomkca/iUdEL8i+Mt7tOPB2nYoU+xh3CwlTh
kAbJUtWbSoxUaBKDWrqFsR21SbwLE9elNG7X3NjEymUYERN7YsB59Kf8a1RD
96OmOin6vpnT+jR6I5kl+Qn6XeqAbZJJTcrI/e6+Thlo2H3psC75vXG1ZJZw
x2nywR45h82lfvHmHc7iy/jlFbQFB9RfMQX+gaBKeZiLzZqfMEaon/ezJTPp
08n4IAzslb8bqM3uXJBlr+YeMW8Hpp6QCp8fsHB/uWp0knVTaPfrF6uPeQxX
/3IMDZyrM6m51KNSwaEucf+sDvr6xm7LIZjXBMd/FJTcocSa0p9gdU56Te9E
3YEaFUqR609ANXBwsSpuw87hdm4j+csvBA3Nd/QE/tt4cUG4LQ7MIX7QaQ+T
hWbN5mCw/VH7Ft/ZUzrNQZS/MUe6LowBKS0eWnvsVIqTgExUzT4dpphNGepd
xEe5p3jEAh0jN0VFhDJP3keaM0PLMNCoFNxaWtrRKc0nzdOO57aTTpJWj3HQ
7sXtWFRJnlYNaaprwaW5dsiH7BGdHG0I+nqLUZXlcbCcisCMrDJJZLO0Tltb
o0GSJRCuCXW0lVS24FnnKjjU//g9MWRPHzBf0lSe0I01aduuMEQfndv/q8z1
7RlRMbSS0Lehvn/Z5P8IkPVcTEnNFwia5VxZglcbg3mntRc4wHSCIWr5lGI+
H1NDkuVezYaxZy7SlYnQ5odSHhVZBS1yc06nZb0hqIsWnaUb0KBfcm+RTxkw
QGaMwYS8lWjUivVtthrJnwTxlnpPQJLkPg3ah5hI/M/A5Np4kvjop3hJabzR
cO/w6eqy+rmgZElgrDpOjGQJ220cJDIYyJ/M/lgf6UI81lBTU9etSpDcPqNG
BPCmpYEZsuVgtudSNAnLNUx7AMwHZwQm157QNJcU4YsTq1A5f1BJdf15Bsh1
5f0AYFq4a0pK/DmNq/yr31JwXEKgXWCupbHwZh9aNWgBXagVnxzjAOfPmR6c
1/ogmUJzLfxhzikkQojlIFvtjNBSoWfk1dGVdp0TM8VQSZCV1i2MaxvOboGS
FLOianpdtUYCQgVtSp16d5M6ZHkMWsXSUAEntCQi6PX1k/BaooOvls+UWLJA
nHkO/VmDczCimkA7ixbl7xECgYNAtLYFag9dbTmfK+TNBkEPpfVZOXL5OAz7
NYIFJ5TeSkOrwAHaygRZGBVm/pHX/IQtU3zRCqDhWQqqFiXIcRiQbCInpcJY
8wwo9BFH0jH8eNTEPCucu1v5wtAIGi4xcJn1t0TCAw5zLIy2I2BWGyshOThE
4kTUBxreZ+1qy8yJbAmmUvjPgneww2g6N17hdROEG64620KfCm87DHcN/VTq
pZrJF1Ts5abJe+I3L6fZTYUpfFjLNRGyCH+y2Qr3WoNYKfFhTOO4N7M6ujMl
SsIIdSN+LpARtD6cRFrKpa1QRkRkm3Gt/olv6m5Ex9ow+BIBan5Jwix1Zydi
4RRFMNUeBTBJ4/91QlcBqMRgiJ2V4fAb8UVXPIM09/hPUIZskD2W0cPWH91Y
0wwJWnyhmFlCcXBN6YM32x5Mpav+OzaA55rTULGWzvw3pRr8eRL/eyn0XbWd
j6V0r2C5EuTaEe8730eb8pVCInaE2hMZRFKDeNc5DocxtQioaBuEcCf5WPQP
JtUUkxucbLZUm5t8k/hpAab4yLSYh3RzsZcFJsaVLtzvMWJyBRcRvBipQg9H
09oebhc7yGbPv9LVL3BNHfCOHNCSvk5CIWM7M9jl71qxnkeEZ4deKAWpOc/S
tcSp/FLp1y2CyZNFbDvsMVc7xVh1N8tC1c896mzAGbJhXOzM7NznIGcOYoIv
4/Gjm+QfJUHjnx1UdqdUnJNzM+KZAC9sNwcncXGN5yichKL3lJZfgj7UZqSm
yKX2BAN4wB1kAUAyEWspt5z+J4/1ISII1ULqZ9YwVkow2VtoVp0VB3NR1G2A
n/lV/o4Kezz/b+kHyRKTwMqN88ChyZmMPgWSdYTuUFyIuqquFjsW1EezVbxd
WhuXC/2jduqaPPVRn0cCpERe0tYiVLy3pSt58BNHPO1OTvmo9gaFX8iIl4r9
zuAlK+3y2YtaluFzSTV4VXXEB99IbHd+ou5TBq+3AY9iE5o/dilNvCMFlEdb
B8/0POxRssdG1T/TjoYoCo+5DVVa2PtNx6r+Rs5pEIPbAppmeMgQPFsu9q40
ro5fFAlk07N11E/fyrIdnX4AhZbDuYr4BC3mXYo2Ey+uYxBHmD8s1Y2FfGPB
hgdcI/c28DHc1s9Nj6wOAHUsAAO8rnjk+9PKLyrIT+Y9t1ch/NCb+UWu4yNn
0bgjLWQyvMLPlUZLGELNma2tCPssZKF+Bf87sLRFDMu5Ih4mawJ6310Msyjr
t18bxdmNxmXxB0ojhe/aoTl6675YtYwiNRYv/LYiMZfbYdyFpFhLoS+DS1cU
lRGaYFgBknGV+pQQFN+HhU3Hs3DmMlEYp/2gUk/rIW8YZ76RTff/eIcvpU5s
tWCmJVZvMZRoR5RtFhkHLPdLTF5cefLZoBJ8SEc0/ps+4ukCVM8YHpWKrDVa
wil/Urs7cxGjtOo0VwTadQ+ekJF1+ANC7gkSPohR9qxU1WgVUENzawmAQ0FV
Pf+FfRfAxkBGcziV0jW8KCvJkWYHsFGoqrtbKlHJf2HVJjI47blXP/bRgXEW
yDrUhVaS2KzcsJnLZze7q1D1vYbTizbVMeO+5E5M1WDTsRJgmMuOTb9+0gYF
YtLtk3h5ITjmosD4c1rFAZRUb+YqpX6knSnBJw743QNokxoGt92XT4Q93P6o
wIte2uBq8Lul1zQKug5gwePbQpnpN688SWyPm4p83t7NfnI2kUNgI1NQBWcG
WQeQfhQVxBcfSpRPACp4nZXPYWrprazW0SsIcdfSpnzkdlgtRlC3Vfz5yjtl
KpMVGUVD2bo4IIwSsmGLOThr3/m6VvJOH8ewB+9Ra/tblmzPLdRGJju56uTn
yT3FAxEgjg66Jq5lySPyku4J4h69R6S62xIE4ZVD0a4u9BRkvYZBPMJy/g0C
vFfDfD5XrszkB8eWKKps19z/mKwbYZXIqONmu8b5wDsWwqRsMgkWb4JgBxI/
iYFmdNu9Azq+HPt2TOl4SK5LcZwQ0ZjR9TtCpy3ubz6PjhkcFSS0KoWA5jYL
Q48cbibMy01dgwRXSLV1G3a1zhK2MCs5/lxWOF/ni8XtD/0IGTFBfKyIc/iF
DsQUwG5grNPCqPBv3dySHpsU//KmC8AR72GrYuLe2t2bB+0/Isi4ndJKL5RA
QfVQ499a9GGH651FZ8Jrt/mC/SXRA3pEak6+DZ8UDon0a6S/er7xBy9s1qMB
jJ8qwX/5f/P2lIwwqawzGqfy7zc6oMKObzz0kaaYU+TsaORHweDJLkqt2uP/
GB/47YgnUpD2LU9d5dFULoZbyRNQT8Rle3ztufl977FaYJM1rh8Ja70IBMQJ
LFmSL71toG1oHH79wpNb0MNYLg68lHLHlRorhtTTc6Ils7YI/z9RJZl/OJLK
aJg945msDzG/2C/+HbHqNiPcOvCubfmN9LbOKvwauso6cA4ZYbHjBDTNLfuc
j7A+CGVsir9U/FCW8vB8xs2jo/uASgr945MtX1v8J3OGa8NZmKj65+aCLOed
xCmisVqOg/1mPTscuJYxhA1mUZnDWZNo8dAIsel4RNI8uDEaxQUziY7eImGI
IvkyT6PaXbZsV1hqJ68EIlAvt4Jpb7Q7p9FYDh+uOGT2MeENlQrzAS2pFmvi
uPs+qivsEDaf+BdjcunPppabzY/7eeKX9EgJy+PUR0gf89yxa8DQBz9b5f7x
0OmVrKuTeKipgSMmMdud3gizCLdu3u3DVSSg8uiblin6KKYzd59hsDp+vfK+
6ABZ7bNUPZE5cXnPLIF2i5dFnVsxSuGz6hRImwsWgCVr081AgVesl/6vh34U
wEbtweY3vgGuDu/zSVPp3m8/hhMgUMRtKsmkE4qbU51x30uZnilZlNn1Ts8E
JDRDLx8FUFFxzjVrJaEtg1psPkDsW7iwMXtZW7KWuZr3OWvE082wNVG0hck/
HoYze/DEL4Ue82n7wro0tyn3JllLXFrL3AXsokicW3xh4G/5DhL8bXp+JVKF
2J5MWZ5dE8wvh5B25Z0eOtBiNbkY8F9pN2VKsrw0DZ5gc+Bh8Pyu2UBkKFag
MevQyE9qbZoYOk+D04f9bRxXAjxTr0QooBP8Ga8+hI7Cl1f/jJ2M0wIEMMS8
L0bzP8ZuyM6/zYbFbepBnnz9SwXW2wiYCOorjr5HrSVA9zjaX/E88/IhV7Qc
Lb0LTX67Jj4DX+HcvlxzPR+uXtMdvghDdMZS2nhfROdUSAnHlMFeff62jn4r
5q7yhNMe7q6ji9fHju26pk2Yi6lJhu6SoBtbvMEPkYwhnTqwvND7NxkbjL1k
HBPCC5WNzDtAmhGJgc/WHwPDChSBzJtxquAkeJ7HI8Ltqy3mcM+qsMgjXx5A
KtRdPzZRjPhLCZ9l8iB8hlcAJrcaa2TphL09iPuz722+J6cSIHfMu2NcxbB8
vNCGUxYEXqWZicycyhrstM7qOP1HfbleOD1UhqUty1mpgZ0s/ERneqICzkwk
U6vPfGtdbgFcxF5e4gTwaUFMACWqBWyaYhI5rMxlYb99w7towIPEqHjR7zOk
jSZwY6iBVO3u6x0cU3PVgubVSirJd6K4h3htT4TKAfI153l9xzg7ibKDIO0f
O3KqQfnV9zWzaLw/X9ae1/OLMAufXB+dsuCYc9G6wcX1485McAhgUqmPGzjU
ZbPZZCffUKOWNe27HmK1mu0VWJ5SNwFIMjXSbVzcwzFq8FuEmeCuJq3qOk31
IltXhy2r3iDuyIuJIkjh3tICQCQ137OQZPzcp55T0HBH8mtdZU80RfnoI7Ek
dt97rT5lb5/LtcDsvMSihJqjVeTFYrFMfxT6AoW2zw+FCDc0f02BegPbVg2v
7ojZfXhQpjVnxLVtLBGEdU4cKQVey31JCuKl4biX66LeGEohd2CAf+8+xQId
5g4pzObG8O6TzbKAwUclmzktVwc3d33qDffVzz6NOsgwW29bBHBkPG7yH0RM
hT/KuR3FLdtTIREPD0vmr9MBiy5QYd608bQwUiT2KQvleWDEG8lEJkL0d1/m
yyNCcSgWr2hFDcUbH2xjuhvuxtKuqcBQQ/05lQVW2z7K8CByyUB5a83J4XNT
0aSnZJmWYJd5FS/mpfuP/EnKiXdMY8e87tz5KB87tRM3m6ikAfKG5wXibmiz
Cn2n+ix7uBmzrMu0r5JVpeNiz7fFVIS+rai5aa1eOQEnPcr9GUfa0DfgvyC4
0gssbEmaBsBiSi2aPmkS7NgJ83bG5IwIWgg98fNW3hdPBJnOEO+S1+saSvcg
JxyJbxEtYGNOlTrQKLt7jxY29Mr6a2KSqUNJlr433JkH7de48184t2usO3yv
ezxbhEzQAUREqtUHLxvbRHgJB1Ry5zyhtwZ34jlUtuCy9yatB7f6spSGB+bj
GD8pctFZzbZn1esMTTT6SEczX9O4ib4PXmkH5lNqLwpaYEGGhsXqVA3XtM4E
SXpZ5iQvCQX8dZS3Zf3bEN2gbeYqMjaTkXtxOwrmxFXiv4ccX+KZaKhGlUSs
6A9EaOxwLaEnVlF5RZ8nafRv3xnQPT3EYGD3hUuyEkuSHL/O1E8PpOanpmVd
9URkhnLi76iGL7nNnr+AF7peihNvr6Mwii54GpIYLrnW+pZ8tgsg6A1c6h/3
zUjS0yHKJHIpnKkgInzYEzOk3Y4ick0dwoKFEjJdEmlZndTesbJYxJxwwg1N
SCH0kqdW7qkwUGJHYTW7GqQ7MRe5BLW/+Q6wxs/mQfC3EJMsHuRddjVuhWiF
286ZAVCqsLz+QCc03wpyegL+BUyDx/2Eo0iMB5lzXgozDyIrTRksIaR5Os5a
49YUqRmPQdBvsYdttWs6ShBx6zvWQClCiJT+evbhCC8t5lHGiWaDJEzJ8nzb
Bz0JpeCMm+h7o2t1bpovecQAcGSSkWyUYvYRMCx46fikTPDw4FacMkcGGmco
FjZ07qLFjjyoZzjxn/SXpaUfa7a3Jv88+6z7gv30fBwf/Ybphnjt35ZtX2J7
aFBF0IBCwgrHSpph3S5Ajg8TYJ+EqcX6LNdWZR9m6jV8sA1FklcrBZzNiTrN
y2SJnBRGegY1vhhA7DHYA8qLS5QiK802xRchl+Bj5wZxKghH43DvyEUK7m6K
1W3ujGtm2vI3uqfy705bfrQbl+u9RWj/092cVvEs0hzVH4mL1e/vCbpjygpF
yph/cri69ReGHO4HMQbqrytk1G2Htgz2u4UK0Mwux3LdiXy2SnyqCzj21h0y
OqT362Tl2RYAX8zsOfEn1y3XexGD48eD5vKbdQKuMB95/zE2XH37WEF1OOff
THKlFP05YFXkhGcWUTqhglJpVw6jLsNq+FY92NJF0rGIm5EYxiyGCW35SmXx
0eHoF+aE01y5RzWvKI29ZRPsJnhPt0KhEJmZKqGq/1hx2QI3nojVNcucNdSH
5l/S1jctGcfSusKRfh/bWX+GpHMsnVva6dzyuQvrNhyPBpZxzGCJ+TnErPJ5
zUwNWiX433ShTmm8TjLaH8BCX+nR93WnaXWm0Doe/rL1WserV47/K++GrQBA
5qtXazG5XCgUNM3ldoUKhBcapffJK0ewFynup2eWrfTVWyguLc4jnXTSFrnZ
mqmduerPNXZz9ndfIqFR42MdyZpl6DJFJhEBNwCo14SgoTA9ZyyMg1aw8ZFq
q+vmt2sBHvmmJvV3q54bZrnuRpcJpq4rEvfLKvMygz4tdyQz/yUExacFciGV
D0UU400N3/byFMwbLJE7354UerNUJeqEy69gimwYDZ0+T5Z54byRmiMzDYgN
GHESvp5SDP0HPFLk11ZSj3VwrqLlP5W90HziRZE1M1zJvZIcBb1GbMRyQj5o
K0oRvlp7rTZ1UsbEpIBvIuLb1RDNVkbxLYYmMJnGm2AYCvRWGuGXlSfDx3Yj
g2VeJun3qLJIPA/TqV+iKsyJOegI0WvOx091YVqPjW93jXFjfIDbVHsNxIvQ
agSb4TTbV5wERV1skmgW58RoJkSHf/zQ+EhTXHpy4qYDhPS2A0Gr/XOXczRg
CkfkyyuVts5ntjtq0tdKMi8HCjguO4jxQyXEYs8Y4fGwFXk5DMbwdbH/5/SG
y1TsXycg95Gkt07TgejEaB1381vSUTQDgqnosAz+Iy/3jVsHC3Eio8UuOfVL
OtG1en9yviMe2GkFdeKPWBndIpE/9HZS/7W4FJNkY3XRbxNC/r9lGaUA8DRW
87T8trPVWXon0AGCpa5J/wqy943gLQngEn94HCND/xPB5Kd2jqtxecLw+O/L
NYVNbreoO+V5ikxCNu8WmA3YdUY4XhoAkylZkPJTV21S+ARhgBeyq/cr3QH2
rMhL4eTq++xQbFADb0D082qot+mUhh38bInUQLNaO0uoy8X7MYvxOwhMB/hB
CROearZzMYVMefoUe5oGLTj+LC3RBnSeQ1+oDa76JP53/JDPDCIwue9a07da
lqHuKAHqy5vZoyOUek0QaV0DXCrHbZh89zqOnanwJOR4C0Z903VDG0Ye7O6M
SVF8CmYEoN13JEQGnj2b1XLcHnzMQiE1SZui8JgXuv+ww/oGiaxdHAXOWOnk
sOHuNvc2mNdCpOvHsFmchuRjPUIuVmtS6nbQ7GL8cLMeXwmd3U4/r45tSSZW
ykgoNrTfHAzROkj2R/OVHRDS2wBK1GCNb6B+rCMWAtq5hXfK+kzrsiN6CGuj
epfI19VH2kL+rtlZ/72i8MFnZOgoZGUQMF51Z+An3OE4ecQ9naSXLQlSPngn
MBysaWsQQvRsPztuSBh2lz5tepGmGNaTK9Mrv3rwhfTvPnt8Kk9viWj2isXs
xX1zwwm8hvrfj9ZEATLxluvbpK31w5wK2UI6SG3ihHY8D9Kzn5tjaIgaSa44
UsWfAVAvQ1gKtnhnwJfZBZ9stm73Cj3xZ9015h3iyVexEO6NlaCrygKLHmfx
SgtU18uxsrfLN3+lcPqL/ip2c476jtvYpRSpXm5/pACqjb4eroxnoWARuLrP
I00wY1VN7jKNfUPP3qWoll8GEGIIf42udFlXORqHdl4SER9+MnpPM/KeZ+Sr
LCeGRh1NfYEQ3Yb4j8NoauU9NYtJ51hl+Fyy80BxyktDaGHDG7gtmEkgPvO9
PwpVU/RWj5Fdk87W4n9sszis57jxbtTkRflWeuPF1jJt1Sa/dswP9HB0+1ZM
bFzB63vIlwHYihsxhIeJ4HCByReAtyqI1JMZgCVr67+kGJzLLXzkDcHmGn5S
aTEBs2ky5aBLY+8H0oOEyzq6To8UNLsUmSdcn7Iae4DRHyyCeCu9Re1L0jno
9nkQxIPXr8K7pXzcLNhOON/Y3sn/NCkymZoHQEa3h8G08PyqR3/ixo++I9fY
btSFUvpfk1AajEK6Bp/uV9TC5AIBzDjhjjFGnqTt/kcqC2BHhReOAk5/EkVY
JgGG4/qyC8PL/8UDVq5abEY6zVnQkBVyr2Jof4H4TSzNt7TIRAb57O3KZXeT
IbsRWh5vwVsZc4+PJEt47ByC37VtTyObpK5tC5LBtThNrxcKxI20/HYtvgE1
Pk+8CZMxNKi9AR+0DPrkgs+f6EI5iPSgHgKG96BA5ogtEdIqVtJwoVJqNLNZ
EaVCqdzZP6ndtSydg0GAcCdh5viUWBOkSGjKT2CudpYSTqq+xyK5QIbSUWj4
1Qb00CEa7Dk2KIOIdrUtqLOHVcGFy20Rg6zz50XZb8kLER5DG15JXnKksCdJ
WVy7+LOj8EE5NB23qCdszvx2jN2ve9v/1uwYbAvgVC01pw1AuOUit5QyCQHj
TWVaOz/N7ogS7OlasCu5Z7B+XCfSymNDC6ochIiMFMKEkf7lxLgQGuSrzpGa
Ky0/d8+9vfOmz+K/lYK6mrFnght92uiibkhTPVS0ORAyADc2k8Ws8VE8RYV6
jtg95uxBTxapCNU6qyaymiO9ZXjJhgfT2yJLgFwLG9QaYF9x4flmZx4a9n07
GLOQ9zpCVk82B1CO6HkkNleSFZxWcQQsU3MXWdg9YFiqV791mf3T+EFTjOyO
7CybkEl4lTkH4IGfkRAuGYlJ3F/TIlA6VTdhmS/eY8sgrsx/pOPbgBJD+iut
IvELuNwMt5nvQJIrGaTUM0+c/erkBFtYfsMWuq70fziIEfcIR9vLeMsmfUi7
qKQWmGHwcFpMoz9cCziVVrPMK8xQqlAETXwuZWGUFIXWuwD9eKRXHLWLeU9B
4uB9tzA1kd5m+Yp+pZzSDejPWSJPwwWXzdnBRwFROSWYtNcfNwf272LfWRtW
maikMzqBvluC9reTdQNNiRT/aZOq4olkPJl3uJssf9reZGFbnmhRJGjsWRGC
dOXALttaOjDgcHJ1BS1ZBeH9F59Cj3I9j6V/pj7j3mWW+nOIvemsOVKFTAmJ
8BD2UWEoet3byqYyfbP/1fu+J/I1iv786H+wFOHfwJuU80jEi7Bq4v3Os8vW
PJ4i4S0EDZ1jkay9kYekn6FlGpDhACYjVXBTunWhBv4CKbW7Zo2ZAzZB+YtS
ztTa36YeOdlmfXBJyh5wZOshvoCj6lrp/JA4ewTqFJfdDAh6pVGWbzO3VlFJ
nX5NSxzdkMzHJAiiYBmIUdWEeLstwUhd1nTRbXq5BlypS/g9nyv1Ts+JJVcl
SnCJAAXRel4acPRSC3D+aQWlWQGtzysLjza/pLV0xEBWU82S0sJQlgI6nxb5
lKeQkVG1S2u7y02UD75dXw8BiCyE4AkWrdi57cyfMKuL0gxVTx5P+5ojO2T8
jkRA0EDzu5ksvRZbRKg3H99SAjm3o+hT1wSopKDypQ5dq/+yrDtC8pxOIo6I
MTuQ/6+uUuZP1QR2AX2HSYm1Tsma0S16xEQ04pTfl45oEuL0uDzgN3zT9CAJ
sNZ6/rBOZU5VguG8OCPeMv0Dfp3GjtdQITcpR138/NHRJTqCJ9C66wklPXKZ
RpkBhAMQg7FeT59ncuMSxRZ1FTu7nTp936TO1B8iXOhVDGU5Zo0XRwRpoYjt
3J/QcrPEYSoyp95MCUfv3i9Xop4o3rTfFNyhv843pXP2/+FW3A/NJKlby5Jp
Ny2eKDz2H8JN1uy4Pvyt0qQzQjvakO267TTwW1DzwwvjMlhyFvQMwD3NC9Et
JYeAZvAsozxCWpfYNKhcaZpVEf1JaNk9nQo3+jEdfmLn3++Os1M0PLxde41w
Cy2BNB7CoXCRRTuDvKIjGnEtk/g6P2VXtMalxpSWolCyu4kahhVe2nE33HL6
EvU0MVfyrGnUqSODgwhexYqkOY3asWSktQhdTIDZKM4q3BT3MX4DqjpXKG1c
RltsISnI+uORyFl/fRs9wcIXQ899EY7OQNFWpK5bCsg7fN5JEEjTBtv+4MiO
FM3YdydxrctEm2IEV6rYN3QD5HVBDl8Ydf4yN8LhN14Q/mfPGbFhqlalNWYm
6nX1zFQe/NYh7rSLNSl3v+i+ZaobukJxOQgetHBrO45j64Wpdyb2W+TCl1Qq
2Onm3ZnEFMQtx9/3zPYo6+vrw7vjyvKtgRb1NX3CJBgbnJkECKdpAv4lhsZJ
oC7jCftEuK+Ix7dgjabTLwrvynZ4RS5S4w0fUzPkyIlGlHv/dGS678noEfpI
AUKTlJpTsubNZrYMRpqatJJY7iISszqi+mG+o040mCj6EV/rSof3RH//QHiP
DW/9QUK1MBq+ZHxMSlooKwwfKEqvkBiaWDfyQsawDr5VK/VAtMhDf5GTyfZQ
ZNyNpTJg83Svh8j1U5mZ4z6lkl+rWDqEm/7UyHQnvFs+KaDIZY/Gpz333O1o
pmkwUM9sVp9xcBsmYR1kzXIebyRY3GUDbDylyFqkGW27jUD1dJ7wfw9xe97P
wKf5gYxd/yiyVyzv3caFy4r2ry8WRVPmiACx/jmxgKu9xDPJA4TbC75zPs8s
nfSbEwHiW05yJ+kkRKQnvSUt7Tu5kzKTI82sZ26hvqA/tqpbHGPEtnjwCzFv
j7vsApcHf2iQ+HgPw+pRtOAvOkXJ9P2l2dgn7rHRtupBwwWmlTOF5l4EMJvH
zBOHJexxw4l8oTPHgr/SpBK1yuuotCSIotYUaKQfylLtuyEF+7lALgGJtCR9
NQ3ET9BeZDymUWtgtFZfchlgB0mMWtw5Zq7CSI8rmvbGuaNB7VQUNgxFawaZ
J166Roq8gjTu2QWvRN5J8EKFrMAX3IYH3Oefcu7DLm68N3tn05fF3P0pHfNG
wH1BShLnSvP0WbJ+nMlp+oQChbXquW9Bkc/vrDBa5dCoHMj1ff9oISW7yxG2
JsiqGWdAFpzJ7H7S5rMv1NC72SFdETEb3CCTGsq9dZtgg02XyTmC+jjCfwcf
EpG+4cUkDbwAgnQ6atCQ8TgJvEVTjTALIOzTTs0PXo9o8/YE8MwQHP0nXi5M
iwSUKixvh91bI7puHHmFPzBQnZcx6aDbwRJN8Jv/WJayVUpc/nu+5mr6OnBp
GktJiBGpqntRCVFkuz8p784s9rl8sXCUCfFcQGiXhygZ3cPA9GV+ZMvHkVtb
SmqI9HtQk7Hr4qmptLP6fR4v8dHYWQ/3F6lSQ04dnCrIYT6CI4PTxMMKbzPR
eSxXjovVjOK40GDL3CqaN3uOadxIi4r5H/avWcKjHF3/gI4gES/jiwuAvX2y
EuQWiOj08Pkg8znezVXOca94/s/BUj4QG3MVg+TN5W0Z0NuaI7o21AVgtW96
BUUK46I4aCZuTJAkPYfch76R7x6cRrXnwzPZMhGJ/1fFGNBbfDNAVQO2dR6Q
06jZoUb3eWBTELyFe5WuQTdhQQ8p1/jNn3yKvaRZROTkoA5G92XQMmoS2uND
dvDnfVqxzSNLPObH7uPtUR0sj3As+TNoPEgVM7JROkV2zdK/GGOUQr9cgP5n
1moCgUCz2CxfdzktOxj8rfFFOw2zreCS9/TriIq6UBKWPniY2No1HdjLFjDe
CQnu5NuodSkjsb8FaowGVrzwsDpbgxZjbtGyAGzBaL2dfXMzxQlyzUNT6o8p
jLoofDvRtZJwZN/Q2jQAaKM+W16J+c1HVJdHq6uSTCI/b30IeYBHtu2DZd9N
Bw8cRQxWnTKaVSxcep5tcWpHoXz3shrh7NqPcz0Gklv+cpZ8/zHnbREhUt5Q
C4+SPaDSBrSMzFz9hfq53FUNqA0EG4r7l7vHKMZ09Ws0lX0s0Tqu0zzw7A/F
tXKKnac0nlbaTOrlSPceTHA7Vi/BeQIEgZo6jaseuCYBACcqwIvM4v7E3lVc
nezb1gcoGpfUCc6poPiZXSO97iMJ1+5hnyEN5iw3viE6BJBboC8M8RWH6qOZ
X3g5x2xOcJUzP7OUmASXlRTFfKt+NkVkiq6VyUlUA+cdxhNXNTX5kBzAby5P
xvX6uugmsqkX39JlzRjKuuMJKrfEGjfBkmrzECcUYCTXb607C9eSrmkbzJi9
X8mDrUHHa0bhbhVsBMVOcx/ZAYczthiBbd8UxKS6WIRhFhDlF2gM3wKJJUQn
owhcKiTxyV1KwnRH/DVRIpWH8OWvaFZ/F2RUuGkzJH5cOyv+ie5R+zmcQ8x1
wiDkhnNwJUsVZLuF94Ko9FzqzjQiWXWs1a0eMTrtBUCqnOfqOqbYhd755FVZ
GlHq4pGd2zudu74frGKEdg2K7yGgiTZUO0mc/rgZKVF0gtJd/EAFcaG9ScGq
aHQ9Hejoz9sY3fF4TC8uap0COwfBL6EEEVNBIkg2jLWd4/Aq+BrcgmD9zSNb
TYyN7q48SipTRxiffVXp3OFwD29+QbRgv+0wjJ9BovcAZIoKj1vT+h9tbKSH
+8NwaWjsQeCN+q6ejo4/dBfaZAOn0BBLqnhzp2Oc0ZiNTOID/OazNYI83XHk
fVi4ssizQViGNUC5JwD8nL+V7OHSRjTSoO67OrlxLU6AFc+FF3APS9aW5m8t
BZcXL4a6PED9BJj9baCP3G693Pz7CTU2a3eDwnxm5cRmuE+Xza5lDfYBt1SF
JNsRhRa67dhcaqWnsKa9A4TT3MabYfAxCSIhPOyiIzZ8Nv4Qxux4JjZ7h8jz
oT8cfKP6MtvTJuASxpavPgWE6sv5xG4Hoglop1hwZNN/5albRsdctloNvIGY
3SGOexzNx8RYIuQ3yZgrugj0A+omQCcxl5lw2WEubrghXaJOhStrBGkWXlUW
0RBn8QBdbd1fnd1HBrcairvbblpRCw+CIu5cJViEKbLnZMVaC3QKuDIYkFky
AlKLm/YfCtN2/7gN4MZDPcAAvPpzGXGDH33BImJigNrAAAaQ2ZWnj4tMCyha
hlZa4+77xit8izlELmg7NbMDcai7Z2dYv77m8RzLu9YNfFiLZxCqc+ehafYW
atN3bz+4mDAPFiRkxYzbb/jCMJMZZrxrCc66JhIrVN967yTG47j4ccBnuT3P
7UxKFq1SHVARmsXz7Ls1Q8+45qcA4+1CC1eBq7ArhoDI03ue0AZGRpFuMP/i
IDQ4KPagf/JXYRLVnKnplG5L+xNq5DJR1wLtVLu7cPYlXDRd625EtBJGEN52
qNrAPrhxiUJ9x3g3+uvToboCr7rbdz7HfEx/73lZ/yt4XEHCfB7WmSuZunou
+xZ89b2whwOygtfuKgx3sbzN0lQ0EzIDuRS6U8jLmFhcGXsti9KPQLRtMlCM
ZnpLeUzr/0BGsttEg/1E8rW/REsOrKY99X6VXPuSw8Zb+4O8Yr74czbDJrkn
ZwMtL6oTjm2FRA59i0whTIkaSdlR057yNXPPCDaAYMEytVwCTfUU8c8eCkWu
94nIyYWbVtNeYi6Qmi0Y5uSZQjilIoE2QXzY3pQOZhTwdiE3EC0zr3+vz46O
6tOb0mUCTVq1qZ6a4AwQdaW3j3mbPh5CsXBRMnNglakn/U8YMP2xq3u3OKeb
rvjMHfqZ5h7qcsU02uToYtD6D5/nqWzYHWtKfCFxWi1h/4hUnu68aTC/ioS1
GUuoj0ZBP3qyvwUqn4jfFQBaJDR7pvFXaGWiTL9eyXkTv4M0Fqw4KTsjiRVU
x+sE9dOa68Q10SYxRJgBeuwxcd0JCYOT2vFlcO8kLlhrumbq7RJ2uVDBRR2M
ZolEcMGQ132JtXAZspxWti4zAbH9imxtDwFmhw1ykw9lW5ePEAvMxhS/bELy
2gAT4l9zqnslC4koasCLlRQG9JxGqWmZeHgjQvSd5V+3Xyr4SFEy9wlrYSwh
qbLBxULfHN8U9vkxtlw1NzJlz5G16rest+b/hkJ5mUqsXLRbdjC/rhzdyoyP
HCY+plNxuZbjgJzr+wNa2pkVBuQG0zJKeSM0DVGuGWrDSTraYjv8+m8ViN5f
eTYtEVcA1RrdCiM5zr4RiJZOaJ7HVpc7TFYOYGNScMmFufgPKz1l3svPHGDq
p43DvPNwhw+5WYVB6+JnndsBB0q2alqvqkbPvzCdpUAgEJ9fF7gxP9ZiHMZ6
IDWUzjjIdJftQHM2aHjZoidLzhK2YGcl7aIYz4Uj0K6PQFLNVckg7WOYPKfr
40YnfMLB1hO+pGBJo0oN1SJn4uAm8MsbNjLVvMViyEOW1YLKfkWC24ka3Szk
Cvi0nHuD/KnvR2h21NGPWam3GBqY3VdJzRlTSt8MOgJBVdeTnBoTI0v3Owev
J1NaWtalJTzmHs1g+0wYxYQxe2gu7BFYgBeXX3xJHHZydnZiHDMmIRzc5OwF
aAYIwFcTLGTpYycj/b/rV7Y5dwNcyz1hbqvciEvb5I+DOTVLpGN4dzkNADmJ
6LCq09QNmImA+j90/ELd7KLJHICTmXGhdCSTPABBgpcUQo1sNvDTNIAQ3Xkp
QuarTK5pX2DCr8bpxVdx8tNQVmIcudkizv//cuJ6HBlYJFF3uRMganPURIuZ
GiViA8mdPWbWYrPY9IPsS5X5NS4oE8sPU5PkfUO3n45TcMjWSTvsn96LBcVh
TAnOisJE3bWUkPnS7OeQM/58XRZUqZr4Cj73WQ+vRviwEm5jduF6mYKyRSZH
8ksCmrcxLlegyXnqX64l+WosZSdOumhTI3eUbdps2HcMWm/03RWVVerPnl+M
Uqx/HUh6Fkuo9r6kcDsmRX+1+F7MFzsYRmXWpo0NdJEAOq74xC71TFLQp6H0
4lvmHYSm70PvIFpzjV/6GZ5E+tYepHYsHNpqE8aCZfMyX+7lyRD7EF4qSFQ+
iEXGI5abiD7tcDqgdM+9xt5kGXN71tB4rELuKowW4h566+JSFjHhRSqMdYkn
gANcZW9w0lXo/AeZ0KGTEazdcy9/GzGVT267KiojNF5l8QfRtlAj7s++SoHP
bD7k/Pp1ic9nj8LmIPDI8f61mh0JFp81XqQFAf/oso5I++b2r5UaEFX/XRgd
SnRmIwcpTylAo+EEO8yn/P//pupl0EGJ/ikX7wTIr8t5su08UvdpWXnvAuAR
izV2bCQ3pJG7qIoFkCAKIWwrZWX/hyTYkbvI/6dW0jYJEeTdCUJ3IWkRqs3K
PvUywgwEOCK5ZpE5uPThtCmoLtj7ftBRAJMBH0+byby/IPC7IA+lB4s3SXX7
ucrj1rC4w2Ow9ThHo2jAkSAlbp1G2zvufEcOqgv9eHb/AvYGYbwd04zohgWM
hulkpO5sS7vaH+t+U3ITcoQCSNgRQ5ufTWeG9FT65C+bgCIqsNMbpF82/zQq
O8eyjkQVzwzvegRRetIIj66trqC8wDZiTrx2O4lPvf8rtCKaDsyYyPd2VuRg
OUadbvSL4aHwcsqoyw4Vsazsl+1eBhfNXK6U20ynVKzUTyEbidC1iP4TssQh
Nogh/pHydEUvs72LmoibWHm1yUcc9DL1k/lE1/rfTnjwKSNtdwVssd23Lbom
ZA9pAYD6szH6p2eXv26rOGsSxzEx3cGJgxCfpu36YppeN89v+K1E9zjqGxG6
jmJHb7H8q06mprtY+j/sBbOXMecNJt10sHrQ6jPnk4ICleE7ui4ishxgwx0J
Cxi64HJkjhd4pChcL77aUtgL2WdI4Rp7mOkEhb8RRFnmwQr4BE59e8sT21M8
qYC2PjUEEBb76J90wCu6E5timvZC9RzRmTk9OVGwz1jFrTOSkggfFi4pPpx+
42fh19var7AKoknCJkcQuNqU5dBQtfjjGOY8aG+TYjwfo8huyu5nPLRxZSFa
Pzk5EwJtBrR/7sXTYQbsv3VhXAxug/CWNtbFLAyAMK85YV23l6+JtKPpuW/H
G8Mv7g+F+tQllomBnM0CnOcNWSjVWIjsahq44WSywz7iyjvL1kK330UROGRD
2klRkpApq1q8qbFWuyA43qibt/hpacZ4q2Vt3Wne8PaniYSWIDXutggTYqCI
cclXfVRLIYUovX4Tqpmm7MrfWvhbbQG+Ls3N6YivcbsCg3wXNHjHzfLicYle
kRukFQ6bmq4GHVhBnHfL6PVRzhWQoBLhBltK9eMbNR/5ZQRajX0MwCPHayOZ
2goC43AH81AYGWBM9rYGx8jgCMbRqC4oB5WgAYh0edKWyOZ5Wm3DuHql1IS1
kzQCi0biGBPEi0/vaIVCZtkExsed9q4scz52G20csWs20d0VMQW+o69zddoU
7fVXuZvXjMunlypn5KN9BQJMMkhjXvNmJ1OCvHz4r5XVbqLKYP7XorUqjlKv
cSrn3N9irA5Z9HzVNLr+7FC+3QMHDwv5ZXnQ4Idq2vLKkv+5pOXFF+GInk9n
zSbnS4yx+MM7wQI7xB8LgkcQzeBZ7ZSbuo87WZklO3ubGmIj036/FN63g9T6
L9X4tbV9Q+vEXdcoDLdQ2m35k5KGiGMa/q1+vhIxD5aOnfuwEbwnwFZgFlXA
3Q6v7CkRyYjbG54Q9XBGKVNbvPRlwARHPhWKrLlnXdVQwczU3SSAw7ONYFJ1
ebWexhHWTt07RlvlrkqApjxaGenXWdC0RbKxFWGJU9rNcMW0iAsDi4O3lMZ0
FosfbzlkQU/bHbIcld2ZP1v/KVB9xfzB/+BfnsQwRfIy3TKY8NDT32F0fOD1
CeyoS1/cLIeJ5iPD2Vr5dc7RqqCIbAioknHogDgCIO6pzrtwA3W6kkyPCEEu
tbn4gtEJ7Y+VRL26Ix5atyjcBqIv/TvwTz2Ib/ZyNNXiDDTysPVhcR//S6bU
u3zaXbbhW53bb8RhH6eTc/oHPmcLY2pVJ/258Yk2gPAig/4jiI61h9cfiFhN
gDH6RK33VdoN/Ljku9Na0AGhrog9Hnb4b0wbe/GcTTQtsplvKPKRAkGDf51A
Q2mu6B3r4OcLZO7WHXgOoDa0IIFcoKAYHabAoRFaUjDyRQmocXVQ/07AAW8+
Y80l5aJubFW4coEQTOm+Yb4zPqHvBo5/DGbRonTY0mggAOhy5gZox4nUbadm
p5K4Wa5O/afgf4cEq7eORk1C+Ggq37Xy00ONKtkLvUeOMPBfd7gEixI34E5v
bhI7S2uL8iFLKfc0MyeJlqw24xYWEwXWyoT7jfa7gZD+HFO2tMm81diltANk
/alL5D9K4iijd3fVaQdBQxnR0UDycHMB5LDfN4GXS/InIM5wdC72v1Ne9O9R
OjqYDG1GD7h73Y1i014v5IJwzU6wTqJO8Mz7C1NEfnkNeNusIigMX5B5otBY
bLX2qkNPtcdz95rFH5z0aMtM+D2+BCBcSf0s6uau5Fo2NFo8MnjLyonRbzRf
+zXnnYqzef8OP0bzXV+/B6Y7Us1NKNBYMHVREl0+BuHjfycVQ4tpAE/yzvn0
0GHE+J6Oq9GSEF6o07L5ghM9z5iiQjRJPzDYG/lacsVgfS1szPGboXXs+ALc
b0SBpag6qSIC4Hc2Dae/Wzg+ENXRf8qRke3hue3g3UIzsoGejfcDKEBRZYSH
05hC07oVfDBjlukJMp7Ecq+budgf1EffLN6HyJEqQThpRXvy9xxjqYoFCohJ
BHEw4mOoHWZVm0BLK5zP0alDna0iGyxP7ZoEgADVHD4vHiNnvwkX6U9oDKhX
mpzdnxS83lfz9FB9qun7qgN5UzZHHnpL8/omwX+OK24ZnnsihgHvZb2JBcLY
zdcD0SqCWeKGvcjoDAFUQPg6A0Um63RvBR9vD4baX9zgGnA5AwRsQjyCA07k
oGSSS59jdasubYpOx+J3pjUfeWOynz2KATF5nm04xKyBnYsqGJnNap3pswmx
3HWyG3ha1qkHx5QuL18VFNxspi0UpllK9iv/BhJeuLwmi+8rGs2yoYVsB8kr
uMwgvQRD3hrv64bt/UKsJ9VUvRc/VbzDmJGg36wI+UWL3qzb7dscrDOYGRY0
r3OKweyQJTBFMWbRXoKIELws3xojZGivUys3fMkFb+MtimslIBDGPJpJZfO4
lRwm67qYfyxh5vtylNV6rVaTdIwtP6sOXbD+E/0zKA8Fhdy4t8laCDP8npql
+KhbhT8661qupWL0cEt4YE9hEIpj0e4Y9lbpLDvdoiBSWWqJAagWxlldqq/q
bTnH899WiEMpUe8Jq3aoYmzbjrmpSB8d/N7PKBz6U+NGDNzkmuxsgezFNpP9
3uEeL1g2/pRzrfYzWNf7de7sXtyNDw/jXlwTbX4SxFWkuHtlo3sonF71ZNai
FskpiuHazzKJW+QAdotBkIMxnB69AswwUtpiy/O+qv1m+5kN2jTZBQZ44cw2
Lm06XAJJnfl8dOZLOts5fGKR7pVl8Q9TE42TagSLIAaVJ5bDoUnfVqIEoWde
YgXgYoNmZGCPPUZUms/dO4PERKabhCvfHutk6vaGX0AFq27cq3mxb5gzfH/U
M2v1zro0LE0STFDiAotl2AhJPffg76ra7M7scoh5+3HKiMKeVTq1O+8wn6TD
YmytKf/ENCqBcGUK1tt2aqICGWc/LRT2xDPo1OXJFr9C4kOmnb7qzZ8uPU4u
ozfSBXdNgeOStkDXT4tUePkLBauN/1s7bfgYRCU2PBIXEiU8MTeO2lYSsY2q
z1VCLZIB2bBHvfmsUvCkD2i4lzHWh2Lc6BN4NnYMHfM19oFfzp8RGHL80irX
eijTmcjPzSxlBwRsBzmavLTZ9zcK8N5KtJ4Uev3rgt+IuQpl4I/2ZOUgQkkr
Kw7rc584lGfmSncQj0Hg7esIQuWMkjiICAZ2ke7Phq9PVJDfb4hkirCZo+G0
tQ/fJCJnijEC2hKvUBbPiiadMM8VD743poUbhgIJTw8B/Bdnmapkfip5VNjr
pz2Ywf9nPizpRuGej/rpSFiGCbskXYV4bx9tvsMoOtmBRdmXUwwkSqrixHxp
/K++WyTdhFht/RbIWkXC1f09VLis2+kRkWbXtcBZDUFjqwj9JtkuJPo8UimF
1831sn3PKozF31E/uxFLgtqVetB78vfkO/WJViLDN24ZkwCxIim2PRYwvdRo
E4hjbVop4MhmL6axsUt18kVlI+Qlt5Ruu32imLTweznAfTaRV3iuKFdweZvo
H5JHaGMf0E1bRgiY39GtZdEocpZ2qoRUCr0QuOEjoJdaLYv1OhxgRJPNWokS
9l0GfGCNH+80zd8KY/Q5HBOYAUlrE3nX6fWEllr8LxaSJ/OpQtcOYn4JgG+/
RLiUZRF5N+oSGxJ86VNifnCnZukA9s8VgZrVn2AhMzcqVIgG8Q0uokcMsfbi
fjdSZSqwveqy04clpDgTwJZEUhymVl+7zfKoSC5bZIkwaijYEONh+rr/LMCN
JM6wVjT5rVNLoMpI8tRzql2UGkp13U8xzHaakWqWhdxApktQskFV5JvI1DvS
zn3BI3KyuOzlAQqi6Gpf+vAZ2QUk9GltmOSG1i/KJ73QayQgNhgBdRKqJ6E9
OI5fAWMAEAH0q9jKt2yCZZokzDAeqZkUBoIl8DdG+md8E82xB/JSeTHn2Y0Z
6WiYI4RrETYLDhcVdnsz0yahR+CvHzdNKMokQy0kb7dF70y+gquWWMC1zk/x
iULG+NF7t5c7ldp7UAtdEXrZvpEt4oTQZ78jEDww0BaO9iLJAUGFZu649cAA
fp47KYrX6Ple60Q/iLRoUe8JbforKay9w/K0sLRiSF4As6PMcji4IRmzZgYL
mmdLQI59oVDvs4r2F2YX6ypkrNBVSbgc7FhBvaT40PaJQ49529H0R5PvJM6f
upUd1lby6xAF8CfJEUEJtDndtasfLYA2vs4cGkGI184Up0IifYE6TJ815dMe
gMatBDmvWtOxOqpJHNmIkVN9pLwJS0VQMd6IMkmveLyqbswDnhTeBQxQNBPl
NNimij+ecEBKv2S96xdaf3eEa1uBME9TO8BuC/YDuyOwFvk/uPxFkAOVZIex
r70XQ0XJ//04wv5qv50Iz+UUlhE1O92P+yMw2DWWhwppxxdrmp2IEQelkJpw
ha1LoWk+adjn6RUPgINQaCHNj6Be/CEYzZoZjw1PXktkrtfgLRRg8pPhuY3a
zMRQRMbohFSC552pXlVaIv5HCA+P/X1m8q0O7UR29Tfjw/zQrhF3CjYD6l0w
JfAFEgmD+yyv1F92A9Y08kwJPolsY5A1xQpwV3HOsyMd1oqrGZ0158zxiycm
GwtEjbH0N4c0vHIzFunkzsAWpvGVJfzOU4bTLPzpx5Yv7GCaROf2bmy15xAe
V0EQwIkl9bOlsQgTtmSjbEa/brEhXp9dFcq3MizYKmiNYP1hq8cvEZH6mBQK
djXtk6N1jixr4B/0HHO8gP7OXOjwz5if+IjOqt+XQtDfqInzTnpdWhY5YJkb
1/dyQpVAQ/po4XWiC1WXjqI8z+yc87fNAGNwjKdQck23W5CZcBTkSnOkXow2
ol3js19wpbpHhWtqPYodJ7bMMzw8dDgVKlmq1o9U7nueEFseNuD8eZzMVRJC
PKS02pR8PAjQULuAUuahprKUHdbY146M1W9O1IlB9NagKtCe7J1+hru/QU5p
/wfmzK8DP6X4Xj8tGWdLJcGB1w/fb3KpMxpsdffk7Ku0Cbp92XisRBdfY9EF
PhhZKcY3J8XHwQgRkkFlCo+Ith6WHQEoxHKTqkoH/DlvZRNbv1cCHfdssHWd
nMBrTgJRrigxT7s9StP25M1kSly6ZSibWp/MPs+kebpoaYK5P3CG2jQU2jil
JLu7lyTqKz+aWHuZjkj63LlhGy3h3pH6f9LvfE8+dGy0883xPO/IRVspRyol
Cx8So8vZK+lyYGxhzr2QlETDV7oAYLtarMM/Wlvf+hKMWXEd1fMJJLgsHsqO
H8qXd3IxL+rAH34ZPu+SBBnXg8l/uI+EpxlTyhSXkd7MzpjVNEPkGMVK1Y/b
L65XOFCPWG4MucLe2W1tZxVPLlOzQAGHLIyN/u8yFBBrei1zgoLEVibhUo++
YU1OOGP0/yrrDLLubJe2K526MRUCjsck/vitO/hOAJ7pZnVZcWcqdXa7GmPe
+8H+WtqgDHhFjJFF/Yu8J+VfIB+Xh0gxz3PYDXwCwqXdycHsU6jtS9ZYY1UE
89YtdR/3rYc1fIyr1HQTdu7Q3m5XgPDMqp7Fejcd4jJbsk9FR2dzxQaXMeob
gKcVjCyUA6f65bdNW3VTJzfc0R8ElqowU9hlZLZj/CEInRLh0NYMwQjAiS1Q
i8D3bohNtnkF2+vdfsTBe7E6qeQXtLP3XPRH2bvbgaQjNVC0cGgwhoOBEHrR
PvANiM+8FsUj2QgRqLmCLacqS5lxkzUx3GeTZF3nhGCfJjHXiDHK4s48LCY9
gNGsFFOiWOD+zpgwKA7WIH5StzxjSEUvdHJeKjBeVFKgDm7M2MIHB0OJ7nc8
zNJtUJ9PLXaKYKnbhWBxfMyYho+geIgnm+oBYsr1cybglFMnRHKVb83jn84R
ThRiJuc4VZibUYyGLLF9XtackJtMYBna31eJbN0zktz+2jcxVr3fhDn2YJyk
NDVtQj+wrMofrGXhQuH3OMmio89Dyo56pYt1+E4mqu66jiIBI8P3rVxmmm7c
Zk+CvAcffF1br/cqb7+z35dsdFP+4FlyKRqvHDv8J+vR3WiB8OoHvqCqZmDL
xoZ7ljbwwak01ZCAqA+KaZ1Pzs3WvhuAzZGYccSMhQYjkmfujlbc3lv2kTef
Z364aH9/PJPIiJ++AK57Y2EJmSfp3j/kIqFBVwe6j36to6UN5ttdAR2la0+c
O1uU6ozLO8hqcICqVTIagtRP/h695b53At4J5n2LBGeLYevqaZri4ZhZuWV2
LhS2TnGggLfmzXqkgr5bNDzlr3SRAiK2Mv91vEslcxUjYKyt/z+R0bTa2QmJ
1btLUgVaxkiP9VYctt6i5bt8y7AQnynp2HMJaTx8/9KFapWN9Js84dQSx9Hd
1DWW6Da0bZ9jN3UC5RNGHznD/p4MYxSFlOUjOiQ6+3x3Trk1AOiBQHs16QVV
kRfazX+1BHeU5t4cAumZGO83SVeRibPx0KlY08hiWor1CpadMlROEYonRV/S
uiCMGu3KXCFmsSk4bebpFSvK41Tg7V2wo5YjDTTCpITLyNss1hlFD5XDbN22
SymaJs85j/aUQQwOFqRgTs3M8HngZFIJb8Qi0gzLX1vMFCaU/7rgWYfS28OJ
z7/7WrpasVuJKn4gr6CXEFWeaNG5ThQ8lg2SkzjIsAAGV3u0jXWI0k3KcW5n
kBugrU0U58k0PpI19wRpshzxGTWb+iSuwXd5SEmIqntqtfeXDnV4erKE+BGX
46MMBiV6KjjO67Zyy1DUCFmM1WhPTVmukmn1nuFdcn0mqO9EtQkjgbI2aJZh
kTMib4fUrBqqZ6tB2S+8I0ffymrT4Qw54ZWWxUQSa4yqx4mHZ918+R9d9lRD
BslQvDmV8k2z9lU7jmCv2y/ihsQ/t4ORAovedxmr+jHIyCclnrnIQ61JPoMB
HuG/CN277SntglCnQbxAagRWI+zXUBWTkQJZL2VP2hPO5frMQijIT+iay2TJ
mVmhZ5YQTAuHg0sXuRGc043awf5V6Wm89ra+29LREye7vfVg+xubllB4pnG7
lMn7gW+vmBXkaktp0tp0Ipd1OuktOnuvSpS4YEbksF4l4j0r3nFo7zkmZQu+
9LC9l/prsoueDlGcYhPYACcp9jBTO/3dsi83W0kfFZnWWQtDvvCajBjPR/yJ
jBGQvUT26Uu51aVe0sEgFZTCfA2Ib82PRMIWvJz5gA3sYnR2GOtXukyztXjn
Q/k4uiQt84xSXpqYNYMh1sPOWy26Kizmv9tamXYqN5lRm6ugNrpzIlXwlzp8
0BzubJmjhc7ASncSnYFCzTfC0FBr1PcVaRmKqbUcoAfioGfIMq4Q8svHMQwX
XJ4KlafA3EOq8Q5dG32kVQD7BbcrkPBZ2UQEBYWeryMbcWMJww90b5gAnAud
6Hx1g0GqRG5PVBS1+Wrj59nFlvZ5LHDghRtS6KSBfe1LulJoxUNEJ/p+aXsa
5FBzn6zjI8YtpgYNNqVDPM4jv9G+mYvKp4dbYiwAHJtGfyY/RxuzRNNgEcQP
vADAzz8mnPNHhc60XG8FKkPQPfyuHH+i8L57yrmAA0hf2zly8JIE6WfHSiju
GceED2TTSW703D0DraZaaC2CDFcrP+RKmHztaPvf+gtHwzZpbRApuxHrIh/1
NC2oHWwWO5ji6rMLcRMrYzo8FFEFyO2RAqMrVehV5K6Dn6SpJUo8Jx0XNBle
xJZhOkmShzKxJnlxt0xVRiLHwafM1/h7GPBR3UvcM4swfqU7y2MpcU40nOst
BFjdDsWUkzb1Ap1zH+y5E58GtJTjpolwI04jZlsvfCNCwxn2fg7bwt0nzMmv
rmM8ZS6bcNTuJFEXGu57N3oGZC20YDYlZ3K0Y/ewIrzQP4S7l6Glo7dfY1ep
IEU7yRYCJrLIbfUQOdXEPZz/DJhpEYea3QfXT+Yr0DANBynmfYjNnPdn8XP7
JGUTPcT7U0AfWze7yQa/ULSnq4zMUY6rV9c82vV1mSomZu6JIdI98qYqYlia
vKeO/B3UbiVEl3kjVNQVjrlrWbznPT8hCE5Pd/7a+8WlCpGoVERrjLKamQ+b
5tM914bY1bzPAx98JFduTv0qE+ZcFVL3umBITAhvCcXFWYwJ2TC3aq3eyK9d
BLtecYmV7ul/OZqm5u1MQ1JxTDE/hRSZjgAXgelsCPFA8TelhaxSRulemRGi
CmGtMr07nWGe+r3YBkRiViXWSj+NzMY0k6NPOqzoIawvu77sPKBvTSQmt42/
uDO/FxFP+d4L83unWRqwCTjNfq1wfipOJhbAkHZzmZUDgLMyd3LKCc0LdCJt
LNCdWC8YzgZVW+G3BBE20NWliUUEmZkKVfmiG0Jtgl0Ms/aezSQyp1XtDVxM
Kw7YnaRND4iu384AzYTxfLLFuOuV6M4X45B0krNcC++AdtCWY4Q2yr2VLzeS
GKedRQNoZ9+K4lAIYfoT58DZ1COBgtkukrt3AIFXb+eU/mboVSwrXvfoziov
Mnmagh2mGgXHxDDSM26JIqXB4eyPC/q8/Y4kHUicNOzMs3VT+WXcNLM5oBYr
jDLWREYRTSn2IYbF17y+8hWVEYbrmZZtMcvGSNPKO+Fl2x9r+3MhK4Jthca2
82Gu2fmnAjh/S59yKeaDir3Txc5jc+6KNSamRuat26DSNEzOJfn1q2aYUFQQ
CmQ5k/0Cxf3tcNrar6QJDHws32rVE3+vCSIX0fE7YnhQuvor+EO6u7bsZXWt
vCsZ0AdAzBcYhZ8AgFHejD5kMYKKqSQlhsm7EPwITDHNg3np5e+xbelIJ3py
VBSOfYE0uOhHu5o95f8WYbYyqLtSRA3FXlXJICio2S++nhpaEQ34OaZ37Z8L
vQp7vBEyDawpGMCxvc/5yqYMBRsoUgB61rxKgpxlTm32auz/FZLhUHq3+z+G
MAPmhovyakAmR5LeTjKFnXgJLIrutgBp2HsKxIhX9ln+v5oLmaY/UtC6qe0y
rUSbMOoaJrE+EcVX3oKXTyY18Frijtkb7Xa3qFd6vnaZMfbb1FB+kHy6dyvl
rNvRJop+hGsYt67kpiDhwJEAu7n7hmhOnnFIs4KIBWenHzQHUqVG/5orq7+/
Ie4alMr/7Vg82NJHnWE3tExnLB44f+ss158tdPWDqmHS+IGLr0izA2t0qYoK
+KA7g1f06fR/0Gt1jlj7ukn/FYC/z1P6iIm9ueH4Rs2eNM1hR3KDrYN/c3GE
u1sAAqZrS+30dLcguAg+eo2a6dlLbx0nC1XO2FNFNEqp+kLNfPSYjRJLGGe/
Gc/vE7/Bm3CW218ZgzlyhMVCPcOBm7Az0gQDWScZsBUwa8rVnFMJSK0TpwET
yqbrjDq3UNeIBclFZYyc01TQLKie0u2piK5aCS0y3ReQk8zSgfti+DM5S4Ch
bRJGSGUagFvgHTldq/crh32zMbgqPfDBoNSSWFUcUvXdgafXsRFOE+Uejroj
rnZopQDkkz/HN16pliA0+8b17DxDTvF/qz6l4SgkbJlB0nJCD0V/Dv+BSxzW
q9B/GoqFpsBfa5ukLrsWlc9PbjnOOKfRo7joravSvqnHMVbospGrUXIycuDW
aEgZ64BHaD4OzcFCAq8Pkld6YFtN9nhRhf2LOSLrJh7AqCJOpEAj/FKqps9D
KFjq0NA0bMGjS8Ca99UI+0r2w1ay5PQY8kNeqJ1bK6wSsdNzLibuTJdV/FmB
tKV7WPIcWcihBrTDWipElkE3QC26ILMTtBW2rpQxly04oqxioPDnKWrhXowH
6xpN5TmDqf+b8F3+vqpctGRT2M82Is1Y+VvRDqm73phpR7lk1/D9bAv2EPBM
2UPiuRhXX0lGf6rpCUIXqzPLxGlC74mV3LYGDy9X4e/N6koF53t4/jCBQMHJ
DRHJzYIHx2rt4B38RVqaDfeSCPR9UWUkaxs35iNv9z+vZSAzbaUcmi4jgT5p
5qPH4CmyRhvP2Wd4OZDp/VoYJkRVsuO3EvsLVgeHvqhEop05xq8VDeJaeaHQ
zEJZeCg4JHsBgmQ3fEkTJ8TudyrOprvyuSQwg0Jk04YxkVKy/bkpEL7prfmu
xiDHuwoptCsXKelh2jZ10Rh3OI6pSZOl9Cg28iwkQPgxXqeLcUP6WevurxPk
BRWnj6cvM6VuPjRlIX+gkuEci+wAiznF9OODblKo+7VOodVtrFnvjIpvsuOO
j/OEOwaRGK0rG6YlqBQQY9EyocIg9EnY4nKicD0dY/TwhePg2xV5no00G4ng
OAUWn96KJlKptHvJhmpcBGK2h16HcdchgKx7FG4gcVQk7yAfj2I+ZjbVzYPV
UZggHTDs74al0wlx7wFbXvSTJYHyY0Wqi1jz6QzQS1Zm4++la0Kx6cbjpuZK
k+1uqSNlJvdd4kA0g0jOTnF34ESGy55mB0AF5kH7Vo4Y0xUqdpO6Tu3D3aio
6Uh947m9n6ZogKs3xtSFGIfgBFEro7EsQhmYJ427br8otijntHecURyXvc4k
a6y5nDdQGiBZoFcroobPGeTrUTHs+MvxQrYfxZuXM6iE08lqDVA5rI5/RWgx
nTnVFfgVpq3mZYXypIAb4OyWfrtDIN6e/bzZagx0bYoCzm/hq4IcBhq3GGsl
3/wbM2IRC2Y2+3MCkRBtBOapPYU171B+J+CVjhauEj8hlcUKPvuGZuZwpowJ
+C9YArMuLbq6bFvVMMu/9EgERfIkvEaatRy0+MTzllfyquFHnMkvcKKNiF/7
xZ343wJx0OJz/f4PJErzB6Y63GDrdJRT1YVfEZ8KXlhWrCHvjkTS4hD1JewV
oLFipALtw3YcV1iBZ4I4hWrnCF6auW/aZGNbmEOvSLdLzqa6pc4Hr8sbAWD9
jpZ9cS2kb53IzEWd4BSo3Ms5fscn+kqT/s+hOfa8xfZGFo/aLwNXQbq2AaNW
4qLyWQaVlQVTdqIis3ydlq5RF2DPjNEFgH1eEEACUFuUme15f6W200DjSk9U
o2PssuINpMEUxtOO2Cvx56QU2nrKAYURgTlH/xJmbr/lSGFiv306iX2pyp9+
uoHkt/lHjPHl97X41jxTpmpOuN31LdynyRUAdd+7UlI+HxBywd7ViYpzVKC0
ArXakWofkjtwNPLRZFIZa30ucodlNUzMLY5cp1LZYiJVKECZagCzSUde0lu8
w13KJ3fJ3560q1WhjiZpKS+lKXwTqXK5OHzIvRWf0UzAGrEV6ZYXRAUmUzZ+
XBBj+EyOBcnVhc8Ka6xr85+AIk/02DTUrY8pZPffLLQdo9FVkOcSHWpcpfgA
6vQuerkxVhzE6zsrMUBGAHnuCBO56dwCClBPbuwvr5+z/8Q3VGkUj4ysTtOx
YOEursO3G6jpdpZTHWFhIlyK9jtfaoO8GsYITjvFiHjqAZTmyKiEcb4VZsas
+XHInQK3ddEFJNg2mrpGVbG8erFaYDk6ZauDvQfeavtTQKd5bUvBL+K89Gl1
evA6tpQ5u2aG3v+Cdn2L/SOVXsEhfuMCLg+4yBGHYdemcDn5EGd3Ij7f8Jtw
Q8aDfGQH6ZiEal5Q4pX8YyvmktvV1jooDqc+MdhlSMQMalkQcrRM1rtwnlUg
uVnIZN5BlAyEW0UCDFJqxdGGlHsUsG2eNTXLJGrJIlIizZEFb0OVQf+2IQzx
5s2C7RV5A6e1K3NvxKzqOhp6R4w14OAPDMx6tfBfW8koIQuGco1em4W7uQ2I
Fvv53ViJbfH7g+ltynk81QUSEeNwGk9XaTgSrUYvkFX78IDDOtYL+eC/w4L2
WqLRzXqDisz+3IzpvPv1X/y5J4O7xOcqJ2phUzDeYcVEarKG3MK07+bJKp8+
rjvm4IcrqPEQKIb7n3c2FCgLFxqEZFe3BHJ43AFaMpgr5kYxAL2jhqeY3eMu
/Mdzdw86dPcQtURRwE/MpAgKhRcZLYi4/cVG1noO72eAekNkoX+iJUKiTBpF
B6yjUb1SYSEBqr/Gj5guJSPFxNjCA6ACeDNZUAVDaQBnpa2xT/90rcTuuZve
quA6Wv11QxQFOe1AFcE5VRW2EWShKwpUcaciMrM4ekwOVsxX68hzYXzYtxJb
9K18jFte8JKNTsEQvfOhDZayMsyl1ixjfeK7qwNOm/MLli5mrsNojBXBW0Tx
san7/gCUkJ0vKWUIt510pu/GRpheZowGLpSRqtbEIYJab7qwV23+eEN09GxZ
Wimx/oymVoOKQvAQ69IMueh9/p1wVmZ6wNjCCMeNhXOlUDzDybKdH+uCTPnq
kK9CYAoLpuYgUs3V+fi2IU+ppot2pA4kaFNsFA6A2D0yy97U3ifak1I7fWvI
m+CZQTKYjK6wJg0CfHJ22mLshmqgRZyRwg3bFc1QtX943DgxLpbCzmXg2xxc
jTYbdZkd5oduwdohCns4Fz1zoDpvmnYwJo0sGgRA4ybdYjjM3eQkKcvypCGX
ZWbfgguomx0558wZQRN3Cn1HVtFImkq661ApmGYYimF/NHZZHgsxamaSQ8mI
Y3wOjD0H9A21jFr33s7bpd3faDhQqM52UpCkr/nYeP/qnDIoZ844ynAdMIRt
dOnQOaiXc2DBtyvKKc+0/VxWXhcWxfq+1cjL9JbKGGRMbFzmGCo8NcAwCTZO
WcBfRj4GuebiNP7Uz48U0URoIvDAbwfaXTev7shX3ujE3d6wfr5FGy4UecPf
pM58JT31lCytI8zbfd/9VWIGqOEgGX3lv+Rzd4gCLPvS6YGD2cB2AUmgKTw3
6OEOolId3ej7J5ugdPWeQLy4mr59VWdmfXZ2VZMo/PzEFvHcK+56FmmAyzxw
e3kkWEBaj+N+bujR+rIHN1j1w9ggzBn1o3+U6dj1jxkwhOUHEm9HyJGBiXPq
9rAY6EtOwBwbmVPNeIC3j0OSRpv3qr3z+Qa6Nqaetd8rNM6WSnZt1VI7s/w3
j8pEYrU5rrCxpcpoGl2nOeRm8dLJHsRx8Fvu/7wQsfTeXRPf0kVz7I9Rn1Cx
ZoFIyPL29/bx1jGmFuPU4k8DV/JHjgN1a4sXNiJ5bJrrnl6Z4bfdhmd7Tx4W
RRaV8v8gcvaXPbqCd9li7yLU+KG2PN1ZAPTbeoPDcvvAXiVw7c9tcTRcPCGN
jZwWqw2oBROycU7mJRczw7SF5elCDjVd5oP8W7sdWZ6F749h0IyAtNglVDK2
f+h6BE4oLmv5mvIQb7+oFkN3kGLcYvX2hBfmfc7xLBDWDA43TxcPsEMy3WnE
MsA3sJCNEJH2xPxPCr3ao7wEFPfVjMzmLiJ9IQplKmsiuPlhOsn7V2KRdag4
R4fZaUbnuKOUe5AhyCXXzgN80CbdN+dm8mXwhTh3PM1DI2MGnjzc3x9KajSZ
Otf1E85A1iDL4bA0abfGewDKWxtBghQRDnujh63qglz7OJ7E2GPF2ScFgPI4
0F5JFhH+NWGFW+0wYWm+jV3yelKlk9NChr+dSXFbCnKrCrgpc83EQxxGFtui
Yenws+8WWtR49ZG/UXqwywWfW+wxsrxgQZV5EqkHBIDuxgdJoPRI2ogDhe83
bR29aZvzxa/F4MwUnqrJ03d6Ifawv1uHSqmb3OLxM4D5CsXfEJhRGr7huttK
BI1HHs7Ml4jUIa/67xzgbj5mLlSBUBGq2Di4ShINI+IfjwgC6ye3Tfz5eNew
RjM/7q6ZQhEHvDUa7rpOgpr+bLUDXe+/R/sV+99f/7EiZw8sQR8AONoaS7WF
tZaC45M3FzMZV804cKcEAj3FnNSiqKpLd886eQ0YIBUyETnfYoYQMTLRWocY
+9f8NxiAJeCeZU3hlpMCW9tbthIPzb5pWWxUBXsI1B67bABFgiBLemD8Jc5x
A9osG9r9ZvMfzUdp2y2yuosAyrTa99PJLRTawlcju9Gy7lrYrvu79cKxsDN+
eP/3RLQ0zHU1d0gHmLZXnA3q69pp/cUBY7xkad8ZbNcbpJ6ueQYh/VhJJE3S
kdssXKGoeTNMcl3hoD8Od/0jGieF3hlqxxBpTdk4eBbEG9jRTtm8b2+Hu/o0
g9FZ6Ej9+NAMeOlpY13p7ZJ8OxSy4PS2nZLUp48+0F3eJJrK9ZHfDKL73CC4
Qz+H8J+OzAZP7A5PsHrQ8vgw+j/l0e7+GcjoG2wrpNe7dl9zqzSqjxJOrl8G
2QWh0AxNXAxzXnrRWwL2AlX2czvpaNPqHMjQb/P5Bu0wYPyx6fPTqd5gqOwD
QzxDkh2pKgWNVikrOEKnG4HGDNjx9gcpf2qckn84N2vXTts9BrTv4oHDLsMh
lwf97bNb7BlUZJ3B5bP8+UtVMoB0eGRlWDqVcQqnn6xOXPOxZPeUWhv9C4+g
FsTVU43QOh9JOpLGUYfZCEgus4I1KNY/hnGGvsAw7mqU74oGnHC35GogP8iH
deLQMYHa9cGy7mkZIuLXzM5v7pkMvWTcPIY8XwoMuNHD0N8dPJh/0hR5gO8k
eVC7iyZMrdBR5d8oF3GrMsPfo/q9/LMFPev3IwL4fg6/0BgEdujGTBjIvLq1
k4IgmcA6sV123rzTpEK369oe0sHILQMGBpOcvkCHAnjyatwMvrdIiaMJNJJ8
Bx93Rpy4yOvLRrGw6yyUFoVTy9iQt80DkNqCsTgsYSjHF1lP3vGfHHY11PZw
Wqt6CphK75e0Iky2ku0LOs/iykBFlnZRK/QbMs7FSPpACI9z0TUJsiykuPqm
Cr1Nf6oX6cjV4cu/tp4YLVGX5fI1U5jw044X8L5QhmcqpE3BE8ork1JN55OX
WLcE+vGi4hT9ldTRgAZREfXkiaxIvgaWogge+D1hyYjgI01NV+j9V1iJ5i/c
Nf05JCYZT90dEhB++ip7Svht2o85OPPVrIXWf2w2VpoumYHvN6qxXO4I4ZNC
tg8Zu7tGgpF3pAzVy7PtRchP6ir9O1m8XkRAdICRCty9wpfAm2MfCHwOj9Cl
aWxIZcNEW1cLzTq0rIokVaVhfqn8SgXpXWK9iYfjQE9gJz7Vu24k+6eMCHIY
HfzK5ToB2R8r83W31F3I6ZlrunrdKCT6XunTUwJtz/ZPrNteTw/VN95XO/Ws
+gGDHHRLYB4RZFqjdaeP+3Y9evl8kfrlCkJfnZ17dd8+AkjTcmPB63t9GXJR
JCwibaHb3Kye6k72ngnRQ5/5t9GHsnCsR2GGx2JYlHkq3MM9TTlDQSNIOn9V
HaeEiSW340WbgdolAWmJyn1alue5/0LbUi9jPItAZMR9D4Mr4mYi0dLIPBH/
+UktEpbACDKmfMF1c3HpAHA16odDdGer/E8XeF2oe65zkPRdd2uovJgqcPL7
G7OkqtrrrBXoqZyMXPJEdLaHqsu9E29bKjnr0tfi0KC6eE5mdMffrywXC/YU
E0alPJcqaYNM0yKhTbAxIB2oxJqVnaEcJoJVT2I2DhqU1m/L4dvLmlSVBd3p
cpFzIAlbXg1El4EInT6WHp4MNklEFEdE7mK3cqSqgs/H9bjSj3Y1OrvF6B0B
P3l/IsyN7DgY0qpWbvhUIa8jNWzqdfS6umBl9YWz/svGB9dad8+9gGbMprGU
6yGfuLXibfIYL07/6BwdPBC4Dfc0kiG97DHC1sOr3/gjrk5dI7Bzrm9tgQQR
jUjjr3wuwwvh46KcnuKaDdDMyK+aEiKPvRppvc39d2lvsfpHhrP7B9/9FEsD
vPFGLkbHvNbtHLoT4yBzTwsJVZWZ/G9HI5yfPPeH+Z7QN2vSU/lvPcSE1L9c
JboBJ+6Bir7Va0f/m07TWeqzJzRmf3MUQ4aiVYZv88byooe+NHLncNBrXepE
esWMb468wllif77RqGPs+06HTRSsZZF50MkmMT0+UQcisB2sMs6jmh5suGQv
12NLOSb4EWUGbryzgy+QRzyTuFzWRdSYaNAqvDL0al7FWbpTvTIaR9qFURAl
m92bKgD/RUNUZ3IYdAh3e4tJ0jHLJSA2Qghe/P3yLpI375izUMjd9s0eqdDd
rmZ+Oejh3G9uFYNtQpTG0ShvGVToEh7bLTUiBCv3bTCMtwdM27/blhE+9RH7
0tImgfS8Nlx+0ue0fnMM1K/KcS3ANv4DGdAbpDvr9XrYjLuxKnqegUeVuMr4
+PXqYDxYgtkyWPPL0mvG3W5wi8ETClqErZnsRD+VQ3CmNQFNcZcwU8NfPhst
mnvOmbaYolYjTvno43yX8MC6PDy0qiVsL0k1ujfX5TnXKHlRrEg653Qt2dco
4Vp4uw52lysd5WLC+UF+gx4fbF7wc2dVT5n/FAWA8DgSLpPlcOydDSMGe8+3
2XoCn64pvIQScYzDwZ+YMf9QfC2eXxU7d9Pn3bpuMU2dRXtzMWQiYe1kPP3n
Pt3vD6ba3uZeb78pynVbwO6/5n74V5e0G/oav/ryQNtv3NfdLqLyd7iYpV0m
bAvo1Za3YDL7aM1veI4bxfxH1n4vbsHYMkFFAaXrkU1fS1aWzYWS9LPaxgWu
+qTR9Fl9w945Vy28UNSVMySW0B8Y12UhqXZLB2rrVn/bHV7OKHZblOai1Ubu
CsWPnyu7i87Hk7r2YCfniLgIWcfwkOrE2zYYU+9LbJTk9XFCSWtmzTo9mvb+
ZFQLqV12t0YOAhi994KjMOtgPdh1A3MelILm2pIpAeall+thvRdPm7RTJrS2
E1mVYpyMlV/sUra3O3oLw9MyyBgIHrWTHFrfs4h+zuBQVFkn0QUOPFkEaI/T
NOIKpsj9L5abAgZekXbU/sV3/wEk/fxttzPWVAlE6sBMFDN26G4wiJjq8BdZ
FCRodX5bJdTWkmXV1fZo0IqDuEKfqCfUNUTPdDGq+nptHV+Ahh4SW0mbYGG2
1t0lRogXUUaPL8kOeF0qUtVBPLq8FISZk7Xr66+TLCzwQQu6HQSa9T/YmO+t
JKBnOx+0RX0ppvBRrppH/zJ3vbQIeumZEjwSFsAbNbb5JCyREFVxyvzZFmjy
In5V3+BWKaAw6+0c8eJDzEYnY2KWVEjKLumD2TOEV3Vj5+jYhJBpZiNfwKGD
JOBsdv2cVVwcqDM/TmvRrJuPoMQ7bB5SbmzuGf5cY1ZOX5xQdTbbolcEV9+Z
WkpE1leIQBqz566t+qwuDMoXbeSZohSaxyzpdLuDixcFlzwT+J8120RkT+39
/Ru/MriKlHDX7QvmVVWCvVRJQJNPVSxP+IDhMakAzmhc2TyKRrv7WMZeY8Us
j1OHfr7bXA4RN7Eaz61yJOfPswCU6zuPCpdkgfKO++ijjAkFLXPLCLjqKsFV
/G9n5m4mW1YBjia2551VleLLAUE+pPHhZmkHz6nXmyJgSoZVwwIEPeGQT0RG
+eJ7IWjPiMRmqAo/TWbAe2/KqX25lsLWgfX6TTcLQirWbCoPyoPIO+Qdqp8A
MOUiONdeDEdHpK6o5QaTU/uK5Qaj+rHFvUHEs9b3P6o1aiFtDnnayP8Ul9DE
mfknZelNI0AWWSQ9+HhmQ4jMzT0xO92ngypoZvdgW18YYCSzSUfecnrlrEar
6Nsongp5Q0osKzT39tGHIpvZMAZnzFNSsm+Dghw0gOe62t/6Q7wkycGP/dbd
kj77ZkhnPj8R7p7Hd+onW0ato5EH8VcD6BQNNgY+DZEZDfWXt0A3kXgXeYF3
npcXa69CK6cbPBPkYcxhtMKLrtv3xY/9oAufMHtPHWTu1/uW2NC7JJpZuHeQ
N1wFohWHOuNKlIGUBsojXjoGHuBdMnQR6Y+Xm7KbWuISpPz1GT/Fq1PMywbD
S6tOatyOO9MC1IDs+Zogx2zBUP6NJw3AK45F+zw/fbiuOIPoAuQ2Vh6wC99k
nJndMwXbNZUAZY0ixqSLXNLa611Iur7RTS8WRxvrWTG3DErrGdzXqt+bsoag
wBrMSObfUSF9nuGjAUAtIlpDL1VAMPbcOkNesLtvsdhJlbz24XJM7Itysi6e
86EUhVRtrNr6jMOwEYMfP2YCWry6HyMAnx8KB04ww7O4K/fXrLmjzwjUVJ2S
bgvT2tDMV8kzR2FN0ocWBgSo/76n9evhGO3miU+q2MOW2XhVPSDXWi735WH9
EixOCi6UCkE+Zhc7+q7h3jjEO355mJZ0arfyzaYVzMgRMejPNkN3AIvYt2eg
umc+p+yd7gFSxnq/weUavp3l1mLVV1jZ4aC5fP1e5NsA2Wa4ECaTAyWJOr+s
L51y88O5zlG+/ZbY1C00mSNJWpytnho8xKdLFJBh+RWL9AFdfKTShwjZx3UV
RVnNBPGrXLyYVWJZG0EKfvC1q5o7WMBMaXrdzsQ5m/XsbkI3WqILcHyUz3zl
1k4Fd7FuVy2fCiPSiqkyG5S9uIO5+JBhCquBthTn9+ZD8noq3mGWWPqTZ21E
3DRsAMK7609ksLvbJYwYohfoAPxvCPgIsiVlFysUZ9AEQGics5dfNGs0TFa4
C2pQTMiGUWNJDgPs87TDrceB3nAXTFnhMuMp9o4OQ54pBEFGOoYSSo3t+3Ej
PSXs+Z7KPlgWuZ0CLrT96ybfUlc4c6UNR2CrwTZQ4xkSA/AHQ2LYxB7kRxT4
QBqDCfFV3QBY04x9I32rNZKGgGhmrXNjx+MrmYpWxZ2XyZeSTs19FR/wy0Qh
I7b8V5/thYOFBGTswaCr0Qoqzst4mEoRaUkA3GK5hlbRWBa8NMKmggY3rgTY
ZsiuUH+mzJBOWdvVueGpf3mHn772tUNFr+Cwlcrm6qeFOmV7OcNkJX2AeQRw
LCnNr53Vt3lVuaQUtMQXQaHvkdy5xtgnqK8KZna9IMdaHPUay3n9yO2bjsmI
kFLKNeg8tPevHQtZWgZuXF3fwRtIaus0oVlXpr8Iw/y0pb1QWYbgKWRXxv8d
PCILFkjnM4xGpgxqUAce8/A+AUOAsAhB1uLmBiA+B+yZLycHd7okE37wxeQv
+IhsHFrImqOyb3lCRlRFcY+XgHmy8H/Ggv+aEAdmI8OAZU8rJTSrETqo0q9v
o135Rn5sRDJ+mRE8U35tFnIduYlmqqUXwxtFCzjEA/9FOFQiSA5ei1NFu9Ab
P39fRPewIzwG7g/Rdwa1aY6gU+vQ1j6DxlWk+uXEFe/LS9pYT49UvAY2yTxL
oCoFLm/sCYkafdiRnEplo1oj8Y/gDc/IEIWhZmJi/2G51Tq02ZIhywEUJ1Ga
8anSrW9q4MuDBKJKeSS08m56cSbKZ9XTZ3y07ouF7yVGHksuuCtmb5rHR8fp
TW3VZ58FJUN4Q54vwjPmcaojvajQZUQIxu/cVKOvKwsiHGq7X/h8o/dZNmz2
n+oyZajqX25gt/a0USQ0+QmlUkAzUeLDq2/xYN+PLK6sKL6uBQ7ZbpxYUZnM
U/7PNewuPiVdb0WbZ3W10xNtFUQZwpwaFXWMEtt+ABrpX5J9FJC1c/aimdZF
9QrtslYYihsrSIjjwvFZsRccW73803W7uVSkvMwftj+dFMcRGkCPnqU0U/Ut
I+JPYH/uiUVlcCpqztF3CU5YraYMhz7a2z3Kz/f8Y22WZrDJKxhppF8bKdMZ
7W5ri+1HI28pDz2BtgCLeEpD6Z0Zcc6zNqyrpYppFARDwKxzWe4Lgy8PqGI5
gumfx7cPEPTjsyoPZikJhstyaVd5YbF8Enav2mfK+6EvLECyuwO3e1D+Lj2b
7c8PdpTeI8nPxo4ujzcFOWWQXRmJ0paoOHRa/DO8uVpMWbWd84Be05m5FKLw
EEpliXsVpKgQtT6Yaz9d1ARhgYIS/p0a76q///eLi9JolAVUsbtu8RoJjSqK
YvG27OMVUtERfFx9D2DxVhOpZ8Ttx8zeS3NeEL86W3IdMyNU/IqNUkFFBHLq
3XF9rzSQgTVvwwZmbJ8QJxmY5b4vK188xPOtcxujehrTy7oXWRWr3TF2y7sO
rS4VNF8AaiSSt3JPiOM/nZXe3HruS5WjOMP9LgRNrWtslMIhwdqnLJFoQQtf
yZEt6UpW7WYOE4IonRHjj/4XvGdBNqkEPmlgqm543KqxcUWT1QhE2bbLSIgq
s3K0jm+/xxkWjFGAz5Dnspz3whhC268wLXP0N6VFUKXcLhwu/sRg9LKlXpZf
Tw/60XxG26zLdXy9ujjHK5ltFoFcfVeDprwfODrqW0Ew/lim7SnU19j80Nfu
XfZS3scC8Q0cP+DOtfzK7a/uV7g6HJGqzlHgSCbtkSuA1bqk1XhE2EjwYbVM
iejyV9JvFyKOoLSPRZuyvjutpSimSo8seaaAlcZm2hQwgXaVm4TzlCf7TeEA
+vrvATLf0jfIVKvnrBtp72DQBob1x4ePzJXAZFdDNVTyty+Nv4ZrDwxQN7U+
g6Fe+rgpRp0vWyc0V0UqyYcfYhnnPKSdPaDUjed8HyytRSWYr0VO15J1XjIr
SeJNwa5gfJfSuOVXNk02wc3QoPtN13VfJn8NIH0JzAvtrEQuHT8K57NjI+J6
zIgAhdKXAVjLJrmOzbEoP9gPHBTiKdty9uPPOjJ2DwJj1QXlR6Fa2w8CWPEQ
s9bhcN+e8YYMJabtvlydOfXbf6KOkRJhml6OxanKerTpsLHBFUUv8UDkAfNU
J69rk9+CxV5Rr3SOrWSAaweZa47iqr/ODuq4JO330x0/uakZ/ahNWDkf4tew
68t8YfrKv52ad8zVWy5ZIBYpVkpdmOosj0UTVLQxO4PiLcSm2hNe0oY5vxaH
+Obfp72lZ1L5ipBp58idkKrzYS7+Jv0Pa3trgipl9LBFNhJbqTrHbSxSM4de
qejmbYPBvxBiAXxfe5YUF4Y4ZsBZnm9elypyW5+yNoVrT+xVGo7ZCFONUt73
wLyWy7cvtD7Hosk2TkYGZ4SOan88bn7TzxTdHfiDDGJLGs58FN75S/4B/1Z/
HZWFSDYbaGPrczmZ0v3PzIK0p/lOwzMxKbm+50rCno/bQ4nZ2Kd3yt3MUqqM
3uMulSjy9E3Z5ZZjmbMx5BFc5mu9MlnaLJSwYfjQJrVYM96D0cX06iLS3Bki
R9cIJgF6awNUC67MMVK9izOzOPYo3He0W/PpSIBNGn6+AAxGAAGKgGbOq8AJ
R6zuPt2vKaSMqUfaIxXOMFoE6dz2A16qwBKgJzE5+H/JFoOVSP+7LJP1JSru
7enxDderb15le+fVOHman74IWifyzZITnQp66N2+P5LYkAJOvLWUw3J9OSYK
LbdW3dX/P07JDnsN8uTDpyYQUEOs2bZELl3rephiMSUhXLS9FPlbD7zqQ9sF
IIyGxLcQvlQB+6sKsDtlxDPVuUi2WtRyo5k6x0SrJ/9Jknzpu5oQd/xr4X2C
YqSbEKexe1t4i1m/qkLlaueQVAW2FCOnN3l+r2chXh7JlTCJKdQH0QZFnzVC
mbV+ZJgt2Caj7Ej9EVestaDZlFdg1ovFaEDuP//QX8lWnshtykFBQjE4BMou
GZfFEU8iVWQh7Bjd+juSrpdLeEmKTIHkGGUx8sgjKEfnAw/Wl/XDFmRqjFnX
+fTrL7fvstV3nEz3TXUyqwl6rHbGD4B3p6mFbR6im1h4OC3+mgSthYrpQUqI
JTxyOYGnYlqMnM4TnGpAJstoNxA6vPU9540aQ8N42aRi7/EqO/7SsOMNl3cs
zdZU2GtvPTiG/0pInmnThqA0SFiFCbVRSxoZx7WQmfyOyWwHfqZ7P6/W3eJL
mAuhrbQejVTuskDdQVo1ood/y4xVwv+7db2DBflYxsaOsADjH4eADflBmGu4
ZPdFd4L2QS9wXe+Xib691Iggul43Od8t3KcMrqmpXZxGrBeeeaTm138zmjpo
87yfZMuLJ0FpyrI5Xq4SdawcwVwmGxYZIcHPxi8uBhrUsTdai9rfMG1UsNPr
rN3h3LpeBbefgI7LC3n3pEblCZxvh5GS1dp50KAoa7Du1NpCkfx4FtDi0Fko
KqXxb5Ko0uE1Pl0227t+4/s2m2KT6EPCfY76Nf7YsAbDslPJXpItftSyORw1
Tj1GF93EDsJDLIb3H2BwTZ3uZvdH4mLcZUst46G4dxkI5OUklEEnC949jz8W
6onJVTDLMsS0kX1lZNQJJSNnQAVCPrfsAf5ZDwHPpTC4mQf/ILVkpNltUaa0
xPYgM825DLFGQkbBDgd6c9ONQuga9qAjsg/VTrUVMQA5dNpMSi7eElyi9IJM
HFg9KsYUtadgFokK5txH2gNdbh5P56m/qToMsX4RasaAy90m9MU2c0aAmgFj
1Aafc7nIpMCt3VYUHowhX2vCJ/325t6M58iBO9arfspd36B29OBqFQbOhN6U
4l7NACD4Bunjc/btpmdVs3CmcBaZZbpU9vfHDntWEU/RAJW7Ekm1Mxn2nkZs
6BFqOovsrFeJ3N/czHQbr0mUuqR+4k99BvYLQJgYJ4pFHbrCe1wdldFQNfft
RuVhqtjhcq+le5bdRgxf4Z9INKJe3aB66ldYMsbn84z2TLJnugVzJDj2UaGS
SAuWP518XQSyFuOR6C6Al3gDZ+F/XY+PlhePK0dWcjUgYTqjBvX8SUM/gqwT
RhAXipTspUAX9FqmoJwq/G29sPzTZMu5ResdjNkDmTp1fGF9xHytkJtNHf8s
+MSe+JsjmyBJsXUcOfhtrAteuhwQKbqq81RCddUNQuEdSrO9M8YMnTPIfSW7
vrwm5m+PttqHaBPpkqVt6PoD57EwBggP1uuZzQ+NNeorrDJcvcS+3s41pJYz
u5LUxiYUa6rf9qpTb6ESCHKNthwf81WZB8gQnF9O5hKRvv7gzOj/CejP07Y/
AsZVkPna2M80nq9pOW7YyvxQomRkZXELtQBO9KQUuJN4j6xEbahs0zv8DxDu
4Quy5nQ1Fe8Nl2RTiqgkiKGcNL+FE8TjNXp2IiqiWzidpV/2R6ynmPnu41Il
SUfCiWFNq+3xlkiQZLXQ1uLOkboJlMEzV9hHMNXBPwQQlxxkboh29bJg0+gp
1K65HNMMDls5oHSMydYTN8kqsRrTPk1kERmU3DY9EmQLs6v1gFn0amLngM/x
4LiijTDvx4W8GvZgWUPpbuLnyVJtcy5e+CzeE2prhBz81PrOfs6Wwjhmx+9S
GTA0zmh5SG9zpVbVE+T66UpQBTlLx13HLj1CGHSaa+I2F8kxPLf+3dI7wRqJ
XOY7PnzVpyww+c11r/MMJg2TFNHPdUiF0XoFeMDbzfiycK9c/nhkRnBJHmaz
6SojfLWc/BoZ5p7M9ZKW9z3T1lVAySJGmoBfBQPnsaSnNSJ05NlCThFZ5oaU
AzKqCvjsavnXU1t4Qpp5XPPc7FLvf9c/UQP4nF6UdCPH2PIy31dA2YYIBhL8
JHVl+FQ0wn2Z7wdRCYaNu6QzNvLs8EPsE2hBr2pKIwaez87aAWamIGWvHUd8
zPTOAr3uHWFXBzGXzmPms3eUICjlA10pI6Rq7ZVFL5fFrezVvLqq3Mq5F6i5
frM0wI9fDlsdvQjB8/U4BQVLtKSVK8KP0b14fRMLwj4hny8BCBE/KWAs1GN4
2ss6p43edUipgbTTfVjCCAMCHKClJU3E2VxLwT9vTfVTJpcPzGUa1QfSFXd9
hz6Yr6sFC0Y1+UM5ebEyMO2Rg8NQ225aaK65laUYoydI27G/Vy+NAUa6rqnI
vAvr7Nv7LC/mBlnF3Jg8q/LFDSm/YLspHjv+cPNjhwHO2Zbqt4D+wfshw8rj
jAgreSbduxB3bnLQZlfICGEDUnH4kwb+jHiLsVfid7Zvssjm4LZQ+VINmwWH
IlKRuN65ohO5squHGVqFpcLaVr+wZoiuN3Z4HNPDkHjaxb2LFi9JqoS1bCuC
Mqu3wk2qnZzwOCHD6NxA1U/xCDnQ6gqebKexBFbkRm6jvLmfbTdAqb7x8QJX
fIKzdo0zlGXGv2z721v25lT8fyXhZ/gZpToRPTE7EB7fMrf6c3FW7IOI7rJX
1vlCx6ardX+Ly36xaGeUsTXhQqEKSOXjCcCVn+x/Ng+Lc+baNqAJ7WYbOvn0
a4BvRRDbS6JmdOejTVzhRZiXbVpjm78EeR7TY+F57tp8XTuOfu9sSn1u11AT
0zRrlA8jScwOcchpYes4R1svseDYPOh3SmWQgnGZ+GvZFbiyQaaiugr+BCPb
+iUjnSXqDzv6h8HBobCHx+QS0e8DW5o8v5Ek+e1xf5o/Toi9uBaTwA3/PNAL
bO7Lwo1nhMYC+EYxRRXxy2xzDj5wECNVaaAL7Xhn+xBKgdaxJ320QJEe1y/U
auKuu3Mg3SutAhq6OjfkvOcT4cR/XOAVkYys4YyCmovNSchIgHoJ3iTHGiTu
ppYVtbsGcdtj8xVBjZMpRuOw9N7zTV2JJKzQLt+FXscws9gFpKfuazrmt2nW
eMbgohflhN2NUP+2q4U3c38I1c0skLiB6AOqww7NDOmDozOz/hYlQmWuUVdl
tIW6WIdpU+wN32axoXKmJLrg9vjyijkOBzr8mKE4X3pNF4YtSUlia9NeGLtI
7TgXlLpnRrjLHdYh1zyXIPGrGD2yz4iMOjGcf+WSHy7Y9lRzSwqVWBpT8a1c
nbPszew78OrjuBHki6LVK12tRDtqIRrjAFcS8e799YAj5jQKhuJfI//q89VR
i8qAUXdRzzE24SGkm3l8VfcHYjqSD1jSogsoqPgoBdcW+tM56b/JNmLOL3u2
b6osDEtwDx3DzGRt70L3GeoxWfFEY9aDg5nb6zkQld+huHZmETCauZ6ne8Jh
olif74S7XeiWyZhO3j020xcJ17Fz2yWTAsxeS/m06W12B+INHRKGPiCuUlwQ
lQToX0EpSD0pOlbvyZ5XPxN4yQei/f328ygqp+jbjym4hkTGvcTqtebNXlL5
vI3ZBrWRAQgYoqJmi04WQ6RkSwIlM3/i/QlILKHDWVh5mEgWgKqMO8bJrVuC
R6Piw2ayau39Bmwc3HMcEWjOPNSqJM+1gPXXlZmiBhhlvDHyPsF7q3MgrAUA
RwPd6Jauwzcn3UdVslImbi+Ck7J0p7vCfZDtU1C4IsP7JyvtBw1YzlbbE2qb
qVRrvW+fdAjiRyfZiWDi7Nvs0UBAZu33Y4TRNziCZ9mcIMQj5faDf2oyT23P
N2fQEv5XSQSvMkwZ326J7JbrVW+sOebTB5OiC/Owyi1sp61uZ6oHsmiolwsb
FCsVu4GhXB9u7zqz4flTY1ZovNTcVDJnnJ+pomHV2J+tV6xjN0J8OdncF/gc
dETYv9DLKsBCzWEgjHQm/7e9iXnzWN7rNMsQGOTCXSKRgBK0kmnZCHAqxC07
G6XkmnLv4B9H0wgCjENgQdeFlOBE2Kn7hKD5fxSo6mwoU5zyxzk5rbtzuFht
YOFWgYKYK4/ZUqkuwyXqFgNpDVwFfwtQCokxlExGJx4gqJguwTijnp3EbCXq
ixLBvXWzbbTjEwK/sJnXF9arbZMoMgxqUI1TDt/JdEWdgJTZRPsmWlr+wVnP
9LS5ePYfQljCNL66GSliuTrj2Trd+jk9wufOKUoSO0CNVWwp54fAwcEdXm7x
0S9qLa2XACMIVt0aCceHF1crE+7J0XH2DeCJqosSBE8rsDc8qAuJuw3R/y7V
u+M3xAmLegh7ZE1U/ywRNECJuqqa7wg0BL63Ez5LrzQNRSmIr1mi7jT2LrfH
4vVdvPdOHjaq8U1Bkok8JamXLak4fM6dG3hxzRaedhzIyxjlOlggVmR/poHv
zLM03A2o0qz+g7hzM14fKma+TQkB9ANDgijJPBO5HXSnHcRQNU40A7if0pvN
2dqnpExVF/HlCbSPRj8jAAS4SDvZ6pDAdbi7lElEfYVu3AmmfKPIuXf/zH4j
drpU5oGgdsw7WeSt6HcYC1PbmBnzF1zM9JZZ6PphsrCo0ZYX1rPWMin5XK4q
I139fQN4OdW6PqLrYjke2dLpgWlFm0c/tSNdtSLY7WZXbrSB+Ac7rKY2DDa1
6prZSoUMK3aDZh2ooxDlsZLq++VTtdLRNYCh1BvI8n5cY1zuqBgUJk30IWxI
/4jr9LojQmwQ6nC1YAqr5RQXiTcVy62AMkBe3Y9qQhj0Hcyoudj2kozMH476
ZgYBUeMXDNeQuva0RjeAf/5tUoiTLenQwoDqBHkWeqVdiOrkU5/7DovM6+Ph
hGUP+YNDm7uslbMV8UdDPbnOp1QXnkjZ0U8zOsdGvePJGSrd8ujXK4bt75Oz
ZcyfvoPuIeqhNUjSubgJVmtMI0NBoD5NS2PoezYMfN+kF1piooLrZ6P4zsvW
8VyweT8T+kkpMT80b9c9XCQYA9papN5wRvehJrCm4Yo5WTVOu6Te+Dwv30Ax
UosSOmqrfDS/MVtSrNv2XmZ8WkOlzcl9H02r/ehzMgaDUlWWZTDcpDtKIXF2
/Zzvy5hZHH8WDGc6ofpEJ/I5Ir1+/gfnqMZ8LCKRPVQaytmiIKtSHfof+AkS
HCaIMnkATyV+zBsnEgpW93bnPgPqVjeJDcmoBWvvrDK3zniRJSY8N3ZGyiTt
+y0rHqO8rtXg9UdfBPzlyTRCRNfVztAs2EHQCOayFhcVJWtcXlEStb6xeguW
9zYbwAqCC6xF/o9IgyaPacgK0i/jsJ2RfFIIog1heAfMDp4kzSikGbT8NP0w
cRNBGdvpqJRz6FDWtr5+pdSxigxtTWlxnAwW+7YDKiOYtjPNJjgCQDiT3p9S
Ba39qd6HAsA0H3bbktL1O7axbRt5OVWurr/yqwo0bWs+9mAPsc8aY0Zyt8jw
4vaS9yuLd1Fh9GbDwqs0a/U8VnS9b1VNS5xn3G8c9H272Rl130GMxC+jm+O6
YKLYAIxTizJ+YEdeSPgUFN6uvgdnXtH7YqIJi7slawCo6biL0Kw5DaYjZ0/w
fcjnqo+ACTTPRc5oguR7tDbIBtDtgvaVbnn/AguKP0DUBndXx5aMXsGQid+a
o/kKJe3X0er+KXsPdyh8k2bbmtbThWvU9VmMyxDXVsy+cxuXSTpDd4gTiFg7
Bcds5NLXiiyF43F4a1Fhrma6HAbcxI42kvOpTHz1WCWUsEduDMSyY0ScA24g
rpRPdkUUBq8lTSL4C2+ABRe47lTKTxzuKFzchXD6y2/rQ2dCZ2AMYxjWauvm
/Qc8EnCMSN6VjNu4JISboeflEaixplq21I4H2CmS/9/PaPPHJmqSV26PCTXg
ry2hVaiiC7VyfMCD1tMCQ27d8EUIX56eQHLGd45oTPq1INI9erR4QWbL8z0w
EzwD/nmAjO1FsX3cI4Q7HVXrD3apn9vDCXlj8DlxE9H3sTuAQfCbJRVMF2p9
g0YgLGLsP63JADn+QHOQtcz2HD+vMhyK35/ybA0TrEKWgpDrBT9lf0tDCXtv
H9ssqJfpXb4Qg0f65njnkRiPL7T3ljaIBw21p5uu+/2c8Am6Be6BspeyEl4L
j6Skb4tgDeXYEOlVZwfp2XRjZ20qyh1lIq2JrOsEI+v7MHHuv9tJm0kLiBhB
ImyPX/0TU2QbizAwnajNlne0JVOsXrgfX8EpLc+fiEM+hsm/Xizh6Uhb9p7r
0kPGjI/1gbC5UULtxw0NPcy4/16kilJx7YExSFdHWNng0jSOoTlzPtn2em7G
UMwLUTa2326iSk8NUwMlNkMkzadtfm/RuBWYw0R0IZahrATfcUnn+NA6kWcG
Qbc1puXHypdvuMUqCJHhxD3BsYsQla/3vEws1z6uth9JRtfc5IQT06tYmXMu
Wcyw5eEpWVJYlue5VpZuLcBoO5up/FZNbuFxMhCex8X7frrXuilImSVAs75u
bB8WdZT17aAlJgc6YH2uDV7qtMhIpeZKtCeM3Wb1CgXMiRcuWSSOfdDQP7eV
kyaTOPrLq/gKvi/Ft8gisn/OYpSQrsf/C+DGJnBQrfF7GFRusla4rXs2Lajs
3v6oVQlKsPkF3oacZqEclJ7XDz0VQbybXGuYWAfvFodYE4E6wDJEQowbj7Co
wEL98oEMNm8P7ReM4ieoe5Ad/0wxbVjIK8mz9zYCM+7Ovy1ogPU2RB0fHjIx
mBZu5sJu5znAZVS6lUlLjE8b9ajZ8vR7tiGU6CQAVpMJAOU8JlnoMfR9wOx3
4mzPZ6S+uON83G/TDMETUE0xQeBQ8/vwkW7wpz3gv4HVDyAstKtuZtEuTcVy
BmKMvUaR/4nfJDvcoOAJ9LOo5gal54+jBddWMD7CmCqb1aE/ZRkMkrn9LZfm
oEmfoM82TcrxUql5iLD0H5SUeSDTszqyM3vHJjfjwfFpb0h2AzCeY2U6Ersn
8Uzd+/BGw51EqAW6s07H2MDkshdleX9uStQeTRm+gQnyqTQyhC6ChwYTh8o8
Co1o65uvs0Ehx0uuEEISkvBXPGBR9QRhKt3d+MipmyFnGvmqNJZy8ihHPh6z
L38X9Rb4ZrqwMjZhSw8ALQPbo0Vcvk0KIWVQkn9Jt25OfrKxwiyTHcz56yiz
yECD1HDnMtd0aQSoYKpQmGVk8zssbLi9K400vE+p/1Wty675eCs7BTSEdB5S
RZmDPJUSx5RbrYlT0K9bO0QtcDE8V7ZhFLfUcM1pHTDx8rSIzHVqF4l50tn7
HW4tHAW9pgmx0q85DxBM5qwaWToLsx7A836mRZ79h1SiQugBkjLiqJ1s7vVc
UhMr3f6jA6KbKZvdf+hRUaM40pqXoc4GuIx7BjZi7sul1kFJeuKyZ4ybAJ8S
n/j8iKQf803Xh1Vi1wiSJF2FdXIgmwEl1tmlIsVCtdLWRt6SVEoLR8aSWfXk
UvmMX7gSDd9ONNcMohp66wKHWNYim2i+nQxGtWXDtlROcXlliIahc2dX35JS
3TYDzF6zck9UJwkD73jjFeGV6rbM9JNt8ZMQaHRd4O4IyxYctGvQeds37ygU
Lsu6iefGneI0C+J59mu2f2xQqDIgvVjahMrmN6Xe6TTxw4ckzE7iw8mUsHBy
A0jnkOUPk1HlQLsYFYzRyQSKzCTGn/MTHr9bL3h9agnSkVZtCdmzIEBOE6BB
Zs0X+iTFAez8jVkx2ONC6TwK14Dq4GDy7aesAVRlxRWa4XGNPpkINtT00wKf
em/wX8nXBV0gI3WYFVgw9j30zs/5k9C5QARufnTrOfOD+NUlKTA5q+T2y7ZT
vr+3LOzXep7WNtn1nvf2BXtS/2sdZUucqrFbb/0NVWaA19M06Ia0QnaBEK70
VnVJW7+u8+aZ+0MosIxSvGHw3s7jUbNovMAO3czkPQb86BBviMnQIV4/ftkl
YFcpM4FP9GuuPjRjFOdPx1cYh+RzouczcK6ndl9BURHgaEm40sKoiz4iuQXO
X7WURduUjNkaWfIWKT6KVps6lEZQs6ASpD+RmRttbdk+d0N6uCNQ1uZrvbbP
33/UGfkfDyoZ1uHbT0sFXO508vqTUatsc4aAQGSznzm6zdAKrHXAGdAkIhMA
wfAUIOzx2XBXTpPbHCDaVnd7V0ZVQ8MNKcm20MFv2aPuaH4d6RCy17+XAReF
9KLvy1eRdXJDTw8BWwkySRXW6zxEB01z6QuuRo4Tr3vLW4vnIqKgGB1aaKW/
v+5pnkJKq6FcDCziWXzX9o3S1EKPl8o86P3aKOxJbYUBcfSFcJua8NOGOvlR
OmePm1d2OrA+Av4DbibdDQ2h73oMSxjYWga1g7AaG8wJ+FNKPVD3MjK89exg
ukvO38TWmSo+6W8JmPal+cbbvI0yK5drRvjawgIEoKR/6RAKkGB8ORtXTuhT
BDhh9pSEoFlfIVE6sWd0dVFlK8vME84xIkGIJ+cufg3dUXgPJuQ3A2NIo9QV
w51NvslY4gglYEGku0cRQyQx28laAC8O6lVJTHb0dTPgnoGS9ySiKv0npXgY
DwSRxNnA5ZYsnpFnYVQ3b44pQbkWSx6ALP/GircXmH+NJzJWhbOLAWf2HmA5
1j2cvQviyzWTdpUJCnaUBDC5ppWwu564e6yU2xeVNpFZoKswAwQY/oCF2TNv
UgIj6V7gMgqUfbWb6Z+51xVmwUj8cJmO0Juv3F/RizTqqPhxDdPuS/8HE5vR
5NLCmORJ5+bGlXv6aivAUmtNcuy7nD/nQ8NYnQBEqql0GipdhA1BsmEE1tFn
Phi2PN/xlZtJtlWnXoPuMZUZO4S2O7X5yKsmXJOckoqx9VGSbh8EOX1Jsj9E
y1DMMoOEsSMt21d/gh3jCyxoKEnZ1VejKtYv34ja6Q9JhmM02R/G3M4pGUau
Iwuzcs1h2ljS7IFPxTut66KCEXSj/on8vtgx8+B7lq/skAV2WJgzPiIf9B31
K8m1bbn7ORv6KVIfBlbcXhENdaiT7bYykHe5wFtNHhEYyNF3SYGThiR8QVU6
TE8H+9gZdsViA/gla3yq4hctH5oSCgdCQZ/1UX21GEsxuT26LIKCL7aKMKw1
7j9vXSNCeoK65AHP1PtKE1EZgLyz3l5N9dC+KJ4gPqQQjiq/m9XO0hnz6Y1k
gFdtvMCKqMT60B1DlT9fRRa3POgVEf2DhiBG9allnGOdtZh/SbremKA8B3UH
Xk3nr+w73WKI3kXxYgNkCfHXvdvd32dIRi0dSfQqtvx66fcyBU++kH+nM5zD
1SPDIFMmR12P4+OZ16M/OGU9ceqDZnarby7L6b4jKdB8F4x3zc8Wfb25n1HM
IqGq2i3GhglcfELpKqrvyL6WCWdppkVs6lN+gtUKtSIaKZA/y8Ih+1stPLJJ
pl4JFIdPJ3P1P0hTWLq9F6ir33Qy4ZhCAy7BQ2XqFcQOKb3SxuDfseNxneFa
qZBl4lHDQ4m5HMRH/rLZVRy3Wvp5m9wStYcofkbxNu2jQXjNq8r01f9shReN
7hh311Mg65Lw+YsmX6FoFMB2uxUge3bDWCbAMHw6EPtkmmbC5rk5w2wwmnoD
LrUDGF91bIBdoo3L6TGeHYkN4VsTOjS/iQr29I1V0aJCnNmnDuFT7iTYjko/
AHtAer+OwgmLhOCtWlj3V0wuMG7TX4OSkwtlI5/G7+cPfGXz1HTuZyfgoaNB
zXSn0QmSjfRLJpvgCoztn6RqXgotMpWe50G7fVD17TCfQyQ4uGjMqqe/qSzw
jm8AmgnTWbQIW2updN6Y4rvRs/iGy+WsDoddRESgnFB0u72gsifqWoCONKCe
yqvXk7o4nbA8Vlup10tuneqitOgI6Khl9qBNhcMUpkZVgrFqVdwZOczTm27l
OGgJ5pNTi4hG1oPH/FH75nozhmCKr26GZ445HMkdB7PZz7Mwdu86MH6jYvUO
dWY341q7eWRDAv2JuecTDYVYIHb08aA+SbtXgBdRe80gnYUFwfHhV4QAgkzl
o4HsQhdBM1C16FW47Js49s0dVz1iJRqYiUVgviIRrJFhsN0HCXq4bPyQNCCG
8v67IqgMm6cty3gDxjBBhACGVBX1sn4EeuAalnB2Xtru5/tNfwaaVsLcv0mf
E7oHWIz7AbWbnpZpxHJARbFIaSQl8qBPex16S+qgWVFXmPdbp2mshDlirJ9j
yENGkkkHqO09eYwfepWxXCSSu7PkTIdbFiKwCjz6rEIzg1bacTgH7yc6AswS
dICd8IX/ug3+v0ziCwn0kf4j/Kt/NghXQf+Q0BwupPy5r7lW2MOqEoas0TB+
jWSMwu1m09L27f9bjstDCiM0Lr+f4d9TFZ+gpKI/MnDJtdbhvx2mGhdY/QT6
Tjhv9BuklIm+FBeXHutvt/9y6lpQsRdXTdCkjSgaR5nXXSrz/l1Hb6MHrz4k
DPT1PHPLGWrN35gEc7wuDAjzyd9obbH7biS0oczLrnya8imnIP21Kggo1OY7
k2SyGIRQdY1U09N9TLKjw4MT1gc4s7BafMZZFljnv7gLN9and/LKmT96rVix
cAtlRrDAq4bxqRA7My6GC8mcpbyoQwaIgb/v1ZeXSuTfptdvqE/a4ZqgAd6y
W93yumJ0VFtGANayHFpX7ftwQRsmm2ih+7I03ZoyFYXJA/IVrQnX/9JxnnXO
817BbbdS1jEwXGe/7KNneyLR11XNQ8V5A+Yrh/sCxGfnBZRLRwYVdHDdERyM
ylFjIRjcRZDro1Agi+VyS0zzeGGHXhVXvbeKDatPYuV+O8LghoeJYL0BOQlu
yHh1FiGxTM9yDtXmavhXqqsIpB3IQrgRH8D+LK43ksmKXEzJNse7uVLnX9zl
z2UAFqi17j9L202H/QhZFitNK8YjOQwFRqVZQSlmD1vUiK3g0SIdxs5zrKtU
K+Egp0TF6lJ4dxjZZo68wpFIA4FZ9YH4Kk/eR4+LGLPHZHwKz8UraJH6W3lh
o+huURN+8N2ekLnqOhp54W2a71EDE5nXaaFh0sWihbHW0gEWty8/3jUgWl12
RZmQPkegdX1aYPy0CrpevBnZJHPYOZvxESUwnBKAsq10M4hVciJDiOzTfkX5
gr5NpyGIZBuu8cKSoSw679g2D8XlTh1E2BXiholjyvBtyorUQywBQBcSEUe+
dRAD1ie1smYT+d2vbHMbAkrysMNCedsZKLz6DQIXz11WLASedADP6TRfMjHB
dupOf4G1g21t0+OtGkKfWZYwbUttzWw0kO5Yu7622exPRVj2A88oaxXqIAc5
uiFfL8VrnNsB0B26MQZM1SOu3KSLhH042mGt9FFab1K5LKJOcgS+b7RAKpYH
2S36kE8Ie9lKbuTV/jPlaQJOY+qP/BreYiv4q1cJszv+V64Dhmn/Uw+se6lq
xKGbTkqZD/NGl3H5b1c+L7QF0eKXfwp2/CF69+faNN4+vWKXaSQWPijQ1875
WExVYmERPXAQB1OH61iCZgtBqU+QR6WOnYLbMgiYWTr2OW6hOjGg7P6Wp4nW
Z2UK/idfma8iTD2klWWATVjlvzs5GGtkvvPRgDUa6Xawtaf2HRfl+qmCau5O
WLFKlR2YIIXYK0ObziHuY89SR7zGLiB2tsky75k/jWj7epvAW3clXbGI7S15
PfB+GqQ5tM+V6cx+NCNfgP5UxfOf/D2KqKZfhrYnajUgrvPZ0jqNwYjmFLQO
yYG749F3cYCuagoDRp/oE9xMNcuX0g3osPDxu6cjHJQovk6bo7XjDJIUohVb
Ao+GuUMR2FrONeJqNkwiSiaatwAPzrxP1n13EK7Y1mk6ZwfDcy103U8k0IPe
UZ2dPKOS0wPvjvwGvT2aopJsRh7ps/86TxY+dj+p1NM1rRJqKntqIsiK3cJy
7nTFFOpeSVF8hUQeGALtsZzs157YBvDXZsctMStwhV8rMDwjPfWDbtID2MR5
kC4lgjBbOVFf0WAiXzQEsOE9U5hEs6IfxxybF1u4y8plNunM+vb4iAwd2z7s
8hzp9FTyjNiad/qCXCSTH7LOeaT4agX4f3q3VsXe+mG+CmnsIkTYUi7H6ryM
vmTJxHLSYPlNZn/7M06sLxcAkgqexTBtT/KrkZ178VelMZ9x7KEKw3yQp9So
UMiozQyYa+bY+MFQ0YAhO02wTSfqcMXMhKvtBSh9GoeLF3MMBal0OpW2TRa9
Qp99463Fwutx6rxGVtQACpa8CNZecSkI2nN0wR1nxXuXD9oxK2eH/K4bUFWd
9NVVsLdx0xZLl5X/WgJOfvQWJRjDAOwNsr3hyfITFZxtRowEQ9kMsN4wRn9O
LHZERarZpQBGfmLll1anm7BjxJBcfUF2jqfG2glpqCZdxzUtB+RDB0rup5Eu
4j3lzvwb86JDFjLW8QL/slsFTo2ud2iqmDSN0D5YDgZS2LV1F5gTlmxGTZow
7qPy1uh6DjqTPKidl92uvkmr49zHhuGYY5ygF+fKS+Z3HnG0xuhLsD3d9e/1
mYwyQL7Vx7I28F6+73QX1UKP6m3wX9ZtY6zXtZczIZcTB+N0ZK442Xma0BYG
yK05ugpNco8biEXlwx1DCNc31wHbXd3mqpkDhgDxv9LGxYakNJVHeTlt4KO6
O+gLSYM0t0JKC/KZGiiVsSmUMIiOBP7Wg6xmSS8Yn3HYXnS12phT8HrScuwQ
e8fAqadJQoJ7wc1WD7coYcQOmgFxvYNQnGgInYyRTDFIJlYsR8q5nm7ieFHs
h8DT/eCMRWSP1DoIxj4EgnWUVUI1qtf6kQQfTmkx4V3rjJmwEL/Z63WMn6s+
/waPr8dvZtt8mMBzwlN+TmYKadRlmqX9cO84Bm1UO2FPzxi+SzW7HmJZBVe+
XH8cf7vmVBjPjMVyDOfeO632HwgKMk6nWAQTLSvl/e1Sxa5PeNFFS/X2snGP
oODBelH81+LHcwKs/p62BpgdVcJ5llv4YTEN5lrxDdyJRsgORXEFjJh55Ghn
Y0zLkkEayYBe20lijbfaJ8Oo5vwFZ1by76N4cPiG0X2cC5H2MD9Trl5842SS
7O0ghSgc1qeCkxeLF0Da2FIgDTyw0S6Uf5mm4s+nZ53cZux5RbTXvCXJlM9b
zeU9kowlixxCKqnRscxLIq2tPCPdiqJHJKA2/TrATmXoWZZZCQCwve9VVS23
icqtu/dYT3gmaQXvj9YY8SeZqVN7UFiozMYQ6TAAUMIf5gHy9ZFa5pNFaNbd
MnqvAxyx3BHqTODWMmMB7t1v+NmUY2QwUlCGJZcN3nTlYJQw4vXr/xioVpkT
4K+7JLW6xuLYUNFRScJKDO9LWh4RDUS1nUhMjACLn7KbUxZtc6CSjywFrD3v
5lgDV5IfEzxM9/kY5N4120aYzhY94f+X0+cYGvI8NZ8bIgGnui1jf9FpW3LI
CxRQdDP5rW9A54CvPgE+g1m7d568AmDEoWAql0VuVJJEjDBGux0R9CILxaPW
8wjLW3oPpSk+2EngB21bMBpjkjKGUyo8rQ4V84hAi0e51kujLieAGROSQQsN
hhbPkCJEpj/kBqKgwpAeGQrmwoJeZ6z9dxq3DayDFDoSfsCZe3SOiqdCcoji
HnYgKGUz+ozfvSOE6l6Y3o2k8bf/BoTzny7ghAlzqVzmz5gqzwOoWZw/bCrf
H/oEVLDWRy7wbinbJW1xWcqAPrOELD8h2d3VP2gS8Qr65fNMEyywHGs7oMfq
b5Te9yQIPrPT2i9YQDQ24h3qEpZ7qiuznhVXeW23lYmD2KcNOMMczWmm8uVQ
PZ7c9WRK9tqFMyZ2/jYw2eDU+Y1GhAgXeg25F4EhebRaUU7Ff0pO2vBRl2t4
c4laEC7JSQzaFLVQbmDWr8K7yJPsWyA8M5rQfiz6SZWVEpkRPMVtALeBWSDu
LCpYzfHxl8ffpnc2/Mtv0bHHNQ8oVdZe3aU1bMjDmkze/ycyJBUzgF2h5r1a
JITQwAwb1NrGws3BrawvmuR7hqvvNXC+/dyJGI9/OFTztYzkZYOTczowK0BO
5cQzuPNMkjsI45/DcfJM1hG6/xTSqmrUYNK06pGxk7+idRtsExKW7M62FXs2
G6xPwvu0mgd72acwYYHIE5P5yYsbumeuTJmF/rYn5D9rBpKwf1aur+NERMtm
wSYbtvKYH+0T8CqmfDQ/jYx73v00ZK/cmoG5rUaqcltnaTze5C8oZ8PoVhiq
eVWCl9kyuQXTLuUOaIgOtT/Sx0SZhf67YlgFTda74rGK/xpyrR4A3eg818Cg
r5UhdPRUB/YH1O5Bu7MaUpu1ncT37nm3pclggFWHTvE62c8XzzJAOQjSKzXl
jNhsh1Oq5cxHylI6rcD9qFoyHOftiGoOgFq5CSkTzXJroXcxh7i+0rRQfiot
4mVu6YTzJqIv6NPaZD6JWjn9W1M1Bza+gDe/BRdQsnhSsKF4lzTCKgmYA0Pj
mzgHNZ1WoySyQ8KXTuQ4d52fINiYUj5udxK3BS+VBl02DPtB1oro8wNZLO8i
e1s+gfRB4K5M7viwZoNEG0RBeEKVuf3eF8DhVZ97MkzBH7Ig9wt5/P6+6+64
dCTy3Lo8tP2iAW4RXKZgo6ocK/PauVtiiFcAj1Mp9SMRydUsZ9sVqHt5RwTE
qUJp46WIx0MIrRhW/pFUNe7R3BpaqC94XxTfQ75YCKEE0y+othuPwJOZYbFH
Kau0JaiePpeA3lzmuQHvqIW1ia1MTMl37hV2+WbSKZFTtCYbf7+9wO7TomjA
iYOfpekIg4m6lN3L8Xp14P+h6GD6dirDRCNZppYy311Ah2in68MKFZZWVyr5
/Qko8IyFdusFyNJS5ksfcrJrNSF84VC92s2mdjR5cZx+Z1o7EGigen2blMzk
tsbkZbP+B7NyMtLkdNxQtd3lD43ZCte0/xPCkLw+fc3LPi0/kiIklrXkApLM
NxvvBE+Q08ew4A6wnimp+PZ8ncPjDF2DxBI8PjglsfDvg3dzasHOlHOXF0Pl
vKQi8Rk618sxscMHumJWFlWoVfR0LMn+gCackc584p72jsTx5Kbq+GwJ+W/V
fi+uPkz/7skP40G3aP0mimJUZcN7zSG7xRQDlXAp/NlwCjyMjut8o89CaC4u
sS85zv3Wt3E3IchgiENk5PGCVIYXI7vmPvXD0lihyd5JNdrQHYUzWlwC424k
sIe6Esy5W3+Reqwo6EnuGWopMJWBm7pyUItiESUMWenViHlRaYzEL6NFaBuH
RAkKjtc/oM4RBMlmnLgRRzlkXmx8Wdes9KAdcTEmiMiLID2C8d0p7WnE6M0m
QEhZuXofnWcMYxKYln8AVeL8UoKXhFuujkwmLUL4YQjHNj2qZXT7Gbe/iloh
wSTSOO1GTuI4JUzGmBYLJSr4aQ7hbA88KV8+zYQb0MPvf81fQM3uH3dSE4cL
EvtjDIGL1q4/Ef5+u3GEb8NM6ihQkOXSlljgOvzFx+ZdOlA9KxxUAwlBXG+J
eNz9ctJ3VUJGhbC5VF6sCNN0Zek+klmh72cCtzaYh1fIXuN2c6ob3Y5LsK6m
t7dcBNgG2N7rdQoKXgLAYG1Simt7yzWYzXMLBVFyvfq/o82f/N77V2QLwcD4
auJCXF1ZRW1DS2EPIvsh0KT4k2o0nytj/w36VKU0rAqpQCNryxrKHCT0ZL2L
WNpL2SKWgP5dF0hEovtM33bw7yZtNcgob8JnL4j3KSPOztjABMt4m6NuI4Fn
NkFWQpRaT/OQ2cgQKzH2cGxujIrIqLtnx3Rdm1FGMp6KPOOCUDasN+nAONyr
EMEXxEAo1YQBJjNMrFk49iMjsXBl86p9CYyrRoTxfIm7I5PoqLOtKOQGVIPF
QbtUZAueUuXBiLLVHK7sjTjB+DE0jJpniMy9ikpkiXTS/FHQMzdV3FOoyHHC
yzFmiZcm/mTMv87rFDbHC02GmUd8iYvfdsggQxj5zCJH88TmjTPth7yYYPc6
5/SUmKHfiuUpoDlIEWiQ/IWhhweHZyYO9yzq9nP6UwQbFHxm0KXWuVQv9guK
MEPAAtaHwU4RcgCk3Yz1a+M+fM6226K4jLJYMLjbq17B5OSuMTWYZTsP9eQH
cJdKMHkyuaKhu4UGU6gh1ZFo1RHw44TaL5JNJ2gMQm4g46BIn8Nxb8YN0dZj
3suVhyS3r0DKQkTy2Xs+iozidpkdydgvGGoPpPKWHAqiusEsOpNhKR1cPhEr
PUrm/zcQgywoaejw/bIOCBQiRHIwkJO42zfFbszhUPTUVRN3UyWPzQmG8gDp
v+xvjGxWRHtOwpZyjsmmDGGS6A6FMhmaFDPZDeKmC8dfrOEgzTc9rdJGFLTJ
2OGqjyTqZfMPGqZBu4/HIb1yvYmxEZXLwVa6fpEK0fbYDX38m4JXDPVSl8gH
KhtP4iuP8g2IVhyp1aKZvpPCB2LQ6UDmiJHdjojZSGzrMdmgiFNNTvTVJ/W/
TpWAgv69rnovYhRN5X6PBgRdGrhegCxegSm0O5xCVpTSJBj+zDPyA8hZ73Wq
OdrgqReAGgW3bU7cjCcvJy+7ifZEOnOK3iMSgMYRljq+hUMIm+tCwaDs6ick
83wUnJnBD9WFQvBYws82AKR81OYAVXFb/arj1+BlDYKu9S2klFcrVSuuhVV7
tDYmLqUbnzAFSMUb7l4qsdZA8VVAmi/xMe4p4HeVlOhgdbXYRp5covhzoyxl
CfhHlF1Nz5va5it/0r/OhsyAJxFlnvCn67hwwbgbRHcq/b7xynxQ6/Kp4U4L
gNmlgaCMHSZ8VCgDlKWniIAQSmqc94wi4AO3eFMNJVsXvRxkNkBxquBw5Q+8
ujj53SsNl6jQu2OSx/I3qZwOETHknPQYRDZSUslDsSMQQ46A4P07MBKENqnq
SL9gbpoXGPhQsMtOahxrJGf6ZierQi01xYRcIOAUV++90PynU3I+alf4oXua
Jp4L9rm/pYkhxp7BWiAmZhlpOyQtv1ThC6POM7wdtrMJDY5cDW6YAo2ht5DM
1h6IaSGyGj5d0exGAHw6TVKqFVDQ9Q8qALC6OfwD8svd2aq4cm0rNah2Ef+r
iXVJAPRVZTj1d6GR+CV/jP1jwC2hJq85Qt5bhUEVYTHOAd8xHjR6IqgY0jsB
8y/T16xMTPzDLY2ljL2DnSyD2jD9pOZbyuUYGenSTMXAB1ldiRyhYScgE7dU
lNu6ljeR9Rg/gp5nlRYlg/yKZcg9yd5I//T8UQ2zKoVljivEl9S4aKmT1S4u
4jANDajUjoIciIJdn7mo/VKAv6y0/xdNWN4LZurRzVMOPAfx6DGTZNp6tql5
XG4waMMuTsxkGMfJuOSbMYMwb/2KMJnCKB+ol0xVQ9tWd/WyYR9oEIDUsgp5
p+OhWQy38Jj8witK//I7kGnKaPeQ/xMZsVdkhAfnytjm9c0w4b+DF/harv3D
DILei8GS0jx5LJL+06fcLjU0MSMNSMOSBb7TJwhMTsbY7hCX0vPZBFp0ekZA
2eCaeVqNgDHbcdp26VQe6Baqmz2U44FYUNitjk6a1X7jA0MVlNVRJ8+op0gh
2bF8wiRsBMoXG00XdRy5vkrcADSJzCw8cG7QGg75ArYEDxkmVoY33m0g3lSk
CGrVvsunxFlGtA6p1OGOHLfMTilDQOnTaynd90D7FxHMIBSTzeDKcLHY1uUy
PX26Sxd258ynALHelHS/BjE758ddILFL07b+2UVwfav6REpOGkE/8We6H4vD
zGModpG0qKb0MpPWhMyCjjWtciMgtG6HPawq8adUSQFvg4jJbNT7zkPN7R/v
J8BSNv9EE642FtsPvfvTnRdEJ0w2JdbkwBZHqFs5x2hwn/bxj70jH3USBo2l
12B52/e5QLGHbeD0HEQr+hRx/KH3Cf6tiAcCyVxuGhLcL9Cd45/DsbRoVt89
jttTbRLh/hcqDJk/m9pMjQcEvh+piqC1L8qwsHhfOTgHUsodhgfahkfPBL1G
GZb4RdWlYsNwHzMDhjnVsW43vEAHRXjqfo4cTLQgkzRzuMMnA1cwDSN1ukV6
qOLksqaRHKvqQOgx0SznvjJSiqMHF0wEQI1LJqVHzthe+JX4CHhoxQDWA0zV
AtU7a93mEhOaIBl4OJQv3efQj6YAKcIp9wv99W1whkfm4UmakpxjBR0rWudS
6Gp52gMBNUjKSL1KYC3AZh0bqJqTtZ+AzPRX4Olkr6qZ9qBglHBAX6lTFvpO
8r8SUT9K37mXcQZEamWL9l/x3euxUMrLZakdnzjluAMFs8cwKCgVgjOckkgN
DL+Wfqoo/BTaDaJZFXEgN+D4PZNwVQJ1/p3hkxh2GvgT86UyweAftiJnrX8K
5TL5Y835gjK9uLBYTlhjZcJJr8kBjohRuEXHPxg6AtPNazlRWI7gNSXb+qro
/GLcCzA+TzIKgVf+UGfSyiSxQE93I96DsqtSJrZwPE25AcCsP48QJ3Gdv4C7
4s5Ep2+jt+B4kz2NotTCGF0kMM+moRVvgopMB/qqn7ZW79b+dZIYoebRORrR
YlA+iltqxmgT8eUK23oRRXMz4bQJqJkvR+552MoldTqKxaB0zFa2P8Zn5+hq
hC3OeGnrwSTmhnZLUbs8j529BAm99V6KSavEvXFkh21aXXw1WYjv1U/TIgIc
867l9OqoJe3CWZZxD03ZBusumtKcnv/Yr+gP+O/AW4Wz7kZjrqgPJ/GwkmBy
NCo+1gBSGb5WeCZKAM8mBHQ2ufOH0oCGKM38QWmqC7BohHDUSVJZRV+VqgGN
JM4FUIOLWEFRV8Q9F0RCTwdfCN1lTHXfAwEtcNuL9XJ5ab9dvIyln50sUCea
RPo7GiYkBdP9fIb5Vcjvyn2Ua0RZAfPSpSIMJD4nIsRALhBxiGkk69cn5be3
/P/+FdiOzQUwk1kd7aIeWXFG/MD/DX4SJ/KlF7jAzakAkoctw0Tbx5LeIEkw
58q/Tf79khSJS+IILdLBDcjjcHoYzWWCT6rZXdX77hceFl3UUiFuIKSf0QYj
WP4rpaVph0mmv5QXpofdNBRSLiXpc32RXzFS6cikmjjlx/R98H4QOW6o1taQ
NME+GdECdAVR12THmMjCZj6FqsjQeQ3WIy5AyGAyF7w+DjvpeN5LQVvG8Pqh
nU/3OaQfVyUe8ov88tfvq0nSaE+vjXo4Y8fn5rRixE/jK+HjYYeW9hhcCfKR
nBBtgvQwbGPQ+GUh+PvNSZ0rf/gpVNRKqfzXXmBKj637ifNbOvl45oQQNMHX
3rhvBBUE1ky5cAWBDnwuUPVrBHfLXJaJ/FEQSzDHSpgqJwB2z2dBgA6kP59D
WOvZJdIfrhWjBDGCliBgZaD5o10xGRZ3MdKEmGwPpcg/RMAVCb612ndZCg8J
6ZZ2tgLNst/cd3LAXHvQjmAuP1F3T2r2f8Ci9Lu7m+fDx68WFHJxroemUCqI
GDRwFZrMUXgh4tSYPVyEh7AdVQbYsj4ilzJ2BKNdBQH7xFxPonV/IFxUAHjh
YvdZxqPmIqFRwblRVUBKTaJX3yOLDZ8umb/vbvCj+WGl9xo3o0bRx+rIT9s+
MW9wcL6PtWVH0Yg9KQgd5Wx+dcHbLWlTHP7deByWRf0bVJmvT3iDDvMgWpFK
E6ySVAKghqNgedZSvyFCDU1H56rksYXfxXKDKDvKX0zciZpH+7wEIPfhWQhi
tDZZ23QvuDnuEzIyskdmUwQPv2LKDA6lxAksoctcNDCdlOZ7+mpzzD2gQjaG
jJU4tDJyWZWlLBl9XRnG/SekwB9/6dgqtb9bYo3QruHhDg2p9TxW/abu+e3J
/g+lDjSB0XCKBzyi3NyK8nfY10Ae4g7nWxyy9tQ5GB0s6yPtUnFnLI+e/XFX
5QecqOxv8UKpLnCVB0qRILu18AekZvyQIFDeLfVuhnxXvnsIHTCFuwrAvayK
YBwd9pwchSQJYB4wkjHNpU1MWPIPmQzoYrFHLO5DXG2zX7qWi4rZ5fNB26Y0
rmT4UyH85EkzebbT+NUsErCN5nUy8Bqniy+uYudtIqOEcqCVwFNEE3WtUchj
4oZxMbkaDyl2qw9jqzqiCcHPFd2NehK2F5tUq6JDDOHi4HyhYmoUSgd0EpWd
mqhXJT4TfgFbAD28fmrAFRBcWtX6MnaR6BfaIoAR2CL7qegTYDN3rFwFfG7K
c6AxPXjVP8IXMLtj8zsWVtU3dOcC2zQAurRpakxNXDk5+PIhMEQw2fXH6QZ1
/Pu2jUz5CDsqgSdYllyU5nxgTcJajSFG30DD97QiUiNS33yMmEvpQ56BO9Sh
Rbw8tLyxSqRWqHQq//HkCq63G9vzAkS7v9hdb5/YHgLXchJP978vnzJXzJ74
jn61GN5UPS8Z2ygTf4IY7lV6CzmDDGU5ZCwXGWsckuQ/yk2GyE0DoMstqz1Z
cyuHfPIJNIK5OoUmu1U6YfzTAkZcvWWmxH33bEWhNaNrr1P5M6E9z7zjGRIJ
smv1mT0msSLDNxu1dif92Wnb0NOJOAQR08KFO10XHWWT1d3O4khBCHmC890O
HGulXr6X9kzPWHYYfdCHdykZw6J9u8Pi/C/Ij1KrYJYy3oYDreDnqvx22nEg
k/NXoXMtgLs+G4/kCxRBzmwLIdl+mqrtOVK92LLj2/HpgdBHpB9F+a/+foQO
hVxf4rxhhOo8o3imLdnatc9qqq4OzXAbzj97iVLfluc64z/oCNrhT5L5EQDR
sB95Avg6QN6QC4ByKv+ufaJiiwYAmBEAF3n7iGZYtaBxOEUkTOwsUIix4xGy
V6w6ecHmJWqjpajLeNqNMVvsda5xST5MA8ifUk64UMWTww37driI1gf/1mA+
2DxXBIzT+mXpbauFQndv6UqglI1pm9JaqaW0yDt7DiiZr5jo2Bk+5nh2iOsA
dwRK9WEIgWx8hWMrY6ZaHAtycsDhHQz1ghKlS8kLf3+Uij5pb3sUK1toag3C
oIdIABazj9gfIjN62a150TUYS7Ss6zN/nTZe+/ClqPzR3ogM3eB10W9WwUdL
WJimAQaFf1KC/4JxeLegYpenlKtbdQVWfGw+x4YcCDvhFLSW7Le9XYMnh+RN
C1ERlvx4eJkx4Vq7JQu0UflKNPFgmf159MZ8KFuHFF2lAb/NKRDXYrDZv4Zc
PbwwJygcFncyohtl+RJUejbcbjcopj0np92VfDD6HAgaQZl85ZHYyPw4tNtA
0ffsfBpRiQYoePtXYN0yXvoM8rmUmmBegtCXtf3aWMUHj9XKhkLDBEz0w1Pl
6UGBXj3W51goN+h8skZiOua363iGz8eExTuHwo7Kv1f7C+aiAYSFC7y3mkJy
Ev/hborNbQJBfwyYdXZjgZs76od+E9+KsURaLvVlQLIMuCaXGALJUm9vRynJ
sY3m/QzPhQ9tdHkCk1UXFZC0b0oyyqyVCPLVw/RCINO0j4QQe4FR/DPCmSmc
BEp/ESItieOZZpcK8XR2HS7HqgY0Y6/WiTpcQkeSfROCpUrQzT7Yu/VYU8BI
NX5RAcoaBstbYzBV2AeM8DA1SAzBD3J3mU16njZa0huIZRYbHvDsJIKuYWCg
+7M0pJwr63GrQx09EJHqTiNZAc+0bHhtGX9GP6ViQZwnKbk6g6D1PDEK2Lwi
2vjdFcdsyn+37TwLSXFQZJBKxucXEbgVhrzE7UqU39QYJm1OC7Pz9mOLQM6l
4C/f/duIVjY+vXhyeabBUfSmI6JOxUfkSQKBx8YjvlST0XVqGFHPGpJHowFH
kIEcMLvmAGLOWQrp1yMZr6sqs0Q21bPdN+kCQhm8UBJqOLFF7RWc9xbQw3Hs
q8e+kgyWvq6j76//Hx6b3C9Gz4EkptakVUunk6pLatLM2QEGewsU2pPWczby
5oPkVDXm9cwNQ+2J3K5anyxTfBQ5TABaMRfYBt1u3rYmDBopxiL9H7C4vOmc
o0afriWWZoyKbTshnFo9q1p5t8plL+ViDWbxbeaZWiUSeP40dPO0L7B57yAb
ffhu2h1CTTDzbNDgJbRo7yw+Lr3ly296k0mwlZNxwGRQgtEnDJIfx8hNZA2b
eJEun0YjrjnqrhIG5775kJ+9h+tqyqD79TJ5c/dOQ8yGEa6bfzZP3XjEK7Cm
gp9Y0ueHrfs9lEZ/frIN4yKvR0cmwvTlEab782tx4DJeL14HG7n25020zbgO
rP5B2BHg8LnSePfJ+EJFXVQ1+aTVuVfxxKvWWiwg/2o0NRLzkSfktmNhDiNA
BNzmrRphA3Z5vvAYrN0OD7EWYcGoXgzVflDhbFvuRh/1++eLfcjDF3aqOfqx
4mytoeAbLZISiVRtZcTOUzDGKAgxVFb2QsxyFUIqfWFMMbJHA2GW+Wmvo3Ow
qFuK+vg2KYugMwaLEwm+dHzHrvLKZjF+aDW9k7nnPIEu39ns6mU/E/lhxj7m
WGH3bXvBm6t2gCeLJbfo2Zth23mK/xuVYvTk4YrJKdQ4FED6wJmFfAi9u8hQ
zCYHNrmtfdQ3Tm+En+I+2F+tDBIExAYRwHy9ZXKKl89Zzjgj3svwAnTdxPHY
wExw0tZHCHlQM7vqTdZ6XDhqOYjywM6TkwoSAI/xU6HhqZhWNdKAIBh+s1xh
WrupVfo7jVY/wptM+UJAnHhMXHKGp6liSkYYbWZr7g7o7L4FD/vt/AwnN8rM
jAn9K9XVkHeoZ0JPi0HrtwQeXPfU6/uzzQqhh/5xY1bhCgVDelKjosKzqRBR
5uTP+IWtJDe1GHXFRCvynaFebYVQVHH9nmXaQuH5lS1Vwoufn/UwhwV0MyqX
6ZeyNIg7qHI+PmpZqumbegUtj1i6lCBLCF7zwkx0k4eOTHBbFtkuF+RX8FqX
WkFnT7Ar0K7nJJ56NJv4FVNDwpcp7u5L+21c2iIu/yyQ1eNS13UUXSCxnNzu
4rcBdw8atCXGsZHBVtkg0E18h+TLcT9kJIwtDcOhkNaqFr/x+bFmpwLLJeMY
jjPCAwkzz/upLG9BR6y53i3yynqV3/KKaOukcETohrVSEjAAy4g5XD7DGbxm
c0H9M7TYKaX4pufcJfGorEAmqgG7Ph3l2Fl0NR473hHoksFIf3JnhQZjndg+
0XtuiHNw1mckmCrECfpmrAdVqfMR5WO3RJFg1Sy9a0KAYJUQi7FP0AaLlQuS
vAkToGUG6lh4Du6YmlAsAWpLEHWJJc6v0XxLYQRKoe6pCTaJK+v6/S3ezgII
KAIjcvnRSWfJLXBDhyWo9cXKVqwkGmAhVXuHTd2SOM4UhqFvBDtWqUCuFU9B
Es8rm5dcnhljmY7cK69RNoZOc/UFvwxw6hXuF2gNRRPfUPDo3PnTQJK5AMpB
jWHbYwUINFz8u8w1Ehv1W5z4UEJF2GTLdpjEGfM8WMZoXev/U5Mp1tQNm3j/
nV9YZZW79HBXG6LDgC2OyRYDSlI05HV9LuaJ1w9SPWHoNRswOL5Wh2xEKxNq
zeU6rbjT+MNNnWs+egBqak5NY7HdouVmi2NcqHqEHo3OtNIxQK/xnM2ibgds
UCndfHV3Zcd+5GqxDQKXU3hB5pi0jTvnxQD71KzMeYzlIlv0NIuSbpKpCJOs
ETF7CX/DgVaccX0UP6Yt4XDhkEzISzYmaAi2cxK6wBc1qVDzQQ4SvhSY+bp0
KxFPhrEqNOYaciZ7/MF+iWYRStwN1BJVlfFyAj3Rv7qBrMNpZou3p23jF0mE
13n/6tsJINvQ5Ppy9zg6SO5Yi7P0eTq0Fp25GJTHgOEatq3HlkXGNWza3/HK
W31lllSied0rLq1/TwxvgzM+iee0F3ILFC117YaXtW93DJoaojfG/Ctn2ZNs
fA/5qQtf0nGuh1QDFJXV8fQnBsMg42EhrlGhBS9e6DA5MiyzsFOaIoO5xjeP
3T5KX49p+/JqcXJB7rwYQZPIZxgNMgJKK/NXNAUb9crw5PH2NZMBXLKygG0Y
7amd4z/OhSPparlI7A/32wtseGjYYrQw3Zvw5ITmTJ7WYkUk83nEoOoCXrn/
iTN47syvGCimK7ihFsLT2yPRo+ROV+eWDOflDM82hVxqTfY1pXOzZl+LLgaM
Kmpsj/ZxWc8IdP2zAJ9MVrGW26SxzJHDmh4o2GJdrHjz+RmHaoR7lHOkOFdw
xlVN/Nn5SHYxMaLhyQltLjSTJ7j+MWYDZ3tKLZ3BfodlYD/MG6ftA6ke6vIP
d82pJbT8i+WndD1LA8Pqu06/bURfcXM+MeOz6PdAf29dcCMoczP0oXebRs2R
4LxgMSkgVDO30x5+Jv4nhBblZY9HFwdqWCTv3NGnXf30VYSwPU9z+nEA9RGx
kTRdbqZ4EnWZwS8C+XtioC7yOyZaMrG7Mp6FcgyWe1XvOhLzz+gmCvYyu3Qm
e1VUxDtptblOLdLyAavuTIEXF9xLmzuhwDuScRkCBw3Z6UVn2UKxky6wo4Zp
RVY6vd8QQQqczseccWZcasNY6wT0Hm8ZjCEk8kdsEv3sOJCPKUWOuXsd9xmU
nQyWV2A99DGQf/yFwVzsCEEEQ5w38uYnnlHriPNZ4E2MykBxvcQbBqZMZEUg
Mpr/ae6oocQ+yzrGq0qfCMxytYiA4IIGbpHF7kZaPJQC+0x219Bg+pAgdLHV
CUnabOYebD4N6nbdoYA5uHlwMvGemVlBynfMNBw3vH+1L8mArsJbvYErF0WZ
1sEAxKk4go5xJF2gIMuFcpq+hS0dunIMyQHG5xMlz10Qd2wLecevxi4vGS6Q
M8WF3w5DSMQ/i8RMovBUQNUEzGzOMHvLAs12mxsILKENAihXtVPv68oB/fkH
4/Hx0DyF8wxHIMhF6sBe609WNxsuZedGd4eRLxCQ2AJwSsBu76CqoqX6tzQH
jwUTRjB4PThZOJtrGWbmTb3J7xW76EmJVn6PaqCHyjcQ0XK4tfyN74Ko0uD9
VQM7OJULCvbzftYezP6O7Q7G0YASD2jzSbk/Dgdoxb6dSBThnNtFOYH7HGCx
VcqQNCZyr26edMemUgPK9VA+RHFu0KKfhHlGwXlxSe/J3PFRxrPNKOU9eN6R
mV+XAYkIQI648wLgl7EVaqanUjcNarRd+ySLiP+eVjpG/kA/NPpUCoCl6DZ6
GUyzSrYaA0ZSX6Jp/qcj/iVMq3h6VdUQglF1+Fi4zAKkGfeC0lPef4/RL7yI
DOhtNtmdfTFoRFUC8Lu7258yWtbvjD8VoBBwg6+RtD5AeASSud7B7dwZOYLk
w6XH0bbC1KA+x3dqupvQBspsOu7lJQ3MUKI9Z8gjvql9lR8+hk1o90QL5I8w
8OggzoZqIP7k5uXnd2eItVGEiJFvbPXbxHaZLn4oQKhYxN0OJMk2d9P9GAWh
y5NLN5hQd6117PgRlVuqLjXmohyXQSf/6aes1CH8Z4bH0gFNSZACR68qQVdY
d9443nL3HXujBQqDCcedhHaP5sXwBxvPUhaPGvj53GEdQ7P7hi0MVo4x5aA3
GqFQXfTafFczcyG1VmzVq+U1wblt7Y8w4JFcK4xx7de4OxJrWlKBN6nUXpbT
CZawh/5egbYVMP7fWkOjZAaTqq3a4swdCw69zRq2hfJaY6PSi5WD8vXrVJhX
yyg0fW38IqmguSJ2dh/pKdClkUesbtzClmDCR2/aELcJom+wzoawCQef7PDo
1ZCv/4Ap8zxdugQfjjh+lUnlJhEduxgRyDsjAXXKlneVFx0TgjPQzlDuEy+x
ojn48Uj+av5019UgVNFM4kfxlbjEbfOB1d7jH6Ab3I7Rc3jBFV8TsUCR/uMQ
pT/I3MLAaP41OmWYRgLu2brG6ZE8itlDaJuQtHEps/KQ2zvbFLUOH+X2bCuv
mOzFEFEIrnVisEeNej+BBXDfpGuLh/C3Ro9BNwJb1Lhoy2fEw2P9w6XUsKeb
HqixYTqpY1KPdyO49yJQGWVgbKPYJKploaFsGSPY5KxFmaF440xbJv0qpxHt
a67t4mrbpMgMbU3/eqK2YVs3wL8e6YQT0Q3EdKkJ7N/WBga5ZC2zgDqUMSnI
Ek3u8+iyS94jQici0aUIJXUqi/sbv1UA4jI6GxeXaFNVYwi3hG3U7uPDD3OQ
vuPH4Ck/OhzURPzrlt+7krkOXhpuHmUYpV4wtX3DqGk8FNxYuhYjg4A5adWB
fi0dq5dv7p0qK6WbYTq9vEFxFXVJn3MV/pRVXFjXjMRLwvWXgbOMXKpRfJmy
QFhYBeuwPxH+lIKXDyelLpgYr0woZH2y/uxaDYsjrT0x/EeeVnGQfyz1FdbZ
lUZycm1UV3PK120BH5V7obxKL4pDKgdNfQ6Mt7bzJck6eL9W453A5nsZrzst
3y0g3SqSsEKcrXWOW2M/+avBtN3ezUJxhcO0aA9w+Ge41w5K1JyQDl8bDFR1
/1p1RFG8sQ90I1poivmPDEbP0K60IDeH19Kv/TMtv+vfqHmT2Z8hO4mVdoJx
jrXhNEA8N1k3qQc0ebOt5kHUWc3O6/hfx6O/YOylTlvmQd8G7ajy19TyoX3j
wledPnOniL9rOThCNRIhQEWhPh5ORJpCM4XL/TAeiDDBMx5388MVZVNk2j2o
0rhHg1xFolk/XpaHaYBnCAtrzyMmKGEz0qJCxJbuIpOWtvyQ3NEOK5FJnHpi
qs3XgXGh49+7nDHrr6e/BYUTVs/4pR/MSqN/w5psgFJVEBQnYSpRiJ9KyJ5J
/xLGrD+wNuMd4jgZJnDZ4hPMkJoLDgttMeANf1UdYGXFrU/tuvWFXj+t9uXC
u8f07rwVAbyn6guJpGZ4VQIToPsJFxU6UxhOrGj7ZXnxbSZPBuFzTinYUq0o
VRzeQmbMmURIYPEYuJguiF+xM9+2UTYszjNAedPUf3h90DuT/BuaGjnbsU7J
JO6rWCGYcvyjVrhCTjKjJABMsk75hSRpJetqpQwIBzpX1rgXY6AdWnOK4ku4
oAy7sUMK1NDFKPM+EzJt+Ryl6NtVJZJ0cwEZqHPdvc0yA9/u6Yr24cETQuV2
u9yW/E58QvGqbYQcAhFcCftSQbAaS9EW+qYB5BIvQYhWsF08L4QdxNlPn5Y9
xrUeTIwBo5ZYc584VFwWq30X7AtTUB2RvXMwhE+KzDBsDHE/gMvaNFpGj2wT
EtlcOfuBc0pYSHF1Nuz9YX0UEqMHC/Pv5nHr1gqI/SNRIdzLtaUhHd7ZX/RZ
iy25z7Zq02KfM8ivzUNvLcIKBcqc8IUpG9zqylrcT/mDJxMklb5OPerDtqLn
VoHzYidF8e/0VaX1JBVi8xTridmb2qdZViPObc3d6Z+qTgBbUwNKdEGYwI7h
UWq6W8Cn+ZEN5RvjtkSdhAIPV0ua34aBB6XkjNGAMaE2D5hLP5O4DWlNg4oY
z6yNNczTV1uDBSRaIejaY97Ggeaqr5yc5i7vGx2XAVIXLgcGTI+ouNXKVUrh
ZAlmQ9t9Y9cKirI9invT5U7bgYnAfAYWPHHV/VevIl1nWj7m9pSbnDD+XKjp
etUs1p+Qk4Q5r/xJJuAry24yPBGJ/+CbjaADNe8TRuc+M7zIlU8RAQdW/qAf
oVqtLUq21kKd4nGneruKCZWhGiVWZk4uE3Nhu1Gc0qfT4yOUiGoLnkLqCqU8
ejSJf4T5k2JNO48mk5p3Y5KNAJgOI5vAJxsGY0Beu70sFQgeFlCsVPtRFnfz
8IulhjAZ/TlHI+WqOVsgE8IGcwFrYJ0xQWFYVidMTFUpZ2ZiHiml5WOrYGR0
bUoPtV/kubwzHEqMCiBJgFyAzQo8ft08IVyN1xtGZlS3sLO/OZHrcPUDdnwL
honj2IBkKJ8dSfAN/dit4WFoYtfvJ0g3ZFvmwt8Tq4pvSpkgU+GK5945ElSO
D7+Hf9ORFo3ka/uxF/LArAR0v8eE2R8L47NUm+BWaWKaR9Vw9VpxMmwUFcVC
C8JDzat9yGzR/zVjU2dhr2OiaP0ZRVABhcPoiMC/BrgPUzMHXpG2auefmlek
k/9fG/5RY7wPts459dwEdomcRD+JWeOTI6lXuozo4w33U7WE4K5ZD2i7U/zT
L5cf/NQZ09dsJrFMW8OQdxpvAXnUkbUJZtHV3XqeDLnYmNFSE5dWA2rnnqne
hxTvdyKe3Zme4+ifNsWyN7LuG0tmXVIG1TbQoMoA01ylHOeBuQm0moQ91LWp
rYNHHTsE5BpQH1apnXSOaKPviqgV3crOt64G4v2IOgjKXimo/aNTJrfua67T
69L/xira8/jW37GqikuJEnXUx+NL5Y96gQnh+QRD00iuj8KMaNwVPVR6beiF
4MP30XTlwFVQZ4W+4VukQKUTSW8fRODhk8wWCymSu2ZXz4Oibjf0Tf2eeyS/
a9sQOcg66bkg66YcRSFoC4w/Ra6Xg4QO8l2r1Cqo6Nnog2NymsKRkhTlh5z8
4pXaA5j7zXQT7Hi2jTbMWcLZPxjgi1Qnliu2tLzn5v1bdyW/MPYPmbFIvhUu
giWaEPwoGokw6LVHBAeJYQAB4sUXeDhXDjVauiPp178bN+ORfWgVBHXhdvvl
cLpfaUZHSMKN6+9WVw2+U9WF4dBUqZCdAlj8Ki4nMxRjlFWqFXT80qwW/kTP
Mnl32boB2gpwtWGwLxyCeI0GHkLNfFKYiCtRMjhzzks5H/Ers2hzocc3Ij4Y
4/niiPArSaHXwxtkh1DMcBexj+uwi92lwQ+WJOaxcntBBP32j3wQ2XpEsDRg
du8O8l7fRBvectojgpupPuk9rL2Xw96PV3KVrJ35enQoF5VVbXoakANb92B9
vlPtyYnrW73/NrEc3Rl2ci384Jk1gyeifyYvlptQGqFKxLP0LlSSSfolbSp/
BeHC9VQgMjmHvPdCByUz25+l7yZlKypNwLUJzAE+wxP6j8clE10M0IZel6jK
eHG1lLBk4/fMXhBZDnV1loEkb4c4c4gGa23Wp6KSUFoGA42sqKdNJGPRaHwf
taxplgEKtu5JUwG3qeM6nuOy8bu3W8RCauLKIpTNrS129YtG0LM9++q1VH12
MrAKtbIUlWdFX7yfi1NL8ydSFp3t23aVKpGtkli5iwbiF8jOgRS0JF+ih10w
MrppiH4+GKVdKd0v/28ooP1ZzM2fJmLi2MxnivEs6IgoAV3cCRCHscaL56Se
SRVmYdvlMUOkadyiEUCqZfMHA7CY4H6coSt6B+Vb/ofPsjFYHbQUXXvtf3Fb
dZyWYLL4jKW8jydDk+W5VnDAlitczTavyEQdckCZeWoxnknun4yBxQkdG3Vb
SJl3PpRLVXEnnqoY3onlTcXn3ERBN/tEdIxonVwWkUruQtE6MEhDDM8u+5m6
TIvkVaLny2abmzPzHZVTziNEnLRRPxzO+PdV+YLuh4PeGE9qwu2FpOcQT6wY
S0rgM5XIhy6lrfED2E2efWEGldNvfqh7ikisdum6F9Wj3wdBPmkyAyMSa3yH
a6WMlYQAQgHlrEuhAHJ+F+ny50xJbdjrDSv+lOECaruQzmw7/zKSUa6DIZwR
+ExAu9Z7EYv51dX07FV1HrcUG0wW2oB0/WPiAzSfcG1gfzDf5s+2T0oOEX+m
uOVxpsAmS2I4KdfZqCBNQtlJwbSwVXSSctzDLdFw/qmbVs+DJcH+0ZEJ+saC
KgQeAK0pWdPA+vUQtZcYKPMTd71dhVkvroL6TEokeCW//4C63GwfXXMahly2
4sKIdG04Sh4vqd5XJLDpR6BgpmTg6WDlxUasD1oVzQE3aQVoM6+67irYcjL0
Wwk/cUPrJ+wbITe/+/iBXIMbJFtGgy60tMgWa4N5tf2ogO4kA+wqdzb4jToR
HGZUfOR9jnTBFBGIRnfiAMgtibnqvMmYmo/LXmdYSG5BKILFYJOJ5ycYwIqu
PHx4tsF39i+BtEog5RcuswVcLSl3pdNM7co4cvC9IvNNskVjxIh1M6lJkwap
d0TlfznI/WEhuE37TPg7+dfycWtyJ52cqvSKsuuJwPwu7OJXHEpmBhtD/WOv
wMe2xarKLlOqa9AIWiy8X0YXDi3zDhG/0uTJt6hqAgTxvClz+vY4wLPwRpcb
Y47dYPA6202i+L/DpfN+FClLvIN4v8VZNitzD9d2NKhFbtxJN1rflOnKOKHc
WvXaVHXC+fTGU3Inui3rE9Z6nnnIxeG6lPBSAKHRvQYAM2aBFfguJFghrW0V
xrOqTW7SQmhVXFak7i4WOiPlWjzWfnm2lwnCKypvwrPTQ5zvcaCDGY4Ng1mq
w5WY2F/inlFgX+SK7BHUVbjjEtxRkZ138NwSrAAP8MkkaEuOqIqEfTizdP2n
a/ZBKaq2QH9yy5kcwuFIf3MzU1guNIZxulT9SxqVZWBOc5omWsPeY75Pc2El
Nr5wXspBWtX8Eju7iU+r7Vksq1GU2NXlTJh0wS8tGC0tag2I/8iOOCBwjHXf
el81ei29+0squJFJiDiqd05UYEVrk5pZjbB4HqKj7ErF/tyFRatlpa9Ac2aN
48E2IGow61DnSVcRy58qKASDdJCpdHMW1KYiByqHKJiP5tUDIV+rvYIcyz2V
g5RJAGF8qq+MhaxiI00VZC7dRNBw05oXVtx3E/Khwji0vKbLQixT+kWMwyw9
OGYKmXv4/GuNgzJAXocShQgd7h4AR1/TbPblccO2Es2Mlqr9nrXx2QbNoawN
VtMFl06R69pH++Nqa3RkAMXlY2cphuKz6Ny7TLKINw9dRPo5sdmaY7ybzsye
uy93U8P1zUZbcgMc3xgN6qp0UVXfYWCOB1SWpMGxbsx3iAosu/AyLdeaHFqw
cO+apiS7e7saYwuRfiTv3PRQ1DTE/qq/ypqkCpAHdavz8RENs3OWwqHJgyBx
2IhMKAnO62kUY0tpwnLOMwoohJm+rFeRnDXozdogNC8uXerjo2wuQtJh3E83
+JnUy0VXAKoKKGAZ670I4eNkloAd1VGsULQjDFMMRAVcumPaesvVMo+f2QSt
78CE+/WiWJiAbPkDllb0IS/k4mXIY8l5ySwYr7JVzhREPzTlgKwIOxDNAwf1
p6SoxQAlAmh44DbVF6gha4t3r6FmIrg8c6eYMND8FTtkvL4mCCk27zGZRmVx
yqO0eIbyh1AZKxqrYefqwqd1hkHWHT9mS/7RoSjlJ46HY5QEJK2ix0aB68fS
vwcur11C6Fe/VZSyDyyklpZDlD5Vq0kzk++5Gc3jMlYbTX8fvWPzw72VaBBi
5l+37tbgSGGtK1WL2UImDuw5/FJEJhp2ja9ba2t5TE/5la9H9PjSuYs+/ir1
tzsAjcQ/1UFi2E9D244ihY8eqBsSYIyA0DRbs6Wi7OXMTpy1bN8aUB5Ss2ox
hwRFDDF6GK073gqxSgvEVWMDd3IezkHm7i+u//eF1JZKb2RurO+UNPgpI6dg
qnhPznlHQxk13Kz3BvJP9FPWv0iK2iC9RJNR6OqAGaDNURW26wP0iGyclxCf
dl/i5huLr3kBsgu+TlwVEvp42Da6zwLo93CYCnTinKd/JWLY96DGGPneecYb
VC89rQ3Gs+1jYG1jKA5TA39OFIOm962z4rS7aSY+wQ7IweQ8u5tljCyzpaaR
lFgtX7P26ud5K9JCs/WlkuJqj6C2jFKBEhIDm0T3R+NE1gbUh5KvcFoR54RO
97pr+JDhFKNEyuJs6sMGOX7ezX/ziv2OKcvR7oCrompJF0h4V5KHbKnMVQh5
+sZO2v/upJkskIi5iOciLS0+/HY+9IhvmzaQ8rDPNPWrB3sGYECLooJazrqb
dxtcpejKdNDI0BPxPsJ/y+rEOzWxZPDBHupPzLECUwuaJWocz5yHHiLxlGMA
BmKEiZR/4wjy9pLSfiXoUFfKTyJfv5Yi953C9Y9h0J8X+rEf04yKUEKgQ8kG
/SYx3InGz7QkFMbIDKheLVzaw4PeN8euZteAu0BAfLiVLoBkhvCrl8nyBA4l
pshw6auLduHBwHk9O7XI0tkdE5T2Ne//PRC/h2lm2K467zy0kfNRC39VeU21
SOOc3BxKb2E7pil6qzScmZVeu7G7XyI3RUSNSI5yGCnv7FDDhRXxAIcMtvmN
U4KZ8seZc9BzNI3t+oZEP+/EbO92rO+V0FLVmnMbAcSPhHUI0cI/ggsLdiFg
baHHPPNpAoRAW/9Vv2euaDA+uo85JJRTpecrmOTdAo9Cbw/L1ZdKM7rrNC8L
Wz+LV4Btu3RhxJJDACmh8vf4Vv/LiXRLF6HdZH42O/OqVwVw0Sz1jpcxKTi7
otr7jFrTLSqig4vmMesprnM8qGn/q8heLTHj83CJsnuNLoidgKpdrr3Fyh5h
mI5i9+llebDeXehZZ38Lk0NXTgT04tEk4ci10guRs1/4o9M4Jn4SL2JGOND8
h+Ry+RPY7rKJJ9CewucrZLHYRZ/ejkMVOKQ2wabBdVSQKHKun3qSqFXKgdTK
TvlK4Elfh5eim/GQ4DI1x6ZDjvnn44JcNkC3stUKaCyN49XOfhtcRdCCmKPF
jmaM/lD4vaiFdZYWYzCcws9mOHqt5UA+AX/ywIg87CL8OJRaNJ8C3MVBa9lo
3o8aFVHJUKTCXBGOOoXqG9TSnAdVu2LuvK4HqDR98rmTycZcHyUnazWfwd33
hm6KgQ1BnK/u5w9b9NXR8GlE53SvCi/5RDqQyCgoUCrYuILXLXZqrngzSZ+Y
n1KqjCpkO7Bedveb1chkYQwKt7g5zfsLhzhlUou0ASagSWB9L+zOITJfaF0e
kAbaTr7RdVT87kawJj//kQEso3LLY9QWYaw1MBUWDo1DPMREwac24FfQ5Wsh
cRSgREeHRZehzDjYqlxvHlpFSpczIhMgBL44fku7cYGerWSczlMg6/Ro7OA+
doAA5XlmqdSQiwoKneUo0FoeAl6A+PENHTMhcdrXRmOauXAJZ9RkUMmYaQI/
lbk4TEpGmFVmUzYqkq4A4/zwRUUkuOBIN/P9Y4Ys1o0RbnYHaWAgy9m5/buk
7ycGVb129tbX6nMNgy9NkLi5SNQofNFNYUNEqFnip/RGhj3gGLN0w3qUjuTT
hGF2+mFmSqYSOgeTAY0JoHVpvu/1sYVjEuZG6Z7wCuvM0rIgG2VDbaicOC0Q
lpOdSQxtvY+3zjq2mi0uin1XT8+MU51a44gMriRoYdiQIreTfzfao177vh32
cEDKkgnkZdwEJ/Qi7mNasLTKms4TV5+c5VKB8G5dnqIf9MXplP9BK0DWKTpY
npWEoNFmcbSuWas+r9dgZ6ehPMgltUMTjTrXpEEnInCZNzn+YfLB27kDkf55
nQ2dQCOwFhCMv+WG/oT96k/MEyIeO90qbTQDtZQ88HU7WR0kXJjsk+dk2aOV
7/XziYtSpuX9ZoaHbgfwLJQulqDyJHPYGR3AwhaBQ2RYH5d+fD4FPXkydHPD
sRxHR5sxnjNyd4Mw5At4ecFTjI6V9tqT7RO8HqdzLZYJIcro4P1xc1o+a6t3
ncdioT3mOL80S5uz++PEGzHrKaSMlnv4rPe7nDomgV5bUrc0hALZoyc2faue
khDZziw0frZfCOZoVd0rbGD0AvdVbBqh0fZTBiqg4LBHiQecRSSI8RSCguOL
yakVMKmOrQzuYtyri7FTXnkDxbqXjuu2U2GZrdV8lGwDtJAEbDSvJ8p3HAL4
mQ5YS4GFrd4CIqEuXJoIxB55uvvQFCp6p0RgqDiV+8x5kEHUOA87lNAZYr9r
/Nih27p6dYMuU79/mzi7oN+BNn98xbboCneJ+xe0G49SC9Kydk8K311Gv6KZ
bYlzRcNHiUXEqPFxRBH4FbfoP5tDnGGvoE3oFU29NSQ0Zt8aFn74YvvooI2p
w39zaaHB8gKt3GxMdLw6xAx/GCUOws6UzrQryFKMt8smIKIT6sv2rMq8taCG
NNUbOo51LC0NhYUmeNrPfLA9VQ9w8DC1e+PReGGlBCpxz/zjbISRedy92OyH
cMrFZwLXiXMGiVTGXlE2EZStxqYQLE0uzVC6zyou7S7ubBXJ0PBh4zl3CloY
xWumWiM6Ill7rSJH8oBwozNEZcFCO5qKFqtsY1Z+Fpum31Ox1P5S7z4D3YvL
mC16aj8xLWprkhwO1V+NjWN9QF/FQn5ESJVJG78s3Nw5jicM2lcNPWixKs5i
uDQdh+fH616P3yzMaWW5qfRzb1E/OLon6fh41CYTa6IrVKSiUHxXFiajDJSn
AKvRo/2vEgmDw/jaTutia+IyusxPLmI0eRDIjxD0U2a6mKnMpTh4P5U2t45B
pZJbKzDH7qT0xJZGp3fmHxYCcgN6c5chKwV2SmhHb2Rc2ZTDOnRhSIoQ9mpu
s6bT6x4qHNpjx8OMEieAqxeGh/RTXfgSccSSInEQVWxPaooKOmKc3YZFbVN7
7NzfEyczS/L+sGePK6zS2jgeKFrPCifG1GksnYPtKCh3j3bPuADopCRRy7Kk
C3oujCHxNYqqNU+FK8aYi4otey+7b0CVkuKAWTCYIpqvgRq0rZXIdFTQ0tns
cs/XBQC/MSZBP/zKpvc9XDgtu5/IMqCVqR5ll2vhacbkoHZ2AYyGt0UckiaB
uPWQnFJiJ5o4FIeE5OZnwlf+xtClcsE0IsNmSrsojsAVIyDdrhMVNIbLPjKm
dqDIHX/qy5nj6n2OiFDuwkR6OnLm8qneeIBWnNPSdla6Oqe6I9/82OBGzayX
oyuN3yMORzRhPXLsNNYaHRB+C2wmIC35yU02Qq2bGknlgFrcb1ZMA7XvrOyZ
lsJwWC7YP+SMSdEiNrglggQxYRmV3PW+zE/IvPSA3dkn7m1zrm/SY4SWH6DL
9T4athbXNCmzfmdQQOWTW4tSSKvVgPtSQFDPgBC91Cod+2Vj7Uvfek6TTMaK
bY0XqEBDWRRnhdwsdfKTytF8hHkwiGHSrTfTwooD/h4zaddHBYiuNWFwqEIO
u48ZfDyYPbYA2saLSvoT1S0mXPgpeBWuuVIDipA9B/lRsVcPrIACM8ZExscW
GszuthdSSQnMsgVZxXuzrjYP89XyEsihrJuHybnGVoiv/JF/NvqyuBINVkT5
D7FV5hcTp7i3/44ZvsVYoVQTf++oRVpcaY+2Lil22OtWO4TaGoBA+eLGa2ME
uLwfQvTlPd0SsxDBSl4tXI1NpDPabNNq12kH8aUZZzJC8Z33SCDlh9Gq6BZp
Cg3hE1ULHllorXr/WsEkJv8eMqvfVbbA5zH+l0X3tcBTuo3KOJEowo6z3RIQ
YhFMGQLbE5AZSJLkDZX83KGlGmZzy98tzEot4TDMhaTt0XfN0jrkCIJWIYgz
tkdxPlPDGTCYzUBaLlBEWZ8TXyERHGsL7AZdMm46iV+pQrYmT0WReEO51DGR
V9tX3wd3HSe6UDTZNcR+es6W8HUzHGOHhu8HiLwpYIUlkmAoj344Bfn0aUer
H0wGXbHcfVqBCMShrNvZn+4Us1edRerp4lb75x6pds9y5FUa2xCx375Pygcf
FVvKMEDDHMDoxfVBGyMpiVjrbWJy2cjrQkfAnKt3nSm7m8w3fiM3X4aVSFC/
CHaVdIMbwBAUI2ac0GL/RT7ISUgWnTmN53+c61dCVKVeP2cEoGHjTAcFqbPz
nTiAvJU1o9YP+53l0Rv+AYC+JWcMi1IUKSpm9b/2OsYowcVRr8bV/LVr51Os
Vl918PYN8lBPORpBzHrNvIAUPKzV4ODhCgq3XapvWU0na+jB37CVQS2yCKKx
laDuh6eRn+XaJldPS/1UPJSCYNf+Qbdsb5xMINrHLmRh4KLVjf0WZetLQqq7
EBxRb04DJWGQ4ubkMrSSlOzRhhOqk4Oe9y7Y6byVP/a3UkgP7h89UYZ7CFxp
vcSTk4UHYj2p8QecqjDMo4++kWQX3G5FBamqqr3mtLlk7w2n02fQD6Tt4viQ
PAp5BE6SYZdcjepa1SZCks6YPcUHopkMwoTAnpjZvKFw3cW0XcQ4sNzaenpN
2cGLbQiLySgfpOnmNW4OsoTZbTaQEtuhSR7JhyqGN3IvU3uLsTrHPzziJcve
jhBa6COZYGVWhCgc38R5+aYAtOzb8setbMMPb1e9HWg25N0K18jPME3EhSh5
EcQ0RjHdwv9cuJBXsqV4B1enXvS9BUxXVF09EqRwffwMVftVHiH0jvXhNewB
TkW5phpfQqryEm2XYanJskyoah5yh8txTG+aI7GlLJx4wTNVi6FUgSf4pM4A
HFFgmBuCY00+8gIln3VJipMDt+j47VdCc8EFiLM15smVLXAzsiAmc1BNp9KR
nhsTAf0oepsGSc9KRRFhMqeGC2IA1SokG9xJh/PzLKUIVG3/34YEYBZ1D6/a
r197MxYFOU+KD2re+ey3DEMKrkH00LVe7ScIkuYeMM/Ob5Mu6sGshk937uCC
R9k85SB1Ux0wGVsxwIEPBEVSJOlQsAUNsktGltCdIEuOgiTLyMZYD+wG+T9W
GLEBqOfV08j9aLwX4Qyhfnm2mNBA5iwPQdaXoTXjwQ4tGPCu5GE2hxSa7RUl
+KxdZ13YzWqDiokuPNhlsIR1K0p6SXdlKPMkPtkmyYjzy/tEsIvDYu47+04k
RFvRBgHJcoyDA0EsmDwxZNSC3IoIIzTEppRX1ol3b5SGg4Dv5sYLOMC2o4lh
3MGnh9pqEwOX1UthKca6+QoASUSmxycP/7Nzv33LjCSIYZEEmY0gDFUbAGAr
bJYeCnjpiVGxWqziG/V7gLqqpR06/AV+Wyl9A5yI+csRZXIEFNnwI/QE1bkp
D43hUt0Izo+9BW+LkvHGaGoCvh3b04njcBPBOf5dOVl9hLCgUiPXX+2Y5YIn
V5FEa0zxP82/aqvY6+AlocqRRST3iORBO59dUB/hAhOOx0rT9khaGgkaVMS5
wkKKnjZgzdrit6ymlcnVPaEbNzm9sxf+ELUDz/VPbaGvvOkixMGYV8O2z26w
qCncHzRllc7EXis/T0xo6g/eG+M6GueIEQfEM9sEBkpl+iw0FCOVmLAdQP/n
zl4Agm3uKh/YDSD8VpSG6gKOPYRIsJWdmJsBC/2P/c3Wcc8krDeJglX/IF5T
xl6jH3mimNX+UJpFk+nwKHH0vjHSA43hnnTBfW5ms1LovKt3sg2AxnQJLGu/
4fPvZ1T09youIh+uO2/v5MVrQCgnKx2Ixn3ZKMWisa+TfSy+y4Fdm8yaI9hj
8KMnzGgw/heBg+EDA5tmI9WW38Gpsu6/YhmDkFRC3E/rjIkX1NSqk+OcjQSq
N5F8qlV1jSqd3IHtVh1GRYiI67KSvRg1y/XYgY/7vh3SIrq2MTDcJd3QMl/Z
4ghVe4WIDGNu1C1vR4HTdHTNJRtZqq+uGLPddZQUSmQ1O2C8kzFS/vmPw4NR
FacVbEc4zoHnjbYb71nrMMwvq6qyAORwBmAbECaxwFcH0VftzwYX4b3PNhJv
RieYwwFyG3gbVgGSlDosp9HInIfUBRB5lWXfbAl5UOlrRKqBT9wMx2Lia/SE
dwifu62a/lrrSvfvEOMljoURsNeCoI+7sjNDWNJYHQpQal7cNsvkImhqAMEy
SQOH3JXQy8vB7akeUq1sgGKSuAtbGdkMzwhOWVo2UIIOEbSF/FO6a5l3dcgm
SqtsFGpULYVw2dWQKiVWi2LXDSkeuKD5pCmrfXNqnAyhnrUpjkbsj9VKt4al
oKihY8qVFFpysLgCDsETKW70DKEmYfGJ7VQK2bgAkLroRifzWXYmCjs5Na0Z
K49ZzRy76+jMR/TrHoXdaa2wJj/PK7AH3A/ZTlKZnB/FEALu2RooYLqqwAap
hopbIxxBBF9F5bJ0RwZZ/v+BaWwkyO2HyMx3aKof8/+rAfRKAlgs3jxnhwRq
OyRfPfBxqSXaoK4wDI3LqUqS/KURI8H/Bqjw1ApFCXAOIJXlXsYgLda8t/Ws
bN5nmtpgQBL/jJMgIia5qbCiVrtDBeK35nkW18HAgvju3vSroRckzi6l64tQ
x+62d/ro2xSzMAmJnGPfx/6qWiYMb+xLzd4e7O7KDfey5LKCQd6v7b208ZmA
jihupFAs9et3PB1slWYgYno1HNwWFnQwo1LiKCIL5oknN27KPZTECtpCCQhM
AIaZL7sfsmsEF8ukueioEdpbngNwm6NoYb+jZ0yikSTboI0c7KDLD1HV/KPT
3SfYi56VuN/agtVZKSMzrcGTAHKAC5DoZy1OAGKHtLMwKAufDDsCeDiASPdZ
b2Tf809XEgodUz76NBA4nFN/yeXh9KUE0vHWHnKbLSwHKFLWVvtegD/ESXdR
DFKW52clC/wiXIjT1GuSX3ynUv7Zmf/oXL9ESPWk0OsUoRSqqGUo+HY5QH76
E4iFC6WUhoSJumcDSi883pgmBWNRpi1fZa9cSB2cRman1U/3OSykJ6xwV3Sg
Cw7PdxIc/6ASJ7mQQKxQ38R3lUL/38BXWjRur+GQ7zbuyfV/JBy3iGtqHiHN
qOULIjqnPPjn1AhfFf59GlqHAhOqP0uTi+i9Bs9Nv1si85r/ZlBFqn34Czc5
NLFscyuFQ3dR7goTWWTy3pNWoAwu/3F5rpGPP8P3rFskZll9ym1wi330HFpC
U3Xr7Ljfs0ibzihSJ71pjbP3XsGqaw7zpfuu8KVoV7IjWtM11acNQ/PXc0li
3YDeEKSCuRTJi04maq5aaf8df8Va3SOPKHI89Bgztcm/rxXmk7c8u3yzkG1H
r1VsCWAj0CoDOiU8oJ+vfiZL2LjtahGaO1p1fA9Xabs14NB9eHFs7/7CBBx1
S24LO3me13tO4sp5PZwNdlSS8dBqjhv8m6/zko41g7L7VkXPxaZ1eCAYz6Qe
5xVA8yThSlwU2fl6vywGkR6RC4t+9UnpjB300ilRiOAj0Osksc877ZlJdU5V
rAMChJyMBeNC8kDlz+quipmKXePzbk5aIwI5UYcoNnCgVuBQrseHRxjl459b
RqVp5fa495cW5SKpABL6yNP1fSkNfj+j6vQOqEnFtMeLz5PIKeO8KTzekXDt
t7rBMpT5GjocBKklD7CaLQz9r9slxTmru74iHaMdvL+wUHRkT/qkxah9WQJ3
iqUIXuHghxutXS8syK3RPTIu0JHSF59B1GIjGplGdU++V+XOrifNquIOCNxu
pKv6azyoMKD6E4oGgtU8+xPGomjVXEAFgLaH6y5bPWZIcgYfaudmuGU6f+1j
ZEsOKjsExpdatsWhnyyzgZ86sjcd1vWaW0zPdsluvknYAell0E8klHRB2A7E
kamK785Bn1jiazRtUmL4JMd9PYxajWwujwS/UaArleC5tTX6mSBj6Nc5ORpb
q3oH/idnezcGOICvox2K+G9jGwtuUyRaAoGc8bMuU+mXheMePH9p9K1RrW3c
i8vbgXBU0c6pFXGAZN4e17fJKDaohytECnGxdqgUGQhedDsSoB7NYU+w5E85
d+J8PIpoakVfPBjQLeU0WY67nsG1gJe09jzRu5tfDOJ0rwUxu7bee7vitY9s
3owKrOMzXSw9BoMK8eT3oqcgm+G4ycqeLft9Hor2qqywV0y5bej63b6tRGK3
wEqxX9WiZx+2255u0gzxFZU65MZlNIqDwp97sj+OmuijMdoVAorgnhvFYC4c
MVzkI9lwaTMNazVU+5RtTX5zlnpSq2mD/a6PYLs/s7z8gku1fK5KXFa/DkLS
RtCg2BUfb46rmDgfjvz9r+r2O1+L+X3I/ID4xdNPLau7HeBNm6Eesw+r5ciw
iow52pcDNwS2RHkHpEamryCzF7tNYEBSMKLb6jgSGj05BNrPAnSl8iNVzvNE
AbblKgUUQYWMvh7pP+3L/YKXNlC7AlGqIQI8fWxBRLH9khadlQ6KOHwo8sI3
GJNrUWPx3XJCtb33hNTirrdVHgXbAaiXMr962pPwyzrrkHS06Me0vEXDIBmi
MCC9yPK2IViwejRQoJ51o6HdOiPJEgqhH+hkVNH+svKVpKwjBxc9v9J+8Yf2
XjREUKP9Ogi1WOg/ui7xoyQOC22nSDQhZV8VgxiDZQwybpbqqxpQ17bl1y4G
3AepeJZS4Zp+jYo/9HJXj6SUbBQZG/TBGI9R2PJnVdt+D2cEQX6EIhGY4srr
9YGSe2fZYAzKz5NfDHdgUIwQBaaVQ2R5Q5mZlzPgYXRNyDYjkw9uIaKWVDM9
ybNNerYN20VLax4K53Jh4r8sYZNevgIXzY0NWRO8yksdi3WAhc5cNpzvjCp1
y+Ckqx+YPZ/dsnTgyodZfyRsY+boGxhOtxInGxp5VT8LlNeV12pekuEEGGCj
U4VlpBfjG3mSpUObpdsiP4w4oWt75YjDZEz2lDMkCAy4YGyfNNXSkdZIFiGQ
o1leijCCtV8IyCdydTDifD8P9Vv0FQnGnV3RsRM8qg5pED/Yb36qnt80Paw6
vG1gVpyCXsc8qS2QXH1+W6HKWRo4hDUE2Fb7jWLhFeKdw4cDvytd9QFDgZFZ
tgqBYQwGT9zkQaJhlI7iQ6Gk8CndvJBfIvEZmdQNvx8FZrhuR2rTyqFAlRgd
l3Lk9jzPKW4FJHMK2FWfyCFnQNIXodO9pmBaJciEGfIVzAM/cMx3LiujaULC
GOslDt6hdpTpDvp7H4bwYKX7M0zfJxvnd/HDyRw3I41BCwdxfrMADV4xzu4G
hIHLQssP/MPvatekCMXTJI5DVosZtPQZUvBHSD+FntQx3Tk5xgFOz9D/v/Hj
ZdHOx/Jx2uwGilqXRg2exj7WhMdK12DYTsY4MLbHYXupSgOG11JJT7HQUqUS
/ldb9HSxhDtmlBqvJ44ypyi9PCDJmEZoI9DXJ6MA0NBQX9WFk2Ritb8k4PxG
TVwasNG3km1V+ETU2hE1tV1lwjmFbiRZjbT6IiOYwKtU9KZEshSv//k1MYg7
upIaCYaNl/cA7KHPCR2axzJNh1V5Bxq7DyLSeh5KISt3bPgvyaOBxCZog8Ax
tQ5PhEU904JuEq4Ld5OIM9FTVDjUjZvrBhx1y/b0UTDGVPxk+3N7oz9P2Yjd
v+1LhLIjFpE0EOBUOaq1A8GdKZe6kIHt9HXQ3JEJ5UEI/wTvx4TmqE5QveFH
af2iZ+w0qXIu/r1/xdAnh2UDDMJ+0P2dUWSm0/ywAqp3EJ8W4jtCCVRYpiM1
tuK7ImKNlu2wjsU/i06YHAql9V8qjatY7p+LheNyyVydTF13SMQHXdrv6Je0
ONdL8R9y8DL72t6zppgoFgprzLjKpalthJRc13XOrBjFZMhZs11uOEtIU23k
1YG1vE786zW4m/fWufpKaUP1VSm2XfkPcgHXkZKQ6kZC5arCrJGp229E744E
is338nNczpEcpwAMuqaGoUgbzk4lT/QUp6io+8JhQSkI5iedPhxJZZEnL5nN
Peh01DcJZQDgZVIELqJppCpc2Qc89vuWurPY0w+l6jNJTfOFaieeBKxurnwx
z9p/mDhfjh/eJ4JJveiPDt9tcNy/0LMivJel+BvYhb82dC5qEZTY475NwmD0
1ZhbuEXBDfNBaowQx3z3xqUKp2/RmMpK9/c+4NAx1VA95A4YkCyG5IeYvkIS
/yYgx4c3japU4mC7goIxKi3BuTN3WtNhqAyZR5WK4Z1DPJ6zY2mIp32h9bcG
z/pEApzDqHAIZgN81ZDEgNmcKwQll1HUa0rkW7Snvo+aZsj7qU3bMb7Iq/Fd
MSe4JeumVyN8aIOK9n1kb+nrtoy4AzAO+ffzPERMqSCxL8/QGT3KwTtaw9gJ
cLp9mrQFsJqG3RZNQxINVZDDhDcebKfpWN3caiv0I6CpoU4xe8PbjgAaC7IE
d+eqDDLPg5rjJJEnQoxjTIt431f2nq8EcvlFgk3ssg8+3UTWSGvifxg3WOhG
kcmgxBvQThJMjxsyw7Sf7uxQ6IciwvuE2A2hPXqpdnDlxWwvXNt7b5/izvVN
bt2a8u7Bhux3ct+Nh6yHdTZbl9h6f7MiHeBSJVRlksRuDYOVc4HcxFfuJW+I
ujCGeugxT0JKMoLwAJQ7Ug+vW4+kGEYpLW+bcoCNtrJRARxQTTr/+gOT0HcQ
NB8nikhmLrZLh70zpH6+mKVMZ3zOJPbN7Np2s1s9fZB4RYBXLJ8sRYlxqtLS
oRtLGFEEz487jEb4L9OAbf8hRZNK+u4gwAcRf+qSdwFQtA9gPQCzaZ+odiMV
GrSbRRO7bDi7HP5oOFCiLQQ9OrOgICQJ0aVCadNSLXN8nW+WHZXdGKXctWcO
83L5zJu4HZ96fVX+HKcnk9lelH0oPhmwh1Ipn2FQCMlbVQt8Ezj8BrzECsiU
NiIZKi3QCB0L7k0ffQR4/kuQPC1me0Pt38FM11sTOb4EE0oRzNLNoqD3Q8/G
KKXwR2z9m1QnNmAOdIUUKo7nDUTEMr68sL+fXh10YO3CI1yE09TGX8VfvOxE
PxdjC9BfX57E4KpxqoTxPvbMhHdTxtLsBjats2PZRaHrTokme8dm/fAZoIAx
r60Ypt7j6TzRytms0Kp8uGi346hYa9ksO10H7mTo0O3yJapSn7soKs61QnU6
+YwLF9QVXFrT2+qID8uzyVII8X/w6giKwi7pwZ2ASYOdNcrlIlp3L/RIXtRd
iLqIJH9arLqJu5/BnwHcy1SFz6sXYSKrvQ2df9/+BVtw7YgDiTxo1Q532zQf
0z1H5FchDpl403mIvlbmWh62UnPU/afYOBufHoF52+Arx6I8429ZNc3p/vtD
1lt/CyXCZ4+t3kytgYsUCHcWpCnqf953+U3QwqZRbCxeTFbdd5LUnY+QHT/R
vyEfn+sdT3h1pqxsC542P/z1KkGcb7BnpMQwIYBjJqFG3S751Ka1xzgi5NDx
CHvuJ2rXjSKa2J/BFtDCiDfLoozbaDnR5CNaCHCKLDFCmkxaQ5JLI7UQwi3q
z0zO0RFpaXSSRayBuElNOHXoDvmULncEosF6ZTah+qlTu2l7wjKBQq91I4h9
vhNvbUTm6BgeSOoodjdElzLCzSL19Sdix6rARIWWw6q5g1zz6MWZLOkp6Wd3
DM+BX0Fd+eiZ6FwVik4nLDOHcfIyoUefUC/otk8AENaEZGjEpsMRqEFumYwv
yezh3vrctQO/z3jXFjwDNsV1ALgWeDSSmOU52InZQtC4ldX84MuVzuOF946N
MJ9+DX0/niCGR8gNGCDTOKyismb8oMtI1yzNxNkH7URDb2MZETkSB7gRtJEy
AFreOmuYVSehGcUzJ+ur7mWM8jNH500MQn5Sy0fgj1i0yWu8O6KYQDZOGRZF
n/I0GoWbwkp+yeGCYw1MLnJK1A3oj52XJ+8eBXbZS55XaFiyzRxKGaBJoQt3
4hASg9SdYGsNbstcgAjtZa+oSORZLmsF6w9QLWUnoN3mQgAEmZITLUNKdG0x
PziWzBdLzYcUaRltsOxqf8J7DSAIlYE52G9dbksSE/pMT5YkOyDnjbxO3A7p
lIrvzvxCMyPfaALWv5Ce5FlbXIBj7xOtniB7bUV+31rAGyOSrW4AMKnnHlI/
KEVMXUepVDkejF8cyMghvNECurshUeag/+cAdlSeaK3qlW1KF3/e2/9nd6z4
9g6eecZg5nlObNmgQ3efKQmtZRqxXBGhHNLgRlmlWJz8CjU0oJOAWiy8CY5a
yTHd7seMoUkJEFxxasHwAPxSO2zuKflCAAQDDAhYkaDf87M6VQ==

`pragma protect end_protected
