// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
YnUsnMKVX2fQwgxn9+wmItJVxsRL2iAClP7CfD6WEPX/Zij/9aORAWs8pSicfNrm
UOlIVVdq20a/u1okw4erIlLTh1e1gpx0cnMD/g6my77XU/pN++u4YFhKt0tgujTz
tpCEngYrYZmLnhowaFcQgSb9iYfPjNzgp3BWZo54SG4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2432 )
`pragma protect data_block
7pNtk1ZLhE8k61N3ekf/2fUyzYswDr/DL7Ijmbr9yVmRYSpieRgSEj8MBTX7ZdrU
Lv3rH0piBEWc6OTRhQ/hzyQKkuh9K6DnGD5cy/d9saSfL5nEKGSdxqEmLm/3DJ3j
w+1IJmiBOlg6fZhXFjghHFlZHieSXXXTe2dEQf2suGaVW+4RptVT4lCvEUSRXTlF
wDU3797U82MDzA6zNkA9XZUFW2voDr9G0UvTSglmTOLKq/neZxWbkxkXmKejpNRt
qjcH44E16DQhV/kp681ZaAit4CGnOMuQY1yk1c5O42h6G1wLyNyLqoswxReWeiuD
yMeasiiDhEbuBIKBp8reyk9eYcjVM2pW/0mLxxJ98Nb6+bHll+NNcLuDLyQ3BND1
2oLy4xhEsHVOfJ6KCOScxQ7m5sLh6VJTRgmjW8/r+lVBOafjiZsQCpMP/7HuQkkN
G1Qi3FNShZcS32dhujZl1gYadyi2o+fQxPMsgrLmSCZoRXSR2YJWTZcxInbd9oYn
3/0t2QLSOGmgVMznMnrdnSJVzkKxebT/waZ/k1LP9U8/Cmv8JxNIlnmkx9MCU/dU
+sB6IdWJ2IB4NBy4DmCTahOh5DPlg7Embehy/OU3qlY/tjypFq5xOHcDms+x0gP+
xK70MKwoSeJSpXi9FuT1yIBLXq/5A2yh7wdlNZxTLwl4rgdp4/OwogZIkE7Hw+bk
R6reIf6MEu90wg/blorK63ETZKZkVxO2EltRI3M6v6LFX3FWi78EfFU20Wq6FZXu
61dRtksZaeG75WE4TBlvvAy3zSBUy+DosXesF62Gaq88z/n5iZ++/xSzGwt480kD
I/J21+vxfkuD6xONjhOuIAjpQPODy9k2QieixLkhiBcoI2+0pvR+qP68aWH8aGwh
CVSvZifLTEb5W9YOzkXScgstN/X7SlModbvyjL2ZjIaCRYipgXUpRQowaDI4BNpl
Clv10vv46RFE6/HmONzxTH2sv92ac9xiRz/rOUW+PoH1feLkzHfe9ET/lSiQzy3C
4NvYuXXcJQnkesI+uAkxJmy2fI14SnvIjkAQwdRII2zAOoFL/EkKtt5KIIwQ9EYE
LNjcQbf8Kn++2aBaCU+C75itQQxNtcmWMsi6hVBXdOoyWG1CG/KjGa3RjTnkCCN6
FlUuFyxNzN6Ql4nwKjAXDU+BBt7bgNhPi3FlBPL4aYC2+ju2ZqARexyioHDhsSgF
yz+39ufCemIUZmLJPtSSearSSw0PWpub/FCrPJOQY1cYabQtBy2p4SJLy1tS8cd3
02p+qK0mNqFqKACirm8j1kBDzv0Xwf0m+o8PemKj7GssxZRmbNHM2xaf617RoktJ
snkhP0HBGzQ9sC7hBwCeRFfZP2H8JEhim2lnpK5e4LWPXDOKyzE/ue7ayoFYv0GR
n/WlSk3mcLWUr7N4byyzX2GDCKcwd84auenPRZjoY7zNxYiknGnxkNgx2kw++pRV
e4344ptxomZ2GoTN8l6RpOFPx3Tv/9CSSQraYp1LJFLtW2Yq7lAAR5ks0iswIm65
QI6fmiUMithdsR7A/iJ+s111CF+AaPA8jD0MSo7abC6f46S55YsC+de/nXF5JMyW
6N2ewAGySA9z8QHwhB/+nIS2iNLjgqQ41GMd+VwbKHjBMGCiSKbiKthBioNxnlGF
vtHFV6qXBBxB4mHjJXvNJNbJ3fvc9ZYj9rH+vTGWfOc/ElkH2d49Ay7nKFe1Hyen
tgWOJZc7My3ucoF1FPeGPvUrA+26l2+GuJLLWGLTQScBSaBHJs4SCkfCKDvEJoV0
hYAdlVXMRp+tiF6F740fIOzp7DZ35iAvehlWaOx/6ndgY5dcymPQOtsYRAq67wYY
uqQKt+Vde7G+DhKO5FWVeSyxqV8Dia0Cf+IfdzwvlYE0dGm1+VE8721Pm+QF0hp0
HDUM1ddJu0DELwRlLEf0ivoqyNO3nBY0DoSYlAotq9NPVhxLxyMoWsnAoI24XJez
he4Fp3eAkX5cu368qt8SmMWvFykvEXIeg5lZu4etrEmqD+5TAvDfcL3LrNf39pfz
MZG0IHW/FvoLWCoC1tPFWoGbUCQpQARQx43O95fyjgFi8rXV6WidGDwD0qqWuQuZ
FA9nEuCDaBcmUkGij9xdYbtdvpsFV2BrLQCwJoudZN27NEl8WZ0tXPXMn3eJZzfG
gOfYQ9EGfC3hs88FsUVgRwQoCInQUeu8MPErWeHUbwucYt96PBsDnPk136iFjCpF
RsSaxwatTVlSVbpbzZ7jUCuS7/Z9kdKSt7pnr9tTdOFpMxEg2BHBT/x3T2/h8ulB
FAOOgVuk3eOHfgVgosTiYjxEKPW9XpPF0ViWRqREAWLNg1ihcGjsDHxW4og5ko0v
Xtqy6Vhm9ydWh/jhABu9EsFVJrWXM47/Wyc/LCcCTrdT5bLsh5k2igXbg5fIIZ/4
+eTCNC1kb9NXfI+5fq+l/k5KBG7/RICpuotRj+fLbWvfvPFI61h3nSQYBrEsVIcB
4R1cu52q0/kfEfYU6I0OV276ScIOoTWlQoHLovTo/AbZ+pWWiFQ9sETUR75et++d
UGKjs+8XLyhglGNVna4nGXYA6drcVPv2zp8zwI2fec29bdjgNqDKPKU2MQFqlYhw
70ck7HCZDag95Wd+IugRfe4jttA7ZG8S4IaJjFVj0foV+avQRHFNs1cMzIZdZ53d
ifAMfyHg6kSciR1GwlOosfrN9wInqNOpJtOSDfI5R99KuLtrFXmewhCbsiRn64zF
wMAG+ezAZb0lezMVXBY6PqGCraYLbTUk85YDqVCnTSJ4pYrcDj2KIaWhD7cAfLiJ
2XOLnKv8FpsM8jjoy8PpjBk1a1MeMyHUvhnVP9ocEyilPHdd2DbFf/YiGKks+hEY
hBYrHx9F907BhiR9BcBR5d8uhUaLueVSOtG3fbd4btWzs75ROODWlWlg5eZZbFUd
lWi99NXKS20qLAZyTUhaC69KpK7zZtBQ6HAdFWIuXqYmDraGFpEglEbqJyzRLizO
hJIDrv0P62ux9q0qDyyWrwpsg3BVAWMwA/ixFk30IHQ2I6vkGA6dEy8QPOEIlgTW
Wfg3kff6gqvtFGJbQojBRmdR9dVPb5vLo+MiqkWkRJENhEZCPSt4GCpvl1YgexhJ
m9aXPo+T1UsMbOvAocIzNtoqRqmLyJjYuqFb+MkqDTfMeQbSlkmFlinpyIF4euXZ
iv38/JAKpK4Hwx8Gw8bnPJ3jLHg00kln7dqpGrsETjo=

`pragma protect end_protected
