// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
ES2eyoTx7XVXhcFh26lglEhgmRZ2CIqlrY5Vn8eKDzznUE+XK6tEqsrHADFGlIOf
Px8hG1CWPJAMIQ4d9RYOeHCLhkoA+bYDzsMoaTRZkhop83HeKrYU1pnB9UKMEKTe
LLtD5St7a8l7doj++VaHWU+ZoFrO7eSADpEN2ZxvelE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10000 )
`pragma protect data_block
Ez+fIR4LfF9sNCZeJZLzB8KW5DczJobdukBcMAeLAYYz+cgPBWTHzoeFNCu+1HZY
waKmoEi4zK0rUt29GsSI+h3ry1okPyGOI4tdi+MvPR7x+gLjgJ2AZ60SSFxypko5
cPqqYP/kXUfVdcnv24npkAcnFytXIQvCZDg1E+zzox5uQwfIOKUt65ILHAbxp+qP
EFbHb54UCjkQ/yaPhWPYowKPgAcucCGQwzqYGugk15Fb4LqEtnhs8VkidN+rG+mO
2ead/6BRpjdBfSrkvqBFv6lZsBgUQa2IGen4sO1okEm5SHaVS2P9xFrFZ1GkgUaZ
uV1YZkLj4YjH0c6h8PulVAtAjoLb813YMj7jLZ2zASOqs6u/9F+nArDtGOw9l47C
T5P2xGAT8x2FHiPU+rM6Shg0TUYNB8qC3o6NJjNMnCaKGHXrRbQ7IT+6jTSlhZlv
QQJMQJn94rMgo52arSZJEcpxTa5Rr+xQFwdm4SST8ZKjoBcD64boMm+hcn2g/9lZ
oolP5Mc8sVBckH/iftKwAOB1riCH3x7Mb9YuvM6MbhRb1wynFnbdm7c+7S3ufU1q
Sb/SI6OCkz1uRKO65+wr1Iwt1EzKEzBC9/mW9v04C40DQxWiykvBD7U3HTCDRush
To+qEep+t7qt/grCfhhJETlgg4f5b0EriCqix5oAsfb5IGvuhPbB2M5scfQSXmM9
msxoICVCqV3u/asRl8V6MI0nIq/y9jcLRE+3saMtmZC5ACuaMEfZVDDcYQkrqHo+
9tKiz+2quzemnckH01Z7XobxDk8eXpJBq+0c3CeT5zSBLQ3vF8FfQIhjFSR/kft+
+fOKfr5TuneTpD+dzoI825YfpmTxTi7kGTcOtB2kQcti2BR/1yRSZDNgNNS1j+AY
SoRpg1qX1rjIH4CUTseXY0/lz1DDsdIjc0ru4wkqmVa80P/yM05eEzvfWzYi+gwo
ime0f/4jhJJu4XJuTdFtckx+LsMYcYcSL67VsMokakrMIkPQh95+SznuM1qe5eh8
nUSpgRTCxZXyn7xgBVX/3AUo8JQ7tHxHCR9e3bleCzCafFIhXYumYZkryt6O6+++
8O8GJ3o+X6L9kGa+YD2hiwU2u6XJFJz4bAGDtyqAHtCwKOxgbvRpBK06xNRcFlL9
LXXTmWI8bcyC+VBXy8zuCcQDdRA+Ur+egr1n3WT/MPzPLfnv8Id1fYPX8qAN8tHM
ibSsTEOGERqq/CiJJDKtKcdHJF4kGgBMeNVwmA7bEAXwBf4TY75wtn1KND9j4ohb
5FWsGv4k0qT9s3ZdAFEEBVnPrKNukg/fuBoXgE2eAhNIfz1va3ocVAmSZ+MRmPY5
MIqt6igXYjG95dxH6jrVcHuy1xl26P3BPcnH2gWnkyQrvMtKgLbHbFTDjYr/byWj
VIhNfD2evgv+v8HBbhLIgVgS73jdu3hivHnXnJJ6nHrWiveOVA8WT0N3rHFSjlma
5/t7XyR/raItwuBJenh/ym1VnI7VwzYNYtt4VM5d5XBvrlDlzB2cFUN5vt9qrR6x
zmMINTiWLX8TiJZioXkjBfY5YXoOyY+ujqEpR7h0udIOg3tAgNJr3jbT/dYYhhgo
bLaNZI6+1fcDzstVx6I/OrL3Uii57wgvBm66axqfpkrCettwxAQGEB0vS9YZWeTV
BFpUaIz5Jced8zt2q6Tg6D8vwxHUPwErYxwTFkRPjs1vbIKtoU5H46Xj1O6Kc/mO
jPOs4kRGpE51o3lg7JJG6bEVrCFQPd+RZc7KYQAoadeDIJ/iCaA0vl6tZa5hC46e
7K+bRnTvPQdZTukpYizU6e1RkSd/kLP5NG7ClTe2ph4u2xvWgMzU6sstQTdUsyUI
JCXE2LR+2gABLm2fC2ETORKb37itpynV6AKJzvBzDHxqfB6Qeksa91TZmVKUn5DQ
RUXliUQej4cHH8NIAi23bQeRdBrpe11bKbueLlrg+3FpBd0Zembsb1+2HBD/cDeE
pFb1O6lgLFUsy9rLwvixyxKcyIE74BDNXQTpBpJYaof2EZg0SGHDhMdbD0/+fXcB
WPomagG2QTU7HWrv7l2Bm/aLE3HG/UOgVKYy0+yUYu6XQmUwMxpCug7iGpp5Q5+0
PzCUC0jo+TmqR+el6HbVfYzxqYFRoUUojsuHRTaQlpZMsuer2K6IcSBHz+aXcr60
lDzN0IFWIfPy2ROK6z/Aj3+nqkZFu0IRXQpXnNm/Yx5qlherGyrhcyi5CtRJHkKl
sP/B4Gv0Qka0Jhx/8IEQRubqk703q9zhkY2AyIfzCPtKCiyJgVTigBjWKvOe6fqI
ktaAwYf8MSBhDH2YzvhNVSt+5wiU5N2+gaiz5gjlylFfPXpqTHPHOMJ0vUhIqWB8
5NjXZgwCetyaGXOSH6tb4ElfGddmP5k3j9Rzwie41aJTinTkBvutMAQLyTXfEJsu
GKr0+NzqzxKzKK2W1awkLbScZc+Y6IIy2ENFSdV3m8iZCiIJJKB6LJfKP9cTMbF/
HxqKxkD4Vjh4JP6aq6tF0X9V3m5NAnmPgtsvnWFQNlq/Hg7wfM2onk0iDSA3tsA/
+o0w+B+Vb263zuWyTedBY49MKuyVjtD2rJCiHnTxSoMiVxJ22oW/dYDYEdFy3NOx
88U+YsATPZZChaG17F4yeTWgIm+qaaz0wbNyecspLqBJ+Td+WJ5SSbp5ULZmHesn
JL680NpDHpJWNeNAAaC27LP7RxakuqIbBBupgXqh0VC5kXkfBlbsILMGAC1RK2vb
79VWu3x7dMx9VXthNCIJ6q8GGd5lF5ccYDckjoL53a7K79UoKUzt3yw01Xd58iJd
MDiMSp8K61qPlhXHk4AcRnrXW2GAMCauQoE4uuZUkAIfiTTMZvyP/3kegJqAZYq9
iqoLYho8cflrBMEcAVgfcBkfNfvIwrdpzfsdUUA7S1+CruqX4kNTBHnifZyvi31s
216VEcBYky/EH3WMLOx4C0YwiME+GnFfKn+mRLlbiYhYETdec843eHQBpgZlabMo
IC5qusSgeDdbF1H3wVor1k0cY4BNDioKUVMCFcpX2/WvSW2TZLc+IPAjiS4m23wS
dw8WEWl7SxkT5YzLoCzpNGqEJ59W0gZMzEFfJxx+3xnzlfBZSa907zvvtspPQy9z
NLNUyLpRDa0Ph3dR2uTP2qaKxPh1zAUDx5mzD9VpYjiMcntiGxryLWt27X2Nq6FM
+mGHy81iy6zUrAUkA9Eow+LbgNBl+xxMrC1k26gDqjwmrE2BGSiZyjTn1o9ZjVKI
xXhOXEjuzyv70TAYYpXTvflkzDVZGSY8PYolEGnSghipdq8CfD3pXn+8Czu5beSo
IA+qa99Pq4QFR+hxrWFKBagzFbAvN9DJHTpjEBH8PI96w1zimOJOF7iv7KkXgpDp
neSh9hDpKH+RAoW+ySxUITokTDxdOU4ntGfP3P/BUDC7fzx3BLqzP+Gz/tDWpPI1
982e/9xks3JRk5emN7D5qnCLZ2ilyCRV8HTVNG44IMuovJrAdErCn+5cNpVl5dMR
IOzW5yxfYVEm3fA9Y4vcfSdaAc00di8UUj6T6urL0FdBgiCjvqzekfFJjovpUeUQ
Ow9oyzeq2Fdtg6K0OVZjQ3Z9DDGnykYskZ5biJP4ZLlfQLMVelS5TxjF61hiH/up
FuOvqTPdr+2GM6UznnU8Ky4f7dHFljEvfStbRvpV6WBolL6b561cA2oQ2BHoiOam
WJVaVjUacXEpY/CXCdVKBI47LVm58C4rANn26K+Thd86qNw9aRx0iNBDjtDM6aS7
7P0ORWA8RSDOKWCF6OJ1hXz79tL7fsKTf1LPRbte2MItQ7HkyN//2FiJf7/PvC8W
aJVSWg8DOy1WyA6w+QC8F1RjJZVL4e6xPqCuT46i23iWXPSydWj0cDG8Z/2EvfiN
skFNeFDFueX1SvK/y5TXOvGMj/lWXzHuQyE15BKFP2m580kCgYyF5c5tzwVcqgkv
n6iEbS9MDCNWbE+TKPs8vdYbKePg+5r8ick6qoGSEbwE1vrcD4MxS32udYDwlsC/
+3FtkOi9gCe6cOpO6ZamQvNpwtGxkSzMZn1nHscv2M9AERoWews21ita2kRzRKD/
+eVAHh10iVOzoaAt8CUDUkdWVAC8TiIHHR3vnGS8AGhsZmG9E+y6+OSIHNIjJ3Q1
RBorN0CnBPlUfpqexyDzfTFFvUJU6ozqvE1G8/aYggIKTaIoqYByc2aWVqzmVFHw
hQFBfsTwCQIguJD3LGo40GfjGDYlYSMsDUZHX5/3c642xyO2bgYxcFnN1o9HH8j3
RqHFMmZHukShaSzDc9D0Xo4FrtKeI5M/2vfQtcZTkj7Q90kMc6bMcc+kpXqbEocv
rewyDmRD34iAd8i+1k3d1JxNo/hJq38zzFcj/w/gy4L3Q5P3nJ6uCfZutueEygwh
5d9WqOeNbune1NGgg7fdWz2uqh+h3n+doQzBqvyIvnMKpVKBqDY7vIebxDHv06jd
Ynw3v0rKrFrZLXqoq1UL/wdoSa8BJrYe6dJZFm9VWPVqOgMWxVznlTQvO9kCvNFd
QASRHF0oQcSqb9zitAnglLFRFzLJ2mVpGDIvlNgxHZjeGlVl9c5OQdQMZOcGgi+a
s+yFN2FMpdHNkca8Eq54iLpMKCV1nlNPetynUkk+0F7q0WVrZlgPtMGfB4MkOUxP
IbU6RVT7QmSKlURGDTNaz7tZMkp3g6doT3OIVCo1VRvJfOVLtCN+5/kZe/PV7gus
WYv71gc1le/0pHcwylPt0ncz0NEK3fdqd8N5uslH6dc4R4NfOeHJ4hmff+b75kQ2
9KZNVg7/n1lZiYvrN+8CuN6MHhyqqCP5A7VCg9n2WOeEVMt68RC4NSG4VGSaPdlj
GhE3FmoL4q3WAijWFtwaga8ZKUTNsJ88jZUrrRbiFnks2JHPG6/Gnr4WCIVRKWaU
Im+OeivKrLIcL8YAdWjwwUIwTd0qA2qfEfCPkyIx1DuyGqk3bArhrdkXPPR1Xsn0
Xd1Xn5p+xjXH7uWcsm1ydcOSdED8Rlzzg6f//bG7RO+GHh/PIWNe11eh+iZ/Nq3Y
6d/iFCrCgGBCyyZDOoRJrNqgv3Rpu/EJvVEtXb1Vzmc0lh8DCNZ8J3AvYGx65pDj
Gzn1Z2piyU2/q3e0YxZSD8UACpLFEWNSvUnr7j2icbmOxp4WjT3Z0brx/TwHafON
bFpgFTiFeVKdVqDP/wN8OSs4RNfne7Z5oZp27v/F+GAQ27JdTZ/LFXhU+1MZRacu
y4p0OVsIcKZL7UCK63iyXGXyTJPJLFanUGSVZKNKDixghACjJJ4w31cF04pyGIBj
Ozd5RDwZH75+4KlIwwhPsa8BpyNqwnbqLmmdak6Z5OxvEn+mlO92ZJGDrNMpkUAv
PCZxzI7aSQh4jUUNjyFh5061I/Z2Iw0R8IOp61YX63f0bzOXnATLCgoy370COp4k
8yURiAdQDHwrysDXwq9qUHOEywb8n48WWhXKqznkrF592IMvUsqh3XXbzP++2N5v
Bi6eiJmAJz9L8M4cqfJ5LKJH683aisH1AdjFqFAizPt5EXz3pM1FnK2wuaSZ6Jmv
gDy0KlK5dPyHDF/OIZpCPZgfWNcF7gFODJTOiOqKcMntR7p9aUflx/iLWOkrPew+
Dp4TqZ4bPsXuDdBcehzj5fhltCv3/l3kmI1gMCFOThAZQDOdBNf52rVYRiwBnMwU
nAQwd9zDiPqjdGBGrMU/zkpcr18/3sYa9nucrzlMQVXyuMsmG+13cKUpEVez/tjs
wj9cx1V2MY7ng1ZDpqw/KK0snd3tiUygR+nX7r2HcKb9I8Yh72NdkMmP7vnGgZ3o
GRmP5DPr80b/JRQ6STxWV6Rnxnr63f1ZJp8Qyq58dSMYzxVmBmU0qyg0gkkq6cVk
eAuXEfLnTKV0+SRByXzDUcUkn9hyju2lZk3hFvGDBqG61bUbTHZy61it7y7wGNGr
sdqexrINqUP8bmIutWKMDGARDJQU/QbZngb9l6ZY0l8U3lughlRHHHgqiUjvmo04
PPz882+oh/A/mueorETM/CcS45+/+pQZ7jDvUk6Irw2Y95V7+Rggs/TNOmQb/oX4
BrxU2ULPF+s+PG3VUbJrpOIrG01k5M1hasXjeJjtrTWWwIrdvPX88oNzk1zXVSke
LvnBHBej6VoLuQRiDbtXFKNXxss6Hte1RgPBNGTHprwUbysqHc1+6uLwKXtmN0Gw
ufZB46fFkqldkIuRqXxV1NGlzM2TAwXj0Z1woLGOpIlvSvk3k/AFZgD0bVVqWmmj
tsVDh6TaM6pxDXFdlEzl/VTEnlph1YurPnwuSr8pN5/eJDcVadInzTwL4H8kdlbk
rnxGrw/4mswKkRAazdpSjKkFziU5TaTv89FXhmP3upc8RqnudaZ8ZeMGsm7z5BY7
HG5Ndbj27RsatmBL9nNo+vlARJTEEJaAubDF/SQ7ZdkvvB9pvD0q1s5DseVYLRtT
n1K/OALdd+Qx83gYMami2icC8AdGZDXsoEZaRnzBRU/kHO8TX0YzAjMufxGoKoi/
ywq8YEiwyuU4w10HpQMgarCDIJs1ksGS19KS9NkCqEBrb7aaz/4H0bK04gC1CESF
SN02yWZLgUhzNhkNw7Uta5lYrNoZOdM7+LFIjevny9LJ+EFBbAeV5fjXRlOgyf8t
jI+ByDvTyz4WkOjNsnkKiUASTccjHvB8O9q9WlBRiRY0pPBj8/ZRlcYMdhl/VII5
bR1++BxkLE3LGLadUPLzXlAToxHORUhrDatZjg3nQA0knVkyd4K0l5Zriur/h0/g
mNhlqrsU03hUtz0+Q5z8zCxWiQ+9MJ/N8HrzouMSYF5YZbliAFgsMbZNR6ylFKFD
PyXO6o/EctJCizQl9sHBR1DQLFjf/XTV6KXGUcGXtZ1JI9RtpJe511SLORq4G+YY
LA7C4It3yGqqeWwGhlK3FOh65IcRLMdNbcRk9QI1R+GeDgqFObJszXO/xzb2Cy8e
JXxBrh2Y3afnkTOOuFqr8R7ERW6v0MD0N6LCyi6Lwoz353JlYMAsWIHhKXjQ0QVq
3TivizQM0vmSvAaE2qy+8oOuO2P4huSPD2iArmyrr0HIPwJ1MxS4xAIz+HGLX0gU
cTh46wbcwmopiEWKr7XvAkjhUoeTfJ0l5THyypVt1fMLzM7hpyIkgRkd2XOsz/fS
jCQ0r0bgsASp3TMp8OLKUb6m4uVCL8+sNQvoh2sqDp7GGnH9wSxpAl8VijD6aWFV
YOQyWeuqE2QJFEjUYlkfBBvy2peK2QmcW+4rmHl+V+2BNtBbx/WitDjyDQDPTDHH
aCpu+FyUyuls0NbVG6Qb+jO7rbZPmPsVae78YboDhuJY3glSiqgioW1hEaABc2A4
N642XNteep4xFYEcwS3xF5S0rUxXLCG8jIbmt3zaxq3xCvF2k/AB+OV7nJ/OUb6a
ZFqEGyeTHg7wHaeGeJSfJW9UTMPoXofIo+emAwJ2DHMylx4OYwdN9BQ7oM/10C7z
0blOcVXGzPl1zEHhJ3ezFzS6O7mgkG0OxuyUklaW7E9xxyWkxddvyu9ZeG9L117/
OmHhhq9cGeUvmEaLx/PExPA0MT/YasaMgyY26Fqc+LEyqBrAkpcHX2kHhK8qPrmR
ES0siMKGjrsJvMLToSWetZYe0Z+M1cR2jh20LrPcSFL0OeHuMY7C1XCfDTcbb4se
4qCeyvaTPalGGUDp1hAQf+HtnqHirLoY+VtTAqR96+zU1+KWIVKTOehIw9EEqmGU
QOs2H3REVDLUCRPmSWGkov7p+40QJdYs3cv2CYyI5QYyU6Ppq6v9i3nYG006l/2Q
HHbf5VaLBF0l0GuPdGxwcrV2HhQLfPKF3LsAOq93A7P87kYp5if2lzHIP5e+2ODE
D1YS3XguYX3iN4/1Vmvjxb0hohMRAs03Yax1meDgLBfxXWGDd72kUxHulHgX8EIV
UDjAQE/eb+9vYMZS3gKVuCiNjhFzuYnXkOpZeQUtX90+dvYGb8egVVCVlJjt5OLP
QCLHTHfKQ1iA0Ie0CBy3/leVPW+93I+1FiyBFyIniS1A8gTfIknr+Ctybz4esyyp
6Z9R5JuisN7dyyUbjDKYms7Kz4dqEcctWsR31TXqnuEgYee5fyGHpr9Efw1WrTtA
gBBFd5SDqWIBLP6eCE5J3R9qpFXG3vQui2HRo5sD+Sj0CKVOOhRsVWYmFM0CIxSv
d6kJkmif745kriGc/XlIhFJ6zzGKmFutUJk8aj1bLQGDUa9PiFgmJUad/CQ8NK1G
B0IG/dnr0bkZsboNDXNrw2Hm0uDC8URo068jRVBP/zkxLOM/ZoXfiMMAEwwdy7bw
4Mjr9BxChYVrG+K8p6Mw4ACh2mq4hBnwWdVDG3XSwwyaijeu3UncRw/skG4mJehT
qNgsdTGyevBq8zKFmywHOnskXJvh5DpRLeXrb76xuqEcsTUGcEHJhw64DW1h+pr5
8YrFKgeS3ntGMU3qVsJNyIIGJLa+l4hzkjRmSBMttogCTLeJ3XGl3LJZdeHWjdOD
9kav6IYM2jTkX2ea684/e8V5yP5AA6Kt+17hYRnHtX/engU3w8ySmwPOkd6veSo5
oj+Dn8S3/TQcVR11YLaD06Ym3HskM+shKaD6I7fS1twCk+UixC+lyZmHUXkLUC9E
wYuQZqSqzeqimQ0mM5Fr4U0LKKeB3Bj/1LqAlaklY2BAnJB7faDb8r9+tcUVHJ8M
CQsMMVfXwn/+/DyXTa414W241W4bxTZRolAeT3S7TLIe9ZPxNskn45Dg5txgpCzW
VQ/sFSWXwbc+JMuTgXzdSzDStJyv7H9U1G69mnIkcO55xlFlwP4A/ZSFCGVtMCT6
jXfEb7r8EkVjMv1Le9ZcdFUuTxxyfJAGSB/4Mq27LsEr3GPJ31ay3ZHR8sJuPQJX
67cRrPVC+r3SlMS3KOssfniGHvylAnhawtyPFxhryJ2vDoaDFPh4sYkpuR+y93cJ
7T32PbtGYezr/CcNvFf9R/pOWA9dKccCdxNh9tPSbKasuYwtkD2WYUPjvBMCk1Yl
DfOZYuIL1f66RmpDuEVmPz5redm19v73/VGrghIAmrXmjXpVvd6yIRURygqtfGL+
dqH1B/8bt3pyBFPBardu3jK3YOP3TToHYtQNETMwNK5o9cOj25Dbnb2qzGd+ov3J
ANDaV+3p/cPen87mimOuQBPYH55vURw0yt2REgswA35MhuGnRx35IVjASGuLKphc
J0+nay1Aj9JBkEHvf9Kb0wXKlt79ikKhCNbqPq4t7MOKoxhTa7qPZjMKHMsRmgKB
ONjuOoQ/I2aFZu36/vDYFAb4O8lN80xIufkHfIIi4DG30lFkQlk32QAVt209MwR0
r694DcFKtRR/7Bx3uheB3j1dzSKIyjKGkD6sf74Gh7IC4+tll0PJREBGCow88kMN
GfcXyk4JpBcILvMJdoEyaXwAY61S57YODwiu2DfyFqprpe1Cpif/fC1RR/dX2gDX
2OiB+wFQ61vFMajooH72bx+act+E20xoi9G2hrrMia9BzqiEMMbgFAnJ1ORjUBvL
qYXrO9rwJBYP2JT7c0AABeSK0//ARWHPBpp+gTVF6LRFRcbIoMysg6OED1uPDL85
TlwlKlbuPP+FjUeXQIr6GZ/xiPqa0Yue28YFyVhsmtrRD3Ax4PJcrS9CoMXfmSZJ
T5ecPegSpzKhyVcZIVXpUnqrCEoTysGNvWYPvGRQiSpaQIhrZ37QmT/6/cRKE0pa
uUEDrFs2/iJ2nTHbrNoTZYEEaLoZIUusYJwKlEV2Ura4KLJ5H8frvyBa94lSOWB+
X4e+q2/mOyHWLMK5Hu5WzDTC1Uc+0+9Ly2UOfEd+xUjRh8Mzk+SlA+V8OLyU3IWq
w4UnQp/2Qh6QYza3bpO1gANDfgI7ayYEuF/yczi4YgQQ/wF9loiNdmEgHqhCtII2
iSVgl8J8lIpoVmjZJLDzyaRhEpoArDR/55UeNm0NF8wekMBXtbu+FeU9Oc463lMY
OqzXd3OoFduKytWT4G6x7D8hzb/1lY/RXhQfRDIQhb3R6hpj/2UKqOCHpbuepItN
fwB3d0F3QUlXW9KWBQVl4w8a9s2iq1aEtwLJSCkXPUGPEruzL5Uw3QupDbeWPLf7
M+rFIwo0qgIhRzVYlrwV0v/BEW2iWpFEahOO7ATIf5W2RMWN6Q/1376ZDKKoLtMs
nLT70YijL96x4Pug+33b4PnPAhzUOvvEE//PfHM2M/nauD0DLGB7sYH+KRSR7p+v
XEeEaD2sPLdA9E+OamRnd0ye3Hb9wDlPV5wWr7P7w4qQ9DNk+lkRnNYWD7aFsLOt
fjam3f0fjzjGZDefgCPymDvidgpu4sTXQVrqACbDjrEIuRBpTc5ojN3zpuspmR4P
UdfB0fXcKFKbSQW5++TCz7BDc/2RU2lHlAgXmJWRdrjCoV0MUnIDPVCLq5u20y4Z
1iTTC8Az/t9/4jT7KdqIj9VTp9Mv8y67bPOf5lrWff+WiFJAxj0cUpIdbNFbKglw
9P5J1PkfALqXNQl3nupfJJdflkQg+s07n2PPIEr32XGqP0BSKRvjuDphlofLBgmY
PWwgxwvvJMS2z9EWtHQtGONPrk506/HrJ/EC+GWL5PrxoKiqB4C5JZpUr3BYkqy1
TZnHBznltiYhaFDgA9DEviiygGgM40o54OSy1bz8NyLkLcXiRKjOGkCgKvwa2LMK
Di3UGnzIdc6JAP2PREXvvc08m1eYhS5PqZKRdXVPzOjjSmu3XE6pIrvvFMeeAoqS
1IK4sHt+C7568+0cBiCcp202W7MzVKHNxWsMxAxk3jXI7fQezJ7VnCapzB1pjw2+
qymq0t4HSwyRhnY+YRRSKTtChGO5FsrZTeNqKFbV51W0KtvcM24tv4w9aBcbepVC
p0a4YBqekYSmA2M+jczP9Rmnov+VvTS1dVcJOBJgPkIStsPT3bCXVHPoZqW7UZ5T
Py82mdXTcY/e2WefppqaCOmQ6se1MQEKL4xuWpHZ8qOPGG1ip9wKPsllAWJgPrcy
f0QpEm3wpiEkZFKhuWhYrCdtE8vZwdp7G0AxSuX4MtNtCh/gGE76jsijivFtmX7f
b0SBLYe+0p20X0V1lm+F2qQQcDPblbNoH1NUM7ik5hloA9+qElFWqGMuUnzH9sVn
tqfSeZRTRBa8rJTxPJ6y821r01/35Ym3v63KqdlcHZbjxTw0bmriDcZrAUX+IoQG
FrCd5M5wyflTtjfCM1RnAu/92CyUdj8AobYZPhOe6thn0CciPuQIv52QFSuF4jSd
7qlyI4bQcdybNoGFEj2BvX9jmJQMn41TURDt0RSpbQKQsqaLSV5y7jv4FN0ehpjj
1DHHVYKxsN8BV7iQ8cuhIDeCGO3tUqn4elF21HISSYgMn5QoIlLLxcwpygbnONd+
IBlDwMkIgP2lNZOf29B5muEL1/+amwCX2W45h/ljdAkiW2/PlHN23O+mY4x8QHZH
/yxortx3fBt9jKtkUUJybggkfVbit4r8ZNJinPI5BgSERZHitoCzTf3BP87RMSq1
I+aGMVHp36t4kvPsJlmWsJDtIMMzL8IoloFQFDB3Mfm0+fCHpJOK/SeLQbNMRtWw
ITCOREV6y7puwgSKacuE/yHyxvAn+Onregye5hsAz2L5wp04eDfceS6z8IPoH7GU
uv4GGbqh7rWVbG73kNaHZe3F58xd2BG1cj+CjSCHzFyCNcMPHbLMLlm6swkgsS41
0fFptNHg/HQ9v0YMtZUl7eliZPHTnZ0w3uJNrBhP9rBJODoGE+WFm6Y+37NKYMsv
Jiu+YFxdBPsDo9qY7KlbQoxZf5EL/yZreRJLLbXaYG+TBCaxLttOfo2Rg7jjW6/J
3YUzUZTuMICgG7GRegIBwAJRHZYwkTIL53CuccazoArzdCnO/sogEk3vWf9jwBhJ
2imjGIQfscdOlnxGlHxExw01vF1GuupDKzT8m/HmxXzjfFt047jMB6aSsL15+56+
mgMIhENdfeHU3A+ylKsIA3Ahpg8CZj3l1GJKEp47ut9co8B32thN/98oDgQyPZv6
+gsJF/ylGEBmg32guidZ+xjsKr+vEHyNkBn5gttxgu3Huj4e/pFEAYAfNxfjbmm7
ERG9L4C/QQkm4gceBGBfWwMPt2ykow7a+MvUD6c8VGKk9PDZArVd7C170PH0+vKT
4xYlNNTcUsAcmzVrqdOHTPEbKGiNHx2giWOdasVGKpzdldKKJMFT8TpFYXEJ4yum
s+z8OK/40F5XojGoQwQZtW11gi1ToYfcYCyn01iiJqXViltKAPWSGT3FYT2Ic9bG
J63GdfvXdrgZMkK6kFeRJZqaT2rvalPanHNQwpdB2v+80/tjqJYY7CRJGfCHNCCg
rnrO7305GpyTt9Nxe/3ELcAZ4Zhby9kUUDmAP6hdxvEi/xABhDNxf3ZdbQI6rfcX
9BxtQSkMdeJYNqE12jB5NE0EkciIGTMBlhzVCpwYcE4vEYkVeChUBqeneOfQlvFx
s6KLUz6+WMK0Yqw1h+q1g+KsQO9QQAgHiov9szeXLge8EQkfyEHA73thdUDrYV9X
JLd87HJ8G9yKPbMgSwmHrsJP4w+tiprG95X34IiqjMD/Xncl2qdbtxi+DjoFl6E0
tQsToRe7PlpaL8M257ma4iZxJxZGDRYxlvdRhGE+7ofv4gYy3WLXVT9/2EZ0qrYa
/c40hPYVW7m8WFH1ESnLzRG1GkiX0rum5O9RTfjv/cQwubHwkpnygEhfFUi+UbKN
yKNuZmEJI1mugkSPIzgAEE2fZMgnTX4evYD4YAn/vXoK9KANKk9jVutfVkjDTV8S
crCvGEuPBjfLa6xQm++Qf+NjAQudYchQhgHNhKbCxxdaSQfCrKNoMrXcFLjQirsd
R9xq2ydLbS5y9KwkI32Mr0HPPDxsUHgIbkwnQTx6Pn2G57Oq5bY3ouLvdny61U53
+NX1MWL7OYjfOcq4xRSdFKbqOaL6l0C1h1NJbm3/FDtVkJZqSNUL7mQ2veyir66+
QZNea7rvNqx0BoVEjaiOUNC/D4IZS/ff6yZvy206ImK1Qjk+DAikKjwfeSTkXZt+
JbOUSo0MrfmySWitthM0CDHThMOXDLDQnxNjkgHr3I48sLC5B1CJZ9mWD/se6Zh+
+5ZdUcx8cB88bpsf4lO6XNz6dVxL/PqI4ibgT/XogkPkijKi+x4mEZ+hsaDFpw5m
aXMzqAnvuRKK0FgkHjQUersa5cloQFIb4f6QcyK3bW4QoyxPnI1rn4l8fmgL2Ofe
9GLIHhfrQLYKNW1UOe99p3vMImyPwnfteF/03qtkS7HxvYTCgkXGH867mb9wGPZ0
dYTrJ/Km7KAYbHpAjUdBuQ==

`pragma protect end_protected
