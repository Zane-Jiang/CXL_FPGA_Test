`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Ye5ndng2tjfEh0z15GTa7e4oAlvu3UYhIPZZztLnxhlhJYtdXGF4pUOBCAwjpV0R
aU1hn9Qn82mTx+qUeqvGm4Ji8SojpwvNxrJxayvNwJT/VC2+owQU20WeX7YBY2wK
l/Ee6hQoarbJruTEwQWzR3PgAY1JS0llJ7NP7vgtkR8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8736), data_block
vGFi3uVlAPdROKU4m42d5dwhn/CkUSL5fGmxnDu8Qc3ivwO3zSWgaHZeqLDHD+bj
gNhH/qd/BIyhSAanGzlJUFGJ5wcOI92Ig6EG+FUxgOrGgKXi7OKaQpMk9L6Rcv3b
qVILhaTfwk1FP7O5TQlKa7ZH5gPsm9ugwNiWW/+dGQVSe0zYw8BP+Z9XM6gCn5S5
nTJRxpchnq7j3cf1GSa5HK7i5cCfpthOw4JVTRxE2tt9sneN0q5HsDv0K8KacgCG
CXaAaOsFW2cGpI6vPb+BBhp76csDQvtV1yTfTJJPrK3N4ff8ihviZ2370w37j4ND
Nc1092ysg5qr5sKra5Rp2f9wwCphHXZ7gJohbvin8WXZaHJreGNdZ0OrJDYKezPY
jY17qQN5f7h0AvZqgXF1o+GKOj1KVPkoJANRlDUDt5b0FQiGUpzzuG+7c65Hh2Xn
RQrHAVEzLnsdmdkz2vDWZoXhZdu/MW8B+jpuPCAzP2h4P3f9m9+wxR0v2nCHCFJr
6T3V6Urp7P/G/5eUNpaHJz45wRpQ/HU+OZm/7iCQEyElQ9KxdT4lgjyzTe4bJrh3
mQcvAVw1ERlqFYzTcAFm6zcn8qLv74FlM8pFaf1jmSEOyGGAEm9oNTnPadYk8l9Q
cdgSH3SyuRsRwnUjRgwnfNOdn5120ZZBztaV27lEy30yVehbeOSXBU0a4FvEjVE3
bpVO6fMUsVEm7Db2Cvioob5OrZ2CBEjVbqEI6BnSVWoDCjPfrkI7sISyIfa03rl2
JF0g2bmHCUxNpSMTKABJlMWomvRAsywUt50nAatLRkPOu1feJG86SxpoB1woCDjh
ZPuKrhEekSn6ZCBYzrq5HfZW2w6U8NLfMV6kS97e222gQ74SACWGT05KRZLhqYLz
BJeAbkWM0CXtk2qrIKrupEOBf/iLLdQwQM7EcdvP1yBBMJxsUsQubbc0Hu4iIVJJ
I5AUAfS2RJdFjkqTFR2d1vQ9Yn2cM7mW8uqSBxSnXbGIKkfYGLLVbaKY1aterPWf
0FuiXVgM3qTFGXuvRqxt2p3tEa+Qhtd9+GtEsryk+JYC8Jdq93lv4wjhCDr46pca
mqwYxA/REy4y8jBpS38R6hwj+QzJDliVOWlk9vK/+C/0+7W0biTKZG4ydVxtAnir
JqWdjIpB/GL/22X/jMqp+YBL3UxEpWLuOxhraALMWCHWssG2f928zRMyNRQ7+TB3
HWDDb2guSQv6n5gfSvadWqHtc59Og/mKgGvP/ZdGnjoxXrgHaMQmmPERTJABPoVm
OC5fILzUrhrujNdt/fU7WhmkEl6IydE3ZDW1lNHNiPWxz2+Vk3a7bTe6IH8I/Vlx
AB0IhFUk0OYulGrBCE8szVp4eRyqTwjGdpmQ4Mbi1DsTqkr9COyFg4rIMEhfow0I
clH7tgIa5uYNUVZq79YfL4qpacd49I1fmyp5ZZfwW+EA3g3XMAoCRCpUqtUkHlk5
UtKx1nSf7abiQub5wGBfuBPBBPAbQPuabYSxAPTEkey5ArHLPYOD1w0bznao/8ZK
OEfeXrLG/J+h/1Pfxu7x+ZxXunFhLm1kiwwJBiYkcq9ZFpjA6pWYb/NzmvzdHOob
4bqwRdb1OBnieUXPfB7xEp4v5EAqanUEAbfSEn5aCiNnT9ZygiYk1wxfGEPznQvy
7rCEnCQr/p/gxo8BxZFd8bsJhz0afReVQ7QD8OqoSuW7o8EeoCYMO091xRwIOLvm
jH7JTuOJhtaoKDgRohU2a83PsUHggu2fpRlRyFJN09Dg8o4Du7uLBzwt0L7B8DMX
BpvQcX4EqY/AjQQ+wwgl73zWoVSDYZUlh++mgRvWiIGmgoYiEsHwtZyK21nrmbMW
/cznTPze5uQ1qOk86uyKMFBLXrzT/pu5x+U//r+iN5oTEqq0JlNGwmbETYbCMj5p
tLslqc2khpG81nvdQpnXPq1RCqPd+FAaBNA0Z8M1dVDrlW3x5EbAiiY+YrVDa7XQ
+paR9Keg5veeJ9RIdJWAjKnZyL6VC+DFFsr6x7TxVM2CudXZNCMRKMGbgzTxvRt0
Izrgneplt1Bghzrq2hnGNqnPzPN9iYnSTaKbHdSiarXs4h21CLoGhVokfcHPLLJs
iw5WW2iKtkpxwbGHiLIbJWhkb1JvlLgBaMl93ELo4i2sW+5v/LAH9P9V083IJZ0Z
FO+DaePTvQebapSJWtjygtL46yvTgaSzhtQjZr3LcPlTCQP+Pka81Zi0M8h/OY3+
3IMUFnGwsjvGg+W1ymP5GDsbRRaVfLqEhXrhG7IDoAkZiByJwuE8HfOAGL4KZdyq
pWiZ+zu7q+8gsKmxBb243qQ+z6MqGunVadHlgrl6bMTfKE1uMK6qvsQeHcJ230ED
H2up+4SIlHDXE/nZCA9KTfY8pNPA2Uq7OcdLcFpSD9QtZED0in97XG440DtfbAmY
ITNX0QT0452d0e6fMErgYvPMaCUt6JzKvV+QUet1b5al5rj1hIRt79LSwVIbg2gN
tjWYlB7iiAfTxgeAJH1/oSdSGbr8q7p3KWeu/vczfsa3P880PFWkxQ1ZUpoozYFR
WgNzyOGzOJsCBrZwNgYvi7HPLC4OmRjNupjHTZv8jrdkGNnuY/yr4CToyLLoPN1A
wAcsDjVmE13eSlNeP1pZVBTHWJtxXQKGJzRvSly99/46kOHlYqcbBpUXwXBXh3PX
kpa9mnv+rRlOVIGFkaB1vkgk/xQY5Ng8A0IlT07R002u+yeGWnqR35kugRkA4ti8
l8kqLcu6dzIUXb5RASErJGtrQtEZKu7yCvzUHnZ+bPZ4eUyALnJhxFN+IRr0HUew
lBt79RS1UZ4Qo6ID9t2z2hA8fWPy12Q9UMlrdFMNdmVjiD0daPSjeD+SCZdofwA4
NVcqjjyzdFcZ/4Oc9YtXX8wXsmTuOxmLCmPOa33rj0SljjY4Y9w/a2Q4HKR2X5TN
5k4yx4mRiA/gGDlFCiLTCboWnbOx2P0WI2g/Qz23EBLQfTqsMkXS2S4sEoJGiN2x
4hfSxgGoJoFAeR6GEGRNARHaZOa1h2G/8Hj8t0Zm6XRsxjhB20LAC4m0AoL+BwyB
oHwJtl7m0WWoZbxpOPGDPnhW6aA/vGL+6GNDXlnhxDLgDPYO/UqHHPqxd30/AId6
FbRsN26dbzZajnYISRat2UNAEmfTp72tmCIQs8BXlwdtxZ2o41pXnKBWcB0xg9ER
RWINXvtWVPBW8NinTmHRMjeAGL5h6mqgpA2QwYiOdMJbjg+v5mQcR2hjrCSXZ1JA
XwX+lkcySbuyVLBso7vS6U21BogbfeII3L7LR1ckHvl/Pm/mocGuoW82KKK+6fPX
vk9myI4A2zZgkpRna5rWfcKc6OC6bgq4M+ufF7d6u/8f4MoDovMr2UBO8pR6N15P
nvzjYi4rRxGqLJ/rvL94cyY2q7vJFe1LrS7WN2VRMsZ7z1QKe9c/hwIGQFWM/6dg
Pum88pB8tkZ5ATczQtKi/Fx88TCtjmz132InR1vtWdDe6tgfX5Q4m8iF2rGBD7qi
UIFxZcrLJTHfCz0omIern3q3cIVDyj8MlnjmvnjHlPXHoXxqaO73EFDbHdpzzDbm
tyvoQXbUGQ9J7Zunh9SkhKkvYRCpikwJAPkjgage/seIFk3mp4akJvDlnfFjAimy
MryoTQIsMmZNMqkZHdXQvFkecPi1PO4uQxEANPDwwFbOpf9Kic6MK4s8iD+I5EVL
2BFJ7Bem1kjDbzYTUcBWOb3KEPwv4SpydgLcMCfmQvhTNBpQ6Khh1xhLCLY6E24s
PHyjG7d6HoS79meWTticBr2Zj93yfeouLwcLKRyAR+S8Jrbz+rORiVCdneEjpsLu
L7FOkUyS0Qxn+3GQkpCf4vZKXR6nqM6VDnqhxfUM+Rw6D4hoDd1xHPQdAXsPPOV1
nRpTgswz/EsvZ6n8/yLpTd1ltDdybM6dYlNbDZWZlVt2/QfTaq1L26fVYZJ2PpG5
xgziVCtFA7NvL+TfjIp5ygcvnAwllIeSajtz21GuI8LbgsOiWT24m5VhEoXab14F
uI4Jz5HZ5SkKzBLxzJgpLTMucOY159fj4BZXwcO2BShcrh+zbCuefoUiTTRgMyjA
RlFuZkhJ6Pbld6tQl4alQtmvqZPM0/DWQm1iMeKDb8xDeEoFCzfVLm+s6pj1b5aS
q0BerzsFt1hdxyvm6FnVzZo2Bzh6XSfSvScYVUNbQ+QH+Xr34pWKjHITEjwcSVl/
NHWf27yrkw0nnua6P/6PzYXFOSSUrbCi8Oxjsr9exmNwfHEHtQd9lb6t93lK9hbK
D0LA5gPI/+32j0HYofrY7psifLVG5htQcEEjf9Hh/vBnOC3lEusxJ6MnhRjp5RpR
ATc036NtnYky3uFf3cHsoiHZJlzVgPo9EjhzTNgvQiBagvzm/ATxMCc9uAiqf+T9
Z38+Z73feNZ/jlQZehUzYul99ZHTDG1fDoCT8CQ8NPnlpper0p0m/YVyZXLLEv8Y
Wmo8eCoomV+ApupyzKdp1jgw362NEMgLiBt5I2gKZ3CpbRuvYjwLEmSx2YMKA9wj
CS5K9TJeueeGdFCDGAu9mvzKInCbYcwVAvxjmm/jG1/rISt14SSEMXnCGeggA972
2bscRbeLee6IQ30JKfGPF9RatTAVlGLTXwJs6OxVSoVTYenZ9K0VIp67Yk3InTNB
8RrOu6uWiGQkL+SigiFb9zbXVYNOsxc+qzLA4SOXIgNMOy19b/3RqlrM07FqqJxS
YMgipIL8PZFhAq9OD2mIM+/pSFOJ94umEYHP5Hdb5NsDoXT75C2EMJ4WBaDCG6Nz
2W6LbUM9xyDuoX+s0PXXOffIPgoyZmLwMWzhXno372K5NaPQJafyJO7iWyYrG5zR
s1Kg2KDgYVkJSMnkEatcJuDgR8U3KFKynvaFypv75cubUKhxJawN2P9burGDkFOo
234h2/8cI0oUbY7iQ80WaAH/BsK1NDU/1mVM86Nxpi6o+eFNQDPumNHQQiIfv0LK
Qivsy6VcvHPvG8JkKZ8SUkb3tyXoaQU1zzQSYhlG7LLuSAv6OP6JgVY3E6kWUpZA
sqx8wUuZDcWxWYwCyNESbQF8rSp5M+zztBLRfMHJEod+uYqzDf0onU1toy9xlsX4
5Aymd/oeWRlXnHOv9VfQ33KKMwQXxmgcDW9YStpKtnnsEKHxLZ6CN/HOtdTzrhdc
jOJXQ66LDtjOmU2fPnAOKQnfn9XsbgR0Xo/btj6Ve+fTmAVZ5u5+NG1O0NFcNv0r
hXU6ggKJuofFbvAHJD5Xl04KuWheJLesZacvweRvxCx7cW3xRLSPXJjjdGaLzIvD
FbPgVTufmIPWo2LtU91pKjbaG5q5G9uyHrns4GgXhXboP11+eH71uscM0GE7S8/W
eLL1S44rY+ssRp81FjpdNgH8UfzU0xc5kPaZBVfZ7riYyZCqq0S8Zqbro6LQqqvn
bUYYT595HMiIwQPJr/pxIxW4NOHG8RIzFEbw/+sNgKs8UZNd5AUOVAAeweuAKDkm
fuHjbU7aQqXRd/SqoNI9f/TI87ewPsE4XqU2Vy86T+mdqbzhs3fw/BCl/vzothTD
7wLF6SSPS6cPUyXiCtFiSY2nU44OK7Yic/e0dr6JJNV8GFukoVbxa0SmCL66BD86
8TRI3QKcJjOeoyw6Tugiy4ayhaFPqJ365delCiXezOTR2aWu1LkZNZpUtlNtVDw0
xvAwiQgMOfED5EXuFZg9QJijl3mHuWb1lanmxjZh3155B56tJs0Juc34Ueu3bfka
c3inGuCfHegw9pYsy6iXhKKIAs4VWFlFBB5tpE02jDTXtyxQrfDTSwPgKLBlNg4w
ePUXNy+qFX+WcrZsvnTSv6Kc2cmVW6jKelRoOnNk1YkE30zPPv4/UwfEW7SfCef0
FlCCr+4MOEyw7niwN3Pw16pPF4oZfvuf/K0jNO+MhUAkJX2t2P3RuGmaUbdm2WOp
any62OHxT2PoqKd89oOxIT415bM1OawaX65YXkW8YFh4BBKGEYn3idYcsB9z1kIh
OKz9KYqjgIvEnIQCub14zRLjjm8dEdVBHGOMdNHtzHb+/67cdyin0iadpBZucXGF
A3MeCi5SgVFwXW7C5wsU2YDzWNv5LLM2oIHcEM8lRO/kYzqaQWqyrF2VapLK2SLK
AM9Z7+F4OcVHMMRjCtJ8poHNiMG7O/JUHFFcYvB28unxw7XTQjpQNWjVpa+0QFgD
H04ZI37CIfkx8SNi3vzt0W8MZk1oO1E+Eae80balTDv+6z35fK6OeORD//NLKTTl
jXyScnts8dy9RqiEsMpEdNTCivarqweCDl8s3owOB6k6N6yO9WaIbMODcnxMZWgB
geaLCf+wjV6yXMZvASWNyVXtRxhLWTn9aShLXwUM6xa7gw3gFLREQ9pBdhHsD42P
YZ+WPPjUq03rFOZDeVCEC0hu7l/G09RxmM8nIDuQbPRMkAmoaYStrKCfzTparXyD
/gHhdU3Y/nYzz+kBuIg4hXcIi009dNYidj6mZNj9uUEUnLqbx0ssdYKv9jzzLdKO
i3AT8rBAZVvkJI0ndjG5oX6aX7KvZy2dnRwL+DEc0lucY2UILrt7NDmdrCqV8pGq
o4pEx3zlk5kp2dXBqjF5769AfqP4B6ewpnv6Eq1NqX23j1CaJ/FFrYS6KQDCqqRY
QJuPFnMYD4kA63QhhNzhMflmeGPPUCx7ZtTVx9S6AzciEneDPq7tzub17xuhj6wJ
njnNtFHaCocd8SDSfCv2lXQlSTR5NIDlYMR1iCnxuL0Igb5e/r5jNBZCHIQif4y7
WUuQEg7fEW/QntUWMsZJe9vSLVKH5f/1IqMQaOjz/fhAFtSdg52u2gnfNxvy1I03
JaXcVvIsB6cZDahGuB85799WEFUCc2tbcQc8TF0gz+D+E9NX86cSlFEIo+Uys4kV
dOEHbX8m2gQOGPSR2tY1t4bL4bvXESJX8iAPgi7IpTbMpTYu8ecrT5JA07qNGXYV
b0oOEYC1J6clF7nvvMWM36jIH2ponkEJ/fBFr6vrucVVDZp/DhJgqnoVxG8JhCIY
p434ZL0GIfu3ePclb915nmO3yNCpRt8YnRbn6x/+c2fLwIowMiVgwbc4S5G8hGEP
2l+V6+d9JjhXdJx1ewoO6jUrpZVyO4Ys3sSASEq+64/fS08eZB9YSxwf+3hTTb/X
dChksDKfwz0hwN/qeJxZ2Bw2UiqMsiJcs0p16h/QfQy2GhxiQNIWl+lxSzezGBvU
+B8k2wYL+7dOhgUhaJgVCNxbpoOxxcwYeJt3kw4W1h6rEVYvnMIeIjPKEbT2ZxsZ
4+QyNr8SDd4prwhx1KAgrv1hkQOZ+JT7rfG8Ujei3uakLn4rVLKguJknMCoxEtNx
I5V+zT3nWsluak3oLy3a7A8oN5xesaJ2ffNdoeIzT8Onr5QZD2nhKYgnxazvSRgp
nGk3qweSvT9wOHvkVrb2Hxu8kAGRA9XZhNSeq6wzVWKnfazqaeRT0IZfrMTJWS88
wRPn8MesVIwL4C9vcNjTlsawfCLYXQei1mLcfYcIKIxGBuBuT+tKrXvVp+bPnOfP
SXZatwEU6JBgjpapal/fx5W1oabqEDxz95QVuwphv242rK6W0iVuXO0qI3mchd58
JlWAccQixh/zvRjjQdzekUHUlTFZEy9ypRjsE9nAze5/75t2DCrhpDpJoeSq6P2M
l7j7AUHtfY7asOpXIK6BPaKwdVctOBM6fylm+NyuI9BpGGZn9WP2UQ5XU/pA1dI/
uH/cjnq9NYeZVdknflnyUgI1zsMS7RWEoqI8FMJf7f1Hr7j4ICi0pauyLVb1MAxZ
WrDho/v834XitFdLGo8xWe66NWYymHtFWtsWN7m4hoJQgbLXYYA3jZTEWgIFnFeL
IY3KtBYJKIRK1mrGGogxFQdINgl3L66H0S5BSIOz8sSXQE97WZg8ekgoHjTVRHBm
0nxNglfYDQvayBFnxO9vl7WBszbBwqecTebt9JMxooEawPzjb4knMEtfzHe2aWn4
nC5zRwplBBEbwu2WgqdCRhu5Cw7Ng3G65WZRFlObm+OAVH/j8c4V86uqws41+Qz7
pd2v+XK5Vf3TO4j+gGQZseQE0X9mkRRPTE7a7I338fHTlZqrzbHeLI9JhQGd9Pnz
u4ZhyMwYyaqYWHCTq6Rg+BOMj0f+xo7dch/EEcGdxFteaApHIv+3iJd9o7Otl612
9IrjmHW7xUqg6hIzwwy/gQSURXJYtMsVwWDSm/KLHaOhALw0Ah3K+WGCMnfJ4i6l
7iq+wG7XSdUNn+XTCKrWdGFpQ6YZoSqHUX0Q3e2ZvFHyngsGlrPU/W3wA28cXR6L
pwGolGyYnyTI54EsowM9zdvhjlotwQHqxGny0K2n779j23Wb/qoPYDpzVi99Zx45
Vm44Bdilr48xsKKcCP9+eFAaF4+cEZcRtyppfAHONxS/J0Yvdj3/O/qkNmsMFX0A
8bgdyAnad1f5tUidFMqyglV6zi/MjFOZxIg2IMrsFqQS+AJYGalRyt0XH+VL3cKP
g0sShkvwpOWzKwzBW8WXkxA67O9RNS7ZLoEHaW9hYlYmEcYghobvrW1IvjS7Y5Ig
BBouHLzkQRTUAoQo04hi+eJYnEyN+bLkLTpo7MvvOoP8tqk4+avJBiCG7mpI8XVx
UQ5ZHAqVkTOSca1SsyNIlqeh5/sw4ptyHucwEMLpDZPZR9lJmMyy4FABnAU/ld7y
UoqJJnHSHLeLPFrenCqgTFiKfPErB8TruM+CCaVcYifVKseBZusBL4zo1qvAktEd
H5/wBPCq/5fjhSP4IVPR2TnCasby568dSUhW4/R8/D/1ZO9fsLX8oj+14hPVLQAp
048PbBDKCNoSuWYi0bV3/pWV/bfoBVST5EY6xDZztGWNGwM1UTy732yHOfGAIRbG
Cd67ADV1ZpkYSdbxbdfhpFMwwcPKyNkjyKZj5lf4vZy6aVrpzHC9x56USFpKqqR6
ubGb5HjlQX5sw5iyXSxPi1ejst5ZAUretdUHjed3eY6H8ZDWBXQzbBEszDJXQsM3
GqvP73K8GghxEGygcFqHsfDNrv5R3VmuRJbgms7MaD3zf7XNyCGtKikO+57mSiJU
xVRcGLPyxshwbxSuGX3qB9kj8JVqTMZDhG6lj8Ri9xi2lEZP9hoFKcl2S48hMcY+
/QAtGSXtG3xFX6Yfffu3Bt/TFIHXod6eBpUSONSlTueD+DzsZDffP1Va8MWO4Qu9
S0HMI9u4MtzO8Xq5iteq4v9czCa3B2JaJanNVOd5aKMBoNBuWULrTX1aJMwyIVdI
vEvCBapbzmfqlmAz/ydJfgwVWpoQI83grkyd7p8bJn6pWfkQ7aS3M1Txuv/arbiI
aa2NM2r6NvKuavGcuPaurOP8dzpQqQci0gajwwldLWOOc9ZmQvm+qMpzqYZw2MlW
s6FzGIkypmZvHtAtLdDwk7+oJnWvwFKWygW5zZkwSzjWdwVm6xDaaWQ0cwHF4A4y
egae1Nw6OKN+THlXHPVEci4StuRVRM7c6N8ltdQMyiNkLjOxrfV81MXfzGWLohRr
6X96UrX0QaPS/UPYCyeYXnzKshz7aQ06ywV2ptXgJIfg9r3xUo74L2WSNtzIjIHI
R56h3yyBxsyj1jJFz5Mab2ilzPQQYaDc9fhrxAz7P8+dPswc7Cvzf45yOfVizZzq
VwLk7EV6FbVLHlauQYWbhbAK5rRheQkW/g7SGP/4sQaTHVYram5h3WjH7ZE2o2sD
Q9mMRO6PPOHU4Ahz8tpG3IO7UOX+ybTwp4KbslCbHMfM2XySbAT5T6f5Ohze7GQY
NIBewiknB3Tb2vcwwQHZHhjaKXcl+bqgfct0mdysTjOBqY4i70wfnpP7Cah42wdw
dWeMNZkdsBtgQDRpgxr5TUjbWL+meOVnCRloeZ2PPsBIiwB3Ebyx+cEPAzbBLzfV
S9Q+lj5vNQHVylYf22zXTSzYR1djwXTO2QJpf5CZYb3K1QTh4g0ssUgQf0sh00CR
k2/Hi5ufkqbMmBwbaZr9NVUE2ZZjqrv8JUwPFn/v7erkqQqZTIhFOE1rR78oG1jf
sjMN6ZKL9ZDakXIIzKe9bxZlVonTT4q6bjSarmrSeYFCDO7GUWPVUC3+EAeqETCC
+u1PCKVNNpN7zTjuFana3QXm9aGJ53JiczIZatB9PybN2QZQx+DcSBoCaeXxA3zp
BCQbTiy4ykGff//ZdWx3y6wR3yCBWQnWMs+KmjY96sYJTAHPJ+tKkd9dsL6+ifVV
b2RGxgOOnswJmrZW9DDu7rN034R5QF7LrIU1IvqevpKQWmmpCmtoJ2A1XbajnCxk
BRAohU/1xivT8BQWQH55yQ5VgY2lWz5RxVgUu+8PQ3xYXIuZFBP2QfajZlSXthQc
hQP5wJZQOpUVSNxVLPpYKO/UibiHz79168aO4jbmmWMrSa6TE1ze7k/u+ynyJkRq
S4IKIilf0f+zy76baiM7W2lOL0SaLUmBSpC/JdjS/V+QV7QuTUMK33twcAhJZLR1
eyu9Ag7qc9MZoSvveWYGEEysSjEVaWRvzsB721wjpd1uh5Dy8KiN0UoAzSHpP3Xf
/neB7AvqrHvqwE6nQN/ryGhME5mzDw4bC6/XrfjZ5ppA6LYmwY+exkXgz2907722
Y+iw8Sq/cE0A+aMKWniVbxuiRl+K7ayQkjtzop6sIoMH90MQHnhWZli8zNTmEtY1
Fek0j1tyKtD99S1ylllBQDW5vVCExjimg9P9FlL4Oi+XOP/QPNjzmrnIl67u0OwH
XRynf5W6/1UIVKLw54T8Un3xEVdss/VNd2b1wUFon1ZUITBefrj6E5D1wSpLmehh
7W7TqzB688Rw6gCN7n1hjcHjJBzNxzHXMAfeNVRjgQbb1xRVvZvumDkCKiAygbqa
ti9SSiNQY/4NtZjO91k73xo+UGDFmmcfP03GMQ57/VVD6yK7xPgzXHLk7WK1S7v5
LacWV6w2n3KdAU+/Ludywcd02CcF5kyiqRlxCIAsz/OcUun/yPEGiZUsDkxRgEJr
HB5C7qy8pOPq24V+fopi9l+5B4XAeWY9VkRvtktDY0f0IMv5tQtm9lF4+cVNR1EB
E0K9QpDvAeOsZCXDDd+u132GPPtLxltfDpGD8z4d+9RSaLDqjGBQnZo8+9YCY3aM
3TAG3R7l0cO2iL2SbK9iaHhBvCmNN1CQAVU5+n06J2ldY64mw4zS9T8ykbW0/Eo6
4C6GTCSbEiJwtGuAq0S79Vimx57irZvsB4A4jbcZeu8cx5KXZBvsKoPrISQRe+zi
Ha5tNG709M4YzhcQ0wilzbF+hDo9SLFwDXNUKBZqJaZKCz9Nh0W69q18O39zx0L2
w3yEWe/EmS7tUUPIA+KiXGvpDWfvQwvgsPbLuI9TJ0z+GGOWxLZxBTuX3nFfroMc
wcZ4eNwXQrNdqOfYKdae2jU4jANTOdMR/WpKKQWGcNGLr7jSdtZljhYim/a8M2Hk
1lQWtGyxQU0cQRJJ2vGl+QrM1Uc5hsyEGgMIp7FsMUTQIjkDmCbBbUVLMD0qqbt9
gKod4XNUZRX4OS1phkzaIglC781u8SeBjhEqYRujDadZXPooRrPwU92iYrXj/vED
KcwxqE62mb4ABuc9w09qLHLFsQMClzcH2HL+IfdxENSHomuD1nSYbmwwE3Ng90fn
`pragma protect end_protected
