// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gJ/QwojKNr6vaNtkZrb/wprassBerAIQ//Uc/ZgqmEwyF160cXO0cYseDjSd
SVjRqAJ3GNaXfAsuMTmnHQDPcPqtnXANtwiYN/MyrE3dGtp9vKeV59SHsx/9
JNGvmhARTj3w/uibbWJZ5Y8/gPiXv5zXRlppVB/SIpGZqVE5sBCc7ok+bVvN
fr5dRxCJkpIVnKOyOhYdA1LulIiWlJ6pBbkQKoxfuN9NLZkqiKvfgRgw+0Dm
N6IcDLrFNooyaTvHahjps1xsPxZ4KbptHOdhSmPgenAN2r+2dVFeag8R0cCF
27HBoI/jpY7bXS1BqwTpB9xDtCct/T/L0lLp1l5U5A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Holxin6R70ZUwxfkvOf/uIH6lv9lsnRmfIz8TqpS/aaRJF9siMfmOIvrD+5L
d6FwlsVV7zmACapG/B8qlCTh5MK6zsCytqcGouM0+eS93JrdxgdKHeXVs/NB
WLbFSfa+Bq/pycGEJHykCjfTRpeXtnFmm3zCRrf7biPcgUiAvrdi7WxJDyzO
WtrMEweVEGi6L/hSqrdO8zNjeaqn92LPKivk6egg3cobaEYYv+ssmBPdrsuD
r40Rq4FOeYf6hG5JYWp1FFXvJN9DfL9OH7PBJ3zZ1ayMDxSlI6ELEAWrZl4Y
R6SDM9Ptn3CTqLbikS/68y8YlbyS7ulpL2KpW2669A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bySbJVYXJFpnH0SkL9Ce1OWd850VvvqX9m1YPA1nLIc5wqUvWyiEJQCuwZlt
uJ+YDN1tzZeFDW2pBwhshvePPp10UrqgBTHYXgwhG1COoTknyMtZWmSo+cGt
CMqyzlCmlarCVGzrodPuYOu/smjURad4YS2T0/l1lqGRLXbjlr+V7XTYI8VU
m9wUgG1LT3edX3qiAhkakPGKZPCa+uRVQtUQr5aFDcGEo1Sdo0l/mzaatvFo
uql2c/VptqXKHotqWgN+aV+EdonAZJwE3mNcCzw/gygNyqfwfh07JmgqDOXb
A7EdM56+sT7S9owh5FedMPvJL3qN0MXZqgQMtSZs/Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JIVJWkCXXSRm6yqi2LNmG9dcKbUEQbQ54fkC1NFtYBxpSM30ttNldNk5zhRA
mtjIVRb6ApDINJaK+Xs2mOqwRwrUixLkX8iYvA13eV9xUg/G0V/TZkBi4Rvx
mO+N+erMvlXw/vQUbafcbo2CsYBAyN4aBsGFecSTA1P9XCY+k3w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mWlTFyBDruunog2Bwkllw4+wJ2xI02Tk4626yQWcCJY1xYn5qPTo5t7WKg3b
p3GhPfqoGELGOiECQEeB6kA7NhXqg719kcjkM5Xbcj1gMQoCTZ4WMs6keTZa
aHLRoC16Ia5nDueDSUXphz4GD1CWHj1FnzcTOr9PYIx1uNYYrnU+gyoLXuIo
5BiEglt7G7D24XL8qZ4TyxIT+CCdVyHXm2VZi8Lnng4x7lzTOJVd50JcFjHk
F5586Aa0Z3506ztu+R1gimktetcs30WBoKpIWYLUcY1Exxj1aD6wPPtTBIcy
QLv53ZNh0KzulL7FNaOzSxNk0XBouPtluyAHOU36tYHXltmlcvZ4Yc2m89nX
4ZVOiniQfSmWBcvE9XQhl0CDdyRUpZXCzetJ2Qrm1YsezXW868h/A4GgBxwP
G0v1JmbTJ41JXh5ZEc18Zl1W8HOgsnc+A4sGlXJoVX157qlQgGxAfh6V6h0w
z8GNNXJKHP/q4hKS2RgZrdJCIDUPtCRc


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
U8eZdiLa3YasJ77sjua7vbFkzDcAWeuVcCGKgTKKdSFdyTCNDmwIEgxWeyzZ
7P6S8h8OzLNb8Gof7Iv7FvTDfDmN1s/lpy9TAT3ol9hLSYMRTD+Ebtlt9HdO
qCEckq4txANcuMQnRkIIs5Z7woJaM7yB9vXVHQCFvrRvRjbY4GY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Qj9f2x42t5tHF9r1sLd2KOQ4/cqYgHbmJ9ibklJFIh0mqV/K4BIRKSJm6Wvx
5nWreWaVYRLB03smTd7I8vlj3XIqa7pzW5Zoht5ZmJ9KBmLcE1gBjq88ncWr
KtGTXwt2oKjeuMdMazwxFef7SKF0yA6tgtFWLd4Fkm3Dhij5/iA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15408)
`pragma protect data_block
UATkInvaC/cOf4TdqplC2aKhb2MFnV+Aew05JKKkGhS9+xxBATdG2CJ2g6YG
jX1v6G3YgG7vz0c1jLrTd1j1dXM/AiiKTh+HHWwnX2Ej1moT2408DMZsiF6a
d/Gki7d+k2c9A9zc9Vm59LgZ7sAiwYHDCjuG15pCDliVFzhcL6ynrfeCINvw
e3CrSxudO3cplOMwiAqXXMhR8geiLMFX5xGFjSniew+wLLcVPNGeUpRIpKUU
4mHhC7jxp9jBuiLVdOg8ofNuj05Jtlm/hg8KKLtV3TmSlTxhHD44JYIft7j/
tQgJLJodBgjHJTWXYk6qHRRmr0sNzJ2LybCZcVnkIRZJzdTOBKqvyFocpb2m
vmyhfAPDqwU7JbtQFuJ5sBfWl1B4OHJM8+mKXB3ZQ4uG0c/ieER8YoVYALE8
mXQxYZ7raQhU2th7LaYBQd9enzxZ8VjCbgzLFAJL+qQM0wKa7V3J6gU7nLaK
4IYKsxJzGLs1a8gm3Xt+bRMkf3yXaEEKNBzmf8EDy5wkzVuTWCggetmnZkVU
ejYI6lfK9Qhx/B0UbHOfdmvgEAfImsNY10Njf3aRRBYiwgRVCJ4OgPWzWPCk
29F9xHJ9kXMXEQEdjWePvdk1I9lvLB+miYBjcMfunlAqEKPiz2tSkUctaJG9
q4VvdiQSS8qxuhCW+J2agLMN+fBBELOll+ifZA/hs2JNXw0tF4XvmWFCyVNJ
8CjCmanythu7OAGyZoHwVKNpdgyIh9o2B5YgNcPpOirKQqiWGpWVOj4BlTrj
SaXLD26nmYRxsLfrGPoCkrZoIibQCh/sAXvl08Qk9Lvq6WhSooWUM/PoUDJn
DLFJVpaYWvtQ6620GRYsAUB2I0DwUp7IKa3SsA1ZdNsvtnlZrItotUaxRiOB
hmjRRXf+2sFHGICdhcNyTSnTteBYEOq3ttUnLorf6Fdx5S2uF+TVDzGweJMT
7We8jGHZxIHvBTRzQYf4RFzj8Popzpi4ujdpHf/o8qUBAD/rrRzAWBlfuIp6
W4ScPvpzcg4BXRYsWXudrMY4XsgT0QYsr0FenWcrTEK54P1CLuYf1roEhnH5
U/o3U/22XaSwm+bSYfSDbx0yETJz0oU3h1hn8Gr26GGKV7B5CV7/eE5VmBgj
6PLzBRL6JcQjzERubbUSW5ko4btNo0zoClTq9kCzsW2w7j28UB8Nz+LvSCif
KFSlfqjqFCVgI9x9a9GrbX9T6aReVy93CjofgcJGKNKNnPFaLmu3TmBFVKu7
afcv6pba6yBHcalIuqXH16TRTaeDBIosnxkMaZg6+N7s4UBgjRuiynsjx670
qJAci14+mm9ebNrhlKMIrYSVXv9BlOtHPGsHmjTMWs+fPI6LpssVGZt6sqHQ
m22BozSrb4zU0p64uZwpMf3nxfxT+Lei1udCwBKu0n/DEZT0ZKs4kuLhtnE4
Aclq+xJXqb5DKldxr2lsSvBpYGxNKNjP2wpL8RNAx4LG70iZX7VWKyxRN2c9
qqF7uHfYjkYXwlvrL4LEqpxOhlROux/b3ICnYqwjGt2e/I1ZNxGmoh4sebM4
ElTKhld7Ff6m2V3OP1a7MBCzk8q0xI/DJd6BmUYjTxgrjoW+YBu/jMhWAzgK
D6p6oyEwbv7GtOfsMaXs4cim5vXhLUgmyv/e4e9hBCrpivawEJhNieOCKprd
uBK88Lu8dGkucB8JyyNOHwl2sLkIPmJrrge0cBFhfSydPyuMGCOQ9onpy2vP
0q7nD28L40+UU7uxP9HjnleZwgXQvhYuudiSdsidPscDv8js07vlRer+t7Cy
zHUhIM1Zrw6dLVLMBiTA0KUd6cGLWW913wNjJ6l8+l+mSCo+WSzP8j5RCxMk
6uwBrVxrJvGvjf5pN/TyeRV5RMIEc25+n4xMahz2ZD5r1KajxbkLl92Oncy0
7899rLFv2UlAATVdk5x/GQXC6M+gI5Xkk8yUgfOJ2UkHCviS6OUpAe7TNZjQ
4eHyxeBdzKINmKPWYBXPHjJkVTEV4vqD2jV6rvIMlaP/lhUmj5ryllvFXNdt
6G+hfHKgesbphfEdxllwuoqZrB1rVyJ1ZOX5pC/iUs80CGii81Uj7kBFc4zV
H7kHwU/DVgyT5xSDJjA2L2zjatv4gc5vbL7beuC1uMuK2l8rL+kQU6TQKzXO
ggOUmxRBxtpd31gND3868g3jZftof2pYE4Sw2X6svYEPinpnC0HBPWCF1cJo
yR6CdukulYQdA/OdzgFvy9kLYOVDsCkT53LGAoihnNXn+vNZwnpgbwpYs2lw
0GOGX/E0bkJvOrzZa08XJkyJzs7C8mx9vp8Sx2P2eoHCgTuODdO1kpoRNMth
VDkEwzCcHJqa5jaHCVkFQ4RoCjSMFPnKNrl9XOfMork2gOvhsbbeJchhPGID
Y+AnR2QlM293HxFjAshrw/rAv4ztfIp6dp1mO0crHCujhj0Ly8ky1ziIxXIC
y+YFj9Jur53FeCYfS2JlV0YLJFne7kZY18mwK+glZL/loL5yV50q9rfOmDQi
9SCJkdmYYDQ7wVDpcUVzo0XRb9rORUZNCi6XlC9pqyPbVdH3hMq+z46UXpRm
M+BChFF7Haxbep+7P6vfSbAB/rUWZk7IVJvrjOqoSi2Oinia/EZsGipQ/3hp
pfdYcYpy0HSbZmzk/eFxOlXn6uzKGE4N549gU/6MDa9O2+WNQkPVR92c/Fya
nF+Sn3tUrB1kTSjIb20+00f9HsYpQv63uVO8CLAWyYHsYUjvi8bKd4scUEsq
O+HlunqAtctWJ7Lfqam5WD7YjWUX8nVt4xMgvfHHmVQb5lExVryI5+et20bO
H1nDcOxi25cNuhdbuHKsn7eWeYek/666cD6p274eoJV/Nd0le+StabfNqcb6
fW8BOo8fatcVwfy+URTaPYagddsLhLaeVJ8VeJl/kgCXpnWel3as6b1BavOi
y71RqAaf8tFbgAAOxUVKLgQpZMo5OLoocPti73yI1rL1qPnKyHWZF0COI/c5
rh3VSB/qYREdNBNwcc9qZERGfMain8yWIgKxX4AadNdUQLUc8bEZvAt8dWoj
Rs6KfzrBRBCi1Sq03bNu2r+q6oPohVlKMTx+wWGnbgwf+5PFxvqIFVhETCoG
4Q0dhyFDPNKsMPlCmbakJMejIqBj83nWNqPCcoHYP4vdOLpgh45GvATHLEs9
QopbmGNsQ89ah71AAy0YEy0XYG52nqhUi0bey/9V65qkG0VtW0S5sw1A7xnR
duAK7n5haMT00KNPwc+lSezIzxJypM1r1P9cXZ2ZTFlLUubVbhIFFDxmSvX5
UH3CimEoMdFUbSXoIX/8pDYjagtqVBPA6yziEXpxoXkYaA4KC95fVy7uo95t
f3kaFDpDNF8zYIIneOsfZ04wd2E5pv4ZOTHzgMAltZPXqS79ssGBhJswCr1x
NEDrDxANFvBnEp7CIedtZ9PmepCEM064gsdOmGWhDZZOELyq4AwMqr4ehGMH
tlduuh5TnJeBaaTMCjGX+g24wbW+5FxSJ4ZUn74eo/imrlYthQdsL9cruzQf
ExLvjRG3ChbpbSf8MkrXIWHq8cbqbsNWDMKosu/gxejD/A8SmAGYKWS3Bpme
3Sxv64e8wK9GRMHpHCxpqNjyjEEXtwtABk/SyRTGp61LDbjFKTr9xd7vKCeB
5MGwq5VFWha6xAEpBPDxHt3bs1AlYzyvsETtbOgs4y21nQr/kJv3smkSFa75
Sj9kjIbSLrfRosuqt9n7kyWRACipJBY25awS/75SfkgcH8RAAq01Dott5kQq
zl8S/VWeP+BfSJBK4UEOy0MB3mEeIp9Ctyg4OmWGQAcwGlGUfCp0EKshrimR
4haj56S4VmnpdC8FOIYaztf6Nyxs8L8OENQFmCJcbMVxP6ROqAK7PlawiRJN
YHE60wBzLQFt2ELL5lB7aBvMzztLwDSJLjPhyFvSQas18SZveF9dxIcznpG2
BV7cyZAan0MCHDU/c6DA2xr9qHsiS2MRm1W+KY80EQJoxz7iHSpopJefdCEA
FBvuVcBExz1DO6oiw7WvM00ec7WuWktmmy4c4qHVIbKnMoiSBjXK7FtRIir1
45+sRKK4oZeTPGGnZ9hq4NZCDJcxUB4+WuRemNZxrfo4DhloCvWrO7C1bvUd
zVEBM7ufIXOoPhYvwZVmaPN6HA6vGB0GcDxRz8wqG0NHoWMSW5k+cCmK+nph
UXgSyFBNRiimzumW2X8t/m/o9OA2bxo/MKMl1d4PXCSPIdR74RwwpDseZSfc
EPYn66aFHOCBPOHozRp4kIyBZGA3EEGRABf+Xc2ZAR3G95S8I9bDPgBak5fE
rHIpKPFfuW+UrdRJ9CY/fGjaHgYdeuPJ3930lthwkwSZ34IuM5wyNtjolIMp
I1wZUUEbdCWTDsYmoAMtvoQnthNUST1ysI51xvbvJxN0+RGxIdFT3qZZpZkV
40e9lIEy0wOnqnN8CWITLZaHEU5ja6c2ZJCcX21C//0iMjgZN2fBKsnhEOsW
1m0O5SahFeSX5PqVBAIi9Fz4NyXGcDnmWo/+yEdtwJvCgDvMnmQEcv0O2svB
RkQotNpUTpw84n3yQp2R7pCQBDJ7CvzkidyQlGM932hNUQw0wIC8fglQPc1J
cO5VCmxMUbZcMGpHiQyvW6sTwxxfR7bcs7QEGmI4rsUXUFBNBvDg1iWZ3ngi
qcou1pOt0zA4y4Q2HNWkOXzAO9ZH0Hxe3VgIJmAskCnhDj91Vch/oPNvZZGt
i505DBIGBcObFo7czk7lhErsTatc1IST8iJjIYnpChfFrQYrh/KY3D6+hsEy
P5NHlVTdqx3O+hMTmmY5aMJy8DMoM5CSLuTB5c5eFRHtQfjNl5LEzNiB4Kp2
b+LSqjJJ2I4RMp/PUrGnv0JRLFFUzQSn+EvprRdMPtxRU5/Y5nYz8l6v/fem
vThRbTsMMmKdn3QCKcO4us6iTYjNjgSgEGy/eCmFpTR4hufkZ2/l1as/2YhA
SR+2dVO1I/LaQrBaiFmCiFwbu5fS7Okia7Rt4SmaJhhwGjpsdD7rPzznLTS3
3t8DfIINMfSwucmVrhmMe3iNPmsFyCy+raA8tyHA1up6kTKFymZaZEMPCUAI
DULRtd1/XiPwtQpGXMXnmpIS6tV+2V5gd5ktkrlXgU1Qwz3rhYQBEvBA+c8w
6oYOYPyS1OKqEiPEPoQp7YFLzA9YzbhlHLn/AXJpcVbVB5k9SaNKlzTT7dgw
RQiSwSVNLQ3AwJG3eiAbwGlbvPIZhu0TgkOWWjkd4Ui/lCbfKd5ovTU9O4+i
amZSUIunhkta7kWKNfo+TLZHkYcFOnhEIMCpOxtDp7WsY/l9E8VIEqUPlmS4
k3nA/bLHTun3ZF+XWpJqx2l/vGTHOlaZ8bbjV/zlMCUzcMbGw/Z48qsFbvRP
uokb2SF87xYeDEL3rfTX6N3xY9MyPOI+9hCidZuv5NhjdAONLUKjxrB93a4L
sAgiW9iSDA/6oAXVkQPbQorC1PMRuhuzHjVDWXz1HRWe3dpwP3G/Ao0oJKTQ
Sdrl1cyvF8Hesm9cnd5cABdpx8lRWphUQC7bBruYBWrOYKAbmaClk5721lCx
9SPyme0tTqxBre0m5GE2Jq/721KBRBlM5ZC3luMW0okfYBRj/8fuqjUqTrqD
Eqc0DCkCLYdG6kJnLxdTrqASrk2T9Yu2CrQYHRRh4edqBvn5lgfrq59KOxS4
PRxQcetFi890xqE5Oz0TFQCg8OcpOQsuZjrVWzbV/WPYTKdXnjR3iF1OhBZ+
/hoY/UxAhYXq7tO1c5NyDqeJoOJLEB5eHw0VTM3c8fOetmUmnTvkSWrawv6a
u/t1PgsknphXgsAMb1Zbg44L3cH1GxdfDiKQFO6p6GYqxsISz/s7ZPH1gSt9
NCvD9T2oEFMR9fvmupBjsicwbaqIZCmZD+dgHo4u3V4jpHmPJsXNmC4X7FYf
pG6hgdEb4Bs5+/mUTj9Hd2ee+7cXKwUEV4I52Ruk3NDpzdFGGhqcYKfSi3UJ
73t8mv4QxZon3qw5gDAjQ7U7MR1Li+mrkJgB+4vDhdTWp17CCeUiMX/PvU0E
zr4gV9uNulZ0rs8X8qXxc/VVLXA8cyhBwqZC96LchAsWvmzJCARIDC3lamK9
kph66YV9iZZT9Mp92HYiNkyWb3IpQq57pBDsHHbQXUjO4Le9qxfkaY9nvfNS
CdGYFgWBx0nQQb9E1RW9Nw1jEPwq0qLsTV+IR381Vi5gIviq4ERWEpgZFu0z
kqXZu6dvLmjR/yGlc7OALv1E3Az9EumXzdzeuZ4T6eK8QnkQPU6fuBgNe/AJ
KP2knEgcARlkYihaTnDYIw5C+6Mj6zO5tS2ghE4OamlIY/NV9bvBjazOXSfp
1NbdZVX3y+pkOwZFLRXip6M7TITF08NxY1vEp9PmCXQjyy6HFkOLZKkGn5oF
0OQ0wdBOe3J4IPUy+wloS42UNND7IhVSRmcCd0pWVF5tuw8GlvQADKjC5GiT
dU5V1KzLOBAugucr9h3S11Wg5hI6a1AQs3g8AZLW9mjaab58S/v/W24o6xBG
ePU91vy556Sw4qE/eNF0KxW4grb6BhopIaw0tbnciN8akwVqxcRtXpMl1urq
BpNFjFybPpIrOyUYT2eYeY679Owp3HP3Dd5UgEz5SRhUW2xnS6nZon+K1ezb
VcF3CdnqCsdGrrziHm//jpiY6AkwyDciZhPPld/+dNX0dXbqcqzj9a30YQ4f
HPrQ5OtLjdmv+S2VtOjGmGtLqZfLcCY8H4LU1i8uTJBO7C0AOGYJEnIdHrt9
FwdJtiTAJ8GCz+fV/ogNXqPZIxPtvqCuFdMdibZBjcvhtFQZtbW9duzgMmQO
wx2zXjvjPK2O9eGJComIxGFbtj9TK59s666BO8WTQay1nj+l2KvwR1olyvJw
haSC7sl7QfUAlXNx9Xo83iF/Jf2mYYj0VikYbYAwGJF+9S4gDdH6BdJd8g0c
pshboRwYdRUPnZrYQyGtY0nfmE564vXE3Y1CxpngR2CRZ5oK1Z/GIstk949V
CjvryXekH+D4balVkjJEhHjABwZOixiaj6z0RjhBZIPB2HiUgI+gSIx6Hr31
LVkIjv4ulJiScAHsUcqBALjeWNPRQam+8a8x0/+dUqyv77xhFOJVn9OzFSDF
DVr8X4DpTWnYg0wOW8UFrusweukHq7XpyU7fGAR5zASyJCjjIRoCt+jvMt/K
OJ1rkutsR6ZJByevXTdDtkX0awXKWkRkBnjNFbMmUQxbiqYK4mBLQoSTapOu
c/UVdzirv/oTCRXgLw9AlFtisKFAL+BMJ14LKb6AV03MH8dqhbsEI1wTxdkI
Ivo01fWbYaPL/ZsTF6Ea63Pte0kwx8NjzfCpNuADSYwKPYEuuld81DAOQhgm
WxNdpn1fNw5ao8aeW2FFP58mGg8fF892hMTrTLHlu4HWxwQfk462S52hBrRm
FzHmMYYHlo/rNZC7oNKtYhYZH9pvbpQ8bVS3bESG3f1XhuguIxUOTuCFUr8s
VTTEMjPP+eQ7X8xVoBYAD4C7N73H2GqS4WNmB4djlKBxMPKWODiLdXkmlILt
3no+5jPBuYzdRfolBHNP+3j2KK6VXP8pDBGnzzYeir+GUW9JqSvvmKr1b7rV
+HnOoNY8Jdp6ShuG3tLNZ3n+RcD2eUpVNQ6E6L+iMWiCxUwf+oGdZTFdEGk7
gJzRX8iZ56wc2UaEMsvRwMKe8HK98p92A2VblVA/XDyLwk0DzP56GQ83eQPP
1qnQeyTTT41EqEAIC0MszUK//DiGGIqbqEQU1xst1RIffCfuiDzQj0goS9/A
rz7s1loZHOiTpZNPGaonNcYh3XnjWPrJjeRFmODwaIFrN2l/VvJZqPcjqaI3
VFQQ6npYmkmlC/BEl33XVcsRyIaOViOLzH54L6j743w1KTn/r3AJtE8SBDYA
SOCqzCBNUFz0v3Sy8Wcjp6xSKu+tbIyXn4tgRUABcpLyc5FXCGeiTUpWLTK6
fwxdfMhvUZ20oeRufUtACMh9t2En9s0hre3iCk1r2CqRy3UcYnIm08061V4H
vg0xVMusMj4PkkwATZDU19MqH8leVFw1RU8Ye/tLnarItZileb6QHVq7H1kI
hhBpp0zUocxAr97poO7TosglPGQJgQS9DTpHCCTN0UmzE81CyDssGOHqi/Ds
AJensalPn7GENwDX9vllOpTUhC7bdDWS0vfoUr06RIc75WbiMfBp7yRiCnGw
ZdpsQDJ01xYdavSe1mQY3A00sTeri7NVOhynA5QYfpYXa4zTFJAkHkRekUgd
0rByQdmr675mgvMrihKc3OjNU12xJElYlws+CXXZiF05kT0Gw/ktkt3RwdOJ
SJkox67KRl6JefSfj7qrVqiAru2duRVD99myLdl1W61RLFW5LIfkg0cchn2v
Z5/AjI+hsC25BI45w/0tVmZfieGP+fSefkQANY/izlAO3qmdHJH9kw0vZnEU
BzPdjeUhWYr82CzKrd7OVUfmUgB3q3tss48bQcRTy0Dqqpo7VVUchELrsil1
/+XI5Sfj+AWVWK3UFTxkdiiFox5/uomZOxX3QxTYdrQ0fTntAm7RUKdY/56h
U71Ec02CTAeZIcINl18llOsnvwCGrXJfBQa3tEINEHZWVchejHG4H3t0JV+N
EbEioFkvKCfGg7Gzg0cywxVnv4LSsgNXWuwkEc9XTqhZdKZPo3fghejIeaMa
hLhSEm6Z/p3Y4103osVjqHdKDYiPU3P6ZOhvCNi36+8kmU6fU9kKmWtb8Skd
nSVCFhoXkaMN1enNGN1qgJsKT030Oi9ahTAI72UjOf1X90Irw5h/wgIVeEsy
zH8qJxZllIXchTFkHteV4G4zxOsqcgnxtLUGNDQ/nfPppsgHscc4IlINnOVN
rG1tVxzD/AoXH3Xrudpog+MNRVn4Xi7NFTSiLueeeNO0IlJSe/Ufk0JAEm+O
RuirbPza3jbddZ7cLJaxeF3kOpTUUVMXtWq2KZohKGDcLlqlBlR6MYr9AkMf
Ju6+BvvVByRdkXlNXuyjiOE9qCE6xyC4Vm0yWOMwQZjAZumUWY78ICgDpCWf
LdBlRHsU0KAcMWtWJvqpKekwT0nAJVcu2eb525/2f4420qe48OQmfVqySPhJ
M65zFoLOhx1PqpJg74AnbSuu2fOvKEpd9BzU6cIhhEGKvDvDcIB+fFjZNtAA
5R6+kAEQI2BZ8vl0XK1qwrbIvwqdLeOsjWLIn59BDdU5prFGU4xpF1oB0A1V
C8kH8JQhnrIqo8kEULYfK3l9Ep85I0PUp7A1LkgzeILUbqkjthj83AXksqAH
fbs4TDKw8NuJ8nLGTeHqwl6DJHnzQcQ396q6ll3f9UWTOHTeLg1tX4oLYcBw
Oiiyp7KmfwL9x2CVrrH7Nb448ujyvpaHUAJ4ufEHPr4S/JJzWpOAF6xlUhXl
PSbFLQBB/+/DxF8eBh9rRNvXXFFlJZn5bw95ZKdr2ruSYJk/stvYNKevGpLp
UnkQSWmnoKBrpjpi8oq58DkX8BToCwB2c5gZfCar9j2c7dnmRoaMaYnbZQiP
6vo0SRjM0RmhF8ltnp+BHu2EeLl5BRmyCGgzQxcNRiBr//8/Fh/a23GllV5t
AZ0IV9M0xtfhD6vzS1qWWbe/0Iri0ZfIRG1cNzQm/TAO/2twHR5+KdC7uLOD
DeP8yJiXbYeVrdmNRlJQT4Y9bv+szowCOnnYqR2x65vPH8SiHABNhOLWIvtq
U+lBip4Fv7ioqZxSjusrDLeq6Z2/Gsy7MhSaTk2jhqXJcOLyQ2qaxfzq/Nro
XZ2mZBVVnLRs6YFdlvjwaBMYslhFCuAbCjUWKoFKCSyqlVWTbHBs7SnKr7i3
q/si/nz0QmNKhz20MpaCu46Ul6jz73Vu3rQUW8LgNH1bsQPAVcMCg7ioK4+m
3jqkj2F2JbpZQqKrZFC+jy283zCerdKmu2SfqmNmDqhQ0vdocbW8LUBK0v5O
9S0mjEq9z1vMdbS/8Ce7WagGv4G9weZLiyzjDgtmpQnO8tSdFlrrm379IyIS
GwMP9fTGNKeeV/pe6iR4ha4L5XD1nuNNvTEnsVzXNjGrS7Nk8G14F0yJDGyI
2NevEPwCvLshxq7e1BRa9k87PobgIEGN0oEtJBcyV6C7e71aUb9Jqxq5UTL9
Y1GEeP73hiWe75UTWGc/6euqOxphZKBObzHi48fy7jJRjCCfzkGhC+gJPtPS
wS4y+o0XEqnCHHLLr8C97Vth/6zIWdN7YGE5q985k/cR7b3JDN05eAe0myW7
SdPr780YYWfO+j6NBlIt82k0rEfrSzIJDIhUygq5+Tp2Kd6m0vQNlYsyFjht
f9FHArG0JRIOSVFHYVbcB20zXvuTcJIDlssMIx6SbYQnDb9H7PB3bdeO+Pgj
PGybgyv+A3jooyMLgAFWWWcC23TP1e0sdgykrFiIhHYzZNRYefIX5gR+VfQO
F+Lhr8eb6WyYvrV7/Tnsa7rU0LiqHz8fewNA1wE4JS7jdLnRCq1y1eXUZuSg
oAIXTv32IFmNZQxjhgXNhoUeHk2ZaLQQ1E9VHTxY1KOmHGTNErSNsXKILSZG
hFhnikXFNEyfzWLE9xAfrLxQHaSAji+sDjSLAxkbbWgeoAQJLkki/8WcgCkJ
uFWIXNnPTr0XKybfci6mEX3zuar5Kpi4JT8y81Kl7Dpx9s5BF9XgqqcGLOsH
V+oeUDrZ0pYPlfQNaZAzGHlPrwAKpCAZM5ccxZQpBOFhOLhao3+QLJEUzvVa
4FTGEdYSjCZYT5MCHQjq25ruN5HSKvXR0w7Q7JmObaje4hhgHiJiKrT3/ovE
4oOL4EKes9eMWyWStqBBgx8hBIGaUNvzUzCOlPHHNjZJ+BBv51wTZOnBX7Pd
qDrtFVc0ZWlc/HL5EphiS8+ROQeDpP11yYv4TxXAjkytRmEYNqSjHPUSmbqY
6IEwqfakqRrdxbohIpqP0eucub+AJfwQwXQ+UxKoFPTTWzVtL8uJnEzQfSMz
PgwFQsiYp2CeuedgDRBm/3Psh1Fqzfhs34htCMYWpLzAGzDbx4cvzp5rlYDo
YMDMY6UdJ4B92Y1m65+TgwjEmkWX7RYe6mxUjMVlWlhV/rf+75YzTpB/DIXz
ukujWpZhsQBg/AWr0rXHqqmeZE+xLRLpTq/Ydict2yaEZO2TohNsA7DeCPzt
cWwxJSPUgzinzPxRicgkRp2NXVywmUXOWECqcsVpwWbNbNc+G+InTc6aNMHy
eF28Eutwa18mIe03aIaGw0IIUp5VuRR0OQDMU8oOgaYgr2yl1nQF0A7NBNCO
bH6wAI4UBxqDnIy1zZUzfDxRZD73DAIC0KpPgRBQqo79udNM5Kd9Bt8nSCaE
LCohmGUYYy+DlUuDDd3oLdg20fV/d3HJvwJZsfFx/PQpwMV0BApTyIYgYa0b
I9PL3Ukl8Hs0Yk9CSBa2CzQPa7z/yuYMR6nZal15HpMqGLN09DJRKqtgGnUz
Cy+/4naF/gBbz0eHGccsZqYpyOwNbXfcCvTueCmtd/0Ofdj52p/+06eS9YBq
6t6DjHblhk33kvnSVuVA1f9pcldO3WV2NFXYJ2MTkrazAuziPXrKLIsBhLjQ
GDpaDF9VgVroCjQeovQMrrmT6VPeTibYLzQzt47/KiG1ocGWtG5CpmJ+Lrr9
NqmWQSFQH0dN0mf7yjhpOnvbtWIGoWYxCg/gSODEUTKgyXY9OWxecLcJxKU5
zXv7S+ReIbo1pRieVpakZJ1DhY/h8fknoo4iZoPXqOm3AabgM6KfvX6qRvOl
9SrrY72fcEFkRtvMiFrdyWqJpY+O2JeDRswSVzVe5k19xBHI9sDZlWtRs1GJ
5xXM+HpP1roPvt+Rork1LvEHSaoQIPQu1Vi7rMZdV8+uLTib23MgRzICYLB1
ZgXKzbcscCd0bfuGPENH9QTgcdDAf69p5WIKzyqQgPs9UnjtkHWtoEgxm4TF
WSXN3JjB1gU3hwLNi2cuASZGLgeYU7JCdHlU5wKlxdZgnVebJi6l5vd+Caol
F7G99nMTgyMHGgCwtWciHx2dwukgM/0BfHCF7W4H4ZdMznG8WV2t3r5maVWs
rWiudzqb9cA7bkHbkAlz+W5ey/tyNf8N/tPmgwPxQ4jP6FcKPr7PzTu8LaUH
XzxZ2xyusOqwJKqzNLK2kdx8ExbfLJnhA4/xEeMMtucMVoamoktSMmSTdhYH
QNoyUIm8W6ElcXBuuz/H5DndRYzWjgWmKeGW14vsLXXtWdI2m7u7wSGZpuZ7
lefEUZ1ar57PAzr8zSVUfnQ93PtbYuFUGxB5Ob7L8LDixEAwxNqSYRELeZhP
O/W8bcpCQgEXH15eTTZEQVBZO+2UmNdqhsXQ/y4VTqckdVzy0oh63mJOXYRq
RuSefuCAtNQunzzVZTeBQ1ShsiPAOuIfLe7nbfo9B6L+pUHIwKvLbBsyuI8c
nyaS7HC0T1+CpM41zLrkC/6KQntRVWtkfViOYDrYzzaXEllrejtZC2sNczYa
bqqp2swbuyyut1zhQFk3d68kXsWk/FET57KRFw5vxojKev9/1oSv/tVp/qxe
3TlUUMuS9rescBGCde1gMGpfmUGDHacKmwwKO1OcqsAuaV83IsoiyHuPsrIX
nZoBggrepRcfXqUPU9ISnE5W7m2DETihauEq4Bvn+xC/O63wrX0d11y0GoVG
HXeL/AZ3iIacD9KpnxutcE8i7IvVKA4ZWK1nqVypVFCMM7j5ZJQQAf88nfnY
zh5CxUboP8DGLJXHe5ZxJwWa3zYTn2e0WZXUcBHJ1f3Y56OyjCEypTpTl18f
y3XL6V35BcLbirvmYQtfrnH7+z1rjeeOB0W4FZGS6o5iEbVoC30seOtd/T3C
N55KDSN9ysGcYs9U2HBPYpB9iaiihBpndR7Owvupd/3exHLQ5l+qjThMthU7
K3iWwuUZ0tes09TlXum2eOSVl8Sx7W28iVVCe7USygNnoIle1EVcP/QmPz+x
SI8Yg8ziTzE49soVu7+O2I7BAZpYeLgdrOXhQmEw410f7P3keneazDjSWTRa
Sca8LnHFtnC2aJnoWVCywU1/SFbLAwUl6hlKl76D5QNOD5fv+RBS+83SO7y+
b09sNPgRzlFab4HjAIvXomnYvrX9iehsIbDnbOMlsdvE37vs/0zKypFTg5j4
lXqBGQ+H9mGq06R1LJ45v7hBOg9d5LiszqTHlOXYX0SyxPrcr2Ta7Wop/7Av
iirhwsfnEAsWeveTH2ZhnAQmrf0GRrs9sGTlhp8x/EJi9+WCkvBRq1ECkrBm
2TQ740FV4VpIcKd5I7QKs4kFiU9pJ9o5rv8QBsrzgvooXuqzrW/D0VXdVoCu
JXP0JCfw2tt1B4f3oIJQ+1QMhdA0lnwewBmJ5aO7+BiMMuEhulOZh7HwzE8T
xeewMujCaW8Xm1NpPpcQveKIw7cHR5DyDczxuxCehNiIyuF7rShXZl3nwzzO
CR2qoO1X9SiepQpjUZ6BxLqZzCJ1B5MxJ4Gmv+jZHcjq5iTIVicqqQbF8gh7
2+usfpP0o3vo0PqniDRT6ugeSoWf9PNNnxEmyo8hC9HVj69+WVfOOgdPf7t3
SBl2NGHC8qsig29bRueO5SHC8W93G7sywwsDgkaKgNgmsdRtUFgjFb2ohxqg
wEAla/Z8Vu7V+ZfQgIKYShSy9EMAAylGfDlvAQMhiemI2n7/bXph8GPwzeLF
JS+kmw4aFvaJqPiHSkz5ye8JTMkx5qwIK0uZAFgqvJJCG2kt4xKsOPJhEg4R
vnYnNeUZ65WozfSKbBQIG3EreShVwz4YhsvNdziNIAewzDdYF/j5OyRYjo5x
jxCr4aThW/iT0VDCd/t9nF073jcLURx3dIX8S6C2XpramLaJHNqp5yqzLxue
JirJOrZSIOid0g6Z16WE2Yxlvv63YxGf8BGjmu4nUR9sskk49jTouhojyr2x
0hpC9VkBVoPcWWebab7X81EbUWxSv0aYMlwVNrD2CSVn5w2rILZDGZBHfcOb
FfomAMP01722t2mCiOpSadDafoO9SwdgPO6fsRiEA4tgQcmdB/4rGeK4Qlet
xcZ88KunxbD14S5bye4x5ZOJ3InfEsH/sg3F/3XgVbkNrnv0a3KDZfamVLdR
OJY/ripXklezjr99EyIuNRcCyoqCfto2AF1mOxxQsQofaAFZxDk3oPjxyiLq
ueqkYTbcBmoEz3qRQCI1k/XG5ueOI+iemdUUumBpRGTPrDNUqnRYREzc45l9
qVEPwUcxHH1Y5kz+dN3oMshV6VWdl8xo6QzUZtalUOzzuSRIPYFeTTUoJKu/
LZm1xuSWybx9v3XYd58Nn3uEIbzrNx0JoysfuBbVmscDb5CMd3jbXhKOk7em
VtmBMJ3YUTpxJxEsSzidu2CilVeZY3/NlwSQZ9mZjDrZIEpzPKzoZ96yjhvJ
J/FRwDArS26UcdZ/nU2DNLVF9McPhQ0LIs0CTgEtizFRC1PafBuaV1Fj2kbb
WKPbhyEaKKpg6otjfLH3j30Uh8ktuI+tw4QuujwmWBaZfx0JK6JU7oW7MIA/
GHJFexC0LAhpqwQZaMFxeY9wQ0OI0+nyt29mrC2zirssPA9zuxfJ2ZIQYgo/
EmeDE3Hc4bS+pwYwuH4OTRO8LhqqHsGAaaDyktEqtHkOO8u4ZcX8sQJ27fcY
VPXm+mOi5MNkUIrBCOeDA0NCC2zIchgFjkpjJwOw98UbLQgYe86MNyE3s5mH
2sbR9NFZ4uI6aEcWsSkNxuMKqampGZXu7vi7pVjicQcycD8Ju4CwcE+a30Iq
HnomHraAs36FGW+uBlI8HlhR2F3Ebx+XDKwoWNnyUiCVQ7DqRAl541IMGu4Q
Qzt8YKuUA4y14921ALjIDFpLsDv1HTMs1IgpXROlRFdSH5ZCf7+SpqfRjMk5
rgsUN7nI8VmLgXwkLAvKITWAALcxfVAYNNbxUxnQbxO5FMb/UBOnh80GLvxH
wErR3bTGKmY0hPdSqVfR2mmKM2QmJXXWepgGsS5JYEScW0AJkQqJZPf7t9xT
0QCAH7KBEFPBuBR94WyIFxHCsSR3dI/nbOJwSgA1nhaUCbV7AFhrYHFTEAYQ
xw30hFDZGWelNQl/JTNIN1LjeSgirWBvaRE8v4UgkJ14XkXyWB9NuwToUOsJ
4s0FQeOKEsuEitUbWGscpwebd7i6SEB7Tmr5tDnjUGoAHi2YRfYG7W18RQtj
R+UDA91/Jma8PXwCw0jxFHFc/zNxhdDoyspuHka0CvhgoWuIRGZiiRCbqutH
5XieZtbWHdkGa2f1r462BP3FozmYg3lSrlh+hvC+BqyDeYwYde5r+w4PcIp0
7QsAc4m7QR3iFlWAPdTgVnTct4R66uP+QzxlWyWt8Ndxva792ad4w7lulYh1
PM0hUbu100ab4JUdGe5cve035WCQfhX8bJtT6cqtCnhNQdUjG6Qj/LfHSbgB
YhqH9aURKWgtt4l84trNrYpBI2+SelbKBS6S72TqOlknjndteagEKbGlgLzV
tbC3q5FtIDxEcH9Ly5eKu3U2eq9nktHUrqVwnlVwuaKGkYaRF6bit1oS1tHv
v3hC3J06e1i36ezFgYe+tPENYdW6pk7PTwnO6kiwt/BuI7Svg8GFaGkjHb9c
d1Tlltr8OzURccK+96GZxbYkRYdUUSVBp59wbjYGyytWLcJIFHgJhXOmKxZ+
ncLMIZ1MNThLsYT2xtHIbiR5ThPSEOHipzv61wb05Yk2GdlnvKbqW51mfUB6
w50yBirAiGQRqSXAsG0sHW9nlKlInmR6bwwGa4Fma/fKjkQkURqMDk1sOwGY
F9Qs7TNhXb97863cOTDPV+s3OwfBlbHpPIwMbHk5nfUXGznrKC74H5B8x8Qj
jPKECmIp3cns9oTI82Ix8DpmyTbB49MtK+CxMQI5tcHJtD5vBhQthokz+Zta
RX0pdZ+kfBqYErxJVkaQRwW7xp6ukiGPvlr4Xn33ZXoM9eILRNSTHEAUm/jU
VJzOEbfHRaavYTR+0L+BuOTnPtKRcS4wzHIgKqboLYXXnbyYgPta7hzpuony
piialnzI4yiFKhZzPJAEVViOgY978yuQ4skS2Z706mvPwA+qBKFo7b1jj0Li
p3OBDkNgLwhAnfupoVwKgKqdhM3xTmPwyf6NQGU4lXvh15X2YuvjXvWMs34L
cTLSPvNqTJRnJu54KkTyUHMfkV+CqS5T1DNsPzlcSh18srZI37B1ae5ymRaJ
SmgxBB8HYDYGOoW2mH8FmzqRyjE3h9ybke2SQOrRgg9uCrD3qa/0HdyrMJYr
ni+4kQhITY8tmVgofEJCC3du5dfzlUekaXFSfKM81MdNIUmbwBCokUqxflub
Fsne2mGGxKdivsLdrZy5fguqRZDnAhM5ZUCMe2weGnplSHF2+RhCaXLT/ZYO
nywMC0Q4EmWF8IQYMbV0ClI1s1nK6on0uWRpm7M9ZA7yIEeJcmzoCe4LFXNJ
wweEn/9t2Fo6mx5vhzfDA/W3hhlDj4FS9AKjRkBCUeDTWJ51zGN2DcECWRRf
HeRH8Lkst4cH0iB+gjywgDMwk05kiAJSTZdchxn5NODFfi17qxY6ix4W7pnN
KmRc08nQOAtj5G/nW/qBp/HKKvWZuTbt1TU3cqpQOySr2m3lp9z1GqGx6t7M
ZfBgOX+4WL8MozK2zhEYsqybP48DrsxWBxRhE3rRgb/FVEwPnoFiXGIeUdpP
MxXZt46boL4+eRtevVTX4KDCC+7401FUJJAgC9gZx4qGhx/d2/DGjD2bhhZL
QK66gHkRtf4DVn/SUsEtrUnrJFmHIc0PDX+snCw/Sqcv/yhctCa2UiQVmHsS
4CCQ2XbvreMY5qSc2Zg6PMkT2Zl7agdKTwcUr27jQMxMlKjgnExEaRPmXPgI
//QNaIJTMjYR4dOtL+pbZ7Av2tPuHlFhshWIEgk7BWEIn67IxUHhIo1VBO5a
utzsDAeycC4J1nNEFoGB0DQborCQnEdzJixe4qciE+rsJlrW0mR6GL15pQqv
XBGWmI6YZ4/QrXkqIzoKrwCQEbLGZX2Y6z/7iLmiZkvHeM47UIsJKgxKEV4q
J8uWCySnwcEVgELdIZhcngPOmFuP1ZyT/Sw32ljwzqA/EvUkOIfqgOgGSWcm
AJUKOkEQCtwLeohKqLDdwXGh1dym7X+xPVnVmCdnsxFyPWHjWud8TG06guNN
OhuJF4NNNNWNQxC6rQyXFkR2mgj5Pp0mSsPrSDjj2xAp0SHgOjT1pynBZfco
cONXKWXGRnvtxh4sSmtn31yFzgA4KYWxEsfxaY91mfpT11yRRVWEIU3CdMwT
Nuou/B/YHzNT4A5UHlSpFdkpAgFwHWDdcvrUDtwXM05OEsZO4S+0K+2f7rkZ
BGqBB2GcOIjiytrYHu/RC+D8ywpEGrGusG/EfPl83q/XKvngvx+AbRkuigCA
pH6egBz+YIKK44QdEMtYagc5pk4OWxSgtIz/yrfVyVQmFkKZMnXhq5mkOmt7
nJgPFvHFRq3uvu//9tUH0udYdh2sNWeEIEPoyPyNBsvbwT/lrYUAqxg0uBVI
yqcjWsed19Tx2ukL9SlLwCr2iBHbOvlHVShBRqcAK0ObP4XyPr8vSojYRXVe
o6F+ANBK15wYaH/FwLpsy8xiVWFtfYZl880J3EpmZWdTkTvm88pKptovjF3E
MJDxL6IBYNCboyKjsCuX5CGS6vOWZawHYfmtSy12rmV9QNDUoPEqarZeWbXi
vr2capt1V+inASCNxTj9haqTjVLEJAdr3gCuif28Gc+EAtZHFc9yWAKa3irw
LsSpg5GIehE0iDrfqylKSrG4m4N7dP+4bTmZbfC96158XpZNAgSHkhDgvmhh
cZ92QMO73Zw9bYAX+T17u4kxCBQJtmyb8H8Mm/y8DZjOaDDoHlQ2WK+kwseC
W7jsfphThyt4D23Grvm+cV5bNBZI2b0ryEI5SAtp1LZFuBSRDs2WRkk0naGr
4fSNcV1wU804IWPdPCOg8pg8ib5JprxBR4jgj5NfB+EIUmQ0p3IihK1qgnbq
4tECwMhjJMXoBagEe4tfuBZLW05h+QlkXv7zebCIM9aY+7RTwC9aZZ9obdzt
XKoPyagq+kWw6KenSxEYMkkonHpQrmK54/Xts/rI6hbDFys5CQWMxu/WN6ya
7Yqalyhaz6sM7ItQTKQx3VthSMdXuXIoV7qb2XRuM7F7OShpdubhpLTDUZ2w
aOTNfRZ9O+igWPWCfNHH5915m4i1oRvKmDIsQpSXDJ9ZD5/mUXwKomKQIro6
QNloz+CtEHvOSetwR7zoJ8FPe2q6GIzP1c02O/84avFtt8EDNTDkRlbInf75
d6cbPL12LbkXpdWjYAcDm+SZCXO+wj0695m7CL3jHFwtPkokn9OJuj04uysi
d0jfv5iVeWJ+5vxCbe9NmG63I5xNqlzF2XmLRsCBwMAWD+vxyImy0f0BoupO
wTuTBsnzYTNp1AkHsCbqW64U2YNtfU+PYflklMcyXB6KWIxNzojaEY1Uhd6K
u7JI57XBS18Bajf8rcGPCSwh0ZnI7tfWwqczUHLnqdt5Gji4RgtNDFjr4H2p
JJcQ6Z/IEP4X4vAaR+d1iWyXddlf8JGwHWG5eBrKJQN1inh9KELiK33YCfhg
fyKSRCQ+ZBiktwlefS1c7PqoUQ8E7Q7OpBeWpesTtcTnRATEe4HP1DwazhJr
+6N05ZtmI+fh/WyIha4DUz8qbcJrgrPlTY5amgTKt4sXxWuFX791fCVztS5g
47uv6fkXCAxufA0HJaZwaHMMxx9ZKgcgAOIi/eTkvfi/q4nkBbD/HxR8cHhI
HyR2bZmdAAUHwYzZ1Pj2yFMLWTz/ONY8ST/sd8406PrU41HP13gPU9NPUuOq
ASvwr3ghn4ieyTL/BSRhi6wA5LJBY4wAZa5BlLvnToFZQUWY7oyzQtr/bWzq
ixoEFUcYwOBRhxf1va0R3xbJy4tvPN6IM5JNYyepWDlsQAQRt6kciGf14hur
1czcITBVHbwdkg+DlrXAjCqb/Wmc82oEs5qdV4unVKzanO5CRTdd6QszKEfR
x/N13KgTuXCCzEsva2foSwEJIn+hToUWKZMR+sn+QdqKTX3CDmNsUObrsrGT
IxaiAV/tDdECEbch5GBzxaoOx9oKfDeuE+rDdwiX4YSdCF/USYXk8+Q1KP1d
2JCu+EdoRxUrDj4ZE2B7x1mG8nzthH6cgwWgi7lSlynRMHfjcb5aOoCviwtZ
Ur+ro13BMOUgqhMxTP3XRx5met4Lk6j7DVotJCWfhw0h2y4zmC8n9AZo/XoE
POJQV3RXNy70UyP/CSjAPK3P48T5Bcj996kZYXu8sDJb7j+g8xCGacda69TH
579tUcRhLGoS+Tc6udooPIl+dpFtQl/5sczbV/pGU3sKCSZRwrVoIvWax6Ex
FQf4Myp/j79bns1JPOud312iil9MFi5GWUN56gggCwZfoPH1qwuvxYIW+ntQ
6b3x46PgZklpSiMvhtB5gO/8HCofp/cxObbQJbxj83pSEgtPXKbUkf4jHfOX
P37OWuxq18GZGlM/B0cLaDwNJ0TlLx1G6opI8lY9XvMQ6WNu2Lo54c6s068D
/nh8JPld++T7mc7ER4YKKlMCc9XBqA5htoHv+ZDER4RH1CUS2jeXgLSyFDwt
dZI+qCxuaBg4MwmI87c5oh+kvDgcivzScQ+1Y4vLbJSCuSB8G/Y70Jne35Pn
zMTmrYDRPE3FmblW9oRd4R55Z5xgB6SQSYeMtIufg1XNfpHvrkXCV1oiU9yh
q4bQ2sYo1g7H3PKxwX68oiXvSL+kAOFaL947yT9eHDaJXw8q7B+rHC31Lq+z
6857y/DvcAqhsaSVbhvC7R6WIeOmJ+qxgTW2bqGlpK1Nsuxnfn1Z83UDVnzK
MqUPPSUgr9I7771JnPn9NSKq+ECcXHspBBCri+1CGHpcgizJj74rzb+IHZct
+YEXbI+VR1CLAr76e8IYOq0gcv0Cw/yauIB3caV0xsBwg7o+UnhC5Y/PjVDx
mS2W09Ndiz8A/KE8oVN4lnicMA9A9lm0hYBnkGJljsod+rTSkwTME2JMo64N
gsfwhG3k35cu+JzzKIn4h3KJUukVdFZ+fQwQPoUq6Jq7oLe9YaI3zvyj4AU4
fC1m0nxOlptA54drPjDRje6vaiEym1Jmh1DzHIc/NJ1+yUIb540AvmlGbwJQ
jouqPxuJD0E3f74eTggeXMiPgRyMddMFb+692lezWUK109+EbL7PYdrvlw1p
Bus5ciidvUbX4V8EVRCiit8n0C4BpyEZfdvtsaMMkwtuXpytBfb3eVSV3X8p
YwvNYuYX9WQZW6KtxGirn4UhleipZ5pYu8K2wFoOGyGOulpDeqVN9BrcG99Z
n8dL7quXzkSH9bN1oCpEls59FL9HGTLVYJq61Wo98laoqhZVBXgtvnnsk6yp
8WbvmrVYIJ8I+V+Kdn+JmEr5f/Ff+jPANe33qH/fA/HIBG592qrClymALWQD
6BTgv5sU++eSPdXQ8gPrc4OPvRZbQ6Tu8WvHN7XVDPh9eVo4bC4CwvWdHJyt
2M7z377T2pTOfPSOYXqkKR//

`pragma protect end_protected
