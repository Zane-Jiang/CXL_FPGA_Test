// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
kxqnNlKEe0/JiRqasQitLMSO6ApXiVejVDC5SS+D4V86FRKMREqybK2TiSO6WHSg
4wRl+CXcuBzwaX5TQeB81ESViXJdqfFI+Hv57RgBapYAq5V8NuJvxSu6aEN5YYj6
fV8Wyzt/pprCaGuTuCVtzN5ylwxUoDILkYYCudtsUiOWsoDzfz+ZTg==
//pragma protect end_key_block
//pragma protect digest_block
O0Qgy3ubn2fmz1pm2LuHI2hUEwk=
//pragma protect end_digest_block
//pragma protect data_block
61AgZuvlKVvEL8NrSW7pM2fKHg50tlN3JmGU89IlfpiXHg0lPnIYMJ52f5yGOT5P
vpIaffqD+tVlrqS03Fv4orjqIH/ojLa2+YzIbd3+T1nT4LIgAarAh6ORuxFOuEES
+1Ck5QnTy/NROMxIxY98ab+rXSO5oUVmNsJ9Herxx2mfcB75Uh+hVyUDvUqerIIc
XzeiVa1bu1a8NNts1kfgpg9GHXg0LJTmGqSfdWfC+GDsYfrmytX+PT9Hllr7GXdl
C9yGKleLaEL0dVF9mTNdIRKJyF42AYITsSv/i/07znDqgVI2i05Ncq7Wdiacb7D9
LBT0ufGHQO4IuNGoNCpJkimGqbR1QKuPFnl3vz9Xs5Bi+3VPoZMGKYycKYJ3IPWP
ih6U5WC4wA5YSK4zDM5QbGsTDQds+ff13nihMTkuR+VKh46A8lQTiNkddQS+KUX3
RDaZaivGAQjTzmYzFAzWtpLbEgBJxi5PJPsXaD2dObxzD2v0G8PNeJJGtwEdFz40
qMmMrtsDyp+2oNbXsGbhs7XKORJK5kQrb2CmdBW14MVAwrFsOEKy997MtpY/rxtW
9JqpFsqvpknt+NQ4aVeN2mDew5cXqs703zjMzVfQ7tLo0jgvHOckCKRLX6ujykpx
dixl1rYzA8c6zsSgqxpoM29wUx1E/+y7qiQjCfKf2lZM8UPxaAdv5nFRKtbNRF/W
aomlxv8rbvaVsNhSJlRE847chkJXx9/fQZz/k9bVs2E+jjURjQxCvOWIka1xjCKO
qccCfGDCuzcEt9VcSh7q8BYudiBwELvgZqO3ln8F7V31xWAhkEFm6kUxdJAUvNn+
17sFix6K91R85nH4H6X0qVSlbBYTOmZKzym4i0X4EkB80NLCfFwCcJNKeSnwJJgY
ZTETyovy4rDKJZZ1ekmw5cOdxwv/dFXy/vfRHczvpfUVY6JGpe/jGv/krrCBl63D
x+EhU8Mw7Z7pKIfVF5q6A7Q067hkQfvDiTGj4LTt5nIX54dMX+NOXPrmFRCjrVWc
eXYuWw6yKNNoZNpzPeRzsOJGqlWQ1Slk2rZPo5OhqQBAC8rFNyCTxBkBu5SMJmHB
QwLt/SlaJUlO9UgH3KNE0UYATFvblreGxQ3cmih2USw0SutyxNOrreBk1ENO3khj
uc3i0llPhtSODEa9Xkb3RlsNlxgquDCFo1koX1b0OE32esW9mYckrQ41jLBvfKkW
EI7c+tCl19keks6fDpLlsTL1uhBIhty4Iik1T24yzbEbZCH93ac5lCEarj6jyzUa
bz6wI8zOiyDnQJunWfSsCiMwZ9NTIzarNnkBRYf+5XmFJpwkLhxB3TlYAmHkQp/f
sGN+UlCIbx1f4Wo7ZFI3aA06GW2tXVy8Bt5321opmKBPdLIJdOLj2HU5NrtRlykX
fg1AMU97kk28crODOmckBWYVO51eNlusLxSzebJHdyBE9O1DFfK2OMVouOwjvv6V
2e3DR9hAZVaG9v109rL7kpRMxy7ZG5P9pWYgwT+TIxJGZk+rFdZQA9aaFVKsDY4C
kHErjN8PAlgCHoCLbYdsi56+zJaNQU9WMBB5tBFe1XCbh6sMUi+Nc01kP7/BNq1C
RBOJoySHW2R/d7NotQq69kq7SVJYHU4aH4FwaPG3ZWL1gH+6BUQGcFTDHaeD5nWK
iRDvhilMR/fKDZoHVNprYJFqVVwxuxv6be+qLm8V/HXYFq7KjyyrT0yaTTuS4gQO
i4Xb6t3EshDTO2gb4r832x6W0oXMMzCGRegoyutLmsMntnTJUNrfkThpky/f1gps
tIo2R1XE2RoTeCW7OC0eCIhxmmyLBx0StddZaE/vVmXXslp4SqKfBnIjkFzlTWkf
DGNjq8RNnYXe7g6Au4qSY6/4b0KfP7VjwphT+thYKMbYg1M/qdK0SBchR5QlnGsP
CO/5bmB8cRT2buJBsoI2o4YeI3K5jbUGCgnSzZcS+6YH/AZfRe04fG5Kd9oMOAjG
zDM8XXDmMLAJgtGhq4VRPJ2bBpdztGWmZogeXoT/cUejGEz0O2JIfBs9uPYWiKS3
imYYoDF4gZkD5H/awY66GQd4CS7K57dHRpfOZCNNB+2ZEgCpmNIZlez9/53jmgxx
fOamLNsE6Pah9eknZjspGsGA7+F/sqEB37jARmjABRNu5CnimIrwEL8kd6cj9piS
lJgBK+XzKvmTmFX0xR2Q60FeB6WkUsIJ3lr34keoSGlC2ycn0IKu3ONpH8Hs+ojX
u8XJD4ze8AyUbd7idVC7TT6DHDNzfBs3b0X8G9VVUDQs25ernrVPmUym+mMqazwu
uvlQNFHLeLKMMr/R7VFrSy2r4uo6j/dzndrTRJYUC88dGRH8isHi6bjYL1HNRYWR
bWPCT4YCKjrxCe1aqHx2MMbmvgn95VSgcZY98qyaMueWppDB+MgG4cEk56tjL5AO
JbjhVR28fvn/4ycnHTskoOpsiVRcynUQi/CAM6gMrpN93H7I7W3Izr8XwWLEgJwz
MZGQQm/r2Gk+SJXr51PmiWMQYEbKRuDa+pJY67Bj8Co0bKqeWRJ/gjDlgduuYpui
eJxBG8C524MsjpVvCJDUT6dgEc3oVMqaeikO5eLNgdAQUkW6hixkok6yLg0bicR2
hWTxQimV6AhLLbVQdvMoTSvjn0ELOWDujTax1VOh1Q4QUTL+MfOHtGwf75GqpFCF
+X/RV1400uCqC4duU8MV5hOuCewY4lJTd/paNy2S25NGMhJwMsHJGPx1TXavnC+A
ts3aafNmco1GOEtmPnhGVdaIYZftcJ/Dhi+wuYtDoCMADUEDUwcP5QjM3tAa1HOM
2X/244kB85N/Q4zGQf3k8J6mmqLufiQrS9sGJ3NjJvh+mBCiy+COFunbDbrs77bP
3iGfhcjVobTK7YslrREog1jJ6SK6xz1wxqQ4jDdwyt/MKiKwsacQsZ5HZXKumPnG
1s0wtZj/grLm99/5R8RUytolK72hI/xd/sz3wi4MAzTw4DtvPMB0wvvY8XDmYdM6
m1LvzJui+iVL8dDJYWEY2/+8HaXwhfOQEw0zeLvm5Blv6HiesFUalg2qbAWUmfo1
juVJrA6rbZhsz9I3jWjDAw+N4kM28lK+X+hVzB13m1Sa2K63k8MNzi7Z154SGjiA
urglsjq9K6dGpbXHL/ul3+q3M+WvZlTw1FAiOd+WAqOo86HB4cDfNjx0Ji97DZ9n
eUccS4sLWfYGoJX6S9we0iCH7PQTZzOvsm+a08+tNO4f5UlpavbIlIGZX9IuWAJo
vuDcqbcSpxalsm9NwV2hsBK1aHpbrrYLwT61wAyia5usyy6YJq8a5l8+s2QfSbIY
NyVW7rXTrqSxAT6UjX15V3SiZdELePWRn4am4QJ/+7CzPiwiV2JxZqxsqYtzhvwM
a0wcV9imk/BMMqlyr35GM892cGvW6aSigwu7UHiYvytHWzVyDkkvUcwTWR0oJDLf
Op22MKFTTikMjVsHyPRkEhftjuM0rIDMQwCDGCh2PyAweXa/HJf7QHSX5VWlkibi
ZxjDYg8vZN/LzC0FubXIoGGgmcv1x+1OGu9TX35RmghlnmkNpAozC/HJwDT8ChVR
bWTNiUFVxAoEKeao70ZZO35ybpNByH9JDRV2Bo4DxIJHLcqR/XMfX4alAVUbhulZ
U9fSIuiKlTDQmjLhcPab0cIFSjYS431h72oJ9aM1uxUIzpIVAUwjKQAcqJVrhmpg
+amOjaK+eDZbhGxg0fnfWxhX5kWWZJvYS8t60vEFnucLweh6JLA9RNjGdeQHkEZ6
d0PgHoLV79J438s9svmr2ToFLW1ofkNFz+Ty4I4Qrjt30oyiVaG8gX3BU96mF/A0
Cq4fxFlmTsDh2V9TaTP1ZJPpl5gQnRQJ2iW2noGWyienKGlRlEUfWfZ3V3t3jXOB
0P7n+yvDciWc66dQPAH+deJ+dn1CSg2KOntn9UEN4ydRpijaHt5EWqJC0Uy6cVoo
NWtbUPYOih6QbTPMDlF9zcpaT/xEmIL88mrKKBo+DJv1y25ymUaW8uWnxG4eWuvO
SPaN6h1I4LLPvzi434ItlZ1xxwKUW8onJClB9t5+KztrpAO1Fdfv+KNNDIYVaRf7
rp3HmSqPRG95S70xcHqGfz5AUrFbNfO7Io0O0JT7X3DvHEqBc0ae4f8nFcp5rxf6
MBPqa/juYlW8o8QvvTca1IM04GSY2jZry72P4fREyuVxoWGP1uR+mSziVZ2ih+zo
wOIz1c7y7Qm2oK0aIj/XRDu4Y/DFdtwOdVg/ZXZMxjTRG/IFxETw8JrI7cAHLTI7
cw6gnDLvXeOah1CkZvWLKGARl113/i185cQtOIV98ECSaLsVCA5YU2B2zOTzpKL7
+BGpkgZde4tRo1e6XEJ96vY+suWpQcfUOwReKqKryPDpoPR8T1Gj6UJc5tywKw9W
A0PPO7pI7GTLe7pETufSnbwhIRrKdXoBhyH0B24fd6/uCOsB4Gb/jF5gPhS3WqQr
8wqC3/9ySbfArNPlBnl8P8BAe4Hja5B4dMfHZDbtjB3F0EIVCHqVF0nvAJDX3Ma9
0bHj6/4FXdomp/Z7X0POsl5W/K/tZ7/dOqx3r/hJZYu/Jz16detN+/kfSqWLX1OJ
aQ3ZwFIbQNIFBQhl6iDKcxXf/OXiiu7r2cnPbVFFHwnZWLHpuzOL4Ribn97ZD7cM
CT+hzz4gN5xPoBqPsgkYxae1WhdsZ9/yOgRSKBHeJV4E33Y/DbLH58DJ3AEioy68
EXgi4iQN2bPdd4jCQ4FYVWR/PcVlSeGJAUVlDdbE5uoFtJ6KWaABn8pjQR/6/x3V
ILMjP47A39bAvHVWHygnPem15bO3qkPX/panihEjtnzAnjZ/UcjcO5QPlab4arLe
VUdi3ZDfJycXqBbyTO0HFW8b0r9cwRxzX+qi06k8WzaI/r4Rup98uxpV707C+iGu
uWQQ4+HAgNTTb4WUxVuVPIUsMKW45FXQ+06cjYHuCeuxU6j3P0EofPdF8f5BUwkG
YA6SmPyS1QXOyFalNXUcFmWTEJAqtjd5TUdXufRdSEbkXYGRxsCA0pvm5ixnwdxq
FaU0IgsX1zBJISrS+Z3WvYYHwg+a7xsVJBNtL79/680jJdfq4V/Clji6GvJG43dD
iPm04aR3GiQHWXgPHpcinwNGgo9BeyqUnEhsU+qdopFtiI3Kz7hhATLRPlePfTHo
RtsNB/KKbbLFaZKXbQ4WW5h/YR4uw/RUkOEaCxFO8nnNRefkbQlYxeJ7bvuQzk5r
yJtXMgzQuFBy4Bt3zZjSnzyQuwxpXYxb2FcvxufiJ9dv/FrEk5dHedtV2fEtY2Q7
2eiokAfah1zZZUmuYQzdE4nrhwaIxds12mnRGVhIhgXq2srVTY9yUqwHuanJafd/
RMD7R46injVbUaJWbgFZvp4PO2y+kp23+kQBfIcPryKciOgezyQyzXJanyZSATZb
eUswZXkA1CVgC1MSQ44GiZRspl4pX9tWevHyu5ggbQ9MReeBBnBodKQSkCDta97L
WFIXLNXdm2OaQRdhfUQLbJUdYWD+QZ9tZV/VzGYLVstU6n//mt3iDJLTk453MVG8
P2+Jnq0BfJnZcRjFnaiZIwnku/CEh1/cIvU4YoBnnaHUOF+ZTgHXxltxe9j9xzkP
7C/7jmsTPJlrdsC5nm3I4OsqhLNlEf3rb78spq73gRsPh5X5jLiPTMeubCxpQtF+
3Y67J7KtDMeDFQ5Bxm/dN7PGpq0wZnZLeM50zJOCdoNEXMnSQk/6JRkLQHBimb42
bT//z/g1EKnAzlZgUjMQTxkIZNA8x4FmSe2ZMEuz4J7db67LyFSn4nVzeWbMRbaT
zcgaZithErXARjYbvDkE6dAM3WQrOOir8VZgHnI+wppeveoYI+dAZWHy52h6Gd7i
IEYMbNl87cCMsvtie2DMNNkhdy2m1RqX+arVftzsjUL/QcRNKzwa1MfZloHY3aWo
SjSWBs8NoXoVi0Rb8EUtRiUbds7o9ShaHmqTlUxYmFczat0MLPWSGQICOl+TtE+L
XbcBoSVz9krRfNywluth/g5R+vayjQwIyLsT3pMOu2FUzCuwBAYItvMsF6Efq9Uh
/BDMavMom9JRuszEs7iwosjsr9/wTQmcJcWTodtU5rQ7cTdsEmVjTR2PLuPbOhN3
toFbXO75z6u4bxe1TH5dOIq5sMlquC9ifWYGBOzzHmMKuxJ1qc2KH+X1I/KSnFiI
HR3XPnkabqlMvu0hf2C9PA5DEBg7x16RxAuFFVMVVj2uKfmEQVVqI3YNS6+vYmTI
lxaNuYYeiOez86JQd5p4kLd9ivt7Vg67+UuN2kzCJSUDmRH6H1B7Qx1E7QtDX+fl
/5UvTRmAX+H4U4rz6XKcPpxMJP9Kr5Ys2zSgDBP7JX/P+m87OgdyTSAdGUEEabeF
Vl9h/cGS1GYOGL5SxqE9/zy+5XmHQ/sIfAr2aA2eecL3AwklXlOLxCLKU0nLoYXm
6r/61bliyF4DvUM5c68gzzZbzJ35gn+jbdqJt0OhagITdoducRUXY3Ll9owEGZls
tx1/xmx3vVo91nSJpw9p4UT92vnbm+h03p2gNOzN903ZOhuepMx6DFBgwRFI/0I8
c8b2XlzsT2jOkTPhzfQT6rVN/ihy2/5nl9h1sGx8FkcOKvCovXdQRvHTzxvf5T/r
htJiKeyy+ocGi3QpG2ockb/kVWuj8skfXYf1UcSd+L1YXMX1C2LwsjJHiq1SiS0e
2PgLZZMwL/bEKQPqAmnVUOXoQKl/rIiTWIOBZXEM1ODP0W7m4j+mRf6MbEdQFaxV
ZnRvwsLXfDvNwV6MIg2myf3rNVl//y7e5xojIg5djPRMn6IQJaJVWxcnDfDY+N7T
S4ebtyzm/GAh68EGbXaUenh0GudLvvqCkvvZsHyVOBIuOPDI0Y48ZQRJ3EAknHku
vLs+dHaxQiuU92edftHL8iZoCFXS/qfnoTuSWWn+K4uMlgp/bmPBncPwoajiaJUD
rKLhLh7rPFKiW7Gg/z6IiHUEwXus4EaPO84zf8Jku5+ZOv/A1nbj9WjEFTFtXb33
gmtaWI6ha4b9VHMaqllCDskD0LPc9p6+crrf5m8GdyFNJzvYbB8OvUFwe1DX0Qxd
LleVMcDYChPK0dMTadvlSyAQ80QpiEiCiML/XxIJ/zE/P56Qb4FcLSZByn3Itsee
274UiUXyYW9UspnrnUBJvnQPeiYCEoNiMOtSXF20Appt5/8dCuezA1prSCeU/Aax
GI97BA+IK38mkN0iaRWylf8V/0W4mxU0/w0emU0oH2yrkLuwc0n1lP3UHtowv4+Q
41UdZ+NTUXxYU1HOgYaa8KKsMG8+EcpodjrE5U8NsyWbgtdyBM1eWU5piq8LsPZL
TR1BCR/upYQ5CzjPXgtHPasWJSoAnMhi4PUCEbzTNYSGg5YJMLL9Ds2j6N/lj1ek
y1I2NEXunZG+vVmPUNlOw5rXn4rWVAQPHYYiTSSK5zrr5I3FQWXN3YMEC2AVK5Cm
vcOYVbDEZ3rlh9RFTs2GDex6fEY0DZp+MQzW6r0CBPQ2nweQ93MHIzNdhteTi1mf
NZmfYjACESQDniBUPBWCAYwbQOiuTPhxO9HkO3H+JtdMXLbDpb+fiU9fTj158lew
svJtzz51G24ahd05hPTovBGlzMRrmSyrzGD4s4hdoqlIOhFBCMv6ekvnTa0gQ6JM
5aOdsmYk6xBbVjKopoS3s1KaaDGdUznQ2061Fzx/pdv985RGQBgvfsX/jrvD4Ugq
qlzaXMJToJfZeljuN8hZ7wSKrYSCbWrhJ8MjS2gy/1bnm5kVORsgb5nw3F3hd4J0
w3jTo5UHt4tOSZPn4kXyj0gWgxCNXsIQyduZ6ZkZl6u3EtbNnnV6WERnZthg0sXu
g8+AmqVUOwn+DoKiSY1kT1v9jFT3/NTOV8nfAuw41Hz810DOQlRYdGOXFQfFzirf
kUm4iEs378lS3zDRAzk+ECubT+mx0Jt+Pd8k4A0/481uA03JGXyJNePJDXxGstZa
iNZy7AxnAsBLX8PrIJnFparpxOFZNiuHyiBN3PzRTGp4yjm1Carvezh2Bog1wTHt
G3xpLGoo96NCGnuR9bU17kiCU07yJnXZ6OiUg6ZIUCaXKSplq4KEWR8JKeRfGCAr
zTwp8qkkG/rxbjLSeILcNcDGlJsPNoQdz7awLSc67LPWMZ0SYuolQkfo0hQb6TD/
8MWG6/9vc6NEAqrq2BdeWxItwGlPZWm/9CYcZdl6tfUVmgm7eD3hmNSk+avkdWBr
BcAofvQGQLcUqChkRDFuDKg7h2xdhVoOw8mLDqeuR4gVA8gYBga2bB08rKwVxH2h
gUN/S/sRIwlfK9oE7/HWSH00efNaiQXdaTeu87lE2JtAlP/DDYhlmXKgvxWynbmi
CTf9TunA9eva8EE5968gcIpOrG5Bt5HIxjT5yvMYfMKQO5cfYiAthjEAH+fFGEK1
dTomW0Cgqj6SbIqeyAPT/vgdRUlwbhJNzmQT97GalSPUqGemJDYOPzZT1DXVOk36
gjE6AoPtKy+D3piyWA1An69vLOv5ZlB/IvU6ecCzLgUtt9vfnmWNOGKC/DoCv0Us
M/HnB1GtWjqFF0EH5+AnTWWgqT6Quz7TW1IhJ79qy05GDI+R4Dd2tfhqG1tNfrYV
9CrOl/8Ez3ArcnDaifKQ0KU0H4SSoQ1seBckBFBLFYy90O78HLnLEquJ8u8UPbPq
EAUIps8o7hs0dg9k9IAc7wDJgjAHnE1+W/3fxy4/GrydODfXI70epP9fvcaPhHqG
buUSNANp3XytZWzYtBInd8gEnxwYYwmqoJP0gfF2KGDMjnPm+RsNOsQIv1LgaDUP
uM09GLzgnFfvyF71cTFSe6QjEaV3d9H/bjRSkQGhLQOvMx7rdC4nb+4vT39t94MQ
AwyV6Tb3nWP1fbKcm8bp/L9beYWbg9YURT7eaukDHeLRsZ2mj+2Ueye/Hqaml0QT
ZQXhn7lVfeKz4XJIlWOk67mfPmZwwfh83yGNpZMxf0ic8WYw0UGV6n3ejiQ+k6SP
RZ46aUflwAdcQ9aoc52kZ7B9ACI8Fjri3gandk27ZCMyxIwaZAlf8iPyEX3xVdft
933e1i6EdeZZW4qTkszhp/15T2ClgqWa3GeroZUTgQFnoLXL/Bbrc/n6eUr/tVJ9
tvtGx5b5KtCOmtj3ShuXj9dPjxB+ceYQs0Hp1UkkL1mYxgtONpd3CFb+7ao9kL/G
N6fr9jft8giszvTzP1cpPZvoVyIjx7NE9uc2PQBkMiXubowMCEoXuhrNvihTBqZR
IRGc2UfpjSCeFdCf+/lv1jo9klyPalrg5b6gJEBqxFHifTE1bn9sOOwPuVDLoM4m
CVWzkYFo+AMg3N0Sa9Zq/dl7vVaELxt42c4R5tuPxBiIhmYJ6aBFz5R62PBqAyeD
BvFYxRnzu1OBQB/VfRl0jRmXh+n4RxyQxZD2mYEXzGUCI7MaTddLPmG1JC4j/T7q
g3z4v21jZEkH1jrs2Cy+FBHhBihaF627DAwxU0DlXbswJggV67SomCjbNQYiE1jf
n7JHBfdfZuR1nVsmUhgcAVZ0VcUzbjKx3sbWizJos6/GNIMyrxFJgFzYhwh2v1fx
oSwVQQE7p6uA92pohi8w2jJA4KL2GqOOu6iaRdyrw1+Reu9Ivjo43Vq/ermEDX2R
dSeR4pGPYmCiEwk9aUaOslCWYqIDXBAi/+ylfzCeTJsM34+fLtWIWu3vPHidkY7n
nnGbzKH7qQ5rqLlq1VgRyjnMJNmRf+wWV+HKIYE94+y/Ud3o2ix14+7jEq9ESFMy
etvAN/vDVLswv9jTdrjNyblp4pOHOtgqBmN4hS0Wt4UGc0IhGLlafOTEP6ntFG77
BDki5QM0SvhCOBzxbXH9RYwEne8Kq0IOHl2dZBimaBVoiO3NW5uoiXo5wHOqGSrN
WeyMvXfhwqqRQeSHqs/SdHX0uyp6KRM5wkN4Vbr0c3KHrFAC65rjfL56qy4VSLGF
5DcfNl1wBGQoYNmaenyuF3mLLRZZfXDglD5TLBMEAFTIbtK090eFX3jGwmP7l93n
8ENXE5klC36c0xI/th0kKU5UBP2XqJObMNt7a39V2HpV8dLBwHh6Zke14sh2cvCe
U4olW3UOG8rffS83jVKmWhH2iagpYneHLHQKjVtrpUjskQ8pE734RuwRj3lxFsU4
DV8gTl/IN13O7Lttwy85W4XS2AkxQtZ5N2wR/ttMi7cE95Wdisiklyna9wUXPp/i
fA7PgiqenAYUpkvEZbhkMdu39xjTW5AwL6oEZsdJZrTaThGTv9Pzto72+qcZHwyj
ycT41f5D5vkzIfkLA8Sd+25J0h0eZ8+BAOYt0V6kAHUlj2py66PaZf6PHKa42Jpu
RWbPmKmv4cincwebdx643Pao3LQOdTYCS9XnWSq8sPT5BDfNnuhefbLd/BcIV5AO
/8JqXUBqAt+xlIo9Oc6R4JdHhWkNFWqT8CL22IS5tnqauz5o7Sf8PBkDzk4sSR4V
hNP9MGfLsqPsr3Iha56abWe0JxnNxOg0PMHFbZL8OejJgV11imBZqs8xg7FzXVTT
JTVceRnJuxFvk7ijmJCtFpFqaOtgmBoeac4/bmg/02ZazXOiTDe5Qax9ejVedttb
T4yKa8tlpbfHnwx214pJFybfPrkw4FVAFbyw64I2UF+Q3NsDfI90yqSh/nsURygr
tMRazhA9EQwfP4RUkMBZHjI22oHoCC3Biv1oU+nMQlsD4wqdtmeBg0V1PZV5gceo
Et8hzCsem43LvEMY3LB7tCH0m6GOwUk3pxAroVkPtRc6vNL5FVAZfCK9I58/ZtdL
q6BPxhJdXwtpa4A6AfYcGEXn+Saq5CapOVx382l71k0OtplVveUAzYKF8fyIZQPW
Wk0NG8K7s6uwmrkdF5pNkKUj3FL2cfzHzMjUSjnzcethoMemkRZ9qxinC0iCyz5l
9j1w64xndWg3wrL92rkYpYHEIMfmkjXsPvYBJUzVO+XU56ch5K12oacN6mEJBrZ+
3ZZ0BZwx4L0XiNUFH9tlI+Rk8snEdnJxWZwR8TARwljAICiHy4yRoQ/8TQ5cSo7d
UPFjHJ+UQOsauXed6/zWEz4VrAV9azWSvKotJyn4+2U2WxFnu3Cw7q8b0IvCoytM
QQSPsHumviosJ4jIa1/67H+4WHX0+OED5MqmCkW/Z/ZqmMSo7QaY/lZDUGnHIYVs
qbFGJBGlQHeelY8XTIuWLuMpTNDALLPDS8TE5NgNr5L+6+neRPqjRLqwfv58Z6Ko
VBCftOqeS2AZ7pL5XuVTTvUiIIRytC3trdpHKhq5qhgaL1E+tjqm0tRIy7w6Jx9j
cH8g34WZTXb+jb9BrO/d7jBbq5EUQKaeytz/E4mazyfFqgJeux+PAv2Dk28JxJZt
obL2ck+Z9SeT2q0X5t2KgbgwVMDMnJ9bx5V9UMR8aQpwXuDUqyyzR0li3tBf058a
c4J2sLXuto5CCGcJ3lsR8qOnsPrM704CKwaT2GNdh94OSzsrfTGMiAKFY2WCMWca
gdwqjkTpnVgJn0x2oBMFU5PU5wjjUeysJd39cjlsOH6Iluzv3hw7ot7jWS3uEOt5
ZWTiJSK+IPcxIsF1q6tEcE0R85+8zIUexyGwE8xBTMlaPJD2y1NSOLL3pTjAX+bo
zM0btZrMD0zUNyHjjvG56LZIKwvtVvoKxdngA/9Qsk9jTUxepC2wJ7Ai1J03HXxq
hMleVXvjSQVON4Ksl/0BaZh1KrUkY6O+VsGlL/pwElTwFKpw97+Itp05qaLX6pM6
S0FPYlnUzqzXfelLsdVf3IcYCoSEFCp6/8GirKIigeqkg5PRBqkBjNIXtC9iPHRk
+FynMKFbFVNMMCyZdjqEtxyS692N7cThEGtMv4Hd0CRxbI2VEgFqdXzv6DYjbsgl
rgpHqA1o3P2hF8JH+EpgkDLL4CZ5ushGBQWAxipKlm4a58iIKYYbQgJ/ZMhawVRE
QQoDw4MmDWpXR9bHfr7rsybK6R7wm8H20+60MMmC0Nv7vg874lD3fDacKYdzJZac
reCF5JfbwHBmdSxp5XTbFd77biSJSDe/SH1AkHZZG1fmNcqr/jBDvdTHLI6zNuu8
kPc+w5BkKa3RJ7WcLqZ6vowR2IXlGJwIyUXZIwy88ZjzpJ/nyypbC6gdFKoOqHGn
/EG+0h56vTbv+9rDN5wxTofCZ7StTvZUJC1/Hs5Ct0rCPvqBgpbCBPjvjll5Uh4V
kCi/nNWeg9SxFx5GI1Aqqiv7fiW9DWKQ4Jy3oNMzsWWiyYO60NSp/3x7w8eloGtg
o2ZcZrYTc4tZa+MUlhNIKHyLYmqnEal0ifcv0iQapQb4DzWY2HcR2zcGc/I3/xlg
LtuwSd6a4WkHHqLwPaLiXM7oUJGfPv/rBPk3MqVYP/grNBUxLoT6gvkZpVKCE6ug
+by6GVr0VUb+E/R73KIoSbJ+YBwV7Mgz1e1YfpBCygNh+QOmMOEY50YFpizVtFh8
ll2OEOSb78GzlE7y7RxxDc9hXq8BEK4Lf4ngPMqLxeZhdJXnbs09fhnGpM26GLR6
xx5KmtncalFju2M8dwKz/FWsO4XAF/fuXCyFtkMnfxPkoj4P0uT7rkpVaCRjjJUB
HC90VsWUNzzeVz0OpphdyJeO5z4UEo8aZqSg9lmxIh4jz6LyTxF3vS24qwL1t2j5
vRqczS1pkHgyqmIq8mPjd+Cx3q9A/3sScqjQXqgtm/UHZOGFJ1NFwfGsmBbHHJQ9
vnSnza2BQZWP5GkoPBCVo0Nz2mc7hNuWJUgFLu6e+s+icrOaxqYxrPyQOTH313Ez
PkyUjpoOY6RikRTG+DMGIqfC+SMkkYsA6JHaqVTdqqKRc524DHlSM47y2Ijavi2Q
r9O1DREK/3QoVG4+zYk1rK1ElhDelsLExXs9FC+05o6AcM+w9I3bTp85oST/CLwo
/V7Gc9E4A8SLR0SKKehQHRi1gv3lWTNL9+gNAUh6nC68yUSuxsTkL8vMfcSVIyNV
1uXpUkhJ8c/+eBb9NSfZVpg4tb9h2vWHlX+79Xc1UmkkHWhT6oGUV5CJiNlZXfKH
xmKARqsnL4s520Mikxw0sizDgN2at464WDToIIXXNCq/+6Y5DuxJXw7DDjMWTJTA

//pragma protect end_data_block
//pragma protect digest_block
44vlFi/szdc7vB1/iVy6765yeJs=
//pragma protect end_digest_block
//pragma protect end_protected
