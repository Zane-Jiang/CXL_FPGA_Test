// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m0Ao0IYn/PUcg3zeyNXga1iHZpqxe8woSYbhjU5iKymRQBiw628xjVGEDjRc
AN2W349tDE4/m+DjnWpF0lyfj0BTIQyfFTt4GwZzOaQpMloUHflBZcGUk0m3
gAKv9KTPQwn7cc7hMU2USoKmEMfAiClHe6jSCRW4t1ZiEkEmWe8qw8JRV+FY
I7VXGyEn3hXFZrvuFcszozYz6dV8zlak/eYvuffA0tDQq6rV0NLOhkGQIPLw
iDmWMtMFQfDJK//sf3BKPVI+nAMs55VI/PRfCOYOL7KxokHlGHeII8HYNr4x
+eyL8h8A32aWoZKS2iX6X8TN7INBNc+YH9/+SwEybw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CmsKAYwQnQgviotSGIUOVkNGDR+5vySFYkMCzbxdexR9EOw2fFdBU/PF/6AD
YKVWxSMSJ47qgyQtw0AgZTrPmi66DTraSZK9m7MahinsXX/dJUDZkA+tQJIG
n03YQ7klls8Si4mhrSJWSIy3tE4VZj8GjmezWK2HCdF+b12TP5Ep3tQNHq+O
EqHw/zoq0Fk+03KOSRtJ2BQxvLrYvETe8jJlh7UjTJeH3uk7WoWbSsWaQEh2
m80YYpRN/tb2bZ1kw51DYjhNU264LOrczvxJjToRRP2Z6X77E7nMsCLLEmVr
KfPGSe79wa5tYktEu+PCRTzO6Q7s3NBlDhOI9vIOoQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pvvTApD1BCg6pZ+zBKTAE7xtKjDsoJJx62crJDe0DQUF597/7d2d2UDJ5NeJ
iED43dm4MSBJL3lOGBebA8LTcq+QxakU/nESNDKgclHWqqenHaNw4LNcVSxs
zbtWHyiBgKAa0oGYZ73xA+RFwdnK/gmKk633KopzByKoWkPpWi6Ktre0ybBY
Q61bXiYBGBdlwuHfntMbQwGCt7vqA2qnW9r+6TfZe5e7uFs5f0kPyCw1HKIZ
0G3BMWR7/akY8zCQ6mYxsZHMn+54x6Gupbknh2tQCrXRl0d4JJxKggCX0Wjj
zBAvsiei3SpkAnfL8Htc0B1EjUc7uX2UvggeHl6kQQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ihbtZLrZ77NmVavaDRLaD2+7/tsPu0a9UYTJY+u8LlixSlcBWqRv/1Mq0/Ik
Tlp44NFgAcuPZDDbKjL4QHyF8h/Yl84RoqV2ZXdK++mFh9RmVfVlyoiBU8tg
/nb3lkTO+61GKI29fwIedrAyKiQz/3e+kHFsvb8B5dy9CLxwS2M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rWQ1/8Qoc7KZLHuDcfnGjXphYGA/Y7L75pWq7pKzHDAfa5c4aCQ5vlp/J3v+
HbMHC7Hm1pDuIk+B2iKWkoHI0VWSlM6dFETqidEmUOjyWC2yi7+7elAkRbUV
+eypSs0h/lN9qCxOJSeQWLWqsQ8Ngr2WXL0e6ncWbi0Bz9wHPS0/tMij5wgi
8fuCO0s0QRvIdV70++X+RR8h2cJK1Blx381R3w+pojvAdUqHkdx2AGLmu7nW
rGUL6g5eqSBuZR1U68pQv/vcmJzknOhpWkN9A+asTsVz/oU18m7NWg+baUul
+JKr3tAs33v/urtb1ZUw1KN9q2oY7A0aboLEo1fCBdUELhTkDTe+E1RInIcb
VbgjbyEz025sc7QP2szn4/ZNU/SLLmz4ZZHwyXloygDfzynw2XaX9IMdF9gY
V4j+EpynaG3a7/ip5oNLXguN2uucHPgG6H+YXjOkEl2ZH3Jvpiy7Rq9DJG5H
2+e7CRV1sq2QQcQ6cjJIBgI/Le0HSNBq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dBuXc/NhprQNa+LmeZXRP9CQ7EDo6xl/5sSYl/YqFLz/uuApEe2YQRRLY3T/
nj/uGI+EzXhMw+EiZyW2xHplJLO5nJJjFxXl1jOlwbVuLhhIk8JqhT63Svcv
B9BRApPzCkprHP9pYCmkawwdV7k7Wdf4Kx9iXsXCi4a34ahL82U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KBD0snsuvZOFFJPnAPN0ji6QEmGWCJqv7YHq6SCzgB3mzF7yBm2xMOvOfosR
KMyWg+YiEdM1UCZBgemtv0u+6WRwzEFmKY38zz88XTogfZt2UfL/yul8hCN+
H+JW6TyOhWF7je9GaKuDB2VrQfsFuU/AINSRt373au+tQ8mtukI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 44048)
`pragma protect data_block
EClybOFhO4/6UV3e+SpcM1mUOgwecbP1sfI8pXhE6qeAgUCKP5VjM1DvvSd7
RqBf4nP3So6l7Ush1QiH6Es6XXBSl1Kx/+oMrV2oatKMsU/hHi6pVsCowZf2
uRXNpANib5Vg7PbkUR4EkUdRT1T/eW/SbdHfEim5NHRcwPs7uI/HrlKy5TB8
/BueYBYB8M1OlnFGcWKKEl7Iki8grYI2pM/t5v2/+/DIjnTuVjqy7+Iog7Z3
ue94BAs6+mtQoNQQvOdjCzhEgo3As/1D32AHyE1sJe4awVEIlRmRm9mHqPfF
sb0rKbprlOSNM2Er/2EswPqj/2//HT4FUfnbralTaY3AkpWjhv8nxQXs38uc
XHlTUb9mKDzSu9ndxOPfVeAjEOga3LifIqNkRHTnCLgIaE0k6+1k5AU6OeNk
85WxduOq1ufctwLreGP6H1ETtjlAAv619NRPg6YlRi324UtIqQX7QcMtFcbE
aBg7x+Vuq8vJbCtTOx4MWhjkWst6JH8sF7wXOxAIoOVqhRmzmrVMtZVpnfKY
OMtibeFbWXJSyLZ8vt8q+sfL8SzzChCY0HHDItUEp3IJy5HfgaG6Kcre/sag
8cgqAhNm/UnY/GAeL5wqyoMf880scTdIIn22OPSUYVufiah5jABFrSS/Mrim
Hqap0GTJrW2+oiaJGmND1FM0AZGNBS+nCeDbr3F1i3TfIqtuxb7huFZe1+3C
DpwXDQEBvFqkzzx6eE+nWiC0/1V4i/Lo4xdeANVHF1WGqZRfCcJ4xVO4gtI4
Lw+XLHdocYykRgnAVijgLkUKFnLj+0oErqE73rPCnsjVDA1h83SaS6eW6Jvk
BYfNz4KgEQAS6iKXTGqhh1ShUNWPNL1HQ6M+RWh739pNHgcWd7zRMcIiyxbI
rT9Jsi7Wssk6M1jsAqnMTZdD062OnQZNuLxfFLbqbHSt5ir7cCoCIXQ7QucC
/vVxwSSwhzUDBeSvcl6nlDoCRU7JkMsYcT27XPHDqFmHMQtdOTpk2w46ICZI
Q5Hwhm1Pe/GJBOYVj+/84sD9yOq8hjMMUMD/9JzhQ0/l5xtY4SjlhL/fP7Ct
jWpvNyOuSBDoE0piEQ/v07BFHOL3aw8ake3tUP0nquwUJudexnxtZ7RjwNOS
u4glQ+j/oreCk2jyu3IEPw1faq5c/t+vxCK9ghdM+BrW4g2wyZTpcSzsEufz
yvMpJmoLvXYq1rxTLQjgmfwnlrqJluYiH8cc78Nyr3Qi0h0p1E/ZiGIw0Pwa
nkL3JtP23o/vVzOkcrJCTanFASWkmMf+35gP8NXdanES61c80ebno7qrpulE
d/wwyk5KOn17HyuI9NVcPgco1YFYFGj2OS+hGzia3ugsqVvok7Fn2POMMZs4
0KwSozrMYpnr5hBmKU3gYjW+c+OE+K7iN7kVAJ2fU7mj5P91W0JTC1pOtVQT
l2qHomsi3gYsAeggfKrecJw8qoQYhXzK4A/GaImbpvK+MvQse9DNqWue4iM5
ID60q9yVD5RHzcvUSuHZ6zaS1a+SkyobL9Zxq2TPxUWmTURVJ7nxzQ08JJOp
oRSL5Davbf7lyH+MqJMrkhN+FuK4GBppwU9DMABi13xURs3JsR/3A08ySCw1
WrqZEX54AgAnvkHh0gAqJLFI/Xauxw48n8b01IxOCXvsXcNBOWUZ+4SaUIQF
iI+lmDk05PCsjI9IR/a2IRaYn98BxgJ3DHjhkO5to64BkvGnPAm77XDAAkNQ
Pf4BdmvySkznaj83OzqOVA+O7houpDccbh4Po+k7HU3nQ55YlERvp2H3kAeW
qus5NCznmXQKhCx8N5jw7KHLcjwBvHW9wuHq8Ua7uvUQTRaBzeUa/ZJ9XIWi
9BgqSMuSSQWzFuSgMdSUAtuKGAnbgDiXRlhaoo9xb41/Qs++5BxLR71z8MwP
vXBVV5QS4PORTvtc3GbrIQdW6ZDTJkGpRHUavIsVll+dAXKqH2OaXt8g4qro
zRXrtTEsZl3Gf4p1vHLHgNcMwebNtt+WYEmfnZvLF4udZ0iz2g9CfpO8A3Yj
ce6PVnlv6yrBdz3EdUdDQirgSire40b3H6JyRqgwZjvzB3u8t9/9kresL0gq
lBR2dV7MtHq2vhyLpswhA+qJWmiGWKdWYuh9YBJQOJlyGDCUn55+ASlTZaAR
bX/QVJOTrU2tT2xGn2iwap3MPQoyriRCWclfVUAOH6/WkiGh+aKlzDDnlT3E
ZFRk39n4mLEEl5qyhLHbr9rSzPHycTV8fDB8J1zf0qlf/fwVy4Iah7ZYRlqU
8eg8xGI4qXYFqSYQ/JRbA844fRrCE2qjxRlk1wetT4qGKv+v4HAeO4SVfBkg
BfDjENpJ4nuarefsyTNQXwdAtIFxH3FkG+jbVoTuGwKU2hzM3Aisk8zBi2Nu
x/pVi3DFXqsldlvGUzWHVkEjkgJTtiePB6W7Yhn6fjoup9fRJFiCgKVAQJW3
VLkoLz1SRSiVHw8ni+yW/ckHAwpqXQp3N9gvKJjVfnvyHTm47YFrLltpva5K
KkBdLZ4nu86EkHQYKCwQSNib/t5IxaToouKeLrecbwZQMMX5JyQuk/8ZgSku
sColWODCE5FQm87hNgMPWpfc31jSjWzxVdpfKg1m9q0d3JkYWOYuWJp7ejd/
Ze5+fupc+5/e9qv8vlASheJg+WZxmXAXLwdcVz/RDuVeX/7oqe469VUWCPHi
jvSwDWlcnoy6h2DShOx5K9Lb8jUXiEJMKs0g2YUio8gq4ZoZa7S3ymDTmXfE
piUsEjyaGZ+4XwR3G1AmN+GOTOPLgFRU5h530Q5IN34bKWiwAbIOMWFxSmmu
GMzVV/ihNzPnNEJgzoIQJL5wh2S/GfqvUFsTCKysvhmVaK+YZUDnwoEtZ1d6
6Z0GH4MGNjkutqJ4ZGFpm4z3qR7A4pz0pHxWEDrI0Syaof3ZDA2Y2QRIfJxP
9mUNarvPaicZ7xLUfGhJD/oWMdzFpuTJZlU9/RSxsrdeSKivfs6RlbrgItgb
xlTcmjZiPUDRR6KUrn4apcHE1jgdH8Y92OyS44QNma1K1EpBs6jteN9vjkF4
+PvBmZFl54rwl+0CjdfiLq/l8Np938/pD0wrUMdNdaZ1VgEPdtcNp0hDhOPZ
ikN207GRFdqqQZ0crfVjdhZWpzHmwM2XJpbbH76/JgxWbTaRBVZypk0Wor4q
AjxMUQJ+qwcz/Flc95MTOELbTNbc4qbaTR+FT5lRY3O9d6Go/1JVHeYYmCma
5YNZgC59YNN+oNxSTBsrQnC0YMIxL3YXHj7EZDCjC1GwxnhIgbQ5ajoIfbFJ
AtHTTijRA/2PO8vbTcJd+uww7Gz2jwA3vY6c3fVCT77g6BA3pylhPOy9qRtd
eLdS46lpIFWKakDrW+jxC17P7iFakYjj1viKFcECZz1phsFvuvA3L8LuLRJv
uuFmaHz6Ixxqa7RhC49x3D8ALIHFbHuqJ5dXUKoOJ9+eUC2ZpQEuw5TWGnSR
DLBvUC09igeaMf/VKwTT9wLXrHIKEuHy/hOjXLubq/bAkQESOUnoh8BA/Dnu
J9J1Px5yv/qKVgvuc1EuZ90xx9v/mxcPCy6W+DTh2dtLx1FpEjGiygMNwPIz
5OrVQtd2l4YGZw6vkDn+IBk59tfOizf+SCW07H1wEB0ejMtdzQFJ/xT0E2tg
rnwHJFVqBKqBB5EA8AvDNYb+kWx9w4ERi6Xr4LtzzFfGYYprbcA38Y//94xV
T6gSMkQtzXqmOXbNbp9Ap7MAEww4QWhxa+RkWekKZcSvkaafbmHd4B3AW4hC
oKQI5xR0sxmdxBjopZBxip8e75sPyWDsZlGkq47Abxa9F+ys2PzgWbUVe0++
3FU5MU7FJoTivDf9Hn9LqsJV+9z82xP8YL0+te6g35cD/OKtz25rhXcy6U7p
Uh9hgME6zcEtIYi95iWgSLv01JTRdC47uJ5GGvjd3XQr64OzHdThKj3spSEi
4emlbs3f1rw4oTqayDB5TGq+QglkzN4subTGEzdRzyYAaFlxFwAPTg1A5G0G
TExwYo5xGfjOBTmUwcfktQK2TNIQIbcTyZL1+Ds0UsncP8Amv+40i7RZU0rM
dozxOZtvfe4P/QaCXNov4pCeqtmfWUv6c4+m5Jc2iPtmL4aV3ucNFYVtyUDG
fXA64AVMmCcL9EstXcgR81WfvRMEEux+4XLovq8fDWcz6D/fHKnHlAZbdr7Q
YKZoi/S+HpTqvcPX/NyUTRDjvl1SHHteM6oK3kWpaUYTet37pMM8eTe+Mny4
WvL0n3CKJ5a674j6ffSw2X1jq3l7ji32rsCMsub9FYhv9Hn6H+oNR0BTLX/3
kyA/UMQNpsc12M3aRvCFqyaX6pe94mPC94uzYyn+L1o+xMrQYgyuf+045c0J
fs6VF2elLLCnD/EPnKBpa24vV3UaAX+Ywhq8lV2IiRNWfOXRQOcIlmIqjUuy
sKxhHvbSdVSbPQivIDaYZxmdTSMdiJyTO+J1ZXgxeDJWjbSkABlyMyNZmsny
9YS82lNa9rVeD1rqp6AG/dt3gcV5Daj53mWFdQwEppPRIJPi1Cp4ATQVjxeL
cBz1xVfEOV7m4c+7AfQ3gqkIj92TmOk4+7fSnS39GKzlpHp1RV48uwtvBSoO
c/zWsaFKQLth7JewEdn5WJto3tX70fC5SlTJTnLdbVJ01dAfEOM+SdWF+MIs
MVVlXciEeCON86a4Gdg0BUpslfkyWGAtHbCc20KZpIGnCudUp7fchr4aGzJG
U4GBgcrF1UDkZwTbyiGhFglN2UiBBDNyShIjzerX/YotPzlOziw5Jb0e8c5g
m7rg95tigr7q3v1BP3v6xdynlitdNHl9BMQ2XWEOeUXm8o4U6Q0GhF+iBW/C
jlwvK0KcZ/TKVv30TCw6xMhxf924HDpOpj2/BzrmjdLaihfAVECVjpIFlNTF
zri75+gtw7kZTRhvdX/oZVZSB5OLzilYujrUKsCFTiM1FH/BqwCaIEbtxzWw
NCAmI03v17ZNLZkuPITNysueiQdRlkrz+P0ga0zfc489PlIxgDlhyI7XCrsT
W0SfN8bbFUC1/rDftjhNYDumnMqyLBhO2YPfV6AqHGAXoW/uB8dzIhL73BHz
NuK/WGOIkCI0dqbWu8NWXQZX0wiFEK2JqZEoVGWk2nKJNJp4bI3QNK15xJUk
vCJ5f7ixzNmb6QsZOTphIll9j6Ip+i5PDqRHF8LHm0qurL2vGZylG3gkqWwY
zahnCivtf4c3LWlEGw9IklB4KkINTwiN+mSfZ/a3f+hO8Ds/5+SAY+YMJMYV
74pp4CLZyO2UV3/zBWLey+mIpsNnm3/uqfHr27eV343GslJuEOcAfBO24DiX
qxHPqKMoIuPy6G5hR85lWAuigx7c9quw9U1gF9gsunY5r1Iu6qRuhh0du59w
fNPU4MTSxn/wGfw6yO6yK6eDNNKNBIeJqjrlLQeBJVovGDGeLdSXHT9mWlvd
VYGM1V7Hm2Fk7ejbNRlNeHtlVhCwYWesC6tYQhL0OesEKTKYh1D7qu5guxdN
jxZKIx2TPUwOppRi+jfjpXe4DJ7yTD9RNu71F/NLIrMpx8IdM0aIaLOayloR
oFwgN6LxMssY56P1sV6o9aF0FUS8DPoxTFxYgbD4lvf4YvIx01RcEaey3a0z
B7S3iXnX49JLs/V90mgAljUPjAepyAyB0IDka5LqQA63QWc67JjPp/uq63ii
WyLMKeRpQobHo7ibngQn81CuXhDdnSdhdouUtpR9quSCiXloP5WWlAxUiLbm
YC8fDGG8n+j4ZEPdcWUUbiIYYdK+3lqUlJOOevKKNGDNb61my5g0ztgme0OO
gY9hnvIdIdcFhavwi+3MY2HD0S3DxpTIJZf9WhWZYLC1amzAUqHXbMnhDbRB
NdHzVkAXOtv9yTDvy88q2LbH8TVL66VvvNr5ai+O5+dXBbT1Wd0K5OWvmE47
58MTSWGfxnKnWCfaEUVdCOM98RjHakvBu0ohYXpXHfVke/T+PtLsdIGM+mxn
ZkKX3OGArNV2iZwMdjr0hnNKlXUSrKJq1r+kmOrR/HovmYdTv1TZv8oVKgic
CilkUtMPYzt3YAPeVFbXKUmCPFC1lcQEFSu8YCaZAGWAhzTX6sxBxcn5/+0C
BTud+aiARaNWDRsxVjbkrqY8LcOCK7gDWisH0Dk09OdvtCmwGWN4xARWZb+Z
baYOZCQsFMnzzqrb6owzJNr06WzjXY2qjdua0K5278rgMUrftoL9liAnEQX3
SGA6oWdpxYMz643uIMe2QgLYfwiaTDfARUU7BCNraXxTNlfWWU040j7b4NL6
45wKzRzvDwm2wOloJ9tvKErSw0Qh2hYx1ojGHkgHZySAA4PFqE+U1FjWopmq
iH5aJvZWsfFFZfPk5oq9WT1dRHr4gGYUxOIOl2bQrESlwRzEpW2tD+Ur+HyL
GSWB3x1oq9DbHOh7HJ/LBZupGaQGXzYUD5LZ3dbG9yiR33PYUnWvELJQLwIM
U2dW4y8O+IfF6EjN+KYW61S9O40JSX5Q77uOMbPr8SsaHX8DYG8c1jaodzRd
QwCyNxVcZqdmDmpTcYqZittgjt+exduRCqVg0g+vWZSuSD0HDk6bVflK+aYZ
FVBKDoEwQ/5EMSNv3bCToBH+YUQOdfGfz9cCNT2Gs4p52U6teN526RbATfyW
/Dtk7GVgsg2YEjjqCsmNH8CNN6JLhuk97ViHcd+dcKDZuPLpNGKoDXfEPkj3
yVCsYccBb0JDyUfLYAnvSA+f1413JVU2FGGca5zKdofOP7FReszQAx3lyNrM
YfWqUqgZG9T8xm+tPgoteg99mwwfhEXlvYPTTHaNpyo/wXIm2TAP/HXaLPPB
3Iek9L7MORlcFcIzZiC+PoMItmTez/ep5gnANhjwx+1KKsdeWPNnxJCeG0n6
bHoY9DdvbysIIXow38kVcJMl5sLSss697bQLS1ug0O0i1Q0a41V573sx7zDT
OiwBBM3u64drzIc9OwBIuEWGULSq52gwF75Z/13xQ7ynR9q8pJhDhvHq1x/Q
58SgYfdO3oxxXJ9aj5pwceyvfEimwRrHujsMS12R5Qy2Fqe5sd1hNtd4/H2t
9bF112tPAH/oWntGsYNjhilpUz74M+O+S6N2k4y5pIP6DZtcWY7z75ChN0XJ
inB+w1d1UJAtw3P8rmz7BIQmt3hyJBj/fXyAWQ+Bx03e1gsrYIWSNZW17GSS
mGAXp8dhVw3qGgnPM9O0iEGO7poWMU2+Z0+seDmN6NQIolLX+IcXs9F5o0P4
VMWIjFge2jB+HWGHQAxDRKJsiLc5CRGjEqL/0+CX7gSt0jWkQ2eQraE6x0Qz
xvcRiN2qT2mBkeS0BJ+370ROeAi9Bas87Z+38TNizmrINBYINlVdgAueqIeW
K6kUKFOkZDsDr/TN5rsSDxWx25AaXt1xNi3QVrcc+5pc3zlFulmM47jHQMjV
bQagiq2KXBBNBY+eob8MITdsHz1H2K/+j3h43to89zbxKw/cfiFWIiH9TjJ+
1UtnBtxCAUCUmrmte1ty95l2u0P2RqY7Io6JBB9OK3GT706duDf9tyrim0i6
q/sOEMdYZjU2sbYe6zw3yj7vRUQ+Dqdq/p5se/KxHQcw32mSan6O3Besd1LZ
YNoIGQCgfaXUadNco/WKmNUZ29j3d85Y2lOXoMoNUboZxD0crS/scB7fD5Sr
KGelrVh0j2qXlKzow7kodo5Gl+RJlDoHtYTPcE0vcpaAbqDbsnvgQXa2A7OW
/3K12EqXEMGRJphtQNNhFFi2KOFO8kGzmyqGwF8hlKuzCU0qZtexzu9ikMFU
q8DI/1xh027jzZrImK6eM2WWVus7PDJpsWAXGCyjmJexAF8Q1hprtrwFu7f0
iDVNn81OHjDpg12N32uImXMhobOYNGfAafC2vqkXKV7Csz+uk/K8ki7MCrVS
dnYIYkHE4chzBLxQudZWeD6v60RaVtGa3LjukIeS99kirEEyE4gIaN46fOuA
8KP7RQDE7c+pyu3xHw5LwY3aJvYqFszZbSn5D2O0i4GCNyQUYqqmPV3EmAG3
niD3bjZid3e8ZLjAEfzVBpH8sGqSxD/vSjCDo2kosblYoJ8WSZKAW7qN9CtD
rsmfNCKmSAa++DpVC58iyYhfAqAlUyjlvbjhSZ6+JAhnGSsle2hKvduMcaD2
VhbV1CakijLf7AE9ogquvTOF3CB2EsrmWZbJQUIeyhdGRkhPZhco4QrOkFtR
SKMqFDqtndCBZUXJ2J60G+LXsonqA7ITyRxlH4vaXQgkm92GsiHimZSHpVHu
V37i/5/055Y3i7Arymcr6F2DSIs05LgHuqiDhH5X+4xmWvJoyyYUBd9c9Zee
i609Ix/snwYq5N0hN5KMgVu5J29qRGXkGr9W/GP1Vf3C+mqS7yLFjOaNxqwe
2kh5Wzsfnfs88YdxQpnSid2v8KzpLziM33/RoOj9pL8cqwxPMJZz6sKeRyBS
O2dp73iqagm+oHJzHIOzCYhDJMvUWqxb69GyKpCh4ksL70BiGbNcCGEWSmOY
O4il7NN86ZNEqVSjDHNRW85wfjYPyDtqcWjCsCMy5BTIh7lMS8u4+aH9B3ZT
efv9pjopHpIwSClCDiln9QEo0MzJK1zO54rtUkq56ny/+pwQYY+ndgrRA/aj
NlSp9+peuTTE37LhX0R4ngmcmobhbNG/+MbLHX7dUYHtHhmIwdC0M4wlnSqQ
GRRDu+HqWwGZgxvk50u8nKVr6hGF+N6/XJu6RWmr2rjo8h3gsLxSo8M/YAqA
FyPPKW047yhKWPaYNKXcu2Q3j1m+dnr5fX0MffG1eYdamjipynTnEW9ikBZZ
uxPNxjeXxnI8L1WrKky+swbleawEAJqEpZvCAAYPtRRz6dXVgZhpARkmxn0k
RoPHH39e46wfANw7ieqpM3QocCNx0KexftbzqdWZylRR8LsNScO6Is/GdNRm
v5m84UMUelrGyQZAUJw9teCVaAUM70OGtlw/boxqQ54Am97hZFEKTwbuKb8w
dPjb5WLvzK5PUMsXTuL6nqHrXlbkgpAJab95MBFrJLaP2tlQojp/J6VHs96C
FHgjnC8CWLSPj949UC228QEXIdN2o1TB8xzfJWP5K+L8qIyYFBRFhOkZe2Do
0RKJ+WUg45LTIiVd84qGl1NpMFN0L2O2XRtBKH5FEIc3Ae+DCBBwOtT/alja
OEcR/pTJP7sNI/4297BMItxhGf4h4/hIi/Sspu35wLjiPwSRu9/55NK2Iqfi
wVzGYZp+wUiLOugtumr8BmdU5sTvLuMRO4Md3uc3MCKJOcTh+8/mPQYL6ZmZ
tXFGdbU7L9cOonTuKPJNFQcu30wplToRPpWNhkhp5kaAmHtshTs3G/JIeHWL
vRFKTlDBVXFyoMumPh0krpYOkb9x96fjNANQK6StNt3GdKiO+WWOsLr7IwcE
dynde7bIy+Z3q9vAEuI5ljFJFdpEUCLfQtpCIdEVgAP9XMo2gyw/cRKjqjP4
FCap+AFGgvnM3jqG3EpqQoKfG5/IPsFznuJh7y4Ol46ABLO11iVUw6QXG1ch
BayvnkfIdPTtjfKQtz6ONVHBhvuGXr+p3BkETJbqWM1wexMsij4VAe5ulgnT
csoB6TCGPnmjiPjjfYYNT6CZS8K2WrTpJhVu4XiSzL9CYbZfBjyRK1PUDPPP
mCRbS/V3AZ1rdUbSarqb+EKhLQYNZ7uuVCMbDJpTRXOz9es9Wh4owM2Bqi+8
R/IyKtmTkWsq268ZnbjhezctnV4Ai9qs3LmMffJc+UbmhoKEdp9DtKAGUjkC
1u2OSpx2oa/XoiVAqfulJ4V42VA14Osz++IF8JCnL91BED5FfOzw5mhad+zM
5Cs9xHBnCORg93LnpEyl8hQzfXn7V16ulGk2iGVlT3nWf1Rxax2zasbfft8J
5XfBJdlk1jFyYpkU0JAKxnf6io3V3rZlgin6WnnyA5LU2uuaXPP0j9FSMOLu
ahrd7BMyLwqKDQId/kc/e99CdRgcaaHiXqwN0KoQWOQmfCfsHoAb8T/Qyhod
as56yuxeTw4NX3XL2jRaTgmNAwlXQQ8kiM36/8st0tzeIDzp+9JitWblb+My
AR/OsUo6Yiz3DClptmS3kwZKfGh4ExaqcRlesp+/qsyBU8QFL9oP6NjHHcta
KauLS0pgzG/MHgS3FBtFVnx689B4vBnPJEK+lH+YqYCyG+pyfuoCuCXBh5CH
xCPFjOwlpqtCSJeJN6XXljLMwFxr3Xp71UU2gJOEtlAYWbSsJRGN+KQZtMre
jgvVw9KfywIXAYCcxcKnfFcnHUmU0hGq3299r/5p6+0sxx9cEtVHJKLstFrU
5elgvQBif3SV5jEfiMWVMnOZT5jGHkxpypflLIBuoKWO9jCFPqlJ/qfAj8MZ
m4ds8517JNS6mRYHTX8ae2fitDCEz3+I3hiGURYZBYcDGwa7j+EwRe6krw1r
LAFUqDZ5XOxhaDFFe9CLsFz/BDl0P3b/kbBgEh/Y62RXUHTGe8TYxbPDByOU
A3oj6ULU5kuSQkFlmzd11tN/ieZv18V/ji+HH1WQhUAkhvHImbt0wMcyR8p9
yPPW56zZ3q7uWR8nWHerqc62n5D0NUesFqds4U1x4kUs4cUo2OI9kIID+iWu
xfbOvqhQG5nSSThjFS65Zo/9NeTU7bPQnnJYPJX8O8jx4wITIPpTywnunmez
Xbs44Yoy8RJ3EBYl93G/PeQAX+xZBJ3zjKeQTWTxZ7qHGXR6iepBXbsSkMPF
r3PvPHeLu9YgQatwKVhpi54Q9pD6pGo6y95zEYH9m/QTQFXoUlYFWpfL0qIU
jI3gTfMtfiAv2zVX0ofBUGfWZ3L+8yOCsp6GUfAeozWKmannwBBMXW2Hki9M
2y7X7I8yaU3ItMaM8Pd+erABsWgsscloW8gOlLhkz2WdxFOffVLx6x/Xugnp
uPzbiPkAyi+xQ2z+K5jlXaQLyVSw6vvlynvsADRd2pFDpbpJOQ2wI/asxaSs
Wo3zXUFhvppRRNs1oovLhL0IF61Kd4sWXd4TVbhi52KpPBwHnz2ZEMpaJrnd
tKTb+9Xuem7hHMhLju2UBeXCZMuOI/c8LC8qa/v2Kn4W1Wq3LOixOmBVJb8T
vSQGk6bcabVO5r+lkcErKaiUtFrMkk0VJhb8g2JtIS3nNWRC9UWhQOLoDqNo
cGeSAQ/YNqsOJvCwiHA9XRl8YJErQv1JNKNQuAv+69yNfB6XB0WzGHBxgTuE
ZBl6+J2qld8KP1rf4swOL8KHogTszCfBltGDuN9J3DuvwZ5mRBgNioVHO0W6
leChRwdXzhti2aIpLYBQh7dJeOJUwlP/s1vFw0/x235u8LMQYQP0fsj5YdvL
jsYuMJgn7tpljIOVc38QmDq3nGN3cvL+cvnN9gWN4DgzHrilhHtHjv1HH/t4
2z1t6yyPJJvc8SeQixr19aB1Va/e9TG47nkr3GzukjfPimQhuNBMIzkwrMMc
Dn0qBI5whAFuvIwPPibIVkDN+l7PqcJEDyT/kqRO5UJL0JEIFkDsp3+F582S
VwpIrC9k9M9S/69kij9X2VYEUA+4ia2eOU73f22OA9y2Yk48P2kAo1QpZ4Xv
mSJGgx8rDkuqbHN5B2vc3CMnPI7zZM8yNA/ipSpiH7RyIaAtqhHtZizGrdqO
yWb+AggXj1eXUCL/UAuKE1JDpE5Etn/tSfNSO9mYbMxeEKkMW0PIOH8IidTh
pVYv8DCqW/68FC3BlaU/AWscNQI/4xbUnNbsyJ3SQimpjGDfRRFiPeUjlaAG
KjbgO4wxqTVLfRaaSyNEwlnhSHtrypovqtyqMz+0HW4yzdm3AnfObOFZreKH
o820lNBdAgEYmEe9QAJ6sEXMWZtK5dcoZq89GLXBRvmqNNruaakE//VJdZOD
az2tIH0FuSownL3l3//VIiWAQ61VH6mYNNZUpTgOA/IEYu0l57/qmfKhGWXB
8j9Mof+RnMH96OFDdBVXvFvAP86WAs2wZTffNlhOL13CYzPwQrqlnQPEX2F1
Mpq8a0b6bjkvT8OBw4CXNZt+wD728KM2iL8aLMc88glDx1hm28x/tHH0WCSs
gAlJ78Jfa8TTghSIcwvev7DWWTk3lQE8nLYfPa1W5sRJLZmCk/ClFgsbg00n
hSI50qWe1+cmsm4KDU5GB41J++CpQzTl7voB4g0LU1jjGOz+S5bGww2NlSvC
cKtvq6yVAUDoCPEjwYgjSvMAxbwTBn213Pu7N/pL0BuRiVkp/pOFKLYitBC8
13gvAJWTaIH/Y/2LFG0pqp4kUANi9swJGeHaVU7Xgehu6tAwmveTT1vvxtCE
ZJzt3VZFbfUlIBNg//itHKd6rOTdcJBo8ysW9oMYo8FP/Rhaa40SlQlHSJgC
yXApGVW9LnSQvhw1DOv8dY/doJFrp69VKs9AweBuSc8BH0GstvrUVhVj2LlO
ERrjno3kjRvtv1IZr4YYZwjBwiI7dRr0p+LMU8/q2IsNtB2E8xHlTMqFaxmU
NZxa/iaAGskB5pzOp12NpTQumdVMiovFpN+GDyB4AMmSFWwCRj7R+8B7SOQf
0g7Dy3zh8KLxQotHN53Wr3+Nt6u2yRXMBHbB4kO+9XH2EU7ORdDKf9uGC/uj
0jTMjap11WLupwEUCV4IUIdpK4uN8Zy/TxVw4AplbdVRvtm1MxSa/EOkdYk9
7FYgNXcccNZPWyLdcrZG3loyu5+1az4m2wDTQFt7Z+w10WXnGbkIpK4qkvxx
FoYpp7GNsAnXA+fEjAj8qiBd0Ra+PlbPHXLYf8mISl8WjFIIxk99McWbKzDH
9XPoALMFU0vVI1S9BpbHHlSnc7SgohkkfdeLqPzEMgqPybkxAUpSzgsEcK4c
UBrpEQwIIL3t2anqLjTER8C0dmlAq130N5+KucusN98a4h81g9OxHwL1/RAl
8i3mASyIh0fFGbvzOTzgYfQP9LRMyBAzGhg4LSEY8ss7/pcOl8QJHdEaGfYz
iOIttHI+P5fBVopp15danzjbmdGJYU0oAmvUdQpV24e1FOtwGVudS54TSxaO
aCD7d9ORe9pLd+BurpNG0fH9nFGNhhnHEMdGwH+65MhqhPbz72OUzsjHntSG
4sh0TZYkna1/in7U+FtrHGPlcUWFsiCUI926QZClOwgxV+otifSpEFTbZlHK
8FTK3hVh/fZRWi8KG7zT6PJFhcPryRPZWaOr3FKUoCCX1AOtZ8lZhV5TCTFr
K5Xm3vxzbO8h+qQWB++YyxiCkXOPeogsUO8jDnoy8ZEhjnVkfGnX5CaIUm76
OLR14osENAC5RqNPLs0IJPmzeMk8jAB8uBoxVbbF3WAxuLhiuW+Nd2f6U7CB
j54LtDzaKG/pPV9pXQLhZgL1ZMPu8Dbfjz9oA0c2yRyKAqJPR2o8Ppi58vlw
IXSWvI8f6vtYKszwih2P2vq5qp+sbesfdtEx/DfSaQeLbrX/OrkKfl7p/TDz
aTzXbLsOSK/y8KTl4ct+Ng3uJ/Hal/cN1n5XI99Bliu08G6Iba8ViS1/RDPl
bJmHaO8yK+F62pVg9TsNlthZcnXvJMePQMrlKyZeL5CxKMUWh65vsIIuPHJY
QbaaePK1BZEyIRgOQimLV97nCKVH/yzkF+2dxGAYgqJyWN7hxZ3vohCjniQc
QpwXB2cKFvFVV/vnuzsnnKKFCPcTm+ZnRILU90p575wUnpJnJLl7RhY07vqV
iWnjEvcne47Y/aw7GEVIH/tN2HCsw2b2lOZHVX1pq6rUCDOV7coYhBRjbeAD
KqTLor7xG2iFFCkjXagQtWz7tLDuNSN4xCPTmJXNsQzymC5LSydgNBjQuhBD
YZ69VoYqyVteqMo/AvlIvfzjvkHWVtlulcQCYvS53c0Kr7XurfYgV3ks+obn
NBTqmjkZhylHlrPt8Z7hWAqIYByhTP0ZdDrO4DLc/7hqnWWCUIwu9vSTmfmr
R+yjg+ZLCsZUPNbVjZm8p68Wl+2oL4ZIVsNCvGBw5oH1y4WR6qWph1VK200e
NIkwAcFkXbgX12DvJ7uAFb3PD78/V7Ma8OWiCljuI+cniWflqZaSZ1r/pk+K
dLZYZmxpZm1/gevO7NIAQ6m/aWDtEkm/CvAEBGKSbTj51xLE32Y3Cm7Hdk4h
YMaatV699QUiAey3hFC1uZU24BrlZMCsnX7q1kzScGQN+mRzdLuvlF1ix3xs
t8I4s4khyen0/9CxVUIHN7WN2uNZGQoFC9DITKmNWo73QJRXw894eZfq/nJF
s399N4FJ3Hz7YIFqfXahAyiAFWk9r8WTnu1OvN0yo+J5vSPDwL6tNmhcaOdC
W1mp5RiAhcM/dk2MTcjd4saa7WKufQfUugI9fRy4REwYkrPRN8O7f1aLzmhn
qJPoUv6sQ6pPJpyOVov4wsSprzUHOHAPF1SZglSV2lwBuj62LNVWVVuC/TIh
sb9porwj1AMqTu3axiYrLS0aB5GLILY8vwIbjK/OJt6vbzXm1o8cgMuJCOyK
VbE7j8z/uAyC/umQITXBy9viSf75tkqzxjt5n92+9DizcBbaujxnMWCmRcsY
zKsLkr3TagjRVJZEAyxW0ynIH99Jye97RQTwtu9GLdl+zPyQVc4ci9tOQ7MQ
5nAwuOMl5Kd9XyGqH8PcyhGCAwyeoIQMqOwz7IU/d9YT8tnhSmZK17GoXfAC
6gsFlyAMKhrdyFYFtYg/771Vxi+CNGvtMLs5jJcFiz0Byx7JaNFsqxxuHmXo
vEajQFR1qD5FnhPO71Z8gSfpFyhVdBxVuqBW7GSHn53vAhDau5A/2jCC8fSB
wd6dsBc3kYvjJuhqj9Mz+uaoYS0cnqGCwQn7eTL2w5c9XBUrTEVISgxYKB3g
k6aSyMmilHar6HynKveZk0YcxarJHBl3fw2ymR04IfcYugmN/8s1oLMnynbt
/O2TW1Dff34Pmx3889mVn35x8NlMm9eCNdu1lTwgQBi1649rAiHer2NPDwyb
hHwwEQIsitAfwykrvQrqBik/HdTvs6Bv4mApTQ7kkgxEzQ4kAF3Tx0CdwYjI
RhrMgrX7YSrB9koP6o/TK/7VoUkT0F2DZFhV48kHRGsDLNlwkr49nFBu6Tdi
KrszTzU3Qma4VbIBjJ9L21nIpVdAOXsNDuuF5dFDjM4QMP9FxaSG4IV/Ft9e
84xB9aVU8cjeY8pT9lBMhpovQwX36i6oDdLPVx/eDuXe8MnV1vDxma7qxVer
3In0caedP1X/foLU9WzBnOioGXgED2Uwj21zXt5pwrj0pucD6zuZ/FM0MVLm
AjrXaVIafYew52BPB4+0Mk486K2YPDfU2Rzh2fSzjOpMjVCDM+hwDRWFkr4m
b4GeDzK03NTscPkYMK5dQxJ9eYazER1egsECpMXp0gGqrcDfgnwUQssex8qu
vy0/u3ZoicLLND+55Zj3cgbuSOuBfrapSauG0ohYP8b6Xwn01usnf4q0y+OT
Z+3nxhu+af8elPywCoGe/C4XTUG0ZLQllH/DQJHuKTOVdhFKrgyK/X5DFtjv
FZxAMZ5SkXcxTpujTnWBkvvtw6psw9BrhP+U1UY1rCpoRPIV20QrKSpeFqQx
Fm3IeJNWGi3wPnC5DMDOliErpZ3MqoliVpTv53B3IFbfsPhwNVoQKZV6abg7
vKqle11GcQGI4OrOF8rzFZytjNpOVE/Juxo2ChOoT+MW/5pdjkHQjG25B1mo
J4MbDhQYcYAfco17hd5IsRsv/1tqChoSSqeRbVO+OFF4WKrj0V+TYssAH5vV
h7OtKkTKtuXl3Qm9NL4HMVO857tYOD0J89xkrusglAhNNP76vTeKlidB6XNf
SLXVJh9VJuFc9ZBeHJ5Ra37DGjSmUJPSkhB47MiJGCSnhOOILaZ2aSBQ6/fx
mPcHdG6O2jk2yI18ZHSEK870q/BGf/3plbril0fNIdkdpVPM9TjQ3LnNifsb
YoNwHVkZBqRkK90HgQkmR3dkcj7kG7FuHOnilCJ01LV31wfuHhsRtdcrjX3b
iJte2TbKhHfApEHvYicUx/XK2+YpQ3lEFgKXiayLLjUG83LOh4Z8XnTHbLf3
JjPkDdgAtr6X+Bceyx4g4s/nnLWYMt82t5DkTBRxYJ/Ccbj5jkjLErNhh9FW
vkbI14eK5tV/+GSu0Kig88JNBwAzuQC23XAkf/3I3JvBp7E/M6HDem/XGVxU
SL+lC6ktPtWJlc6DQ5XVoKYhj6aDyqzDWPDwcTaW4HZJpJk/3kJwAYECrHhr
tKGk4g8d41YNuk0JZ8p7qTQk3OOG6u7pNStIaQ2MXU0ryvjVpwmEsChqaFNP
w2yyHCxeCwZPCMEk/0UHy00kj5zWgPLtHCIP7cKDX1uOG86y6uCC86U21OfP
e9FQ9bUq4C7mR9zlq6wW+h3GuyvQxamcUlJXxQ4u4oSpfO6M4jRwFjZ7MXGo
5VO589Cex7oAq6Zpkjv0EsOb3ZhTCitIJTs2g0Xxozp5JyGZVubZm47MRxMd
I2T9damHDlFVLXmd4Xc+GXd3XM9fZp7n3Oz26Q5ulUilreTBrGnGqrzCfhfH
8pBZLKUcfhor2OR3AJ+Trvnhw1aGUeu8sg4a+/ghFCUCxGkbcVHxE9Mxzypd
ELKDA7mpp42Fbboc5UpFq0eIGh1dVwZ317cqYYyaQeNyQZ6Lh1BoTy6ic41b
9GydSVoUCYYkWRYAfBjfeV/GKh8TyrpG6BwxegkTqbBJ6jqTF0ftWFghX4k9
HybnXVelH/QRxIXtpXnBZ+bdqw6CXdD/AmaRntu/O3Vzy0NeTeJrAYm4Uopl
Fpjvf0WezLn1uyEJZ1Rpv1Wzkf6JAIEiRTEx6+d0see/JwyTpi/UlLWSsLAh
QqEdPriM1tDnEKsSH6CQze/fGVI01bp2wSLbravsCQpqudfUsTTrkHyoDcv2
5Kc7Ez5D4tBKwWN1KhplSO8vOtumrsQah9qNT/W1MDMieotoNXT3/aiIcZ8B
vhqZdZQN4gfanNbvQUILqKGprCmGEDbbNMrL8ESGeZnbfPW0TLasdkhCIaQB
Q5mI0GcMkVtQ9KDxddVluMPBwzg+WIZTUUDsHxVR0tSznypHeoYfy/1h1uMy
cHwV2U+YJVN56lBBqa5w2wIYNi9mmlf8FMtffS/8H24AJ8FmSt6ektwZamP/
PuOMlDpqQOjgnLUTKDxrrdgg8ZKNkOFm4QpIiuyt5mGq4T+qR7fj1VMv8/QC
kZMLyTGr5j/tF/cpyD5jUX1dnbzfaOn/9+Fq29/tQX6zGBZ8TPdlhTKLmZCf
Zc7Xc+/gStRn8lg4N8mdD+WxDqktFdjg32SBiAjjZjcCO4IHJAXS2USy5K7V
jstk+tkDplYJYfVj5WsfFpfBkKYhEUjjBG1GNaa+UK3cAbIRk36CfhSEXX10
glgpJ6rqnYfU572bjDRoWrELUF2jZmfCmjaOrLCBuLy6WtvUaqrH5eYstvjr
mqMW+4Wtx9LLXGTECePIPAu1QwRdamsmEoAp88T10zPmHsB3AWbqdw/9qnfG
TFJrEBMe80uOYplyYgcPJnXXBv/mNvc8/sVTZ0WrlFLNnKovTPdkXmYa+Mf9
LkASWaCwZ4kNdcGLFB0VKk401+PoCMxeUXGY0iUIN4U0DFMfNOsuGLfNRanw
LhR7Fgno+znLeM70bhoYlsu9wKXmn8czUQCNj6eVWQPg8HpN3X0pKW3DUJ/g
Ta52IITc+6HkQdKKm8qaYRa28dmjo9hI9lNlJJCGz8hv894/0h/YChnDl9z8
k76vZ0174NgpmukUJFtHT01S1PpmpHRXEn7BU1QAysYmKD8Vh8/QuBRBNM4u
QUSSJuRf+OdWGE83GfJOp1xnVgC0rLhaKXDz3DZzXRNsNMkBie9UwsUUdQNT
WYGOz+7JO4Kse1AA7FxpqqiWi8qQDH7LI7ot46qYERR/C6yzi2qgeu3anCqi
tjKJNLllbX+8JzfJdX8BliF5t+IIc1YV1UHtSaGJsR1NIiSPCvpYOf4CJtih
kmtBNge2fPGYF8oe7iwwRIpIeeXZS6+Cyblcm7AfNqhTPdaz+TFK1yPHqfaK
4LkBirxkkfV7AjI2pLACcylhJBXK+hJlm5K6ia7ex1GLLS90OgGmtxhGWi97
0ofn0YM7hubT+m6g1pK9erF8TBI2UNjan1Xh3PcnR0ZbGn+ocsOnHiwmuhjQ
f7ORWhrL/LsC4QGQ2DIYV0itB7R6qzObwyAgp5XE9FaJA9zXp69vOCTMRveO
SFJrPUCncYbP8pLSH5sjcLN1sfBKbeTx9mtpZq3Sjl591kXb8tQEP+Jr4ZuU
gWZupkW1NcOdjBldVC/nTrtFqhP45Tx8UZwMhAkCy5VUchrkLhOOu0pr7I+P
XkYibXw+QeewIEqSnOUCWQBSCGuH3IQ8Rz+V5hlnp2etpvNCHfQx+h1jInhz
gJg5/IsIifvmnZJNzHTZTT+NFDV7WQE1bGM9JznmtM67xGqlIPuRPOXEpOJA
m43RAoYx2CmH5ph/jlb5SssVu9CrDScUY3NbEFOarM6FpvWqQdPidiVZWyGn
nwH/PM1zmXdwJJMww4jZ+rAqvqB6vlKe+B1W3kYC9Y0mcJAfK6c5N9sq34iU
TJeYg1lOZY6UbVWti2D1obg+hsBWQZGaqq04uRkJBw9+r1p6ALMTwdBkJ/IU
mIExOcSgGgBxK5MUKJGo0UmOEJD6LjS8ZJcOVs1jQOJKRmvD8seczUWD8pSc
Nz/rp1jIL9Ayu6Z4bQSv8RRQXbMcXvmFmmTJjTg3CFTegSCZzjnZG38PGDEE
GTAQ3YWQgB000ucGXt3QK2QQhC8SGFGFMY8tNmpCccc9DidavfbgbVEaK4iH
oS5Qi8YvfWnZ4NpT1uve4rS6aadFmvhNbxoyYe1dFECKPJIx2HtOnaud00ck
YYQfzXCNgyzuV8HGN5sS5YUpdk3bh0qoaw3ilYOCXbhASkypffAy8BaUhgMV
nHAq2ROEheeCMzZv+wGRgGkf0ZsLMkZlHw/FKNsjzrvQrmWbBJevcFjiwNwG
tvXnvpIsWWUXdreGH83HgrYujfZgMEvNwxSSJIZFi3AIVcDCqwLbpHQapZqW
koCzCzNO3I86h5zzgwOehCQwCGO2yw2RUdoSWz524GMPdCJTrkFa5ox8y1jM
WRYz3U93OCrzxapXt0rCABFY9onhX5Y8rJk6pkYBLLOFdUPvgJAQ/Mn1XeQM
KOjCJAzJ7LlcVS9WX6y+PJgkiS8w6TCi6/OM+xw0yEXmTqVjYTUqigP7i90F
vRkQlACNgGp2IYb8O843Qjvehrh2YEd+XvYNhgniDbbT6M1aSOVOGZ15QDzW
zWhSIe99ijd4w5KaAwWx1fEk+l606D0+LU/pV9GUmBxsHyXtuJzun5csoYA0
uKacoD+KZkGp2uEAI0Lr0grYXQIF3894W6kevY5zEROtMEx4LtlHKYvZXzHZ
T/CO1Kaf61F1pBa/m3UiwmsVweymNrhF3pyYTnYW2TXy6U9vcrmt9RPcHPmZ
Zcx242zP4u3KqzqNoXR9U3i6/TzkkloJ2WVWtbQso/nT/Zon213Eo03RoSqz
1NhRgER23yNt5n88KEXo+mrie0gsG88XBgUfy7+8XORwAjq8IorBKYnMn463
GmIx6hCKiEz2d1nvR4qEitx6OwSKbGCIyyTEoeRuLJja1d/jXiHouCCipXHk
sAeIWTyQisUC2nXlBIWz2vEXwxTdZvJfvD9HtfYY2ZxZBuwp9/A9z/yYB/Xq
5f0KMX8ZYZ/OW4ed63sWp9n56n129ng2Q8M02H2B1UUt44lVVkAzJ8VkPja/
DiQqt4IyHk9hkmNDBwRqy76moXXuaaqi4FmSpAHLd8h9xqdeTx7rBirD5hMH
gY+4PgtjtusvGpthdxi7WxD35HcrDhh+h/3v6LNytswHNc08Iq1hb9w6bKUe
iQXKKA8kG7Cd1694l483w7XbM8VAzdRY9tWR0ZyDdaeUKzy1QFJyyxJRV6vQ
LoHplPCBVJ8fO2C0RK2rhcr7As8+y/zT9VPs5oSXw/Qaij7xY69DJ6D12zhS
8zP07wlHprK89p3C1EJUNIBuJzKBlhUJSTQkdJb3ZBTBjzA0Vwi3CgbSZnjB
gHrDQ6CpgbZvDk4dk14F+maK/lM38XHzk2xsdggArBu0J1kJwh/WUdmvAbIJ
jvnn7JHLzYo7Ojo16nhpVh+lalQL7gCqOmDz5FrmCr2ICHpQkS90GPKpgFHo
NoOJ0EFVW6R3s513no4rLyQ+RA/Sohs6xd+wY5rmQOh+8vq+nnQ7pnByuBDh
cUW3ZaxQkTRLwYpkWov2mXmfcZ4gowoIZO78SVBpMQIj0v2kd5hwwNTGCqfX
ryBoFVcCDGGZoB1L7moyw1YCXsJ3z2mKdXWkW2vrZlrBkt17iCntTieXwhRu
xmx02XfJnonmR6GCa1bKWdq+zNJhYoIShFaBCSfgSkpGWMgDYfuJtoRWila9
WSB3qg7iukqkatQz5ajTboXaTSDVrh4arRiGeaXDi25t7qHr/5v2gQe9WGS8
WM5hZGU+Gk2vq1FwZYeP5xSg3mXTP3JX9Uut8xevppQS4JW72uncIFmo8oH/
IPeWw/NOd2D9x7QmfDC+naJGXO+miXWUvtE2Qs9layP5jDxtm4ZuoMrqLYs1
4Tmf+OXGT0GZ7sG+B9IgY9CStHkwwpWay7hUHwmBU7CjlKs8d0aUCLiU7UpK
GKDHucM0DpJV6PO4bw0hn4TyHHcWuNwVfRmTW6GrZLzQRGhzn7xUiDqUTVsp
R004G3viioFRbe7QCUz5z1n7+xrOnb7xyzGLRnzEP89noQbWe5skpj3rvM8F
gw8dMyqDZRHPQHeTBV8AJaflhVUMQ2PM0GVWWywDewWrNAKtzbXmzP0xnPh8
eSAQyenmb5Tf5OYR36XWuB7VzJdVsZ7cd8MMb/MuQFy10GTGG5O7TvbLJKjl
b8//mqEj8swBG3jNd/XAa7YKQDnoHG8fAdqA3AbRedOPWpE9hdqqFOZXZSFI
iZvcKe0pjzXeu2DkAn+XrRheOpvwkzCVcFNUCe+UjvjzvfVdn6XKa6duTReo
CP8JAPN4pHkhwygGYxXR7MilG4yT/FWZuwscLPIXCVpmMdiCVnjG8PV9u7wd
xt6Yify7YZ5Jf35QvD5doT7WPc0AX4KRt44iIclOwWFSYNkt94Jswb0451I0
jXBr8nBovfh45Ar9lg09d8QPq1fbz3jVQp6cMOgWPQZb7TNcD0IC/nUXVBD0
LnwOP1t2IQNr7niZoyFxVb6IWqEYZd6tuX/T2r3m0G2Y2Lx5FdiYZbrX9It2
+6Vns+DCg2/u8qE6WM2jtDxJlIN6ZSA/zu5ZO859wrFp+Ef/s8rEgGXzBKxE
zvvKieGPBZwlotUh/Ehik3OzAP3Nos46qBDq3ovgObHWq4ogGW9zh6ey1/3K
yScNuymbtmJJR70ARwa6UNpkmIVewR4KcNyOZR/Dt9Chvt0xQP5Ko4w3Lqbo
KbDwEey4MdUBV+qXdbIfHA6e4HQDqS96EpfHdIFbJAUGg+HRweb0o6Z4bzTB
8OGtYRgurDnasK8EUKrJKFZMBYfv/N8wdHDqOsJTHHdpH6wQa5AOlhtsq8RL
IJuTV3Y/BXK9OVHyh0BNBa9DGWM7pf8V/VPbWlCsaPO7bBLotU3FociKGOQA
0eQgIg195MSxQHxSFw2INbJT6i9ddAgH8gdHrt77oVtBhYxnLQV+m4Dg+abS
MSD3uihMd9JFnTcLFU5JiKTKc9IkGt2hsfpC95Asn4oL51AkG5tNXaxhnEf9
figwYBh5n6LuCA+GnojvlJJqlHIkZ8JLmLQVHWmUqdhOvEzsIoWtTAbE7ZRt
9tQEfBJbeYRl/Dx4bSqCy151HJCOVOnPIMAzcAVCKdIoWxlY+JCzBVjZbYqr
YtyGBU3ZeK/i7aZf6Pm2JkI575ZQWuQKmTzacSsX/j2ujcIir+tk9ZOIyQo0
oiQ/X5dypWaqa1jmh01n7lVG26XTN/ueZsMu3+GKc4Cpd6D/trARvna5dYep
MfGPfKPx2D1Vnq1iBYd00jM6otyMF+0o1X4PKkcUs+Cr5Ai+fLpUdbGJF8Gg
LAGNXE9JwJYxw/QsQ5EKfF2JV8WXahXSyM0OXIIIgvC5hHeaeJQjsfW1valQ
f4EbLEi4EVPhrGtdjZZg8EX2zb6Lu8/6QDALMf1lVaXyy6jh0SIGPWkh6qvi
fRiz1MT4An8JI59TMbM2BvVQJeRNkopjhZhFS3lRgv1mE/0zZKU+w0oeihxU
H/eX1m5rvXDdV8cWZbZfeDF1keJNEUrkw3AnQ3hVWDvvu7ciX6Kp4ZlL67j/
MgImnvdkq94Qid6+arAjevzE7X52FvVgAziYtuaC/Vyi13YNSZ88/GtPi+Pa
azU9wk1hrhV9bi+aF6XAwEU6jQbxU79wjDtNvL1SRD7Bpv6RQvFHfplW6yMm
AVd1QcdpkDiMa6S7CDtHjF7acmXdLsIQz/ORBHjAgpQf6Vr1p0osYxuHVy5z
Qh6goXIo0+NTG4KtKV0nbRZ4VWSOpN8mC3sL5atZI3eYxZTsES9Wgm/TKBHM
mFjg8GaiVaZHKVVAuUFDmI3xJLziRsgEKnQou9DNvFOx0qIOz3RHm3HNUobQ
Av37kjgeS+TctLLziOfq/+7Qp1VSNPcHSUOFrSKrBXe12gA8DDh4SAhRmizy
AqlDsmgOU0Q03nBG5+zWs5Y6fVABp9RqY3sKyYxMmCV5krdvIZCbykQboerb
XKV9jxKzTm9LAWEQuKdHtjCQ1PeMZEOOpSQO6O39mSn8OeByj3uk2r3/4cpr
Souk40CiA9wDwnuVbrn+zNE0mZoxaVCKVzGPDT9VE6BBfZCV3RbYRguuTexj
XTKo6QL1VMwLzfma55Xx01Iqy/YBsq0TE9US3FEip6ItmlDYbxoB2JkKM3hS
bEZP7M10gFxrjaohL9igTqFJPL4qDZTlD9Tgka7UajYs2+DIP+wgesJhbtx/
JbMfGCKe6kYav32UgcvyK8gqzGqlO59ijYA1jV9q1Tgi8b3EyUgbFOP66ZOG
SKYkZJSr49sLymQDDLqZV5jgsbIvqL0CqIenDMMK0pX8kRILWGCS73kGerfk
JwhWIwFaUPaCSEF2fxu0Pdb2qTO5yN1AiCet9YHqSoZsEwnJI3jCeCjOgzPC
/wsfWeH7iM3TZF3uP0je3dJwf/SKmhoUqbSZdxxGylMu96NDuiCEebTbpfCh
vGYJBEqUqehhc9gs6gh6oakEN14KuNHv/Oxfzsgx8lPd7RGVV9Rz2KtZ/MJP
kd4R3CfYxnch4fnlHqc8DYm2eLBp8pqlHCtHN1PbXtsjrFNj7s9//wf2oVch
ZNnCYEhmQamNCctfDLyKXQJoXQBM4kf354U02s7S8i+8hjMdCHZ6UYUJTkDF
UzJyyu2H8Of+4hQZll+xhP5FhRAhthFWid5FGW/hGTZROZmT6KHCdrdZaAUN
LhDAsGqxJTeFdqAuv3SgZxDLJwp+LZ4qJ0o+qf3+1DWY0kgvdP9BHnP/f6i4
/+dlDM/1mLDzMQKPGvUi4MfT3+nIDGwEyN/vapujXRmhp0Iz6kVcpxwwt2AR
I9PfkUetm9yNpICAx9XU6kvbNvF4uv7okyibBCVzTDlPeHpmxerc7uMZmBgv
h0sfpxxTCftUogudIPWqUaiTK5o95oePFILV17URXSoQ1kA0FGDLj8bqhabO
OQPcY+U1GBQEVYG9YcklU5i4Q05zplM4entzRga7alCYn1VOYLpLtYsp9Qop
T1NYCtq/L8TBnoXVc49rCqfS1Xj4fuq0F/5Dz940H9mhegM9djBSrzpvlaC3
NeqajzPz0lJzWTOOwgXJ+ZNfo5nJ9VPlhiWLkh2K9vXOT3DJHVP6OZVlbH1A
usZCi0KWvxT5Q5goODbh4hPQe2r+APFsfSOcRkOEt6lLo2+qU+Vqu8FgpSvm
GLetPh0p2Swn1t/5eezogf+ZTbMXjy/mnYpfotER6XPnV96BfwefTqgiLvcj
uOYSQcuWpcily+smE8jQhb3qFq7PgIoe/8a9xp6wXZN33mKx6h9TPpkTICW4
14cZcfJ+pmcicvwnI6yIPifgHtxbiyAvaLS+XoA/dfcVIqeubdggIKPCwfKw
jXjlFmpkzmJR8W0mNlJ6l3tSfW13uoleSlHYFGOxGu2fbOW7nlwQi8EIOGD1
gDmPXJ7XokdhSaWXs9nhPc5MV8+dpjOvmcFzNNE+5Q/4oIGpboBLk56WhtUI
RGH2P3+uJsmeKEn17X6CcIaDRn5U/YaZ2nWtOPuzO9xiHciO2lWWBLKJPFGu
a0CBF9E0iAPsm4tSMGJqIYK+8idiCMOIBRPburh9VwRH0if8nyCmvl4ArUlG
ldzI+v0sDDqnsDs1b0tWpywX5AGlsjivGi2ihxN0NhMSjdmehV0GuA+vGwiU
IauCJwyPWw6WeORFcLO+8HTJNlnqc0I7jIDQYgKsD3MIHRutOVdhxtBZMd+0
LLEl4WvoEzcVNVGxtgGeAZ6h1SEKOysyN1NuhtV1DdcVzEseCvhFk/X1hdWF
UJLviPpaqaNuqxycqx/09uil7rSN12DcvcnusJBPZhBWDieirL/BkeBeAT0X
nEmCIl58raSNmzqUBM6Woi4GobV0HVbeojytCrm5MCpaOuwzM0SaCHhne8N7
qkFkIWIA0O4LguxqyuzRC4xWFuum34PgSshuriwR4jwyPdsoCp0KqCvJeRK7
jl25FVGu+ha98jNHlUngiCVudioHvO060HXb37monKJqiAhrgPUOavcfjqqd
j9at4hC+oulJfiNcr5BYMexzaVxPjVyrR58jHQekaMbhC2ZN7isD92HI9Knf
hnDgZJfXMHoPzgL64kfo+3iL1k0MJE6ogVLNPpcq/O6lmSElSjEv709TXGKq
nWzNtZNjfdXljoYAwmP0JKLt4g5X1eO4mTRrQkPugpk+U/8xYSRd4H3vFYlc
qA61OaDekT6ra6clcAj7el6vmc+88C7SfmWZ25AEt3qMfVir7Ne+ZjIz8+0e
ZoleGCgP4uDJmPuLsbCNBBDeh5x49vhd/ljsZTSaoy6PuET1Edly7ExS4YGr
SvbKJs4r1lxLixI17IPgykcRzzadhKd3Zmg0oxixGpjScSfEqFtD94OcxSEg
h9XaYP3FZlc2gUAlgU2BRr9MiGweNHbgtAflT3E8bLAq6rmgg3EPDOygqEUe
2/C5qdL/CASXe4SVsqA91CEiOkguYop/GmmYSu3rCysLYfZBVBNlq367sn4p
KbmWDDMQC0P/e05mY2kvaNAwH7YusPEsixcB1FEb1rBRB6rLtFf0eSP8Rx9A
UHDNtTQO0RUVc1y8jWwefhZ15k9IltBvrsJLv7mFMEInuSGXOC85r0jX/Icu
i7Mlclzsz7EtKiD/6R2mFEe3+iieGs4ODoctCwjgWjV0g2w4wSyIua7nqSmA
I1G28Z3H/jt6d7DU51/apOex2eZeqUoYdSGIbrzCiKbW0A1zZ7x6GpUSjVnX
rAHX/SbOG4QexwWi4hbNcA2gagxQb0J0KKv55GELVaEAXJPhZe6WoETVn6+q
oY65O3cfmnT2XNpuLWxAJTHMxtX1Xt1gyhWsDeKxRl8Zow/OsxTeazoDS6Jk
VKwhx8+x/lfJi4I07+ubBXwb8gd28c7osQDJKmLh+8qGwyB0KHpFSEgnHpZh
iPKC0uG8gJv9pD1GvKMngy0glpZfDgjYsSCX4KnNabchPXk+9wdHhgYa2mKN
SL5e9K1ZEAJTn2vSUp272OxnB2Iyhq/SRLj3IGM2yP3YsqpfJcfm2FNONaCV
pmrcNDGjSUgj5wPwjrCTSmBv5P5mx0OOkhjH5BIVIuih/i+eLL55gJlUwXKp
aDz2piv/Jstr6ikZzCv/O2KHckf0zZ0FhqT9HqG5CX9rT1g22TBFp46J0649
yCx3R7R1LFoZhiHCIEpEr3YdiXzhL1XOKjOwXcdLRwvPHRHlTRktExlV/FHn
/hHjjl/hNcS3Ed7TEOf66D12TyI+vaK8YY3VWX+IjQz1C7yIJGLrkEXe8Wia
GPxxUjbSbjthO5VPgykVL40Kh4efb1Jl3yUv9nkKtDWgkpNNHpOpHzlL5LeD
zB3MB1LkFhH7WiZQUyQX/doCLJW4q0LJ6ejpOkunajmqYa0oYm+0svFEV6/K
4HaRVtR7aJqK6sQ+4I8y7nBTy+0La43VkEVVrucnH/xQjhoIggk8ApjuMYmR
TuGhExUVeURo+ariUnlk/NJnGI7pu0+fW5B2Qdaxjm/CKhumaPU2/JFBRdyS
thZU6MI9nxSLGxz9BJ7hYOa3svsLgrSdA+fCn0h8iBtZNII1pi7GpnkSSimv
o4Y7OBDTA7vOI/r2I9P3AEyV9AJT8X6zIX6YlpmPsCkgC56ZoZ6pVDj8htYV
QaAzHxRqbRPB7Qj9YzQDsaPUbnYwUwxUVj0VZui5YU/gUr4KUH8tyZOHLk/Z
loo/RBvyDKODXlucWAOlrn86emP8An67VENGI0HVRfdp4Qi5QasDiLfTtY6z
8T9LRnfpuwAfx7NhtYE0XHBdIQpFX6MTO4A4/J+2SaVx5XhKHEM8VsoHAS6n
WJY+ylD44BunZNL8G4UDcecuphyxtvCc2DYg7GlpqvxgTPYuJxm7FHtOwYVv
4dbmqRhv3zBTIeifAyDIlqO/7jwIlWnLbh8YpMH5ZHN4MrADJ3+LJFN8l9lh
PbLWcOaYmOZqpRmv/mXrglJqFhu5U0gRN8JU7XGkGNg8kqrLW99cW7EbFQ+u
2L3IEDiv04Kw5sjeAlb23Kb3zAf1Ojk6K9pkqXBDzYp+j8PyomNRz9dVhLXi
Pn9zyJVS4Yd4UkMU2brG6wzQf4gzHwimhJ6CdEM3SJWuDX03fADxsfOhdMRL
uZDVXB8Bs4CM9of92f6lmAssAt9MO927oNjSS45nmYShoTkxNJawk9wcbQKN
kh4SWIfOQ18QXbbf1dP7YcMtcWN8FMQY/qZqCzPiE3z6y7hzW8AyPqagBXus
BI2F76zjL7qvNldCC5C7qlaibeeQWfC4OQzF/68OexozJwE5MwWFxvqYPqvA
BdBeoC2DmuvdO4dJBMNhkDOSwk5jqi6qiQLpz2mzC+90oqwA0uwObqtOEQTr
UVhtiHl4hBCd4zoEUTvhYOp3X1JEDYezbTARzV29Pr2V3+fqCB8/6elTvwOh
40BJJN6OncHd5Vw4JH7cJk+MKECMc4qK1DPo9HYbgYJQUjNDzvfQL5rOoYhK
2pyDcTQ1LwTfJ5uv5SW74jT/XwfgWMSjxyUNbfjHE4QM9yDtFg9lAbK+kf76
sP7Duh+kOOoECxVsBsSN7yoGpMqfJ/c4Gr3edp2tSuU3VikgYMxkA/CeWFrw
2WXv88BY9HlXDUNn0wDE6KS+a5PTUc3972+cvltoJVFlGo2ggwK69wGrDhCx
d8dkIDhhAy2oqoV7x7JfB4rzJQIvljc+tnZtQ2PpiFW25qfDrxqy+LAfukuU
nFx0BmkT1HVXiyzoWbB0MqQYd5klk8cwsxhtvFzhkptzIP7Xlkpa6h3KZLAd
PWjrgpCYUnXjOF9vfkx87kPyiSPNLMwfSSwbZc5uKxb/o+7TACA8nVOHddOK
T8VqOgr0mWEXADNmYJYyZZDRrm1Wy79V6ANSiCzUQUN3FMESp5qNTrLVipiw
UWw6KkCq87iRT9A7Fn6MBOf2lK4nmsWMpwN7JknP3BBjJYgSICLEZut07rRz
GOQBxk96X+MgQFTuBCsvZi1h3oETlUBhOw/6+nOeuVgtlxsG5Y4gjnscQBBz
dfi4XXGFCNKGlO6py6Z6n4G4L7C2wfmNfD0voUxke55H7f07B1kcAo8u3fVZ
Y3Uhlyc0sJXjcwmvSbs9dWvmODArgtAcYFAuFmYt5OB6Fg3yErcAlIkUZlP9
bEtmkXMH49xOXtZTEBpHz38ENOdhuDVeIsNTUwNzJn+MZxd//3NfEMrQAJAD
/Q4VkEQETiquIpn9kG2wnUGEcmo0Y1BPp1SHEjYakmekgM9qPAorSDM/OWs2
4tJ0EJsd9tSD1Wao3jSeGxNdkNThF+BvdDZ7beytZKkwAZ4iEO0Z+oIm0GC7
PMxQ12iqA53Th3B6nj6o01CvNMMl/sCjOv1MS5JXnjJ83rMoffGP89tN6Lun
8J/5jRW4igPuj5SSe+yIxPnxpBj4/2yVAxKNZOW8cNAmLbe4IPA/4+y1RrZX
+1EnnYibJsLYULAAO/qZUTKiU53v4R7m6AZBdleh1/WxQMuyhuGxVDLQLPiS
ZUXgV2ok2NFztfk70w3AzhlUkllVtG9YmHUS3GSvdQ2ikh07GfxLmYgWWvjn
Y8v9MsLS5wGuv2c17jnmQletkjfS4Cwl60HuCS+Yquni3h+x2Z2M9yC6A2/m
+mlRFoyIhYJ4nnmNDy45ws31thkwpbbG/sDB4zn7e3Ms2mcB4O0JhAnAVelZ
+rbi9O6lrJrPnLIMu1eCkjlXgbwMAplfK4e5H6bPPi9zdd+ea4yGxIdoDD07
6T0xCPucG5MRQOzLZZ4dbVuGcPdsOEO7nzaNHn2AXEEnbPlNmHlHpm+Qv/XO
y6uzSWuRm9cAnBTUQdFg4xAbz41FlGQDokSpGFlbIoOA/1PU0r4lpJYmIuci
l6INefk2uqfFV+FISGC0A1pJoqj/zlCZPaZfjNIbSzcfZWQzJiMKaiKEwwwX
y2gOscdZDJ8i3V02qtclIDFFppjkm2sIpmdCGWsmMOaCngp66WrxIbI5Q0hB
ld+Q8Gz0mQi55qiUctLQCjl+uWmg29vyv4npDNNuTEAVP4QgfQQrOxL0WZX7
o9dBUhRc3OaFkmdnXcHKLoXrPIXQCi5dIYjx1jASRc1LIJk/4WeIEBiv9LWs
K24xrSRGFfw1UAhARX9wAJZTEdDD4i/9FMepAHZDxwoNiXbPl71lN/LOmm1m
sOQJwXMjp5ITF+BSppiQupqanSqCA3DTdTPbPnekM3iucfqyjSWz/27lja2v
GpLihDoFmOEUYqsjof3bmcwKxkkLd6gav8uknCXf1chEzOFm5H/TyMjD6NR4
Kl+GLkN1MH5Icg4a2JO71CxJLE8GjwdtJK0sJb00kg4vAg4xBzDv8hy+K+7b
7V848FdY9XYFHYH7qcUycxcEZp1kToCOrTWCqNpBqk6a4gF/GnFDI5H5ZldH
1Wqw+dyZuX2yMPjYMXcjnprpsSOtmS+WuUGguOaMaqrWD35eflhl4bi9kGu0
qLvaoKOdNTffxBIM3wwGRMHFbxBgkLaV79oWaHBV57u2OZ7aGxfLjy2cgCKD
bOYk7ODFae44kLR77YU+53d8v9e/eQs04Lqowt4/5fg9fEMwmekGqeXK6hVm
sxNcW+UG5bTS7eoW235erZ3vQmKerWcWd32UnPkosek2SBty2NHbJB1cJ7uq
BLZ8a6OsTOmpvXMq0Rgv8Sq8T0tsj/rMqlgWv0EpPMkVMBCaLIrX1/+mVtg4
grRkvRENxAdy8+aZLOQtqwqC+MHVzIzqYjY/skHsODERulPOeM7/WqsVPHBu
jh98HISTabp9WqYMuyaQhh0gYkHz5qicO3Az612ekl74Pd3BrGOqQmnCb6UZ
lEXr+FlBLKBMHgh2Av4dm+ukn/s9jCooKiypa+XxudaR4Wcftuj4ah3WRHGI
7rJHDbK6agjt8PRzPuHtxqELigNv01DTD+2UbqEVBRXvDj+5oz/4f95w1ouD
xAnRThAFdiY4/OPv1+nckqy8iUY85359+XMUneJj/y3rJNwI/DHHfr9zCCjB
U+qLo0cwL1t+0sZj84IJIlT/iMjgx9h8x0m5wn/o/DsgKBiJkUYtbXWNrA/4
CPElWmEy9mLk6eDi+nNd8+k7jxm+fO3GL8PYApQJxC7rgNsMUoUvwpBERgM0
c5z9H57pcTxHXhuQ4C/fsUY5oekzG+SOFhjXm5YBt7WTX5X+uljFL0y/PuAD
d7M+Sz6gG858rHPn0UqkWgx6I7mw5LvB255q6yg9GZwZ/tvdpaLoiaNmbbr+
Ci9JK2pq7WQsVy2BxaLvONHWmTL/jXDODN/lpzvIAR3BXjkpMFGN9QAL3tdO
mswiWz9MEm6MlhEk/PFNntWY3+nrPLy3/WTqA/0NKrz+iPVT1Iv5PsfPc/Pw
Acf+hXUZwEVGzZvFqIsXP2IggoNZKXw1UNdbJGMTbwFQgYW78SqCFan0XpiT
4DWPgyPCHguQK8dLZEY8kKsEoGCA7Sv1feBDG+4zHCrjZcPn8BmXL0d7gA0d
Yp+fqJlLdaOlMnwq68ajfQAdftKVykWLvEqJYMjJMBesWGWGcf/FoT8XK+Iu
/G5d3Wfxe5Qy9Y96XsxZ0DZQ4uJefZ6nfBJQwmfcEBZJt6PUZMMDKZZQ6kr8
fLPO+vC7rNMVVIArl9XpUkpXiBo9y9tsGBRSsFTftulllHjEwgM31wgHSPGk
m0YOzdUW+uRUqNG/Aw/4mDPE+Ujy2BtNC7CRN9SorPJK7PAbKUEAbx4iMiTQ
4u8TekteS5YfG2sWRVrUFHfMetIF30Dx+pilbSVwHtgPabeNFScSuddBJnzu
NyopDicp/lY3IQHAUtm9rQ5tm+WFyiZG83EpwRkSNz8IEdtPLnbz0jfshOqh
Mj1sEsVbe6TBH5S7XKWdMhVmD+4/zeJ6NyLnOIHwy7n3UH8U4+pOCfvUaWzU
mo+uFvNyTAaNNwWaFvRW2SBo1b0mZnINhd8c5qsA1eVwrjGEJk8zq/F5TCSW
o7BzJKvAwYgA2gOAsolxpvXvrnsx5n8jPp4lzPRDP2RDMojpQsTLliypaMpq
uL+tc60Y17C3wfZ3OVCULAIO99eWW5zXuL4NUQpfp6rGA1J37RV73/PsKa0C
T8AIKTL1pxd7ZCHeupg1lPg8LFh0Wn+S7dW4OQ0IpfSBBQ/bAxp+t8kOdk80
miA/NJfyS2teDgmkhzIZCStXFPR+SX4we0ApxBvOT9CptDaGbiGVobH9NbgG
oBJS8N9lOfiNH/k7rXnDS4IJA0WvxWuBSzx5qDHXK0M7QG65wVl9ddJzufzT
GJmnY48fLCAZPbYtXBzU/rn2t4jCjB4uWI6e7XOEjPTlM0Qkn5CsownCohOD
oZFjK+Z90SL8oQ03me414sNEIXlehyE/qcRL67HKrBSfZUHjZ3Utk0NzWUQp
RhqKBjc8AwnzXsDtFjrkH3X18dw6dia71hKE5l6WO31UbvQhq/bVFBo0tWXx
MtAPR8uNKiYH+c8w+hFblG7H+lsVVkdfIulznVx583pDSUIyqnYmXob1P8Yw
QU3JAOjBuIfGhqldWdfrhCTW9cH3x/YSn6uucxhrEid/rSPB+ppJeTFEUG2b
GEhS4dElOXmzqXVvMFDMgbXziUyajxVv8ZRxG9ENAzWvsV8FnPPQcq6CB9gD
Y9NGao+XCGAJlTVUV1MvStTN0JVgY3lRbaxHmSyf/WMKRan8XJBhpcWCf9VP
gjwVvgdXVTYQbIextFjR/MTidt11hho1aRQBLNefQE8MwjktWcHFfIhvRMOG
oiq3z/Qnlkb6BSCvX8sIWfr3nP785pvwwK1VxsIgYGZtcN464Dt75V7JwvPv
UoYbfupFu4g+2+i9neBcLHUmUEJu/7SUlQsJaH/VwDBPATdVreuizqN/2tDY
4F4+yoehASDyj+Yr6P8+aA89VwWJ9oZHHq9/M4mPbscEh2hCZocksQpm2bvI
bhUM1aT942IlNmWnoTHDzZ/jqgARYKJEocN1Izkqv71A+NO+B4fTTEUWZIEH
ESuBhpFJVfFmMPLJvHQTlg4IMwCGweviulFiLpNC85B0WPcy0UfaU/Vzaurf
NqZi5nWOj81YZBZ/KKgu/qF635s6ajhtyIqlalndQdnvGw3dMRCSoA8196Ib
m4FxAhKke0wztsw0fi5chV+WkNVnALkMQVSLlzoDosyErYhZ1+Cfy4laa1s7
Dbp4V1QtSf8+Lc+4GpXz2TVXc3y/aMddDX5N+k4wuGJFpDke4kMrkgtKFwdu
QPtGPl+FaJAVvlYlygjpHJ6s5MMyghcwpMaogIjP2VVRvVdjqMME7gxJ47AW
z/TyCv1cKxztq2AQulFDZomZlRGyrhCaXiHmcvbJOQA5nZOhVKqJXh9z76xs
ChZlRsSG8frjoHkXaG+LjQq0PotE3GErROqfSF+E8gk3aO+85qZf6aDbmFF3
xB+5cVTgFFSTW/eThtCTFp5c9IgAJSWP+47NAG6jl1YYKP6ssEQQk+r3wgxI
naBwT4cV81wPXFtDq0BJhS49vPFFDfqPj2Sjk1gQ7cu9iFcOeEIGTYB7D095
ljagS68vHO1FTMn4fjZX4rZowTrc72oqIPv5znyJ5k6Q725pS42lwPieJ564
MU1EkA3wj37eGiHSDERC8SaYqOSy4VGkm4taSt0u/TjzLhAluuMGFYeNXACc
NZwhwhrfmz/9xPYey4GdzRu8eu6hSckD/6LjxHjaLah5b+DkG+wfI+8PKXHk
NAcflBWxRHzbUYQ/0TjaxrZhAeCgFpLzia0HC4Y1+HQaF1zNju11vyl71UGW
xxaxxtAUNzsW9QHFjOiRkfseefC5A4P4HUAwZ3IvQa46XXiq13uUqVM7Y8tg
PPSk/qmW2VYpE8Wi46pGxzvdD2Jivyw7brqLKs/AEOWjDtqRMZP0p5rpCkTG
kgSIK09UCrKFl2gom+EkZLt8sTQoXM2uo9n0YU6crgh5pdaQ33Y2+xBid2mY
m0gm2iQzxghbV5+bsr34EICc3Kz1pjKvSZxJbD7E7pRPmvestkYStrixo4pI
7U8E0s/nBaz1ViIZRlj6/+qB0d/AHyRaZ2giyxIr4R/GRJCgNhIN1ccoe3/7
Gb3ylQYpI4ZLZZggPBNdPSBI7tXt0ZGwBehuUbqHKwb6S47z6Z9uuiyYgGor
A8DXuw/67OxRxKg2IeWFv7LQiZcF+n1X1aOwS0GY8sBTERFn6a30fwkaFbct
l7hSzVRBpGSNZ4WZjq0k4epeKNKRrBeD+5vy5nGRYJBPLinMlZ/7WTxqPcMy
uZJsNd0UjNEgH+GVDU59YL6+zWd6RLYYXQiGzL4WxnSNomgqhwe/x4WPA3nm
TuBSH17KmKejUHi46HG6whgPzOzG8Hc6MLVEXbHaVuGeqmMPv3BQj0tXGR9z
XEEMmmfGhWbzYOSNd25yr4D+vFQyuZQCqzhOk7EVb0W7giSH8V4EzAQCJKFE
cZHUmfKqv57Al2C+dyvGYjUjiOxLX9W8Wo0QfoKgcmkRIe3/JFjKFBOFuVb6
BACAuhWCaz4EOrwqzvFFP0NXFHJXI6OWy1wmPDe7EsdApMGQRWpYBzgzkgLs
miYMlR7uTUokxkvDVafwuZcpVOuE96+kkxIsoRM/4X0koBRG+jvPGJA5l+ud
0L2Y5WfF4aofgFiMrckSYUVPnIdy7jOdfFkBV7JaN6+NRmiTycfKWlJ0TtFy
3iR4Ubdp1eCQ+APwwP87nYTBHYyEOLv+9XerCVJnvQvJK+XpuYDhDpIQlYnm
9E8cAWTNopGeHsaRMygDA2DUjCM2xt10Z1wQkrkR4UQcdb6V2u6jJlQkRG6x
VvNxBjQLXliB8UxqwTLtNiWuGTKujvh/zBodDLLwRLBzDaUCCvsyHJaseqJR
4/YRZeeDayXKZb7qv9Jnq+/Ug9/ZK4mx8GX2JZQde9dXUzUqs/N7MarVClYY
/OgCDu522ZF9optyIg168LAwoAUNrh9l6he3X+DGIm/rips8XdFaC9uUHzGX
mRzZq7Cu+Xqx22SHurS7R1yF29gyEp3kFClkg5UmJuErZTBQHigmT7xd+UBJ
rJrlnlCy4IMyKFq6xebWyPML3MNF1NHghFJ7q2GdVezZRmbY0VUEUrciEIHH
mQTPgYko9NLqvZGBzSC0MdJiQyxmWU8rYkYbSEHg7kMD5rHGYhWh/PCGcaG3
ycL/LSQNbfbN2Z0/FUSNJF1s4Z9nRkF5qZQZfcMge9NA97uyIBvaNonn1LBQ
SXIU+9/1F+fch5frlrGvKMvbGW7Z678viN1Ta3D7qfOwI5p9Qe2Eg9+mE/TN
zCoaJrhTAxXoOirzOCD1HTYMs5S93Tj8/GPqpjifn8fPO2+cRKpKWnMWyTkJ
dVxFOt1P34MhgqlDpaDYIB/DGZXRXucGJcQgvNaPmbGUMlMXM0Ipnj1kf8aj
lf5O9/9atxdcewb/JYpkTFhRUm6DjnvnT/9rFca23N8LzbqivSsMjiswcDMO
hq0rCc73GFmP4UlVuPsaJEZ93rERfX+dJaQ3F7/G0v4WfpC7JQMt3aXJgpih
MYg0A67cr5bg/CmU9fYek5IbPe3W7GaUTjMUs6uiSGTpWNU2EjZOFv1l3Zvd
gXXDzEm77rD9PnEGBm+H8XV2qCOnEdAF1mOj0kP69DnEXCvbTgqMBJ39+lq4
oDntIqNU4W6M9XJQ/TJh0Kqhbvl73dGVTFbAfvQonYFBZYr+RTBiyijEsbdR
Te38DC1RTW0XvpZidPbAFnVkCzWoIQtUgCyuaqS+MpMgeCacL/u/JJZwgbiN
4yJGfwqknRT2vDhQptBo2wofHDY+Y6zhL4Y+WczcjmHVcdxmHveu2Vc0ZNU5
BZiZuPzzpTOP0lbu8i7HzEO+puAgcKjhQp8bg9X6wREuJy+Gr1GzQVVQsFXJ
NyXuKw9te2jfXXAy2jEXjfg27LtOZl8nkIpF5ej8U/4CJnRWB4C95AG1Se+b
F+8tjrL/ivDO6TtO+cbN0QBYOeqXChBNJYb3oFbTJZRBXzY5fOLxMLqumi/q
TxZlOjZtCCq4/otENW38di/LS3IJF7l4w1Zcj38uIkZ+46kolWdChSdlDiZM
VnX6qDeNdIibJV8VTv/Ud/W05AC0chEdpvoLsCQhn4vV1G1tDUQ4gLSGZ/qS
pb3Cdbz8FZFaRFjHdGEZ2ID936WfUPDgCVwlDleSDWYlwJQH3VlgG52q+qKa
qbAbCZFXnsQKlDuPOvogoTlV+lzky6YDEGj1V8F2lk9MuDsuTn+w6SksJb3p
8i1oBaTGJjgcs+qKpFIS+ZApFDxJOibHEiBWQE93EjByMAUVUHCqS0Dx0bt4
0IRiqx9Y7is9vBrr0TS440eNtogcYB2T25pDMFL1holSi8CYGqIfwctPp7Ln
z1QERPnv+zfH6+NKejwsxuBLkS5BEaui73qa4jdrrTO3MvCvi7chuy3Z18/D
qglyAK+Tjrmp06eYlwGz9axXIR/t3OkZnq1gJQhhIl3Gx1YS2+7SeaLIW/yH
tkNRfXgIU6swh4g70uDEMwo/rc45RXxVckbX1fv6EooxYwHelO2D7NJewzVr
xdU5z/wokPc4eEXu3gznhCaHrbhK8TO16sFPgHrw4GJPESYMSEE4wqOFZVCt
1Sd2Gb0bV3GBf6FEftu6a2v4dfMKtiAURsYfvM7RzHkbeMi9TTfsrLWd5U7h
AnmCm6gBGzmi5i+PQoPcG7ybLiXQQxdb7FGjzIpYoqJyP2EaA43p8Vrpp5Na
OjqvcBHKyn3fzJC9EFLOWdDs2DvJgD8g/UK/4G8X9rYLtnRrTimbeQWEz3Gm
EOB/bbDf6dhjDB6NlIYup+aSlHT5MaRGg79NXSAGnce6bBrTsJNY0PjFXf1e
LOTbHH6Z19vnCy9/sp9+H2fBN4HzWV1q8DoQxA0jtie477lb+KZohDpIOlgv
SJu+oN6XmPb1H4jnuz1u+NxdDBuKdqtb0JebCotOxhRWwb/Wpyq3wInMsWAl
ZVmvcYBWk0hpwzsGd7f6KnA1RiVlXXB1Me5rdAZqxrmiIZBAJo1ASQmiW86o
uG9eAUPuaLBCyumqC6I96/FRR/vdBpUTrxg2SUogPKJepfZeHrRjqeVJWCba
hMX6Ow8cCNLwssv4VoQIVk3jOyFbT0PXffeofYML+07OUjw//hrcSYpKkfHa
h+OGCwH1VauLd7vNijgLLFGy9UEJb4BwI8mjA7kDMX1uqSw1+ga2KQ7G6704
DNBLQlHQIc4D7iwAE3N6rcadCCLmmkfps+YDOUFU3WNrhZhvpK47hgubMPL6
YAf7bxG7zfKcpcy6nyGvP3FL0I89R+gkvMJoqB77Qelm3g+E4wkbFHl0oHjN
qocV8kIjLsjK8YOaJy1GT26HaNWsbdvGB26LmSpwN9j9v8Trtpu2W1twaJbz
0ZSYBnnW0nMtw6R/zZKhly9QC7H8X9CNkS9m6fcJ9v18OHIaw3AzYES9jDuR
4GRa/QJtP6MG15fHvkO0UkYF6UX+txwJ8TsBWrklxNXE+Nf9B9GwUwXl5eIq
RajANmyx+w0e/ZhRJDf0RB74cFGhsmSCjtdv020gjgTxJsShkudpeFbTJbB2
R1TGWObHWEVHWAm6Q1vHkN896tQJ018CPykXfge9pKSbMobIor11W9zaUn45
+gN6Rhnu0wKAb9MRzlyRBnjapNQraN/+23VN5Sj4Sticdwfq+6TR5WOt/oeR
cqVdj65xdcTo9Cn9gawzlHTZglGDbIU6bzGukk1YqMVHM+oXCWWhdnM7whx7
ETPVbtFDRafCLI0qlxoTs7NUD9SoQmEPBYFrBEavnwLxCryQ2lAuAjVkPVli
GHgKPDYQno3toHiPSeIBfj6X1tAd30AtgX/nbIfH2P03cLdJZS1j8bN0atgk
RcFqGAIuD1lrGgcf+y/gRccUyLLtYQzeqaRKtTG1AancjXBl0lmbikYgdam9
NPeKYSUfHxrBdFgeP4OGRqDcqYkXUyiX0axDG4CdCvd/Zv+eqOMwchP2Ca2P
exlI0cn2bsbWFMpAjC4TdIvWIyhaLOTnDhX1n+4CmX7LcDAhcPUcerInjUgA
N+UPtgLQJ/nu+rW+7txW9f9h1tJPvQP2jgAzrLLpoJ3qxpElZ5vaQljHuhSU
yK1GbwQ+kUX8vWg1zKYMEOOG2KmUfSnRB9gd3G4tfphOzzx5/nC2KpXaflVP
HGeUf4bHql5/myqO+zsD5Q/FYxOfjEA3S//zHfLtIqHiBGhrneRgux84CagJ
9PcK0Z+EY5x0rlh1HkYGvWYDo+fVt81lv8aFmyhzZqF3Tnjv7QUNqpEi2R+E
BD7k5s5t+TuD7H01CgOLNu1+lEZEY1ukAGUBg7j7M1RxnLmOs4yjW0IQHkx2
r/mM4GMdELidDIwPfKUlI+/QV1Ja5iUj0DDbLbcNRqTSOdLmsZidwkUwGaZ3
+NewEi3cBetPxZQv6reynQ58mIpk9qqiWH7LBQLc4d+C/cRYa2rBuA5n+maX
W+56bkLSBJwbeo51Vw9nqwGoz5WePH2mWkjXwdzNBPz8nEo+x6xBJUgQmIXJ
4GC9yygLzZdr3DfSBygen3VVakN2WciduNLOQ4yCmOZvXAqW+fz39wlRXZNR
7jnJSS1jrPowQVNi76TuxXZF5x2fPrb+M3XqdsvQcFgXN3xiVsKu0OxI44pu
lUcp0KXin54E8ud0+dv4yooD+uue1O48ONCeoQ/4aFq0YS46cyaSRhp/hHsQ
S1P4dEj6z/CtopyhTBf9NFJ9mEVl0eAf5bovaO7H0IDoRZnL2n7MeoM181ZD
M5glL4w1518Cnm92SMsiB+pcgehzVWcH+paLs575+HnGCfbDjmGGMSGbfYn8
A0RaPiueg4aaPdOyrEOkJCLJt4oAJOys9E6SNWuIN1Yw6I4QTUJVmc60gc7P
9JYcrHTKmmnucO0lKfHMod9Jk7ZmvyW3IfYTR08kN/XlBhhgQFxVS4QkZ4WS
J2Kh0RkEA0sfzehlfK/jR9K0S/Mk812SikUn0K9AHGANnLEadObwmtPJm3ir
/i8D13zNj8bim77wmVREkUCtPFjQQ0wNuczEsXPyKjhenurS66gP0U1SZZ1y
K9A+9vi22TDaLAEsNsNLQRAWJQafe/Zn/sMF0TpE8EMmQ+N0SclXYN2m1bkz
AuN6P4fwxORKWF6FlywLQBwm4xqmA02n/nVP5fSKTiW9vrTtBZs4YPUlbo48
GXmDLOg/sfCpUspNQ8HmkJO1v1zP1tJi6Vg78iLdQOXJXIMxgqNP6MxSTePI
PFveYl0/dJCdjQNZ8+b71ln8g4OGBFUv/dIDHZVXxU1CwL9L2cet+uP09a+a
QHigOXWyUDnTyEr/9DfqyAXZOOwYHSnTaZ5UnD1RiSftn3JDhpYb9iaDbtLB
gezTNk5D+6Yv8tvCY3yNFyEcImqPSBsTuGJ8InA52BHlHEoEWeIe+r3BNnYx
JP0OG5Xngd0JdVvh8IxXGViTfeDIh+Ww+YdqsADhWeUL4EnjnMo+31nCpa9V
2cpnYX82QQYa8SQmOsrnZcr6BfACzZHSdI/5P1ByQdURfTxvL3IPWxQAzjB0
VEc5fVjav6KxUY8Xtu4k+8SrGZfHFbV85nIaPdsoE6H48d0BXG0896ep43sv
FtRFDHrG19QW5pWdHX52+8Ej0fgwo3LACny30hJODd/OFMkgPVtnJR9esEm9
H2Uz7wXq9w/zlglOU7AwhwryJVKQVRD5XlETSRoRrK+aHJUTHhYtsS68G4m8
86xoE1GtTpX3vf0PCc6Gvd5qkY/5p5iCY2MZ214vyKVyYs4WefG5fUqxyFZN
sxJuRUxyIGCsa5evGldYDZdE6tvWdk60bWbrypwLUs59VDR6JwbQgK08GitU
O8yW9oi4qKNyF7iftxaEtW1SeQcMXGUME7yhkMriir5TkSAAtT1P9GAJVanC
fjLRL+MpLdc1JfXBbl4U2YzwW0cK2UxlZBL8jRsaSSFg+xHeiSc0J5SEp7Nm
eSxGAZzud6UrHg4yfXkn5CxXk2F+LG98oAdHnO1pLDSTJqjNlEhhKPNnOpOk
Ok5LL1TGfu3unxD2VVaR5b6YhIlZsvLrT8rrBw2NItkM1rMFp4zRBEClE9EB
I2W7XR61an1v1IB7US3TuV56Y+yh0vUKO9xusixd4F4ZYfANsMrKsvCKlO8t
sg1QmyIrfgh/+pgFYfB2aX6+bscTj4QX9aIClRiEdjRP4RS6w9FvLChQ5lhM
BAMYz5Z8Gu/uwJcE8ctsEfl2igBqyy8I4UCDCjf2p7tIVM/dcOTsv793tqwo
T742O0oLbIfYP+lDHYrUrWNYkxs9KA5k7bDg3aSLuUpWvD2AAk0N0Vln+4KX
bwC40yr0lZezIunSUHP02QcvCT0cwtRY1e0AaXhfI9v2i2AYVbzre7BPOyel
kgnbzmg+A/282xup94qn5voGhwHbN/+kpqv0blzW8ejMNNsbd/6CFVZKHl9L
bkAPdPOogiZbd73Yq+qrUxYGVm353UMVs3/2lhILJaIsfeGWWT4j8wUeqsgw
K0QNUttJcbPHX2box2AEcn20XFS177KTbhVexnBlf/DroDcd7vmogRIwkNRG
cRS9c+Z7TwEzzaF3BYFUrtKveuDgUaRMxvJw0NrMD/riIL7A8As9TUbofdPQ
SjzgiR+1pBt51hIAGR23DcXdIfAVPaneis4Ag/Lv1Pk6vZ5D/h/6B9KYMVSk
ysdng8yfFJa4czhuXan/MQqPaFIyHdkQ1kOGaY4U+XCEJB2+oLzpY2J/qOBc
H3GWOu3gMG6xAzuthKdJIVMgg5UXj/Z2hBkilnRwmuIfmN1r9ZfJxu5p0YPS
XiUv7D++BOQ6t4MIZHTZPDqT6K1Upgu1Fai+fj84PlX+Nup+J5+8uoZn60tl
cqwDuz+1mMXorWsw2rKvwo6RKPKUyJvuKacaP8oHwlrkmTDvowyO/c61ZoNy
1vfQ7HBUBYyUUAipBIOO2cvn0CpnO3IirYeNYBgynJwFgeuAQ8JpkftTZmWX
zNAxidHihwOerp5NNS9tWcwyk1FSDw9VUmaGFz7YlIweenoMN/flXtsT3zbz
ARn+Hy/5wjwLm3bWBqC9iOp+JOT031Vt4KsXxm1DAmo1u+arFB1p82H8PKRi
ZBue7djrw29KUHwDQtazuf49y0YyAId1wXrYbbVhnZFhzaxtArdJaA7GvFYa
8kWJMsu64r8QAxq1bOIHUzp+AXKVAIGQyoelWFDrXT/w7Well4C9kO2sQYRK
4CXH5N6nRidUiPrcnwgtUk413+u/F+t2LaauyKpZVZn+VKqsnqFCiofjBRCS
FhJ5cltlCL+zRT39ohApwafuMaQSL9ZKdcQVBMYrAEw5NyBbSKOF6HTDORav
AtdlN+GtRaOLqAII9kHjkrocXfga8+ZIv4UpYdrJhMkwBtsswId6B7eH4AJQ
s+WzjSzKjpc0DPn5ELQbl8YuFOkrvjxjM7RajT7cM+6Mn6glW6f7DX44wz2H
PronxDbPCU6lwMGTYYJaRlXw9u4FKTDDKviE6b9owHuiIo0m4cTzy5J+AU6l
POyD/gssT+jc4T4xzPaMPuOA9qzooxkEQd3omINaGF60gOH0xp3OT6O1lz2w
SqLANvjEPcBvxZ0Q+Cec27VFkV7KAqckDUcPPMMNID99WRh8+mDsJbASuvfH
mPqNbO0MyjsdTdbhwAE847xv35Rtx22a3z4ryrBhpUoxKw54Ame0EeTLBi7n
FOY18MvqNbjJpaccpqubn185N4sD+1M0UbSk45ViwE7IzdeQ63zgi0QjC3Tb
FmXCEN3ihNFQuTD9Pio55AHKOIDO5EprJh60gagMTTOINIXI3k8cM1e53LWf
WikMQqbyZPd1wi/aX3Cb87EuXACnK+inVqhnXlcJWbGVcw7r0fepqg5PcXYY
A6mxdptRcxQ+JOkFoojWNdVdJiYg9OIxcId+QmFENwJ1huVH4AOva1TeeOa3
ja/hSf+huPiAKFb+kf3Nb3TsMLvRQoWZcTXEZyNP8cptAf55hAlos8rThyZJ
jqe/pB+URQihBy0ia/Wsw9Z+coSVwo00pwpWjPLhaq5pBaP8rqwigP37nXKQ
sevYeJELUSNew42gNErYzj0CFuvoZVjkVkGZ7vNHPTERCIRXR4KzsP03EJWt
kC7QoEq5nEHJQrDha8FiEKEfPFkmR24WgTPavxm3AlbNRiSkegkuI/fdO87c
RrfhNVcBi4gmhxCAjfwxEml/OdzManwUrzRem8LbyRbsZKeaQlM84TfePpSd
UlGFcttpGvaTE4u8JZpqOEjKF3uhnDAer9Rcc6aJ2Vftn4naGVJQXTcQa//X
R3Kw5IyqpDQZduUM9c/5xVKyhR9jFRiesHwFmRLAgXD4daaDBY2ovwYvy5Jh
0k1/xacGLwY+OdEyQsV/v9iOJrtRKTSpdVnZeBunhyhaibJHm7vCmwPZP5f6
ESSt4k/0XjAyjDSphPTOauiM9qIeTOwbqcub2PWGwy99Emoa3Q6ebFiXkVui
iuarPLevOfBT1CgmST05456R3ESywvmsgosMuEKV/qlqHlcpvNxtHqwAc2k0
nmglDGDjemO77niMp5I16+MKm3R6zdwtU5xdAqSp9RREs7Fx1HrFUm8R+r1h
WeDDblpW/v2a2s0UscEdJsMrSYXb0PPVTnXsx+tTmke8bRTUwAYOtnzql7fE
XPn8rxBtsOBXASZIwIA3RxHnsZvs3sC9pcbT1HqjwMJj6pfO8B1D6Cn+2IOp
GymNwVQwvA8I7A5pfPaeU0xHZG772/WGrZ2ucqw0crSYRb6etZsWhHGWsWzR
3TQ6Ga+mmxCm4zLFB7zACq2ic69GKIYVNrCcub/q0hKEquBWlXUvxJjRU1bx
RtX3OUcCbL8rdGRKPEw3P2Qai+S0YTPdSrZZRpDHXGdAD6lWodm5jdXo1Cap
ov1y9yR2iP93PyE+wcXgu9ta9Ih/4uroAyWNVQQ8UhRP2NVZYsF7rztxDaop
oxVp5HIwb6MI/lPRNHpfTfdps8ojR9zRLmaDuDDDm1uLRXlNOxEy4BHs6V2l
nof7RWCZDjvVDnxDIDfkgGIiQ41MEFNEoTp9QPY6x0XuvWJOvur2PfsSHq/z
UTyrn3HviNqRdU8bOw5oPrXO+Wd7VRkTn4oG5ZSRhBkTUb+sSlJVRQfJ965p
WYn7c2GmTs6wpeyGfMl1K56UgM/tw2Hb6xzB2qXTw9cNuFXnXbfzEyDv1FPg
JmNINwW+s5L+YWAtb3+G9WET7toKyiNtmYMn3vTeC0i9eEI3K+fW2ZP6xYjB
swFWvCNxUrCrWmZji6nx6S1sz545gjGigXZ8HoETv36wziMy1GV70S76+4x5
0d3bUDVNaM4qXbhctdb9FTQX8C/Lv06Wlk1mquBjLm2rA36pJTXtt3cR9t4y
ykWqKYSwtQU6t4jxZOLZu0k6R/n4W85ED6UkvASYtbMNSUGKhG6gH8Ef7qsm
nk9y9iAq5zEcOKJ9KnQHHaE6KW6pgmdfpqpM0tFO0yszNsmp0N17l9J5ysyQ
YSss47YOvMuSnuIhQiDK1m4FM7RgcHQWUxxpk50md2dGHJVeU/N6FeQuW6EU
7z53XKdJH+TZOBIw+gtfxeRw0FalofHYgImF9iVYb8SAZcyBqR6VznAEl6Q/
14ZaF8QqTFGnWMw1aXLhU/YS/lII6rxbKcHBevPfQ80D8JNKehmPhzNroXFN
zikcVFXik+3TIAMKQabLrYonmWzfUQQ+oCADUUFgZj165iUhSu+I8OXy8zR8
GaY9yfHW95K5PY7Bu1sVVp2Bp2CncIGOBlzuqf0IGg2Pj7441bKr5FuZWV9l
j7gSC+1tzmraMBEwoYonsN4EC/qo+ycb4RtwgFiI+E5YFMwUsOAevLPWy6jG
7Ggn4qZ02xguBvh36FwfIFjV5Vs+V0I5kKIgYEQooW4Drh9CR9ct7pYyfAHH
D0tVq6ENsIbOOuqaBTrU0Ybd8xvazYqUj9FslszTPvol6/S1VvGVrfc8mJeL
ifrmGp4VUPF9E7fnd2yNKhDCmqemOGb5IDGsG+pIsKe7zMOz2pTwr1yHFbtn
GqF0AHo4bnec5SNQQZl8/aCLHZWzkOOdLzw2bNGf5H0FmylGBUpZQjideAfI
BS7LTfqh07BBUuvDAuqKQOYr5Uq1K9kCwwPIa4b2WO13oV62bKDFlD0BK/P9
E+0P//YbJKXyqVCS6Qcmpka7rjbbthAreKp30fDycjEtkYYGAc+QLOwXM2iX
EcKKOXkKQzwT4GECWbKH27o7U7CKlx6deeWHvC3IRifFLrnef2XOz5GeIT5X
797cZMDwqQ/Y8fj4kKGZ7R49l7r45blbctOir67d3mFrbyaMR4q7VlDXba8v
Dv57ICq3BRGcv1byfsD9TZjsu7PRnPCRGy/OW4xVw/OrFFET1/LpweO5ibnw
KcI7mSysZ8edgvCQai7/q5WDrELFD5XPI1oRHZ8vjqQPoqA5H1007A+Pr58g
OYIFSvN2umH/l5Fw6uKouKe7Ev9ie0NuJeNw93aPcdaSr2vXaqo62R1w9+gJ
RI0sV3RGCqsntYW3eGAxdFVPCY29e+6sH8nJyh65v1vWDyd9ZCdiImsXgEEp
bq5n3FoXVmmPnvvJsqadryx65iahTOvjGNWLhfSesC1OqV/bveVfnVozyM9Y
BBxBE4HSIJrv+3TMy7pBFOEyVq2y7/ORlsYjWo84Bosj4z0DhB76p/GoHIRK
zax9868C9rdBM4vytYlfE6QegJvJeS5KS9MuVYIGhmr05bv6LSF84B+IeA+W
yMRTFeJmlTg+xGYAeEq2Lj7E7AO65hRHGHeNH1CXh0J/ywKQrk0l6AUSVaJw
roAr4jAatjUmw5RwlV5kS/ZkIQMkJYdpeyad8FV7QDva6sFI4mjNGCJ1sfsQ
Krq5gy9ZDFDXJ+v2jBIS9oV5tJlXrWvChfPDqJpMvH36zRUcQer7489omagE
dipAO0TmiFQK+sbE2d7jBNwDrYOgpE1hSUe4iQWcEKnRZzTagSRSVS4lOFrm
LTcOhqL4GlJoWRHvAfpEuiEvT+G0umBuJ+wEIynwJCzHSR7UEWMjCdN3j13N
39fcu9Aq8C3cuf31BuyPaN4PCOiPCxgLMAYMunN3vD+JcgmNKbiG2WaNHQ6T
zWQ+0wZqrX8XqrcxW3O6WRSb3ge7/8GV9IX/Z038mYFpOiEpWas8sujBpnuL
LHWAkQxWBHPwBubqmWcYZnsBghEO11kE8nfbzVy1BTm2meC9pqFR4VCUw0qy
DvtA4UmCC9hyj6Yc+pMk+KcpfgAkgQPRUcDl0/X/27NqRx6lxQ/BWDfCUpSV
k+oXsq41nUOXzOiZOng8W3DvMzZTggZgIKJn879zpT7e8mvDOLO46r6peVSg
88DQOJ8rEqYtVdyyYnWZdKv5/nyZLKeYq8pRYvqopR6c6G48ngGCmYIPuOAH
xlkEOmzcb3JLWZz2cvGn68qs2NDSyXtrY79hu64fTFjOOIxbR6F1EoRJMWnJ
g7BBy6/66LwuSl6tIgoFbwTPmsAToLlJ/3lSQBudi/XQ4pahKPCA64tIWp7S
q30WnMhNKCBKVX1SqwSo/yuGPWmu0bgdxtx+AHBEd2bw7YUyoMxTqyax31Ye
s3+JN+HUfNvP5aPDHo6wqEqXXa3clwQb+AfNcFljESBFgrBx7Zn1eVY8xDf9
+EuCFyH5kZ3NCSfA/loPgabuvUgmIrfriHu9wpdC0f6ZLvCjyXHvQOpMoqxU
wC3AFLo/8+UExie6oG0fioUuyNIXbE2nrAR910AidMuw/h1q/ifBJy60uClF
mJL/PZ/fawnepzEsf+NY2F8GqNObfkq6HN9luvMorUHZ7Fd0uq7fHe8qk6T0
eKJZ8kcH9tdmR8kCL1YhF+D9RGor5wY/TkgMgzhWyZjbGxF/RAKtRxj2alG4
M2TH9e2XGUnHKW/Mvnxc7VAl/YAf1L/tzLW7f6gH6HKC1MAU9cBQjAuX9B1R
QtPHljayV8WMuv2SSKOGl/LJ6RgtuGr5Oq+F0vtQfnzOQKAXWPTODvwORAem
IktXuvEAarXT4rX0e9fIPDB0P8LKdOyTs26iiZM83eK1Xp+U6N02VtgjlRow
sDS0Hc3B47JMHHUuNlYOwRlZLB9geSp7OJwLR702kQlUyk7cX/gVtGD3P1xX
zqjND3vRwAfzPKD3w4LNb6gfbM7kBEjKEk9ttu0hKrhJ5g7CUpN3bh6Z/71Z
00t+ReReKO99G9P5mTMiDAbjx0Y6BZCUzgMVvOEOHHebj5MMBdepE2BemDG+
P0DGnQ3eeNQ9Bl+Nxq5LWjUJmtiUiYS8nPcm7jwbh9Hf24eGPY2gMeDEH9of
NKtTyHFNZXX9he/6i1EzO+ivDgBEKlAfj3ukc22RU+88R0KzkGfR/4ixdK7s
+vEmt5weFJRPz+bcixD0inVBw4qFTtIpTV9zPnIjQqdopbOCo65r0by5Fyh/
u/h3QP7kKYd9KuyeW54nRB3GGoVuB1f2g6+MZSaHQm7liwewpKtIT+WcIr2Z
HZvIVEQ4BzaI4whlqkoGkfAABGQGY//0EdJt7t+GMRTVHvirWl6HeGlnu6th
VDNapIu/KnUx0eqDnIrwFIDLVO6rzscc3CGoqDZKYlHoJyzr6FDEwZdMkCKj
TR0eGFNC/4EIvm5Jcr1/R/+26RRMEscBnma0jXFUlvzVj+OsMhN4v4Q/gNuO
IpDJ78OQo1aePGU4SGtvSlkjIw4zI7tT6a+uR8kXb5xxC3b8sn3SvaV12aRU
pdGKf7h0lV1RcFAjQMUk0+8u5SF2IsiBelmGpDcRPcV/iLTN3TkvJMqU1x9C
efORy0GRZVky8fCSZXIHj+3OQsXU9hk5pyMnHkhq6y5r2/Ss09BCeamMmLwG
rbGjSg7ZdqQyvKvx6wSvAI/Oscsl/5R5v+vNkeDOlQTC5+/bKs6gBZVZBMQt
mL4Sx64ztef2Andgz91LrkMhoZQUdxp+PQhbmuxTC+9Dcrv0RIWZYrxBBYQW
8KcUaNMQBikf3JnmWMKThmUhHx9/DvPzAE6bhcdynMPPjA1fCohevTbgR1Ww
rUQOByjsqPxn7H/BcN6bt6rSO/eRUUqbYqqIpn0G4r4/bCttScqgTHJy8e01
6SBuQzmyxD2PGm472bCLhKUO+lWbzCjCguwNg1Vqzoxlb4oVL0JVuSu/DKeD
H/YNa/Y22dumbgtA7n7bjch8Uyf3z/XH9f59s7CyZd/fjcCtb+Ae0PIf6ht+
AVB3hjFPOlRGvmtVRR4yUkyX1dzXkpPJKRLmDngTV0HWD5qtnfWsWi+AfSwn
hm5RuUtXQfcH8H0RuNlczyzjBXFN6Pp/pIU6fECMAZO1pCN/i1V46jr9QTU2
/Naq0e3vufiAXYH8rDvBbz9vclwyJ1zC9F2FMWQh3Jvo0kQg4pz19doDXDdj
oOkj7NLD03rP7RiHqRIeokqd6WekoiHfIPD4JyF1+OM07m58O7ikMcBBIz5N
luEL8mnbp07/Km/vprD3w5Sj0EAPYjRt1JwR7EhrxD+doRwbDuf6xDPj2o/9
mOCzVeakdUT46StMsAxp/WhOzj5iotbu8V5gki40hu3x4XmLm3vJKKsq8x7v
bMAMOSSVSKwRSfPUI1H/OacfyU1z6xGTopqa66Y9tOjxO3xiXwaMf6NICoPa
nj9AzGmIWO2BnN7bGbnAkTNVANkr8OmWTSGINtmnyDkJ2xTSDLevWJruonJ7
6cxTX8x/NKHaEAO8D0H1YsZkD3hCWdeYNO9rzkjCevn2v5bdqSJ2LUx7xv24
c5QAmKgIxkTu4AEA6R+/wAPwomPaGFA1agcL1okHFLOonjfnB2fmJJE7D7O1
xRZY7+jMb1OA1DCuPJIbk3MPhaDfk6A18oVmamTOOLDOBkgnER2iE+gKkzx4
O9InaaoS3PUXXzBIZM6RjypH2uMSCE5DnhXmfeHfe4A+ZD6PhQ1bOOLudvqD
Inpw2yLSI392rieQzJIasY5Ky1or9Ag17u+YWYgyswRE6Y9RCsq8m6xF7Jdg
hgvgCKuVbCX8anPcWc4YBDW62Oubax2zmLLHE02mdm2dgTgN5gzWmE3r67sn
7saCw6B7APWTwMHTZ1ENQyV/+Ublk+XFzWur/ibiPuwO/dzGB6+tkSsKZ62f
NmWnoR9mJEIdcOy4DWneiFyUiOhNL23zqZhmIOGgLGeC00/xmxIfXkfAilmd
+gVsO1SvQMhOynwqmHxYsnsWNv89kFzz+L2hPJYWmB3aHyiUTwVXs3V0vE/4
d715B5M/dntJB7v9n7UwlSS1xXZNZIqJqea59MOta3GJlEBweM49S3+YZHb/
zknpr3BCKJPI54O5sRw05eOPN5ThFXaLnPxt8oZcGtfKId2zCtP94yZccTIg
qcfPRmtJo/JdcA9BqqAE87pUESIJRkcwZQbb6rFV/WjHOr4cT3JlfMitpM/K
beG9t7ttjRStxMWaSOVCyc+YfW+9uV1jh21Ks7I6X1eHKl8rABclsOwKNwPc
z/aPmFia+mXw1JxPI9UDuTuwr+U9IKJ3uSE+ZVbfYk3iRsq41n2osOhjVCDM
HqcxsjDR1Dt4IaWNFFwUeNvN1DTU60typpdWypj8IkCVRlZpuAb/Da0XLmcK
mlxH2VJ/z6kyR+zNiST7CaFbL/pzOZAL5g5FnjufJ8Rf233jfA1S7gIgDWbz
pD1FDn2rgKu3W63dNXq81Y+pbkcfN1CSjb1LBYCeMTo3r7k+UetaXp6u2a5e
qU2+QqLipdVNnSviPUDAZuyokqbpxsTiPk+onACviWUBH2aSfU6Tsbv3AcAc
BnSHxWCs/sw+0y28zxw2f9I7Ni9c/V3KT20D2BsHJZwX+1n8Ck3EnQY3j64t
DffqEB/x/mcz9Aj1zjLM25Ko2EJd7t0nSmeAMPo/7F4h5IWviAEmkdBBYgX5
j1bsmSIKuZDGvGw5QqNY+Xd3JunlZRW+b68cfaUaYpBEjf1TCT/ogUdrBNnS
3QAQqiZSgnflPfR5NZIXKlJwD8Fk2hzoac1uhdIy4ALa/B1ZH9Tm2QogJ3Dq
ijfaJ/v3y5mgCGbToqACVhMy0n2pCyfGXsGOFXYPFOiQ1yWk5POoH49eZGn/
pC3i632nMXTI0dqrrijzVQR8DLZQzstIwoLjyfNI6P8y1IQcn/IiySN39i67
xhjO6eitaFo3z2m61rfNcasq4EVvPWpe88INHbi/A52J/UR1mYKxBfyK8fg6
WtBmCrG98m4Z87TmorKdiNmyAX3DrRwXU6CfpYDfUujXzdMu2HGOHR07Xzle
QwQUY7A9IdSYWpLQ5EOAyZv1RFJejQlr9eCaCUKUP7G/jnVUHPuEfAi5sDiI
Y7oVn/WLIdhg6W4RjLszGINUgN7sY0SSSeC5DvAd8do1Hts4P85io4PijQTt
QXnXGotjuAbG9RKz9WlitKwxUPWa6ltgfgbNHFr6tzqxbuQRS1USsghoLvUC
bkFQixjafP0HSylyvJnLT3+qgs06HiYunuBT9E+QyOq7w56H3rWt7sTibrG1
P0iDDS/4g/ySbiAOHJeGDLJaTVDhhVk1eRNs+PEx00QjinLqC4Y94KyodZyw
vCpq7qyJplq0HUBmCTJR7O78LKpysirqoVR+ggUG8ZkBxs7s6rCtY4LTXjab
Ud3P+X4o5BDglQUKEOB4jv442+m+s1px40eSeLmbGWo8H3CQkyFFU5YhPVoE
y/gReFT1fRQJHDiblZsR568dp+m09pDHPaUH7miNTWfMeGVUaSmgdlkCHj3v
KyPil72h9egI86IaWl7yzuUiavebe1cwSscgPWLu58pVtZ6D00gOSQDuVPvd
EXuv4ottcV8CLLD1lVHzFVnnN1FL48tBv3ONWAsE48n+upIOXu0+KRL2sXTd
/BTvuml5S1B7yVjZLZC0sqhZosWnH2nbsT0VwnAwRsj6SLWLmTsNWTFwgLPX
D31HE/2z3rfiqZIo8YI03kVkud8KrBvg4IoBpHhteYEjB58BcVSJl3WgY80u
xQcZr+SMChcWJsD1udkIQsRKDIjMETOG4St20FfJyDHoEpItwuIfk5fmZbeh
eV/LDuml/ZeWDColBUkr3Qn8FDLYM7AotDD5s25fwea3GWmyrvJN7Xoyn68k
oxx3F65vpUDuKDti8uoug8yk2oZj7Fe91pxi+vDJx9NhPcruuuhUR2h2A1BA
Mw3bRin9nBwwWVuawcvdO1bvcLAolmanedOD11STwitiJ6wotJGFh4pyfb8L
4s9lYjk9RjLsMS+oawLehURVQ623l4dRgKUGrOEKOqmxegUPw+9OA1lnq/um
hNQNTq1gqj64ElT/VKHr3v8pnkdU+ZIRf+dtqI4nGCaDL9jDa5I1U0laQFde
ZNoH1r73xTDZAHX2aHRiwdVzBnK+CgWaUPMzh8tYtOSernz47DpaSH4IWKhW
GmjPx/TFEAep+P7nBgONTKpRoQvOnGa15Y+1GN50mFLFHxF68LjDKmm4oRiQ
cD9YzkAtaG/SCDdm7qvgMOWA0CiiV1RT31Sq3tGhbNPoqr0Rcz/TwBKwZVhv
Gcmn9Gotrmrkeo5y7aOGN8PqP8GYEQzvZdRnMj1PU0QqQXaF3fv1owM90tpd
wt8bSLkkvxOyT4/v1xZRe9YnzByVSTOI5s3G42bhP2LP4LzrK2+Pf4Vxc1RP
56Ue5mY6hr3V69jbd5/n5iAZY5a7G3Eolcv+dFyA5K6Z3ILVfDqHeax0VX0O
WRZLvOqfHZ7w0zSxsqAjHaRXJj/ol1wqiEomSd86TOxMZpZwv0YsEAU6LTHn
qUA8HnPpndwtDXd2SDniajA2LdGgnACZrKZ8uddZDHtU+e+Oydi2Pb37+ku9
L2FF2E1P2xCwOFepX4Fij6GL66a8HzArPgtlCzNRJreKNFGpz8Nf1/j/I5jV
LODqwk8sLfqFVIkZNyrpiqOEmwKl+aSWIwE/a6pzcd6yCPfCkoQGWwS8b/ex
t2bieNZuTLt5w+yyzeSc/Vsmpc+U20YuZdtcZ7uKc12MBdI2bWu+DhuOSYqJ
bd2dMfZWWn1QhupSG8nYWz7uMXqWBUi6Xy5Uwr62akc1XXkc4eT1nXgPmwdf
EtARMVur4ylSZy9jne6Xy9ACj6jqWZAMeXzimvxsiCptKBhxVxBERDFa3Cu9
RtYBTYXf49brHoyBmL1fcHjVeo4dvwxqQ960GFoFWA6VoAy75Cxzm3XZ2bYx
GeDKjhOeTbIQ7IVXurfK4L/8as/am0AxnZA9GBrUNUEddRJGF3RfLqSafHRc
RYhdZYWFMLmBt8uEVxzllRVpsp4rJEMSl0ahin36mecZJoUGLzC3aP/AgqD1
Hq3PCGUvnnM1P+hWJoLNMbQ32p/UKpQJxn10YdzOvZ4SWpNuZLSlY3T215fj
decQeO3aPRWTUYYRGaqJvEEMPIaKeTmGsH7nV5dpi2IEECZmBArgcil3HmFR
LdZOYFH2ETQGjL2/QrlvqbBQ1swlXJl2SaFKkAIyLG1QGfnXqd0uuR1LMqN/
rHZtjz6DqNnM8N9tOu0XOVbmnMI+44IUntf9WqyD0g3OuvWF23Z/yTIZs+rC
PMh9mGUJ/pOJ6R7JJczLyrPNOul0dSpcro23FABdKmYX3ZdWqwjppSdTy3s/
YIPBncLF9RfHTKiK2z3COEYLOk47oKh7SDFmOZ85o/4wLGwfcQSgEa6KcsIU
J3yXJgbi3IxI+/uMKCmEonPviT95oifJmZ2POMlhnihTOShczSVoDA6NBzyv
UHx+V8+rgCa7QBoblU25hpb7RH9Z//sK3n0xnDsN1SHoLjwSf/CrcKzQEoQC
dmn25jvZkHFTWV+bNpW/sZn07gofJW91T1PKJtgNZA9NhZaB0euAz3Nplh80
dpjlDdwLw8dyRU4VYnW3bHYftArXoSeOT95j1zeGA/XtakMPm941BRpeT95W
G2M6Q7lZMN+taZVRZjYJriM56p6OhpXeT3e1t7jxOeIWow/hfxmSHhiJ0may
L5XTzeyIW+g3n9BcVPBGFJhucBMInaHk+ulROce1SUHL362TBYdqOSNj5NX1
XPlb5yWaj3eoW76Su5yLysg4mEXizIISVKklKjl9wgStEJ+jL+4sv83UE7AE
DU/v4O1uuF6CF5bs8/8eFZHoQWxWM4OH1/lEQaFfwFfoU5If/vtLfH61e6oy
FH/y2eQjc0oEVkt3VuhZsPqjsB4u2Bi6cZMvZ5TQ4+tzNSsBAQ7es/SAzOxX
68JYazJVq8J9WbTpdYYfC5BL58MGas0cIVvntpKF5EkybOwgOswygcfFJdRk
tKZ02p/w6Zyqh9P09WCmY48kooTJhnYsThZg+NpI2++Cx2sOpz5pkdN1ULfv
n1Q04RciS6PsQRq246xp17b+jc8w8+8xpn5sAn0p3MiCzjhbMaQjw4zbYTA8
WIEdmZenEXcGGnWH+GuQy6GBx0wllqklYFaaDM67U83Kmen4NaT5DqKRqG9f
HFrmmi+A850iD04IH5iNWvCjtbj23qtSrMnEOTGqNg5BQel7NapfhBKHoGDf
wmQ8VoIM6HcY3/MHo8lktWxcxL19OLfdcFbwKfg846z1J+Ib4y+Pq+aooFTc
Gd1mhILzKtKq8d+suTek2MtPlHC/Kw80t+FEz4cOMBAfL+w4mpnAc7kD3mon
Uk1Tqv1uSYhtFk8OT1HlNjFLo+DqFbQmFC6qfr0pFVc/YOdEVyQCSizsFszc
eO4Rpf2Z3FnIGj4k7KxaZdw8IOWDewk+nK1jQjzJQTVE+h7ZH7r1Y8FaxX0J
N/rlXysI0kgC6B3LEwg3me45W7fwb2Py9m30oRpNlfudBs9pBwM6hm0Iq2Vn
HukjIoOvufogrF4rH2fTRACwbNr0q2cEWhf+UEDdZ4T6c2/5qEEMsShkp8gK
cW6YPdNxaObIE1oXZY3uUNdKDjX2xqJttKU0sFNb5dbGpqkGa/MNwuzj3QWR
Z6ebKc4XzZAphAiFsaJne9OFfQvzySzy0swiYJBShj62fKR8UrnprF5AsUGb
xnP1y/CAksD5VutheEPjNyZevz++OUp2RyvjOR0RbrE0+3vQXyRf/t5QirNz
jkbkcu/88Vq+vWzT5VD/Y9W4dk+am6OW18zViwxRn20hS9zwiakEMra63qMM
OfIIuZpP7PFkMjaurBTZbElMh5c5S6KqyMXpcV0Kq81XZSbj7+17IKGPD6yv
AwkMEj+078UZDXofZwvI1J4OZ5hiprIqiKQQjC1LFXgPB7oo5IAcG7ReTMCm
BCUsBV6on9wlsVYYloTeEUtAlqzRFw6IZWZTJSzYqDcnlH8lR3PZahGM6LV/
+TK6S8go4FgXZYX5Skc8Fs+9MaGZC44kyJzyF51qJ0SBdI96cYAYweOjPryQ
6euBTcKfFQ57oFXwV7r3Ohgp6ebCvGgm3BVVGKdfLas4PGh0M8wPU1CDgmr3
czmxqhGiAeKJJ1/913avs6Xml7sm+djWqnQuCTOweqldIVHtc6y7GsDnx5+7
28VkTC3AgkbQnQ5z43TVFgQ40T9abssCw/oagUSqn3dnGcXeCKzdTZhnaKQt
aGyEv3+mCIqbyJZaNr73TX4zW0XE1gdokkMzmidnoe1Rj6Qt9gvKDvPWU8xh
DlSljpbl/1Uv5JmkJ3nX9Uxp3q6LURqCaMPBI/zmQu7i5ubO6xg2b7xLzlf/
aaW0cS+73jBbI8tkoTB4MKB3bAJMNJmPLhM0vbmyXuJ7qDvp5fcxSKw+8xUs
i5VHRHTtsBfUp+dF2VP0wTZlWxrs0J+6HnfQgepjKXTHqLMP/PWtNEmBKha5
W2Wi4+sTppkoLWaDNAxtV0NR98MmvUuI6mL2eJGkxszmtnI6Ok91ERUge8g2
0TyfV+vstgihggvBbA3CtW0v0BFfmGa6Zfah8NvpWz/8NnPYGPVu+muvwBIL
kAX0XXZ8mk33/M8bNuz87MRHmTPlhG32ROvx5ZvMokjfoUX+ngI0XLKWqJtj
tCUQLg2ZFsxSyI/Mgmbot3AgCQT2J2T/cZBIFb9bTlhtIxNdanm7zQJ5WTCW
CCNnOL6Jk8uG1W2rWizMLjKMAnJY0gFTZcidzq6eJ+j+lZLPyiYHSVkPTNy1
uN47Ls5zOziISxD6hxLyzaYQL+Jvc9eBNF00Yehvizau18xy8AtXgKCRJNgc
gV7FL/GuWOGSsFmNr+EwssbeHeGeVCLv910pP+I9KkY4vDByQn9pViK/xtJd
xpD8rRYO4GXWECe+sOisfyxr6B4k7369UKzZubSWSWVgQldspBr1JxEExCI0
j46qXEs/zyyNuoO2Uw91fkQz0MWfwoYsRXsl9wMofGQLKN6HNTP6RQ2cN6UH
1nrEk/WqB4iImIF2s9+X0mj/Dp7utSt8DsiFFWNMyeftfoUvbEkWMJLBANEH
9EumRzDnN02RtPyUroJJZPAVyT0BvJa04MRiKXAsgU9P75n75/5krGavmX7x
keyQFC+Gja88tYtV2fiEUDOLXnkXY5Njd+9Y49lszFY1InZLVDFwPhUmlGzu
PM0XUZhrRlaN1ELa5cLM/zJNREvfHv/ZYF901o3Tci3CwYR2B04aB384lpai
RwcxRPuf6/V9rUM0Xv8fKEuY0ALkTws3wNNKlUjAphVNI7tq1QGQ/tEQwp8d
zfg33EguxuQ5Dj+letCvu8Ac9iy5hoPpQVlwqbPGstMYOCP7HC+6NYdlf51P
h0QzBMc4mRu1qi4OqHybPkXIwiQwdSMVTft+M42KpnZhSkTmqeGXCr2evhgO
vjFBm9Azfa9CYvwaHJOHzS945xrfPRXUGcKI+IDLJ4lO2T7GkqPgsJ7qwwsC
APximlP72XYUEzc/uOFRxkRN4tWW/jVYVz2Avz/XHOsv1Airlx++fWegQHUi
jgBx6EOxhhuXLciFJYiwoWNIQ1v97puhFBBctpCTFUrtMLBV8AiDA31WZv7Q
E7USnHvpldjgz8/NMU0Ez+dIxc1daYtLg4ssVFCwKatBG2ThOWCYpCAzGmQx
YsWq4VG27jtYLH9Fdv16xBl+AGD1P/Wql+ozfx37Big8yqFL57QtfN3OYRhn
drV+BTSv3G9A63zMr2yNiwt3zPOczpZ8eFbzlqfdyNAr7xWgvvksgVPdpK44
C83E3vBnT6bxhAhl5C22hEerMHDA+IsrL0PhuJ5SSdBb0zBnqQmsWcedQbVv
xamqzHAUYM5lt3beHRITtdwBcY/lMn7pP3jUtovWv/p7j6scFk84uTMoFsDU
DQfu8YAgZdo/eDx1PnuaIaflNAZ9VO3zFmVXJAe9kPoCF2B6cF1ip5zzoAbt
UT6GDzXzmXo+hFHS5YenTXGYYfeBB34Vaa9is3QvJ/I0p7MFKEmE9/ziLDFA
eNCLJ/Tf4cGwAdWLphoT0KcTy4oBF7ZsTVS+nVxi+9pMcM4VbR2fi5lA8biO
ZCT0fhXD5kwoS1eZC3sHb2YedPAj1hwQLNT3A+ZuBAQU+dYe+5s5JziKbNm1
c6axL7dEeP1raaZNJB6pVn90W8JwDWTw2fPki5jV/+rAJOzeWWMfuQd3wGbD
Z+WwbDI//p1dGsp62KipVxfDabMC0Fd3nLG0l8CJ2n69vU2+7sXjykkK1LNy
8mf8Gzwo64SU89/51UUGvCWjYnOiXMlnT+rAmUo73neSHvbGbprPykQbQmLX
f0OaDkr/NxxHegC+9rNll9DwV1QK3xF687bGyeKMSS4NdVFTT+coUbCHj8v0
KWHMeHENsZAuiR8iFKdCZGvofp4X9l62SPJ+cXZZKfhTx7mYxROpJYBhYEAg
Ljd1vBJhKixCssCpGWvVj9yhTMcG+qB2w1167HPYnfooDXtZNrDOWqkyPwKE
aTatMqFE6WsfRpuNH6B1gtDsqbng6L7vZBkLd94rVIQI1hjJKwMr9wvxtgHb
EiYmWcUaXQnK875w31aCUU6lw57CB/cGPfB29mxqGMBNNp1tMOPCWPEkFuVm
437dTl/j1eKh3vKqodZoOneuhqkdDJ9zG2ec4JDUxhZN/KXjLeMFl0NoVkwa
eFU2hc5MqNV8JfYBXbl5Vpus4SRiNXATUyOikrltnq5yqs438WvxnK5hRsoB
pdkXhqVDZPSsVBAftuJVHcB8WcvwOUb02r5OsntIDBvja0TC7SCPpZZiMyaN
PeqsLYJbR1KGMU99DVjOn0nwBKAhV6KGuYuDoYPefqWaLtCtdj2PqCH+JL4w
3am9jFTsq20KmR/8yF3Ug7hsSY594tvzggcI+EtAvGFj2dsc7TcP4+JPeKPL
0R5NwzlFqNJdkAkz7UfiOCZu6afvQqAsdPMIPjB/LXdrXumgzLishXmmxgB8
aj6kfwKRG82qSFl0+Hpkcfy+MhsqjXh7Wn9HHitMUWMJ79K0YoTUz4VWDSgt
U/34PeeOnWj1RHdQ8e17ovLseTscUZ33OxLTZzI+xReIQrB0GDZU4uiOLi6c
wEZiQC+8V1Vz0fQafAXJm2WKPPyng+2toVHCSlhUF5AnSFIQjaj3VzpPlfLK
x0jt+EEZVxCI4s9RE4QoqyQblEhM7Zv3c54PzurIsjIL8ovnzO+A7R5SBzfS
u9/Oxcgm5oDYSV45hxcq8NuqrnsxY09wgXXtc7gQ0y7tfNK5CWFErrP782Ts
N+7TdYh269lh+b8K38sbVO767oPLhu6QCb0Ag2JArTuSjjp7M5K52ji8GMkE
kYGUxoGKMQWoKu2FDh0s4dFiqsxxq0ttHrfLSMyOVtwYOOwUTZIG0Ux1bU/K
JyfoHO6cpwR28aqppH8vusO5M7oo6xe/HNXBhAdHjNr4LHlbdL0u/r01jOyF
oT7ps5z5v4atanNc2upkc8V95aGcNjgVl8ftw+hBfLNJWOG2UaO2KhRg6+1L
Q43B8BteelcaBUCF6IfZ/CrgE99uBEQqi/EjRwG3DDbLQWixC5QARCvowwQ3
z39HQaN8Wre8nXPhdcX/QQDoADx6PXds8cYj7AsRxM6OG1ChbPRrsy1cXMDV
0z+/vpp5118V37Nroq3yPLGXbionhzXrHi8+yrOIKNIYOlgzBTZT/2qaQFw0
Z+HAewT8TrGeccSVzn3lkz6hwW/+LOmGV4e6m5D/vcUOrv1dkj8eyPlee2wC
BpimpjrKd66/yr7jDcnkOQxVraWuojf2niTqBG1/VEqB7MJ95GddmDDAse3s
fQqNfaWD3pGoGZemdGucRge9CY7yhdk+v+Z1gimSKGwbCJCKwSQ+pDHq7Ddq
ncDXtFRlTDZW5L/BXDAdJznfJ/vZXPxcVzyBkAo85PeLstbnruWtDhYRQUl/
1J9tp2QSPJ9J6c9nZv2DdxpYouq3O29Ww1REnweCoS8lmFvQ1Rq0C2ihm5bc
+CDwAhKSom1dNCPIaVMWWb1S91Cuh8vpo7gpKwgxuRtzN6rplxgpv4SAfAny
Lim6P8FqUDpXPKBZfDb4J9/uxYKodq0vZbqW2vDlyHbnqr02e1EXbegPxB7v
s/VR14FpvvaJ48hj/u2zDuOVijL238TjP32vURmE+4G/24OYxQyWoEWTjEya
dZz6AnjyQFwkExL95rOvZMeHRl8OuV/Jy5bjXOuFs6ypDHX1L3WBKifz0D7/
mte1X4z5+r8Lcj4Jd0VMf27TiyXoxkjZBTO/tbyMgJQb66L4r2Az13bmEHqe
ZXuPRzUUgyBaNQAR+gkHNv4mfeF2cZ/HFwkiy/zjBY9SzRsbtQWTnnhgdGLO
zUs+SdsUWF934qjuuzlhgAeFfPAmxHT7X4zl31tPrMZz6wfUf7AiyKktBvG+
KJINGjVh8QazB0KnyC7bL3dRKF+5L0Wp6jRwJIusgfRW4XrOXEmv5SyFa8RW
IPGwRLHE0KtnHppl5wMzL2LRGDZczNGt3THJbtg/Y9ViK5DucaSgHV1RhwH3
/0rPEKT5eYPM9mxTHxcNPpXA+e+fy4XFgRHjqkxjKyP6yn3CcmRj64KskvNB
Jx7bmM6UWPZF9d87WZxOtp6hf28eYidPhuvgg9MsSeJF6BP+k/lVMfcMgxHN
HkehmvN3uOya/h4tdQPtPXLYfE88GLiZxoMIlDjCs0Dy09nyBAtEYMcaBB4Q
0hjj7yC4c/NbbuUP6msLRI1rnQ2tOaqpKZpkav8RuxFtKjJbSCP6hYFWTvBt
+ZQh4/N9Ldel39AG2V14xD7Rj7l3wAI4q4M6EHkvRtXxgZdFcU99jWO2vQgo
tTptbxlZkufLneAhlngOSntuUZaFGM3rZ9ynLFbtTDdsOl13Oxgb8GmlIj/w
4y6gWXOvFPhw7cSLWwiDskXeXzkST0lHBhO9Cr1BNOnnbWTZ8DRscnWiy0bA
Ny6gLiPGTUqNdfP3k1a+4OzT+MmnCLdsfF+1Np3aNp1+LXG46U5al+EwC3Tl
pT6QIkN0UkXBW6WPK6ob+c1U+PTrV69eEuYQGZERzl9YMx0x1wwl8qm/e0Wn
K0ylu6UYDv1+JcEL1vdPByUtFbatukHS3J4BJCK/JufMS+A3LkHUDZllCnKK
3/uZEaj92ADPm7dLKNEQiQl8ZdHyWtC7jZmSTHGtsZl/yk+0v5T67IqiqQSV
76kUIzJOB4/UiA6CvfJILo1bne5JTv/2/MQD0gTVVdy/iwjcfEbNnYR6F8Sa
06/l0rHE8FUIY4kvd4ueAQmuQRd2ritptH7SVrtT96ya7cAi9Lk4x4JTmhBH
vEHrSbKit8zR9345Sic9bopvju2mvaxa9EPA9Eq2eZBJHPQcYz9ZdT8S1VNz
8tJ5mbWS5R7lQyPVUW5D/qt5im2sMJxKaF62xlZHTIe5jlltSgBsitnO5nvb
aa8e7nPQo/aKTw43Z6VCRsj7OmrrwkvKQZcT2EnUEqveeUVntGGcX0HGDizA
BKopfqAypUA1EjRK6S1Vx9RFYQt4AwfM6UmPEFLiFWyfiuGacbAthuZFBRQf
Fcl71p4m+uqaZ+35E72NkURzH6JamZ+TCCJ2GtuV8JQ+OuuBgD9ncQ1EOo32
Woy0vXUXvSiVrJU7DpiHPnyalwE+KbWWlEqcJHHjAfDKfVmp5ZYmTh4NNtAS
0I4jP3oFCc3YTa5nSPIKceFUFYerUCRqxo0J7EMqzMm0TpsLVKQrNP6RFg1+
VV2HupojZ/ODApQ9F2EPpjNKGoZtUxv315K7XL845c/Yt4b6NIBDd8g/0GMS
nJpJ3gwGl7ws66copdsHIfWph88oXI69bKkr/wT1aZZB9pEWhzOxDIKCDFrP
hsGHYB4E9UxH3y2wgd/Je2FRJlC/BpMSUw77yJuz5CLMALVTHnxRDsani2gy
yLsdSbcfmUm2KFx7JaA/QNA7i7A/tj8rRYWvLHBVF3iR0BF/tDSHUtlyHI5C
VxaI+qFr8rievRyEYQhbAMp+z/xyu1b63eTU424gbvIvdT/e12gGKTGs/l57
6D1JQiqAlapulugCppmSTZrbU9VqFVaN28VVwZhU/8LupNGMsDnHwMEHNUCh
3z+/TUE5CCc3gBQGDIhF4YgYnD13M1eiiOD4NXdG+WBEhcWxU8O7EuANfmZ9
S7vFyW5skZZh+mhERiaHHxx9dK2BglyM8tjLWyRDJkCLPPokur17wzu05cP7
Oz9Pbluokz6rUo0LhmijblJnm/vim/5M86hRR8OUjj+cU3yXdKDLg0PT/6Sj
Ff6jANUOPoubra6HNpYnxJa13s32+Hse0wEU+/+yGjM0FCbXrGvOtDrcuv5j
SEyC3BiGJamzOyrGp+tFk1BV2fdOzaOz2EBxU0LqvQvOpUAVwlx5TSmRm/4m
kCTEGArfsh2Xyh0rOL4QHFWpMWnKVWwKZ2xeKnVLqTgQY10AtdwjA9YJ9p40
ByXy4eHeIVGFm62bOfhsglaL3q35yC0/ZrBEq3OFaVPsvDnoM8g/KNQWf/2z
BxOij6hUG8KcX9Z7A7SCpaMJoj5aBP+yMYhst6Umbxhk8UNrjGDZpSY+9Uwk
AGj/775RcOklKgPGCgnNar+/Op7O5eQrDJop+q+7gs0eQt/ObI93Tj4fFSjs
mgbDwoPRp65+CpoXoyzZ7sCIWfeJTKWWhcyfJvjY4J++Eeox4fBP0JdrZcK7
Cn5Rc2zDuYyMu+Q+IxT39I5z+A5RnMOX0C9aUWAhsqnsFKZcg5I=

`pragma protect end_protected
