// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3CyEu15MVnWQ6KFP9JHm0mD+eroEAXjd0Q/b1y6RzEumlnO7uMzk7106VJsgCpHc
3sJHCVttMybzLwHtufP6mEpvDf3whlNwPA0sNAUqqbKVN7SV1qFD1/GdvcSC1aaY
xKeRnH8o3N2mjiC4e1dAg9iD8DuLt9ndyQ2Qkqqwp9w=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 3792 )
`pragma protect data_block
2TbbLsczkV1WyozI4rt6PolvZuGf4tqwfWQO6PfoQHTyPlnUtpqPqhXbjPkNzWVo
b6VJX1rGU6x6jKjZcYr3bMGbBG36Bz6ajTZKFa9qELA/NNPP17KZ/WhC9XKH96Ze
rtYHRWILr/W1rJnvmaN2x70uUw1aalqRI+m80j+NknESg3lCXxw7HJTTvVOxlwgb
lmwHZf/f4gf0IxzTrWXiLAM5s5uYiU5lakOXM1gDA9ozHWE++ZuUUQc/DE1dogJK
oh+yITl5MNuT2E9d4dWCHLhJ8VE9QnXSa+JU4tQn8Wt3aB/yhFnGXNLDLL3HADwS
1bfGmJEmIEmex28oFf7O5n3qmCsLot/42LfYJptLzM4VmLF3aneMC0Bl4dlaep9P
6l2TQekrs+VmkFRcBWyc4L5ktc1uMNmU+rN3q4vKUHjAcIlXdQ7nltPS++HjU1Ey
D8d+pRLJtwM06CulptSi5tJ4guLAlII3qYIOf4zenl64ak0E12BkH1yf02bREWXw
pncfoaNNjoPNVSMAYpjfVEF6gSCsKa0qfm0Fh+ZJDWCjepX86M4XQ7SiAx37bWi2
odABqoyuPdfUuIeCqhSJFSsOMOPpyY0Kx/unuFUi/NQEGlB6pgy1bT49pkA3nSGL
UJyfxXmDZJkXo5ybOEDcIjw+Z5IopfTF+67esPO4JdtT9xsxbeCr9SuEKucN4LXP
aleXlKhoRGbRx+V0rluGc/QuXexriVQEqMPaOZaDYrfREZ/HarYM3t7MP+GKCazK
R/fHbPUiZARSvpkzvf+lIfIOVsRpRCxRxVEDZ0vNOagGcHvcSVoXOLtu7kg+u7Bj
h2q8ea/YJlxHmeWKIeWm9UkKhWwuvBiC4Y8Rp8P+ABH26zjtdwS6fSODT9fDzHwg
hRy6N4A6wxiQOB1bE20djILDBbxk0dh/SaBHCeLkYW0foaaGEDTc2oRlybZDdDuD
u87hLz/mw6y51cMF6of8Xg5N7ZDTCmnX9F9oJrXi8hTaHvpMbgqHTPS4WM0YjhHx
OOw1l2PWMPEbjBOSmEkuU6D7Ea7Fo8ZT5XfNsTfmTPPJP7yxIdo0yezavbwQFVxX
K0npUuLJp2If0YH5oAjSi/oeJZkiraTVm9EulJ57CUM0dfIkUH13zAK/sitE4Yyr
2kWo3pSIB2rtshv1PC+Wh1Tstfjp03CFYGI1Ci9zxJdT6qWz3fR2YajInPxIcVQF
A8uwryFk3w6hR9sLALi9fvAJQ+YdjYV+FqnZCrR/pBcu5zy+wpYeWMXCKvEJaiuk
FA61xiIN+bcC21XZLvAVTqjknjGVHgYyMiOasHNR0/O33yr1wtJisykKWoklRR8Q
41hiNMxItPzDEBIf0I7uUIzdU3H6D8lxFfDQNuTnu397WIJ8LLpXyY3xkb6KJbiO
dXEcCL6esFox5Zcpd+puTlg7urPjIlfcEFtrOJ62o/ltE7e1gXKSsMBqx5kzdSmw
aHGZSP/NB8dIQSYlBZGK9L0Fer0no3LNOvQ6eHQG1tPtInm3PooifZk38uAVAxD1
DHgy2v2uSZlI0jBtLX42hFI6/A5yAdMvbI8paQ/Zkx/qaCD3NreUOHuJ42ry2d6v
JtrWkXysfY67+WaLG/ezAFsDtfdIE7mjjCZWmbJBmkB8KhxP3gy2OdmrIT6AeugT
pFCerMF0/6Fc31BrPJD/DzNVGL/9UYTqQfzVOBx4G9br9zpr+sYkyTVyS0oK3lF6
gjlPpYW+Xrpcmuii8eAG740aXoMOILi91XQcnwRdTXBGwnagY/PjnQUXxCyctVAG
XBSnl1eurMAPUAE7NbRomzjBtENQq5GgCE1nA4oQ73VgMEiIjfrW0SbhZ+acSLTd
kZ08CfNdE0wX/RYSuuWR2DIV+/j6wKXd6uIDnQQEbossT6aDVhrPbsM7wBdDU56m
M82Ex9nH9dAwK07o5/aDGmPJaFbxn/KU1RqfF3mf89fsNlH+RRr1GY5X/aYQeYbt
uL2GL72hjW9tK1aeC5Y7t3tsDLaln0IIHt6fub/fDyWJc9du8196ovrewceXDBji
ZJluGAnbIMA2kJ+FwwkRZsP1jZ5T9x180eAcLAFh3W0fLnT6x4I3x2HDsEg8dSoa
BR8yJIJp/mL6qhEKvw7QwLyxTKL+H3vJW9FGJuSRlIUng/Ao5zoEMe3t1iQyq+FT
ePdasZEkWyDnxlPEtHn10ok+fzzjW4nAogILuscSYbx6tAGo5k32hn1TN+ZRD8N/
eq0C+YvPFhilNuj6gGs1mibBfhIO8tKhMb4MQfxWaHWFrHJxkS3XxzqeMHQwmcMs
soLFA+fdiT0hOUJz1FcQ0HgtdNHizCNiiwrFDLkmPBFQVPwYD0YRTa4N5HO6Kc1V
AqDWyhuNpzwTh/ebk532cyFH2LMin230twXur1jn2uMVqxomFhgsLlHY8+u70+Tn
Wty9fXyTdE3wd+tg+nsjfH1aBQab/Af8b4GsJI0q+97EuT0d5ybGgBznI/fRJWWf
O41Yye7xZ6lWnII9/xe3M+URaJxOvdMmxd7NneVaHzhC1wznKwpPqPBHUhfCNzTj
9vQju9zhKaQFlB49/h/N7RZihvl2FRv5cp3UbsmsNTM+eYk642A2ucjTXCKa/7U3
xZ+oyUhLo8MIfOT2PjpKBnAND8yj7BThHJI0r0YI9myh0ntOU7HodHi1G5jJ76WN
Kwd9I+zNIs28rYE1s4ttfSP3y2iHdIG1qpmcwk4gTTYdRNip9ju9WrETdjKSFV7M
iS1aSD2yyGIO300J04QZpuxsNYrT6hhsslya4sEUW8/NYu9rjm59tXdWCV1362Rx
/xOPZCWu0MqXwkFpD0zKv3hvPbo576SlLsCCRy3ll6RtFrPnuY3LZKOCDVVIIWNL
EasF4cN4/3iqw7ArCc+z4raH0k4ors6+SP8SJvHaSnRH7wDQPFJa+MYx0YDlCsyt
g7k9iOTs1XKOPefvHqbLqQqVJGDKAd2HnSpQRRjoHhALambNjuUDXMoAPnl0Id2H
/IZ14ufqcFSouy1zYqWfbpfi97pCbTqClcwiVEnsA1t+3HWc4vJDsup478zN3yhf
AlfTx+dJ14IDfEiByqHvfr/Nvfde48zDJx3LrvLqhLi+BRftV8DFI37TpFPk0Okv
AkxXxz1iPqEyg8Z8skIdth3a48jvd402f5GG+Jxhu1l6NpJ/8aejhJX3FRzYt37S
GhEz7+0l0p1OgUu9gTOoJMYz+OWq5c5pKQsgTk+VEJuSDCoPDi8OllzdzPl/At9D
Fa+OIiaq+jtqUvEZzwPEX2f6mVOCmn9tkOUxVpXvL9eDVg4k8R/t+A/LU0r9zX2S
e8BKlr89lv3UIlRQW224pxGFqlIZVhDk/E7DQK0zI/+C5EfnUn8vKDdfRVRHsquA
JFRyF9f/JRtMtY6dchI6HVGUZRcJlDC0PUZJLMiy/peghSpZPPhUOo0oS4gWc6VO
4LZati4lwAZ8fQ2kD2PXGp1PjomxwL63/dNSyrFYm8lqUfUpD5rL8DDh4fqYySN9
HrZtStYe1Mq1u1rMW0uC7VLlDuVNn3T5J0lUQJ0WBnYjVBaoul3JRCsJT4jthTrA
HBmxOF3GHHgPzMJFU5N9zBu90b14q6TmS4BHzFUaSivl8B3tOh5IPgxrH/tfS1MR
J0Uw8KeQc/fBmEiycYF7LAwF47e5UizkO8CzW1byKvB3C7KmoWI8ASNyU9Og1pLk
pUeSeb2+ZkGTVyeKqZOrL5be5y2m0Z5dm6Fd2nHXmdZuRrX5WWXju4BPtvbKIS5U
q4LVp5HUnGODEVCeGduq6r+F96XWEy0MdTgxbvyPcs63mQt0stqowwkwvYap83t2
6infNJkuWSxb6a3a+bxQJBqgO8b74RGyBojKM42jJm2740dlmivayKAh/ZZS9L22
RiFG/nugv8mTOPrJFFijW1JRwXK86FmgEPznQ3PQUrjA7O8F3YLgrVfgmGin2UIU
yC60pk7bK/9cYdPR0u/jAGtKLh5loZpV+edpZSE+KL3FmhG9p4ZQE+i+/O43Sl9u
qgI1R+rrpyKmgSBFTJ+54HQ6YYBuiaOslc7SBoAPax+obrdyX+y3qhD23ilxJO0k
FFoQ3MC4nc7Dl7KsWX0HhnxUTiLe1QSO1EEiNPW82oMmcjyzAYfglSMfl23sVR7p
/lh2IqIghXGV4Dx8tb+4Q6GVylTr0pNupLBGWC8hxdXcTOqgNdVinPAu2ihJMD7s
M1mMGLku6X0zWsKTNd9cwyFC8i4K2UNVr9R+8rndqR22z4Z3cEXalCvkUqOBzTbm
Ig5Pwqdm1/XAj7FXvTjeG9bqog7KWkXFbG/hCnkzfHK2j9ojO/Q224lDl9G7OE6/
C1Mtz94z5RlyPRXCwMt4gs3q7FSe1JPgGnmHZe1YaACqzYuDx81YIq9teZqnzwZw
GTZpJFL5zi7ptt9HouGboAVag5V67A7upO4CB3pTyAgQMHbIX4lsu6U1A/XJKYCe
vdJriDZKGRlTnrdifn8Pk/v2uS0Gv4MAeCR4rOfMd45BaJWHu5gr8CSZ3SHPBu55
ZHTrbLGvOFWz7gnJzXAkl1MpRfCXc9yb23RM/7RepAJ6lFfNCAfc+nMWSq0wxNSf
ohEMZOX0C/r9+LJp4B8vzkw0NQ12tWpBfJeLSDCyYOfCwB4cEJmsntJrzkndxC4J
2qIEiMMSljUAOLJN2JrV7tLq9vQiUnU7GkKbrm9QmYiaUAijbw6Hg2JZg7FBPB17
DvfaFOUksipPIUqjnFUjnFFb9QG9YBRJO56Ui26CgIlhyCn2+fTcQp/Du9isdAQd
rUyyqMRUTlyIoH/RK8ej6ermigh8/lXo/QydX7Ot0q2+Kxxe3LYaffpBK7Zqy+CN
jstvaegXkzkTy3/IuTf8wgm+uyRrIzp5LoebkdiimFj7OxP/lu7aPjj0Erv24Py2
jOWAMXoOaAJ80Zim/gSbT/GEsJFjGogdwXb3TfhRYm+i1engIuJr+nPPx9y+bHg3
1pJe7Y9L/XZWoCmIV/iYk6zimnIbW568u2J9Ge9x7UvHPn7QQzXUM91We2X5MwXQ

`pragma protect end_protected
