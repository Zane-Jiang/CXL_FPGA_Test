// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DTQm5kINHKB8d9WHQBVp39je9Oi75HoI+kzwS7ZcleITgBlpoj4aC2esU5rv
FtqOa4jbLMJ8Tdq+5QeUsGkECGoyok5CQMWck6jm01qrPEcSUeqSMxfYIe9z
mRhDLIv+fIagJEbLCfJSrk/i+iHPZxZHaC5w83LLIyBkEGy991xtEDqZYYIJ
1PDF+BTWz6t3cnf+MV5XHADV12sVRQ3wv0bDDv1MD73Sc4zpCqBMXWDUV6aB
W2iTDuZFajUcFdFIj5/6BDfi3U4YwHJRu6Q+032/0igINwfdp0UeCUh8MNqK
EK2Qmryxo6+UnjHV9L0kfhNyCB0B0K3/DourHOXTAQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DKaHbRPeoC+VSfYAmV7VjG+BTGdEgGZX4L36Q2Vo9okMLoMS+SaoTyaJ19xp
6Pk7vC0BSqDft5VmNdHaOIahK6kjwjFa+TWg1SMvfhlfFGlh/cbBIHsvrYo1
CaSsGAwVLkMblD+6zQ8cGxA3E1mmJklFttjRZGixw5DAyf//3RHitwFz1Pnf
QuNZl6PF6zdnuEzOCpjtkvYPlSh75hmCopWYKU/O+epFYvQw0D1pyyxarCjJ
hZhkmQB7vJTn5BTUBCSRy9mHjWf8ZnacF6J/+2YSZGvylc87/9G1/floIIJ3
ntTw6p6uiBwP7ubAn6o4+jLc4wOVZBRHWpcXjiSYaw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EENEELP6AM9BrZjXYYaF0Gxd2OWBPpupLqQU/qqtBT/WKH7HPsgjSNFh+FfZ
ctVlHWkhrxa8/5nBLUibKN28cO/jefpfBEUmyOAXekQVJa0zqUPiZsr/s6tD
bzcC1I/nL+zilxITjHDLlE8PH4caa1LzLUKdc5xSp7V0X61FJnszO7IUxK7J
c0MNRLfOXhKv9lL1kEuFsfR9vshgRtQ0nuz8ymEJ6YwPLWQxwA0vEfBW7gvt
6Yfb7yjxB4YhwwQAjiOBqt/rvzPGXoB/N0mGmdaM/UK7grPdZ8Mi/XkaSC6K
j13xgIjpa1GZCgzTayEONwxUTUIQz2pwV6hToOw7pw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rdR64PCFMXcZGdvOrzFoh4NKdQS5qchmrnN00iGmHW+zQMyEfB47ySQDd8r4
91ckMSnU1uaxYsO1ZJ83etV7lOPCSKJkuBP1REHCzaTtAmfO1+djUPRLU5hQ
kO7ETmdsRrthbIq/p0bll1gmCLS0vxWxm8MR8DPP88i6wTUcOyA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pDOHFyBjjfNy1DHTt8mW05gswTdrjM9hYwGomhCVPTB1N6AKvYrhyXC777OZ
Qjz7cLJY6glz9ni7z061EHnCGm2g/A6hihIi+Coeke5v9SRaddvG6rFJio/M
ZKFjMuLFStPRfD8Ei/LUyXHRQh5/Iwub/djYPMUnYHjH98FksqG5vc8O2VlM
iee3mZw65AQGt0wAIJeO6sAI4wUykSX4aR6RtkYC90sJOVn1LHoLJMrpr6xS
cCATLHmAu0UV6GbVvwPvdpAfZgBmYEV0X9Lrtjmp90XA9SmpZ+7Nd82B3lDq
qecKNxWDbGYQGzMwLW7nKLoXFtfdzditAN6xs34+O5q05Jn/F2hwUFmZ25vm
Ky9oRfXwCRGMJsDNeJHFXfzShuR2gmlhkdzDOKwO1bwALrtiH5Nro7ZMJoeY
8ESj+HDw221GXIoGunCk7T4SwFDEe/QodHuq7p1Q9U9KU+wbQQZLSrxpRCQ2
GNsyFTykjMLvyLUJdAn2GPYhVx9hpLjY


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ClBoPqH2kmG1Ug2w/17Xje48ITBOatx5n4iIRvIC/p8qR0jAMMb4GgxerdvX
kZBZ86msJZC8V6JYgXTz3a/X3OsQcFavmW4x3lch72Svc0tmczL5mkWB6Tc+
PpIKjjA4+Xt0fyccM7ROENX6Hnjr65/Vvq1B/GNJMNV+Yim/Sbo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ixyBzS1/VyVmtXBzaN7eKi/y89UOAiXdfOb03l3N7SICDBO7Tu6iawpRkcDd
8Xqrmal4+PHKoWzm3lqspgn1JWTM2xZK4KeomrUhgVdawH3FEIj6zerUjXRR
isOBdneTcaIJOpJM7avES8OqJEBIWvebTq771xo7Z9VqwgxyYrw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1456)
`pragma protect data_block
C06XkEeXshVwkD3rj7/L0F95zkUpTRYYWoXgQF0k1tN7njgqJOY6P3Fsu2DK
HZgJk7ViX8OGyqscTB+RQxtU13f2lqp7DD2yF1EEUt7CFUn2NqdEJ94o3N+u
HFZ4oulOa8bNq+uFap9ohFFLlHILFkhxfTSIrfm53zHENHVyQRPQ/aPj9DGb
m8G7ZAzWp+m9y6Q/JSU8t77Z/XpeiAJ1geNIWPK6Al5aDOy8+mlfpHtHtgTt
h06FKsroKuH5UPqtCnE8fPaU7P+nNw+Wq1jMvhvwOJRXvnBQIcsvmKk62pxb
T59OoFO0afHaJ6+58EZO3q0zirMB3vQo2jQw8r7fh5OErl5eV7ixjV13U6ST
nMCQH+lxGptkD9YFDuEHziGFVcZ2xhaO3FF2JrUkeQIpkZkRok0De+W1busZ
8RIzhOrUD+JvOvfeaW+V+De1Dy6WN20ZkkTZXpyS1MOvBmnSPv6z2ncLBzlW
Sb3cSCXaGc1AoM8+KlA4085KxCeF/kPqFv8B3H3N2rpHahgVFFrqlBmOavdj
pi0sncgPjXa4q9/MinZLLfuuA3AWT43G2QOpNCf8fFhD5Ga6Qv3kpaO1XiLR
ENN51IWTJNypPhu+MzH8VxgJ5EcZkw57mVEFSQscDah6qm+/kZ8QFO7N+VYF
Wez8rT87tgGcikOBOg22KyB4Sm+W8V3/l6RbyHputz7gl+RCN7pJtZlhBZyD
paDd14CzLRcyBLWqCmJ0M4ZI+EmzSibaCCZ5BLoeePHTi1/JQwmZkng3JRsV
KQaFXJC8RjDSjje3H3CD35CcYMUCWdKp+jbU0wR6vj5ocZMNtEKdaiS8f9YL
rtpkFkxgzkJE884kxidZLv3cc6hrTGquIZrOq6/r482ygHi8YDygov+mftw9
ISepTRwJCh+H423hw1oK5TZiLHsCcOtvfZY4eSUHUZ7PCTHRGLFSDL2eFKx3
jFwNx8m0QepJh3TdnGMsrnCt8IB2SkMoHC/dCWXRyoRhufmL1/8SoxVP+AqH
3jnPCiixKJv7vFyU7N3q1pHufvBIbwaKGhFYxuI+7b5g0v0Vbsipie9eFDvi
tu6xmR6ZGbYqSQQDCCC2jaJqz3uy7RUr2bPRr02tINaFXnLL5kL9SHIAkpaV
0wTsUTijJqIxh4uottrZSuo8pPwS4DXCXsXmy+kd32Uk3/F5GS4IgMplhGm/
wYLLRYdMdEjw22VFJGy9jX1LbdJuXxxEQUXTL3asE+5PIyOz4JGy9CnplmGr
qOSBXER04qPSnQYXNyBMQvO+j8tFIoTvIOPqBgSh9VSQ5C1bJPoy9W6kBswD
P1f6PkIVucXQtBtBkg4o162yJUb/ZOLV0c7wUKOMz4jEcge+mgtgmUTDLLzN
HnYpAyXC5IMZLXrjOPhKurxZ7Krn1+VSuW3f0my2er56/h1oSWQRtQs/EMV4
NZ1eDFixnB5HvIXn07S7iSgtJEVSKnjMiAy5xdAvdR2dXRFOmCrXN27y06BQ
ec5PDibwkPck5diOtm1Rl0BrhttEylmUdbuWlbVvQvziMBi+fAesiKYn71H3
F3TKrSEKxOAcfH/zHgJkqe3fejpNeTFEQarbfcon7p99ztANk6MbXW33OzBV
soblF7hX5vcrXVRaDb0d1UcWyfoKG5z+OcsiIkHwO3K95pml0dkfZKDZlNjH
z8pip3KWOaupNvplVmo9iE4f5DXoaNQ13l3GxzpYn4crqiuf3C+B1ALOeICU
g/ZqyC3u2qWX5Z0IFI+GMje4mf4l+6lsvAfwopWlQ0aics0JmSf0wFKI6tXP
S/ksHDb0W70ykSq7/Xig6YyqzVZTR2SIVhJQmbgzUK+g9xdl6MnPsO2/Ps9W
ryUBETBfGQtM8wXsRqi6iW+q48ErWm5dLlj3rXnoBG90MVs/5hyj+cdq1D7b
FdS72Ru4fIMvLOql00dbsQ==

`pragma protect end_protected
