// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
g7pZWJmVFK5mb9j64OrJCFdod/8C87GpgYARUX5jwM9VHQ381waEzn63e6/v
/3D52LDFaqN2DQBdVa+Klpe/K0VhAe3V4/G65i/zPiVZHMI2fuwxSXGMW5Rf
3LfsgP0Nyb0BSR+8IG298j18n0zHicqLk1fx5BMSWekdbik3oYiyaCbw94Vj
kHWTYJSSMc6Vyv7BkW+zY50HFw2EvQNlQsd7+Q/NWHcoUqp1GB27hz7UQo9J
kL4OgNQOHVgGSezuaonLjb/HPexfsQpIkcyy0D7fLsFHZiywQIpwwf9ffhYg
U438Z2VVOIGSaYX2lIAbjXNpBeM76lsSSx1V9uu9WQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ani6JpXs4lbVOlqkEcyZC+co5Wi5+MEqaeev/3khkmri69GG9lLoLbnO+XC3
GktxeLY2XVWpAjw8AAtT34WCxWh56EfTI0f0+KBJdO3BtmOvS5AGaU8byHPr
gZu96ZrINr/qzRSrQzbOBpyFTJCN5PxwhnyBPlPA0v9eoXNqXN9GOPtOzuEj
CIKzVZhm4zKA7mFW/KU1X5JiWGNL0KTs9ZUhQVaRSNrEIZ2VhnOq6jR1mGJ8
QV1l/lssUFgIrlz7f0YknpQ5SCYCNyYWhRqz8+5iW0HtIAKuvAlN3gZaQ5Qc
+zEK+zuhtrL2RNeGGC/CYxL5le71CVhIKHW65bjxeA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
e4Y62NnSMaR6T2bpeTBTMw+e7SdnrdTxmocSj4BvaprPgWhO3r0V62pTSIXv
CB2serEkxhDukH0uocwNQmWYuaxA6wHuDXnbc73CG40L0oluIPH+TNqe7LJa
uJV2mtvaCv5X8/M1F8/27stO9HuIwFkdskTafSG0BA2dnZQnpDBpcUUiVV7s
PAqPGMvn2Gsc25TIbtAfa/vUPRzAY9qKkbzbDVe//QNs8v8AM2siaP5VJtCL
OaJe6LW+XO0RgX8fY45Iw1fhjJrk+90sEttit752Nl0DaOEJd41AASd7wkhY
zwRAb5CZ1vIy39MRA2UbvAyXO6ZuzxL3BtBoQmWRbw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PgGARdcFn0nAC5GbSUPIB8aGBHXFwfv9nGGtqHX04hnwOFiC1KYcepmdubKg
fJjgG/m1Oqs1KJJmgt6QytccJKmJrFhS76UdLTZwyUW6W6mZXQgPlKnFuHKR
MnMeWKLn3QsE2rBcn1CgzCu8vUO5xG2ml2bOnuYJ0Mf3jumHQCY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
E5uWmF26pxJn3fl6LGIUivc4OAK42cxgEfm68lWKZAXoEPXO+XKpApzhFOX8
70CeHJfMfjELRkcE3F0Oby8j6fBoA4xIpljVMGBAYiKpKRS1lgfjKbty2NTN
4p5Ytrj8vAtxdumDbeWT+vdXMS1q/q1JiKMsR7u/fly8lrDFgKIDxIaxTEDo
tt6dc5UGJVe4/eiV8DnERPpdZc9NqKT0/Fpv3sdCajMWAPv3LSjcBPoPJ22/
SvtnR7j1PD1TLFK87vD1VkSW4hpKQnuew4CKXjr8ObbRt5w9tJpcAPewjHUd
uszFK8KBljkSm+YadojGHnL3UtJk2l9ZhcfAsnrap3Jj/MwrsH80ikfiJ3XA
Hmwmws9X7nP0jHEev364jjD2BvaC8lX9ev1+PRoCfTiPKpFY8sgx6Uel1/Tt
+i/69ckiZuNZxgd1slDhu4RfrxW/aSlYFSjKLbzjNcINArB3ednAtF2F1eA9
z2oSzr2raUJf1bdUSdFqD6oAJOz4GpaZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tOXL+chLvLW9O4hVraHoSptJi+1m5QmYb624pRRkNezy1SHghfTnUgTG2LTv
V5Twusw2k2VQjI7M/0Fpao0gbruWZf1G8/isbeh8G5d4Taf3u3xWIAK4lAd7
Wr1N4ymoCquuFaHiCOjbbXj9/MDn22vunvBbKmAr97YFIxF9CQ0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cQsZ2Rk1uRxyiJJWYkn3f+kL17LHw7Plufw5uoxA1O03PD6oXgDqOwZrbnPQ
f7ae45amuDzHeeZUPhOQ3J/rR48WECm+ETzyxICoa5ErxSRNEJ8vshIDK3i6
/bLA4oa4OKsk/v1UnxuUhWptLWrRj77ncPM6mPZeFlH5DF+PGE0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 49536)
`pragma protect data_block
6ImesZ0QUgJxQNBDU0CgBGxq1UsNOBJKN6kxu7o4ycT+ELIN4Rawgg5nr+2+
w42mwSVZC7U1/pGJTyh0V6fsytEsNyXzvrsj+SufCDwghAfoAdJNDWeQdf6v
vpAUlRzT3nvuL2O3Gd+I9ts3Xve3icKzjfMMG1mXTaFDsBlvfAqdmM0ntlyo
WvK4S/Ahp8USlKR5L1ep+NPvTHcaXWQy1jsG/nFYjWlTmjwh2Vs3TE7aXgd3
aXvS/B4kd2mZB5cQFKDtcOAr8OMSzUCAKa2K8zHB2+HI2kOaXXeS7AMwV0eM
JcFdzduhPAecGRi41Qt3QCKAb/PXGlilycDF6DKlUghDKrUyYX+dTF9UJjfb
oBhWGemq2zE0Kn5dpzc6kAxzMRrRupkx5iXWS6qMSRaPzqpU7V8yXzytKq/5
ZGtwZNK2pNYJoCyMNCnPVC3u+NL/K+u2p+1PYMDQ94uvWnQNf2PltcE+uXGn
PvKAV4IOGSMM78yPHuUEBDlItcr3C9erp/FZ+49TcC41L6OGTcD6v6a/fNvB
PtnZAJp83H967I2/WOTMDJWdXFOrwGSVU20WyYuHtVJVED5b5cjHwJiK2enz
H+3XGnkfHFLAwqyzyCAaBBWtRnjuhdzg8hAdTETKU+hC96Um2nla2ayYIZcY
Fr7j0YSKiPVRJHvsD+i+VIifXtLULzVrRMagF/5TtUuIyRXInckRRB6gLbHT
4/ontBAEYBIUvYpz6E1sb2s2W4/7noYpARm5CHeDXuxdGX8AbQk4Co34MaBA
I394xb2AAzKIKAuEDwcp/N9dbyh2iUDvV7CuOexCfeRbWRyr0kl13fPIMcOA
mvj6qAYj+II/DtRcaE8ARr4b5u8HkYePAbldwpogi37CFkiU/lPbBasSJ56r
H+f9xEpIEtzihdA+/6ZGGLRxH5uqyIMWmsJPoryarI+bLLcRffxiVWYbFe9E
0H7gPTVcmrsLFULU+/wChxbi1hiyQAdjf9adgRCDthu5q5j3jq9Hk3j3AYt2
MbRFb+DIhErHFtB5C8pL6DImpyDhCFASp4h4u1CH9MYEyiF83xq9mi2tp/kT
dDF3wLWGoKkzp1YQQOsh2v/iDvHyPMexQQRi6EacaCiVfoz1Ru+zfzujCMQo
RUnTI+cFM86klgYHWfX0qR5/ey1z3Mlcvieguc4rWJmr/tH4LHn34Ma+UeCH
kL6E34/GkaNTA0wlbjLqhAT5hon2kRzQqXJFc/MyQ8WhE8XewBok/ZDCnIE3
Rs0evA3l3JO2DHaHGLQEH9+2IvAy6dXZcOmmlQX0LHIQZDC0BJ1ARbMd4ltY
l05FHzYmHsDgUEtEdBy9B8qJkKFKNkYa9kmmiw9nqvd2q7uvyo+58ileN6Ya
UREwc0O4PG7Ffm2av56Z+xULSxR5N1tKSArZNKXQzn3gagTelJroKByjKMg6
3ulPGpfxRFe03Bb0pwuxSgVFCXXuo5HheVmYW1RGKXOe11wJr5p3ebC2DX/b
/GcnyIh4F1eeGasW2pi9BsyrX60DluTM6c5O6dTt1Surd808ck9YM+1MvVd8
tyCgu8UeyF2kzTCttcHWt2hTzfqIiw+Rl5YSRz44k/g8IVvfZ4zfYohPSWz8
zD5XV9PGqxlP+xs4qBp0hZMbqmiinQJAg0wn5v7ozS4q2jl4nel9j5e39yGh
PZ8b8Yow5T0Veu5IQnl9Ia2RsIbWPWQd8Nmahy944sm+9SxCzkmaKB7CMbZ8
HUJiueQphqjwxxWpO5XHjMg08AuzsYq65alHlH69KSEGV9oB0IdlQcYosvxE
EsJfP4tXO0l3itaMabKjLnNnMFErVxL+NIFMkjLaoutL2L/NRr8zryjHsxQ0
g5yaeO8RA59aaadvP19H2chYUZJvlrZbfN5c8C+Sqolgtbk+U23awoj6DOrK
VqdMh0vTcvTV+GNPq5NlcOQ7JBt4/DOGC8J7qghcoPBeHX5JkSYGiE9SnIiD
8+j/eFbDdVMtrEWYkW+spC5XNHnn0U63ACUY8pQVxNqcgMXd4V6oZe2n6YhB
QDa0Ec1KnrwkOq0374N9b02QkDDxLBgfUd/hozTPbRFWjcqiw2SApqBVa0Bd
LFxSpDd8SrBivO+yVjROmAm0qcaMixoqlRFVOBwKAPtkSQM9eknVpU98fHyI
6qBSaDSZH9jojXBZgOxNmA4pUoyKCCaIQaindDXLFk5JvvQoZeQdGweTT9Gj
cfQkkyeYUJflMPV9ATOd2eD8hPZfODxcQ77G62syVSMr2UDB1lR3BpY3V4vs
UCRqMU/39wVwn1MZrjWjaROCDL8MjJiFv9MZIyvZusV98f5CC9mqK2j+jwNM
tQkmuLLQXSVFP8m6BW84BabCosrCv8vW++9IVYuhBNJKm4oapbR6O29SlIch
MQ6g20UT0fSwxXOm6Z0ZutJ7L1L5IkcB6D/M15GuWc9P4V6YAdPoxS1WwQur
yLzGv2Mzkw+lHa01lthaXE6jr1MTlFWWvWTpeVckzAZyn5Lgnz3VjbVcZqss
+X12t4607naTgtVfgWUY6l59qaKJTW4m97gsxQep/zpQfO+BjR0MJjM3nOTk
UYZCclNV1jFH4OVRNl5UQ2EhEwUOjSCRafUI+3mxCq49+9z5SfsPwdyqKbBU
mqRFWDFxZY9PR2DhlDDMe1Ik/hQYPHvM5jqOTeOgYXzrhpUrPZ/8gBt4cWEx
L8qYHT9caqufFmpUiluj9mgdtaKpcKRpLwKalhK5fLpZHbA0HEJ6ajz/xEB7
Jwuq31rQc7Ham8VcGj1RDZ2E12r9h6bkVrE+FPUpNMRLaWOSmVSIDkPHahP4
HrY0XaTtHmx939nNrdk7hWnAa9XFAnjEEX5HZpswarLUGsu6/4WGkkClHGAP
vF2eRDTF/EI5jLuicUfnb5rEO+jFZme2GZJuK8tYgK3je5Le/JpupTBLZfBC
256wvkHYzdVOV+g5bXC+n2miFDTZgjJZwWP75t2n35uAHWJyBXZJN6m7tVwA
aWc8q2JDhGMvAI9CtF1ob/ALRDJ60g7v0tsskjipZsKwdHuo7clqdi8Fq86a
Oj9xalxHWvTdkeAUNSiGNs5VjV4gSV8hddK+vMkvzrcZQSuR7Gg4Z41nVKK+
U4S8wc9kwUKm/I42tuUF7l7lPNoIQBMY2WTu7HGKzuxLfbqlO89zZM+ybtc+
dK14/B4f/BhAFCAcftn5h9xiwX6+gUlQSk3HGwFnJqkrkceB2fiff4hJ/LH2
hi1TLqiG95E4esHvancJLWnV7S6bmiuyuA13weSMYIVRLMW+zIDTVaUocTYf
ccd4FOMRgPtfuvs0aLXU+908a54En0r8PcExMq7aJfY5ayW/Q5jJDGFDOHSJ
QEEjs2YZKgQqvUVt6uU0X4pGvyMP6awtD1oK27PbSolRAvol3iFZvz7iF39k
+vt1M1fUqCD+AIzc9cqJTlSL4oZbNvzUp26FGnOmHbRlVEMsCbTlyZZkcTlX
hDO5IvKrKF/+r25+EBRey26kgtQX6IxB2C21GXy7IRFsT+QBQ+6exg1oadWZ
weVm8ntwcN8omsGAZYtgXXTQsQ7/rix8ubUsqLhssqFF3A/stEa9/zctoI9w
vGZeEda195aLbNSpEkeduyRC3NRShbK3/CxQT0Qeeb/9GXGNJLvNmBgkG0k6
v8NOEv9tTWuHStqYIX2TRPsjy86SdQ+GC/TCd6Mp0QMcHQSrTmwxLzd8axH7
LgydvRIeAj3kcCOAxEAEU7iLjX2ZhTvCf+UCpZCagBjPlmDDimuLxSDzoiRF
CvZ/rOfjvjMUlnynIL9hne1QdVGdCB6gJ/bAcXnsRiOq1LH878++N1Ozk9Fu
AMgDFIFNVMoFi/FTVvlhKiNgoniz3i54FK1rQbvVbde9mdY1LWwZIabwUilb
dJLHVlc2ivZg6T1He7CQWyRFU+UVl1XmiPrYN5SjzS0DOCcF643YrsL+mQF2
YXGmb1m64BYq2Ad4e4nu8QHIv9nd5oJnqGwGwJGghcxZS4F5kyq2uqNO32fw
AryOi0pbsOcQmK1ei7neM+mE1FaFr3Zn/6yh1zSImdFgkFMDBqkLbOQ2Ytvl
wPyPuYK7NMFpP9DJLlL93WhZtXeElniwDWN+Ra0hYLJLs3vk5vaOGC4LKi89
m8wZ2lpzDBK9Hyr3vWrMKNFjQWXVK77IssaQx0kQtBRYCTCRiVy+ge+3YfJd
yAMrFU3gDeLHdudqa2z2P0skiQJjQrga+wPFc8WYlKGmEXQ+fzwSLGZWvcym
T+zHN7zetyQ2/WnqnTp7ws7adqQ6izqHtSjx93wlTNjNsGLWO8iaXyC8Dodd
Sx2s2+ka7mnYQwdQIaNugIaccqNEAG44zvTlSZa3zEHXuR98C2zG+96YN00v
YW8sIOz6TW15xXbRl2CuOCxk4pX0UaDHss+5oiuNikpNBj1Uu7iTZGuIzn1b
Y9FrpJ6Q5KCjttVHMpb+ke6j/qhvEr1STKlSfniYHCs7q7kjxV6pl9fWYzY+
mxpWq13JJRl9UGdfbvj5U4fwcnaWnrmJAkz3ZKQFLvc1Mxf4qUTV/PypPwLf
oxpJ49oWHIHvtZwhSMVwPEXYKQEH23JnAWarGpK0A266Vz8QtvNN+TxDz/yM
Xu3H3suXNgoHL331das3n51WlQLzrHLwR18EfH8uoSuRKQEzeWYjLNguIEXO
uF55wrqVweUnKL3d2C0c80JlczAGq3rn3pLMGYVKAD5DYleWkVhlr2/l35C+
Rvp09tiOOeYFV/4rocPuCH6RlmYXgsoE6zsq4iDjVKDcuXs/PIjTZLI9wHk8
jT7VgDdcVv9DQMnACODPKoMr75doCM4DoaDGgEAQUX4Q5uSBVRKli0z4JOUZ
37saH5cQgu1pty9P9kqE0nSB2vEY2LDz0ijaBGDjtXvyGlNhqaBdGjVsDhsc
ttC4d4eL1ORjdoyf8JueQpcUsBu8gEtvjD1YPbbdU1/rfHl/1j2l6aAKk5nv
bqfehqLqIVON0B7OCfYHi+1RR/x+fSUtUlF+I3aHLqzeTd/bZHI4T4ht6lAg
vbQRL3xsDibMs7F2yMAq9p8+brz8ztoZJ6C0bwrMPfqKq5Nc+MxW0EiVUJrd
II7YaV7PXNOT9vlpf4JQhdvwr/Ss2/CXGqgHqUy3tp+FqcR8Nu1aPJ8nwbh1
+7NMXM9MKjlhp/nuiGH+vyouAjmwv/z/kZ7WNWSOgcstvBLFzhKONHYevX3X
IQxF1Gb3nK8CDIkTeNipXdBYk/Q2Fa4SPCk2nEM6TRce29z35/a758TL4duZ
ujX49d3ZtJXgvxWCJKZAzKhFcDtKRJWhUxahVPxwVFNTP+qXIKYTDY3jN+xO
LB1wniCGAYeqAV0Lll+VntpsTNy9Mr9S1a9i2syofNC/Qbf5q9sacSrGDavq
Q7PzisZotcuggo9qIRxfEpqFFuHW6tNDVVeNfpiO4/zL717dp1QBMW00bNaP
83ArxjpNGHAitNUcF3ISuGZAT4o4alwqZcqPAn/0NWdpXGuYzSr3H2BN0yZ+
oNVvyV8+zHlWLbiiovsJGPA0LwP3nKBozJS5dcQL6Wt5dHa/ISXLSabiAbo5
8hiSEfXdAX0r1U2x+dkHqmMYwx9SJMamGkzcxOoPhUZ5xXx+HS3mEoQJLqUl
0jmbvjXBPj4vBk5RWiHl1IzUQ9kY5wy43WFoBPAm5GEXB6Wm3XHCC4KBk+uP
Uc4oi6959un+kNPgYQQdwaakSq4L91hOswth3+vEdjTr5U2swytSMuzjbOhB
SvVaH1Hz+Ts0ReCG25wKa+OTOWvWpIut/YTDe0/OA6lHILRvp8XAbPDqPcOW
vrPQTfMtHY/DnL/U6o1H21kRIrlKz3MccuACMJalDiXihOPLvFylyWHH3qy0
dua/NuqY2j2tWdiO+9bhyGfm3ErVfsMTYxWalNkFDrraiu2qvuWsX5mHmA8b
W4mbD0V/c5XIpL3dGcSEYnkwc4FO6KMpa1pD6FAk+2DCVDS7Ept0oVaUkFsf
YXclKmdL2J0V+m4U7Os+P/7PibX1cTheH/9uwKVRy1cvr3wdGy9cTGIwVGt0
ujsBQKD1iwzza6OYUcRiu181VWZAT+ZBaNZK96psYq10ppzD7sV6gImt5H9D
VwYbJOsB7xCWf2az6LKC4hJMXB58mQVPDr5BTMf9XRwLMfdpxRNe34JRcc7b
Q/QwHFCqapVc8I5OcqJ2jrU1EGJlzMzrVY9+6fXPKujSishypxVgRj4snOk9
sYxFqFK2ORdGt6DN9HZtSiCEvD9ZVoLPTt+T8kbWIyBxvNE152+niz/qWG5N
OeNwyPZxxx8iS1iUO2L1YebQBGXIsfTvrSXzKriBp2ZhlR3qhBx2Nv7c58kI
FFqi0y3h+jgxtTfYYjh2UORiCGIceu26nv1F2NgW3ocu9o5hZpJMl3jqehtV
OHxU0XGdaO4lJJwtJKMpfE5R1RD78yJuIDZdMi2lWbN6LoRHI+S9SRogItJF
YNJ1R/gmBz63fWC8P5W1xhVfAgmAnGc1DH3+Fi3q/TsffSH6+YyrkkIfgxFk
KpApbmFbErbALnrOnW/b4sYCTV3/IqToCuzuF6JnaJe9hr6PO+L6SJgO8qnT
M7lQwckf4r6T8g/5HLNDIHN4orL4D7cOL+VT3vOAVC/TxRCTG8PFwaWbUAca
M7TJ2RLFTq7yfFURiO7PYiz/2rw7za9cfgG4fP4nnovIEGXBrZLh/6Xxjpik
jw6jFA8HztEs4QCmcJPcnatCUfy1E2nnwyqEhBuflyfDzsmbBNuyX6fZK2n9
WCH4Z1eRugo3Qt7dCkQ+L6V4UBQTlvrQ70bhm/NwnoL8Fz1cztSiLJywtYhJ
yA71maOUX045/32KFB2jJNvKzdnYNv5W9eaDcm5cPLMlKh1GrWh7d6/De2y2
1+M+CW7FGtodBvTLKFB2HvAF3mQCpgwwITqgl3juf6m/XZ23j97E9rJAMkie
n/0IJ/78M79Y/oGaRPndWkOgQPktztZYY1supvBkmLS+SSzud90gNKcWPCVY
iM7Y+IS9CaXYZIVkdPONqs8i2nTu82uRy6JOl/FXuCPqquqhC7t7Bgl8dW+n
TCYv7kWGK8HDqfMvqmMRn4ef+TbixhPa2AeeVzKJnQsSHDEEllBwcgcqaZOc
uBtnV/nQRUNg/VM5Y6H0lHs8Y3OlatmE5JAnLX5iu2k3mE71lHngETjHOkhT
RqU5MXTG/mUsb6BD2ew/aZp13paTP/jDYvLHEqBSy5h9MaTWEKe8pKz2foce
uEBMeyC1Mk/E4UqW/Ca3YXrPG92qz9a4Mx5o40hC79bVjGdXINXyYbULEjDs
vJLUb2tZvjpNnL+0jxQd/WOWb/fFLCMSrGZP3yg/YdVka2TZ3Noxl+NqLXP2
qgCKDl8qQmwrC2t9aFtn4vQFkQNtrzyiODfXRwpeOt5Um60RVZKMpdCh9GDA
L88VELV/Uc/1DVOWsQJ2kMIheMfnWsLJk0spUSxSWA5U3e3b2iMhBm4GTE6o
9av0es1tyG+8REiWrqJzpQziGkB+vKLV/bJ2NVCuK+V3K9GMMgmxPJToIqo8
UWpVENEqLE50wzhYpqGX6onjL4Tj70ibX2rPftwJOeVEa7XsWOj4GSSOoUCo
W3QqXwDTYo0NKM24iDshRUUt899TMwgaww/3eevJmE4OaoP51yVfyB/eU/aQ
cpGXjz2tul+8upp/YfEihywsG2p+A+GlhyquZzE4cWGsGvyTZ3D/0zLy2SSI
XPlFYx0k2MVrXPnest+Y+8lUIbiVrOSmUqZH2cCj3HFQwbtV1w8+lT2iHsiD
Pid5zMAzFkhYNbukhFmkGYdTrd7WPXHkdUVyS05jLEr9EIO9IHBivOU4VYQu
DSdG9yoFXmCNpVzYu1IuffzyveH3VO+VQOlsqOWSxkr7rpyAwQ3njYr0lfqg
tM8re+DDkIFP/1cuakkFjrAcDV1h+em6n711JefGawvpQSiVokMJtMAn9bPR
okbK2uzit5LF8foSE3+AnCCDno+txnWh8y/7fxpVBud005uyJ3qmDu4zDhso
g27vfJRKAx3PyEpylVOC/cYi9D5FvwB6LxsPiUAzOlNIB6L8G2t+CZw7hIAE
08+hUB+lIs4JIwPiwfJj9aZEOEPHsZzuDma+hnikl70DEBOBu7EF/GGliQA+
8NRzPVQqLlvZsbwwoMXrM9IMbwiTPznr0HVkJkrgPBAO3S9M2yFU4RPmmGh3
Zh6EejDSrCti+2uGOHOWJ4XsiPSKmyrUZTTEmEgoywlSYinKgHCwllY/LDVn
czu2QO7ePQzGx+q8848r+XwMS+BiwImozv4QdZ0hRvHlsg9Kf6dXQHX5yHyk
lbJP8h1N/rtLDk+P8GbN2i+CjFwN3a/gy05uAR4RL5Gqqq2lCRy00nKfCbjS
zbSAtoSYyI0QsXz+84BZIhnD0DF0KU5FI35FY8X3mCLxghf4p0ZFDc47jyqQ
3XieMISYlFcrsoVyaKgPMP3SednvCdDFE6casqmWf+FUk3RdBFJyu28QPrhs
7vRTGQFukn7VW4km8rvkDSnM+rTHqjkWkxhhZ5XMRLtwYr8sZt3GGP5CJXJD
aSKOaMtZbCjFY1RqfiR+Qvb/++Y4ahUDD4I4fLasQyiynmAGpd5rHP+pcmbl
erUkXb7JAll7Bwj2u4ZTBhqE3OjuCFfqGSchFo1VC2Zgb5OeGt7+dLrmmK7G
B65/J3f+yyiH3i5KXi9O94fQnm3VGLbpQXk99bSEGNnyABVzwmnzDdfzVoe5
QtL2KF4TcQ+cd/c5uqCj5OkPvFWf3q8t1h1Wr9n78nud+hzd0hrREL7w631F
iosaPICqKPHFnp6MSYkY8AdWo4p1sgSma59MdJj2Nrb1uQ9rA9ZU3mzIDEO2
T6tERBdvp3bjHZEgCZtmkYPckqRaANabGTdM1WSD6dMGTSwZed6P7dJ5jeS0
pHpKVc++cpFlotEUAaERKyHCYXGDrHTTcsXTyPSCwi+REahQCMuLLZj8xcj+
kQf1sSqihNmqLV+H66MOavC08/ioOyTB/MrvOgJAqCE4BgpI977n99wIwghP
DVMg3x7zSVxaQFmUefhikyuQlXPsFpyxM0d7CJ84nHiYYS2eIC3Vh3A4zhON
9OP9yoOXDMYu7qNl2+arHmQHyPkhKFzqOk/nco+lfiGzIOZk9wPa/wiLSA6g
cTb5+vpRZDdWLKPLForgU+rLxERrR1NHeU0w7UB6gOoULdkF1i4NyhgQd8So
6q4ogwtsvKXmjLR7DkiuMuK7+Zz+qsMZmoKCcqtB47h/hIjT4cxCtTAS9hKj
gzZJ8PmQeuQbD4qK3SDV1ss+CjiANrvIkB1imuK0tSdggyFhNFEJ3j6MpwAN
Tq5aY8NtmHcsHtwOG+kqC8LgpcYIFb47uh9KsPfMuTLXsoyoAri9WLMH2T+N
ucaLdYF9SbZmxqjNSBBBeXvAh8ie+R1Bf65hZt6ikjvyGJCD6XX54VUWlhC1
lkPr64K8maN3y9QGppMuxMtmLBkvEIzdhW3ECSxceh1SocFMxSpZHthwzIh3
aS2rkDEdHksEolcg3pupGaNpemtfBC/p5kv9lzVI35mXr3v8JMajVCe1+mm0
2Sx23YqZmOM58qZZyrdGvQ1bGBrBI5xDGXgky+MFTof+Am6KN/6yNrULriUe
fgQSJ2vQswrOHXZ7jRlwddWaMec2b+ecOflMSo6SkDcujYx58ZiUdhLxQ7/R
z/dza4PlEwqfJSg3/qHObYRw6uzEL3UfOyXUBcngeVkdJ+4lp/lif2dNJnqR
t9loxpiNY4PufCW04JnHhim8CB+rVwzcIlWXY1UnR+smZCeHHU7eJcVnKjSD
8Pt5RydnZMNb83n+uRnnKmAw4ghNd4VH4R6KugtaBbuGCvxGbBthQ7C1th0D
/8ntQt87DgqBzejmch+W7wDFQQ4w25u6uepi7Rhsty9fpObalb/TrLse2eHg
t3Ym6yMXW9xi1nfdVRNpsDTo/IHTUPcYK/oz1CPYdhAq+c+WQ+NDOTrf8MTW
Uw7UUDkq20bOJcbDFABfxT0ZFDxAypeLS6d/zaBubsIih6LxRTntHx2zSW5G
2HIUPWJAajPEHG36qcdju+L5MhgluMyOlAbHlYfg7hRKdqSU/1N4VFcJKQRD
DUkF9eDEBkTUalCZEIiEhJmq41aaASAq5fI5EWeC6QfAXjqH/GIC8aWRVZ/G
/+zVwXsPCk8wfr52aiudb1ppCbGhsw0NLEBI7/EmW7ElAcQDF702o6KAfvQC
4+xOFXkX+nSrMA3rS1Vlv7gb7J+0J8nAoC/jYaz4jndunvLv95fBUJsUo/2F
AYRgM86zkeA6jgEOhD1aEq/Y/GHoHTlWnYjmnJzIOjF6Gm4gK3dDVPxy4QRJ
YxZ8HBxBnqJz4UsVEx5DBnesqtb1bBLiSoM6Vn3mbc6zfCdb4LsWI/5Ued9P
LNB3hyA92Mv2hEniTNfXMZYU1s/BrshtYzweHKu4kOl9KxNDSgSuCie1ZqNV
6ZmEXFjCdyN7639iSq/lWrBae6+y7rOozWxxqBgFfWkg7zWtwOAFacXi5vww
7trtxLHvSCbM/jUUvkKrhVB+SzdKeF6d7N8KAisS0P/Va+CDhd7PC99qRX2g
I+HJoQ90BmwmbY/uNN7HurQiWJepicZeB0EvGbwivUsKOJjUVIMYc06sPoNc
f9fOa1vmbeCHEK97dRMgBZyWAJ4nxn8h8e0Lk5z1NPgboD7b5HMuv0ctUeu3
zdvDHuhFNX6I6NPPLy7RtuLZOKPbKCip+7BOKaifx7ZLIr+EQN9OVlTBsiHc
cmOsKLeCg2bDo+ylB6Dr81qKmiA01SJKvAyZk76vc4du3igx+U+yrJgmrJXi
fgxMdSLk5+sysrgVHlUXQdXPBWwZMAZaD7DonV4iA77EGJPXmm4maiPOgcCQ
xzLkyQQyIiYd2ShsxkGvFdidhki6g7ru/wQYOZu+rIJhn/rTwKT5DZPYcZL/
fVm75Q76zACJx9htkaeaMNB9uVLbNgfCeD6H6RTdfUjhTQq+H2BQkNoOwbN6
w+4fRv8BCiNyCTthiq3gVLktzcjME7yffew8CeshyHcBFhXAAHAUjsW3bXRu
otSbyvxeoOrlUBR2LBY5Mx/GaTU4aQJ4I3TOovLAey3HXmtDRtuqtXY5emu9
nAkmdDgRLDb2iagjtRBEmBffs+tASTYUgWjkxRBc1e2kiw4WurCzoVPeSW5b
oWyIiTkwOtaqz3AcHtKnTJN8/SezD9kyARMyWDtbTjBVvI9C0eET1NhA7KEj
ds735UlE+x8FD2OL61E9tAwnA40XFbsyQ0JX2cl17VNbz6SHKafpTnaECput
b4oVjYqePpWwyhkB7ZeALjADK+sYewhvHiDGCfdCi3ck9fL+dUYXpSS644O7
F4ppP9XFL6SWfAER3xuPDm6b0w6mSKX+vjMdh3ksEJUJf4dgGFjj2cIwaoTi
NOf4FomzPZuZ4XEU1qrIuohkMVP7csmTwf5K+6dV4Ef3uPr2fMjW1zOzTEK5
PsAqf4LCN4SbypBnBXyvsFHbrpzcalR6ZVxYexckAPkubagxzVfvRDaBmbAl
UfWq4X92RNYcfUlPWWgh5QU9T/W5oT8bdsTnKPTCflndrEsQXBXRDexeqYtZ
vulACgm8ej4Lgjy0QK0xuYQhAk5FBKgVR9J3VIcCq7PK4TkDpSut0JlgvBQJ
jlx/HsK/fUHLLWASHTImusYDWoszxkj+L4cBiM0Q0P4XnmvRK1xVcxDFsP9e
QkbrU0gIHb/Ze7zhfihlFc6JsNZOLL2XKiGCB4fD96bPGNvpX2SwQEQa5G5S
m2an9uDfEAm8FR5uVi2ijgWuCX0szps3nY9whGH0jzZv+1O2MVmhAV211sue
wj6f2A//rP3c1WEvuPkROqX+rwMkYaMifn0snJayQ4RrQLCwm4/ZslidLnB1
iiZgnSvN5N7qhZbqkyRxWlCwHj5KCciJjc37V9Zs6b4ZiQ/kuO4+FJ9TPGYc
cVJajZBk0WKtNZV1ezsL6k26KFwEZh9JRvrPCPDPEOxuErlCRkNPh4U35e95
RcNayCqbW1WEeXi5QdtECZktPArLuSyG6Fkssk08dyCqxZ5w50L1MKBDL4iz
BRdRX1/gY19gkirXfY9UOGJIsSnoCbcqtUssIwqhzntIdikEFCATEkPmE+DU
NmpiKLrgMcvJ2nsGbxU5ly/ejACSgX8MTD2U89Html30DhMd9m59c2v8Px1V
1OrpB9kiJXzVN0WkPN5UG/gxZVNlihbSisqdAH+oOrwhqDszW2dgSHqVUvBr
xCadqqIo4tv4EUl0tG34IfKGlo9a52yv00nobbyF7gXgarWuMXyPiUx6vfGL
QuSyRt3r2TUW0zEp4lIWcT65/vlqFl1+aiIDSBIt4z6t4Dx6BkSeFMsnF5oP
MlhkkWAXW3O8esZ1hJKFX1ehibicvtRAEwMJnVw09Qhws/hbzkPppmwfiyDR
JfWJLrPoXhov5C7Sg+XKcKi2PGH1HlqeBxk6FFZfWuJa6w/0H2oNS5B+p/LH
dlJzxBp1JahDxw6oAhyh4O2rHbndkGJzItWX8JWKqihYRzT53O9lQHPaaQst
W8rXHLScC0PudtxzvGc+oVRYcshgS48ouE0q9ejJCwQEel5HiFNp7TwpjFUe
0r7ziXMtfcIpBwkIeZY6hR3obuyPnkWcvRGu6iYG8H5zr/PUxwdP9jioILbi
i6GLsPow5CBpLrwuuRtXLxIY23h9IKWAiBYRN2qagiHREg7M0XVBi7LHnIUa
mQDGIvvEJ/+bjtM/8gk0udAeIDTm8B0OdPNMSwGMr8vqswnfiSNDc01MySEU
Fm4FIsUasiiRnX0fdLPkFotC/rmTqkzuNEMcFdsLREE3oXlRyv/pnW58QIrL
gKvJQph/d+9qrqmqWslrCeF3veB3BmmOMxUEHi09xXQ05kPtx6oBFxKVHuxD
8Ufsg0ZLrE9d0A1sbSiCVO1esFZb9Lm9dYZWrE8JTNz2FQ9jbZyxmDWjCRaI
13NC/IHRTZ59JGTQD2Z23/yem+sf8bFbfqavBmFYYzWxIqqyiDdZAkZVmmr/
4uQpL3Uuu7+kKcfp9DJc444XGpkFont+TyBz+Q4oH8YcU2FOJ5+srBs3FV+X
rt5/fUFhQCAk1OK2cKuy1Ee3UHvUCtuAk2hEBL6rKyq6jYJV1wEwb9GnCfLw
C+0c989sm4qf3gmewcFXecqzk04XrzvKnSyaeXjrVmbmEVAlX2E5+ivAfUMl
PJgQC1lnqS72qqcA/mkiFhNJuyXq+rRAuULprnNjaNLq8BzN5y3f/dNqgrox
AVZqP0osNpjUweczxjRlXn3N/DypTJpY8ZBW/toDmkEDkJ/euhC73e3fa81r
s5NAYzmRovCDT0JkDOlWayEUmw649p+qGkJAmQE8jjkUVR3VyZH0qgZaadaN
05WhMH4kAl0kdjt9Y8XqioAbzqdNEzH7noDWP1EWkBHIr2KJBiqdQ8dM2o9R
Oeo/I2lksTeGJpJXOc0/c9+NSUgl/GfBwq+oIz3NOyieJqbvmNzoDMGN9SnL
X+UqqjgcTjpeuqh+IZy7JjpMkEi1XZs2DEH7IFbRFiFy68l9LjIz+EFXgVPc
aIw2qCTDSDsHlY/XjRvvmx0WYael8Ieo3j0eztKkShPYDG5nmSHl6dBT2nZM
ut1ZHPWldwTpRyU0Bu0tgDyjjiIFtHxoU49M9qKyq+INTNVsbWc0yRWvD1Zi
oq9rJjDFZsU7wM5vTKZH4HL+0pMH/HqhK8mn+hkowmSZ37Sgxr7mbHwlHYVn
Raqe2dyuGhwAtr5Uj7ddAygGbU0/n9Gxy6BbsjnixKe38DlYQpueIOTAPHnF
y9y+bsK+fA2uAY6fn7gdzwaP4DCjSjnyLcKvVxfd0JWYqtO/SQHnr3cHljWi
85rVcclVxdr23NHy2I+D/oYTu1xcwdtVjoNRUup8GHc+GQhY+/oZzi5lQY9v
9H5OyMxePB1XILMytIh1Ku2XDI8NbcIVmhWn+OCNlTP/1Q/O7NrKic/xmoI7
S5ua8zKEjN44SOFU9RWOWzdUqqKWlJ7jV3jbJX/oKlFaEMABEnGXn7hS1ojN
eJzGTg3yT7CP56/VhdoSWafjgBhqxy4sx6LFrYXAMucExwM54tM3f/DuNsTN
82T/IJliZ5wEfcXT1SQmd2lf42+g+YRrWlmAM6C5KGgtmXuIw4yz+luvLV91
TcWO9WUdWJfHoOwEe4ZGB9rpGQF96rr1VlzlOG1Q+P4MZujlhqLZIxV2ppSF
OOqq3cbXlP3I/JlcWQStwE5u6lAfot6UjETwc/jh5Fgeeofx4B3dZX+T3rzv
KS/yc1UCpW3PjPAW63FnZW76Ld5aHrTWWYK7zjbtufS9H+bd5rgH/AVu11/N
HfAV9T5n56zrO1A39RdI5ijobeKJbS5T1+0c+HE4/RH4nkKv9qNSp6DAAjaJ
P2VLdWIQZN02FaSVq7NvtDL9zU7qBqphuRqcNLmtph20atlzlLQbmJSL3PRR
PKsrtA45sfgd13i55Nj35Vb1ICfBay8QdDM4xPfZ1wGcak7EtOAgnyXby4V5
BHOOqLDDIl3O8Vv6vwnn6yija0xtICD1Em7NDJUSxA6vaNzgSqFLzNT9EYB2
n+QxZ2TKNwZjG4ESid/qo53kHF7fpi8Od+60QOfYNp5QyArp0iqFepqWxnyz
nWPopo92JxE2nT0cnhwhbac3MgUUzO0vzSJnxJsrNPJwZ/4Pp1+uuHb9LmVq
Ia3U9kUhv81xelb9wnz0sOhy9Lvj9Q5T/PSkxpaTefrYBgDP5s3YpFgYfiuH
KtqNy3LKRe78/H+TfgAuuqNptBRV2WMFlOw1ATOVkWhzEYU9QUktVLpu8S7O
wkXHfzXZ3mU+IrtnC397XtJCS+a3q5nh/40lbvOeHpyk5cd7b4TSsAWuBxGA
3pF2G7+HTYpsikUyXhrl1KnOZBw2ZeVqcxU+WDXwmqYATXkz1q4bbzq6lHU8
TebCu97hXdlhPXUdKRADifFMVnp4DFmTBYEpaZznn8kzOZXLh7ashoRl2oki
040ebJOBRdOMt7W6PwCg5YTr5EdMS/GB8SjvDRSUzWyAEtQChdiY7v73GtTD
LF3dzQvpI02rOdEvP8S3Y5nDTdE8uN9aHBKyswTatGCZT+FDtEzwZr8xxHCl
0+YWu+/vmg1AeOADtMo2hG21mZbcl4Z18O7Ct0A6oQ8Qvfw1p0nb58XfjMsU
nvkJqVEpo5nOyfeOxditks8u/xYITn9KWqcssTQaKNyLmPDfe6VOdLcvIHTh
Hprcw1RVH2X1GRvVCKpcxHCWU462tM3pwyhoiw8kRUdEIzyUmHaWesB2CnJG
TbkDSFcADu77TAowCQZRy7kq9gOrPIjc/emW0ho56dA+raCJKwSRxcBoXB3e
NOiN0C0eBSEs/1Qzj2MmO9PURaRhaM61RoUqOfbPxJcmGyyj7Dr+HNaPyyPm
1YFb7XD+m9pxEOX9gtaMcDmHYTb3CCcp3jTWRCDiG1yo70lUvQm9AGUu83QU
9MHi/e29yYw/Dgaj64vjCtMaGWxf66XQk/AXJhscHwoxf47IKgFwsWRJAjUx
it/ItVS/TeiI56baxuvrNcCGOvi/r33bO7+gd2qAOOlETWPsljYg3JHGLexY
JKUzlg6AnVcnGJGA+IeXCkPodrR5X4JFT+ZUzwZPh5BvU3hnrTH8x9Cr9vPu
4b21mNBi0jAzvAQeppBJPz0G0sduYv3ml863dk2pjsoQTu84XPIVfaoQnqJd
zgZJ40k+QzDCuDZIP1CBRVO82b/qgVtzSk5mxpfFyfgU/JLIm1W0Hf12K4hZ
Wiz88Ygv0xGcXlsJSO99flDYDJ0ii0BRapBAyyBSxUASRveg43Hc92GLsIAv
K3vrLZ+RsUdULMRZDsjc8tt9034KRiwE57753ZPUKPNpk14Pcq0fh/MNbNIf
b66datO+PlkqNjKnU0x1vQXdbejD/TXxSYaVnX3O2S/7a25HrljUarQuxzLe
CJS2uINhNyhefHGITH0PrNmyNDPDyYwyD6+PTHVBrAlq6mWw1hillV/epIrX
8Cfqjh1HAXy1p/BAl5MpWkOOULFLWMyrL8TZdKQjNt2RAWf2QNJzrQJjUhvT
sgZMAWIsg4hspF/6vI15vE2Mf7ewk+9cT6s/9udFMXSEnDxNv53+yaQjoqdb
waAe7OEAJhQEAnPmegrgGUPCOR/btMjRMeUhWX/jHCJrjTvG+TXUGz4Vnvfq
LRjJyZeuoIXT5VvIb9n+xQnTbUwRINlAA++Q41KaqAkMIkItDk90jw7a07MM
ZrZNYHcJ4AXHWx8izbnJDeLO/8R0EeQaf8d8edWdkX2GG80fqm57iyzSixZx
50/QFkYtzhY79Iel0RC7RmFP/t7VWGQDQBLEd9s/On96SQnmV+7RuQdfeJB+
aioMTrSRFvKXPqdAtWwPfM5GERJkDw0/j6wFz+IgthwSE/1OJtnOXOp85JW/
rUaarcRnUvDoKzLxeENWl71ybD6m1sZLLfrDryTJree/q/agmhxATEvtpTBG
XyNtsv9uRy6gax/RzjAiwKsQ1WCkx0IMlbzpwMsDd1LH90KVto856QX9zRHc
xqFM7nm7eCQ0cmNn3cOWOXskExOsjpURl8bXlH9w6nKwGgG7totxEFncA5fQ
jwvQ9beDW1uy87N6aq2afBKy+8MttH+bfgBt9+I+V3vjjU9N/jptlZok6GW2
pM/ggMVLbZNc6Nuv87mfmyjgQdXMgO3qQ8DmFHOppdKVimycfBP+C14gf5WT
VQfwHT1TYPpuTumEHF8VqPr4g8otYQs5vkjMJlbLcXtHMLVZ2S8jStgzHJr0
mTSGZe7m7z/3Pbp/WFu8L9qYbr9qBv1ATArBqJAwK6HezAncLIOswGgfO3C2
40P3f0E4n2/9mWEabnk9YNJ5pHNrIFyj9af+WSR7qehKW3yMQOz28CFSaA+k
He9iuyaLKn9nckL237oUI7gXJd54A4+v8prtJvad4b3el2JKPw4mvW9RIWJe
6BSyispHQPR1eifVDhFhIL9pf0Zz1nZVdE+2ZlryzDipLOoETOkGECEt37c+
hzZd7l/+/uPHrJekWVi4qy35892Y6m66n4Lfaqj8U77qGIDxs0PWlI6jyEvc
+meypRLye2S8iog5pnOpzUYAoZu8+QijcCSmxjZ16VRUprOas6xeu7gJq06B
RP/eCg62pIwDrNLUgYA2fFa8C92uBTmQGYbmX8la+BleG+G8LBMEZdTd11dB
7MZz9+pYAnSNbVSxKOaNTtwWaolzGf6kw/JZbpCTPrtKsUVrt3GCltxhL/zQ
kQz3CfXPvBRwOHELRABhCiKZshENFnVdJX1pZQG/d6CzdF+JUPYsCMDquY11
rDwL3sAELqgXxFSi1dAuhe3f6iNFodU8ytuyu9T5oBa/J294MhHuBkU81U9y
RdRwafjS2+8BTDi63AcZBVCCfoyRKjBdaVlUqXsci3xPiqKnPUlmhjLpR/de
TvLDTzgBM8Uevyup2oyoKg4bhsw4xTJcKMKF417rVh6dfo75uYA81N4ph8ke
HGENbczybpGVCsemgCc2D7l/HT/fbb9bUIu4hKutVZwWbFaLnXw96r6x8h4J
M+pvG4Uw2jn3b0TZM4YMr//ZY0h1emzw9QR2H566OfrKNullLphGGnNbplyO
fMe3NjWTV6hlOIIqyKD7wCMcrFoNJHAo/TXRt7kmNT9RfFkMe4jzEj31npcm
HYvzTAw/9LBXm3P6erS5r7cwbEAx8BtsHN/No8fDkl1BAmGGCmOy9UZYdtxx
gfqiRQDnNKjBGtBVMLaKcOU0aW7Uqq/XwagjA6A140lDhegZexrTx4IU9TqL
oN9+15Rdj58xjTh6H02Cs48zUEOjLsGyGAAX+spv5Gji6fbMJju94cdktHwX
4y+/gK6r3ubh3uv8NnqoFrPxWdicE/SpFT6LOBwzVqkzED+wBR9Wk4zL9spH
CtTWYbp+x91f4meOKygx6LN4KtykZZ62EvncUcl8mBUfYdtL45uySXbcz5Fb
Ta4yzpfZPsl7HOtk6pXfDzrRyQBV8TDnip1mrFm12/8e0iQXvg3thhDhNLSa
XbhYRjpnmP4AnyoaR+DEPS7Yz7WSC/MXQN7VN04ZG7I91upTuzLNvwb2mXbn
JypZZlet91OW55C50LcUdJC7yMaAOjiJVjmh+AJEj/Z97myRGnwDlAlsWgwp
KX22TOXcaKMnTqDfh2aren51HEIEX3s4H24hdLvp4tkE0/9C8V5JhjFZGW3E
ALNMrjsaOq2j9Wnhrp6/wjId8Ie1vj7yHD0YGDPBA/w67UaQIyEfCE2FpVpU
P4M+nRyZVe7y6/B1/DV4WYu1ZVOcWERZ2FoFgS7b08VK5Svoy/OtbMRacbM5
mFyX0gHg6ZTyAsHfD1Qt5fN/MQ160hVCepW95A2bAYB/RiVzAcqmflWoeV6p
axfpcYFgEHHH2CoeiHvMaLfK953Szi6o1tJL1J/Cp8lSDcDcQOyEVBPeMjHG
dz3quwgZ5DlFyT7/RhHk8IN46i3IKazIQ5Soo/41oC5P1ciNB0zzfp23L913
NgqCPdf9ym/pQLFpVIvn1oocOPc17Q03UbGGhB8N+zitBvSXrGDvNFXqErzB
CieEdhIu0U6f6KE2fg+Phzz+ApecDFDng19N5hE83dY7DBKV5BrLePYs/eAz
Viu1VdAITZNASIYCFsgStvPMPBVIsTi5tIUYNpIqJDQocAmNFUKdixLtUyfX
+OSalb0uc/snRIYs2tHuhNPvb0c0ChvzmmWrbBA3ZegpLiEqZLnUauGon1jZ
fTpxpQ2oxvmzy/NoU6hDilNVN+W6DAYdvAPJLTFRmM1PWcYShCWwWNmyNUrt
CLMY9PIdskWTlI/KBP8LEg9J3De1Scc3OFSutCoZG0mlOIkXrGxQ6bxmVn10
xz1GaEiAZXMUkuJe0D1Eii76mRa5E0wkKPt3W6hQDbHgJvVNxvIIA7IF7pJA
34DsJQ9xHq8QWZD9VCf1vnObvFP62raFO/aW0bmUJo9tBPjH+KcijkmdJUjL
AkL3FxK0WeDK2RQaK+7n/Nt9yXMrNaV8WhXbAdgVnohnJBFxKqBT+47m+g7s
HpkHFbKaWDFq3nX6dxZq1ykXevFENcKQbR4amA1zcHf3R6WM40ADmtohxUfu
M/h2uwbfjo9u5WVgTpDg57DX9n00BNFxN2WDseCu89enB1QWzvMa81obkCBI
VwZxOtvlBYqr7ud9T4YvH9IDpC4wXveKuidNu3xKSeu/5bsj6wWKM7sPeM+v
hwEntFxrtw69sLfzyl6zwCfknwzmPiMNrSZTbu0DcHiK7cXJMZdu4oCwWEz1
cyLeuhrFOsNFyMZXqApkZZ4o/32dpFCuDJ16yx8V1V9AyDN64wKn37lRYiBs
kXEZNu+03VxRxMYgBWV/AKViJrrvct6G2Z+Rtk6PPhMw95LBFFz2RQva8EQu
tliUAQ3rlOxqrJuCA3zQuiThVoUb4UzHeh/x1/pQ/wWOpCXFh2fbBYlV82ej
PX7w65+JSH09vhuzYEdw1Us50Kzut5lHL2kTypf6n08zBSwZewUUK0VcHeDa
+gnDmHs0CYo3Ac1Fe9XJTub1JwplE6sTyr7auo7vHh5PEwnKlmDJH1lXFsCD
uthayfQz5v/BV6etmaLTtPBQa6tS/CakijfTKIwEqvhQ/RDKkTpH41FP10ED
FAAvFfCq5MFYFAJqwV86WGl7rgpq+POuWj/IUNAuDM0WOhlNpQRN6sY/cYNo
8c7bB/SnEdIbRPybykadclv3/99Pn+QbDEsPq+8Ry+K6e6O4p6y6s/coyM50
OzVpsipyM3O4ekScZ+7XJjpdWaROZgHAYteSP5E1DC0eCPjkAp1Z8l0rNa+/
A+xLZ4nzk52eGShQTjUIX6i4b8Hz5nX2URCEs8mi7aqwAB0EKOjQfmJ6Mpmu
jBONo4eTIFzIuKb12MMegfXFAzJAkF5/gObRw13e0UX9kQpJ4swUx7q5VxHL
2Qn7TMfVUaXqBVgmaNPWg1Lgjgdts5JiExAzyOUKfp7x6qNBx8tpR4SIQlph
xwVn39xjpkDtqxXFxhWlZUTV4fFnMGvD6mBv89PLXo6DLTvSkDeoNDNyZEIR
SEk0B4O7jP9ZNWIz3lECGiMEAd+ruVYb5wAyoHwtTUmwYEKvCRiB6KUtWg/Z
PltILKGRf3rqnZsXAJCX3doUe0GUAEJoubnilgrpZ/W/sMvm/tmoxDHyHzRI
8n0AZDBCpWyUBjyoBTerjRW4T6O/ObcSjpijGKgjosmk1BrcKKW6EulscwbC
osWhelL9hTG1T5qvSsXfREiT8pFOzQlPh+sU1dTInFFP77WAgc5l3A6dSmV5
IT4E9EspEYVmhT4EVjIowcYI4cwe9uyYsq4Ln8ig586lA3/vgqnuilvrfrql
FrXy182/QRtgDt1xMx1I0eWK1Hc9lQt5e5o0b8RxbX/2cgrKJMsPWwGyTutv
8WO7xmDUC3ypnnjPc8z5ilBNeDW/riFWQGdnhjBacg/QycJadMG7JDj4YLUm
7WkbY4hVM8kWKlHzQgCcr2P//eDWZ319oYkMYAiMHrEXyISOHSscjpuuEPY3
dwiYnLW4U2NF9S2ckTBdJw6NUqMvbSEnqLUyRM/ZjX4KdBn8mKwdZo+cABNJ
dXEkqELt2yD5yMJKklQ+4NjhdzHme95rUHRfovXIZyGDEbvEjLS9NgPFe5/B
sgPyfFHlCNS+YOAZbAYyPccX2LJRhvSlRNnXpv/4mZNeTziRh225u4/QFZNs
5xcGLKhBr3+jeZEPddav7oxugnYhTPZNuNntn1fClkVOp148QLmuLoItTjBp
85b82PzlFFEXLJbWhCgSs40YWLV3iL3p2GFwhqTIPJsmUV37QT2myvgM310f
UaiPcjoNeo0SY0kE82jv+LIDHa/Iq6Wvg3xPGZtPkNooUfXkEcRhme0encQz
b31Tao+DZhAdhvW07fQn/YhMtkCj7e/RDmKnvs5EJ453GoCwaQDEG66UG+Ef
2wRm/THL9YvmuqsVaA/Aaz5MjUvZ7fjshzjA3o6Mhk4eT8iAmJiEt3n9kzXE
Qjs7voTLsSkUPW+TV4PrDBucHmwE3FlRsaR+kyjabrjv5q93uOz+4LeWRSJu
TZ8fupzltKjmfI5zIAOZxH32EtGs81bPf2+pzRPHHc7yV2ep60aGyi/vzu49
Uv4/05lzCCmIPwW/KQuyCKrhHO+cBzwGET5DhKEnpmOc7cHN+i4T/ZwgPCOs
LDYPY7ZdVzoH8uX8oR0IbtzQNd5/Fa4TEjR2721enZ4AcPb+W7uF0yMc1PKC
2Av0GV+DkFsnuYpb5yM9AYZcM67S+HS6o6lJ09ukvajSW7a3C2q1Mb6ilmMa
xQhYSM3AvPrnpjzUFmo5P/xxprxvDPQ1MPI9EEVTreJ8TL9OUbv1cF4UJYiW
SEHtgiHOlwkTiQDSAs7aBijz1BfdcjlKVZ/ISgf+wG5OfCJeRLKctB/cjkof
4c4/UhVnymVbGsUgjCIUAqIUK6HQm4KydZAVY4IO5Pd4K5rudocW6GrPiCyS
xYcMGya/W2ISb0WbKUmhM29bopDZ22FJRPGwk9tNx4z6Oh/WQVFL4erJHLAO
Q45mZfIuSDfc7OOE1k//NTLtiit+gLuywlgw1munZdvcCb5C4yR7L8KjTtoO
8ptzz3wGmL9BTsje0a/92+FsZZxN3//rmqx5wlfmALZ6GZJkAUU799/D2bsr
rXz2GXWN/vmU3P6/JDgaG+NA+pWvjj1Yopsd4Kmpdnl5m3K902U9+XKRpgiU
VCh9Qe2Z83ZUmUXSVUDDH1ABAxC+7/K2ib951ohmxd0/y5tGoYmntYwjkQon
eg0tJGw+ckB1qFaLEXqolIsIWXCLPy3oT3J45pizyoqPj7TBU7ZPiwRrt32y
FKrgp1mf0em885lTx7mu6FUHPtGHwin40dyWtW74MGMnE86czOnlDbrkx4ih
gHvMHPo717qkDzvdbFmiQaM4p+A1zEg3RgpGWpOuKGkyGaORQRLymKzh9mcX
RlXUUbHA1FrTSgLU5y34NsdZYkEq6OpO9cv1GC25zFdg8X0MPg8U7zVI23nG
OfV6Svap6tqmJwg7j2WhcYnKB/QUVb67ygdstYkYu1ninwIT2xLfOKVDsDOa
ksqH41G/a4hw1+okDPS6uXw4jzThZ9UJUQlOQomUVqrlVvIpfg3iYyGmzFND
DVmRBzie5Xn0sEDrB8lrCJ8JlFAJnHs4of+pBWK/YrLzMABdEtz4rPwUrdTF
qz8Ki4kV74j8CEwGikNl0AqITHFDUUSzGt/dFNk1NABKWOQDAmXhrL3S/8T/
jiVOTALceDkyyBQmnlSeDSJVJ2wMLO+xrNYzbqa+VbMjwab8we7jFs08Aind
dyEgnSHgpPMMiibLioW1R6IyNn2Bi4ltWFYHZUfZxKpxhn5uLaEMR6R967Xw
LwmEPQLurrIEKNu6miCEH4BLJ1FPxbnZ+/MUltFPyvNDwzMTQ988UoZ+XN58
fYIkZIWKv0gAOPg143deHvieG3GfG6jCdHMJFyS+XbbAFjU2UYpaI8KkxBHQ
C2nnaYIrLcUDqiQ7Ul6ojMXrDTfmqiE2Gkn6ZdMjSvsnNl+oAxUMpwxp+S1l
QQY2+tjDQVZVioH/t/r82DyqDzfpQ8emuMNs5GiVN/x4Cedu9e/9qkXdJLZV
sZJy8mHlt2wa9IRs7voJGDmZGfZq46DmtTzW1F+OS/ZAtIYS4nv411oP/t84
OOVC0DtQM+Y1ZX+HD7YjehVJJIjCyS99rcjJgHAGlLn4smRh87D3Lp2uqFVn
Ha4RHJ6wZVrqtGPJUFdXzX46X6wG+GLqdA9VwrYLCdKUbZG0lVVbBjtHLulq
mhh8Tyc/LSym4elE5USBhJ3dA72P6YtIk7YOMVvtJiUN8nqcgmvsWtLIIfH1
eEWcuMbuQubffHq9mjm7Qd5z9CxDADei/hfDscQiZnfK55fngeByqGmvQ8ss
usAe+xKcQHQq0zag0D82HeekUpHZQTxdinU+SGiAKle2U6P9YgyelBkYvIBK
QeB+ejAwiaOnuVi2DugjPTrxyDfsIGXAH+Zao+VCpPTg+a11d3whFiHsgAYL
ouGzzb/2D0TcCrX16VGrwfMrvH5xR/4UNAfvdeGNA8w25Z/VQhUvAqlbZ+wD
/hu2Vzc5/+wQhx95lV7vgKa1rV3nrIiSb1EadiSTqzxyhpVVpntxa+Upq1fi
QqY8HddFcpQggxH6MYI2wEQtF2V0zKpUEP/qokKJiuD3sATQVRASvi9QYxq4
8ui48baOoDsnxxcq3TFSsJ/7+yUVdUHH+YvKKPBzxDaJuEGBt0CphX1EFVMC
YDGQlxeb0v0hzjlJb4Cki8Giafd/PvIiT/Tf3ogRq5di45PZxSLURqIWLD2n
biJHsE/gcVs2R2BwEsW4jaVH1VkdyZ5GFcJQl+ESPwOzudAJuhfB6JfKIosp
yOrOco7FjaFofP/KT6OzMemz4FtvDWRE2/PTqoORXqRTZL15T/6A0eVfgw04
k4ij3SOsWJxKbqaJqbNcinCypWHlZ2gr0i6HfnXR8dtmplTeJ9E3Lwi1FqZK
G+OCNz+vUx3wZsfilTcf62HF1xkKxNHTxs9fU4VlkUBG5t9lLgmhEn6qQ2cx
7sXUDWxGHmQcNYYHoDFEMwnBfp/IMbktL6QcyAqjSgXTCfWftrk6DkaRdE/E
iLOKfvrwOEySHvj0D3rRdYDTpcEhlzrhfIZ/t6zXbyfPpSsou07j41WpLYKS
W8nfX0CrD/1VPSJHsavt1eVwvpG7FqmG4901OxejNl0VEH/e0W7/miDnzBiW
uuvcrLOG1QtygEH5HA6y4duv9r52FPDRRDrhsgVPQ2/xs9uYP0BlBxVnA7f0
oS9071MCDp3XUqKtxkqj79tYd4MR4M+WqhdZTAuH8KIURz2+g+G89G0VjPQ2
JCiNSdc8NX5CI+REUGUByiOjC7Mb9gazcg5PsCvAuh6q2gl5W5DOu9S1tr+D
1+YJHD2eTMevjNELDWj00PCuD5pKrGf9RVpQsZ+8kbUdaxceojeGyBHdkFkn
R+FlCnrlXiD9lReKyoUa6dTEsuu/1WXv8eH35v7YGUOEw8ETXdNRvedqO2ye
8zw7+7rpylVlQiUcQ8PAoXo+Ja8K6KSvH+6vWQIaM2Fo2umF7aQDaZl7OJb3
4kQoI9WD8ozRtanIzMCVIQkW7EmDQHlpgI1VKY7KJjq7TVckqkJtgA25IMtj
ZMW77wtuB+tEVJCfJWIkjbx1sCZqVZjHfoWnq3O7C/G0WpfLsh0y5cxHauH/
S04m9eRPucK2FfN8o8FU10CGNdf6PP/UHyYcS0nznR96fCZF1f536pLjKHeD
GC3anm6rwsYMbJ0jR0jfsRQNjC8FdGH21ubkPDo75qy8c61QyuADOw6l+E5H
1e/FQ3sXhIX7uBjlATnq60jAIWiXkY7MMb5ARe2OXa/X0Aq95XWoQG971M5g
GkokfAs6r49+4wiIdnFva8swU4DVaXUOUy+blesTagSNUhaNt+MEUtZwKZTD
4cGnpkLSoIpRbI67fB2vxGcDYiiFuQIx5eTMfoPA5H+5zCfSDyuaJ2t196wG
c+YG49RaXFpFG4HQk/o23UKcV4duSG5lRjmtNyv1ZTpaBo3Cx+iHQSGS2S1N
/Jp9SsbyQFyOedQ0C/DY4pt7/skP6mPybO0Z4iAEdCEmk11Kr7gc6BpIjBjo
x0twz0uWZ1jmPc8s1rDiaLZmgFxqg/Ba1q7+SaNYc3RlbTIKKq06oF8tMDPX
tTjLg8PloUF5x7CFUKzOV44zr+Cf7LrQ5B5aDewnEc/g7+SWOZPmYJJONS+k
07/6VN9/tuDNhjH8wZXjpJis7HO2R1P/I6+4R+op3KDYO5EDbFvGTFgp/77m
WsTXSE71PaofRqiOVNmUyFxgrv5YXW0m5VeFolommGyJb8Gg03AA8bcDYjxj
sNxc/uS0PDLxA6bN8Bhewi0bIYYjHK4u1CU0518n5d/G7IFfgfpo/KvxJeRz
jYZtwrGUH0NtS4CKSCdYJj9cwM4rGKlzOlxniwZOhhRFkkkoFvaSs1Bx+RGa
EqcYmsntCLWzAh/32XRWYFj4FrY+F7XDfJB223yzlCO0otFDy2WbHXtsODMI
yhWQ8obM5TUCop1ZIty6AT85g1Gr18REzL34gxaFo8I9jZtKdMla0fnYm9ck
Sx8HtXzlkUoJzBdJ824ILuCtBqK+oy2IyVJ8S7uINiJC8RizEqNbkB77tYmg
IZkomCUYaxmHIWIAkV4tQRGCa9Zq08fmegosfdMyZi6g7kA/xACDltRE4jRN
UDnSUyTw7YyW0a01THixGJ5MoFnZoMo+yrQEhgVcodsEZ5KeLFsMSMnx/0zs
Hfriu/TgrTSWcylqZAXRN2Z//7dGtM5oiYwxkx28uDR+pNRGxMlhSoGgITYV
TjwKIhucZ++0SFO+lE4F5nFwu06v0k6pGOHsrk6cYschhy/P6JYI9TtfMBU6
1/fnJKttDV6ozF3RhnYIXvkBf0j8houFIRRv7YfZuVTfLumFBWBrVwnQ8emE
3ttSNIrYvBW/ff0QJo5NqB2gVodu12pm+e83E4ic5bSE41gsEWCTGNC67Tsz
DJAKfe7CWjKmuFzsC5Vh+omfpAObvyfiYlVHJDiGXDhGABTVwNQJGZoAS+Gq
ru1qRd88ti5cGcduV1fknNrAq247wtVX7eHFZZMddNkGUEajgdeuwgx2vf6C
Txn/zz+XEVMfdT9tCaukd/0aeWnUSN526dzqv/VU/PcxfCHzWr8u9yiJM4T0
UB0UjIdFR90l8tPj8bRemoXxwJO9pMfzvD5QULqEu+QMbie9mzcCSX/65mHd
gOaNO1LiF3kG9+U0h1BWeM+W/IWW1AdFnWUzawvz50KU9IOwJkUx1Rib/1d+
sn8ZHOGTt0N+kH8R35Vq4joDAejRmiozQ97j4fVBgZhsj4K7BVpvbObYFVNd
QQi7v93NXzbmUomfbDUQXMhWdeHuSm4JFelE0RdqmBzjjh9NGpruoPvPuqfR
OeHIWyRzV9GmkRx/Kkee1K3doagMbSxRt39bS1aGpPQjRRle12MBOCAL6QcU
1r7BV7sTEGzAINQPn1rLJ+yneX/9e4V2pz3l6u0DaxfiRUeR8twlPP3T2xeS
C8FQgz9ZOCcw/muOe8vpVrj8KRJbKGJuwnz2nJo7H39rE1jSaVpKJhJXl7LX
MYSEZg6FNiMLY1CxsInM699sO20JEYqmGZ/nbG1AVELzyds/6q50natD9Zwa
zXhnrey0IdBhPiF6tAoSgZ09CcjjJQZRe2KfJo/TLbbomrS439ePfzXghYna
ZrYr5i2hWXBkbA86QUtfXSyNFMK/EF3o+PJ8WmIAEwEvBRj14x0pldpKzB/R
u+3UBV3BU+vrEO9WMa+tO1P5xagP4w17est+F9Da4iprnfYUvDIacSXS5JPn
GmjZgKX+RRb7iydivjmTbk7m3RcVJm/pIvCYLs8qlkxMRV/5GA2GSQ/eaifJ
DyYB6eEwMzhWNKC5jZ7+8cq+eX2iu/a+j5dqj9EXUG/aMER1ddzh32xbGl/H
QQMpVVeDOnl3sJZm+481n+LKod43zXciD+cG/3K8xoqtmyl2CBoCWxv+HBuc
LAONJ8zAm1LYQh65FMpWgDAKKdJxM61U1DqToMNbtFmsplinw5xktfO8TRKz
uRDGJJuML1g8a0TMgCsFhgloHWkjt0g23A/KerT13LtlqF/m0EZbmrdUBL18
tGURNSgasy/miUU586j0xIfCJ29Fnm9bgla1s77PPOEnxAVIxLZqhw7puVma
F2HkzfR9LFg0bAE7iVN836/Iy8o215jcabQfwY7qzXYA0uDRiuWSl8WxtHYz
C7ddXyOLpZ+l13JoAaDMFn4hBfkcYzMfWI0aQz2YHC8c7zd8lSEcHd8sxj1f
JYJuRf3b97434jPpsFhGJw+Zo9xZqEyOfqa0+kuWlogsTXCvy/YeDbBbdW9x
6OHafDNy2nimygQqoszX80plt/txSYJIqUH22U8r5r8IPyRzSdUdf6YzArqm
muFFGpByiLWCv5yP4XlYgtPgjoyY0FTjQKqhba+NAaVdXpIHRq0LuR3dFPv1
t3Nll+dWExvW63HlSB5VABWX9ovsvqvHM4Z2ka4wI8gNbsuvK4/YgTjEu1FN
RQQGpluitx8K+SXKen6Eq4im7VRUnw328DCNOeZoPeKUJktfnJdJ+TQwtyGW
b+OEOb9RSt6Hu7eDcpkYLdgsIbrB4s6prwSejIp7938UuGJUhUNDZEjNlb9Y
9uH0BgVKMfge/TEplPqkYvgwUioFNi663p+jVutP2MH5p5Q2mRxzBO6Bej5z
AfNA1Lvc+HkM+1sPY5ZICxhUF6VDkN+eF91trmgJiBpFEA5RDMgl0Z6Rci8c
GwO/DVlM/iJog4zEY35rZ3+roUzVsvgam6MJH5hTgZlFUN0R2WCl4LqqjR8Y
hKyR2GQ17R/w5qiNfCz9uz1CPJiJg7GP6UR/M0alASxmwqF6mgrs/SL7axht
iLEgoVetWRYhrkdiK2UR0+RC28Sb13iTUxXDRD/eJvpSFPfuSeVEn1S1XiKa
pfPCbtOZmQd4u8RYkl6jiyF3z/UdKBnb8J7QZPhCxpaCslwAshLBGFeydOtQ
VzVbPMBsrQNbfwyhloViq0TDB02q7wJEYr24hR5mzKdDQPxh6HmBclh6rVCn
iaWIRXfWKqxBI9KouDukOzoUnUpTwJSJ8CETg5NvuDbCwMIJev6XDu1AzR5A
MQiwcjTVWOQdsW1k8qBPcuDlGHvV8Z0GhfkS6LtJYOp+Szni02tmb2MfNwnJ
/XRJBoqBsdn0KfXjM3k6d+HihQMIdmpC0WkuOtj+b73K26NTShkYD1r/MlIA
8+F4/lUyQnRUbxjl9jqOp+J7jK4avNJhbtcHOh2vWdUwFZC6jhZl41CWnOa4
MAI42VLnrHDKPBEtDVAoFIF8fHHhgk6cq5aFsC4YGzN1CL5q5mA9TpnkwN6F
C7YDVG9bMbHVxP3N0meyvopUT6reyGyaWUiH7EaQ6OBxl9un0BJsywuUrUyL
h8vMbLGhM/YXYcT5fIMV+FVi1pxy7S2uiPUAUXNS/0UNKSbA5fy3DH6VyTdF
NMqlzpB4sUfvg3vH7QSyf+k6fypb3Ww+Q8nWSBl/22nk8+MJp1JFSEuDRG3c
M97ND6u9jUlPyKsFS1SjNvXRw78rMsMphDWiaWVxUn/SDmIJpQkMUxJze3Jm
RYcIetnKDng0QI6qUqFsKHLGxPFYCjrdy3fOzCVOGCcuYc/xquaZt7mfR0a+
Q867cyHfLvazVcm2hgSskpqITNMRNMibi2GuyNuO6va9Yas5xywqbjh8SB2z
oNNsMC8+LzizyL73JwGIMWXIoKLF0ynrW7AfIg9ld4Mdo52cklSM0mxzV3Lk
ZDWIojrGrBhTiXfNIbDBmb26gkldl4wSJHY1qZa67nZCFsKK4xNGtp6E/XIG
65mXPgKI9jOu4bfBo6OzONdOwBmpxy04eAWBFyaylK9PxuMeEH9636ouvbZb
5fO5z5e5yQuTAtjVd+mFLoSlCu5m1ywfJNPiDJ1IyEo4HQrcPNZqYXAEECtQ
5guR9XPnGxFvlOu1xGxBbRdFd0BGxUWKeI3OTgBBnP6+N5OMsXguoB6W2sWl
Zstiu2Je8xMZWFjod8RlPIi6atUh5P+GZ+u9tER0Rmi7aOAfSX7VwyXQNy7V
Iimc75580r5qku6r3kT1mrqoDsW+v8nOHNTG0X5ToGgl4y7U3yvC/dVE0HjJ
e/Iznp3XubmEpzP8mblMRBdbGK6K/q7MRBAFQUrEmzWg0PgUCy+kGcPlu4Pt
CKoqDrTPzBlBIUV0yN0HBOhbxo+kFdhnY0vq9Pogs2ZmRnZDziCVEOrjDZpZ
iVCObEKD4BhmsDf9izsxUhYUbG1kOXfFSCCZPpquivgIB9RWMzKm5xYcXP0d
FDVVDd6W/vjceO1BT80zx3SbHwDEnNaGUFN54Av1vdLDNvomwLV4MdTQtdSI
zMQP3fcSV2nGh+PT8gYYPJXQW7XyR9IRVC+OvEIu3q9w4WvxVHCxqdm6aP7l
tIQ/JdKbbBEnU9F3ZxadJh37yDAm8S/OMqyWCXvTkMCRpNVQ1CxgZZ409NUm
QdCSkLzi6WSL5DNkH0j5YJXt+bY7RU7FeVadZZnJ+i0FxJmIKGgeVphyjOrw
mToMZLZP4176wB01JDM3eTiOiepDBTkIWrJ0uN8f9D6vbvLimu4aWBdMonNb
UX7wPpQo2e/+QHLTGua9phtL4NtmJGlogOfbQfu11KC4raZH8EXDBOSdbKdK
j2BAbP+kM9S5bHMYikMAFHonofck4HP/UzlgID20sginACMf33JVR2V3AKYs
HtW80UDyqTuL3zDrFqHAHxY6kkVr46vNJgs7tC2DeSgmHiZ6+Yzevb/nhxPN
BtGEdsjX/3bqOzWLnVrVw93ESsHyGTKH0AVQZAopM88yXqYMP2IG6JI3xjhD
9paTHn1hy4VJ45ComUJXLgZGqf1Hzjgcf2mSHpDFQsOLnY6oapezu3MxL3pA
j86p1XTqZ4YHNS/ayn/QzBd88ZqWW4tGtw9X3dgnXEfSP2hPLJfEcPVVzVcv
EkQtQc1pTRMQeRNzml2GyvtCXWoITY/WbY6nr6CcwzDLKpj6g1v3FxPoIDOs
LkUf5i/H1LQ8Pd+t3fs9BTkOXjAU49XhB2tut6oTgBDe5zXjiA7DbpwcR/9b
13uBi+hfg7PxZ+848mn5wVjuLTxb70a9MFr3DA6rWWHWz5BpB5Gqb7V0G3ea
5PuHNLrGM4fIFzN1/z/+IywVcQyN4/kNm2XxqZa1SPq0LHvYLuMVoo8dvhaE
1MO1czUOlqJ89BYcSyzkpz0ejaPYQRkI5RC3Kle5gW2m3u6g9t/w+XJJzhYW
+mzi0LEUQkYDkS8MMIyDjMv1xiSQc4BXT3a3wdLFwQMlUHJbuBXY86FJfcXX
9I8ufYpyv8G0RjuOLNBcCQuAU354V5SAab7IQ3HDmF3yxIImukDDnPZ/KU0v
qQTi/uHv5yhKRvPpJZV0TTb0QNMa1JxNgZm8ETzU9NBC+nFQ17VKYCXlugXJ
1kA/G94RD+aQJspyyR/IMXfzRhpdzNszDICmSWuR/Eom/Q7CmB+WE86bmtxq
kt3Nskh7XPYFkBMgGDS/1Onw6+iXCe5K0NgBdo3t1NkxjCY+pEf0t5Knntsw
LGpxOynat+h7CzBoAwD0UXt88R34bST5yDOBqhnXrAjYWpemYVslTBPByuUM
+FIU3wWAVkZtL2RRe5MNNPnBQy5Za0vj473pfscj5vb+irYgn7fIZFt3Kg/3
LtdlyRFCoIUdyIJG969NJdGamV6WxvCSUOnwW/hwlHxbVEtN/7AEUhGV/2Vw
LmDJrBKtnnGtSn5xgQr2OSOVGIAzkXCdMjYBRvVAnThlGCNbCY/aEIVpCUSh
jEAeBR4StOOkKeVx/iLDdaMcRn35Bd4t1X99zHKMyvq1OaXs4YRXojtrnHJK
YZ0WW5PyDliYbXc+jSEdl6lFq0ixu+OKrlZWC4L1Y6r8JA/IM6wzH09sb6+z
aD2lTLd/hJ5CACkng93SI6lpXVkZ/xq09hG1wGj7QOko99wkpWMh5dX8tJnO
tLCG9lwwKZJ2/Z9rBo0WhYWG/BwYJhph16Wn1+iI1lzHlHja3w8aVDPg8a/q
jmkiJQrYNYT/ZutXrAs/cqE+dKGU0L7qNmIx0jNYSJDyc4hB/ppCxyZDllmU
g8/KgUPgYOqwXnCtD7zwu/CiKde8ir8s/PmyMe3CYxLlFYlGQJNWQMbMW9Nz
OWYRFF6gLpAZLXiok8Bhs+jbxcurKBOCbgk4BxRmr4TU172WLWQNvGjBFPdm
nT5/M+OJf6YRAMnaVHxYLHABt1iUGacmcZE/oRoAHoLcCD2hjJrPg3yXvwod
G8Ka2UUxGLiOBN1qNDQa/giYmmrScrMc2oQxhMsFX54KY2hVCqHo7ULYV8mz
4nYVixYfXDF2TGK5uMLx2dDF58jNiO7sESxONjXQIBe9h0g6yXZ8BEL0DYME
iU56ao9mmLl3mvCjf4Ed7nI2/cXEQqWwKCzCXbytJuRMwn3nQrox6AzHHNTN
E2frIObBwft1EnnGYK9xe85TwLDpyUUy47uPr8PY+rXVNPhtAiSB1T5tXMG/
5oxEznrMhSpjeEZdMrWVOaXp1nIzGxpxMj2/UYRQI4dvhTLHK7Z6W5drvtp2
FNrW/kDZ44hF2XQgqB+4YHaxERVp4YwkbdoP34qp3nTrvQKJWm5GQPWm3ou4
2+O+s2CnSWbzMauXOt4fsToynzOE8JQSYwE8wOpu0F8O4ofRikBd6G9Ykn2i
JCq33s206WtoZ2YCLagxSUO5GSqsqM8MIVTFVwfP2uCNfBbQNKjDCKWiFtn7
FSsZftFYI4tZVLpHQj9Y+ZFaXnnzWbqihQQy45ljiPZKdSM3CnVFFwARnPgK
UKY+HL9rBwk2tp37XwW8GomuEoqI1gC69ANXCx/yefQeWJu5e8QWB1mwy2sF
W+KQuk2abOpIkeMNhLZ+1N8Mb3UatgL7zmtEtrVAvacObAoA76Z6hHhkDSKH
oeg8/tJc5xUHf+o0o4bY4C7UtVo8t0WN1iaJl0nj3xNbUqj6hGpGNG4VRseg
MWoe8Nz9pzI3Wu+SBhGjacyT3mKcxXprfjqJnahNCzEHbxznCaa8juVTHCKt
6Qjg+FUk+ajYr7+BX7ngYkXQW3opCbZlsvpsKfM/q/HPPyBWucdzAIXkrQAp
yJAxQjt4W0wiE3apefdHZwFHp2tRcyBowfOPx5AlpjMmtTYFvTNfd7xSnslO
yjdK2QTfDQv93cqcphRoZxI6NB+cubp9VF7K5Cg3QA3liCErMo/eUCsLfVEb
3sga8ThGnk4K49B+kflrpE9dqc9dfn2xunUEHsl4m12NMQ12+fGJyyH71a9J
dqBkNj579T4Vc7jMWnHnpLlLemYN6SsALfD1eCv8HTV8GTPkElvqMHh4C9Nh
H0kk0FsuCmIW5ViPCgH9kupb5s9GJNFQEzE1lzH9OUtUwBDbXwK8Kn8wgFOw
arpK3FJkx9DcCCoSrMgZmJKfEqfnEy/FO+ky8NtX5qxVtaD/s4D+cUPeHmEe
JioPOorvwtl9xAZ1++FX8EUXWlCBhS9+y0dxe2MLFqDnyhl0ThlphyDOyqv2
3Wb0fx1O9XdEM4lw0PKOtb8VtvQ95+RyKziMvVrsxA/khFUk2Lk6HkaATgP/
jTmwpGFuoONFZ1fTWedzu66hpEGrmH9hA5JkoW754+wHtmYzQ+SkEhZuZFwm
dxGPgizyFR/5e0blSaGTWYCs5kznvhwxK/adSEqXXM/B6l1dQOrNph+PvScl
utF13pvRg3AmJsuN5Ia95ppOCvXM9F7YEn4zsypJmvoEnlxpL+b39YVnRxMO
QaO9Zc/35Sj+YWyydKSUmcY03qRn80La5VMLAcKv1WaVN8XYdUlq5nBs+fOJ
+y031p48Cs1Q7ZXQtUMS2eiHWjjBN2V9WJdSEMUjJFOy5kJCR2AROLBXoWmH
GWcE+7ZzQI9o3Y0ptXNcLncgmS5sN6Gcptz+ZnMUGrc482ExPZqCWKPxjMtA
DAS0vIwEZOCS66Qa6jUkLM9EEwgN92Y+W34TTAKaLjbaU+kIg+PxOSErz3mt
VMPq9+FZnMuOI+Beqp9wvHnSdRmUEapB/Yi9rIOaddnPmaBJKF0t3VzPN4RE
niuWSvSDG+fFwR0k16ADI8ODOWPsytjwErJ1Fwh01vlznlp/YkFyCGyLw9WD
cOO+vo08oHDwZtKFd1DUu4/Z/tTgRMYLw7BSczTXbuNec3LCkDnl1T5zT0Ar
9CzvI6AYU95UWJWycY//I8INfrvMqAOs1BaSWy7D6wfDmMkUl/KD7ANwBQGp
MWnvAyQrpNN/etHtAvep0xYieQFIdUSZvGD6BIa2szPo2lYYM8mfHBE3fUht
8HglO73OygE7xnExaVKB7zQTPEm0NyNZD0yZJscHgT7b9iv16tI721C5Pvhv
c4+FmntyQvUZB07ZkvFtqp3yJFQyFb+KRatZ1Ay5kenxqS6cZfEN3KyeDua+
vEGEUFRhPr9fu6MONeUCGyZTB6yEMR6s8BcNwbeZt6H1eKDvzrZ3uzuHNq3s
tfjwVPyvmPWico92piounEc2njJWNe4sVVsnACZQGHjPwx1yM52BTd/idYpi
Xn29EcLEZ9gnjH/QuGNu3jySN+j9DQID7NX5jfiNSyvyjeNeZnyZ3Nk89agv
e1BbriDqMdOOE1ySNDhHGNTx8yAWaaKdlkFw/TeMD2I6XZoIKGC5GSjq29F2
tezhobZDke1wLPGYD876HJJ2mDGQvweJ06Ggw8qtZnjaWn1gPrKG1rz+i5BW
wLjnigDpTsrZDZ/S0fvo3IpZE/3Y63sTcGgEZD6BZE/AUBS4Qe6o908L3S7S
hnD6wwuyRKAbDHASvtrTfYHMT3DaEToi1NjR9yZboBR/mtIUXyPa46jQXRrt
FQyDpdrUn1tQUk0y7gBexZ+i4vGRqBwVeZ8GHAEeIlKbgPZ+utq+ldSQ5XHu
Se4FPCvCJfO9AGHPHQ6qjF3Y+kQZE/7zi4teMCLd7dMBuQw8r8cHQBQjlRrH
kBYRqh2cCvygUrok9hYn0EpJFbDGGz7cCJNnHMiIOmzQZmIigGlq2H7FApCG
Wka6ExS2HuGvjpH1vSb6oAmIkKcL2vEGgrxgMUGLh/TmuFE6xO9BfSA+9C4l
K903LWGTAHhmAViWT3ang+YXrbFA2/Ic1x8RWkzVcaYcd1T+jkU/5RL9aWqr
cdoXl694+pWuPIPE6ZIa6KC6TqVD9YJjz3hj6XtATwreC0X2GlrUGin2rv+O
LCQteyPBTcdlq84DWEYMAQy6RKPFGyszcHCMVz2M+P/fj3TF4TD1UJUwF8fR
IsdBzHZ08GoTfWJrUTv37tkbE2rpi8MQeMtjEavOZ7QgjiM3Q9OB9I10C8WM
w0oOhE+5M4QfpfcucFz8D4v4q8tKSHrkbjSXo6myMtnOiTwRbw1LPlPko5uB
iSpdDvv2ZM/bwwecgOC0HT5iU7AfU+WN6/MV2QHQZ4IxH1ZIrern4cWe2T08
Mdw3tX4A/cPvSVUZFEq5o+IWDwUhKbN4FTTju7//XDWa+L+MASEWgDg7x0BM
NRQfVMGUtEGxTNgqHp+M133AcAEqegC0h6og5Pt6ZNTonJQ2vdvLmtxHWGWj
W+jdbVyVlv6jgPLaIWXXNT8ExdEjtYvwz8kX1hKkgM3WedwZS4tfGmcyXzqB
K5LkW0t3IKGnBKRI59fuhBMNa0+2g1UFHAuQKNVBKDWk0G/tX8wFtiSSyf/C
EJ6IbzTCAETtN2Au1rM1mcNzlTY7yrquz4hqwAPgHaI4bUjjV65rNuG0xLB8
naoZnmeSQGGGjk8uPVPmBMCF1jlpB0A/umhV3ZRE+yskN0H7oUCa1vfh+r20
MWOpgquzADlkl2E9Ltfi+LSuAYX34CVsBPLxH/4MCRu+9zT5i/WxGG23VeFY
Hr20qPpDvQuuXq57I6dkquf5p8ryzxQiy+M4Pnq+q/y/nvBhLCQayKpRmvB4
GrO3HerGLxpiO/o+883GLvfgCp3AXvaDCIkSgJgLMiuz1SL9NNEQny3E4u0l
nO92YvFU7hl58LeYmZC2ThNF9BXMj5DTZRAoV2vq3BQpMVDLciQ99Msh3Av7
PNumHtSZZEUEQ8kA5L0fLPhyTU42btIKbc08P3ohTO9aFKWXUqwWqBiUdzef
SI8RGd7krDiIwPJxeeYk44vHQTDZB6eXIDKQpkIv+lEA4IMean+3m/zQImpn
fEteuwLyGc7Snz8ztF9PVX/H3KZV1BUuuKVh3xP1CEFz/tv9w/ClqLw4wAwt
w1XrUfMVowxmLKrLlo13yIEezeh1os450zHM8Y51pVGGyXrS3NZrtXa001BK
JFHxY97/zpJFIbONzRkfZEzyeg6RvcOlryVbFFyA/XFbebhViAuJCW9f6LlY
3KIuYc0F0jtqO6SQOyI1JR2nwHjnKQIxX9bMAhpcQjij5xUW0y49IN9+jTbG
BSb34dV+MKsyEECLHAYkQi76bPSCR9oaemu1JKDZg//mjgXTDu2ptN3KolfA
x0/eUE4xJ7QXf3oh1OxMiXBOvcqoSlbSpOmPTSOa9jCjsEDTM4CmqA/U+iqE
hQlgQhF9EOsEdSWAA0s0uolf0YGlp4R4tDf+QRH6fwiO0qiRb8mbcM693RG+
F/0rJ3ra7EKwIYTKgzK6UOT/dks0hdA7/x25PuO7RlznFV7zdhljw8j/Ii4V
WBru3v194oZi4vHVuOXKrea1UR0uHOwCHd8SKLjieskmllO75FkyDHoGiUk1
NruM6PsUPVSE0XQnYB0VfGiOrB7aGz1FdZSF8C0p6uoB/zwXfn9ScDYrlb4h
/AjDtD1xKsYsb8k6iGJBMnZOIe8IuTPpRRAzf5RfnLR5ozkK8Hoit8NyWTZf
MLI9sWi21OznTapgs6CkcAtEV6MJNHply91BYl4BSVNOwi+R/b6GT/c9rm+J
DcbyISUu3c48do/PkQzRzBDtWuwEXM0u8dBWf0IYVO2ytScX7CfwATwZHvQt
QHprfQ3uAt4jGUlNqJf5axIhDj/ys4G1SXcGRPIi9j17ZDxFgVvp9D541fLq
hgrDjlYmdJU/i5oBfNrhWdH/jt9g/qS4vuv8SAXYiPrzxbaWJ6kcUywIJl+t
9nNUTnHSi+3bCqUoXSiymLXAijOlzhWucJA55wvLsvptFetG81uId7XagsS4
BUq+qDQMI/Hb6zIHm31gSFxBsxTXA5kSwqZdG0AKvIp0ZFgu0OKw+FeAeUbT
Z+URIVlIsI179dR+BiZ8HFH8hAtIYDGyv2rL44bf/HDtsr1kJNz9hEL9VZ0m
ECQR+wgfI79OkW6M0eiPC2sjOQ7qIiEfJnPPOe69f8PDqZ0egCZqL91YsL9P
3JCIKlSaW9/x5b4HArPa5qG6c8FpzPAtAju//p0xYopaBGQQSbyvQ9oEgYdV
LzWxxuGnC7njj+UVz9W92GnS9TSURo+k+EQpSYfFicYbZTznoraGgpIYyRvR
2nELXnu7mBC0cgB0OzxBmqz35WxwRmRq2p10+XiGGiHQM3b5A6eXhexGL0uM
GYNTZdP/46gGx+8q1SzTuWL3vsrSWX1nXbSg1x8z8aTt9XC2Mbo3EGPY1VHg
dGIR6eTZFbTfrgk+UKA5jtqQY8u+eEdWimxd+nmsNxiYMQQtYl770aw5VSfd
E3lNvyxX3u6YvhauzNaVbQrKjL/85/u6N1mIcbYD2TlwahW654xipfzxwquS
ivC6U5fhff2c76cYSRmnFOPMr8mZsixRNZEDrpBcoeT7z0/tCN0RF6QTQu9Q
JlK4k4avwibYjp06N8qhxHy9LQaXW709mmEEg9JLw2hW5Vp8LWe4VPdTQ8k/
Cg1A7Qe5XTOqQCH1kBfjN5ZsuttZczPwCOQzrc7FLSnT78uub3SUrB6gbxAe
UfZFDVdX+MV4oelNwJ6DNnhRerWksjQaJKOOAiRHI9kNdgnLPA7p8N8mtlSn
V27zGZ2bv1DDTB1jzxaa2YmF9Ut9QAG12e31oMd6pgdFSxsfHeoVsHK7q8zi
KR5Pool54MqD/OoHsd3DA+yu4Zc8jduU3hJVr4QDzEOg5tMIrEbKYgweS4MT
7nT2Hy/ebqqGtqO7b/vuld1p6vZL1xbW4dhKzsl9TbRSJoFEcsXbtlNb1jHU
OTWA69VH9MvtzwgjOzv/hAt2eBXdY8leHI35rN0Pp8+cV7ungyF5ytr+oCeH
pxfNE5iC4lADq1NGwluN4MOUM6bsWwXkGfdpKVIZoWpyb59Xg239Jz2P5If6
PAijwAOTfQl2o2pSBz0/xEnwue0x4sg+VyGiMoAZ7Jp+x8LbWvKhVmbu41e/
UvVl5E9qlbfriFKU1ktFZpgw90gWX0QqMfvElQ8NNpNpxjOVzG9ULi9iUVIk
TADdGz0e2HMIAl/1eajmcFvn9dE91ZsM1KQx3NozJl8G68E9519opfmP6aNF
RC//ioo9oglXOTTEtzDX4Wncz+Qw6QJnfTRZNjAJk8zaGaDKhei+DtbI8yD9
F7jPW+0jGbc5auUP4n/LOkJLpj2XzNF9hulFTZWlYECemxOtcxvMgwnKF4fK
+fhZFXITo+O8zb15yAaaZ4YGbvEOOS5nwYHoXjlSoM6jw2seXw3x99Z6G0Ra
mDMTpbZXgRUr3bXug0QrG8B8yCELURlP17NrF78BV7ZY+Csjif88UicGl33Z
f4g5t1W73hy9bY0oOT1H5a8gWXRm8L6yZGdV11YpwkalJUL3xgecOrp7ij6J
7VUlJULiW29YKu+flncG2YM0gdLydviD+PxDCsssx8jnom3HwKl3V8ttTJ5F
Fre7OMLeBrsdj/D9RH1aOt+3h+DvC2EbYYSF9eVmAGNXR+kjdr5OwYneJv5U
XxU2Xh5U4TQohj7xKiPHh/MYOuAMrfiJ66hhDQAT609vW6Vn5sks64fvRNGM
r6Vnv8NZzgQOZsKllDjDL86vG5UPk0MMpKth914JVGN2h2X14021UqYSI00E
nAJSZLdo9ilOGTyzgHHcRViTYist7chUPX3sf6Sf+DMvIVm9BpK7XG3cjC9z
QKuE43LuIsBfxDFwe2NWmUHbpu5UVMChHUqEJrJQ/N+meyfj+o2/7LDEjJi0
+L6qEkR7cfYw1vEU2z8v4c1NvG7El7na2ARolwm7D0pxNANTJ2SMRI+7U6AI
hVMOHQY4cZoqbNmWkbvXfJ/Ypc8YyffxLBfIj6EU5NyAgH2Fcmx/CwlpI492
mS+Favai40CwhoOk9nAdevbOOGw0o0ReCGnXOJp8cDPbRWXNsXIQqXSX+1Ow
dJfDWcy2kIfa6c5PksUr7LDTy8T6BkczDfHBdrGvV/s/q6C7BnGoejkepTlb
7EGtuf/l76Rz8urnRjeQTno4w9gNQWBMWl1EULMNeRHooTcbOZA82y6Gm9Nv
Kh07CJr9k/IEqnE1qOFq1tamghBlA0nD1EEyDMAQFlKswbA7vY3cixEvfbob
oDm7uaNiKcAeZNpTl4doZlgF2y20rcAN2LcA+Hv/fEnVtcsKoVVW1pBtfpa0
ECKH8+OuHiPr30vrEmXZ8ABBbpkRpjUZK3PTLApFQwPJ5F9cI1P2NvT4YfL3
MQguX6kIYeWB8t6UsQcaVTA8IUwXTp5sife4lntUOcilG91kwp/2KnOIf7FQ
Vd8D5A0fsLCu0cosndmPC9z2EfkV1jnkGK4wkNjTdOQGvtXzgaMvZwsjIyUk
c9GLfxHUSUJXEkbKxO4Y9+IBO1n6QPHAmnaRKsse4xqB+021cJqZuCkGXDjj
5pPLxtTOS/gUlW71Zz9+adbzKM4y7/CCmB3x183PUjdKPzw2yYjNPz3D9nH3
gl2IB4OQJvSsKlL8fMvClEa1LeuHd1kuJVeKsXIURDvTR/CUvk6CobwQy471
AjJMDNdauadxa87Qiq1lHnQWHJAdEwSuzRasxB3xygwBwSiUN1iRPsn3kFQX
W0Ek7sNiNIiRWJ9FWqwLpTY3bIGAektt2fC92T4PqJOaWODblbHCixDH9p/5
05HI8PAfb3MxPbFN6KSZAhnjnGiVJJQDUoDTuMScyOUYnWnAU960jmb68gq9
NlCsCpmY094Lg2W2IMNzAZwVaOgpp+WHQ4W/Q5ZFrpLktcKnGdMqq0BvfXNY
k1YZAXmP7QH6GP0lpj/qTjxKU28+PHWw4UTPuy5y9j6b1L/KcOEgD0/b24Tk
IGQw8JkUZmTvZyPgn3SgshPwaJTBX8X7qdpkNzgula+wXFBb7TkTpu+kLWHC
0q4Hv3Tm1pYePjJRn6W4Mc1+9//5uXznadhNPQd71KnwauEsda9zAfEAms3p
3J7QS5P7OLzErbdmd3ABCwKqxKcn4cuO0FQycxy1mmTybRpyDj9Qc0zFDSNW
th3ydQgTRnkMCJdhxh9SkUVrQW0AK48um22pZeb1L58LMhoLcIgu5Yt6Xfn5
Mh+XTpX3KJYMdpjYQlqz7Be84ROE3QIy60uPfPJ6wdvPNCW7emdW0ertrL2e
Sq9WA3Edg8Vs1VjKEXismYNNJ4ywcVdkuCOqM4CSJPo0Zg8vjWDoW8w3Uo3L
3qJ6nA3pYdn3jdeEbdv0hKtGyCWSuZcBFKBNRIQkRhGmvwBYBSNItvcU2U3b
/Oox0l32SjelW7x1xs+csQ+rxSN6tuf+blvkQJ+FUhhAnDyZdKXacZ4ce1v+
cQQwYkhSCNpVPeX3suW4cO9IS+wP7nOS1R0uO6Xmj3K8YdZx1IRZbtvs+XLf
4F90Mox7DRh5k/toCi5rF9MOH81YZ5AA5BmoB1icPKotYa0QKDHZ6SKlWJAJ
7q+QruB47Z6Ku9JjzXXb2G++k3HAH8XBUMKqQ6bJSIiUe1vTwkQvW4wvYuwC
oqu6OHPoJIxVOnXmxpxbocNjC+TYEnEEpbCFdriKILD/CGZISitIw57jACkv
EX2eoL0nDpnPtPnobhL4GiGX7seOlFe4mOjNqy/06Ug9dEkXjeG0qKKfqOwm
KCvpuTLvWXkEU8spQuquU5yoncd1wvcMtWBSMXPO0LBxlqLk3mbX6WUTJ2wr
iJ7nDXIlb0UI5BScZ06yplhpDq/gEVDsCOnOsEAGkrgvEgQSLR7shof/3sTW
UkyaAjxPst/tL8eAzriSwQORrBS3FIn+UNlEK9odEYNVnQZNAHoAxLec0vcU
Ybuv7qf5Xrv21Flo5omtU2Q0Hs4JUIHjZFIYWVZ6pG5f+OHpHigwEgQW2+nP
4y6ypCJt7Lul2l6EZfmeZoftuPIYi8L61obDdr1tNvQJqpdRSxkvPTv4B74/
695/jwEVoXgFevTBVW9oytLPLluasS8DjZoYpk35buGggVX+MnqCz2idEld6
NnG/G1gLBwDqLCwdTGOPpBznY2Gn0FTpuWFVhZdO6q7/clXJZbQlK9YIkQ4u
HKTFPuz3QpE1IoYQTYjqp63Oz9emq+7Sflgxa3meka1Wc3w1sVJdehr/bqZx
OTd+I9i8TH/9F4rMtidLMUNRB03xZ/wabUlPtXifQvFp3hcbSKFzUAcY6I8U
oTNHYWv8aJBSIF1w4svSWTDf7jCd+CfFeiL0tAyOutlerA3J6w0hprTrgK7f
cySRcdH7+KFRt5yXJfePj4gAJGbM18reCCzZOuCqOaCszYoF8pI28EnygRKf
ifDx7dDHsJO5ilA6AshTeqxi4cBghblcd/Ez9jPMPMrkM+fxMvQoOJlsKsYB
yIdWTzF7pEIfHo61+exaiJGh5YfhI3i9B42Ta/Sh4xo4HuGvFYnIYP59RS1P
rePe7IbjWDBenK8zivgJiDKb54HsqyHO4UUGD5VUw86FbZNrrts7sAtU7a/E
ySdDVH48Q0NOEwtn4gLL/GKe5vKsgKZqEd62FmlspOA9KjuUGaL9Syk+ewA6
H8tGxmzDPPu3pfbenhvDA3U3iXsoeds99PTJSIHXjNzxBlUxv14Q9PtpQacm
9FHMxOo5nXO/kPAZe5TON7r4hkv2yR+CWnVDpSMZQ8hUTK+y83fdwmDJKLWL
5VP0KI9EgZxHWTshUmTETCC49R8Izcb2gpIs08eYuhtg3hwdNptdCQk2WVQ/
Y+fqSajBvrvSfgVhqtt0Vw7vctYCsMlaw6y1Dg9iv1lQO/Kg6fIJXT+CSqw6
E1aPrO3r3YYj0rA/HLY7xFLUDwcKq2ypQeBJDtqyAwuRP97iS1KWgHKLaEwT
nDjmHVY50uhsr0qqupmxt0GHCnlPqA+2SXForhW/5xT1KXXlnk2ycTcIpy6A
wV+WWkekTSqpc+T4F1ELcASpHIADcZG8N8zxWgLO2mv+QKPzoZIRqc8VNULr
QBdURXnItEv9MqoK0JH3KjdBTT9/ljDsugdQXKYcx4d/SZKDrvPEBGNZqmMX
+VLl1yOthODebMDCKCfRS278NE4eLYFnVeuoyFSoHM+FEur2saN1oBYmG5ZR
7lgQqabeWKFJkpevFiHv2G9MumHdgOZiIouQDJB2xfw+X2hHRdOB6B39udNQ
LfssfiPt8mGsINJPvG0F3d1I8qYcAjnrnJyZdWz7+9dKyG1FJwCoAX+a4NrP
tOBX6H+ateb50KjFxzRUm3T8vUEz4LeOgSOr/+qoxjSRsmTF7BxIpvd1fGgI
iD+QobOirCT+IATvdEyKAgQEKFEhle3ayst9Eg6ibeYCrUZ9+fUERjyfO5uO
WBJ+Ek7O8uP9KKjwHPyjzmuU3Uqo8Q3buT6EUXRSzbycBSTl/zJ90XkvtLm4
iNhbBqH7UR7izFQdkeeGIL1/we2Tq3dpPi2Ot8mpumxQJGZ57GmFCqxRphhw
3197SBj73EanM+jzrxkIPn21m1g9Ag/FJHG5xPHMfJ0pwhxruQQyTq4Yf17I
LZqUNLuKKMfZAscroGHH155xL91CvlWD2Gcmkjn20d7ek6kiPdyb25QjyTje
PzhMUCWl/mprpovwKKK59oUWeRsp8ET7Kr1l0DzC8HWRnOxQgSF7tsqG34sb
gUfdvjGZFX4bvjbqrhNWA8J+X9agbPSb3aRl0X40NAe4OoLoIW8FSypDa6J1
GbvjNRNxm17T6OMUZZl4e0HA69IR8tXqPFiuwlTN5t++GmDC2vICBz09tu0a
LahESpcklmPw+irWnndNdLiOJcs3YAqXQnEH7mtyPHbFumzGhaBQyVuoFlFG
GAaUK+hit/H0YREz3+NRpChjd962DyysXSb4eWSuxx5M9q4HcfWVTF1487RS
uVYILIBMCuVAKmJYee0aN8XBE5WjWucdJMUfamlZH2UCIDL72Rj0RE5vrxqV
L4GRV7xnieT5ts0CLxNoOT3zyUbfXV/ro4d3EDA+x5JmoVxroN1pWU1j9EKM
zuUg/uDXkBiAX4iYfvJffA5cfYrwpjIgCtQzmB2XH1+hgiM3c249BjyucMEP
k2Nvvc9ku+Cp7y0JL4Qt83xVzswFez/u65i2+awTANCfG6ZIaDJMFEci1OZy
HYANR0IEoXFWAr70KtNUPTovuahuE1ec+LwYERxlC3m8Q2sKaT/kiZcGY1BV
JW4ifRpYa7LGOLsbAEnfT68X8GrtEOvw9zbIydOZrJswDCNAY5jEKL1g6auK
cOYqb/pt3SfxNKtUDFE+c/HjrOEd+0Lq7ZhXHXEnRl/CmRytrFnEF7nPWCty
uD+mrAL2/GrfRv3L+JQGz2JjOVSz/ZMDV9ibliQ3RTwlU11+vsWlOCQ0FvMC
GPljvUhcSfA188RDAHpyZqEZkzCmCwcsc/ZzJXdwwXjxLpdZdCeVpsgzD4hw
BkOSJ/zI9Z3kjhsIrHoCAS6F9VvqICPd/DbjCcLxUw38mBjcAsP8MKXQvxa/
E1h96KpJPGvijh71dZFLKL95FkHlOFtR71GzCFz39D35o/o7HVuvPnjVkYTt
al2RBHuxRWAIwPg/cDiD9Qipz5eXBOTckbzGDke1LcVJbjS9nk99KUv9s3we
NtaHAgi+Ojqr2XtlSi/uw4HZHnkDa9trf0auraxmf42NwaCQPZUw6cEfAnOR
5g6APNKBg66yJnirau7tI7szSJHGoLo4/eebtN0vysURxzAPpxPSmTctPglP
Qy7Jq3NnFdIUMfNTRuKjx+GDW3tC7WVqbIv1XTkcesqt+WQp5l1U1O/A6OOh
W670xpoaf9hhIeCK0RVrZXGtrzj+YZWAJi4HAk7RQgZr3x3kdA2p68IwQoDN
m68V1VkRl8Ztm5ghEd6lDnafNBxbaNezf4viUilAiDqrkH6txxD+QfWwMgHl
7En6tJBf8T6/PhId4J5aqR3tNV1l7hyTh429aOi1xEhT9sCkH/kSq8Fw8lDu
y+2OX1LhNpoCUMWYjmdpoVnWy18X+abybjiIQlYunv8MKXoPvwE7xh0wmLnB
CQE7EbhBeIJthTQlxpGiMuDtOAv0EKcKFsBZYHE902uX6+7yIAV9qqvjvK0c
QVx7qxlTP6XW0+bFZIFD76OYkS5/ihL5cWTR9YEuSW3nhia/NFwEl1cWRvS6
JdZtUVBf4+AjBh4ylCxZw6fgd6xu5yLp3oDhw2L2TTHtJgidwiYjLx7JD4Dg
di0UM7LrS0+kJt69upex8Doq4x4BmxfiRg9NJJt/OfHC6S1DqNQBL6wlMkhL
1KWf1ozx48CvEHvIlwiGWQbQcLvryqmkTWgLcngxFwYUQ/8zK4oMTRIiKzV0
3cacH/otLxEPJlu0FfO6qkFnhtuxD/8kvP77x6dgKqSVP0yjm/gHnQ8JDEYa
VKHGkW/1ya6vJa08HcX4ZswIKiSP1LeehqU6PIW+Zt3GpR/nNE6tGbs6fOyt
aSULH7w1kc9rLHJjjOYvUqlzhpqb3kD0p0YxDw1ZmKNGjualAMnxgVD0XeMZ
OsnjyvvfUwy71+4EZ4HtTcFczF5+tLnJIxTXiK3ex6h2Fc4EA7Qhl3GPPdC2
MLlNN5kBmDR041psTDf6XI7ktrBiHyfyFl+6/5SXw59E5I0zmrur/J4yCOkV
S9i/FnSbE7BdDkfqGtp747/GhXn6EooDZNzDWwYydorq14ghzDcBU1sXKBmq
Ys9WHFhavGFfxCyJ02YOj4dqWd0Vrw0R/vovZ0rR7yNJq2kvj4I/0f67RNdM
bb5IvskuuJOYl3SYeLWBqspHao7zwY+bazi56NUjJ8RtJWEZsKapPZ3wa/Aw
Il/ez9JqQ7OE3R/loiODTp6kMhRoRRocKp55RGD1n9X5bQJ8a2xVCXUI+0kb
o2kOnEj/WItkx/sROB4zjXCSh5/PZoCKk7szg8ZVR+XhTbdrN/jailLvlMaF
Tkz3I6IHyb6RsOsb4ODIlRIrgzHpdonsPa0BvB8XlSLhb2HZBrclLJwAGuH7
bcW0o6vdvsAk2Ytg3aJg9+dUO29HITR6/vIEfXgevtiZJSW+HU04nIOk9dHW
YPeILyHXFoRKmtJviMFExQx2ukyfW7lto/oBAEOTIwK1BRjjz8OJYhJBaPwQ
CZQ1inMF/3YRUXpwiC4f8vnepJDzsmxvpWUUTdkTspADMJgtp/PdVIe7ixxq
oKuQQpqeqdyUUILTZoz79T8Ijd05enR/9nZ410AQWw/AjB3QPQrzQRMKJcH6
2ULlCtYIALBLI+FrWnSKQvE1FgsBwxkhU28rQWGNHkHKOGyObtfurAr251p9
2PwCkiE9MrNupbFhrvTvEkKGCPTIqlntBe3gZld5WIEFtdlo4w0tcsYmvN86
2v9o8w9M581b/CV2SGoYA+kUz2hlKsbIQ4Zw7gT0qdy1i6P2GFIF7+DtNy1N
gd0gA0eFKlVInN1I+5yLU88xX7fNrcEU2Lm7J+HRont7YHlZN11I3RxJEMKI
nJ8OvSuq+EOkT6IO3sxtgptjeLsXcF0QoGFzA3fx28KsK5SfCgTGvVg78QLL
05c+ZrqiWeFW9Ey1Y4bvaw8NQ2OjMfm/87S9nA7ouZEM/9r1N0Kd048xCqgM
gTMgpf/oUdOGWiEV52pKU9BQBmtyWL9sbT+xu7DkVpxDowPpP7yHY+lJ32fH
kibUHnP0DGsFGAnh07ur+jSwKwgSVWeJ25yHhC7fag12DwguvWPGKzI/nYcP
2pNnDbC8+A0imgg2VsYX4elDLuwDLPFpgtWEXDrFXFB97li1w9khOWRm/Jr8
0u7gpPatqDe6po/sUNB6LB1LwkomXfBYnbdLCmu/zjfAVLxDPOZpWnTjC9kS
WYk76GHFRcxZDYkCwPelMB/DkD+XZUdJcGlAnXI36frFilFrz/LK3XCGxjh/
yXr0rWGI01rIGvxFgHV/npa1sbjzgxOBwsKG9VkbnWlrHa2dalk9y4St6TuG
y35OU7vz/bV0U2rRmpKlVGklpbS5VqJgnVUcKSJXCY0lngY3Sec+Q1suBU5Q
wmGuhjrC3nUyN3NnOWOBn7FP01s9NjeUylwSQaXCJZDCUcx5vYqMCr7pH331
cy6MhlJ+Hwm+boh8dgfXPEmaw43d24FBKmLO4VFjx17Z4u/RkJAsxaZY04qg
Bmgp5AgoOOT+gfzE8fZRiyrWwxgAECgcMt60Esr814nERDasrWlYvAOK8oeE
M+7tZI0uRHtXOCMSR9mjrmBlDIV2SPSQ9TH++zH28/Cqt4yTQn5nBUB6LtO0
guHq0KepezJnFGTWEnkjrkrF83ez0t70qYHx53K9Y9mxYRixFbg9rl0hxwFM
MmJmi/KBeqke4qMzBzS8gZUdYxPM1GC2Xbs5C3NCHy3zXOTo77+IjTeinSDF
0WYXSMayIexKUcCZMZYX3nhEeaF4Mnw1Ev56npYLj1bxGWhdGAOZuFTdFY7Z
trQbKH58DN1lF6tE8DK2MCIrs+Lsy4zaj10/8affQNC+qC6r4P0TsTTvQZKG
BbWI2muOFKpAX6bXyINR/jwHVTNOg/vz2iGEZ+sr7hIUielTJmcxKirZoeor
QaVLrqBXyMgSLhxe0qSd8tPHNGsM0PR+oIAsePtbUXR+f7LUB+8Ue1QdJAgm
ozzpc3Zi6Ct/z/wJdhTnuddvJ1iTfcooYY/pfWrbMdWt4cypPswnQKlxRTFc
4a3ElwdFzt0wWcNXjtn6jpkigw1eQroMfhnJqqwSJLHA4ee/pbDnUrFGmKQn
T9NZqg5FN7drTZsZCFL47MQU3fMHsJNtJ1l0vcv5y1L1jrbfFJZSvLP2MwXb
XjGUc90SqqgXdh2fosWUBzEe+0HGZcOtwuxFpOSShDgWdm/zMx3o8SNssjKo
2x5dLBDjjn48tRb371mjatiuHlFAFKCIEGqzMXXJwoT1yPuDpzytAPlc6RKQ
q3NTJ1Rp+3NQ8O/4ruxciip5+adgUMpd1Q4NnwIQJBRqdf4U29to9p3icQo5
sUt8qkJBaEPa0js5z8Bk3+LvP7+/7uO62EJLeDHM7J/lH2uMARPLmdulQS72
88rG2tRF8Sz81hsUITtLjrz7tAZm7R/oNdDp+ajvSNAnYx/LZw+HwUDzMlVq
5phFtH0k9suTuj0q4cdSW7TzazasZW6Mm89HPUNeFZMtGGx30VJEmVo36+wa
rMpvMGtDUzzrNqQQKwXW/vZXdvpLhHIS498E5Pqq/K/ySS/ORlh5FsyeLodG
fYZswF1K/60MaGlrI7uS/v7moWPzY4tgSiUD3Fn4L5LzrjGEf1v8ffECmhW0
YrBaDGFJImIyIGT4Ob8tfc69kXlQrde8/Fg7t1hdPBJoKlAOZKAaOAY5iozQ
lKcuBin+kuPvdzIukQhtKpHyDsvMn+NcQkzcV8ASeL8OAoTnfBQ0U9nhb4Wx
0yiltgPKugDsrBxdekFK2HRp2VSirM5mQt8OPhDbsYh8QQQQ86ifQcPu9Zhe
MyLgW4gvbV6LHszYaDcrCqXh/5iinfpP3a24IiV283BCydG4vKMr+9UtnsRq
ochrWkxt55Ele9DG9dW1DJZcbnK4aEdK9W74jnUruc1W05tmLA9UrOnsKitu
1q1sLh66tVbJJkRWaca5/KRjwOaVHFlK4Y3J3KpBRGm3HQbfoLdHt+nNBI6N
Km9wkqk0ybmDJgvJg0pWpSJTknsN5abnLjM4yjbK5qy9iizeMtXLhDlHn4PX
LD6PdYQdqWcld0LEOAkeN8Y4KWY9teiY+EP0wp79whMsOPkOGtrZGZm5dhFE
1sVP52gSJ/4tkNZkmQ65DcSqsh43LxYqDjNP5sud75vMb2bWw74Hvtrrh2Rv
Gp0nH3EmDmB7THDdFVwu/m3/w8y+xKJEKKSpKYxT30qCjv4RJD9QxJjHSF4z
0i2fzJScDsHTVBHOtoH4mi7yV/LOCVqe6pXXNgdzq3zFaH9Q4vszjt1qyOy9
nkkxVsNuHHraA6MhyLzlZwiai8r4kWkaBeqiJKAtyiZQol07Ij2iKTnyV4Zt
Q/C4gR011EfZmDZrlEA5CHm1MQDcMdbYMjWDIkvOAlDPNP7v222ir40suLnx
/8Spe4ghkLD9amDyLYPZKW7RlHXBrvW5TTfNBYHtBeYe9YYNQBvMETy6Leo2
IIRRvm+Smmetxf4xEEnQ+U0pXOC0HdhuDL6069dbVi+qQUadIK7y5Ht2lRXn
ek9VrnXjsCju2hR550u6oH82T/n0GYByHXwtSu6ik7vYe+xR1Q+HuFZKDKY8
Tg49c5NT6+64oz4/BNwJNlgrru9SVt+r819fuoikOK6aM9BDfiAM+cuxJHlK
+qZR6RinWh0Imohz5BQaPIYxof9VaVaGICEjBH5Xkw6EloZLhNbL+K11N5d5
VEMzzJaD/lH6s1fzyK+/c8PRDcChTq5SuJHl4D/tOVEjF5YCx2rVHJrftkF3
yp6UOuMLhF6pGR1NK2Ov4TekRaeaZMr5xHbI69b60aPgkMDo8lXjZ6hRB7Ip
1ME27RDkP7RU8A6EB7y9sQwgqMtTu2r8GNrGzA5YE3V/Ag98GxiUpO7ApEmL
THaXlpme0p0mfnSB4BCCTo9IaYfUvB32HXWzK5dX9SU8g1XRT1bhgK92SaZn
8kQzFVfpFaU2tZVG0vwYt/gDudv/E6MWJ7aBcdfA3PxdL4XS2mZnLN7Fr2W/
SUkJXXIhIP6Speyt4/wCg8d+VWDTdFdv2tNmvh+Vo5KSevmai5fYW2Zpi0d3
bs5w/vrSYmn4rPF/e4RR0aPcXip849DPxStenpQ6KBarrGLNxhz1Iii6SeIu
sABP/oWugbXq/zE4VCGJYNQOlaF9wiEt+ti3+HLP0zY+biUDqoSgRWc3nEpk
LX+gGO6sDZdGf8dgecMZ8/1O6rL/DOGSMLNQrXDDkdvfBqt1xdohQ86MESOt
7blCk3P/n/zU1Ep8lRVOfeg6oWzXc1C18qfFzdlg58AVwKVFRqW2AzWbpPhM
9JpH+9Vb8mh/w41mF3MGXBp4qvnphpV0lQ3VeSF+yjWSi2H/VUZeuXK4jdRz
u5NsoEtiZakquZVdRtEoIgUcHzmjYufUV99k0iKu8W8Momu5D4SleJzX6sfy
Xyu2DhWHKBVyO0T88elZ6rD8Ytk5BZhn2bmqrAT81VPl/GaSNMizH3vyd9/V
6ner1slwW8fGZeDjxh3088q56enx+9jopM5XYeVKJKF+ecCWBEuRXyco4Veb
i4/2Hmn4VBJCrV0fhJlMCIkXXwN1Unvm6N03PteZ049WG7RC2ayXVd06xZx3
QGNUAHElIuoplT1zYCoXsf1XpVlmRojscRiiBaPmv/Zabi2Un2/i/Hq9q2Ny
w5YgnVYt78rIMnRQL7E0RF6tdwtOlZhz2aTEa5eiAfLftsJKd/37xO5RgIhY
56p9KlB8+xrZydu9RtxuiUh9apxd+DzqB8afEwwuauNtIrarqbpEaEscwG/7
91K/8/PoP7+ExN5cKfCA+wfZ5ZqpezSX3H08Chkq/56oxYGW+/w3w1zGbsnP
1G0j+pxIUb7KIlrU6xIItFyMwzj+YkJB2+jBQmxUTl0iwV9lWtI2yTXDOnA2
k3qZPADGnhkiRYLBYby+EnY0pAQQKN/4Y3BhU9K/3Hb3bNMEy7TiU520PJ/3
wDL8I2gYkhWImH2BQ6J888QWYLhWvGEcloutxWHfGeV5oq3prOjmQlAWwj/3
JjnWK2QrvmWSGZo8/A8qZUrTwM9oV4oGDvKuuS2mOUAynYyPqIHF90mdhkLF
i0bk9ms6D1NXZlascfuNvktpdWibMXKm93q8U5n4JwZYiC0jXrpMTmu9NgHa
PnSCAcsKmH0LLZ9SHpLpmg3NZEttGrKXG2oScUsiKud3T39bOwY0oGHq67Wy
fmiTWVA06gQDccwEoUkclp9r3nGkhIQxGvLxFMNTf0/ewwtluk6ejseONC5F
zsry4SZyZQ3wir46E+33ZkVD0Rlzr9q1DUxm0N0DXncad3WPNx3wZQlyVl75
PanjGh93lR6Eeq28CC1QswAXs2TgVT2or3cJ/ydhES1YFUeiDNhvxrB9c3Jb
S1xUnmiavmVXv8MRo/1TTXKyTakdKTb2YFZPNtbco6SGYiSyq0BJL13t5/JX
X2eKhOJwLo+DGj2lEHDaCtCNSNMY0NkEv8r/4RJ/oyDGDl+D/MBA1cRqCd53
cCDunnCdbZLWKSR6wwufVe6Gz1asgUKZrmr2nDvsuhoGVdQBNpu6OhNPrjjY
w/LOIGkW/oclRMkrL8DJSnPhPJxJ6yk6YVr1NbGEjXrvRbaQvHHWeTyyiijw
iq8miQ9tRZArDE/oOnwer5s9wAt4e7tLbwpeot2KAvCHnGy8+axqXnucPDwR
nYajg71iMOcIrvV9OUYclpMA7Tq8lLtZ2DbEzI/b10oxMZcinMgh1paoXawo
Bg4b+uwVE/jTx4OyRgN2VL0Yl3nhHfkM082k8TWRg+9yv+oQR+S6SEe/eeda
KJFYie6PbUb1Mpw4sx5dOr6lDE3erdQ09npzfXTyPYvaqjhon+Fx6wA5w3o/
oTyuK327taNN/cPPYOCjPBWbSx0DTC2QNviFIwu0reQw3ABQq/XwHBw6ETem
JPlBr6zacBlWqr9mgOgh3Zot0BsxcY4re2BayO/LRZ3r9gD6ApyJkK7gMWkv
c5gf+dbJxV7DcSPGTzwdP6W03IP2Ug0gO4pD6tHEb2GFsbIGOiyZn3Tv/EYq
i1gfqNiT2OvM6eDddJ2B6TxUHFQBaS+h5fMm87rppDDAqjVmedYXB3x6WSoI
cJrHADqldcxrsc2v73xJ+i9mx4penr7/esvxRJNWv/AOPOPE7C7qasy5uYTJ
HjlPFQmom26Itw5Y/Bm01fAIUHBD2wRWCVyMz+EKrlM7mfct5mIyPX3plN67
QLU0LbjbMaKzrATA5OPJxEk9TavwLZyIU6Ol1BRwbeiHMewnItVIV3/Idv1n
qCcnn49N5SnnhtGIVlFC3ppPi5Q5eMEgWupILYcEg6ADKE83NQ4apHWdonj5
T2egnbRhctT3Z2gLgfZPZ2BZ08swd5zrjTb2FLBRPtIZstSJwufdPGe0tpLl
/u8czdOReG16dWp29jGJoaPRwhIYRFXCy2aotXItO0k33HOJQgYTwwIZS77W
KDJ6SVezkBtxOLVYkAbOvB8DFeO+fMUOzwbQnTtly3j1NoCh+Oq87OXl1DP5
gMVRW9YxnRrAvkjiX/FGn4OoBXyoJkoW0Er1AABVHLfNP3/eweEQaouC9072
2hVxGDfwtNnLyMPWhjIFKHMAXHOp+TRG5eZYHy49jQYiKqjqwYt8jEgzNMMn
DkyM40XBwqJV2ddjzfb9NTDKrTdn2S8K/FLXJyCEIuJvnw5jcuXk2dZ1UxPM
8Hk+qTRmQy87Iuml5ZYQN/qKvCstRyq/hhJVQ+SJJdejYkTDQghMaF/uMvmO
i01b+WWQzpfCCqeECPURzOoRZw0xLCv6hhqb9JSHJZ2RNFBWcEqbyL5wGXJS
HpdkZ+3Moc8u6XSe3xwStVVS4XjkLgCuImqV8qeG4SZZ/MZ6g6XbwNTC6lCa
iVYuX5PU+zoY1LbFaUkwbgsujr5Weu7wmioGfIXIpnC/1eYaBFrRsY/pf9MN
/vNEsw/YHOsbvxVVlU3im2bCWUyU3cCv/Ktaxy78v5EgLABUIpdFWaLdupdc
Kcv02E6KigBW8tB80K9JlOnhnZkJ6XclcLTjhgRs5RO/3U9QjYXQblAzIZYO
LpgyVeBQQy6iziT6b5pLOFK51NPPOKGfF8A05hs5aJw2aAFRLusotlZL5xvT
vaVTgZxIgqUAoI3FXZHWJ8J8aNNKpAUC2JIDC2MkQUJXTP/wNGXyp7zt++pS
gK2IRJkp7ADHbCP42hWPdmL7MTYKJ5u9xFK8202H0vfa8irmHFtEEhQOj8CQ
+MA/YetW0Upv/C+x2Q/mIUHSJA4eyXFXp8rqewkCQGQ+JBkw//IGX0Ovg9bW
uDuQTylapAKw60w0d+7KXjXV8Xuc2VdLZXxLE6C1xvLmKMMjLTIq6p+bdkrU
mpyL2N0wxj2rJI8S1FhY6pPgnNBkRydPcSvSPo9WTrnMJboEvd12mma080pO
Goz2yqOFXQELjpafKPdR9ObIVKPRN97sdd8A8G8Ee2rouGWY24BICSj2dRjG
UOZtMxcUuzuEddbC9eHCuEMqu4Dq/yOJ05dSTH7BRmcHorWd9/mYyvBvNHnr
JrbyC6AudjTmL+C18aaBoec5o9PSPwmNbHteWFvz9wvVKmVG690cWmnv73PM
nhJvYB+bRawi7aAdnyw1nrpXuN28g2ZrbQVhB8ulgnR1yKWcmap1RnXPLO7r
KZNVUN2ra/GwODj44ECengv8D2iAa6Gf4A6eLCMb2p+yTBMutabxxEzDnsec
fmQ39bQ6vnJO6fIJ0a9z4Jfjh5YDXA2HjCUhdUOdlGs0a+expJfERQNPhsRk
qk5vJZCT/H97CThH/6ABgqGdJzwwgMMTaJYR73wN0R0i5YNUA4RWli1GwNvQ
DQwlogC2V6XfEqc4XhMSSWbpZ3ceGYyMmE0j38fp22yKyS85HOcCsQAKkjyW
GyWv1rPhIQ4zXt7Rv2/QkcqmHaLLGCvBy3hpfKEKQZCjimTmwKy8y0+Bgbz1
pdM52TOqL+eS7lfKFvFMDMiQJ8ETrL8EU4kG3/zbEQjieh8vnvRAVNnOIsrO
3U9p++dtoUvDycvHI11gsHmB7xEQL+VvnElPkL+mqAlfDUrhTQTb9n7AVDIG
gc3MCr3kzR1+qk2y167+pcEANR2WiVuUBtBzdF+y9cuDLdgqb3cCX0lhyu95
wrYsS/8Rq88Qj3MlApC1LD04/Z7g2NUcw7BNt46J1rJOwRN7wSh25KhcR19W
2cujGLy53W8w1FP8jT2sF8/nqAwn22JR//nUWD0zcCNxkEwE/zt7izsCg5Op
J7ItkDCTRC7ZtCCyGmtEzzXBuNnFwy9BGhsRtoPjPc6gaAnpdOIi8XEXo7IJ
Qu4H2PQ8EiyV4D4qcAEDi8Kwh++eYuy+X8ga9BBV9OhDOc/ZlUFyrHnVrHvq
T2d8ATRoRFdkain54QaLupi/H9d+2RmnJCgi5Q1fNtGgojZzo6XPVfpUQn8e
dDiVhQbTClgnetfJaO5jPaaqAIuL6zBsLtHgQYITTv3BzlQ8XJQb4juheA8H
AZnpY/pvAhlIvj5pBTGAxLFVVK2DnVVOAmX9NnjsHwy3YPXlodJSaTntp0A+
Mp3WN8ilsWB5xl8mxZVHxROZmJn+qQsyALQKjT/LZ98wE1mtsTumpD+8ee2A
Ro21wW2YWsHXYR6TNVGOLsjRa8XbYFUnpYZt5SqmEMjyJntcAx9s6aKsT643
Qu7XLGHVyABSDcovTBigHrOLa4mrgaCIGIRJX3Pd7jtxAq1ka8+OJ7jB2WmA
bz3MLOAEhompAogIF/vqjKGtNpJ7qcEDWXojU+Q8NZCN6gP98uLtcL1PuibA
VczaOPikXqMVVyIfN8JnG9DcG0tFaF/qNZGR9P/AGPSv8eonbNDgz/wQjXyd
ypcXJ34jp/GUOkppL+rHy9gdNAiqgSysxfgrPFbHR5MKC/EZfruezU2bXLAR
vykqlsxTJOw5A3+ij/Iu0oAZ6Y4/nqzOTthsZ/tvm9eZKiups2Z3a+G9TMge
48pd1TUU0rEPSPojORuUYCmPVBYtqqLdGsA4ZCnKWNkqDKRJn4f70UMXQ8rg
e14mKTI8Bk+nZAROjixhZ4M95II5Y2Og16VslfwO7BdGvvLrihumcfcEKpnk
rIT2pVB4Q4ffwqAKsv9GTXxc9Ce0MV8yvLYNN5Omd2OXKnBtmyc4OR35sGlR
bD+bmrs6SNNzrB5we5ImuFgzElk/RjvYzV+5D+yIg4QugWjgnwXgMFe9LDCV
GAfNV0dcwZrcrM1vLQxSoQbxx74/ucRtdZixfEDRYS45ULsmC0KCtGHCMxwF
ExjGvOkINkjBbk23mKHSJohULWsN2C7pxPGkqszvuaD4tajyvhev1St1R1rb
BpmS+qgBlpwT5WRRoH9ZJ6i16gSeyEvzfKqVu8NS0DYZ6atHKELL5LUoGBnH
wwrDNxI0ZD1G+VPZTeKWabdV+W0SZ3Ef3WykRKU7GO8PTM12Wzf9eN9iRZkW
dAflXsIRuT0jOhpKqoP9EUYBalEAtVzgVOKsp6JLGoCyysdFLsdEtKSbLncO
o8hXVJu2tvYWiIWzTeAELAnsj0EBBjVXzjmyP4cvhCV9y3uOWkybi3654Lm8
7asAqsrVMIhKY9oZhaO7JHVtY1PFATyKm5m0yUZI2DCrwt6l1y+F21aeUy5+
2Lq2wcb2O7w8CJgi3WUyXLBodP8F7UZFSYlRkrCBiwNqYxzxARLCMalZhKqU
TRcSYT5ZBFjt9skXHPx1A0u5efzv3fx8RvaJCren3mb9UxxZCIQgCFIua4Re
xo067GOlmF8zEHiTXT0EmRdtAP7kJRqu8RDKezJAOwp9fQLiECAixnb6zr3e
IrBRzU3L6BmMBvpv0ZaO8A9y6KPK2HXUPDUC+HIFjfDqr/q3e54QvG08j041
SP01rESYqYwFW6Eq/DULQ8GGNd+E2/dATZ/ot8Vikv8HMR8ho24Qjf/8PdJd
FWMovD4ZsqfbLz7aUW6stYS7JzK496D1gsif+NV0zUjz11gPHovWefpIBYkz
egWXb5DUKbvj16+r8NMKJOowb3GDAu5E3T5Is4tfx+V7EScdEm8ga6rqrn6A
00JJsOEYZTwjmZsT4uQBdBANUsd7E1k81FU9cGDQZ/fGUH015qP86IKU/OmO
+Bx/1aFSfIPQx8Pehu4MVhgDaKrZ2jHdL5R/n50ny19QbiVJ2YE3iS3fzkEu
YvL9G4JmsPZLeZDdgiQ4gHF6GDkJ41gCzdCe8SebCjVul65iDZdrfA2Z6GnY
lpT7ppmHwf48RBP6FljkvGMjeBatDhxa/RZz7dXcUQk2P+bpbtJ6XyrhA9D4
X3L6+7LWWVt63n2x0g8ctxDUSNi7wSl+L/8HqKDLOuj2jPqwMjhrTFHabQAv
jOawVJH2aSF4FIvQ2eIshvgWOaDCds2FxVg1ZJh2t2y6dzChgIQlBbfEoMHj
5H6yYxmb7VleLisjD6zh1/plZUCrsAmf3JmL5eJ0S7j6D5iG+CUjK6YcyfbF
8IbdaFjndit6OI+sE3hq6ypdH2AZlrfs6LIWs8kCVlstx2HfHDnP6ZJxCQI+
SKHkCv2PAuXM+ynnlECswHH2bHy5al80Ru4q3k2nAVh5Iubmkty8WEVI9AOG
O3p/S6GRyAMgvMl5ZQhMDcPDQHMWWwjAlCYuqbc3keGWuz9ow9Q1Xa5xUUjZ
ZvPB1MrjEDS2bqOADg4QXe2NwrElbQZ5gQoFdXNqLkoPfkWzGxUj07bdbPev
WuH5jaK9XVQs9PTkN2jUv0+AZfKnLl46/2r5ydWXM+Bp8Ab9yWldk6Xkkowb
8kNlLAoDQp2dql03XM6uRwgNUzevmOKhLvi2lpKGiMM2fOkp5bmbu5/vAIRX
N6FnSZGNK3fMUQ/ULsKXKqS50XMaRpCW0b8YUvrK17V7IEOxsjNrRqT/C7cx
GH2+j7b03wXfUT/wa1DhvGeei/va8OwCAHZHNMztK7qJHLCM74ks5AZPKpw6
/pZya91o/qcERxvJupT5b9/34s27i9k6AJ4oqd6I4JISb8nmmsFRh9biHso3
cOV6cOXnSIe7bbN2fWNVXB2j/ykwzMi6lXfPwlCpUtaFn97Yu0UMJL/gb29A
XXCzhRJRadnCioK5z5tv/WDPehR5KzJwxV0sVR4S87xsWEBag+hEXBr5t5U4
870/gmwQuXEA8m8LHwZe5rnK8/v5yEM6QMnaLHkb57DV+NAh8LF3IKZnPdp7
2HPyen+eOAOH0LFKaUPm1BAOOJJ7MWUdSUNTygV6v4Df6pp8UCgqz7cqqag+
97W2EAB+ynYPRvsZkzzkBCJ1jC3h7HimC+A46pciOVuUFUHAsjQun2/kixr2
BrjeSpyI4JhVafiLQe+2iYbPZTHjAXD2RwyAwgQB38vzfY+YE6Ds65T32vEh
/2tWxAworVu3RGIs5d5VJ+Ew8AqJx8atCEAxPgKqDB2LuZwjaaSPygULZXvj
rB3CRwX2KSONFlXbHhJvOCUZWrua2LN8winmf/9vJKCeNl9Xvb5Cu6IsI3Sq
HIcbCRM1YRjPxITUxbZZgwp+Yk1Bg8UR9VXtT9ABPm3ZiQWL6IFGd5Ugf7w0
LceuL47nXQETafIcL4xJV/lCBeVNa9ppYX3/ks3bwYy6WfRbMcx229AsHTnN
+fK/Dfvb2BHSfj24GyVjcsNSqDF18kDBlcFucKurN04asQgKZ8aRairrtJgm
d1rqVQiu1BEYujy2qQdO2Y15XYpsKzreYR3Bt5EG6IY+13Rn2+DWWI2qa8eU
x6iHJ3YSVoFWiJnZsealQao0nE7oiwnimstroF2WOPtJF2udRClCGdGYkI8V
fB/fnsXhadxNNL+ucC0WXbjzuBZBR4Xyrd/DvzVtangWOVvHueQ2XBZVjFFB
eCbifZfdt4cOqJFcfocnKeJw1veGOq+W6HsoSVzdTftvtAK3lq5lijhocXFB
/oNfGNqngUFOEhbkHmFE5KfeWeuBohwxoPRYOq3A68M6BxZjUgwAc8DD/rNL
ndGw1+KlKYO/j/Eu1jjB8LtIvF7Ef+Y5GddK1Bf59zutY3ZTlHet9i0X1KXr
bZ8qiB4jr67D5iRkV8b1QKPWIDWQqy0v1E6206zTLItsjsr/BKyH8/cOE0+n
ZMTwEOsKL5kjo4cuwbChgv4I5nh9coEKqi/nQ6VCak47Lvq9bl86wpwpCMnG
1CsArW+MIN3fxyiWq+uOlv/Q9MMVkYcDmW2qERn9fHGeP+00vHKhYF8xa+Ta
myheb+W6sWQX71piA1TBx7tHn7iTm+O+zcjegsXjSpHZSMZ8XMljcNx7ThOC
4G+yLLt9ETQWn/alRhD1rae/Sh3ksnpLN84Ly79nDT/LmTvqpf97ycGuKHt8
0Kud6Hheba7dbaufBUV9h8qm0l+7LreKysdshZsLNQJ6UMrmX2zGKkNpSFFv
CcxUEv0FNgk2F60FT00YVDSZ7cwx+XSI4XsGqBtAvQV0D1nVV6RtZToBV40C
xnJq+yhxdk6SsGP6ow9YM7WlamNeAi9OcGD8Z6YkJVnvSwQQTAk1q5koFhyk
9f0o2QOEIaBF/+orzAWAT1WubpAHQ5q8jRZMGXYNiEnffbbNPe4QyfSdhs0q
eXPQdvhLTKBKBBlB8ZpX4ZckhIc1cL4KC0DPNo1Ryrscg9Cbm22wHsR1vEDp
9OtGhAWHpFCDYEjQiSuU5f203opAhA2pj96toepGHyRMZInWqlft9cBZvsp3
wkOBMQrnELAQ74K2jTEOlY8YU0qLuZAGI55QZ5om79nv8/nO0w2Cyrn+UmOi
63rxV0mSFmEIunVc4RySGSg6HyzLUAMLYUYZV5xYgjH8j+3Y5oPLhS19cVLO
6+KxtomEfifpY3EmT+cLW3moe15YEZBN0IT9xeqD728Niblu8yuyMWNIdEH1
QvLG0isbCKMOsJmj3byxmVvFYizDUCZ4lf8o2RMjyJg2QO/itD1kDW0a5Amt
gdoCqvV3NL36yC+m3OD1uo9uZCns98lPwHygGkdl2aMfyqxXMQ2VOkeccbXL
msT9YyF2LFoN7vlxCqn/4zLq8y23eIfDwUm/SkvFWnKyyPaHLR1Qd7ZIuXV0
TX0NQ7bbHvJFgptKZLOe2Bw4QneDAMbV/cODhLtdaYDKa1Ikfhm6XT2BF4cE
RfRO7oy/CAyHVjNaZnkbijQhVYUWROljTAyc3Fz0/PytHLro2v/IVnQLZXQb
aED5zTNzhmHPEzlF2VOksJZXTCsnGWkopFWCT96plAzoPgWBHu3UvGZuhpCn
vWAphp5WaIbz5O+eCJIkkK6cqn/vmze7Esyi1T7DyM88vUDa3blm6r0BAVhl
j485NNRzinc0WBP8gNU90QYo3oJdI4GlW8CL0ewPy4pj4fdq8pGkcQR4aoHT
I284xNKUZgNvRPpBW8UR27EE+wozzt0RxJdyd7sHWff/9JmTLvwYyjq5ytdk
tanCl9TCQw9Brq1eW4er4OmSA8/sHxp2IcCDUVA9kp/861SMNuNrMhqOp6qB
m3gRe4HbZ7eD3fG9TRtTn7HQGyZ4OUIygbPBImXiubtxVl+Cey2lbkALBTQ/
C/DNQY7OFL/dnfciI9uA44tWj9b70No8qJBwn9BS6O00UBMmvlEK4I4mGACQ
T/9q2KO2UHVZZZ1cjgTeuxZxINL5ql4KpbSUoZcHCYZ34t9zZqFezNWqBSaf
qnMX7+5Vc54/lQqyhUolI30PTTq2xOQdhqjguvCHSUrt1abo6GyY0/FkN8hE
nDCMMQmazj2Rv9o8pMO09Fm0rGxqLnK3ZXDpNmG2yRP1OkJ3kXtY1Ms1kR/E
O4GPz3bPfpkSN8m8DNjGl2ocZ1lr/gKoFkwhjeXfKKQw5q+TvFXSIXBb7ddN
YwLmLVTxh0kFgR4hgb8RTqPvstFR7+XUg0f/UzwfYFujqLnblc5rY0vMZYhl
6l9h4TLKLn/iDGJjZrGJBL31B9/8Cg3RhQoCnfTADvAu78gvRzuBiqORPJmK
lqxq3zoWD3WIzpeG3GsYzBmMTOomPoIMM1hRTlw8v+BtnIvgrKeckPZUOhH3
kuXq1kFsHyWmAwi4Cj8+Pn9vkXMdGugKEIj9A4UEwF5CWJnWEy+dsjbBw0S9
qXQbxK7KoLYxWKiB4yU4iaEVNT4gQXfBn7JECGgCUPMyA/KtcAGDT3YppGz+
M1AjUPLAqAn0d4Bvo/bP1IlZKaeC1b7DOJdXvTfGOGuCp3M78gqnhKWru+8t
8Jh3RrhVwd7mMYNRLj/vLsTB3RgVNNNx2krtie36d41NlWFWdQkQtrRY6qh6
LnwygSLeZgUA5O2jgniZqImjnkSg8U6hLeHiFj2HTJFdzovkY2ZmLHEww1BU
xSjWV8Rwv2d3Cfqe1kiyrFcBHmnfMC/0BdaPVBr2xGf9L7tHpweoZ8qzEhwp
AU8HdXzlhEjxCzBmdD86/Qj6Te6zUcNrLdlycms9uIjmcqGIB9XAsE7dEgGN
NdAo+b/Oy4I8fNYGxqqFgab7S2I5d0LVQt2e71nB4g2RWP8HlR5dMTADBtHn
UI8LYk+QNnDoeM0qjA2ZDlS6tkeHSd68nQZ1ncQUgUuGh4KB4LEz4qv9eSVG
XKXlQKPr7hxE1ggrkngQgIzupNhIolzl+2Ym9tjZ5qq/cqHk4cqWwze3SHiX
+sgqr1rVYqinlJJocDKLa+l141Zj/zC0dr8yra5DClf2C2ojRjieQBQ8j5+3
4YDLU+pTx/IH0fwlUa0/BVQBc5ZH6guKgI42PAvym1heZwjn1wXo5FwNpHdQ
VkHmzOf2V295JKbC+95WP9Y+xDQUQ3G225JmRTKFZi1B9mvSOQGjSvlZIQp2
fWiVzawpJ11aAPlNrxCMlbPTE/Cf8NBPbySWfFH+Puz03IZJMxJO0/sBLfhx
Kmdg20NsCtjDkRGz1l8CGzSmXZY5mYJLjVorRV4nnUrHsJW1rshckTgoG+kk
bRtpJpviVHf5sJlAGl1KgLijaODiDrSX17vn/WlVPr/jtNM13ArrjdjgRopU
Y4QPf+pjMY72ITIt+Hcb278z2V9r/uIdGS5wfv7FJQ3pWDPTPDemmeI7tRmz
Xz4Uo6NfREnqO4rFqYW8aScteqdiWDCSOzrOnCiLhkScODRYr8afctx5AFG3
gAMjpimKK4Q3hrlTLfWpzfb+636oxdZTLS8ck5csczqR7BGghNN+FnuAhaBK
P6PaSqewWMLoL0+KF+fAzstt2r4PEAABFy36RSpZwcZDOd6JKgGdqh+4M+Cd
qtUuurRA3BdIub1Ute9Ux6Y4BHjj2mbSXaK4ajspfbZcU7VixANlnzPj17HG
8HC5rm3xbbAPK/xbUj2nsSWYj8PB6FO2Qc1rRgkt81qS7dll12RBQIGBnYtf
Uz9sYHp0EI9ytOxiWbst4zSVx3TDz3mGCLDFEFsYurMW0Ua7jzX/PZ/+lQP7
XAs1Z/STymwO/qxqvSFw8CTA/j93pdGgb5mAlW4AMeKwDWxpL3xGTVlsM5lg
adUrPXU362IV1FdDD8FuUn1R2uhjd+TQqXQk6m/jf9+2NiRb6FObfR7MZbfg
riLEhMWheRFrYnKvBbRgZ9psg1d1PAZdB4VcjA3w9En89CNXVhWLBJK8JfX6
oNdGrLZ33OSn4oXIIeOlMoCeBTqayUos6diz8GeogiTBWjw0nP1rwV3RDggx
lBsZb5eeKVKYN7HRDjlkxThORorlAU0mkoYXCgByzfNlSd7hnM8InmDpMEX2
BOiySyVTZzqeDALHiAdNZcqAPsuuXQKZpZPubWmNQTR3VmaFSADeN4GKTftg
q4+ypYfgOK3iyDiLEajXR9GxpXWB7E9pmrUIeheWNjhCQ7bZ0qqV5vBzeS0d
YsTqlED2vQUsT7dUkUKmhybqbw+NVCLqBragqWVKyI+TO7rKnutsOANXpV6S
+m+N5Il8LrmtEzt81WBBwQGdgc+dStO67GN3PCpQ5RCkEPLXf/XkPi/gVt3y
1GaXfWyxRcSiTC3v4degue+UpK3SBACsPOdXEaVePocv29gFk8wpS5C53Cwc
GrVo4z3bAyxhBLFEcj8T9x1xMyDBVxi9QHaSjX8ao/8vZ3zS9PPyExHeHDzV
ah8oU0BA3oT+ENBon1ghWkeJJ8lxYYp9rkHfolTA9N66qr7KXwZ7I5IaWy4o
8twBvGJJtVqjCcFtLJ7vCWYRKjyx/KYOo2TFGy3C7HdCEMtSnQLUEz5x99nH
LgCfa53Zsl5Q86+dylsgDSXqz9uMxM2NZeFEwMedpEvDPv5ctAaS/2hSxj5y
ZMXi29SOsq9WC9AREV/t9hOWZCxDaVopE3t9gobrv24ZPoHDO8v+wT23ZbqN
hxgtKqSiOvtw84AQFHTmPQXGY9Jcey6dsWvIW1gkoeDor1Gi2x+Pk2TcqoUw
ojAxXRHLVAwLnMLWDi5zcvjX6gLp2WJWkaknjtP/crhg9hj0dmSyAlZ/47ya
GI6tJMzsdDE6Wkz4lf8RdRcG1Sr2MB3Bklz3bJQnPmYWI+Gf2tJhCMIA7pq8
JrSxM9o35mE2DNZnOiNn3razINCNGMNoYzxyj1sfySbdLT3QpoImL3AKX/RU
lwhkp0YbCWACIXNDZYtzq4IxJYv0ePKGNsrb9DUAZCR14czXY39CPTtA9GVk
HL4IxKpaPd93lGIwLdB7M18ZyBgJQVE5kjOj1SrWgJ6UekAZD/0sGQKsolCL
+q8ubOxwI9m1bCl5mkMVWzxCywGj+0LYJVbVhjU7ciU326UDrdGNdrATIMyZ
Gt1cBTOY0DQDomdDt4CjAygZCOoW1qkXgwVdXjmUdfXDxk3sbdUJf+MqEOjU
RRmXIYLaorqTVJ7UvScexeGOqApWc6Xl/2KgeGojFFjzVNdHzjpKNOMdat/C
rcG7T9Gx7mc1lRBlPFRBdVefNU75egIucrMtUMFtbRW99vhhXikFnUhxEXfe
xk5yylap+2hCCnnwZtvdiMj49UfcQK00nq04frnuQMHVAwRXidCR3TZ+Kh6M
mqLXLFPil8D4r71+f7EQvuNCXBAxOhaBETwUA3O+6B8NyQTyDy1Bgn/KHhK9
AGic8n0Rps53RN6BwcJye/Bv1JZ4/ArmIBsTgmPmTHZlustgCXRVGTPwMRE5
4NrWuHPOk3tHivL8E+H+kL5bjEtrW30SNEoxpTkjryzqZrlXbDXKvu1xFiPM
gfVt7/S0XQHDiEhnDN0jGsfbJpLPdtpLrBWeVhVz24uSdkbc2NOcGFaF2AvR
tlRv7Pa/mIDggDNRd0iGws3dVp62fiKiyuHv8G4lnGDZbrVM+/u4k4rLtrjn
9iZZb1BeNmZoX3boRwZoUekdaUm1pa6kTPRp8muLEDg+VDZvUPzz9fgVBQ8f
aikvOL47WT5hnEV8+Wbrhy3wQZYxbSRseAwF2uQ951x40VmBIuc5QxgadGh6
plOBTaTtsENcK9GenzKk2rqbBCuFIHCN/hkbD5oLJLMcHCg/AdwPTXS/Xy4Y
do87vJ1KyBrk4FfeHwydUa7jzraz6MEsy1Dv9sdjjGjvY5PRgJYs1CtSSQQX
U5aIDkPymh3i+mrXlPGrxzp3GghSZlU+fAmU/n/GqIj61RR3/q5T3O8+vJJQ
AncjEVZ8mQpZrMFWNvjrxQIyRpYEPDV2ifAR0SXaHaY5CQ7aPrebPvygcesn
HKTbSYPxVxUcvkINZn3o7skBdUV+frA0x7BeYJrMbxvhLeTEOelC1abU4JiI
S7lsmGtmAsylc9F/b2wb7d1WHbBzats7FKAe4DIPZ1VRR1PzbuIjZrL3glEI
cAWAsttdvuIONVdZZmZ7CZ8muvWKfLvcQ4VPsR0kNkP2vwXvgnahrYHoc5kp
QQ2B+chrnVRDVkh+nlLxP/O8zHZPNxFNdllEwIZaAO3F/6+DaXswfFk1H51N
2+8zU2FeWlcwJZXlcpf7yVfn52Yf2s+BfMamn256CecYt5wzVR7EEDvTseto
rXV2lrq4Wf/pL0dXcI5X0IxxXaL2nMfvGasYiwmjrbLpEamf7iP0JLg5nTxm
81T4GY4Mc4bcCliN6QlDBSkTvw85YNRlcQF9QBWNBqQNgiG7ak0aM2LupsUw
ORVgnmvJ4OQodg7tQ0M1fvpt48sGcPlIgFFJLzo5H+g80DtQ2jeWxn1+Et7w
vaarx+EPDsmYZsX04+ACZmukvKXRc6cHozWy6ApmrwcgDu5cKcUYKquV3xcd
E/OWa6AxLBGudKx/seDu5icYYlvxG20J4npoMNRw/0/Y3QNEl6mR3zOzfjYZ
ghFPSElO7uoNeMqhKV7Ho4E7Zfr5T4Mfp8Yd+LBtYHcnfcTtFRIw+5Cxn2ux
3XlZBLdSAPowBTXPhDCaz7Pui7b4R8qzHODjTxu0AVI7DXZDZdsWkjHlwTV5
9cWqOX15ZzH0fl2LJULWFRGDG+iq7cwrdPHOX/DNlSrQRfvmiJviV1IhUd51
pcTAzjZBvjPW+eLSSlVlY8zb6lN2Whw14GLn/o2HaFGNuDYh7VKxk/RvsAKF
gKIAzs5xS2jEh9Ob16hqV9wGziLNK5/0DM3N4Aqz36K5PVwuq1XsKkKRe73u
us20/P9vKaE0ZrWMmd1Axmhn4iKhAeSHYsJBRyjrw4X8HXBCmdqIFS34qWtB
xzLNFmilbaCjgCwT2ccXPlNt3EwX5fRW/QZvCGPZdJ8zmZiBQXzdUSZpTT2o
olvbhv/IwPbi5uSgH5piWrpjpTdhkFatptOAoGNtXj/xGXIkdzuJjSisdmFO
OaOBBQXOcbZq58ZPbDsiQBguOg/0Yp76wFNM+HoTtILY6bG+W7wJ91KrV4mD
116Eh4qZX3qLAJ8Q65/3Hpgc/njgjZ05WtK9FxobEBEQN8TSfrev2wubj68z
Sxf8lXgavcNpyEv7+qDcQs2xuxb3YULJhp9+3Fyodho/3KJfNYkpTKvt9GTj
oDp4442lPzGkGntoRdaORmICC6OzupB/jiVajysQBvF/p1V+bH3CK6xeTRBC
qkWDE3dk42Vj6B8VwVMIu/AIH7wa6Bz6PpPniEMTuxq/ByzkqfQKncF+/w76
5KtWt3DkUsxJyVWI2ER/yaQ3sQaKrHtx7nmcpvIJTJ5xv9Lnv8yxMtd0lRKJ
Cu1XezFZ6OpqzEgt38SZ4KO7ehtgEBqLeMB87Nh5Y901pNOZNoamRezo1ulY
MJ/YY+MBeBjDd+0ZiSq/Xi0LGbDOMA8KEV9A0qiK3bK4PqxMTEDXhD/qD2JQ
ZMyrOC7+x0KH2eJKYyO0QJzIl8nc3ZTS/tKDJCkstdz/oyaXBya5B6n7ek9l
rhEc3HB1uUr5vMt1kMe9T+ehjEaoKA+JlM9GQ5xamtGCJ9lOBKmJvN/g1lb6
MXDuuETmBeCO5r9qU3XsZzHD+cWWSw/6gICoC1oWovBIem4FaGG2Mpmjyu1o
NLNTrqbjmqtSePmFhDMRvG0SN0KHk3iWr/MXbHiGPzhpZG/Y4appR6FlfUGB
+O/n9SWQz5f1WO1+KkZxM6MEYGv/bEfqGVYSkSG0zPe2whEuMxzueNJ5+vhp
4iIDlZnmx6vcqpdRQX6NdvHRJTmCcM7Ec5WvIqkiv/yimxsuYgfh/eQKvEnf
j8x4qYQnLb5Uqd1ejMeLfqCowp6kTkcg1IbBBJ5Dc6Sy1JYBpKOwFPB9kSPq
oJrl4yta6bglSS/WZqjwfwNsPKQtsb1G8nR+jktIBj46ERtTJcaNbQG0buFP
USkzlhNSFbIiaylZuAGibPEyLgXtjrMsYvVXf5/DSS4BADKkIu5lTRZiP3lY
prq69C0N7eIEE7VwEGMIdYLDgYq+XJkUW/bHc+fL0I/NmbVV4PR1i4NPECVH
lV+9oELCNy711DV4WcFOJTROrLe3VIDV33jRnRBYQsBfcvtpX4S+X6BXPOyq
gmpKxPgLy2cvC7eTlh23Sp6rRpXBGYxnrLHe0YY8BY7cmGTV1D0vwarMEWUZ
7/5odlzwB9+0qpUktiLFTOjvonNVZ1VUhY9dBYSDtgGf9B3KbII22DHEL2oh
nWNYFe/jL2BBlzHS1cYmgMF5WUlPpUyPwrL0HZFLev4i/m2fZQVMoS2yaMRK
KlmLvKyDgAXL2Gt5RvkutM/J6O3Qhp2ZztqrfdtzlSoPJ1Yz7wvBEGPlfWKP
oLEkUgvKpEGsRsKF/cMwxBi5qkSJdVjN6l/CvpiCk+YyYXykYnBfdRSs0emb
1CMFV/nhM0S5UmwURZu3u1365lV24ufk2/LCMcEpAOmd7IvNBd4wV0/Gy73y
hoAevFYyhihQgyHr93EvZqXFL2yJ33LrvzLAp7zWNXX3nMGIsTBarnD/i9Xl
9iXsOwKeVSI3W7kGPh5KGfeOAOkw+JFahNACr2UGLjKjlHUugLYHZHzCh/5F
1XQZ/kKmZ4AWcfT297Qjh+7DSgTrPmN4FBsJkI/pyZqcWa9vb9ZGKFHIoDwg
qoajb9UvwraexuEd91fVTh9g11Mx2PChGrJ6L34HxEZs2PySLK0aZojCuX3L
F/qYiGzTgz+Lm2orMa6ba5oPfNV1vWZPaz0wTxNOsZpPzqjuDd1MoNXcx6pk
0ewOVTJR090cEXBSNgvAoErE9BppySSwEFB64dpNL6cWUamwIkSIVORmGzGS
0RQQ/dmWAJRFASSLHdCu9X2nTWFO2uz/7l1rNs9yiGP6Hg+2M3l3KgnAp4X4
F1NDuHfgM4OQRa7UDDtW/koaC9zBNvcQZtsK5fuhUUBnhk6JheFXAtlMwPzF
FAdfWavfC2kiLNed+bPZ1ddlaDzC+mkjdKrdKPOdx49Csu5dd/kK+Q1zDPeF
LGtLNFWTJvy98FZLBsieYBvfciExFHF1ct5vlJFsPkp/oTCx/msX6PVXQwKm
gqpmS6Wxi/7TY3+JdwwSVMM3xA3OKjpG2dpkdoY8Q28UlveEGelNP8ZAz3TT
rSWMZldOQmtuHl0dVebcY81VnQmKVW8XE5JHkk8VRPKm8kzqN1jKG4ZiT+aR
OQrCeJxf/GbWaRWUpkd83uE81h1yuJPNmVcFqQ6oAn94c72XJH3sfnHEaDSB
aZWHUhyHT1olWMzrwvB3GdNbomqREkxLwsCqO4mlCAnEzDeS/JMgdath0x42
pf9wfUXkPYZAIWVVRXLTZcF6nHWiVxi4fghocaKBRlNu44Hy61MWFHEEzxNg
y8dd80ISiu/gtUH1YYxS9RcOz3BwphI84i1KoFjTMuevcqFEEp4wlnwrrUqm
+0K4y1TtW3R8PscKr+ED0WxpTrKvgWnFT8U5NEQdSXf3iKUe1W6Z+LnYBYk7
NV8OW/qmbDh8e6BtN1QgFmY6H3SSAC42I/UXl46tFUuF6oOx0JT0f+oXFAJT
jdC4x31xbEuNU4EYj5nKWhjqk4RaompHxeh0QTSPFJa4diF8WdM117mib2tB
7aF1XSbBo7um/qWOjSB5BJO+NqfBN0a4n4+kUotw3TOxHnszfQuvMJzR8YZz
XGUr28bf4jpq7HSpDrrxjwhl5Td1Ye5JCZY/e9FaYRcYprnDfIc4oczpM286
mzW9T05acvlG3JMJVzKbWs52nDlEyNeFoQhC8pft3xFGOTx007m2JZ0JAeYX
ciT9fluG0s1R4IGI5uNlORnWRV3uLe0FVAd1uNkHktv9VD6iAOHvqQdldUeQ
LkbL7hN43Z4Sbgvu6Id65708K9n60EtIdf9agsBHg6xNy6qj8Fyqf9IGacX3
79MUPF6kR+SdM32qqInB8TsvXnzQ/FBbacVvJF/y8E8FTWc/fLxPl1H9yFwW
agQ8fvRQzERK65ZmtY6iNywCmoI8hiInE6B0JTk/vEiBPJ97VvnY/fDhXJMI
v0rD+lHq4H9E5+9xzlW89p4dJJ3kFDx39OeCwoD5EIVi2mlRr0fTJ5aa0IL2
ODgnc12fTMVRk3c1wYMGXS1FgzR1jNEgdseMYKsoJMQFt7nAQAKuaAqX0cnT
utRtKdxTRWzVWhecLyhCBXfVMPvAVoJUFNNF07QVh2z1FWsA3wwcnn0jbw5f
/jujHMj+hBGwbA/NaDcHpK1jY0SuQMhoHFtmiAwGIlBoVefbdGmndEYPgrMH
mpUcA0Fb9pxY76XeRs6yw3nyMfkJu1rZ2kKioQR4yef1cdfOwhORGvhrrbtk
DU9sWc/STZEHULIg1Rf7eOlkcxYWElKmM21D3xpLECQ1psA90C1NaxHnqHfa
q6WvVkpRi8O6tpCjfciL1MSJmsGA/kTA7ojDD9dDPsuyCHi82N0TxOc5bKD1
WIJktrD8j6yjjP88NGUF24DPTn9jZjY3t6XH+kaSq/z1/DmNqfqClqDrW4wg
zYtHbSrTuEioJAIniqSWKziKK7flpS363dbUzIop1rDW9+1c0K/SprDtsien
AC+Eb6dl/prJRlysRdHyku1kA/dRRCE5whNEb2UQp6FhLCTYg2vXaFOGvrWb
kxSlI+SumWfrkKI12XWUsaiuf5KhNqJuP4lZSa6T0NGs53Sn

`pragma protect end_protected
