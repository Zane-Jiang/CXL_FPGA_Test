// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
cWg390MBjRO0CMtyeOcFm3BRGKfSMJTFD8Ytuab1k8T5oUJZT+cJIf1DT+tV5e5S
oUmE5rL3OTElCUUi/YLdK6jz+q1XpTlUW+fzP+fqlEoz/0O0QXWsx/KBFNBwIv9T
bB2bw3jAOUWEUcWFi9AQ9a9uvEOYo2mXMdTPZY3395Yg8aZ3eorDvg==
//pragma protect end_key_block
//pragma protect digest_block
Q1qVfk8nkkscIY7Pw/4LGE8Z1Ck=
//pragma protect end_digest_block
//pragma protect data_block
7npd/vauVVX/pbi4+C0/pAsCfQCKaaQNa4VZTedMmOxPp1c1znOUCbr2Vo58GG59
/A57xMBud+71g+3dM8sft+olJVs07VwuvyPBnSUS32XjrAvR1ywRgYS3dkSirtiE
uSf0Bhe+uEc4s0iVTj7+mKBeu8oGVVSHIAbFXYhJF0RdoFTbUlK6+svkFmOa2cgU
Liq9YNBllf7obcnwiFV6tmmliYstkybbZO2M0idcoJvxxdfbM1zCS8VRkO0GG9p/
k5HTH55QhYwvc6KPqHODI7GiUXups7I4nHkA7VlYqcw3oJrHk77EU50G+XrV7qH3
+FgDabTSfbJ6ar0juJ/SluirHyLgyOKzLLs7HfkojDCne+xIxLTN7lIPFSSNOt+z
wrXj4oyEejRKunTziB53blDh8nD58kT9sivcSyP941ibJtauiayrYqHmg5kSPWSm
iL+N9yphPfCqbO97xTY+zyxtG62X5ee/ltzGqNKrur97gkOraFmt+0/x+Xj0YbdT
U+GOlhdz1y9jmeCkdKJcFJNzvZiJ9OVaq3sB90/SDUDE4bU3//xiqWB23AzG7lK8
I306nIZKYm+nD1t6tk/tSmELEJXuLVVzO9+dLd+r4WvjilKJtLrgbcinP29Fo1T2
9xZgG3cf26/ut2W3uZ9udoRxYI9o8vBLdfhg35wa5WaZYYX33tVJj32NHk8Woq+u
IRWMJWE4ptc99C9DqcdDli0tZT3hS5ms8OkdJ1GffxsOboQtoxKMJb7VD10O5iHQ
8/0CVwluDR/rLR/rBHnUmouc4TMZ+NHBnDJyHq05IBD0SxbdUDHP/K0SZ40LKj9h
ill3hrOcfh2UnA5tsb6dTaqZ0N4PjvMF+XRsnokUqrHXf861Hsuq1edUTGRis2Fu
QTuC4ZxWtHhsCx3cx6y/oRp3jFEzfF+aHjAtr93sIOqmYMb06V8wRJWPu02jbiND
/VS3T9Ac8h4jSm8mBnXk3hH49nd6RS5weDHEhnIAofiphrPbtj0C63uZhg0bvsIe
Yd1TVzijfT5Q0Fi9r4c4jnEoiisVJ7ceO4dOSa1GnEa2QAm2ovowP+42t80zPw1p
55IipbAEnHEF4u5asusqtX9ZfZQAwx8UjAqQ0zRteZVLkxKQE9MCfcpA3sFPnyEM
U0tpd6lOZF5s6Sp0VqUbyS5oHLbeTBQrsw0zIvrM+ZcvXipItCoUtsKwc37XKx1D
Llk2zU/kEbKPpOdmBtSD5Fo0Et/dGofXbXiockasAwTElnTgprJPAu30YjZGwijy
cWeIuTdPzGLepOxuFlIcc8qxlHtMIuYIaCYY4xTof99F4gVtgbM3Vlfa3owSRCk2
VkFv0cflpfPT+/Nt+ABi11a+vadBoZzjeBEkN9esiZrCKY9irkcqjO7Rj/hljuIE
GLFASotypdDqjKP+MfMjMjrwLjp+cI961H75MNtTuR5qtBIUIkW00ma7Y7dMnq6G
EZ5Ha0+c+9So+jZi0aOIx7qBBOVdL8UC9hs0V1EexJINu0kAYUThGdQc+OgjsPnW
dY3uricKvOSd45Lk6zpzlRF9hDmbljPnJIYqQGP4PdycGnPNDp4I74epCjFg9+0U
2tbNZBoKAzmNgZhiQi7DRtnyIsMTj6L/IcwXy+DM8AnTkI6J+fXPlJmsDM72kpD0
7ILyVRix5adkdWlLaLrpnxJGkPOQpId12oAl2HOg4YK8nlnKxTX2NG8ZuPZhA/Qo
5xqNCc6Z+3p//yLgUYZWGIxpGvdZx3Ubj7jDAIaR9kbv90xv0VdxXnQ+7+ilWn7h
pOmXBSe10Q9GxsBl4Yt5cZkAvCDi4tz268yxfWx+VrUjWGutlz41P0eayqLy35RH
wywCstCR8OkQ4FK1nu9korYXM8gjYgP6RRWpCZvKov50zb3wWPjx4lr/9xkx5Vzo
7SMQ2X4O8MIAeKqYN+VWG2X+N3IGpC7gRq43s384hNx+butOXd2FuXqzy2q/T7nm
pII6GH/IS9/PEBJ+jXColB6fSEJwXbfUeo2A4ZEXd+wULzH2Z0y1ZIwsCG0+sN/6
82zDQHNulkTEi6hVVoDOiy1f9x5Lhby1CPPVEl2a9IDOK/zgMlgIy95uCTOnOUGT
Z7RXA2zrXpfeJsWfL3eFmbp1UpRwKpNtNILXpZMomD6MP5luwn/9A32ye5MyvSmG
Ve18hfEStCl6gZBPfInRSnDy4rOfPjyfo3kYkuKtwYIJXH2wm7SePZb6+6bxnb2G
WNygJiGZMDnaNnNcyXuWnBKmor7q2JyzyOsgwyKzo0Hrbz/Ibs3ka5/JEHDet9a8
5Dd5BuM9bShEP4ProEG85F7bVExhW90J0GzZVh0xkfluje9PZS4DxK2h5qF9NTZt
c79AcxNNw7exBCxBqKFcvdrkXRS+Prx+4WOY/Rh9N4QDm6pA7O6ZBfiVRPpv0VSS
VF9LF8cLDsOHEdOv/p2dNyEBOmJ2Eo8rd4Zs53RsukKWZdKvNNKSl8rA0NuuN+pD
Kh9UKxNydtMgAtKYWAgbjATduJUVuwGsvmmP5zLlkN+G34dDM1rEVOeE0PUtcNV6
gbWayrdLRu8ULNAsAr23LH5T1cx5XyqLTtbho9ZRlroI0JRVh1d1ucS4HRyEMEoy
SSwX58Chl34AtS3KD8w0XjMhX8e5yJDL1TEwNHXQTEP9VisW/VWWaR2goY32QCiJ
DtKWv9bUZDQVb2kZKHPu5uxZbl2aiHlYpdu5ID8zw/O9ufbcZ0vQtft/y3Iu+GSo
Ri/ygdCU+nlRwY0tkapUfZEEo25wDY3QCKFl9PHayJ6fHLtFcjKioRHHdrHUrhbi
1DFonJ1onTZBCYzSckY29pwAC87BcI3sHXikz5NfBtXnLhoUrPAEZlZA+5fAUkIv
hAWgOYEKpbnYBTMHchzVZMJpxlDQk1Z/LMgtgoOxmBl7Oa952BFwUSGqEK/agNJx
ZhqYhunMmfL6CYXEjBtIWHSJY0pPefDADgZ8VtWB8Pgn2URXx7T+8czXCWMIP9O5
JrUjwQU4Liuzr7EQR6ik+S+ttKUg5D2OnMeL0hbt2GrGEA/tJ852+WszIFsOwbhU
IjhzNNwAbRVpzJw8gFzU8TasOHvWlqT7jb6eYt6UNx0Vd0m8XrygJks0OG0KkDp1
L+btzl7sCkD2XSIgL2xRk7pWQBp2hPwy2lyjmWQXLF/QGiJzI4saOnbZyZmAgD/L
cz14SRAc0dsBEs0avNyGnmFkWrD/+lIK7Td7NnfwewSNjmAMxhT5VEfgdiy6s9F0
o9hyRSjjC/kjn3srGJd/oLxUuML1983LwybvFnTRvrLJMLuVM1kr7uX0hFTbVKH7
DEjoeBObeXmRPQmtyKLKcBwkJHOmb4K3nrI3rtXzaMPzwaEiH45e7Q+e3OqTdEZO
/DpTZqbQHl6t5E/e7b3bIFP1ahKEDtwRBtQkreau721YBwS5gGE1sCjEBo+06t7P
0JE6GplZIlo4BoCh00Kz761BThToAB1IyFET3ks8NTT70Cd8V9FIhM0R4fKvvYXA
9jXJ8LcpT4wwhHitVUrn2c91vbXfvv9MWOhtVMIU4Pyoc7TS/55boy8z1Sk0qBAU
AkhTaZUObTGmLr1NpN7k27LWkGGRX6TlJCp8ZvwuzamU+ddUislesQgOmkqOSldC
ua6lTd0Q3Fk8/8SpsyHnnRLBcDxLcZlvmpTNNPksDcQnY+kI+CkTRLBdkHRM+00Q
j2CVOAwrdF7j+odh6YPExtlHkHOQDv1qLAZxn2Db+2Q/nNg13TZDUhD9zpmcgmOE
c15UG0/P6X3MdKJLxMvcQcL1DdDIH02CSlFoHuQJm29tNqS9vbxZO+zRbfE9Vw7H
kTez94VClLUKiqaDzZttnr5v4R3m9cRhHYd2yBWmoCgAvbwIW3ULrVO0x9gDXgDI
ktQLzmC/V7dgONncgDhxiQ1dsRaJ5FV6ZjmSTObT0ty8UPZQ9ow00AY3AyqnPsu+
3jXm9HaibUYj87gydbytxuAF6ZgfSq0vyTWWKJC8x86B6pucODhA+vpMPRZxs2Zi
vGM+aYSJVy10b6RzRzTNQl3z4dZ6rPjqBq+20VKYVTAG0taiwQv1Zoqh28Zk4JBH
ijIPQ2JVNAGwBOtf55fz058YnsOA2ICakZGXVT1VBU5c++ad3TUeQp1y2TPGP+c0
VFqKwvH+bZMEJVyubGiRXgsjYwe6ZY9orXCqP98SJtZacc8TGsth/wW1x5eGNcK1
Bx7TQQTVacWRLBQRyJJsVuPdp2vgDqPZX8ZMZSwFU5DyJx83pduPTc+fEkPCSqAl
m2Diy8+Vva7yKoZrqNshp929a/d9bViPKQXE7X8VoXMxfYhkJp4Zm9bdEqzOw26q
FTlLaS8nAhwl9RVk32YfOHpOfQmENajCMgT8XdJON6p3HCQkP3wgQA6yfyivOcQq
h6WgPxxpXkDzRZhgu1RruLl0m7zMkhiod1YTKluPfMrQ6MY683W6vkt411gkO6bf
OMmDDHQsW3dohJ6L8vTIUPATAxQP/WyBliIXV++y6vltZfF/bbOEz/x6E0/iurv9
cjo0yVteKsFEj7s6W05vHkTXRYgpYOXvaki6mlZXO4KCfw4eTnQ6Cc9NpC1dq9la
RZQ/qnE3CRkGLrWFnQFbo/eb8OE0t4/F3UdwzV2d1SojI2JD9SYxGgUnee4S/Uya
gTcFZQD0nnUCdNas+6q3Va/EHN1HTi1aclX2JmyzeOx32MitMmR1Q5IEKSBw1ddH
NjioE+J2OwvtfZbcKuIJ7OYcSKiVpYR+o+wPMVWRROpbX5cfJY++7+sEwtbvDZqZ
/ccBWP0L7xlHitOS4KAp56GV3eq8yRAZ3U1T3Bz1sukYh9JvxZdJBC7Gd2KLmH/D
J5P9dUMqtCOr/bd4MJtk4ZCnoMviyNrGjzIeggVhriDlhMcYcfrsCXjnnzmA7NQ+
annGwWTOh44AEp49mvBp2YX2LGKZBeOGSb5Ml3gR0dNv5aRzpKQsLgGScdPaqZu1
7WPnL0bNNSeB7QhodDW9+TIHcs28Yv3lIjbpFEMqevbbXiTAVfDNMllvr9l6rwfX
5+IyUT+AG7cqL6NGxRIpa6PZwjG/yHy9RgWzbz1r4Ld4En7597/TDU9fcv+YGvLr
WtJLQ5ocACK6c5yQZwGgBQXJCHhbfw5E/Uc26uio8rS2rUYnTBetcDKCc9vWXLeK
X+hWC6O78bzPaQCaemkQG6Ul0cAbHKihuqRbDEU+nWeLJi9RhSQMzcPchmqVhvw5
US1lYcNilnkJTyQ/ja/AiIWajeQskMhfqZbmSF3JHFE2s9+Yd34F1m1BMOy8wWjR
vu5hMlP6z3rjHqHFpygjxT8JuH7kcKafPlBHss0B39tU7d9n5Xwgoi5LTA7KuHss
MpSC3GxjfkiqO8ozmUsne1LXBli7U/zf72FS+gy9UDZEcXermOhVlbwrUMEFYt9m
fAKc3kTj/rCBMytCnsBP7MrmzHJZfVHnWRbzfmKYF4OtCCgGP1Egxt4EikrhU8nb
OiffXAnPXxB7OErQTkyS+TK1F6q/DgjLm+p+GNOMrCDrWir9R4gjgPpZrQddVQXN
QM9VLuoJMFKlHcR3FkQ8qn+3XXeHIt9Lsoi37M8XnFDPeGNyGYjYpIQP1DF+Hkf0
qLMV++5iDg6e48qb8zCXINKYwaEP73wxpJnQbTgLhoma+u8ppNOLavKmigGy6GXl
IF43nCSL5iB9UigR85qx1dzk4vF/3r4YPbnEy5NOU6nyLK30eWWWYkD/bStlLd4+
NKxJX6NN8utCgZBlx732Alqw6UZXHVoO7gLHZDqs1t4y512eYx4tywobNRSRieQS
6h1ShGX63OS3yq5lRreqhinNYEA3+defWFc9AXMfpjPqyWozcBF88pAqWHf3gEuO
Ufc0aNXTPGBuOXsADqTTqmeJdJZdMPp9Hbr43x8Ws+9RwDnIGnhJsMSY7/naic0h
0ADF8wzl4CxHghHHBzH3oQuKN4Y+LQpXFp4tzLK0aCFBjiZjkLEac8FNKcGHzxvp
jntH79GOelIgQEnjG6Vw2CFlLl4Li0uIfrfELgeDzBGsNKIMs9XDPJ35VrbNqcUR
yTXSVAhstmSRJ1ALc9w0aW0j0Uily7g14+UfXt1hRhoj0/HzwSApxgRlELwxTT04
vHc/hdfwL7QsljPKRJudR29BwHwKFaQpCe9X6j4+rqWUyiv/dxtyxo7USN2xOb5x
1X1xH/KQBjggAvP+pkjZRGYlK3QLZo6lFqstcayqfOcBrJiJCBBYqQ8RGCrshQZt
qBG/K9yOSBO2SGI8M6+4SpqXB56VkYkvjNKqgR/d8YCMtLP9rgGnDMTioJEO4eb7
AG+l+MbDwpaCu3r03KOi+NJnIkQF3Mh2YZR/IlLyRH3OlWADKm/G6WopSEpjuQG6
xlGPvucUnOeIMtApRtCaiaiqtddcbMkp06vacoBtgxUbOuKfmI35BK7c1jTkaoU4
IECyCN047eObS+WIBo8ooKj+dDEVzBfcuc7OLZ5bWK8tp7zzyJIM0Fs4u3deRb6J
j9xQtOeK78LB0Y4V8Uv5RRsVSNe3zh3TodD4jEUwkz9tnUu5eZDrWxTUna/U3jlo
10f7IkkJQyDiGUymW3GWdlfnRHc0h/ZaAE4O+EF2jlnjHR0olYCF3SaMw8JGmzb5
4Dbj3vchSXyt0neJwTR6xGqz6rx2aAQOGYK9MgCVi9xct2Qx7NZF/UrDZKMCK5QF
/DWswZFT8jYGjzJ3mcCVTKG2HWEHT0LplOF3Q/kSskzgAkwU9YEuy3yPboK+GK/u
xDTr606fRrrsbzV/LMCRXWlv9wcXKkRxO/Av1v17pwTRMWkYVIrv5PI1Is+u/Cie
noQVyhBQ3VC8GkEbzwJ1jdP3bbGMGo7Dcgzt+LaXoDF6vfarEgyem29mAySe5pHF
HibfczG3ZhktQdwRKT8WV5AHX//ACgodkQH0Zud+bl+Es4a4ljlNLBv/Dokh8n4h
DQ7dVxORPT7Pl9YgvLpKRBxMqXlOF1o5tazHf9HWafyAuY5wbozh7nmVUz/TjGKQ
VmkCKkU56VmLxijO7r9x44J0UHGVjBSZC9w36vVgmfVm+4T2a4iMLc+NJ7FAlKsf
+lNiVrImFTgm5bx5U2Ht64kCUqYQzyxDgh/3mqKCZcZid0PLWG+87EgOed6I4xdw
EKKmqMsziGJpCsitSiktz/sPWbSVvwRVJZxtZkLzWHqGAOz5oxVoNHve5xgVDisH
JLtE7nI0dehhkOE/v3bIIIVwLfqVOp9+EfODhntGPKES1Rfr7tlcscIfQJiZMZ5t
+Czo77LUZFYDW3RPmhT6ja2Fl1VuSmlVQXz1TH4Ebcbpe9BODYVDQw+YkpOHGZ0R
rNU0yNoXnY3O7os3rNICm9Py3bSDC9dFN9qtaAzrXs4qQDpeFMEZguISKJ7DEq1b
etPtkHbGn6xLlD1yDbnpWUfzlRTfcNKsTufVDDgzBRCuEjNQ8Wu+JUzJlR/q9cvi
Kbfzgo8oy8s+froiBqbjvsyeVQ1w/3FQMlMpONgBYvgnYqFoP73y6vjjUmcMJc8k
Ar68PZ52NXbaw77IGY0yLNmb2CUD0HJ5TOONLDjqvBQ0mWxCag/mGc1cgsDbi4pC
e9qBFK1IzBppJN7fMEVoFsFEgcJzzahAfVXFZlPul+EvegtrAg2RuqD+dzMJtvZp
5pBgp5ErZJSZ6gM+6pSokQOoAWiYed81e46hpI5eZmDHwmyfSjviWcnFGBdoLlo8
W0/jDou2Y88qQ65koWV8RX14ojMlvwakkqcosIyugohKNcpbrA0T8zaZIZpXQ4Jz
V4+1t5yRvy8Ju4+v3HT6MfpTH1UHX4l2DZnp4At0Y4CYswpUZ5XD5y1AihdZdofh
at7xGNXZGGe5hrgMj3VaimV+P7aSgMux2RCRu4aEQjXwVSfLVlQEYFm89J3Mkdt5
giDbNVo8xudZvjVw/9dxDmf5BMPh61a5sD97MDaiFnqOsb2gD0JJVfc1sFQUfjAt
2h8ivNJMjLxsAMJOLv29WYNwpA5m74u8cTl2rjp37gOzIFnoVhYc6neZ7Ukh1MnY
iPG8RYQ52DOnh+HBEtI3chq/ec+GPsG/sFLG96syCvh61gw5CUNpx2MJLqEiN6Dc
panFKJqHg83fCwAqRO97s6V7lodw1G0GRjHFQpXCLdya9C7qLfTRSfVPXjbKGXbl
wlyit6/tzz4pZJqIzWyIX7T3bCAu376D8p3CMy6VdsVB2Vp7kIqKC0nwbYSxnFKE
OYGP2vAgYQf+AERnmocMhEftdlCjs0bQP0+n+3eE1aSnvZrEygV6DgCKPIN1bbQW
v71Q+0y8JZM9VtLybIk7Jxg1bgD76yfuywmCEiPsARnLWJL4tKnXfBKkqqhW1c7D
quECpRiGf1GBqI6p+OAVrBhJF9/VyKEKEyLTcD1hMoBEThIWfS80HWfDbLi3JfuL
hysXm3qav8eu1wPjg+mQFXCZ7qrWwlBsQjcxmY8z/CfuK7AfYiEBsIZJS1VC0VTA
ejdY6DDIoYkQhcZThdcZMVKl0OEwD9tapimp1dlEaRjL5WkmpGseuSsOjg0MoiYu
7LjD6Kt7Vhmq4ywTQwX0JYP7MxxGVgyflubSO1mG108jM22OPnbQh48hTazdMv34
Sh2pQJ3GSbkTfOyPgjPFIpZWBhRReVJmgE2kL0lIE/6m+Ck2pMKdEJ0diJvcrlwb
O6v52tWL4UjumiVpp87SxWOHQ8tel7AtqPEN3j/klyY/kyj5anlOZGV49D6dpRNV
3jQCHRzCtVD5DOZboJA9OpWNLyMnIvnqeBxextQkBS4NECY/STxpQWpOUgTCafzL
BeCtlaFVs0zfx+KcJB0HQH8wnqz3whaXaOPBNZ9RDleZZBHuwMUiWzTtd/+OXbDm
lzUPz4BJg5DbDSbTrl9rj1KLD908LEP39qNWVib+nD0ppEzxrXoIx6XnjEpz42KG
2dyr0KoEDqjYZARiCLqkm/zY5FH0KCVV+wkwE+LZQd+qPLp/IE5x+Yh/Ws/J/W+E
vXgNkErdEp0otb8fKaRoyoR+Oa4v1MJnCeQtQUO2qXFcUW6UZSugWq+I2eQlJ9iw
93SePDjCjat81pWTZI4l3Qbc+axYLMfutahctsI8ZO7n739cHQ1/X1a1DC3MrY9v
PDWnCwYrR8PwKPS62qgtkla0t0OrdYpuZneIc8UEml/MN8jUXavhAHGUwxG3Uwmu
GellVB77+eeQSZXcAgZvRDAFJd12EJu++fzpMhxh9673C5jU7tMU46i8VxJzuvtX
WBFmmUQEth5gsZU9ml7d26z3yAFwooeh9HXM/bSiqKYTFigI1Qy/iCAj/AVVIIdw
TDrVcwgKrHWMd52obvIxaiWqgtfS4NkIW5QERCfBpKhCYL8KKrTSFYHYDKWaPJhk
InBbvyu+0Ab7ZCsY5dr2OcwpAx8cLHwjIJ6LgUl15Z2fYM8cldZppetjmB6reOe2
i2UZXXypEY406LWR2uDRUJM+zchlJwEhCYcm7/1A+H/qPCgjkSn2GvxfbJy6Lnnc
EbkuHxtJV9r/oLP9+OYSkHK/ZggLmWOzxPHDU33d7reXXhb5yhOmm873AbnfvEAf
nihK9QpC7n6NrP42hdLCRUtVLeJx0C/XxoAz3FJcK4GZGeHqkMlzDJjE6pim/vaT
5mMLp4nuSzDwcQlj5TEKJfW+SvA7+Sa+G5A2y2Kw0eNhHDgCa0easDgfzuLjp6+t
x64JL/9eH1SXTAjheTty2lt4onx9EzxAm6+80Sq4RWnqzc612yX/DVogTX+0zCQt
DPX/inxgNql2JzX89TUtP+M/tQg10fAOe0cYl3wfq+dXnTq2r4nfFlQAxLOfmhVU
W6YhFdH7IGjfy91seRRW3nWk+OzjEjIkFcmgUoj8WpddBTeA5o2zFAebWGJ+jD1t
OMNAv9JGPXAWdPDTHBedjctNjKJvX2nLpjUu7i5FWeRCNVHDl7Rs0i/0A3BQsVZw
q7Bp8dQ97PaKMCQ8sJm0uKmnqtu7o4GYVatzdQEIN9/ibTQSCTWxuWVdwToWQj/Q
+O024btmY0gEQrt98o3X0V3MVHMhrofWnTCIyqDjiUb+6yl2SUmPY9ucT6FMk71W
LxhRpnf9Qx5xw+wy85+d1xQPov6mTCNeJsKtLPEnduTL3ck0/JMqZvOMSB56Rj6q
ZuiEk7AJaErKfkuhaKZYxA==
//pragma protect end_data_block
//pragma protect digest_block
6+BomaFoMMTEnMb+DK0VC4Sj7Lk=
//pragma protect end_digest_block
//pragma protect end_protected
