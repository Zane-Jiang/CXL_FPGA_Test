// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
GuuPsNQ/8Pvd7CNQvkW0VbL2aBJo37pBWkSWb3nZUdPBlLb5Vb/GkhSa/ia56Hxz
AcX/rlpnO6mH8OuLO2llBs2vAKIMf3sKL6Et+OLUneci429XyHE7SnDYchxe1SZS
O+ZVcU2koRikNIvyneIPtwNsnJrxMwrP1rMt98FaNnk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 4624 )
`pragma protect data_block
eEKvzCKN9COHFwET3fs+gMawugPvJo7PzSAmSllrjJTWm0h41Ko755AtO/rD0Miu
g4BjSvm65N88laFNBLk4lJCfCorKX7qGMnGmUE7WqcK71ChCCbigkdf6ni61OaBO
DtR2AMxjM2FMvkfdK9p2jASpPV71A2kvIQ28Hju0pHp0QriDTgHaNHrqjoX/UwDM
C7NpM3CyPKN4rRVHZTZC1X2cawOACxxBfmmXF5RMBKAW5WvlfTv5KFY8hKfCka94
Q5WI0aBGbkXYsNtI5769vyIwdABqJ+x5Xr3NOj3UMURIhCvboHcchr2YeGMtQSXh
ubcEb5CCXUsuBsQn9X28KixUkpwTV9FK51HQNo1heR2uNTBeVUsGV9Rik/3ainif
pwg8vFx3AIatibMK7ib4KobkRhXgFoG3xjA0+xS/hPhC8xNKTtvDfHGqKnCZC7aa
PFVmVjt7pXB3bvRkKs2bAac9M33TXoWUDQRvufjlMmy6x/6ZpHRmYCD9x42QzyYS
97MRZEPRiOZW6/E9qdtz2qdYmUAYgYcnKhEBBXzZMsAk9HvuNvyTLVqWTsOwb7B3
sJsUFiJaFs12VosvvjlZ5B3++RT4DmOn+LlDQ3I6qwUNglf4ASPHAu7TV1mnFRyZ
MwVu84kfJS1qNfdjR5omDmvX8pPtttt2aBPWLZsBr7LeFMZYNbI2h+LTLdOl9lmI
1M/GkIY4t5bPtXAj9b0TuEXbcVvhOfgkySSZTpipZrI8e5ccP8XVPGuXH4Z2IjIP
xlZ9IXHS75qw+kdEdki6oRzwg2PdiHIVZoFuXNXEugwC/cFIZCM6tM51pBUEimwp
t8oDOOjXCoLqDNavHQLBPFQcawfz9K4u1hV2L76mEchhHArLKWRaH3r1Om1gUMQZ
s4gJfgBsWpB9Kdrk6zkrB23bYrgS+mYglbLxax6nEk2iuVwc7wb8+ZtUi5OXxbDU
jHE44+yY2Se47Ij6QsZ212RTLoiFv3y231NfgPejVfR5x7q5EUeo2DEgV8scoKf7
LkgdU8D+Roshf6YBkN6AcY/aPZTPOByBEFER9tiG+wvMDI9bplDDXgF/HD/ey1VQ
2ybfiNKf/tJTDaeS6BGZyr7dAJB+PCCtsF/peBkfpGFVx4NDkhA/dn2BIKNdbf+k
Z4CcZ0L0RiQpmgG1M1pYQKvcP0dsl/S85GNLzRA/GBWQWn81sbJ3UVQu+9W+7wxw
48auTmuKIdHDGpbAgsR9/NIZ+DtB19cXXTGYuhT7lcKeloLBrDQ1rP2IUHfK87PE
VsYvJydJ7nbp5H42S9bpXCMYsb1axKg2YA1LK89m+kxrkhzwaWXpfXt308xT6i8o
bUbX6WYjtu/CZ20uUFbvuihtHhCZfIK1NFCZz5H7fjfV/qlOJZx1+7aMhkVax+hd
LER9+bY77AZ12r0QjOzvF66WM8bCY6ip9EJw4dmx3wmv9awSZ/xasAm66MWN/khb
SlqHhHsWqO1UV/EXwmISv2SRsNP8MTm7U/Lk3IlOHnert4XqjGw+H6NZUrGLvFfY
AGQSzBO14xuhxGtxcEmFyPmOpcAsatq5zFL8aRaraC0aK45SnOHyoRFuqKnBbKbL
np20sq7DMZ/vOIJp1wFEb2ji2lnbi+avSD7fM6mbaorFm1lPk9B65WvAdjPsjF2l
v6BsWCuUGaMbBu3niCSDdohxDQqSNGMZStwH86CLq2qR7Khx6Chx8kKHqvjnEtdX
8RYl/po5uG6sDL1CFx759QYwkFKRkX8t+NQvLEGBNHzowSZX/YGfOcevHuFe03Zp
FxmCpqIi3OQlndjznrqN+KU0fUe1wwEAl5iIrjN6coJ2HAB31I0lkIc2kBXIj3lm
JBYTX0De48OUhQ6o4ka0NZSsNRDaOWfVIyJC90Gq2yAQBhXqsfFGhEMQAAKTsKR+
EDcElX6v7BBvRKIhgKLnELKMICKUHC8C9IRWogRETpq66DxTgJl+QiYxtJnMor5s
LphGFKfI4xODjlVMmET1txZqnKVnqQYYWW5M7SQPkYl/PQVT25CepJe9WjksNYoM
WO8a6YgrsMTYZpwuk2lDLgjaVpAjzlmOQnckrMuMikkcOxVnx2tr6kRXZO5QYcSt
Z4KvQkUQYFqXRHKAfuTOGC4y+u0zsyMu+kWGMSamXFpO0cIEYp0D6xaC4Hu7cau5
1XB7Jth3djIX7/SXw6fTlH3sP8ka/ZzAbtSZR8Ip/7CeMCO1/owb9FjoX4RrcJc3
pvM2zfm4BRzpUeiYRrKmySaV3bB7LxfYxJ6JbJDji+NhYRfJqMpiqjl/VyPCW+qf
kDZkCwl3MdhJ5SbeGmR36ySuvxNtnegxq9wowZ838VyYqaWBHVIgrbN036OQDqt0
4vLaS2kCCBtBzouMx8gKIhHdc+YE5oIh08sNiH+4mbVwNnPFCBnTKi/ozubmQ2iJ
PhjxXUgvl8qNMIMoNaM9wrFeqN2e50rEn7Jkjn4dsxt6WCORD2u09pPjmdQQmXC9
P7PidGCRl6OwnXBESdVkW5vqJAOrWLIHqniJgSxqaRfLhu2aJ/pe+YcoXIDDl/HJ
vs/vLKhmdyyMVDzvq7pl/An2UkhmxIHgol9VVJlMwT4E4T38KyVTUmjtLbjJtscu
E3yFezK53RDc6IpDjZ5Ag7pIhRBOiCh4lUKbRvdKCbhm2ZdEl6F/Htw0oNhNaw4A
SP/1BzWJWegUwo7skfU1F1/5L0RHZC7Ep9TgHXPkSwniPujSkAGIdYfSzmB7H/zn
JfMnCBqv1yqxYXL7xtvenUgjZMvlVfzE3CEdFxlD6M7y2mXMTIduvHXdFGGLRuGx
TKUI6h3Elh4mLXW4vfhA+/2I6a37/2Bhdj393H19O3WwvwVL8cuK00MYPBWqdp6s
Za1tRxOKPuUxdy+/71pQVEYQwLUOf4BtFNod7MJc3swBlbIMqkbrAyZBDrU1bJQN
rscc0wAGnoMSTDF9nMw89BYOP3lFMZAj+FH2+XqcLqWZVNMF59Dp98YrwFcY8qKS
H5wrXRJX+iLme4H5dUOU/GxKvSgco9iV3zPu37CZeMK2+YXRSJ0a7IdVXRtNMiwi
wUJBsaGBkf9k8Qf8LhQ1Aoq4OlgqVDszn1pBRIM5f0SiYSR53YK1Y9RhybcgSbTY
Byl1YpxnOxCRBmqUBEYFtNG/+gBqlWnv+PEVAtSqamYVB1OvXt3kFXIS5y/isSy+
uaiP/eoUh4O969bVLLeky3U5Iw+oEjlwIco3RaoGavfX9qH/UXwdRNl2DRx72h9k
0nN6Gkn6cQfm9CgF2nJWWStsyVrkqMwZb+a36gc63ZowMB4dZb7OrKUOy9NV1T6g
LgLvITembXhVevbixYIbXlFswE5kT6lVTZw4TEzMVsNxlh6VXn6ybac+tQm6k2ao
a0Y1mYcTBu7okHLA4fjrt/fsXYKdKqC2VQNWkHFUm2t/OS1LySsYYlWasFHPqsvw
+NoOs+7Y0bbnNYr9QRGHAr7O7Ei1x2h/+N4ciykBuf3cihUeCBZY15sILObR3mf0
HBco4di4drbMar/ZiWooruQfIr+NY1IBeEepAMAPygA0XTMoIi/5XoDtmu+Y4JRy
k2l40Q12Iz0839JBk/jNHgChssZ/t1UEW4VwCX4X5uck4r4UmOwsOsFH/4Vs6LQB
FNXOrNzGtSplQc89FqTDUI7iH4qjxYxc4UvEGhiqhu1wmig4h0Qgb33u8K/ViO0A
Yw151JZe4KA74zvIOh1PBwOvs5i+QxjGvzbc2i18V+VC4NK6kRAgpL8xr/kF8eE8
TMfekEL6N6H+O3JVPakIMqur16tRmckW/+tApF1LjiwVBP5f8li/+yBWecheO2XD
2bZSraFQD+WBMc9GeEn/Hm8v/vMBmTttAufN4GPoimoMxp/Ij+W6ml8j1Z+KVZPf
+QR+AaGRhIeG5KR3m/RhXRh6vKjCGfNuq+PRhMQHPqags3iIpWfLzaZRFa4Q2pTk
0e2FoIPvWc0p07TdDIFYKWRin0P5QlDWMpYxbbUwXCqEcwK8MkseK+DSOxLb5j1H
kUhM+9eUD9teTXGUfhOoBj5vzH+iiWGzj1etHFBRzBPgJAzUkByFj5UftcaWPMsb
s5i0Lp75dpCQKC8Q/amTorL7jM5YKweO/Wv6lF1Zzkaj0b3ZHieNj5QzxeRFRosj
TbX9UuGjpNWPdB3j/lrrp5tswuQ1FkFhfSyS0v0Jh6gbuoz3IH+hsbkWzHVTkh0d
nji1M++151YFyAl+5hx8BdY74LaTfKWOPftI0vWF2Gs4PBYnuPGmR0ZO/S51QWcD
Sfm+2NImZ/ekntQyoAWTToLL6eiLHNue6VDeTgw9ADMjpbALWM0/RXsOo/87mujO
djBfxiLuVETPC3PpSHXYLZe+GQCnYsKKqE7QHXrxHUPkCX1uYutta7gKwopnLFnp
IN0yIMxrQjYybBQmkSS69w9QlKaCBwTWqIy1SA4p38nkD90TcyZWveDzeloBp1FB
nnylyQdbFciIdFVFBp1SIt/C4ZVay1dNPyQWuHzjJM+Q2GI1GmN5Y7RKUAzKq8Xc
glYw/9S75Yadxk2wbDPZLwjJd5n+4rrt/KkAGYTvakqdhDbNPA40da83ceDgFpQc
U8Ai4IjeVr3LK8Roiqat7Retfo8qOf40RFblBFv1FMSb4Dto+65I17Rz05LAH7Nx
WnL4wSBi11/BMNeG+DyF3vsgoyShGMOb7rrhWLFQtL3Sb1Ao1PidWQk5XdstKVZj
9dqVmOqOGzMraRMphfm9V3NV6e2CgHqmugA/iyZVoG9MhKRyKsbcg5jMFMGO7WFp
AF4Hkynue4q27lH2gEPnPVBZskbeeN1Qxj4YrzbQceTeg02PULFqaa7FKgcradjX
hXWKH26cv52qpXTXkIfkg9SsAG92wiWWQrVyDUx5/aUiOEkLHlCFEWbmNuhVq5QG
kTjtR7C3PACzefTLi4CXHxPqO2HxxqCghSfSIDOJfOEEhtsCVDGqQDnTWPIamqAp
FxPD2pqLFWcuXYQU4DmpDOfRe+uokhIhZIrB+g7nQ8bqaiKdcqUQGdkqXkLOCtKW
S0z5QBwDJhZ1NxQr7z8+zrNPFA4dldv/OCBsh3EEYBDV0nn2jWo2EgWVAT/3fu9L
Y7+HgZ0xXXgxZe+BNQqBhVeEwZ9fI2uXnupsbVE+dOOyIUCb481ngd1hjjTStgDm
6xDNXQE7G13rpiFWHUtkwFoJJZbLUkbj/FPkbyYORK3dNr5QpC6rfvPIZK2ZILYk
xUG78MSu8ExgNpVO3TRP8m4IVt2TGom9UzwFgGcUP7R7JaBgG+0PLvbzDBpMQX6g
AdODv0rdEqmgpPSujIuqbgmZ3lKpXIZZr4ccT9BshLyj/Pmwupf68aFhRFJfSUUl
I4SzjTQMPEKai3RBfGgJR2NSfzn0v7SyEThy1GU6Oc8NH5QHefC9N7ERBWy0El2Z
zM6U2IjKM5DngqDP8JfMDXYUsuB/zvFBLND700wC9s+QbpJJySEFoak/2jQa1rKN
p+hWsOsL45hN2KaDsAhIPiaz/EjXYXr0nVmFJb3YpqqhUgJiFu14/qHIkkiGLKjB
3UO4Fb8bSMJaYrMW0I8BjY87sV8ZMLJW2GaQCJlfg8Io8+5/hz1kDROmVR8l7xNh
nO1NqW3ifx4vGDZx80UDeD0+fuXFrQlCYFHVhSM4C0Exjat3BHQKpq6VEFPNOTE2
H03rQorEzhzKxmIo944z7tHbVFlXeYifQyOsbq7IDL7swvTRDIS48seh6RfvqlYG
dJUTbw93len3Xz8+j+i58f0Bqt37TiHqwHvdf481bi042BuRKOt3qHZVuRL1Xepe
z7X+PPMNV9wF2KbGPQHKgZNYZ7bF8zWOZCprVFdXnFRllkjHZe2XNDwaS5OvKHSB
EKRSCcUwGCTZjmUP0anN8AvKLWNSvqxA4o0NRXKo5erVr1oZdxzlDCtGaVQJ7iX2
GWa7LXowwa7ewwvCbQ6HQqvqwA7ZiGUR5Emu4CB27FSGwYY0wmfxbigNu9UOlsVG
NpAeVnhGwFj4U3WBS564VGCFSTC8kgKSTKtYAYOGkjTYwRwZRfqfC9hIvP9pnxiO
J8y1jyvWQm2ZVk3AMLaoMdsW8QH/EJn4WgJsSKNSirQmt8RSYEdZwTdEcYPtncf+
EnsYFVhpokxbej6gYoKG7Q==

`pragma protect end_protected
