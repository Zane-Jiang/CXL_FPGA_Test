// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OaC6onkeiRZXXyEO7GwlfPNpW4CkxSh0hxhtVWixcF39wUnNHufYeOIx+Cic
5Hko3azYOEej9e+PKFOpKeCIhoWcwdi7+mIJvb1JGJkISgOwl9tBnDSn1L2O
6LOpfIrkJXb6Q480snCYGmTIXPsqLu3ZZYe5PLMaDHMnk7nyLnDc4wCxJ9hb
itzQRdUQLmEAre8nW+OW2ZFunIRdjYW1DNi0+e7gV68hnotL/JlKKRdQBgQU
y4ne5cB2ziJK/1LApJOUc1BFatdKl12ckcm2AobPeX2JblQmkChSXBsqRnAq
JK6u8G6GEZHHDh2kbGhPPw7pYI3W6kiQUaLLzpGnQA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
plFBl3FQhUZMhr5ry6RM7JlI5lovqGnwrQdaQLCo5w96xtrVcV9+TLBBsD0g
QvmbaFMjanGRtKJ5g1mHSSbzMkOQaPTI3ddvJov3ByzU0BhNiy6ai9KWz0Ue
QP8LV8JCEPhPwEcY7Pki2Xr7dkRUhbZoeHqxkvtYjuJcT7eVjREGjSDErjAE
HyPChqpQvkunM09PiZiOO+E1b/JmkB0rbazmVnmPgMTxuM8hOu407upoNZny
IV673G8bxxhawR7BN2klPs7M/EkoQiHGIcE99BNwI8voDODF2iBJSs0cGAKW
gUtUBRjEnmuP/9hm77xsIjYuPNQTWTD+BQvfkjF4zg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oriyoepzm5Zcqs9JefzKfaTYXrs1aBDZYuiDEoObLJU5H4gF+biT8CdbnLRw
gymGfCa5r8qNlxHG4atthU+XjD+FhYb+dZ6sviKzy9hyBPoOrjoL8yBfEGs8
XACCRL2sDr/0E02Ns2JPtl3lqgEZdSk5sdZ5PPbptMJHg8uYbGf9dCgYmXae
7UxLsd/H8a6F+uHDmvO4x3YA0Fxd4gVzfA9BLSiZSBK8NL/T6IEO9GbieXhk
nQDugqhPN7nyKGnVj0cZtKgC/3U82zlp30bdEswC7waaPBOQxKK+o0IkONcD
6SWU379qBIUkKcb+Ayu0yUqj3Un5lDU9GBrBn+upUg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gUFCLN+kSRKHmq0VNFIwo8DzAFVIEVLKMvEDPGzrMUhat2/5aAGm9TzYpOd3
E2QeaQHMlH2EACtLSLzpAlvGsKw4PxQTCB8gRhuVm6quKPYsDDk/7KnX67yi
8skl1Irv61UW6piTz7jeUcUswW9+elEAbMcNH7cla6CLwzguL6U=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
N5it5Km3kAzIxA+i5sjHCHNMQCDbcckqiwvrJogkt2UC7Ho7rtSI7/QmXfWV
UM7oam3Takq6QE/SUB3tcWYPV76LQLHp9pNtvP9dsFhUelIQMSPrsyhg+frV
8flAcbirlcktm26UxqOSymzWYEKKXAuaUrdKrRM86Z4lqvQ1ZYnaGsze+hAs
re9DDkLmnTq6ZxCzdz9BlXGMcCse+kk3ZDamRDIs1y/oakQwIxQvWWzt4Cig
X5OVuii5ertEJuFYMHwS9M+FVDtvq2VT+P2ZaJ3vpUZNQdrcbCHk7k8oJQuj
fACWeeaG97YVxyrJcQZJsW4cryzUEEnf/ox7qpoeQriCH0YpXAJJb7bUwnsV
ckQZPsCAULRDbf+2QCVBCKGWesrUhNYL9frRfWoO3nyh+5FDwdjkI9s8H8H7
pvpfn0aUWFVEMnLwiUd57nMeFI9Q8VZnGT/GjsncbT7/xVeMTvWG9LvGyi3T
9XGCfYVxFUHWNImFNVN9QB8tJjDU8vDR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pQufPilcvgUDOxe4AQ9/a+ngLVWA2VlzwksEKmrK5JHzLSkygMMx5g4nMx25
OZXb+Kg87WXWAMpVQmT6CHmKwAivikYJEloCKJD7w5YS1j3xky/oZ+diSZ7q
Z56qsV06tqxRXSc/x0oEJgciPNpv/UtOICKTevyKShnkDOBfKws=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YQ9bAQXnnyq5UIHmGC14o0CE0L8deVua0IuNbu0GyA+om4gYveKGrS5VCmZx
uy4jIFTLgrtsbHZY58TNWBmChBd0nQldEUqzkvI4suGyJ+1dmcaIxhV3Vtev
h60HQmv0CygsjayEly+yKcJVfXOv4bTsZ6nrhCNJoQc5cGkqQoo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1104)
`pragma protect data_block
Tko6IrGQLnRx8mZm9VtTRt6Ibh0jZxlxICrPo7unwG9F6a+ReJD+A1UftB7M
mWOnIL9u19tokJ7m1UtGQcjFxF8bazWeHkbqs91C5Ogl9Mh7wMh8mQ82wVLp
yw2WmEky8n1cWKl8TMTmRb+6Vu1y20+XYmqYUhmlUXT1raKuZl3xvYWpJ6S5
0SjdcOWrOxfuD95LyAU3BmsDmjBAPFtHSzxMWcmgbr0M0vQAVkTyvwjerskW
v12vl8Q+OTnd7m0mDAJKT+sof8oqDDIVxGYEZAiZD3FaERZIbyF5H96RcpB2
ibqnsl6XQ8uEo2l7GXDkwPMiX3mbc+L/UQXA1fz0Kq3KyAL9MIjO/Xhe8pY3
q7VJvbjM/66bEYlW10YbZ3qtwxl9AFtO8ZGcGrEAUtEz5uxa0Sj2K4iyJamG
NAmKevg7BRoJ0uNcDhjGMsfA97kOChRZvMgxLtlnDly7nOlau018zvfRaAx1
uD3fOxtKEYY/jmiyWP6dTYAf4vF1njm7DCwC9GLOm6wB5JBroWcA87+IoWau
836DEGRmyS3USBIPQmDqjvdvPBcrn9UfeyL41lTzVN8+nq4f+4iiP5qsLF7W
Sn+xv9XU2XXTEshXRldSjA0POMIXFQckjfcGZXS+IAhHV7LEtWIuFNxyRJS8
Uson3mb64Fk9Cji7ShRg7S6wH5XEWrCNRq+/AkJvwqLadNiuCyQHnGFf1wLw
YtJTRCm4bQnLGF0Gc4bTmBOIAjq/T0M311GZQeNKfOzzKAA/90DLDuF/jtdb
6Uy2EbGpeY7O02fjEKp8Gepgfv8yjjriBBoWiTsZGC+68MgjLGX871vElTKt
0anppKcWwcnr3Izz7o/ej3XqwVbzR9W1PAWGlTYssUdP6EwSMLgVO1Mr6WCi
mZje7Vq5xYU/yZ6eX/w0mpNOds/Pk8d/t+AD2+MKbE1bFv8+PshuEV4P0tiD
rL1DvJm+/HQ7ZAgOAA0k29/zRFITW0xkN1Gr3gnKB5ydcRo3LNcXR6C40hRk
KuV2MoiYJ7i2t4Mpwmv8ThSYKhd7Dei5WKopNXIMouj1HBdbuSnRTgCoJyMF
I475ZNCHrhSpDuRpvPoACOc6m/9ievRUbFjOKcdB4xQ2OdQ1JFFDarIr+S2z
SUWhtV3dkjAbTUMK837H8JIwpstoI9aljbI9HdITQL8wcc003FUZpPT1X9vO
xBY1eVnb+W7M+TXSII9cDk9+XNwzaylWFvlc3uqQqLVc5wtpFvhZ7ehyfp/M
xgeXFK/ukjFwTGgjEdSoDC78ohqWhaWqd3D2tovKqSa16rkYeoEf5RjJczP5
QE8aQM6ZO+binxWCcPaQOz+B8lIq8s7zuKetcHFtskviDvDUWi+boRj8ljS8
6lep0fS3QxXXwjOPxWjZBSIEm9Y0CtmkBiWZCLvcZtcHbzy2txkTN/ESZmon
yVo3Rp5quQSiU7NCMGY79t1Lb4tPhxaE

`pragma protect end_protected
