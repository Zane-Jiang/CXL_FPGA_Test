// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
loi7lWEyFunIIgTOFu/zYkFcbXJpoF6/c90I0Iv967bhosSCZPmGo6RCUAj3
xkoV10hSzRfEhUum2JB3RMmGA+rgeRUHWGkWaS9HJe4/yoAUKsvA48SwTAHb
fo5RypTZOcJ659MUl9Y97aodv1vy7uwuFp+XWjJgvYg9zoIKab0ekNBbqBmD
ZJezbdCoyl9yh8pO0WnxG/uinq3DSaOWPNyVWNlPEk66QgajPOZ3iH6nv3Xf
akDI40gJ0jaUFX9JN1Y2pvovNENkqvRvQMSVgXgL1U/f6SiPFFAR4PxyWNOv
v8Buy3RYjh1zX1uu+KhaG/g0qqBUt1guk90R6SYIIg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JYpEqzBBb29nTHpBnsW48X3smUwFvdFdjAn1tqfnMwkfob3JxrEmMWcRXWdK
PXHW5i643LObiWt1u8TgM0Kq3ImzbcO5fdExk6R/35b4LdqxoGXsOviqZUNE
nWB7z5Hd1D2OULMSV1I9SOAZnKWf4REDh4plbx1xs5CL3Z+r1HNe/zE+B4r/
hl71mf+nzrGBSv/S2BoHfGeBnSvDCbQdjcOFtC4WFmiMmAt2ulDBIGHi4Whr
xvDwImDmyeVuNeTGovujmFLfS+VqEB+SVubdpNSobcJOaGo/XtAj6E/TW36H
9G3m5ThVs0fxSQ6YgAlflJFM45L5EhaGHsbytyTNng==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MRfWl+yKSqdVU2prZ12wZ08eBh5y25sSI2JGD3AFTC7ZZUxg320RADb/4XP0
cr6SIZ/T+0YaXxDn+84sRxIHaINMIs3JnUGpL67EEYip5WwJRt17F1D6Hunh
ipRT1xEVb7WRy7aXQ2lpxLd6Q/5fh6Cwt7lZLHw2LU1RplHzcYXBuObiC9le
ji4wxrLwherZ7xLEhkd6KvEIqmp2ezj+Ji7aM0qOzTFC3UkYL8SWVoBckDKf
liOLOkt3I7+Po8dJfbruYQIy3E1J+YGUOzZWYXqxwymDKdEBbkSrQOxPwZMD
B5Uv7ZzdP1Q8akvAwnkI63i5BeQCJjwfXhmKs+SLUA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TbR+HJAAIB1S4BH+8QWF0jcnEjePKjTOA5d7j+gQkssXVW+aX9TC+566kNgB
81KSADlzV7BNcUQDVDQwVH5TEelU83em+xeqsTj6oUnAl6kMtwDFl/bAB15C
GjiUb5+188/GfMAVaLHG349UpYXrD0Hd7LVD9ATaV88YOGs9uiA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jYBTeaIzq7bJ2UadavRtnUWU0xZqSMoNTrg/DkuNKkKBm9BofzyTg4zffsyv
KnwNQz0zCq19ijRBcoAKK7oRtBgCtc8BZLyJ9wTF5fhZUvMnS51pZhsUCN4o
pInIFmzpmbM+sNebCx0BC5Jp/g95M5O5+Zd02xRlvH7ut/UVOjF+ZsnrfrF4
icZRTTjwnaGMqJmiBcDrm22E33Bu7r/xkuOBnm6O3eihCDlv6qrqdPaw6yf2
PwbNw20hrS4sYrHjB92d7iUOLljr2rj8RDTKOUHTXqT6O7sulYxJN5pQI2rp
G20ILvX4JU8Sr3JbfzttKalMoLtRI7Rs2cNXvC96vdET0il1jHjvitqgzuHa
5VpFq0GR45yeLlSwB7QGgfmpTpeOIhB4DIjrCxFwTRtxRGYhgmHKfzJfxhq8
C7K05D9R9CVm5EjHKMvb5q7hnvOOI0jzxlCbx0W75hNa1H4n93DnQ4aUVeU1
KP+ytSdP+bzEzjgCeGoKnFWdBz0fDzDs


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GloqtSfaYCP9mlgEM9yF7X2yfDpMaFsJOH0Y5pG3VI3cqbjJ15kyVCOMyleR
6QJ4H3N8ecsYs6EoPwqko5NPly6OIFJ5zJ+RlaXX+3x6+aJjyDIM+QxWo/TD
3hpexThTuh2cNV2hxGxP5VweYhkBTnvRuC68w93D17HckfMpTDc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZpNp0xuAIsBDikaconIYMFoirxosRHBGnD5uchewgXyCYRx12jb1cBRNxsdW
G8wCRkjvmhJ4euOII5ypsIwwJpMEAM1Kmh3vsJPmrr22o8T9uylc148fabLD
Zv2xz5hMdMWpyqWyyVtnh/V37Tw+nTwYyAf6OS6wUH5h8znF0OY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1104)
`pragma protect data_block
dqn147Dsv5jKZYu8SiK82XU5QbUlCgOjtQMyEF5CtCI4ZW8bS0YiJV9zQ5X0
ZCUg76igGxeZnKyvfFkZU9fidynF+CiInftAjjlqUON1bmp3Ucj+VPMQR2kn
xFgf4Z/wE9ZCdl8XzSxLSRkhG4UH1+DkZCdDl2O8CdQcX5CIeu3GMmCvRhAn
Kix/gL8gDYH16h6fz3jyxYnPz5/5IKfV4YfOskVh/1z56LM6lZMuuoKdISvw
BI8zACFnq1us4SAJHRcR58Pqc7SepoXpXX72EYc029smKz9Ud/db07OS//nU
JBcNT+sgwlk1nUTXpG/ncL6Ml1Fr7CRONAP6kfpyBBWqnsi4gBsTlfz9ruq6
YW3z7QaIEOGh4SE4GP4sIG7PtLXr77a3RNhWHZol0dvHz1z+wDPFCdGZX7sL
yUC0iHxBJDOXpxSpkfGRipBCazwK61xdALL2SRteLBonWGkPFeDjun6wETVw
l/D2fdBO+axioN1Yrk5qGZpFgDV2HnfZSswuWC5WMoGWtlqKcrhc1VvOXRTz
J7tfuqhR5te4adDYGwAELlHQyvDKstfj5P/wSxtYB/pzZ0XKaFxNkFTe7oDJ
cvR1yMtcqUYKUPi/nPnQ8id78pK5W3p3Z2RC1jlH6AlunyFnFDWdv7UO/bZF
avqcREn+ECSjzTqJ2gX9bILa4iKnrzqc3o/3wjsOjVTNWO79ozjFZjAmCikk
1bZfVi1UFypA6na0y6Yc6gEbUipFaUIYt5u7YgLFXx0gHVTgT5lzRZCzNUV1
hSJZfsfUh56fr2eWRDJ7ckriMa4owYhawDmcZd5FWZhkge9G+SUDKrviDUZm
+Jc2zmkfjqXe0DetVJ33jZbg+6kRHg0qmlvD7oQkkqF7Whj7C0wNdjh3+Bod
wc4KN3+cr34iBq8FKKRgRAVmrNhwmeTU0SdgI8mDesroTn2DDe/E27NT7/0U
H3KOeemQmFFxFCBEFMWNREFr6mbX/ufVOPOYWxo6BF0dl454EeiAbX0dg0cA
Cvw3JJ4lRG7K2qpYokW7nXIb/jIrYsEbklti9vZBQAwm9YApsywzOV4Jg9K/
L97pAFzhvNMv+3OPukQwpgY4fIu7YS9iRiqID4EFovDMhzs+B2fRascuUVfc
q148e99Y8bsTkILTNfwClELQzStCzbmCuZhxatrgpzq7fCbDE6eAAoJ6QrWu
ncmopGy+8pIUlryUn8WDk1B8VaxdHbUKhOPr+DS/q6QJ8I/iAp+ZQRTnWPtS
0Q5Pfi3rHY4JCCee2U4Asopxi5qcYKiR5ywjdfeCKm5OWLmz3yKsbm/qVh6D
ZHw4OPk3KS4uXD4hQaf9L3RibuTjOBHYhAbzjqTEc2ld5gEZkHm6Zx6p9yKz
g9c9oeROg1gg2GDsuic2cqfNXWKvmtAiU3iorLD6WWFnHHWMAXXiQA6mhaoy
9CLujDz50+LxWR1DPM9HpG3i30JI5JCk

`pragma protect end_protected
