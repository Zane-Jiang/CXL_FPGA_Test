// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
chQxZjQRLz5fjor1GAIlxwFJ1EnvbbhfUuR90FEQc9nZ+HtC6XSLGfqkYr89V1wo
NU/17WrFV7t+n5CFWpJmMKU5/H10yK3Myw8nOlnv6Mbv/gGLx2wtYk1JK+r4kWJf
C/xQHebb2qlPlp5qmZKhCrkL5Csu6Fm+gvEL8jZwn5g=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 37104 )
`pragma protect data_block
Sdh+9AwYYCj5Q5wuxW/PysW+MNur0C8x4SthDa3z17I2BQ1C8wWO2tioUHB25Qdp
NNPQv0JtmjktQ+h7vACiA03Hr6boKlKpmW//Ui3ojeQ9HCCGIm2OGlB7XDMpQPF6
pLiWLUAytk9PPMVWjoYwygOwxZswJXb81W/TPPc2VK8Q/hGw6Ivek+6y0283RE6z
iWLEy1WNgg6VGcpMYSCW4WSnxMejyEXrnpzCZ4pcv7KQEjbeDnEFUIMP8P4YcLTP
wZAZbXsl0z7fWBxLZ7zrTua2zZdHDuKjEUJj5EConpK8GuUqP1dDINEQ1ZH88E/W
lDPCrgjuWI6H8+4rOkivF9Hfaj0k0jH/rOZ6bn8pIqIjjGiSBlcN0HG4k/bzJFar
Gcjkg3/RxHZN1KFeUoFHlQY/R35KBPrvfWLJzZnmg2mDTcJTz0a0RMgbRZrdc+Fw
RMwQddo9RrxUmiakTpAmo1s1w150bg6fY7nRrQt2FmXCDGJEordXxZSWXUXnVu/q
snuyLx44wcNey1O0VNqVJCOKSO952Qitlw+FhA0GFb+hIUCPBcx1ieSj2frSBUlH
EG5NfJoqrDVfEbG+ciJwM9eNUhkxdonKMvls4TbN5ie/k1zEL+H7Aez3BwI7Y0yU
+FZJvqLBswLNayQ90fPnfyl7lhW3KrTmfiJDElZT1lbh7iktb/IkyE5lmMKWfCxt
yDyXsBdCmI9I0S0zN0bR1OBbneSgPASyWZ48ssezm64Ivvlc9yFsl80VjrNBtsn0
Jg0ZvtGkH0aEAAQTyPOjo1Blc8YCrnR8/FgowXH49rh8TCDv2yM3VUZFesxnnH8J
bYh/SvofbQHKpxYhfOQ00i5JKzrya1pyc0+pZcBhnFMLSlnBGjdN5iypxTfgWGaC
LnqOVyTtfFNM0J+ucNdmW2AdnkFNoKWUxHpoQqKJnuQRNP3M85zu347VSh7aFZ5I
3hcAlfprOgoXFyDto7iXMQsYfFLfaqOpIHpYoN5Ks2msJMcNGjH7P72B7LNkEik7
5opKA+4jfFesPVRtzFTxr03ArUg5+/r3h1WTVhphRGxBo44zGEeveIM0P/n6OI6x
SXH4tMgnoSBMU/VmFnokyrhUXlP7521BuPea6MzKLPXpszh2KEUxEhoI64YgCV9N
LJlTwmeqAhu0catkEMem01esjsrGh3AX7eOJft0bEldnMM4/qNxh67dU2C78xqEX
tp0miNo4ZUz7uRNl892iq9ApTU8hfQbJsf3QWiH0XRRb+zkTnEiR5yJVIV9fh5EJ
syqYzWVsm0jMkkMro8BKoRMTfGDgj+AY7r5lGlIaLKmuYxhyl6u1oDHeAjYt6nQ+
NfFcivh5e+WwsFnoQCCCG/bBMLmon/bRVM9hAcQUpCqtD9oGel6XSx09ZrgWPjlr
f8MUWef/zWmPBZAG2dckavFnzYZ1X4ImUXYKCjw9APF77fiVM2cXewkNeIJK+jl8
yuRdbOUMlgXWFSh1MSj66asviHB6To0m0Q4hHCaho17Uck7iRKTFkeZzNU4+0OCP
fHletYeVzIBxpYYB1Ob2gUl5STduli8R573mx8yLZZE56jVKmv4M4Yr0re3Z5eFz
CMN2mV0XJUUh+YIwccd55vDt5cJsYKL2xtrr09kWh4drPMlZ0SAhbu3ekuw9OWFD
cyiRcA1cWXzjYfX0p4YwrGLGkZAyoeYfX2ExVnwAmT5fMLGFhph7ztlIxgiCbdLG
SMKDDR+AhRTMKR8ctv8stn8ObMDsTo2rKx/QwAXG07Gp1TlVaK5754k76YnAJVRW
4Tn4nIcQi5+LdM472zBuiZj+dBtPPl9jolKxap6SeF3C7TW/75YbKrg9lFN8faa3
jTRHK1HhEqgd3l8h+3gqSh7/qtBiSCm6l9x9OCpEboQ5cT/0BK9WLzSUIrmPgX9v
VRVBU9f1RS0vOgX3Spzo9Nabt55gFTBCyn5Y2z+tq35mqW3hFVTfkk6D/7XMjFEF
iDBd3j8G8g/p1VTbG7g0QwZlXYHeDL6F/vT6guEjmMo+CvDfiNLZoDSMavqkzSC9
69s3FxIjyc7jfkxYumghZIMyKR9RqPxFQNowisrV76HPjgZRiwv3UDLaZjeqxkvq
Weee9kJ4/n58sMdpVJDv+OpJciFadjE9q39vW6i8tOiRC9JFMge794SC38AzE+6j
Hzg4g7Jd3ajZzfDNbc1gvqRRtNEsXGngF3mCWRH+D3Ejt155kOoLCJic4OzdkivH
WiAzup/05Dmfm3zFmi9lVBqfQYGV3C9A563M1TqlToV2P6kXXrQB+wYtTeAVdJAm
4SyXBDep5zqrRPY8dyUnerLxBntgjttA7F0nURektPZpon9M/41QSVNPXKYIq5kA
BKZRyXVEaakqgqORtkmr00NojKHz6wh8S+BrDiBNju0N924ZMx4XgGJdYCGS7xaQ
mYwv90CHBIFD18BA/yQYC6S31MRqRdNiC7I8LQG7c2lvo+BHBzVqHAyfb4v3rp5j
gL3a142kI9l3QjXIugwlVa7TLF7aZRwBlVs0+GjqPQkomYlRUo9MWngX+YlHbN5Q
4JSWJDDKwWVxdDJr7Vuf+YiaOqaZFDSp+vWZSTUcTZSR21Ndifcj785uVQurR+8J
sNsbbw4laC1mlBB3aoXLytleiN7Jz0HpApZR5SLcYHGGgGixYJUiwsxJrXz1VvEu
q62FdfT4HlWcAJ9UcrBpHxT7mmj8cyChgvOLw83eTQdDl2nmRLGWvwaXHNd0QfsN
7WrDQLc0Rush5T1Cbaqo2T30cUjTERmwVOeIaw0CpZapfoSg59MrjQZRuvdDE7G3
H4MO8JLOmE5u78hAex+g60CF6jvYQCJF+qqliMg0/Qz5VzHWM/d2rhxNoQGfNDr9
15DEJAk1c55uE3G2znee7wmV3O7nfqHOnMt4EOzSNodmtfGZZJAt8ezDA1pXiP/r
LSl3sxDRIWW8nWY0nJIrcnUSLWGEJqpaSFjeI3iVqDyNLpVq2AvM4JDkufu25ybw
fFWeTJYMEBRbM+mOyGi4SG/TGVo3GN/mkECRZQm7ZyRATYexImtQKVjV0VtPYEGo
kvMn6/EW/1SQ681hfYLMNDVNbPkqRvB+ttklfK7CbKZOrxRep/mCwtDs/IZA6GPw
rMxZU8EKpcqJGwupk1D8yrEfrTgoisj1m42zLAR7W3Q+0BOqNN5666kEkymrFwXx
qUcDRhGcoKVA1PfedZypNIX45j/ZH/Wd/kkTpPza9/2bscD+D9prUs1/vTJ71/QF
3tZfbZyFwnMTulUetlG1aochcsraRKdB3ENT5t/v7c9Bir/AvInNlhoeruO+0I/p
8YVO12hqRoW+MD5aY2S8lMC8kmauzSliiPM7pg9qJkcdA/+YiH1O2xgpQJM+JBfE
fQ10tbx8KRzZjuZTC8i4pS6ZIXVgPaGyDlULLYDCtZ59EuB7QucF3KGeYRN0+eGL
8xnUzpu7Brv5jLxJSZVigNc5qDIdzq05Pl/AdqJr4574IpSo74qT9CnjjVOpqG6A
LG7GLHkc2B9GQqEhRB4HQp+pUm5yvl7ociwiUy1eisI3w6JgcCmf4iLXT/zGpCGu
qjkzl9Q4t2AK/yUx/ftTX0Ij5Yob4Dz5fBgEzDN8jqNOH7IYryd0VCqbl3mP+25n
WCe+xrkokh+dbOYhQX7WYdxc4g62YwR9bukc6C6cQCf/YdkxlgVMZ0c3Bf3i2/xH
iupkk6hne27e4IrktUjR4tRz1SKeCTA4Wf4xLoevePIxQVc7k8KP1puaY2fFjX2d
Qxot8PTo/9c+0TF47kVR+TmIhncjhSIiSKWkpxPqiL/NGlZgwqFdsQZsm+vhkrpD
CNBZhzamof+5okmOW6KdWl6lm6WraruDZPwZlaoXqoaWTRf9ayR9Wqm8c2Rl9LXw
3nZYXViryUB4TB4pvopc73GNlMgIUe6hnunBPRUqHwevc1wwt9ubJfnKHSroQWS6
Dyxja6zqyv6rV/bSU19Xlh66xjx5z1XVuihFOOKrrjlYfiP4MwJzhc7f26a2fT8k
yKAYKAPrRct1ZL90Mdt1oh8wlJ6/ThOJ1M2qHpXoQVt8WwCZ9UCUCiwj2oCuOeyZ
WGfw2LyB4Hs9UXDF3H5AfZDf/GJgRsJBpAWnYJOTObeIVsQiAP12SO+vljgeSrai
orD/06OgZfr/dNLSPLHPH1uC64qM+z57mzHlIekeu4v+BsjnlwJBNJZeVUZCpLv+
MwNfpTznssj9gOJ//55uQKW/EgGv/EK9stWFUE9pTAokp39mRY47Rcbbwk2lOMZJ
9ASL+t/GNkLFas/M/5puyOha+jDQMAvPwN3wM1qnJZZb7VMtvCcO/uCQYMtSrDW2
dYTl7sFCY9MHt/8XxKkvOBDvmQjbWJ4nSqNdAyJ2P4wEtJiAhNR8lDhO+Il8UmIx
RzhcWJbtsV3HDPduFuHpNgjq6sdk2xVHwZ/H8o5Amx3mhl9dMGw1x7Fo6HxRanfd
lGrYikK/rDSMaWjs4VSrdtmqYw81aY08+x4oJB2yaqqQckHiBjHeZWoPc3sjxZIB
PkUYfMJi3DoMcoCK7YnAKr9yYrE3Mja9OJOtpIKqUsKddKajEjPsHtBPuQD7aw/b
v6dgxMwv6u9X2ZpUnuKuCjWgR53c6T7V6BvO4PcczpzZvq28QpDil4raURfJ6tkN
6QuW2wv36XMawwqay/FDQk1AUH7xcKoeYI60RtQ4bDe6K/JyrZcn833FaK/w4zq4
7ofpNeVhoPycs0lKpf9ugstE5UNXlzbWdZOR0DeVjO7PBlRec4TL2ZM5g/SOtbKR
1Bje7ePTmrms80cyehNvcYg40tl0VfTCqsmtHZs236VRhNG61mzRlRDfaUKKzp2c
DKnaYlAqvK+hMr9levy2mXthSc9IU8V8s8hmYYzyW6ZDtnvaEtKDEqn4xiOuXGcS
8bBgdLPcF65TbXNdx/QDkXHnEhkPIioloBuhElh36sal6pMJlKRoqfBP/BTVwjIk
3vJpftysonzehivRQ1JW2/hrcqdqrbwwG5ArhCXFTTWGzLAzZT2SMgqXi6dBQxtD
1T3vxA61zXRdR9g3VW/Coc+wnLB18VYinMY3s9eyGh6s6LMM8XkhpaPzoMNr6Iuq
5EwjyjWDLPX/EMvI9nV8baJZnH90GWit17P2pxkx/7VGOFo9mAD4pqlwkx+eMh5v
z9dyQvD8cyJNKTWCJvOTi1YqaJ35L74FvIQIZnyFeJZdEBV3KT8EqHiEEsSRguys
DbHQ47HcmH8sfAJvvSBrlTMGBUNC0FFTNMzfpGnEgGoM8eTTEskdtrcY/RPDL7xq
TsjXWqeFVm/kWj61OWVg2XAv5SLFEffsUsQSv5dy0SPWNaip+MypvHWhkeRxUVNq
tCbc10LwYp4ZwG4Rsq0W6DSgOVdVSLc8i6kk+DJ/p2/hL/fiQiVUvLvFhUbY33h1
zUjrAIVcg6ymoKU0UMl3qhCdfxLxYckWZlOdMnVlbltYZor+Q0t5MOvgSRNgYhJj
Qq/5iCvS/Ut7dyLN2xKLGaBM9ffDLQB0LgOi+bIOalF3tqWwACKv149EBY9Imrw+
Rp2p2kBOxY9Wa226vDOyLAnmc8rDUWd6SNcujVCE6Q0AiDc9d1CNUG5vug76X5HA
tVrJ2Xw3xi6iHy9vDDnSLaAldOZsNrTvIySg++3ESLBEvWUXq+1rD6onT7AyNpaY
7RE2EnUQkE0G6K0NrSp1zNRmgVT2iss8882u2hsw90hcBFLhmYA6KFhEqGDVhDfM
5/rYnYAP3WlMqye56MTjvBkprxionzGgR1uL7qhxMlRI1IKSOji+o686PfF9rOI0
XA/YJOCbp5UDeudUs0O7tnaA20V+7jHZRu2OMG+zZ2HjhCSynUxE6+n8PUB6jpl8
Qh2eR8ngSAw/ra88zJnAmHr+Pcr9X8e3s6zPnEIDl/Y3h/15u7sM6kXTCA5n2/9k
4v/uFqbwBlSTq43hp4swFR/Bt/Hkf+IuI6r/CxmHB92C/JpawCd4ZQAlTK1uQWP6
ixosppdWRmjfPgyUQSFH7OZUqY+IN9Hp3xWLaZvy5k8lsGo/6vTlMdT/zj/Q3Ktm
IT04mp6MUICenAeFhYWfxqORJv0jJDVIhGnQ53wBG4tHGDNMJyRL5rAz7ApD8nxw
nkIazNSAFVmiiI69ZjTjT7j3Pkxo2fw4wSSrGpJSsbryTDLqwT6cdIiZheBP2Nun
vEHb5j8KAj60ibh/vpwnHy+ARGsl8VVMN2tdAvx5eeKfIDh6IHLglyrR9cBBQUHR
367NZrLQjds/5skA1YmXkji7lRcgI0ArSdr4veUpXPsKMb52dn3/2CigvF1qQ0/G
9YefUf37E8gTY7y28jI7SrHUbJYIoFLtuYw/ddOR1GuPB6EmV9pVq3wVlBA77lwz
kfeg/oorKl3kKDJCoIxItOHjcdHKexcxbvwzPouPwWEZPuZ6//EGHNVY9XrSLuQm
m95YpyDcSL2rsvCxZdcZDmEf1yOlzN3Vqhm08BOVhl8phswOG7gV1LmEMcLKcRcY
qiIp1mvG2OVN0L8fZA+Yp49ph3vvryJT3VY4TqR1bpkV1v+nsyKNQX56hNFE8gXk
YgFc6bDFjAC5hqCrepDp+J7RR8fV2PFyBah/4qp2gVaov9PqwuGfirwkyaFTl20i
qdYIdxAcbY9DY6JaTT8p1u1Hq/R5FRPJScFdVLLXgEpKOOfdpq5APb5xP2bI6DEh
CRX0ialjdob9KzLydN5JgpeEEcN4FGfL4gNeIjGyBLchu+tDZ4gU9bFSg9TQ78Rd
xQER1GkhfiWpNnFpISUN5eYIBgoLYOs9AOZSUg7n0VoGOhVnYGXhYq4F+657PohH
yy8IqPKRLZzS+PQrfhGl2//FSxYf/DsAliWSGAFwcevP6FOY4vlfinhnjYfky0F+
GQ2L1TXA7knwK4ffoB8NB2mDcJIYrzXCysV88KJS6sYXvadblFklSXQvRkzkyJea
MDDCL5DqoMYjFAlRtXfyA4c15/BkHKEqqdjJ6pPhfY38SgnXnFDH4ZlEVbkbChbp
U/V0KjtTf2XQuV+7P3QX6r2gYdEFqbFRx0xGrxflqVEcY4ybbuJsMO2bPNgLd/my
SsxKGrz85TXsfU8sfZ9BuQgz11HnwSU2KQkHg2LoDSwWZY499PP3kVMUGEuZ2tZR
//+wiqMLSxlihpfKeyQCvS1nKQDOUgkCM0AsXs2tYRC+Jb22QZh+ELvvCvAOfvy0
Fg/2ViNYOC4Jdik3q35+5MZaG6qJVyI0zlhC3bfcqR1rX8PziXJwFq8hvdt44WQ/
OhNpoAy681i7/O+l3v1j4xrnRWfXaA4jBjk0wAR9WMIFO1/c4w06DYXHPJ4A0CIC
UbWKUWacxiTX5pkIIkoxZuyqByD5/uRyZNko7v4mZhzlUDzyJNldiLmiVdUDXohg
TbxDcjOo+2EJvtYUHLSD437az20kZ/1lpWX7jVBz2ixfSUU+R2rvhKRYlWLOeFZl
j7mQlO4ivcejD/8jSCW+OeYT/hKJw+WYu5vTrGfgQwMZPHwZeoU6RpAkSOcXH9TL
X1OXyh12TN1Go4/FEgdN7EV/W5Exmf0WLMIrvN4C9sWxZLA3xRWrPvmPc5vclsg4
pFiRbCS8CusYQS6zquxaBXIoAo+088uGq0yMzzZXIt4o3Rz/wOQwENUkO28aBGc0
am/oTVZ06s4z9fY3eN8ypUGiZKz04tdY9dPr0RUTjKzfDhuwqWHwuDTEQ20pTsgJ
F7R+QG5E9gHUbDDTZaDVlAQ3+dMCjkA5B2zCpAdBNDjziVhgUyZDBpqqo4hIlaUs
AjnjSeegwpfdUIF1LLVFIiAbE8Mn7NZxZcofuxzxxT/Y901HYigQa/2gTGzmaYCu
5u6kLVTOQsNrGFeYnlSf9EiCk00HmirWQDhqbDrJpaY9P/9khn+PqWVR3eA7e1aD
7acmCEiNqsMVN3mLGJtulfUnaiTt4vAY+M3n3Z0Sd64morAa+z4DqOP2XdhsOJDu
y5eAja6vPM3V7knIkWQh230r6qhn6yw9etdDd65zlfe7UzcXYBy5eGD1wlHC4y+l
LXu+EtC97AFEsEJt4bAh2Lvx8oIAP1CdSk421w/u8gqXfQT+UyWaDs8URbG08ryr
MdIJhm7K4GCA9CYcVkMr7WSUV372/T048wSkrF2Fr7UGmmocsBxAxF6LvT0C4oEt
vEVtIJHGW9OjmqEXKgWNBMpgjwt1Sicurs6LEapsiZ+k4G8r+O9wl+jWjDDxGE7y
iT4Cl3AkpVH0RHVL6yB0/E8B2VM7Q5rEk8lTlCDZhrFoIZGATawrEKVZq9VYwPBk
PS3N5Nj03P4H6DzcEEWa6xCjKkFbeRrvsatMmnBSmLdtRH1iEhE28GmyXagS6lY8
dgcPuK3dJlRVIuhaG9Bx69tVGp1CBGygN/0ODB9q3oilWuivmAvNGkTJmv16+R3S
6DX5qISaxKYwQFtQZiLLYWmBqiNGqT/IFuflR58EPpEX5ialw1OzMeyj5qLgTQPL
9KbUnD29clf4XS2+P/6ctcd94ODqN6hCHMbAuHVO4G1lk0Zx01osSzGIYNpdPehl
k9/UGuTOHkUvqxDY6QtRsCOdJNWuQSNSrXE20cqdyc8NwG7wVVNAIzPcMErBtEf9
OylwGlymjm6Kt7CbFVbQTGAWO6Id/SCBQg6FzmgHrjyes8dhReda5rqJFHxSKrdh
hkOxlXMn2Uc1zdNq9eEfBRLUKgEayI7vTxlhIBeZ8tp5FU3gWeid+Gj1TovJo+wD
lpVRXmu9p6kZYeZx+Q+uG44OQQSuu4GX7h1y25CQVOsTqlOdTLAfyyNXhAPeCcm1
MArQ/zuy3AmRn5mtlBn4PVAXsZZLT1RP/2koTZJ/No/HCKME4vSC+ZDxeec9Y2xp
CN05AAlIiv5tQMtjWhsZnipOyLlDNG4K1KjbikupHymTmaIuCTGZGm3ldoNfGDA0
cURs+8FpY68t89HstNrOogQ4+j5BBM8KljqWkUljS3/NmRJXKXwwCpJVvbRQxedO
his4rwepJj090rVVfV2+nLykotKto+StTiosQhCzkxNQrGXHdz3t2FDw4wLnrwbS
OfRiws9K4+opr+tpDyugNVUFYN+GSoh3j2645fuZYd3xm86j3JTm/th3Y0U/sNTT
G6SpFwjqlvdB+rKTZgEAzBqgBTOFCzSQMJGuvJos/IBgCrS9yJNV3U/r/HvBF5LU
1kXzOp8ZUfk1TxTyvKNsDpGlruWz10edZjfSlJKsUbDW6h2TbUgUtzrG4ggOas1L
DkfCRiCbDgZxPehYjyRMOWYoQakkenrI/OOeYGK0fnG3olHvNrxs+O6xEs67s6ce
PppbobGTCG9XKGNVj63Cy+dokM179fmPNGDhU3IdTmx1FoKYNDq0FzKAXaolMEbx
Z9ZrSsQM1WgT31G+O9i8TVQtJ/miC7DSMpyjWIamqHc1ghYkqJ57rP5abO4tKBHB
CPv0gjte3hYtnIRbPuukAAxAIRG2Zc7JjG2l46vmnn2LHpiAhCh/SCdLAeohhLGC
l5gdSXTEJW1k7eN7YzXUZYOm4lnTJSqI63zoFtLcO87/fTtkW3u8HaemgGuUp3vj
vEnUdC4SDLYKLedBdCwal4O7UsnU0QW2d2/T8LenYwf89tQWGnAkeGTuWxOEpL1R
/J7L3zyUYPgMW03tSElYxiZQAgHxEF5MwOAZGt9UzMTaEu69egmJxCNUPMqd8ey3
AKXFd9hhHnS1ovvrJdiNzbpYNeLr1B6agPwOqCYQRSAwGGNeiGn8l3SE/IXGoPb9
c57mrH7psVzgVbLz3bpIGhazFCgZVQAFsBVgB76hg1ieo/X5jHeMkR3fkN09pOZ8
cZoJK0NXo3eKwJUeVej0qJ+3pIlpheKtwnTqu7lavyjthzni6cJVmi5q6I201ONX
VnbayqvD7SWd/0FgfrfH4LwIcLP4QBklFBnNUq8q1bJ0Rxh3jwwCsdglmLZh0AOV
E4UlSflC9z5BveaoMVMfPAsQmQqylRnLcsM/4/mq7vLUrjIMdNxyxoSrEGybHAAu
UDnFS7pl52SNYUpS//HJdwPWYFTwJ8iB7LbxyebMXr6zHJ5Q4uy04iJ8pKEBM1aS
/e+6NdzKBUoxfvMvHLVDsyU4/+jiqwEDy8v9SgMJv8tuPBYJepupVCbQh5GUo1Ck
5tXnvWgdtYLpn1vfzPHNlZYx6CDraK07oRDuUzCnLHNkwu1BKNrd1nIzaDETcMME
0lFIp2l3RI4hh0qWB09F+cnUEz+NniTVBn+xaa72rJbvGEPYDWW9kF/SZSC+0MjW
DMNFdsN2+it5RqlbYMwBpsvRNPpoML8/8BKximd2+vWjOahOkcXP4ux2nh9G/5ZM
dI73Z6qNX3lVywJWrt9tnWAtU/6DLaxPBHQ/YBMeZlMzVENzqQGtas5pVq/G8tR1
uQHGbxZK6/NFYBV617l5aDhN5JvRa6iv6Ew+09WGeMPjRYWauE5/aHpcxwDInTyb
3b3l1SbsgGkoS/nhJamRPjWNL8NWlPq5fasqMglmZi21jMNvrpmjTHP7eJJFABgG
T3KXtou+4IsXizC4Vr42MK+gaS4cthinu4nzyv9XpV0e9WgnwBrfqK0mIvzoxBMk
1C2+yKyP8+5ewy31+hAlZbyWnBDNr8D/2+CxGRXSCXk3wYpCGk7ypWuGJpZsfe1O
/cTc8XG7iX5pXaFY6ZTsQ5hlPDsrjLZXxXNG0UOgfqOxjdR4qYrDTZ+HwFV/4p11
by1jfIOnrngDxyBg+JNAcFJZLgT6JOxZDcxDkTBg1B8nmYU9TzH3tUSkYXLcNeQl
3Dlm2ZSuZ9aXaN8DnJQrJy5tKvJtvETEOaZ/fLD7nM0adxeeWKozqEf1KytzgDO5
I7vW0EKDpGpe2NY1S/nKFw0e0xcG4f87/5FJMHFeRJ3cyvzdRCEHllyk03dux5h9
IA8+AtA/X4JEEF4iD9jZoy9MMcnl635R1hTCzIX2UgDy/Tn/+XG4YCdfVyKShylr
OkUcqKqKEnfcK6zAusd9kE3Y5W6wOAd45YsYpoxEgOb+BXv54uvATOsrBfoMTbkb
sTe7cNDIp2cqQg+VVtpyfGHouQIKgOaZCZgGPbIcgZSKg8V0Hssel6hsUDGnEzxX
YNB/zGbNntoVi8YhqGN9cPP7JEUSmzsqxpyLXJa6sKS3sFRLgK+v7Dyf2CmR5Ii6
iQYDmv5S9Q8IjDXlZ5Cog7KkejtV9JMAvU0taImNwCrapKqPbcX9YlkA2YROVN78
fdnJEY+x7VuMR9IEaCbLpuKM9Mu5l5lWcwWjDVOC5h8+HfZhvbCo1m7OTmEkEd2X
WStzA9VyS4GEadeuoLrF3HzT9nTSNtfoA/zazBVVY9bTJGn8iBp86SNKQix3fpoj
qHfv8HtzQkIAginRlHhZCmvyoNwLRp0f4lPvGr4JagcmTPEhvPwKsnGghZcofEeG
HUvQZonlpMeZu3hO8BjOYo6Xw+aKeuWeS8j9FnwMe3ILVCHL6FUWTlP4TbSlf7EQ
WaC5/8ZpxOCoi7JmG9ZcS4+EN/lJWrCjV02/2C54bsO6NipsjREQLCejD+I7kfYB
/G1O1YK943ZhN4qtXvh4aJ85jGEx4ck+XyOOio/B0DFh8ra2uXFKvaDW80nlRCu+
rZD3MjPGg9Q8gaUbhLTQi2RFUhdDYlXYGSMFfWbXBH6ZUEANb29QKo7do+MAuAPD
BMeJ7YxmeaB6vunNgthqiQ+drwo8Akb5emBBGRCydkmkQn3cn11cVBam0P355hsa
7kWJPY6qJ69APVT7scWZ/qTAMhYc4IbMUg4UqKXccUtnJcu5igHsOQzr/nict9+X
OKVCdtJwSeoOkKAIjY3dWAW6VPb/pP6HpQubKhGC00x73ozLrTzH+CJB5KXktJO3
2MBwwpGoToRt8rdyf54XFWzxD0DO0aTmbvh/7T2EmLXvBsaKT6CQRSoWsQkaTYai
O1uHNmIfVFgufpH0OQb7xNAs7Ep6RDUcGzRulS9r901+dwBfLmkLZyYTDx/b8AER
aAARNFcOZpwzZUqE3WOzgDNz0sDqzxTRZLioVDbtw003qfUH0/r1bHS6ZAooIsBf
l1ku5zLp8CkZ9dRbntrqR5enXNbGxtiOz1io3Zx08/ROdzpCvxC5a8koh1tuckj2
QD/R3oI+aQrD2LjZ8rbGsjSQ5IynTeAqoF3l2vOrw6ibKLC2sPzYZLCX4fxlGs7/
palOpSwQp/SnE3rRZH/01zMGz7zno2FB45zgUvfamCMasLqVeFJznAr7gGjxRPnc
eXSQ6DkcnCGAlITWRez5S3G3rLwcKdIThDMmvmenNOHwSO+58t2+dCXVFPXk9p68
iGyfki1joL6NfoBnH2PmKtwM3gnbh5489ZBxG0T9IvmmN6+IqDnUEJuSUFQPsCPS
HD8CjZljYV9s8d5zkgkjgc4Ai/k+3fKnYoKt9u6+w85HYGO+jygVbdd+GiCSiP79
L6TTTeR2WKPKvbJfbXZVwzMYaF5Scn9Ff4ffmgbyF0Rb4rp0knj7Pfe3FhNwRyJ5
oRvqC+u2koDxNP10BPPQOvKI7QV/PnLDPdAHLSRqae9YgyVap1LUukx3mVKQsK6g
r4iZdlryEfvsRs3UkDqU90RZAVmeJb2FT9rYzvD2mzu6yWfnN01+E7zNZkiKtO+O
M36Rf8SLTzM+Z9qo5mGw6AZJ4iOFHroIzEzQaslAiJGrRhLclGiX+8nbcLM2GCFJ
QwgiTczHmmlxL+JgvOakAH+hRUYKh8QkXaNzudDZaPJPlgzIwzPMU0/auIadKOu9
mJlRXiGNoJ8OtXnMFFNMNX74wE3S5oqmWlnAQXNMZDDXrlsq0bkJ0+CWVIJX9b0I
wbOKdkV6URN6jWEhFxLiZOIxaJDAYxhqJdWCrx5GYsELSPVoo0aI6bt8Ng2vFwDY
lJaJ60DsePQav0iALyZHkuKN5dkGtXTGdKMSxrLDpkTNSlcRHryZ/eXnDxo9mu99
FkrzAHd52c3XmA5cxZTG2yiwP4IpPjc3zA4Eb+e265upRy8Ije5QfccrMKzVv9sW
9RyTNrYkfqWW8HXAiErnPE4i71XG0H8OU023hky69mlr1TXsRLIMXJCXdI5NmzQj
HdQSISAldFg37KjqDJjB9s160tM+hHsmswzYGNZcc2MWii/xpriNOamS7jGo/pjG
250/p4LYjCUIvF6KbPnCQuNV+wcOValtXD0Px+Ow4N+discYCKVkP94S2fL43jcs
mMIyaQtOm5MkYfdz9jFDOOPcSTa0UDH1OlpccVijnbDatp4vAUIKXY8sp1hfLJqU
7qvTe5bO0kWMjZV7mRZ57bASGV6lza40cyk5PvQIbFGane4BAJ4zks7NALNbny9C
z8A/uu9Q3MdpPtz6FITMooMOnY0hBaywSbAiwO2XRw9gqtpcQrtVv3B/AnPWk4lX
9sWBoH7+rqHwFZ0zXMGzAkeLN5sI0P1O38HoNHBiOi+YgR7njL2VuIPaUTnxMCEM
6CcxC+FCVgki1wlXUNrXQGosrOKlLwvam9pucYaaqf2s4SxvBXNRFZ3NL+TPSAWk
+i++NZs48M7nGaSwqeB93+Qrce1aOY/QCX1ZbiMPZraJIV/Nqa3zRq1v+XdgACLf
Nzdle1r4D3o+efs7lXqAN/AGVptwTh/C53QBdQC6FMAEDNdTvq69cZmkDeY0wv9T
+AJKs8SqeUhaeghDbZUsURYePS0KJ0ovBo4dQw5k4zDTrZttpX1PI+CSL1NvsXbJ
dKsYGG20fvReKK463I95bU+ikkaqPQDyh2965id+TcGFzJLXKv8nJBVezyBoQEl6
wPEwNW/MLFoXalBiKuDqNM0m9ZpeQXxMWjlBffZG4UwTw0VhdT2U8OdqCgABVTkB
MYHYB56pV3L3tEP9Kdqj0bIu9xjs1VBgikAXgmqlBHZsy7ywtZP928HSzBmnKCFx
IBhHRYKanVS7ere3B5d3VIfK2vDP5QNrgfj3yCBk1Hx5gJ+uEUU11tgE9N0ftazt
9rRw85kP/WiL+h/XZi6lglP3LrxelqbYACRQVAB6xS6y600k+QBYvmw7s8YI8KE5
LnPPqHsj7OT/kqf6EZuP2aRl3dgvpF/WhzPERqAhv7p/X4TUcBYpNcFlnZFuN+12
XzBDFFv/NdwBjI6zNADp4KBuVy8v+C42wyoXgVvbuMZfDecS/Yjl+2S7fqZIBm9h
GrGnW82Xii3sJ6+IG87abF3d5y/lcgNXcpOzCKg6YxhISdc576a6kVf/eKt1kww1
V2+3FZshUsdzr5eGII/JZYkJCcMuctciCcnM0DZoggZqxRyKy/GxXwi4L0dgh1kZ
nq1tbHinFK/N+Oliv6owglFolMc9DhtApKngRavxSHP52caltOHnKuv20wrq1tpf
mXKGr3yjOYKM/tuUp0D6Bt8dmKvQrYtCmneum6eVWV1B3CnygH00momEcLadwGeE
NcBduzKYZOJRcQmqxM5Y75SQajWVaDPO3rrSCHl9l9bc6Pz9FU0xfjkByZqZwx9y
VdNGvAaIDaTOCXC+LPkPD11jBEHLqEBzkW1pg3DDqhZ+3Qp3iMupcRAwLwByv0/8
mS7ZppT2x/MIcggKN0S0pbtTZVKzafeum9kdEGFAzYphSVKN2c8IIHef+YAQTyWt
J2+rk/QgAC6sFRoRWT29ZKmeCHJabsbntY67Gwl2SLmncFFXpxs8pr30btWJT4N0
vvVbJijBBilbBebgQHTYNCqWopnTqmBBVXVPwoBf8uaq4biGa7PC+gLZq2jsysmv
+j6V1Y6jdg9PwdSUE0OvsbUZ91nzUtSGx8HMJWC3665ZkcR739WImFSh4qZDlGjx
xfXCeABlqXIzTKJtOYSKQ5LckpMQtDfRidETepFJRDe3nyUxBKkGxCOGMD8bxuSn
ahsZ9Kv/oZGsWaymzBLfp1PdkQdDT09dq+03AwzOrT/9BlQxdet8yt0gsmKW2psJ
o+gvWYX2+fvS8VNblcAhywyu4w/+7nPDY0SljxVS3ZxYzP6cgQux4IuN3nC0kjWM
yt814FRe3u/ijbvba0YdEkSMBVY9i9+fIHwDt3SE/pPVXHWT/D0hbvIOP3f3qX5w
4k3sDTO7j9QNzX0RQ5p/NK3LhjfuiD+x6ssDRjc2BiwtpoouJXpugd97q+OJOGE8
0m97eQxlSzSctIA0ofIFy/xQ1Ju2XjlCcoAnAArMvdnEjwRGX5M1cW1AkDFI9cyR
mY5h7bCAPh3drrafSPgnWU/ICYJXfCh5gkD5XE6owmkRUbPx0qHQJdVvbbk1xWJ2
pfhV/JFTKn1mgwM4v+DrdcpC9iVOVIFEhCOPTHARwr3y6tlg3xPOOuRk7wt4hkqd
thfNW1Y4S7NpEhhTpMBjBLXhz4QPrGx2+NKtzkRM2BhYUa8WrKPrjZsa/ios/k6s
hVVoEB2fsRcTS3po+OPlPkcUJ6lGsP6b+XMzH/E+AG8I7jC7n7s7Ck3L2B91s5Jh
/19zHyXeDswn+0n8fhMWJmgPbAGQjUpfkqCeY/AE/R5u2D2kf9JPk7yQyVF/2Eju
6iFgVJZIECrOQJfHVr6BCmVq0CmWkpkBJ21WLvaQe0Ce9+XiXXogrzRr9qA4I++S
LLO46nweimGYMOk3haNdTczesMghKecRZOnwxS7UTS3lgTgkVu0cbQYUzJIeWFt0
G64DVYAjl6CDpoW7NFFJl2jsSYRoBCDdrMP4gKKfG9qDjkf50Ox9p9Bo3T3hSA2c
2HL2rdVwacEpYlGlsn22uCU9hK/UVyim47mBY6qTbWSLKjpNmai4CHThA/X0Hn/j
PyW6EJBscI1qKG69Afv+ce12fpljxbHkG+bGKo5RbOmxpOg6OtKF0okxto31Iafa
O4gGnBQ9001ks4g4QaFOSBBwNEdSiktC9mOFNaYX7lUWuLsaDPK60ZA1BhKXRnVm
aoSzJHhjeVKKaGp3UCygwHqtdZOEH8OspReUdqgF3TeTXajq4n8Gl0vICTE8VRIN
C1hFw1lHVUQ/Yc40BUIUheySIXdXb6H11Tki6QtTNSkJgw4cz8io8+JO8AaPj93I
IFj35Ch84mXr7dhwPS5jpjwVKlk2bbwVjT1ZD/ExfOJkaJ8s59LWl1Ro4IoX9PGO
bZ1CFjvqFpfH4r7uNSu4KcSFsuUUqy+9E3tTXwjIfUBQHPjgrNv0VSShf/jMGES9
0c9pWW10gSTiEdsTt0tV+53bHfdaH/mMTcFJ/U0WJDgDdFmjXs7+ouAhxYpWTW2Q
CySBDo0yReeJBLgSu+3atsIxpRb36XJtg6snBeVF65DBTKkCt2Vk9F0645xb/5pd
IpW+C3hR6kavRBRuHH0KB2tqcbQWPzd+GlsHdtUhF4I8zlFUYZFohEX8GhI+Tvxn
NxdzIA+78/KHrQ1dKfv0x9RX6dt9SJmLk1jkqSNwrrtWJzb5wefvv5FFfTgyLGtI
kGER4BRO3vxgVk6KM1ZqfcnkQHILOu6CL+93nq75lrQXkqgXMcJ0Ghh38xzafztV
hf1W5rA3m3OWHLhO/Slxy9nfMhrR7Y47Xv/NmuITqTugnJvub31PrsPDybkPKwrq
1/qYr2xQbKvCPP4O/v5XZomrmLx0vGXV6sqNz9ZgWKL9lrwczbTxjhs3kg8mW/46
pTHvbMTzDvzLuJD1v5KGdtHMA2ei5QUUTvOjcCHl/8z3uVFLriUz62hN1nWKrRAm
qTSOEBK3mXg5Ar9KzB0bWm3UNtZnfG/uBvt3q5N/nzahrhwoXAzSXTFJ0b+t9jhw
KK8X/m95zIVxAc9tZUK58hNPEs+ZDF7aOZuoh3wlV7155aZmH9nVJ1xjdKJlHzgI
z6p0d+D3wwsN44KECu1XSJHDlKxTHRnhWV5q8WIEQNTi+xc6tt09EqekiVyoIDAp
j3DNuFUec5P2+NMTKYz22/gFX5StWJEuxS2MDdQt8jOnE9OyNFXu0yPRZ7M71mAH
4j/zDcLFgD3Lmcugfm81q2YhVOry0ZiAT8jhGJudBUNVtY8+10qj/mG2/uBBqGS9
+LbgccTszqplQjPPOCPZy7NOwBRSeNaxqveUtlcnMUVKhGck01BxR3sdYO67e1Xn
OWI5ysSwrNii/9A29Q8EXfI6D1WNKwPwvE3HK2IS0l7NGhT0P+0a3YwyGjSngq8w
E1FwSQov/atKSn4CrP66gVSW5F0Ueqxmd+0rCJqWt+PAOHxC7DrHYQFdur4zUyIv
9mjrVh9fa4S/9sUjr/y3u+SJPLJckX35QS8QRfy5nxcfWZGcNngcOqQ4UxFU3/6r
fRnh5Cb/4i1bk6HoUwUMyZwTBVn9C3uOlkHL0v1q3zuWInZixNe7tjcJC8ghNSGY
a++KySxQiRN6EIynnYCMFZsPRC/AjdndX9jGd09HkXIcNqQQnapNIB0RnjS5YXU7
Sl4X+NVgBlOnlIWdFtGc1bYjj/BE5DyL/dPhyULp8Ym3pL5R2sUB0Ec3KKsM73Ez
J7tXWo5G+fUF8fNqV7J8VQX0uVExM9ePjZMvDNP+IWKSPVfyukjucFhbgK7o6V+U
W1T6cSccdXlvgPjv5NAO1evI5DvzqhWQQsiO7kmLU4abx9xwJa/lEQslYKUTaDuT
QqlrqaX7IL9xsj1i8sa1jJ6we1kiZ6vi9oC+pkrgcX4+2r+t3f3HTzS8FBliTydT
v89jtX64bth66e8rIir6PgLTt0WSYc0bPhW+6EV/8gZl7aq9EalywBFxdeeA75Hu
xyNBrdboeb5OfkWW7pUsjI6+1JYePK1Upm2KqjHLpdkj4OtAOazC+58po2BiPKlx
BWI3M0F+iJwzOVTIHua589jf84SGqm5cZ1WCjzI8sPvdIzY4Dto4zoacjcbMrs/I
ZBMFWJNhlwhsKAe5Y9JKaEjlUdf7c3nfaB7DXkfIoeTJkTA+IQaK+MzZLdIoyxcf
ABcIq/FkNCrjMH/nro2YrCBCDl2maGFYQuZTpoLJEWVd72KedGN5ro4/xBn/0MmW
xr/eNTt1tJorxkMIUSyAzP4U1jshrDmPJYv1J9+40MCHo56pb7gQh+gB5XtqYnpY
Y6XFgs6wzr1dcODnhqFIn7QmdpvtGP+JVZgpptc4D4V4I3qmZwSQwpE3ml1geR2a
UbMJOQ4qpnNnE4o6Frh9drU/sGX+8Zr+TLU7l0K7D/vnkbeLptu/HVpDePBu7jf4
ZgIQ4RKEkz0qqwDrBqFDPq9QFbsCWkBzw17E+NRoUlDb+B0dlt4fMRKuTZK+MyN+
UYQ3NwSaf6IE03dLJYvFiu54bgOKprkplIGZDdGW3eINYnZA1XPEWShaCxft6m5K
h4PjiD3IM+Exxacr41Vpkis+A+wicPeIEzHofdc6uHfXFOz1l+Le09wtuYFh+3mc
wUJ4SLpFWuyHF6XQUTJq7YjJh38VZhs0RCuO/s9PgNKj5sTlivp00Tth8V4dssRC
ObZV/YZVQu7siFV5XQbjeTu13FNRcds7msoFsn8V47DlvTHSvjOgdS/ezJaJfJmA
NVxAhJSw3jR4o+JyNcJJ2PfUNJK/bFuuAInMGmIT54B1airFshpnet5HCNiU0Znm
pvED7hcVW98MnPynHOR5HqjcFSvVZLCR5SZG0+jbbj3K0IRXN4+SCAWllfqgDGY8
OOoMhFtmoocO6zl3Ly9oqN7BzQZSlYVMA/LQ1+QHyksOLst2qOqpaV8So0FDiix3
/FZSHqvKJ7NdPLR0/ylsMBDMoK/7et7/oWKO6YGhIovm9Q++7L1Cds8Zr/9jhDj2
nqZ5kj872JgGyHLPH7ufwD2nB3vX3zTZ5m8uPTVPVjS2WTkT8ynIYgE5MMZ7quJ2
SsDC8XYc1UXOZQMFqYa2Z05hKts6OMJDOrC4P4SCIjosPrcuQUSuJvHHGf2b/Sbl
8ELTGwOlNiFVtuXxvsZVg6n7pmrmM01F2WV/QUS4hFLeFS1QDzCesXcaV4wwCnhD
1KmnOj2RuBvLg4++g8/Fdigj49IoT2LbNyVr/EEmz4QGevIgddenNRGpRjlQ9mA+
5DRVni8ApBXlNW+aGJnOXgTdwwIjnO4z3JotlgEFHzkNIqYjkajTnOSzXn4uHlGP
nSHc+meIMJxYW5PDtdle5f1oopiS/BSZGUHPEr7lo1g/aQeR5RyMhDEvVPOpPysy
J3QWTIeiECgrvB0ruYITPfLwWZOf9NKeY6Xw9M3p2AVC2foazDEvu48MiKI62tka
tjTOBHU3vCqGiJ+R7vj3ATFprxV7Orpm2vb1e/rNoTvQRe0BfDrOeEbgi0eP1ig7
Y68fVF8UEIEz0bbhh7LrYBgH+Ogdi1fkpfdTSE2XzkKGj88w+r1/2LoDRBNA5AxU
Apoqx+b66Oqc88edZn0Dv0bUICsV3Wwd6COd1lx/F0q0l+kfwjJ5et8+ARt5hZxz
mV4hUtP4iB8c7R2Ms4Esv3eDsdgEGvU9LPJiaVViw2eLv3t34FwzgdArO9V1XaQc
Ic2Z8S40s/FWuJYLS6ubr4XugzjzWI6hfpSqCtIyfAkw1xaRPxB6pThbnW0x4rg5
33ZhH75m9GfxCkrZy66u2EUNoVkPgAXsMkRuNVRmoSyprMpdqzuwD1MwQx4dNw3b
/XP5g/tTq/NTBruMy6B5LT1u5jd5wldPHdFE/k9v6XNv7Desfg12FO/oE61M1nPC
+jV5UOJbaHBWTLRrNf+4o5fpem8YvE2mwvTe8v9OJ2qbcRMnqHfBq3Nfo+N++M/2
EFtRDFMmWud0o7xGZ8UvPDAAO2He/GbZV6OVL0EvfFfKTFn4/GyXI0WoegmKUhB3
UrIyRtemmCUE49OUC4fb3De/lDb9u8nBZSiHR0An5KOkUKCHIgSMM1XzX7sfP4GD
DKkzrtDtYzgkuq3nO2AzgdRnhw6WQtv6c36Cz1zEQuUUJkli3HOhSfuT22cd5/t4
2V3Co75HGKrVgRdNVJJeq7rBuMOsYRiXMLy3kzeq5B7KWkTYoU6Dwyo220y83GIT
1/i10ATV5cuCNjZzuG/mG5qXieM+Zpe/KLUpms7UvSaHY/hFcqIUpTnuw/qJg75x
k3EQlIo5/Bn/mQDWiidSZxIMTmhx3dFDJr3tYRINCIZCUmWutieSwGQa4I4kIgOi
0ZFBNoBccFOeoNLbTKtfGhDT2jQP8INybevsMgqjDWkTcOosSTs/yKbTNrBoHvyA
KYMWqnc9Uju7I9U7I02s3mVEM9AX4LBjLKVT47tq43q7QgAy5yPPoIh2TGhzFnE5
EzmZu6q+552hpdCzH4ezBnFrryEa6WNkHjHWsngiQ1o/jFI8YDuW7M63cMwE/a5v
amRcsdDLr8v5taiUFB1RR3kRwrtLUvrS5Qe9xy4b/VNFVsabDEnPTi+v++swpZ2n
Hvuva3kcY1ZJqhZALrYpBzA5551hAJfYqiaF8ryvUP8KFoLpkruuF0Ht0hexxHsE
fhJP62bsPlyaGl+R9HnjItm5pw+LDlXwr3VgEJPvffMYcRQ2T4BRth68Hlf/1bWz
oYjqT6B49NukZks03eJXoS1ux9vh7NXevBeJ4feffVrlxVd2CuxuPVV2kV8KTJ0E
dBzDyLkG7MSqcY56MVRij5vdHwh7toEypNUlI7a4j1w2lCVlPQ631JpYzC8lrc06
Vr7iw7lj5BrTgRuTC/wKK3hxTjf1fJ/jlz3kSJfAhhpelExok+18LNdemuwe29lW
Dpin3kdQFO4V2S5XODJXhp+LknRXAw4ggaph6MvAr6g9FCqaqQHDJ2aU3dXirPuV
WZ/Tx6wfv7yJ+ambJ2Y5wmnmAG0Z1DUzr79m6OIyccFCkXfCzSbZhGe1UdDdDlnu
3yGtBS+KXRpsbWiHbr1Ikt+xjiR0qIbS+nSRydX+y3hLtKAAXw3gGqJtufBpxijS
Apvmmp8EWAeXxTpp9KW81CqOVBQpJ8i/A02CUAE/fPKoEvy82JI3VJGe2WGXcz9k
5MV+OXvioqqmgePUmJqni+JYHQFlgRziwDQsGQBvdrRsRm6MLFst98S2CTbAv57k
35NNxDNireS6uql9wXq697rP3xjGyxSmP5vNOGN2v8z+el4uf4/jVGdZCjK+qQRQ
1peKGnHyCkeOPM0HTMunhJWRHOFVZaVgBMkicoQHFj4u84Q2/Ki1Q5YWuuVoXsGm
pv80bSB8ieweqGR3BbskcaCANcRXiPY4SiBr50X3MTRRiW8mj2WkitvZmam5E83i
He/gUG+/sX5SvcVkZ0TZQmSdMqWi0N9uaBJnekNpo8KUS7ZigfE3xVIe6SjS8dOJ
ctd+Nef38Sz4bYpKPo66gB0LfRzl6Li+olxAyGS/F244Rf4TbDlCOVRHKEIPHiip
ZkAjgUUMb2r4vC9CRB8bdj0cVZ5AnUmT4KsTwD/qThEJsNmSHh6cBagnmB+ZSj4w
yjNqcaeM8E2D1mUHfcawfskVml1w1rvXX9N4U2ZAf0ruwrz6lsrfyb69WfKhxUqV
v4j0CDWQkCOlX1yLqCDIh4MpjYlt6m6QsyJaymamVCIbr7ytsustSRJ+n3le5COa
ZMnnwZIdKPQ0uWGtmLSumIfFb3MH4KZjgr/Q5Xz1iFK17yZk/OHzKfW2T0nAfBrQ
wD4sv1NWcTzeF62s86wjK+Q/PNHFiu8JDjrXYDmNsmA9/SiNXIIfGmt9fesTzRAm
PKVPSMKGtraCQVncyC229lDcH5I1ctk+T4wdGwBrHMs/Z2UgnjeGCDrE+q0T2RoA
Et47oN1ojShGFC65OQFAdB70IDBD1zj2+zduN4Rq4K7ICocL7UDG1SquY45dCQRX
SGihqDhe7OrZHdPbSw13I/Qq7DwnuEAni4m7phpDMM5JQ24/TivReo0oTuKKoU8K
hEQEpSbgtlDUmx9lOjmSMPm7PiSHmrsPWVQLS6n3n62dpSuJK0NhZCHSQEG650/8
tyYoDa7vRm8IlIwxSACmmdcA72KjTQAEKPXhWDCjiWUmAzVzDZhSFH0q31TFFPC9
cKS8eBQY+64EjbdYDw05n3toQ/5N+c2rEg7ukBuwJ9u0AfEBTVnzHgjYCapIhWKu
Bld0xMDyUP+1lDdXZ8ADeGAeac1G1qzTqag/0V1PIBO6xk6mk8J10pkxVCvBl1ld
wR3PD3wdT5pFwHZ+4J+ZwJ8GSFedTdEfMWNJCco/Jr+D5EnQqBAt5EN2PTrsVS4m
mcfzbd6fneVwFA0pTHHwBn2AKJX4hLFYtuhStMYXmfGXd97cn1NuYXNoHiV3boL9
862zgiA6hJthBx+qKRBhOUL10qwJmTrGvVjhaFlqQJZeaHl5sDgJwqcKAPE0fcqs
ZWVOjKHmUYo3PPDVLNxnD1exOQvhGREiAJ6s+pOr5UePxg7ny8JZpTKWNensu6IV
OGQDE+ALkMUmA2xQdvjnGYekBGleyArk+0YMpl1SWT/ChmzBiLXgLI9HO5oynhWg
ZCt9LLqM9OaAjEmW9nvRkILK+w7h+dDYyihnx6QhsAAfp51+5GlB8WuVnIF8wH9E
yl7GYfH5KGqpfMu7dy5frsvgNpSNGfAy++fh3ssrKoWxeLqMSUhVVx0dX6wmZ6gW
UA5x+FiSGXOqXEn8Dgs5/r/bcU8+RP5KSAqU0RHcT2tlaqnCwpI5zWA39XWaJMrQ
KPs2G5LpASu8LO1r4jcm+Anak0moZ3pQ1MyfbJvQfvfLuLGfxYM1WPdjZ815VqKp
pmszqnCdMxYcSH6QxrMlMF3CYBZ74YUjDhiroEZgcbztfqo3kMyBl72XQBptcrgE
63LZOzgCD8DEz0wEGJy2LEPLmgnlxy0FIeojqceR4FYKCJmzmtBzKUeWG6vtDkbY
dBE7pE2e1M5asOUrTG53Ap6S53Bqmd/2jnVnrUi21VRofsflC6ASA3Nfi1Fk8eL9
KgdSkDpikUNUtAv8mT+U9p6+OOgafyFuwsblGbjA0OuZSTd5LhS1uip/+FwCVio2
QEGIDPQO6V6yb8A8A1WE7mphMdiBZflNnpAR0yP9mqcTySQN23mAS4f9tyMC5X5c
35/bViU3WYttaEeZ2Vy2YbaJe8iNe1iALu2puXWW1roEHmfiy2J9qNWL1bE6g/Y6
aQBwitEfNAv1m0UI3hCBcQ43+QrBstqiTEyGQnQZ41JvuwDITvffj6d4NHfGAp4g
qd8oJTQACsckmi3dFcpqLxib6djUw9LKdYpNBTIxQ1dX0fN47tAGSV7QFzRUrUXy
dfxKCdpQkB4fW5niirlMKJ9/2qcWVwWtpBbB5lLK1ASifhNuXOkVaNr17Y9jeR9n
GwyQQ03Q+Eo6DkPmWfJ9tCIW/4iD5bdDxMcpETDrejjl3YlsWaWe5vFOyVfhis7c
FHSZMi6xucxKLwTdXPGDb00rqVpjlW53exAVFpYgA+lpssSNctMh7gz/yZ5bsF/b
yK4F3lfoftqhMBqJ/x25cfENQkkByLQo6P8KH4pJ2pyyAdcazRX7IkWuzigJL7PO
WsvPXgq5rCYkp1mXwTyjzlwpEYZk/b6geNs83z7uV7qblBwh4InDOscDn0SbfFfW
TaLfen2gtaNFNoAQ6EaEsSidNiUL1bKb0qoqGw/J7w5nqBgDf06+icDD8FMZa7Kj
FpyrwZ4RBbRNlAmFwVOCa+2MiBdZB3zrrLWHWILsBt5tYh5rEu56jJs7aNk2aazm
h6bJvBqv2TnwxiFT7QrhZUphKalDX8mVRST5vj2J14Kr0e+yYLDF/pay56l4mN63
0TYRz6uknOv9+fCutyfq9VDQ6SyOhzoCx8p4LbX4UhhF4Mj4HpHDNSnHqywx6M7B
akDuQyFLOP8djeRSG3yHNBCiyyaUq4QX6bgtu6KHWDvPut5IxinsrkHlCvs3vIow
eYizlDdYs20c54nozLym+0ImgpNw0SX33jiTHLIfpGjD1HwHNNIHiM8ykyTsNTbh
5lB7vwmWLP7aNmpoXJ7pZB8fumgDWck2vCSBmSeaxwXY3mSwNtLTb6Krau9GNc3d
furCOIy58bcy/YfoWUfcmpiDzKGE4IgCd80Chy9aZBELGDDNk/39mMEjkeak0tq0
N/Al3xqUr5V0cDIXQKa1xjfg/lVg9F8DcG3S3YF0jKDMfiBQCqHtP1t1+KN6TH72
2hc5lCIpHrhe6RWTVqS2Q9q6pGat2pPjyQT7LaMCITFViAns9D5r3b6xw/WAcrmS
gqfaV+aRIpifeuc451SrOULgFd++F+996+oy+Scr4BXkL4jjjwWlj9h9hgOJbQtv
LIFOdNEB/QmL4qAyY1HugRF3l4Cf+XIWa/Pv2biyYLyU0QbZ9gqf0/Lbjfo/ktSx
aawgIMusRyyriM/MH1Lgmq4s//O7JNz8u4Dd8r5mbH9GDHvlACGL+fkEPNlgIT1r
nckfFNw63Rydka2XwilP3moFfKdXClLk8J4XfZPXmhVUj3hy/gMzNlUHCx/P6nrf
yZqecP9xvCfl7UQW81u7zYpGMhnNjkJTKGjS4Rc6LcDeIp5zqygev2rPtCXzBc7u
wQ9f8ZdT/PcjLO5eC5aS1f3bIJzTneL5PRxgaPE/eGp1Q+sMXhU8qQ1zOcoUWwgt
tfBHESGt/pvKRDLso0dNW7iBuBOrmtiZY+FkyLqQzFGEC9EhstB36KZTDI6lDKlH
1l96n7n+SYLAwjt2uuDXdoJndepAZXjxP3IzfrqvoS/yXdwuAIzGrjtz1Un/R499
k0wATAL6MyeORMdV5Cq69hflau6uIb9uX5jON3ZnNH7YfUB8CaS90bMiorzTU6OU
yu87WfeXeE0+SDuGuSnA5MoTpvzD5Fsm6QzDR3jGEBeMJggYyGLhtBobXgtVYh57
Y1pFezalYCjzQEXMSFwo4kRqWKWoNf0S5BMUNDeQ+HJteUP64Phq2UTCnugedsJY
YjIFR8WnNlPzqF1rdsoIwBmnpXJIFaIYf4XQb6PPk9K+R15zHznjqvVWQ2RtLEek
JuTQi5peuX1G/wRmQu6E3gHiBFqYnQJyU8gox7Z9X+HhjHutD5eK8cXAY6XfTPPM
g1MR86lW3161V8OYrLQiaRGn75P0kQr557E1PR6jyitKLzB0OytRcIYtZI0ujK9N
m4iHJVoxDTTxedb3Nbnwfi3V5hI05UD1nBEENzhCls93vCcgXWkPXSpOWM6AIaE2
pJE+o1y0vdtPKlahp/x5s5yFfN9oE5gSC2PTAe5x48X/7s8MSZX8NxiAtJDx8aYy
h5rDuZO3d6xyn1jxML+lG7NW0kDrMEp2kj7KeRa8fYLKZfiiw9HL6jg/DrfSxyQL
GXDi3Pwc4vOZgRRVeDxLKLQZBcCZg/BZbGweKGg9NwkpgsdjwfGB/1fTE7R1YO7G
r2hN2/X5WYNjkB1sEUyBZYWLb077e2zKuWyAZxM4JwZVquxUAJArZ73Y7NgyVDhh
CGcHJcexpGpRpcI7/P5teN2QzlhHbnccvH116yxHCSOyipHndi+++KhfXsOSuQLo
U9J6DtEa3ca9cbAURElnAREjhLDZz50TIIlQaQHGViqUybgbQ92zuWeF1vp7diW3
OPRH+1YetjyDBTN9qHrpY8L3YCsds0U+hvZc7eCGh0/KAW93+blF8z7j4Ko9CyAF
I17Z3R4EXGaXvlJAqwEWNz5prhJkLEL++22kX4HGJkmzHcmTLCKddUC7WR2X3ysO
6jNiVetc23Ap9h0KuAWPTkebem9GJM6CdluraQZkMrUGJqRRPfIuvVNkI3r+Xcke
BaUAw4hjVOZOQCqI6ZS5wEmpWUVjepREPnhZ99RorJWkkz4WdR35TfpUsxlSwVCl
3SAT8goPVciBsBfZxS9T9E75ULXSblfuw9TUH+olP+uLW3lOTxHeh9E9d6E5FwQh
8rTQ8vJ1+lTAdTpFO40QgNhDMN9Q2zJMJs2OsfdPOENCnLT+msH69FP7XVYq+n19
qAT//DBygPg3AE5F9SIGVKIcOKzc4rnIFQFJzM/cdHWCVmUwqxsuLg5Vs2trsolK
eFy4zbuhFFxnRNhboImxon97mLDhTPt3iSe2e86sU6xK6HTRSK5Se+imlPvkAb3d
SYDxJ81p9BaGGPtfbNbSIrCE5RkWjKkCMBc4VClCgZAyvtEIhWoNMEs5fE2+TQHf
4HJXELP5O8zXazHATaVxXo2ipytzcTS1pI1ZzPIFn7Lq25EriH4mRbrOyynRvtaI
skk/q0RBKEr9dJ46gL69h6rIFJVNelu78/0CswLv6r7IyScTGbO3HxOCx2xG8/8y
yqIGj2tS8DKlS6Mrtr411UtpXx4ePh9R+GPh6lf7Jj2Uof22MlVz2ekg78oitngQ
CNtWmc7fsrbmy9YZgjIvPHs5EUut4EEI1sXDT6B8bmQ+OvejnGuqN66dZkrJgF03
/rIzP8WSZeKSGQBz39fFPQrgrWaozrxqNJwzgPOKxgQlzhz+y8ZW7chzSjHP0Fk6
CqDsNPWZykjMehDaZp58ORhOZmWlVtApC2opTRv5H1IA05e9Zp822ZNpb+wXVqDP
WEVjkBwdBZ/bsG2ZLLpG8sFUCZPH5+n8k3gZ+QjsF6iMjfJiAjTIiaGJMKQ7ZNVY
Krc13TeVhyuLV78H0EaYq6HrR6PrsyJeAKezxIz1IOLZuhcZtci6k3vbkZjQcqGE
wimJocGtIj5WUbE/K2USZorjuzMINwWDHItm7PzyLFNd+xV/AgAPMR/HPQgbgpoT
fetUVsXdt96pcF14IWX9rU1QrnBCpsf+XpDuePLh9Xp7Fq6xcCiy3NXwuQxfsNmq
DSLwT/VdD3rkgkvRyWig0NN++6zNCTDAvdGvWIen8/FKW6u9IrD5Yz1yNMzu/XK6
gDK9Jvu1cEM8pvxYOdCH7Vq7QjGYdE4cCSaEL3e3DTliXiBqeTeO5XfI3hpaBd17
Rv11j/SdmxCrM7SLr+bawWsZeiSwg/k3xDWd2V9QOn/ZWBAmKY9hJ4CH5ZNg8ieE
QYayBHRlvPxN/L3lmiNHSsO/HBua9YNTfD7dPZZd12YIpuncQR3uAtt2TSfOETtg
Zun/e9CLQQMMOvCysU38Vq1c4/PQb1d5bwLsxNQx5fUP5PM7e4W4BeW1dRQQV7Ss
F9YlO+P1v26MyzonDgHWtXNKKGnyimSyRl75eJX/tDPYD2/0HSQd2RbZoMEn1ZW/
zwA5o7eZMNeakG6MptCCMv8gkmetxV5MCCyMsbqk0ii1NIG933f5jtPEpaidhel1
F1c8+/h30aHWB7YjNNvOwK24wvMqTEl9Nvc0YxpXsynVdT5GNwJunaGQqf6SNCVg
lxSFatJ3mKdu1Mjncp5GAK1WMWlRbwqDUPtZ5hLwF87Gpi6R3vjyhuKtRvGlb9kg
FFHsYtLrx6AdV8LC/bss8gAPrrDbfxALHi3OltShen0unLH0HS0UkGefmck7b8sz
e2PJsM4UlmV6cQ4l2v5xSFR8hjYqEbMoPUv2mUA+nD8DV7g9gzVnwBbjkOp4AEey
pHeskknZqhKZglujQhkjOG2JdeiAx8lDksB9D0a2GH9HBhx5jO0cxQ+3oQgkoBvx
gACo7/IMOHNWXsIzshtwJdvKEtS3NONHugIweM+HNtlVKYSRDr0T9sHSSaZk1KuW
SPHU4IzE38bi+fJ60E0ZzI0REAle3ZPiVDxXZs1q0pyhgBhGsCTtK7SR/mS0t1Xe
Iiv7vzT8b5b7kCzQVT7SEiIa5hVRFVcbpVBEVG2WTgl8CjBfxojExfEdrvaeINGm
sw7YRMEgKOkkbETxvUW1P252I6qvzc4ompIPvSbQOewpGbt4nPfJHjDju+pMcIN5
SHjNxXrm1vIkIW7/sb1mhPmvqz6G3km2YM4zzU7nS55JQp4koJEeFa4biDaGgXaS
87qsedaTLUbgONNeXzGzXzf1Nbn9FOqewWWaA7UGQUiTF338IOIaBDqz+jJ8LHVL
8U6Fk4mbm92KdbcYMXA3SQvhUaJv2rm6oGoB4LbtZsSPLHSE7eJQvJZzxrBYkpGi
TU3EFDdBW28oG29Wg9xgPFmsTSeuEtZk0Uu6oH5upDLE2rZreI6Mog/7Xb7XZxIX
g4QGMekQdGEEC+pwng5sh+ajAOOrRRaYbvSgoWttZuIgtouoHcAJnx7jDQKXi9om
83dR8pG5Pny7qgK98TUC2b1eK68C9F9NzCG5FRWhfqEYqlnAxVnx8r90GXWiLV0y
F7zvxqX+QcteOjJDpoN02V8y8X1cSZtijWSBYddL7BRjAdrdtEi0mxMTw5kQ/N7N
i87+7BDO4SmBSod34DbBu2F09OOnmSIDQfQmhchmGdFohUlyxQYdvKCyhamzgwoR
gV71ivcCvNSpYdwgbb/ZpqrZ1Yd8nUr17z7Bm3KchZmJMZr6GZZhuPzOod9q2LeW
UmNPFEsJpAT0RqFqLVhEuuvyqX7YJFKvMLEzwMSO09sj5yHwo5UAkOy9wi/HRydF
boDchgiEg6Ef2YYkukoxz8ocjpScJnjhDptd2py7x3agyY04yNvCYyQkdroIru4z
skxwyCx/m/q6Ofoud9CnVPlsqmFis9xKCm+B5qMMThL/pWWpzIb0RKqj4DsSMXQJ
YlEUlecScNcttFuNZh+Rfrmv1zr1xjaUOqFJshur6s5RwJj29OZDPEhjw3d9166s
z6pGktV5Z/4cA16etHYXEIAR/1fq2/kfynRWUsyvhF3dAFNLKV/MZIr5e2+htmrR
ghwwt4KaQAo0B+gYeHVcxXuDMicuThm+8ZTivjluXY+9OtDFY1DqeIk0ZstC8J9D
USbNdjDDUzTvxkipnaWZjnpn/Nrl81Woq5oLmScRBNkBoJJyd3QTEyRLFIlC0fVK
aKsWsXv14dpyujF93CrNbSYFveEy/6yjjFPwKFS4kL1Q26YUZ/Stf+hrVCXNFSGy
tS1V9XIvGxfY7hZKRCGTXNkDTBNg6IHQahGo1s3SosdWqgeVny9CunZ9GgPQOLZJ
UNroFcCJHwMUt6l1pDfxroeQESljYLmBL/x3N3CViTS61ODLlfWwb48qePqeDGGA
3/v6/UCxkZJUZUES2tvE/aM7qtAFENk+23+yID8bM/25Ch8LOOCHlfjXy4uWokDd
QWMs8mtyfS1Vd0/4Gyq/41bmA6S7SYd5SIjOFIcwoFzpluJ4SOaP6094aK/77ujz
DmevkAuTBXqq9RmX8AYUcFvvQsoyw2eX2gTeXDBfDuIDlOlIsl1w2k6yMEHOStwO
IT7Y3pUugGvok2p4eDMkE75AQ00y8J+Agdlgjbrb6b3sJNCTDCNO6uWNdlqcxSAu
S7DsHvfiGvEqIia+CIC4o63tp3YLqL9+wHSfTnhJ8+0uqtix5KEqUbCk0Olg7Fq8
rl6yQmgwM6gj9EeFAupHVJz82oFjwg4UXnWqysIf7SRq9oeWwYa4jEdzCifiBW7Z
60ukR1ZY591j5btoSW2bOQjWQT4ogkke3OeVbxljIJRnBaqT12N84tssbQMYCu09
D3MzYSmNlkRLya5slWmZ2u0kcWG4Q88PKbgQgQQKad0FEvcVcz5Si7cxR5ClJUTN
SulC/ifGIhuRV/nBtYNFj5NTagSfpkIj9IuIKjHWvwxZ6XChlghh0yZ4XZ9dsHj/
9+t4aTe0Q8crzJQdvAWe/EJiZts+mrunojTJ+xhdbMR2sKxrSKugWigZUgDgai5k
HPOj/RNZgHApyyIOleMYWvsOBV1EPd70aezWLveaQe8XiahJ0L5m72SM2OwZDVoe
srFsO40gMy6ycG4Z3FGy2VjRxYKgqUlCtWNUKePBXySv03g1itlOf3KQ1f05WSlo
WBHxNZqAJwGQS1VWFiIEz5LqtVsJj2SnYFKOML/ZPTnOd7tAepL7CWy7eAOQBeNu
S/VgWn1EsjgfkdpkwP81bB1N4fnjXP9nmLScP6JKCHfPgIw1Dtg7u/vRH0Eg0FzI
poVov/lE9b+oT/jcY3LZaAvCj+wNefMWe1Z/SKvCB3xSsM0TZcQJuyE9I8LWZqq9
4lQt41Cf+G7d70VEOnYyeQ3EzPDV0mJKis0PWyV+iR4U3nYA5zhyg9mlZP9KVfNZ
rxP2owXw30TuJiGWBy0FbFsQcOSDaG2Nw9AcHs6vhvmI9wnPcO5gVe9ch6W/VEnt
bO+lEg/Uiv0tj85/pT0cDPZpZwgh7xEAJ8p/FVCDtZrd7ooXOGE6IjoC+EploHX4
R9S4ZFoZr/5Hnj7LI1tYJRzebjqhtlw7TquV8dAUvEA3eDRWMmgq45tEbbwg0Nd2
hhD/tuAA2ic0xABsPCoD0mWiuias/WtjHIFKFHhQ2+hC2UW/tk6SYDrsIR0u2me6
uH7QvawXWQyKZV+bXcPvJPuqVvoGodpRBzYt1jTiLQ63sScP+mdfk7Tw1B/5P+GU
8ejqETTb1XkhLD5VUX0CVtG+kAjtya8s58BJIaT/fIaTHvfCdcmHkTPfCCBl6Czp
Rq6DQrfjP/Ve9PX0C6efGA2lK88SIyikHR5PW7ZvPNTWatpqW5pQ+3BaDdj2LSOi
RmShKR1dzf93TiYdSy8sJB4T2usH/+HIB3Fk9AEWgDoOMXsvVlLzb2HPdTUTwEXb
lAzcgccIgC/RyoAf69yCChF0MFWDyUjMHQAauhvYN43J82NuI6UJRdR/JHCpgF4R
0pCTylX2AJ0chQgnuMTLxSXye5TyzA01oUruZCHr/B4blWLZyyVYTxareHpBbHPK
HbfGcXlraRZgHCcdk2kOxBdCXW9xbfkryslsnjoSEOWw/tEhA48OSFiT/LIo+Jpi
8xSKWR6gNFao/2FQTczObuz8O9KlsVe8QU6n0H8zF+3p+AIsGnZjy0J2n9gx2Fhz
MOjWV0AEsKpwb+ypTz7eOayZz9+qSHYn5T0Wwd7ZCsTGUykucCFymi6Rw2L9QSbO
cX6swMWZvfJEYlLK4Xrl/Z4NBhbjMvsWjVAasjGwGWXsCQe7gIpens4dqVgts4Y2
K2P2wLsINT5rid7CUFYdVV8YAdTOp2gSOzf0AP4H5SeP/PZbgahVqtBMlW4o1qOF
m0NqCgTEzqwzBfSDQuobsPW/REcXM9rB628DPoDzlImVRPbidgPAkrzT+bz4KjI6
pbeleNHC9l7hG9Y/Re+BmgsJYan4og3ho75iFPUuHyLEr2L8gEadd9G+LuU7w3Ss
X85kZxCZOwdIb+c2gmC9UGsUhA2Bd4x9EDjL6WXVqyTkYrOfIw5XsPw9IRQa/epe
w6i4EmlSsDQGANM7VS4qZeJ4S8xTwLyKtx4gamrn4FpdmQCKfACJ7JYyuuRXNera
CYzB99NEV+1FsOC0tSQqUjdLNFvEs+FX2T4RqJ6Sgih7rLvBfm3uYXg2OwctfL63
qSZQFoBAy8bBJu3P8JNZQwG8FvEalDa+d6LAJHNTQ8Mp+iIQJGbTXGNYnaMkIPWI
mzMmB/MtkTITosbI7245mmrzuYgGNn0WJHl7fD49hMLXgiHFx9zRl/UZ9niKEmjr
yAkK7caDEOwdfIJr5TIyTP04VD7T31Z3ZvU6Hrjif3r7JQA27qY5JNP2z3Bbt7Tc
3E+rfwjQoMEKl4wSv/weVXUQSClGs2WolZ3EhwxBFFtwU1irgRdYEfFHg385Y/Ga
aP1jVOY7pvHLuwf+/Pw4HHnbHYWmLJNI9iYOWXkQa3tjr8jurTnBjsj9yVBtYS3E
GfkuUaKOoyTN1yjPM/WqGq8I2/GMRmEV7zUK2+19NZjDX+45Wnm1NbZp8zA95W5I
jOqDEVQVW30w93frSwVrkjMWmvkoO8SWpVhZ5vumWXDQ8NwRyCP6UoHYvIUfmy9Y
nHro0a1YAK2UkrS2tAvEoOEOBYD+cfhAQPRJ8LYinji5tRV7efdgk324ChEYPz6T
b500NSefzDmhA/hMhZtp77/xPsys8O0gkqID92aQDzeVRVZF/P20ki/QCpD8X7Zm
pKT2f08gVD/wUyjJalGVGjhBPiwetum33Ks6phdxJ4CpYJVFCgiZG1OHwMwILUTA
vpztyKQWnX2T83N02UJbuiQ2P+o6/awSgri8Gru6QQDE+kPA0gGhX//Qt/6gMbkD
jQtK9PO6Hvv1c+q9S24nmYDDf0SdTrmWF4MCTrA55Zz0LiAFdUTHKh4KE9dFfbpJ
MLCUjSOpWLEUNAoFAJ/5P/z7IzJvVW6Vzx8FJ2mFqz2HAwuGRjhOn+0iHAE3joBD
hoABL4KxkVJw9p5u/z7LXg4K5hwvJqP/2SH8VN+UkZ08MJXXQWM50Qo0OOvAKVje
a0zJmHmwVfVk6bzLcvVQhJgfL0bd94WvfkIX/RYxL+2DFvDEU8raGyz5gA/dpdrF
6slSlzekvmh/yh3+bkT9GcS9FuMKLcZh5+nBUI18BUuqqDjcfQkOTiTrwKmV7+Hl
aqeIln7QxK5Il91Xf3ESIGbrCqscK1dDu5KOK0T71ocltcLNt890EK7yBRoVF2kv
uS5+V5odRznruj9q8pEPpXUlfSK5TRnWVgwY8/bLHutCOqkVXLwxeCB8Ye6Omff8
Vm13f/2XljbjmEo/OsKJ/xvv+0X8kaNWhPfaZ53yuUE057plP0oTcFD1O5Q2KstZ
bgDLoFH4T64PCFro6k9KhoMNBJYtBhcRblggLgOfNTguIWh1gxf8ZKZSs3YJnPw/
xbhXs/HGy3DkR16IkzS9R+I3XymV1rLxDNGevhELx2GpaZmPAl8bOWeS4yFRgd5q
jgw+F0Drb+vZjGGL06oh4Km5/IpPYmYm0DPHMH3AqCsNofeVoAKLoWSnXVcUrVc1
/udlUNC2GHzpVzalRb25njOYCsAAHhgniSv7HRN08WzxePJAbA97WHDqG5V7YmeQ
qRKdwEuq5Vedyg6i/eeFSCvI4+LH3mV/9kvYXceb1WYlaePAm/VRHkLp6IYMSeeS
jZcdRTABWt9txbcBiAcONQm94rHUrebXzNVAHgwmrEd9FAjQjW4V+2U9IwBTGjaQ
hI3b8PtYDlHRkTb9/fxjbnPCm2i6wu1m3n07haEr43TTi4/vUcW/AWZeiehf3UaO
89CRKB9W6JYzu/bQRnjAjzhBDM82/NtuoKeUJwaHLmo10iM6zCaC9pSlYZy+uv3O
dwi3E/shQpvAgTyrPjY6wuN77fUeXYH1u3r+szD6JsdCi03Cfb4mDC8cHrQ3xbNq
CASDMhxk/hu648hY+rwPN+LxWVG0aRILjooKOK/cRxJRcxZXrLZ6PvXT9PIbvtEI
2YyLvPrpU3y6zDJ52UN3DdCtwe5Z4rYZwvO/+/cFO2CW4nsV1XO30Jh91mqjMXsn
mN+X58H6uCaexOdseE/5AY+I+FcLjUXkNEG8294T7LqMyeqEF1/i1YY4IkYKm7Tz
P8qx+eaxe/zHNtmkyG/RU6lGpTNAW151TYeVfrqfqvyKHy/SVRBGJVgacztQCWxW
LvlO7asES/ILxv6Y/ACb2jy3zGigHOkTQQcwHe9VXcvU03LwKff1Y88Wl14i4ULG
YElv0vRsw6+aLa5TfMbKl7DpEKJiChZ9r2Ixf0B4Rn04KGMWNWK8EtqNY30oW/Uf
V+S9Kc6zfciZ339fAU0L45V7zie/xW+ck60yMDz4E7r6eYmuE8H7amyhkjC6Ht+L
DkbBwDulfPYAOiVwL0qFxfs6KwiwE60m6Haj/xDT19hgTiIMXzTFQPztNBMwRGK/
CzdwVDWKK6hkI50qn+9mzM7T/545B8nIexLDM0c2dGhTZN/QADu/FB/6L09ERpW9
cSczj2f57wUm2V8pox9I5JkEDI0W5G8Ta7gs0asFln5MK8ebowvdvD7fstG2NzPD
l5maugVr+nfPALQUwrrmkMwqNLUd3ZvmIBROjeHpvr3fAiZJnMH5+NZoSIKrZ8r4
I0Nr7UmVaUCi/2yMcdRfkpcsDU6ej9FxUZng78iMLc3iYA/8SEwNbrEyu0olwMak
n1Io06wlF7JOBLEpLc7EQ7R4rL2eOjvKdcgbCN3w+Sl6V6PTh2D9/KyniJDRdzF5
KKLoZZ0hlM/jsoIMv/CXbicomKO4fzRU/GskkQGOyczHhPHmFE18KnLAifuFLpox
jzH/yCWRjlwDrMSHdqSB1aO7YfRll1E1RD+jC2HVUUUKHWpLQeIDJV6ez97Zsbo6
Jh0iY7/uYdh/QCES2Ao1206INvGQDXf4nHjiyWjSJ8H7on3kBLGfC0mgttWzMEaT
hv6XiI8W1BJ59W1UUH0iFKXTnA2NyNHH9aXyu4jSofZI8qiPt1XBJ16nWKMm+5wr
9Rc/MH+m651Qq0G28jEPcBf9lE+LDJNWN4EnB8yixPB1i9oXJj77tbjxWT33AByc
eZ0TuBbc8wgaZRiuTwrdu8rK7hKjGZj/BA5bPBjrCtx3j3QYjk/VjK60AWretmqr
arcel4Go+rwTy1Ud26kqs88mYmo8B7JHDrvA9n1SXqcbxXaiPcf+eSFJwxMLBXNz
3pCI8BsK+rRB6nPnh2ljdk4yW9L1yO7yCG1wodmBxCN/6uxzRO/q3gFQtg3q2wlv
UOrtLsHnZI6GR1jsE46NW04thTunkLXNOzOKJX5gdssa25LCVvOSKznVHlYulRIT
kXGzryFqgIW1PdWYlGy1sztcXOTxU7qT8nJXN02p2hDFErMm/DLXRCSpooCWbef6
RLuvVWU8ZfVeQm/5xSLEyYKWnAsSFoiqjr8t5Uuwdffx+8h7euNRW9dbOr4IfaT3
eemwnWpQUQ8WRXCyR4Jg/apSIO+FdWNDeVQzoNrBXcXL+8yQSuFUi+JZN2rk06pO
3lz9z+woMr9/WxV9sTysynFdKgxyqjPFHoWwUz6hJfccLDta3T/DUL3uxQwRU5wp
rfjrqvxhlLqtZW/ug9wQ/jYyFc6860/erZVIl2DLhrGR56IBjLwZvz3WipHftMMO
9BvouwaGtTtNZkBKy+QWSdZR3h+o1eOdvqDl6NRVlPyo+HnHyW0XNbfU8cHZl8CO
XjmIJNm8hIVYIb4w/aBeOZJESWOwWNG+Wk3xIwzDpINHc4jgsANVQdAZ3PIpTeny
zW6w3KL7I+qD2S1hIgTt2NgCSWwToHd+1vyQd0uxpQ2q4P8CwvdxLxL8fpFY8zsq
3evY1x/QA48RzXCjf+IExjV+IJpAhc2zah0nWuVXN88j7cdDRgLFEI7Q/3QGpbM+
ZskKCVld/GGc8OW4Ln/Brttt0JJI3fmBcuj0EsQ4CSXUv3rigX1kNY6U8Y6yTmT/
7ypf36KeoK8hGSHA6+3uLalMU5YmA2l0yjIc0+KJprm/1+EkEDLxRsuvQf433dfx
G9UD23Ayyxd/whZBCVhoBUj7DFl+kXeBghYsjuQNyxTebn7vdy7xrlINoSyKOuD9
ilm66qc1LpgsR126A51dl7UGG3Suqjim0tGViKYgOEdXoTusAE/r7/8xHCo0W91c
0uP4jd2He7/G60Yd1qkenxcT9mpBWWQSwaqTARoamDIT11BP571CxwyWQeeRbh48
DnpThY5SwyJ3prtL4FcP6DrbXvoITNTdJk+MoQgnoPodtUTo3wkzWCwULm4cOzNb
zYxCo56Ws1Niq8PHHexlcjzYyJorSvhxZTu80HmiPpV2MH/JaJiF9Yg6JftcMoJG
3JDKn06+tNeEH2AZBP7DHhYRtQmn5oXnkMyqmIkROL/1zeEW6jpiFZVjuePXcE6n
JG/HtNh8L7q//W8RjsJlDdsIszkDQELUaty08njJ27WfHMXByFjA/cntI9C1wSRn
IHeRxSA4vkbcsbUFWLdogR6nyKOqvRdUDqGRZtwF+sMAD+2pvGX7+kMEw+YHNeys
idysctZwo8MN/FCGp6wtgjlqH74Me5+hYvMibLK1c5n8C9fF8hnDpdfQro/caWAn
FhF7kHplpw0DqFGjmMxnxc6KgNlUTTQ8a9Gmx4mAajI96KVsQLtO2Hc1Y3G4tvpa
XydhhbZ6cW3AkHOnWnsmI0rrs64e4B+tos4nxinzm8jeTZltEM2C82AgMDNnaSn3
ATP6jxlfDfrGLNTrFmeTV9eo0znTZJesNlFgdLe5MxUeup26fQF8y4u8CSihT1M5
DAVav5bsHVFXgR/7cctIav9eatXs05FbxoK4izBIVf8TW/TWgpk1eCvcieJqxEHH
XCtoSY1iuMss3Z1JTxFVSfEDRUKl9aKvfxsl9yJreEIu+YFzmzpJ9IixyjdWM5Vy
jJmwMk7LdhVyc4ydh79MaqPRHLDZeoCyAjQZ4Qafa81IoySko8ysEUQBlfPnIyIn
dL4Xv6sZlAiSVD+o+EjcyYZMXwwqEkoZWZB4XD9+YNoF3N/vkYy4t53+u3t7Smwf
CQwhCuN6QCV0nsmTnZuyqrVMJCwSAFBujZ8/SPmIOSsXdrJg+/e+5V8ObpPEiNMR
SbBM3lEZGnPEQRdSoVTeHwKufFnqC/w4tzrDhnT0YQp9X/4h+IyLKvg+L1YCV5WA
q6TFh4Opyt1lXwILgfYdafwVt4sILseNAZLOMcNN35Dfj3rBKdCeDQMzcxGPmioM
x7XdONhddpaCQ3Gb7OfCa0fj5ywJ9LmlW6wvdpNIHpzQZMhIfAWjTp7WMlPKo53O
p6ug/A3YH8CvD5t5nKlBpVIA0DYpUl7K9hD/RGrmonJi73jdWqIRIrXFhzWoRQtT
6FeU8S9FHPkYp0HhdEAdfzcf1WP8kMXKv4xrYZ/HjH6Ce4rPwH4eaJPqltI0Z7HK
S0Gyu6s8yzoin0uaNQZa6wqiT8D7Nxt4nQYLYb2JJWozYIIQIvuy+aa+WjS84aBk
7bVn0Vx9ZtffNEbrdoExo2YlWijE3OzAt/ZQAcd29a+186WmPPmL4oI0x6DDkGS+
uZ6O9DLQOXwtb7HLIyyxonNsqNQYg4C1GroM1ZL5clvVGhDP0+Ud2uhIS8SZhkxm
yAsv9apX5U/irQhKeo7owkKgL1g7N2u0H7wdU7Mjo/SWhVOLI4UKoF4db3R+fYPl
q4Cp4zFth+JikW16QUbO78p+noMnahhoMQCJqwePsjX6jS6/iZaMJpjG4AHSn22x
DxWBujBo27LEXF6ittrIk1hqGMJyEyyAs/MJi0G5rX44WCTeqkGsAMu6AR36x6rC
X+eIdd9FDy8t8/GheS+wa+tXjJvJDJxFAaBtfrjXNEFHMp3+Gzwh6xFPp64/f6Hs
jgCvQUxO4GbAF88UQcD177iCO9UxTCpOx7dX5JtHVGbNSL2oExOkaj01BtRRk1G1
PGTiUwIRMmw6q2zobP1+bknqWa6TPl4veERUeyzqsISdqA6IOORfGUPmGCgIsMCT
fNglHJ700YJwyfoYC6UHQCU+xjHW9aZWKTdo4Ua9x50eFAwWU7+rGX77YGzGFXAn
8Sp7L5FGBSskSnvlbRspgpAmxTSuLPmbv2xqZDQDNB0CQwCrwzhW/QPhbnPY9+qB
rkvc9Jhn6imigu7A/zQtubs4FQQ2C54wUv7EaYDBdvyISZGD1W89FucHgT8heHD6
u5RWPrR4tn4bixcihRqKEdeMCfnfwhBz6LJ8Z2W+Q6QAhxOTAhQv2ljZph5AGTeH
nvNsbVrNxsBJPGqZaPIF9Io5ErhjIG3bVN5aMNHoqFwvAzeyDAPwS9M7MDhv7PST
PFdht9RG7i2ykUvJ1eJNvrxoT1zHNrvVN1C8+MaCdJQghc2WyWQZh3epNQ1tjiqF
lU+/q9FyxN7zh6/c0QnXgctpGxfkZ8I6VZtxIVS1MDPjqvPTAXNh6TYtIE9ZpubU
J+Ulz+WC15DpX+eZomc34WA72qQfbJiLPf8FqAsVqUJMw/722xhktRqEKP8e96IF
7tdmhCTJ6ERPiFg+u3tmnb/7NL1DiY+0e0FCgOFkWTY+aEBEmZ9oMUr4D3t7OP34
v/lVfbj1dlLumui98EONSI536iO3J2yIfmOBRFsgqUX4oEWx0RAQ16H4bLjBbQNI
vf/IIkIyum/ZqPOlaokwq98Cb9EUQgr0GvaV/RWua6HomtykFqNGIAxuweboCEt7
hFy+Yl+i8bu6T2NLVSps2Og6sWKhczHg4sABczJgxtd4EOE+ymSG9qCZxLeDvZ9c
37i4T64zGCyfp5v4NKnaEmIf41CNhXvlT9wt95vn6q0aCICxwzQXksogJmBiNKbX
18Kh9k0eFE5vpDkKEHZavAYOZAclZZ8/WL6ICX3Ml7bE4w0q0VxfT4f+t70Swdo5
VYKsLchBRSHO5lSj3iXN4StelxvmJaunnWp6U6b6iLnACZVWT7rOK5cay05WO78I
4dNWafoO8eLKwsADm7n9YgqJ3+Z6WdjMxGvShTZxP0Cy4C0GAVfix8N+EOQa5McY
vghsE/JrrilmPf+dZoRfsmB2o+V0JbB0KlHE4KjCCeUJI/H1t0qdwSPNw0nalfUT
rGAaG1K1ZJYiwrwR3oXyuxht4H3aD5Dz/jkL6l6l9nLwu9s4ZQMfTidDKg0yPiEv
lB/SFlOqZ4CCRmdVjYvpmC3YoPrqq7ub3MrGKwGULCPrKFqWN+iq+JrTOTt4Uu3v
KeTYyNlsTQuVtYb4HZwsjQKsBGTkMRJ24NZKv+KxdXD93/dY7UjmnX0Th/Gwaj+M
IMRFrAQNnVJDLATc0W56zSSKPInK49mVKHCMVnGIL0AD4Ody6OXzJWfIL4uoWEMB
G6wwtvSXERLAGK4YMn/BHewFrEjPQGtwZc+Y3XUTM5Iuu7CCqy2XwvNq23XxMOEa
Q/OIo2jmwp8HlHhPB4/TXxQyy8WoabuXMg+gBVdaKRsUM9mrWPOsJ/zqUUXj/yLE
Cbk2Vw+XWrmLqwxl1EBxVavSQtFaSJPodPlkUT1QtQwT9r4ZoJs+Ozd1TE86txXj
MJgdlRbE2U+8n73sIuc+0wjljA15Y4I00EsbwMmBpbcOyH5RaCwoRdO+nyY6f9eK
yKkY+1R8iGHYU0zm0AQVLcN6rr0twgUH7Nzmac1gzduiLv9/yXYCXFL3TaNONN9G
D9Bzp3L2ZPTQ3jyRQM3sCA9h0Z1s4mOAUtE0CSturxkwN02Wv87u18oIlbYHnGhy
+yObQtHN3VshGOUBznkCPUSGtC41Jyq4NtHSb5E7zStqJcW3kE6CHmNJxONRvJ0w
tpXJv3OCMTBo1s3uoAFBf5rxZ92Mb+lDkMMhGxXIYXuloM45RQNAZg+f7yBt/HAt
r8KCijR7JKAOzUv6EpYesZkElwaWTgjvnbuT8WqPKKU1qiAGDgMxsd1CAHvMkWuj
iPXCA2j4aqR7CGklW5YWJt1bUhveqyI9lFBn2OKiRAlDAUO5E//g8DTP96ADri4l
PBk1NxsJwiUH3QlIdRtfThEWi41IvFjM0Om7v2+ShbBMm6M5cbTgb/8Ky89L688L
iBvsRLKbCUhwDH5HgvwDollb0YRAGpEyi40iStrHcuEL/PnLPKgZTwZl0UvyJX6K
/7IqeJPpqjA7kBSJh6Z1aueqna+vHDfdsxmM1PCrAcE9E+HlHuDXLIB8pHFMRXHj
u1O1k70NbyjLYa749VOHuoZherSEvKElASSh7MQYO1k8jQhNjlkyLutEfD6g51XL
/YYDoxpw2XpepsjoBPkHMRSX1ly7id1E2Cq/4uAWg7z3R+abGDPkrwMJho1yNFaE
orFMB5hQM7b8azVIRawu711iSvNGL9r1Vua/Fsba9B5CN6eOIV0Cnn4SgkLWobb6
65qC/uNXRYxARypfyfPqrKm9mgswuFcf+n4doNz9J6NpZIGT1/4aBMLvonMyJH75
Z4IyVYIkjnVKtKHojUctBRpZhzZXFIrc0+3spV2RcIhedfcofC4+nMBsmhcBuEy7
5nU5vN4HgR2NmOmfwg6bxJaf4FB7faYgoZBnmiSsIcIiJ3yfmTErsAOE9jz0S283
cKL7GVu7y9eFyYaO01PhNtZ6oSFCUjCIJjm0YVRGndMAepeyyCyNQEyFLLkr6w/W
prKpTdLHRI3PSFMEkXXO7S/fqmv5UxhTn3VT8BXhFg9xTHo8BASeUIHN2/ab0Owv
7RXKC3VPc6UbIfxMY1X5IkqLlXpctlAZIZWj4yT9sFn4wgGQA3AuBnSd9PUEAS5l
L/3TQrCpu6iXy+uaV1a2xU6/6jTLLz1U5IYg9C7Syq+DteBgL3++c322sdwlJEH7
STLVYyL4g8n+H6WaTdM4qCr9x2iiH+QtvGCoygswUL2Ttbrz8iWc0ugoyZoe3Dyo
QYQXfXE03bQJ/jDvPEG7uIuRNc20h6pZvupjcFfQIvkLM5OzCQaY1yh+XGh3bWp1
PiGV1+qdkwxIjuOucd67grMQVbk8Nj2fCKw/H2vq+k19J4rayczOkD9YAwOHh1KI
gvXNYhqZD99mvoiLvYTBA66W5gEC1s4KNnT5QxXIJ/kUHpyKZsmsLDkDi7EfoP6U
dWusFQi/pIKusv5Rh5GnJGPM6IuEHNUMRaaTSp/e1lFssKCrgshYQhZ5Sq9JmQ52
CGR7RpZYhcdzC6d29lgaSspG4f3raVYSqtus4841fLUf12yu+zqSRa+xDrr+N/x2
YWElwiFrX4Bz3ipVope4E+tS+HTksnTpEmD1+87aN7JsLDom76g/1MH17mbHJ26h
ijK5UNprm/0nP0+CTs6k0CHtBmZ0nagMS99uZVtjjvsRAiIDqzLAdbe1qsPH0lRR
Hyo2k5/p5mUFhlR24KXSQNcjOEA/lfUJoePHhrdRMAURs8kQc7TpUdm2y1Rc/vqQ
8OlOaDpw8ltRueE7v7gEJ4x4qUCu7GU51+6iK8hf5BSZKZoby9C/LUE7XwSUVsjH
3LFQKXeFNq/uei2CN6g+8xr/LC/y9THAJf/NGZTWC8mb8/b0GxhU0bFPsfweOoKU
WD8OzWKhR3hKqkO2kS8KooKsNSOH9sbEhgJN5zH0JYlyPAvu1SKO8g6gr4Rurd7d
9ucS9nyHqGTeF8VmNIOnaH5B86frcYN7iKr1bHdddPaHrQhWjQowsuxYxymkE3SU
jUjuheQr5WF7jORDPn2EshnzLwYavVjd89ZZQWYE7tX8mapy3F2AYLoOgDIg6EFI
Z75pcw/KUTxWawm/OsScKy4E+X1N6nUcOc3cUmnIRK8HK2Bhz7MSWutvOIlGP1kF
+TussLCzdDtaQM7Ev1/rfXajM07ihom7Eg+gr8yL7DyRpPTdzh8UEWv76sFee8bi
DyDIbdVY7SJYtaYylXnWh//qpfwdY7JVuoKOJzGSTJO3I9fRfJG81UdeJo0Bto2o
zgx+js6JTjvuuPWxajmYGb0PSE68LE/qOh3JIVYWBPQ3KvKq76eWWtBxoi0zjxQO
ERNn1Qfszl+fI8ZU/uKg6Poqx8zAMrqQvS51EQDG+C1BPKrUO5MZQXKYbcW0Pf71
CmSMFbMJQgEYnbfPcy6wkcNx8ewJLFYzogz6Yz8ZJkaUjg5QUa+OMq+Fe2eX8P1U
aGa2RrfE7TDP+bEqkmWXSJFymo8HjA1M9tk2lRRwgsY+GICl1G9oAL3Beh7LppGX
S9r2nHEEacSYSlVCFBYhXKgrvQTVDYu4eFaU9B8enelNMmJvRbZvTvqB1K0qjWVK
/gwKd4zWVNTH3p8V3A4jDFD+shCNfSqn+/VRxJsAYdPqA8UTTgLmifjs2F/CX9jR
LeYfpYmy+B5lBdfwyBt0We1SdbuVapmasz+HQPIoUhCPd8qfDYqVeb5dupygLHho
r1G+oC1/E9q1cfeY+ligQfs+WVZJesyuSZ0U5x5dS9zAiUNBoV8Sf+/WoPN2sEzn
NDtrnMjblwYPrdpLA0rAicsu6fYp2TFvznZzAb648pUltks/8K7iIgmJNi7nRWUA
PGZF5zvK5HHWjakTN6K89K7CVNzFXtHGsgAic3oeNW199pbDhrW6teHgFUvYU28B
MKHL1N3RCNVDasexCIdH6ghd0scvGK2HQmiMUHfPdLRwuqkw00q8SzTNLcDzL77w
KFdn1U+O92aj113NG+Kdc2+l2TJQVCFqeazwFaLTV+6tVlVD1FAJjzVN6kSKaSXO
G24E7wzprWFCOMiZoWTEKSEvz6Qh24WBR0IwVqRzmKFu09lEdJfDVYJGukk5KbIG
zHtKdgZ41Pe7CBoJfmuqMGuL3DvFf5OcBNzBoBERDMCIWAZmiIPqf7tnyJsKUqri
EkTY5ygVgv/5/tdghsbKgAdZBAu47O8btvOu1rvCmmYLK32SkTid709G740Bc7nR
s5++1reBZh/Qfwwq588v5D8zNSrgWzXWjYqUPEpud19oSU45MGV3ZndnmxZDwDxA
7t6c93yZhDgOL4HWV9ZsXcnfqHUb5F5sbUkFH92JYk7EsTNTZ25WJHzh5SrXgJAZ
rrjj+x9hwNUNtZO5smU3zskEQl1m70cEbRnuviLNGmvQV6CowTLciKKa2oZa8mVx
74trmRex53kXzKjA0dXNlDmd6Rbe1nJXUNmtjaKWEC7yoQPjvfUubPLCoI2rK5Mn
9YnYqJK6LK00+7XlZLM5+/3o6ECHaW0eeNWFjIN0yQPHRM7Z1cS8d1dN8HQ21/SA
K0R4AmTvtL3722O4qohsBvto4u+6sW8MfRjV12eStxZ+/x5dWIeOrvZbj41e8qoG
o+PQl4rdg315VOTemIsmfgkoy83UcVjijZP1vr1lVsqz8+tbHWKtaIApUqGGE1pN
pqWjAUzhSl96t6pgF9u3ynINGTdqqOql+Dke+OGmS0GNaS9LC6RGEWttrxrVeGFy
Ry66EZxI/XvkbpMLVlDRfLhiLmLiXUsIu20zoo4489RsXdAvkP0V7U07F22JAoXC
slteKg/2mTuKdNVhhN216mTsl8L5ESLrX88c1Lopmwly6Mg+zHjKC7QvFKzWSv9u
SviDjWTMvxo82yHPSrMvi5wf1k17hCm5a/CV4a2PdVdte5+TxBa5yrNF1SrpmwQ7
jQlq1pdxGY4ttTucFo++HKra9kfNr+uaW5w6zoqsSX3/v1Qlfb8hPnFOi/dIpJdI
A2R3NEtrTalyX3xQ5B01mW1kneC0Cx3ffuAs2kVcGs/3BE1QxzETwyLp0Li2vxZa
eOV9L0h7y6RjLZhKQeazyjhzgegb3BK+3u+Ksr5R2GALtDQn49pbLQxzr67NGmty
jGFYuQyk7nzwydZLtmmLPu60VD41iNpw+1u9ZqFNy0keXelwnI+6SWdCpF9WmT4I
mkqanVRSKdGAAs3dOibV4URhOVGz4r5eDyCZx7di6yvLKtq0Oq3GNanv5G8LAcce
rZHfAI9ur40hukJaIgmtyajLQGREULKnb0E8z/B7NVwl62gJi6if2x7WDCNfKxUi
enKCnjdvxzeOVLfqWXt+BqxtqlAlTwINhQHt9biBXJMCirUAbm+yTIIPV3ehkc7R
0xgjfhOAD97Myr4SQh9QrJwh7cAlyP1ReTF9ZGtlNnqkDEneyW4PaofPewTo9zsi
hHUdU7NMxL/sjz+gA24TGtPfhYQTGZm9VeYlM387ETei6Zq1ea6LRrtoRdO7s3/5
GnK0XLZQGj9whsGGO/g4uj/YxeNYOFuKuFSt74GBVZLzD1lPDL5E4AZIHEm7UY2l
6zRoqdKQ18HkduiOn9C8fgAsgwjmgdok8rSoKidmL7YK1LTMW4DnOGmU+v7tkAvV
ZxFVsdwoLC5OyV6wuksP4vwsC0DT5Df8X2VYRFJ77s6ARp32DO0Rc2J1DY67RogA
xka+vGhSlGD8sMvLGN4tppij+v1EHdviCMtnmAEKOYKBFV2s86YBiyCtrrFspIGW
hqPNRS97XRWC5Sn9rZrdFuwh48tcqn2TgCpzrnfO8RJ9hCA1fqOCw96fBCLpTGza
9a/CcGzGN0wzUAFtAR7nIll8o1RwQIJavD8bzqvip2eWP6SHgA2s9kovM8irGnDC
Nlbfgu8JbrtBJ3gTFPXr6SL9a8w7CepEr8GuAU+wtB6gSklXOO6XKie6kEIJIiPt
UsJubBmlBnkv4cAWAnpvt7RbBbPSE4nFS2WoEA+QKGMswh9Z+yONBmaaA4Co6sBr
6Ra10avRP7NfIu2cBwybx2TPiuObpJiN0bIY7aZCFd2ZMdqp/cace/r/XmW/HtcS
NjoHXHyLmI57+9Ib03GYtxw/FC0vl9wMX8KDtMJHYR5QzRb2LgYJudfXaoG5GdEd
dNTyeTLaZYdmYDRkixWTIecl0mo0d5yMhk26N2v+ZpTjCyXEg2pP3kL/tY+Xlzox
1XYllyprjmYDMbjaVpj9HNXKNHoToLDgFXF0/5RXpsp2w1NznJb5/0xfke5F6tTd
m2wZsDd+1POEifx3m/21cVNa9LJACZQ7W7wJB22Py052xMgJcxg6eSw/eq7ADBpI
cFU4XM4LBlX34gut5evJbtUkm9kG+e7ak9ou8FCwPiAHtTqWzhsP7nMVb+gC/ciX
hEmnew66w3xlOz76HJM/pgKyzMUUuKeQfqBER8aUC16jB2yIzBhcMeiHWOR1QLj+
fiR8yjfAq8RC33uEP2GqXAx7q0VH+L+rpi87FfpfYdZEec2Y1GX5Q1BvgVC57zi5
ZB4bwW4aFOFQS8KY7G4FFmuJ92Ftw9UPJGA4JxWPybMEXdyBLRYDgPlCE7Wup5yv
Qq/A1wPY/AbH0kFyy/D81TBjlP/a97JMGiZEQ863K+cTJap6ffgjsCxrgc0P9IaA
c/Bc+JLzrYLbekZHl3pFbCSdvbqDhVdUD2ehlkwR8i5US9R9nPbE/he40E25l15S
KaoRzmv5XbAjLQqYT6rGwGfIOcxk/di9psNUl68PMKp/CCLBq9IH82gqULuI1DQh
3yJdy/1p0133um0r6bL1hRBom2vVmcsAg4uXLYcTM8wpY2w61mfqz2zYWGWUMbhD
j1TxbrQa3VlgXl99Fam4lLGgAL9s1QbTg4GJqkNPNCJuHTmrnUYj/Fj3zgRHQq2a
0dx3FYCIYgHUoO0y+wzI+/b3MQRPYmY3PDQibAEcCcNOVye8ZuBSg/R5XYZAHVgb
R5KIwHcemrl2wDZJKeEQrlhWtJKGSK6FCP5vE+VEdaSKF3CbwpBaz16Zqw4i7k16
vp8ZHru+7ClAGeMzyQKqep3po0WXv8Ksi9ky8o1TkPT6x/hHFEke5ri/FVDZs9O3
FPYn8kUANzzLB4qo5MvBwg4Vht4AdSxNvn8MuOwEv2ETG8sc7azhux+/h2Ec1Cf0
6q5YewMSoHOVVEUXQqZTYb6xO/GptkmEHDF6Hpp4+cX9OOz5H7wEsvGiKb6w09Fx
IDZ60Xn4Z+/DJRYEMdjHwWsmWwBbziGK1DSlv2wodX2ae6abemq4SxN/aVlLamcx
1N5xK5D+BXOVwEZK1lYlOiS5MD3AT6vXdhoEn6jDDHlKB8v6xUVoO9SNO6YGvqtT
TEgG/g+P/XYRleTjBSVsTOfFs17r01NwOwU52xaxpcL9LXkZQVEGdaVPdE8lK+MP
SfLMz1zlLmsZsqjfZSCZIrTnjJl/HDCO7VrNTRPpH/3eOe0TXW4KYIL60LilAq6X
Qutljeqd5kNHVIzq4qgTjZoHgPtGRgsc7ZIikohXYZng99WzyB6NlMzdBq9SqRmj
eDdabg3J+9cjihD7Pqd2cbTrHODcvBcNliiq34MqnLC1vRl5DnYQMCGTW6IUzw+3
O9EDCrWdu5a394AhRHpjLB/7414+QCR7mCXwM8vsWe0mpbFJgBcg83lueqshgEty
7DX+AU7N/tFPUGkYcd3eb+lWo2SPKdn17sHhS0MzUluEfBDDjytepDM5cEBOvGJ1
7M+BoyvH0muR+6DDBzKt9bKWZsHxEettJES47w3iC87Dz315an9u/HiHBlwMuBAR
/nyRIwf4Rn6jRkRIX2JamhpWp5tBMiLXfwAGc9GY64AKswf+xtPbw3X3BccETGFr
e17XzIbzExCph8Q7IvUcXkdpGTCtqaa54AA6zjhi1U0q+VHUeXuRMLsqjvYFXbrV
t1jCpRaBxrVHU222VacUD7xthCcUJeZHIFpOBCQkJg95sodvPc/Q1601Gf/rxbwO
knLIF9sJyWL4t9NiycRPWz6jjF6KlHbRPX4TVR8uMi3GC8rsWATdNpvUF3rwOu9Y
VFneyGXoCbXM2ZMXokBHuq+chB+91JUnZMA9v3WOo3lTXvc+GKYQSdXIeJlWAgpO
scOfSMYn5sXmH+iv6SOqzB51bODWLxm7ZKO39wN7/POizTHKqHxB2WxgajKZq3ba
Zd41jkRyGnXWAeqkDZ9/nmCMgCxrcrEPy+QNLc/lgEEN2jYIHz4Kd1ghzJO/nYTO
+WCfST/hRzPITCGRIzQ40mF6kUbUV5s2tE8y7+cXj1Il2ojHEgWkwtnelne7f8rE
jy64J8KL2feMT9k8hDfhmFNKMkL727yU6BIiLpcuTer06uHOSWEq3H0GiGFsWOOO
BYmm1Gh/SCgafEDt9tyvOr7MBNMUoDCwtgreMZn4j2Fzf19IxpPwO7DGY6Ou0xom
ZT95cxCZ6YV2pVFgBMo0v99J+XUukqS4+IfzIdRNWYsCKde6iUy50U38W4+/8hpw
EEq+2jwZMZMku55F5TTmTssGV/GbCDNPdVJltx/BWtuT8UqLzPEWDQ5shmo65xKS
ckHIbqOib+eYaeLObuj5W+KBuwTI6AntVGMNSNHHMBW67bSf2/Ym028aLWxRy9ut
YrAV/8tgodVhD9zXT2nF/CRYfDYLcJxXGvPtB68WW74dUsSq1oTCHGt49Po4LpEM
4zCsFVrWDgp0c8UM4Da/020rb8yOfoVQTm2uzVBM2Urk2BNgSUp1TNQG4s1A3qHi
ftvJNzfm6oc07MmZTA4I9qQeak4aObzYx0u0maVdySKegXu0eSCOPbdDHg3mVELR
3H3dEg4Vao8pnsmjYPmIog3yDBoX29oGrRqtnkpc6653cZ8FROWyO30qrccCku0m
TGHoL6L5jAWMWRVlW8Yo61ShWBfRmMjPmgjepj3C9bahrlkhgsfLWCJHyVpMaxEu
ipAajyEKlVy4ShopA/HS5fvqK+e6fEhW0GosvHpSXFZqsOpHW0uy1Zhx9pYG9gu5
HV295QJHN5uHdbg27PPrT0iOZUTxSluc81N83xSt6YlIZbQLohyZqSaQL7emWTYe
NDmlKWmc6GZvuSYJPoEwwblsJGcg01q2ALL6Krj3TK7XNrSzDQ00xgxYkU7b5gYD
BnPKegk/K/J5vd1X8NZMQl9b7xC7MGn11hjVfCNgpcMJiX6K9DO9Dr7NpyMcUx9/
G7apj5mku9nqP6UOvyzxdXy4u1RWMAYSMekbE1Qz0PQqxDIPqnidVztsRJiQgd+I
pXhwOCeu3kNWiq5hS4tFW6YV9qTW9EjlVNDHLX65avgHKYeJw47XFQcAz0QrJ36F
hS4fWROB6okzX+BQsW3MAQwRNY9HR6CrkPzIQbFYnJoRhQryCeDhquee1hdPRbzL
d8IGzuTjPY37bT38XkIgTzp/r8OUBMMdOxMM7K0SIq8utxioqphoBErUo8xF2HGB
S70MLydXc9If1ULOxaA0Hn47KOoravTEqf61xespdHLxIMBV7klhlvomE4betKXI
BvDmFEoTGChhA9WFsSi9S5rhq0Taq0KcyPfMmRfHr8mHVn1FuRnLQxWBbzPjLC7V
qJ409Du6jASfGb3u+sZUoz3O1NTesjclkjYEk2ZiYGvWVDGIFqqnzq99PdxJNjKE
YkMUZWA1WWseD8PbkSnSh18O52AVsQbuqnuw6+SlHl9aP7Kg/4HsO5c3Gf3OBtNd
eHWfU0GSYhhHSxTN46W8cOBAJhlmhzUjoG9DlmbR2wMe/9lx/8UZn16u1u5Wo7NT
yO+f+9HqaEgaSTbPAePY1yGQS2L6ihJBBiWnrcc1X/zUoHH0vRmTw6v/fci+4asI
BabCHHEtvA+SbxFy4GugG/OKLlqTgNSOZ612HTC+X+RYaKfkgh+JVcNMQjFZslaV
BzhYGQXKkY2VyoQTvC/sEOWdpwRmepALwEv2e4UsuUZzHPv3W37y7KvB6TvO3T/I
2jrYQJKogi9xQNGzh3B9hIk/bJ9jASAQn1XrkOR508SSgQehCf5mgeBZQkUCZ0OQ
OK4J0mPZgQq5CYonmkIxRBcOFLOkW6ULwtkQbDTsM5+VY5H1lVp6KBU+oGJ/G4Bm
u0EQs4TwKixz6Xyh24wSPR80WLNx2k4g7YrgTKDAh3MKdAevAvxcvepQXzTh1q+Y
RRkr8wEs0uVx5c5JRZx/GatPQz8XtNQA1/Dm9hHeMvDbQmAucVF/VSyLa/NVRafF
Fr4b/MZGoYZQbvzKs1V/nxgeMQY4X6q8P/iPCNZLcJYQp3zKIfMiNxXzrpaOby9V
a2VdYrv7gch52QU7Jp6tiD3KXJlpZheYmhTWrIskqX6K1W0W0RbS01pmQ+A0kaxr
QQlDNoyfoI8nXRlPXbbuHS+zVWpW/l+H7Igt1JnB8Y08HineToC7Loa6k+Kaw6ns
AkgVYqPM/2tQn5QOUnGBfDJWSvnICYaDLmAVF9wjtr8urtx6mxiCVpZOu5LHTdux
5UPXb4f4gG894D8K4laqYlt/Q0S0A643pkHPUyMEEQXH2g+12gGA/69U4DckkeG/
n9PPGXoAZEWYs2ktKQiEfjGhE+ZBY+scILwdM1xIj6n+nHbHXEPqozT/PtEo2n0V
3onQ/a++wroAPYnYlPOdvfRaEpfJ/xmfJ3AcRKSnc5EyZ+dG3/zkW98RkPFYyqL+
ZJY6CEiGP26fN/30CGJFj9qV0RmRlz0DJywscC/1DF2/oIOn795TrbbtBK0ifCQG
zvVZzW0IN5OhKBfvKrJBa71lErOFKzZpP6J3VT1tThKiHP5OFxLDkVnatLaDpjBp
jpZe4ldzhg8DJp95mM2XKmSSUyE1whvEuWWaGIwypWTmewM+S5k+Q7SKo2c2T4KN
rV8P4ag1ZlJrxzEQLU6iD03VgaPPJg+UA8t5jFl08GUGUpncaF/+TD0bL2q511vg
gkAk0F6Dh3tbG2SvcWKV4kcFptfEjHi3nfT3WE1YMI237kCU/4Eb7ODM0WplKeCB
pNnuUd9m324ZYj3K7v3jRFzT/pPgMa+UE5j4XqzsTby0XsKMDRw2ubgZNEeMib90
8Og2oNNGQrS1lhWYN9hbtRKiYiz4yuwWKrH/HhrPs18pHCdoTDJ1o1vTN1qEvWjJ
3dGZ2AnKIihKKTKNq1JpjLTVPZRILISy4sKTdhCKfHKd3zmqzXfkcXpzosB0YtgY
J9XLTFyCUfWgDL5McMzyJKNH71INbJVOAjQSf2gBorhkV5HyNwNxQQkKmUAL8Q8Y
vGebzGmn74hITphho8jQveFmHrUXAoUCpkQITnoMsVHSNMgLgSAlrUk4y5CXvBgH
BOKSpgr1J0f83EtXu4CKpNm0ZhS1dWtxULZB1XBYIQmx9orHA1PBZk5frC4cywJj
gducV7/NJCSvPTSjHZwrsBNuj+jwRg2+r8x9V2bxjlzDZa5vprdpCofMm+1s74mk
E4WQVLb4NZ4eTIdrup+2UhwjF4R5/VpYR5LI8FkqJ4Qv4NZCx19JLDUsfr0lGmL1
1dDgeocyPFiWP50QB1TZ9CUHGA2mXsSLBwL2z0IZqIgM+BGmf+a+6nCWP2z2DzvS
xvxkv/WerCQ838LaXdF8Fi3j21O5O1V0rYDhKke8oJTx03nN1x8kOaOmgj9JxM/m
dwaRyS5fKHjcJWZ3fcogop3wmoH/C+vRNLUj4mjQVo+LnUotnX7A6kEhQn/JqpGp

`pragma protect end_protected
