// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o5roZg0nm+YkGjVA3I81HqUsawVVlqkF8dkBDUQD1ghahUCcDUFuAiJymY/O
V9zChSSiyqkgmzObBV3E/vrWOAtwvZ+vSaQNVZHkl2aLbvAtmvPUQUj/AUnK
X9l+WEsZ+Y1hWVXMBCGIDwkL30M9g/Au6RfF0lguHvIEk0rE0uKW0+0pfxlR
BmWg1xDwkrjlbG+SuG3dPPWN6fv1u0LGHubbwDqJki1ctGY7LXZ0Cgr3nxPu
YcGjbmWTPLM2LLSOE4pFvFFP1dBZF+L2N0/hC159wquv8OIt0sV6HGNzv+pk
KzkbaeVUVYrxosmxaNGHrT88J+MGWCyuf9MmdV+Q2Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fnq16YNMStilUlm6awpEYafmlTQY08qxz6ZWUbdxVuUaGi3GACbU833bunmQ
hGP9m+56MAQlKOvPLugqfNreHos15Ec3F8k1CGmHvWjBbTqQ7FW6oP0D7Yd8
Ubuo2UGCQtnbfXE8nAghhZW5ZTW3co7sDvc+jeenB2wPzEQR0ZGQFHxrbPci
GzgeqvB0reLfMww5PcgU5llJ3XvRTNbpVvHtTJ+GAJ0fMyzT7D2Jmeo7gPKQ
aB9+khfI/qXo+cOICvNiVwnNAOpb9cHiqDl+wKG3A1nqi7Tkj4nP6FzVdRb1
fi1pYNUAkmljCitcoBjW/fhegFopYikK9dhTnsJjmA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ECh27O4aICNt2AYgc8rqFD3S4waa0YyFnsq9GXTi3KjTv7rDWXDje3IPM7DP
Qbtxw8VyvDHK72L20NqWlS7pizr5NoQGsaC5P5mdxkanF8duohFROHDUt81+
hOKKFqX3BsIAokTYZlU9SDek+FNHFlQFZf6gCNuwtmv1eCQWPGlElKzrXeHD
3kdvhMNnnccxtEG+kqgLUOyS3IZXgkh+NsHE7i+qydlgE2Y0e1ZHCWs+MKZ2
f3SUZ5Q+hMFF7oRvg88hlNL+J3THG2XhiWXMazdfpOh6HShfbSNpFQuALlVL
w7FomKQkKGk0luDZkUJ/mySkM6gD18dV0XXCNtk24w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
l0WxeDz/Ie6hM/nHenXSPMHu9Goa9gx4OB3LQHDAfrVwxTJjVDDB6sInDuFf
CleBZGAFGvp9TSplXPrZGvusMTr4FPJlOlOS/VTZxjDpfmyE6NaLzXwFFs/y
Bhmvz3Rofhf8mAUmi4zu050juwif85xB6wxBqQqY6Jkf6b4Y8m8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
UBJZrWm4BVN4GOx1KcqV6WQV2smdB4vffh2eMdqVEDkvrYHQ5IG67ZKEWs/X
hHqMD2j45KVIEx7gtRHHoqdzF/qQeYOPczCCYVDlNcZd0i7fPS5WkS9NVCft
xRFamZRLyrhM7OMb2X07jhBvt14f3WiGjT6oopPzx4PHMHhz+esqgl9KI2S7
KE6FFe4GblMOqGUGc+eZKiSohoO4B/dDlD0QZCwCIeJCL7heWw8F3+PSOAJm
pixy9Cj7bJKSolWpjGOyATyB0klUAeqgfr3Y74HfO9vYof7guVsmEmDV7aJ3
S2P/embJ15pULf6MsBJWlVHkw2gAs0nvxj3UqNQDlJZYE7g6RIysTbiqa1LC
dXuxl7tFC2vaMN38ZvkgpOZuFWYVLiYb5WZTL1dAs/NtjUJ72f6hibpAy8Pn
qpU8dUh5Yn7iUk7wGGrjzgGfTRWn8S2+dYG7VLQh63704I8hcEwAi27J2vtS
3S0pGnTsaSRXEIVrc5LZN2bDMBo5QOkv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OOlp/VLiviAXXm1ELNlQDwpn3SLgSoD2TiZ2QwoEZVVnK1WtQIsY885lezud
awZHa3zBoH1cp567bS5pso3IBGUyMTtd9EG8MAT8NYKk5tC1j6ATffG/uRG9
LhMVQLD5KlnGX0MPldxAeEQ6v2nps359qKs1mjn9eYrFh+6PuHk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eLtMUCFMB77cIJ+noQOTfTJrM2RRfLSsz3mdRtOjn0SWgLXKoJ+xwZXNEMQo
4qEYQbIO30DtBZBU3J88dpfgEJ5YeaP2BeYXFmSpwVqLSXob8GsaCKcLSKbg
3NSLW3q8VdRiW40/qwj1+YyAISN2ZZRmpiCxd6QzbeIoq3rwbTE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 50608)
`pragma protect data_block
yjwl46pRaY5JC8FwLPMpaEAg/S1uUypPlE8RMa3Ud6s9cVd/FST6qAgNPgqK
H5d3ECLVFt35xCvlXDq0eAZBD/abXSfe+/oClxO7IP+zBbvbegrAcQPxmKgC
FaL6hXl3SDfkX1PlzjkdrbtgXcbr5o5SOB2fvoV4ctqJ/HYkv5oYsHlCuoEu
d2EQtJBUP10+TDjB2+sb/HkRB+QqEOxZVtpr8DR3izag35EWYUecoXIw+ICU
bPix5r3U6z4UhQOpOj//oVnPoX85uXS0Tp34c4GzR7/YtxIlYM/tpzQg29Gi
5r1tfWibD8vqSEBG9UJtlRHPohGYL5eYEVF7NYzrGwjnmtA1W8f2cRL5ifP+
IvdUGRh5oiv4hv3YbRnDacB1j4KPFAOLNvmcGJvprygXy28teQTOKdY3zEP3
v26yk1DwsXQWF7Vhr2CnfFRUcVqMCJn3/8b39kmV14bR5yjj2hANf7okjfZD
U7YRTvI8f6fIzjeFjUZ9mXBNPFEncSyl47k4svbghdMc3qNpHC/UqW939Ju5
utx+8b6jggADvewTiGGUu+LQ566qn38CypZhs/PqUqxi07qTVjYyFmqa1nez
AOIoPBcIt2I8JY1ErWGtFebZftK6T2N6SVzp6PFuTE8CkY6ptRIJXYCBQBsZ
f2J1795z5vdCtwSY1QtzT8a8G+h7nNieUtRT92TsQqt5wRkE/HH7R3JkWdkU
PrjBzFz/+mglV62cLbAOar3Gkdr9v6T9TQqTXRW7c29qAQcT6VbzCy/bJeWD
LAMgtkbPpXEevbs+PJBkrCvjGZ5qpfW6TMGL20wnPk2iCCPGZ3c5vZ9CRLck
L9zzKCdPi3YRQdriehbYQujofUzjb3b/x5LZ/1u+1uLMRfRzAfV0j+tLMpU2
bdY6dfGULwY0OQn1Gyipa8kI/sVO/cBqP2NbsKmPMvfbPe1HZ3fRqr8Cdbbt
smQ8l5c4XyTSYE6RZgfq8hTZdRd2Q3E/zp7C3ntkW0OuApNJOLHOlQtGLXbc
X16c1j8XBITbftn+a4P2USuMjSf/ryzvg8FQ+2AK4TSGyGjM0yAOmczCix/r
VwrKiYOsTQnU4HnpFxRiDp7lKxdRcCTOwfRnAHrT4Q8rpIYvZ8Zypdn+dFXr
AW4ny8VuywDea33te88TlIQwxUylqbI32JfkFhuL5+LM2Rk+aeqkik1P6qKM
V+mtxEixNhOTjfqJtTz4wev6CU3n3w0ikvm298HNqN8zmbz0UK1iWGi0G7h1
xZbz632IpGwppMZgHn7DwZOhalkr/BgMg7q/P/0rKyEYQJpnMugwagnMcHWF
7/VOm+GGd/uc5/TgLHF/LB2EfNZFpsbzzvlON8duIp5WXBJRWS6k0Glth380
FfBbTgU88/qOBtB6PWeScZIfGYSZC8TpTAWCegUMgDZeozRQGEGlyQs8PGdO
LsdUww8du4h2rk09Hbd8vBUn/I4oAdaUBdZC9UujrtVlDVgsx3oSaMUYX35h
ClU23Kur/uJ793tZwkGF6/nOFlUxxz2Vl2pRUkVTW0X2dZNafiaNFCVSlCWW
HWs+MEgRzQRFKiqXmPk/gKRvh96Qo1TiQv8L3IYXRRvPxG2NLCcd2fzy/TD7
rZQ8iZN/T12vb7WKL9BuQw4UJ4tFH3q5F96FxaLxtBnggPGvXyHS3v6LCyxg
xjlsc3ZpbSbSfcJ5zonX8laeCs8urKnj/g4yHVkSepcnXEwzfNSeTy/JbegL
m2M+4jLO3fmPW+9MhseUUIb6boHgLm48xBWxbi0SIBYsfWyakrPPx8DCaORj
eCDWoSFD2eTOYIRFDjN96Wmhb1D2WeQ6Zulkv7JtA9YC9GrylaUVJr1/Z4ID
ZBBwxbfYsCwp7kM1CUQai+wxPU3H3bDlyfafPb2zW6O3nBHI73L9ENpPig5z
0tEEYpHshEm7twDfV5+J8f5UHkIVp1DkYGe+BVdqevgySireCV8AnnzN8H/a
frMt+nwDHSmMm64ML3XL2Ay4CCI58JINsniD2ACC78T2WqQ5d3wPfFeahhhs
oDCkqg/w/LuMAvJfqXHYPog+U0LTl+CN86p99gAPUvi8kCwxKrjM9dHA8FYA
rRFhot01RdAX+mX92Or5ZCzIJGIc48gz7p0omnk2IW7rKRw9OzgcghDvnDNr
WasK4tl2YYjFJj8mBrWIUzjsWAddrtb2Jpg7lQ5pNaWrzEWY3KhafV5WNLyp
ISLwkPQfGoLWSZg4ThY9Or6Fu+/PLdb+OhUQ/ceiVhCEo4tsmoQ3+W+xiFy8
/2OpVqjf9DNdNQDFyWOvZN7b2BrVWL4gpmTb5bCzWXpvy7VDQnKVSe47Nl0r
Wnr5hKGSP8/KjKfoLcQxFpJ0wXveC/9Cc2vazsGVQXuHBL/6doEdV4mKeaw/
DRpFIr3JUec2+oBjpocWr8L5QOZeHbUXUkGyJAdgkgYnLlLcjBHPtiSScEfh
LECEnIx1QiZgeVSV7J8XWi3ArHWcvrCnRCrIQHyE59ST8eiA99hjtmZ9YDVE
cnm7a2gFo9j64rGcfKpCZ7+WzB4mZnpFEWxkeHOBvlHEv/W1iAxLH9hN9BWc
ZB25+I/iBRtnh2J0+Sfwrjw5QjTD8fG7+KQNI9q+RlGnWl7h1W7X2otg6ttU
dCh3VBdlirG0x42puJwoMiAXcS1h1wdNHpfPrxlWKa/bXfDkPP58q8jfab4r
T/hDzFM55/SW77ei0Ynr6hV/gTPHOEmuNJ9oHnOHtjyuQ/uRMeRMCM3j/8WF
E3wMKJ5lsdU4Lssb3Q108uSHI9sQxvwCmxKVb+2vULgQRo75IteLfHh7kGi5
nWVerwUD+oEafxbb6bP8V/EUO3GNIJ3A4d/Rv9XnaRITKQfyoby66F33xx31
qfosqRfICbQX5YPwjHVH6WuAHYfqI1P7N8pE2WCGQrAV1rkK/Hs+1YcmTcLb
PTdndjri+vO0zLaTRltaZ/zIPTo0i2hYeU9HURJ2N3w/KMOTUiff9sf/5KPb
0wqA8EqvqsXy3cg9vBWeVilo0Cv3YYYk9rQGJgoUn2LhAWiFkiR+ubx4xf6z
Zv4Y9yG4yTVoM0KWVZ80EsQIXQcrQRow/p51DzLY18h3ZpMfvzFK6X8C28My
dO5u8cBkzhQ5/l6GSELodGkTFJkCqexIN3MLRihEX/p0WFBCEtGSTI6zZsnn
xHZUUUkebH/hLSyrhmaX7M157MbcMFEagPsMVsHODrG+qUBXLdklywwFqt00
Xq0P1QgBLYcKThskOmVTcxlsZsMJJaZO4sjnerT0MeT2nd3Y/kNmO9kpI0iy
anwZm1I/vvBQNHSwZvot5uoWG7Bw3bABMl8L1ZQZWTUP3pivYPVvbRIV+NRt
R2vtasWzwILtzxm0/RCtS9xQbNkTCGkPkyWRdQr6F8mADG5PKPgPizrgX0oy
21QipFqN7cWDya2SItWW5r3TrKE2mGDVvMcndC4xMagXoHgyum8DvNq0GdKX
C+n6uizecQB359LC+YeYewzrBeNUDG3CISHwpj1U/A5I5XyL9bKxjDN21N8Y
Q1tl8d94nRzDNbb/gLwLzShYb21npIqfZLnpJcyltVMRGzYgXBrreS0eMIYU
L27mQgPpZvYDqtAaJpvoBA3cg9wytL9P25RGRy/iOJBffjWV/3kpKvgVEJaw
bTOtFg9oLmZim/vnQADwX2GttOglIbwYbxwm8JTFAkRwsh6C2Iw8dfJNJYP6
crOexZKi3OBVO9z/Vg7cVL+eMG3BHyWOoPc9e3GwS8Forn6YxLC/nn6USg3F
WlcyPSMkfjDmaKoHw9lQkCtDOxgeLBWoTxHVWmOMBBxA2/rHrSkY+MWoSi0M
SBdufYkQIOsKmxaIHmsrMXEzsD75OYlltPCBR665Gx/akwbQuz1ZKGlGWIU5
mPpGF2YUkb/wzIwxVtazLVzfygy9G2ObKxrHJ771pDgVdUOtmpuMmseMQuoR
AXJLl7ughC/VAnxWCTrw1ZVzCxSML4ToUyFpH8kATttb/ZEobuzmodQC+90v
P/qexJvxADocz0YkCnQQKlWS9/qBTRLQaxvUiJ6Pt1P7AVV1tjxm6KdXyLQO
0nCpUR+mNVYB5T6a2QlRefDSWqoFWIJAAdio3ro1YgV0nzVIO0pkc7sUMyTb
25qIOAD6y6udiBskkMg3M9Fxc/h6UDc73nqAQjJ3c3C4G/B2Wm6gwPNaOFFG
R2AwdHNhNrLkszVC4WcqzjWisqzXEaHIjxxc/V8JSD4rDetTaKXS0aKEGPi4
3VPgoQKQRUonfXmMOx43kh3kdme78I7/FcUuEJLm62hTaISvAm84HXeWSHNp
Vv4oPknQf6GtiUB9rDtTy5P2TVioK/N2kIwW7e5EfMWgtio2l+WXyjd74e9P
MXI/9OtXwcwkJnhYYzznbSdahjUeAyOGMwaX/gw6Lo3VIcFYgZ87pB7DqJi1
8BlZE+HKUkrWUJytljeJMpwR5rrvaTJdcZTIdoMj8WYlEOGMyhVKFwCCur/1
8mVxy138d6rR2w5g2SDa2Qce/T107wFJjJRdXUNgY0Fhi4Zpr0htyaxfR9xw
FWBWavjG/mdbXZTAt3VwLlEvm6O1ha/JG3AkO6IGpgoy3v6s5L6g5mKk4TUY
eZxuErcfd8Do3GXmaPRbvtlGnZar6mxqLdUH7dYd9W1wLBrgMF78NI/q0nab
50SjBRErtq5Om6+hIJkqpCaqTOLXxD1rOzW7bOqzW+c6kDLTnD7o1z2kcHRl
BI8LClfDxr1U9TbgGWfjkzWuDF4iay9JDgrMeuMi5DrtVMNHYoNNBxnPkVjW
BfF5agJLWsbg83LYiQqXR5+gIZ01fYKg/ltw1jL40wb1RvtDlT66lTCBn+IH
TvWSjeuAlPHLbMYuXxJxYsMDDa7SuAkZ35bkW5yqIzkVQkqBRmadBiuZdGrS
v9i+bZkUHKC+IS1DSE60i9ad8IS9UkumwJh3dMp/evqTJsI39L7f5Trt4TVO
5K9WmD5Du/iMJmiwXvBMmGFci4qTLp9qHIO+QlN112ulmzdqrXbm/ARPWb75
VAHqU9fxWWfBQ1Ai0Q/AmP34VqiDChQ+ZuWEEs6u2Zla6z/dvZxtbzpMnHFp
FP9JwPCqunUFfGjCOznltL562mVJ6gnP4061ApJ2uNeFqRSx924OB6fvFqpI
NSkLoVBFivObqH1wILZYlWBecDRIU7ofEz34TZq8xnfYlGXsdhkoVcvUpjdU
DE15zjyYkE5WMTf9dFQJkhQBGtYYQdiBnKeFhYjNPQJzz1oX2FES0TTJ4tAm
CcoiIJuLo1Uwm8G+172DHF5EZvavVNPnH+UXA9jpkueX/M9SWvFK4DXC8kV+
hsF4/QdlG1ihBySwl8DSamXtWeIQtBW2D/Iq2h6W6XtwbB9XD0gEtygiye9v
8xSZ8G4/r1llJIn/3fB2kZjgONATAnY+7//peC81A7iu1MwMbS3p1ZxiE+KY
of9ZWSgjwpjeEeAkwA6ayfVMz16oxXoeOlgosJFBQlIM2eCd4izRqfjDrSe4
66n1cWusRjOho+NEBUu+aoMoUQ1x2pZcQ+DaMh4sKZ+PKC9g/p5IXDWwnCwX
Cnq1m/oIpge5au7AJUUo+y5Jr5dVuosDyOXo8aHq2l1Qht+y1qkijIe38lKk
5W5MjlhjWRNS97YN/pq6jRVe7+I7kS3W34QCwsX8U2cMDGodFOLNIDsDgaOC
DYGNmK8KWT3u2agHITIUD/dAMpqM2vYlko7FMDKu9Zp8NkMD3AnntrbCSXz1
ewuv5A2PkUkLDo2yFwcUyJkMU9H/z6TsBHKaJDI5SZ/PeqgJpzzOhp/tA4vV
RFBWbqK6RG+PMoekn1rsg4NBRwRl4fMJtqXjDsmcejvwg8gG2yBTxh95HsZ+
jmyQhR3EORYwmCR51P1sjMUk2QgL+/gPrPNBS7wdTX+cKbzEUrn0m6gLFK2T
rbT85l93WmlfyLy6amPNBuhOH3B3upcChhNKzAUpB4cd5aAqjijSUX3huj02
i+5UCqsT4EPxmDEHPFChhMIzPfB8JcxRQgnvJyShKK3ap8lz1W/GFeh1e510
cFbcPQovSa4bvYwNEwiUNCAH33AeZWueUsp25dUuHrOE44AK5o/Rl6GACFFO
1mC5FB8zC0iqV4lg5qtnR59EmQum5yweCZX/bv78IRPlzXg0/vVvQqesaFb3
ZoSUaDZkh6onQP84VGXHKeXLhooiPuV/8mhm8DdoFU7bjvIq61DTN4+Ru8vS
Ztr9E8UgfvFBy7EoDCbQQFVMUhasjIh/Fix2oL2VuxMFeAdcbSY49BkiT6Gc
k+QE3GyfUDCg+S4bn5MUlHRkz+ZzBHo9t7lLWajRRInntv4vj5b+8HEGcxcW
9BVmwjtt0PFFeAFb+5f1MgCenDXdhoqiVV6/suu3UiHF+oo6xso0KaKu5J/J
hioMnUDZKa9belm3+Ozr4uedZkkil4Q8i0tfqT2CNoHXCUkVhgSU/tto/Xou
+DSB6dhOoUlUFv4B4CN28hkSFMx9aEOGkrYuO8UJD0HJVv7/DuJYxJe7TwBJ
s8VJrkZ35UwkCHD+Ga7dkfvBrCuDB5Q9bWkUWvn0N+Bqiveg0/b2GL+Etg7e
6m4el3MPpWaGbeIVi0zv4QikAuZFbVn8pM4x88WBF6jS/ZGqlpx881aFeo0z
Bqbb6l4jsM6FjN5c7O7c1vI/cyKB+fD1/ikIToK9BEi1jvpkLXDg8v8T2ptD
aYii7YuLmHJGULvTbbc2CLOW4BgkF0oNVKXbc43SOE8lJhICW7hO5DXEl4pe
ygszPzDzRq9ORZ6rKp1SKtbQrWgFCrzWltvasFX13deZjhM/R+/SH1wsXvo8
Fck0rQKpxgYOC3wLvYf1k2sZWF/QP2eirbOdZXXPifxpMHQZ6kJHcQO21MXf
/Y5nRtIXLybnKAN8ErGTifG7jn/wc8dT2CmxF53zG0zOYEu6IIij2+ENTVDu
Z1nA0xm7JdYukp/S00eQZDz+PuF8UHPp0pLPGsicbml8YqGGnbfIMGD1Y3j+
5i9FJ048Uhcn9lfnsAnpKjyjhjDZh7KGqZ6Lt6ll6Ohb5XSDcA0cSh549Ceh
wadVL4c8q+Zhl3aRvdeevAfLBLIZMRbhyMYC1GSdaLDEe+WfI92NWt+ZYo91
zLtNh6XOWSdhXm7ki8DnH9Bv7D7+BtETxGuhwhMQ+Efp7zCaTyV1Mm9AroVX
lYUkS1cFfvpeKYPIOnaCvliRNC25zue/PQ2g/HoWcY9o9TTsAZbcyqq3XCmj
ECBHZ7JL2vf/q0/Fa4LqHRQ+zevEALittC2YHSYnDNoKxiPKLdE8pKogtCDA
ze08Kdbn1G+qmj7orNiocKsjmuYMyeQQFOHpLJfPiquJeEpyR7UbFPct6OEZ
f46reLV7aVqCbH4etFJigIH91P5qiYEJ0DwFMHom5mgS7aEWTxWsZfSXxcE/
2iWhAf1NsftVtzYRGt7jIAU+EZJyccHO7W3Jw/T2rmZC0MgY+4Jhx5Ih5QKH
ZoTq/a6d+iFYmmI/YKM1D+46L2vxr2xcVfTGii+8jd243p5qoWQPS/FQWtAo
n3QT78W+GoOFBvVu2y373MHVpJE5aKTOxtP8Z7gAcjt+FQ5NA5PSN7xTuQLJ
kzV50TJqNgFs6MW+NFGVfBJbV3L8wCiEAj648FVxRFMARNOeK0/DIWUKkOtb
qbmb3AnZzGs41x+jCFu32D9uXtoW2Exd0bqYGCZuOaFGWqhLDkFrYhx/JHHd
7KakPCsQaPYYY3k1Xch9nZRuc+la9B1OEoD8XA98zjZQgZ1FPYir6Wa/RnEU
oaTcf8jjTURbaq3rKyVgNoJJBhY1shggaT11pW489qVAn5O2ctRR2ewFx3OX
9HkYL1deAW4oEVmYnRfR2bYX/J7Nf45YTfq9wqvfzjIqh3gagRB1TDNu6myQ
cQkfK/23iMc4vc9Lw+AD3Fcnw//WHU4BHLrb1pvHn8TWCBuPKxCGPyi61gqu
6YRrCtQqk4DVymf6Fy/jwHBezdZLOnXBWTslO+u6I3mvnHDe0CYYmfyjcCGi
YYlwjvCZDG1XPEqAhn/m9wwroxRtmZc61Sc2UuaWeWixLUMJP8vSn9OGqAl8
GIqvxuFxP/2y1+lLe9p0hL5d6S468nof8G9b2BZ0UycYtRrWvMJZViHagj9O
QDeFCrSp8RzqjdKaFSpdnNDaPYJTz5POQ93o4DmfKEJUGpeTqhX99W9ZoqUI
T0fKV+2Pld5AGiETnANJ0ooarpOURmJbkoXfQFa7UmzfoEghOo0PcOFRbxIt
jcye0J1l1GhHh9IDcqOLHBcRZJipHewQXirUnTUzrD49lXYhuBrIpagt9G3H
YF19cBr/BCXc4N+ziT1BJpMl3dbWgn1UH+QkulNYWlRhku7/RSswAwi5tEK7
nW0LIHND+sInaXgO5jB9fHLA9R59+US65rjP71K6/xiXLAD/+kqvr5YViFyr
npudKviiLcMWED2vySVYWy/+ZiWwm50tnKLAe6j+rmA3YSwQE2E/3NiRhLNY
L/xVC5DS+hGKpgS3ErGOc1zCQ7WXZknEbY45o2wUeQEY9xDeKAGenuEK3Vjv
OcXgow6XNL0WqNufm6h54Pf63yKcuA1mACAoztJMx6Gno+81bhtDxs4eKcC7
b5iYWlbb+ymW9BTPCrPdqhfDf7fX/IfslyDB4ImLAqLpbK301cE053I8jiU0
yUNgb7Rn93HM9Fq+QXVHliMHD2t0n5jH5gonMNK3cnqQGw4XBbdXZuZcaueX
USiS4Kny2HKelkZq3OkwRZD40O6EGWBrQfmdndZ+3d62OCRxWnRS4Ldt3ggx
TvYmu1/7LS6Kkx+NiJzE/Fjjkh+EhIrS5cVXAojjd2E+QbwRU9SBJFhJgMvw
YX4srfjqVGNdvXWArq5l516LjaBN0tO7WKGtAWr2qmuE99bOUlmz+ceBCqzp
elL/EQ7XfeFEU9UwFA7771CJpoYM47aGGqxxxRqxJAV5wV/wzEZDdxa2ejAK
sRpzo7K1MIZmCNkkKM3Rt5JMsmM4qmkey1RezltbDObEatGBR4lfDFt26TeT
0Is4It1OEdMxPkRlD437F2wBS2SxbWKAaxXio0JA/fh9m5amddLd/jf38Pb9
iJSkkTDN5ZZCucXwDwDbfXZ6OJ7bB4lWgR0Kbt7I36023qgvm4G70GoZH1YH
ccbS9quMua2JWDf03ILgZYF+NJgfTQvC1tXrVqpBGVanjgijxWp7GsKDwIKd
uPST+ivBJ/fkKWjC5KNAuAObXZosODxqU4Fcd11WkiAleaBM0PgPuIGgQp7C
KR2/qiVueqbRsx2T9upg5xW2UBgNOYGH77TdGrKMzIfbsk51BfcXCPGL4Swy
k4DI3EW6/tZ5GIycD2YgzrjDyFrI1zl0D0xKIlQQEqmczyBSUmlZdYPXF02F
ZlxUfDdgob5biQ9/fGBAjDnUto/0S0RJ++JJOYx6H/ZqTrAvZGsCctU+qiL1
9wbW1eql3qx00glSUfv9SouFx326ZWF02jQmG0wZpi2xNh+AAvPUY9jQ5vNX
+NvQE5hUt2VN8wD2CZ7eEkSFIrSdkCAi8Iifrs7PfOqRv1imbfYL+Twts9WY
iENdUDZvoq3ZNWFu3I11+qulAkLnjnn3kpEob+hCuuJJ35idu4jeQ5SW1Wis
z5mTJH1SthxERnmCEB6kdhIVOUTv5uSf7ULAwnoWJAOg+KspHI76CNl17G9p
ZWTDP80NWGGF4Ev4IZGY2vz4nTef1VszsOUsuQP7TJKGf0cvJBLm1BBPAUHN
8jYLqPx+fgybLBmqsNoGkoAeVGIpeIl+2DQZqqlfbo+3sDFY828zcWuJK1jk
xRPAJ/vrPfExt9l8qXvmYxUp2uxoq+zdI2Z3PyRLX/rR1jo0zES18VQvy3KQ
n9moa5kA9uSKvvBkRT/vAIkQZKH5+dY3U/McR1yz1y1GSfYuGRr+uaQmaBJe
zOl7YSxv00tIaItzYufnlxfRSf1gKsXo2vKlaN2f0C+81ZrqMcSWZp65ySAS
hSZRcH4kSVhogNAEB8tIBczxkzT2UFKWceOfkRQFyoX2Ec02Lp9CRzG57Ppb
ipPKNOeFfklMS1YdviN4A1AggksNZFd0HCAOb2ikzXzW9Ou1WOrJNwcg02oS
WzuQx24bYpmp3esCBHNXBNhhvS1yKGMhcXoYrEGX+gahFdAdgJUYP7AtP/cu
gMVnwKwISXleNrcRuFtWJxD5VywDCHTTPIx/+nUbAGOKlt3p0BWpYO8VCIfQ
ILVPm+Q08d5wMHEdaJaEUUGeuvfn3nvK5rDUzQevOb+WXKkWR3LOAETcZl3l
LEtVvNaypaW7j0cyzPK/+42yPwSDguwtdzdZrxcVsZDejY/tRbMs7HX9Yw/p
BwfUug+2TxBmNlfkVtJWnCXVDpvBT9XT4UUhkb6Rwmo239ZspL3PUHVfJ2Zo
n9uv6dTdIHa3IFwekLIS+yX/jjpcOzFzz5GzpRlDNFlR9XIfW4WIDHDuUB9B
bR2mntOBWAgueli3UjX39uhd0gipdHPSPxI/Tfxpw537Z2uKfSdff2ET8Vkr
dX9D0pO5BsUXtn00rx03fkVyCnjP/y1RJz8iFzsVMsWrXMcjBx7uHMVdQGR7
/K5EkroNfyZ6ulZruwH10rZPCAvrX31QRWh0arsTZz4p9VAxtqJiwkaIW1oB
i/C+IfILlrChH/q1ERTQYMry+wF6xZVbdfqQE9M5eQDq34mroHci5Ctt1EBy
+SMnHiQXwvxlIHZUaU8OP9LrvDybD2XBCYv+bzDlLJMtkefP1D8hc2lnOcs/
1MKofsco1oRoL8ZNOSqxAxFCg1LnOje85jmyfRAnURCuFOZdiBOyta/9XnYY
PDTkQhwpWyTNzBJvBUyPz+NO5yi4/3dUFlIpAVO2zyiz4tt99/ezkXaiSlB1
I9o/LPFBEfR/O6lBDtxFDlzxaMoJEZfDoVp3huvXJsiXkiVUB0Ao2lMfbZ8U
JvOP9HkHQVnJa2uU9UXjPGtrCq1iny8QbbVANh60iHh5L4Cu/UHMnEhBBCKd
A88q3F1uYDhi6xbAalrC7TrVr9BEQiNEJ/QzRXVVzDFCVcrI0bdbCpqDupKt
cFNMYEbi9l/0+xr/TMcAfR+ux9bAYkB2FoXrJwBPYunlE6IeZAueA6xk/eK1
EIcROfi4ukNefAGO8AcFax2lRwgzt7jqlXUrFiAb9OBwLFDTCHoHHaEDtlF3
x3nZK2Qo/xoQZYIosCGsje4XY7wA7aLeQVI/se6OOohlW5M+kxL6cJEgIyTV
0kU4ep0IxJqDLbZnKAfmxpRgobs7jOjQUnkHVU3W2I1Me55Kh5QZhZXdTCJ0
sqd5hpOGVIyabqVblzM0fE424YlfgpyuHAipMAG7GVFWxezgYX8XoWQGfc0N
9cLiwkTFgTepVEnrouwcBt+WO37qLpxwQZXX+WTA42Rr90F1VOgkJx2GYmH/
cP6L+uFU9aLqe9CeRXSGVnLPQ3Q6rxCvKJTLvPS2cg099/gf8OZDb1GKH/7d
7kBBsZXzAkgyybMzm49I/LnXHH6ew0pX+5iRG+hP692as9OV89kzJgvAgrZu
57gsC71bjD4y4SanSjODbl+BpxJiPSBsJev+nxQczek2RK7rRAsIvtI73/fW
YQRUpJ8l/aXUH/rEgpVFmp5Sq312ly+CU0rSW8sq7Rk0Qf42yFGuc2Dc+TDF
YJ5wDdfSp8IJemGr/tM7cmy2cocjKLxQk18D7MQ6nylujExSOZ2ca+vznfHW
Xz8fiocwm7U6dFv1ayPP2PoynLwu9igR7VCWkcqdLbdGUZ4fY1XwNzjow/nE
t/ttnV8fD1fDbiUwvTT7I1ApbbInNBU3SO/v3YaYVmcTKQ3zrV3eOOdrsheO
XeQXV3RSxV6+991oqX8jCOutyTiyJUY6aIxtyw8vGLtCNBGGu25WvzvUjdF9
PkW24lriMtE8d89UAC7e+rhnNbSIHYVNiGEW9a6WJo5yVMCJfjlG+fOk4wNZ
9kk7JmAb4AI7ILIRy3yeT0xGgdcezCDZy3NqMwmrjgoh83lOeQKyy/PeFgVb
u2pna0SFPXz32MyET2nqmZR9L0HdKHtfA/5UncRqpox15KE8AtgWCBE/qv/q
1oCeBzpAAcjq5kN8VjcXPGSSiV2t4xaScDzfzxz/jykToS7aXJlI13L3BT1q
Ob8tjNrK/W1f5RENM3BqIzNkaB9J/PzJJaWxA7QIJJ13j/DWL/f5oc5dUS0s
wBve3qa7jIyHOlxR16XEpv6vk+b0fJP1iT0zunpMlt3KKfHMOkooULnp9biI
v8v8yeBxPYIhNsJGJd5uCA44mTqQtjRdqlmjl5Tp907fshtyS0q1sJnOkYYw
MPACqeRrfT1BbdBV5dmIdPL31m2sPynSEvZYRv5HiZwVsrBhMs4cUYrbqd8+
eM16qHpg8ms/N7hqpPpvspsYiZgEiI45Wq14AWsT7lIS6LGZQKKMH2B6G7Kr
xpd1+3KIltJHTlnxXFrten6zPriMHwrSG2aVGYPe5kmdeUo+9OKoWA+NC13m
JL+L6zjOjv0ldrDIgwocHr2fOjY1KV1jXhdbeoO7IPBxq8cNq02FyHxhqinm
QPGfsSjbSW4otSkk6dRICkXhfBFsFTgC3Yj6a0fphLsNeBqHnkXi5dcfiEKZ
XGTagmhjy+IFWb6v9qwJJE6DBhcMLOb6GmpU2llKAkaPxbjQBiX5TwJHYpmL
J1U3HK1QNXJGL/JAjCnDFw2ajaDX7MlV6d7sRjX9W1exAcS4qe74XBsJh3/h
cCbJrEitkBSUGXviQuSFo+27OoLVD66Aew2JuRd8znsuNKKJZSdBwo2uWjT+
dkQbqK0M1zd7+Z1GA/H7g14z66cu1EVbBcLxm72Mb7G7rgqTwmDedMKjGUFO
5TwmoKICMU5b1wGyT+wub+vaCqtJ+M453EB8m51yxE5yU5F9wOLgVC8l6AYS
gzCSHO5Uof0zuNYN2pasY8BtDyyWSI1LzuNNF5i5MauBtWTW4ConFb0n4En2
jdfhVrJKAoOnOLDuOM82LI9K3T+yggRmSrgAltjIlCpK29OQRhCZkiq16JE9
1RWmUDc6wo5xdplXtvdFNc6kTORKnC5frSAsdKy7fe5gLUIQ/ehLnruKg/4Q
2V0z++sj+oSA4RuCWK7g9saUG7c2R5mLMnIt9ymFC+IcMlNSNFidOQekEp7b
JSAtERnIhKbTDepXCoe2b3LsN+VlSKgNkhj49htSvARbmwpT07cZ6RTQrktg
eEjaqmEZU+foGXqRW4rlSwiFI6gKjEXcI1jnF97PsOBZpm2dQLdm8xipKbc0
Q1lISKK+WKrKvT72ciaEmaf6mlCM4RfjOAWTvXJdWb9/sFNnYZcacbr22XZd
SpBMXstM9XEmR56qGLAmWrnK0NcWGwqslrZtZFCoLdULFY3OkYd2/ZWzjCif
XlAcLA6GgjjvfAf7KpJAFZT4IswfWycFrYjrmsrLPxd1v7ssVV9+FX4lNNSW
fTGXGgmbQI5+dSJjq++GFGWf7IrOoSRGPlRuMa98nMK9mHqLG2IvHni+C0lc
knr9r+1DPxsZEpif68+j/pSdJDVmvtp3/H2/N8n+HCQyX73ciJMcP29A5KHc
7BSuAGEiKi6tOvfFABYt2wTCQkEquaX2ScyGoghAUVRKow/sUM3m5YYvgLHB
Dlmqgj9sMj0uIS3YCidypWdtzh3x88nMsAXlDlZInrMNf613AwKOJeyBnJhd
pjfr9B6L6R2WRILV7cw2BLxVpgI8p3TMmrOLONqJy4QBe44zkNx80EVdXbTV
Ri+YJ0T8dDIKdVrlyhVwL0O4/TRJWyfFR/DFyEh3ANh+6Y5/O2Za5OqvHLxg
QYAd5AHpfgy36HAafGcQmulb1qaLRnqj1vI6wcDeg9jSZtCQD6cqdCNDzKp1
dskpiWoXJ6Kpvw0jhrRbyRkCpfRhzDqrfDhCWN7d4Az9szvzQ5WhEtnDoUTu
KCiwFjz113JFH3SdilxcE9zQXbxTaeA4rBoRDe5+5IO21I+2CdINeMfrfYzN
juBnC5XFBNMZ+skOPQXPCDg2DdYqM4JSUg2dJntnPQFweyAz87nsPCHpzIgU
M4B9t1EH6KtHvcd5mCJbJ+WTC7j4nKtdk1bKwhMP2ptcjlj1wLQE9vX8621b
3U8TyyTAFWTi5SZ6QEXUKs2wUfIvUrapHI0UmRE32rgXb9TkTREH/2q89HAP
WTWDQizyXy14D2HxhZQHhLG783tbsVU7vAqKquF1HK95cMcoJro3UNP1yteX
KtU4lCB2RFkw74AEC3k/og4et68Dzr6503/zPXAn66z61katwGmVQm8UTszQ
plQDnSb8Zsxh700GDirS1cyp6KPrAYGhdPhNdM1G5dktVCbuLoupSxabPmKg
113E2ky6jkLRT1Ch6YQJGUDQtb3uLEJWpgOqvQHWcTmK5i+2byQBf1hl48ze
uslLaajbrQm2g35orGo2VbGEP4qooSw2GVrEsrg44hqSBOlX1dLZhYMv99OO
U22oFbilc/iOpgjMyrgLRaMi/wb+bo+hWKjjLt1UBMnc1dl7Hu9aBDTNVME6
ukAkQ9a3whhxuQho97FIRqJHkaECHgPVs/CLoKRLyvzrgZlTCejCivW5qJWm
IC1mwyCwMdWlVuwyXuIp+K+fHe7plfRZFng7hIWuHOmR/pIVqTUaLAkDWujL
qdlj5vyjK0SDAZ7zq9etHn1MTUYdBMt1Qt1aeY3vEdG5AuNzas8Z+itIMXso
ChOII2A2LGr33PSJRkLmim1HhV39L01fvICxpBUsZ2VUERlRN7oGYjBesW4X
ljDKIhnm7PC1+qtcMFADBj68T9RISh5F3cIIRwtDOxai1TqhWDczvNgCewyt
yYV/koMNvGdYvP4gEk6+ovX214TZbdqHvfNrZiTmDo6r/Laul91cOh8SxkxM
qjGNjIyHqz9igSqPPooR1BgHVfz8rHfDKKxh6OI7HjagioEZGqGrguzhtkr6
NdKOjHTkwFNr+UB3Ei7nP6LkX0LU9WGrG/2vbJV69ZOORweIT2AABifAkRQ7
t4foS397JNl2hcXxWazeCQZI1G20FZFN5eyJ277UmQrVCWjTZQ3b9Gdpb7g7
MkzSAYv0uIH/JjqqyLDRH2DzECtE+7mE4h0FobNskZOaiUniRCIGt6UkPaIl
SfdDCSTh/PEObD8cF5zAMft9RXtouGz3+6uyjXNywIeOP85LANvFWKPNIyGD
145qVdnNhc2GiDnx6kwqBKKf1xohjt7Wf6iRnSGSeVHCoBWvxtOhPfQ+YUMy
jNI5mw1OITlJvDjtoyA4fzlrEf5Fmo/gOe3Pc4/9FfBqihz5C2Dxquz7/StJ
rwH7XjxcTvNJmL9c7gF4ZPcNi064w0B7tluAbLYMu7rSOyXXF3vo4dtino2W
eVRJjZm+ahX4Q3y1HdQNnTu9kbpnemYbU1mFDtYpyEZ9YiMwvseyHKy9Tcg+
Um95H63ehOn5IvxRHm9MY4uxY0VTxMfMKI18Lj7VvS4QvMibaPBGxi1ctsSH
hZoOvdxVMiY3ugya4KVKmXm+ATdI9YHxg1ELZVwPZY31TKcDf9C25KPrQQa1
qYb1GCFcD2wnABcxZtL+4pwRK7hT55qNMEv2QS8bYjhu5RItwftiUIpMGEpJ
zR2bolnkdqRaqc2Je8WI+RdZvzf8g5aS4C7nPGwKY2Gc09TN9L9XWvIJpyHq
HH5IzYKRWJMiwJHn9yCemaq0KrU2WXTfT/DHhLr3EmIb+GI6BfOSRR4kTbW4
iCZwZKLPO8w0CP73sFrTafzFVNoRiU2Y1s1m58thpmOUjV53g41kOAsrCIxY
Euh8DL1MVtCqx+ohcw77s2/z1SdMbNH9cR8iHBna8UUs+2GyHVQLnb7/2iNT
IzuOdFA1hTLylGl21175dtIOCKVLzsaM6MycgKwUE+JKGy7C4bD9ZOzI6el0
Dz7IoaBZi3uSJW7B8joGS0cWZhTQeCZt8uoA9Nll/xsAlY1qmSsrc8HeMccL
GZUWQn5QHi2Jvw1SJpQJgwbJtIJG9I1EUGwOsVLoGbFdWHsWnkZUuTYD+RC9
FzlA82zfeiBKC67zYtzqw6Yu5Bbo0yZhDoODNNCpCWNspfkjV+bnT5V1yjG1
VX3Sg7ZaFcO5Sy5Jv2D7rcNX7owVkcPYhtxWY80kW28su7LjL+9pMwQMu4LY
T3vuiolzhBzxBqaq4+dfkRhFojoRZ00Sy/CEamsmAtN9/WdXR2rLdcHZMBCD
JyVcMxTrTeQM28CcC8rsAWwLFxq7cHUDBoVP8yWEntaTbTDAkbwnPDhlnzdr
EuYkwJhfVbjzzOhddQJ/oR1hBYhRwhdv4zqNdIu1xmOBlLLZ6r8Rj24vyFzr
rGw9e0ETBY3JGTmUTHQBy9U6WP9oP+7khaSc1FCRV71GKcJDRpbnYrowXccY
g+J4dlVDL/eR1Q3ogO/kFXrahJB1sG4WrgphwW0sPw3J9e9fPARPvLmLaQHv
jRtQSP0+E1QpflZ+j8dXy6/LUE2E2i55n6D2jE/rJL7kgsPphu9yK9OJjUPR
pgPw5RALBbuxEyD+fogRTSsO07MnZ5jxqHmiUDzJxQVjC5ibtz+GUA7iTEOV
6iCimkn+uXqrD67IW3uGxuWsfhHQETXFkqIOlPq6fR+H1ftnI7rOmCKrCI+h
QYum8WCSjPWroIYPCusjarsKfR/5srqG3xwasSi2A5xe1hG0Yafcduo6+f8Y
SvCfYQk6O/YrrVPuFwKk8KeuuzEuQAmg4uoXkMphs4TdC19M5+GGvqqNkZsd
7WOF901LNIMXFSJtKfQejazOK+LTWo/ay7oNYr0VmNrgdcBWMkvO/nPUm8xS
uFGujEc9TON7bVg2jy3zKT3e6SzBUgw8eKXofQ/QIoy6GfeY6e1mis23uywk
F3ktb1OtM5aotYqcBKMWCuxo7J1K7vw+hDwHQ/8wYQlfY7zTtcsFndLbXvxh
cZNYsvkHxgmRq2rLSkeD8PF4f3V8X4aesBh/NSs9hXU942AIm3luAaJ5G8pX
UgarGXTq/huESc9xZQNP/zmWW/56DiWltdHcy+jCbZCrH3qM1R3ALewsbXLG
hc0G9kf8O42scZPl2aexAP5quuDWmYgo6UA//kvP/UsLLZQ9XLuiknwkQPqp
xZOu5NRRQYugXIRh/CwzKsXEm7uTJ2nD8BrlH+gmnsm+TddzHyUTnKhJhtwU
GcSkTiR4f4jDsvgJKIlE7sSKYyp1qf1jaGij50qPJ9KnBuBlQSxI4uVm30LU
CY19Vvha1fnPUPpFD+VcMEYcsVmeRsdM2YwDgpM7LaBiYx0v2pHQwKHNmUCm
6lbtfM/uuSSPXj2TDGyhe2e0nRBMubODHvcl1xYJ01688qM4EnZzsffbI324
weUdIupmjTFDZhUd7Pm5xv1s5DQbamH2rBTBFMCMy+lete6ILNecNoSM1gdA
kxnnJqjBblwJD7MG5Y2y8+VkmpECAcAc8qk/9uAcd/lu3jU+lwJstljJuyTb
ZFRsfS6D4sn6nYgEi7+dr8e/1sCCkofBxmCxObM9slxyL/+mxcLkDpngK+t9
AJd58AFAYqOt4nCC5kSMuvHrFsl+8G52SIP2EnlTAXssoceuuHiK4D/BPRgg
9GuVBcbY3WI8+9abE7mRjIYcInKLM/6+VQzEdRXy8eNJAFjUYzJ8g2z9le2Z
IOO1BctSEuZlCIsjAOyUkwH7xFmQ9JzmfM8hyNu2JK0RAUURKnwoM8d3Nym/
V5e4gDU4upWckS65aeJkeUPP9XaFB60fySfhipxuWAyfrhYjZtDdFjpSu/sY
A9GDXiE6irpncmVhtdVR+cyfF2m1+2gxYM7Phx+iQ6zBo2ntbHkzhs3xkPbu
vezFzF1vdmoVv+7LumNkf1wr9JEqrRhiA5fnA4eeYSvLQscylE3bLovSWH55
Luo5wwCLHrn1hHLLni2+IRlxnYlcftSKspPGSP8aMNy/6Ujv8w1bdyCunJyE
AxkQ5afd7XfBlSdpi15M8gWQXguNyQBFPbiZmFIHldxmJL1r6wAow85FxcTp
y3ZuaVi4uAwIQTolZB/tkmYjlIq5bcAYn+2OZhYZZzvcFp3d55x0uqiKGvq2
KYesksl7ensR3VlLpviK+oe+yTLqoA0ujA2sY7LkdGdJk6BntHGWXgAdmw6f
B7EQBYtgffyTDwQg1JKgri/uFWvjEi55K14yv+HHHhISLbfGlYBsSdtajwQQ
OUfeSEBuLp8Q60Sg4CkYSlJmProVNAQOx/4frY+y68MHwNMR+oNZwytK+1jt
2T8CzZtJBI6hugoOcl0TSNP5xr+VlQ5N7U0m32tXfIYxCu6gVxkNVDQC3dTP
/psg6JZmmgY7k5qB8Jy5GHmU4n0jk8DVxOnNYW4Wr51t/Vz0nt++Avo0S4Sq
T+PVEJAK4KZFaS/UJsP5XKJOz7uplnggro481rqWpm68QNC55sfoEl9EJFjD
Rt+516vZHMSIO26nYiDw55wN2BOEA4z2G2LkjOjGVMmAj+9UgkaQNHJKLLYw
OgcC6F1d26/IfXg9UFnQFWQq1pAaojv+o89otSi3U34/nQ2pFBZWw1SIPtzC
NRn5OhFTzVW1SfMBeKi2d8SkGWgMb0W8CnJwUXtbAM95rZu7p+VJecHwtBjZ
qZ8/bzmfpLUlNamRQAy2COXjl7UX+w1eNzg/4nzUjvMRo39dE9H/bcvIB3aN
6x5OLCmTOi7SoEF2etnLY4I3KRlvED8T2ovgVTbaSUo9vtCOuOj+shnnxXNJ
ASOkn5ANOStrN9XU+sXEWevye0j5Jj2UZCNbdFfMK4joshcGmjtdaAOK21xJ
JsV9471GfKWGOjtYqDDm9chyYV4oTdf58YthSnbZGBDWOGZBeWiYRde5ZzIP
eUxGqd/2km9eCnL+Lk8v4/3L9j4ah0Wl0XdNRIF7wmc11cvcexLUr7dyKYFL
By6lSrbGmMFdz6G3hSA98iR0K+Ddf6LnGHoHp52eLHk7DlxVmfvUIYNzf46X
agQmuEaBDfcXPv1fyM98fwGz8s0KJlz3Liqrmc5MKVrbhCwn0StpEJs030qx
wI8EOjyI8N44VwFd2A05nvpXmlW70kE9tU1vmUDtuGr13HxRLlkPHB7pbee/
rCPIAPmPq1pmL4kdEbYCdmhtdIw46E945qNchaRmgDZkRvvT5OJsHTLH2qRA
fygv4/j+8hrZd72QRPTWwQU/T3MZyDr7pqlvU49V+x57QNbkFURAr281duiJ
zqAc/PH6h1rgsAJ9KUzeEw2kVTorlo01zHs7Enw7widUCK2M/hE5ivnsFw+6
seiXCP5G4lmj5iADSeH049tQcNoSJ2+b/Du5V80AG/gei/JgKVsz3dTAsxWp
Izm/mUO0sPg7qoCCIxwlnkxDezm6R9BJMeLrEhKC49B8UiKqXkbhAv8Yj7sc
OU/QaHbcKk2gmM6c3WU2ay5qVM6UuFKKxQe8que9TaC2cwy+kHjtua9GnZYT
wR6eCygSEgAidOcUGfvBdORD7NkXQ2SK+5XBzWKglbimbaLL9rsewDrF+wG0
du2nPgTMiM17Vclkfzx5H74xEMl4XuEPGGszmOeb/kh2fn85171uX0xTd1Cu
o8UogBx7HilAo2mfKANDsQUB9GCoWVjNY4lIGXBgSIqHH20tKHv0h7DKPgq5
zU01RRwN8eHh94n9dSKjljYRhNY34BBriKSHtP+Avfwyex7rflyMZUNkX14N
txqQKNfVCsGHKE5Yl6qsIwYIg5F4fA1N5dnD+jvtW1zgXWWy/ep5Gb+jBzEO
MhddfOndgq4DdaRsVGXy1aODdfLG2i5SKya15uXTMzxsS5875z2OR6RIGTOe
N96e2sOimIc+FbLFXKqEBSF3y7UyoEWK2u/sm5Uq7V3LCP19dCVA2S1KitEx
96Oe17W7G5YOzMUV/+OOwPGyl+rf2KwJzkXuMqRb9qITKhkY1ECU630Zq+in
ECKh/0kQsGYpAmWq+yDJ0PCR/S7O28sAPCY9I3dQCVAvplCx2G5puM6zjuuZ
zMvqoul1F65/fYz5kVX6Lp+aYaCjdjc8tT64+j5F5LgrDkEE3eFbHHHX7AuG
0IgGpT0cSKRD9siLZEakUBpcBYuIOBmFGx0jpBonXnolGyDGh+cX4VDj3LPv
yebQo5RKeZ1toz10K3ZtwflbkVdMA+xH1Jv0g8iHlw5ZKAhckTzdVQFacOgn
t0MaV6iTEi6Nifs1Q9lhfpIMYu1Yul3PnvjiOhrGPqz/rRZx81DT9gn0nAKH
61EBVqTHWJvHiTaubxD0aXs8aA/UFeXVuN1nN/yJlj2jZjgvhc4oTnWAVbAe
kJqtoaf34NUnqk7fl9hMiSqPidzle/aZ/prcbL+ArUrz8piYvTrGqM3pIQul
FM/PXjRqtt5PYmMgnFzqIK3lZPuzqVvy3Wl7PWDIf7YBSbccKG5zE87R+LI+
s020EUd83vaYa4Ijk8QZk+ztKQyyo24crhdYKG9D7KLhN30vUD687K3t7gXo
MVas70mhbiHnm7fLTgo75OeTElAzSCh7EXwpvTbKbgjwZaFIx8r+YYscgsU0
AUqZhxN37EyIa7ZVLb4x+lGkcLbOCQGPvEGIUSjhTJ3YNk/RHFVL64HD+s/k
i5Qdlirt99cV7U8G3/ckCaOc8sUbZLznnuPmpUopiOS/+/RraUcVlOOTuHwy
8pKwgiV6vnTWVDdYOiOI73UXAIC/VV8EUtDuM/CSQZPzJ+yFyykhO+Oqj5a/
2egphNtiQ+vLM+xPCldXi3ts2w295Whjld6irFtQIKq2sHzQLQANamFn/nyV
grxMBQeNZ3kU7zYU1iknxV4OsktC6Ec1ze52zouZVElLKIBeRQytzUV+uAhK
3lJVJllA0/G4sQ1zVcZHzkBAHmeR5wCtlqHk1Rum1bF4fFRqW+SdoLjyCyWQ
IvGdmrrEUfmp8ZwX0tK/0x0JqZ3CuexPg5SUzFioq+ZWfZnkhoYRpje1fBHq
oo61ZQyzgZFMLm7XRDDcbLv0DhkpcBvbN0Necvja8ayKyNUxcq1Ce3bJDu9k
lz6VrjMw1uEXhji0M10Z9FKNyQb7GpL8bsLsF8mWpZJ3ZfIyrwLcAzDTfPzb
qNxs0+B77WW2Vuj3cryAfqcbTyFs9WIYrNH2X3V5qxCzuNShuv19Ygx49Z+e
945UrZumJ5Frp2d3nUG86vkK+u44gOYffzPJwKvrHhZWIkh7LzI/gBCT+KBg
4c8/02yL4XjQNUYObsASScAoiSADBFttDukLQ4zBcnOTGb65EXjpv+hKCNX9
wmJhD4K5tWZjUL5ceWfvd7OPx/D0pmJKziMn5hhQFgeOrQrwtl03222oMAxf
RpPbh4N7Mty1+RKSYCSnJFeYULCniM0iw4ohA/zvGPHq9xTOxxJmgnSY2H+G
gz/uoJBHY0i4M1lyaiqJtd4XcKNxIGyVlxTKwSKQJyGANjVQgCHPhcKWR+RC
Lkj5GV//LZXBqSWlUNWDL9TQSEL9qdvFCzfmCEHzkamFKybfV/R53QvPSf2Z
o8G8PiqxMgCqLnpkbrW0e9XelriUsP/upKkM/oMvS3WgFa4Q9JnP2Qs0+9h5
JCs9T8WXjsbTnViIMrzlrNQMWXBqyt2NPR0zetaEZXrpO4FyfD9dCwUv/5OA
kwPksfX+SEz7QB6nJewgJ0NkEUrqxAaMdnNx6EjnZg3uVu+SNZDwZkfMn0h7
r6ZEmtSW6Q+u287AHcowxtYYuro6gKsyZ6G5i6Ht3nTgJ7Ur0K5yODh6WloY
tWEyBfyXge1ZA4GXn4jMY7sJbUcX86TC7C98V/30Sxo6zmFOHVN+vsvNMhQm
mP5MDoz+0R0V4gp6irzpC2RaE4UQg+NWMfJ0uP5w9U6No7ugZRa6yvSYIwU+
4Dlo7jHCyEXrpUM1BC1MflOS6w6myme24yrkhE6pNWjiNzPcX/a1jBNaKi4O
tYcreNAOqXwl7B8G6/JuakDpVFUZFKFYJxKbrYGSd+G1TRaevI8u/Hk49wK+
IfFQP4cnTDrXidRJ34gDojyBYVK44snodOG5aDEXpmJm3HcSYNu7x8OWtw9N
qyoaLU4ibllbdmxQoQHCY4xJjTOrdozB9zkDtB0fGR0i+eiwyPg7aLMhjv5v
wWT+4DDVLTyg5vzpQB219pfkIviQiilCG88y4gMKy0whJykg65MsomvtYDoy
5QZLy7QxMbqCMUgjhZRC8kV82DuXiUzK8XiPl71U5TerVAcF4CHAMLozhmrD
BeiF3ykAvw9UjUZQhF77LEhAYWrioEEPLi5CN1JWypnWeibuv4lnntVmudtQ
tG35hBJBmym7L9QBdVyXiSiseWvkwCOTRpAb8NwEHZ0qhRQz4QllmNX8LSkU
STmISOjonO40GS5fK4ohd4Crgf5jHHVik+K7JCKYDtbVaMryf4adRkk9FZn3
4OYjVNfU5PlWjvQxa42dbSW8YX7fW3Hkin55qzQUM8wTbyuhAeH8/MxMY8xX
Iepbr6QLONZjeojENGeTjOa7wuf91cEFeLys3xmoDoYMEPfKTnD1v06fbeQD
Ie/X4kZsU3E3DtvE5raULS78aUnwFqycdqmr8CUQfQJMes9xjl+ZFQ3LqHmZ
gDbzLN+1mDAN5U3wCuns/5R1gYMy88cUuvEAwR02rN4pR4Ln3XReFlNqhXKs
SxJwphwgzD51s29NTXyDwgjxo1vkUqYQ34QBgjzZWlDE2xeaXDd1nRk4KBaV
aB4ckEqlj48TKYO3dufSQTii/GA2NvGDU+3/pJgCC4Ta0+v85mpBFvuXWA88
9CDFnYnAltBJu7N7N/AudxSHWELBc2UPyVA/k4iB0U0rl9e1fM7dwzHCrjmO
FfsPEisf2OQOD/VPmY/XarYQ38AkniUsFSYYZ8vlhRQ8oqF3m/re2Z0HBLaA
pyp5oLlblgRMLUhgKqSg8IX4jX83JWMh85lN5keUOT8VRnhDQW4jgxGbgiSK
LXMyR8aXGkd5DSGizA9rcVKxWFiTl+a53auQjHF256EA0uL6nuvHUW9yH2fp
LJ9kG4AXo2CHkIJOgPzCA4cAf7kYDZ6+MNJOcts2Tyuhw9DYRrkEVoOC6IHG
cNLY7LHca/jjEtmYk7+JhKRzg1yL0VN4PhAyHxpAf1pkE4GrINkz3EESTc49
dRG4czwVa/B/HAy/jtcObuVEdHVpCQqR1O+PEs4mujQwyKgE3u078MIhD+zw
+xbvIlWAi4ZowAuknDg0DadOToIDHJov/q8geRa14I/VXlaD4CEOkxr2gxIK
68cf+Mw5Gj7n63aWdNoX6Zu9uTaEbC5H1pBbTO5uVac0syS1ZbFgFeKItS4l
BWsApGSa1zA9yEfk+dDDWCbdy+UdgvYLeKDJWtW2+BpkCGEGNdw1OYg/K4/m
5u4HHJn2oEu8ZU0TEFDC1sra4IFent/wO632uCBpGAEW9U0mgxeYzR+aWRk2
EB8SaQSLwxqofKMudP7CD/dMPsIID27zbUT0SIXJpqXG0xneT8uqBsUvaslJ
F/HrwzDsQRo4SAl3l2XI42oGunqDv19cGlAZWSG2agkNso39X41zXJ8gMyaX
3VIgL4aGtH5KCMLs/eAwkXqZEoF+Ow0yU2ubi30PNLENYWtrT2WJ01rzVQv0
yzv3Ttl+ghLDytk6i1A40id9QdbCTtvQeYS+D+QAFeIUjpK3US7fBRFDILrz
LeEwlj4Hh9kaoCg9ae/mH/+kGjwXKPYtRvIJXa027nEFEluNH4o7qO12uJoL
H7IPfXWhq6VNEvZctSC9Wq6nejBPzCCVNHUomL22bjK7pUpfwreJ+sBAOguw
r7+AMmhnWimqYUCApkjJhkqnDD+NTsrUcbSyFdZP4GetqwifDZ10eWzrxaHR
D2n6bu2vGpl3BXgAOwe20BAIsr08WBdi57dII6GjmF1WA4B7OjJRLf2YbHvv
m/FxZohjpcXhOGcbPV5i8lTf43XpIdQbYCDF1Cm+XrZWY15IQN+TGvcPXb21
3uNq6MAxQQndSXbmX5M2H+VBIWGqsqxI2DHOCyVsOrArjzNwDdJrvxqjzMka
33Hd5JdnSnEIFjeeLwbErNJkAvPhpBlqhDFcqHKlJjYZ9i2pLiwIcsIerUkj
6DEEWy2A48fu56p1m+hT0IKvIv2P+jaVl/cjxqm5DwMO6JQdNyI7QJls/iXJ
0VF0cOP2YbCzRXKL/q0quwUur5GTbxnFmju089fKAAhBqFADJfAuTFFnTj31
snivVMhTQyu+jYuQ0rZToSWhMJ7RhFMmF5ephPUWHRRFZAwwz71pNx0KJ7oz
SFqlXRoKLI80UyVBMtUDCjXCohYREidbQkSG4N0Kc1hAzrVkFX3avX/e3FjH
8RUGwwzyW0rlc1NS56Na8+5JOWCaEdviTFIIqxTtf3TFwHzshpyd6ScZGebz
1QLUdfH6yBp/iPqfM7Uz9C1oXuN3hAZN5CgbsTwssjZZc7gRPd/Zk8YAuWGS
AGJbkjDG3eNZmC1rab6lxSyCUabOrJeucB32kytU1+rZT5PlDJQxshm/AvTa
7nj/JL6vSKM4xsrnQdr3Tiq50TRVRwWAXD8Ki66EVO1c8mkoQJ4ECCVjaqV4
Y3FhSBqy6bwgTFl8FDLZklvaJIvxKeDka8/UGXcgm17Q2guDS056Ptg3TLvV
iVGQAL0FxgKMFk3Qokw36pkORjuXrsulgIDs5so2YG25B6W0hK71Icw5hiWH
jMkNa1W2i6CJTT+ACeBAQL3UTiqRK/y8Wyj8DcAKysIUH5C3/i21g2ZoMTsx
SWDUPvUVHpmS/4t6U4NumoqfbZWfugveiLwGpE+SMs0OOJPV635I/B2aFWOD
f4/S0ojsn0EPJROQdRfOpAvSsElEg5G05uJ4m6pLS6yM/xrA7RQhnKglzguc
+FCJ+XbYGwJadw9AaF41FGj+OD4w8L2vgCcVFGt7ahmtwu4VILNwT3Rp/O2i
JMzTCop8cfWdO1W8XyoOqhKpkIC1kDOjLVz54EvqVXPkyS9XBOa6XM3ImRjq
VnmF0ApFrVrqBkskh8LE9zM3A74MxglCdtLAu2jiN6+0Vc08mYLHt4Vi1e7A
fFWWplFypgl5eXLlIWyBJLvjLQrN6shf7M1SZvmbkuwhmynOUv7NV4NOvxPr
2P2HDDlss4jLJY+g8tJrCR+be/S/PdOutwMvWsWHTcEZ7mLk19Ot2U2dQm0Z
aohJNx72LvYAWOxcFrOHPKWy0NBCKyaRk29PvHrFktEZe7iwzeaKblUlQGgE
ee4UNXbdYHQpDnNyzVkjEzOOpnniia73SiV5CWq+mF88BEeUnPnDEGlXNoFh
ojXYS0DR6muIOyHp7je253ejSnxiJ41nWknmT3AAF8KaNbQ0hx+Mqo/aILom
7O2lSAMPEEx0qVEBEJZSrdUbRY2SKArZs0RtpEAXFMwzlppvpvEEeD6apypg
LMIbmaQWB67z7tpXEx8L1VIHXQhn78TwAL0Tf7CjA7+cfqy+zuwfRpxCdpqc
8mYhc5DeXFXeHrztaTja2+WQU0luFWzlcUSCLMeReqFfmsonPLJY9UEkshkp
orxI98mzXAaFO+tmEOBqK0JO/eiSLlivMEM5HNnzxtkpRleGXOi2EmcpWXfS
3SdElVsWmGZh4D4jiCTv/oqOo5e3eJDexco1u7gX/RQOoZaPo4bHuzXSUYMU
l1p1UKqtTUP/YYEpZ0yro3+LSuRFnAL8vKO/r3fuE4Pt384L+Ic3AR4AF74R
BvlLMNrVsgaL28uWf9SdtQi/XsgEE3Uznq/ZabwN2p/w0HTLHe/axS95Jd1Q
ljxhuGDe6U6NsLbM2O3q3cE4bkIQIxfbtBrr5D+BMGK1SXtyFWM4ZUWCcNm1
l4djpU2NwyDFwGXkTfRPAslGKue1I2uQga+rhh4lio79/4HzQTeeVRzHosGi
3BV0fQnPI7Zo/SPG9agy0VqRSBRpobx75S32hiTEfyR7SKfEP31q+TR9BceF
3egOMNSvRE8gPOSdYxCQh6Z9E2k2JNzIRwM/nRCUoq9Wi8+jEWOQ1gzWO9Et
TOElyg+e5bmlhc4gEwVFb5TwGNT0DpXFIBv1giHqCA/jXhiNobv8KyqPVYYo
0wpmMZsC6yXFiMP6UbSL3orZSPRFlew5UarYlJrq+oQWYYcWs7Og7nKx4U3/
DI3EnTJKOek8SxEB3F6xg5nioqlRSoJhAqYeum8CzzvaNSXGHkv//nUkJqKx
Y7B/q5+Hr8fpxxtN98SmuVEXq4JBRjFk41fDT+AoU5+rkSIrihBOQzkFXT1o
PjYTw75Jlc/3hh0oERp4yTgH50VekM2v9U9dUZI5gSRDhQqfSaVUvASoTM8N
/Aq6zMliaMvrxSQ7JcumJo58LHdUrJaKkRnUPDzUnWnwv+f+T3+dWxv5jZvk
CfqBsP1zusdd+dNInr16fsr5GsVtiQFhvuSdLc0HCbBb8OHO4Yg8QNFENt17
1RyDq9LzXVlDk7wm7l8HIYsaIQe97uiIjT/tm8d/v8Oq37PRg14/O59AhzeM
jhWH8OKvH+3buSqLQAudUZKbchNyDcc+Zr5XJZxD67AxkrPHbrEeKit3SnSn
9zZ4dBSDfgblJqWTX+2VR9rz24aE2f/G9Z+GdiRmemVdPnc0PJLA3v8VHdhA
B5MIc9Jg8y8nQMEr8s6H/V/OHK3/LFvfomyQTlAnF0CnLSf0Yqk8Vb2HD88n
67JLLuMqY0g1hbJuqm+RwxNKzkZuhAhYxzvB95OeCXTA0xaEcUMJu0pnm2q9
iyzFImdpdbyYxXTpvPbdids7lTWg1yaGD7qvpO/87szG0tFCWe0hPlDOVyNE
MP03xFn7DxwvpOZPAhy9D/3X4MNCRTXK3VIyWivRgMTPzCsvsRWCECWiC9SI
Y/T8yYgE3I4RznJrmYfGnwm7aoEnuzviW/Mei0A25JOfbXZMRrB7Iy4Xmh86
NVwzxNFin6WjUnRw5qZg84fGk5qToDbmePS73fF00ib8YKlwcc0adeuy928e
qJRuXUyA0+EqiOoLIqMwnGC/ETqhmph5GWQq3QXIiytjzYkoE1LmJlVYDWXm
zw9w2Mhoxj686V002QTLgyr6Le7iwfoXPe4bvKrJqSJ97M0XlkimXYN5GlRl
B/9aYC2IsjanHE4oLpNH+ttKQRYPlgawjDlAB1i80VOSbz4YzLvMrQQ9nxrD
EUuMC5Ut2/N+IIPSgsiHqgfUL6hYSg1qfUmbliMIafVhm1cegmC/EYx6I2cR
fV1ugn5dJofjV6Y5tEEcpeGbK7AS2sPoPoTOPmSuAcHvCJOPVfgO8H5ndy3H
d9TbOJBPj9NXCI3ADrciAA2nZdrdm0OMYiRVLQnAzR5Xi858rqSdzXa3Mh2Y
CrwfpDq6YKvtxHya9nKe1tEMw5YAiRQWBRRVk/VV0l/ams2I/9AhoYqmLBNe
xC6mW5l+3CbjkueR9kbvKzc0eOT7iyBgT+SccWp82kJcqeRtwJZgSSCD27hV
1hOWyRpF564Q2uogKXHqVqyfOiceA2D+m2fhUEgoFjAANFyVdfjA4BT3Xzgz
w38T2j7EiBZCioi0EAggh5LCacT+pw5s5xfku9RnetUd8TzcQySgKabG6Xsq
mSb0rYRtEV68THHQdnjt44awsOcMg7O3F5ayIcMeerD1/kt6eQFNWekTiICM
Pi2KZrGpZrr/JLMu8ZbIY0PN+h0JHtMPTNfDVbUFmANzmi8hWfKReQjp4ogY
EmdonYVMKSdamlv8h70YFguqlpZPS9CY0N225tJanL/yEGhucoeif2nZUZYm
Z7Xe7pDvj+/Y4FAXElWlky2nqSgmIzbTQeEyWewZvF/JGlOaGrtrlv9DBDk0
JKqm/UEWpSbINDLmTLmwNegyKFa0AEp7hWzaS7/VBq2kR1yRp11d5xJdMBmS
6+oYaHVUDWQw08c7hKamuR0qW009HHBDc9V4NJSQEgPtZUeG3qjfExCOpvkY
9kAItHIS/f+k2bFONmGxqAi+/AXBIDnAunqFfnlHuxQ9LmuZPNgg/cfneuWH
eSveA4+bnPl6UfqiVNFCbxBQHMAzMoAUIwJFri+z8vckHRXzDezgPwYAzQUn
Z00k51sGtIrnlAFs5GA+63GhwCiN9TPzGGWXZaE4BzBNfqk1u1DdUfA4bMEC
+f72ii3kW+SzOJFo3lDF10xXNkWPkMlzg9AMV03T8gqVq7Cyi0+3o8aujC3b
h3RsGL8RbTH/XQMzK54bCqlixzaEzGfpQ9K6yMjEjaVtp86gIQN53aeQoRxs
BWPBaVMCvpm3OQOtX3M3VNohV7j2RioGlbNlWr0hW4kLWH1ZiJ9RLzYgYWBl
pI5wsfeYQvk4BYrs4CuM5OBS817+fwIHEkCFh5KSO6GvGTtZIo5kSRdzcEye
3Rvv5mlThbEmDKAQVnE8ds9WGMFJG33hQdxOVAQkhY3mSChkvp/qL+eWm8+U
9Jy2nypzReMO42oPCiMAYEsRGZIMeArYbs4ypqeeWgycmf7sKyw+2eLOJH0y
c3tCFPM5ySfqEZaDvt2ZwrC2GwVGkPzokfgjSsRMlbWwWn9GHkLhGHopHgrG
j9zk42BhqzBpf/jOxmd9XjtWP8QljpMGDr/PE234gaLUznwEvn3V/oM0+wl/
iNbfLMDBaKtKMyyAwtBiuvQB6W+WURlZXn0KGXiqLn1AT/P3yV66UnaMORrd
pkY1rwh5BB1y8eHtmQ5Q+f6WfUHID3YeboD+2dLEV6egvx4Ph4kDFmHgJvCE
JyvnTzTEbBq1jgLwfnPCtzV/sfzbyBIHhpeMny3rhEWtKJ0LhgPX4zz5VPnE
Y+zCFXfe+QpAyDk96lBGg+S6btv7boLAo66LCGrxTxILkX1nkyIl4RAlqqDO
x61Y/ysHlhGdcfTiX2SmmQfgEC7zvyZkQbrR0N4HaaI3ll23sW4BG/sPV4lD
AeL7VXkrRBrS8UUlL5XB6JAhV+Q5JVTWNWSsStmh8Cd2lNZ6Ghip7+wLxNHr
OYnKdSY75Or9kdKZxtSI+BH//Qehs9yNUna8CyHE5uK0RzsYUoDAjCKwVlxM
VhJt4UhvIeTMrsNMkyoO3Eeem+u5AKi6Ut5nad9wPSNrD4PUnpblL41m+WGw
PulalNqiqBnoGRkhBFPuLCKePoRi8/EFlcv01Dn+Pll9i6QuAWek0hH8TtZm
KR7PqFoBwXeYADNC+07iCRnuE0JCC3YkNwRgRIuMKBGHYwbLE7+LCindjJL2
u8TFZP2E7sWsXM0vjELr4uhOgRPWKrBb0qvBdOa9gY2zIYl9FeKTOVHj7V+w
USUGstcPyLORhtJ5Umq6yOybwvw3V4R6CWjJmAi6Zgl5zwh5aFa+q4TKhpiR
UFW1ZAEJgJjEzQbryTZvFuH6eAejYytfoy4baStdgdouKIfDcr8mrQZTnyPZ
CFipa+tE1kB5LUfzJllnKKNz1MadfJqqK2IQ1dLYiWnTddnzjh48imzuWfVw
un8SyMAhCKRQwRmmpv/TWLmn5cYlItJQbFcGCFQzuUUAwsuVYFnHwhNnmXvd
QXA2lTcqXl52CVe57sh1o9Qxfr2DgsIIJa5xymZHguWtM2/5kySUFE5gZyf2
rh0hF9k//PvxG20bqSbZXip1flR2K95H36AyaDEAmDBmOw53PNGC7UZ/a1Cc
RFtgMFJ+jV/VZQwHTgCce9vEaZZ0CILjgBtpIk3kSbjrsjtsppJmzgQCxEoI
RLSEcdtsRiFiU3i8qKThPov9ar45VIEMqnvz9oMsad0QrZSbEywPKFiV4Yn6
IAuy6yH7ACSRjSnhtRV0sgAizMZfcE/4u994kuLsYCADSjMf+z41E1eynrNo
E51KOPDZcZQQ/+8+vPB15ETREKmPFhEAeAMSjw50iiMFiSONnc4v281oWfbJ
+ZJddbSAtPhmx5nTjb0zF+rDiFpav4TETwp4eEj3zqxZVS/xgFQ3NFKXNNwv
/5k8XRa0WjsjwXIo+fe+KEaocPdp7un/blrB5IYLKL4WrwczZyYrEJu/XNxo
dc8VAgroblI1YhnsYHjn6yFka4Yt40TxZBQwrOnOVk6Uu5aIqkhjnyJsFlhB
N3ZocdCLkcT7NMoyCDUr77FC2x3yQd578vEn4GuKsdMajWcQQD6J5+v1HLfO
N3mS0itbX2uZr7uPlPUYCDFQ6wIRYMY3j8mdD4ptqojGxtwaSqkPfz5aFbPP
Urikv9Gxw1Q+vJpkzOAx1oCuOieRVV4icsdZXjuz25zUNFSsUq/jT0zGnWgm
yJKNHKmTx3cKsJLAt5QPH9dYYs5A1yRnahe+bBpnk0vy73y2DGrHl5IgnsAp
CPY5NLD4xADzVCfEqM9b09t9V1fS6XV8L91HCWhmSzxxQdnqT5SDYXK5cMwI
djMObKP3TB2mbX2TCd8nqG6oZUR+6wa71n6Mctor+A66ZxJxgZtJ1UAU4jPi
3AT5oSSA9I0JdiH9Ho2y08p2XIWxpHifhPAxvci51o4mMmZjhbAC2C1ghMCN
fWIqAc7UjbqAvX1VGfkCjzTCRejGw2ypY1f2xICY4+Oz7y/wInALYlCqwe+s
fQ1AP/wyvGhK8ubfYNeSrrzE9JCN+D3oTLFJANiprfjO0odo0S8LsJQdm9GK
LuriOjACuYxoC7UQz4nfnW0UEbJ1ibzOZaHmYpzJiWXKcP9Jw22P4WNLNJd3
JRd3qnlDq7y0CM27NNWsE6vbbDAM3HJx8rqOLB9NjDOtxM1WAiziYyVi83T4
CYfk5at4UFL7H7ALHm/QLUG+RyYR43ZaprJAOkRudr0JY2Owx+2yIbkHX4vb
Fq3joZ2bG9Tq33O5EQEQsidCBjnFFlP0Y52NpRyQ5q7jRUSeE+gmmX+CDGwj
I790jLKD8z55OSo9qYY+RWLZDfF18et0ExdY2SLso5bvGDVkQ4X8HnoC2Lkp
0J2VjPOW57Yo9W4KCSIna6UJ5TGcSz4XWpz1HLIPNtnTsRBqXKZn7OBQ/4tv
iK5Kf5fDJLXF1c8Prw8/4JgNw+MwK1XZQKIOr2yATG34QZSRwC8uzn+s6JST
m9X48RkeevBYCz9tCzBMOHtkGA0ob++FbpOzITvh8fP3Tmcy8CDETjVdSoyJ
D9OwdhAKCu+Fhsz4weYpSbue1p+x1enkLwWzIylrQ3SJ5x8lzy8Uw/sg//yg
ucShrCz2HemhoXGhvjY1kX+MTrZjeESeAuXe/77F4et2+V24OiDkdKr1tdTn
b4dtyP4Ya2I/bOQDFISYvD68Amz1bVarFC+WLpzo8Lvy+ZblHJLqDDHlu840
wnBu1o6Kaa6gQhh2SLzZW3f3OVHIIKYWtKxNoQy79ivagTcX8UO30VEnJtcu
FmAzBB7Vlz781aV1vERCZswI0iDk1a8tpQEKJ/wDEEkI7khZ7rnJ6jJ/hpOj
4rrE3eb97n/q0eff7SUnZoM2DmzjIYoD5AooMkTMvvt8OKWx7DLeXpmIyy+a
AeFcjV3TixiKgC29/I8V3V6EhUjt3yrVOj3MIOXIdUZKUMbcC7RJXKiRdP9u
viVnI5hRKETUBoHAnnGipkVJU6nrPBkADTkeEJCRFsVExSAHFbNJJzqctF4D
lsjwTgWtkWbkn8+Y3TLzknijLQRgO1KqKaQokB/tGf27p3inWCOqtg7YmlDC
5j4vh4kdM5dqOwD94QEUr2J5u5Oa6iHhNN0fl0eLkk8VR0Grr+Xolmuup5tH
fsCrkTBTTeUZW+tQEqQsRvk+8btKc6qQ57tN7M+Kb+zE6871qO6y15xWRkZa
/Gb0ExaiVH9QfReEKTA33+xQUgZ6AMrUT8JByLCSm/C0MAiOuDsYSgd1haqh
7R4Pz7fY3HgOjjU99xotv9hpCd7YXxwmJhlEbKyxftBR/8nlcjxs5A8P0deO
CJxLt1JKnkIWKa6mB3TRsCWdhhpTFUYn9i/CG4jEfzLmRjXhjcnt/Mgah7s+
j6Dgr3w6zv1y2h3znl1IzmDXMreraVsXVCIzru2X1jTd3eCFCgD5u1O7nLUv
8CRlu7SM0Nx02EVRjCBLjbVFaeL+gGO7pjn/Cs8UjEEsAZ1tRM/TFGS3tAU+
SR97JklyFKCwwH6WAxiZeLq8j8eO3r/1MnrZQIwbcaDj+ZpLdqXqJEe5ButO
hMX1ahCyorq1MEsYkYsvjL13aPd1hkRGu7RWmf2g8roQt5UmZGfzbLM8V295
mZPNCWlGDg1BpAUaAika2b+z/xL92nmis8fwHM96VCtcoD0Dno6aO8v/CEOC
jOuAO8f8lPEnCPYwZGHiKGFlwQ7xiRc7RPHeCcvXpScgXzdA/DZccQNaoDEp
wj0TOVmaDvhSSDZGEtzs1KnLIIUzic2MptQ2bKl671nRoZSp0iTGr6BSW6E3
uhv3qDsPOZb8NAPGFuoszq2ciDGbVczqfpIm8AqWtlVwl1vj7wnBNT8X6cDC
/BQ//NCpCO32/U3t2ZNRfGAbFPgK0SZHcyPGpqH7VQAY9YCnwJLA9Dw77/5f
Kif5PQu68QARsHhQcLz5udYrV4lEaN93yGf1+cc4U2tVXcEd+IUf1O2Sz54+
3PSfYdVzTuLqGm26IpmGRR0b3xhVn8I0gydl+Gkk3VJ3duv9U5l/Db2Qm+Tj
wI1fPw1RmW8/q2jaaab12EY1r3deDZnL+JYXcrCBJHHdo4atzNPhDvYJBf2R
LaMZJrlKao2wWmACYUlsD15OP9SX8DRO1YeHPw+4C/mnxKZlI0o/C7KgCrCd
8uLF5WXt+BqXUO1e+y585RnU6vkT1pbmxmm0EvCJ/g7sYtdlUCobmoYKnTbc
4exgbfW+6y8G6XxArBz+iMYgy1wNmYdT+ab7faQmLHSQseOmCBO543v6UFa8
lgnTcq9ZtvH6XKYrtespauOBX8eNN2U0r2lh7zM/KOv2+2PVcRG4g69YcHzh
tUjSw2EuZl75yL6hQjjlXPq5Abx4Oh70fkCC06PZ9f37Nm2uVrfEnVMUO1md
irGnvRuIA1RQySTEfemh4cHZb5MiXdN5opuJx+UiOyVyI8sxqegI598B3afy
AQBigXsUo+pyiq0GO/0ZFzXKPNDpOsQ2e0yHN58HkaeGoSqcbZwnc6nNW8lq
iRoMNQUWI7gff81fyYJ2QsnBxVDtepxaPTSgcPbwkmezWjlydbFNc0L73orn
l6s0zEG8/9R2MaRn2mVEdah4Or4bCGVCCViT84I6/1Rwe0crf5zL2eRKFDUf
1/xoLgkqkX+Mx0AdLbXhg79eXRpWS1tM4Z+QJmps1kSSytZ3QMHs4zuUSgQM
FDLCRhCEbKIT4f/8+zWlHOYCUBL0zdSowvBfPFxaeuD8CYqOhdp/3WYbsU2G
uaEtgtGfbFmO69hGbmDfHc/voC6pwf5XtdfS4stbptThZO3sWfw2ALVH0NO0
+hXpbdRg3Q3383CU88gaE20E8giTGPIUMzhCugqaCvnmga5plpp19SFE5yW1
7PoMbSEC1HldVs48RAWUAOssPlF+yUj4cbAtKRSBghwMWxIu4s9We18kkOB3
7s8F/SK7+XgJ7qIc+rVoEr25/IbZNQUYEKdf49wqQhKveTJAYYBEUtbm5/sy
ogJOuCC0HXf8CbbG9oBS9NdiOK5ILqPsRnlE0kMBKHqyj9UKOJc+zPzi2a25
dA4ko9BgASlGrZCIdXBNIcxbF0ZoYbOUMbPrJoPryJvOb7O7U4ZY8PdklFRm
o2aY+eTLsdcwEMgIdjGdfayWpO8E2emGbpuG9LTyJLhG7BV6wQpmbY6CW406
RCI/ReMj6QN1JzNcXUc21NC0nD36Ebt7xHAt4FRdd8H44eOi/TJrutMyf8YO
zm/qxzGo1jXepPbFzl7GKY8H6hmQsywxKvrykXDCX350gjkxMQ0quWwOoJIp
wuDwchZenACcVOtH5Ll50V6l20Z4LX3JgMvUEguEHGO6os0CIc7Zl7KLTP1+
D8ahoQNR2sobD6E/H2RGUdyvDjz+bmlfAsY6Y0CWTKW6LuROChqAzqkUDm/r
vmgExQ67Ldf9qixPH397xjxqIDXq3LolQbhhRFGfS8W7CpI7G79oEdJ7MQGt
pJ8V+bbOaf4s63VopVJIjyUolpcat1opqJEzDvmY1MwOdyNkB6B9sqGsLdtz
pKWe/2wI0M7a93qL/O0fzW0WD1MotfGIg1O9vGrdA8LR5coVBp1fy9fBFlBS
kGPWN2cssHJYscV78vlw4S36oHh3TSDB8dHkJYQVeU0+n4gPl5vcXeG0PTIU
CbYSCjlRkx9kL4KHuFkXeWQBAd7scAQM4t4ohY8Q31UB40hB44Oyn5up1Z/2
5TDbSIb/e+2TxVoPaMrD1lct+e1PYsqB2hjaUoUfM7tubQWA5ZNt/4CLokJC
er7wriFPdwDPGyizC80kMVYcF98R+WVDIKZdqb+TO45cY5jk9257WgOK9E/Q
4Inr1nqdLK0TsF4p3n0qtZDiDx26oBq/pgwAo5Ei9mAOgiJfgf6dO4XqnWjY
OiSfTeH/j3jZXyfcrF2F1wiqlxSn9PDkVeoJ/U1Hdb2tHx9xZG20bFZPvGd2
E7A9A6XmYJKWIF8TzaVdhrZ202t0AMZxlvtPsPSKvw1Ayd7r8L2sB3RSSp8a
fHtjSoO0P8egSNN1WiXJ09oJqJGlcJtsH6XbLtNHWReuoOSGXJ7jiicYcT5J
5SAVoY9CDaBfuWM1w9cr2om7id/fjLr73et/1Ac4Mw4RKXGJ22GoNbYdmLEU
iWV6u6Hb9q1FmibpoVLj8eVAjPahz9W1yyAUto4UevwePMvVVjH8jGmlhOJw
PEVhwwrqYVoLX08XAcPXO1VMhapxjhTLCQHnR3prq8Bl5TTiuvhHNPmUr/O6
YH8D5WVKrjthXa5gdAVd71eKXGcc4T4nXhcLBsHnT+78KjPczq7QJ1l4ntGl
oIwyepV8Rp5nh40u6+5bLkTNssAKczhfDmmo1NXHtuzb9gewQZI/ON6HAjJE
KCJQ/NX18BRShvK6tA3SnTu5rZtMLQnsEIUcrRP57UmYMSCL7iZPUAc313jy
7gQQ/EuZDcuyAAPmEbyXpBOiULyP3om1EvTK4fn1CEh042jrnQKHSIeLgG1+
YxvE5AsuuONqOEzjhRPV3DUVxoZgd44JWHPibLLU7e2NZjI1K8FRjoP+hM6+
ibQYFblvDDQtJw3tc8bTHLsPRwpTv/xX/QKcmKFwsycrNjr0mMl/opA848vE
obcDdq4T7QdWQu/uJY7E60MMbOHkzaZ50aTsZSg1uN+GyjyC3M6X7vLcf25r
HdD5gIYiEq7CVe0AaOWOh2BPleWHaCrXaWJ0kq3RCGE9TqIl2wq94D1xIhtS
yVa3E/6H/4jcuT46+8aMvTkWHfN4f6t3oQNDAR/0Z2EeUKX9NU6aAQlgJgJo
2zh4jlChaKYA+DQB7Pk67cHMC6H2iQQslqTEu939UtzJmoT/qW9G4awb664v
KjPq4Gct12pL1u19p8kUxwcwQcjPESgvmbeBELDk3g7ZP7xEcQDgzWoUBkwa
lXKCJkYoDR6j+t1bujJ9Vqd7+E8MjnYyj7u/RRzk2Nh3vzhQ0+fm3/Cx0+hI
tCCSiLdeiA2ToHH7y8kYPa3Ir0BOLNTKHRfVOq3NFOoFNgcNu7kLiq8/4I7w
ncSIoHL3aRMwiVxo2TSImUmxS8mvTXXyciceCG4QBWL5SyOlR02AztoY0mR3
Dt7Hjx63/WIMdc1ysnKZQ54ahBurNyKtuVanxbuXdYqK5qv+ECSbPEFimBIC
ugPIerUimfbsHQ/7hwHUb7BaR/ie5HeWjQK0osETwgKNNKqYzzuHx7TwrV89
lhnhs4rr76e7akoQfVuBZjC/5qPkG4U/Etj8XJKrlLutukMUG+bjnA0HGLEm
rj7BHd0ZA0TRcKVkmKX1BjyKslY+JFGDS3f+uOr6EpD0dCi5ViSM9BPlxd8j
fi4c4FaFkS8WpwX9t6ZheZ5OmTC2vBRnFCIl93H53A8mn3GrwXT9M7ipuobA
mSB/p60HrEgALYUZktCzEynWofyvI2GxcoQUbdQwlGZMMWbYrIPwOoyvVmN2
1i2rL4ej08+o0Z+vH7XkmFmIgPcR6X7h74pnZPfcRhQIIIqQh/aTCjys1G2Y
CDuM+paNwOi8UPynApek1xjgF+iFugcl+cuSKzsOfrNdor6v8CE2u5Ykt4CI
oKEIXdBBiZ0qslkjpJkt6IqYdcUdTLVpzIcceh0Q59JATts1/WIwpVXrNm9v
8qe/b9XCvSuoRRVr1HsBofI+OSk0BLm6DTXtfl9o+4TpEezUE3HKmPbA/wcD
NZAFPUuS2vAGPpSscdb11OJ9MgzQD3kGuOl/13nwekV9Bm4FNhT5V/G6GJIZ
9x95hagWn9Pq9466ZkI980cwNb8HqeFX3u9cRqpfnj5JtR7TSGRp/pwM1HJq
Fx76BBVN/j0FEqjPnHgaIrbgyusMf+cceqfv6eBENn5ubXwOgc2/xKM4NO+3
R2LtYZ5JdRFkiD0MTkpQOBBQ5HE1g9J6WnUCULHBt+JXpfXbkAloVQ7eqkvI
3TVsAKwZ8lqMbuhOIlPW4zX2jbbPDbqeU6gR+0+HWXirqJjFc94v6Uz91/3t
RmqZcxzIReTcrcNLdqHBiVErPFLEREgq8C5WNeSur2Y2jA1B6KklY9IhpEaF
mP7qhP/zPSKTelbcMR0aWTYCpAOEXHSfySAp+ufe0yE4yVJTv0Flkfj796Gm
rxtwpfbR0SY3w9H8pcI5bG3WECRN9ZEMH2bBBQIVKvP+US9lFbteuZYOVV7J
2dKoMts1IJbya2hPHMjkrfU0cYgLNYznTC+0CYHAIxYDbN/WlmL9EiiCzfa4
KauhbpQdaR/UQfsILjCS1IRWhN7hLKlBwcdTv2rJ9GhgeJWXtqmzmoVz/mz+
a7dfVJaTNUUY2oXW+sSMfIl/d1wgCabqqlXdIg/I9Qpj/sa0DFfIqRQF5bFF
LPAhpA7Loz+1hKKaczGSTdyEAEjaWXqMXCkY2L7T7yCnDm/aZ4O46A/e7LEx
Vt9sWwDmPM3d3mklVQ2kIvCiozPMjV+nYkgkpwccDnC8vwmgtBHOiglT9pVn
FiieYpHkhWt0e66K+h07rinwQzMYpTf86Cbedf6zJ/vZL2rSnW+WKW0uNtcF
Mu152D6rTAsnZckUDz7a66GtImcV6AYYJZfR9z334k19ImWF1ij0Fo2qXtQf
6KzSebqqEjEC0LztT6V11rtteFSdvPiPI4KMRWqv804lIObRHpa0avaVrMrq
5JDa6XgIN0dQUE8f10h+Q9JhghxNCFhGuoEu7dHZmAr3Nu/Qq9i+5hpTvnMm
UFkTIIk6PPvsIDUJ2x/Dsd7bqfX6YByUIhWBQsNpp98TxPmxt4SWpbhlIkww
QcAF8WYKIMqPCoef6HAuzvai870S5vhyuc5/vI98GaXOHmld0Jw+X9ewBPen
zgi/TJ+VRQ6WmdO14BZ95Y9tWpEkHmgIXaQPX/Mui/rVQjqIwOWXWA4h9ESQ
ZV7EWqNQ6V9Z8QniEd1hIQ5weAXdbBCYLtCkQt0B+UmXmIjpkwT4T9I8/5XL
oyMt9tfogf5gWy2obG7YuCnwBv2QOcxHceZLsx33ei8tZqakIaqsvnTeKxz4
2hocYe6qXap1TJrlEJ0zNMKliDdZQnUeL3ZbDp8w9ijfFc7aGZ1gVF0F19sZ
dbKt3UZWwbw5i0SYnDbCzuthrR5eZjwUXyy0JipRCl1E//eEYRch73sR9ZEU
FdkS+0YWo5xRDCwuziDpeUkF3tp9mojteB3mU5zNqfU54YBhI0FnDEvEPNfX
/CkFvW5Teuk4ZqMd0NRzseBqGaPJ/XDUansLkr0HkpdM+ByEVNren0LOrrhm
Fp8NEPn4EjNKIr63BsKDr/UAebTrE3cR/wq34M7WG71faxs6mI35t+unuDml
nIhXg1kEipLqAmlbgFM6d+YdipTzc9/Pgf5TpiawASBHkUPde9Zi0KceWX8B
WKkf3OdZIAyaort8pQqLPlCOenlFRLT6qrK2Dax9++kE+28T60nSdJms3stY
UUoFFFNAMhBOj+8IB6Y1d5gNcab17sKCOgYqOn1527yL5RizoWynyNfnuR+t
qbhF3lm5hxA/a6kCpAD2pu871P0G4F3PVr7H/U40GmrclkWo5BN1tTnlqE6y
eW8WMwPhgIxxFKv0a+i58QgSr6f1L6Ki1KbT/hUjKXCjpaPi0LAyEoK1rg3Y
VZxJdJZrJlwrg41H4zvr40HDyoCLJCaWyhKEt1P3AIYy02rzaXotVSF18OU7
l0soSLHnv0tkojxsCieHdxtHfXxRE/+TXwqsVytIs6Dwp7Yw1dF6OzN62XlL
U3w2Z7wQOkIqdvp6ZzSjpWQ4c4qD/DUNL0ceUenb56NABsLZxhYWvoGpN40v
ZFGM3bo2pYqJrKmmVeOPCDhvHVqAHyCHfxat1d2gTm6UWXVlKmqV69LL6I7R
rOFktf+gNln/mdGblOMtKlDgyNy4MZfNWD3yyvhxD9Ld94tzsTWFrNIq10Hi
eECdgK3A784z8KmCKnFQwpJBn0TDTGD7IJW5kX5wmLlhp25tdhLfgUh6U5vF
mZXrGRgEDsIyniVcwIXkVFKJHCHEaoaW9B3bsSnX3AAsWr/9lG/s/5FCK+6T
ciZkcLoRtEJDu8QseajxDiQstqB8UL9f9PZZntyOy3+VH0hM0C0GmZdmikES
j+gbt6jwwUUNddH1EUQLeCRLnZsUqRIA++K/NlwW6df2/TEriYl0x3x2k+uX
kjt0XOjv1lhy0FqFxLVMYQa6+Bt5Ryo7RBUZ1/UeHWDBjOGLQhwd9VJmV343
AompgXHoDnPLShh/Uetv05JNJtaN2V8T18Oh8IvuM/NwqgBaPLhr7JcD8eFS
KZhVPcb2HOidWsDKtWPqVllT/1rUx79k/pkF45lN49hyYfnnabnid3r+t5pP
nXUdWgHWpE1/qaW7MvJTpznUGHHvkIWZenZWuBkDvCaxz8GcvT0H1iLUltEH
N7kl0ncWjqk/pJg2qJ1HLGAnMzqkSvieJRX6vYvNtio1llP/xzUgnEgljw8S
0eT5A3DgVS0RCJu8qpuQ0tv7zxkUDd3p0+9k0hBeDBAbDjIgwQPbN4cpdCsh
gUxDn371W4/cbxMsDqvxFA5t50/pJI+oYhkzVnCWogVHRIMWSBC/6IZcZK5X
+ScVeIxdFVD9YyOHbpfDPusrbp2pKKU4KMRV2NeLqt8tOiJ2gFtIO2Lf3rvp
CA5Gvk5aUbJqCOnpaaq1UXRuC3j0JmRwgCAfTgS09N/kMwtPEl1rltjP7kkz
aTb9pOLd5WkgewuRzmm3Vo8ijCdAY35BFtSUbEADTDv6Tqh5BZW5xwthZOct
9LSRKLT4rW7UHJivYYwsR3TXDBXqUqAvNA6xu8WmO+h8R9FAi8GxzZmUJYL1
HfhKPGlgmHKETXezXvbAuDJfw+Sdp3nmuZIoTD0BpfpkaJY0JRIXP/CLqQtU
j7vHr20gTr0+vAzMelYWt+OexaN+mDM/aWY38yiZiOzNWvYYPzrKDGjXX67h
Z1wv+ykWgB03OgcC6CqHrTxlIOUd902iOwyOG4tleyvVhGo6UMLucu6lclCy
9JIt6WW8Bl69CNcp6gIZMdfXAOR7ugTJ1gkOhZlgNLCBWqXLrcQfqRVotkP0
ueYzdXkrI0rsodPp0jUeW6otf7rB9H/VdhYN44fxbL/JfbFv/JgTXyaabYtb
yewvHojru1V7UW3bExKgIW7nyyLWknZqcMkcdvmwsR+SXrkMCvgZnIlB4JJF
6zx26roDkvElhuC0XeaNSLnohS5byio6AVbTMO8s85p/Q6WYgWG5KZXVG4ib
lq4/J2QDTHkMRD1TLGxNEjoASifB/euWFoWqKchk4+PQlL7rGgjenPAWGq2j
Bx57X0sR8ULD+o7gIumPVU+lebQOlrhA8wItUC+5bG7NkdZG0rS4TtgGX85S
ox0etq4Gwb6vqQQo7poeUdSdF3HO4fAKQ5nWmLFfFi11CmoNBJoyHWfbi6C+
h05/Y+w6T7jECXO8MGYUPXSm6dFAJH7xDbpJSoycy8dN4y/fknhsxzB8jcBB
+FeHzEXVOKOd3PY4RX4TlcXyeuY1wW4oPsKawdDmf1NDJcY2ps0B0biUknOz
x3B+OByGqDjK7Wfm0ien6Xp0u2QVF3maq3ZAA5xfjTh1AetUBNBsno0Mczv/
f+PDARNep5CfLVOg2r+ZpISrrLI/oAhVoM0j84GjQELO05AA0WpBDq7NF5kn
NaVAx4FR6gIqQu/FHcOvU/S4HUgvskzn+y0/5rjakAARvifCCiTibyexaa1U
/Gmq/FWmmSQWt0ICe29rjjATS+NnvC2x/TIsuhgu/VmWl6HVGJ/JEaFkxvbs
v4EEtVjOujJOHWxG8yFYIurZhRNSSC3nQ6VDzEw5CqPCdvr15dRcrr/+rc8k
h4bXmkz+ZQB6SpMdjVLvtBR5bt1iAL/t1EgvbwYeyXQ3DiVDaeHbDrWQVDOE
PNouARl+64fchH7g1zBI7OkqnZxtDsCnuNVo6L52bRS7cr9+dqRWtuxF41cf
OkmIpzYSf8oRaXX5q/ZC5eqlHCGbXgg7N6V0wp5GXrb2qvy4hqjRO6lh5UlY
qDnaVgxhsB+hjcy7dsTT/lx9kWCmbxD1fAQcZ7Ml+DNdOAxrUgmUYj+4XdKA
Xu5DqMTEF5Bqxgv0Ym1FMLx4OwHWiKilekX/XaYXeMWuSxCOAPR5IE07mJOx
TflF0s4AelUU6wozl8bFVfE4Ac3JQmz/ht/Iw4D7MZwq9qc1qejWo0qQyHQ8
smZn3YG4IvFRtikLECKRb+fYaZ1kiGwzzq51pwhCJYlkCL9jgCzJ+9FiZKXK
HDbE72v8sgXZzBZS+eYuossiF3w23qfBcSCt+ksVu9kbYBksQdCa0UoXCS6v
m2W+9DZnoPBWDAxqr/SrF1u77rGRHKgEKiGmIxIiMlfdk7ubSCK1Aenhm6pZ
6mv+Xxu4HDtChAhuJ8cAyTK/fC7jhtwPu4nUOueZBzQKx8DWym4bkRBtFHVf
IWdnfiK+xRvGVlsZxGU7/ks+cQuIriFCLONQv5G9PmGlKk/ZVuv2J8MldM9S
TlwC+SzU+2ejQvOupW6DxcuuMkUevrGZfZ6njdLzKcurVMj5KZnhhRH8W8W8
LNXQ0B6vtx1wrQegVtPavyyiVIJUNNmB0on5knLhY4ZvX6MJM1/XBQDpHhUs
o6FKjEx1Lx/3OGirO0/uMYUuq050bPcRXIZE9SdGhc1Xkt55rpGhyIduVk0Q
HE9oIB9Qbji0ynxb4skyjmvo56dlu6OfZrfwC6XTxDh7aErCBa0CU/d97FtH
Yh7ieTPsMJK2b6DOIX89A2IjyIJkmpfYJqn6eqO0E1Q8bDbVmjMPfte/vZv/
tjM0yxiRwPUhDG/tedjRtGuCQqSlAxxR5E8H8SGS/6nOeOedjP2SDPAa2P3T
Xt4BlJUKEdJFZwtRPxiohTXmiZgk7h/F9ociPFr83HBsaFr4MzPLw4CtCTPA
wtAwO664Zd3YH9njAFkcTgyvM9GM6D+zy2O9+OXt6PI+aMl5ilxLdjWFeINs
4/PBdISqroo4Yi0xvAXzenE4eTAxY4BY0Ly75Ao2GeUbNsIORzKsV+HNbIq+
NtaQlj0dRpUja5hzbyN1Spcv9nm9ikA3CDN7dPw1lRFR3/5w5VzZdn/CbbuU
rLjvItdKmmnIXdwRdn/VpuIo8Owh9QLoKcc5Kvz+RdWSNixkrrct6v7OHtfB
p2XsPgYPdT495U1WTwK8PqQ2pp7ixSlzaPjFuf8FddIidXIoZTdi7WAMb+N8
3pI3U4gQ9jQLo3XGI7+Z+VnKjo8XkSq4WlbYcifFUBeCi/wh0l6EYeMSH0TA
GgCgR4jD7Lgc6HLPZmkVsOQhaR5830+tmVnhY07avBEEFZG9FbP6Meadqx9u
94WdoQZgVlMZrwppBOeYGbmAHbQCx5qXTf8Og8/Ix90lj8MwOb86bZnxjZib
zFaPqokWIeoLbXRLgYiokZEKRzTtro7e0NE29pXVOlxqrbwr4bWbkKlr93m2
WHl9MB6gMJ1KD3etyOM4lAcYQt0mFwfJrk4I5KqQiitb/4bH8FMr0dLz5puT
1AGNOwHIxnDhmXD7tNm5r5uZgiDEftgD52xHMmkGSHHYrPtz64UElFqkm5R0
Ru9pt+qjeLl/5xb3d/TPxk8byOwU2hax6qzMVZucNw6W8K4fXygLy+nUzkHV
s2PxN85am7SwEQOhY5bfs5z5ZtBC46do60abhZtHkJaB2RDj7Ult3E7W2PKu
PB7m9qcqFrEbC8INuqtKfWDUESDLc+o/g6ob71m5PVgc4mb0IvwtMArhFB/4
vLl7zEfnXDd+4pPOE681e7ohnIyVzddxVfQi+ZRsh7f6Z2n8ks1Wb1BRWz9k
54BKL5yyKB0rOnH0SVB3We69IkRVjVnkR5gIY+rfQ2Nm+xoyVbgEweauj5MN
bCcmpETwE2Q3qNDjQbuo1WNV2/H3yMxUitUZqk+dAzy+ALdO7JdQf+QyomWw
FwBbdVz8AKIjTBfbgaeMDbIRzGdbROhlFSvnxIVQzfVv8v1ejEfzrU2OiVbN
mejGzvHnT9+6wOFav1OpFsGnhi8SSPKaO7nSfHFm1pqOvjpjVuo3Y4qHM77p
7N3J65AHBp5IP7oGhtlyJgyMVsOIsOYlQjrlGULzxNSjfMChZPlRvM+Con1P
BERDXMndAJJfajIfKkeFQyH4gP8af8whJrvy/in5S1dg6ZbiWHCzHmafj7Yd
CJs4SYa/+6EkKcB6LBSE45gRmWb3wbRYJbdM3nAbnibCOOBzmEqPuBh9K7b+
4Ouiomh6zGhjgnnGoxnbZua70nFsUZSm5CF6GVrOS+hXTk3Hyyqhl3WV8OYr
6jhkIhuHXDYXoDoYwnf7fjsOwM1pvZg5IR8h0WGQVSzsUHGG5le+aVk6w7Bt
X71k/JCusuwpbFu64SDwFKaJs/Zv4of8g0JQYwqf+bhis9LnUnSrMMLIBvV/
0eXQdtqwRDTJDlWkGAOn/aMe6W2fZ6msioTApK6rtnVoDdOvaJ4K+vAw0H4n
ZFjsRddoL/Xa0XNwdqygn2p5F8lQQEatjhVajC5RGrr3i7ba1Q+lXz1Y1LL+
nOsgZ41oGlA6rDVh1CXobitzX1SmRjPbBWpG6YJCqk7y6IAgtLnX+/C8wUQW
LggxbaGX3mHSio6r3o4bWib6xOHv5Rc3JRKTAfmMa4kLDhZO+q6XBhvQPIL8
WnT1s1411Uw/+Pl19grGGstlH3IbONukiVrtR2hLdmUQNk3PMyq6RTVRh5LM
ZIw2fhSJBKyw2SbTxZZudcrcR6Oc9rvQ6hnTFOjreAwQ4/XQ1LK2/6l/MqeP
mftTKlGUce5l2xG4V46nVZiuffkgRf/icoEIEF/URB+OBsGuxXmrPaLAPAfY
65SzmO7HBipsyXH7Bxl9afAlqTnt3bWkXveD5HT8tD7fVP+v9ZADogARtPnp
V6jBwTTx0yjSYGXvR0728Wi/wHdINq/l5kpBTgvEz5R2+h54YSjbn4lB12wz
/2zrARu6RjC1128Jo81PxHBxPgUN3YrY8OaE42PjZGmSgeaxeNRxuKOBUOhd
CJugx6hfDk1aGFc+fSk1OL0ozFbyOEZgPv2B6oITYXn3IJc2zkf8Jg2+i+xr
8TsN5T5H7xTqLcm8NVDZAvBjQ5HGdssPttg1uBP32poPcINQ3ocWiEVo/CF4
BkSO/Jibf0cFUOwE2tJ7hN2eUlCq9Q7DWKXQq6L7BhOFmwJrF/E8bFT+1bjO
8YdHrLjJN7tYU/VWJR6DYjCSVXROF2gWwP/f/uPeK/OtYyImnzRm44Bi9PQS
oHDjXcyH2tq1pg2CdjLD+3nKEWI0u1ntvaPO+HPTU1+1Vs+7hfrNznxB5CsT
GcvQB3F0e9w0qTRFPCDXem9HBSRhnOU9GWIyIoFdGpjM0/y4WC4KXMQFpjkl
KIpijMxtx63KuJSxEU1vg05Kj72M/CUDva5BOey28Gl5esSaswKc5WZnT5he
FMEh4e6LsHnIO15TNOLGU0rrq+S1YCJgtacZPwOkYluwqOxUJwL5+ynhaxQk
P7Ud//wEtIOfMjQFEFc0XnIy028uzvW1BNVwZz+GyziEnL8W5EQucBBcvCW8
ArQ2I+mKmx3aS9O/qbLu8XqA6fFVMDjHaIazNN+FgRty7zGXVRl3ptHKPyMP
WSouelTDcWTvV5PRpbFg7+cUASTaBUvsQGn5lUwjqsGH0SpIvnNObuAJC2wg
d4VlwK8DTEVuQXOEZ7nosEsPGpWg+IGfsVaG8T7tfUlC76CUldJN0k4kzJ/v
8uCWRiNomlnbGZkah1XwvWa+O7xBm4hBluizTAl1/18EASsD4292/ZJ2W6c9
7dj0WLw4hNf6t7LZdlDaCTl+apz4SL5VHD8hHrgoNK1STFyrhis71KMdZpy9
zSOuMoqmdn8FSkJqfY/EUmPsxTjEJFuOCEeBwPZRauKt4KLyaf+q3AWWlgeE
Y1arpH4P6cn174Z2oyb9fpuwpzc8AMFKJgDpMprAu1FXgae2OWFls17gFB0k
EVpe3DwtWwXt85AvN9Kf8hDQjfWP3tuDKT9ObbMWE6eOt93VLxeG5X8vYKJ6
P9G4aAxG7G4iR/5JY/dG13sHafbSljYgRhUP5C6tCeZbPHOgefMDXa0xb9tr
UoGZbx5SBmV4GYTrkHXYu4K6wfjCduF+Mbd57aFpdD5/SaXyoRvW4s4ZQMmD
/j+g8/962M9qAIf7BvEbrRMDEabzNNrXvaPPog537hppJi8NkExfo2CX0aC0
NJyf0dbOWmvOJTejqFlaEscGtWRFcexfabMlOAWnGuwXEe3IS5TW2mpdwmva
m5g6M8xk31BuDusyTxt2RgJuaKxw0reSbcOa43y9YKWVvuqiMag/Op9qdcsg
LP1YIEDZXOqpXn8HKc+mErumvVA1mgRjBxsmOYGVaGb0yEJMXFs/9EF2fYs5
D2ye2s6HYvM3l4MfnignxtQ4hwe/1vcxdwhX5sxxsUKL/RG1m26toIuiWSYN
r8H+oJAy9xfWLzR2fLQeo5pvJShw21CQ9Wupd7wwv7M0X6GPC7AmXqxu9P19
B5bjDKv6bHdq44XytcCCHwwAaI+qISWq7CrBhE0bYH7wvVyrKlMlMYLueHGj
wGNwJbh0S4hvD9IitXrg/EEyfUHEXXwNMsIa413RbOAbbh9fwMO3NtBIk+lW
8/d+MPUXMYEZIGTe9gO/M+cA5Ihgyz11Xh3YZZiSL5HPW4s0/sHNZuKOYdPG
8zUuViVbCAXNm1FUCW/VVY/wbOyAEIcXC6s06Xv0xxQ8REtu2pQ/kqiDFbcW
FG0oVxJFilrXToS1/hQgYFiRpW9+VhAMZT+6/YJ/ETRkGEi+Lvf2XrPFebJI
5RdZpz57hxhPD52MYuABxskvV+AeyjocbjrFN3kxNt9+NmPaVPaKsZJjVBqZ
Lx62PNb5E+KYdhDi6DiFQlCYMr9wRIUzNlrQlGBlPInsoOR3Z3upftMPpK2Y
IMM9m1RtNYSnkGSJr3bi14LdL8Iu6p2l9XRlM/IszVGc1zNdsECP2qcqme5Z
oa2oq52ZUoiTXYujmR1vGUcO12MeXP58/7A2SFnb186hcwlO6NriY2SIzifK
5QJ9qQXUfD0FQ6Wkn9sfmhE3qB8Kjy+0zNOpw0n6SjFrOf6Wr4cyRiLaLukg
J6wJLiEW2Mj9NEKkjnDnik68yAmwh7giO8qvL+Hr0/TrhZ9hHTuSNS45mzZY
Is9sxqdHX/rqQZF+/sjvv4IJ0a2khsQzICohTPvpqCNBKJx4xPSklNq/RWBk
dLVxbgI5xkSl15hEySRBvhV+BpQNL0K8HEy4SPAOMWSfUS5pvr+OHR5spwnz
0eOuYB9ewc6zTdkTqgEXF4DYspfLgR8iB3ET2n7R8Y+Wu/DHFlIzJe3LNX0A
Z3kgJuAOVGqno3Xihmm56qBjglToTmT79uVR8DqnkndyWlvt9MX8fgjXNET5
EOctHwX4mBwG/McvtyEwLZT7veei+O0RIscTxsyfe17+0D/YUc/l4uiy5Pf8
aB2oCNeU4eoj/+cl65illGbzk6oLsqPD0k0TV9SkkjvLCyHBNSD+u9SB6RBC
zNiI5kqX4baNjHvkcgOVmPj03gxdjdA06a9SsF0YEAdgVELqra5OqUm2/pq1
v9M45KNSCDmTqnVIsjWVqLDV17R/gs8GnyPMAv91sxQQ0PowLor5hSorLLzh
vIc14morwQ6e/oLEkWQLc+/cALLKgmgEzylq67C9j3ynNaGETHgfLCOdoSOV
+6/RbYqUuSZTSLFc3yYO8fdmdIG0xnqaj8X+QZhtCwkWqujzS9M0Xsbjp4qv
0pckqI99RTFh3WB1wdD3Xarnq9hysnX+MgMvXNO+Ny6W3rzs8sjZqr5RAcf4
QGita2MtldL9Sm+Eo8lA7ATmQJAYQAnhpR80dmLuc2YJm+25DNFx+gUIfI1A
k6KcDAgFKCUswSJ2sPhnJYdyQTRyhKecOb/8x6u6a1qP6gVl3pToUlnFUmRW
GDkxr/Aadsu83bh+5ik5O6Iv1uhAbxg2QPQEaVDUYFVXLMsb+urZC/fbw7WK
4BFkavUZemmxbuYiRNVvFMdW2ZBnNjdDlBCF46dP2zix0k+z8arSGGBghzye
AZ57nMmOrF4l/EZ80F4GPZP3LZ0Gtzw3GpK4NgDFNCeitWRSZu3nPJNTnrlt
yqB0c5XBX8xOsLu36L3duFxGFLJS1eUF2/IC+X3XQfeyYlTzNH0qWxwYXBnk
DYIFbSYVkdOGxfgq+dyjjIOJXkkf44Ryqnpg2xA3hqdeqoaS+AvjHL1wdUbx
MZJsQv0WwYzx/YqzE2ajSZR0Je6/kcYa3k9Eabtf0b+MZCBicPGPqmdsGQ03
dAmrK4Q2hGO05CXvUNfE1AwBC+Og/CbM0XRcIw2uRaeSM7tdw/S6A4+zqk9O
ULiVb0uf5s7VpR3WAt2tWLC0H0eyrJatpOonPxeS2UzbqHzqmaE7aJFDlxg8
/I3IliWVAy7QMOqPqfZBgQYhXvMWQdfhBKPrzhCDJy/n3wOKFlan45XfwkIQ
KFqo/oyIB2DRUhdt2+rCMwXqNCw4JiBvypKmlzXHi1BDD1QdgGO3+njMTSCf
asBRaKci0ZwexWD+X+pvQXf5vG6luyDXdNbBC6jh3VYD1St+oO0C+o1DAYjJ
RHDHHWsV//yot33ybkUMPIkTvrIwnjUCkNxkFs5kHZdGcx+llEd+M20r9+hF
1WyMNokG1x4ZpXTh97DFi7ooIFMi6GkaQiRsnVF/FOGXjzZ+Ti8/RSSvHaHc
FKnPmHkVXr/vmhqK8nV0Rj8RD1+46I/q0UB8F6eaFY+KSZP4MMn01yR826Pt
E9jBzUCmmn34QFoVXsiXPUNla4ppNMpeqL6p9uMYczvmcoGBvu7a58FsF6FC
jfb0dmpiSPC50K37k7IDHhyczifrTUutKETQvAoEEQ5X3DsyFj+MQBaXA8rG
JxdXHUmz+m/okJhzsi97veS75Aep0D7PMMqfmH/ZHDiy8Mu9ZiLGaKDLU60O
Oprq9BUeufYCJflHxh+c5HJs/V71E++gIjuibwpuUQebMhGvHIIp13sFBZ7U
mWed7qi4l8H3pKMw95bButzoqVLL0gsDjEDR3nX9oDCXxBxIgv2sxI5uH/CG
h5snqN/TI/bajyclxOk8ugQKaru+qjylu4LLhbgkFQ1EPtROlr7pA5TL+21d
V7Nc+6FWQC9Z2//nPbEP9hv/pcZuL1wTC2SxN7bJDkT+qdbWEIKfF0k9dVgw
xLHtx+OCArkUF3NbTVp/tNL4HP66fgyAdLGXR5QgkhZjoZ4OSVijOyZEbEVB
6wDu9qYr6tnq80R/kmya9cAO6S8IUV938EKY1PvPSvPm+CPsZ9csix7cpIIw
vwD9iv4iIl0l1f+CkURVQgnx6IrRu97PubCJxi5gAmf3ndEufPA8vDSARK2N
PPv9D3AdmOX1t8FHksos+PIf8wsor5FHaD5AzZAcHYb/e/OBfGYHqD1co3WK
w/Tdb7OoglFsj4sQNGMn+YrdI6j+hNLzuPzlWhKyqybtTNXMoWuiv+2oKg41
eL+Z2+DQEK+XGWQlIyqnRNFDwCCCQaBPskaNklqtbk7GlWFnf6mcc3KyuslO
GIBAVyLLlP40nPxDzoBtw6mYgSbK4dnzGH6eZDzZL2hmfnQo5eno+M0QcoP+
Z7l7JG2f3kPIsp5Jn1WVXDAgNepEoyDuYToMz2TPJlLuKVLZu+9z8tBr6M3o
0kXjYco8RHfXORdNnQRrXN3yrtsvsWd4FWLbk12Yd3dtJYTKzbRnBR1dKKg6
gg1R0P6GqLUoJYCfWzqUI1ud4k/Kr87apqDPEaOV56DprBx+6AwSolnb1JrQ
DNw310LicAUiipB1VeqHnCJtZwEZOmFmMTepfcSDSZh37NNeG2bRIRQmWHSb
dZhFD4Jwn8Rn6Mop7Kr5J8L+bafWvZVh0tPUg56yxDyJ4g92Djr4bqywoB8x
v8KyYdLgV1PGToqdD+UOmDiz0UPqYPRSyqpDRj0UHaf6SgSSFmQqQyYCux5U
i3SS+R+jmiVAOdIu72JUVnL7yvM17Oy35DMNS0x/Vfxy9F40RrwWJHW9VgfM
Y6JpN+YqK5UKBVGi66utTJEFsTggRDYsHWDuP+RuB7o6vXXS0Td4Bh5fTL7S
BtbG7E0Bjs8pyPXBfI//3M4x9eL/oZM5K31HXeixcMglTa1lmKfBUUKAi28s
i+OXCxONG7dt8y0B5Ad8fEah8dXpPPR9QLOyKEynQIFgqQISVM4GhJa+rPKD
NxtyKbS69jtIzaB4yb9JwsOL1uRCkT2mVHAb1tMt62ltnimTwl1gw7C56o+w
5CpGMS475hoAUkAFvhIvYxcRLV0zPWDwD25zJp2eepDFHg8jDr931A4AI9iI
rePDl4ArXjOU9v9iDDR9Z3by5rjuRKu7qw5OxTuMgM9fy8gQZb6Pj6SGYqTI
1wxk+skG4BEy3UEHVbqoIJ3E+2CGzpFne5vCkGB+RfupKYFB1ab/Nc5wp4e1
Z5/T2bQihnh/qEPN1sAnahtsMEcHkLOrdFlWlgfkJZ9ZexyE8WisKKWmRLz3
14gCKPe4Dvwr4/GBmR0+sVCSWDL8WlmI+m5ZnbmUTLrF47AWVQLm45xhgxzw
p3xibNt9PudVUrf1W4pR3NCVew5VmCUieUCSL0z7HtkBSR3K55o/Kgqbu9ln
hiQ9gH6t3esY69ki0VB7ixgNEEsSreseIqoQSPNihfXi/vn/GA63fkl0AyLz
hWvJ0Qo5ftubWc2FpZT8ewlzNjIrhyE81g5Vhy9vX2NndeT2/jTY2cFwMA+T
twegZ7cHPcJE89YpQN/V+rBsURCj6MSJ22N4h2nv9/RP2PUa7vXYB3ev6xlO
VWXoVTkSFAtmjQUgHpAlCXbQZh4dD02eION/OBJ0rPtjtjlBukxpx3WlRvZo
/ZHmXMFLRV8LnYVZr7/O/eWSp2oRYYKY0eFlFGr+dZtofClKp886CVk4nXcm
6535ko00ev3Wsr3yH8N50dXrs1IUrHM8cV0g3mHFIUs1hjKy0eDI0kIuXmNj
2+HbkjaiSsJOHHCx5Q/HvoV3b0OuWonQS+ax25OophhLLxUWiBn1MFPLirdd
JARskGCg3twPl+ALDtniOVaQLfhjS4IMvGNAbL6038XZbz/EyaNmZjMETmdu
7znWeUX9KHFIhHvYg0/rfv+UCnaw/8E6zI8bwrYdiDMNeiCvQWIHjlFQpJmu
lzigzJtPngkbVBe6ShsJtoceak6ajj3UgqvBto767UkxvS5RKWsts/aJK86k
hMvN/3fJsiEXG+NtfdfwDuM6jHrhftDvAfqDeAkd1aDtaL1F6rVLQ0PCCkqb
zB8SzTIfu+MtJD9HxJvQvjBjyBnAIKEhY9UbSplt1PP3XpqNCHxgH2UgCLxl
//lkc0FGBWy8hcHzS4rsmqYmeFPs9IxtCROuzl8Ev9aBIADY7XwWxcah05JP
TiTJw25jorhRVfhWBVdVVvtdmlF10sA6dYHh02L50AZcZmx4JY44CaOq2cbd
uWr62253cD0JHPfLl9ApMNjsQL4rcVyoFOZpm8naRAEUnl1CH/qcXvoC75CL
94J/a9gQcdG1S/g+15sijHnllK546Dq9Z+Im/2UkD4pW6NaJ6gvLPSiJ9QOQ
go8vy7TKMA+aC7oLtJU8cmGNNhYlxbHURtzidjOsmSNisjYMUCCYbksv6l20
KKOrxNg0YfOmxDg6QSO+naypdm4a4oKJsgL4IWUHqKtwhwPvE1dvZHTXHM82
hfAToKx01mR9XRpxxvKy2mfr4i9oJNo9LW7lq2+n+3SnQOp1TnQ053IfC2K8
w1oAiKi4acXu/kOoMLmkLcrQicWNSKqBHYVFflUgcZq8BZD3nrLpCMLYKCSM
X6zx5MLLycytpDK//N4kM0519itYmnnsBkZUuJuz0acNVhQfwu9zljCC/Ycs
lUceA48V+fSOjQ2PFFv0hdRRTatLnWlIqCLRTOxfQYnaNmi8RaKwxrRdfluW
uGRJ3aXyz+E2Pvyl+0fZMSjv1fuPGDb6z/9R/QdLaiPAKJWMoXGThKGmhGL7
fWgLFd3k60+H0sWI4D0EVf92VifVvJ3+p4RYxOSELshLM9aDVtc0UuefRVHT
tthMqOnHxRLtxZBNxM4iijD8X/hq8reTMIY+mFIEel1q/EYDEl5zpr7emYkC
hNv4nUAMSSUzgosVv/hMAl5+XtJf9h3BDODzd8XatKtoJJhA3QUbVF5r/OYo
SzBkPiYNPitoXWNyILBr5Bf4B7qPC4rVzSV3cc2487j+I6HW7kHBFm+2Shc/
SDdbh+RIhkaAPIokkDh7ipfSGcvkbWGa3Co6gA6NQBffV+8XODOB0hhJjV0J
61L+DNdyAgrNCdsxbn2H1OfoKZFrSvW8Kops6XXVLHDxSR8yxub8eXcSx8b7
WYnEsG5BAB37q/N766ZvW29IRaOQIAJ+AvDeHin4um7X7X0dJs+tAsxtD1D9
vMKSZh1fVi+BLIhybZimg38HHdmi2cU52Ju5A/qnXV+JW9bUu6q6hDcRVG+d
jj6OYKJGcPdqrzoG/TWQBVqcLXe85eZcr9QH4OiHFXwNfKIqxgv6v5oWDf9N
8HvZuw+jy6u4jCvetICZz6sh7DEazGzYXSHp8isch8eidf0Bg5ksnPoXFzp3
oPhfpC/z3cfPbkqOJhHjkhSRkXhMADoW+kvZyaZISjl2s7lXa7NoQIM6kJcY
1pYKS8RXlG6saLLJFwTB0H4VrXjeqoE56NLk4bGsX4PfDtr6UWqGUJm4BQNu
m3cRNtSpuiJClyKQGIqQvI1L6JUSmHYFI+oXk65/5JWLLgnqiwMwc0OiLswB
s17zsH9wbxyETD36sw/vsQZ6q9MSE1AH081c9sL3UJ3qm2sVG0+sMBb/g2oL
qcf8Noml+1mtvpHhku6KLzphEaJEtPjYF5sMPisrKfETHo9FzQ4ub2TexfDo
Ob1b5xUEesEhBZDLQz7/4c/TpkEqUk7vdabRt2O3dFnCOYaVLG0qI/qkzJ81
QLf5RQrTDl7n3NNt03Nz8f69d1LCFCKOycOuHHxXEqiJUVQUuUawiiKoRxn/
wrrdeQmGbkU+juhXoprEAx7i2M/aY5xTvDpj7QXzedLTux19MFAckVAQc2ON
o3sc9oUQbsZWKicH/Uou/2XpnF0INYGJyLgClvlgYf2H1qPTPTXXqLJBOdL9
hAZgPiA1KjEM1iVAV4SgeXpUTQDXhwW3dwZEQo1YbySoqDhflbaQADoUD4hO
K5qlVF4A65UFafFtWssj8RjP7WI7PewKDogU41AhzT1A06P3u4X8Myv+NL6K
mn2VMu6lhQxMffHlMQw38YX5/g+ReKaZugFADl83H812FFFdAds+100HO1CH
m9c8osorC0+LO93R1sg7j4rZnDIbkFpc6rFrBgGtMSanwV0Erhf7F7DofH1Z
nluPfxwp5K4i+Ds4mZ2xNwwpZGtQNOFRicI537jVB92sGtoxUE+1Sl8Gq4jR
Ypty3HsBZ7qNBf8Lk+2BQIznb/TIn6AjhKMBLJz/EAu2n80XSPEmrD8szapJ
6ynFQrTVdus4YAJpdtIWyzfdGUN5sSI+5E6+2yWlvcWXzomxprBIkqtFSUE6
fLoypqcBjyLbFcBYoT9qt6tfcudp40sUheAmoMjqOZTG0XbMNjMHs7QfcMbW
sGewKJlYq9FszFAox9cXjQb+aZUNaN27dZPDZrvctOUKNJBe4v3dLw2Lb3oi
kv5H+UNAjwe3yL91kb912J/BOkhM+kq4N7N9iUgjXAOJAsmqA/dcqu5eQreO
3yzy9SKT8vsDW8G8KOfCnv+LvSZ0lNIIjnSaUH4/JTXGXOevsEv+4GNpE3JD
/74J5ROh/hjoRxYtApmtI9K9WhOnWCjKI+GoZawgaU6GAee5ho7Wmxole+5y
HDHolJBhyRylU82RuO0GgCkToYyRqTIvfzNMn5xs0JFO7tjbEf6fhrVKqfUH
kENwJRJ0ur6TIekgDtop1hRVUsfqBonrlWzIifc3jtZhjrQMv1aYlM6CbZvj
f41AwzDXUZB3k/udVyzTgG9FSNBqB/eZJ5BmooaiN7OVuZUAan3nyE0jaFM3
B4eWz5I5qwC8K9nyxZdWxX8OQKsSHgtUrxk4l3ScV6fUZGD39FxIjohejOPJ
5TeeqlxDj7iOYEsTJ7/bUeZrj0FWDEuwXQYE0prsT/iEzB4aIRNCS8PRBjZu
1fbHIjMLC4iZxrhY/lgJpsMz2L5E3I4r/q8HFefhqokomlP5Dhj+E4DiOJRx
AQsLKnCOPCh00c+xyGIE8Jvl6rJ6ZCyiYFGHShOr1HF4ck5aSaKI26nTAtqT
IFFkT2KgDeau0T8KC1DAEreRyXhedQb0mnnJjJodygyuj/wI0u0PBcRQyqNc
LAkGfaeKrWOqNyFiSdlMFufesCFHMqlF3L0CmkdB8nMAZhPXN9hbXKhmHIqf
v//0mQzXMd5vTvVpAI0rrlqyQxRwsb8MF5xcGB0DfWrXDq3P1Vd9y0Dt4Z44
Nnnfe9lqhNoTolPWVsY1BYXyKbjblzUyqkTKVysVyyg3YrirOU0m+pp2j0ZJ
z/k8AkjBul+MWkrtxnY8vvjXagm06nbilTU0miokGeNjXeHqZxs3Nwifcwbq
yaN0YzLpeAlzxgi7iR1U8qZJ1M1+L6o5b4UfJzHv2+G7MwVTzcj/SSQR/J5/
LT4MQd0KkOxvZ5ZvwnSsGgduTwXsi1UoWiFXLwVDxsCw84P4SHjX38xvKgQe
xk0YbVL3bnzcnq9v0D98VYGrLHLWsgipNbVojmh+369PsY/EEgBl+2qTmzZS
OORGYmew601C+1clrMlKRHpM9CGUpmp9ELApux2pQFuhYd+vXh6PPNUdACxo
2VPcShv37WdmlDPw/d1yKAzrO/xblEDz+UKAdMKYRnuiOGOpjsWbZNngcZs3
myT14coAc8BVmPI+lbhKN0rwFT2tSrLV7TOhrS0dsTODCcy3OPBpI3Kf336y
xDtcK3w/GkG+TT74uYHwOH/zc/IIWuGh80T2KVmLK464O3EiKAm8BKk3cLSb
+1PIUcEIixhz6jT2sng+uFHcaR60115b0+T4NjW8Ebavz4VL8XY8JzANU4Ci
FHTtWcgUD7nUIjHO8VqVwLkzFjqAq/6kwlvn+56F7TIsmd0Y/AhgPH/KPcTE
8/2NqECQhvDWmx7pSW0aj4i3zvuxujRgZYi0pn8zebh2r9THA2d/PtN797uZ
Q5sJ7w5WSvL4uNR+Xbrmk5h7l215iEY5hXgyG1Eybijo4fBVicq4Nflpf1nY
1SALlbLhCSDNbVPMBPL/MVD+AWeZnYCbk13W6NaRFcVO0RIeM7dNDQUauD8F
Ethnp+W5nRikUlnorqFGTJ4ospeH7jJXvWltwdHi4/v/Fzr2F+sJWcwBPJOu
/MytsY1/NwzxxrS8A+r7yb8cJ4Pfo6PyczCfseGBhcdANmZKOitzMjIwzpYH
O/d5RTlPXLMpLBKwgnOZppb5qqqmnFEifGY+2cA4b1+l0IYpSCIKYNpf5vox
msZPcxf2UErrtxpCIpSoOWuAbfeq/aJgsiMCvkxUn1Ih6AgRLsr3bXoNW4yJ
ZDg51cbkdOEyi+dfeeuj1t23W3dqZ0jUegvVP0rA2pvGl5TCEU0us6P4J1ZC
hg3YJj18nT+lsoteRg9RKe5f8Y6+BQVUAqzppC8dqef/GF0SRclPSvEOLhQz
Gn3W0la0M8tMXxTr5y72Ynfpl7qzV6+J2hZxnKy8XrWvmY6loeF8NwgG2pdm
gpWa/GF2nEsb2VehqBbsczZ1sJ1oT5HY2cl6NOAm6iB/IQ//ZMkf61ytC3e5
GS4eVi16kskHfAQhsusukyruLKlfQQPhSArOz5KO/WwryIOkJLn1XrGsKCt3
oX67fSMzA6qIX4J7xgtj/sCAp//p8nYgYq/DZsr8fcNtJwfg782K2U/t+UT8
oHBsI5gyMsbKGWoZB3ywdz8VwmHh2EoPbwbsCmO2o/j2mnXXwGWx/yLoVnfv
5QkH2992h4WdxKnlbYmUilIwQoZfCsP0k2wTUt8gIbF00sQi8jC8Wa11O6/e
N10McpRIBIn28DNhQu/Z5j7GHmA9uh32v/fASLr1TwSWjglwxZEuRe11itAf
DLr6bW2mkMKZyD+yBseasBOtcivJcyv4roRdgVC3hIEkQuWK86C5pbMOefcZ
aenXnnSbGczSbIH8BzNpdLQ4qQyffOd6cModzIF1WJAbq84Ds1tIMmIWueq/
Hi40ZAhs8De8uBQWAWuSEVQOOLWOLSx2HE+4ogDN1lqAEc2qtWl9lJwEbOa9
41CdFToOGNHbxF6wqFOlZSv7Q1LDfPTG8P6PwuSIWFVaU7lUGmfLZv1rgFeI
Qt8jqpKEgrgPJEloIy8dzZGFHNHEfWMwJfZPYYvAtGuJ9dqssGyiZppmedJ2
vkUKVtXCCDr4dpOrrmMyHOqs8lVFGP7gyYtYC4452BLH0kOd4IeOGZ8G0paH
CrFtUJrnT+yQCMorKtNFLQezB93UA/cU9tGeUh7JJ9KuJGovRjFPk+NmdQnb
R2v8gh5LWG2lTz2qwpIDEV6wQOQjjRiKWXtyGUEPOeKTOdu55aEE0ZtV5TOU
ZyA87GteV8dz6/nldDlNdUXU03FucbeWIBST9+brAUqwzJ1WYrMEDp5drdzh
53D6Ya9IP7tVgNJD6QsssVMetuO7fP/1PYK7UGjBCkqe+SZY0k+4L1LRdM8e
1y+ZWqF94PrzdjHcefkuVpjqeWGhqg4G+CX6ZwIVWSCxMiqHybsdjjw6QI2d
AyzS1/ZKhoKEnubVLtAqUPzi193GXSPsvPLI1kijcr6J5TxkmE/uiTgDiBsL
chnl5gQbwJ2B2fXjoKR2qClmtrz2S2Q8GRumj01F2QQdsKb+mv6dq1Ty7l8D
wshXg3AvxbVW1nwQZAo2+CBuhe/kZqcFTfDgcoGoWOUqqIr38GJVcxm9c5tY
fTWViLb7FqTpi2Yq1rOE0MCoi48qkHqRFruODAAOhtOnZpG+R6FxoEZhK6te
R5ltZYPDsf6qPGiKLbgtW0rHRgZ3/tBGWDBnUuNkTaQErJXZUMzt0U1WGKpn
k+7C7uHv+cXi9/hQbh6PS+tNbG+0MAAc8yTkqvzCTWp0UfaD7w6vEPi9s1Ts
tC6k2pRtQCCkP7koViubm7TmpUHmIacp9TbsIO1Ne1iTo+LkyVaJotbOh1Oq
o9LgXdQgqYfAbjq36qJiz8R4ZNDqheb5N8CQ5dll8on40nzOOI+UtwvXowmN
/khl59g3YldHbZ5dLs1puJ7mGsvB0Qz3uvbW83hdN471MUdlWlWIBkOK6Ei9
FqbyaaK1rdWOk/Yl/o0w+eUfqLwi7mgTISakiu96OmJc58HpAWJgk0iLyvJe
VFxdM7a8V81ehkXhvVphA+z+0wgSuaXHeVfGNp/o8nJoB5WUBZHtmjPJIVsp
YqOOyEafRq02y2xWI6f8QX9MYM0qGxsH/VlY1kkcW+SMxSqrZ1/XQs7uEDhi
BY2Kh0DMqTtcxHgBZwxAA8F7+sgsHQC5+fShuep1bB59PyuFJnVWT4dYhlVh
0+ejSsuxKw0UXUja8jjatPfbGCEbpwwN5oTieEg0VsK2Qlzz5ILhJMFBwlLf
QirkP8S8kYtiNKCLDJM08EZiDTl4K2M7ZBjKNHkDWmBHOwAciOmRVzwyU25u
V0pb4jur1220UPTw09tYaOuTbThDklg6ZbIW2CrX8Z8Yxh7fWeOL58FpTZyB
llXAMOB0S/WaITdpyk30m0RwhXZOLbuagGVgW3nzv3fNmGko7y6NfJS0LRAP
mM/tLNaN84NX71IF7uYMzETl6fazd5LexjJv3bc6c3y+P1YXxsSte54Ga9Jf
A6c6Sp4BF+iZrwC1ClP/oTC2hPrVmRwJe5u8tB4F3hwwFUDKMA1JiIPjcy37
oVMprju5pccs2q43WFF/cuVl258aVKRWMS4OM02Ohr+oZ2XwsIqQG6irXNDe
s2Mojdohi1xMSwCTrWChW3/e9GR3ybosR5JhwgT3PR+L9FFDmth1Zb/pnyNT
JO3TiswBjG9PKwvDFwbRhPzO7KsGqDie84ix3WSjtOnKFIykOBvVd76gBott
RQ+VVvCG4/wxBcyL5DcQCoKzdMqt12y4uiKqo1D2lTxxy1vAsw77+OP5Ki/l
5rmhLoiYApXjPLTgoDoJAl3nqc6CER3Nx9TI+Jiq3yVKQs9cSHIsnAapbFwg
Qz9/KebEZxkygNOe8cjUbdpO/vFoQ0gnMDd1A6KaFTOKn617B5bCk2U2wAb1
Ma57FESnaDG7PTA3mBQflj0jhbGS4fr7+TguFMm64BXerC3/ho9gY6WqsTL+
uniJVenAtYRapQdaTcu+FXK4wUNiSVTR5TZcZcWnqoz+ZNtfMVUw+e9xdHaa
+kwgPCzog5Rbs/MGwlAfYSDloVprvICtyp1saUIbvSPhwhTUfVQf0CltPi77
xm/LuLvVdCemdT8rkiu6a0nvYB4OaqPI2JvjcdwJsnvC5XQvRx4hSeZbE4n+
6wiHeWV1Ng3hZ0hZnk82FOMB8UImtz/UeJuw12PBWN6hPBIbO2fHgXk64MBW
Dzv629Euwq4+FNJvhVCKr0lenRlmJTBIQbQtGgVDlw/rV2KEKuW1eFKdsrra
8KoQ3omYGRZhN8DpsUVzvqBg0fYj4fjavcvD2gJO6VpDKYECOnoY1z4Dln0t
CRLIbrAFNBBFYSNKlly19qSYsb+Zz7kly3PeVk7lTPalmCSCAah3zAMIbJap
C6DiEbAtzqWguo726XXQV8ema923PwjH0OwGFGoPY4sbbwJaZOeTmolhY4xC
pe3Jvkk6Rtl5/KyxXW5pO9h6U3LjQkZnYrrKy3FNMECF5obGXTJPpZaZq4EZ
xNM/qpCjAQEnvVJEHQt8XXhgH3bjyVtP3aXN5InX/DKQ1YfJmAqqJoct+3jr
MD+D/RSNnZtlSzEMYeIK0Yd2/hkHG7z3QkGj2pIA/k+o+aGFM9rN4pt6c1M6
N7biGqGdlZJprc1lq3QlxS/BP7e05EAz2wwgyRfWTEnpbcw6UrDrEciC/wNt
F5QVzi7j0U4ZTcGnoFD19JaVEoCbqHLgMSH+ECuUk74h4IkiE3a7uQDinvdR
MYvOM6AXxGLv+0juNUrUGc/MEvP1oUp5sJtLRxGzcZ+Sz9QTQ/GUzgph2tCf
QEtMdp9kQWmcxCcCVIDFyE4mIIq0xfQaaVxZycd/SQ2pMOQ+BYlmtHxj5k/I
Y8fAr9lDagzIIXpcF2CcWZBnzSKC6CiQHRtYcIyVZTfEZg9JRXT8Fk9Q3cIt
ujEHzwhuxHwxi0eCUVBRRl40QPkV+cLMTkVqrPj75DSIBVuzmIIrw0+2caYU
UDJQV3UbvdC+YqARWeIO+93GeV31ApDRyuPDMLPN01NtDxZ3AkrO/LeHxMdS
FtHWZaNyB3eEzRtC4pvvr58lUd68vQDUEmCFzJIvYQcpzruaIBhGGskkhzxE
WBaiNQ62z0lA5rgesl4YmPJrU0oDodkB6VDQc/c/EbZjm7jGcRHJSBZuc+dm
PeyEfB6Ow+kTJSJ1nFVLatZ7TreMEl6PO4zBxOMPaC2MlTXgcv0814HnXfIG
mcJuadFTxgLkSxYpLcFXaUlflN6IeWc5xrjYuoDFkbf8oeMkCbXlSiEJ+3TA
nW5X5Y/7cQo5v2gaf+qrxbBaAoG4LTBYGireFF7/mYKJxjG8BT8Koa//Equu
O0fclwa4T2cqaFIYXYJrnQ9YHPRDcA6J8TavwYeakKiS0EzYALkfeO49yCJ4
P0ccD+w2toqYCnBPFpd7GEf9+XfXgsMAAB8bH8kxIYiWPDF4SPbKttrXnFRi
AbrvOG4ATA69D7SsuUUgsLcyfMd+YXjmRnZroCWMHvRIR5xDsX78fdDoU4pC
kFvGjOSf+okA1VdbDIaG1XGCBVgMB1JpMA++LyymEMcDM0xzO6fYWfv2YnNt
GrAHd70PQraB9VcdIzbWmw/T7JRyjkXNWJz+5UA3jaieBYYNzAkB73g70Oau
gFlsFZ5sb6pi/AV0aTi/Kzc+qAN5XjVNKJ5qj9V96DZ1r4RYuocw/YQhvyyA
jN38iVlnlSyw8eSyJ+LfnXA1wvZpMCrZjeRB/IUshn2jHrnNcyWk3wYNiYfl
Mt2e+TsEUuwSv6SHYbRA517Gjl9cWSH82hfTnhY1PyJIbqgkJCW/6OHvfzXC
cAxf6eLHKyff7H9KX7/hWsdWmukKKUv+0U0zgayAtY0NPqXxhtF2lccCWACz
RYuuUUsCnuKrjzJchWepYXBdAUfuKHNADyQEHoK81PdBAS+3UCr2yso9w4Di
3u9bKLudlv554EuqTwbvARi/WPwyf9e98dLouNwhaHgfTshgBOwf4IIKAHCL
5flSq7XS6B95DX9LE9XnQ1YzE2zNwtZ+uRx29tNqX8nOM77NjBqBa9QWBUTI
wLBbrsP8OM+N2Wy/117a4ErgR71ZnkgE4p7u69vdwtpDGJCdbzUhor+trN9n
x4rIZl+OagTl8t4RptofEFMdWR6PF0gmeoskpqnlZKAWxz8MxHBdHcjHk5QF
mzK9wGBbaWbM0a1uxRijNATwCvnbvwbPpYo2Ieo6/D72ztcpIrOUmDGkKjcz
DlVBS8YqOAeBJPj9reQ4oVPU7+M29atgckyOcSFpqe51a5le6tIUCYV7FJEd
rkqWbBa82iRwauCl1S9+MxViuuNMiBEa4bGsIko10C1ztpmTf0LG/iqoqUPQ
LsWr4QdZIfNGvLArIyS/XYQ1R8kEr3n9UoPCJelIBK7Br4Q0Lhvm/T5NFKVN
L22k/Xj8FARpVu+iFh34x7DUTYXyWtWlWgYV7H4j09X2d5v5cUVj8Vejbc31
p5YJ9T//GdE9VyPtSssybcTSTcm+NM+FZ3CPXfi5nM6RTky5DM30gzn5jj6/
tK4UhWc7ywUPchcoNZnvTkUVJhmIfMtm3zWx9cBrm85kRKzqgcjGLFrGRTKZ
iOIsSVIB+5NIZgt8Dm/IPlHNwGYEfZ0sgh2TiVLCaUt7DReKDmpmq/lTjvMP
NYhH09oIfE7FbHl/y3pShFbal2GAz8SPwVoqZy3GstK/S/JZydn3lB6ML8I5
VkYepZL5OwpWvNreFOOaAHdPhoKdoUoXbXnO+YJPu6JeQ1oaiwqfr8w+Vohh
wMDoBmIGlxzFgg0TyWi4awyHhTUtikuJe7sOLdYpbNNqpr/vwfBwWzqFDkEc
IhxGt3mB9e4MC+KRc4ytw+IGSyEk0IH3NWpcPUB5jQAHnPJsiF3x06s+Mx/k
Bq0Fbyb1CHNKmlAQjquu2TfLkcYo5QPFwqSrvB3nn/f1ERkAwBeNWydFs/eU
9NxleU6fKqDMul5Yzc3U0sb4RFgUdX6a/Ft4fUENOBuQetSN4QF759bBw7q3
ce1b5uUZVS6ADFBQzn2p3gRpBY0YdVRpIjmnU2m4hHrWpd1JnwLEuc15jCEz
RtmcVs3NCCUE12YoWiSl+de9ObRaerCOADSiqafvl1J9zQ1X8R7Zt4HBpBl+
L4mUAB7RDXePdkxhO5Qw/yfQqfXiBTxeHDpk+vRfy/V1S50jbMk5+SIasyIL
g8iMJq5Xnuqs6p7wmOxV5GXT7pQK8KNfUS+jYiN23D/rdWVpwhfmL3Lf9oLb
CVHDZXU5g2eJ07umHwxZGCGDQ98MU4braT4SV2bKBDbCEz2WOBlEyrj/cGhc
1nisc0AUmlXDQjdmM6bA7vvn4WzczSVBWmTM0zvEyo6UFJQdg2OZSj+GDdDY
HvajknahVClsWxYc6f93qN5XLsh0/CVo0VDhyNaOZsfN5Rk38kkGj/3JvkES
FJ1PzKoOoVdszm1qFmQEPVCmj0weqyuT+N2NI/cDOG56eJBdRdfgwa8aX35o
Zy9okVAH9UoI5rdgApxfhuh3LWjH/H2eVJyO+B4yS4IdcL48MG9iDMwzEjMU
qQRquMjTuqDpfU0uPQEhbRbnE0jqidvMSFWIipJGkL/TkztXzDOwnJB3kTOX
j2vXaxvSRHq6ddBtHYfeSPPg3AohXyl+mmDY8jOJx/SYcR01zg2SB1ui5isE
98guOKL3p19l3ta1KGUbWP8sQTe+52UeLMEMT52pBtKBan9bkxtkNJIfc8Xt
yFlGr3BK5F/7odlKSD9Exo3C47WfZ+95Gnw+5tE5s2fRAGUJcJO3Gs33c+mW
FoN+D0kzA3m3At+GFX1hk0O7ET0+HLh8FCN1lNn0OI06bH8Ogf93T4A0BtXv
SOkr62P0bFRGJURxtKI70YlnceIPjOqfpTetWNkmGROze3npXg20Cogh+gr9
WKAqxq25ZYNGq4wsn4QDClmFH12V8uyJ3EI4uSpCFQv0oxGXt7++6Er1gJcD
zMFpohJ2lxpa2XU7CX+qWgo2x/QuAVzmj6nmv3jA8mxGBan61OUdDBU8e6Ux
DcbzAXxeXrhBwLo8zdvIsu7PKkenfRY/liDF+EG9SQxKHEnDv3mhQYlIe5Zs
FFsaJDD9OgOdDzSUbou1iBMzkJRfcp+381Kf4aOoOXkCZeVRl/HNgsfQk2y2
Wj/nm0+bqiClpY0RcXzyTXzj9SRStXkvnq7iBv9Wb5RHMHwAtLCAVA9sbV9D
UKtGV7obcmFEDEsd79n4fM0vkdXVpoq/jHWCUV+JgD3oO3kKmMx6Ppxwd1AA
jCZWZ67iC9nnaf+pAoULwK33pMlU/RjyrICC2e1ekO1Y57HM51E6cxfFTt4E
ttpPJhq5mZncedorLbBftZCpY415AX8/JvWAAC3MgENrF3wFDzF1FVNYuXzo
RdfKbVlbJVMHP3k/BgNL+nQjO6E+8s7WgTfrZVhp3W+A32Mqfn2H6tVo68+K
/cGEEMvdoMTehMz9dzNpW8AOeRLN9l+/GChoIq3/cdd1cMHSs4LihvxkFzGz
KaUVONbfvY3DnDGHrtCBoQS+bqw1uRXvPGFEG/5REOc+QJ1uhJpkS+RRQ0HI
rK/XfWMsMNGW6uUjxaq0IojKZPXg/SmEppn4yFQY5ck9hi4b2xy84A6jsqyV
U/bSUvjzai5nriTk6P70Kh0F8HNI9enyQt/+YGSO5iYHBZBzrXtFj2Jz2ifA
2x+KsIs2T2ypOdSkmFePx+vZigwZujPDtcIazlk82R9B5ox09k7Z1MLs6Opg
+e8AQIrNqlum0LymBFXiB0KLG8le5XJK9HGyGibKIl1r+HUhXtFAxgSPKXgz
6PzAxz5XEBtc6sP3zZpHzGXRzgEskyOFrzajgSl8JE1hniEt+NqUgom5/K1Q
hHruyR5vcd6LKTWJIxee+GoEupy/RnANkRtm4oWdlOX6Cw9ZNpxratICUTxg
Ob8GVwnBj0H+6Zv0VJbDSlb9NWX38M1QxC3gAOSl5XpZWjMFOpuELdmgcfHH
35VpsPBuKiFkh1mVRAV0lvSxOAfggajWdZWNGd8V1vmIUliJnzsBrHqHNyqm
9WU6cazwX72yLKODZOIBqPEGKklyGTnW3rLwKOzb4s4rJNqi+ktT564fCSE9
LYUQgVpRvT6xJCatKRmzQiFSXAZVFfcFWac6Mx9vKEFMrypEx73O0eSkH5HQ
W7Yy/dbJ9wXz2g5SSSXss3nTww4jKjUF+vWmM1RM0Y8jZkS5C7PRT45dpg43
Y1FQyVyUi7A+AXyAuYvsIUg9MLwYsPCC/0DONj0EI0Cpd1BEXCUstF5fpVfj
uXiTFrjFbAR41vIAAKHpDC2MNtxy8jB3JtG1tGEAMFgwM8DaghJsb+CeTwAo
JK6vf6EXwi4yuOLzzFyVxVmhH2YDeo49e6ABH0YWrnBW8Dha1nk8/g3NbdCj
i+rtpz4x7ahUZA8J9Goqrem5iTHSdSjJnGgbKnoBKs2F4WyR9I/jLVWBl0eC
Fg+LnGY2fh0R7e+A2LdDRUNaVYQ1udZzA3/O379jdS/fenjiV6+p+Q8QYlly
W5crs7k0GbYFjcZoxUJu2TwAS0v1ZJEyE0lLqo2pCZ4//41Cd6BESo7egIF4
2kK7RzTJbRCQpn/SYD7MjyRX0HCnF55CL6qIiCFPgSpvCbgOyhwYqyyVI03h
50jJnJWUGopPcS9dIqL03Z3B2A6Oc0ARDLt2wy+pdkA3LaXT/CoXMPtE024a
t8i64KmcDzrBPd/pblnzAssL/r/yHQcqaHUPKRaz/XiZuGLU0WdybXb+mAsO
dqdt89vVJja/oKiWR0k4OXuGaFHSR6k7691PffNFzg9To+BjdL01/ad5P8Bn
mNcin5asrSXbu/WZx6tNZST4KHpdw2zHZcG9vK/D7J55Yg6kRyxgplVV+wI/
EQeHfpG6eKeeIAds1Q5V9tBOBH0V7Y+H1eDEyLl2sDw0lAEG3bE5pJ/vq5+J
mcWh0/Oowe0QbwHjzKqfgdIu9J5OU/sRrgggN+UWINBceNcnVkq0eEIbwV6w
jrmN6//qsjWQ9XGICsJArJ7fiGvAYL8Iwzo+N6VPa6mHvwvcq2KFjIOcgsTV
4tulErAkc1OnWHErK7eWyyfCK87m7kiUtDy5+Cqx7Ct/qrPbpEjp6R/dqrhJ
1JEyYQD//tg1QVBWELgyTuqgI65AK6Bsd894Zas+AKiS1EHKNUHpXQ9R8Mhv
UELWeWcPlJA111H1DbvJ+yRa7J15tgMhLnHvpgkFc86RX5O4mMviAPAEPPYR
0TSl9eHfh/hsbVxT/I7ox86jh2lKh15+9TLKAps+ge27cGd2OBUDflSNMPW4
DQ7qNAZAje8S+nYIWw++o3HuMeYlq9ggrERENi15QiFNtzM7sxTIRKwRv5E0
XOO2FZ7FRQH/JhqaCeLYCbOECpjCUyfE/TxCdhydS9Xtg/o7X0F/aKvth8to
aqBMrs5RiPnv+jKR8IpqnjiTMbs0y159Q0/+H5S8AvNmwgbq//qQc4HmtV9N
6893aT6WPusCJP/+N/T3Xw4avLgzs5iR6M/bEXpiq8favXZHJqSVhhAanBu+
BeMkvMPWPUNsWXLbkHSoV2CmdmIoQyHgT2ms9OoPCJiFHB1CElzy13ZrkdY5
ESSUtadVjiS1XEaciLciAbYhrM9IEvcTp3POcOdeYiiZ9JLoxztqVWnEU73E
QeZXhfJkSQcL7Bxd+ew7BIOSncupfweg/qQJYdyuG9IpYVvmBoK1zRB/5BLw
Bfr+nq0VqHQjJhwQuBCjwLZ5X5VKfHPovwJOjo8RWBBeRZ2cB3YsYzz7DMSf
vxL2eRLDpPwqg6QWTJ4im2MlydFPsZwmiWTWT44K3y88vIC0BeYIT489dVZI
drGubIKNFd/p9HNr+ln/aYOmsOI3OhuuCIZ9Gpn03Ro4BtBtJ3FWHc474MbD
aRb2W8kFxddzfah/UK4kPJ37Upj/OhB5EHcM4LAeWrkJI+AutPY1h8/1G4DZ
YhxDgMT06Lk4TLj8grybXtLnFPZQfc1JRIXS0D5kj3IP4QpSnjdVWizMBlu5
yYAFLMY7kjapf1BTCgrQvDBzkwjbPvCuPeZ35O+BkXdXHfSbEYNtYVWVpj56
Y/ezeXGt4V9L1BxqC+AeWtSNbJZcLHdMLTetVErBQKrLWZCPI2vlcWLluTt7
kPDdB1wIsfFqJfKTDzM89kIkW6udXlsi9Xbd76ip6ki6eYm6J/gO6KZUFQXA
73khC4gVUVGc60qfDC0e2oYCEFZNHXKkU05kbd4ITNUWdkpkiHzrRCVHPBgw
hlYwz5iVPUuUKu7ENsy3OcVB6vNOvnw0vnRK+xExTIvfHeWEueNkMu3i8+J0
BEhaYBOF2O/wsgieJE3fz42dgXjsB2z8Za/oai+gDOFsFXO7n8OEhZj9YtDI
W4YabdkxhsgWK+6ObLYejHpQB0Rs/3EQ7oepXN76RFYc8BONdAaLl8BYi3zG
S+GfNLYupRDGw7LwZx/N5yzRYXdDohOvVDNxWHO5Ph0+jK1HKhUso+jCa8NC
nLmn7W1u9vXfQTQctE2cysCmHjVXVxQepS9TVZOH45VHQaH5Y2fj/B5SbXTN
Jpn4/CUwqMakB3BfGlo6f6B3fEJdtfGG5vgmXt5fXhNMEMnQWO1bhFkouKjO
o3lx93xu8OkbA5bQFzm/PWdIBqHAi53q4qPX2R6tOfVhkmLzoVmSoTFXiZDI
KBu7v1mweEJDCxFSdWHpz1XWAh2YJrFBonfupoULglly9q2K6160YFAmE31c
fi6yjZML4ZGZcmDo+XdD/saKKyxa1OGwWLNqQkNYL6dLX/YoHa8XG9aiZB/s
hPHprPOC3Lu/aA9i+i5EnAKDhozdVxwGhEa+5Q7ikrLMaGdrElFp+Xv38VpQ
brCpdb8q7kKulyu842Vw7Vmw2O726cPqGBA63ZfuBooxdqoYhwopPs9/Fy1x
J2wj9gqKnihHdglYpB9aLwFbrMwqu6ABD2XTRXcg1wLFeBA3ajMWoZNLHxM7
aCyMQrZGE8B02/Jz1iyNe6d0z28tfbM/5Adnbb1Ue8jdUUtfLPHGqwIaIyLX
vM50CxpejvmiP5a1QJPTyydROxMXayFjG3L3R+dYWYmROAB+TmAfO3zKsHP8
U2l4bSAOxBwG9v1Vx9yIB0t5Tzx3Xs3aoO9vQHARiEGM6X3Pa8rTlzQ66Ak8
ZqnuOwNum43GDpNqcXyFoHtCqDemKYNdfeIRF2S4OdqRhSqbt31wlDeCbPRf
FP76uhMHVBVISfLGn2mHLb9/C4THCC4XQSrydDmRlL/893kw427sGLF3hvM+
l/VF5fB+Bn3GukTnRVR51M7VPW4x5QrbeYUSi8L9w+f77MX+EccOngvCOJ5h
l+btY9g4cVfmTZ1RJox1qVsSWhjyOAT1HKh/ajnr6nP9oNmaTR2zcpu3JiVt
sk599ltNPngnNPqKlaVXhY5zgmJP1Q2XPbfpiKvRA1yoXqaqsWijRvVN0g58
5ayFPFkCElShVMCMelKqV51/RC5htjjQB3LmRWoRW6HOcHpuNnBZkbdByrL9
OrBzkuuazLwTE0Y3f2sTIiKR7Agaua6HkSMFRZcal6ZGptgkQUANVBoZAGU2
+v0oI8HFKtlcYBDuL8j9eOfwBZ+ArmauGI0guIJd8nVUfRS/wgi0C9/uh2gm
TxMIfTo9xnrkcd0nlk0hUoZBAqAGTlRXjNP3TBqJ/rZY+sARNQrSG/5Cno7G
dfpBvvSIvPkI4t8M5PawwUw12Dzrnlbxpkm/Fzu1PQSg6ZBXHBgBky8nKAHh
kkpmzYdz3sekjiHDtoaeKG4Hux1lmdcVCN5gnbFAF5K8dVTa/xCEhSf20EBP
B71Tf9o9hquO9W9pj5lTU24d51ITWYBAJC+cyU+1cvazhgq7FHAlf25T4KUg
p3M7P982v2dkaUQ2WZ1K78OQAe3Bx8FNvwQuQPmthDgg6m6GoOF9NpLkyux6
BcHQscHuJik3uuEsZuFxiTdITxm/Pp98mHwcrwJtw7dEsp6mUm5u0srq0qHR
QW2ny8Z1A9RYzE1y7zZWiYE9AdW5kLOyusJyUkZChKawPWWP3wupfOkAaZvN
MkQHazb4G3dJYvJS3NmdDVB+kINK88PJLpAFGp/U+FTxKTrO9tSECGEk6NV6
gBAaKnnr5KW6pncn6gdRILJmvHcrmHK7wxuCendKtF+ExWUDmI8OlXj7Utoy
TnMXeAzJgmRiKHyvoOpXHr/8nNeammcvdIUFxdkkcL/SOrMOBsZFMQrY2eb+
+0D/4hCKnRkCp680aq7WKpvLAt6CYYH1/vAemRVWAHwDJ3N8tkL7jWLmxaPY
/MzsvCBXtvPAwG6Uo5vfWW9yHYM0UT/PxA5BthYvWKfYbV+fTADz6PkZDmbg
HhJfKkny+ZAJabVuepK2arWTkFCMSMdaFEx285a17vIchGmptS9i0ytK0mFD
wcunTTV/p7yhYoD6ahAc/G3QXOPXwRTiCg93EZWuqIec3fGsN3UCWNpDbZvx
jgpVDRXpmsy8xadIv1/K35DC4T1qE13n0255zRIszj602AwkUf+0o+ygTqsn
0Ppt9CWjF/im4yAEnFH7TwuDt58eba6H0/9oBeSAACN2oC3ksEm4LFnO1zn7
IV2s45stW4/ux72zLa9AKQtiBD1LTphVlbiJIlhZS5EXhdZ8WPWz8ZRq3lBK
xlhwFc9qDodSdDrhrTk2/lIOliTPwOv41VAsr35WD5F+zL0TsliHOZdUuDHa
XRwl0NIi4Gq4hal57C29Ej1efGlcVxNWtLpNctcvcyX4ddcTtnZ4O08c149z
oMkoqP+tpQjM6R7CVfh8BMknFCdzybzddmnpdyS3Q4lOkF0DBzgyeoC6W5fT
1p0IgFNdbmFOOgs9FWu0+YlnJmXJD/Qx6gFlswo4CL6WaUYZt6T3oBqG7CcW
kRollmaMEH0c6uYfeLwbxeOHupefWX9i5NFXaUBFBZdSmbRzddFOIgUYFKwz
GZS1DwZ2uncFdZU/EQR4gK5BM8J3N4af59hgz2eHgxrxOyNNcwv+adMTbt1c
DoqZ8G/6kFUj/JWgCIY/bVKEfyjZsv+f+7Utvnj2DAiBo7lK1Agkgyz7KPNn
vN3KNuEO1Ru3vEYL2kXwqR/6Yo/v0yg8lhQNQRmMi93kAsk+MYLGOP7F7w8v
xWsXnNSI4bhviOSapXiCd3AjUnU8iVo13fx7AkISqZJi6KUFmOBAO5qiGrVd
xd+NsHDyiqtO1iXpCnCh++qnwWgw5vjoaMTEXTnHV3AFHUalK21k4NJ0ZUFG
DkYk8zqhKV3cpq7dgbC0EjsQb7FLcAFiox0SrLL1QMK1jcz5Vxu8wXEz9phX
dsE+CIq9Fnc4LpxTO8LwDucxjcnBbvQzgmGD4kr1c87M6INvfEAoDKcOIjLP
DpWoa1TX1dmYgvgdFIAAlkhxPQHjKzQ35umQjBizRdBXPHeL/EZVJhl0GCJU
XdwQnbqVCNIRGei+xYgX2aQ89+v5MB93PYj4Et/D0Ha0WqXiyYKw40WipkD+
g07Qh5zMH7k8TfEHqyvdqITCR8/PJBTDjmby/Q==

`pragma protect end_protected
