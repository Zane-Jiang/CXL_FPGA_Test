// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pa3mbIO45VlNvciNiKBDc/5Z6Y5PCMG6UMT6/KXR1VeNPei376h+F0zlLEkh
2X1L3Y4UK6TCyLhdeyrfRiAkfbJP+EAAQwAnimC8lDpAvNhQ1NkMgPwwSSBO
dKvzru95zHsyBfAlHPjk0vW5ITnZLI3uGKHJoW7AA7szgVVhAJOBZ2rllkjn
QQeuAqU359IELl3N/GUuqLx1gqydoU9FA6m8S8nCwDfmTJFbCT2Qva+Pzkpv
ZB/rfZLAmT0gIJxh9lpWVGN+Fjwzmk3Pm0TtxflJaFU5Z32nyemk4Q1gXwO0
VHaRK5stciHIuRtuiGE2kHWateMIvkln7OWHRILGYQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kq0iMq76cmI649fg2m87hodCXVQvPIgyIjDGqbI/Mv+FGCGzaFTYXxqm1C3T
qoO6giGRYpIATfvpAlL6ahyctL0dZlQ5nys4atfXKcLIzogI//PxJsTw19Fa
oMAbfYr+t9CqnGZeE2M8XwHagtY3V2z00rgnxGePOgy+IoNM/b68GsCRIO24
jQT3Ngkth1IzsfWwtL8NyDGfnR8FpLcpg0zY7kf2uBJ0mAdU/NgpGfFzvC6+
mjNQIlhDYf+h9/qfg8ia+YnaLC3JKHJhVPsaKGS5Mx5c+tPx7pQfYkn7FrwT
WtYiko41ahObkjXj0F1aNYkg8zt7SA35tUGufoXU5g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d6BrVKTwOQswAqheYe0kRRHmr+M7CKXEzXbh1ai7R8uZg1iFj+JEOcSYaRzF
srL+Db1Ie6l47HA5ZOY11V6wwID+WSvMSvbSdpPre4z7SI88AuwqKW5BFTz8
1xsddniFhV42cE/hzxEB7XI67GRPyuYb4EaDnt5+GkI/LBEDRk2c/KIASGA1
DLUta2byiK4Dwec3tHo5wdAiW4QvOXqxOMsasYpmsdDfmtSF9nCrW2+qfefC
LsST6JILIeWZUSjFpZDX9S4jqZVoRgy3vtfyPt3jAIRenl0j3r5YWZfnAb7f
vibEd5T8gZ/rU5z7zBaBCS4BC5LK5zwoYqA0+nJjbQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p3ie+G6A7kJve5wjKPIJbXuGuiUNmPVZzI4nTPLMJD1fxESHUfD5gFj0NyiC
390OrSltUdH7z/OXtyIO6KURGZ7txLzmB6ZY5z7kFw38w6EN7e+UP8/jYlg5
FcC90GoyqGn+chUz9yT8C0OgoggalceT+vImXBSSLqmyp7Njbe4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
A+5VFBuRR7RGa4Vmzs319i/c7climu4umNrXlJN189Jtcn2E0cm9hXFsCyBQ
vl2zvNBJMi+5ghFPVDxSjWxmEnwqimgRc+wWX5i5XDkWkm8MQht2DotOReqP
4YP05WlAJoQ7yySQLpDIH1hnTxvMAg2L7cjBHkvLCZrokZfGhwXMYrvHJyV/
qW/PxwOxLeY0X05HhZt3YvZTyCTHSyeIC4WV9tINJbKdvrnPOcN6PxQdAbio
LNO8eyE2tPqexW//LYGJw+PBUpt0YKTiXWtzEM0NjqR3JYR7ijegBA5eA38k
btpdGgL/+OxznVlA7nFEHDGdrXEO0JE9su5D/TlN/z/GtKdaF9TwvJzolPD/
y2ssUtxXx1bn4ueC7OwHcWqsgTJWq+CEeJJlYbA3cZYVcmCC64Q+6Mr20B04
P61aEfcLVmYNS+u5H13fdf7NgmOcnI5k/34A97VKAXp0bH4lxypj3ZENIJUD
Yufd9+M1IzdbZgUwVylLJeXmUUKj5mmp


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
C5MqdO8vj3YJ+JMLSBnW5Hh84L+86vi0fS5swoS+t+3tsVDijugfPnDf1icy
B04HQEnaqNthM2DLWhDI09IbxVybgKFykp++cqAhIDKaws8Oju1378uS4DDX
FLs/I8mYCfNGIRQ6LGxaH7bFpzW0qeUOCzDXQmKj7D6P9cl9sVc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pkGWdO0FYoF+CrHdWpBdO9xiTFk7RAcxWIZHwbTOEksU14gIOaiMVOCwad2n
UpdGSbnsbDZfIqdlqBPK/NWFD7Lkg/GVs7gfPKFmCdS/RLV2+vrS0ejCQ4D+
/UkxeU2gHRhb9QQb5jYkykVADfB+EQRe7ZgS/45iMrtNUFScLf4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1344)
`pragma protect data_block
FT1Jz9NSQ4iT9dqo5Htbj9HQB2H0mlLEnFCGfTRf3V8VNVZZMZGXA5XDJrfE
JPzZDXx3/H4MizYy1KE0N6S0KStcJIsQQZPp7eSGI9BBHMhV1TTvbW7mdLdD
JIMXzESj3PoD2zss+UbCm8w+M4bowA2yJZPVrXpXe41A4ckMrrr9YGrsp+fX
Dplnis4Z7Noecgcd56SoVl5XGRU1dVNx3fvyfmtfx6/AmoqN622C+MITo/Tf
uF5VlvMa3Ka3CKeoTyH7y4ROr/lparp+RQKk4eidfBb/orL9UAa4fhFDAvz3
N762mSl5LjpzJN3R+MkfpxO1WgsTsEOxArkn9uPgJHumtIGK7vP6TimAuaPX
LTytZm+icnMPOPsHmkdCt4dLTdEnqgLFPLEXv1ucEBNTcI++I81z9+g0+hWy
UYc5jlFVwaR4X2j4inqP1hwhRBkxdvy0DWr+BIaOosnm2fo/aTRcRM9usi7f
ukZJHvVS95GoBXcFqFOlHoN1+R+i8y4f9o1UbnP9u7uTo1yL4Nks6M1Dbnkn
rf6RnX7g12iTHtwxobhLkJ/DZtVyhc216Hx8k0d3FtvE16a7IMqx7kNjXDlf
zEUW3QahOwldhdvPrNCipLD04pAfZjN8Sf+yxp8BSUEPbFAjCH1ozzxIOQ9G
jq6zELmvmhcGkWUCkn3fBVCxILIWz7QRbSU9XDWKEf9J8gce1XeO24y/BGpp
j9d7ylzboSYblN1mkdhN502dwP5+Lr0fxQjC2eKpfOMlofHy9ke3ACcw/+AO
yvpPbXVrYGAQqG8epJKk5Koga4U6i0MZ8ppDCe11ujYCB15McmfXU28K1CQG
7QmVogEJdp9nZrkL5dEiNTLrtfQq57BsLU771Mfz0aLmR2ObH3Y09o1E1WSO
BoUG/gxj+KxS7a5Fx84bPYRhGWw34iFsZEp4BFWbX62oUMDzb3mv9FBu73Ax
6qrMUfvABemXWq9iyvwMB76u0CylyQzy617h1w5wwaiuu66unkTWM7AgPaYk
NRE8n1kH0Oofop5NOu82xcp1AxdVCIJXazV/Dr2D1MOYjrk549tmfziKg7Za
Ba933HQoaioLKiga8naUYOSbzA8t2d5Agd9sbB2ANXv8pK0tqHptGCqmQnkd
euxzlTFE17Q6bqtWC+e6ud9ohHUXsFj5KNBq3dl1RGiEBOSlt9UoMpBNcl9g
q2A3YyAFVu0cAfl3YYZrqIWcwIuGdJIih46mIcTiB1R1ZfJCEpuGVodyp8vP
bnceW4WAdbYvDnuV8EkVvq6edzd7nNRVmEPdtfrTZ6hXEkAlV1x1oIp65CCa
T5QqpuDChuCZxf2f+WdTkVRTtBesP70C2COICPj454PujGV+40yAUfKRULSj
4o45soCCPwVVYOG7jvR3ukKuYzNcbINZmdgpkXNDMmrQzvKqAHDD5UCC+4hj
whqC0EphpD5gNRDTjsLTHFeqwTQUNUMDpNWwvz6z6dquAomy7K3NM0g0HM2O
phXj9jemrrMGY+8k+SuhLv4RZ6vjYXqNXM2T2sL7UI3KzBBKVmwiCrdQswEY
9hrmKYyA962TK76P05F0MWGMPWSn7NyF2rCHgg7fhepkGdBrFo3Nh2F1MNz7
6kLtyIlNH6PGb8I43koCqrjvxsX0S13sU8XcfjpmmL1KfQG1AuKcgrCtWE0F
p8tf+P+VZzl2XtYeV73PXNuBj+hFi/ZwmOYU3pC8uKK+XNNxisM1RFxAukJu
QEJ3bjZyWSnAla0IS/ATXmMFtmqHiGVK0f2SL9GJrhZvHh3+HpFJ

`pragma protect end_protected
