// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
SuZ658awRKYNDFFowOxa9crMwPUHFtAgMkZXaqolw1lw3HEOXDNxktlVQjG69BPs
gCe1wdEzfFOckWGmyDdAgBylo4xJhuDzY8YJcpS2MVGxzIi3CILlQb4dT9ohcFUB
fYadEvxsbfLrDl9rgdxdIGJgpjde67RnFMeLbodkZ07P8+tGmNIidg==
//pragma protect end_key_block
//pragma protect digest_block
M8LPWZDGD16g1GDQ2qCG9LUA7qo=
//pragma protect end_digest_block
//pragma protect data_block
6mAZWKgCa0Nc2FCzfKIB4mZdiLTDZWYw0pXBwBvean+bFAEDI50oAOz8SwTx4/b9
PeeToko07KKgUFJAfn19jsLRVJEASBYr3zFz/G5nCNgsIDX6cKvEugl9rmtRGWqV
rRxN724v/Mn/WlC4sCEE57s82/Ho7zv/+SBHImPS8+awuoiS8i7qhF/bS+DvzPO3
dAySyEQ6wOVD5iCbU0+Pzhd3nQC/a7/cuwUIAFPtmORCbrVD+eDSZ6gx3TMgSWNl
OPYEvjXrQsCIjtyovdik65+RVv7Lx+uWOOqv1dWgofnczy2vPSrqfVXKnywHTc/W
sUlNFPmMsQkE5qpTpuJhl91UTzpDFzYSR2Un+0bxXxQ6r0xxELMAvBTsQOVSd6dW
rKb+lodJ7HzMw4BVFYLGnWDj39ToMsgFq1NjjkzCyBZRDU16HlEEKQMOvFhBkXbv
1yuhMULOIrTaU9350zfM9sljomg7Or3rodfTqP0D1mavF3A61NW606WVAH1T9i8T
cQeOoLDH9k/n1odM6VX8WPnGhI1w0FRE2pNOjVtWrEFcOFaugGKYzHyEmSQTkswS
wa7YfjfgmX39gkD4ISyRd20QKRzxH8Xll58FvxD8seOi9KyhVve1RCSFtpiNWuyi
shlhS/slCY7lJZt09DbAnhk+TVMbEoMc6tHE8Z/Y1nxNGwoUP/RcC7utgYwiTxzY
DCKz5RP/QoP92PzxPzVwpg9OmX7dNVyxVrK0JxqgQxZO/ltcoP+7wzuOLv5VWsIm
43uETspWo8y2HPUFGPB505yXGE7x5HouwdBQ00EWSteBpXx3+M5dvPVk/JQk6b6C
7ZiHhy+aRdE94JGeHOLFg27FobCwil0khwV5Y0KE06lljv1rvrrcTW+9cHN3Zcfj
HnJgRGs0EYtrf4iLGQBlFKgqbaiVdNwcXuBdsH7aHudd3XMU+jndNwfEcglfsylW
H3KI1s2chnTYw/S13erCG2HbibRjKcfZKraeFW0FqMt+NGEPBnOm7HyPPOINWNsq
KPbWSWJco/3N3AlFeQBe5zg2aGv7a6OzMtToZ+/w9KqgBFDej0yR3bfA1BaYLbbT
9106vWD/gGgB2S1feoym7EPGJItTn7xFd2bS9+XjaDus/VjBqVJZghZ+MtJhjAEU
oiAF54avD8S8Hm8/k6Qy/ZjVv1tIxkteUgVqfcpQdaZbj06GnHOtXAndhmpVCfDW
NJVy0VFM6X0+hoBBTxayBpqKqBFe8F9D7waVakJKTbsAuUqmwt2UHeC1EMLqsAHv
MgVdVhEqupRrO2Ue9wHp+YpXEm6iECz3ofNDH+EurGz9vri4ZR2/rtKxr+UL+iLI
4UMnzt/wH7Lb73w/I3tqedvdf0wMxwWD59Ml3lbsKaR6hNPi8SJe7ax/IMN6FC8q
NE4D9VU6InkcnBdEizHx5v5RUZBIXcqOcmvpht16HY8MaubdIsan7CdTxOSJahuL
wwoElwkBWtDbSUL7DQ2nbPTeAcPjqZRmK4y7Dpto1eeUwq1Bv9iLyWq5xdkfYUhO
5hmCgqsgflQIbFO4hf0uIvgeby+q/cbznCf2ExaKa1rkDCx0IjiXy5TTA2Skyv8z
k5+4d12Z+UvW/Wwlr0NS4L3XxDl6RSPZ2AaL/NLQguOqq1rCZUkHn7WqdcV0VJta
ZAqjS04u43ikHxvKX7x9g0Nzfq5XMCTMmx4AL/mBvm54JafAVGKQVlbZSAgE1caQ
fDkupW0DjBTxG/RQIRgQNFlKlX3C22+19OuAUZLGdWqGKaewei9Pdsc0X+8ZZpWm
/8v/A05WPjeTsGmuRpmrbgZ41Bkj/YhNNs+cWFV708qLdKNh4k6AkSTElVjZCCCC
ONsbKe0taL1BuAXiovtCv4VexAyy0qp7gRfYShjv+ES1UD/ac1m5Hf+ADZHL38oR
d0hQUVjYyccZWtNsxuFutEQLxYfLp67wXjWAwhhg0PDKYoXT95Grpaqd1Zz4eBuD
FvjRhctari+z7wUC0BW93srhTVxBIlyku96znb/pkOWMzn0sGXxSJEorP0hj4A4N
PUaJ7ObcOc7JDMUDPOLrRAPRffhfTaMPVT8WVIzWoN1w4FVaP3GJ8JzQ9HKg0T4W
SdPUXORCv3aYucYzSgtq6AZXUDfCx13/j2KppEQaSpMt469stYELm8/auaLrnFkt
3QZ0eoxxAa16MmM1P5AVfSGOeXP+vUvaQ5cSMoo/ZdaRL+GyZ5VaMrUTODBxk4tN
7Me2Xsx1NAWd9T33zJBq+vyEFzc+3L8JlFRQQnaaZGf1uGXwitZWzIkUFMYJnO1k
zPNISdD9gDXbGB4yFf3n/N4f8ezGgpfbCOpWjcMNxjvnTO4MZGOQDgMQ8HUbtV1Q
CCEzrpXKTAtXCuOPQ5qVSY317+fAdLifiIcbhdv2rAEpKTPTRgMbY+Np6NXk/9mC
ymSs9xX/iyVX2OHNhFA0TT5rPCrksVGB7BH1g3SH26cTlGs+d0/P6zfTitC5LuMm
sFAlCMWTODDkBu90wbxPx15rYJeL+olugOvMC2PBUJ1wLx0LElln03GY9n4urjBL
4Zd/FNQkTs125l4GC189+laMEoVdck++dP137SV0O0117HoVmEmqIkiJnxK269U+
Qnn8coN1Cp0rL+pcHf8GYAvm7zkFzD5NakQgCR++4sKv9ka0GCjBaSyYQm7e1HgR
I+OPtWpb9Xf1CuH4lSDg0Wrmowrl0//kORoDP/UIPlHp7NhLlP0CES1GwFp0udFi
gab75pqriiq5D48/2C0qaq013WsekiU6GeRpNFX/wmA3IFv3SaORh84qAMfUQMZY
kQsum8Are2Dkg6jfC472EF3Rv3lfi1jx7pnO7QrgQpOpWuyeSMH8xjZIZayIWXjt
ICvEz6+RysfSH3G/w3+XZByJhAWuBd64c355pZS0P8vGeOCPXzg+lrOwrOCtSLZ3
us5ChUjINrSk717kO00rFWLdouHUsP0cY18y+m3vD5o4kENfT0rDbaQF58EPh+mt
00GCCtnSKucCw5q2D51FUrZMcmY8yhUOFIzEruCtkSvg3OjJOrt7ZBxlLnUldnWu
jdu5BW/Q8/ptEc7xFply3yPAf4G0tO/paUzesO3TpzhsVKm2+iUe7aRW6avW8jj9
eAlkSVtBzKP128Ibtcq3tLifQdSIhmjoJwIh/e9qmtfEp6p5NrpIO6VKbToqYzch
U9wmfsQ9hCd0ZhRrd5PUlxeR5vYQtL0Rx/nphajsuVlvn/uAkk1/Un+A3ANtwjDH
Sx2fXGheTNx7pe8n6ydVZ8AOntGKe1Ai/XfsxJ7A0DMcNfw2VB1wtoJpqAXPpmgx
0BqDvgZszfo9A1qnEdtGJOGRWHTTC8G0t9YwNKjzQiDwRKkerQ1h+6nCzTxrcTqL
QR8Yo+WUS64EvjNih+oS2Z2QPCZs3ZxO184e/aXEFM3EY8ftnJ5vNW3tkTrc+y13
fPUGJmJni40hJ+DYNFIYwxYvI6Bb8JyYGdEyZcrPnCuc60dI9S+ogmoVbqnPejKA
MScmImFy79XS5GVgHCAx+fkWezSzvojPG3iah37Xoxm/3H69OpghuEL5M3qSaEmi
/MHUSsoVuNI21O489JHgWfIMCPozKP9XesVw53En5hCZ2hDwc1ypmbgTnAhPjix4
yEwQCc5uh6mVBILVTG4uu7ruxBqDvhoL2yE96FYNgH+8kjiGFiwXGL0CSSwhTKyp
7t7LIkTX6CrkNPZWzBllzKVuEuRYMuGVtwSjpYFC5sGJdFCaqiRt7PHarkNXoUGQ
ICMWUuLifOZcAu748tpTYnNKmn7CMYHbSPpNORGg2+7mcLNKC8Y2ENzvQnwA5hEJ
cYwrV9J1zv+x6Ub0Nl1btxWAv40gttr4NpQNCV9WB2aPMtMLaLCGPWQhI/ib4yhK
5DmOWNe9eXQGw77GZBgrWWjrCZFvm1sX0UMbntJcTagwlTmrkNCsF3+EkcAKHD8p
WLU6PiIwWra3cNaT1Kmh2UxhFvBm6qj7LI143CEydE1oQKc49GLREEVxAsUf6wZg
vW+8suzOdFZ6wdE3kuvg6O1vhcietyfmFMQFLLdjxOXYJivCOIIzmG3im19IJ4xI
VfG9wDGY0Om1vWfPv9IZpYUGse3fAhi/KrCj9ZyUWFomu5WdLvFeGalxjIUoAd+Y
y8xZVuBKGPEikw2rTRzE28H2Os3K6OhSCFtrh+7uv5/w7L4cL/PwCdEobbO5utc1
aKC0ubeHQM3pY/crpoUZfMTDLIHx1Q2SuHleV7JcEZGcM+E2gS/3wahdI6Ky3uBF
mXseCmwxAibVMX2XubjRUHUqhKew6MJ7BONZY62wq/qKNrbpybthRmwzKd66c4NF
raYuHEmRCXZuprn8qE4H99AOfwqClwxH7bXmwMKQKkxLTi3mfPmqkebhejqVe+o1
thLO9rRyyFpcYn62AM5vCUKQf0PO/qE6oBXyfB2RxRTG0F1yXHeL93nRMK5sClP3
+vaYxyKGaIqPO542IFwg0scoKM35yu/vzCm5Mt7Z9HukX63IFWHghNNApVP//Qxe
P7H0d3NYb5CgFnKKLMsJffZ3ZacyNDZGGNQdbE1gYCwnYP0/5K8Rigup3EMPbrop
gV0qiAqIbaL/LrOua/FLW+ORHQo32Fkzy7/WpJV/cYuOxdfG4QgrGyFgou+u8JJe
iNB/dhoiUxRGqh1QCaeCJZwuQWUw2dYgmgbioE7Qp+WvLiWqkn5kWx1Ow9BnbX+5
Gu6oEOxxZOgmIXLbUl3732Kwl9+qdvkAySMcmWgRI3Cim1NetZdbPTZP4fI97L5A
6pzZ8pMWW5gPc8HA47nM/s2wKnTSHHNDG8o2I4eafUVC/vaAhVgmvkmrAiqvNO6b
Hp+/gWC33Vrx9Uj7VqhvigvZUqTJJm4xvM/p8YhEqpJsrzjmx9VqRkWto2eW1E0N
1QN4idbzzv0C6qFTMMjnN/M0w4r56euMYrhF1OKvTe3IUrEbYhOa744T4fnQGoA/
aVuSsExavHNtyfedpgbj2eF71K34ia4GCpb9lEpf7f6C6zuOcjymLfDmg2qNdTzt
AyF66NWAHYnPxwNhunHCJnBCn4zgkzYbftDbEPTVnoyjsczOzAVWfdsYAGazvnwe
7z08V+DKChSM5zfLHmvLspAOGWtSMFqNNHOlcqFWBARMl3rZ/9ecO4PwRc9RntCd
nRrY/jYGb8lKKvRFLbtDz2XowgnbmXcFex04S0zHdv82CcFo0E2ae6Lyxy3NuDFD
ZI1r8FxSaXlxpFHzKBMjNQ5T2tet5U8OjwTdBpCG4xtncUmeCUftTfX0NszdhIUV
HkHxSHUqnTQe6QULFme0kvqayclAhQMvem6oJJ6ntPegBiCnMP/XakMMgMH7Oo9w
ffYGFeVINK+wiZOBT2dc5XBVYV3z4rYHEDOFB7JO7b09ftrPV5enQmOB6OPTepxx
lFZOMGgBoxAwNVjGdqOe2u2NmOnld9szaISvig4tYHzKO+4R8mysvLi9pUpB0dNH
D9vL0qAFXsrRl0xBGrstFsYbbDMhFl7xjpRY9HnpeK0nDzb+lhaLgn4hCJL+wnLk
Vh5iPPZOEq2HeaE+n/BNB1WjEiRjVzdwQT9Jd3eWHcLTzu6L4FUyLlphe+o14+06
D6yZ+wGpTG2x4NpPQhlpOTXuNy5ji2mdA+S3jXjGjnryrnO5ECtDY5IJEIhuW0NN
ry7Cbg7TwHr3boN8KZaGC+eAcq+64QXx6y2ujAYbnuiFUUMqhuF4YbPbjZxchNO9
WcjzE1U64I07SuLirMPI1gway6DJTkiitfS6DLgJUO9WJ/YVfnxZ/aNM+FkUI+kf
C2UL++8lCzCOaiR+UvFRd2Ew02aMtf6mkTcjYoxsj75POY4+BsR+Qjbrv8mAbiDI
NHy1knE1fP9CxdI+TDHgK4h0A8l3MdViGNH62h/Cax2AnvK2Mxqa33YpVCem/jff
1rJeNDg/1feqJF1gG/nvyfHqNgtcS5l+hjgTWBchiljHFGEIGamhrxQP4Oa1XqVJ
7fWzDXH6Y9ndaSAvBrs0wJU1uWSAZk08bmklUqxSHxHwccBDOVv9YuzCX3vuzp1A
Cn9yP0ycTudPXvUF12kgmCFMzpQGMeQOC7s/QW6DeeMlycbM99ZsIgH/sLIQinz5
eatd6X2ah3tjBr9UKbnz3BPk0xIeqiOyRBCKrWoTqsA43nHXXSFy1oegrpuGuq2F
AAtacnq+/98L7pEbpw2dkERRsEA6lsfUD0sh43fbFD9danBhjkTjZOATaTkaQolz
TgSSYxzGfuyPzc2N2QY9xyaTQEN3z/O53ySwmkB2USev2KRCPffGhNFPu2lwRSNo
UAZxE/Zp0Q4q0g0SDwThtkpmCL6Dy66/6KuTh2DVw7D81ayVvExJuvQc6Kj5FpwE
4doIXeIZbmxaCcHCMMPQhUT61O+mHGGdL1CN8++6Hc3KS5KSwUtXZo2/b0SVz1yU
JJophCixCAC1Lr6i6ej/Tid9/vIJ092H2dNwrfJ5ZfC0L/t/+9b0MIqnoJNd4IeC
eCGPTmyZxeOaU2rFtGR+2mbTNqFbBrCpBGakNAkf5PJ/L4lB8zWMm47D5rTrRwCw
LqAlEhHpMOt6ldKSKPqbTP9u4x9IBUd4rYuAXiINJlQrdaX2FPOaMd47FT9QJ14H
XOSJSuAOx0HmAKjxmBcwld1AnJZRHzSRFjuYm1aM8EOoo7h4g1Si/+umbNr47U8G
IZLhsfLRgbYJ+penVrgG4JtG6n9/g8p5CG3KOeX0wbmCRE/TBIFUCHsb+FuxtG4g
eEqa0jTLr3oE/SCaNnlc7KOmLewaOMOLNlLSmMRB4E/bmOC19kFA8kbBZ2H2KJ6E
78iuIWQKjwnl+aL4A5zKdM4eCz5cnjm5qbgJrr0uHeZ8OlPPxP3oS9IHW6u9cpyL
WXNn1tDe1+beyXnYSBerq1H1MxBujgXfS5DwpPhLA6vZUnkFNpQYfiWo9AaAOkfL
s7zcC1veSjLdnHpvIB6ViF5b7KEwl7wHIjIb1de//gbaxoUTls0jCHPFDsAGOiBB
4oPNFoPrL5foL4RodbQPL9ymXfC6USzCm7Rk5+ZmBcLJ0Itzsh2NdM7VoxhesIC5
3uTWvTn2GAeVkqdZ+EJolPA4oZH5O16hedRXYmMV0NfIBhH9Amskoss2lIWRAgxp
FnAnjYFliL6s9Ix2mDSk6wjjX5NR8J3tqnvytZU24lVbrmXf1bM6bl6JJpPP76Z+
OXu5RLdMeVi7s9UnIAszPo4fiw+ni3EuvkHAlbhDGHqK8hWF8la98+bysIkC5Rl+
ZOn/Ti8YWEJDcNc8Z4T/8iOpJIAs1VnFJW5ulbJRqCgqdWbl4tNfiwpWf3EIkwRo
inFD2AmTBzFYV/1sQ1TNm2sDP2EpxKG41UzWZRbtIa3+zlX/pJagLH3PNFZC9fEp
hT1idxQ5NVDtLiTe4BNGTFj6ggHjBi38Lmx0YTc2UZfVKqyIaR7rNB/RqqC3At7s
ikvqkvZBT/bCL+hr2m3ESKr6bd8A/f+sLLNJ+1pbmXn45/+0bsu2I9BV52/8QmJd
rb62k9UBdIsFGqLhnylboRm5o2/ejudbRcePQBl6UyUgWc4LywQUpo3iOhv7cnGl
OwiPjQ5RML2G5kgrYctGEq7VesLArnWO+kjlz+4rRRkukv0cANCyqLm9VHGVqW7X
l/snwTkFBruWH7JNCuwhy78K3IQ44plEiiwZq+tuFY3/VrlSh4zyEwnaXgvtGUq3
9n2LJepBuUZ0h8s/XkHDA7FBn+1AeEgQSr+1rQKdUKnIlMSsVrt/HvynlijHjqRi
tjPyPnUzWdmgCclAgwCiodml54rfAK/PKGchYmIeof3Qn11HIxygk0FDsiK/ab3Z
bc0k6TG+SjbTo/oiRw3JdwkZ9P8sI4eAigxY7VaNa5C6+BhIRFG5AwY7B84kDplr
HPQ3ihfE7R1Lcb1/vp7AvTIddn7bfO/WKLOk2cy9JGPTsosyj4kYCzKTTFmjcv2G
xYCFqVzZ3shmq3uJABTQPsYavRkZXDvI2ZwS3Kv9ac7dk5kmg2F5XNtlte6N+yZ6
I2tuWSSZjgA+69/OgX30lBa7UTFYalUU4gfcCMBA7da2/bG94i1aai7DNaC3TO4j
RuP7xRL9TiD919Xjv05/e5lT1CM7RP34M3/ktbE6L2yX/2elQccq/1e2LIG/5NEH
JAr4D5aZnpOhyvbNCUBS0sqV925iQcylFbOlfPwTuIcby5Tu/RZBdJue1gzfj27T
YyMvWW3zL71PibEZCgrM6ocWMB41INvS0z13tIWusYgQ6lOihpTzUXjUUXa9xoat
PLVHn/lI4rHIhkUk53VMnYderRXnMMzaKYdQiwr6ofahTipD32ML5R4UtCB+p35x
JMIuV0PXR6h8T8jyGQrx2DPCEp3Pmel1HGV6Jrlk6mIi5oEuf+mxo97QD7jc2YHT
kvdXMdeTM4Uau3q6pHs8h54er7SUXcmEQVJcsZIZtG5wAnB/3EpgGOmH8iSEFzxv
xztUoJSjx7a9+QPIPtPkrX5E2R5nnDmSaJZp0I1C9t68AOaMjPYfO7OGgAdKcEGI
AwVdaQzLHgY4wSHz4iVX6mqYR0BuSF4SXAJowWkvKnc07XFFdLNhY7h5/0ApBLPp
NaVfajKFXu0A9YAUP09girZ+96hxgvzcJXt/2aPbG+3vfxnzdfnnVxSzAGEe3ab3
fH5cN7lmC/67IqDIi2FLruSvgzNF04lhqRMPY7opxcZAP+ES/0V70UHCsgmO9K3N
5/vV4bYiohTTIMYvY/U4nhRG18UrwRJQFk1d5ELACIU4Meg+4mWRI6KhBB1kAqjJ
GN1WCsggPHc95Y+NNdNY9rt1nDtJw3RQIox14f+VOpCDIjzntL3i0o3J3QR9est5
rTpMRZjuKaiT49Avpx62GVPzsPDOK0coLnp0JXXkWjyYuQQeHpqyWj8PtQZKPfsz
YmZToICYTYUw+zfIe9N1qzxtrxof7AZOWMPRUkgPOdPpW/n/NXvkIp/JEfyLqcer
ADewoZqKHwEy8tT9WhVV/Z4v6dNCm6wo1vJ1dXePJGe5wgnAG3XSYuSXWxXyXEuR
TI94jBikoltOkwmAkCLMCnNP3AZhHqTqcBIT9gBogLXKE8sR2G6AmW4IZXc7onyl
0b9pj0IG8FKCm0+iDMW79g/mXmPUfKIChNoilLFhBMxzXJlWY5JYabfWs2Ekf4q2
SgnYWI8eveDSqicrWZtBMHuw66mi/iOvTRXtsIKEiK9eGE9FgsomX9/2HzSdKwfY
BN1QuQ/h/R8T1PXiV37zFkPOp4q+rqweGOx8g0eFI33mdBI7GW4vP2lxYbjKwq1V
ycLRsIrkeFNWGDY+8zNGMAHzTSstIG8DYG1vjARH8+N0fCf5adGPqB8tH/EF1Exo
NEVbMn4ectKJOnTJQDYeM8+5LYGZQarWMk3WhBK/2eh7bUTELuQ/1lM2K+FYK/+W
EJisY+jxB/PiSKN94LENZRA+Db5ARJevsixkNG0opFhTMvFWL8ej3IENBvrG/zzB
0EVoNCmlMkFv0rSUpX2p7+AeQ47/wF+xFrfQkjL6dnO/WjwB8FeTUeOaYHuCDu6V
p+HrIZ7/cyRLzc9F23hZ7xnVqAlcod9txjEy3s0S030fUouq4aENBIG9ogocGRna
E1N2PuivqZW2s7vuDu0oOa5qEgtJMfhVL/I3c2TcdUfIhsEW2StE50kU2Dk4N06E
p5lxesHhSPHo+KcOwAKekoDNpWHDeqiWrtUDBJjt/Uc9tYviCnH27ebrneOUDwDA
NJ/kmDCd7qI+CJYmH2iLAVlz6AiHMWUd/Kc3tD1a2iwKocCi9f2AHBot39yYkI7o
XScC493eGKfWR/rcvqpJtWgBxLNcKhIF1m5ZDEYNB8ygvffJGbn4L279cUzy1QYr
FXfDnIKb1Vq20O0Umox0yu7q9yYw2y3WcDNFr5fZXSigJEuEwhuvrduXB6UfDZvU
URWI2V9264dhCqbHUwlSzohOwXw3ibJoWDPlsGJRKYOe2Wmrh7HqKLLtNMyrK7e5
4kFFs82mk9PAw/eJdJpXU+VUVSy1qJdtD86Q3djngPksCy8PJGIQSKEX//bCbtkr
8ulAIUJcCNAVCneGS/LMOhSTjSNkf8vbllurO0t/eAKQaH31Upmv+0y/LkzcxZvs
iTo2HX60ANj9croVkS4fMuzserGOmyqOCrefHukODpiwWEAZ3h9Gcc4bBZSmBuEq
55AEtOaYYGJeBscjLx8YQV1AhIRYtsDJbNea2ZYImJO76sTA7FGmlwSESNiWAqpV
B6eG9DMcCOAVEt0y+NRagCt4F0FX9zEIISav9gA4vr+LHsSGaHndTA0BfuG9bd5m
+GJ1SmJHmTZcB2DMxRpKG9bZVBz4C+W70lQE2rkRlwALJQrcQegOaURmccb53JzM
6Q6uiRP9LBd9CnEqDMAxCKHSsbCltvgPyivTEs5FV8zOre1p/XaHPacyDAH9hta7
wnBPayo2P9Ip4p2ngweepYXwS/V4jA+TtjN0BBaosiF+MlFRavbUmsgTPMxmSUft
JrfXxZvzrbVvjy398Ysyj9KXmFhM2KW9KhlYpmNUabGBuYS2a15G/338mKk6kMLv
7PZ4YxsnLq7kj0B8aZTHx6m1JYV46AU+PgjCVKNTK7r3CNLjIv5S8SKUkX/9N1Ub
R7rtXf9WoyLaCBEOZdyK0GQZPiDSo8nl28cHzXqgl4CLk4iSgcL1vivFpj+CH7OF
cH5roSy5+zYmfdOhb9nWohsFsAiKtXyn5cFgEWPzDSSb+KSQD8RDYZbYLvgUct/N
sCY6vikhj7mYUtv+xol1ygHaf+cW9dBL2uIGXiTeVJMUFte+7kb857/xYCJv1Z/j
j4bPNmdl0SUGNZ4GNlKu7fl+A9gp6NdbxSsDZ6AL3E7dj90g7b2qG6Nref+65+1g
qVG7yEqSphgKPOpp3wOAHRNG4hNPih8Jxw9KRxtgvUVD25hvhoQgNTjcGNxDQ0zn
iU65v045LDpj7a3JNa1tYEylIqCGuiSYmHdCAmHX3E4rPmh5rsmvRs6RoB94mdS7
eIk4Usm4vLS7em/9pgm4fDjGh2zDPM8JQUUu1NbtvdENyhFBGDAWxAwJGkBmqZJQ
dE5QyUscqAbxMl/MjjzAx72nUaNCgwNlyrkiR/2E3zdKLJkX0cNfAJCnP5wT9hB9
IgNVcK2CcFgYFvVgfq5d3G1J062qa3MRzc43HpIXRRj8GZrX1coIFFsrsDc4lfyn
phSGd2xzrivtxMEZgFYgjcZmGZQb4WpBVRw3Z5XGAb1mkcm39QPQ0ymDPsjBK0gj
MXoy3PKBIgfdlDl0yMlxPJFe6el1sQXeS9zZVGIMXHvtuLNykBLKCtzmL2jXaXFq
X0J92Uy4lADpmdX1SI3AnFfb63I/pKEzXXs8W0Aa8jJZ3LO7jhmoUTn7BVLyhAJe
n/mrS6iV5IkhuJHxmGk6lVj+W5gaO2G6rhhM1oerXcr/wBz1Okmv7Cz9rHxs6JF5
LMGt9niy49vOHZMxPwcHcQlpyTsH9fjT7+JgR2bNFK8dyvIcims7RAlISIbzo1fh
O2763Dpk5BRDPGhSpyWXitWnAOtGnmtcVsO8UnP0Sft5gDVdH8MjyZpERN4lm/nC

//pragma protect end_data_block
//pragma protect digest_block
PaaJiUTNHZZptLV9Vj3s30giMOo=
//pragma protect end_digest_block
//pragma protect end_protected
