// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KSgMWQ9RP8sLUBWPnJsApxLONXyz19NujaKzW/ltIo4qkhPcW5wfHG9TB8wW
Rq6LH3JxLUrx9S5nW7Pyay45Cz5No4bKG9N85bZyGtdGlv2R7t3iAlT8O/vY
uHB19hyYN+wk0feqXkrhTx+wKXPme/fapho+eyhvOcTaBf7o8cz8K80/MfsU
130g7JQzp6SvUaze55Yj3SDc6kGtCsvB0FL7wZUzpySM5DMAtFJCVWSzEKW7
UAVEWWia8Y9QySg5/5EMzZhmvzQOv3fqNLGdQmt+lShmEr71SvrCMY5Hbv0X
Rxwn8iDfuo0L5OuQ3iCKTjzWdOWk1BEZgqY29bnruw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TvJaGY9wRPFsuaA0DOTyYwn+pgvaTt8PisFaUGxtaqdf/PQ0pzDwmMGuWfgV
lLtxaxfYNa6WoGbaqBqLAkmnNDrQKS3gHN71V5McmeAXtQWudyVebm/3HhsA
rpFswG5CJd7g9nzczcC8beqg5QyZuhFaevVsr36Hs2BgTzM2VRb96aQ58+J4
e0OUg71quacPZBLBEq4Tjs6vKMeLVa/KT0JnQfUVOrfnjR7R54tXjUz7pmFS
rMxCRx/5Uviot14ZmO57A4VJXwAVV8vTdzo0xbMlA3KmIOph68h7D1r9vnS1
IjcatSFDtMYphZxfU6C/1U+ozV3oB/qUcWEThXpXsQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fThp9gVKvxKvv+2q0281Pdd46of2x+WJmAtIP+7Pv3P6SwWRPkyrm3kbeNw6
5JNEfXwf31OP14rj8S5q7MmqlvguGaEHmd1EH3srtFnTxtwv33m1ZicVgJwE
hWGtt27wsn25wd5WmNWMapq4YKJQBvxz9pwB9J2CcRg913DhGjesc9+EtlQu
IPbgaDk4Gkk6v7zRsnIZeV+ZTurohrBGpAvnaCpc+wZ3EOQ2SOa3u9SY9A5f
kVyL3aVdu62i7ie1hv091b+y0tOtxoW7o8nwxX1wQkHv0e7pDs/8pGCIkw6N
sAKM953velT3z9R++xnhhI9Br7HUFJqq4feq5/IRYQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Snwpiirwofzrslg1Y5EnBB5MCCZovyNpwtcCBgZl+GHNi/T2BVP55Mk5TYPG
xHPPId28EH6mFZxyvf7bMxtPEHNOiNWQajPYN3WlKM35yzs/eTs4H82F+2ei
gsKAUf8CMXJ4EHZCcVZ1KCibDNZduFUkU8dl0gdhMtJBVnVGS0g=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
khjHT5Yc5VV0ZcL8uIp8/Kon/JEY1Dgjq3QMLr9k2X4cY+BvlMONtvDJ8EEt
wTdFVyE9cqM+TIQ9xGG3m+O61q5/ph/Cy+BfLfN+ot3uYmQPvUyweR8a90Ks
2O6m/9ywkOU69ueubo82t1JzcA0wTo08AeUfIOtf6pqO14FsQC2VhXGKUizM
W7dmR+dg/TrdDf4aTt6FhqbJly7y319NbAzKBPZvIG25dNHG8VefMxDC0d+x
WQ6i5GcocmLYhmW8sZ5EUjARA0luqqU4DXnpBA5z0GoGMvfLK2BLaybsrqd6
JT+GxLJooUS3EeGbMSOV+aYqAHeJK9HA+wVQgOtwbAx28W6cyQXTHlXPyKqb
wwMMz3olpFAbO1nAU4ILq33Q8Ug46hRGwGlTu3drY94nYCasGYUmcKn10wTF
9e0Asn/XkdsVKgVMz5yKKvYT5IXWFp5N5eJWpjGeulL8p0f+JPsBnDtQDkDK
ZD9mRovCUAPyPUhqpuAmLBE5bA/Gzw0Y


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P38JEQM7AWezjGw2IP6Dh+KTLUFSTTKyvB2cLO4IWhpFUbDqg+z0mrtcDRZu
7zq8T6pBsbmq0p8wBX1kFwX7aaXhN8923jbn7L/rCLGSWEDo5PiPg6mcPf3p
ncrg3+0Mh437fWZryGydK6UQG31rRyVWfuIs3Mir3QSJOix1Pdg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pQ9APHHvZnnkoYeQSynF0cCYAB3xrw0EjZyq1ChxadLndtdpNBdzMd9L6Ec+
DSz2EgLiXSSg9ojS3PLd6yPImoPOUW9Jck/U1zJQ7CCnihxFKHJi6jf+PJ04
uWvBYHTNLlLKiMmrUctKkAehQesfzN92bl/gzioGdtRLqRsCmI0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16832)
`pragma protect data_block
ftS5oPdAR/IKD9nud3XAFEtHKmehZ9HnnDS4gdcvos9GFkP9/o6YUFXb5Ebw
cD81Z5365FF0RafLQyj/My0qx4v/cRkzrq0OJtNr+S8EuLey68VJ5R/C8spM
dRXJXsTQhyYBQIMyWzoKGea6NvRT3KE8F1WBDiwkf1TuKPtQ7fsyAkR3skUv
puiqRK7KYrD1fe5tdeIEFNjK39RV3zCQirtYsEVHMGPsL3fRzKrkTwgugCkc
7mTLUEHHnqeAQhhbswpYzGYeK52LCMQhcMhbxr0mkvrni2M2UQnXiKj8Ktkk
TsdgRi51tmUAyHw2qjmQMLyDe3KmBVkDH+gz0nKOTdao+WnXrTL27KTCKuE2
D+6PUslV2JLUw86mqFnGHfia7+p5RVKsYZenEZBke3k3+tlCNgLyLoYrHqRc
CpoZwi+W7IgVcLXtuLk6qcDSKn9sqwlDbBpnwcTl7rzrgEn6Kf+J+9aRrSiS
8d10BGgmUsZv2/18QMJ4YaLJrpd4EyXJUCdVVDtBlhISYJdV4pqfJ9lFXYmM
mgU/SQ4BLIy+5cAJptBY/knlg751Z3vBz4BSQLikUfmoSClkjOlkro5sh/gE
GFsjI98zQj1ryeu6e5z7GTiok7M4FuOgtiaZ88uC5Vq+MOIY6VlzNOGXo8Sr
oGldxqyXflPKFSMfCNDC9gTy35XoSZPm6csXRYErlOvBf44gKCQGlX7VJFGi
FQ+bSFWciI8lNU+n8vS5da3K1Z/DteGVnur9Ym15ctlMmzUoDS1LlwLne9zn
hT1KH/ZpvjsTtBybu0yIBIO8Ui0J6fnA+MGpYcHhsX3hfHSTZOQIkujcYerD
LXowsU/kgV78qcUGWX3GEdSzRzX1cniZ+umEZ3JXxEL340GCky5IbX0ipMQp
5Voa87WUAxsM6+6yI51GK63ySflEC81NNHOz4UN/dwXWC/4Z1BACqLnoKhJN
7v4jiPbcueJFdV942nXVG0AjGxwNbVfT9varCZAHnyKQLYDvudJGEn7hCuvV
K2jS0coalZs6X1I9rjGbhRGlBalLU9LcVONWlp2G0mxUF7lE7v8+2AgF84AP
8yTRbmOO8h8Bq1YZZLiECuZ8xlsPjxmqLo3fMsd6ER0SukG+4ncytnvonfZO
uHoOlOONOQceYaOQC75BZKQek9n7g7dNHSB10UX2jtW/RtSkSGv38Cgu8JM5
xjCmqA3t2Vju+eaxVGsPipOpwpDjN481OWjxJw+4++MgGgKW4pV7jyawyxyA
vM7kqlDRhRyLXtg+LidKNL8TycJ7M4mhwa+pTaFZAE45bA+JjRbXC+Y8NR/2
0KXIwmD9HXQZcT8uRGRPF0EMIBJoXH/lLcWBXQuUMWb6CvxXlwuZE+uDWTWH
o+bij6C8S47PCtOngOLjTRps8yNoZubVlrYNwjckk+kFILJR60P895e+MRgY
YMDPPsizHBLqBmSeeRw1lnC2VP9czZc89Cmb6u9V6LSBIxI9eFKg6MoZTjtH
+mCQ4XH5baoTaHNNu5gWER8MMCSBGHErfhvXPlnqDNDm/s7gB3QLgOCJCAqH
9RcEau9q78Hg3ovwZQEWd8bm08ULQdv2YPfOWM2okCunpVT/r14rtXOCLnT4
zMe70DFW1Gn/2R4WzsfGfXCGx1itFzlugW3Fu8kfY0P2pLMOUVeS67r+BIIG
5IHeHaOEYSF/lQ61BRcUtfr9t7vftt+Yu/fadUKC94Xw5Cb2ShLEeRoR7bV0
H+062vKLO+IjzW5tKFMPRbJX51tt552tMsbPYzILDivhlX/KTvp0R+W9oIj4
v5QeLh9lEs3v6ck8kkNEvVtHfwH6t2fo7l0Mot4idx9YoLsYadpNPyZgcFKO
aU6WC1vexdIVUyItxjVGV37cI1hoVYDOB+WYac+chG5RkVrO7c0tN8QP+nr0
XEDjbXZLFgY7k9AYmavfvaFqyxckiQco30F+D6wdq8PChDdzkC5dijqt7lyi
TnH2TIa3ZgBEX+xza40mTdRwB5pVm16m2oubZ0vvJr6jGzFVBvQfGLXdTjLV
nU+GbetFHbflFwq/q2NmRfhf2lHYvfukYTXVF19bqaI5l0DgJQnJXCBf9SCV
ChbM9hiV5D/DoqIVCkC+oyA8f09S9wALnfXaWXyV3WX+lG4Cw0+Du2Jwfg6s
iI7EGDuuxYEIVXvJHG4068pWsY1oiMPdO7WsdarU7dQOsY8oIAodwxP219hj
aKZIjDtXbZ1NuiyWnFUmOQS/prRyb9onT4pKze+x/fCcnppdRgdU4v0DT5Ku
IdnuWULfqBPfVOZa+29YQ7OSXbLDb2xjFmAc8SqWBtiFEnsSYUckvxiqCVHc
raoZXlCg3xuFx91xNq+xhwBZYdezW1qT99xafMnAjzSpvgAnvWk/snyJfbVq
h+RykNYzTgpErOGsBUSANGaGMNOkegk711VLyfxuJOU0W418e8xE39eVhDIr
bTEUiJk2ZqcVRm2fofoJypEWV56bvFHWm1GjgXSNb2+UklUJUbZBFYS1YpX0
nzf/QjNSsEC2ZuCeiW5n0EkCXqUGUA2iNIlYFuXl1R0+kkE0KMYNqZD+5Ohq
JW4xa0vtGh+zH1q8YLKmfM+Z7ggFr24WvuAnDc5JMs22on2c0c2NTVDKDMT9
dIlVjqje/yEp3t48eKZJl8XxSjNQVsuoo62Z3anPAjGIsflZFB9nhtHStTfX
H6m62vHmaSA0IxBCnhJgqWLpq43kxBPjYHCJSAhc1BCJn9bCqHADN0JU2rlD
KxXzFuiS3FoXNZoYRX8yJjxdMctf5NU4yCtizpqxz5oRz/VER/FpsCVQJyn6
Q9zpwz/xtL1x0S6NWzwyc92x1P/xY2LFoZnXHrDdP3vBlrNNA2LqYqC8HkxT
7ZjwtsHxnYSe3780bDPtuCrOEYJ0bsyxusU9MBrJWAzL99Tfritsouq1bidD
OVgg0rAep3+Mu1MCKoVpneNgVhn/Q92VOWTZqT3f4VSIH5PqoKMedmhCX3ea
TsHNRK7TsR/d/sjT3s2LABIXatbM5TC9JxkfwQvaPzjMn8lW4UIi4F71spYz
q9rhGGAKk4oBzUIlrawk1Mv4jhg4NB6Gf0qPo6QY9+i3vKIC/oHrjheuK8HZ
Bg8yEqqF8QaC/ARg41B/8pB2HCbJU2AWnWY0ADyjcQYvAVJ/MAuW5bBj7SSj
GiueDYJhsj67dmgfJJGvSuuvKKjhO4kzBWo+el0fbWPXNXggUNYpIIxOm32U
Njd+65iH67pau0WriB+WoMGB5KVa3J7MN6Al674mEhUtAb4lyKC+wXI/JUGW
Y4w8dgzarjF4fU6gCvJmIi0ypfVu7Z30ArLNegB39oezKK+UTWTreMtIgS6R
Q6Dsh49fRIoyBubdYJqklqVN2HotkuWjThamzvhlEXneFvc9Q7rCCBi4BzTC
d5hqsz5g6+yET1Oc/53xLlhBH5SljfqhDZW+2GQj7iD1eRyPjZPPUGJEyMc3
SKCWodJqKpGr8/+vW5Bo2yMywYrGQxauoaaN5CUk1aRYkkT4Mtxcbwt0rkDJ
uQW/0aa4wQcb0aHEoaHLTNLqVmY60bniW+xapsTJAg07wrJxH9AKhf3lbMUU
Q1iS82Q1wfWBfEHH6UptOh61RE1h/8Brq7Jyb9xSXRUhHgBC2Uf/Px8Y8eDU
PAhAgiKeu06sWLLORLNQOGCem86NkfVu2ETn7iGMOH/JJJUmAcIr3NrYu4n6
l/oBzdLQ4YwPRdtOTukJFVtd5BzGmkkgfhv1WrQuTQRqbS7QoTCYO0jSiYyZ
eZJL0yNOMLrFXc1v9C6B0nfQMgz6XWTSZUqi7gHV5Revgon4DnSiUHR0EeWr
VaqO5A1cngd0cWVU9hzjl2TWRN/oPB7ZVxsCEHwOjYEac2PKAn43C7kTLmT8
2ipFccC6fVhfFqqGtj3tyRFd5IPxLVNZtvbQoOnj8ti+KSdRPy+rU/wmtEqS
Ng7HbwnKAAs62uF2fwh3XQ06Y8vqawx/WwMNuscIbO95ehJDgJ4eqQFjVPlu
61TPwYnSIZ3P5XrH5/DE7GU9nEtop5iBB38fHb1JxZM+dcslNTpmPSuB1A5c
DKZMWYsyAV96EZTdqhHs7nfVsu+vpCJkGB0c1f5/GIW6Bu/bricgb087kAB2
sTFWjwOm7dCga5JevzMblPE3r1YjkI0RDMSspuzlWigZ/orzP4q2EYNp76wi
IN9K6dCqGQ8Mijciq+1kIlwxhe3hzmBNXNdyErPKCoF8Bi6DypEnC81+49NX
1yZAKSyxCZZ6xtuwZVXx8VQJX6k2W1KU7mixY4PGy1+7BP0gXyS2p1Jd0Tfu
k8Y3B5/AlbB2pkKp+tWqcuiHjWZVUFDGTItcH2rKR/V63bBBckksvogt6ZL9
svJSXkUMSdab1MpmQgXnzcGZ2ltY8P9OMhQhfJ10ke6eliKPj2MBo2axBBX3
9SNXNKz0FF6OExmpAFfpJ2Xqb6mmG3dMFmdMpgBUo8PCJURbh2cMXeTqIqPy
OPkPWXZqMC/6nevaW90Eb7SRMCcAs8D4SQxtfjETOo7EhSwf+ifZf/4WpxJi
Qh3L/TnRZgABoV5c1eQRJbuJ5ARovUp3+SJR1HQW5MFbuDvXPSz/riFlvJV1
FCDpJEJNSez6Mg4L25/tHUGOXfupRefd1oCAZ8N2EGzWIrJnRE1SMOpYuy7G
Tv3k00KUgF8N0BFO5KI8yHpvSDCZ4hdBNOngs7vrNzt1TY7jXA8WfTLtoXii
XJ83QIbIBhH8xxo1OAZTrOQ2oO1mc7SJQNCkGfu6Ugk+8HA7nU3gPhbeap/G
kkVEWWKj5exObZCo7l9GsI0uA5UCbT5ebzlfzXKd/vQmMxkCZNdDZ8OgresH
PwZCdGFrIsB7XqwxwkbQCW7Oc4M1iYrzYDD9YN4eNFxCUn5BjuSzO7a8lt3i
ED4VuETxhoXs1SYYG4M6tRbxepraeH/hjrTPZY8MwpbQFXrQp0qJ2+z1qoL+
hDNhtp0h7DNklrfg4xI3Ez7N7Dtj0jciag5JDWzLoJ+fhfZ09wOz4qs0FLr8
NVaeGeTUvid6O8Ih5Pc6k4YuHIeQy/ADmBdGsXcVVDrqlSgVS7JT5JGlJqwF
JNZr9hV7D1EaOD0uD6aD8dbq1qQEHN7Hjf/gbhXAwJLRg7o7D4v44oP71Xwz
0sameoGls8nmkuED2xAvszdtzUsUifDShp6xEM+T2GhlXtIp6TozDTovodqB
C1WcAPbSbvjU2JD1XH5xgdAZTL0NSEY2OEitisEhUnMwLE0/eCSKcaCzXT7O
eRlTCNfzMMd7aCt3aARmEwWuv1eIfWlk/bB7GHXk9fUwXoennHAKO6whSBdI
2HaodXDZYuvMk5R2GXqsco5Ey6UJ2qA3qGjbP23OtPvQw+NKAjy0li9L7C6u
YM0DuSZX2AkDjUmovBRlSRYO41pH1XD7+cttkQrE5p27Iw3Nq0hI7FqZ4DpF
ei9YJ7RbHTL0HJ7I9QPCc8JSMfc+qC2bHDtfIvViSSJLeGyijyroORjLK28z
xydYBZ3Son91oFc8vQVUK49tVCqtU62f9aqhPUyukPpFROsLN20ABGSevLub
lFHeO8W7bSv2sqRkITgP/PfglBM/GBZqWjRyVhRSG11P7hvVbnKIImMSPNP1
v9InrzRrj1Fn8l9AfYtVYZR2ZcfHc01XC/jQ+/NEFgN8SJRT60TBg2EZaqxq
kwDDKnKXeLSSXTwSyZoydJ5uKAqDL66eVIueX+0ioopv7XW/yk9KFAAI2G3N
7pfCefeNt9gfKrRY1rDe/b+MHNAswq6ClOKQao4uGBKauGZgAX+y3RM9IjAE
oQSF+VC7p1pfXg+cjyTAicKk6UGUG5V//b8KXzqWQaUBjysQyX4Mm+1/Czq4
UzhkiYnlxlpr4XfEM84xCsX6WZ8tNg81URESTmiUeZxGCUKiUGJIWd/HwsTl
rNcDqcr91kl0M98JwrWIhcVegssdf4yq1X3C4RCJghftlorYojri6dEc3DSK
KHD0pn20eEvZWjKE3qM1x+MNnvV91y0HtgftFJvnAzmZk85aHhYFhUWNh2la
2TyKwwDajoA4WJg1mEopa+FpnnrO72EbcfTDZIZgewTL3vrbnd9vSvo3lri6
RVHjirk8iHLm0xom/JRBn7oNPUHLJMs27U5BPdxaIVg79cm+UbgjeDJvihiX
PkOSoI4keG+E1QSUWQij3OBhlAe6tqlLDQY6qCgqK4K28nF7U1DbrEfmbxFK
lB4feMJAScDu/lTXy0lCgftc+bO7ZEmDejqmRJkzfyYH3gNIqO6UBdtHSi6g
cf8DsJOOK5JLRj+nBaYOHjxkMDUVid0cQlMqC0j+WagDecQrBv6fZRUfK2Uy
jTReegIsxzaxwIZzx1FTWnhhnXPfQZ8JfGFWS5F656p6G+manjfHEWsOpevW
PwYeyLumNs+WsdX5EAsGfz0XqGLD8CzxqX1iuLpun8Yi+/b+S/r4vssD0ved
N0WlqBMzYs3qEKGoYlmBc3h3vlUXC/zzp7yLl4rQkbMfJXAuoRS7ZLvyfxpD
ol4JhaMUF5BfPT5PfOP3GTjhi3JEMu2+0MImyV3F1oGoIVkjO/kLuTds7Kf4
09mZ5ZUc9IgTjTTe9E97KJj9y5oGks81Afg4dJehct3aW+iFnRZWz4jMv5kP
TNDRm+ywUAqHamj9ZB1rGqQSUu0h37LgvZAXhABt07OtUlYOh2Ff6r8jcoeO
BwigxV0UCfj9rGFqrxcpgyl1cdauKGpNa2dfpqWoejgsapYJxMQNNC778usS
SEWP7aFoExvLbMUIcfxtLAOY/7TKl8+wUAmzdL7LDQgD4YD4y7J8jyrsf3Oj
OWOOy/GdB4cv7Ql144lXQTYJxkTSFcNVEap/LCJbAltiQZl1E87N7USpuzlv
Dgg1hyyIgHeRYrMnWGSoGlf45hvRnU5u7Qw2qHsNt6wWwAphnVVP6kGZMwCC
7VVUtdfIVk1tsb7zoAAEyTvRko8gNorx4geDFRAm/5EgDXtRPqZ8Q1eo+5Ey
oRZPdGPjb8OepcFu0d1bfM0+Vy3UAQUVrHE4HFzqvbxZFfPPyA2EgRLkPRl1
sI7mDrun1CNxcv6K2XBTdZhvUsbCVu0TRCn1WDyi0UNkIMzy2Zgu5hO3DFY4
jFToXOJV+EYGK8N38x/aAaLTbY9IzU4Q7dqz7SpQQfubVmSvnvi7LiM79nK0
AiE7ajWBvmMyMfywVAgV3yZcis9WbRckinwS+IqXZ6JHrnIwF6+dvf9DbvUz
oY+dbI5y5QbD570KgNH2SPiioldINUyuOqxYcrdDiknvdOUg8mKc9mhRkrFo
+lvbKtzmJr3Hl9A0pWYP2QXDl1xMnuUJTyjpwAcOPZXSN8+Hj13nCKXQvYK0
l2Jf9W6ayQc1Cn45GswIiyQWsbIyZDkZYd3Dj1n74yUnJBa272rFiFwOc/U/
1t8L80oRnrMR3k+BoVDfYE2KrXXdHNDxTyFFWCyBdhpst+56Y30zkU9TSVB9
1a/xUqYXz1yoV/UpOgEuAW5Ix6RG5GkS/YzUrGsvezsiKKGR52Uo8lNvix9c
kogxuJ0X2oVeGDoYNLfHtubMAhu7Il9ndyURGGUCFWidPf+MfTF0B4OKxJuZ
mXkBm6ft2xrTebEIhs/bC7kwSWTgqu8Gn1L7rztbXMD1x0wrTXg23r/m8trH
38AFey06zrNJOWskR2sERHQndGM5D2rqnS8YtR5JfxUR56bhT1yn2ss/1jVW
nCcGbC83o3JwRvVCsF0pat+pWrD5GRczQTCzWwlanGpLll57xkKtx5dxcMSf
eHSGTRx0x68B+G5PWHvKJEpvMzYQfJylPheGBlAJ+VPK2zhzFphw89HAxKRt
I+bXiSXXgIc4T4yLDsTZzFHcSq7nF66GCyOS3SMAN6hy+WsHnBneZOOq12qP
f1JRIm1xVoq40iCT0Lh5Q6z9G3qRyiv6LUx1rCeafPfeVLM1bzF5hcZ4I+Uq
49KOSdCiDFa28HaT8aIoPTSstDD3i5yQva6emOEtTSt9a1WCHjTsE3aCMnNM
CmnZA75B2PtbT10WgTm1LrnV0vwnRWEFO74BwCexMHGGbCr1h5cnb80aimaw
Dz/O895qyq+EFVbArYNAAlqqMl61sRLZEv9FTlJKtQgcwZwWyTsion512Dss
c3zB5n0971kAVvu9UVP+7q1biRvRgQfcqnjjyTCbH1gXhdEpD1zTzLMwO818
SDLm6lKfoZdWXdLlkp6nkuIKzHZoz5JN8VCbgewGHvT2EmlalQnXYTLR6z/b
8Uw0/2uTTCaSBbW1ZPxBEULTP6Sknd5n8lz563AX6Ib/VfcRutDuOOmVkg9S
2cvVVFtSJKggIYhudqJGz1JyMU1VvjCizqeus9fsTGRKsuF34Sd8yugMxpKa
uNcvYnCWc0JZcwErBQXMEldjE3bor7jB0NKK5vTpSgxXx1Q+v9OElkDzo2Op
ABXAtqRVMdJF63EMsqozXLuRXQMGnu7RWKR3IImEtKmsMC5GjSR9Nojdy0+E
KaVc5QtML2xxZigCaBO9k5qwy+EROOIH+zJCkLGbU4u60HX/rJ1dZfvKqOnC
nJ+yJw8Hbd3PneZIGeJueBzx7B7BA83k4pmsU/nIrZ39hPcXCLqDnIz0LcKg
dKf3VYG0DKE0yuXLZve+jn0biARerPOGtO8+FHvFfguwZ+MALaJfewO6gfBr
2PISMU7OBC6vTavpLpoOMPTWLO2YrUHbysgXtxLbR8E43bRZpI18PB9kmWRu
BWD9QwYFj9H1QiXQ5sUWAN6PSr3gUkKfArNymcnwq5xEVfGfjWpvIO2UTCOR
FLL7ccdeCFn3rTqIIkcv/NGH4iDUVV870W7OK2j3pRHX46HjmkHOVncpVyHL
npmtL0efs4VJpRFMvEcOPrx1EyS7hCj1Z54ou3OpXhSHutlNtnuHv0w6s5BV
IV5t5CBq8edD7BOlX3mp0NY6a7AKWdFGdaccfLmmJvQUKFMQT96/9jmDpXu8
gJnpkZL+F4/AhOUgY7is5wcYCdi01pnQTqdp35PGLlSjBOItCIqT1BkgYlTx
Q4eT2FbAy6B6hQzM8hKJ+o1PtZOX+G+azjprWptsIrK0qu3jsXxJ5eegp0aB
67jHVz7E2dFF9CAdVGXmy978GvMUy01ALW9f10brMc+ybDr3k4lumKtYhUYp
91U8t3G0XQ5GHkiuUI1uA+6QJSgix11AbFrc5OeGToPkzs6YbJjW6xonB3QT
7mOmsQJ1Gb2m5LPHvZEDLMMZ6yO0S8E+5qeRnOeti09fpp1/UtVgyLgFpQ8P
U66q2m4xMPEadq2bV8ymY4i4JJ6bSo93l2Koj6HN+4Uranw8QqPrZplMjdOd
QkEDdij6SCejptrGKzx416HbrfCQj4Jh/2aNmXjKErv0XHfMNNDCZbOZXlUe
eNG3BohXY841iRTBaWrJViw/R1UjTSjaI8/u93REfQ9ZI0dz/FtAoSD1wbzD
SKaA2/PPE1NXAgcCdDjzNBIDTPm2UwX7Zul5Z9sJacXkwcszASZ+zaCKrEx6
l9NQkL44hIvp+XZ/XRPo5Nqh8xcRW8Wm8TDf3Vt0Gl2d70ey3z2xWoR0w0rc
TzAoLgxaepArOkHH7FHCMDemptNvQ/uw22rCb3xpkTETRJTkw9J7UOlL1M8b
zbN8TjJt/reRUF+R3PGM/va75iVQ6Nx3EOa07pcRBjRGHBIr24ad4wr5zpXM
z9mhQikQivLhaZ3FCarjKCxzosydyDZbd9O1PtLEE6TH8+c32AfouTBHX9d1
87PDDvuAorUYevSvCScAOdR7pn63vc5HpliI9BrHmGAwMKm83TJdS4bRA4DH
ilyhJMWEZ09UtNZZabwKJV0r78KEH6pfCSc5PK18AF2vL+gH+GphbIFdazlB
bkYmiL6MClj+BDW7gvDvGlwV3IZ5QqhkR0RkCmFtg5m1DiQcqxP0SDJQNS0G
Q3DymGuBe5hMWzAWkG1uJxPG+rOkimS6uWgUW2AmQqTuMDZxQeVKnU2MWAVd
Zv8zVSMLsVTdce1+JaL1Sw5Nath32Zjri8U9MXvNQnQujOMtGCInkzlrWFiI
zEnrIxTOpRMqsfooTH0Hi3uY8KmdiHbfrvndHIuWwdaBKWAl5vFfZLXMopow
nKSczrsLHPT+q3Rc7uakHwGNkKk4oDbsz5p9hBZSSqmddsPdB49RJxg2djRy
Gcna44IHV7qjNePv+BiirkFXvx4ZstakbI/4WO+veJt19fNIakYFZx+rlKFY
YMGd2zOUnvwHkxlh0z68WnFnKoRXzNfll2+Vbhlf3tNW0Bqu07dWwHLVW5o3
0VG8WYa1CRaBQr7/jXrNVBAtxD9U79Mq459EVymDlOtg5aEmFFOLwJDNhdDk
sX+KA2hYYKgzlhiPZaPFnodcfdaDfI2or23Olxifgka6PCoO+oDMIG1O0EkI
9FaGMd2/fC3Pk7GBKQQpC4Qd1rjsPznD4vbkGmNMBRlHbCpcNcv1wg7LmXTH
7l7bgF9YaIuAhiQCdLqlbu3t65u6fJMyg4PUhmXVH/I0BiD6MFwmsRyIQZ2t
aEeGKrysEkz0JlbacEsi8L9nHzth4nJW6oBDIooIhfNagaDv6A41RWFr9ZMs
b8rL+5Or8+ONk6ECq3BjX2ii07Y7mrQucP0D0WNs5/sn5uNNvWN1FdvKZn1b
7ok2mLx4TauWOZ+iDDd2aq1auThm/NfWQk67EPCwesKmmGcAQrMk+VZ9USwA
lhqdClQZUTrfuBO0Dn+GhK6eNC6LsoFulKGuOL/TpQ2pG57J/V5zUc1i30dl
cq4rvWYgCoe8iOu/nxY6EIV/lRE0Fvd2uG7rXSxw0uR87Y36zg/5GiBZeH3q
nV0wSpctc+d/0gih3RjIUClOZFYoWGC5sk+55ojP6TQX+sB/h33T4uWHob93
SCyxf4qJNSGqnfAATht5ygAYc7UmA63gsZZYmlRFT8B05rsBaK5jOiqafj/F
atY+o8OxBO78QVR3VcF1OxHuHn/vvjS7kurAq8hC3xXS4lPEf4gCvyzB2Nrn
miWmeHvEixXmPXCn/FowMYX+AZQ2UfcxZDVabUzhT4399wFUHJU2I8I7Y+un
IX/jrvP8C5Xz+vUc+pyMeC1V5Hx7/fFguKEFN60o1Nkxa39mIeTE26gwqH2I
QRx+nzone1b7gwHXWjiT2FyTvBpe4286Rf1KP2RBk3zaxsILt9QVdYbePbCi
yIfMYjQ5NGOPXq41QdezTdvcxLiQUCFvynO2mpOmTbHwzyLFohOe7CZxkQkq
0+TRsfcvCAEyxfBU7VQz0afysSC5gbBCTqYjh8pEuWsw07WT2hsYgt/OSByF
mN5DR9fsG2WwewyOXYbSqfVvVU3BIREQEBhn76YrcsIYqRJj0dyMtamXqe9m
KkrSscM6HT3ymfl2XV1YiZaG8o5bpCWdygdNETTJgbLJLXrwnm+rQmTtAEfV
TekbmW/7uMKJa7IPlgFYO0FWcTvPPz7801V2bwGWakLkeTCIxEI38MFGn0if
oOS7Z7g2hOqyJ9JOt97ycYPW0DycWZ/wBElBXot8A4z2H4f4gug0Qk0uq9dk
hRveZanx8fdzU2t8vjCNW2vtcFKECpInux2dRLsh2RIYSIeoo9FQ82QEBut6
g4JsFtLgjL04CjjZgdS3mddPiUPvg6Jkh9m+GO14HK5ejgnO9k7OUtazjdmp
LFIcgdJcXiEE3L2Cx1Kyr/kM+bXin1ldA7f6Xtm7XoNXAZMMnfpykVcSNqAN
ArloS56IYg1P56FQv0bGLhSOUiCmMqRihls+4wAVX6xI0yih60n6w0iKV/gx
9/UVNi5JIU/rp/2OprbkpWTXFzSN0CSRoQwNKx9HSa8tcTwMGPNbRmRb3xx2
FkafFSm02s4cek9aoEXM6RqQsPX1M6ByuvNTvpisqHbkV8YShTK1/9hImc5W
Hfkhu2WTpDPQb5lNuCHmpkq/cAkzPfoKYzaNBZ5Ee05Ls1mt6BXjZX7y2lBs
MNOMqo8N1Ee+EwoKLRs8vWBflt6x/Suy6geA63tixRO7sxvwo2qN7yxqqiVf
Vw3dsf3cIEktHCR4eS/umYPIwExRu1srQ6a7x8hhizRRDbiec1NJ/EJZIA7m
G4twnyCJWTZFtAkiVCY4W/eVNwp23jpKwg1iPY0pjirf9jjkInJ1U/OF80Z6
ldRaE+N0dG5ryJ5mgBM00uXHuTBBDS2P8jTFMgLSyiHRCSCENhafC/ctMNn8
tI4ROinHbLCSNa6fR4dK/s1/ujdWtz8bjmlc7Qg0Aa+Aq2PUiZrubsvpG0N7
HMx66y2nwWu5PVZ3a9LWN292NYRXLm/r6CmkPEMEDgYTQHtgvOwH0+5CqziZ
Jq28LDI54G555bRsnrVcPIoqPuXc+xe6W5p63e4J5luCTP8ZdP8ToHGkZ9lI
H7TclBYRb4jzS52ci9NnCrYG+JDL7gAfHaIsLfomwe159qRB6+Zg/dr5EvCq
OpS37Tqftl6LzRJQVmloH6/nYtfMyqbISZwOwcCQ1Ovj2ld7v1UL1UUqjvja
/WS702FfXQSgJubCVUCjEg1x8LZCLt4R8mfGkW0xeNT9jzDKpraYcGQueYHz
lVoTqyLcQaC/cPMzim1MYRu0X70q4pR6pr7g30oW39Gn7HLkuqyJysBJHA9q
xjk4brfAkS+w/9+0KVxQP2zJwPMQz5e9OUXXcw4ALIVYuYB6HdO13soqO1MV
prPkJQZZTmR6oI07oGSY60To6rvmjkJtDVN0+BK/u4mC0OLIizuboY1sMilt
/VEqMf/XqtaMTmFuG89Ap9fQaFtC2zw3tZBHUW2nHCKxVr2p1grr/WaJF4rv
H2gq9f/mjOCokkqO71SCE0WYu0SMpt+3DPVxakoUoQsrSvEs1+VuNxDK6tjW
HUv0W5yAkGP0q45XDsPjjoTww+CIFHDN4S41erxS4TgQQy8bwBNB+dhv3Qce
lQlXA4uls+DsZrqwPqe4p1FVAD+8sa0kws9jtRjmUMMay+58h9L4ja8BnXfL
lx55rZ3Wac+xjLzwjw0gC/nKOTcWb/9YLgljfys2SPCbr0p9h8W6R+3dkPQa
VOyf82HZe/LV/4xyzbaWQn3bwp4L4E/f1tWSkaijcCnhO5MeR/h3jsFoJAqt
tWH2IZmAZw2uPI6AFnbLFv82Dv8h6b1rpvZkqI4PTdlfBUz0aV1t1pFj+feD
qpf4v3v8hWtQuSTdJTWEiSlnuUaIqT5RgJi0aanIOMu0wqRqCdONP/rzy6eE
1k4ycGTLuCzlsRYf8gCurPine4Veqt6qtqwXdTre7LER42wp3RjsVQILChfq
ooMFFa9N92f2+zWDYS6+9RpxOGnYva4QbbfOGsw+AUMcN8OF89p9s/wCiOws
LYdqweMl1D63S88sTHvXaVQEW2yJ0ZhN0dixqn9es46sUMR+VU4Esg65xcno
uQrQfB8IAR+0os2cciAxoBIzqcpfVBE6+9j7iUizK8+Pu+LcvdayAHyp9CrU
JFrJsn7XZXtEAVY+vrvP4maGuaWeuZ9mtl637tRjb/iPC5KWfkQLlBeM56bn
Nz5TNa54RM6abDCOHO9ywiHwUH7uBDXzcRnnYPPslfp9C6iOlKJOe1xjSB5P
PAHJcM/NSOFs/Icz8ElPjoozSfj/bvt4jAeLe+nbBVbdykjxq84M+8GdHEY/
sBf7VfZoG3iWO7hVQfjqk45B9W7W5WvbCJsVzv6lPhjTM4anwqief/iQXAf6
qK1lTZVsAn+TeRZv3IU/8PAXsECeOzEdB/XwtYD0s5mb4EjLBpee6bU+sQFT
Ol4QT7cfgH5qpeoLsxOz1Ledf6ki9SOd+nD7DduIHOR/T2Bw4bbNvnRyBfVn
pvw7KIukg1tUiRHD2KYwu6uXsHJtdNMlrWhVfOinYs8MoB44LAyg4TrWBphq
f1Od8P99Wp3ebyuJdKCwffSIGbhyI3V+sT1nZnodbPYdHGf78u/zt5yF3pbT
6yBVmbWVlRD5j7FVR2a6b2BZ0GUNi3H1DLtOo+5jwsXbfwFplrx3kBd1TGKG
4XpFBqQe7v48aGs2Joq45L8KhqkvdWfkiZo06xHJ+6hDNxsuc6xSRpmQF8+g
CY7Xviz9dTbqAjBl5EiqlsFEm1oCpoFhnNaJDeGfPTKNgOljp1UxCMtV2ryx
u2JUBMzHQx1L5mpqySdSD4he6jmLLiBBSgQzcOFhxLB3ASaHQTr7z8ikl7w0
X+NXRfNWWjCo6sfYd3qlPmwEd6mx5cX9SGPCuqhn2lBFjK6bu7nvT7OVvYYN
DGHB699pJ7YUo5imrVnys/9KA1GUiJaiGWZ+w/nQlBOiQxzsTx7zbfF9DV3m
4Zd0SxpDWMuDdbpOUMCJyhJT5Iq3FGRSS1s27d7c6S1HCTrIFgXzmnOZLeP2
C9C7SXDNMhmyai1uF3wy0Ttr1I+ShhY0V/LckdzToyBcK/6A1bzioKtE7VgZ
kvHAHVYLgikQgh0rdGS37hX0IIuzNW9s+ODddnnnvkIN+p8ruCpVtvGE/q/e
v7TSoXT1JvvvPVARYIVlJ7FesI8yFTdK7KOMtZ1jpd4ugU6Cslo9D6iU9DvZ
8XLhAlqT6Tl609Toyqw1OiMh4JZGBxIaey2MvpY4SOVZmxKokhNbdgQwB8kz
cai+pJHRMaMm2mcZc5ljU6Moox2Z7RHsCTkdHY2Hik0zr6n3V4KxcnoTnIz+
lYYZcJgZZbOfs+ks3YPSpWcjm2CL3gh4epHeHc/I+dq/7lEM9SAMPt0iEA7a
hd5/J7xirJkLw1R2oTz1+BnLeIBVOOO+M3dnNkKlkcqOtgQSRFcjeCd06EQB
IFAgdCFQsg5Xt8NKIGkec+4BACvCXGNizDxtODDFH/8bC8nK4q7NDPoxvzQv
/9n/OQtCz6zHlrEZYlsJsgsgLIv9mHXWiuSHOaVandkjrPiTLt2H+2cMgRsi
J1uBot/Bt/uD8lB+ONA8BbfeICFrkDufbsvHEci/qBa/mU/ruAHJ1ish8gT1
3x7ZJVnmoY92WF0dhXSOYo6ou2VTd1aRDg9myw1PaE9fBlH+z9EO1N7XB2E1
P1l01fi5jaS9oPxZlZqAaYuHoEVGz6I1iydWN+ewwYEaMzbyq1egCQOm1fA0
7dYu5wkg9MOaDwP1LP1vGUmrV9b9SzMTEsZHTeppx80equMTg1A3K0yWQNkt
X3WcWYM4r6YfBjoJ5HhUVzwpaweFQFe02vlKSRA+cN0Wa60uXaX5oiU2X5t1
wYkZEqiatFI5dxh0a4aJ04ZXbdASgMO/ueToizF617zRLZkkytD2J1OrFFol
f4Yi3Z6jiTF+/BvhBfe+/DXlhDWm5TLptRouTR+cLTKv3teJMVl6ArxX65JQ
Q6uUo8IP5HHfbQSJkGKncQoecoApYvkgGC4T1FANa0JJO7zrjMRoDwNIx4qr
joo0QDoOwQEfyOsVRdxXhb/ufSK8xu63F+4iWuPmfzsWe/qDztYACuhqmBpt
VKi8RsXOaDWFbN8XWYlu50+z64DmdJHo1RGByGD3WinaTVsBTXnxGxDPbDDR
T6vNpHu67BTFcqWS8U3O57Wg9wkayouchilz2tno1u21LnQj4UU2VGJ9LqCp
HA57cAbjARkBVBGIrqkLRn7SuCGXYnjNikKc0vVX9AXYZcnmHonMuWoqFz+k
6+RRl7g/1hfa2j7diSJIPINcJJtxBQc/UrFj1HCB3/VK2sXciTpUK6b9SCNd
IMyHNYO0oggRYOMlUYmHIke2XrJhRZz2P7JrpIVFCJd+TZyom+m8PEi7XtCI
XW+B7bgUajoBSkFs8V0dwax3cKcYaw09KGNrsQt7TDp0MlIPv239bVjQGVJN
xvQ5rfxF187wWlN1Ie/1AgiEBsVpFBLNWKgigBF+3eqVLnVgNdCn+EDJZrsy
wr6WAuIh7BCzL9zMe9IoU+ZiFD4MvaEz7B/gc6mCjhhm8K3kh/RiCwik/CSU
3J0kgLgumiwatha7uAm8MNoDq37dljBRM+c2vUIoBBUYn/Ozn/HeSIqDRO40
KQbn2izWW+UBFuLxMDn1Q8fMRdKNho0nhwAvkPSAGz1ewCH8tRf+4tFxLCph
8yqpjdB0cOKT7RPQosP3G+F1NfP6ZmW+8d2oy241QWMGk1CCH2g8SDcuk+gL
h/soTNyC6sKQRt2IPoUNdB9CUXt+hDUi61+g8VOpt7qSHLM1RtLSdnwZSKhw
Sp8iAG4xdiMItmcpMyGfOEhL88CUR2i6G6mm6PwXYm3FQDEvcG2y4P3pH60R
UGIe3qt9UB2+B84grBSFixehJky4M05YBHEDIC/Qs1hVEIQl8OzXNboVH6b0
mwCqlbH/r6dGDSKEVChHIX7ayi85o2QAnv/+kNMUumxW79G2tBIKbNLJsnLf
uKYtQUxV21OSNFhBU8pMfisFkea1OlmQrvwyWuxt5zAEYbunI8G4y+4mQMBG
cgGXqEu9erNi0kFpI4UfEC4kd5NTPReu+aLP0SKbWQoGyjZzXL5PWcgMXHLB
IfY92QfL3KthrZ2+14WWFzW5j6lRzwa0dr0JTMA8izWphJDuVkWwDo7sfy5C
ZWv0RXYND22IyAB6h5pDGPa4ccnNj4nPHzMIx34nR0DQqkpsOBho9RnrrZj2
SNwFkpExQ3LTK4fUuQW4OpU2f49sij/jBIZcBj0IBvsy4yeLVS+D7lY5pxlk
Ia++P7G5Xglb9bqTfCEr91o5yvV+rg0qXPdPeeDBkQAv0bEgvF05WENidnYA
xwqHzlG/wmn/S9G/oEgUl8ZPAepftRjOmiDUyJrO6FnKakUI0Yyc/W0WiH6H
s0ALsruTc/dcPEz0HyZEhhr60HmzqkzI6Tz7BDYxotJxCqkZ/Yj7GsRg8PcX
NXNsSfwK/ryiOpdD89WoVT2MdF0vsLdRMZLm/LcAexWE3FQiX5q4EdopFJ39
vKngZUtmq/PSF3WvmMgzUNS/BqOIMcs/B38vW3bkPOlRImZbY6A+ckb1hL7E
aXbwjTXc+snjPkBZDS6iRIWQXuQyjRQLVPXiJpYBrj3u5FDlG1XG1jktJmpT
xJPIfBBIsq7EqGGG/Q33ud5U0sB9OzXIYi4zqx0LiMGjMDiBctuB7hSugwTX
mhiCXL8oNToDZikPDUONSbhWSojixcAw0r9cfFfVraMUsoRJAKY2OztaEozB
KTLoZTlaWPjNhUNSJO6+oE/0Tm9ulDyM8xV6IqyzjZ4YJtpmI3uYmiQRHTqI
NtBs++r01zfpaB6w4Tf4mqIXpIbqx/VJB3uzhyPtmEDsD0IiB98Gqrh99WJG
ijbcD/ZwszU1s1r5pTtbiIsbxtWM/mkWoeRmnNB6tnEu3ozJfE5ILjf+NMtI
wco4TEIHHI+szqd5cgaFV/Gd2SpDOMc5s9F4OP/PeSuaeDQyT3YHW0EUfs3T
EqjAtFm74UbVC5eFGme3nG7saTS9b4pJ+DX+PLZdUOq9NkcmCeqKIFQlQEuh
771LctWZk/QDEJGjooQayABjilxdG1S1LUehY4ySAliUepOKHy0auyzXtSic
9xF1wZ0zH/6pwG7qypyAUh1mDt8DsAdkuqNgxHmneaq1Bmq4tZ2MbhDooOcv
qCkGV68vk8cxfZoknpU8JZVbADe5X+74gq22xaonw8eFO2mAfqFIOCtrHPHN
J9pW6CA9GcD9+N7gy0IgxWFFLK1PRfBRWY0KwN0x7iLKnzM9FLMtjFyUm9IJ
Rty13viCVWX0ldIx4SAxLcFVwLt6Fm/WPj4UBuk/LPBu4XIlqIErYsPxDMVS
bNJES8tE1wpPhotn09e0e54mm445vel6MV+U0s4D9Lo0p72z113162xUtVaV
X2dujT3AnQytVKpTKCUqgsbrpL90GWg0MxDyv4nzUwAF6dnsnmXK/cPBSwwe
psF2WYvpY3lULrdh7uAheZ4nvAvw5zCuEftaQjXSJ5vfwqjGQVaFWoAihwQB
tBi07kfKdQtTi0t2tqpBhFAiW5nO4UE8xirAC+g3W+OY2FNrlUcepDdmqZwg
7JTsYRc4+JnHdA3SfiS5AYZEaOiqyA+dhxpp/xS4AEtfVOFh9/iSpJ5xC9iO
ps/qGez0ES2uFZkFcHxBC4NG1cqi5GwLAr/Nz4bPWiUHiBZQjp29BKBb6pdO
6S1my2edzga4eoaLPwNKweTv+TkAl7T1B0ELsn+6CYAuOvdVvTd34ncwIhNi
GNhsr59luUiE3eJvfGSgmzGrqDV1qjLcN7j5sRWYo9ochSyQ2q4P1vfKWYQj
f9/5rcostTBtTqq0FFSmi9kAY7CzBpkN0DmzEmx3cASzpviWXVAZzF3ZgQNk
Cl0gTxIx6H+/Qk4zSIIB6xztB/74a7ixFxf4WeDC7bBHU00fFGkmR2zjCPrq
bRMQOgfoF77lNWG0gI8lWtvbshMetUx+n1+NpDcbuzuk/1ewJI3aHAnWBf8d
E4Kelp5+0DV1McAO0PW+Ow2TZ3pVKAl0Gg6+PbMabmYc4IemQpc3K2UIvydS
cyJtg2YDHvCpRcFPrS63/kYOujRGIa60EKZ+G52D7hdP9oIIGqUJp59rkUuB
BIZIUaNmYdZMyXCiZnF6M4S/40neHpFCApN380rlXWOw1U6nhsxDGpJVu8wr
B7Y7LHoxwbFALy7PEcxSyrGctveRqQeSC5Kx3pCV3AL5ltqnN8rNyMaw2ENa
VkZ0/fvOYDhLwMLsOJD7vVcnpcfah06vWEroUkpwzt4Yz1LXpY5Awf/aeufl
EcAck1ROkni3nxdRjvR6LeasOglJARgdtQ25TYqWcwrsmEID/9k+6+mtN1Nx
UsFxB9pFDem4Jz2TIo12uelwQOdtnXXnLWgtxkuGb69DH9D95qiUZOX76SBP
JmH4uC/V1CrkXuLnlaLF1u4p8zT/wM0AOOghKY59/UY82cKa/YGxFnPVk38z
lfQMmmScRk9ybjvMHw0HeEDKLebnSJp6XNU8oGcSSS7fetPiH0fXxDM/r+BO
AGMBUXOZJDLg1crOHFs8DBYGX4Ggb/f9P6EhJ+JVLtsp177y8J0YHYqLbYX6
nH8HjOCFd6fqe6J0oV21T2PWd6uR4NDcJzfZoKJcHswKb4+hsWyWFLwyQu8a
xxPE+ddYDzVc2Jh7UHfp0lTvsEDiP6UHxZxOfXUtYwAcbQq8rmwR1APW+SiW
28ju1zW+R2FQNGrtPAsnzWSWfwDJDZe5S9vrMNh8mcS6kNAqe7bQW1khaPrw
bi4vsBcv4/Sc3t3bAVLf3yPz7aZDDsoVwfvyUrdins7e19/SCRaHb0Mf1kM6
x3dfJqFoyxgOHTbk/KJ6T/1Lj3A+PKJy25atLlJGi+G426W0+baZ8u0tj0yB
6Iibx6T9RSrHoRVhEmH2sBX9Q/7B5PR8Ks/qGjnqLrlQXCkdG7A5j6Vh12ag
FKfy5kq4rMvMcvk1A5Bz7zB3UHaAUc+adkg76feFjCuBtV8r4YMXw1rPXbC5
qrdiHuNLmWrV8bBH1UeS5+J5s5Xbp1ca+wtc6qTrSDG20fBAjVEmDRS7dvDd
gksL5Hnv3R0EOWAn3XYofGfZP9nNXmeJN6W/RC3e7Zmj0uVhBPOY8/BSDd2Y
LZpDEg3MF3A6U/qnL6UwXCOLj35QM4FTEJHTScrKwG3sZm+pFMh8zmoOV/E1
GTffEuQGcDTTa5dTSPWVSJELxf7xnB7bb39WmonhCku28kB1pmJ138DXMnFO
h8kTQf4BZSNZa2UWnwbJYaRNXUk3/J0DT9k8pJkKXuGBvvjMqIKraSSvMsb5
wmTRFccxaVbHk7v1DByRt5U+T/cHBH76+Eo7L3qXLm623oPyI5mr3nE94SUB
cxqWCqJPbow2tl/1uz/HrKRFcNepMEBTbAzSzkaMrZxxLN6oEtDPI4gRR8zX
PoNSoyGGrpJWb+bDEk0mreevUfZq5CwEe+ZvfcY8xVFyB1oFyuH+BgGRUQXk
VcahqCO8LyHWHMbHL+AcBCT6Cu1Xtpmq4zXcpnl7F2UcZ3FFLxvoyeyF8tGK
87sxj/nraSQ9fqqgnlXV4Dif2A4hsH+sx6yj6m/TUPK1emDghxt/FumcUSQH
thW+NIHti1N7caN+2u1n6BKB+URL++OwUSyb8w9jzKiAaTS1QOdQhn8tjosI
QSRlIZJ0ShhmVDG0mHsD5SSMLEElSNPlleD9dNXyWEl7eJp77TCVHZrW2hP+
KLBMm4C6gubGsWh/QlmS3tvo7LGJf1K0egsuLVeWnOhPBshW+FsSyDrKnMpO
I70oA7ANq3WWEvinxAAcFG5b5G2UysdDQC0z3sFxvCPUzpuTpUfpUc6GUht1
GAn01OTAqvbLWlQGxwGc5YdUXBjTg7ClyjuT1OFFUvNwYSzzuOJKRiJkNuMR
ewHHCLuqBldJ08bBnVDhh+jK0Lxj4T8PPvK2KkhvGEF7jD2SrFWXpqoQTzpb
BY1CVfxN9SEmiMHxl0GonJQ7KfySJVx0FhwV5cpMwSOgwLYBXhXfWtBKHE+N
VKeP/42nAuSkqMdN+/VzlhruXgsp9mnMWUFJnW7OGibkEm7aGH523Ra0cZx4
TLg2n7BkGSP0tYMPcip2inUJZM3YtJoBbdk0+rKJCSDZMXGO6yhSddgBCP0c
uBo4ue6y1YbtDoNBFwt43q0gr25PSYSP1OvJRlXk73NcAJTriggMnQlGYMrE
j+6raacnBJjmWCLAk6JGj4yFgA84Sv6W0NZ8amEYUL9JBrcTG3aiBZQIUlGL
YO1SLs2eUxqUlOudO7D5VwyogCudGdBnlqYG0g6DISh/tDbLkIt8cTJZCV42
W8GYEanpoMLFunEgA5IKHIVDxWfcB72pwwOs19XKi/Vyns06lQnkMm5ap014
DlkWnzQ3Wh+/t2LxRNbq0uUcIvEP32eoNXO//3se77mp/eV9L6dcuFSr0lCl
CHlJi52vbt/xG+8uVdTN/uaXtUnDC/IqAce1FhG9409N1i9X4bhD22n2eBqT
RsBXaGNmkmPYDmZ6SUoKcgFeSzPldPTQEXRGG5fAbZhzuCwzsNKYpM7zEh7e
rUP5vBJPJzi7sOceox4Lr7Ygeg/biaKyV1q5mcXpMjzJkkKmNwEwrAADBiEY
/u8tTYa5H4m7ucVIMJv1rGX6D2UBWct51cdqXO5WymODt+SCBEW94HFRtpvY
+GckhDdLyV8b5HBwYeXlQlncao8Ahh/K3t/v4aEqJx7hs3CcNjfNOR3seTSa
6rO+sCaRR+MahMuSoc1DKZtKV0pFoZntaKhsyPj2AsckwIs/3TmcgWhQv+rz
ZJTZnKFoR91q9p1hiHu1srLRSqWtjouFqR0QbhYs18Fds6OOb2rqBnYETfJ7
hsVuoUg8aHm6Y47NC2miYboiq8BDIy9NK0kBfr54w4dEN6tia6q73lagbEKL
5d5tve9aTDJOFFabd22lXmckp9AivXdZsEus1qXt5mgQrKXPOClVT/SxHYhD
E2qKJjT3Kyg9sAdlIBW7FB2bqbWL9IgTyUBPqHKChCPPePWPRYNoZgStySGl
5YzuBKGOrRVhUpnlHfklEQ9FmhiZCfpF1eZ5/nb1hmyde+0PX4xPRAUTq1yK
cfaZqzxjxrkuQMiwks9YiIgnsBWfugWud1GdTQdehKtv0hHFAx5ovip9fSMi
X+ksWAg6tJe1CyNMz2WGE6vaIMC9gOmheAjJ4Z7qRRyQT/BtRG4tVGpno2cY
LeiLgmc8BEqwINZgkhom2gHfWt/+TE6qeE8PhhRa7ng0hOb7ckgC8Uzd4kit
SLBcCkUef8oT60MByfvItI9RAS/z/wzL/UaJV0+FWxWMFykMzXQLD2SaaRS3
9li9/MAjnAUaK52h/6Tb9lwhKH5hqTnLZKRy7rBYi34mpAcOITV3JICPTJGu
3maB6pKTaWk5//zk5FuiN2k8iW21ZERl5PKlqGSjg/ENIeQ5pXCuJQYRx0KS
RHou35K6UG5qbseuYePqRrzTi6fE0L1A4W5IfWT+dBPIrhUDMS1NNAmUx/lz
VnfLZaXXACbnj4DaX6J1UCrNNLuDTt8soVC6aqrMAAYmRaPE4H/wC9p5X6JY
CBHQrqF8PVsazCK4INoPNdjgh3x+7FTWa/BwAE75FVj571E5+Jw2hQeeLmSV
AXJ+cVRsCxWWSILQ6wAN/IDTx5q5A6csC4rj2FuKYzt6YFmhtoDHpDxdr2gt
TvYAfSoFp56oHnM/AD7eZ6vBN8yGBGg2PqnKK5DTV/C13EvrTs7SB0WD+pJy
tXuf5fGCw/aVzginOBMPfLD1X3jki5v3pJ8pBcIAgPqa/BRMgVfnHszTPOnb
fmPnSLZGad6a7njPCOKNjsTFFqGbs+H33e6dIGm2IjrlZPR3RzdxuCNI+9ZG
ZO2RR4D1X0hGG1SOqAgxam/ZQ0G70jdAVDsUWM1Td5qAqfanBZNoe8A5EGhd
COa3zyjDWH4ww9f4EzARq9BvR8uNSvH3L6bqY4RCmZH/xwXtL+x8KedZacJh
tiI=

`pragma protect end_protected
