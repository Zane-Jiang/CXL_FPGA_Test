// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pgqouYvzbcKPzYCxI0Xaagb+P7Kn9YEJLLKOxMOr6Q2mPSHFUF3pk5LcHGTN
cLiTZuehojgCHyYtV9YgDNSLIdrfTnWKksleEUjDGrle9gZDacnQKaNwZdKx
Wq1mwUjcbDCzgvWDZwFq7jhhlDo8vG1oJJw9pfX/yhw/GFfg/HAFlPxUaRbD
k4Jp9zwjVOpg0tsAuRojTzelEf99u5XxjMdQ3jxUKYsjJwMKSIUVj4E62jgm
oZjXbsatNg5v7IWMhLLacwlNQnXOEzZUnB5xaxR3SaYcE8E0pJgvozol6zrM
HZuxjIoIQu4sclbSNtAggySdv8fp2uvKid7IiostCg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nIcJOP3fSCtEUMsLsHmeLHDrXV6pMCorXcsXmK7RNLbUiJB2myKorHRwiLlX
WuIXhSGy2aCZ22hXGRSpf+rTX4j4CvD+oJYLS3IIDnvWiH0KgweZ9H1EvalN
KssOCdQGTGkvSi73x1ODiAAmqOWFitR1sKQZajXYH8ezUpGiiCbylOcYiVFY
uNui6lhkB8sw7bl0Du5carwA7lO40gd0mDytk11cssW71IqkD27YofoobX48
5qQAjkeXznyJYie/mT7s7FE6N6aCEpaG7HTy+6JxRuRL4ujTYxGqET1Iez2+
Dk1dBhYM8lkr3WoPFym2kUoHU2hZwrF8nbdyH6W4Rw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gWFgZeg5HrO9iZLi2rIcbjMYT84gO8qcgaqb6S5Di3pZwJJRRulWDFpWp5mA
AVIYUC3iFOXHAWgQw1mVy49s8IkCF0Oim0tl3srPJudG2XZbepzUtWLtCtku
cBieYQH1s9kjWpxx8wOJy7hofSelHEFRNYvt9oiXE3rJe2K/enADII2/MSBL
lPW9/KEYIk+/c+K+t/kwN9YamZw8JPPCPhtNbNpvjsAF1BkB5WFQzt2GUGl8
O+of4i8eAXSi9wjmPISpIYQXYTJedSb2HxEgHGMjqLpBor4WrY4QTwHpaCTc
CXu6g1At3mRJkRNeFhCTlIx6kl2XzHjog695nBTQ+A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IRsKks8x4JltntVlewx3Yn2REk1o4ioggige/PLDyQ9YnAgiZrk1wJr0DDh+
Q2/xCQTLwWwCb6En5xCKYpr+ZWhKreOLsYT8Zq8ksMWbb4aLahM0/Y9nmW9R
F9vAzP8lgpBGypdPGXZ+O/qkmQZC2lwiKm2JV9+kourUq40BJ18=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
TKVPAo1+kJ1qidXmRC9ZsuY1AzO/r+rlYLlu2r38y0VQZnAKLlhiaLbXC05x
zW8t9tJX/Qp6lzwzC9sCP5hRiTeMlrtdBw4Zz6oco+HVO+VUW2DMm1qDZcaC
Skw/kp06QCs+7aK+99CbdFEyz6pRhStU0Mu7n1AuE24pH2ZNHiCllB+8ofG8
liM3gLS7iFEthqdAH1Rlq245mQ7mqqg//A25boewZtZrjfYwiS0Qg1vABanP
08WTw5/STz8EO5fZIZKEO9eC4TtR2Tyo1f6QcDrVs/5LgC5+NPeO/acL7p9X
CKWGQJYPJg+K93K83bioHXgLrriUagKV7ndd4WouY3cRXiu/GWcJaErC0MLI
h5XN7gZbhOK4dm2VFn9s0cyIVe6A74TDcpamfOmaWQSVZWJzSizdsLUAeWVE
giSFCMejY9MRd0goLltxUBOLPaDkNuvOSsmDMYY38VmMbavKsc7kjKtjdTgw
CsBB2mUGDX9UIYeohBfwD9xcmOG3ixKI


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VwQQJQXfIuImbsAXIzcv6yqi03YAf08XQyYUJp3eW/f8OLzsDUZvFD6N6787
SWaEimJp/FxwdOT//IivqegQ4p7xibXGOfnT1lArw9fhqQZrx8zQ+V+GhYss
Zkk0adRRT3ce1DQ+h8CKCVsTbKYBVoJJG7CMwRa7yn/qgkr3gII=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k9KzNV6CahNynhwv038vn5L/8ZhvSbORrsPf4XbASp/HHniY/jJC/DRhiIRF
lJILNU8yx4TBhb5rp+1HUyMBOOVrme2Gvo1+67zyukqI0VnQBD2gP8yWrLlH
QaphwdKj+lQ1AgMLCHaVIKLKRdCqU3jaKyyyeri/OqMj5+uh8y0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9584)
`pragma protect data_block
jdmS7ImyVxv/Xa7KT+Jgpr+sbIghgjQGSq/EeX9G/XlAHfGpB8eDBJIbQzfc
OU8VOGK0wHFsCaOqwtbl9cF9V90tZWSTZYbX/khOSf2YP41IBXbQX9mnPCwf
WTWDU/++M2KzlezBhpip3W0/fmNEFyAnHc9SQY+1jF64ACr4gzcqhqCC2Nou
K51LCfQhemolszS9VlpGHTFL8PMMGhUrKlJYiDf7p50jSmTNCDZ6Q1iCUnoy
TUClSxxRlUEx8YqGFp/JCM4rxyLCMjFMAQC0moY2dSiZ0oHvjf0QxxkSv0zW
NdrOdc3nN0NYuNPv33Ln4GJGV1TN7V94/fV1lTheCiQ75MYWU4r+g5Sg1Rek
027Cczb0QXqW6LWlSh8gghg2bNJMoGPY0cyRiy/J0enypBcmVgTasrnvM4k0
MY5xiRa0rFPJtXWqNPuqombnepyOZtV+HMcZwQ5YLVEkzjAYt+qpYW28D+Si
++OaMy8QBNQdlc3lgwURIfC0R1XOrSd2ZGuihSB1Hjjyp0AOrl2E1d2Jksu7
D+WFSY3ZdN73rb60lVeTFiNcqCl3ijZi0UwaPDISJH3km8jYE6K/7/urhL7c
PfGr/XkraO9VZ4TFh0hWXax1SBxAxySg09a1Z1sAJjRsm/cCpFoyyCW0XTCO
wOw+0hPu9Yu315XDgMxrvguHGII+mlfhSd9jqK8icnhYnALMZrzmm5eUccpc
OZ62bMAFuE7J3CkEMc8QahG3EIyPVH8CCeqCMtQBEYHE/kZsOnNbxqUdE0Ui
cMRDYxdeK5JXzE+TgySZk4OjAZn/EJSY8Rotd2N4DpypZD/bVbpL5jI255qG
opbhXIuvx/jdEVaJ6rLavQ2J2q8OGqbX0nBgSi0jfD1Yki3T/fMyh2tkyo5A
VgW869dvl60ZrFH7Mg3GXuNB04aejQkDYSMnbflB5+MuVaZ6HL/ffKXBDHoJ
WaB5j10qOFH8meTlDRmozm12qNK6xGMnH5G3aFCT8uPjJnF6s9053XrmbN/s
wEoXXqA/Lp78t0by3SiV5V1ooa8F7N7Tfq7/Kr7aP9MqVcvsUnNE8KmhAjhG
dFaPnMrHZ1ETF6lF8Nznky1i73g7bIgA4Ip/o7W5pPKiPX7oqIzZrDB0VP3Y
aE59mxG4Jjo28xQBwrJM89dj8mwhnWO1NsSUAyQD9ezEiecBMBGxtXyi5XHi
5MIS4jVTEHhKT1a2WCSt/mCVy7mzClU3N7SpnHME0cxRGtVAJxUk5+bCBa/d
GGiAW0kwGKXJa+30X1tCF4vKw11sryxWraySDEc+zGdbT2lDz0/+0yAtEbUz
cEwqOD+r6o7SeC0pytCwBIbfYym/l4b1UXoV1WzXwaPKsd30gWywnx7HxlOd
DzSh8OV1y3uIHUw5C0pjFKJj4Ovh+OVtKWUouoWaOdPv2r7HUrf3JsAU6pXv
LotTjAGXF1RljlSX0UXMuSLDDd8Bp3Kczc1dhsC1nPn9MvnzezB/WxEiyKrE
9xYufFOdA6bat7HPfCr++SotNsCKyxDbr5Iz6qIViC3Bf6Fsq58+uxEgoigV
+vzJ/A/r4IOq7tZQZ1D67fW0mO5v00NLVk25kk/bTlYlwSSG8kOt0oQhQhjk
jnEt6PZitGtQxY2N35wCwu+8BWnbgvAigKHNxIj26jvlKqNpwSs0War+y5Ey
G7AO7TND1aKIw3ZxJA3V/jBZoVBhpLX8Ke2ZkrXOpd0Q2ViM1mkrgfx9T74r
4C/3xaQxU19olCO1TC/RJ1KOxXs1xg5dvJOTIZjsjstnaVDfi9nsz2Ukg2Lx
3MRQIVEnt76DvNGvodrYxWOKWmPEZZ0cGxsg93RKJytt0aT5GSSxDtcr83uV
TDjV2kRKgOM37QUk09eB/oJttCiengStFiqnqGr1xkFC3vVkLYCdtFtWY5J7
o/pSdlpAO/uCZAsceUrZ3M3NkdOF2Nv4+9gETlJTF7LikkmgKXLik5tlbdOc
U/3dV6jbmrn1vNTdC4zXY0oCspMwtAMZSWTmzHKSqelFWOzorSkIJ1zZysWD
KC1J9wngcdmfWwQ2tuELt7Gr0lcs02oF2XEi103tgPxkAp59UPVq5Hef1kak
EI92Gf/QToqVRys+8M57s7/21x7uJQXWG2QvfEybZ+GzOR2+0CGjxcuyXvIX
skKDWZKTcqTlbjatNJmZ60/Dzgg642rw8c7/e+lV1X+mX4dv+kqUsETm/SIp
1cxjsIcbQA4yP8YbNp2fmc7SvvmHfpLKOrh+2APbQ4DdmheuBovrqXTatWZi
3aduRvCM3QKko5xbssbuOhqwOtHjGAxz2nlv2d5lL5GyzgTP8SvNR67utvkS
CgQQfvZK6HPDVwN+0869tBGEiXd9Df6ceXpKoo4o/JLt1AFJMixLWNpVQw8+
r/qnFBwNbgEHN6P4H/G1/bLrjx9b+tJUDUfrckB70/bb0Sksk6ttbCiYfcVd
jj1CO+2ZIWGHB0JX+GTb2UC5oEmxxoJsI+w362yOosNPtxcLgLucYjoxNz+S
szs2rjm9RqQMQVVtVlJ623Sg3qdWXkIcBo8hRAeZVWqiYa1JyMRrlYUdVdgF
ngBlU+7yMZtyqpa97FsAkQlFF+xLWtuYSUAaclntAXLtmv2V3MrPcD10e2uD
no/1DaAkFAQYkA+Annk+5th0YHq8kwYuzJ19rsOenTECC2XJLDrkncjwkHOQ
c3en60wxc24sapNh02/3w0//biD27WyKOjDIa0MyCq+2iNlvLFJKsFRhl9W9
DWGdc+4rKWEMrstBrolBbmzGwKq3OYmF7JoGwwnVZUjNKLAhDcATggES+3y/
0b4rqoMthwJG+M1eEmd5pcgNg4pe1ZEd/eibeFvcykW1IGvMk/qoH/bjoMTP
mKFS7OvtFyqjieNcz/Xcv5l5Yv+JqAMJTLyaex1EUfBe04arT+L1XvVWVCpX
D5AyvjPLyghue/FKPPa9RHSr3fJYPNn6//hFdcGNAQkwCovZbh8CfHxswrw7
SBWgkJIdQFyI6y9mj6AGxX069ZXeluj736hZhZ5dAOq5swVdaNsfUDVzaMnn
arN+QeMNJCxSBvQ5R8mzfCw2lcZz8lmDiSX2/01ox7tIMqvV+zSpDKRGql3F
UymBr39hfZ/k6UTLXe2ASBcR/cuDepGxUZkEeJTK2nteGw4X4AwA+tDPfRLo
/jcCe+RtfPhMmzB5NNhROq5gMF8uc7wmMMOVXK1o2/PEXRsbAGgWH1nw0J5t
+Vz1hVNMvTXnMXRXgl+qzxw1cm1zQahKrF6ig2P0hPkFK2yvTVyaNedlnqdq
RVc8oVhOFARuBimSAe/QCDc2+cLK9wu2Q4gXYNCrPaxSQsDRb4VOxiBrVM+f
GpRrhvYnrRiRG3z3NWHgnVmZBIbA04fHogUCZXO/Ih02HfucpQR2+XXKFT4X
H31BhyxpuEl0McbzNIqKIQ6Ng6HbgGfYGbSFRr8mLTNJWDzXxDKL9gCP3pHv
k89I4u7cgqXI3ii3TVtmKexBWEYI9Or/MsIOQnzUV9YMlXY7WRY2X3Z61W52
3/eFiS4VMqXJYslelfp/syMNAMTbcWHT0thzBy4rkKerx//UuwAzvXr/Q2dc
8s/LrkCbkKMuh/O1kFsxCBbqXpKvqQyj5qXrKfAlepTMLiLFQrIAXvOLqfeu
SZfUTAlcmx3wrSn4Zg6XcQuoVCrDFpyYiXJdIymTfmTqsPfjO4suwikzBCEE
106XZlAjwIB46Pkt/w6EdGZYIqyNgPcdkjNO+83VZVlWunOxLMT1fSplOw/8
+CdpXWC7hEaNq9AJgEy9Hg7ivoxWxbLPHL4z6S+4wxZhx8t4hiXUciCOcvci
r9qqcFGrfAHnnp8m3Da1TT/R9/hRFaeYSyCy/zwZNdIV4xnFYu9K839exc3N
J+qKQ9LwKlqMOMg1aWuZNAJSkrQIWIsQwXySzc7/icCBerKc7nNCuxSSWXHL
aOimyqwRVRh8jg/KAz4KfEBmxbNP0inURr/qShb8jkC8QoDRaMjLlax8vgBw
9+kRqT++KVii7/fakUaLEcBEw5tAVfVwGHeRBwpECRJQxXMz5od3MzzhVYKT
DFEifbdsCsyhNbbjH30NFKS7xEixkJVYQTj/SUAmVZnl6BrwaBQgBJu68YXP
NAc1hIKl0Pl5u7cb90F0ZhjICE4N7Ce1sVZovDFjxsPByTseFPDUgr8yH6Wu
jPPWtwo06YUN0y7eEUyyl4339XHOkerFsID7KJF7frF0xRHEXcuBLIZVdmrw
oxMpGfnlrLkO1mgPNnQz6UbbrahF7i4GfSeMIyCtmoAjWX6cQNgFPHum8Tgv
2gQaswDWhM4wjjGlM6WrwFCNs9tYVmMSqkjioJMe9ng1EDDM4cMCgB6SN84s
t+nKmvpOzVnO9q0z4f/aB9/vlgjDgsvO2NlSMxHGZ+paUwXlusNsJCJlyrcQ
nGPknmJ/rF99vP8b0wkk02TsJGjWEEPBXMkjIW1tmmj+UyT3Xv1/tbIs4Mkc
8frbdeswMQ8Ui7kEd0zA2jYRpO2/H85acwwyk4764iiCK9m9Hv32WiYTlBW0
W3ukNLRpdKR/1Y8EV2XsaI5XW7lklA5cZgKjV1cPV25H+lp/EKeME8NjQ8n/
qfVa8PLL1QRKAroTTUZx+7d2Be43DMOgtTfZipUI5iU2mC9lg9wuKU1RN9qg
r+PGsNzLIFt4mEmsc1tXNizvU7iDj7VC48W1J41j7CFx+IYT2h1BHXJ1VZYG
5YQTGddjuMURfXrfongv4M/Y7wJtBj5hBxDd3nELrEvt2XoOOVm9L8fPbAHu
KmFY8Ug0WMrOIcLSzcecGGcNGacW3Q31gy6crtcTkaEUFicFyUWZBNO9Cr7B
Q4bJpyP8SWchHKuWE8sRj9PXzoUitPK7V2BFPZrpcEEgH3yLRJD4yB2gwPhI
DJWNpZWz7xaSBtwWK3JUDeZAQ8VDkiOwPg+K95/EGdsco5SbaehtUMVNQirO
SvG9nj+KKfFSAaapyjwerXgxmiKgS21gx/rs5O2Nj7Xt6738+aGdcpR3VwBE
jMcDUmw7UXOs/HaxCU18ksuSGyPNu2OmGVKilqAlqOO2D7lHCJ8OiDuDHMec
O0QixQBTnnyuLsZag/+sa6RZ6+NSqoXhExmKD/AhH5nVcDZzEzxrtKIzyfYj
LSIdwt8Grou3MssqnzGX2mXk6S0grf7Nc7Sgmw3lrQPxnlbotRGJbIySm8su
RkQ1jLoyR9ymc9kxArmAsHq142FIjPgpSdGmu1yCwfCESddcQpEeoLTShjEv
R53ipoS0+2JDXQeuOWJzmMPz5UO9zTs/3VFzWG/O+EZamsAC19wIS6KIDleU
UagH1cz13pL44jG8+1/pcFWgFuErPHRrCekaWhRP0U/L1933pjDwfNI1S6rZ
SyEErTftlYN99RuHubu/XWKnM4vsIAP6TltnJ4w3bBE89hRwnxc0mA4L6h68
r7h8hQ61rn8fcOfMBK73WqEgYiXjgPcR48fO+1H1Ms1xdaHOmAh721m0jhKF
pXA1GFkwltZyhtqHO8UooXDN6FeGemJcvhRg/ZpCXmsKXBAIxymsk+1D3Cu0
ZCfZ+PlGv4r0czuOhhDFcawNcuKTbEwHvD1u0HL97War83WkcGq9MgE1ZyK8
CUHezSYZi5VQhxWggPD6wOQ8uWERkPfUfkx4gm0/Lz2BlXwnJt8XGFXS8oc+
kxhVAcMoMAjsibs6Ut1guHnjF384sS2DsjdqsghZBryfzTXYeBMkTsXGPgXq
bq0aEqVCm07MFtX96UtgkHrCuaxjfoHM+NLkHPFhe9/oJWrkW/5xkgmI9T0V
mqmHGDCg5iWi8vTMTjMWoPjaMlNVuXXa5UbUgdm/08YDsqRG7xqJRpsP+43O
LzksrGqHHN0ffB0oVMJSz7eY/tq8Cnf6cg8nUToZ6hiq0RlmA6OTqwjJDiHZ
nZG2ooVYgJXIzciMzc3+6JV2uzULsqZdZFACMYoXm3H2TXb1CgMJZGxf+PxQ
vKBwCrnjTXBoUOp1oPCOajQ3bBEvpM/cll890lH7RLwJUIKmpQC6t7Mme3Nk
Qj72AG6kctyCAfz1ex5VUvD1qEJ9/zN+Jm4w4hBz9YCUxgT2qL9mkjNb36E0
ApLg0BFkfrNfqO6i3+lsVRwnjZH1usl/nJXjYXz3sb22YSPxcdXLWkcLxhVB
jHj0pkyQXteR18RsXSP6plR7jJPbMzJSjv+6j9Ra7PicMYboknTG07iOVqrE
hmt4M0536pnZapnk5ZK9OXzPipOajGa9BRqHUO1Fy+XbDbWqykkJw8zVEIqR
S8YbUygfeP3jrc0rw73YTtqMy+dPy6s0RWhQCchiT9s3D1T20eLu0KnyKTYu
l0XNr0syFQ/bC8U27DiaWebvvlq6w6PKIaL4cMaU9UTcEIHrmoCD2BJoruj9
tgo1nrGUv72ktIamy/9S+t7I01ujqiFZccToYJshW+wd6NVwv+U6a+uwdV/B
miMueLk5unea8ioePXu3Hr/r/dGX7AgVNZymHlIwyvZQW4lu1a1hJS7C0Ou2
PtEbo/Uy6IpMOe7EA1zeiCC4Fed7AgBVjL9rh/HMP696KMIr4P7ZLv8xq+JZ
4sY+XNgk4zFcSiVJrt9UlYUpfS4iqTdJGe0+hsp4yD1xVPdEnZN/7S+wSSn5
9O46g4bdbBXOFoV6tCKb++VQ+Hm6M7BqH6i8VEeUkM/xBZk5KoufFWzedweQ
QuHD4WrLWDTKGdE31cEwAl6Cefuu14nn+KgHRrEwfKALHqfzcfudnuMFM9fm
OtqmX9hkewjWB5DS4LCLNKB79biAfwZxyTS0Q+XBAnfABbOr6xJOY/1b1rlr
tNmIlGbtQ6I6kuPuXzPRa96krmGi1MNIiywIiFSXb+OgbYxlmSwO7H8b44p+
ENbhtXMO6DJd+Wxq3z2ckoFucfyN36Adjig/WmJwSvaerqc+xpO6q+otpCAs
kZmJ9T6MENKhdOyDUc3A0VpIn4g/IGzCKZsdMtiPK9m3GCDJ5uCd6knO5Jfr
2Qk18nhhyc5NoY8mGPY//KYgb55+h8Lw5SuSbFxFGPxGSG9Ku6FqnIjs9NN0
9gbuFd1XyYZuKlkBxHWrJr9XKShdMgFPTL+FtVAFMg05q+7rjgRnwEjQ6H/9
eq+/siU1K4pboX8I2J51+CwZJkxmKvggrbYp4WmHpbAd/PS+NQaZIFZ8wAvK
7eSdLAXcihAUHugi94dPpvO9dcSD7DGMJdHz7pNc90pCci14lWa5JUXjZKAG
awgnrHAxugVSHk5jBf0DMgApRWkGCDUvYJ0rYUY3Iszkqiw0nrwp/Te+MlCp
whRPQRywRuy8wcOi6X8qsTJTgBfjZ2JfY/yMz79/c4/5rcTRUrLVkPP9PBTi
74Y9olrCTvkduFuMn0+gXr+nKAocoTDG3JE7Bdop7ujet5a8wt8Sf1KVacin
klSGb9cmK44asby9em+SFm/G8umgKsDKxSAU0Me2ZnP4OOoaUUTk5ZqP3bXU
pjc1oOzrp878vFInvJ4xD/ZFUmV77XYPfkEhDRMkQzgoQbEtM+XcKQFicwd5
bJn3Fx6Iydm1Wk8MMBMrIwvRop+/S3wYoaXe45t7PAk3uJKFqZyd0Qw187Pf
+28zwPkoGrcOi4yFLbhRK5DzMHFcifwRzxi5enV4Oj4JsL75Y0LN9zOgxsg+
sV/exNGYcfdz16atxgQ1OP2DFfhpOLsRl+Vx3zutL6bLEMdgACEBv86e6xmo
QqGCGTWHzxd3bEcgWDnnxqA+XbasWSXkiIvbnntXEob//Ptbx1Uld9wvAHvK
HXKCpxtEd3yRtpLzUqqvdIko6+PuKeob2tV5uznQSEFDQCJGQ4xIUcTAargz
r76aqcYOB8CuKnRuV67KNZ06M0Yi6aptzbOeGdKP9AvHXN0WS1+gtKnxgp1V
Ev5ci75Qy75sQktyCdfjrNfGbq1gJLYw2YwDba3JhZn57/NUzpe9MuF+c/rp
wWotVHXlEckm3NRdKXYkFdMmylrpypsYxe1DwTZuqdC9NbWwvK4ORaTWn7ro
1IQVWdpJwsGc1nl/94KiYdZ4Vf2AhmkrUuRy9vXmFp36NoISsaD8CqGZXHUK
xoGJEeQ1mYukw2Kx0a88FYgzlIZgJgyIPQ+8D3dW5lxJKHv5wA/BWjZi781s
7naCmeN3Y8br2tlmxosset5IgiHi5bnrsenQ9csPUWnBer8FCnPGVIa1wWWh
4/KUXjM6qyLForFK/Bs75k6JSl412CVDWn4s5fUf76m2+sKI/Urm8h+AQWaW
TqHzG+NpL5/7pRlSjvAUsnrlH5jTVkmFsFK+cuN5H06YnovpjbpDXYAnZ5eS
D/rLfZorfTFK7qXuXRikJGvDn2JPaXaThzZgWS7iQLdPn5DbcrlNjPwYDXeY
iCBAlTfpv4ysBu0ThtcDwkthZiBCl6OABQt5ARhJLdw8OPqISssT0iB1jTjB
6qlzk5jsr8ybLG1fq35EfuDYk+mTj9OF2NZ2x0ArmVdqwIQq4oo9v2yVnVCN
egwN89cn/F22TKmGpsaZ/KDzr5WKvzHmwkcs2oDSORh3qq3rFYV5dgggn8+y
v29e5aX5pVsAS0oL4Q2u5GhxZ0lHU1d3kpsH7FITlsG6/ZAbrEF2o45feI0u
ooLhjqoTlgDthJTJaCJX8ll8LeaEcGUmayEgWcksJVpXFG2BBvcZfE20Zh8C
yLTl9GXMcGf/KRSas6c3b3sPypeT5OKjFa97Y4Ghh5qkbCN6c8bT425u5j1D
flwLGrpsLOq0ihGyHKJfrAg7qmImUgKZ8/eTtFvDhF3V8YT3xz4pQZXSbLGI
meMTnBTo0ulrngfEJLFZbRqvT+zV0etXQ/qS1Wb1juw0RZ+qIaBDumjwFdCJ
9nipTxQoVFJ0T6bu+a9tQpttkhs29BquekDcQ6z9+FF1MEuUbVq9gJJSC4JM
OUd01aMiLokL0qxqHvi/uQgLmukuyW0/w2EGXAQ+w9WzSmD33qhOhs1XXUa7
QH1hv5EsQXMZkSu64IinodqOXEVJfTC+hKZs/JGO59kjJyJGLxvO6t7uisDU
bjSJA+V2Rey7iUL38tkIpi99qxMb7zoDjBmNrAMg5fuhu9Bmtf9q3oZUeOA4
7yyOE117c5xVn2mKBfdGrrj66iF6CU2FlsTlNjfShcT3yLvV3bNTq8aF6nxt
VSo5fDpgQqsqL4oZTHaR4rSRAeX8e4ww1LzWmaSGDIJPTwO74ULdIQgc/u9L
LrAsD6jlEZ/vpwMy5ihENplJ1js0O4MYe3z7PJP2eDo1MbX8LMqaI8s72lqn
+jSfJBmKVDW1tvcw3WKfpB9IxkcMX9zH1Uv2NSX0uSQGGvZJv/hVnRRfbyUY
TkQ6PgZhCA6b7zUvA/OSEhDaI01mgzKY6beNVluxcLnmNRV7E9RmLXzjXu7a
v5xZTFqtr2HbWGIs4zyq70Ttzo+s5k3dvnM++6cu+eAtEBADwAP6SMxJ/ZX0
HhsMlCfi7EoMIxyBNfX0C954aH3dbILLvcQHuEGwRLQvbVNxbqnuj7MgZ4vT
N17sFvn4d3/4WKIA2NnNs0SQdj9jBUp7n4h66XloNu1diuQKr3e9cMVLk+Wv
xl5wVzYgD+ZYyqP46TJfyrOAcUun7mYsgbwcK/bzCY15oG4+jBEdKqe1v6To
XluIKhEmhX0JIPlQLupHTGnjpquuNRW2rjFMneZhAkbbS4ghx1uvBP3ibsxJ
Okq4hS6qQzG0GXCJGYKljlj3fQfHMqAYGa9tscMJZB9vwJ2TF7g1qkmTGkeq
oksAoMySwD7avHtmVLixshQQAJKP5b3SaRISUAVcfOrFDE2GiU74rikb0BAB
On3nVARChVdIWVM/5nYDmoLquk3vrwISBoc0n2u1jzbyZq1B7SCOX4i/XazJ
mwOeRz5u2us0YbdT9HJhbCK5s4B84W4nrn6Xk+Vc+Np11Hnyrh/FDfmGEjFO
3/X6ox56Oqh3nDiTTCeuFViJ2jrlGWJWyGr9n7S4hoTV9VniYcvMck4V2Ro1
6SKZY6tyIl+h+0dS3OUy/CDDzf7GZTpbbYXAVfWzfpPZ8WNcIpWjQE6DAl4A
YbjyaP9HTJt6S31zVuH0cZxmBsq1XPPtqheabeJ5cbf+mrtF3HgqyzzopHuC
Drt4wN50mCZrZJO3uoCKNDg9q0OCK2ern4iwfq/SVD0KWRtYf3YVWJvBI4W+
EH7trt8Y0hbGH7IPq+s/upVj8w7YOXYfQ4lm/hwZQyWa/QaBGAJ466UALmyM
UwXoL3FsECLpUHSQV+lkw6fdouL40HBkd/bKzNSnR0XglujwrIG6viuEkMD/
bkxPbaMEXWOnvtCkyFtauMW/f7PhjIF6/74p9+BdhIoPaT0j2GWXP1+E8KZs
X9ujKfFkavKmcd2BkaJXYYiLGUeOSuumgYNcS3XD9qGZJxwIX2eKPaxvCmsC
oGaRQJhBq5jRuVUpO4sYdZZUDRNrh5Uq54DQY17J1tGmCvz0+DbJ+eSFRQQH
CPJnNG311e1BLM+YXwb1rNSg1MsKohZQcB3vWxYAqpZoMEsOkEf5+jceYF/8
KSUvaUD36SclSjyI3fMHE85rivV/Q+djw7IztI8dfEKaXcB/49GvCTA+pYaV
z3buS1wujJF//HykqAyD4oMuBsvrrBvBXyCtuX4rCHs6p2O0rG7PxevxBMFO
0Grxnjr4Bemggg3FqtcD8Y7jvEkF5Ede6Y9FWrIoY7eWmI9U6N+TqhRSKF7i
08pEjYdd3zh8G2BqRxzEKG0pq/VCXtmatoEar5JyOb3uVvLA3eZRGNcAF8mr
CdZOS6DvqvnrsHpy9b2lygvyWa/UWAEotlCmv0ZaHUYUhrpHTz8mGo/H5Bdh
DPNmlqOGrA2k6xCJ5XQREKfLBCf2iKI5daxmkmKNGKzICGKfsFQfGtffYKGs
+4qO5zb6oM0Dp/DkRccniIWtyOdEi/zIHlSOHxuJuqhs4SWzM5Ma49p+daNX
PaQXNtfVjL5YEw6vc7lbQyegYFZt37tGLYV5CWzWT02QhgluzzMd6eE/MiK4
DqlxaWtl2WWHfV+0qKBqnnlfFd+vMbUUbfjA7Hksh5zVySk9jbfsNFiWBNeI
JwfmSI5SMHmgmU78s7UgC3IQ/XYOsjxaHtlWiOJk89G4PiswciueYnPJUl5i
+J8XcKvo9GUwa2lH9/Zswva6dhw8wn+J3hYkQnfFKlk4m0VxCncr1+QerAeZ
DpETpwr+zNr57OfUHfCNCBtaAyZmXtGIMClODuRfty++KrdmDxPu+AHGhcZO
RzkhZ2dGq7EmbkRyD49juVRG+c7ivGhsy6xxnPNxDda+7hBtq+gqgkZGv2G7
pkluahRTmN8BsIsBqT1bAved3fasrlqRnoXnJDxxBwFOVPm1Y2MgkQqfzZtJ
HzkNbB34Uu69fUVmQOl2+wZ6XObC7G15rJW04yspsy9kQnUoHz7TZoQ0IlBz
fNe0HuT5e7+A0C5E9zhbpOwgB7oCG5bAqgbzBkyN0LlwzHKjNOX42mCEjCZI
WknpE4cOqONmoKvYO2ecRpy6RVaFE49cpatTRoO0SGiYNfzSYWv/pGlB5x1e
jBSvbtLNJUPFVO1m0iBzPcv6pSwdHMiSchjMgILia4DSaGI6PKuzVjZvUbAw
wcxshYnk0OKQwJURMOVMF7/h12X1SracmD5OOZ6qVtPN5w2yXr4NKEqNaHas
KI8XbSFfvfXXQdVIIBv7T811chlqnWHN6Gbr5+NtQi/HCOChGV8Im9UkKVN2
SX2LJCBuYzIvMNnC352RtMaLD99fiuxCB7X+0DSSSPaZR4BIt9/PezWDO335
uErhxM3+CO5/BiPJTU91hOwNlkStR/ulQTSI9Fh9HIBb598cJsvbjSO65UTX
SXjQJTrD7EKBBaOWi5tRtBdE0QOaZiavO66LHEn/syP/tamlMAPqhXMDBCcf
zf/OFIKEBEkyhjBFZ0aKm2Jm3VZPRGXNPpPgAutNZxY/3IkPmIW1WfFVUYt9
4jFexy5cnd1z9UGx18W+UdtIFo/N6rgA70Z7Glo9roMt7zJesJgFEPUZciUk
j0X4A+waM2b/FRAP5snsiiHFxmWx8CVVT6mzCpN8St6TpsnXcNeUUHhaVKm4
0zK02PDckLUHjp3+iXEzMjrqtKO9ba/iGPTL3iQ4gDUzfYSpZw0GeOKPGqtE
5kAlH84tJ9i2luaShmVQfM8M/zbnAme0VrFn+AMWt6wNYC7Jg6EGqlrsaBs1
twwoueC/uJj365B8Cf0HBOVVvHNTZI14igD3co0Ycs2ywEaSymrDETpbqFgj
yetxri6jmf+WGKHb5bDQx/ZTkS65Lts3GE5zEz74qCwPh2SP68Xb0YzRPMB/
BXJy50DJa7udI3i9PRg0zbIlX4odNd3F6ZoR1jlRb8bgWL2RwfyLw+YMVgX7
vh8VJ01Y334WJ5o74WHO5Iq+aOlx1VlmbyTC9OJrZbJou3RhQ5ETuCWJi+D1
cquVY7Y/NScmzmWSIUjKVAGXWGj5UFmWej5BqebWtSzz/RsARNLUAkuMm3VZ
MhoY9hHPKSy6eUp0rJkODiKdLTwalYscV0cL3cl+qbYCIl+hLTcirCCtzjZG
/UuPeAmd3eTDJLE/GZBjHTXWeeXgqiDeX4tj95wjM/kssKgi88dDSFvLXOVh
q9PrOB4rTjRn+TCnXwO56rFKPXr+K7qbPwNjqfKEIe6HPbwnCCWrAUUMNpqu
vOWR/rf68M2mkUpFV/TUWSCoG4F1OtguumBKaV6IxnZwdjXrbw3WVoJBHLk=

`pragma protect end_protected
