// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
F6nsSLCVMvmb4uVOilPbfeHRxNopisnIAKK3B51ff4jZRhpj1fP7C3uH+RO6zQJP
d62L7Yc/vjr0ZaMaAEpTsMTCmfTNgYPhst4A12a7uIfCF9h43t62W886wWkC5AdD
AONqYdGKESceAZIAsvY3AX40tWElcdCWOGQcVFDyjfE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 46352 )
`pragma protect data_block
3UFLTkBcKwySb7iu8ibMl3dSP3W3Qik61mTM2hf5AcqbXsiprcSKl1tMq+2PJMjl
KOgVmOWuCqNaLXpPHH/31ysMU0GIMIaUVFIKBtwfUPGi9+eifXcVVUdl8eqH9skN
iLxSZyG4quqgZUQTU8gtJ2XOd9YiI7FqjymmeSSouiFFRjQLmiAYhBgejpZcuMUV
3nCN5MDjnpUSwHJ+Qbu4xn0st+fcEkghipK0InX4LfaRrAJRWk1fnxMcE/EYvqXP
Gappf8JmqqX7M+W8uKeW5Fseb2pPHjy/CjqG0V81A9tz42nmbDCwzZHwDZ9oArtc
axsmC2yFuI3cieP79HJjJc6ZpmisKdV2pN6+cq5W1geLrtN8MZ5QPeWkbbIgMywc
ntnmqdToGjF5UjkRNIJisRiUzi5ux6c+XFDv2DoO6+gLwrZEvcDqs6Lu7vGJhj5/
oU2ZrA2Z67kXSrNp/YLA4FcoiF+2YuvS8NExKlajHoah/QuXQ866SRTuSw4uvj8p
Xlu5LyJYtvNb9YSJhzzReEH8S0/n5WS53YpZjupGCIvwOeYtvs/kkR7nlsag+QVh
I1lVGqd5MkP+fU/yn6460AHHaS4tLjFMMXOxg7dmFZyobbQgOmH8wNcNVIfIiSUx
3UCisBInwLQTnY6vmS60vNgXZry9FlWrTwfsXlsKMGKRa50hvpZTxh79EDBcORiO
WSodI+oEYR3LGzExMVLM3CGhvFQCOj6zlqPGwq6LKLfAtwkaRCkWWnu5uJJguGko
+ea5EW61EgwGxRr82UbwS57YWW2NGneBcbu0viquDUD6trTRI4fPWLCsno2/i3oy
lOBgMX5gusYqbc9/bwcTIW2T6x1+zyJOTEFkdIbMCm7WYqKpe4hQZfnDZZYjFRge
SP1hc9ewfnLqV+tUjzhAixz7unVY8oliv0xcL0L5Ud2LLjL931Q16imp4HnbWbKb
K+BPqwWfXj8RHz6B1dBqc9UG59aLfiW7GrkHvBBoyQrzXKP09vrAphoLIYX7TONr
ryjSBAshEO9V3f7O+1jm+N3BQT+6CCOqwA3LQeUX78i/GNQClDkDGe602/dOV2+P
V6gnocuG80GsBsqa2P+5Nkb4nz7nUldAw891p852lmM2r9SU/i2m3PAfoAUgF3wU
YspZ5bckjEyXG6BbqjGWkqq81FJDMNbcj6Hq2sBPObzWzYY/TSiF4ZinB1JWN/UM
x58HjjlThGhTG3Hl8Mh/Uyast5e/QY3cDEHNEe4ua7p89cqFOGK0ozhh0gGCdjDb
vJTlZsFXQf1AKeNPExZQ7BWeGYPdYHegcNwo2UPtKOuFimwBCAhYh5Fb6BnBEcOq
B8SW2k5tmHAG7zzkbxNkp1E7vp6rWDlz9MNpFSXljA9A2QIJYftpaW0mIrNgm4Yt
LGYamFpc2EEQGU88fzsIQpY6aRN9WeSUZkZVZ6BJ3ZuvxNxhuNnCoBURqzaQ6GUk
MnaVn96scGRXEGUFxW1EmEoo4OAsigJbnLmjonjVwvkYnyLGjUXAiVdNHNF5kjI3
VIpYzKfDHE0lGZu9/QIo/Dv0sKk81L/rWYvgwg/5sXMvLkc+GJ2xLFB+Fz33Fk0D
L03IVbRXfbpl0+jy68OuqQaVV7dJn6Twuk2AQT3Q3iylSUvlBf6CG/mJdVBsWwcy
BVu9oZ/34vY7MtLTrLoqkYyUR5DmWnYXHN+46+9vejVnrJTc8YRGYrnMszqKhBth
tnE+HHSOdDW5ySRduJYE1wr3bkUiFXfv3u4FuZ3/CeB0C366t+6uV+bIyRpHPkm3
8HBNGolQmUxBwHkuTJsYjXOR/246/bUASheC0MzAaPSO28AdnHt4225R/ug1lb+G
bvZu1TKGapKUnxsOV6i8UzF/6H0npSW488yAAsYSbrUXwBPa7iDK1P1QDeOxCbq7
EUvB5ZUDuEDOIrU7g8mhq5KNezI3JWmxk+V6lrFxojvd/AulQQonTPcnGimvtkNM
RVOpxZxO0ZOKDKrmYE58GnmKyYc7yYufPwUPQz6FNg1ZDpg8w+QSksbHwzkpy70J
wNrUosfZv9KHkImZwLlSphejhoL22/n0CwcYWPP9pATR1jDdLmPDKLD1s82FNEvG
hWk8nPEnuu5iCLmPp55ZkNi4r/Bb9D5CzKGcMHZq7a1LGHpSaXlgPia7dyzZm2ex
5GNv5BrJKEAfxP8g7GGtZo8J5VXaiFbEbu5EsKrME75digoJMdt7Po86YF0j65mz
ea+lJEHfIenCoXyuwoXIs1AgjcEd/Irh3mqsm6FaFzJgvCYmxpME0TCOS7+QVtJr
n4lYILD2c7rZ8fBOMm9jXD62Ptxtwj1ZLhorCA06Q2Q9Ocfzim2RFlMoDDGRcB2f
UMw8IBclFqMoKxmYQSJkOkSP8WP7+m4UMDftHL/ztDe7ATK6p+ApDn+j9oPENz0H
v9nGDvvjKFpaYxwk6GSFQBOG9VG6y1qIN50AfKEE3ipx1pnCx9nqGEgopoRXcB1C
+2AuQ+QcT5CGkxa9t2f0wu1OsUc0a7C5Qflb8H5ImJz7IxQ7gKXbJUARnB2gXWog
m3xZS0vw0cMAMOk1IrtBhSL79lvwkBhHUgP+NRW31/araDJUK1hObfhpmWr/ic6j
AkHX5JhcSUOdOllnc1pTb9X0Bkv4/tILbzyrQDOgZ0RkEXgA6DbDzjpP13xnrvge
/tmZf+dT2eVVKa6WmzQXwufCgRna+CRxijnUjmXSUGy1uOh1UM0MuZR/snzCQ/lm
Zi969iUZs+bdDaDVIxiyB6lxJdlomRYgCN+nicNkgEuCFDk9qiATEoOzmwBrpp+L
/k1xoCrLCDjwf9lyoA4RGQdYoKPujCpCmabyWZnvm46RLn2xMgBKVtDvDkhL1GuT
cnNXKaz2xbdREFhjC2LsGemmSCb+cKYGs/l8ktHG4iP/Ktd9xwm2PsZwt0J5mE4Y
Ao8xfDPdOnQJuwG5X/1P/+J50dmUHshIYLLHAzs0g/HGdATiZp97EPA4Sr1usfMr
u22pUk9nuHMYK9Z4kXDfGTeETnAiMzdjgc/L4X+VBiz9j8Lz2L5SMoukgjrUM84Y
5pfRUDrE/A0ASpZY/v8zMQMgnGe3uD6bNviWP4af+xzmm6RjjA7MXzAUV3fx9xqH
uSjBJoShRT0a/QNMRD92XoaUPnkekuBMFiaO0gATznvhrcMDwsMg4LODLkA9Grgu
JQ0Wziiq2QZXsqftUOrq2bVJYRTiHiixTpKOhViO5NkJ2C6qQ+eR9ACvtpK0gSMV
J7WSHPai+36efx8VrNJ7V72jc+aY9gMsa+emMViZ0RAQ2v1KiVJdiwtasroT+l/O
LiA+qo+KVEdTbfMg8GzSGYCwAsfH4GVRw6VGz3koKY68z5LhjpscZYJxK9kNoQRI
g6Y/ZU3KR2XQxkyOIoxmBwEn2Idcir4OpaqVLKFzcVdbNrJGvMZwXgWTCngbf8t4
vUHvJTKzUhNQIQdTE2tYX6Mu+MULF9twFdg5wzR6muGmE/p5xMNw1C3/VzrXqO5h
nhjw+r+rboi2QURIYFPizLW4EPp4tnfYk7hMRE969BsaFO2EPNrjHzG+TzN6M2R0
P/b+N6wq/ToRfTd6Z8FoFMUB8tt/qij/4l3Z4wMXMr31u9Vc+3BPrBlnzvsrbiXm
mLRFySBWGJs64r9H1GiT2P2pOoEmjr8j6+7q+QlnUm4ScjnuSu8X9X+EFpNbYbq1
zBAvQ1qEx6ipsUsj9PFQ158rlYheZXdMc5lyxEDgw7JaybYv6GAS4mKbICDmQhhC
E9ZgCr04KngBBPHhWxHH+qFnrh5NPAaEKKCtBI96Ep4CZOG+2EWIF9NSV+5dq/TH
PYT7g34vhY3K+XA8/ynE9hsOzbrhaYlgSWQV539EA0ZKaxeqUB16ytbXsr8JUoFR
a8ItdAP3ONRW/OtDsIoANSkzU1R6p3yciM1B7QeuPjBENseuJCaHfviMh+bcxLAM
0XNvP03J8OuZqu8F9TYNdfbJNpHeghQONrrqQ96MdiyZT1FJZJ5uX9chgOIEK8gv
bY1YGe2mdCKuHxztPtXZnjhHsAyRmO2GvIANv8/hRxC6TH90qU6m2cBN8SEHWNc/
GGgmvc5Qsqod2E5sPMyaoVSUjoeKcEqv74z0GX6N9AVOfr6dNlTLcso+R8WDbbjd
7U4vwXucPypTU38G5198Bn9etq1ZDdJEjDPVEtG43haDCV3jQdkXg59uiKwOp0Wb
d5HAcIV39JigRgeiBaWQ71BeUSeI2MOAwojuh6++Qqa83xxQbqetdjxce0v/8351
j5DkKo0f2iH04UcHNdNeVTAagHBrG+bj4ikQz3rsLcBehc1MPm/eyESG4rzQ+esi
hBwUd5jeIZQtB1k/wAoJ472KsTqq3f6gg2uhoHTz7qOwxApO1v1p8V4nBLXw9kGo
QPIgGSHLWkAeq+9XEz+oSsBV1Cw7sXLbceW+6oQNTyGozVX+wc9N0rrAUXL7cV4s
UfVpzVZcQjcDbHU/6LDxIU3ZR0y8cL9XURbBzEuNs+1Ngi09nXhjxBjzNRzyvQmh
GCn4R3LuI5cY3DD/vWnRhG1wkxj9lwaIiluh2e8ACnE0JBeMXRI0gKxsOPdJyhDv
t61wLem8z39r80gEz0dZ1yINUlSQoUrPq3pV56u0rxL9aY69XAwAgW3HS8oi5qxp
qeMVRSU6qGzpPo5SWunjc8V6r4an2BA5MPKOvYLswjfCUabjpYQs4n6J+U6pTTED
IviGzCls5Rv0XV0/xiRKxiTEXpaIcN6XY1pR8htySODAwM+dotYfu0AqdoJ+01Np
HD359O13ABRAIYccqAqvUGZWp8JiyyjDRbWvcImeFb1NHdmgFa+d88yCKthzSITs
i5l5rN16k9ch7CJYDuAxOsbkmyqxqX7v3/vOFhFwkI4AAlG3avZJU65eEqywq5Eb
q6SRxHLqRq6I5X8UUNWs2R2QxK7CWkLCbYsQE+yTbCUAjAObtgtkakVzIj8X/ZCa
fD7jIL507YpHjWll2vBUg5/zv46NQvHaPuvMDwHST/B8vU+gWweuFsXLxO7Ijjks
fCdFKAdtZrZAK1800GXgeXWLXrSlNRwTlK3QXg7iWb+AC/u3NY7H0tzyoNRbXnT2
fH0HFke0JqxOAT5eVEibJI7ApzbWPl3qXKrCTFHH4WcT2hPuLo/V4Fp8re8svTPA
iTLnwapPjI055D7F/+n8vXP1nAD0wovjOT1nK5Ujm1Or+H/m5edLUM74b5vuvrwj
qiwqzMSp+QzXrkeGAwdNFDYFCrw3vv0yqExVm2uYZkdnlYkjZvDhRZmWcORtGSEX
hUsELsxm9ApWrdhuVKJaOlA4KfSIQzj2iWNYamQEN80xpeIdf6bbgocAMoCwwOlI
XFsn5AitsD/pILovmrUN6MUfGAsw2lVmwjE85pinGAamrUHAuiBJkrdTBy0nqnX5
UkcmolnQ7CQ3nmjQGaSYVP5SngorwW9bC+A/7qaYcrjG/XR2VvPbjwxQhD6+iykM
rMUqHn34+jhJdBaD2opMAobe2XPW7AVkdEE7EOV0f/pIpJkke3EWDBdtfS/SMUEV
Hj4goCLS2AK8/sIji4V8ejTpuBixZHLFl4xVkpc+gPXsCEFexYF50hoiKzpO170z
x3AIejWy1VSLpNDAi7cMqqwHEMpsFWwsxlXw3MxPwjnSS6okOYumQlUJwmieLYQh
qtD0+UTzv75yIqWPly0qqteoQGTKct8gYl0B5vMEdH9YtV4CfH7aebLU9sxkSFut
spiW8IYe6yO+WkjON6L2YGhVVoJX7yyOMiyNddZkPdEfYHYiWk/y71wlHo8S2ssf
AmNTy4HFqG78fzPZeVpHSJ/qS1Jb8vowXLHi/0mNQj7g4GZpPxTjMzGYytFw/Sxf
krnIoHJP/OINPPNC5L3T1id4tadssHbhfu/Jzb2mcCgfCqt+ZeZ1wZLVmEy3Mw+c
Ikw2akhhAI5RkLSkJ1695p7WhbopkWAjYOvrXiNF4BH1RqTIl6bNcEW55cKG1zHt
41rxEb8db1LZfxo79OvRj2vuGcKjNUZAz3bvhBJSl8NId2fV1XJ3cmzKWmN60iJi
agNiOtfcRQrPaxSrVmTDih0J2BKlFFuGZB7r9PoxBe8p5896Id6an6BRZ2io0eYM
W/hr5LyYs4bRSpziVGtaWdpxIoJP7k7fl2XqtsrzUd9UhTJ86Boqtz1mh8M7KGN8
pH5Sy4Y9qfoX3AwLiC6ShWUdEH5SH3QBsluJtYYdmxyHAd1B3+qsFy4NGEKijSu2
cxqHV+t9oE5MbK4l8eEAOLcVY+VZI8e+DGcMJ/btg+QwF1bd6FS5hlVz4P/LVQDc
R7NeuwGx1PmgZxm7joKx1p3xuEDBglBdXDoVvIkndN3+0iuXGh2mogaKK80bXEqB
ut/RASCfOy4eKqwmwP2TS2lBKykH5IIpBsMW6r03oPRWmZQWswgclw1CSYQJ9sU9
f8LhuOWpTMJn4lU+rK4zODUaG5EbPX/zk2Xs2t3ZARkx/+2Av4Hv36q0I46fExT6
whPNbCNZKSVg2hzzVdwW56KLLRh8NwJ0yFxAdA75kwtgTdsop5IBo3MIOvHiUPVF
qnAoRZvLjmzo3ecYEFmobLr7osviPXVyZiYWXwE4BIduwQ2f7G2AU2+973dbmWAo
qZpfV5nsbcBi+4qoFjOHpWzMHfLXmoIG919L9+JxVEtJvySMDtM2tBFlh82i3hYE
4hCXJrFt3Bgq/nA6pxj6Z3Mc8k7h0vhUoy8jxoF1x3oQio6V0Gr8kn8gian0DqiD
AguqXiObKuomZn008/UHqK1rj0e0JNAgq101Ieruf0fUKJ+SQ/Lmo0jQMZiLqaK7
HT8gpXwrCGMLzG17yN1YOjogRtJ7nzJqGKG9P2FZllbVUFFyKqvEvq5NHnjsynEL
ftocbh+h9mg16OAXjeGfrNJxy7iiBEcH80hYiseUy5lTcONUmFr1NGp81i+FcYsh
Lb+lJtEvMU3VZGo6o7Hk8GkF0NfoPLQCOzfR4IcdoKY9HK6t3QF24pU9LmhfqZ/v
EsCZ9BRXWin0N5M7qYUP4wFM3qoeo89q8QSxhesFANwfO8NfcsrbXJFji/wBRfUX
ifXc4Hw0IKyDY1vZNCrFgD9GAbFckgNeLd31kYD3SpcYecButfSDO/4vH3jPaB4s
VjIXgd6q4qUrQCrFARmN8QMsdfGFSNFfO676fiezF4HQBjHMiV41VN7vJBtrn2d1
yuHsIdyMXV5TBuzOyOVz6wrDpC2ix3qU+KOukpFyC5+c1sYJB1/BM0l+C1ypKqrp
qJRF7hKrHkBQpg6cgyOJvgLr00gRGhw2DoySmIKbiIrXzGR8r90WlE7iLOKYXKDo
d/ypg/VGizllT7dO5kQu1I/bVvmZBEd4DS/irJYqdnFBmN4pPia3eT9FSbvt/bMn
91KBA3WgwwL3BhF0YHVHNggSR+ZurohDQv6oMjEd11XB7GdvQ+9zt3x9c3fogiwI
E8oJ3K5o4Ch0jXHueLNt3iZl+C+A8xzAiVj5sZrm3e76SOr4BZ5ebDg9JBuSAypm
R2eNndTbL0uCPP9QXhHx/xHv5zfv1Hzl2NGO3ikqA0TY4h53veE75M42YfiDjLtI
gLNplEMMiTnpu58DmGd/Sr7wfwvKI+iqEkRLXV3ASklBORhhkQstHgKlNryPN4yq
dijnq7+DhxQa8V6QnDnMDNs+ZfgoNFt4pH7MZYJowctYFVBqIa617yzD0UqwaS8/
A2WHwer0qKUvc8ZvJZKcFqnOFYtPfu4gtfUjmgzeCYThUXlZnGv5LNOmQoEGieP/
G1Pa0M61A16QbIRfc0sBlehG/0wTA0sEHMdCMarN8KYeqK7TKs1A/hHAxnYhfN2l
PN7vBxX1tiMIMJK8XyMfA5NEBnzFi5Ch6TJYGDGvFH8m/Vp426zCxWAvcYORv24G
251u0GavmebZ8sAnbl0naA86+Ot3yiuW2eU/oD5yia2n1S5OLHk3KXmYIcGNw8xz
oqOWSrQrorDf1sEs52+W/WsBaxslxSsCP15lMe27T9thAuxfan9N7J/xqFPhDVtL
I+9CkTkQzB7DUd3cpa55rLq0zj7RdizHoGHANl9mM47G0TanWTZX0hk41T3FX3F8
uo/MtRwY26sV8w4BT3KI6fxmo4ym6LXIYxpcd0qyz2UiJC3U3EkDM5FJCbihaub5
yUn+a6PtoH/Dj2MfJLwuUfqb6ivBYs0JbbJSmv8Gv//oknHpGi9Naw80H5KJm3qD
brS57EnMe+v391whTt7FbR1s+O+Uftpx/tK/TXvKKMNLPkR0QRRJZF0urXCeDFP/
DTi52+j5DhfvtLls5oSVAKyMmg8D+o5rDU94oz+xPeIgeaoDBiYuYnq5ROVLsiaH
j1OYMMLMt3JMW/06GkQjLWYL31cXClMC2TLh8Mma1hoaeI1DmGu/rIu2Zul4zhH0
7LaIXEFHj7hx3gnOweqc3BKsi8G4t2S6mZpX77K2JB0J7oRDY9R7PsvdNMC0MaLa
XvRiGHctrn5x61jPCppHmRR79uynTPUYsC6+iJXd2D2u5syGUBVzWj2LNT3M+mzk
MZT2Pw8Uen2QvtrIEcRnLHw4jVexjA6+c6p7KtHyBQiXBHdHfg/N942CUNtfm0hq
I1cUmtoB6k1H8IWDWU0Sjn5t00tuaBbKJt1qaU+DT2yyEq9zGi4GpuEw4pl62jsN
Fk0cFzdShdy62FUENDbV6lK78Y23f55C4RoNcKjcmOAlMZIElgI/IVVHzhSm+go7
2WXKzdy5ks8Q5GutNrVfMp6Za+EulqCVUNavZUhADee5J02KAtRN3BTo57xBvwFt
DaVqmBqcVdrLqdz9Zwv/zEkzUMhppSCEtc1oc548heJlpQR0iX5+mEGouzeRsafX
mgTjEsms/bzYoJVtrIV2lMTAnj/Gg7pv4wsjSPWKWdv9JBS2WsqmVbW69BNHTu6u
yeWn1VnZP2QYdUrgehlu0nX12tqvJMk6m0Qz/WoAXs74DMuvU8RD2uYdKEVJXIhB
TV8i6alC3FW0IyKNRsCBbZQjRmYBaUoJzQGJQXs72ttqCgvsP3VY+9loHHY3ozM+
DAMiWsB7UJLbe9RbPXM/iLCjGylwk0ftyKt4vajaxikPwkUe9uvA39xbMEMZL7KF
6zR9GqUGGcnj2pheIo0PYxHmUOKKp36YdQIrqw1hGk/6GNSkM/XRCSrQhySfBJXw
whOBc8tRGe1kslzWYEFDNQaKgV47/mV961q8+yOgITwRyws76hxCxiKXfuiGeHF3
sBnUhDB8ALKYcCCBPSPHFfVGHHLOpLbA4EsSWn65UB+UcG63WGajjruarSCrr4qj
FBxYDjTbPV3pRe8idRrBHdx7jnJjuVlplf34hNgTTgXLKlO4vS17KfCQoiSEv2g0
1Fc+kA/sPPNk4WHrn4fJL/ewLoq2ESa27KKQv0puzBXYP9UBPOj0KDqy4gdJdMsw
xfhnDItx8B9wvX9L6uzxYBqKjAfVYtZxQ0jM7JJORYiDawrkU8qogAbGkZXBz/Vf
7ENer96gMcqC2V9hti1XIzpeZKG2rra2I6f4bDl81Ctr9gvE7lkxtZ/Coo/9aKT9
ltChBQqAYiDjGJNqy2zJQgJDQslhwrDRNwIZD5MpKPZiJhze5+R2LGfc1tXOD+A+
UdNeXkRankxFS0RPjCGYtIjBDzR27H6F9d2w7MzQc2ikm6LGT+1cctH0kjTYtgVM
UExCbPBcyRFGyj3iI1S9lSlwpUewqOtsVXIaHj3aIe3A/WO23ro8a2QkkButcSJB
gzONUxORMvLVvC5Ihf3OzYq5N2S1VXRVrbOU5hWWGlvINPd+tua+byEqlnN2xUSU
0ZuYQRKMVBoO3/T3qtjLh09a7lNcbfA0Du9L4G8UuyZEwiuv0SWCO0FxnotDS/af
Amgx+ObcarXpCVKhM+Kvtr4z56VQQ1hlk1hNJ2OhbLzm32nLV5U7S1OyFe7F3NNn
8FIUdBOh+FzqMEL/oydmWUqnMkATOH1rcyh6ixXPL5xXchUa0WCxRplrjXuqkkHo
g4Rufrr/xrp1siK3BU29C4uKeSb/eWXnl+jhmnaP1PCvmR7gww1Cps7Ll84jWjsT
pmawdya9rg35DD3Y/yZTiyxjIzYYZDwqyaDyOZPH5PD5kl8eJjvfCgU6nIYxo8Mu
jxksbundaoztRIbFRc9AhefgcJr7SKYPsbFtndRjctu9iNyerSsZt1Zc31S+CCAc
Rq3heEftzgYNdApBeLCVtkN0LePFiUEWlTqPCQ73N84s4VTEAT6E2lKYMARI0Fbr
GDqCyo3kEKQ+Qk/HZsXaCUwBN2QGzlYlHftcZQ6tn2Tl+98KP7CXeNsw2BsAnv28
qWa9UFk4J9WeZfMiweCDRyV6XHoyFePqpyLSqWVzvTSoUZsxE0U83VrZAB3ShcZ2
Aujv8/s4uRcy4qOEOmPhZVBZ/KqBbudR79J2SH8kX01eYjJXK4W+VBTsL0ls2vir
cQYEmLHzw9y3Q9FltbTM3b0+pj5HGTzHd6jUnKVUQ+d1gALI3Ausi1G9vt+YCETd
3nN0ZQE6PHoR2fASD0QIIiijZIA2iAJIEjrjShlUNVhDxbgX1aydP217My1N+hav
EcTo6LgPGCwmUtNPpWYE/jDE7N/CdOLNtxVxZG8fx70A8MIyqJee4K7E9flwXhj8
1iqjGjYbVpGrmWIuvcAF+KhOddchJuYuuhDxURHEVfHk+oLP8P4B/N6ILy2v0+WD
kFa59ixqqVXyFnMLdeuzWblnKqT5o9rozcIZ0wTeFZ2VqC14Sya7eK5je7ADBeh/
jVrwhwLFw0C7EXDWi3VcwqXN/FP6FOIxW/vfYnYX1IYH6oPRpWwIlC8zODRlJXBi
+MiZsWHvPZBX6zNmgbdsiXaF5I/LVFQ9AppmtIFlqDbkp+nM0SVzer//IelY6Zhh
M6An8RCT7g2vfK8er0H8EAuBl45g4dLZcii0QlbJrQT17vSv6AOIzOrap9dLgJ25
BThZsqZafS+qqKi1+J2ZF2TxU3Bq7BjRHWFNEBkFCcujlTK540HcvMyWPdEfusOP
iYrA9Hb7+plWO0lFx14A71ZG6zaZbGnCEFnGq283JnbbBdR3cbIP509mzWUHxi4+
AcVu2UVu1xwaSsV8B90/YXNCYYuJyX545g8wVFToDMgmntYtInkhP5TkZXPc+CAH
hVBDuMhhIj01DzUXq8Gwgm7DCOGueWklhX6v04/NTt97o774orOOgVFY2RCf5sq/
6UId8cTfrb3l+Puuq3vHeRYoi8UGbkFVYpBe38klqBX6nJkCpAGIkPpDvzcNPMzi
XC1wO2WlTgTvaRkt7DOPVx4SbmPkwf5IaXe7rMgxqFKcNFeRjXHdb6R4AwFhNajk
awGh6+KMwt1eWQJtWRo5Tr0s9Ac+pMfQyfpChFxBvtcOzjfb5nOwxUZ+amhQexmi
TZMgPCHgUKfeNPyx3XGMO6pSxgDACJ7TqVjGNqDuknGL+IZPNKBehBaXfJzEFQUc
H1smQb9G6TCCO1Zn9gbukT/NAC3v0lozWIt6MDfO1fRCwqEoQ4PU2oczjCG0tdD3
Jz/Rlftb0lLKxXvU1zP5oKlTuj7le3Evxs1ig62qO21K8l59HSiteJ0m1hro6FTl
2bmiXjLcrzaomBQl5fRoM6OJj941j69NMx6aeihK8trR2Vsf0Oy+0PC8dchsG7mr
w3ngeSRj+qkrAIQS8q2xg9YkVc2LyI30UH2AfMMM3id5o5X0MVy8se7W7RlqSCu6
dhM+Mvwmyi9iIzkWGx+nePip7fdynEeJ7VLB9PlE1tSI0EylTSM0oP/ipOvTXd1P
BQmfYtqWIV2nGT4WCgxgKRmkJOtJXhA0JPN/piw6aA0mAMjUzjF2Z49UmyrKC/ke
udcgF2NC8yX9cNPuwFqJpe4DqVh6KO5o3SBwboLvJJ5kOBDwl8u+4ynKUykXvxV7
LVNeC9i7NaKSEbpgWJ65BXA2/hqsVB31IaOwqUEOArCybJNFD8DwZ1claR4Hzx2c
2w/LMujpR7k/lyusKUAeViKeLHmgQqn9qSdMFhHUg6n63YShQRA0oAV4QhT7+bm8
gmyooUXTGf7HYZYEdcXNAcLLUorFcwKwy3CCmax9kAjvrV2KVsovuECNeosuGTMH
A72WXaEDpexCDMs923qbp6t3Y0AqXDivtwPRz9vGdpPa4D0+mvY0wCHk7B/efYFl
NHSfHzbGK7L6gVpxbidpnr9nQv1ZTGCHwq7QOPWNewCYUORsXVPMYKho2s+Btfsp
7CM68TP4qBM1e6m0u74jURUOB7Duz1748AYIy3WdxpNtr1bRVe+QYhK++ix2FKBo
7TGvPH9/81/mREWjXxw4XiasBIVdMVNdFnRGU1f8u26dgEtkGCfZ0X8jAkdZUSZz
8b6SF6NC+NJAs/bFqEz6ZyAxnK9xWjFcfvhNIjl3Q/RkoiNdwWOb3ir0faYRLnlC
ex6s5rN03DUldgXf5oP2S9kH3vFGYqe7FJshAdrIeyUaa48YP7yxgIjGuc6mr57K
k4lwv63BfV6QX/lstb96AmL+xKL7qBsyqyGP3+N+60t5lEOgEjFupfdpfp3tfwXu
qMs+RSMd/Al0rtPqrdUnTsk2belBB0oHLN7bEiTxAz+JLV/ZhaqHbp2kc65eiH5a
3fWK7A70m7vkx6f8zwOTmk6/CZs0UBsI5HiWKZDcAyE4LpaVyxe4+qkvJcPhZ64K
/qwVowqvlCXrlMlmOxigKrTVQUzzP2DXoMNaODMa88fkVpU+vjKkUNFRamSYvzqT
dCVwfg0CmsXmctInyza8Ja+edqIzoWjjYrn6LYKxSjiQUjKezZ3RG74/Clo3WE9D
IPnvSfYMWFxOqlz/C1wgQQKlLG8MSrTLvhjWyZ1veC+kDrgFh8EyOBBPe5jtxjN9
L315pHqwjeIZqbyhenGpIP5zoD8noz4/4BgftxYXgohtuB5VWwDAHINcuiKY8/Zj
A+7FTjdXCkKU/c5YOR5OB66l9sdUn+eI+lcYODeSXwpjrTyRwHo7lExye2hpELk6
sDCxJPWo0JWMDo8UBQu+VHNGtvCU49TE/SiVseb8LJQZg+TsbcIWceXEK/+mvPwK
Ct4UdIr1j4TLKFyyO7HpUHWBZoao1+rXBqEsbJ7rbHPFqjNjmcdRfKiXmMV+WsD/
IWY1Wr9NbUikuynqU42abBu61aShyQsaQ7VdJgnL/AlHSAWZsQ418CH6riwc+ICf
a7PrT82QcR6wyIqFAkJDlHMDmlfSHljIlIU2+qJ0C1c8GHSUQoGMYzdV4AFTSSuJ
IaRXui7GwQ3GcLInqdx5PGA6BoqWZ+5NesAtQeHKH0FfJjQ6BfpGK2f6yC+61Xfu
GrZrAMMY3uUDSLI2N2zUoS6UgL3QX40aCCB7PGBmXk8Arm50RMrF9wTTTiGOzoLb
DdwF0LzZqy8bELxM9CVcukU1QTF9FRVN+liBKBbARfQsZBVNIVCUXIgPE9cH9jrO
26Mh6RWgXbeX4MEpdwxRkOr6C2Bty1fSGDKa5ELNif8cdeW96UsvpMMqdS+pVdBz
SbSN3PvU92CHpHQuTWsBcWXVulVvSPLnCLPPxAr82Jb2WzD1/0Uv56Ot98KpLVQ0
Vuft6bdiC4XDUoZ/2NGGmc7nTrcDyCXJkO0eO9CeTFNFvrQureJiMUQrLyXCs38Z
MzIuXK0RMLBjidCdcL1f7NvCZ/aiMlC9U5R2fyeRwHKEBS4WUMbnd8g8RgToEH9s
MhiZAoo7XaxYRNwZLd/jk6UARFeIbuFipWmfrwjk7dGctVa+2lkCzEsvMxSbAvdA
2md2pmHUe6FASgRhYTR8+vExhCNzMOBLAKRTNXJN+CqZ9lIPEjfJWiH89smikPi3
Q732xv8DtCmDRWr9AY7VTBu0dVfrtS/XjTnPWlublofbfdSFb+H1ieviILuWal/Y
/swJC/sktdGpxqooZHzKhxRREggfox48/sXTv0f1B7EJ8sbxtuzmLg6Y9Mbq1Jv6
LfiTBvNCbXa2rznsRvroX0ENjmAUjQf0FOS+SIp6fk+VZGXDJaf358uBbQ6HbdoW
9vWpGd9gQpIct878VmG+CHUt53QXdVz1pTBGYnAqTHtfI6YDlH3WE1tjV2oeXzzS
sxiZHsBBUuWlYykrzHkSZ62IMXCA2WPAUbNtVqbHzgNH+++a576OWnX9bweeoUI+
nJg+OZ6Y9ECDlv9BDbqc4VkMcmmaq9cJdhuQ39ifikcSyn9VSkvjnfTXT/LPa4ML
UCem0obwe9s+ysmpK69NZjWmRadK60wGR7AmU/cdjsNdsjzn7I6ye5IdFvhxS0JH
rhSy/l47idNzmwdrsrqkeXqNj7Ed0lV1fG1iF3Pn2tb6Swgm1Oo7vBDfv22YfEI/
EVgeGij460SIBaHdpIIFWpU8q8SEINaKgj2TXaNrpDyHI4UgMJNT4of99Emo8lmn
YfB1aaEK5brLhtmehGKAmVwjk8KOgBr5qAZyx6jUuC87wH1x6tCaS+nZ87KLv1Ep
ZIjGEmbheaTP7+RAm8neYq5TN2QOzRBYoP3CBcbagqyrKiuXIgDSKbpuPNShCo5O
tdKGhoBzlIZakYIL0mFhUyXXy/BM/bL+eRXM1NyNI5fRMhDdsufZuw4jh5pRT95Y
Nkn3M7yGRUL/juqgC84AeeUrSe6OYZRZvkQLHEaBIjBSQNNXNiNkRtO4gFydFi2E
KLm6zhY4ey58mcUzEs2HQ547XWpF6phasqZlw43TtQeiQJlZZqaGZCte0SSt90CX
WYJBZ3UdBE4bvZTzHrVmzD7FlAVABIwR1HVJrJWMAd92wX65US2qBQ7LAlwc3tPs
zUVXjR0F2vhE0FsXZI7G+0zor3LCar4z/Ep/xzEMdh5eaOHUe3ncZYncINvCu2US
yUMc/nTtVVeWlmnnF1dZF9r6VtmkAi4tu8xqVgWRfsbjCxTVEVMJLgef/nA3Kx+0
PLjaece5iEOdchGR2+8H9w0bJLcndN7R9Za8TmOncS19+VferIDjTM7ivD0hyfHf
DBqu2ZxhLJ1gEdKSkyQHrtEPy58N40IiedTWxvZXPl48EJbY38P97qCMDL0At+YT
qtrEZ9SWnb1c/bB9MSwICouUUnNbVT75J1iHfLwA4LT6y1Tr3XGGsQzsEVS9gYqM
AKFMvts13AlQR6Wg4UFr5+Q/2TcVOzNS6+e0RLqkX0f9V9oAgJdxP7Em3VA+ZFeW
vg+3DL3228wjR5UNfDMK54nSAT7RjuLltremWAzoW0Muw0EzX7Pl7mM/g/EqRPh0
nlXseR8plzWlA6dhlZBN3yrtlwhY8NR+fQBU4VxmtTlFWk/9x2i3dGvZ0oPttvRw
q7FRcSu6J0QmOa4nP2oL2ODvDZNVJRuTz6vkrE+yKduQGwtfxzyGiD6rIeNvWRjA
IaBtBFaPH//+lCtaPbu4bRQcewDh4oI+rstFIn26h292xASfLj6KXjndlUIXZJdO
cgFveXZMcmrc3LYNBm/ChO4mxptAXfovvJq8Jyd2Q0lwg2IattKgf4Ymx69Lml03
GZeKNsFm32Nz9+YpcbA5i8UICSM+gZ06c4Am9lBzMXrd458TVD1CWg6ukjGmNlAv
pU+kbE2tk9AxPt1VkCUi9ProGtqWVgDY0UVhicsXhSjMalwmPiN1SPBIBa66aZCL
0ODg4FqaPlF0ZBrKVcYREKyhv9WOE+nJDvlAStUQBc8ZCoSPyOd1ijrHG5FlKukE
iSvxKpa/T4NclpvQt6NUz7lj5p8inMO+1757RBcxXMQhN6RhVJX/9SCJ6kqk0VW3
A6Y5u7R3Shra+bSQkx7cPRDlWgRWjf4wN2EKTOOVMhiBFmf2Inhz0BBsplV/Uio5
4d2hBCxWwWXj3O3Rlgg46BcFgLoKX/uugGCCmp6AGIR9HO818oeJNlPes3GH0yJi
SaBtpiqlg+YZBAsPYQjaU0LoIuPMeQPhXhs/Fq7eIwfIdFoxc5eKUDVdgOdS4Bxi
Rh0qcaLWZE66k8OthlvvrK+NvixRrFwGCA0WcsGEvgzAwRXvDmPwmGkVAmiViZPD
X2qrgpQGBw1cOTTp0qfu8zllVCFneoeCMqPSlSrkwrAYb2PeBQeaDYUsYD14Hc4V
t+f1wpNa0hSvW8n+c9ehtk6PDoyD+NNorf1yjY0LnEnGP5+2LLXwYbWAm+H5cGgq
XkPuGBzEGueiOg49xxHZk/pDAyu8lDVNPJmMbzWDxmYIIlZpPIYi6SubKpgLqUjt
AX7JbVnVf4pdvULmx0+iQn9NwOn3o/lJzjifLRHeqEOMwj+DXdMhw6RaWomialSY
795GaC5J4jbaHm599wNxyyotqu8dhQhjYQ7014DGF7Uz+DrymRSgqromiyAqu1zn
in2hsz78Op59Fqz4yqt02bUhfjiIWmJl5htjI2XKEoBEXTwZV6ruci4nB1RdtlCj
Jj3JfCpjizQJOJmNAFKCrijhDH7mhPBnWv4peSroRY8QVsNgrmLCiNJSpnDDAyEQ
Ezly1A2uY68YG+jBbyhYEJlDp3oC56GM7qBeWwJVc7rF/mA5o4nQmWCNgqnAoGW+
FRnGbFis/WdqWcOrbiBUenjAUs56zb/5tz7GikDJVBb6PmIayfczfB1JaCI+343Z
9F6CvHKQYVkIKmkSGqQxTWtyKZrKVlrooVp87u7np9ThH/cJAayVuZBgG72QIeAd
+aBDQq71Ufm1Xre2yLMuPf3Mm0nuIKAEjGJhfB3UDmAdm2RV/XWsZFV/Al8A/JCR
akRy8o2NOoA2j+H10d8PHXAjQbbIwsKd56mCqpM/wqMFr4D8N0EEJTs15EzlbZSA
ziSXKwFm2L3AHUdjiYv6f15rhPgRZsmLC+Xd4t+xzF+36H3H1MPNvCPX2LxfDODj
g78T5gfqPM+M3lWTpJdmnjDhVwCdgoIx58RcNwmmG5Eqc8CbtKpN5Jpj51xsyrlb
0m4mkUxq1gHbe+FAmLMx/2jocx7gNAZo8ZkIBKurc7efRRyTZzLLq5sF0Gc5sfc+
7fV3XIxmMNvTSCHJKc+QGWDIFJFZPGHDtpTuTPOJLMDOS8EVB8JuiQ1oq4abLVqC
7R8Ggom7OMXQU37kyMFWodtWTAGMMwuHBJhJ3teNiCyZ5J1GDCkWlXEL6Eow8Jl0
f+oFty8SSytm68oi9mzFM1jiS2dICoOLzwk1agjWMGXVdQw0VPOHiQbh0R8ytPKq
wroVvpBT3dLCHzu84pFAIyPjvC02d68bBA2w0LDW455s0lo3hHgVEL6/9opQqh+O
EsfQNJTgApRhjRcV5WyGPtgPtSe77j21TqkkAoD07t6qM54rWpuLBhSPU/ASpK6k
suCVWlFVtVRuA7/2f6fVA+D9+2hMxmyKn2aCVj9PLHRmKSw1s7I3lQ8ecSO4JOrf
otD6U/vjBWy3EAcCwOsUYMqAgEPPDjM4gnLbQOWOj5Ic/i+JIdKZpBD4wAsjHeEu
iBMW2RebKLOA4Gh1Lt4sIpMCrcaazBlWoHIUtvOKRlkU5L1oN81E1q4Yt1mefwTq
QO3Aq3gs5whjFzxzMbjBBpSAQhQtZCyp/3RpncDM7OIQ2LK3aS6KF/s+RPHOadUC
muehBTR62qnD8RlFB9MhX4Y8x/8l1edtd5mHsJRBS4wEK7KfWbyS4ziipz5nm9EQ
2peAdUTJpYNJzNXx0Kr++zUg3Bm/FL1Ztr7qW91mad9NoOmqUguejN2jcAH/xzN9
GfokzhhX7Cdvuaa4/VfgZSdx7z0eVGrTs3+2tJaN5udRQaITOZDZRPcBjitnGNvj
2mXVhQqyflbfu9OKl/Qje1w2H1pkZv849UKaFSw5Yx5HOhRiInUcRo1ZlKQJJCfe
T+IRIBmYwnIyZ2l5jTjAA11fFxt3ARMyN+e5o8SdE8W3hvoEpYmwetpfYLNDYJkV
QfmnE4TxTtSpArFLTvcDcXJGAvvjBkViaJcRf2lesEoTRMGcHu+FtZz0Go08CXy+
0o1c4qJulxFaXYolNPJPtYUuZZHgwW7AhWDSoyaxHhBEPaordb/4Ccnm8NWQR/0E
6Sb9bB5GrWo/MqjK637g6XPGFzWYaucWEa6r5df6okuE/D39TD9JDRW7sqWmviF3
LM1VVche7ruDy1C993+Xnt7AJZ39MZOY4iZiYpfPNlH/qtlG/oezCptVkiVpVVwe
qA3pCrFZD6HBBcnhQAsEIBlMHwTx8fSgeECJh0gVR3tLQB4vxcB2iC74wyTLbgBK
wBL9tim2dsc7uYPZBgDX/3Aiame+5LSXQEXQVjYLIXd5+t/r3tMF3NKGj29/53Ju
1HY7QsXajFaT6yv6ToRF/TQtDo05ZMglSTH3A+1tdx4nyrT5rUgJ0oKbnBtr2mOR
Z9TGN+FqSAxXgv+INXmauUGFucF0AJhZyd/2qc/o23O9Db8WGBVoZMEbWuyX/LOA
yZUYRlegRSVc5pcsdgWCvQAymGOkNLBEe4Ieiv25HkonNVYp+bfbRqlipi4Jd1F2
Sz5PeYZKsGkEE4+OMOSTb8NWxUr4CC1LzTpAScjHUToKuSsp7vU2bXTaSIG9n84O
g0ssbGUXDiW48VyA9/7+oKfBFidPXCp1mRanjyC833MvQ6q/kX6XNSqVJrUXHAN3
l+ywPKmAnPyfdKtynJWTW01teckIAmWQfG9TVoUttntm8YeUk18CjZCNL2dJM9mL
PWwBYXnNJcecFt5JB8M4kumX/3uNUyTT5QNgIiyVIz50YvKjvxm6dUy/C9Mv96sV
naJo8lqXNwnjHNe9zlARq1cfiqxBPF7PaiDnz+nUiOZ6iaswM8qtXNkzwlhUEiBw
a2bn6P6na1gG8hCqy5KMbOMJzAsQrvZ3m9EqROF+z4uVrQZPZaznlnmZHqSMSX7P
TSGjY2+obCrMZ7B54ahcVzKtZhs4Zf+w6tIRVIFbu0uvddc1fxXAfZ1Q0zTv+ufQ
FEu4b/n2h3v2TNyUxkKGRjfs9PAZt6MjnqaI4RtvTyGwMrjngYqJPVO1LZt3yTGQ
uyy151qKOGO7OYJhJI7HVXEqZXPpjzn6e0p8BtxB4aWNtAj7jqcZ0EdF7yyyUSYv
lETCJ0ClFxme0LLpRxipsAT9HeZNkiEFQDEyE6pFeaqjOmG9tH5WctqjsgqOnr/A
278vKT7KRK9v/RlIVX0rLuD6Qib6KiTK7fU+0SXpjRGjVRiFITaSsqIhr62ypS67
nYJKfl9cLkt1MiYHhZUVl1CouFWkuxEaZiXMVPLqXFnE/Jay4C+3VnSw6LBk8rZk
xzVvAAdBRUFQEWxhXGmXDF2CSP4JWb6L3b0gP1Jgz1aXguGmI9zFDD+vLI+ID0Ln
69RwDs2jwivzsUhoCUG92SEblen7fk+GH7tqBRh5yUbETRSnbKWiY1GszdGvnNde
kWzk6A9FPRfTJqHAHf38pN5izIMXi3FiNWzdFqPq4XXNy68hqN60pTaIJo/S/Q1i
JEacvtnXsuJeOFaUAV8ZD0dpO1Sh2em5Hsvz/rqQZuSlj5EQer9Qmi5xCSXtL8Xs
rT3EB7z1o5LtIrzk4dcQDzv71uLe/zBnQV9CG57bbj+BUxQQFEyAJ+g37SEBEsLG
kowTy4LrRYpU3AiWVuJkTLvkz0KPtQNTkQPQh/nVr/eMZbksG5idmGOAmmw5Gj86
y8DDmsf8US06fAAm/x6miZzH+W4JhejPhpXdHY8TU8JjtFtZ7aOSQyBOmnX0odBQ
mRvVUbdlbMbMsMb4kyEIu83s5zNQFnQFXLyeiRT3xNJfj6luGY13ouf378SI9eqt
A/+LYHNdYnyhD2pRJQhndgNIC4POfsAhTiCn0nzpQ0kkNogMaE98uAs8XsuJQbW0
WCvdkUO4Mhxj+POVi+raTFuOTRpkTdl3XcVZGkYwwHxa+2T6gRtSWIPRrnLWU1wF
o+YwovvTX+rzesmlO2QU9PN//7yLDmzsKhX2T0CaZWLutq4zYw19+A2y/o/AvYEG
15MB1BiJzeRxURGuNuJSwoDf/kdGznlZRPTUQQ83bKsnmgdxkRW+6QcYsGaD8teD
BVZaKCA53Mmxtp1NwSQxC5c2TlEQdpKQaKahk3BV4XVFPK8l8+TZlbgpqyKTQXYs
YefFyCqnHjt8wCLTzapOYTy8dNFluAgJMpPlJvgehf2KRXk1o9P25YlW0y7nh2PJ
4L5K0/UBbt2nZMHRB/5bk2Ms5EGOhLfO9/ePNqnIy2K8LqUWT2qoBMEcmzB4xHRB
8rBVk4x05XVKW6iB+iIjxiTfuIbjLdb/DLMigzInPT417YKtEmNkz3o1Do6WGjoR
bD764jXOL1XskwaT119FrO/+E5vvSVpDRZgiK/GSjVXKDwvrjWdbVZVxQ+ouN068
Bbg9s8O2JZ8AOOViVzqlTKp8yv5R1qAMU3XWR7MxYE4WuFjQDO6kMnNJB9RdUNBP
HPpieyZ2PiXTMSP9wx4z2GCNNbjDkyaNX+JzUT7SyM3Po8I8QfeJTp7arAGday9P
UfKGdhS9g5okpx3IZSixtf+xZ60MasyxhCmBi+8X3hjQW3UtQ8f+cOn8pTMFRR1B
Gl/IjKNrC3ml3PwtIdfiMxip4PTa98x3AXbbjnGPjQ4o/FcWmFnVZTkx+ahcLBVQ
yCYUSB0a6G22/fTUqnNeK+qkbpm4ZIY27j+VM1abJJqRMjcmwn53WnbnxALBOpCA
KBmd9jp8T1HuWFgOhZGJLDHvSnHfHMArOndYHx0o8CTPKBjIy3I6XgjQJMTT5hae
b+FxyrvlFC4K+z4SrbZBn6N2zWpWmvBDT2kwRG18Pj8TQDv+rM7ZA5sCyHfb2a4e
5K+LY0boSHh7ynuj1BKG+Ek2LsFd9w5MF0f5QETxzBS2nPwlL5+HO8zPuoTAuL2O
9R9e721p9W+ic81C6bZbFRnMXz8AINCo3rFn1Y2MXSSTNtNxco3kb0tkN/x5v6gN
08l9eeQ7bUySNYNcA558+h3vShgEn2+wc7KFf5CyFMqgR6Z4vi96wuX1TYfHTlrj
JDSB1Z8CHlia/UcUT2YCB9nU82YvmomisHfN/TMqoIxCX7n6DIPZTlP/bHHYHc9m
PymVlzvX5NekohzyKxxnLFmDhGK8J/QWWXiRkPjuhoXVjM8G/CJXdzefu2BnvCzc
2Yq4607OpCTwDP99aA8RGeYugntMWuTKTtg2vNmtY4YLZk6dXcdo4m8yKfhiz2nE
+lpy5xPKd10grKSazc5iuo1iv8iSSMzOXsdxZT/7k+qW3Rti5nV+nEAiE3vgD158
fAHwHt36EgK+t6jyHI4rFAxdeewm4dWlVE85Ie/kj5cSWw1NWig8yEy3EGFY2QUK
aoHrr6JOWZYijpYlRL4OnNFiNJyhjMNK37SVbGk1jwJZDx/q8fAJOWVYPyp9yzYq
30Ei+gey7xWiVxQ4/2dZkHTjxxbzFxHfcKbPbfWGbzqGs9zJkqjYG/tfLp57KOS1
CIPBc+5IWaAAKqduOG+EFsejgYKmToASXcd4E4w+875gDRUrrwm9cK4MuOz64PAE
C/ifAyi0Avs7OKzDBi4RH/zuKbTBTxnKBUDJw8Mcqv/gdtHrn1ETZTbxIP2upY/T
jsNqmF5Lv3ZRR3vAJDvyCpUJJUizWXU4i481J6UBYMF5apqvMTuf99KdLEV/YM5p
kT5a6sxVLroV8ThgE7gbWZCvmxbhq8HEQhmlV3Hg21KebzB9jxe/+HI9lDbY6/xb
y1SSG2pmmC9yRyyhEom8X9F1Xq6rC6d/mo8YrcWoBUsgwEg15VTlcioMlMgSGi0B
gsOey1jE7gi5mrdfHop8GpU82RVBLYvc7j/9KGfePcQQCfmKAFupaF5Wj+Mk4YfO
/qoUSbvx0q5pTvztgZALtvpwzvIT9BPaTK5alA5G5IKjiiBt2hs3S7fzKa1LiwNb
aiJ8a4UfxI1SuGtJ1KYRD01E9WYJyWfmZefBZCWl7MsACA0UVokAbFjXS6oeu2nM
vKOgs2yZ5iapcGsyftrDeCzHFxONgxPuSUzi9aiI9zxKL7GeqQdNHiaKCi9YcGCR
aXZz7gCtOa4mfsTi62xI2RzoE1J/QUuq8xvuyAuHBUWtM3GN6tKPT0B3ebUWxa4C
bLmRvFQnovu7LDZGfWFZHf4dvsl8lS58Ed46XKDOa6AnlMOG+fKgOBQslPqb1XYZ
lqk3Fk7TQBV58tHjHtsR9dT1PuRLZfZ7RQrrX66HLWG6kM+exkkFYcCDrmvtYh5+
MNu2H3F0QOfc9CiQNqwyBDB1kQOvzMmAUp0DhbCUhMxjsi9IV1+RSrj7ZDYmAaSh
6YHXvsrslQdDSJTiwjj89a+UNI0FSnhz5WTCLJE/RqSZYqOnRjmBZ+4lDPA9czLE
WNG8jmHiGW7ET4gEAMAmBzJer0FvR7DJU/IKPIdN8Ipr5AazgE3ssOolI43IQQPH
b9waV1wKJA0tNBgIKT+K9h7LPMzs9p2/MGITw1Gp0E58bIg19FCj5/6kbopDUd+1
hCFe2AOs6FkqIwWAeU0DBwUQ2/gbK58jgwgHmlfaOjWo/iN0//hGiPxvpf5TztlR
OeJFVjGqDj4yPyoOqMbtJ/8fl/ECvazn7HLkaI4R4XESs1gGRz7PoExWSPqi3XFy
2CxcFOOfGHR1yqNMuYtCZmHTinVdJc5dhBey8X8U95+yASd5EfAawVkWeyPVrl4e
9EG/fVi+q/rEuwNWFh/tTYXwZDXgnvAiclK7pLzyLDkE7poKn54lxdKu1Oj0DY5w
UTbfyfkZ6TQRhc0I/HiWxSTJEF531yI6w5G4zU1bdlGkpS9D7CnFhrIYv5n77cQJ
kLxO44CdIRJ5+nfPIDqIzWyQVF8H/RwmgEysw2XySkChhYFttb6YEItvLIBolXD5
qPZxZByMc6gukWeQ+rvmylP1/cTbDzyEY2quvn7n+ltHdyOm2vx16+5uN3SOO+MW
nXv63xKA23U0go64/k8QTLduOQupKKe4E9ZPjrL/yQpC5AWEDu//xrcmSk5OojOq
33bUtKS0XsS+tHH4KzczlZsqAXg/AKC63ri/5oLK+j8Q2TLvlMo8zutrbHZMTKJb
zyVcbtmVzczm1VI7usx480LrRZE1xCqgH2vO+pQiYcDwpKHkXzlZfb6nDaVrUmV/
pbZC2pCxOE7kKLSot0wNj6cR4OnitV3+NAeq4tRQ9siNiLnQuOhMLFEBYqXQSuzs
/APTWOM4TuueV8BTXoT90ifm+qTBhCdZ+LSPNq3f4IBQnt7yvI7C6rS4v+lzibVb
xqGvqL3H2vxunqqCE8vxZiFCu7I/J5WQAoyCankVExsSwQ/4rrSOiksdB9++b0PS
ox2xo28LGJr5Z6jZsLNA/si1NmQAgX4LkL1x5kh4QNvKgykBx2QsWNh6AvvBE1lv
rK6ZMcVq0osdIfb8VtLyEiTzL2uYkFTQ4E3PSKRGVwkA0vzsMIcGS4jIT1MCEe/G
bUBwgnNT6pDRAt/k7UwOF3wYl4f8nEUse+dMtbuo0maNsViBLkrgAOEEM4/hKEr0
XbL7w8qDV8SowulMdKykK70EKB2VrMbWXxcT4SELb464L5aBXZS2t5anTOfqVQvc
NwUMWQs2RiVQeezRYDKxM0t64jPyE4LqajqI68HhvFofWEe1xCRu9ORYXRVfmCcn
UfhTAmy5fAQ4hbD3NwipYC3I54CX0S3/rfDlKdzpDoXiItIkzSBJzlBMtz9QGBE6
ErmfCA4kn2wcOq4dj+0rsbIo0gV5VQ2ceqEwxllyDW7GJtpVJnpRxpsv+gGxHt2/
rxvuOtb/zoxx2fjmbHyRgjdouvG4jZRhMcMtO3ggCAvBoH/F0XvKz8FrOYGWm1CE
MstFnsGUJpTF69CVAYKs6rIiK2171zk8MB9KLFeARekyn5WMdeJdvFxHVNi3zwvR
Hp2wziLdiI3B4pBswmgYRdwOUYPFYfFjhwD00km7esi+j7NvQZuyIG02RwWvYePZ
NFoCGhB8PFlY+OGU6r14+p1Ifmdiq/nKWyKRpaVTaSN8Nm7q15MHmzrqs/BiMlNm
+7vjyzWif46aHSIo4gWWkjX48PxI7Y31bEQiihICAgsB9A8NQJQMSas0xpeObyqy
xcZ29zTUd9owb02GgsN51j+RpQdmUPrxfO+9tXFT78iXk7nZoPppHu5DYV9m6P0B
qYMzzX4TaQWZ7TTN5ztDO0QN0cIHyWCPt6nlg6WDR0i2KfvU8GnL+PxOaubbythk
2DR47FhDlYFrTSZLcgY0oyR9IpDxjAVn4y30gdHuBk07GZPa7sYDoWb9FEHHgbOg
PBGKu/lnLYAg1QagUSeXgodc2LJLHQSTr59L0WaKE3MzoCR4EB07LoikktJ/KFdh
IUGB9xqy2+3tj76m3E/1EHU0cNEhrP2TDTLqgR+4WyLLq3vaUZAR4Rwq5FtG51gW
diAwhSbHSc2723nCFQRlNzhe4ywMPc+seJRqBCS51cC+iZhqOtKUYjVaxGmuQS/D
M1dZJOLibTXoKYcXxz9tmEcF99CN8h4cv2fQXq36p53Vk9Gjr6XMAtb8+gS6xIlU
vdtfjenmtV4w0td5EefQ3Godvy4YyyiCUpQI89DJ84upeIVQO3/RTxmOS8vZAbaD
70kW4rWbQzGNMewS3HGWgA9vGFmbveTnqyl3QqE0yuaQuq/3xNk8i1Pgd5vTWb9N
egKZr6UAsPbcIZw1DYzROZG4ofWGIhAq73wFgvipqFjQ5pIkiMRaKgZkPRMi8qqr
+5PCrPk4kZYvKp7EcWlFbBkTNwhfX45DQvCFxa3Pa4TRoEV2+kX3Fal56/BeMJLu
l2oM9dI71lderqGV6jHTAoqGiqvqP5N8F+SHiIWAc+Hc6+MJCyAIN+qnU74iwCW0
9i6htSsPF51wuKEFTH5EKVW4RK8szE3ukkp8lqaf+MPxHA/q/ADcqzkdV5O+/4ja
bqhanfjNA1lrU4uu4ISgttVP5HObEg5YqkCoG2xW0lhMizVgUrBofaJ7djFIminA
fs/vXwaSt+L4RQcb597lKEOs5XKKeB3RGP8ETBfnAk2ZmKvwKHgolwEcuqDVA6W+
UA6XcfDKHwjuNtWF85l4xL8yR6ZyJHStZInk26G7DQYzSFSVJaXLseMuFZdv9IXU
w5nb7EdQ7+zD+g6koKk1CNLfjJYyo5FY6XtACAWneX9qxZojSzhmT38TSpmPrJyr
ziIWG7ITVEiEhUN9OEONhrZ9zA3hrTQ/rer9Xicbdyrz24iQY6dsOlNP3lhWYI9S
MvrI99oZZtLsP9mFFsJTNvIuUiYtvLHjheVyVrB0eJ3SebmV9XNhWRaiIvBxLKi7
/4stcImIsPEQAajWKtw1qo3LvyjIe2rGsxWWFVks/osrPkAmCf7dEeUOeCPR7PDg
Cc5EogeRYfMrsLe6ksVGbrlUfB8PLeQT5bveZ3PDB248pU4ep4X2nKSlv4f6IV0J
DZ0NBVe8fhRuw652X5QarVxqdOx0Cia/w9ldhCDGeVEN/E/jGh78I7PGYz1MjXMr
xadHV7Fct7yAxWiVwYYk9J4bfxJ3qqDNFCKPS6bBqeszcRilRvMWdAT1JjqL6CxR
zVPpkqidhDTLujskT8BX6VfpUDZJWckTHLSV2KZqaQuksQIMFARoD0iatP0hV7eS
e9VnYlCL9Rwo70M+fdWeAGvGFJaRYjE4TkCiok9hFgU3WRihWf/y52PCmsP9TrS8
hcdxTrhHDm8XB/hfJRXTr2nUchwNdXMunn9y9zLeMJ1VWAlo6CbXHU6+TCE8J6dZ
k8EzrURRIrHC/DAUdX+diFYb0MAyCMQODEprGXnqNPH5VE6tqK0Oh55mae3KFO1H
czOxaIym4ccjCInenCBa8fSuqjQIRhHizk0yENX1MtlpmkS3aNXfWlVgECaDeXQs
sbfWsmjga/BR/jpBqCvXAPS8mqe/trGVsIfNE3gceztRNxEejmKtfif2qHwUrwj3
25kd42lorhN2AkB263aSI4Wi2lEECxUesK54BKuzmk97qkbOfB71gZjWe7eu1bwX
egyqadghFKOkznCrodHBwrPHgfL7hiZlfIlw1UZY26VNoq64pnKWYIxjlXI2Hews
pig/VfpTMY5NGUb5/+KEjDenwsQBUMJvQuiy01i50AlyZv/gvQFYUgM8jpRtl1k+
A7tZeUx4OvY1jO5ckyIm82dLO64081eTxSjO1zc+GHMHyz7DIplXioz24hOtwTCw
IJdaSC0jwC8AWS02ktAR92MalFu7YeWGbT5ftL0tp9ecF1rdQWmwh6nHXVq5r6tL
21Yfr1YSby35Z/W/OpSTlUOZSGO8mKZBC5o/K4ToTitzBiApXxahuk2EUkrHugi4
pnUevz4jKY+s86B6Pnwsv/Oqt4A9srOKBPcXZUGq7LzlBlvZTQbJfJ5RLmTX63lO
djsmwWYKXfnoqg1D+HoGimnYwOlztMBFRVYzz5nMf2tnaS5F11GUaT+P/4cbKGO8
unaqPBZ2dmckIURLDOfl9hDLujzEVq9opQddMN9fZxhPMj9/RA/644rY/II55CRE
tld7cJbV++F6fU8AGuteFbG193Tyk01IEsMyH48tOkefi1Vt1ALTG3qsiM6jGPI0
zvMM6d1hSdhZJP2tGAEvjgrYTiGzYcdttLn9F6ygsQD7BRgH7uK+Li2Von2kH/pA
Zn2veXyrnaUbToPnrXn8H5VT6pyaarpd1cUY6iN1pNPcweU7BjLU+i04bkFReQd4
BjTGv6QsdovqNzUH5coAskAu/uchArNvPWas0zFgKjgPT/lhGVKnVaJ24K8zJ9My
fn/XagSlSvTrH4a35jXhIDiBGXWu3f6zOflzHjhkXHDNlX862WZPA8MPmDVnVKiL
vUlPC1xWQiy7yrmDxK20WxSOKfSjDL1mdbVoLi5l5z+8P9ciJW+EBrY6mcr/8MyE
56Q9DTi8tbobaE/HixUeOhBzAy1ty+gd1uU4MkMUUBhJdxrQL1I0GDFUnLzJR0YM
4wFwc7ft6ZtUfvpGUtQUraqUsAhvOqzYsgAloFtxtihunDCjJWB5CECuAsmQqHPu
Y65JcsOCoC1B57khwYb5iCQCIski7ApcVVMiB6oIKlxlRR0ZQNwJkzlCdlOeWwB+
gEz+qX4wNREnkPMnB//OkISpASS7mk1LyhMNYmm7vqL7OvADZqIVGFgs2PgGBSMp
IEEp9j/UCxcCC51APCZL06Yfd7aqpDZQkmiGnI5aUGmpdybjLkmBRTDO2kRMy6Uf
ZIE5TT7Lquuh4DZczRTcZQY271G1ZgzDBQi7/b4vc6Jb8v5kX9nXkWvytimMyLdB
qLNvZfKaIYzdhWjsDA3qu4BrMmSSrS4d7iacbxBC3bp7bv9APfGuGLDY7uIiWvYA
16iYDwz2dVgItvK0AVZvlPzRtrLUYeTIc/5oUHhgtkrFjZ2qiarVibbqyv7NKtZ5
yrNX/s4nhYAcRXAqdoj71KI98O07Nrfvtj+MMzGY9QxbKxdwumCS5UZLSdj7+1na
iKUBtz0hwdUZayfOosuVGj0rgsM118cYbegx7d9Plr+zKjsQ+cRnYrqhcmhwXqvr
OPtM8WaZrwSsE7Y4nnLX+FZ3T/n0hRNjHD+49YrIhOj+WYBFVPUiBNVEnYm8RuvX
Wf8SMNAT573800c2gdcOHcpJ40lvI4bDImmZZ7OTTf3YOb5AW2YAtv4CjyIPDMfu
WU6YJM4V73HaRy3YS2WUE9zj3gIpjnLFNggJ/X5yddPhG0pCvt8h9RUIkkuCllJT
CyYJk9YCC1+KIzxTrtYC9SwngX0T1lgK5XwRF4+XA6HvjvrFa60l4nM2Lv1xQ17J
ufPgtE7PbVWAaFoBPEtAzIQhU55as5NUVPzyCn5bLex8aNGakGwWcSWSCgRt+ZB1
IV9Hc8DjY0N3fAiGOR751zbyhalkBkNW0VB3a+32ONVs2H2TDSZ90e5qFnGPpFyG
DVKvAKjfFqFmdvubUPx3U/Q2bDHdi7Oa+b5ueQuVqNuTSQgEf4vE7XBoWSBREwML
LXpYV2MB6hN7pBa6BCeivIbOB3wH9uspS9YHRg15NBr+HkUvL/alkBhubHzupgBE
XgWjKZdvXbRG3eBFezsX4ae33mqW+++bQlkT20hfAfFswhe4LvHodqoMAT3/V7/d
zZJGGxvOn/pf+G6Lb2Wg9Whm07epwslhq4z0uBsRvIIKTSPhmxiHLw1V0bmkXZnC
NBCaPnkoQ+61JN2ut2RMCSRwMjFGH7fdIDbhKuKntxnmorjG75SqrH2BxaeRRpGK
1U3NacARcqCKi5XxtR+mVq6IXhHa7N0I8NsljVa/BTA8ikdlgpobJ+HrSbiLtYeI
m0VEdny4xGfyOG+o+TbESe+DIrEwD6G+vrdJgfB9Rz4NtbtX3sI1KlLZh1r8TIrc
DSmgHWETY4NSw15vIoDq4FM9k8/4qvOQVNrtAmJFVrUym/EPCpaszY7b/lfQm+ng
jz7tQwCA7sX2KxdIm31wOwVEtZl+IzCQSoJLrawKxrRR0+tB9hl2994V+TOjvg0u
RiU4qvt8n0HWoz+K8IIzVTPVLyg/4guf9c9EoNVBnjhQIuhCkNteeHYDVXLCks7V
bca27EbxjXxWj+MTgSUtoVLzmFC+llbhpVCy4EHSPW3fEh1eFpNK+RB9dWDtaoH0
rVQx504jcu22PRRaV8PbShllio/dLQwPGQAeMHDRwveQCdxrpE/5vtMQZ+zBfy8A
554NeWqsq4s/1pcmBIDeccZMFZXzNIutjH11P1U/370RrwUmvtdvFwgF1zM5N8KK
b1j6GKuG/LT5QBa87HL+apvnuNJINAeE8GPOTHOZ00AOWh4shhZ6wx73IdoBgxqZ
3+KVfuLKBJycdYqPNgStPVfrkasEKh03AXb5KauRpfgDV3Aoi4jsDKrMeMhGwmuv
XgiPkEV1Ji7tIU7/U8Lsc44R1D5fUQa9Y3VCCvaVl4Ms/2zxg2cQ+HLpqKyaDs0h
yG0FJqXu86a48yeJGA8WO48sred5vxl9L3Qc+sG2lpAGIXW35LypotKx2Us5Hd0m
7pnO6pHynEuOK0Xicgq8n/lpfL7q6CZ41f7i3KSrDplcLBqdLG6ToPEV6YoVvQrh
ze7dqI/dCUYq1z0Zd5mBQ8HQp1ukeewLGLh1Ds3vnKECUvyMFl0X+5XVNAk0CvgI
RYmMslgftf1FthOnrNE05od8DvpnpEUKb7TVtNBPcIGTY5F1PeAz8++3fWZdtPYh
L4m8pIYGbAWgptbIxY98bL8KBFalN6ahKaouQk23sENcqjlbDiVxPTiqYVjLTUh+
xTMNmsksbE7oo+FKCPacQbYrMxnEFadxI3zZx9Tuj308+7sa32ZnE4yJaQsDeLpn
umdvIVEtEq4a8CmgcR4Lobe2t29yPWLLeizNE3o3YNOMipiPcZ+EIu/ih5wa4tDi
TXKmQgqDP8HWqSFmRSgs6GZdhkWkR5h+QoBm1rbAcJg/d4n3IHaBU4dHubb4wM1i
mYCYDNcBMeJokKYfFWJ9BJ2diai2yhPtz1IYDR0xLBbYg43ehbV1sNRtYrC+rYeA
mC6JtKzzRhmiF2I5syNu+MBIYID5F/10CgcbFWOQIx9AT3PHF510RnnqLHMVHrhO
8GNEgdMwSUgRt+TgwFoiRsBUXLG2U5KtHB0Cd38O+QEGuE7J4XHWz8le2zsqcv2P
prSONxSkblBbAXd6plOEsVZfSeyJp6YGESFEaeCLKfzNV96pBFfAoaUVX+Ir3OI4
IFdU0/Ge3Sf4fylcWKrFB1g1ysI9IEyW5ItC09hI+9QEtWz1SGrVMgBubavwWelK
TIRSiC6WP/PEUP55dhr6EbUIgaDF2Q6CwVBabEaOK37loDM6ic2fVhir/4ed0HhU
G7TvMaM4991RFVpRWAVGVX7apGsqA2I3vGA8Q/sJcQuI3JWS09jncpj82MdxX1J9
B+ebzbzlv0p0g8A3nUabhSCmDN+iKXLkF5PiWRMx65enKMoUXEwS4SxgC2TClG4K
eaPeb9nooUu9a7Wac9hirOlaxBRahnEA33ERCzNc3BGr3ekA630yunsiNx2z2m9D
8cIrO1ow8xLvfO9LGztmLuN8pH/OleAOENwrvobTYaoJOoDG0QaNw9gAyPoNdFOK
0G2EB/oA6JtpiHHWUblcUilahwTACbediAc44CAj0HB0mDYuSpnTft6Cx+7CWbwf
ItlQ3GieD24ZMBTUIAJCuAIg7TnDoDnqEmwTzmUgp2YU0sG8dgTs7G3v0fzm6sao
iWcU4ILszAgjEe9i+pwl+c0u2Ml4d1FaGk0MboLJq19fPrJ1gdQgVJNJP38B3fLl
XbGfNHBO+YU+iFlSSb5gEiaDEUmN0LOZbtIYNQ+fjAdPwZjRMtpyAlkjLL11/R6J
+XcdHW4OUH3XM3t7K6ZO8sk2L+Idz5rPiVwkeBayvS8IWbCWOVPrnS7m01CIoR9i
4rsBZJ1FzJXmBgt25/gFY+y9J7rMM5Y77GrpfxYltJ/6dEN2K7d08WEmVrPNaqBp
Z30Cgi3u8pxqo3dArUx/auBWE2Qv8kwQEa6McXhLkxT36t9c4B27YwdavqM8Odq/
IQqSh9ddaIijwZH8i6D6/oM24fa5uvib228YXRuY+wJWEFH+uvd8L9SBpXH2tGHz
wT6WIKbsRR3Cqx6x81TZ7v76j/pteZ4CnjjbOY0cZ9+XN+my0ilP65nLcq4/vVHu
P6Mf3VvAn3toHQTMOB00t8BzTB6qQHMM6DT1GkK0pv6BHYj2O51rbdoIDcyDWjJt
Rd/KBY3ZRGFJWKYLFxyvhReIBtTDtGZDDgv7tLIFDg4Nge0vRzPnXh14NynoiXB5
/w40qt7XaF1ALlDUsbRFi2+16hV4iShTPHSX5lYpvJgg5vQ4XGpQzplZ96c/r+K/
ig9wKh+m8fEwR1woradDDO+naBTbJvnKiKvqbm1CjUWHcY/0Iq9TVMRwc8PWVunv
32OSu2N7Y2pTd8i8JtV081u6rErWYWvxpLNRWANzePcQT4WxaSY+ai2irL/+Pgoh
SsHlfxYpLeQP/4hwH0MXGn0PPamQy+fIVOCkXdhzMYefc/tb992VTHu/AjAo7n3I
3VhIPfMc8fFZDpRZNt8ZtpQAqrj6HYeAL4FLDza1JDsEo3kho9BF9Q3gq6GoFj5+
9iX8moYgOCGswAYjYf6kOxSPnXIM+fcp3DkUa2juUcx/L47eyBWuSHnc2j9U0how
nI5iNajIXro5okJjMZcSDOZvvPcq7jy/drYQRm7XIT2eydavSxFmKGc3qislbo6g
bRVzK3mUW4aStG1bWnu/8qVC3SLQIn5HgLtgL4T8q/So31iP9MHDzi4yK9a8V8wP
KROpjHqJsMT0eYfQcVkpU6hJ+DUQCrOfRuUknSXHkS+EWMCTxveOuQVjYOmGaGqq
PSzmHVZf/dxiROf68H1Kk1n6vlXrMBxbiWCd8b8in+2ZMLM6kEVEN5TWdkfzQWxB
q9J5j2uEr1aNF7Ffh+aE/ywSyuhz+FiHW1hRu6joKFgZGkcBZQI0zwHZsozbpBPI
sKDHrAy4cVhhfpMb5N4DZa7mZmQwcs0EEIqZk2AByvJ+C64mm2Y3OmVAj3MZcVGd
zg+FMNgYPOecWvEvcFf9yl6vs/ezO8piMxbIbaRhN3cgDbKVALlsoU2CAMmkVsIJ
GfPudYkMqmE8dzxy1krG57rRt0/pf8357WLwXY4xMGmciHs1zo4Mge5B7it8+whT
N9XjduYMUEry6xF9B9Z25SmwEHM43JQhYWv85d7ZgxtWvJGe5xtpaptGJWam94iT
EkO9+V/N6bm0z8DYr3UOFpaDjafbNOf4v800DTwoiqXme+dJj49IJqMJMkEH4VbM
F3FWUToWTftYhHvD8HTzmXQD4rqUgG8pIEvGS8xKNJ4dS6vOqUmPhGLpxUwmDm1G
1jWewM8iYS03o3MCLc5z7fgpHkzvXLtaTMhLnUohWWwmzN6rtCiOAMRofzd614IU
GFFuhX2mJFOwHikzGu9lNMM2OeUATWZJGwOsnFoWFfKLHzpchIBbt4WtysTeOOpI
o143wR17e6zre8GHKmdsSxRtB6a1sk3IU+JXUoxyuc49IZqigGKy/7GhWWr8f9Cg
sCR4QNtmvPisAZxzBjhSVIiJSX5Gykh5ZDGayXoODM8YFJaOpI47ZhhnDN5W+bJt
ring+1jwTcomVaFxyViVrMlqbLJesnwAIjM69PjrOeGzSb65/zw61L3NHUp9LmE/
skV4IBiZBbnF0yjEHC84zlvkLh/lSYi+xzxZTvsEn24q+Vxd4c/Wrs5uQcvdYaJg
Ysbtr22X59QJs/cclwJO6k+AWtx4o40xACc3aJLZMStWiQHMavBUhKa5hIoV2QQj
thtYQ1VM5GfQKk2Ui4oXSuABz4Ffx1FhBBN26C0oNHayiAfyptkDDQr4dsikRT0A
uCCwLinKFxcbf6FQvP9/fOwvir6E8Y40O+WF3gFgiyxdBCqUvxydWwllFNn6TE7h
o2DY7671s59/DdFnR5r/+HAAAkA9Xj90clltKzOH/FcSjjB1ZIBBBZYX1W2TAiKC
QA6A2BDFWTRgSwbztB4L8kj30nnniczPcC+YmsDY+4SXs+uW1kgCYKiHJx76t71R
owyhrcfI/bi89HnsmSYGhAoYnUTQo81GKS65NVmspOFaGFyDPETLR/T5r0TiVx4q
5j25S8yTwj7Pmx91lmOu5aWs4vOHnqZI6bEqPjKMGIlZBfM8XKVBG5w9p8X678qw
4ZqVSar+rjz4LbbitVZu/22rP2lgi1dv3RYBrw12VApWgSF/UgOumrDoy3gpPbVD
DBBHoULaBrJB6BMFZy+NJd+kGRtDbolFrfjdfnSNiMQ/dNrxzpk9l4wcDQUROz3+
ui0TK3hA5X5hZss6W3KBHT5MHgEqhXqEhU29LFMhvRp1aNqHS3LIibPCw4VpgsKT
fsz5Hc9qgHYMMkm896Le7o/wDABnzv4iQ0h+vyFKqsX15i23yTu6pKgw9Q9ZoZUv
0JM/3lgv+uc9fKuz+zySmacjRo3Y0J5y6cXKCyPIaXnOzxKACw1ZrwloikyZdQWn
FT5c9CK77HvNzKHpJ4/5lPXuzIwMPbZ2JNufzClp5gBF3QLfg+vqftUtUnLC+SKZ
7sULbKMn5s3n6O0CPThYzieqAqEZz3FGvN2f09UHWRXXHNVOW+arr6rq62+iVWf1
88Rj/m4/OsKeIwY5ubPrIWzrnRS9LYfKf4GfwdmupH5hRfj44nUWQp5jSOuS1zU0
nystPEuntWpPRfGpdYvH1Qn/3bDCWT7osmygARtnbhrwhgqPSpS7/Mg+Cp/236Dx
iPE/Zxnw2428hl1hmHrQTObTh42JGA2QsqNoHang5Uv2CRRvsTltAH4Bc8+uzDjE
WoJxvnSIdq8xW7pF1GDKTOD+ClxbDaxyzBC6jo3W3IKnEm5SroWXJ4jR5d9g59N0
g7SC/mUXHHnj0YVibAJU4rqUrEqFWevticRktYhfzu+Y8yETXfO8nSoQNIf6PpgV
YB9NyjEmLpB5YFS+QNr343JZ3jvduyfc+gwS7+xM2Uall33cnWJTglCPXBdP794W
AcHYUM5b5iVrNdY8xf/d+b9AhxccK0VAIKv/tJDTT5swEoLcxdXXf0ykdpau97zA
Fa7TKOw1BUhVSYHqDN20gfDjaPc4WbW1Ln9Hw8k74Ao7Qqk50j6zpHrVBGRwkGyF
tWEW/JwSRpv8mnPOgj9XuS6T0hL4fHaFkL0Q5YkmDTpVf+JWQkGkoxOW4a9qMcn3
QAbGNme4W/FeC83tTe+gNxPXuOlPBWqARXQJV/nyq5zJhp6hWNjA82wuOHMswRr/
IA8Vre5Iv/hfR1bvZD11n7cq6rgckdzOWLxYCHSHa6pCXBekfCb0llHL1LFIpFWI
C5xMtbzWQizrG34GoYuxAgq7Xn+Zl0y0glIY9BO/0ptT9op3ZYQ5w7WnJF4P/sPU
jhKOCItv0SLa8bn+xrlax19W/Ecv4nVDQstX7X7Q+6RJyRZUaY1TCV2jld19mlAC
g5YDzY6UQM34CRSIyHxD/eTkeAN6jSsZ8JTgt7/Selq6wsfkChkYmqK/KuNt7KjW
a2HnPWb78HM5G/Sse/tvZKBl67naTjbGAXQK/5X9mTccT2cKE06pZsjPISR9fP2P
wTBTrYVXpeeRuGQZAA6SU7msUee5fXGcUgjaGkImLd4ZoiXcHTeOURYONnSrQNSd
iHipcb72MBguvnsFnYWoKSKF/aA4F74LMNiY5fY2OVv/iLC5IRsUW/cnnC718ta7
Xu0Ub9CzuJqsGDxZxfWScaSCP/I40MAfy8E52KJdv4iBZafyoAyYIOZrlq8xHXh8
2bxcjW6mdH+SoplxwW/zEp6ouWauHgaE02yAIlVntqchdcxhZSVRWboU/1p/ksSA
+NDf5d+AquowyZAFYTom6TG0z8CWyajc+pc8T/cQomxxZ3bZA7pKf+eAanKwOFgw
xdjLYVfjO/8yj7l/RfyauRfa2ferNqiXyIiOnLqAZ/Ewcmp7yHQR+G/7dHd4PZgU
dWxgFO+morR6qJqM+WObJLLY0l6801Q7Ngs11hSHWcknL95YVgd8nWz5e+2ByVpg
Ru9wkPCxT3z5QfcRMfVqWwx8HcKGfgHL2oSw5qJTbcudkOPqwH6P202T4webZ2ij
99TyBr2sSX0iW0GXC1GQxFJKdV5mDgTwnkkDNA+xYbP5+lRHQwEJzItvQ/wky/1g
Fe+VWk+PBTQmcL8GZLWJWBk/0k3ZlgNCeJaV+dlTjKm3bBZ74lw0jq4qYOnGc4f8
Vaya3KvAQvBRzthZtu1Kr+U2dsbbplfpiwtJtSRqoxmfbv6nelstH9fKDllIe5Po
mDGYjP/kts1Tpo+ZqpOvgcGGLtk2H7/K82yeX8khMsEzmOwPNCOKqhkWLjNRZ8sC
C9VHrN8V94/ZMjd4VDfcZwseIZr/+gzsQkyJuE0lGosvwxmH0Zdc3IBeOIb0gH5Y
J6lrzxjZ4pN0YfYo2a8SlahNzqclahnvOOsbqZd/XWS594vrG1r1mQf5PFCltZB4
63EjspP49faGOR99zZeOYwee9haa3u0oOyOwCS6dIMTq9+RSkw2Ob4JuAvnXT5xk
gvatGgTExm6Ly4LxAYJKS83BOuKZr3KKnEXwzYhGfUS9gKuce7QBj9mkcB5r+UOP
3dlBC6Bk08EA/K0zRFROHbgMR7GCjZtFJl2VF06yK748c0dI8biTiu3UA1w/U1qY
PP3cSRncZ9CALhqTreoJYx4587rFhDiiey6HHnE+I3oBGS+gNVNLELIeUbLEClX4
w02Ak0BKkhSu2MktGdSUJh5/faVX5I1j4GoJGCIYRv4NFLgwvJm0WDqk7cbrNO5z
TwwiA54CrJ/qnbL6xTyK6bkVvNXyKzCcofZ/4bNN398cvwXBsn7m+0OkJ4dsO2Tf
OiMDAOnvm0ABmgnUmpZdkuVcbXxzV2wuFmlz/DXbWZzpoEyDIVCgK9lukL38RyW4
X83J6ulFxLc6pTiyXag2Q5NPDpIniah6LLSnoAop+SV5SYcNweIz/FAQwGSOuaNU
fSFkGtnQlIsjoFvw+HxuWlqoiZDXXD2kh/0W6ip0f/6eCyTe1HJYnm4zmnT/820a
6aQFyxucUuUJWQQqeEjG3fuEX/SQqk/ExaYRoa8rMgLWaMuNY+yAUH9DZMt3EcZ7
PvOSi2EH8wSQKdN5Wctky9vwDrp/pjJCrjNpq0ebDxVuI6D85ODkcZK4apcEYqEv
WuX2AOBZJWJ24YfkoIhMJMvwtBqlbAdQ+NEGLX3jQhSm6QFwYX8Sq0bR9aCPB62O
dbzEYBU5DqVajrpijxsE9jtIe1y2vif7kGYmr07A/Z4wfK9SXdbsRm2kgL6zWINU
JZJA6dSk/HScr9tmhFSwFVz1dW9VQ1kk/ZW3gykExuMA0Qu5vp9m3wCXOGNcGE7C
Ug8G4Ccz1RQjBGduQ+qaFLt1uHJ0XWVld6M9sY6NoHG8M8IpyNpcBnwQzW/bg9SO
H1VcPqLTc8koZM777qNXys7J7fSgzdnYSbIFwnsk6/ie0bXGyNWI+ZCv+gudPIHG
RLVWttkHfS3gPNXf2EuWV6Y7QxvWEa/vIw0cfxYVRBuBS+H3HI3sfi0jj3lqfB3o
ab7cDfsb+j2R5cTMAvQQ7aC6lWdyrF45Hsc4AcN2kCsQM504EKm4k/CTy1plVWtp
Ny9Tn4Qw7Z2eA9+hCtwlQAWgOuBGvArPynsR1ZlvTZlVh+70l3mvFM7iofiXm838
H/ABWYpT52rLFs3ZANUCVtwI5pW5x3of8Xe5SUAUi1YAcOSx9IwUkTCYd1/1fug2
S9mJnMrTbqey9HoWZwZt+vVD6U76AwTXQZWpnIw5pf+xEX43Ciarn0Ovt+pZGsE+
bL5Shjs6lDEeNpg5FxME97R1aV9bCaulgV5wqaYF6D/ufyMe+MMRiq5NdbVA9Jex
5GoDBaDN9GAedZhibFEu/oWTNspis8kyZ1rAvMzfG+3BR8g5WwVtCVVFgtGOkwJj
oQ8jf8M1m5GQRGVe6+9R1+d7FLyzQSRu7z/l5Ph+Y77li9FzHp95nyhpqtXEkPot
yO/+ICNOsa+II5UpiaxqL0AiRhJBWgCPtuUKhO7MXdHeEJnMNCFuoKBY4KJ8/eYP
C9VV7398Oinmopub/kMNQ5HNDR2rUc3Nvp9FQQDFJZVxZDqLFcGKZblxiLTuHXjJ
WE/2su9EHMn+W0a+rNBbBq+WvYdcA3Cel1bTwI3G0fTDoxEUr7WpucFbJ+na2mvT
Sxb8f2Lqwn/xyN/9F3Fj1QBG4OWTq3KSmInspaur5QjVqfMTp5hsLkbL0uW8VHJ5
Omme/0LDAq7yCOmTMguKLzfcosN4NOzyG+qUmk9IEws+Hi9Biyfb40/xhp/Ds95g
IorUBD4JPShByEAM2jRTv69QhpCJWW2H7QfxW7F+HdIoy5xFFGmvfUF5THtcc2Ma
kGbmZfXLFLoceL69OUwnz5fonQh4EOjw3dJmZ+LBeFuP7dwwzuibzHoGHMYes86m
LLdVsajxaAli2mJetsNAReivu+C7tMk7nD/oMRQEtP6rOnkYlsGy+DhB5DQx7LtA
nAf2x648GXKYP0RmxJ0cqjrcoknlXjiArdgbqVvDluOXh8GSY4lMTBM5gmxDJ/4y
9UOlCpsQ1tEQ7iU7B5ds8dXqDEcUx1q+hKDG7BwjjEiitH63Eu2+dMxiLX2bx5YJ
i+9X5TQqU2lu2w78jr/cljTBdOGtV8C6jMrLwePJ3l1GGV5/mydoeuAHzbUiDNs6
a3buCEW9dKp5rt9VkrK2MNRp0Jgti+ajF2Vc4+HkxG63fVbFTQ5WFooaxTSqMd5t
+xDx/+DUP0+1KTF9vT+IGIkDk4Xf9wSeUNsxDxpmkhROHLSCoZPSoXETPGlkKKWA
6sGjFfS4oR3U7Dz/zG1zVOe3q84x/EHLSv0ZyJq9znzeo4qK1dzbz/V6RsFmM6Ls
FiRnJ4k0C0QqIbk/yZeBqyVZWf7hBbHhMzfz/FqrezMBjL+IgocemE8iHMmmDjsq
AEcYhgdGPBDGUOKWg+SrYF3vWL9DDRoWzYd5J19nFWOoTuvSxdeT0N0fHtiVLswM
W/JWHEDeeWgFhMGEgFM/5EHzYqv81HvRn7kSC/Sxn1DPyI28he7SRRs/hByOFaS9
s9mOjZTtNP6Gnhmi0mM9o2UsBOPMQfEtiWjUTXy5Ezn8JoGnsy/OSUo7v/Qd/nXf
YezUqPlF6GGGrQaOU9pqPSf1owjSjQabUFFCFUR4unwwJK/3LeoB6O0RBCLMorJ4
yG5j+UiIQp2vBv5k+dWM0yKprC5iEfiRL2bpARpr8G1hgt8KeaNIsIvDDsy/mUzC
ImQZMoAPVLG0eDS8z20lXkC1zxybu65JVcLJEWuFHTqkv0jcT7j2/b7/eQxecNdA
kNyH91NGhLUeRx5TRL2d86Z8c7xhFeT85b/DazTFai6wGRheGwrspjncLpRuTSQP
bTwE6zClcKT1c9zo0BzkmQ8vtHrLOeLeiHvj1n9GmvUzuWQRT7Ec9xedHXxm7v2L
svGDP1cUfW7Ywmp6AewhKxiXX7OooYFxQp0Vanx0kQOZ0ftqEhmNPc7a4MvkeOxz
VxC2E7/kcGC17pRMFntajrEEo0UhinFeqzY/4FGJnwloeMT9ODFP1qulbgA03Cs/
6ftoUQhDCJ6dhoqxxfZQorWZL6XuE/TcA6ESdpvVWMsk6H89LTKpAFeViSSwSfeB
CC61fcyBfZQl3Ag0fTj47VVQaVx3pa55rnpysGNQ9VlCE/cjS9qHZce1qn3TGnkA
cYqew7siQYYKnG2fpBKi7OLBEW5AQJsjvOOCMLrSy1mVDwa0cSyE7GrivtxtYYWv
ruQZdRuwAvKCK5ficLqfL7MkSNMjX6xLuQOfBB7hVqj8W6ZfYqveVg06Lo4WAqKI
CXuhQ9JfXUYe7pGAsgoGfeTymytxsta1wQvV/QT+GMiMusJ2V//qNofI8QddyNnv
XMvRlSxqeEvQpYsqU4iNBsqgSGtXyQ1LvdJilKlUAlOaoxSazFomIrONKplV7qgu
S/uwUpaospqq3bpFAPpDuWPplKJr97zKsMxEXg5+Sm61YOGeiKQbrKxR1PTQV1Il
jXXxxoTEsFDU8AP7pCyYRukhoHyZPYcG/EKV0214+62rIFcfJST1II0KtXKsZb6q
HGkWiCPCCMNHqpF2r3rSa9Q7Se5PrmiewhvA6UuIeE1P2L0O4MIzvNrQisnyZTIg
L+W+RdeRDJP0AE2eBs2dydT4AT9aGjFiDyPJr4C2mTMfnLTEZpKgrlWCUr9a/UDD
19hCb9oZ2eUhEMSeQdGDpHoQBgsgndmcaNdfjisUHOxpP3nuxVEhSxilpyfJ9uyQ
tfPL+n07rN9NCm9UTHdYPsJ+6EbSsxtv4tNJ//jQJtrVoBHnbRMw05QGAllUDgI5
Hznw75gG8gGLO7alSvghoR+TlTEtR+6qhOXSzd3TCHoklhPSf3UYLAK1X/BToDga
6mPilIE9efR0HRvbDKNzNWVo3qZXJmiNdMiXQSvtlQ0lKPqMb2mTULrPU16S2yFn
nOp7YqCh66yBuvK7XUg0xvasGvWi5KhbHr9k0+t8yZ168GgFYJu+OvdmFyDLCj0c
Fr9Mm6zwJd+EcrNSXPv7dZWXEvGH4vo/LE5vRYQlMLYLzf+oPuojZHOOc/8b7N3q
ZDRyO3EzqwDxL1EIz1PNanKNrE1T5X5xL6IDb+2Ck5m8DQMcDWTm6Zs6njz6aS46
nFSpPD22KD9pm1YwVXje4//MuR3lFITnf+PE1Q0UU0DAzzeDLvY3cFFmU6ZWItqf
RiSMg9gzdtJeU7x3w0FqvTKHRZncVHHf1M6ivehDoEFXz2cAIMqMn9fRhWnymNok
JsRmp+5n9NfsLJ2Et2rsfrwzWUZoFGnRk25TV278nL+rEhqQRi/5tVEQ+TlvVNhp
FQ0iNhkt872N/Si4u2agSWStuztw7n5VUnxTRAO+qt0IiRgPy5EdFE4dJwihplqs
GdWRw8RYtVA9l+1AsDlCzcw773HD6F/S5cX6pNjB7Plv7lQp5IWfWfj3JxI+6JB0
QfyJ3m4COWfaM7PgYuWy4pAPCtZH66SlWHqkfSGv00ZHLPJ1mnxtPsOxeePwNL5w
TONsUC3D3ffBqmqTD+yBj0llZ5fnMrqrlT9biGqrrfpdD7D3v5DUacriP5lH0R3g
Ihs/wvR5tvZv1isgn0DsWWOSZi1MaYzpexkrimukY028X0H5CQp4p8I4QfTeyusj
b3HEYehm6OuVbtL5+cn2P5VF8csAmmkRdOXra+tgu7wFjTxI5vwaK4nhgAkeZJt0
TOr1ToUfIFUOMrCH++2NG30v85exHfaA/ZbAkYI5wFfqWiz8ByZoHyX2J54cuMuK
Gt8g1jmTtT7eCT/e0zJXGLgKFg7tyCo/qBaALLQ22nnMDTAOl/DPhdZBsEsswKH3
fTSgvrAvEdsBmkWHQjtpqx4VCzqZkl6+Ci1JIVehCIGYNz1sumfOzx+yU8xaO2WC
wqXzwZqEr6Ai+baPYAnJnl3iv8iDgGukab/jUS/Heu6rMA8YgkDp0xzSA6bUR+hb
bGo+gxLhbZUN7WhACmulLj1fICxZN6GbZqtr2jSZkHbvzsUNMXnfjg8YqR2sic8H
Xi+ll28mQFXZxvNbOuErx00j9vYiniTxDjpC1wL6G6u7+tcRQi+bQIasWNAyNLx7
hHbsIIjWxCjYqVJZk1Fg9THi9bzaRbLfkqwdnB43mosEhktBSXz3SHBH5Spmtgjv
fvsyuRVkpZidsukM3i8s+SjHq20ygLAEaqcCxA81TKrj6OAfPuRYQMIlvYvS96CS
XYUlCeFUUF4cwQMkhmx6RTWvlkYB0a9EcLDDsfq9csyQ27MuUDRKi0T0dFS8Cmfr
cAOKqOGKXadmLpGgbdjJWjOPc7prBa6n/xvCktL7kj29UbcPZmmIpTK7bpVaMG4U
tAFaSsYMAIILFVKIeDxxQ4SFZA3aW5bkok3VeqbcxPJtXMrBaaXnMaCNYUkDDc93
tHqFDovklPPEz4iQ/V0gdsqxbNmYYDgdCfFaDSsCOn9i2WuhiOTFr1kX05whfMhf
pfyt34CdG+4shMBh3Xb9bEO0G/9l7oSP9tUk1t8Naz8SaBgYKqEtL88e9PeGEJex
XtK8wAjKSwtJmvCCETCwh8MKhGOowm+BtsSVIswwg5H5/b4uR2az3fNHAu27HJXD
TlOuc3fWLSjsLX+JzAeknipp0d80CO0gP3lz4qRWJELGR/PakPXb5OMr39AIhCeJ
zbQTwW0UFamE0MIUkEnSKjsYPiR2J0Ji5kLIsawpimvbNmZgcER7MkvkA7QZVTpE
lBTSb+wOh7YGO/K/1zYtaO8QdHvpX6+jzHCMJfdi75SpjbtfACoz30/1UjSSSFfy
VTCpstzebk0O+tU6gA+Aqtm9TyhxRLitcg2wmeBSm+Utr1skBREveUThFqMgWTYO
txAx3G6eMx5Gui8JGuzHimuR5jr4BUKxWWHGzR2OxvbRKkOyNk3x1u3hW438Lff5
Ku3IISgkyWR0YM04z7fy0gJOI/HD5gc5gl0pUT/dctKOEtnaVocDLuc4ACvHIYiH
Ee8x+qT589QDHDZONIbQsiVJKI+ldb6OBhk9lLh4kdTvYipxSYg5j+IcQkHpVW0o
8UohWUMVC6hzx3STUkX8oT80p+oMizoec8t6EcBkH10W/huknYYsLKtRnUix9N4Q
GBFcKmYj7cBujP4n/xtvASBJqUFeWqi6Derjnk+MY1Cdds5JD7r1xZNIXTGrwxj6
ZkkCZZc7ZXmVFEU4oqudLORumwOFXgy3wqCQQkOkx7HlJN0zvZw6JWNy873QxhB1
AUfi5XqXypOBQHvbFmw71sQTJ+nDV0/GkTZtqJLuQjhOE86DA0aW/92C0aRW+F2/
jcmnDYvLEEG3skfcAmUUGmrVZXcBs4dSKz1VgPjm3hp8er+Fia2/JN+L97kXX3dV
Fkltjzwz1+hjDERYK77I5YEgMH8gUaVnIw6xwAfczxJKtgnkXmRA683qg9k/OczH
FyCJ3wWAwIifAC5XcOY3E3G4ToKtXk3mjEAmr8cvlCz67L1teuqSVHJQX5S1FPRn
Yn5yzkbdSydlbggjtfDVhy+0XWuy85YcUOE7q5AsQfByo+/hH8umTfoUpl3Se9nk
hZ5lONMCJsmUON3lcM+t+YbJPXTltCchQz1HzoOGEuPSUwifxwvafI6eQzwAXe6l
nTUgDUUyWQSF8NZx0VoH028TECzcpRx1W4IwES5GXdeApPU+Xs9TxE/48zS9ZAZh
Ilkh8bCKSXC0lGJnmgo70OG/igtRkSSV5M1DKCcBVKX+bsS1bauYK8qWBxOjzgaq
CPfAVfzeOB7mdztHJ9SXolWqDACILwzA6CdOub2VLTXT1reQBmgk0bbB/fe5V31J
r1XiMh4X9LBkhoL8LKJ4YNaWeN/Nuwmf2Mhz3Et6/vNZW8ezE+l9y8Asn7INKrIP
JB7zBD8Xj5gfLu6L8HM0vc75U6+uwVu33vm42oD7tl7H6gcIvaXudKIWRI29RRVC
/eS1nX0NDSwD0k/HfP66iATNBFex9VeiZszZqIOBQ3K8eVYKSbnyZ5KT1PSiTvYO
U8mKKreW2OO670TNELNyKTTTTDvOPHrWO95JrxaBaNSYGFGUrbe7CW6NhsUQy3B0
X/PumdcBFRcMojLQph0KbHyINiUuL3LiKo6PyGYMQJKVxQPN609ve3Svgmn0j7cW
+ZMAhB4mrS4GOICvOOWgKqUhwPi99+MzxGPgM0n88NTguoT5UZJV+2pWEnwH2Vyo
nCfRmXYMtFf7sKQoMhgF/psf5qubzbwEonaofCks8QeORVUqX5MLNJPf/f+ESJtc
WVRTzrg8wA3sPuCrH9JNmemqrZCKgmZZAtkOz8/BVFiSashi2lTc9oUGFCYXTvIP
CN4OpcD1O/zOp+Hy3FmcLRetTes+W8pLmHQuf6CNfUIXoHiYnaOf0FDG5DO88/Rc
BfdEY4prUqxdCm+yHSCpnAApbCEbrrSLlGgF8h4C/cTYijsWreoMiFZZdBxxMvbM
q1hTBAvbvKenWPhda8qu8cIXUvx9517AjCJA1asaFLJFGdBi8lGjaxA3xsJsI/Ju
gsFoUEmYEfY6xCWlv4Wq5ZwKqyaIFOHM+9xHNO+6Ks6U4otFZ2M90gpHHdLhzNJ9
hOPZ6jMVRChv53eyCCt9L9a8H1vJAG3GZ63KYjFaxz5Nh1VqpQ1rexOE/Q867P7T
UBEncxbVZGLJTBmgdMx+45XVjAWj2HhXhy0WXgPjFUOusAzcRxoYVk8iAQe0Q663
TA+XTlUkGRbcDqgN/Wz8oQz3mecGr78trytpTw60WSd5lYUMCqZ0U9WTuWJQK0L5
oQ2SUd5Aidh7N/SjiI5gOB8iznQDqyDf9cjehV9IT4AwVOQc8e+xh5eHE1m5/vsr
zj61ksrx8udkdL88ffHYZCBhO4ALiF5A5WjmQkWuNXz1hEIcO8KyEeSgf2KeNxeb
CRyYnQQwqn3p7Fz6nAzQCKF0wsNHQAFaywt0ZyanKG5AOv+ZMjPT450H/c6BHJni
4ZaKpMI6+N419qjnDx3ZqFMiUk8VQaPR65P+JKUZEmVgb1DpWBkRzr6JiZjIhF5C
+ftKpnHf3V7ztRoJakMh5csRCUFYm6oJirLZ4m5ThY2nW2nKZOnAUniUFWfARtrg
BQPMzS13dralatZrFqgcErRmhwap0Dl3B2pU+eCVR6yvnErN5q8Rd49YHKh1wjqw
HvWI71akayE41tOSuJ5Kg8YQH1XTHjS1j5vuc49ycGQUyzEH+S5alg5JG81H7h8c
enEU4kjdGnpR3LA4gbYsPib23NQ1x+X7TJrDqiy2B6x6h66zhxXX+Y2QBtku/6Io
i85CF8Z/08C7+Fn8DlME3pSo/glpJWcWflaH+k1RbEYl4N8YwmEz0htdFBgStKtr
qcede3K8ENJLYw+9lEYun+tMipXejGec2mQyy5ev5FLfXwR/g6LkPl+n3nLzGnH/
m7RZMWHJ05omFJh3CN02sW4bMgVaazWumKeEqoTp2w0xUPw1UaPM87CELs4Ld+/i
ISW9YoGLH3GlUBexlb5nLNAstMjOM5O+TWe3Vp+hDMv8b2bCHbduCmsO6pC1E2He
mJvutQBWY49vHYjHEFtCXPlexUZy93NKidfEj3+ZN7KH5KtV/hBn+U1X+cmzWC84
L8+5ulGs5+bzO+IIb2pevRNS2+RTpeqeebf2TU3xviF6ZUOaI+sEwaFcbQAe1aqT
AvqelGFz1a6jAQfRBzGPsi7sTRAVjRzXZPpwOMXuAyB3yHNG9b2r+kFe7QEmMJWl
Ns2z+jBUGy+bOMLt0mSSIkh66qRvK+OGGxW6I6rjBkIiTGWoRXOmjqfVwUfOWsaA
nsb7rL9hkXKJFQ+Cp9eR35L9Jn4duKHjATRZHTG4BW410OVfQZI9K0hiqOhU3Lst
KJUH7rGpvgjtwU2+ha/qJ21OfAkIrPHJRJYbxFmdVGNiuUQhjytTQrM+u6L68ry1
4xGYYAr8JOr3PUxew/tvfv083P2csP14kDgXxlhtC3XQGt/pdLYTYsWBhdFvtbGo
djA+kJFFgtfu4EXgJVIiGUWPRepcHhMITzyA9tsSjnwuT3R3t4CjB9PL5IpP8QIV
/wrhdCn1NnB8K8N+0w2Of75GNEUUmyf8dbyVy8ITcnEzBICo9wLICFR9okeVS746
0+20PFfHDP4sSGt5UKGKRLHzRBvmeqk6fBd2vbXtQ4+fJ5NCGra+WJqFOTLH7iu1
zEgZQro3RN5uIMD9RLJwkiIvrpa2vnAbY+u1IdmJ0/gS3b3BB8UaNNMCUy670UUf
T40JSJWF4aHAqaNCxhrQbJuvSN2R+ipfVFBkHJyzhoVhPblQ6OF+zfZPXOEvICky
sQB44A7LBNexyJuThw7KSI5+kOsy1wrZIPBRmSTnWLHaNzn3vB+tjW7NX5lENLb+
XvHBvPSr3PiB8aiSFoii211OXs3RHk+Fmq/lyMlk3m7hlWoQLLnTdz99AVqkqMCO
T67kDFLPrb30n7J0AFWBTdW0XOOv3yg7mWU3ZUllqzHpUOZcU/j+g9+H0OXz3OwR
bJ7FMydFVNodG0aWLMfs/2H7KcD6zuwMkFVuhUx9dioq8Jbl3777DSyclG6GKNfr
7tzBXXCzPuhZlFst1vDzk4sSOaXDRCfur9ddWTybBEtY9tTuNDx/V8ALXB6BfHDh
t+jL3Xc7bv5ZN4clWyYSrbVeNWoAjkNndX++bhhhGgnjQHLnQcaEZZkFLK6d+EUm
eezqV6MztQHazLp5lGpYfNNTDEk1bLttsv4g9ecZIjS5IqsS1vBYGmI7vNm7+6d2
jZy/kuFE9CLc/E6ni/io3LbwZT4bxyPSb2zFgvTMeM7SX2DzDvSkl0arqow20qYv
Zt3RaY359LxmDoFGRB3aNlnBWZLln7xhnQTzPE4hrEXIa9kDD5bMyTwTsl2295Mw
9RFI7nSmtvisG5Ghyk68JUFRW5MNooTFO3DJ/2lDWf2ke+jkpXaR3uw6Sf9HoGv3
3b3Q37yAH+zmnz4sF/GO7VCF2ExUYEwFsK+DK2cJaOGwJoYL790inf34hf5zW5RG
1/n7yuGs0Z6pszFJJRTk2Re2TxW0XMdHjdZd/lgoyn9r/WDaborMORbf84rrwqhU
vwfXnXJiQMimBnepc993fuf+gn7nClWCyPOPZhCTGOEdyh3O5E1n8T/x819UsHnE
lmHQVCLcAMU/R0Whtn4u7pek5+xjZUyKLrA6pYkFr2bkryieDzzFmeAoJ97rlv2l
cTMxSR7BioBrdMwVsZs0sI3+4t6TuSn8pHU5G4uZHQ1Ba/XxJ7oPgyTiDQHpN90+
UKE5LCjRjp7HAWn2MojdvX94NOHMyg+V1emXKqKDFec+mw1R8nxhwTkzcFwR/aEr
P4XQkklXbj83P7LJfJFTk6/nc8xoyVC4AzJKlRaKTUdkBM80wYFRrCH/2pbOk/0f
NmHpkRQuO1k8BAky5WfCaSlUZ4O10PWiuGo24762Erx/rBlFTS2lv+R8a5qHZ24+
SMk0bL73s9THYcjMgt9pf329HfkzcaR/XQAdhZHPwtWpRHvR4c2F9Ix+4YrGOQ1s
QyXhiVMApFR4mUS1IUKailCt9bV4k57Ei1lJjFhiziV18waC8qnQz9w2VbgUw9FG
3Z/7flXSwRoJ8jyFmZAe68YGK5j+NGCRHQjGDtfT7spDepcFdxYFMuyFTtSn1QX4
ef68KR2oKA4MgEwxF65QWNnMYZjWZC6FlsRIV+LMe4b1vRVtc2PvXu6RRKf31KrB
XXMw7YrfHOVLwjIKteh3JOnd//WxBUSv/159kiwlACMKQ4a2KnKgWLf0S5oMDuLZ
zHziWLGX5CEjB4f8Qmcj8IS6ftpWHsw2yhQxyNlmA86aD14BYolamsgw38l6ze4f
mI4wMzFxRaATy0uJ0VUNJFKmm7R4gvP+XAptRVzoifhHDlwcWd1u0bnX6eK0ScvG
+O5v2gaHY/N/gfRZBLa8doPJGmO4Z0JwqJulq2rFQIhHjP6XUVBcWd1qbfanVOyP
uFoBQrwOAk9qPF+62CAdyadwDd0bJNWMQeFlWFQ7HSMxSrIwFYUdCjtFU+oyFhXU
HAD9cwmEHa+bR8Jv3fSDFWfs69yLhteXSRsrdKiG4r7FUDhxztbbFjKRyCr7IjEQ
Y6KEaMi6JXErFVd7THfqjV6ked2Fvl0VbmviGikzK1Yese8/JW0UmVWfRft9UhK/
br8FQkEzkfch6ZrzAaIVH8uDIZ+wzHaGs5v4qe7uczh1gGjOacVvygfa9Zgom2sa
SzPbxFi2V1uebn4qSW/7dNojHppkO+4APXZHJqVY5QGEaifecQlKBcLECNZYvN7D
bydXzdbHpchrC/VRnGKKF8Cbl4OUbsIAYa5Y5K35b0Bz/91YySHB0zsiGawfMoqR
rwGNtF8ybBAwyhWWBLyZghyT/O7yfaTmNeMmwMBPnz3tuHRmxnwnVjeUNNbwe+P+
kI3nU9CKZPk6vWaAsvPpQyiAUNmNhHfMiNOAwBDtkgvoaR7B2YcOCZ0FhbKmsOBW
DETwYbKcjT2aBTmscg2Sc0BWoQYzkFXyfJaYXL4OF96j5EneBjzzrqEl4JEI0urw
2RGY1uEfZ7FyEvgInusDHCV6tXMJe7DNPKd2gCU/e0ULPwpoo3DxZ/3YC3806lvP
Xf4tzMeXnDTO3xd4rf9Nvhh6HsgE6KZ/Y8SHuPQ289wwsygcLjhvSmygM0dQXnt4
jcO7V0vc3+gfmKZeHyzbzEBRQhssA3gr6XXkYwe1PlwnUWBV/5MpO/SntEAr6k2B
DSlOu6UHMEThRcwM7SZ4nSSo6+MYAqnVhpTedUE3GTJU8g2xyav75ELLGASCG28B
XoumtRIw+KmXYw5c1D6jaeJnBbfQ7SyYIkWJZ2Co34OEOBNcHkgiOXiscKy0GhYM
E7oRp3xnt5F0LvkioHNoMruv46HU3OFubWt4tkMuYc2EiY08VikL/rrwDT534sWF
mwh8GIwnyiWI/1kjvVyNy/GBAHNUczuzFZMr1EOJKg37I/sU7MB8/oiAiwhJWxYU
BGULG9Mmyl/6CnCKXxU1tpmTKOyaAoBq4K3xb2w+rpa0AQiFk9mrvfDd+F/wPDL3
gnjXjZap/HWdBOFpS04PLl/rcE/1kVOJEktdzwe45jIkdwFmw5YeMErRmBPkhQoL
CegnXN1XlQtob652Grd6qO6LyMSiFhNosRS3i5nl8DgsH/2pe1rQgm3nWRxkpoc9
hgxH56cNw5/UPKxe8AwhfkB6vz2WfeasPXTH9bOzYS1vB0ttmx8uK/uoZkMFJhN6
h5jFiB5MIl6mjqJLOITC8am61/QC5joZT5+DYurouvixRy+UAw5aC0oQLzD1QrBu
1viELfD46BingoqVUArbMng0qNV9Kr1sRa5VLGRUM4eiOeYJY3HI9lNVgC4LnEEw
497ZikPujBlJaEqetNSntNZeb/4P12bt7JO9Jy8DuN5Y6weoVujXQIiUzwqE1AWY
uGrXtWdNq6h+jyGQkSA47jU5YSvSV+cGjoLbghBQjnbwctxkz1xITh9lfUuPHG2i
avF9hcxV6xnF+dfneoq9l4UE7Y/UhEVgtUwzGyqdr4d71IplodnIU/qLG3eduHiN
ar+QLP8gBHqmY5pVMj9KjqIis6EjCYKIgN/gT/ypeJKn5mfb8Mbl5XoqMkZpv9jd
CInEfLAZLzQWq1ZCHgLA+NO3tan2UDAxtxfDTfplCozCEn3kymnrZVtKFwnmiHHn
SiStBe4974wVeAn3NUJmOWHPLSKqPCy5w7bpJ93hOfphcZDdxOkPP8WdggfE1yx1
ldOh6t9aoqCRcowhAM7i9poIO8smFyHbG2LztdHZYtoOdVV/7EsWW/PltLsRGYSj
umqwFML4PBwxrLCiJ3yWHnLlAnZDCYgWq+hFjrsGtFxwhImlNRFt0t+82iuI8Ufh
EuRnfs58TA5dOHFpx61I99kbYEMk155p2o8go4OWR2sL0yJjhjhhM2614at/gOE7
q1Karh5+8X8plpKg6MqLtMjIQAsXMvrKK3XeQFcgYgYD12nqAAmnJ3x2LJYfTCjp
VLwCcHvn7KcYIonlHGOaHhl/UfD0/JzH9IGQBXWWsnuQr9gQ2CZGWG5ZCBJyiWgF
p8phsgOgUPQ07P0X3yYjbPcgBz8kNYR4F6DBVbc8MDXXAyVhBnNoJKqyUy/FI9dK
xHPrALBuKTB7JY39GYtVgWuVFW9U/xM9GTjZc7JkSCYWDEiTTSRE0OdiYaG0kops
MbxWvBsR4+I55Hjz12RgYpJ5Vyg5hX9uryxv0QxX939iF/ZfFGM4HSH8owxjwVgu
IDgrGLlq2nbVD8o+PdwWQ3/8FqzHc0V1cLfe+VcLRir7p2wkKWqm2fxFXeha6q20
z2dnvTOF7uTvQrk02X3Agt9CsAouShDR/nFDLcFU1PFZJBS4zm05s7Tl6xuLyxks
FYVw/mfhsilkP8t4Mvp64mOrO8vFSd2HeE48XeJ6bQ0+5rZHbYakgROFtPe658KT
Ho0j8SthEnZ/NNaW0QXqXsv3eX/gw0lgb3XADySV+VnMEGyeXAXjCNRMMFtuqU2F
kWJmkimKKQtw6gKSl/V5AknRrnDhQjJgf/OaWxsNYvgbIUW4DgV775xCEhH0UXBI
jgJdO32OMXF8c82L8QhXpVmRJeVJLaKHt9SeVMNwf8ZQatAUCSbfroh2XVE8r51J
hNa71TdkLo9BrkdGksp/8xTRnoL/uP/OK4V7F816KlkYBsxN5zNBVIokohijpNVM
vVkwu97lCdeptcACKZT/Dxhvm3sPckUwQUSb8WqVKtDYIFrJdYEG+i8p22K04we6
evc85s+w9S3PowheUeRkL4js1QRtlC0hKPsbe7mjP64KxvERk8YvpyeF8gmfzsiN
wD7fyRqKyaaxbB//kds9GaUP+3uTlmrxixBqBTvH2KyUnFXOeP3QN2t0UwNud9ML
PzaxC7Qt3AqSrcZnCIdPE+5Xq/9nflo4z/INvnp3FmkhKDk14JGLkgmp0rItpSYx
uZ3hkdxb9Yfqmd9i/DrKXL8CfcvWqrllaKpvJbQqL/rahwnyTPC9nXxdHgg9sMXw
4v1bfjmthih6ttaonn18+FB4XSL7Fo5djwX0Ut5kymG5A0OzP4cQkvYSWtYJ84Ch
P3g8uAqtzk9Teb/tx8o2vyJjY3NP2yY4BHI0WMt4kHyUSBQ7YMAf0AQB3gesp7lp
n3CutVqbEMH4M+3zOSd+nqap3NlCQBe26lcEU7hofZgV7w/dFWN7r9VECaB59mOY
ybpEv4ThmNIjHqAitaiHKFp7LrqZ3gjBdYLMrJFOaXZ5xxNGL6sPA0IyZ1XsEJTV
qXadbC3QinxcfB31JG3T0Sfp8RaLCyzC1Y3UQVSAEc+3sdxNwgYQxsb6s9/ESd4o
8BUpZjjOy/Fr6wqcyZtcXk+gVFpyYbDC+pLNYZlfioq64/f8YVu8aijqfHalqjqc
rBbaD0P/tQUIS8c0CCVsjK6LgWU/hhHPIJz2nUCEzQyMpoSgtkO7Sl28eFKzQhut
14SguV8SqXHd7DELCfkbZss/l/7xCZDlFqIUkrszfsRAy7tgooHsUBgyT6rAGs23
hLfakHxGr9iT3JjfD2amDGreq6/3S5We1MoZDbXocZkopMn2KOjFPWDjC0bau0Zt
ESguQWGKu/k9pDLkGWuzezBY8Vw6/eFroV1Kgvu16gOK2gHKtjWvwGFtZhfOC+wt
+NGFZJRKbkcD5H2h3osUB6SzyeztDOnl41uPXDmgitI1f+Cj5ZLGahVDWWRnGvSR
cigRyiqPUJf+PZ13LbuH7PHjhNHBfhT2Al/pPJbAEdKA/ktH/KXzVonv4W/0aOK7
E8t3J60BuLhkr8uzTh/1L1KCt+aLMAxHL5nbfaXbVL2MhoSYt/lPQbhBeMeGyoLS
7IQxC33MGPewjwk/VxbLVnXmkNuX6aZKVA/PCGI7xK9zQ5hF+UWITD25LKcZ2hxK
jo0y65R3pFyor0aDF9FkJJhkRKA6N8qdK7dh/TBa/7h/7HldYSqYDCl9XmoQrVlQ
wfRxldwCOvhlOUxCcbOmdY+LgPlQfySzcxiJ6sQooDk5w7lOT/DJKTUWll/vHiU+
AJH0KR0I9i8qgPRE41dM6JbKotjDSaOG/9scVcVGmJ8LWRaksiaMELQuz4Rao3yw
OoL0wpRfSn1fYR2kIj0EZCzhaOoZtQ7on9tSq7B0kSyS8Nl5TMfKLINHZ1VPn7/P
UIkXo4V9uUnX9kcYxPOC0k1H8Q8DxGK9W11vklxQNvMhs+Oyi8lW0L+jMDq7jDU8
i2fP2KsvOOAsRHwcEPde08fZGewXS/ejJyY3nQ9qQQpeyp8vJ+PYJ2w0FNdjt3lY
GVZPskPlf7y2QRp4WHx42+rCHGOpVWZVhswbmq145Mth8za1nACGX88393sDvcTV
opF1c9UImGIbsMqZ0IdoeE6UAByatPv4VMSQ9MraUmhr+7h8EEK0N6Jc5qthFs9D
6+0gXHbO1jAzdybpiqfLxaveeJ2LxPofizUTLBg/hqTA9NyCk8L5spYC8nvFPKq6
P7lW7J5hhcyEf56DOTZ4IdPIA17OI4r+junvVbsfkh40xkoEqijxkCgsO+KEsBBy
szlebz4ty9GunQde6jWY2B1flUW6PAKGqxxE9cYT0S8mCkfHIzIooDEPph/X5JP8
Khw82B3maQLo+cGmWr77BUsFW5CEr7S/HlYDWRaYaCnOZEXfvOynqdAUpJTHuAP/
CkxfN1RLC20Q829LkG6I4zWcba2+yJq0Rh72B4xV7GBVpie2z1ehsMTeHAHWh1h6
h2g2F+niirgCWZ5nC+OOUuXj53pxnRDxOVBirJ3QqL1/Z5jlO+CDATt1Txz47WDQ
0OZYUgY8MCr1gI/2JEj4ZC9Ynzbh8LXJzSasuzRe+Gh5+HMWHbd7NDy8b3gJWsao
vASGHAQh6mPmurx0lhGw8PqeIlCBWrTC5KsGw5rqCOTRdn81t0K6NKuRLvhVqoVu
tOs/AzyOAsjloNmPUqLj3epiRFBsY2q0ZmLKNdxqDrS/fmOPq5CjkcOIaCkWHrkO
H+l9b6yoQAKB0uEyPGxTJkKJ2IQM2ey5AXQugCxW/XPd/DEZCXQAWGXt5YEhQN5X
G6TAKWPY4hJHGL5H27O6h2vigb4DAF19CmdQq5h+KzwvPIxCHAcerMynAMD6wK15
is8CG71fv86i3nePpRBPyaixcLEqoTvvdqXvqJOQ9Pd1M1t4zfBKuyE1Qma9lypP
CTeJefogRORAT86k2uTMZF1rGbIskJz0/8LWMg3kWg3IuQdoS+ONqi9f38qSjfaH
2dbWjJZYIlukIUD1pi6KYBPkH0mnEYa26h2zvp3d0ujg2qy/m4J2m++HDggVGKqj
z3lgATdLudYlBvfEIaIFwi3j4ZKu00m5Db5Fy9jA7HJWQM5P9C55mhHCLxll2GCq
b1NLmbrTygpkmfIcUE4tTFNIw1yUOMi577OIwvFn0capVwwrioS2Hf3ARkooZw0K
deAESiHa8H5bNePsK1aR4j6SY+uD+8vK/z9UMDpMLWZneywCMqkA/ylnSJOmNgoD
PRN6JUY6sx3iKxabsBJ+xxt6xQsVAXasY7w2z3PqrOQ2dc9MpN4HMbz4qsaZDbt1
CohQ/bLnepyV7MyP53fG3lbGqJFCqFDViDv/L9QNd/isSD9lkg8uDJrv04VEmHzM
RBfSXCAYAK08W90Ec4HTCWnFGQL0iem6UUSU/DhNvO3e+C87XfU2k9r98JiV0ly4
vsvUDnmVZekcmE4kycrkLbBTCbe18aO6PIl8CN4pcyyO9D5wthO2Z4HrPoeOXjqh
pOnE56QuvXA6atZCF/MdAz6ghQQhcsQw/PfimC9XT4vLSnGOuDDlvjBiojnV5nom
HuARmLRCxjbtFGV6m4yEIpNuC1hAjvJN+TrYhOSRd6nHVJtNWGlQDqsRkXAbW1Mj
/T268l0rzW8u+AoyKQFbLH051WtiC/PmA+768RcwbynchOhGJgA4vJkopCTgU7fV
xgJqWww48PFrer1Sx8UcMxJrhI6dAZf8nZdiQ238BcDeah1C3DxN7miJ5gW9N7gY
qb8FTTRJcvJtdZZXxaOexAK81Mt2hPq3r/5EvXWhKHvYWOliyfD+6Pdr0lcZk4xk
h6gmRmnnzkYLcHfRCLxuRwT039BI57Ra6IP0SoNghxdTygN54FM2d9cP0mc8hQKY
Jw/RK7YMCc5tYYiaJbrHhXVfed2zRetz7D0wsRDWmLGa425xs0FghK7IlwBnmAOQ
bnjG7CQX5zMsqVqZxwFnBlUa1DKU2jbZAi1sJ3+Ilf36edNen2sxC2rf6lzQB9vG
MTAnbKqHjloXZbnf8y3atxqvtP3lD3E440trulPtB6dHnL8ZZz6CqIkrvt81snb/
p7Fru6HqKnygGAogY+fuCdbjyxrIUXgSVm0T8jyWUn4L8XbeoE53WIR4MsrC6KuV
Y03NdIqT0+E9+5sknoUKdZ8LMZtr3KfEECM2M3hqokErNXW0sfWa+ptfJSZcLjqy
tAbxryFOoJ6zZ8Adj3rjx6YITZAvawuAKlq7YpftInrApvfNUpgBLbIxmAqEvLJs
FNa33NFNC87ex+e0ETlUNI8gXtXAfcGFfMEGgo8U3rNRz4WwRvLf4Oi0seZPPKVi
wGRvDhAR29dfNcg2+e0ORGJDfaD2Wvl1f0DSORyYMNXCJa8Gu4L1fKLinHSYw3TB
u2QXJLNK5Hdp20CC6jI0/EHdIbizMqC2e1yBlavksilSpKzsSe3QAEigp59I0iHG
DsC6f4uPnMm5LB0GOfWNf5PqbreKzCVJrtd0ZNyj0Mn8FSH69R/m22J5xBjAFNAR
stF7PaK/LDqaTkhoZDv7n6oS39ZvZMbHlmLGvda4QhmbV2u4LLrSDL9NfDtZq35r
exB0PEvRu6iR3mhOVrejOY6gxqDuiispBODv54iWaSU5TSzKs0ijRwNzqMs86rhN
50wFmlTgl1PW+ztJJE0vz4OIZqNAEpxBU/bW1lFDgsXTc4XFE8ISBIJ8DSipPVY6
aWvA5bi0AipFsCpYad119hB5eSYPOoClKnszzubSX0tPI7nY64xX/66A/q4cgln5
hiBy6WOZy6MV2PqH2gW6WRqqDq0shD0Eh6/liAggtT1UROdU/zaU9LrmbWWfi9j9
5IKojgJ8P5hS5tMCqk6VStaJenC/pAmUBXdhqh3M8IllMOOa756lqGq7L+WWn/lZ
mK2+4oEuAHCH09ZlAFhDjOev/od8l5jbB03AV2AsZmR4g8VL5+HEkUKO7Q5ZuX2c
im0QqWOCJR1yBr81Xgp/pjDt8G45H0xAYNQOIJ96mbo/G3Htmha9qpJPgR98OTw4
mNF2Tz2f4VeiZ+LxY5+CXXm4VohBN++P8DbtmtcVHkTlJYTM+wJWNjp1SEVVDLcQ
sRttBgdlB9PsKh/TSX1FyvMmSYTUQTwuy+7Tk+uBWA0kK3vWBV0z8Fm8lmz9XeKl
xqxUWGO/u7f4VZdLalM/H35mpciiQ7w9btZL09XKW9v10/vi7qnZt+Frn6Avthxd
3c4izONSDLjkdWR/thYlx10svJRBggD9OS22Ie/APJdHOZ+gxmLwP6NNdvsMfBd0
ZnvHkMFsEBufffeD4zcSwDCCkh+JMpN3jhCA+OUjas8Csb+DikhGI3E/tkE83FWF
yiqU6hhyIg2MT9s299tILO911DnowNIN+nSVBH7Fchblb3YEI5Sv5ykhCFr5z9KV
QDMLRT4tNtsft+esRFwzPZ2XZaRLftvG6FoZulOZfcGo52z6tZb3YYNDYNzHsBOe
Da5CsSpr02On23ztPYJGHaOaDbA4MGp58sgEtxNwoXPfbEgFeq7YEfN3YqARq/Mt
AqhBDDQtMChf5J186CHwqT8kySZaYjjOHcovIWv8Uwpi6yE3jFObLldx/ApsEg2d
EdUf6o//nOYqgRIpa4zuaE0tXUhPLvzBtQXirUmUiR536MWf0vSUiBvS6kGZCQQq
atfi/e9Son8AQfrPF5arwgIiIiNCMaGwfYj+cw73ofCjbdGSppPBZQAGxXfKnbd0
LldBLMujzlQk9HFSds54fszXM5Egv5SudJ7JLipTgcVkJN305+RWB5oi1ReOCYAL
hhL9kHKjMXir2E15Lkcfuso05ZlrWWB7pVOg6YoP6ozLUrWDGJl80OmNBtFejmjZ
M4JDZhOGaCGMFGoef4BCZDQLGqlnxQrMoJ7K6FUWqFK47i84yq1K3iNK4ko7qa0U
Yv7YTFGuEl1DoTIzrbKdwH293zhYe3hF+UOIGubap5f6dIZtjeBE3c8IvgD8t8Y7
wKvfh9W0p2hStKQ+55XHXIEAOQVPDsGSv5MpPsBlYRruoxHn0uPX09X3PPzz46ld
r+JW/ziwMixgHGeTg5dQo7v7wWXNEm330WL67giFH9H7BU7rs+AII9gGVceIxb3M
W5/36ft5nwP1t9qQKUfC5vorDT4WKm+yGSLx9f4yESE4BuT/Hux1JyU0V/hKT7Ww
KTkh4m/+Guawxg7+DQVAgo7R1jkmx+3KKgqJEtQy/C0NBsyCZKBvzBUuJQGgmJpc
55mUAHEb/YIkZEHkF1JSXfEkwwXs3ah/wm6tO0/eUlvj8oPkaYkjUWkhamtgKU8w
axiYZADcZPcViPTSU1kkvbGyaEBJHHt9LwBXH9H06DuSewv/cZApRBC08V59tuq9
FJNQ4emwOy1ETmJDKSego85s1ribPuEY0nvt1F7qe9ykvukurW3CPHSlQaQNI8yM
BaQsDiSC2WkGabBnhqsoSg6hOFz6/dII4VZf4MEndESzc8FQcDJxO1U6il65Urmg
78VzccQKxNgiMypcEH/BjqugOW7Hv4jFZV1mN1bfQ1tXUYtAqACHUsTvfLPzN37a
J/qCk5MHB9TNcslJeSpjevaF/GXz1N9z2Xyq9TcH36BOS0cmnp7MlHCkjQLlc6Wm
+mMzcxQQFDiIhLCfKtAmQNmVC75nNumYttaFRswIJmbrfExU/24JZvU4EQhc/d/k
+k4fTeYzAyabNC/xRl9zouh2P33oEy+jqhnQc/VxPf0aB9ZIuGcXknWC4bPGc/5T
eXLWV4o4rWXjvAm2e8kK5Kk2coWp0yKkMEUOr2HS80/qcrx9I6vEw5+FrvDRNz0+
Awk4S/2HMoVyUdiHAJtGXmLtpbuFs8+P880MZ179h9UI/ug2sztWWc/ugFOk1eFj
aVEhrjyqCWkWLNhvifwnch1AxrrhE0su+TaEtvrDL36kPJaDBEvYFG1dC7IQpEmC
cD1EXby/kYIG3STctWs8xeEh740vrdJVKRGQKyRR2AzDx33vunJCZDNp8IScks6A
LP03NzBXMBFnkRV7ULhNMWUkQG/HV9VYGYto3uHx6XCRJTBHEiUo+MhN3Bcci3iB
5+bmwNQSoNEwRBCfrnbGPwheU7Xnm2KVVaqAQE5REDlFp7VUKdViUQbeBVjqGBg8
IVgTaeLW622hOuhK0F47plial7JSjBPwpVQSNFBPPCIBPTvp7KywOzlfRgbVLCpe
I/NMYw273AAaEYXQ4MHfMdZDI0sEESz23j1yTUeZYeh1GqgP+pZkadFCc7YsJtxA
iw9RC6mwc4IafXACjWP8wY7ShPZfjZ7ZH1TeZOiZwEOgOKt6jV6Kp5WQ6NmLxHus
qQWU2G0JYeWtAhfVXrfTuCrQ6TekdKdm1vTzd38BETJ7E7XjQNRaoy3cXk/4VXdo
6c8tFZGRjKHzgm0Q24vzr6eQ9CH7A0MnKar/MuTIVIHKAm8UzUZdvfWiyY82JG0L
al9SPpA34IjPMPVQpr0S/ABpF0b8Rbi3JRDB06hQjLGKYX6dIr73+6qMmOuQmHaF
73oLAzrvQwlg+5dncCXYus7HOpljk3IGgHAQoVtIPKxJESyZe4Gc99xuuxBPdV+Q
E7NDVKWiEmPs3mLDg0OnKm3TLMNqyMYkzyoujo/dqPWV87N0WMCwJ+GMZd/+IgjX
TRIF22KEX/ucOfCiSvX8gF/I74xmmCzESDdKonKgowwKX4CdCd90t+tuwQiFr/m8
gDAFqf5lRpMj6JNb6qTJSzihzw3zOF68oWq4d88jFD7SEBWobu86NyVN1UQFdcKp
jGJrreIwLIpFNjjS/kXyBRrOQihUvYhPckQochvTxpB/T4+Hq8sYy9KDQxpJqUKC
kCTnvi0dFaEOexcUydetG2dLE5HC57vC7W7gpwonM1IHo9kMQig+HwFYglAvIyh0
r+uvb4WHHUwUZIUul5DIXmjShLcg+c30F4t5Gg8bTIwqe6LtghbVpA7YgEnV4U9H
ZCLCIfVFYETo9UbY8403X1TCilQ783ld5YznWCWZxecABMHe8K2/ehi5g6l5JSY4
i5u1TdVMHdHAjKNW3ckdyTWdTHOdqCrYg0kDA2z87QNuJ7vhe3WCG6piFbCd1XNg
GL73ru2ftmHI3DKKBY2y60TagzHc69DyZsvdEoBY37AfYgRIauVApik2QFX6DJ0K
+JSzBnc0LR1SP8Tw5H78hu+nOClhcvZCl7VbFqdztlbyzAIUHRAHGSjhUq8wBwvn
Kr+zx538s0nZERKj4FAu4IyNU9sc3MS1Y8qVP5pSGkcSks164noibaR+HXbXFydz
LljAvurVfemRT8aucyA/Qxrk1AURKdBP062yZOmsAONic4drAQPTxRRMJun0ADMq
2qfwOmDUW784ZEP2HHBJvLgCaXjFvXeKgDObXFWicBLbCNAfbchYU7yD2TGIE33n
6e/+QoW11E8xc/MHINeOUvt5iv1orr22P7WGUSlgYdFJIa5rgMageTkO5yGF3Z2r
jHRS/bNT2vxVcv6OgC7nOklEGovkS/MKiNBRUhu7MOnqGWlTg7bG4VRVRGPgtr4E
3ZHZ8BaisDJHS5XFNZOzhtiwVAMOhwW09XLXwNVFHFV9AF1kN+95+mS22MmhQKKE
cAZ14IS40GBA6P2ofoIpZ5VVFD6hnaib783eqGTpWgUE7b5ouVOejSUZSanCZg7/
DfGOG+XVAGvLv704j9QD3moJTHXY/9EpnOphofd2ALqKSYKGexjddzVOtda79FuW
YG1SCAcBgJLky7CZkrY3Ltl2v16CtWZ7vTYOgR4iYJAfMGA1idF2bM89dlHNGeIP
VNjUrcE10sSRvVdCsWq2hm0CFneLM4jAKvwXqQTrscwm54qhWvVyw6A6Y2e3fubR
2ta1uRocKk4fNIVQdIKTvjjCSgHezknDw9hb2K3hP8RkPuZkV6TSScakZw+R3OXt
+nICiqjaiFXZRtCxipbVhlUGUkntnVdHsZHTF/uvAM2Zp14nzRhWUpQvhvKGPAEN
z/fxGQ5jDBnFACICYA1jev7/JWKxSMDHnif0q7y5jxar3rZ9xsrGrUZDwMTam3Hg
Yl99j5O+RMx2Kz1O3E0/ik/YuvwERkg5qKTfFC6FosExGB1CQvAakj7dBK/xNN2x
qFuNbeLywOCFYeTbiBll58F9/Jd+uioK5VVeaXx8H2JtXOqzRj+GfSQoVa1wgpAX
+enfr7MLC8nOAvKU9L1MIhLZxriXdE4EAeCpQii3+qxRou4WHR7OnfacJU/AUqdR
KM4k2+gp5eHHAmQFvSQVIuwfPupI0KJxaFXr0dY7jpjEkPu+rNfA5mnM1TKKbFVm
pYGO7bgwvnYjNlkG7jkDy6WT8n2nm3Q8TpaM0wwA4drYMDQKtUwpHkBZf0C4uJmm
/jNhJbmDKGuCmgJk185KagJ18c5nFajl0UdkEPbuZOhcZ/Zcfe8TtQ8g7Vn91fPZ
dmUd+aQBo7D/6jqa66NaIjzMM7cfgpeyU82g5qNcrUKUEwgJxSwI+QY2evpI09Hh
c+sqh4dHuYLYZZKZSS/2ycUxC25jmM4w7axEWef5VM5PZY/4TE4vRHio6GZerdKU
SI+gKDmj4WeAe6D0+0uE47djGDOHTe2eNrCOkYutN2gTQ3cQysFAtG7rXqQt/adV
T6DFrtIxnBTO6w33IPQtm11GzNxW+oj9TREjitHSEAi+lN4jdVkfOTwNeRvGi3Ob
IYIgqaiKGh/dtw2DJinH2pDcYwNmPpkAfBsfu8Whxb0f0PDeBcOCG79IcWIWFO/j
2stD2I7ejQSEOfoya82W8PLnMl+12l2a+f5YSv8AUl/yZIvGnz7OhIg5EiRmDA9v
YzPhfdncYkstEU+p3eECR0+8+20+2SwxhDLA3somOe6LPZ7UW0b6rCoOLDDywDoq
zyYOL8GQ8IoKCVrVmfpF0gzNQukJL/7RLct8bs9G/JFpaexGnUj4I4B4n+xt40eQ
qsPzFBQDWNs5pQi49Vgj1XO/MlFnqaoDBgFqVKuKNSv+/TLZbT/Eg5EJDfUJzkQh
iUcLvqylUsN9Vdbs/GEN11jLFwH5BagJGp8+ql/yy2938qBTJTr58Mvmoy3m6koX
SX/ODTPBJtraCWSLqQ+pVMNkTY/qdFKL39X6LRz2PMNx4egb8Dk9YRVwwDq2V8aS
OsTRw4kpbK02OfBCzLkPieCpy546+atytUzZJvVasWSK2xrxmFoq5efvp9Ap+2r8
O3SddY/VMQSBl02fcLl580epH6Fk4n8jgJC3DVkgqq/IDBEwMvhfZM3/9qYBgBy2
5EXnEeLO3YziD9zgibd/261VQy9twwwfZdM93seKyAeRH+TFzz4OdkilOnBMJdyf
fGu6sp/kz42pKJKBh7/wZudUZ43ov7aOjzQIMKJJk/jdBxJOEf3jJtEwRb9E6ZC0
jkNEggwEwjoR7gE/P/cqHFWHZ4Bw2pP8EsJoiW2xwD0KqvtGmnPD2jHTY7xCHyTE
qlIpTfthejwEJrW3ICQzLkFHSBQykisc37sYXH4D8RfCCjAaDdjcmAaTZjTCS+sj
fkj39pllURjy0XN3DQwskOA1XwzPXak/qRLCN/bHMREI3pf53Rs2tXTAcy9Eetr6
mTHk2mYue2aYbUfbyt6fZ7l5h2iStdj3Aztt8ZxVr4YuZpjYLuR9gIcaxlo9PNR7
raF4fJ3pJHWMK7LUVP9xiILHUyv4eponnRUCcgsax/WHM2h2nt+tIQvcqpzvnsnF
c9fnVKoZhcmBk7dOVo6x1gHIvzTUKbTON+IgskqvUkM5RVnDw3p1EvZdKA3Jy7To
YcSDP0u4HBKkKhY2tHSW55jaqFTiJvT5/kw/jUa6eBIV92omiINOpXXMqnQGg2FG
b6IqQIRfHeIJFXilrLDTAx4cWL/54+hHi1VHxtwsIra8GfClERYWMcgLFLBVE4SN
yyHjGVWMj5BkQEEOCSn9khNJq6b29Y+G0fJda5p2lR4sUtAc5LmWSb66fwHnBGbr
sSu/dddMyzQZhLf5n/FHiyrXbYRitgiRuFywdKP4hsZJIEZ0DTkuVMcncvdOl8g7
qoldGuJGwy7DeWSGIGS9KBCfAzjQmtn9/Kv111NunBivrKruqfIHah9fZzvxgQI9
rdj52aObln9gsgzwTWkeDvT+D0jPwgOZ3uup6+WrcekOYZTgY9la0/6QRWn4ZCCT
xmN//54/YK4I2YWuGyXj89vk+oYNui8HPyYcZdeHgY3wiA1gokp9QuRSg5Iop5AI
j39XI4O/TKqf8DhK1HLy/TXSc46x3qeDCJATbZBedd8DQCXj53ijY5uqik6QkvcX
HwNKEShw3I5bXr4g/PGLQMUEl24fV6I77XPDb6EbqUofQfHYbbawjfB+d+Ctq2PJ
Gese11LQ8sstqFo07V5KVB0GIYtrEspzWs16K4E12u3rdKHTO8Nw7WyfsBD1Sx+S
i8OB7BqpySsgEIsQcIxiveZLYHP+9S8B8CtITcyYZlWdeWuxwJ85mHQZKhxG+c70
FgPITtUOlh2ExvjzIyayYgL9q+BiKHR04WnKLLVNkL9dJaOIFA0ayCH2yjeCP216
beVSjJcxbEzV6cYgeeHK8AkuJrYyjtJA1uD5scIK/oVz/SskNDZBlIZ4sj3dVyU1
+S7qPNaf9sH2AYNe56oyt1q/038gYFxNgG/LKu1DuVGTdN3seX2ak0mL3y8YvyDu
LxRZFBUJAsdd+4Y6nxT5eollokY3ay9nnhIosjholDloRqHYdiIpeWiPjX+PrjZB
nwH9aLkXVne01V8YteWZ1lMdsxy0Ww1JYK2IhvVoHlyJmMqEcHik0UdofdZ+oTGb
DzJboZE+GJKDha1rJCyViV/MmTX16QobqDuqvtg0iHHRyeJFJEDMBs9i8zGpN6AC
qtLNeatShBVdR4FZd2+qZ17PH9aDUjwh+w4wR8uB0r3XZTOKy2cYvYJeB1uPo3xW
ZG+ZwG7pPVj3Z4J04mQc05Hfj7Ivy67HP9hNsyEIswbTQ2BYRNxlhu3ecXaxcTck
jxooTt2O50b82Ed4z1d/FLa+7G2KxdrOyrORvOOAP1B/jv7XFMznzcg+20NXVzpb
4xbVM77MroC/RS00h3bTWPcH3TrC5jxY2cG0ZkTWckmFtueV6SVRRbhdsTD260qD
IdZC8/nRcFJKSUwyFfgebyeBkaK97vtDayl32l3nFwH42BbUPA28c8n4h9RKWj1c
zKeA3bq8hCBZJuWWMjW7FZWeAfYHLrXCxrNbOHrnsIukgUMaPcxiiRBwpdKRNNr3
Qf/hF2xu/j1x6+yc/N1JHqsDv8KO5Dc+J45MhwaAaoT+NxoP1SQeMDiM30bvqDrr
jb2+r3gs3Ps065DbJchJ+3wDeDGduZM2tDQlwbdmC/3Q/rVhBDk5zDrany6D6LJZ
bIUw7Bu6zDgZDn544yVs/dueloXaoV4Nom//JhloCrwqS/cwqF97BnKBKqUhhGIs
WxO+OMFmFdKzwKrE3wwJ0oPbHskpiN1XmAGosvZZBCzGMxcyiP+PiQGUst+ws3m0
AZmg8SfQZ4heFLW7g27o5SNI87DUdlpK0dYdZo6iNQ/F2SbQEyzlsw1JIF2Kc2g9
cbXxtRI0YvmQG4+FhSMT4iSQGwG8xU0tcY3yhetRDVO/XFiApJtxj/UEPNDYKLjo
/opNQtV6+S1o14CgBhpqMVX5WfVUdPMm0bq9YiQBtUFp+nDfU/lBsBZrwjWsQ/os
tEzgxU/VuwtzNN0uJztX/yGhP/GdvNnr3Tt0wPHovsCGARmpeiMo2RZvH8Gx3YXe
cQsq6saA3Cj1cJrQXc35bWY9I2qvzyKd1ae8RyaNdoU5PAuYDDbSntonzLZGP64y
Go0ffX7GbNFINoaiwcmjFJJceDNCmKelxN/iWiawO/1oyxTjnJPxq9L8gXQnAMiG
L/oJT9YWtXgvLDCA02vWXXcu3I6aBpkJYHsyw2haPHCZUIv/NzgKS6i0QYBdq1YI
tBdRB+1fVfQdpQA8lr2PEDr3AjP3WQAMG92d5zWoNIjS3bS6ZRXcGGRBaqtP1WcR
oxmTekLjmT4JzUToUHqRbQ7ZfEb8HmFE1b0lL0UBIjpOuJmt3qlRFXgbUxkbMb3l
Jb4u+3g9KIB11V4s1w0A1soaZBMw04/WIWQntwUHuxuw5ChZ5abyx4f+Uzp5f4Uc
qne2wOSPDYQGnjqcOBhoKd8OAMLWs2BWUwuSkLSU5n1JlV6qe4YiBSpiKwmqGWLr
Bmx1tX1E2XpmHDD6gS1C52K4WWE2Ri+8QFWLNpWLnmLE+1N8YN1QskBURf6v/Te3
Os2C7V2Iv961EEbNyKXek+5vwpQTxnOyRHPsBnwBCNGh2/FlaoSqlsxGYYnPoRwV
/NCbmNilrpJPmgdV3lu3v7qnqsuFQA2GNAWeXP7Au3s=

`pragma protect end_protected
