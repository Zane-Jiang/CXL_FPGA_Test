// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
sOFG3IoPWQbtYPkpSh9Op4OhRn5iAWrhDPpXEVofaCM6RAKILo5dXLo9Xw/Mvi3h
5Ch7M3SinXdwXOcSvbP5APk2JLszfHY2FsuJbNB+snaMoAOz9rUtu6zoJy7c1sOU
SnFE0RfoE8q3EBXDlJj4AniExwPujWj5uFK3k3E/ADE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1744 )
`pragma protect data_block
pwB0GNJkdJ/rhWD5fHE4bi4T3KQA6MmiWlrzRLhyHsCJEn7sDSvDbfqz45QdacNQ
SrR4AyMRmtWF7Qz1uWfS8cYvhIJmhBwGTmTPvNsPzJx4yT+rHlZlZb5zOddBy8y4
ICNxk1QLKhm5/r230R95OodAJ2a1tGQ7lOFniRJ0PtjoNRa4An0STTZziw33b+jx
sdq/48tPwmlxvjEb9Tcg4r0ODsGxjvX9HeeT2CWa0+ypgiUv7eXLg8jkKkG7tb5R
iVZe+p88FFgYdAuuDLhVLcATFURZzGRjqf2oY3w/5Qt1HL6/l8dTTWV+sj+xaxYU
ckzfxgobqCqRV2sydkli0fuFwdo2swy8SLVSnjCPNxBYmoQlBH4TJLWPAB7eHaPJ
ZDMiE3HdZ3qBjcJaOMVb8jTHeItqQl9InlKl+Wkjc9KCDfNTc+a3vZNTD/O+aM47
4FBRg5qRZqBovPvWuFiHGOI2Dqbe+Fv9Jc7GwzbBlj+0q7XQ0q6bug6WGLs71nWH
K5Nz+01LcJHsyTfQo5jslTx0dBjWTJf2J4bzFx+iVOEGiiZRJxhWFJScEdsIwlPu
jJ9yUzcJGdMIZyR3uadyA4XMDdA1Ieckfzs+BPB5QAh2u+PPY0cnJJXCP+5jo/3s
NpRXqaEEN4OV4ocJDZiMHEaTQHhuFh4aMsAN36Cj7cOf6OpSOer21vL0u35F6n1I
a+WxBy8/PkQZtFeqDtq37OHUSJkdxCoJZDPVnYU7tc7AetWotcotLWqIp49qxR8W
MddUDkNe5DHP4ZYgRsnV0O66DL56IYq3UQuR5bxX9riHNg3S+lQiaD/IlqpHlcFy
4zXbqSSoRFfJjZe3jlDky8I0oNkxTsco/aCIM4lKCWNoYyij0a+073oVQZTs8D7l
nYfBjVOcazp+aXnZI/Oht/Ys2ZUOCSk//nOA0ysTlbC61AUXkBDVfL3lrL+TbFJk
urLZOnvqfZAID6Cc93Jrm58dldX3BdQNKnnzIo6QYHJlzE/PsPiXZFI9j3ha3oSp
C/kWw8mUz1fXNNL9I/CTKSMD1gtyu3ltpYtbq6Asu5zSPDlE67Y+OJCqShL9+VTK
H8LyUhQf6KcVcaS4nfn1OzTfwb+zTd0Q2EQJ2d+s8JbZbczqk8LXTR02rUX9xDL+
CE10+JVBf6aZo8TrfZMASnb/okI9+h5mzn7xdibKmKakw9Ywn78J+3kl9TpDU4Cu
9ZtTnQZoAeWN18bbL5HxHMANa5AiO89ie8o9laNvWm3FgZxoRYEZ/VntdABlOv8F
9zgHm+5zUxkvEM8DNfp4CxVjA3qVLvfoldk1XWSFeBwUfnsadCWRl8h/xlZMQtRm
Wy81KtfySnZv0HuekLw9EnqZdv+mpoUuV2F7O6ERQtin02k4tC/OJVLSwIsY1FUQ
4H83X6hBYV08wFVpqKrhVADLG65QGmJOHgAoZNAFDhx4pdgW0FURb9rPB/AiYJHd
bV/owy4kmqU79TZJ7Fr8a8Wey7pQRI/jzO0N4FitlVVfnFAk1lVZE2BhI3/DH0Ca
yqeQy/UPRpwdABbCSxHRsLUfTNKw5jwCIHdA5Xoalgo+XJjLPWM1AkD3whbI2HvU
PFh4I6K2Tk7yRb5dhyVblRzFj9gwcJNmVNCzBYAC4RbNEwhGlYZ+RkCyp+c6t4Ci
lf6DA3J9TIun+xNnbf8f4ZehOl9JsuEmpjS/k4QzGXoSa27Qyg5oF0JNqRmYq9LX
bhl5UZRsKlIvLcF/G+UmsDPhdXyKxeKKr9TUc/tv2LD4yPEIVqRu+X/DuJUmo4zy
kWYcP3MGFldcLQuGxlUvfw3ABYTR7XRWUOxC2tK451kX8BfkZ8Djsc+DLWxZFv7p
7RhntjtHSZtdHl442Is3EHvfi9Mn/XMu1n7Jk4enWRhCobzpgp7UWtiFngIqdRFU
Dp3KPICmLdRd3jvj9wLjruROXjwiE+Hucxfsg7ruDaJ/KdnO7jsfq6wRvkCzeEpk
nXH//mEJLaLptsJ3LdhUJftRc9a8WB2KuCSiw8HYygUCnNsnpgewULvLSBt5U67W
lq0rv4A5mxXPyHtXbOkGtOwGQCWJkGkVgK4xeowFFNcDOvU/tcK6cQNI2NmkB8R9
HWYCniq5jdKGb8PatPELXYr8ZpyAJcLilZhyu/bEmXcE/tZi8jFE74yIsaD9q185
Q6EUHbv9G7ebec0aBA8ticqp1Ino0+8ct/pTRzzektbrVD0BTu1jRbW9F+a0W31q
8Df4OIbbRoAEtxHsRMG+xbUprcU53L41+9bq4ZDIZ7Q7I+AZ2cQRY9WqTzo2EpwI
QBg9t/1sB7VKnwDjZmsWfA==

`pragma protect end_protected
