`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
epHJgUDOx+YhonnreEH4OzVbRyXwjedFyUoAox+IDKPlKkS44RhLcuLRXfBiQ25Y
Fm0MMsti8TMZF/Luy5dq8ONJAekaV8aRvIVmYnC+O0Tny2V4cPDzg/309ldCg7+/
S6uVjMB9KDY/EI9K4rdqUxl0nZB4qevsdMKKWEyRkEY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2352), data_block
R0Fd861aFKETGzHctFFuMiogg6K+PLXFEXvONzWr4bFbBE1m8oEKt7leddT+GYgx
Ersph6qRuHZpEnAybaN47q/6pboRLeuJyn9xftB4w5AIqnzz2BzlERV5D210pby7
HQIafnvMaZsN99/0E6aTs+w43nO++7Ypn7m5OBaVf3GO59wxzN4X2IPOe+ziTvE7
Giahj+uqQO8+OrdziEUIYnuv1Bgiv/8sFqcuweQ5021rNS/cvTsLp6+nBozZMFhx
Ze7JiahFpXXJUrU27+sd6UT82h5cbl79o9kxNP5EMCaqn/gRwHu047b4Yl6JfgC6
wUfymQFRtAtOoHgCon+5MrkvCxVfmSQZYjvO6567p5NmCEJxqu4bkeoBcYICP4qG
W1y26vhSimLBLLpfwwf61x6IEkMCjB6D2Wqyof8h2iTuPj8vrAUnBitq2IuaLqbl
CgXHL/Gu2cC7JmsJFjSMRQu9Qo0JMBc1vcb7P38MpmyOavtWb/gYXmCFY6CPitSS
Uzf6f3Ic10TfZM5OWNYTsRYoTMvaODUa5pKv7BrvrtljDbl1zIFqhrAkMDMnMEcJ
KNqFNzsDsz/3wWH1H4ZbVZ0yfuCXdQOSWzi/ABGnVRX/MkGrVGgOIM9k22geFJo4
PzFr1a3ZUfgeOT9MV7mzH9nSO+SeB45VuiC7nATK/unrStoZmObIifTyuHERkSFI
FMCOk8TZ5Rc0+DMGQyzZpC3v/PEvR7zRWHBon371895QUdGzee3BGT9Tmol4AuJO
BM3ywSOPclXEueBjB2JTWi+tJZ15AVaH143bgFssaVuTm1vT9WW0B17YbXP4mU09
/r5mC5FTGsJYYh6bGdEI+iPsgaKYFJwC6wAsC6EDaXEryw08eaRDeZPuCR2wq9OJ
qyhMHto26uW6pOPLvbe3nGmVPU7LYblUP0nR7E0GS//gqsCyhlQ+8scIlHWboALE
U/K9VEMXBF7/JF5KdA7HijmsaTHPml0kiNKoH/2WwCTwPJUi4k2fBGIorIDlhWVS
Vlb0iPCKoEE6HmP9iQw239aEzuBdGrBRLyr0Kbf5+8YwkGBJkKkYYL67xd82Wn1U
MGgkURfgT0SRFe+cpixP2rf7+etrxdKpnoxomE0ZfUoKiTnmS9xPcuXisPsNygU5
uGXvsCHcUJ0o0x/cOYkd/kCmwn5XAIpJ+tvdmK2X7VnjpsyBVhTbVxmlI/AoYT6d
G+TkLQAIuSkvkLN9A1crbcmO81U5l34a520A81rwmtfKIPiJawktkQ2Z/5rCS1nm
/KFBn2h0BT7BNdq7GYRFT8CRWF8Eaa4JLES7MzLblwsk7rgEErBiIrRX4clm5idw
XdeMpAQdYICbqacc8uxmmgCK4LOhfDT7awKDZinddETKeQ/XrhQ9Rj6TUY1TcMbK
N56MYG2hhz5U2teujBrL2kr3eAS/JKo4NWTm4TjFTvYgaO2Ik1UlznjXi+2DeR3B
7OEajYSZt4Frz4tg27fm8X4yaNrnujg/huTPxRYsk5Dijrf4+MRR/GLvJxTrmYJ3
O20S5u5KergdOvBq3I3T2vyQ9A/1Ld5ukIIs3jkwfafftY6yIxux9tRf0ZRxyUN7
SW9GuVtEgb8LKvLW5GILSQHeqxbdqm+9b4tgMdtBu425AgvwRJ71Vvi0gQf4GNlv
3r0e+9uDzGw6ANnivbyp2rnyN88dfhZuTct7laTND4ehtMBWAaQzbemW4CsIrBAo
fholuax/0SnYhwMfWJgpG4l1F49g4BuwHSnl56iYoTkLMh5FYz0PkcXNj2+TQfNO
dMIdjwmccDbIRdawQWcOww4hlJJIBOuiNNHVHKo3FbVsAe7N/9qEt8AWyblPMn+s
TD79TjYdbsvqTMKYPWEBG8R1a5U9Joa0mnaDW3vJqGXiinzJTIDY9B93uE6REKnq
pZYJNztq8H9JuyXfs9rbQMfzRhrPJViWY8YONt+tbZh4RsMxdKDdPHALrB2lAR3H
2fVhByxXER9/t5nuaMHcD8WVKls5ymhzIYPnyU60S9BRC/+zeJmADl4jTKJPpC6m
s6o9LzH4prxLiRZh9DDVVeNBhu9tBqSh8sSLzSe5CrrgtJC/sU9BaigY06uWf5iJ
GS9l2JZbke/e8DTODrtC3H5Yk21+t+Kv7MWhgNja4X8PclmCT7P23fPADrk3/XtK
i47OJIyO3mqm8pIS9l7Q8jdItpPlqyhObJoQ3AAC40NsaEBGefTtWyTwWdqJVbNI
M14H5hasibBQYTmYC5jFL8KRvuJGzmDt4id8vTBgxKG0XEJ2Su0e9oYuwm0xME57
Nw2Cwb5PocIeuUFZsPTWy3ZdIWd0Xsrzs+76/HzL0cXEDQZ0rpjgNwf+CHdhwcsk
M7liqTtU37VIT81MTV2g6Rxla5fQvO9tZfuuaoH9VZO2rENNrNnS3oTncRQzHfIl
k/GVBguyZURkDH2SXUPUP03ypevFudK2vn5z+SUZVStj6C8kilwIZ+yid73UC19p
ZcY/z/ijLIbmrHt6h0G8QMOCK1LbC1q7zfyUW883WUi93tFWjRzIGgSkQ1WEZLX3
gMkRJRKrTeps0RAp0+eRSx3LGwRDDCZXsHXrrE7YWdxoitu+roVDquUUO5yFyhwv
SUpvAYYs1TlBgJEEeJw+Wa29DA48edCXuZSu1pIHxwz5FO1K07DteLlm6apkDpX+
WlXoXn1EGqa3uVHtSrivCblBpzXEQWao/frn215RaRoCY+I11hwqf2WMt8fId4P/
bUqI7ZkV9lyw3jOS3ija/Zvvi1+Rk922/1CjvqJEWxawkqzNN/J0G5qkX+LJKaYa
eEI7YEujjJ+It8Azkhhuz2nIX+wZWsVIRCkyF4ZrEyvxapM9vD4efFdqHIOQrPSc
3pSR7GT9JpWtSUaQcoLcEzCRCjUTYF8ZHuC7J2eD3vKf/h0Cgg7lhVw7vHHpXZls
GNbNTiaHOC/DIJhn4DKlJa192G29aIMwi+alsO6W6GAjyv/z67M8bMmD3Pf/OEjr
1ghI0ZbW0jaNOYSG78/vP3MR4uwoDVLEpLS71sI0ktQuMNfl8HpCtAqqcAUsY7BW
smrMI/Uj3d9BHcYeNziyVXpLmsR67qzPwuzNapSz0pT1Re1PJxo0WnrUM35t1RDv
`pragma protect end_protected
