// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
XGIKzWoFFOZ9HfgbmUKja9yedaKdvwevqh4DvOzKnJ9mw4oYru0JtQATnIKahPJefE0nudCSzj4m
njdaakKTJyGxHqhGtOPOkwPThn79+rYSA+OGpgWpbsFX4lR1uLk4t4qGkO69LyWJkgUO3SkFX3S4
vP0vV5DRsmAfeOTnnmfg2IweZuTRMVQnFIaW/1RO1ILmdAk/mW5Gf2NuXhkz4w9G8dtYPI0O35UO
roD9/vl5coOzeH3WXmtPORLDajtjGMb0vtsXLZ9aw7bquIDLiEZAzZO2EE4AtCRkh5xPczppMJ0P
se8vkU/n2tqEMiCsdxWothGu9MMPadyTfh27WQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6144)
gUeTU53TuNV3Vdic0Fwojq9NbMWqy9glyY0QMcMrJ2AtMgfdSxRK7njrw/3zFUZ55QqTUe15awtb
/jHjYaEzjIJWFMoUW1SKo1JOSDgH4EMSWyrOPORd2Cz76ThviSqjJlxdjetkWJYZ6TTYxmuOLJNS
1LJPaaUBseCzPMUE/hhjPtYv9uH7ULiGaWYjdCgtlWix4vvVD3Ii0hhqmjbxNdtNXQbtiBh8Ie4q
Ip8rroMOpkl7sCSqzkCW3TAxcZJNvLJ2ZeS7yRv4AQbD2zNGwsgJIP81GqnR71q61ZQI9omFkzwX
ThBlyAvFJOf4ljIRdz74IyRV9wiSa6dbotSYxDxuPW8Q5Yb865q13a1jO1nm7poFueJHRN2U6x3G
N0T4HQdG1AjFt8g/4HQJQPgeiMNDj4xlqlCR+RwnWviCB4BlUqsbXKaQ4oBZ0po5vqSNHNNopJMc
sm6iPWKLrqWhBpAb0wlzCRhLeEXEWo/QoY+22BEmPtmasxpH2yhWgEMFkh5/7uuIp3mr03zDFI9d
Bc3dYiLYHMpObGCDKnSMCsIpkECcrJmOBcghNKoErSX0FfPF/whFH0DIdKmUoXkpF1xaDBDn7w3p
2otN3EcoQOObWBBCX7rnqtR9fxI3lJwvH0bpZwps6XMGb4AxfH0aDpDpBnNvcElq1OONt5Ujsar/
ETWMmjAglijajagB0waHocUE7NtFJfjzuHkXjihfbELagW2V5PPVJ3XstpUmvlOcst3krl9fXnGX
+oxIJiTHdoS9n7J1XQ0a2tfiGrnvnsoSfd/9Y61vAYe/LXb247Ctq9z+XSESDqwYVSf4gjPmtMSU
jOrYkOt7TVBRGPaWeVReQFuSc5+59YDv/yiemnnh7YJtbnc2vz8GVCD694s+z179M0nlDPMLd5dj
g7J5igcb4u8UuhR/U8ki0Tm+WpmHTynXVLYyg0C55oKXmApbtwBJw+BElhWyE9bY1bPuX5JfFPo7
EOY8IgH5k/KqR+SEMBrLC8tVqEsrc4FytIZuvSIH2kp1g3Llxn6JPM0SeECho7wrvpAhDRRyzeFl
aRORWXsijFSWCAhl4UvZnZyszYdMnnQGBZ8kB7Iqk8sLwcemoCQBj9Wk8/2exlrOxhLYLUSEPhNT
hSCR69uXZVdZJS/ObAvFxUjJ1GEMctT4V8OjQ/QnmvNKwXO5B97SyYNZ+VKP+4a4WlgBEfbCf8Ji
tbXhyJkM+8acNxlBORj1d+gzGyxNXtqevo9zH9hqi4mAtQ7LQC2gg28EdcRII85diCnK+RFparcF
vthWrwncdkjHB3jIvbAQdg60meq5AeFrNziXuLr35O0Mg0virIwD08fqcDCp17PRjkGbqYTHv91G
JkQLZsw/isU736pic51OhvyTcse1BeO6Y4vWhaXuWKNWdrq+zaRs3mi7RUzl+1zuj4y5vx9hiXmE
DCvEUiMaMm+Ym3ijb6KAdVr+RLtfgRZQd5FdTpcxKoZJUJOxILVuFeRS1hR+RAWIibpqoLA25I7r
8ziikimTIR7n5rhkSWotM/F0rs23CyiWUo9CYw+/kCBSm1uSIvCG6ARZSYvRKs2xkKvh4IdKsh3P
N6Wqi4+kQXSmUdUNOECAA7/koyWmdUZ62tmIyYaq9TGCbArVcyJJdUkIZxcZssnHW7W2vrF3xlUH
ZxAJfjzruObLEmE13g39PJ6Ad1Pps94+5WIfMA9vaOMkGhsst0azRCiJGRmkewka4RfBRT2p86SP
AmdmLfg5RF/s0DoVEW6mvDos+Ef9W3hDCSA+p0EmXc7oL6laQj9XZHanlFDjAABw7fQ42TxGrITe
kYvafbFxXPTqmkXR2gH/rcPOthkcFuSA+PVwqViy/llAydKe3e4zh1uuAVAxUpCgFuX+FOfFcW/6
qj/VmtcWKwr7dFowid1o16m7A1yFojiiWQBJLRe9sQVg1bWJ4Yxx58+qKhXU+BAhL7bjVIfQBoZS
1b7Yry2uVk9GWzl2XaUl9yNq8EoBt6KDXoZPE3WmHLHCNaXs3o8u8fYr+JRzpcXirDOV4Cfs4ppd
goAw9K4XuoDfPjl3JK24Qk0wP/hsbj5GnH2++Ybyxd6x3WT1McNLoIY4Qduqis+ys7YQ6rKpNJZW
eOgB898qDOIXR2Ou27d0pNqlyYxe9OsCDoKp+zAxIdg8+5zLwbPjIMsIyt8Fa2OJBZ4AuJOQkg7s
kBJGhr7yhR/RQgqH/AmYTJTF/KOrUTQvRAg6q7j+vV4i0dzvz/cghvaYue4xRQkK2vAySj0wKRTB
tRBU85xRLVINLT5f7obYA0qZvQAhq2kpqjWu2LDmM3AC55adlrzcbCjTjh4HgywoxumjjcJThbRd
QxP0pbVs7qznrHwCqscTw7uAjNYhsERDbNNoySvqdi/nsJea0+JKKucMeU3V+JFsQKvWCduQZQGB
EXeckj+PGCIIq59oc9aQ8i6uheKs6kL9H/5bt4nhnTc7nAjAAUm1jaUadfwAcotWSGscc7VdZhRq
+Skj//joAEKHdSsRcz3TLCk4GnWdf0RtcSnwWa0cHX3DbE/DtCCqxDqdXf+Nbk4V+PTiVW9w/f/R
VJpwN/MU7qdXnvQfZ72q02e0VxmpFIIfCzM4SoMjiY//SybCvF8NnQefgi9Qpk2F4CbjovT07rtQ
2ZJBK3w2Hjzs1xqhJobK8To7nhVnrVxc01ZUAwvybOBmEgUADYSDe+vbsig/k7DjN/Mg9HlsCVOU
x2z21XhS/XqgxNaQJZoyAIgE/Dt0kIT2mLCBqdq3ZwnxkDK+bjlIhetTuukK8M8sbL0R53zuAiql
tMtJqYwmp7bZl7+xZTfMdwFlxy900dib67dGC/XP04hlXkk9kV83pAbrEFV4G8vuY+w5nNntTBWW
Wfpiwa1o3wiZIPjMmBabUiVJ2jzNmEnAsY/8nuwMBwR64CrpH/RVN2X4tcqJqf4ZWoiHen/aceKq
3vhax/WMIT+Y9AQTPHsy5lWnxFGYg23dStufsi3v4m3bLlBF0jAmtAGW5iTHiI3KXxJ1YK7WEwzm
uHipdmU5sIHkoI0lIs9M4yo/x7H/OJ18llPa2K5+dIY4EZTTlEnSku8PnLeerSBU+++F5Umd6s1I
7/dTuj0jnSboerHv4XD5tLberf1Kf4jXfEtE+Opjrrejs1kfEtcgPR74jV933Ez9IvgqdO5stql/
wzY6l1xVCOmoyw+at2h3gs09pe7bXoP1VxhcxdNMpZqPnYAzV4ag7PNHvtjVcikKtayeq2yBJB2x
6OATiDB7/ZT1qmQoKBfoZ1B5TgO71gQwCwqNOFEw2pjlqpUaleV57t4zSV5SdPFDBwABZRzhR5nj
iTVAfY+kUtuWisR0G/1DQYi0bPACNoDnnCN76snQoiyePZv02SY3oGz2Ab5FCW9uoDeSbkYihdo+
3r0Ek/RcOI7inBMl+23jMntXWcWDDrFrPMJMGNrXr57FTuJWaHl4HHF1lpk5/EfYuYkVPn0jloV3
2arMo3YwJV32UNn3Ku7dL/g5Ot81/DJLH8QpbMi2wPQ6JD0rp2JZw3b211ZuHvn3PbzBT9JHdVkx
n+1nttX3FrEKCJGcISb6rKBqX0wNWUWuknkkg3QCK5pF77P0HfuhhEUxmMADwxKlD1zg05i0eMGP
y9QnFSqa5QvnjkIUa3NQLfkwNej1E5YMibsjAtg6Gm3/CE8pG4jaUdcrfJgd9z57AJr+t8gXq/YR
aXjASqkEuv8vIGbaK1CyksDeto07PMU6D3nToPiYqYf2mjsbTUKjXexCqXeQ+1E2viGU0MkJPIRF
3+ZVw3OHf+lnsXgqaUuF5NWwwK4NOPRVHTNiyVleFKDHkE1LB/BUkl0S+xCGBTrOtFFe6SiQCNqS
3QqTPD4GnjdR9CaHaXesbyAhpzf5bML0SwAM9hqCjg1MVH76T9ZLvw2reewt1jQef4R5iK9u7nEw
z2fAUxEcnsgJSBqDd/JvxQG2Jp6SrK6RZrBX/tsfFb6OVaBNY4M2ba08hz34/eB1VkSdK/tIXy9K
6odMYbimv3uI7rXVxrOCPTpgej4ZKT9wyqHQ2DeOnHTy2HJiWHaEKL8joKQhq9GQXVoWrt1c2Xko
s6Gb7mtY+RkYOuJfU0oBDjzIwPtGC0cTtV8B5uxMhceYVPcjgIn+x4NWEPOXKxfvUiOgAX4Oc7lk
DLKX+uf5J+6u714TIGu8MRoPMx6X/DFdGdCj0zf9kTyHkZK0un6GuAfN8izZvBCUcdatjC1GkT5M
ND/+CcdRH6f2taV+A14tiQuwo6+g8EpIQUHGt5obySkEkjuY2tiEEN/ourW7+cqv8GRwQk5fy/rC
RDdFcWFX85wyTZGNK3omgk+XCsFpJpHH7DnlhcQ7h4NyXgqAHi/l1mPiO5C98P4WUPMtnbl/0O3G
qeFTo9Ilh5Fj4m4JQfzn0XoBwec23A6TzzosaEabDRwCeuDvx5xgRZf32tOx9LESCfJrhnNJ1k2Y
o9zuz21W5KCLWwrFPTWb9Ot7QV2EUZsbMo4vkmt2Arx+AULo5doD96CPCri7U8p/pgXKfZ4Wcn21
Vd8ftwpqn/wuS+nliHM728lBWghcH6klsF4ZDv640Irtn5HpzXs1Wef0QuqEYtLdJzrrA9yIr3St
aodOTTk2oLpWFAWlr0ON2RPP9qWTM8M55cMgSvNq+Tah6stCOy5SY94BrYlp5iAAK/QBzUG7Dcmb
f3EfpXYNBkriNZou9Z8lKEqKChhefmbQ1Ab/ito+Vq7WVKk4lAOoMHPVywHDzjc8vTWkup4iq0F0
RVpf5uWZbCKXvTUbld5LViCDAxzIGDE7Jc7YUhCoJB5GP9UqUvQ5aGVr8zlV1CHgG8zhHeC+IJJt
vw4Sre+TXF4Pe3+IzCOA/RrAilGri5d6wHqdPJJvafXp4B4qABbyL2KSRLJc5pvh+F0ye6cOdTqr
fx1/HacXdmC2jHUy2tcTryIUEiLAmsgCLoPbeNrFIuPrIp8EjgMzGppbbGsJvim/qJJE8utSgljz
PJKl54hdBMxbxe+GrB8tTC5Ignl2fj81Jwaq/qlnrpFxHPkdQSKNzyLReOVLdanAe0WjGyLgzc3h
v+Ly8kAljJcMr33/qD699540hDkpbAOlIxMsRxl3N3nmhCJ/aOfBj7t2Rsxrb8JWXPB4QBVXoZFb
sjfjCQIbwBcsuVKGhYKErYqez8KI/wPTQuC++1PzfW0ZW1r794r62/awusr+PH9guYjURahOGxGm
+g0FljfE5C2n9BLVsVsw6NCuoQj/UTZBNhCOCyGzJ3EQfSCts6uLkI2w9Wlwq+XEnm/rHmDL7jSj
+5KK3nbehbChzckRQHjQZyUGqzPypmHXwplFk9J1S5Hkv1lwLhGQk4ePpe199wWf9kblYU5mk6AL
YJo0NPAej5sNP0BNrRdc3jq4dhjyE7NM8WERK4kDqFk5Ui8FuU1JdTohuRUhv+tPHDLsRzHMyfsG
8PbZywcKrgRtNnA5N1uv75OxmU6HJGiMcZ2kfbnshpkgWnWC6MPiS2EAJvVysnHpPu0LFWEEPLfa
/YUEzU7jGYJKtdJ3MH3il/ghqLr+f0mkT59fWGPXJqb9VGbUu4eX7unKrIUnehhmgMtDyK11JQvW
+q0FtD3I73Ao7YT5k5I4HIBw1Jq8j51ggRHxhoIld4H9aJvHwS+Q20nFnTHdZghr7m3XmyyoNrPI
X7RdTIicdRDPA8YhqHbzKThfhji/yWwx0t3T4n+NoVW29fUS8WU9mp/Wk1wCL5yFrwEQ8wZhVrTv
TRWqBUePK8dH4gRrz8Me44wh18eRoUdoQiKtnK4ZUbuGLtScMCcau9f5LM9QF6aDcc+nc4rc1OGO
R/AHoGLiyma/n5c+0PEH39PxWvQz23QT9L1ljoI8K/4h+fwaRxTRoYZPIO5pBdJH+rk/ta3hl3wZ
AzNP5mse2kogqPvl4vatvmF8DObzY/rHl+J0pRdm7PTYcRTsR6Per28k8sBgHzIvc9iZyKhtZQMJ
w/JKlpi1fmo9tM81xGhguw3dfxxmBLhTjC5iEHB+IrKxM0m0AR5MlZNW8Bh+/sSq5PaP7XzhPD3f
inSuNZdS3azK9DvaMd3TAPjiOap9OTlKEc9bsIfnTtFb0rBmmzQ0JaBiDPRXeZIJnxeiKxXIdCgq
7gKcOCnCpLVXMLiciuZXMfGM/w4/ULl9IZywcaEWLsUf422c3EFO1rCP0X1m4IICljjElWF88wgJ
Nt7J+jsuD/mQSlQ0n/rBHSmDGYfHI9vN38rHhTdOTiqStTgTVeMDGUx09VCcjJECYnKtDLTynOgW
CVl+KMlMOwXCg0LFUyf25ioqyug5yd1jJWrToGAXcQjLczn3PfqmAH9a4JKiQQfg9XXYTHFbH/K7
l8pRCR6kIkmM+0H6+3VE7RJcZA47NO9U5S0jISXBqn4k+yOHHOGopiPQx8XtwgetLnEuDZ80wBZh
kuI/3FzXrBKKs6/tEbWpHQe6lZecC8Dr6H1Y0XILUr2X8xWceNz4dK1/9mCA2Zg3L1zV+D2Uxarq
YCOWXAqeZX9JScIgoOF9gXtl3fzTgMV+ZbI15ObPkXtBSuSt5XouN42ALCRxiSaa8qXZzAvBieXf
colksom2xGOIwJEChJIazew1WfEuUFUGbH+pWwBlRIakApxwCYE1Yd3hGQcDqDwqe0v+853TysNm
950FkFxXkiKwTKO4y/XXJr+3ppWKqqcvwctpuRc6fr2HXr2GTiYQ6tPPsXjtaxKUG/+9DrAXZOcX
P2C5JwSbQuDC+KvNoJVAnJ4rkl0jxn9OalQoieAxvIIiftRL4Ljd0xaVAyOrz0giSj4XtMH5MJvz
jH4wyGaeBtJkhcTmipDRr9vEFqfmK1G2+9zOsVhR03Mg9voOuOqHD6F5AtPjTY8y9DxLke0RBExt
dQHkYpd4TGzuPjXO/GzQ0r3BgO6diA9ZipPHtcIzV2bdsfDU26EsPaVdTauxNi25HWbCKD1W8TKv
xJsJfwyFv36kN4PclKp9Wth8CQ4JNoNGwD9JlgizwYD6yFVw4/FaVQ77eZbdEIYiBnOomdup8xZo
RNaaUpDE+jvEOcn6YdAkJiYxlVmdD8dcLXSkqX3LqnGY0sL5yt+iBMjagfSv3G4DtkXFNzDOm+LY
elKkRSKiBRePefdksinRl4TmJRb+nyaHTRolFq8bKbDrNUhsAyipeiftPjmZJxy1tgWBgpaugHtn
ox4im6bJirIuxEPUQUSF7D4G/IgE78b4mWUhDQDF2kXd5JldBzARcEgAFtlpa23TGvv7wCn6VnWl
Mq3zdoImu5bkvVwGATQNoXXxtXxNocHAYNsnPapmTKSI/Hy/iAVVvsyJkPIs+xJcWpwuOX3vAnBq
aLJCfFRX3l3cbID8rKLQ/t25W9BBb9RV6Py18OxgV5YaaDUBfR0tzaVqzjuVnltK1D6MlUe2uuM1
BPv46bI2MlAAU8QJqMtrxlTDaIjIj/dCzUq6euK1ecwHobXBymoAGYvdy2T1gxjgkqq0X6hZPMkn
MeWQpZUBbePYjx6ShiWs9T3i1EA8QQ+c+5D/RkUI0d2O1YyR1JPaWgn23HG6Pbps+IMqeR2pGyju
jV8LoMOyzYasX51lDnv3Un9STmYI0nDJuX63s6pa662oSR7VKwl1rUi2Rd90fglSFWjx98Iuo2SP
iM1ZyflW/psdAI3gjmfirvPjN7y+s9ORI+6/RLKrIoEfWNrZQ5z0yRrXIowEcWpc9rYXSKx3brla
kD3lTxyiYMoJikLdgPPlO+1ptLqslPW9F3ofaeQJnyj0ulc/9s7XnLyi9+SLbWVqZbdbbX6Eaf1t
VAAjnQtPiClXBRV+uHF3iOi94GeX3fQ59AxIYVh4Xr9uAS0/okXRM2Zt+o8Pxju9sk5DTHP0A2cF
SPNTs/rFJ06ImXXy+6hF2hgJUfw5IxYSXam0iP+KIMg+0DLOd+D+/w0z9yMcmxF0H6yY35VltAkk
m4dwfabUOA7l4op10FJVKR1qXhdJ14DEjZ7lnewq8/1MW1JL/XEs/u8H92v0i6YipMF0p0AIBQ5c
8BHn6jD8PkxL03pYs/yMSPvGTSYMMfojVyR1eIrnI9GHCo6QG6ztYzlUBxINmJopqqFxrxi4ZMwr
E/ufeh10tdR2LXYSQMRMqCBScEfVjUB1UbLaKo9aevfXD7FQWTlR97cT7I5l
`pragma protect end_protected
