// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BDQLqzJ8vhhpwBCzaJwZSUewT0jqJhFhXHJybWQb2Iarx9A3VqjXbCcLuJEx
2WwgiaZN9XK0o7ru+ZQMBozn3OObIxMn0E89PDwDIYltyYeKD+hwQtC/1SIO
peibJzxPwy/L8AzBa/ertH8L/o/pBzgHFgzSODnJkjUtaUi7LaJHIT2dzB/C
NoHIDo50MC0ktuO/aVBb/kHjXZeLxFkG22AH1ngB+UN9y4YWsRRzojv+Mhlm
FPimxnf4B2ieqpB66y28yZmtnOjNEz2JVlpjemdywzRyBfwpbFHBCkoJiuTy
53H9Rzf+QmO0ReVuJ7yt14LyLtvA+Pn6EqxOfTTgaA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
es2Pu1g5phSCKiTlix/dGk8qPXL6VPDVMxZ6T9WXscOsD+hXBqRjUYNd4LRx
WoqrZbj9IpFaFIL0PJe89n6lezctFizh/dxrwQ7r6U7AupFta73l8SBeIxso
1GoK7OKoCQ6m/CkF7/kMqa7SA5w6TORWKHivsfy5B9zgMP1mVfteKw4shyIn
KvwcMKMKeZfIQmur0igQnicumxCRnuRaKysfNaK2vMzmq3W16ec5VGMLBt30
XjeHbEk6niiWQgYQD6FGDNGscr/r8+Ok84kkDp3HNI/m72vAayw8yPuIeC81
W1obzSGgX/wGF3ukO8LhP07D7udcw6XFRefOpeO6Ug==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FP+mujp//B6a3X3A4lbMt0ZB0eHfrJrQeDp63PaU40PvApdxdZf6RkQDR9mB
+xMYcw3xf6Wq0u3yy2Ryq2AvrT/8rDm4wMNYh5cep9qVpxLXjcNTE165A54O
xfbS3wrJf6KeBZFr3aAnVn66/FTp3WJIp5HjGGbaOsZ9jJZOD0+vpX46F/r+
hIENqe7CInhNLt96ORatsVQQ6DIn2sVg64qmXPPFQf1GRvM7Rqh7R0ZmDH1R
CIzMvkRXJAN1SVVcAYTxRUrDwQ7SXOJC4ihDeQDD4agw+Ea/UmL/TrFpWraZ
1iZ/cTGQ83t7pKTi97oz3BWtO5b9LcnNeCBC0rdC3g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
N7ZW//xGMA8W8ubRt2vZSCyUS3mQOLtxYio3+6NKxVhwTF2ZzZjWzW/hBJYt
AE0lC5GSEo5iHs6zYKkYfilYB3awNL92I8YGYLbqTmyBGlm6XNZ5tAnzf7DR
2GvtalZ1ILhqJiHoSoFvdmdfTp8/ahzla5dfBSRge9Q2ZQvVdZ4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JJoSF9s++QQlMijx2MB3lIrUd752BlpDzxYtS4sQ2xNm3Y+TDj2W9e9aBkKI
FxsaLXERrHNPPemk9tGbzs+PX3rynAPir6MW4aG08NzcBrr23ZQTWfm/oIgy
klM+8NOT05lFU5GS14eQPpeaSaztt+A7UZm8wCRMO2RDhoZmj0BEZbtc2wJs
buiWOp3fYTrhxCcYYUHvp1oe1JIGgwC41fSYlpYLIkqdiR4wokwtHhGrAWsk
ZHDXarn3/vWdsfXkom5q4hupW5atMXxNw/RU2zGrrwqVcpw9fkybNcNpCLzB
V/cQvkgyQL7FAyILb2LCg4riEM7cjOW5SdfWgVLkpSnla9zVtTO6RZtRTLR7
dks/q1sSX/gzel3N3WtWTHOzWkxyFl8dEiPvAinH3BKbRQmHDzIHtEp8t91K
ygFcVVHq6Ql4YdY82J0yDn42MP0/JHabCnUuL7sNQ2WHOB2c4R8ciD7uDVBe
y2IzyFXWPcQ98S+6aqFhsGM4V4eQcMy9


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GuFU9rk4s4tfNSco2u6nLYgk5kVH4r5L/n0qB6dOAIkvGY0Kz93YaR1beRQn
635nnKmup2eapoye6JZxcYOqFY2UeThuRd9Elk3e4WSYWlJaUJLjgAHntKg6
XZ6xvTgHmq0oS+TUnbJ5YLWWsVY9NJCoYg2GHM9z7bMJ/B+zSf4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Hzj5Bel6UCZaSJVircENUBY4ZUXqG//6d+Os7bsfwsRn65e09o2nUJvmdL0e
YJ845RSpdeYn7Ky9J5KgxcBZJ5gkrewwT2NzSiOcDzLQUZvyKIg0b/3tVTPZ
xUTK1wY0zGEjoPjReMg85FtZPnyiW0UjPo5PuZgK5hO90TgQp00=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 129136)
`pragma protect data_block
9Vesi/tTpqyQlaHclYWvSvbYWvn5NW5X2uDD3H2FxDs9KgrXYAI9sGbHIkVQ
7MJkn/8DjvWoHUMiOAKykcIF7q/pcJBY8DfcHdIBf64Nynxr91o0I+7GdXja
QaCUJe86FkHpoT60/ZuYg+xiUbv0vV0PgmhJMZf+Sy8jwAy0JJQ/LTODslEj
GQUxuIAUocQ+8jxrS97rswpQ7jToEtGNpD0X8mXRkF0kE8Ya2NHOwQwm9bTk
PfC9cfTCksazEIj+AHFDByPZXIV4NBKCZZ6p9439H8QAlu7LIfWl7Uuqn8Fs
Q77KNH+PcYhGnM36E1qpDKdLmHAMpmXNTAPK69/46ZUpmI7FLaIJHcrYwotb
2eVxK2PE/goKxA8SM9ek5dzL+pMit+ANWDhYDHWZoGCBP/zi97MNeWOr1pIC
TtOeP8hySUDbVVWQYvSTCj6Qh9KiN8/tzPsF+wMlw+NT3UZHasoYnFbYcLsx
QQF7SJx9+6K8iK2i1hcILw4FggTfsn0asH2fX+PTx4gwjoRUQHMdfVJVuCFY
wc6TSU62O9hmEQQDhkR0kQEOF1Hr2ENLzaFe92YjTcTYvdaVc3Hirhef6S21
2LJ6cHV4n80gvObQJSsq6OFhuhMFtsQSDQmF8w4cqph7dmAF2ZvaiilNe6VU
Ol0IBVbQAK1sGIPFOndyuV7N/ZONnllNMf+3bU77adO0JU0TKTR78v3jzz/e
QoAw5kkjMkJavMSAMdRWBHKeF+LUP5ZJ+K73uF+NDwb/TlnunEenclJ7b2hy
zeAFOV9ckEfwv3mQxqEh78F24dU5vRByhSj2avCLJg4AqcdllyxbryT3GH25
lEp6cAldwrdS+tCiJ0vIloAxib/oEM3CoCx4KJmNg9cznTMwsZEpEM/XdZTn
oy55InNoCEYhMn7rYzbZVYeUo/r7B5XSNXeZQzB7n6OEuLpirJD86JpIdc1l
CXhWM38OTR3FC+Trf6cC8LvwNTg4CweWZZYjGQ1xP5qhjS2b1IenuHodMZ+Q
99a9CDdeYQFn7HpRhL/K0e5JSW0FypKNP1ZjjDGpzvBPuel7kNOkjUHKNpAI
5RmnxFrH7CUc793rvsVsRkpvIJLYWxRySMPmv4fP+CTEVAMhEQWk5t6TFeBq
+154+Qweo48ztjNlkFsM7LfzMvH0pjBHT2Gxfjuc9UMOpnNQ63x/jw6lv+NC
GHqM8vl287DrdaAy/LXcEQk5BltiwNEXP4e+xJxFlXy8y3BdKI4vIUkP+FVn
MZptW3302YEiqtcrbSTuydEQzf7Mz3S8Xwe6Ny+bc3y3hK05WS/il0IUHMVn
U63Wq/U0A1SZKPmdkpc4arv80wxtB324ewGE3K4koldGpqBHYfmEKH/au9pa
y4MSKFIt1zlW8Nvw3FubmQReXHIC5ClAN+hiwPGnSbn7ZQvFrwEAyzpF/3XQ
DxkT6IHy0xD7xF15SR/5oJTHTphsdRL6bnFeHP0ow5uY0/eSpe6+LjSteOj4
/puXm6y/ieyxVzxjABG+i36rrmCgyUi/BwvqnOgkYOw2JzUBXpg0uxqKOykW
Bcgu9kcpO9dq5zmq5fRI8kp2OLUHxNq6sZ2sT5ZJKS9fWfS5E/sXx55C2M/e
srQejEvp/GE8fVtG0OqkIbaQXAP191z0Th8a5upL/rCoLo4RtaIDVX6qmh7b
EklJ3jkYnuG3IS25acvEmen9Qhr06Q1qlyiT0IbZBIM0J7NH8i8YIIvyq7/n
7AmQ5IHpAt+zzuN6OH19dvHqIEzaM7q5M9upcvPTUWBkZU17q9tNXDnjPVS2
0bNfa3Crom2mNcXOiE4ReBSML7ww+bU5rFGVGGsufzzr0+uh9xluqbdeLGsp
MIRQbZBGPP4BHeqdZfoEjW6Qs+mW8DLk9l0a7rj+dFwvF8TTL61f3zHIjCPw
UVNhXvW2koAgGNpEPtq/wOoWPl/ObCigYbMzORxxF5Cid/GCLQXnlOsTHZNM
/ovLSs1hvvQDaFz99I5mG9ulSgpW/Xb84MUCKV+hI1IfgFlh7EKKY/eoOrPM
IYRvsdwXmSiBxQgs19VIXAnohaa2JqF6/W6QidJBeaR1sxxXefze1hPnAOU7
SEmCst9n/Ehe9MsCPnPFWFJtQbaGWJFVqMNWWetuphMv9METalFTssdE6AO1
1WZoRQ+k85L3ojLTEYC1LpCOfv3bckfj3GPJcpwtL3Jc06lJQhVrbE0sPY2O
pArYTTatRirAb8Qufw8Migq/LUB5jld1UhGbdzJ50yS6/1AQR/+mRSXxsHKH
D4N2IGnC2KE1keStzhS15XLuo7pZbxTVcJnBJCSN2+mxe2NvtDFGl9jgelIb
RkDd1b3nD0FXtLC9Cp2PEUqfbILxUYKAysPAXI99MGAYbxxg86PshJkuKypF
VusCd/Z7tiI5aW/9NqTx526aX40D3cPOi6VIPVod635oQD6DGuVv//dVP8gy
/B6pNogoI24dMbf8wsg5CL4xKderFPOedKAd9ZV4MIxaB5lG1L+Ogl9z2zSZ
a8NvSAo/7fc3ij9WUzX6Ww44pHBPdBmmEGTwGT0zoTIo0yKRMo1+jdEhzazZ
+slp0FgMiYbtlihPyXJB2sLQS7kaGec0FqEZ/sZRg/fAF6iLshExDrbSSG7n
9O3U0/vxmgLdLXjTwvo/4nhcRKmJ2gUZ1ukBhX3GpdzjauWcoPUTnsr4qeaV
k5tE+eC11U42g49QFf55Ew2ZQSQqFStQQIJvw2LFB4VVmbyIcQX9EaovvpDa
pHGxxun3RC8ETCEDCnv+rhubjd/OFvZxXszWLpoFutSE3Or97qWLnU80hUhK
osyYlB9bDEWbzJdZN50FYxMbihhLaEkKGkIvLCt+hnhxFxxEIcbyWReQltCF
EVnbr9n18T7EHrjDYS8Wkd2pxWi1RL1BsWm6bpjHlfQvbUbkxOyV45COTPkD
hppVVEHYopvZbh4i0bfTQlzl3315tH4dJkRBYjqnm9zismQaNcbz74fG1fQU
ITE2zI8L8fiVizFGcx80bbduQ1fufFAy8DRMCRO+hZjRkX/I/I4+aEfeKAwY
rDkaWA/1qCnh9p6mQaKMjvvG8iygLB1zawohZptGWG4K1Y4lGs7iYBrxvzC6
FLcKDx6ZWcJkogZN6cVJwdz+LYy2NHeuroRbQzo3rCDX04nkN5Ght8Bvl5HA
ds3tkYCo/yQ9Tn0cp0z3Ez8L9ydkY0kulohI5fYn6IkUZeUAXXnx1LiMHsKK
xEzA8Bx/xg5TaFdFoB1X+Dnm9QxhqAEEBY87xe3CtSOGdJa0DyTVw+XEK3mu
DoLCODe7Js++4SrZiYQ6Ayi0G83tRTRGPrEQI6Ywo/pPUNJE0bcPRjj4wPLk
iJU3MHXZNIo1F/hgUGNc+tRnSqHTS9g9QqW+hSuPt+fUZxJdsmhURx0eemlm
qZDBHnJTcYymOTPff1af6yIoz1BdTeuMKbrgGjWzXU+juaihTwkGnXsnSyPx
3ok6Mw05GRKqq9pgys9gHm1gASStGFvf1XkYkanK3kMvNyq+ETIb+qm8ycHx
+b6Qxtw1btAnVBGHloBJ+L7b41AMmj7HlGAx5ISJbZPRu+XigQu5ZoJvfQND
B1FxBMKhrrbIFNapHd2j8rDuyPQwa52BM7mprZnkHsBfDT9IXs0Pt7/N0qGq
4oS9BOb5HxjJCOMAIwmgIDSEIxU/aqocDgzEGRbTg8Zg9ozVRv+H1YctfkdH
Nf8+SCBWbIPnu9h+GrIPLnssZQH+k0A3fuX6ezW04irvh9AUilpap/TzDpEc
J8eA+epI2xcG1zkAUoxBxyNCcbc1IxHBRrmODB2Xp7Re5DRpk1/MYRrqAOW8
hMXHanNG07k8JATHHDEI8kHM8jZlsbyf+bLFU8NNyJYDXYWIxWzpk+wuZHcL
N0EtGra3bdRKGGPB4rBr2g9Q7K8Kt5vVqXMSKU+za0zJf17jaZloh3wZyR8s
Zs4CdbJcd5EgoY/KcIxFEBvZXueSastFYf4bxuincOewxnE5gbDasbgnWd4O
TrJMh0C9//V37zLZGwci4bJdZrNZWpANzxNUGy/KEZtJP1x+sfyO7GCe+o7o
ruAixN+fiQlTv6RC0Eda93fEFECTQx7NN3JFnOJpWESpF0sY+eGvIvpayhu1
ckACfTay+CSVkqoWvtzUftAxxnEs3G048ZQcUSGvPsuhk21BVthwjIx0REKr
Suv3gbw1nKEsuesG4F52zlpDMuyJHxr2pwX2q4EiD9y2mFFgGe7GEaeh1qT/
FWcjTEwhJBMCN36I6RFVxGivgEv9GelEAzRBDaHE6yHpwX3A+eWfGRSK2hJ1
bJtxboxhzOiLYFxGgZa/v1vM/SoWTGLjwxvxS0hOGpbr1DvhIpCCiuKEMRJj
7kc/2rcZKmFFTTw9Km7ehgKkYaEMDY56LuBM4TS+WSLEYPzlkm+cTeu3a0QH
ACGPes4fE4O+InXwTPJa2ipQe2ofYM47lRGmEGw9D2CXIALqrCTcK4Vq0ESQ
J/trE6TJWP7exdg3GycDZf0sV/AcsRdQuyaF1Z1legedz+hUSHGfAk9ZKUBq
9ya/BP2Rq3//9W3KH2D7uoePxvP+nB+KrjGjn7tlTQ3rTJT/56XUBJTNS3xS
XpHEg7dZZ0AoFAkfNVI0StQmuDNyKjedeKxkne9FXdpnmYmm7nCXy14XENTZ
Xtu7S4yWxEnLrzPClOt2lHDLuoWoFlBsIv1HygEd0u4rQa6siAaDSoQuhYeR
D/mi7f4KngIqtcJkTQ7KJuTWZmzCz7YwrYrGmFvFGh0ibCxSVPgGswbxu1HG
B4RVG0KELQ4wk5gJDmw3aengDsXqrQ/9eY/4emxwKDKc4yX5EG+tXSxosxMV
qopKk+fcQ7WClypE7Q9jopQRLDBxvmoWMOlWa3slP62uldI8KHI4CTwlpTJ5
l5z54eMUdUjfJXwWLpTtnJ8E0sh02mghZ5FE8MDONZdgolenn7dvwk+AdaNY
Y2Qvb3r0eYFh1tuJtLkMPYM/YjZtNOym0QqbcUCSEtwjH+yRf5ZzkWqzN3rR
R09Pu6u26hKQoIFgcPYji5p/+2CTlGqXFvEc8vU377bSOeXGayGh4oj1+igd
aNpxnGFj9ofUQZOFNNOMI+OfuDt3/z5F6r1CjYsEvFNaAn46WVTUo55et3PY
TsFoKIgmAxoxabSd1RTLU5x087sXzaPBqvJJNALNB97MsdqORlWHoOax0wwS
Uy/0bn9JOfmKGxwVLeGkI4non9n5kBc43AUTscWKe+5rIiE8Uz1XwHgCetMn
G8vSvyTjSSF2+iskRtGi1thqP+itKTbQFvWqhi/YfRZ80FCasy3pHsqjxGbE
YFw0h/0rBhUidLa5jcC1MgyCaDi5ZIWVO3iqBW9B7wGxB7yoD5CVsgYrd789
DGAx/Z0TO4LUJ/2l+7lZsMbhSigmvZ+xaU3yqS/WUz4EoWCzCkcniL+mFLG9
mX5TqUhxH2Lh68+RLnY7vlmzvlc9/V+7gLZJxRxW1IlZbHOu8GGiFwnJvdkr
FEQD04+1B52uvMgwgbEgjuwRDjsRlWrcWi54YC4suoixEoFIAX9eY0K7PXsg
RGf1vMffPbOZ8FzkrlJPXIoXkxdaUffainbeWZr2agHHkaTkRL1ecpsMdSe0
WNbfll7LX5RNxkd2lc5DPtCI6qFmikvnKw9E8vbhdmaS3gxuhNOXdFUidrZ7
/x0lDBjX/X3zXg+NyqIowLtlsKl3Q8tpYMJS7px9GiEhLk5CwK6PzFSUqPGe
vhAaOV2r5Kv5n3gE7w0NkRFs0+x9JrfQncuT/f/QHEYgFA8pv0Q7i47QDx5b
mwJOmy8Z6p+NrSVPO5rpWc7mEYnamReG0hE0oXz4yFLINA1YOHP66uca6TuZ
A1QGotXMPKNLYgb0kbxMWRay5kTQe4J1Jm+zdHs0HfTP6qMrivWqQkZQWDSa
JhLyIw0V2oVGFPVHCneHvRHNw3MnQmJMuzxEuFCrLqh+RcdHCs9Xp3mu5JHC
3qFOfSAL7NICzdcM2fHyGATYb4auWhlaWZOWjVxQWnPex73FVcYJ9lNQ7rHL
L4UDuF8V2AyMeLu4dnLwYpcHA1gnVMXB5uCAdxBqjQc3UcNLcilhlOmUYIpG
J5tPtQvMtCb8g17Ie09wuL66WhnUchI7axQoyvpiT0ESR2HN6CMgQpveCnTK
7kic4C7J+O3+8y9YWF90trABbURA512GJyTnn8rhkm6nzBfgUSYTOoOb6vpB
VTckxSKCCzYH7DUNJJe6I1VIEVn42spOJUNj8oowAV3hiqOiFiHPCqjx8Ypu
64XQsMuI0JIfoadiCk67GImRnRdqkE1hGZ/DBjmaP8KbcoQSSRKaY9Vun29W
FB9CYDu8MDoOLV/83Ie93+h3eMYQVp5frmXjBQRhWWajQMp5bblzRRxXcgYH
x61Jpkjv8J7vCGyypzZ1bPEolcqURt7yhgwzhwpWv49wigeBb+YDpl1uvjiC
TOIdTbro9A5zM3AWBaUe5e8gem9eHlUztVDlQ8Wymwp84dKdj5kPrG4HhKTp
DDbUBcpSQSyXFBtO85epLoZ16JzrynKDDTd+HBxJMvReiM5TRlILQ0EuW1hP
+8x7JCIsS+FZbxwe89ieQIPYnUbN2LAfqHlNTfN0jRtmRrbJGaxnPMXGU79G
PGJiVuUvmscAEwuVTlC4/qsmsULaYSBjsn0P2zGHzQUGxumMDYESXsAAoVlR
3ZApEtOz/u5NrK2Y4nWvTq6BdRL7rp+I5iH5yb6/33BsM+EYkdvxUuA1K0Oe
wDmBIZpMMDeR+a/CjqMecMBarVrjZ/oeDCYRAXFnXiEqpZjTC6Ae0AcEoZHB
4e7ab1aM2eE9JCiCxpu3DUGmebM1HfjYUJilZUhlHzr0yms9Xh4YO9Yy5Qkw
/5qwvZDTx5CbtxGxFnqBqCfXcuXYvDCKyEBBFkgKuUYjRaDqcyGJE2rCorj8
KBLWTwJPuT96U6hPcmQdHWQLsguI9RLim2cO1mk7rkKnB9p/6ri9tI4gMZJM
iX/JhxEvwythAa4Gh6dRxr1sLGFISbXgY26vmZ/VsFhvub+fqzYk81sj+wiT
mb2V8N3yPcmxFnlpkBexm9ubXM2yg0AMjBwaGyMF7nMWHDQMkvDzY1iDw6Ph
kh0/K5ZUEYgbWkueCtmOg0Z9HhmQevFvzMG9Pd3plUMS3reiWfp5KO0EYkCK
1BfulIMKgIpxFitkUdn4b0+0iRVeOm2c6+wl0gadvzSBosKjghSBT+e7/udS
5i0UdqDBvSCN4ckyRYXE/4aJxWyslVggYflTfODZ26gUsqOUwoSGjZZlO3UN
5p7ikrYTgV06HCuDIlib8S+JpN5EEkJZtgfWIJCxTcfrqanI6etDCwpa713O
EQaEtfvJw6gdbVG3U0tjOotBctpCGn9bCQWeBGHBU36C3LURFCgwfCp/rsbm
ZQy5g4TmzBWLS4m1DJ+9jJj3PxW4f/uivEKy7tJaEdwb+jBGpdvxJJaaas8c
9gE8Ap93FA4C2ud4U7P2jcCh47aah9tXKk0Lyx7hMEUo3betsj2JROy3yZ7I
DjiQoS2Dtn+P1Rtn7tm5083v0h4W1WWJ8jNiYyeD8uHB8ZSW7vDcMUngabDv
8AgP/N8kPKhNmhLkgz3aumPpMzN6oywqI1wFO153LZOTNKGDt2g2o3ejeiGq
FzTlxke7yBoqAZoahDGdRRVxFeAk3+QRstwoQPO4fqXHmiNfXoBXyL4i8zvU
XNrjZp8kN01MjzTDD5jInMgUmjwyn6MZEn09I9yosjoarGHmd16qy3v51NuM
/Uas73bKUbBm1jxF4WsEXLS3F93VTVvLZo8xBw7R0XpUgLXVHa3lOniwaAGs
sV90Mz0FnuTSjlQAa9mmP8u7l8ydprFsyBob5lXMrmro9jkr8egIKkSMPN7J
H45g4C6k04Fu81OwTdGKVUIOHs6hwRwLeWdleyZFYCLpX1k1dVvb2f7cGInd
mD5Lgn0GMg1RUA4ogyCscDNSXmRtoBQJxrfJZipJvkV9ci18ygomgoX4Bqxq
1kVapaxYifgoU5wNnKxGwEXKFeD0DciDmDAfY6o6O76YzxDbaJ2UiLH1mI3P
AgeHaBoYKpsE3Vsi3dHqrqwf7KFh836XHHIwR8mOCmG1r4X+9fZriYRR2Zr1
seLS/SRVoZVcgTfJHUrQIHX/qLOKwi0mIdfUX1bQ4XzdCm6y9DbhXYunx4OV
gE7O7KtEYnckXac2iFQ+4KKRoj0tewVwOrqKVO5gKRFrcwvcLZYQxZGRrtJw
q5Zg5Dv98YSNnlFUudRIVRwDHIZrhUZWnUm9+guvK3lJxJwxBEZhHLm2OfR1
5LwBO1PSFDeF6yBdGHkCaDQDa9AJf5as6/rVeFME5LJrNwWs6xxz0lbpGi6p
KzRakby9QkUlWIPJXmnEUI4nVnTeFv00BTQ69DtZ1BXse7feXdp1+9EN27Wa
2uXtW6NSaXkuKz/A7b6mz4ZUw370+YNrcpJKxZ3QdM7paSZf3ToOF2Hxi3kt
6vzoKK8qGoeyqrNonk15B2HY7kyYc0mEYk1saaheEBKlA/kvchs5jsNibBLO
NlphTc+tK09/dVla4538IegNPYnp2TMQi1yrrXkjW6mYgpyY8YuDIObvac+d
YX5kvz+VNmgw8s/82Y8IJ0q0xAhlJEtix1YR2nRhEp+UQQHQxuqCk01Nuf0U
Z1NHt0LYZyRxnw9AQDhjfivqs5jE2f4J1giuR5y9PPXVgxuhxEPXDh8gIief
7oVsDD3B7arS2i9e975LjjfK3I7C5ekLs5LaqvJIBR5X35kjf0hlRfD7wqsq
Y9H1pD39VQGoAwmw9YbD35UHgaH5MuRPI3FQsp8TD9iWVn0SK/VHq4cSJs9s
qOZl9Jrx7FLDW8Vp4S3s2PlcjVbEIOm6dHo4aYLXfnbcf4ZR24qR30rARfMj
QpuciPqSBNXvECIATKC44oI9GulY3Xi8qwocyD+WXVY5E+182lDSUn4jMwHC
CH8FV1dhuCO//T2F17uHLtDt7iQy1TEuyznEiQvnamGGze+bWoKYVFxESPja
JJNE10UWwjHwy80rqaD5PwjZZl+AKrNpKIILCj5rBgijJ8HbFRrDqFe8KNyK
dKaS4ImIpjc5Ul0o3RjhU7V7FokM6QgSDu1rMqUEmTj1enpXHSsCBYKJg3zS
pgZMFKgeGpNbOkC+Ws+MVzSEztZdQsPHsNnP863Oa5ZY20MicoIEUMvpeMc8
WfRavkti6ZL3N+SWV0orWPJJ5sDHsLJDiwvr6OnWq4vRDmqoKymBsQO/bkn6
jhPflP2hO+D9MB9yRu7OSKNqDCKYqEF63epxxSx4DBJTlxnBWE2XK7mwTbUb
+UVwrnOJfHf0VfqzeMc2cKj8eUv0O/keI4DsskEJBN2hLB2/B53kNFU7+brI
n3YG6pU6Ocx5nPDnS52gJ6rmy5RmOQEsxTTj75Q+MMBQYzGqQG1DZ0HrcFv0
CpXbDltWIBaXucpNIH1bh0jqMCIa94DWO7eAy0ZsnmlVGniS1M3iaxYSR0xo
1D6FZ7YUUIgRaH3uu/llz4Xhfv6RBD392IIoMDLQV1A4ydkzOjiWENxA5Zne
pi0kIi7PAhzYxctTyrrdaJ1aONg2bf1+/Fv6enDLZbWzH64d90k3SqlD1eGT
OfUOTTCHAA+1mkOJGAT6ScErM3dc3K4rbPRpTyzEhvBcGrHg1OizBhs5/NDo
LGhJaUK0OJFOjLe4pl7qod51h4rdelOXyZdI1Fwe573A+KJ8rrWFAumV1mN1
sr1P9QJkzyqHfWDpb4z78iqzcmPoVsIBruwJpNODNtbnqFobqzgIwd6yX/Yf
jxwZV87T5C824SebX1OhImnCjUbDGfuvKnKiXhH0yZeMT9TuQTssKO3kHDaK
+OB88M/Pirf3nLsWGaimdWwbFYwU3N7YckSEVo9oAgvQWgIxtdmURAuOohB0
ZX0/wmdSui741f+aqukei/X7CL7g2WYvmXnSEPs4TBXQgP5PKzHhLfwesrtb
Z1IJsEaNY2S23FKbqYyo6JL/jxZFZB6KItxiN7SWkw4Irng4ihWJkQrQ06rX
TgW3L3qKjIli+qTQwygWcivZ5AKPr8MJqfOrtcHePD0LR4E4F1BIk8vHi9sf
ZF1Vg/o0oahxETXJpEUalejbzdPJR4O+lzCYnBzOafd9gFhFQqwTFpG+D8th
GxfK5xc+kA+K76sqFOzaZtXxLVprjNEeG2x4aM2910MCS5YnhJdnhqvRgUMA
JnSy63GGFpClNxe40b3Po8byfekX7KSC9zpXGb2vH4M6s+AEeSnfnZW61MRy
IEhE3qlFF3AUCSj2DLDV9SP0lgeMSvHMFBOMkhTTF+gfM+mOoH6oXsxwWmbL
aHrxm4dR065neOgzmqD7NCu6nXERm/7Qu6st54/0bozTgFZ268Yc9UgfxZMr
2UVmPppkH9JFh2hoRwG2fPP5g7uWiHQIAeMVCf+N0NYA2XzssrWEXAfLU8ID
mtgYCU5HKHwf/V5AdyNbUuiDv2sddZeX/JntB4oFVBQxBajvdooc65RoWiBa
/OOp78zIQc0iYqBG06IUPlQ5saV88b6vspWtHs5AN4htXFe9eOrS5wqcdJSh
f7oNCEmBqkyu8Wb3JAfGfUNcHJ+z/W++5rk/6nSFZSvt9Z/eXrq2S9VmdZi5
+Lc2bg6WegNRqgUVr/kjHpGxWKfAuIodOfcYItkJv6VrI6mHFs2FPtGwdlZ9
pu6xqrd1DTXpMonD/7WwMjKJPxOQ1/41VX0Ssl1iV4ykPHFowSClyihncXmh
PqjLAkfyRoVJiy962xFc1XHP6DWgkFPSlIEuF9LVMUc8fB/xueIOT/oGkL0l
dhZhi01vWwPJQeVRC5nNpdofkkyuGmLK18gDGzmCen2Cxbt9E10rXrvIQiVO
Vn/36X24PhDBJqMMVEu9C94hhoGxNpymA+eR0fuz4i7GdTktfAIy85jnVzLp
hqXkLmYxRz5QyMWtNjD6UIMiRsyjtm/3w1HaCSQEeZIZntVzrUXW5nyjVlZJ
34vSUX2ILR9iZEPnmLk1x6JWs7LYQJPL1xlxtPp54PswHtLR9fh+RhixqF/T
+lBpisvAhGxU9lLyzAS9Im13eCL+b8e2DNK7AOhHrcXnmuA8yt+4/3j6z3JD
aMIyAU6X9AKzsb4fdEooKX9gKcAWBss+i28ekiKyE7IOROK3TsZYFSS8aIy9
yR7xyU9fnZx9BGq6O5Y2Cpvx4yyADPbQjN1XHR89rElRL3hrAWDo2DkgrEbD
tcHmrhWWoz+GkrVw2IBIbYi3mead4j8+hCvS8wQp/4JhYz5g0mGYoHdxpWqs
dnZrCCkn9UGNgAF0ON/heWERxYvs3ns3zEIjuS3F55xSjXROqkP5Mou7NxZY
bASiP9wybYbQOV6d+JBdmlcZucIWjCUrEawpx9UIUD548Mwp7VFoHhUXsqEf
1Th7syuTP8QusNztbeZs3i7LCdslHyNm+32G+IzyGPezfENO6nfs/TvDOU71
jhZPk5upOFLFNPOo17ybBdWi7l6M0BRBVGoAsAE/9NbVwAHDNBUosdR255za
zcjJE6ViR5KrfZlmArqXHzdQXzCue3Rbgbiee7vB+gzJa28+gbO6jfXBRWI2
QMmFogsF7LBCUUJT3oBN7qvI2udv2PyM7ns+wGQc59G+A09vF0jr4FlGM0MO
OcrUpPebZZ338BpuUznRL/34QoXU35wOY7xUzWqXBZ8fa2V9Lewz0bf9+AmE
fLMrBjSJUJOnanSo3ppEiq+jJCQ/6MWIO/6QsHm50kGRSgkPD80pHGHhCHz4
Rz2tChciqxkSGIQo6Dntbm5rZ8ssvLrylcJfbov1umPKVyu5M8p6wn4vozk5
fPmFCx4nL3/XvJOW0Xqur0fo63O2dzvPpozP7TgQY76lVH1cNUdlYagGywcf
HEhFuV39eT+/6Q2M8/nebk4YzN31bK40P7OwVzHxtbmqM9yl8X6TaVDzyrJ3
zAHVQqZT5v7h6eBKF0DqW7XTNjy7UzNyYbzsj8P9OGa1onab8gULQxefVkvb
efANA444oBudE8xRn9JhaMpBnZXw9UbpeTz6dbdqTKHo6DowN8UIRSWBYmtB
On6F8OngtVJlfnSXiVxoLpbov1QZxtP9YoyQT3/4V4BIzrBSKKPj5gIaJ6Sm
VPmiASYpwAp19YAR/Sh3rAAsZdusPq+xwcBUzH9+nW4KfZ5yJL9Rpf7EaCe6
nNzEFQJm6ATbL3ExUpicuSEfZpXwmZh58ETKOp9CDEGJ+aMoL56ppuTrllDO
Gm5YwKTnksrfR90OaOAT59s6nh6Ok1dBp2ozQTp/wJMlV6o0++VKkL91BjyU
oI/RSxUHdpAdgaMysxFIqAYsbI421veREwqDaEPmE6PZ/KaRSLnj1ifWOCyh
9GheGTw+4pxU0z2ehG6Y8L4fK0RwivCg+E3YMyP0Xr6bjSSCmbj6zSLdBATH
g+5WQ8OpDmHG3Rt63UqMzZAhJEw8GQolAKoeRaqH/9p3wCoZ+v36O5iP8Obk
SACK7KPyMZchtD9bKvwhI/FDqO6W042uwaF3U74UNypLoxfSjg6t+CYkNOGh
zOWuVo4OHCpn+g1ATtPK18N0s+37LX+8t6DsvHGjmoBgr+ur8CW1rdxptqXf
JCmbXor/YlKDOHhKW6T4o0fNVd+PPEHU5UGGQBGQaJNAXdsF905AWa/j3ZBj
hhjOiiZ1p3mhFsxMBxjI/OK2cuGNykZ1lwzg9+5f4TZm149KzZ66OzEjwc7t
oGWR4DFtkoUuzpI5yPGrHJ0hXfTK0lnLH/SdNViao9537MvBcfpq9FA1eLMA
+ARR62MiQyhtUBwiREHyTBWKKzlNk1CCjXU19dxb+PDYMPJYlBYEJoiSF1MU
Nu4ghkDavEyu68Ck5ftA7eA+0CFsszibN4QEUEEH3B6iAr7k7vS9q8LvdDUE
stRsL4N68U1qTPeQ+DROqmm3ox6WGvwQbQ8YuUcMCYnMEkw5CeBAxndsQjUh
qzYFU0ChfIg37PKrUyM+xYYiqZvf53RcEDJJSYsWgg3Mt+0N4MVLDxAb/dgo
xhw1BxYMmkiyDhVXhYHAIdQ1hOrE91SeBRTvPBkhneJCBql69GMYsO82f6Qu
s1Hh3qIrj+bwrXiOSVRv6VHGr5A4MI8qqDhp4+ecZBOJsZi9oQCj1Gus1ebd
7ZejdaFYnJIzjsPHB6rG1Ky+1+qI8TxmHc1R6b+YRKWs8b7DpYCiYV8Kz6fs
f5Pkx3mAyC1s359bjoC3NlpgapFbi9A1d5DlEQuVWlixFa7d6U6XiGY5EPI1
EfNWFg6dLJvXB92v40AdhLeKO+FO4KY9iLmiCyS6Sbzksl/MmNc4Zk5siCK7
vYSN5J6Jb6doHumFwXdviaaOJ2OL2CENDY8fSzsHnNGZu4iey+3i99eQcd7B
ZFQMZFS28f646Atmud2rXvN0wJry9TB/GJcxMG6hxlbFlYKdvGzGtHOKBANS
ZqfYWYN7+QTJJoD506KaXISICnzPMcbXXH9x8YbFjvkRcby+ougt3xLrlZBr
+vD57EqLvhlEMdgFGynhRH6fcS8D0OHyrJFnUgvRHff8t7C2BSNpyG9+shgK
JjDjwPsQZ861hxGHOkX9x2aT1X+uDcbtH9SvQ1NWXpKqiz8wZZI0wg7Tnipm
Lisn75aCY5VYLuNk12S2nzTu//bpRbSOB4R99hgG2pgD2aeyLz8QgYSkfXTx
sEAVvca8BY1yxF80YdDQ12hIIWKx29r9OtKrG0UwvhPevjjgaC3/ripKDznV
O5s8mZULwN1sfizEKnipIJjBgx4Eh55th2LX6jiVOk0r+sUAYrWSg4OegCB3
COxupCmkxCA+NtYT1l62CeLPy+DcSXft1jxooqvQFk38bYK/0HaCfAtmUcYD
lvtwk8bSvYsr0KgbvhbhKZSysNWC1b2LdIwFe4y0w6OHlH5OfaX/eUS0nv4L
crz4/wgNKf1y9jhOsFSza6JkRudIY0cVIeYnt+JS2Fpamjo1cLyUMZDciXHU
dwKHqCMPPIBsPGHbxW2U9+8N5iNiizYM2nM48q7WClJJEUaajg8PcnLTyNsi
Y8oqx120Z0af0gg+wkHKzPzdfcVomX7QHmwKEJKEJswj772YrybHkGbJnCRI
SdMPYJ/YvgAagliRFbDSSuW5Bf29ApON7KGneXk2yqjxlIRuxL6qzlmnZdR9
RA00afyQsodm0C0YwY57btDOdKCW32830B6wbc+0SrD8K0iTPDDPOX7F4DWP
aWStewoC7qEwaw5YhjkCi4WQjAZYf6L1Ja/Y0aIbVog74wSGR37g8hm+X3rb
mBm3a61hdLKkkjw5vDEh48BQ5XMoXKnKo/4XwKWORjq8PRrGt2tfU7lNcuHE
E1Z0qQ+tZUDFYkpYuK0yoMez8fxsC6lOwcXYf1NxZB84PE9dZYuuqLo9MX9f
oCT72lXqR2wb61Q0stxIERkvSPeSRpeSbtT7fMXQ6HeZGpIe0WJGgfo4wVol
lhmxb5w5PeehsaYYcuq0CeKhK3oAubZBJa8e9oBZ4dBpVZqsT1zAVEShCklP
q8ZP99R17ZjL1NF7ow4AqYTskx9SvedxN9rL62V4+S4NOyCR6aZPKPdIC8L8
H7c4uEU7nOLGXnpVluLk4mMODulzOJxPZ/aTZZz6v34MwfUWrFwXRV0B9jfr
888Dv9cYnABIz3iUZAcjbiRS/fFXHqRqXfhCl1l4r2I57Vb1FdpfFMIGBLkM
dJf+3HKfUvwd/1ehXyaJO1s9tSd0O1H5jZ0Dkhm7oFI60jSXZROxd1ZpNK4A
Px36QIvCdowdEh1/onglBMzWaeg7wP8qi+weH+Hj8YGDOSeWPhTBZ7dttxPk
Z7cR4XUcD0oc9pXz6Aa4wYuARFNfVjaURmAbcqTzHKAAUZ2/ytZvsV8QnOsP
C2XF4Gch2wu+BkL2praAjkhcgYnhMPw/rWois0zkMLwiZeR47xfI+jlyctqV
XNgmWwW5CwkfOVJUlO9zp80mgiEY0zN3p9n9hEV25c44s8bQxrCGRvmEJNxm
JVzUVR+XIvr6Q8giDt+Rsq1rapHYc75fNQpSkrjm6f0h4OOfbwpA7nOFvXSI
UbhiJX9DB+hmJVJbT/J2dcd/qqhFi3uzyp1507+6dPxM7ZSkj4V9RM6sB7ur
ahJOJu8WxtUcXoG2z2Bu46LXbmLceogEylBW6pLYzKIeWT7xpYid98DWmFGN
W6lRPJ8Z90SCCjK788ZWpQtu4/X8fvNXajnZ3pHLZI6ZHeVFXwa4KpmaYJ13
zCL2aiwfMalB3O2o8EmZdrX1Eo77w+xezm8+FgZsnZVOGatH6aC6VkdBY19o
gck9ml2PY4WvD1IbHFZFCrseJCW52hxULFl03DaAOM4TGvl6CYEKqe8K4E1D
R3A9Iznq16QWH0g5LkpUp28DRDSrmGjSwvtRN87RD0JCAkqS0Xa/8A8uNYcx
eaWFibAAw5dlMgpq17FTb+qpJwNvZrQkCU5NuYmxoITqRlXc0b82uWlfCnyG
HUiixYKNzGro9qi5mgzeS5hS3izqOMwxXO5oRdQUE0nLK9/Th+z1M+kPFYb/
btMsoJwumc9ooUbcERfY7h8ZqjDZT2z28cOTcfxZk6VClfoj9Djnz7S5W+Z+
olfVDly+F5T1j9YgAFD/AOJpviYFZX4aoBhoXrV2JgF5B1sgAaTXHDjzIYM/
/kaYWqxJrnk/1Mkg8BRccZnfmvrmwBj81A9Ew/OI0v0SdXyjvHfPCNzxFODv
Nt90REeHK+2Lnp3B23rvGZg/eo6BFzV4Vg7FbAsKUD7TTZIFCELIdytrkawM
P2iqe2oOgG+hdNSMAw6JD+kxdV8TNpSYFcJlFQWseKZME9KKWb9XyZ559tlV
mF7ZCUJo5czVH1EWGfIpMusdju0xFp3PHB35GMpTlnNWRT1hQHdb/YCVWsGZ
xkt6BkjrO4+nLOr0loH3LgNlFxHD0KvbAyyRPh9wCb+dmpB2FrcdsrpXb1kP
M6t7Mm/PZGWTNTfLdspZn+FYvFXsFFwz4gToHRF8kVnoX9R+YyyX3wJhFlNV
ppezRu9TrSInTj/ytv/e0C5urv++Dbon6EN8wOIdP2oJ16G7UPBZuX8nxK1v
82sDVME2sL0qMUt64JlBgqjHSWcK1TkyF3INBwijteaIJrOEPh1cYpAkV3u/
7zKi0YzWB1MFNkI5e24ug/s2kXebH/w7TjKxOSpx34CONAg4w0xXBT4mklPV
PHxfBeY3FraiGcmlI6DzSbFCF1F2+DjQrhKjlvN9HRjQQHjR5Kt/X+sWqLzO
rfOZwPwX6BMbqINYzDpC4Fan1/bydQfAmMCUvFhs6V8RgZ1kKozPQt77Ic/h
qMBwVDMnUqqbvehxCXcXeqb17lUXWalflzYeU+K75cwU0ZnIBs4RBuErMRhs
qPOiwTKZjogmub1vIX/OZPPjRUb786DqulawZ8s7SqWeidLgKg5QrUBeeB7A
xho1wU6fgBw75767jD4oYH6652gY+McFevtqNRri0OAjOh5B+2DzgHBXP7Zm
qtWggUuE0s9mqW7gZCMxnd4eakgkPNkoPNPJt8nLjJifme2Bss319qngvg+0
qlzdrCpuBj6kFxe/W8kAQNGhuxMWg3l1p7xl/xpBbKuUEUHMF5ZDP4TpXStP
i7PXcck7YuLA+uhCJGZAM28Uahe337lfBsfj8MiOx06VgZjOTE8fC+J+iEMp
jbwo5H64PjIA6oIIOX0n9jE78xvVFcvKbbIYbXPDAitvTJf6swq+Fl4ELGM9
JIGH52iqTvbJR1l9j8+NqdQAHJ6in83hhx9tsr0LjxkkQxotiUdZkBtWvkc8
gfB4q/mzAvvIPGXE95xS0u3MgE4dXoBjPGHNzzmH0Pi7oeB4V4jNEePTYXb8
eX1ByojwCZhaXulLEKYy4jnYif0DWDvkakDRhxfOA5eP58hWMQrtREox9vNs
aFa3IWtKAa04ipQHCQQsr3b5WLf4PdBCyhE7ysbb4sGPZXBJq2WkA08ebxpJ
6OuGWgGnQK+LCvBibro15Es9f/R1ygIQ5BxP9gyZFiGQLkUXCSvUlhtpdDpu
ZDgbAkqB6YZpvgcLTuAOoV1x/nmV4jQjeCnXLTwNyOPnMhiu7FnuZ9LPT2ww
7GfqWGK2OeTUbC1HAlcZKdoDYLKZ5zs9JHHGLbr4HZ34Lma9hCCIV8MCdGRK
7/3wGQNvEh/kQ4SYxiM6fbz5e16j/AtbgNSatVc1074caK7BNFmV2PxHuMsy
HzVFmCR0WaYtXr7E+qaKQq1wxrRH7qc3HkLeHQuKxMlMAyLPEwTN9Y2Xvo5Y
ZmgbhL0lKhReCUSSujGn+YrOvB2QJbr8F7Z+brBMpmmEeaAaBHsFR+4BTkmW
myZUTuBUvpAmdwM014LfJPnzflXq70uWtfETD7Ibr6losGLDunrhEtqBdwKp
JLlrTP4LlbqmIrRPyhF7qcLXLU/jXCDceTX9eEKTyYwUhe8ugq0DWYVuQ0nl
UqWj1z44tYzsIJWG2NBRAcnMfiZK+IbLNWeH6VeeaNnR/QbksSu22rIiJqOh
bUqVj2g4AwnBGjrRiJkY3Iwga4wScJO7WHKgLPW8Wp6dEleeeQl48j8H/nDT
5FEQRzJZc/K3qqHgkB2N/L+7ZwkOVKdKQ95J4XST+tEH87/DLKsBDa3XdW9j
1dauDigIKTou0Q3Xh3ADv8jb8Exe0OfeQljdTZs/NaY7G58yQZSyympYKFO+
HgBQFYwoNOY24YJF+RBU2Ihylqqd7uRTx1CSF+E+5OaZcNXZ1ptp2OOxT0Hc
YL71Jpm3vLgZ3WB7KHnWb1yLXdQm215pvWSf1mcTkuXS2k7ul04Q93b/gzWW
gIhgvF6SzSBglsfpQv4Bnf0Vs0rBR0es3iR137w9LZItbKbHB+96/v6zALxw
s4a/LXXdrRk9s6A1Hp2BycesnmrXMiUSSuv9zQPwPCjaPp3g3ES+NTekXKQ2
d2dhyI94yyZHJjOYzFSbx0gDFgz3MjCGoh16++YgRx5SEkX8gNdETsvbtoYv
Os9eHj7GoSf8xkVBlefM4v2csYk+zR6IyqbcyT06EgVQWl8BEieSJWDMfl6k
aghoKHtpMfdxfNZ4u4SSnPASI/cCINmZEj/DyhRR1tjoLnECykBAaGWoLJN0
nHs4iqh6bPMsklyHQOjw2trG9MrHpZcViaBYMPkNOA2+PeynFuztp0tI4XZj
7VoxSgyoyfn5jQyEYRb6TznH3xXuGtGmGp+tE1r+DtHZih2NX44SIZ8G4Pap
wFUtNsckHX7qL28RNfIUh/Mg3y2rmFNYUbK3c8EpuPE09i3ztH2X5rZW/E5m
4N29ZPWpS99tZetnVgXjw1FlJSEPnRJPU/L0TvF1Kwb4wCcDCtb+efCIEce5
A0AthjBWlg0KHriiEPhH/UUcBsWWbr4iK/RJqeLKOk/7PU8Isir9J5Yr1b00
vrX41vpxjw+B94/aw2V1fZgz9BSuNdY3S0DmLKotCZktYasnUvcUEUfN05Wk
PAG6gxIPzCLgQLuMD5oIoO56lNUKWbeRql4ft811ljUM0IJobIklZICTd5nR
rsj9F5xdabYrKehwUn4GZPllnLtz+z2muelNOQf0diZsFb+A3Up75CC/3et9
1g2kCEQCrxUAd7ldchpV48A7Yx4Q7Ed6oiaqvQixsVMP4hpcmeO8agMI4Lk5
oQg3TIZ+Tc5t2bfO9trrUl4C0c5YsGH/n8y6UJoHC1nu3qbLTPTQHocLe63K
ALpgP3zFFH41pqvkDDLpApMlrEnvyTI1fMuVueLaF9+lk150EgNdzI0S1PSc
zxsInqkTIStNYI/TWChFWjO57JQE/CRNCAInIxlxjKlCTPQKLGXWtb7uFgwy
U2/CQFDf7I52U3+d1MoNloH0bMveJvwrOOkGLQn+xTgTVhRCzRUydSpFoPGi
LM9P4OwouZJMdWy37geYxt4/5N2gLQpOZ9Bt6fG7WweJo5yKOf5p+yVkQIMa
gNhvWgTdzGANAzPepinwq+yuVJ6x7ON9qh00ye5Uw1OnAdRp6/eLetg7dcxC
gASxqZMJTyBd/iW5m/HUNqFJodFUMShmw6n1UQWOKZsKpihyU4Lj7dKoxVkr
zDw0iOP5l0Yi263mszorh/O9vi2vimnykKsn6lvQtsbI41G0npDki3dJEhpI
ldREpaUgJNOHT77ghAgpJB759ZrZRMzqIkc+E1KZp0/mGMVrkc1jvZp6NkgS
RT5dKeEXhXNU6lAXWHMH8XVH+3bTPKaMcEjPDgUagXLcgKF5XDwtnkzbVZwW
V3k8iukuRFXFRuuRERx+XXSKDit7VzzzhBp2q5LXQ9ngIIaV/tiOJ/31YIwd
2a0czVSJ43kWNKhiV07avCnJ/o/fWF+6ZiAe9ZKLOQzK6LeHr0andaoerEIg
FDSEyWr0Ak+7ns/1raSthRbzs2C9PFzxCJGlbIeVRmRd6jtyjfYykaHK60ZH
pBIOM3mnlFMea+54oqucQeQPgwP1rOk/zXkA+9+Xwxg5Fwl6YpUj9JIwz0Ok
cnfQVaLoy37MvjXmND10wo7MIE9v5+EWv9LFc1IPXE8pklE86G7v8Hk/ul3L
HflsZZGzFjfayRyIHNhroPk6DWlnPP0LIr4YzFPt4jFaDqS3lKOnlKSbf5L7
UA18quXWaGE0cm9LaFf7lH3C9mjJOxumexiMFzaucZ6l+H+PBb9jUTJFSQm/
7jrVG0sjeCNt4hH2gfgnVwRtYAkxQEgvoy0TS4wAppyc9dMjRCf8NgcmAFpb
3jCadFEY5sBpbfPAE3NyMtUMUeJPBb5pHQMrU10WQeY2SJ4RcyDrYY/9KumC
XLxRHbsaURJaJpk+kTErxFdW81Di2+NMFhZZNkTEKzH5P5rOBx2aKcYd80wO
Bjar6GLFJefE61JEhdb+KmYfeGCrkpX7gTGFG1yu+lJzisqeZpYR2v5KhNDK
sSKUL8TAJpB+SulCLAgmJrZNyG1yv0x6Bce7tOWyi0Zgj8+2eQsvPcsqoscV
FnQv5Y3BzASV8C/+41+6PxVk3e7InVCIofYTG7GFAmONSEWn7W2s4EW5NgVi
kP5FqARGQgy4K0oegFPTupaR65gkPonZxou0ehLhQpMgmIE57Cg0i2n8o5fP
Fr8zByhfbwzYxZwUlk9TQffgDPjr1aekb8SLbWrfbVP9KCTqzuGQ7BwnE9n+
7033UVHzGMo4gPPSaKyOgPEWyCE+spo1BZORaLuN9RohLxC0roWk050MuB0b
5XhYH5SkLZkASjiUAmEKlMXX+mDC4vLDOCISVqeWSEE6hDexbw+S1Esr3pGG
X5H9YESBIJHcQ936UJwYArNJwKTr5Vkqmvx/p0LlgBFC7napR4Oob0UZoTnK
0xSQny/inKgD5OtajNkCpE0eNmcnSRDsxcQYpv+ZpKzOWReWUiRu1SiEB8CK
UN/LF2bhvjz4EonFlk+DuBdo5TV9Al9R7BH/PmQ+qfhvjhkKLf5bLtnfBoPk
p5uAk/2f3VfCbTUMK5Dn5YXoxxRyjqc0sOOS9jFHBAVy3dB6Rctpr2nUmTo6
EszvIB6VvL3tbuKYjRU4jt7OM1owgZ1QxOauqpvRIfUF0qHmMJkC9M/orGm4
1ZGXpFRayAB4xw2MIV8LvF8Sr5Ozv2POofST0bLqVwzR4jgWnUkato9i6Ve0
9om6FdjsTk/KWE3p6e5KaYXUTMg/sJKXei53sLnbsTwtgi7bEKUMUq8FgrwU
n0b+NaGprlJjOnvSt7RqjEPJsT7v5jCad4sjPRNK+RbxOTkhZDJ8C/vZBL7s
4H57AfrEXiCRtl1OTOj0dzCOsMT31ifANN2hI81Dli3vbBtgqfLqypMYNTUl
FqiEaEdWC3OrwQgKUte7rUgj9UAPVSGrBKwscvdSF7ZlD0rE60FQVE920f6L
7E3dimTlj6Fw1E7z4v+MWvz1gIsBifKFQkO+IQPmXcSq/pgg/Q2O97NIrFgs
Nbrb10at3Z+g+8Fa5Ct0aLCX1IYqswbW891ZGhtIuhJsP2LRoniKeWh3jWzN
dJolClMrXTj1TIziRt6IiSqFuVuQmKnPzA6XiYpCvCFm7+oyjb0LGsuOllSB
q4Phg4OlX9GAjVIc/joKjus7lGplxnrYeJSrmQdCuwGSyIv5T6gFvW8Pkwpf
dnWqm8K8HGnlUxu6LOeQQzb+OUa8+qyxvRZa3uRG9k+DErTDrGUM7xpyozSx
fKYt2UA1sMP5qM6bgLM5/yV5SAo0rkbDzUAnkAuv9at1swbbaREHIgImUoBa
T13ofuGqg2XxgulRGp3D/5BGgV+y8KHo62jvday/hPi6WWd0BV60vA8Hq8fJ
5mmhcy0engyMyhbtQf4G2VPqCDcQ7/HKH4HJQ29ejqAGFPSpDR6f1olrb8KJ
k7AaBFlo7R8oTidmXiadH0t9eACa9dvPI7jsdYy+QNRngYOvgoHhlCM2nUdl
mpP6dG750OUEa3X1RoHpZxmoeGFgxx52RVbVz/aT+Sufq9IaNUlcNKrAaQjK
CE85ckq5B9wnQccAvv85QUVcJo7LRceV382SUzIzkz3W3diFMWUJsaNU+Wr7
1bll0rMW0PjzfDQ+jyDQUxkBGnp0bzRmUbbw/N4KubbmSw5ZDoC79D8iflI/
lkPAHap9NA/TfIbJtat4lF+3WVqtuXeyhYXE27ZCn5ybguo5os7OqKyjMqzh
kVWeuGBOloRle51azBdlBo3N2CNP4wODYkWpRbM+HCbchC2NGfs1hjKuHa2z
HovJ0pbhs3nuaeU0FUwgAn7RA0dSprx8KOOJvYMZPt05RyIA2a+Ohl0U1IBN
KpAZui0wx6l4ShJ8ayIh2yfXjC7mEVzagDY6/dQ4U7LB5BVJuQRZknuh961p
OsD2tltfcu4Qn74Aj4neGtWPBpV25qzoEJUnvaLlyBDuybZ3JJgEA1M4Qtkz
pxQApPtOQotVpmEHu7ISLW6/hth6r6GY20+hzuGBasAHdiFD3B56zn+/lYCv
Uy0U6oF71btm6qta/vbM2t8Af1BCxYAkz/jcnbgUD0BECH9tNHUJpvCBfTPr
ew0EZ2uSZX5pu0/cNGGMW/GmIMg1qyA0ZbZX088ERhWdWZIygNqL4fHsPgEC
/lLu3I2BFOFxENdF3DsR7cx91kgASlFGTertXWporMFgo3N4RxslDV1H+HjM
I3v2kyxZL0Lg+2Vg8kMVK776L/CPR6HhaWCToufky2sw8iOqFxFSm+1VuM6f
Q7ksHq7iJilsbTbgYIr7HbY/BqWEr9fq6afe1Tnsxr4yznCzDKSKth0tGo9L
7omxzC+Wkfr0qTywVROkjheVJopYLj1V6ySwj6eZMpNr0Z5xzqtUuBcgrNy8
m/9b9yCw9G0BdTjod7OL62DN6oYcmaldAu7I/3ZZy9KxeIBP2a0Ct8OiyPDC
irNmMApwazPKG1l+wfe1K9bgdiosP9Y4OBwWoDP+ZzAvqRMIrwXnY3LzGXdn
CgAtNFUMFvBLde/nm6kZ/0kHSTSOBfNnzoOLsNKMWnaUHR0enRiL5hP7ibjy
84vW0pOBuY30Dkl+3e8zNIw+wcxmcrN/1tPFlgl5Uh8+M2Q5ZUB0f6N7KPM0
I+MyOrl78mLxvjjpfzudothpHA7MPMgd0Ylb3r7KXbFm6DwqkxmXGP3bDJjg
gRJkmH2eRa6BX31g9ZAFW/n8+wGRiTRhhwORsH/fcTgxagpaxBD4X4y69o/H
JbDmQXw/ZCf6thfmNvF3XmKW5qybHiDoO7cTrYRh7dqIKvG+ltSjMWQvbJ0h
kNiTSOvs2J51YC5RaUzAtVfm4H4XaH5c2vtE5vMUSg1E2MDAUpwgtGPUl3Na
n0V4IMIuIG20D/OpsxPW/fqFtHkJyDLmHQQ7jxEBd8HNyeJL6zqiDrAJNpC2
J/9GvfaD2XeGFYbJ+1DxusBpl2LcdA8FvfGhz8hh6OJXa7Yy1Y9f4MBBvOmO
ylM8QXwC/ZX8lJ5Xk8xMS+DssmsExZvDFA2RNmDewmKjB56WlxCtTPJG4SQb
A7jvwpEm6IysMWe+YJZP7Bb3XuqVL7G/AvJbvLbMt8ujP4ZSqS2jL1mQiSqM
irlhgxZAPJMgvVGFV2XNCAApQ8/2EAudQXU8mRLK+WziyGtoCZOVvb6bS+aF
4fb1Xfx0uac2+HZs7PVaOHVnmmbLSKp8YxYsKwxrtUAYaUfjyoHZLvllLmIT
u9CPjRFc52n3u4P5kjcK3oND7opMFpZEUUU6zErG4hjtS1FuuQKdJynAV4v1
K+oJ94GC4H0EmGNRrYH3m4SlscuqNC/C4LLcbV7lNAuOVBnK43btMjoDXyPU
bai4GhczX1ByiCiL4cjMBknpwdz0rscOmTT0MNRSy+AbssuNPVungWTHMw8k
iPAIcdIFzwe41QwpEq6kgY0qHJW2oNMvcUiNFZ+Xt/f4WzzKYghDvUZ2dffX
pnFu1A9sBrraIrcZHW0icXoB9hEwGf/C4uYovF9EdmY5u3V9JhzGS4TxYSz+
zgKbXf1y+yFsNYa+zOjmqLpRxAR9sqWBNpfmAIq0PN1Vl4OhJ2OGCYUHf3ps
kDvr830V7d4W0JOUDrAgqo/oQWHJNblGpeXBAVU0PxYzeot7NEVs/ps6UWYD
ouUUOAkGoWcI1PVUneo0eei9GYPMTUrtMpARF525QDyVBOQJDAZm0xTw/v0g
73OHcngM2VHdHyOhZSnW+IixBk0c32fMvL8a0FgFeu2mMMXx2/lBWkhNxLeq
mT5lo9Z1fzr5Fbm/T6fjNnVJFa1trf9qO+j+XR/BnYxjfLeC8KABRRwOIcYV
QNV6w+nIE3mRz3eMr2lxEyVLrLmFkgnP4RR+cbymy8om9bVuG18MpN6Q9X+V
WOocTmuwFLAtTqktK0gYyu4D+w5XtIMlvriwHVrOHuhFYs3EcQ7IJwg8K5is
g3QEyIM4waMaIZ0B94xXcugk64z+1SqtHLEUXvJaNwhmu9GPSwYZ9awa6COy
l8BxIKNgQe8wmZnwZblqyOgUAYvpIVpy6UVU/V8q/REs+7edJWZK4Lpo04ua
exY2ujln0wVqT3SBP7SfwWHekuoOOopp09+PQIc/IYoFrgKZiZAjmvmmC0/k
2TGLeAQTbH+KN31ihthyh26BN60k7PTkCJzlkWp8WGqOQnyumtVk3ZS8S0iW
5jDwDQQHPzDFWd4ZP2IBaYS4WhI+Ma/dnih6MdVkrDwV+q9WJBR64JzvC+E8
f9p+qUAExZ4oH4LyKO9p9l7F6+2jhwPP3xLQg3qy3f7fU56qBBlmaiy3cxHR
quAJ+NLtpGc0jxIcPd3rO67TI1mIVr0K9MQM35oEB4E5pqJnzXl5iYAjbqjI
vwJTeI+j5YBw3qWNWPzp6IciehuMANI4CIJdN7vKyTsN7MnSFDoHdKj6AIAX
KP1NqE009+kPVgDuc+D/V3tPYpMOM7QQgDPVX5eZsr04y5QhKe4jX+W0dh+b
ew6VKba9lcTU2hbKwLoVomC70s2VwCmUi7dG6rQdVvhVqyVDT+2Yb5lPaKU2
FJW5uWYQgtS01VtQSX/Bbr/Xi6rGojroQcSoqv2OS7lpUzldK37li0vLjmdw
t6ojNK8zbLODHNXjXqsqYjzi14LLiIeO4js+DVvVe7J4nmDxO+tgSvmmksE9
BbY1bSbDzmDSdjGdPU7ROOVbWNioY1/W6vWLSU1jwqbZrAsLyyahOHMWuCAy
TRk57C1WcukY5n83zUeaq69BA/cWeyNDgwdaLdYL6PY7obkLURzlKUuS8XOs
KZIHMWAdo2+rVuNFgyFI7wIC+7Ky/E+8+emkFq2jdo9sA0XA1ykNo36IuDp2
0tk5uZLcp8GgMq6h9wZr5b6t7S64pvx8jZyZzT6Q7Ko8PNQOlpQuU0f/WJEG
Usgetva3KxqzHFjueRqfQHNBKk39nvvKZoSQteZZUq2YLolXFr5cBPntvRNQ
akkp/OMcdUj/qL8sQ4vveqZBkjVwMbWJbW7rUvNsowz5OBs+SAyvqWI/obXw
RFdjAbYoIRDy4gbrEiuDGqqbEWzdahy5KxtkLrmlkglqfv8dmg/hveT5QPTM
DeqgdqOi71OJf4gpxArq9n7pmpMFEjzhOBRK4X3zRa15/Nx16xlrPyl8OGoT
UrcenNH2k2w+3w0z1xX1fWHs3FaYcoYfLKBM7T82/2P0K7PL16jmM3e7WH/9
P5IXKBzEyjxnkfFsrBrudTANOH81RuCGqPJ4249Wx/redlmYan8pMmIlyA5o
XrPRSvyCLzcLx6OG3QAQEgKuFghLgGD01gY4Y8HaD7hsvw1IPeG7B42zg3il
NFjKFaKi7PUQNyAZtcOo+LiHnCh5jZRj7hYf3HqFyRy0/fFWoMeVid00VTN2
4w/N2XlJWcl6+cY/ujbcJUaSCPbUG0pXEB4yWxskeJO8JQZ4pnUOkVsRoc7B
bizA0TZAHibMrVtX1L5jUklS/1sihiZjTKbtLrkcsyv+2+JjGkubeoqVT1BT
tr0r9p7FyERTFEW21+2S9DwutC4ZChjsKYls9U4V8m0RnnOjegX6RTMDBTq/
yznegwskFm2oCPOp1sxaLkvpAaXf65mCsfbnfdfHqPfHLJaEeCbF9CHbrwJb
+m3KPXwmEgldlwhWCTGrdCXZEQOgXV24RPrbY9wvHfKdn/B3tOjyQN1nBsys
8Fpvn+6kPxUWB8WrfWx2O4dG/usD80aR9uJ6NC97AGjapjactdggCKbyBjI8
n/LA+YFuRptBtS4pBmiX+D9DFzff6V6L9GjHBg5+PU03YJTIlBfZZZeJNdVE
Fgz+fL8ctMol5bGV+kuDNfUsxiCoUekdVqOHhf6T/zG5A4kQfLbshujQyqvD
sR3cXm7Mpuc0mz/OIgRdaimvYXP9bHW+RGw0i86GR9fK4+wmbVUFvm+f7dpM
zs9vZZOLvoCAh0AbF0G9RMlQ9NsYrFFAVjWsXzo63fFmGstxd8MDrDkdFhvY
p1TNHrDkTDTZseRzIt6Ox1GWTrb+u2Mnp/0D1dW2XYo91sRbtcqn6lwR0idw
shx+u0OpsELdwwS4fepk4VrI9Vp3QHOg58+z7VKvPJDfo0MSPRVk5zCdSqJf
z9NOy73+WFxMN82rNOjeWNzH1sYcjJ5goxpm7KSy6NzcTeDDl5py02pIvIfN
Flvhq6Svc7NJ+zqniILzlbvtVGGj6kgJSSNG8+bOQOQ2J6ICk/rLDRl4Hggz
FvTB5vuEHDSru+cNACoTlYAm+uI5Tysm3MX+o5Wz1ez5CwyP28tPTL6ulHjd
y5cjsqSAihJa5/fTAJkDaNRgKAPbPNBSXnv637/fSBDBpbpcVn3+k9xkcn6o
nGENGBiEoHl9DOB3iQTRFmoYf5RqSKYuSgtxyAmsii0ZdxC/NBuK3FSlthXR
98Z6KqUF9hRZjUE4aM8Dwh1hQVa1GJMryMiOP7xSPkulFfebOOcE32Y0gk5E
9OooKfsatSQipK90BHCWg2vi2GRyGttG3hUiLWblR8LDVNmOfZyRIzlubH/k
QwQsgy0ZVjjd1zHE9UlaqvryzYQOqFc7q7alivsTujDp0K9pJPFwWtkj0Pnd
gHOjeMgq6Wxs59odaVWZnybTXQR5oXeniqEgMNTDzyTcoGiCgE88lkWQRN6p
7SeMA3JejVAL7+cV2knaNLobaeNSaxoXpXYE+KrK1VE3KG/GHJhd6Wsgoe8d
XWtY0TVXjOCA4PF+4OKKk+R8vxNTvHNhsrc0DODfiyNNnYqU6SK/P39JmhTu
PsVr6eflbbLGiMjxJrj0G6q+U71OnkNJDyMeazPRHkNXhMpMfs1v8l3LHuSW
lmhnhd/1NjTwsCqWzwnUstoEyCmfTFrGuocH4VO3ua1h/yimAtHWe0DNAiJZ
G5+W6YE12InBVY/Rxj1Yjf/gKAmlcz4bF9gGfjMxrFeFhGnPMCchbn1a0/0f
eFlpzMnozUFbdT9ACGK3vKVpksPkx4gIW1OQpQ1M+sGmJLjNQkNwzedlkFj3
1YniO0UeB+2RT51qDOrx7RhhZluFwuY888d5pLu/pp/IfaTcMtORL9kX2/uv
da1U47Jjlxyxsx5Aep8RfxCNI+ZF+s+hJPqdb1ha9aCC8ihDzn8IHGrzKNQh
PRjjui27sk/gz6M9KS6M1cSq//458nqR0ZpnkHQ/mC/7i8U7maU5yWxlyPLZ
Q7SLK3QBearJ9v67t1mFG8OWeHsOigMgTvqYvf9wMXzHu120AbG5IKbqMXJL
YKVteljIi6ZaEi6b4vAzlRbk4rWu/+HByBdJ2A6RMuK1WEgBasD7SJUVRwvp
w+fORGDsPhCbe46jxEfTEDL0LA6zMTbFuqz6ltEvgMxVsUsPH/B/mESczkA8
5JyCjFrP3VTrB1aqPT9cZhw9ONwkVs8U1DON7f+wXjtP7891Ee4r0KSJir3a
vER7kTa255Utqu5jxLhEyscawWmcKPr7Oqkpj9WbDYKfSHIhFZl4uTtPyrRd
Ye3BzD0gzVvUj3cx1Dq8f4NfHq3Q5GbWvxgkFuSiUvlGTu699kDzGSdHECsJ
cMUwKpGq2POu4zASR9H+OML2GZXqXtuKTOTPBgPWmi8ZnmdDXrZHLff6vQ6A
7Yg0zntEI25hkQMHR0CvkGpmU8umbZs2pVzzBLEyGpyFWLYxx2fNQu9Gw6P+
Uhwli/CQclxBaAJPoLzhjmBc92EKoI9+3YFTQoUBwI2LUSYjTNznZr0XZ7Mz
n2xXz0WM7l8XmSSHSLHUHqnlYC6K17Vus1ptA/YCZJiJD0WMXGwpDsvMCJqX
WLaFyRZXpd2UZAaqFB+uRApY0fvr1WgUzCg5fR0IFLgFwL0mWbxJ2h83D/Et
0oQEMQZsf3XZG1M9FfYpMFPERBL2F0NRpgoe/vM4y6FhDQf/eCnorBlNlu37
WGf4WTqK+mgyagTs9mksxt0IerdK1Q4Pv4DFwtIG+Qg34SJLfDReQfVQPIF5
9Hjn5q4xzX01iFqPBDMwBa0BqTnuJHXO8HCe+eJXC0hhK8HYcjK8cyc9vlMa
vZqE8UcKa1mCc7ZySPT1WWiRKageSU8Jq1YfOSbSlGWvtz9Iw8qwWX8iRjCd
1UkgRsvTutQP16bJ2ANXQi9plcIUZg8lfNqXXP1Bk/7dbcMmdwQgfezUx8mo
DKHNJaO5rcLVBi+AXFo1UHupaxjP3c9rl1kxDlEJAg53Nbk8grphZtxWoxK/
Se2rso7fqVZEcU+gg32s/MgqJ7dmgnaqOs89huYJfmPwYxUSw7nlPnCqdh13
I9YPK774f0E0tRQ8a+/QZGQYQwQUzmSiCcuv2ARKXIJFdlajcIxZk3v97nij
cPIosyVvCX2rKa4vJI1eoLs56dEWf8iHWdT2GWSponZERIzFbsPqw2tnlPoI
xFd7yOw2K4PiAHH16kuRC8uI9Q1Xh0tmSSouJcSDcH4oc7O/diAWNg1rBTi3
TcmaUlUdQkwgu4QB429YLbk47jxG2UonlhaPYc4sdLfJ7tj+dbIGY1dd4nUg
zqBa/x+09D1oRW36IIKuKLuhldrwU5Lq77SDOvtGi/BSOXNtl3PoswYRES8k
NfbZrgpsz12FGZplKqIy2Y9iRjB7TW4V/iewBRqWdqVFmZRrbkh5npf114o5
I69eAqNIVjmakfQ/10WjXYdx2DSagiayFpCukP3WXBeKd4NYxwnbz3Tr7vuU
fy0R7fUOYFgvrmpMOr5PNcTgvk3OMFiz0+rfKkfVduhYoyjzFNHVIsdvuu8T
9O3tkc4rhvkSLsFYTpemcijSO4ZjduuNl5lbU9YQ4E8zY/5+vd9HM/y41Qj9
IQOWzCQ1FeOsV2mfRf/+FuXdQbeBaOeTot4pckz5RlVA3yul2w7/2ZjxE+Mt
2u1YRvUaj2Y5RuxfGmTEfEU4tVLoTgPvbNH0+M3wonFnOuSNCM0TlnbxA1yE
72wiQFHXc6ePGQhPQ2gZVwwwzeIfmmJChmSx6P3folkB02UNjWnXMlEn2vWi
BnwcRkKXc1G5fB/xyoiuT9F5kyypkykcp8buxtTggjer18MxRXq5rgzxwjaL
BYUdWwmjLiJxQilxeQ2p2JJlJbU9OuqKdMwj7LcuQtjeWSG5a9rOQnTQ/ZwR
USvoh0+6XTrdGdWv307isGzMXuuvAirrJD7nByW/Z7b7pbeXi2otqPNcsn1W
ACx7Qh//HHBs5pqGutyRDEAf1LcJ/xfblVW6aGr8JHMg5KuXpTRdzaOTA5q9
eme1rHax7v9s/PMOJtV5k2gWe6JY26J5WgC2b1NMQ+EKi62W4h0tysOIOiRo
MlpLaVx+KLSxSDQKmbl6zimZh/RaVps6r6ZOGdvZXv5hm32+dcP9GsZ/d5cz
Fj5nKveaH+aR4JyBzjp8szEOW4JANPLRXLyEI0IolMa8b1X5t24eD8qvsMtc
athUaHQlaYZf901RRKqAuL3PawtOd3LuKFECwY8FKb48MUYKoVr5keJOo8Ye
DHMBNk61kZdhGB+/c3lsh+ENRk4+YFCIeTUSJ2t16ec5ud2E2LarS4lnDBMy
SpXaivJ95O2IriH4BYfPEB6yqcCTrDuX4tS6iXoDEKIdamW31fUeFruQRcTo
Bl55q+RAuwDggqlqPdMbBQT0WeX8i/PMu0AQkyxa9VH8M5FARsk2nzc8CGfb
3KEat5wzm1lbGhRqJAUlmZEUqkgBnzsz8s93f1QyDDmeiNM92WvyPPA6qX+a
+Mv4hIBwOD8zPbZhviwKcBRVfJnkXmNyeLqVAMqbN3rHwEhEpa6P9Zy3Ssag
7Rne1f+Yy16bJLI00E3tjYdYkBjMlEV4NaXNJ/pZFh4cQ09wWX7pzDGthnXK
z+W+n9T+89bFftNoeozYHgjA0WwxSgzfXEtTZ9DB5ASw/Kwdrh9Psp7SrLk1
KgJrrwculMK4YCfZyrtDOwVxxXMYl/s8LMHcEaKVvX+JccIMWFuA9Ga8crgC
Sd5lh2PbWY1XGaStxxeWxN5ZcHcDGlIV/rQR0M7p1oCtdtqP199zQwVzDxNm
DQk/SPoDvc/eYzG/y9QVnl6IxR9gGWp27WzFJn7zZGxSUrpwUsXiG9VCZOTj
a1L+SBk5UgpvRkEQ2my8Hbmb93eRaIqCS3RyR6u1tshI8qmXRTE2i4oJbAvu
eQXh5HLZmitAY6cqspYdvb1Bah/ZuW5iPZHel6g7dqkSgdReTWXi7kVnU1oO
Mgr/7WMEE+qqWHKFZ3yrf8P6x6hynjFf3cfpnFBwxJJqzC4gg7L+EZKjQhMt
svDAixNK79EfpW+6I0bpRGxzOCTGuUwHaqxyUbCc18vkI5OCNSbM1B399mcg
QPJdtdXkVFCeTwaV4QdrHHuCcnWWHXzVlJEf+itkmYu7a6P9mP+ImWn1BK6h
BexUkN37DrHn54gYVy1R45ESLAsHuMHOHVozaqkxP7gKgOEsfl4PAUmKaW3w
hwLr9Lxi2fWrZPpmFHhjYcTIBMmtUG15cP437kZZKvWPdt0LKjMSCoKP5SgL
8A26XcJSvWk9oq8g9abLyAW6WBZEkeTws2Ux31Rx4QNrwrs/QcJJ0bXgtRGm
xKlQuSirPakQcnhna2AXkqQYtYX/OALoT42jgh1Vp0J37kByIetKCxMv4nXI
7Kh8T0a5unh/d7sABuuTxvG5uiTXmATOGn7CdtCydz3DXNu/d1yR4oHlMb+d
xbVSmqaXhnQ2RpxiAT5NLRTM/LPDjuMJL9Bd6y7sU5YxA/2fIVjtFbKdQVQv
rLBTl7VzzKQP1lMCCh3WJZBAzWMsyh4p+K3x3QJkuJqbe994ZzRsEsigx06T
Zr2IEhjL1uCmPXe2TCWtHKAKdzhu8BoSuHe5inJ4UEBXOFg+tWR5kdCj2WWm
OJUQB14Kw7sd4/ASz2VH7OZHI6mUnL6L07bFooKkrJqNdPNCic0vYLP2Hjmd
tfvORQAhoIwLzVPH/IBSdDCzdz7NtAoJjCIOOvF541L2DRVj3XLfjyfXiix3
IuMfrtj8TNPweinX9yMuXjH1jA+viEY2CZHja71bzpYfiPDEWA/WKskvqQr0
CQAmRjmQP5HP3/0SoFtMpGlMMGEIdmodS7f42bCsvcxRuX9U9Wl4phBxAQAs
jnYUlJz37rGlu6RUYDGXSI5vQIJaJNh3B1A0Zt4UT1CA7qlzvs36RAtk8vBy
5DF4JjaCI8xva8uWe/maFiaZleVcPgyoyHmvNe1ZFQaHmUkKWV7xgNxb2yfo
YAwRItlKDzN96OKv2eoBct4wjGDWEn1KYqwyBMZfOZ82AmD7YgYv0ndKfTg7
FOwlhq3aVMaKfMscE+c7LBmbreaTvPnV/JDb4gK0x9tv3QHKpByeXLisgRXa
+QFl2mbTsCSzUYyWnKBBQydN2PHnHMPzhCTJERXs0ksCfzSJIAFAhYZfzpu8
3u9ch4xySSy02h4CbYVNbh7pX599ZqGCvvpEfxwuzTLLLRqi40Mx66fOa3kB
fnu9lZ9+XzsOxzYovRb3H8VnIhkg8WqnGth3VbGlIp/qL7RZmFfkoy09wUbs
opZMgshfEBRKRMyy1o+jKPqS52I2kzCVyhf/61EIwELpdZic3IyAXJvgFR0D
cjrKYNSu//K08CyQSuiCIyPkrnIgdL/ZybuPSzxWCuV2Z/dkm7CkS6lgobL7
MCi+aKowCI09c29tocqRjmcNXH3Gj0hWbE94Gi94/7YMfjBwltIz7Tu3VPPy
JNgIV+QYSbRM5q+aPZjbbrpkeRzOgjiozzNLZixDwLN2VVofBQf/s10Qf61E
lE8yW72YPL/zuElb6C8vMUB/J97ez7dweKN88hSFbqW5g2Wuf2ydqtziD1aY
/SwPz6yH6nCd1zNlbpDWM9RyAOuUg+mtDuEfEfN8Z3e6VKeK7q/7j7PGiaqD
d4dnWOo0jH43CZDv/cOh7SJHdLaezSolGhC5nk4VwCUxjin135y2nFBJeDf2
wYcYgvyFpwKufx+4j8inBceILIPRWqsm7O0FoNc3KbtIgWyHBI5kC6S9K4TX
rKL+z3AJrQSeAjMKhc+RczZs+53yp8nhYJv6nSNiltqU/DZP81On4ax6iukm
2lOSrQxzslJz5vwgLNMsq2VS2ZDrgx3t00kQK5wAZ1ud58Yn8qb8AEXffuwd
FZaAXXo0qZbZONkFqy3666Rqqrpxxj5DYMMn4bM9k45LOfZrenlG66BmoWag
hvEiV9+HzD3xqUL3FIGvcot2tQxYRllQbp/B7JCnEBK8IGyF/qKEka4X9Xww
MHDVFqnuPyU1w70MKD6Wu+eDmSX/O0cLSiR3nnY/tgChZKup7gVLZqdaNSJc
vMz7RTEnLMURqtuSxo4nF3Bbw/uKzyblivmfZIFqFTj1/yyjqD+InOkRMk+5
fPupnE/qArXEhSN/yZAVSU4mv9Q+pTkbkRETDXr49upclNQOArVexPt+azbM
6iWl7zSn4x/Up1JLc8TlSJwRhRyG8Tk4wcHuZBKVXqegI8J1cV+HzKi+40MC
jIG53WEAzKDgfs0eOJkCn02k7Wmuaz2xr+5unixjoO2mGNEPoomTMCJ5+Bd+
N8UiBNw4QyMRElTnzUkk4SO2NYMeFXkMG9WtrJJ2+q+BkWfTsI8H4H3b1W7o
Frn4OLbSXhUmZz+thGVXTPawUNjS+G7MoYmE6Q1BdmdxObAGpXM1OujMjcB0
tbZHVGpeTAfP1WKgfByqPXQNiDweAWYuUtZ6yZpYJGraojFjbJhiBqTtTh7l
Dqx6La6f96H60w0Ah6zTYJrpXRxW6TscNbtiH3hq6y7x3ecUntBB5GbiL97j
w/B35wMWox5Cee3b/RytOAFo1JZm5W8DwHz7Laox3EIYvGK6BKXcmej6euWY
PqCcyzS58O5JHbyC2U14B7Xu5Px1jpaE6UsPp0lt15zV8QYuD7qQEMBq654L
kd/EkLHy0Wez0sDgbDrq7z9jrfz/Tl8didwdZy6bGGf3t55JMJDMQSxCWZQk
Cu8OP4TuN5t9w7Bapac41G0NUknKq/zONNF+B3skSe/mDIi+BHM0nNKdxQbu
wT5xWe2DMEwFMvweIYSdA9Y3ZXPZnrayQIngRmM/IIuyPAILhjEV8nUriRiF
E9qBKbiyZX5JSzopvhGt+WpqS0RRN1benlE6NHON43XQ+A9iGBWK5ov3fZf+
OrTOZXLSSUfgnlrU/14ML1GO3bwuhi/04f9ZQvgsvxn0XixqrgkwcgDP3H+D
8oE1/7xg6EfuvoxHN4lJaUbThJh2vx50A4FHBTu4sRSDt6d/0IAsaU6sYKku
LfbpmUPsCMRq2ovxmh4iJH3trz0BYtaG+4U1jIv3HW+Ea0+M+sRoo6Vno9Pe
ZYuBoUp/7/Kg70VLEMVlk8u56vPskoUVHzg6vIhm1be9a7wIlAfb93s+C3QW
W4tlj+YnvysqxbhRIVrxUSTlOJha5JZ2D5I/PKqVeHsYrhQNcDzgvs3ooiwA
+2xukGIVnGVDmHKQyu2D3GqETqD455XnrB6pYOUk4HHtphKYYx8UdhzmNo2M
USrYXH4v0nCRCi70XEtr11eRORNRC2AxZtgfGEFQVEExxLVHWnBfWtcO8iKO
8TwfVqT8nmC3k74pGIcYYQYfM+GlcWJD3Bo7FDDZNCBebWwE6Nls+C0mToYL
uGoAWCI73g+BkyoCpFXvx2iS66IcGnws859eq5Pnb9R6kX3uoSJko54NhRo1
W+opGlf9ejH1l6qg1jR/uQVC1KU5uf5I4e+iCJbXC9qdo4awRL5XAPzIabQh
b5ITfsoi4lXJp+4KeuwofNypqzmftVpHLXvEE5qufmvgim65XoTBQz1zBTU3
jkVY48gAucdRymvsLJ0+Jzl2lGwwfkAYN1U/gkguL8EMBQ9zHm/OiulqBAVk
fqRJ8+MqOjWh3rmaE6/2PlgHZWh6kd27k3md23aeJOMV7azLpxtPW/kJYHVF
PSaW291pMAWGB8+xkXW2IkuSo6BaCMKQFKEY4KAx1i8jVT2YqYMmgQjMcvcj
PikskwWkZPN6AfnPONmKv1BACI2gy7FtsnMBE1c8iqE1wplv+TjHCY8uHTsr
P6B/GAVvd1r5lqh+qbWIP/ynuTmwkx1VxnaWHrA/6TKuhje/a3kV3leDDnhp
Mu3z17fR5nWpb/juHKPL3sRbFkKN+pwW7vgjCKYX51DKxjY8a8KkNoYvyIol
ammE7PAsQh6HVoWiRcIsu2YaBfPccKBHswwtX1l/u0TQkiBbJWnIKruBPYj/
CBZjly1wFFkgvYwt/SXDF1JmoBE4yH2/SicnathnH602Il4rA5OyR7VKkFOb
NnBYSnh7gUwARcX+DSDBzyFusnD7rnsscvQBuKfzvAQyYChrSpBoWwrS/4E+
ECasrkS+IIcIfY+/oZTg8hWqxrX4B0Ym6BVinxvtPS3RLDOI2LmnhVKyDN5E
8PM+290Uz16/legyfOpTb5FyZRLhH0bKwewk7GpwzqY79SiFD5xTCuujnUm3
n5O0DXfL3An5ZykWecWRCBm/oE/mHxQAVTYXNem7AtdoiFBr7roV2zDDHPMQ
pMm+LZD1euP0KPKfGkH3VH+i0jOe6LPZJi6Pg/DUENH7Cnz2LHHd9Lmzo/qI
hRq0D+Xhitq7ZmKSIXl60g8EqIWV06xQ0uyH11+pNmDqs7q4lUV7ltKx8ryl
NfouGSIrw/wRCzHmHKyeCteX1wsMj3P2n+ZaWm7ZpU3XOQWesQBRO8diKpLA
hXxWMvLw4hL9FpXtfaTlWrUHXkYpAUO/uU+QN3wA+0eFUf6VK/xpi+d9A0za
sJqhiVi+KIyEL7gWEoisZWfPcOe9kwYJdkL5WI66CR1IuLSHgvWFLcI2EUn1
uj2tx7AulpH5iBQqv17Bnm+qFp1WCnRyFv9xXPu/+Thnivtx6xpVRLC5rJk/
O8b/Z+LE8LY400MbRctl0cCDCQ5WbJn7LRg3IKZtfNiAKPRpzSj5NbUx4VnT
K52rWncOiV0IV+ifLs2+ndferll1WOMVndTd6SnuBduddGTxLXYEKVnD2c1m
DHiH3+70jdoET5Dsw8RLCzK2aNU5HLy6W//XA9tzkRn0dHfZCcPVsrcjUEXY
Jgfiz3f9Vjwcr0di7jq8ean+G1WCImPYwcNC45gudmxhK6OC9Tu673nTyYHK
uTppaT2hYHi2FMgLeETpRlnrtC+flw2TzLw+BP3CDGJ0Rmf4XVZSEXkOc+I/
vCwl8I7u6twWow6/AranIdtDigvg/RfHFwRXQGtHt7eXPhXmOiAerplJQShd
UZ3Uz+o8I07Nx3ZNl3RhAk2sChwmdN12EiHcENsrBRl/w0yHk/SZjTLwhFWi
Vg+2GBSMjNmFzHqwyWYDWjf03S/PE+NE5fJvdEh1s5k+OJHLXRxbcVGNghlY
Wn5TwaNjDCdY0i9muISy5zGM7HARDPSIdeVDlxvTO3+ywmzyBnq3qpWqVFnN
QxX9IDw/n/BIVjle9oLV/d9NH9XTDhRyAEbjsEA2wrBcXjvNTjT1o6YnDYDR
jB4a5Q2dvVztFCKJwg8/FbTfHDw+Mw8mBagiYeAMdJPeKhnVhcE1uinFV8nd
RpkmK1wnKQ+//XonBAZLyZDWDCNGyCOpwcjHXkLYq6Q3u9xJ9BhxtUjGPM/P
VgeoMsJGD5aAPMeIw/NkEBN855MbgoBc/HkUT2M+PjkU+AznFCXtcMzyUROp
yd8jBA3s0NuY92PS8/k5B/NcnGdY75dqlVCZ4/SiIibaYGhakcDHJz7eJDab
tFOfPa1EM5fDtkSCDLB30sbhzZX9GxQrw3YYqrQyG83NuJtdjXnPak7JM13f
3rU0kqdb2gAArthE8xJEN62S9IKDm2E+VE8J39xObwIZoyqRB0qjLynDmVeT
8AYaNtUW0zNFXt5nN2KYDfchEH/0nMFNzXZuTovbdU57NjuP0hVzBD0kOmqH
vHEKeQ6BI705jK5TdfCydpn5csdTvu/Gtpn85VVFcpA6XuM19g0w2i3iqCwB
odnFtDqnf6GsedaYKdv7m9aUftBSfcP9Dv4NK3er76cPx+b1ylMaYft6fO2u
9yyOToq/z8ks1tIhKBstzqspyhu5zLa8kCV+ZPv6Pff8ZVhWh8VGBthYuwsD
AHl6drBv2gtC/AQdtMe1z7QC2H1wIGjwMIKHVWTdsOIldfS8euEDqJBizpsN
vTcDBy+BbD5LgSAyUjEVGXjZ5c2Vjgk43Po4XSPBwFKdFQGyLwFX3KCalF9C
93HzPFJdklF/XSJ5wZv94wOpSVl4l85PaPYm29fupdZdGXzmNzeTlsY+wCWN
U3NrY4pk7+YX/nFyEkwuYqeCntmil6frxgVveUkICoR0gMa+apGeyNucNO/u
8pAlnk0jgz4SE65fCkAjnWmN8y4eNn1KuYFQtNGk7UfP9BXetE3pycDKe8w1
YcVyLeYX8mzwxhmvAIyue2/Q00D+OXNv3XxamydcObIqR2p+7cLTxvHSuRXO
lAG6mTnmAer4YjMnoH/0QZyKA7vYdLCjYk9VYFgnobRd9aiAULNaP0N2vnJl
f4znONuM54GEL/yvYdY84jIe4rc0qdK+Xk83cT4CliskhZh+Z5ixiJiZJkWJ
42Wrr8iWGEAPTuhI0gx7qwVnWRdffBVCErUn6pHePWGRfiIjywd3+xClwF0u
4QV8og8okT5cUtZ2F5EsQYDEH//gCtjU0hcHn/eyKYKop4tFgzR83Or1wrWW
R2Xm40MsMEc11aWFz1lksKngLMoKyrMJlrH/TuuLOIJdG2JWEXXIczqBx1sD
bWtBkKDiX/HgJUovIeAaKJY4oCyhP+huk0mPA3vxuYvS6yigk/LDM3NDK42S
BRgpFmIBbN9V5dDps8j3CKBpUvVBF8qd2goCfE5T/uqfEqby0iL8xuKbE2Yq
1JNsuzxl9btTCTh9W9EeRst1/z7AlVOOB4OE05/r6mpBnlteJs4PHCL6Y8sa
aQMP5czBJNokzU7YHxO10AUYfb62rxEorFQFXRIzSfuauSRn5XrThjPELo/V
7hsayiJJ1PW1hOUuQjmqzd9UC5rI6B0s9LlWwuXXVgoCRUl5eoCgHfGrKNRG
wnqLif/1jYYMKJF8Bfm6MtpYlGNcrdcNhyCL3kT21w9kRmdSrjG5kRHXNXd3
d3gcN/yvPSFPcDgmGbJ0eG4s/+MzBKWuIqAjQzpFNrBNF4af8st0bTw0gFlX
qUy2zlNGz8cce2p7vf2QLP6ODLtQkAKJyhJ7EONrQwPDsudH1S569mMsHTkV
Plz/ozjt3Jn93GTDk9VAjfcwt4vhe5X8JBNT81w/iSHjLlsqfFS6uZmCniM3
LsTix6wnnXG/Gj7EwCEZhj47bLMKpzl2eJlVhktnJWd5zZw82I3Qlac1RwNK
uQsqGQQ7qwmMFhhu9itMM4BzLM0mjKzozxgc6lVr2Qx7Q9F6/7AX8vGrCgDc
1XJLqHLb4bMmc138pxjaeO6A5c5uyMFJfT8EHpePmZLc6LGeSKvgmRe5bezu
STq9paCe603NSBwxCzl1RxWLIxM/fJSnUimxYEnemKtWRcfsZ23sowjz00Qz
HIMfci7BCIzQ9UZ4/8GZy3QLWpl+HeiZDCSiBNNMaV/F1i8YSVIBgO96HV1M
sfAAaiabhHZUCDrR3/oyVxq6r+0k+zX534PWLbPBQuRG6Dlt8YvU4PGbne8W
/uigyiaAA/USmk9hWeM28e1KPf8y1wFZbyPT2idC+pwOjrnvfnmQDZNdLN1W
fTfbhrGIHN7/X69RfQoWIg1/4Xb3BzL8EpCJ/tNI5O6+hQItOK5sNG9haZJM
YeQ08hA9IWxgEIcpXXybtdW/XEa5aPhzLsigBukXMCCAG9kjhWNOnJcqhIny
3ZeLo2MWndxL+J1BywxwHYAGl/vpSmS/arkcJXKKI18wYXYT9/+YDdnBKeZw
Pt4hsaRYfG5awfDliUzuzqEfAw41DEJK3GbrZ5LB9A6wEQ8GTQilXq9oGTY/
5wZhYpsGMoSpExAfekogWc5QNqZHRExEh8OS2NBXeaEuA/tuDcq35frqlw9J
0YHL6Z4FXs9JWUWgkaFTtVDeHqIwfvzBjC3O02y+r6+Kx39k5ukwx9Nm5hc6
FE9aBF3KNUIwt5FrkEVhq5AiXFzopqkz7Y0/WDMOedZ59ekwl4zbHT7JKolo
7QtEaS/LSQrHBLjoKSnIaMoFOwsVQjEV9/m+4Bk6UnOsDRLYx4uY/okti4Rf
aOHx7/bQjO9WGmNGC6qqz5NDb47dK3SSTVesUvbA/222nvad17d7TAZvg+aM
JoF6Q0PqQXPddURsX4VDpyMpTrUf6grwrvf33Z02sFVLlaruKxjHcpKknDIi
jWtStKd7qgpL2T08WxLhgdH6yCpUYYM1gQOpFzp2h1Vf6H2YgIp0aeW3BeLg
Qc1m3iJWjFzWc0qNMLniX+CRScWcQhEc/J2nL1Zwk+yd/nm41MYGa5v1rqjw
bCAgYrZdInY+M/WrHrJk5x0FCxlqL3teoF4un5h6vqOArGKsMjLvwwv1P/oT
L7LOlckNatPIkyDiAyXEt3V+v4MwD4r4qxEYkj4Ef0hB9W0CyiqChlxFjfP9
27zQBWpWTISYXQpsPtlsYuxHI3kfBeQMxfcqPX2HuSrqR0YSGaVnVQnHkklO
mkRIapPvmpqK5H3hikBXD5E3tbjsfKI84ifxENtd3LJS3MTGtbNS4GrDHZSE
UjglFDxa7+wvxV+w6tYFX5/7Xq52khlkG7FoW0eaPIUXtcRb5nFZ0kUXwGJB
n7oGGGCmyM2rhrmk1Ox/5T1es5Nt5gjC77BrF8O6C8hncySQgmDpPO0RnmJT
/09mKYkkUVyRjrEnLCQiDNkXe29JPz6LWnujexuILiykdv4nzD1R7ygO7ghH
R1xzxmYJXn+NXKSKDnthHBnLrtHz+GwWaBwX/ng5RdY9hec4D4s3o9Tm7cfR
4fbhNzJG4Kb1ShC8WhTzRuOAW349isVqFTjRfH1OuTPgWdbpEohrBcK/a6vV
nJDBlBoqvtc0tums7Ac9wCfrv/BtObFqUWwzMZ6N5lleU46cQocMjPitvEPs
IhZR3alDo4fXR2iUlf9xG9yPrPWLwCPX8bJd7cB/KHeaXTBsAH4Q+eFyq0Qr
Mz3L2ebbBAAY+y6ooslTtBT6PR/4ZNCNruwTGrczi2yJfYyWdE9DLTQsGpLl
pN1vXL2OiqryjgleQCbB8AmJ6kugkKR9qFRF1iDNYqImrwRiBUxiGel29wql
czvlvFzcS1aoxe29CKwRJpsp50h4B1fx4otu3ooqzEYA8v3nTd7HNk5r8/2i
iZnBSV3yfXg5rXyCgSI985iw3z4TLQ8jLC0SYoB8IWfL0WD1ZA735KyDSmHx
9uAeGSYkIWML8IaNiSB8gzU1ri65pzuDvnwWmraPhG+00QZEy973kPndR/RL
WiXsV/NyTUVX8aQP0vVaAecPuaWCzXfDT28Nfkpa2oTDwhBcOFk+h3HlgxEf
RW0+EjXwKDx07mhr83yCkN2nphVOmbEKn5sAT44xmGIVLPMGMWKxlfDb7tY3
qHZJPQfjoMyZpR/G0BfQNXKIzxu/FZ1p0s7x0hg9+lltN9toidXaNGhxO7pK
Ua/xLQO98aGISjrbGLtvXKx+wWR5qpl3eSkDKEdhE7niWJpU0tFPRdQFM6CC
NuEa8FxxSSY76zPH6S7SpJPDqTPpFttjsvaaMe1k9JnPLH15mA6tJjQ/6Obv
ehKpiHDRuajaTskHgNEiptbBPdWhICPZWYN6a3QrXaozvYYeIOGZ+r844/bo
vZE+QnCdvatQMGdLANXJgSCArWWIoJ426pADmWwMnSe40HM5wtI3DQds+uBZ
wKvH/Pcf4phxuPq2g42ZQpi8FOE1zNrmvl5wV0xusnlcs37fAkvrTEBaeX91
CnsI2/BkyJltQXV2TdAxx6UZ1cZwRPhlySgO6/CfdCTJ9UnlB5WkqQIn8duX
4uulJtsnN04mqCVhQDOscv0RyfIG8c1ynirLOeWJNaRQ+z1KtWb3OfmU6cbG
dmDViKYLifZauqdbUAP2l6tfZjIL3SJDDBNIG/1Qj9wK/cirNqtEWjE3ZihQ
ptRgj6n3aEUKZUNpoQfo3C19N+2LQy57jAj6PJK9zI+laBgh4vfiUUu84QJU
yC0QFtdMw0+ACY1ptqCQRp8lURd1NeWfVBd0zE4OQDCQu2nBl2TmTJoxQms+
faYzy7hI8/mk6wX1ifKtBbtds811oFPPnvxfOdtlT189GtD9vMLTTy7g1mkz
087wUnYhRdvMRmejCgKcsuOkfY6EqWgspNp7VZ5vGhGLzWC+UjDg83fJri4d
pGooSnG0rU4Ho37HDPl20SwcQs2TkKBsdXORvcaMxJC9GV+H4vlByNJEbOJG
mlR+XwBg+8OveOxFl3TZbHrf61izEau/zu/WigkeqU5f9IG7CnxnSBlwBe6K
0g1iW3WlcmAiXfQCUGw3GWD5eJDg9xl0M0cJClYE9Kh/VUTqqIYSv+341Zwd
SfIiUef4/zgazfbD7nSrJa+JZUOR8dJQJRHoIMbvGJUckkNhUcXwuNTL2dC5
zcOK7Ez1XDkatCDawingUpYMu35FxUYtSD6UMpmTEBFqGIxInCf9yPYVdgQT
JoJ3sz29RNQV/VYNqEg5ov3lNfod9fAu3TtmjWx+crZPnro8xtuwV1Mi/2SL
cMIu/sPM996AaHDIpToluQrFewcfSWEKYjDxxX/CHnLemsTsS855wShd+0Su
8o36q4AEd+x4SLVp+pO/M+p06uZcO/Vw3u9Dvsz0AgeG7LL7AFk+ltsp0tLA
Kzjuj1pNXPyoBcBpKbDb8VK/ljCsdz4pi7b5Nv4ULJWy1/TXGCqO9d2xdlzU
Q9GKY1fNiRtkmf7cv4CxiPgVTkSjFboW+jDeIDrhnj32PM0mPcJyCv5Fnq8X
PG0Rp3jlzEpDLxn6P9kkSKmLi9H5OJ2LDYnBWBm3rDBvvUs8akPWCOzwQn3X
N/IZ8ZwDjHNaUlxrDJgexE7BDZ8RMh5CnRSzL1oPHHdm4jIuZON4ecj1bn88
4EiCRbzUenG78tVsnLNK0yxUcO4cM2iqfVS9+cuW/Ul4f5OpERcM/XVu6DeR
opyKlHgOdAmCCemCrqLEGldPP+EAUyI95bkjquzwBEp25EBj40ZUWq0GVDKv
TRjjM0hwElCFm+GdkPgG6J5wwFAs3F2bPFbNqlliEOxmsfyEGMjAEX72YW5w
aQYN6R2FIC5ixI9dfCOdxqFe8aSDAjYFeKrVu1k14YMaMiy2ARBVJzataR1H
0MD+tpgs5cO6W5wlvYa7C/FB2dPyx6RhhQCF/FnaH3WKYj2/L0tKAmnbSGxo
9PmHRw7Er/WmXIKlIPhPPAQFGgk3MvkZVYlhKzfbrttkpx/N5Iszan2qJ/GV
pALSxmhtG46Ieo/uBFQi2opy4EZ7VIYWxKXClNQu6g/b7mMDxPtYRyxI6H4X
ceRifpt8rcM1wLGAltAEefTxvZVHZ8TLUJBtfJS0K2IpL2CX9JT3KWW0OPcL
mxx7zzgXtBrFm915AfZVsWdtVqXPqTJrjvh8UzC2DRXJYBTDhMZH7kOcQzYE
XhXLgYodElGnu6uHFzR1Fz8R3hW9NHESS90qhrBjCAzlSyimDmOGFsAzPvp7
3VAhz7Z0oED9gJReHFFeujkQDGoVVaNLfTvlojJSZSSLn6NM+qEM4Vl73mb5
7Njnk5DtWnxF1BiNE4TTRBI7nthzFkTMUv2VqbyHEs3DpIwqVYdzIeZcwR1F
j/79MSwoq4T67vW0JIradz29C6jseAqdQMO0tP8asWlbGGLTzc6V8RAknsZe
65khIn5Fd6MenIJ0GK8k4PBp50mBBrfRStl+/cjbqLe1tua9r1zxpMarv8AM
5sAtYpCVnpatnZvWggNqlC2MfcoFB8nAwOS31uqhn91CNyAOxBysVcGXPdsr
V3R478Gnk5nV0RMRY1j8D2lW4OzwBOBEF8f3D/sVigwx2uizFiJPJZKApJZh
6PaSs/5Qma/Q9faULWn5c66cA9nKQhCmEo5PqbuUI/AYb2va3x+My8KalTOB
Ll9lj6xVFJcsTURS5ipxcg6nLqyGq1KDPb+hbQG/XdCkwE2lORSQumcUYmc8
kSFPherhfrdi72+l60HrJpGmNJc1DBMxZwlmd1uJXiG5iDqkGi0olXG7oChJ
UDAgCur/9JrsWHud9PjN8mNjbd3WELSqv5ivRGjHOzf0nXtCqv+hVSCmY3DL
f3aUDCRqA3+EjB3GPBy597HfRLR/wW6yh8aMynmiz6MZa9Ei0aKtn88moLWr
FnvwygqdOKWlABz95xqg0dVPOpUqIP4qEmCpoTRbyHdsmZmK8yTU6D6XY5CV
lhjlJsKkBkLZ9ypbchteSFvDSt5BMOv/k+OwyrIBWz4h/CHSv+vPx/YSIZHD
X3hke0HOTeWNk8CCQO5fhfTdpI5puWCDLBj5t3PhR82JCFiuJQiD6NN2VzrH
WX/KD3oykbhYax6eDHbEgTwoYoOUVRLVhk8T+a5K3abK5WSlLkAZ5WkVJdjj
874UhcbFBsalQr+DloyLebp1Bmu3iyB4DePKyyssHU65CUSbREz16wz9LqcT
Z8SxUXn0Q2vYGyRhikO/d52oR754gJ+oJnE3cqSyiNP4V4Ph/gbTVE1y6MAt
BhMRb7KbeWivpbz3qtHwiJiila2d7FvuHXLCkRCT74hwgUApjbYlG8F++YBN
Z0lyGS9CPZxFwa66OfPzVQWUa8nKQsWeVn7AnUlEIEHfsCOmvK6yP3RL84F9
X109JFVNzMSgn+pTabKNid6GwQ9mx7vycN6Sc5uF+Acux1cTRC/ooQyRNa35
SWgbX1cx+lFb1fWw9yxGTUwe1M5cI+ni1uLPik+oUennAxSRFuZThu3XPH76
yYNxGk8qr+cCl+Os55wgXCCxFFkFTyLQSbYm3/WNlBG06+FL88ojzXYRI/gd
42ox/jDTvVQXQmJzhMvyYBlUe6AGEai6984vGFPs7KztQI4VF3ch7GsfyN9A
TBojkQpS0JrxSdGNR4Z/eylQtLJE00qa9AUjxVCO+ilKZ4l03nDn1KjCGGHT
gcMPOCpsnBCB2NDTY+SXoTJ4ZC3PFKGYS8YpWshLsZX835iwcktJCoRxmSLP
d74u4cFB+NJ5e/cazP1sCqgTtpHjmV8hGfvLs5HdERh/P0G1KKeRfGgEmVt3
/iG21GL/GlBb7g01NPrWPaaJGbwyuDP+fSO7qrjOoAdicbk7Ug8XsaNp7vxw
tTsuvdFsVbH/mWD2kiYbXBLCmL6y4hj8CE4ML0J6i5bK+0FX1/k7YRvNW8KX
WDxMhRaqdawNe2QQGvzOJKfaY4OkC6VBJqNRw0ex0Op6oFfDUJMtBuSpO1Jq
hssylYMdnS9t7f98rkcF/ocQVI8fozzJHYEFzUKGtdb3tY46Ip5+O8UiH4qI
3kNXH/8Zo1DpbvZVIM+gnhyen11XkugIUi2KtbEHp/omsT3h9rHzsy0JKak1
fnTcbzvxfqQ8JKITnDXMUM3pvXy3sX/Pra3Dlg/m9XH0NBLyKaqV6zx5xPmx
Hwe99Ms2JoHomdn6RgsVHVJ3D2OgGaH8PWiy7dV2Tfb4ODUJkgcOiZB0s/ZM
jW0CpLi84AMEqr05Ld1U3GNVSfAxhZqnaYCCbQPnFKsz3g8g+JmjX3mxYQ41
c4cFRiZesWFCHBMznf9BhWIykqCO+IlRxhr84b4o/6hX76aI8MbruT2xsCJc
D1peGKN9gPzK4ZLMWyLxIO1k6LllQX1iqBxo2PyHOM2rnBpp6PD+SkmOqliL
e0ya4+2PaYsoj6+MLgPeJOvTeWnkHSKzSEX/Oa28gZ2KA5RhrJ1FUt7tVObx
54+2PSTPfw3t73Y1K6470WqPQoqCp18l9Cv+yQ/5HSY5GGrUWNe/haaEKunv
6su5YLGXJcT/R8ZSczHSTpDU1a1hHfnUdijx9gAk6CINAl7e+5x6UTXPJgF9
boQpAOePqbhkojNipLQT4fgme/ZI00bJBOEYV1lOToLgd0GO71hhRhKfkZ7g
ZAp3OiMYF5m9YSNgTy9TBr0Oz8gWSl3c5Y0zH8udPyiCBP0Z/2CG6xAUvhFk
mwJMmO/crxZyn4qC4qu6vArh0Tk3a8gU+tqvhAlH+8jBzzM16QYdFDRsYvZe
qjscNoOoD9CobN8xhfb7r+EZRbgfPhvX2Jhq5U2xzl9drPcjXP8HH16ZtjUq
/carErElt9ia0J0bV6RdwIt54adm2DqcWvRpEh9diCW3yFdhnuUniujZapyw
FKan24mPoslN2IaYnnnYFg0t6I0gsPtcaxjIL5DuihVjRd1wguiOvuoTfavQ
bs91bUFJqY/5ZTAeo7PZqlE9fbqkk81SaN1zmLV+MofdG9li07bb++xJI59C
yAle725+mh3RhMiL0KI0ttBBR7wrrrmWDsHpPkyCb4xATmpVNsZ3v9dKJp65
/QLp3rMSATNrTcQLvcLw1JU+4bWd5zmNq/f2YvnAlqnljem20fUiAnAfLDQT
ctnKoZhYGavBnDO8s5mdD9jsdc+/QzKDbRRfHi1g9KZwKUKjIo8QcrS1mZn2
aRuwsIQ0wyKGj0efRDovqgJgGASBuvvzxrSs/IpalLKnnAaveedbax01TtoJ
K5gT3FxVaqeXdI/G+J19nIXfChDR35MeXUf2342X7ITgX/tryvpomuzhzH8w
c+P8BnQBPm7hNZByR3SBZrSAq1syyiEDMZqB9KgHkDxx7EBJv/Q9Bxu55tR+
rLPAAIHYqgcslh7HEAIncF0oQR63Xg1hxDZjYQWYwJg9+KcrLWXkn5VilfW2
+NKDU0Z0yEJxZ7FPjHUfXlL1LvIyFaFjyV6scJz/qXtzTaDlMXfWGfTaPjqL
RW8SPE9i6HsE7z1prcaIQFE7eTin+UZ1zXigF3t2W6ZfrAJt2p8gVNojLhv6
cxKSGlmMnpEZAdp8w/QJ9dZiZBG2Bfue15v2mGk+td7U4J7RRsn2jueN6vJW
wBAf8F0yKyTOmoZZGb/IQweNqal/Cj1TWS/bROFzQIK57hdqabx57z4UEyPt
QJv2Ammqryg5sg0Smk7jxmLVHIA0cDjrHT2BATsXRZe41jIAxZ+4f7nWGPHu
SM1suggB8VsNTbHEH7USpi0QhlaXrDxSAJb1jVeaNi/mflGC7mdNLR9luWYl
4mpEosXiUSUc5Hmv4DeoNt/epu+jJNMQIt7kMu0Ju6/4Pq/J5zav03PVZo/g
LO7JFuLCsNtYiccdIswIwwP26J3ORzG3fd+JMXHQSyAHS/uUo7Pq13osBAR3
hGQaKgh6lMabDiLiicZIAUZuPatPayZE3exyOca3m83haLx58JCCD122wbQW
C122fMGE93IlQP8fhDg+e+kjyUOSjl41bIUrCxOQdNLpGWLUgJEjy9gI4TRx
kkg6UytLnKtYGMCwp36AuPg3NEQQpycJgZVjy3rbn652A+EqYj2Fpu2Nviwb
90DAX8YwRdjnBFDXZUoelDk+oCGBJa6JFJasT8iVVKc31Dd2A4+LaxZuAnw3
bD1ZN0LFgw4iSCeD/cq0XgWI7Okhg6x6Gr9st7m66zBTjrx8toqH4gwkzojB
a9d9FbTjnSy4S1E8E/tK8TRkDDbB7khi9nAofhuPkfE6TxFIiesj3cgDxT2T
LBhE9ndBTrS3OGU65ZVmMJyU+ye865XcFl6JXn/czX0//fL2LcKaRz0FWfnq
xc9CuAtn1Md2ow0c8GlRCnpDMVh9BnZ1WUCGwtr3h62V+rC8MzXTxfDxo/gO
/AaeZFNnYRe17dfI74XQ/PtC1N/pvdeIyoZ8TzpZff0hy2fnabDCVKwE3kTA
xapR70Wo/FbmyYXkODNIGlbDBxMEodmgBLZpS7UJVRpq4FjIPPaIe1Fp/rNE
Ade7niBZWl8JvIsM3rlFTZDhzVuWR2SbbEa1oXPtFNMuPMBrYe4rxING265X
NfbgZ49YFUJBETfL+cq86dF8sxoLq/hnD42TClMII7hpVLdPb9314CrbjxQ7
I691EyLlcNNff7fRIZTalPlxm6U5azV3Yby4pNyHYN2pwFDkUK0q3rg/kb3E
07xgx4UhQRS16x04qHx5gyc/kmDZ3hPQYoIbltKTpWcRXOW9O1kAl9hLKVCv
7G7HOkGD3Yaxg0e5uD5ljf996dDKYsCt96uqsFHPQyGtLZfsBtAbwu4EtKnL
McOOXjpzOIiEjq7DuVd9H/tIeGhFCaZDLvKlj4SKxbi0VRIJDfdfSZgMS9je
DEBGFcvDFS/qV9NdqGl+Rp/6T9o4kYbYSNCjdi+EnlYvRx/U3zGHKoYbwVKV
aBjUdDQP1neczPuHKXM1PSMafBNgzwPdDBOIeeue4anldN2ke2OOGvmyy5/d
kOtzp3AGSCn5oe3aYubwIJxyZZjUe99mAGZo/DImaQp7ewGc+f3F3iIQTncg
iobzn85Wpw+1eumMkceUUBeqrt2bvMpISHGnkH1KrmV8/CMKhtAEerWerjVm
Uq4oo+ucGVb/+zItVfwEbsLyMk9gMz/2IcF3ZZOIarwvK/LN3VI55Y1mK9TY
8kegF2ifzPLUBtaLiv8w0721CmkqJfAGEB5fd3aEzemCjm4ccsK1Zn643NCh
udbtu3i3CYPPmShK4PiBxP2BrImt2eqgXhD5L2BtGibO6c2fR/lMRgI/z7Ng
dh5D4UCFq9uU8R6hhjxQoId6iRMRXc4myDJrqoFosAc03kgOXmYUbhHnikzL
FqTN0ak73PgXjMwxrlUSfIMIclfRODlhMi9UdLbCZo8QnR4GvM8gO21Z5ZQM
k/6jWI3QnPl3SMLeVHBILmi8zsWJsX46nmcSuQHQgEqHr4nNwRuDGUyjzQdA
IN4oQZx5f6IjhjU1+PNXgM+4SaBGJZ0q1yYt7uBlAUu6DhlLdPAxLlRzhfOY
KTqFwq9rIX0PkPt0gFr2Y4C1jrstzY/OC56zEKUoeGim2yAxxFWmI/lQVkoL
gVfhATUKABXAlivvPX7dYsw64o2fqI3v63SziPjNKuhspqaCQ6/QBavPBw29
YrGtsqRecnjiw150glstPU57uNWugi4YA0ZEEygzC04ks5PC+IQs3N0khgNv
GIBxVPd6bJ1VvMxYA0Pe6bmrkJtms5i/7LsKIfPqE2Cgg0lboqfgsLk60BM7
8WeFm7Vvju3R3PCZ50thYlb2UNXXQLWWbCWxPHbWY/FgfQAi4em//pqgd8jv
q9RBvaaWUoQNExqh+trD5zGEe3KcVDt0BHoLxiEPdKIYdJUhRJ9mQpbZlM8K
Teb0BN67KRjIsk4FGCJ8xdPfNzEUWGftq6Edjh+siRaVmhgz7qSuyOD7pU+z
NUnh8bL25MNoP6DKqvMr2YxC+jzHvTfzXxq/GwEjD//EOZETZlM11u71uKYV
jjxPh2JFmRyNCG02TUAMy92bAxiY2dOEXKtNV46t66ZnIVsrQQiKMLVzkP4t
OXKCPQz9myde4NIT7vG47LMMwa6y0xz0WOeiA63aMqmwed3wMstS/Js9GP0K
/lsTINXCSeLhq9zs2+t0DCLpRzdHy+d4W5nPyknSxuR90PntEdbvd+vpU8Yo
jxN9VugKPDzOM85zZ2Gkf0i2Ho1R4xdoA4kK8NSOjCEg4X8eOWc4h9k43d/c
k8ITD2sIabJD99G/N9yvwyw0ckXuts6PWRHr6v6MG9OpQD1Xb240GVCZ9/U9
ukZma4VjP+FPWJi0WqZGZusGlR8mz1LRcButZFSn/24t6ecyDkuf95IUscHL
s7fLDBOVgHaHlXA5yxTde2qmKJG4Bq6P9YJAencmLMgc4V9zNk3IcXRd3tNr
Nd/SsBIovMcMz4OpBcPMa5E+nALQi7+3NieDY/bLcHQ8Erx8dQsnkNetF0pr
q6TCHJ+XnUAvOLlBpZpRJRXbnrxTtoNyt9B4PSSn4eVmsiaziCoKIlSjtW77
UP5wOYWOtfCnn+FsUUUFju31GYitImFaUIL9D7alPYhyFaSEgwERzJzHUEsY
D99bK4xg3wBGYkVqYTlb5Y6bcSPJuGaVSsrYRPja2UnNCzDjuCx0429Z3zhm
/mIYiaZo+VdeyTBJIG3RhVGJQIfiGvMXi/5PnTRVZOISr4b7JirXH6Vaxflz
v7yPHITJ80UVoPA3ma1aZRpnTvml44nJ5vBDe97iS62HdWo9N1m+ubdpwWm5
K566p3sexb9U80jMVZs5LIlYamXQqK+xHrmmkplzYqhkyxmkB6AJrXRVqyJV
+jDYnx67zTWRAA3QNsCFM17G9RIs5yi9ReZJIvxPEAoixGlpvjExu4alh4g9
TA0etUqCcKztMt1TW6cIlwgkfpKHDmmIG1qoUKawk9gMzr3YOCCv+xgP/M+h
stt+tMui33oBeMLOCOCSh84xsE4ziFo2O8Bsh1qsApDdN9Bf4m+f+5I4ZeG1
9Tw96TEQbwgklKuYOta7WCbUXwgmsHJbjn9/qm7bkzwlZ0z3wwG16vxmHMLn
/tm0ks9StdfMsv9OuckIxS9a/ODAJckMLEZEZadYpRSH/mn8128A/QsYT/BA
A5XrOceyl0gpb52osoFnhMBqn6woIXuY4eMHglRcYy/tQBy+zi4YQs6lG/wJ
kp1Cfkuv92hzPBa1AWK3Alk2sSrf3c8g/d0k7S5JMHT1ZMr2bVse3ly0A6/y
DcdTVTKLIBOT8hSnHPgpstldtVAN5cO/vZ70HPXnOJXi6Fh3XYG90xtcNNTS
JY5bFNR/nMUduJfRpHRKGdcqR5M4eHLEJ2aR1shZ7xbEsou+hFrdWXQTx48y
oVw5ase2Oe8XhVfkSx27aM2NipJbrESRH4HUPxscADK7FdUztjvYGJOV/xhZ
JnDOqgAzhtPr/xG23WXvTFcmnP+q6jx3wFzyLWSSuXhQwEwyz0aakGbr1iqH
hEup4Nkumy6gLUDZ37cb5+/WMHgT9Uh+6sBt//vCWnColLsYdLO0VZgvtnBh
P/lcFrJ9sGLOvfFDcar0Wp0vT4bGqCX0sqyJB5S5hz0qcdnYjJq6AwWZQkLc
26ksKk12H94xMzPkuSNvF4vBW2AA57wV0JukQIxkKDgUf8adm1te4brKYZUX
MH5NnMfP6go42w58FkPFRn8GPNiNisWwMMGavANr8fVPvZDBaATDZigmPvcu
WyC7PLB/kR4IYS7K5Obwc4JI+lEildsMFnfZP3ANU36dGBHdqEm3b8X9Wt9+
YNhbVUBgQ2KaRVtUOOEBO9R0N7JH7Nu1gqnUOlPuML10nO4soiqOeSSlQkQp
5ay8b5amoadeNtPrRCG0YbLh2WW2F3FHMzEXjeQQ+kew1Lrl1fMYGfVPkwlW
yRXza5lg6kCg/hc1kfktWp6KhLk2iGPfkr4riRk7Mx+8GCIZq4KgLfEtmSJ/
an86KrcSjXWWMTb6EyKbueqdZz7T4jJZ4DvwBCL2+Zjyfc1cM1ZQSPBYY1ST
PWCTP0El9ZZfG7EG5cA4pvXagMVlB2GGf+rBKhuyP77x2ZACeYMK0R6WAxj3
/z8jT+tiBccpbHBXlCdoOgqq1Gbtm4AX2kBzo1psXx92Cg+pMHCQBV1T0eN7
02VCl29YYMv3eOLtUJSN0JPmlakwN3e1Yu2aYk1W6K0afJ+AR3oZgDvDBT3Q
6SO/Bv6fc9EG3eIXCd80s8sui+fgM4Pw9JMdSaus6NID7Sg7rIUiv12z9zCk
2LZPevzbdE2JnB84LN8zSuzjU2zd/6yoS5rbZCWm87GFO9QPWhe/LvqiUFoK
XacsZ3Sc9p4ckimMm5D3r8MQbiiVMtfoi6s56PxtpmIg2bHY4nqq9X1twtnf
KehT/F1R1Rm7naMNjxfUZctDujylHkuaaQM0BaE1onPWfgz5xox2+73lZczx
3Y7IpTb9BHU3iBPZNtG9r+IYjwmutt720IWRUDsTnOhjSb42tGOKMVO/FmdC
WxR/u55pg0NyPCZwMkecaz+cEJgKKJzTGyg3E0z6d7UpFq6m1LgTWiFnN469
Q+TgVY4uChWpLOTxL2oAbVIe0chRwAvEgi26QsrjElWoXMMgGawb5NKKyD+x
gIb8lrnI7JGuoCJ1M3pkTyk6dDiLBJoyzk8E3CPjgODn+432Rr/E44MgrUn7
+gNGVPrB1t03qemW0TiCeGdAtW3tyAZjq7A/yiy+8iaeHNASVeUdaszvGFlN
rnw2kcTnELTHrhTIiG9/ips5vr4+izyNKzaCcP7Gt6x2igm4OIrmwXf01mb4
KlJbg4Z0Y7q5Fh5qoITkRQWAwEM+3HgPPHCKBybEGGWGN9ckh3g3xtD0V/sc
avMp9Vwoh6GS79EcF/DFN5IspJ21AQRdY9xYh7+DlTjlxnhROWPZgTg0dnF+
dX/LEoYaaLkOqFG3xI/zZnHcgjz8Hp1aSH2Qqn64ORkJ3AsPIIHSvQgQzTvg
80RPLuX1mZ/tnzR/KwgJaak04Uuzko4eH94NS1iLaHVWksMUXfT4/cW/L8+S
TNj1c/cDECV8IaTgHozPvd8vqDOWcpWLGx3XmZPxjZKbW0jfT6x2DIXgOtdl
F9t4fsc0zE+QxOwBgmA4ZJuxcqctUeFaaUaz2DSCP27QnS+jfLDuN8Pwigv/
TLAfnVBLoCdXC8R/MxdASpEUWdUU6qDzP4Xm8KZiw0VvBxt2edlNHksMYEMV
V+V3NWiwXxZ0V+9q6EQjbKSxNXDXjOdxUbJS58NC3STbGsxEzDFCn2oSDtzE
eIwsBi2bFxlXLFr2Jwqi4MbRjmWw/yJycz+ebaefiGxVE+ATSgAZrQp78/Ag
Bt6+T/uEGYw99fxkX93CPGRvyaovbZDfcJSlpLO3Tvke31fWaBVUp7m9e+6V
FTsM4w7lAa/9TCN5TN2dEMfBB3uZWyXvpt+xrebS9sXAh/BBiCknAJznKhut
k/K4+WCnHyf2VhIwuZvrVACToxr5BeYFNd8vGhPZHwywh3w81U65QvV1Hdq8
/bUCUHga2lijnFY4lioVYEDexWGB9dX25XBe+sOg11UNOODy60CZOSa87Vwx
C8gUV15mBeyYXv3SUFt2IcnRVZuesY4p0y8tqnrn9BPKz9she2JFpLcTpap8
OqtoJpTr5yB/0ImfP32fHn6uFxZ9F9MnTl2+PsSZdmN5JUxuXRyO2nZv1S7T
ejJkyMmrZERZ7mnmewySyjxs443swka3TsZLDj+JwwAMNkcbHo2Iqbwsoz2h
Ijtyy94hVi4rrbkPD42W5rkf0cWz3YlNpuKxmVm022cddr8rqKf8cb3tw6bj
I+vIRnmiodaSOgyS5r1z8Yx27ElqGmYSYauEmyWUpX/JB66SrWET0FwhkmQh
Yng+24t0JnrlTvr/42OxH7LjS2rK/NhKrREA0DlZMUTv04bzn39JfLbZpSsh
tUl1GcxbT0l9yQ2PI8QgIBMhDtFOJUmvaXAdGoXWH4in9wwe2L5NpCJXYjTz
ddELIQ6ylK50uT5wicnkXhn1eHxsaBC1LequN1V8/0FrHkaKy5umhaUopTrc
Ovxr9beHVcJcd/LO6t3fDXtDx1tocHx4Cdu9pmluJT6RtGDRG2f7V8b+rWJ5
FFwO7DJtO7fpDZD4aDlbKa69DYt/98m8PB0ZAniLiw7FmMhYCCl32RFK6EMo
NNZ/Kva6sjAGE9PIWKz5oZ7tUiliZUKxqWUfz3cchxHmvdzWhzTtDP1/H9Nm
Lwr/dKldanvTTje1tCkZeJpVvGycyG/PvujfX/suv1C+miLJus0RjAL+VJOo
L5kz8VhDwf659ijloHPaElLad93tTzXeXNNs8jB4CP1iEwZ/kXs6TU8fEgAe
ZZZRwePHEqrSBXrW2ESeo68zJ2EFEtBjVSU3W32YFmkTvEPCrJZKc7qA3NZs
iyworJJVQTqw9NC+xTDqneRQ9lDIihZ0Y51KkSK5SlyU0ch19imSyTRp+JVF
psMt9RRV29eLPAc52Ow7L+FgPD1LvQszYz7tXMKSY4Z9pmd1FNO/rsF6YHF5
c0qv5lobWqgXsqQcFlwHBXd1lUtp25+bdq2OxsMaoVknbaXe9S4vayI3vSi4
elwjWjGyLp4+sAmTHUz/Uackm5vnJHHmpkpHnzhPYLt/246dRPWsEYH+ETp/
2XjS48Jb/rGroPADWBcoWl0C4AmLi6em+bTYluvrlGEY1hKDfGXwZ1FqVRbZ
Bntoeoe+uDq4IcflBZ0YhnEUWp1PYOpw+34cj2VQNZdI8yrnDDn0+zgegXAQ
fxkl9JoU3v2Aj1RczKUd1C6EytaZ274wSHexlnntTl2gyc0CmhlQvxG6P6bj
UqUqPHO716JQKf2xHwb74NJXv4hNME7LgrNqeqymFJF9seNgzG2gRIBTnb3f
apC1220KIcst7NFrBSsmjtRclQzM8pyZ80PfdUYlaQCpMp+jZYEM5cG3X8AQ
k78BCReLpCEzdLvtcwv+l3lZbXgX8o2Pr9eb4H5qybf+32mht2VGlDp0lL8T
tuLSYBfTGa9BBDzNEc7aQdzxCpDQGBJoY0IJ6zjeu0lAM6EWCdgjZAemJLp9
ZrLZ0Hee13cAj1QujRb8TAiikhreSRtpANVtkxXRSZhKlQqrxCGNL7NsEUnp
mScrIuQY6UIiGpHCrKJqSHZX64mHPJC+97897Qfjbo2goXp2R2jEe/Sj+n2Z
yHrHHLnvaEA+fb1+ExjCngeyW9IFn8uTzUubBo8VCvt7JT9XyteKI3epaEYp
m2SLru9E8agTmWY+iRdAc58OnDpWp6MbOEBA6aeu8WQhh/qijgURsfYS0cM2
fAbP1MCVzusbnzYej0C8CYvBoVM4tgk2oyJv5EqciFUJ65Di/NPx0U+2z44U
tT5HY4eN1TsyEsmRLE99XQU1VVDI7CZ7azy2xoFLCzGONbUqLJSQun4esWep
msILRNrlmp/1Xq0Vqxu858GOl2R7IwbPeJeu3/1eQheVGQ1Ux/4aI4Ts+R6p
mciyAST35E7rSBRZB7yHmymOgsI0SG48Vt6ifRdgY7Um6ryr/JhZ9u/0mKy7
eACUOw0xTtZKh5lzqvGwmdPx2a/TgXVmFZYqnpbA3fVYHD7zMyzgeBDpitIm
UMnqS0WxQmcH4cfnvaJL0ReOgDtrAlLQErjaNxCcPNT5siyFENbPyMsd3JkF
P5GbfWWZJ33wE3X8rcg4TyBIgZgqx0NmgbB/F+g7ZKy3NBRL5NBSEijzLmFT
O5j7r4BHU90zz1Qxu6ZaHV/iC/adYVj4Ogyd79ZCYQ/WZo9RvRVfk/BUB5aq
TgR030450JcMZrQCRkfrfSmd+dwsbysYtMRoT6X/zMwFxfJsQCwK02sjCPxv
lvUH0vDEjo4DTmeMUxFQobcwRpsh4Vd5CgEzSDK44Vn9g7Mn9YYW1fGDIBat
M1WH2VsJCNcoe43f9aGUkHlsJBC9uyJUYGe/KYpxoel2IM1SkUJtaK8QdcTs
HToP41EOXnzqCDqOKb1RjTSJOhTrs71xohGxInCKIRfqSDOV049pNK+TQuNm
r/d/+AolJQ6jq1AdampXr186cUQXs0ssjwJg+f7/sg2FN31qjjndGRhsFBSz
RoKFRWejZqjU3LyqRAGPHYMQW56gIXx6Mqh56cqQocDphWVJX1PQ7ila3J7D
eCEQt0V1yR+D7rvJS0+NoDj+mkyL2NjJ31x19Tk8NCRlNAEJ2PqcojGpJze9
O65+CXM1oDP0jtQ9wRuBab3CzSMYKiDUSNSMiVoSmqBlNrtG75peWsBDFo/W
pzfSHzkTXQOg7w2MfqQd4+AS/JQvVTUuanjBgMMyhsbRTMNMcCfzrJ2oFfDw
+tTiHqy+b5SFId28TZNnuSGFtnFkiAj5AyUjFu2LhBOru7KYD5kWfUh8ZS3g
1BS9YH/MRfDF4Miu4xDX0+jguRhfV2TMXFfw7XhYGCWAdY/fIReFDlMuAmHW
IpsRyD+UFOFOoZftWlKCpmeUIyAMF8BIRZRiFFcOvMEjuZNvi1Qc/QsqAPxx
yX2KpdqpBl8Amxj8ppnRhw4fltAsuOkgpsm4HSsoWoJVDpo1E5faIxbBasKK
to/V0DnC2zEqF/V+4KarI1K0Ky/Gicf/zdiRuL1S5cvGkDuBeuTwZBCVWdhw
j5m7QbWKW8FD1iizXVH5jVL0XAdn/Fi7bcr8WqV9ulV730MIhnHmSb3c0vPV
C1QkDmheZ35Eve1LT5sKl2lxU066ZJ0f1ak3WFTRnXrH+9uTasaXKuW40t+i
meyN3TaRETSu5JHbylBHbBJmHMhu+p00eor/O9aaCtdMjHMhXTf/JsE+0E7G
cgbJd9koDBk8Cww/s+mzvDhtd7k5fz1ljRdif0iTHrrHKOHaYMULAdOcPH9N
S/pjKEHuyJ3Y80Z6YstFeP0QykfrVOVbpASB5GPxVWXA+aZbNeu4zht8n2YE
XAk65topZfsgph1SA9MtVgUopQwiFcFD7M03rk6/Vr0I8O//UDLmw3CzqejX
NB+CgGcVW5imVn17lAG4oojyWYq/ZQaPO1Uqy19FfF8Km/5kxTWYeSB/hEvp
B/UC9EN4OqBTcWcwRnO6aGMG+mXNT6280hKLLXzEPLxDBzI1amHusbclADWC
heCyKt40935YN0LLKJRZcgNJWJokW6kICEl91/GeQAzu2km3Vr57wxRpNE9n
QQgp7hOjgedrEmMOwJgqyOETgYP4bERYpKnqdqQ/ACqBMSsSCuyePniHzRTn
WHZq+T+lf4OUyM9J5cfklD+Gpwl0FXv7yPDRPwFVSsaDnW5yXNBwUpyUsXSN
EZiVLaHOXU0OaXtt0r/St0nfBZuAeotlVKsvIbzWAD++ahS5d+a8QG2H7JRk
P8RktwlFQo+9gdYcVzH2Pn4SSRjFDeNhycmNKnfxuVQrhmvI7ulOW/s/SGwe
SmMXsYYsPFqhjGa4eG0Lk0DvTzP5qx5eZ4yhz0Vz4i/OSlOgTo1NawmQLO9/
CcZHTJKzw/zdJETfgW37sfp3Y6fV+ganK8OjAvZmh3ojr022xzdcpR0Mdf4D
FumaR4gjBA7LIBc7LtUMDpMCyjz8NTT8bAKjOx/FTuZa2Fj1GWCcOujcSOyO
6N96dh3ROxF34bnrJ07tx93mZOuD89+LlACRCyG1E03JuXDQvUURepUrYY2C
UolccgcM8IYyBhxUXxlOkeRiEVYLm0cbXY4hx34mcwWFgRQHHD5thP9P7twz
MgjCcNh9XRWBe+I44v7igHUmYTHoS7dvfdBoKjaRQh4bQYwKp9HNdva27U1M
/Nh7UQQvXCLVfBjR31/cvVAqOK5AakRTSCJ783b0RqAqWc4uE9BSkuHgznfa
eX4yQ/FiLKiTzVVW8Bl+Mdi5l37zMe6FFrva4G2VS3ue/zI64i23+WP+Vx7J
Ycnxf1qX1tACp+VCLibp/sKS3YqZLIQE6+l4fKOdxKTNSawQkKTGhN7VAW5g
pr7HoxvbEEGbat5WKgeZSne3lE34J1p0gcpCO4pfB845ZbZwenxYYJduQrX/
xmx9AuxkSsaJzER0zJUYEJdm8hudO2TDcmvzJcCUGJfwyVErUCLSVgVWgU/W
I8VQN70lxBdHeQFeix1IG88s1onWwAmW6TEyAq0hKxE3DeuEG1hZQ0vQZlBx
6Zd72FMnaF+fpSFrplhAjehZo3SKnbYFML7Ls/4F852fXPMmYv+Ut/nQzlGR
G8pHQlZ0GBldzZkwVjyfckEABSyaI5WbScJbTdX8GnO7RIKaC137HHs8Vo9H
0NXMXGh0/H9D4gdRcuGUDWjzCD5u1V+9PLNixIo/WbhWMEHj/OzdhsoGpoHE
EfQMwkjxqPAZsPKQVKRw9DdKx4/rFSDzlcDDCgSJkhj+60dEBYrPv0VGMJSF
L2NFTepVbn3L2ccAFmgOtrwTSUuQO4KffrW0em94vU5jf8YFJxP7p5o/6WTL
BTf66gtFwexuJE9AVPSDxBDYpYztn8wUYD/Kj7fQ0fY0mM/7J23FZaSOqpr0
EBOs7XXq3apPQHv8OBnfXH3pfUBTs/7wvh09rqZ5042aRUaC2aj+MyZF7mdr
fjadkDISFbqIufN/Px6BBOk/lO3Km7GIw+e98txep4NEiV10Zl1rET1R4l+5
2fqMZA6/wh+kdQvNGq2HV8wybyb19ehNskQkZLvre7P2CV8NX/F+uVGTQ5fX
1+s8yKZH/cH5KqUsqvUQvKPEjVoCpKuCLjZt02F2blIjTtv2oAdL7HVNmMTs
sDawwFC9AcnasahL43BYxJIi2mlUbvejYBJ0tZHinfEtIS3BZ/WrLCTm8Rs/
yJTPZpSPThqtV/JhEtdcnJp3v5xoN5fKPcrp5MaEmSV3hIdc9X17fOin2N3U
TboQqHExGO1QZX3SHt67sezYoakoEd9Q3f24WxK+PrC9laz+hCIZ3knPCSC0
L2uElP9Xtw3H3Rj1XBoCeIqnI+Ieaa5f6PHltyrdPWrX2zFMaNujjY1mbHmq
OmfP8B6Z9D9USmonHCoREwDnbm9EOHRb0+YaAk4GmSl3kqhqfscDSpW/Qxuc
RQkjFlPCsvsfa/4hIi5NDFZG06bX0msJaLqI//ShALNEeF9mTpsvaCKbrF1I
PxtFQrA9PpCtvpdYWk4L+IRZK/fgLh+EDMABJInb8Ki3MRlaSH/j5rZ93x3E
ISiO+Tsk/qcvDYWGUqxhWprhUbMMvklxHm64949izbpa13antkpjLRBrq8u6
oNJ4dA1XmA5PYL2yKyYLc/lJ/hDKrhhPoP1HIpY/i1pq8WxokH9ep3zWJvJ/
hCEo9dlwiV8jU0TDpV5h4dunPNaQrnstca6UYNfEFVEbz1u0ydpSGNJadXQQ
QCfv+gMqDZvRqwKy3Cv75chc2QXz8EAf3eydgcV6NkS5fh+w6m9zzVmv3Zmf
sHpZzMrCHVo4J/+CXpJnY9+18ezqO/+LumvXYwRRl1Zai4M5ATzlw84BJe/X
c+jehFlTu7EGp1kXbyvxT0bZjnK+RCuE/CkSaryVD8ho8Uk32Qb7MPgulZfN
Snzke5GFsKOkvOdajZycHhDuGDFEk8FgIfc6Phpe+LT+RP0H5jPgXCZllBmc
2emzMJgMZmGe7Q+rLy6LsC46tYnZ4N07fzLn/E+wsR/NqvgZ0pRmUTCCN9va
87287+RsSinxLy1HokxLZzVWlGPFeI/01kxYsZphZic6PKXihPGA4VrcBODu
5nQpJXz+gA+Ni091BGhjrN9XvzdiZQ9D/cJQ06vS73aiEgi3opFh8e/mV296
BDTGfmOCK5/v3Yc8AFAI0s2/VE2+upbAJoKROcqqnGiQCQSsH7e/MmCIhDQT
YhK2ebhxc9ksPHmEjHWI4sT5KBouQ+Ihse1cM27rw+kq8pDixbznkQUn2wyi
QXTBoGE4q2FP+e0GWqpHW/XhKNNjU/lDEiWtx8OnTLGqTBlqIMMYje/Q7G8U
2dgNv40PQc202MmvuUFI8lBirUYpfkbYLnEjDn3wURP4feX9ZTTSVsxkHDyE
QX+/5pLB2ibcA0he1F75Jljmh4Gags7t+OcADDk/G9/t9pI40+JvASTKid/2
B7GPAWdf6LMOlNaj8SY81qeeQHbTUupAtYTMgyG2pEOGZB4pS/mdpmLW6jUj
uNi0apQ1emxh02v0bA/XyONLjzfCyEiHwpsf8VCFtzQdeZWD4Wty0NuD6PVm
G8Xtv84rtIL0k9CRU/q7JMKfn4vF8ceH+jQDvMi1BdyRXbWltmXDIytEoszE
Vu8xnhJ9p6NRI3+fuXbynmFkXvn8NNo9/WfWz8P1z1nGe3w6NrL1GBiEECn1
67DvEQZKSc45mKSypZS6eNejR+17C1FmaXjLizgIIPW9uY65A6pv/dV0imXC
76G2J2iiPhs5vgZG/gSsFEbPiCrMPUvyAJ3T0OGTLTI0TgjhAwYB7j9MYF0r
tZlxna9JE/NvbhHI396+gphWDaJjdJ5niXQyFTEYoFdWGz/uof/t2zVpBt0D
YlBEkSRm6vFo5NRP5anNqZ/8pgY+i94fd5HGs284PjiPFwmmOoYfk5tAMMtd
XHk+RaCKVV+l38FshqXU8JtXXDfmdshBDlw+2UH4s2MJfFAA/7o+qP33pX/i
xX6C+9Pyr3mxTdThcSAPNk6McTzTV+tz9GKNYrtUUChuYDbcQRygl5WhulVX
+ET1bGAnCUM00fPmMsWwCtJdhms7M3ebcD+9FSlYknFhoSdujzlLfKMP9EPD
0/u/lMN1hnRqsJtZkK9gGwWZwiCSD6uQwOKG44IqutdXN1fg+1w1t5A1Q9N7
wMz4skXLfidpiJ2X8Q9Q1LLzo6sB707L3UrXnM86S9y+JAV5LS+KJnrojK4p
/akPRLa1rXhNioHOvDR30gcriHQRaAk6/vsXmh51jye9cuYcA40suJ9TU2Gz
YRuJgsdTCd+Zs/Dkd1MCbrHmo4F0X5/P5xLvM39Ir4yuLKHevDpAZZk/UHjv
3qEH9Qiq3oKWOS+awGHCHLhmcfDt+YGXCj4X2Pz6BvWEXhXuSwq//bq9sy6P
DnFGPH9lW0GcLx7/s/2F6bWf0SMiOKJn9mB7B/IkQCalHaaX9TGW35BqiryO
xW1dBX/ThRM3LQW8iTAu66xAtX2cTKeI9aER51Qwnj7H34NXjGhV0xKnNdL2
3cWaq08yWc2hZWVMiY86dbtlulKKdeavExOY0c2cbue8qORbX8mHGS9R8Ah6
6z37HvZa4mCKoIewXJ3n1KgZQ0m7VUPTOpdreafKefJorthKmS8aq0vjSS+0
dxSZVor3P0ULDplW+0/vgW0LiUDIPHtqYipUdTgmXLWn/6qKF/gVz6esluKw
af12HrNY0u2bk1P+xYiaKPxtbEu/Wi9xFVFSOjvyXoZkw/vhPTWygP7vnif7
CycA14v/sXw8YrwtEkR9DsBnjECpeR1o2b+h61fHiIIkPc2DauxQRNCiTbdV
oPiFOmhPc//zGWcEzKh7rdv574dsQzhymbSKfpYJlQw077hlRN8qFxEE9cve
Kbvq7bdrzeRcoGL+tyu8ob1+i4//Wm2eBqE18J/UJhRLytAc3rbPjzqomk0U
2CM4LoGNx7mZjA341mIr7P/cbgfD1s/WYqbPdxJYi2Gn0vC/fLxMwYXjcMy3
VktdPoY85y138iP+/gsvpWnkwtBrN15DeQIbguXQgk8CgWDXOq+MzeTlIIg0
U8muVDX5qDcJycBGnuvyOj/wuno8/cdcifxfKv4qfPEce0GZVAWm+wTxNr1X
aJpVc9KY29ul6BO/OjbjlcukQ2AdAwqDh59DckwMbvkM/8UjiYDF/2hZkxuP
41TXM9qL8wJOY4eiEPZDm8K+9DAzdTw7dExj4QjevufOIq/BhQb+F3jmy0KJ
qGIy47L7/vvoFMXmJ5mAdnpkhqkwHnB/g3Oeb1VM7yyveD4TPsgNyV4ZDg2a
rR8HcTHh0qortvXe7ul2SOec2GXd8N6Z13yUyIByOv1NzVHjvrjsCWXTEYeZ
kfC/tETbTjSFE70T9hhgP8vjI7QnsGJVxhY7gGZZhplW0GjUEFKkj6pQDxMA
DbISb0OpeYUZaHirRkUM1makwRDEQe5uDfOrHDDcjueh8LPUWGgyvc6z28wF
WJlOPFb8RaC4HeHzeWKzjcsI8CQJ5KprrCA9jjecPOM5gCGsoXlJlN62qiB5
v6tjUQzGI78uGfG/rz62BUO7jVrGE2MvpYpMbFzH1XFPfXjkX17aMtyYDiAj
uddE+K+jPq/gUhFpfQk48n2MlBHVPpSby2LqAcuk0u889th1aTCvE+HPCdFh
yGenBRRJPUj00gZ9b9tqLzEdn8GjHq5mJn6hHP0n/L6s6zow8V1H4BBds2xf
UrwEX0h2HUCvIXX5wewF6Kgawci2F8hF1SoNPQ0HssposPRdLHXP6ZGKE2CV
klFXmS6r8rKkPGOj3rtVlOIASSA1axF8O9tbfpvZve8bRlvB/IZ9BMjkVpro
C6xvKM6GtusNQJwZTGhpgI8+BodeGncSF6CrwkswS49bN8LpU+dZZuT49vZ0
Vx/08Ox9rcnE0R93L8zzR48AEzlPKNZuZ1twvP+lhP9yiPJ6Xh+r4FmP5iWS
4UrvRjrhqNQiCaKtaagOLJqc+hC5/h47lvQii+GtGcDfiMD7IW3wVknnNc4w
sLPO6LHAm6TzYuppm8HPJXO0/wRp3pt+ZuvQtYAtFD9jtnYGoefT5O3oamni
cqaIo+FeBfzWo7qD4goeyTwJ0Go2TInOqtnJRmA8v+V9F1DLLJxpLmH1oQ04
hjUANAmfwJCPq204lrMUsmmrG8FC2Js4Av6+vT700S6X4wrdmgW1C5pRokEA
zvIy9Vf1w+I+gU9mzOS8AxI8xOjYFeyugUGyP7KrjgSR4ajwcQw1FbX1WNSA
2ygOLeEYFyKNxhLB9dbL9r3NhLXXsj+11LLeFPQErNmEQ+dnQ9g46+Nb2fdm
bEDTmtW84RCPDNhXhIJ6SASvSI88AIS0bpES/QLHtTkipd2mzKs7mVC5ZVvY
TGj1AuHd+GEtggleMDg7K5zfAXVoVY5YQblFpuVLYm5n8xbCeIV7S5aBGGIU
yxWQ6LqfAPe/8qxwIPmvQyYphQ+LzpcH3gRj3IvUSg3Pl7XS7EH2jaDQG4vZ
H7rLRpz1eC7kEt0xGGYT5Bjd9u/yClrmbwx6HO0RSXesiVmaTSpjFiV9Egrl
v+gkrLydhHueQzTaYoCfcYdCKXL5BV8IHqQnxBn1dSIY71Ez4yTIvzUsFmyM
4fo47oLYASgCzHP4Oai/9IftLngk2QX4QJhSxcEcOnEuO4IETSyOT+SiR4Sj
Iw/j5/+bT7TV2Cr8lQGGxyiAa0ecB3HzJLWjYZokJomTV9bhQKnCrDUfaF5/
nFNenjPLsBAIZDy0q6ahEqHQ6lHe5fXDobYAGqZ5Oe/q/qyjzWqsiEDtu1wl
/hTBCjwsvGJy+jzoVP58EF8WOeb9auIU7w+zYB/FW3Ns5mg1A97+hqnYf2Px
ceH2xDhIYFQhHhZvELSL0tHl6qctdNr7fhtA15L7jsjfOq320cmMcDmGuTh8
PPM00mq50RO5fIawJTf/e7R3h+xANcgn+DBLI5WDJfwjNQaaUxxbX6x488Jf
QG0eWiHpSgUSrY77VjNy25P4oEHiKK50GQJY4E6Od0L4M2slJwr1Dh0Vo6lF
UTDMQXbiUK4eo6Z4vaC3bSIrfLYAZmRGrSLOg4odbiuCw9PwRx2eCjsD1SI/
IyVJ/0kZAmeJIvRGstv1qNBEDyjUEsxMyjlnWDKj52ZZp/9D+oWOreL9rQNs
2oYQ3JvBEogDS6zskqNg4iPwT2lfur0Kmssk5f1iCOOaYCeYRJUt4nkPz+zc
9XQig1+vZqBPQ71CuhLT1vboJpA6tC2h9axGODRkrs2vkx8oOtK224VFd1Qg
nqt/idzJZMO/MsjhKlTxqHmoKL0e4KScYJ+Qv61n2YIJy6WctXw3mvvq1ZS4
S0BAdoSzALDS2WxLnHVNIbUQjHN0mIJT6z8FukM3QWw9ge4KMe9nD42ySSVa
jGFMQ1n/2vckm4EfkaBXBIi6VZMD4KLk/iWR4VyTomojctUrkC4NNWVc9MWp
cs4q8iPy/6SW/F1ZfcaUQFIoMXmgZAo34PQoliH0GdBwSs2P5M2Pcz0LSZv+
nW+WVzY92i9sMyh/KJmDqorg6P3ACQHeu6fQY+Fmw2koIsJiV4yggJfHRPLA
+11op9sQ3dROEE6GW+Lgq1S+7LerF7eVeua2DMUzydBUneCsAWk96Mrcj1WH
xH4Mi9LAxRg0jlUyKnh/Xc3XDXoAf1zVuQDXX4RGi7Fl7KIP1kaIeKSUxbl2
lGWHB5DMx0J/O1EqiclzdNoBKLAvapKxgOTfrl4ldxc4TSdccPqNdiAshi5D
HI2+2LxD72shzQLc1DEMfmnDSLW515i3o+gn6NDeeGeGD1PO4kvc4uovXBcR
TDFQeP2MQykoR+zE4W6dS2ZNbxzptaEd86MkGm3Rakf7OZxk8W6ZszlFvl3j
2najhJJDw1/xII7zHnr+gms7kVYsKUXo9Vnj+wnK4vUTaAk5N8PE9+E4noI6
tHPdRv6U2eyfu5gfLY5rHTFOaOIIfKHXNbc4zagx7DQveqe7l24BKYS+vNlF
clH9XxHFm0im2OVhAVF8Qv2lJh1h/Ar7PuVDLAU8yT+CC1dswh22c6Gnc2Dx
j/wyY37lplDiyuMjkNVOWQEj9z4BFn5vQdYG2vk/qrBrtz2fmQKUN7abmfmK
peK66AyfUew6vBvgHnTVoR99JOBGJtFOMWwjtZIFs1b7IpiVrwrKGcxaZRzV
nTO9TiaeeoiZscr2/wfvjK7fNSslHAiPVKpKhuTUftla/uP4m5ciRLHQCLaa
f2GOIXX+Bc9Cl2oPALjIpy/xy5Rs8b1ilfPsfIunX9Y0XU8t4I9ExP9ORHlM
y9jsvAAjjcAXlWPQlQSsBuQV497iQatz92SrFIft/iGJemg0nroDW86Z90Xv
jidIt+lBS4DFDfrCFWe33lamTieXZyCnlTzYGCDwMJ+ZnaCGMPxahcopl2Oq
Q+4ZRF0yd9NFBG5ufvT0ogy4awYTJ+5O4dz0FkkuhRG10rFclliS82HXogY/
SM6GnNP4sIUCq+UK+Rv96MK8OQ+MZav2DbCl54tfvWIjQK+Mo4pzt+0HIg8X
gEH669GcWu+EXD/TlE4rOQKY3arwJa++TpiJpJN7HdfZY9a24jrpBZqhV+Zk
FbZzktJflYYgl2DRz1dupE1KDEndwnOnsLqteXlOeoPXsyLfO7dN4GKolFe7
WkvlsleqQ/30fNi9EOyjQdc0Vnb1aE2IGulM7NlgPz06eqRWExqq4RrW0IOI
RhrUuR2UVTgaLeEYhjvI44xQd4dbwrosV/HCtVm0TCIkSQ0cKBb02XkygMKk
Wa6p4ft0BNUSvEJEpl6j4gSm4HKAtH0Ao/qOQWmOnbDgDazq4NPVgsLtW7/t
PxoHReolHdLpKfYjqgBm9xQC9Sd78e+wftAEwTpJybTggQBJxSzrxjmlwfNc
8ZAr+FnKt/HDOlzlbxhTHU61o7NghxbEqOgCw8pMXpXHFUTue8E1tvpQbpaU
9JR2bVC0S/Yh5tQyApiPGD/1ppdzeI6udMz3NxICbijk34QFmRi9KcNSagds
sM5wAJeePopFkQ1XSpfiikk5Qo8PAx8g+j+XOnGRgplc/3FxPEnP6zXknRBR
2LWaPLDINpB6MiRnCtYwJxouxyTeGGXpubaFcemVhMLYymu9gJgUKUJUwXzY
a8zea2hhYqEYjY7q97m4oMOTS4cCZ8kS+IZ5RuJGmWz4NMHEr3gTKoxDnvwy
dXeBHUOXaX5XGy0eAaTPnWdpewNZ6zI5k4A2SPscL13A8MJanWovE+Mg140z
i1I1NDsriA5aHhw+bhYGqe2ADK2qkT9TzGoxKXbkxLpMX4PIxOcNu8IFZW6/
WO89aenE1vVos6MXvrWFBDn+74W/37BU6/PYm33KYH+puQIPcZSPD5qKSAnu
wyq/ZMZlhzTYWwXE5AV5MToQB4Bf7DyJ3+Byq7bana1DOZOMxke8xVW7VkHN
L3QoJW4FzV6I04WE+kcSx1UkmT8E3wP6s8qLLWymeb86aSjdmJ45sL12VjKJ
lpEtcJR3+7X6gQAOZihle8raPJWdcoRTwupUsrbSov1iMxC/z4vMLYVwuYTJ
YpeeFEeqTvuwpgPmi2pn6AHqXBbHf/syxlbG2fhFKac4r3+mbpQEqPGaNcNr
iq8ujlos9VPW3Ej9ZkAP5rpcL402G4DP0VejI1p/5TgS0B95PUrBrNoC6HoD
JdSVrS8F7FCKedQXJbH2y1rXbpm10SSqay/jtoHAdTE2zbJNGJqcGizaFWj3
MWCqIDPEmdFjjj4URuzGbDlLQzuq8RLie9C2XO09I4cTvcUdOsmmdLgYMTzb
vJ0GP0T84Zl9syK4eU2saulS3PSNvpIVC0WvGuh5lklzpCNwGS/7c/4dPgM8
rk0+XNggVN02EUdi4TSWIM6gyXaeiE0W+yZk3pW2h892L/AdP/OreyKTFIly
mtkuFN2wvi6zd0MLjadLvfQbfA911Cm1nyKJOjFlXYsMzL+EFykKmzN6jQIh
s70TB4sMfTlR1byeU541CKPiQl+f6wOcb+u31+OcMvul+724B6ibuzVTCH9T
upWzfV41ALn7EfxxUjJ/OA7ksoFT1LPmFQDEuh1wZrczn0zBOwMQxJOS/BNV
4Zs5tOewYBfzevKe5jjbbNZ5qGTDXZGiDcIpiJksfB+kg5iPDsMwTS2SpCsf
NxEnivTaxTecwfpeAzhiIu7HbF6BhMAWgU5R5MmB+keV56cQuSJd5f4qYHdr
c4LIdMAc5OFpMRPc+PyjTdIW14PpYDFxmSd4agIxdhFsGQl7cwQ1Yc2DVntx
1xhe2DSu9gL0BN8dsT5wgZY54Db6gZikriOOE3A2J9IxIsBz4tczv72Dz8U4
1LrxbMNzq8FHtyrwplxZmhbRJsm1P0dp5X+YLnzLabW+4wkTe7frN6YI4SN+
Dqb+gV7PvdjuYWxZksFJbA7NhDCqMzKBAErxFbu+GhdDr9mbTjeXxSm4I/Wm
0n5/sg5MYHKE5DOfq0zBJzOJsYGz7R3Rjs7d09wrM2mhGisnZy4+sTORntzA
AteXmIWryk3LD0ZK8B6xhAXTtEmZ1cgwD6LTeWvjJItfMO8vtLFeNltD6pgt
GOPmv/MGCSOgWwGfYTrgc00LG6JXSYLKCTAGVlIEYsMrj+6j8lmAf6EJmFIt
m1kYZEmzycailUiLhUnCGBQWK7SZynpqsI1+km+VqzpPvMo3uNMHJF9TUu1j
g+s7ihb4O9WKihxq+RSgHm5FVqJ2Hy0hm222mfWo3tMjm3FDTOfYkjI6w/ed
qw4FLJLpmNKiNETbmDtsvFKCwOwhQTkvPHc8JW/jx7YK/HYI2+RUGgw9hGWQ
4W6g8l1ucgSsfuMbSPwIuA8DFE4FUflPLQL5CWeUVdZ0qSjmafDcUGROAsuT
8nzZViekYkfAeKggWEaE6yCemFzbF9fLeMk0/bDctN8mgKezhd30jeG0F6oO
M8fFXkFjFtDVxXIcC4pNfEmgTRJMTxPjLbhFi9n/i2zR+7tqRC+CxfVnSjbp
BS80VpxmYytJ2q0Ygz99XCjmz5zw/BfcWjdGODDDIl9LbP8fwW99YsghmhWG
+InQFTox93cqrm3ia+6E5ODdPOQr9Ljs0o4HxFFaHVU029IAtJ+abKweMagK
H4QWsfBIxbOpqqXKf7cJ4DGAkhGA6UsIkdxZwr1uC2ilgwIUeUjDSzd/Dhtp
NXflAPx0yA4ZuvSms9OH/xJTqo8qQQr39f7IHtgS0avPzwR+5K6uHs0sWBgv
AvjmnfcWNMyABcAfvQb/OKpFlHtp5PuE9v9O6fy9ZyF5HRAGMabvCQLnarcq
RneyQ2nDKVDHCHnxzb6/HhHv4VFsvPNuXVStzSC2lraVNBZ5B4sk8OHxQnq/
f1cwTUmIkCRcL5fEiO9zYMsnkQB+m1461E9CTcY710bZ1TWM+/Ek7NBoIFtI
2s2smLu3AIjotlES7GtJcPHPp50W2hV9N2no6zOTeDKah0nqVe906HdMEN4A
XpZB2lYd5tR5ExNjMpTGD935YzkhBSrZh7lnrifY1dztZZPdaOnN7V13qk0d
E8dcnqZkhrlMGb6qPMPFY0TBqw5qZtI8G9njAJedUszcXmHDa939ce4qTkEY
QMNukWzGaH4Dm0osXWlPsMm8CCPc4ul69ftywBfZZ0wyZ2SUEDOfwIps3u9j
24aSd4DQySr5PQ4UfMQ9sJrf2ZwddrurpCZLOiXq2XePnXuStCSlpCxsNCht
T3vRFxsgfFeJuRvsVCw2yXlDYhzpGRfYBp7wxANWgVhERz0i20gdTKH9q1Bd
HJSlfQR7uvTZfasqNWsJ9eS3pElogYaCEbkOiR04CdF8235524ZF0v38MydN
M5DUtQSnXtf0m8Hgae2jPjNPGwdbC9ZniNDjIvw8KVmNBycw4sibdREyj8m0
vdXR1+bM+Ji4jEpFqRbqkqsupkc4YqAlKy57a5baVpb8MPyxzolhQX91GRYY
7qZRwzVZT46VuKUJ/7cc+DjjByYW3NPDP9nRanVk5RFWD27U2SbfvDQkRQ6h
v1Pw2xiNb5RLcAo6ChgQOHTzw9+NNsTWAuachVe8uEILxu1cSvchaPeTEmLm
xh6kB+h1OXPcaSIR8CiEGpzeIkqe1jdxCUizGAYDi58OsfFa7SLN5g9KVitS
DLiMBz9vBgwAw0EOLD06q+xQCOVkeKppnP8gpMNVpW4QLo7WxSshSpI144Er
YwOhzMXKHfoGXOIKIZws3/TmW+GcZO+j3EvZViGoYcM3eDJ+m/UjVvGHMKzF
0OCbA1ND+QZquDQ0ZfkmbrL//aXUI337ImkvS0mc3omXr9unxiLUIDMB1I/F
wDqFCJz3+Oe1l3aIHUufmGEhRXbQC/I4EvsaDdasLJoZWLUNWnZGj7rHWcFT
NwD9uyJ1A1a7ROc88bNCdfWFOg6tfBCFGOHh7dE7i8VYf2wyVr9z2p7V0HLK
jXd7Lm4WNs7VhUU5PLJkWI4LxPiVaPrS2gd46riCbzsy2yZTfEi22VIqn/vI
A0g08C2s+lXvYm33CwvGeKAZd28QKy0w7QsxbR8Yb8J4+tl0guUkZC3LY373
2Vhi7Op6gSAbato3WYKbOR+O4xXRdbyS7P09+UKnLJiN5/lQv2RuuTC8Tf7R
7Cp+tkUVvf6eOUQ6T3N2LuxRg3nsbBuRDgqh4y8KnBvmUPQRLRFq2N19KgZL
D0ZUj8qJiYHjTzs+88rJ/gyq1la7CpFmQAJdT+AClcJBGCsyvB6jYXbNYOFf
pi0D08fVgnFXyoy65iNq2nJCDRu66KcoIHdu26CwdevgQ6MI0KXDlkopZsgh
MM9cawh0qPUPNE8cyt0H/hmXx47Yv4wsfxYqXYCIbNHBIRG64bpedw+CuwAn
5VtYw6qAc0zGDaRk37QUHv0ZhzzxErwh43CuMN4G2opDAOlMS3qGPhe0j85n
Z64XynzPcdRFyuMiT+ZkO5BIx0mduBBS0W62OBSn+pPcapmDoKKkMXhdefCi
JfZm3SE1NihBLNwTzFRrbApiXRPFVM3MlemKL7P0yis2jZ12Vc5YY1vBZ3I4
QkXkbzVM18qcIf8K0XTlHLR4ole3Ywy7MmAW/+ceufVe/Sjc/Z/I5gKNirNT
CWGqHxrzrs5158qfNq/dYq2u9hZlgEOuJ29LQoJBaqmklGaggMeZGcbpkw3S
OF10bJhXdzBDDXLroPpf2OagLrybgzvApvkFjPEIUMndNd8kzjQzkQmNSqIs
TTPWP2wZZSzJJ+uCkEhWi7DA78TpswoNbft1TTKGdsojRqJBKZ2UiURe9V7A
U3gekIJki1EvyZo6Za4+2zN6WRx/zQGwVclIFxvIj45y/5+WfgUs5BU6gNeE
I0Jy0/NeCpcXT97DM87wJ4ObaTBgYFuZNNrCvWzytfC8ZO2fyC0lvQcOMU8U
HHyz17cGf0BgfrMmMkb42m1tdEqlpmbx0KhRcewD55g/xXOzF7h3c8dY+PEZ
hJqt4UAp82zHrVgmjizy0hz9GPtG1UIFQoN0Xq08TiPjMEpTscrieN4mvlko
3qdfW8xVWKrVLQhwU18SBJkGtm33bfID3sw9tEf9LCZ+rSNq2+l9XM0ySUYF
bGJtHApizdDZwYhsSqJbeNpDa5vUPeOSyWZsAtfxoDG6ZRbML4xt+LSSxjFq
f+nWufTd6Sp/zZTsw54fRCZT8qAdjAdhGvaCtW2iPhkHJRX4Zl+LFNBl2pru
DywHazrgdzQISk7Rhxnv15IpDe/4TjmaW9zX+DBT/grIfTUazIrpTuq6oi9n
j/zOfft1zoqpCQiTlWUOTZIqFK/1HDBhzneFekvsoCNpsdA/trPrIbzN8X8t
yGv0mA50g93Wjc4Gou0VYie1CJYMAm7Sp04E/GTon5QZvbWJp/BCxmTGNrc2
jNTdp0+Cfz1XNeXtLiKEwugPtF+91qPStEoK1TZsSlhIuePzZbUdZxgGivD9
X5rWnNqZL0cWG0jdR0kFybZHSrHyyMTUzJEam4+732wv4gdtjDRgyCEOVjes
o/nOE6eaqtXJpk9yExh8smbIsNFPKuvc8GIfemeM+fkMifNjQgaNWax4EbmO
yWVCNtl4GpEuVQm1442ohVO3j1ydv3leRUXBBDRcTnF+qwbbBgs/7G4RxUnK
zz6BEJt29J5TJMrulzED8RD2gxl5YaoO/muJ4uWsjYW/x5XTqX3Z1RmAUSE3
r3SvjYbqzvabTSzf7N0Mk88hHFIb12MHDHvNm3WDDnHCiNK42OvdK0s8OXoW
pftx895wWxLe87JvYYIoWZCJK1Y2yGGIRcnEPYt0mwI0J4bbYd04mLirDiV1
DF+5dWB3Et1m7gfrvRDHHdeOQ1d+Qz1zlew+wJTBoqV3M+FXwjuvxdchh2tg
6uAbW5OfRRz78XNA8wcF8bmMWKv/JeGCMOiJbDXCq85ODMajZxWIHMTp2SEa
7yn1E2v8RYZxKa7FU0D4HMkR87gYIF6H65uwsStFs0709h7ENCtM5FhI8H+G
UQUQKftGKe1XRJFqHGyni3IGcFjCchbXK6jU4QfpPS7a6D69OgQpMDbxyHbc
3Q/xg0/IzWy2eM5Gh2R2uHC30k0614S6NDdqIepmXm26d0RioTPt4WJjBlyv
t/q/3TPgMYC77fn4FSwvCOFAJgD6NavlpcGbaeQA/b2fkxUtHb8cYBYmbb7N
JU+Qlgsgyzfgj6cXUCQFVd9IB0d7ApA8gmdLisUsVXyyjL/YE/DpD9bC+okP
4a2iYmA0Ia+IrOfd5L/eNa18uc+kLEezwGP466Z1dn4Q6sv4FK9hsUgxrQHp
QQsHfGYYW8FHePyyj8M61dkz8bMJ622IYHXj8X+m/0BDnLUIkz0kdbBl5hF0
Tn4mhjG+Nm0y0GTF/SyoPOyR6svW7/Only0B5pt3y/gRpo2TYY8JfqvIwAZT
2eUEjtcrKHAHkQBbBczEpI2my04AtedJ/BtnKUyJdP70acpCpV53q9o75iAb
6LNkTI5IOEbCPM3DRKxeFoH6Zcsg7xnqWp9q8ZriFiaChHDcEUyZWdq7WiOp
Ql8jnkTWrrHvqnpfJsFezyzT2Y5bfP32geD88TmLXsTQ10zevtiH5f5xVhpp
U4xGJzOo64xmvA1sZunNuGlxVxxQMMJXGZVW6MA0i+eiGaXSkgmQPg/3Etus
cAy7s9Zel7MuNgaMQ88AeH+naf8BBw017kkaCbTxeHjm3a0MXPVmCYRNpE5A
LjCWmvXqeRXsIvkYPzDMz/RfCFJxSsgemxJkIPn+xlVwwp7a8SqF58L2aqre
DdV1vyseTJNPtdIrHFB01RPdhL6p1y5i64s61UIRR8wy79cv85d2mPaDBeWk
Ttpi74JNmt/igTIobj7FML5CymPWspzO1VORsU+EiJXW/eo/PwkFfAUVAguI
1jL5FM8t7zUaUm6K1IDNj6c1eg3CSkBsIg3QmBj/9U3X4vYCjaEeoqwfIluP
17BO2qnqH42R4eVw1/ghfR048se/gQOJ0EYuB3559cQsMGYJxW4MjK9dWIu/
tuRsTxHNDPfWBvTU5rcFyyUpZwJt3einWqn2Pvz/YKB9kwEscUyqetCFN+uj
EQgr6Gqufoq1DTB46yrPqwcqFjwD1hpwYvIiVdPXIn7vVBbYgEqMWNCoD9Zq
2Sx75dDsV8PiBm0KSdRFpbRfUdEIf7QA4gv95ZPBye44bjvrkpKPZ9xNtj28
xAC+xehYi8HIUOuXFihFCItkIyU7gBxLWrpx5qgwD6sScWpG0DkryIHD0OCM
y7N9BI8Nw7RP2rRjE1Cjsv10T+p9l9n2BI4IYkT60m1s+T3LjYsvW3DpdsXA
3DMKYqwIYBSV5wnJMSJtT8GAmzAnS1JvIanz05cjpVpTyr936JdviBY2bCMG
eXwz7a+svtpIvR6wnWG5JQGz0FMZ9i25MrPGRYgvwEjk8XkhA1ZLAoIEeUDj
SBbXXrvKcfAXkaJK5pAVeLEXQNWQoCCWgFi6zO+2xH3sMUfkdWlDN7d6cKxl
wOJ8/E9+mNEUSSy+FETvLwCMYolRUyucCRivePvnd1REfttE49JjeREXafrp
UXddoQbDP3K3+FQUCc4yhsf2ap2qfHtYXnk+nUdQBnlXhUHZffwrkQz/tSTK
O6oXZxQ1aQC6PPgkh77rH80OiHGIzCuIx9mgb23GqgJXy+dKqrkzl+O2LsKB
dhUf77z9Ld5TtzRgWKg64nJzFEiIrIRUmCytjb1xNHQxcoX9/00jtFr3p6G/
0N6oG+06Y2lH3c5YEotCLdNGYqelaYkqLkoQg+c1bFePkHDVg3VDJskhEeyz
9xcdTXE0K6NI2+TqIA7w8+iVaJQtMCz3su241ZrLvPeemCUbZCFCZ2Niwk/L
FcCoReFEsEitBymmQMHEQ5cavbiPiaizLGy1HXPlY1cMfKG74aev5xyNF9sd
7TMIxquW/uEb6IGgGee2bJPVCvcpqLwF4clGmk11GoZRW5eOKGo3GsTmLAv8
9RQGawF/V/Hq7AyD88iGajCft1F/L4OqKifR4msOYHnG6jAlo7N0oawxV4mk
/eoW3121SDz0F3lHINQT2M77aUqGpsf7V5EcYmv80IH4FtJ+LSNUZpvW/7K6
gOfKm00bhwt8Wpnv9NhXU4DXgALWR97x2s0JdK8EOhfKDO/ZnfsmTHDb3S/6
E5GG7wEcwAAPvXNpAkDDD88+R+mnsWwNpZN2ykOhpdpWngcaiWBuKTcTjRYX
cMPZgfVcvdmY92g8siQHjsFzqZ9uXmssI/oJtEE3q8sVXFKDxMGEPdARjLun
gIT+lGogLT+RBKc/X3NTadexE33bSQUQQgwExhyTapPSAuQzh0pmyCPqOsuT
q3utQQSI94SdcZyNlsUKyaHbaGaLMrfbLW2qXDSFyX9MCSHRbWfmYyHxBFjZ
GzDqRKgntHhBKv2DvaoTpBBejeDpHiQ3NXfr3dwAEdjWaFZcCT1NQ9W6wDXV
b5M/rMEh6WUdbeEDaj0wH3zkNINXNR2BoO6dK5KLE7qfXy/RCikktr58BGsf
JQekE7fBtI3uXL0nZ3kePho20hy6aF82sPxXxKpH0S5RmzA1SbFpDJRI6++m
g+Vx9sbykTHUcnnA8a2C+peLFkYsuvB5vtIuAQSiyisC20MnY1AfFQboS/hO
zpZifqV0T4E2EctoFg/vyIJAvfAbUG7k2r+vLGlzFELFKEu8SFkBynpbRVHU
z1OFP6TfgA3bQ4VYeV/39Z/ASLCta8IV8CdBDd/6KAmOAe/tOeQwC3WoMsxK
j/J4Bb+k2wBOyPXAWMGqBTcEkA8Eof2+UVDjEpjtmqp+0ny4OhoNbl/O1N2C
QYVC/9gC6Iq4mV6zkpFWk6FTsqiCsBV2NCCurhWX2+HoAVhrUmt2hIh45UQA
CwWhNm0pN+GcpDn/J/pCjwTn+YyFOyYYsbJhDjQADiqKqZVuYT+rV6Kj3JWo
0aACVjIHJoCM+qtZosdHqtyG+zCrbkNyxrmQYELKY+q+j+KE/+CwXiiWoMhc
eXNoVk5U+RgnJWMzcSzsJSKLH2XRA8/onUrjYYKe5HtVT5iKC3otG4QEDU0C
ljt/R2LJRg/R03upuBzQBMOodY1/WUrHYL+MjtPLnJxR9xdvVJCPDiabYJeo
gKQc2feO+KpsBQeyCsPLlwglACLICx4Nb9BVHYfMkn1ExLkyuDG7ffMUoJsm
qZ6cFN5gmZGK+hXUztagzfwXX0bul+uLqd0lA0NPmMo/WF0N/IC/Y4OE9JzD
do6qEU+yoU5xa5NCH27JzIp875VsW7YM2hZFO0YbwGK8Zk7DlL0OI/Lc/hH+
MBgqok5MaixkD5pGNX7jJ5iBlsF4JL9AvEhHvGLMcsuA4gQ0iPVyLhrVMIcy
WFulHXk9xO5iGgJqa2W22AM12eOsEjMupkF4ksNwhOjsZPQJfX8TIEEqFegj
gbzRb/OmvYEnP6l+hO6etWC1rndYzaBZszcJw19OMEcf10dUPfoDGLXGy8w3
HwzvYG7uYxJtS860SGa3QSypdQORwOBWSBE3FEMV322l497eSsHKzxn6zbuk
CH5mgA5Ou/DYZXjoO7ZGTBaZAESCZdkMIHHvNdkihIZCpyMroqmTyjiYkXMQ
Ik/5s8M+i1e8QJpyXI6aYCdZjvq98AaXJm0t7Ir8WOrT0oZsen0vjF+Bi25M
zbk8lGtdsv5FvcuhzToppa7TRAEcsWneqoRLtSdLDmSVjzdJqjGPALd6eC5Y
de0JCJ6jy/3NlmsSJMR41l3lyP2HihQ++NcM8zCds5ylra1FAL4SbJffzrb9
SFAvg++qtCJ+aQFMUOglIz7Z4YtBQ2BlmXb+Vqfp1VpXhGU6ACcshlE5y35w
oecwOTYAe3In86NLMVF4dn9DXSfdiyN8lKqfjSUykKmo/ZEEflS2s/qc3lSI
nXAdEFlRW/zLLivQ7sXOuJj6KTfhtftGP/g/cPU3N4mjS7+EDLu+uM7U+iGd
b5XSNu47QFwyXKpXNmf/GPxLR1vT8dHwupENSllcAfqLnYSy26o5jFyV32br
8M1cgzjTytxwiyn+G85b6y3zeVxzZ0L/TOX/WxwQSMeD3Fa1xS1d0vbHrGOs
Mc+bwsjUVSrXs1fj0n4EFw80eZud4lN86YB+YXO1qfXgzi6JqpPjJJrkHcqY
bNkDhlhpY9agiuWqzaBnnZGbb0kN7P5+XcqXeVoqPnKGxgWmzCEUmXErBzcU
lm0eknxcvoKlf4WZ9TWWeaHG/xjhjRe1MCMMMthHH/KbEbLZx+3YVsOM7zGK
DS1E20/MZGOIaYGBnkszfX0UAcBVlPuWffNsMY/pyQOjJgMeKxolo8zwAaU7
oPf0p3WlGRzMLN3TiWXTM/HX4mC+kCOINHx0FKI8V096nYVMIInCLmrfR6gP
V9eC8Ac773Uk9D0pQ3JAIxmAJ6huGqawkwhAHpNY0ymnFUTXwtlkZxnRPPAB
NBlh9Kzoea5Pu8w4wVDcbTEcudsgEM/Fg0qvdeueBPzbzv66+u72URp1aVDr
aRQDBogaKmcFuJ92QjIEMzlIH0Nbdey+qelinnh0zWNkFaGBISJ4YTEtgisY
KVHFSEAia3ZsFlSpUVnWNx2y21M594J2pVTjvHPW3zTvmtLDREzSnhgOXuB1
nARZ56lDVQ/k4Uajd8ie9Gvbrv3acgGb0TrMrSndGf5aRDSoUvLY8nKCEYYu
evCy0vCFSF3v87pEihdc22YkSQJfHdYafhN4HEJMKp8K23nVpAbT6Wld4XS4
tucg4v8S51kuFntkVivtmVZf82hdvO6K53q3Gh3jMBiDM3BFaC/NVtNciVHi
fpuTf882su9eFXG9XfsOcwHkD9/eyOjbGq3Za+2OdOpfwDX0WCC/TvPqscJn
QALBQq7pW4pLSslYIWhSOB2/vjkvJ269VMwP7/7pWjNGlr6iDZQw63GtHY0A
YaZk75XIcYxgrGYTbv9xJJhkRw1T4atGXIhX9+SSeCeSmEzK0/ZxUo9PWZZQ
+4P9QI+6ceVcaUJZekDbFe7/qPab/4vl5S4JYLBxjCudh3On+iBcK0EPXNb0
Y0t4skNPixEvYHpRfMXbBc+XANUWNZAReXxdwd+k9QXoCqE+SdWVgxLhRGoY
f7VkfTlpLmCDNxoCykN4CAxUUJqZAF9ChyaJFBhgQM3gwbwL+MSnEMIN3Dv1
cXXMoR7ShpJF7jNRwYEG3FaOAO1ocdxdxfs9nu+/l0iW0ACHr2MFhb/ARsaf
XbHyLHrmN6icCquFm9mFxpuyNVwH4iwKPT5mxSKD1jpLHVJtEp4fiRxQnD8b
AYo/RQrRTrYLVfB68aK3Z7xEe9GxiU0bxPKFwDFtjVoLFcRRTZMFhtbxCCbK
keXYvCigs8c43XNjESp4zjs2/JE23X4dwSQr/bKb9HCWj8/xFP+FGOCWbgf9
3R/gOVVBzuKqghRTrT7VLFB0xbPQxvPwh6RPmMYdmuzRoV3VJE3O1twMDK0w
as9DQf0DhyfI5DvJFaMfgjvZ87re1uLfzdLhjtMBsQ0B9fvBS3cler5JoHwT
k0AKDHMYljGsjqsOR1Gbp3FhyFToPy+cx0Wh1pxCIL6N8SbRCkRbp286UFG+
OIdoMa/lAuSxTTFd87wzBQhVT5Sdj2D3g5XIJ2KozjSBrlUIrNclaa95Dz4X
jtUd82K/0hpnQenOpVIv4trjOgsQ/4LrJH2LFsOJ7O9dytVNtJmBCSaae+Cv
aFFPLOrwBSizrrpwWNB8bXSUPaY7O5KpDfhe6nfbP70hQ03fyNMXE4StQ6m+
2UTBuoChDQ+KPwblo3u8T9qNEK5w/jlT9aRypV8sHIUMW891swMkcR6VDUnn
5unJ6vJCxTtfrCQ4qW6uIATJjYyNQJLyTqaG2CSMkZPOWjN+qTM3njobtgMl
7JdLj6fNyrAM6Yrj6i7WtvhxsyIu0e/unsQGu6XlWBt1YtVIi/sg0Ousq/3C
Kq1lfvVCM56MwJ1XZn5mhGVXXwEEKnq5VYHfs9y5OaKMb+t3o+J/xnFMiKJh
G/bqctUEUJYnlTymeVztSVj2mK69KHifkS2m5yTdFuBlKGx/8zdP9Jco8kjL
2EcAuo2WIGDm5ddIrY5QgTs5ts0LMdgxymjwJ7OYhJpjTQ7M+eh5s2t8IJE+
w5xi31jY+dK2mdMXwWwMFKjT65i9r1JNWESHKuM+juKVrxbsDB/meOARnIni
IKoZy5l/Q502UuZnrifq++bAmLYRf+H9yBtCt/R1m2fzJrOzDMOjR1jSHq/A
PAQeLp3Urcd5TyKRWdz4frj4xoAGGbRBcjpsvFvfrCOKMOc+b1uxiK6w/eei
RF57w6tLX0nx/C44YGWvMogTMy1GBmxWOR5dB9/Z7G/bFnalh4XzuTwSRdlb
v1jcQ2D/AqED9YGXE0jVO4CKr2zJqhg3a7I4NZwya6OJygnLxbsctIkhPluN
ngwmAKDgAmxVFWMLbAil5GKahxR7mxJnnYpLiuLzWkjBt7TYfvQ/6lT3773U
PecU0BcRw+4F6UqMyBrwGWrheT/027DoHyeKMjpnPUoSHj8H1V18sIfzg6lY
vn96Z1BxJNmx1i3aPeCcuQGInJPEAMEUdelDPRO/pEqMxBNlKtH6+/QOGJOo
aITegvSKCarWr50WfHXnyve9z3B9/28rO/Db+HeIFzyJNcbhAY7tTsD+ZaOr
rQDeBkxa1/rJo9HMKouZMKGKHDNr4HtjAsW042EndZ35Zu8aRA3CYtfTc0J6
6Ia0hran2/PD82ZWZn1Ef7nmGzxt40APpqKugNgHmrT6vDxfA7VjcawmVbmu
WJkgMUMzwfl+nlbBz6QuWXNtmQGpd6CY5dijZ4BIXTBhXdJ9p5Pys4QH+qQd
hA51LNrpoe5yeZqussZbsUk7ozWQ8qguLeqwF234pfc08ByZRWO6yOBgykRM
+GRBYg+bnhpziW1tcA5kq/rI0PPbDWhUFoiJkCSidxRtC//gs5sX38FoRfLt
QyORMy18uwOtFpUGJg9MdHHKaxBIGpPaUFBQgLSk1GGZoAs2nBAF6ZBihNNE
dzK25lkBfnqbFMpH7PcHSTKkh5Ylu5ji5C2/OVkeXpD8HDrHKqX1jm4LE9vN
YdJqME/Tuog/i2FaElHCRHpXvSlsAlY1GbuH5D0QTGVlg88D8Cqc4BZzdPoE
bq/VbDP3bHhGNs6xTKEq8lgQ2Z25Ocip2sNZRvqtPfejLlD12rpe0GcL1mks
BCjLUtil8VzMQr24FvEVOaewnCv5AytP40HLQxvWfzu9/76YoNm0mHDK8NuX
FxCDT6YfoALX5VMGwmthtJ3+jzh+ESS9sU9VNeUfQoSdWM8KUkStpZKx6qcI
umE2OtNe4WRxmajR0B9/2OYGzW1p/bCLVb3CSAVMrEyuQX3QNlZce/mkR3XT
Y4rmm06JJBHXVfZFL6VPhgJO8ISpnAhwSOZCmZV1akw7FL+4jPb1kE3aaXA1
72wDVEa1TAUuYMRxblTTt72YTG0QkRF6WN/2P6RLlhyVEWAXEupgSrpcPGwg
8YgjJpveRjodf9eZLoWavNzsPFhqv/QFOEQCcGNIBLsDF7o+yN9bQJ/ktffa
1ARp/G3QIwqlXqN/GeZgT+Uor/o45RcuQvwduy018rcMlU48Z07q4pmZQ7mx
HkCFVAvoOqVj+GkvpeBAlMJlDm4UxivQVqNb4XCzIyd+RSUMrSk0IpSEzHz0
1qwH6qgAoUJ4ZatUbkN+giLJpehGwy9/qRGPUyYIWr/ykx2kPNN/TeheOfWE
S1SZogbL4LVfugFdozTYVYDijSR86HcitNY+0cANfXOOcVDGZ824BXCJ59pe
2ZuemQECYvaGQhGd7d3MM6R2dKudwOwysa8A3rxJUVRjw8bksKXnXVpJrCHE
ylZOAtGRqrmRrM6t5aLSESeaIZeWBuXeyKU0GBFXUaIlsLS2UCg6D7aAUTjV
XPQPpvDT35BsfMBeLC3i82jCMhiz9o70K//VZ7J7yOIHwX905/Pew7Cqsh3F
CqtXYQ3DeJSVbhCTSLrCRTnr5Htw66jwIcONmI4F2IFApLMUHb6QqldSb8mp
wTZgiFIrqgvV8rrm3SH8cYKlNaY3Ms93Lj14ontJYjVDlFp2XRje1b9Wa5rd
xmQ8DiOIEfsJyyUfxNj4E7lcvfdP0na0yxoTxErtTEwlAZQM74xWRvbaN/pU
g/yr23iVBRXtsPb1GP0kSD4MvrND+KH45qicjd1dN/BZZAk4Z2c35RHjV7D2
46bc+8eFEJYWqrPzSpFJmSHaA8kKMYUIIlCqDFRDqMMEInhB+SKOBHo0fSQA
g81jIHdlVMutAQ3edxozbHHAND7Ch57YazSX3dwZ6odjbPUOOflRGE/ENl/h
hSjZ7/JRX9GIXvG05WGDbkMNRR9eP+Q/U3377P5Pg27IhW5JLrvyDtJrljgu
AlKfe33h+82PBMQs6Qua7e4tAObbi6pf76pSM/gGi+lgW8B2N5GeIyPgV9GJ
2IfY6bGXWmG0KFK124NZqKP2NqZYIRjI1n998FCTFytZyOYBTKd8IuxWnnI/
sN8QgPHtu+DfENnXdbjCroZnfq5WoUzJhYT4k56yBTootlBXrTIjsT5anVt7
QouaPgZiDfygI2VnamgKWqK7twbc+WfHnQwa+1T+ahIcXlMu+6T0HGxXE5K9
ql5Xw/u7ZtsnHglce57pcI4W6hO0coZLw7Z4zNlBmwG4WjiQqEHHQG/yEy53
ZWaVcpmQpFnGc0ZI2AtQdY4+6OuCmkuqchu9tGrP7C4Qf/4nR0sjF+DpQaSj
2bNYZQvc1LsOnDZidc434Pr9rPNUjWxpkx5ikgwz2rlcPmavRxoZGNturzPB
xKiWC/dGNW9PPkiD17wY/N6+PTv6gvkkEGRF2MZwWIdboAEvoOFUwnKDkRsd
SvRaaxV2ZFexLUtnPThUbqZsl8TfgJoTDYWtIMs4MsS9LhXEFvuGNQEZMe/c
RW5ftuUkE6sMsdlu5lHrO598VatXjVv1SrW6vAV8gv4U88RHg25Ae3MW1BLp
EDp4V7v075pWms1G+uni9Y/g2xH5/FUUeYX87mtfXewUgK5R7SxYPNaZHiSP
3qY6ufpjp/QMoG/UUSCQu9IWZBO9n846Z78qgGayF5HBUYSFyQNmkwQqCkg8
dyuoh6xfbxBkIWq/lL4i6hKVQv2f3WXVH3dJLjNIrwqzmXTzRMzScnxScL+f
wyIcZrxMOfO+VNBBdjSxszp355rLtify6r8tmz6aE+7LhojUa568VvLTOqrO
GWZYC3viddAy/PD/TWVbDZYZoC9xXBklLjvdimBNOBJkDabiSgHB4voymgRz
uwy8YgQ4/hJaw4Waw5pbBcwIyUYUXx9Dy/9LN0/ddxOfAwaobyXsEbnXi0iY
y/BaDf6R4m4HSbs4uKh1vopMhXqXT/MP1H52hquG+VfWVkRrw4JkRHPjJ5i9
D2OQOnwHv0+5Bgt7mSXhHJlde+FW7gSt7VU29pEeiGsxY8YviiNCcsJYZ+bj
Wpw3+YWNp0r/iZ2YkAOEIBbrT7bTwB+exnPtqVHs/jLZhkVwjCUzZfX5/3i7
T2TH8UKF+VYioPPNFgATUAsRjzw0BTM049hG4vc7aG3snClmNyez1YGYbCw2
1Oc/E1CEhNPJ12rSE2bHEhjCJ91NAVJRE4o/RP9oS7IQYtI4u50gDgg26IQ3
QL/ChvDbT1wKU2pKMneLLXmiiG3NG3hOze37i/unOJIb1q5NcCxv0zsFXl5f
KXMX4jMcvcf51Kjtpzhs20UH+mgY20/z9uGoX6SACTxxbNdVHC7Uu3fQtcKS
scLUw8hGWPD5ltxGh163O4DaO4MqLtv0R66+dupG5ent/Be+ryVE39beebt+
fBcd0dguMAhQn1k9SxDBaZD31Ey441wQwrbqBuT/hAlQFyMTEJwZsm6PagvI
WOzk2imq3umxPFtIeHXDknL9Jtb/vnj8qUWpprwZPLxS2gRxVKzHSy7KFK1V
1Ucq76GIMPHZCk+kHpCRd3ACZCC5QRCqYC7ETdTM3WMnolccCt8CY30ShUVi
+I74auhuU+z+J3+aVX5Vv+eWDbf3XEUMtxPtajspowC9Z5iWSJpHg+HmuZEw
oxTcCBGKZ01YsYPfO623RpR3vsyR1rBMOE10GUIBj6lLhjSb1tnK8ldOPuI/
t6+xKzCiSM5Z9D7JzIn20G4K/JOfJoM+L71f7HasJbAa/usLF6skZygJcPaM
XbAruvT3VLo9I3GsKw0AmuLJZbqzaGw73+diWnydFNzZPPpra/3QnNUbGBc3
R8xohuWKm++Zb+CVnyXshjVINOAkS4ZnMhvXjOAr7IIjkTdQ9Fc2uV5I+XHV
EJojBrM673FfF22qMP4wzHJ9+baW+ZoyGjT489e4xD1xOpeKTG+safurlkyY
k4kaujpO+NMZPrkZ5njobg+EG1KPfR6kJQSoVNk/VTkt1KKpYvVl/ozS57ym
i9s32B/Fn8pazA03UiKKZmxkst635qCpeG6/8NgihRvhvAJYbGp3NCz31d2T
OvWPbTvwY1pksh7Uv9B8GPX2PdnGuzb7+lr9uCb4mcUj6H/k4VuHFTGVwchF
n+SBQXdQAivYr5T7w3tewW6e/eQc9sknRpGrbx+Zcm/QsJZgITEJa47CiJXt
HfDIl5rc+yntg8usCCZss/A0Mzr2OiUByj/l9d6sti2qcsJAQRFU+fXZLdJ7
XnnGn7Q4/+zIVee9gwrAov2IemdhRT2alx+9rx8uZJSdZ+7Ac1fSpMfxA8dH
FW61mcQRzZP6SOk1o/AQ15/uwYisNuoiWwp5BHuzJYhGvZanTeG0bCagq4rT
xq6D8fFsKhwWBwG7hf3Rr2VvBHvKId6N7vEloKfc53Dfs40zTnzbFa7tx+1g
d81/qkCkMWM5uzBmhBAb9YuXDjaz3QWBw/c/dqNbS9dgqvYF6Rx1ipCLGIbG
P+RAOeesttcDkplXcCSvct6Eh/5GgxrRSPXnSweerSn+bJzXZuklI0rJBBjF
mE637RP77RsRu40jPdTYH+p9Z8ShdbnVxTkbZ5g9pGddkZNUT5a54PNI/FBJ
WseVcCUHgz1MyAfiKa4qx+rgJUthSNMsTNWe/wW5mxxfbhsA8fbwTUVnHxfG
NGi2wvdnnUcbG9H5uiILAhRZo7BM6jJCMl8mOJ6ftwkMTQSiQ+ASJTyf8Sy1
mqmKzPGwk25/mI+nicmeGLKKr/ZHFwPpajUrtzAQZ8WQZCs+z4WlR3sZqx7U
Cogw6kNxBqyoQatYfe8NgnWb/SRN8BtewmQeiACuA5k6ERhxZjmtNRuZ3fcQ
2KNZHmC/3rOn7AODlJOf823bz4a4VJdNeD7UiF/0fNj01rb0+al5bu67WfQN
sJDOYqQ4XX3b9nRWw//3pcQ0kEukgk+Wrn9be3+lVDM+90jF0KxRvF7vKQiM
xze3uc83fZ9UU/j9g9fNUSSLxbcb0DBmofdCWhW+TNeIkbYob2cyzCg0sWVO
eFfRN2ee8FbYoeSrvy2Kpu4vzHcVzHtyNHcl2/4aCdyLuDuGDtcKdtlnaoKT
gEIB/y/Lu6DqsML34tSJKJ+kIpZptVImOdONdBDsZxV/d2jqgmSM8m0YA86w
mFEIr9bCF1c780gtyCUyGJgYX929u5tVtQgLTGyMnwLG63PNFwxxsL0XOQLn
mTBklolVUxmMl8COwRs0AFl3kUycfdx5aDFXZtPgr+R35vLdesO53NDuBBaD
MZvFkGQ7Xfnv4wuvZoWTMJNwUoXvyhszuZh/4yNyiL5n3K9TkQ7Kk5unhDsa
6Wotsf1Eq/L74ZBiwYp4g9dALXaF4sw0ZcaPHrjo8e+LXEnoN0AWhVhpOqgi
U6ND4Nls/kwDV1T7RhICxEU8Ql7q7qksv5uWh1B43UHnt/X/Pr3WIUmQF20c
G4wXepaXVlUc2aiGjxegpFrn63Oq7C5Ma3FLeAjj0O6bigj7Q6JiwET0Cxc5
hgjj2sE5pDKMewRRgt/xpNXWjRO2L0I1o8gXX+qcVq50yTYd6tbZST76Vaii
0bzBwV3LzqEfAJ+xwP4hrgo8ERz45o4LtsadL8BKwB3hWwv1yVyYA15aXfSc
r9J0CY1Div7Ll8DBqe8j7Bu7rwcPNGt2/QLgMiOjgsW4aMgqAr48dQMlJDzy
Ut3q4UunxZ15RwDVKSkGkIep+MsibNtqOZaro2WELFqiA/EhAXgM+/8GmXAG
F9Es2xuDaKoUrCVFd/CSCuDbKY4X9ekh4lxGAiRdeNLfyB9Uy71TRmI2AZqn
q4E3/NoOIvLLZHcGMEkWKqj/qY12n78sNtkHlSHkc7NW4WRl+QHSPCUpaN0m
GN8d/R1Ig8+KA44Q3GVhJds6q83xt3+nRnZKoQuMY0uX8fRk1tZluGiDyROH
6SlnWrVYiSJ8T3FN+W5C3A7ctR6gLpt/5hYXnxacgCq7udFkRetKNx6U4/Tc
ufC5bxWjTiFpTNlhtFlaIeGwJNS44WcqRXfq6ZOman6apUa7pMCY8Q/OhyHD
ZojgEI4/PlTkBBHtKOeXaPG74e+nBFwXhqBiXxMesochzjICAuZBx1llluad
302YUwyx+bcQseAB649sbXCWo0gXJ8iNa4wwfJVzElDxAhUpLJ/d56sPMKj7
DF/9gxd5TGBQZplao2UE4ji6NnsXbhmGO1FWsmSd3DEwL2EcMVbNBXfWXOY0
uYR0SDWw8Y9DdfymaMoi7Btky9ljl1NH5/Pj7b3ccl+8/0QgQMAjFmgcGl19
Sz89sSH5xn9AA89+jBey7LF+NsjjFAnPS3JK9rR91gT038uGv5NlJGY/63I9
aqqZJx88KVi9+T7NOA9XWGIBK5Y9xvi8cBXOIoP6+tJjvuMerAuR7Ex+QawG
ijrOyDtTSQ52HKiHm8WbVJir5LKR2u9svRegGYawzKEgx7N+NowkeAAX+6YD
sRZIwnpp1ohz5gOLqe5+i3LDkR8O9f5Gtbqpf0onE/vLMFTHia3lvqHLz5qz
S5OkjpK1aFWD6SW/fbewZ+9ZalLSC7BKyaw3OHmEgj8PXtJOVi/gdD/51Xuh
i0kh1JBxdrCxX+WzACDazwCFTTEWBPHY0zTaMSLmQdk3ER5mSl6PL04BsZjX
gcCL1/y7cKFnJPhtG3HNDJvaLMOtsAkfRMKk0YmGAOGQQVeiwYZoFJ2cmjF/
PL4t+9EB0fx1AcYJ7794AK+PQNYWlFH+qsOChfEidrWEPID4rbBuDigUXUXg
TLgB81AoTeEI8qHm9wji25Qu2TntipbrBliR5gBHif6Srl9yOKjBiGh3tubR
Ya2LBo39IM7zF5O2fGldlWRaiYnImvyE21ObPQxdESfuC/MxGayd7N/Ub4tq
yQ0dAp6IW7cq+mQFYWdJ843ZwVIHXa7gc2fjBnLfqZcLBf5R1K1LBa/9q+x8
DpPuxi3dns9rghDHqUcD+Bd3IV+orjWom8nyos2/Ye6EqK4SG/kHW/RzAcVY
u1zi2PerVpOJTk6LDAcOXoR605bwmBEhvyccTdCyBOB4sMu+vGtwA5w7jbih
1ffCkJB4rSIH6PqqEaZcRLLmpfmjGzxNnzbj8eMuQXINxp+s1yqnJP6lKdmt
3jAuUAccDq9K2nvOSo0KrKUT83/u8mKcguPej/KkG6W7/AcUGRkv4I0ZgNca
0XintXMPEWLPVm7DHLFDwi/FrwmxiZaVMvj5fqvjit1wZnsj2OkPcdKLdHpL
+BNmdL5Smknv4S7aIzzhQRYZ1sLAE91tbap2/3l08zZDOrCksyxjbW6lmG1B
cK/PPMxcZqidzFetkOWIbgIJWtM8xpC+d0F5KW16Lh497yibIJQQ7g3b3HXb
jxjKYaiGLKVHjrRI819pFOVSEKnYCtH8yPEBlnGP+zUT9GMPaYotrkYPF2ni
en3G3U8eVWDa1gE7/WB2/Zg4Vei9nckNaeM57tGfDpVIsHMVVCjbInd8XZHr
WbmyEtFvKodI5ZDlR/xhXAYx5TgM1ycosNoCZnnJBcAWKc+C+v9oswZXDx3M
3cDWUu+RX7rbOtRVem4h8Y+AyU3gHCA5eY0X+nSR+AlgZnYBjs34iKtEN9jx
i4qy8g7HVEJtV5RajmdoGaZEBV0EjgCHiOpG3rWqWnuoN6VVUAa8CJTzdvyV
TaYsLb7h/nszEdhTtsBhVhEQ15u4I2rNct2rcP/zJJ6PiQTmiP/b95Rj2DN5
xZjd11D71i37Gr4Xt9BDviQ4ikhH0vRaw48NyplD/ODaUP2MTEjkV4vwa82k
fYJCT6U1bIc5+x7xT1gRwzI0vMviVZi0ewF9ktPaW9rboY/BLH7q8pRP283T
cu/T/b99JIISOgL5pffl1TZFHPSaAQMDDpyNsrwwoUAS+5PrOmEnhH2i8/bL
Hw058cxWUemhatQZNVtNM/Qky0UoT6Eaqa7eNnl8CDcyw4agOeD5MVYQ13Dc
+izUmPHTYxvvgUczAQcz8Vwq6PyBIb9AR41SRIJzi3kPI5sRY9R8yHljPBAY
PvpUQXNVgk5kEwNxq89KrwClX8MDL/7juG14sTNtwkMYRpJfTGtLXfxRDf1m
2t9ne/TvIPRbj31Hf0kLXsSAPjb49Tban9dEap5p8gd1vOAg1ALDn0mEIibH
IRcOb4ynHO432PPM6V9L6uDren8N+JflgIVLWFyUdQoxNdVJumTCpL21FDac
PXmPNYQmVOGkV4gI2BdMl5/ZjDusQUt+Slyz1MTP4MYo/WekcZbYFt6VGu/j
QaAm0NTri5joLOqIPw7jrm5hYMBhaG43xE73aeeZoQdc7M9CYO3sse0SMUWs
Gb6WJMB1eLs6YxSaFg3GSGEPxDFZn7w1yIVtLIEyADcw7BSn4QjB0BhAYoY9
FA0aIa44x9uYw+IK5D5tXSaSkruB5yn2lZrLHouTZ2hECdU0Gqf4/r3vDAnq
tNuu8M3aI77S1YUrt/jXkWFDwCLJ7JQOjWWlbKQ16V4KqsX5PXJ38/bWJMHN
WqSS6ymzByJ/RipT8bmEJ++Q+tePkvS5FenuyFRp6vXpoxjSNtNoJdFoMaR/
nmp9KdI/jFK3eUQmti1xPlxkU7cYeEyIuzU+1pzqb51byas8UAilnFrLeseP
61A1wrlSTFhSQ39pkidhsFSv6kJ29OQsxWFXaCauZSvhW514oQpBQrQW6JUr
rH9Xu8JjjLHc/wWXEjRqpzALyKj4ibyg39pG5LGYxJJUeRWKWBwqqN0BK6ji
pG3t5qv6Or6oeGZk1SCPwcHNRH3c/zezTMb2WYztIymMEG7ZcQXf7TCPxVMU
THDF1p/uM5OMm3nA1ZnCHveDNZiCSX3UF7Gbjctne0mdzs99B+HqPWUhRi3H
83zsItoFlI6+pne30dvDM7sDio1mmoHSL7vuo4pKpezOHZs0dzYMrGOUD02G
bXxdYydORwjWuBIWIj5LoJzInHVI3Jr7+Z44dt4hS6oNd3y/BLUqw7dlWt9J
l9xbSE64D0hdmPTkRlbJFAskjgn/7XPVH50ZmwmpWzxEXsinXLK1mFk8dKA7
k7gJAAb6y4GeH9tFG+l70dHc9iqV13nTkhCjJegp/3lCxlhMrMZYs4XoMq/K
05B8vUpSk9WHb1PUbHBqCk7kfddzJnefd0oawD/e4E3K9NFj00o2rp9IOokA
brK1F4zV6rv+ZpZ07qtcGHJ+jkfqUzNomaKdGCqOr/0d9JDPeGA2ee5uK7KE
dVDYNdLcBo5cCs+uBbQLHrYOiFXbq8tlN5bJkN2IJUmeNRmrLzwm+94I2ofu
R/9qawr/AMNaHT/0IVIZU897rssh9GWqLbXXM+3drYxugga9j1CZLv+TNLA+
92rVXrBE9tnU4qw0oWXYva7Ffpfh7dqNuSr/2V06F9r13uKSrgyc6amnRJ5D
dbGvwK/5/6yitOI0LRmBZMYDXS0aSKZG/EVulPdWICmZ5qHiYz9U5heTMmJB
y5VO3eQu2uPYpAECO4vLejppmzclLsXv3KlUqO+vjONl1F+/TkFOQyWSL6Sd
KVEp0qVy6YWrnvIfYEti50XLmloYuAAedzHy0ndIneGrNMM3TGlMOdrgIXUU
ccmXESEkuO3Gp/TRO5Ku6np2djR/MGHY5mqJA8hYOmL21bpwx5rtHmN/yh6x
sO+YnFUHfiRXZWxA1AK43gg+Afv/5LDtSIhdQbpAvLcvyQLX/1F6vpvaHzD9
1/rNZMwbmF/HehExjrR71jDpXoOibS/cpctere21WmEOir1u+lgrk3fNSmnu
bUeyEX67j5IR33AXBo/ahWZoiPWB1Y7c4z+VMhP2w2N+zSNAWLLcgpwXiV28
LhtNFGLQ2g+38z+QeC0A7/TmrIWwPbHJYmVKac8ZPYiteWuFxzxYYKN0a8Id
7sIjchjNee0SraYFWcoC+VkDavRFaRSGfgsxS9A+xLMw2bpbUGuOz9yUDpIo
mDemrBSA8OtOSSIDUTNfnxCTqnmqYqSBzYo5yQ+vT7PYno9zp0Su0Q2kQ8KI
rPY28OCXqcH7tp2Vvn2czVB9bf4jL4ZG/0c/6JBlRVt5CUbPZXDoC0nDfGd1
Odauz7qOePkZmoogkH7rsB7kWrbRXvEROvAhRMwbZHV4pgk3e+yVzgXyZQlq
3hD0IPNejrjTzRFUln0jnyJyA3RiClyUT9aqvDzv/fwUHA1ZLsRev0QbcG5G
CSM9CcRLch/SRN4wpOV+ofZV46wUagZVGJw7vQggq4YVgPG0GDCP8m7XHNsA
UnTmSiWDvtDhAO8WzLnPZ3qy536k5cPTd0gb/7C3iTAb71N1m74VDfO3lZf6
+Abnknod74Kyizjc6pyn/9sKqkKl0RVF+M3Hv2+E+ejUX+nsI5M8eoNuPMhZ
fgECvmko3HjW7VKw3ig/Pd156zGKTvxX+BlU8Uw3Jd4i8hyrT4EVtnZmrMsQ
S+ChMYKfiltzZNQ/TOK/K8JuVMIgiZBWVRSEHL/KZcZsvOQ/rYyaUAgC6e1q
C1WzCTzKj1OVnAFjc86ypWQ6zNMaDxQqEUHq//9rgvmFKgQpwvuvYEVU52E6
ie6VbQuWTqdVgIIcZunwjbh7l34HPM1JMVJralrhvktey0pW0IhasvsAQoCC
hverUEz3Dtso25YikO8yW9FhrxoT81pH5SdSowY2QUKKJus+7QwofqwGyJ8f
/KocF063AN5/sbTe0w15uIBMx2V58Ndv5uYEgG1oOa8QMbXMV56LOIY1aqiA
RjnlZ4lDG2j4qy9phy1HfKcMQ5Ol7eUwOGfhc5usnc3Ks5fgjCVw12iLPkx3
g6or3ryHDwo3a9fwhOW0VSJ5Bjy7bFSJyDMtEoRH2IpUtUDfgVEqmsH4a8N7
5Nsq5MYJjWzWTMsmIdgs1RlTZrtWUZtOHmrpIdRM3QEMnFqdYipIyt6G9Pz+
4ki9FzMZxLo3cjkDghK6avq9M+m7cSy1RpeSiwT6X7XZTxyJraEBlj+8YDGX
7ZmiRR8EYY97hWYYfxE8WHwdgE+LWedwxN/hCia9HpqChIDo1Oyx0UxzuWyt
rIUfwd3bNDHAJH+hvQ/WF0c9aAQIQFPPWjbAlZghvFIU1GOj8bS+UZYHBvR/
USIxjLBgvuhY42UCW8GOORdbBI87ezkFFtXXiYXeQvIgSF/LBXCYk8fYVIwH
OePF7k/HXd4VnsgmaZxiH8fhHW0ljcBjwwe58gk+huZ/Lz6P5iotliF5+WVI
MgNGv7m1qefRarVmUji/NB8qtyxJUakl83NVpIcwkRQuYd06X9pQS2Nsg9+F
wfdMrjhDTzvuCyLe7BlbGS1lCdwSnW6l+4rp8dAIfxXlpPxTCjjvGndraxRj
bESRh+qwSbYwMLhiXXKJJ3/342rb++eUHVqhWYU8m7ecvoUCJIloQ6R7TPQR
2PJ/RmXTTDrl6Cz5QOdpmI8s6vCmKcIx5hGOh5efDxwm7+hyTuZiv8lDusVw
DyUxyz7V+wUSUseWh58o/i6UCGaXm8uNQqeevgAdgMuX9ujiTrnbjZRw7r15
kXzVTOiz+FBFkvPSHek/+Uuae6uELYKWEWrmNl0cSlxt5cJ7V7WyX/hBwwKN
9pY9TMVbpyj09HcOBNRvsw4cduFubmKN+H2AOLpIwtssWtGAXJVr/pcnAebb
IvyzzLzUNb7WCTaqdTrwLQgp5DRqkhkephahTipedEdlWyNOouwfp4q91iCE
kmmGeWDS+VGVfZ+y1vIJWfC49ahODkKdin0nZPTFVKlYcnPXvae8oo+UZKWO
f0McaPA+pLBkyRlXnln0n7wa2l/LnfHsAuXX2hIUIHBBUkC4sc+NomvAOC0N
8SyUGo1KlmmjiUlVsSH4/5sizawh3GSKwPfn+k4DqNxVontJQLhvq3IuHIg3
RUkI8q6cJkR+elUn7RUd+OKJxGATtw230IJmr9WpO1LKpDEHXI0prq7aM46y
coKAm5VdmVUpoiEYGdRQAKdWrUX8Echgonl8NQvWp1hx4fKq7xcDDbmfI/oI
5MkdnTu5tZinP0s84A/aTgvRvK7gGiMW5KLdr/9D2wu4Ret/Q7rY/NU10aEO
MHWWz0Ty3DFwrnHmicn0zzf40PN3WKQU5URnN5Q4Twgmou975vl3pp3O8+CZ
s4f/GodXV1NbY2Tf2hCRyiz10zYX2UnC7Rwo9aAqmvBGzAaZcBNy7EbrIE9D
r8gYXr9ivQRX1S+PBh0UOA+vIFr8X9yx25rc8clr4GIvVmyvaQutRrAXg79p
v/ybNjMpORk6rwpREYzzg+AJKkH0MAE8qCT6jW+xK5V3MmCgETdvRxNljVTM
6qUyveOhFZnByrhy0FnaIOV9rX0EQxVH0emEhMTihJv3UIX8bWFUlk5oiqiW
QJ37enibvvU1Ld0ChNxDtvl4DPNsaEbxjd8IL5Hs0Ifcvletzlk8blWsSvPw
cvPViwfCRvgIcvDBch8j0aYLAh40pSmLxtGTh4hhdETiWhEvlJBAwOe8u5BJ
LXT7goQbFuU1WlTnJuJQR4ehMKe20Dp5aOekWqWRfc18At1KTCyYdTAl96vR
t9YdNtQjO2NYPzeGZclhvB4s4ca37w8VQ8L6B/0Im6ZbgI5e8bPvDxRfd+jd
y2DRZ7ST/PBZIDMYTANNLzhcuoV1Fcqm/MFXdwjTKaTeWfijykGwZ1S8HDPy
1Gi/lQ4jhYeJqgzNfvDIxeWzGgTjIg9SEUkQjh0izFmLau0A+0veAXCQGd8f
Yy7lL3EuAcmfkIxeQm+B05WoU0YX+Xcb/5UxEWIlV8nXuvR8joSVvgba0gHK
uwFrFYUytqkBbSGNfpTzsLM4yjXPF7vcgPDHnlkwkF0GWK0u+UxYcYRe6K7B
JuW9fCs3xcaR6A9o5+Fynqm8L/fxBUUin1MFL2YIF89BRtnW0mVyJ5TYTJyZ
NmmIgKHgFEqlVKyTQqpwVGcn7PaUKSmwo922nQoM26AIXCmS9rgHDxRoheap
Gx1apwMiLV+bYtbGihLo4EoQt6VmLLsnmlQdLLp1Zcz2QJVKidx4DqFni3PP
3ZsWEU3YlQ+DUdvzqQBsXoMgPsVF/yIDQ+ksDdqUHxmhxzz/U927To6lohvp
m8TPm1jYP2d3aD7kL/ApIHpWL2EhxKPJP7O3pyA6hQE1mOSIioFgx8uPRsB6
a2kH6s1BVW2vsGOXauXGMHyqdcRw5zgEdAL5Sbg6+A4YZ76HSXgEqk6+0YEj
q0/aiGgELvT0MCb3zyvDTDjchoBqfwF1o8cz4XE7HI/QkmbapZv2O+HeANWr
+mzheLHU/O4v0w/L+H/x3V5Zw23trRcGCdhSebroX3fjn3S4HbTa0dwzu51r
T3hxGUFTQfwlFXZrV/z5HeJMwt4J8osBGQkLBK9HtknS6n6P9+GcJSKAxtBx
ba4JCv5vHRxmXdG8+iHPcuz5Tmq62cX45onoffZq+4bJPAH1cjMx7uT7EB0M
eQ/iTBwUHw2MDNCWog610sfbaqxA9gylWXh31oGp4qeqYaLsgq6aCl17mub1
bW0VIXBcBRIAeD7HPhm3Pqd6eYSCglpp7nO2FqGgUVOhAjFjrL1ZK+XURjlk
clMET7JLsRd60M7JIQ0cMYHcmPXL2FjUdgeViYs3QYek3am35ackky6f96xf
O6cbckCTdzDRhd9TnsqQVJpBAewhD4ASKp9CZnZQ8nzTjJftcEVEPsKPE4ht
y/ZeUbRo7jFT8OAyr5Z8kNpuv4hfx0DkOb7k1zTZLdV5pzQ5aamwih1J9L7f
HLvkjZuMXOxaGsfrEPq30QkRw2jHqiDt2/ZShA2tLJepUb/9twf+odK1JEr9
g4q8s44NhKrSPWGeiERA3MM6ObB2nAXcxnkZ8Z+ltRTThYQPSAsHwJkashhZ
WxMH3L/gHa1irJ3MsJC9VFrcG2Zv/Ew2XnDBk6y6WeoLy3y9uN9QWR+GIUeG
G5ylXoXE6LiIfmTiNb3LCV9Np+Ayr/qV9zzlpBdUWuOsGXg4xGp8F6O0MrPR
2rdnMmLwgJkyqqbmA46PgDMO5KmWVYPvK4Xb0M46UaeISEiW87OSscNjaLo1
s6WgEWf0kMdnZoRIRpjNhhBAq/nHigViZpkWBr6byOz6nmQZkE2FVZQI+Xya
xrWxbPnEPMj2sQgcyuT0nseiAwjL2aHUNuOE76Vv3Wm9yJIyzLXrojZ2VJuY
3HA+KJQhNZcAnZtju2hrMrr9nKIBVgcxwzH33Um3KKUDLjJQ+SfKNrOVLhcB
DITOScm3bJ2F4PkYz/X2aUp2kopuPxeC/IV4aog6Wiz5aqkTL+eSYYvDkOl2
sE3AxVX1KQtUNzXrEoYJo7eu3afADWIOKH9/rWV9Gsxs1ZOFOsc8AFc0Rssu
taf6mVn6mALN87zOxHfXxLF3I/qlY0JN2oBrd2qkl3BexaAxNmpPNMdURZt1
YJTa/rN0g0Mhy06dxJiZmqEDdMjGKxaFAn5zYYZIKSp8t/erAMACzK5gECk8
MPbqImFdPzC2byC6x/1lSE+DKIOJKxG2/40ux1Gl0VI+kBUZ8RSZXrukwv5u
FQ2qSP5VnqTeYMxO5v0U2qY4aEG3GpVeiD1Us/3LZL8MhOpK2F1Rn70ByGvq
4MhWFT+joYEjRHCLu4t9ty5MXW1hGcZX+X7hyDvqSVa3rNnZEz1JSVKjjGeT
tJ2Fv6hGlQZ6Jg4I/L3YbFkTuUFfhA/cyU81euAkKidqoeosbcpokWz5QGHC
+4SLo0rSQuJbQYEDnEFUlhD7fjSXv1d0wnx6nfQY6JWCgTrwTVByGn4UfyZ0
aHEU/7xp23aUb1100mjcO35yzmjn4/J6GSH2UaetKTGEviZiM9bw1EJ/lE80
Iai1QjQLWG4X5SaCA+OwgpzOI51bah4lU1wL/5uW9W51BFkBFAaDlKAqaOQI
kw8pEtleIprv+SeAkyGxzz70PgoLSSA0yfc2oYZMmPK+Wv/UQs7pglkX7+Bk
JeKpRU1uoiffQVDQdHMQy0jIgbVExeBwic1zwjeslgu0B9e/g/0pOl3Ocm2e
wp10uWpXd/K29/N9FGwrwmmjR4baCFbksR6fLfGncTKrJvRd56uZP++nea5K
6tGRjmYjrz8A5EX4lB9UGDCQNHEPZxPyzZRl2xs4pRFeCrhQZI6kd/B0aU1O
Lu/In8N0CvJ0UqVzsVgj0NmwZAVShb3oBuqzLpxczZs1sdmdf9l2ZrXgEkzG
j/yu34q3vrVEttN5JuKIFPsKZcQJ/ktt9v5NO8aS4CHZtPUIEcKbxNao6Cjr
Q4Lma1tpsAdq01LnuzfNpr9NwdCRmAEr4aLYs6s2kk9MN36nxIFqcVNPFlgh
ZIyMo2jvBhh+w+ba/bonKb4CqZ9pbeHFjjKq6IlQuKDXGV6HRzBqWih59Eod
+h/PI0xSkssTM3DiivQ7EGKtikt+ZdP5ovhmVmqcRhwFL5LIFgqoCz2ulrpb
WdCkFuzgUKMir14TiWVdcHyUrEblH76kmGcdTlBFHKCw9ndS42TA/hvwAzec
Ble7ol1QRKqdxx0EULG8L5nHOJXKYHhXuSoeI1z3dYUkQSBx2+W9t1MOcd2W
e/zJ5CNGr+rBY5vDHvpnvm9aZwvFyAbZkBrr2X76A1IasGyskaVnTRQJqimR
RTuqFAnTJIFlqkmolZe+Xj83Zrn/9to3C1BcCbJq/a/oT6Z6UqeDx+7rPTJj
Tgm0gWKj44UbzUrweJcpLenUiD5rkVcOChGm3Xbb0Lo1SNwx+GaQq+FgNDWV
jIch2zGz4Ttv0ZxP5sf63sNEpSTBk7mGiDFvGiFC2erpA02ZuOFQJplyFGNO
zbVa6UR2Xi6+v4vg8TivzCGtvBGIQzSviz5Dod/RBlyAcE1nZCb7oOmkARqs
Kx6rZwrkTta6EHRjleUnxQK5FwwinM2OTperwOi9sPCmvG/34hRgGAfhyenE
JwNaBbqe7jZIGSEdD+FRNbbVy1lniMsql8I0J02wehLLky3isyXqoTuGtcWp
J7/oX+13nM0z5WGXnIo8hfTPUB4WTWFONYJSL+BLWkQArmirpsnfBCcp3JJ0
6abb6QI4FWc4dm2tqmazlanVt1m/KoMqgCqfw8gpEaHFh/f/qxy+yTClok17
pYxcIUk01/hZsMVVmdIW+WeMrT0R7/zwGZcJOOKc4vHVaxlkk/xENcTbohow
P40gCgKrkfLHgCxU5PVblLRf+g02xub2xrs0VyE+0PJ+Lmhup8dALhHIJ4al
hjC1FHgcXlS6JraZiwYJe3kzEPCbfm/823VeXpLPpyymAg3QCAD/tliRHvMK
HcU393PipAPoBHNEoO8GPX9F6aMMxBCb8MWbsUIN4ql9qV39UzAiWZkej9uq
aX5DhPvbp1zZHAgvHOxb7XMlxwf3lpo3SgpsmVSvbxfgHC3mdnOWB+Rw2FBA
qiViJq/ccOHwu/WhraUhltdI+b6s8cQHTHFiAeZRuh/FhxjFPXsW340bHn/s
jG+lJWr2VOk/KbyUKa+A5PopVZu5hjIF+CcRR9DfZzCpJHYfnu+N/ppTJ3vd
bfvjMZPLlF2Nt+7b0dG2bDJRkqZopxkLCqgeSx0QUqK/M1+9yXKAdqxh2Dhh
QL4N/OyPP+F9NJI7xKyDl6/8Oqj8AEIqK79AztYnGM+V/mE1VVCfiTChsTjB
lLY+YwKVfZ9aCNf2DAVkZAn43scce9IauJ5LiUomJVescsvKvhlRzvQc/U20
mUr61ZjeELAlI8O/V7OcLOmZm1aXurYmLllVucw6RZyLAvL4aargdDb5Qax0
ArB8sWDV4x/zq+qVPmMG5HTo4/OIiCRyit7h5b1pT3GXHMME+fH2sv72mYXy
4fh3nPOoQn6iZt8UUxq4MNOtRze9mGJTV/kVTaw1+1su42p/3T7cvQJMAtMG
J2xkxGRYhLRwxyl7+x6EIusQjQcG9UtcVY9dFirJS5JIoOMRlmoEh0O1tlxW
gQFSJN/+94hnU+78IFZNYCNbozdehncP6IB/i827gAtL8k0vCHqi3p/TeKwl
QktHFKqL8Rb1/fsnhUSF6eHHo40vTqk3XpN8W5XMdLioh7fGkUcFAF08oelj
9kuiHlMFAY7UYM83cTEl9Fu5x6qkHSY829WE1CsF25zarSEoBk+j53tYRxn3
tV4SgeDuDgYB/Bb5qBlkC2VIjwMIJdiNEuPpSqx09VaIcRtXdwz4nNW5B2zJ
4HeNDldd8lr47Ex6uwut+P7ntnwBFoME+P0ggLCpeUBIIeZTRYQeFmnHpP+P
Js5LKScO0uXVhTWL9+h7G6su+aFG3ln/f9XC4h9/OLeT44w9LSHYz2oLiy/d
vojY8UdnKtqC+vXakkUPhqma175R7N3SOhlhmPqnhmLlOvh4lUwL/UCpRmse
nW1RgF7A3egEMnO132yfip8bLi8JeUxRu+d1kcIrnjJ/0tqC+PcKjjtrLN4l
+YXFMIvkX0TS90mlvaHEvCwNeo+17kHTdIMUE44atvfrtPSMwEt1ijBJenLN
L4uf5by1dhF5HLxbR38v9JzbsjvYDzRxY9MAQbrVX49N5TNHWimGA2EW7iuu
cvjT0cCnPgxHptePD62ug4oo+2EoIbviYbo7v4sllFZzVS7WoOq5Ec7oYr3l
jq+LYMxtfmDXP3Am6d1O+8OqifH7KcKAH8wL9zujpUYgoBNi0GgFkKAnHvac
gqktU/TS1YGYceq2sjKWr6X6uW9DKcAQU6HgOzE85Js2VL5q2gNztAcKER0L
eIiwZl+gA4yAMZ8W6+sQJRZMsdRNX54csKMpvRcnso06csSXoKQ5Pu4hnFYc
gFLTXWknjh63VL9ZlkLRW6t+BJm7+3gNhatIpQhT7SA1azMmcET0EtfeMvZm
phWyO1VavsQb7wqLUxz5toaKC3XLMLzY+MKcoVOjRYXpGHOPiUKZ/1ndRLoR
D9GeJOq8H6HbsfA1LL8HCzvV6+tqCliQufYJUCvHxVQsPmkyGpDbWj+oLsIv
AWexc0xadB1+XkZ+pwrx1rOth/bCxtNxlyiVpRhd2RnJDP3BPWf4dV2XIG2x
sMSMhZ+CQF0vX/6DVMhIC99X7ULVJL9hFXz7UCddplwFcfGs3B338dymdhHs
v7gren4TOHi+XkD9dQijSZL6b1GIUMlAJCp/jhinmz4UX17lQsEY6dGAEZih
kilo8P6S/UoYVV2JVjcJxpOseqDwDi6Wz+8HD/4irKeysdQwJbHt/d2CRmOq
qhzNLEqrLzclHh1d/c+PiXP5CYcAK0qYyjWf+7gZnyyL1zJGci0hdS/HlKw+
38RVOAbSgJZXLQWC2YVIA7MiQLfmJWHdCDI+FWFvAUOFm6RS0FHom/BnAAt2
37NKnNvSCCBz1i88pgJd+BVXcDPgkazjkiPBD65WIONN7EreuI0LEI30YzBA
hipraN+/ymQMBP/wP1akI7jYLjL9a8hc2BUeuPAL7fZAXsPhRTbvjS+x6BMm
8wAzFSNMc+6LryS88UpQAc2CCd4j9w6kAPR3ygJmohpjMBy0MJdhDizhb4qr
hJL3bxVE96/Fj15a/0imowydK+iaIwm3UqXJ3ljYKWtqQgaZdXH+a/SWF9BI
Rk3MHp3p9HxaVWrGS1Znhff0jnFj69vZV7AwFeyCTc1OLxGDoBfchTyzIRqL
ez9Zx2/6on7s7A1wYTzPWa7RpxpyY4gFVDyrV8v86UicBTxLsqjCE/CTL/sZ
D59uShEabpgO50YmJOBbj4b7lFe0r74/hyJr5eO76uvDRG/Hhbda+PjLTeYz
/GLi6gXTvSt9Mlv7Tho2YE5XxBj9SPWNTlkPbqu3MVcRLpLH3eiO3GO9izw6
fhUrEf/46qwQd4CiShZ5NvaLnObHlfggW6RrYel83X3NtaFJ99n5avuiIkBk
yyNdBirR9wM9aQAM4fb02dgU1OdMxAAxcwIXc+ZAYaPjx1TD8fvGItoqAOSI
Cmlr2oh5kY/wFOBhe6YsYAvtQTO/QIN6/UkxNaXJJ+5Bn7Gq36qptSMMmPWQ
CrnN01uJgXTsfh30g+mE4o7WufraVElUKGxJSiFxp976aaA3qx4GGIQGxMBQ
u4dBBocJwwUo3fJ+/wljs2K8tR9CacG75GTSGAHC+LZgqw910ZVknQefqlTk
MHh3m6aYr3hhIH/Sw9s87HAbZh4bqu2ntFvCzCxkUV+zEfaouRc05fPMarSf
VFtgoPebwyD08+KWXrlgos+0DO2dKQwVhdwNBUx6uoC+O1/TlBllU1TZrNMr
ADEbXLjViqsqBCDLWyIvf4i/uqA7o2ZEHHrfQ964uQ251hCsamF2o3nZlsut
2CSiliqNOaqSoXRJ9cFBeC5FPm62P+U1XCYwR2drXabnv6AfFLcoCr1aYDcS
oEOHmXYMwh/l6msIDPKJzdFlru3o7Mbz089z8FOcu2QrvTw3j2V7Gw0uGdFe
q0+ffcHZgCVlO+Pb0yUjMF7/1i8F5z8DnvsSvP7HZGC9vNijDKJ3NAOQEvDA
tzk04OHNTou6Pahtakwana5u8mF1UCzcWQwhpuKrijNAVSXeMg6lp66WWSy/
otFxg6f7BQtuZ5p98d0wUQgHI2+uR3i04FdIwZBGJwYFL7zpci16Y5qPFfu5
2re8OKA889CrP+/oUbleietMgRn/FeHJHV4DI+GbwCnOK76cykPA8a66OjuV
CqiF61RgSiqSx/pJCizOIwTK4WJV4XJNgoYNHL7MLbBglsvXEFmZ/3zD1IFY
WDK99CdDlO4iHURD+kRgbVEs/9/zDCfjWOPT49uqhYcWDPNpcIOifJqz2YaX
4pE9eoeXjgE1EwQ35jyyuoaaWRtTNVveVe48UhYFY1h8LVlNfwMDnTh1S7+r
AEZJzo2MMhMWEKyTEmunipFYWRkr6BWAu7PGgnXKq/8s9h/SlwjLk5oze7G8
tl3iQ46dywBFHSz8JWPnVsRpQcdaKDfgYRiT8i/OZcjna2yzGHy6nGXZsfpK
beAxKhcKkbSMtTJe/MuSJL18tdQXBc4kPBZYP0Itx4EFTdxAjK3anw51FgGa
nY+LmwPObJeRHsLpvF0D1499TybLX1tKfpAwBrxZ8Vh36ezPkeYHKlNtIYGt
6Ml2oq+41kIud/Of5v/Nl0Cp2HLKz0PQA+odttLzHT40ou/SEuFh8XUShOaO
96BS9rX7SJP4M6ZM7A2rXIQlUUpSmLuPaP2U+1SnPZe9oC9ZVJPGgv6JHPQQ
xrbZG4h1K9DVWaSYmeBWF8Hys1ABkhUJsQfrxFfK717zePKAoKqywDjpED2U
Bi/wWJotSiuh8UvQruNF+2QdYeImSBpYdXh756tANX8eM3XhJAOkAWcVDQ1y
ZqIIunO3GbguN7GvG603dHzfEpP8JVAQrZnQfacXo3P8YmocmBV4UB2InSbw
N7qtz8YL8YXmnaGFZV+3XyFMcysGwDY4z6gBYrEqjkw6HQHBes8Y00ZUztJV
lGxN+oHO0JYQ3ANptj/6LdSEVNODvczfXOgp8tSc1tALctmw1mmC9gF+l3pc
iSTjI29a5fzcar1KYFJ+voSH8OjEWnNZFZCxCOFmA2pknZnj8rAYlmNnyowk
2vN40wzQ0ZiLmnrHyxUiobxlWm7HtXw7OyZd7JW2qyT1IZGhl9yWjHs/jq0/
vNuyBZ0PF5h5zuzdsloph5Y5yxEMvcceiRwS2WinxYVa3IJzN0/ZNxVLAADi
E+/CkJyMsoMweAPygM5rTb1DMXNTb2jz9R3UMz6iDyRbgOhX/fF737CZcOoC
33jmxGV650Gmevd6NcQvvTBVHKPnbawsubE4KTbtPSiwyN+kfOO8x6W80F+n
RCzS/Y3qSeHxiA1nAojjTl/nbRUYlvMgTSBZDoicezNofn8m19JlZdobPihV
B5+UDrmnQ4NvmpeEPpiL4nYvSOgEQSXsen3ZAz2deYeL+xS9M13h/O7zAUNu
Id9VXTtlaWaOiy6I5fYGsH8tgxUWBw2LVW4dqmRNtj8YOWdRMpTL351BuYNG
KdR51/UyWZyJvUGPxw4yl9ODfWzvVPWmhBREY+idNp5uBzssXSL4Jf9ieXNN
p1q5iWWN2ewGGYXlyTpmzsf3QJoGiKXT+l0dS+if8Xpf29OdMB3BPZtdsb9g
bZcbN2Qpkv5Tul1K+nMi3Dr+ppsiqyf6HxzyCP9WjGrHsylumXdeXJzu0i6e
AVKdpEf6D2WtltrUAMpKOBWzxH7FNxm+pSfyXGs7ewfM71Pn61ZkiF2WqX5w
IKhVI1lsqg9mNFNMqtw9dpfJnaEuytonTJKeSZwUrX5gjpCKh8DfpeAZUCgZ
3OY7QaobhlPLkDDpaPY1m+uxQlmkdI/Gp8HM/ZAfwUCd/9qdzqIOHhoxd0kO
Md4hqTmCC9tfMZKlkihXhcSCW/jEqxmwiln0FK7M86SnF6MeSDZy5wCN5HbN
7FEG1ywE1K3qCfcBHAYvlHbPkKN52E24r99siZegGbe0ldJadDwdKafUjTw1
6UyOTsRsGRfbvRPqHIff4rcN+crV3bcex4k8VUCaFz8Futw9T1bp7Gh8hrz3
nvnxtZ3BxR/4SGtW2/FIi669TzIVlqwU1ams558lA/TbbHZDseDSI733YvVg
c+kBHqZi3g5SXui8Q5LAOhwv9AOgZq8TwqhDPBp6QU2fVOB3+a9pP5g9kZ7g
aaYew7c0tpqOx6YQCGxO5Y/IHiOkxnFrVi3B+081o0Fk0j6f0PDpio3xYWrB
jaXpgYeUv/v7xbEFDK6gA8DGmNI6xgjlQ1kwyJVkFME/XNRCQqA3gMxn9RJA
W/CQoeoXZoPPHsVtr6rcYCt8/u6H/lmrPqVAAHepDrEcLIrakNoG6Yn5b5/Z
g8lliGfW9LVQb9+Kipx/upRNw3decQguYLMi1bXHQqOfmtG3wCwrT3VFDwI1
Vdxautxvr9tPKN0TK2P+/l66Fj9NeYz+pGRFs2j0j9gARKr5wifWEfCFndIK
vVG/pFA6SF1ZhFkM6wFi1cle7LTTZ41X/F8I92GzqCaRPnmfWyJOisNzvf5n
KTyFgNfk0Sl2t4IwVK0w5RG0ZNbKJVSFy6Wn0EpEeCc8CWlNdKgsvNdEkFHD
qK7iKGPHJXW0jtgv/8Ux6Wqpa+BvbIdYj8EIj/3tuuZh5/vanf3TUrJTqSeH
vpzD1RsflXjJZojvRrm/ANdXMi20mw19rNWVCs6pTB1sk+HCb8SmE+ueZCld
g8NWYcfPcGcaSzNE0feQco2XGYisMU1MBw6mklPfbIC/mVRt228ZA6Pd/Qkx
bebLWOWNVOqsLC2hltVz54ZDMQVQe0LUziA6NL4Vp72gCT45rrsQ0N19YC6a
tnboENSVCIZgPMRBTKr5OqH+bP1b7z54Hb9GlQoTQHuQmBzQyjQOX/BmeIlX
yL/u0Lrml5eQj/5VJxzzr9MbkyVTaWnLSFfLTDQ9RUjnUeyUGj8OQBec9q26
ffIjBj95Ltz+fOy0JsnA/NfqTbCh6E4nn9Lw7q2r4uNhKwLyJz5AciefqhLM
QHS90ctodCEGNkteSHu5gZ4IE/3JkFAagQfriHD6gtoACO3k5sPYuWaI0TW2
cP8id583+JtH37UexIQEVOKIQdbk7YOcjjrkOcG1h2kr7DIjdchjUmBxtx6j
xIXNT/GkXtcVfoG8DvIXCcZlrQNpMIKG5ZmZS7ZPAFOcwZfa6z/w5opRknkA
PcfmWC30oc3AhQxfeN50W4xugCzwoFbHBTv0e7Pr4oAORSM6LDxmw0xjj/mq
iS5D+MSlDvBBdMjZW37LpNRwL6coJBUjOa9OnPltjwBe3rg0mwwmLhm85F8c
4LEuRxBUQZQDc4tGr7dGnbW6HA3GPMnZFIgHoaH79JlSSf3ORI9pQzRC/5tD
KVZVcBsFLhvdTpaAbyG9XmLM5N9iYkTOyqcxGkOoKFG6HcFsqBwAytJSTtrm
fn7qX8Clr0rHybKCPN/mrRJ2wKdgp1ZZB0lr+oS7tUXqqIxJwDJTiul44n5n
lbBRwsW66MtqzD3la+e679V8z0/gLd1sPMKXVhJTd0rhyxwp9TPC7yqwGsy3
bEbuWpemKPKvkIQQrFkyNhnLlp11wBD8fTFlJOyCBO388Y2X0xS3MX+bRH4f
mvrOEDlMoTl0fTjim8uX60kuS4kmtuoHDl3r/B1Yb73Bk5eN7wqJyXCUKXMu
kArhgOkhZ1h1kLB86Paij4w65agEcp0hR0T0xnH9Ak2vafyb2LWzQECOLU4r
KqLvH8otZ0IyPGVTj8yvQsDn59fpl8mGyHVsqXwRTv2BNY/FCRnisftV92WN
WvpLcnr92XrtHsietb2gvxyBOK129iWmOH0N5xV5GmEMeNUfdO9RhlUEAnQX
xjk5d8d5S0pcA4DirrCApBXj/kZgkdZfG8B63VHA1QoMWybkHl97SMCMXbEs
sbDySn7RmDybbXKRc5P7z/BjY4LWQTOvwdASxWAYk+YP+Mqg3tOFvzPltzvc
eqYVUh4jgkFrF/mkTyUy20T4DReFReO/oIex/UtP6ueJp+s+fA+FD//h1X5x
53YuY30DRKeSl6EuVPCT+LlIse0kBAITKUbSKks4mEexz/IVLP+0DIWl4Drh
UpqP2HoPXlD0Mr5/Kw839W5xlyKNR20OVahuk0wu8K7UODK/FRQgWjCc0gFd
mH67uHX0i68ARd3y04kOGEcY1w1sASfYKw4uNuOg5nrtzCaLFHBtH/BLHkDz
ZM81GNF26VivByKF5fTOneauZaNPgYtP6TGL40NyZ/xvH5b9+Fs6De+I7230
TOkgWuXrTu61JD9vUc6tbB/eD4KP8NYMVRDRRb8eZapBGGcIWww4uBxqqsP5
Fmd+d2Rpo0x8Hy95Uta16mrste7MWnEsa7xQg6d/znh8RDwQYIQduS7JtANU
sN6PhHRqZZflU1CwbCEphgamyYB0nfeD46saTGluNHrw1aZBtbZuxYO3iiad
sO9Lo3ZDQsY97Sb1NSjzIDVvvkJoLyUMiT1WjekTMrIXM+jjpOjezOOsKzfc
Mn0wRU8I6N8B4H2ckce1aMbT0NlE8MqKud7BJm6NmRVn/j7yEgBIGgf0EwEd
pKYNwUFiayPuv8HcrUCveL8a6LnqkLD7ndzP47ObgFdowZ6TfF1oi6B1WSf+
WtotTKnNz30GiuzChZGEng5BBma4UvVmtQumaZh8FZNNZaMAzOVMA8mKO6ib
toDonijefdgHnQLFHAtDSrmNGASW6ZpUBruKPXdR7HoiOv4gAwgGi4AKcTpP
x51ezRxC+BQTUvd/BBqqZVrfXEZWIWrC0lFg+5QcKA+a2WDsOHA7CLwcRGUK
QxX2c+zJ/X4wVHpS4uCPntdz3rKr6xyZ2lmLHthlflHhX0CRX5m8CwbnmQ35
HwF3FbmR2WvfaL2+jtZmPrl8A8AWOgTb6QA2SEsqjvkbFtKeL11nYYPv2ZLf
wWc2WhKUHNfPD6tmEjVHqaAHseJF98kYKm6/dLd2WoEnzKR+F0ABpPXlymPN
wivdMQ5mn4ZklMXjXNuZDM01tGeikx+qvBm+iRCy61s1QsSYiC3vOdgyxUP4
Zemp4Qr+wZaPalbqwkPB2HnbGlGipqNTFS2LBsGdkZ1wYEecRAxWP2B15t3K
LxdwKZfcnXbbu/hInoUG9FS0IQWu+wk9+n4YGPwLL19BxJwze+Mg/DAC/+Cg
7Uw1cebukWk8nICLLyH7zl6MChJSmPJXTFbJHrc1Z9ChhQjK+QZyegQ4htAm
A5RVGGpTamE8e4RXbU1YkTC56CFympLEeiA2fjOeEkoPKKkfw9HKv7i3elDv
L5JNNUBnxf5z9PiHnU0VXwm77gvwEbgrQQplYoDRpFgdtACIvpk5NMbG+7iD
9jqQQzTcwhiscnUBkrcJDh1q/aGKFJN4INfW3ZqnnjGE/LqnloCPFEHpihtb
KsmvQ79+cf1HZDjg/kJdAyVGawWDdv1adXFZrfignIbQxt/WYOZ4v6+ealiI
yz4Q5GURIoEfB++VgyhvHX+POYY9IAeVBHd+LUNXRGzsSOqdy+NQPbI5GTCA
QzRdktf2FsZyorDeqkdlgKz2PjGWqn52eCMh3tzBItAhTPBAb0jo0pAcOQKH
EL3BSF7LUGeB78z184zj8ZaD6gMUq3R+fi8bCkAeSf/rsa4uZYLuJZ3R9Ob0
Rg5uBJ2uRLXD7WhIGmViznJ0v0CZEu0NPBMFo9uyuaw7gACAHQy0+hqcoqe9
oQlr1S6vRM1Igtuj7zEIRxKkWvYpzW/0sZBzj81737onlwccSvBr43NCGFoL
WPIBoAdfr3A7FZ74OY73wC5vy4cPQB5ihSa+vr+V+e2bynMHauMApaL365a9
24QsO2r9V4WS4mB/odkxS8B8b3WSDD2sPkkY4iC+NdErk+gYS9KVOD8llz1O
o++Hk4IbeunShZtdBrN0w2WkSDYpQIFtkKz6i7Nx1HMFldaePECleUwsVFMu
PN0FnVpHFtLptc2e7/W1twHYIkm5f8ZStbS7B5LH6k45AjHgCIEKR4Yr8C8y
1xC+kmc4RLvJ2G7zqJUHuyH+FOBDcpd7bWbdEDBK8PfRewFfeb4lGq3A+k5X
O5rPKws7UdM5GrHENq6UdGPD5udayLCYSpI5XGzoUixDqq+40tQuzR2XJ69a
r9zPf+YCIbU+WKvjSQLseWLsiD5zFfsAIW23LEFdQ9BDFej8rxsb3/wQGPYM
Ku7xVsM7jSGUEUfBl3iactVIYgbsvfr/UoP02HEID2irjyv3KfbwajMBh8hc
Akzv3v22+0z04KqYoaFRBZshx+i/ThzbkFoTz2pKqbuUT1YReioMXeJxgSmz
L8gFzHCsbb9WzK2Jg7ysQ7MqM1k122djLJWdZmFMJv1SB0eH83yd+FsC1IsQ
YZMS+4IpfXARJdv6bD+yxe226HfHQmxaINc74WI5yECyd5alzE2Fog5qSA5F
RiZTiO5oCrD9f6sQX73RZXXOrBq/meSfGPAxejZmPS+LClZU4NceBPUolOJ5
7DFIaACbA6xP6kJ8U4GsV46hBHb7YAMnPDg9QT9nPJB/tLwXVVduXoqpUMhx
jlN8RUPKgLGykT1S0G6wGhRURIhOqp9zMUj8jPmwR21rHtr+OubOlAllXiZ/
x01U7yGtAPMKUbytV9s7rcvfwreTod7KhhugQDwiNoh8qV1eWbY3J8ENqrFq
zTwWkVnU23ihgU91hn5dYzZUJT3HvbfHhtifBifrl40a3TxYMG+87QFnjMIE
ZjbU3Dw4CrggqNkoXeFm9NScqObKO2d8qThaTUGyn3IHQUtRK4aKdcXPn8Cf
mdgYcTFmvWJjQBg8zfw58WeWdmiJUqa5LiVW8ID63/iikIo4+5lVvcD/Cjzv
i9tF3FzxtBUdgymLCjNmyuc3FRy4CtQTXgoOeEIoIesM+VecIq8dFtj3mw6s
G83HK2hR6lWRKq/7Ex4DghkCOQnx3Yb3IHKK/KBSUsoaQeGpV6rRkpH/pchj
RdWlt9vHFMkDb2O6OM5sCLSJBB568evjpPf4w4d42i0RGf+bUPq30WzQMtrN
OOEi9e+B24rrVwQv4apIIgwrnpSRGCTqZidiebeNnWW8Pt+kkz36dY8ssD14
+sj0hF3NJBCNc55pIO3NDLuHMrQ/mSf/LZieqouolC+JXxu+eknyo6vcKHK5
4p9/le71hsz1cdV9eVHeo5jNgGzP4ix01zcSGhlk2CYHnFKnYxWGPkkkvUTm
3qT6cirdLQew14Md+a+pJ+xks5mfojYXmHu/Q0A06cnstH2/E/8pjaNuOEb8
8IX62n9B/5b+LkM+TOR5Rhbvf79G9+Jb9lXbGW/4izMHEtaYZ5+oM2m0Y0sS
OiGymXh8YcQ6Poqvg7FDURRBDMM7daFLbI/PQ9nToSwgxWXSNWvKloTx5aap
Moh2/T3LK18beem7+Bz4vJ3GG+LKH6DpLOzbTcp9ospOFZ2Qkn/wqFtFE9r5
pvv9ulHRX2D1fBNXWhVY6trE4WgWjT+507GiNA3nC4uyxmr6w+isMw0IOqUn
oixJ0gQMWvE3ePSdXBvLLScEDjhnKZ/gRTfCrQJPEwY9tI3qlTYSqZleCO0A
d4A8ETmD9AsyHsp7htShEoDoXS5hV7cMmcN8lKDNZ1rCbd4Colrk0MwI1aDb
Byy19eta0wK4hEAVrmswNenO5qbIHhhsB/71m/KQpCepjcpm0tb9Buapi62L
UQWlOGjM67N2o96DU9l+Tp0G0XJWojRn3UHqbnv/AK4S/vzhm10XEkwRBX9h
B8z+uvxMCRvsH3Eq/BvVUvmrrQPts9qSdS7A99WJJo0pMfIdNqnMexillky6
kDN4VMWJxL3wDWEksDe+N5G2HZgpbo+XXxjp3P/vcYJDjnIJnl8GCHye4PBz
jH6nVF9+BppWdFQei1nAPvVgcBML0emg5Xlt+SliGTpfAvqPp2tXvkzJgZcv
ttvWG7JLVbS4jqEngMVoprebI+PJ0AcZGH0LqNd1bXQez2zHeVOqzVwyddjH
XhgqQomz/oSlIvjzoKApgL+854INsNXo/kg5FRl9o8lnAeHaVEuq2Zwe5Wl+
3//7yTo1eG77NSbWqFMABsBd+ZmVwMR/caNpC+Eb7/C2/ZzlLIsK18OAjbcH
xs+SuXcdPX/ozu160mcWVMrKL3ad2hNNfLmnfNfhdsA0Qk20o4G0fuO8nOLb
T1MiYFbzM6RNpDnyYsc5rCKBMvAN53zGrVbIOEx7Ut82TtcQCrnjQE27ugoD
kjJQIpw/NlRa6+C19h29Frzq5X/37sxHH3bs6eXg8d8dbhhK+PBrJ7wkFdUC
CQZiG1AGFaN6oAOSD97sdZ0V0sJsch/Nsaq58GHRNTnC0x9/XvIlAW24Y+wJ
pNBc9mxvprytQTm6a4fydkD48biI9ZlZG5/alezOSygUI/Pwy4FO2GweKQdo
QTvcwelMercO1YlTgw2xLQKEWSVbNi8JG2LmyQXpQO2UUytorFbW5c1pnlmF
rtGo3U0lESvrESIHiyyO0tBGB28IlUnXTZORRk19Eg+XX7XuSrhvoF12pt01
VFs7i4VxKZ4EG1LD1yeHV8GcoOU1PcW5qcTJDT9qcMcaEJ4DjvC5LvgC7o1+
yyRmllmZuRnGi2ri6f8j0F48dOXL3apogB83wlqqdeUio7zVzFaIbSItgjos
4/nLvnbdWyq8WEYXXvo6UgeyAwnfKxq6JRg/6mNLq0H9ngodZJQQaquH+Cug
xBPwo2sZxoVfdzrpoLt98+4vZn/p1BSG2STxJh9P8Qu2pP9m9qT5TkrA5sSo
xzk+9VrIj97/Ev1LzFUlrx/K1Y6kKZeApS6wnDcdE21yu34ij65sgwNSLkW5
TIIY93YmRxZTMVAGg87tUhy/YONmLSLmLPvJQsyhiN0OocQbVW4GlaQwmz/t
ruVSPvcHv7ounkaaG3z5JdEOrzwKl52IW546lCU9IM88IwIV65E+rDy91VWs
8z+Z1ihXwRS/kdqy4CKDW9s84q1KD5usOkJAO2pZgq7tjMtOZ63aEW52fmqI
HI5eTvkas9YfK4e9ZK8dPDTJlb4TfSFhP9aMT2pTaPaXfiPNH09wMjNjuzCX
IVBvKmSA4Y0dNXnoLyRdsx0CAcmVq1s6CcsjHA67m+rJHD1dP/Svd0cNt7o9
Zms300TB9vzdPTYff+M8MnCV0hb+f9lECq9KOvfUJLYaoYcTQsAWtC4ImES6
ABUhKUWUqRgw/Au5uiX5o3WTICZFKhOMUmY714QyVxgK33deEOXvoFQRKKx6
lVCG/vw6waR46zS/ZYRQqc3W2ZHqSP3IL6k2NRd/ubi53lQ8vslZ0Txnncm7
o1LmXPt0rkBJ//SUdBZR4lDJnKSt7M16bVB0Mkvu3/xjUEGlXAb3615nKeQe
J01X58HYSHrqjU5JgZ9cPeOunzqJuaDnAlVIWhwajIj0C1KVN2+UUP0oq4er
JAQEV4ItxRBmpv7ZQtDOGBzq40lHoDvx8QHAw84fa1dBGs0CNvLKq0cGZDvD
mRhYN0Fqhs8sQFUcRBEtfU6iBtCNs63zCXR0qMlewQwWnk7aCQtn2bARZ/bM
eHNgKIyaaESG5K7AfLivlAd3QQJU12L2lfHmLRoVBfa18kzvOSlw37kncsy6
EULyaLMUBR8PmEQf8SFMTWZPrjTovqgqhMizZWdGGgAiB50aLfRtmhor7A0r
LjcBq5B4gJQh2Tlo8LY8oBO0FPOWmO11LdZxMiNdZIsZGobWgyhDnR+lRkXE
C005moIV0rUbdfQAeeMhSehvhc/0BKE5WVBFB8t2l+IUHPRMWK9UYYfjh9TK
/RAjnJIJO2Px9U/nh405MlRMOhirAaePuBphz+BVFjY0X5a5FRiMAYBsqbe/
1FZ999EoHTdU9lStQRpUCYlrtj6SdcL6WRT6XCoT4yGhH1EyANjNWGa86TZa
uK2wRmzz1AMpK358l7S4wbgDYWK4FFpmmFDO8LMHd2xCShSB54P4VH5FiHuB
/BjGU67VrAaH6A2uj51FS0hWYn14e5/4lxIGe29wW2EK2bQPRG3V97Zoxw7b
7PIv06xqrGDXCKdYCNY6SBB/qWeSrHHd/Wu51eVx2L7V5cnAZ0RsQu1JH7ok
bAwWeZOy+X76St2cQynC3KjL9qGu5tQqnWFPUl1SXQahc8bUyGUypBJquf/e
QeZtUlKrCfH3ZLC1sU8iN97cG8gcsgm0Fr5+W4QcrR0I9kYB/e5MEw8o2yx1
8XoHTu7O1wM/0xmML1vsAKMGBvIv6sQQzOfYfaraW+dLs/N8TfwchAaNgAsV
Nk9GdMwHKtUHF3kYBT3ndnNLlfOh4uBn/3pfU2kOHomDk3rsjqK28brnQ9tF
K22BjCXXk0ig8NHCPiYbNMxOUb9q3MveposRZPN1xQ8UZtdCcU+ArxZQcks+
OlGqlUG4ILTgz4ojFG/QxtL/ne2XqYLCvZEt60fu/Ja+5NFhOg+opadoXEqH
hTT1U67+w9VEwkESkb+KBZBgrO8TT/4WTJqDlBPr183IqKMiPrA6Z0TcaAMY
wiiP9C3X2pWERL4CgnHN8SEM5OUbDEQD2PUM4jJx05F46yCTtT66O/pEwfVW
RNu1BW/nWYbetpXL8Niac1rYIAdaGNZLzEy+BrL5tRIc4seB+M7Bx6Dll+6D
Po0T58gvmy2S1ooeI229d3PTCW65kW8dtRJKH7H6hSph+G+KLI39SvOXk7N9
IaygxE5xlZOU16MOuTYSpXGDWYVKO2X1Y1ClFtYa/dLZ310SMV7VvbWNCCXz
WXfg/eALH+bAMF4/fqlcK7rmf9LdbgPcboZA/t6Z1p5PF6ImqKU6JVru6rkI
Lp2vkIMDpa0qipnWQj/KZ+MuPWukWzE5NDkSTi5R2kCLHYlofZ7GnFbsrGdG
YF/8klBy+Pzz3QZQ95Eed5C+ZgFQbqECTQ/hXaEX6ma9490vbpjLI0dPRV0A
3FNeiV+fCvCQzn+dNwx8L6pIQtFYMxioXrc8AjUVV3Ra7Yli6RA+BdDwj0pN
uCBE9EEYQ9C+PMHcE5NuikK+ha4YVpA1/Q9Da0unLRPt+U2uzAuBNNZo9ysQ
kJOUc6bEuzYO6SD3VkjmzBLX46lOSLK/o5adbHW9lI/83PlKeSyWU/ZJI0rD
cXUQDmKGvkUBlavcLN91Fz/qGGSgJf8qtq0NQX7IKGvPMrK5FX6QbSJFn/x4
5MEJ8rbRWN6L5x6RTQST01ToPq50a+Dt0LF6W9jWK2pJ0848sJRNQcwKmMp5
onuu3qSym5y4hDAEc78ALkWdJ1sxib8s5uH8MqJbQc/X6E/thuTAUueBs74m
QuHbEYbwc6xH65YC9fMLe2hl1HKKIiOILwWlaYk/z3fEIMZfLUQM3K5vLyzL
amz+fl89pxjWqT7gmSBt6f4Xz7BjKETYp3Hm6dnWabtrhU+4teA2wfGT3VUl
QXZVDL/dlu4zx0URKrGdnk9QsWugdO2LcBlVFiPZpRnl+zi6UP0gPEasYLXA
a3sIV3KQznoS2Fkw1BiMcT0gSjoltRakxh+d5qaFPXRa5ncbwDfhpgu2eOfx
7BfeRduRo/6RYVbboqVT+gpKlpK3q6NTk0vt+vm5jZP2+kAz1aWIStYZVajh
WnyTcGpsnmzp3A2nbdIa73sMZcCI/cCdL/3FKHKNKAtQmfYS1Zx13p7uxU3j
ACiz+1BFwgpRXbzMbKAMK5KDpzu11TtkGlG5+hJZ4N3F11voIXY6GXaPRMoj
i8FAxhg3slFclS9oM2mPCxOPzLrUfeUlIZyJVp9HWYmcKXpmit+5YiUIyeAF
2fVhGfg29/ZkP0t/Ow7r9zpSoS7L2lV1gj1d6grINzNs7QxH8LjhT32ilO2o
R2tfWnFOmWWfDFxmFdPPhsdO1pci5lumRuW1U55b0F010mv42Hi+Gboaps6a
W4VLFuUDWVJ4H6Bo5RalwjlW8g8O8DMUg+3leHc/+7Jbp+N1oByADLNCwYVQ
WSi4RxN6+R3Vbv2SgBsLlcBHPSZvmD+PPylDuCoSWvdIUPadqGfu1sOZclA2
8bK2K536P9yPipfq3Yi07JtZ0vHD2AINXMRLNK1I/5PQjVt4lG7HDhe8i264
GcTb+SCZ7pZj3HWduxp3i7hsJizyTrlyBSoixtXDEDHzNr1S7pzr+lCs2aZ8
4pbl67PYUUV3mx9Gqow0Zs5L5PYpk38XXg9gjFuta6xIl06nw1cX9eEKL9TH
HoWkZys84vDun5pwmVFrb9zZQV8M6XkBPNm/dn9W4pQWK2bYgUtQzKCuf2Wy
Yx7jJ3sC8heLd8283YKR/seTeWBH8j6L4q5bD0aSwj5y2cALFcTYlHoZcjcO
2ni1AxqOiANzEUAjEzqAS6gVktWTHB8Z3/qyGoXiDCXAtsw9rknEEtbeGutf
kOSGv9g8zl2ILKi5L/pmwVbrRQ7xaLmSB0Cdquz0RHOkePEhuwYjkJHQNHV8
B2EOsT6A6TxXMV3d+phMKc60tl1sBuZsq4339xPhZL/FGVueYe9/7j5YHMnq
3+DjLywpZ+WMapr43KwsvRvwxN0QGBrLz092cOAu8PCnZLRyUgUfWvD9bNhG
vcrrJAulBSh/KCOxQflmkiExRCD9Y1U+btPNZs5lbTWFiWhjl96swGCruvDm
JZdWfRlzW1pFKe5wIL2bJ/mAXtmbXZWjo6c1kdF6WG5ESotwIRxtZZoyUyxF
V3dV/ZcdJYCrX7UUhAjaPt0yO6/GBOkanTTxdLVnOskhZ57AiTePBuwgRIWJ
1/mUEoIdBdq3tbKbAO913ngi4EN3nOcHwCv8AiwIebekG2uApaZOVUYFFmks
8zBwqcGBcGfzGilQkugvCKi+4QxySZLuMNuoU8cttdW9HLcsE8v06h/xhYYQ
/SDf67q9P39iBoZWmeWo97+sJ/n4DrcQSWHmNEGlyIAwe/kkU4RZbTTtTbQX
6+SpLF5D2FxyXK5nL3hsaNVjLJ788Fh5DkblNREBpbHyvtZKf+/iSLIFrp9B
TEmnBW8g2HayNbxmGQMCVAMrgPqFoWrNIsYFKEpdL/NDnsN8EVD26B3ZvLYF
dKqSZpKz3kDkuSbMXf2TZFztt3FRFT6uxrTIoDepvtA5OAy9PZAMR7K0/zmE
g1diRQdHhImxgzqeUXf0GrOwVbtnVoN9x7k1IIOzUuI0zT65fB+zBdBHTCBG
H0Ba1WfZ+b567c+Yyi/XqvYKJ/x4NsgshZz1332L9SEEEuxaO+iAofoVGn/C
uCOXvEBtTLoOhLaCehVBRTVvVQ5aEHS8axcccZY3SEMwslzv/Pw6TYCYWMqP
ZK6Wt5uTJyX6mZ1KZ6j63WOCD66LqBzU7/C85I7+snGQ39oD76K2D+CDuda2
+QNLyNfnegzKIWhoEjbVb0Zr3nZnZkNmIjDNFTMFY7r6jPgyorWSqtWMGBHE
pDJhUWjsBv/prcEt9y7/oLLqgeKVk9t3X+oYVvajk0jOQAYzPRqh6V29zXs+
4gHKqmj8N/pTdUIkLESuUTXfylP4DMS43lHavZbrlfVbkj0oXwxk612rrN6x
2Ic+G1gkNuYbtSmUz/O1u3P4I7lRh1Prdw99K2m5m3kiQkVD2UiGsWf/a8o9
5eA6xDX0mhLs0fDMVFKh58Uhx2StA8K5+GUErfPeYnsja/imU7Sby2gnjexO
VybA6Z6MzY2kBQtgWcfJZabsJPJJKupD7NbFVxFppMb2kS5QjRLabvrqnE5R
2ZHE7MHC6WvX4WFmkCUJmK/jhHsGZ7nDYOHkYVYHbkJFkov+CLmQCOxn0Wia
bijk0fD8QOasNfsFPGrBUpi8/mxpGbHmjNuN0IY4Va0st5Vc0TF2aXht4lyB
t2OOrBnsfRL6KtJipeZZdICZDkDCB7V6kYwKFdTXKqfUxmQUe1hG1Xd/V2OA
kO7+wRzk8dehn2FZJBK5TBh7lvg2lQHb9x8JGBt52y1HyslZf2xBUauEUdqk
eAZzvHQ4F1Rx1zc4DY5gCSSUkHu4GGFegEONVVRv7UaNq/U3X9dYu3o5VoQe
eo62ReJ1zpz8AjhJTcsfFmQdoy2O+n/0aJ11CRiZ2popeHLemiw1geM88CEa
P0dUJyxClbJVvV/QHDaUVMiW8axmIxhNTqmUIqh23gJJAf9MUYjZanYDodr0
1crZT0xU5oKFPa8xwvhLjhLgcuw5FXYv+Pb2ifJyRaBu7QCS++NLnOVNhwld
iQ/c47KmMbc11AMa5eJ0AaAW/BkEZeLaatkVbWza4H3KtvgKKO7TyHBc4YlL
sq8h8kDKIBRcpDpaNo7CSxqPidie0/Ay8yEY/k79rI3iw7wuSpDECegIBx6w
xL/MFQ3AUWaoYGzGZRmM2bZ/6QVzTQ+qiEwIT4GPurBxbOO49wqkaYVFQRv3
go8Cu7UJcN++2jiTFUMyQjIb76UZ8EH/15hwEsZSt9j7Mk2rrR5rbW/Wz6gO
L0Zf2IZ/E6SBXdZF1/G0BX5C0ByKjmfbVmBWwZHQBkZsx6My/4k20p0oUs2I
/+7HQyowUb6mUgK+jfSJvoJVZPTrha1/Gf1/Ce4mH/UqH183TZKNcvA8EiGz
D6Z5Nsnbm2FsCJp/Rtuqe/t0gIrL+rnIZqJo0Nq2nXlPoO8xKNj9YfTIpvSR
tU7BrafSbKj6Brir0Y0aOuEYAros47xDzfK5F7Q9ObQ6hvqkTIQzlOoBI0pB
FDb49I1VvV9IBY8r/xDpVW55Iz/k/KbKA1HNuUt2gyiE0AF/gGkdV4uDsjAs
RmSXbtfIAQLcmQFKR96amgBsWyi7hS477fPg9KtrAcDiCyyhxa1VB32KCyXj
GN8bCk2OaUwnBKGaHT/YNcHPPBa0lNimKADcHtfUlQrCbc7VXxbOuMAztCBY
9ybUxvR6PoJ+DyeNzzEWqFBEw3620gZAzwh0UjpTLugJ5Tjd5V/tWZYTtTQ1
6RC7OC8aj4pouTLQ9oMFMmY6TALZ9J5W9pFFpBq6c/wc9AfykHSu0BSr1wSQ
FsynmhuOn6h1l6dR+a9IV63gD4/Jg38r2Cc5nWlLDZwNYpGRWO98tBf3igBJ
EHKDAizrW1m1mo7ljm0iunarWc30ioKSSu2MyOkIVyIDufkgl3ULM4ot5uuh
HJPApiC4Hqrp68mlyhf8VDaLxfe/rdpfWEzL8ABelK0uOvqbl0Bb/UhtTPxk
24xCEc4JrwawLmWP0UPPrXy+Zrnu/x84A5srCOpB0JyiY5ElUuvz9Xz1VzPJ
lOOQbgDk5739wu4KVRDqGHzwKniGCUTW7ZyKNzbZk7nzMpjD3PwzMbpcgkn5
9ha9/9KPFVaBeBAZ0z0ef6o8VUbJNi1rZJBn3xehuE9uEiPryyCDd39CCtQI
ca9Lc27b4WmDw+g9Oib2uWCfGGcQepYVgsjm+PqYZHj745Fv7dPvqkwozyNm
foRUXk0DezR6CiMjonOa/vxdNhEkoknDEyTIYbBBEFRO7GP6mJiN3YwCHw3Z
MxNZdHNSuXYfoQo4BoVekhlWp/gg3Gnf4gzi1k+o3zB/HN7QUn8sSlntZZ0m
PsEar6SqrJxjj9giuxXFudvoBHh1byYQ/vkuneMD2q+zWEy9qEync9itpdpo
6IW/67dYCKbXZHtXImvYQMUw/L2pVKEqArs2KwHl8GVz09jZ3FfutmzvbUyV
EoDIVLeKxEUdtKJHJyknG4E5BpPFw+g0RHKQxLyosZtjWPZ/gVZFst/LCEk0
4LgNl3CD2sDi+Od7eIN/5NuXOwD2BIVbKDMfuHkYUw93sf1ToVOIShc+eFDq
eoiwf1i5dcGNBeX8hwa3N7iC55gSeO23U8CMDnai/6A4Nmyp3mOwqLsipU/t
rjAzb+3uLXwPxLvyTchVUpRVVAh7uoNKSdto8gBVFOVRoBw7RBhKELoPGdtS
WoBMyI4OI1ZxPlTX7znjxsKuE1qLQqSogx4o9U/DeKfEGQ8c2P8Km+6iUYkz
TopjgNeDbjtznjMjC1RHgDfovwxoqbx8MjsNVpsh50JTWtsNhWUGXYiAChes
4mAIfUlP9qk/LiZ3gf22ScHyFxJ63XE18fjSeKhjc4d5TzpFqmcG5sOfphTa
4oOihBeVjGsc97RM1JJLDH/pgrq0hO0FyMSWJWko95Jjcea20Yyhaqnyrqee
EoiSVNMNJGmI3ZaDQwyVBlKDHA5Zx4rWWH5U0kphuXs5yVPc2obwGFqlBgwr
5lA6tphRUA3QdvIxS6hHaVsxM8ZACfSbNlSYNL7yRy6JyoAj5QT1wQQ9yZG/
04H7ti06yHB5B9OVL0ULwfvF2xhl5jKqNGrKvJDLPIROmqwN1/X38OzoH+Q4
O2MrRwvVEWHeAhv7upy2HW/OWvU8Oj1t7j8UYME3/qSwX31XlQ6irasQEGnc
5MO2xUma0zINZKgTiHxWru/TY7Y6qoEfjhHpiK3cx1jtrpAzVjHSaL+jgUTq
G95MJIl8ZsmeSZes6zxeXaQTozlXSAelMK/hvWago3eNTixmAl/SyyJF15LW
B6un+QOIwzYidfi+PYNL0TIIEB6b2/HTT8KeigFK0VofCfIzxGKOWfY3Zq50
KeixDkledtloHTyQSdN2Ht4rTpLISqJBRri+ZMl0XE0KqaMClMGao8yyqnUD
nZoC588gfXdeoTy6A34hdS/889Br3VQkSan6KuXYIaXvxy6PtaSGW9wwn7rA
GHmFx8SW87LW8Tj8Hnc+asUrdwvCTbDyLWEffmMflVSXIMrrjUQOpMDOmhJb
FH9a/iMtaoByIGQWHC9IuzSK1efREzOqFJWxmM/urLRwXeGSptp8T8gCv1s9
JOzjH6Vmh+KbezLekuHLrbaQha+6PArFGqZqeXIFM7maBZpn5ECU5cak5iHS
TH2UCtFVt/Mw97Pq3DqUpc/CwlSRn0QECCyP9prf6r5lYpDucnLRS0VHOMK5
BEIq0oG2KGAPvnk9Fn3RpybnYzL932OsMHEMgRDoNrrxbK/55mzU3ZGUBvwb
RwfGmbbt0hi+r9V/KQiW43EyMbRyfljLVyGrJJoax0ippHR5KxbUTM2YeAya
zo+EV/nbIApAjcQJjPFQIQy5+6H2ypAX9tQG/tpe+GsMSByQCtmwwBCf9d/S
JqagNlLUogGlIld3r626QW9Z61p8pNZE6tIEa0ugwqkrYM5fm+nOcptTbFx2
ELFX5OIoHIrsiYrD1O42e4A6NDey5Q3QvBbpNua4O3P5iltcRrzrK0t1ErHu
uj4qXy9icPWc/pr5utszvVmyh9cM7KcHxGi47BG7J/bMhwAT853a22ZTrR+s
xleshAGH++k0g4gQVxt/fTp/XzRGxHtitBN+427THgX8/A6B+VfmPcZhjZPx
MaWfqjQgdgWmtYlcYuhzly0aG3DwlU9/MmMoIzSv1PEzy08mU5OPM4CF0n+1
X/NvslWkpvAbZkv2bI3I+9f7KzKI3cdAqh+dnAD00OLMxAbED6H67dX2Qf7J
IVtXbmNyjIA9ext8bdbvQP7bcfcNZQ5fDUtp0+lvPzlhCnugKBOUYG0MpvS4
zmUc/cBCTdspxzs1PokWIw5WZ+etmx5qpgF7KsWBDarCJleprGFqVMZXrAmN
w68RkRCaHUO4anUp/v62rPHkvAw8X+M/IppQDOZq2jAqZfljaSggMUlxAd+F
+hsN+P+Kh7FCPRligZIMGAZ14Po71Qt89SJiN6F2aTsaXhIOZL/32dNYFkml
fGVayRHstZCwXNr10gVAIySYviRlMc/5iawTCGs4KCmBm5I/OuxZK+Cj+IS/
4S3hERm/Rt2gqZvquDxrNgn6WKwKp4AFWUfcJXRWuw77IqAhRGe4DIT9kbbX
UEouTDoUF/uyPEvstsCiKMKRTsPyPcTbwH83h6TIDYdpcz0eIaKK90ONnX0N
o0msrYxXzoi2uswpfuRWaa0F+HHCcUhnIw6psPoKG9SX5Ypr8rwPfAre1Gpt
cOpTLh8FUVWXkkKkb1Y71D3FhIE/GDEPyIaS87sBb6/6WOvjmM1shPpYQxpy
lIgvY/DnolDWWSckAbLV4bcM5aEvByeXmNVE3ttWI80b+HqmmcXFcQNQuRnI
fT7VLZ26shooLG5mVpmc+AUAold2y1WzsQohvdEbwy467c6WAIGeroFpmsMx
QGozDq7jsyEo9dzU0f6S5rLxMmNqjFjWn+k4/5IqRcFg7pnlCBsSxOFBsUhi
xaWNKzwTMjdLtGSWqrZm05vH/KDLzqvlGdWLCoay0vxAUqJMl9Lmkx03aLiq
4awSHE+0UdMhr3v/SZ9ZH/7KBKgjsjmdmlKSCkvPhG+KvwrxHzFVMog4EHPc
pn+roMEty7GarerDDGkIKkjphnkS8Y0eBCfHT9JGqkdPZb2zDFCnXrCKo0uW
bkVuDboBP8hrc/Kijh2CMoyaoo2MER1UrY1LphOJcQFK9PTHKfwraLuc9nNp
jpmUCrIyFhPrmqH8l5HnJdkumf40Ol4oyhTgdB5XY/3+DOFwsQ2/TmG+MsoH
VhXwOywNea4FP1zMNFH4qds7JxVfNnBYwjLVOl02vvf8Flb1a6MDzIudMvmU
iKUmT7d9aL/OEyGSaZ/qLRKumUu3mGBqLUAIMvco07BK7KoV7oVweUbI6KJZ
qYxQiMPP/WL0G8rUFvFD11FSgfEc87kQDirlKXuftlhCozZ57CMQZYNQE0WV
EB/LKbO4MBYcXT9dMxKM9tABrt2tJRTbiOk6tKL2r/kEZzhK8X2RWyxAsJUQ
1/D8xLgNFP4ijHsxTDtcKbK6qXnC/Y5csi+AEBOMNojZ6uzS2BS4ZOs5PZAd
VyRX672DCBZux32NVfp8ZYahG+WOBZ1tVVWCYyYSNi4isHj/zYNJY48jCUps
lxF0JL6UYeN7jZco3h77DEFHW4QnkmieeSfQc7TOCHODMSs91eP9xPbW1UfG
qMd2fxb/+vpOONSP5LJaB21v4NWykhnbWCb4Z1izLFe9agcyU8VkUacraRCR
JUZlyb6W5zQDmdUtqDhu1NClrKIVpxb+0Tk8Y3a/cTU9lD4syxHArOVUC/9z
UuGa57IcFmI8zeuVsINnQxjvGsDBogKg9n6ioXBCb8N+2G8hfCumAp9Ax6f8
6XEEkJHWJwDMSwn3x9HKANXvE7GQB9IZSyT58AA203EWkdTJ5B2hZiyGck+f
m38Np+KQhjH/D32VoxWNKLflkYKzml934V0Do570ABIOrFQ5Fbmzbu3XrOn/
PkryzU4HLEieH7XGsuH+m+1i9vPIQfAW1cBvL3EgVJs1J1jjzXtLXyqK9Nj7
uFX1aHUGNjSrb3LQWm627zTYyfe1Tpbam3oZ6zPMurWN0oaBO+2u78/s6tFO
CFU6G4DEkRnmWvCgQ+XxCa/ssGoqo6ZeTnleyF2RHuTmwg1clRDHizFfBDl6
oeJbUWb8lFiz9/07OzTr/nFqMcg89VASmn6LLZNtCkOTwt0nWSlUrpI2DHWZ
i3fnscYtu3RpEveqeULep0LnKESve5NZt27NrCpQRr2pKpq3f2vcA3cG2Ou7
VFr2sLCLZnIFWsVchCHQaCZrZmX77FzawZK8Syk2OZXVyRMcGxpDUxuIwbVK
cJ1T8G5Ad6kNfXgcYk8v2K5svYVF/DLADq6Y3FRYlYUYf/pfAxwG9M/WomOf
aJO2UIdLLy2IP3bbt2cMgzIkmo7GD91PpNF55j42gtE8LeqTmDqoeTqUEGEX
GeFgx/MMDKBnvg+hat8JRE77MZPgmyeAnN/skAqmymE/zHk30zyJNtNo0N3q
agyDA9vYx5ALPo67xp41TDMV/8wl0CWW9oRtf0xIB7Q8SgZChQHtfwJKuB7K
7XU3X9Hj1ZzhZ91nwJw0aLzmlwkiq1JTga0pLYFbra/Y+Eo/MJKZZmDRtJTL
HOwdqdhFeeN6X46hbtWZSgFluvxaJSWgaeATCCGhK4a6vnsdle3F4iEyKzDK
UiFkV7EIAQG6lNuVfvdY4p2a9dwmaPXUQXr7ZslmKTKY+L49MBobmypLSGea
md4YTbGljETBl1J9jx67l8/frS065wijrxKI/LapX9osCCHqghqCs0dm63Ey
t4Wmhr4CiSy5BZoMkP2Px5//myEDOpGzUkWlxur8U6MUnTSLG4Cxf7Sg5sAv
PZOjrSedBCvlxeDBYNYN3QvZgmhaLHh4gy29DKxSdvqmms0/SDpRdQtpLVfQ
8CoZiVuoYzmHNaK2FqJfGHxzA05AljiHUUmVETLUeNc47XO6cFrANGlyAr+f
8x4GessW4B282rD+o93x3FRPLJF75FS31KLHbuNmmSFv2a5K7MGio6WdlAhC
7duHRcIVjVdOYMapk2G9fe0019Wjz5nkcYGOU/7pvDn0lTDbFprwq4dcy2/t
JSjuqtrSaBF8zqijiOHZ+awfNh78PxftnxJMxnd7PWp3Fm4loOcD7ivS12xd
U2DyZz/PLhMKHsy3vDkGW+lhxl1mRTwW2mECWnm5TreDwr0jEy9qwRYrYhpQ
K4JVUFmDWvBnKNpwmazogxXCPv1xGhCaFeUmfUyGg5BD1OYlV9rLyBrb2pH6
rUVmAdI6L4zU0l/wwjmzdtXfpAgscxKbAZDTEW5xWGgDKgCaeMR/SLEkbmbO
+gW2ts9xf7PF+zYF8J602wAqApKAyObmkxM57uYfWbPCW1DTD5CddNLXGRoI
/HkR1LjP0ohMqAkXQ8Eedq/SEZCaBXSC8jBecDBKTkABJEGvqy8KyEduFmaQ
fTxJ1kroVoTK1zOkowfnKowRACu3SQXcGM5uJZHmRV0S/G5XRa0UBEQ1kPwv
X7x9+lO9eONWKQAgAFONZVgAJRUiXy7Zuyjfa+dRYDBSejHKtaVzZ8g/20tN
jp58CMLF8GXeqP1HE6laRbGZrBrw5ecxm408vCZDROt8zMIh2vbrWUXrY26R
uxKNSoHzrxyHrLyxnP3ZW02KkLY/y37W+leeREfvbYdTsuDhb0fkHmBh7QUB
80bt5cVJTMGHDXA6mvZJ7QixXCaaCu0mmJi7LS4Q24H5gv11jme3hx37IEqa
RXL/lFdFQikQwucEhgTRqIRn0jWigQ6WGbzqCPysGNYM/zUXRbtU7TEiIyPf
Pz4jg5ILJeCew7v8U3dgdWeNK/k5rVjz1an8uiQa+r52ndU1f5o8Mz/1vlkp
P6GfdFQuU8yFpE+OG/OH3AGqtdazUlpYJWk7IzHizeFG620qW1qcJUUefBBL
ckboe+VTDvH6eFjmT8LCYnN4b1YWUwxbpE3Bu00wgVtLrEuJsqL0E7enL3n3
Ix/UfEkP2XObEvUcqT8ZLK9wPMuC3fDg1owRo/7zQZZvqRn9TgmgQXewhRKg
k8oAePzoEQKcxeajip/XbsOscc82lhF85X/C2PGndxDfuQhjfhM5enB3Fvbe
XuxCe2ylWDgmsmH/4KS6CjAC0LKdxwbQwTxWRrruCfKMtE22GZGBmwhvhk0C
J2GKjAfqwcUq6qDr+NOYtjNy9v7mfdOI4OyX0jssdiV5gfuFxNVqDnGwOWfR
JaqMsBJGQdH4hhJ3n9oWN5yV9E/XNyruJG6kK9q41fqy/o90TqByKUnPdSEr
cG7B9ihiw+Ue0A0H489zXHKDp9XR3Q3LlK52V845ut0Cgb09G63AdCH4HDJt
3xJ7R/zzKHbZMW3Fr/QmiHUXIWIUc2PpE4jhnWxt7Hm08pkjA/JjbyFyTfop
82FRj+NqLsGmueSdc0zkHcOPRV+g46A9hw+NXgiD9dU0nYPVDmGSkx3ArZgp
pikpyVLI+yOxKn++bk4KBiwbfKx8B1U3PIDo0/PZhYkGwACmIUe3cd9nNf5q
dVEzcUW3IpkrbUXLnUhJZJWtT8iHHgE9J251eisd+pROo9hX1ESgmR/gTTnk
I87Ep+cnl4GKCQx0vJTezaZAYE9tqRFyE0UJoL2w2bBR6vKjvb1DggfkohVQ
aBRx7bs7WrZxuk4H9U6g0Y7kUtJKvIpo5zra/g6LHAv++Sx0ZI7YtM9/Ndk2
OjY4YAO3m/wEKr9H0AYkTzr16+c1bfWqQZCA1DeiAQeFjtLvrplrR8+7WlWh
eo/Een9h979ysCPZHnLee/erl8hj2I5BrCXx6YP3i6zmkmKGxyeXbrgg0klI
5/LAIooRkJoGtuTtqkK0mmZEdhbcR4m8CgJja0qmr4zgmQyBPhD3vMPtuzhd
czeKqYCvR6d6vGbWOgqb7ydPyHmM7vYuHiIy9S3gDSxO8Ob5IEyVcECrcMms
xYtlHYet5pdkSsrYGRqU38jG8EUofa8k1AeB1ubtHfd76keFBUqKEMoCZFoc
mWmC1shrXqZbiHDMIMKaviaGALoprarqHvAST0ZqQAdvkh2eew5A+XcNt6DE
TLJF5md9OAuNwuhsmG4nVIDJ0+EaQRIynHFzqNdtUVZKRYMnlxXhgnIRnpPu
WmL05ZLZHYuHueczEglcDlennizV8xszDx4eZEtz8JOjhgKxriVf5QeBx15G
dfjUV2LJuPFTkUm5Einhputbt8XI2nTcQykLWo4VqDc3AUYGp+cQi/PATYiC
ySHPDAdcS/Fof153SFO4TZFuuSusnty0XQpsaSK9lFu+x9R9AsMz+Y0zEIfN
7WEe9WnltnQuRBHOxBucIoWHA2lKILcQXx8Oa+2DHTMSXowJS8CL6T/Zn71a
6Bh1sXjN40VzdptfjdBCnkI3IeKvBuF58MyzWzKC3tXcij7ZFbGM2Q4plZGf
jgUw2WMNbY1B+BDO8aA6OgH+GSIKQl3fDbZrL/HAl8mZwrIe3FuCXZvjbT+y
zBUd6K1sd4JYSqMcOuxc5kPfgbbVjEEHv48QC9m5JI8iGpne7w0rfWSjI8Ku
FXGlhEfXxomB61aoPgraKtRRR2ClvT9p5VPbu4fu6ne8sA6cr11RI7L8c414
wmu4Mgp7wmO5vdeadIFP60fLH4YRb9t3VG+IRDGnmEBtAfJ8metY5PvOm3mk
rlZdhwRVR/FUDg+YRfv9x4jhJ0wjXZx1ZsK8TOLm6bUWb8jZZDTh9q+Au1bU
o6eBz8x1a9rC6XVqKT1/FiQvt1r5ot99F8Mb47ZVYFKrQeRR3wuYkzu9htuE
lLsw7M9qBRR5rhHLletU+KdQqLRBLris3cdfQru+gt/s/wiJan40pIe57IBA
PpKPpiiZO7Jv+3DrrjHkffMxqhrFusL48W/VsX7//oR0Q3Dg0/OUvzWI5f66
C11ZqoW52To7EsNQNAnk5BSi4EMjzpf0JVE9lAL9uUdQN+Mbmxp+kaNV9Lo3
WTfdcs4sgCA0ER1V4OQYONJxaT8JcojMdZwsVE3VgOfaigtKnyHI2BvWOPxW
qVmzLppPVRqI7kTLYcPhDbhxR0qJDXk74JIPkht1TVV5ml3MocbP3ps7VC6/
E1JiMgtSRLE9WXnjEPvMCBhXgbafu8FF3Z0pb/AvXSxvyXrfyqyx6qR16VBg
M/G2lvy2VgojpQ3AhzlqhgzxUCLsH5vC/vY5r9jX16h79D8dj/TP2vGfFXFO
IKhFF0Q7tHMLlx0wUXy7YCZLOIXV4V70UsHNdxrdQmRslqcnEksCzyOmq4tS
jecKiD2ek8MbwX8GK4SW8emvFoHYQvdmT6rUqax4RrM1oX2T6+PGYHk/sV/z
+gUG66nIda0OlawUXSjwcOvK6fiY95Y5hWZzv7uBYqvt0TSZiwqOfKAoFTQ1
972TmPPeiZR63Cy0nYKQCSZ+kJRCG0OkenawWesX8GYS3+CaG5TENfWzw95f
SrzjoY/RQA9FKACPpyRm1jP5MEmp6ehWa+TxHZNPpeEvY4jsB9YBm9sR1Gdi
vXAA8gslYsPQH0PzNjS7srqzOXr+ky9YIR/NkxPtah+rzsyP+xfQjRHh8C7Z
oUgBoydzcVpjJeZwyWNfQeMJnVccDqkb9dnK+eb/ehuFUzBTvklXxxtS2Kje
GavEd9nVjL/JI2T27Z3KTtaAC8UQ78AUw0qbBcXgHlbXTvgxhECDjRklePtc
5v5M/30aRhzi5xmpg+Ly9Z+2Z8saffISp6RDjulj5+T9wPr3aqJRvLIbewG6
m8F6/CyqK+nQKj/Q2y5WanUN5uHIzvEwkwCtIUNM8YToWGAABllhZNyuim7f
EbJtTFa7S7BYt/VW1d5GzntPdKgyzgEbTWck7ytP8AdO7LO3G4/3Y/0xG5GC
Zu1GMswgW/qT57GqyceJd5y5RW/KmXpeovq2utP5qOwSNE6GDai4MTu2vnm1
h/DYeV5PHOlzv/3d+l82qi+1X1BRIvbOm4+9h8lUfshvAjMZD/x9dy0ZRfqw
1cMAR9LOIvDEPo3p/OFzKYjjk1KuCl1jZ2paX7TQH1PjAQ35DLuxS9UnHM+G
GMp3SAzXP1rOLX+gXQ/ajUO54c5RMT+ARnRpLIr8FeTAjI0aaOaBH3YX9bxC
E8674tzU0B626PI9QV2JCK4voH7FZt/P662BTCGT0zJJ2AqklwASOaXX1JbO
A1bAQgM7fPxAXG+KU207bLyuT5+QnyNSm9RGWO/Xyg2oPlcVuBpTjKOmJ844
x63PUmufRUu3FwXfAmevWIDU2ae6tnwdJaGCE44cnDSIQAxS4AckuQ6rDOJI
JiCHSreFypuFiF/J6OMOXLxcunxCJT5XqCDi01Rtz9BEI5GjkeWNwZdfcscu
uFwEO8X90iTraWvAMZ+B3JRNKfx6XhmSyw1+HMWECHvT4s8m5/6rssXGTDgG
RaJR1jVz6kTmI1PW/5+6+Nd64Wrv3l5MFMxCrdcN+dyKQ2ttNOA5fkH1gMCS
tal1DoqkwNAiVyk38we17oR6EjeFu6OGkWxXfgtAMujAweUbsstOYnS4vs/H
32Q/hEmunr11TXrBfe0Ps/dFeTT29rlUmHcpwSLvsCXt6omv5y7f7fNIf29M
DS+3Co7oy9NOVT0u1ujRNgWK6qunqha6K+OIOnK1IU6uC4Vk6x7CrfVMhuDL
Wn0FZBENmeykH/MqdIv0LUOZdDAK6QibDAn84vo1WUZz7HZ+qHt+8X2RjP5J
X32GWdQhPTIzWiUibfHukQvysYebYZCDwehwyjRLXqzDRQQ1cUQKPFrSBkdN
Vs9zx6hfZh2NRr4QlQTHU+Y0T1KLo6+vg9bE0MiG4/SVPicVjlph9r0n8h7L
ydnQ7hAh8UPOT8IMZ9m7/jt8+lRLW+Y+Gx56Y9S7IHAFwCCeN7dLxZZOa8RZ
6zviJnFN8spXCH/it04xZDxAz06237P/W3DndQI3x/x7eYiyNbC61QwG84YO
qRI7JbrPdfF1QV8GktDdidYIADtXhh7k3qDYTgYIJxvkBUG49cHcZhXuDymy
wr6z8JX6Npu4P/FrTnIsPbx7MRJXdVKNiIfiVu9C1srlwvGijposg9Gu3vJg
V85WY3l9fmmzADSLb2nEpg3QA8DJxCuTXlpKflFotR1r6peDklLOvcVPXZ6i
K5n/I6/u5dTPtp1X+N/3CrmSWA/AzjN2dtIAtXOTWMWW2rvijJPOIvT/PfVW
DN1DSBC3hKpS70kNNrupcFmlyxfV0qDXMlxfzOj5TdiXQqPiXsDWMOoEndhK
e1TNFVtlwzcOH3ffq6WLi6QAsYdcPevSwjaVkzPF2v0vosp+1Zl2iARP5hAa
PXxQOhvVXw3zgx9LOwQRvbfGkG82R7rems8wISTZ1tjffXvHTR9T4UzSu6ev
eKRN+hO2kO7KF5aDoFASqUN11bOgSPSHUy3bFanBCAgNjr4ai5XdioROvtXI
1zyDDvMh+BfU2klxoCB3cll5PbTo7K2haDn3jUf7RxtFlFo0t2J6m5jrJBuH
xdYBIqc/88RL5mTz/WMgr0hQBfzHodBZr12go5Y05fnvxh4mXgiO2oPmesEM
MGMfhpXyz5HsZYygG871d2hgA4+UEJgKpccgEmKRNkqP+MAF8weS3KyaQdpQ
dCbuuVOmxJaWMzVM21TC7quYZ8+A9fyZtOCMzC5fW3OeGLQvlGWQhD/TK9hk
PinonJ1Pr30UcutklIuM6/WIfu4XazZGEoV0iTpXd8Z8sOJh3ODQoQDggEdY
Lk4fpkZenage8s/Sb38Ow09gV9b47qUCIjUeVyCjM/GbvrJdQeP2wnfFwKqq
I2DGdO/JV8lUruI0TCUcSKI6ISnDnClBUsD+dzDbZapRFmt9RcqAWu+3Qfgb
UpVGXrDzEmZGlJChzx8mNlCo3FHTMKH+By25iO6OQWGwd35Ikb8LPOWgpvdo
GuL8szCr4T4az7lIFrpFWAcdhKAWZF82dx84Z6T7TyxyVNX72ir6rzSvVoSj
O/J48vPFiIxe4KIpLMTNLL9RQtkKsggyzK4CfxFVDeWD+SJZ1UA3vWuNeNOM
koDsCNfGeG917EdDFa8r6Hoei1QlUPLuJpMOeL7yEZHjWs8IKkkxg3uV9r8A
OI1rpIkGxFXL3pBINh7ekrfreR/5U5rSvCdjQadyCWrB17oYYvnAcVkjYD2Q
JGj51gwts0MwXbRjcW909ZJ9M/x8zDWGUeUVoZKUEnVyT6vAm0SzpSJPvxX2
zHBMbTInejQnsRXqosqgXAafJ7bZZzz3vMMuQ7jz+nWfAOu2ni6xKW3/rQSK
b+7NHhDyR6yAGNTKKh+V2mh70tK7JmWDOSWoYRKu4/ZPo19KZIDMgoQRzAjL
iGNFtmnsRa7Ts/tqvQ6FWv0Sl1IickZOJSyO3wbM1rvwrVcXm7vFLsBPbvRj
p+Kx2lS0gftcX+Cy/g6SKPIOM2b1YXWJPNSVCfws4tQ9qkw0g6Yc/aYBEwmh
nxBKNXhzMpo6ChuOYuwK56n1UyYlp2bGlK1T4oAJ203uy5687PMzGJ6xrbSk
QLJzkMn1Dz2JajQc1Ex0s/u+qLYOY9OMElhbiq36i8onzp4ijdnkU6Goj0jU
MojdhM3Mcm2OdxAIz+624qzblmQtwt+9VBlw5GuDENiiw/X58QY4WfKWy1ZH
WEClApIuFAN+XJic2ZYRkiJ6jUTc+O1fLubpkI6wE2qz/zFUmD3Apu5g4Ssj
R6HfitmaCbisw6JJFvoemHCL1xitiCTvQoW3xy5Z8emaip5CWPkK+7pvOiAS
Xkk4Aec74E6brMuXIfl/Jv398KSJwvVnlVXbPNvGjS1cSB3H26plnP7BQT8t
9EUYiVW34PL6W0zdI94jwpJyirdCcLjS7aKRV8NuLU6AVhsCvTasy8Bpa3RQ
y8aoX7wJWkpU3ZHIohW+KsAtau+EbxPvshxbLrwSuZJCVOOSt1l1oYQtCFiP
te/QOvYy3liYVOhB8LzaD+r9c19CeOziFjMka6oO4561hr6ixRwiAgETuEGM
tB/69BH2/3hz7x4XLD+y67Y+keGwtyvA5VTUrbFEgC54E3jhzAs7Td1sKEk6
4aIU2oIzJ53Cfg+noyNmYBRNsKHfTbMa4+5yaDPImzVodBWQtgszEptH5oTA
9+Qp5oiKkk+nM0bZf1ZgKg6EhLgxUg5jYbaFVLjIBzJjKUtSVo7nzZy/1Whq
ifxPcfq1b/Bcjj22jGCxyYPrjjtgUN1IlBCDIivE61zfJLNeMnlNXBaW5cGM
5+69wMzmj6Vz0tbsP2I6LpLscvz7vmX/jAFIp+7ZsAJUogB1aoYmt2x+C9S6
GDCTtFxIWp64wLwkloHmktMvDh0cntpNmZ6TlezM5rbNeqNm5SXEeHAazOLm
bSgo/a1LjzhIHnwdVV/XJIfmGLLzclUihTxvO2CU6TxjVFRr3INmlJyhvcYd
HhGxsXQSPVkd/G3U/n1uEQJ8gLTp8oTOYomgRx5qdv9D5VGl3wk+gisaUGa5
v/XN384idvQnEMgni0ZaYHBSIwP+HXS8tM+eGW8XxMM1/GAknqQA8YwXCClA
NwVGTJUo1kvvJbkDQlb6HyEAwLl/cTNiGyXAOpyfd//+mrxS8sj9cwqY9Rx3
WrX30Rp+S+fLIbmOV5PC7C+D8IRiQP6H3kq9gOQzSSx3a7IRJMhr8GpSAwmr
4t89rkHA0Bo2/2h+p2Mz0TZ8Q3wkQZC8H9kWR55deO4oWvLZ29Z6Oin/JbfW
jSTyZNgEJmO9RAB6wbTSvv/IqhpZybybRjZ1B5OvjKbtAPAU7xa7qe8rlt3/
kTE9N7f63SuARNOhLmutm9qv+HtFzon4cSwgrKFFe+1SUFk6oDudxg01j8ST
I8NxIcO5QsRRZd0qnvZVR6AadIq7jFIh/yshVjqQ5Qe/K0BwyHFvjVBhqjim
tvkCihDOyw1iT33pvT+XVPFMyEb7gC7IzdhAOxMApDtSjbtKPAbKAHeJ7Jm4
n6tcPBZmszQZZ57dj2VAQejucZUcb0vDg0ENeo/W7yk5/b2zgn7ufXZGQu7+
ZqyzaqYzcjtikA80XvWSXSR8M8jfsHb75phDp99mepbvCdzeGf90VEljAO4x
Va2ypjsa//sF5R7J3C5TYg6zf+b74IViKEHCXQUZH0fArPRbf380oxm967P7
DQhlyPnb2wpUBIxy7XXPer3DkPgp9gRH0dAWmtYDCcWpjKb4JZYssu85Wx6e
Xm0pHTujXbxagH036JXjWli6wZy7tsKZ4Y/847i8fqrL2RgxaZJoIkyjWMrT
rys2T3dx3RRvlEbWvoJXD8ll1pv0/MYXMwfKaqGn/keYjlTneydhdUjWf3LC
nl2zXSCLz/bz53p7YVzW7TCZkyM9vI/JgK15kQxdIidWgkT1ZsXXIT1AFUMn
qpwMEiOSwtbPPMvRXRDTHgeKm+axREYBj9ksomYI0+T9fD7xF10usrQQUZCy
MTqSdcDdzQAQT0/GS1Tesf4FBTwVppDFHO2iohbd/FL9e3ASKGaMd3ZiYmcq
rT7kN1XYrNb4UwIxp7OdiGBwEqj/RpnKj5QAQTKqtalgrCtaJ/7ZIKpDa5jh
7vkjQgKa6tOBcsYqkzNfK+U0lrJWIM87qKrLTx7v4KUBKUdIYlKyQ6RPMliJ
/MeXVT+3wQn7loGvp4fTDRiZj0oAUseUXukgZ+8zOdE9gi3nk8x7irBhNbxc
HtFma1PjltV037SJOQeCSFAKZ4gkcc7hU9lGI9iWqTYwJRRskqpR66mrJt1f
YkEYhUjsTFNUnOopIwaYtDj7Dr0B3aFjkZztnB9TBSYPG9r9PJKsOPaknsCt
uLcql1gq7pjVeThu5rDqeO6ukTGvDPA0YIIjOBbZOqfl8YfwQZSkWSoY5l+U
E9jR7V9JHGr6h1s0mnwhI1NUc13/RtXANkNpiOl2uKQKVLicKJ2Yv/W8gJB6
T8nsJVqIuU8d/dSLs8eEAbcabUXheH83vzb/BvFdgoipqdMCcqGNuseriP4H
+5DuEtqpKXuSt+1DgdV2N9eior3wofv2w+roUN2ZhMFam1y+WFuQrG5UAjHY
FL4Zkk14VwUrapjXW23xbj2ceoLg1mn31+E8rvCyf7JgF5M2roXjFqDHOgba
E45yokMHcQnRxgOmMYTTcu1uqQWM+Go2v1qgyuzdqC1IEz5XCmEZtSEVtOhe
LRJBUo89cFwcp7FMf0EDuTIgKsDlgEldpbY3mF0kScQDSHynoYmOATiHXpJN
enHH8r3EHQxGvDJyjsJg+/wM9np/dYwl//S3xpBf1ZpKMZqP624DUOAHxC3X
3EN60/ZsYj/D9E1mTUZ0tenAGK0K4p5zhtOEouO1LdAdhVVgzhoyf8ZdXm0n
QM29hhv1i6uFaqbrZ+j49ppzWNJpTV5pYHRiXhXlNlKN8MXnpxt7HMhfmwC1
OvYEYwqlsfHP7AJiL7vdY0banYPiWFSxU4leuMsn9Wrpt0tldXKP7hKBXAi8
K7k+EpdL375L+oCnSlryGvWWHkbKCPxElVS+x/lae2d7KysePUE56223GzLy
W6g3GW9SJzRzXmTX9qdNcpjqvLyOG7Ly9V21SQSJ85vtpUG5X8VyweViFKH8
oS4HxuZzGktzGddmhEXSv9L9P5XwXRRedBk/fYRtwaYt8sDMcpKwVSCYjzg8
0N58x+RqbkR/NZ0l80Fn3p5vhUuZcZ/JOp4eKZDoyyHN1N8RM7PiQNQvYl34
NQ1/DHYwOgW4N+VZihb94G4XkRl3kTUFMVJqabvjDFnhcQzjjo1sWuu879qd
tTQ3y485Hxmf0hC+pi8vba1hvfJeqJK4MZMzmKd/zArYUKpPsb6m+7gXtJKA
o24rSBpCww0c9o87mvU7U2BtrCf6vwb8xJWolygqh62OcJV8ajH4ZnhDtNTW
FmEjOiM+Z3v5iDLi63/yHSRsys1QGr5IKG2TlllyKYjMLMb1vlvhFPyeD+hn
FcwY1xNID0ABgJ6q7eS5HGYjwQ9ILGgmexhKvYI/WT3VHuWasRh4aV7gczES
Xeb6WLXox7hXmXwYXsbrk7Q8xJwFPhbOQCmE83Qk/bqXG38ryLnyYIt+NHH2
+MPC0m5m6tytVGbIdxiHSLHel9zP8DNG840HSkRH1Di7GbZFlHSiAfZ2lsZ1
E2wpYtnnqDhd7rMH5r/L85Sxld8uxmUtkUy4uC03B2KvTe/BgSM6isz5aKZx
IbktzFhC9HXbS51FvMYdUVZ1KJVoO/Axt7XR+rABTxbn7BWsN5c3FGUPGVSf
Pm0NQFjC5T5eRImas+lEuZfaqqrleKAY89HUjeiCJtAi1PWLQusEJaiMfT9e
nBoZxn3FdFkxuIpMKMsEQ8KCfNkD4YyXxuy0u21UHZIDGCvvldCzQCgJ4jxb
w+qxWLI6EUZcN/mWYGA3etiSPcXhyrS2raIKH47VwkTooVxOJ5JTbQvFf2KG
cRXEUhghMEN5DlS6rgL2XkqrC9zDGuBemLnXMRp03EJb9DmkMtg487H80ctH
AvQoBGJyGQq10VyWEWGPeK7r3DAxxn8lRjqnrs/yd9mtn6/u0M6yRlUORNq3
j8mxfd8IFt+h4goV90pGUyGj2GukzMa8mfX1+0U1JaMp+S/CWxtaNZKDdeEr
vUelHoeBEzDz+jOQDsPObIiWCqV83W310ZmaH+R+Fff6p/o9eAr06+rmySBK
IxeSWlIrVqdkqI4dDtb0nWGL2NV/RWYHpde77yZZLoL0TaWLzQAQablgsdYn
tv2bHbBkv5JliKk/8tfFamH0O3jKhYbd+YKdK6GyxXv72lCYagBu3HMU3rXN
7rGvEkIlRhRD+/Qf6JOT7OkkxhofvAErd6h27w2KLktejJWtpOWYdxwBdXU9
XsiZSw4SvRJp7bypq9zFncOfzO3wHKh4Tp0dEi98zs7NvrnRBZ14DDr6mudY
DKiokRpLqif7Giaa3x8EZsW+bxubumPzyVqsupdKuxt8WvLoEbkrBOy9Z3EW
xs80unxx6Jb4S0dfYxzCjQxQDQc53QXm+FsvFSZ1JEFDInlAIVO0DbC7X3cC
nJALyVOIGfQ38kim/jJELuEbVuc3r5unrJtLLEd5O2de3fF0mBMv2R+VZTT2
hRw2Hu5cdFx9+6rsXi/Dw7DMgcKBXLc0yNcHEpuZ9HdCbLz9x67Zx/eUbNka
xFBFpc+RBH07bUeU3GRxodO+n3rq+vR9lXEt3EUkzAE7+kLK/Sx/aZF2yTXB
KA17XBH243NPOz0FECOHJ9bWuT9rx++npeMiCQBL0NknHAV5scMStOjOGtYO
aFn+mwQLlEYEzWARYfwLCVvtvdkkpZQ1FZnxBEEblmMNZeAaWIXmRnfBvwje
wF6knNPAAqOuwOemRFJSldngAF4aaaS0/bJHf16uimLqmqhJ1u8AbzjvozMr
qJDg+8J762i1I1x36NHLDHdsM/vTFDJqZgCsS9v3uRioeAsdDIRKBX2gVyqc
s1GkaN1L+dQoguygQNbAIyuV6sU94vns27vx0eWn0mv0KiSvLXki5pwH6VgU
GAeOeStorZhkLQK9ajT0Tb8EZFoR6U6HpZM2bvGuAxtVTMYskyg1mZuHaruV
RqZqw/AQ9GLncE4RfAGcAD4hRC4UJliP2Si2xw7hpfS8iz5ecnEppT80dMlx
ShIRo+EzJzqozbusR74gcbV6WtYcs1zX6rztI/B4YBS0QZgkPM51DX6Rdxxg
pwxafxz1eCoMRyPXJtUueT2VtG1GMAdS3+/Vh9g8OAm41skPyEDaQVXOu66h
RGFKMGHMFKTWTK6fmaRH95gKGsefRsBPJdfENYQ1F0ODT8xV5bcCT+rym/BZ
akMb+sr4aHYxDlmTEyjm5QRVX7ezawVktkE+WQFNIB89sF9kJfeHKixXOwt0
MBgdcNl+dB0CwSDjfpqfUvuMK9zo8dJnzJ8BSF7m0N/DSE7ahpxGZnAf05uN
EEtv21pkHiHgEsTzvspJYoNlYWCW15QJYxZ6k7O73EQyuI4t0/nUOBhWN1tU
NAagmt8BPixuLTa1vPYghYdWnFNk2ZOjwPFmP3iLgg1IkuQhoum3+Lc3niLZ
quqtMoPwZNVymc1Ft+UNKy0HD/W4xL+dLgF4kV4NeNYSPLObfBbBElthEX1o
veaM5O7S7pfbVqNfjVQBojlwehOcLNdCLd0xcpx/Y+T8VteFnPDP8A6qc3bW
s+6XS0HJJRMK8P2KvcehQVLjOcgGW5JtKggGhl6Nq8PAKi7wyvC8fHNk5N8b
X4fHGbP71eA3bIyFI1ASnAMV2pgfyua6GABxgBvrCl4L3rVmW7c+Sh6PtlLE
jzq/7zzPCX+EOeGQs1Ziox10KqpNfNDAkb2HTcKk04wbaZXv4O4bck9gcOpj
0w6sq2arzPwZr9bLF7m8CKEpThb5QLI3otYsKVEb0v65XaK6MFfKrl7dShiK
4Q8CFRXoqOxTgvC0GdgiKhwTY5tnB/0V8xuOUlXZjis4Y9lkav2DgEJbaOGf
lEJXAAzu8Av2KvYVZSNxskzO9Se44bLayObcq2ohCxm3BhBIqFIfOry1+m6Z
glZYobnwlfcVGzvnJ4i1mCGYbievs/Wq+pbpHG86QCyOdDv6igM2LDbBxbqa
z9QcVhoyfyy2D3zRFp9bZf9QKtmXo12GjT862Kb4Bx91a4zIpe1NG53o56aG
U0FQ0fL1tir/S3JdODuj+DnFMy9lLpO/G8cvMOI/Dolgtd8MCnRpO4oe6FyK
zWZz1Zwf+8Aapva8+kud0DP0oFA1CCwaubBWkZbzjkYmfoAgwvpf5d520nzB
n9HjpBHGVLoNBfp5FES3A46uzQFDijvDhnZSEp3RyE5S3S3fD9D9PIijFdP2
Qfu+nqcg6dTMUM+E4VUfVcsCONw79RzOuRDLc1obW11vyy/4JMGZMnrpd/bQ
QNJjwGzDBE+94hDNLHnawULab1UvIwVzY7E5mQPrSiWkbf5wef9vOCs/7Xi6
R9YMEDN04o6xzP6U3sqXCT23rz1g8YmtWNOzLHnCZiOx3QIpANThmnmDl1ub
Y0n5ivWlP/yI0tZOvMGiZPn96ZwOusvFOANO65OKPsY1NjvSR4kvddagHQNJ
EShRBHcR4CM0PInaHZbVuJf/LuDssUGZzqgcNPWF+My7mfx0SBalMitayhyj
q+SS32UV0ZtoAC+pG7IDJdG7R+w8x9pJGrZ56sTLEOPCtmFMDhG99Lg9Ozm8
7GoUUODKNK1YY2hL+II6h9VEoD8q2bfxog0R0HhM7SPi43YCxORU9jTqm5Re
IOOi8mrAO81xeTIbqtBL1xZZatm67lfctJHRUjR0wUTFcxfS/AHTwW53QHJA
RijXBnSQ+bIe4NCMFYZxa8St+Scy2JsU00y9D11j3++WCDbhS3zcix4UsO7U
XeNzXqcLlLkb1FPZnsE5O5PZEFaMY3SiEsBsrQreLuyzoHzzjHYEB6n7m/ps
bVTcA1Ab6oBE0RZldxdEVGgyEWMgZjKEkTLVHTwWPknv40VdGCcIO5AjV1Wm
crcBeWjYp7zp2G1esAT+XqP0H1LFjbAYBMZ3SpbGrjYkx8O7tOEQT2HI+g3I
mYucsANuAYvTbIJ+bNYF9+GyyXE3lWj/Hbkg9CHNjDuL3qq5TEPLSnvo8f5J
tfSotRgz86quzEHgYYZLpOfSJUze6Q6yr8YUK8WOU19Ppf7eu6ZZtJ7KB4Fz
g2FcsDqvxQcDGJDweOG4qSSheehM3j2iRodiS3fQtwXJII05cun+S7SniyPE
0ijbbWUiISSzzAkpwBO0hWEaiAdaIx8Mvz6OZqgCBEkLpgovUID3mL4rfLeb
fmrRP74xLuOFj2p/E7gvPrjKDUBeXvOUYLYo0sDznqQEYYsnEEy3ElfWQVOX
W9Ot/VaitPGPgFpGKnehugboOLVXN3JXJFkghHg78JpTCt4fu8mBmqObPmru
1Ap1WecLGQahwjSvPuLsl/qfDd/1P52i8+a++Zy/Yf+mcMK3lKoM6MeBZA3v
Je8pFNHxp00Q5M8r63EphYbepT7/o55dj3RBA8TFbCIOEUYrup73vQmUrL8g
LaBr0lmKyx7IGa2lMuIf1sWtEqhT75D7yNvSxlsbCQ2DL/5/0cg6ADrLW04J
EB1i2oEJWVX8KecRyzQE5Oz2vygiL7BrxYGZWF3KOvGYS8yS7XgvFFVMv0sb
79Sw7cqqpYV5HRcVTuAAIlYJIEa5cWRjvCovp+xFCb9BAkkU80PDUIu4jL7P
QJ5ZFzGfdO4mOjWygqwuAm92uHdReCYiSWQ0OTAQojJOkkYY2JWhF+z7byq8
R91QG+mMLd3tMDYBCWTkQogFG0Zx3LxjWgv0jnpE0JUa7Wb53lMETcQvPu2H
Z2uUhOcu3ISpVMLwsHisMS/LJSgW6t6/PDTrSBLIldwvQ7D0/Ar5Nrq2EC2R
r+4MYdaQ7u54u5mTpAxfcO7UJROP+T1zl3Z0wbDxq0UvxM18gFW6FSfrGTtA
nvqpHFI7LuhJBO/S5iZ3haKaLrQFi6L9sHFPsiZx5uebq+rEUAb8w6/f8qP/
00mjSOgLuTyVgKGQrPJGlkpTXSSd3sV4YKwBgOWU6HwzlPyqfN70U/Of3Jgj
zTTAbiYxlLKwa1IoNOT8pC8K2o74MeE+YEC6H9x77+rnjNNEMERmYwVWT9JL
dbyr7TIW2lfhnphpeP1WrHO1KJKfth4grOlkMKuBp5WGP4BoPdtb2ikWMqJY
D5hw0yDF0zy5FCI5ecHDauoFbFLnwAXQOffL83mlD25sG4h84JmIfi7p3AIR
OL2O2sfH5nkQZBj12wHiBPmEDkwEK/q+R/keNUtQmroW4IYBgsQRFPZYRddZ
0LjYQnZioTm8sRG4rSae+D/7B6w4NPELa1bdiVUoGR0g9c98srWu4OiEOSUc
EvXYdK2Ir8r95jZ2vDZYgr/UQxSnQQy97F5Re2aRmQNOxwggypoo3TM/qN/m
4bzbsx2sCzfevO9+UrCHyzy2dEIDiEU/r8NyIrbJg8wowkWtO/5Iaa4uy5I6
EofWzQ/CkbPKXJ8Q1jt7QufEglJV2qlfDYxjBaqej38nz7KID+SKW16nRuSf
I/na61lfWWeepgybl0o940bhjZgjX8jP77VU5/KNYcGz3SlkTdVySc8H2qF5
KOPm/cULSMetlthLcBWsD4Lcz77tKqsZZEDptizFaYbC0ChOdyOKrq2JKqQX
GXEbnmyeCIjeYIF06ZIlzh3ucmZQE/07CNY71U8AuHs70g9kJ1WyH6TP6Hr6
FXRoMjDt7d/Gt+pjEDvjet2lvn0/SfkMVCqF5Ommlfe/eDyfJl7sIqV55poD
o5nUBAIF/x6+on0r7xcCg+AjZE/WUds23kTHnO+GZq6z8XUCVlC42c15vSMP
xcsiXFMoj30G9VlgNAk8p7JYdqLqIZ39uD4t8O5+WMctP1pSLHYJqbZP3jHl
3S9ON7nWQNmIeKqJa4WPb/k/+HEIQRhiRO3S1MIRnsG+s+3FgwkQ46qL020R
YvpZY9qVkHcoVL/xYczvTzVwaNzYeIWxlvqKZqhIA27lj48t5yys4XPV86hv
z6Yb2lvQP2ZVUHH/JpsLXDMp1Qb8ra3R+oQ0rGEM0DJ5+lwWDepCb51kFDnP
NU68JC6Fpq6vRUyN2Q17i1eIXhf7x6ZrxvOtboRl6WuQfV62aER6JoB+s1w7
oeNq9MLrXLknjsXUcTtZmuQpYF5M9dmQ0eWuB1G3NM5U9FQZOee+Zd20a9NU
t0PDcgPfnjLOj1+nX2+SRZaGik4LVR1ssD4e5Z4fd0IJZzPLT5xdIV5xQ2e2
3T+f1i1u25xg9twZ83lNFqGFhos9Ml4eeQe/A15+H9AUP6PMbyeQAneGMeX5
y4wNEcL1udvROQf+pvCcPzb8mkduuM4v2tDtm484z4NZpCe6taDBosYOFtNV
DhvxD6mKdA7fG8QAlzCzZcEGNzhYQ2WrZr5e7cnoufLRDK6aQLanrxFT/QaD
k95dL7UOsq4jjzaxGdlokv8keyvG4Nck8QiH5aTDkvuDYBhDeCcgAzhE7j8z
oP4mK+VtYmNgiTDWtMleHgiofPKfG66kSeqklQDNPPeUBHHRcoNhWIeSfsiu
0wenUd4IitwYiaNurCiwd/5yz7AZTv482Cx2mhysVTnd1T5bS4gOh2Lbgn+G
Isw82jJcdavydHgEpyfVT752lrceWDZT+fpq4zBD9bYox13nMuFsd/xR+PHw
l0HWoYO7aLYZbvc2CWQCxyOZ6H6ZTqS3ufIDCqPAhl8YY4Mwrh+QPRHP2qtS
pVAMxw/TZr4kePTiVLmN1DUVbUkUghEv28t82tW6xU4PDNSPMYDYFZGG9FoQ
CAXm1J/XtcnOz7J0+rWwgWmsFJdAJGt372DOrT+bHWS6uAH1aes+iEGutsHx
uRTae5G6jabzGsgvPIC/qkzXnnFuTE2MG0tyCoGFaNn4mmclZIH6Ws/fGW1D
m9vzryGuuWTd5RB3ND76nJGp5+mtk7q7GqZScxMisBxRg0I39OM0EqRBXUYl
rr2MVp+4dMEap1gYxEfMMziKdGKXMxfQOdG2tlc3bmml8bRuwLSADYz4YScW
F4hMThdphptQi+2Ljs/jup95H001DOPMM35EGTxihDVSVuFuV5tXIV3Z2i3u
G52tqRGSw0kQWx7Ki9G3TkZ7idtrVlOck61KpcOa+kRMZn+EPAw2H52ji5+z
rnjfgjU/55/nOUebdmzb9mPZFn2+ISG5d4brlklQ+496+cxaz5wxLPCEtInF
SEpEs+G/0w6L47hYQ3KTKelBviJVppegEX2E4GxddatBOR7Ds+/5FMN4S1Xh
HCsE687Z4AoKBCE2dgQZ0lf26lcAE7ZzgJv/BMElAtpNJg6iQn9w8sdoMAvA
t0nzLSf9AOIgcokbo23qRFdSC2pyfY+N6Nuh7yW9BzSdLkS2zTPseoSi0s6j
YZ0u9RhYkbRN+7GkwollMtcnrTCNMCFTptCcbYy2mEETeD+aBrAGA1USK09R
bBINY2LhBVa7KF0Je1Jau+/mmYYE+0k8IeVyye3vtlJ8nOuQB1jaTi2SyMnb
DpsAt+v86qL6jTVp73eOD3amvkFAacSyEGmqxvOlqU1s3GpPdxJB1rEmece+
Xgdb4aqnKHnVxQnZ7X6k/5VYt2zAAINton2ptYPUW62x1Giau4fZAXbKQOJB
8Yv9BXC+YRUFNgmogcdfkJbdbP8zdudQlBAKViAhsZUJkIAfU9nwQt5mj+UW
2KMcZr14S1e6yh3Nw8kBJ3ixXRXniEvoKwKpx54gEXYsKZwKnPnvdplakgBM
CRxPsqtz/mcTCa0h63rTU4y17PZtaIxoQkXffOVAHmDJPjKnTbzbk/5RZlx0
WnW0bvUhxShbW0hpYm8w1PVoVNgO+hVP12PCzR/CuUe9yt5DmidRj46VVWoB
/gcFuWmEq6p0IrX46prlTYP8e9Lzp6bSabHJ2McnMjJo4AuApIH6fglRFckM
YmgjgcRO0BY3w4j3qIWYwD3mvgB2cGYTm65Ec9Fuey6LXjYs7hkNkvk1Zeae
O9htJNJTkuRBPmaVaxxgp+vhQj7Q+ueAjAcVagTWPi/XMaB/8lO0zOLPDKPt
docFtG3RcZav9ydektzBWmYJqse4Uy1jcjdss4XPNMu2jrLsXFYBLBqdVv31
yfVQdfDQyKf/0iS/V/+fGc00KPsOUDygZubbT2gbLnV31DXvRGhw1TdbuZ9z
vY3/jAYheEBypkU/JTbgVQEDreeNxsmO7OjFXnTqEX4zrmw5v+FxfzaqKGye
kjEi46tN7BO/HMlk8sUbH3W9rSbd9ujRr+GdFPbbHkovdS0GT4C+aNQhxKcP
tPYynyAsCeu/9o6+8SNQudZ05LOEaabTF2pxqKzNatMMPaNMtlQoO22x1Mfh
/GapH3vvuN8jJmnsrZ7PSMh9SVKQoXBz/+JcRUQMHBI5WP7XmM+QDK1/vMnV
vMCXAUBg04NRPl8FoJ2KXRzaSiHr/OQRSEUVmOQwV+335lM+Bam0CwI4Ao0x
+S3jGZZpggpoUhwMNc/jeuSmPHU3rGh5C8uDotPoWVYXu834QHOXPSlENJHW
ciFptRtW8mDauNjUfXBZbs3Ohge6hG2ebHZb4KRWpcyLeDO0RQw7ybMXLBMO
0Hn0Z6UCL/TYNpuD6TXug7pxbT4trCikMKgZouRFyZlxjKZti4dbY+cVNEhI
KyanfgmF2gLJJNpkwdQ875d64893dqrmxjBptzXBr2VvX2aYd2/jd11Zy2h/
BgB6y5TXJo2j323e2CRZs19AIPvIbKyS4r4ItW0idUJELW1+QyoPIGzYjkhe
4hX9LrwiVsLSYC0q4yfs4twqn9y3QyAtIurzReClE1n5vzXK3ZTSCZzSkHxF
sX2q5ECtMMtqitAT+shN1HdNNsPSKMIBk0WNHEJHzfohjyE841vomxBilOZW
jVyj6lE4fOKFPEnWw2BjEmsaBdVZsjYsqolPhaO8RWo4v2tra8f8/slFlkB7
uTGmihMadZur8BQAXSyShHcuFmY/53D6xGpbx/ZLvCJwNsXLByUmhDq2LJNf
Cx2DdeKxBCh0iiSLkaykuWiuThy+3CrxyP0v/pE1wieU0GMPrHcL1Wt2O2gb
qT/8zMT2wP1DNqgDUi25Rngud3BkYwnzrB9jfqGLD5uRDc7IEneYsOtZ30+p
XT731RstpXIDlDneUltojl/5hYtpPrzMNtq6+B5hB/Aq0kJhTMqWux3mBbl8
rJPGdCkMK7YEFSQo/aP9LidNiTvlxuXngsdrF9SfO/Nxq2zPdsfN8OeVGJIc
VjriT2iFYG38T+YvagNm4CaKuUuFvkz3GExrwkMMhIfvXONMStHdCd8p3AV9
d0NFknL15NbF0+EYkU7y0K6/87OxpMFHYa4DYnkMlEGViPBPEdgVTMXMq7cl
6e0mfhLbplRxtLnNIAKFmZC38o4imu4Huv5DJIz1bgew8ihTp0Nmz/PR6EcM
Q3NOx/hPpP6td9zvYlUmCWMZEk7YooDE/YbGmtchKY23zIEtrtPyxgZ90Fbf
w2FlEvSwWF6q/ePWVf0VY5OGt7u2rxHlosvXlgu8K9CHfXNhx5G068dGbXsq
p7LqP5O05ocZUwW4Lo3s9RmoEiD0MEpzDCaT1eW9c1AxYk5g1drWur3jwsYJ
IeR4NrF6crQOC9J220ohj6wv7SmSVaKLOfyhoHMDRDGNDTUUOoyrBV8s0tXO
VHL1mjm0x9P/Irq7115EMoOpgDnhftrTEkAdZCCxZlPOIcZ8RQdvZy9PaSdq
Lq73KdF0qhveXDneIVnaFn8i2nvHrAxfG9SLGD3oyO5wxI3kWt40V3TAUvEX
i9pcOGvXcSlmpw5pktsH0PuD9cf1MlaW3XMbtvRXQrFsYNx62Ldqt06hTJ9f
no3MHX0nnQdXdAs9GN8FA5z6fxOQ7boSr04NatXUmJpqGVX1g2VcClvo3VoP
ODxwY9nZItNR042hss1WegLNkIM2Bkr59+kwEwdzq+4rEi8XJxW+ktdJsFeW
EaEUlbuGKeLlloQlBxJFgTdFfHVpZ359IWxEcqDjg0aOuLLmOnf+IrqfdB2F
DkvvGiY1DjaS59WnB9vDFYzeTuh0/NnlvfuTtgy4aqg4g3z7vt1XpZUL3wdY
b0iVNKs6EKTaQJArwu51Fdk1GzOteVo4ci35xOHnXO7nZwF53EXePFML7Ik8
10CkRSTUMrg6LG88LAEfYZxc89NY/cmDwaTFATPX6viN+d5w2+avP0fPJ4KS
B4kXsrDgNnlgaH5AOEa9GWxATLzWXm/CiTk/waK0sWmsulm3PqNk1y+XogWN
46VY9MN62JjN2Oulc0zW3JFQdbs1498tfFN/+tNTfi76R2C2ktbvUR93A0j3
NJmJW1bP/dZxo7elJDhni9FZRuV+CciO5fkObZPlZPAOU7Y7z9RIjictZh42
J0qRWNYtgHVWvnPok0Bpyj3YL90GofiVli3bgAhupytUAbHAModH5giNbKV7
4+RB45+jo9VFQu66XP8ty20Fpv76Jt1078+srwMdQMZ1qO8K7mF8g+5cs+WC
VF4woqPx1z1LfQvhpE60Lx2++X5jP2d82F/vPCs+6NknJqNHlpn8cFs5DLlF
10jB/IxjhsVBsxG8du0QirGc5xGlDhZP7Lw9FOlqbJX/3NzY+ypUf21v2aTc
w9WpiJ3vnWBGkMOjs6q60fonTUh9g1fAklFuQpMtRy8EqmfycVeOXsIYNeZ5
5Miu1qtsmLIdghNN88NVk9Ee1/CDTgvP3CBfH2o4KMHvVl6i6Cm9OydXulsR
U30txgRIUGUdvUnbIBLu1Y0SZtNe63gYGmCcgsnof2bhQNqP7vi4csFUPO9P
vyDjMykBoxNp322t1KAM8xsji2eql83pTOcEfRSx20xNuJOTXV5WRsYHec7F
TIdWp7WFJdLCrxULDEIYvPfAGLEa0pjWKPaooiXBsPgOjGGkQAkRF+ym7P58
mQ2LfqOPO7kMUmX9inobtg+zwo2q9Nu2FlgoFvw/Pdc3ojQ2pmbGowPUg9gd
TcnmFdCntIcXx81ysWFQMbbdqZX4XgNZee2NRQ7fEeDGnOCVZ0Q1k91Wj3vW
M8PaubAnOW59wI/sYN9Rj/xEJJ11OTpPevBmF0UeI8/oW5dPws8GMobpWLDE
e++CyWUxmHh5aSfL0tJ0wZLpcWIwRgYjJoiAPSOIJL3lU1sx2KCiGdfXa5jO
LH8uych5S/+8WRtFllegEXJcqTpFQH3qrM0oQDVVkT9JKbPlW1IEHSEApDoW
psHJ4hOldIZTWK7dk+dpjKIkiW5zNWuArrAuiGJZP6hilszkO1juKW6EO11d
mdchPmmrCaOez8GNR1JvNFjNtQSnhx2U2gKCpQYPgVd1De5hLI7L1kghyp7+
B6pmUNqRY2DvRdHEp69lP8pyyh4CrpwlUFInLNQSt0pYhl88vRo2LpJQVOSy
KpQvYaLP36Vzn6FMkTHMkw5P/Qnsc2aiP1BnwA5c4xAxTrro4qN7c0W0FzMg
e4V5L6ovH6fEEhS/xjSQn5o0APWgTq+HgF2covrEXlyZT+U0aJeGiD2ZEJRD
Kb9U+vMsFRGA6IiT3PBjJ8GYgloAdHv6bmDYupNkpu/wM1ns9VnlLgPdCpmd
0xtUU8l//qN8bcU4mUlTks9yaJlLXrx8mPRC3jHam0AvOO5ODcw+ilLli//R
kM2HQGdNa8IKQ6xePM7QhaBWEEfH+iMccTwtBFX/FBNVvJBNMXZ9gEFdHP+Q
MK3d4WPMAn3nuTLLdKbub0v7vtWqMwdWbYb/KSkmlVCRSImNPM+maXn/vHxI
tqPmCQJUEwYR0j4Onp6jFHSPXkgrFbhfdhsnXUxLn+CriYAiwyxy93dUfJbY
GlrlNBGoPJr7oDn8fialVaMJLkxwm/fBi1oqR/lkHQP6lcmfn8b5aOfXzMzt
GBa2x0WbuJnvYZpuY+fS42Kky/RAdX3gDFBfqLa2Lf26vZDg1EfktACtdy5f
M/eL0nQZaFBbvgynS1KmWPax7dv/bUS6pz+i1rqfECf7lhl5/cS5e0DIBz+d
zZQaNeNBx3qUYg1L8ncBu+8MDb151HMOMlGzqBrFzyj5KAUJmnIpSzlTKhVV
R/e4A/5bFb1EmS9tzPE5VxwMmRaDFK8m5NHhJzS/UOM0YaGatmR/nrq1YSda
a1pH+YnS/9bxRRVQFAiBogixcQ35IUde+ryfhhWFy7aSXKw15DD0t/eCtvC9
lS4KuCd6+wUKQA78OavKwndqlDpYnihhoLdINXRHnRD8QQRus/kv0MrOdHQR
B/KT7MU3mbqAmMu22AQyxSmfYIdVKEfw4+Yv/3gAsJGcJdVY2zc7VAG0/gVm
TF+/GHzjYPs+RWRJ3/JMdAmseoKh9mRgWDY01r7BWugybKB1GPkuX8GwGhWy
tiEbbeug3kyJtdQHCbE5D7/5LlL66eUMsItMJs728U5x+zvKiHTVArzs4UIF
YOOtveKT0NGUYLEhdktuA8fWoL4YYVNa5v2PtxVYmUOFtOak8s8o4Qs+G5wi
KRoSsOKaLm/TxLXVIFwV7tpYqOy9pOCT622MOn3vGq6OXSWDn2ZEYZQpfoKS
WW63iT+vEZo07NwZHf6fSujVk+DOK897rtWDt1VBVx70u3bSC5VudUEP1OA4
EyvfHBhuvqZMrpZKQ6rIcey++NOFo4KILrVpwK6IlQIaBbscb+dxkpXJwx44
9KcXrKFuCIl+pIA+noHVG0gEF5TeFW3TICiGVPX7/H4X684QojLr8yhX38XV
Oo1AfgpLDrWhSEgGkuKQW2dl0x0Y+marXYMS3/Q62wlito602x7afMWzSfeQ
cAzpMJajuNkmngBI8oXPzqm2dhc0xQgPQPgmVLxF0aCfSFLobxbYHK4jQjt4
8/fmImkEkBlhPX7niLwTGpJ3038gb3dW2yxYHQxhqL0NQYwX8c/UQbN+qysR
8sCZJjaFN3rIb3FpUZKODMfmxUu9/qvB8AUZZ+6FPzmurDR5XRl/oFFX/aTe
gPQh6lnURrTQd66Cm3Vg1ITJZl+oGYpC33z3NdFdzmbU2Croi4bbWai7g847
FQjSpjYDFSJZKJrM4TXmTyhdzffRoRP+YW1bnzEgDjg/jPRo/cwcH4sqkxET
BQ2injUMlTIiw/SgXyyLpGlWIFbf4OhDdOTc0g31VLpk60nMnrzBrRsGfEbs
j/j1U0lJ7ag3HX3tK3UiS6YXJzynAcUrHZTN3o9mpwhHOuIkElYOzrS/Lsnw
cUji5Jna/csTgHoIl4/t4pS7NXel8jZ6DAVYv48w7oO6J5mevqP0kIF8RofC
sf2zexKlyVb7cr2PAulAJMLE5d0w7hBjbOgW+okaTBnwa6rSeZfVgGFDjQ9o
cK9Qd5wCvU5StjCzQ0TggKt2weimozeUIzJJWwfFNDTZoo9IbPlWK3sh/unQ
r3cG5X25Hy18jvoLLMyV6Ao/wdcnFlBLsP/UpKMwk8S8qBmJffei6J9aow5v
s1NKZ/x1AQ4F2z0F4lF3bu1aAm9+k+NtHQaD5sKnlWW37TbvCnssaKguTFEg
ORPWC3DfULUYCtQj29vttreTR9yUUDHin9zf8LITF+SxTH3YwiOypjngUKt+
QYH0SeFnH4gQwktCYN291p75zN/fb2s5O52q8Yn7PnhcUFcbSEB9ApNj6/Mu
XPv3nkFlLCMIVAc4i/KZiQ8KuFT5fdEgC83VQI61s25nwTkmmfpLLaiR/Xg3
ZLW3uJqqUWSV3D0hE3BMThz0DPXo1r+wG4cmEXmsFvYstzn4wbth42aPsUKS
OCRrxDyg89TqfBWFiImDMoFsX2Oh2EzLQSt4HauzxIQxFmQ6UjDyouVypecz
2B3Vb8gZ15NRmDmGNKqXY/3qCqq3iNAkvwY4WPgW43kZZuvr5Tn+tWfCq7MQ
f7AN/CVVMiJHv2qoi13ahOVHeXz5aEFNXNOuceqxqKE8TWK+g9BhuJkZGsvY
K0stCRjzSR2KiYESY1dvFXwgLScC563EVOcm3NCt6wBPUhwEgBH/c0SPaktd
zgnmnYyHwhHR1uM0m1aK4KFRz6D5/AjLdY+whvtgzBA5rMsIoLtGie5Q+B+7
ufpygIruDygU1+BLwiRzJbxCa1n+Tfr3Uu/6ifbB1NSowWUCBc5JFC4NZ/eR
Ozxi4GqvaRlNEsMIkBcarB6maXzrdhLEHBySGEDq3qvt4Q8kgydPRM9M+ocW
E8Ur+mpceSSeTA6q8QPWXZLXeIdrO6fTJQ+QKuLjwxN5Odt+7kv6sYyklCn0
CTVLu+C8wx/2+KD3GPOnh0TbFSGDzbjXJTIMcBY4CT0XZQUyG3GlKDySforY
FPz5X5FsNpQSc6kq39HLVGeW04U1wTrqNM0QV30zIY+ZW4Rkhzo56WMOd/Jr
tQoJdCBnduCjdoUEtzgfwgppqaHMs9kLUIiov1WBhnSNnAOr+/WcEFwPM7ye
4rPhpWVB+E1r16EJMBCd9nM7hkcrBxl0G6a0LxOiGAel1B7A8i4HpwQS3yPa
rAatq6lRqzYghGzxADLZtEWcbUoV0afoObVYZoJUA2nTbAoZxp0/3V9OwZDv
QvCAhnPnFs+oJx7gxE7vwztUTsrifsXJrkuX3S8IqvtzMXfiO7ygeR6zc/GY
f1+MHyoqDukjSrtLA70rpTegRcYOg51D93/NRIGlH301bo3hyE2VCl2exaYa
4KX1zsU+9HG4eqWlDtUQ7QMHfUD0wy0xAoqLeq4u1FXHC48YeFrSIr6ZuGe+
kAbiAWT+5lu7JnQJHi9vNBrdZi5LWNp29ipXL+7XWPDkZ5RSNvsj1VDX8yTS
Bm8X/KrBMGn6vv1I3S2VDxa7N3u0AdSYHvUHYnxGQMBTmWOlt1HoZmf4giVJ
aj3IiXGk1LVgpX4F2m67/HpNopc/bUWnN2UxIyYOLx6M6o4mk9+TlOfj8mQs
kc+Zwr/LVRr1QC8TmM4b+fW/nA7vRz96o+KSYby9odJgYajz5tP3zNzkcBeB
0HA0ovTRtj6Je9gSaL5Vj/EvCwkg1tjctNgts00GFyZ46QTAQDE/MEtIxRO3
W0tUsvnVpsP1ZCMWz4is+FwM04ohaFvYRNjdk70Hh+xJvEOzBDrwMsc6ThtZ
T4eIqsOyVtQ0LevouPT12JHMud0F8RopWK3REDYtn8DWXdBseFZs5ZLy7h6X
JJuwJLpx/9ICP1iYXtVRWXuW9JmBDXynFn/IHxZKgrvMIGAz/iXMr6lVHbkI
HIsagoveUpPbV+VYzu2PwVxyS5k8r3fAdLwYkLcVG/vkP/5yy0aQtR0sV8tX
SZ8kcw7vsYNvKk51PekzBgn3fJLsOKxI3u47g833yG9jvHiBm2FhzEpCwbJG
9bimLuwGMSdDubR6XE9D7PORnRlEHw7HDkB4uvoO/4R6tZCD2LqumVX2ysVC
I0rzPCGoN3xxpYqygv2ps4opveet99rK7rSAIqhosKwKxPY26bSIyXA6sNbK
UbXLuLA7lwnFq9k6+kN9+2nHBFMWZ1ZjyUnZcWfm9ZwtNWdIUiNreJSun0zX
uyxOW8Dr8hwkIgd2Mpb/mK4aR+6Lc75Txwd6GKxg0ee5SKCle3b3rXFxHrl9
Tkm4ui+ybKaEUl9Hy7bTibmgg4+CY98YkjS+UYr1s0dQwIxQobuyNvYMtX4r
v61bWJ0U3zXu31lUPCeYVefshgZg4Jmb8LL2kAPYIJnKqkQRnJisL5HsOpap
wcH2gqdPT8n85NOabgs4+g+5xVXYioClnoOxGACFvxShzSRnOqJcmRM6/Oo7
Q/BNKioLhUARtDB2obOxAiI7y0qMh79NF77JnJaZBxJ6PqTYuzEa3oFc2H+9
cbWKlClVPqeaUGxJ7QZM7R0/UkPnP5tRW6Jn3nTw2wS6ejM37bKnOkT4z28E
kH41tALPG4M4ShUMvwdDLBVEZfYe5CrndczrXaRWYckOMGB4OLgbvVeFYLZo
BdwtCW28cNEMC01mpB03hJYNaXjF/2j7Urkx5aRG+gVP5ZoBDjhYiZH8P230
QbFpEdZBwMFfh1RIM9RR/KKah3cp02BGMuV7qpAtEqL2CE/pP0xTD6nzvOS7
nHQ2s9IEMQqZ/3YTPb5xrkBA38jspGwsldI0cZAhNCl3/WRM0mMVT/PI+NH5
TIx6DCd+YTC5Q6oZX2A8bwLRevzOdI5R6iVv4Fd6FXKIHVwwKyrVDIEgw9N1
YL9NvlOdqSLZPqqxT0Q4YRUqmSyHI9l5QJkLj6ZxGRzgOK9Uik2KbwiW0eOw
cbEiTBlODOsLPd+3FYsy2YIX48dszY1aYLZlFteOGXJFlYkzuX6g5YiDe/jm
DxK74Af9qsyp6CFYoM+2PotZ2J2Oj4enVx5stt8oJaAUxZ+LwHwkS0ojp7nH
HySV5zR1OVWtiqTk7Z3gUNZFeAzOG6WMI4qwkacTthNFLT0+xHn0gfeTmfRg
eEhQDiDAKTg0RKCd/4riKS+lZgk+YDPEDCjUqdo3awMedNWYzP3sN8UsLLpI
N6zniUsIiLMWtkwrR9PIj1vetZSMrr7cmE+gPeZWOAAqiDwBFLU7zV0ywfGy
/8wkeQ8TuE+L0o7qlFyYRqRq5QwX46lY/FhOorAiuehktvMfOqkNtEubQakR
eMV/s8mnu5FPnnXDyUYo84fyLXWxu4hxYWMZv5fmXoMsup9Du+/x4SYLfAC9
VzLP/TgMIHrDLbObezLTIma5EdcKH18nDyML4fL7H0jDYxE/YhldSVi2+YQm
3bGP7wM5Yc8n0QsTg3CHDzosMqDO0B8FD7hnoylMaxGjWZNFQlbyE2dlLGMg
KaMChgZoBZCcIV2dIt7rZWqHF3XxUqJ4/6nasHvxud/7fDeAV4yNWJyEVc+x
zOv6RMFbH7gIzc4e7mcFztq2M0cGMzlJWFufqRwQxmPOC3O967+fWuLZDi7I
pPxu4K2NKxGghe3mjFB0eks6jyWjgIvFGRfoq8YD1lb0U1ZXAYsRytPs5AsH
5BhZZQ58e7XasnxXtYQnlDHAnlCtdoGsRHJuu+JP9z2XDcjEbNAM5HFvHRij
CLzRbwps9kNxHJjMfLqBezQFi17m2xm9XGLf6NiVHyNrNPKOaMLppo90yS2R
LSTEXaYR99trU5Aq9U9iOUExCewZw/DlMqwxkfWs2rk1uPOS9hxsgnCx3UKD
PQqlUHiep4uObGXjgMJmU/3aDBWQq5Ecxv8l0ExpjcSLrq768RxAXOj5UxVc
aWluJNAj9yetcft2s6PsbcrLE6WkyG+T0XOyTnkOS3/QXrmaMWVTcXG52eOp
a6wdIQ8iQECqwIJOYLB+7Sdm3lqP9TOgsKi+wnZPmXCPQbbpk1oWNuFfiwCm
zlqxcsHjAxcyJcCzLY6fVwCkMmycMQcFvDA+uE+pxLMef6V2JCg2mKLEfNMA
XXtGaUFRIAw1aPdDvwYqMqsprO8QCl5+8jB4oox/Ous9O2TNDRTmxPdmeP7l
J0UtKpGp3Z6xNOTy9dMazVA6pmBJ8Opej0y6cAe6lz4fZm/6+ZN4VNPcUBbm
m0cpM35yrcWIjeII2PxRjqKAOQef90f74Vwe6zD2oIDJcCDdZBw6IDbJpWbb
WcIjPGFnIIVcf1xXHxFCzobnCMhs4V4gkAIzW96J+6/ejP1Jnpur7treR+q4
sIVGnNMC+vi+1Dy8gX0Lb+rMxUHLxyzGAKmjCK7aHN6aiGbs2vujArHRxBIo
0twz43/N/WHFu/uc2fZes6w4b/iu1HUxvVVmrO/Gr+OXzlpS9rOVqLFb32WY
TeLfmBO3SKWjGe7OoBL+XNZijtjj5IDFgH24bllJG+lSVyI7sVLuIVchVDQs
GZztxKyNdq3pxXt/XFS8gMJ9IR1qcj2sbXIBJLjJo/e4n0a5IZ1aK0QS5/cM
jFFLAyNqTW5uMsj3ld0f4sNr+I/mrB2T3PsnFiRsxWBr4bJVj4Krjxhm2OzW
VuXHra+pjjofanf1RDdySoGg73AkWj88pmecjziLp/qOKOEIZBrXGm2QjNDn
HDl6Z6Amwmu7pnFfibMCREpdMPm1MVVYSdf4DhhSE1iFPo+rBauBfQMJ7p9d
Ahna+8m8byqz2zQauIVewMTTIz/Q61+tadygbVgZzdAzjkVtdhR1E8a27Q+8
OA/J64s7Rj6AcssDy76ulOQUGjasTj8KZRc3bqM1NUecAbWwBsANVVY4SUPr
Mad5oDrSRXXLyffIeDAMSQVSvBpySZrppdo84dvV8OOyqqMm6cIY2n/JxmhG
DsjO24dSvy3zmZxYMO6WcPilLZamUZAmh8pQKiqvYzJaxL1DslKyXVLxPn9J
OD3GJ6wGKPUvpX7o0VNZhcfIKJgGXUvB8sXgpkwI/XFHqmGjmR3APK8avfpl
690gPuPjMXZ1Iguc6zVFMIdJUFso2OiY5LUzMb13czkzmm4CMm9OvVa2lf1z
PcWojdS/vW6968eO1UEvWtdQG5/OpxG+/lieDIJjSL3MVZPlopiWa4+ZhfgC
0YLbhKiZKrjoE3vdYTvqFBpfkhgOFdP71s5blr0GyuQo+RPlAtiDTVlHz/Gk
v57XyWtLjpXCKQ1D16LV0T0cJpwKFw8nRVBQM6o2Qc7lZQhn0rIyzzdBbO1B
tt5iY1fhNtEKGUJPk034UldFtG/p+bj6iqm2RYiLCmtcYKMdfv7K7rDFONXX
CnUsC1drJ+txYDmhEz+kNAv/BoFH6jSTLuFcCI6Th6RmMMGcjKIUYSRq5G9X
vwg66ryYn0cKecLb79/yQvCsKvTASePdV/RMpsuhCMD7qid+bCKMdn0UCaPi
5lH+TAcnrzxAFg4J8oLJNekEye49fyKVR39Yda3sY1Uf7oHkDMawpU6oqska
z0yOgdQdyadSjBAh2XyKQa8e1DJE4qkER/1oYxHfiZ+L6Nx/vWOuSbFnqBAs
aBIKgC4zYfKGgN2jFf4Hg481mFvwxQhldhylf+/JdrusOElfRDJ4bVjZZjFb
lrFO+hLINZ6Q7ClKv1uml25LDm7IJd5zU+Id7JcXWkMRLzhqWaw/idc90XY7
a7r3+Q6psqyeHhRueV9XgO7ZXjAtmGYhd40+imT9AmdHBFkkOafJKBUfAftL
d0y5PjxZ74iYm+xG+EhLIowrmQjxKR0netHwJ+NiechdbrDEVzB8e/9X1Ozr
6JXFrj5yQq7QZKDekb1plTz9y3Q6FqzEXdZEc1j3creLWZPTeGnJL+bv8WjB
4nRfrVNBwZo58c0oWaA+SHvG77vSowV69McVueeniYL23WhOyOm3yDD3GVK7
IAPw0n2HbirXZl35WemYbmAyfWhyhXh9EBAZbUJcCGhcaXfxatjL1y4WM0XW
xnY9gLIRk9ku55P+jWLpsfWTrkQbe4Z70W38VQZiBRnS2KD0fnQhOH7RyuUs
CrNiHTWbmjl1IWC7+T8uh8Yc6ZQ1WeZQCl5HMp1pTYAXOFtMEpmAAEJYzrx9
ESVSb6Q1o287kdcJkbTpsFuoxoGSvYcEozRRDmU4DuCMSPrlUXi95ZtDumkA
v1FdTAlFjPJtBB+Rq/1ENNsngyeKLQLOYuvVk2+eUvbwk54jMh5JFsMWCIof
R7JyCyzZrVgD28WRhD626FW51uiiSL2Xpg17vfjFEP2QLY/+IbwsqgaMEFyH
yDjMU9Pes5E0EKnqFIJ/bQO0IUfZqBS+o54SBpLbgMIAWLt/aMqbKtIXToFX
wuxnp/aloe0bJrOfrk5tDeYdHdv/ZeUXZETOhv6sqk7wYpwIiKT/VN1oOUk9
cv2O0p9ml4gDQ4dvZePDgGwqWOCIeRsHW38kBWzA+hN8N4ne/xEyNT9A36Lo
uMbo28KiXXYbn/66QeQnAMh6AjzeC4El1E6D4JCEDMU0bO24vvSoytePMiF5
t2busNVAFHAaPTudbQjGjwD+0RSZZoqpq9oVPsVrr/jQb8ET5izOChBk45VV
D4Zn9nEH4XVUnS4Roe42Fmu7PQf0hp/cKq2uHmTeOWGBiHqI6rASXuqD6txZ
/Tox8h6E+BcmNvYGIjUKkYt+b09kMfdNwmfrSbUTdLiRC3ysDlpn1nQK7pnc
vKIqq3b7FQOXrwuI9l77LbWypHeY6cALPBTRxtqO9PVxPlfFqqX+qn0nEwYe
Ew3TqLgA2KwemJvlikoa9c6kuFwugStFllXd2f4DruIgpy9nR8bOGzy5emqX
XQoZG60zerJJWhPi7ZV7AAZ7psDxgcWIw08O/jw0usgrTn241AiQVN0YoHN2
x/9qfR/d66CxVK0IvKpUUFUxjWtpdtRMvmTeSLQ3MjPzbLj9Zb+WBe2PuQp0
R1tv+2AnSgi9qDy9K9Z9h9F6LE5aXxcsfnTE3UIvm8X0U4gSWL5v8FVZnwt7
cjS1YwR9Xp9ey/xpXKBkRnTo/INPl62UJ0H+QDrf37OqxDJ5fjFZt+i1AtNG
CpM5dtcgyY6bhDE22oaBkOzScwx//RJWFaiRQbG7mAL+FqwGI06bT6isAFTx
ClycNv0hl3nqsF/Ftuk5YAO45Pm9ePFzYVESpC+tOPmetvFzp7nNF5iXrPlo
8Wv6TTyGYqOmAquDPqGjYJHejN6tO5bzIGt8QjEICuPy8qI7Nk5NTm7afsSD
k5jLh1/ZHGqpjV5a3eQhtSO1zFcOjbUddPTGoQXAZJsvPdBnyvYIb+20BMUZ
Q6dTynDDrbEweOqBSpghC8qxPYmB6aBOLUHEf1UJW3sQsFslc8jVwliZ8k9q
GajIjCQgYDp5UjXj0oNDS8O0+xUWY/kvd1ZeCQ1CUTpJd6hPtQkInwY+BQkz
D4o1I3MUYUcgFTvRvzy9GatM5+FMz7u/1OQXE5tqy9qYSisRgIsj5IJTv8J/
o1qtOAsAXkszTn/dae8GKqWCOY2eE/Kh9ocJ+75sYPDAVkZuhocbeg18x3fE
MUi+OmBhpHZfCQf3YkeEAgFd5SPS7o3Hc/ieA81b5KIZe8DMEKF1cS1HidVY
ox8mudO+oZpTAXBhEeNZv4xecCPQgLc6sY05z+8VoHxCKfuO96yBmJ19dTI0
B31na/6noAt1pRfjGfOClHPKxFguojIk9lTAlY/BHLUUd92cwzvdfTaxS4JN
Wy0NNHoY9xRQn/nD0HG6y2sDumWIOIIY7t2rLIBLL+/na2osQEFTXeC2sUg9
vbomYBtV4ufsSUEJlvE2VR2o1fdTSZbhLXyvq6Z0dfN7wjLel4lfRStfOO0K
MvWx+NAcZJ8WsA1tkJfAHuUZU3BEyeRFuBnwC+M85Q/dYmF1hIj54TqAWQj0
HJQJGCSsRSHXVYhCeWnnce5WKw+1ZQLq1hVjer49fm8dAiimshCIIWrLqowC
4+Es7jxUm9lPJ1GoHJHX3YjxmlY0vbKbyc0L9x1EiKOTxZIpN5ALOwgQqv8c
P0XLKVduCtVbMpVP8jBUBkjX2Y5fnBO517dXQB0lhrFSBkn1yl7+SxYFv/VP
Fe5Pml7to5SsLb7e1YRurflNPKypE2uqEmKjhUfIni2W7dm0KlrjntKNKkoX
XOZuHrYEs1r8CkrGo7DceLrPnFs3y75kwfvndc0+bUuKqOcJlAsDe/9gzPj5
83ryGsBfAGXjk8zRBxLyVWa9FGuhGKHn2qMgdwSsCazpLckdbtOKOQnkv9lc
6tF+ovKordjlY2UgzwYVDyBSAMYdlCEeG/rqgtIrcR/kC0fWIhffV2vlkFV+
bd176cdpALvBHGeBPF8wlW4z6PYcIlyDSc1KpMTDgC8wi0FscA7FvtjcNGkw
lUtwhztY31Usfi1rpXdAn3APa7Pd4cvO6/en1hJyYXBoj4ez5rWIoT7u2md8
410L23YDy62qWGDOS6p58Xpsq9JwQC/1xrVBx6bj2L2qFd/Z0pGLh0NE+H3e
lSuz7iRWx5Q5Dp30sINOaD9RAvuJF5E2IN6daCj/gmoO6FImbAp/Dr/iOh5V
Ep2EU8F5vOwH17vqPF7DO2ss2C1r+xeC3pYMb6pkeJ/uMkeNliqZyC20MfPV
DGALRvOcSK3uDVbWzLOWJhk3vkMIbHGUgr15c+dNzGop92lK+ka+MIDNNd83
z3NHbN+jxunQcGqboRi9dsM+P+jnujmYUSUh60IjTUAdqBP1CjQcoQVmDWdR
zanhopoVbFDFnevgvB+9fKk/i/gpn/8JX0AB307CZGHWed6VD4m7ePb8wJ+0
jdoloIAzySfJMizHC/JKFya1pRyY5mmNuhZ8mDBbFd645l8e4vDBcKc1aBj/
MmyeC9rCoWCmPqYUCnJ2BwkZNMyOmqRx2IRVZ9h/X9s9Vmhfxtu8EAyqzSxk
/4hK+r0CZNj43ORXaH0bKZZClUdkXBp8WI4AKARVU6PiicnCLhtBwExt6/Xg
kODPVQ2yvCX3B86jrt+xfoI3ezXwMIUmZiIyWO+Noaqj/HImUBWBfH23H+Dr
AWMS+ZPJpzzGDvDdOs0yxpSvD4p07PdKl7smPEMJPwKrCh5hHW3GT2G2/Mwh
7ZVYAX8zipVsD9H4F/WGkyW6ZECNxftqWi6nMvbn9L/r4O9ZAANlp+mHmFlj
FF7nNVCytqkD7z6Y8gLLN4xE3fAOsh4vwE9fsZEnHw4CK8sBHr5hJtwv3VcU
EQvL2w7l++e4+x0nATbQIzUfAS2+jAbwe7njeqbpvI3R5pGIsefDkdToLRvb
wQeM7/Foqt+FYlDIEmRutpT3P/dsgQIqNV3XAW8fCNwobUoUlSed0ZjmC21i
VL060pp1mPeY/W8W3hzoSBMd6aOD/ghN8pGjMudN/0mY2zcmy9hhGqJT9qFz
eidA4ilK/do9rsZxC2K8Kvmf+SudTvalDKr18eNIZXg9h9Ou8GuZZRVNJ76o
1vnrLW9VnN0a4yDemJq2ORPwU2g7MugULnT3UO4Lngrki8bEozLSccMk2kSI
YVfmOyS9kEPFVqMObnapTIWhqwSN15uqvTO9+iIRhpnKxTnT+N+EGwU+DpdY
Ui2oKEoENdMOlgEPF8q1U3VJtJUiEwIeSwNCw9z5KlibrOmbgmb1mF9YwOkC
NSfXbyDpz0nvVbM3u0GQWxgC4iLAuA7BrDH0/f1BzuV5pdun6gE8rhzYtZZI
thkiQiDLyvO1OtPwHAphhTLbghilkQ6RqDLV1PqmNMjt3fngr4eSRSKEOsPs
0NzU4B0RY1IWGk1MYWJBXZlgxReWw+WWNiqa/LplL95Jwdc9wEMjOjVSc/L0
e5ZbzrZf2DRQc+OKN0AA0NvQgK6Ny/G0+rmERpBiltzM4Ee+BagKTQAtC+y+
v95+6oma5lTe/LRr9sk1Kd5qhUHQKs5hkmEOzIvtyGnd4qN0mIo5sUXmxBti
z1AvFdWnPNflk4fEhW88bNRfd/qGi36j6NpCcWmi7UsNB0AIGOn4UyCcr6B3
1Os1cJOqHxylSnXF5nl6SFbB4ejIVPYJSTo5c2MJcCKNaRv5V7Q42sv7iVF8
tBqO53H/D6kAmgsy8BIw8N2d+iRoC5Z9asevIBREOmNBqiMbQO2X+1N+RMVx
PCFa4gGwcpu/4CDODC7oeDnw+QlBxRwZW5kxFWZVY09rxwaHW/uLzL4IdaLw
UPbOJNikbu5JztmxTWNBwL37PIxS852TjsSrdxKzilIcYq9FKpGSHH7vCtJQ
ROpDikrPYOfxuTy7psCJcgsSM3f6GB717c8Y58evHRNGHCjVY9N/rU9touxH
LFn4PuuKg0gyLtc/CbCM/8yvVCML6bXk9lisaj09YdOiwuK27d0XWYBDbpBI
By7dK08vqEnRVb7vFYYfETFaCS5DshgXg3AFmv8IZ5eCCzTmFdwfhc/a9r9T
zJ0P96ozLecfTxPyCkxRdlwLyDfnacjKucwkFNP9hFFxN/99Zdmt/lLVr43H
O2+xXpvPavbL7A79czMkKkKUE08IcH9/tOpZof5zehMrgsNEoA5iKDg47RXK
P9ML/+EIsysryhp+0gdbS+CJAzoFIa2H5bI7BdTPLMznHbr9WYiErrnLth+F
q00Zqb54hNCGZnLYRsAJzkuxz72xbvKKbZfrN/5zC04dJv+KiStYvPkaVjjs
Dr1bkZeNkjdTSLTehbvzal7yGC8OVnurcJOjx6OtfzaQ5N9BVQuYokpsO7zH
YH7z7EZ/Kx9aOBqWV+ER+0t8A9OoIsokw/xhJ1wfBHCWk9FBOUMOiI4yeRy5
iO4uH+l5Pr1x5V9oLqRcESuvOYtxrJVILP8WhGs5hd8n1uRAzdRdSfe61opW
ShQQ4eLW60Ft1BtY9c94Z203fbgbfdJfBN2lee8rBVvQFRGWbJKuKg9fH/tw
9U2k+8MpZ4dRPtnwhyfimjnS44zmDZAwyfFBYNWsS+wL63y5IiIuMnlhlg/y
w8yZ5KfEQhPBPdEaAug2HioJWwqUL4dz+JxyRl5v3nz3pscbMKhfhDwqNhbv
wp8vghoyoldYZCo0JHyyLgpmAxAb4IGVHDwE2+7eEiG+sb7wSmku9WcO4F8C
YJa6wSVtg94i2COAAGza7oNe7G1P0Z7+QBGFigea+cwS2Yif0CuZ4f6dGy7I
t2BOSyTY6FYZDZNXfRETWpNmq0eypThtw+xMuNQzxxDbzW4AH88JGxfc9j2d
LHLtPUQgNeQRPqrRCnrjHJYOV4Ga6UD3aFo/5kGK9GQvTspJVRJ7Grr1pmED
0ePJuC66N4e2HrlQRM07ojeTi2cPnOR9WlT6ldS7NaXkvvrxUbfj/Qx/5/Xg
4sSWKQ5/MeHf8X1H0JojzK2wKr7/HWLzIvr8pSy+0IJevs3BhkIUBqC5CTgH
NyJfv7/L+3HVi5JFb0GwloqlJuYLzPvebCzxbns2Hq60OgZadNHMCUb/uvJr
aP6OxAY03q3304p17t1o0reHSGCPXnMyHOyc7I2ns3OorCxUUEA6047iG5im
k/qQrjTvQm7myKnqZ1dkzrPr2N9+Zgz0BF2g3yvgjJxNM95BCw+6DOszrQXP
OddqAdY3T4gFE1WW8ahcEVu9EXlNk2mVnVKUb6aR1ErZFa892CJ39mJqFQoM
9xOcV4Mf+lelJ9LdLAIR2j+boMXGFSaEuyeRCD0TNzbUPRsDieEeyHCJ6sJC
ondel6XHU6EY2FdL2DrvwvsjId5O51nzVky4vqx323UH+AlD/VuT9S79p6o+
C7Fq4OXMKBec1zFoSMh1ro1mO3iXZUkHDb5yHA2/utIVQAMJLxNsKPqTfrMM
qFAC/KhXVsbf/rASw5doDYT/EAZG85ck3HIzO1HZwBfXPRGaKYAF+e7gi/u5
voDmc8AL3ynOFqqJDQNHLffOGkrPR97qlIjQ/z0jmEGHheWN5uYY6vt8hbBc
VpqGzNeKX8by5shZgfbEjBGAffGHtxhoUEZ9moIdge27RJpq9YQzBXMIpr9l
+zZBL2aBt7QBSmrExRE5+s5hEVqeMpPUCeUSKgXys6ocJEhUZnoWad7ikGxx
dWL5oIn+xsJp9hjsT0PWwQFBXoRMlGtmVcKdvmoxjCQnZ+k1Ri9eqMyoWjVV
yRQVZsTCxbQlC+PaPaMINe2U1vxQc7V+1x/Z64QaCtENa91XJ3Dpc1snL9Me
rpa93Bdh0QfKmnCgEhg5to3jHeIPmM6ZT6TIq/TRYMiQkT0+9XA7evV4Hop9
/FZKttULPvIFpVFxGRFbI88kYxX0/lU+JhsvQeB9OgscGQ/8BkD651ts9EGe
WH2QzQcdl6yLPhk8Hf8w/Y5DhFMoVXvN18Myatc367LpISwU9Ly3Wo+CKSL/
p1aTtSn5zLeYoHFNstMV1HtytJRYMWci4ss77d8kH1haqmke6hCaxdaDGPFF
G1M4m9UzUtjVwRqY0YAnNX4Hy2vIdDxRYmV9Pm4V5weiZmhjZY+l9x867jlG
0yQ6jjbp26Wr50LwUKjaG7lkSrJpL5u6NTL9gunXY2qF2DHQu4GXF4AEMVs3
iFqu/D5QfLKZ4R39zbe2sSuhr/8UUH2kEVVBv6CM6as5fZnFEmw6ZeAgUvAe
UlLanC+l0qWbuai2nYPliCBlO6BfS2V7HT1cu35TemZBj6s7oXtNTl2dp7Ns
OJRtrl/YzpGD5yppyOt28eSBoF+xd6nEMl04vVi0UbJ1z+LmuSWbM+kCQAQd
SFr0Ts/jKQCyJo5TDqZzBhbwzSfkSXYQSwP7ESxm76tbLGxOobhzmNxxAvUx
hZxFgNKeJGdj0oE1U9FWB5SbFIE2dfDvhKTt8uvQxIWVElWfrF67dN3BLJg5
Wc64zeYba8D690w9wfETSAMSlTPvV5rV9PDExsxEUygnQ4yXSFGGIOB+gCnm
L4T1q5Py8kLh+IB5yWSuSvZrIK9RlaiPfpubKe9CB495VNj7Um93oBr//Ifq
tuV2DU1vJ8czXe6R05Ea20OmlgI+5JtZ54matmHzl2j8qUnzeNs3JTxk8ldD
3D8hwTXMi65oiTaLKEOGo959FR+z8l4B4VKpcE0zTnMJFFnSCnjMY4HlXZMV
pOYMffW5v1jbbpQR/nEQrqT5COYYXzbXowdL0gFyh+4xbWr+7Z/kKMhBbM2B
YCDwrqFRNjTpsXD1EaWXA6RSaZMcNl6jcwUhXOp/T/iL/hhq5i1fDFGTg1Yj
ymGImlB5YfnYrxq2vNM3kvwWeM9EjXRBLMfRRxDWXgBjfAcoglKRItKI4UA3
f2aH7EvJMhxOn1OW4LolK/zThSoX2SawRh0fsqvcRBA5EtJI6oKzXG/Qyy1T
7Oar09srLOZ3NWSkIlF4HIlrH4HfM2S2QfsQZgJwKrPBn+yiU3JdKGdhRQql
o1i/RIiUsY6CTP8A+14p3wek2qbHvP4WXHK1auU3nAUSTJp3JvboStaCiuuV
XqR1Qv2IXNIZkZ9nTruox3j9tiaPk1723pVJGM7wvFdkK5JrjPA/iQn1hf/C
23Uew5Dh1JCLOSucJ2zFtULQBM7y5FJezTnVqJXqHcB0LNLlkE6WBkXgTKTA
bMbqYuXcITK3DsdM6GWKecRghdWYwr8h1Iu7RMHjjKlMqmqL8Z8pwX49XJjS
OdMfnqHfiWfhzCu0zhZfBnI+kAJwrIidA+yKJq9N/vhC9y6RHFE6zmdwzmWZ
vm/wkrpFG5bbPoey5gCsbiSzsMyD48y8IkPB1fq1FSvXkP4P1VeHmmwsqpLw
eUwkAD/gEzLFnlMdSlXomJJSxwNOwNE35F/cQ+R+FQUkyfm+upX03tnKMxJl
mNaLELNIO7T0trgAG8Y8UcTVYm2g7pjqLG3sXhK9AWLV4njrrDdVT/38TvCj
Ln4u5ydQ/2imr1jvK8H9wDQG307eUBYieLcPJl+qgHHhfQxHl2rOhBkLL+en
7/V7qTgD8hXrsLMXaJjd/nAKWNvpO2lKHzyMUwRxn9QaQPYEc1l9uYhHnMBP
bBISm/tNLUNqKjOjqEuUct5q5e5wfuf/PZF0I2UY5CQp4lti+DCjz5ltRCuP
br0DaqU18bx6vfy8YKp47UkaCdapMb/sGAfw1o8LWp6iO2GhOjWjeOst+8PX
3DD2Buu2xu4F+l3YjHSfC6MsUTT9W1va1aq0CZCKvXQqEumQ+RSu8yoLZ+XE
z4zNeyjb23Ki2QQFUdHPVqZ1jhTUNhrzxrFXyGEVwdYOPuFCd3diqqnCoadz
pnduc9qWZnosSSZblCsKzsDvlOzKzqoz8KM43rVB8Uzo3IDgi2GN4kBVSaJc
XB+rMJKahyvxIFEv5wXPOme75yJgOhk1qY2dTXCtGq5EP5HBv9hyGi9z4iOV
hi91ii8B+WrA8MM5fmk2IIMLHbUO716SBDmOm6qAYG6aFFhVOcyEVdV5dBBR
1qKsRnU07Uv4yXFnM+svfxdILn1cdhdcXA52zG8igTcxpv7yE3AHVxaXJtKv
Kf2zdgEAjkRMw9023yW94tHA6JOKPnJxCQNUDp+g3BMlYiLQR3w25/0Lg7Ui
TTucVfOSZjpKl/+7zKM2F2SbCxrQ85Jcv95b4AIqP5HO0qQZDiq8691uONrv
5rJgFiR2wBpYa/I/jvi0JqAn81D1P7YZZcoPVZ0rtGM381Py8BPisILcBob3
egsgrAWpHKh/z1dGdRJ7yiPqvyUY5laqW6Ssq8XJBxIseVeV5P+7jemCwsBd
wJOBKBrICyGXQSPqLAjMJTAEXPg7bpPBB3fOenY3qQ8QXPPfqmQ8+DC8+dLw
wRmSv5sDKoje3SAyeG6CNQfjhtANibTq0s8aDp8a99fG3MI3Mat4qagdZOR0
05LRIMHuKsF/BjYJTZjshfBp3vlFj7VsOO8VDg4cfQfEl/9NhmYvfvDae9Y/
h0tfAc3Iw5LhqbJlRLbYUCzkkHYQaSalvhR03dRHCvBaQFVYPle9aiNwri+4
aKIQ/tAjYvY8ZKgxWIMb0JlREL0AyEExSk20D8NrDeWOKdN/6pMd2FaUbeBa
x7ZY1bXp5GXbs2BDcgeOcdyLDN5KJAnpsUrFCdu3hKiwonrHlSA5woMVcDxJ
+DBw3xfMd9+urRLhEZWWEpEQ77QudpQR/f4w1NRRK9piqRsLjSveGLZMvF7Z
0GR/B/MG8ZPXN5nn1p1jV0jE8H7uoTEeuYdQJjdYewYwSV8DRmYEP9IqFt94
U0yv7dQKPpZeJU1FNTk8w1rk5cOAaipatfEgUxTLFwPXjHwsohbEaGQSPk5j
6qVbQSUTaO/RIr7vWi9mBkL2wDpij3efq5A1CpFQGbahNQg7ZCptFa+Bt9sB
bBsp9vY+fz/UGkZ64HR1YA3bq6kvHjAy6PhNibGq84oMTY2R75E7zJBdSJPQ
V6rvQ3dsdV2vrBf4WKvwwlDg1W+tSUMRboVO5I5aJSJwPUBUbnLxqUFGP3zZ
72DZUgV1W00ghUtht0qQT3yNbEUK7OLkeOicbScoJ7D9h+6OKYGzBS0BQsAW
gzxpx2IDJQlpvW6ya3l4TsVwGSEqdmbSCytbBbv5CNfg/Uybd7dx9p00oP9i
IKIr1EuCe2CU7+ZHp6DVT7lFzifNEQ/lFrOBEfMFBf9AhNm6SMpMvkp4fqce
vqUkreIZgTvU3jU64bqkk4jv6N3nBS05cnSmBru+TKoQFlrISf189V8LKc/3
yRemiEtPrkhUF+OreYO1EuvbT1ouxSmvr6ajJThi+IRCvC2BZiIwgjmChT5i
dv7OuiW11zkXHjTwuICd/8/VMI4SVl/ei9yp/GK/QJyONXGwOMgYh4KCLHm1
0JmEbRZ0dFGoDQT02tK+yLldIt7+h6mXz1niNW/eg6VZRzC5o3z4YjzcH/5X
mN8SJRIUx67E//E6r98Lyrb/mSW6SNbngNxtc1/6CTnMo46gAgv/xSRm4pLO
G1qxhoG4lmlf0hvvHxfAo4t3tUHGNcB7jWP/UiD+8xrgS0hkkK+yG4jCf1Vc
IYOlTSJRy1mPqQ9nCd07bqKV0DYVg275GA+m3s++FnH8fzGaSnLTos6GcTQa
MvnvXl6rhLXbnjT/nVrWTOTkld3ygsWRko6RA/XKQfaLimwlFjJmpXAhHTHb
KV0hcV4aX9s9Kv6/njkgy2jwsQ9UkB7YOO/T+872tp7fuT4kkVua+t4OXAVC
n7nZMUrSeGvuBkwxAzaXVlbLzA/kB9g8YtZ1apJYroozH/yJHTDQ49e1UgQ9
RUy4Me8lyg7F4hL926YB/S9LHk2/+9DwW0uCPR2P12j8wLiaERzhjY6vHWNM
IrqAxcYH6u1/E7g+UAx0he9Fz5UcbHO+NsPNrMdNXn0TpudEzMXEf/9yxmKO
Uuh5Jmihpm6Z0/wldcSNaQwWMQ4YqTT88TBNPt45EOwMKqPGBMiFKSW1nIQ0
WytzS06Zu/HZj//OZDz4461+6S4AY1YlLF67tRpaAuHc3/2+NNpWBzqEY0qZ
0wkDQ+aYaW5+wSURNrBG1Ues/pRJHZPvX+JtwXP3e4CnZD02S+KMlSE3aeUW
0Bgo1CY+00mS87Lrw9uFPrZqscSIGTSEUynwC2B53kulMWa+mOXyg0BnW4lt
gFcSCjA/oZi32EyImJbLVPHkaxiIRfgwvxBB4ShY9f161Fu5vzPDGSk3Kkc+
BZ1DnCz2m/5z4jVxiumFEHvUyxRAbdwJy4SpDg6GPsRHAtK2J8fpEnYclwss
dVTtreZ7kTDRazMJa+JeW8JIU5oXRpcOZVpzkHFsZOeH7Xxyqqh3Hjt0w8TY
0haW0vGPt1V7W0V/PWmMviCVrEMewaYADOS5AnM91T7wOxOZ3appgFvgmQGp
2K5OBBVgQo9I0rHFvkRdJbLGLkDnja9ZwRe3NYvkaUSgsMW3Q74ktRMLzT4F
AehMwFtGSAYkB/C2m5ofYW1r6kI3LH9pvCHoLCziaX1PfojYKpwQ/yzGkjgn
SOY99xGU8/A7YgUzyPN/z4Wtz57VEhdE5Q+kqMDcAiCq0p58vCJiVETutPaw
7WO0RvyKqQJz4Ue0BknOU/q0DI16Qf64zuCKfyvQkSeQ77g17dFgk0P3JjUg
+HDbLEs/0d/4q7kfcaJKPQyJxPwfITyovIpT/XuK17bF0T/xamP8a87vvpVJ
eGEIAnjDtTNOzVm9o8aP5gSf3Td/AAGLdNq2NiBSnhDNjzZ/6n93f5uEKgZY
44yOqLThgqjnkrWa37u/oaj/P6XMtYB1Ny77mGYGvHLxMAlWgBIwdvo353Pj
BIQAiKk1FF+TxO0nNjxtSsnL70sApt4VhoPUsdfrtic2nA+9dkyAp7w2PZxc
5i1n4KzPv37MgfB3ZQpMXSbaZEDX6356pSaWdEO1BRDH6kVkttfZW7uWdm/Z
XhrytZNNOOqh8VqBPeD5iJRLjUE4LwC49lvagaE/J0HdJAApYe7KVCmQb8HK
3XA2uxJ337E9biCdF1MDHOPH7U6Z6hVOh+WBkLHOd7e0/y88D3rPw6K/9Qwq
W4EJDKtrH3AAj7y3xcovr9xqERTUb5FH7WLxBarY/4mBfode9s9W8mmk+BA3
79veh1JZQbtm/iw4rOazTLyvugTILZf0ID8q+fYj3DhFFf+dWdYpzsaZMPEw
35rAFi//bTph2CoYh3f00rCZpCceIIbNUzwTkiaU9zwJkF6oVKZSLuog1+5X
Ju8DIyck6h6GZ47hIpJwarhLYGDhY0jjwWcbHDGm2W5k9+d/Tab1UyrqXPea
km8E5Z4KEbfNcxe6q59BZ35fMynG+232Nae4AYUQ+ldXMirrUlIgC/KFlIf9
TXW72LF9p4rn7TC3+eZ++CQMv6MNo20ttj7ArXVqk/VZAN0NzMW4hSPQt5y4
aQJb70pVaunjgiZKNjZomV/+GKPgj+i2ZBioZxlgx1soFTyLZKTL3FDzQxSX
MduOtfY52AiaS6mHjGFserN6UddD7QidBCyjmQ+QzOojERrAuJ9/HGq0Xn3D
1KnWEGfnXUOIkoP510lN0yuqNUPalrlMkfwgICAZE2bRGpErpHzwaZsE8o5x
lpmk0kdi2wno25dqBfVyzZu0B3SrUf+EC8v5jwU/YV816ib0K7nHnUbpciGS
kVGQVKDdXGF+yPVoXA+X3JxWrNwubdX1b7fiVghY8y6q2a5qE7dSTkUDEX93
Zh9xMhpPxbPOsgH3kSLA3vPN0sic7UiWZzZOL51TmpZhQbzqA0TWSwQqV0Q2
+0vEbxKIqt/3hYNFGbRjxmd3zN/7N7qPLSJG/QdLyndRPaR0vfEsPX38L3Or
tgzr7sETTXPr9ApPR1oci9HzVoK/iWZTx/kV0c9tbqyZ0BXc08Z4lK82LSGu
CwF3FGuID8NXrsdJnqJ8p0pM+yspW0pghtZrfq2sXKduQbImcWEYcasaUkn2
nwkYa/HhtSv388vd4Urkq5HntK7eieujnqRADzMGyuDdxeoIim8bqD+1VxFY
mbpowsMGxvLlCX0Eo+tgs5zvFCNwdAQ4Q1UXUQHRT87HFWvRZoim9To3915H
0QZ4LlkU3uNofnPPA8edikTGT5YD/ZDEn/P/ANJmlxaQKBAZfTCpVsGuDiIO
fA1CW/5hugNiP6u0fwAzlgRnygmXZsh97jUmiKHIAbyiZ1eUM2vGP9k+yWMS
vQARuObXkhRrWhCwW0L1qIuLw+6wCKt3oLo3Ufu8Dt+JMtmTzvF06qTm/PXo
vUFS66YdHZqhX91xPvDa7s5eqAkswq/KU73BJAFpd3iKa8NvBgjPxqFN0gaK
jp+cAzhQo709ZA+Xtx7p5racEEbe4hLJyJ/7EM5k7wBm01uv6XdMW6MHAt+/
eP+DWM4xyX6rus9auTCYPIMRAREb/xHVB9rV/1ORj9rOvs+ACFaPNfW2ruKC
w0GwzsluCgvibGqiyOpSGcQGSWKr/oigN+LyQpg1pNXuYodgiXJH87NHBkUu
3xYuO09t2mpQ2MBNCt/C4lZZNfqi7CuVP5IBKR6hcUArW1hbvllhOvhgVuwm
vudr+OeXNtx8pP+iCqL14CwjTrEG4hPdrHQRFRvaolcDUbiPu54XvWg/1dyS
sJ/SyyJW1/4K2ZNh4w3nsOebE7D0FNyusxvsNg/mT41Dvrlm1EIQdzczYSUL
5fZaNfsGToXkT9h5xCcKuIh0xCGCj62TYfaE7zeKAo7HxtmNjPPyJd62cYvj
3kTzQuKN4VAlRLD/n5KA/IND1HgUQx33GHKohstijwJC44lr3deWQO+ZW3Qv
s4vHEguGPVcxVPqm6SLuGP1/R63QR8O+hJyep+SVowtkicx6uAGL48x2ApFb
THhjx4wnWycJpCepS8BOnVBULvh2+hu7qeBPvoH9Svfx9Dt10cyltUiNvG1L
eQiod9T/tVscrWSNqDqsSDBC97JzZappNcT+n+CjGnZyaeW4JSjcepqsalxf
4zztpTjQeBYK67CC7cBjjcSniknOOYyzGXJNXVYuukTG/kRCE6QLEVXWkoHn
W+EmTo3oV61nn0LvCnCC98Fv7dxa4ST0zF2xDPAczZpg1k3ij/cIR5nOFGsh
rW5NSEE2PFoyEYFLKvIryZMCA/d/nSY0y10AKlHD3pkRGAlVT6MUNXzUtWXp
k1aHekF8Uu6EYfObAmA4bBJqC8oSqbLefmrEbV81KherDcObRA09UuXhblQM
fiOtymtS4EHLWtbuskNXhOh2T6dPZMyooUodBGsXHrmh8I9iMdbVWZersJyC
g8AnN/PlGp3sfc678FG9voLInJjX3ieb1eHLncLCNsG3f8h4KOgwSo1EQZ3a
CLawjz/iVQ09BGrwlnQzinxrFOcMY487ghZ6fHIPZ6UFiybHqQGIx6Cyjyqp
BXCrCek7cF0bDgMnSqZ0YvS6I/omLM8bhGlPk6+THgFR8cGMVv5UJFQCQ9Ft
4wpjwARfbeeilQcFE3jZunzV9BVXxS5VLEjAWErgCdtUL7Mp5nqkhgG2RFAh
GQRt2tANdGzwjtt0cmKOXS4XTgd+nygZl0gju8fick8UJr752gh9FTmGWC4E
xqK6jp+Y+FW3Cg46n2ul1F2LRKk6uuoOJw42ZGT9PHrAYyzNFwdwc6613fFf
Dy2hG0GTRJrCB4lTPKjTXgFHxxHkXUEG/cH8tpDPGjOlLNjFQwpdV83iTWjS
qWClU2KA7mOZBSJzXiPGjYH8ZfTx2HXPRWpj1BFqwkdaUlh77P4CiJDt58bL
MbcMm5tHXePllbVgAYNRbRG6rIfevbYpIGDzbcP9hzpEzT3VEQPMK9d6wNeF
nO/PTAPPCWp504kPLA6e0xNBtZgEt6yf+OQZOVZZS4A/LrTctatqyPRatmiY
GhwKL4pFoO8JTafW59M6jLN4XL6ZcEHi1lReNcPUwLSDoue6KlqXK3g6f5ZR
3xMAymXTKJ6Z1R/0QWEqCVQWThLWvl+52A1FzqzgK10ltr2eBGQUow42ybez
tc4GQsUMRlyJBy3vhraM7U2Us52nfYBKYRvzpRfYy+UJGj65/DHvHtRTf1u2
0+B1zqNqgue+2YCBtV95Mk9dp9Z3kt8gYooNjNqZv/jPOmrpyv8lBJG+JslI
ahxvuPUqRGY9ZMUXsOtTrdibtdNgh9rGREF1KMVWCWQzfyPKShsLUXRGzIpf
YKUtp83APF+ii0RILO3kuvn23Y6fMPLy15EU9iEEfXfZTxiXwFe8sF0X44MI
bAdRwitUpXZs1Fy+bDwUL4RK9fJIz7whqf61KTbyyicy7APobAwHvLKjwlAO
U4C3QzIrKWFXEMxfK59/NDx8pfpPpGYyVFS6XxKu1QSD8GLEcTxVgRejpM0f
4aQo9RuEMdJocm/VqkiZXlIdO3x9BnPFruMq9BYIvN+M/Qf46x+zJGBHk3SC
Kjb4xmiXI0WrlOxknXL5NKjGG9JNq/EeN92Zi+BiNR4vaF2OY6Qgl67fIjhs
lU+JNeHS/aNmLvBp47OJPqyvP/Qrr8qVwZKbNfLrzXtpI5vizQCaOdYkaTHs
GPbDLr49pW92F4rio+hl37VISdEwcLxVWAlGooet4w4uHGET2US5VKqkGg4r
lZ5/RR57dEE2JYu+NM2NgTjL5N8dc0xzQ7Y3grHoVpeu5mLqlv3XI0rKclV7
3cJ2p3ufWfcrFRJKKC0Mc+G2JOwKdDgSypV0NROvLgsV5IgbUaDyr41iRWIj
Sau8YdGCnrK0SQIulXqCUyDZljfmDao8hJ7PRdodYRC7L1wJgywFQVSEUtt5
YIdELIrkFhB1rQ1lEKkPYNUSKT2MVCVCehOZXLMpzb+Cq39QywIys8Ic61zo
9pi/hwppv7ViKHp2mTyGHqRD2vlHyjwpilnaM8QUvDf+tudvYShXOU+w2n2b
WNRX12TZOLZiV5wEX766C26SBK98wmWdxGsiMRvMtmRuFCIw72qBEt4q9laY
LzgIrBh+XKf1UKhVqo0jVHlpB3Np7hE50ALF/elRkS7IyScUGhA5iSKYLi0s
6x3YzbtK/p5AFBiLHjRNeYBPtdgzMZlMAEdePfQrk5qdSWhzNzdE0NZJjXvg
UyNSZT+u9C3rfPh9aCTULz824n4fqgyTZcuzAUIjEI79K8KMt6Iy/BBC7+vS
dw/r57snWq9hggDqAu2TYsz2joEzSx3EHScK/QahGyF+mraCBT8Fa1BRerzT
XMRlREPeF5vLSMqaEfnVW0jBbuPKHh2t4TPJFAFmKZ+vCbL3Y02xEXDE2bmt
HpBx/zHYw6rJv2hX2adGeaiuCgXHUJGnfL0OzjdN/rnejKeiiAbwNrFJwCWI
ts0wBaAv9ltMvY+aa1RaBrHa+OEi3zxVWiKkYbCCrZmOtYdJqUhiEjxd1Utk
DuE9EOuYfcp6HyHyN0mXV0wjO89Y2qmurR4uuPAQVDrZMcaGnJe1xPtridfx
NGYdL3avnw/uxRC3c6+qd1+LNHojyr/2J0UtccIWDVUj+6oAmH7kF2xkba6H
JdbjQLz4yqkqO8HirTvqJ8mkTWBTV+sbAPUfvgC32QxJfFaELg28+BCRB/CX
fck+W6hBOCbrZc5joCmYYAEhB3YmHwEFyWamaNN3EGvOcPCOtoVu4bMt/Xrf
pVloncbFXLxvhCcYzLUWyEHC3VcmnUu/dr/vNtrAb5iWK9YFhL3FXlB1QBDo
K9Le/4urt7C9RfTcjl8NSu6kqOOLChIewGdnwLPsFFHqjpmZ7dPROVo3cgtG
uM53oOSJzG87WdVluzV9nF0DS3qAHEN1AYg8wITaFwTOXcW7gm2Qh0UDNrEx
SNwn0YRhJ8M9sM73Bie9ahRPRGuY1knGlX7gBGP5+Q7kjkGxoV+3KjsNfcmc
wuZ246TfoaEGj36C3jDFwAqBZ81jnTnU28XzT0SRgJCsDobcqCZJiadOLQwa
oMqhroEBd0jMOQYeQ63L/p90bIhmZybNwslS2nK9ChblCWdf1yz1doPgBcDn
fp+bndttaVlZ1izXeiqQzuSKEhdrJ08szep5h1Yy3TEYoEQvPrlutAHRsAlE
agBd57qm1fh79eU2+VoWQrFo/tYsVUmidKkUMe0ZLVy2mI8a1EsdnaI2epup
dzBTc+0pIqxrGaKYw5OjpqcMHWocBG8mIjpUDVhcjqCSsJ0DXHvV0pXPOK7E
mgWJJcz8sMcjKb07591Ifr4hW77Hs0ZLac+yqkLnBr9Q7/c8X4YntTc2CHQY
JBet/3Q3WeEdARtO3jjN/e8d87Mr6tRRdp8t666igXTCTGiCjHIgI0iudFZ8
tvMBssT/EA9a6/eeJP9USYoi8Yfk5mFU9wya2Ge/OTGHa+aFeZlWrZ85YkeW
Po7EjVPWsBBPH0XzrzsPFo5ISS6brsDKosV3HMii6qjCf1yaw3ogA2vSTikO
kTDwtRd5FCNzx0crnNKKvJ8ruHo21wi6Te0d1IudjYZd30wPzdA53e7vp4fZ
k+WeKk+S2zUWaKTGbgbHnXT645H1rmS49l3lkimOEqnmV3P7tLwsq/Mx9WJk
YLgPqZJJ/rJTxDvSw1uznweA+tx9mFsr2xKgiDwiEjVsrX3zlh1xGpTr1i7L
bFtouoR84nPJ+dMtFSapyhrHD5VRT1J1e9uFVcVk5NZsNLsdK2xizZwiCMZA
az+dfbVS7sno24wS4ya5mqWNvJhk2t6JMAiCYqwdTWg46OslDQTJZuB9FBu+
MmLm4H38jR35O7Ft+Ee6T5sIHIonaW3F/Yw1KuRyS0Z6OPhBpqNslkm/P260
7HpZXI9SwYhx4Rs5XH5C/NfIPyfos67Faedp/Iz+xA6iy9xTmiuFqvJDlVHj
Hco4g0qr5veXPBN6LkFy6Q9xu14gfnlvd2RT8QfZ2jxivvfoDkXIsaDV3pAX
L5Z1DNRrk1wRtnW0pJFsfO+OM2VxJkSqM+F9A0Ov+CqEFINYEGS6a25ALSs5
D/Ive9JUZ96yxCu1JoCDj6Dul/FlpQ1HQR495wgK5qWQFT/pFCRl2YkLZoRk
pRkpTmVuD5D2/jGJwIO7ta/kOV6frYLulqIXV+ll+R+LOEyGExjdjEpCM5Gy
YrFU8y9utVeMFxWECm8ANis9EZ0knHefX8tk6jCVEg4jURDFVZbbFdlsiRTo
SJcwiSqtb9j3ipeoJMZhDKo884YaAle38VYd0RltPU+anIjknOeG8KjVqI+3
PLqqOqn7/FXdN5PbkZPc5iHjZEbRlaCUHGSk7qb4X4FVJioemzEQISOykFNU
WTc9kdNJY/THQBoElCBA4/qPB02i9CNv505ywtf/HUvVRXUNENDIs7RUVaAG
4gQQfgPwKOBj2DVrYkQ4huqlARj82CwrrfMZQuvVaAg1tA8MFUzKaq5frxRb
8NbNKyDk6k27uCzae9ZqlMo6S3/ixHiu8XXzbe47FW3B/rvXFEm97hiuEI/g
3zaJqa0ESUXaEjrEVFJY8UBkPXoMAafnwBTicZRUMuOlozediuW9YjU5pSgw
rnIIs6prhhichD9tRfcfhPneOGjqAz99zn5GhIiIrAr2RY+/fbOZwwCcQYPb
3c6YqL3GnVMjB09GgRmPJg2uCANmqpTHd7BbC6tw/BwYZQ4MEM5V2radC0BD
Npd8YTOF6rC0JCA9Aq3mbRi6ZVcoMuBZhCbX7eIPiNkWNRM//Mrumabk/Flt
HSWpJG7wmpxLv1iI5jrfTfxLn3+xQ9ybS1rd6jJkvwcf8IvtGWaXvEGGV9Vs
i7Drg2n8MfmX59D+45WjMGx3d4T34QBD6rgeIlUngXM23f0aXoS5EKhguImx
jASGZsVvwbLOXB4KYJHqxMawCNJRu9W0Tlu/t0AyD7Ou6oQo6/vvYN8Zq8Ep
qAemPgV7i0xQB/DYPxYyr5UqKBS5nzqZ9eKIl7pmtmtdgHh0jAx48J3nVl09
7CZGUhz++Ue3HM0+1LhwF6Ts/+9Ls28n02G4gq9PTq7ue8Y0IqyeeOu/cRuE
jKRlZWaUeX8QCUd22c30QDJcblDuqJVEKxNnFVGQtq4JegevMk0k3Pk3GdYn
L2TqO6nmFDiu/c3BWjDVSGMSnQwslMbnZJmzxn5JPr14mDSV/Jordeh2s4eN
ZO0OQclZ7t/o+yBOw+Ieu0FnV/8XEbBLuxpTT0x8kC0URGe3bGkco4DVicRC
LT3OL1IIIDaMOw5hDSraZXVrSvj/G1kcrQPyeP/Asz90H67ao0yOED5VKYLF
r91TCy7dkEvzhm8h70C9b7tjzRMPAId1dPoutkVeY4R7sd1qvFi+q99Js6/L
RV6n+3iOkg1B8C5C5D244aRvv2jM0AlcOIxRjXv8X4rCEcNkS3Tr/DFkhNUs
AQ6+Y9O+JZAWRZkE+WWeFkkp0jGjN7/qozzlcxtxcaIs2T6ii1PzWkS6sied
hW/5rXVS/YJZAJlpD6YYQqBAWN4AwWEmIhIVkLA+Hj4mPUfzMZubBmVXIpfE
sJruIZd1kZ7UEmi1Dq5it8JV1MLGWmnX7buWiGRtERvhGMQBkt2+EZU/W56Z
vM4NVUav3YTSUSrLWm0H4iXt2n+beh4IbSK/pFTKghyCz4b2DEVN/J7vh0o6
pccdbK6lFZooxSbWYLA8I1QZEfPfd23KDfZRbuOtVNSoioiAggPnuQywOs+t
lujLkUrp8Me6eeO9qv0HVIzUAhx36XqHQvGZmLJN0tb7rkeB1/P1Fh8MfU8D
AJoFh+2cNudGUUEENdps6nbZmHb/ZhTlGwIuHSVYnDbRXDtxfgEpZfa8waKl
HTvakgfOwzZPdlmH3otoxKY52M29bw3m+pdk4WC566sFyK6m9pdd0r3gl/Ei
7TtOcRLi/bA1RpBZ+rfstGfVwHPRJdQUJ0UKZeIpDH2K5fvD0Cm1wirmts/1
I8ZxIFBraDsp9WA0M2MZjSpRQTnJb2NtaIc7GVZP4Ln0/b35fvtkHV/YCymO
9Ly7fLZPhHMtAhQY/TH8OsX2NHeTX7u14nvSnWXxUo1eYxvTXatyx8ia7E0m
FtX/OcbxEWAvObpY7zkQot1Zby9Oja/i0TLIZxFvintJUPHoXiJiNCrjAoUB
xnIPiOdpbHbr3HhfvIXC4ocG2NEdkv3AinC9RzDLsLVMFESDRI5hgG66Whu/
iNWpnXX/0x2gTYiibkDJy4lpKESaFihLYI8YZrqNdx477cYVGQXBF7swA9QN
ff9/lFARcg49srn1s0j5HyMA57FsOKmq6DSSaqnSR75kSCDhHI1UXTDfOgtu
j8OOI5wfN+/n3PMsxWj8S70bgkll82f/n6Q6obom9oowwo9hMkRpBtzSnNiD
b5MquwtkFV8kKYIXP/OHkthZf2GVKO5dBhRqnT+ZfWte+WujxmooNCTGMIQA
+Q5/bW/ZuCOCyCdaujeHPYa29KmlselXUCLxBO8qP5ykIxfNjCecEg2IYYd4
/2OScH/+qWrhTmFGzQ/VxG+MuBs8lkw1fjaG2LWcXmvfrmTnJH2RzH/20BsG
WIPX07KxPEvbl3UpaiuT+yZCWJAagfJhBr4dntNiJW/GCVMIW8HrAQDxS6bH
p+R7ll0Ktt1/ND5+uT7nBwvIQc3qNY2LI378TGleI6Sd+qUZKqGD0wzZ/hT2
dsMPfY3Ml95Qs+18jIwrSd2Qm7SICz3ZYQqw0pnw+SQgAHh2R491GX2lXx7V
6DSs0twYejLkIpbGFjTeWRfDlpPvNV/w6vRLfmTvh+au46qfukoSYQtFQrk4
DT5pHWcmCw8Q3Pkc5/uyeuCbW/GiC6VqjO5FGIhJ6qVYvZHSBKWZD81Yr8AY
bhHXdr0xnXY3gplM9ze/lhZEbGktRwOsblTg/+tdkYjVCRn+bQOQ680Wd5mc
RoDxcDxrQXQ7j5LDqilQimAAnZQkTBCiSlxmhGRy8ZPVf5di4P/79ttHAz67
G/Qt7A0IaMCXfg2ZGbRu14LIxz3UeqPJ5rcHu/vlS6MWQHCdrirC3d3FZ7kU
lBMT5ua63CR6ErNvbrALCs93c4d4b6isH7f2TIWMgLVRQqM1wGF6IVsnbzsR
oQlp+aU8/nCLBcTBd30eWRjRnA+RYYyaoshybvn9fKUYxBrCymCivij2eqZo
VRlDk/Ohd9r/3uXFv/gKLexvnGQE1f7HK0LDpxhCENTxQFKjndNNIMI8q+Lu
8qtoSqyxDEpVrA4HXq1d1CoZ/JB0bctomwv+ganRfh66ob9y48SkR3G6U009
fgmNDUe3h/7JNer8V1wQzizShEJSGM39kL28QtVWKtlhC1KFOUaQdI+ewTTq
jZayQcRWR4MIwkkSiR+lhEoc8wCJ2jEK4EGCXzJAjf2XazIJ+V/rHte1LinE
6BrQBCLb54AMyqtZ0++boOq7duqE5ZFFH7y8kc4TRn2/7K7pT/yjdsuGhL+p
d+LXL++dA/AENVqCoR/Zm9HK8/iAjIWtMwdhzZhozOicIG6YLucKH7rdYl7d
Zg+o//b4mjco0dIFica52vjHFDROoNkg0FhdNvC2mVOAAaSjbA6+Pkiwo2Ft
KX1WEQkR2iMDPBOPTl+vLTdZELhdjKR+e+tdtr/H6MOMplGdhp45C201yK5h
2gWx3coPeb6zXS6VgWI4hyxbexPFcQIW3jBLiyUGgb7v4DLgJhOfg3qpwnVp
0FDEmu0tuI9QVwFR4/QdzABGAkyoblrx+qygiLI4qWVPDgsQb1C4PuVays1R
Xyn9l9v0pXSDZRPyfhau4pzsajOMx/YYmUTRG3IHKdji0XCHlWDindsGE/wU
oqlSbtI9V5hkTI3AdIF/pNQCk67Q4eGfLRNBRcCiHP8/6BXMreIGWlx88cEg
EHs75y28SrbFHEXCAIGA+9In5MBpbEpxio/NFL/Qt0OnE/6M+JOphR8HtHg7
6g8BM9AUYSya/jAJ5JRPFPU6Lhzk9+dJPcGt5rCV2xcpQe0M0hZDqRNHYNyv
1EqKjqrx5l5uXZj6aDA1vb1GGODLbYisvD9k/fKmJIjFrF5AhCfqXpGVOZAU
rmXSYkwD2AGoEQTdSLoKfacIgR7Pp5wH8bI5v91ilnUGOV2akBBYnqaf34cN
7jSDb4Yknb3J4atYFisZDjxd3lFQ5Z3zV7HrLJcXGBr7RSm0WUr9GbfiwOBg
NAh5QQPTwtA9uKynqHRY9DDBylB1C9o2cbZat9R0cmGVc6B6Ddve6Gk3D/tM
IDHV6OwZQIluEWdsb44FS2T/KHMX2y6yGDUqMsvFSUAqZQhDPllGuH0hYPYt
d44Sz5SjvyUah9rkn+nPRII0ak5hq7vpkHzTagFoa7v7twxLV2GmpBrERiAp
zIdfuy07rSbJB+wgGqTL5JOdTaVOvOIizrCH8MH8/0fe0D7wyd4+by3Km2c7
xB/efADLDhcUFeH6uiMXA2B14gSur52AicNwmrccaj6s943UPBLdicHwcNgl
2jMSiFE3k4GiIc8Z02OmlbNiGtRBW6ttenUA2QV+b54Gfqi8BK4SkBUfAETs
I1dBbqUWY1vnE2NUsgGj/zdzAdV2JqTvVnF1AIsgW5WagPPDwyAdb1AhcX+M
gD6yzvv8Zpqxg6ORw4/1mM34QOpY7M2NVs8+JB9Uiq73TeELrBsxRUqANMVM
wYpAEV4HjdWqEP2EMWROTNoBykOaAvadD1YTwiAOTn92a4N9431XZNIT5Es+
8bqSAQDUU8LaNt85XAoku500D2/SOHxq9Y37Ll3TrGuq+dBmkNWXH+jupkHU
C53t2I5+oK/jYr/ptKfJCAIwp5uhgGf3JmyIauV7n1TUb/weYihTCmCus6Y3
8fbPMys7TrQSwVp9dcWOUgE8NmdSPJ3Bvr/77cr8RoCk6PVqhY2gxebR7LLy
gnM5zzrf0Dh6yY9TLAlqHjNnn0urs3tz9VagNUjdEQp5Byk8YTDJzaMnXqah
ql4kO6uPljZfHBsyYQPJdE6mg3C50BKgHd3nkg/kbA1MqNAlFVB/rF+JABZz
q29PwWulQNs2JYMuajfi/xGCJlfBnzTKN0Px8aGk1kaVd+c6pnVIhWCeMfMq
l8SaHy5iCG6PbVKWjr7DMMO+h/kEzvkJTSpQjBekBktoJhT/+TSA3KsR9ZfI
Qo+qpxsZLL63zIpRMqD0LizX9SpR8SoCIdwVacrCc04a71K9MTzDyZ39J3fg
YSWt4xrvznKuMjl1ItC1CCs9dctxgt3JOvEREMtX78NW1hnG9URRdRJ7NZ8r
f3Onx5iZdhg2/n/qbWHUJsx/fCFA2jqJ8WqyUp4fLe9EWhPKWlDWLnaoovgg
UhD9Sg+tQ/12ZDk8fuanU5l24I6Emqf19yMeaSCavFhf/SiwqZTf/677gh2+
HBA4uVhMciuZyTbumH2sLkFLbiFEpMC1p4ewlN8aWBlX7gsCvXbP4LKlR2hV
F/TODj3JnqSOiKWD/lKCMGjrLdkyD9vfvzV09fEcWgZP+Srl2GCILncTLkXB
L7ivBv9gjujp+D92YuhHBNqwQT4ZrmPJdasbhQI2b8bZnzzI7p9ihu9KfGwq
Isj+/DeAWry49wP8/c7MQp16uZvhNr9RUJkq2IZ/ESiYbnHe03G15XlakBPK
p9avmOpTxdOdkqVDGawhJHlW2kYBFJCLYSlnwn5Bd0x+wtWW0xBVa5KwZgmN
ocvTuXwM6hH7Mr+qMlyiVhtQ5fjS2JC7eT5TX4dayj0raZne+sy+ORv9BdZQ
orPalkn3rpd+FzS+mk/7kcjqvidVSi4wmVNl7V2rtDQ06JdpWTjSaTHefs78
eEAlUPQU+NoVoCEMT4G3MCEWiV+QJTaP+VFitaiVqv/WG0qy9bCo7hYqfXpT
y8W6i0rnB+6tkKxefN0w0jIUEuvUl94CsrKQ34cuvY9XMKlWq4TTrha0k8EO
9ZwmJhNgMTwfijko06h+x2hJPILpkvlswuLpfSbI/O/SDh1eoYnKPecQ7DGz
7dWXsDK1fZUEJxUTeQBONOc0xBjLDzB/JedkqHtxPz7lFuLcFqf2j4ftAcvN
kh+j0sXn2I7rtYD5HDPZgaUnKl+Vl+vuxScdmPnAPiCI+38D9dHsevLbio2l
ij0MhIuIeZo2XMBcKSSq/Bsg7ZxETbaVIWyLZQwy5VxyWgzchKB+dAbWX97Y
73hI2M/UiIe0sxg66i6WczmIlKbnUvQ0SYev5DWPwT0IS5deW7O1FQ1csEd9
yZfiGJeeKAxUt+4TL9BE49+0OBpZd2PTVw7SNY+qKk6DleK1JvWBzLvtb2AA
FSsfFP0FG2gjAzlXod3Q5Ddh/FtcaJOYwxTHdgRl5GbVLmeMeChV3y2I9GBo
qIbAeDK60BwuBveo6fVQ5y2V+RHqFBp4SzYUYtCrUnnCGbuOSvF/jlYcQJs5
oztGXvQrUUv3DCFNtS++zeKK+T+t/C/+v9SsUY/vJJf8l0YYInnJTmIo/Fvi
MaacqsW/y519EslIKHOHQkhM2cy9iYdTmjJY3JJETAP8MRTktdeUk8VKTe3g
G1bZjb4+uZk0YM7t2cd73EuI2bpqMAnqumOGI91vpg/iuEUf7W12W5cyCFtS
HyWieuzAGaaRsP9tzXIWsRGOo6rK1G3bqMCfvItQz6yhTSX/kwP9uku3dKLO
cED+jm8CMcuPryFqNKya2ahnUk8VimsSIDHqV8oA868L3fGnZwZwzD9XE3Ml
vAoiCSGOdChkzwiekrDyDbln/QNf/cN8SxZ+dsZx4pqUwLpebs/kgP6605w4
8NUhjt+noy3C/NuAjIS7sHPvDb/w7RyohPAr76NbyQ8dYez6DB7DhqbaZE19
V+zqWBkRufYXX7t+U9YIE9yuSibZ7RZ69mCIN7Uhxm5GqBvjH+OT8WWgap2w
q5aIHipFVCx4ztjhac+9g40pWcmBGBjc3A6LDiIy1fuulUxrijdzWmXSTzMb
WkZ+fVF1nZW8Lisl0zolPqk7nfqmOr/twhsIQK4Y3VpUZ/Z7vdWmiWcMEfoE
I/y56qRhJVsOpjNdAPPtYpQnog8rhdL9YWHwgurzUFUgz+/0byfZX6FEPM5O
ODRvFbQlX9ZT1pmnzP4BQ7Zq7WdqbPG4REsIdTVD+DIYH+pv1Nwl5+XauBYC
w9GzyVm5x9dzct8jDQm++Mruyvv2Plnk5uuvYqzWayeKbnFH3nw7y+Ua+pOj
DP9fyykNE5Yx4yImvbYDmiQ2O5nIbiAJL3DiMlbb0YD0Dx8tkozWhxbhPtS0
IOkqdlPsf015ruf7quNtMEIJeBl77Yb9QvBgM8kg5Q9xy5RL6btKg2E8MWs8
v4v0zb51S341zerf+XkZyL+XkV5O2epIlrXqQf984Wt868Tc1HxrkLF+Psib
KjKE7GlFsCK/SgSn+X2dPnGV+sTw0FK8pvNB0X2LvmnyXL/DYtXF+KzQizpi
8QPGftmRf3SVJ9IYpkIOLZFLTcobtQz0l9VgmlWIazG6BKmuqs37L2nIOOn6
uoPJTv71V2LOF+KFGaO4uPLxodT37sSBdPiXdoB/iVrTB1Xt3ijVq8e9xotb
xCIlNHjEfJvfeLk4LxtUQPfh79NJkvyf1mHkiE2csLAPgZ/+0/z0R4TnDExQ
VSeChtpuroH8WMEcgUzN6Eh3eh/U5PAlXvzic+eE8rkYZXbs9oYZ8M0HmhSh
sF6YmYPwxdywsfVmEk9g4NC/S6YllOglZkaPqan8DHOQhaDxpiGc/zeZlZau
KiPArvaf07pkr9NOEsYxVgEM155F+y3hEFdst44u905M/Mubh3+0gBAqIvgb
knn1P9SSHgFNV/+BpmvEioWK+AU+vH+VCb1cHjA5Nb3QE5RKoN4OG53cO8Lg
Ez0tqvQvNMjhX8Ij+wqbVvD34E+zUlfCaSCqE0FjafYhitcvJTCXeRXZop/X
uU5cJS8gL2EtE+4R16BudWg78xEFcNFHOYyyzmqraQr6UuS1sJSrBoR7xnBU
WbkXhpddsSSkHmbXEqyZPBAAEUlzlAtqIaXHErEYidjMrO1YryN2q2cw9q2B
hFDdt2/ZZN6IcnPxmS6G7BmT9tfq+GB3vaWF5s9GJaur18z8y5cI1CSiSoTF
gLM6iqDkGAV5Qb+Tpust6BTFB0h7NrqS1GnXCJON9mXRf/4AMel7tC8Jx1Sh
1ZlFhbHNHPRqE8pbpBf0kl/VsL6kKQopavjhRdRG+h0jbZF9QkUaJog5f/Zy
5rmT0u4ghTMK3meORxtAQnZ5JxQ2s43we4GAW0FW2FRXP+8G9+bc9CGtxi7f
ExEp8gvqKsMNiVzTRzgHYnj8l4pxBBfBc3+qbhXSWsTZ4wwwLc2D86GXT0DI
w96/AIYWo4/NwSRYaNXPoE8tIcys8FD5+cawgJJ/vFNC0/NWjqeFl55MZC7F
n86/ihFjNU8SKhaIcknJ9gAA4AKWOa0p2Hd2sgBv8rKjBet0/vaI8bCpNJg5
SRcDsmNRdnGNvMyYWH+XMgcZMfVCKoU6HmkRcBawLqU7V5SbPS9WZst5h9FZ
eta3QlpsmGSt1ulKd0xOfC99DtW0vTD4eLQl03fIZ3/9BgW8bjk3OMpnLQcg
YaVDQkYQBa9SA9XPke+YZtxHzAn/GgUvZDK1vAE+0ZlslRkjFns87OcPHnl8
FXZ0Ge402nqIkQsb0MNmO7VRGdQ9eLHZ5fE+YrB4JD/C6xc6gmCh3//8aFBa
+6az1LHGJF9+TNYiUZNRp5K1JX5TerHUC23KeyfAiUaZmcTZyMDvG6AFC/Ox
pPhXwFGthQMoD2sb6u21B8h/opPGOTYR2nTCzAVtqsjGo8T06cSDSTlUz1+m
N8S7R1HChWrfPWt30NJnBROOS+Wwbo27etphKG1osew6r5SBwHlFicr1+4kb
PLrFUr+Rc8aSUrzYtDsdOVyUeDS0sYzQ4rrC3NsH/FvMOXf/TDjmjKR/DzBG
fec+HbF5QUJCKGBUhy4ZzcXY6hTc4v8SCQH8Ffw1tui6ILHqNOrrk6klYmzI
odQeNE3xz9h70LROZE40vdEgXh1L1ueb4V5oRliX/Jb8EyvwXCWUDsq2Rabv
WU19G7xHsOZoBzt8KAegRk4lYoQcQd5Lzwlhyf4kZEdHQ/s2QqO1CrGNTh6p
jZCjOTV95sdjDnGdKj33K7hfTbib+gvsxoGuRIKJ97itz9cceM8aEEytDSI4
cxTzpDy6DILx8JG4y/UwIF65fiY5y/RVW7VOWuddzghTmgjz+GhgWgQhdy3s
bPFUviaWAWpoYGYAU3XbtA2PAxbJZcV00v+qxgO5fSl3ZDPn3woun7ekCJmc
+vOH2bRnKfv6fVvD0pkosS2/gU9ki6jSh0QCobqjG8h8IxcdRixle0NtS4az
EHyUNy8v6ZD1zW/5nNovXiTsMP71GORIknZCMK2AwUV7LZJjgoL9x+Ezufz6
2e1Uh77R7zUml/UXbVsyfrdsPGp+N2nVy3xbUy75oQdEfBeLcY2B64hTFKV1
qg/L5ASOC2dCm+BMfjQzTnY7Zgk44XotFKXCH8eOMgkajGpKKPMf5pIqAmYS
FSFXhuinRL7QTjh8F29Tytmej1zD9Fak3PLe/sLYtwF1tRRTZc9UASNZzAzh
8WDcFF9X+sKzzq/8zx9KCVwDXh1LxnVxV/8o7LcUWUfsC8TYxD9xpZ+5rS8L
rXtcInaAhbjHfaPMPcpLVI5OZossIpxYMJT7HgGpD/RSRAvjGhw4FNC74Gby
+8UCj1t47kZmiEFnrELXsAh4QhEjZS0RAVwc+PGA+rWtnG6T+8ICZo3p0SEa
wKzeFywTVdrJpwFaw6OKo99fWeqdS82X2hfBNRivF4z9cWNuqvmCv7UAzkUk
gn8VlH3b+6Zr/nIhDhcolg8ugl53wYA4JNOhV2QH/6pB3XXYJNI4SgcrlWmv
gf7sPdFZZd1aGzNdLxRD5epvayYtd4jbCJTHJplBvF6B2PT//n2lmFn7TDiV
l0ixXxRe0mXym3jEPqFKfL3WBrHmmnEoJM2pKJCo7ES2RLY4TxGM7Rn1mkrx
uWfdAZKbah7oZ7iSImgK16afFwyy3iksj7dzH58jRH9ecRbbMhQ+rmTI7Rb4
c3nxZQ3Yi3mlI+acSP8UFBBrD84ftUponqq7xK+AJc4v6WVdQGsaedL+NbkL
MBLmVBOUvVpV64UnwHNE0AW5bpocNaQngEhg2o/G3NhmrW2i/jkAx8J1xNm9
FVrM/XeO/R/QV7NLDa7OFQ3eDfo6PsNPYlfs5gwRTvlFAeY7PAVOFMi6ytif
GDsopJ19Q6rNchPHuY8PenEQ4AzxQPuoRMhnZOswAOPzTLzfOuk0/vbdZVmm
4e9mh+DZUcpr0d1DOYcNxligkBWLrw0DVMeizLsZSHVqTWh1V00PA1NK2WNj
BYjnRnscv7PiWLTau7dBk9uy8xXrdA3l4T2OM4haxUIBBvRuVCPB1dN7zI/a
S/+2NgYKZ3sUyjGaSybxhAo1OEU7jN1zMl6mfnCwkBIAnx7c2qq53E+AZajz
RpavubgMUlHygJvUtZo6V0R8VI6RA0fRN4PzayYd7rNy7DeeJE6NM8QaKhiy
RhbK5rTqxaClk+/rUYn4/wa/USBT45MgQ9YfXEvFd7rJ2xzv+rxqR41e/IiJ
i4hus+LM4NgORefU+8azqmiaEP3bAJ7Y+62jpLe+3IwfjAYKBZ6rBU/gTj8n
wvMl2NcBOBDkO3NFRzITyxAggBBdRSGlE+2AjpENjU6QK0wVOZ2NVzqOXLRj
t/8aHQbQuEDnmbnOT/Kswcu47M3827q50X0bzHlQ/LdVzuQhd0T0rgP9MMLK
jf+4FJEwduF1xLAjVmV5mc3y2VUbEVEqNtWETpS5Ky/5gu2LjefZnQPKJ3ks
TPR5AxO9JvwZ+HINvxlkax3GxD+pV+QU/AOGT2clS36Iwce59Qoxq3EJ+HbF
b2De1XPYh15MCKz7rsMkYf4UxjLaSGsuZtgJd7OOh2D/OwYzDAWj0AeP6gSz
i0tJJty0pbo7hETHtAp345GrU1yOyFnGpxHUV1OD0FFi+4R6SmZgbg0DGOfY
mKpiEUrgBn33xW2OdTYAe1i0ayISIeiWbWZgbFknHU/q6bvPH9RkbNl/L7eI
v7yIEOB8mCf57Z2Mv0paGxr9kCcpDGxhXen7/AEx3vZReoauT5d/5JSwHZEe
PYcxgA7CShouXObwkCOMvOMmEIPOG/YWXJAmcTD2zOa9rmmdtJKb690RQ03W
3IgdTKr9pbndYce/Kp/SqCOL0+85ZTrU9cn05ApeFE7S25809zFDVi5rfEJh
RgYWYQ4bZ8eaG6Mmh9j8mRg415ALcRx6QRbKUk52sKl42SjyuVOtCDUSaLpV
hc5pfARzx/S2X7iA9s/NvIXQNpIEj1ZwzDOjsDzHak7eJ3FCNTnH05ZC8Q1d
X18rfHQzTlfDoT/Bf7BdvKSVC82RcKTK1ItqplIuREv13cnRKqZveinxsnlB
3GL2dJi/ae0bMR7rbZ7JVI9Dr0aO8h0vsd5fskDnFdBr05cjiUfa4FVTo5Jx
pN/1BsqBdTHDnJyP1VzgpWP2ilcRjkw531l5miEYRXwVnl8xBKxgv6mzgHi0
0y+3ps2M8jo2JqfC8Stk4EdHd7bvit6WqtNhMYLWzA==

`pragma protect end_protected
