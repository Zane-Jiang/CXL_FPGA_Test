`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
IjVx2k8MEZoz6UzXM4uE+D27TZGcoGm+8qu+QK1vxkFKzNF52wU78otAtrV5zM/T
IoXgF2ctG4iyjO44yvdXmPe+gp5Jd5tV7g5CZ8RYH9x0YgHF7hsQvOu2mCKcbtJj
/cjJk8G1OyYr4T6o3bvGo7RPEUyYGAwQugRukjtj024=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10592), data_block
b5GTFAj0BDEaUhgL8UgkMfWghBd9A/I6ZYDnySKez6B839SS4iBSnwSAOEu4YT8l
twWiRjUkG4BTQCn8i2vH8QrjI0rRspBhkktgr/uXSN4q4R4I3D+GiB4IZpfE/0Jv
hN1fTtQYU21snca02/QCnXtxK2eXwTvmg84SNBTyOhxXYPRZoiRslKzkulZpIShB
1EG+zJXXv2E0Fnu1Y++J+eBiI9W8Sfby9cvyqeksMJLneIzw8pjBKj+DbSURFxvP
Zyk8vcpio3Bh81mg/mqJJAqt9eV91VxRapylzB1P5aArrRTAz98E6rD5+A2Yb2H5
+LkmoXsQ+ckNT1YTaIezukPMLtGoeZ3EbzYJPF5PwVv6kaQAvI7ywnjLktJUhUH5
sFoqkMIOUI1Uq7zRudYMXiNWo1wW87CqQSmgYW0vhcXDKuBbuZ/71rVVvBoBcxq/
1Na1BaSirRqYZNh4icelASuVmBeZh794wqUksqHFaZSxj8cQPmMe6eDw3EJEzjtL
3CAPcb2HtKZYwPWx+Lj3RlQJXNdbC64kcw7H43ZtiPnnsbT9/a9xoXgTCM3gdh5S
ia6fKjJFfaZ+HWUsecD4JJsddlrx78kz9tiMmdG0hg2KWZ9uiXQoxWSNB44ub+te
Nx/zLJ5FUsQVfwSRHintR5gajzjyH1A7ObzJOBincMhKKlyx+vLok8aI+ezQVpgw
+AwJXO79tghls4ugb1MOocQoQd60GmBMOUc1RkdsIT/F25CTcl/xTNz3KJFMP0so
6Y8MTFnrRgNyB66MiIpLJvrH6Vg4ed4ImMSTnkIYQ5bc68kY1gxaGfeyQP17i2Ma
HTTJh0aYeqJXG2QOKNS2pyjXcnQyHd0iE2qbYgMUTw+TLGkh+RzxIxxgDNCVZmJr
wevshKElg/gZi9IvNEE525MqjGVh/5CxKtxFUhGgv4K/no4Vi+v9fHUxSzALAz9U
pzNiEsOPLi9rFE9F/GcCCPS83j4UcVD1kHgUwxR4dP/pAdvOvWsaDLtgOTPc1Uzp
zjDd7PJql9icSep9bgtrVwV040aFJxn19MRu3DQ0Q6CXw3CUo1oti0T3BsFA8FzX
xEDmyQLs5FzNTHXD5aaFcV2737+3asjdrA7T0Wq+WZIcNOcde0yfXhDPW8Br6qnk
y2B0iWObLFBQl3yacJm5hbnvucUMCYw07ll8wZNvUiK0K9JNrVRFPvRGpfBvr+Bt
3zD+XSx5ijmD/7uHoQ3HlCcuKsxtLwGI46ywsS6fSXvHkRkcrV7Fnt26saRH2kIj
7vK6usfYrqwW/sCTslozG85Ha8PZmg6/gzZnYGlrlj6TOCaJspYro9AYoPOoHZYt
eEm4GUxq0aMrjbCnL77ftxuOMXcsQVKl48b8OQOXlFwTVGTVu07b9VTquWOv3Zil
OLE5/V8w8hhvO/hq/pVAyOpcP908XhK0U50HF3Dv/r8uSDz+QBRopfFSaRbWHGKZ
f5q3SwTBSwf8R2IhsDwvThNO073B6mnVLbqf38zKGUal861DhL1mqUvzWaKLrHS4
LYgEnqoWWUlaUlrWT4pBjK30sCyDPsh9/c9vT2VvkqI6yXzV1I400zcQ+lvVAS6B
mus0PLxVH5CvxqqGHNY5dMarlF6IAXVHz/cmHppoxtP6z75xNA8UK1XMZnOYTYAm
oy4bHU1+GY20vbcIwQJv56OBFMRuy/cJoqKDxl1wqPiSdPta2dVjyj4eyMuatAfn
YLwAOwgoreaTwKgWSl0zJvbZmBmTc80TM06lwm6yOF365ewgYjcyMLdKjeHwefze
3HLVTL0cXbxgNK7vHgBi3eR5WvEk1GAbCqNQrP3lFzvNeKdk5HwUmD2OSE8lzJlj
dJTXY+rBI9SZ6NhTsK20miNsyVs/WCI0wMWvPx0gksYJcIL5tRIOl+UIJ12q279v
wihFBlI6IW74QYSDqgRxg6yyZ1WIY1y+ljFvPCQQbR1TFOuyaKlqgjfpi7qKWkUO
t94qzZwFlxfRDlSIMuQS8wWcAGsiEV7/RR/E606QaUeVVWGvegPYCjh0okAFO2tZ
H7Q51NrARvYm1ZC7hqK9GrnwFLJpUYknKo6ett3c2zf52hh+Yuo54J42WzNWE4QN
fSXvNgIvTfukkrQNvILOGwfN7r7wPxTMj3+21w2cjI6obzJ+CxgOBDjlDaWBPzP0
trZn2nbwCOFdk0Vd7WWa89xxSczv/Yn9LkDoh+DqQOX2BHQGWXcnPXjrmGEQMEja
GK2VdvKYEN90CcVaCntF9Msszhrfamfnyl8MipZfZlTpqogxvnC9s05cnsM8SSyl
FfGfhjeWpG0GqF5jZdQsZodm3xT1V7PnMBTKqyGBFJFbO+HbXO684dYj4ddO08LU
Kl7wBZdOng/FpGQ03jAbeqchhwprEqQzJ/2/L7AMWsFLHyfKL1LtXnWRwl+GcOLp
RQbhsUWeT8Ot/S/AkA8/Tfh8e2QnmoQFbUxvIIhVl+FpxLJS91dA9tzGI4CfP/aH
WMf+Hny+buZ27Z4BDmEqhRkd2u+kNTkVA9LtnlhFrrNFIfc/Pl+HaqykhIJOKmF+
ji6suhwMmHwTrBA1YQLW9cnz3FsRVMqpHiN0wewamtioWoSQ9w4D0kazBPAZhQvB
6haeTrFk0GKBhuUU646NxmJA7dORRovrSNVCISb1zwwrKLrvFFeHfLnkcnnSRkSP
K71RDyFrWk+C9zXc6BBJ7n2EgJPUqFzOehoRl1HIFk3ZZlWGDPqWDZyr/hvHwpb/
yzMwS7CKgjmPmm3DgwkSEWqBJ9KXm+kkOwoXOWeeqV+qBgfEADtvpnbKwL+Jf2/a
ITp1pWnnNKmxXCQZ4jAJNgQ4eEOlAe38ysqxQGC1i7DeJAi2Q13NzsMjOwzRJE0s
UFqoWfQT9eVC5rE+/46DQrWVh6XxbSFk5Z8Qotv+G4mt1tUlmLr6kIVyNDjWGElV
wdsFYwbcqC0VFG1kMAOoDuM1JFUQRSpNipbwZBVSoQva1lSI4N81qbl6gs5MNdlB
YRyhlk/arCW2giGpf70YM8q8m6czEEj1IYw+O0+zXgUtvovTkwUEZNgvKaPk0X8L
xe5ADgtALYzKZC2wIe8DCc3cx2b5rCBLQeAyBfjDXMryoZJW7WoASpjZPXkFQmdd
ZjJYTQXmOB/gAYvwKH7HjVOIJN88hv8VLRlW6jyhpZgIPblwaMKCef5FaI+BZFDP
0+vB0zPHOkiS3wiq6MmBybyy3GAfozmtler5lbd4jgMGF/7lodOj8qRRkbDZ9sJK
wdtMNEVooGveIcsFEXksOdvLyCNVI+i0ZLyDZNU4uatFDUbknr7JwF2zQjrAHn7Z
Qh8SagzrGHofE27EVuYBSk4VeBL2P6Y6jU51SvF+xNFdq0nK+ssN5wLJ1bcseYHl
P0KPMBopMF5oh3/sybVeyn9RfP2YZjo9veZhSfrFRoKm2PRRDdiV2rWjcZ/eGZev
ymmYSJYfJfhROQMqMDpyxPcL23unDHOjsUPuxAJDYh0i2pY7vomapPPsiHj7vauc
t3J7As17AaNSjjg6aR1NyMsbk+p4XAGRtGneehFGhx6tL7CuGXtlja06dcYchxA5
udV1LckMSBHZi2UgMRYKyqqqwfiiGik+hu3S9AhLXqgaW1YbShME4VK8Wxh5znVj
iq5MUbR31IW7avhfcAgU2Of82kZs4BfLYrDUQjkcwfdkldoKvKA7s0QvZ6EQ0gU7
+ykRZoTmTI9aNa8YBspNJN5Wpo/KPIiuQPXmSBi4N7rsj25JawBnbu6Bm330ANGn
pKcuSIf0jYsW6U5yHNMsVK+4QQQCmSPo9uAfmLS2lmt164YCmR53tH+8PwcxfxTI
KQQHC49uCjbRgE3+zf2OyBkl7jpOz0I1XFzUda6jqRTYgFyjQXYcG/LZxvKWU5Fg
KWz+EuMpgN+Q6h0ve/6OMclZ/VNCwJu8khmn8S9YZdEvkdJe81tohA2Dek6qnQvw
wAy/NTIR65BlIlXJHhL68IeK8KbqF5I8ZkEnlVfzXu6fvmskllsVqDW9WK63YeTh
HfSCeraKKE4qg4YT0ZdWQUdg0OnmJ0+is7ZxfUl3bNAEj2e8VJ25szZ8Yciwy6aV
2FgD6L4pYY3wwxI1u6G651T9F7nL/43lajN6y8wtasIq9blBUpXCGntBSdUbBc7P
fnI/OslpnrEJpzCTwSCpmGiGIMDB6q0WjKiQ35/UHUK4TRNy4YcCrv2jsNVJ4r2f
8lJdu5BcZp3gwBMGpjdFwS84hssPo5WfTFW5iVkbaiPb1neJHH05527f5fKUA5T0
O8hxkhPJbCXtEFuPnBjFMCde/YBS3M7yN5Ws2MZtc3E/p2L+q1dCGilqIVGbRGmZ
tpypCqwVIKdQjtVTsmu/IEVmtBWkVO1X481B7r78gTcCz46h84b0eIK8gKc2mOP6
sZY+SoaC3h38lDx8oDACArDLDkVxDcO27EcMaDe/C/0CMhKzAqjnd5w/YtMPvGle
4pe1h4Vev8NtVyL+i4heyVgwUeVTqih11pUIkqnWQWMNU/R2Am84u9zeDE2y9KAs
RB8oWYdHQMGYbp50Le8zaARVbrxMJ3LjOjclbOxA6cAKaALH/ExrqWmWgxs5V4rj
sBW3M7tR4bwTcvDbg4kIpVtQy+7GnLhJDvS49QKpatLt2i2HndLXPWa3U/+jjuI0
RMueXH+fiCrk0KW7ciMaokAPVuSjdfnTzBwVsQSsx7shwIilaqb3utFZzdcxsfSB
I3uliKxRlAqVghzFmNsReA1LElwrgpiy/OSkH38AAns8VPDdLrR8qfzdCX5fCLYb
C/9FPnQ/BSVuuLvjiKph/A4lvgqX38qw8pMlObhjG7R4VFdLHuBj64HALl9oOAiC
oRfg3eDcyf0Zy0KuOdPmSMu715SKjMzE5tZXa0MqbmB9Bh1bERE/m8kaOAVmypwj
l0VTij9GEgl2CQL7BOULjgXdKdhEZ7hrK9pJMtTvAmphEWaLWAnruISThyG/RRkn
1zmMcz1SdGNBq6ETEJD8wO6pxXAkofwroEBmcEYId8ju9no6VMegQ668DSBy+8gv
EfOsXGoTCOtYBoiPYdjypr6MtGSbDZGHwdT19gVFTFuQoInJikfdFU7M95uu8Xz9
XgGGOrNrcz8I0zFWAXFLVnQRCJD0Gsy4uBrHOv9BbDRl1UrtljbXBeSdnvo+46Fy
6rA+egT4EUhrG/WzdJrOAHiEbsM58ELnliFTp6oeNu48wg/l3I+X5JLqDog8Whp4
ApWY58/3ijbkSk00UOTdohuHtsL6RR0z13P1wSR2VGUpU5TFJzSpx41+PnhvP09q
TZGkl4qQ27PZDWyQuTDerUvDszVQ5FH6FuKhOHck9929TUFNd+o8WnSqPW22RS+u
wAgBXyOUlFm24VQu2a+yzykNVVZoXeUjckmDLhsFsZdyuZw01wKF4bS0t6UWGYd5
OFt5dK9dia6lZ+qPhaBZu4TEoizXVPq+6Ua3HHY8NRyc1j8oa36J1D5CLzluQ9IQ
f8v00CJtceiZXI3+4u3rOto+1RgnLtRJHnjdB5jVathzEkDwgsyWIrhw+YzlcB3D
iXlb5gjRAfFYCc3XiaJNARnG2jIGYS9Z51a3OgjCc3sIU6Y54jioQTxsqIp+LpTr
6OEfQUBej7EOGZhIw8xt9TweOTzXoiKKAYLBLr/jEhfJxQI8oD0pwEb5lL9ViUX3
SkrWZjXDuaZYAzkqgIPv4e6GHCFpwh+/8p8UYYMqIxAue+UcYStLE1yaUlvHcedc
YUKM576nVM8Kz8wOwZ2a6/qROKgDi0jDlr4JJl2Hb/pUFcsoKFrx5Hzy4WnwsL5Z
bmtpStsB46ujPH3bkDaqGmm0B+VbINw29L3UzPE0NMu4D2Zz/N13Fdt4iVzZL9/5
JBYnidchIrfJssHz74hVShdeGjrWGGiU9ZFtdfSKT6iXykLz6SGSe+6wdDLBd+Sx
pHhA6N+itN1X9VR1iDqPdf3U/mf+3hvsksR/s8x7qkqTN0tXbKIVk3ErJAyLZdkn
RFsGvaqy0gn6VOB5qxBA2Q2ZIgQO2nTe4YQ2/siLtoPViRuh8e9YhWdhV8HMSb7D
bmfmBfkevLCcy380LQFN20lyyFpcIY2BGVv0DF3DXda2h3zgf7T3TcaFQ5nezZRE
v6DGN83INJApWqGEJCaEufhEu8Xr0jWjzWqTWDJFQG1fqBSaGO5wR1uTph5AYc78
zNWdSjcLWMo+uQonYofxsXxxQ1lK42CWsAXQC1/bVqNRrKN3s8FXXKvt6rNZXMVd
WgIqwQEadNpxbXaICLbE0F380i3H5Ce5N8IYvbDZoRR3K5tvLv5WM/PG8dlDdX2m
9yQZVBMtAp2aAmp2HCTNSyjE4fNv5QaLn/BnyJn8cBKIXgFMlH5ytn1++igx0r7e
6vxVuZh9p+Zr/48GYd+Se8skNKE+QJLcyQgj0fVEMjRgfx2onilbNjCGyyqHTrqv
9piWb/6QZsrtt+PQ6W2McmmQwONv9j2bZV1tFK5IK83JAwgD1W0yNouqjzNumDnM
m2TaePcuBGUFS0H52dtu7i8kFCVxtoePnbpwn+TaM55v50nIZ703XkKhyQBR68C/
2t4jerwIG0J5zWTh5kd8bNVUGpxzzUNYafQLIHyP9zdwwFHA2X8MGtcUuzsDaHWQ
idcB5M8lQsubDO1NkYnRZVUgh8EeALz81M/W6/V+/ZGqQyOCz1OwnQr7eLjIhr7O
d7x6HYc635wDiUZEQ4SOWfA/ky/ABkDynYM3C3xhWTGc9kwmfNQrsVf2MjWwe3qB
B/JkgRwNS7S9vXOcQE+w//6QmsRvebbFXnLTqj3/NG4CLvKg5f3qqHgLFtLKaMv7
N/Wfv02bA8e8KA6G+As3Vi3tZSTww7VfFvVyqDTAYemLmLj404sARtvuG7tz3gyj
H3wVmu3YwVS0TgyT1w5EfinrKd9Xu9iPUOinIqU7rJfKcp5p+fsX6f/ga+uCOkj8
Prk6mAxAIOWsH39hech8/0KryGNk04/BptuAQaJUUxDBxAzUSi00iImRjVfIILun
FlRrYWEYo43ZDwimtzH6G/zY3NugoPttRvPdyUjCfsmeoDNCR8LuFfBntDAmGK+B
PXpMp0KWb8Sm8x7/k+BtlPvHrp6cQxXfMFQTCZsSBn2VpO3BLeoMLt1jdtth6nHd
33d9mjGw7e9Zww4Ef1j1VNx4ITWWjjXMJCsh91oXbawYwXyKw0nUxh5oTUYdefdh
VYgftxyMO/7R6hDcWlpVWwj/1n+Y2VlD7IhRFbrXLJ+VEkA+yFZ70AodF/A56By9
HwioqXbaKM/dDYVw0TubV7UuTmoVCuvyr+Kjow/+Hp8K8WDa6KFPXPjBT95Nqxb8
9iJgaq/4mTymHid2UQ0weKKyeWgoceTOVYnnkab/yyXdRBMtPcJUN9CnwuKFPPFP
hOuU02Ey/keWH2MRhx46KFRmPc4q+1IyVgcnbuVG9Ow2BdBQ0EAroxIN0yGo9uUE
20+I1K0QZee1l5wWNbYbmKlC1vYTnRWzM8FUaCl7Ctl+TxOcyEfv+UiYAuZQVeRj
4Pe/TqJv102kzkN7jNQd9AU31iji985I7PNmr68loGVnZxFh8APZP/F9UxUmfepO
aLCJakuAYh/H+pgF01aeinEepzAVH/RlcYpZQfyBTbAUyBr4P+RBGnSYRwbXp1ce
+1OKtO/93dnjhWaOn2OmPN/gFuA6Q0Nf+72J/HWgMOumfgAxa6smxvwWzDvdlMd5
KA3I1Jq74EdS+cny/okhl94j5aBnPjRwrTyQz5ptnNWqlZJW9ITCpkp944sMDuRs
DgRZyFsdq9D/rdz5jEsqKuMPLzRB9ZwtRl/N/sB5c4ilg6cSft5+iGJw78/3JixE
YosiPtsvrxdKknik8jmNGxacQ2oQokEGNS3pRXZ3rOSujVavwXsKmnPUzLLrbRqI
4+nEuBwv9SEtHHZlgP9GfJORXnXjXkjphC0Z8vLpPhKd7E82sWKVhzRW2KWiBBeF
3IEuT2BH3IZF+hI2oZVSgkGsQyvQ7MqH+fxK5Cn3ASqX50deeKnmEm8F5gD1XRi1
XJKCoK/hGEVOpEjs8uzeAvHfnbWRDzrSuoYTu3A9/1LqvEwh+i76f1qlGvTnxLQP
tn/EXrHLHi5KM46oM8w2f6pfC9nUBYFJkC/4cCSZzauxCAmK2fO4b4hJO7FX6EhQ
OmkmSwWcKJHMmKmeYBbhNIkhOhtBkI2w+ilB7r6H94Sz3ZivneRX+cidhqEp+tHQ
DpydJBv7q4boo++YJwyxutptoUtS/syavw6irzDnImYYEC7ChTPNAp2r8A2kdSta
TUO6qho+mel0Bx6ImzwndVi8lHqGfQ+Z18JZkp5lJ37uX1g6h8ICANOoJM46PSXz
P/PWatY84HIOUUKtxNU87sLyVP8z5Mkc2EN+eNXiUjDE0KDcfXOIKmq2dGVcuW0z
otZ/t2GL7FaSc/oH3mp2Cfq4hlGr+DNixHe1ksN8OPyRyF+Znl91AWqGTOfwnO8Z
om4x+Sa+KDjcv93rzMsHrtJ8aQGuI7WY6tAZ+SCGVQHdMkD9uibkDqCmU6WJ53oG
2HX1GlgA1eU3RiMGKg/rJRZn69R1tZlTz2gefKju34gOKfxRQ+6nO+Zc+XBcj2U8
D4o6AQossJQkaUBw1xRD3pxQw0LnvhkPvbUwNDeGtpQ26uYzc4/Nds0jEiwY7PSq
vNUGySacBY53tc7bJVBznE9CellISjkb/oGTIsvFF6XAyKzKnVN7lzmFvgtN2Hnd
D2M5TR0ZVXr3XyMDBHZ/KOCFvaw6ClANivw0tOxIsR2UeVBCQjcvSpKAaGvPKXHj
DW0VSbtqzZEDb7AD45WdbnIsSxdL2CyjM8LHrr4nV4qb5LgMQFz10hanNV694rmi
KMrJ6wBe9hRVeYA91sJJiGfcjvr93AuFfn9FO/KahExjli/ABocjtFWxT4fcTUyW
2TdLlYa00tFm6UdkYyTTLpX5pyuYA+YmrYuuOWmiwDc2A//UmmaI3WATnKQZzctz
umrgThBarWs82V5e79ClKiFUdGlkbVx7f9bgx339BiGfUeC9wo/ZEt42ysCvvJ2Z
yvSRGFqIIXTmYACVP34kkGEc93v2dIK/dPgaw4X+KJu9yoAK49C23m6zTuT/uNFe
lVxDyHrtv7vyVpDny7isSg5uQe1y0pzu7Vybd3mWXC7XXozSNRPDXbfWEYpLD1rP
/GPDwj0QTDxCBiZMAtg/PwJmI/GcO1XqFEwb8mV45g9Ji45wgFhKxx8ISHbmNQ3p
P3lQtm3DvwVhjfG9aejiZns/G+SiVBQGwgwsYlFgzbZHX1sz94rniCFbXBnnMtWL
xH+WwXAoe4FTy4hEKojROvNduNGxzMB8d+CEshA/Q87LOG8eS/igQBSRiP+IbBG1
L7qs3Q75MyZ2ghvWALDSuvMloVTZ+uiQZtBlAUfLI+vGBkJzdvnzrJYWG/e9YLo+
bcmAfq6bx2sYBX5OOkacka930C4Q34KxIB4736EWntBwDJon/1yDFoIwEqT7DRaB
x8a3d/g2UVL9rFiyLToL/mEroKnuJC6ytIkl/Yscbh7ThdFhaKIxRDtoiMvpkkiv
YGzeRJwRq0kLQklxDYtt2v8c5lGru0lrMV5CeiizgDOMpml8lZBjCLaiMfk1A65H
fJfn4tWUhoJu2rgh1zXbhzHbj3533zuJhZtUCDOOpMypKhYPyFPcFiaBPmYMeEvH
w0t56aG/mUsxWfRZZlNwJpiizu3k4igfZ/SajtEq0DXpNr3tT32w/w5H6pEhknGD
pZlBSUZN0eXALA0XCMjutHpyp+8u+O24geokrPKpAREzHYS1dmLxyzmPV38yZwqC
m1rDM4mmgInn0Id0P6he+d5sJL2ZZf1GPD7OqscmShhbGvvEM/KHLvyY1eX0hcsI
+qRzPmbDM54n3fRi0FOziRNjSD+5KQtMKhzHAqcQEr6ffxkMd8ITt+R0dyRel3rI
pzNi+K4pOX73LCtuQgFS68FKqTKsFzAfkHtzk/8rkjdP/KSE1M2vBa7heGeXs8S2
eQhfpm8m63trJ2OGk3E3TU03TCbh0esjwMKhJFrk7kIpVtChELYKKnl+kszuWvZI
hvbkOgh0zFwEkn4+B3hKY0O4k7Csikypp9/HSsTq8X+KVTAInquv99MX+CWkfsGT
nLfn0r00r8zxd9eIDuki6WYQmzZNT4R9LELx2AJcO9+O9gln+Wn4q3/ap+GYTLt5
PofsUlMkyOdNMTMnqH0/pmlr1iTK19WOgR+cSSLlsiiZ2kEPyGjzxtWgZkBzX62g
v/JY8pfNDp7+jzRUCbh2MhFBzObqPkkV3WwemPxOu7eMbyl9neu6eDTkq7zjZbfW
iHShlJUOPCHqEkwI1Q803CVYHACS3gJiq5kh81UfW8opOh/iEj8NjKLvND3uqWQl
P7/0ttTigZlZejpUmog7VWXMbaZ5RJQRuDxgV/xO453akjbc+JMkZGex32CUGj2v
LPvW2fbHElpBZT1092jhvklHoANW8HhbP6txWW/JaB7Y6o5Z7m4pvgwvzWnq8uhp
M5hB937abT/tjbgG1lgqBU4WbvJ30J+7J5VyzZVtrepg9P2mQvlmg7pzUQZVjMF4
9BsyRUFMFMGD4VRkxMjWwcM5HDVKK8P1DoGL+p1c+8X/ppq1wh2Koxwc3JH5Qb2z
N8CD/8qhKuopRGEhP4EHcR7RX1XwHCRtaTG5MFhzEopXPVUqy793nKvzKxhZwZAe
641lf40NY12kV0u/OXyV6jV7vFV2WMvrLGFWXI3TLnewc3KIm5y7zebFByyHx2QS
zxkmrRq5mYX3EKRF9blKZakPW6iuIzrjXzefyG4JnWtHlqXVmPdrWTyivQrt5lhg
W4CL0deT8VIy9YHatKTqvboomae4mIqlbvmUN5fi15b8SqU/ykYsnedFcaBppSi4
2Av3WAz2VAZq9RelRiEq7SJmhim4zaWUB7vKG2Qu57robJiz194QK1IiUEQL8rts
97nTMPGPaoc78Pu6Pc3Fq17Q57YJJqVn2ZJNPxUmjsFFUZ659qHiWh9B+1Crkpdf
R+ZSX71/kiuYbf/CMQzuIZDiZKIo4dsFS/JLhn5C7Fioo7NuGeVC+jJ9qI1xDF4b
YA6gNfV7Uu4plZa78u1d0no29nLdilhDXqKUNl+yddpLbnO3MfILvuNALoyCLXq7
qJEPruVmriMYnv3FJZ5eHDVyy8e3vm4iw3JDoWp5Y2XwoHhZBMi4MGAk3dpay7Gu
SP1cXjKOfFqbQ31c22yByZLYI3icv9bMWlehWX0EWRCgphECzLLKtzz0fMuznNHg
af6ABrv+UJFNAd4iz33YoBc+i1eLQ7Bl4Vjs3VQwi3mp9HSbOmF0OUpWDD+enWHv
HGQPDphp6N/Cfd2Esko72TBSd88hxBsNL5vGiBuo2OF8g1W1LOk0Hujs5HzmH4Id
M25s8brGoNetY/xp2elHFri6xkc9nDy6nLUn0xWlybhMiyBJO51JyqPhifiqITEr
/wUCcHcvYRIutZz6e/8t56jQbxo4sqmvk7PelksCBvu3uTBLiMJ33Z+vClbh4/Bg
m1zHezpiLiYydWlkiPjcNTWVye/rFzbkDw3yL+rJRQwdB+q8nCBaHQ/bjmMPlnQN
+pPV+ztAZRsbP0u6HE6PzhsquXLA9MZb66j9AQ8eByoRBRVa8SfOghCiIZrIZkZF
8URKIUYkAdnsS/s0L5iz5C62qbiG0JxEGl8l7SAL6i85nRScu/0uL86nGIBhykmj
exao148xgiPEZKoIX3E1UFcQaQ5vmPtrtn8HINz4fbMRdghtbC/8++K2Ye69j776
pVThRNCyJywEdcU0kX/RclSrkTEVPAUBK2imkllzTeM/eYLCHFIh8WO8m7jMAt+2
pqhAJfmrLF9YEbsHOR92T1yLCzcTddoiOpmZYJcRi7MGZCDBNjYgl85Frdi9HZja
PRHJrmIBDaHs7PfGyWcdlnMYCVSL6k/5jqcPXxeE2elDQqqEKh/zcchYbiyD8wa3
MRvLtUizgssYs3rGAmCtyO6EIXGPn3Tif2KEyduBGM5Hbs0/dWrpvLVUwum0TshR
vv4ro+9ju6Cf4EdplkGF956O+BurTu9kOvJG42uTgck4PTeJrzbpxuetgEO8e4qP
plnVVfGLBFkMozx0pO3kpQ2KQMFDVMyWLlo/vkBUMqCqn0kkPtsa/XKanZ8BAgVd
IvJXxQUznXbwZdd4HAsmLPax0KV4FA+SumN+uxO9ObEaB21Fs6fr4kxXs38cl4ti
h/D7RWXdLOcqcXW7VTDtfJVKHlHsE5a3LBJg+P1OE/fLHMoMsrlR7/CCijDsQ6zg
zJSuwzJGplSL42IO0F0ZNIbgevki1H4mc584v7nurjTg/jxJp9Slv2FmXsey/1AY
G9XE5M1uOsKqAnJzu6Vrz+tv6lx3ra+hwoQChmPqtyDTSpdwEv64G3KupSuUGiCe
UoStZ56r1H619DZBWi+j6TfP2oUQ2tX9+mk7ogwldd5g8bgJxi1oKrjrd6wAzySX
SFoXb4fs2B44a8OT4VIMK5IB6lpnmTZh2nVj8es+w3XaUyi+HXOd4cVJ4SNNoaY5
T/GCTSml/eoRjkXKIbVKdjaWhzb2nOHK3VWSKWtiAiYt/OiNan2X9NLgZxQO/vWL
AUhfrHjMGudWek+no9kHefU6po1ovPBh+PddbXuwBuYUztwozHvAuy6v2a/R1mwj
IALRXJoKqnUV0GZItDhHDStNI2lcSJml4WGHUk5jQmIoDFQJ0ivkkrAjnzBzVme5
hdEXN8y9jeAux1i1CFtdgeI0QEZ7X/HpiEOJGR9GpB4WVdWxaoNvtQj0WeUw1pHz
oPfPsgHVZ6v+tsnJTe0ebH1+HFdii0P12j3X+0z8/YO0Lk20pphbnvIIQ0GqhZtG
omw8vgi6WrpzlYeACyLtjTAVIGO57zxcuV9cCqUaC2NTHaK80GoAAjm2/zVuf4W4
5ZUk+7b5Ktu8SG0dVa1bk4AAGKBy7JQRPfZwNtYG3yJQ/0BCysa8O+6sBlSr4h7Q
8Qam2DF80doZOe+DF/za6b5tq/lKDYwJVK9tj6Wk+6AMdPe6SbRmD2JmvV8Jr5Ab
IZ9FsDPmrvkReya9Ghs25sl8rkMtYftXnY+k3A58vNg0iNSEvtFLdhtrsqY+piFE
mYNGWjQw/1ur/9MbnlsUMZKLOLQLmKM+BI64paKemf2wTppsqnVze6o1kQ27cs8h
78CVVht/lGOpX53cwrnZqHq/TxDh0VnIxwNZ8fW3bXzvcbuup3f7kC4k4Bqaz87J
olZg43xrQvtmJHK1IqjUSdPF05x64i7TixRVXjEtzBOg+64CBabUX+lIh10KK3y2
3W7wNdrFzfMevyYvbbtaTKBLb5XB0KPkkc9hnIgRpP14VIHYxTTvFbE81cOLmPRL
97azp2AiWdl5vkcq4a3+JrWFCIpcdaaqaIMyZdEK6Ski+SMut14qo+aBW+e84rhO
oYrCbS+CLHWDsrDqNou+tSs8qx9Zp4GpLbLruqJTihP3QwLuUljPquM6zljKWVzu
aOUNGP8Czlco5Pvp3akjdYoTV12hgFZ9zs+AK6ZroQQjgIC8OFtM7kNcXYscaeQr
nwbAXEJkKeQbb3+us/8GyFQsn/DMOohQ6WDkpH2d+KNyPsVG50gQ6YZmf/LhFZ7e
cqduYY6ycm6/0jOJnBlI2oxd4SwKAu5tTFnD2TmdyyjLT0QcIyQwEUFbjuz2clHs
YBN9PsEx0uP4/FHHGZ1RewK5GlIHRHbwU06P+NHYcefT3i69NW2RzaG1r6vIhMrq
lhzkhmxddX6TwbwW4LhUO9czE5brYnlcZIAzFsXQkBrsLT22fCfwRkaxzwgnmLrw
doSrl8AAiQ4jghli4+Ntgna49GWSaO2foFjvUJYLmZv4HPRxyEpwAA6NDPuAjyUn
kjmrwiZSo9yPsSHTdvudCEgXcaopGHcdas2/nXAXBKlADyd2Uigl/nC6cqytVDHk
iID6Vba4+7cohTUZzIR1VZ956R/VpsCHZdWHtPhTleeFJcPvHy2rZvJB/+2u7n6G
FlJSv3KeyROU0WCJ7VK2oC1HdNKTsTa8NqjvBnlGy+s=
`pragma protect end_protected
