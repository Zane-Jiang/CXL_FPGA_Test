// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
PrKhR4c9Q2PuEPBsDyiHwyY36FOXwU5pijTM4SuDCJKKHCaAIqZDA9zNLYmY/EfH
GQr1e9A9VCHS+nk03f3gs8Xkls0m0nwBBdHnaU0HUyKVfwB1hVPrv6QdCpSGhcnJ
oJU4/4nsJyI2dbFpKDv9qh2PY+zULeQ2SU8UKVBoWBNC1g8G7CLwEw==
//pragma protect end_key_block
//pragma protect digest_block
NncTQZBTsQLiTB0VvbDhqCtzsJs=
//pragma protect end_digest_block
//pragma protect data_block
guG4Z8d+t3xlyvXsMuDT46zYKDZ9TMlqcbcGo/xjwzDyeCu0Bv/JkahZg589hzwa
DRhVaYFldT5Y+hszYzbxJWjoyRpsVxcBX0j6pK3aOm0dhpCL/Cb/rWnYvOURph86
YkfdWa/zyptMHtQ3r6jOEQ0SR7kP0GHxxWubIUuVjLpdqyEJMT/VGwH7VgNk3Qwn
YufiwSsoOCDgos/wawPW4L17xkEqlgEJNDfa7U/oT2wxKLQzB9/0c9KglOVDqPLO
B1gdOnZeJJYSAy5UB1lY8lVbRpkJ9axYI1KjfqnLUGwixZkwNNK6vg3DNO5XRO5p
/jtTnRkUaQETzUU00f1HnhU6udrJR2U/z3/OkmDn2l4v+dSLUrdGnYmANPIV3WX7
O3jNjtNlZEgqd9Vb8oKdrH6owNztpz3ENR9rmYfm+xpCrC7ijgiycMneO/6nhLwH
kb5GYBvJmSNkdYr4wAiUtmvLVb47QWsE9xmBkr5xTZx9/56MLmwSebVDV+Z9t2Oy
BZex8ARw7V0XHMTGHU7ZLEIt0C9d7D/rRkhHmLEMI7U3+ANEH/tJ56tT9icC6opV
1RG2uAyhO/HJ5QsS0PBXsKDWcqsX5lnjRU1dwzJjgqpJ872MmHmm/DEzc+u7iJzt
rWf9FJO9MHd0ZqQNBD2ZVAS8HElMaITzeI71yENvKjT2tw8nXbZd8OeCIKbbP5BD
/du4V9bpfnBTu5cM1kxUAIN8NauPkaGFPNIC7p/XZmTxji6TpLKX1IgKv3lmGpmf
BqdbGrDxW42qHe+wveGZe2So5nynW6Cc0ygLpnexuUwj63GssQ+IHnZVkA6kF+QM
G3Px/4vWfOPv9IfmJj7/S3ua0V+WO3I98uK5CkhTtNXH+1uEE1XCLdRSiZHPxnt9
NZlPVdNYIwBC6/VDaGazDI4ewfWmQKpP02zYbctHhyl12yA2K4NuuuYE/2+cQ/B0
mq9CFToFr3ySTA35cPoMMnnOH2FPltW2J8gF+Hwr9uSGuSwTL3sXmjfpeF4KM6xW
x5YGXexon1r1MbX9kJW3OulJfQM5pnA3NIAThBlfA/uDtVbbcdOMJrxCDFyhCp9T
R4IeL2Ysc9/m1nzURMDytLpsJlkoDbJrcvM2nBpSCRhTgfuP41TCpU/TW1eERU2I
hfypqEe8sZJFssF60be9jKzOWf5kSdbTxwMW5V9mbcv4ypH4VaPWKVZsxyaY7aap
QELAkDkccl82u3i5/G2ioMZz+Pm77EycNL+VI/oOkqTYb/zSFvfpI8cpO9ABV8IJ
m1oqkC1piw9yclDM8xPtfJQ0dnv75uIKorIYt+uJhPuOvvsL53jCPGJ6/SQTvexr
7OFHtRKkyT/zt6696JMXXN8apOD5Tq+8PrQuVUGAwNVoVYhgkMxHuM5dHtKh4IfB
5WJp65aYjWAL+eN1vmKEL3Fqr2hh1DlPiBzAArraZ/6Z3DhAhUeIl7Q+DrQ3kcQT
hg4afpjYElg52sFtsKF623w81paottgIKTyRIYrMpxS6JscTIGOXAzPzS26nPzxt
UbccdH9vUOaZ4JE+sVx1hcGu4qm8Df5SAy6hLB6z027Tx79D4doRQUOIxXuhXXuM
m/S6eAs++WzbPGKRXRd3DCPmi6HpZekIzsve7WVP8PjNk/mqf6QJDXbAZaTD3dXB
mWra9QLsR7U2zMDzIWy4gppv+uJf1YFaA2az53MpHJ/gWq7elmxCfU2tt+5U8tOo
sEGAGxM39GYf7+l90bMjglPMQWxxW3WyXsyWQlPJvwoMOUBtfs4xUHY540o82FA0
b4fLm1T0b57RJrjctW/OW7WDDA78bjXAkB8MTcdfXAlK2xHH9nVxnjaw5NOyIzMO
04bdywacW2oL6aIc/kcooxS788vDGpcikiE+6lsaAHCysaQI0xdtbYEzIfISeUmZ
i//fDKlB6zeOChKcAy5Rmt33QgEBVCNUdsQHHi5J/TTikZQBiMBqKRh5kQp/WceJ
RXs1w6TFxUbbLQM62rUk9VEFTT/QFsOzBBx1PM5My8IOw0WhNqGkaDWm4kqdX1Zk
jQVtMY4tC6KQvhhN0szm8svETo69XF3Zr/+8oh0TUfX70zIP8WKox469rW64LlCm
BdI6EpRv3IjGig5nQVhfM3YzDGMrJ9BB3x5mUdflqUM9wsVy3skGRmk3yw5PmPpy
VDPDutYSMFFH6YkVJwtmh589/L69iWTSwSljapYc6SO187oLp1bXmSAyLlOQ0j1D
P/kmGguHQ/KkVQnsLMV93anoXPZfA1c0myOvZlRzafkFTVVl2w2RQlxbd8fdVNOV
mXoKi23Wbv1UepfSJawd7jF/9FGPhJIoPXOv0wBe43nWeh3a08+7DvwV+YphDbdl
eGTe1+gpjdK50Bpq+hFqLyV3bwzXIqpCLP4IhSaj5gkAwfLxc0aGHOYVWopAJhNz
4enjMm7SMh0oCJSPaWimLMjQKdPqe0sNIW3losujOFtNHW3MiLO44Mcp7f58Y7K9
zLz8VX8l1mbcjVRamkT9+OieD3ASRlGRc327WFFrt0BGk6OBDKyCVzNndxoS73rQ
L9hcPT0gK+sltq/BTsZ7gECqT5aTC3OdYQdYCddQe/MX/iA/MW4fBPnf5ma5mqE2
B1QEagTq3ARxVvh0Y9lbVDOv5vLJnZg6sndAxUQdXMzwXXx9OR3gP/aHUzxRA0/J
DRZyX7/U2eh1oTI2oPCYbhUCq3WCVFCgKFkEN1Miaww1MyZvhxuVopV26S5JAehB
Ebo0k8OHJdvl6cihBLBZZbPFdP07D2YcuF9CWTuVzffQvCo2IGHHxRG6PiPgDs8y
ljI9cLOY3me2IUMfvRATwelHdz2/SEeeKDWRyBBiWDyb2zCSbwaqQydJGL/OgRCF
Ot1+WtHGo1U7BbsKrmO0kbsZ/1lqh3USy/zBD4AVCTDEmND2aYqrEpaeygSagszJ
vKL097QEWT1xzxBPmStKcLEDX2KG2piZgud2sGLZQgNHnFZw5fexzS/5aWAaGZWT
7XLAOzqETF+Bu0Ej96ATfDLK7fXmLDAYvKsf2isqxNOioPnpDaV3n9yjNDHbJJ/L
muu/fCJM3TpXOQT4diQuC7Z4XeYAgEZPo+PHDy5azFtLGTD/RuxuTKrekAxo58v5
UbjzyOTNmXOTHfMgsyqhA63LKAsyyUq9vTC/d8nzE+URYl3MJFEXlN8oK/wGJdOx
ADNO6Yq0kG2pp1bkMOKoRj8uQi0w+ewikMKqAMhTW+zBBrYb7n0JQiLRVv77nQvg
rd9nfdj4CC7A2CEt56qedhPrJugl/elpBT8BRDuLK2U9WrSP7ysTuKuu8w82sgAR
KGV+KwknAYDbm10fZFiICQ0ZZtk17qMKBXs0GdF98dXejvVmTOFh/s2i/VU8WOGY
cAcgIeBj7+jS09S6YEAV2sjq97aydWGVdH8JWEtB1TRrFp4H6Pkd/IidNpNaeX5G
sXSJFEKhQq0JSXBWvQs1/E2f+PshOdCW7URn9QdsziwnfUdFjvJBYnYTlIAQUvK+
Bv1mo6F3ovAesKZQDCBZ8N0e5+SuO+0TlDXfm5nZPAksQsEXS+ypYhmyUmSCbL/z
1dk7PXcrUO8q2W52BFtD01BfT+FdzkAP6CyKCDcT+NPT1lMAfSdUoKJGhqTAfxkA
HhgYaDr12ZUW9uT89XRYZxoUzRX+HfaFHtWa/uBngfnLNLSVaH4Kp5bDqowlYrOA
mj3KihY/5Y43NLUcgsYH3RBzWWeZCTe3PyQylizpJCEtStzCbPBU5c6ZA2XpOa2e
2aScs6qSdHEatgOqpwdNJXq5rC7MyI7PpZ9oJOaO0KivmdsUopnv4iTIpdIlxEvJ
EM2XkHjlmcrqiArgkGXZbe0K3hAnawWfGwPN/fjakKXVJK0JebNhBU8Rf1qE+Ogp
adYpLJ4a76O+Dwh7VuKvRP9R0H5g9hqn7ZUq3xLkXLoPAA81a5qPntxqKLivIIte
HKPxq64Wjt8sID1zdFT2xjQfOUolVR5cCngrchXKGdIRRGHPd26D+X0KSXu8prSH
6AJ8oZ2wAR9B1k1sjpY8W8JVq8cotiY1a5pwJwkpcS1vMzrhOBaYOsOI8sRI7tQv
K/WcU8Ow5CPxtbioiVh2EmLBc+TtMIyj6ycBXC5txWo6xCmQOdyTyVAGalZHjFf2
r55AKF1kaKqSssKkSVPlA1TfDU8YSECmAM5WDL5Cw9zUrW58McWxZIQ7MBTlp5CX
y9nTcnBnmqLJwqbkN0H1T6kM3NU6fx0gn70Cl1/0rdWSa6Z4WAnchPLQttMYAVWF
tSEY0I2Rdnte8kWrfD9Zqckt3HThf2gSWZo+tEllfXZa1UPDOYk9p5IEhPTpxWX9
YaylgRnr++3wcPZW0MqrOaT3TORHjd/TmvixjF6DF3USx+XlrUq7XlK0wDUQc2qK
iNbmdxEJ6nIhSW46jxdCVbRemgptw/9TZ6Tl5PiGzqy3GFO+joQl3u6nbDyGyvbY
7sBuTtyH3WSKSOOs/mP3viGCG1zjNiD9fylL+WL1wMVitMkpSUo1MZkAhkcngDeF
iBx5GJMc1QPuigDLu4jlKxNOSTmgzwnSu0cNN04xcPvAitA/hBJyPl3RXi7MIGOZ
lSHBqfeHzKSSPcEUwckFItBlWG/YkmPHvHonHUo7/CX+izUS6Kuh7+J8eW3SrI4s
zbe2eP92Z4/cWzjHvjGGVqRufdwZPxhBJXf/O+ilOAee+A48Yzv/urLF9Snpq5I8
LTxwuYtaXwjn3OcNkaR5Dm324PzN6k+y/gBSCO62+8CW9z2oFlMwQF/+hhtVpDYc
SDVuPUgkVqJ6Bx+shqBr2CFpr8RtHlU56sFXJBuwYy7h9ZlwE2Qa4ZhrZBTZ2PT4
QSM9m4GacP5JpoEprKZMtCVeuA18xzGLLjzSj8kWghU2oT54WCAiT2FJ2BSyNiEE
Ft+/LI+eUnAsIBHwnj+ycPiWZ43gIOTvUp+9mzx/LAML55run22y6tJp4I/6JYBP
oHLpia5zwVPNY/ax7d2ssq9LgRWyAC5DVK0X4Ml88sNZSs9zZeMykkA8VGm0Czs/
hYRY8Ap+2HzPdhmqzj68EK8K/g3+cyDMerZhOVPhlLrSFwMHng8ANmt7EHh5ahLs
skM0CsYaMEFrr5vxU72QQownJz2r2KJu0UMSJ452eqIcQ9ixD9uFnfkHEYnXsWUb
LYrBtjL02e2iUKiPv8eEme+0Kp9fg7e18fUUNqUk3+gDCrFj8ceviFg0yBYZdBh6
H6TGTforaHRHiUwX6HQYkm1jmTO/HP9z/S1VnPXw/hvXvDppRkX5VMlDqASJiPiJ
F7Mkb5mWWxkkaL0o7pj4bpd1od+aS2YrkXRywYvzyCpaXo98omvsC+dcUWeejNRt
192NOWmtkqk/sQZtZUjhB+FbWGWPX+SMdI3CIzahpajI/zzgqzORiaPNaWUSuWJ8
bg5MqAUz5FQlls0KZQzJIkrz2VPDHLGMMhvwxB+Rgi+GnucZQ36rdFv79U8Q4TpU
VLYfQMaY1K2J4v9ARBik3gNsyb1tQEyReytU+9hJ929A3dC+5HMajcTon3eLZV19
/nBeEif6v354PAVyZHvtFb0GBk39SviDMPE8YTLm+DItLgemuV2ryZ039pFYLFXU
6a0xbFOB0a2nBGyEwfkB4PRqx5Dvi6V6eiBHUIHtLDur/5Nh9yvADvAenI7QB2Mt
9kPyvjJlUNFpnuTRz6clXV2naHeJ3BVFsh2k7MJsjR2Yyc/XgYePl5YacRVJlJvb
m4Nol83pxFR68aG9mFi6z4B3SMsyTRMF32mS3oZQp2Tr1x4dviMPu0biPqcU0zC4
719n02wZIjapq0Xmm1A3NX2EytUD/F301OjaUFRKfLipvpn23IklmUjsJy9veooH
6n2HmdrY4ZHgThiS7laEnaSOpk76OHhymE8zVBeQ81F0KUaLfOQcrTIpquAkYcgE
QaqybBrfUxTm250O1sB6bEUWZqI3GBT/+1uwTTUdr6sU2l/ynjSSYHMVBS4SyDCn
ibVHXdoCV4qskJ+/Msabg/fblLigUEV8kZNjci0YMCHLCNeDE/OttFw7Vmf4WLM9
eVZYSf8/cmA2fhMBPs3/MfYk5pKcuvGi1rupCrDSBGvsXUAAOkUsYPAMCxco8h2O
nwnHYxT9jYNPYgQB2UTvgTil0ZTcQuRBj2eVfpYfGOuC44Qu7nMCnjXJmfmqYF0R
taCMvkPYuEjZCXLUsNQokhVP7LJaCMVi64UofxuxwoAHbQ31ZznpA6xt2TqJoZA7
lkeWDv758vmS3q1Dh/V+yA7xGPymNMCR0frNEFRbQmOG1pVVIlaZ2JWJ3/NcKFAm
/9DB/qwEHpb8btiwjg7Hz+dfAMypd35gJWS/ZiQM7/D3RycGHYcCdFDKFd3b7g1s
Rvj3pZh+LobE2QXrqR1vMlPpN43i0/IWM1MjTLZE9SU/isz5JHV4S+YlCBZyzlL2
i5b4b2KKk0GvFQiarbAKzAOgM7DRsJhz0ephvLRzhrvFhEtW6hgnJH9R76peVyeS
RTX6S+UVJVYHIdyPypKGK3fqxyRhOF+bxxcUY3u6ax3k+MdUBCyH/OjiXkQoLYEm
PuPNNVUI4VRohDEY3SMy3AG8cgrCrYdmY2oZnqYROFXmPBfFD7Ru/uCkQT48S4gg
/t+QqATHscKFJf5ky7vODA/2/Br9DDne1xCDr+XOmprW/LM/IawUeu5Q2hq96r1Z
vS/cAZMI2553lOpEvOa6pi2x3EX+emM59ALnzzks+cc8MZnM1eVQnUiv+yhWueRf
IiE0cbtLUV1MT+6+XLJVmBcuVAvSu0eexTQBj/m2zz/VIxrfUInOr/waJTHQoYW/
SKEXmZ1wwKR81LNvsb97ccMvzrn+oieX2FGPdAXD8we+YHq+WB8+vZ5NnGtrnEWL
YmxnA3CajmuAV+U74nS5RFwnLhq5jdgl2DFQShB/0Fo0COfHtnjU/zFUZHFfP5+H
OEExTerDsWLnISpUgDeBP5+J+/pC/l2X0L9HOOPQdIuNLO8ZkEUhm4X9GedYZfgY
wPKMYunuzYg55BpqjrdazCM+9nlMWElwvHAuzksgtIwxRSKnSO7JVA9Njh9aLar0
1t6sH9p0CocfwHGnsM8H+ZXwhi/Hn3+5wP4UTenD39lqjfr/PmuyJuol3aq6gVyj
TYdqsIgmz9MGOrnxUKQqSLqknk5OGZC9N8IrApm3NcU4VmINpxNA6ud8ntHkCDtO
xOiTawF7OYh1jgg++wHn2iFnd926Y048b+Q79PKQKOCKksC2rYCHmNGw4BkuBFkH
qMjN5CO/0PGOrCYF7EYK+2k27mUfcE4zksE/xCBV6Cw53iVrOYbSk+rZotG1rXSP
ZArHcE93P8JtCFp6Wsm9dJl+R1i828akRjNR/ZBZrkEatf+g/WvtplM8jkn+s4Ks
4rn1O648X//6gitBk6KiqlstIQzfVXWKA5NG88HNBDVGhslsdD8SfurfhnO52Kmy
F1qezBuwk5n6wGM5Y9UsDLTSLtHyD5jVELfIsZVdhuF/TKEOA8w2Tv7e6UGDzVPc
p/qj91gZ4aVheMVidrEERvcyNXg2HhU0+JOqam1c+608bHIg+kAJjFW4KBDBLnEA
qvlVD7uNoWGMyyzsPkr8IA8UBCfjuTM/5JoDhKNXenHz6Rl/APWBJKUuvJTZqg59
fmg+8O6jZtKJIp9HjecoPLfny9qH37q72gLed/D5MKWEtYq4ddo81xtwy+328Vqo
AAb5PpH1pjtzNqeAs56PDODgPkVB5Rjg3/31pyIIfZ9K7FSSnU3aESAN8+GhP/bq
SGkD3G1l4OdHw7kbsEJ/Tzd1HRG2xB/VjRGiD0N5RmyipThO1FdO4kB85YnTL9Vj
nUHPI2X2lXK5NpCc7JqTmxy7Tl2bmRj2eA//jBbFbjgsuwm2DVxuE872YKf7JoQL
bnRfqs7yq6AHAwhBAyXbhXghhP1WyTZOHdn0w2Mpb/efSKkFBjRAff7bXY2sScUc
sqKweC+Ie12PJxQEf6XXp/eVZLHFstW0kK1d4/p34Z5wSa46g33BMwQHkpr1jyOl
4spYwsvcMM3BNOZ0YeS871/3whsDYA3RZHYJGXO+2ELJUawjkUsqv/EGdr8htLsS
HrsAWTmuhugdVEVlmVQanCEx5ZOI7nikBrZJ/QpaX/2J5je7z13jDR90Y29YyOi6
DDoNPc1hHQYTBH3fWiGJr9hFGrX3RZhXEasyYuWeo9cHk3Kraawq4xIkkwUEAtl3
ratB+oHlP89TS3+Vy0cQhDe4vV08ZPgn97+FBDeD6Ui9LYFWtF08IHlHXx71xyOB
q7QkeZiCFd7Eje4gk4cQ8Zd52xU/XBBUmN0p5PX1A3kacjQICYWZ82I0jz8zdhQ/
y7iDRhZl2IFaNrgwq29R4QWRUChwoaHZVafbkaGvqJpVpF4ZTYNBsFCw8od+6JfG
gVTkUGhzH2ivUAnn0uV3byrWx3nMYeNksDV06xetNd21phSxELkp3fW0bUqnyWpO
5+YWa3eIYoWoYPn492br+SF3AvIceVBNx2FVLDPtCl6Kz1lQwWSLUP6Us0sLPAVO
fXw0LUkDJAhpWD4xLX1xtlUzbLFsBPKPSd/33iMZrFVr+kDwzO8tH0lF1qH3zzEA
C5L/OHjYbQ4z8RWSija+3n+SeeZHIALYDMEkyGei+668q08OUo3FwU/6nLdawxZQ
fqhU9qrrHP5ciaJgZWdWUhJqAiUTv01iJHQW6GjkjDdhjWzeIA3WrPCYEnJsRurE
FdEhvMXH7wQwC3h5ShVR9RKGxkDc9Z9SO4c+0hhjmY486nQoY/yW4KIXT4y0FKTF
wJ0vLcfwCjFdsa+cmyy9EfHr015jfPvKrtes3pHzRUOCFEOzZHb+AHGPWokl2TUy
1YtYCgqmGf5j4ugva0j5ELSDCjqDSgo89BN9rLuqQC12PtruT/BAw5PfY1KHSwaj
9/4lnxdLF1A8Mphs7rX7HMXXqT6QWvV2ZG8g2IGViY1nyaZrzmJSe997x51nf1g4
QG/J9aFS9+zva9j9Pxo2JMtEIn9CZCmnopwW1ird+UDlhMescLdG2tcjYSF6TkIA
RJeqTGFrTt0rBuJL8o+ecT91kVygkdmua2uafEGlcTuHQMSPDHjT/nj17gmn+n3X
7X5mX6g2fpqA6XTzRMoFTnV+Y0XOwNFSJ1kyF+LwX0OyNhVy2rD4xBTX3TVhR9ik
RWRIk4038+b+65Ud2wqAumG7XIR49Aqa6NwEs6R2tji26e1/kxu3ee8BU1rjqQZL
7KPGeAQ8PDVJ+Bpp0B84AkNWMjhQHKI1PINIAQ0gYSpkLO7uS6ac8OQ0RTFi+ObN
n9sOBFnO3NIkmJ6iR2mgXqLAooVCp0O9on1PyJfoT4nhNiIGbBIMB/wYhuwzpPx3
NdSGGCVHbNeJ1gU9dLfpe5ZZC7YEEUlHjOglWv+t1WT/MEcDQ8ayBrp9+JbddPI4
55h9hIRK/j5+eRr1Sf62vt7PS3juTzJh/0Db5CIaODlDrl5Y99smfjDlOcqAf0Em
TeGxM/sSGNOb+Nx+cKnr3NbKd1hela3D3hKh91+L+bzdDr6OoKjgB2yiwjww7ouu
A6cHYUA77pMdZULOK3IS51qwbCj6pC341226/YUzT1rwzrUvjCb7wViR5xADao3p
WNjI6eVsmJ5IAhDhX4YWbhiDF0RNtAiGiLz6v46uw0Q27CvL87yfxShE46vjq/Vu
n7kZ+UWcxv9GOtP4jSp7/1bh1jjtwbf2a2uj7dRCX+CG1Fvvk/5/TvEsUpGMoPpH
aFHuWIgjdKnWrAYVxuHgPV0qG1s9UdYG/qCtbZo+bsvYgNU6bZ4NDSEtiq8AM/CM
Zt7lEs3ublNyyJBuocitbr+POiF7pMDQUk5CGXyoEStWP0n7SDgE6TOMNTSrfuY0
WRSOOE+dSvo6RBFW49TomDEZCVESsN0fkdcxSvbglD1siA5RH+TCRhK0B3g6vP7K
Z2edcGMbGCR7H57mSYQEwrzqtU4ckZIkH0ohAR00NLwDmUF+wvpSokgi8qmP4/f1
Kz0s33RDsYpD1a7XWClhjyBQ2Bff2E+BfDAFfAmPzcZDvOh6Io2a+6w1UsQnHJ+1
+isLI4uPuudRgZCkZ9EQMc/ePip1EKlebt59lH8KHqhfBnbVA0qcwjhsypgxizYS
538XWdLxtp2eWbV+BEHC8fdR1O2zuXYfplEwwNTvO9/E8f7CyIJJ+cR00YVzXuNk
gvOT7QxpFu9gzSii1pqwFHFlJskoYOxphecREyBiuMwYIViZYypXbfZ/QWDcLEnZ
uBFumLk1tiTyDLCoqtYFJIEuoOrZOztgeryxM0As0xXJwnZJ717AQ7DvuymWhXha
VZ6zTGkWVtLroqn+3eCHFSn7KYScpE1n057OSHWVz3H1pHTRL9IL6thwPYVN4O1c
C2OBz3JrS25vpUjMPbL8Q89m3boj6M4YyGBHgwJvTmTw6E0LKgN5qG2UB5hez/CL
Pr/0XrIaMtHv9CiNQ7301+TNGR2VXYhkiG0awKURvVRN86fzhbN1/akojzuzAyfq
7/k11X4m7KjD8d3pyfB8U4pdpfVJNzWRLJYQ7XheVA+8ChZQhn8iJvgLmDB2ngSI
cYpjD5dZpP/RzLujlmE2TJ5V5a9Z2IdaXoY1/mIN5KBFIs8UbV8dPARIqdWox+Ck
doHeTwtiMaA0zG11UEcVKIRPY1KDGnBesrJTBXhWxa1MkuurYXsBHpC31WXgSmr1
11EHyv2CREzKc0WXiMhl3abj9JlG36uaUi9nh8pvP1GKsbZ3GnNDQrKlhQOg9cPP
YKi1VFlH9/uopCiNg5g8LV+/xvjoL39rYax8r0kbu6+E93KA9bMd+K0fNia/EZTh
brDBm+pjSC3U+SLE6I1S6BaPRiRWO/yb7QlUbc5g24o/nTQCoUSIH8lJrLlAIvRw
oCGwmCf4y9mQZjDoSqwRZRz+6zBPOz8bTf6iRH/tdTbn1NCc5gRQUwAcPYRsQcYA
Du1w418nJZorVweoLQGh65mC1E4PTlxkQcaVUoa/8Iz3ewRa4X3EuLmgmS92WyHL
dGXC6IWIpSn37pZkiuDDYb6sZ0+6veaEE5Wj12J4v+1Di4lWAru5PbguHB9wMK9k
Ruk/ATPrIM34oP0tkYrtB/TeF/4Okr9dubuNq24D5fu04VIlTNc6n5oT56z7FVBL
7XGAEwimhF0nVwu3znGOreBxz62cFY3HiEM0xX26aff4Sb4HLlu6tWDOCahUKh+A
paOeT2roed7BrO+ZFBuOAZA/WKLet0q3ivRGrnC/U70tkzxyXmQ3maJXYLasOh5o
mEVrZdtGg73Oj7SOm5BNLMHi8iyyMzDvZCU82n8G7t0hZub4oCE+YeQ/gjcxULFZ
gf5jlVnt1qsHX4hoGW5Qj0PYSssHqgdib/suQ3E5dEAa2LsqpfbV30c+uebidZIN
kiMCeuoKOgm7O1zDIsplFMM/Wu9TdYBTiiuqLXwZbbP4G/eRTLKT02Gkfuz4ja8v
d5oNpAoKRbZO0pzB+bC5GdFbArsEpFPfgmrkAyqkev4i1lnajF7p5k6DmZzQDA2U
CsHB19sK4wjLkBD2qchr+i1Ac+Dw7fWLSunZsEBP0rdxX8BxlRkAGmZwxZpatoy7
EMi4x/MxFk9CebUSWeraDP0LiaBhB5z14IDealGhVv+z7FdAwQ07ovuAckth45yr
STbhsndkrMbCXShnbh2zvDpQNzk4y0APcKKLiHxc8Jtp9DQatGs/+HAaaY1XfAIO
QW6T6KER+ZwqJxmr0zwcYYaa5csNWByUwtiHLChXmY2Yn9HyhF8EpHyDdf6MN2Kr
qwXV6FQEEI0YAZLlnnXJDpV2o4y6zaDg809cyaGlHVxleWp84S3HBMyWhr9IgJ4r
eAcSmXbV1l/DP1jCv/Q+nuXwM1vD8qlp0hzNnsRGMT9o9S2pAnpciJz7sVPrHGlG
V/5h2pujfZBHYAyNqC6qYQ==
//pragma protect end_data_block
//pragma protect digest_block
wBTvdCH4dBn1rzIKxH4k1iNZTFQ=
//pragma protect end_digest_block
//pragma protect end_protected
