// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Joda5BPK/UUceNxti2WibgdClrDpmD2nadLu68x9oVF8et6Som8jVUBwFEMX3Xri
vn4SqerNJgTfxMZoUWhybyxc63YNlbXxNXBPAlK/ECAz241iugdc+iW/3ge8BYAi
IFcW2QgNf7dFZmYTSZKs8YmATUdH9bFkN6tg7yQtjo8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 12272 )
`pragma protect data_block
rOsKFlB8rXqQBG4LBW5MYL0j6gvZAsjLVKZI3dG0w+vuU8m0pxKSFWWllRWuJL7l
j0pJxVElpkeA302CbCfhpo+eJynnPofKEzoA5G7QZq7SVR5juByyz56dSVuiV5RD
uTTljQ/QFtHBDA7lpoEQJfa3ry9/DXn1R7WBSbRBES20LYHyjom1r5z2At4fowsw
zcZyGqnXfcm4nOooMnanlmGO59Xam+zxSiYpYizY3/tynLBE7SwObw5Js8Pf1QC9
NAIa1BV12gp3f9kYzkfECgPGB5821f6A15JfQRiC7FQxdwQ64Hd500RJQeOqzs+1
M+8HV40BSTrqCJe5vbyAidUMY5uyeIPnkZphae2gGVc+cyWu2jq/BIZYtyDp67U1
PYoZ5KOsj7sEM6xoxyDn+Vsql0HAjySQ3d8sBZgjXe7mR2FwiZ9J21JMsIbXz3pA
zSC5W5vIt6N0iR38wgCHBlst4/+HEaLUrIqkhs3aq1wXyHH7WCfUz7ybzQvMGFtZ
e+9iFCbTJcgHCRNlZzkz3wgx2ebWEmwWtjTSiTCv9arYGuH9AY4fj2nwuA5ttttH
uVXSfWorjLBojTJ7YYGV9ZA3YuAEQYfWAjxZOxEb70S+NslpUAYH0A56fr+wpP1N
OKTaiVXG3TcXCWoKuA5ebox9vH7xdDOijFiMpUneA0e6+JXB+df/chFyuEypOBtv
GwW2XxkP42QavfYWIREeA7duLSxrpoyhJvZ1vjqs+WlIQonHkhwMbS9As+VkgUox
DcpJxT37hn+gfcg9VftP+J2OLe0B03aJy1g2FIgEH4vLS4qZFqzpx6hIm4jnkBOo
8APv7EJVKCiUTdpiGYu42g6kb4mxI56YOiDqwlPI2cLDviuV464q6iWTkYYz5yG0
PjRc17r3RxuL0Bvd9dJ0BX5xrArXjjO9sNHRBDpcIlQ2flXwVYYWsyTU77Im3zs0
Y2HEvc7B7boZtGBYqjdk6EkzXApvTUT6lpiMrJp6lu4uaiD9AobnukVQTH3OdUf2
E/CkiwuqnBoe6i2j7OB6hMWvSGi6wjveK2Q/V34Htc6c/iVa7QkN3Q7ofdYI4+n/
gpCOT7/8OK3EHq6qSOkmzl8Q3PU6khSs/bvR53SelDt5ld7DkuWy19+oevkYSmux
YdcAgnOE2qFPy72vcsTI9MhrdoPtY7J5nHAT7hkKSqei2pd59O4A9SV0AQntrt8+
Wng2rZQ5RTeHCsqLrAysOzN//g231e+AM1SlHjT/8LBsA4tIqWn2Et3x426FnYty
oN29BmV8sV6ivK5Fkz1t+p3+IHSB0jXYTmPh/R8A4QtlkDtszticHavC0p4F9Tt8
5WgIM0+wRNplLbuamNvd76v20zlAQmcK45CQmXXZjcf3J5Z4p/hNtkCMiqokOxUr
8ZYc6CzFGSNXAGbLcvfCjR2KufbireKIZJTgI1buMqSX8oedhV44HEZeQ1ZCFiLR
X67YsNOTf3iyM5+w1cHNm2MRG57FYZsGLBl9rGnMQSuUgTHpG/5pytkO43TadDA8
jU43dbulqBr3KQtmna5Dxn9rkZdWvIODJUdYLcOcyiDPwoE+sXb57oGgpcU5Bwm/
PMQblGVZgPaomYLpulaEUDryifFGhDRzu3Om2jCjywHJca6mRvV1aNGaSokYl05N
BJFqgVMrT8UytYIlH815t+QG4Unc4VmOneVyU/wNc5FakHZsk+lNl4O8RMlMg4iV
fSezIn3P9p1hheogv7YW5+I921tNfNXSJfx9nSdavFrSS7sxcxhFieoktqB/Ikox
7bENh0XR1o7KMG1vlmVUdSyN0OXNFHUzWp7BT4v6asPu59zbDwBS3MElV7lvDlpP
6/RKxvCromopw5B1CLwETlBBbtdICXQFKbHLBfK8/LQ03U1OPKEyvcCvwGQyasV2
taJ25GNEAOVtEHBLU9s0e62CMKJpbVCm9R3nRQTkqMlyACWxtIAAnqrjwGE6TAFg
OxTHFJjpbhlWf8vUMwP8+FjPTURTM3B8PEpJ1NPEH29CSnbT7cDdpEl8dCtH7d+1
5TJ6vXIwVl7tHyoP0oKpmb3xVH4cGrl0xtFB1OLteYg0Q0CCjSc4ZvHdMtI/+ZS1
RgbBimmtoKPjkp1oZm8+eZ2FIb7QngGJfe7aJEorB653OBSU3L8ToYd5MsKWKVt/
VLmjuQslQ3YbPk0mgs0HmFx4g8jZMpMNrYQ+nzL0kP4lsRoHIgZlJFrb+V9qJmRP
CDyiBEOQOxJyLhjPjzqAvAfmIQy4+NRCbV48acG33rO5iSj6eV+LxtlBuNybadOu
4nh9b0KDVUNpY9+rpeSSe/t8/znjerMnOLGwdujIFyp7O6yHJTSKsoaO6qim9PiU
MkK7t/ufxXzA4sTTD9zqZJXQC6BudsgXcgw0xCJB/9o6p4RLGXFSuhVnOAB40KVv
fqDXgTsbrnQJC4lNMn0iGEHjudD81TEf03lCVjXWhsV3VqAB1pX9OJVkDJQXQQ9z
/2rdUxUKD3J46ZtARZsk2sFkZPj/swHXVDJ8SsSjVePx3EKtXY0YHiWTrhBq8LLo
i8V0BDXjuerfAIutvDFXSqKFYtdB1PMxkfaZSGIHOXyPaJChgN5Z2GgBVGdU8LPR
2iJ+r6ehI5N6bf9/0SgqzpZ65AKdhLyUiZGehRFWBwkQwKxXjclSVZBDTGtr1HTJ
ho7lBwlYI410immlIr1Swuie+13xWuTkh1QtPyJwOnOjqjl3iKGLhZawYzSTp4l2
D9RtcYlb9GUxprITO0tjiAYytmReGqeYoYuOJNWtE3/5k3E/MvdZ6OTfzEb+oUSE
6UhKI1I2oqCbe7+ceqeKZRjb+DZzvZryEWeX0f2ANpZ1zFn1BQNdlzFzc0T47ULx
sNlI+6LhT2hpr4IvWeDkAeNweGetFDS8iU3Rnl6oxRw+0A16Gk2gG/rseU4cwTYX
Skuq2WZEzT746ecvNkSozJeVGHUCVSIoX7iVIc5x7KJk+IWbNgzsrsrJD4rhgF6c
SWNoLihcQ467eFAgPSnmHEsZeSO1eZiYJ404nX6Uptafh9x1eSQK51dGBeLU1yBf
HxB1Ib9QhzOyM8oBa8IhQ472rqXcW7jeN68ix+50r5v/TbUS5r0DIqlTQp+Bs5F5
OW17fxm+8GMGfENU3mTpocTLYKv4u2j4gkUZ4qWyMPUzHAUg5K3qX+U6nT4Enqzh
wqLOluPjuSfEUZ8JEDcQA80b1ZKiSyUnVFSQM9H2boChg90SNyOKW+9lf+Vkeua1
QTqMSKIWaIgOmC6a7l2F+PfAsjuMsPIryYMMQX673aJTkQrcdUeGTCKuvP8QesQF
LpeyxK8AUJobWSTkdeS0rrrOqo7idCJQk+KKPcO6iO0MVxE6IMN7L8z2WV/X8J1p
ZtCliaWjwXecO5C0TvZH+JuQ5YHQhs+YySTKQz91O0Cm5lu5s/NJMCDSIAvO4Jn4
NCVYvjhyO5+OZnOJIxw2kAqcQF3wkKtgVAIuWzCLzJ8lTRqoAQB5AoXt51/PM90s
KNkfrzmM9Jr+nbznhu3xA2AjzmMOEsxlApvNzrndPaiL7ujK8Cp/DBXdPHW5TD4D
ewQlyuaMFZuqpPdQNAPuD9qiIAEr/IIEP7XgU6znYreyoDnBNTdiF7ApIIJpeHIR
ZhK0BNEWOu8S0ygI+8no5vOJtf1RTWdw9XLgjDn+Q61756UEZBwyY5Nf2lN4m0f7
Cpq7pCu5AyKaZ2e8hbFi4kfjJkfwadm/3+0iELPLbxzOP7hk96Qz44R3md7SsvtZ
epYCbxDj/IvoB9YjP8DLx3vYfWmtBVtVwrBb5XDidEpJT/H32XvdjUYnFX2TJ5V5
Wd4K5ZlzBHseGn38rLURJkc8hK2RIFtBtLmYRVWmebne/IoA4L0Swq15TX36tj94
Fw0dsOkATorK7tk0Nxi8/nNYsmn3scEPYmw+lo++O9RPmrlzbCx3CGf3EHwy+5gf
Wz77OEA/4gIIqBvReUUDpvWbSIQPbihh00R9MK007TiXsehVIUvQXsmd2wKJ1Lkx
aKsHlCCAITndrcUrhq/LtOKbAy9a4GjYnzNbeNmAOEGJKXLEgLtRzI8ZmgWOqJyQ
HgymKWtbjXwg6h2kyJr407uuRhOwzFybZuaktHHpBAvvUdnJfTUwH4Iu4hOmJhWY
aVtyF2/E6wsR65bIgjeN5/3lnyD37MlOXJMBLyoCfZ+FUVCc0r9NnPpH957lJIaR
aklDAvyj68QNN/YCUDVua2ikjbaTi9sAKm13I+OzrhVltKBirzCfzB3qIkzP4khk
Umdt8FfXCnLCFMBIaW/FhzfnfFPh814aiVGWnuSc6zBbhe7616HgLwO7uSrdbJkE
xSB21hsYkmg4oYBajxbrxzrUxFKkD13j5DC8kgZsqceIJ6UiAdqEVFGE3ARwOlQo
K4hPnBx2fsyJJjtkvqJedcdNCDWklGnV5xjbxPDTW/LlS87oue71aZxcc/Wut32T
JNSMe5fet2HsUH7alrtuTcZYaJFF0/H4iqE1bIseUi774TpsM/sVUGOLpmtCKQqC
gl24XVLHIu2GMfOE4jDWkm2K4ERZeZ3wD393fxyBKTfV7/eOspuPUT2UitE4naa/
W8xqwGBrO1RU+rDVtj29ozT80R8nwIL77/TggeEqVSCWFoiiqY6ajjZQ30aBlKMl
tktjSO4PoCcdtR4YQ9TGAGmT31EOFxcaokmHVhdr0RykaxQNdDAmEfBfP2Ic07nO
wQt4DRNR2oZ1U9ZwbIEwEr3kr2apNVvbf9K/TmM9FdATK1TAHozo5pdyY4PNsVpd
jiqsF92zdhmWJ6b634tV9FJS1YPw60k648imf2NzUXixD+bjav3vy7a3vNA+7e5/
CXYwd7r+JZmCyF4pCpKj/gRv0tBsbJL/wgtgLZgTR4+1n869rbzvAmi2yIZn3Nfu
/u738MmPisgK1QmLPnvGY0Ec9Ol8bOcPi6pVzA8+7zRikxKfPHI/M9VV+Zx0Y9Yx
4+l1kW7qSOrqXwq4H4MS7AZ10tIEACQiCvF2iL1hoFB41p2g00XEIRF9ngOD7j63
JVE03pbQIBq2u4JUfpihn6m02QpsYXIh/TLB4aBurlq7Mpowfz/PrjsT7oPJZzrn
0vifgwwir5AqcpLgJ95uHHmuuv3ru1RlviynAGVbjzEAOstmblffc+1qvDjQf7E3
rg639L/CzBeUjhPH5irOWm3T8SKnvKbXLGqYXJ+Vv+JbeBP9UwDCYLEHfDrbocyb
dIVX12VYAyIHyHx2UgIx4snaNqwjciCt4n/IfDEZHr2z0QjL65e6aU0/DBi6r1+k
XQfyrma5t+nCxO2wXg3BMkbVMp+MxycMmsCoFESMzSiSh1foMu6EzFWkwlTWRuVE
woth9tHCKQoDcbzFDquS3ec4YUz2xp7cvo1EXEX5r4uhtHqAEx2Adz/cMPoVnHxl
RMt6lUQUl78gpuTobS7SIvwcYTpZ/c7jHi6C5J0wGPKGSBOvSPcuUdzgojKxy3kS
ePOn98XGDMsyQGQyPG7RbmLPbl52pZRgD2NCrasxNlXBV2bOiNf37G3ymWhRfnho
qq0mEKIpndssBe5HKEs/Z08XK4/JZwo+zqKbVBkMukV0Qsa9/ab9gTN0hBBQ7Uir
U01lOLgC6OYmhLlCeLdcLn3ZP/NbPWG/X6oJSlA2FM2lON4/F/VB2OnUnxAHRiLn
YE4KhrOJi8pTO6DjheyEx0APzpOWEMHwg/hPUasNJwVLoTWJ7yqsWWFXWZot67et
x4q+soQ3Wrp1EtyiWJp2/2Kwi4yn7RAKAsma0eTZNacWGwFymGwEupXfi8DY50i0
54jLG/3UlMA27/ooxyf6Ct2VXh+3Fd+krI8WcEP8mL1ys9xbAb8RmsdQZBQEq42H
IYmAaSxmeYSVvAWgSRWQ7G0G8+vQI6nwGL1JhpVp3ilMVPlrVS2R5H6ZXut4bXOf
qPj3ese/7lRoSCYZoIuA+TCzhakdu543vwQg1fDIRd6TGNXLdWYczp03F3597oBD
Sch9iCiUE2m/+XtCV2f+W9AqzrsfHX3f1mxjI82AVincrEvFIEKfRliieYItz+J0
Ao+t3dirFyrG7ivM13pnXxMrVwERA4DRiqO3PurTjF/Jxgk/atAHXK9hnekEnCLk
6QOdOlEzEawihaC813N2ItaYK/Rwn76z6yLp/39i+Y1GjGQzfr/6hFXoc4ltz/0k
7cCMhcgnhjsoS8ryl/UPYAh0ruWNS6tzTSUPa3YSNo6BBMy1wrVps3auMwlu/5i9
+h0nWNqRBHDxD5To5Ta3WRdayqyQjmzsfX+Y/LHDKKSlY6JkOKbYVWpb893BUMUM
P+OiZBx6eN2Wn8guiV0rkBy7vLuAKz+WwXRlBoZZQdnthkDZLnY2yhNFaqmHJdGN
A6inDQmwxgogxDvy02Y9oPumNuMyr9yYGIai9s4aInZyH0qgwsbEFu5YPtXdeA6x
hy6IS9x6IC5B7ZVrChOmPGA6n9B5YzZd48r1/84SW33syeJ7224Lucm3npsxDI6m
pG5ih33pDwtqbFhhF3rIo3Ql3pbggJ7l7maMIFp+gGPz3YLSvDwpDKUVwXpG2keu
u9ct5JBDWw4Ll54bKI+/cqF5ohbovklorb3nN/8g18tkmOYN4vuoTlSzPbgFa8B/
HWvRS8RjR0VX8R7GgqS82O3pahqmsKKY6p7146IChDAZ7ilWuPyLUiq+70rCN9mR
Gn5H/I36Q+Nt6ZP03296fCeHnmlBaFITaOvFZettvZYClhXazvSXeOB54ugMNGix
PCoFiuxaNXqpaHh917dznxlsmysvZWbTKHl06np1xM8Ig9k8yGGGV7dg7CtMrWyL
OhuenxdIy9c7P9kpkR2DnRQ8PgJDY0+mzuzXhOm1Wqf7ysott0z1ZvEqsB5aNfMY
s6qvcwRcxgFFgr/n61TQ9PiCHiDVEOinNtvTSawJ27kgG1/wckeYOc9Y1qbR0hao
VhcbbHacLjwrKQOHK6s26if0NTiARnlwJ6I+lzq6RHEafgFEWuSP8NCw1JMbOAVQ
PZn4p1gHxhG5Xm1BQAuUKTIQsR7Wu4CA1I4i8Mylr7yjEKdt3EkDJ73mRr5BzAmw
ZGkfeYkIl7xI3SPTy3gWu/p9y6sQijbjYxX+2mOj5ourh5z3YRygSgAz1+i5zuB3
8IfHgiqK5nAxBR9mc7Ffa9Jb1o11cuWyhWfNCvOd15hIs9gDcs3uh7+Dajz4llbD
Xn5IwbQ5/FGytVgAkYK0iUIe/lFxQ3OkkWQPV/BC0+lfdhAqzicgqm8wv/mWY2ff
iwY3t+0dZiOBg99tK2EDDSrO6mpeVTYUSFyLv9rty6rQyRsvalIbkZQT4pfWHjbs
mT8T/jYjvLIvZqX/YqbZlKivi17qKvGFVUNlzzLr7C+0YQ4DEXRlO201jtn8JVmW
UW9d3SPBu7hG85YO7IWshZ9jV9fDvs2rDoBW5/wFOVyd2ETU1wbCZhvyMVHJRowv
Km2O+eBxRB0pkGEKnxdnvPdrx0HDcQtZqceGZ8SlpSisdF1lw6xFFfGXKVjz86sG
vEQ3QXkyXWm+HsdB7kB+u8w8k3rOBq/22VSZp4V8DVadeICXXhdY875IcBojO0QS
GBgPmFKnXkfxEpL9e8R3jyj3SUYSME3on9xon5hMq9Ld7W2/SMNbnuTsyZnsexn5
xXBG+9dviDCixz8wyNl599Eqsdk8BMCmEILs1loBHOLYc0yKMcne3HmuxQz6yIcG
nrzHsy9AY9sHsZP4qxY6M2tPtxbsnquhtlWsvr4DBJpv8TpC2oN1GAz1KrydnIA7
jDaufSe4HgJhAkdmDRsKMuuipk0ctKjOSsAuIydsPOFOVkvMj6vuHw5xdSQaqXBa
OyXyJ7Cn/CWfpbTE+P4QmQOejzdlFp7j0OexLSYnqPsbxluRNgblRcnk/YVxjlrw
44Ok/zsI9NXl/WPzX9be8ztOim28HHZ2e79XR9evkEmCcG4Dy+eH6V2JAHAJ9vyD
Jv3NpJTDmIyQxRBAqlnN0HnbhRZq99q3npr6PIcNH8gTOB2kxdKh1XC/NUR0rqwT
AZQNqT8tNBOTgB23Uh8Mu61tLcHSbfcX/Oqx6zNtuJ11a2EUwqhbPAZc2L2dHyue
+uTT8UNkyZVsdOxqTV2eEEKQvojjV95BvNsa8i/cM3Ohx6HL/vqqmKqKT3mp6+5F
loZ9L4fKX3S8sPseP0PbhG+z+bdUKND8rDIB2RepHhemNuxnYE3ub0C4bU+PnG5B
tnGy/QC5qUqNXxj1kqn7cDVyxKibKY3pHvCHZ7toM0lYzdiJ/uL2xAL5pDwKD/fi
MDkBYfw+q3IdYE6ci8LmU+9U8ZBHzosmBFgrdX3nb3HXr+/0BfssxFY/yrHA6dbu
YtPuoNzmqD0CXXSrpVVl+x6qacR6bMTqWIx35SpdlB3cHtt5r5qQ/GfvcqkHLIGP
+IjFAmV3fs2SxwQP7cxqfxW0+j4zC/O9DP8M2X3loYHGRicAKDmtmvo2v9N+Boz+
3XMmuVsAcoLhJPNA/c34RGwRf0JcrblfyUN3BUKALtyT7PYR1daDAF2k+poPbAD5
Q2B0JCwsc1xqZmcvkkvvPWzkj5LWV7NwYjwqPCGj7nLvcQ/kQh8kub8ivWt10QSA
gDMDZtNTfzEhiEmDYSbdlN77D4nxXTub9CHRmJymPbDCQqIvhZibjlcyfJIE/JLF
iH1w8qWApTirwy53wBC0RAPECyzLb+829xOIvQEYlvd4qPO1UyHAJyOo8ywp0lvA
8PPeSgX0YGZiOv3S12pFBgFGsIMXqiIuQr5opfFoKAyA0eZhJLisRCcVPmogEOdL
gEx1jU+yqw1O0oqFPFqJUg+aeqfWe2AWlQbDn31+nM487MPsF+JVmgNNfJbvXh7d
ID5GTCoy+SuJC4n3dRJIxZM6wcbC9b9Lc9Wbea4RlgVtIG2HLjKnPEI8ve477pmx
Ch/uY60y2UbcpmuRPS9bjik5BTUxxhXU5LxtO4xvswTNGxSpRK+xx5QL1iX1cPkK
JrJ12hZut/+KfZ5/oRXgQe3/1hLqFUGxE3o4QM4sXEHFIf6kKr+HP8iFib1uZ+aT
VMEBhAViaBBaL6v2ru0oUjuqG2vNctFJ1PgMEA1+7q7Ryu0X96QaCAMe+Rfn41Ns
AffGBRRxB/m51WsIuSko3x0SgLQtstevWRngac9LhbSh02BfrDPmScucnu8uE81N
E93QVe5uApehNjLvkoIVU509yUIyDtkEqR4KyB+EBGRLGreClFDR+T4BOnecVE9s
szFz2YaDuYy4enefTEGcSq9vaYeqEOQXPvwuLXmSc18aXHjyV/mjo8/AkgpYJKGS
1/g1GO/WkaCVdQRzfSz/F7yS/MwgQP7Ag6czhvrpKK0cFUeAFHj2kB86sU93SGHO
D8xJnQlqfcjP14zly2+MmTLKh5J70JiMNVCermE/gpmLim6cKSxncQ6eeJNEQrr4
n0w3Nhwa1XqXkm//f4iXmcYsTiwIzT5JIbfab2fsTDrTy9KqzusEEBga0MLRvj5Q
AnSWMSjHZUHUllH4kfXUw8KPF+7Le8vktu83mdj7OBq0yCWj6RJ8hPG7KSsazwLV
dsbgFZmTzDWHWJdK6Q7iyYIVd/C6ELi/L/fIm0I0i9LtDx7tuWcAanWS39bqkYCT
jNIY2wvoiYIYap5Xx5RkHAr17RrMS1V0QUju6rWdaeylkFXuWwfwb/bDfFctYwlS
8nmmIthQ54RrHtBR6fIxok34Sc4MQJBnaJrr26SZcmdtW/OGEyAMhI2VVPk3fUZM
8iQzmWyfWh3uq1QSAQrHGYJ+SpWNEIFgasMaV0MPZWksJuj2eU6LYU+LtDU349cz
Jl+X1unuJ0mqlgmq+I4zzZiSGcLF90b1HEA2TXv0GbdARUHD2KE3xLMknuukHsBz
0UbBtHDQZmtZ77AeEyIDmD/u4LSmJcuk+o8DGcGAOvus3LsAfZnWNXtZkWVJ273c
XzKbwFOeCjnS932BwMFB+voU5JaO8dXh/RUinERzNarFgNVk/WGRXUPatyvbkril
mo9QToKBQro68tukUS3PpNGSqAb6FoTBiIdCo01e6sCGl6UNFk04hCEAebfiE9Y4
2/V43uhf3DdCRdDoa1IGSDidpLnccbTjPJeCpHBse4Qx//mGyeB8N3+b72xMPXZV
pEWv+27Gihe++5cm20vZUgtB+bQfp53SKAW/AXp9HSsRYCbiEh2PB0AiwPFKVpFI
mDg98JPbqPk8Ssg4mMu2akzCBP8OADdvxKwVLZ5zJlvfENGzKjd6iie65U/Y+WaU
2AvxjfSYXuhSYYLaPosym4EpMWOy4KVPx4u7jEyHNN9voGhFVRIZ5DwKGhdhb+6y
9RmQCSO6OAFIvqYekOHu0HAfInah5SJl2bHVcQ80FD+fHkMMBpJcUVrMXOTsS+Z2
Myt9PrDSf83ElkZJURTABn/Yu6o874CJYmjxqgPj3XQuZ2xboEICZ8Uk5qQ7nT+6
MNqVwbUJ/0cowegWjbKJQhSg7sIkz0u5SAEGLYrFwLvgeXFHWpLUEa4JPjKqgDSf
I8uAV1l7xxMkSV9glaRuNb7hZj6dxaelGjAXTf4n7MfTRRImaSvbI7mletTLy5xQ
OoJjBUMbAC93R/ijFzysvpVtWJnwnO88TakOejjD7YpEHDSdca7iQggpLK5bDmX+
dEeC27H/7fzrUKNjaFXOhZZ8L2HWyqineaW8dDF9VclHpQ4eWfAjvjRLZKBsNVJi
TNBjy2FAnY6WgvEmCoePrl/nijhJjtvenwI1FWCQh7NWatwG1xk3ffIG6TeA3+Wd
OVHZu7eVunua05B+FVEc4O8+oOovGEMJA9JwsHc6e2vDBuSKylsbGbWmSjS3iVKo
uoz0mpSQVQlrgRXbQ6zu3E79z0rnJeNzYLEwbqge9O6ATLTbv0rrDCLR0VSUaFQY
1co9nxB8OwDpmie5ecxP4VQfBaseDS/ZO1b0ems2jkbgsHSke+10Qe5mBIW8mJQV
TfV18rE38ePgFdtZJj8h96A17luGDXhYaLcOZ7CVvwqzJ6pXTpfwt9DJdO1NjG8V
XJwE4SCKU90gFrv1yuS+SKO5G0fRySmTPBTLqNieBgS/nQyliD+6Ml3js3xFqJUH
U7HraZc3iQt+8Cl+l+37Da0BzrUU/UMbeyBDI59fIfSVHvKYNRNdJ1g4+lvtodVV
I51hxMKf/Z6Tn46K8VZb5rPpbgnCIOqU7XrAFfP03Lr2GG/AUc/9EA6U9x0UNqpN
uxUltvT+Q46CyEIizWT/Eakb61S7QZFyobi410KpZTiRm5F/OM3d20sBhZjCO7kU
hrhc8bZdo2UIff1IQvrjo1ueACBUJHyOSNofGR8lQSGRNRP4caeR0vPU8mG27h7n
D/3nivvxCdaMM96601P9vmW5Gw8rtGtfzg0uioDUx/2pb5stupMBfEgduyHaLoW5
0a2NGzT+Cplrshu8IjvmoHAwl1D/QU0jEu1WhNFqtyqyOIlnyRM2kqDANUd4vZTZ
GDhCmh2B2vQjNLswvhcyi8Z2FlZBWioAvVdNNyhIncVvKN34DDC9sTvIghfpnUlX
r8ATzdpLdxzByIS1qOPiH2iw17oG+ulakncCwyr8YWoc1AuS6KsT5S8T6YHSd1CS
IZCVR6COG5x1YJYf80pCq8xB6zKm2Ru8o5KckhU62r2wBWuAVXKdQXoz7/v71cFf
T4Lwv1S8MTUhXLHAolh6AhrPn4b2smky/my0l8wi3sFodBwgfSue8g8PzM+Yg1+k
ahg5HMtYi0F83onUgL4PDKfZCRZVQ/TaPOKvpx1fcBSbEKudHuds+JPYh/UTALw+
2Rd/i49G/+GDhLosl06DgQ0p9FVkoGgckfl5fxaoFGN71hTsDlhvsnmojuGTQAFq
e2B2nXV/3r9Rzo20hfvJYCOQXEGPRnS8pQFcyubBBLg0GspAxi7tv/RMMnOFI0YA
W9qcwL5igMas1eze74AQPiV+aW0R85gtulem24/LJvtuGAfM+hfrDinrVCDL9zfd
nmhmYZz9avYQl9cVUfoOAk0yGACnhv1qY0gNxkGoDxzxjiUtWLKkkiYPvEkEtR5K
J65EtW2wFNFfHVXYw+QPHhA3qUCF7big7cyBr6Cm85y4lZ5uUgfEVNhtxOka86Zq
yhCP6LxlDB1vOT20e3CaOQ6Ak3u/8FNurRow2uOdZDhEMVGWolkT/Wi8gnSOv2wJ
NdI8bjDeERYDcTkVbBBojIRC9IKJUyvz1B2/VeGxE7b8Q/VV0Nf2R+vk3qxe+Gze
QN+/Qjq8593d6pQTPsW86nd0nVDKJhUYkvMquuTgvB1Mev04Ly9dQ8FppuNaoEN/
1dfgF7QwgCZV9aXESmluoD0Sedh0rbK7wP9iYV0FmXjjjto4wBWt+Alqlk54a3+q
cWiu3UaT1P3W/0qr5x7pSRage472U0FUuXgrZu0JxJg/zNKhHhQQLPjZoaxJLCP7
reV8Fb0q86eNpgG1XVtehUz51UP1zKIJicakQ3BBt5cUYfvp3N3Lr2QjCckAraNS
QkSGJ1ICnoaSmkRh80d7Yg0hh2AexqbBkM6voA4ev8WSnwsZ6oSsg8lUKoHSVQ0o
CymynT3KffwwiZTjfUx6AQIln4FCao7spCkq5RcGT8VISC/VD33vCfVeLoSzx9kD
pXYEY8yBv8HwRcz8JcaFaKuHklD3EsQzI43e0doz8NRzCdaajJWyx4Voh6QnRdjY
5uUpBUIkh5MJyoc73RPuLKpX9oGtf4kUDN3YZZ8S50jaZciFE+9Ta2FEfUrlzMtK
Prtlaj0pHV3ox6NgZtlX5U5Vc0jfagyZbJHTcQHaoDGnjpXsV0iGYAwTPEINSNtW
HHCNKxMYtKm0/LJ2ML56fU9dNoU9hQTM+RjUeJqvQrSVOsEt5iEJRMngtUY84tGf
sO21LLWD5chzKMEsReNbx1FSLjJdEFCdbA0H425dT3tsN5evb75Lz8C2TtvZL+mB
rYfJOV3xLd9+WB7dyp6M01800fP1GHYzOZ9dOW1PDX3MtyuMOIGBMQUSvW2v0nq1
2sg1kl0/oDCrAUpgb8GgQrRKhG/qJARIGLTkPpmJOu3klo1Ji6zw+4pCr77c5kNN
XOcny+qc0+oWxS73392OFa9nqSKo1i4J2IjSm7KTO377Cm/CRuz0FnciqZ5Ilclj
AoqWj9DD6eyFba5oLIuri+RyS3geQB8IC/Cf6ZUs39W4btiOUInT/rqo4HlsitwQ
u0gP+0gCIovW40fov40MqqYlorjvCsA59hDCodNr5MNkGSrOQPoyK/D70tna8IlB
7KIKHqj0s9FHK60RDOIDbcXRNpa8Meb4pgfbo1IsSoe/hL48AM0I97YlrD9Lkait
DhSQzGezBOkI2Qv7J5C+R+DiQU7C6Jvv33v67QB3Mj1OuwBkMiPTWHOqXJCFPlKl
a27EpCrfnEGAJimy5oRp6zt9QQpqC6C2K8ZEGKbVzgyqYjWVsU8FGXb3FrF4tnIZ
H/5J1g+PxB0J9pfPH7Q/0JFUe/iuxCcynbtOa6WxYQiuRQ07rkZoq2sVNvYFp7NQ
SyYg7Lq5GgnmHsIwhyQv7HPlumEEPdfGTexc0rYAkcllCLGRBMF2A262PycPEOcb
96/3Bj6bqCNcAXOmXBcgD21SnoZk6QfW2CV5KwtbywNvq5X65PiejVJrk8QvErZs
O+aNW+v0MiWw4lkOLq+HaxP3NLrSS97Bla5KvY+iLQObOUEQnciKRZ7OaVz552xC
9Yh6MjsIneDWxXcm03pN8KH5J/NqTT0j4M2+6vzhxoHepyIJswd+PWf4qx7QW5yg
lJ+PqugjryNmTo/5IXGOjsQYNBBP9gD0iAslPXT4IOcBHXU0NuBbfQapua+EyxNz
n9GbQNl0DU4jcvbOVvf8fr0xPWZk14xTl+lCDNQ8zWjPw/N/0V5NA+bMnpTGUu+q
t/0eEGCaGdJyoqJ055edlxoYbfnteJRv4YwH40EL6km1x6cMhZbbvMyqKkxFzss8
wVFNTmTT1jYKeHKhsp8wIoVFyl2QWHGFGTGiEQ8gijTjXRJkjVTZ1iZGApTyDOkn
1mCd9XNp5k6bUJ2y+Z9qrs2JPzSpRsgWr840/udpaTrQ8wZK1ti2SyrD2NPCRikr
tPISF235vf0/y4LKy8tPiFH7Ni3mvonscO4Mfv0nsIcmTAnEf2G+J9t+6gFW1foi
xETlXCfWfVpT9o5pYV3EUpPkPTYuBKKjbD8rCcG7RedDw5Wh7rzNUMefMoqk6wEf
sFA0Vsm1jxQh5U1AE69ZDaXSIg8V60SP1cVTqW+Z0yr7WboHIJjK4nR6dZio5fQL
8/x8U6EZiguQDghJU3/SXWdvZBb73RxSvb3jrH+E8WNarSC/eA/LaZwb0L9qh75c
HrM2RmlgGUyUH/yiWE1mDNFfVIu+xqwpP5axm+jmCduFVd6i7BcKGSbeN8sOVMR9
dT/hhj5ZDY1h7B5ucr32qEpmLHmH8HAPnA5q3DjFyRHuuk0aysH8Kf5DOBFwlLEC
CUZ53H87UxD2CxQNz63DTP8yW7XAv188HIh/ACILrLGYeRKsOWotnQuZYFc0I8TG
hc+/wQfwbllSm/lIDH/R48lyowtaHvzpfHaJGrrx96r3ipPJSkl6e0DF9JVhS5e2
fg5Ml62PBgxeMj5W4yq81bo0kPGnphv35gSmjh2gukPvJfjMHV3PsdDaYXTjmPjk
J+TE6aaexiB5QVrn2ZRZPwZ535go9u91NKJ4xO/fgqDxhBtm0falFkia1Qpj8JJl
jqN8Bv2fcROZhv5tlviiZuZm5RoTboQip9ZKYglno9MD2oAPKFPltg1PYvSSVVx5
kT9YwqCBmqvogkR5MNBZvjIl+Oy0taGN5LA4hqgYvwaOuBEBK0dQ3e3aHmpSEM4w
y93wtinngL0zcL7WS+UmxevDdQiDH/QtnzqF5uSkGzchw5Sh4jh03Veg8xAt8tmg
l2e/A0mzsSM/NvbInuzMxJOMOnPnRRmBoAkB53GqGeL5aEJoWsMjiq8sjnMSv/s4
MP3IQdLxrlzN9PnJeX9bCFIX4jOpzAsguIA4RYt0C28gZXfi2Ya3Bcg9F+hQEeP0
YoONiuXrUAB+0I6FeL5aPhwTWBF9yknm3o+R8uFHRHGUIY0qeTFD733dHz9xZOx9
71SE17QMdu69KBquFvjfcqYtJ/MK0Xu3cj57q9C2pg4iPKQEgHk4p23ne/Y8mi6u
pFn1ne5hzHO5L/U+ZRk5NKh/WfeMPDQ4PRXe/nwJwKbyXD4o3m8Ta12MH1Q5/JK6
/P/PbLUpfw5v8xqj5pWeBdlC71IR4Oo3KHvt4Ujp8JD2A/QebaCmBJLUP7Nm2Li3
yuz0HTVJ41rLMHqiDtaOr5Fi3fMdPK4vg4UVCzW6OcpqVz1Kd4y3bbtQh15j/zFs
ohAmApnld55BkuOFhheVXmZ+DleJN3wAF9qJWs+vkiKcywYxlHIEQyDggRxzmqTe
mhaT4I0A/e0DvGEXC8UGbLSwBhsQoQ8MB4WYsE2sszXe0mHhXlfaQcC+aSxQpeq5
WYR2g+mPb8lSLXSuFNwUeo4dCs5xIvQREDDLhOZVBhz4AWg2kVtOFXI0NYl/QRFo
V9IzUke8yiGr7HS924rMAJk51AvK4LE08Dvl2NNM+9KZU1VjXcdCFpHWDXcq9GIm
o/qx6RWPLOcqK92WVBktN5f/bs2wyWkJPpeLIqEsc33Fq4+Rs4Kh0bXeBf0joy2i
sHgrVsIg3qlg+7B3/bCsxdcS2ysHllaW0fNfk/BflRv39g07HsFO6cQRVtQFCVrD
GY5eGDdjDIEB10IrAsHb07fHTGtGU8Y88yGVJykMrzbx6yyleRVq9RznbPTrupv6
LqhE/JNUj4wsLIBuPYeJmJhHaTVdoZBt8s0vZCSgtSfsMEBFVrs7EoJHw2D7uL2h
1PHGlA0841mr8xMhRjEuYXNeSdmrAsvxUL5/qm3fO/epGMjbicqPXi2elMVfjsEq
JSSSk5H1J06cg5shpz1Ktgb0OK6tqqtkeCmi4AYTYofGvy8rbHxCPX2mkjMNfqrw
eEg5SAr10XnxVbt8S7cFYR9cbvk60sncIWKXGL/ZE0ll2tLukn+svSJwFQJWZvU0
3+z9Zkb9lNVS3EESC8XJp9MdDtCSu0TzntSI8b9Cja2Yvh5Hy8UJo/DEfvgwDSmS
yPegHDvgmNgymWKyJpenTq7E0OMbXQ7uLNFQUv/LFJeNkGxAf+zQpnjrXIvyuNk8
Rm1olUykoBd6/K++WDlBEVcxUNSaohtnsXI4YPwEwMcLQvp5TXtlhXMNrOcKsm+g
gpoVRYWOnINdakHeCVOZmTEmXMy6o9as0Iu32FD9Dz0=

`pragma protect end_protected
