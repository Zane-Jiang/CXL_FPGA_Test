// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bgcytqHPBXH5L7GfUBbFPJAWiqssgOFCbz0uZHVt4s0qFyl0Sjwxp+srHsNX
+YR+9WAFKwUcaauHeQlFQyaTN9l8/qYiK0BRPJaDau00Dd0k011QDDylPxxx
t9Q2J/7Uvzfw0mYC4XL81GrvYsGJqeEsP42DEwSIF8TUDywQ86Ifk/KlK/Lw
qJrgskNbKR/kdH0u4XphVQhpI+hBDjXirZuB8J0640be5pyMjj2ntaFZCsjD
Y8s0kyCjfP9yakFEcH69bNLw/zbXu5fg7f7kA1u10n1MDuV22B3MGkbgdy3i
MfK2VynkvhtcVaWJ09G0k0qvsyT1HdrqjNed1TOC6Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Da9QHcLDaZm3mhRQI0U9gNdaNfW5yIj1RaXsfu5UokZgm4Ewc+YlYff4r8NL
sLztq6954mLzeUratXbusoMWUnxspdbc2V5ywbF2jbI94mkDlnoqIChTGgxC
oDE1Kk3CHLat6B0KiHE2DKFhREsI5S1/G7PtrsjtSnfTOIiCCbZRo8V+CLx2
x5xJp9+zrPvdm70z01SsP68A1ziwuah9mUclxwDGLPe3sXL0AYPzmclyg4xK
+4Ul7FPVXXIDCDr0H3XlqnAH498JSVFEqg9Rp4pc/QsM2luVx9LbQu7hTaAu
P56JjsQfm7dmWU7CWe5tvH5xvZRiUaTHh64pPc0SaA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S3anGXu+sHqiV6tb7OaUJ/hHfLJ/Vc9VliRZfBeIFRiHqKj7dzRbqf4UkkiS
4w5efpfQ988k9PDK2/h3u12Ayl4nuiOmMfC7ggMqkfY9lPGhacCZQ0dan0DR
HpiFpHJbUo94pmoA6gLFxW/mq6AQpCdq9MKZJSvcmVZDCu25sw9VWNUy2opq
MW4Sn+VWuqbBsIslrHAg4sSDdpqtX/oMxHy5BxVR08KLWMnudNaJiWu7FIg2
82TF447n6sr+BMLGTKbDJejva0QCfV/4SEhbrAQOHOxixFqR5CdUIM9Zuv0I
Fy4+JsBUnWFKFSclApgCdiMWWlGKws8oWn7Ef/Gb8Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
D4uxY9qzEiSbDQz03PMRV9unwRRHjngt1jBqlo0BAxFyuOhm6f/RPNvP4rbk
C2vhbDmNdTiheNphmxSQ2EpSG6fhbQkEMmxlg70kQIbw0y0tJfx7uh+dl4Hn
PNIhESHUgo5IyWuYOzT7PvIrfUqiLdhxQXaQZbfQg1VuZ5zOukA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gpAywL9ZZD0/OM1iFtfk1GtLRhSZwmWtjcWZFnzjbwv/9nDooDCURZ3/L1Dq
bqlpKk3cQqxeEPrf7UgbMbP8JE+7/x+97sXAV37ma8SrV2DgnBV3kKVKL8+G
X7gDzvAnplQzSf2VaFlIZVqQ3NNf+O7hRb7hA1daYUfAgI2mAaxRkrAjG5qf
WEJfU4WqIWmkwZ64PihxXdYa9Z64NUZmQEZjxSHglTnbhM0R6s8Erv6+SpA0
pLgMQuJrn7x9vnBpjCzl1rtbutyIoP8joNKXQTCSHIALRsaCU+v2SlkZvntX
CgjEdK2BbWMUK38hLPfz5o8bP8B5rFEc3fJHoKwh869T3ZC2JO+C2oKoWGwP
vrklGzaYS6S9Sz3KJysPLpo6mP8U32sTQEsK2uAUoloiruJucKWv1FVqnTQV
eKQRBlv5GB3Za2oBJjgdouDeLOHhFsnP9tXmQyXzh96/+JEhqlKhLF+EHztP
zuyeM11A7UdkhMvS5M4c5dykI0IIOW2l


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bwxu4kNFIfahTDavJj7BQ+phfKLF87S/NLqavhdlRddgRBreo/rVoYedVODl
XRx7hcRysuCvINag0ATkE+O2IhJ/xXGoBL7p0pJQUytwUXWLPgdAKGLe6RWO
8GnGQc8IX3sYZjkZR+3r2ppnchDiDeYhpR855D6/FQsfemcDkbs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IZUJhbMauLe22a1hOk0QF7QrdKVCUBkv+GKigQ/3Y/NGfVBoz30mFMMPzMhW
tnen9VN/Oq9MRElIr+ZOSlas82pPPNpVcm5A37H86sgxczmu4Kq6WmDTXxKb
9iyiNxIW059vZvSwcNET0Lx7P+5eSS52ICpE1Dm/diKI8tUR2b0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8944)
`pragma protect data_block
y+HAnFNHaD2e7BpOrNJlTrHaoDHoOmr4Ad6GmBkDQ2BVqHOhBhvOh4LdzEcT
5k5EFGYpMzMuZcWlFscayfnIYMaJoPRjkN/XS0PnzCvRIa13+X4/sfd43zHJ
SwECTDXf12wWuf9rWbECZnW+VYzoPE9hT6AkdmLXcE0JWpA7YLwoHGp5ki1L
Pa/KwzXng6AJRHCrFYNLNDw/5rutFe2RmE7PqWRidzUpVgv9+uYdmgYhLSW8
l9LS1+rE/omaDwv6vVsKrBS3zqdkpJg/v7xMofNVEfSabPuXt6ek7MuE66tH
i8MUvrT2dt+TKtp8wbH6zTDZgVytdaiXMhT3Ua82+PTMuG/g/rn1Eo2q4zYL
ch2VskF5kVqzbTIgnxo4svn59lxubGvZlTiErOuKOo3+11IND+mgUTsTbMcA
+tDEP90M10R7LKu13fU8CGy+mIqSwIjxg8P3/t+7soHBXPm3FiY6pU6qYFnc
UDV7bF5zrqiQGLjKR7Z3tpxsPp+WmnUIRiOtGtlBoEYmvz3eRAsEMjCmBsYJ
p2yTS9r68p/akNMe+sU3wqCxmNVnblgZnpw8geFIf3e0buPABkeX9auLqu0G
0iHo8igzbsNlNAmKK+nrQMu7JW4tq/bGo6agpWQQ8Vvab91+dzu+Jozgj0Rf
8AzypnUsz9T0gPSdtzpLxOVM3uIUYZd0d4++u0I8JA5xPS04wMPTLm1mLQjl
uM69yZDEU5FzBhKswhIFkoVXFcLqKawiyC3cZtVrymuzWOs7246N/wyBpp20
zaMgQdizW5SvRBlB224mklhdj6JnreNXXJAv1dfvGO2q3WVYUpEMswzRJOiX
NvbEaB93wXx/lOsxYD3KftyfLBUBfA2rbluhh5hHZNbBqoPtuiT+28clqZD3
ACQYQip5vPuzaGDCTI/32B+UFe4E38CkW9eW2P0hzZufkowjDw+RnZMCdLZ1
uwI6oiQQYbs+Vz6QKZzPnm+t4VghgORqyohLPIcqnHTjZYymefCBDG6s1csH
E7PMutuu8KyGFf4PbpYR1iG4V95hjtZsUjVSfnRS0iw7npFBRRE99pWhIzrq
YWrdhstTg+DjK8gdi9kSmkPR0fMDKaqHQqcSRlVY7tb8QC4fZ3W0I4KJuMry
lVEx9K3mP5/QIiyF2pzhhFMdjIhV/WhfJvmtM5BlvdM29QvvKZipZXlvnP1j
QrvKTVJwFqsK80nNv2a63AOUqO7hbsyaJ6aIDFvi0+99sRfo+tZ5YEoMKQqE
uCrMRbWbYEi4KfRNePwjVseLE3NuX6sCJteq0F0NlHDVJGMRWfbQCbX+N5am
Te7EBMppAoRIxkO6dMhrsljgvMw6+N81mwHXQ9g0f6p8BFc6qN8E/yIKgish
p8cg6f3N2Ugb2Az3jbHAUpK4RI8gcoEoYYbJux5TZc7Cp6yLLcbRLyYPheN9
88LF8nTOHmJeupg8D9+0EsU+W+EAtPLOWPYfMoU4XEDwhla3hgg8PUBCvaoJ
wcFyx/22IPQvYTMKtobKeo0EQd2sugL1RodDfN07KNCZCXlh5hHWjKkB1ZHQ
kSBTK4le9WylYYqoX9Jm7VJ+7hgPS+UQNwWaa27bUp1oHfKeFwF+D+jANLfU
G7zD9Ho+Gn+kAVLiqRvc3Nm66flvBt8gmBhI2TKmCAGFNrgSGDrUOYRsJK0T
JSGOUsKBhuxXlQfnhmHXfNFGSlvpo9TrVR6E4Mlokq8JmmTqCwDSD6WfBZIa
A1P7p4fp5q8J8iipU+KkfvM7ewT2sJDUbpCdPYdxRmjPvJCtljDPVyfZ5pml
/jnTIXUAy2g3BRa1j5Y7Cyl1aNtewiR4l+NP3VlDPkJ5aOnEQHRJ3L1IIdQ/
sxj6/h80K+0XH3Ar+86D7J946yjuyw7JCOSYRKLTcqX7g658CqYyozgSp0E0
ljY8KSoZjBMM8LvgeMS32eIw0U4iA2HyOlndTfcm28cwgCl5uNCJglEDGE/v
yPHQMFUKuoUWy2lB88lmhqga45qttVBBq9IdPxgdojdKwPh2498AaRsL4eoN
RdXsZUTTNGUa6fdajKlbgPOtuw8i3go92qZtGra4J/LeHcrkEQchquIbZOkr
eRUE9nsEwgtO2EYDttvo7bdBfeJl1jmlcE8M+h3fGyfQ2uq999bBY58hT9Cx
6qKO7N6LnvAK2JvdE44MvxiiN6rTNV/zK0hs/j1f0PTObIdSdOk1F45KR9sC
R+DWOxyleyzK0PZY4GH5odV8RDuBG2+UuvjVhDchqbyt2UIiLbV7bMy+Xwj6
vvtaKgO6tjDH/hMxydy2t7LjkKE27rMuF+SLK00If8QYLYltWdcjlQYKca5M
wWUhuY6NB6B0nM4CwmwrloMwQmYuVrs9NxP3oATQ4fBjX0rL/ExRvgEvimlp
xKkXvpBPNxyQWA4Lboo8Rhw4jqyB+nC0WsKtyFxa0mIkeNoy42unbmbQLC8B
3dN/t+W++tj6jgiXF4indtoIzMQvbcdVgxKA/p2mjIVwmHXiyHzlDRIvE3Ta
FCWWZo7JXULCzbVPQbmc7NqtXd16Fi2R5i65i6zSSiHn9Hr9YnwDvv6mblys
mH1WwssDCLie3uiD/44qAxV6EGNiQtGYgiIV0nDSgeY0XwFiD4uKaLhZHfAB
JVie5ZJzmWD7dbeXotuySK9BRObCqi2CODndOZjQqp2cM5EuAMgg1AAuQPth
7KR7PKnhUbSTSlk3Cq3wjpY7SmiwJSRHlRR3xPXsZLbSi92/NEkATeEujNjJ
fwcBYh2S10KwqrVwL3y7PJq+ZMuXFpwdHOjFEPQuDhj1dCi3GbiMXEnuEwkC
W+Ufbl8AgB6agEHZ54znIW/oaGn/sehBQMg0MRA0rGhX6HzviVEvrN3YvSvw
o1yV0sjaduhqLEkN1aXWI8eEIXNV1ZfbjZxRioxpIY2lwjSKKx6qeFJ9bHTB
d9z+1M3vK2hIy81OD0beUjoD/OMjR7tjLE0oMAqZ2caoQ+6us3XxyJhRBPKL
N0Tf+DH6UBCjKKBHEJ3Gn8zcflDqDHiUE4m9I+QAfCWuIDep3sCX+ZfTfrZ1
zmthF140O7Q0iNgiFkrrymNpDlA/c7QK1juaDirjj8Ye/XaTkH90vrUC+rMF
qZ4AJRDEe+AKPli1yqnh2Rf27tHqApjKh+B+n202RxZHDkS76aAfjwjBReUE
/wGDhd6HjCftA9FO+0zuZWT9V5AxdHFMh+9IdBiPdTHoqgT3C5ppM+NexOTJ
VhDnIuPmeUbdcpa4cEWYKzr2gaxkbj7zUsKnaKaZx5G3RKUNLa75h0OGwRMv
0L+GfypSp2GOozYs3TLsKUYLFrWyOHrM+z9oabCr7fmsF04pCi9CqyOj2nB3
EK5gIS9xs5Q2aKW+AoZxaPxZ8zM53X8xIS74lR2cK0N5cO578xzmU1RWJuca
z/shmz5We8iL19RMff9HYborwTXRLhG4AaCQ3z0wyIWvVJvgktKvca1YkIdy
mhQprA+a5Oo/WFl6Dmt4f1VSyoia4LSLkVWnimGgwINSVrtGe60vXGW5C/rl
cMON6uFw+duwt7rQz4D3zdUuRv8fpCF3pTkLu1oJBKGUq8wHxgxetLZzSiU1
H4JSl1OHFzPIwlRSLcSoBJ5fNG5ecSTu4/yBGV1P0fsZugqTpI0Tzs4F0Hnj
Q9Tp2+rJUXnB0V827ph1GS2bK3PJRYtE0XgwnqgGUNvmhOO9u4FCFwEbF1p2
JzSW0yARMTaTCqi30dwiNM4D8Z85FjdnkayDwYPWFwFaQ0hBYWEl/2kL+dR4
1f4m6ZajcKPUeh0lKPRQuxigDj3SYMGlFdV8J5/r0BE/Nmdnlq2NLnA6jhJB
J+H0oPHkn8OsB2CJ+HLSK21UdkvKlW2thlbwOTdtapOAzE7d5RHyyhnU843n
tscysgk5NkcGTsWoxB8P3N2AfpMlqmTpNbUfKH95m5FZYGziyQGR47wSMpnA
F6VD62J8geD+WMAJmSRTI+phh3ojSMhafZRvQU1xKVvBLyc7ptkBo5G0YOiI
VOki+qQYkUfQXHue0bsGBIl1+fSbzWAoQEo9rU63J3Va32frPsjhVddt8shS
MkVcQ1xnWj7eJcU0b0RcHIAKosSJcltkaHKIvKjkyALjAG4NoonSsPHvobtf
/8KuRz26orkb7padTMj9svqf7YEK/GU9skLyCf/jL1RwZ66YY458VTzJAcjF
pAkKi85/E/g1pXqeDKeI7wA4dlE04v7yQk/w43cyNsv9U180KVv+gRsu5eN1
5fHm91wNNuPinoJsxuiFJnd5qjnOWrKhbGuS8ip/cxj77Yg2t3Dvl8reuZcv
orKPxBT6Tt0X7/kUK+Guwsxe8jfAWwDTU0HCESjHTP3Q5Gyul0d+/08bJCmN
lrZ4c96EHgwwoXj254MzFjD7r6qh10eiCcPAP+DPh+37yO/ZnYPvEAZRsMIV
ZQvRffqPCr3HEQP4Jb1ng82x56u6yI7Aj/A2ieVc7e7RwWoHfKCeaD2BWBYD
iunhzMHeVxXvhQQwCcHX2WQoiukw5b1eXUCHTOFo59xDVk6uV3/UW50xhJZS
V38bFlu0DcKyUkv4bT+NLpx+bxvuY08EdTpTDfpzrbfDlhqEhaPXaqMRaA5q
5AZ77Rf0CqWVL+sSm7D1NT0qhKiRUMy9e6FQDSlaLPLmRlcqbQ+yZo8kjpi/
s6AleMRD0Gn05Ru8usGYuKC76lWJWkJD+KtdRbExtTD20P5/dI8YrOzQx9pK
44YS+31z4nWa/kKLfDhSX9nUhxS1ZhLI0RP49v6u7tLsxfg9SxkwYAq3cOhP
Bq6SjwMG2eIxI4ihPFa1vT1BwglcMXnX1pNxbKiWpwrkHEz9cr3pGdPAMc8C
waVlpg47JzlHgo0ULsJcaqUGRLScklnsAbcpQcT+xEz2lfYm0gUuKMzxiSTu
tYXo2ag11WrtNXbbnVwjI5B6m/0mfnS30U+5CtDwxjiFp8ujXUqQDcrgjf+n
3nLANajhw18wSBSi0NWG3d7Ct6OvkK7qbtufBUVtWDfNrBzXz1aD1NypOv6X
LR0nQhlcfbt7KB/5sYtpxtYR8QIS5NejTVfdrDLF9k2TXzzPETvWRJoYLaGF
3YlTPYFh3fluzYOK8lHdUMDfaOedv43B1SEsb+mNliOmXxgXi4FyTYxM4FQQ
2gIOxySwqmvIUThHhyU3aLksln73YXt0nqzEiGil/kgPJh8yiLlpKAQbjFN6
oY87b1L2lRW5mBzJHP/KCDEccEDlLUQ52qtm3iuq5uHRGCbY+4pcHlyajaNN
61ZQfY6JBaNQAf8h01PctZGOFkNqAdr7KIUixt3tDn0idaaUjtlr/O5PnzlZ
9xqvmPFF3eOmqbOrocJDMJo1mShXxAUjzRJz4X2LzJf1ppKLCCGjHoipQWdj
ZsX3/tsbj+B1v6fBKlpoJhjM0mehQx4VOzjuA5ftTjwYC8U3Vqh97L0tXzg/
jYns90FyIG6ucbPtt/lNxtJfDtRhQnkGF3K5Ai0dZvM4c8BVrYiHq/qup9yd
D81frY1SiDIzF7lAm0GWgwckDe6lz/cJnX57Y0fUfyXv/2i3ODKPQ8B1WjDT
J5fufNqjYcIrymT1vrmeR0znq7wJSZJ75+zam++nPkoBdzkWXEvGoMdF2V1W
CheHpWcBO/XOrOw6h/9WYq3tryKoKNXeQOFZflb6kLan2Kt9SJLNEXOMcIUM
0w5CR66ojsqpJk/PrLLxMFUcnlHGJP+QzXnBZPKTm6oi++7EkDBt4F6eoelO
WC+h6Sb03MMpptmcBWaN1wG7VB/YHW6M7YkwXLoC0zEbVaxhBdbLKkU4Pg54
ARrvHY9TYDRkTL09scXTTfaTRh7V8GNtGFM53PF3Y2QqZCuvSOf9H7e4pFRK
LZOPkiYV2CTJ90emip3qcrbY45Bgwi/Dgf1S2zOa1Is/SQiZ0WTysm1Z3xxt
g4THr4j6HewY1FxY1vMA3Q6ba5XheqpSF99mX3TJcwJpdlqxdV2o+jhMwsCk
n8M0Y3gqIG7kMfQyY1KV3J9nwQ5sKRlJbX9qHf8b2Xb1PTw9Vxt8G8xvOFkX
IooyEbf87LC9Pb+Cilw97ZhbzEBNBwP5CBU2lS4hxIOkS2PKSdYnXQl0CKgi
vxIUlnImZWv+oyaVK29YkZuODgKJBzOj+vDTe6VLUo8Scv+tdQlXMZPvoxfn
DUKnhYKBthwbdmHjzPGVRbZ8olkE2awwx3a9Hb003/rGfzuia6HB8HfOsC3F
sbf3U8vLw6BFFO5ciqbHQwykAoL+tg0R1jNKDKMCJgiNyWA0u1bRASqkwwjv
owqFjy9fxdaucHpOUSIDDaH8Iro/hjOqIFdaW/ft4b9xkIWTwpbvk8lqWksg
QTlgyM5Oqdqxe5wDyC4aDXpVrB/j/ggrdPQLj0EUr1yeSDZZ6iQHt2kkwS30
uqBV9BpBUg4NvsDlIUTXgAHmEiXLRki0PEKGSRzGgp16Hh2+BCM1OdEoQcSZ
OeBMJmU/YxjjiRudwhBM5YNC+f4BqGNITF4M0vFh43rGOgytPobim0z+L6pK
ziB2IR3MV/gEOwq0m1WkL7tN3MqsyiprIN5CD2hW82SpX1R9sxMdJqdjWlYx
Vuqiv5vbKdNVBnu7VImigAJoRDwjh9AQzorvnX2w3gGv4YdCy/fya6Cv2ftl
UUYa8ACv3z2hE0Nq/JNb2BpMMPQXOTg6E6E4mghEqIYcUrfyqHK6dAkaJ+ii
pa+yvtiKZtqmt0r0Db/9B8/KDv51h4s2RnU6+y6PGkhgOo7UFI1svQWqL4Ve
OmKdQ9qJPlaGR7zbCw6ed3IfCeUR/3YexYKcvydIEAJrHxeKINoXJTQz+g9y
Pl/jK4mJgTVIxc+jVFDS4Z1SB9YOaZvtEsqS9/OoH7Q6NcvV3BNVvSc4K7O8
fo0ulERdH18DJ3pyHXL0lGLni9/APSDLdc3jEw3lEMtMVcIq4Rv/LPVt/mJ0
BlVC4NmJ4apZiJeELAGs7HuFtf0uovOyu59dJ9/1YMeulu86CjscAR4QFIdV
n8oaS7Q/XTwcFOh9TDXlF/+vKIqjiah/zsoydAZLSvEB1LGbpChsanfa4mre
3qwNG1lYKlX5NM6aPznnlKq/d4g3QZO0Xm3MT4sfJZW+LEWXa/r7k6JaSwnA
mLyQrqseHoMDh50Nq0TIdiHP2bZmy+J/lLLcQ+OHiuxz+ymPEhTQbmvqyEDf
viMZaaZL1PFBw9Zeb4m0Vvxr8/m4oDIndnfeNs9QSAyONsjcAx0PPz1BnJQN
G6Mfb0/YppvCMSCPV7YH4ju5RiKmaOVRVbOY4sYseB7adb967v2d6tcizpw9
ToxEJ+mUtlzpLKDHrrqy4LxULAspPIhbExO5CNzioOt/04dqW+HfYlY4NJGD
keNDo0i0f+BkhTLKnpwzUQOGhLF8sKkxGFS8/bHryCCpaprcdntw4I0loXD+
Gl+elHE8lpUMRR5gvSMs9oAo4xSz9Yt0yz/fGY2OHo8Eroo/EU4FHUquDyaG
kCC5njmwaNH1BQnzEpxgOhL3ZcTa6DoP4AOe0aLd5Tsz0qGwhc/k8gMVTRCu
RDrsrmh2E/wkDCiw2rlXfTDyJ3ylSc7uTO8NfaSbTynbFIr0lMDSXhTSXLQ6
mGETjx4EaTTmCliUzfv/W7FFs/7k6Q20d2zDng34y+gWBTUy6I6kqWVzfIGw
PjhpTUpV9C41pwBP0aotx8aKJYMZYxoeT4tVybaYVRANYdmbkGNHCmcfEv5i
v6aAGb2JC4KkVxokCuukovpoNERk8cDgHR479RqsF6JXiw/j8FQ/c0NWnPHr
6N5WUzei/PbnZpjWe2mShwkEhkSEcyJEE2qTrLs78HdKmCNBIYX0sWBTQ3SV
csD+FiQy13Tq/dNOByDPHPy3tCYKk7xkuQD8/ODZo8XxATGgElWvHy8qokUe
SW6v3j8cJGWeRkF0ajkwJG58h/ovL/LNyjnFulzByZDYv0wDgsH+GoQLbgpa
/jz3Sill0DMakjtwY9VNGRmwMK0A/Yt3Q3SgITIYvhrD+epaawopb1q++RQZ
PTelJcNVeGeIssWES3APNGVTyiGsTDEyywvWzbhawKmnHh9jkElqCYhIJcvm
VO+CZVeGQOTK+O3AFRXJcQw1DbI+gI8xUHzuoeF4qAmDwubvD5YzkgRDRNml
IQPCKW9FQndwNZPo4mPr7E8ZBzPA9NiT7ANlrV3yvwcrtdDsUX95VdyOq5Hw
hQb8LVUXS1yj3sDqctY4V+LXX/4Ux3csZwq79SI36+BK5iKeFXf6z/I4KjE7
DqriJT3XNp+j14dYAqd1t8diE2ZZkYuos63+VrGe8YymXfrCjGqCzyW1dbvx
CzLtiX3o05gkRY+0kxX017U+wp0NW8pywGuauAUpRCqd2SWQ+XRBpz6Ayf13
tbQPjRId8XFXsMnOjAgBSyBUmn5ihGI8SVzHIVVI1YgB0kqkYAIOOgJOcluu
ahlZ0d7iwLKNGvXm432t7pg5hRlRHfGih+xLl+MoecQbmA8T6u8PpC2BBkz2
KiTU6q/8oT7bYbyYWITaF5apr784WNMLIORw0hfLwls81CH9WDEgEL+6qbSW
pRYEWMa4vdYaEIkcHzmOWIi6SEwkfxqV0loZ5JZgSPk2Mf3sFZE1d7EoAS1R
b17mSo7rMdmPRYMOMMS5l28ZhG+C7CCu9ojnzzoVr9vqU+PXKgb2BdYoDGFd
Koljb5FtcWo2WN61jHSKpvmMIq1B4oMuYQMVsSyQcGPyRetSEFTnXceYgKPU
wqGhDG3HyYC5LMpGH3yzsggRTowi+TUrr5IHMoxBNCgwOivlrKlQqc7N87dI
gtgPpKUoKJiYLZ4CdgGsE1tBmsPu26OO9VtN2d30hzzw9+WLC154rlSDJ8xd
/v4sSd5tS1aMfjscFpMprUzBDq4+RHVCbzYdlDZwO3YTg7Mju8yTVNQq5Svl
8DPr02UIQ+QYbkvxWZqpZjfl6gbDdshE14Qj+DbNm+8e1L10BEnfYcLf5eCU
kDwHq0CcQqTsO0YAy+nbHxiPkB8rWK544T0EPqDdsu2GgXpfnit5acFKfQU9
ibrFLG8ARxJVzK+WT56wSRqlExVN+vt2TA1oxkrJ7hIRpA1Lr61HjwDg70IX
bGBpl7X0rVA+FZZnotPba9YKl33PceGLGu/W33/gBONp7ZyMZh1/m2i/bpJx
QCGbwnb4OZhrVl5Ud+hnb5EEETr5PlQk/JHmNipzhmipdbpVRAUKBF2hmX4S
tMjPWKGN6trhOtiymSheQWfKEL6H7EqQjx5+/S58wGlBb1ipn5VF9MCPSwfk
OJzLc/XtsJmihqiGuykKNHaukLbLsropWNsmnfi05addADK1HczpV+9lvcBV
H+iFq8Ij4oniBG3cgwmimVMNlFNuZ7SZ9JiltCXERx1jcaykzO5TMef+2nnR
MhL16Ktsp20ymoQzTICTGiF2owjIWeYCUCp8nr/aaAjbc4c85fSVboMXIx47
dyfuNMt2/q2SXJpZfgFHshylDEda+3mYcbroC8zf2cZpCzvIlou/8HDGV5bK
pCz+jL0t26Xohi+7CweZvAn5TuGdrz9eKosXSSEq7jJYSzrTooyKP8v7c6XM
XF6C1i3OYT0c9j8bQ+KrafwopWz6JSKLnYL3yzE9Bnv8yZZCqBG6v2UjtxFX
NJ8ZQ/y6y6lvHPUPY11yYOferrebuMtm2EKdVsUcojfRqnlJCfm0RQsmub+9
3WPeISbuB9gM/kOB4jAaglj3UucXfV+EOnacr+k1k/E1xT+kwAxCl1pAls98
0qbhlwuoJWHh3aYCiWcbLgABpUKNg7+MvH9URBQocimRLW7fhW5q1GVmjjj+
NFry4xGTUCNCyDVW2xWYSETE0ZBHzKFXxyfVCHcXaRqdJlm66EPVYtoo2LQi
ICSN6wbZktbKn5qy0v+xDiIY8U2DzeKo3u0qAtq10cF3W9W/uNE95vi7zjoI
bxFRewhMxXSRLR6k44RuS/pgL72b2NNmau7lmZyo8EaQVP77JlTE6St/VxPd
qP5juN184BgixqKgC8NnsUHIcbNO3Q+to+TZJBRfftilXALeImsVg5vwieCP
h5uUsPEH1CMOoiSbICpY7cw6e5a3NHQrwD1QqKJ9PZIeFI9ei6xLamHv8EQo
TFaXJobP+I6BkVH5vzXcQSYSOqRrDnjmDmcWRDbaNFXyXT777itTqxAYjCnK
Ttlx0q/xhes2mPnnyjo9Tj2uiO/3y+PBdvfsUN+i+3FNcdLNQnY1Vglr5LVw
Z7/iws0ijIZFAReyuZpHAy2JZhNTItDVV1T+6Y3Qh+aMErRuHm2KFwm3t903
ajfLWASvqD4jzXALtv910g/tfEZ7M9PqRedNsolaUIag6wXv/LlCKi5L9uZQ
qd10BzvR5BN5s+axzyVLfh/aaR93AMckZnFGLBwje/GlqMZbNo4wHvatFMY3
uF/R5i3bWmkhvHe/FLfSoEBiZoDGH60ceXUEIktGK9en2gf598knbs1PGntK
OAWO3tTe0aHFELOFJderwUaawgatPYEKughwX280aBexlUdgI4XNKLzUL4SU
+8D42gLJRUT9a9Q3aaG3oEtX2a/SlKhTIZEyd1IKvWNGZg78ssVHuPK7Q1c8
1Y0Gwyt8Gmlxp2/n9mxIg4rtAAc2Ti56Gy5C3kdA4Pqp2WRB6ghLaKwWy5Bm
LGtjAY4H0MGlot9ZZwD3dbfS84D2PWRTKVVYt61lJIFQNLS3A2BvTE/jIS63
s493UF7kTSCsZHEyQ6zb18YFbg21Ao9GLZr9TspEvYk4rzE4FqwcIWvUfF8X
s/GWYmSU4LKOoPsV0UIUPwXk5ZS/yBISdDnSVlpGUcjblHWFzG4hThnVkvia
mUPFkpMOMK/FGGslZd4SoJ23QZv2rT8CD5UsvUOfJnbRfMvA7QYCFZo/Wci3
9cRj/6/heKYMJM2N+EIft/aRSsiXEjLj378eYWKEgE8wCNsINqfhLmL8oKYr
gD8EDqDCxerfaGFYoLHnbC8Y/aql33145EAITF5iiLwB8w5SB5fUVoDo7i62
hrBYPixkvkKL+jqPDd782brVmG1XUxJAwqBvonyPmyXJ2L65DPcMLf6QSoK/
s29N0JPqp+DfzZKdQIHciui/xvFh+hmknjkVfnEldwm4q8Z/+PkCGc6560r3
2Xk+SLKric5n7TNcL1OoQEQAQ38bgH98kfk8nFhqZBvQr8eH3TjPDY/PrfBV
v1XioonbMWNupHaCZbJhubwcUSsISX92hrEC2C0muYazUFeUTyZjPApr1zYO
y/PaQZ5d3gIDAwxu7KKKcG9pMfNG1IoahEzPoigAGXTFabKbNAm4wewj2D94
NK5NKAQoiJGOqVWzbE3UaToB+99adv+SbPXj4Yevh2dQWIMAfysUhh8/DfZy
O1HS/5ELMp7RjBPL+NgPVVhzo0s3b9hD8nZai/IqZO+jejbbscL1xMPZMXui
uLANrmxwDaTtIq6q9YA7IBAR7DGGn5o6PCvJHyPpyMTf8eqaHrYGuPlNRy+N
uDlfpirXgAgjZWpRL83gJjwxHZpi+P3Lb70K6hJRQNfY77fAqBR8TAAkCo0f
STac2dSjw1ci3ZXIAV0EPaU1BpwP8NtJrE5kTd+5gA1x+VIHLUfSM/Y6P4re
nDXRW+jKhb9gDg3I2NGsdKjjF8WGmvQwbv/Uv68fvQID1W9njTTLlBroVte5
WNqQMgvqi9pEgfEy4yl0LsF+WA4UtDyXpz+vY4cb4dgaS6xKA0hBKZnT5Vjt
AroQVAMYyWmAkk4syFIBYkEfRuRXe74Hj3T3TRjIL53UCkdfL996g7TARViO
kryQKu20gGDU6bH8bxwmLjfTGAdDAj3ne0x5DjHU/vAJsURfbZGHb0VLpM7E
8LxEgfRy/1g22RrHIOiFL5fOBs4vELj5o6ZipUdqsvK61w==

`pragma protect end_protected
