// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XymUfMqk3IYdKrRh/PFFkLbvzKhsmMFNqsoRy0xBR6Z2gJFzRL2zegqswnL0
g/tFEF66ricNjGdra79dpJf0jCGHvP8hEXWQefkRHiPTFbx5wzxXKa5s9++O
zhd7UC4cxjCj8aeVFJVOIsxXjR289XH4dsDGTlfr9UeIi0WcD7KBc0nRHzx7
RgtIfITP8Fwl5AmyGj7BJhYpspO7vHUfsMZxFyPf+r2sl53s0zAT/tWhJU1G
P7Smo3i8ExjlZ3YlksjC1BFhf30+8NpezuuHaa15fSxtAhanbj5zk/MuUlnD
4StxwX4KDSKPkH9+6RS1Ne9zjO6j2fnRmGxQLmhbxg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oKfF2cT6nsJv6uTGfEQKWLcVeqYTZeYNmCpd1ykSZ31rEQ8sxdi3CG0EaU4n
ia3ITjnr9y5oB94yxQ69vMohA/m3PHaMYKClrIT6ZkgLnXisutJ/v838cRFE
J9KwG50pthu9VMVdB3y3PDLJk2xCBWPf0ugXbH/ZX5Yp/TvBEwPew1RHf4J9
6wyb6ETYqB+Nqg1L7IGFos+CEobwa0wBmBaLCw55sjHW3+AJgBCDvu08NO1H
58JmYQpu3ilhUByBF8x01d9tOPXYM2lqy6ll75K/dInbOFm+c1F3HSDGfhoa
fUhGSm6nWu00jvqyvZcjaeq2z0J6NO/gwG7Yaw+FKQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ejS5UwTSt9xeoJEzJASgOEVVM9Nv+U9T3gnxxRNbV8xVRwIa2uiWi8GmKMBU
SoTRimdmgKCAw4vf/0Wm4uAwSVfcnFT72ezJ4HrJgZAtD1kLSLwV1XvQCLXZ
cB5GlFg5LEOduRZjckTRhBQeO+OM5CBKd4QW6MWCeK0BKttCWytoujTjpza7
KrhUW4K/hHvZ90ebrDhrm91+z0/e8wH4cUG7Ts8xlAUwcIuupiTFlkcexuPW
iXipCzTtPQ+ZeKe7l5wqpSraMExA+4ttF3lDB6EoBCqumhcEHzGNZZG76LtP
Rpk+WIx6fzVK7A3BZIt17hs+WFIWzvDZWHlMwojB7g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Sd4ZfhR3CtYmPieFnMKlquyakINCJt7YwGwagE5khNHlPdEc7ipV6vbTyHyP
OhmDZmAhqeSEG3T91KBb8l/0PyidhO2T3jIvzAtVCYsVCgrIwuEEut1Egqe9
i7dP0dcX0obrysvSJnBI3NDOW+ICkzNHF3oFE011N7IV7SDbZRM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uW7goNTdurgeA1RBKEdN0IsgBlLxkXzBBBQ0Yp8HNHiDKbHtserwkiawytia
XQ6KOazK+lqt4I9C2A2yMt3hnkiB00XyEceN582RHdTGnh97Yx5R2pSyTK2J
OMTLdl5N5y+26Wc/Hr/E0ZEKnKpiBhKvSUCqe8kZeIcA4gF8eaqN5XnZ0Cmn
B96Q4dQSqYI6lYIndo9XTLWYk3pv0vhbiTHz69/KYtj+ZhsVGG/ngCJlHBEq
kvQkmIe4qjA4sWpo9iYUsh3KqgSWzTV5nWX+Wi9WKsiuPiLpFG5XkxfHIafR
Q1WiMSMmpb6SPKvkiGbtpCNAp+i5iDh5rA9dSvzVYMK8OUwy+gumJE/BPZXT
b6K7JZYRLFY92FR/VgD7Klan/K0gxdkX8qeXQXPul+fGktdAPBmvjxDb7B53
dni5NR1mrXL0hbKAzKqEiyXS/7HPMKdFGeGz5cDYuySWUPSSgtOXkF/OI3IQ
o17EKyNANLInQmwNzcjaZBBGxdx2RkA4


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
o7yHoEyWuE8quXh+jCxYsUNgkOvePghqH4IsdMDTRcjrUJdmtGGgaf83/xaT
fWVrAH/1YACJu4j+DGsjx5GylxaWnEAjeCyfW+eotyuKs+X1tkjXSZgL9xog
fga058L2GZhZwLoklqcE4xYbpuWDfeIF4hq2mW8RCnUCpPYCg8o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LGs3eitgIBG9m9WOjzJuJi8AS7ixQoUchZu7UkwBmvW9afl/UpSbnqeB6Hlx
9COv0Xs5IHSAWEwTVaj3JcQHotjA+cZ2V5/hBqgOfKLcR7apydacagyEBSsM
Gu7GG2dBJTylGB7QTCoiZMJMHGx0AbKiGw0omRAodZR7SOAYSk4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8000)
`pragma protect data_block
5x5uXQTkJCYeY9Dw/l9HIuMMQ6I76JHJ4XbolRjesE+ftDvm+zuuAEHOPJwf
NTlH7du54KMOD7Fee02BC6soEeFw8buG1muXR8q0MnpRqwquQdkcZwYOQi6d
hWgwcrDlB1Q8QwHXgCyCQquqje3wtRDCn9Wj9eJ4qMRBTk1ADdj4N/BmsYuA
H9Up2ebArtA7rI/0XDIpcMpwI/9HDv4/JIEByVDQ+7olBTykL29LEqsW6MSE
4jVBfg3clTDbgew/ZuNgMTqjcnKobQ9wFQh5LYiG26vC8zMLuNmp4UdF/Hps
G5BsL+qr6vS4jquyz3TmxIWqdtI7PulIt9DyfqKfMfGOAapiwBXhMZ7io+GY
h3a21SQHdHYRq0aXX3fmSPexEwTcF+TFx86ntBtuAXpyQVtPLvC4DBu3hpfn
ZYG3eWkG5uIaXXr4yRD52E6mHf/yTxWs9OViyb+/bFiVzMEfC4xI/Cso5fNy
0XVvYhQSfJd0Tz7NlIubGfY7gGZpWv1IbzmIbQuWEo0/I+R3zMt6gB6++b6O
6MlgaVtfHlUo8oHaViyBVgQ6UKvwN+H7kjZHCMBrKI9fFzVvutB8w1XjUV0c
UG2dlhjtWb1Dtbx+zK3gQn3yM6/1EyKRKO5vj+81dnpcmCTvwMHeYTnSQA5q
2ajrCldm1rfiGDghZMhBAQCtkhgSiI8kOVqjO70AwhFwWVgRaCt9lBYS/d2R
i0BKeGRqc8tZcb6xLIu8vfPcdYYztuxV8or6wxCvYlndNPoKsRfcFzwfqaUj
o3+WUmkUKYASuRZULy7+5Qc2NPbGqvpseGkoNQZbtI7iLIvW1XJXOvwlgOi6
qM8NoC2dOQRMaSxmbqDEJNBOyuQrXQYWxlCp+wbk/OBzh4srCREkHjU6SGtg
IUogiz3oaqzOgkFO7SfWtkCudfs9QSdXR5Zz6jZCopxVfdeCuwbnZnScp8/m
T0TQXJRhBNiwIHkaSZvmC61O5Yt5N1vt/zvcKJuJ+xnzu35cOC/y+KMjvkmH
OfMGso6XTKwV/bo/9NycjYdLPJUvlV79uOojHq90U8fzgODMOp+X4H0UIlL4
kXj/1zqBnYZ1AkRxiYoX3IJi24Nm597KYEWAac9qE03p+Ss0xVgYWq33++R+
dX1XChe1nV9lcr0Mowu1SYBMudtL+vv/gk3XOr+YFHj2lOLg1IAIgbHj0Trd
0TfpyBezppM4qYjoDoS9wiZ4uBggaG+Sy2JgEqTlYjiObY7blFiSrWNlb6wA
EbUWHlTumb7MFmuWaiWKKCBJxirQHAvm+mg5DE5Zd+ArC7shI6m5Jh4NH3s0
uo3Fh+mkKUAnrglMGcoj7JtiA+YFnhUUxutkVfFEiPzNbCuBtuaMtEvt/EWA
j+7K7Cw2+ZX8IdceIiqWpp6xqa0RiFS1wFyt6yLVBoids2c0smWEwGDGB6j8
h8QoqRcyAL0f8/tojNfqJLXh0QS4Q4VHoDSUTGqxQmsqOINKN4mjkn7rq7Bb
iaIj5z5Vu/3KSvBACdotHUK81uI2oeucPwr47Htnv0H+RoB2zHEYbBNJchAA
exvfDs9VCEZEVjxAvmDK50hgOUJptBXkSepOdfJUVSQ7aV1ELRNoxq2o9sfD
WJAqjYYFbziiFwjHQSjaU7DKbmCIuE9WV9hNKhrOu0lOdBpv9CS4tsv70/qc
84sCv2eU3/M0676t9tCaITOgAQzQyLj+lKw+ANk58SyKSs66VvD+X6Dl1EXE
xTCgnl/EZrUbyG/bs6nArg64kVQr8QMf36x61anHQ/PPq1XsI0miMSrT/dsG
AkWzen4zHjCCVf2Nua/Nep+4KmxSDAU2XyqZV1vuXG082zZbHqyO0CuZ3Vr9
h5gSVrv1RcWohINJDzda/UOnuCd73+GGBE/83JsbX1vLnFPwUcb7CK8YmtK0
X89lvvTWI/OH8H7gedP7Q7+E903+nP3gV3yS67t6F0V9Kx5Oj0ZISn2ipLxr
MQX+KmdKawOXfannZejcs3+zad/azbWvI2gv/84SrfD0TsBQ1lTOGpJmicFt
Om+V7NwKj9rKs+Q89q0gcRr1l00U70f6tx2RttnoFkF6ksSegN5BMqWigQAY
qmqQrRAmt2U0patxYhLPaw9TgIppGPjJKUm9x/cNloBFiS/4P+HrS5IQ2QDm
h5dszMpysUXAT0MQWpRiSVIoW65JLlYN5IwsqBpc7hxy6ECytelI8P9fOJKC
wYqF1bwu6eArK1Fx80ctPepe7rHH770IuSutEGi6jPAyADdBp6+Q53aJsJTn
U2SAzDckacQmrRVlQ1HL9c7VYSiyUoTv9jlpUi4LTQhxglZJnVg/1PQXhFSu
pM5gYgKBA9cn5y2H6evmCB1djcu4hcIfaB2CJTAmYi0vo63/MsQi68Ovxhxj
FBH3aU/ClbTZ7CD6kjFzDH6UqesAPPobSznZmyDd2RShgEUoKqYZITUF0brC
qwrz+CEvzt8J/yEtAj7TMUjE8GoNOrJZFpPFQxR2thQieLLP5/4E4HAw/Kdl
DgJIo15fpTLKyF+7fbBpe02MUNFcbkWlFDlf9ik1fxyDe5iUh8/tZPENNFS+
W9Q7siUfSlsuAzsvu26MTF/opX8VtllMOAnrFaF9ZXSEExlIYIsWpV9Jnc0b
TXwPdyhZbprTNTNtE4hGJGx7MzBiHqRxT0+6K7FN4LzpxtBT1BORMzvMyado
oE9G/MIUKtEXKIUCcfZ9TZetvBvWbYPqAGETjKCGDyKyYJuO7bVPe93RCKqi
m3iKZqY4G0lB5kiK+OwP+FT3Orx2Tbfv2PqAc6m3tVlLoo5mTe9oMPYJDQeC
MG97Zc1a0awzLBgglZNIuYlVrpVrf5ysmtMZoomPTayhtn1MPUSRf5P34rsh
zCXx8x/AsXuGJBewke1nqG60nNZAB1x/FsWou8Lpy7J181MoOsawmLFKpHVz
Yv+lgeC6AFbEjcqnX31LE/CjgQiLojzQpU2rwO1kWeEPsZDfJKwoWjXTlTi7
YVe9ksvNGf57yfhYs330hw76vXxBWLKnC/8bTX7HA6VPoI1C937lVTA/k9I8
BMic+FRo7aLmIPhWLEyjvb23cHZK8R/R0UghTTcJ/Yzj53gb2V6mWyJqLIpi
7ZoJhMvzXOhcd09zvntDHAV/ZZRLlS6eDNJaCQ+P+zCqwAWgrENK4SUJ0Bnv
jGMhOgHXJzUJMzxtAXuJxlO++26IoYyiVXFK+k6XoWk3j092Ut6YP3uBnHlc
7sur6ftTY2Zc90Pa5sieAfmZLNnj7GXINK+rRuFL3swu5Rx1ju5f0FXmgASN
WKU9vVHZW99GvkrDJvotuP9AZNBlERDVx7Y3T9W8KJZSHTDpqIsySVCf2GUi
Rsjlla+PeLo+NGST2TRCHHy6HKO50g4Ni8dBkP14yZL7ki5Vn8JtfvBIPQuA
yUCa6a2SO7dj8amcpR2tURhRRqXHJAc0QPh2FkJIwIE6/2S03JZZqyIENBwO
a+L6uhH3I6ljnID4RHVtkU8p6TbHMtBp6Vf+gAdX6DKlXI2vDqDLSoxrxuRP
cz/hdKpu06JGNGC6f8FqYQBeWaIDlsVdQSNoDshCHTL+jjcf8J254F1IWShI
UKDEPXnQIxBLH4qTKftsE1Vp8IASSsL6dC+z6EesCRBH7ae4CHVVOHkKOBVW
TMmd7EBWlFsvev2G4xOWbqsupkRcQFT914taEQFjWEpdO8YuLIOwZKiuW5R9
sxiMt6TieC5tgVNCZcUsBxN7Ysn0Kiz8nfXXq7mKfLC0/wOKJrrLveKL1pod
Eo18ATkcSFX58mypP69ySUlq3qe+VqtiEEacNPEsSAJsi8Rd8Ruw90RzNc9U
KRIl9dzyjgEE+X3klTG+DEVNDMphFiVOVUCRbQ9yaq5FNSIyJKL1eEbsXfNs
WFQTiJESxcnsFSrJyFVT6f8FWnqYgDVpLR0/ew445wKbASbqNimGjEakbye+
zGt4dJ5pDnYXy3DMWy775HSzccAIWX0/NBgVoWlGkjSVpamoKLz1AFpa+xZW
doNczPcl11+x9F7R18mqTnKDKeW36S4qJ/ztF3sioy9Zk9ZRBWC/kDv6ve/E
2TWcT511dNfeGceuRys33ofm7RXE7NzhqIT+Qxivn07b0GQj+qX0rdiFHmEw
ohAQ0GIVnkilc2fmEBlJqZkcSyvOKNI5DH2SPW1MV5lfhDmAjJF9S/E0LaG+
fpt0BYsuWFhqDOrJ13rEqTTmYXTWul0KFJW3c1A1TAweccg0rqiXlnCUu/P+
zBkOBABSgZidGEQMftA9VoELKGqaQ0IzO0WdP8aaWqI7gC3y505JGe2JnW0/
8cxjeP014KblAbHXnTYCYxQjOj58M+XPXCwuoW4x8QdQu6pnDqJyGOc1LQKT
WTUAn+1esRUJcekzubH/f3pheYFtbDUXIzWb7xEJIUMTLCCgcpm51SEGWtSL
NwIn1hAip3J4rmGBEkg8exVp2DXTnKmTWCamLQprFcQO07NqShnt2v1dhIR+
vU64Bpeufic3w6NbEAN/qeKZ9GkEic3fSkrG222cM8Yu03dkAYcYbNYPUD2t
VBvrPcIPcNXMXCantgoN2hKMhJ27KSFFIQ7XCTyDCPlABmwzbpdEFTyK75rp
Ch/APG9383/Y7uPc5MAaDlvTwmGtiGcL3HDp6B+MfF+ZLJzNAQxZ5I9m0MTI
4aab98i6FFW7dh/W6CkUep2H0/LhuMKiICNOZA89ATch7NMHnz/oNyba7Kt9
0yw5POZ1wCbOjx8m2yNPX+JulfGe2lB3zRiegWLZPRT+jro8Gdo1mCVpwNE+
txNowaaY44hUKwVJUrD9vqWkAITKrSupevwkt61KqUr1wXZRBHJJR+ve0I+5
P4Q7LN3wt/xiaWETdf5pwBgqLvzvUSO/X37BIWptd9w3jW3PS1ZQE3I9cOUi
dYVEPuT8OAy3+pB15hmXg16/n5BU6MV+OlQ6fMwrEIe59jwdQMQ8YvViDr+A
HgWbx/do2PJJZhetPHemEarS9xQMcz64xFveobVGMVgge1UnsUos100n+uIA
xgkiwyA12Ujg31Dert8CKhJAn0CPzz399Uuohbu3Cmh0dggMaR3MgVl8IfZ7
6Pj6q6KwORNYJrfZaByQ8ogiSw9mgUjZcGYiJ6aqqzrcI9cLb08vI5H05HDs
7+IgdCCpjHHsl0q7YBf8SVizvbryUNeLzfJUxZRDaZvZMpGMqf4ZxX3ZgrJ9
1aoQBCcMr/L8kBvla5p+2VkbVilR4BW70Z1Ex7J8xCjXoy73WgiuYUG7Igds
13l3xZ4fU9GKcUazcNU/RCjNrZ4Oe0U9bWjv5CuXNCYo9U5e750b+jyuUfmP
8XNgqVWrpR63YgGyuVtw1bxDbNgWE1YX8hukgc0SrIpMKNbhOCijE2C4A6lX
Z+XIVinVzqrG1qRwhqDK2hL+TutC86WpLG60HI+gDMdbZLQGJjnowGipF9l3
cTak85OpuqkfAA1KYutB3cOGH7vT9gCaENBEcsYTTbxlla/J/mjhzqh15wwC
P/nGwOE0BiLphYNs8xGFQuQqRYpSwO2sIArkJNw4HgMTxrU89DgBGIwoaxym
Ojxf0WBIUaZwSgjm5a8pYioB/aiRGg3pSCS3XnipVOOR0Cu3jWwWd05DDpIJ
rXX3tZLe1t9MlvagMSfyaKJdIbdKn2OBKOYEqcXIUOI3iosXwCeMr+nmzgFe
PPemk6lEYXPOK+Xc3sxgBfaQnhZj8jrYuAojBnwStR7tzZlzybLikWTi3bsx
2B2t13xsrLV6Y4f+LSy6C3okStNVZpJhRvpQlLFBI/pqfixZEFFuEcZnYWfo
Mz+XKyefqnck88omYMyI16BjzdFQ5XUZNg4LItYqpS3DYwmNgjxFCUzTTCDI
nctuCR9/5SIqvT5Op55W0Zd2OB95pz1DMz3vAg1WP4uWKzT5ibWqhJzYuNkL
dW9fAxzgS+pJ8Y+CQGbclKhy+QZf94ymjTxgB/0jqVj5INCTsA3qXozpVLL7
NRb2EjxqyFDCksMIyGIZi+Gktl8cve+Sgz/O9RlKJo/q84qRsBTw+RndW5tS
H0rguMJWkK6sdRqHJZsUx3D11gzDO4IrjrmDE2DhEdbNsB1qk/qgVImr0x2J
8CPh5loIG11RDJni1CiOhJGF8nj0IszSn4LolAy/7zRjw4sdQr1EV0rmCbyg
19IiCNLcFAaJ0ID4jhIolNwN5oEpXy2tUMe6VijEL+6uR8MSiacaqjltH/32
uLfoMs3/47D2/z5k7Qi6wKyz7H+ssC5/U552YRNNKYIUL4UIfQPmDY3BpgIi
bdijODleh8/AxMED/7XfjHJj/K+F6Dj177JOlL0Q5+f758xLzE7jxpGb61qb
mtW5CopYAWPnU0TR5vOhOPc+rZWFyZxsWG9vyPOUokx8GSQhvBNkN9GMvMaZ
9vVyux4qElzTXX91/xYKcJ0d/q/8uVOjGUsIhkxbItlPpyvK9XPm3qRHdqrB
Gs2gXpn/bDR2VD0YSrtA2upqBV5niwtP1k1X50KDC3M0P67iUhHliXoR3qgT
XgZ6G7FXL9k/afeCRePYlmys3gUZORyTvu8Myez0Kwd8Amgt38tnhBnB4e1i
VTYszSV2UaCMhTkMOfHfKbEDJ5nciSy4NPt6ig07zRjwTVaCQarPL8DMfure
NH3zQm64PXZY+44D3ED/Ghn1iSsODQgIqq3CUR0k3A2sJS2txzI0v9mcACxx
6vTCT/+Z73HJfM/9xf7UcsTsIWdUwOrvC9mX+ifFCcb1+tIshQIMHDnoIpuk
W0hm1dvMKtmHSnf6TMsFe57hjl/UUR+gqtIHC9m9o1dK57fvTbqi1sHVieZH
ExWwxjwRiZ94gW9WepxCzGhrRW4sMC+hpzOF5vaxX4M33ZwY5g7/HbfY+Iom
u3ugmcUZvXpm5+EqzjOROU8v/Wd+3KJdg3Bj5Q99O7mY8kYATCIRRrQ3TPey
VTVPIrxV3kIdEqcnIIyB+AwA4bWREBRgC+CVNA/kjR21X2+WSr9u13ZFBh/T
UEJqWGJrBDHIRRvV/aGL0rNZyfZ9s/RIVeQ3hcNfo0ZjiDu1KFGVcJQflsdR
SrZY287+si4pGaoSE8w01HyrOVm0dL8/B6pv1Z0Pw4FpKQV48ktMa0l+js0B
XxwPdl/n8ZJnwkQ8ba+mYQH/yZmnyYKpB2724RLnHT997p0w6gr3vVYc6Ukb
SiEInTwvF/tXrTPhnkdhH2oaSmtgUk4YJEfNOrgl8dpoI9diZymZOp44o8Ni
+3lll88K+Jech+vsecKXnQIc+cT8RIdKeKiFuUHFCK2CgbV21wjTR7brdQXS
vAmvWYiYsyQjk1bztakgsuoZqUpxnuyqoo1ICM3sHgpiu1UoZeLvWqrFbStM
TLnWnpkL139vR2uYPSMK06115jrmUkdv8BhuMx7jabFc/lpQKXLWR2MyGKkh
X1qs+HlC61uikjEP5gqLJZu/X95iTWownFkk3MYvMkjibzGhFZTZKLFsl3kv
I6GrFsrVdCbmA4g2Ordm4KbZq01Mf3iqMfxPF2gpSgjrHxM/ih/6KgsLK1Rd
KCPR0UoKAHPuDIiDr4KTkoGFfveq62aiU+j8tegIFRucS6S99s5BKFglAFXB
E9/ot9gebaYi6H69eHtuNZ0k063pgn25TZJgXUOJ1dVETagwmMO4viZ4xj8P
AyJ5/EtmCmTgzNhK1+y1CqTMzTkXwKg1mG8q5chujsuXeb745hyGOmp0NCyr
a0bIRRVQxTrstxi7LFrXakdlDkbb4iZWgwaXxN5JCwElXQYQgvBBhghrpUJ8
AVUh6/f0TmF+NzIvonaDmdp5FbfpWwbPXeOR+iGb4beiosp8SVra1dUQcTsx
ohhOYVvSz4HuujTNrzOSPbXIdLUzMjOZEppqF1HKIoFpfGRQiHfsnsubfT9O
P5xXs0gFLEnShPPIFqbpMMBaV5N/AjaK50cJC3oxB0InFp5E+pwmOpcz83Wh
N9qNqjtizuwZv6GJRWSTMNads0+CawWyUiC++ZK9HPBs6ktRCye1odOPjvRp
LktqzfJ0TVrfkRufcmNhN+2dbFYYI6PCDjVdd9MhomV0ps+6iATNuth3e4th
R7JAeCvatWK3H99YwfW8KncZW6WSIMSmpeKcYrbn007siptkqPTV1a7Beq7c
/6aLVlclO1GVZJBBGsg7BPMB0p9Uydg1EdtD8Q8Av1SytfJjoDB3AlJYLR30
5uJrXHS8HlmWDh/v7lKYnKFFY7ruvXvhTqR1JFXhdSPdWe+QM9uP0U1NGaUZ
NlOQTGCaVdqwScYJCkoFu9X0AiQH2XHtnrWyZ6i4NKHF78aeAttM0rvRPdVR
ZtZ0HzsPwMl3ZvozBvLC2aJ/KOndQuyFqqfCtXiu6kWRkl49yFGV9EQTsFvR
sCZw4M558H0xd4BH/OKn7rNO1IvFPXmzLu9YSEDMsutR3E97c7cf43tYzOdu
doIt1ikJqHDq4LmudBWD5JaFmUFj7uaeve8TjBPj9Ojpu7ejRWGgs0DlZq1b
CmNGtcDjFlrlvaUPjljDSa/aJCiVdfPHrsYzvFHKtGT/eOImFp5JoSZYq0cf
rH/qzKskMh6dWoHKq/84f913zZBBuQU3ZBB7ZgEFypcWEdXMEAjW+PXpg3d2
+rraPjNfweqEUDIOOHQE7dUhTXV1OQ3yQEGF78DZJBwb+0Ji/uM6g7Zwr8yd
qVaxVZZvkS9qNpM+CCXa024XjSfmfFI52qGySHI3DOIj39tnZrmvgRp78EOR
kSpgqTWIw2/jrErNMlxm8ZFoi0+K9jFueeEbpn6d/aiqY+S/tqld4xo8A/hU
JbPEOLkUa3zAAZj6q1lyKdO2As3+cEeR3PfGwmzKeA2/BzMogzp+AUCM5gQp
EqUeFiyZy/oxnETDRk4Iq40ovxpCgNOx46lf/7I/jYUfQAAPpJ4f3iyo/GJN
H3V8d4uvOlVWMqIKKzAXMWMleYNjnip+IeS3G/c4VWhho7i0ZLF713YPKxbK
RMAmN0/AkrUuU5Dj+xpmNSnusyhzpI2rY4Yafoy4g52kt3psD4u01ohzjx7E
r4cdA88jkSc/chhvuW+TceGoRzS546s+0qelvy12qyKMryQfp6HjX/r8O33X
Fwdzsc8+mV3kl2D1s1B8dtIhuPklTqViwoajEl1L+FedtjFaGmPKGR853HfX
Dek/fBsXngsf5IJTnMBj9DeQ0KL1M2zWV7786sUSE3RFUEolLL/OoPtKMtiC
Mf0RTJB5H3JJwznds6HWgxgG8SXoGp5bKlgRMeyRv/+iY3Yc5RCIWArzTWE6
hgQZNFAE6/Nol49WK+7XbgZrHkUAn8y1CxZzeZw+yajYHt9MgJ5BZCAXfSbD
taTSaYAvBGsNxzWntM7RX0mwSRLMHxU3DL+R81KQTZzOEGJGEinCEYzyZ8TF
gBEyHTxXkNdkQNwM/QX3ze6uaPB3Iy028bJCWfY5NZLi5bniTeCSqtVef3sg
ldk28vc2EDAH2JGMogTlmkwYeHXVxOuKNZRAMRdRbl2I8rnxNxu7LO4WbgnD
H2hQh4zArg+4nKJSfYGZPWr/vDR62RouMFcnGUrJhO53Yd6ESodiUc3qIEM/
hiTrvpptvPqQkC2mD3VtelH/8IvD40H196CGiyl/mmZ1z7uN5DbzlkojEBuU
KDKULcifZwcMAdD5QDXzA7fDqSHucih136+99QAqG1y+RMeo3mLo+sSEI60+
k1ptVeUjv6NRTp1BSofljrGRjbemSJQezGCA7CdzszVy+ILL6mSIu16kvgp6
B5Jxc1DEFFumA1vMq51TfVqyUrawwRUk9VCWSErkcPVJnILkoBJi5yZ4avbb
oBeg5CE7VRyM4O3b5ajjisngGf+GpoMJdxhwQALbG2z4Jo5lZYpZ4KJEwm6w
70+sggGgLjbjqzWe4m2rDTYcmkJSKrTajSWRZ8BSRQRQpY62yuj6TCIpm8Im
jeZgWuWk85yYf7u84gvnajl5yzk63AGl48G42DYK+fj7shaKx1Igp3rKG/AH
X9jNiny1hGsvK/36+zkho2DtPm/5g/8hplxFOV5amAOzIhkpAgzukVLFmp+A
1rnHlru+NmXQP3fj2KPR0YE3ufF2pfG9XiMpNbajpbnwWvbfrEBrBd5PRDH5
jORa0rADKj52DshcDlimBl4yF1Iff2xnGRvJSDp9N7Hr8FXsDDUxCRxxp3iN
TPugYH9k1wa0JGm7cFYbgELH/ja4kvxed0EDQJTbVWEv5AtCIrGzvfuiocCg
WXOgRlasGoGQQ7jPZJk6RRaWKEfv4Lt6CfUelfc9MQHJNv5p34DbmA6vOy3K
b/BGk0cmLos9ZSjwqoBfab37fJx5AVB5o/0FKbndjjGhOlIPirPO3fmpkB7A
rLbzQ2gdldNf0/DD+VWSbggiv7zJwvxH0oNw/zOHp/ZyjYZSB3hKL9uNNxD7
AQ0QnChO9fDgPXBhGJKWiRBeFlm4kyfUSnDrEWe6e6DTFH5BYM1YvnqYWA0a
zAMwdg+fNtZiUZ6u8ZXfo1fLEiUHRBG3Umkj9qjeELvF+FT1blPiMwvgPmoV
eKZiHwCyNz77xab5QZaFkQRTo22dWmD2oKTSEiGNRDHab1kT5oBViIMycn6c
4x41ld7Iao2gS2xkqzEEz1uC/5WDef/ovC2V93w3HPvSj2k=

`pragma protect end_protected
