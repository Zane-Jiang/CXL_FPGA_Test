// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QKxWFUsE40Ye9287ro4CQn6ChbEzH8ooo1Bpsu8RtFqtgY8/rAfhbkZscrjY
qyKg5xGEkCOeAeFG638RcgM3uUgi+bygfA3r1WuzBVImkLfML5L1sosB+vkm
qAzPerGyWdHD5TfRt1sKL7PP5e1jK7edi0CyVu5IAI/XgvMtgEtdTypsa63W
FXCJNv9/yoXE0zpx4VvCtIUHQUQ3ZXOcotcaBwtpE+uHrj7sQJxpyXKkhzaW
Q4879AiZmhli1d83Kqrm9RthhGzOJQ8Uh8/luK7gOZZ9wvARI5jobTB8eVvr
cZGgncfDNPpbPWIO2PjmJB3JmKM532Uv4GmpO2KdwA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mphiZKzE8AKE+aAWMqsMQZtz37fvc51g+yVM4Sru3OgR+dK8x1PX9wcC/xv5
Uwtmv9L759VYbUK587UAfRA6St2X5qoVsQKQx39Rbh0YTkXEj1Prjvf7Ljpf
Y6SZ0nVOTwuTvRS0vZgKEdO8HjfhMzn8kZ1wFUQu39RSEiUQikgQVl9oVmFr
gzOJ3+BXeeWy5WCTIO/BrYIuW0w/VgSt4OQ5mt/JCPEed6i2IVm90MTLVz/m
3ON/0b1Yt86R8j8cuRlYaqHiVALz2D281QmHJoU04owLpM/ZX1tVYlAvyOw9
g62f84e9VMycpQSAkHOeweAP60j/9N5mVe2LYYjBww==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NNbrwwUiOujQYV/rL29yVdEF9ewcet/QYFwIIyWPV21Ir7o7Y7rfw6GBtGKE
+NPgwocDTgUhqZ4OU/gqiTaIUjsmkveu+KeF/T4sW4mXaRoPxr/E2hoGup37
bUJEDr1KkAjx57ADvGyW7uNgXAOw1dgxURUjrtOu2mt1od7bxLURHSPXG4ug
c+k64dVfh0iYTUN2kBSniTZCkIlQWOAsC1UbD/hUTetW4ekwzTMssBfSk6CE
wlMz2F3VMLlxOF86z2cS8ZWiKZR/45occZ2L+UyiN6WEruClLsGpW/5Uizrn
2H5ct38iw586Pe7pX0XnkADGMIOQiqaUrr7CjiAZ5A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VcBS0moG4ducW7sZfpV69eVMoXLAC8DL4uyMAl4CYpGIEdUEHTbTUszPLxQe
k2rmFIxCg4tkAJJ+LnV60Qb5pchmswdyGYVttDKfkN4Sj0JNeIzAg5gGwGJX
nA7aQZNg7uxNKRGWT+84o7KOY02QYNgZAF/kXNYVikqBQDEN6iQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rBJ4sqK55y7tNOr5tCWAT5M8rkMr377OnyRQWMPRNCO/PqB8StH9ImK4acS/
j/6V8CbT5SEyL2FCeD0Pd3azZKKr0/FeKoMd816gX+AAeoVEnjtz5uyfoyqc
8TaqKpJAqM0cix1aJNusD/RCTcV6/jHHuPlk045cwAvKZwV8+BmqIceinNk6
28eBoCA/qZjc6nsBtqA6pPo+1qMIj5Y1XT14yXazMwqarotUALIygEb5utgD
VsYkQ1U9b26MK5k7xEMr2petIeP538PGogBw52TsAgppdsiSlSKkUZ9r/OK/
H/kLHIwZVTtEZ/uMpEy7bmW5x543UYEnq3PGoVaJfnorDb1VYKSVAcJxJhn7
GJ8AF9+LwKVeEgA9ExibQeKl+00pTCj8VjNESQMqCNFLekzC1aL7zgqR0H3R
GkEO73sc3kZbVJZ23yuAsQN1f4z30luEg0Qe4hp41hT48W0fDZMMdpza+LnE
R4CmGR2s5GYy+zKijdb3/xIiBFZGGkUo


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cQHGd0Rbt2+LNqfttCg25X3DCGpiTmvYar9lX1ZsMQ7q2yzD9NIDV1GT1AqP
6RdmxKgjYS+m/hyfvojtfZSlOamZaMud2ixntIdaUCgUpdfKzNgHpikbjmoW
OQW2/7Rb80F6tWDUP75gjBHGBXvg2RbETGoQYEkWMlLGGG+oso0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nvbhBSUAg0XOSZK6fK9pyc9nTyjNmD/viv8+5y/PFOP2LpD44qa7f0vWd+HC
Km3zlHeWr2yo1woHUSHmY3uSULImXZRhhOkLmj5vbIt+d4LudEPNwzAo9hUl
OW6RvILY+IBo6eXjbXVEke53RGgios2lWLTKtuy/z/NVtAgckZY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46672)
`pragma protect data_block
VTn5xTX60zU+FK0XqLnC67jz80pEp9ERYhf44SbbX+XsStRuPkaGBJtz0ZmB
2ANhJw1+NEHo8opbwNBDYozm414RCYkql69agNvL37JUXN0iwFeP48BBypXh
BvI/Rx+Ataxy1nCSYoO77xHRXnNTaLDYiTJ68IoqWOZcgGyb50dYkYoJr+WE
4fNMv1gAdP5IVbBtdGvnEJD4Bzaz7ffgkvxzEvupCN6ZAksiIZ3oQY+xmOjr
OHwASNw3nAlUp5flNEZTO8b5pnBYGLfFmHY0yfzZ5gMFN83flcbUmGznnKuR
q+1tK9q61H/uzC/Nd2FVewRve/7bWhcCndbm2BOKHW4s52iSHQiKgIh0biBR
aw4yrjKPG1s5gVOeIfSC3sfAnJ1DcybhwO+5ko7ZfBMDC/nWreWUeeiGSH9Q
ddSFPiZiZAQ07lC5po4gHGYzubZkYkGklBQt9NmC+2sy8Gjnk1D6Zy+9dtYI
wJZ11ETAM6AqbAD9avcUwoiRYY9KRmDlp2yXTMrBkZy31V6ALQGYWRU0z2FI
DtCPN9xw99fRFpVHJeveQjjSLjOd0kPAIaFWhk6xLXpC3sOnpVPVoSmxRtE2
fDdTADHHzeiSNOWcJ/JvJUsHxE2fbL9+Yo4skblL8D44tCOzH5N+XCqxrbRl
cBL7xDJtRaKeFD1/GZzXrGri0+8mKKYtM9NhzAMqsQAAu1jhwjXveUIxERW1
st2vtBHqQEEgMB0mbqK1SXZlsYBK3dlXugVkdNQfu2sxFqQxF/YE43iYGP8L
ygw5YYFCRZGKIHaVps7xiE9hC6M80cQWlLlPA9IRDubK7pmlwNX/cdt69yuo
ISzTO/M1qhmnYqHYNfi8g3RATgY8NZlzdlkMLUItHX58OInb9VZYRJvqwPe1
hMu+Xttown2SC7LLHgqJsVtS36VND5SrMdtOCfkDFPZEuHhQxIDX3cXs5aMZ
+SFaPDRxQ9VChczuMHKVrTuP2xxgFzehgdzKDs5HsxkU9lCZmlKWVIEHk9s0
Xa3HgjKBKzsddl0UAYk3x/RcCKbIAOBEFJDG7X5BRqZrKqTSRRr1DVZ+lc/Y
xaniJFZASVEtomrw3vH7bveHglGZzY4ehcqw/PRVKdkEE73ByAtI188ed4zU
DzYY6TBOYqiRxsuux6FMh28Pef8vrx4ykUhQr0fzGY4IOUDkO+2l6eYT0tvX
HvOYeVyxD6LeSOWjYh/wiBqi4S3l2L3A+pAsyEwvFW2h+wNYl1R7A9Yyg0Xw
rsJl6uD6PAbDfDNZppmX5TlLrntko136eyENR5/BPzRl7D/gORnkuHcMMi1L
3F3I/fMUb3AZhtYhL+c4SeAvrvEIsR5zs80YebpSMjzdjV1ZrOs1e2+GZSXM
iCTRBaLvJEy/098FjXY4dwKl9P6fEUZtcn7uSluMD1jyXX5gEwXQZneUIitB
5Vo/JfPJqEkDlTJU0UVD8odg4e/F4sP86d07+gm7RPy2hIfg+/cqwZE3Y13P
K1XjQUXRdWsgY4tzqde6aM5KO0Ud2fadfEudUx/nMsY5Syftf0FRMGrqq3BD
9lvcRXGRGRnR5otkcl1axPcUuAEy9UOEisTlvc3Iorj77LgLiWETQaaLM1Z9
uPFnyMXo4mhrMnY3xOJwkDgale5h0pOV5fyU2KNOZpJfde/emzPLpccr+Zhk
6Z1OU9E6nt+Y6fpHfsWSO3jdZhT9cIPzsuUymzjs4xjMyKbv9aoI2l3k1eGP
JQsGRupa0DMjdWz6yhlmdOPQ4pfpcsTJdBNv8Nt9qr1uXzaC4hl3SDREZOTB
0KS/3iJPNrEpNezlD4ORDpo3h6ysOJs42EMJudDHdSbtywBrPs5mnuq3gQGr
NOvUzig43khCEDKODxSMkb+zgWmFl0Ya8oyZrwJG+NAd7A5AY5fzCHJL6A16
qZbMEV0hrhiA2UuNXPPaH5cmkU5kdxDjyTvONxJDyLAqsasEvxzlWo3FWzcV
FMIm1wb6uP3ucQOzN3WDwW/VoXPAZYLao5o+YMhwdEjynE1YVdN+xGV/c7fn
Dt15QuVejx8sJqJscmt6E9exDAV/2v/4CDO+EWq1ZLJ0o78Co6bbRnPyxPng
RO8BT0oG2bJAgxbQwEClROIXgXTcdVhkNGfGTmfhqVUE4Zi+ZscAG/uyL20l
m30LTsCH3hfXCOoxkEOPV48Xq6Zwl3FOyuJnIR4/PaPUTnJHkQpRg6vyqqgZ
/AXxrjV67s1L089elW0UpVDQX3S69DnWM9Ic0WPdnDq8Q0yB24fwOLTqwJF3
QRYkTf6BjGJYUGB7Y8te/sfSTwJyx7h92jqnbq+fjd9Ec8znukSq/FJb3bqq
kzhfwsXyiDR0ZVWhNqMhXjGSUHVAof94eq2h1dP+Sj/UfXMZShEFu3OdLVhK
wjtq+qDJgSEjcT+S7M3DHz6XOFntr392n91qH4PWXRUAQp9Yd+YLJG6u7FJY
nNSDVK47XsTnHND7qCTgS+MAVRX8UBnF5DAK7KUQjdiTfz6gGKj4nY5+3ONB
axt7B2lhZm86AXMRMaCcl27e6NjGGCyHaEB7OPlPAlWNhnLDzmksKVS8GTh3
5xHM46I+c7eqaCSBU8BFOxUawc2hlm9U7TmQk+yynLv9QV7psTjrS6GWRau8
ElcSaYOaFfzAbN+7R56sJOxW/pQBByAB4IUhQBopQR03zf/tTBNxaVJ3lInN
FFyydkf0zlUE5p//vVTbpN8NbHZS58cLFBOpY9c9BIhgpvviNDKS8Lw71i+B
9c/+Skig17ClmhqZazRNz53AQKnG4rnauKUnPxWXYFjNopmV3wUSy9WFLiKU
PK0ZNuFe79q6MjZFXdUQRU/cSz25Xg3mhvZOtsYs9tODaL9BqnzExRyuNXVa
3TX/2C7OhWUdo0Sq2GwgpWO2mPExD5/ugnmk3szfF9Yd0U2RcAzOR5yY0Rra
ap/2yjZw78S144xdEEHVBuaPrHkUNE9j7YviQmDv1sMMuW4i6ydGjHR38ZYs
JIKJBnxMpO+5JjVv3A/cN0Uc0xULCR8ZyO7Bkl7hGEQlfhJjlKxIJdRoPP8U
XkVvjyMxohovOTTyKPWki8lalNGReCUZbi5fA/bD6Zd6iUYzbWkwiYIYKEIw
ZXI27XNWdhi6m4s2bO/tnsTxTg/iX2zx1gWQ7JYXt07BBp4cXoS0hvXO/I+l
p51sicJlX2tFSlSFp1bNErTHXp1/5Q4SIenb/HcCZVTTgPWaBXcs93rUotfB
XalYB779SwUX0Jea9KUCQ48beHCSHXPuw+bl5iFlq8JU3iegvIjvTPPO/5c9
/W8mZ8F2Og0qd61b8VhjHuiY9IAv56Zcx3TLEaKlodxNCxT61ef0VxiLVb76
P3vEFSqgSGqt4RIiytJNAL6WeN0vts668tAzyhx5lQMvmTamram16tkbFYX3
YAHlrdiCbYFe+7FzNddef0T3R4CrjRv9scbp45fPdcEl4XkfXtW4JGFLI5SY
FaGHSixc1BpurNq+Jzw1lCpftFr6LP1IKqcZtbnpKjeoMHpWFLUGff46puMY
bTl2Sy5F7VGDdNJTUP8JygDIoyc2QlZPu6KwjRxfCg04o16yxDj1ecZ5cjDF
Goe9/gS2jabScq+kueMVvzVxVRDs8ZRqAklkEj8J3J9ReG34f/wmChVGYkFK
mEJ7QtpavavVEduN21bjbZRlfmsOpVjRIODLm/alRMD+KkRhIOOGmTQACkAg
lAkybcLHvUmuICMKJK1r/ao0wudHSth09dmnc6YizDcqrAkYRmQAwBrJA1aA
GDbyxr6Gxj477hoUYdgZ9NnqXjDZ70LehlpLEAQxyD37emWGQaEibxD3XWyM
Gi7/Jn0pPsY2cfihoeBkDH7SStAf4sdlQY5Qx4/kPkJPcHv6Nm1YiNDzTg5R
O8nrhB17hlVJGUGLNuX/Z5nEZtuotbuuPWxZPtyKPyTUFqqz2aDSgA/XZKqR
+foYoervgP5KVoN3tyAHdvBqOFqD0Aj5+A6BM+dw8bvROBPOjj8zWpl4856w
u/GnrLZCjMjPpCUlyOyIRDkRBUutCdQAGfeGv0SPQqHH5JM5V8sC4eNcz4dV
80BxoH+DvVHf1zZnAl5o/8/9UJBXtbVJUx7B63B6FX7K1oRKeQsH9kla/0k1
dh+LXRr9qDxD13LkRwKicXJJxEU9HeRTBDuM/6USzMk/BvCNNNfnTxbHjRiW
uKAiINK7EBIJfsKLwkAQopgRzPcDa7O2hQuWXk5l9gu8R3LsHEFgezpDjLnv
DNgsDb/nfnWK/2dYpHAhNBoZf0vtE4N/spmG9NmAJpsnuAOUeb7aGSpYot2o
zc/58A26/ceTfXHslu3QjLh7QtfZKqAE0w9Bt3KU8YFj30QSSiVAvaRe36U+
R9LNNRhm5WmO5vpPTq/g7mjvFAjt9wWw3vq7+uT9R/yDUtgiBn/1wUDz6jQu
toJTN5aaGMAGDA2OqAvyIvd5NiL2Fiwo8Be53hGbMm+bQPyqVZSQ6yGbqyUt
lZYlOT+87prFUvp3ThLxMpr18mTcvG2lrHJ6NdmCrQFUA77SwEIw7i6ulp9Y
Bga0G+DVQzNjLe2ih6RzMl/9ztse76RMI0/ndJEJTjSl6TChjglxqnDnHsMf
D0ZCPmD9Q7rqQr2f9MEe0pWDnyz2gqomjyq1fm+rhu4DvvY2tJoMFHoSNxip
ARoOFtqXt3c6SN37beZ3yASknDB+hXhfVxLXahpcAS9VnUlS29HV4qiN/QW0
5Hr4zAoWYa3hK7IetTDWU2heSoZ1JDlgDUE9DvxGUBo1jC3L2R4PNhc9rXs3
aUl2FOa61d9DLgsMhH7tORkXBEyWNIsAZFzvlwV1IuknUw9/gXgTyalVf17p
RTQkFp/Ono4ulVf+TLci9l+FUATMbvx5I4iJW7Wde0Aw9WYOiGombtO6UMo4
JMSy66tIVJBRqSLW3A9E+d8E3oKuOC5cHASD7Vg3qzNvgd3lojKoFfIMqmyB
wc1j2h4S2FLUqGkWJcpmUND82oLQJOOTdRJ4842/MaiiJI99Lscf+NnGLM6J
QnUp3cEI2oZvA2UoARuDV/2c8XXpzeNVQhlNnAy/TG2JrmLOg22KRdR98l/z
nk+14+z7hwf2NJL08b1DhgJftssNBr3y6z/ZLf1cHnBrVX16/toPyB0BD87x
mTMQzUh1g7TE1t8x6/nmYXPxgPSvrcCbtOplM/CkuqrMNHVyX+nXAOjxL2Pc
xJRWxhMoiuzhK6mPERJeki7XVeCab4D0IeWdX/yEY6j+joLEXa//JESCfMHN
LsilDRUYHfOX06oZY2jVzZEKwS66+hZFDZ+P7o7x0pkgfhh1MeAjpeyBOEA2
ppr/REaMfMvfW4fpP/30SdNBiNvZhdpmNV3BNbID2ZbApEVJ7MmUhkf7y8uS
59wWwIcEy82w2JFK/cztoZ20pZA1URl+2II/mQUvaveRqU2bzdrjU3TvTGDQ
xbFkN1JbBxhMakjVn5OfnNw+x+CDDt4PMZYztabaFrTiVWONPsmABdMfQrvN
Cm6MqH8UMGjzzSSX8TtUZUt+OoY1FOtt/iEy8kGiSEfFQxLBlfYbjbUUqagh
D5vcpRgwLw1m7+5SL+VY+1hMENuHI00SPLx0ZK/1Z/u+QV9s/1ePogQKEdud
NdZI1FpqAIOHhwD8hRTIbfC4GeUqYXLWJy/f+BOeU9RPNEQmL/tUxoPhPj3V
pRTTYTT/aVqffnD3Fj1Gm/d/+m/vGZvn8vnuQ4XrCjO5IOMXAMPvYPmtowpJ
E9qLrQRox7o4timXap8X4aCNLDno/7j5lewpEJF5CuU5E2k6Np1+d3QtJAGW
l6dN8xpvRArH6hSZVZcSIWYC3lzOweINItkOms67b/4+XgFt1gDE0d4jZpOE
9PsOAX9Z8jCYPHgxUqTZxiuwXCjYPiZ9dM/NyB46YWEi+hPHgiAsVtBEKgdD
TFiEi14qheuGN5PW0rnbpVAkE8up71J4f9m9hyXDkMVpOSL4kjYK3KI5Q2vV
7+4J3uvfBlsNkvZ8+fEKwpk0ErIrXIocpITDHOPFyiNBCZyhp+Vz//weTUgA
Vw24zNjJ19WJXe2gZBVdUSnen84slL2rgUMJo/os+iLRpRXer2ksxNJbgN2U
6aHs6fVS4wKFb1Rcd6BByFtXdNkjRIRs2W8kHRc6wHuJMnR1Wby60cUGWcAt
tpkO6SyY9ItgZuJUKaiHd5NPHuZhoBS8OZrkaTvNtGTq5HP3808lZKhkiHFb
K4z84eDh0nbdyUoTGJFRqFodRiuqftftMIXZdGb7sUcNRkL9xAAFAxwy2q49
ZGdsM8AGk7TPj2DmOFrs5J80fleHisg+ztEWYbnZ3EYv8/RLfWl2dwTy/WVv
82zPqwZWjdhZrkUmFWDYV6BYeFRgIKINaf4ME10YD7t8zs3cuWEAqNMlDWfa
GRtfBFc5bO79phF7cJcHntXhlmAdLTKn8tA2dI9Rzn+EJOvjqeu7KuMae61n
eZk3fUT1X/zXV2lpRyeG4m9WiVl4+ukItd1AATBynO2iTKluOcfm5nLNCxIT
lYioaaRcSp5COgTWe99WYeYgNMhWJ87YEjp2f+jsDRspP642ErAM43o1YUCe
YxwgbWsMxRj0ytiiAof+L1rgavD47GZ9c+qfr1kK6qt1uBKDCxT9mPZgRyOX
XZWYjwVZc6DwvrV0PVVjCYJcWuBDB9ea+7Pa68IpUgv7fSzx1NzvmNXfulkc
b0pdvh1EqwzT6F8WtvflTHIAqPbStq0OELylBCENKpYN1tkwH+H7HqicgSyC
R3QB8qOwtBr5zLvLMlyB0ufwnlAHic4lgx2wmAqFr0F7K7rSlhUfptmK6wme
xCxaY3PT9M7IH7mGQgznAD+xEZp0h62B/zTASVDxueFqszsxxuUNq3ZW+zeq
uVitkPecX0PBLC3gdof8rHOprXtkgAsyWercMP5tq5slZygANaJXwTdwGm5i
IucA9tRnuiDAUg2rc3gBymovab/UB1zbcxN/O82VAUg33WrTywpJNw5yt91B
vnxmruJmhAFcC4MCRCgaVrS2U9pxB1aUPTLOEHnscZP6oYRM4mQ3rfRJARGx
zTV6q1nUw3GYI2oZ2u12JA+ib9rD7ZeV68QHhcY10dLGeZbkbIUs6fo+k8jl
KjwJb1GtpJds+rI9bAakgzeP2keJ3HFMBO5GquE28wipRGV5cMQWUGc72nsP
pv5oIh2xpLLz25PPkSI6HkU/ITRXMyMdZQV+ZPulsr5ctMMummNChgUVezDb
Nm9n83u7XS4Agm5PEqZDIedovLW96iVz1cE3Lx1+1B/k8osE1UtpNn4YQ2NE
KR1D38Ax7nwjz0RSXMAGX1Y5P1UvZKkU4hvV+dgHZfz7HRk7mc4IeEe72cDb
eC9iFGpL6HT/Y8cnHyb1cQnPZKsX2IP4wIoPL4TabfLNLnpyPgvvPq1q48sH
qfK1YK/EWKIKsPG4hN2mbJmGBKZAijMrua9WnjCVJXrTZiXZacLzg1qIZsmi
Uqdp6Uc5xaR5x2a2VYA1Dw+4jqh8MXUm6xL62jyzms5fn7KDrQSEzNfVVLGH
L//jTYk8ybwAbtlVQ6E9Yn3/lZtGN1hiYHMzFL2ni0a7lHfAJEfkqCo0cLy9
Evmb6Mnpmu5XFvbDU2nGPAswKfyVdixmjMZ4593pOne6awxuJ6Dlsa635cB1
6HKrtduX0IS8zXpa7OgFGSi+BoFgJWzA3d4eGGWfou1jchkV2Wch8lYxxuRa
vhV1bxH4X/EVplgQJFzlmrMQUrsI71lOF8vOzBsIi0XKXc99iGDoAQQwyysA
YfsI+EijhqzimLNO8sPv+WaRSE/wHtoAqPCxxjvJ+KK2YmZdkJ+HZn8CJd8S
H5N2iP6/1UdWE4w0rQFP+w7/H9uJ07q7p0ho7LIZhG+MlKzZJU37sPf771ie
+eKa3g0BLEz7Vwxzx6Tcp+EdvAPFbVD2bWQSfWo771UqhJ182uxt+1FcQHcY
JTFlqGqLP9yYZULC7WKA9QVKeEnZiN0pb0tRhvEbXxvDp9djgC6KM1B9oJ+A
GCJbv+fnGayz5Nc3Pt3xuSi3PW16QNzpYTO4ywXDKA/+jBHN3Ln8osQ5wum7
WW6lxjaenIsubl/jaG1o8/yYd4mr3Nb7ucwzvhm3NOr+UK0Xr3OXiKypeVvU
Qv8UkDvhN9hEof+VqwS9eTVjG+93iUx61nTCYJ703wt0v0Z90Sgc/XtCDa46
HQXO9u2Ktq0B3qSzKETUUUPLwICA3IM+86Hyp+3dPPD8yKyw6G7q7kzpUY5F
uccw7+5GFGtvrX7eApOTs9pgf2evkUV8ol8udFdAf5QKHlV6kDvSd17FPFUy
LQprHmaQMV2qRWo2hrPDqMH3fKY6onCOLnmV+5WyBDkDHka/ol9vNHtTwNnK
+tXJtijXl1rMx60A7hRI6d7FjsfoDzViEsOz0U60ZSeVMqqmr5dedMC5lDBS
R9tPd9gasslNLYbWvdDcuvGdvWTnpAwcq+WFK5wIjHCS9ZzDdzlnKvbPPmKP
krqaLgYwuIodN0iH7bhEf6IOLsXI3cOcMqaBtKPWN476ujSku+s2JOyAug2o
DNhcL2w6tdRHkc1cIZadlm2LZw7AY45jmLacxOMj3EccFe9iYcC0nJ5t1YQB
aFgcsluJAfRBtu+4xLNbgHrS6el28fY3nJXbVqhNtNw/rYksNHD216F03dOz
+djB+jXPjTYI6EBSiT4tO445K9aK4lAvCtVE0Ns86XjUSPrsSNpJVwB9Vuku
0sqXONhFoTX4krcLtdXO/Z44s5eBzNRHUWgFGafOOJT1yFUj0YowArHoBfDz
o+mBwOcpJiIuorp5fe4rxRjvGDlurbUsKZtc7GxQUvx5dPjMGHrnMFzua3+T
1NLIWKmpLY1knoF23U7SdN79mtVFnYN3LTDye1N8nkV6oz4Opk7orWoixQiP
1shifOktbOGcp3O9h5WOCFlZWbV71YRXpMFgo5q69L3zglBy1WTMcPa56ECV
jv3yWWigkmtIzlmgsCIza1srZmIUSZ03R5iw8jveKJzGryvhyTJQjO6i2bvF
iVERxiFLvGCQBbu9jSaUoKl0d4itvllm6p+GVNJ0HeTOh1QoOlIy9oVnmc74
TpIG3pHuqZX8jOTWkmBKb7AqEcDgNHpCslZFixPvKvJ0/F1xV/1zdVp8bo75
jDKVH5RJOggJMEBnzGBOSzlj2pElZu4UqJ+z4n7qFPywcGOoRVyrGKmvwdt3
L0bgVGszDFFCalaxQh4xxeP5fqIH+zEj3TMXpGGvydnTN1EGcE96aZgQtL0Z
+boAymKP5vAbKbZyqVlwnza/t07Vc2Hf0PDXaq6rdwtlDsBitHKVCjVHUz5M
8e8FeigUBgW9BtRRKQBQc9zrRZT1R9AT5y3pY4qHhBOPI6stM4vxK57q0jJK
jbbh193ptfo7FbFhU8eDBNKDG7MGeljNARnlFJHTJGHrNREat4sevWU3RsDT
eO1bQiUbW6sgwdKlor4qXpT1/l+SM99wVXPUMRqo+XK6p3PoaSkmTnigpRBj
lb67wGRkZJvYU5sv1KoFLf4fKw/Hm2RD9xNfSheatfypidu7Sbx7KqFxkqbW
39XcwzdqpZevb9VkDXHlKtO1Vz7l0eNcocT4zKAaee2jW4kcJU5UX5ktoW02
ZyGhuG6QQzfWKWZyKg/aBPfUdxOcDxSvFExi/666WGS2xshdIxxa3Nh8EWNY
rleqFjnildbPsWkbRew4F75LODTNW9gM3109Mg93byJcP/p9yzWcmOIm72sB
RtLErdEQbfsDlsLAugJdQiAGbzUVoUPPcsdzXp+h+AiQ1l6dyxbB4R1CXeHD
IfuwSZIGWjbWi5ieuogxz/wxPJWiveExt7smBSsnTSduQql6SZEx1FlWsJOd
JIqG9MPq/LgK/k1lalH5xwSpd/Cpr7pYFJ+1Ol5QFcB39RewC+e7yt0cX1FU
Yp0SX1WuolPcJrIQMMzjG5dV+FCTC9FsqqdKvNswMs5900s/6IDQnH0stwAg
f9zU/JhpL/Ww71XBFAT6nsHCBWYh+5l6FIw8GOvdbD9ViWcCJap7JCAshS4f
ulRr41IB6I6/75sE7kbN4AsBb+QgiQHwy/B3xs1s6zA7tacBWzDCIpQj9VHI
EdecTT23riAdwDJ3L3ILej3tylvoBuffnXWwAq6sn/8HboINKRoiEL14/F1T
Pb0mwHVxwcmu5EAk2+ooNKTuw5orKM68eH34k19V0o1oUXdhzLrHZRJ2s56Q
aR88fLaBtYT2cN8/ub1Qqnp2eKEfSjEiKaCVZau5BfWC/WpLDbgToh2JD1pM
AbwiPUbhbLyCLfd6sDL9OEMmJItoYGjbTzQG3ZMdBsdQhGps1GXcTTFUwmaH
JsusFWaOQ7DpHV+8+KnqP9FHNLOIpIzSlP1r3RFpqfbMPwPdKcD6c09u0waI
1HSg/WmZSlXwT/XdHA91rEMMs5zqolaoW6E5dQQ37CbqAyuVIz79eCnkvTEB
16BnNER3lIYjpeZtxF3eZUkSeGgodoxD/Flkq1v5UkEef0tK0UNDvvj4XYZp
qzPvmIEIChYk//QlwWPQkbj7tLjkfGWZgCJ1ujx4kBwJf+MkvPyPmLOLHTlM
8oj2v7nRxH9+kc+lR7CfPBw4QJN4UH1tIKUWXR9w2uY53SkaLcEk293s/NJO
pUVddUh0L3Vsqpy9o4ylb4gRqoF9fy0Dj4Hm4QGDpjHj0AGF/FEYV/MjUJSE
5tb6FH5eXMhSTcaT81WQiCmVc/tFlu5OaIao2xZ4RGmTPjl6uZOhq5foruvl
JVXifjKPZv3AjCMRZF6FPkYv/E5+YOhDkb22/rPEnc1AnL9CnN+DXpVDhp9+
eOAx8CL0becntYlvDYRvdeczBVjAJiLhe7nxis+x1c3Zd6UWR/asvWMEnnCS
DG0woB7EREtH7uQMYU9Pdg3Ingm/2uTupHGTeM4VzRAya2lCMW/muhX9MD/k
Tme53jEm7ATZ/LbF5kCCTA7jhBeCNMpbXurkzapg6Buucxf5fwGlFF0AMvf2
FKyZjiPi/J1M/EWx5hzs8o6kHsL6rgbjOCH7uNw9UMhBOeleIsUUxCFiCxhG
+J3Ynw/TSx9JL5tDLDZBB1DR35JT/J8AIgnwgF/GNvYXn/5w+LcGo3Nnc1vQ
mtSSTtNIst/h4o57Llb+Dbu6PC9mEJn2zi/RxdaXdIR/Wax3gPfcseLyMtVv
9XtDJun/x6n+kACYyAPEt+f0/25D4zOFmY/xxYOinpT17pC3hIRmjkm2nrjQ
0gTkOZtn1AY/2U08msMDRJ/PdHrzQ5tSc4pyO0LAg/MF6u+c/wheC6yym8hS
CrCGOV3HO/xT9dxd/vd7ogG7h7VAxMfsfvon/y0dGvOton7e73/NY913alpF
Hno6H74GkTqs8Mx/P7BnaArMljRwnmglfGh1XwT0tKW7nln4UxVn2WFwinhu
nMphtteyUfruOMHHK/wBFQL9TVl9ldWcmjQ3Ku4TvojR9Zi9mEj/UDoZYpQe
7yfHt8TPVb0qn9R/i82fUTy06raHVAu+pALEUY5xjxuCRPYrGjxIsY2RVj5b
1JbSjyRg3IJUtiO5oOks/c87I5lHunDfUD5p2+KJREAs3XjOXdVZ/+ErhgZ3
Zzwu5K+GAgRn8qMKhj77oBbNG23ZJ/Qz2xwIIF2F0gwvqs1Vf4nAA3d4/S4p
fuxZMjTuCnvJJbQ0vEpjX4c7tRNvwmXM5FY6T64qEtxAPmDQOUSnGs/yrIIQ
qlmTUUhXE+34tWLNmWfwyKEJpk6N4E3U+rIorrUJ6SU0J/jff8FT1Lq73Jv/
odcFjYW8hbfAvB+UFwLY6f9sNaSx9Pr124LPqzhNVtQLYBzZ9NUkjAryqhne
NwinGxRr3zAVCTHDbgCsRJ7I6DgjjrePxjTg4D09ETTMHXXUkrxpmu0cGP8T
T0nRWF2hNgUtl5YUoDMkT3cppajI2SZZU07w4uU2/fIqLUg/gShn5KPYs9Oq
PEOi30R8kw8x0J5gvEs+zj5bNZ9boA4e68QODTCb8mU5xh5clR/SV2iEW8p6
sHIkzrdJaXAMqxK7pPpVolZ8Mx2P2xIGHjMYQ2qkW1k+JsQLklZ8SvOAuU7P
rwMOUn72jVXKOSsOSYQiJUxiTPpeNsB866pZHMdb1ncPQMNyd0k1Ai/YCZjq
UQPUGAdkuUrUpIbAqe7bHNAAg5QT5QK3w6r0RfEn/358AQx6JwUgJ9iWG9Sd
NjGUxEwCc/yGcLIaQRo0L6XD6qtseiGMKKF/btYKIzUgvppsTa7P+bG897y3
XsTfWeKpcePD0Trkx5C2xcgHGORA471mXWQ6tfM3iQoFKJ1QirwXbuEANBEf
LvvxhQc3/d30ljgF3tl9ZCgKjuKhEIWd7axQ9Xr1XfPKOGcnOL3ojCD2ltKH
hr6vkZebtpLra92bSvr9WWqaKD+wCLyYwqQp6oc4bNmQtKdYi+ktBiEGrCS/
3+xsudWd7PgQeHqglzJ743+4XLMn/gBwntwDnvmlTnX1VoGuahgvnMUGFnqH
fAZsCNaUDmUXl2DBeAWofNjP7uPut6xfEj0ye5doN5557fhICFyC2xaattQe
FF20PSIKda/ESRgcJ+oojbbEHrjg8G4eT8ArKKmSsvHEh9VSM2GsGTjH7vsr
1ALL7C8IEXHZuEDuTIrmbSINyoG2ix5FTZ+xkj2cPiSzg3Ptxo5mUWnohNfY
o2uAb2G1HcsI8PJCypDEC7o+LdJrr+gXUtik57e+qDdy008sD6gGpyDIk4+a
Q2de0X9x1RTMyZ/yg+dequ0eNf3k+S3DBfvD8Mw/jSXWYddIQKeyW7yh0knh
LtklptEp7k386NBtQTlIxgeqAGStF2n/BKe4f8btIIVVl4B1mLd5ojUvPHdE
Ca5y/iB6YcWdB3keCPj4Scy3lbw8Xl4PcXwW8cASposCvhv/jtOtt3WZDdw5
ToKEaH+ib2W4c73r3Vb+5fjsQZ7VUbuMpASfMxzTpH4GF06DGJUo5KTVf4L4
pgb9PiNEEDjKVQyACVViDVHuMlq//ksiGNugpN3A0fSO+0MLzdxTOhX12vrq
MuSE9Ud9COLAhzOPochu9CQCeDcRIFby5pS77cVrS4iOV7HazkOuBFafySou
uqYGI94fWMGaIDFpuOxCC0ey/rIjf9P7MV5zb7CznoaiCSDLq0MDF4wj7q9X
Ob3cSw561DzFzThHslhhs7ELN21HB6TNUXcNVucrqwVbxayckLYLMKx7nCCT
PyYwYuArzJ4Qxk9byYPsr0R8yO/nk7HaldZ1APE1yBMsYKYDgwamffv8VULH
Vh54yyLPDbvsqmTNuNSJLrY4DftMWDwHRYT3Rrl3PgWY4W/E4GDIWePXXHR8
ls1C8dJLiOED5oLK+Fcgi1mS9beVDJCJzLajxHCuql8SHMkW8dr1lGAqj1Eh
FbivwAB6mRZ/ONXoasjP2wI5OwEn+OEYnSgpJGz++zbmVThHR9bAbDxJJuzs
u+6xzMSlz40BwmC32XHlKyiYNNZF1IE1JiGYcAOClzgh+rM1aUgVOLNR3Miu
Tht/YGlFIhsXzZEYBQ/o3euFmi9hA3sq62HWwAJVVQDDrrtBo3C7L+Yhoa5t
fy10D2toFlUL9diGUi4AUW0qQgQHn2t3Ki1RfPo5yf6uLaoc5W3RwBX7WnGj
WNk0ZRN1tq9kWwa4/10+bKUG5uxad/BNBqHgsqbNDkL5Pd2bPvc0yh5YQQUM
mCM93XzzCqJWRDvkh8wSHFIRjAxomfyShhN+vN9TUAUZ1+6ckrl0qIct+CiK
fUpl7l4f1ehuhmuwvaHH0m4/ntVy0tIo83Kyuq4Dpsr2NMSoj6g0uShPc/YL
DkDfVW4eHj23X1gS3imDiIm8+At8Kp0VjCyiEZe4z/AVhlBxNLjvaGBF/GQ3
pM4eUuZcMhpW7vNcNmvEkQTcUS/60OVCZ+IZpKqlP5AoLtScm68Sj46SCGYo
mVpVaLGMlaRUZ72wGtKEPX3j91qBYknyNJw+F1VrMmR1PYoNkWmCus9LeVEA
i/nWE+TF2DQKnDktyHnJ4HUCDNAsEFz+XECJFkB8cA46fZylSHLjUbwGXC+i
z8+wlWgpOFis8SHNF6jl4bnESNJmemLeFXP7WqfyKi4H6vhRGlJJYFqywSOM
U7jqaKe7sEFGxe7EZGpFKoUI8XI4tYVKMiEAeTCaJ3ziWBkcKAsWZ1jdVAf6
J2uXRwvOfrmtiKML4mqrnZ4AzeyiBzCOvyclYJVXYbvq0KyciyTd3m5zm0lE
tJn98FitjNYX22Y8SHx68kJu/KGd8ayKxqadIPA7JLxKUz4tglOA7G8OgXKF
3st1S0FzmGpF6z23kZvNf7aVGTVjk8d27/jmfS5s0rpP3WwWaq9uBumZ7s0j
loN+UUI5n1N3MLAB/5u+aQQSij0ZbB+rMXjeoT90zAX4gh+YR8eoQ/4dwq0J
1WRpK6+4CGlpVe2kfXRZhq/TzDgSV2wQeMIV/H59grBWHcaSCb5r+CH++a/+
kWMYisSFOq+1ZFv+3m/JQLlWaPSD+atGTjhDr2lBS8VsEoz89KXXaUngDVHP
wO6DYgp8oAytkAke7lwi5M0sxpoRpvSMw6uKidUxlcelCJTjPi2t6uIeqF/2
OunRC6zP+38mSsRptmksEyMs+N47easFT5ZXnh0zUpoEPX/DbMdBPzj8EYWa
Lo5ogyuvxmUJehdOydnOmAur5DoXKR26JuS6jh0GGYaZbJ/kEOnVmrSDsAWc
zLK19inawEqb60KOAFWxtwM+YlRTIJu48KC7YygNdVAOh+QwC6V7HA+tdIFt
2DeKoz1YeXTev+gGMX04dhOzshSEMgw10lfQ9ElRGhQf3tqdu622dSFwN0vS
b8UoY00Gfd+bqYJ4HCpGPLBNEeqI9u6YDF9yIxcBR8tvRFO5bQ4haNpb9k4C
8yT2MCs3qxQqkmCpuR0jCs0PP2INxpAKfTeSlPW80MRTC+E8yEsj7A5Iy617
Kt7k8Fg9LSHa8NOezK8K24Jzr0AHfBtItINfV1xg7cv7hOHytOcmvtYCXxyN
mBjiyd6C3YwSExXcVPG4KEEhpD+C6y4LnGo1NwlbBYR9Ae7BhS4si88cFpQ0
vKfAsb289s1IPuvxEUuI/wG7cW9L15SLkyCG5Vk+HAKplTo7rR5uJSktCkKB
vBTf2MDAXxHtoExYRDMUnvap1SaW0dA9hqog0UuTvUds9pL/+JV9wQ3+QWap
qC2RdBQpOy+Yd5Ea3yz1cZiil8fJqyy63f28lCQIhG95onDmS4XfKNtzEttq
LnT0UBjU+TTJ1QJjaIB8KNvFJY0LK0SyWzt5HnHA9JArD+d5UjgrHXKvr2LJ
WIpAcB7VcT1JzH2H+9V9NQBM7IkZobOny2g/qGbBxPuRH/FmtppZmGQgdkFh
ZeUAXEpMaclqrgs3yctWkOFhDv6L1ZIKgrGdX+rndpXLv6Omq4rKytj/xJfi
LkmLX9MZTJK65hsX1FVsuvnMbfjmt6BcmVCOOF7Qs8mejY3jgnpRSkysMYDE
wriNqqvYp4qv4XBQpo54/Zz2LW9nz3zBmCRZ3MXdPX0RP9LY4TqTfYk3mFjf
Th8A6K9InTQDEVQcVPD6Zi+DendbiTlRivoSlMSNRPocoO0ISEb5ZkY4LbER
qdX7ZVfUQM1C9vxOIO1op6AtN66O9pK8hFrvr9+s3h/xrE22EM432TyLDRTC
C3wm/5a+PFTw1D4FU/JWRdznmp0fN57kdvZ0FNEBUCyRCOSyavsW37C2V4MT
uHytjXvyNjdEGTE2c+6bRp4aca4ITgS4SpkSmQbJO1dHosN+K+YGT+ka/E1S
5jvw57yIkYMH5rN5P22IR84wOrEfjohkeP182lp2h6UOCxmlbmkFUy4YAY11
WUd4vhciXOqe6LF09MYWJ0GxT03rUkczrn9n19sf0E6XJ7MwIc99KKAzGQXD
+pMGr06eh9XfLAZS3EylKSPi6oa/zTxOX0PnuapXvZXDCAnTZI/EvOV3kAS3
TeRPgipSwC0yJcCipaVXWyBUn5Uh8ULYsZvvWhiMqTGsZJXF2WWFrEJSXCII
Q1gtf95eVtfBBM5guXCWBRYlKIdWOBHCnX5VKjWSJZt3ugy4GfoM7FBW8arN
yKTAnjFHZ+svfH7NE8xzR+GiXbcwlvfhg67KMuWfslDPmbhpIRt0viK7BtFQ
SvBj7rBM/+e6BC/t5KDhbg7DdoMXvXY8BbZdg9aZmEbdAJyYJVR4qkET9/u6
rmJ+7haZxmXJvS7ZljTS4hoWMhLsn1evsi8I4yyDpMdQoB69y4L3swjCZwh4
D+k2fkwDANgpUHcsY8F9GqcKwnqszzn8U2/4+nhst1wgGQw9/4sl2lxdgTWn
bNLYDnrDANqKS37scI/cU+w58GJr6keOF09QxgcccDNWbete1O4ojtuC/hSU
0CZZfmfBwEmjVfHzcHkAaCyvASKiMMCcdPQb9N50zk/yMIGwL2W+ohi2tSRh
asSVB/XtUVH2pac1XO6saL5Ubg5d2FIifE1/CZlZaGyU1wporBz1Tvq+noC7
91xRMzEFU0rmhHF5TuA++GK5N9uC5yhLkCS9UgPWkcKmpBVBGybLf7/3jSoW
MJtAxH7NSaHgXpQndjYi23fzRKqSWotGKpmz0HYzIQBNL2W1Kgw5jOc60H2n
dM3CoIR4+gSmt9hTS38emMEX18ufDyYNWwxAtX+nA4Fd7z4PluT8ViNeAKmi
pdiw2EFRGt/6e7SJ3ZVVXOpJlgiIXiRN5IEDmv8caX20XyxMDnvwB8V+Qqts
koOVCWwOckCK8jg1/hhG8QIwJhpC4cn0I3hBIaQnx/GkOHIrG6pb7dopNSkz
Ph3AwdT5AulIqNZXvtMAhvWd6snYHdcOu0X0SbiJn2MA4RBVA8G1j9oNtvEK
W2AdMSLf6wOx4xe0DA4I/XtpfNMFWDdfRImRoxnLuNWC3tDhkVposL/FC/rM
Wgxbs+Z43QXuGjY5IrWPL8sZyoAEHP8KplBcdrYerevRQ+/fl6UAn1UeVskh
wti4sXmZl3+RMjM27R7skEciQ5yWh8Ph3ZyX2bzv4p/XBGVk9RiISpiRgymu
pK07NBIFETTjSzpXRd1yrhUDN7vaSdfpoLsq68jD44oSHh37NdymyefpmsIf
hJJH6Orll6iqH+gSofTISDn/JlHU+kt79nlaKz3oXgppVNGyO9BJnTrThIKf
0g3KKJbXyEhKFT9CgMyHXnJFkvkhcclJJm9akgfqImGZu1FH/A71lAiKrbjo
tDeK+xodUpOMpUTmN2cSbySkBzNfBtw9gG2rlKjusQ6d1xzXZeZlw6xanj/Y
7v5Vpg+Kd9ByeqtYhzUVRqSkkmaoqfnmoet6vvzvDoWc8yTv8Qki1Kd8ckw4
QLeCq1OTW8I+ytkCMrftwSHRaJQ9y3gJL3WwkYxN8fwx/kyyBay/w83qT198
L6ej4Y/ZZAZ9mylhIhnYL63OE8iuakc0xb6gCrVqrT0AucAxGvwvTpksdKfZ
iQ1tI6OWibqoCNB1494Coj+GLMC5khhbt73BUEWd6SYlao4G3UhIR3GrHYVW
rwu+V1vr3xXARgBDNJLy5K1GMUXCpSPOZzkl0BkJx2Vm1Mpl906FwZZO7pnp
QkfRzAJabWhYHwsrv1b5gXkA/SiMxES/QppTT9pLRWfAmM2DzyNHo7Gslo43
atGJVZntA3l789F9DYh4pi4nipRh1bU+qRxMGMsvbWmcPujLtJodfPmU12bs
qScrt/BjGj4PWu7ei4qi7AZDSbbMteojWs2yQiNgPrkyHiJ3qSrf2/g8RoiN
pBmKLm8v1MQLHMhoqlbHL8BmnE/xfUbfa0lTUComzdnMmmfSdEKqhO3aoBk3
+UGgcth9YGMwuc8c8q7r1iQDffQ9g18nS5D5wf8Ho301iWST8WpzyQMGHpqE
dXQLo9I6N4/6A9V6Tlx1W+J8CKBR55aGTiCUyjjAZubyRLwMGbQJ/I53eFkl
bqaJyBXJEPfC02Jh1oqdCCBDxU3/vHymxFh3G4U8CBfEHZn8rj0oiqts3el9
l1DJdxKJ5VZ6kjoGQfbg6Ea23ZIUOyXrttTZTeOVOTAq3o62ecHdxNi5a4Jb
fU9um/XKUDx8fZLws5z3INn4CaX0SOhsJj7yjgnRqDUDgrd4gp0LkLOp678k
ruRT+s/5XOamA2+XZkmb5Avbkc3QnyzdlF14F0JHyLKR5X+abZNyX9zbldDO
+AxEPHLZIUsxyItE5/NoZdZYXQdSnZGozmJe55ghMD0VKE9rX0dEnTaMTyI7
yXaB4xsDHpVPlNedG/qTmmAcSQgRxEIRHgtCI4jSG2oekKta5+3+msEPriJW
k5IrxQb2fYhmvWDTR7uqlGd0Nn6sL/IV37KENsL29q0i66XuMxYPNVG/wO7R
NzMWMlHlEi56PmFHS1Jj8eJbQnHe6fShbyPw/Q0leOsQq1z5OphdPO4cbxEF
w15v/BPSGfub0E1c23YvVVE2hySm+OoMkMbpzoC4/ZeFUoOZ6RnGs22pl+FX
CzEVLxJ0Fsxbv0KhgPmeBGke4aD2cnwo7NNK4HxQVcNPR0Z9KuYeO51OhBHR
AV58mHvBmy3ltALQWuwqV8oDIbNbS8ZgrvvyWc+QELMhN2cxHq06s+GZmNSv
P9fL8/NE5r2Izqacly8cim5O2tSZ4cumZAj54ouHSX3a1kNzJGmJo8OXRpFh
sm/bjrFUGdzs5sDgCyKlLde3xNOF/ZYQISjUnAzAnSng9L46x+ljpxUp/r3+
LyNHVvp+DmPpgjmynOayKODmP8wei7RrPHh1ePcp21fudADZToW+Z8EVCHAB
PL0J1LD+kYFKU8YyaaG03t/Yik0eIv3p4bhmonRwJbJjtrH4T0EBotUQ8+xS
RG/vjlSaX2D5DOsdf0mxeyXjEw4quRpqZVFTW3QBQCVpBYSk21IlnL1333yr
iZXRdjQTdxpV5DcPdPp00wknpUiJ7Zom1uEFQy9Y2U7fkhnizyA3Y/WkWXAS
4ZTYqLqv716UoDr9TMh2cQJIF9XWQfoeYBUu3z5fzEp5cuOnfntXxZFGU9Y+
dhx4TizcGG3twyiYVUXIsJPfWKKWhe5O7Gn8uLCqwUHmiK8QC1FUOgt1Xm5j
erWm/VDDNpMm0ROlSZEtoDm3rC4liCz4wlGUmzp+i/8JGkVQ4CePUySSc2L7
0Go+4ybp9LjTSOSiSVSilzQ+4K1K7y8/MPyAzwij6SNEMT2+QYUk2B7w7VyY
rtCN0LA1j5cxeZW/TsflSl6AitkLt6yaVUwwP139v9lC4M8iwbxwI7CObTfz
Rl8qqY4Rfd7cRxON/ynQqmJNroPslsI/VztRL2UHlQeisksQ6acbIrq0MaUW
xwmTjvgH5KPNTgSOhMroph+Dtp9A4EABCwKes8Oid+nQNwxFd/lhoki61KiE
SSRbCuBVW+KGVKvUYnJ4AIKx2zaFUoeDmF5dwlLLjKN5yKVx00zOXNBnZKZI
8PoR8iQrnZBg+H1yiOy43g4Yv348nwoGnI8SkUgf8kvHRKjSaBIVlA7PtHmW
nVquYEDLUsW1+PvAfcOiuSkRiRo0Ez/kydLBnxDBkeVKcZDGqffKHkyQugKV
rscvwwizuj3ImdqCXsMzUOJDmqRg+Y5aBsjxpGR1BmqDwZAp1SY1eg37Kezt
hZEYD10uS9yT5RKJnnbwpKCYkhwXyOIUw2PEpEit73YDyIK5KU1Df5Zuvmp0
sYg0FXLtfhgE7viiH/XdHMbeDOSVAXh5O4iIwq01zdtqLfV8hUMAAE/Lisad
DkUZrlySNE6bEVs4pDmCd4DSvaDUvsBds2N+SQgbcuRpkpc5J5ty5yQwGY/U
vii7Jpy009AIyEoqEkZWGi4HXOkdPsxntF9YT+We/Vd9GYbEPhKmXvDQH0CF
O8u+nwxuPCK3NX4dnkYs5us5NgdR1DyvUMtoOuKhKGsFr8NXUG2zsjgwP2Z9
dbm0jV3qd8YNB8MO6YINWL6Ox3ASb+98EHKdoPP9wE3un44InZDqCHS0LJmI
EDuJq6T2ViKXM3ehdUr5KwJfb5+YT3IzrY/FC0HU27+mepkQ7Leu4B6lUnDk
9e7veKXmJ9Da6eDKp6V12X/CTk2iYJ5Ke/saSuWTseA4LbfEVxrCmWVDLG9u
iQERC5xI1760TMDn9U61fpTNhkKp+tXHUwwIHnZHCHV/LmYUgBFzQ3jGLNhf
ZdaUn9t86FP/Y+TZFgd5kLsWCOmXXL0deoDJv1V+Rz41dDtbIa+tzo4TyxLS
Z+vdErfwCaYk8o0PqaLxTEDyOdAxrbxavmqsCYwyKJi7H9RpmiXeTM60oMp8
iKxQp38uNa1xOokGUvEDHJCd4kilGQQKgMErgGu6oAbLr531Zhy7NkOOzZ2F
hHNT7zSt+tQHos1frYy1/zSXQn6pfI1C9Pocs8oeELSuTHBfx3TuFeegs+ju
1cRiyYZtjtXkFzubRq5JMZUIXfSpEfLBhA33YnzhyxpZrB/zwRgz+HydB0PC
WD50IOKRVSWcTJOmtEDB93ZANpW9LbhqxAAgwLiUyjmDE8xcITbiwydW5u5c
Aq7W5a8v6Q/MUfPoT3Bf828pOkE+TwKQXpAKmpHK7TZxfh8SFN1qQ3quyzll
xKAK13Y+eTsPld+VXozZeqCTNJ/7Nc2LW+Ea5M16uG8iEzsYq5uMnnHI+Cjo
LDxnZznxClleiyOLBX/juFOGVEga4GhvB9BzJXXGP8UL0pE7e5s4lOztI3eE
cXICFRQnaCfyyhebr12k4XpUqgxYiInaooC1HFQN7D8kUUPtD/p8BxZO28OU
FckxzoC2k4LqVObw/tqgJ8MC1CzqSmDx1PG8Onh6qE9Mt8ka64lTS2kO6m7Q
C3BBkG25AD4tf64OBYZ31LrZztc4FdQmOoo0HGgyeJmR/Z+YLfxSPnnddCcP
sFDLvSvjbpCa3Gn8BLnKRkLUZXDpXPs1ppKSubJIIi15p3oFpyfVMXba3Z61
gj6wc6ty6BMbzf6hPEcxzLHgucke88rKutL8cwYK9EHPocMNyXoIL5OlBWwV
2QdbX8ASoJSRc8Zr27wV38b3IQayvJ9kLgz21yuBk2QOAUHPl7jVDuqobMNI
DE0g9nMhSHAOlsNsnVdum3bA1HcjSB1eYD5jcwbOg+3YSLnUU8d4COSIaX9L
3L7jfTU9A8mVJteOI68JVPLC6zfZrYOwW4pBnCzShziyWgx+ZLEItmHpBmji
3jusesd5Ch/zD4oJ1AF6QIl+xym0O5FlZaOkv1VRadVKtCFSmVpgdRKZwfdK
CWul+iRFHNO5sjvQFqZVlgigNYbmtnIUAndAKoBT/FzccKkTzHymDXKtFrCN
PYk13zlZZjBG6B7BB2yjyLZWhQXpZkW1MvS5eixyoIfv3dysqJWLCUN4VEAZ
x20WuqiLegxGBEkc4qBQFa2BEBnXLcNj4GSF77Q+djXH/GcBnJ4HQR3WkIiP
y6VeuhiTvUc8uyY3F8S8SHAkwfTpkyK9kNP1/+f71QJB99nuzchVIImhIYor
PL9G6XgeHtT7VStAHrJIYlpOfW3sOhB0Z6jp3/znOh02ra86u48GaRR3C93p
kDyjwEfZKLgXesvfh95/KM7r8PszRytotnFibSRCcwuHnv6BA9Tp2TBuQn95
QFrQn7H8KW/p6s1WvBvZnOTf0pads1PrA8fX23vF3MZf8kdeQ8qzulVVsWRV
AvggzuB1ptF1NyHELLJ43bT7Njheo21Eal2xZv6EfOuI2Wh1+QUNA/1Q24ly
AdqZ52ouitCZFUbzYf1J/jPfokcIvRbYtm90dbTpHoxXDbxT4/bJGJyzg0Xi
w5BvT6SlzPDba80Y//K5wBpF6Xd/o7Lb28PQ27R/eaclYxs8TB1pMwYRJV4l
tolSlaD0t293K9yaEzrvE0WmQfpHKwOdeBw4N6lctiMNstEBdGVH1IULrYlX
CvlNL/t4IEgo1S9rJXps1rOJ8XxwJjA+yk9ahCN5bYXAvjmc2y1f9HdqEYE0
p+mdHlY59qFA2KH9coqioICFe9nKx0LP8tU2GtBEmR7Ftct3En5UsALSYMZd
Cqprr6fyAREI6BNZ23sxgoEu7Z+omeSYXeEAAm7d69pyjlE03jIMRAIOOg8G
MoPz37cAZEVflWIkX+LdUN80hKauEF7nZ/lWXW22Vhrb756Age1VFWwQhDEV
QDmB87Zmb/5XSd1dbH3tkjjXsHrS+RjMIHh6AXXM1M/XMY5KOx29viG8h6iM
Sdw1cmtrTBDqkMEyZhjJX4wuc8sU6QfWfGXtUpzXkt9HvrTeAF4RHX2ZjrbM
uIkJ9Qabr2nSQCm8x3ZRDRvQtvmY5hZZfZgd8v7D0Er6PQ6NGqAOjd8jungj
LXv50tm/9yoK6GZ9TFm6e8pG0Ahav/EHaee80BFZodbBHITGNY18wVKVc1x6
gFng9FFotKaWHycIrmh7igfBAGD6fY57hBcsx0MLAsDxS/xRdRSq5JLWSrln
p3d90yCJQqGNOJlKDlBKlZXZwgKZbmbIfdEyaXmxkkbBudczekSBQovqgCiA
iBxapwKt0i6T7aTLhJ7ZaDiFRSu0BfdCF5hCI/UST6AwBflRllNwxg1vRXuq
ai/t5Xn7CPUvoEekJvtdbKJmMEyv7O5d3/ebyTSDuawuJ8KnFTf0vz2lSf+D
vElFaeRn4hhQNzNXCiFyjlti9ABDgHmn7zvAG62wjodFCJwKTggePH5PTJQv
0eDLS4aEZCJC2zYxC7F6G8JcA7ydqzfLtiocPetuwSY+4flbNwEM8qtIPx89
yLyCLsBCWPDM6oPv+n67EY/28Pe9zqen3NCsYj/a8DfwqQvsfOHpQTXuyvb3
TT79j3In9huro3Dk/b8TOqTyYjXWb/E+7zeAM3MXm3xdBqVvNODUKhQFmpyK
0Z5jBm/A0oGlW8DEjVFuNWE1VS+PBFXnfqibywhfW0ITcyMMl9Y2YMFusOTd
GquGE3abxGG528fL1jR3zxLGtr4OWkQXL92cExvs2ilQDaKiNY632oESlPA3
hKmwaHjg24J6eYH7iJltnTLdt0S2cOIKRkkDMwlLxPAGBZDY+sdmo1xvNYhq
GgirtROkCmZH6d79weHk4NEVL9PuQ4WuHUTot/vjLFH2caYftVVZeVJKy4BX
3ZVRHx3v2zL7wyENGsi/9kbcgooENmz1gywAWDEBOe1Nx8He3/ZmgnAknwW6
iZDS+71GKYLpfeUTYzNBUtzLvwU5+C0NircBErHo8g5OhIoOP546woeox+RE
6CEC/BzCv0v4n93MbIN6WjJF6anSfcGsxfqOyyhEoxF2V0uGyjFIxXLkd7pH
0Km2a/+FpTWIJmXCXPosjq24zyUN6KG2Sn3OitqwRMeWqE+cX/WV9GjIbygN
ZBDf2j9xtMGSQZoePbukZY1izB/ethSEbB8Z8jDJ7G2N/NuVS+g1xanZ0H+0
bAxTowr+Nq+NTm30w6EPNZqBOjKrzxKLunAwsNsC/HCHaF4oAGXr1Ztb3j++
8So7lOOMu6rfJFhG1sh2CAhEZiKAm/Ck8d3bpbSj0wrgDexzoEaU4dFkb14p
ZrwwMOwTbnzd4KRCWuFy9FpKYcPgC82bg8T63P1YrXiya3E8k7aY4jsAA3wQ
i4r7Ey2EdZFuyGXi44bgbqOIALY4tSOWJPQjsCCqAoEa6eG5HJGn1RjJ18W0
dlPD642CsXOL3/Q3P6J2s8WHjWJtXMoLH5Xv7f8/PlcVm7864s8zjlVV4W7y
Ss02+9cvII+749Sm8WrUsXG8XIs+cT4MwEq1W7j5sCzgoKQUkYKicleHUTBB
pLWjDyIlSfkdkUpnfPBLvzDQE2orDkxwRRnRNuKMNwTjPTDVCpBtwuFEGHX4
FZ5Kfq83MgEICy0nUz/n7C5FU/ugVTWa9k8iReph2qqhg/Mg3lxgG/ZYbTkb
Bls4hICLUu1bdcMTYWvo4C4dbMQA/Wb7chuPsLlfqJfitmiC0+T8TFSOpaD6
nS5UOezH/4L2Y7Vzj8RSQkYZZvAWDb89bIrJm03v+CD8BNQuiPj8GnUlwpzV
Ni2b261XG0DuI4O/SrjO0x09w72Q8/HpAnfhlnbDw3KxMQrhTR+czjZofjOp
G0TZqrGnjg7CR2V/1xGbsISorNZlyY1yqsFW3BVWBBIXNkzsL7/H1pr4CRHD
4qsuZ53egO46qfB503i5PwSajj50cWTNToNCgZim+Lk3j/uPhs2V4yj/iQpd
LHNEC4gD/uV+C6/cx7c9R3On8Xvzl9WLOxuPD0gQjqYlSibueDSGyuCmpyjo
8+kErwZzkWf6oMA19AqVSnphzfgaWkMiD1Phsy9c84ig7bQS9xIQ8CCyqGZU
tmO8GvhI1qUdzzgqhARvor1ZltxLRQI1NeJ9a+qhj/ylcFwNuPLfoWj5jiu7
uDU5H0uKTqi/eylZsfgcVyrsxq5sgbBG5s9Fl4zu7ypqWES0DKiqzAkx7PyT
5W4H+N9G/JHQKsXvf+qgORHiK1+m6VuWkz6dh+WHe1akSnMt0+il8zPQKk6l
9gOroUyiQozxMYQDskQJCFykao+AdVeGKLoq6Vq+/3RHPtF6BzcYW0/LJwzA
iiARhb/HrUga6ktjhSHqrqZes1UzyWW+ojPlU4HaEnvIaj3DDPd9F0UeYXVC
janK0UJ4bJsqLGWntHGRz1fDSgTP6F43bydt8LQEzm5xnndzol8XSM47v5nh
C3AnYu/5l6L33AHk3hPd2A1bCXSqni50g5O6FOZAGKCt4qwSkDkiyBKwGMJu
mSfnawVZdIxNcnRz+GYg3i0pKGTpcNQkxtmlhF/6s/ub6us2MYRSpHSIjxjQ
FpxhxDnh6mnFYj/UgFxPLKjcFVPWfma5iKjCSbVVIhwcEKSirCZaJ28elpuz
p9pCEFhi9oEIZGnNkgg6NymhUJOPdu2JUUfi6MiSI3GZh8SL5wED68/r5pjT
Lar4TmL9C7iPbVmEaYP9BQaN7qHu4C2P48xli3gj8KUp/V8eECFxw8nkU0ck
6UjtFJc1ccqkqWvQfmuRAUZ47HUiY+nJnI4voIWnsQc/ZWBeWGlk2ZBDNqey
1uqRUXRKk3uxR+G+JdQvs4HghWUhVzXUEz8/0ReHUufI9NfT18ZK5DL4yinA
dSHhx4eh3VujgfgOHczjSCApWx4X7jZ5pVUwaDZy4rQjLjsfr2qaramO7XkP
9fWI7GzXnxvf16bCsj4Sj84WcZkO8yqdaqNxzi3Ct3L1bpMOJBvSP9fKTxXd
XPztzkrlKK4+Bqgjg9S0vbqWfEW+oML0a6zrkesjxfUQyB+ugJXb7+ZyOa8p
2ZRBZA/PeVyPdF3RxEYt0fmU1lkdRkIqpItJZ1dZ1lGt//fg+d3vJfdXdgCL
U9PxZuEusaIqsDh24jrrAsTJoATEBgcb1u2PDzVKkPQJkzoRE398as5LJnlf
6ijUiPGGcSmdglkdqzc9foymIk6Blphs+oV0xDBsGkRdvn9n3lxbH2s0Kj33
XuEZ9eabaT6JFYT74dBzQYz4DbEd9RR8flPXAz6qv1A8iQfXaI0g7c0Fero8
tfw/muP3Ct3G9aW0tNV9IDz/Em8K0tx3NvM/REbXpf9Vp/I92O6usI+iHyX0
/ywK8iefpjtdEvlOV5u2/Jt/f4D0UD1n6OytgokimAkLL11DEwsXjhKay03D
ajZqEYK7rFBkSyhsj+cfPP6VGARUUTI8Tg47gO15uhEXjq+uL0H8ElWvjHXr
5r5jSHc3a8Gpjz0449qWsyhqaBMGj+VcOntTDjcf9QqFlWs4hGXvRVCVn5Pk
oLJX3NEz9FCl6ungN4cgRQSd5NZzkVxYtus87C+elDMiwbMpZVNLp79ypRp5
F0g8q6ILYcM4AZMs4cW5KMkw30W+h2wzIfPWIFOsJqq8wMsTdEvdxzGJcyKx
itZRQoL9KDoZtbZ3cduFWwzpkdMwkkriy5ANGWbb+T+x1YybrtbYDRmwbGYO
DPBfz1XbJd6nbVW9Jbd66jite/PdbrSPiF9jNU0l1DvRx9/m4L2rKJe+e2O/
7CPba33GLYLv9VwBnGBcc2xyitsn65a9HUiDE7KV3pfmbNCaQMJEE9WY/tu/
JUzG5V2oGUYvYte3ct39sgo/p2q48/RhvT0v5DJDw1W4ol4L8N4+YqO+ME36
+zIJBS3haZ7beSl5YmVLJ5RjX+4AxOyv6lLV709f0SqhyqQh6juT8qrIYD7U
KZ5UBMzszO851lriID0HFn4oDPinpPBB1HiBs8SyyEKzA3mFR6ldjug0lGsM
EOe8czYegMCvdOGd24jq2TLHwE4hH+1bgL/XCAGQwWHlUDytUF/8wbf81vDz
THKbt86rrjhmkpQCBr4bZiS5BrSSLCF+GleI60f1u60/2T2qdiHuBUfhV0mf
bj3u5QkzUhscvxvlyBLhPQyRCYlIwNZBRLLVTinarG9fePYCJguuns0q/dJj
v6OYKhtoGaNc6FUOPqsASlAYOjwYZNwSlNvFirsCb2md4JST5n9bxEcJeQye
qKTUKItKhPexMzq3CyFDH+57yzJn04aRIZ0cGZ9lgOAte/n/3JIIXsfwo9PM
Sctmlh0W7McVVu+opGBItmACxvoiYOiUUJh7BOeTsxGowW1meI1A8vZ2w6q+
SFF236TWoN/Fudm9pa1zV0nSRtJc6FeqnXcX5KaScvb8Pz7gJjNCLMtN75f8
1+Rs8MSbilAUBNlyLRimMegmndIPS3uMSSo/K3ea3vxW9S+KaOpoPIPFHRSj
1nqpWIWMS/oqktwn3K+ID4H56BxLiHiUc1HgSmo0hJAW1Dv+6CW55sMZXBjo
cOWu/US4K5GgOJ+pCYDjyFKH/b/9dJLhwP0A4PHBGZjEs2L8eCXfeUOw3xzl
bkf+/bVtDFKmUeo0wWu/UndnbMzamxRR9RDCs/0US9UtJa1lrId6UWkrVxc4
9P+FC1j22PG3j/DyZVbTojMqS1T5ucAMHvGR5UgfT4Krj5szwvf+Vd44edK+
RklUQIPqqcJez6MjZNdO8YFpHcs9V36w8Z+f8/BjkKWOo9D0yNMSJF2jf5gw
ZylyTw9IkcpD1ZofAhgzzdDjokMBy3M1BKj10H32e6/M4NqgQb+q6iv7NiLq
eQ+exBjjss+kssWq3flX/3bov5IVMLE5EyBq12n5j2DI/tM5Mq6YApqSmzgz
3N4CitlDr/lOmZTvTGaOi7Ya5xMWo2a0NHofGNBK+jhWN562fPxObiX4H03I
+1qRYX6JYmRTPHlcZ2d4sxrSQB+eMMCj5zEKD6n9RBGaindx27U6Xfpmbhuc
5T+zbUN0JOBxvhBZs44otY6cf0YTg97zudrdKf8UMiHSy01NALhyyqj3EUvG
jHCpyHv73uki3579+2WHsHUIPOdOmznjInoD8L9hj+9nbO463bSNeMscVmV5
RpF/N0PWtPxeGdqEAaddneOeNPFgGtR4yf2dEUpYXWD7lxLQ1GB3f3HUX6eU
vgpWTRYbDLjY3ZomK8y1DKIptAP9XPJEhrA7c7JdaF2ImutvSPq920bnNGpg
ou4ed5zZVcoySfI2bXCzKqAPUJcRjtQA0oWUn03EPV6qUykuC5KqKOrCtjl/
UT5Xn6ayNFEexyCZJ4y8nJZEhC/GaVJdk4c9zXCgT9kVSNnLNzer3slByyXO
Q4WnQJb8dj6IpDIiNM0SbrGOGYLmJ36wNjMIcGNtpNY6iXPS6zTjWuhX5bKB
GDW3YMmxeVGzrBV8X69/albxElEB8j3TwduXr2wMk7l52bcXDu4WeDki9kGa
i4GTx8N1Pc7P4BrzXC4PghvdGT8wYk3ifD8O6AdSHVhpuo9QpYiSzEG7m24Q
BwETeWYigr1OO0kwXv/TzJmSMxYfpvvdx0U+2JURE0Y25XLEsGr++ADqm3X/
8Bc6V1QGvex8eHMsCkIOMY29sR1j6fsx+tR7+9Wx/L5Een6tzZNw+lOdD2Qu
9ukP7lMrF9cCdj/GnfPZHDgKoAgeYCCG1Jg9HrOAxZbEF7qczcO7DDmJ1lib
Qk2skXyGEAfUlEXkkQ8GsqK7z4UWxo1YfWHT33ClG04V5VzLtD9GjnOCzq6f
9ogdVG0P3MH9ACrwqbS5mJvPB7pBBP9Kw+9xC3f8KNADc0uBYKTzOUqjB3TH
DFgm1WJl/4Speb/C453sYcqTXvubL62dJqGevvse56+6SdBtkLTx1/M8ySQV
55pP07zq8MG9a8AvwkGoPggQPFhGOGE/09mBq9o9wjoAbhbF9V4YVFzCB+Lg
Wy//Zb1fVwlGKqPTATVufQJVoQEyLaC8QcnynRg8Nq72cco0xTbpG24/n6Sb
ZHHxD0f7QscZ6S/u/xpgCUFQkVcEES1Ua4cq8snfD4rVN5HjIXibalIOGG4Q
Sc63jf9NI9Cu0sDIXFHLlDP/x/+vFbwMbR+XlG71Nb0vY9iCaeCVtYfRRAYi
mQARljtdc23o8Lcu79NGbCycEhF/XXD2oj0Ji3pkwcsbOBGioqPaQn1Fs2Vo
e4Qm1nrvO4P/GDWiKGA7Grz/gUn+EzzlL6MNhJW3D6uE4VkxQTTP1FNo3X5s
a38jPbyG3oXDGUBNK96F3l7JJyOanLHXzT5XVp0HnZW+sxvd6+/ZfnZIjaCZ
u8kM+gZpUxY0PPSy6EoWF5di1OY1NhRBIifPvvmxGm+7HBP1PlbmRJkuyJnA
EwduQSX9EkZ8CaWDZJP4XLn/y4CgKwjDd5qr8kPLE70OH5aenNdwyxyf2ldY
iH6n+mu6dS2iOCTkCJt+8RDJKMUgliKePSFKm/IZlgSIn93byg+R7erm1FhU
qGyEk0Z8+x+KBx8T8RQlhzf8rbyYRraAuaUQUWYYpN2OeSJmnLQBhvMKlEo7
PO89WVATd7M8AGPhuDpajvR16izZ80j6zScJvaNf6LiWpjOlo0NgkKaJ1Su9
iRUmXcjSxv7UwZusneOOiTExZf9tsTb3RX/cNsNC1hOx+ZmxbwORnmQWT3qE
vl5G7B1oI7Gr2AGUj2LoSRDtOP+N9aMHTnCnZDQg7RICCQiUdEH+sQw97tk8
8iBWKxS3MvLnKjbAe8GVd0jL5Vg2/bP5q2NgBbHliL2QbvumwNhAnDF4rLX/
h3BNuooqMI5NaJAV5D9q/YCXuDUz4FQkN/BFM53BmMeaT0+PhFeMLpKWkPbj
te6SJXNv7L0/t9ZpP83fqprWXIXmXoONMzSyei/RHk/hbH6IvGjxEgqF0Q9k
iFBVs6gohBpdrkOsCr49Of3zPh6TXXqADxjVWoEDiTaQIaxro0pF+lyi7Cfi
R83lsaUiGu+0XNUwyM36ENodfPPDc/DmHnKdb8dWnTWT4RjZvX/xTJGRanl1
mA0ieScgn6er2Xsi4cLnHImRlRq8oIxQyai2gYzzPNvi7JS0boQBq5vaMKAP
sRXgl54fSGiKAXbW2Wfo3fWdgtXj8Z/6bAgcLI2OyYX587Yyc+uTiJWcgxw9
AwGZ3wH4G0Xd0DtaPY7pW9xTsgxImYniHRZeHLA41Nde/z2VnUzcXfvOoo5q
oPbGB2ca3hh7llYPkEW+tiAiwhU1ePJJbfeQw/qQQzrobDU/UzPoWqFItyDK
K+D8iRWrQG8BcvW6pVtJDMxubGg8vC47yi6rixCCja8jTMcEDM/q4ll9CWYQ
T2uvop484X0Wgnlk6jPv6pPizf+fl4yylW7P6bUKbI3uIU499fpPM7vJCI0N
ivIkXAdL26Uit3M5nWrqgo4IQ0IHXBLIfoDfLRH5pXuFLkYPS8r7yZml52Ek
ZnrtDCZO8QHQdaVoKyHyCNaSmPnqVQQupsa5K+IGyVoTEOPgbRDwJWZ+7KCV
k0xaHMvTdu09hgZmLMfiaB9eTEbWDnr+hvWKjSUns/fkz5F2PQROVHslRVdH
zT0aWZq80gjaS7q0AvGoILKH3fMVlqXHJTo2KgrVSKSETULDYUk91xkc97bB
X4YXgpO4bSYN+QigaUdrEpiDrA5R3xxGTCQLyyo2/HqAvmeZsOC703seSW6h
WaI5nXfed6pMbt41cxP8UkGqhTrJp4/HCqUO989x+MlgfAr4MW3VqNFqx1sE
+oQtzjhgLMZ6m+3ymLW0lpfHccqjjB0pEW1T5rkGgBoV4iLKSBWwyz5aZU40
jzCZ0CjO8AJmERd5Tbpr0IuB/bRcoc1Y+Jph9nPLWoOwFd+Wis5SFBgrkB/Z
9MAM/SJueH6TGLI8QkAAFFSPgAd28TLOlWUO6SaIIJVKFXKgadVvpsMmi2pW
BiBW8cnYhd3ohPMXZKbqTm7NLEtHp7P+iwR4vRZRMCoIK1uBnOo7N2Ne0ZZL
fNemZt3SfFgzbFHcVM5BfX9+oKgXq/NQ207hvzdwH1qlPGbKRUzxTvDn6ioE
eBKwqOC7HYMeamqr6/qPHcoY2WSyfcAKtE0pqGo0isVbclcTfbnSnEa2WxsG
UxbpHyu74mrYTaiLGpXtI2fk2BCKbDL/bCXO93zBXp8CX5V26Y0GXrNcEWZv
bc0jHBz4dHYLyPzN0nfupYO2dUhvgJl50lC9EpJEuCKNY7UDL5260KKkZDI2
94aR5zNKuOFtvQ5tPRz/OQw98EEH7LxSRe/YTWVU6S+SQZ4kgcHtKfT/kuBh
HOoEScNPk4TVtzKC9qL958s+5XWABTqBAlBT6TH2dvMMk5aoSJN9AUTcjCmy
oxNeOy/ZuawhFoZuAvh9FWsm3wPk2GNvYA/oICFzovqJt+jvOaKLNwlhaK7T
lZ+yDMGd5y81SYtPvpzb851OaWANpFxF5dx6eXQ0omGcEzzubfG3WgT5lCdf
AjmaUIl+Id8ZvKBMjOWE+Do8x1xTLN8LFlWEwBljrQEF+WP0/gGfw5oLNxe+
MRRqKku0B3Sw36m08w5ssPTaTG2KyQL+tuR37hwKy4tQkm3zFAL7yV/Q1Wia
ciPZ+fglaHmw7DXG0nyGpasnVXi/JM3q6lYzTSDb1HeQEigJIkk/3eLq5cc8
KTQYPYtnsWKiUIf0MKgHCjBtrMaF0Sw7kRk8LauiBw4DZHJigwUwYSRu0STD
/F1i4ytAU0o0INVy7FjuVs0Wt9MXRFKaGRoevEkBO93MgsZDJjeAg0GJ1KfK
baoXbe64R31eYFXaAFY6j99g/vPR0KpdaL3VSXdn1jWx7Yfg377vjRfilulF
BhqW89l/thivCUqj+iiviHnWnia8uKvpf9EXm8kKQRHZEnQofN4MLCT5g0xD
RkqnH/xxEmFuonTCazaA3Q1z5gyuY7+UuZAtnJkIoXi+FTsVRPbojgWyFLgg
2WIaeWpH2g40jAhIWvvUfYPoBz7W0xUbbHcLcAq/R+iHS0wr9tQKJJQr9FTL
qJj5nPi/usgACBluAqrUG6/qJGl7IB9g4cUZfmXSEJIvx//AsMGpaictnjeN
QobosZpSxuBn3uLULM+S/29kZMtKHCAmIkxZ5d0u8v7/jIFS8/MC62uCXcZ9
cd2l1eyz8Soeb7ZxjlobjsQwxjSdeSAm/o03eCfujRjnr1ENofg+31bK78vh
YryOMuIBnhsKSytn8sZiWCaK1Orz5ZH8yQKAvb9vjFdfKwUG9s4HjSsJwyqi
YDW86mxul05aVAW7mq0IaNHCybAfclHCQZaiWtyyVRZk6hqdWrF6LYApX+mC
KFLh8VlCs8+Rn93Zuj4U1q1/a+mFjxAsrrfkUX/xOVQLqlkh7sUPmjAqdvqA
KUXp5YBeLOB711eFY4h2dye2vbf0LCL7W7R5EP3qSdX6TfvbQRBc/5uOP7L/
dEOlpjeGu3ODekBe8gbqR8etjQEWKBkG7WJvn8jH+wWgyr+N9Dofq+bEpPUj
HFnycAI5TprIJKTYqoH8pccSPoU8esJkotcquAaKtov0eG2ojQEto/g04/Ne
Y5VkcRW/1lU3iKFwUeOnhu3v9lIOwnGq3V6S1M/6Spm6+ucOr1lQ7A4soK2Q
LLu+fyYUApa4stFd3MrunZe70wt+uqr6YzT1rcMeHgteMghcgQBnaLRsvc6I
PTyxsiC6hpAaJl+JDH0SyVQheItg7wgK3aDwvXL2oA+0C9x5YfvJ1kj9P0dl
90/ZYcPT9cty7EeTh85Q9V6MoRSuiipruYZ4n2D9zLVfH5mFJu8oOtuIzFC6
RGP8KNnV3FXWyXCU6cEF742Kuvoecj7Y9FKUgzrRzBSVEFAC2QtthDrSLPp0
nSJL/93n+R4CeQ4rFqZU9OzKBVnVzpgQRRQcUutgO9pW5n1452fpC1rJ73+2
Hn83ZtcNRxUn7v8UMmmRQHUSDL9Khglmz95/mhG4xY6Os5SvyajiSBHl8Zpc
3b8kg8AsHK3/g9kuui4ARzJOlvKqJss7hdmqrvkw8Mf6iSD9DYK3ISC+r9MM
OD1f2xN9jDyOOQC+UsxbBGFwhfNhFGhfhhbzwSsiQpN6r8mpn0SVrzag4fHx
VOpxDJPixvbcxNnmE8M2bhuflwF7c+i1c+K/NjVGHg96ELxZEe9/cLNPdYFz
Azgy6w6iIuTwquo4fYQd7v4hcaCyO1VXsy8V45lNf4iVs+w7QIHflc5LsbG7
5oJZI4BfTaKNUch4IW+rP9Vr7lusDmpR0OPKVhZEa+3SjjXlZE57IJRzJxES
IPXC0RYHJNIZQwU+FKS32Gm0PTxjf6DoXrYCpoyzwzVNXR3/1SroSob0+Ct+
3hy5HmdCi8B6Qu9WNdmzHLTsv3yKnsPwp7nkKNvMI8QoVxXj0JqoTxo9XJvZ
NgFpfMoD3Pa7J9oFy43uRy16uRNeFI+86e2GRJLsD1QOwSVILBWzg90w66td
zBK09DGi22/59vTY/W/5UEE8dat172h9WSP2wG6tKp80sEAlYEK+cxeZLbh2
F0vNwreTB/kdiVvJ7g9zWQHadR7tooPcucHDj3hmaYYwUY9r2POWJB3HdYcv
OnIoCe0K/b+IvKRin+XKV6XrsGmq5cqTQ0dnOm8fo7HFXqxC9eafG07MRFi1
7zE3g7gX1P93kaQG7XvgMYX64MWfp/HRAMU3ujja0uFwCWzRo4bVFDwGxWhx
rWBxlsN8O8IMkIYSfqUUVE/KAyPJ0RIuCiNgJxt92RMjGR0PpTx3gcIkYevd
iIDFDsGhGezIcvSVXX091PKUSNFJ9yG+KYZ5jMoDr1ietAHdC5g+nO2giLBg
zgksLLaH+KPdDb6gt8ooGpFAesxpugWF4Uqxj8Fr13PMkThV22CXOyxm0hof
vCt5AeQJ1mIR2JPlaKnSwE+ZOYtfjx0z4dJFsagTZbfgtVqkB4l927dgLMoG
Ca5wmycWvGQRQ/l9mpgMDSodZa2cmnstVwv3qCPnl+D0qeOM7xntWabNvEab
fNIcLfcOsmreujSXhKwK/xmRj1rbvM8lKISj8Jx+WJZVlRrrO6jH5adLwcFU
8BYO5bwhC8P7/dbudxZC5IKwBpQuH3P7Oudiac0sFBzPEcNFXgqaPmrdn8ag
Bbo58f1rmXh1iTl/1CUQDM5dxZ42HPUCUWWnNvN/2+uiiodph7n18aeT9txa
Yt9/Dal4X8Oz5NNRMldeTn8uK7KXfWUt+843YIDp97lQ2I9E4vj97yZ244tE
TyRZYkTVPDkFe8nf2W/Q4BuU5fql/qeL17M/PlTTWwFwitZwuZ+kMduy7SiG
qxIN+Sc20YAyAAQhMM0nVcooOFBLN0Xo5zxLxoc2fwtK+16yTlSURwjQycto
iQBmHSunued/KBUCynmigzpToOJTvt8L9Y7C0Sa0/YRNsKnh+pB/ITb91hn8
2F5T+WBZGvJ4aPcniOJGMcEgmfpVkKT0cGEWDj9LrB6eOSiwIr1p0f7gpYnG
RbQlbVAIQetxVhOn2fH9Rv2caM7gQx67LflPZdn4igCrzaWHkzFuu4NKz7t2
ja6enq8LwRMh4Vcq/Er9o4TjFsyVRi7hbiKSmS4ba6e0aCk6ffZTjUGLbAr5
lmfZheOPLlfYdVjMhKTIKqQiHFKChUlJLtVkoc9dctCxgoeRnVHgylpO1Y4n
XSYrzuZt/gIk75eHjwCArknjAi+CH1Lidx/isHyeK/X7DB6tZco4D8cMecFK
CHnJHEMyJxWHv6edn5I9wTpfSs42SX2i+Aef0hRuedrbVYi7x71EFfGHU3my
EoRjtQOIuXdOMK7RBDQD3b4c8CwIiH2aCaqHOxJP0+v87eUiYQzzaoBIShGa
oYfh0mQstX0Nmb+c7Oj1i1KvY3pgXcRA2mOYO2hEaEyU2ERhk2iHxGLgNCgl
/duUK15ofhwT0kLhHBpUcQI5ct04rgvgSRsZemgxmB7mhlajrIU6DedzmUlP
37x6UvTYXoJhYj9ZmiBX+5hYe7nt1gIUNDtkv38NX6pJ02BrQorXmleQNeBW
E034FpGiEVEEqIlvDEJWUMSwS0qSMSvJhgr1uKCRk9fb593XZZvpso4Y3YBx
C5PvS+GTpxQkJ+XukuGO7LLvjmoCr0tP6TBkPVh7q+srqKVDP41lDapVNMxs
LSD0xxC1S3fb+080A0qt9fQlqLQjYtpuxTIwtU2oea8aGQy4gHixlf3MqiOq
85nXImma091U78z00fAcB14s+P4w9d3vBySBK4fpZvKsMjFudeuf6KNcr9Xs
yM5k7XyXtVHochZX0Kp1qtP3CSgowizH3ESTjl2PGXgOp3HX4/UyS0UYMZko
wsVbwtgnJp2dRFAyJjX2znBDrcHzDeOzfxvhu79rY2eHcBAoeIro3uw+4OpY
0wzDfRsOmC+pwb5dS58VPUg01Oz5j0O1aWjYfRhXomws1IYCCnadu/rDnRiG
Bh6pyy/Whuct4fgmx50eaElgHUHX5cJtMbJ1xg7kb2OiARqXh3L8BnPZEPVD
s2hfGqFvYLS1z4LjxVwdxORjEnUfiIDh4Jvn//ZGq2RA0+D7eFti5wuINXBW
hdu5IEtf5449HTq5mpiXqVcZYRCJnYRPD0Ag/9qKdwtxD6dw5AKH8cgZlo1w
uqIL2AGeAS6+9qPOmZwJVdwshqf8VIWwdG341lV2n2VZs3M8q74MP7ifpKNM
mgTEPEQGyQVIm9k0QkyuunUNZF7ZHa4bcgrO7s+R/u8kMncZMYffIat9CJTR
3/7d32/1tJXFPkdDsSbT9KeqLARw4wtUiGFgrinMIlpBD0ae2GK1lZZ0zV0G
QxRb12AGMaineBGeJDUBPwVGgCUuOAhK/yeoIIyHaxtY8+nIa/p/rtxEq3aP
CAQnLmUVf3NJPxossWoBvDCr9p4NUO23IWMfmp7jPV/swvoHK7b989iHm1LM
B/V3XRbVlzunXxz+In9z7HVFyP2kKai9FWtytiB8/xpdGBZQdktr38sfyr82
jJK3l4cAtTbdS1jS+VZdJmq/UB0kSxOSksgbSil6x/Ewn4VIShMQ3li9ybiK
HRaqK6QSCr01FWDG7Ss+ycw/KZ8aLmuJ8powgKfUpLzzPwWAvpl1z/554vsx
16d/nIdJb2UISKZTlnV++ZIEXG7IhwHKs08qlZL6+FVVrf9aMGzx+aw2P0w0
foAeOVNVUaOFlUhRPPr5r04Y03vNZ6X/q2zk3mBUFgDTMKZxzps4gdcQl311
QaSbRt521QjLLCHJ8hSIJ+26BZUGPUGVw8x3s/i/FJqUu/CzIfdpJbTkfJgO
rdsLdKduQ/lyqJHYxcY+ePL3ma5iNqbHGeby2dCN8CRI8X1q05g/qgiYNsR3
fbUVaQJARbs07RQXTYnb5dRqfKDeAhRWuI/ICapWY0PcllL/bi6Va7nT2ggg
IGESzIu6zTvQJijYyoBpvDUkdWWgltzwcFynzdTTavD0Zh2cXx8usgryJ934
JYQBBE91ZPMHgEHHVbMHgafTZBsTQb5Z8ii9veKcNCd1bbOo2I1q4R3r6pCt
fbiksFdIV5+do8a0vh9KbpzHrwX5FTI6xBXpU4ROhZNdhBRr8sBXVv0kF72L
gS19g6uoYewYZedI7sGFc/ZEe5sfDu3zGgNcu2EaaIHNGX63uvkW9gSmRiTE
r7oTtQNwXqxw1u7iizx0drd4nCCxdBhW1OBxD8+1QCQpm7fkYkAGQiPvRWEV
dLOUpUd9G43JBWlCSejIKmX4xdxKc70Y/pkNKyoT7yjgrpIDPDWoCfGGIqKm
yvxBXHYMhJ/uc54v9CCXZmOqPc2SWl5JtYIhglfgazDQhfeW6bCUxqv9Q7oe
6kkVtZuPXQsMlC6vAODPMUrXln99XEhZH///zend808ohkRBp81R/nNwIeiL
1L+6fpxYnW+HN3ZAHt6m+CpqlLiAImVr6nBpi+XzvHJ9G2cBIV6UHGHtewoB
7LPjkFBi9U4RqOOVyoq2xNNo+WjmpSXPWv/RHVV5p8YeeWH9uY5cdBqedq3z
4K53eWKSTr6I8zLb0VKjBvlDBZHQvSVcth8uTDIWMc/HS1SGoqZg1dvQCcV2
E9muMd/QReSrO9wltalWrm+srlY3TgqcZUm2qKKjF6VackRydM++65ZSI9VE
YiJvoXGcFMfDvel8L9iiOj8JUqO7sSr0jhTYpd2rkOdrEDIecpJ0GGBFObv+
Vu6EP8f3upZnZGL7rpkZw3o4BxmBLYiADQ3j3GoQTqCtDdJPsn6anc24G/Og
1riagkAB6Y0Uf5FzD+OkGvroOky3KX6cE80xuc+XSpUu+bpo6lrmzzSpvVan
Nvbnj1rgyqjyvr0pb+1WOTan4VrYCZlRlHTnOYPBQahW/OKgZHMtnnUs5m98
AQ8mgZBBC/+9pELI0YFWo5vHpMaJiZiB6+N2EXye6qIuyF334e2g3ao4bgXT
26lCYlnntc8xz/E6pxzGTHVV9sG7c3weWvl6JUKp2vFWhM+E13D/ET5xoTMx
Dtnm39Fn6XhES/Z2UzWGbKFizH+nvngK9DLLRrc5eQCDSANOz20ItI6fLjAA
LwBw/HT6lvIbqXCXWF/13GuLUo7SLrjLan7NrMYUbn56pr+n2k7d++GLnoeE
KJmWwRHgnSAl+ZA+fUBX85iUJfUwDLby3n9Q64lUY/9MkDDoNyKM47YR6U/C
4pAK2OL0e4Sxs+aGs7fBHw06RZvYeqaOYnTitfdw4ipmTY/Fc6W3bbfH8b+e
0lSonHbziPyXQ2TYAS8IUIydWoBDQUZwzcWQ3EhOKi2PsLz2zLVK4GsLKfQa
33Bob0RmC83FmToeDB0tc5l1/ksAvMlL2Uo9mqULF7bNzYhwzn/MdLK2YZ4n
0iJBOL4gyjUp1cUrKQW9rZVtzO3CvaPzpzv1psksflM0WIKLn+gEgV5iXOJs
3Y34SzhZYEjvvxk8tBX0lk8W2IL4X2Gu+odSIdKppsaKxj0NL2VKE6rQyFKv
v/zpww7oKPpq0jZM6/jcak1TK+9ZfXrC/LgdmMXlD9sfyLuV3yPBA4cY+tP+
6Kzs+PwFbMXqG6MkFBQWRSlBfblg4vdlEvZbKd0aMuw1+XgE2LJcz5JWfAPB
XrmUcL0eEVN0eNteh7n78vBgiouliE3OMXQByz5cs8ticdwJa13gC00qE1kK
HeVYFTvfTO5wD8aksqOdCy2wv0Y7JEjeLxk1E3kty2g03bzDkrN8b/Fvs0Ia
d5fzXA7oXPE8mMtg5o1IekstOhAjOXWZadvK2o8pYxQFuuIAsnbciEZ9lf0C
Fhv4Rc19hxGUdQgARbFd0TGyiz7mUkU53P8mPYe1fKCEJ77lXbIqP/MlsWd4
PVBCqidxgTeiTgwT4Hx7EFebVVeaTZeNDWfojfqcHRckbg83bcSF6ZQv/VXE
nOYL+1Bd/dDQucrcAB+2OtARpCvdcrjPfW/60VmcRD4GECV594dCRIMHmNnh
dFwNrIHmAVTeD8U4HbS07YLltkiy+KqZ2hKMvJwRvpKwd15MAvb1Y7Mxhe+W
JKAC1cuv+u4Q/JCsYUAlJf3iCpyJmwjBUCRD6eOL2uUp5OvMj8/+QuRPR2My
FW/1Kx8/eiGAmaDWluAAfR0KeohgrlHduJW/x/jjk0Rl139YxeIdsJYt3YhN
Syt580TpHBFpRe6wVYKRRxUXyCXgY2Aqcih5iH7jbNk4cVvpzOfqL3fvJD44
pOXROa5yqUCzFz3N+H9+riO8pnwmC3o1RSgmLhTSh4Fbdwj0ihrXwYi4z5+r
0qEiOCZ0MLSTBEnTTf47K4vqyG0kmFpys2wPb9IINaKrEAg/WA1HtmriUjvV
RmVVR3TcDFXZd4PP/J6NxbHRGzN45ySJKYXw0ITBYgA+EqD7WfUsV1CVPXqB
K2eXRBVuO4qXfA9AjMZxoSI1PpJtNYGRyhaVuxMyDuDS7B3sSl5DtNR6FlWn
x5VwhEnliNJG8Qyacvaz7FXdMULREqSpNbArQIBcjKUpANdkGOM88hR2lFLu
8nSoLfCJ58E9qUO7vRt/jAVswDjvzUu9kVPw9Ux/1D7LehkQpj8ALTSjceiw
OypyHqmjWh2IgLPMMu+HzCkXTl6+c0+oT49bl9Fp19t+HkYZxFYXswyjRKdm
GQTql9VQrtJOLGiGE68SVWY1BL55eLWJHhLa7WzEkR/nMVm2meNMph1y52k+
/KUdEluaEGdy9gwaa+tUEzjQ4q5M7DF6BFCFd2cCcfjEQzSyidpBAfbWfVk4
C7X7lPLIVNLVX/RM9bir9xaqmiCQGoDFGz32KkOKH883TZWGIVg9GCVOzJLd
X69n9NmIPubk7RrEhxkmWSyNSFCUD8fOZz8Z3SvRrN7YgtlGp+XpklqdNz+i
hi5l7L+qKWmzn+fxjpI9k38b/CGTfE4g/fSehfQW/caIkF9GYq/7TJ8kpov2
XyAiZHoaMkjLLl/jqEOzxUmhNv3c0XOikeKHq/m4s7T0phwM9j1j5Ef8MYR+
t/Poo7iDkZBmwgTUiVcRtZp9hJeRsjT/FCNhpzewfMIOB+mNd2HzlP/NFtzT
blJWLZDUOe9zaIaGDi8J85HUxuzVu7tdax5xcI8dE8BaTGkbWx3+Xpgosszi
jt+3+7AyX3MEvyZViiVhL1q41SfZSzyRv13DsheXBnoyEMv1Q2sba+6bamCa
jhI8gslevz/jjyZD49HD2B2ZBvMBE/VbU7xZ42c9Yek9VJArJMQep4oHxHl1
HHVisXrQbn5cfDqmskZHIRPLKFJ+ua5ytFL8rNYXkoixFCE4DQGXfmDTnZk/
p7kV9qEAo3nI7xYk/ErPsHeG5bSwe9J7GxDho1w3YRAE4s86awvnADAS4Zw9
iCXB6oubNdG6MMR2MSqSs8xz8KSYKl5u1cZlpDYM+utBzYPZHRwm6cn2RniQ
96eEcAk4zB8mU4SAd8IYe6tGmT9ENV3QktFochmPiRqO2oEcVWmenl5HZ2Gr
eZVJjg/AczUXt5GSXmuTJ51RVQMYwEaHNvRrEJ9pObS0Zo6mEQD0FPwzSWEv
IPxnucyYCIPKvkEeNsN8oiM0LfY74NmBBzsI5GK+7qUoC1DvKqZE6W2CqwSz
H6sYQYOEuXLqDK9hMpEnYoIXtz88K6G0Sh1F7am1skLGvmxHndL0SJpLMYj7
r7OhCmFXGhWJtlAkDaUtG4h94ug1BCvywBr5+OVDkHsJdXEpbpKBe96HcGrt
+gYFL5ZIf5mCIIo30btm3uiaXQwdVsZR0fKVcUdJKN6zmi6vGE7f4/eQ6EQ6
9hfCelwcMNXLT/KHxIzcwGGsRna8ZHGk9Xz4NxEjYH0zX4bmZFP1dYl8HLHv
WMy4yvmg3kvLvTge/oGsdJNC66bGYQA1BzOWZBILSH9xAurspvBwuTpJUzvh
ht9fCD8goGC0GGBaFIuo+cskMFE4YRPbal9sXKJhOYD8TRSsTB/btkyqLroS
CeUczwkAMrM199a8BRrnvLbB+5pkvRu5aTp7anJ21C6uW9GlCaGHdfMzqg33
L3gnxvcJHBCcMolxGaYDy5W3ThaEqPlh7Rd/s+zXq5tmTRjbuGa5nM3B1NV+
BLPd2OpjK+sKJqTs254ZXyj5PPn5SxFCg/C+KkhWrGxp5n1rOqy5DWgDpCh3
W0wf8tti1ZSDsxE/nmOX2nuJ2STQ3OZLmEEttrmAkRgQcp13mIH9kKDnUaJx
0N2WrZlasytNtLGHtLuO+9IQejtysV0dfhkhnxdoG8ZGabCH2/zmO7MCb7cn
oD8oDb4nFNBjcwy9bDbpa8klpYFkJwcB0onaoOt0HA2EkQcYIv6CsLp5xDUW
4zzAd2cbymwTX+CibduJpAqJhhJwxV0kxfjkDOZe9cZ/lGEu378Db4fOrm5I
bkJlR2nK/2XWJF3j0x0rIFzrxMqzX/Pg69JdgOVIUjyb8FrGLr5oxlbXJGxr
BSG2yFD9fubE9Sm4e3p90AblMsylIKBTmO75IEvz60fdJNvketrl9rBvMMo1
cfmMjiuYju8QpW3qEgTvoFw6jWZyw1uG13pHjJMzYQ2OpR9whrJhDtZFK9Tx
qFxFPeEulzU24z26iazq3MPfNSCTm0nCa4yVKCmKsWFUXq7GVBh2+pV+VNfb
LCxrfi0lDuiDBR2BtylPXRae1BtU1NlKx9sDWOriaUDwxak251qkFvwcYqo0
tAeEHEYsaieqLByV2u6oL7SRwOlfJi4pdHP+9wazdowCRbMSL/9aNCQ5MOdR
lipGIkpCpy0LFxJq1s9kYUj1L13PMMgUSpC29oITpB9NqNM/Hkq1VjuZW+jh
UX+WLv7uJq77bv7xpRkZeHtfQj+68yTgw3887szl9oXGBxigltz/bWRvUSYG
pAwrsAJoGZfSpwqm0EJhmlr1KxJVhXHCPgbOy3qhlUH9kolBQSz26ejPfVx2
927EqIbT2lKAxGq5S6Qw/kwCJk4Hsx8/1EhIyGfETfy6HYq65srkgQ7XUsUu
RWhqxu4ieGNWV7PoPabRu6ycTmvIuvY7BA0ZqyDXnFP5KvQGx1OSnLdKzBSa
0rxyl2bHYJOdOJEpLjWcS5Gs61T5sShhyKfsaSWhdSxQt/jWZd0PLRrFNKSN
0WwKrvs36O+7mx0NwDGPYM7ccGw1uROYkjjFn/tc3oPa+46+93Gt+qslnMI7
wxteodK03U+Yon/7o57TB6Ms6OB0/PIxXJXGQd6zM8Wbzka2NH5HeSJoUZAy
cin4XittovPfzuxoidAK+0R1TzxUT5yw1a2s4fcza4kwpnTMp10lO0hrc+Qy
RaG7itbk7vDBBE7L/GhvBszi1RSbJHG56DP294/mnAbmqJPATLyJ9LBuWtEu
X+dlHjdqNmAL0+b2EhF3h4Kuq69Vdw/rkMlyUxQZEibIqNvv+IeHR58BvOv8
riITbsGfHX659qRdGYNKw4rEe4B0TBZ7k/df7cgo+MHfmfWq9vO6DkEENXTA
Y5aRBDnux4p1bAtUFxaZ98Zj1GJ8LQvL3edpCPsppqrDX6bWojS1CG6g6pMH
ZwMo+hS5Ql4ER7xSqWt/2L9qrafBar9c5O+YveqS2ZcdglAK8pbATv8Qqedl
g7cWtej25LYtLBNlwRrsWDFj5X62ZIVhD2ka8LUe0IRziMVSIDqdYvOTZoMS
DyCzzAURHPPTO+HWThf+l4jDRkLwrd34XuLlu8yv5dK2jaZaucaLs+rDGP/Z
hAGvBaxToyU0O1SFLW+XQq3QzzfXESLO1xlMgocKzLcAijqrbAxSeXrnoXlO
0U/fbdvO9sb6lj4OxAKTHSqb081CyDoMaMirp+LBHvtS5frtNGNJqC6K8ucF
yjUlbEbqx8qt7tkWqOLlXDOv7JY8w3gT/rQbFABRwjWX2cQg6FNTY7PMV1z1
mHpBDyVOd5/Ubh6ui31eAIsqSJ1XwXfXpk+eW8A4My0tVvAE9dP82UB3OFS3
NA0HkodkyyLgI1UuzuqLXumPhk0PtoYlt1RYzb2lOdQUGFXhRQSLXQHHMG5O
jINFXP7vUPvl6AC6h66U94Aj8fqIpHd03BvfR+5aCyDArMQTdkbaIpBd+6jj
bgTiNGUF6kb6hAXaou8Ot17p5ieRPCwlFwibM+thP9FaOe4ITPBcyUo8CAwo
W0nvw6nZWpU9ossuy7NeefMpkV5xw2emNbXNN0AtmF/CvZeM/ABEf4cd7vvz
VLM3deB37I1llCLHc4203bNP/s6UPYthCxxXVH7uLtV4/hhtFme3zssKYJZq
XmxkVgoW0o7lWGoBUmm6nBwpZGrb5XKud7HCvT5ZgQteRy/ovvrxobUbSm4f
mKFGrzEa5ArYRw+zZeg/LQcKaewS6TMcrW68X7WX3H5lRoovkB/GgVH7xhC4
tfxni7VqKmC+l9BoeTIJjXSYFpSIxU7X8XZOoAPgvheTzBEPR3I4IyKWZsMc
DwD3DvLdGAQqH7wKAO+HOkRcoPArdUYecPpLnaIyZ0jhvKzDlDZ2GSqOLsK/
kZ8apw8xesCn6Rxr1mq5D4Nh1vvg/Xi5gxLF/wrZd3aWonejIjGF6E00jAE3
zyR3iqVfoFvGMOO5ZLHL8OT8xuOAF65700yM5BXioEFABQKY/ek0eKkMn+Z8
Uoqt0SXtojF2o6AAOsk6cSAk0LFPgx7MPMVFRPfbO0uJEOwktah3GVDzoO68
73fxNcnmxd1kyzkH6cRdb5rQYLRO560mgL1zninypmsHiAYKwvCmS2CqiSdJ
EyK6qh9sCKAQKKy39bv1+avsVZhQsoWg+wTNo+UUVubQ6/gW2Xf1P2HGZoab
J+4xPhvLgNkw0l/jV5/33IVGUDB0zJQNLHmriYB0zMEB2J0hrbsmO78BHwYf
8iR1B5fXPjzRrU3aZeA4/NBz6Yih2/Soa4hKCB5wMWy6qhC4VfVekxuT4UEo
jR0QQ1QQQqtlWsszqG+KaQAWW53eTa56eFhbNPRq+Gl9N6DT9jfHpIxx6AnI
L7eM/Lx0mDQ+s6Sh7bS2KBAxwUQ9uUYAWLdNoeN9meIAfrpbVj3PM7sDH2jk
XQD2OeTXbd41RiRraJn0Bv6K0XkNtfLd5lPG3sBlrS8WPqikXyW8xWjE2iLI
r8F0IHd3Bl/FAQSAwiI83LTfVRzJeNsM2AZr3b12PQnbQ7nY2n3ntaeB3R9G
EEAfOdgJOZN0sgSg1VBrHiMSbV+qQLOQZ3q0Oe3rl7Po3T/21QJvW4vIWVrP
osHCZVFWC8MgENEiWEg4RVpgLtki4eXv4laqGEUQm4/l5gylfmcO/PRx6nwI
jxd4iGewRUyOsdy0tqq0memAKhM57pume/N+eQI1MpHSA5AO/FlQjUNJBiwN
4TZtLAPo+iUakSCejF35Sgy3gNyHHQBbQuKiixrOiQ9x3yZRM39fBoTNGitS
p+/GSKoKBTLBV+LsVdVhXeAdll0cJepdWlMJQiGmG+4QEzM4IYe/geC5VeU2
aQGFNKwDassWkbADHvfD4ttIBL1BN70EoldNK6+eyKuCOfGRf7ykyG57FzBl
KIekSq5+He34eR6ffRZWK5m26apYg/WiSEzyvNLMDEOT4nsPfTohev3wg+BF
1aFsiUOPyo6439eD495obtRU26G010YhZ3HZsIkF6uJ3Mw4ZMyrbpsNkvLCu
GKf/DCzP6+Hd9bjxvmM2RrjQXehjgaYluhByJiRIHpYcufbWvQ7VvzhYgq+O
NxVNG2AtlFt4d662bVoRf11VrZYw0cPVjbu0GEBeGfUpS2gbU/aLzRXVobKe
qONTx2Jmhk7VBbbS5BS8/9Fo6zF9Zkv0YLnoLgh0mTuwDT7USNiQf9e/d5mu
Nw0d6zFa3aSEsN1P7HA1zCAm96hfRXZVyddJU74uvRplSGP1kjCMf323l4ef
NtPUYo+X5lPTWXDPyf8ygDMFPlJK8fPeybmrX2FLX2WPMBiwEhH4zr2UuL3a
Beu1skmpKL76G3m5IVDvHgWCxhV9uiGmNYFO0/RLL5E8NvH7XH/sKn0sHB70
ORUU6i1kOqZ2etSsCOGe9NUl07/NEKyEbxdxfDNKBnJxdYc4nOxSWXQ06BU5
cvVBQ2kcpgeeasneCpfdDMXD+fDW5zbQrUq0NIVnF8BWDxLT5Y4zUCTQsHJ6
aWb+uwUBXaR2xm+YSpPXm1qK3tkOowiu4OHmirTUP0J4K8rqR3rpUaHIwYFp
KEo3v19g5rwHc3LWuFyssbRvndtTXbaeA4Kue0jV1ZUSyvwXRdoM1L+s86Rm
8aqQRZ8qRmoLgUO6znZDX93E1oSsqpBk9P7ogrNd8VJ0OmSLZuMMJCJxQWeg
rZysD2joltge9z17eo3AsqGxpdRK0ghqfcKSKuh4FzomaoxcAKbBplcu08s7
x0XBpPyq3HT0fIReG3XqOSOr8sToz0Lo2ouNmCklGzSxz5EJaiN00LDsNEwF
3vOB2cj55Kh8z3GMmjnP1Fdl7pS5bS570iLbcWpCeAoqMTSevw8p9gShSsj8
H1b+swTj/u8Jz4i+KaxcNe5CWarblOJcHVaO3NHKMaIAL+ZbuOswTiIt1y/Z
KJ9qL8S8yXZo5wPzQQ7Kbi8mSmuwi43z4uXgxgbpH8d5UWCa46hBS9Owys0J
Db1pB7s13DQxnBGOPRoFlHBTNEZMVlwrH+HdjEZhFvJ0T/jyEHSL9kFsEDMx
G8T9bm6Q5597adzwBsS/l3wyBxrwjy12hqbDcCmch5VRE0iOZt353EwDnZgC
N/1e4023t/l8ixliX6faRFYMUR/3epYPhtRn93UrGCWSmhW654AxqkUbCT3j
x1Nh5ABrkqIj8HTmWDvUpHKjH24HhBayOy2MjgNeKfh+nswy/j7NTn5+c6Lm
pLwtvdYDMmTjD1NxcrX6P0xvywjRzOZO/JiX8ocXCRQH9gk4ofeHkc2CNoCq
GnOVPDFhuCArR5CClnOQMup+lveaDJVjh5AUXt2fFVDuRBub3Ya/QON9QvAO
1vfYSg9NMb4PVQo2MBw4H+zkpQ/GkjoY0ZZHazZoGRKsLFFpaOvyNcYl7H3V
xrbrLUz8zWJLJ+w1o2CjkxNyYrbx/mgnSVjnT2JHiRL5b4xQ1RvNuQnuF3bN
LZDF14YRVN6PQ4VV6CcWONje2hXOAzBvIpWyuYjtxOS9rgF0Y2WxnXJ4VuF8
h1xn2lEI4qwVRSUa35y6yUfmbhgiY+yMAfksQ9MYJDQFIUI28c4PaD7ZReGq
JohTtfnlYEMorwXh93yD7KjfuZuMwfg8IuUtlaCu0WyfOdnpvcJksrCn7HnC
llN4YIplmneJ8HfX36q+XMeXuoKrnJOdcySP1fx7QiuaaVP1aiP4pYo4TBxC
YY1K7xK/7Nij7udL/lh0YJIWSpDGKkEJkBGtTo1bkcZnGdovdQttFtNh7Phg
5LfHgeAQwBxSx1nPoVnzAlQRey5gXlkmDluzVDu+6bufQ9vlQ8IPVEfE3U1r
Po4OIEovlxRtKMk5IqSEHTUrAWKZ4h11eTin/1QlZ+BnpZx94n1S6n4BBsvy
TdfQFghjvtw3F5oq4wPpyPKkvLCABavq01u79K94khIiTFD5b1peRCMxgOzT
a9UqBGXlprYTIytZOieUM5vRlKfJLdUXw2yUXcSOjuUXaERH28D93URX48M7
jnlugZjUVMdsdBsw+ntOuV8IDrKfdEWziTBtg6Fw6kQexwQHLqT2iGZw+lRU
9znVykspHiKW3DqXnMuZtUeMtMXqh9xEgi6fJysw/SPKqAN+8RoI3Ioghyxa
ROOB3+fv+QG+tR/5vNnVuFlZjrACTb8NRoqYReisNJp8WE5fB2QeiVsh04NT
rpwcwY3yQEF7HIM6uYNl8JrXCRE9IcOFJR6WuSccU0UNj7PCgneQDOsITqid
X9SvLOXFQDds0hxhNbAdwKlkHXRfa3zvPDzwTqu9xEgT2z/NLcaF4sfYqK2h
Gxsq0nMD3SGCbJlZZhRVgNBIYMgWc0mKXHacXiLIA5Tuco4QnL1AUq6rSN5t
sBhmDnTmbouoML8G3/jxgYWgUXyjTyEJl6Ha5mQDcfTPOyJ8PxGP6nFXyzkC
Eo2Z6V0nCit4DaUTgT9dBiIjPjfxSI1T5+HxuMBTjANL6L/640Kys865DINV
8U5gqIb/DqdhWiHBPv6ATVOLF5ffUK2I8rhPPQ2vf7MZ3/Nvso5U6oVLLJgc
Uzeqm8uKa9Q+Tis+4uqQbQMzaCcEoEmftSdaisKY8bM51CGrlVZCKhwEEiF6
knAY6w/WY5l7sPV6hWukktEquQhtL/b9czl5JU9IvztPQwjH7YnUr6DQByZr
1ZB3d2SRjOKbyxGdugyufpRHqKuFb4ZukKTnW47F5vzQsTI+tTvwl90Af91Q
aphQzWwyg0c7hhB5mv5LFEXmt/az9VFxC+3vU+ksBFC9QgN3FgQrieSoYce1
1LZcR1axzDl6f9NKlzcKxmFfhPU66heNQHQjA2wgX2cIgJBgq+2/QG4n7tf7
qr4BM3Mh0FEf1BAXdfR3QhHokNx9YWsDzYyMJ0jboyHz971jIjnFReBP5/OS
l6UPgz0eRkXXNB/n338KTJuQcdX1NUYAcNApqdd43jn79RkjqL0QPyYRgD7c
hIHXoBzkN1YxxgK/r9iRxrdwrcxs54dMvAMhU2YEhVfGUhjFw/VvzVIvgoLS
4HwzHbUEqZtC54umDNmaaHNr7f8be9jMU2IMb/OOgpnY/PbyxUzOF678HaPV
/ddCWZOLro62qEMIMBVfEBNb4/5JtDpfJEZvbXPJCx0u0IVUFw3cnJUEQTxM
KSxZ3XXveaT04K+imsoXpysbJptrrnQh0bGU8cTVfoQl5Ii56UqXPopEQwsE
32loq/FYm2dmp8CA34mZFQ3CnHyzct2xThgAWmqPpr/dP3yA0ARG3haOsJ4Z
ATUbjZmlMua0gBIadI8h5FocGNDf0SxfZcgeuNkXs68dGqx5gIhYpSuDMqf1
8oIszUt4oWeZspimc3T/Fkm4Z7WCDPzCJa6AFCUsz1vtj53Fw8O/i5qDDnfS
pbk06Biqwkcj1wXSfFY4sCfs/Rr3QyGW+XWph/WwkIF5qtX0KytvSAnT+g+9
nHSDfFzJmeBu562YgL3rcTXLnj0/MzVq4Y0VUimt9pVqYDF5y0IaxQBNFzSX
d7kteXJL+IU/df1A4t+0tVcqSTMWVwdA/ppdp42Ichlv9VK1Mp/M9H8KclkX
fqNlDysN0qci0/4BMP2l9igtx/c/Ixer+RGzo1xWe5c/9HdzAZIeypgHw3h8
viwVyNZMoIF/IJF3YJHdCR59ShXDDUjQBzs2sGqimGz3LxESVqalr11hNzxd
Tw4T/DJ6KQkmupEROOkogJx/v4yt82g6Niualaj6QdRVdMnTIXHBR6YHjk36
pjGj5m5RiWqL9ovNvantLWRUUmoGbrCuZXbUzBu52ghLiBkZyGoCJ7y+WgFQ
m7BCDsLFr7WYA1RJfTpq3qJgzmjY62/jrm2MULW6HnBNumhiZ8liBryvw8iC
ZCOvVS7V7CHw+fJ4JLYAma/fe27bbP2wi0ZLzAv5byQsXrrquWdoT6i1/gzE
f8pvayXzrVTiditJ0p5DM8PtyQ92mSkK1P/L1l2ZfrbUVvbv6aSHEonch704
3K8nXtaR8Yeu/WwusbQzvhw6j0DN29uNfBd0X1er3vyvyjPg++Dw+Q0iw71x
IeSrGvbvz9y2uu7DG9zdLSLleCe30pMfI/2CKLjTFtOz6VGQvhNUr56GtzOm
7mmdj0qBwe27zuObSXKHgywoQAnYXX/j9FwPs69NU4dtfFrAg39JPUUjJljR
6VnjPgtBfnqx4Hd5zrGMEvkcr78/vZXmmwTybodLNsA11/K6wGTUejb6Rsjk
VQoLejH6lr11FXb81pbEtOg08yHtSHgudi0+wKgNyp6/K0pDwtuZV72AXuTq
8+xJlBXW4SFFnZcuRqsaDnXqBa82h8VUuxoL9FdLk3CwOmy1jX1wXqqQHKql
7Nvcs5tHg5FgztwOBSqBmD+dKZlLe5gxJHq/No/M53r1w+HQlwc8fYQ0dmIk
3Xe0XeCyERpMlm3k6bLvLssuuo97gb2zeJWd/xqOBzE86uLnr4zCZIrBQK8H
uR3WxERsVHaMheBViilSGuxG8tykjYyQp894AayK5fDMn6yFX2hmUBMJJc+8
ZnmB8JQuXzAwCpmPwSFcet2IT9X7pJXmMUNQKzYNSLjXUH4qiOPJhe4xzKuK
cNrs5AT54bW+jqMj6GWbZ0y92NlKOBcGy/mZqXWQS0wqMmCqnTq6ybpj8SFE
rdoqafwYaQrzbjG4R+O4P+R7GAMzfiAisdCjB19aSBvV0GolrPgqfw8MuiHs
8kkqZwikJi4nFaJyx1ENdqVpbt8oqZSSpwYj7SXAmeevpvzgGljV3ugJOdNH
vJRdWoUDlAk24vGn82PrPc4LjDe8SJwOcZ+tARPaWNkjdrNjxegN/IRXEkhX
zHnoL/rn07VM8QQq5wbpd1cGBYROIvIGhSNhyOClwUa/uVWvC4ji6zHA19Ms
T3bm/MWXyfFih25DjBBXcKzybQWA6PUSme52xouDOkqsCgPMBmwAKL6s86cq
2WdMqzGauIgoil6pZKnnUibEbbBea07Bs1VvMbKZE2Eri5pSM+a2W7hHq74D
g9RqLeMrh10vvoNeZkc/pzFYfjONcUBm1Zp8M/PCqQAiUyg8KLKvvZmdJ6b4
kqeGEj41UA25BCAWPr4gY+59+bUlggLd1IxEywq8ZGwk2M7LNaWBfdkzk+oh
GfLmd1hc+98n2Xfr7OtrN1zhhho50tu5ph5IuCrhztJV65nfr00U5FOgJkZN
fmyYonViCRusYJCymkWV8Q968uwGpX801A2VGGgwNtHEfBAEf3JmLApgIEvN
Q7N34tBGVSrhzYR1iibBYVve6udkAWAu2RgTzMfwQ1w8KHQv6Vr9raMtj0kb
dbnPfrCXrcrT7OwVtGBjFqyRA/T622sfZnKtGvoQ4rvectcJ+Gk/3ItGwunM
IyAtfnFVlV5d7n89U/F/nznQgVFzvXcVKBiV123xcBijcHc0DmWCyyUU+fbQ
o49rlFOBUdT6N7tgAz4v7LlOIb98QwILnTmXN6hRpQQDuUrYkDoK7kUxzpTN
C0DByCTvvIw9Gxg2K4SJL7xJU5dlRWduhC/b1MHxGfhXb5671IF+DqRrHE+H
WlQO1eQT+oRsSc/QmJ/dWe8AdP6EhHL3vcQyOPRKTD64ZT3v9O1kkNEDnwDK
GzvqkvyHm/w/0WSsX55Ylhi0A0iesEz5LIWTajhSSbOzjJdUHU8xwjLArqMJ
VIq/gMQHthydOB1OmSrIpCFrWpAHec2Al9Tv8nkeE6wj0fPbUmlzGt0f79qZ
ogfibxehmGIm64nm1YgB2Il5XdUUEqyYuYy6VTbsEVKemj4VqDphHkJ4iYUs
FWmeMMMyqMiLtGg/vQ1ojCL9HL4O4mspol2JkDMleMzFmlXvhf5qBMhOGbuW
g5RvTVXY2GAK2yvJT4LhPfn3d8jQUeMzTVLK+v4gctHI6VrO1AqaPWlJOTe5
/L1/H1LQgJ8uWHTpN/wS6KtrR8uQS73asl+9Vr+QpzT6CNi1iH9YvYx5D5fV
iilvv0JcMNQP/hQk3E1VoP/qM5tvHj5WNan0O1uzpq33Yd1cd8WXkuVKeU/L
flOVGIcRSIP7Ob6VKLiMiuRnBAFTflfU/Ere457Qb3idQk33980A0tWSqlf7
ab5lDgGgC/4Rb6uZFr1aEy+qmIxeL33Xy/lQxxSzkM+S0/9Iz40us1i887lW
3NbZs9joFoZe0y3MIWpU+C8G//+z7++k76NHKwD6gQxeClPlTtxYo9E6bhCo
wRP+kcYKIGyFyMfB093PTTLaqziPmRBIvE81cYUN21k+0FTe9gxFxbcOFAMt
vZgJj1h3EbpCsrRd+huS0rIYPBPIsE0jhFYdVEeZllI1YK/k8qTUSM5Os9+S
5YiriY8geyddJIjxwdcrTGd07l4TVIHU/jThwmL92Al89dpYuTKbyV+BqOWz
Kbe/8kSUR2iOuxzphIAqai8gVbomz9i5gx04MAHLxf8wJ+M8+eQ6p8DV2j4z
Zht+26BHmMICeKti6grczpvNpLB2msZgB03V4VNH4tDTBVrBD6UyFlLmJYFu
KX8oenwChmLXHhC62SUaDh0fV/4D62HVd2zVvWnLEGPvlq0O8xKp5ngjmA7L
SJfc4hwXumzDmm6MDMIFpMC6UILtECWWgdTLDFuSHC9SNXtYlXZtSXmTUtAH
bb/nEhI/D01iihEVtIL2woXdFkHm5e9fNKSmowv826buGZwMv7+hs0AYzL3Y
bbC2Q78KjcDBt+Adnn9cwUi7BNxofN/ocXm3D+Zxq01m6QsslHrFzZzWPRad
fWSH2Tm935ppWRnl/BcCgKAoQs/MXO25D1lQ4l/IFm4g1E8Uk9hCdkhehSv2
fZnBIKcq/FwXtny0vnIiTDmV4sHYZxRH28l9s7YUYlZ7jKL4Rsyj8NMdMmhP
cHfZ1wNFlb8P0A7WFkHiyzdX4yh739jp66PmEf33j/HfVbMqIA4cri8MgvyC
WPxLAdd6/b9JlMp8EkXDMx9Y4ufCgsopA61hb0ukpMI0Jpb5+OoYLJ1EYJjo
YkGGUkXRWvWBiR/PaLwIKbxwgq/AK+o3Vr+yV/NXlQGUtXIWjeCbglc7UpnF
+NvU19UJ4u4t6RBIpzW/XesJKDzUiFNO8S9dSV7+eRnDohd1CV8QHWweQzfv
df1NMPtKRQIQDdAdkYtYFHNPhFZbMdfFqLYmxPkF5BSxxQNu5s3J6r13RsXQ
+jibsB4QlOLD0KJW393CTmwN7zYK8A26uqZ/V+J/Rqh8A/0r182EFhPTzGf6
FS+ZAev27TEDxscE3Cq/QYOyN2y4WqQJT7Hko/65tR2gNd5wl4TN4d//VLu9
AU81tbjfm7pBFzJ8Vpuc/EBCqyym8wHJi+4trDl6P9weu9Ph7ODleSQFJjOs
hqOXW580/tfszQg78i/1KuqCQ/1SAJXyAu1qgDKPEada/MFS3xHdjXemzC7A
goQaRM0ezclSYPSWdY1UTj1XGihx4yhF+zMyFB65FKMHJLr1SOLSXKVmvmYm
RNRqnYBFy3PhJMCpbqOdxj30wBDMvMktJ1iYCrsB2Uo93BAIfiPhtIzoOr3n
qjqxgFF/bLymL20qbcxB9XhdVocOQRbFyOiH88i6V7bYUejPKNaVIKUKu64G
FkdHThqu37oaPdXWRLVjubUb2J5fkkNBtU8cdS+/kSNLTgzmtA8bIh9vLDpV
uCkfrPSH9INFwe1FTYdNwKMAPeLLWw1wUWIVePBeHGwfjqBYA+xddNo77soo
prxdkGNGJFzI0QNhDQ8NgdH2puyvoT/vVcZXAVdPlY7tL6yKF8+g9uAkpSF1
+naT+J4a9QSsVqx8YkqD7BtePcmR5fEb5Upqp1QmR1M4dJffeNrzLQux0BPv
QWDzWz8TQ5WJOwk8SLkwf5bnEv+yAkT7CmPgsZSyI4wXVbLRs3ZnD2xlB/Us
medi/j9T9WiiTxLb4HqURCN2J6CI1MvbRQh+uw6X54K7OcIRrhknja7UnYep
GzTGTMUVxQe48F7R/pT5+1q94rUcJEbIT0IvKbXTBsx0a5etikCbtv9B7Z2K
8IbE1qu+5jbDlk160dwqpvezMTQ49P94w9frdwJluWqbYqXd3O5QxdU6uVqe
LMDSngeVudaqq0L71QsqpPyQKGx8bSMOT0rWWOf9dlFIT/BlNLCnNW9oQcCp
psyM9zdiXjcBcqIeGF9SQsRtmw68euWhTJHxG3QSKNpCFCEmKc+d+2kYkWG7
FKZ0PS+waZwQ6wJ8T37zQDSDGrcpXQMWcklZoD3bQUPXV0DakyPX5O2yVH2Q
aRzrV2ACQZ1IRpLbPd3ELxwTXfKh7azeIKA4/jvdGriEIEP881GVUgGQrmXZ
O4yXT9e5ixjG7ffNlHgrutdupkSXqwldG7RiDa8UBmYhcMyOmi38ADI/dwrG
GKmIl/IAEnSAc4H+KHQWx6oc4m7P59Um1uzK+doyfeVWA8pTTyi19JYYlrNC
hwHahJlZ34QX6Pl5QTFnTZ1gWLHBUpdMA6/eUfUIjHgAyL9gPFAGClzg3LlF
rutTZni3dBL208+t3ZPxn9PI2UGeOsw0fm9RYTvk9K5ox+XbUpdJqHGSJTxY
UNKk8mtkemfC1pc+aQ+eYezQ5k7IwH8uJwYC3czsvLXq5vhDXxQgaexX0KcX
WW0cdrCGq4Zb3q6ih5BH+NV021dSACQh36vx2TgJUGyHXETKDoMaTXjiTSnN
cH5DuqKWdhdRa1QU/hlIWyJyGavfkDnMCT6LIzP9Vvbvu0U7cdd534c4AEJY
i/Now/uepocP6Y4ZQ6Ofocr79jBfPKAFQbFXtEoTxw02Ikx718vr9+pLOe9G
DBrto0nUVHUfA7TNw1lb4AoMaCO+Bip7G4VNHc/ncGeGnbmN7R3qoV1uv+gI
dbSeKUq+ZK3H3zjHKM0Um9+dy4c6awRFJzdIGp6i3ke7eBX6dcIPa/z/dGRx
E1dHcfVhR0CQjgjy+tgNfACcGt6XHsX+2QhuGlUaF3zWWgtuyeUT5zji1yK4
2i71XUf2HztRCyvaKnDJLVWvompjbjgKnQaOV89zRbtZ/Gps1uUO0CqSiOuU
+Ik2Dx19N+OlkNdpdoNptwapcY7FAYsqHgIcynKX+/5/6kZPbOHFSt+Fz9Iz
8uAgkznSuS92Y+qn3tQqSVG0BO6OkD3cJP1PuKU6+iQW3v+ZRNv1oRfYufbQ
ocha3GrYBxT5Aj2NS3RMuDxlOB7ZhybRSZInjwOv9GvyyIujYWQ+10/A0EdB
88Fhb5PzIkeRTr2Hunqs9+oGDLYSvKw6nOV2HekB1b87nwilWBkPZKB/CRu0
yUYoUdHEPx66v3ZBfT78cADKvLjLgCOYDZazvr1gYGz5dFFfvxfae/VN/xaG
h7YmOvF4cFl/reKBkrKPBTB2+IXl1KUFNf/ahNmBTZywKwJWD9s/NpwRE9dF
0rZaO9wKsoF3m9rH3C8x6mUKbHHcY/dOLq5oHd4TEu3G9rlgI7QruoZDrKUw
n0PLIWyggx4WiffDphzp7JEc1pHlEzwLKSiFNeqER9gFM6BqX8Vq1SuMY905
8xamxBzyIUsqHRkLs3ZOGLYDJUSlRHktq48H1lHurqoZO+eJXKqSbO6lBRx2
LeRPmS2H2DWd2BN7Hbn/P9TxYMtZ86gISpMPDSVKDhxkx6k8mHxFJqlGAncj
lkIyNa2jpAQVG3sMJnrGRwYTH2+PrwZgnTE+/EOX2fv96dAFy98wQNyLQhlN
QCBfiHUOL3Y/Tf9FOiOdFpg8Mfm9N0P9MFzODBtskpShz24sBfjv4aFWs0M1
k2Fc+z49HJDol+NagBC3PrWadt5Mzvkl7uH3W/airGG8RIQPTBzFcDYqWa7R
2dajwRyLCAM9em9uqvOAn/KaDyCxO2+HpKvnl1a5tp65jcFMGOX5fLDppTJk
PnMwcIDJjVu7AKvTOHn10VCQ4vwxw8LJs//z/ZrbTJ0NGff4Kt/nkqdEdRLh
ULvYbLx8OvczIqDYcEJ+89i8oJ6Xpr1IKSmQ4XeazMjcpd3qSV9WJlDX3Ghx
WIJCL35BatG5VwYtOn0al7ThzBNNriQmLrjcxvSj1pOJgTfX3TGQfnN1bVKF
CLtV8tgRnwGzlUp/AiK931o7stW6JcHC7gbWR55bqwMZo90JIHxb6n7ZAQlr
dlsm0JjFmh07u/Rityo9UMaugjTLnWNRqCkMJKQE5to1FONytewAJscB/4p+
NLBNqiDqtvRrucPJyzylLL6UCRoQIL0SKdXRy8vl/sdC82SXa3ON5npAVrDm
V1FyE1wWA4lwiTdro9L5Q9gLT8LuFe7af5cuTOUDud8WPgi1YYzNq8+sL/uw
8nu1UTs62CKOhBdTG160V6ZTkHUQ2wd6sDZh2wREKDKYtNhZeRLyHntGmf3L
mfOpuSU5S/exGDRD1Vbr2IbjxqyuU7z7rvqcStCtp88fbBqDxdJfFhBi8lDG
AyfCHsKkmCYRj2qCTMlomUB4R3zDaxnscMUIOGboN/YOchnSR2xzkuDAbH0o
qRL2ZHKjJ8fVotr+IqxgRQJwA10Ovw9c2xEZXuhZ23SV+ogEleDp5sHz3OBC
saaUglOJFEsAo90CYfW82zmZlJX9Weba+bD3P/6ulW9gSFVTj1PyCS9rsrtc
wZtLW5J5pJPF7WSdWGOBPxK0gsxd2RcpKWQpTdNLHeJR1ubLdBjp0PjePY6B
6S28khF2xazpltvShBSKWp7L9wxHKIL/n/L9Ew1MmEKDoVRD2OV82AFtlBUo
IAN9PcgYqS3GvpJcrDvkE33CDWF44znaPrNPbYcfd7WgwQFw3JIGPEiXwjrc
rzi5w3KiP5dzRU87XZByRqvGxaNPPYUF6B3QVDMs5bfo3ufzGM9RpYEmAcvb
HMLrHuO7oNlqOjLa7PaDcXB+M419TP+B7H/mFQMZN00TQOJD8USGsuNFHvMk
mt1u3QH/mQg0EZBOTy9GeMSEIKB1oasPzHKh3vqbPrusEXppCN1tEPKIL+ys
HMhIk2lGCkQp/jK8MDpKPfZtqOWgZ6KE/Yb6NPtbZ2PGXPYOoLr2/yu0tvNV
w9DToZNpfdzpDI+vdOuhey9iG4WaG7xG+hwOJdWxcw5eT3Eo4vzn4xqKrtJT
a2a+h8doObV+Uqgne2Gx3r9Obu3dM7+mmuw2yZCLjwiuMmwyssN+C0sdGbVi
AFcvQyGtVfMdl4O6pQ8VIeAo3uZO/U4bj6mmf2Uq09kPtJrQQvSWBAFxF1Da
yx9qJr44WvipChpDVLgmlJaOi1cjJjkvbFIOzbuwHnAFXQgrFb5uhBlgJaR1
MSLNY6rj12tDSSSd6OtE4vLKqzcN05Bv1wvhonHAfzYZoEaE5brv5HYP+rG0
py1DvtY7gUDQqU0oySkIyLi0b2veUPENraqmd3xIhgI2GneP9R6pDKSorTie
Pp44ULd+uJfHdhD8qG065hQISDh9r4lu43+yMyOa+8MPRTw5uXQe1qBhYcKP
ulJmLaiIRBn5EgOBOyiGntBQGEAnJeA67NpC/ltNXGgo8ZX28LiUR5TVRgj9
oK30tyjH0DkJPIT1QObR88yzVcWttQVHirBmwC99QTx4SSGOVe0+NRppJLvM
tHfEme+Xc4V68mceGBJDwdyuYZkY3byE7FB4LC15NpUBRdPjbjOa29Pa4zWc
8Fi6eI7ELr4Vfjdva57bTesQPlQLP2OHhJ9i1hbwSdUEquce6y9zrT3U7/dt
4R06HXjd99eJLJJijk1PIAarJFl6cP8Cnd0TwHwDjW0wf8hsMGWL9/YawvxL
5azvN9paSiueUmR2iSOYqlylBC2BWbK22sUTWx6GalmZ9aHryFGLTB2SNxKq
UfXEm+C2OVORB/thT3UcrEYnVUc1uSQq4f/j8NuLBgl46HyL/t8xsZS3X95u
d/eBOuP5NAbtodzzdogthImznEEgBdfBwe8N1OzkqgxnBXX0mYPe22UUrwvr
riikSDJF4PA/K8T8OXwF4++tVBvHUALiePGx5xbf4loCcfRFqUJSCjn1TvVt
JuifGHepGcl3ao0AkkuP5vuxd2ahF6p+FmYYmJxfRiV/eEg2GLQfFYbj7zTM
X0NwqN6wdtTuvcSyY7muWAjzSBLjJK2OrdI/16YL8+5cs6zyZGtrsR+SI255
YSS7L9OeO1JUarh91PoXErn4RSa2DjhgumXpLSvuKxmGFozca2ebinAVqRtI
urKmUdfbHw/SdkGgQ0LObEEJfNAmj+9cCO6qAFCXVdDGYO4wBarK/+4v+qkM
RDEl7fSqRX5vnuM8er/P8Lml/Foa57NXoqjF0sv30pyPamown+nILTJsC9H+
VZEroOFwzxeoUJ2QNjUUI4ggW6GCfNVbqWZKttzmOWf/jsHyOZe6m8MkaZUB
dkLiH+l1/Pb0nds9zNGLoh1VCSKiedWISm8DZU+3hVNKclC2oYEtg0bvwOCP
RZgiEQST1KkX6GLgTa/IgcxkQeQxS+qxOknIMrS4OuxwPt4SPJV9B1O8ZJn/
K3+xMucesmHL4dkO2YtPEwnSvAdWpBKBDJkWjWoqa3HwC1BLU/b9kxqZ3oKu
pbukh3VPWyJL/hkjwj5y5d63zOc/WONOpUXK1p4b3FLRBzeZxfmbYIWCS3qY
XwBiGJw2lZ5EWwPv8h/rmMu4Ai7n3OWKCQRTnosM31e1VhC7cUMMeQzjQGA0
/IwQare7pCPgtKaUJfukg0tzgcH1gW3ZCErduAaR6su6GBx6VVrXkzuTPNBM
ryql6+xBscoXVh9YAftVIMITyRrS49b4EJvA3oik6hi5r/c2Qqf47Yx3oH2w
todSIvt5ZAGorLala2f5XKHbCROtZaljiFcUr4IfUMxKeq2vCfKgHNFwBuoy
RMA4AEi9mPBbEFDAhpkGApFCSA6xxPFW/NDVOjIswMkh+hCKdWxndmIyZRZY
3+8bR8Bjtyqln1f0/CUaezFYBxMuHqRFcu6MwcAbfxQWJreBeUJXQe4yb2Xv
f5JoLW9wvgUNLQRtcymLOha2w7bMy1YwW4i3XfTiQagQU3JjAEPJl+aE6io3
mqJJHNn3pacR9yrepfLu66DrCX/VfXe7phHZyfL23kgOBE/RmSSDaYcXnTHk
9fweURJvS7T11Le0c50+q1jKOfzDpy6qwUjdTqqdurcONwkAaWE8JW0d2mLc
XdTVQ7brzAGVZzoicns25EAEV+9+QhiAb/56CZXDuMTNqSD01gzkDlnHIKzH
LFCHe3lxnzltqunVYjWXntei/f6AteJApoZ/BGevG9bsOLR6yutIqOBDz3Sw
637RHkUNVfYCxt2X7LNHtRP60ii3+T6Gpa4KBu9HT/s1i8bK9loSHsCAk1P5
mw6sFxirRiMlB9usIKr+dUaleecth0Amc+HNjTWNfgm3675l0wGOl709KYDh
raMV93mhGsfzEyQgVJlUgxUTLBa7qSeOMMyBdYpbQY8ZOkigE3ZhVAgo75U9
FzvXCZTe7zNUXQkXK/b1uBm2MiFf0TQ9bMAUrFupfdhyNYKlB7jRStvs116x
LNQCItTkCSyC5EHLnT7QttXeiAETYEC5Cxwcd+BVlimRhDvl0Iqj0gPo55Xo
kKY8NwLx8/7BeKnFNTVd5ZlHSqduMXdTsrqmmKpH2MmbCRJK9fOL1s894v+w
36UuY0wRD2vmILv4yK/okG2jzYs2evpofXsIDwQGnxhd9nWwhtCIi+RKyt72
LXMT4BqH2ivAHHyVvNof1L1NyUdvMOzUd5BYPPVOnOUi8OKu3amF5XZ6etmm
EpoK2iWrSaj7STJiQsJ642AMCauOHPabR2hNHvGGAUN2g2enoFqpKJYdNW9c
Ni3SQrIH0EsT+Fkhy3xkd7D2+A5C+ux43I4njOa1a+7vuXEN0txIYE22p4ra
LbRZZItngjFXw6EkhzY+FmL0+8USp1FgFXFNojlVGVvW4sjjCx3G7TeIbsQc
4ITe8Kq3nk+U7NCHw219GAn6PI2m6I6xtigNmM89wdsEJ4ygPfTqceJ7yBKz
w1WBPmrxrNH8r0OQNNyBAniwx1PPvOQW8F+umHeV4kVBnpcAW1svw1/mS8tD
/a76X06OTHxVJaAcGXi3wgKvBgqFY4faXYYY52ZvbXAYujI+oQw8vwZg2WFp
/j+WHsb5f0RpuPnXiZeFI76Dg4nTTztp74cxgqlgydJ0ij6RkwHLMkd5C56T
4UemTvNkQLfyLPcbv/mZCMopg98OSIzuVZu+q0DYyeI1n9iyUGKe+lZ0gWe3
Z/LdYBQ00IVsWLCj9vb9HzQNaSgra5KvO512vGjjrU7itQ6+3ovlodeqBpRN
uux5MMR64YIJmPuOp7IR331P6NYfGBg2ko7Tm9mVQilvHMxgkjec6FG702hM
dy8wRnNqq6r80ME5W6APVHBpTdLqLyj31WCvEU3ZSMyjbGO0/5Hs/Op2QWpQ
iCWsy2+EfPCldYySS3Nh2REbt0foUfM9A+Ura1H9Y+w9BA4n+SlRCQUd/cnl
+sh+/PUP6mlvQ03ng91N1d97cYpo8Lu0XlwH/1sp5ZTRi5TdryeyGE1VOXq5
PR9DhSlZ9iOGTdlyT+eHsk+LZoV0aQoSIUmQnersw+Qd8OM5M6OJGwmIOeu3
k0UK7B9JpcFAd4GOEqvZXBN6H5CJeVd1VyeDbelys89vGVvxcAuPj/1Lt0Ah
jq7IbNCKGI/IGltdljRxcK/5AY9U1XVa5USfAJjaAO7nuY7NmeOJmzfWUNhF
eHfI3VlE+MKgZo4e7KQxp7H4owjkFGiHSPdubKxr9JaxeRbSBkn/2hp4+QAL
IDfoyPyc7S1bcxkpFBtuzrpBeUWx7PxJOu2hIHtpaV8tzkdfg3piF5D+Btw2
kfmlppnQPyqrVPXdwM29kd+7lPFc2zpxWKO/TWPEy1Iuk3aWprvUi5x+9bsS
xwho/n3TEu+7ahr0inyvKgtZJLb2NESZuEwyVM+MaO9JPVFPhIAntddDhSfV
y44B+IYIwF/gQIwmXWcj0TF27ElOMb7etAGmM4bQrX1sAFE9IyLpgtXOMLe4
Vt86Gq9DVYxWUsSIjfZuxx9OvidaX23reTVTeh7qnISYF/DXlvVnSqfFZ+VX
oIx5qt1HUiKaekH2NCe+M1Hr6sj07AtQxzolQEmm80Slyu8N7yLus/tD2kgQ
IZyEFWTyyB3rwotB6QB21wYBHXhFtkI/UTUkjWUxMdyiQE4ff+jN+tK/WkAd
/InBwadCCQaax0U113v4Ppg/qPS0c9y+e3zDc+zSV7cDmNcoKuYEbXgOBi3g
neZnt1lcCRITC8TbTKqKHf5Nfz3it1zT6zlrjCDH6dyJjycPKkCrnOUX/TaW
36KHxcL273tyPjwwXAfrp0cCAwcquWQTQzMWEstUq+VAd0ya5n3BYwH8oGFm
gtR1nFDgZ/+GaYvdGgsFgZkVwOzGV3vUXcmYu+1nHuLWhtBYYyC77jziiKlO
7HxAeAFkwUOEG2YPR/OgPVi9R4kBE9MCNR46GPlilae2pbURpJPabGRfiH/p
NnnTTWA5GvH6xQNQ9UlH8ecPAimq8NFgRIDTcIWW6riI9CZIt7Wt6+IhNsAi
xLJD6rmkCFhFF7gGSzeM3kA3dhWWWRF/6wcHCknadCqJO6NapqjiyrU2vxek
SeeETpwIrD6uBBuF4ATOtZ0VmiPZDA03Mtd4OJjwsj1bOgWXBBqh1F9accAe
tviZZacfXL1ohhPKWDQW99AOzrYDkKzPvKKKYhNg57HizWsDrBJD0CZDH0Rv
oMAMMpiz7aBtKMlJQWMYNXujUQ5bg76n9jtCcf44K9KyT0K+ULjs6TQHBJaz
4m6pWF32yduJfYY1L6aWlp2xkWKQAeB8OLqiu3xBH1F3nHDQxJplFIsieD7j
PcGSy4T9ND+6vlX3Ox3iX/J3CW3EQIJehUVgGSuSiDB3gqy3jZSSPJORJE7H
8JCzA8KMwUKpIXZdHEJRuTfd0F923jBfMvHNSMv9OBb3e7yhE4RtiXRr8LuD
k7t160B99/7sZOTYpgAFV4FQesdGM1Bo0mDHaLUi+3C1gFYuoHfm7QzRgX3P
IXhSgybxOhNg0h3M0JM7UDSptOiat13yYkOXUfUvL+XTPDU3le6jRSdHoSuP
iUIUiKGMvsJnhHpnnnKYhAkcIs4IpuxhCpeUk5OwomEERell9ZQ6Zotf8y44
9OuqKbYP+Y2Gz8XCEtwoDF/zbZHMlrQF15QNmBsm2z+r0ZIyzQ210pI6brPA
/HrMiHaHeJYRaa0kn4HEIaQs+2pu8wdXGNvELelTvcf0iaywBV2h7uIrMTkm
oFKw9vXRWoC69BWcnILFIkb2YZF7Y4xn396lZvGujBPvZqdtFlrbBLrMeSOp
3aBhRQNtYswoGan08AMDYLmlpS0UQrTr9aVGCALQCakR8wL5e6dcyRiuSadS
AGTYTSAAohI17xpYh8TRl4vk6eGr/AnRU4pit1hKQuzh6aduTfVvJuiEGRx6
qSk2MjQ2QoKnvOsWFaKDV169s9xPJ8CKs7tjbMDqka0ks2HshTedWDLyhP9k
DwvqddCC4lEQbXNlHcL5C2sq+v1pl3v+HjVmpmY8Kd9znVw2XcVoZCGS7N1Q
EpUaQQOMaN//Zh/I788C85oJHz5/yajbiDMdIYSZemZKEoP0rQpwCRtp5YqJ
P0+7HEHJQW36gqRQPdSLPd5FBFdWqhbVf+aYhD1vimdRckYMypfcfVe6hSuT
sa7Wbht9RGLsHY+FG/nWLTfIxBY2EwnvCG+L+bM4WhN1/4ttkKcOqkolAQHS
bA1qZzWWSXxLJ9gDaX2ELvK94sWx/TFJhJjdLIpLdwEAluRrJG60jHGeeaEl
hma525DwmTG/RL6V3kjBZp72PmCJvcwdpGV19u6+UjgFrISCMj+2tAndKmtT
4IYvmvWghlYIhrt1gP/E3Wp+gEDRdxyR/AGiDqm8XwlkFXacuFsI6MnVaiWw
2BDZIVlZydtVmMs0PmIGY1qkBYoucJ142XCLk1lW7XQJdwuZ+/e+0wIXqsOW
YKhXfr+tG43aL0jL9xPLf+gYbi3q/uIc8zZs5+ecXf6bFIVUBoltb3c0qKN3
9lDUaNKn1kgEUQBQsZIsb1TQkAslGOZ/oruhSvAZYOCsUAF8cQVK2Lie4Sw3
rce4FEoweG4utORHn+HA4Udw4y/IcdoyPTqILhQP9UTikSZAx0JQnLAeeCFt
7hFhN7vWd6owzCFMPTTWnX/+3GquqDQmMFCl+5emrfMhbMmyH8W8y4sSj/Ka
YfzcG9UCAo4dsGJGVW5RbOeK6h/HiLu1EHwzHC0Tvxj8ToWV2fIxMJ0v8ZpX
WoHoA8r/L8gbWWnixtsUl1Krsb+2mfo4ILbGaDAPe+amkY+cEWr1zXLMrSaL
7tPWdcCKLfPOxsZ18IU93nHQrjuRvaLmfA6IqLtRXlxMNeRn7TCHHMDE+4ik
FggdWM91eTpBb2p91rwGxLJ9RSbDBomx/Rh17Sy28ejWkb/7p7vu+YYRTDKU
teLyCYjEoyE49su0XR0CTIm6VAL8viNobQRBzGJqa/p+buhfTBAv6ss6QQl+
06zDH6zVSzcN5hJBWegbb+2oTvcthsUQpT0TBZcknh560hzg8tsuIDqlIwE/
LtphcwsfdEkKpvVKiYuychV2nDIqnFkUWioBWwMgBt1JBToVvS5y9vR9otUb
jhjzko6TaW1YJVyeeqTJnkKj0OS2uV31INYpVTRUu/uWiJrUM3CfqZK5TJU5
TkJXfAhmFZM4H97lE5jzvVyaEgYXaG+0yf4+CSgHcYA6z9TARQB4Cd8RaA9F
xxz5xsn2+HndqvZlwYsM7uX/uuRORh+NM7OU8XLcP2KoIRLqrrtnGLsJR07v
I6pxLt97hBqfm0TTh6dTdkeggr7KlTB7kFosA1H1RRm7T35DiwZ7h1gULkMn
M4QBfuhv5vjJnfAypFUYCsrchqTLwmTQ9vQKEKxBmRs3amr6t9c9AwsKVxna
Etr/5X7D1/bFRMRu2chept4aa11NMPldisfWsCssirI0OAiS88ivAz6MG3+Z
PZpHnYNowz5+hBmwHQzbt9X6an7tmzXpC2QG2wJBTy8fOqY68GutvbDB+7Ps
9dfOBJwhPj9m0h5/kKK3MsLQUuXfKF0yvji1/S/Bni9n8oV6WJkx5KwlxG0G
OGVd66WarBOXfvDQKs322H+xYcs6YtzGxXcHKKe7arsg/EpdwAbJLuc/fhE2
MOaLTM1oraLPcOZ+lVze+PbukwrhQaAVOY0OqJVGPohDh2tG1lFuQqz81Q03
nnQffxea2P9FbMuIiQ+nyh3cBBxqA9I82wwpHxl9hXqsfo6KYn6XVVlcRXbg
zlesE0drSckmdxcN2B4Qkr+/AeDFGrKxfX4/ccn5XYwObxxjoFTqgbGUFmx4
KghU3TJcG0g/pUfotqIHGYqh3ExFxqlhBp+D7TBtXOTOdOPPO1Fn9jpXu7Yr
maDxkgeMS+zNyK7OsWGFCwmjHTmjmQmwaVooqhfrTsbvp02ykHFnKsXk7UuG
PcPFIAgrtvLVWTXVBJTxaFW4z6GoILMsW8DpxF8mgZfqSkvCYTN6InUWBkeN
Gkln4egSepmfYGrhjR79J3lnYUCy69lIQBsKu8N3Vq0egd9J4dxuQRBgXSEH
NJSrGiBVTYOg4JD6heTg0kDbAswCyD139GEcBcvpFOtyyehvJKjBiNVcvphM
9NxsAOYDiw6Ky0maRjwM/ccMMoFnwo0s3jt/XGp21HDmDKrH2fR+EJeE1bC+
J6xJFWwsQDrJrntFS4Uue1LFc7cgE20OSqOXXRzrbVWCZr9W6R7ymQwcwYIo
uOfLA3q5VaAQHifyUD8CQLvE4iIX4UEvsYwvXjKI3AroLtmcE15sHOyHMBZA
42Nu6fy37Hhg9K2EDyRkg+e8lpoSney3faEb6n6qruwoWF2Y6Tr5Hmb5dWGI
/ikLtnjlSg==

`pragma protect end_protected
