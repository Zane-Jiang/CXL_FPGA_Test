// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
gbmxj5YQLFkKqOWkGGmcBvDxshakZH8kXKXcwN2xAKF1XsTZWrRf/Ubnq7HzOmteIC2ensF92Hsg
U106OGKooHJGtz0jXARFKTi7+xtxwV2HUlAYkhyZ4/6wIjV28mn5RPTbZKFDAUJNFSqgoLzF11PM
cv4HEJn+BZfNczUKP8XmLWE7dpK8yviNLmSV/+ZPC4/zthHzshdhk46bll/JVKetLewe/CoRxYGE
oDKa14Fs1PxLjOv6CXBLVLd5//QDQM4Lr+gUT+BX1Ba5PRuJDfIV4De7DhqbOLSOOkMjl1vpJwEq
7Hse/155L/TiwIZ1KXR3/gDzTDKMoZgave6UvA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22160)
/fJhaO8mYWLrkHFQQlfn7IBy35SiG8p0Sda/1ZwsWs6QZDCQ1hGZMfZuIsVy6cSh9jvqPkq76RM5
V+QRNVK0Y4iPppCbMWX0vueT0+oJapKz8/p/DFoKWRtqsPILZX3auwl6EWfuoPLx2TTedK/E14fQ
aVGM2MXXPQGVWD2+6nkZP20sfb92u48iT/RwOZworcEFgmzsuY7omh7d+yM0k28lJ9UGIemLVJ4Q
F2FDusa25Bi51rDhTEMJL5nEMwPYvBw+fsfzjLiDAsYNywFwRYU4bbEOOcdqjlts068/MovgQLHo
uZRWQ31QVg86jhhiOxjQu2wdpNkOiEraA9ZveLvZbPQ0mdid4sF4x65/NZ/tA9xr++2jHo9Z1tmN
Mf9hjL1rNboA/n51jJ+vDlkRxvIzBcvyQrt3pcjdcD8C+DHbUKS81smwYkhxKzK79zWawqTp+KYF
FE+8wTuj6pBYu/55ofvdPlcunIERrHcwwZTzuKMXH0gdRk+HID5NxsWSUCc+K5dhHxVLPdTy88X/
AUvN4XJSFBKK5pxcbzxrM8qATpedN21Vt+rDPZ937ep+VqXKBdWsalgmOP4AAtZRl9dXwR/8P44/
stHdx/lZ7vsJn200K7VaOjcvTfss2ATjRC2ihq2lCDkk694fBZUdtX1ThEGGXqLxlbfY4K44JDio
7YKwQ0v/S/dJgByLammXjBK+p/VzpXspZJwGqCf1JOr/BWn+Jy5nEsr8fXK2eGnUoKdvG6tyU+J3
JhtHSByjY+fFfuUmAtpK9EWVg5B95UTG1PI9JYX4Qeb6NdpmJB+N1Z1ZjCuhRuGaSX4XXnkyCSBb
SBvEsLJz+UrbplK0WjKTtIvu0pUORBIyINJpFu+vx1Z+idWLLabziQCsBlDekEp8T0ZeD+zAX3UH
eBRDA9eetfAXn6QsyX8VOWjdceiT6vAr7xMigHwF0jLXQa4fJa00GqXCRJc9fSaFV9QMg9KLCPcV
YBBar9uBILft/tbA0aYZBva7vv9rU86ZqU2vcMJMFQKh5hMiwPsra/7mJZSudX8sDRVOFb8DeloT
R3qvbVVJT39Ua2KxsNlGTo8lsHDJbBY/wyyKcFfpdvtbLPnrpj962hasA0Pxp73jSrLaOaMhbjve
ZjJlfEJne8fGDjLLNzXiMJdCAvxp+0ufSvuCHeafNZs8v2c2Kk/AKjBgjGSCkykESqbdPJVdhVCE
De53enhr+BAOQQW/dq8tZyxoiDxJcl+HQl+XKmkuTD9zJ/44e4ouhc1Vp7koU7NFwHg06k8lkJdo
KjuD9MfiTxGSsikHEZOq10XvtjIVPEKqjdytDK7g6y4jehJOPuY/OtKurORRt7Wya1nIqxh35RBc
naIzbgz+Oq8M6oJ2rmeXuhTc4FQiouB1wjcMw/EPT+09TQxExiukooSd89Hn61zCScOnkUvGQFQK
YMzoRe6b3/doPZP7JGxuxtvMjUMkfjzei4bf3bO1Q7B+gaFOhKXwfvzeREdKLmUKG0WjinpmbO4g
dhLDV6X9BJgdyW2hTyzc/DpjgDH3rkdx3iWmxwxPrPBYdLVR2lTZvylGOlQ0J655lpSmFjXw689O
fBg8eAFe6OOeaSHZ6JDXAuLQtHUjvYmrIqLrl6Uxlmvf7Wd9ck0tokHaNtz4lrledCaf9ij0qbwr
/F7pB33Cg2MJuyfWxoHX4VpFh27OJEyIygv3ZwXV3ul3Zl46b3ExAh/j7EoP2FJNafEEFNCyE2DR
OIiW6kk0F78n/JNLo2lelxa4h0iwZ+eertrpCLWfQdCUywUE+aTiCTUAfX681qdpdfiiicVLziCl
GTK6cpV3CzIRKgb1LQXN81/u1wP0JwdvZpKOD0RnS0nMWWfSVqyEXJ/p4pel4kQAwxCo03BnLZwV
NmaIeYDLwJm9lUqcdEl8AJy96Kon4rzG4e5+FqjiofyL/Ib++5DOKlJj5aa2YPGpch9JCvHzaZYo
U/RDAEut7T6n1epf3olJMDMR1imHXlfd22O3YW58RlWNXRTg/f9xgc1rTmYr4tLJDxlk8bVMONOW
92Lkz92XULRbw9q3/rFyfxTsFIWxfKYPekqP528RB/xksKNTPUkRqsqpfU4FOaELVLVMQ5Ta+Cv4
wwyDpY8u9TGGJVejbflb/9OLzJqyHR3stONNTPexKfLIOtV3A9K2cmYPCNMb+GtzjdwmRM9LALI3
fcfRO6qTfcPXEs7jZ7+K79Rmy5zn92lttR2kSA48bxvjPPo9e1sFqNLjfqCRqlBHWUrFjlgvLVDh
0+kSVlZA0RVy9R54pFRdgEAyIVNhZsiyVcexj5fk6rih5u5h09MsuR+GL1vxsiY+jK0t7zW+eCg9
w5yUEoXQV+SGhmOF14Ry/WXP9GQZ/euanm7dx+I7zPhUIWO0ZJC1GFMfdXwZLs9O0NkD17K8/3y4
avLHPcmRY2FfqlHF/2yVWxTf/Hy2XiiuysqdXsvzB+TIwsTIgtM5wvzTDdk6aL3rNOGWzGpGb1cI
MIFj2ikEdlwxu1q7YEd/3goZus+WtkSIwULcscmDIwurH8rEvJhAmk2zttLO6DGM7m131iyFqawg
2aDtewGOiM2gzKmyRILqxR2j3V+rSyPYRiKOhMybr0UgxaJlRbYvlebV/9BMmLDJZKiBP9Cc2aQu
0sKjlAItwtSCaU3xWZYEWiKW2X0qFNAnnt5GroeWXT/FqW/4010uDi0qISmGCFJEVxpVKtwF5Eq0
2inxZAKGVH95HaRB9M1x337FUKWLM+3lWgKIaYpiiNax6dDDVzx7aXRa5KtaZdjznDuxt0sxiUIj
vyDZKEzjquRW3Qbnx+/X+En8XLdTx9HVN8JvexqJnSliriy48B/DFiks5EXKwAxIMBNmrC3dry/T
IVjmijAJv3jFzNK0qVbxHMSQ/NCcnvmqQG1vIW7nxWbCESPsSmewl72urfHGvQqO/XwEqiKe/1XU
uDeViu5XGEPIUN9FYCZX4G74LKHL46WxPlxqF60HpXxA6fUCr3vZuJIrEn1i2Rfau14jJFD1i/+b
xnvZ88ltsGvH165tnbsuc2fa9cOH2pqGLO/d68bgBbD/Aa1Nuz9wbboX735tZCQ8pMjSSHD+ohFi
TzcBSw0SE6iQIK3pgxlK7bZxY10+DGCQDqepJJJNL7eWtyDUTHqplbZ2UA7jcaW+zO9EIipmPwwn
zqHLBXOb4nrhjgjpBNhs1eyPXFGIgk3MlUZ6qy0hRPZELVLU3Hchr7l4E/m5Qr+jZcDy56bnzjnl
MHO/7klrzBkB4G9qKGUOjuzYeS5piTxklLnu7/RTTH7hSyJeLXJRS/D+9i7KsU8Gm9RMp8kLKyP0
xY3iO0PmotiZJjj9gJzqxty6bpT5h6rqqFX4AIanHXOzLjgvitHPTSySghzxklrEzbaYs/eEj3OU
091uMQwdtj/I+evamgUybUVIzbN6cdQl90bZmxlqdMNk2pitnf5cze1jY1yWvlx3IO9LYEcGvzoB
dIPvYtFJJatY0Z2sM/ApIYSmP5JVlCLMYdPHNV0thPqRRNHQkbNn3YLwvz+NtdIgaupkqw1ks3oN
WBbuiKBAkxLBhkiRr4kTniCO9Kz73+yFiakpFLWN/SmGXOHCAlcAxziNtxrD4CGxhY3ffgXemwOf
2zi0BQgAPpDv8OFW+XZBH41ID4pyrghlf53ZZsMj1aD5qp2vdhcRIuSXjWSNwNFaGTAtsTkqt31z
8vsUT/qZKGRlPzeePowYEg63yrj5V/dFz4GX/MgdxfxFU2Rwtn1KSEf5mpMJ45AN1BHiPMsoDiv/
OcSRQOvB/l0dVX3DtSBPOuodG9SIOX57ngvsknp01W7B0GkDMXSgMuypnF5C9DlJZ4iFpLYzM4VA
26JBRAESjGFtDxFC33FhcsjiLivABh5H882pFVfnXFnNO2Vo/wDer9Z/B6MJYw/NAk09TceYjNXY
8Z/Copxok//DSP6WxTkUYlDKHSreimDpXFoulPXOobS813ChRcxnP4mJDDTyoW0t3lpZYX37LwbN
K8a6ZOuqM7d/8eHOExvUFeGApviGz+jNXdQmgCIa+OaVSfVcBHIGffHMCCEUjeDgld3DYqMg8+0R
Qu28XRiyevBd5JPNwNdVdlsdeNWxqkCRkOj6uIJ/uNV3OdizTn2YBGHh9lZV8PkbBMLBGZUi2OaF
RS7XpFF892KO/Smk0xDk3G8hJGhsshgrku+oKcovjqjF7d63RtHK8krO4NB4GZMkl+uhjDzqO45f
j2UEXVIqFRuNttppYGDT0MXlt8c9XI/LfbgeEsFA8vt6vPOoHB6nwE4WwpdJ1mFjVLv0LJuHa4yS
n/Cb0dMC1Nu8t0YQGTOkafk0jRtkf6CSh1ZimMKq0GZlhKBzGBMEOkEcwusWf2CJhYx6v5GZCX0j
4SwKjbKsYk6rUaD9T01VVSbZaTlF/6EdoiGmB3gUkqjp8k5ICqf+aKxhxs5HnlFeL5HVGwP27WZh
i8P5HkhKFsLjjrC/xDP6qZI9u7HhAqnI7rHRUNdfYsKTT4bWN0z3fNOUeRFtkJN9rEjZTAnfRAWT
Y9Pl/mFzAODW9r9bK6DtYZObsv+UUnkKZA/QubT1JyBWpkqXJUzEU9VPmwzxr9g8Q10w6NSJi7RY
kWCemeJVqx3Kc6I4d7ffEC5sqDVEpI6HtIewM5rmJT/19br07drX0j2jSjYGf6kQ13T+D1tLqIzS
rnH9wis8OI+WsgQVeoMo1UTooZ+HmegWYmfIS8c4hkq9XgW3oMVlwPBmv2eU/lUW7/GJG+moKWbu
hqQvFsv+azH0ZOl3HY1TGqXH5m1Et8yyev5nYa+Gl0eN27He/iyorcccAWRjqrKPP1YTH6QJQBNw
tG7tRuCEI1YZWiU/7CbG4N9SJbfYiqnKYefhcLv40UvxCcH72CGPffjq8KI5xJQl92ASXrUuNzB/
wI3OO7KZDhbUaAlqy62zE8Ixsw3hrbckMoIv9TfvemngkvJAmEQMGfqHLyP5hhEzZgYZrfLac4KI
YI2nnyPolb54pu+G2brtBZ2FI2PCY4a+RAX+Jkt37MHOXLZ4/kBno5CoUPeoTsU/ZjEfpzXrT7NZ
W3Prel9ldDCpqgqCAz5bJGHAbMQAMZxSxGZt9lxkxd/R9Iqx0iWTHmeaLIgcvEtNwKLE0N8/EA9s
MnRQDb/AcI3FTzPi2qWSmvl6VMmXtj/3KFgjpoqhK+JIaSRVQUemyiXJ2l+BRPbkViTp75QKNJoE
zgx59lHG4cuPzM8kza+8K7ZibpzpXQye+a4yH8rTDwVbwL3l1yBOH2JDUaVo2V/Wnz3sFKdcw7Pi
QCgY9tJva7/e3W8fy27PQlwlUFkgsFr7n9NZ8shnQVmxHa6of/Vx6SIplyj+DX1ChYrbiVQu7WCx
/f+G30R70BElnPdNuJ62dR/7M0l0Q+WK+XsaiXKlImDHwEU+L04riX1/UI33pRQcBvJCXv4zYYRB
TR/NU7TLWdor04bGLkOPTC7MCCKfinOI5aTWSun+HO8O4qShEm9pGCvOXoZXSeSODf7KPsERkSYP
k01LvFVxZaMZAsgQisNiZRqkDMTKCYMg+rsy6iPKlb/2fKh+v/w8M2uDKts/swvkN0nnwIoqvGkP
cHN8+/vg+iqTnhs1jO+vuzynl7iLt/lv298FpiCfvUI8Y6jF5JKT8rv19H6L72GSRXiepA80sZ5C
XhBdJdXlFTvSGZRVWacM37AXfqG8Zcsjg+fa6ni/E2zTQtvyHFUJBMvBWV0nsPABxkknjedkxiDw
7MGiqS92fSiMsxQKTK+gFSDE362b+Jm1Mnj+0Hh7qr4YVkr0u94Ra4m9o+LqOBLmiBXa/t8SQ5Us
Nx6KaD+f/X2hz4cewu7qDUP49ZGqYPaVh+Py9VW3RIabE5zy2L+HrVyLBWmoy5vuCo6cfl49jnOE
NYc5yV4jP1EB4RhZME/iop+CLPiqCjqgInisr1VZ/FrV2QfdMrdkxSKgYK/uAca7Y5AoKUPfYsAO
AWlDkU7ovQmSvLTOcUp7Re0sD6zzvlT2+YMSZcrdMkMISybipgqbSBkr9pWaD080UOos9YHKvLH0
BgVgiLSCTU+ZBdh6LpPqvwbVWmeb/UXqaiaZzAjqlJC4LX3VVcV2f8hJa3dIWF124Wx/v2hlUZRD
p/nNazf/GvvtZSF/gReugKXFTsC5Dz9d9LXfIFq7xNVoLw+hmn/RZ/dLGO0u7MmWjdb9FE0tujXZ
VMyKUz5Upb1RZsIIbhaUV1rbI385No3EISK8hTlbsZWc5omJqOjLYyMEsHB9tqQJ8zp4uzfWBfru
7ettE/quxuOt4JcBg41zXl2CxX411WK0170ULLbihHFszGpwIIocW5Aa2VQ8PH6/2BmqC88oLuIt
fU88y4IpYibxzdC342A/p5We5zy7miBwQjAXflbGo//zeWe6R8XJGx8gY/uVPxvxQA/bXPsupYCc
M28ouQv75hMVoAxqOGrr/BoTYuiccZkO8jjuy9ZP7iqMz3DBgiCYFYUwsqvHq0D8Z0usXorRJpeC
Altx0w2npO+keNzHJ9JixkJqGFwPCxgY1u97qrTE9oScUSW1Z0DWT8333tZpFhmjPsWcejke4dpV
/udDkniU5N8QLkYDizobtli1vRGmutCeq0qsbg+iiVBwa/OZYb9YX3VsplKgkyn9kMV5JdOMKsbo
q9AuAJZF99VjxXU83GYzTCMbVnyu2BsPmR349o146Q9PAhH2CrnUIjh6jsW3yPbnpORk6BuQNwSq
/SnHk0YDpEhbfS51u0LTLVJB15L9M8Jttxr6INvrDHPPIuPpZtMM3KP2Q9CeA9v1JDiUn2su75Ma
/EsvVrF3HUTgHLbvdnbXXpNy9TOaeayMDbtB0B2g/btW2+dl1STWLQJta8aa72B2sTchB1Ary34E
SWL3krH3SeNj0wooW1QwGRibsryR6gnhIVY/eRl+4+A3jJF30WCLTmjDXqv617XhmzSdfIdiVhwi
kgQroSYgBgqZos/mOTdLObuQP1gDNbZvsTaDcYwBdGJvvMM72MQ9ty4C0080zfd5L5dPhC5WjXQ/
TR+nf8m0ysiuubCGz85UY7QUwhdQmKKzhVjmL2jMuAYBBdVTH8aQIntTZriPbBf45TaYKrTjfYac
gyIBAjDDaC7yNgu/eUUDSj96csFM0C44XbYRUsgVV3jaHU7JcCw57/l62qTs3Z+Bi4W86GI1BGCP
oVf5cg1mafbnIrimcBFecfykuxgPvh/rKELQEZaNyXCRbNXmWQIOBQHKp9Lut4ZFuKCiw3aoTDfd
RaaTUX82mJDknbi03vWLv+SF2nkvOPmDx9ug1UaPaQhxTLOiCfePWIZpKAUNpnHSp+uSSKmowPuK
8zQE3fJYC2jm0zWqRzcFEf5fcI6RE3oyyQViqS86sn0jhxk5nyzDiZ7S4t3wW82qNDmRR/77gMzl
fpA5m4EP7lu7wBAri+eEZDZczp/cJLJaKFmII/Ha8A+YNW/eVJespG26JTZlYBVVJbpQDREC9mvK
eeJ+zNTr0lw9vhKTM5setstPIAMKhlDxBwizzHtdHI7dF5WSPkRriKbzJg6okLaFSvpWhdyWW937
mvY5+3W/PTdNvv9/70ECvdu6tPy6VipyFaTqud4B2iYKOLpZ6FOmeXkYifoYNfhoTWzJfgvqz7z2
jGLW3+lcNBjpcryftT3sSz3yUbVUSmgYJNjgdRoHq3IDNl+T8PyNOl4S5oYmUBQ/Fih1VoilRJ/3
aJrttQDe7dhBmEduSF5Z0cd+/aEuhpWrT0YfXMC5n1lAWI+CVWMMD6Wfk0XGsImOUUng8/7lsNY8
YeesEwVXgZ4xNkR555Omq+Ny9+ZIIP1gFzte4ISnMmznYCQ6Zjylvy8bqKg7qd9cWPrN7z9Go9Ei
FzSYmOcnfd/yWEagsOeQiMCb9uFcqdlVPLAzCyMcWhOP7A9/DlP6mslZdc6/UHHsudCYj8yWlpwi
+IUGgOUOHxjTcxDUI9on8ZgjG+UOUmsauE5ZxUaXODcyDY5KmOXNtQ346ef+4lqikcbM5GoMIr7K
kYX17O5f8gzBTIkQ/Pw1kuxxZCLvwY8KFYH4KKW22JI84JD7v9X8vVC/DeHRUwZeSLTeXJru5evi
uHsHaFhrzA7V3pEyi48lHYR5DY4cdGOF3hnqPTAW+QPmYCkuO75rxByvG+BY0463KEC4po+rh71c
oO9CeEkz9HZGXYpuEs+Z+Ih8arEqIbG9nlqURTGKMpZgxR9P2NK6wr58znTnmhNqt1Ok2H4E1OhH
K5Ip0Rax79Ynjr0/S8eoy182a1T/M1jRC6+ImimF1jTSRMqTQ/wF/9HeTRfgVPp9jvu3jGVh40fg
eEw/55cDb/DVR1q/Lik4evtF5SvWnkU1Vui5mOon5iiukMR0MjraJzzTPPPHIxiQx2eGHPf6fzrN
wwzqF3w1dmwKUeGXhHjdBfh9czKUaKsTNHzSt/zvsBbCqd0D9Oh+btCCdqKU2D5Vx0F1CIuVKyoo
l2umt/oJZacMM4s40HcL7Pgvv/mL49/YLpIRzPaRVktsTYRk/xP/7fWiUWAVaPD2KCkMTVmOSFlS
+mnuapbQzMTkEPnTyftuu9GZN29zl3fOg37B94ygupcxCUD/dASs3RP+JVR2RzhJdSQaC5g5mWMA
rbv7NXDChJxKDtyPviYrQ0XX17y2KMrzFzqGXtMHoe8x9g+MON8vxMavDOg4SStE2d4Ep5HOPegD
HUk/UNDs/hjab6q0suSeKv93aPC/JPg9zZbvzdCFFOREWpg9rSWbCbc4gQbQL9jaUtth6eKRqLod
Ec8lMeQkZ5Dt1KEMOU27dJRFZA5RqmSqdOLydthGsxPWk39PYOAOcadf6UxE0qy7C6KrIoWEtiJW
dTRsoWSezXx5yrDbTulfTZ9680UW8Z7057/7GbKIB1SGi0bqXnkf7nVSQnfeMIiYpt3bmbXu7Thb
fV5XBwanhGp8Rv2B1uw8jWdonqa54yZ0tH9f+2UHp4hadvcSYXSAUwrWbQfjwOVBOaf7x8Prwtdd
bK2O1iGM4ispoCE9nlKVPVM/q4oeq2PRnQpyNF5+ATHC7f5wM1J/Ua1fkg0NC73JxbORADYk1s2+
Q/UZR1Mmysgzjbvpn0p89VFIvwzBJ3VdrBdh2Mg7RiyngGahkJFda63p6J6FaWQwEATMXn0Zs479
eC9GKjAuAJ5S4bHRJjCj1DpV+mr7xwuSVu2TA+ar2MMfwllxXzo3FUgcsbfWY7D8Ld5FEKMZ/0Ce
BG3Un8oLth2iYuJTU63QaZhe5yUvzWF/hj5L59xQqvpLGgao1R5oFMxDUlDU7isxD4mo+z8YI13Q
BP9yWk6QpRbhIZ1y7Fo84I0/zLHgTlZwgKrMZIo/xezYK+Y5hAyBRF51+9JXl65cP3BZnzcrSDxn
iYFR1XLsYfNjxwqaFcctMFeuzxhM3k9pXjI900q/Pzj2v0+zNCsCktFdP1sz3ONHD6g/8YLwImlm
sAlWGsAymsdK9p8s4CrgFeKtm32Brjxl9GxllZO79bwa6Py7hOKAhiyP8SUuHT26oGDc/kuOsd6A
1GRJf2lM262PpLHN3DkM80zsxJ0ev2BBwhXxMmKcZR6wa+sPniko6Y3p5o0fjxIOdv6CaaKOav5U
TffMFn0kGpb+YfKXAyZuPhot5UoriNyuF0WSUPk1A4qo6Y33+MiaIAs8HK2kB7MzsevlEkKJn7Mq
kHIzAlhCh1f+bXxzRD08fzuyXQF9Dzlh557dqHnZ67MM0vDIkbVsIaeKWvWZn9iUfqljA1i1uhjJ
kOZpyzfTCodHH+n6fPfT7t7Q8R9jAuWHkUlT6GZAEi7RaXFh1yiT5HEMevFw1X7S7ZdoCKn1od0E
JNZuCD29HtC9K9dfk+9oEJwjPUb4evlZUi0G6w39IXB9FPEvaIy7niaJ9SBSOc6H3Vkv3u+nPo70
kc9pIRzCeuerEgEZghKelVtVSOL+6+/WmpneKlKSh7Xk3Qc3NZE6N55FdxeK8Ubi69eTNOlHIgvQ
avBG0Tp6ICZdv9eNHT893aAlNOg6x/dgMCc049Usa3zHaHHuAiZJgmlnd7IW3mf0R1Lea+ZAxV7B
y5HpsSIHx3KkNPrRBFvp/PpoHZiu/3YKFMRGa2cgokzQo+OpdhC35Dyj4pR8GwBR9cJd5KYXxGC2
vyHE+AUNYKDDn0vwO1pmjM42lLhKw+Jxdx/onB3KdR/LE+R5zLM64/8SaJwSqaYHrHveRN3bEcSe
9VkfLSGQThxbQWGsRy9fIx9XF3+RCWALRRJtPM1DfKGNln+jGRZADoi3mX+GiYYxsVX9ynx373F3
H7IMJTre2nOA5gDRAf+JbsLv/XNV/7ZEHnOpiyl0NFBcj7WUu45eTTU6LJ6EuI5w21qnfskFyTig
qyxIwwrE08jwcsekoq+jdMV3tDIbmb0994epZ0r/0+aZ75qqosLUAPRu9q67TqrIS/+uKK6Fhn4s
rT2GCm0sQNvK/OrFBVQ4g2ybY4CYtR2RZ9K7lH82xtYlpeCwpCAapttS1SqZmHR/ldT41+Ux5BQK
gvSs8fbKQRVi+XkkdzUmkhy3z5pq+1sw8vokm1oCEBSqP16iDebaEww1eTWKmRjRj7baO/FDZdIA
7ov7q+MkwsGxDtiMZ30eB4T+AQbLa9WHe/zAdZeh/aXgiUw/d5ftUL68FTLVur/17Pn1aL0tvk9e
9sCPN2JOYOS4oZyRPq8267VzvPx0eVfO89u9gxp8/NhB9eOiDM4p96ZRoFDuHtHBf+CpFUjUo2EZ
9H0Hz0yw1S3w54ha2YvqMAH4hm8icexVIOTYcZIx7ABwloWqLQ+UgW1KeQMWi3ckXhUui0YqlpRG
SSraJR0b7zvfXuXgFz+y1OmSy/dHwf0ttboDxqBARXOjW5W94XJBCiLjo1V3rjpZfQVljtR1TdhZ
1iJ/CiZxjb2sqzZJDwS0eOct6ULvzlGMsbhSm0GYURIemS/zZX3L8OruxCO7SBvpnvEBbwOgRv6h
KTOb+jTiQ9hz7rQawVLsXEYR7Amx6XKu+AuXfHlMoPL1XvfvnAREnRZkfGOfZzY62fL63j5kdvK6
wp7BIqsACOXTy3TXZ1Z1qJxnOSn+1lQ2tVZ01xiEfUdmDl9AfEUw25g9SXVBlGcbqCkISj7Y78Tb
AOMMbdtVDczZqJmsR/Bx0TMpe2Y7/RpQmlFSigGaRtj9LjqeSp719hUB0WuUg56l9yqNZ/IVZXsU
koAZHSbpLldhR408+ZQM+HWJvhZ0+VMagMdlTpPNIXZXKzdmoFELERFRQLPTtfwbYvkufnkSKnI9
DAaZSCv+L3LFECkukW8qUf8LDVhpQU28QBqHeyyYELm/4kkvG9SQ4r+2bT2H8xOIYqSbLnhyj1Gu
hn3ww2P0QiDPfoEQbaGSPVYWg3p+9p7vLnvVYrbXe7x9Fy+SnMOhjK7Bjl9jqVpsAivl7R16ngt0
HLNyjepK0kxFccM1TR0b2/F/kIw0oBTWyk/ZIuUSSSJkHbd/GK3jCNdypMkNjHbGQZdX5H+LNImI
18gmxC67JqCVz4gZ6tCikgJwOFB95OpM1JxNH0HXbTl/j0ljtFdgy7YsoU1bOXNdHeZ0l3I23qHA
9VILB1DI6xbfV8PR1DORnVdYK+1zlcS5T3golX/cz6yX48lX9GyhrU/UmBiYiNSMlUPoNSpZlyRC
xORmXgrUPQ+lZiGoSxw0va82ng3KhXVyp+g6f5BEOeXik3AoviuK9k4bncIgH1i6XFefzn6Rn3w6
+GvLNFSImmBhP+jAPPXPgx3IbfcvGlSipWW44M966qd12bKsfvuMNQDTFOkr6Q+vnEil+DgBQR+a
4gkZ/8uCguJMfWu1hg5eSiaozY8uN5Au4RJ71fb+ApaVwi0pQ42MsCfzyRlW9EcsagjxLnrKvWF3
z3JiD0o6A/u7EDfKcDPqPOz1gDuWrfjNcLS6rKQ7+SNOJaeKWu2gl1rEzvMB+/HZ4vzNQWb0nJhm
6wZbWwroMXHRroUumwD7kKAutVmWjOksYcqenzyBa3+L81xiiYpVWpwHwP3Q4ycX6E+RL8tfmuZ+
mc7WnhKsZsbtAG+8cQ+Gof4gEwGepKa4lkTl2Yr5BhkQ9cWoBAADeL4CF/++oGttDK/Ys+poeiwd
fWW3BUhV1yn5t1FEobIx+SjrRHwNhAKOwEAR63SVM3cpsRDX0HN99HhMXbZ0QAxClP+HBHjFi6OM
tHlv/WmGX2qmLt/9Z6IMkvlKaOaZaRi3A7y2dzBIffPULUI7j+xvQHWpJiYtMAgFODXmUWVk/u9P
gIcwSS7E6FdkkCLz3me9TeitaMYwIcG+O1P4xUxLm4TjbFutVsV0SlXsTyfRdVoKQDmbX3/levGm
QCzE+8rTJRFF7oGYz6+4SgxlE+H7gCA1ErNbbMwVvn9JmKUBK7tA6YW8/qjbJm9hgI71ZSKRoxOy
LR+ZYv4jWy8u1OzdS7MFAk7EIgkTOodOzU1cbsHtym+b1/ZLhVZo9adRXARs2gmO5kDCsLgwiTA3
z+sSlFXXnrEVbLBJStYB2LvWXLTf2KlW/2/9vj5e0uPSMn8Y6+Jk1YQ9Xj5ALRfX561Il3h3zm9I
VOhK49OQFxabgtcNh+5nEnvJReaqf5l6/J7+Eb+h2knAQMRiBVs6+EJvuTKfNXzVajDv47P1P0iD
XL9qUZVAEA5oxit1iMJRa9nyVzcfOJBm6U9uN4AOsAwl8fdpfue+HUpURFVsMa3v4JJhQvekox8s
sW+LTAA7k2zvocB6+VdJaXbDLuLNNVpJK2oHQzF53CwlPzA14qn1IlPlnMtkl4OmkYYFO2uulzJD
gIVqmvpUpKZFxiWRIFSCH0NAHO+BNwss87fT2xqTMF1a7bvGF/hv6sLtUoKnLYOj2F5b6jkeHJBF
MwJTLa2Vja2jJRh3ujS9WkPSPx6Gt7HvS77MsWOnAGehmGeftRSMOWpZGHxrBN2OfuQfrSHNgZyk
llLldMl2b03Lp2W5gzdHsTme3T9p8RHgXbknategu6lLvpbthMhS6AP9h+MQvFItxpcsJT5mHFFw
HAcQOg28IXpo/mXGz7z+XjDMFL5EN7pCK63j8qeHxrbTdMSX/vVA3G0RuqRBqJj6TcsQHQe6qQVE
ptZKFk+Iot7/bKPiccMQPDAVhVb7JN2jtSZjV23LILTeqbjvz6u57thC1u8jOSMUvol45mFAHntW
NX+P3rdgqVHHryugy/bpdZLeQ3DVAVda1GcNBgQn+jRID/ENd2yG2/JbO2b6D2CTubc90JjCGPxG
LLYEj6HUAjwInF3CWM/4DbkUmjt0TB4oaj6zpSmqwmsWjgTf3pvtFsGqMjAGnQXOVdGGtS0/UcGH
gMbWft7Lf6APhgw12/oYRcRCDmcdTjkpViJ/DACueteF06TvKVStynEJkGjm9y3eX8Jr8qKPewdT
tNd35zdSbQr46QFXu8kC/3RdhzFyfo36TYYSuAgmMiOFZf6GHCLC+mKvjNqzPEJOPtbfG+C6TDqZ
E6uk0tzmYHQqkcMVB6oVy8pE6HDBjZP070kbFRPhrdfAKaTDBZMQwGZ02+C5fpgpw03rIJcyitlf
AcxcVV55VLkjrNZJ9Dt05BFzO0yULcjWV1cTE7ippL5WOEwCv6EoH78oHSEy3LZ2Xe7Cbcri+E9d
Zqx6f5mOnhrdxIuRoQ+3PXf7Jj/b8e54JrzzlNX5bfTCMS8OBhH7UPZa7pkNj69wYtqgcnvKP6WZ
DxxF6etIq33g+fHFzzBcPHDes5lN0gQaq1+8BMsdqkkQpxbGlb29woCg6Dico3utllOrg/KSg4Wc
9Dz/QU3XJSZ4HYrfYAZmTgbRPTbhSeLosRj9foejA5MQtxioUQmZNoRxxQnj+j4i103MjdlL7oFe
+g4Cvs9FmRYq4EUMYcavwi5uNlv9jgR0mrwT0fmti0H1UHlCZtVoNIkGZRafSilbeQ+ee2NalmKX
kLX4ligLCNFoUcntPdYqXCkTQ1k1EqTL2s+UvO8lsw7OqnlPxLR9hg1p6ZOPWlYQ/EMYX26xBc1L
dc4nGzK/9FK31+u8Mcl8Qk/0rJz7RwyShGYMBVqnXLhcaSwFnnLl8UkER5I5iiYg0RxDj6Fk7GQM
xXxwEHyHBBWBBcQLZnEZga0CcBflXl0GfUYEMy3+4KMAvKgO4pO1Axdi8b0gG72w+YiK0V+T89jD
Fg5GGkuxyakxCv0zhxCbPRrNfNAcPJDnzqoCnkl0Ay98RrJ8KnqFiDse0uHGdpiEpQdS0ONAAagV
LcbmdQPUsvVzo92FBrw1baF5B2QzTEehgc5VYOYeRiGxKs7I5nOLDrfOsV43RkA6vkFtJ02zJpAm
2WH0kA9WSJjhyPzbcv43rvwtOKV/LfwazpubBmqzMo+zzTdr/KYx88EbM4Ae5ZgB9zPnqMhBEVZu
6nQPGCQIaqleBjn9FXWy8a6Jd+oBp4i1Gzzt6UOWY3pYGPTl+yvTjBLn3Dw7xYOPfregMmXTwh70
eywBZCqZDJz7LtujCSZRg9835aEc5vbbuSUbqlYSi0DcerLrI90zKTaOL6sOyIALsddiVP1eZTvO
xqGq6O8/x/HQ8sdmoO9/PTeZ2LRUZmSdkzuMyZj2QgH40Lm059uIkvHvxE2Nfl76MCBC4tWjX/5R
t15+HBYlGCp96KRVwr2LiUaf4dLR53Be63Yih2uM0t8vMbw+vG289Vrs7sXI8O0fHu+cb2HokTHD
OJ7AnB4iTsrFPuQ45mZVuINBCl1JHdsmnqINZLVdzNwJGKGfx6pf0CPoLEgr5gIHi3NcaSZigN9W
fhlrzaWoHbAGB5ruKmXmPIqQrrhn36a+dj40mv62CxfwRV7luyETG1hOlwIZ8TDVqQWvI7IZH3ZH
k6RN09EvvUBHDlPMBKn+r+9ET4w14y/aJAVt5/BqWbqDqrbFNM2CF1jEWp9rNBHgheLCkYY6NCJB
78Jr6iTezHx9tDRT9006Pm9ihG8fPa/1gyCsdu09l9EUhwOndKCo9J0Ew06EhexnkFIMnMtxOpga
8AYl06Oohveot0jVjORYjLs4CJAHDnQWbsCcuTZI6ZyOD4nVC2FiPPf1pdx5KvgVl1we8FBo0v6F
8IJZOUSZtQI2IAenj558mhtbZQCwt8j/SJu4U4/WhTXCrEq4OXpJFW0PgC0fkqOQEGjmUTsuAYkH
w/ypqRsf1EHmIjVeCbRiJemLNYSvVyaj3sNou+3ZO8OkWa6uMMZpf5aTwC3ku+bXZVEJO1Y1h8ME
9ZpK+u3FPeuhX7MM9It5cmYeg452R3CioZTcxhJtMYVyia+YyWd+aQORcCoysbs89httMTJ6pJ2x
mHO8WREbuKJftxR4tuZX+cTvlu2T0koiPn7c3I46jFBUAEtuYlKEbBfcNyT99alU9gD4/cP9TfgZ
nUr0h11sTeHBhDVc8ADJ2QMCE9jGDLPGvgIUuq2J5uYLb1rTsuJQEjX9MkMv4UFbkU5JbjQfX2E0
/1EZHnS0BdXrCEJInFlitLi5xX3NjA4T2UHsnhvb2yKq115K+/23BEHmNhhZmfFg/D8FXx8gOhCx
hFMFmAVjCPT4g5jerHfOygeTfuUVOrNSAy4grSoq7Ot2U8s2mlpuwwiW3xEynUd0PzvSiDDA0i+E
zOvVuHhOi3EiUb0bR+SPCgOa/waskLgOksF9uND9jPIlo4uGio3Cpiru+lTKh90IaHMO22Ga1xe9
u53N3R2IuWbxe9ej9S4OWMlMdZaQmJ6ItAmskuGT8zdJOwjLVEl3TfgUt/3fRe3rD++2l4D2U5Is
hptbXHbbK7quZxt3vLJeNCqFDnI9RNU3UxD+2gCqJ/RjYxTx6l/c0pk/0r3UQTxKMIaUYZtBMM9C
nA6Xa4bUHXF3S0hcxaGMxp/qsdIgmYYaQsC7iKf4XhLLfCmWOzmG823lP9oxl7t8XWheAb7uqqfX
Qk+phKAeeUyzj4Poqz59Dopp3BxHEximrIp/ozxhA68OI0a0p4FGYMUgclKEZN1nRW24gYv4jk14
K2C2fQFVZ58AkUQQQ2wN+QvUsrn3eJg3l8EZvIGKOVVgqEoKsYiYitB4O0My2P0xtYxlM2aBypOv
sbMB6G4N8fC0Fjq1ekEMG+FtqJ15f4v2cR+uy4Ix0VnKcRsgdckoIuRrV7eVz9Bppwsll+u5kh67
jYnZm457roeoINZtsi0Fxt5B5U6TowNC07uh6Vh4/IqQiTtZFsgBOcPhp9/vQHtjLnD0m1XH0eI8
2RSijln8M3BUT43kQBd0n8jZV0RoilFpLNdS8WZDnJMhhKdIbxdFLA8Kc7M6rNpLdl2pL0Ph1L8a
LxhvdlA9PshUke7LxHuf6K5Bx4Om2adLft2eiQRRsYq6YfTKM9TlsWjRgUKk8KuM0Q97XtNIjbzl
FB2V/7dRQCnKjqIOImyOxOcF9EaEXoLmb1yP9Qgke3mO5DzHL0e1ss9GgWaqPEi1a7diGyyp4MZ6
0+hIA7L99NIJ8/HU/31DORe6CMCN63PKxvesrAhY6ZxDKi/RU7tHFbwEr14uwt5NNDAdscWWuLk5
nxymRkLU8THef37jVZ6ZmSISH3qy52UR5AO58lrLaS3v7Wg4NrS6Jp5f7Rnk0EzwEjURxua0P35n
Yvi8MYHW/L0xm5gJpBsXS4i60SC7cjEciBuASdJT4Q5d46p8lLzEFGLo2tL6NrIyoZdCb1R5DEWP
RCTAnjYt6pQhg9zDhQgNq2zykx+y8W0CLagAYCeNu2Fq7z/Lobvr+EciOD3Z8d7y0HeIiVSlM0jz
1vmzCmvUnhFt5pXMxnEmA2aSB0X09P5ehJcCublG1K3ZHO93jzdypQQIF0lUGYarKk7yumaX+p5U
hVrF3pjisdM8b+axv/ExC6nWChpkeTzAyBdE78pbAvIPxmXyFssWLv7+K1twvJuQkaXNfiJC+Nuj
tgkkzR2XQMDz7kwEAJuKuVBLKJvzNK5N7rWxo8XSJROFJrv78IZrKjmSeRokz4jHl0O5CuDLE01t
RnDugXOwLVDRSsKrNz7i/uwjdFUYSTjRZkm6fWOwUKQzWz+j+eDqNz9NjjlQ0WJLX/CkyWSCnNYv
HzVRA9p0GEwOFF3r2f+HtGqw/AD/rG7ff34xfDzDFFYiGy4wuwWy8wj1p/s32YAWY5VVMuQjXJ8A
WlP4XqOzfkzYYNMY34ZMgi2Z+9s/04DgmayQ8jqMcZysqKaFpYlmten6ORiXk311XF/WafZppB8P
1mpTBNvWRs0ybkRPkLYDCF/mFk16vyhWEp6XnTrvEQQC/vsdzXsvbeafwikTRhjM6rJ6bFJORJSy
eO1ysNicoGk8kut7wu2GnUJq2tdtJUvoU2LvBtMLaE4+Hu/awGh7HuS0FAyeV/bd/PsbAmrziMJe
p55AY8f9bKihlMNiTro5ZZJqLf8yI7e6xRrOpFJsa9PtBPSLNSGtEsN20MwhbqzHmwN2m1AOQ2Du
pGjZHn81m38LYZVx8RDTHUndyz7d5wPU+r05gli8ZrpZFHiVri14eUy/1KHtkURxAHNT7XCSotP9
kbN2ba38PajBghEHNm+p+3L5SuLGzW79Ck5w1eh0ExT2zrr1dkSPstkoF0N0XAinRRmYHXtBn4e+
G/5vPMb0H7iaRBzscaH9Xe8wqMI64qEaFuFzrU6PmDbtkpOUHU9GN0cIPintcdrmazn0bBrDAM2L
cyNXYpDJTP/6e0dkxxC0SBRnZM2ryzc/sqRrsjVZzdHRg4dum2mZe66TEJe7D7nhqkgh+sZIB6xp
BJdsOq2c7yE1aIo1m3CvURoijO9KhkPOihFcodnzuS9uPNitOPKtwF/uSW67BMHmGyqXEfp5mOlx
rtsVo65pbWitri6zjn38Gdsh9hwuwTnrloDO/MtZCwOX+58UN7g2kTtC3qOyHXriN7uiPZGbtmYT
hvvB8L8URGWgAPPJ3zf1sJ5LPiQijaI0V+BquB2jg04bpgeRxnbs1kp6xz59s2TKknZ7B8g8Y//T
syJNLhdhJteexu1fq0ja3izD14j7T3jdyXmFRUucWlKawymPLXVc5I+27W/fOYHRiD7ZV73QsjKj
nCOb+Z1jvIvxiuTaO1/pjAuC5KmGN4Gs8gG1ZSvlOpbGSOaNKgwCe7jX8o6fam1r4UoLFnx3DiQu
jG8ODeG5Kg8hJiPaPgCFvmxeBY/4YMdE+TBoaGEyS0BKK4/js19OO01T8VWaNEuavBiTrvzjhBpp
nbdkyIUzVREDmQ7nw7IwTh/X4COPrrKU51GmO9NPK1tOJtN4zkPwwhXU5KDkinIWWLprdtX/jvsm
zFvZI0aPT8JmqkQAGGtXr7ztmvxj1uL+HHnl86HInPW/r5vXBPce/qySx0YnV1J0411kL4eZZizd
vgIgW8U+qGBkYFE2LTTc9CEYoVlfhtp3RmcG+ccTHqbNR6wJ4nPKGiixjbnAlOxi1i883DQO9t93
0l4QsvlTrWyywYhTKEGUcqQU6A85nMIHdNTazu9nbTe/N3J6Um6DZg4khZfLcijDMkeqR7CEHfLA
6F8EglqjPJzG4HMJjBxXwJ6dhKx0IvfCQi4+ihp1WNhjir+ojgh92ezJjKZBzK8UhsP3qGLcGja0
m1Qh6xM3G8cgjFFzA0DxKPI+8CUf8AKHSSamXRu75Q1va6bhZJpIyfGK91gzd3Xu0HfNKV6rxqcc
Vo3xr2xooWPoyDMjz937nsW/RlZxsLGr1yOLl4EwqPj41uLNXl6Ruz7T4qcgUCj18T7BSezKACr+
PCYAiZ9cc3OdBvOVY28EonjK8jA9vf0+K36++KQqkNxXfrS890TnFzn2fyO+R3p5+U3tM8XglfJm
2Krf+9q8ZbCOzlQQEev9nTpK+nZd3ImC6PHzNnP5ToPZF58i/R9fbG4iTH4LoQH6lj7flJ9igWET
6U6UVVV0ejtBgbg6M2RLZL5V78mqtz/Se5TUUmSsbJh397ttu7mP5wdpFyFMhEVQ8hbY9dnuFT2K
hPQp/Kv5O9kT6gzuLkAaV7v0mci3CDrtSqZKXZNX2dqyRvWwEwsA9hN5Bc6XWs0WDWGJDADinonI
k3skQdst50dl15MGNB0ctzut3Kg5OVMvRiMyumlhA7MIYYRjzgZ2mA7Je5dTwuQFFOqnt4E3KcuT
YoPEaXDL6pbkWX0coom/0/MGhBliN4evDXb7h3oAbuZJamvVg2eRa6/vpQUuaYXUDK/+4PJQYGXA
az4HXhj+zm3FmowWkm4180aMQpYy13OUeWVvv/KeVGwxZ8XYPvZ+0lwNy+OYIx549AGBm30z7v4a
E6Z9zHNp5fRvKCQ4NCRBtQ9iIYaqEl0R5nOdhB4VYhI/snOGxPhIox2aTxRGV2OGQEIlu2uHthaU
iy1tQrkqaWQPHERBqRpFbA6uD9kPyCao8sQCkrRdPHSb6dt7muLi0QUlvIY6pvfj7nGenOrDwftF
s3NtUZWCYwSxxeAgdIvFUlkVzGRFyu+6rHEdlPxx+tLOccNfiQLTDQCeAIOwB/mg5g/GG/9jkGyb
q+pBuIOEKPMt7aBxjOS1DpJ62JjDY2XiU/CGuA87vW30iqHYK1TDGlgLaYjAhpMLFeLRTdhmBP9+
HcmzCt0oOKmv8Yv0ucLr8iLaoN/LzEI6F/o86h9ip69Xa7B+UsrZFI2Cuas/ZYT+xi/ekt1cd2Ux
Nc8bqF9dm2Umktte62xR9WxSfOJBhL69UAmf8d55hP48IKQurX7LSVzGp/hbAXEdTC/Xak9nYvQe
A3fIUpRTXctVXtqbpp29mKyM/mtPXCi5IYUBr8wxgOlsGKtUnQJVTU+/+LHmoQdQPL8Cl+C10Dgp
Jnfd5nCNi56P17yUCOStEYcKFPy53/F00Rv3QqJATOd2H8nHqt1RpPaLzmNh9zjkqmNpcY0/dDpN
rxL145gAm44DEP7U282sWknOQbACaUcMQB43hmi5B9qyAQpJkIVFqhHKLhEemxV4BApG6PVoyx7Q
GBED2cNguSaXQ0DsuIcfJEToa2UWdDrvM0AEsRu7ln4ct5e1MM+G41iV91DwD7ETlNAM64SVmmI3
0on+XBZxfp05dGmL2GDvTVNdnV2fZSTUatCMSYbHl8dp7mEOE1ByLTcMfICMVfS16JjeRgYI8+ht
L+OOGSRCZiVffjjT2xBF6NvnXmFmkohY5yKb8aWJzE/sxA4Mf6fW4lerSrI6jgLcZB3yS4wcjYfx
ntqJ3YSXmrNa6CI581j5gTugdT0qRtx4FnR+n7H3/uRUDGuJgCYNnaXdNfRFob92UAPQfICxrXDb
lC9K8qG55SA9VpQFJOOKbUVyUvZzfrif8Syqw0ps+AzvXOH0PcDCNpVNcVJKvMJOzCdnRgAcYJjl
b6AD5aYZEGDCskX7F5uQOXc9TYfJ+iYF+Epd1X9hGsP0q/vssy7tRqhIoxppn69a5bv3d3ulJ4iV
rF2KPMRG1IlCZwxUG6o/tpb2f523S1dHWoHtpAnoKT/A5zkFlNQhJ1FxbfYlqNa88lHXjrpvO0w1
oE6I9K5hZh/QV8WPDVhHi6JayKfWiJhmEKiZdqGq2wLvhe+e8wVoZ9vJh6qzJF1tOHnptf2MP/WM
j3wgH+fi1iBUyZVWxSpFzbNKoDK3hUXGPNeFud/TrYBJpV8EfaSj7wCxDt81tNDEJ72Q6rzBKUsA
mr9aQKw73sKeFo0rlc7AQLB7kVxkk3gcNUgSag/udq7QgbjCGpszPuaWx/aiDzAjpFSMif6D8bOz
q6fwWgPGTw8g73FgEMwqmlEjF0LHUDMoDbUzSJES7YdxGKdAbUmlgF97u7cKTRXncBLB0fOJkLvG
44xIvhpo2OTZqnkEuh5dAUzYPjzCmVMFPQ1RtzPobssXDHNT4ejXkpsIC6hXUtdkkHYcjB7k82Vz
kPWUmpRdS1jq5eAKBhuAiFWAXhQ24a2kbmV+0m2vzHY3XIU3vHE5MeJxw35O7/OCvRclImcyBJ5+
oN1dkS6SxKJKnQwbJk9KvGnnjI9PIC5CQOawiQPLoDEug+wGmqx9lsXR1u19d9tSXKZDU9xXHOcO
jN8sj2CVn/uZB1BL5z63DprH4aRAIQflq/Lqq6Wq69wSHMn1IBqD3Ug2lfakXfOB4YM/dCnXIAxI
BYu/hRdR0FY44WFRqMh+s4TpMfbZXGmOEPr7jdDUmrlGzexolUa3fMKoi/6HkdVGpAscFLpt/x15
E90fjdI32zl5Ul1cxozaPVaWp4JJQI3jvWtrc2YeZhDgE4QEE69Uzuc7KUVclCNRb7+mr8bOrskl
fz46feZE0P8iPD7QdJbDUumVzKPQn20VwmK98GJVeHdbIJdiJQRD7LnXqtoguhhYFgZFOg+9zcD/
o6MIpRC5xDzjD6mW8EzPdNn9AlwUS4w0qA25fVe/ZPZNXhKVQHGVUJ2LkmZTUplCzwD9Qz60Kuei
cNfVN4aG3BPhU+6eXOCWbp8/eBGHn/ILP3xrMApENLlsOf3YGUI9lT30Mp5N3uo1+SXwhcUgbDHG
frU92TXnEjyqVB4cABujjcbN8WugFrLZEgXftlpIjV8KoZyK5RRgLnwhNLNniZCtkAzzZSrrtPVw
k7TgNfIXPhl/0MBVc1N5DSvnziJHn2hG3P1RYaoU0Wa1PxgBo5F5ziCWovMlU/GGOUB1zf3sVUVK
JgrtX7O0yWiRUfSh3VWUXpROUkXjZI06UnXjc9Jtz4RL5V2VS/pFWtIJqx1V1vDq7qug2WmAwNM5
uiuBt/0B2GlaQRhmfC5LuP150keCRPYOPCL29KtmDxNiIQD7dM2li5J84KalZvNfd7bgksSC3waX
YoHnmrfgc2lBzHYcQCL0sXnO2gp4mHxl6UHGCJNakT+xhcvYWrG1195diBnxQvB7Emu1cTBG6ihP
w7XmPjrZa4Ux1N1kd3JHebzYMC0DQ8FHeCZoM8nwhEMoYek7dq+QOPoMldNGDVFYRi9icfF2DGSd
XLM1J0F7VM4if21vvR1jntq9rxpuJCVDP38crPyDAv3DaTBeKDY6kME0aAGh+uV4pRRlAwaf1+ap
9OgsMiU7zdKU6ya4e1ZfVnM+bS3t3vBL1mWl7KfODudTKyqVHxK/XDMKtbCs+ZRWx+gUgf7I8peU
HFBdZzlXZ55WKWoUN1VnItqf1Je7mOxnxExwOJczKk4Wv48v4ZqtJvVO1o2KMrLGQ0k2kV7YiTo7
CDU2kLvDy1yGGATcfopqTqAKnara6cqTv7TC33O0CGBwNfgqHP4KKPcFAYCyjEOxGGmk50adBMTM
Pec3Wvt4ICVT41uv8V96BZxVkyvyqk3/k6Zfaz+tXMa4sOI3rBo8hbFCeknn7QpwpL4/jkGAuTis
6e1J2WLcxEphCerP7dmaJ+Sz5vdDKQ9XBCZ9HLWx90+JhdXY9A1CgEGgzNaSh5YtyGleCTd5yDSC
GdQ9IOUFu0UW+fAQf1h20Z3BwkI4GDHHK0S5fENXw0P2HJROiHjDUS++X3i3UjRenFyZlG7phSWQ
uGbC0ZYz/YBQqJ9Mv6plT6vtYviUVFqBYNaKra+GeM3QGQHN1rPXbWBpXYrjrb6JfMaCpe92xlJl
v6sarkOBz7mpE4+VU96J9E2gRRq78qkHt0GtLnhsjb4BmDuvtJ+b/5wD5Win+goQW4VCeLCiYLJb
OJf5E77d23wfkKyxK7uv62RrLdz23i23McdwpPwjcFqBenvo0eriztCLvsVI7q8Rc8luUre0B5XU
gVjyEEYaD5RPpAOuN/0FYGXkTu7Y3CMPLyqSQQSEaOftIgcRu/iq4jzF2XX9j/ixtMAVuiV8whUN
HZAtwIJeUW16k7z43qfQdCCFNnu/AKG+tz7NeWyfWoHvvmCli22ZmPlpUarBDfqRe37W/mXvVJrL
7OWBifP4W5xxDrjwP/K+jDM0sUrJR7ysRM3K8zfKCAaKnuvwRrCIBeLI/7B8/fLbJaTOcFpA/d9H
vn5HE/F4E3eDoaebYm7zgRPgZ6Iyb0VZfKdZ8mFFJf+D5/7I5lYDtGz9L6YphHfLqRQUITs1t4t4
L60/Q5cx1BHvaDEsCpa9dS+LMtOkNkpMofBMr1NlAalg207H155mI+rm6XIuS/Uy02/LcF5V0Jbr
X1WRCtEJY/s4GLqr4Ar1oQJGgfsjnd8M2RfRc0dYvW90NW1px3xprSt5wuAso1Jj2ZtleXDnbi17
Jc1AvLFcn//QdmcQ6T/Q2ht1FW5IgcB0B6F0613kZ60aOebZYR7bQVYKOi7xPPv8oUNg6cCi4bNi
3NMU/S0aROe6b/KZ74oDLeM6eGC49n3BeimqIbk8s4aX0Li+8hSpYjYSoOxaYE3/Fl9wx6hvrOLo
JnMcVxLtQlJsP0Q3PNpPalsprucSkwyv72n1ZvmHOFa0Oe2x/i7BRpB028IuMcdxLmv8lbr5tTch
pYWUgwZlP0QrQ126j+5V04Z8+eSIDy3lBACpiBtPV2HlmmCXsdFBPWrq3T2aiP89RauoBlqHtq7v
D9H7V6Sp8FEnPo6UYg2jAwW4Bcs1JzzHOnCb95evU2R+mTTggxD30N3xTKC52fMDToyx+3hHtZPr
L55mxQxdnzrRJQkLI7JTjPhAHVSuTSaAjYGgAiE/kIbmvhazSbsTGKxA6vzIA0QFyEvSDAdGwV9b
GqriJHIrzZYIjPxLHXVXGsz7m86Fl6nPIqeLmNutWUPEgGQFIkPH8Iyfy9P6y3uRpGxn84ENkI+k
KIgNCqjDHmWRcHoMfwmdoXPN3XfK0wSz5RThuA91UdpmGEwEMajibxa3RFlCgYjij3Rl9xyW6QHF
KHhGmlT7SpxEM4n781zY2GVMYiQ3k/tC2i3nfdsxT4t869JVxyrMG/l31KoaDsQDc7Ki/LYg7D/Y
vEjsKHy6Scq9EyVD9FVll52NJJbx0nE7QaDZf8Qo4UzDNPQd0BDu/xMrYXmAhwY4aC8ncKbhZ3cL
gzb12K9t5ekXnmrV6jBFXZgaRk7e5I2eNHNKYw3WY7LUvnB0SUpzj108As/oIpxviu0cUUbWAdbK
5tyzeaG9+hwiAHZ2WL4uF9E9mhrctlFVp8rTE6RP+mTXtjVcWFp9sHcbUupMwGmg2EOLInzk6Dy1
mfJWCTBotP8sqKxhYJVP+0FlDtGWJrG7n5Qv8gqcSpr4oZIMPL5+d/fdxPKAv/6EeW9UoaVN348H
FdDB8XKu+5oMZBshnx50WnFMTS6hBI8rXV2f24bX7yl7HP7Np35H0YB7B5lc/QQAfb/lmRdwG6C6
PodU/6RjyKCSX8YI3gI5CkziOiaRweXUcWqObm4jJdvocbjzGrcGW3Mpjqf5mISM1GrIo2Sb5tOV
H9R37NEcK4sYyjcwd1moaA6k70jnFJmyGGmiT8jpFIsu0YcyvMuXSUdOAaVM7vMKRga2ZCNwQ01I
d5PaBXocVWAgy8FvE0es24bPXJHkxwJmi0kseU/9tiYm/GMomzPZhhuk8UnEUKDYousx9Zz9x3Xv
1SCGH3SzXZxoIT64+SRMaI6wDB2OT24NFdqxrYCtPHU69MFgsumy1uuGNp0DFZF+PCiPl+69a0cu
EfpKIJ9PstnkSSXkYA/4HyTmBEm9ny6ovBiPAOWz7CiqqG5XBZuCj2PKhbqioPBIztBPOoClIO1P
f5WS2L2tL6tjF7AcP57152gP4CINuJAcS4lKfqCO2gM8AAADq+rDXbugyLGSdd0jorIKMFGza5Cm
/ivuTj15JZfuCUlaoNS00LrmTXWWoE6zNXKTBPwzHdqh3d57vm5lSkpvIE7U/XaW3yGA9Mz4sP9u
EYI978vc4zSTHAJNJz1Fbwb4iRcwwmU78hYcjq2730ONIupb0I8q5vXYlBkebqCNtIaNO5df2wir
cu6C9+d1pEieFcwGpgLn4XjqSNNke8eSPbzcKxBs3fCveXnG5KYRlGxHnH9bQxjq4QujUOCWBhtK
Wn1PhLPQKmZWlsb0n7/CkgTQX6HCu2iFhUymgdkeKhFQE/ul40OfSm4YOJRxvP265mDZNGMKd+q9
A8hUuRLzsDXO1rgq/ifZuDW64ESruVQ4YKNYD7N29YLYgMFNj3XxNBx/whkKHi2P2/0q1HQOADaY
bRXMSuy+z68aRnl1bqX6uW1TXilKMzCSoFLfLxbjsqrsu8hJldBICV8UBvQAVDWrMVH9K0wox1O2
5LFawHmTFJxKysF1DGX8uCdsTWyZ313deNq8ygZEG1GPFuttnn4WcD2vVL6DBl3KnKluXOH1BjGf
r7r8fQornKe1XnoQkE9J2jqlTsQvs2x49sliBAtxvv7rpUu4ELyqkoZwsnITPHi0pA2b7jhr9dgL
wASXmybu8cQF3thpC0hDlHw/BG2etoyOjiXDWgbs/WvMMy5mNxEsgs18NAbRg0GJpjLsPNUlz0TV
sryS9pPzCRDMwElRz0NGewVXDVAvl8xHa51Xt99p1JDHy01QHeOptQYUhuOaU7dxZtqsHR1MHFmo
mfLVnzITt8u3sZ+PYDYNwYBVRfxb3RWqCH9VtpF4nzI5Zqc6FnIeXHAydRNBM9o2Z8CP0O4nes7u
9rfo6s5059+BMG1dgAhGL0buW0JqghKu3bhvtQ1hsNLrSoupxMceF8MAApKa3ZoOMG0pvUOQM/Nj
rOKcmQOV0YrwQzoffK0wsXFBs5goBv/Ysy7atV2tE1vADhJRZN737zkvLKg4BNyyTyPsuX9Gb2Y4
CMi1j6TlQko+l3CgQNW8ghOZdD7ZSk4oNW9PV8qlMO7hBCzYICILFJ5Ry8P1jo9egx1JuaMxWvoR
Em8rCvelC1IqZOK12U3/hqv23ITGQ4qVuSlPRSDgdMhIVPir9PsiDmiaR+Fdfk5qyU2vGmdHkHVo
IcI6U42sUq15iBv47XpWke/zKiN8fqVjdjQ/cKdPuj0+z/H1DvGaY06ulVYZADUwsOhQ2rlyadoH
2w1zzFOisHWWPMbGzDxyMgxKKP2rnkiAhk3A0aw7J+d4hRt2I590eqWM5scADRP/0DlCT/9yLhyf
aC6e61rFO7rWxK3lwZXmGL2JVSqKDP8mpYJc4W+YZyDZ/ZoVPYEXfSc2e9jjN/QjHr9UMOVOgE6L
QY7FnrQzaiSsL3m0SK4PmAuk+anZ01ae8OL8ZLTKEYcp4Dow37lxHrNmSk/+hZECJ8HHbYyde8GU
ML+0uLbjHFn6EjuJ9RP4mqfYYN3yoqB0koYXFumtXFS0FXWGgPBk892A8PjjT7AUNp+uNTeZ/i67
08gPVtw/qvu1FQyD3qVQvt/VjS66NsvF6LJABC+1gy6O7h2yYOieDYmrABEI/l4jwWG8PVYtnQcu
sq2nNi8RpTbqhFsXMI86ONsVOHbYQwRpBd2QEpFJTD8mP34JbkD4LB4SS9fh4M8k8DSb9OZ5oMp0
2PF0nZcow/YD7Y/tLzHszWhXcwWGaBOd3ESLSWStBSq3iNQNa329qpx3OcA6pEESHqDdziZzkh6W
BBvHuKQzZbekcdOwW8yMXDgq5+bHSfRilF3m5rC7Ivc0AVBFJ/fmMQ5MUYfOXIfKFexYnzs1OgDn
zKuEIpvYcMz8MkLHM6Up2IE4yFJ7lc6NuLEA/LXWDNBn2t5fE1m10QD2ovJHk8d6R59PfL4Yg4ap
gE1ISBGWIGFfi4zAjeGDA9HYIYOJrQEXmZTcIGw5wULtuipKTnk9Nkvk5soVpq1JFqqR3L2i99xE
vHxKyl0mk19aU9kCMatzJDZ+93i88kDMIRWyaJYqEceHUS4QCQfsF7bC3MihhI6vLSV1EgljbaQd
fWpYeMILy8Eod+s84n96qiHPVWTMfLgXlTlbVogeDP4uUDvWmBTKY2coDHK/ePJhyAludFjluJae
seuL5hOgslMbHItt78/JDF1fOUDuIkifuZoPAUhrO+DU3/T2yrjgGUORm3+ZTtpSmBknawVJ1rNJ
XsmJ5v5dsub7DJqABNpAn8zDOkx6O+FO+0AtzSvmPcU/l4mqKF9lPlEZNY5s3bEbyu0dg371RRRX
bFGvI8a97Tjm+O/g6BYI3tKrPYCw2eAue+fXo9wq75ddwexaIYWOTr/ygROA1tL03GSKEJO0HezB
vcamn+RBHIiEiuu2QTq6NqewZ4riUMLBxICU5cNQJbDBz47tAeXgiqKJ9LjOAfeZ2iAc2pOckFd+
9eu2fKKaq61LPHdK63B06qNMFmbbskgUzaMnBBrFOl7sxaEAs0fD42omtKXrK9TVBmnnA/T/jyEJ
QFHc5finJDgdwmClPcw1pLzhVtYLGEX3VwKrmyOR1EgPApI05KBN/ljl6HnDZQt2e8ljHXC82S/n
DRYec3DLbxydO6Ng7+kmgPLzZpPb5aSDls14HxsZdJhaZnba7X6fBYdtaq103rbkhqEZGiZPnUSp
Ofa+8m9uy8NhbnWEGVqc0NbSmr2j3Dp19tR0Jl2ga/ZdQ2dikUFBUFKACg1ykUEpeaDY06p7itfd
ITY+Xg155OQ+QMKcKvkbS8SMknifNFvjP5/h7vzVXl2V+F/APlNFniMRIjaLZoOGKrEFGxKcVNGD
MhSiYKnf+/PYbAwOOlQPhhetUn6k8SisfENcAiC0AJwESCFW/UtEsAdev7xu90vOoMwD7VbU4xJu
0qWVCgynGcoTT93Uznv9FYkP9TDoO+UA1rKMsVIPGP5qz4Yem3MmYxe35hg7K7kFT3VWb3jDkzUx
Sm85aFp+SDjtDbGHqGiyldNVEKE5VnH1XxsbaYQDTghaOXuKn34ha8rulsk7lCes9g2bo1BsYvb6
qk291Lbv0M35lw4YSCAbYSeYdqjael6Dzu2/XWKk7GsrIaNv+kxzjU3bRxk98xGf14BBnAYBRaBw
4zzin4XIXpgYwsb9R/BrnanKaZA+yTNUYyvuWLj20tYMy7nCoIU/h6T/Betkp7i48lH+S3wnthAL
v6tCn3o4iN13KBvzFF8Eh3RrpbBEcBIRlpo4n7IM25npvbrxbFKYhPhRcAwuFZcnVrMHRc5d8WjS
on6eO33vJLeqnWTvSOnGcC0coOyYRERU0PhZfuQ5Or3k6pRXGdffqL0s9GIGJtSaGRW8OHc/kM8W
/g30jNQC0S65nSDNA6LGE8ZB5+z2texjct+hQqO2RAz9cExtPgpgzdR21foAqDv+x3vQYUw6dPla
El11b4t+aCrAcTL9t0B3mt8lsRoiyvrJd29wBYFLBExpe9izsBjKkQKIUaTVD8NH49F+XVpN/MqY
D08Ny2YikuDik9D0065N+XsfrB2feqbJmCkyP1BmS1dE6DL1geBkv4yfV2U4uSSiBzepfxHovmqC
S0aswx9rI8kv7BLwIrWlueKkbnVmwIjFszp4enc4guOhlirFFHcYs/Be9DpdmAWjb4UwlRBdfBdh
OhlN0ZwAtfZ2ARTVOXPUvvn59OOfsE/SHhZXw5i5mGr3dtAxSKlbrzhWLNPoEQkZ5a0c23mf2L4n
8mhqcA9+gXPZLj1R43GghlC33pg5AukGAdBDZXkddZwnSWx/S9w+/ngJT13fN420h0EAIsu9r9Rn
pJ3rJhYNpy+HzrWSwxEG/GaRLJTt2WK+MJESX4lXAR2GZ0bvT1J3UB4FE/fBdmCONwAnTPavt3W3
fAo15IMgSzZdkOQ89noyaN9lpMJGe4nm+05RT298nUYDLKoNhNs87UB4L3Y+WB/SeNTIJoVwjCvX
dcW1gO3MEesFgyceZ9Dk462Opxvu8g4ka1QfCT1ZO1B/8LlnvdYZLSDj/u8jLKZtSL5oKfFj0F8Q
jPaWPXbBrnrUuS93U69TDFuV30UNCXDr6HnbIc438nRO8omDcSZtGv5sCCPRlOjKPZUU52SiDX5o
eFzAU0BQZiuDJjTPs/frfksv6vQJIETrDT/fYsHm/ON3B/9lRIkwJfaY7YyD68sUYps4pbwpKUrV
bxDKpiU2YMxyU90iUQHrHiaorXy5bwcjv161eJetKu7YvjLYAzt+UkG5z8UwNLlRyVLNXK1nJU/b
MZqKce6iB4EqyysPTqQtbvC+a95YIcOko0GaAycOo5VAAws9nTFWuQswEH67N0huxpiPCM/fDWjT
lsGJBKcEPht+i7q9a1n+HR9TN9kaSHhpjh0hmpK1RprvGiXLr1lyp7Xyoim7jScW/LhufQ2Nk/67
YX1Bb6MWsvWvgB9AGDV8+lSi64oF7LYhzqCSeSqUvcUVKw0s7f9XV357/PCbwyOiYEMky3nCIRKD
HcNLhpOAf4yI0rpR7OJWS4jGLA5PCH67+IerGBKep5H4e0382zP6jJb2K98lIqYkutyLVsftLBUx
VeNmR2sfO+RgE/CRsPKnW0UTKAGlcR6wAd8cw8AZEEImgtgGw5rmNy3MVZWuFNdTS9qpd2N1tyVp
jVklmAPLNyAe6FEWaKShpA/OFh5/7y1EznyQ8CBs15rdYBCDuBzfZR/YIDY4oE5ACBFFFLx2spNZ
lVSL0UkkY5bbRmrmo3paU+IQWi/X9ZMQkjsVteJK4kdAwfMu5KJIUPmCREfVaBNTL9QBcxetLs9T
zQahJyQ5piHAj5OynzYcdCGHkiH7i2A09zGrenZZlWUC89iK/Th6kwo9Mk8=
`pragma protect end_protected
