// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K03dbU/yfL0ocU9ivqOliEZ4JiIxpNx9IX7qZ6iULIwV6SUfNjKJime7D6T8
Uk6GmgKivvFBQd+PYvO7B5jK+bSE8hKE6juYS6bOYOuck8u5yrgOFFrqvZ+W
QtINn2PZ6e6DpMw61TD+Vun/qGDfwewstg6dPqZm/gB23dBIK1C5VW3qUZxE
xvLTAj3DSVPx+F2fhU+79IQCnUJuoQGFhh2qqmyBwMk6q+bWHlwxYALGRamB
45q8uk+HPwnaiuG5OzD8CMGb/p0V0As/H3zMbcCHm5aEOzXThEGBvdDvLmn4
HRsaDAURPm8SKilyiU6hO11us7TCUAGpIUi5U9vuig==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S3MBRfqSIGhKRZC4dqIoPcUcHGnXiqCE43kCKmn+AtFr4FGkOfYo2IhBVGpj
ZfE5kFXcxCAhMwE9SW7VzwXYX68I5xkblDAgopG4/5UMiVl/lGOrBMn+7uzZ
Cqp5p9GutBX4R7bMkIE3u4r90PN5HGsx0+NHiE/lGwp5lHNp6RAfYoGkm2WD
YGAKeNcSsUVDKefIs7tnOrYh9Bp4JdVxl6sKEezbeMOFka6vA6QnAsYmlxfw
NzzoYB5U+j5njZOQuFHO+JLXEXVoHy4HUH17qnsL5x+x/rL/sAMsr/JUXHUW
X/8j90GcYR1S9X+tWJevY27iDqdlIaW3fHiVIJ9kyw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S0hvmtiB+0YmEzHTXQT/tWLiMUMyD9P365UED9VnsR+QI0L/TmmyH/JllhNu
Yh+jwhjsUZ3jLwSge+Sa8xn4cky/dNzJmgXaW/MRY7rnOzYvYxfboXdWJi3a
Bo/0Lz0lZiqkmxFKzksiQL/qo7k8HG2ZmMSNCHT8khx4Ikpgbu1pTYCSm5Uy
DsYh5ExaIFa2nJF2qKHgFBkXmFFZz87Z3LfXVRJDylCbEw00qNXjppLd/ea0
SikevbbiPs5ZLVS2P6x9AMwKBdU1AyhUxeo98a7XjFvtYD6pRK6aF/ym5N10
0cQ09pXkxRydql2XJDuiyCBXydfNha2dWvNL+WqUmA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DSIyaflQF2+PdYbCEptqG37VGrb5RjaA8L2sqo2UOfNztSHOrV03A6lraOXL
xAcU1OzZNnRjQWfAVTxUgTr4ZG3Ydj/5Qv8Ov0D+UYCmgd12AM6lcUKA2UzR
cL0Eri9b+8pdTDMsklPG1k2uBsh/KGgNtwl4pJIk4yZhJJ+JG9M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LZLyxgoHIVfLEGXFUUGOQEshGJILis+qGwFINIk7Q8K5hlggMWz5tGRIn2Z/
8zETYxLee/kEWs8k3Iq2tFah+MII7vEFeMHen+eUoGd0l0y123avjzdrWWVP
cQlBJFr20xQ3RPhDmVe8PesBCF/HLEsZ/KG2fhIFcPmtMS8nFtQwBJ74xewK
ZluezYN8HzOHyokVHTXTp9y2LI4Ab4R3XbxRuKmCn0TWP88dADegVZLLsMH5
HYdInEizlJDRnfMZgbU2YLDRXC/IkwhRhKJfRSqRcYrKnL9Lh0qeMWEqAvXZ
xz4LIVm+osTqUk3VITewWPcM9gKW0fGtPTEO94DZkwQvzo6scticpDyamu3I
pz3dfgkIwiD7bDZufu56UuxT8TbLKIA0h/S05a+Hrg97+mtpgVRUdbJiJU48
cIy3tCeZLXY0s8/grLVteXsCI3k9njuciTfgxy+lVn7ul+psGtUFhIGP1XuB
g+YPfFjlxfZn5hYTQKRNFM7SVlDDsPt/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eODxDt10aop5nMp/jy9MZoiZew91NfD34cAMkXyJEJOI7exd9vQfFU9+MfPd
Lii8tK//ukQ6km/WUvEeuTgwrTDp8bFOQ49q4+gqDQdX6m24+ttf3nqGsrJQ
sR/Wyh5tRYhYk2bs9UqBDXIKMkmDn0w7SDAl0MIZZYea5k0saes=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oJOMWBVHXj2SvGDXG7ZY9HT2wJr3+zBDBD1yl2K+QkPlN9dZGNFuKy/ZFPBE
mPkWedkFwTD//fvhk2EGzySxgMWLWD4zcHH/MTVEy13jc3GxJlOD1TqHJym1
Uy0l5EY1CeYkvQNeph11ibMnvCTGsMoJCXslC27YS9UNFdv1nyI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 642064)
`pragma protect data_block
/tyL8FDy/RNSWlcXrvHgH5hxpdSurgdKNBaTz4+o/9YHJtL/KwXpUQ8vAAwL
2VPR4ibyeIZOJzQegJs8zypd4MqjP1UdQIachRu/ThMp7sj4W78L1vfa8N2+
/p4E7H/zglckZ6KTzHdN6oul7SCeeS1XyX/Qi2a1hntl7HNA7fwKR38K9Tny
begvV0sI/fMh8hVnr9ieP40yg6IPBGMO+WlKFulQ214Mh+mYRezKEQ+3MVEG
+mKtCkPpFmFdnR4Y9NN4OJ1pesl/ownGwOGCBFJgPKRhxwx6srsmtZtUmzNY
ARi/ei7rVK9d45/yMN5mIP5iM+I8uG5jFZj8eQYS74M2kFn9xavN9og2Qs0U
s+LLcowuT7AC85vyNWol8erPC1HpqxxUVT0lEj8gaxaPoR9L+eh+9T0eZ5R6
HfnwziifRcXZkbtOn3GeWNesiXrRzEzu2hN6S5BzD9YPeI6Fp6l5KDcXOLO9
q8qPz1B2pPNLoHpYl+ob+dPYi2AXvvXTYCdi50Z2uE7Fig4M+7XPUu7ZuUzl
fQzkmfnkmCxXpXRQBQyJQfH6zbBuOZz2AmPPTFbgHtMZOb+8boojH5wJNKJS
6GedwpAWl3+XHAuJrbDP3utYIvpIELLGKUC4rAq0JQaxmkW3RAwMIlDd0SE+
qlkDhFVEGxo6eqzzm5CSrOMB+K17MM5resAv35QhMk91fSlhMFkfncSk7kpQ
QCmhKjTNdfcnmbGvFZq5j3agBQXAnJ72kugX0Q2UXpVOaP0/xR9idBearhM1
9SKybpewrfuncZyTORwhrq+DJBFtSR1V/Gf+uP9uSsgzw6Zas9Qe0PLNY8V3
aeZEVEjThNsoYVPe1WRLOeLq347c0+Id672GdVmqvRp+5gxn/M1AXdCcgUAV
m+9xoTjPoDqCKJbcOCdhlxStl7SttBT7S4TEksH31LBh9x0XBPm/eQlUmJBo
d2xl+hit7QA1XsbwSMJA3JOMibvmUC3kYZdVxD8+Y/uGWbLOfRi2AfmiiczG
2Ni8jLiUALGHTyl3TLzSlny2gfR0cPJZeojfTUQzyIK25h8R4g0jpLjDZkbI
YRRxsFDbmtj4PgRllkc6RvRW+CneUBnZ1wyrEZuwap8iRtLKVHR7HR17dsl+
fqk2XxaKiVH6HL/xTcODRJ8lUceKImUbwDC8x6kW+YkTVuCUwhJ29Rg+M6vU
M5JouTD3dQ9uW5bVDibs+92bL4Plbe1wYCrRUHJt0KfwjySXGcPueGxH8mub
3pwOTjloPppo/nLE4LbX2U6e0ZUbbXJookUeFCltFEWDAlcSQ61I1BmCgSCw
UTxxEqjiSsU5WjeFsDeH4NwlmB34Wrv0hpmV0D0H6W8grOxe5zzgWOd7qBvt
RAIyvojFtGho8xZoDBAp0o4v3BJcW7OOVGhvpN638DDzFBTTjm03p/UTAcpv
fGkfkYOJRHA63DgW7ahNcjhfE+RNBxV4d0HdTkefBooBO9Hz+ofUBQFP4vdq
D4cUbLJZsIJazYlJzz2ApOuDfLzwpja2G1/FsNKTNxLvj/ET16pkAOe7NWfK
5k1bu8+UVNpPIxOi1catWk3wwU7XKwHoiyU0NpTOQ8fiNAYzMvrkqG57KISn
1fLxckX+LbuPvZQzQbfV8Jt1EMY5bj4lAoUt+B/y0F2hZxJ9Wbh+NWMkMgBd
983KT+cMlY7aZDF9gi+YgOoSnfy57aJYEfkVImBwyvIwMkjlA2YoFUI6XXQB
KDLOvjVqLVVBxeUbOwHg8sG5AN7Fj7fdDXrlrT8ASo7WBZ4Zm71Zo6lNrd8Z
oFXeE50RbkKLbPVF9ujRK8f7Eqyoi6ViiNOnswQzlPc0LV/BI8ybHW+Jkgsz
gEvDHK0wqRkC6kmpz8AD7lK7xzlD+NZOP5CgDCnSAlVCFcRLRsRJhCpcIYBy
OwzA1BVbl/07i+Mfymy+PfAj1935xfvQ//RpzZ+VHN6AM+FuMRAx6rwTdB/d
BYzyfWo0wGkWQtdBWSqykFwR/P2pkEf+uTy1s8L0YKjFxofuI/vBALInIpIi
vIcO58XSy5PV7CGBepSrcDIqTIt+AaBbggftK45njGG93E1Llp+yRjVo3Q6W
C38ZvXHJLuTxsTJiqJpbgr0TwL7Vg6yIxhn0qGN8CVLacxhlJbYdtB7NO5mA
x5BALwmlw57S7Dgd25QVOlA2X+DbcREsynbLT0s97SD092+I0yLdqI1aU2lk
CYzOcfpmlAC/fno7ICS7BSISMTRCUZ3jlrcminkbF4IMj4B0nfmBbI4OkinX
NcgXdChzHBPrUwsZvMoR74PGrwukoAtb/kCkj80gDhwjelHxEGsEaOtPfhLW
esDn/DmXYFb3mZwpGynsQzx7+PUzO0r40aOGBLukk4V1WztGqohvsbUBq8Ns
234IVebzUfHn9QWz6hEGuuvHZlanXz2GtGsiWKMgWohHaPa+p9noP+Ili4hF
4pVje6XZyRLhENcOWMQu0LdkJ4F3KaKzulmOwWQ763LUZb8ahHxEQwuufQQy
+ituXE2Rqow2W6WnZoBU5V8zbQG4S68AhDlOKrIjbCM8LUshBIofDF+ikh9P
JCHQ5vz2lqdgEajkWBzrEVTRsdF598v+6jrR/4bi207K5Wq7RdwaZ8xRjD3X
aZ3S1GpmhTTM0xcvKjrz104Ffz/J0mRrObcLJ2nMTDEj1rmj/4O50skf0mFa
AT+eVWdvPneDEYE5zD1Gwiu5xAfObm2+EKx/5FBsEAVkfH9uYBwH1jYo1cfn
jA1XIinNwUN/Tl+bLC736erWXT2FggCTBoJt5SHpAd8abPhi6cSLJlcEXnb2
zh6+enwIXhhDYLIZm3ax1l4dzx8yF8JYL26WPJUVDgwrbK8l0UMkEQgvjkBZ
2K1fLl5lO1oXtM3Tgys/xtR9xLI06EvHKpUoU3K1rqXN9JwNskfHhKxKY4DG
AQSVKiSp1XsmZxFGYH4JYvUe479FGicrbbacTEWizMsIZk4/tAZcjFOj+viC
DWnara5iJ+7mUxvCgAVJO3i5U8MnQIwFC5Hy+gN6HZa20aA8YE7ZKnFPGoRf
xEUWO1Xm7y5ltTo88xyRSuqgiC7vt2Ym+i/unuhud+ffsQVECT6DVfZKrGHH
lDUzxejHdWdhnu4E62QJ6iw9gqBM1/+QdYAvOB6RYWsdFupiuEmYcIqH2j58
P2JPUiI7J73sGruO/vjUhxb6Pm/tT/hRVl1fubaCCmPd9mVAmNwxlaCREbSu
vpnJG6TGC9JM+hTNldA+q7dRPbHU0L2jezbgq1TU4v9fHZKAMsXq+jOVnnPr
ftDmFbwdzofvz77wY6c1DPx+r+BZabx4ik+N+M/Irvjf/l/JZk051/2bbXfM
H/W5cpiP9A21Tp7D542HgjLf52AGHgaqf9/q4YDX+/f3Nkkyhzu3dZVMl1E/
qgINJ0C4v85r/Uz00qYQsrD1PngwAhgSngW6uuyIKnoKtynh4oUDECrWPUm4
NxxMQer+YG+Yx3xAC19OA0t6phXmQEKK/tGKQXwrL+oYifntNjNysfUMDTO/
2ZLTkfPm4+II55QmcRXM2GG1NDcKkzJUw6vLf4cQ1Csc/XNHbdypx7BPjkBk
Bgq7c6kr7z+Ej4G/9EtI5aFr/QA8vkOcpyM7IlqdKNMKHyc5c47y6lAaQ2UQ
Qs22e9qP0cJxw97Fn9hR0+28eW9oU4naAYmaOAod3J10BC2AJ1SjBjno2dMd
mcxJpN1xiwIJ5hqEeu+zKSrM/kaoEn2OUxpKFza18sM7Y2DSi9njRvaz5xk9
OLFFQVakhRlFuyTX97CSij7Zn+Z0aqiodNdIcjPK4N1iQsAjDDBWHWgwLBFZ
PCRhu+J+LFMcV53m9nrTFcZ4vbRpIA2P5jWl5cd8UjFRSgbqnc9+fymb8HEy
oVPapEq5HGGIP5u5mop6YBy3eShFCAiCw2y9RdWDdVDMkHScZjJADG+hznnU
eMwEj8/1A55ioFO1yDtjM18iaskjSqraofKAilgMXABqBHs1OOem4SAd22o0
J54AVm+/u/wHeNaD+rUV/tgJYBVnmQKhaLX4E4yOIukV5KtwDN+nEv1iB9Cm
aHJs3RKJ6PSIShv4wbtuzmEOdZ0vxQQ8jKLAJqKFI5Eq9t+Qmb+zIUdGhl2z
Pcn0LvX73D3Hy7DrJxcNUV1igI9q52J/CawuSLYJEZt/UMQ4p+oDJJQpcKbq
MSeREZIgEJGHstb/AdyTDHtrHkEgCo31l5oXTCNgypFX/edNVwz7tKHoNrmF
/PCBKAmKKQEbxR9Gio6ET2fbTWzwB/yGQEK1KOaQmry/hid8SV5T9k/twzhZ
tspLkMDOlGQocGkcjQnk/xw/yX2LQi0ZqDSZJEPmKBMnZ8ecas7DZaULIRX2
Di7tKZzxGzS6ixvRE8DEl091E06xty9q1OerR4VwgMJkIB9ZIWpNciIgcyW1
vKaR9HzP2T65cnTCRpful1ViaY4lyRlR5IxmIpy0J9UUCTGFkyilb3QriI99
4GKGcZhi7vu/0iqy+6ugz/ACF9ak31vYWyTbReRBsxWvWStTJ/7DauGKOqzY
k0yjHklaUYBHgaapAnFfllcpRIEs+PBXbYUru9ETY5nuT4JgRGHUI6YdudZ/
nlBSCo5Rl58TbrlmoRiaU87veiH8br2zckUvIoFLxh3GlEkvz9s661xA5wmy
79PJYbWNXNkiqnHp13G9qMuD/nTNAIROY3VQYbI74NzdsqVN03b8M0HmO8I9
zeFB08r3QRsx6FJItHBiUljI4CmBhQrNOkHaxtlxd0YJHTZwtUynHACADfAN
4h6LqYyAwBXWr+RWtMkk4MBTpGjEaeS4TgzLdey4DAu7UCoto2/FFZ7CGOzN
44GIh0regqbU5SdsZouyht3m8+CQCAD0SPEZJqRGooyZdiXPqt42xk81hCe7
ipj8gdS030F8eNodOeWdnK5rL5k8PoSAx5+jhIGo2crK2ImfvUGdzbE5pI+5
1yiKq82fxg+5aonXXw3ULQO8tozl4CykRusvLanMRK/D49E41MX8WcY0XkA7
dzk94QmOFhm/YkSRcTfODNJD+CnLgMxw5MgYiazDPH8U5LOX2sPCmTW34Qsk
ObncWCHHCtL8s/TCroVk57xNCmK3PQ2UDioRoDAlRgW0X5FKN4cBAjCXUI1X
h98bH2Z2uHluhHg6nAYBPpmYyNOl9+UhMAj3Iw1VGsRzbk62BUcnuX2QneV0
QEYEQFis6YlqS8Y7rJ5s+EhsjGcb0wuhCXrQoBMWSths/SINuIQMCyKX6cuZ
pwdM4fkX1BNPttSlh2LB4jaSmxEClkYTrGA4vLAwwCHpe7V252HSupIPOB6N
f4ZIPSldyIuqk3QYp/p/tJoCfeAGobdkgVrbRSNT3MOO2Ky08WUHKulIRYPw
bsARo8QueeyGrim4JXyDBU8TnI0BnUxLAM2mtuRSyZ851tdDbkAMQ1q2kjl4
bsKANBjpressRG3kAGUCB4/ao5NzfaJ71kfXJu4lM4qa6xSKjWVb5i+hRL/r
+qPPwrsjB+yBs8I6INyOFP3O+4j7l+wz7DOI9f2ttWLfEFDcw19YtY1zGPLi
KQ2TYwF92xbym7nBOF13AFGocGtveWhP9qoPcFfijpa1sMtDeD6owQS0bYRE
uBz24tS8K7hCxfU4epgVbUQF3YFGCwbwGN427LXqMJIV1VtZWIJZXKQ+Q63O
UQA2qm3PNF/tQDmhYon6uK2J19O4k8XjT6nemYb5OrDzil9vhCBOHtCwMNda
T8DqqD0aPGaKcB06yzuyDY8ilPHgTC7urK1gI1KswMn5lBl/AxofRucCFshk
PX4NK+uZFWq7mxyskRJ0+3Ll4Q1yIBzh+6moLPiWXDPx78CqDSVVMtLiElD/
YNx4dPq8uHRGntCcQdLCN987nlxEIROcdphOWihQp5pM3zrkmGLscos+N0ca
O+0sXQZ0Ix7i9Qq3K/EGJvufgDdrzM3JSntLL1fKYNwS1TNDSB1aZLBUz9VN
LpnVL0xr/5fmrvy5mIHvDthrS+7sExat370mR353ySW6reMxwewb9crDzhbm
HE2RM9aPww/R56jJrDk2U9IklUbmB+254PHhZIl1I+jnB2HyUgufVV2Pckw5
xepu3EQAo+U0n3G16r/5gy5B8hGZSWccWT81Vl+Vc92jRwtca0svoIQRLzaW
Dub8eS3VQHbrlMi2gD6FZfcrm+EciD1SwnvDbuHihHEGebKQwk33Shg8X5xG
Uis/WnkhGRYkG+hJQodZP5ef/3LWbWfhy6YU5Gyqt0EKh7Jd4Nu6qY3THrqj
/ISrb808dpv+9EOA2PZzIpHHkG5o2z2nL9cUL6wVPHmprGreB5uiDpMLDUTX
SeBSpiLLXR51u0NL7fRL8A/bq1er5XlI3XSc6dzzvkDUxw2aV6hw0dEsGmwK
FaC64Jg5aIdsIXzpJA3mAWGh0WpEIvk1KcXtp57F9/GRFmxZEpJlB6quvN3q
e0ekcke7DokibRDs6OoERsIHjrdLn/+Ir/btKIY63ebFCrYXfluCN9GAGHOZ
wTB2PJhO+psK2+7FZoRFgf1iewTr2/kF4Cm9H76xV0BBWZPt1xE2sg19g+En
7B8IaVSCfrvNJQBJg8DO3PTVPzKNq5zlfn8jXBE9kYTe4FNX+plxtn2JE4i6
7Evt12Jcoh+VxZF9KYn3OTORPzVrW5wrMS4mKmhEc+AMwwuiA7cy28R5Q7o4
VP0AivjFQVP962kv2TgmsVohpQ4BMs4Q9lj81eozRyEbyGma3eq/aVdqXW8w
d18vKvOwPWXXK+jNPGld6kSMAGX7XOblWi3+NJ1MtMhIUCJUWNFpw4qXq4IB
0G5QTB25Jnw0Y04bTDy59pOiZ9hRFaobQ1tMpChXXDFUr9/48mm5ADmRx9hj
jsE3imM70fujLnuOYe7mSfSYmavcA0ZNjh4vub/fAA98zzrs9DnEE9XcEuFP
tAha1WHOs/0ml9P/e5h/YF6oiMc2mgiotGs7+9k3/pye4yO9HTniI77qmW9N
Q1RM6HvI7UgTltJTd8DLCuNvefXrcC8h7ydyPE5kVYpZR89ZQDDNovPK1RC2
/a1z8v7Dp2/rpZQHRVNOwgeClAXIVAzeHvB6z1Eyw7MQIa3edehUA8q40HSj
z/YuoZNxDdIB0USxtYws3K7NWfOcUX9cW7Bmu6PFWcmw51eH55ug7jmV32BQ
W+F88Sxb3/XrsAzSR8cztVpiv5KFQEtjovM8S4rvp6/ZJLsY30D+fqc2xagT
TrmDnaNSvCAOarORPfLXiT6WHqpsZVFbC9CmMkDY6dAuPaktGjafnlqOPPJU
CP32wBdIYdJTJo+Bg9m9qvKDOZjUIifRvlWKqGNuepPW73TV+1TMkkKKCXe8
Mr0d+69cXXHcxspoHuzAqMS3VR+sbADzaecTwVuvYjKmbWNwl4MIoNYr8EjQ
qg2NLUp7q6D+1KmS/tQrKALllXxuwhQD7u8boxlubZqVpVFT4z/tRneYj6VE
hsEsmp2hWM3N0I3lyORx//v2bDwr9BErJPbNCIpXUFQUG76u3ZKjNwTu86mA
n23h1eR6y5AsIAkBLU9VhSRmkoqtaGkH3b3a1JoM92NyY/Ov6WOoNXD0VhY9
hyF+ovsv2OfC/Juw/Od2rl8sVnIERPcqvvRDE6P+1sRFcFjYJYM8S5hNOpbn
+UkJ74RCqdGnwinGJFqNPZem/VxKYH6dxcqEigH0w/9nCBc7yJkdG/DgA3lM
U28mugsvobhaE+08RmznuGgC6Ty/ZI1gu4LzPvUDfquwAIOwV3RAvl+JNYzO
UvE82oueFujKYBkiw3jfdzElQP9mUGZdPSKaJzRI7CsZVirINR9az0I5+7ad
IdJWfvn5OE0EEVssDGJLRmL248PniYNq/hp13eiUYoGMWadoY5495Ke1Ck6q
803sIR15+BpW61WbcUagYssN7GqZsVyvj9Qe1VDr91O4br1PUchBoMdwhjfK
9wd0TQHjvhggRVQtWUSvZmiCEa6famxLMsZuhRX/7YkZwXnP2UsCXAS/BhYX
I02s0dWWCp/AhXQ2v/tMaSgSlgc1yPULiKrmKK2PsAyFKWA5RcxadW2PFMMr
861Pd4Pnf8+7aZOYfpGI//FMWUnFIIruSMV2mrFk9NvBbjtMwbnCwDW5zD8L
fg0DxivH+XEfffGykuXah6GmIhXB05h7gptIaW/owyUtDT7gWbkT2sPJrt4m
g0ZTaTSOHFm7qterBVYy08T5FpT9TG6uzC7mVEKp1DaUVwW58sJSxLkDXKe2
MG7QnZQSaqnBi0R2/m6AQviVE2zg/Q/cUF6lzCBuJS+5VGXvrUokSEFOQjIj
wDH63TmGLGvlECiptbcZ5FzTSDDp9qTss8uGt14SNtVO+QLc/wbNGdM9IMN/
76/Wfl1NqbKh3sxZfCOa7YO4wiJgdMrHC7Ph4uYQO5kJ/KIomIV73MtiECF/
LJpURlyZSynsSt5bv/dd7YOQILOXmhG9vr3ggFz8c7gv/TXteW0kWRKT65ul
LJMe2BBhf9AupLxVSBqxjFey845p5Lq989T1rUP+GUA8ny8JYfUycaJXL7zE
9Z1V+kMI5ClXW3qKOdYuYIBFNhIlALZxe+PAnuoR65FtfePANgEXR1zTBbR5
keVvBXBO2+J4wuKDtdmej02G8cT+diHlLBID5iQSNrI3Zq1qS9G5vZhkDesZ
nCzhgA9ht6W4kH5oqKN9UHXtfLL40Nh3RHKiHyAe61iD4p8YPQBbB+m3kW9n
UWGXCeesg+vKkjwWwPvNO2FZAyRtqPKAQxfupVtFjrtCCnQrBIDqguJDxyka
lqaXN8zo4qo6VQZbOnDgjfAl0cv8YXSW5ruxhnJPsYLUGpCBj/kR+BXuATup
Z5lJvS8z3UVR2muuIqv5R4+qHnPpxhkZjVIXBebQ5cfGTk9YGTPl1GnkbLGg
plNfB0nfavlbqbE18aFGlpxt6IsbkLYp4L3dEfZB+NXNNT9wq0Le1JIBHYyu
mEgmSKbYWz1AOH4vbSDxYsikXwbpqPkonI5eIwnQ1/9BrtmwQMyDwuRtP1P9
Y/Sr3Vieo743tEDkHIkLtTgIdR6I5HE4ljJ0BI2WMR9LZ4m5pociKhe+Y+Nn
kAeG7hL2o/8glHAghEPuOQqAYdU0XZaTYcR3xg/7P0oV2/ZB+LZhuXZ6FkKv
FdN4JQ0QvAOq9ZNODf6osfc1l/6YKpdynQeHZbjppTtHrjkrqIB3XW1Jta//
ow4Fk+p0APPAKW/NQITGROGMmudOUXsESgdpSXrpvxWyYva3pN7JmY7S13cf
+YAjjz5BbZ8iOjFr4VrCPqI6IMHBI5GKwqeG67vJCT7lzMaNBj7aeMmw4rHf
0bXexSCH8mxXoJ7VLzXFWwg/+/Phrddzq9TCa0e4SmM5QOD66Uj8/sQgyjdX
nz87RDnS/4ruvGu5kfu9EVR9tnr3RDYy1tNyOlJWSYvkXT2HwuDfbJ8SFBPd
gm5/tK4m+4lXnnspYZBNIeYPypERz0ejhwjdmEfGwAl1o1VugxfIxe9dz4By
IL/3K7m0p7cpgQQkG6bGURSzT9NFQnaxnI+BjXbwSAhUwpveqQy6sfVktxQT
/EEu6O7QJuGvdOKKo5OcM+iRpakC+zbxH4zOzX2bVX3JnfXVSC1HjXCsw4FN
keGkPNlrkvS30S/R1Xf1V4urKKjU+DK+pngGRRKryNkKRvZyVbYkcsIHFl3j
ADQ6R7PeXlW6z/mqUlVPsBvjkhLOHlCnjT6Kc2cIY8hcW44fitkZmtpRgcPv
M9GnX2m0JH+wkL9zKOBuqBTpXKCmmVfRCOcBqxdrEzggP3wSxuRSM1XJkcGx
fQFQE2UdIvv34SF5mzjSvgGCYg7KYPUueCVmzJDXplQyqIBix2I7p5DW0r/5
aAzROmtObQ7m4LNK+hlxtwo55roufySTvs0BRErP5Hxv38Un/uqxmFULL7h8
EkoTCQsxJ+gaJI/FcBSjTiKofOuRhuxahP77BM46CwyWfMRoaWbl/5HOh/Bi
fV8O6DzK1tp+O2zRBzZERozC422k5sUMtBpmsFmLuM0D6rI9pV0tE9F/cFXn
N93HExC8jLyVS47IjDITobRfZEutVdFjdJVjK6fKHQ4IVrUSTy8c6Vq5VTmO
yX1+u5UEz5q4yTjrQ4WTQwgLyqdXZ3uJO4w559prRDigfckZVyVUENUghApM
/5h9hUDFEx92/IjTKK/PlDg73NJ9aIZ/jayXLcu+586H0+C3C+37RKTO0TR7
6qzPjbhvVl6Yb4ESorahE62LPTXD1oe6LuLMbAa9hzpcHDFlj+AkVoFwHTgO
2AYEAl3fqYrKvpTk/ASUjLNN+qSBnE1BrMzDARGXlBl0GyKubGbUkYiQbEuZ
3uzHaI9l47tGEM9aq5yWk67Dmh3Skdh72l/J5t+zm9Q3vXbXflzHHPgld8k/
/toiHUeuvFMKVvXcrWO5pFQ8bksvWDz3yWqnpKxvWvDxxzNOaxDWfX0oyLix
QtXKIsFxrW4nJ+9FTUyVJAoODtNOp6vXXALrlhhXpi2vI1j5i98EDmsLSrIB
TpPSVTKc9G5b8IXwly9itwwsh/Ov3mbkNjIrI+0JzfKJW/ACgyyObqIXcAak
hXupqS+7pWeNNTwzBp+P14whpFDMcRN5oEgmp1UhqW/IGViVb4s4jmNoZK09
R0i/dF00igyY9T8+6j6Ea/TZXXoNvVZHWo1ckqsvpTMmYUmQBWwWaUbDtGBq
2bxxG/LVZPio4AreUY8blc/CZdPk/foKISsxZXY+qWyJ26pRpV8aGcAgZtsC
aJMAJWWOcaHS2xkfIQObj57V5EMwURJqqOMlpuxy5jIMnbjj07c6xNeDd4JF
6ntnmpWwkCmO4zFoeH78SuEj3GUvVUuQeynfeBMz2wNGcSrgF1XBKf0d/RZ6
rFt+BBqeZ5ggqpPrngNqvp0w9Iu801C/ZkfOyM+hOsYR1wOveKtJpW0zNJK8
j0ojjcdoZlFxxphe8z3b4GQJ/zWHC+2WI9sHqN5o9XwXJ18e7yz38LDDBKWb
j7+UbZ0HzQLVzYFHdMKCUbcxp3H3uo4MKcvMpd6UW011dokWtGMaU6t28nex
GW9DdoKIXaEKIKbP9MpIxELezHcm2R3srRxZ1QzVYRKEcj+kP27hVNPmRMLj
7+rCfVUNABFtaocoI/lSjg8udc93bN+9C01xO23A/M/KwfJ0ZTFgRyey8pBi
6PxLNVPL3tQJ4LaXj/Zw8fKboOfmaxgZE2g1y9P1OQRYTP8R+NRemThyxicU
pprXdL1Nz1KvQRuaNCgaK5WBOjHn0TYfRlEfXq3xLGJ9ZmashwSTcNYMf5E4
hDvpkof4uJcAAKi6XqN8Vxl6F1vI+NSrx2wNXFfMv+2Eg9a3qqL4/NjPF0fv
J/81Zc07XYiFRWTPW3td+L8/vn6gA176DFi+iokiuTdPs43BWvxTERPlxJIu
iNv3B8KH2xE+cRvh93MGkJ0BQKo32kBYVmFitDwLVWLm6Vkh3erGtwLA2dmW
Xyg39Op/WMqHoQ7j1mxm7r0zlNf0B0wPS2tRbKT2NKvb1OmHYukegULUgAce
1L09vlacJUZXSmqcgRuObjC6daryV0EDcLdlVf07mmENzjSgDEmsnZeJ2LEc
Aobka76cscXJtTqFwARMuVhOvtcJjow4IhgJ6bSZ+VsIkk8i0gWYVTZXad7d
q7eIp4O9jbgej3JPWmM6zxSBfj8114oArujq2SsaCbYb7Np9rgwIZOxmayo3
uSk4vAvxGUQRc6vkKxbP+1s15japgHPxGGYnVh7fFoCmhF4yZvmak/dhbX6u
dfd14V/dvKsOp8kWkiwbTrsnN9APqKy4k4Z2UaUzYqcxb03bR54JiZv+2gwq
4vB0aahqO2sq3P35ZLdkQ4ooBMiTrMKxqW+MjRaKsBuVqO3Bvm/XF1Gs8Q0s
V36PWH4kqktvYHD0ue3KwF9UI6F9gMGNrSrZZDVNJksWTOf9UHHrUPD8um9E
2wdaHbnZa1oAyi2498NJtQGA+ThNjYbhTl6mkMnhOQxNp3GnFrVT7ZylxnKC
WMNOjmBLu9nfUMqfxrHqi2haz8R71fdrirS/r52TNglfCOkBCEqbAi5D6GOM
oxU+T4+BIhmyEC+YeM/5F7eQ8D+kbHxgF71NCzrK4LsfZK43hkLOYrRvswmI
eHUgiMDCjFRAnOs+VidxHVL5QvaR/Z9bWt4enT2cQqqhfOAx0PwE89ONYUVh
mapXV9NMUids8ZZbZbNFhR9jQSoEB+ohWI1eY9iOlRYrVycbwLmhYGyDRSlq
JBl29FXA3QtXH2f9KGscNEqxafXCPzqeniwmfigzQ2t/2u3wrc4ENmU11TlK
EaSnnfl2RtfLHiP6lS8WA1mffTxWl2yr5SMnGXrDllwFQftDQz8x/OZgrwE5
bUYfGe0jotHDBBZgyGhk0Wj1wctbd1UFjq0HkPfzcD2Jd75xD3GvM9yxrHqI
a7pQ8yD6xoKbEo0QR3A9wHUJE1UhfG1EtDQpnG40Uz7+o7d/XMbXqWFkqzz0
LaIKN8gcPOR4fXf5fREl/7zi8WaHHk2mBaiBM3RPjTAE9UaSY5JCEEc0wc+T
X5R+Cs278Frz9pKnpRDmrYns8hs7pvE9Q+1ZEkZHyiuqP+FvDDAn9GFmhPSs
qTV+AR7EELM2ba0WvxyYQT+bHiTQYd/Zo0Xc/pcu97gdSvhDDzk0qU5tUmyl
FJ6yAZp8FWXh+9Ghe8/1oqgC3NaIrVQFmy07xRVEsyiYAGxMtavlZtjHQaDc
O0uyezpxGTqmYU5AMkUH4WKnWEa7FSFCgy69N6VnA/fwqmV+5lKBJIpq1f+S
pxvMtf13xnVSsXnd0MsCy8pV4r5r/1W0EZb7T7UtiNUHflUXGINCemrBG4bT
NfmeUzjk40MSpsk3XieE0VrgOsPqu7do44DWLaHt/3GPg4XpyqB/oiJ6j2bm
kkI9JQYHW8pTkgD5GzC93q3gXbtQ/6y0NIc8HkM4n7K6VSBxqN/Ge+abez9X
DTpSNxjPi8QOTR5N4QOJULdq7pMyLO3+5ZMb1q7HF9sDNO0X8nOMwXQRaP7O
AJzZZA4UK6KYx2oDMRZo1FgQt5SszBt700Em2uC/6AAlMSgNZDVRsQ93NZWv
cT2lNuNWU4qyuKhYMrHsZBazTCblW3icIiMEkxb3C8cQu7o8ZsPaVHvQwbzz
SuCCo2e0JuSriBSu4L8UhiNb2yoi67eaofST/5JhCAZv9iLRyeJzqeIB0fUj
l8UnS+3QTp+qrg3vGjXyQdbb04v7pmzQU01ULWb7DVzRwgrSwLKc0ANXMswc
lLnWukVNWppvWxBbv46T+B+IgE9JotymSfB2X6bu/btmadAnflG3ZALELBVH
TwODjDy6jo5lM/NkqeFXqMCUPtEBH0KBD1EgrT3PaeTM9PPW9kiSoW1/2J13
dEixjIRBbkd2W+8HP/r3UIkja9tEzRL4PgTQwRpsnV29Vwt8/87kGXCV/k9q
odyT0gFAaudcs2SiibHuKSR4e0cc30mdxUoCR7BjEz7xrKZTdREqz6HnXy8Z
W/gkd31rjT5FtvN6AFD9MVxZ1GyAskaN2gg0Rqcs01MsP6j7qcGn5qByasR2
ochJ1xqSv6xmy6bjIzazmuOZGCCGk7NX/3Sa/M5VJ7i+HhLT/vZAa/Is6IsZ
o34qvIipCkAYmqeKGPhFkyWZ7+irSsQvGJUKAKOlloRsO74NZZFawI8uZJa6
JQiGOUh3hwPnf5uU5wwpdCYvov04q+DRT+MnOJiF9jO+yUDyTy8C61TOvk/k
v60uBlfiMfiF1mQmznpKXgxY2DYE58db0jmOOGS9q9I11zVJ3rniCw6awgv3
PCqZAO45FSOF0fc+INl8AnUDnnXYit8rX61SOVRCt038siq/6DDx2iu7u0ku
qlyzfJ2ZMZoGKDNqlkqu9tGTZiciss/J0QQ/OcLgHGC0YlZJaIIXb1JKIc4b
HO/TB5aL5m1dwPHTzsbTu9HMF4YBAlS6l3TUYL7BEhjyMBUCvSq2xNWiMPbp
Noek+vvpNowR7Sjaato0QyFRI6oaPY3zNkyKJ4QLv6zyckZM+kAfQUazcgTg
ZxBoKYtJx7nzDDmW6MHWLfBfRmEYT3JtZdwLmwkQEsOZ059hAlZEBfZJbBpD
XStp5RZR+1DvAwlbCn5wDsFPrjkkQNS3pZeEmRX65Bs20S8LC/VHhssnCrAi
P5UZm9GVOa6V8fhrjad85si1Hm6ymgBB7R0n9n69aGk5Mloe/483OfgLNikr
l4etYRu42/z6iZBZTK3cTLAJQQmJaq7933lQNXUOuDoN4SpcRKmkvj8589Oj
aU+Z3798RwoSOHkGgbUFGRBA1skEAlXUuVxJHHVewfGyKo/3QQa/JdZi1XxT
OkFOLatF53bJkn/BPSYrsd2So21lS5ioxGH9MqAXDscqtBrT1FtERk8aZXYk
O6FR4N6N7+YP8IB4wn+kLyseHdDESQIKugTmgC202BGM97tRBYcTSl7HTt9N
OuKOsqtHR9gaEEqiO7JRQtUQzbbsLlvtZrGa1ErlpG7mMWXX5K88JZ+BMZP7
K6TY0cMcxjbceLkiYrZ1J5sEZWw1wEBrcU14z7pIYGNM/ED125ZYBYvFHFg6
yQsf5Cixf9YtT29wRrGPpNwHV6bZcpiJEa+m1cQEEDNG+JBtPo1NF6MoNSYn
PEsmnE7uG7r2lY82QbBkhEOomW1FCh06KrKU/PTCrq3eXzVa+Zv+0xXxA180
9k6NebJqWHnQufaH2aK8A/MdKIaF07VDI5Eoe1TKMO9TzOGfV+RmYPyPWSYS
XnKWrJyQ2o6y4QcWWzhysQ5DmOEqQJDzOKODe31oNIdTbF3PPwcYwcjOORxw
V5dB7tCyUsRd5NPpFq1H5FeX17q9TqHvEKmQaeZhtfHNkmJT0wt8tk6lI4yC
/BtyYD2qLxq9AvELG2HQZT3Byut6/TxFi9uybCOBLM5zu+3y1awy0eky6NUi
WsszVqhV064BTnSchou69S8TjRKkGnEH70lbwMNzKQqW+kAi1RQw77yitwVc
2DlILqKwlSQI0XgEluhIma9EpJZnv2y6mGdlV8Uq0kl61VpGk++tl0McotHM
bVE3yQfIL/Jeoa7d2Qyw9hrlNnec+/7xGREUEviqGvU9GI1sM4J8GzFh936h
IAi7TsoyZQ2gvcbxt77CEqpTcsI5O/AqQfVhcOe+RfgMQ2OEFb4JFZZ3/Pq4
5TRiGrDIb42PqrdGsZsulbDAvbUoyJ+7hF+XxeY9HcziR/c08ltseCZcR+uX
vT/6GUEW6EawG5BoZ3gj5/5uwPnEiwecoGj9p7hr3yTLmsTaaCUC1gO3/NlF
/6v8im92WDXvUI++cAqvvv8KpT/18X3WTFCmUI0AuOUapeP8M0oY/x7mWAG5
eoS4w92hjbpnVWCl23iOyG9T0PnKCzYOA82diUxQ9X0M8PpYPxXluVZB5gss
6aakRRf3TtKOS5QxUAvzIlJDA7X3xsT25y14D6xd42imEP94PSk1pi52e96b
q4l4DGM+u/Ilz4a38/pUiAvj8vgXz9tXdYNEdC5zNeEAFOiRbc5sZw5B3LQ2
3Eu6lwe7deaVh00JBoo+5C1uusKQzsEJJBEiJxv1BWn0WAgyuiCPla7GDw4y
cccjgsEDzDfhwaAdbAgcYDOJtr5TdpKbriP5mQJQOukVYce5IgYdCYLkIpAF
8vIgxc1P8E94K3/rgfueGmEQjyEjbVbaQJCDOI6oA576q3SCxHdL21X54stQ
iiiN5u4OaRzJUSXpq2PEOnHZDC5hR5winD9XvuhAvzbRyxjS0dZty2pmhkak
E+WNEEEXKzaO9GEU282NVLWdLXUH/rdIKnP04aOVEsDzdCrwtyc+e0rYvrIK
ki+AO8OhGLrQIdwcRQdHsNWvbecFiclyngYN6W+fFAj/+tLt/tYlSTuRtTM4
l0rAaEK/Er2wsol2zORTc9Pj4DFGKJoAI9z8IP0Add7y6iK1b8euU/h+QbSr
UDiOFxZacoQv6bEKkO6icxVeqJtpmjMUOCA6u3IuQDrdy48lolbO8zMy7zuh
wW3bmkR/C26cBlcLvupz0YHCOtwnO9jx9B9VMc7sKF/wKzH0Ca5QZyR+EQzs
ESroZTq2tBM+v2rPNRRft2tQB+o7XGoUP3FsbMC5902GhzhbB4hw4CW3pO5R
+5rIfr4WnP3Bso/+7uty1bnnjltCrrYNNRVsv15ucrCWZaGMwgoNWGOcVRsK
IeNwkH5RaouCnG6rwcJ7qu1QH487RtZqJoJidrXWCI26KIbuzuogU/V7vyRM
acXfstso3Eg/K1TtfEgNCJSRyBl9rXk6xKR9ihd2AZ6kZFg8mN0ibq4+jtMg
eAQm+jTukl3tR3DCDwfKDL8xjajapUcuc0X/nBJGWPYsfQpacJYJshauVpyK
4S1tePmWhz5YIonoY/YiEZSBxi2SZBpQ+toJeo36Qt40DJ+vTY2hsTBFdEFj
CV3tNOj2WCBvei2T1vBfPcXz0/OZ5qrpjka5kLkoJuIwlVCSpnW/Sf3HfAeo
k/V+EBoYeVegeRioD9E69qZ/EDD3Qu0yrp2t9odShdShy63av4JLHgV+iS99
Z1xSos+ctZkhDd3fZw6G4xjMRgGTuez0qUXGO0U9VA7mEKPaKWcpLHmGYNEX
NqSDFSWojyTqmdBz8MIXqaU79gKi4WI1bv4XzP/9/zz0sD+TikTO9xxVzMpM
PRBWeuBTryNooD/XkKA2xhUJiB1jP+M99hfJXBLBA+NXkpmyEqTHh1abI7RJ
RUCud9p8o1tTTwtlXjoq0u770wN5XO9nQaNcCtlDzZ00H1D45wSeUMu5/0/k
PKKrznK26MeCc9zZF9CT7gx8MWqyK9289COHwz5svMN+3iaeYBAP5pk4jH0o
eS6tpC3PvvwIIeK/5MCEBqTbG0VjsomnsdwN+65PvWIAbvytQBxUUesVvFct
xmB//4AB5CE/pNupNJrL+oOEOY4ZyutMZQ6shInPMauJsioNXXUNCBenGcbF
23/dQQJpjN0AVA1qLr2k+HCjV99HKU41vgxWc2khImELLjg6nVeQjGUFTRwa
bM+WCFSAuGNJibES/W/Y4MwFXPkQw+2ljFHVtqE/OnFyYh8ZeigbkrQ5+qvB
ICuIzcy6d7PQvUBzX0PQst9ryun1MatothoItXC+5Cm8hpg8LTZoXrviltLd
yMg1dlFZAtFZvYQDmp/J58QKArAIRNgR5pg66RSs9/hJH2D7sB0wplj5/FbW
drv43FFLgxdpNESk6W1m7jqtUh5c5WVgQBlnpO1bsto+pbYvW6Mib6HI0/HU
jg84Ppq9Nr3iDpwfe8ga1Cd54FUTOzh9mzHquWHRfVuAP5blbXJAyA9sUqM+
DLzB+LckJgFntyWGpx0kH7RMco6jS/3w7nT94WW6WFsQXAaBY/c8m7iQak3d
dfDNZYhjz5QXH4SGhsGFbt0xXypwG/2PMSjrfK1uinNU1db9ZKSnCyLp3eD9
QnFcNdzmXEirA52YNPzHT2gtLBLyf2ne9b0sVYlyvOOP8SbAMedidW5fFERT
El4PlhVuwsr74o/FfCGrOPRGiapgcx2IHvfV8WnHeGGToObhDxel8S3lUr4+
BAAXgP510HKfp8wKARbd9brJza15fymP9lHzhPSUw9GyXEnRc2GsJayzLkF1
lz1rVO5Tk7B/joBA2EerCEn9oYsM9LwIVAg2ttNraAETVAGp6xewgcq+JjX1
inDQE0YEV165dzZz30ZmknrLFHHEH4+TbbFEvbcUy76nr6NJOhrLDeEX/6A4
or1XEu5fs02xg1hW/tX5V2VMdx2bnvVAUkqXOmXCoZWMaYuOkxWZqM4IhQyk
4t25DMX7bvVHhf1ryADOR2VK/yJS+0AC/zIH/k6sj85JFdapgXuehen5XjlL
5qkBzQbR5OcNy6iriLASqUvcdxy3qyHB4SbWhG1SoUX494oIwHqGkwVRXGr6
2RjF5lLYPnhEtvcbmLjJ64syi0d0i+cz2zIP+kHajPIVkXPDQRiN126kWpRE
BfCCW6zxyYbvefM6zEz3hBvqsEAQA37D/UzaLO6e/kFuMmptteplLGKg9nsf
Z0OGmbNMRSfwy1jI3xZQWVzpMWoo3ajjd+p3rEnw9IWSdzx+xkRZtQmkeDug
K4Yi3Ar5/vObLb7QkbNoGNuYaCZL8FXal6pqOTBWcmZZ7GGFI3L4NZI6/6KE
KNobntAwraeHOedGDuxdriLLuntJ5qJ2Y4Diix9VXeYXTCacIi7WcZ6+kJZA
dP52mbIl5fyb+5TJyTJcoxUJ0cOKV/tHY5a1Bk5IkSuQuYbJ06rfdCRbNEvf
hg2U6JTRWA1bZTbPsA2iPlyhx3h0MkoIBzxPrtsvoPkEIGJOwpMndT3yoW7b
HOSdhGU5nd7c0HgUg0HAaLOge2fewM55mYnfp1HYxMaSBBRGQVOy+90HvDL+
d+PCGCtk2ZtRYwGtqZeXZSf51h7XYx1RN3/Gbkanje7/2UPsxyQpewDEw54G
BcId0GppSX8IERavsi4fuoHFbcI8zOvwqHAfKd87VY0/svyVRr58SWPeRsVU
nOlGqUjYa7eWsHI3PFSwtM3Zvnv2T2BO8BACwIYO0VTh5Dkxa4ceb/Zl0R3/
5JehME1/xySeFdvyycmUGeql1CFQESRLiQQfTdCd/+of0FdHTtnb8Q2XiVYp
xeFeu3YDDSA+r8xethEsfvRy9GQvnaMd7iXyVF9qRpVPFeKxKrlPJPZjeVuQ
DixKzhHRjb5ikUDm2IDWE/SLOmHs6hqC/LnTdvtBty4iOKdMnRXHVfSU50G+
rbi+clDiVw2bfjMHKdVT8x1veHi6eC2HXeDErRhox6MWMc6Cx2OlTTv+6gJo
QsSBRDL+UYoOP5AzGVjXDXLQduEZTjGDnleGOjqWchheUWOiznH4JHWU786Y
QAhrytE0HPjIrJKWTrmEKsN91tREHB6RNlYgZR/qrUibOOKvMMKe4iBwpNTk
fSQmoHy6pxRbtj11z+wh3hVuGCJSCQZes3Hk8VGuCNYQdimINySHaHp5gtYW
sbZilXa6BJ3sTc0xvgLffeFVnb1+b+OeYJTKAxnAGG/NVjXBJDWLugMbt7Zn
xgY/4qLmKak6hVXWNzw5HFCT1oP3eNO0EyrPUintofAEQmSldK7XChZCCRUv
Ejb4ukSW3nskGnjMJ/Qere7Yx3cp2YhO+a9qP7WHLPYsqykGV5MkOZ9I0/cc
fJ0MD9aoxyj73Atr4TvfqxNk09jax9cftzp5ArpPAt6UXbfuzdFEusa6P42Z
z4zXyAuIuOgoYbCgBbTMjMVN1vqQSAyPqMC1Qf3Q/p4s8Sa5M0aHX/1SeFV5
BOTGfeCtopclXu+IDdIqWHTL8YenMfPYA9S3W/hqAG8bqzZO8xghbZOARt9b
ZG1QwF0f4aYFZ+6/+Kc/nXyvSWTzKk4V0tBH9qJbprhyca34fQdwiDldrpM+
f9eVdeyW9oHXhuPqPZKqiA7oXsz20xbKa3I+7hFnWLhharYuwje7zf/1y7xs
NrAXXXNuefIou3Dd/YhRM6if/o9bNfzMIgrOEGo1dWcHum6WhPfFuHSqaEWR
PIulEsxnCyvSxijh2ANAXPV54vnGnV4YZNM6YKVQyLSI08i0McLFTj4nBlKq
OV+HeKpYjN6Tfr3BBnHXq3qk1kbXtHAB0eEQ7i3phRac8EdW28rYLJacUkVX
Cb/LxjJ7J3To4L3z2VV4vkbPGDRsOJp760B3BFzIcsT51eHBFVv46oFoa29y
tmQusrr5GzPC9RwHjxNKYyZE5N8An5RT1CK93XCLOArAEOYsuxPF73wxK+jB
3itFCTV2az99vXmfG7W98+0E7wILLGVwci2jgrjTXbAob4QIHjLJGjoXaTVg
1J4nV6wVBAsgSXQdFebYE0MQDw0O/nSthyq+BYyxdSxACPImJzeFMJ8iWTry
iTdPhn7JN9V35ZXl8XBJMr7RJM1xgXjL4frIVi2zz/4FTH1jemFGU8SXG0J9
oxjgCevgyMYhqBvuOm46CdtPTD6bPxXy270MIxsfP6sGZIOiocEYGUv6u5I+
Ftxw6CfO1jjT0mfiDYCDdKT95lwOXX+b0fvhvYNuRHNbLCgX7bTwesAYOTEv
M3AbXe1UggO41h6JDMwNNqe9ao1voXJVlBVtqBpevUwZB9uPFKHpONfYXp19
pA6skWehc1/7NKGV9uX/37TSZYSjfITBMrBABjx15j3Thxfd6+f+MrvtzMQh
jBhpkYxJvEkWQyjBC1yWgAMMbW+uFpdug3lUW3KU0uDY34PyxOdadiGUvs3P
TGUeoO8zW0thMbJ4wk4OhnuTMj1jaoA6eXpu1KJBNT9ne2Ls763q4bqiWxFc
VbCHQaX8bcCAWpILeV+PGZs/EjGqjr+47QqMmpTxU3BM75gZKaNKa4I/A38T
46IwiGK64JF+xrrwf52fX0kfg9ZhXFt2Rbdt3+7onFJOCcfV4e7GhrgGop5a
rSO81ErS9N/K9Pd5FxXbetCNY01T+78byDTIwrvugEW1rk1ZCS9Ci+1LU55c
Prd0+uPOaOZzAKt93Nsfi2YziSp1fB5tuuJ2ODwehn5ka830OSoZZYmJ8Dtj
nd7IoDRCKHsQ2aMDM9MXzvw7o6g1LuvX8RYqr9tGaI01V6jKenkf0eL8Tw/l
EOSzEDwKYM7TOdpn++Sd26+dTjtQiihX8TgpwRZ5NBAmutQsVwd37+kvFC3I
drDZluLOEG0+XofxBBpVVcjJhg/Nji4BiawCoRvzCaxD6w514QbjVychYHZH
vAeUDCE3cmHpy+Wz+9oYM6zIRBkRJRqBwQJyPRuai5wolnCoVhyLmNXxdhEX
jGhAPgiqh5mUGN78AMoqtTXbT0RwNYrwaqEHa7kqJLWFLY4XEqiKfSfO54L2
W0tN+nvvKhxQOA/pPaUkA9AurVlJAxd/D6kjVUgzJmONDSGpw0RoPon1BKks
cW/tLFofpYmZsdgjKi/KtBYiNtvUbNyL+XstCASde3ux0CoVW0gZ+XZjtmxz
KZ5ojsb0F8Iv3/EkcDYM1kW/9DoMc1sxiEe/z9c1lgPwl3ib9V0Kpy359zfc
sLtjVnZMvbnC3aDWH+f2HC0ymCMdGSizjSjrthMiJ1P7q27yx5e9N4rDjmwt
iHt8tC8PCCfA7HbzSDRJ8IFRevVzsKPu8rRuGd+PgIy7+1gyxyzwCtUE8Xnp
fuc3wAUVkJXEt60KExrV0fhlr+tBc6Wn9VAAcVgUSLVjjmMjt14mHwz3UvOG
kBNk2c4N/GPJWIRX2Tttp0wsnwA8pBH4JsHtMdZQ/JKhqlZGtb8Wuhb6T2zR
Y2OuKcXmguOP2HvvgWldYTYmHi7Ivf+azB66UzlmlzTI33ZPCfFPfEBx3tfj
hvcv3TG1VcJBMLKSDx3ZGcbT5liJMpYmPAauKwwA5Os+F1ysH90cXu8FlFjh
jUFNtcTK3srJpj9FK/uySYBsGBQ4CcdE6+1Um2SzcMug4beXchvCOyep1FKD
45BL09Uldhxi22W8kfUgE+arDHjDRoiDTJ+9m4f0+lYPpHj4EAUMh95Eq3oZ
QfNkj9lu3Vj9vA00VxeHf/pnWHaASOovGoqChjQZavwk1/8dyJc9RRaLvLTe
APWcGb5x+d+jg09knZcwWawcqw41YYA+k3iJfG++N3stI9qXA6D5og3+af2n
jI7OL8FiYNUR2DL+rziVBZzbzx2pzSpnhEDTSMmoUM2LWI97DMftp4LWLVQS
6+tBSBKu9mN3KimzxiF0zNj99MCYYtxEbUS2k+nybzsDK8AVfUcxm1gwz7Jp
fxw080mhhF5ZETZrBieSNA1v2qMe1h6oKd074dHWiP9pLo2bwHSxWozCU6Fj
HSutZ2SIvv4LRDsBFD29bNSaOwoidQfjwUYcTVjatNwGvZ2gjn3YLbgNB2my
wshjWs8UZeTkatf1SF/KGAEgn9+jD42HiX/H3kqnq6+yFbSwVjJNPEAzP01J
GL1L/Cyi3m2BglDBlUEjvm/2/dP8ArXw9lkNQP2BGTYrPKYEMlkGPrDybCKD
NfF8w9x+Pm/MFyqXnwN4M9Xy5FIB30LLaJtaya0ohn8fFk7uDcS7xCc4KzrC
oGG/0u4X8Ab21XWnc1ScnSfW/R8Z3KaIsVIEZK4GAxvDJj9/8b+6ogHrI9Go
GZcM6S+a+ZM1Pek58iOOLTSWwjsdjIziNIKydyN3VqTFqP5D4O4M7giDMHiU
45nqKb0w7N9IJ1bxGBK8yyRdAKnMl5AdzA+Gj7M1DpzCRh6v3gdB34BmWILq
Jl7Z3GsIBRRebmiNgBWEHEGbDav3LZx5eAwT3tDq4b+Os8WhWzYc9pZOGKT+
JoI5mZz0FebSLQrJqHd0Mid1xuiyAZxEbA8oh6D/UnjgaBL/qUxRgFSRNDVo
PMKk6oa2ACFqUfEmTx5HDO4OsJXn6JdWEMS1PP0j5pyG+HfR/yDwNiyFe1m1
ed9rMOf/KIVRD8Yf2HqE7N3lyhRZBfaTLZC+IqA4fgFVMRnghYtC5IUU/rL7
gJTz9ifyGlHJHbQh2nxpohrEKXqXD30RSHxfcB2n3CNdQYHs/jaaM5QAA23J
H6O2/Iup7WKJUmJJJLazaOWiaxHbLlAnqv7vigPQDbT0yYze/7HynSqcc3Gq
2DxkKOjX48d2PUGbWxnQqCm3Xw4O2s1HBM8XcNHD1E4K9nDl5K3G8+QWWZwk
7m8C4ZURdsJNFM86IVLdAt1VoEvIUW28KxLChLEmoDyMwMnqmQvb71Skz5Ga
XHeKxxrct4yoj8Q3K8giomELeY7f7U/Ihb/jtsjUCov01QqCu3mSdqI7S1SH
bYwhMsH99mAO/NV6LXiNwlaiSDyuzcOvE7NIcK9BLiR2lLTX0ksYu3QsCaEN
JQ4IqAnKzSQ/vpRtZ1IGK5dPWOcJ8lbCr3/epsm1x5cg8JEZKCJ5AGrenOsz
nW+LHdckhaqLbFYK6ta94ywo8gj1WqMpI1QebC1XxInx2SB2HvqY3FcO7NPS
1WPhareqxaC9aA6G1cekWYbsBANGZXQT7gqXUdzZCNhsOFfHh+goqDHW/cd7
LvEaq5icbshRZ/OWVG+F2m8TpgTYVaxYyuCvdt1AH2QDrH3pwz6iAkKkBQ5Y
DtoZHbSbu+L84b15tPfk898l0RPPNj8mKnCWAMjCuG2/1HljLBehrt2EoDWF
ttQob5Y68tcQnExznhzFDjSY0siz+LVnemx8tcfqBfVLbuskTDCsliRVDbr3
iWjeHIXk6QAr6SVqKwTAVxT8GtzsWU/5GvyMJwQlrzojh9E0pz9MOP1uDy7k
XGmbLcFcDJmOMOCtmcuDC5dEv/na47TEuae2aMoghmgnACXBIiaO2uTXMBG9
3RhltcaxGGsXCzJXiI7ldZPmGxZV+j/zN+EDK0kAZrslCxhV2pswzX47oDX6
Xjh64EbBIt+BCnhPEFZvf5A1nxv9IuzLaGEYdoBlmHUD/hhYcjh5yMk2w+fK
JAR6WytS7Yh3hh37H6313Ru+qQU2UepPKyZodE4n20N2wOKlZl2Kx61IAYtX
kKBDpvvp0vM6Pk6QjV5SpNXjTdNmtIirm4i3zwJsr335eOlRdlaVz+1YiMlc
bKtaO54xi18g2TsB6/CwzUwqZcTimR3SHvJW2vum+NzMiba6drsOUcKwX4dA
LvZzir04uMdOcsfep14ur9qVtE4zJ2StJMTcPFSIBpyCfcRgkqiqQ6soYQoC
taoOF6GaSVSA9N6jLmbGOopZyha1piBUXNWBGzywX99bnXs5/+vIlY2sieYc
6eVPShikZ7+b997f41X29K+l4qv5mBgqptWKQr6aiuUEeM3ULnFiGa/wu0R1
rK1ff3AQUnJLXI8WhpaCjOLNpztDOUztRv+HRXnpJbx1dRKXclyMG4Gurg+a
2OIf2qRrZBby4lq1nP8GbeEkAUPSj7sAutiB+wm9guPq4CgEYsSbhLt1Pw/6
Md4Qod5kWnYhZUZx36caJqkaz85PFqVsW3rNk6L04uio3M11rMAfRgJzMXKt
ZqbJP4i5HQPu0OIl0pnzKc8e39AJAjytK62yUMsbgBuNClWXtGP+4Qh9fRjZ
gwxMBgUOUVAoTtsinOXEQVrNXhadijIU7D4Rm61LfAR5afxqJ2k0xJDtzAl2
D+QwM6qGPhjEeyPwDmSUiK/+MCD3eUYFFsHkyf5wXLA0RVrO8a2yefvjBRSp
3ztIG8tyrpTDNIKjU3wsDogkovg4LVH4sBAepMrtBghxwkMhSqAfq30CoD0p
83jjYNEZUcnH89q1OOFaZOVvRYzkUQOHFZeUoJ5vecF9fI3YOdG3KRXiIwOF
HsjBjf5GQ0CTmsj+iMmHyoc1oSEOYp7aVXaoIbLS46DRuP+/ZNblJqxADKvO
Gy72QQb6cDqnlg3QJyp4GkFbLraOTEQ1/zJtUr/MnjVe1xrGlbnJqzIDMed8
n2q+MsA9l5E7ApIuWCnpCPVKdUj9KnvNuZTHz+66EjmfmK2+ljDtHGsHoy64
lm6yQY26SWaswEtz7LNVZluH+NnBJM0rLepSg1pvpsvxZDyXkWJieXE8Qa7J
OHROk8xtGAxFrCzqACdVAn8gitiJBJa56v/kbIrJqtt+lp5fYYjoE0ZjpZnO
bAnJxwSZpnsotCRMLMkxCcPDxDYCU0ZYa2ItpYUCEa2tn/n5MRK6+MGkNDDA
tTu9u1PYc22X7NB1S6TliugNa0wcIDerGJmBJ6FsewftS2ffifBIjoX5HEBt
Dv0znseur+FuaM+FgZIBWBAYVGRhkhGVFkavk89xC6vfenN0iEF9vHs7zXEt
zqSJW6X/bDo2JndLerTjzLB5Vtkp3ICJtHD6OIjLDXh/h3yUopTgUfsT0RRQ
7UMTVkpo4OgcB/Sp6piIG14Fq5JUavF5/FeB7N5x4Oqu5mKqmpr5d9uEor6k
cgV9QPItNKTxBhPCytyVhasrk3dASwh+ew91mxmH95kzv6dMMNRebwdv5wbD
aWGdT5jC5oj0Q7BBou3cBYmnO5fsw049pmeHo0JKDoAg31QKsh+bCwNCp3lf
8koP4YXE+nJLuvccKhNp+KPEDANsG3TsDcbUinnj1aODG9HauO3W7+Og5vYK
buVccMM+LwNErViUcOxUJ48NYG8ugv9NdNP8QwEiBgv6VFzN3BRcvJOXcokU
0WCmCVyZE3t8BOxDoyB3UzPtz2G/4BLOmuiETYrlgKTixALEZvGFFDYBrrjG
qvotwHOe95GX10+B73KwEMxeo6RoXkj72P8qyk7j5RVU79FqBbLltTOZRVkm
PezwFZfL8NqLy1j2l7YJS0FsHuKfyGUlBJUYyfWFwMNbwQzy91kQlj+aORFc
8X2evET+KkrQ3FVRb22X9X7e31TPaCEeaWSRHVWEsxE3W4VXFulpOQYWISOF
hy1Je/VY05916yChQpv84ColSA6BbfpRDINfoSXXzKPLpQK+tzk5DGM9mGu/
5JDTRSl7HXNzrOuA5xVQbk0eXGK3tc8Rkq6hD6JIK7NSoBfMCW7jtO+ZUNX7
eISWEmCca1pys7wVDAiZfBnbMDvtbCVY2tEeQedUk6r4+sVVVa2j55HdHbD6
Sw761jHDjHiYRO5/MBZK8xWqhkRwCmE9iY3Ahkkrg1VQegoH1ivzqXcPFGWc
3z4CYpyp5F2M1lziUlaNaBfajQdQc4XUqaTXQDPZ83feM0hZfojbEjXZN+zy
vnYcgOjZlexEujD16DRWel5xHkAwfdV7/dIX1SF7XjqqMjbUK1yKRcDEfpvy
Mj9TZOlGBUrEqIU7kj1spwfwn7TLh8w5SywriNhgcMSjcSAI15x2+295Jbxj
CFC+t6eogHvA6PQrDLFG63atXpmG7LrbNXLBK4ZLfO0DXa1svfL0wiIGbQ1j
981t3scaYy6gGE7cTpcOemJlJZwNhIdMb9WN7Mx2Rk08zA8r5+7Isx61fyRu
Oy5Y6n4JqWJbVNMn9LnUecJ8Fe72jhvCTROn01CV6fFOkz07tEau/WzIeNLj
gJ+8vwuPRD8w9vIib2mYB1gOwnKEhJ7oCDlLgz7XmRXw3Im/ILbVm6JsraCt
bqQZFvFHiQlrGuljIrByGseWQkSsgif44UtKxPAHqUXuvaQ5qoTVRdFta+85
IpIrGIidtbsZ8GOmgZOkP6QozPQqYt8fdN0IPGxTm+wrtw2lCoXudwiKRKHv
TSkM8HxdxIdRmglSnnTf2gfooWfGjgmxVRpogyyO3sdubKgxZwHymnxNxZYW
snx1051I1CkO+gLIGrrYE9vOJhTS4LI57K9g9fhiLYVdd6C5kDtz9rHeT0HU
tRYyuIZK97aaRsMxe0emB5rI8cGVBDYo3h/xBZ2bduKNHdGJFQQdPxAQ8EYZ
x5wCBpsJ4ZBeORxogr+GaiebZu4jMj47KQeTrMapWdnj10jt0vlK4Nt/OpYZ
Vy7E1UGD4yNOeRoLpAmiR66vAaZUdkIInuS+pSP0AtM/oDVaFU0GBIHcrXPA
cC3vC79XIVLSDSCiw0UK2g6syUNcjJznyNXVMEYtAFIdGvYrZjiOndvhSmdo
+aLpijpnma7lI9CAT39p5BI0Fv9xrTT0AiCZvNI/Hh4xMzU9YWqjEJMLPlUK
UhAcbMu9cVQH2ckIBJ5eKkbrpg6hvJURjOS09o4UbnpDoj+xXrFPmFrhf6pD
aCMQWBc6eOBAdTE65XBlg3v/NJ5LfDpLrcQwJu/bc8hYtqSJH5CkjQrRbADn
eQXlSpHqvlSupmwbpyTKUfoRTc3tzhN5PZHuUrRzRzJgbR72g/6Ez/t16mii
xyYYbRSGSZPzrtOAlj/Y8whm5/ipVqUT1GtazKw75lZUKjpmlUensMNtoPAb
cLP8nA9H3sDW1Se2IP0bdDGhJS93a9TntP9ABUy0XD0z8Hw0vk4FHu/JpLdp
mOe/ejaK31u2SN2cZnIJ06mdtKAyYLcEOfQyztU0vxv5keaQ3QxHDz8bm3XJ
sfZt+0zJo64KODXMc/nQMeatUi52o/n+SjPIo314ZBOqjphQgiiVuVGpjmfs
PZDFBUK3S3zCdcrMQmuQXnfdwn/7dWtMMk6juMNePeREigQXzJXaqS+5qt70
nbY/r4DmdJAg6XsVdsL54Stv2rSbG8GBrW4ITXAF1j5dJZIfcrkjHeA6rN7s
9Z6TASi3x83qBiRR0/94rchMJjXJHSCULLuLDU9CKxsB02FLKrcijXtNbmAn
IUVQJaC+0Os2eF6F8sxtxOcBhFNXx/ONToXryCquZsqg/e0R5N+BZ5ggp+M0
du1UriRirQ8eFuwW+7L12sqfaaL4dK3y+1n+4ejXBBSknmGlJ31MusSM9v1Y
PEvQ6khTWQ0/jvb/o4oo3NNKvPxth0PLN8N7GNtRF+8KGQA5WPROj/zyBily
sscFzm37vnqh7jCvF9lFvnTLPU89mKMWjfAJPZxqS1nLO+ad922VI4aUEW/1
I4mxqMc3GQFvs6Bmaufhv1gbBoj2XjBFV7U8ukpYVd8f8PQ5/XUTigwJ7HQ7
KOXbzcRSNB4tL4ureJzJqPty78z2qAyOKG5ier1ezH5zLKeWTpRN9e+Jk7We
ecbfbhvKSTaU2iZtYZ7SW/DpyF06iQGS+QfMlg5p2UR651eEtjZrqG13ppqN
kYG+WW2aJuNw81hsWpt79v7yBNKAYNlq+IHzGfhnndED/BUQrpPD4DElMzJf
r1dnVJEtE37d6VT8USa2DChjPgLtbrvrf521Jb3EDmIZX72Vav1rxxN4o2ZN
AM9VoGWWs5s+J1UVfvzPaU7RJEajK04qwgc1Q/cWHqzVCEhCk0+S/9AJwnyp
VlpueYcddC4gY+XOanFLARhqGQMYN+flHfacakulgImC0Nnl3QA6HzPtuI8+
WCNjSUxbryn/enCElKlYJ/q0G+m27zEIxnGwPxr0BlEIteNjBsgGRGj3rmBU
76Jpgq7CeLVXYDMgXven6L9bTIXF0pPiXGvALiesf0nKnXaR0jFSrzF3NSud
CAHmvO+lXBJuEMTc83b6zFf8G5Zt03NxwnMUV92w5820gDpxwfFggW04XuxE
ekWo7dc6FO2RHqa/fIo5Oab1LYYZUjkP/LRf7Q4XZuZRg6R2LGPK5zIYUuG/
SKoOld8NYaejHu3cJj1LL9VsU8QiXCkHW2WUkulrLUz5UgYcXsrnnhAjVLi+
dbG+t2WLnNSBbOI32F/VupQnm8hmOpr1+iueNmkoR1tiwhCbSIHj/ep5pf0f
d6GMARxxim6cuq4TY9k2AnvimtBZQ27v+ZtNPeWWzha2HUTrp3xhaDARVR1V
YyNxGLOfF0VDmZROVTURgU1qfKJPo9ZwR8F6A2h1BGfyOpj8eEXjCZmJTH1S
5RecyB3RveH52YjOy9PmiX5eehgCtQTnDnoElDSiVgWV2cYgu8hclhzunZ1X
0CTLqm6V5TR6rGqYeTvGl9zl8Km/dGGAvwT5n2yQkfXlP4MAlnP8mOchUOL+
gbPNL9SIRShOCqhNtQr0lBIcYOfPaNm4eS3+0acqA+J0O9KsLzBYMoMUSPm5
Y/oKpLx9mqnyfEwoz0yw/COhXvCoi6IY/YCVZ9dXTx77ym13dJbzjlg/SZVV
r6Ox4ApOrQCPfv6PtoP6pkgGFFBlNKWToF0/EjO2bcP9FBcWJUguPkF5Gcw5
6cIJgxvbTr0WHcbbpGu5uwGFURhnA4xiqSzSOqP483mvFmGii3VbbFlqVmfG
xW0R2GKQuyDzAb77MUIFY6Fw4EPAaSFXYhTWZTB5kQuWHSaJRMxHRecZpI6L
TpWtDtwxrcUGnfrYHAkx9VVmmhysjt1MNhiIGnzPJR5m1NU1kna+L0SSXdcv
DHsQAALoQpvo4qBoEJQZs8znyDLllGTMyxwL1+Fas80f0bQIEQTtSBp4qlbi
Bwh5Scx3C1Y1eFCy7JJqFO3ykxyssrTBsiRwgepF1rWkCAChDnZgdpDB99Bp
dYjWqJmzvyHxUqlD95UBXBvApIHm5gwv8zMKCf16aWT/dexo8CGDyFv3KEts
32khu7mxQT+DNK13GWvVA5f+U97L8pV+Mo26kGDfYOygEUIu+vPBD5AqNSD2
ThJSh8oVEzUFAMQvtGig4NEL4xaRcdEzRDKcmi4vLFeZmdWmbFf0gmmhbs1N
eCYzx2aiKQ79yzPPSrfGKiWEE4f6CmfNQ+M/6HRq4PrImFR2/ER/HIBAB6po
k/USSp0M8qvEueEEgSG/iCyTNLbIalx8JhraU/GCPzEzkjB787kHrGzAON+/
+wRSofOi0w3e7x/DKihrMCplGhkJudGUtdtwQ+S26MBJkErzYpwfC8Ds5IH1
zy0IkySFySF4/vWQkT6ak87Jt3gI0ycqaij4KIycBWU0pG83dXjMcYFqjnNm
7/crXp4dd2DV2Q/ZpGqSu9y3k0gECGZoCHso5cNEQHdn1ZDRKpgz+k5VBVda
UkELLh6Eu2KZVqgWGgzdMoRjHapf6RbrAv/Ai2goHsQM1m441wJkDvhrkMmh
0CkeHBri7BWqSTGrk6OuiIj6Z7HlTP5te4ysgXJ4C41vLEs4CwB8epXJ7mtw
7gJ/wBhrYV5liKXsSFMpF+p9g2CB4aHeWz3PE2OnYrm/1owN8m0dNPSMvBXB
56CH0DNDWkqnSx4NofyzTAMEb0MTgKVnDH1IDIpwmYX8Tur6XAj4MeevxNw5
Z84wRmxI9tIkL2JuFycn19SGc7DTvXxFXQqbfurIdpiucubL2vylq4BGdI02
K1yBVzg+ua8KN6WL+XESikezUF+rLNtSmW+TGBO2jPOn4He9aFvgKAcKgD6J
3dVy73UA5XeyoYmOdde/4q57RmIiHXgpEBKDh/KUZm/EiyR+n0Do1tolLeEX
7ptvIHPVbCXXcV8yF/7rTzWLWzNpKa+8kc2uvw0DS92Ex3ZPQjmtRlhaOR0B
o3DL4hSkyI0O2Y76Lq3gbmAHCgkXIU1lb60vlj9Lf8zcIBZAl0kt4Upvvud5
TT1dCQ9wPVzrPIKeEfMUtPy7cT5zRykJwIlUBPPnc9ASVYrbhIdPBRcCnKTS
DMlCBC3NkBVPGodHtn1Lx/JpsyGqC2WPAgKSsN9+EZ9RJXtR3Fwq/ePeDQAS
6r4b7bB0unWAHuPYxVXtKM+uLNazwMmjlpAOApZ9UbDANdHXzOVzrrLudsa9
62LPDnzKS1wRLWt2W0xnP1lHDufIv3CZ9OWpTTgwGp8W6VgjVQXPc791r396
dUn+GQH3tbmCtozBkPYvmuOwUKXJVTrr4H/qhbElT/1Po1fcFHOY8ncdByua
yhNT9yHdVlTzoZFzpCBWEJxTI+AhGpib+lK3c4X8VYAzO99XA6ERXtMXxkkK
mfmrcqJPa8OHV7MhRYbZGTXkelpO5EJ8o8sOKf88A1EwcgXmRIfnkzkCpsII
Jr1LcKKffRtPAWi/lLor3q83ENlj+OOJQKK9S/PJqUUeW7L0i78ey2lS6uNc
/2c9DCQ0xMsySPPLn6ZExG3IipEN95yNYBBMaFlgCwLQudv8IuI9/aXWNH50
VLRYkJUg61clNFT3CCO77eXbst2HFCUP/jPvrROGkRf7HCOyqMlfUje43qHw
kFRcyr9Zp9MERClt1kxqTpxm/d7LrCZtxY7s1EOWW7S/bXA96/5uZmkSOP5H
gDrJLlcpDsyO47YeikYR+QZeo2dFPJ2buqKBsLnJ2ShXzo85ZziTVAMRRv/Z
Bp6b4xXfZaMAMyd9+D7CamUK1KxJxBlDUWlOuFyE3FCoeULjMeFkJEcNKtK1
a4CuGH+JYfuLWVrTRoalY9tP8GAuc4YmHC5OPa3B3d6fJZGuBZfEZ0c9BAB5
cv43YoXgUmuoS6mon8vDARpYlnluwqfsbNt8yCY7zkdG+gBVUuMy7NnxeuOY
f38dJOft8+DBO30S+GFh5PwkqZ9VnpwlPnBqDLfRVoR2TRx/Uax5yjaRIZQi
j+gy0zLcfF5j40g7zaoWzRLMi014+zFLBnccuBp1RirWu97oCiREJbXd3yv9
jljpT8zmqBjEsrRPFv9BywDLpoArk0cRsOC/8pzaUvvzzbnqW4OZ06zE7Wpu
BwCTUc4x7DcHPyUIpzrsf2o9X4wimF1KqZbIJDgY7KzZyKkGWyAvwK9arv8w
MH9P1c51D79xsgMHWYCySTdW8TyyxEbiWaJT5iAzY6rTFAlavM6v5yV/1iXz
44jMKRpL8ewSL4bUF93aZvDMo7crScCVWpHvReCL+f8RVCAXYw/3qDeqIOnz
cyZ63Gd8/NGZYNF4XwuKZzT9z0/JeblsnnPZzG07UbB0NbbB/rV4VpHogwrd
RTRiAb0bzSBxLff3dy3FEe920o4jMi5FLYUJ11ap2IiXzc16U3XJclyOxvoc
ONW/z2R3cWCIJBvSosKVfpDpfj3QAM0CqexYp9na05iG9666KopNPxExqLcN
mOvbEFSomylQsRrvlEaRGuNcxokFZWOk9iTt+a6SgI8mY9v6RB58daRc2Z0g
BA7uNF7WdE5XKloegzYyTjblvlY4g+J9VsA3MuSWDrRU3a5IqqHKL3QpYBmv
AJ0PcGz1k1zIO2gzFyTMzUKDcRN4oWA5U/R01dfdCeflnkG5bklLD+HjW+35
5lMYgFEiWqbGVbPpV2oO/L15xj3+mrtuhdE+/7kR6+t5fFVHBHfPF0NhPMyS
Qbkt1B3myIlaWNqS7fqd3idKL9IuNmafWuN+4vDDHtFTQKrWb1x2rzYVlg8a
rdz0lkgEHUXjL1e1f/2DiHS6dUZ7TJXO1VKFp3bOeZHTUg/tKcbfeGgF6cz4
roRxDEUsMnDtl84gek0T6m5z9RIfje+lS+wdnGCJWsv1Oh1EWR9RafV3ZuAk
YqGmeqDUPDZzV4i48It/cmTnh/owTVsn+qozbMj/4R3obCZbCTKVWklqcrGT
yeX4Kx7FxorNXoYwCT+XWggoR2RIWjphVw/VHguK+HBP+aEwsMemgKoUJJ4Z
QAWpmGMDv8lr4wjvLae+rOdYicEU6/Jvl8JUfdntFXI2hm40b6jFp4GMKYkN
0qOchFFkP/yxvoFgxwzs6f1ZkI7rhsP/Zs67Xbt8alD0ovZdjseGY8409tAF
QMfToqk4mYJMCLMXvJM2nWeAtgA3Jbc9U1KLTLzbdJJRdkd/AJB2RkIVFD50
cxr9Y7zewc5dBjz+p8x06A9PbJlX2c1dr50cTYM6YHGuN7mIOYAbyqYgBSAP
D54oMvDrVkPNy7EulBqtb5SKlTDKFxxAUcQc61d40XxZTUhScEUurauomiZf
t0EvqMGj5qDD+EBcrALotKvM/nPS4MmZCp5enkzesKTp+EDp/ZiUdUbxu/Mv
ahqm0JIN0/zMZVzgpCsuZm4ZLrBXSDVAMtcKVRRQHIsG0MJrxg7dq5JVNNKA
0eJWDGoG6SflY2vzA8xuqvFSA3+kp41kHSEnoQFvm6I0iaJWLPLoUJF9zagD
teUeNYDVDPo/0g4UGN3z1wKdAqtOISWGN7qXLRdJLIzSHViX2Gpmd87WlUFB
+uUeFwcuEqM2i0BBneWjR14SWYyJZSWXDZ1RFv8Rgrde5I0y/KFk1M7nLGKl
RGF2wqWV2xJ/+O6ohmArVnQrMrQBgtVnMrZtSaSMwNHSQwKdtZClhxAz+Rw2
3uDEs4/MOMIO18KX6oNSeggwdjzzLmssyiyk3xweyCR/F7iOxUmrWUyqjP2o
9xtPPnO6eFPoKzHbDZ7m2U5jgVW5PpkK+4ek3ysotQSNlbu4YTHGv2+BNNca
YDbdBYtIJogj6EFPgoe9v5v7ApTG1r8aS7aVKzagTsl3FKkHhw1RGNj4HRTs
E2zrGJ/r6VQWzo/DPUj5wcQgYqak9G2hn0Qhd+qFPPtI0bwbNQsP3Jf/EuwF
HxTWTwigOunVq0f4nN56bxAf6vALImywSLODkNto5kOWRK8GiZhU7oPsOtfx
V4P6HIkVyfsU2vT/kZWxQ8utyVDbu+gfrjW/wPrNrRt6DoCd5kuDpyadKfgP
iAWYX/Gz/95Np5l45+qlJkK9MwpSEbFPLRCgh/sZ+y+6Mw3uG4WEeYFpMu0o
TYe4T3RAuLbsHqZzAvSGqdKgEICVCFpB8PYAWuGSlracQs7fCKIdOZ4HXDAW
Pw9b7kIFEwIeaU5pmYZZsFdElvpMxR/KtFbXTgx2aOOzDYgbferCQNVZBszF
xAFabuwe0EmVU8k5yRHs7SBzq6OwNLisZ6EMy/cMaEYVcZ7zFF20ZnVZOLmG
syNNKYXTSUxOBBgHk0kli6M/8H0M/lYwGlA58lMQIczyN5gzoKzAXSYHkZuN
sy3p2hQQEYUOs0V2h00fvoP0ceThb9CiNnji6BbY2y11VFxNkPbk9BA4Bqc8
wzCgc08Bgrggye667oWI2WfR/28tSKPhYraMw5P7Mx4Er1zLJFiYjOwhCMPK
qTc3lP14HgtiJsIv9gS5qhlBnll5WSAUo3rEz4Z6gLpJr4m0gngawVOkxXuG
N9E7gXCPwG36OqeWE9m90A67SeUCE6n2W5QBnmMZEtag9v/Y6hJYuBBf1n/j
eee2TWT8kpn1FHHeNZ5UrAzzPv8qge0NdrRHlk3sape3U5QxQXgppOXYcoxH
YqGuFqy1UyKm4w3lJuS/icF7TjYP+ezmecLtOStYMczHpaXcAYc2/Z58x+PK
70Eid+qwQ4jSVOrIYhdFCj5dUbPhu7pcirxfMM7eiU9EPCjrcfnfMgfqQ/A4
BvKWqprD+gG56SfHZ3wG0SkErURKYcrnWh05s547yeXSqA4IHQvO6dvaNXbV
VD2i/BQsfuW2wkvR9oTgxil2+U1CZDLUz+lTtbmg4Po7+TaJDeCpCa+ptLDn
fC1Mh3fdjL5gzRgktNuXIvEB4a9CEHHwSSiCrvNE1dVcvqHlYuGqSErDYD1Y
yBPoC2NldkBHUlQ00Ve7dIjGQj7C4U9UJijrz+/62nQ5WWUaXtrKsuIMJeKY
5F1dYXkoD1roMKTy5GX5HWxqYF5IhI4vdPLMRgvpNvk/QOug5zykxqdrWU5/
8udJRxYTcRTBKp+Bl2ZcVZNMPDy/Bzydf17RT57yFg91o7XLn7zjALb/ipRD
VfB39/FNHKmEb8smdr8M+1Az2Qxql9QI3kdx4Kw6MRr8Rt15N/flt8vMlVFW
HPp8vHdxVbM5XSqVxmzWpAXAW2N1BucNwdFKONTsJKRQzmeYo7Y+7c4kQDK5
TCNd1r5IgT305yRd4kQfPD9+9mnJdgXELXPQYnzpY9WifEhVHjocsvgrQZV5
tuxplN79wyM+FeX8Pd5EmhFGAZlP2LUVJWU0pUPpf0scBFClclaInYMPEoDO
oC24QFFnW0CqE0uUxK3+nunXa+sWAc/m1AnAPHGtL7H8jnmVr/DmG14sU6h8
3iUrVOjuGfe8mdATHP8z1sdqVtxuQf4Aay8Zhmbl7OskP9NWTJ15dVLdRSpf
2Q6RbjDoJck7Kcix/yWqM++fPA5AVeZlRXmDNrpFOx5VD0f5401GfBAN6J4s
hD4dRP4EDXzA15XNO4wNA54GUKO1E9dC8OaKd7vq2HyhkUhkOB59QRlNZ5CM
sJCEzZ+ClO094gCXukNcUpKy0G3lbad8s6RSrDysl/Uife1vrYhmZ38DptpY
DhtTqeilhHqlpsv3mxIAMWD+fOQm7KTBLu7Fkgk41WnEgsVwKcrdIfvTQ9gU
/I1/74ECvo5a6B2Wx2vD31vD9r7NGj6gttDgjTB6f1m7gt09uayATMWjMoEp
uamz2l0TuMqOMr9huv7yHuLjqntQKHTu2ezJMRmBgjuH6b35gt8D26Nz8cWa
qjXINg/XUfunf6F6XmYVSGvZQuSPwB3MJdCUzhpWl7jmpe+OYAlwKZzhJ53L
uuwl23qHXg7f3BWLwQFcB3TBhV5gTHZf18RZ+juHD7IwUX0sY6Nxtbc35EO2
u0Gbuk8vlaz1Y6swkmNMdItk360CUKNM7yMbQui3erLu1LyFDWeCaQADwK4b
hUWtXV9h8bHDr9LtFUQCh5YQ/HnUah5xWMb+ie644BzDSvzQqZA+a0zvd2gg
lT2X9FGOaZk0WfpJXClLkqS7e6/opVhw09dOBMsdZibU3OaOWuAOaq0skAjn
H/45E1KlIruY/uib1ReYOElN7f6AjkpwQxjPrJMN7ERd8ubszJGkNnbCsxS5
qXpqbvQc6CduVGUrNo8wFwvY7/KtyEahUObpx0CLGcsMZbYo7S5OkoscSHTI
C5IPHMUVveBSVIwbwng4khewzXeYnz0+v5r1c2cI8yBcwl5ydhYltjuVIgdB
1blIvRIc4J68eUy7OJj6rCjpvG4G3seHWKcjh4RNlRzYbv3b/62S0rTWPt1C
vpf8T4gWnS9/Us+Ih9JuhpGUWerNvcNmtZCd0ianQEXniizyUFuEDVfoeiTs
v+fjb7wwDFXjYO195+b9a96y9vmIzj+0+VzzVdJz45h6dqqaknuQRBG4g2CE
XIBISUaLg4rcZTCOKkOA223ZpThxI4Rduucy3UQ+1GjEsdaBLgVPUwLzJnHX
tzOnRQlRPoV+zEipjet5Yhwj9O6P39RVsq+x23FwMOCxhyBcSStKYY1+0y3p
ZXXBcip3hjZr+ANByv3SXfHCXaoqAXbW/w206unolQsTJciBP8Tbmb5IkBxY
LJEZWh0ka/kyuPvYobuqWHvmPtGPsPth3lxiPS70nw+HbPOzWSgxynYH8ryv
lfU70aVTWu+ndYSn/I7GLzYDvOfZccYasfLWAoiiO3jHufZabeJKrWiImRV/
5ugCDwhK5FyaTqPwPvXLxAVv+E91dPeeYRJbY8H7Jv2Hq5uMOR5O+excyW5G
yUsVi1g5m9Y4DknLjRHTT0j/Qm29qAT5HuI1+ClpNaCspqO/mtulM0IXg6WA
4y+PjQjjM6PIb1qj43TWiK9oZRU7FYUMFVWduXcv72X67TfDSV436eWwl17q
YjQH0p5DxoWlFnEH/VFPvWT61snsc8bVONQP7ln1UoD8FFhmQ0UP8x3CtJeq
c6UXffCnDt5ps9+JUEcBq82tpvyk9s95J/CWxFPi4hijN7x8Ox+Uflgl3Pwa
p1UfTpPlLDj3wb1ZL+xKoQAo9l1YXt3YscFmLDlTG1smL26V0O1Q1Ld/vLQR
B/xu3yPEZOpPFkA75Kxtws250bkrb3qmmp0wwTdHnjwLtXH8LqAo4GOT3iRv
SacGLEcQF2RkMHOUiPsI+neNO7Fub/JtrVb3d2pzwlKOnRqkosFTzCbTfqjC
zSV5vC8R9TSVkvoE7dMHfyCnCT8GOAP4/3TphMoYV/XLVjhn//gSw/C6v/53
G79GU4BcolEP1MsY6ZDxXI9hs55Un/UtW+h8E8SMbHAAyfGw8dAV22vZRE1A
F12Exa/fMVFOinIEfWC+9VnHaZmThWBIqwe/dOs4CDPujYvtKzflemFRoqgO
Y/6RUCxO3GbcwIXvV4tNOq/lBeeZk2QUfjxC6nKQU0Ws1k4boFGEuIHE3klG
F1jfnlPNyvVE21y9sRpdn9EadUM0HGxMyr2sXqAgGRrG4IsI0e+VYLvcmESd
CVsojGl4g3Gt68Sqyi+xnYnCBhjK2gVJoYjrF8ZPZYV7id9k2zLSwI0uwRv9
TDqcBit2E+rxYEagmelAu+/RGAHH4I6YCS5p0SHbbVTV4RNuOOMxKidbzgvI
yDdxjJJhF48ICW8N2akd4un3CRXajI/1FjKoo+rZMA4JaIUD/d7rojEX9dr3
FGUd3TqPecjXKu43v7W94i8dAwEGO9Qp/Bs6a3GqLHxekWJtBHd+0tQkswqI
8Lm17FoMd/BySANj22WYribhHivGTbNqj65Eb4w5Eyy/t6El3QaI/LkeEvy/
WRQCU+JA7XG1vC4SRE9KtC/vgFHyQLNnM3pkllhwPJfc1sIQKpsXsWGRNEe3
1kX3IKbGm4HffDv0dGDwsdOjdMxZMxHdR4r45QfiEvb/9T0/oRDy3zfqQVIC
hu51uPg3ZzgAy1e03/vRjQDpDwGRrwsiuyHZ7xM7JQj13Qj0B/Pevjz7+iPj
3shqgI50SyrbFyZ0i8mv07MdhVxKBA8EAar1rPdOV34FfDQDA0IczRGh6sWd
HHsL6CEbKs7wkTs8XAjfrotlHXPDJHcgDWy32tkH3eecuhC+Dhii8Xz9xZlR
FT9hTxixQqKUG2OV5wXxb+Re0t/TyB54RCDtnfDFq2YAAzog8MmZ27t8W66L
5Ru1G2vQ4CC4pkIHA+2YHHuuGXdm/pgUmu9JpXFSC5LvNk3Tl90Y0ZvRbDiQ
sDPOWRSRch6pHOmExy2vYG6lQCt6tHdCtNEdgxnlHIImfa1DEULagku0mGqD
I5xcIN/WB6VDImMWZxmWxpzANuoIJTV1K27SST9sWDNMF+3SzYY8QGA1Nid8
R7vcGlMPFbyRVQOFwSQ+aucm/Bgql0eV0DSHRCPZmTBwZdhSmbCTZsSN9W8X
8ylU9L/0qcbqlje78oVncNQ032RCMwBEsb0HhNrsH5TWlI/bCCYoKNs7iin1
8YzU+y2BRYpI0Meiyr4ALUmFam6Sst1y51NgC9sHn2/5osiXCyFkzCWQVxyq
Y7M0RYc/OQ8oy7aVol2NEbHxFJ6efKNM2XNySS7NG4kYImusOhLA0CEnPRFY
mKjKcplw7HgLMFHM00axC4JNBv3UPSeYjUcL5vQn/eq1jdZEZKKp3aNdBqkE
7B1ZP9/x0xzb0RDj2q4cwKCZRLrSQCn9OzSuSQQX+HvIlCuzqxOf8+gDsysw
sDXb+Y54lK+aG6CCQa2grHDdvIClLiaA+N71itgotlaRKBitPsx6Aae2ojuy
0Z4WyqxgGGI/stqFqoq1hnTHDB0orjNiNMosD+BysqivjaTF850tK/EoJTa0
8g458pRL7oS8bD7HNsgRdKO34mkJHGvP1I+BhyCkuD5IQwVG7bM7M+f7gd3K
P7a8qdB8WrxhiUmh0szk6hXh+5OCyvP/dpCqXyCOs72Qa3dN4OeAr01p9Rbe
dVsNikWTia9ovUL9WGDNlZ+veGIjFqwrLr6VZBVTAvNgxcRh7c3AptY8PNlQ
zqgFEoBCh28fRW2X/8jrMXYoK3UTc4yNKNUDBq5RkZTlJsTjSDosm7Skr1rt
3Cm1ASRc27Clcr2fpyBdVAElUfa+j/nKk5GgqB5AQkZJVLhOFI9/ziXyoIpR
H7ydkre8U6OdMm841yX5bzK5VtxQj3R/ygdq00VYYgQZm/Guj3SHlupBf9VE
//Q1SzSkC+eKXXD1nmF/xhLjjcLS7nq5t/hk0uSjNTLVlqgUtQJpbpVsN9cC
u6RqozYWfN6fWgvUxCmO/IrD3Y3DrMqdciWkOHaYSJbf1RciHL1vaAeZE3Qd
rmIFPMr2oP48iehbZ/nNfg5r1B/k468pVQEq+Hv+Ed1N0Xvq3uXMRmfgOCmQ
SVJ54bMBvxzPW19EAiX+RQzEOaw+ffsNWqj9RmjMVxKw1dyIUs5/IwFQM0vr
ZehQDuKP9bHpvHJXf1bqQfqmO/N2clU0zTq8D17C3tSy7+CxVoHSYCQzqtDE
paGROZEpvW9Nz0oiINC+KhT+tQKw4ofeIC6m3E5TUHFaEX+seP04yBQxEjos
4hF7kNTmQ6Ml6ns9wqq29pUr/pTF40s/zBHXD9VYUWQ9AvOtBsMawSLRu9el
EZCOvsidJp5xp/DzENjl7WRJlF33w4XPGRuFSc+T1cE52/H+zksV6cEwf1Mp
NwD2OvpmXtrp6A+d3OAXVjP9D4+HRe22qa9OeJ0gMXas5xhqxWK1gunFh0cc
HUHIL4pGG9iX+W64+FBdJHZiOhV2U2rj+Kt3mFY8o6Sa0S31N91hHXFpJhRi
+cB9yEpgzD8bLcmOVq6cXieAeTgF4mdHWLGNdT/Tz9DfmS+WncaaY+0WYmyH
FVr6cJ3OElSXQw2NYfO9AsVSArUYiJQafKCQ/B5Dq2dR+Uo0pqjjoLY5KlTe
ZbJzMANlW6hnxiEZt2IMAhAoSlPcWdbBPK8Pr+RS0h5X2DocW7TTcAhWh+2B
OZ1vLWK1jE6sVVKVav7JG1caMHPnC3clayRXM09LGKi3MpA5QTTzojDDaBui
NIhsuz5GWG12Y8j7J7pwgXb+QBZ5bVICIGUG03qqBDJL+bJ714pb97RQxSKN
V05s4Hlt7UB98OPaaLYiiHk/iXq9Pw4gr1vkVNjhhWbKR1B89sQNbZUVvKgI
r+HZYGQx75K6H1UMOVQDF6aYIwtGVFyLRDYuQhTdqhNobYtjKo2tl3NngWsH
S4w6Bv+JL/jAVhEfb0LkrZl1JFk2fkfSgz80WexQjDVdYDEVP/P2NakrJfNn
QS49IMHbAXSQLM0d7kc5IuLK3SXgoenJezOQFurG8he4iIRDxYpmfy3NyRke
uQFVhnSLGDzsqqEvp6Ts6cOioLzxbVdE2l75VnHe0CRSl2jwxdsmhSZefUn7
/afKVUg6drQ7T+jctsv1cZMi4rz1hteSUBR45LutDFRRe3Hy4HiFPcg+PBaB
zsYuAxKwr83eKHqa5GlzyUr+zNwzdX8xiqvv+r6x1x5IJ5wplTjAUxR0RK5o
Abu0jxZhXsTmi42bgcQwuh0OJoZCzRyCQ36mFgjhfh2htaJqEkK8Yd2KVuwS
BKno/xQq1IMOu0L4GKVd95K0AC4Zuw2CtNgBlKd9yHdTFpdpoITncjq2l4an
qcWmdIXYhOR0nOQ9v9QP9QQEb0yWiyZ2636qqkM0teWJVpC3IdSWijtVm3YS
nvRSsJ9ggrXtiy7MTEaueqLWL4PvghVlZPtCsa69M36Hu2ypWL7I0mWZcDap
L4GxzZEHNTP7tZDYHJcbMO6qtQutUdSKTqiE4cA7Zrpiul8Cl62LPHyJ0nT0
BDo/kBSa4BX8mlwcrYpmedq1iGpqpqnpEKckbCugaH5UkmJfUo5a2PNHGaby
4My/S2PF4my4DgvWikRvX6d8prQI3pFiuOCpQAJaD5Wz4myecUhivVNVX99E
8EkRuDLatN5BMz3LBld3IE+vJTu5kEU+1qe7D9i8LpWIhgdkqSqPKRPXQqb6
+7u9z9sDa+IWZbmGk2bcZLai9rwxq+6ulgS3C/uiquXjRSZUw+46OoOOm0Ui
S/Hp6h9FyzFyVWhtJoIDA13VzeqykBvoibzQMDlk5ExF297+fjgDFYsp9tVU
9dBzhKVikFq7FRxhbpJMkgL+B3rRfqamZ/dEk25wSYiRQCr2ZH4X5ncqXY5U
ljrMw48XJTNkO0gSKbO9nFagc/dftqQpbQ+qwd/cakSxEnIk2BzFzvw3UrNs
HspeHZYzEBhFLSdgjgOXJ5Yhwp55TdY3kLcUfNWs63kRi28S+gYZTybgGKSi
UMpU0btkjO3xNkltKDvSgE4IUqCcu4rXQHiSA1nItKQdzqIiJjhjNfu3m9Wm
jvuhdKkkJN4R/1edi5gFW9/yIxtxUSKbM4pGb7r7TV8N0w9LJBvcDteTyEbQ
fwR0MN7XLX2JkMOMh0jOFgzqgsbb2+huPAZA0xRj/R8Wp2Ol7vpFVx1YgnEQ
syA5NzWKnzvhdY/fmwH9Yx2WKSCON02ZwbNkQTgoywT4y8D2IBCLvjMA3y/c
/GRwI1w8pengvAxs69PCgRAYKq0qkgP2ofyLaWpbVzfw0wXMm2GIGe2iv0Wm
mU4rIZQeV8GM039V7kcGRKtbSgoFg0p9TKSanx2nK31uBSqHkMLpURehAwl3
tXN4LbAqMONI5m0R52xOWWyqGEoj+Ha81CqKjBiRypZXLxkYGSjaZJ40o/3h
LVnxA5qCc4SaYZO4/EsHWubUZOui7b9VixSr1tWy/XfSWPthdebDPDec8jME
H4NQcJpfbA53/R+2U1QZyU3rVWCh/zB8dvqUGZ8W8kGehdrZ7y0/DScxFQL3
v4mN1QW4lGTfmgF0RAnZLRYiGATtUNKuSZX4Mg3NZmkn9YI0A0HU0tMHnKQU
XBKcWP6nkahpu1NaMwp/MQmzmXjKyRzyWXkVkqYCaCCFsUYtd398Z0ma5jTJ
+GkQe94cZi11QLVPEW5hTNWE6bwZNgrpT3/GHGxgdmrE4cKU+jrSBqWA+OnY
MdMYqggLkHyTTfzUhKU6sSXT45TgUft+mfXHbkex9/s8+h+jAv6qnz1uR5Ko
eyYz5U8yvxTk794AAjFnI7bHQjxzbmqdP+ZOkvc1sZrpz5pQYoVk4PpeyIiH
EUA+HYtYzJBUuasDzhwLI9UVx6sRBABVSED5ZsG+IXj1FTuKteLSjV7+Z36C
A1AO3a5KKtGbEdR5OXPL+3Flw143LDOqV3Dw3jWQDaPGCintOPev9zADKsxP
TXOZFCOld2q30sMs4jl5ZsVn9pzNavweEZGScNYFQj18BRl3rywDefZPS8rP
tkGgEmw8Bw/eKO06qVPEewE6Qq1LP9Ry+RTY2mQZstHEuEJb5f71f7NCkPLU
lDDRfihAarkj9scO/H9bK45Y+XDQUCGRINmf4GuuSVGDHZHlkLznpzbnAn5e
iQOdHLQtvWkyu9OTFWyp///s555ZErlqlmlnApKLQFafH9EIv9IdFPJLlIjK
Wxx5bIi2wDAhK0BZj+ysc1+hbRjF3bjuXnf/s4nIO17T7bNrSCkFR0UqLNTA
cABq652YCDrvRokVf6tGHLhd4F6Xgcr5iUYz9cXUfExjBt/AGP/Grb7VC25P
FaMS4M/EoZQVDdEtjEjGvR0HDB5fRGDReAHFCWHOQsvOEe4bK8E5ApI07sro
tdtNvEeXN67vKJIYG/CN8Ayu//d9dnaSp7IMp+Ph/KKmcRNeuseqsUHlLFMo
Cik0a3OZkKOVbMAF0n057kDLAxYFwG1djYeVE18Md0PZulRjSNOcU+1P6ROI
WEFTrof2XAx9zJwek5zhm1B5FZczeh8oeXVhJFMquTgA2MOXOMckRtpWZvRp
f/qGLX52E069BVmFbmpCNwpsv+2moMokH3OFq2MPH6l/PhKDnPLta1ERfkeA
Fpq1MYf1J8YJVvappGt7otWBXoKvp8rT8u82gLdUPw7EJL68k6OwVjINVXsD
pQBH6nOfwQKCcqYNs1hhRgY62PbuJV+btOHOyC2lv7Y6xUsQY037ZePfIoH5
3N1xIh2+CiFOP7rLjoxzGysropnODZcaaQzfOO2kscLLdinbRoGjen2FU9Vg
qZs4ymhjVtPNKf9cBHw7t8TVQNbF41VrV+8UlKuGn0okqYO1UAnsjXZyau4P
v4PLAmaTfqnTn983ShUrugSGLvNe2qPTN8pGQp/frDN5KC47ar4N1cgtWxsr
5ZSt1Li6PEELgzrBK6Q04VGc1U88GelfFQUo4wVF4GXyFiFv4hyyiuJ/8Lq+
BDjTdsP9TzYgc+7I7FLmUI/HBmzu16sFTP8McZXydjlDsBuIyy+K5LXLfkXk
V+4FuVK8ZkNzqbXzSgI2+lUKubf5zcp9AdoknVxJ+S6CgGx5rCYQ9qyXoXIC
VQ0nTrdZeDWvkWDOuWK5B3TTDLjYKTJwyzT9/8g6fwFCUqmIM0Z1uGX/bSz+
AQvAIwK7mC3UMs3AtnWTzYOKpmW7nl93c/yCz2nqp8lx3U/U8nkff+7yoFct
ByOeh7uMoWWHCpCHzoj4X/QSR3QuTgRvHowZY+z+9lCldRQhFk923Go340fH
unjA3lxM1590sDaCvsJ4oe1HhSn4k4r7pdj/ClxFrmJN7Axg7q09PV/yr5X4
KhmoXeat7+JbqvotFweqq//QUO8pG6mMGQ+uNoqFaS8lAFPdX6zH7ZgNzojB
SLx9q64j7AfA3KC/qNjuzBMO04Yk3O9YUb508EXtDVBzOGFwuwoxIHtxhYMB
cxBFKx7JeZItHSJ3z8MpgGQg8XSgUoIag2D8XyRBfGJ4ZaDmOVcIsKgHFv3s
AkJzXEfZKhyu1Shnw3QVAMcqWmbLuHajaIV61sY0Bye7oGvCbg4h/p3USJLC
NlUGgBTlvvpSeR4KnbpXYreEDRyDsUH0GdeYOdGEV9ITNdaw5ZrTfsFLZjZ2
Dts7AeuscpQao2/EwKkHBVSdfuk91g1mBbJvq3EgbQXqY2qiCd9X/VHiyyhl
O476prJiR1AmJATuK3Z6uMzjIEPORoOjIaZUXjPzNYLiZm2krXxVeNE1r624
3n0QJ79hmr+NOE+ebl1EwYUYD0nj+QpZnd4cylEU3oIaH3EOwvqdufIs6Ni+
Pe5DD73wenNd7aRHDZuL8wmfDJEOK1scCvOrxHCOyqfwF7i9nc9rBw9Stopj
IJbATVBdO0DjEk2x8JvaO+LfDgMxCrO0XtkhyNE+JzFYgyolzcNtenhkwXUn
PI3PfvWEWpukwT6/Vg9XaLos/P7b8MD9OwpcRsPYZB3eIs6GRCAovlDwW/ng
bkZVRpjIH6JLZQukSpD+Grf6qIgw7zXbhK/+nkeHbjK9GchXWz3OcZCAUNu/
9to5rn2iNpMhVv1qlU51QqX7yZkYkgrwAHppQU91XQg1CwL6Lb1mm9G3rMbv
6a6tFKpyjGuBHQzCl3v/zs5o9hoAIOBq6koSsAXTh8u9sv+XOB2GR/RQzBQO
jDBuEiB6h8aOyFRayxWmfWfK7htb9J6U8TSx04DMrDGeIK+dgcZLaX3Qn1an
yEFWDMknuqgLDfo5sH2A6ntFMlZ44adtKT//LuChCy5cE3SIdWwOIEqZD47z
WtEvk7ikqq+xY4lIUbykfFaCbfRF8XBbXr468SLuoTQ2lt48uGlrk6+x+opy
Z8PqPGfXgzQU2eBoCm6uVRCqAVZiuThqNkxw3iN9Y3hxxVQSlgRx6IcnTafX
X4UyX4s6ihvVZPSjdPKWWjo5U9zGqlqvzB1Jykdz2JgwJIF6IBBQyzcrga6X
LCyLYMhsq02ur4y5wnJPrYOmMmTFMjT/5etp6N5QNLRyg2GrGRMd93hNV/Lf
lRJ8EE40w8tegqBZ2//J+7Jtx24fzFNLYUxjlM31S1KYubeq15E4IMhW6Wew
d9VyAmblTf5D+IUgle9dydlD4YZs2+LURpyWOWPccMR0ur7XMBq172Siv0OW
F6h7bnDHRKoYqP1SyAJGrVThYZZGVOCrZ4p1K4UntERF6FXPIPmXTmt2r9uQ
FzrgRLCdY9AxfzQaU7tdYhEIsIumA5TEHo7fS35MVH3HomjOHqyUJYvZfHFQ
DuP+3aOTroGZSCXdehUbfyneCy+3u0+CxrvBjMFrBJPYuM9VDTxnXpC8pZzS
SJRCxy+obvlrxNZPwKbwSRcacIYsuWPZSG45hfFjJoNb77b6OGucIjx6ogwC
mB/AsEwCNaV+VIHfp7ZYMLt9lxZ3cPNYP44lLm9Rynb6ZM4BWRwY1B/vZMQ/
cgox1Om9rJ3tI5SDC4Z3mwXcxGzDFyHXhsMlXD9pSk9zrwLdcI992VmICh6m
ntjDbaUUUTaMKy7Y3YEFiTaxQNA9jJbYXjNNYfgKwSpFhvbFhuEmYBXsF4YV
j/fxW+QNgnan+Ld1eSNJ7EIg9RrmaM/PODRfPqTDBHHyZRqpTRg2U0SyaXQs
G+pq12ZYqmlp3HkXpg3Q3bX3KdyivwUGlP/VNukhGx2tCO+VwMuYiODIs1Po
tpxs5hzeJ8exvG8PDIyOFd1abCcHBVbs2GM2Rn7j5vOV3pSQ2kgiazzlGaY3
+WqjhJJddZoy9oSoFKf3mw3O8my4csT/HNqshlCbQNknt9CGuh3fAjO38ztC
JBYfb+hdrKf8Uu4cyzUnEsgELmUQ+rMWA08uTmWiop6PLAYTm6amYtbet7I5
UJMoD7z56QAXYR5ZuOfothR/WD4sZX3unm1rVXwUu7Y9qJ+VmxGLj36DDlU4
ZGPv+urvXwuUg0w525IVX4oTb48nA3n6cBsnmfwZpTNjfSlXbcIa7VXiVu1p
dias0Tj0kuoU+dKcdpNB2uorR8E/QLKTH/oFh/pXqc5HWcU7gYbwjcQVC2w/
5ZNi9BjdaWIp/+r2iGpLBuVhE944+fmfSZ8CMr/oerPrLuECWsqECEL86mQ9
3txf81HEmtcKXrABjBwwUbWaEk7LOwxH57ctVwNcLiiSR1KwGZP4TtAajHH0
tOF3tV/hsSwnrZPUwZ8V1/Zcx7PSO909vpKQcGrBh8W3umhx5Jnn8uD3DUpA
SjmnOA0473HEjosFZdQX9lPXJXLsguPTFU4LAja0gUnMUyEUB7U6ZUsLll9B
Kww+IqbyO0fLHdjG2NwV7YrHv+sTRgJvtw/Zsi+ObiNodqBm2X6ClfunFuQu
cytm22lR4y19Nh6DEWLkr65o3vOzqQYb9GtNHDOW9W3x1xj+WwofDCQLmkum
Mo7wRQ8FLkOhwF9ps0bhyQFYQe9i4wpaEXgudM/sB18vlMMsSOX+NHCUjvgI
Ob0vsxTK6UO4PCg+fiHXZGJK2szSJ9tWqXBUgGKmfhnLyobfvslxZ5X1SVgm
Hbe2UtMPVkJHMNrXaw3iNqo1VNckQ++3Y+Kk6ujH8L4kbbMzylBxCr26Keyw
bI6VQnHVAq5nhu/wzgW8RxyhqLtGED84nP/e8trTdlbSXumuxHY0yZp6mXs5
xXweld9J+nq2bCvILwL4iXPOFpeV+ocEyXXpcvQXzXsUSHXDusqm4mr1v49Y
9GVrUkA6kRQZR9lpo5+87gWM5kzFzEYdptndDpkUMfSZalyxFvzSydLxeI6x
zXfImKNqRG+TFlqW1VwBvd/pvrdEMZhTAk95bABRBJwYyhD61oyTGPD7NfGC
mtTn+xPSRylgbn1rlGLW9Nf2AXEN+V1d5fGsd6ZXuedk/N0I+k9/OtI6l2bV
e2EtUngW2RGx1RH92QtSt3CHC5JTrrOvU9Wlu8PfrcqMRPXjABzlT85mQ1eF
XtH3VhVM3Kh7XPpVpJRF6Toq2ZWX6AGaDQDM4OS+afMXDpAeVv3oL9FWSdaG
js09HBnbF8n3yC8cK21x/Hj8mrHugRR2k09FduAFM+CeBlhMmg6cjVtAVecz
mcwftRev/6+npG46noRUA9NWFF05cV/qNY4Bvc32HKHAo/vZOg7IhiWR2Oa4
LNKd07zFLObxvP22BJve9HWs6tkVLCawwPhejxGOSDEUPuqwW3VHxEW4RUD6
BnjCJC9YZoaVrpYP8932ThkpGP37Xhf9lNbAJ5OjZKuWsa4nTJXSTJ+uyTe8
Cq2mivTe1MQRb4V0SMTcLfHCZNm7kk77AHfQ7gd9/wPRllwtBtrwBmRvbC8q
xGkyFpILoDSvb7N8pDNuivPqtHP/mH8k91mJQE6esDcZBx/pkMJN5RRYRkJX
sA1PiOp1hICKUGZNk5SXOs00qWbz2ARAeMGffC2Gu3EBKj7rgXLlT8UrqgKp
qMoDUmaxWX6Dgio+VIdwjDdCxCNFksFDsRwUTtVQ0R1CYJZEFrSxHgmMdIsT
djdpp6oOcX9NNhgQzHpsKdgz5TmAXkGuEr6DhXN3RyaATA3QST3Su+RBoTZP
g5akoxMs+PDWQAfVp051JBR9kvy76dL0LbYtZw461Iso8xwxONQ5WzhuoCMZ
jkiYkSPEJ/knPmefotfEVdpX7F6UwqxAQsrrnL72Nx57B4+lvkwGTJ5DWOl6
FBbCjd/fOCHCvqldz4qST4d0d6yaW2pv5Jfd1XEdOqIvPKcgewHipRsT9bd1
nx1IaawmN/3gsh6U2Gt8mbS8srg67wYh9qGp/8vX9Da8dpEvciX9B2pucZip
YTIZ5HZT3g3vkiPlHRiM/MsHF18xDu2xVD5ZN/agb4G8gEkE6a143RziCgU+
feqaSVCDf0htQOe4rGNeZjLheEs2IzFeiodg58ZGdXK3L+y7z/01WY6C7+F7
5S9pOy/V/CtSEDcOk2J15hmH6RhrlWQn/7HLtF6vngOfoaPSOmDaE2AZsKaj
Zod+i9q6h+k2jQVltsca1YPPENcngImDIGDJjev0AwmiZ1KmY4EoZOVdeucP
cy/B9h3awE7BCYDF37wsHlDG8FOIiONhy5+PNczcbMkEMjwNxn68nq+Vtn69
y3pgpQshHUNM1ARN2MWzgsxckP5CaS5QTnAfd57VYqeliEgrZRKlJhOyLb3E
7/TWFF0vTSDKDWWoJa9DBCgicxA8BL02LdDyr6b6+0tajnTtdRkMUPRBHwrQ
B34bI/wIPrS/huHkeTa3D4h4BUCs3Rg4ME/ru/BHHW5J4BS0F2l+U2AtqUil
mk2ugE1ebPewyp5ayAZmAgzKjUv9RkvOI4+FI7luOIhpovjqHIUwzK2IeLk7
fdVs1OgPeVgeYY4f4VDRfLDUSCQlkg3/jrHIYuU099cHU1/OH9bzbLPqacV0
0qh665NsGWKn66B5+qbgrgoW2ksgPgyUAN7GfvXzPTVx4obRKcLT+P5Q1muB
t0NsIny+lWg/jMmr9zm0RNP87jTXyoIgpQOx0n/04YF5XUWjsWIOYQyQYApV
8J/WKod/SAtgwMjgAwe4P0nvSafeuJWDito2mWhoJDlAGurR+UvLeF7VuAm1
myMUBW9rTNPGcNmr87t53acuE8MAu0166MPW6cOvUsEqWYYWqm+pEmnXa1Ug
vtjA7zt/9UF+kxtMzHv9HqMAJqk6p4gUwpNw1KYdtWzNStXNYEN9p55mq0Aq
zsrBYGc2s4guAUNzRS+55w1mQDmmqxsnzVK7qao2tghMeKkrp5dGPVGt78S4
sUnyNLFhBOu8466taptej9FwRMyJ3o4gLv0ieD8arNoOermSmZFrBVNDbTxj
mIeWSjEfEWIhF50ugts/EpSQ9YazPfYAv+nGqfT3FrsiauxI5ejqcBmWi0Ov
6NOFrjU23xosLPf9vW3CuRdQ44vHJbAmI9BqhZz9J98VgfIqhiURo+3TWcQw
FJShRPKPICP9I1P0AY+oD7er5+b76JUUMDGAhx9toMFHcSRqryTnAnvZsmCR
x3t1yP04eKlg337wzrwa0zo/CmxjrRyKux5Esya/d0tY47SSMyiHS8oOxuTi
HsHznANDg9blRJDsiU/Lik4inTXq9O5NNJcR/EclQU8ht9r83887xi+cTXJt
sHXURNM6tmRz0Bnj82wDryY5QWJ5K9qxF2fqXrA99H3l8JNgnNv+tcEew9kK
05KEwJBA7Jxvi87XvuS0nrQ9byCoV754+wVUkVgD9OlY6/71mi9C2fxJ3adF
jAUc1faEJwHUzTeKbWW7KJGIG85vXh7SXNO0LxDR+ZsRl7YEaCDkPGO3/tFf
HN84BLK1u8YSwHjSvyiz5PRPIkdLJbcro1M3jdiuMM2nMTimh8SAe2T9Ii3W
6cRUULIkbJS/gsTA0ZbiqfX0J+V6ANHd4NdyHhQwe9gVYHLAGij4hvj4ua3V
mAuiKd270NbBC8YerbFfVSe+PNFgcAWQQ3FGVixru8m87rkevbscLKvPANcW
Ow7ZZAmDsWNdJBnHvfNWAET7RCJZf/zPap4mBENgl1GXsL18MDy/fENSOcnN
d5n5vFyODJGz9kaSHP1PEGKfZSWOwBsyagcFf6whfwcWL6d0oIT8bMdYXIif
b5fXuFqrwC1BW4apIcOTGkDMsuc7Vv9OtKFT8Ucs2K+9ed+YRPNOlFlVf2Bs
31KdhQbvYqwYoqcT2Bp+YNYaHzrMYKsb+bO8Yu0pVSkRG0F84RPwHZKT0ozK
0jpXqnsedNjykAUDiiFs90tW45fUq/q44siGoXE4AQxaSnfp8ssi+isIc4m4
Nw+mYusysR1AQ5H0jL+HUDSWg5yqPisbwOe0NTpqx0+LTILlNRO9Dksn8OOx
Rg1b8usMOMdv0RrebnXK8IG38KxQnAokk8dCj7E/y+l6UXEQSVeH1hWv2RdH
2w0BOmMvNWomUDG+ocI8TL3IcV3L1kzmZnI5P2rAe6aLxVWC6XioSEJO070B
ALw5UBHwuH1ctw5c/hBxO2KuOixcH0B02iKlBOAHbcM+9YVgjmqiYo1iGinT
ZrxbVhwCMTHGCwN+ySEMlTw8cFK5ci1GwDO/iI1odAmiAW2/PR3CpeCZnMAB
5QQRG0EZf0TP+QSb1ol1GSMzYgtL65ybkWxe52Th8IuGeVMp24ysb8FJdaAD
ma1sG8VpMa2iNxKNFqKwNLNKcDd+sBs6kP8WP5+lQPuiD3YR4TRuVYAEM4LM
v7DYDAwbiD2ReUbKXbfu2CwRB7l7M+/iCpabmkIPpfqMR9Mk2+0oawt34lUV
c9rLt/Cs0EZaDCLl6oaXpnFaIprp9xJyICxjspQe96IYwGlbg9LW250C/nQF
cEcr4ZQ9iWkh20mzOp2lKEtsBib+xrqv4X7z9LQUUmm46TYN2s0VFUKGIxb1
IGYE04EIMlbGZv+5qR29e/VgUnCo2HCKPHhRGhfWG8Y69CxxCJDKsL3ysRwc
g1XZIZlQNJQQ7PFwep+sVCIJRZYn4E16tJ+ARQqFnU0mJ3iGp+plBjszi9Yy
xNIHCswnFj8JanAZ2+jviNKzHi4fFFxa4hPIQsgZNPVtiphLC6m0ETpmVuwW
AzBAGd/zbS0C2qVqkUQvyR0wCPvyj8eJx5yYTOLYKz27IW4Fu5nyDgXQs+h1
EH9I6iyb4jRlh1WA9d1IMI0UOtWIDLl4ceypTcaUQsKUnguLPGQkQ6yt6RY4
2m0gc4uKbp13h2NdguOBsgHTqKJaWj3QiRYY/FrHOq4WJNyztkAtro9gMrar
qJ+m7lpzxwH3rvhFCg5h9pb0r2d8qo1miKjUY8E8NL6iW1OR1mfN/wiP1bUn
yz5uxVRlZ18Y2GigaIZ7eB7RxsHblu7yl+cJIOR9ZGfsvv+WuhJnnbjkEViM
tKwLOTcQPw4Pb6sIujCL5GZ03/IqZbMHmS45sVF2+Re7rH/zvAbbb3uS5Fej
1WvoGoWiSzH3bXp/yi4SiTnNHhcGa43Ympap3kJdcBs9HpqJH8xDculwLu/E
5dADQz02MUBB/sR+xL4+E7ZK5Iltq2QXRsNJ/2tUTJiKTp+DqWxQPBel5Rlv
RuSQL7VYU4c6NRUwIUDeMCKRuvivbc0DcivZcgBrG13gGQCG/8r0PNqD65Ig
2vzagDYiGITWawTqtWu9Df9ldicptX3EHonyjMh/YFS3cKXNM24+62ggiyRc
X1uZOD3AKrRFDyES/IuptnUMZMbnV6Scnbx8vCgW9Z/jN24wHilOWSD4dRHH
+o+Pe/phQewAgDaSYUYfbNwGRsBEAUnV6XUzw7QIzpVjYIUOoBUQ2zQ2OpbE
BV1tVWAjXmAxygGgSAFqIrY4K6XBpyQrR31ImCYsq0I5ma5rjhzmTiOT8TiS
cb2mfbem3Rwn8k8B7tn+3big6d71G1mrPXboPn09NZrBXvdBrWy1mk6Gbk6K
Gg277wBmgGo5c5Isxt4WL6ET220k7owJr7w7pjsMhyQR1RrQsT/TLrnlj3pZ
JyGy8/udci6JC95F16y0faPbUGYa9mvueR0Q1CHPbqCYR93zqUdEacP6+pod
Vb32S8HEm3FGEz7yU0Ea4du6xcsxoX3JHe9hjx6+n1lZIsAlrdaPFNbLMQz9
QoteArkc6F9JOHc4zUrtAbwTQn78HQOgwb3+pY97TXrQR8pwxYFdTuByS8dx
YY16ahP03eYcvlRgT3LpJhCCJU9sGWbwjkPEVcP/a1uuyZBy9WzbhNbcMTYP
oZ6kyeZ3AiO67bBeuhM+90DmBucGNXeR3x2ZCiPaWH6x+MMewwAQ91efPHDG
I1Ti7MtTUDKM64SPEhNR5rHEs9RgOjiWo72cnYxQSpJxkTmZpWAB8z0ZSQKX
s6JYcT0vMomKmVrxG6wb0SDTlrwdrhdRf0BZB/5MPHc8iH1f8jz+5OhG+leL
JTH/T2NrCi/2eAqDWANraOSMT45KQWUT6UGGMesG2g77E+V+bdqVoAeppI+C
6P+Ier/0hS+xUGUoebEhrF5SHK7ZPLGyt837wUcx1clWH/kGWwiNFPdICIpz
ng8QaHyVPiIhJ0VJdYvaOdChZEXGj0bJ9xHdy4AP9st4+uzr3gDhGynNcItP
HX/LslNmc5OIG0BCFwkMFjMJiA8HMm6lSs5+i6zEkxzK2tVkz4zRyQLRSFxN
hEuwFRVYeEZKgP+Ye7s43miwUTpVO6HAuAdzqhmpLD75iinnyd37ANrcGv4d
n4kw5LLPtIHkC0fE/qohrQqnc8y1d3e3SdKEIVdoo1pZxD866oG/c+3d6G+v
GCiJm5/UtXG7iekebVL2HH0ZuNc2KY+fdq6hRUnXgIiH0CMgLYO4/4JM7FtI
cibopx7khiXtzQaJeIg3T2KvV5rhBOMI1hQuvhu2qqS5Kr97tC5YoKobmrcu
8eHZ/3/RMcJyZmIIcAYcgAwJKC2/XJBnXCLikkkDdqep1oXwBOhkJHo3POwD
6EATMQj5xXLciIVmf0i7xdm6sda4b9ylAfhX+/wCJH95YQP8V3+ekX4cS7mV
D9RKBoYpCJKh0fM6chcpvGiMQp4+H8JPwZhpS2s7ffETV1EpnXfzSAKM8+Qx
fTVU3vY5bhc2ZwYz64HIxfY3CpuHOa0omTtte6atp5k7eeTWI9OgqI8aLxrV
mEW8IdN7AycKXCzuNbi5xjuAfc5PUpyes75P/ny7ulUsfrfPedaYk9uBzUnR
wIZbuMbhaI5y+eU0WMS+wEFzyZacFZrLYN+UBIRZv6aSdK95k6JuRaBzaHcZ
D24r+yRlgkvAC1LftyFAwoxpzBgFvbU5Y5d4MR394x5XXyCX871J7NKSRL3a
LRHoHd7Dhc/1um1ppcDdQWOcQVyU+0oZOMUEGPvcCLFwmyEroLmSKfHult4t
Xpanho7oXE94XGUTOxjVKTxvYUgXfPjH3asleCod4RCJB3zaOpjApvOI3x0D
eI2mdTGoZJxVZFOqm0uN5amfswqm0Ohlv9WqUNm9ZXgweqKLuZDoWZu6oa7h
RUD2AHqVVhl/APRLec3Z7ySpDArhwqNd13RTm86FTDsL+Q4u5X/iJgqDuj5b
WLi1M28DrzWrbR6TMK7Hw3XWKXzx5FD0dQTpRg0P60H4tUvqabTvvvIhQZJc
1m6CWmbQMBc7ooHVwqBEA/road5dqnr2ewxJyS8xJUs1RyTxyAtKIsBtMjt1
L6TKjV9dlwaIkSLjkfkf13P1zn2b8fdZxs4kzsqkb3ATsO3LmT6iAOcuRTca
J0on519uSK+UHHog0rwIqOSVij5oZ1Bhskog8C/LIB46wFOzgk8SyraiDHir
UVgs+En5gOyz0/xrcJDo74YzLpW9dBcDpKqyrsomUYXG72dce4LRO/iZufgm
BEGXibqBSb1H4coos/5rBGy970uCGb9/i/Aoksm6nWwaxSx/BKbBDU9E4vB6
aPPzSYPoI1tmRGreMM/fk9wPAnnFuZmG6op0sN9ouOJyVt08fBaWlW/IvF8c
Y/4Mo3J/S6t+U5GdMjLAyW1fOxqhGOC7uDUl9vg3YYh1JuZEKDY9JBp2EvHZ
PNuJIK8ZEDbU1WG5lX+An42/8EsxN97SHfDwxOxDgn4by8uVwQk24Xj3KEez
fy+aRn2rcAX45HlF3yYr5pHMOqJP4Fuf90kLNu69R1AFPVCt+b1q4VxggJO6
1kW1vhhDajay3fd880+xI62/kAYrDiwdZicphMteO7e68jD+wxnOjQ+OB5nL
RvaD8aM8FfV34I1oAkK085hYqyQkY3M/nwHRXnsWmXdYD99CS0LAa5wvzxrX
fG+I2bLoqwaPdqkXH3RzQqQPUocGbXpyXEns6xuzeMwCQvnaoNgXf4972p1e
72yimfDeI30oFY/5llBd2yzux3aoY2a8yJD2kD2KfkaYnzu0C99Xv3bTbFec
6+6JxGFxf3ItVAWRTljJtIyPxNR6kH93l37+5Tmkwk9piLjs+q1yPAf4kF2V
wg/84+74KrsGgJ5nv2DDPqiGUZKgNZ2FNUujh3ZSCtlP5xKzdKRC7sZ8cm5U
9R2xMl3rcCIAEQiOzsXQb/mX3B5xfF/LW8XaMHAu1AeDmol/K5XRmAB/qf1P
6OsMUAahX57ptmd8dGVFY+0hlAtSLMBlGCsYFEg+QbAE5d9LZIlYKpRqyqGV
d0hzvkboeMEIv3OsjttxwUCWvpi3lg8m2nuHK4FY/CPOjU1cBvsGFkceHNmx
h1JKd83XO2YfrNFq6GAXaZ/K+Iy264b/9TXZIoyvqEhk/Z7G9PrR11c3FIdo
NG+VsCWrCwg4LilQl+aAVpflQpsskrkwH8H02TLXA4StqLP4ByP4+VgZOL9v
htMrAcPvWM7Yd5em8I+T/M2ioa3CfiJeZ7wx2U7YSbgVxN10wPk0hhZ9xedO
wtAL20YPqvvzUMnOu2zdRLwPQKimpsrLCciUyGM48JxtCO3xiGigvtq56rcj
yptDw/i6JVilAGJQuLrwl6+bcRhMTR6srAsKz2xQN8X+io+/NE7J52qcbw1z
5C4kB64GIQfJo8r1t0ww+1yuHvdxsLUUUdOSehvowKheSYZ/mSJgbNxg8tdL
CMqHGUTYOna36U/dchYgLz4TWnSbNZjzUHQxQGQEI+a657YTxq8LbRSXU1kZ
9fFhxyxIDzuwvpEQdNHn3zt8Bk5xyVBin3uibLWgNGFXgSeDm0h8M441m+mt
/4KPYJbyoFyOfsMk2+oaqXI9CIKIj4/vHfy2XOEfEtzLvKLgvoW7DLlpYCTr
tJptUxF7ipo6wrfprltnsHPqiXIhvpoPRKqpz9blA/WAUTA+kyyOWGBUfJuk
yrbR49A590cLP/89cKjm6Umk3p3chghwBimnB89TQkvmF3DB2+vXZfuhYNKP
U/TJnSu/K37lNkeXQ3jylaSUi/IbhCwySVEvCRWH287Sx+nQe4Y734XKD4iv
b+PhdHf1wz/2wFgt6BqUSh/TMK+iWrQ05xrhUiXfdi7nCnUmAEMkLRbHKDv3
3cKmB4Us6QC9kAovDAsDYFHMt8+zEjI7Ipd4BG0KyXEGtht06qveeakIgsD4
sPorlv2fAwPgk4xtJsxjaGJsexaEc6MGKe63a8l/hxB+UBSf89qPYMEQ55cM
eMgMSOliCP9Iqrqv+hhMXUXZcCJoJtWZxr1nE3Y5vsGNmCTBgDdT62ctrrI3
XvyH4lvudBAW255i122naJgZ0kJB7+FsAZdeXWgTgVXkENrL8heilVaGWTg6
kfBlpxo25PeTQVFkZJocUrb4pWNxQRgMFzTcyC2AcPLSVSQsLZjmHr4xHzFT
ukZaj/ZRuPi+yUgaiS3qGc/i44k6N6LC3XeF0PrcakJ0OB9y07NiPdNdjZI8
Rkf4sRerQJFe3yR4MzTr7xcxcFX2Bbit3FU5UvNTzojeJYGS4II6EHoDwYFO
wgGKUVgmg5+taie/GBUNkUQjYG1qS6Ylq9Pi2AISbcfbtUkNPk/W5Tkt4z47
ti6gpOPkOaIOl/HXxoEz+5mhg59jfhMJIfyhZ+L8UCqOiJhLDOZE/62klGQb
ZoyzJRh/eFMtcdZF/chyaEIfj4egh6N8nuji+WT1BmsDYACLaOhifCGHAI9P
JoVHfzm33y/nW4x+sY3PxEYI2FfoKiL27zfAYk1ZWyNIkCDZak5hDxlaFXXj
u6mGaSLA3Y6U2n2yTlEwoFSpATltXU7emW4OALJwTIekTb+Vk2WaUVp+bthQ
sq3otUXagjXEwAiSYRXbJbt4syYh8rDjP0uuUcw2m7JotW6GuSveEd3Cy8yN
REXJyd0XyTxNXZ7r6GQ8sLGE3Kjd5CnB0m7vJZrsVpkHZOArL8m7UVuo65ec
Yx5pqua0eS3IafhtGIjVecyTFnxdb0y7rOmrpJpN5JVYjJXar9eB2B346otY
dBAZnZ/lDfdhLyqvvA82TTmG+InyXNU0wPp7VeQDs5YiyNSeRrknpk0M2pKT
WAkf/t60CycH3oRfmV6hXfjyl7vIMirtkC/bVwr9+NjIo8lnrfzdLvqML+Ct
UyUxKmkh8G0Gwd+yBKWAGeIzSgVjb45Eiu924DtTcAHyFJhEcI+X77PcR6wK
ektFa7qDv/5aoB1gkrHUiQ/ozsYI3zoBQfSuOytiNS92Ty5ZsjAAl8/1dh2N
IDS4xbagxS2PxmnhS5k2tfICcOQqLvL0unQsBZ/fwgEZOetKSGx/E2KI2lEw
MJgvqmpIwQRWq5a/hebLiPMUjn82xobi3KIIlmHdTpQ2m4uzTHx68CkoXySD
FUmyhyNpRmMSozfmwcai+v/1Sa6rdWx5zC/gMIshAx+maOioXZU5ase6/Bke
ejqawydLSr4fFpMOFTUuNl2aWw0Xv8k3U4iv3CD3keqXo8hACwMyln108+BZ
TUuREil03Xa1WBaDUvic9kRjEf73LmNAPPKMp48pNKWLQjTTWz9o8/LrejHY
Rp84WMuOxZf4OeCyK+om95o58m1WOZJH5yg16pjzd5uXfrjLVpkiHLn5ORSG
XSBrZ98h9GnI17vbbDJWSHN4EwVNSL3L6aQvivmOGz2Eg3XmqPK8pZUdW/mZ
x6H7fn0ZMgk+bKsja+1Xx1hHDZvDQILAcDiAoCn8P1Kmhrf4WoSu71XjlM/d
fdAPJodhietkcqcIcd+jvcEr3LelVZWG0sen98zN9bM1RQEpWCnDovtwyHE1
/erihxPS1g75njSha70cgkm8Gg2PCNkS8mioRhmfTK3ovJ0n+nPpSPmwrO/Y
PSdTJP0D6xkFu4MGWXMbjlx2m3z1rSoLNJ/cykoKbvWaGX+OI+EY9N1N1V0N
PYrrHwEGC8c3GeLpuQzgt+zQpwbkK3Uv/fGgXp2YIQSXBOB+a3+DT3YFH4ZW
usuQrJphPM9U5VnEkma96b9x1O/+jppoqG84Tnqa4d0dx+SUOgb2++euaTi8
ss6kISqMHL8hrV3OvhUml2kRY7i3cRsFHVNfRMOeItIo7tmNK61pfYNf3N71
uujrh06Bm1XG2CpVR/EgqGNwRWdMgbsKM3DLguLR80XsrZbdknhT7o6ZVTmy
zgbwFg6Abvhgg+myPEd3tBWSPEGtY3D3JYT1/YxG/aDzcMDhGn3Cc9GTbq0p
ZcSzTDcVyjcgS1V4IGnwX4R8GMoZosyjB5WVRNeUn11HJYI60dAd1mjD5DS2
Uv7fXbKYB4oFojHTOwRfSnULQOHzxxYZCFDKNVGgP28Fkvb8Ihm5pVkWCfXb
VebstT48ulIwhaStx+f/czEVTcyl+8ZbY2W1njwGF1Eppii9D7O7LzssE6/d
K4D0dj/H5dfcbuwxaV3Pci7SFJGxbdAcJZ+brrGsJA94QveCmp14SRlX4i9H
cE0G8L3Fa38ZJ1VRsW2O3Uj9rArn3HZ7NyM2XlF9BwdzWtdL6Vhj7ov1dTKp
zSzf+JR358v2DdDAkBKMTl53GInj6F/ct80eypa7OPpyimFQxZXDD5PaMOH2
FBLwcgyokozSuaFNIo+7s3pd05q5srUmly70sUKWtMC4UKqt1Nmi56wqa5Ic
Aja7dljNZZWtAovLzj7lMbI219ej/J7kdpHD3BIOQ/K95ddKXViXecUBkoIK
0GkSQukjJnzfR8iFdcTfDBtfo++5NHHEr0/c64hkCWlEVJKYcz9JrttLk4op
LL4a+RpasjiaMY8oO20Z0GRCRGyfuzBXA73xG7fmrCPk9ZWjXlhvkjaeuQUD
eMbKiT3ZhRMW4NAv11Gd4tNWO6ZO/rk2aqFJZalH34nAMhoOExfU7n5jEO6D
uv6YqGeExyfSAFrvCSpscn6wry993hL6+7xEc5QGzr4wS4jdCsOdWtq/vhaG
BMJAnpKIaNgPUKZmnfTY4tfna1EaJVuvKuJN8ZwSQw6iiUFNiNcPBMn0mA6W
AHRghp6mWIf7rjNPMldiOZNaBXNHoB35aC8fWiG8GlNfndSSwcmDko31VvHc
V8Tf132qLUgO+r/HCc4snUSrZ8UR+cQ5Uqk0fHIIqke/cPF6QynAmMezlVmO
Vv6L75rxRnD563WqDYgLwxGIAAY+OLRFXQiiRgg2nWounn9XbEndPjxaWxFM
EzbBb/N8U4Yokvy+b74Bnhn7Rjp27KaOHQhl1Wcx9EWsZFmKic0t3UUPryoF
nSxkrlOYMuzWN4NVnMqCH9hYkdCtok1UJY3VOMBG2oyu84422SzAH8gYZci0
5g9InZSlrwr3xldeEYpNJNhmMYoKmtssEdxWzmGuUvffCr9yc96ZT1GFbUSk
YDHAstEafD4eZGPlyCS6kzvnM1SWonpDltKVe0lpyLzgTvivsE3CxkPqkz0s
UIAdNUnmi0Mt9sWMlRvM7+JYX9mInzX6bNocaSoYjozY1crHXAKgILhGVpc0
Cy5PMnTf84xMokVAUpr6mp2CYsrfbxFX6+ydf3w0OsnIy0RGkw+GI4ltXPLX
YL/TAiJLoEYe5xbh0GaCHM5puUPkAjiiVRGT32wFOjITlAaRdJjiKS1FzV0p
SKiIT2dZJ3lVZR20Jsr8iBXc37imP6rrfk38A4Srr3ZD9X+VDpYZ+IONVpE8
WjfgeDE4F10blTGM0RumnERN2QjD1kYZDlXlzvrLIi9zct31KT2jMLnGwaeS
9K0+x+xN8I3NMwUP2trX6WzwTx1Au7VVfsrSoVYUkD6LTJQnp4y01M1Id1iw
j23AP7ozP6crjwP5wmbWVJkn7nYXRjmmdSF2x1AhsbPT3ROcgjoi4csrT4x/
AqG5qKCg0vpJ/1GYDNh+rMvam+KpAdPbqlaIL9RhmLHZUtC8o8NTtWsIVx4b
KRMdR1qozunD+TtLCMgjiQ+ACCc6RzzZdU1iJRqespkqGNRtX38JH9tO21J/
FERc7HeUGf6ULpYf05DYLFIRWVr/P+4Atqlx9MoyXJC5G34rmpfvEdcc0EtZ
ySIOoh2sfZTRYgXb1c6nhbQD7zbbBROIM+mJ+Yerldgsq4ChRRg0waw/f7wR
FESpNw9Q9UiJ5vceGsdkSMNUyVLoSgS/+p5anxV3XT8Im5w/sMxtWfwW3qc8
wIcdlhFENau21tKV0Oe2pxBnQE2f4Ki83gqCVVepVMqLkLKlRALGNXaTFZIk
6emOu4djazaZyvqYlIIsW/gfVj5MrZOQxx5ybiis14GU1KWvJDZRLezlLtb0
3V0sORDLB4//4pp1jDwuPF4w50kbgTKnKIQrTHyqXh2X80yCbUtwWBy+56dF
X+plLzDD1Tl1ymlgy8l4sr0NqIytNuNOUZaLt6mIL3ck0rlvoyAPJyUbWCUa
PXb9fk7eMDzkw+Zdp6O54IIUrFZ0OWyeE5xksFwV7fOI49jjYyIMw9V8VPpH
OZ3jkhGIlx1g32dpjiE2VdNIV7UaXDQli5VuASufj/d7GxrMWIMIRVPcvdfI
hLhGCJOvH4nCbW+euEkz0YFkTfQVNO+HIiE2dht3LP7DgyOisOjXct3n6Mdn
bfkkJp5jqI+Eh6V0+2e3YZ/GAAejyPVt8dRGbGyuUjlj9+AYm1qXyZomlp9R
nR4nbjhltcMC+0XUOH6tWxxC4rq7i2qmPyDqGs7UGlV69+4tczUDyePIGgHN
yKrW6bKhpKByvj3CJoTlYFFGCsPZWDHknEGkqiwGYWNGMsY6RNVAPOCpflHr
EGx8x6KIzgCxy4/mRDmMMqy4DkVYJcRQesf8W/LkT/OFRRHsTnMhN9SBWP8p
LrRvu6Tsli1MHnSrjV9znheTqWtD9PKSLAecS595yOK78LFJLbu0A3Ru5qqr
rT+grC2NzwIvANQwzhhIgiTKVMTRWGbMPMoHmD5JBKqmrYk3KXBML5e3rlil
P4BNvXhkvYLf83MjAT3rlYqOB19cCPPBmxrSVIK6IUW2Df9d/EPWn3zFKBTE
6Y0m4EIBDcVztU7gvksgh/bJV8zp3jk/I9BFZfbV/aHQL91NgQyvQWcOWmcE
mD1Q/N+1pXcTmSH37m2k7jjDo4aq/rxM/hul7/YwXyEZGeYyWerKTLoBS9ee
+nJQNLnVWz4l8ffOkOmtbRc0uJjMh010BafFq8HIQya1za4vGPMht7Ezpjyl
ac9QP0Dmw4/eUyUjM6NoDZsTkNCIqkRmzWP3anSWr7iS0lSGn8hKtofMwk+p
FGNia95UYDMPfihkG9ovmucwyU6esKmILZ8/f7LAa58R0FPxfzme/hCj5l7x
dc0AJRkoKLpky9A+JIrSymG/ljbETP+l3sYFxZo2aWU2IMnImI5gCjMOqjG3
mDlAE5WcMhJZCwMwN7ENkCiK3VqfIPO/ux74w/EwGoIm2rygfJ3uP2/D/kFO
Rdz3kQeBz9+rV/Jd7xxaj3bkBBy069WEQ2UqH8Bgj4CIqVQExxqntSkNN71/
o7TgIcRV5HQQwGBpnWtq/0PfwUkciiXgTg6/JshBzn+vztAPPOlL6wLlHeNi
7JrfuZ2YYl4VLqz+KzO5EdD58DjcLMc2MXjIyVY8hMno99VezBpDAt0oupZB
t+T6ZocvntyzVKGkfpwEbvQudMzeUB9gyOeal+Bnd6kwjMnkPxbqKrxNyd4a
qbjspVM0s75W52qgFgafN2OrD03GbkfauxAqFadcPltaugmKV+fe3G/o2cfd
YHoE2edrTIjfqvX6xr1iTP6EyugvMpCoX5v/jFIcJw4ZjQWtRfae4wosB42X
CLDQDQsDHzjdyemv8Ks+9zkdIekk/1Pox9j/l1n8YBkSNaBbmujAn9xPAh+g
HZDW3OqOz+NcDY398Gg4zz1gx+GJyPBJwH98TQ+lm+AnYCKdXH+WGC6MAH82
E+FCv1693KhFDq9pWFA7NUf16J6T2ak1JMyQo0sB6SnsQUb5rp4Ca2uBkrFw
YXff7OVBgxj7RONDcnikhenR2LpG5SxoZzQFyGWdOoiZ52nELYYFHSKYKuf2
GyVU53HRhvizhScqB6DK601SkQovFl22IKIn+4G3i7/zi9JSqurh43+g6Eyg
HzERnA7LsDv50WeyePAcSVG3Z9X0aeNkX2ITPgF62RLelc7GceUrT3sDhrs5
5FCOvbc/jseRmv/U4CBOuHKCRCaeBsLo+HQIbaKjjCKCpTSpLXzVRmWo8bjw
Mr0AaAsIr4MPpQxAvkCPFTIDEHSbjGh62QLODSvL2VntEgZvepOsLnGfyffz
s69ipWZ06XxtO6paGLZrm2qC37W3mJdbfOdLBh/e13naxVFsAiVCw8A4i+52
Gzy3xWCYPSDDWUAS9nbb23JF9I4iRicfzvoeJzNYo7fpUPPtG+H3Nk50DiNr
vHyMR9QZ/1VoiFlZHiOTCl0y9sKBH0qGvNueTi6tSydTh7MZDgiUN4LNKJ6e
nJUrUUVrf1xGdQFJKnLOA9v9KLx///j4N+rYsYxgMi8+xGed2WMnFzoICbXG
EgNM7/y4LmdoeiiEDvixR1nnIRV2YKO32bCa3/a5owlH6n1804Njvb/l+i1R
gUQxH+WlI+YzcUCNLZQbZH9kkkw7KT/nVNVwSqoXWmYGToacXOK8EnxM/G4E
DMr48CFTsxuKLaF+mkO5WXuykBv6IZxjCP+CCSNIkd5T+CQHdtPrA6uEUMda
UWODVZfZa/j29H2rVabXJ7EZvw6Dtd1vuPiBHzCSO9hPXoi/HPvCk3XnA0c0
fkXXxrYK6zyRoQzEtUf16cq/y4rq2+G8KzwAIW4wTVXhk15Lc2QZf/w57yqc
nom6E67c7McDSowI9PYrCCLigVHBxXnLs+Cjhr8cZsaKhdpqscHxvfXpc/Qu
BUr/paxNBVPR7CJ3Cq2vEosAUXNL/4kXpmNrGeEtnXXHvlabirvu9FY1gkJi
RMzY75QsJN0Dcr/VzjtDOpOP7TxwrHTekuHXwUsJok3oktcAv1cxlAis+ynv
jUdmF2D0iZeW7tdRCE0duISYSWcsoxc+mPStx2Oz+olFUnoXeXdng4vNncgH
9CyrCGDxkFj/VNugQmLFiicu3UOXpHM7Yb+5wai7sUDOZqG+z5EZu80J2s/t
w06zidbN6R0BSZeorWpjo3YsmKd97TEAH8oSaAkGuzRU1ta0PF/64MFcNahw
VYZ+v/5Q/QpOu0dXiVsXlRLdEYpY6JYCYkI9iuFWVTiseHfmC/y8P4UX6aoN
0lxEi6gIWfr5gTIwedwZHsgGVAa3GtvuIqK5u5JbliiDKoM6d77U2FroCPTp
ftSzXgF4XG34kcG2YVQoqki5Hmx5klIsaPGDwXLWWznLkg/GPUFjQm3GRla2
Z2Ie61hKTrwMWIdI4z8Ddngy+2aII2QJ2e8uQoWUlijXEgzW3M5qQGYMv5kH
OxTB7x9U5GiPrBWDQT60YYcU1YMeq95BJ8stCC0zkHCeVAfQrEXv4rL9uryF
hYEs/RLelR6xo6vP9Xpc2avKJbNY62jiEOpm28C68YNKRCKgIiCVoUha/6Hk
f7HDW6hzMxXZIpJeYTmlhB8+Gi4r5t+2SjtdIieQtNFNC67J9CRwK5QpgL5m
zfHIll+TaFLQDZgmeX2k89f5/j2JYd2uShe3Q5su2vpHhP48YlOSGjGPBGk5
Vc94BV+26uon4Edl6zieHiro+zYpWgqqg6+jh3ZPvd6qApQ5nxkTkS9IbvZx
92J+mKugRxjgsssTWJ/I1Mon500DewUOAcJHHSX6SEvwTzjWb34cLzyoMKLw
MbQToSQz2KcB1yoB8xkrA7a0tZR64TeChKfI8GKS3uBGUj7xQzbJTAWk7jLp
jOwZRwBM1Kae5eBsDwr5NlY694HFU48rhbT57fKpxzjKRHNllw1fEOu+rk3E
X4kmJd45V/uUnErhFFVY3UeZiMiFV9ZJ47WJHF/QLtjMwQ4JXzxeYrauLjoe
dSyg1qVndrvAbs/3e4/wMYbiBzMI5TjHhPir5ANogyjUipnjdowYjneKFAfo
XRrqAj1wKn/A6Kf1/yMEN+E+2OH//R9s6ooY2QdcVT8at5aS0pQ2ZFNzXX/V
tcEXaXWFOoeBq3aRhnSEdiGhwi8EuF2oEEYSYgqaFyOi2gQqlgDSsviffkQA
gJVo3HtiDO2AAAfvrEUMHavQ4kbwryLsmfi0Gm5F19pK0zJAOIYudYm+ozv9
G+ENdnK9ksWj5MlmJjX2Alf+wk5Zf9lnnvOsUcez5wW3ocqxeT/iqWEhV9v5
9V5PSSlz7K0e+EzSwgQkWcRNmtdZY3VZbWdxcS29Lk2giu15mQAl+UAmCKgG
iY2EBvllYRyreSdftVJvoFzaPxEKHgS1hWXW0U6nZPI5ml4J9X+WPgIQhtCn
zREFDbVKFPblYksg56P1KbqXDzE+fNsclPMLtm1Wa+W4yNV7JolgnI0NxQVt
04sQByvwN8zSr9YBV8rf3nynFS03UMI3KE837ZvRonGRVTy+8H68gwDRBiKG
HfD0qQwWojk/tPRVupqKNoqd1mlkvo4fy2CDO49kXfCG80RSA1WO+gWeecWw
/m3C3WVKLDi0oD/GcH2AEmX9ujHg1ezwtWwLES+EJYLBDyD7d9luvLnOu3IH
7UsYaLLyu2eNKhLGfzMPFCScvhsb9/O1cr64iGuSVfwF3MB3mICqmVrER0pO
rtrr44lUDgxPCPin6DdOA0+VEGsrjMwZb/O4AEPxQ+nrVPr3WBmMYrQFjP50
D0jcTLjfk6FZdV6VF/PXor9D1zBRp87cnAfvbm/BLfFL6uO972d8RVMX1jDM
gZmc2Uos4dGfLWb+KAPK/RFzDtx7yVJBRreHf3Te4Ka/2vVwaHSXa+Y/cH5T
tBX4x2ys3WOw25Bt0+JnocFOoFja9lWSR9vYer0ezMTVZwTbLhheTBVYgN2v
E5QXQ/fQdXEjsFZXUBf6IEN6R0sRsYyE56jrN+v7VzsrXbz5/ePiPj5ndStm
WJOQdVCST6E5+sBQenT3oUZkNLPu5rjRX3bb3IAbDP8dtq3g3YFQA2zhJX8Z
87WHBvRDycfkLmojzUmezyrOfPE0MxaOZmbWBhZlRAxbmnknsTVWqF8amUq7
l+D8wZ4QCDCvNPWf9lo0McovA2G9CxwCXT8l4lUgz50D+RIczXUDhpTRiglb
bhNfBrBwywov+5wKSUwLy0NAGh8bSsumNnCVK9xKZtiB42SAjfN1x2hEGrDV
RVdZuQ7V+ZlDdIr4ceWkS+W4keODWnkf1tmE5VO4u8vKo9q3vvP1MZE/KmVq
6q9fnKmxTPQ2CBIsA/vhesgRbdo4PH9MijbXWuB1AcIaNpKYfLtfFXHFjTO+
Zmum0hCNvRSKJVnTc7YzeFVvhko5AQ3TOhQAWjFkspiL5J3R2YjoPkU+D7wa
ei6dgi3oeSalRf6Bt9uiSwDTpld/vPfcb7Tbosdz0xNPpsphnxgDWlW+IceN
k0lvtsRsii3zURSHfwhfCLDLu4kcLtD5RcJmws6zjMZeJZTmLbspIV6r5l+L
+/jSGNlNDNS6M0MNfF4wSzjYhwDD6ijTeeVf2jEtUr6UInYhk87TrMnq00Km
y0q9PhzHayF4FcPlN8oyxkR0V+lXCGHxTNYeokc1p3wLYUMcR53kiqpjaK61
Bp7EHblO16iqiVNgnY4Yk5splqpLhNIS/S8aZKj2+mwXw/I8xuJZCCTdDx1I
di8l3Y+wm1COpPpxjMkv5PJa9DAQpn4Hn+hBjAUwBb5fmJqg2ERhz4rjHPle
9/DhslqubrhIi4zmvFctuSuTpQ2UlGPm1qLwR+2D+6KxqtA9jcnnUJbA/wbK
sxJYmsrFN2li9ajy1bq6u/VVnBPm0sS5SH5PD7tKLcvOCOx95NFRZ+1bqd/U
rsJm86vZqQPuKgtC+8F4tU8noj0JvsegU89cwQ2Qgp3WcTl2Yo8kOv1cv5t6
MwA0Ci6Qp3jZKAC6q2m7u0tpeVXlDzcP4mRHRVixqdfg3ZwSCb5ua1fnE1ps
mdd6ukgVAug/ByyBd47b8bTk3US505J1H9F9BoRjHVO31azHlydM5SITE+3F
DXWO4VXW5M6Nkks9O2gUxBT9xymTot4DiIDGUrmOK6bFK78ocA2F4FV1qK9F
nraQFuLblNLN3hctV26XkGjw4VSwlJsrntPM2sjIEQTOLAfffPNV1a2oQzcX
JYqsNJh5JVGlkhRLM0+1ogpGGZUC/UIo3I/sSyF7uAdCKbEORG1tGufC9aFk
T4vRbbWIZ43GVBUS8UjYt/wMP1KeqpcpHRY1wqWjiAvdyydQz8DKxri1tDpJ
h8FeNdYATW4VO7AcKey4J7qWbdKvPYpWWI8uC8qYrs06YibclP7gD+OIVvwY
ZzzoZ5FRfnD9aT8uN4/hx1y8xMdaJTsju1NGxLBaXr37bt2T7SfJT7v48XHd
1T9qfulf2bpi4ZT184HYe61w+I3d3LLhUSepuUXqJRfwMeCKw9fMVozJfDCT
stQIoTaRVV3iseGDoadYb1RetqDIMYxcjK+j+Qnd8mr3YD/xYjJfB8UOFUvC
EuaZxJX6gl4p4XCdNM90hgosOTzb9O+VuUL8ef2bT7YTnTEkmF5PpC4qMfN4
FJw6sz3AssY0UrpQlYC37Wo+APTmx/z/6tWpl+9jClCQDzUfsSPs7To2pRGD
pgh3bPy0D8uEm3Xm4E1Sp8pa92HHFbkQyGvOKdpaRZE8T9zxXfng5wNxIdLR
Ggi0jubpLg7fnYmnrgk8t3QuVx9geN2TO8cjHyfaueLd9eCmqR/jtF8Msm4B
2GYBFo4MsswBbjlt5T019WDa4l2NHwJPCcHUimraC0GvFCQbg4kYdy/A3GwM
LpkSeya4LpPK94l1dRXfYFpl1QvbQ7Bf6vy5xeXsA7GYQupcCOJvfCjkcII7
VKNJh1iqnvhf3rBZK8jtr487vsQWTIPsU+1aJIIr44EMG8mhh49Rstzd6t0o
EMXAMdqwdmhZmmbV1jAFMlTr/FRZf755/tFZLlZ+IAwtDN/rWR+4jwz+IYIp
wUpst1rF0pvERe+E77NyoaCN0pYbQ4+LbVhntCbPAG4X2VwyhfPYxGl9bFDd
3vsiyvma5Xk18nSIbeqvQ9Aohbkn1PecJbDzkhZIM9XNacSJ/OTuwz6F6XMJ
HL73Dcqzz/deaiKRAbj+MckxdhrGmDek3wHomnGb/fXhpN3iGullC29cC4RT
83KHIdwaiBCOZevOvlODAPZzz7dxDezu6aJE2rL8dMz16Gj/LLEAqsVYMnxE
nxDy1VcW78qJ6g7fKfoCiy+/sYOQOEabVFcrMOfAOouarKxNzb5jEFFMTU3c
hi46otS/fBB0NUuyAJs+zssjnwHR/JLR2B+sSXMpvTRyrVGP0ryt5UfVVDZ6
IUzBa7112sAgeDunpvHVWNiqdN2FSKRqdC6Mqu/zA9j9zk1rjcjNAcYXBh8y
yLWOe9Z+Us0Nq8h+EIu8kc2BWXDbdcAlBx6UpTQH3KHEc7VpsZctO/1fdkwP
W2z/YvevE2ogEiLLqVv0wI8Rm1UsyILQ6rL4/U9MKeprsJPuYgXMj8RYohxl
FR9pBX5A1byna35qg1NzTgjNOXnqEvO9guWAqaPVFEAjXVDyTuIq80cgQcwD
0Kkn4dJDY0jl7tMnVV1Xh8qsc2OM8jb8/igymZkahLiCW/IYdH2/QmsHpJmq
ILJeXJRRnIT+c8EDZJWs21qHuFcJ6VFxwb6UyKAReLzZD0xjx9/I5miIPI8C
ioc9NAN7uYeYCQurFdrGnppxDNDTiVbChhUFxKjMrFO2jDY/yk7xrlYlZIJG
PsSNAqCwJydz7pPFsiTwpD0fuFXfDSjKG7xj66SvuqCy2XOIUssE/wFkijEs
xLiXAl2yxPtrN1sTVM55NiE8M43nOoHEPu5Xe0BRrXctqXTE3qHPYIdl43h8
ZDXiKtaYJGzKbTSQ1tXlY13avwHZnGGXRA7H3oxXTqOp0wE7pcQt+CDBssJ+
zZbgL/78yv7IgxmGumk9CYzV6kfMYU9Ar5t3hla2041ARsCfSauoHMK0vwVL
hnrE7o2R61pbYLVexXCakC7hBERKn9b25ZUOHYg3E+hMbEAseeCV5eVZwjWN
az+w77qSmBCZ7Ex2uxiTOVUOfHzZZnsZCF7xzweXUhOt7vt//bY/XFdm98Xr
7/odCSyzKD/uYp8lG/FetxgPEjsBdXgF3C8w9iOGVZLEcw+oIfheSex38Fmr
OcZ+1rMviKJ/rIrFOT/oh4EhK5w1jGNCufbb0vv7pMGuzNPEJ3vUbQtaU7ul
GU3k7gtk35pYH1cRmWHqtpLbofP82bSqIz+Z2Kv2c+hI+wH4uEuEKRgBY9G7
uMhvXUiBwfOOs7loeFo4Oa+OVU1vNya8p3INZ8k90YJ6rIK+xiguZ0B84K2a
2NE6EKWSqnX64WB7A81Ymn/sBc+yZyzeV4y18C9gvOM0p3zrxaNsOSef4NDq
zsUmxeYAjPYCJ9pdNhCHA+wI5O510WQCJYPPpy0M+BRUQThWF/3Cv8Rley1K
Sn6RMMpSKkjP2WRUwtiyLmDvrk64jDJI4BF5gBeyd6AQB36hacliZyJWwlOX
1Px5UUzhfK2bB+XuwQlTyIlVJ5+s1GDjMvnmDo5JF6BgTsuYUUjONWY4TPxI
YGCU5vcqSbSg40EsjKiCDq9WH8DGqwVwnmI3rZYe/prR1d+xSpJptGz+CImZ
QoiyehY2RCYgZYk3ObYwgAAJG+JVOr3bdOn9OJyuAIugaE+uKMAt/0zNg2j6
DZc/bH0RnI/3HTKbb9KNM9NKa2DmGq/4ES3XR266+10+EhL/RIF/an9EJRVL
oPgI9pxCVnPmjJKsSwOmEx3OnftbWy/LseNbltzLEXL2pZy63eRaQb6ImhXK
mo5AXTnkeoFAaZw0oHs2oveu1UrzOz8QJOnx0rWYceqZr3W7y/VG7j6MURQ0
3ulrs6rgspCNnlR53+kNuXl+gJYFlpBSXEkQmm+U6FevFG0v8cc/hIgNXUol
atucxABl88P0AISK/1milw8endvBKzmoezhpwpszIW5dkVYjparsPyuSXgJC
0o7bEE4Ikfm+Qpu+8dEtO1caNqIvmV4Y9HEjBWR5QoUH7+diVcjwLSKbRPab
BXKx0xzgkG56gan3fG2M5WnMTXPxdbgcRKw4TGifsCvX0V5kh8Kg1tCy0xSi
q6O7DHnhZWE5IGsuQanCQe2PkPEZi0gGm0TshlWr/NaNVdlMx9rNGjBrrvrn
OmZL+vDlkyfiC2AcAnk5USue1FVO1+gsnanvW1nolf9vzY/St0C71lyNz7uL
QYI9yzbaIgtAccibgDf7KOa8nH3I3LKLDkHs0+BWJj1ldbUJO15Qi3k5fEzQ
3GiBZ/C5hs7BzWQ2/wL1LjPVlJj9+InaCywGAjhB4sLnuCYfURyLywmpsyf4
I2cqWQ3opZUotJGx90sJkhLauzMmghpLpBb27835dmkh/o/49k6p0m8wkpea
hnp/d2qdI4y7S+83dg+Cs1uWIftdbyPWWmOk0x07KjNDhH/zuVOn/CrDcq8r
59AQJ5hPpz1MSn4SjemK8/aAbKt0oEaFxSv+GMQQY1bC8MqS4gLP5/ekswrf
FGXTzKaOEeOmuLdUZ1PSHXI9ighR0umAFp3IqpBTJot9gM+NBOeIWIzZA8pE
6quNNS8Mo6YZhd3U7mwm+POJ/ERGumSq5Fa1SDUfx7wQ6nb90j3ZUT8dmFak
8U5f66irsFOxx1Z1tzZ340efu9pxub6Emgbx2aCh6tjnpTl7n/JVnXGJyGRL
PPXC/f5F1/0gEv0CC6B1Xm7ticYW3GtOeCyf8BvPMQ9R6FjLKZJKJ+cE1BIG
z3OoojYnlZiBLfQIs8uU3++3ZSmOqivqcWd2wnYKrwVuBd5sIqM7Zrq4HDlk
NqjCVkqWwLDbr5k0xBHDPPGnGI2gJzB5QIx6k6fnNXIblXbWlNIiY0uXjlRG
uHTscz4A/oXNpSVthmyCejB3tm2HV1rOoEtVq/OfE/qyatF7MQJvOPvLqDEf
WT2zvppRv1AvHKy0tnf714Gik4uFqN3Gdea7cSYW1czxgpGw3CMJ77rc0rqk
PsQ/5F+gR3oQyu8M/gnKzHqnFnLKXAsEb2RIVGAS6sDXcxJLQ+PSYIWOzw7Y
vbo53lxMsZ4h/osjHefZ1xkM6oXxqD9Hwckif82tbo3z+HnOR6CmAEMHrffm
mI35nUitd+O5KTAqeglpw9/VpMXnVh/MLmj6kBEUNuF8qicViFKRUhx9F6Tn
gmVckmN9uNN2O71uQ6XavdHPYbxwV8Gy0Iu229xbBgXjy9hUn728yM3rSMfy
fqAQP+VcDMq/L3Ae1bMHuFBDZW9zr+tPfrk+le910O0oZAXkv0KDQEJX3QKs
Ao9mRvf7y9i352wRvPuNPeDaxuHSMVdCVPBSotmSQxHcJKGF1O5j8Cc/3cym
6P7C62lvnVnEP2TYj77d03Og6tG0rAxYe046LGDZSPSFs9tWLheKVuWNVYO4
xDwOK0A22NbzDrPS2C7e0igtedU24id0clay3RZFYHgBij0meEiEMemAEz+M
DLpfUAjqFTHYyph1IgISydw13Tdtd1ofQ/OxYH16PW2jBIGyUklfKKadaBVa
/C7wcearrMSrt5dDu3r4uu2sr7t6jrifcgN6AS7Ow8G+twqEMypg6yVAtQH1
HWSyAGT/N2hnglg9+xuF0qidLhKCyWkhM5GK868mZzsp5kOJ/zE+MZA9TRh/
nW/HQVM64B6PpbXL8EqTuPW5cED28B4Hkx2NdSn/8gjO7UxG6ebaWeWK2LKa
Pn3wLb3VP4Gs5IRYoBzqEg/S29UnIunJiO1ksbiDPJCyydLJsQrOZCSh42pl
U8HjdIp50dKWdm5v++SbjsV2hS+6Koexc5OQ4L0d+gdvDQ+2HYaXjTrRoezp
ZtzzIBh2lTGdD77Wocp8WEA/TMGN98qX26NM9Dz9In7v8GnR6IQsG8WyvCNT
Ie04rzym0oVW/nNnfJaitVBg5fPnPX8SffK/5EqdbwrD+uOqgcFagUjRzkH/
UMabXBl4ki2ymgcZnkcs+t8WPx4sMuI2E/Xi4UhXRCUj/b58hKBloTlNy8wH
RNiwDgMlR01+pELoBYUJ+6yE2LbYwWr4f2ulAPmTUYlN+ij0DPWRBFz76nCC
8peyCcWoH0WgirbXD9Z4hzoPZZAg95TyVpLmhXkaTPR7NqAACHtFU+23FZmF
VCC4+pdG2G6q1CYkJy0y8NbvmUe1T3X4l9/o3HFuUSFTJwcFHl1DyUtpC/15
m6NYNsfH/2fX5HUu2k+xIbjRcig/ikk/qOGFqgK7FNJDA3yu7tIGIaEFsByK
qRbLetM12qLG/zDAjya71Bud0JhI1Ei19cEBV4YtMqdvXtHQECnL2xDQena5
tPGHp0kgOAi94noz1VeDnSrhfxKbUHFuIkc5ZwX9NrwS+hmjS6pF4HY4PoIY
FH/m+urQsc/tO27dcIXHjGvxmTjwYd1EKqrhnhnXNbNd+If2qNdfETcHcv77
hP+9i/D28d7QX1NPQ2QlK+8bIGC7UDgixb7bdLz+XYf2rlnUFr2D2uG7XH7t
iWgnyZ2uaM+bE7M5oUx9oV1H0mAoF2uwt2Wc71M9umsA+rl89GjHUUpPPjBC
/05s+Syu9f9HmASxkF9l6hB6mAVaAlMmejQ6Jvg4r+03v5tRZ3VDJfO1czWC
eIvKdv2S32cQi9S4yK9fEAMKahRN7694dmJW08OI4HK8O2qLJXvWPAvU6DU5
y7JxGWiaOjQnDZxT2fFcFwU4LrcZSo6Vfk9Z8Ho5CEcaQDtQt6z+PZ3+8sSw
0aMRzHyJEXBxD8ShvwHp6snQT8gLQa/Po+s+MN4/M0Sa787xzDINxweINemS
ysa7hHbghdQFVITZLjyNeXCSjzDw8ndM/94VC0zGohxSZoZ6McD8g9qMMOpF
K4iyJWCIACXz+cSzNf1v7vybxgSizCvcuP8yJFL80zXn76IX7aN0YA3e+pGx
pBATxsSNoumLYImDNlV95vHH0q7ATNyQIu8InPcP2G65QMh0m4SF2DxEDkO0
SD/UWAW3gZVGKktYTFBkMNSkYRpDANJsefLzABX77yLvE6hp7JCNX1eoPB+b
2kzgeoAyXmCzZc6ED7QTQlqXtBFks4OgqFuKFP8WPwKATLdu29/Ik9lpOEkK
ByWHySaXO+X5uWYimXL7p/rr60GUYQ2LYDjJNqvyi6bGr+6tc82/QXUZ8olq
RKPdrquw00yN8x0NbcqgTH4J2SJS7VL97uUDzaiHuRtQMhZ3o61vo5gVInGb
LpQxbHbL1yVwqy8HPi+FbEBG4OAaZCIAi3A9shO84cLQhkw17j5g4xQA4l5z
aiK2Bol4UX1y6dwfBvIaOqWM+99KVyRkSsx6Wjf6uCm6zYV8DC0Og2lqwhor
hToB8CVunXa1pyrfaAeyAWCfsEE/1F5dGQMl+gj6yU+t2+k6iqmOBFTz94up
o/ZPjkMR7hbC4hfIAdU7cnkCv9jxB90YKBpJdsIBYlXkuso/uz+8aSzMrZTT
ueSBCIMS0TbT57LZbyAHbRsq0cf7Tm3HSkFCTWFJPXT1A3EhEZiF+VmyDU/z
3YLCd10BXuewK4l8DHLJRmYd9S7Tqf1fNNfVjRJe2j9ra1mh0affneC5LbCy
+PBjJTk+pJDe19zWIhI/SHZjV2I+g68kp7ezbgr87pbh3GK8GHyrChXhsSHv
ImD8vBdB9nN6Lb2yCtB4S/6CpfelciGzGFWcjO79CWhIxdJeMvWr6Fo9KhIC
NhNNNlK+9qY4ZSbXt1awUqu/f9c9C8STHc8jPYz6E4HUz84ZcmMGa/t9xnOk
C7B3ukn3X8BwEQhMZu0xUmXcaz5Ew+lOjHalqA+O5sG55I5UiZHa75cxcPZv
yzTe2oXdFFLauliaIvgr5QLrVsHkTO1tipbnd9Yc35Zr6Axat5glPtxjo/5E
cKNE1Vs2MtGc5xhI2JZZbMcJ46U+xe4K+kWHKlrFKmP9it40XX1k/veNRYQJ
2IKc02COMm2h6mK6ugqzRP2EKg0udDDlSsB+EKqzeWKVradvuO+RovbJi6nE
df96jFqqjvcgEh8GC1Ve+FMbCHiClGy+US/6+iWkE9z3YMxBPhatsqhIKQbJ
7+KnLsxoyD+tRjMwyV6ld0toALezJb5CMfWNON3S/bSvmNVaXDCtRtnnIaof
RufRk3G7L9x7jkh/wXJdUoRzuDRaUIfL6WIy2uDNsIqiIPdJ+biJmz5eh0IG
P2KVyiYSY7rnUAYoNmlPm+9WMohG4VK1CA5+IW60mrxQacKZw6QL/lq0MeR5
m2zIg8xnAX/dm61jWhEV+GvnDMLnzLyOGConYdUNMPDRaZnLYb5bezkPBxLR
rhJAaUvzuwoo+Jo+JS4OhFNHnVCrPrgY+2MtF9+IrTi9hjqfx6FMCy3fEPkn
yBpF3+YIHGsa+p1gCwLJzVVDTE0tok2SYXcCV4rOrQwdOsME79dTxi6Zzwci
xvcQbwx5kWLt2FpDrChgWrIRfY8Kvia4K04mtxhXQ8jEhmMFm7lG4Ge0n169
QH9tjS80Hc1GbKdYq55PgNS+sgCTBZFTGUHaChGmnVf7+qBvnD8STOitG5m4
MO+xZGGUanvSDk7xKigjK0i0WsAyTyunzetz6Mugw6YyvbZzyvr8ll9bGzaP
4axiZYQ6J/bWD9RQrU6FAdczQdqTaqoeLbsf68x3UTGqQHpO4DIyMrfBIqcp
CYp92bSOyEVG71et0JIVCGap5qcL9+gyGMTCzj9gljzN6gvH7QL9b2OPB75c
XsgwRKQnC1aOPRT97TMl0XxLo8N1PWrqqCyb1sYO4zb2hnfbGyZps6Bx8Wkf
3qA/6C141ziUTnmeoKKKSzAvqFeon8W1bfj9+9kaO+bgHNQ12oPvnDtiPhZY
9v1igwtV7TVxzhfwOp9GjjlB0oGmnzxybjjMcA657ddJdUSOX70xVGLzVV/R
ydBpnT7uqJ+zOsFd6nalygfIGD9Rnt4ZXQodxXeamF25KXjBZyuSDewF6tvK
qZGsTFQqEImw/nnyhVRnYI+hIt+PrHGzLU7+8lW/Q8fSQqebEWjLhberhtJj
HN2VByLtB8Xsfwx024za7YugDB6vC6PiZshsNIXwTDNsToWMwCFWBZJ7VA6q
fxFFGVNFl9sW9ajiMAG4mY6FXzktagtX5Q/3APXdb9V2iwFFTAmyiDZWoOeI
BkAT/0QmHZ2GhEVheQLz9ekn+uY4MfX3q98Lk1nKoP7Ts41/09yCXicVSBEi
elqYPuLtghDOvpXiQZN/Pp8XF+3Dm1iUMiPwH4S4mdKGmn9VRtL5vBRTscj5
ImUNQBUm9J6CcM5DenEnOPg0AilWYpzrlcdFZkDAFLP51f/Z2lVUVnDm2Dmu
y8SsEHWJSkidijXpFtuSXiACl6DA6zcW2RhaMqz18esFRQetG97mwJdSCkG8
mMWN3hiqLUdcIIHMnfi4CXijgJmmJRK4i/jG7Vgd232XwIGWmw9HRsDi+bzg
RmfAzt6P47zNZnszzIphiexxVFjggMlM/a0Tk2Jv03b8cJ5Cm4eGNu/H+eu+
ewoAKLkL1AvnhG2WiSLhCWs86gDeiHsEu7vw8xbdNnOrCoGmBSHKMBnG2QG+
wXDxHPK4TaGwlUtbA+wZLxArvJ1EJtJAyD6+iId9KL4cH8I/pSJ28O1zmDHk
SMrpLirgqFQbTpFBttkEqwOgxPKRjF+C3qULFKR0PGqfOTxiHuNJGIABMIe+
4XGZk5CLNSgRcB//mv3Y/jDNKxPCJ7IH2K2Cose3BFN+EAQS9ZnxPRzEjIEh
cotwpJJG3BgfiRp3wlasXA7RddStHdLMfkaNv/sdse2MU7GiNyGH/FSYNLRV
YAVs/mD0dc/TlfjxoPgr+8AVDtkaENyIdOERVwpHrQb3nfn17MjM+ar7EWzt
YNmWVIQMLcaYgt+ozBRmuI1UythNNB5VNoTmEjp/jcsK+7J5bF3zj5JXe8HZ
H8xt6Ogu/D7ODVPs6suieQJIuboOCcwao3+t0D4BiK7BdkrjyMsQIZxjEUxW
cOzZEmbdgUN68hK0x+YT/Ad5Orxn2VG194S/PRN9db01niTsVyIIHONuLTH8
J8M6g8LgKk7IEB47NsC8dnk7sCuB10h3VS/gp8+KRBKA68G/Dw/g69TmdhMW
LEs8qyI5HIXJUI5GUGweWjX+rB88ajF+/9zsv9tGaKp5XGL+pZwpqgW6sioQ
7HJDRyVEEVpkq91DQo1Btw/WFwmdDQWMWzh247VndpfUA7NlF5+gRnsFmit5
b8h54g41alpGTE3nU+k9iKwf+YGy63BVu5GeZNQWLxMw82KUkk1UbnneN97m
ycShTO0YNdieg80D5FY+1NIiTYcQuf98Y/kgdFg/HMlORzgX0RYLYQkBpGD9
eLr1bSod1gcBOA4umZ3IisTGfZqSyLFsfVBK+hj3tiGHQ0ffjEXArUS3Pvxh
eznO30crFiuG0frkX510+fqGg+V6jvQJ3AKS2VvkuAn5PA/eWvUiWhKdRj7y
esXEh3/0Nj2a9WL6ONggaOEtMO4Zu3m4Uz+A3Y8AMh0iMSTMPLzug+vCXwqZ
uaw+7zi+lus3AEagCxyy9NBDWyhGrq8B1txWzigF1kL51W3I5qRtPkrwXlQH
gjqyixKt0eGs1MFVujRlbKTAcYMS06QT4HJX+0AZp54773M2suS8MpdHY8Ue
V7D8bWNTSg5DWUkuryc7nHCylxzUna4q3F8vriEV/a/bXEZnFySkIxnPdl7n
NHL0WK5rx+MWdb557sgPEw0H1nVl3w8gkptO1ECGKqpGpj8Tmca+PkFC8fa8
FP5xwBjb5P3Jv3CY75/VgBQNzntGKksAJ3igCQOWtJPWgaBAhkZgrIi9Db35
WBfoH/eu+tjHvxNgrtjvRb8mxpk8b+KfMJXDfeu6hpfvhtmwWfRC0RsJw4Kg
2/gc1YWr81axqvfr1zWQ4a6Jbr3urgbwwK6O1Vom8EG5fFNG4/a01X8aTTD0
4p2yHRduLrNR0xcSS+elg9jF15QAGKUxKoiMg4AYutwNpZfXsJZMQov84QNZ
3JxhYJEUtfnoJ4K4lDNAJQaXuZpN3hZHclsa7Ssdjy10BEXrghcmHXdeN6sH
ruHnVYxeZnZ7AzCLj0EK4muA7R2BDrlc5WPZ6AMkiSM5qZBVGnXLeXMaZA5U
9LMnuTbqWWnudV3E2gjBSdiLcOm5dp2KvgjtMs1HgWTQq37EGAn5vo8dXKZW
FhaslK0ijFvqyh3kfYKTJNmx/pKmzkP+qP8wWm3KMDj1RHkuXBO7r1SmzJ0Y
+9IFa7bKEStXKVdX1Adq4JYCB/npMGTYLhTtkYFCgA7e/d9sc+eLo0n1SRoR
f7CnHJ/FUkSsgzwpkXA6BqtD6XIGGYMW5wag8hPWV7uNmyVdtTrQpm//lNHH
7b1LqS1KfRBY6rRtQKzcHCJnZgg1CFkId6t4wNTavqDypF7CPR6h/XsYZzYI
zEuSbwQ5ev88R6wU+PyAll+hAiQgSX7jq1/f52zREoq62rzG3Ie453m1zm+G
EFKzU9elRD4oybx40xOAQY+nBJ1ilHvZhwxw1uxGhWl1B6929Pfnp6fMGrga
qEUj6JC9VQv/QZu9HavJShAH03Vx5fjeMBnicDax6oa/AGbCJcz66uRCZgvr
GSf4V4dXnNn+EyRefzmBeevW74YnDncvOWyw51+11XrHopKH7sjeu3On9XGd
zjqnfeACNiPyQb3tMPumGoIVE8gOGKtpJf6SEcpnksQiHFnhALhWeB7HE1Q6
Y3f1mW9sBUdgcOED9lWLwbmJyo8aD+WO/0o6oUrXALsZV31WCcp79Tno8gdq
+KlgHEwWPn1YnB1urwnFdD0/VzZ+2ESExGM8uKK9jC/kA8dJE3UifJlV+VMf
tMnilcfzSGmoCFvfgFsOfUi0w98xuXdeR2+Wd9zOqeuzIqDjiSvH420aGqfZ
bo0+GMnCDj0QtSugqENY6G4lHbcXBmdlHlJ0N8OTEtKrICJn1mKUoiWjiz5n
3WBPtBiCa8ohwbvh18xMtajkUM6VrLadNFyQW6lJhv4rIyVsQab2AxC5WRJI
iqIZA1P3sCerG14nHzEBmV5/Agqzj0sBRMgP/Ewk+m9dFE4oreYUOVqDconE
HrXcfiSYExwa9YoKdrwsiC56kR8t4Zxt6vH2tfbSDxQo8vM4sQRpKFcLYlAK
UUwQM90Pe50mu/wWDtXjB1zhD/09ffqY11q/RE2Y40wvOckzdH+7NiA7CaZ4
tji93p1bOPCZpDww75GHau5OsWkFuAkESyG/d0oTC7c9DS5bygDriDm7gm75
wK6rdRS/hSlVelTqjJ7c+SV0JTbwcD5r/5oPSpFWPs9/3BZpH4VbA8mxBRoN
o7QJrtMffcbJFkIHKsTti5Htt8wZpDnvi42Szb1RtqHwX5JpUARSEmhPAQY8
w99xBE6vpayzWwmghPUk39iOWdkbyAauz1SK6GQTQOVPj2mNuHfgtcJqiUqP
iVpYT/3yGWfPNDVTIhJkW9rpHJEWZ/jKxobl+dPNkbR60HCCzkxCdcT4jZX4
wGiI6GnXN4QGDMqk+3+TllxM/9TZEp+n4wxgKAykW3z+Em+PKC16mnM5PDad
jgzdexNvlPWBkOZw/9EGW9SRSoecD96B1yUemDBbgYg+ARt1RGD/EzikX73h
qQ9SiSuf/mpW/fEZIrKKgZ/LpWJy5cQl9a/Eas0Uy38DWGfRyhatIblWJUWg
SKstTUTtialom1EAeNxyTGUPceUODTTxt9HsnAVNvQhjQ/QtTTGIZvppJCcY
BZ4z3H68O1ys4dD+fXWRxTjl/vh0czGP2LcXBaRCKcc0J0/uPH/AAHnJ52Em
PBieOPRlQzIrNgMNMjFIW8ua459zGzPjoNMkzF4kSwQDK3jMlnRzd4/Kcxzc
VcrRFCcB/MlBR/wwTOe6TSZ2v1occhaIFY4kOaOsTMd8jJ+/686Vd8n95yTF
JED4aEpJWC2eqyzuqTDjtXqLlRsxkXF/f/U4UpgePSYRppN2Injt8hPYZ5/C
ozIKlGzCO+156UlnYfOqniZr0iVJPUnB6cBOUFArmIWfnHLXI0OpoehQoMNq
A4doav7jpk87M3mFxy8T5J8EydrSwUlZfe4wwgWSlyCuE9ZYPUgCVGCusrC2
NZGam+leqqgpGXSFkVEGIilkpK65GjcgAuh8qLMXHq5wmpMwobq9lTwFk0jb
AbNvHsFWLUdsQMwB+8TIiGnWP+hn6mi4WLcamLV7Rpj4OSvAltuLoa6MbcsT
JDJrPg5hEhwPNglHjKUz/JxUKpqQjWB67zYRL6BoUZ3WsIIl4SyseipLyKE0
sN9YD9OtgfOWbSVc9alwUjXMLRtQh1yO3L+wJWWyBb14zpCId7q2fQqRf+xt
0m2r0mx8N0/ts++vzqDruiGtWcA8ERPU+lByGG56F/TTC+7wkkFdSJl600vh
GZyJWncKwrK8xzXQzaEfDeS3bzaTAjLvlA2i3goAQexPsj3kF1y/nZnAtLhT
QzZJZdonIPvWl5lyIPsI0wt0r92z9yJD++mk0ceRTDqswp/cumcMslP/44SN
PGY7Fp78MpFMq7qv5IyFJnokAeZxTlU8nzP0ju8eR07Jt5oNVUjqok51oYY+
7NZArt3CoS02v4rUQhw3wUmm5mTRNZzY52tv9cho3+SfTp/U1gBt2Fby6SaB
IkXTN5Vcv50XtPmj7KfqkZe4u5nvNqrEwG8NL5wsnOioVHrCid7wuE2AtZ03
Zt/ivvWhKwCwFKa9r1iuAkZmmOubWz8jXGXcShhQabosHHXJoLB9KVerS0zb
BpcYj4x/2qwezqKGT6jA17n+Mtyzd8RqSyQ8dVJJAMOV1tSV2gye2USyIiw2
G0QlTXAmj/o+84bXgqzqfkzIpduNS/Z8F47NlXce8veiA0qrGTpZgcGjNZiA
p2BVrWwZO7OsGENnshc0w36m4ofdDrqwZU2dcLaOVKwDSrYekIF92J1bnvHy
GsG/8/jUZyp6tqrUWRu7m1RmfD9y+PD1DTGBDEjQgoZjiedziqs/kpMRsYYV
dxfw3bDIIu3eB2UolfulEHNkN4BO9hXUFbPeL3aoOqSYrHvYh7EJ90tvcQ2R
AGV8q846iuft09QnidO26qw0tqszPQJvcdRAozA5GTIya1XvNn5H9QypgN4+
n9Sb1rUCT6xohtL8nwr/zRh2JpSP40ofGDlkiHBkblOWx+37tfk7+G075Hm5
vdDl7d4oCs+nisKTDq2sd5kcVoIUrlKmIdwWt11+f7LkdsmOFRJf+6gTe3+O
VyLbVzZ7IEOKfKNCokBBwU6HrUmifKDnXuYyAcpi9etHZOTi3iUq0cKXudUc
a4GvlK7Ge8XS3wP44zDyH+qgAGQLCKkSgBDvvVZwQ4cdIIX27iepJxGW3sRY
1mHhFZwABzBwM2YruVAZohDZpQPdhaeGVfsQ0dLaOgFrrC37rRzZLmX1qV+1
bFvmg+1sHHWosY2WMMTosedPAD6IlQNF6e2FIzWrlG/dTZUYlpVJRdWjcDQm
75DphhwGtPdwWRx0X8QuIoHTmKJfigx/G99pNV+r4Bpoy14KWizXePYlnJ01
jmSq8q153gij9H24K9+oMlovOCnbV7PpOvCozC8emVbkgcbXzS0evgabChtU
nDryvYci/1r4fHQosH3gIf+h6fDZip/TeEqhXNSvFi9tXcp10NR/HPNMlua/
AEz0QzlAOJPmr76E17UwJQALssjvgLcp5sj+3LwQx1EvSifzniRTP2X7F3PH
mUUvYz4fzp3Jj7Svlo+Bvtp8uo++lMzvaBqChlnZzk1YiOSr5VukivJzPA5w
BThx2L/z8Dvth0KsS4Sv38I/2X8+p6DKE8A72txf7BOf2nidTlI3sgoKEftH
6LSqeCmItdo1HciwR5TGIIEe0jmrGEMUYx7hPwgNgWFiBpgX/vYCxVlSKpUa
7OH/USEudfKmwoonGYs9s+HJcetYYcyPtjgqIR9Xns3G4r83NHFX3yJVmp3t
UMjX1rdTAGewp5Gh9v9skaXBUuR1o3dao1LZfynRxszlub0dudzC8TJsPSoE
ahZGSwQPwhJIzWWkSTy7xsRq809d94K7CXpL/ySpoRRoen4GOFDzlS4P18Mj
Z1XSwpDHN454IWcx8HYxcSnfoAtSPDex+hb2ekyDI0WTvO+rBVbK8JvNHx+A
WmkoCdJTlrVtBxzA4f+uiBuU45iCJoz7Ly8h4nImMWhXgdh+CgU/UiwC8zpY
G/edRw32wpsZ6NeMPh+LiaXWWzai3EsG9yHQMHB7bcHpJefDcNjtuHAz2Vlw
okylQ+10MbTJXT94LibqVoUhQg7iYE8WSq+m3cK3CijVAA4jDt+LT2wGGVIF
SnJnnQrZFq6LXAwfQMAoRgCWgNYva0dP6kDJRzrcOE8rR9BtEN9fwKxKEyjE
nrcHTIdIxhUTzAa4Cf8Po2gWGiBEK2cP35ZZzRZb9Q0Y1OvDAdorZvKBvUeo
v0hsETMmpLK3tH6KHLsQtAtqpwyGjmeEMufBACy0t2okyfG3fw3PmgUETShi
wKw5ZDkZmUc27vXUAo+xZFX9bqJY9DTFS+UM9rxaXjUjYnEzelLpBwwwLa+F
6b3s+b65XuMcEYqa8CVdT7/5Beg4Fa6ZKGrDo6Mtvnpc+fJqhpJZNZdf6gAC
QdFsaeSkoCEVYsEHlfy+VBEG43wSOaVouIcaq/AzJg/YstQO8UZwLPpRbZXb
QaS1tj/FZH556kBkVZ+Pb4PFqvjhhlsCjD2g83sI8dIaohHqfjfGNN52KbCu
SR83vMUe4LW3fQgd80FTdbXUFDILyzUmxETY8j1NmFeZLMWSwX/mac6Mhrx+
1ngYG+yiDfrXv80ubmmhYaayVhuS+dNZpUZyMTKeDd5amM9lE50QZvk09gx4
lzRAzaEtq1VJgObZXBQg8bOLSWrubd+4swXb3PzG+sjC8IHqOi9bdl9uKVVH
7Zs2IILYfIkVP8gBpT+78/Om0NdT03ktcGztNPGLzxnf3nm9VoYonUxYvljL
9Fp3njIpZEk/nEvYbQi7ly0cEENFnpMomHH26HVP6sYnyiY12GG+iFSKGiMB
OqsWwkAkMP/3hcfNno83arkQj4sSWJtHd+lgr099nHd6E7AETphZIZHoLE2d
4Zm2XEzLBe6FOS4xkK7dMj1gu47ae+Z7itkbJdplVo5YRwOrjzhZ/xpG4bWc
vOZDA52z4P9WtxdzxF9yiMbdfhxBoPZMnGy5762fb9Ttgu5RWruey+8i/uZf
x2Zrl0K/z1cWUy7Rnc7YedpCvJ481oem9ygbJvA5kYNkN1RutRcaQR3FdfE4
NnbCUWeSJcKiNiOxZrgsMUcpjAaWYd63MxNMZGhgyyX9nTIcBHRJ4op47CsW
bM0WMpcZFETiqW6ul5Fd/kt8uN8/DPIFs1X1jSggDUqFIMkgFq3GTmlaXW+G
ImgifYZL/kzYqyHxDIw6tJAcq5f01Q6WzFpGByjlrAQBmbgMI4wJI3w/z0oy
gpByVq/4uwPXN7sD2Bwg1+DoCXCN41M7wNrixWDZGVlv2kVu/tx3dezvZHpX
0GETC6Y2rkm1WdMOn5fVBzCzISsU8zmQTKfifVRC+XigrYnJ8KF15wBizZyp
Pjg2iqbfkTolDsRynu3NJPek28RGcoYSLpRY+ott+BKJdvne77sWJIrubkeh
39efb0ALXOab/HlbeKq6yIH7jcjE/+qPo4wFNIfZSA0AukjAplHwxPKMSEsN
QbS6hQMWBVg5oLI3t2qmPXGNRzyM0CgyPI53s3yyy14QR4FO0wOHIWowurAT
mpki9pxMnZ/4a1n4+AunrZXyeoKFwuuW8f49XHEfn+9H+4ZhpK4AucOahz/h
9qlMdaEr9dudPtsm0gqpCAo2CgggdoEQMPJ+2td/BXSO4sx5twtM8Xv0Mt9W
bnhJPd0iwbues6d0C4QKzqiaXpEKPv2C8zCccJMj//ryZRRxzym3DDWed8qg
M857p0XHKAyp6JzXnWD8QoDLLEnLih4srKi8LY95tw4gCjZ5oCqTtSexDAkp
eg89yhlQXoQrTU/BKOu9GSst9FYPM0r7yaHMFj4N1+f0tknTJ8VQMU35/IFo
QrI6MS4VhNU8vWmyVFqtkCow1xZ49wXcU1ukyRTNXKUSZQ4sm1vC84XYZhra
odxjRMqKztpi7M7sKMe1wVyYy/WmaJPkXt5d/GHBNLcDJ8S8rPkgsLE1pxnt
biabYXMoYZK61btVU7xuHSFczQUyNACFh9wdQQVmxdkl21Lw+83QTl0pLV9G
ioX5bLoWO98JVMr56OGcDqwY/4h1+6rP6wUQwt7mbi3ffgBkYCcQOLD2cc6m
5ej61cpfaa+IX83/27fStvgGVFnaAPd4q067G3R9NPBaR2k8UsaY54I6aisT
fjdPdNRyyvSrAfpp2Z8IMvlBzmRAj2St/KYcMjq3PaRSm9hQEfJLvLbHkh2W
Efl1JQyRy2L1OiZS2M3zg8rvQh8GQJgxwy1nUO1Tab2j1PuZhzJ5ds6ZPCdY
RQgiG7tBOMC2s6e6y1SI88b/QJBBdRC82K7Eq58AlZSbBogEJ15REGkcyXRG
6dFKpRceuuZPX7uMJWVh8hnLGNri+3uDg2Mp/C8qn++/zOGXw1owjj2VYOh+
yi56DKBusWgzhLd/8vPPSBlM3LMQlgw0ygsNaDGvs6oGTJyd6TY3avI4i1Mh
TN/0vLX/uPT4BL68lLpsfcSCEP10WabIzB40wosV8h1ZZaGTTgNjbghSZ7ug
gDz2e6oTggIUFRkQg7RQK9ktxmuEPe3W4w1Cxt+G5qBrRwtIkkUO4MkUKKDl
/+BtmvN2r8sbLDN2hSV1lMAAOnOS9rwsdxuN5v0pw6/fh+RYScn/FjAyvG7M
IjxZoFl2fGnOt0aMbzf3HiTGqQix94XyF5V9A4uOhIxX9zAdc3Scn1aJQ/h8
5cvLvXDzg+6FBmU9N5xCMNgZnKGEYgmSlt60NohTkk8xv8aR7HFP2llMQgWM
IUrZI0wHb8spt/CrJ7+Qpnm/Dn8Gu38X5svkMIL2eKB8goqh0TOoXqDF2dLj
wJIEOZVlxNyepdBBElYe6sPTNwJ9PN7Ie1xUeHLCnqZIlEJJ7b+qdcxAmWnW
+2M4aEqU7iS4y3cJNQ2/Q3tXlcwxV8dkOcFyri0NHrnBR++sMXj1nbhy6yCu
WF1WZ9drjqzGeAaEGrjLkerY9MDXO8RUlbesV1RMFwSF894LrP9I5w3+OryI
WTSGyXW+rpavAaqdVorfwGWnqctbT4rGBqK61nbTB8kUvEFOEMTB1Owv7nOG
jf+hJ2+iFVEKXn5ISv6mqXIbEg9SVPVUZ2IO+uS04fT2y8zWr+95+KGokqwU
vlEXQmSiOEmkeYBgmNCUkfX5dJEWt4f6FVPR78cJZRMsl4og64c6daPzWxJF
grZhcn/d7pxebrSTcdmA5vEiCW5AyPfhgOaKefYZhGbYehmcR7ANF4QCZWZm
seH9wCa8rVI/5OGdvj9jZJ0Q3B1snRgkLS1nyz8/wWUid1KdvYw5V1x0dS3r
xD/65DJqIiLDZO90akD9HoU3G0bi/JE8ykdhCDV4oZN+E4zfX4e49VeL1QKN
eU/Pa+H/bZamX0zl6pS68h8fYYNbc9XXyxnnnL7gnRC8g+L/2qaazEw8cm6p
YHHNbcmLsEjblEvTj9ozyKMbKZkU73mZF4lSFeE+M1vJqON4NJpJf0A6LIOT
EBUflCRpMMExDpDGjlybpp7mILEWoEeUaU19KZXuQyJXH9F9DGeLMlH6g867
vi5aISLRp9yHU/g888c5Wd9+2W4h3r/vTo7ZM1uKvO7N9uVM0GSf/L88hwU2
3900dwDiotbTENdz3DC14FfwU5mQVFdPhgxfnk5n3ik5xT5AqOlmsBnaau41
h9JPFKS6ujsljLSDYr/t5R/gtX2rbRa4ElR82AK12OpP0iqBUUi5MGWfBhVX
/CLKt6SYGt5XbX5QDGpC9JTerQrJ9LsgJEakHJgAzXQnfdO/5bSEbI9xV1Mf
ukMF8iGysmioZNAuPmHQACUA5DF5jdDVeUgZKyAoytVOquQlocNQpsCkLEfV
RiSlK24G62BLUBnbwA4i52uemsOib+G6COZgh1nekoiF87uQlOYFguit2wcQ
HK5ercXZ2jJa0l7lQUrnS6EcNVlaUb9EuWW7rqSnOpHjJQw7iqCREYcVawjX
Ggsy2W55V/WF63Ffw/phY83YVQUPKUhA9E5ozfLb6aux7X0kNTAiuSDBGYw1
AoDGVQbd3K8SQbqTFZY6nBz2/loxXmPsNkTM7J5KK1ZudwKp66DuXVpeZZ8Q
9dTasUby5garjsqPDbWSMGBrtFkm6mz8JxDnZvOBsKM0HcwnsSxr4OaQ7JCc
Zry5VaWDOsEEfBZYn9giXCWrocDvR1kNJ/aNdrVA74xlOhX2Vy2dBJP0GL9V
WIl4uKuWQk3DP9rNdyZD95DmPq94KJilFIJ+QEF8X9lb0vgTOnG2KnEbKL4J
J+/i2iq3FeCZra96s77vkVFN7Fwh27YhIXypf8m0CiBU++R6umbmbkqwZquQ
5Deg2rXqLvYiHlJiVUsglwPTl5CwWUsqpalTIk8Ze4/VVpnCYDf2SpivNyP0
X7Oajqmke/Ly/vpReExiOIgyGUt4bSWBeXp6YpActwbBZjXguwfpz1BILQcQ
KRfY9DgdgialaGAaKHS2cY8Dj1hL7pEk2qajHBIla2iZtHH87D8XXK3ybnR3
gtiXdABCknkRPgwS8dmltqaPGvKLKHqlfeFTWlSAGf+V2F/JX8pcMkSzjhmm
8IqUT8xTwzXuUBLpWsXADro9N/m9DT1TXi0N3iunhdklv60YM/vUq5/A2npE
nB9fis3Fv4b/Ztbu1H8vauvKOz3n1mPOSHrTbUhz0VPOadxqq+cib2vg1e6h
W9hr7qPPze70xR96WUSUq+x32SBK0CLgH0jwls126LbwiOsfhAY+4MU0KZeh
9oHXPqTr+ovh2OnMn8ZiK3b9IbQy/X9MQub+UqLHjNh+ED/O+ntOuFaNhQbI
223s1CsBxDLlEYLBU1f3Uz1gIvbCbrpIuMJ7WxxtFA/EQpGrrlZGfT/BUFOL
L4WwcScZNPhrs9qc101pVeZXgCiHOFFE3XMxpupqhGpkGVEAYIlyfGnek8Gs
8IYgQ+0cY3H7rweEIO5pTvZH5hoap39LM1BzHgzEjFHLcLve5H8JIbpvwg1g
+Qnftds1tfylavq41+Qhg1HPIQg0ompTmSCD+2Oy3j4F7v+YiNbR3HTMlm2L
T6PuF8uP1LR4dJ1UIOpn2p93+Wu8KWBZnN+Qgw03S+5kZjc8O7F6HqYEpszP
r4PX51R8dU+M0viRx0yYKEIW7lhFg4Ew3vfH6YKGB08xGvCkv1rcuDZDZQIb
cwnBKgBA86AA/nhHySGPHj2dL45QC6irXGAh8u0osLMZlCBb9A47HeNhpaMI
mPg8ZgYajfma0HkgsEsEqqJ71TMayW+rJEmW+G9ufxYiEUH0X5r9d5fjuMqE
Xoyv9R/CTBMy18+z+bmNRL6rOR8mHksfWfeFVH/BaL97iNp6prCeI/bAW6cV
btTsRc0K45fJpnVkMs/GS+lRZ0mOCvZcTIGdbpXZcwOg/dLDi9vd7unAo/RX
ScUE/a9TeHfzQHvTwC8TAmgpAgLrmYwDUlfgvIvVFzJVtKLvtCV+KRq2x8KI
tj3VYy/Qk7Mv9/YwelhATmb5cT/DguikCNzu/RtAz5yTYCXSvzgGq0ZEtgzK
9FA7vv30C8+y/zISmtS/GMt9cZ/K4kp6UtkN7xfEPjgBB1S4Dw6J20N2RTW7
jgr7SIoDu7VlkWImm2BjODuopwqmsH04ED+wYljfjaksZ66JMMprHDsXtqR8
Q0wCk9W+TCfNb8eBpnIs64t9hDx9RrZYXQina0oBiOwJtm0dM5BRd/oaX1L7
tUR1PxMgdu7uxudGJiQH8ucKA4zoDVOc9diKuH87KIMcDmtwd06n4dJ6HxDF
L0tAz4pouuMjfhH2DjEHJkAOex9IAWPbHQs08ueHzoOzvT5M9OJ9H05FY4Cd
yrVhwyNyJTUmfnmjVMefeqlXnStGahjqMg6f5Ja8HyCYToCSTm2jQt+M3xC+
8Yx3cdK3i5C4lbC/PorJJcWqgj2tONGU+oJGaaGVz8YLeLKDOdE3I19qRgde
VKhwfLkknZYX4GOZrgKsPkUJIRdrYEKTynkGtxZSDXDBvavY9AYsFU87fu+z
kXWlskwCXbdsFVaVTd2aJhLAwqPb9ZYdRJAL1SlUtnZ+Hfz1XuunxtgvKzlt
dHSE5wpKeP/teJMgLHEysu3rvMEElPQMKHUg/4+e/dCV7tSXXTwT7Poxg7GZ
YVw0TdjcS215rjPzjudFWgTv12aD/PIwjfN/6NKg6F03bFsUuxTekxMCLj8y
PjNdf1xth6MtZkiPtHuQCS9OURx67wwKOi1sObE532kHay8h6MwohHBhCZ7R
5BALDDJM6GQR9nkw/0kKkRcfTJHDL1Ef42XlOPXx74TnyWqVn26eTfC+/VwL
OtN9Z2inIWlhC0wpjIz3sGSVu3jb1dqaWbrMIy0sce8HfTtmr5yfDrN4eHgc
ogo6yEMxkJd1jko2JZCup3dPBNp3Dxy/C7JBEcPeKgFki4QsuQOwLrVM33LL
IxfTeD6Fu+Gbk/fPWEl2LZj7ddr1kl26uwt1/BY1aBJd4owntjQ5vitpWE0I
Ev3J2+6TO2QGwsOniOWDR868gtk9+vibgxEcs5wa9RGdeLGs9R9fVLo2yPAY
RC/QwQIaKvQWh3cvefBqsK69IS6K58y0CtDKr8zcJL2qoFYvvpzFa8WIaPoC
VKf8hsTsqPqoXwHCFzLC+Phwrm+3RcG++XBDjzAgbRfHHsE6iugc5T/HTE5k
P5cmg9zSbG/byiTIt+VJWctqn1KJ9IYhkMhFip++ihplSkHSwLHri/N5xR+5
24AwUicsFxxvEGxFxYOS9ih8H2IpaVyAoy0EmvPbrOJKkHiyir+M5I8fXSfu
F/mvrjdlHf9CQQB4sznqZf/pDhvXItscq3KOxjP5UrqSFrMnhWTy8ZjNTlfw
M6yR2XIG6qSEYeU0DFp31ThtJK+WGqR2JBDodF2Ra4IBxepnm9dImQN0Br/I
/sJewQPbmhAMb4FHHEkxkYr9SJeXq9XZdAF/yp2TV6n8CkEB2iP0xyhDZxzm
XiUh3JZxsS0Aw7s+l+qvIp6iS9pNUACOjEAe+nG5T5HKriy+TrbrNaR/h0Gs
OjUxlYQ4cN39rozbZBqp+ZAFpzSkH4XwYWZFtMri1Ig2u/y5geANUe3spWXM
EblWdMyXQyLLOtpggcShvE6WavZD9TRc835IioZKs0DKX8ryuIH1C3nN3hhH
VIq1lGhOJpJhvih9kbmpgJ/U6zKmBIH7kXbUCMtJ+jDFL+RkXQfJ+vcagAZ2
tGwuQc/pdn9MSKxFRRd6gDaurzL7CczAyZ6Ao/n+WhpVm2PKcTB/IQ+rgss4
XM2OncKdxldqTtA7V10K0Vf8q8kHxvRJ2XJUG6Reg5g7tq8TBgt6kg/QAYJ9
5qHHVFALjr9s76Y2369LQrjlLr7sqPRlBAMUQLooIvTxQsB8qbz9h6z5N2t4
9XgA10g86ih5H5FEBuldzTsbJ3hQ7ajyw7BvdA4WJcw9pMyNA2TUubDdnz9J
zrJsiucDvQHtfoEFt0C0ZIhuMivFw9fYZVyz4t+LLAgNoyy/oeMzbsPNVEwo
XtZYmYfxHxHPubU7YNbvn9BVv4ZW+3JNTtAaExYsPbH/o9aUfAKMy/AF4sfI
KL5m/ERQNew/nHmrs+JdB9vyGpvG1d3xyODSqMG9uy0fam57zBimUVCISwkS
OJyOOF+VwfpMiW7ms9a7kSM1RBBDNXEl76Xma8xVM7ubIzpusnkniIAMrPAl
lMcPCTYnfBFOpMwz6ZYht9qC5TQYoHv/XO3ZkCw97wUYBSyH0+ZKTtAUpEZu
Ocv9/vdlrOmK97yP2kymhvqDgFyb8acRKQnOcoAtNXvY1oKcvZs3roA705YZ
qSAme8kwzVrCobS9QDTdJwslDXbSJ6V5CAw/m17JPAUx1KXBp8uie5jYT03i
ThdrAvza8jVNPgyM1eCvMjiglzyPZQ8xA2Yylpr5tcIUuF+ris60oQhKu5KG
+UZ13H0o9m1MgOZdC7DAaV6k2nJpjJVAScRjULsAYqY6OtWW7ipBHqdwYJua
HJSJAAMov0wffh4MHICkgznkw0CTy1gU8SThXHj94x2vI68sT/bTQmEIIs00
ryIe5EZUNyFcuscDGU197s2oLizWi/D7y7BQCKA8awW21epvxosQfJFsTe9R
8yswB1rKq1ieTXDat5b4bvIwlfNit51ynt4HVNv2SX0a7xCsMKriUSDhmSE8
HkmS8R7JElsKII8f6EM8JKKkRxwy7q/hHhKA36cfsXvUox7mTNEFsk1wP5+F
WjQnehSlotEL1X9vkhEMS3wmZVhH3fYjhvzguuv9A5yCQIGDgPCWbj3hfe1P
k8690qje94bq8FvKnzC2xkGyPYPS01D4AwJ9H5KNBJ0pzmIyENgnmHwcThKd
iucEzVVAgBwnnHKXSStfxWX+Piz0jnCTbsh4uZDi3tsm3d0KUGQc484ektpz
yaXEx8haNWPfbGprnPvTEqkpvUnRQh3rwMbutE68e2258gInQY7hinsC+Gxx
7MIoieuTtU5ymRHbBsIjB6rtT/Ql5SFFAGyBVVNmOgbQiRKA5uNhRwBprnD0
i4pJVI+wfzM18yH2tf+iM/7Mo4egXfdeAiuc/f0Ejy4uOGK8LE1tisKJrBdo
WqeV8+Q8gQwvjCxxLsmOTRm7vTJcGCg9fGZtJJyv19eoiVrAmyfIpNa6/8PJ
8N/MRaNA/B7qc7pZnxaWjgJbCXa++vdtijrih4ShSMcn+CZvG3uwpgOa/JYY
0pPf2nRDDN9aJ6u1UrrL1pQKea2C4mxtzfimUszfc4+reXQXRHnj13HxZqBU
FVmkgg2XifFGx7nvxOet/ckRiXgK70j7rtjw27vlFCtYH6lBGD1ZSpTue980
1BUdv3C+9x/531Hb9KeX5SfL86SMlyhvYNeo7ZidhrEz0NLlytNDKY+ODtpP
2NVuyL6LCDpy9lbqak96v1lPkhJ5bwAcHzINU8cQUGyPISt1Gxgvf/46yvoy
DS67tDSjn1XfkpUSWQjyUExrv5+5uwXcwVb3076h/TrL7+qdpM1nGeh/l6LZ
4YBV/PjzeTUWSLjUEir6R37BrqH0O2S/xd78fnj6AgJCrZMIgRH/WQBORRgx
abKXVxuBnpePmwZxvuAnXUY5eapWNdyoqdFLEtN6u3yxQqO7yFouLvKWXTcP
rlJwioq5pEL7iURogAF609xxPLkaXLPVksZxrX2uf1LprfOSM4CyBD5ucgLh
DlNtdyBataR5bIZ2PItBrcAJlKgaXnOLee7ZBDz18bTHHQa9uhKRWeLT4v2x
R+B+Gs0f2axQsO3xSHW5OuJ2Lo9g3iRKtfXNP89kk7zth1UmhYjwTM2r0rFb
4KhUyXd4X1NMt1vP5kNEbUCtAifB2UgUOS6BEkAoy9vkmq+wrjklupoa22vk
Gy/1HttwGKvY00ZEhikow1s/K8PyJHTHLVFG9GlxR74q9reAT2Ei9ZVm+J6q
BTLb5eJZWcngtq57KZmf+HW7zxgVCqNSJScBUzefp5Uwm7o4A5TZP43fqX/r
HmWrYXYtVMLsXCjO8F7zfw+divuifNEM6LMWS/Q1ZOG4dgdd0OVA63bsbEVF
2Vzw7pfECrqfgZT1OSh/CtWhKTQe4R8xHDb6Xfl/Xt0rNlLpP+JYl+/Gfd6g
ct+rljyUO3gmMwpCpYyD7CGk+IU87uTBvRAeKB6u2mwID124heHQRNgAodNI
0JTJvnDKFQVWMu9IkJUyrLHAlrhlkGESaEYgViwS8qddro9AfAvKEgMhh7ib
fRGY50+pU6xxe17folUNFrAN4+5yT3umHpm5Spd+9r5cK2pS+gaHxSeS/f2B
+sZ3MD4DSzEiqyobX5rtgJ00fRIBynj7EaeDVLmCjWAq2D1OHhGRZrhFhN5i
yQB7XuItokKmi9fiNvoavck0pZ8gfc71S4q74KLKxG8pVGUc5vp/fdHtz2/p
KITqV6aXLPdPqEh2znl3AqrJQ6Q1SmE5cc+LQA5fMyhuzVcdQc8J0WUfMUk0
Ti3rM5NWIyrj8gzXjxfG8KRecen4UdhT0BASk0YUSDWaAbJF/B4j5qRWozDL
geo/1h3nlG+cX4qWhWKSpnwbFPkp5LMwlipeXtv/fr1wVC0qMUWxo5o0KGhR
x8s6r/hWKyTI+LzvPmkpq79ypdgru+q/W+9s63C1iZ9w0ArA5fG0481oDvcX
0teKXkShaXZWo0DR+bk3cwv04IOE5ikZd/UVdJGM9R3CYagBr8iMwDOXDwi5
i4Ho9k5U7CUdUAi+ZzzMTzL5jpvoHjhag6LPzdK8/D2aCN/0S7ijlQL6VtlT
2aODcYE1zlcauuUUc+DeGOfUZ0btm2ZWs1QTZMO1bDdspH40LV5YFIShoYwq
/jAqBGY8o3SUJgVQskde/r/WSQDqq9920SiVTINVgdM3yejfUYSLXGnOP4j0
w93OEQSYFYFd9Nc7vj1oy3jiAjjPAzVoAWFaSUnHG6HgNUnjL9jkYSfRx9yV
GcJywDJY1ATaL4rCHWBhNjcqWhz3czA0KC+PKWbCiReew0WmG374yfwKqTos
iphP1/OADM1fjUSOZyulRD1G6WCfV4Cxkx3BEpwWnqRiNe/E689S+9Q+G0pu
fz9xsxXpHkc8khXxfFigk7Gu8swDwQnyu3frM1g/L9XbzglS3k2QK7S1samz
okAFRXeB5RKx4SCocDU0G2TuLt2sgoxRYCpObBloP9WuanU9un0udJpspzmP
zvU/7ef4yEiAA+y1RU1V7j8nX2N6wlYyp0jtcEGRJatioO616gMmgi2kDdGT
u9+CHUejDWtqDcpX3rxuQYz0gHfowpENYKZN/PEBolgZrB/s62ggZSKFbA3O
XmW7EmGT2X1wPEmi/5l+2SUgOZ7uReDJDH1yBeJ/pkVvS1G+JIZOECs1cLEt
IAn3AZVlG1UaYuH8ZvtjA4Av5R9OjNppKFIFzWrVazDzrk0XO+yb99vFIcOw
FF8Cb6VdzP8Zjqb3b+Sx0I8FPyFkb3KGM+TR9sabiKgZtv+1FPQPkAh0vzUq
zISUPEksTE/geMKHn4ufGwnUHNG2Dw7evT/oGwRHxxLJKXepv8KiQsCR6Gm6
c7wYT6LSMfadaakXT6usRcDr4bLJpVUxTS8pkt6HERrhiDwqKaMHPFi04lxt
WbI45STStQpUHyMpYV+sWRpa2B822tfWKQLtD5kU/d8P2P/kxTVPUipvFOkR
d6+k9etpVYVhKrMgNgoCAt8r5Yh9udARp7eJhI+CwM9wgvMrMEVSOmwRoqO0
GebLeZZFnbCFocMHUHgg7uykB8KhCzQgMivArn1kuatMKmIa/kD6PDJ2NBpL
oiLWBOZ4l5vjzVLgyaDJp/IEKo5zTBc24rHqFWzAGRdf2WocRjbosdK/UYXf
YIKoZ7Q7Mty9kZ9Gtd+xaimBXZllqWkXiZy208UIyKaTGSQF6uPa4k7yHNyg
7YVwKKvfHD5L0mc6ROZpO752PyoX1MsucyJhGzEgbpk72C7cWSvHaUjlJpRm
i6xNsoYDkiRqNP4FX8fdmM/3EASdF5seWOUQk7aGRpSyKwBpqgkrTQOCtucB
oSG9MJImuZr2ODgak+G5k4mWG4ChwvXFxEs420FBKWiX1Nhc3jqmHCEM+QYm
sA6nI/utWkEwgJepwOPP/VZNAXj/hh2lAylcYsuK1IXp7Xl8SHh+3tk3/9dd
u7e84AgSTyqZ+rbyKkUOvWn3qqBfn6sz8OABdu1ltYbMkMGQAiPctzqR2oMf
Z9HOhXTJQ1G/fBXSqriLh7t4viKdfjdCmyf2glAHSQeVisLZ4KuZqRdzHJTF
fH6ckXNNMXn6fk7I6z/I98HlFLXLXH6INHVmVBYH78a28gFVONw0hHBvL2vf
7gwqK3lDYIH9d/UDVHPYQxlKUSWCliokd3dcbfvVD4JzeGMTJugbI0J/mEW4
EJJYT3WJ6kOoPuaCjDpaggMHjWGrNa/OuK5u9Z0MytC7bXKdDyfenCF57gtW
Wx1gzz0M6ya/7Ct9b/7PmVft205dIx+C7jBamW3GcHDnDIe463ARl+tIcRcV
3a/L+k9kGLtMlmFKsmvPiRqyRSzdvjBpX5Yssdnme3qdfV5MOW7piBTl+0+B
fH+DwZir2YaYtmuatERk9xfN+DgBqjVbvr602xNpOHWVtN/4OjkJYWwyj2Sw
oWNvF732rTTC1t2S2TwltVGmVN3TdEVnP7gCtekw+4aAXL+z/YUBKq2wBWa4
dHsIygm48WHuQ5JoOaqP8PBL+5Wcei9zQdZd31dzp07loIn8IVd7mMovPK7V
aqiUHRf3Qdsu607oFqja8J/PANRQiyZl0MEgp4aPsPs11e8DgG9WOAO6WjXu
54WbgezYhiad5L3fr1khhX1QbH5n1Y9KmLes8QUU32hu/w9PrCkwmzvYDSMf
OKzcvADJfnar8ZqtBwhkH9j8uhZ9UwYWbwA3BGgVpTO2tcp175teCA5zvUge
DPpchzLHf99iB2le5IvRLGT0iQXEa9bp++PrxQa077iODdUfGpJ5BZVAW/8h
C977ssDueGtJYm7rCNNOTdZX919iMMkgqSGvSKdHoRofC9p945g56UJsf8Ln
Ckj1jKlS6sURpD46zIrv4lT/UnP5v3kDRt/7xxWE5K5BGipF26NSmGoWsqIt
M7yZBmAj9gPHA2JvbNMgZNgiW1wIWr4Z3rcEraU32+kV1zERLmuvWFUJ0LhU
RsLZ3TC5lpYhms/AImXdE810/ZvMUJE4R5eW2TPjTe3s4RGO3EcwOm4pQEsP
6wWUJGw181OLDw5iOjtJR2sLAuSopV3vqqz4dKr5ATj4FNuQJSRjo35G9VaY
9jQ5tVFHr0oCu6iR2c9S6lMwbGwbsBNXyWahV6Rz3nv7yalToQMB8FNK0jLm
/afJQRnKsxQqoMNpDFPm/97Wye7S/9FfW6bZKBxnFfasTWfOpIC+pwqFt9fY
+ROnxiYWSBvWOJlZFxpc8EVa369SuLvYcO0Tv91D7+429gDPnuIPeTqS0TDn
UIA92WnyTLuKJWSonE07Qe0eqxx9VoeUoI4hVrgejZkJfBr1sdlsaADGh7Ae
w5ayKfmKuMD7Mfh2erFA0D5olEpJxfVS7/4IggW22ahZRWjnyAdfSti/K3+Z
hXncc/xry68/9ES0ETZMg1xFTlm911zYE0YlQsmDC0OIpKfZu6JjtyRH0Mex
O74noE8ZMdxdu4ROdeoLCQoGkOEnQKkwtMGtviEPr+mMtorAF0amx9Jdj0UB
xLLod806wo0yzFh9Y8oD8i/8Oa8LCM9ywNIIozGWjo3Mb39pKZ57ObgwvwCK
eh7XQJWD0R5JzgtuTHFEF0GqftHO/u4C9sQeHJ5AxOxq6xCx+MS7GS18bPmW
/6lDrN2fjCNwJ43xphtzM3I4lwSVS1gL/hHJo4Jym8EtotmOdSgTBAIIxZgP
/mClgE0RTvuRaw/BTtxHh55HFQPKCrrIq8zen1/aFuFCASSn8Ol3eL+WoRDc
YoFGZAIbIwW0eWZbveldGbThwxu7S79397bpCH0SydhgU03lns2hD+JpQjjr
tpUDVh+FmGhRHpDznqrJaA1CNZ32w1HAt95R81pF2qc6cO60Z91JNHeAu31U
Ye7p57jeue7NfcKry8IT7b1tW1az9OxGDz88GLpm5k7QlSGHWywf0J9rgDkx
aaNxAp7NizBJlmdbOvD6vMcW2OWL2kWZ1L2S4Wm06s5pe4mkHsDcnxoTHeYR
JZAcqTS9r7qrhIQ3iO4bfBJJfQjiuEGgZojNEpCbi+DJ1oMoMO9diMNeszms
iHv3OtJ4XOiyojoDn/sy8DUP64mawXRdVaEyqaQ34ofPZ685UbGM8Hozzllh
KRE+qCKStYi2KAG5KJ9fXOQXAyF/2NmowqUZ+qsDa12AG4YprOZsQDsw+nXp
dSAu2OXb7hkNibtrFZfz/7kwNU1Jkt/7n+V8jPoArRTmTrwBu936I0sPSArJ
QuoSl5keypDF3RiKZvFMT/9z7+fRvROBxJvKPq24ScsPExwKiIWnPYJ1dtP9
qwLaDwpxZoaNoHIcaA1h/EZrTS/sfy+Y2xjFCLGg7vluzSWCzsoWCcdXKqBP
qo19XKkK2qy94x3LT1dMU/Umjh69jmdgG/M7DUL6egru+Y1yRvcYSwvNum5M
0IC4dAARWr2utTsP+F7N2KA8kmXjyNKzDMqwn6/+9rTiZl68PF42K4AW1FKv
NOUsBo/ebzmhPHVU4qw7GRNyi3CLDS8jLFZAnpCNlUZ0EWo3XlISk0Hh7hc2
fwhZZnAFGrb906Pto9v1sGkeeYqyoCApwtDSRrldwNG3RkcvHdzE8vvWATcy
R1kFJWvrhMMPwKztXPMMbBT2sg9BiQF/zMECSLhKRXS7iYgtMlN4amjKDnlU
ylzU+14QbW0hHEQ4LRRKsKBHdmfFQ05WJpKofZHue5nMYLNNJAyzCdNbst5Z
cFw4fPJG2AXliq88q5VQ4bpLuxQAVsK6BJtoGK5UACTLof1+yYbqjxWAzis4
DDk/V1DPovFhfrG/e8FltimteTGP7wLWoLeScBBYdBQNK4RhObMAhkjwDPjJ
ImBkw0yOQ6LPiUtH0OTcOMOPV4utWYImirCIiAugh0By1VtAYtnXzbn3xd9e
JlLQrnswITHhGHpjrPUiTBfv3v/HeBqk/SoePEEEEUN+lTclqIsU/U5NT6nT
6ZCwGCbcTxXarHQJJEhZ2HaTRICXhtzEYR229LTfgDrxjhrOhjGJ7UhphkYZ
jYoQGidGICi61ljxRywC//rlIbOjpuk317XqjNBpBz1rJxdR42FvbLY7N4iD
o72jQ/DBE1XUGycidtMATtECTgqi2AeXhMcFT0O5BBQY43qUlILT+COVPCG+
YaYsEyetxETt6T+ckBKl+0Za0ANT31/4B3NKxJD/stiCbg8jUqBLUkcEj7o1
yV9cQRF78UktoRUbVv06BmdYh0yaSTE1kK5cyVC1fOI69m1inL2tnqOFNpMC
xPP6Tbd7MHmsQjcTU14h0njsddsm2M7M6PhHmZvAbgudk4J8DCzfF7QlgQKN
kc36S4Prq/vpgMrD9ZoZAuDGdjDml9SNatBKLihn+cE+FjidOTcfOtAqMZyk
ITZXm1JjVKsCBPfp0gr9bcmja3iS6IohyX1O0ztOCGHqz3IGVnwBlVgl6xh7
h9mhqbLXSv6jXNIqlW05PosizbCWJ/0hJe31ipF5Bv3R3LQa2XbkbblGtvvf
ExVil2PbIw9N9U0pUzSa7MuOspVD/YW0KTNk5qLl8fAniPfZfelkw2obO3DM
OVfm6oxWuJhHpyRGx4hZvJZcHjhNMlRABUOrWzj0ijWwnKICQ6sKqb3LPCpc
c6ohIapW35gMZgUBT9GSQz1qfvf1tZ6R7avBoHkneqaF7NvOlR3P74Jw0+Zc
rnhOMszFeHHef/0P6ve1Yvzs/F9AOBBz3i5/EvsRfhIUHmx51f4un2zH77uf
R0gZzyEvBnn4qhB0lgcnyVdzGtOvgl8gzLXal8vQ1h+Ke7RXrYbb1i8FEO5G
ZBeklq+Sx8kwKYhYRHxiN56Gpv8AzrDIYSsAZukBi7qu+GE8GgrC9ZUF4TPt
C+/GsIks93BCWCE0to69j/wdwSm3vKPMLQmGdz0E1d2Fawfl5MtMecQ0G09y
rfkzyl9TEwPdPFCkav571bdoPPwIWPp9b6O+C58bm9bFHUHeaBe2zyHHvce4
QxxqkTh8HDar/e/Vj96R28uSp/eS23J1juKVCnBQ65Hl8KsOUHJUIDcMddGJ
3zPzHs8vDvr/brvKcDmfgHrRCDjDWbstPqWp/E6B8rOeG45dmvdqowGvd+oN
/gWgHMI48Pc0Th8D5BMUG0icOIMHusVIoqNKiM3xiEW5OwluPH07pTAc7pAe
E7BOgvXeKCPAjqjH31k8g2vQRam7nWEAD5RqAFxW/ofn7Zw5FH40F96I5c7z
uHROKqHmmaS0vjzq0iSQ7BMYdATQzWWVhwF1sCHL8Kj6FKZoI8Rf79I7dImX
xDLjlzKAAOdcORtTNCJrbZVO1U6PEV4yjLnI2rKYWlXZUjyB5GmMO9vfwwWX
njcMrtRVLmh60qEiMWwSNtQbmj1PF0Kw20GVYcbwjZeDosU6FGrL5sPZAfid
HFtfIhNU73x9Iv1eUOtqG3vAWBs78RNKO4iRIi6s2V+Y1ahwAh+UWXCT7dd8
T2MG2zRhGLUT9c3iQG56AWZGljfKPSGOMcZF+925ByF/jrDYlpcgtyiJbT9S
sPRNHYZBa9NLw/YFjXQ7HHbMEfxcs5hQOjQvJRlTFrKxgmrRGlJGD6TmTTRR
ZS2+kBpQx4DTFE5fqxdyFaRLwf1jGQRO/n6STGWG9Hg5zSZZqtadkC9IuHg9
JE/kLq/Am3Sgz7gq+B8JkGxmX8uzGN73n01i0H93fJAPKfyIh2p370o457PP
/Z33fI4fk9iY+zCuCrIzo+y6V/ALrVessz0EueUxVmwn8PlxiOTVbD97GDUE
pone21mMYQD1PfOTHvTkl0ui6Q9kluDdU4vPMwZXvyy/MSPnqOjE0zlEBnIt
FIl+ZHWcZKvfWFRVlDFw86PuNbKI/Q0CdEjoF3g1DwOLTjmH8muABCZ9d7gX
elqECrxwSaDBa8tw5Iet+l+d1Z6MlgFxn4URFagc6icmxt30N9Qoc3BDmbQN
A60S5wHtlrhfHIUy5JmPXXb1Ucc1s9ME5YEwtdJFzTErTffiYG4MxA2/Hw9P
VR+qgq7DeByzbm1/OOgFdE6uhRV4wg80HULiCzpPAqnl7dTTPXGaLkiLjjWk
SFcx3zg34xSSyZ9MuJnfCthf1UHcDluskBfCqER2N6WpQ6NfLkQhzVb9Hpib
9q7cbwbhbSQiSHtWFXdOQI8zpPeI0fEZB5Y43VQYX5hwEATXv/37iIEeyY73
ernvoVZqEI95lj3+WfTYtQRi9BRbu6dKCDKeuNLFMgaW8LLOdWPxPwzTss7l
qvhQqjo2qDpiZ8FbWiTkUDxkMC/BuDgzyU4fDWc5mNo+amStKHJsPj7n+H+z
fxom6gBPxQ7sQLDNCLI2LCxX1OWPOoLPLmgcn4xWLXo+HwCW4fNdlSvLf8Nm
Pzr6v+BNb03hkLQJp8KzL7/MkaPGGRoHyEWmb+2gMBoPD6DBbDICv4ym1qmM
wbnEs+fgEik0v4ycLkzejv6aPyvWHO2POHbS1/1XqcCwMNgmNihBeHLeOMsM
qHPhVhuOpb/ROVKENL6ir3VrPM6U0lFEK+IW9CC/OZ9u5l2RIP8D3DhHuxet
/Jr8NKzgg6PyWllheukRrfAJtV4zhit8LaWmZHPOsjHDee1Xnr2WWzZOhGkM
2V52CfLlwpRg7ja9vBTNJ6WQFJneDot4d3xMlYLEza466kxxolCWfB21zdhJ
3/xaJIsjjr/ikdbC8XS4FwrlV7omw5K5wy/93jthnxLao/V3q80ncfzMZyQx
+AmzIQoyYpNnaMYCSGXBBb7DelV9hNGucc6VicB4xp1Yy9SiZkwLMcEZAntP
NSxqP0x7M8LlRFVY9odJOxY/tzkLE0HJrM9m9fBx0k9JA67YU30vAfq1mJ5w
R4yUlegOKh9snMI56k06jzvnrubo4b/+jt7iyzvZ230peNEfhduMWxIU8b1M
Ua5VZJH6DevWU4+XqjZph/CM0ZfjNj/4V3tKm2d8h7PUElYJHYTcF7Gl+x/Z
Z3MxIbcETt+yXT0lPQP1cDrJQ1/R3ZjzO8nqeCK9DxioyIAn2w418h2U/R0X
CGE9lzdcppyjYMkJu07LLS3YpdNqY/Fdxc+NP90/1y8fmMhj9estYatgCMgn
xDDah1n4b+4tGB4Xwa5fNzKJl6Avmte7XAsJlQR+NFLY/3zo8llzd2x0EBd5
+Oft3FbQGVF0e7NHe+0lVwclvcVZUOmlGZ4aa9F/2GqOBw3XGHnXh8GQhun+
NvFtlNuDrikCHq+D5up0FOaMjqaNME4jY9vLN1IU0S8vBWQGGohPKvrdi+pY
1dCNpiA0gTU6xc/lva6lDhrCqLS1OfHkiXfjAT3VE4pL+nhCFs1LOcH1dpn8
sOuXaJYBfDqCZ0uG/RQBVUn15pBlwB5AjhekohRpLeGmf02396BrXjIHtkHK
1Mtnt4OONBQJgVwjTUyKNk0+0vlCY4XvNKyQirYkuTBxc7CRP3jzGOddB70h
ywHh5xiK8YANBb1NFR5fbcGQu7ROyd4GeFw59afxcha9mInIGNbDIrE2vONa
amY6W2dWHSC+7uYnkblgjJtzikoCF744f0oC8eZBa5z9tM5x8+/gi0PtCEEx
REr30cLMsVwo/oOddT11uGe/UUPVKXwfJQ8wTOmoEjVXRyvQf9i3rw6LsNG9
4/2nbCWnPoxSJ5lBV7XYc9ntWvtp1QXiJx3zJIOae1WGejDqqSWVDyEwHOY4
Zw/bgKkBdUV/EJiGaMuj4Pn+Zr3zLDxicSbVEsPSZUz6N9s76zhN5ueVNaMh
pTLLycrrHpG29VDRtryInvLTNeNJdw/gi24Wl8obDIbXU0Em8Pt+IRKw3lCW
b5E9s9jZJ30hmUqMqstwNlZ6Di/T93cL3hAg8TiEKS1Kza5MGi5jssIZLt+A
rhKDdi8hbldz/EYgdawczCXatzWIYwtdghMRELGopOkUq9FtXoUJyWttwRrb
LNepX1kWwZWnyRzwreKiKw8Mo8l2ZxpUKT/Pw9eC1KZ4wq9bTiFGayJF5e7I
2JMY1rrYYlQFTRnw7WKoPP2vfGsFasETncP1KefFj7IS7mqGL27uoumLqOcb
CPmHcUmTJVhlLLqFUzOnELpdWkiGkapb8oFYaIDOdpJmCeEVWVJnn1g4+DTq
NqhWCBZhyLjMtjlmd/i2QLcpm+C5/AkX4Z5rqBvKHl7r6fDmHmg1prfDG+ZS
sw2ZvOJVufXfbofq1v1UbipxUxn2EGayKRkO853dWQYxrgcIy5qNAKDUDbRv
vfYiZeD9km1KvZgjqLhh+ZHVWx0nv+kYbYCK023zlPoJ1lkd1JEJx5283kLB
u+9UTgrFcUrnb2CfrrxXyJZZJx1wJXP+T1gwVHvR0GFqwwWdNrCrZpRve7G/
jgzCgeLP5ZXTHeZW7YMkfJa6i0pfwNACLBw3oC8jJCHi0rLOlOGSAsgTjMqh
5cpHMtM3uLnJ7VPJdXAhnBSQCrxacwa53QSPNgrKbec0UMy4ufFRkzDa1paX
H1ADXcb4Pst2AqS9mMrBQbjatApIM4AOy4o6ugbACGXU1AFdPz/hIr06ByBY
t9liwVvpJD2/7iAgLS8tqlUAZ7rC7hqRZIjFrCaU9bSmnG4/8851rKxCnmfx
QUk+AjcJlAJX79iaM7G7JWJBp3Na6teu4uNLzcSceyAX+8zNkGlPLb3EJ7JP
9HAX/drcAJHT+CGa/rJenaoXrBoodf4aoE0xnLlbMTDaiq0hF9dOJsdxP2L1
AbUUMTUHkFKV1yKrOmYchnB++Bv5rcCdgzbUpeCrDPnSGGsSpDZ2ZBmV7CeB
raSqE/hO0kKjRit0MT7VTqZy1fFi+iAhf0t8KFYYQlzohQkuCxRduEKWfS7b
c79KtSIO5/4NwUQlG4IyUDXnKzPoruLV9ZHX1UNLyFA9ZGpO6A9bpiiE1tpD
8SetHju7NklG8XLzt9x8zoiIbANyeLN4PvAXlaM0W2ZZjHshtnsWkMEbJlxH
ZmcVU7R+1UNxdixAVwH1e2anbgjSCpiZi3QTYHx5o87hN2tCprQfFwL8PXhr
SWpr0nLrpA/e1lUTzb4QbdO++kGlxvjU1cLJmxUJ1bLIrzqH/replIyryvhL
cvZy5U6gJnRubIyEYZp8R5T7vovK0fqRpEKJaVd1IFS3pn2XYPW9zWILwhXc
uRYVGzt578Fw/Gp1PcngP88x8qsukuBeWb4jaPm2d34qiwAS/ODJ/42+YB/1
RC2g5MRRGxCekcWQAJ90brsRbvRgYT77r5DhDCTFHWq4fLu9uCr5hKaG0czb
aaMY66Zpa/YQS05D3MDW4pLC6FFAIeJB5aGhLc7yuDWXIohqZYHjxg5YaUEJ
sdGJ7PrXsHFfE6ePqU/dLXD0AyVB9JQkuUEcS4mvROyrqjbtNZz3Ne8+XUp6
px5W6ZbRMwN2Jo7OvTaU7yUqzN/FXTXm6yA+0x/7sAiuhcQi53nHtnax9ac7
uUocBPzCqXBoMFsJUzYEwc7vSPIhAK/cLLX+2qOMAgjh5Y1EVelY8OAclU4S
F3wXU2r4jc0m4oeRgqnhtF13KvFyDP5Qb5Ge6j4912lWlOFfOICuh4WRvwh6
3I/eKT/HjgTJ42fyE4pNTSBql9qrgXV8HZ4MeXVO/1uhwASA26ltewX0MB3l
g2guZ5BORAfNAgXZypV381FpVLCr4/SUZPF43L9RTOcby/CKALcjdS4eV/KN
gKbRe57uQektnfHImatUwhMzkOxOrxf6QGTgVbmbPezGUwV/5PPzYDxAMsrM
/4o0N4Uv3ZJ5Cc/MZjoDnozmEevq4wKZ2KRoME3W8pJmAJOz+xoJ97JcVyu/
WLO4oY9gxM0RNJmQQeA4B1rpWULqIcxVPenVMGU4BdlacPyYJEEvvCgcBYEt
ZSRdOwV3zHUj/rL9ofiNnbc4V1ac5bu4i16X/6ptRtAZMd31DK25Jhm/qr8l
qOanUhubWUAUX3vr46PpUBAA+GE9W+3TU1CSMh234Su2D+MrN25JlYnl3XAM
tuoz5Se9XrSrjVbjDwNoUVIbpMBMUSwxR2hswtJSwQRTNVqNaXumZNsyZkJ0
zDX40tsiiwmkVFa7q41JFXAEzNVRthr0oDylr4UHqki+qjIb3k07cRfnsaKU
2sBXjYeu6EcN6TsVGTI/xpyBjIZ4EXvDwdegd+RNL2v93YMoZwrR+iNAaz+r
KYlE2/XoyU3qtlIw8IUpM7rvK9slEk7XSb7g9QgaOjTRzmyuZDooS1czcnLT
zbOfX2/KUMGd4b9zYjKQRACi8+IN5xE8alt1LlryFxlsq+79TWN4KmWhyRDK
9TUIUVJ9KXq+Fz1YCZt6F7BzgH9gl+B5Dx3dArYLNODaZ8aF9E2hY5a2WIoY
sd3S42/Hw9C4NWIZZNZXZBasPGSnIAwux83Ncl26xIQqK/s2p0EeeO9HzJGj
YuO9vhtBokOBMbGG3TUb6Jbpyx2NWVHFwolLhHGxIFa20UPkvTnfFTF+q5qq
DdvTEjF+2DatA5LZElV4Z+BpqhzNnRFxU04fmKljeWe69tyzaNlMHwdBp4Ac
TSqs2qmYgQPz1WGyXLYCJvRAgftu6f6TnOs0gn0xNs2C6KonsfxFihRUQhbP
4E+Jhwm+JpGtxx47CsVdMPvE1hmLfVgcWL7Wzygr6hHP0Xqtm7XDf9vd1HzG
g0DzaVxwv44NJ04k6iC3ZqzUXAQuLkMoaOgwUazm6y76utmTldBIhOr9rk7Q
rOVEt4PAvRNLvPkIxZExPfmyo2rcPEjiVxluQYswnPp/Uza4pOlu1sJsc/Bw
aJFrEVov67mSbCZm8cvno43D71GxeAnQJwq+Lstqo5icAV+RLIeAK6wje3B7
SoC4XwmZBQHMK/vStelooUWbeZpdRCIQsRz2IdpV/vYHEjllj2KpPRwaii+i
8s6c9Mgn26MxjvkQ+I8VTbvIkjvv66H4ThdD1ja9zjPnCXB2cPlPTncYOYpB
/MfhSmp6URwVodEsMk+pMK/PFiBMTUPtcPemv6gpKrS3Wm+6R/wdkQphhwEz
PPdnenc1mWbdZcEwugMqNVkrsdNoQfvVUBjldjC+NXGlnyQagCAJgszxhdo3
3bQPZeID9iR15Nm95kdkhqSMEjLKcVIHhknEEvWFWz8zjPlhzEAE5DIi/Iu9
MMzXcH6BiXODqaiwNQu8chHUZ/Knrs1HS2UA1IRMes5R1JVcyGyZax+OxhMn
t6cLC5r+MxM6oqRbvyKldxYm8YKs2sTPZgIbVobuoMi75OjjA8jgYM65CW4E
4Q1WumbRObNCdTSp1QH0fAz4nOLdCZLEdDolsQlpQT7R9/a0pxTPg7CwkjkO
Znd1j7+aE1ildcbwjOG1zMNpbxrjEsOa0Fyp86jVD675ltWMylr/B8nS7wo+
bStq1TVd3+VCqiLoZN77XHdHtC/hllFGARqeXD856l7SC9Rik2ZlfKdqlmUB
0QAnxmqRQyHyetq+2XpS0dZQP6kMBV2Ya0LCwwYNW5YymZ/MJfMo36l76BLd
yb75r1fs5k3bci2KNkzfcQBJ5Msvb3ohOJ6iWdxI9FQUcE5w8Xt5DXXwKnda
CWE17CR5E4tLopbq8a2IZZ1Sl9X1+SXgSz3c9cZ5GpuXe357lmuo24AcfEzN
xpmYX+GOG7YXTRsFTdcv6XY1gEUiQ/KnxXYW8nZfVgDRNoBVIfQXrVmZ9mcy
O093qMmAk4+uiah6TXsu3h2t8sUo/E2EAw82w8M3PwKDxJrcDydocMJ/S6Ae
FNZ/PIYaxzhH9dB/c06dP1JfIO3t14FC7ztSY5FV1GXUwnIWT+ZUhU0/2HB3
h9JosTNQW4HltNiX9T30mHoQ5PhmMnv6/c0IagL2Tj45FS2Tuekd87qIfSJ5
yoR7biBe0jaPw8wH7OTJiy+o979d9VCY824Ikr2UhcwVmem1Ex8vL8a/tP+7
TUTSNamRZtjUB7vpV57wI52KvN83XBGM1KRweMnBU1CMcDlMxIpKPbRbQ6ui
7qvy/wz16V0bxCXDYh3xaH+FsrijV99nyCaCg+X2ygJqu37VGqJgItOFcNfO
Iej35GyH2V7HXm8Yq7zwd8A9+7CT94s7mC4CHinVELIrqRH0JW91FkJWB10n
GZvYY21vf+DKXZDfTBXwS3TnSmCgf1eMZm9o729r24rjJ5M6lMLboYh1vESy
yh9uhzeuUpr7/SJtW4D0vhUYegCaj/sTGJzKjUp5LsJ5mt69+il4aVmSEZff
YVhDEFBdr426AAduW3x9N54txE0IDllhYmFzCd9Z5wqCxLx+fRmkXjyMJXfN
m/r+Sjc5OA2rKQOjFezUZb0ukhmdfas91Qywgqf9YuMdVujhTAwRdLerSgcX
VdJkj8lgZ+Bs8PvFxWYqBhsUBDCTLM+FoncSVF8SfaUvtURBYFf1m8rhJED2
Lx4jyYcGScwi9Nl5SxwJXTO8pVCRhWzhQpBViae9HK896IkQmKxAs9Wsb1rb
Nn5mslffiYlqKlqKcQ3Ww18sYapklARe2uEe5x26bnxo0e6CwP2+BiMz8SKt
gVqrO7mbkAoQF+wDXA0j/27PhoTho7DZV1KM9bKwdqsntWaiUQjTjwJ7O19d
WFig5xbdwjOTFu80fK6TeJMZ4oZfQ5XUdP4EbS3o3/bNaXkDx6syJ8tPBN4/
ohI7yY90GlANQslSKyK0dIJm0dHaq2xk9hjCsHHPJzQeHGaCQ3kgovw104D8
+nltQEmM4jhb1NuFx2hy1eOJpPKWyillS2guGczgMGrZkl+divaZdX22V4t6
igORk8aZmigyA1/Bnc+2GLq9T6ctzu8V6Rfx6czqs+4VgCNwyEI9gOgzIK+P
krUhE7cWVG1Oqnd7b9bsSuNk2ip6yFTEsC045DgqT5OY82xJlEcf8rTHwkzL
4hkeE1orvb6xYHw2uTqs0qWm48hNisUMFuLXRJBkn4MQ1Lk0Y6X3pgTG07/b
l+lNrZj/HE36iAPG8DGNrX65XOEkC5Wzqeh27zI84YB6Au+7Vk9me6qY8KKi
VlRKWj/MDeVC4cp5iSYdX+fOU98+nvuN3UZjD3PxLrycnLrhh4U+3htf9D1s
OU+Z4MQth553HBkU2VePyErd3P7E2JrOzzzma4+vhjsCkMAF3gEiiNK1DBk5
dyX94QS7j8ts6jpI3FvKDBG2FoKkCwwOmx2xUxQzp23VyXkM5/EkxV/zTWra
2G+86qS1l5D36uIJr3idaUasF9cFMtu2bGEDFa+u09VjWhhqYE7Ft+/mRknB
6TDzATjJQM/pjrSWPq6p/53NB4uPdGs+F+PlTdzPYegxq3oc1W9lbFVsyp4P
IVHMcdNavgTvV81L45C+wV/f49QJc3PedviSHGo/apL8ehwK/JtwFaFdm+MD
cQuqyGMFPXalzLxRbL+KEIYU4NV20K4lyYdoBoGQJTxg6sBJlOYakV8ExKyG
6i2e9B+cqsITZ2FwnqSJbqzurBkDF8LxOVkJbVqsDmVhcM5nAh/oMuV5Zy/x
ppuZCh/EKpH5I862lapLsLEKLLSCxPkXK9K7Nyj+5j7HMAjFv2x8GWkyV00t
+OTy9nXSRb7o5CZx1cEJKeYYv8unKpg5ZtiInpxxhySdVi3sw4tOKRYqhnnh
rXzSa0e4cKOdHLttncR996Byfy3Xh7P8AnzTf+4wAIZMGpivRSgKi0ALJiwu
Vtaf2lpLKQlD0sYERtXFk9WsIgF98GmxvKvsvVhte+gdrCzcGCTbrxvAU9nW
6++r9bJeh+ZxNEDMg6Z41g6cUc2mUxozSV2AlMa4rz4TV9otx4AKW4e3ghds
NAMika3geqqXviCsvWis3qHXaOk9/yilMURcmxCBAMQyGNAzSNhLvxaneDdL
Ve9XqEbTWcSMOy5WKweLE36Tln/OaT9wcYibfFKvA2Kc0VEiL0U37fcep9I4
ERdxXhmfFyXhYy+ilM/PdQ5TtYkhu6rkxeXgxLk5I9xqhbeakoxM3tyCusbD
PRLrYwl7HbUhq4rDRvE1ox38yEwqPagVGQsSzjTog/bXZqno0tI+eM9+bEyg
NqxwdT1oxyUG8UWGeNRutO8oM3EumuNNyywNjuDx8+ztQs+xsWzs56lw7SJG
K34D/StXKwm3iidNGUE7Gt6G9Qe4jat+vsEqMXFFVRdOH/s0PL2bp1m6d3R1
gGzOvaUK3YKAi/T1ZvSyQ5eWl//j1+ZVgvSAcJ5VXl0QQrXdImNgBkFFrTFg
4GMX/PFAoSXo8SIZgI0Ta12GJaljzN5aAcLYGy1fPBpsyGsg/Qdc2TWPd5Wg
amIdztLwqNSH9QJ8NR5qnTCfo6T9VPRKSNfzgEVj16EuA7doQvYgKD/LHrjQ
lOuYweYxt8OKc0b7kZLpOZ4WBElQxFLBgOh1YN9gbdmh3Q5zJaqh7AqESM4o
8aBFyBxLDkq6HEkNfsJO/XjjW2ssGHGGGuYm638w2I5s59QsRlsG0bS3ntG1
+gx+FYghuZPSTWk0PRvQDejqsEcwY+P0PIEWXOvCTP56JMkiRB6qN4FpXUDr
y628DtFDWC0hVCKmbSar0bNRswy6FFnEI6+nUl8aRjyB5D95eF0F9qnJ44fA
HF2Tdhf9X2+xPODlEITXb86BmlHA3PrdT9lz4S5Ij0ZV5BdtTWTcFSdosalw
vXkXenkMW22iapsF3XQWDcQp5isnIGsqm+w0KdNP0VT6aDnVPlJ0Tn6ieWq3
kh7a0SlFufSGm2AtJRlMEiwzmo5Kq7HL7MAesg0h2Z3yE8SqSaZJoPrj0eWM
ZQeZZBdFdmoFZVHvMbM/DhwDslS0paYM5eOxz/c0AzJjYyOCKZflSBfCdlsu
wXD9b+XDQCghalMdEhHxbVXyD9CBcuNZAZ33KtIwKFz3uN/QXFrAepdy6PWD
6286e5RqVGyQVgrZH3hN6+0SegZG5sccja3zCubLn9NpuHQHAfXquW4j3Er0
qrSEN28x8uN7yW8xSfPN6rufoyedx3zYcbE9v44kgd2mf9+blxyaNl0/mVMw
WBAXPQD5gEd1amImLgrD9jjV8ePyB3v1o84s4MdRmTnhyZKLrOzIZngZrT6u
FatH/YQVRB1hTjFLAVFyzrn56Wy5K6wlSubpw03Q7UDW8LNaP54Or5fWAtxe
PtoXmHk4H26DXWtlF7rS9tWt9VZAwP0pjPC9tKcQ0EmvTIlMb2Hi94zsFVDu
xhIDH70tDaogg8ordWy5KWBWl6yRxKX9urqzxf0xF01LXJoum+gmIOxpL7Aw
j48Vbrm5Sf+p5YioZc8JSE/U7wEfsJArc+3BQZnTHd/EtVBbzcqmDt+56a8H
t1Rn8lZiXIY+oZisONnsRj7eQOJsTVl/cTuogg7aR1NfUNIk3Ezo74gdcRxy
QrszP34OG4hnzOfXd/S7wnV3KKHuEujdFn9Wjlro7hM2VrJe/7Wxd8WW0fd6
qBoPW7T2beaMzU18I5WPNOBdsaJokwdMw8jMZoRgpZidriGDX80ElExheXAN
NlLQAi2Vdn+u4V0tm1MvixNAbxPSoyHKnY7AcqUcTRcQJjKHu8Fjq44uSuwL
gYHURMPmZei4aeqGfy2pBqKd/yFkxEhxIlNc9zqELIh2lPURcKDZtm6zqjsa
agJAwUJSC8ZbwhAcAwDtdA/jC3hR2p/z/WPIbiojGdJ7ePVQrWFpiGrpdm7Y
7NWUkHtrVyldJntlBuajszDKCBHoFTlPMyp5e/cPu0LQooH7weOOMzdrXzvm
M42ohOy7SpSuM7o01F1j9oqEVyCgs0IOlNvvGR3YZ2rifDFsa6szZGSJkGvG
ZPoyGv0hb1tpuVS05gZseMsBO8VrfbIFrViDS4s2RBissLwgsWRBoTkHYEOO
KwBZjCXSQuhF7fEBlkjgnL9D2izec+rFrzKompk3zXSBwlCcADxinZkkldup
kkaSM7Yv3tOvEfuXcpF/RaOWXH/omd5vQ1/2UdX8vSlvH+iMreQIDbM6a93B
DT6jFGH32t1PxH+FwiMIaKe64fhRzV0+bgmQ9HdyQlAcXK2hj75E6G7NzpA9
whLLHLYkuIrq70XS7bV3KM49Ty6ZKxpcOrF5FCIOIE4NXBKEmskQRFhjPGuC
VYQe0urjRVQ7kFCBZT7jjVSNYHqChxYr3O9VPYwlISHHabS04baFxReO4odU
Ov+MlNzH1lEllLlkOgj955F1I0X1NMx5iCLDp5XAUYY7f2NQNd5cZnnJ2nYZ
lt2KY0ki6JCIZ/Bnabf7uStlLRtzW8vZFTpW8aNj2h/11aB68CjEe1SWeNEe
NJG7YrfV3y+Rz385XWQYGxeYyLM1YjgMz3zT7jkTt7OawQYs3/Ab0NVuzSqv
j7nqFyRgTa7+9qUCF6v/Zs/oJrJpQV4tWG1bHYC3A0uGyAbQol8Id8csz5oU
3Jq6Qh2DQ2ARTWMZDu5JpDgXUraqIjDNaC5v6prg4zWJuo9gKlOtIE1/sAal
RkCjPwbieyc6NcsWH/utXsF2O7j7KPczJJtLVlP4ztZR+m3SB/uL/BVPu0QT
uEDqDU1zQZ3EkOLChgaARfhE9VFTfi68aZvafHwpt40uM+V4ITbui7pFN8dd
BT+nOuEXv2wFuHiF4e8ptlmZ57fFDb+NKz77bHlJlTlezv5AEquPn9IFH/DY
otHx2NK6wXVu1d1wFPVMDj6tfUkiSESmUqZzmgD1T1z6ok+wO5kDLQBlUd65
jZUHhTsTVpZefwdB5e4/kyRxp/sdYvClSitQ0ZoNOItWV6GOs1Tyg0hiFNlY
hPMX8b8rhiSev9PZxz2jQwvtaAjzrBDtXhyGcpqVzao1dZsABOQBxALlWijT
x+OjpxLZjHscw0Dxih8TZQxnHsU8I5u6MvIZY4J2tH/Dch/VT2r/HBdQuDOp
ZYUbTIervv6drXVXcUOfWjYvfLB/q1WTCVC64De3htQ6phB5SeGTeby6NLPg
MB9sHcOWH0o9kcRaRJCqVBvaLN375NCfh+TGnU0LjI2bzrPsCXJRO7Bzq8U4
y2tQs/Zi4lmaA/TYgIJrcCG9hSeT+eGHQzlySfwNJGb/+DC6YQ/K44JSsTk8
cpkZSbmsjeGy+VVqXKcy6aERuz0M9b9tTqw/V4QXdtHF/k7E9jeAPDCKgG9d
EeqBVY8i50gy1D/ULhwiUDTpub0op7KRcTuW7VqoXaG/hYWHjRf/MjjFN/zv
cZOMgMxg7Wsfrtp5q/AeIqE4O9P1RUwhd3l0pq8rdannW8tG0nTsRavJnD1t
SotQkcSv6uvjBgMT56R6FdkELs6kUr0tYxyBYxpZAPYFlwKtjYgLrJdrTpbz
smp5l2dTGg0Et8fRH+nHh07D9HYmwVWW1Dt4NgAwg0rqfOc/nruo912yWN6C
yABkXBjvTF4h3SlZF6T4pE+jOTqm0uSaKyh5FO15YcuLu9LmiwbsgJe7yRYE
WRm8/4ICLTLBji+MbNraaUTU5YcvQhZDAsz7bXKP9kfH0SccvS5ll/5OreM6
TrmozpzGJWjFMGWz8vlij9FFuKE4MsNQJ063NbL06j+P+WqMG2cGp8M8qNMh
eT1Vz1drvYjJNt96R3INeUenoyfH1pnUK9pn8FBvi7BRyaTN4KzNUUliDF28
t93xBNl319mra+MAJ3Yyzq0MvhReoAy61iPv/59hE22zX1V62oWE6WZdCnUE
NBKAFLlnZkWZom6iEbj1G9rp4T3sg3Ouv2DVSBEk6HolOjVi6NYggeAmfeWa
jmreaSlgLpOYxShyRUN2BdfZv31Zrp7gCPHm1v7nbgIsaHCdqfbL5UKVIV5+
VHlxG2n/e+Ys5z6Cvu9QkoAYbYpQtrNeukme2MGd7YtwFKgBXw51HmmnlMkC
7e0u18gqQvMlH/EUxFnxiw3l6eOp9ubYX6SOLtFRp+rj8voFU+rTQ6USu1cg
b47+ViQCh12yVZnaPk9PPR5/xvkyUJevIPu9yB2V7DcPOVPQlNOVt+GRMBts
9INrBlFN3AHc6F71S2OJDg+Vcu49ZnuQ/FKEB3g6fvz5/XR804YqnqpHXJvZ
dEG+ft2KNNr36hyZzPyfJuUlXLN6Oxp5zr591WNG9bDdtbKEw210wDVF+lDO
mTpjGn0SIqPWXO+v96IU/LPzVzAgVp6FlUNYFSX0dF+vqWCv5GHBW+2UiiJJ
yYFcTOsr5rtxEzM33VCbrkXEeIFHn6v1vMCnQLC0UgSQguTQZXkro8NBllAB
zdYD4eDUsuR8Xxhg+Cp7JP3sO78agY+lHbiD1Lr6M5NjbSOqISDuvHHTniUK
5Z9D/hRK1PuGF7jcczVbtK/xyRgKjX5LGclw3FHkTOgMHCNVjrC5aAJ8iBm1
fM5/iMtoabcTJ7knl7q4/pwYYF/I7zhA5Xaku+vdkFmEN8WNLnSQolvbPSQp
xQLotkuyuDmvB0eaNfdJOxkq3Qj19xwd7BWt2JiApVxW7As4oQwye4BZSKey
oRkUxSC3373E4BqHo6mv8eHLLQSC3yAK6Qj6apai2aOFqOOZbusFXuusXFcu
e9wTTGx3ms5scI9JctoR7iz1K8tXs2dpgfrtlqqHyTe9R+R+Moj7X12rR1ll
rdp+4xEgjLp+ik6RQ34pwV5GiA7C5hOd4l05ts+dVBvAU+gjNYRbbyxuM/Uz
MtwiWP2M8fjMtEzl/FSvMjWjnwcczdFWbsfZ6tz+6zn/fp0B7PiIOMGwWQT3
4PEROSQOq6fl5tsE2o4BaOz/S1d/uKtLOeZeLI757F9TAbL7Lz8DrijCUqCz
UT9i8y9oKXdL+ADYvkgiYYqkX8ZQaDtW9RdPr2VlP4S5oRF4GipDIfH4IQxW
dmDJnKGeHxtqgzAEbaWu3XfMpbET/Kdy11JuG4oafvMBqXuFdk9RuU6j9NW3
2IdC1CQRemrnKWT6PHmlPjwxxdFEYnbp1B90Ijf2hkcISCHsaL/KFCxiZhG+
L97+dEqlzoEyVIqDhQH140JeL7hN3cwuCxak79iN1unEBggNOtUFKRkGl6XN
ChVcRbj/S+7QqEUSPp+N1MNAoW9rY2dBHAC4eTg0lk/7r8O9RmAoUCEjWiou
/rLkseENBsKyQZ1S/qNd5efpPGOpmsCd6VPRYn4R8zcByG/u4BCrNWKJFHWy
2w3L27QPObTC6lnU78UQp8VOBbq0HMPvT+3UTb9cWCZaO6x/UU3mPnVnd9DY
u2L+BPi1LPWa5GuJ/Jiz2JhX036ZA20t+oJqFBWqUTYlmaBDcH3zJgVNGDfX
n+FauizFSpM0m3HZDJEr12qlPK5gkfVW6EyxIJOZrcHXxH8g0AwAYEhNy1Wb
HkY++ySV7B3Jm0sk6f0D+kKm1vYQ/ygomVdTFvvMcEPJXIZPSUrnemJ2XoJq
nS63+FEGCtQL2BLlQbM6WRqqQnYv8q6aoJBUEldq8LEiMNqbvb3+JU+A2NvY
Ohb6qDzOKhBfe4cSrkmqnSjw0s3RbYLXwqBYrbNafCFwScgvFC9IhxxpJbOG
A+PXOUy4XEZ5YntgTtkdsgvFX7tqDM5C+Ce2iaNwXh2WfXnPSxvTN0VRXGWW
UU9UzwBlXNZNmz9qfiLWzjjYtX5qXUdHlLjZIYFT+1L3yx/XAwtsMFbwkcLE
qoVZ/A9A9G1t3JoWxbgiuWFzgwV+vaCbBTxtBwF+x4KQURHnk+msq7+DKQhr
ryilCV5Pku0BLBIHygb6mmtXmoGEu04uN7NZmB2SKLrsTdXGrHYrbnzSji1w
o4TWlsE2ankFVflybCCV/I+iQPLXqAwPDgegOqPWcAQoRD3Iw90KdYO/yTN0
NpSdo4/LSVs6i+xIKvOwoP+Ok9HJxhzkOORq/oU+Arn02BvbreNbve9ctB6M
Eqatr5RF2wl1cWwsDZvrC08KiuEEwBRvwTbQzY5rOuIKCstX5tMVf43JjTvN
Z5g/xmGXorW7mReoOJqkB9Kj9EOXnqEcZ/0CBo3mwrpDCINB4fR/ZetRS2yI
q+XVcMzraWcPP1gfRHbOVFsREOdrG5SiuFLlrL2kky2Tgdi4zY+zdqdh5GoO
vehfnl0H8XjMwlglo/4QYTr5SsLdv3E75QfoXCCQUsgYXr6G+3aOe/s2hXNJ
VUK0GP6sLrVgE0MuQBO3ftZS04RKh1QYVYtSIFbvrADyf+bjuWM9prtzoA55
0eDl0W3C+GZhxsRlmTDbxILiuNCaWH++K57L081vePVMrfW4yZlcuxJ2nbec
eKVEFaEhYaYkGalTaPfGk+VjY7jdugcEygMeuhsdsN8ooklu9/UmxxDMArVf
VIq6gCp/7ktlgVYzPXOPftCWiXVEp0LG0B5KRGj7hXlrC4aHAcjOmEkl2Kv7
i8CSRZeZIN2XTjvIduSPrClmWK84xpz7Oq+wfK8XPXotMnli6CIQf/Kfwlsx
cEV+Ag5Xs0emBhS1iD/UicWTgt+3roMMHno4oXa4me6sVwmsHa9ORWPM6vNX
2K26RX0IPmy6Cdg0iPdRsqNtjgse97Y8k0KrPuwW4FGk9TKAKfHUSM5Lh5LK
2y6eh3aiELhU0YvyZH4E1G5RhB91g416nDoBZ1diCYsvhf6OIAnrTwr3J3Tm
/b24CfHfNgx9dMYYbtbeg2zkR4W35LaVYQhEA4tcivYiT0awnyCDFv6pTPCf
crg8qemUpp/w2goKHHNXTgeyMZxb2m++7FLhZBjjQ7Ht2wzb5sVHDoOuXfLG
dl39Aa2eTTuV47dwT1H3bb9kBJn3QAZSHx3TbRUTrjWsfk3rieNwwQ1gyDkY
voxx2ypsry5vtn57E/QsFvF2/nBQxaR2pnyezr5iAq8akbldyDgdB4duF/OI
k9D0C4cL7gH3m60GQQdGaazamMRhBwbxsu7uQo4ytVzFs7ZZjQXPUe0sMqq+
jn9/ZsGoIco75ho28fvJmPnOnV0XCuwlWtr2bsk838y5f+uxmxpY+VfMOoWP
jQ4oZrk6f/cn9YciOqCkWQMmU/PkLUkv7CmLo884+kW/RFIgVyA9uiEdPcSU
I/pPTKf6AVxUnjJYXYAeAAK6d8M0uuxDKP3F7a7lCb91JbUGnzheuNCSHeYL
NmA81XZQAvUiaoPczYzSalI8/8Zpvs29s+1s9VdIErfGxlH/JmwqPZhS8vDN
IQ4VZF69MpokHO/IfOtJ7sdjmD40ZOCYaUW/xAbbF00UzmfpGSjGQ6hJoqfc
oyx1U0Te8/aY/lcWw7RsvbWrbX4XdSsw9RKUp1GrfQTR+PZplFwGekXfufod
aYOEQ1KJL4BX3UVRKf00j4wDN+MtiAdFU+C/oybYtkn5o4RTQF2DPndLFyNa
McJlnJACNmPIqyFQK5Z9Ha4RR1/QhWWHxXfOtB9vxJJeKLjp6TQp2nk9VagJ
H6qAFxDiGe1FeAssikDzC1eWzWhRjr4knBS7/AN2LI7wrikupIDSg5k+8uPd
p5oiO0Z7SGay8t9o3/wsvLDSKqKLZ6mmX9CIfdGmUT/WUMuqsrLHc/CBdB9Y
cjUvfWc+C6O0oPVx6eCIw1wvJtY2jrQSLOXWXwzGeqQIpSbnguln4wOLoXlK
yBpydJQ8OfkCqyV005u5KiCrBDmmU8rgtJZ4kcz2+FTBW70m85aj9QEl4Y5A
SrGeJ2gJedbbaxsoELK1OvWnoCi8Rmcyjqlwc5AjJK0V1iz9YHsA0Hoz/obk
xbZY8f0bg7+ljTsbs65T6BAA0fDAplfsXg9mK+yFVcxc0bhZKL1L6/r1S9iy
6zVFjfRqWqUFOnbElaKpIz+ptOVxgBSlwZhAlfnLjMj2S+fleo7atKTaP+Fj
9lUb9y026W1gD7MzdJh2BNofip7z0IMyI370NpZNQiYr6uJQ68p/XmM+sjO0
eTxPd1N3YZMrJHHHgpk1P9DqzYzIVWXYT/B4gf0cURPUGVzaww3dEHz7wP1p
w8S2f2IuiaiKZUlL5Bmbj0rZbPwWokMVhMepFbluaAVCRZr24Yw3Mk+Xl0oA
Ic1MhsLqc01qrsLhLKFlDK8nnRMwbYhcy8DAcH59fodivh5ZZY+R9BdUvaPM
Ud8GhksYJGcBANZn3nDycAK6zJjw11XRGZD61x/c+19lC2E6Q+CRl0nZUL/l
AG3ZjrlbRx+cossfF7a0cccEb8advo8nZiYh9TZKvs9hmmYftmwdY8LKuOm/
WYGaOK7t5p+0MwGdeQwK/YUeL5arYx8tZjgPKb7BspuaprKqD7eKojJi6CxU
Zgl9lfKKvk2HOnt3Rx7pAPA23tmzpHgtnlFzvIIPAyVMSn8TYKa/knp9vrqE
0MdlCUCMIjL1amg9oR3dGiDvdCPUuWTzOvh+YMK0ZeSoll9iJ2apJzq8fNv+
GGdB5CKjuMnQItiu+es9v44I1CyAE/obDae6+EXEzFJHjaT464RkolzO1Y3n
ZH7EbvvxFB5qinZsBnIns7IELr5Kivy/LVTEZgmPeI1tWss94ePLbDlUUKU6
MsbNDJ4cvkY9snlNXgAOyU42hDHXDCJdcCSgQKzkE4kLlh27eOEgPFpTo4TO
S3XQsNNslqVUXGzIUUzUBLGv/w2NgGe0b2wef/p6jqvPhJoDUATnbevQMC1f
4ZLfQsQJ42EtUcAfYhgzXqguPD4tGju4LiUSAiDEUJfuJ5p+jpXAz3Q5cdw9
a9HNg1YYTaFrxdLS4Z8d//c22DCrezQ/jyQot4JFPjfSpX3KtrH7BIyrvx0f
mWYEASfv9SPTZdu7jbV8vqB42s4Cbsz3KUJzPRlEGbS7slfLq93iUuddYRbl
zsyZCJigkDAzRIa3ez6DvSdqhxVUTOjG5TsVoi9D5EZTAxPVLC4Hgikuo+Lh
1LsCdHXpm4Flb0RCioeP0U0Pw6K6KOdlwdMGVbexU7RTWTlcD5f/wX8LKoLR
zNva3dOYECfVGm+tDKQrplX+Hvw7bOeyRCABkQ2rkY3DJ6idO6Oga0bhNmDJ
0b4TLDaXTeQPil1JAy7uxMLTdNr5kroDS07Eeqw3GXJkQcshqrRhXG4lQcop
NGt218ZpimVdcIqHJmU16GLeLUZW1KkvbfMdG9H8uN6TGGdOWHYROYLb6wBa
iNx8IefTePmhsW/jTdAImpiREu4Q9ylw0LPWp3VWGCeB9IXB+QPEfR+r7LA9
KaWcwBKk5jiyzMoWs18yWq3XdzraVmcYNDhiwnOZIUO1xSJW1XZpGmueTUjM
a1l4UUluMiulyX2JqXJTqAyCDaK5gYQb/yDSQ4btp2qP/DeB0/7ADoqA0ntZ
dHIR2wAGtkcOueM4B+RVrChWyM2yMe+DECrXNUhtv7LcTjOzzIjgWRgkjZxZ
cSoT6ZzzcMDhANC9IvIcAvxwstrr+QfTZt/lSpcsGknSqq0CdpOx9nT7tTBR
DxMp70Zg8v/OrOANqUXYfMOA0sDlw3xJUoO+IVqwIu+BIDjRty3pXKZLhn/A
Ajn5w8wkiZLFCHCh30D0Cn7P4b7KTJKf1PqG+JkDwM09WmzyDloQgVfAaXgp
cczvPr6fG8gSwSBfhFmtZzK9juK8UBm7zbbp/5ZCXKSov4d2+gdc6MkZh0HV
BX92++xXegIf1nigqJLb5uwx3BsGjgYZ43d0W62qrTTYghyinfuZBu1NGGvj
ti11FbIr2B3P8T4uO35yOssRkJynb0G07pZsUB9Jkj+zMJfjIjVLDGV64nMi
ZJISz3y3W5p0bXHuGoFe/UH1FDsq4qI9kKW8jN5/5tpQmJW3gXDl45HGCsac
M7eo8JVBpXTX2Z89XCJ+QFV5r20nkaKgCiunu+B9dwVNjXcLQ4mUlXfShNuC
VCc4PM5NL3VMIMmjLqkDn+gHILNkm1e/y7cU/ms0wE68+bkqK+FGLn502FN1
ULKrRIFdDX/fm+qf+azCeuxwY2BCPGngI43rHjC8pEOjaHOiK3sJw0CZuPMY
lgwK1OANhD0KiWRdwgF/TKBMkaqQrjR2Ob0vlFfY0hjyRNuXds3ikICKpchN
VrCLj8eNtBc9OrNcJ9PWKVgZBfPlKbN0FYhIi9qLEzUKSjpHFFEJ3EFkz9KT
s2lAIXqS1Az9DUrlAiz5fCAoZOX5lqcP/bLWGD5Z9Tf2XEG86YyojHKT/BuG
hmEWHdPs7it2fcNZ7XHg0OOuyampc25N9I8XiUFOeEN5e8i2WVYX2rS947WT
8hKnWYMTYlcNt2kFJCPTyd01b3nGhuT2DRDiZGaHSg6WZRgtCzV1XHLj/R9J
Ksyi/EX8s/YT2AnZAZg3CxsX/4cKAOoYd+UucFs0ehweSFmW94UInkhB/BMT
q2lwfv5qkPQKIFnXe5pxLVoE8DgoVIt6Clh6VFKdS+tntN9oUD9uRYWgsdwT
6bq//3IWo5F7owlL+5ra3006sNnBhPj/ushuS4yodAn1hr7DtR9qLCJrAfS+
9K3GmlxVpdqGpdQXwcc6LmEUiSPvUcEqrl5Yx+/2w8dtuRcwt6YdUlwkjvCJ
Kc+QpX1n/P+2y0/uXSJbom6msg0WtS45r+9C61M4wVpm1ZDChov3RxFRUUiK
UQdMs9ibJLl9+vL7sBiHbGCAG+URct+xoND4zuqL/l5juprTBIjxsXh4M/sm
7gHj/CJpah04ILg5JyGMKXphL3qoOvR9wDFO+7x46rR4Eo5/OCEEouu6sMeO
/RQNrKAhCu92Fuod/7w9ijcNspxhD9X6Q8gMDqmaQxseFguQt6/ReACipjSM
+3B+OXubJArCHie1mdZPSSth+E+9KgOm3XmhMUQYeSnlpZZw14ARoHqej9Zp
T9zsrbkLHxGV+1n4iAM1wi+vFRHecAS7x7rZOKhTT8nw00KqSlJ5q8yGokIz
vviFjeVfGMez77Y/zJvreDZ572o1rXLrVGHs38/WLPbDx3gQz2DMrPFtLRJ1
7iOaifnTxy1KlZsMqhdPTrR/Id4bkD76pibyP3GTwVboC6CHbsQAyCz9psaS
3eQVYEutqQXFmLwb7gkZ4tU1Dw0CLAKdQWoCph8FvtIISz+ZguNstsOM7EiS
RjJz2HEWdAjYM9os3DiIjt7qBU4RaxeQVhY6aK4t9mIkjqIsx3OZc3nznwDU
BxgCmr4cbpQkz7DjDMtG2sjxtrmh1jnwu7FMJcDSCnuy/d3SpWZviLuyGnU6
r8UVkR2cNveTvOoKOTsvAvwuTjvAv5Bs6v6fMdj3c+MQFIVTnCDDmNm51EYF
RqsjcSyPmTv0tWZlEBHLeV9XtDtR3U+y4dpRdrLgXg6kBxCB1MCheRDNkbfz
fWFNzcvuuYG1tPGZ94jqIqzzys3DUhryZFfdr+Djs2mx8dDbO9MwPslwfNdV
nWWIQ5oPewN/jsv2CtO+FFvNkYmm8Fwh3ynb7/GIa1Ea0CAw/NVSGwMw5UQU
WUyJkRQeBe/Sdb9SwYxympnF0e+eEj6iF5sssvDuQ8Rpcfu0/J002QZkma8w
4m1YIiHgNam0IVO5gKdWVaIPka7EysmKcJ7i9/lPe3Y1JweOJLs+b/A9hFBz
DPxsAqsLYYpJTeGcsFjQLzdvdFwRTnREVOPHe3AGXdlr7kF/faZiGBuOBwgG
CbDI6vnV0Hin1bk39MGq6tkR7Ycq+ZldarU/i0tCdADcM4VI2OBiEhsQGBh8
NgT+Vf6xLNGX23HGD11c3BlDSjiBDlAt2FoVXyr8mI0XfLBb1oNzheEhizRM
bMzUXaKZAWJ0i4YOmLVATPuVCBGONSsSEDJsfP1xVZXbbWPn0UgYy4kU8lZP
HmAcdHYZRPjQPV2HQ4CFIsLMJeuBZ2a4BU1woquwKtFkDVK1Y7LX5Ok+5cKn
DHQXlezckAz/4wBeB5nRGDpiMWsDuELEz7U7pl11fDmidM4/yBCqPIWubwn/
SB8t4WHaco/N8reV0x7SDGHjlNMQzARVikKmBLSE2dI2+pbkQCKIcpquAmhj
jTjIFybcoKk9/6XMdHgXsV53qnmGdcHB9gORUAGiJBZdWRrZ1YcRHt1A9XZI
Fk07Kg+ztchhpL2leRw0mPLOJh96HLCqPSdhJiFzdVOKOExn9iL7aA98i+O0
oWtzZvPe8fLNVWxoVX5DlRVC9H/sJjcDM1hVMN3izyN4iJ8UBEzvNbSlob1W
J+/bxtF0fO91mvPPVV8Dt9QCk9tgRJ94lJedT31s09cMwxyX8hZe5O4IxP+b
iqK8W5liod52mSzKAu1ksg7S5e0+BivvtIRa8hxO7yR0fF33DA3/0SYICWeL
6kcSfd7tmgqhVH28joevSN1S3XqkhDSI6IJJPTxzZYW4By82s5VWHlYr2iyo
wGcYnUXAVwFpOwkKqWiZsaCE2KgNZKvJQgXKHkwNiVd1Kk5Tlz6iaBOGl3zn
gvjeZGpN9ToqsbVxdfnbIfrFjvxkfEPz0cDrM9fFDz2QX6ScJKjl5cl4fBSd
HGJ07E3BJRNPiwgKxs1/FFvsXcEq7cQFTfnsMbOCnVJ3SGaIqqvfbJhpvi52
WIlOSAE7F4xHVlIIE74kPkPreNOQn3OuVF4g3Adws1aXA0/F1xJtQm/1VJQ0
xoVJH5qowS3TTs8LkEhYg9WlcBkp0vVHqakK/qmw2LAlUmYeWeA9uqpuLqyZ
It5zyq5tPkKqW0jP35LBs4lJETEZXP9Gxh+QvqtnNvjMnz5Hte2ZJ8NgYsFA
Wr4PduNzWUU17IGSFsuNKclS8jjkVfyDZgSYYXruhDPFGRnoPct6ar9iL1vf
CcdKKGH6PUes573YWBw9jTf7CAcoNqV4xcpIsS1v1KwOGvFeA94NmrlbymLy
88v+1PQ1/siSxwWyTAgM44LfYlYKPz4bwd9HcMLYqcxqN2eYFs3RUzgHbjfB
I2sbR8Llc2Ogqul1t+Cr4ZO280/UFuR4EPa8TQI0XRuW1nXUnpmLzVt50EMY
CD3iDlAnYfQ2ynh8SZc0QhMr3zDVbycjHoCJZIuxrzslLofNWSO57riF01qh
dk2ODMZbqS8RoG6/CW1tcjwLrarMv1Hm5k5DGMKQt+61zQgzA9jM6S3Ndppv
f5BzexqTfaYwKMzYLLtrlkRXccDeInVy8Ug4VwRMsmKPUZI7Hn/dICMSWrOT
hQatqA+ddPn5y3UY5kqrGLlz1TtWy1o0uKuKSHwLePuRpahOGskoEYU7mh7V
0mraJw0WsBqRKbbExrvieqFu6/qmWjyQS1ewF88OPJqUXPdcMGj8usTAMOfy
fqlRwFw7OEK5yAaad+R2iTEy/KipUP1jVJL+jY+BTj2AJ1/+O2n7qE7vziZT
V1YkvYFvPkDghh0zyrox/iipE6wBGN5t7M6GeQDAJ1lkd/54fQFbMVofeF/L
V0oSn2llC4Ijc+9F8Z6vGpuyOvDVM2nZHawbWmRi+I/r77MZRaLKs2xaElDF
k2fVvIH/p1RujhF/RWeTgSQqrVFtEhqIM1T7wWSOI8H0t/b8QyhWtLHaXImz
2aS/STrR7UbKX0Q5n+wj8rH0D4FObod7dtCErHAK7XnY9Nc1MEU9NNCGSWva
OXhpHTgF8vJbK0x44xXBg0FzJwmpMRS36NhMHzpOazkaZ+cJEVVuXjJE8Scj
DkqMw8Z7+N4wnal9Jw0ypxWnDon44/g7hZFmFwVizmYADPjf/TpTcN+VDyf1
B18R0dCsuNWt5Zj4shahYzHjKoRIaEYTopK/4Ic69EcuzV018JmZnNFLNw0m
uOvV3svvBwIUvHTpx8WJ3Xe8aQXCT8V4ZIOgmFZRpvW+r0bq0v8RkI2aPcdR
O33C3r9DgZ/R06RouKocE7f75eZ5GgaZGoJgwZEjKV1QZH/zFRXbkkSY8ecr
aJ+ONG0LXXXonp7CIYFwxKwGwvKZp1u56cWKu53zKEDEGD6E26kNiWSo5lV7
n8KskiBrtlxYaE+WzvOHCIWUV7TZAKgCK5xdIv183eFA47PMrykcmq1/wxse
5IgIe21W2UfgSN+YJ5Q9m5u0XTTLaAtnlTbZnkgs/I/Ra+lataameRSWyOcH
VrcZsM/hu84PJhx2c+D3WP+2ElAqNYWctx+WSPrb5YA6SKCrKOQ+zyx57X4r
tJgrpTQZl+hP2RgUblhVmGE6VAEuwRFAPkzQwN/eIrK/mMGC2hYRyX+JdtLA
eaM2c4+fQMacBLUvnWAGyn8+7Pg77CdnsSJ4/AHXw8IE9u6TYPODlIheJmf8
wbgaJYx+K+dqCPMkIZU9ibKJH+U0amu7nexDib/Gr+71qWj+SFKD624AlnRU
mHOO6JtzR5cly2xOzOasHDMoX+TbsTG8+j+GcRwGnYl6InJCn61Tu0JKkQWB
FWKeT9mIEyhfTXagQ4eAQl8mSzJ+vuaB1j8DiMY3bX5wxwOAV0QVh6gwJc7t
S7J+U+emmWK72lSFK5StFQOp4+YPGGSFFbG9w5N7TIFvDk1GomJEmqohriGy
dZ4iiB8+DeU0Dj8rtRVhtxm9hm+WsEG1oJV1sdHHB2R6oMW3j7TX87XI81dJ
czADXH6MlfIAF8gIkpokwnjfhZkSn5JlbBKlcZ0DDYBHR0yj4mXrVpGqzCEo
4FC3e8mIN4bXQGcno6XQNPINYhTdpQ3IxOHEuIqzyrb9hKg1rQOFc6XJ6/qV
v0DhSAPpTsytIstUR989L7izr3bG3heJHmc7Fo4K348o6FP3KMuiGbW9ar15
5URFn/CvO2iA2r3yQRW9R+HecSXkMwJORlvnmCLtMPE6IAPUGQHcLpanZC9b
aNWetRGOkZenQjDGQDk01TyrWoSbMg6wAecpPbys9lxhDNrH2l9++mgtD1U8
UBwitJt15D8+Kj8rh1ntoWqXU4KtZbY1xNa5QRqEQ3wYRQoIzPOYCm+EOLae
mPy09UF5G+uitSZ12R2e7jT36vu8U2ExOcTVUepZBzodPfA9QVTFnlLuOFPr
EkASThbWlHtAobF5EJ2P/HpJOTsiG47jjDGiknJqm/obN+4YINAGNH3vpU8T
8X/1wXzmGjN/Lxpr1qrF026+wpltMpwlU4Wn0PNVzJfKy9mDzNhC9TBWn7+z
1TGOcIPkn0uWZeTXwDSMm9Ci1OVE3XRKpZFsrnUZDAVDP60ndDDx4TSWc8Be
nd3Zx1xEwpfykB5gelSDbwSGUrrt281Jl1l0nU6q9hJO7JH54+6R+82MaKPg
5b5mrTA5opdA1oOJwn1SLjCGHyy3l0ocRdl5bo0/C/VWZM+PkSUWQ/8q1cp9
j+NwXu9cpN82fGgSBoDdbZWXCm3PWxgimt88AghBrWT9VfvTPf/Wl1PFzYm1
krhZNbwCu3QbOxo4HHPUMHLgNK5+1Ylgc89Nr14TXsbCsZDMR8Cv3ojlyRne
8Zc9Gej0MIQxlsIrgMzeW32JmpV5juRruXArLkQUf4KMDaUh3+GSzJM+88BZ
23BO2i1rAn0BYUogEDIt+lNF2QCQhXss9/1mVw5Xr0hNRvNnpMZP0JHprh4O
i8x0+zw9xxliQArR8bV/cDA3cCFdf4VtEOJDmDzFxZ2ZUk7wCrPrHJyMG8J/
y8JTUpamHbcyJsb2pEXQv1yBFnIpMKI88ArnXAGCpKvTdfFoG/8P/aAJuHu3
EGoBaBoY0AsizokvCSuCZofdcH699oC9d4Z36bWnyvrQQer6hDcVfLWEdwyZ
jPSGS3hN0C04TnHQcqEfU5kpquETOXqr7m521mb1YGjYrrl7cK/kSvnVqh1z
a05VqNP/U/S95lF8fcL5WHFJHxT1zuBpVFvvd6/drjy+kYmIAnxia0iQcCAq
OkmxvQXylthaUB2BxqUAQodgSc9TuL4nTNMIkZ3RKKBE6U+4aSEqiiTZc+rB
i1uJ7D5kdZlfSVJHHBSLT+fGWK6wcVwGZXovqXrzwzw+H5Xo4e6BRu7C0mjf
JW80uVMjDGeAjUVc6PRgK9NwQSYCSDxvcFkaSGEBc+hVl8z+VqAOs21+Ay7u
nUGxcL/C2Mp3QJ7O0y48KIwnZplHkEktlrd80l7vU4Du2jhD/9ooGrt3pGjv
6z0G70SMPoLQu3sBErCuDcH2PKHbmLqxqGyGLjE8HxzBHKVB8wDGTBnGDF7z
48AiVhkOfMpV6YtDfpxJ6d9rKyA1Bkqbr/k2bY2gqP6omu8TFD7wtOqc8Lvo
rJ62fdB/CwFCT13Hz6f3KsRkl4xtalVbxHz+9nU2iTk/doSrdojNW28TDCzd
rKX0dXDsATcL4iSleTVDYzsH8YvBK+Z+rRdOPnG+rZqewQ4D3YCwxsPpDj/m
Wbc/iRYtmsiEvMSgW3GHpMPmTmCEXQ9hfDJW67+gaiP7/4t7M7dWl3STPodM
Vk87Y9gZV+fpdLRvaEAyftlF4yXRyq7bMgkaLioOCQesYRuRlHib6AOTG2Ns
Q7ehkAme0gw0QRhhO4BiqJaWAe/M8oeO5gyOUcyktfLpCBUiMy6EgBETkrw3
vEuYBBLW07BUoqt7tHbZsFJs+WoaNKpgxYr7Af0qeEvf4yoqtXiUbOljPiBD
TplwyDwY9O7uDd05TcTWhH0Nd5ayHE3NsBtkM3zGLu6z+a2KbyZtc2FgRzou
LKPGm9dqjSmgEys6yo52JOZxKIorQ27RxQglPL6h47BdheV2y6+709TSafgr
yZbFNUNs5hdnj/Vvww1syshIhNnxXN1I1ym5YwtabYUfMTfggguY6EaiyHNt
T4sOGtkOHpwfzQARMKx3GrA9+WL9mjJWywxoPgufl7SBY3WozT3CcdH1Jzbk
hCIzkm90IKwrTxhDCr8CNhd9vJmi+cf97ZPnoSxBNIdZeJty/jouB1T/HCT/
Q2w32Qc4rH5ciDl4VTwX6iILrJj1dseqMaVGvs5X+bGNO4GjbpqOCUveLSfq
VxtbPSgwgpft2UNjoZId3cKHZ/jhYteSLMcK2RimUqVcMOqzGZgXfFMulBzy
PmkhyY5FvsXEZOAA0MjF6BE44EsqAssoRMqkEySqk5j9Oexrr2EK1J8yKwun
vobphXkjlSFWhVUEoauFkF5nvTjBOi1+s+pOHlt6Cvy9O9b9LY62S4IU6RWo
2tE/0fBkOZhlpjMiYjjCL5s1ZBJDB4IFx5v3nueYUEzelmphb7iy00D9YfoM
lMkTqWZxq/H8R1vPreIP27dz0bkrayHPypHBso0/isN6iQqKzm74bnaCJ8B0
pL3TH4x2OxcIa26a2pdL1+RUWiV786udBe+G88o8aXDPg60LEoT8JcB3PNpM
hYR8oexAl89YodjDAsA6+sWTlvB5rjv9g/TjtNUZxO7hLWcVoNl8LfwY5gWz
lrUdqRqEHmz9zkvtxeXDh+3uGqVV4YjvgJ9GcA8iVL80T0z8iZkX+W679d5i
J4CXd1kiCLG/9GI+ZRPBXjuPFzxkz82xTLVtplcEUHYD/0GkTTcSRD4fjoZu
oeidFtLTuLMwnh5s+4JIHySGUiM2a3OCzndrfdQqfYifyw/uXvZFIsZNiM5X
oiGVbyQG4kY1Dnh0+4+kLWFDOjbbC8Fup8xSxGdVs80/3+taP65YnyGYNIln
b8Tvzr4bDSUzaODjEUwKpvgqRzrCMdr3HCBvYjlM3D4P6h0a2uf1NON0KULR
NpukvLgY9JdxYR6GN3Qn8EEDnhIUB3vci1TR5LEXgAltwDOsa+DFz4q8jllU
FSgRyiHf8XOApayjGde7k+dRzCKvBh7Yyhk3OxtjmDGf5U7KP+qbqce17xAE
2xsl7juX8f8KpUTETuN2Y5tHkDLVP5t+SR64bjcEsHZRJ2l4YhL1UzKic12n
8KyPHyudHVl7scfrgzA5sFX/1LnUk126Wwg4WnzOk2nwsIdA+u01FP1cwr/3
VunesJQpHV15YzZiW55tCAoPmi5I8TjhHvBou4MpdHzrXLyW1S66XxIzQvc9
I5zvdu709xtR/tu9iNcqGFm3DksfGnkZOw2pYmS36cTB95+J3moMdX9rTSrD
5Cs7+IJDcac/n6iKsEIEdt8JsAd7D4243eWAVdY9R+JsPp+AfgQ7QDaOkH93
VaLmgY7Kr3z4SxQSXNxHUX/DFnLk/D4fSjLPK+eERNBaO4hM88T6UeTaOEfU
B0STYzW36dSm57UJLiR3Sma+ahEZEK52mWhMNNsc3GRdnxZtfIrG2i8tjaNS
pH7lCelxTDlfivEZIRAYH32MMBY96bqNsIi+gx0CBnZhwZatevlbq5rLovnc
kUbVRdkxouHMJM05MKqz6Tv03pVU2Yujog5/b4Fu/hACtKaBBYIjQkbQFtbo
57ekuUVgCjl+RkkfIx5E6LnaIJFG840Je0A9PGfMuEzVuVU3oe4a5bPA8GWB
L/A7Jrdp3Nqn15AncZfzTjTTUfK8soulxnFKxV2xI/2XOsxRwmlQdETFMbnm
PRVihqHPfIYWIFaS7sGvrBxiAKDAhbhGgV3txi0ZvIjSwILnLz1oq/cAQYXN
Sdq/h+zd3Eaxdv4zFRbyCAQXBukt/0334yWu6CYbqtXYVWdSplnSIlHxO4r2
F4o+Bsoba8sT1QUUgKhYAV8UDKu/xzIw07V6p4jykv4gaLIPXk8fVXhV4LDS
aua/4c63PjEc00UG+bawUrrVRXAPzIZbmBCwcsGzaxxEVJJ9OSQEF2hfN26w
gtNrp+JvkL8HkgpgbtZuN5md9lZ8hZUW0IJcgfCcFO9fJCzSSmTudQSgUvVe
z2DPPwFCSwyA9lY5PWCoOfaBaefeWZnZ1/Ybgg9/jjChBhZlVmR2Ri/A8In/
Dkv+ji/r9K86zU225HC+Dj2gjHhkS4FNntf2m/T0r5hDcTK+iL+CXJimSC8Y
MbMoi93UQ4CQyOj8x/ulTRjRuKr8tlwoXhxMFr+92u5+SgWcKUEm3DyM3T73
e8s2+vZ4FfkSa/b8wP5Xh1zpcsIGaRVze3obAuKmBBWrdI0wXzcgzalPisvS
yZshpA7y9ce2nS2SUjB+UIHfyT1LJLgmC+Jlli6/O+3qn3k34NPHsoqLu6B0
aBYHheaBMNNXkjAIU8BqIhytYG4Yr3/dsS19dvIVcGCfDzE6qrLNFZtkGxhr
7IJ0DPUR7GCRUmt3kQXdMI2Kwo3QEart4mV6jGdLriCW2lawwlqG8W9O9hB6
xKtduUm9OLIgLgnuXAQjLEIb9ejaqaHNIBzB3Vkqt9sI+jcB1j9OjnVclLtP
qM4nm8DBv6JPahiLEQGcwLvqrCUN9R08gavjZzL89hCxKR6G+ORxVbxS1T+D
qXWV2Vwp17jQanoRBGWlkU5OMVpFIAhYxHfjytVQT1fn9zbcUg9XKRCz9Zs1
f4f4Upxu6U6tbfuBWqJdjeAzmJcKlIK5EtsnSTV3vK2cNCwyR05Rn3AuTgN3
spQOc0MkWwrtGCoJW2hn7rFOIUTYWyfAZbXqZPaMBiY8sLIIJmNiNLmZSBK+
A+0vLXuOkwpDnNprv0YMzEQrQ37EjIVshNnYIgzVAOvN/2CmjCuyfrswFx90
rUNJe34pXQKJ9EKF+Qls97G3IIOpI5wlm7iJCqYk4XSefIqvbh4R9XkcYRRC
YqfIKwBjzncdYhtV6p1ZBRT97vGaoacPyEZePwaHamh20UsWHJjMowBJkRz8
1H+aBB8eX0K2YPLh9lbr9zsQngajo9vE6M1OXJOv3Tl8mRTYnljmnGN1fg+A
VPGwEW4iQTN3/mooLg/9cva6Ds+v/EJ8ggm1sEFl5kH8iD3plLoQYAdSRMII
rMOcedS55LMzD1DFXyiGQqA8FQL8tBXXZDSJicar1YY+VfAkqHYz3QLno7hB
Jin9rp8DVrbUmXoEwLvG0cTRwmoO35Eew6SUQPU5fXC63T53oDW3pGYGmuxw
uNlKYY+ZwffgBA1k3qPXmMetorB6YbzpXievJG3yzzKAzguH1i+zpYB2PxCB
opoF4pOg0CP2XfBktIpcLer0eL3FjN9o6R1NObyURy4WiLAu3A19KZtKTeT5
jmaH6CN/mTmCJkmDQWA/O1z5ufXCPvQ8IUcT77F58DH8g9Ul+nGmaAv/DHyU
cTyL06YjbIvDyyR/9MZE2BoUG+L3ENKF6gGl8AuYLEhUlZm5F4WDPqGPRuqm
laiKiR9JgzULlNpq2foRteeZJPA2rSvfxJ70lgu5OSat674FgX6el7T7guZm
I8GGNG9X73g/jSXz9gKdx0H93cHYWUFR7O1WVZlk2a+GnjS95H4sBL2jWBl7
yGvKyUMzXMS2Zp54gCcXGyBsmTmiED80cntd+2fIC22WwmZzL6Q5L1UtwlKi
2GtFeGbvVUhN3hk7VNHkTY38k/jFYG9LOaKZ1t9xnJTGgLEp7kVubAWK6Osr
7L75rH3NXGwDO9KQYkN6zq5skEZgCalvyrTEEbIxffBJ+ddBPDCKzzang/sh
JSy72EAFSbWGWy09OGYJXkkvBK5r1PgpECyUP70rFodbsdITvjtFNTwQTM0g
iO031aR1xv/lcBC8HjkAL1t2GS/2dJ07BnwGY99JPCv+VdIt8sh6cVYkTveY
hS9/9kIw/yj8x7dhhiuoZNgt6s87zZLr7mMP3dbZQNhmMhYe8XpEHzL70zZ+
Fv2OKNl4qJ1JzovW53BEBGFn/9jdqZj0BrT9mV9w7q88gDJHTRk5hu/OGQ6S
NEh8yLVkadoCXmc6ttRAZEVCedaHmhGdfR4+xcXLEfvj4DlOIn1jwtJeIEZD
rrRjh+ior1gHomEQ+K1YvJ/Y8iGcIxtq/2Mfj1yenszi2WSey5+t1BGVFzox
lCyEMoHdb2QnxW0Q64jhdF/KEqmHwZ8/cBzY08Onkm7ZL+F4E7QktDzV1GxT
UNluKSVgHDmO82yql5UUvnMOz9Y483sVTDe5Dm8doz22jpT9zDT5wBjBF/cU
i9qk/96b4L8woo97z9QVPqirgtutk2Mp0JZN7f8r/8O0bdVoeWppUZPj5ZyU
XmqYiEfJWwLclZlhigfXi2OJ1NNdBNG03JXlU8BVm0fu+mzuGQPK50H+vIr8
5t+D0G1vLgFlqwrH9zFH+Cs+TJNDV4n2Rk5/x0lFGloBr0tAYU6ENV0lvSXE
jEV8f1UkzqxYlJEQVUaIZONqiibbJlabs5Nice0pbEtg7nmWV9T0huZDUtAX
q3E8JJek42iZu6mVeCTXsrlskn0XDYbGsnF/MEQivrAFg7TJ5H8DNd1FpUsy
8Qd+98QoYZtSAXkivhu6cVzLNWimhWtLc8s6bhiPr1QCiIkoGi8aBcz1OqGT
7iM6ne/te2EtXEeB1HtDBjrkaXjlOnvpmYPNlvYmnkjJn01rLCDM8qn9pbJd
J9gmB925xhRt81yXwGYNXBqfbwSkVQt5NiCip3382lz9OlTysnJbreKkO0ma
uL5CJJUETYBV+opuqaJejO/XvfnavOLD2ICeK8dDDC2Q88uIZAfMr0aoGEve
G1cw5NR+mmgaSf94zyI1j5e3Wfz7ZyFa3rKO8NoX1azUPObAzSIZ8+6+n1WZ
ajZerBgjh9oT3Vm5wYHToyLFL36EUQ5mG2K4o9wxmPnQ5aZxavsbxsfGhpa+
JUvvFlDcfI9uko8O4ucqkZT68TLosVuHv0PEyBkseRt0BCx1Oy4bDa/u0E99
oxT1dM8qtbm+f4W8xDKli+LaYAdsZmWe5+aJhX9++ZivYBXxZ/e3A42mW/nn
Fbb0cpGqPOl/yE60V0iPQCnVNF9BRdrl2a0p37p3MojbbUUduOxqEGv/NhQE
0G52IXMnNjW+KyoRMLuJXhJPoyxhcdzzM+VQB4j8P+pXcMnoFTvFlpKReuIP
2wAgKP3e3YuBIcB8ynoeamhvO1Q7DvtOOKJrWcLUZiSoBkLF+m/HTgQWO2uj
usWo7/As7IKgqIT9cV+eO5SkjOg7YIwBDlMbRLhZTZI4V3nRkaJXnDUHh+8G
obbTNMUGItMsqtJhwHRMjN0wnYe4eW6Bo1Leajnb8+j92/YhFZhDhxn9W2I4
dZbKnlokROrw+rNkClgbGji8lD5bnNsBELjHFcDmJcK84/2GECdnJTLMLIo6
VHCLEbdPQ/vKLZSYMB9R8u7+xLbqQcDoH4Yh4pNaIioH2dkpGJUFSrw8YdXy
qTSgq64Aux1tx8DE4WSrJ3d+5koyBT09IcFxbfLmRUHIY0ufyEp+Dk2UveJs
DN3lF/DplrR8SQbWHDH9zsjNsFNC98uEjbLwv7hmuWz2nZ/3s42q7FfIWRTC
xk7/7lLYp5zdBPpE12wrgBoxcLtIopegR5NselquRSjHKONhscLztCuPI6y6
l54Ur4R4d2cGKyFZZmokiwQ0ycY9G+KoUXZHRQki3GKXdjr9rJwDu7KFuOsS
6IHm0dNMl/h0FpiZIxJfHq2ALmhkiDLKgfiRnjfW0CxpEqiU8NkL44AO5TRd
qq1rV+wzrfdH/gniVHP68FvnumZEukaMHM3iVut++xn8IN6WdCv0C4flN6Jc
4vJcVCqm01DYedP/Q/+EW/JXsH3e+2dZGjmBf4perK4W9rEsBRY4kXPrwe/p
0XcfWB5QPDPb5RDpvcU/sI0YZ3URxDUp72es8xTFKV3XfqYai+Z7+E9TIsQ4
w9G2A0SXEbzscgqFqXgw9IT2Q9s9WKb4Cxf2ZPNg1PeLD7CvltGaf0aSfQyj
B9S/GThgqrSfkCWSzc7uvgCuv+hSf5Y8NwONE0GQCn/9JTDg8Puce4PqeG+1
3WgJ/9gLuYjHb+O6CHdxlLT6iGup0y89mBDzNl9+tqmFNGmzJ3LzMlVuiVaU
+eiWG+nqzt0NVRb93Jf9ZKxlwICwm+8ZXjv0vLABtYAFHtDNFf42Buvp2nM2
qBPaMGSFPxmgHfVxqyCvLSknZA/cbcMjGIM4L3p+EMlwrKy8U/nXWjj73yPq
oeG28rMiX/QZwZpxlcvZbxSObOYplCr+Z4mOD1cpBRT/+PmVnYD63hEEYcUd
LUMncMziDsunNhEDtDOqBZ+INuhdNDMJTEf63BGEsHfvPuvbZvWTMtQYhHYe
BGLin1PPSOk5C3TpUmwtAdXL9s+eUwQMCLcvLY/w3QBf4xgzCJfWJaptwB67
cGfs7v/VuALY+oZfAHDmS3tOPyjB8p79R50PPqDdOKfYs63RKaZ4PYySM2uO
8st++JATNY4rkOfrw0S0A9LnwYa2UJ5Y9UnXVXhwJsKExKxRfwIxi/x4we/o
YVWcbNTlSNb1aBuASkx3iXhAQIyQ8j3jNqeOWDtbCfm6tTSVnOt8QzX08Epl
o+AyZeSByfX+e2Nl7euh7wRu4StY4gpb6nKxN0CRzxM9jK/WcSD91ycXZOqd
6R4B2/Owrvzt1feGdkoF1ZaB3+Tf/wVGhLmLnNJpNms3lQCVj1/zSAy1VxVl
zPyC58PnY7odSCZUA3GzqPftCXVGhr/YLnzNIbObn0gSa3DVAq1oMQekMAcT
HvlXcqDXaNKp2AGAwCpI+8Y3TrTCxuEIWF3rpChEjz652ZwCQCeBlzrZw78Z
GZmsRxSXfsFgjds6LBxNIv6UDSFh4azPDUKtofT+WCTEMAwEX0Cr4TcfkfJE
ciVaXwvBbaH6uZ3KcmC8Ywlhn8zmMJ36pyroeiiWy2KpgiB0lDPTUKaDeXxe
TwROwaKb2YD9WCEChCu+HU+6ZNPBumQZudyW4fh72+E/allP2uLyJOXu9mLe
aLrUX9WLe46l22AuSfrqdAVbLgRPNRHyOVXtr+L/5mIkxDAsb8ogGhkviWsu
FU0jdLiYh1FJ0RtONnUbLU3HEn3xGQ2WzP7ScyXQoi85z8pCmPUgsp8875rl
Z3X2KqIFexczNkb+2J/5IEFJ+JbZITsTR+fe7ggTe5JDOxq2X96HCwgPELJC
yci4Ba2vh8UoGdCpJQ2AU3ywd8p/vOQXXU2WPhKUxFNYLhfjTxQD/chi8jFx
/preYnCtZUXrwbunEN9dn+Ym5lORTUM45kVgr9xudrV0WhSZWw2D3HebVX6n
4MZm51sLRPzGVJLWRp57tt+Dsp3t6aL5eWWEcexYo+U1UWlR3usK8cutbErc
bGZ+hSQqSyn8Q674pKsQy9nXs0yDnBIh4swmZDqF/nSDpO8ZqQyTU9ffUhwD
kYrp1Tt/qZsHYzrClXSgLLpvvxFlDahMW2foOvpstwb1XRll9kKwjpnk0DSK
Oyn9f21hC5Y9fOQJcaQfWVS8LswlXdQP2bReE+OmVQKVz7us/G/OCEMi3eTB
KR5TTbVmg6zukBltWTFaHef6owf+OORM1543YznTGAKD0AKXRGMbad7fnP6T
hbNATVidyxvFhdy+30fExQBinOe7P+iG26MtlOFR0/+pX7gDMxA0iYon5/eu
T0IrQWrgU4KUSzpQLAvOWvlnrhQYkoqAWIUeJETTgJIVBBAFNLg6v/BsEnIy
hlFc8zaVnBCzoWJyEhXATmOUnZngi39pvZmneWzNV30s1cwq+9kJkelS2atQ
5Q9rE1PVgy6bjUt48IfWNOegt6a1CS+7a5Kk3W5Zeljcy332cIWnzTHBUabn
eECiRxgN2aPia11l00+LN/19jR3nk85NmBuSb0gwbdJ83L9t6nPHXVWj3npg
Dq0ywV2hDlFBmfa+DlIJkrG9XfFrukLJ9PCJ68via4Voqft/shUVkM1SBqse
mCwZXlvorahuNDqccglOMNNkhoMxYgQrufDEUMyfajcu/mh2UzjheUHQT9Ff
gdbKwSKMmWgm2I6eUVoN8sTP8FRfa/2g17rX4E2Tkz1SB2dwnJcFNp+ApAe0
wwE+mrsY+MMHPe252NGg0V8T2Cpv8tPiFR/83yyyQcFJii7GqiW6j3eLRbpQ
14x5pg0G86g9QbNLU45FZbakSEmRBGEl10LRGh8Dfukcia9oDFhDCpYfm2Tc
ZpYkZGRLcngwjc+Ep0IkLN27/A35ctf4sRFkfK04MVUymmnNBY3I6Ux6Rmyb
/3z56F1ouS+b/t/F1XbM0r7+1yk7TNAfPVNbFvZqccxDAZ3yZisJX/VJcisg
Yu4vkiNyQrgKYQh423AqELHxkhuO3sgWXPw1L1qlKQjVJHqIbX8q4YRNU1v7
IOOYIEGOW+/GVt5XASycVOfujoCdiMrK8RhU4BTu8uyB2sGzoSV7UpZrg9YD
8sTEDefUX5Z6WWVd0SxaPQgrUcqtBFk0989ETAVTYB3iLfwAsIWNbUD4ltnT
vfi+hpX+NinEuz15aBU2u7yDyohiABANGM/m6/wAfQOp0AZdPq7vGa3FWBjd
5NhWvCAVeFzVcNMxnMO5MYUk5/S/ARDRdp3ddL9zCeoqwCiIiEJENlKVdRFJ
/DykdacguS62+uwltMMHdTe4pXp+4zqD/X0o8tJyGTLmHQHFHHc9c8fJ3Ik1
SjXTmwVStaxlBVJ9otpWxPhjAYaUWF7XOl5q1akv92GGf4dqgC4sB6HDXV9N
IJpW/HHysddgP0o9n+BcbhfrWKJU56jcjsMsaNF6OQorFvdCyGU8/2RHCH3v
KEi+Lj7xhmeALYo8bKsxTZSBZMCLfPVhlHDrafb2VJj/bN7zpXb4Xa7WEMtT
GjrkROm3V+HL8YFSNun7wIasR/O/csm1emPFZPHXUF9rNrYuaJqXlhrkCJk1
UzoDMwi9p0CYKWXIgvZJqz+ULwSUO9vXAh6OzeB0doXn5ApSWYICZI7CtZ7R
KTWihz9oBrAlGNFGmodVOiu1p9irl9Gh+dKcssksJ+I2SlYiSMgpi2zlzV19
iuPGmq8UaveUWbQmCc7jzpF6HnlPZdRm7T+31wG78+6oclzZbesoTi/AT24c
keGpKffithsIMmikGzRBWDzgN3f05fYNU+d+955xtc333ep89V/vb6kjjToR
AnjR4mBaTmCsvXrKntrGXACHVvmDFYuZoQNpaislfA+krbrZm8fvEWZo2M6v
heYkTxafrzhZDm6JAzrZuMRygTn4d69DgPW3YuKM6a3oRyQDk+c1HQfNMjtw
5kEqUeY4z7wb2kvC05mGE7CJx6xU3R6lLZuERxdCDf+NfZKQ+mZxqDaQ4o53
0sJHbHr0SECtxqSG4SRPkL3XHnKgupbd6LVlQXUhx7Z/+GaJkDYnmssGYI+P
dGamjMfob61ugp/F9EvfuNMjD5Cf11d9ohP8upSBN+IIqPpYlU4iXDITjBOp
yaeyeZzA0FMmsT2XMrOXfqueH96o2LtUDjQ9YmZ8uY+Lhk/Lk/rDOPCW017/
IepQuNLb2C2eegaGhO2Srw0ulQ5e6eXtUuZjxRraXIq1s/+IVEIkjHjPFXTu
8xLbDX3A3ptQq8D7d1zkdtJ+VpVAp//zOdKVhjm+KApoDGpIAUczbGIyUNe8
4ewxWQHS3e2sb6GerGJtUfRBU4ACXH5upR0u9/f+mQALp5r4KGNIpRK2uLpR
SCiuiS5S0nGIFk5Zp+NEKPHtORVDEfTCcSJg9FEsJVpVUn2e7n/6tmN8U0RV
I7zott8MF5ZaJd7FhxvEIrYTd+tuWxhBqe+N3NgKEkM9UmCMjd8cm6pGFZ05
0jtJkPdXp8rFsqLQ3dIIchdWBOje7pJQLJd4H8+SnqwGH5TNRAtYR7UPz1nq
k2fX23L07/MqPPth2nb9J1H3wepC5FgAuPi6hoW6kEATL1Fm58G+ilMcwRrH
Tc2WQzB5HGE4Gx1DDDpuhKEDwYv9uxL7c45tGJiLM3l5KqJM30vKRMoUjHb1
u3TmQzOvM8xVBFPf9nnx9ufbLRV5FSyGMzhUKg339CcNC05gO+muqbCHIbNJ
LUisHBeu6s7sfSX+EB2oqV4RinGyToQ7gZ4K7gTeJiQw5ytby/OuHFO8R3wu
qOieiGJt/cIhKPTex5QluaWw3mq8Iy9gQxCzt+mQV+V6ulBxmBdjeTjR2sDM
0/Pkwv3cTEiY32K5MbmtmHzvFN1lHu1zVUhxfSgDo/8zxwZVyp5lU83Lsbt4
QNrJkPMy5+zm1YAczVzKlQCmbi0dAIax8+wfriPxKmkeEbj/cL8+Zhh1pPbW
29rWZBnDR1c/8S6AEoyF9ovJ46GdUIcYNYHcuDHLYQtnYHsP+UKAhn7aESD0
AEe4QKdktt6gRxJqu5OUxwaucSr+Y7WA0S/x43ZmcCKRftfIaSnTYalOd2xX
A6adUssd+sgDPQRHnLUI2Oc5fr+Pw7V3Z4xSoHDBugEng/geRUSqfEQ8+9Yf
7bTrsZH8/97CNvGS+vLQwijcR9Hu+5/p8xawzDHZP8WAbzl0l3QjI8YlzErM
z7QzmzLc7IM76uTkFmhpPLo9h+bwTvowmUUmeJ4WYoVLoc28FnHfNXFx6uog
0PSpQlnNShuZzHnFigL/7VhxzX81QqFE1taf48IEoS0CKHAWWFJYw7y9u/XO
RI65sMq0Au2zelcaanE99alGJ39goMWam1sy+RRAa+oc4zU2YYFAE4kzkssd
tCLW4miFX5VuHu++IsaNdoWJDiIYnZoEqb1UlLtPsh4stPgTcrN4r7FC4G+8
NukYGf2gJKE6IdwJrG0Cp/jCLJq0RbzXqzwLL1LPVwW/jSp01B70szW63VtR
Y2lcYpbFfH1A/AbyesBa6cY5FHRbQdCEIGvrlDRAZ3jLmhJ1/PQslJNCeZrq
TueROWEXSS/b52DRhkHduTPqKZbs3JLN3O0/KtIaNobDXzd0Oj13oTVcrcRO
6oEZbwJbs/KBPcZZE+0jCW7a8adLDU94D3t4uezwUxeI9aTT3cRVPHxDNuiK
XVGuWeWOP+Hed5jPnzlWIhoSBv5x3NmJlOh/0iVrl/68eem8Wu3nVrUNNE+Q
gJQvRtZv/ZsAbIEzNtYqUAlIUJFRJsLmc3MydPnRQfIzcw33Gung3zYwQcu/
uNoZAR7HNjNY2gb9wFVZ5cBSVVo2qcKivRdJJX/5HOildWJqd5h7UxqsX0LV
U4ibFu1JzLr0g9rsVvHv0S4WMMS/EYH2n9ZoyeLB8aHyvlWxYEjGn5jxT9tq
a2UWU1JS+Id0/v0fL9jzPfb4tKPgj+iWVv0tvVun1iIRQPH3+Ltpy8gsnhPj
56bdTn8TGYIfBZkcTlJMjdNR2fQ4dcAjDT17TBLQVEQhYPGpHKD6m7ChNIsH
S8A7cQnWwnOEgHorrb/ImIV155mNC38t6c8uY4ZvMNFJdnU1uqfu1S7XoEMk
P3xUhvqH1UEvVqLMd0P7kdJGo3QRJCJWmWmXuubCx6wEbiiLIuKLC8JfHOQs
M8Xjqrmaq0QSSGL3K1Cw4xezm8cerCDo/GMqx4hLwT1ENt1aS/uRbS/Esqvc
LYLAw3uh3LEZnvap4UmlYay6JELRMIH/Udov4SPrHoSZR8C4bpNTgxcczmkr
cp8NRJ2aQTMlkmPQQ92+BFPwaQADY4rpBviE4vtG79Yl8FFtaydOYjBpSnGI
4akhJ5XAUjVpYBXlwiYBBvtfbY6aj7sHqXDIJcsAKhx9V329oQU2xmyplm4G
yg3U48E0ijYqagxJaErH1ApC8YUys+RcOVef9vL3WQALx8uh6ZacGFzakpIi
XdOMXKBbygFeaNYGXrkXdbfWQBBf+7qcp13bL358QBy9kJRT8f+FKwOCL3eZ
dX+Kx7cSHVO3TNEy73c1f5QE/NzTLlIID1yNQ7YekZEWf5RODwqHrPXzzfAU
IOkXGYpecStzXfx5Rm5x8FTZcoIzFRWCfNYq6z3rUR8HVB77jzJKp7Zpgtbk
7yJUBKKruOmj6WwNjUqY2KEEi089Zu+pO9zlbTOe95Oha/6mF7D+ONXGA7rz
zcPthw0J4N+aM4jKDghq58i/MaALqhB5oRlw5sq+jYG1XG2CcuXBjcl0kEl5
sjstASGSh04AEqPxSES9sxAVR9AW0vWqtj/SWQSakrDPJb5J7jFyAti6x058
dVhHOgGP43BI5yCuvr636j1ZDrOqYv/49OQ/ZhsybRO8PZDdokluNzN25cok
fLeILaS9iYrgdZjqZWm/4hPlMoyOwqc8TspN9/XCxJ3ZrFHpmD8osPvttMSL
CeHT4HxYf5fwJi05dqKPsfSizgAqFQdnzI8G+aDGfARrTfsoAvtF7AJ4uo2X
8z/LCyUIiWDmj9C86UsQlbD3PEHaV3f44QtY5fqViU4nlLtBFBd1tQJJsr1a
iLNxirkFqhGKAiuQTUkIVSE4eEgFhQrviBsMQtVqx2CiI1i5sqo0vOakxf+a
1BCNtXTnhh2sV8BwRN8QxsKdRu0SBndgssV3JS5NPGZsX1EWNob505zgwXjb
zB3Dz9xWvaur6cwqG2nzRYE69A6X7KqEAY2peR7NM1+SO36oeVrlH6eq+q1g
/Nx7RWkhKVT7+U+kcbnSXlfbHsCaIbCkkLZs/2++jkCBxcL1fxpO+3/FV2kj
KO+g4bE4Cjcwm59YlRBen116LsWfC+C570R3JWNeuBD2Ye6TtMFHHdZTgDUg
6oejH1TO9rhaZqArH+nLk+GHl+ZVtQ9icide8prg9v5m/6gNaE1scYwqyI9e
hnnslYEaM96O3F0aAu/2vapK1sJK5aDyNEor2vtXiq2ZUWHZjAcKPcMzqEhO
4KPMS4NdGm2fgVwoykENJkDMXzKpm/HfnVEicfrl3diPhyTQlFnDEuozLy0G
OkAeiagDBnsehoFCkBS0juhbjMT+ZcHHJ1dVQ/stKmRYtZYqlTECnocrUnAO
q2wkjt5fv1iSMQTiEB8PVEUOCAOjFikLLiyTbRMTgkQHDAR1w7mFlu4LBOvz
XtfzLecFerMTOswUZF7YvQ6Oxtsh4w22AeE5JGcDSwgu7tVBeMQxJo1MuSZo
DfIN8Niw0YSRV/sgwXvSunzUZKVLJ3JmTA9YSMIN6REtMRp2PrNPhcYlaMVB
gi6K+oWwb90JEC1RxqWNJPtBO4ARbt6HOPtEbe9NSvNCNnhEqRDpHYX82KIP
WRCNHqQyBZNvhzsFGcxI0ZLotPBj7XRaASTjWU+X5lritG/IERRIiu9hfuZP
TmJbBvSCU1hSvvlg7Zec6QLk3/IClcazEDYY10l+1dPLBvbTGcce3dnqoarH
USCB0nIbU7TKn7TBEJc1DO23Hvwb8NkxRWIvnCcyyXqA9aUhVT0KnxIhdGeE
4gJvrUcbU8AdHH9TM/OYNhjkbHNgKmvv14vUHZg/Ya3BqNss0tXX9GyuTvh+
bE9N1LkZLXp9shx46+Y2NBjhO1xpUCc5ks1rdEbBvrK3FCKwvofa7lFyLLHn
J3MC75dYAVs7ojvMccyH7YOJiDBSgA7370EmbVFNJMgFjSIQogQqhV7Ki/76
LvwsWoewJwp+AjAG6hG/DQFUpGY+eIkn0YiSEoEkhE3xwtVCYTzv1xtdHxyc
oPdhdTkWIrVnAAEFu9sQkuwfGqbAT2yF4o9tgZnntuMabNfIqwgA1qfVMn8a
2ue77F6Ge7rG+68BmWao4ZUZTprKyY0EW/9BJ4k0glM8qtcteK4WBXzuPe7r
D1QhwSMN1JKLGS9F21mG5vxbzCuZ6dcvGNkQ3KJB2wplSPmUjEeDYoAsxDvB
0OFjW4KB0XFXXQV50FOtee6qqPuCDNTwHc+yzKndKWNQ/v/hdT2U1vVUtZo+
4UY9S3lDAPspmFLKbngsC6tfmZDlzIcBmCFvWKPQwqBo65hNnAMns6R4ZUh2
dp9ECoVeQiKR8ud+U77waxiSJtk7WXrdHR0loXVB+U4Kfs5DwSbPd12SrycR
nbzmxMGwGrkG0qYL5e2vsmycrjJXy36ZG85dAV7RBfpRDErzQ4TrSz+127Ct
tXIIO3rswn/3WueihSHsratTIUV1otHVQXy3ZGphUcsM/Mw9MPOJDBTriXyj
H1cCc0fvEO8JAcZ+NPqzhzrakijNNpzOi/vZvGypVbGh4fFiiyvKeEs7aolC
AsS1tA7GIrJKl+PKeTa2qZ/tSSkwJhSu8gPsOVfszrMdXRhbiewA4e+15Eg6
j401d1azmpd8kUrSCq/8tS3kw+PxVR+cb0xY9z2R+ZGQtf+XpDhppaj1B/0K
uhR2LeA6fGZEs783Mfq1Q1g19+VaIYR+xxBmWKA+Sm2IQt/63G/InN7EFZOY
HxjHmG0tLt9fSDQ/xc+VSIH/GnipNPtBmGFo6n/e5SQDHGRzpjoJwMtLI0PE
TIhX79SySs8OI0ibcVoAQMkYaD07+qoh+kLp6IWuNay5QMwR/Cf9QjrmF8mH
/sAlXfSFSeUNquRbiWziBro9zU5F7VtPkca40FFtQWTyqr6dH7r1ZF9a7L4b
deac+u4dzriFmlDmf79p8m6WDs5iCtTXszhbUkmAH46crVnpXxrAw0kXSo2U
6XvCJvcIEYQN1o/1N2CrN1EIxJOtcqytDvLrYjWERgUZ1zoCzzHu5r3xgYeH
u1JK+JNqrIw9oq4gn6R1xhSbDiWWQusI005389IYvew6mNS3n0+hHqnatuRx
tZWnLb39KWvRSy+Xfn7Kbztl8SheoZjGcMRcitGE5Mcq6KR969O2twgscJDR
81xw84D483dQ2P1/HdBB4vo+1x17zXib9Di9u7O+pYlL9MqQRR0WTCiNx2KG
UcHLQwv+UOLvl+85BpfUv+KM2WGWKIkZcM5VYi90XmfqN8rsVYIFIX049oUo
NV5JjjD5DLqAyERMQTH9p2bYhzkQ/RHLfy7c2Qjh03qt4OLcjh4Um2SZYLLY
uig6Zh4oau58jHT4Dqye/gDvsOkffC1x8xUOWqPiWxrc8POIZYfvvVhBQT6i
sIEyuNoO8cJgfHfUm8yqA5zpVfwk2Xxe8TIV8OnPBcfOOyqWTS7pjCLVEgUJ
2ISKlEkVuCgHbQWo77XI3lOg/6uY0/yxBqWpKmymo1QThHVycvZlThy3Ncwa
Fmy2OCO9o9Ip+U5kDf8KJCtebSiAZJmnHNsePXxZ11GXTTpU+wy6Nngwig04
FAwK3yjfpijLKVu8Om/PJKhhMyN8NUxbg03JYVHaudTeaJmnwPlTlQy7PQz0
Fj6xbUZTXCFjlTAo+d8w1AMH8lL8wX2ejaTfGaDc9kOYSGOdCTwdJnhBfu34
7Vj2Sb6B2JgoW0zdi03n/Fcf73F8cFB/ly7uUZHVc4j3ErLxF9cHo8DB3CoO
021MjJ41UYpHqgdESj7z1XPXObcwdcuPIydnSj4FZdRHJ+JTfbCfjI9tOoKy
ldN7bqlMQyifhA4gFBLwh7pwk7xMBF1T50QSExvOURxDWcGNFT4I5NaBHa9Q
1rGmtwjSGz8ecYkBCz5G4ie8+CghbF8JtgRoajRongcwUFUduOBgTZvwLeee
j5wMGJzPYCkxE0wCrRJNC5C3a/my/25JSFOIdIBo4PvtMOHhoL/lzxPjHDP5
ubrcRVdfdgEHJQyItXhCiHf7o9tcv4PzEmnFMsDGdPN/8I4tlNg9g8iGnCgJ
lvO/1HtrXIa5cvtW3stWfzqT/7X6CiBsfvVUY1/I+0EJ9Ce23nmn6m70AjkV
b4m2d0ydF4KGcvj276m17u81MdrNXL161re3aoVzffyGu4XfQnUPjqKMHLES
pfN79Kohhc6gIEKW4I1CPVYudctHkAZRSAfl5fFM3ap/rCB1FAShJSb7bvmP
ZtTDsdJ8yRTuR4gQoI2ok26u3fvWDekDbstxuQt4PsSl5rJExanRNcsbLO6j
CfYnq2VO0W2oh+PU/PLyXcf6t9y6+tDm/P7oBPH2L7nBFy6XPKx8KdYeJMxf
z7LmT2Zm+odDFRHh2+HcWm2UcRANW7WWMulpc2AvifhpuzeMmrDebPNlFvP4
ML9rd8Iq9Uluu3LRqb2zIDZTHCVm9XRkUfqTRG68P4CV1NvBcx1nXeBvRRFB
xY1sthpMiUzDXWrzu+iOBkFfXNlVgcH3himtqcZVJGwnE/Bvea13hQ60K9td
bHG2tzB+qqApUxH5I1faql+ZUV6Cv0ESack9XFDSwcoK7609av1Tpjx/4mDL
fz6ZfJ2fw3/2e3ZiSO56Ndb+4nnNVG+FVeFz7sqhJopVOBIGPqeno/vNhBKD
nITjbAR35o7oIynorJOGkLsH9AJurI2zw22magAxEEGZuMKcVWfn4O2s//j5
SfLRKdffM+qQStTGm1uBfcC5tgqvv7fZa7SyjVniElcESDBocwRAWEeD2IAh
0WabE0dpNmHhwqc9YtZrmslr361J4qLi6330Zvul3ZoD1HVGTj3lbbsqC5HF
rd11cvRgImOvMtbg01VPQp1o4RSaRa5vLSbTUZVh+G+qpkTTA9QRyVRsMqYl
QK+QVB9HsQKF9fgkdZYt/tGaWS6hKs6/vFcND0K88lRRkbUlmf3pZb2wjOW8
IUdKI6KlD5M5XfMGXsh3d8SVVFS5Ga4fszrMcQZjLKu4vBScRlSbLHIYz7/I
/ejgDcweiWnZxRLStoMRMGeOkXhrAf0p/tniNQrxiZjIuSLabELHeYBz/jkO
He++AlnFYJQWZW9rCUPHxQvqN/bXaQCmDzJF+GfYdBV0x+YhegLMHIT5tsXH
3e0D9vc5zBa/Y0zxVJfLX0co4gOmq4uIo9Jd83WZfEOWaK4MfiKcnp4B8mJJ
0GGzarnPAQmNYXbJBE92oMecqIF5tF0pVfcLhznKykQIQkCHfqTpEG8AYSXg
xwxXPEgSgK/uRqUy+5Gqnq+A1I6oHG1RCiaxhkszhpCpfQxJcQe41iJjKG1B
Nj9NW9is8pmxiH2FUGkENsfH65e4bCRwYrM0ioPY26PAfmm+ZrWhMveZt3ef
xSYeNqbQeWSuCc0AW+eOHClHZvvA+h9aGcX2fDuFVr6vLmpaE+BsM/KmD2nX
JQvNLygXC2G4kt5i8GaVQUP2i5qApGTJIG4zn2pPWJX+Q8vtcr4eiAmBMi7h
Dh5CoJwxA7jnSk1zpjX5sIy8Sq2sh5Kub00DsGcgcODA/wHmHl6FE1GkK2MR
dvnCuC1N11Zfu1HKIVxyZj3qmCTpADziQutHnKOMjBcrzZe6leBwoPImUXR1
jFd1inCeC7ndvHWJDHiKSODQ3oDTpUEjGMCI+JEBTQAcQPow7IEabcPBGIDm
ixJI5MzgJvPBIZXBsQSLQWrbJfC5q0Kw67xFtkRE95UsfPLzg20H+ZTCqp8P
ycNNh74ppwytdxEIH/A7zgKw4NIMuE8w9Z91eXR4eHal8ceC3Ya4H8v7T/CR
mD1zESPe5FyauHqUO5TPWaIAbqYhdl2O4R3tEggMVxP1xfcGO8r+SDOZc+hJ
dBeZB/BuvE8419JbqhQL7TgF6BeeBYzUHa/becw7Vw0Q2cqtn5Wa+XHjsYwh
f1n9P0qHZT5TdhLib2sdZAks2OO54Sp8tKgS8sJmwNZLuK2l1q6WbkH/yaI5
Mvvd0/zKqNGhDLOk+WtUjUZ7x9ic/pvUzYsRDXDMeWWk6ztSSSgHTQoD/Exe
qNs6gYTJE4MfzJaL4O4LPwZsFrVzi1KnEDUPybbp71zOiSYw7pNlMfqQ1W5V
Ca9iIQgxRuoeVhLh1QSZsL0upYfcgKE6JAMf8hGpwv+fIV7VDu/RGHQ7Cyvo
2dS30PCIEPs47qmUkB5oPEfvDdW/W7PwzIFjGWs8qdw2D9wDQIdkP2l3/N/R
AlMu4rvXc6+LrE77BrqCsiN7jX8UpxrKWu2Qh2wTk9VBHiwcGcBMBej8IRRs
37AwBAPGWhdlrYTghKDepmSlNwWLn4Iapcb3791Fbj33dqsz8WPSIGj6uf6S
HLioAebQbj6RzrTIWeR+q6J72iqKhLTa9Hyf3MND44Es4E7LlQf6QelVwRwS
xLJ1jFEmrKG5H1vFYMdQIFCdZPGXLdh+HrS5Qu/FPuQaPNFP4ZIMiEg8E0fG
N8bil82l/npgGsgqA2nrgwV1weQtVycDMKRV7oeYxl2JrkVw2CRkV1hppr3F
AILG49yKYXqgcpcyXU0iEVE+igr1s2QjIaXl5TWbifHhLSrgfdDMLDCUqoxo
REXyRy6iv29Cw1JNAzVfgbN0Hl23Q71lh4Rv2lYIZDc3dEKFiWfRXuH6sa0C
4W4nTqw/sumvKt7VAXJBjGhdAOLcRwpeKmtddnJ+mxSHDxMnArxjE9Gaz1oS
rgOTZDsL8FqYWj6+mFk+h5PebnaW7sZWIr2BlSfDhIr7Z61t+U+f86GZp5Gr
XdXKhpoXaGcI65Nfx3LYqXJNNzDoGjwm2DkBsehftcL+ETsVf7Q6Ther5m43
8C7cHlprpNsV38FKC2xWTXRXMq5nWObzuviEAb3iQCeayupi3oa+ZlAZ3Ifd
ZPLVO6Ovg/D2RJOSwvX4iMHOR2gdF/MVw2OErqSqy0tp/wdpqu2DssOYRrB7
k91WsVqDwq0vYTigz4XCqepTEEbB5YF2XqjwxeX2STjzyXeAa40BDQNeN2Rs
Qsqvl8kuO2hUFMaEI4o3ucoJbUAm0d/qxTpkYcUHS98sQCGqSW7pFjVOTFU4
RsExCir7FF2JVHA3wQHOu4Jk9BiqxGba+nwqhPq00cR5KcnYFrZZ0keaVR7z
g7yoGEAXWS8aag8wW5XXAmdBDKuZn0aKtSX9X6YtuYzuvXdDhRlRzOxFIUO+
lmuvi5ISboMqmKZpzzxKPZCNrdr/nzaKmUbxzcNYvc9wWNPqVB/sBATY06Ai
SAcJxrrRZRQ4mBs8XHaophyC2HbMbD98yQ7T7aGLFZfClGrPbun/ua73V0Fs
8sITXFhDHXCujBvcfKtd0Wgp8vZy0R+kTF8xgTDL526HDvZirnS7+t9PZTKI
AebXhCbxGTNBSJrE3Z2wE5UoGw4chu+235u7j6k/k8B9EGm7ufJhKTgigUmL
iMMIW4Q5MzTSjlYooX0Yx2A77+gaTfCbWmoPy8cftF2xGHLd3O1uP5SCMgXm
YNgwz3QKxh9Y25KjHK2SxT2QUxxNpow+M12jHN5QURp5R/w58kQhAL2DIsMJ
523e29wffhb01q1kNX2cMZKZDfB9VlZeIH6bzz+75hw5HUMGP+SYFpopF/ut
+boduTbW0nzALJIQTFdnlLLuQQ+TH88fgD0q/2KdyN74D+vRdwoGzFtMrdZ9
iYSj3pEOei5YaDN+QR+h9nCKw/ImLMIhsKp/27yWwv1roeB677YudIZJC1MY
wDGTwFWux2KNwXWc9qjk+ZYcROQayf5dApltu38xFL9xUz8aBfR2qtDykt5D
u9DQdtaEBOWg1LA9vqotUAnQ8nr+PTerF0ijethRLsZdBtKQZh11bgOew4IM
h+utt49z9oNWjTV1uxNexCz6EyDOu9lvhNCU9jNAmyCdfZdTeveEyGksL4rm
192G2649iaffKSK1AebFVfw5dAQZSUZWPoTXkAX3OfzqKwYwvnwQxKtswIL8
FfFD6kYSn9ONrNQNV9II/e5gQFzgqAPocNTx5HFPX4GJ+5yQyUaFgYI/bBl3
UpWe76a37g2PywdlVkK+y7CTBe3WQdDalu1AuCfzi04mr4JBHgpfOBLYteMp
NITWVBPjgB8Dexpe2qcXjeMQVaDfgzlXw6iU+aeUiSo4OvfKaSO39DEYYU+m
4yg07xGuxRrlq7jpaJGUNpYvZrFAITSLgujey8VCgeS9poMmFCQ+HLvZs9YJ
VBrsommBvd7ScrCcRE/Ao7Is5cuj3DAM0LeeY4WUNRbDtQ9/gkmboRdvz/iM
BmnsUQyq7iNI/qI1+pCEcZRoF4sWuA5+1dYF1EYTKIx5bLI1VWtG7tGOP4wU
7T/gKALqAH0fPaOZYCzNh1XVXRLNLLqIDjOtkk6VivgGxWzM0N56TeACBgsn
708occ557EHm9aTR2b5jMnAM9D2DlPenFn4sXStz9O2g/8UxqssmvgRxoqTE
Glyc8gPuwfFrT+LyYFiZn5GkJEqlXjKVEXGH2V8G0rpiqYPqFl7gkTeehlQX
QNcVULcA4IB+aEsJLoRLgM5ol6XpywrPIBLxmoeYEjQP7+nMni3MoJtg4/uW
PigK7jq+RjC2Ov3plHo/CFbvVdDxStEDRQ1cJ9UOpN0tq385zBwbcMLQukvq
7rifXhdP4MsgxZ5XTllRVoG2kcDc9AbhGALdkjh2PogIFmQkx9CogJOtHMdW
w7l8uSSjRgqc+IcBuNi/tuvNwNHK/K859/nI287qYJDSBF8J1mkLxBtVXKH5
+EfPzRVgXPaNKrNdi8mcnyi1nTYwLJtmt32Un4hCur54UJUzZxaPIhhBZWwA
AxUkfdFkFz7fvHD10YXd8xsCxE29Emx1vhfTGgnb720yATOLX/qyxuFJCjGb
A/rD3EH9OkPr9fnVppA5DYYhXei9bunxaE5egXWEc5CZSXCo6kDhnkdxe5pr
4dkSGWUuPe4c9YF2ZeBFXYXsxXjGxu0kKBzO/xYAKWcBvFDpoR9jMnGahE1I
JI7s6ek17f7NTaWKb/+5fjcb/UX6xewfixnezr/hAmXwJvz1vaHitrmnHzi2
8gMys6BzAtGZKf721tjMySbYSxBTExcuIi1WLYZEfxemeKJm0pSqUPa/6I+l
fYlpf4vrIV8vD0yOsSjPqdgiVYjFRiYA0QGX2Vg0tT8ElESAF6KduNv1IqEY
sZ+7mgZc6O9ZsQnLNNw0JPBWMOc4XQOzXLxgFChFf4AXiQExGhwy1miYZbwC
yRBzx95RBmYzKHI+bcbNjsvUihD6E+bZr9f5rfhHM+elpG+ez+2zXWQnq7Jn
iY/7Dl9UQZ5o48wfx7fjUP1PZdRJYADRbOekfi9uSQAk4x+PPdiRG+QeY4ZU
auINfaxBJjrKYwQl6t98JcLYJCAqZnq4jQ5q59HnZYIertRbX+EtzWeJX4lJ
kIeQ2e+RYEjnH78xBp201aafgeTNysj3VDsl7TPPGSw/dY8WapTq2FOpuxxu
zYptoFA8yWBmGQNpq/kmC4RPwj7vKDI4oHXqy2A8/ksCc3kVFbj2vGfGUbTi
PAE/Fwhb7y2FIe7NI9KXiiRM+B3j5VH8b/DySPYpzLt8CBwWZV/I+zV5J3Is
tfbgRBKnkk00ZuMzl1p+bHSTFAm9w3uqN/wcOnYEyI/ehcax3MMjx5C/V5M8
d6qAz8jm04w7DSV4gY+azzc8xB391DOfvzxHeFMLn6kOsnZHiSYkgEQw/wAa
CFcHyFd2GzwWkgi5ahSHkfeeWdAGuhiinBiw+hf1YZXTr106zEoMXz6aAzRt
mNsH47aVaFUvrya9Gt6zFncWsUTiFUnCje5mgyiwGloeT2dm3iE94rxEiTYL
bCmDp/tbUB9Jh4+VyAbi/XXBSRT2sEVSAUujvgzHUkR7oEwxc3zPpD9lskTU
D2T7x0d3MvoEEPEFHTAcARLmpUdP9HHF8m2aSBA4ONGz1LThfkjiIPkcokBd
CBVyM/NyHzjOZUiARYfC/a+B0DWz18lcjaK8VdOKnTV+uUW2A8edRlAn/Qhj
tljQI1YYMcw+S6iJA0caG3UTvxwRmAeld1P4hQc1ILs5c+8TPhxNDepMOs9s
vSnCQ+nJ+d0158PWx6MXWVHD4cff3aFKkT3+0z9lFMV5Xgjn8K97+Is08cVW
vnbuoRJCPcEjZnytBFpeyPGlwJefmxP1w4rLzg6BBaZy5iCsZxuxYGEbb2cg
JEi3QaUj6oPKrLyV0yT9MLGTipLr5K2tt4T8bYEFevamxYfEedRif6M6H7uU
l24mFf/Q7u/L1E1vkRR5EDtuypq2Pi/eCRFFS2lG4UQ7L+UyEUDlb45WoBce
fJThf0+zm4Edh80FlbmN5AmnNUgVvoaWqH0S2gcYV5ML0a3mGQ6JFfV8ld+I
i8PSaqFzAlxZ5xB0xnEjZYNsNzYNUtR52uNtNUfnv5T2u3axP1m/mi5bWL5x
bbOSfKV97Ou1RQyW1+Fb36O5MoHN+ZaQCUdKJiS6yDXP/+Sdq8RiT8HzQGNI
sr82LgEhee3HC2UB/+ZO7H5p/hTgSxAQPz0cKIaYgAsIdTpwQvKxqaoNAQkb
fRbCfwYhXAUAfiwbYOai9+gT7lelSqbfP1QmRCAqspZ9PE8BSdXPFVVQc4ca
cLo6WeVJFoG69SXqaVUuj24+YroTAvoVOOp5PlbNaEc6wUHbRaNjEJMu8Nct
NVp+l0D0sSUB9CnM7HSsvweAkbj+jo1stX2YmU4kQfveRbuphAnZMcRZppaA
fuitUVXap5iB0XY5PBqpXT/I7v6SQaNv7nG7plHGCcorZYAu1voOl7K/dfCj
7Is4zlexiLei90lKCBfcll2ZJRjK662ni6WRa/HLU+g3obJzMgTWzO1YNtYp
B1gQoLvvb17YSAok9AbJTsiQJYgvOHTqOnqorQeozAltRbiTW9OXtuuj6rVk
ac799ZUUtwuEVwr6KPugoeJP5/5uoEvB4AL4O3Jw7SOMfb/th7FMoCuGaKGK
pBs4VzmD7gYxkr+tT790Dhnr0YoyRJfOwqwbU6zysDWNwZCzdCHIUwFgPjJj
MOJWLJxBtQOxniL181UvW++62HIcW7bvjnV5KW+VoImtIJyNQQFwnm3coW0i
gZZlzaPqkBJJRwiTTsnu5T1UWiPNlOQ/WZTzaHGuoPNxjY4gIsFxLztwLN8E
mZ4wicn/KWZFoH/1ST8NLKdijhYtFaZc5j1AiQfr/vUCV4pb7FOFX8DWCR9B
s3nTwG2HhIlGwuIfSoCbXhEWundL/CmQYIw9r0RBmOlS/ZNfo8rxvM49vZEH
ZRPA1eAdjWoFgbEFNaGSxiy+BALMSt1CKhnK3NrGGI1ommAe6jqFSK1d1C1s
nMCGjqdKNiuWhiK5LyEr72P/PYHmHRB3Z5jAt0xf4UElUkrWwtgSv31POM0W
XwJldo3KcYtkzSNZVOf1xLZxoJpEkCHTey9xmb8BA5sEGTzYm4urfGzMWv64
9pvZTBGWhYSvv6W99OlUiv6sZbH4DpSP3eFGMSp1dptwcV4nXuuw7ABFYKLW
Bsr2VhIIAoOitoO5k8BjX7IE+48WqAP4Z5bPLNiyd4aV80/psxoKKwX6QAQv
/ge05sXjfpy733I1fdBmC93BcFI6GcrAMUxsrpxCQmBzkWE8lm650XWfE0cV
9Jskqw9mGKkY48D58CFs4ibC189jkv9LOau5l72wLJzhiaBCMmwHa6nzEdGM
LgV6EdyCQUAhrYAxuK+EgWfjYPlfPOl2I3QOs4c1Nc5CG9fglu2w1HuY9Dug
uU5qoQRp1Bnv/EFbQyQk9+p5TT8WBtPUTZjVGIj8NLsGNosTDn1L28/1Gqkn
T8QI8bKdG/KAVb/6I2vVeipSADlpkntqXINt7gCEeF1FbEIcLCSMRDb2EDVc
7ki3eDyb4qn5J2fHatl4vUKDdZAzazApJjO+0izde1uoJ87SpYOyA4N6Cdhn
MKuWrbk1NpLemuU4CSfwrqJ/P9eFRtiNewhcMyyMQlCKIIl13gLJj3da89bT
d5xJuOvyDdAtaYdjhhUcPjmQNad184VJucXDvdMax2Keq+emzXCuH8W0efGL
PZ0v+xTg7epkuLxcuAGW1VchrysW4dwosuix5PtpNZftzlFYZ1pAZu6jtL5P
6nuaqn7xulYUEC7ndN/bvkT4Q/cuEh74AgL2ycRMRO3/d/gRR1kfoDK2KnKa
O9sJA3adtIJf9zFw9Q2vqPZ8rRj6zOZbQiLjpxnZfFc/hOoI3RhL8CRTujEo
2U0NvG9J53gV9TUuDgHhRyi3CoZamWG0izWnQYGOQ+ZJdvWffB4u21ltjRae
BlBdwBCFy7KvclVrVjRu/k4ho6Z/8SAE2SU89jIIOOd2ZVCee6QzqR2xZJbQ
mhDGSHw33dCbFNrL2a4LSW9hEPMXZqRr7D9BoPGUCNGZM17I6K6yJIEea/gx
Ar42RzN5YU0C8Unb/bWIwlgqJx5c8I/FfCfHNAHpRKixickDtJRw+scAe1MJ
kmwUdh01UkG2yXhc392wF62mS2KBJGRCclzibVEOY/pX6FGI5rUHCScrj6gV
AS0pz/0Z6sV5fSr27WArHiqTPFr9cm1ZGQ3jpFEs2qUvAiTf8U9KOIhuIltW
VB9Ft8JzAvwStdwpNxF8F+LVAiSGwR4qIIHHOvPYbd70F3ZXQ0nXH6l4JW2a
HZWpzf2eDnQzsqGqtqTjyO5TNIhLvsiSKln/5Tif1qcVYZneGTdXiZCr77u6
Dk5bD3WK9zOV0Ct/YQSYuASr5lrHHOrOSks7VC6xovdDhwRqROMeTnv9yYm2
ZiSLSQHjQmOuSxQxHOv37yrBNuj8YX91HybnU/3m+GTyJ/n85uYTAID88SD5
kaFs14EbI2Fr/sNHrKxkdoYQneRmw7CtL1HfSh1l3qdbRJFmzn2CTjF4BYEQ
sYRqEph8NVuLotGETTUg6ag2XK/72eHKNgcO3sUoCeP6jqBXr2TDzsAjLwdn
1tYxviQkbCUhpb3ZTnT97IdMrvNjN2wej2YHFFODcKdF/KjppEj1+A4WF98/
Z3MOTSXPDUL0edw2ioXIWVvdW4PWX1/K5rGwLMKA/GijP7jLnGWIyX0tt8HO
oVw2bMKjTl+Wwt2a8tZ2ojK7I9CoOvsYo3wgbZhU0/4KfsBzQB0jbNfEUK2u
vcgIW/IO5tB+75ytcxfzeVtQfc8mPNipeeftZJK2V6M7Puz4bKzU3kkoyLJ2
Sg/yZp8jeKZrXTh4fgCH+fjggjRcwI3O4BILVJnGS4rOZ+Er2bQdr7D0tPS6
zbLYBHrKdiP24aJGjeXXWicguviiqCvf9EcDuh2VavzsqkBPJ2zzDwx+d5J2
UK27f6eRPx+CcRtE5yBqnu1Z92Gq4RZSyNWArJeu4NCLzcdUZTUA3Vs980vc
4twi5Mg0RAAJqgDmuq4q/ovYn/cF+lf2uj+EwtfiY5adiLtI4jPp8aJsY3Xr
m4BxIFKzznTgABP0GUeT46qbWKuSHxlOHdQRHJQmX6NqjCHHx1oInCtDGSty
KF4jjzxMr5RHEkciG45aBbgfZqkhxnRRu7CchwfK8HCQtN0pFY8bJhkwb1+u
ntrJYmZfwoXjEZ7lbZG6UeVt1ASTvZvFZIHFQFMi5fAJ+7DjnD/nRzbfK0HS
JtUhh8UYroXRX0m1IViT0DtSg5hpXCjOqW0vlRGQ+47uet5RQRTx//onVYY+
TTu6WYqa/718B79IlQ5nAKqi/rOFi1FwttGVB6x95+uOucM660ijQbHrOS3g
2YoiAYU6jLrqpQGLPodHq1ullbp8jUrr7EAvlSx+h6JEpEWIBVB9P7MCstVE
mNlW36UZsWftyKd987Mv4LMLBacQ3jhSuQQGZvFLSAo3ihk2acT4F2B+ZVsa
colTlNpjwekMUJ8+DJnZeg5o1O/LwC4xtSYH4J+TrvdPTn3A7ZH5bTzA5MBI
RVf5FCMB8eBAd3uTt1Tdl6l1MvC7oMdm7g9vkXghadpM0RLBLdC5uXKxmPNq
mEEWVCsjQH0bzzyD6eiepXXjQqt+LYPx8hNv2EWGN9jPV1b7A46Knum/koWF
z+lQ1yGhtvaIIVtDzHSJjzmkl2p149o6JvEXyTqM0oysQb5SNBwiWYCaTG21
rerXLqGDguqnMDSkpYWNoOoBboLm6vHLXfnJnEfxvPWByPePk04l2BSkIF+0
QaTxvMhWsqJavuc9eyst/sdahPMXMIVnr9zUV+I3XGYk3tqby7E2WgFWnWek
jjyULELgGhp+KBj30psPiFa5mGQK7YF2F0Q1gPOOOpxqLoZLil2O8z6LygaF
qsSfRK7cXgQPxtTf5U2TBjVrCfWJ0XbbO48bKMB3fx3wsfKZwhYFwvQTqPW+
80vu8O7ikOhTFuBSO3p7yvl6b1yRY5uImoROVmXD6iBUK9fEQVq5Ix1YwjKb
r7IsAjOUYmwwn97D3gFHQ0lvyY3lpmevZ3YVMQ3iMf1YrnQpt1M+JJbMJGNt
NqjxtAX3JvJaEAD2Dh+fOWLUb+AqFbekHU/odja7jysye5dbZbe9H0u2lXk/
ISIcq0hF5cZOcYMeyUIb3i2j0ZjFKo0VIQdoTexVLUOc8jAIKi2cA8aFQu7i
FaHEEs70qSFWcmIxA4GAKXC/9m+qgCXgtBlmHZExoKOuAnq0pGrO1ml8ivrl
4tUKFssLykC6OISG1sNOD/dtBv0wg2ew/m/mhgN7VfX1to+u/K+hfBVVP3+Q
HTiNNY55CgmxEnYrkiYRMMaYZj5i/pgf5+DEmyZ1C5gU5tp5D+jqbTioJvLc
+FUtPr6Zu1ydZvNdH3YKQtK/BbJZ/fjXCNT3XmiAoQEpR/5PW4yMGUiMQy7l
gi/WkGgTPXOH3K3RUTh5EfzM74zJZOmB/zVCvgZqiG81dytA3ZUuZJWJrpXg
Pi+I+EyL7B/E0ltyBsIuiyFJMABnu847PVl8OUsAVqDztwzHA+kw/F17veuW
8wLe89vsXzWnXWn/spKztRbHSzsVSU22fipglcLd8yJzIUYGdtEcqdfPpyxJ
m+LJIvJs5wY+nRpl8KaQkZ6LKQ76zRRTkFAdhEIdtOtXx/pFd2VBAATwcBpz
0XIkbSh7vo3bcn0mPRncnB22Cyzhr9fJ+trZu1Bn1ghESIOm/X+bLa21BR/c
7Rjv5HptjLJPGEqxJNPpSOMJI06NF5cVrH2E7o2Kzw8kmnBIY/r9dfImGWRR
WzOK+gImykjxEEu2G4mDJyhuCFMcC5KUflbRrPF3EUOjqyGzDfbkz3sHgvTT
lsbF7KXClwOwwYrmxZkDzLoP7dxQdn8zUI/3NC8aRDrET0HrcOvMu3m1EawC
oSd/YsaOWSdBFHyGYMrMP0Lt2x364rxFhYuj3jW1ixIVasjEQgS+04+eQ0dg
EHnYTvE2dM4D0zAY2xNY/mvwpnoI5+QHAw0uJK/DetsPgvHAEsVOFu97eDC2
rS6Rkk2yOhFQpX8TQlbc7KyYr9fghimH8yYVAq/nfKQ9JXtsMMfM1IdRm3Ln
jOGRkOkfICEHX0FSIrRh7KdkaPtPl9NNI/BXOCR4l6Ko+VMAP/kslJijXs2F
2NUvGFn2B8BvXutMC3HZXZFFXWwMrx3HepDwOPXgg85Wo2S6iB+gHGLEzTjH
zqm2qIgzW38DwbXagcnRQpkAnb6MEgyu8xA2pxBpVygyI0wsLw8Ow61qQWmN
GFcYFwOFVmjVtYj+BCBwUtNZneS2KMdK6IEExSREC/yGX5qspUfIU63w7wgj
2mA75PF6ISlNyIi5TDcUSOXp0t7Pw/wFhEH6ULWra9CwfdIA2cPc17agxnyN
hOkYEag9E/ibKhIzyZWPcqniQwxjodTzRK1Re9UwkhkP85HyqFE0lL80if4h
hfNXsiljAaqRIVy5KrOahpS4gOs8sVeDYE6NIOeJB5a12T/WnIOmrEOxUo/D
yQiV+mhxdR2U0+UlAUsABsj2/sLBbOcWh+8lw1sDmPHcl98hO1/4vICDcOFm
e42+w8w/Mi5LwuV4dtOc7sGfywl+C+dHFKzcB/DO5UgtOQblRwZOubC/LhlW
/N+ZVYYgua5wLIgbWmQd5BIjKZgY17Ewrq+cBB2cNBzk4p2CI87ipHYCRErG
F83N5qnzAs2B5ah+RTN7JFbCLep+iPKoz9wefVbLZcgxzXyYzbMMG2An644H
Lra71RUmfMJFe+yWrAEukbyqg8ckzpHhRelfAlDTCchaYyiWpLBadyOxbWQn
OTtSjvDdZotLCwS+J7yZd4IOWpMS4NY90dPcMvdoJ2AqbZFBehZnIkTHn0qC
WEXjoOEWp30VKX/OzHbsUTZ2HTiVb3KJLsPsvBxKkkLDo6QUv7TemTbQXrCE
RIvbVA7Z33V0jtfM6PS1geqk36+nfGm4SPwL0UA4zX2KBlf0fB0BoRNzV8Ux
msfG1ddl1CzssiEfqMTXI5xBNdAcLxE390YDvV/YOqbHfD5APLm9jCX99eZL
21Ysk+L9FD+iQjb6hDv1MpDGMDRw7RhHVzG6AiP8pzzy5s1OGWcTsSWI9y2D
96P0rrsbdcuhptRRknveYAGosdAG0z/TvTQltL9cqik6Nv66mqVPR1+h7h1c
eZckYTw9/njwV79m6KeprdFsjocebzHq1/RSw/qX+YKPONgUXNrPWGDhctEM
/BQHiG7pcVJklpdVSZz1+64fbpkp7+3g1WGkQMO4qLfNapCIWC0LIgm+hygj
JYY44PC5sQ0OAgtvxR0xsSt/aN2s1ruOucwutdpgvI7XlPlkUqetIZG8utpc
E+17mUUSLDiEZVMUgIjKVtCtne4BS/OzlDdWyKLuAJ7qR3uRBLcA1hVrHcF2
AfvGDv5yINwd2BbuoNk/Ed7iW0jxDMSAdiuOFtXNTJw7W42DHGfdUuiRcJpR
3XwtiZFmrqZZLQdP92+uLVMFsVL8OI4iM3CssfB1bnH2L6zMgH6+Mi21pv7C
7BZvCpyRgl44/8/l6MyPZPPxsXFp/fHV24kf4E6inrOyBCDGfVZw2XSjTSv1
H5Br7GUJqHSHRDT7ECzdejQJryVop/l99Ou3xXj5kqjF0GoQfhwz64sYEOdq
slNegAIw+O9fuuo/ll1An7v9F+zrbPG5Bwqmp6OOxqsAHECIhypDUKWarkjC
r3mag+W9Ucab8h1Xjl1SYNCl8n5sZIGeT4EHi9tVjzy94QzENpr9JnRkL6+u
ylEOHJMFYY1/nitPv55FIE+CiF7iWZo6bot3xoNHgFMojK+3iUDQVrWajk/O
TE9aQh/Ef3PVr0HyFc0kvovbaI5D2qpaOcK1fnyr3Gjxv2wveXZESy9+Rqyy
mB8HKYDMnlAy8Rayd+oKx5IqCVMlqLoTr2qOnPOCV7yBtTSUWPUgaquzhyeU
x8/KnJzmoGXE3l+vKvYH8LOH/aIf6ljnvinKlcPZfPRvzNBNJl2iBlT0pevf
t3y5vsFBaW7XM4qHH2PvXRrROgYZ9xEFz09D0rBuQiRzk7Iblq8BqKFnYPFO
AVfwld12jbRyZTtDgeLfo54kwc/tgOwaos+oZGSVR8202CTForW63At0DvDw
JuBNnypzlMiyHUvKFFGsktagqqFthAE4b/IQrRzCJA7qc5U+Yz0eL4E2J0Lo
Q0hNiRgZxhp4+nlkrZDCIkqOy+bszKLIuc4FJ7VzowDvJ8f6t3Q5PiCVLSWU
+eGa0jBXLB2/UURZ4TU7rnZBRvpJkd4KH+hUvFIoTUnzNfaaTZCjak3LoJRk
TivoOix3s6cwSvwgtqCelhUsPxFxpnAqRzwhBSfRTPH0tJioNDvn037SJXxC
TLtkEADKkqMbk7J8W0Mv9338zf19Q++DI9pJI515t86zZoCNaFRgx2RQJSd1
AhV9KczVri6MLGN7ROZEB9W8Rft53ybiBEURg8uN6he0zelQS+c6ovfiFjnl
y0v7vZ6EJPGQEUbf06q+FUpvcRKDh1mLhDeGnQN/33yTM5bxvyqqGg9LQp70
2BFxMPOIOM461Ma25uFa1YZWi4fX3QYiVWOejTeeC6GLzRpvb+QFd7Fe8WQH
J1YfwBAeAVhSVv5K+iT74DIw+EEqv+ZnA09+OECo0MdwiZxrNAfd7UbVbPWs
wq62R4yw7KPWrgVhfh8wbbmcW3yPe+ZW3Zn2qvW0fXb5/KsE9FAj/jyjXynz
Sgszc3OfNz6IxBA7m+z63IsofibO6j8Y7+dmGyyEM3mXIwh8pVj/ZhVRo173
qIDvCUA2hfeg9HLuiWQbJ0W5XBfDYeHwNR6oDA0D+Ttlz8oyPCmguxPbtbd2
poYkIahYVL2PB+FbyK2O7dgsJhCDC5Zp6sR0OAtsyGQSLyAFHKSNJ+Kbz6cV
4mklLa+J8zXFd3wi5osDaFW2ATWpwKyQkEpSnE0niuyOquRgV5JXr3WKM3Tv
QD9+l6gnNMkz1nzkb5Wqxvoi6BJg3vRF4XiRrp+2XgUg26n4QApWQT8MrCaJ
7ot/fFKZjEwEQ+32e2AH0FP2PXVyEZ3t8HrZgAGBHW6S/3bI6AHaNooi5aQE
JN3JHIqFXmRxSY/1qvnBPNiyYNFmidsq3NSx/kJ/WvlkQJM1Ln2oBoI4Ghlm
dvYR820WGicUEV59QmVZjKkNvl0K9ugAxI5XdhDkzys9CCqqHMcJ/s7LEnC7
DcnTRRh9eZ27F/ADUB8UrKS5gKHgolqlDDAKb1A1wQ44V11VgcObV6DeYHAg
54Rr2Obycv6ILw/dL5nzfi07wNtCrbqlLK7jpPORPv9Y4GetUQrXlpcgF2RX
wEBpKcVgO3uly42W7HbIUy3olzvWJ81jOFv5OYxME1kflNtHC2HfbOKpIIEu
2oqfG86bpv7s2bQMSE3ZM15MZAF9sOivRbKqHljW1Z0f2wzhefv4dZsu6WJh
GEsZwtkzcqB2uuRQceDJZX+URXA9KczxTByLXWErD11PFdB+OgbHbzPvghwx
o6PKXPfjCTH66ZcDNVHr90OuwgVGnrs9hi2LroZrnXol3qqR95o0kgsq5lBA
MlMlzXU9T9O5gHmj6hrwQy0qdU0mCrbcTfFsQSjj0lq42nnGmZWiQv8Xqqqi
Z/pmqU7rjGhOD9manQs8BENSRzgVwi+tDGUzgRobMprrY6d2CSejmEuyD2A5
rDQ5uAKpwCuLJf9RRrsnZ1ErfAH7ybuzPhE+Aowu8cYqUYrwuckob1S3IFTy
mXpMhOHjB7jlIaAznNAsSckMYSO/2MRik7JvMvGA8SeApQBCRSP2xf2jHIpq
lozPcsi5skRMUULZYoF6zGiUvrKkQ2wAQDOT1PJcyG/fuE5nREBdCVYe3cx7
DxwPXGZIC0jrmFXIjZqPvgYJnzG6fkGLLF30sp9Obzkpm22fm4uOG0ueY/f8
VJpZ9DXvEk/uad4qb+lG2tKic2IUdZ+enoPYL7dFNLOmDsOE1K1QhUe3wgdl
GHErAqx5B41Ok36mcSG7ZRZawL9Z3i0SFze8J9CRnKOlxSr4fJwuYc4TFQWa
sSIAQa68oExgdEVsBkcKuBrzjImkP4cEc2Ey0qlc0bh9Pt7NHijM6GJJRzzs
5IaOETDUM6ldoPoLCBnMUwOXEuxPqdfH79dehwBYJySogycXQTHmjcs4S59A
OzV7HL7VoNygCo1DKfYqLpLzZNOA6W5+N3SK4yeoGYDdBY0eGf6GXNJzna2S
WljkA18oAHdd6Zd2247G6pdCxm6d805UoQeVb/uTvwPYDTVWTpzAWntluIY8
MksBIN0VNaOSi4YUC+Wykwrjn7G9VBz/1Xm65WbM3OCn+CkRQ4Iev1/II8Sl
SwndYiCYpQI7ng/avKYSJwFAqxAPvRJkEYnsnqPPu8Px7DgLinddhgoADIxA
f9jrdd2sZEXg0gB6I7FiQSBifPTaZM5LaPoRwCFp2583GxAN0EnrvFRgxdfz
l5hoebEo//FuHqnGWuhcL6FBYzfqpasvLh2o/+sIbypp9DwzE31Y1EVP2uZN
mz1pe1Fz/HTA0HFWrO26CBz5JHlz6kOsXOg8hCRBXSFepmIsa6W64ZJU9Mvu
JwXI/2snH5xDj2ybpdlWPYT9ozoPWX7aXPBjxieF9JKUWsjccXDQlT9mPG3q
nufdUSc0tBFXEe2D5POaedjcaws8wfk1bgLADfjT/MVu6cVvNQfzqOcznFq+
5Zw2mmhh3x0VSWybo4tZoXantu+rwmD8NNXET7FZc+6pUdJ2R/QT0oxq5FvC
x2Kun8Sj0Y3l7Uw0xStuES+nVTwaKM5g7EkYNCGOEQ4mJ81Gg4+3e9QZbXvK
SXiJbENtuAyPnCRt+ELEtfgm3wI/zJbVURo5u8Rb7469Xpf6SFMfhGU47WEe
jWcamDf1eYYfYP/FUi1IofQAriFiAPbEbe+2XUFqB90P1iPKbuiMXvMIHVr8
1pSczcPOpOfafYFBGDi/D7VrkTfYT7rb6CPSsOaBksyaK1vSBwYxlGoQTlJx
fIM7Emc4h+LJrMRzQ07uZe0HQDphgFKUAxrzD5vq878VswZFjn4znvXzMYbx
gR6/Xnyyg3Jx9DEuR8swbRZaRDcTiH8rTT5krduK+IKU+n2BDuzHOo7Vjrel
/gZux1MHWLUPTFdgu5iQW1Zexa3STvdNH2fyGSrLzq2QnDOKZ4adExskNNoq
xgjYHNr/lHg3v+zZ7q9/FOkoEpIiPUDf1273wqedLZZEfIqv5lXcw7QTNMMN
gwYdhGwKEDua+YLAoYo2x5hqkJv+DLJTrbukZAqHjbenzPF12QvUVdSKf3qM
NiFp/x+Q2LQwi+duUsB//zWJCv7AVdysfZ9/UuyptEo8PV4Z7UrK4CtRZqHE
v3zSdseZ6uRnrXljrDt5w732c3wQGf08p9oxtuNoRs2v7Em9fdai4xJ2qMRT
+2ltLwYwV+PF6L5GewSvmDqYRDgXzqlcA+5dqIEywXgskreIdiBj/LZkN8Ol
eVyupl9KlIjaPtOaMUyPf8Y0cw4kzUE0dpuRl7Yv8XlhxKV/xUNeI3/+8ip2
V/GyfIU3GK1synfBGy+oiX68cZmoSozjTRueLVyiTrr4p1lRorjpu3nTaRR5
XAzdXMYekSzT73LrbtiR/A5OBCGXYrsC/0mv01nwRznpt/o7d33sGEHWxSyQ
ceZNjIEJnhwSjU4wyo+aC27SWhoJcQAfySkQBfVBXKoNNvFZsXRZY4ZrsUJ7
3TArqtI7e3Es2DY8Dk7zDc6NgSFc1E+DZDjQpozmYzM4mZkT4i1DpgGWbUWI
eSyn4GykuwB4AuvbhIMJFTIR9u07UqzaXpiwFJ7QuJTOpl0oL/KXAQAHG5Hy
OuWSwJMzVRIhwIhGWmkHlsbWoAWSA/IqHSItEGcmG+eynkgW4YY/H8trCQQJ
X3jPr6xMLVOkSBDIij/bXvJCFxpRlpT+/sxDxebbvVhehkGfcYV2bSimxO4I
KxCM9lbdfa5wE6Roa5hLvhtst53sjYSthq4tjFMVtZXBO70p5/XBlzCovyQk
5j+W3CI0n8UImK7Wlh9+L8ig8vDiprvbAYjc0zy8bf2jWY5ppAYI+zGlTi2/
PD5wkDkuv9mySlnEFtkQquJEwRqhMUWDCi+1FhjVzfnPp1oli4ly1USa6Tkk
h+5GId7JwYOEOFYfL58D0Z1h5hWkIDYp1keyVU4LE2pJOrj0O1jnT1Q83/QE
c12AdoDtiZizTP7NPUUHSui2XYCmGmTLLf8NXvGcsIsO7WRVFwWkUjj9kLaY
nSq3PRJcydj+VzI9dGM9w1n8kDlVoT1rhz6gVXnrLQzotMbnR+YkEBIqXqAS
NjX+oRzf+B9hzShAI6M5bi/gcNeWzN+o9OJ9Hjrk+mkxmAFLaIK5/dFI0eSl
VXcWcOCTVnbEanlf9DPyz1Ny39w1vpPQYPUwQuT5yEa5/UHTpyGXvpumbMnc
gPJfjQg0YtKf+zQKtDXtpOPLvCmssiZTzBnCtag8tm8OCAh8Vb3K0Zh53gA/
ezO4NvvGKrGt2ixJC5v50KekuY8/1xjhEgx99qWKOaGPNYGmVjrCR8vKanTH
pkY2tRSZKSq847nLNDEGlw+GEEFKEakLKPuD+uiB7VQN1ECGeVlEDtwBRr8u
EI0RBgFFCprI2tbtVc1YwPLcMe04ccyH2no8dHb+shx01xmEcb1Y405HyhRg
jZMY0tBDERKZmml0OPWpINTiYLwM1aUhEaS/zd8ipJoSFpDH/rlpggozNG9v
D4UK6I8qCNGLF1SJLgpN4chd8WZiBLDuGr2/GgX+MTtAD95TZ0Pl01+V9ETP
6Ygxfbt16uK9h/zDupfOpA4GIuq9VqWH7f2hjZdJclxoMrv1TOt7O4wPJyjb
krmWFZ+OaSe4PuBHoD1jC2SsyDNemCZAek4/9cIO2BPMMm/RnEGZZeRVWbN+
OJdAY6X8pFtq3Pw1rUDpCat8gzeeyQMMAm8Pk+6vud5GRWZFWAbT96yIKA1O
e8ZlbxocfdPYhK8N0HSXqYyMU3lw74vUutI4cwcTcrBT1ZgMwEOacR2cJeiB
cPaHG3gIyj2IcZcCQ74EF9FFBfC7jPeEjAABmPAMBGsIms7IgCvHCKqALYp9
yFOIYlt7/EagfpRhYub9xxqbX1gMZMqW8RMjqBlKqjfduoms32mKYypjWtpc
CWFgPbv9GLM7yCZG99eFWQ6t1ipOdCgHV4sJrUPg4q7Le/ZK1Z8xz2Vq2yrk
KpAa20GoHpOCIIdS5vT3VpimvHEd7Ngnl1gg5RM6EDXZBiYdHSQ9eUNDrYRt
5CW+tbkmcBozkBBScrbGga5rZNoVeMKlGTEvZXmoMX3M0SGDlzyGIPlACG/K
C78U3/79aAan8ecPplw3w6HXPYIAjFF2dJ9g8zp8X8VVUVmyAmb7l8HntDj9
hK22QYmsEzxn9+E9uv46RSdXwmkMsgESNPEWZIoxhpVXTwXegSLsL4qUZ7SY
gFcy1TeoWQdmyWdYu/1Oj3HLH5fSDKWkc0qRfnpHVoWNFJ/Fc3UZzU0TfgXv
/q8RSfUYDZy89EORACr32WUtHg2UyFOmcPp3kVapn+uHNRxPg+ViEyr8JC1I
Bo/ruS5qwHIaZIxzPirJb8Wa0hzuIleYD6DPgH5tSLELeov1liLlMfJY88QT
WLn7EWrFp6ElzoC0jRcnJMlK5DSATOthgwosq/2iFQIsIu6Rxudk1egcr7A0
GOqWnDlvmbixPk4fGBhIKdUjVFhrCxiskjoEEsMAUfMl1LRG+3fU8LVAvZaP
cgZN/xdu4y20Nwz/A4XGQuyWlAawLhqynTRapFtGUUPtV474mFl3geWOOJwb
oqBwczeyW0q5Rx73LQJnapZys9Qu6Y1DjBJsEkZg5IY46x8DpAN4OZOSyKg5
hA/OJSiD9Gz+YqpmMgwDonybz9upAZ9vPe8BFwyzYgzzbtr1leg3mhcyza56
MlXBhWPAaBvAqI4asezye+47xf9MMD+boH05Y2DV6rvzBW+Ph1TNgQIiNMl0
hwv8wIfgLCL4bJxf+7+rk+sYLdA+ZCtblEWDBU/nEPrtCTZV01WqOdHVo+vX
dbHPhU5SQ0++GxEFsQhdYBc0JbhBMIv6HbjJmu+eHrlBjogSbV1nSiCCOIfp
cM2FkpZnSrAuZcpX6wSqX7v4oyfzDr8anJ1lOk7Zs+pXDg0HGDnm1+VMtxKs
IuCZ0Jkj62li9UuGC3hRzQIcrvrGxspFH5ZzSq3IVtPFn84rgjpGJs9dvPcG
lfH+0g89SQHzUt3likjYHcLVXlQAV7/VUl64UoDB1mMiYabiaM5fX08vmlDT
YdMWupwLnvG+LjLx/VEohl20w1XsoZnVxzpYsje9ktZLO2bfEQt+LK18lzjZ
5539CUXAhRNikfxYqVAX5W+InSv8QzXJm0Jq8S+cFufJOXF0gP0AlvYVbbGD
ZLAz1m0OBX7m/5u220Wj2P/gjc6WBsaIVd0CSL8MVH7jVC+ePop1ixywn/PE
/YTHr+xHXdYi/eHQh8WCubJ1DImg+yEFIZrYWqdetj4+aXHx9AMXL/1aJ2Wi
S0Tba7xlWmhCW1AH79chtYBufbNyuFjjos6PoCPWrqnF6MM82IygsLB00d+V
qVzTR+u57uoDfybms0KZ2a7lbFmNLiCBbHXc2qD+X9Rp56RSFk2eH/xWtPkP
QaXhVFv/d5HjYsgk3SKcQFEitMHZPtcjE/oz+8/rOet5Ktl2AkcVjQNS6Cbb
cnNHvK6jN5L/IJxpT+cIMjNvYcmEZkwftza+obVEgbgxlwX087t48Z8iJUdv
xslEjkYZqHI3ScmTVir6b3qZHN26nNDrGf5cgJm5pAjnBs3UzmmPtEpViKTZ
Vti2/eqKE3SNAqx5xAcs7dcoJ2hHNpEMuXSrMIDsCFhuFOQq/xcMCyQoCqI2
3TVcyz0SfxfOghBQKt+00Rks4Testf92AQst12vDqcZ6n6wQnmjZBUr8n9kx
xUxJmrV7D9ErP4DgpemgNhG+yNo8ZRX4GojiuiSVNPo1oSWAvYNXh6Xz5J7Y
agONtDad1CFxTGStD+/K+Jow2RWZKfqSGTx39NfLePGCRNQYEjSDJeSBWc6H
rL/Kts0Mdhnt4bbmYG7xMltv0zzm2zXfySbXfGZv54P6/ZPX/0M8A3IL1YlJ
YKCtV7jnIhOvWupoH4N911y2Ok52RGZlWfLfsGpwu0+ancsNa1cveaoVbuhc
5VtgL7hPqgPNEBxRZpOoVB2+hpz1Q7L8ezOXVdA4wX5LhH8LLLxdSX5P1mB5
xQRujOPPT28tql27FISjdBlJxyWhiAtP2xiPZF2FEMiyD5wM/v85nGJYitv2
aMpX8quxAB34RKHPCmCmvCuIEIKAyk2i5SghJYStt+vsgZeFkG/Rd0lG7nBR
/GYF+xds+R5UFf3SRq6bYhe+u78YIMhRU2q6YoU+JHJhZ1McensyPA1vwwog
gbbqSDHgxoLGODdXxsQUylJ9UL30hnWvhNZppd4hbwk6FvYvFZOGqRVk0dF5
RxaKSDO29UPLA19zQsaXw0/u4kqvGpyqUM9ttTmyKG66ayseMJa7pf3j1upJ
yA1dnudItNlMykZzdLDu5U6AA/DXUpeEKvrQizJ0F3PWFMfmFA41y+G94Dm7
Yd+sQeKhC+WjGIbXeayP+yyN/goSLtCR3Bg1cuZiYNoTAPSno5LEWx2dmkt9
iD0xdYBY7Q/921NFGnU3ZFgz05uyZMXdPw86IrFR4qM1WP/Fbgdep8B+SJ/s
1ds0/mv+PbleYpPFoLRu7iRDMYEN5psZYvFCCCUkK7+LucbdMWYsfHRwYdRj
Hoxi1JRfR3/zqjhvfZbllrYzF4i/QNLxQBx413CYbXtHD/YpxLtsYZv2mC0J
yjDdlucJdYCRVpXLgL86rNqSPmS4C6TspRRNO0NSxVRpd9zlx+5grpsyERKf
8oKNlAXFLsSw6Be05QoUNN1EOCiXTy34OWKeJC6MmHi0uKgb1eEzpZq+o6wT
ArEl9DzROLRuh/nb8ra1Ii7jtKLq7hvINthuFRzFXTCtUXrKuS+CQcPDXhZm
fYnZXQgr72X8A896VMf04+bC14MXwi9mQluW+P5xFiNKoj+Q7SsFdRxbd8E2
GmsHtydTDAONmTOEVVteW6PTgL8vysTjRbMIKu4Jssg7iCrs8RBX3KNqUJN0
Dy6AHaV2ggN5To8sORxLt+1jlo223hf315bJ4buxK6UD+gBotMtRRR+rV4Fc
IUb6Ozql+0nf20ot55qAqk6reQNGdYEE3epHqnjczwFOiGtaUYfOgLxWG264
ClziQ+5uPdQ5uoESxnW9nXXrM17VMD8qqoRq34Ov2NlgrupRn4TZm03CiLjI
wRI7frwdSwDtapiW4zR6pYLcEZ5bbA2VWDYZQ7mDRDcmBEVs7/HKYbQ60UCG
io+0MlQPRA+5f/z+zr9END1CjVU89leCCXqukZyYLAG7r4CnppYKhpwkkPcw
m7U9MHAhtWW1d/o5x2vwS4u6vBhtRDhe5BRbQZtlVVcKXoPtHOL3nd+my9yG
SE2DBYb7AmLxDOZRKfV3NLgPlc9SwnqFYaxErbNoKxPu/GnV4uJhynPldiQ9
eg51OdyexHGNvU3WfsY7QLFdD5CDraJS9UjJ4LmaI3xuMI6axzMt5TA5l3Oo
wisNWGv+V+aYnGPs93/ooiQoCZn+f5H/79KBvdpsGmC4GQ95R6C7PHrkJsJf
tNx8gxYwNVaBj0JcqJ3g+/3F3QfWk1BSlL3lwp/jzfe8rboTDwX6M2sTpcE6
MF23+7IlgpKKT4J9/TO3Y59ycqmBj39+zD3p579ULLXBXkQ4DVX3/temewyP
/mndXAq5Y1yCxqbPmNJH7kcMXK/9OCiAYeeEYdMP16dznC/SEtXYpUnMkYCT
eADbskL3qgxiMgSlEf6bgKVSc8zDzXiWI/p8QmPsE4S8EkGqDb1Ef8Hm+oKB
UOORZdWCVM19jY9jNYMHLbHOnq78wQ3/sedNC9HsAUXjstIad5lqltgsqCDB
25oFiUIgBeilvGl8YPkflGdxZkWKERaibbIVznC9uOz3a2LWkbqCSnFbL3OP
TyDTF4cyz3yvquJYqv8xaR9h2L0dq+Y6IVxPrHunmJme3t8KYiJMOWGlDPvn
7a8af7AtWuBtnuLoGWbU3sjbAwkm54QK+yfC5ZKjlLw5QwFKe+r49/G/yn8H
oCBcl5T/cyLM1FA5Nq/L1Yp/D69UWqn6YimuRHZHxnHYUdhHp/TImmZ+uI1f
IR7bJ3eGF8RilvnNA/wGIwAq173gnqVzA3mNzSCdqUM5bI3pDqzIDivkNFW6
XksaEgrrtVGaEXvqzdYVm1YuHv8wEhwg84s9rP9VG11gp7mgaWy7kfoOcHIb
EtAO+JsKywej1GXARrsmLEnOQP0RAwNx50vHnVTY0ZCv4IfyP9ACxhOD9EsL
NydlyS4xkx4yEKvgasTMLiU1EeAcga2YEy00m3/KYsJKy1N8YdlOe80WI5o1
zJJ/xl0BeDOWj7wvlALCsePNRArgWDvRNun/rsS+mN8YkPcY0/N1yCZI70P6
RG3nN2tYIhAuAw/EMkUewrevSumHB7BxzE1LzhPxM7om2evKW5+b5oNjNwFz
nzF300aIvX0+zIG8gxGcDShF2+P8EI+c9Quqi4JphpPDZlUoTdHUCm2QrKXb
x5FJ3U3laeBOZg4a7F2oVuC/Q4PJekLTxm/E6qfKBWUtvN+KkG107I0YHjAr
WMpF823J9aBBAUXusPLq/l361G1JUN045vgC0R+bsuaGGcbb1DylQn3W25i6
bpOeIyWsirvMDw0j5MAEVGvSkjQRryjmUW1cSL2Hq7QukSEv4RWkIaYEVXsR
gxKhk2ckvyA/+KPl+2HW6bKmo/lSrfcOrnZBTTxf86x50B7pnadMsPeqK762
Aw6irsvptaJFFU3K+ZqOTz8GWWlJ9tTRpojptq0MM8zqZGQgXf1n/ywqszl3
ylcD7ErStyo/bRYz2CV8Pn7vEHFEPeC/222m/k41/hnBMsED4ONfFgpnGbZ3
WfYNDxYPvrZ6Q9DylWfonIElVgqolyvnN9m8e/on80ZNVjapdx786pGgKGia
lqJiChnK8eJjQM2KOSr8pr3htEJ0MK4cf1kEF7dzZZ7sYgX+fmrBQ54OvCcu
juJQEfV4mdXwxDn102ETCVvN+dgFWZJVX12CZuDWiLMhUQ1VXuoSwBXC2PdP
5Kevb6xSKhT0JQJg1gOGLI8tKJDjTLNNNp+sD5hZvXOV/4QVWOU3psLXwos2
FLovfwM0/qJXIIaBaQ0DYrK7KgQ8n3e9Dchi7/noqCr1+kM7+MwOoexyIpXi
uodLOKWv75ijhtlrlaQbFgbprkNj0vb+1+54+AZo5OR6JB4DgQZheiAEIMU5
GuB4BQLti4osWXHjsg+4eteCGEKg8KHtHmqnjwFCfNJtSMSdgT3On9CBcTKJ
7k6oIqafsuxtt5QNk3g//ZRnOEZIMwn8Hp0oheI7lNhxFHnW9fdYs2+o2XSj
loaz2spPPb0uDciM8W3//7O1j/TUf0Go2YDXH8AedcRREP/diGF8sEDabOQn
4Q3opycqG8pD6erICXHFy3yZbNVDXVDMYE2jFwZJYaGVJvqy94Uu1LhrfWr3
cM6hluS0OGNLuM97iLkLUr442HFdUMlAtjuGx/Ax0NVkx/xKNVHL5CmmbtNd
MKuUwMshURINbmkRfTvqcyd/5ZKNEl26qJgifuOzmbAekW+xRO6oi/scdNew
Jvx7MtuJxvoyDk9GTZuBC6hgUhde8FuYVh71m4rRKTbnsIrgCQg3fvPzlOWG
b734/p4R5i/wRd89kq1RbxbD2vsZYhOg0b6UBGsegT8yLJ84951Yr7rCFB9c
lUuammx3TJQASnMRJ0h0m1M/o7V4TBdqe0uGhSD6JA6iuR5vfuQVojdCS8jh
qWmXaPXt72mhzueAa/fsxRlq8Y4mQBHnsCRWyKy84Vu8eASQXg83Vtdgvcfz
W7X2MBPfi4600J/aPSwus6O8ngpHaaYo9AW3rtiOryNwZexAbd54ypjsV/Ke
LHJ52YecyG0bLJmZjepz9vXr8z8n8TRdwGDYVQDgdcrjG/wjNtqavm6gf3B9
Vba9o/PfmNaO/Qy/Z5db5o2e2g9rWQCvkN1/LNhoNhrB0WJOtimTjxn78rOZ
BTDOS5siNzkg5K4AeQK/e1Czrq9p2x9LyceOPviaHY+GGyVJOOZCAk+5XhLV
ofM/dGVO88vq79w3qyWVY5ohuO97dKkqZTQFYwBzDNZMvetoU++Sy56lsDqD
SB5PQj+YP5BvT5cTSXw15f1bfR8ccSRAxeOM02Mmb/Q2lN+NBrJOQO2LD2Y0
AObZnQyqkH48SrG/6tC107TVA6fJlWs9sm3owPBIwRcjBveNNxV9gUsZuwWK
VC3/+VI+sxxM32PGqk29ujlGthfR41mhBPDuskyXAz8yVjMwOpGCkzsaRXwk
L5R+niu5fxQrkesQ3RGgrdc7+7RGm/4runhT88M6JoqNACTSXfWvcHXG1Zo0
ro5SRcn/JQstY/7BRgzDU/HL6ZZRqm06nYS3fvHBdLB8Grup00ak+I6mPgSl
/2FFyE3G1LrmGDZGqMZG4YySXwS4VRA97UAaDAAmZJ0jc16slZviFa8ttkRi
xdBBb6jDWLGMelDReCXnUpK/Vp/K0qUqGMXa+iB6WtTjnzw08WST75NqYNk0
M/pAx4qJ82GpSSzX/XargFFKoT0/5XYMzGlHqqGCzTADq9neu70GzWtGDiqS
wABOYvD4DEZpDTmPJAUVNq4Q79WfTnz12DRTf0GaICSVqzK8yiURNrYJAgKA
QgJvjv2TCqssApWeoL275m+2h1ryaJXZjju1A6QnfMCiaFHe/NEO+PUy1t+c
EUfh5xFplLSisMlKfLeAf0Fkn/H+kFq7YWLuFRZKF3qxmpnRj3otVnA865QG
OhIgDtqPPa5w4KXd0VsB65vjR24p7ucVFmVVZURLsUf5AlKL2fsnI5UzkVuN
XkKHpMJJJQqsd9BfeH4BcruyUKAd1STzbnvkbNN1gWz2gFjlwYaJh05s1Vgq
cQ0Ag4oyfkCntsm+Fcpb9lLfQvXNmRtAoUGqXI7J4nLdGK6T7lVre+jozwcH
LwHnHOEDF3rVesoA/7cU3ncOFSYdLP5AkYbgzIYRtWHUSerhfdTe2N/wI9ZX
O6KIqkhEaxIemRpqwJ97+RgK0mJB8O/YT5y43yFGDzO/i5TE+El5itNPscH0
G+hCBM6pNVhPqUw7AJg6Dh172SRAiMsg7vlqhECl7aUvwkpiGTqrzVK/AF6G
oeuNgGEXJiQMQ1Q/pI+gZD1a28si01vn+O8gvbtO1KJAZMN053RYywIu6wfC
H3OJ5ueWFjap82kTh4lky1pujEVHIrzWBNumaDWcszFBjdgt35VyC6OHNkO2
nyWayfP2C4p4pT4DA9eb0+iHxZYSbZoSHfxZlStupditS84KGetsRS7fK17X
v1Og4O8WZ9k9UpSZj/MA99B0BmtPpGD5hmcdpFOzTXWCgbl6rFj8j16/v01t
A5Mtmbs3J9UBx0F1ZNbfD9f+P49VLGINa/snPmiACcadX5aIZQ/2ehWlyNGP
qSDpNqnqmX9RZ4YLIXTs1fSAkyamSi6E6oN5vXEHJQNp52JHLO4vMaaQ8lPq
esvd1FHmJKSWHaSiVBtjz8INAaGyvBA+HO8IdvsWoViIfXyLBrbS63JhRyte
vBVS0+TST5kk5e8Wws8+pZXQoJ6LJ8e42vsNOT7GhBoG1qDxpbx46nu50u9/
gEYm8I1VXYzu0Yn3WOsI5lJsUDGXmzr9kPZElcrM1OUi+aDvLv3IQss0KuFB
UJu1lGyslqsewV+zrCm0lFY3fqUP3UAFDbfiWS0dl8mKEgetaLb3kFkz4Dm+
ZuAyA9lENiCbdajm0ZWbWM9VX9E7J8Os+RsxCVMveH6LdbqepZxOK4ElH/vz
8TM6BmOQvcT/53SqBSMTGsx8qG7MojD15TpBHpnrk91apLNag+oG+F7IKtJQ
Tp1aBDnuj7fQrPR4oGnpOfPLmPUmquYK5/kWsMztZNoSG42D3g9rWWmbQyir
f7sbijVm2eaTFo5sYF0Ocm3x00/P/QuSZbiXkpsOsYKQu+nnjdQr1CHnbqTT
EDIbFbg7j23+XKSuob6fSAWFYLobvVLXN38nRTY0OxOlfWfeBDu37Gho5cpA
fsQVjY6zZ9WxdXJK2yT3ruGJ7U9nHxYbhB8lFiRVcZkuxF9DrLCZRH8ZWEbL
LU6AowmXY3hTXCIZIhqHzm0NCyps97LumpdNN5uV6frIVQSUVJBF74DDj5+X
9ARie5KyG+iakVh5U2v4zx8ZbOwo9vDNXbQTu/3dKmGbeBeq3l/VAb9JTJUX
WmM4sHur5bMzXFjdCHXA/1zrE4cI0Fu85Tiqu91Sr49NV9ZYOBjlASvQKGfK
2NE+okk9gLqr0MCkp+PN6VIV2+n+HMVxgeWQ5u7g2/KsJEbn0f3JAW0+hPq+
6tuXLX5yuXS9XF/YoRk1DF/+7TBQwmpz+5EaYy3/7t3eNHJWnlvxUXI+qJSH
1u9YxqxseyWFSDBYy1feIckc34+1PQrH5nk38nZ6qGM1jAqMZZf0AO1101ie
/ksugPB+bbmw/Wuf3bAg41xWVYS8CVe0tmsiS5yDA0DmL/dJXAH8CaHGqwGd
bxHB2pXZnJK9w9ud9DoAunyl6oelivdzA/vjPTKUkK+aDtMhRKpzIEls0L2Y
1uvq8mOdEXc6bnFvyemVAsJ48nZuZh2RhJ33txaJ3cat1vaHZRANRnfmm4Q4
l3uqdtqitNd4tICfjNNXvY14HMuNtWs/rwAAprhPYtjXxVpMb5tW0ICnfIUC
BCNZ/y71jpHQvdLp2A9t/Q8efOCTXll+U+lGGHeYiTAKD5NvAIk4is8wwIQL
Mrvbe+Hd/wg6tiiyoS75BC3bfoRwdm3HGIgk9+Y81wFZBrJ5U9miFg5qfdiP
diuE+TW1w7z/DjTd5aYfYr4BvpQ+suYuslPXUDD/qDoC3n8LC/uxfSoBgzjo
q+73qSax9pu2N0r4gkB1ujOTwZg+zNXNBemVzo/RRBJddmJZYPsQj2KY4csk
kXugxdmjwbPImxPyTDHN9Ypjh51FxBk9hkkJ2ceKjBv0F1Tm70GoErFPWpWr
v9pvcoUbd/VinYTwrJPrxZzjy7SEwR5QhE7e+OUZrZrA80dS198hV3N7vYBc
JdpVJbXIweUkzm/qQJBXTfhjZWrxNe7cPvnA1fi5dnkRjf4NIEW+i6OWErRj
Wgox23wYuUPt0tsU9oOiol7A6bQhc0ZF0okz2DSjOuwk1P4vWwnmjmCuUx4d
xoTABMthX3xzuLsIN8aV2pceszOaWF0pV6F6mbtT/LCUKPsuY5zdRgqj3J1J
UIuVceLPdvvJOa5GicI7WUqmqP1tMSIMZHHNzK02g02E5xZl4cxnU5048Rle
B7U7EGlAPffZg7OjX4IcNe1Q1+vmwppSLvU1l0rgVxw3GTJZ6iYPoCu+U9XR
00cSfn0ul/uR/J0QFCnQejSfNfiN6sbIjuzbEWA8bxKtqtfQh16au+uIZtsH
H6OK/xMDq0iunSjjF9kT9brD8mknjvEUG3rAEf1+4q3BJQTv0T++vftCDk3u
Yn7iWHmfF65P/NmokWCCcnhQkoSvUFzTrUdhVAkx1rZX6m7bYrBycEhE0DLw
p5Ujafyskfyahur74v8A7J3UkcqXwQoMySUIdNN8RClSYdEOYj86+EWEIOPk
OsZ+IvPxvka0k4EoZVF0oldsdzli2QuzDLMRxqyqd1t8zBm1pGyT2EjnqUDc
riGRRhwH8brxrY0anzzcWhAGT5WcoZjM4BnaYu5mj66EMXkVc6slQGfthFg/
RUqnXHt+7PWkR/bUAUi4v157hJjQ1aA9AxLb14h3u0aoRo6GXUJiEcDRlR7n
KGPo6UpVGufKFAh33qfRmWF1uuUjhXuFolZDyvXnoX2vj6ePjN0aPPas0J9X
s8HOLSKQXplZlMrI9BvsOlxXksSmUqHHuVR6OF5lhEA6Qv5ISAbC/HRI6NOm
qVOg6vmVj5FVb15ATVZBArdCBDPb1iF9+bpoKzw8qeZlFJrW0Vls3+c/NTZx
DHR9deRg26A1/R8QRAZCg78GSa9eB6TVAvTTIqEcQosgRYvYHEiwjHyxnWr5
zqzfKrOySdvDLsDWgFtKtjvUKcv7XbQI5eIn72g8bmn21M0Y7zibstVgSIUg
wI7TARzsXyK+ygj/y427FyMHkXWWDi3WsMEybZkjsaLf4PA//SGtkVTnhpz+
6P1ADZKVEMPL+XFoQwiwQyUyh0J4owoM0222Ppv4qOeoumkO/Mxjy05iDZ/g
6ZZbDCPI0NYq5XulqKwQ4iUHcH68/czSW+A8t2EkQcS2vbdt9Sp3fPPMoAGw
fcFHhAzbqPblrWXXU9gxGlzgU2ftXl+OanVRxM0DiudH289Rwj4nn6zkakHb
ViiMLBMpn6HQbEkRFMVTGUc0am1q/j3vtX74zwMy3GuxGdk6Mw1/1V03m7Vm
4B2+zOM4ul17fdRVrMI1SgAjH3hIOxet2Z7ohWOTXXmH5znTjp9DekFHFbS2
6cPCMiurNochPRB8DY810IWchlLy8IabMrj674nJ+BO+2rEuAvKA3uOqaZsA
2CE6tkDaHfqrA4Pno5iJ+rck+TddoHmrKgdQTuy91WAs9yh3nkRS89qNIB0z
nRNVg7MFHNJSc2jr0EVaN0oXUNADaq1eNWEV3ckWOOwkpzcE2W744zPfTs40
kcZiBHx+akbd7n5ywNaq7Is7cUxXJrvXnOD9l5kQ+q/+VXZDyTcz82PjeOpx
5DJh0xaZpE2HcgQq2aov6PFM+2q1OW2jhEtyOYd4RkJkKXT4oDSUCtDl9g4S
nh9hClMk7nztvfOMDx5Ab9Sfs3uCY2NDHuLR7KrQbrZ0YRINblqaeKJi6Drt
mpQ75AQSt/Lfsko1gCBNDUOC0wEjTCHYjUAZd7bW3rQvBm91PWarVlCQw9wQ
JTQ0Bnmx7Gbfs+g/9go7UGytKHFgsZb1ElKY5gBDqCqDooynh4BoLElo/gl8
uMaxV+CJswOTEbaTGeVc85wA7mx+4VJc75cvk3XfQmllldkh6+RsYFnwrUMH
wZr2zUgHitFxtDiPTc0yhx+PAV5Vx6wPIEXMLuLzTFDpcZnZj8xQWys2YvxW
Uf6IqQTZnIL1kJsO1Ilv/+SRcXFTQm14ntdVAJXRVJXh3295+bcSFXAT2cR3
XibRI6t8dmRUF4q143o3kjr/ba/fv3UH8zWqwuS6OtUEkr8KXUG85xq090L2
0eZyq6NYhQFeaba7sXMVE3cMbUDLTr1n7FytRTfvfo0C2duUr6fhOiwgCbY+
v+7zoJLBMK6Xm7xBlWdwimEVqzpvzLut9f8sbC0eY3Ie8DuZc+fGKVkttbNC
6sSnrT70NmwikYrPk2EF08E2RAkEXJChTfwzkEgpMxbfBSDAm4cxIJ4qr+Aq
zswTePkhYTkVPKd2NlK52D2snMY5mhTuXXdd/j1AEtpe3FOGmZKGRiBfSM1L
8yjUbQ2VPgqnm4owZFMAl6mYpPF9qQTTHp60dtTNpX0NNKKKoH9mTitG7PeR
S9bB3LpHZrl3X5Fk44FPZcTwIoO9Z+gkWACB8YjzaSI6r/A0Wxun1Bb5FxFI
66RmPgPiftxZBY47Rx95wESFJtIaa7HX+oacCzYrehP8acll/Qm/ODiu9eFZ
HAlJvyNGbET/TK8bQLjVoxDm2T6m3oyoKiLoY2ksBPXbVf/poj7armUg1QnB
HChRdIUCMjR378LE520WM7bsq05mpT2WB6M7oKntE3MOfrgxUoqdFIglcCjd
jpBDAtDKuxqTKkxn76p4qDeQs2wOVHV2cH31I+MwHBWO8bttkcVIKL6egVJE
rnQ/adNZ6HaYkwSta/8c41xjD54HMaO40+trNSQv90QzW7MVK3fYJSUhrGyk
xNgghx4JmQKpxfnP1hgd9k9E0ioocFd6hqTdsU/ap77vriePXGDm8nwoXJVo
8lOYt7n4SKuY2Jl6MKoxoW0D3AaMdXbtrvn6TfLRqPhD4EasCVsi1JIj55E7
dQd1GN6iIiBK/jFRMp+rclEplqfngbxrfyO79gOTSe8LJm4y96Cf5chSt+kP
L3Y7aHTlqpZoTahnq4Plmv/xH1+I23RtQKyqZ2FBL3didDebs8o7aA6EOnU/
YtEnfLrW/cRnN1Ehtkm+1kFPNNFBiflTug8HxTbKTDluG58f7rxmb/i3jNH9
m2rOH6UACJiCNiDJjhm45IoYBE9fLMTdCrCqNJkDu71Q3aZHzJwgft6SFf2K
Ou2v9gDpkuOPLh8Ebpj3uwj44sH5a8873QW9/Rmhn6zqh/iGNc5GpitlN8na
xqQ6+BuH/r5Rsfc4LhkoZM8uwx/E7HxDyRV4EF/x5TWkyvx++o2wkXmqfDOP
fM347fggMyCEJizmmHBuTPYvFwbNgFfJ3A8ibShi9ijK+kA8zXYruj+ZHBYW
X4pzOiRh8waPAKp7gtgkGtCi+mOh3LG7xmbuf+gLpUSIX3YWsykrsb6qiblC
kTE8NsI2yVa1UrpyB8plXA3BKlDp6JUh6lAi8kQC6g3Mjo9h1YIMQdJIIp6n
fKIiW5ck0Eq+xetXCjg/2fK30BASihDEA5f3/jsKdLKh2pgsH/AmSrV8Crnk
TB+35Q/nJawMqXC+/+x+UWkp5kD8J/mKKWA4POhoUoFM98pw2B54YW4X4PNu
erlKqeQ+kB2gBXvqo9HbfbRStsZfz48T6lMf1K2M9lF0QztAg7oHCe7WQmZn
KLDC18P79ZO1tdll7sMbBxIMC3lyYMsBgaVB+0ySjpK7RXrxP5Em2CPUeqiF
kOnZn9NiX24gpOTS6pvGEgRr93sHYhz5ZrkMHNYyRDsBJE2X01xd1NLEkNja
qCtnfMMUZe8XMdxSMFog315IB15sM43H1MAGuaRKnnXI2P7SKDqijgE5VWLs
+h2TJZE8AmfuIlbB18+k7alqXgnFJAoFp9c7hHUw+Ucbu6yfuiSnwQxa2bGd
693wTUUFm3JKB7evXOvKayrmN8KeLuKHucz/VQID9nZE8Dgbylgle+UP9LWq
2TQLQ4jNc2XzUQqW/f/WEpseoK/C7qRJzuE+HqW0ca+esN19cOPWQ8JojqgR
Hy6s15g9TSL/8W9FZANiwLvgzWcO1YkpO37hYyH7KNtrxuQHeBjXFBNbGF9g
l8EJA84AJIy+rD6R0RV4Qc79iFWNBUZJ1A/DNyry8nAFnt9uKrv8C0tWUn/l
6m0aJiy477UyL5Qca/b8yEi/3swbYvOvWE/Y7+jyab75Ayw9bO18zAAdfSOa
u+eIVIUGmkGuqoQ0wsy/BM5pqOtKGwGZ4gQjV3pDkokXFeKj0rCr0PtOCnFj
zsW6raCfVjETBmJUySpwBrFg8G83wmcz9eYs1HPlcumJl1MBLnJG9uwp2Bh/
hS3hScIL4Pg/uc39cDzU4+IQCOVAxa+nUZFpNuUSalc9xN9C9qDFdVVOnSHc
f8BmAxPjIJDFZaXXsVVuPo1dLZruDS8VzISad14bbHQlPi0OQvaHuAj3eHPq
0Ks4VxiEl093jzndcm5d2LJnCrZdOntGf7KoaJt8Hs/ixTyc1Mn+LQ8JSrxb
QqmVZDS0HS/AUSo0GwjsqwmddbgWJSM7+WRAU+aqL3plAcFcDTp4AbY6Kaxy
M4JkTXS3sCRx4psCZhEkgJmQv3FSSzeygupAYCy5RYLBEXaK+fah4IQgTadu
jCPs6vDc1l/6vXk4WtfRb89rk28NcJN/eECbq2pjiYOyjdSviErk8mh7bpyz
2VVeX9jMxkLpt4pJA/mR+eoBTO6bvQVIyP4HS+Ol8Q62F2n638NhoKEdP6M9
MHsGPuSHewQfhX8FmWC+Qhr8TLBl2bTdiE8fgkLWvtwylxg7z4NaGDLxWJDG
wrlwHea2CU1j0V2/N1gxhxd9T/OrekStTovJCZORwi3haq4UmkZEVPPlnt67
fSBct6UQeKP+ClncT2T6NTGghSV5veAe4qdd/YWnLa6R8GsE9VSVxZHLzSWq
8yly0gAbEOxqo9GN0NMsxI7jhHd7C7m6NprRtK2ghGLrWtodGGGGh5gVoM37
MhcRCxwLuKR2gNnUv5i3lrCbOM8FXHJ9Jq21eE+xonnGorEHw6elNbd4gmHI
nopDh8niSG6WgRPrsQNgEhGHJH1a9LUGhavv3i1c8PiWCroEkQyzsmtIEBYM
Hz2wVXmAu7pqOE54CYkMNm2QqAecr9cZ821A62ARu+vhmRT1Kx8VTb+bHtx2
o9vQ8FwrHD6ZsuVWjHA6sFVxu41YuhG2DVBiFsXRRjxAuCt+PjfyhaoCSiA0
jX3LRpC6HFp86qr7vqIsssrXpwrJDJk86505X/0wqoDBaGRVniCEM0pZgRpI
yHmivsib7w5NPbn1Dscbob478zOAFyUudHr+CbzogXJn6DqAtSYKfw9jOqTD
ySt42IWEVNFVQj/+d5lzXM5DeYysNdkRdD9H62TjctY6QZxJgSVJT4jJZzNf
pC1HTEkHtjWwAH7pkGaS33NCeT42hESBy9SDf7AqJFf6iDsYnkkIxNU37tix
kSAeVnsPLyyIkhkSxYLWjpzFMs438eRH8CCnRCNGnzpeABwQqmo4sGXHSCXQ
/9cLg8foEPOQuy+rOFNuxH/CHfB3trBzhEICyuCe76Uj3MToeBZ7jgt0ECbd
3n1Ix4INXmf5NI0FcPKh9Pc1jQ4kkuPyNbv+NbrI/rZ9VsNQoNJjqAU/MckT
1FKufSsV2dRmYHdSlJ3v+4cM0owcPtRlbjR0mpXu5Mxa2Ax7ycwA6AJqLdWZ
rqnwxHA0XYcYIf6aO0bllb9pGcvYHUUets4OGX2wm34L2MiYbIJ1Js4yQOs4
8udVc8RVK0cQmvRBFtFbur1du94ATtW0o1eogOy+O2o5LDZwF9na3PpoOWuT
vBwecDVX3ZX6E+a36Q1Rf32G6HKnB3WTr+MArfgF7/FY7HEMOzpoqWftRzoO
CNkWkD8cnZJ/9ytJkCPvzewG5/q6Ft6RZX/2LdZLQaDP+BEGD8+h9W8iAegv
JrxzveUBtMyNAwQDHrkqnFbn/VCdLSfq20U8FiMVkbgsBwoMgYMMmd4Xrfbs
S+/XvIab7N1kCl96c32r7hrCwRDf/K9tvtZlvep8M+4a9VZliGTddInEr6EL
K03HmRTfrP4WjernhEBsuxV17jUL80cruzrn+WJrJBggeJ1aiWGwvh3JYVtd
wIIhRK554CVWeKy8FU8QXw9Ltt45bPLDgL4uTr8R/LkUKcP0ftqcZMjtKTYd
Tcvsfu8Rz2ixUzx7JUMIGGbeN+ntOx7ab4asyx8JtDP0sLcCPpz88eFtAbVH
hwBjZUCopYi9q1KDj34sFuf95B9nZt6qglksmTZb8mjDtgJsIOb+UJA2iVh9
Vhx0R+BOe+j39dX3vewR/Oodl0SjBmNTVWPw9klhhICSqlYfMNUz0bZBe3fG
Kiil9sde5KJ4wea7+FlpktdCrbirxlO6W88mP5wiAsmtRCYDMIUSlP2SK1J4
ZetueogrrQMDzsWaBCuWhinRf8qapMsKZg8ct5RTyfecx76ZMlOQNEdf7xm+
8QzGx1I+AhKgOnXfGBQdgZTdKU32LdC9vqKW9YoagQ/J/0LO14+cCFzbvvCp
m0QzsbzifGAOMBYcY5JZeQe7vnjhQ8+tVn4RI17hkAdB3I6/uA5U+qnw2Sbj
4vPPthgreHgQakpRjNMgnKeYcgDgiH3lB+Zq9FxGH30r9Bklo26RUu5IS9Cs
g2Oz255LGbjS5wucuJqggc5ZZiZXShX2f1wZBBetvTMFd5HD0om0JjKoBdk7
N9SNYQ4WyQ0I9pWMR1EJEZ5ck5YkbTvkM8HQGQACE7KNOV/3Fr+/5XMhIJzK
Os7TiN5RDenO/EbeA5uxn5o8joGx6h5ZIJ7cDMTBhrSmkiT85WVCfWkP2nq2
xuqpOygSjY65lUj+LCenMTsG8drh1EX6tHXY7V2Albm183QyIeFcR/eIMge5
YSmBB3xMWEAibs7UcDLMQ1OajCHmXPY26QmdwHN+zvjcDe0FETTicDiE11TE
35lIzxV/1r3SPGRr22HbQX5p8cCZV7fWJ3f2fh/J1C24yCKk2fD+YVLXAAFM
fwCNImhcCwopgOgyLgfx3ZI8ujhES8gccwu3ZEOuYbX6DTa2pxTEK3cC1/xH
rYWR3rg1PFjNbIMGoC6DYEwfhJUknFq8yZ4TIT1KdEZfCT4ICkgtfJJnX/p7
5S1RDj7dysn8go/v4zkgctP7SCRRe97F28nzm4M9HWMwz611GoNzg3BVY9lz
vScATWHHsR90U9LAssG8Jvp8em4S0Q2Vym9DeEfdf0UXawWj5jLlZpGmM2I1
w2vgpYgGRxemn4raehBCL+snIl4QxX3qmEo0TyOZTXcOzaHm3AWHFCA6UXuu
k0QJxYCFToPTJ5AiuhTD4epz628z0G1y6MPbrPVKofAHle8LnCjRkgSMKROa
qFE8xSPcOZMDFK6RX9JIWp1wD6JLVtuonlgz6gp1u57J2iwsLXCJkE8saY9o
ctm+vskavZOChOwu1ytSfx9+cE+8BMdaETccHQUUxx+rNjPlEorHeehBeHiJ
q8X9E8lWDFe/KtxtNFBuR3PMk8qBnJKyRu3xL6TOrslCkPDsM2WnRw8/wsrY
La8KTooochLF5isoZMeXclS4FFtH42UyZGYHvU2hiVbWkz5MXWA18t4CAMi6
z24MGnE3FJ2d/HDclzQ/PmKHz0ok5w8g3mLlRJkdEbn+3ScpNHRYv1jWlrIm
fHPLx3A4I79X5RmEPWOQ8U9pgHAGfr6zZzr0iXKBANY5oRqGGwWCQfUSMoht
VQq9LDFrcVzli1/mOTfCbWoX4wLPQDzLUdtfqHBjA0MyCaHuzs+AI2XcauwH
/1sWV0+yNKWBZz/BPZ5sp1+wsbjHmGVCZOeGLgDkAPDpwsNTk3EnYntmnrup
Zpx1ulfyvGg7hXHz2xYUrRU7RV0GWf3hJh2CXI3VqUw0+pC3aG2/n1p1ekgN
V/ovFqTHLI52hPqKZHbDj1fYiBTmyuYlgVTKSlslIgCzeRESCqShFDIwU7yB
kTnOUXLsZ4oUDZevdWL6sFLi8pwOkDEYwzBjedWnnxsYlpkiqHBjExCm8EbR
IiYDPNIEt8o3sTK6sZCZYl49qUEBce3ZDjV8JQBZSBes+bvf/xNZ+5ID04h3
3XGGS7enQA0t4y8k1dxDk5aBKlla0CPNq09rPH+CxDOlFXKvwr2r/XeKlvua
G0djQkNF/uxJsnxMCrG8Eak475Qzt3KM5K4Et38Zkplt66ODCd/LgIx3HrTv
RwvEfwbdrz5/yGUyCDTnx4QvApw46pj6HZP5UKF6NAv2Icp/KyOkNFkSkycJ
/E4zcG5RS3qd40QKv1tiXU6T3f1d87UOjlMwWVDFs80+89P+sqdX9gZ9rieU
08xLHRCfV7Ruwj+VpRsVCj2JKv5KR++n9zYMDdRVWruOJh0XMH64SpzqHxpL
BVMd1hcweAn7UOHo6NsthxOHxvXJy+6JIurXB9Mw4USqhmQBij0Vu+CzcVcc
WmjqOe0IN8Y4mYDu/OR/V75kkYvrXgSgvkjneoM3WawLW63TI+YxySfm6xvj
9wyvt/AT8O02fj7ucAHoqj7d9R9JYJKp/s3VoAw51sX4eSd2SgO246vYjVtX
21Ck0qc1cydg2a5+g7glimEMJTULozpfrLPL8qwaNEhA2roMkr+8Ur1+i4Y5
9f5trZSwRM8cg6ELwIQLNtTO9D/R93EcidvDPqtZfOWChhpT+ma1AB4hqZA5
v4juCyeV7aOiIL8NlUNSWzPJi1B9mc5OzJmj6Aym5F9DTV7qPQEqqEWdQ40/
JVDdnDbL1oTMLzd+QEWTpV2uzTIFXrdgcI/rUlqJrPpngJS+pC22LhskIf/Z
T3KCetHQgcfQ7GwwFL3Q0nye423KZ9eVMyTGnaCtOZslFZcGc/t1JZA2YhNG
s+Wcgyeb1FDV9clkxNBOsDmXFwPHdRziHfuF8W1YZ8S8y+ms/hqcwZNCNbMG
3O2Ei/YF6c0rE7QDlxl2qHAzXvBlR42TMrA+/8713fA7OrIAT/CO/JdQc+ZH
PCFXf+vpS/Z0ZrDdJGEcHU9+gVqtVsc9+4O3ICfjf90AG5r9wbWpr1B++/VW
BCizr1WnOKm6p/iKiErkXvTHt39qbrYSfYAytQvz8bq5ueUwNn1hNr7k6NTT
6bV/ZNFMg7kFnbpFV4HUG8IyvzmZ+FRKugwOf4HVDlbp7Roq/DzIpCf+xxeh
MLo55HKVyA7j4REU5ka3sqSPQSNwCl31n9UOJBxxNA3NksYWqU4kVjqiTkWL
bhyO3KEv7gXU8Suzr5HxE9oyS3EyZs7Mq9vTj0gE+ubFemqcCfKJpWrWBdNs
ANVcGzFOiJ6A4LJC+7ca/ysu3No8HCLAq5akkpcNBcZefYk4z2Nei+E6yAel
Sc+MV6htVylD+cFnVSJXK7+ojZFRX0yLTeAUkywMdRnZ+UBwRPKaw3urHlJO
dRomDCyLgOlkbM8d2DQiOK5S6S2oXtWjWikHjQwe8B5n43O0i4nfKQ2QYVaI
eHme7bQv1R8KbhKo2F39X1alHpU3Q3tkdXi2S4KZxk4EKnMJLOqzB0gS08nY
bugX7+tdni1bQ7pMgObDx9j82nTmw2qJdbj07YimNfMjuJYYDwtmg3Ylf9+S
zd5pFhd95pjX8LpH5SlyW1wSxOU+UsnNRMN296+C9fjfOVQqsOw0Cs3DhF3R
GM4U4ZE9MdRpdhVgw3+kSRnbL84nnYbRBvRQVqy6YVCgzax54lkBmtMV6VG8
qqklpKuonYdEXOyao63KfDRmYtAa+94OTpht+RDtodTXQFA/jAmeP5nvKEcc
qyo6dwHlk5t3zARkP7b75Dy/Ki3INAALeL5abqZtGZfVdBRmFjdq32OgBNrb
0f6kqvA+SIoDgI6oMECrByBjawqx6PH8Dq+FkjIVoW42CFcoQ5x+kx7Mvjw/
jNkGH5Sq9KPFn/Xunut7uf1GpG5Pe9cdDiB++IsdtKTvojvjCTjsQtgSYqTy
IALS+Wa8zFB9nHQky4cP7msEERF9qZlEmWtsHGM++4X1qrAT4jJaRbDZNcZC
cgCpPXn3L/+KqFgFuoAvAw+cHGfwQ340/m8C8quDQBut9enJIxjQP/q+oGau
niDIhtrZ9zhuRYaDCsfMpy45g0OqUrYJ4CYB17xw76RXmd8PGJ/XpqT0CFU1
FXReZWzImpsmkmpf2LL5NzmswejGgrmTQ1xOv23e7Fzdk9fz1axgI1efAFg4
1EdvpOpr+6VfpvsOfp9utIqwox0zLyD0G91YNYnR8vc+KqT+iEd5uHnpwp3C
K8f08UO4zgT36YJSNdK1u/KlI6uOIxYT5Rkx8e/YRD63zPRDjdFP0fmBtLPh
BEfZgFKvVsr/TH7dEpMGa5oPYHe0A3UAJHvVUUGyQlzPL0z3fAnAFpb7spmy
rx4G/n2gN/wzb41E4ltIeEXFzR/Tubfej0TvrctYW+Q5Fh2HSHwOReOWCG1Y
/IMldvxailwPYaxN53fVhhd1re+QWgiFst616ce6OHKCfA7ALBOGU1InttL2
yBrQGwV4pJ59FfSKiSdEg4xRSYK0E2HgwcB8HyvkWaMgwH1AM2sOke/BBse5
vdT5lnQZzSFNdRdl1lEqLNdUHVT/Mv7V6ZWQ4kP4N8xbwGNzEVD9Gbspomb/
dGn1eQ+ftmTm6h/j/FpJGQRq9s0uJOmixlFI+YHFi39b6KdyFGAUlVyt9IUb
iDbzicy94mnofiFrf0yXb6GuslmPcnvRfqia8CWX2in0ZfvNG/2jpoJbs34C
IkFr2XP5gZEKG+Q12+YijxjcLbBGyTOBIXHe+geIk4SHu0Ss5/Zvm8vS62x3
EcV0LpsHWDmUWavnQtyY03uKWhMGvz84YNoeEu2ERS42stTZkCLifNf8i/w1
dm9lz75jn+1oKbj6f+O/sYClgV54FTIhogKY8Q8ARI7ZYKmJ/JCby6kIkSkF
1kgVMqL4L8zjT8jbfR800/lZGAsNwWFfI1FRNEmm0WUMI1NkJwfRURZEqsH1
qFq4k9drOWSKbI04mNUQjcH8bKB8PbmNvXUgT9dcawzrrVtP1djFfiCCEuEi
f3hW4ktxXz0ObBNLu8rpigOxNzDqNBEb6D+G6PmzBNC6WSR8kxfOG9UNg7xs
5wLMey4KJFO9eju4tK6IZq63LaJMd3M9fdPZs4PcSO/wcTuJzcj5r1IoAeQy
RacDd4nsGKthF22ZwuPJpMSHJDuipKIdV+94dGsvqmxkzmQMzXzy3pWCvZci
ZccN24VY4duXnCd7Y8d6RUbX6i+b8F8v7LnI7a9a9ltHeIxjPaXsOj2oBIgW
mQZMpQ3RYRPGorLjxYhzwTdXoT8LOGnaGzmmJvac4yIB23bjXjqN1vQ1Iqa3
bbYjj4TxHz6QzzOA6dLjzqJq4Z1j0L8EBdchZlQ9drWo5CUyhSSaOSOvTPhk
ckxw+tFBYp5TLasQd+0/7e25oCvJ+GmeJhVZfLmbP8Fq6rAOKELh+yIYDRE7
bIhVliFQOtE/goZbp2FjxBLEu2bLXPtP2TzRnuJQO28rXakSCvJcw0i65CjI
8IFfTLPp/edaX4dyBiFELEnfZeFdUicWGS9VOVAeRzalqcSVVLRuYe9eFw2r
0k2qSNo23dJmd/lJNSuARncMHE4FkH1GjWJ+rp/mkUnAOY5kQF+Q0lHusjts
pedSC6MbXlGIY3WMYZs5UhKjjgGS76mwD51mkUgN+1uRPF+AfFdcMSXDSPG+
APGYIbhym2TrNRNfk8YMD5dYVfFApN2dwe+zqYzv03JdF89uDbPP50vHI7JX
ldDLm+OmUIZrIBAD3IY4RrCYI60PMqH+hVbEvNdW6En0vPpYOQccbuh70/qR
UBK5SW6yGxkzvytNNsNcUcIq5WpJ3g92j9p1RLGimhcT969s1EE0rzwvWR0H
Ia6F3fG2RtjdMpqeEsOoALmPEU07ubNxs9EjQEbKy5/cFjBdBaEMOOP7cpbS
JCVIYmD5uHp/MkSmcijdjJrNriBrQsJUgw2+NAikp843QvqE861hpTvdtGEw
yaISD2bCRoYwF98ESmud9HVYkYPpOo3jVYb/ulU4Ast8PA5IGIxnKd/1pSEv
2UFIgAvC7GhEj8dswybljD3Fx/xXnWoyxqzyOVqXHL1XD9VSBA6iulzq+Zrx
0fp0L9K7bmgAl6EGoAkvxN9SyD+PX6NlSZTkBeu5xVhnM8NR0vtMAFpRgPky
xFi4ZpjGzujSLh7wqYAs3yIAG6ryLzOpeE/D4b2vGrgwjdLTv6rL3XE+bYS3
L76fAFGKTzSjg1xjfYQEqtAIV8mZ6wNw02Onur7MKNMoRD5WHTl53JAGlXSl
bB3hxCpr2tMU9MMOx8hWV1+4i46vBHFnN8y5bz6AnXydS5yvfwHyyJo6BXLz
HnJaL0aHEpuNxxf7q9K8jJh0e11zxA9rbYPFCAI1syavcAsvIEq+Z66cNyku
c41OH7AKsk2gWqIRSZGl5A/+2GO5ckocex1MtxGgldMCxFMtcH8S74l0aXKS
R2w5UQYM/ejPe3V/pov1fXeM40jE/t/FEC7XF39hL05EtS+MNhY6eyA4pR5z
R+kBB5+PDeIcHZEJunYi4DZY2o2eYQezE8b0K5WYsSzRnfaXLj5YMRLpWp2n
XZ+cCHYCjqeoz/8C+1J/hd/lFwEphh4FJt0eYEcXo7s/WKsMLItdOFOTeOWH
YW8/r4FL2LoVzAROHSZbNUlb4pB2r93YrrGd2lhhogRdE/vTfSOO3TaXfu7S
vW1Bjgp1H2ySNmi24M9rgDsdjAqgZP7kSApQKXDdPnzpxz0gfz313WrCaMYU
N/JbsGBK+zUg3kVbeEDYTRsy29NP9JaMPTcMBLksLhFveY46i8zHqbOrVpQD
hA7VH0wileivRrIypSV/0zdV4T4hnCHxpKBvhx+HyheDlQvCFpcQ4TX/kihU
qjD9jkw1YT67dJlJlmMePcxig0axEHmjbsBSTHPG0Jw2MrNFQiEeKWxqaGhg
NC3lQ8Uo787Np8EOTh/4gB9Y2sZc64tPq74DxuTkpq7Aub8RIdu8xkvWQ4Vp
b6Sdya2G92IhahvruFKqBR1b76iGpywMD7djJrKV14ikGnQq7aJtJqgegc7P
BRPDanvDIrgdyPMHmD0mnT/FF6m+SZJ/ZOE/oP3iggb97zOnfUrmDMRDMOo+
KYzKdfeSgOALmaRZPj01/udFvYVjNh0xUr5aDBWBFILquXXTxiE6ZGt7DkSE
egF3B5irxgks5TDBCGBu1RG02huhnDI6LLvn7la3nwR//9W517YYc6U7mnE8
rlmOeH2IS0i4dpfqDk9+PYh2IMb0hKQLIA/tV0JBCwzZqNu1Xl1oxLkxEozp
rONZT11cVLolBCT57lMIP3bqT2rQlF0YVtQkm66mG364NKiv+PsOoLXe14Qd
UONpFR26AT0gMhiO/WB8gTM+shLGs7QDuO47WkqZHeliVmqHeu5PLOxZCGYN
H52LesxhiEEsrbMgGFLorJ/fSCqgkPZ1cZGcJ/t4byyp0ovMC3nGsfABKAtf
uvazz/OThHFv+55ZX9DlOIZhNdprncYgFLq6OLE+qi1fCGnLKu8OVcZEy5Xw
5rsRItmded1eIV3ZdCTNzwGtY1+0o1ZoTWMwYO9tRDOpDnJWNnIJGxMORxn8
Pft5wJrjSdp0XEaALxwQtVbQoRdzBeP6RlU68UUx46crgb3rVr+nal879CBv
4peAYsQZhAiLtoG0932R9LRBbHy/eCKYPAkWYPkDDBRPOmQ9h//58aeKPr7o
kOig8ScGcBfHdiOAOMrBUM7CZ9eR7s1x72b+cJMCxF/LiMiog7GF6TWS4hNu
6jFyu5I2WubLfm7EuZcg7K1mnyVsE/UxRIy2bQ2RjWuUPLVCEsjMAya4URif
Q21qad2sGVNxhrS72C0utIgnqj2uHclGkVeEaeTxrxaqbkv42w306CH0c6Dv
9TF508nKdgozSbgMp6jHp8ozGuTC36rKQzFtAMVZlhV0/1hz1U55e5BpGDb3
+XHPYpmzSx0CVWVWMR6b1AwFDiNtDdTC8Qqq9CgWyEfub8dDfKSmmjEXsxhs
M7/yIUW6yTB0uLHuWnMrRZjgB4bKzEOzVZXszasou7Ys0KCMz2cNzhAQrnt2
8DGj3CcjOh+xTOfBGNcmN3Odq4xJbYwYyu9Hoa9ll3FPeXeFsbc93/HYaoX3
L6HiVQvDwPuGl5w0r0ZCm1L4C4qtoe7p40lDP3nVWIMFEwwF8TI8bLAs4Ybu
pcIdHJQyCzmt5m0FAXbt/ak7LrYGi9CiCnTRRQcq/nSe6SCRyn2/N7begIj2
03VG0qcYuJq/XH9I7C4NFeNkv060FzbyNy6uHv64ffOLtaIkI7Xfs371K9y6
MQhd7A6huBRAKYymRw328Ywo4Bo298HzGhRCEyCGBV+X/DD4oXoudjFTqUmy
SkWcqpb4QtXSx5Ia53fnm1GZfY0m64xOYcBDT5AIxV9+J0lzkJfjbTmdQxCu
yheyUUvJQp8/NT/x0K6wbeqOjftk/F4+8fRRMAE6qTO/r6V85dpWJhIZBDzZ
6i9LBxssoJ5Y1dod1cmfgvw69hmEG5bzEr8OUVt8e4yWUPPSekaPdetdV+OJ
Pb6PkC5jRnRbgBAk//XZKiOi5X9NsWoR/ujfFszKIhco4JRRdm/iUfWY+rrH
q2TzqXO1wQ5+xdYHd35WLsEBA66DX6CyJ/MdPa7ojZPD/xgpQBS4C0SsxB5B
0rz3sur3SUWxxXIA54gCMhGPnT7LZEseBht40yaPNRYda6sH71PeN2OO89K4
6zTRBPF282V2MqKq090oE5WH8j4OVbIGBHmEAO9FfpRgwvfnrvzkoeDFpe1u
rApZgfq0EF6o3gVqjyHDoRMBtLzsIyy9iQOBMu33bpjT+1RSiiy6zSQqQhL2
2YJcS2g26vgBGgpY3uKJf0Z2mmIct0HRIwJjBFH47/wdjHURClCtYWxoh/yJ
qvVqz5HUeH/jTYcUoHk3XttAJPl3IZkIh2EN6axQeuV8O2pxra3VZD11cuCM
9u7TKBXUiem0aNtGvPy/ZKcjyOJSBJ3Zc0XUFei+V8Ds8Bcz/GSfMk9xYnNW
kWugimFdFoowjb9bAHh9cXX0MGhGTRHh4i0VI4HY99xFZysmh0KjISzPj3AP
5Z/oBybKQywVbdZiAttQUfXu8wk8g4N6Wg/RwNHmZb+HTWRZ+NuZkErfXtvw
3GZIqh3F2ylVyYKS7hT0/tBNaGPUxtSMShdgtPkT7a10q2NrOjFJpy/yG+Xg
FpkSGO8LV52RTqNTDC1nrZKSr3o4FJBodOQ0xRNlka2SeKRkuezq9USNof2H
NbMbqTReNRwsDG3C0rInq+qqVNeK3Y94AMSroPvI+4Yg7llgPDH3qnRPMn8A
/pDBZXdgpjLphVRHIDidx7oHnSM4ARMtGBgItzR3YsBHd0qb34tn+RqNS9L/
/ULI2QQvRLIgeiBM2kFKBb0ytVPY6jywQtShAYlkXNNuwCDPdLlLz3P2PQ6g
rTjGjJZo/OgKfk14LKqc+hFhQ/LcPa/FCQE3HiWXu8+rCgMcF1MBOJ0BAFTJ
qFEsUwwvUBdtZpXT3HFMldMI0Q6ukSmoPY7Jd35gr+Reypw1Qe/wDPwcAJZK
R0H8zVQ3kUaih1OyCZJ/mekM9B6HGWtLsJxg1Bnf6LoluFwqzFfqc2nGCMPD
5q6EompYfatkJAu2lWYBxiTHS8PYfZmK4Ata0+Kaey0AFrAMEsRv3yIy1UIx
9oVBDls/zI5kLLyecP2WZvXkgtYspYqhDcmleIXFXXQBk07l98jHkdVRgm0+
N9L6as8sgTJwa4o5TRb3CjADVbFt/MDvy4sCEnvMShMUH/qaQ5Nwvj80Doma
SCDcATQjb+8+eJB9hm25ZvghOtS9UMdgYdWiun6A+EuVzfiM3ybKxwOe+Nma
H9u3nZPt8jdVyzDWlK5zAi4FKfR4Qb7hAUDVIBleqoIu+s5CNrKwP4E+u0/R
qpUvy8KwL4xSKIUp3/117Eza3HwXZhdMk1jYCtrgrCNgXOHJ7m79DkMeg+LF
XTWK1sC9VwdLYn1zLCyiho0dv3wBEQ26aXMBSyYqDjZpws7RxkqgM9T7P7W6
ftrAs7nmPOOUWiqq+8wAstjTONiUna6CBuo2hTyVgMlJamNrfK1rZLKIP3oa
U4XE7T1EEeuQnmPDQpn4YQ5Q/8XAGzGhNs4VRR7djJKlZGC+OpoJO2u/Xikw
XOIrJvGF9seDJUnYnlH4jvrr6lHOhRnDPaTb1avL5BhZ7X9tjz4lv33d2YnY
i//gM6kouQC6Lk0QrSIkITFJTTV+gvezDZucCdxF4dApwXouzgoyBdL1+4ip
J/Oh2cA/1o9TwnAQS8EW5FQ+KXtrlnave+/s3NmiwKGzWxUsUM5CZ7RazoAW
pQDWc05k/eJlg5O/roGek8yd+KdLGuJ5dUx/0DnRIZDth5nv/ta196IunpVu
2w+Y7DdBTfcU6JtuSsaFZX9Wuy8lruChLSeTdD+ssJ4sw7KXuAU7k13lLsXW
CQzdbFDMvmWjlAFZNyAuDGKAmDlxSkSnNqqUfn6TVgWwD+E3LkTmKG4wYxcZ
TtMtV0YrZLqxiKMcOG+RwufRXT+GdtHLg4fRohZehibU0S/Bu2m/Fvj8syXI
l/HSMebdC1qJRTICyl9wiFAyl6TskeMFN1+YDofdV6bYmhmOA0nb3rGPSqzc
QuCkPaKHXHp6Vjd2RXxIVzJTspLcDG61wO1qp3a9qMsTozRnkTlf7p+d/GEs
z7LWghVqClbRCy+Y3eEyr4OXZOkUaYC0mZ18jcd0E9vXnDgIB4atgv8Sxb+d
earDSxH4f6Zk5CVUCCqqtne1VyaHOJMFJCYk8Ivi4vlUPL5MbfDgQjGj7hVr
Xxx13QCx6xHLBFB+6W1IfhPsD6iH04gVrEJeaUL0zZ/9bHjjsZdSyxcHnKvi
t11ADkdMaTT0NpKtTOJYXY0cgYGUw9ssSh4BuuoWCgbc8+Rn8URbxWuy90fg
VHEav+bxGkZLbL9mLQgcxpQ8mobNockDvayHsu+VkAS5xxsumE3vP3g7094H
lVfsVYqV0bs+KAYaAN0dbEQ3lWTs1P1XjPq7JBH+FZGtQXaktqxIN768+mYY
DuESYuWofzRsAr+Ci8mugRFa5leyLy93SW4m1UJFHvWEXEAPfeTEtTX6aGiX
ibOuOPIBV9MtIVSrzybPtG9zuR6eJoS675yu5VluezTzojH06RNN5bSTrcYU
6lnsM55zGQ24q4L3u29r8qAeCBHoVEfNvuWVA16F2Lqb0BBvZAp/JAi6n5gU
QTOvYEbOXBnijvN4r8aP4tUyqlRw5P2//g8536yv9SJg76dCpAWmz9F9Q5ij
nyxISvhCtnWr3xim/pk0EbB4Sdc1ZIa1NG/kBbCXE5K52NgL3Bu5yH0aBeuw
TUD18bKNMVBbhLiDasiXQU7x8MUkMV+CZajTnArX+L/tKP2/PWxthn8lYyIA
JAclFGY1j0j6v6IZYT3O20tsVCMaWwZ0jEBxb9eMwWdRAIvx7bpgxWyCwXnL
6AccMabOI0ArSi2qzLKWzKQgct2bfLW15YYUfgVGLI/Dlx5rSWTaDEp8TZBx
fpY/LyzZMklS1oEr5776jpApYZotOhIdJMLYu57RuiGqva9y9pv1JgAtyrRO
OhukQ48ZUxQUNuQwT7drXu3ZcP/HV+Y36abWzIzlSC7sH28vyD/Fdhcj2ql9
Eag3S2UWe70BR0RgTJqD3tWVWznReyOKemFClNxRx5usq3zKt6q2bk0Xy9q6
xPlN5lCH4vJfkcpesbnWd/l06bC+EzJlctdl6/kNpRTNzlHbC32eyfsTmfU0
4MvzZ1eSmogrRfS2p+1E2M0CXI9R6zuNUUHX3jj9oylP5qA2BcUsjhMxZjta
JXVOUpBCKzbEiqldiKqHHpAuOCX2WCYfUIJV68NaS/sgXauDVLbExxuozMa9
j5lViYBpY1/TrofLyt5cI1t3BquMbYf+PIpBQHEcKw/eZy1VXvAKs/2T1/Dq
EH7vEiTBwFdixAIs5XDJByPk4cOm/h631GqeaOjhdTVx39Vfr/eT6h7vEyzu
7NeGkgr7hrRaqdlMemTkYwu45EUouSJe7SdxoOYzOtKYbOmTHsuCG7Uh0Ksp
7K1VKWjvLzfAfUUgfziUe7NpFOItPzzgIS04iEMdKt7/wfvoeDfM32drOdvP
BwGEHl/aI1WqsaPqypuTozRk89Saj6Bhbqqgtw3+gVPtFXECfluwzOYzVG67
ZpcwYYDNdR0ah0+7b25qI530X31d4PhjI32CWp6R2h/fqbFv4OGxvKoY8844
2nOsDwzPoUeiKyAGdOJwb4672d924Iuh9mr153AhXOhZHcTXXULkAshAiBed
vFhTI8P5ug9ud4WzXRxDSQqTpMyTAB+anccM3hcI9twKcacQKfwIUzXhJa1Y
bmVGa8MN7Q+Kts/Fjjf0faQF5TRM0lRwiJgtTjrT/n4xfoa3lWPn87YP+FiA
CC849hcd0qMTwSltMEZXWckLWnJpoEIj3IjUz853S0Kp0vCw1zx0DiwZxuT1
f0wxcVdq9+XLppErpun+Rbkflrturt2fPMYburbcjBFZLqW2JSCikWZ0VTzg
+jMx5ju4Jb2xZq+MAg6ev2WjJjizxjkR2gbNr3PXbG+bl3cYZGyREVeNm0cQ
F6PO2y75yyFA4Pecvl5pBNgU0JaIpb5f8CpphvXSsgGf2G+rxqOQT/OrNdGT
A94E6zaMU4EqVCetjK+xCWtpYNJqaeR2Cr0C2pD1jP1VW1nsSDLXYOs4Lnq6
0/Ui/u5z1eG/iGmdIod32RM8kybxDeN4geC17clwb7HLZCZ03J6rV5HQSYYy
rC78UVllHhUPSNZ8ErXiEc+jzdv4PhRIJy5foyBniizy4+0OM/f2bd6i4H7o
2Tv85Ln7353s3ai1FK/2kospOwMvwvkSEzJv9mdw/cir8yQx27j/G3s+LWqa
NWnVzY6y9qNdVP4Dowu0tbYOSg08QrXsmeM7p4UZl1EOx2e/usrrDSqQzF+r
11WEkwPP0fBW+63dXQ0O0Y1/mwimxa69GpEdjvxbVfHDFPBaGpbNyBU8aXwS
oO3Hsok3imKdwZdSgs1sWzk02V9WpAPHarPnJWdme8JDAQeW1qRzNwcjcf24
VrfXUlwayOmzqnzjBPptnYqhCiKa7RdsMOQCENQELQcdOL88INed1/Sqf1rq
IGxUfl1Ve+sWz//Mv2EuMvtGQh5A15EyAt5eNE2CJ3rS5r4R64RFzVWb9htT
A7iqscem0XKSxsHPdaX2C1ftlZZv60bKDLPezJdQvDTCjqI1Bq8JYt7hZFqt
DrcMVtYs/ibT9ofhByG9ohNMrekttdZfbcD6zi25CQ89qBYORsy/ugXmH3c9
r6C12TUJG/D0zAyasW9QBdT0Kj9izsa+u8MqitW3Gj5cf2pAQCDbtvbdMQvL
gVHgLnFWU8TrvqLX+C+S5Jm/K9FetAYPBbss2Be8q0YCHwb/IOXWJgTwgy4t
8QDmk08gTeavhCiVmTVM0vlQtebH9Hy/dCH3hmp2EkX05DmDe7cd/bCXLtZz
VcUFEYEAWcwgbw2A7MDvS+NrmTuErKiR1lwmT4fy3YdCOQodRh0GFcdb3VZv
bH779xZu/mCgINpxH5B6yLXjvIS8gm2AS4PV2BEzcO5fc28k9h25/F+w3iYc
GBGHwKxc3A0GbcuvL9Hvr2V5olJ/K+4t9c/A1OZwZBOvH7agcwrJv917qryi
On2x6v4pajfPJm8sau/ygZFlJUQ6erdfjiyJnQ/HjRcUIAgQId/REaXJ4IPE
0IZZGImkfpUoaEvfeMpn/vAWutwXk1aA/tFCfkAqup+zXIIxLoZForD1HGSL
9pIDlnBWszA5CEinEN6/QRwqgIJoPYXIpr2mW8PXnfzDAQwwxnnjRsNtKKEu
/v8fn0NvRE+UdR8auiMUbwVRb4yBxBtRp3MKz/syuaQqJ5x0e9cyjIFBmxcN
UGGvPzUxdx0iT2P9dNkgw7ZEDG+Cj6qGjhIyMo9BO+iyoZPmc6Ufrs107zac
ejK9q/XpBcyGNe3a98fW//F9jA+NuwA5Fg92EdizMevAxX83CiW2Pji5yRzf
aR/XWClIf4VtYPxqkXyx3jBKK28mYCgGXG21U+iqgemnCW6UwiEMuyH3VLjF
UxwJQARSY2qomVSXrzydN6zAI397voOUrPTedf0ajicmxcB2a7cuadq39gwn
YrxNkNb9ET4srYqmniZ/oX/10Qr76MBel8ZFpb9qAhFRiRTyF0jOo5ksbnPb
FQeB6nPCpTlcUf8m5xWUO2NH4Cn2PBRg9UdS0pg1BSYYQF6XToFLdYmYF7LP
UrfrfWA9kxNWhuojmZ+PC46NPr7w8AShA6DeigxEOmhJO6bjvOwmNzukUZeK
x3QE36YV6pwsVNQ+1TRyjPVe74nySHl3Y1FBY89sS9fbBB0qVNMmUgE7eQRo
SYcPGJpL6RBAcUcNovZXD4HuraM12Q2olgrffY5r1kAkfeNSbmgWqpYFLyFv
vRr4oot5iPZ1a7hti7mENeChgjAKMzHyfvVtAKgdeKJtynjB+JBOaRmXqXBS
HRvgguEzc/h6HhuQsIMbaorsNVm9fVeSffuCf3lNCr0sJpkM/lgZ8u99IFCk
JYpip4NNPoKRO43D+rofHjD/5BYerUM77+fUFnoDEbHyYeB0ptayPwkz+PSX
AI28D2C/tcHPiPkj7SWf4S8ymCOVD5SvMxWD6XFwOh4XZlgp0wiHuSyi3Rkd
dveH8C5EbMlDAo99NRWAI7WkLK7u8ofntuo8c0PIcX3thlK2kBqZnN7/VbPs
hKGVE40YIfb6YOXCIAH0G4hlelNVhLHSgwmX/1y7lulcNBQgwov8wtdsW7wf
gqAi/8wZSlRi/Ru8ykglEWMaT03mE7STzdJzxBnwOkOxJ9kW4oR/mVBwh9Df
oRCKk8LXX9O5Fqlx5ifyXhULQYEW6efCZ1oF0f8sK6cEud3WtWvokRTwHlbq
lWyyO1TePAD3UHgCZK8tpLc+VDapGFfxZgdAD+o9ISyefxmw6oORwTLGzoiG
xGueGHQCYE0x895z6GbRvl7yaWwdgqrDOPV2/O8sF+kM7qm9sOwn5dvpZqHx
ZUmJZz++IPBRN18ycb588nOpZmu9I+hlDlgX/+96a8GLVyAeZ/Ariph2omPI
4aRtQOBO+iswuDNgl7RVNGxfEUg7/hCbgODszXZ8sq5DJrANEUFlOENa+eUs
Warv8xyw07O5nip02annhX4MnIWzLmleK+6UC0KOeIGfteIM3qArgbE5qaJ+
Dlmc9GBemNCqumE8Bip2IyBgP8+S3OLRXkNSViAdVEO3+wQ6BDgRXi/A+3C6
tu77abSHTP3o7+8Tj/ppPH9a4g0PIBrbXbrGzqYK9L4M5nK4TEDbOiRye2QW
8XcOiIecIyq7w4Vsp1QMEMJxOK26mK4+ETUEt6gh0nM5KchBbk50LGnEk9ZX
dWFkbYREoA+2gsdaGzknSRc17xuby3K10PPW9Hgu2GeqSa8YZi3YVaZyPu7E
fj0Yph3qpvibHhOuJyE9OXUK13dVNjXRa0bvRd0HIYLLRYkU0Wt5s1IrNOY+
nThgD8/jLan++viL3PmrOvsHOcMESsOk38m0CHZkH/vPeDQy4Y9GZE7s6FSK
pcwQuKxz1Basi1u6BB4fbT9u65HS1R441AarroDb62xxcpkZiNlXd0dYNtJt
fXXXJ6NSODZvF3TddebtRzxbsJCJGrPZLdvd4kWTKRz7DgbIhMVpDJJDaf0N
dNRpeR0olw8zQL6eWCEv8vUaN469DN5KnSw2raR2ddx69tSjVaPnGEOHzDfP
rLXuRwEc87ZJVjxOZeDqWvwabr3wvJdGiw03UyfSPw7C8DKkZc5rAY4wnQDh
+l8LwVcGBfMfDB+0FeKOoyXR8uIJgGuiFj0CbJBwLtwn7SCfgVZSiyiYPXbi
ZO52JjJi7ltBQsr81ASmlUYBf5IclwAFX7N6DasGJBY+FVvQc7FrboVyZdzC
T9ro/7O6SvJ8i4zdCSJpnuB0CU2wN0jyCsX+qxGFzxpQnghxQFv8W6quFgSF
9Iy1eaODiC544U+rNIdo6Wt+/tPwYwjo7PedeuBXUcLd1XOlqqMhVMIB/dv7
vqICkNk5izezveaWXdkqRffkRUzYIxeJ7rdL7x/J6oOEZ0n4MfDm+jAFYiPs
b3NkmsPtS3szpApdEdOk/fxenTnJdWsSF63KVVzFbRPqNFYQ/PNY2VzRujcz
fMpxuSzt9ESWYfjyaSZg3Bydy7wcMa3m+eRSugqL23EJ5v+X0MNEb57OJxo4
lxOnr8ZNqYyK9KO8zbBZ3UVzH3NQvTvm8r7mBrEdwu/e5lUziRNAe9KZ4+in
FM+470JXLJZpv/1w19RgA99dbIY0/27qmIfDPWZaYoTON3NlfGyqCGm6NoTH
rNyRxrxslKVTySZb+/r/COijijtDjugvlI0K+zVD3YShoONeyDsOMYQLaR6P
ZwvmnQQOUf6e1eOwWvCGJYvIU180jTTUTZ1pot/yAHBQeMQVxaZJ627VufC7
eTJ0mLX8En+eWJ/b+s58OSpUPHY9uLhE+aYY/lU5JnRhzchb2BTrzj/0g7Lg
rd/vGaF+iVlytWSoTGtG8xMSfzNSWfDfBPHtm2KHfB8L6uHV6cHGSfMWPVrX
a5gSH1SU2klKnGC7lF7uP1/kHjwqI/ou6g2oiuezNnQxB4R2cG84HGBIfsj9
xcBSkE9MTl5CBohO8aW8XKSKwfnDn2LPtGiyZlWzARnDRpGPXzKPFr4RhoGg
4zVFX6t5omj1JuLw8WFl2YkcesdvVdDBvpm0aIgjJoEmYMQn8P4gACq9CtYV
Bnj2tLcge7QiPXKNmCJKNf7oIoa8d7capMlYda1+OKDCilDlFUs5Wk31eGX7
TtV7T5RV60dddx5HL+i77FQUmM02IMby5kkquznG1OXL4704tysKJYgwCCif
laqvH4jtHVih8tbl6vPEwL/7bzNvihscATUiwtw9x9beCVrQ4wXUsnB2/Afe
6ZQ4RWy/6T8QcYUgzI7d4XN1MZoj9dQzhSnIXd7ufTdGk/hNtwzK7C5qndBJ
D/JTRzf9iMvl4HNRwrVcR8/vhEJD3yYbBIoE84xLDdlMZBCnGxH2/csueLSa
NUcVHas0Itg/INiw0p/yFve6Y3QY7sB8oC1rmdBXxjOR5yfzf6FxgXGt3zcr
Yb4ryWKimfCTwawTGvLHqLrd1wcRJp4V+ccmjc4e1BSDPUq4ZyQZmbSHUwEH
dt9MWy0V+EliPAhUs4W/ag9IlAHBLAus2WCo9hI7ERHKOx2tp6EtfwUVxY68
kL6fAoOEsBgjHZLLIJBUnNKZ7IOekTNyy6/uH2HPBdxnoiLDqU1flCILla/J
zsYYF/g1OuD5i468OmLlFPia6zmexb27bDpa+69ZBiCup3B+pj3Zg/ti1G6n
RYMvWp5s4ywEPOzwuZCcXLiGAiSD4jcTJwTVtZJdH/1NJPHRmnxSNELT/Jvn
VrpgEov4pr0YNpX8uAS3XexqW1N6Evg7WIZ+IJq0SgUQfn/kWUayNS9Bqy7d
JqmQSN0gJnpEks/DGTtjy6lj0xyb1LO2KXKL2d0exlgfqFHZPYtXlfCE+fL2
yZ2UecyfGU899VKn1/OZepxEM/3XpjXRqyX/ytj7cM/Pgfes1AROWwUbjYlM
xjR3+2WWWsU4Q09AQMW82dt+SmaTCAAuyaWv6P11jc7TKRz6Mkjksbs/6MSD
9UvaWUtP7Bkg06zQziJGcwHyYd4x62PI1rtWSZDPDHCtx5+EZ0rZr4wtJSXU
K36QSHr/7ObWXBHwiJpWC8N6GJlwvnEnzpIx7wjdgmC5FHKd6bZMneRoEd1X
yblN4xgbIXUkRCUGX4qWndJ9iWrd8v3jwo9vuXP569GywJBsVtwb8+2cv7sB
efMK7rjBZJsii4jVasW4yiVkhshJkcLqLMBoyISWMbZjJMGh9jWJfF4MTPJ1
63arHT/ncfNEFpDJojuWdIkdAZssqNaZKol5qHkCXn0r5L3rEppLyKo2rRAS
jgpeSDgGluCL4+YQ8FoHPqeNU3bPUbqL02dae8SDwMrMj4tS26A2hkVhcv3h
XUygrhpNP1pAmdu+/6kfRHEeF5MmTLjtY8HQoJJ8nuWiu84NboblxvdTQXT5
/sCevRNfFO+XFi1wsU2iMScRpRf1qm3hN8+Y5qzc5vSP9kloeZDYUcBna7n+
1KQPs93HDs6K0y3dVdFIHs0SjDJCFS7G1OdngllEawV8yymZC7QK/dCWqpXT
9vuReCtGYgjI+PQvGMRqjh4K+4QiZ9AIVkADvPLcvzJ8pQAVMsXgJ5g+AHhq
Bacl78bIhQYmEdDsMWSdx3cxfl9eAIW6XkwsvlWmSyK8IoaufaNjEfVcOLgV
itC3NHbHRTbQioOPS42xe8srNuhBNu0bhYlVp1a/w1MIMI/wqsthmPLX2Tqz
YqQcRM2Zn/t+mBI7A8xIy9x/jhdigHRjW5R2b3y9lwBvxmUV/KCbA263vBdf
p5iPzUisbYgUTy47qXZgOLFOxgNps1VcRZABh7zY6lyYHs1kOzW5Wf5zv5Jr
ksdF/2Zmrs7L4EQfiSLmIJRrv1uHJckzFmxZghlk9dL9LUfFlrmclfUZr1gj
G87JrOGu8Fw4O3ZrXh7Hz10tsgm+NJJf9Bo6Fa4mmj2yShqTdlHdJk+YmkHF
fZX4m1TwVXP0yzxKCeB9tkgWftEeMZYLCb2N+nEVPhVRLDkxsOm6r2k/5IKF
qdHjz27EJbJ29pnp3OSTY3exCGMr81G9ZROwYhK6O4xzWm5cc/0mDeKjecNb
3RYzJLEn0B/0QIllTFPRga6S1dJfdkFjP0ENi54pYm6XpPiwPkF9uS13CMbz
SiZziA7Y+VVuabugGZSZShO3QrITu7r9T/MFBB/w/Bb5bYxVFV0jmurWmDYc
rYLh5H4kkgR421jTWV4dJJzQz+ww5pbiZ20L9rk1ySh3+KS1gV6YVL53rbcA
UmVyzz2tF+e7v/ODEvwA1PfxExc9w8teOHVoOVfhdUQeM/SV2Vll7C6MydOh
KIlSZzetgMOw6K4AKY0BUFDC865afBh+eAookhkSC4l7RZEz1uZADMH/LnjV
LPKv0cnvRKQsb29+QNq8P1IqNdCs1Nw09B5+emjev5Zhk1mmjRR9tK+R+Hzi
ORMHaP7ekTCttjYm71qS6PhfcKjQH+Ut7sMEr2+EPPlJq2Z8UslTz6ImSyLB
URwSp6vLPhcvJy2YGU2XjhX/MT1rtuFqvdd29nGKbLNrxtCxj/gOTnp3RbYC
hOq8pAxQaUA9czU/6WLlcXhxd9Hw7EssVpLq3+429kz/rxNQyhO3/nqsOwJ7
HgHSVt9EsypgE4AUeYASUZyjmo4x5ZXPgBI9V3bQbZZLREGxR8tCwXUO+Eug
IhaXecJ98GNcz/XNX8zYrfINA3C7xHlmQDPhBe0TVC3GQkFMrva4SSnT/Buj
ApVn8G+fqfyj0k1thpu4mC280zfgFpDzVVX49Wiss8pvJh9rfV4PHP8jv+bS
JvHC5lvceJMqHyCm0k0lVtt8MT/khd1d8wfvb2w3WQQxILsiuyualDDc8AMW
iDcuy3i7D9RT3L26C5/DVISYSAA7U3zkFqvr/Yxf59jcTeTF50K0Fa1NXW0H
4BXH5eF2MHc/8GDTBTO1IOPnNZ9zzPJXmfQhbVZTAVUhhzSy+rwMo67KtNy2
tIknzpeRo/6SG0KKy/sQwkT9UdccubZwNzyFij6/vbCPTrng8a0+F33sZfjc
Kne1v8Q+CqKzFpbBNukrYd2/0PNiHHQUfBPPexbhk+QQl49iHJaTNlW1+qW3
qct6Gm6tC3sxXKDSS6OWFeV/YZ2F8VdmYX/5b5wdAfNTr+rEVmMrnS4u4vf0
4JUFwaYajQxM5yapJJUcxVnj8eoMh3wvDud41qxvz1rnF4XafSGJSbw5I2Xs
GEUK/KNquheYlH09JpL2Ve8OzTHlxtoqnRqFNPn2AfhYhV0S5qtDiC1jWsub
bCfDq7VzQqPJ9REiZp6X+XqQ7LuDfDnW6Ev/fa5Achiy+yZDKkfAARHVBTip
vO/3hC3LtiWDn2KSzbaZXlEoDI4Y9j+93D54PsWhhrFRbl1SK4/RBVlmtRQa
eabfLV9KD3kMDzcQDGB0BFUU+ODAKXCklQIGj0WlHazywof2lBqbCq3Me+O3
T4vswH14uYC3O8n9oXDU/+3jy1Iu5DSuajFu/kOUwncp5WBMwOzKngfhgIsp
yjnHWGDyKSoadDWU85T+VhiwOcvUyFvr57TWA3ClKc7W8VbgEsNs7GyNIHOj
0SvDGUl7ACuFVX2G74WT73G/RW6VCtF9XAhe8CoyOdoqt3DvHMwZPxobdJO2
7iLTzliOGSWVoxK380MTkV1C4aSUvFTjt99S82//Zf4bs4PvR97AHeN2Q2qf
PrZZCfkCXPuLFAa3+wVN/1SqB8pg8gkOMZhnRHvBkuGz021aVyIprfnd75nJ
jf175L9EgEFeQbn9Q1Q/eZnLmulWR8BaZ1e1sQyGna7BrmZfac34famNirm/
n8eY/INpseIByh4Qf0R4no/5hXIhqV/LgnmAeZY0R2CvcJvuqHyGm+z1WpaC
m27cQE1QkM+MprrEu+xDhE+YpBRTWrzBY4xM/FbkeM27oUbe3BqtECsGlmse
WdQanXQY5LODxTv6WPRnG8089/9vwPS9yOjV3LSMZB/AHFEJvtEsBhj/fp0M
gYJEBldDYO8jKFny9WfhWg/MRn90hvnCjgfQugj1cJDpEJKVDAq+oytf031i
z8NEgu8nt8ejnUeA9nchWTiwzDI+TARj5W5FdMtbMTWxU951k7t+/lboivCn
DlhwGTVq6vGKW51qL2A/Cn3tJt3rlYZkbw610aH6ZNNh9qICwnO58GVEn25M
skPkBB3wjuai+OZ2H4eGy+8CsE4l4LLCMnR/TUkGD8cBa9qsOwMuDF9ZZ9CQ
uX5BvW0YE9o1CxLWDpKX1zdVFtUcD35cmVHuZw73r/tL1eMSSRa9QPScfdaw
QtIe5yzDc0f/SejWOlmoCKFv4+O+u7m8Fbs94poY4wozTxEexzo7QKKtkx9a
Fn9Aqtm79Xuv4Amzle8bkDI8jjUgT4UiGp/5VbnYjEsBl8epoO1YTsvLCi8g
R0QT0dIvMzSuhI8cMQZiLMEb7r1UWSkNnqPjw0mlFnlWC/do0uCwfKax53Vp
3rd3EMF7ipF5/YF+Iiq8Lef1jVYHs5/SPi/Khlu4UVG6XtkvhE/R0iGe7UxA
X0EVb5ZtYI8NzZOw7zjMSNhIziouyF0RtBtsQpvb59gsjaYvmymj4KayxA41
ip6JBO1KHSh33VovI6mkzeUzAbc5iahWUTb+0DkCb+HJgONpHBR2oBAIQuRZ
dzrkuo6CNccYSbkrWfeEEd8AMQZ9DQIciygsj4tjncaqoKwq+rvNw4L2KIgd
od7mefbJagy1C4W2k47YUJzjRPgY+uaJAHiUNOH7PpJO3rb5sIywy0zDqjc1
AOIvwIhW3XdrMiKQG0v9pLAN1PDHZlX5xANsPY6CZXLMHxQqUfhEW+8rH0p2
jzaTh3bJWQzVuyaO8e6e0gilIWHxugQYRhwuMq8yRMeB+QAflHHL1OMconRH
ZWe2xHXyJGnjVSnl9pAInoOUOEnEtYFQX99OGroO7kSAHYMLm2o/cGUONu1q
QBZJJEfaWwQFlHxrWrHBLFSKN8cvxBTt+hz96XqD07iXJ9FOPmV6YfKmpvcB
TgAwH1lA65+oKl2lvc1gjgBrEwwClwmANVko6SoBszKKayp2PbFQsXmsJP5W
MhWLiB/XT0NfOuaM+UmJIXh4VFguXIKPWipaAs85RBTiX7ygJs5XGGFGm6zv
vmfWT6ppdcGt9SROnQjXRS61GPxESjUQ6TT/Su/6b45PMMkqdHMWKgTJXbaA
RV/p6PuGzSnB332x1hL7U9U4iUYklFDLH1ytJAY2db8uDd819SjFcASnD8Jr
1TXT0u4FDbX4DbZNW4AVOkzxKUnOqGzEqMprHysr2XE4QC1eAeJAmXPukj0z
o1BD5GBpxX5d5IlRDkK6C//eCnYevx1MJBJeZAvvbM76frZZF/pRhnr0ZGVz
IP9eACf3hpbGrx6YsLbP4YuF9X2CYXi3wPgbVXQmDp3Mp1/rHZf7aGGylPJ0
96m6SkzdFgP0py9Mqidvv/8ro0la1/CYi5hHPgyunXEziwg5UK3QNQ8BTo2p
z+ARUKxe80BC10vKOY5ceuPW2CL4DrZ2l/k0onp4lMi5AWXs/wG+/Yl9xtYI
Rpm/H03Z3Y3IHSl5P5O6Io7G3Cvtp4Acul4Ze0IzseCHS+TYs1lotN8k3YKX
A7imLa4JqiNrPVp+qp4+T2+bOS89NYrRSqvRWo1KBtVkptlGOx68MAfq1B7Z
/195mzarHZj0JJNPLnKrcV6/qPgB6F8LPfxBD/Z0jpqPamTh6MiSVNGuhQOY
dL/C/Olwnmm7MB+HZnypZipG8ymapROMv+RCJTUBlh1M5EAGFD/MucTH0YWl
nlWyo90Kp2Y5U9YvH+QKr1eOGJwBP3dgUDMkAwMLlYpcdmF3FZx5iIACwVW8
gBVO4zszMsLOsO86kfVARq0QayaB9Poi5D4Ukp6i6zc16OMyhKmTR73a1Ovo
7fEPL2zl4+EoVVpR2b5iSwrqdE0YBqHq9avA0b2sZVfu6Jb9sEK4YSY67G+7
evlxbRIjT6p6bMZCFW63f0aMaNojiHuFqoeFix0CDy8XJa4we+JVkiR4yTJ6
/77gcyWjyf5fM1hONePAvAiC3DRP8V7yRmfB3S2z4nyiZc6wwlX3lvPIM34F
3o63Y5iqbq3ebZMb/EeXRUkTN5DCR1EW5IKk5ma1HG/JGlo0GSp6DvmQPhCN
XLmCgTE5njwjzNc6EO5Fr+bz8EjetSZenfwLvQSfJOqjMbQEyDNn5bjWFfOu
4066TshwrFttlBEuXyvTp1omvO7DAtX3AWUPmq0n2Abf30QJiv/sx+4iV8oR
wX7lnm5k53cLU1XSqaPBAJgG/z9AuHX8QHZwWTyyRXkKrAkVpeaf1JKGO3fh
ExBHVnWxiI7eeuZx6kb5HYNAxhyTsdz3zdIREDCWhxfk7Zi1mqG3q9sNDi8g
10iqe9voJY6LifiNN75ogX3IK4DucQoUL+kjH2ZEXKdJ6IQRSXd0hytkxTdx
lyaa0SNJVKwuDLOSGLfpZBG/eguMq9OJ/Q3sl2HoocuxSjGPVy0qz4osuFCG
60PwjkmJe75ri6SMDwahZWAXs5s/IjP9/nxrQfYwjajJCs5wr0YcerP1I7mL
4de65mWyerB6BNSeYE5ihuY1MqPoaskDfJ0ytFVgyFKtwiG4u4uyb5LsbtmR
W/UZ77bCfL4ZF2llA+bzaiydV9/kHjbV1hGKp/tNb0MbOCfBO5NbL75Dnc56
nQHRA0IIhuNYvHAbm8AsbdMpJnTXB+dKH/Ux30vcbMbPiGY6lWrV5h2vea+B
T6t20cJA8jZlGnbjB1HAFeDzTDU97K+BQgX+pUPs8n9JDJAwvXkw21Mq9YPp
eNUlT2pFWv8ySaEKg7ueLbGs3Op18hsbbMXqb4WQBJa/iQQGtj5sNSEWvb0i
4GTsOixil9OU+eBRA7/iFJpWyvvW9IzvdJd71D4Af7uqpk++HGSmPP28Fa4f
lJZCYGFERGa/fWFZA7qpZjvJAdTFzAK25N6LkOVvo8CwbHmYkrXqlwQ3iGFZ
Vc0BkbJhpD5O2ddhZSnzl00RRk4xZWIenU9BWYOfOM75zOo7Ji1275mFrhgh
SJmwBryochYi735pMsAKfA7bRwitpn4qagn3ondXUjYqplkNJ83blViWQbsQ
poFWLJhc6fhRSgBfBooMFk+Erc0RWNcodHqk6GGnoiNYfIMsXpIjlChxBXBY
1WF1Ukquu3jfCsO1c2uEbfdSQLDCNHKnRZVR/mnV08CT9lGd3C4jDS+Qnhx/
Toxztc1UROUCoiacKXIE8Rs199mDzb+/DKa4wslDr0W5GIk1S620lSq8/uW1
MhldBwYKDCBUrcp0RAda/lDcT3Ua3azp9UafQqPCMLL5IRk/yX67VppCLhax
miAzj0Jz3FIJSCreyYDahfW2CqDzBqu3aDJ9cvvXQ1jy0beORciYWrCLnhC6
dMkzlpDWqU+rXlgK2l8CU9oruGGIot3pmE1c5NKHTJldnLWP1oPNsMGLQs8I
KzkdIBv2VGSdZe/d+OmJ3uBoejITZDwTK5zMvfdCeJQNx9ZsCgoFIdQSV06t
xX6tAOLv/9s4OLlz4nWbDfTQGAhl7AKihUlLAtIrJ94gqUi1PBjyCNYvO063
UsYBABUpm9wl3oQBgOFuiGPy0GstVVZl5qgiko2XPaSK2xdeNLgKWjZYagel
2EmKEA10uorfcM/B1J7OPxPLdHBojoXF2e5o+bKlIZ85z06G/cUeF03FW3p2
vLN48UzR9xj8lZtAI9Y0zUQ8JiWveUt/5nqQ6m+5tXi/INKTFWzfZWnEBLv1
SxdrBvbVBPDO06ueCVvOyEj0nDOA7EUE0GjfB4Vt8Hzi7bfOHaiywvYEJ4qa
XHAyec3htz0H4FfRqXqctz8a7/hvXnRKeulQx0t5qVLWp8q/90pfBqkTssJJ
7MWBv0Nx1InkZKKKzsq0bfvNGfo8CHxBI4G9XuRswRSYjQ/KFku8P42vlpW/
uZcKFOwaixw5FF+CuVluLILrAa3uOLgx2KiXMNsiI3hn/8JlhfEiKAVS6EDW
2M64HoyRQvhU33KoxkdtCc2z6bVVNbdMNnwcQCSQT0J1Cee3d2hjj//Jy10L
rFpj7ulbDIGAxPMKKBpq93nnTwNgG+0sKk/RW93HAZlsSWb2UhlI3XAiPxBP
QRpK/z1DbE4YDR5JD/Jhhuqc/LkTzWK0Rcrc1GOLZd4I25o4xr7q/kA65J21
E1LToKhxEReDfq30feaUSjoKmSj5/0q38HkSxfVNRefkbWQ7CiddzejiowEa
S0+dJ0qKxe5dxiYfpIKhKjb+zSP9tkgrRY/+6dKlTUYhheTPQbxAmI75ve0N
G34/ZPwF1reQOdVmeJio8tXHWq+YSS0nf236lKN2nOUh0O98I0XqrEV19HrL
bSR2SdUGTd8FouQ4hj2dL8w6UFlKs60fCucS00Br7CqrWGasUdaSMrYDrPbs
vGo6YoStwByQ2BdVENHG889m1oIAPxchOYqMYfpDFobBRVLEYmIjfEPpnimQ
28zC72Nbd9KfSPeN347hohKfPAuC81Q84Idg8JlyURP/eBgWCrWyzgr3+TwR
m2WX8WhAvSR9DLtxZZ+C7jRo1Z+OcwqZqL3RC/aOO5sIJxaB4/I2uv8rw6HS
vIbZKtYOjQoQ9Uv/C3XBb1WYq6dEwyEskgHWC0hZvmZYfeaQcXpDKdIbnmMi
6a0oqaEFtrEOlrk0XKASmDhjZ39MVVwTNVpDS32FqMZMMWIFTX1wjd6wRF7A
hwxEWriLjpPBzytNIFa2Jk5m2S5ifJeCIu1ukWDtBZBoKn3LG8Y6Cbbr5z91
TESZdbYVgOSRXOmGLP97WN5MFXlz2zGBEEtL1hwKtzIEaFMyvmNmT4SgvHlm
OEKxpDO73jy5XQsj3oTUJGT/UmWmZVpo/pPyjI06EJFo3p/5HKB/pWuV35Va
+EyWfo5wHq8GJcL2If1gBVR+YLVTn3169ykPWZiXNri5ZbqyrBAMuQNejyvZ
mCe4ZiYbI/3AwaqPrHcjzNnuCoMl73g+wteXVjZ2IIwrfWVzxabzmodwJQk+
Ns075zED93ETff6XMvHv29jFhTFJYt1hxLa751aaphfeaIO1MZhehj+XuZYn
CFfOwRmCeJ+ZZRnOa4FjP8wjRBTy455d4d7/FjTs5w4gD6XRVxu48fKm+j41
kcBhp3OaTH7w8tj0vnSyFeTKBdtJT1xaoLCtzoAwjO50hdI2lXhSGzqMAats
tdKLDTbYolDpWlXkatsj6YgHUEvuwbFRrBTa9F6Hn/jmL+Bk49Cx/RhI2b7R
776H/mAVmfBMzGUM+Dfr5KVTIbyn1VJ79VpaO8fq+nRj0O1ZLYCXtoe+2BLx
r5sjwYYDWBeBfB41UHU72QpjW48LXbk5DDqrQBM5PEurSB/1dPF5MIf1INOo
+MxTgvNKvt4PaZoYAT1AHnkMwJS27R6fTscnO/0VKPZSTSFxNcBriGwkBqeT
o1OyrhHz5pxBZ2rqhR7Qv0OzjJW1780elhmd3lzHxiodyAXFq/zXF0gbjNOm
qN6F/UmQ7BbAPERlFQwrGWkh67+RfYc3Us+oJA46IeV/bcWW8+u0vCWAz0mq
OKf7m/2Ihs0xppOz/v5Q8DkLuwOoLr+g7rvrK8qRG0J5cCFNrZCDYScBJXHJ
RuNk+TwdckZ5O8XsZTZyNIGTHUhk5jIoPCF1kzMNtuUN/fNQju8P2yIYqJ+O
ckZYtTgHFGOrKiFS/xg5tEx+iQ670D9zsbvVJ2lAuH4m+ZL40xoETboYSWr+
dK1jkBxT8DlNTMw79JeMiNy4dWPGz3a4FQcQww7gll75E2S1dOW/P+eqP+zI
dFl/EKCtYw/EX1HYX+uWEbkjukUMC1ge7IGg9frQYWXd8bJaqjJkJHCYu7uP
lSOpZ/hbPjVlm+cV2OdtSwaG6AIxyMLexU3IN+TKnFXX5jHTE1mQerFo+XAU
sm8IMQjONms3kfVahnUSQTUIRqJ7nnSUtxJafX19hzTJrSonU6cic6GYfd+S
8/8IxxSeMAfr8m6lcj0YMNNGUN1evyKwUcLNcNH9N4limNkImpwkhVINfJvg
/wrEKS1EUOl1TCFPvyWiWHyDhdRsihr6LmyizEgUc1kTwQWW8JHQAcemUusN
ZCyDRteZREpHC2Uz4FXQEIYB9PkuXqLqWST9wxOtwxUYOqxWprdWD9OrmvtH
OhWQuJAx7Q8kZScuaMt0lSBgWqIJjwibWN13vi+LOfXoAkkjU0Jor9IPi26b
HB/MxLVK/Iz/zD0m4asEjV1ryaDEotfP6X3uTF8v5eRR0kE0G4VhZQ7pbn+y
uu0z3nQ5ULige1WwCuNuBGM15onWqvt3z1OrRFAxGh3gmF9ZsH8PDMC5KP1v
2xC2ZLBgK2cjSqJZfI8tjB5qt69n8ipdZqNNT7J5JvlA6KgmcnkyEJBvmYML
GylNinnIDSk+5ujK6eSDxeRb6sFA8VuRqCYkc4z99P7f6S1z07hX4nl3JSIP
aF8mndvVCHr1+9lAH0MACwLh4K2bMAFuxzlrMqzf5EV5TL8d+wpP/EpZT1dy
AKB6fZoN5jchYpXQqr0+Ro/ecVfdqHS7RkfmN/4a1/58SWlpBMDymHph1O3h
o2peagLJhFTQWrvKyWw5lZdrzCwhnh1LirVi3MiWl3+xHaxTcNGBuI/mJlC/
MoZmjaT3Js1bNlbtBblc8cRU/YG46DcMdgRRitPWuENmJgR3HejLLEPb9iHV
hSkdsBJ29j7cPpWuza7l2v5SfJgU6Fh5jOqlikIlYqIbKr/Dji+U2AxDRbZk
jBsjutWS2RHGZaGpsvP3P+nA7v65gygXMiV9Xkhvj6bOSbD4l/241qeKmY0q
z6azUmmrMVkIjwTb9YEcKeQPF49/ALf3c1hmwlHoIKDlHJAy28YNSGkO4192
F5hSRS96V0B0526BxYt5lECy9r4uPjwNUN7W1YHWAv7lh3tTCPXVbXTCADy6
iwavFbI7eXwc8hFXz9zjXu+Cm+rkFYHChxK11Yg8UaJYoX6fA4TbnSc3Z1mE
F/P03bvEsp5x08PRZ4Ljc8d7ML3zHStVz2ZWLYQXAure199elim1Z6NvnpjQ
/q/HN8Vd9sYetNIAIUxIkPkjLgTh/Ne3M7E598CgV1hJ9ti66Vux27mopglN
HigDwVzQM6mR5sQ6syQ7UdMu4TyP2i2FZ/m5piXQCgJ6Px7V+Ma76iucj3cd
Ory26VmGWdUfhmdhQocrHDJew5jp9mgGga48qGxD2B8RerkX+suyzP2OoyYy
Gjti3r1gp9FVqIkO/KfzgWnmMXXiVRA5+pljmPvS4HEstZRrX1en/zUtn59D
Bic0fRaVr3tRecWuSbUbYYMmc/VhxVmhtPSmWN8YYOndTDn5zPUgyaCUF/of
l345SGuMRaCTC0sUH3MysE7pG3fsGPcRTg+AR/gXoHMtuk45sSdZQMVhLV+L
8gNx+ZnMmhs4jUctnlWXV0BoMzOw02XIyF9SVsWmz4NZBJVB1XEnBdOEPzSp
9TMeq5mZ4a2QVrQtFAZcc9tukrO3T9XTtV5e3r/0o3rwJMyDgpQadm4lo7e8
3ehqyF4xVWJ3ZbNOOE4BQkogSeg6w7xkpaWB1vwAQ62T6wBMnjRrEf/smR7s
ehIU9QZrYfybiVkHNFVaYIQTOj7R2PzIMQphWw7M1WTUUuS8rANoV39xtKVk
5X71hhuz/pxCA5S/pee5Wuv2LfembWo8tGYNWZwnuuQB9dWvaB1lo7IhIIDO
NVQ5yM5XxKzchrN4WS3dRFIt6OKh/YLoSKgHDcsbpUmH5l0erV1qvxKk3ciQ
LQfi98nXEWOeLrKPSjNTOCvaXCsJloNX2YC6dFED8oo4F8Gm0XFDKxJZ27wz
Q90kbEUg+4+XlXckmhBmgCZxiQy2DMDS64O0/GiaD9vgAeeiIDyhv1A0cTFs
5CyjfstgXen59iU+1QZm3xNA4wuf6GbSsqN1hdlcU9V/dwhGKdlAty0UNApH
hqezpz4fI7J+kvfyxNa7rd0za65HKOKJWEq1WWVY7th2qLPVO1xTgBF0AiFj
NeK8LJDGDqrqDj2aJsJX3giK0Mqs71qy8jQrib0ocXog4WpQsjd8/lrH5Pzw
3KCzt/3ZswUeWni/k+awwytOtLdQcDAe03sd+8K2vyUYYVaQtMOMqiJSIdf0
oJ0wmK9BGHhROe3Y4DqbdSrtfGXzXQxwni01YpsybGRFwzJgVQgxJtgQknER
wSKoLoqX4vvot+VSkf3k9tB+aC9Ol0sekqhFOTC2OCKy8FokCINZMjrDX9YB
esizBYkfEAzQl6Uc06hTg2TK/9mWGJmC+ByBD5sVNiL4k6kyxbeDDfKbZmGu
fB2+5w1CJzhGm65tU3kokzoRS82V+HmNHcPeiU6r3yfDse9oavJa6SVrH2F3
UE4FvbieCigQa/e1AXOZ2qoEAKI+ldUni/h4eXgQFzSLfVJAA8JiiR5WkaXh
FY+FrtsM4m9wA+D/7z4SPFnAy5fjoedRsYkb1RKyL2eH1L4C6P71YD7ZZkj5
2N4/k8+1PwLkGGregpqxNhbGrhlrMMT6JbQSFV00NuZ3jvB4QpxTaN/SCFmk
/s5Qfhgf+7f8BybabDeUWQQRF05nWAPgERb6KtJ2YMc72V0jC7/PaOVwocTF
O8EnealR+LZtAYrYynlqpoNtOZSiYOWCyYw/vUDA46oBvP3ssCEv0BgYZus6
IEgEssH9T3r06IcLmaSK7Jv+REBVDpeqegAvOdU6BOdnOCRo5x4WYNBEsn1X
yq0ebp88UFlCpeeqIumMd7EEZgEi39bme8jnMO65La7EI6VQEoF3wD0ymGU5
OLdSdwoYgtChVN6Y3RKiivz9JyZeIOnMcy4BJ5gDnCccJmSo4GHW9TlYLJyi
gHYtJ5RafAGKA9C8egj/6HlAH2pWOue8bkaj7ycLSuN7/F8HdIh5KCxfytXt
w7szTYy02hGFqnUwMdkBnWBOz+CM83tOzrWdh3aOERFAbfza0ep5mShdal74
c+WW5soCQYiDUWrCOGe4V+SphFwJx6KavSycl5yEpNc6Ys9KCKFB+HdaV5bq
kRjpQbnbdQCeTdiWXtHpw77ufg5aQ8fAe/crMVkfjZvKZk7LXlyTJ5Ojszf/
dBD4wvuOqMZOl1u2AY5oRxrPI/ZF1QEhyQMsqcX2Jv0ornSzUzJhCns63lsC
QIrDBnEjJ8p2aqzCaShZf1jZeBYRam2NEAXpHdytsitAsx35ci2giITXUPkS
nw9osowWWcxcExMtPNp7LoT74/n7/bSc3u70H2UlKqVcgHtL+xkQdxJAZAEL
+9uH8WwPSeoxfIkV0/SRg6qISe+4t3UtYrQUvYqicLxJdI2KAOtwvX3xLNvE
HyfqbkgXQJGNrYqs9jfzmRHYn1kh3bjDinkEq/qv9NpYgPzhHTm7Fc9x/EW+
u1OxM5AE0QXcHdG4scY2kXsxTAZGy273rJCR1HFwdBjSUahRRN0G45OHQ0uz
EvsIo+DT9t0WE4vWPpMawc8/PYU/uU/ohEm8BD77w0vuUOxXatuMNe6p6fqc
eC8nz9Ja6G+NHhJihxfPMJ8FxYXPLTlssTE7dwgaW1Q/JLdnDJiafPRngN8u
Qh+x3PV4pRBChWNV7FimCC4pnxneeVnULd0/KQ+rfAKpQs1VumXxKyikbHju
sCZYYyfKc2TJl32kVAKRsI0+pFyfjIo/PEMpVvCS5sjZWgCOkqaT7fmxMqb2
HLCbmwxmoAfnkaAyA2fuJQnnAqWKBwR0zMZOOR/i/NF3Ek19cCDXblhug8Gm
bIvZK/3YPzAXoeo4BKp+QWuk5jwBIoD4AeF+hXlHornnLI7Em/yi147g0ose
0vMuvUtoTK4p3R9ChIWYldf3PMIk+8DZTjCVo0kMLObP355ITaIjc0HxzOY4
W+Oi7a2L9Y2NPe8hum8DE+v7Vex2yBX4fBu9pItqgQOs5eFFUQ4ZGg6ffgHP
qyNwkCVQVdQB+UtebcdGaWlk6MIQ5J89KW/PBXzHIUUBZItdcZOun5YnG6fN
CRBztwH0XQFgLf8niUWuSAP0Y4GHBC27Ydnri0rIJPGBPWDpDySuKX11YZra
s8M//GXLyAbLryzkn9MqtUZwPnwuSHHuhFXplvYy7WHe7Gjm2tWTeyaWFH6c
D22uiuExXjg/X6TB533ga9IgYtK5bk+C+Kas+rIwXhIBV8ynaOvX5uzFFTtQ
o3TTbNbcGudqGPpZItWp7UhTXakz5Z0msWHMGc8LNVOHR8F049ECpnXIyPr8
ThIPHGTMk1ehMCR0wSRxzfOetlHUqAhOzGE9r2s9DJct2qDtpLoPBoOZaE0S
0F8WlEJHrl45aIGZ4BUVVlSBO+m47zwIZ1LDKRQmwddOrTAipMNamzMhHBzm
4q8xJRGbin8VVONOv6mdgQ1BQZmHhDyla7OX3UMyDioJxvJNvZy5agOsteZI
RIDeU/aJvDW6j0Aepd2RhCM/jwM/K+MMHkwpo8CexbIJi28Z+7csiWeAuIOF
Y/57swp9jz1j93GJJj0QUKUJoMiNWMW0YzG5f5zgp1UtDjunurd89Q0V/0Ws
EYXm1IWkLaQLJ2pjBnckhjjuWAMWaK9nsKbvnMewsIe5BNe/Sow0yYw6Ys1B
GFST1NZiI9yUBPgRG5MW2/u3J8hLbXYoceifko2eABPH2G/Es4Ja5EX+MVnY
CDE4BcQyxpKKx3+10CqCo98YZjXQ72OqBqvQ/GwRmG8wyJVNijYFPB4kzzT7
++srdfbdrPP3Q/L9AVjYFeWB5qFg+/3mYfqpvpHgSvUrDBYDRZGLmm1qgcjJ
n5eSVOqS1xUfTdgo6aGHfCdD+Urezzb3AggZ3KjbvQPokfyIXRnvYGCbNV4I
HJgWBRMxOv4PUxfkT7NO1qSvz5sFGvrHIVnIsqmCqyn0JT9e/gzTw+1Uz7ly
6Y1LCbijezYDpz3Z8xl1JnDDhmr86tihYk/ucZ+7KxyD3K2W0SXn6Jt6HuMw
z2DK+6CIt05Tzq0+4IFbN2kAibzp4Nlh/PaZ0UIkebt0Z/LNs5lHJzKpABmO
3XFysycFqzI/CjIApgKwdVGitww69GWiNm7hT+hxiDLZLHzHY4V5Yb7NBEcD
M9mbUz9Oo7Qt08IvBjhnWm4Q92l3YRkvVuAY4P8mP0Rzt8WWmzUTYqooa61h
1bJvSnUpfczdnI9SclDU5Qk8GYjUCG2TIglAAWSoUkM64KBAszzd2FH000Vf
uJa/yg2jZD7hHqwv5KLk71u1oCEgEVbwIroGgbGTZUTJfB8hT8StcmgtByn4
n6+xLwF6gk4DPnFLa2qC/2S5brIqKB5MjFHTwfMggvn3LGeCFGU467GW501y
LWWjLk52Q94jOP5nn02etV+ArqjGTEPTrJcmLVVb+Ewc8YgCL55rrEgWNzVP
FpL0k7koZ8CiNSe7R7bpeuJ5HTvafqHPoGj0AuTd3qWgc8kkxwyINZYh6/c1
8Wm46brUnjr2WXeZOZ6LTJ9VRMDrc4tZD0gI/oOwwalzFSPoHF8o2Z3T9Q5y
jrKb5MSvUqnDRshPF1mxf1LQkrCPoQhTkNN4jX7woKhsVFSJNwPUUNldku6l
9QHxWmlFNeuTUr2svm658w1EiPR38Tcu/NflQqvKnLKCr1QIYuwacqWVsVoA
ZIU4SUu52iZNyTrdML2CgObezCTRRMgXunnoSAKUEjlMtgACL7P1GNJjEZZ3
JSEOc4rs/JxBfub7OZRdeTpiBEykwBX8OBeDPYqOhH0Gw9dOkGAfkCFy/dMF
srKitB4UYi20J8B6oEG2LDj0DHCQ7NV4PtZs77rakrZak8xUual6OdNOMO6O
k9ELmhvB5GBCUU7mgTu5VYdPD8bnSEi6OU1BBNXmQ6uAdhEOugcKtehBMnnX
gvC0fDR6rUwoiLentIRdQIj2qT4FaB+KojQBOCR4ew0E6IN9R10UIuzLDigZ
xQ0kHNWPP73OTWUT4JkQBE0Q5ZzXlbtfMXruesDoVuRjSyltpvU5wgZsSko1
Ac2TTMCht/SGz4IqOTGsoptXBk7nKpfMgH3PX4NUx8tkFKWOXK7qR7DvOcth
tKz7iVshyX8DfGrJ22KfV+CeLtE6NRwMfUOql31iQQOvOvQVRdVpxubddYX2
UA5hdy9QtSwpeD5WbNcgdHXXO9+v/xtFIArZUZYPrNgbHXGqQcrQiAP1eIlT
LcIYqzxfMg5Dxmn9+AAX6ybluefiQaxM2sZ7hI/NQ3HFE0nPrLiUJs+3Db6q
dwsowSjNIFj4J2RVMuxwOtnPAMp5qFbqwX1YpzUOB1w8Na3KtO9DbBBgVc/7
nc9avhjfrngLrv4uvf1W7FH5zaCNWZSnsruhP36naZ6ofZd8873GRYCQ4YNQ
q6INWOFtYSfcRie9ivqJ2GhNAKAXhkj3tRBjs74iH9QScoAW5dnXRsrS5jt+
BbrIbyI3qGAzYPCZV/B7rYEo6Nt8wwc7M7A1OkBQ+Y09vHX9n+jDcHR7GgEJ
egmck9aBieNrAXt5oPu/7xrueuKXLEiPZOluZtsNJ9LjIlodJUlMxinlcqmY
sxKTrm4ODajz9KsRDnfLIdA9iyYPHKe/BVEFc8wpETxOG5IxSuT+VZUM+xe2
hH3Pa+z4oOv2c97juLwuGmR1wDjhUdXtYEYOx3RIMd9Wm9VC47QrSO2xXcIh
ERS2kj+8aAgbnq8kzSJy7TeM+MmzlciMqzCIyZlmWWc6lFFpn1GmBLRy92JO
fU1P6hA0eZtofDGgdmCphxiNUi+u8Kb326TIrYizeaC5TxthsAOXWExixypw
YTGMPDQRPmJXBfo0urtFVTVkGzuxoX3JDL//C/5PHmc2HiBBGQiWbXOPs6rT
KkQw4JdVWjakUympHIvBmZqoexyad4KeXLP5NEqSt5RwZg1XxebXmGUSWWGJ
0jgIT/0DA4gVMsVVDDD10oAeWxsigcxsJ5r5D2bFL1MhmjtJ4uWi03DYimWE
f61gRNnq2qBcyz0Ad4uzfyvg2xEcfCpEEeoZ1pjuSGUSLPe3tFR7Zmh9ywXd
rNO2CS3MVG0jLKUj0vhuWjm4s1Jtv+q2LZFzD5UFBPY9KC38GE8Hy4B9v2RT
ebL+LhU2qHJlkVwLF27ig0UnjPes5vVavzXCtnI30t/X1BC73R2znEFH+dgl
bz2whY9QkjBqOMH9Rah2FqwZ5Xc3aHSCu3kQf75VGwBkwpYwifycyFI5+CNr
sEmUxPhmtAiyx/GtEngUBfdqr04dUxch7o58I3HEmdJfZykI/F5tAMkVvOxc
mExUjbHtY7zehGbUlZQjcH8vThvnCQxHUK48bRwpjKQY2BkTUz/pUfjwo30o
h9PQPb3O2QLdRXQFcX89cGhJyG3IuBAvmiMyKOZRjCGbTw8kQU3S4ail8VbO
4/zPnWz92i3IlwxzQnFXlj4ynHO4DjLCQwXdgAEWDQhRS81ENw9JKBdQrcls
kg9Jfr5MQS+BzloC5oWMQu3bl2pixcNYCSseKkyFIAb2p4AooSR/gmaIkLzM
dUDUmfmHClO+4IzVQUN4frpa/huT6yckE8Pz/qp7kkd8K9K3mMBBnFEJchss
WZEUFUIwC8Q2y9Lzguae51uerOZR8Npuup9F0RMvk615nLlDd+qPByIMGy+C
0jQcV49EMnzYEmqSkWvgb9z+6T8iYftEq9QUxZTPK85hpM0BnovhIAHhnGuM
AuXu5UJF96fAuZmfTagJS4n921aDW4iWtERsknQAHaoNgps3XQSrmuGLF5EH
+GwxFO6kmq/P1JbPTkBh5Uqh90EQfngWSBplvumYu2WKVl3dRJuVbqv+985g
QL/rixwkp3cpUqPgV2bU47+esWZU2jyniUP581a6wqCJI42Llbn/OsHCFWo8
HZvTAcQk3wjsOGZp35F4ffymwkyJa6a7BMuISh9nP4GlkgykZmeyNK9RPBdS
GD9v2Lw5+olbmCt18MFm39dX+v9eDZM8Dc4Hw1yZmRkicM54Bo8xhw/99iXt
cGUr0uINpfsJrDWGZ0hpf39brasdLudtqoTVbiQViRxD+Lm8lodS8zTsMGwP
wzfUzt7ASowxZT8oM8c1RMkqsjAvxctFTgAwDut34/1wLuCQ3eTUaP8+RR7J
AYRr1zJvWHMokFB4sbflaMUtRnRM4SekvZp87IZkcCl8BYjX4//IB9MR5rKY
+ftbM4JbfBoXrUN9cxfE8nY6/58D6NgwDhSPByVgqA1Su2+tsAmLL3egcPIf
thRp1aA+RnjVNQzXLE5BG/2ScANZMU2UST0gmohBR90MOuI+SZcaKS1BqJhz
Ri/QhIy1S8v8WDw7sgULN/RGLFUDObH5MMQgXQsZ6nrxQpCfQ7PiSWvAU/uU
8Dic8LAJVByKwTeQD2SFd9i9ozPKxeD85yfFPMxBw/yGHukZT1h/jidwkxZ/
kx6UTsBdCqs20MNCopbG710K4RKN/BcHgXub7GVvimy37aPPlXcaoX5XghfV
pBSPpWR8jwQvAIo9nnqndLprFRyKOR8NPUtM7ab5iPRVzHGZytLonhQ6V8yr
UF1k0khzNbrww60OV5VNy7R9J0v0ryxUZmsY4U4WZ+pnNwuPs/658qAfW1IY
LZAMB3/Rt1W1cb4CzXmbjvQYc4OBGg6Zg0z6WEuNmCptTNNxMR0b2pP8O4jc
3xon1bZw2T5tKI6/LWHa4g/AHo1In8Ujtfh1EaHu3QPkeXrLkG7n6SZLC8YG
xLeu6tYVS5xAWYzHfKT+CX66t5qbgaKURbL4KM50t7ubpSJsg57y/212gbbE
C79Ld1h5GC0pE0/JT2ojiRwXY53uZbg/wvCk8yS8LePWdkjFQEYlGTPCx1vx
d5PbZqdrn2MR+h8orbkUbI8sRHVDBlRXsK7O1+7kdNEle1MCqcsxxLoXt/pt
VcuFEmMf6GgIzXGgG1DQ3Tx9RsOsnnrncatYB4pEtuDIMekHnGm2IOlg20uZ
Ii/c2idcLyEAoQnrMJy8+omODcszV3hOJSqWo3pbseXo+oawWlTe+w2lWX7h
nqDzIMbkEyJvTReaEAQeLAL73HGM+Lu+I+27/S9mZQvaqYeaOHVJIOfxdyDV
b1xFe5HRfHtBotM0azXcm/p/uqAhd6nbaIsGYww4Kmx+kDHPs6FC0W5oad/d
Q6uSinGXxJD/tcYayHHlo6wlysSANoUuBjw255m5jIocZduH3klol4rxiTqO
vr9jDGKbt3QUSxXe7VBeCgVJClx6LVYDncRsL9uh0DwJpKvHg8u5Xx8i7TRG
uexs2moHKk49rsOBru6wtx23IdsihdZ58fZ76w0AUS2nHtmL+sEk6YQkj9zR
OBCUH5UV06RpNbpi4v4tuRYCCN4mYhwKY4wyXn+fU1B/n11tJpV9rM5/RP7/
nHLvYyJ6l3VExQ8KYXrOlBI+Vpqn8EoeLPTjhvjK5MOChJktBI/abvxkwN7z
cst0wBLE3s+XHAl6hZ8jn5IvOBj3gL8LbHdTeI3hxd+kE+xafltSdWFProW+
VuF7xl8OwQLyukGq7SrkMYZNvBPFsWe3TTvyGGe40Ji/8nBQOhHUP8KPwJ4A
jTWo3I22YWvn4jwvYte0zBwG6YFAT6O2wBGxepbBvm09i0ZhWvyc4si5bYzc
zI2tqHl/zoiVm+7KJbM+WJG4HmBhOEJG+6l3RUY886e8HOgsEkA+gEgDo65o
/0AhyCOtXdELsL1ZPnl6mStCDS4UdTXrUuY4PEFsUIlLpNgY2hPImEx9z8EN
0qbQZy1X55EGBQZf5M5Vxh9VQ7Jb27CmdTA3mYH6PUOI2Yj8lVmwLfrxsBc1
iBVadK2LDyJW24kFdriHq7d4ck7jKameoI+paFwT2Zp47mDSPxpwkx7glq78
HDZVJuxLjn7juS0DlRX1IrvJjjTLWfQQNdblZzzoEXdsYkRgEKgRSx8rBvXt
+LLFM9vvj+eoW9Qjhghr8wcadKCjLRQh4VAdV1eZ/hYYsYmwNsxaE07l1PhV
0XKsZkdFyphbgvpO/RE9pIBbVhrh85LbHojr9RWYYbAeNpj+PzPfC1ocqQ1x
gYj3tQgkbvwkYIDk7hE55pu4yuvsOFGVcWMbRunAIEzOZiVxGkC9MzhNfR/C
VV2MdNyrc+00wbDDweYg0s5yjpIZ3i7Eoeh5EO31CghvHVwL60sQd9kRSXbW
qOvfifcw6Bh0kjeWXYx9tUoogcu0NlkyO5vB1TpzLXy4jDjkAZq1ywwPsZ9n
ABSrhgfqLYylX1hE03CHxleFzJhULdUoWNXfXIfynO7XOT8CtXbAyeDKH5oM
2nNHTdxDcNcqdbgo+dC+lEvMV7rOlNJNPahojHq/7+NOmCmb2+O+G5BpD2Jz
G7h96v4zmFYxj4PwZsga+W8Wgk6dNFUS5n4HgP/+mRI7Mwu0hJtOJ0c4bA1Q
jxAGuLGVNAopDHS8VKY/JizmTBrLJLzrz5LZXrJMV0I8/QnhCf5wpsHaoeGY
BYypeb1Z7rYskUF2f3tUh0wn2nHD2oONkzxtISUPXGwfficQaGwLWnEc1GL7
8vDdcWJXD5dkelS5gjwGL50qDflI4FkdEbsR6hqT96rLppqaZQh9C/hJPnKG
K2qOhtI5c8KPLPdicdBwQNHdm/pL+yEVCidXM30a8N64SdB+BYGaQkWW5viJ
nfoimkfa6q4453lMMsT8122hrUspKbwHAsarMS5J/Ee+vcUfDQtNrfn+wOYx
fd9wok3J5UxeRo8W4jTDWqgmfD3uZP7oJzBZ1PPBrkjhDGBCGoWFpGujM6Uv
LegaHmnlBLtKyk6GdwrWqbAE9xyQQk8feydmaYCf76jusWA04j0t5apGQcWs
8WYUfT1Hm2f7mkJQentvXGHnbuWatHHVnwGnVnmJ5yb0R+ts0mNEhzYe1Sem
8Fs//pn++M3I577iCUDBapLRH9laNLBMMziSwqBLrgwyrfcWuJKkB+CxAwuu
dpnhsXD5whk9incb5IuM8rp4lHEq7Gpc+tDCZBeNpY9fi4HS9RpY65cZ69ml
kgPPEv4CXjxQN5modtycV42fybyUQCcHAxUT2L++UIP84h0hJ5iAtvcZvHBI
Sgq2bMvIe5YCH8tvEpEfb91NjWtB6l6noqqPLQFZTUKYwok/cen8Ob3iW0q5
9ZuYDcEm5v5GoUeOGetd6lN/YcC4TIucamCMoWFrB/h2KPqK8I7C9+swQxSL
mpoKHeemHZ4UuCAIKW3LvBp9z6jo+MocwjbLTdGMq9NFG9aF5ska0vsIeeN0
t6i2cpqM/4Nye/SF6LCg22RHvI+w6qbx6QSJLhH222elpj56wNoIp8xV/OEz
ArGRE0M6W2eM6FVLsFm8+mAagef0qdZcZoZe+E6yctE1AAzQZfA2yXvw/RJB
oOdmFAGGeEDGWxijfYB/17kpwN42omFt4Y2AyY2zLRZiPVe98+ihqExpxCFb
c0MhPgtz/UGaah13t/0QoihohP2wwRKzBck3FTxP3NPrvy9yD6Y0v1ZgoeLk
KaMttVy/P/pcnJcg52XEZz3K7LdTkqn4ZD7J7deF73B6bzCYPzbYV6QuUITS
fTlhcuQLh71AUB5UIm5n5wRdPbP+Kve4IDnmejMJyUv2cq+1R2AghGJOSV19
Hf5vC9K1xjCQhHoVVLrkKROPWyoEObTdQeAU+YbaUdcu1cqlIP6IfIiHuPEm
Z0I+88nN9K3Z8DmViGxLKJ0qTFgtPMPjfv/HnK6swEpgkaxxcr0Ax3QGOq5Y
QM9MCH6L+zHhLk4YH+lTfjgXzMVadJlv/lRqjB/YItGCyIYzREUghkHBefZl
e8hKYXLffNAR44NW00FPHLqHsEVnYMwEPM8QXs1Z3aj8jaFwO6psT0+geJEd
T33Ke9/eB8cvflXEotjKrTFNX6/EcwRqMwkZQlPpzyaxEoVEd96WIoDs+ZCF
R5jqt1bR0gLG86Tf3AcKHisvfZ8JQ+xoX+kAaQ3MxNtXBj8SwaFiaicjjlxL
GL+T5t4I/TMp/aU/i/4Ch5aqBM6lUwW3adPud3mOfGrvq4Gg9q5cQUVGDfc8
h6r0W2+eCeLd6Si2V76h/gmV0l7hj3vi2DGNyYuLldMidejzV664gP+1DJrw
vcpUoEmW12kPzhM7gxGucYUipGQoVFxAMqZ0EnY8Filqzic0m+OdrfLkqqXu
wtKNY5D0PtpKyEJbcvr4pHmt97IKNdG6uVanx5b37sjDu0rQ+PWLDJl3Cp+C
JtM+DdOP4XIWCFLoV9YaSl0jgDQEINOXU1zjUnbvBAyCCu70BzMEPZTLHrC5
Y75bcFk5l0pXKxi5HDGnsq7EK9QZdurpdiS79038hntvEIsORX/zgDDlaswU
wtRMjebMbTI76riX/OvnKRxIGDN0dzVY6Y60tVDOqCbwNprwuDHDDYSNG/gZ
FErkY/Kc07yQwUYhobrOpDN9yZa2veCMIAo6waxsOKgCH4ZJTnPn2Xoku0d0
21Kvw5FgCKa8fGLZ1hIuU2tI+qNGhpOIxIqmR8zwRphtdyfXi78meog0vF5N
/nBiOyMULB/3wQkdpHYQWYake7M+YShRlfaZv6HT7cztepmBnQmUKZ+slolw
2GSPhZbxbw8OOHEb6qok8wb3eSDBeh8ZngSv0rDVHs9+XHBVF/ge6yPShN3n
YAgB9D/VKThUDwdNPo4nWy/LHihRDtA/iVZLWeWHA0JYoM2P1+WLk6G/86+m
YppJ2ArPD8/Ffg+l7ax1Rp+M1yKndoB5ub6DOTcle+S7XU0yq1kpUKdZZ9PL
CZHm0EiiVZHr2qMQI6kTuSQ/tyC13TptnsPwPYEUw7budUhWuebRIGyLjTr4
2npnctNfOH/3dLM5JIz4Pbxviej1iqwhbz4azBAe0wHMVgIyP/foBWWLWD5g
VY88zLu1CsxihkQ5c2WHwyIxyoQrRAKugu5uleLt4X/9d1tBdsZsNfjxZumm
JTNXMbvZNRTC8cqF/Es6rBKZKQpbTuUYLa5L0AaSlif6Y87gIozd3mysgWZL
Wovd0zYrAtZS/v6pFcLv1w7pNkpoDVShWwT5JM9mcZLIEYvLlcwXhO4X1+C0
JWAXdK6QyUoThDNmzS1HdZiqwXGZyeObZtXVwCOWhTSqxiq+jPwAeQpsMBQz
HVN4gPSvHUTVv4LhuFNWZyFgFgJR9o3sKR9r2rkOg5p2BD2DSIDXZxFrnQCD
mRdOt6K7Vrr8uXXPG+DeOc2a/lEzmcOjVWRa01KfTTwVob7uWJFLioogqNcD
iieFhrtuq6sm7NJ9FRzLYFRxQH8VlZFbZcCDVeML2bF3PQBDgYIWf42Bkj9L
QanwHnZbBMAa4cO9K782lX1LNYr3Ui60iSooee8D2zVOj5Lp1ROfUD6mVBBo
VDfrut21F/1xOPv0MpdEEaxiohVMeh1D+MLLGOC9BkjDZmwCz6CEDfWHFvnQ
JTbf4IePkNY5klXCGOJlNpwxDIRUr9m/G5agfJTXOZ9Y/YMK2LqGrI+aO7Ua
0SWNRws2CTibQ8TFJyBTsbMiSPN182hbUG0NCw77iG3hYYWpkWfQZx8CyJnf
YZLIsOssPWNIrT5QHz6SvmLXB+sB7+apS97cjI07RMLk3XBwI+k4YIid/np1
HZPKg7u3/RXJzpj+7CjaJexpERuv3x9rrNusAR1z6rKKhZ2/UTa7DQkYHlmZ
wEfHEsw+E3dYhE0Ds+UoaqRoBEx+k6sqmiQVyqIpl3rUkUYxrPkvHdS4HU5A
U5rAm7veFUnK8u0UG8n+YAB09NDBOklc97Qtec3JZPC6I05kkUZNZE0cEu/U
P7MnbF2ENknoeVAzv7vFqFDjjNvH4wN1AEGVezzZR+hM2KNPjeMKS0DULrN0
jWTb+4IyObsVPS4uyJ876/xLoo8M9L/+aV1SBS0ey9q0wcUgoIXbVigyoVXj
lo9F0aBwFz+mh5pcSx//c6vMf3xXxU3hh8I01QWyXuwywdmQEREA5/s98RM5
xyAYBsXADDz9+njDXcHj4n/4vQxQpZ466vYtfjKZEPiRPRDiIBfyfsAmDfwT
XH9Ct7AgS5jnMFU2qijOch5UuDz26Q9uwKhi8M75dFMumq2/sLjfQay9z4QZ
sT2qHN4BP2fWbEpZf8dEEEaTw9UjMg6Z0dFA2Q4VllJJBUsIsOSHTFDiuRXG
gU8M+2DNAzjFnj3ieJoHaKeuhtmP1VO5DrnRwmUTjfXyB5XyL5+ryYB0GgF0
Xa56TZa1arWk4dpilXW5dhCUD5tcQ150FyOzfvD2dQ/PSKfWuQWa7s7iU39L
b8ZW07JPsFI9ww46lfKmppFEQYUoRE5gTaWFUXOUEFRuEf1qeat22p7c447T
WwTXDpX1/oDsLWOnCaME30eLoGP/HAarvB/YdFLRDzoWuyTKb5XjsKejYOyK
5efKYvd3dD4NGViD0kl93lTUB6vdJe0OAPGXQ+Q//53UL9ldHPyZSRSMSn+I
vwYWoOwOCDPpKLx5TpM9UwzIhYhKrbHfipFJ4u2yJ1lPoqBZ9vV6DoiENLIP
jvJeaCbBUfWd9Ozd7HVElcT7yMIjP51sD8hLkZkpPDq9dZ+LzZZf5NekGjSG
IzHx/jtmiLbG53xGv4DSzWxWzMf1oJkRbqbjuJgVvKf86TMKGI1zgbHaDIIe
e8vK8AeoSAAj3p0cX8i/+0moogDYqpGj0CEkw6y68TwlgI1n76dk2l8epukw
/AcmOqIjoCFYYjFUvjcMgM34WgjicFWE2AfzAKM4TN6JWSdKfrNuD1Msd/ZI
6QdEvqhem0qknXoaGQv5a/9D6dGzMYe0m2lFX3tjEFBsOWJWSR2S7Tf4y7h/
rSEIHub/xOoFBtOaCzENkS4axOh20krT0qTnZ73tCAlCxWASrjakYOp5Jf4Q
aYedeAwv0GxsUiECpfQSP3jOZcE3jmnTnLlhutN2wx1VtGk8EbuZFfixFaUX
gIuBuLulnj35Uu+Did83GsWFEKnr7NdIyTgr+JGywZATTfR0ZJScv9JiAI3S
hnCxMueyWZ45Srg/7Tho5438IgJA79RIHoZkO1Hh2i6pSjVO6LeknLmTV61W
BMspuAC6ItfiZkOKUdNncIU32y9LpP28cbbRHtTPeHX1j1I0DVxzUQ+BeBLn
sE0IGbWwTE2oYoahCTwm3mlMZ/MDmAOhSIavNjIymlm+sQMlPxuru9tTFDbI
qrWVrk2fhsAbfNMZApGMbcp0r4zeSt2kW8VxCcPFIQuTRXYesN87lZDv+q30
a/OqgL18D2TX4wNzFwWgmxk2TWuzauDo3iJZ2X2DXEAk9IBKdVlyGgyrSJjr
1FAJWrPurZ8Xa6vWVJI+neI9rGX0YhP9R1u85+40Emiak0S6kgqOIy7EG5Ev
3/byWXlILUQb4dbpyFEqe13SBeWzLeYRSp9y21/ANn1O/Wc3EModSlX8ce7j
nZ3vEd5oFnVk/HTYggqc49Y67NLAGze/G4TR9u0qJg7oFeFxTDemegBASnbl
42UpO9JXpMOUXbuQdjqNbpU02QBBTlbPJBSstueOuz2Y0RWA3c9pkYxCdR13
WMiCk8UnxPm2Os+iA8cOskZ7B+fyDJVBe9F06ZXs93U8Kh/1REk6jvIaeA+A
wVIVsXCvLvxVxrbztdvPFF3JpnSEbViaqlBK47yC9cBZuZ2/oXetvgrbopqU
/wS1isdhFvua9izYx6/5s9C+jCZ++iFiPEsbEVmqblwuk8FN1haT9UMgubXo
BG/0AkWQKoKf1atEnl06ZgiGV4z1YdbgBE/TD3Y1l8TIjCix0Au3Fy0iTbKO
rOQYVfSLmg9AYyCQlm02ZtlCN11I1i3QIjHjSrlgbqB+/IMBr3yRMFOoMkbI
piq5+sviFtNQqgWsoe7ILsfoGa8/jXBtIKKb6MARepvNFlsaqSgkFr9jUX3+
RD/UrGH4ZWgULk/Fi1w/WIl/OhfMSIOlFtJWGSoiVX0lpbP4px4TWvatyBYf
SIZJcLDMdqfambJJ4KmoIRpP2APse1iGLAeD8LVBH3UL9RrmR1NHYYQt6dUA
DNq5z6eInwF7Q7TU82K75Ul84S+XrCHQxrd1lLLihgIOX6j77p02+dyBEw7x
WgpYLIfWrDay6880ns7+qsSIkEkttfG5bv2adrOHfDEm1jXgl8bv2/yyWI+9
u1+FFzRW3yc1KeIr9S0WKCuW9jubxBNuLW8OwsgGQ8VL+oYv7drhNk6a9uO5
0jCC4WLhQ5TmLyMHf56dGRl1gWUk9AGwn4YK0qD6NQbeuM5FfXhVyh+oXwjf
idwvTW+hFWKrKj0eCpunNGhqmc/lq7kNvy3aioD2Ts9pehXpiI7r8gmB4hLE
87aka98zHF+wmCv3D8QpMuxYLiNTD3Dh1yGZa6D9IJCKH2ZIJgNuinQMOQR9
Wik8Ot7FuwglsLucxwo3p4yqnyj1JB73Xt4SpuAsUKT9uYPbSclRoNcTREq9
SJnd38OGUe5xGx7vCDQY6AxvuFhz6AAdnXLTv3c4CVZEp3XXwjoTOyIc5X7X
usKepcYBj/cygpdfDTV2vLZN7h9Owah+BHtogzT7llzfsQ5RVFWQfTzjI2B4
OwX9LumbB6qWXwA4se0ZUVYFoV04GKeu9bWixorIFv5B/nugMk+YrXZXnWtK
0DtIFQXG3rXMqEA1Q1xh5NJ1fIiKArzQ1iHRA2JlZIJhoPBbAtje6EKwQOrL
9fWLGUp/wAkrlhc9GRmReyFLAqZZRbEQvJHHV/XtKPent1zDgkNcAyyBQi6m
9I3cVoSx44NXXlaYJv4eOSxFa6T40Q2iGdo7rbLvDrfElcENR8u5upUlPyeg
+ebbjNSquhThUFdr8ahHtEMNk0HHzWG8JQ+63J8EXEQ+CI0RgRIcoYXPiveW
JBdO1oPZA1346F+S9b2ovMNYlMkoAMcb49FInojbU7zJ0sqD8GK3zB3OAzdP
VWbsyjQ9ZC+H+ebLkseopWX1XHYq+P0UEU5yy74y+OiZxfLW+w7SwMXp0Ifp
KEmcAIfII5r6vj8vcCNa13at7QQzfara+2QVzHv0kI6lDZ7Dica5K2eRbZDv
pQKIYK+qHLWYqSHGiSlrdzvKiSYQpDhkoZbGBnUkg8HusofCPTugXLAl7iSp
VDfegpaMheVel1BTG6qbdPBMv2/l/0zv6OuCubrh/gNyyVMEAlDkx2jDXEWV
vnfoCqp9bwi18ewwkkK/X9+RQdpmXbfMUEcmcV8KiI8tTHDH+b29NdFosw+I
emsJ0R0NbRxfQfJtF3rJr6jpsTfufWF99coJ/UaYAYhy6dp/GE8SF6OK5Qkq
PoVCw06GEjIJvFETG8q7pOjx6zdS7cDQdYtwoPbb1x7u6HuVn0Qdv+wUvb+L
Z5U6nlS2m/zrxNPeOIwtKvHgbminCRWl65qBt1hBaIY+/AgWpiHaXnZBs/ua
7iF1eo5m1Q+nrLZBRYSx1UgkjqPvr8iSV6dBaxQk/mEu2tQ5k0Xq1NP3qisN
/B1PDhr7trbds8gCfhCHTqiRWqelcnFs12WVJzU4HrhEjJXJzfhFCi9Tn30C
tnFys/rt0NecyropFVFB9Jlf9z6YEVIqM3jvkdgUk63VZGlBxwmEUcyf+7MD
pe6g7Dx+wjGBcKRgUt+X5mn69QKldy9cq4xqCAkpNdz+qt6S+MH2h1kIVjNm
4GxNTERsQCIBboA0cLPn9LoRzD8WkpfLX+Qq69SK9E7ey/c7wK5EK0IOwUVO
LjkWp9Wj6CNc2c/dbMP/Kd86uz/htsN4+iGfnUQ58pryLEnArbrcJcRAd5Hx
6A3FKdClhxXtbJYeh8MnCCqRvVbeNzpTa0PDJQEMAv0Ky1vBjaY8AGmKDjJ2
iNWaWJFtP18TIYIGlQx9Qrcnzi10Do0JonRJpWo3p77mxa8NeoyXIHsTqwK9
cPQQ6rE38rkHXpW7o39W9PYFcki+C6sUY1ahHUgesT3Hcvxudt1XqMSjPVcE
BBrPWxmLHM/UXIrnkrBxFWPzn7MXOp6OP6sj0se5aa+ihPzhYWxoq2MwIPvd
ulFm8vv7MakzUa5BJJATtEotzCWznHTPL8fU0JYPMHM7sHIKA81MRnqJKgMV
SAALvJ0m07vP0ZRlqWcLZQeiN+720c++hHGR7qnX4fZ4VKgDQz0GwWPQhZVK
xFMrKlbuc5ZwgW7Qy6pUrVJjZVH/OEGQIemr7PZIAnLZlVtM1kDqlLeN8HLP
E/JNr+yfgVUsO3h2b4lS0FhIqzi6qL1LZDmuPtdpx2Rc0zDM5ZjizhI+xPBi
Vxzw1StAW2j7Wc5z+SdC3QlKx28iJ8iP+b3jmCD3mtFUoXmW3822wbM5Mlrl
Kbc1oo4fSw049k7fBXlQFeF+CFPMzI+/QolzWZymLra27ZAtrJ40bYmwJMIV
6YlOa4XGknIS/H70bZLZNTYfuiYYrg+8fagBoG+K2StgNtvYtF9L6I1n3WQk
vFYBpFg9ZR0gIqC0wxz2iIhQhNphTMCZ5auLgRE6GWY4uueau2gyDsVY9Mcp
U3U8eMpqL1uvrgXtAZhszjJsrQg0nmnyzlmHtiHnJ901eo3gnTrIYvqMY4D7
knc1TYtolmC+5Aq1SVd+OtZeko/99+Cxk44ngvJA35lnjAsx4DVgPp79o/y5
lAXQaOQGv5rZ/vu77vIxVBxHcdehKj5AhBp+CjfE4xZRqwgzDXBsdMBJ/uQX
NJttsNBiL4AOSOnNIyZn1ViwmgSeViNM7RSyrpwd8nVdgi/bteGCTGqqMYKs
xe3XZmx434LY09tXZOfYzfuN7/Lc3bosWs0vGbZqav2XC7VrcGOS/FN080Mk
6Sj0JRMl9fSaV37H70plV85MXDfHZFdpT2B/NxGON5Ykpw50LZGkOtmIlXbV
w4RNh92/9hQlwrJiR8z6lwUSbuUFF83oA4FxLezbsahS3No/2Lpn7d2iuyzg
/qER5KRaRAxkNSVHaDuNH7zVwi5j9oLlM29fIkt1d9uEGzTsYN7XoIGbEwXr
x60W8Dj3t2zfc7XRKU31d5jzKEbQaS3UAa4Nq6ogJ05WtiRjSjea45xEOsnG
bUE0H7mxkQbbW/OkBnS+sAF9ARBglEFypy3WhkE6nXNgmjrvGibgiPAY3QLf
gOjToPDpQOw8PGl03bzGVzRwEknJc+pTW0xkcH/PBuaswCWBUsFs0nmO8Uxt
/6JOYhzorZSaX7/2Z/m/Vs1Yg49HPQ3+QkGrPqpI91aCZNBkNb4YM0fiPZxp
ZQ3SeZKE1cIPpy+ubrLCmoqc7SR9g/YVjxeXJiZVzQ4epUKDP25GRUokThQB
AbNp3Bu035m4kRqSPWYEGW6llTMZinP2eDkjC/4gEVbMMWdnxFMazSUt7Hm4
2JmSZiY2brGArvd2VRLhYW0FQwrI0wb0hV8jUFe+gXJ12D96taVcYXPgGwY9
mp/KOlCbe573A+dYYR0PgKCGAxHfm6bFByeWf87EjiUjyi6W45TBs5YQnryV
FIAJVslh4y7iHFkPJcOgA1lqu7IXcmfAOQyzxrhmCIrEmAU07hcr79FV+E5+
wjkvNqLmBBX6JOx6frRopGTbYx+R5y5JKHMi8HGpLggcB3uzVzKM/d+u700l
kErtTwNfrX1GTpD0WZLkV8jjsLfCvuuE6UxUVkhKiX8c+k0HbLxHX61HOsXm
qKVwUHV2Px/QziGRM2uhmdru14gE7TtruTJZ7Fi/kN9xNzYAW6q/Q3Qq8xLq
5zGM/3ZC3i5+PVKHttklzxw8BLaENYZoGgxBJP2JVkTZPlPb60d7tSRZZ+Ce
kZeALOSujjDnPSk4/sXHGZdfCwU1AYinL5+RPKWYUbzxtm3zon31FU02y4h2
Mwe6G/UD/QEEPf7j/D4Kw+rnJ8V7fN3cpa5I4Xedk/H9rX6WcYV0aikBrXk/
in8vQaX7SitK1Hi97Yjf2AD5rBrP7Pl3j9MkoOaCoj36M6Av+7MapX7+OcA7
5aPjJnRB9Lc9ynMhWBmeYSHX7THSygbJnsJDYEyZ2CQoKqVL2DqAQJxD4RNu
k0RYc8QYK9UwWTzUsd2Auaj5FNv5eCkzWQo710QOmh6zXGeQQXlo0y0bE0K+
U6iodQbVb6t1o9Mhq+l4uUQby15Tq9SqzOl08j9WcCGZozb3LW8YIihHAa0n
uCHoLKRW8+alT7pbRpWA+MKNgtGdJYHfEcxDyl3RF2VS8lr3kvwAJSekv0e6
rTZExTXLScsj4VYnOnWHtALT/MYbnsBD6899tyT7QVnFOHf254NgbQ7NWWHl
lCZrCYROu/5JkTWEVtK6MotE2Obo0+bYmfjsLDCYPZ1bx4aciCWKeBeJi7rz
8fE0SoVWoEgHtsoHwkXVZ0THOxeq0/5vqbjJNiAsbjTXHxVkQcLbZWGx6Bs1
HEJ/q7+CnO0xJbFxfl2xk8jwiLz5yCd9ZcTOkmS7lCZmiqAOdtOHA0bkvZCf
NJfabvL8RBNZccZjaZNXUuTIvr/ylwuBCe6pwNBOHjLE4NtWOsxzDjHcd2Lu
OliabagoC4T1YzJQiRSzx5VeJOpSPE1/JelT6gWIwl19EgKVjuyTp4YFzrqV
qR9Op5XJ4trZRcla4IGL9hYXNrzcgTk1cb1slSwsdiUqWHukb4WLJjbdDcip
UnZ9j38+md5vWLI51M7/PM6XUb2u46Fl1cDBXIpxw3Lp5ibRSurxhvqLYILT
NSP1FKv3nPQRQyHp3ysk7VgEnS8kECAQ6vwiMbLcBNtslam1GzV19380u+Mr
8UnvEZeiYKl/2E+PA8wz2c46cRBJqFbfoiRQkeAr9frEakbqBLP0+fQ9SQwr
KN5EXX0t88MjoR67tACqgwYvd4G5fHVU1JuYMYCy0O58Tlg59HO9sZ3T600S
6YmZ7GXpGjJFRk90NJh8Fju1v5nqdCbBgerTELTxPejfLh3r76XfBZgsy35a
PpnMnvr6IIRRH6RkwKn64Zg6y8VGYyCD4+v1gem2/iJlHRq3+6TJb5YikWZf
vDXL+/av43fbYpkIS/PWq2VXvhMDfpYqyQfYG4l/JBWdSDHqSLbeuECIsPyy
sXHgofvygXiDWVotQWiX614C0IEKuD9/pX2LUbofsickC1dGm1VtgxaVWWhM
R1JYRvWOFRumyNt1Y1dnNTlg9egfSTC6ObmciCba0L8Mwrzavan8tM6BiEVK
Vh3G80LjHTqLmDD2KX4yHQB5zbr33+hp0lyjxhbwnjmhYTHeZOIWdwe6ncN7
aVRJCMlRktTvjH0wCoifD4wU4rVgul2v5AAg7bJymPZTHFTE/2AL6R2KShua
crOvgMf7yb4IuWRDsq8BVTD5X6sXYe4ezz8Wx2q0GKg4Qb/eKN+4B3Uz6jIx
FgeMzUk5VvxKgEmxNhp4ZhN7bGaZVKBJALXb5e21D8+pxsWLkEIikUCwyCXA
vQpRk68YQtliHL//VDpobt+Ct3bkcpEpwn+fU93qkAzDwd2kVmhrSNqCIUuB
0j0VZ8FlhNM4pS0e+rq0k73Rixs8SlaImH0O3IiO31l0/hVgzWswkfKv6ZPK
dsOlFVaqOOdx7R4O6R5ZXMTRNDsMxv0So0r7yll8lrSoodPQXUgodKMdfYRG
6b7xT+mkOVAnlopPXgJHJLCsr+ozcLIPgYQcRYpqyA40E/Pw6/2sucaXCdUw
vjZeftJ+jhpIL1i+jK2VYVp3Vj9kARq6ykP+yZd81fHu8wFhs9lUoiiCGWOJ
NVEBc64xpn6FxqFUB9rDWD6Pa2fgKcKbviZdDOTTQG8l1/tZ0g6dYlRwvJWb
O2V6TiQeOKvZ0Ulu4euZkdwS2Yxkpzh2A1PRI0tjB8mo1h3CCPZbyYhkklfr
40DlCUsheGZKhzFeT9wMvI+kfOgk2fVRWUV9+0+/De15LPmHW07wJ19tJ2O0
f0eFEAih6vzFsI6hIZ8yDwqGIwwh1J079Ep3uGDKKpv1bfbXzKY9S4Vjw2G5
nJbtBpr+HAcHDnMCFivfxwD+ElVCNOj1JDvC8BZCmIVIkUx3q149Vvue48lN
qHOeIdPlXY2ZOpP4FF5AqKA8ji0zOZL0TAn4fKYi8s10CNQP6/g5aACwPTAd
86Kcj7ECq99ZL64WIz/do3rC9a16u0/yPY/Ey7gO+p4m89+u8X20F26blWy2
04qS5cMlRhP04+1NH2uPMgxEyDK8rex3bcD8u8K1YVgxAotz1CeHnyX4R3Wy
1zuENPdOVenf7q7h/Spo3J8dunk8r9IQEnQcZcf4B0AQKg3EUVwZB1wcmQhe
JJfP89MGvmcMVGH8pwQLDjyOk1u3NaFhebWHvI2I6z4p0fE0yxVV2kSY+1a3
Qf1dzmelry3nr9FCd5GJ5aMWlaM1zUkJMcoRFpB/S9r2xvzQSGUsbBkFy7g/
lGt6a6se85pUvt2dyFOvySOJrSsDrGw2GL25oqTHfkacW93KW0y/9TF01/58
Af/tWcoHZAmeFDYYXffRbPsy+i5olw870wJh4XFNmSpWaxb3qRRV8hCXdmzk
jrCCBVziqtLSfX0nPeAMr8yr9MlaLo1wBTq7KrYKyYT1TIaNXQfqNT/fAguK
hb6LRSTUuFJeAUtA938HcgiRXej869V5thogU4C4mt+cfMU6txn1457moNb6
Lfs5El7vfBoWSsXCQLmnW771hqgBiry/kzH1wdwm7gGKjYtIDzAjr3EF3RtE
rFCjp48ptT3tFIaIGtqO4ufLzW5jq92CY8hPgskUDKBQOoQhZEos9uo1kgeB
GcZZnJkUZ22JUakY2oolxHR2mgfbYwD0iuW2ZtQCSN0f/JbKkIQnPpACkQF6
LPUS2Vdm/xwY9Im/kLnDuaUF+slnRYpeehK8r6jZfgCHlLAl0cRh+U1S2IDy
3d792KBcfgf71ttto6eD61P/fDHToW6iwuiw+lk7SOr/tf1V4MQXppPEMld/
yxklk7JpQ1qTQo67pPoNQ8gOuXrjT4cwokKaGdEFs3jYlK+YdtOPfG0jAm33
Z2Ji2M1YgMweJRxW4X+porwufVWCIckv3QQDGAcSYQTE8r7lNMSzV+TW1rfO
GZ+T3cgaqzLXa7hFRGd1kZC6r3ntwIp2kgXrgT19Ztx0D7Q2KszT71hShKzf
CUYLZR4OwzrVlG9fuSTsCWD3+ZY+fAgbzAoo/S3/8V1Xdvbh60uwj3HOjjRp
PInBAlcrI703JocGqDrJy4B6mqz5l3aEyJO03TMCDjnAht/AmDE0s45NBHqr
6jX9kDpPn2CIouZd8AS0oltJhk7GgR1N6HYu2TDCx/ljFZC0qqNZOfSIDPrp
qZn5VZl5WyLzjglWvlx+SR6rfoKyltFgh+uDCrZA20SJsT2Uga7sXG27lRMe
+Zb5dXGhc52mwEmx0OhKlPcZVe6EGP8aMKrfitUQg9YQRoFt7eCpXzwaMkgD
QiardZLIE8CnBZcdl3yZk57HMT3VXm6DekC+jW3rtXE3R19qgo/UyGFx368Q
Xj28ULPoykGP0F6bo11LsT57Tqp8yvechRHyJyOJMxMGSXGB+VON2r1Awh3q
NmJ4H/S32ag3m+PNxF5jwE9pqgg1ttqysIY7DG2sZ6fxBK8qGXT4NkeID0Np
t1TxW1181F3/tU7YEphzR1DRpNaOsSuUQ/55p0woWs47ZQgPJVtPbM3/HOoC
lZpB57upljE3dYY3FaEpmGAerLSw/jXNzANU9KRCDuiID88fY/qn5CT/1Taa
HoE886O7PcWuhxLMI9LwE1gVD+SyJk3mRpOq8T6d4wj3aQLoJuypEQQi5kqF
dlLgDyURqgIbUOLfwv5Q5lmHuJGu1TpTxwPjZu6cK4xnKVxb9YPvvEX9lKuy
HTGuAFlZ/g8Cln1VUmCiFDAOzNLfbHoZvc4qGHjZa63e3GC58A1Js01YYDnb
yty+cL/8ZNLGGczgVj3eZqHchPsiC7SQfNxXZuTM1WTJt92ph/Q3GyLy+3Lr
UqatDURz340isVM6Un4MktNhlZyWEaeenWMb635y2fGegGUtHFRcnwyfx76q
bEIVau00ZovRAbYy5jMN/hef7Er2g1a801l5nuBe5K8KC87m4fT1q+RwXAgJ
znH6Ee0icoQDZlFwjixbxjfysIDxdqnzsLbnTO1ZeKZpzufYDPYbqBB4Jhod
KESXluicuETbLQ8ydhP3i7ThMHuCSuLDTTKVYLXiiRAHFwSwkqdnuqdzyp/w
CveqW8i57/H+LVH5DLuEekFh3HjlpQCz6fw3TZFf7mtiKtXRaDOIGGPAUhNR
3MocQ7t6eVXiTScJFd+Q2mCd5dsMq/+g8Y0BL0YZb2kx197NgzDHbj4v5Msb
jBj0JpRcuv8Y8uxWwYTyB0FJuA1hKDL1tQsOmlPyv3wCDnwFMOohcWfweSr1
Xf2c2ROWj2DgtMS6xQ7hSYqr/vkQ7FU9JU2xgn1c/lctmUIEMJAlMhwUc466
j5lgh6TGw7ZpnkCa/ATF9Z0Epnpmu3gJZcv7GOF0FuSz9m0LsLIo+HCpOT0G
LCL2JkWXjtWveVCxw/QaVO69FveepBR6fwRDsb0NBkHcbUadgWiXErX22eia
5sFP0SQymEun/6qQ9SC7O9zrf7RuZc3tZQsBiIn9w23RcrJUI1qLkizfWoCD
6fVpCfWEBeKwFpM80rZHqrxHd2E2kooRsZZu02e89Tikr2WDQa0ti1da250T
GLS0210FI8TqDzsOcdIEK/bZmvbQaqbrN9jQvZcAXdBlsuXfzx+ZcDcvg9dg
McAiSuIvfpNxtXX7lGV9Smf2hJQtB93pTDbVixoKTeG7S6x8etg8Sy4Ygvp+
JJMiBW5WVrW//iD2PPtw/dSiTPYvKY2TG9/IE+x6s9SppEUSPu/bZGae6l8c
Bo5rWxZdbVz+kb4BJizXbfY13PHp574M2OxLr/xTKGT2AV8tyvyjFBIgke4a
EtATZMCQFhRSdg3dAYfkMxgY6B5aYnB94u49c3qXVPfSWgeLqt/iTVr8xDFS
Eq/ISTfc4qa6dzu5v+7fySbea9loNTQSUia1gYLZn0E1Xv6qNYFKyvEik4BF
52o4q8Jc5JtIPlgA5HzfkTsHRDydSKRXBStFtXbvmpH19OwKW0Y1PNizuMLD
1Gf8V0pfv6awPw2GEGcpH/HbtIEF7XKF8YcxURyTbTWK4SP3XJ/jtzQRzOWX
04rlMQE072AJnrVDfywzl6pUVB6cf4Tis3v5LWllAu+4peH50P6UY+n3Gfid
a6CCEPEWz4ngsNLMrIdLDU73jhdYlRNNhglf0+A+4VRWQJ3DQc4mm7xLW6fD
fA7diUZ71p+n6QvXTpikZt6YK4t+YBObUiULGq2NtDNZNO1cPOSAB9GwldZx
5z36hjXxAePrAsbFSMfGj6znI/wjLqs34SqGW5wBegKa2nDT7gch2DGxmDte
bH02uj+D5jsDBs7JLZuwdVXdbl9Ngfa2+5zyiQKzy6mkZdWLnfcnfiP4ZHag
JW+CO9csyboCPdzuJotx4Dd0LNypgWu0/2xsplYF8a7/y17HI/6xnpve3vS/
mPxybnWb+CSrSDAAhCOdNA5QhOa2II+XiD+jsgCxFX23+t4hR7i5wDTZJ4JM
2DS1EAWN4hNJtnuPjCwDGbmnd00C7Corq4IRR3lTIvSQ5iaR3PDNKyEkAg2e
fXgRud8ylU0MHQdmtIOKTJQ25MESFsoBZtmY2+/XcuiBO/hCJWtcCTI1/ZAk
nmI1pAJCFAgIEcqwof+ioFGgBe5yu71xRq41pSWjRVBeSJ9NVHo7k/yRpW5+
C4Nl2HAKnfspnGQHUrBZN3RVjvJch3p4ruJ+btczFBYOMconE1ZWOz51MtEk
5+wqcQZXL5PCasoAOa8FjR3w7ETFxXudY7yNp1DBOt1gyir4SLEsvxagBVtN
pIVka0z/Xb7fl6vplthHJxFYizrUrHH5axXtKYQBR1HiaZx5haHmnuH56gNY
UT8Q0x72N1iINHpdJPWmmgI0/A/gBAKHI6CfaLHgjvXP3M7NBLKdJkpHIoWO
2ZJqa/4syMqu3EcIi0H7i/SPm1J6HX9kJiwgthhLceYtcqs2yIJcuxdDcRze
5yfhhdsKK5M3WUr3HWzHMM8dHz5tqeihGTgYlH6lmzHL02rjpJ+d9pFEQaSj
CrLX289Z6TBzIdKVCxyFVNHKWVOiw4FwAIDtAFRfbhZR5ok8UVpxIwLQBtAi
q1AVg+hYPnzS27I1u1FYdT6DSd3YB8vQAGdyaE8+U3viQcIHP1q+bhgbR58D
7R1QEwycpJ/M8qzBY8H/7wFrIS2aWJEQvkNLruwml3KV2W0jgbAaTnHF3O/k
8MYeZRCzNGKj04ZaBLJyqKIhZxKcG+jLMrh+kNnMTkG02egz1i7Q+rLlilbL
OyLtFkYZukbyFiT6ZOdn0YLkX4NEXzw9akLDQ7Xk49WDPuTgt3HtP13oSoQc
ascHp0DZB481mN+pVIyG0SZJxjfUYBwLeg/W67KIFxVl9SivXjSs2CxDLA3n
FPINMCeBoonktZpRjptKonEcGE6pkFvegS6ZUyICRFSZcWpFHwQYScYB6lHx
2KOYPqxI/ecmWZbG64keJscsRrNXg/CfE+/KFvIDD1+Pume+qJqrOWUl5BMN
d2JwAtebcMchPBXeY/+GRoXb5L3nMCsN2Yh81QmA5skSffZIUaXCIs6jhQbb
CbOcK2+AQU+WP6wo3ZF9b0vHlT5PD9W1iH75EKhmN6t02Wy8Vv7QNBL3AeZx
mxNxtTq8S+b1yMq1M6XHOl2PLQCzanqPvdbbN3gX+l5P0TsdBKTATm2rlMJH
4B76SCb2WkZWpBE4Lpkh4rSWdbcxI3OPPrqts5ylj0+plM/pF7zP9cv7cIS3
3P90p1N1FD2RBlsGXY6Saiad5v/+uOzeyzkgf6uSSl2qs1ZOgZEu6UD2tDqC
biIiaqdpqTRrIXp/0elVSOkIKFs2qSlKigQ3WRnwKOW+piju6OPSbI+Z5IIz
RsSYoZrl/GFwcVA0fk8FXJytnW11c7zsAcvSxLuvC1m2eVkMJXhp2m4TauFt
Y9q0EibufCLCUom00/XJi/GYHSSQaT0THtOfpwwJk+FJ3Zw1Aa6YhPYo+O4+
fr7U/E2ZeLWvc0t4JRIEAxcznu6c879OoCioqDUPDdt2FDq1jOQ4ZfIQHTVL
mAegKvWlbNKX1DQ657ZnSD6OrmdOB0/LiX+AxchAyTffn94CZOOLtIcGDoDh
2+llkul4LDJnOmgK/UHmbrQ4VNxamOCmNy9w9yWGsC/wQlp/5rs5rC+llKYy
LnJ6r/hhDZ6RQMJxDY9xfVmtXglXTsAqK8fIZZT02sFcUx8fHA4+LnZlR9Dp
aKc6Sjdgd+J0FwfeiFJQrLuBoRwYqaCbc1m5tkLU0njCC6ZEmoTOm28z5RJa
fTCkRxrjJVaMqlpLCVuh9o66hsss5lA89tEah3uCDalwQIO+JJUT7F8+CY8k
DlBB5z9SKmHYWEt6w6U5DXsj7wytEQ4+idQblJALoIgU/LqAdU+QpOpEadFu
BL/J6tvTGbF8FERtLCRXMbs6+9+/oCLF62WOpq2ob/sVJYAqHQr+uYzsQMU2
rW8S0a3DqTrsg+oFTm3THQF05r7jaOX7PBcuJeinROQn3axlkYkoH9k6LBi4
3IHcaeiDTJIUdI1WmMD/WqU14EXHZMWHr2ItK0CJ16VT9nCl0NsWUtJu454X
jKjx2hupL+hbCrGmnxX6xUALo2AwEwVp1UEeporfuX2pKEhsVXDLrndp0crY
aZO20dSvbrq5QdF+nsEZe38Es57qT8NXiKjwAiGlza/pxDVnzHz4epDYY3OK
JLdgLGEc4MPIZx8Fg6fHdn/xKqaJvW14yNLlad9ou9d3T2iSpBysfeSuWmqZ
kuvtDXSiRYNrRr6bPdDxM9Uo7wwq6A7cKCZ2FY3AUBPjlnWsX/ckwdCdCed/
zZKbAQva8J871c8HpmJs90nRZkAeygFAOpp8xi6LtzMQbeZg+MPVna+NYPYZ
2h2UxNweSskef9C80KVKWbPeUlxjvWWOPD77fCfquqBcuQTcen57pM74MHn8
3/4qgBt+lEEIPBgS7fVfTH+jxcVAavdZ3D/R3qM4MJhJLn8AA2KB5Gwf4RSC
AHj5HAFjy9/KISFcGG0D9cjDAT7jPslQKM2S77DUgw5A1QLpE4XPGQmV0WBg
dccjgX6LF8Bu4206g/kqTrp4yCoqoG3s2T8OlcX2pFfJpZAyK7nHwcbD9hyA
CTvqUDtIQJ0aDtqV/nXL7zYnbjVckLWboa4qoYYLFbAmPUJiVmQDbiVENJWX
VGdqufxJzDfqePBd94/Z1tVgSNsjmgqRCcAnINMLbFEsHPobii0AhjFnlIDI
udDYAqupNvskPd75mth7J86lucGW5IHj9XU6MHjO5H+cQpSXjTx4liy7R564
uBXDAodFp6dhVJg7eGuq8gGOU2ccvy3NHOYMok+xRA1yawC+cxk+J9V6Cn/b
t8qasBjKcQDi+ANOSQhcrpIFDQQPIU776KN5XLij5SjjIJPA0sr0f8n4xzr8
45xaywT3ccZgz5Im9DsVsjMtldTzS3n5FltxJpkoaB3Vr9hmFpxzN/cUuMrb
WMo8Trb4uIT5i3tz6DEAHxCXDZPLqXAlOXGhIt/padeCoAySb0AaANYIWUrl
N9ioX2fONvzhovMTVHTFSrDjG6GFZ1unYqqmV698LjtfZD0K2SBubtyPLei6
L2E+5iPBXV6FjVJhSju87KMuyw1dE1+iLxEECSwNPtM44dLxaGXSwRfksxpn
3JDLjch5tkqxxZfzJqBjqRKLn4p4BywtbXQlNdxlJ33tWKQeGZV3Jjzof8Ow
IHfK1Fi/WVHoVo1fZ7We7L6RyA9MvuhvQ7My2Qf4veQnPKHiSmxpu6D05NMU
TrD5jploWpFg+hnNaDUoVwI/ZZNKNuZwWq2kYeEVCHLTqThuBdsTjq0bVndg
/r9WFXNXwvuDIqN0qae4f0IRpxxtGhDqRu5R9BX07Icsu/S6SaW66F35TYue
/CkVIwvlUup39uwoYrOmdZ997QcVIQkoMtJB95g5SH8Z0YQm5ph9tuDNN7JC
WJSinTU49CyrPc6yuYkEiwbLkXu5OTwYtisxIug8o8Kvu4k3k21F/fxrtVo0
Qw1AzS7+ukIr3Sdgom+W0HMZ5Uakd6EG+K9wKA5pWYBJBlSOc435YPvnMCLb
rfXoH1C83o4PWjlf8v+HtzTKRI0nIBV7HMyVLH/ydePelYgRzY53Zhgg1z/A
Aqmwr5bdynf5zx+woBXPjuBqK/TfpgW8//h2zaAGg2i8JyDCERvezcmh+VSw
JK/QUfKU4NSDcPaGf1qGFdwqjYz6jBy2RBKc/8/MHrLKK035Eef/i3E4+OFd
vGxoSubk+c+nAmwOhVvk0TJj/7//tSwZbuBW7Llp4ST7pb+KL5RlUdALgbip
pnvQa4bRXg8DMzWtznzfVzwCfusnoIr7vW1prKDmXN1T6WmYyFN350iiE467
pISiNhkrQriw7ZnJR0lhE/4trflP0gqVIEWBSWs/JBA9SXGMNy3NxhmghJBo
Q9lqTSK7bqh7GzGyDCFUHDUzbrEsdVusQV4Lxci2N1z+6rB6H5oRDoO7hd9J
E8lk9QyRk96wD4NOFYrnxT6YepgTqcZoBHouw+rEkKz0A0m2Do9ecRPeHT7S
LvHnNqhq1EAaeWnIw5fjk4dE3uhuLS1eUaOK9PLHja2I/P3ZVK0dsxHSeEvG
FI+cQ7jCmotLI0y0Ugt/qxC24h38XrWFqOAqz6uYemJhO7CTjWR/Il4bG+l9
/H6MORjVlW2Kj/UFmHuX5UBLanq2muQgCzovb0FUa8UTRGjnDhM4YZsQrcM9
fL9R6emYiI6uShW3DNkMBei4qALRqxhg4pstbD5sUcJzAxt7TVm28HOhslTx
KIu+UrWELdCMTZyih96IQNwKnehVcz93OyjjL3rdAeI3ZrYb2i2bXfV1+sL9
1JI+/GvjMYcWbB/pw12FQJTnNmjJtKEWy4MxRrY6FHZxpfKV1QLzUk3inIop
fxxW0LmuX1qT4ASrar88W76mBGbR2AnjY1PeOsOAItt/8ofJCTAmhECpwVyu
DK7irFBpuH69Euv7oeNjvasf38T1Sj9TzxI7AY5CJrgcjSBwPYFqs73pktwt
JTJIK1r+2wX3Fh4PR360hW8QUA6BhRBGT98Ja1JYV+ro3NZ4M4XDZ4Jz+5rb
PGUVz/PrtC6w6aqrVJdROpb0NmDb0yDQGhStCrpl03J+EE6Z31V0PoQcxb3Y
HPyo56e5Deep3aODPrLEIQneyz9enX5dZF3jCNYaWSVorhVWigiBxrDaaaq+
Qy8qJuuhfseVXg81cjI3Z2ks405CcPfSgxZBc97ouC/NsVjK/+yKajMLiTnc
Xv7SU1ySx8nuNULIvdbkDlxJ8YYqnr5Wf0OpkWJ14h8/sdynjt+vs+DTzPu0
q1wo4lhqsH94kQBja9mk/76GP9Fa5xer6I4fQqL1vzzf+UA75SFug0qVNAie
7XGb+74AgqjEUYxqolKMNr998//L4NxPTlqnRTmeKPcGlELQ3qoPIgdla24E
ou/QAsQXwLWe6MnHTcXzDe0HLhl2OUknZOrCysCMTme8itrFhRMSysaFAY4D
hh+eGOGMIPp1ABTPTLeP90Cn426FqYDBBQV12uB5Npi2UxoyrQsb96iYvqEI
RCrK3TIm2ioO4TlMoiy8dMNLOHL07fXTaH2CWMUwpHDAOqDMG9h7NUqAsxXo
E2q+XXT0Ui6TL3uGub9g9YExqrwh3kSg9/cIoWveCgcdNc9JZOTIFww4geqB
81lMKWrDWQURLAvqpEfrzQIE2W7EpHl3hWVKPWLBc75XU0L08wc3bBOcIWNy
nSRsArF/Z8cR+tUHMlIki3elmZqQAAfNQeLMx/ZqGmp6EmYwzZTS8D54LMfY
0H+MiDoO3+ERFHcJlL/H7PsMSpT6JHTrjBZF6XasvCzybpqF9qL5t+XC4G4r
Isbx1sQ7R0elP482VsBORNpDwLYJWi+1N1lbOhYvYqRgCL/V8Jth4re2ixsa
Ls5Tla2CN7tkQH/sOoWgMVLU+dn8u6q355EzI2JLkqCfx7ALtI+TBRti+0g3
B55wQLGhRug0jtJyL9zSLkrMS8E61PLmlVoRWyD9GahRWjGKEocvVVcYD6/a
kFtXhtDvnNRNvAi1vx4KlprGlJHlF/ILcIJkbJOrjR4/wzHayDMlRuWNLSFG
XEBacN/FV1x0zMNE79ZLufd6T6II+oGvypDOjzhap/S/n0vcswJuSejwI0Fl
zILCzqXjCkqo+6D6qBVf8cofIo04LN5CAcsaw6+tWdj7AwEDHTjgtSDwwRmb
+KaNGCZYqmipeS0IJOr0qUwu1MqOzu/0NTsl1nfPjR29lh2MZP9xjBW7AFVl
Mtw4wPKXbV8Z/556W19JiufSYclKgHbaaJe0Y885avumgTsphpTbfazS3I9l
3z605vT4bWXUn1e9MrIcS8RtaXNiPN6J+WnLSrOE8lNOQigJaiH2g2aJUkUS
cQAkvDs94Gn8AKDfP1v7grfizlzuKXzdhsvt8Zy82CW8mjA+5cCbL3Br5+OY
v9OoGgQflmSPMBU4d33uWzja8R/MrDZ3wBuSlp8QODA0nTW6G4emcIyGFDR8
KSZ9KzrNFEQukxNszokyaMl02ubwRoJzCHFYbfkZEYjBQ68TzMXg03RE/+5r
15LevLZIyzulrtssE6BGDsYx/kB7JIyFai9smDvYOU89PbGXVUz/jhhDwmTA
x215B6xeMB8RIxRStYaEQtwHPLbZipNdWrWP6RF783yDWDGxKUZ4W/TgSyLA
v/jT/LoIq5gAEpXqMIRUxTqN71ByEL70nnqHevY24fFFMrLei9TbQakvCepg
UFi2d37QIj4CW97SZX+9/Q/4nTxG+oSzECxW+GXHPPVcFS2sKbjRFS01O1kK
SSU4sz0HB8GnfLdqroNfSYaLtNb4LOsPALlYNyHwp4e1k6+auXlECZnJ8zD7
ujWSigPuELbPmudj+EPMnxWU7zZSfOJEqEi6cvZlJNJUp+Vy4CNLMhyfrab6
DBIFbW8Px0PEUQhH1ax9mdWuYgbRZlD0JihTFrLYw5mgcxwQj7RRf/VDGlDL
DZ1fOXcpquSHHlzsB7dGcLvOYHrhw9Va59S5B4yAgmtrtw7rbbZptPad6cTR
j+zB0ZKGEiS4YlagGigWNm1Z7aLVR1ir0uNBdCR6f7s+cXReLLkuV7fmbu1A
hPRCcYvRmAWYxZM8N5DTcKkCe3kOjHtWfAXFgpLhkoQDrrw0Zb1+G181Fg+I
OXj6PLEd6SNJb8rWZs0BbrSMwrjfWZjqETtkNm3WVxA8jDRsEWUuiDHlqYFJ
kRgnzfqCxrVuP7AslkDsLJl2ms6sP9TsWMPt3J1a+XiADlCiqQtxEMt9K7ZP
UlaoRSK7Nh/8zGuCHbWLSeCm1XDL82vDDm1A/BjLltNZkbidBLkdNcPJ2Tev
MdU78FaPH0U1L3kLdLynPDzsHdnGfZr+sLEDxBJDmNkxKosTqzzoZ6gZJITK
LURx3HKYJqpSJ7BD/0F2EgZuYDqCHi4D54cdUj+dg7LV3qYb/X8Ve1/4DEJ1
FSnTMli6Bmvjf149enW7UblgKUlfDT4itqQPJt68bFD7HkTkPXsSVfI9pYUd
/VaXN+/mI4kRGGg+HkHRU7cOn8aWeqwSHhQvbkW/84plLbmbhPoMRGgUhcCt
QiILWeOlHAsFc05fmRvzuXQxfxOIbj+qIpZWa9KWGYQLYHnp1YMjfxVSWXev
XEEV39lIxD4jpNtIL792RTtRcsUvtZsV5Srq8d0CFLXsczM8c6ZSV5+nqVwl
WrTULjwGrDc5Xnm/O2kBi0492PtEMZFHVpOmvEJS3vY6ybmDExi/iGlAhbZY
ccArvzyWEYXu3uCAXOQP3RPeDpiDanCJ/YVb8i8x9VgpOafceeycLwkIZQsu
jNufFlzR3K/JRigEAqcmeV/RAjEVdWpnUjBEpZPIhqgOoNt65gk+v2JC171l
Mii5BLeEsZGS5EivsA/HLYNE+8Qsofvz2J1NUzLbKNG0Qk976vjozQg6fBSV
5jmAsA8vq4Sblx4nBKHJ03OIEvg/kowt3nYzyfdhiQ5AdnkwUdFTUicaRrb/
dg0pWrYfRMZitatsFbrPco7+c7iHP0R5jDRKCbNoLecX/rMPNaBwSVFlY+jv
tUBHKcBz00tyrCZENG1USswQMI7dkB5GCGhac+tylitzf1+Q0L4wMwhbcQ3t
Oez7AAEJFyb4uHqXVLQqLCSlSzHGgiQHGA9QiH4DyGAaWJp8+T31HUZ/n9PW
5P7M9HVlrs8+O49ZSVbkyQGoAg3Wi2UW8Nim05piWyS45chaXEnGjITYnt9X
YmpnhPOIlwUtqz8vABw5UptdDLdEdRMNNRij9xyLUm+nnExOBBhPV8qnw6Ip
oxSXE2Y9hC/z939qL9bXEtqVhoSBPoDCvGDCqzQ72sDow5JcIfHWteeB5njT
NiGqeNUULLb1Vf2DQ6MviOUOwrC7xuUxnQaqNwXbpNZ0zuxdci8rLvddESgR
6gqmsHCOF/e8X34ETKi0MN1n1WaAszQSyhOTolxik873ah3mBTUtDLAxdg+f
RRwUqW0efJbXO3Gx4DU7j25sALQx2ZvJboX88n8TuajYPiKDDtI9LJl2RSWr
tM40B8zj2/X9A0BSIz7BqIDw86Xn9k023JwApGLjPkxKx1QVps34cOt8maDo
C7tC1nJkoOkeJQfJK1BlqKXiGose3slxNwOyUn1sZ7xALIVLnIMVdDtbkxJg
F/xiwF7rjUExEEFqi7XwFZTVKCiW096MOht+DBXDhBtNditGiB4/Z3HJTPvc
4Ye4xXQiRH4VHDvSRMtyzIiTdBV64cGV7Bip3Sa2d5g/BJv1SJ8GBXTSAAus
xBdkAbZ2PC6ZsqZye+WZL2zetDz/6pSz3uvhiux/Ic5ncZbiSjolBsl84Ezj
KDkzzUVAHGpBIqJg5KbhdBoPg+MgcRh2hV7jNlNnBsdqcfl4y+kf9oQkURf1
oCgSxBFXLdZybNvXcqMSzG3GSkF6W/li9Yha5OcahnIXduT54jLeuoVOfHpR
9kE1WTobTBzYnomsUeEaMa+F6pGftoxlr7J/j+ROFz0qdr56HvgUjKfmkk1J
/w2yYD5nWaZ0E5ltYUxzGQZue3H9mhjgBlU1MGM1O+b8idDUHbUh3GXdBGcA
faC2PiMd0IpLNNPvoKNcnd/XFdWF+Paa4MNIXrn5Po+Col1skGNakj26r+6z
Rvi47sL3jb4g8uh3OU7oc8hantz1wyeh4ihGL2Sl2Svbnv0WnMgx0xc7MRnV
dGR2uqFQAhs/08pNcGmLgP5ksE+MfFHY42WJP6QMBj2T6tS+Ag1KofExbaKJ
W3Hx1gjlZpFI9lQKNc/LMNc+wInIm3jzTM0sCoUK33CLAxDj5NOK/lXR9PpP
FnWmuxGCgcf1lVQtvycyxpC2ky81J9peuXhRo9/eDB9NKDqYqxA75dl4BlK7
S0mDSJNhKbNA37YdeVCE3B8jYg7H4+uhtQbYv12/gf6voVowFDMMY6Q1D03G
7sv1qovOZWhF9UtnRuDlBbAsq/ED4dFqWOQhCivNF8TpF8xQgSLK7NvQ92Mp
n4KcJVNJmmy+/b0FTKvJ8/d6XtpdOT97ysuF9i/0NM3nOsiC1yM0KF9ICwUq
hHithFsBNGeCszKWgy097N/17hXDjlTh+queeE1pThERN483Yze5HYzWkBLc
C8X25KDB1fK25zarUgR6M/D8Tdd/lSHmsmlH6EF/LLDnoly5qdMU09tC4XVi
yHzUyN/8jMIAEfeOCfmrzqDJ8GpGjHTaYEeyfaQzBhxGds9RjpzEtOPKgier
Ai5D8WbWUtTKl2VqjqoBaivIbrwACg0cHH2iuVFU67aLxpBQ/yecGi6UFhtZ
OmdAajGkMmnKBBckzLyDdc5EPpjIYKcTBZmYSQnd2lNPVRzgKAayKjWLYq15
DOLGU8Hg+g7fLwV68uRXuD3U1mdKF0qEkTkXkXe6NNWhBbZ+g+3njPDuOWxf
2CVW6dqHntxJiP7XB7NSHuUA3V7FDRcmPebw1SMZSOUVa2SKV3KvGLF6ouEU
o/k9D9kq7mx6PpeMwPMupGm/8/3H1WorBibm6sHPvsI6xuq1pWeZEBcb98AN
3PHu9JW88HEMxy3KFp5rqmpfsEslxDAlpgTdIUqMEV4atneond29PwNulkmb
vBiVHzyTmxtuYASRljE2b1x/isz627KPRsFTVORH+AlhURC8fDNzK2z8wWN3
PRXh9hLx56UwXWOETOCgbhCCaDHwuovkn6K5B6e+l+qqbQWW0EKkUf4PqHOS
IZXF9XjisdUlgHLrCl+uHEnMr2/VKGhQZwNnYDlYekPJfgAiVyICAtIcTYkn
2lUBNsvKC7Q6g3q5creYXXP96sRZNj5TfDvNOq/JrNXLcon6+g3dsI+kKg6n
DiocjDlEpaAqDOJF7ByuH/v8qKnhx410/2DDL+f9xKppZuaVPJsMFkLF8v1X
rUVqZAfPrcUeZHrtnEMMVvRUeUuc68mjXTBMg8j2+V3EBcsa2YB9I1KRPYrl
1UPdIMmu7MEwhCdLxnLqp363gkEJpy+advw+4dghDF+5te24EXyhyWl5UCMM
4YiaARHRgDrou/gRLpXFpJ8UIK2oiGlLBJiOPTf2omP/WTo44UrzBNKtlaVc
Y0XXw3Cbd16+HAuRCuTziZkpqMKcyIn4Q1AYTYAeZzWCC+TO0ovtqINz7HWR
yji/WrVwvUfsdwo41dITBkmft94OuRIkFVSZGrKFcvVeG3TZmGScX0ezf/aq
D6AnKydUnrBtDu9/cvcZ92LxtdPf5BStmzeSLhRdszlmmzSt+buTSesvH2Sf
ouxG7H0A1HhDgsahaGbRvQAE9Mg8bDSvuuv8IDk3BzQEmLm0DIGDG2tDCQdZ
sYSUc151XCKcEZ+KX7fUy1D1te4IsFeHaSZKYeYvThg6G6z6sUZr+26fWMDp
YZ9fn1yz2yrNX/yvexOAL5K2wyhaCHzOKjz8P7oDDes0fGyqSUOS8Y/uQpVU
AoqAoNuqvgkDxQIcLnTbT88mdkHxHKWQsOTbBWD+/sIIQtyXPeD3YgtvxUuK
bj8xpFVbZp7EXAwro/Jc+M7gsm2NzKWtO7oEpHmy1p2R2TIiw0TG+/xd5EGg
NKKSfcphjReGs5lO6VVsKq+ikTT3zvSquFFnWJjHuAvGB6k1L/+WGUCa2Ywa
RZntRmjSTTHYN4/zUow3YBJrNVr+PSwTxWv+Ube/wwsd27F2QMeo4FIL8f6J
s1skqW9KOqg0X7CFneulQkA/1i1nvSuVE665PAdBI4qYw3yCoQw99cTQqryT
0kbQrSMPltxq1S5CQhG/ReCZ+521ASTXLNkwOsHMsHyHggPR+5GSD8qKGlj+
kLPxqLZwUM0WCJTNTq7JddfCCjPDjKRIxU6N2RnPkUDH9orhFUjqc70N/8tN
zlcTc97ukX7nJ5gcyUvtnaM/RYc+C2fCJRazbz3uL9SsHSI4XXmt8g804+E7
6wfHTvT8bFiMOVzmXRkAy01oqj5fIKKFFQnYEzg0CXMAHZ13ajeqAheuFuYX
R5uWTJrQYnJZPVQQQOZK1VxCRbJ9fdK667GEKzRrsgLB98qKlYQJJDwhf1nI
4W9z3hUbpERBvg0NoQgLQppznnhTbWYBD08cUqAX7zvxZvWs9B/gMC5PSyrR
9o8wtuRQN3xgAPzbeDBrRcJR0KJaKzOYY5spbGYWanEDC0rfu/qaH++Jbxxp
Ml5KurwQgBb/ByjeXg01vMb7LM7oyo/kvnp+ibWBt8IZhUtcnMktuic9TTug
GArKG/rQCm/vaAV2FOzMmb9Ser1jN3biaq+hW9RDBlPOu0rtljOWz68NzaQD
13CrWakRiV5mLANM4z5sGM26G+sM0Ew3nqy+y9CMPJRrXPUKNC+EQf0zxHxQ
PjKe2utuGneqCcBbgDinwTPdgmOfR25fzHiJsNfUg9C3gZ5X0f6fuNIQZfve
dD5fgbPPnXGpHP7LRDLdVu21XecUAZ8dwRzMGLqxrBOpm7bdahif/jfVYfzk
9KgQDnZRg2Bnr4Tj05QpYzx5tAFoUoctc32E8ZuyOGG6++hAKBH+qaPvybwy
ZOu000cStZ3fFcVWBsqIt/GvCywm8ApaxskhJkIK3DswHRDM10aF6FqBQNpO
E2d1vzwLvCpK8WtRw26hfXBpwdJKs1YATD95SrwkeWTORl7DFe+wA5WSI+uD
gB4piqT6FLcjtScuPWzGfCV53oDFXtw+AxJwmAE746oqCzsoLxM5DgRjtI4V
GnulYAaER6CkKnPCix3kHXX6rO4a13KZrMRhmzTfKpD1J6PW3g2UNMVwIIbK
lU2ULKW4xY656EBCZy+pT4ip9Spz23/Rv3FDZHeKpewNrb+8S31nHhOLTx/s
e7ZdnBOudgtCFdC4Z//zkpgfB8atpCbao4C54qBzK980aIlmQk9KB16uEHYL
JxNrMNEI0Vrt9xJBJKxptqFdQjBgRRHBQjEEZpHcu4tXvT2go76+WJrF9f4a
b5j4rZutO7CPLuKGeSulMhont5lxWIOrB1nX+MKjXho7MFu4uhXFNCA6AC/v
NNHvFMa4rwUu9KtPSx37nNhDdpIF26RN1i6jcBIpHlyxzBxwqlmmsbU8yD2t
pJbfykOrszFBvn5ZS/ZrHf8TY5TJpDV7w3o5ex9saFux7yXlfhNY908YfLKp
8ZE5IJX9C5AFQHs3rLd/4aWql8YPk0d1EB6lQArn0r/BV82FrF6gdb27Mvf7
GIhYPaBEf4P7uz6RrMkzs7155IfmS71UAk+oXZk7799UX0C1XhecvXXuIRzq
S90ln+8rEpaljJUA8ON7OzTD9LqzBATn5210aKIz52eJqQcAT/mUq8sFEonU
yLh3tdDWIjdawse13mgak9ADDfMekrxQ5FcSlObdeI4KWD2otvypkBRdtOx7
bcRcZ8v7M5wiaOaMxh9h70aejwPAD3+GLp28FeZwz2/noMrR0hIHczHlTEN+
0DFofTHogS/bXeOJDMhvarwUaM2olFRp5pe64Qr7mmcNt1wVB2uGKBdgYJRP
Irv5gHRKUpOy/1FClJqGSU2fLnDgQ/Ok3O5mmJlVb8qmI2dPYfulfMziID9E
lRuDiksxG0B8mxkI2wNAAO3SZgUIKbDa1dYH9X8MWAOrlmKyU0szsqCXX0eQ
3FQH+4gDrG79TemKEnmZQiGvt1uK0tJrvILm9p1IZI+3jEb3cnTBP47EG3Wn
WAdSuyD7ewL92fCbFDBj6uwszgDVpI8TXIJh7s4hBwlpDUQnbjuShRej9+qp
R+XSVYxInQRbCsrk+4toPiyGH2uQeI7BemFN/WqqEFRzgXM+1REbpZXpgkr7
FjISTJEGKtEUq8KU2/iCg7kZQwVaxpEib2m9oCKjbDoK/eHqV20WPpvld118
Z/mapDjGErjIR4lNnuLn5iXWy1/ir9X0bjMvZnmxvEtQ7Ze4K2n23aEfPHb0
+NQa/HRQ8UkKczW5X8Y35sEoNpUUbpRwRCRjjhvRP+Ny+CU3am2LroTRKZ2S
Zie7OoPU2SJ/B2RXR5qOL3ccZUcPwmV48yA+xXyjsuqPlJyq8ffMf1yfw7EG
IPhF+eH/u2632i3E6igpaV7Enin8FWJ/LNVmBQRjWBD2SCuqe52XIdCLPWvt
UJdizrJbOSgzpDoT5gXwMPCBEYiwapcaniCYXf0APKWY3uwGmBhkUkygvoA/
47WLRR0XkNypBiIAb+t04TAYMYDfc9CSklbj1ZjCdp9j4fduTqreN+0VPvBb
4nJgbVGHih0LzQ5TYCs66tnELM5cI9vW3tjET0uX/V/BNUS9VeNVDY+yCkmX
jA4F5T9ETo0CwSrZBv7us0CVdUrx9UMeXvrrfmCVgcZzQ1NCO/XCMhMaj2pF
ZvA4LXnksJF6FmRxUZMpizs8cCpcNcEg8lm8p84bfL3ID6/1DhTkBtKuR1RS
qxZXjKF8QJX0+LunaDxPtwb3xmHE93cSEWTrGzog02TLGV8m/piVTGaHUQR3
BS8kjEBbGtxrIb/n22x0/cm7Onis0JGzVm43C5d052+zASCoFPfh1P0L6/YT
yMsydLO7gGjMaBcpMVA/HpZd8s4m5exIg7XrMZR5x0pnx95Xz14bjSo80OiF
ZQ7p9+gh7I8PR0L4iCPF5UHyf7W3OKX7QA1ywAQKIanelS/TcTxrkfN4A+b7
UI/oQ97YXgGDHueKsuJzy6pAy71S4BBD8BVn+/vWopzCueQ6bvPqcrgyrp6H
qbBltVOSMUood/k/N4mWrFeCJfCToA2jHecrP07PFoB7fTA59br6+fJftojg
2PvmfmzEY61hlCtFPgMIaA9nPzGGMULEq+GG7sVrtESAM171QC17ou3Ig+M9
Y/OlAUffPS6+Ua0t5QoCzNhqvn+mjKhIeL8ZP7YANzGE8L1EZCT/mwt0nUA9
mRthT/Y10O8/d8oOlyUomqU+HX7jiSetegQEG/0M3b6oW3RzcGbPr+2xy/IH
Sorax2cKos2m1AzJ2arYdayphN6s4tXqvdbTpJuqndYVWQUSykkdPmBklZmu
BnFrYNaPjrX4VO8wBza0n99K/8eC6AgwKM1lwxE8qUiU9bJWPWECOS0opiHo
akYkjd9iqjCP3/uHxJd4tH6d54eBNmOHxY6+l8CPErLkoJ6/8YtsPbv0blK1
/HfqQKeig//4SkiqCkepgNnxdjt4q3ryBq0osstvBZbD+++sw/ZKSjUlPozD
N5uz3Fl7ZQ3yxmquSWx0AMbmW7ETV0d2tPC1S2xytCstqHdr80baCygnbFrn
cfF2jYiIrsmaZB7Woi1n/n/0L6r0l4S3j8fza5U2L4dgu0KbNcq7fpo2L0tc
bKuB5h2Ii5Le5rr3PavygcUGT1kLp1VQBIHxJx73+bJyINYP9xO4+wAcWyES
Gt9vH+3aNETfHl2M7pxnCZjTQH0JiP1RMBaCRL3o0JXMmXu+XPOvaXOsqHBQ
8WAc8o5w61Kiv63DzkXNg5VFh8z6LG0kXck8m7dwqOe3eHzqTP6h5d4B0K8m
Ayc0IiuBLR7vM8jnWGmHDFlnM/uRn8fIwQQfyfpEhjCdd1/SJ9PCGzDuN+bb
1eGX2WuNAKASUZFKQjrf2uBTqOL1Tw0y4qqe3+XCkHnuIXsSAB2bOM0lC9LP
gqDzcwMj5bZvYAOedHjT5v9Ds4uW9eqgrzUK664al3ogo8WIjMkuHRyFFq5V
d6Fr7QeVqNjSss1cQhvhBBfBcNNPHSjgrDhpUFNDTpkVZiikE8uTMDsAh/99
vVL/OI3XoKgd3q/g4JbYR6qiWr0GT9NlvzH7RnwhJ8xvJP0/X+PSmr+NVM3a
MpoW/3v39UI96HQMLEtlVdQlw2lHwmbrwtVP6pAu6j+evCP/DQxuPp7St87Z
EH1iMS6Rh5dqZSN6cyn9dLiHYHC2KVLNIGhOG16Des5EbDSxelp4PbPr3zXZ
pPZRysktHFwp3nIOEpzeKHDWiVohQMPgdadqvlhOa2fMUbmSkhOEWisJDbYR
kbbXz35tV1TZjpvqHJhaGii4JEHCBqpbqLaIOObUiiVPXeaCdY4pWU1GKo9b
Im5KfRFcreiQp/OE+b9wUFNg/ndmeQ6/9hp5GNWWRb+ddQdcu8c+/Qcq3Xf3
zeTJc3CJ5p8noR7Rtwzh/7MeFKkakeIFlNvxivdxYvmW2kog8ovAQBnqU4Jm
PizQurTmqsgpAC9vDkPVCLgLYQBX1JF6eQ0ThOLOeEpJ664gJnKVCUOEX8KT
l/SN93RzJekhxeNS4VmDXvwgOe7YTRJh5HcMsULMML2zMz2VhpqwWoKr44S2
pUxCrlbrMpeMVjtgcqjF9XGHtCCpFd9I7EFXag4IlCGY4ySSlqePfc2SWQln
+6LhmbWeI7xRXDem+L3MCJpLa2FECBqG+F+8G0+ct2eRq7gsq8mzsgUD3qOd
I/vVS8LKzFiKvdZM86g0NOxQv1ntxpYtLY7JSKg1hRDkgwzB5xT8AM7Yil9Y
zhPSI8Q8s+NuphnkdCvvRAeyxlo5zIA69MJL1PHLX0TuVgmFk+uNgcAftzoH
nmbQIqJc9G70BP3nUXorqCpQsc4Nb5ZBwMQ8RYWXgNZIOb/vKpwwzK+5NgD9
OTZlrYu0I3tCvQ15iQxZGfeIZVG7err0Gtz/0wx+M3E1F2vNp7fKP07FjYDj
5YVKBSV+esM/d6LL2bG/oeMPWHB0O4zwCaN6YPFTvLCsCd4ZMLu0P+qgM9Ix
ZDC9iuFDig/P+5rIipyNqJQ2udwX20ybgTXjPtNjpXCRNdvMIJbD+Kzyn2gP
qTSZMDwRHvdNqhnEygbW9zPfO4KVdPzOp77SIMHM1EsXBkgDpl/yUPuy013L
23HHE5EXXi4iD25raDu8ACvg6ERDBhk20H/ylvXBWhNWFWMJCRO/67pdaYMj
0+6fHYg5RV7G8LbkGs4bfX2bmU/8C/6OR0l9JwcDWJAq/ub8o1kFMPiF967A
d9AKNuZHm0n8V6ecNbr7lTf7cBWHWtesCa7Z1qs1WusnxqUIvE+X3m/gMYHF
73vViYF9fmQnA+ILP4Y70E3mQWBMLH+kEtx0bj9vDLepOizbN/u3XF+DOgTZ
5557YhVw5t3H5Kdq47yeRXd0Z17TVTdVj+e054PjeYc/frgazGiNj49vo1Mp
Qzk02Ta/cgPJ+epetkl8ycPNz1US6cdhjHERtmXUK7ELXEB3hQNMYxUV+1OR
qHDToqIqw23t9x3lFxvBzTCMSExOlMMRvEzmzAgBExE/4RCHS8gP6g32+uU+
EUCdhi3BG71NVy2pj2ku5D12E9zmxf6st30Kat0ddrkzCEkl3motizpyfcE5
AUL5UKVbCGnAirjHK3h0mIjMPIQCQFbGjYBVh/ses33pqMwUrSg7EYbyZt8j
jr2kPHymUcb3KJCrJmw1hwIh5YstekKOvpV9BvolGT0yns11t/3OwjRdXPEg
8hTPA1ayWeUkM8ZjhYgW7pjdeZEbXgvy9s+MjT0kzYu8VaM+rNG3ihmy7h9e
kq0GJbENWoTLlYnPLHJzLLDYZz9CxofEdNfJGQ/WFMV1R4v//4rWDzljoz+q
ILKN0M3S411PoFlVvWsL+6wmYjcPNZXqfYmMnPJCGK8GxfGEAJs9alWF+7Tf
jbluVdnQtdby+eS/sj1fDJZzieBJkbH3If1XieZf1yrHj1DoSpLmJCStjn0f
H84cDEd8Bx+ILF3a/EsfffdJLDq2aqhdlGd4+Tiko8M51cVnhF5CC0IbCmJF
YxJfPySCwPSuynvscRqMDcdZrbyQVMDiRe6gf/4tM0+4x0A5RFtvk0WiYU8v
Pvyr9EnmT/vAbJRCyqks2r/n4yCPJQw0wVspkIZCDGUHuKBGWfbf++uk0fMU
udqXo1vUPzYF+E8u5+Xr29oWOaETcsEfb/DSlZB0Z4dpHIRMWo7niPsiBsub
ujILvfNm4jxFEmF3SYIzGcbg3LdGC0LMYZ4k+y5SDI20wVcLsQ/E/DOizxaE
3JQqeDdYycN+vDaSNuY4Mq2zlNS7et+/Czeb650615kx8pOwIdnruRh292mu
RHxuLtx879JS4XaLMLFO7SIwNahzdfprOCFSIqDvAHbBCYmDpZod5qSAGelq
ZXe+IHteWxfawWNcMuG5j4xhybp8AbH0ArTBSd5Zh3VcQxF07e/ghJuz4rmQ
p8dkK8Pw9KcI+v3DD+pHhV/D9WnlG+h4zznN8Fcg1me9RDg91OgeCS9KhRPT
FKhpcaFqwPZeS2c12/jb2SNkaLQGIOa1PTJAcIFTLipatKWhCS6yb6rXSi+A
wJoAVRw6qAOj7bZK3p52EwMvofv2Lq0bBAtX5H77i6LSyJSoDUVIlSlSz36c
JAcwJb8Lh3GmzpP3grjSdb0kiCpeDsBKOeF3Ly+mgCByhBep0aYYmpQQF9qa
KfzPbfqdYru2lx/nGhknQvePlw1eDY6NWvh2CjMmSt2JVVmwezqs1ODu+X1a
Jj8g8HeQxstlP65Xfe8GFaNxRpmhmWx+RUO2G7EV9bFZ/aApx8KaaWNsTEci
gzwGYdLKuicb/sp1MmpampZ5giBNghusmGa/v4eDePN2lnKFqbu6l0GvUhi3
x59vnzznU7QjB5Uw3KjpaAZCL9TotRaero02emPHzGPImht+U0ZZR1ZUS50l
N4ujoHbTI2mvtZKXz8q7pKaIjzVKgbK/I45BeQSVYPbd7/eMhfFsBNgQWwI1
suTEeklgbwf5a8Cfx5cKyBw5CWnX/+rfXTG9TeEZ+lBPZ0gjQj6p/r8F14wG
JiV/B6psEQX6jn3U25RKeqilgxtoTsBOeSo72RH7GbqJm5BIM6tW2Tx+hQ6Q
erEd6G2a8iel6nKpd1lMGTiOm3t2DpuFnZlq1eR2VUpNPF3d12V4EX9nYCKf
Hoec2yMfosuu4Ez2zl0h6MwCSFN1oXTgW9cb8HLgl+pNPrzdYhxSTM9gxKL2
e9KAPh8RyybrBGSxSWgEbjW/OXKavwZxmLtJpbcTN/1OORBN1NaFW2M6WB6A
bJ/r6BQBm6qS8cp9/WBQPDFxn5g04//F8MKhXgqpDR054GsVBvKlLVfV6wW/
FJfvzwHd2VhQ2d5pt5HRa9p7P/L5mn20ICgwHBp8+VVV2VR9hwnX7t7GyFtu
iZEvJ7Fr7u4McDsTkqsuvJU1bjVqMXAmqhjJvO4SaSGirASstkNhdH//w8VC
T1HmjOmK/JgtuXz4E3Zh8vkxTxYe+Db2dkoUsSw2A+VHAm1nRcssf+qZVXjL
QbzA08WME4wJchyiJXZ91AUDCQVzoc0PWTk7dNclQHznN3n0jQmg0usvZ6k1
SmIidGu1U0jjCjryf/FJqj/Duz9SeFEJqklt7ZwZBL7abvy9YIC9ArJra4Pg
cgJk0M1fykSIpmEx28aSJSBypuznWeHK5un5DTE8enWJpeTPZZGs52m2Rgrz
fDaGLMnxuEYOLC0lNY4G+amqJID1Glwbxa6TzpxMeVtojft0in0c106i52ln
h63YnNjSxbHl2ossYSc3WCU2Wo/MdqfdNSA31q384Iy2YZ5STxkl1suZ4/lo
xO+i/noWoSmu8kvgJZO2XeEdJBGB0Q28+WJA8C+K5qC0s4vJf+2o1oef+Z7t
O0PTvVuLe9asHURfwhL7WuOyOUuAeBrWlNV/d16x3iSjkDcWhdJ2RMv1vn1c
oOEZLk2bG8j9zN8xkYVNO4USqz0hCYnw0kNPf27sr5UgeGlJOzY7yqgsWpOl
K5OMgQaBRVuviAa9zE1HM/cC63fa2ON9rUMp8yw3OFt7yHJuMFdxL2LkpFwc
P7HOCRf7YPREBjTuPbxGKYabmtDmTO2x4hebinf5Jilh6Ionx2a/dVvHQqdE
2YG9iWapamwRIxPs0i8niCD4FPCHsoZCrm7jCmnWp+RLfaHikJxFb4r6BITO
+3JatXTO1+D4DAtIDyRsBdm14O8xum4MrZnnOu0UYeSnbdrc1QDDdRdxjuII
HQCb7myhNY0fYG0WwdXpgglKcpiSGQUDjWx7bj5EKrk7W+hKXkVubCL7/dwG
DnXgOB4yP3fNvUTkbfdo4b0B63rIqDhTfJ33/siVvW3aje0Z5vcXaS4dS+NG
SSxoFE8+xVhGsGdXVRPMkya7w/CNxKT0eTg5FwN0uPmTH1+n84ZX+rT5W0d4
AYVrqm09Qumt2/UOS6mVIShp6OW4ennywrPSqtIX9wQeZS8F9BLAfD7mfMaN
fZZdPqcyP9ou+I6jE80e6WC/bblOTJ/ytos0Lx3fmrSgBO0849TQ0At5Uo0m
ypzt/EnmU2hkdatNKo58YuBuu6RBhEsKWSsu92WvELTvT/KTvHARrnHl71yi
NcsYezJ1m6uIMWVAPc57RRghhTEs45DIXrauABGRz1lzM8WqjIW5dBVUfBQG
S7fCv/oT9D/5p2FIjfeNUC0XbCsspb+CV2QgirKXis3ybf6bUPiycLwcQXIV
CIEcSsSkuAaK3Iva2ErKd05InYrUWFbZ3RP2OGzbY9Ilgl5O0jAt0nDfqPbm
wS6GKa62wBtIleCJd50VESsJzgBLmw6BJAaS40MgaCI9BpTy1pthhz4Rz31j
UcQpheBL7L6slMeKhKZchRTod+CpWme7tKBhF0B3MSQ6ZV/VNi5au603PvnW
lWZ3ahuzF49QjNDgVZ9bobBOP2oZaJYc3wi8Sh5XldnaYqzedqeAI/tjhyt3
zipRLuUEL0V7oOEOrZNZE/aU6KzXAYtjiJzSsudWcO6EtrNeJcDMro3ICYua
/RXA1dNSWi5FkbozRzZ1oMU4QR2mccBKF2WVtV8g3DY6gjiJrDqDko/IKiFw
WEgfhsWfb26mda1TyYiizUeqDQet3vzYzkh/uOUjcEQkREfFgndgEjdivEYn
v7sgjK2cgtXA78jq7vl8+ngL4d7FJiKC1ULqcoqPWDoP2KNitqDFGjR1+uNz
+PuTvy9P6XqyegItgMbbTMiBPnHUMzBY5yFbZ22ZooKGEp5gery+cbETSfmq
pxfFILopYHILQXRlBM3y//GB5hk6XN9YhBQATXqBwsagfmd5pkhjuP1fvGaL
vf9+qetbJjIV9Bzm3W3jERanosEE8KguEdU2aSG9aPf0r3EINJ65JbigHjBx
1p4mpHkhnC46mDi/P+Jx8jIPVnpXctn0+QGrf/qDBLIP/3AVBGOj1sK5c44W
e6LkKBKAWRM6iqwt8HB+tnVobTBmh1zpJ9gZtjtUBogcMZzP/H+dDMj2qetF
CbkO8BVvQVIPqtD4mMa0xq2mhozUmZSleQT609vyZ8ZiYE/X6kI7EV37/iSR
t5pYPzf7NChVDqYArUtBeralEffRGpL5rJlPpa/NCWTxZqsf1/xJvqz2FiWo
Qo/fOiIQcVK6JxClJxBxapq2J/LDbkRCdc6xVfLvjrHzKZxQf962DzuCP6M9
fu0Y0eRJAhkV41Ak0s7hKK4n679QtCsGMXfiQUFxz8ErIfNfBM4p70dGc6dC
IF9cRn3KB3zdYU/JEle0VXLm1A5HHX64WZB/xNcmPbky27U6fGak22yG9lPi
ac9jQcI6RrOs/QNPFmMUUXIpBuvkoWEJGvS8B9+sD8LgUhOvcWoB2OkC/AOC
dtqbRUozdYq9izd4xFN3Ozrx44zI6B37BiIG3nnocH30k7garLl+R0onnDHk
cz5m4wIwn+1ovG7lfYq8wgX/gYLOgkEPY7AMUpXEn/dS1JI3igGMEuHXdxFV
HIPa6bUiUeAUSnjyhWhb6469kSGcrudgSg+CebYuzc/mq3S9+B9d0c2kRWt9
z7Y47ogJ9O8gPZTxU2XkW1WDRZVPHMV0D2Ea3ssSNTL5F0OAZhLUkdXGItPg
wSweHqH4B/CuH9bct3GFMVcMBeiGKOIoQYi+TMDmzzIWTL2HthlM2Ibg/eu9
XBT/1peL8Fo8GIgpY6Gjd5+1ANTO08AqcZHzOa34Mu5eZDTE+PgEylFtK3xw
n7rZHzqqwt0bhzS2i7SJGHHMye8s2WJXBg2NtBI1NJs8o8thquxTzQ+UOTmn
fdloggMKqljWQOu2tac8ZTE4JOKON91EKxPvOYKGR7p5sVDOQwSg51QbDH0P
cQSP+N36mZP7VMpJoHLeuDHCzuF9QQr4yzD0sT8fNyIC591EQKsvOhgGcj9B
AJnZSSv6lLjTx5XGYP0TGFXNlIWBo91uXGyCTiWf+QW06jmqu3MyiNtkHh5e
CApbGg7XApP6uOgRu6YAvCO5FdTjDqBCJgS/tGywMyATsARazks4mpPeYa1U
enhm3penB/TiuFqmqTw9kwqEnEx1lrfbEfEeL6N6uplZYa/Q6KzzV0nIgGlv
sheXd6K9YGhzjV+A22RPDUjBuN/533bOXBiFYsmIV6declDgP3ApBkxSqNxj
rbCMAj7JQTwKryHtt44KVh1Zy3PIXmdWwe6fB14MChPmfo9vOxd0pI/ZPyiF
YV27lJndIB+L7WuRYaJcNS0M3fss9NapBVcLEvOXd6nEVh+2DcOE5ONz7Efs
fxRbPx3R9sLfU/12KMzDoHwaMftIIygjY/pxzsS1+BghroYqoMLUpveOR9kM
/XNZiZP6BSxzBKyNPk9jZ/mAOOKeDYm9P+vKBUHtxZLKFgU3aY7aanRwu/9v
gHaCas4a0PB6mfm3DR4/hFY+POuutqrNXq513gy/9Bkcpj+2NjBry2zD6ZMf
6AcpwNpbgUlqwqp5+fcIV4QYo+8+NV+PLa3UhfLvjrFsoOW4RJTNc5qTWV+i
ycQ+cSftzt7n8bZYHmNyUBnSJ3NsNOox6NyynHh8Wj944nkfFgipjWygE0kW
5D6SqXg48gCVLegG5cqd14sO+nAfLCiIOTM1O6RNs/tdcSObJuVDvJd2eM/v
njYALHLc7rJcRwZl6NDm9xI4sgsnfI3Gyh9eOQHhvRe0Z5XB6hqwtbLQDoGa
mz5Go9QSB8k0EP73Z4wxem3m8cu3zzFp7Lj5tEFsY/IlbY3EOHQMVnnGFCOA
iQw0Xod4GEB2s+dG7+jkgNtm9kVYT4Z23Gh3ILIbdppfbS5yHWek5epJ18F6
XfPYZPGFt/CyW8i3ijd4mKPd/QGWvIILiSWCsz83tnbutE2fZMDV4ym8jvc5
POpb9fqHPa/69PBHgxYvbs5tQal4R9Vi58x9U2mlDMU1yIuHKWglcPQrVhzD
3ggxFnjFENkBZMxiYITf8J7jwp7+AdLk0H61p0ASzEy386czPCJh1UQdwnbD
7Vvu16nkMPcv/cZ371cVeMEYSnpQsjJ35EDYSkoW4ITNhwd7rkcKMqflPwQD
bpcSOtApVf0j+WBjMQxQbo1llWOtDLuhjitMvya03pKJEVmMazIupvh4XA2V
/7ABae1+kmtRUL0LDLqJi6gdPH4/T6U2K9Nqr9i/rZvOGXEW79VHX97KAjdp
Gvcw501D7peVqn443s40dykfIhOKtFB+YnnbJkOLZFNaejIQWnrxv2RgK8/h
Fdrd5j1/BGD2+Ayt3U15qTpXlQ1IGBSc3EdBvuq4jT0kD7VI2MMvUSmusu3C
OXuVIKZiZpF4X2LNhnAKpDm6XwRC4201m6r0RHAfQGuTA5d6J+xrrf1ROAii
fzloNI096jqR1Y/ti8xxY4Z5KEfDY6bVx/BVnqNCLWuc9OVLBg1AwAyeJe+E
8aqX8eWIlIx2j3Ifl62Dm31QIvVNcFbcxA8dzLj0XRKHP2Kpk8ua4L7WxYZ4
mGneTxz+gdTefhGRleDlVQiEIFmb1t+UOLD8+KlpTlYWpzGD4rIGv6OML6oW
oPUAktZIkA2JYgVCTun+OOFEg40q0GWV6DmEpaAY/4ofG7aX34WW7MG75uBS
K4xrHOqJAUgNBnH3ln/Xe/1xHDN2i3LEcDoGSR0milWl36Y2uf+sD6FrKCcC
gdeKW1dOud7zzbtqv7Db1Q45d3VhQhVswY2mhsuuj0fM7Eejhid4a3mGPqBP
icnSV5ErCdAaA7PQ4zLcz9OuOvdU7P3ro5njL7dz0Kqu3r7JWS9mI2nAsXgk
KBNlrOG76eSpEG9S8cUdSNB6OOM4gbo8bnZxTIKxct7ezkfQQ/p5IKNetLSJ
MeKunyjlb56/l0WtriBIhrh1REQKzuWoFgGJUyQH9+b/cRjRMJ9IYdQthkKV
22dZkWC0pnBIQOGE7L0qRu+Jy76sKFU236Bli3Q3l2ebKkp42PhTvDFGxHIc
IqYxIpb7V/NO1orbdhMsmz5B+sr77uUNQcum7pi8Zu+k6QA+P6QceZeOVgqx
1TiusGo42fr/Y91/fRxhrG3VbBp64AP/KoOsVVanvfVA9Fhn0po2UDkWYwZv
MwDH/EKKVSbD3isn5QqGXJtPiS024U3HJdXbhxhN4cr7cnU1CiVIuNQU4ARe
Y0mHXIDNAiVaP/rQiuKASnt9OW51viSIIVw3qT2X2R6X4RZLd80hs5sp2NFm
ljaYMzFNMgR8vpGp3bEviftWCLcjw1vo3K1GCMpRHR1X5RSEAitWtv8ur6Ey
8jLB+zPqtK2S2fOeA57cHTonaw0SIOfj/fT6IQ5LRla4zoQfjgW9rBjTfizF
MhxTYbzrwSMk783QdhExnN5oTe5ln2Eln3GuWjwZnYTC3/hJQot19DT/t57G
CGE6Ddh/Sjm0hyVaIt6yMzXn5mQkImk+H8v5trA+RappPWpAr1OL/2RayWYM
M66CqNhiOv5HR3lwLvYZmNCTCIFYNUGG9v4EqbQaix/pAGE8U5292OpWGtPg
sMC08hVqeKbYImxgKIrKXYBUpWdlLBSp2NvLEZPygZIlUvRhMewm7Suqgmqg
bWO3yGyPTAHFoeA1wqlgHR6WcQwuGlhVGlWMD80zmhbwc3Hstloh2JKTvB5Q
GZOs6vsWgFShu85txA+vLwQy7uVNHuybvQ7SvIxILEiW8M5PS8wC39L0d8NO
ItCLMBVMZf+v1O7fkldC0Z+1A5bUI+P3qyzUiHeFJ04v1HZZrA5npd/01FI1
DV93zqYsL61AX0D59ONk93QnTpG4lPPH4gqDtAqIvPuzJg615aQIiLI4NOjB
txi5KEK6fwYOEiNDxJZwnAraB/c2Y02LvUfHVAwBXpcIkSv36WVuVqa5jc35
emCbay6Lxom54Krx4eJzHMHHmobEvAVE2t1XuXBNJBWO5S9m+KXQU/PV3xrB
Si4YRVsT0Wm6ifZeDzw5GtFVOg5L0GHFGfKW6TjMaWgPlyDS1aw1aZ/VfrNv
k0e34B9r9NFT+tiQ+9aZuI/JTaf/1ovTavsjKrMk4b+oylYtznyF+vOHtz3P
hkRVQ9VPpwILu+KGxnY4oQtryD4A5WDJ/DmEnBHwY1KxOSRGCGfGucT4nmM0
Ymf2gx7CZdrYfiZCl+Sdx/yfJ0EQ/fG3dKAvpxzl0ANhrz4Q1pkYzQZ/tGJJ
SqQdBjNV82M5GNvRgvBmdR57FCP7+EV+FzGbtkGDZ3kP6q3ryNnXpdFYQSCw
gjOBht51/cFc8lqMCCWUm7WtOHVDmMrnJI7MwEN4gMiqqD9n9F4XFK0eojmO
kfOjUETeRPWl73wafxShrrEOgNyDDZMjdTCFBF4uemj/QBxBGsWSdpI9L7sF
9QuZE3m09xwSF4apgwXrx2Ncn9d3tX8O/8nx216OFu4dbrcaO2XApHYsPyIC
0zeDEMDijrI1EX8rHTJL19SgDjvtejourHyo6m14tgiJbDbyXoJiCxV+x6MR
snN9C4rZodZu2M9Nbmmg+dhkFqNB0TE3bjGGxg3WSZWfQpnvKviSl4d6U3qB
IAF+Z5QkoxFMP5zBl89QEYRJbLVicZsEllg9KU5knq088uDIOzErWt49q8uj
wwxtPNPDU40G6cBLCEC5VeXyYku3B3aiuO8N77CQWDMig0Vol901hnKMOzFQ
IIrp/HiBAJ8d+3PY8feOioIsKrq6qvu0jw6CKxRWlOrVC7QPphw3lYytWV8L
ekB89gZReMFPNKd6t9BLa6waFo157orOYAdIkd6UURrkmHB8Cxmp7vs3bPC/
RhOOKHqhF66VE4zvVbg9LutEkLP4EMnrRJcuzMnP3fQZrgLp57pUjTc8twIK
SAgK8lSwAI6sy+Ql2+W8Y5/60JsAibiYGjLvGIENc0eiis2Lggg0s9VGn4+L
Vs/gOM2kXWTGbfZBbGQ8Z967JExNNipdKWSb5uR7iGUiLZJzlDtv2MKOm7U4
/QV+8eqbKi/P+Q3PD/L8tgDYvVprFxHOjLUSHT+CUKk8PU87nOFbuzWc2wvc
YafKL4J9kCoQUBXrXrLm+FiF2liv79UaZQdK9IMG08j7WIFT7w87s+sHPAow
2wYj7msGF2egXLBgbUaC9kqMYBmQTTQ2KTyY4oTJvz1hKyNPvTTRAWAB3t5X
nPaPYjEgPcmAXG1ZdBs7bjosYTAFW5jx/Z908hCMejONowgmwgYFP+YvBUEQ
iObBu353dNNtTlJn51nJvsSYrewyRfnAy/dRwuo0b/IXtWcEswAuv4bLy67A
W4nlIs8P+J+9BblkUHYwZu8dv7WqySdkGTa70eEvDlmLfzFZDKh50hEHnutR
LuMq+8g98kyIM+9+EUaGIP77sYx1ExblPgj9Dm5Bd8q7lyY/fbbNSjj2pZOi
sSzmXk9DIcOAhEQqATIojX41n1+8IMhlZzS+AJ7GuKe3UbZRjddFIq364s/h
NvtnUniewyA7eu3sTOwi3FEi/WmFan/Ib/Vjn5TAKMTJG2OD5Tv/cu5ZjBAW
mDrMBHWKdtxnYghkABW1jXnt+5iY6BORSijHFIBixdfmtvYnCdfVqnh9oqyc
BIXlL52Ln8GSlV/la4voWQgkVzQS9QNEpTKcxMdNZAGWmj1bZ10Kj5OIaSmC
7xaxjgFeQdjSS/8IcjJLTAieZ3B8BIVhVKCc7Bod0fs3dWFjyewIb8nviJPf
yeaMIjGcuJiJk/9+abL+DeCAuumbMs5YDjEXTKt/8Yj3AwQFORqRq+RBrNAn
ZQkgmaQYIFLlSXs3NbwmXnCv8ix0WciK2yeZXfxsn9x/IXKNW+IpU9UDWIuu
Z0AjX54FoMqB1/pTmIygcxd94U/AMfo5vQqMtpmWroQnlFWms/Qpj0OLpi9Q
B7XiIhvYyIfnY1BMTd2TnnWpt9+gVhAM+dqUtphpXeBhPsfSsBV6uBtOmhsq
+tF9xj4w/DlTjXrVlrGTx8rOKtCB7pg22DgF7uK3nsEq1muE5N1rNwpfGIjk
TGd0bPYFN8/OTfiUX4TiqISpJmvGBQGb9h9ynn2i3ZTG6LPB/gGvTcvAUZ4k
BsfDnnyief0De+zE4ZgVpLRd7cgflxhdRN35P4ykkSAzbGF6PzOVGSXkrB+R
woJnNEvKwzZ6PlW97SgLkQc+g5OFEwWoncR2nm5sSDvhoy+NjEFekYzvj2yl
ctYrSQ/oBpRw8ZZzjPDWReN1FzpKY1otFMl+UgVhVjMpVKDItGjdljc1y3Nw
JECu1IPBO0tbA5ym4Jp4aW/WBCfyjPxyJcdauld/aknefc3N4UUpoUwxKnPn
OhqlD6EeCV2lZA1tHRPvEL2A7yGOlN51cQtSs9GyqjQwxGgsugip/WuOZY/C
ZWtMFit2BQISP1PIRfkHJhfBqxgl9tPgajhhwjiuX7AM6K7SfwHRFV9mYYl2
ALX/aVYvZkdTxhCSq0hpUuhKXpVDGjRzdZhkm9Y9Ma2KXhoGT8rt3iQEWcBH
5yaOhvCpl5NXxrpKmjJOLlxZOSauvC3ma07yJEE/CqP9H/C76EkSmq0Kg3PO
gfb44eJIOyo0HxpDGxI+qp1BRTFpYFFR8UJbFrb2uXMi3QuowAdky2aNulJ6
hFqBM7SLgldcE6n48ndq6HR2thsrZGMNLd90EUIdnD9QiCJi3W4ofzkO+1Mt
5yjrIKCgIw+zAixCH/YO5RxKVvFVzCMMPxDFparipw7knaA4DoyaukmW9YZ0
6An1SHlPVG9d7g+3wxeCs/Ilc6NYcYHXgwZvxnFGBnYpWPFxYrKSTPnaWT3d
avoRYxdLd9UZdIKOa2KWDhMdFE66WTmFjFQLyxByIo95nQ+qDEoh5ARoWP3v
Ds/Uu39WeDFzNk9axiOW55mloitBqF4Xxis5WwINnk4+VUicVyoESD1dCZRd
5itWp2QMEMz4p7cvL129G3j6+4DqrxlhTZYknA+esmuDxfqyp7NOIjpnyBFn
rTD+FB2qK1FsgzqXht9FU4Zp+qNgXB64uj+bFsxU8BYbzjqDrqN9vf23CFpC
ngd/YqtU5MR8qYAgCAf0up4PvP1XPdh7z+bV9Ud/uxN/NDs93C+YJtQqk9wE
quZWwh0COWSOdL7yJkPuI3edOLREiif+7BoowCmw1Etoi3bS/qGBPUBExDxh
nlLQOqDfrTiBLPkW3optIvs9A5gmjunw+cDb8sZRmEmoH2a7/STCoxC0qBBJ
GAaqL/PNNXm2YlwFevXc/XQtDHXr0C3UPpBa8sa4qxpYu21/2mA8i2F2QBjd
VQA86ERescT1XYJ3xjykwJE6AlxnJZvnXXc3L3SUIRbP6bAO5CMrT1GPKLov
jcGY6FGd7Y/llC2SXFncmqiSNXsebfPIqMD36UUPA8oYXf/A6YPTSMzRQRD5
tkpD/I/1/WW1trSNKjhPCdqKQ2AqwVLE7hTftrAqBYuWWf4lP65DIsJe1BA3
uWAvrEgW8Oprw50bdQ/uxp10/6NM9RWxLDqil0bFvt+6junDSJuQzVL/8Gq5
mqJ3m+EAYiCgYz4agUJwSPrr36OFbMbHycmwwxqAiz+LviGvyESRPbYCgSK4
mCF7Am5975VRE5n9PiVItl4oBigR1jrlAnKAbLRDxbrMLxu2wBHK7/m2O/xh
RVgaxU+atBTJ/sVRlcDPGrV7+bAOzUpd47SOOcLDlZntJ17+ddmQhbcbCnYX
gmRXSuLwNV2UHYkzSe47SLNOkLnHb+sHq270YSnsdYN+HOcx3ySqszpjJe4w
qPDxHTAq+4wPtrTDwGCZb9zfYNbj3r0S5Dfmx77thgUZ6aKr+gVHXxNxTPrZ
df/bqXqHL9VpnwJylWVivBc/JXpPnYXqBwDj8Omx+cYdj2AsrAVv0CebIPjL
LRTwWcrsRiBlr3gdCsgvX+uGZ+axZ3oSCR/byv8lpdE7dw3NqsMjbA5cUCF0
kkpDErVx44XubpJL442/TUcSQZQKB3mCtm7B6VN/dBnVn0g9mVBsbYc9ycew
VIaE9cZU6L5brlvfHXjtfXeWJZ0iea7kZamBSnVfVgsYWrjMniklyizxviX9
wtQYceDpznDWy7750k3pWfbzV/p+U6UiazTREzeT6c6w3R08GGlXATexIn8U
D/8Qmu+fXy8aQWv87dxOcvmhM72LI6YrpfOEoHgYglxShoIU9HKFxrQSdfPi
wBvP9P1j8e9TJkUDj1wDd7bH9bzLxv/O0wLm0k2EQRnKrAK/VvsFiXVHqLCf
hx7DILJqh3OruAMk2xLP6vRv4y0HskKJsVCGVcMi0doiUTuZ5AyXFo21GJWD
9HmGUwkGDJKABX6tBuceOiHv2/JTl1kRMR+Y13ESNZkhgnueP7S1wfscH7aW
5GyIU1m2Zedpbr1dtOmwX638l4RmpMOG3M2VioS+URn5jwPBngaucswyteot
NblhuJBjxQ6FIESrLZQtsxLa5gihpeTBJomdpOjfvgAhJXPldnnwbb1qcdeY
rv/hK8h6jopiSUcIwXCwkKPYdLyGZICKUoScraS1Q0wcUSmuDjdsc4Wq1ffu
E/j8OZ9VkRaTerdDfpeu/6+XdcCBjzpT6W4nzaeMrE46AsWjg8Pb/u8qyQkl
S6VK8z8z47eauTywS81tfSycis/LTh1jVF2k2FHIsUDG/5I0stCeED5prQ+2
HF5iTG3/spw2Y+kTaSdtS3ndntQSrIJ42XtclM1XbGHhIDIiD7pJn3Zk3GAx
Wi8w6leXKmCK6H+QfKZquJD6LecSYlSQ14w74mLG2nAEDZKWmrx4A0ZLU6re
Bj8q0ZoRKrb4777Ogq7bajza7kXjgZbXc0E+PgD68pylxdLcy67lLGJw5CdO
EK3BdtljYnX7xg6VRu/HT/h15V6RwPWSZQuiHUahg4zgnuY593PMhh6kOb9x
dhxBucz95yxgMT4kp/NLL5+V/7JpEa4IQaZ6wcKBRZlN/WMH8efdOX3DK0eB
ZU3c8alQjomwyukepAK68rGSFjWAHZwYxgRjEgRCKrxlNWWSARQxCGVUSLot
Myce3lcBUlPnhudiginZ/bRXgn45VPStvetU5sY1PgOQj63KJI2TewK886gC
PF9UdY65YHNhpoy0wzUp9khcVRCDn/PYJv7WYHjASNHX5oxH+b/L8pdnEBDl
yVb9/8/iRkcHi56+PaqNTEn0mRQv6dYYjxyJv8YsM5wrPRUYyaYbhtocBE4y
WqGf50KpycD2G70E2t1QLMjnpsrcZMCYA2KV1fYCK0bMCOxExm2/YKPuPXsG
2KDgmGj7x0rq8ecYsVVebZXgVwHl75xHP2bqauGbDF3J0yP1hWwFoDc0/iSM
RNHUSoIDZlbLQem1cJulOHSCrUvg1d8/gzr0a5bNKDObcBfB7mSX8AoDhl7v
c2nIdc+TtitviAtag/WYtQkQZwxv1fTyw+9viaPf8/uC2U1OqfTNG14dO5Lb
C9EfktBA3ngyX4pURq3Z+Km4eq9dFBIemYGys1VXCCMli3qnuPQ0EAUML/cH
sxqvX/UksD9ycCOriUKt5xP2tGemTANFAIYY5ZQ0ahJTADXiVGmejwq53/sA
gaGxE6lPzcdxnFt3RGlCdrKPFqVSCpLiHs80QLek0zWuv1rYEKzE8ci9cB0M
gFwC/tgP7rmKdtxnlIb/Q20v/WaE8o5XsX3Lk03CXNb1Iq62MI3Q8vdp26nE
T8GDIzhr9ApeKs9g0msMPJHLmV9HeXJvr2woYD6brqylT+lTHLvj3EgTfe8q
6wvQTgW4YLDr5hrHK+vRV8e+qkUPVR2mh7QFfMjkAMVAx9hwWnQfSuTlrz5u
tpPkHb/8ZtqdrXT9sOBqp/UXmJu7RxGJhNHlhJfTg3GOET/keCaM42fHQO7t
tQoQ3estLGE+sj2kmaq345QxX+KITm0YyY53l1vO5SMrLcyB+awg1BJfs18v
lLf+FdoBxTzx6iDcVaO05fxLDkWj6GZBKG3jQs1MjK3nJDdMxFoyzOGdmrqt
fP/yj16cj4rJcPQ1Aj4xzm/uzgUvzKOXW2nzoJPghJP4JXn8D8tggKQAo1/t
LzeoQRL69pR83xksAH3SGqi+niS9MdpItHKvXI3tTSpNJpl3Aa2fgMmHg0Po
OD/0hElZjG3PmCpwrXav10ppAKpZ1TPmTbwm+XwR3mE0fnnAg23M9JML6bae
2O+diRCftprTI4NfR+wHKQJA1gEyej9aA6Xeq3tNowpQyY5eizg6TQe8iv7C
bHy5/fhSwjm/od6RTFw+5a7FhADk+uqhmDzTpsGwlTSysVjKCU88UzVjJRyp
/K6ukNDG/8TDOgQZnfOQ4he8ilM6xpxVDLkLD8K7f10/Xgov6aAwnYuIpAxj
szVM4CfMPVkIeSFOpIuuLVyTRZ1sXsV2tDzmj6Vap18FdMFNnBEHhIOlYkf+
pX9m1ESz/ooTELIGXMmeoPXp9SxnKpuznClYCa/657B7u8RN3imgzNmAbEUn
jJp9ZrDNzmEFgkU+UK9vm2w/D+guaZOuBKheUHhLjGlkhiXK0dtizE8Fkt5U
WXGU64YMEnKIhKteskSIX72YcRV60Dfd2RTvIjInP9djXdswS/J6C2WNBHgT
tgCXuMzokU13gctNxqSeGNTrmXEjPb7uVuM+XN9jjfpjynkr/V7Eo3vhgTOR
HZfh8kSvS695cObhnWf/8Q9XfWAHUjDHcKstWqsX8Awo6lISENBzx7RRPR7Y
zvkULGVoAcVNExrCQcweS8GDvCCFFR+XYyJEQL+64ogwdcmvS/Xp8dbqusRC
UhsUbJC7dTeYA8Cut8uqVPfptuOkbjqs1E8j+KQgaixCjDz58T3zLRbAOvkL
CuC0XKBgngi/evEmblWQxsHDc0X9+reWPvGY8+Q9FvvrVwGEM7dSOsW/P43f
q1GDZcqLI81vKyFMDBa94a3xazbd+ugROderdyZoWbW+Y1dRPNjVyIMvV76z
uXwQak4F68T1spqic5UYI1YHEf6Wk1dKE2oE9YkAxGkHTwnrwD6BfzHgJwHs
7h9td3uxKOyys9KPgMC5lIQFSX0CBlEL2FW7RKNXM+uxbvJrNBUVwKtrB/yl
bACdB/q4IDUMdN+qtSLlvZOpISKdxM20SM8whGfunQn821BdT7fLZXsAhCkt
nZCjh/9MeBLJN472jStF4eLi91Lvur+LkLeIRwiEpPNDz/c5rQoBMsrViH+a
Gn7V11zODvYcICjcp+iWvHOnLIPky7iZ66DWDxuosT5c+C1PJfEQI61f/Eem
X1sc+atZkxwpE9EVcDzVXxRszxfBUK0wXFs0QNankU0L+dfkOZjSwhoPFgiK
FOXDQ3gUQjQbFHhCgLi8V1NrCxSdXVK09Y9KXD35aLRCh3RmJ/45SUKsVVp4
P5HN3K6+H92dDqsHBN7d3dpGZYxvp8Wlac2W19Vupp7DOvXdvBYywHWkc9Z6
r94KHiat9Bu1GcJSCUyBP6yWi/s+b6Fyz1scq3cKyCvybIArENLgsXn1V4A9
EqIW77ff4IEPXxV1Zer9MDgh24rkJiVlzXThqZxnoAvhMinBxKbzlsXiLZUB
odcAl61cHZskwmg8NKPyiA2A+iVSEDaIWQOq6vCLCf9SLIDyj7gwYVxC7FyC
7cFaRfL1hFYnByqHGD6pShFnqyGtjKBY6MerKE7OD1S3rklblwGHOTGSkkHO
nOgA4KFGzW2ogWqj1nCpN0MQulR11qMQiVGNmCRLimQEdL+tVQQuFW9FmM55
WjFUQrtr4Jr8BWfQODA1Zqm7+IaiO6ynNX4WpCU2urXS/Zbctg33Yt9s5ftp
r49R7YEjM2I0jKZERCW/D7OJyuGsEU6qH0RMUZZea3BJmt7rGBKtfgUrmqjy
BmxrpxXGBgoj4gVcCY5Kj0iDItbx2kSDUfiPKF4dvrgOMZRnGkPa4HVHXtuN
4eApdu9NdytjY+TwlLkDdZf9+Ktj1Ndm5G0toeNXG5QYbxITC7HLhvJIZxEL
5zeCTacMK/etPh0W5PU0glQm9SDmsBfsl6R6bcNxNFcz/YQKTqqJcfSsvzK0
gxKcEQWcfaTeD0I128R1zs18IK9r9LCwaAZPL6190x9HUuwHmT5DHhDLtj6t
MkGrpElfyw+CtWUSnqtUhzC1tnrw3v3TeeL+MBlL/cg7XIEungj2YHVXwGBF
lVy8AJdU4RIAAtn08Teitb5nqx92xQnjquTQsxySXWYh6h0EXOCfFQZHrNA2
2h+hrrIqvQ2Fokv8f8Ee0HD0Qq0Dz4VQ3V/59eD3/bM5o7OkE1RxvSe819OC
N0Je0vKka5zQKrB6HN+0L//UiNp86rQqqUkaJfRUahIUurKCDlPvBw0kvjIE
i1584QiuTeT9WPx45YIk7nqernM2HI3seuO+x6UDrnhHy9qAjFZsDW5ZubmQ
yh7dL6RPLHy2TsuidVBYko8UgE7CpsaqO4ZzZcDTTZIibkLRXsOyxj+42bnO
9PEeKP9zClNwULAy+62RfcXxanBwvvlLKWIdQ4V6FBYBOIH0QTOGvC9jgVv/
zA0dXUGywIcvBoSDYEuegoOV3Gr8iGwAdaGQw2iFPTh9zz7ao4NlvYYsVJ6a
Ktiw226gunuOBB/LMYkTxU007+FfNUyHnPM3roB5LfBCHzwLSZ+3e+hH17hU
KULmodW2PjJqf+LBGioxqP45me66Si1MZkerMVG+RVfV9SCwy5REklACksup
ythRWC9oTmJooRGkgxGNHuQvLEFy2DQxd+iIO6jis6tLXITDOEloPUHPE19a
2O14lWX8GfGtUMR4BKp28l+LhR0L2PT+AhtodrSVMqIbgQDLN3ukeWUUHdjt
TIrucTYEyIyEJwqUOvriT1LwtCzXth2h3PgEOfmFVRRTw47MV9TI0Em6WYVa
qn2/MlPb+edIYynO9moEU1x7gekNvTankYFo5n8WoB+4c3FfMACxuIwPfwYq
GD08NParIUOVPMmhfsrWS3dfIZ/Ck1ncOpEGBPU0FqErSQS86tFlF1BCMXlV
DY0GSkJpjq95IvaB9ScYJlzOpIMD2VZu7VcMH9m/CtpK39jSYABr6KbmBEDE
jDuDf0NyaacXOWwNc+UZWuTAtIv/aSGAjUlWz5GIjjcmSgwULZwyVYTmMwJV
zj3M1uH6HUfwPMlALC3aNPigz5QqC6uYCbJAB/VIvR4zp6J5Fn02zMzHTcn5
iR0UD8e8z5XxlDvIKIjOJQtO4b8jzcVkNjFcOI71dSfpBTOYwVVCr4M3UO9K
T+VEJcIQxv/laJRg6LeLKWyOdODLp8pE5trZZQxdXdwh2kFV/QqWwgcwv/CP
Cv9MoVuiJ6K1u0a11YLAe+hDMqlSUfce70t9/8SMiHc0gCRFkn0izCsWh85q
8C/nzRevU1JZOUWGkQnCi0cWQ7zM+xK2cIZuY4bjaP3s+hbYpJE3G098As87
bY7klHgPDewUWcnU8AEx16XX2Mbv5bT+qNvntzPMeh/APHfS7YsBoP2485EC
2hILV/S18g8D++rpoOsE1bUmcP1H9TYP50wQNHBBiJ+XzwxvTdjYW89RmDae
TNDV54IN1Uq4QjgAqDW8OGQ/jce6GmdvqySa8Lcuue23Eg0poA0pb2HZYy4g
MBwbTpNGFfRAgJ0rVHMIHxeHdSuXeW0oeeMqFVJLP8MUQ9jdzCGKug9MTmYa
bw9gjEp1+eZA8/MlpRvXYRgq9cwQEZgEtBXTvO5ROvkdW3ThkUNaUNO4N/Kl
4wiiOybPWVFLWN5hX8l6A+WiRMzSqdb20Jss+16W3JqPi1V48gcuDi3ftboU
UHEkN3uyavy3zGCGeACfq1Vxhy1J2+7UJhuUDpjtArrv/4yGocXrq3u7ot5B
j9gkh0zFV2sHbGioeWz7Iww/YD18e5aBZDPMnqLRVgauDKy8LIO8nPI33V7o
n0+S+/nR9yPZcWMUt4HFqQRmxDkIxcxWAevwYV6k/nhTup4aBdzoifkBR7iy
k7s9xvD+MaRlK8lf5ZcrwyATLrkVi8yNo0kNRerJDtCZWa94SMpJKu+hxYmy
0W7uj1f+YVYwaJRpDAqrRgH0YQth8GlHRG6PBpRQMoK4ifs0NSO/cd0FOvwG
to+C7M2Bk7E5EW/ICUdI35Lb+3hwlGz+fesdoDJplSQex5vs0F8WcSXPdT9E
iDz4SG2kJVK5YIeOQljM2d2na3bCxOIUVdRXCQPc6H/V0OuNWq5vufcTbKs9
R7EEvzcdD1Th2AEniBG+oHAOvb0+iNs5zb/I+cIhMnVUzOhb/F7ScUOppZdE
QjHnONpo+4bfYSr58TUrkGHYUBKzbxfh6GA6/dTRB2bDiWDxSt4M9dWm6X/5
SJwD9DyKiSuEgS1tT443nGWw8zpbjRfyrleaUgue9VtkG+5Jx6+MiyPyutnC
3JMcxbJikNKgk/n/Pr/tXyUfOaeO8DnBbvoRaGue++/1a66m6cNTavJd1VIj
sdYbT9ZOGTqXMNEusr+A/VTfnQ04g0TC4zQjIdwpHSwUi/IzpIA6CTn6Up1m
KFdjgfLvgcRKtQ4JsSHF3MFwZ2Ee1qBFSEiR4oLCo+LMH59IUyeDsdosSdBg
X5sfY6nalWWNIMYMf8RegUqBGgLAdOdQSNtUmpmsRdyOYbRaOcrWvF+USM/M
IgOZu1SS1u6lFh8tEHe08hw2pkBQHDwkBWFmLLM1WWgAVFkWK1rgQWQn6G1n
LY5iU7ccE3pU3j7D+TOXsCGAAGFPqH1c5FilQz2BEmJcSmsHiVsPpD7P7fJh
B0h7DrO5gMTYcDbrgVGtpp12P78TmuauzCAK3vj5ssIG4lfEuiuxsZkIlPqb
UtCgSEJ3sJH4ErvSgqtv+Wp9ZGstlThPfsTiGlVYbZEDUIrbyPQGMEZrLP1i
sOZoI370n767cMw3ucpWuNMvroD1H/64L8i2NPSIhi0IW64NNTyShT+1Uyna
kDtQB9W2d41SgAqsCfy0FunqUIsvZLXICPJ7S9CeqOC3NnVqB0PeBV2mdzPn
ub9WesJj/4/T53kYt+t0hHPTGkyFTCawNuyOaJD1FFSB/aSXG7/sxj+9hHM8
DU0c4gF4Ug5dCMpWOk8X7LI1g1NRCm8Y+4yUtpnJMimTkCSS8lJrN0aylsRH
GB22LcOQef/WiCfMHoc/yqzhWLewJqgeHW+Mt890CeH9+lghFNJEtuXSbUg3
wVRc5vX/YF55fTifi7N5iB9RatkzEiovsN70KtS/a7t9HkLfIv0YIw1DNQft
EyREaJ+3QnApg+gbJJ/+Hs9LWB4/9rmnOyxs8U/8e9azrlQIPAYtIjWdjmzp
8sUaE6ChoetLtgcR4E1OigRoMs5EPcqvm/nJoY//9hm38uZ7Nk8J8i1qPolt
SBGll9EOKCBrUZMT0pUlDQmGjMMWB9T+4Q3j95bbTIa1Mir1jmyl32tlZoTM
QqA+LTl/gV4J7ORdRYI2Jmm6tg64psPdK6+9NY8KbLGz7+CobDCIU/UF52W/
ykuKa2hJdnMbjGGyuNflJ22jf2diDQMsPyTzFK9mM2V5a39GL/YTV6303d6X
8zPPZXOL7nizU3AawKvG/aOmjcFzImb5riDrC6m/ODtUNYKh4IyRhwtjB+rI
MnTgAst/rAguHfuDorQc/pOqJ2W5uD2T6j3soiwYUmdhVXWgBKYqYCMd4toX
fWL/bL6/JGMzwat0DodMaqEOv4vFDsLca4W9kdnmHx4hlpWIBkBQScRKw/C+
Hn+WrOHslVTZ+OoTDXsrjIDTRqF4r5m3ueAPhwT/tCE5yD1vqmh9zZiLHSSn
lKsjxoTqXSN9w9osGZU1yyRLUWYw/4YbYchp+qm2mkv0uTjbxTxip4QjfcyV
PIK24PeT0CvMiWLXGPt0winGqohIx/HTWLk10zbqRa/afA0isNsoV7o0iHhZ
ZyzFdyo1nVzupWVnNh9+UkpiLEj41j/ygVM86NRP6Ieif2FSzBaE5h/sTVTk
Z43ynfWfoUg/B6BP4PUNU9dmK6VMOoly+8Ms5lRtJ6A4Sb80bLR+XdDluOaH
kl2S98wheEj3YTx4NGgGCCdDp2gKt1YzHu6CCA3lbJjdBRfmTjCqdvLbwn7g
Z56/jOTJwiS5DW0cl53PqQTCYbltlSVENvbpSvD/gS75oOMRwIAp0nQ5uKrR
vE3Tbwvm+bcatphiqdfi7sqp40K48cj4ki3KooFJJZ58IQn6xbnT4ZR+zjDF
OqX3SoJXoBwbYho/3ICn0odXnDWr8x81jVFcx4mIlblHPCVaTu60E3x7W3Em
TdXs6mEvNAOYsu4OzNJptwOfEWF7UMDyqQt+ACa/6j8s4WTHYoXUmJyz7Rpj
3On30dUsud++f757ngA4PKxpw4cOXbSDZ72j++vupVKBseLBZYjvbhn+GG1B
+zsCUbGMEiSDfoz8iWsSxC/DYD1OBd4HEHvutUaQyfWnGt9JUFSSFvOCXQuO
KJfGjR7NHp+jCqz8IE13t599ZD5Vqz16bVhnWklvMdm+zTD1YaCSBklv+1FL
XleYnTgowIRtc3YN9pZh1PPxwW3wOXNTC0bDnmhxTlvbTHHAH+OfG71sKBk9
Caf6rtmjqayk/R7WCfyooPs0TgwkC1X4yYJ2Q1DfjGDQN1VATQoWDWopruoQ
HO0XQ/GDXHWSisQoyP0DeMV5nUc83bn2yBxqIPYY+MEnlR+DxdaJCUe+D9wr
9NDkjyM3Ef9tu1/INupkeEJYE7Up9ad3/YP16BEJGuFb4D3xbD1RfYPYrz/S
wAIt3HJuM7V6YBvSsaQxogDIcGCL9dnNCtSkkt04scCjyo8TZsgZ/STDCBJr
X//xV2lUfmUpjidZZS8xf/z5+WHbyy2iMNRk2ID5I/4EE4iBEzx/MFEagNlb
Kf/TOrOiEpHwtT3U7qYWFcFzb3ao/MnzBrqo1A01jrcbYbbvw4uulQssPnf0
paQ+pVkHXBfg/ARG1TZ4RLSeNlyuwqM+8Mo3NfncPtdFFZZKJv/cWNsAmveJ
7E/kDClhAMXy0KWT/2DrKkC3RuxqKlmGn7Jm/KMbkUuRfp4eY7CxZBDgl+g4
bPoCQbemxlYFxmDIx7zXWRnHv5HHTFKHHXtFEnAVyA6RzzvRMES05sbGLafC
WeVgCzmetOeeS1l3f12qMsEOsfENnzv9GxsED3gqfZbATbD36/DR2R3tZvol
ndngcNVwuMJDe9Q9oQdx0o+UeAuCr1BrxUJ4Ns1pHUyT6cjX3AvrevyafLcf
NpBQMh25HdVcrhAlqHHwhd548NoeRvfC38Ph8G59MVXZFhLa7rbSRxZD3NHo
0fXkp5URW1DeImDDLtMOSOEgS1HIoEpuu5L0/qkZX7fy0rgn6ONAMNBC4NR2
1a1pny34vsgiumgdBQcHyaf9ophg077x9snbIaW7ix7N1rdmL0bmqjMeUKky
t3QsiA5Kms6xWjczWyEViQjMZButadzSVyd4un5sw/RhLR7TWNGK4DXIaFmt
wI+1QDMa8ga4HUXIz+q4oSlKgSXdWzs6sdASeAhWUj7Os6oFUBi8QqIkx+lX
j3qC625rIu890/jl0P9qFrbStbzK2g9uBd7XuAdGhRQvBkM4fhDmGv55J40A
MoEu+6EbLIR1HLXfolnN2k1JEKec8JjD9/bvO/8v6lx3q1fkjMop7T41z9Ax
nNcdHci9fedb2CoDIeHGKyrpuMo0q0nwD9mxxTQNqQCExQFvvMHo4GkkEL5D
s+c6cYV8YBhCDprV4SybrdCygX2v4EkQ7kLRMI5qO0fClIwerTUUbkEQx2Sy
aFshtFxLILe9pNEwpIz7JSEwEnKz8Q3aGbpDFffkeR1RsGsQzn8VYRUtAGhq
OYxYHfn7CsC/DnpjM/YDfCQl7GqUssS5rJD917oI74Ra1zRXcGK/KEjImkSM
ytS3e/i74bW6Uq08JcyW80uLMitzmYeswDb7nXHMIhYgOAwSwFWv2rP+CklT
KZa8iaqpZilP7sphF4El00hjFfjL8mFjuLV5nqnAuQHxfzX5Ld8npVFeTtm5
gDeCkt+ZNQwmdtMT1DA8w8PqGZEl3rYl4y763qwwaiYprf/5mo8Bq99/GSg5
A5PprIytYNNr3sXR8IC7uO0EgxxH6uVGWX818gBKFvbw2jTQ4RWwTSd0e9SC
Zax/YcGMjtzTfTLZB2yRrlk1QLTpEBWdMw/nCALOzxMmyDfrs5RePXf2rm4j
Nn17xW/tkfW+CYldfnqQ9XLuDZ5smvfAZ5pCJqpH5u1bbfwikh30tpzmL7MX
kMAyAr8cAt4af2s5Kyo8+PG+lkH3XA+vatUDgvFrl5aF0/7wQ6rn9PoeNsbQ
2E4xDrJmn9fJ9h5B8K8x9uKIMvwobwdCcCzFV+QGCquXkWSqFwssFaBPAg0k
Z623FUusluu6G8USAcJhaxB92zwcVjx0s0zyf6ms9+2aGiHkuIM6xzq3B4DM
2K6kVYXIVtgCoxbEB4IODqiUjfrhKKucAlfFvc4vk+9JJWKlt43SSvCcE6P8
hQltZEhGnoj3jb4Z39BKR+0qnt0ah1MSUgvjR0xCBuaWiF/CM/mvZFNNAQ2d
1KxzxnO8gj80KT0Z5Ny7EKjuj7HASCcSa4Scj9Bi0sE3KVu6sUjYVTeH6PzU
k9utepTPeMGvoU0+GG343jgBOrh2HONnfq8Ezopwo3GdaORe5QrQeCvqAo6s
vDc/QLx/K5fh8OgUcR8a+IoPE+CT5o6XPWxCmwhEQBJIot7iN3Xxo2aAu3mZ
+bKIGhDlsJG0VUhoDA7JHCU8000hS/lF9SvXxt5jbjgNF31jqpB1VLwDyaWS
BH3F96V3hTW67iuKPE/BhTnlu1hxOrHv8pXlKl2kobmMzr4TDZuUe3tzfYop
Gpwxi/BYxFVnpQ0yY6DrqpZUwdMNlDtLbjymIMaZV872k8IDxo1iluuxkGW+
QEQu7cm9leW5ODG19XUm/qWld4B5P4JOApgmnv8Ujepmgv/mGzx6zTeMtoZz
SeWzitdu5IMwOgd7LLP5KroY+cUr/qIqvh47QduZZ8goC0wfXXP3D+3WfdK6
26hW7njzN2dc3hWxX2vQ/yAsNcW1mUu6G4nu+wd3j511HxWbXqS3sOD2a7Pt
9wPZ0CLzgkMyRCpHP065zDouFVKazUK+PvO/qD2mZ8iQRRDEKSY2sU6tvd0Z
1vRlhkR2c2SfqOmcvzpfyZDN9QSXwK3z1Kk3MCC7tcbRSNd2uyIhG6Zpayk0
YY+J+sEsVjjSdMImawG49uyjsDqVgVLHx6l9HDybA0g2JUhXEALDM0RytDqA
DrtW9f92PpEzEpSvvBBtU969FSRs8xuz4QqbgYzKhJax30ozqCNKvwPuBdWU
ulwHVeAYnonucAwu718HZLSzYZeos8eGyrhcUPzlTVTYdHirhomkZKL237cr
PKl0EIC9SpLg2lgmbVtcM0CXuXuctdP7v99OT0M6mZW4fEDy73MckuJK4t2R
QeEo1jcN1y5sNN0xqOM4B/ebzXYbVwiAfnOsD/Meyo68wg7JPMDpqECysQBF
SJJS1+z4rHDTAMpKzGCoffrotVF0klR3UQzARIsy0w2vybKZwXUIln1DiURR
FXxR8j0TEpiDdeum1vBf8+lmLI968VZ/I6LRfxa0Hldd8W9YuPaSkRw2LR9a
tR5B0Nosysl49JcXl6wCn1LgKquOzTmzuHX8+3KxiPewKMi5pIjm0OKwx95S
qwcSwqussxI2sjanfioFQykLhf0saqbTi3VgoMhV1GU/VOi7XjtumcKdFhda
Xe8WvhZdNzoMvbq1XRoPRnieBTtP7CVvkL4IbTZwYG+GwkvJu1hWiTcqVTf4
Gq6MjduFa8W1YESkHCJoWl8a/HH6OHjXl/5LeNKrFldz2ShccFazSEAfKV0r
HOa+GtH7SL3ws3Fj9V087qVpSk+2ZqmjXimVCHNxiIWLAnJE+C01Hvd7fg7A
PoKBSTs/8/Wh47JB9MavzWRJvuIcBuvgKYVlisuc8Wm9MUFvlWNRJ9cw8Jjx
GZiLVotOBGvYUrppp0ey3VxjRfArOCOySqSNJlAnMrsmJ8raSXOSHmLO5+hv
ayAN0Lx9Crt2VzFH349HcpmyyCEdy7u/FK5bkAaMbuNhNEfPeDojzCQSsZV2
NlcmZqSrFdfj1X5DXjZrPskULtZHFMQbLwOZXaczdlNI8sglmiW+bwxhWfRW
tIXyDeQ+GVA2PphxX8hn9T1MzuKJsSo+va2XDOAGKV9tNOG6V7oy+fFzN+7W
0H8PJIaUeRPrSfjh2HltTFNjdPjKp6i84BIHHLRLOL3qrA24pDTiV319tUhU
MBnlo1qHMB6A31HH8XHuohBgJZ3Gsp75YzY36FOjmBH/8ZKs6U5LQ6oX8ouj
rjlypICg9lG1q7wq4arsJpkIre6zpxWtj+p6VS26wTWF0nI07waiySYUju1D
4TSC18V+h/qTs0exWh4rhPHlhWdnKw+2KlguoL3iW7rnfLhBL16T/wUJg68J
JwctBwRqiObcZfB+QRQ5NxWld+Im7uroOJYq4n3IVAXlJOsvwGzUx0BxAXNe
38jW/egWz6VENdYG4r3nyTI7a+HzBeOV8noQuCLMYHamBzdJRLOt+4CXPmRI
G0uKBTli540Ou7oaOTjfxdDlj3vCEhUPKv/2b54hHHEfK2OGRj87Zpg2LIPD
Qpw2Dy23RoyvdM31pfAYxAV260/sTEDprhh7UDRFoKv0lWQxtVrtbmvyp9IK
luDvNtM+CQA2xWxkptVU8rbhz+uYxqhrooXBPDTNL5r4/J4FrKnV7LncwIRr
5sG2K5SzKXqyPqXBwymTgyqa6pJW52bvrl1HTG9WOkQtnL3pwjOGB42e+24J
9YIeB6L8bSYXKlmPS7LRD7EivDVTvm1R+59OPF+lOHaI92OxZ4kx5CT42ZZJ
itr0HfvQznRIVwkh3U95De/bgJDDx6/gevj7UZdz3tyuZ+SESre3ji9/GhIm
HcqV78oc3hFdGRaIRqZXxCBkFXiYA9tx2bTLSmqAsCVrMUjLXBqp0/yq99js
GfjeqH5P1Vs7pAf+ojE1VbHUq16VydDf0JboRX+DEOMaMU91Do0q6IsaxjcW
B0FEsg/vpgqtvB02NtJf7DxSOgLnH6jJEpqUEboYefJ2gHAFbs3tD4SUzcv/
9PHO8TxWr8/eym4pbOdMvBroFv0OrJOexsGWojNpeGfpgULfTUiMWmDNyXCa
Z3utyVJbo8RrsC/y4aLrERbrLCBuC9+xPlxIy+/o4xlELoI7wZY4ueavxJUr
JIkPwGLo7U2V+ESbZGO7pdFH6tlTRocQ425ZNuo/k5uZVoJt5uLTb5+HBG/X
lkoXuvyH7LS42pbyr0CrrcKmKBMw2oQqWSaB2Msr3yeb95OiLsYFq9iaUQSH
VMEmDQAk3d5HMTpdL7/oG4ftz2CqsPYOdOF729XR8pMp4aPUthjTuMJjmLy8
jj1gQl1XtnySjOGDmtSFnLHeWpYvcLizOZJV2XN8WB65DtHvADaZUCL0zzX5
D5/iAMVa221jy6j5VEVYOfZdh4PKtUhZkBmZnw3FzlJ31Y+P8N0zcc613X6/
2HlRkTZi+9rxjmziHuW/B4MWUj1fMIzOTZijhe3uGZEitT2e7kH+Dik/o2kS
axL4pD0VCMjzxNwoo56Ws8AXbRPH/YEBzISae2fvgxbC/4f+ZxTX1zc8Z0DN
WRVKSfcp9MEw8JFJtzTzNWb+qtYqxqUYWIzCZVKAj4TtlHikVsLwlLetNDQE
2AfJq6cado6IudM+W+mHO2cLHM1FjQ8OdGha+BOHN+lYhLJaqYc6OjMrb7Bv
HEOAFQu/ZnXy+Td+8UtJPMBH5ACGt6ELis/xDTd4njo3LqdaAV6XIExAwLsO
DyzKiFAxqbkS4eIUs8TYTWPxgxx+GZoh6FwWOUSYiJKfLVkoLyiwWiqrkIhM
DjHwPLMWUZ7okx7wEy8uTLHj1BToYJljGdC6nyYthPWcxP8OVGIBUJSSozgX
3N3EcWlrFS4n3jjVkDjY3xvu+RVtd/CgboyyGnaDgFAwLs/nB6T9adgmG5zu
fc6nXdLRt2zXXLhmk45n+pdDlQmaOFvMb5yxEF0H0tvjBKsH1T6l1InxuDFK
8zFLCXPjAMfyHJNzjuvZ3sJEwJ/1yhgo6O/aZWrW6j8F40p4eGV8JERRyWE6
KDYVATd96MnwiijylXx3NY9y1vhbiepmQrHFG3tOjGuScEqYhkElrVzp97/S
Mhg5iQi5RdgDr3cJ0hRUKJHs9viEDS1r+YrNEkPcIvzdo1096CKAqkehjITN
t5MRlwP69OAT4+vOusjpbsJGZEm9wsYrTGrzM5VcD1Rp7CZWv9mIfwoQzIoP
zJ+Nan8Abdi/tPqPSq7Ke4O6KzHHpwVIBMYNqTdY0uixMX5yPjlebI0oJ/78
OwJfgVIsN3NuHBQVba3ebojzFt61v1sC/kqCTw2hNC7fbiw1/U6z+X9cM4Ix
mmpU5pstmNIErtsS0jdZAc4+VgjUqHtu9XV0pl2uybAuz/LIz9o3O0haVF9Q
J2Apg0qPM/ta27wZ15oelCweakvf/8Q8SczL8llQ1ObAQqjyp4ARf9hfQUP1
OPBkT7Be9prPwwwBx1aSza0yl5NjLvg4Bdtn4YYpWBEgZWU45eFsD/srhvV/
qg16g8TZOyLaG8nO3brSJDeelmb5JX5JdnFpkAhZGSH4n1c2DhR/9jLyinMR
5LrD94Zp7IkDP2ZL9iw+5Pb/pjGt6OjybGUt05W36LGnns9TUL8dvd6I3ts1
8rCLEpEzSv3B13SIePktx2Nd/Pz0x+BXZddxnpcDdbwMMBmvWJrck+9kmEzk
0lIChWQt6r2ELCJd5k8adyuFhw8dwn7EaJooSx8bs1Dw0BP/OTX0WKCB9JsW
igb9fCiH+hVld/sKdGO2Fogo8J2rFYmyZRRHLboAhyUW+Km/MsWrlZoIn/O0
f3K7edMDRrawrnQjmgTfDpGUeWeNVXEw/YH34VAFi/TeOSuPmT5QEozHxG46
1hxOVtMUPkhLmj+aUGayJdUXpy3uNBRiOVllhBIUqWAN8UKvvoDSvt5kTgO8
rmDx4sAjk7SNpDFdNnZb/pKq2gpL9/qiPJ3FlLcCr9uuZfR4wAALcENAj2rO
FA71zMKYAvWCHvBE4lrrBcnVClH9oAyvgN7DJi6tCbwdREcbPkdOMbMsc8BM
pmcXuDr4PtjJ/xhjAoYPYa13jy4K6zftUlCq7TuVT3mcYnnvfN7gdlRT2Lbr
8Zi9EzXrVMztSHgQRAUYB9uiXv2mUP8vCBv47gGEibQK1zCu7liqhc4GRxGZ
M7nR0yNODA/3uMm8VrNmflO9SC0w3SMari7sdMoKWDh+0SKCty1jcmorrevD
JMcsZAiahDVvS3dc/vMBqsvyUUk7l9VTddQG2+nPmlNfPk9ebCaxOfby2axW
jqbP4Xj4oW2OEkQZugcJVZAYDjEvQThLdmMWoXK/uT1rPwi+8Ct9ssu5JYAk
OEZ7rEw6YVWIWFlgCF+BseuDorHKwtYYxvI4p8ZMwPtbUqswjvXTIchgnOAw
E1ysy+z//J7tR9++rHjFZ4Ox+0IQr9G77EIaHxjQUPnjP/6thrBGYYU0p+62
yKD/Fo8Bq43bonWCioNNHi1iQCUm3Pl7iR8qUojbW2fHNZYCmFB91RuY3JMK
/ZJcb9zYH8nEpdEqW8YuVm/fjlaHJTJYXkEWN/xaR2vPKqHN4K64Yvp6q5ap
DB2xJyOPCk8zaB1pNeT6ZF03ykgPYFf1bCH8pIykjBRqPYaHxzYSVGDP+c/4
nkgSbJoscOhPGkc2QluzkPVlyWUuVIjAjg9BXtFbIdU1UJQlZ3rW56ESQySG
MWU3LU4nQW718IBw6sXzNQ7IeaiXov2drTH2z2jNIM5cm4RBJjbcTvL9OPzD
YQdimh4GopCc8hIx1hGRhPWpT1Ib9YrM6vnqh31s4htQtr7sLGP5A4Nyi4A7
CZSn/987duxd3ji9QvoSeuOILFeW3xF8FUMq8xINWJIQbIX45K81ePVYOV6o
VlwzKOWTKxZi+hWm2sSMMqWX2qeA9r1JHW/ieNeXsXzynqIspHZDGcU9U12m
/lczbn+k6BrxnNVMCP4WRE+uuwpqYpZd0cXSJhjy5mje3zSARLL78Tucj52N
A1LXF8AkM775P3LafbOzct85dbe5aKAF4vuwLmkcRI45TgJuL+9KKLrb0Vdp
+Y7TCVRqmWSkhFrOpap4GXDmDRzGHPB2rYj1pUahQO/q36Lq15a0JgydjR7W
888Fk4estT8HmMXTdlntT8Dy83N5GHkhpAXil4msDgoF28uVJUm6IWbYvGTf
BXdhqCapb3fApFTWhcCeAIhGsyHyuRaPrgF1U/LamFWZUIwoAS/30527zM2M
Gl2S116nHTPP1nrtKfju8OsnkzrjXIve/ih6AA57NnGPi2XtUKkbl04pr0vU
9FtHxijvUf6AlSeBu61o3M6fHrIwAEeCfTLLeZVfyuAC7VUx7ZTDHNTI0ZC/
elWVhI+V87AyCLse3gkm2ik4QaM5dZc/8OdqoOXyP4lPEnfQtb5j+RaAnCDI
UQso40zjZr/AU5SSBscDbDqJmrfGT6apD+2hxNWhnO9kvvssCo+F7K3U9ddk
uBsKYwWwkb0zBhV2dyrK6qPwLTrWwoaWYOm+tLNmC2AYVy+rTLX8mmNvWrwU
w4BC5vyEXM2FmbG/qmWbp8313guRxEBc93DLkt0bNb21tC1wjLhoVoElt90v
7zZ3gpcuA0RVLDVhEc3qLP7O5p2/+8K9yPpTeC2rfv7gB3tug5fnGbpe3cSl
4pw9aEdnST54mtYEu+EvVAh594VkgtzBzjsW83jneoBrXxaS3kJPwIp42++y
ACtqJ5iyoGHK/OmKCntPV6kWjH3Mk4g5kX46dLcq+Mg3lSjgz1mMxML56PRy
ICxhRazZPXTj49lFIvnSBEDoNPXOMEnzmoloezFzCHJ8K/z1pHmx7+qAZJRV
+Faa52/jogMcEMuMhkEVj/t5ecwyNfU/622CIE/Sx97dtUH69SNArLumv3mb
aaT3gpHdQ4Tlgefb+wh4TL63T/iLTxFVqmx+AlgjQcXjv0nbHZXU8A2RV9qn
TCHWRE+BBJvbqhehqBrnqrU2/02/gJTp9TsEjcTAvKTqVdtCisXVAHpAk27t
bQo0fbzPmUYDSNKW42sjJ4+iROYcJR49ZKYI1cGDUnm69QGg02DJyM4bywb0
ttW27CUMBgm92o+LsgfoU7qlxxDkp6b+MOBoOrCiZ138qcNWJARjSyBHGAhT
U+u7ulMmCBIh7XYsikNZkbKxGEO7yuXJgNw1+gtBbD2GVslEjA7hZIKT6wWo
e9MvHiK3vHbBgGwcDWOwMNNJj+Bbe7OYKufR7Ks7ek0wk8bHI81jXAkX+Muj
+fSgt/YZ216ltUbozgVJYv+7MdGGVKM4DaeiV1m7b/Xno+OCcnlxRDBvuLDR
4W0TDoNopiSqDC1jbCdjjrd3c8zIyT54y10rOPSkjzBLWwvPIOCVh4lxO8+o
PB+FJPL0yaMW4cHPEhLt40wXDBOVYW7SyiV7BwwZN9WHRxgVfA3qlNB5YJpv
exJSXa2zpP751rSAzWbrTmIUUa6qM5lYAUgh142g3jcp4O237yvTvwRAwKKO
QQDrvFDP661uPFC00fdr+ovfkztTqRgdPHXRhh/Rghg1u/lsP13GyF44e7X8
3C8ItXUGwGNC9NvOC5xQvROxW47T/Pbdi50z9pIsRzuNA7QxiKmNgARqpEGc
QWXNoGPZrL4sHAsRYuE60PihEBoBa7Mv8DceSJD6QEiPQmKrXRgQuAC4//zm
4H5xdbb4xTKFSbnVYyxKYa658kzk1x+DZ5M031lK4sMt0UirQKq92yVSuY49
FsAisC82WoIkHbcFzclU4EzTViPvX8mw1nWLCPujLYeehaEm9tavXsOUBHdW
0Er/jhzd2atPr8+MM2x1jYDcPmNlrXYP70ehX/71W355w0WHl7gEuKmWqRZj
0c0XPU2BYLWO8m15qPwXo8S9E1gV5+TYSn5uGuD2KBefc/pYyYMKsY24swUY
tJAE/eleJAlZVsOfu8Uq3oDwReMWom9TeTGGvNTl5yF0P+OZdkUAQD1+HPc8
hkL1FtoFTviBhGJXJNqL4dMuZAWgYQ9c/c2Ivdmg9T7T2tKm21GX1QHkdrja
ZDWIVkRPMG3ITQIST84dst5JGo0Cvmtjk3OApfy+7h00vaFBCm8VZegs8+Sm
QWeOoAPlejJiGbVp2KZ79QVSaZrrOmJqYAsDf21u83+IWbQ7AJ/NJTNbEi+m
YOUIzTj/4e++BTZyWW8f7KzGKlO5V3r6KtvnNSUYRmK6ACnOOJ7ZjRfYmMtZ
x2psEtk74Yu4agp4xjyyhs3vkjyIZBkHkt+fCV8l5zd70H7omSdRAuylZiLb
bznjxSeZmyHrvlBd/nm8pkUJN1dXjFpKeMaHXLOK5czdMyvwkFbPaJ5GfTct
ApC0TztYs4imUQ4ECKfyvoAu4awR95rVpTfoMyaApvG2s0PvNJwuiW/7kzw1
e5WGI6jgp4DulDT1hZ7vwMSKE7FQoQVLQFInUQqEN1MDo+T2G7wfr4nuGyYu
J7On+kRA7FsieeAJ/+VIjeY817brD5wknFiHOI8Sp9ejOvP2JBcfItuiLsJG
bSuAHOd0k8XMQgN+BlS+EP5KxMr+goEwZf/VEb3lbQJLzRlbJeAddz/2s3Ly
K77G538BQ+dK5W1+F74yQOl7JKWZBotpx/gpxzfVZVdhbIhrAtH2gTI5YJkd
L6SZONeQN9f3s36Kq6X5+pqgGHYGUGJYqWELZlP+CWcwK5nO+QQ74FUlybd2
mWwZeHGNMrVdHfIIbWRDbRlH52KtuTGmTlI7RpNFWm5CFy7GG0/FDpU8K5FJ
hVzw9kNXU8BW6KJ+u862Zz6j+I3HiL211VgTM6qo0tNrBkInCvjkkAqU7Wmk
f6lU/DbScjpZ3oC3o3mnxqD1Sr6caSP/FEqlgraJbuPButaEZ3F6Nps+PfUY
DPeuiYRUCJUi0fKah93x3hAMp9V5XE94xOpePgQiJGUwA0dQw97pWrBD9mSe
Hsf2pdP/iLBNexiIFmOhzdrSij8EcHtiWljlgQpXsPYtGUW75sjbiFtaXZOe
M92J2IBxxPEuH9FaO7IenAMv63C8cNGgHTJFjECWST7Mx3p34GhAFWwSEoA+
VOR33OLkj0rv961pmyBLpY3fqan/71nvC/+qe2L92n2sBFrsUU4MdfmSKrr/
OvoyXalAbzrgnFXKpvRnkIQsF67WW3/wAtZLtPM2+eQFwrrFmu+LukxELSUr
q5i77sTUUDkRciIWDgoZ8LNvPz0CNyr4UFDA3r9GI92lbjNq6mcM/hbMOzhX
tNvwvc+f/GzQ97mjI+hGLwua8dgHavHAyTEDvubbC8XfcU0uWOswT+01cKs+
eP8X75RE/cNDyLAnBor2ACLr7s+t6mcf7GcJ298aYRkq3wCacIwDP18A/22B
82bHJklTGK245O9u65uLDHU875sVrlqWDCoanP7ka4dtAJYUZnwjG/Cls4yR
mMVQGIKyMi7QmpyFIjsZnfm0+jKeBzqHx09Pya5xXIJCtV+kSqzt0zgRoK4B
64wjL35TDHE3LZNNBZdoqhNsKeU/ta8Z0hXW/7jJ07UP9EYbuXsmryO7DgFB
4/FDhmqiLzjwoT7e9gqJ6w8V6FQTXkIp3ZIne1szmg8YlmOewnvI8cMMqOcI
EzAgZTcIl4VMCUj6L8l1rpSC6TZXLQzIBVQ0PttnWyUM1P2cAEndWNahwm1m
Lp3XWTVHWcfNVG9x34w1DLKuBr+E95rZwLJXhzwOCeuplcBw2aXUK1AAO/dP
u5rS7sN0ksKmioXXqiZMqBSmBBX3imkK2mq/5VDC9uci4ciTUGZg5+55DI6E
3uPowG5xawKHqiWUn5twa9Z/brcC3PZKw64KaAjV5h5EkllQZO9HwjybYSya
ykDBU6d3xZc4+VAZdODvLrwZyvJnWO0jTpnxKzSem6HKTkw0u1F5lI9yzTqi
g3LgPBC/Fo611DDBxEE9ujpfb87R9npFzTPEPRZmElCNDQRarggjowV6ShA0
bd/xEM9vtCQkJou5txIUeac4FC30/qLlM1UiGH0a8FqkkaQqp9uPibg0K3ak
Ukj9AiM5gQwXIxj4v1gzManE9wqyYZYXDfqjO+z5GkSiy97a9jf2TXAvyWB8
iOanwDH+oa4GNnEFtGuq616Qxen0s7gH2EXG5geF8oaPqQd4LJUI49ZGPc5b
QjwBT16UIZc7KriwxkWRWQP6coBRgn9VGEFfJB68MwZDzddjCQRqVlAO6iAk
9N5RpEf4Xu9sKNDNmksALfJ2K+OM8ojLYYaTYKOixMs7rUDLgv0KH8EiCG5i
KvuJrm8I9iJTyhDzG7LiTgBXdwbu7iKDzEaj7yVfw61yxkAnPTg+og8U3VZs
3aqobKROpyydJWTWazPM6aafWSOFkJmW6qsbwMh3jTkHhdoQAEYS1XTpgnxS
gUrJA3ln7QfyK0a/u5+W6QxN/cv6/BNm7sCsApDLMCgqYcWiTqsB+cvSFrTA
Cizb6asluTFh7n39oeTNhWswK5ahDm6NgNna9r7E9aCj956QlawAsWrlFgph
ig3g06hnWeaVwssM6qi75Y1enmpTbJIh91IQ4NkMfSid5LZFDnthyBHTbwIY
Bm+sMIKztrNRuc0/ZOdDkr3FaPIoq+mgliegaBcnLDYxt1tx063IyQ5ZDQyo
cnWQweGlJhG3rt1LCCSPvtdPs80vvfYLERg06oc04enE7CSsTx9WOfaUOkR3
bReLlpLZGCIom/NGiwOUxJIsh8+v3Jnw2rc1iDcCFxdU11xw7FOtpWj+D1pG
vAoy/3DlXFj9euZD2sMGJZAZc1Jgaivi5xRRDZPpODIjJ0LyW96euFMVHDRv
fygeaZnbpXz2qowGj7ObBxegbOw/POJP7Y93ZaL3CyZAi3fQVlcoTwB62VUH
N6XsiHaZrZrLq24KJJcM0TYajwpywF2IToOhj04owTZZSqBQTJHaMWHdrR0K
W7a0FeO2+ttL4uZjYYOvYOWZtAms8S+a9Hd8Ur6wtxlo/Fwxv6Cd0XsbhRR5
FXn+aci/OCCcFcI1FQyDFAisauP4QqHAUbOFiCb+SAOi0CJDvsauN8Llxebk
uRagJ7Eqg7Tnrrj6kXK04979iEB8siXXwNdpRWcePYnhN4y3/QUFokfWeUgU
T2LN0K4wAihMN8S+a1FtGVBB8IpvpGkfe087pbqydykWmsobowO0zAgxf+br
DXHOPe723k+lBEKFq76Z6upf+rCQjIaW/KzeQ8N6mtCogweRSOkQ0gOlyN0K
1B0OCkBd76fxFPYatua8UIr/Wftw6pWNdJFZ2jMHCANYTs1wa4pG9+vM8qZa
qCTNd6kVu/y+qay2ugnzGETln6BMM9/pjR4HasFj5mMxK5djTEWmLafVjfrr
dWO8hLNW9mdv222qCWQozAKgYFPE0DPFP6JiUL06DYFzvay150RUHAwLmXzz
8c5sT48ANEw7XsKT6eN5DeykvpUqh6vQsdSXXdqadXAv9fVV5aMiHZKNgxlz
0WGu6DMGOdsGGqmOY6dISdZ8ATDiSBB4XXAgZhs9VleDR+GBdpRSg/WmL34E
lmqfuhzIKmRK2kdY3IANtXAl7HxJUjl2Yj+w9D3QrTvY6jbOxgwnZDlWysqC
Nh13YCfKhFlzthC3rlDEl0U9qokJfndNCdAk84R51BtvrM0jNISAfAHvUinu
JWjRY/wR5tz9HHTb8rBCr3HGPnVxNIj8OZri9gjHg0Tu4R8Vd4cSayNRbIxy
beCzKPMp6pMbwEuXm6jZyJxcsszqO695e/+4RGhXCtNM7Rh7PW+CI3O4e21o
0IdzuCQcaYw7aX0ixKRe53YcYj5V1ZyFa9J/XOvdycvuZOacdEQNV+h31cXy
8M7hWlwwpzBB4sndpAFvRZU/cRrkGlEQg+HjoHIJ2l+//8jd3C1/AbpFztdT
BohFqt1T61Ul/kfUnoyKO+Po1nNbG2EIXjU0kRQjyNGgiP9ecCoMdoM0lopG
jXPDfjSwFH6hpKtfPey5l+Tw6efXfWSMwj5dGbMReHQfpwyIXQBcxEAi6pFX
mnwyYNrWxISVkCTciHH1Lox339FgYyOo7swJ+3NTNiLnuX2rfvbivWhQSVbM
m7gt+ozHNaaCmInD3Y4vE6qVrU7SwSNbCwMBCuQ3v4HrjiXSrHywr2DgP4Wz
OFWoLExTr4XVCOBqhy1zuQqYGj/upES7WLKC2GA+aLt4Eyjxsp29eH9Us1dL
6fN0MmK3OXt9/Sw2Sc24TI7H0YEQhd67Ac4cWz7jn0R/Pa5pMUpzT+FZXBgm
A0ZHNFEq0Xx7NTzlLXajBKk4ZplKBnvKKmK3r3yT/62tv8Cxal3dGZBN5R3a
9zZfgwtuGtcpiVFY2CKCUlIjWp6I/cGXf0HraXNezmwoN/ugXxear10m5SE8
NEU7fftm9EiMPwHiVQjieCZxlnSgZvw6NOXrWd3UrF/whC2Op64s5m0svIH+
PIJgixLzLQCNAny5ZQYP65ylq/WDcuokLfiE7n82g6kgL9QWy7siScuGDBh2
169cuR4txjL+iuPqTZD7T0G+TJviCxOfz9RXodcY2bYKa2jpi44euJgZcbc9
mGVO6O84wF5Gv0hGHeLjdfI7OoTpHzOYCeBUujhPP+LH29q3VecclAUN5kEy
8dk4REazqTfezw7yrDWw0kbty05LE7ETTdtR0L4JsHEvoQ3q1buGiuBRDgj5
tchubG+cCJjsXG6kI6gianAhyFsit3E3Ld6TQguyKZ+z7eDuU5ssX9ceCZiM
a8j5n5x06H4r1PLubLNKtQoaC9CzPCDbLmod3GPdK3GdVBFcqQgewaQuoj4R
ByECFRu8Y0skM5Mr4lCV0c0rpg4dEd2W2IYmjSQKKUMLM3wCYVCYQAKicCSg
0G6Jn3hCZG1u1qfqkVGLjH1U5FRYOrNeyem3vPqZtqZvwa3R51hvZwvf0Gtj
wyyEtFEV7CWVi5ZZrlegYXodCA8cUe8L7yONG3RHHydXD/76K0CTwtwP3ULg
OVov5Wlag3Eebwh81ajOWDdZmN1QF5Dr8oY1p7GJbge6JT8yRVab1wBofc8S
7aMTFpHMOX2STVQwxCkX4Es3Oro0bs9gQLZJt1W0tB418FjtvZ3Ky3QO0DoL
T76I4M8xaDSrfj9IlWCvW/4/C3VfBvEwmB506VaJqrrKecTb4BW6gv4Jm2mF
GEtQEsJh3RqanCWHQlCfFkj3M1pen1gbQ/y/Oqnze4uEtKtBh03o8l5VjpVp
fepUai8/ym8y2CUeQCbpfHboKUEmPu+r8KqX9dD7MOXTTm9D46oRygbZsuTG
YwYWgABEWIbKTu7YTZE66DNO2Cv5P0NwsmjsnYYIXMjHvsNp9xXTEPH6Wuos
pkSC3GygRGPIUnkySogH0K3Uir3FOHD5TYwy9J5lT1lwHqIIgHyJeJT5RJfQ
bSVqSf7SbHZRrRNN8Uf/+kH4G24rrkuvJJLwwqtPNI1o5nKJUCd/HZKNb77r
kfVrIyBAeNWwbCQwT8nm4onmFRmyH3ohov9gyWZ4snad65Vk3gikxNZTU/se
Y9zo6pjO/Wa4B8E+WZyRTHEQIdyHrb/r/T7pb5DMcXaDZchiwaklmjtGPlWz
tn6GNPZ2525uqVoFEm3rLatxkwy79ruPPKUqAB19D6YfetlFzQDnjjEuvleh
EN0iQp2VMBbeta/cVYwfD405Nw9I+2iNXy3LoucqKy1ondfdmAPiBcyq1SNN
G9WrVIFw17xY27BDWqAfu+sTw96f52dJ3Br9VOs0J4LAr274K1pk0aAUyj6k
OfLXrgihsJIwXs6aKSS5elOvB53J9iNnVM/bvWGs8ObEJ+3oZV/Y243iURwh
hlXkcJzFFQAzZ2JQycZmRh0zEdJTUpFCkF3HZpr3MRoRaKjt1lg4l2NoNlRN
+vVHW1yxnCn3AESQq4d2fJQC50DUJOsy0e89soWpCITJNVLL5tGIgdYauaSP
CiC8Cq2sXxN8uMEorIISg+UTELRFYx+0eShescWWQPC/1NlY+eZnel0V815o
mhydqu+Erkpsf1QQ8ScZFZJfAMFp9KVwN1VpcC+no3ZABkh9dphyxLHEvXzf
whWQiagZnsUte3QkVNWXNLaOu4SLa6edk9YELsRrJptMAL69N4Mki3xvfR+s
/m25ENiaYolt1uKDhTLoYydXkpCas508VKkXyFqfqphaET6sRbN5h/28ldwT
FMPz4+M+gl2lJhyxCeZJiUudC/rmv+rDq1Qz68cPY3vUkiJh+EJUHADUKV1b
a27+6b3s/M2/v7SesT9BFjUgPTX6LQ2o2Yx/Eh89rb2MmNMEpioMJfDpBNGF
IYOhEXMvCNv121uIcc4axCy+v9NVdhP/WKnvUCZaJGcShPXKTmRyHiPgFM1q
t66/2FU37oKC+mydVUT84UquQ2DpZjcc01ntAp0w6ZAbTdz/ouKyDAks7CSI
+iR1p/ROtVuRolh5DwU6AVRYXMRQIuHP9Al3EiNve3StwCwaBSrDbu++2S3q
bZTjhOlgkEL6RhIY7x6DScnLHwkc5lFA9OMJoGsZ+CVS8ZjBJZbwKg5hEE6+
/30mPCzKlBJJK/AN/qV4BLzdv+QcdQ0OGuKN8eXAEVHu1myfIONr4qqfxIrH
s+oAfsDKkINwj0Z3hzbADzIkwk7b83VxiF4+vRwRoz+jhaKRc5EA8QJZVCmT
zdva1EvYceIwi8gtNfSwulOhkpaMOjEWuvm855BnrphgI5CnbK6KWsf0ZvOP
jqXHCBq4Cfvm5kxT11xULFjdjo3JwTwERujYhOOsxuayOz+mHTDRs8YXNumP
FWM2HUVbmLWMG9tpzfxOJlweEI2gKh5STIUBbJBy2l+XgYhohtq5QyCna638
2Qr9YAdLaWxph8ib8i8hed6SC7ev6uE0XSmwQrQei3rqO2nr5wfyS/kvlx5/
DpKIUrPTCY+gM9r0+CxJC48NKvHNrNZjDQu74C7AcNlVXHsJjnXJ4meb/Yyk
6MTzb4A57L4OlWHcJRG6yiXZvhwGzk1Wif7raZ9IS/Cn9ZP9wUftNYnGiXEp
rOegpHFrXn5FfqMNv1NQqpSO4GvEqIgDs9ddgDCGlZqBZ35tg4gQpNeAbjGh
COa6wGbj5CewDSM4TfV3G8X0jUQVDtb+QeBYhhh6r2KIdUCQsmky2V2I1Uk3
HdLteNoMejfN3v4UBKOkB8E6IgUGExvhOmyqcdkiJ3hoVtjLhg1MHaDpHCzR
LmLxvwYb2TZ3r5g0AbzzIq/6MIISEf0HVhyg2ZdIABTyW85UlCqVIb3pdYxC
OKjE18G5F9r53xzGl/P5HaagBXaXWk90oK82CtAYCbzwIC4QFRtrphXsbWuU
JF0fMfoGy3yIwFytxh7ROfLuKdMy4BFPL7tPYp8hRqfSSYXvWGQO2wzyhyfc
+BFBxd4jakiPB5U0eTgmfImDThSM/WKZcxcXawX7L3EljYAP3yOQocyRut41
LiaonocKyoMMtsAdu95wGQWblBS2ygh/45K7lU6uBxwz8Mv3rw3IJ+1fau0s
E9GZKUyklG7pJSGJ0AsSrc5JRY5OmhK19wkLldQzQZHSYyuEuQ1DJC19gUDV
a9KwW+J4m/+iTmG2IlYtS+2bF/SMcqpUSlObaWj3OtmxJyrWdqXW9Y5mRqqD
Cq3BZ34lXVZl3lIBKLaOAKbQKcwZYengjfLIDRoMleGwrDJVAUQ+eou3WlXY
FvLNyigtvdFsL99zS6yMQAPUgQU5Di5uzrZXV9WQF48d6SVk/VC90G4KM5AK
v0K/cnmR65AaXM1qZZEtTQD5kIQUbQFYld3ifwA1Xid+vq5EPMvBjC4NDi4G
bCQtqRDfVz1B1pD/oZyK7YyDJ7jlqzO3o+Bxd6mAnoxnydpn+taq9T8EPnK1
IypYSTUoPueVRlXC6PG4hdMH7IV01JQJ9lWERvsdBoBbsnTd11RXO4sTfS6l
vCL2lRDOb6rjCTm7DEc3xDdfARtzwC1OD8i6ZtTqCjx1X+Sm2jRMioHbF4yv
7JeVEp3OotyPm0XAhK6XASkf2cFulZAcxkm/LRl1TZGr7c2kuWvSHX521j+z
cOzt59WdQjRwEgLcfPWlsksd++I3pD0u+jRvvi1SUjG1t/kWvBJSQmw5RynV
OQFtF3ayEQNzCvmBR+fF1jtgzcZrtcwZDrvb02oOMKijasDGXAEeuVAywo+b
aRkq1tvPMBDeUy/aNANivMjOxpjUpa2Y0nsqE4vq26eGHu5c9dx+K7ikh8sy
jlcQ8q51tnqELIydSgvGrJNwyZx/vXcusSegQHiAZslAMpqjtIet1NoSxu7F
nLyKdu9zMDF41mTfGoEJD3/5v6OjwU1tOLDESuGW6uLaxNAWn2tibrz/DA4/
jckvUmyuCNSFys2tyQi8WWStiTxupYqWijNKQopl56PfFiOMafH5loQDPWQE
kfNQPSXTsW/Ua73lcbb/3E5Sm4lnbRH+6PCP4PGc8wXldt9jDy/m3o+Ubqc/
7xNqORqabHXjnbQHKP8rSZzAxjCuGgBR7pudAbkyth+qfovp5TybsiVXE9dR
CXxPyqsXqM5JkfKAPSXVcsBjfDFW1wooN5QGGEhBIth2WlCCWf0rAlMjns58
JCfJJAHW20FdPcgXc4wivUh582eK3bjWQzvhu6/BI3GO6DLXIbWx/MJffPCd
SETQm8+FVwwveVP+NanK0BZj4KC4p0dXX1mBt8G8IgcsIedb6+cRjRvnA+xS
zZvs8/xUrQ3e0TAhB7Z2nBZfQgvWLK6v2HMG6lvdUoTFfjiQ0yRU54WQlsgp
XAunge1wnCZ1UXhJacK91tfIhVR3WKHslY8KwPRa3iZyOiOJGhWcAJCJJ1Jp
oe/mPm94pecN6wtGML+yHEikL0NZ2txbAbuyIiepfVw48C7hUDhD9L5KOf4n
m5HNUJa4SboLiupiWCft4uBc91pIYC0F1qzUbU5ZzEyxWlTcFUoAYFSCoQ0Q
QytwS+RHgzQju6wi/use1Ac9YWkiUnC7J9LefYinNR9bO6zsNAHFpqY3eEQv
n56Ki7V0y/q3sBEu+5TaamItihGjgr6xoDHVzd1q52tAvdUYk/kRqH0CuDPm
lZSsIGKlUapPRMofI4vFevv+anShBWI+ODxRyb6sJPnhiH6ZxbcO1SSHUiNI
RK3xAfzQXjRh8XkHm0gHwxfdlbYki+v6E78SMXC8BiaLj8X6vUJQUYEQ2Zxj
uaTFXZDYkVIRVvhqgrZiepqWhWXNDGb59TyNRRSJqpdDRzsWAQZzVMlRzZYw
RlgL0b3MXJ63rjSchQLdx80RfhRkETSpsVR8V0pfOpAJjdD2YAVMEVzJVLMt
Ynjqcd2k6+9SlU8wIt2fG8MNZwtPZCk1QBffoPjMHYa4pwOWYzo2uMw972+Z
l1Ktt8jmxA2lTbgbPNbaVfbVHgE8ZtRGmRXj/r5XjMHYdIaonGwRodwvsK8d
YyeTpNa7k4x0BVWYHe/GtpDpU+0g8kPgLt7e9VO88aPgdZOzqYQ+LQnbxkjF
qv7/Uqc6zWNSsGnyLmUPlzs+VuTT+ZaLH+6BZUoiArpukpjzlkSnOkomeTiE
12B2ka6pfuPPtHksUYMhwx/mFJEzMVOIRTp3BKqM35wtUL+AgBJSSjSwJxWr
7k7ZEO1cu8LQEobMj5XYxKC2w0QhHeyFglY/B/PJdNfCk5qBzh+PZHldRwHQ
T2gCNwhFOvh+YskQ6Ky0LvwiQWDq90PecTaXz9+SAkEdBWXZlfuXs1zYKKsO
bzqoU+GwsW336aWiwuIwXZc5Pi+3N0lpovS9nkTPfGCKzhnHnAbjqqiPiFLj
SDjl63EzXEdEKvv653gERlNCfEs3aK1I5OGD1zBMb37g2KA+KhFtb4pmxpiZ
JzTufX2/L8MBtd6Ns8QRffxDMcuUi+CrovXDvI+anCUzcALWOTQZEoUNhQ8E
arZgKQXYSe38xreMkSJqEO/5EC1n8LKlckDcKo2GOmj7koLnXLS495AgJZWv
+5ZKZkYHm0c99lrnqJw7VEKayxH57ErOY4TSWQV3zW2J7Qm6rI8/AmRAVIXE
JkY5hBAhKH7ib4yJnfODxkrVqkF43O3ijWlSV4RHGNP9FBAgpCegxAWCqP2j
NKsjNaLNpBOpkAVoSVKtqr6CgRQUrh86G5obfiXWT6YWGLy4EAFmjR8FIW/3
flTYbz6NarCL+0jQY/rzh9L0vLDuNERyCwt0kh0Ml1Tf+w+jHeBqMVemb7YK
tKI4nhOfxkdWQqW9bloNt/04y3JTPwWqbvEzpG4szCscxhK+rPf17Dfi/d47
oLV531d9wGilE21QA88GkyMWl2u406k/6wdYALfB03vA4D2ZYXaa5t+J/NVo
ggcF9fCTZ8gTa83KXw60B2k+l0tjPb9/RntqjQ3jnPIVDguULVNqNBMi3Xoo
mzu/STsJggaZAWywIdmoh8zyluVLXLWwwhatdqDU2QC2csZ5XYTcYJ9G8abW
iDaj+JJX1QXKQYKRCOFqwgimkqhSb4U+qShZ6Dsy0AM3UkbCptL7w3bu9epA
Ys+wc+9cMgPhdeRsEOAe7NmR84j/sJoiwzthYCKbHrlIkOmNaWCPKt8X2Z5u
g7kaAG2AyStHees6/6LHYOCMWx2zUSkGae+I4VXtrL07+88NwngsyknItZbS
lPW315cnURH48wU7ZgnnzOgcpfkuc4qjRDLOc0Wtc1IYJS5AHx9czftoguB0
a7jHzfMMXyRd/1Txqp2Nvbcsc4mxSQsl9Z87Q9AO/XdPmJ86jATJDz2OilG+
IX2D233B8HO4Zkb7ruD4pYI1tUzLyAh6s7BpH+/QBNJsoektcakhMf9qlX+0
E16Mn2BKENqEXZ3OLRxjfkYu1vgF/CYydWvA66Ws+TByf4Ca2AetCU1tnMeU
qr9nysuEd4XqBA9uHOUB1LCWxmXBAr6ORsT3n58JMmjhHnXNLzcr4l5bImRO
F4jfXOR1Dcq8k1nDlSK7AtD0DwhUkz7F0SJqsWgscB789s8U/VIgHsdYUbDg
in+Ie5kRTInciADdqArBCBLjqLKaoIbFzE0ZdxD9TDPNye3tVMkaMAfyEQod
86toyC0NYeOXnJFoqHZVJcC2RqdUs6PtEBsA9h4z9lOssUaqUJjJUKv3i2ee
DxGYDY8ivYHr9jkOZDDFD50THKm3fiXHRoUHm9mMAKwQb3Q8rImrxBGclh5V
BZfP6tKNP/Q0MasCH1QONvjjxG4IiuXW1FgXjscfwpwbgXsZ6HJodIM2B20J
qYt3nH+MLqmZeq8VEJF517WY/yXPmKPm1SSD5dEkMuqfg7O7GS0yx6uwpkCX
DJI3tUxLLqzj9LZ4vjK1XhNq5Wrdcxag35s8KGakVBsF5egeRyzZ2Fi32R8y
Wr3TJ0FKlbVNqDVTbChIoRtczEqqYcuXSVDSx8t6fc2Y3qkW1jpPZvhPi/4N
p7HfVoR9V6ppkACu7LVaGc6i74JzIbLpylAoaKUX2g8PuIESgS8keuYVLYbn
Gy5myLKDJRmAcdpCGCrGUAbRHwa6zuYMvrBGNRImZEIpWEZPylmXc8ot5fcm
rvY4x4txiWY+f1nZGWWy7O++TRJZZsodvGOmOMdsTg8c8fjlfXhaQI5BqF8R
ens2bb9c4vKOJvvKq5k7kUYhsgspoohUy6trwi1qMdVltkei3Yq3u3T9Menp
B8JpxgxZXJiXwkYwDRb+BrdmnO2dIfn/CPTjyKzYQ/cPXAt7k7xT9mXcN4l6
WEY3ii016INepugZLwCCOmnFrSFNfYWAJOeImNS7ceUQBkAOQZrFCRymE/0j
TrL8Iu71eQB8r9qN/BBzxd/A78HbAD51wcXCRliSB14Ufpu4v2IqCuPLUz9P
Lbmh4sj7A2rapNBMSb783m/7qf4bzpwFPUsCxGAZ2wFbOdq8RJQTzOdQynVl
u/5SwOhjIPUkDxMZesfYmr+pudwNFsqA9hvZ9xQjrSgmLEAc8DsZnDJdbrPX
jSXUXV6SIMp6uilWKZ4Bve2sF7AlzaEWaLVw1PXTwyih8ThAXdz7m/X2Vr/W
rHrTGvu0ZmzDOclfYh2wl0o8Yeauc2nqCUauVxRD1pyLSRSw6yxUtdgz5Ay6
Py4SHsPVnPZYMPhqT1md9f3x1c89O/ku5ur14naE4oPUuXYXmbirytKP+XRQ
pJ4KRATyatQw3DSQU1bQv5lyhlF57jeMjeR9tAdmn/edvFkgn3o6YvIv9Nlf
7FFVzYCriwPPt678ms1DErjgvYCE3Kxx42u8shB/cCBn4jF2R6h8wjxwOSds
lVFHxM86lDxuX3qtZQVc3dDPRZCE+kX+C/wYm6rD+D0m8m0RW6I9srs9H0rp
UFtZlde6RYwnvSidC1dymkfk107SGxRL/hFguII+rPd9IanSL5JAk36QiJpK
in5p1nU5WgNBcVJvpYQ583Am0S3c38q4c3ahyLI8sla03ouJofOWUZ+sHhBJ
pKHOnnAfZL7yXyq0xR+c2nOq5CEkKiBrrQVrrruWvudbt3hcZM6xHZG3g3W6
6lFzGdyFoyyzE1JiMebXt+faCr9pS9pIHM4f7AgRiZNOpHpRiyIAvvDbOKYs
jBw2c24rq4g5rqC6uhSJfcwRscqjN4fRTUGgpxv/pKryQSY2MeUHzHeBF8rs
d5C8jafIqhOMK+uXKb9FCm0piM0mwNGPyIHacPZh7NErZSpxvdtbX2C60eau
V4XE2ksvkm/WkXyitixGnIql3+IlAyr9PoSMvEOUN4zuSWCL/oLcOvfmwiZa
JGrhaDAKa7HIcmknlZ9M8L3H12k2T8Rn6lX9vRrQLFPvSGXuTRXDu1Gb+VYz
NE7ZLlITllet9e5LILIdTpTjACKE7tJqPWLwVIkE38xR9wndGHHQQTuxUwEt
vqSsrg1JkZMQNE+Y0pEbYbB/ITMM+xmLZPQ01pahQdOzyCoRDAg5KcJ1Ihch
TwlQQIosUc6BRZP/tEhiQKETBN3+rr90l4bjaGgaUZaR756lWRUg10O14emU
yH4hQOwXJIiO5I46El3UDV8v4BusyvmoBoLflJJlLW4olntNcPhvhAppdBkE
ZHkFLGjh4u/MBQFJqtzHxz9mwBrrykwWnG0xEP9lcJ8SZM4KvfjTaMUoDo3Q
P909P0YMGQISo0WZin/iYv2QW9fXMvRDvv4fecHNCHPePbdFvsHYrEETGWFk
gt4IobsMidKmZjlwLaOepoUOIgQRJfZCQ7BOvQ168LDNDpfEoqDH9/zoiW1e
kMJGbuw5dU9nuaCQKH06wi9AudRHo6feBnbT/JvDGEXwUBqFCaTCsYmN94oo
YiRCxrcywCseIYJW/8x1puGdFZUVRf7lqFLaZrT+rjdOYml5rnBNKmGciPDH
XxhiQSdBMihXCRJFZ1LH4+L8O7gPJeSc2+I4UPdCRyO9G4mmxkvxNeKf6JY9
zL5pir9iZnhXbUDR2No9IXpMPYNKYj0a6XqXGwF6KLOfYGS0A3+baRx9p8nh
ALdB3PDRC0wV7WiXH2hdHN9Q3VCh2BsQ2QRKF1+Ljt4LM1ImBFbMjLnKhvYG
qysUOSJZT99HASg/5UKJgiKBVOYH2E6UetGNYxsSCYNu0BbAAlsd7SfrVeQm
iHEaaTtoZcZg5Cnbx9gtTUyEJyFMl1gZ1/XGqydXvqne6hV/LrLrly1AdWRi
MTYL5JqgkU259UhR/JYxYd8xe+h7mIE9b69guzgej7+FIIcIlNzigkDplVVC
jO3dzsndq9qBJ4Wd44wJci/huuQeIGb8fkLC1SxEa+cXQMUxOHoj/F+I6HTs
YBq9Sulmw5bnbQheGGUCgODK/OCdHkMb0KmNxvHt6YM40JlA/roVjBoSCWgu
zLs51SSM0zHUtQpuwCDT6/sF3wNaXhY7vRAsK1ofPVFD5d4Wj86+QJ+46n/T
lt189q7FXDFlga/3PqRceF+66NeIkFEgAFZQv7Pn9AYUtKhKSgVY1otIKMp4
/6Li5VIQnQyv9Brsir6L6W5mgNlDtYnbZqPaag0icLEdKHFOWb2HAI58sZhF
HAMXH+Gmxz4QHkbrwSzCDlsLARRCUEy+T4KBzQoTPznbd958fp7C1ULv0dJw
m0bbHHCkmxr4AhTGcDs6yNbYp6DSawMzMcifWXynOQ7rVVwiEtULL2plMDwr
Ndgd9ingtgg7LSxwIQBmpPAZLVXKx1p27shcaUz+niW+S9E6Fo2rpPquaw0Z
PIqiraTLhUllSNjqxobojjwdNw26ne2AU+5bER3QzGpIpo2U+LNwv2xyiLH4
0rYnG4c7UBRvsKE12gVABNCSDgXMYmW1GXWKz7TvDNIYfU9m7ge3ouHaGhDd
zYle62vlnxVUKmZQdEVNmbLzAABHdaPE+l96/3jXaaZshIphr4qm2zmK3gmE
Gcf+/5IDOla9mQIt2nxSgp6LfG0AC7gpb2QCamRF1RF8wY73UnDiNcQVJZ8C
M2IiyM3UaxLw9YZ9qj7XSX90UMOkAjRt9CtZmpqp1H4v2e9ZRVVGMj3/ybmb
mC6+K28z28Qx1E3oO2hmalSapCUrUvvRCAec5g6EeEXjogGP8HyEV+m07h11
WRu/X6IOq/u5JYgcydx9iWovlezNnIaRtK/N60pp0bvoVQMqUBkxTuB8uLwd
c/VqsG4svAE+bHpaWGwUqwQOJ7pqBQAcMEyCsIDQey6IIqMSinMLTPxsik0H
34STYg3XZpm+N++mLAijek4vVmJWrc4JKBdILGGvsMpFvtz36r5+m42ZhRnv
jKZK9pysVaJnjJk0bdZLNksFjT4a+qgACk6/MQI74SnKdtMiF4Ee+csAv1Bo
dIUb5SWJN4h/EvctdmADYPlRGrwZ9eE9obfssPwYspYj24UXviTRcUoTc1rQ
wSSGPhOq/rVQxKPrP3JJ9K9Th9bncnlhsZmviTVsMJPDsAAFzyWlOfta/5sX
syUMo9NYvbDccS7XvBW2BRCUNw646VOb/GBSydPdcy/in5mWyuUWHC7NAgiq
jtGcqkDQkuI0WcWVFoBOnOfmDNgHO73KB4j97HmY2GeLFV+CDR3Hvp1egTGq
gwHbLQPNTwySNqJwjehXITC83BLPPpxpZJU0rMZJWoAHx5QkbhM3f3kEt7AL
KPkounLHOGUWEwzX4t0ZXyhIZNGXQ9WA3us5U2G8Dy65RKmdGVffx+nGI3lV
QHj0y+9HPPCsqUAD3u+dDQ56aukG4faNI8WAc8ATgzpj2/4wU/cFxUXgKwVh
RVqaHWhQ0dFyOIsAPPFvgEyQLu57xR+vztnXOQjDFB50asfWBo5HTxETbyhU
kZpebRmxjLklFsjNR73tQvVBzwXR/C9evCRuAvGGacmUJfwddp6utT1hxWAt
WS5nP30sFcl3BTLRtemRxhAsMVp5UnHoLyaHm66Kee/TKvKWKFl/YOB6U1qu
qOKAUA/W93mDPnrlcc7EG7rtjbYjjaWoJFtZW4M6xhk/RMwgHl0fCmMsxpuJ
feuXJBmh0rH0kRZNEIVaU7QvMp//0SX4wUDMmiIB00VU+iV3VdG41rTJvco7
acZcIZooR3LKTVlJ+2jrXCY6X4uD/PJ9T/KgXbC4lUsoo7sL08QC1kbo6bXc
zhXNU5It9ySq5ptP66rlH4JIrNQQcmNAK7lGU26VJJjtBTlavTzVnXz+nSfi
G4zBDIw0yFSeHU29joQdESUTou0SE6mo1bWSeFPjuXUPMfE1Ec0JwTqZQ9RV
YWQDPesTd9X+pZQDaDUaKtDsE5epSJQld+A9XjLvuV3mJwulA4vHgjgNHCyc
3NBbfFhMee+cKjdz9fZjH3+ddgxlccenkOFcNBtBEShcTQsO6uB9DDpMYcf0
1yfdjCD070rmqfkGZ4FDd7N52uaBuVlHUryQ1lHubXFcQae5K8Ff8gt6TzTD
y+fJD40kUbYN5cr9Vi5IY47Euy6E4c4wR65KsOzDEkv2Xx9LEFJ6nx6SfNoK
ZfxbNX1S1T/MoQz99Bv3S5RKRdS4P1xAFHyriQLDi1PoNnXb6lrOjPPkzQbB
6y3YSS7qELhR+k7+tWZZHcjpCbFoKHWRQpwtpYhbrlTHvR9rLgeqURZrae4S
ay7hWJ++m/rf8XDJwdG+1MyD20+5c4ymqhsuRHoD9WT0cLh/+AUAL/lqnCDO
NbXqdiB/T+jNam5UuSDbPo517SeL8+PU3cvZDHcobEskuzdvQmCufMus0WCb
kdkWVk4HoxJ3uYR7uuOU4LsPBiWmWG6GI3kX/Yn4wfLE7mZqoeMy2YoMB/xK
N3lw6TE1pmB9hgbPqO6hz0K41YWeeFIQzXsE0J5w9fWIDOHW4BUIUwf9/kG8
qo1Rh7yTC1Lf9EqICfOQ85l9lswRYNryBm69BItYk4T6A64RN491XVhb6O+C
3BrPBILaTOI8SUTJrRoBZZOtRiJxYTAxw9tox8xlVt9O9dcTdyzGobfo0fMl
kc5hO48GcDyuxD8nQOXTuf1a4Z1kzODlrt5ElHRvt5BkwjLuRJoYR7nJT4h4
emms7ZkMQ1P7CYQyE470HUO3vuZ1DMd/oIRvxpwMXWUU5x8q6VtumtaKHuNq
GsTPP4BycPWjsE14Q3wsfspPGmLf1vcbH5X2FN2T66YtxCKF1edxRWxccdXH
ugtGOcbCejRR89RnNz238h0b4+BSYwQn1QnMu8HVRGn5tMR1m3FUve+iSPvg
RyEnACNa3m8DEJOR+GJfb6PUfX8VnyQWRvh3vfTzi2asCxSa6Q0XvV96YZ4Y
SEKSNGqkz+9HLm8CP7BNUzOIcOJ0Pg7+u51LhBumaNFwJCMCXeC4UvFJVXq7
V5IXKM+y5OUvXteorFvK90/fb+Yb+QbM3zMse2vBS2+r5VeEcHGHTxzLJHje
yaii671+F1p6gH86M6kLrpd6eonWRAWeLxYAodA87W1iz9pVNBHnq0CgeGOT
CaWPnfMpCIoJGAYRqeBo6QxkUclaRx4q2tSD/KbtsgC8aDR4kdUKcTCu8Ta7
apW3li9JWZN7ipyHlwIdllNjuOkgKd0gD9dr+MWfAy+aL5mm2Tr5z/xOnpQF
yTdXYdjv3cxWWPntrg3f8g3hlpPkgbt+hB1SJc765WXMQUx2UmY20y7R7uQE
1aoJYclGrDd99FmV9/D65jiGUbztt7gejFSlRGt1ahMWa4+Okxaj0KnxT8WX
gWd8SmMwdUD6Xj0Ak+YMSwh8aXd+BkHeRCeR83CuvvcKDv2PfJyz3fsg68gy
rAhwexbu6F6m5KxnQA8xOjNfkK2TwGswWyJ9XQi4y6NCRpd5oIP4ivXalWeS
yOWtdmIk4tigyjhP/AYBVfcGKiTt6421xVHfB3qF4wUgfcXvL9EcG6AfK6Qu
uFD5M88/5lcohfWn3CWGPZ6HXbhW0A1T7QLOQVUxuQz3VoatBqvf3I1g1QUX
tAel9Yh16Q9j1ArbfR15Wyv5nFib95/6WxvwVex5CVWvBiw5jm4KYokZB9hz
Zexx4jOfj3TptsDSJBk9aHdttoLvEjIaRkhq9hNAIXFNTrEC+utnqXa9OA4b
WYRz+OwXp8R0z3+Kr/4RguI83HS5KA41+sbke/M3YqyWCqKhEC8WHHuXdkx0
CGakWkWQBBRJ8fgCqh8h7CYZxZaprruUje8KFtXTj8sPHRzYJlRuU0DBY7ky
jOIZZ3/5+Mme4Ng3z16bhtR+IkUBpJLTL2I7CKlISf7j1LqS48QOs1VYmdBY
UtGDAU5RJHlcTzmHY2cJcVFJhQzaPMi35titqr3WD32eTBvNyq7WjvDx8HYT
yUHFKKN1vwmQrzahP8GAlpjck70BwRtWCrkHk3CeYzRC9YoWv96hBluhf2uE
B9zC7GvjOCjdNXTMshC7FWpsFfD/dQ9usZFYGOxmB9ZYLUJIn2fY7AKiXSj/
kDW3fEOUagB8wd3Ok0CVykTjtRhTwlPiaJGHVPCIpFUeD/t2EmLspGjA7c4s
UBfCWp90GvfOrICRdO8xr2NVrhU7ztSPgRZZZ0KelKB2a9jTN68pBBYKZPYV
a2UdFPlAJPQQFSXDkuiqmumlUUpx9+W353c8ZgoOrgwX6m0Xq8rOn/byBeTM
XN/47SFv1tfkKS6DFrCcV2yWxlU2covuwgt32QVEjTQ6mAkjhMK1vWHxrFgG
HNgp1+EYGQrfyUPgSPuLLtBzXPxqW69y8k/8Vf2qQzI2BHwl0oebc7zz29vo
soqVIStFR+DHT7SJoUhOi6NnnNx2dmkj/Fc/2RTpM1pmCQRuqN9D2kfJrbUL
mgD6xScLMnrt06CfVMRCzQwVWlZGUX13MEAh5H2zpnirg8/jp6t8gBL42m4D
SOFefC4pQiJlGIF2dJRpL02iSZKPC5K1s7YA57Mmqg1JPgyF0Ku4xjDE8d4X
JQxkmNLpVYam7qtWTnk1O6q3hF7UjyJwNPmC0UeXmBsnAYd8GhxG+bostxNE
I15dR7DRkHbetsRTL/htUlL/qeH+6+vbaRUJDndbNfuPwAdT8ham0hu8hkCx
aRLOeudX7D+1ZmwlM+B+tBkoHTnBtnr8c7B9Cy3n3erLmUSdgtF2abWlf3dA
43tk6uT08wKOZrodx0+TqR8qTXPfcuNcIhE8zddoJ7BQSdU+L6jUX1hVd99T
blOd83c9jlVffzQOBGwXwcMfeqQGut5rH4BggDvOafNeYDis9GJfMksxt0Mc
eSJOc8TVnDlUGTZqVtwJqLmSeA7RkFMhaDCgGadL+DdYHr6Pmbpx0AASm/nu
RNgt0bHjmG4iSQk7CM3g2V4jRqJ0fogadahnWM0gUvTnob8afw3KtrNxiTai
eKjN5mppvB3f7gl/A7R0Cq9HU6BdScp515sGiOEsOKuJHOqeGGZSsLJEBSTm
Oo6Kt1kGxkHdphaie29WDub2OFtAJqvawRECWSa9iArUpKwy+BFp7HkXvfNk
+yxBcTVDjY9YvEeA8xfbxZfgHfTQBJHzOazFdeBEh7cd+AsL2UoM0ETC6gBl
lpNdkbw8ga4zc09So6oaE2PuG6cjZRxHhVsfOUfoHbCQIU3wUXrRc2Fwj5qb
fvOzSYuGbESjQ+pImFNvmVruWNgdV1wWxRlS0ZzY4OQcr7LsQS9eF3wcsJdp
U7v/ENF1shk6V2H5LCx9rHIAhdFoOGIlNhV/awD9fA4uPGwQ7J07r/eTWyLT
oTNPhHWea9bntnljryg3BeQIwVAwhUI0seMRx1fmdG0dncQpBdIDtVAZ9Tk8
f1yd0SjGLA9fXgmQrB4z4q6GDZLl2deVNcPt3R7r64aa2pfxDxske+kgztp0
fWvAbkztQpwEDyYtvmh0QHLUMTS58ruSXB9EQ1UiwWGbNvlBNepJZoPlfq4q
4r0ClUt91nUqyuJES8ZrOm8FwagmZ/NwY9kn49a1+3R3nR+Bc5vB7lb3eSak
KFK1xCCtlWMp+SfVbNxthnzVenyuL2dS/djGsPImBs2rDx5elTuXa6mxsIBz
LLU0woAqXAoQSweskwcRrZGDVJFgVHe4FDWZzyiLASSAeU946Rk6vIJkUZYl
XzVSIEXFHaAKgMGI+7ryHJxtgSivbaZ8y6AOFhXeBdg4rNXNlnGFSYANSm+5
ZkhhpdVQj79Hh95/S3WpmRBf6Q5l692AvD5uHA0jOau0sNiQkBnOzxXdcwuU
ZIPIJXQy1ljohYA5Z4FEVbyC7KJBbSviWeRNNeqVnwEG4I3+HeGwu8hI7wB8
n+14BzlfTvSzLQ5g9ufWwNldEtsue6qFQ0gRp2poXLrlTIxVhNatcQO9Ttdp
luEHPys7RHWavJTloqFUUwpLnB97W9Io9Ng76/ZwY9lf90M212KT3i6zwisD
JlVQe/RyXigZzIDqrET43YkMSixPyNfhTV9X4Od4aXKV8Cn7UrpvEQhIvXrW
L23j8+rKRZzAU5RE3i74T2GJnXPLOX8AAfph4boTVrqzUwsyU8QL9mPBw7MW
cvCAgotu6+HjR4tjKRRp83YGRCdV4EjkGLlOjAUa3S+jH/pjhUOZTt1zAFyA
PtINw8tepD8n38slQPt7CLpLu50LHjKl2ZuxFwb658V9qOZYgFoQ6B4QNaWo
q5tj7orHaHwXB5mdrkjD7QCLoXO/fqb9kH0mgNDfPK1NYFMXrdoRq0DEq29q
YcMVm2LMYsv5M0t+CFsaoRQhMxIIBBeLmZTI7jdxiASfcVnZvu5XuH3JGHMb
wwGYwN5IRMnA6s6cDLWKDWysQq4WmuhBupL36SxZb8ZxEuZfZ4qI32L8t62e
GR0ZDQXNJxNaHp2umwD4SbY4rSbOf4xzx0MPi87/MtLQ1go4tLx+3S/JlpiE
FQRIKTOoVhbLfZXSUriQQ50iHMcmKA93LXtKnvQZGlNR++mp6COPyw7KGS8L
iRaIBbKDTHD+dhiGov1j79VgMwRvYeVXSGY9RKPmR104kQvsZrtByoWOSSKw
hm2higFzPhjykbBEuhor+BHR8x0OgSJylJQ7qC60X/eR37URSgzTcGjnpG57
YZmqs8Ai2/Mllw47mlDZvBbGwj4gPdolU6zDkCpaPbIsHv2wO3M6xgBn7DK+
WtFEIT72i7x30kbi2QU9pK5L5rguj323g+sq6YO6aSmXBvHZ/IaCHE/BQxbw
sYXQ47yAL+zpRs+uJu1YPCbdsl15Syt09g34zLuRgrFtgQ0FCyE55gYnVY66
MJPUsr8ulthFHR2pULQTQD3UGX3RwTX5MiZ5wmWp6rbxDe99dZhcS+pQsihB
ZZKL3bVb0bpVoK/3YpSeaao+liHQXl7pwrQtwNCxJqrLIFwToomaRr1NbNzs
XwDr2sdUjdUrgkaTGkJew52xFHtRIIDEgG5EPcyvJDteKAT3yzz0H4cfcjL2
Lv3QtPrWw3yProAJaKKxz4jBOF0NWNobIBw6qeRBiWMAcVOZ4u/fMd0Lr8NB
g3QRDkQeIu5K9bqOLNRgsllzG5Iqte+9RPjei+hJJ1iCWPgPA4a4BaDGFp0T
Rt8eYpL1tCrWhHKVisodt22/71hyaj/ERe/72C8e7sXIc8l7pso53SNBrH4b
FDQE5yUUmEoIzAAp2/J5RXhPU6IO9neQ8HyMJ28Wjm5LlB625gx0vO879inP
TuzLHNp7u33XDO+UYQm1hXSK4vDnfUJd1Wn1QQFDWWhIYUlBEJSQAhJ5UZeP
mXgQzqZ4N0lnpE0I8jkVdG+SGqXWRyAcQI/TLms45ey/LusICoAzbtPUaNlo
F1J8PXurHktSPXkeHdTHq5BadgW0l0qy9lKtBwmOMq4RrQZHUyqhfMlTtBsz
LfhSOu89bxL2YjgdK/qYX5NBMPsCOpgFIct1/bOtF1JqJ0q5WvVN9AqJ3jRn
xaVsugfIK4GJl4g77SCsBcz75sSfolp0i5cC+8lOdJ8Y6FoMVVMYTn5k6qBq
SEKiRC23qVxz8le6xjx4kRT4BYH0iuaLJzBp9LtrrGF2sofd1cY68yLUokc6
2SCRBxpv1QVgHWX5WxwNCF7lz5q3Y1b8Zc6K+zmfNcLFqu3w6asv279zKJKv
X7/EeK9n4SKFEa2z0p1DbjmuCFeB8OYpwZe/hlO2zMFd2B+68/4sCuIsD4V1
Rt7gf/Y70m1AHfAg5TKhtWA/pFESUvLbSmjarRMpR2gA8zZ/7pauui87ACg3
yNU3AJyqyruXliEcobhRORVsBMvwLNiCZZ3DOIJuckpZLeK3+3dIcIgDPsET
IbPtqQjCU54G+Dj18ab7MtcncrY9CpILYLXlhhkpLSuKioKXc6+YanmD6+Aa
rPTy3fjfdon63Ivz4HtUAIrOflhxA750LH3TpiqmNiWXJKUwdJ6C4KBfEFTh
sZ+wxC3YkB2d96sG93HTv+xZA3dOCerPqeZqzAoSZZ8wCWdIscDRsaLj1lc1
68/nyHKLAo0QZeGU1lXvD37lmqj2uTy2UsHyT9A6QXJQwl4QRtvtgdLrxZy7
fPZdDfuVZZHF0mIt5l4eU/ElHQd5b5S3Nz+HW7deg2uxLlMHdIyn+e5ild5d
Exu2tFqtpkVPaxSMkvZrO0iiubhYy0xNc+lNYCStEfqgIjYRu9Ijt7qKX6OX
+X9JjkSEC/zOpQPU30CvdRNoUuI/fdBYxHBbxnuC0U/x9DKHGotf9y7e76PQ
gEFYcxz6jciWEOO+EbYr5FmZXjB9g6HFzHMwop7Gd6KgG3uN+uCjNHKpF3MA
9OH/O+U4LsdJD/pqvW21F5SBBVWFsIihtWqM9ars4aPZkR6Vie9jo2lGFBtt
EfeVG6VhEZL49bH6cllJ0dnSRIunbvq7YJhc+v3MY8wloKpQ4PZT1Q7aMYgN
eFZ/vYxkHoim4EhXPNs8mgmLmpK2LCF36s587NsHSmesbJyG4yEptfn1fZN5
Nm0P6HvkN4jXnaafsFaeEreHK/rs0zyDA1vWLr5U27gbyVA4p9IPs5m8tNVZ
083vV5B8FzVNJQIpS9SOVVg+S1APPW0YNgJ733yyvqhNJOLyIZCtlVxmqHwD
WOLrJKAJY2VAYmlIsP+haGG8KWppmSSyJl/jNHS1vEk+xvzTpwzkMBq4kC0j
uCFTOnZMSKq3KKH+JXKFfqfznT8pE9m6VZNRiA/YM/uGeo/07Zz1UFD7+KAn
6Gu1wgdqfmyfKN8OLYPbPUqP/BZ2TsuqUnEcrG4mCys8dW7x0RvvLzfTlY6o
FRkZ4SJ/57Ut96W/gEcXRIiLRg9Ac9ktt8KfQyINzWyQ0xWP3bsR9Y9TeU8x
SNfTwf51OTeLqu42w8P6wTSa3XjT0uB9r1UhtONU5jmpYwhzzuyuqZAmKWRP
yeQXG5luvtdymrKbBW9SuLdt7WoyLz3/hM+7bPu0MjEOvOdJG7e9j0OxNdIm
PWk+JoCJ59HCqfGfBvDZzs7522aG6cY/rf9OQ1muc0ecF/lGW+s5utWmXCRA
D8+VAhcBUsau5GpXPhDGGyJo67ecNnaM1wlf+cYXHOZS2dgCj2zhIqkyeMLP
M+8Ss5eLhbbVf7vzkqNEwwilETEbiMOaqSJm1sse+0tsmNSVDlgSTMw3+mTG
QwMMdFIik/jLrgx4IFx8KQ92v/nXWJKwJVK6anliKhvBeOH7CtH9/ZoA4A0r
PVQK8aOwkOl3KVgAO9OKmp9eAm3naC0YyFKwyNqdqjFIEMnf9jlbiGBXQYGW
AnQpMma9Ikxrg7BB5T5lFWJavvxu72B0UhKs07aqpd2dPvUqJJSMsCatLlsj
sL7BrLxsimHwjWMr7IzhQR7+SU8OsM6IqX9OWSb1gQ8n61egRu8FZ5pnTPTW
Kx+ATnUt7U9QB5oD0E1zMREMbYDZSUFqngDkCV/CCPTIsVCp2HxpEd14AgM/
1JMI60GVMAmKUhn2wJwMA06FpavNGoVyWWmNmDySsERG4mu22hAZf6jbflg9
zZ6QMnad7uZID9atwkLKMXkAAc8XpBqqgj1sb0ecMRR/ho24q+P6oVQuPOuK
/OIaGUASd/La8EXOTNrs2DlqVqsrto4mUURgZ70Q4Qz0GPN7vrFvsOn7ZwHi
V3/bagW6AMV07T7WvoSVF0/yEqt9H6YWC30MFFFRKwQ1WEaRcRjfp/Tgb1Wi
XF/iqxRlGeKohCLi2HyZquWXREbf/mVtsjdrVJJLpdi1rtw74xHndgOgNwJD
tltk4+WbjRDScplj/KFktMl3SyN5tC1lSmRvpmSMvWgPTyFFoe1Abep/GSYP
YeosUWX/+vg/lMellk/K8Q3dCiZDz+sOB9AN+MwXtx9tALu+6Zn+KAgwE8Co
HhO+3cYW5TnsLoATtUObzxrSGs0/aQa1W+wRsNPT6SVnevBz7B2umMBGFiA6
JDXrbniHiK0JuF5PQI0VS6+fAx1E/wOcM9dKYm1GAwpZplUIDz/lFENKZhyn
GO60upGMkK8Md/IjQTLPpv5lb1nIsayspuRlZ1BfCAbMY5cUWarzQlzFfqS/
DjrwLVHOn1+MkRhsGlnIRCfKB8JERx1QUrhzNTtGqBk6bSl+N6GnzkzOoQez
36RTdO5ncPAparPuacHbvKJAcNxzmaxbv4h66iY73bjd/A70ugo1+Im3s076
kv98XEK6iThoLtQZ9/w4e9KtggZZrVqsX+j4mz5sJBk7jaOWJcri25U1ZVZ8
163NS8ZXyVKvYF8rNKUoVD/yJsOSbSvkTzQDkYoOpjdDADpB0Hxx/PRzcWJG
ohxbST3kKstpFo3Ok4QgYEaFfrXf11Jqu2FPAvDpuO/t0aFSQ+7EyOuMbd8P
kNEdQ9Inp3BsSqWwSzjbQgHFOosqYi9HPJBgSzGxRKozqU9rP5iB+PhDS8aG
+NXmuV3MtD1P+GMO/9fuIvCGzDza06McM1g8da2v8qjsSkteHwGgjDE+VDwx
mVHlrnpktDO7hiZS6D3utCbd2gmNTzZSq3EQMCXU9sf0r9FUb00xY0/ebNzx
Dk5SvsBh+EZ8qYDhjmV87+M4Jf+HabxpmVNe2j1H99t3j5+IhCLZXYGvlBL1
xl35/ytkgyWhIm/aDZHp9xqtUkRTwKwlhVyv5erfkZC8NpNzQKUTYoQsThSF
Kj8GEXnbhf4SaxJaf/VO+Td20xrY3sjoaZ0IQ3jyG1C8gCbQU35mCvbWKNWi
EzUZQp2+wOrMtJWUlvTy7a+EF3wKni+fiztLnHGoyVaO8ePDdNpbFWaUAIG8
xUw4aSuIt/w8XHCdD2MhcnFxJSAdA4rZgU3JukRwGoww/EgwhGCuN/ci/X7P
4O6wnq3xujzIWCACVEsqnSCkE87ion2rpClmBwy2maDBbv0ctAN51QVAsn6t
6A5Nbwh6Da6kXxoO2DtcmxeWjfDsV8rcQsOXNRitIYh+ApOFBahzO1Fbw7o3
jYTkL/SxvgeniDh3xyVXx7NuUdImXKSB4H1KRFS4Y/GXi/OhvMBg+B5pNlOl
/O/zdShBUCq31aY3xFmHN75H3BbGpUiAv12tliivfX6Mh158p1+/dOnPV3rG
bHG9LA9kDKjxBXM9tSChCUYMEwwEQYKrM0qEsPj3E5RcHmBPWWIs704HEBw2
B8k8xpRhWCX5Tde1X19NU1kl42xh0qoLZZo5Wj0fNT8KJsE/aMQsS1JIDB8d
aPeoJl1mysrfglqXbdHVD9maTdxPjczslMeHkey3+l7JLavX2W7iPy6tNfbh
QMF1SaPVmle4gEtghKDhq9Fy62DYVu2bUmJ+PBGlTzRxfmOv+dArONd8/KJL
I9VGpIICh+RCyWHsnLXZqJ1upKtevuJK7zexrf6lTnQiI/VTg7Eqt5HtP1BC
h8oTu/lyeoA+d4MiIOgo4QW28aqI47GC0jN1qJTznVfEcT13grKCyIJB5ez4
yrkcNekwwiIfEz0drTdsjcvF8hBXL/mgtSXkzsKBZZm23PZO6a7kFN269qjr
zQe4TkbKZIWwr/PI0yPZToL6afAo8N/lgr+nlOgZIkSCGcDo/gqfnOQeEpXI
/AG9B0CVGb0plGWqZKphm5nrHjSG+ToYArpO7E5QmCMdHernzbj22DXlmrQo
2BYZNNvg8J3JD7Ryebi547pzfw/1FlKimFr11+wtBDWdUCOle3XC8EBhD3UV
sds3hDoQOdowZE12nowvGd1mfkjn8QeXNxl1SSw43NV2fG+ez7pw01bbe5tU
+O7jW6n4qacR7lncW/zTZ+sRTXdYCbTpfZU53X+zbkGRYw46AK0hhm/MVaav
JrEt4vGNbi3DMaJ4Zuo8umZYFuX61zz/o2EqJoq29Sd4ROeWuDlZJtWDjTH2
pymVhGU6s212xoO2sFO7yNo9ZOSiBZHNOYf+SKnaWDXNRBUJ8IpY+tfM8LEO
8EFA5KTJ4Q9g0kDVt1xTWESdUJBzhcIeXGOYboO4Gbat5eGWJMkXdYetq2uF
I6bGLQeG00npqseYml7lpnyFsnBlaHtf9ejqj4DMEgvXOkb7318YIoQl6xZo
1ST+NzhRS2KDX5MIOeCA4D83koLYfLJddZtcbk/spGSRQKFVg+TiahRhv/iW
DYS41jed7M1yH+zNpSd/vbHgoHNP8MTjwkVUjr7tPs4USCNIR0lN3h74RrmS
0L6K1OvW7BcGKD2+kzcbG91DwD+d8+Ecb6a0sD5+1gsHzXybvdkv6fiN55rA
h8QjufjpRPd0BuvdpafkKud3lBlVKvHpaZzgFm7H5jyQXSZmNb1gSiHdXs1i
9CO/fGnK3jCAQTavkTlj3uswDqKRIz/AaRIfS9jTu8AyMzzbWMPuj5Be3vST
6vs2CUvIBerVFWY0Mup1Y5xzeAy0htYh/ktRIieyrjqhlnyD8ls+cl+5fXjc
HMGAsxk9L9lDr0RZsW8Gn5rH5URVxb8ZffHfu61fMnRJ0SCYr83LL8FYgb1g
79ELW1OB1y6+Hi1khS3lHEItQqNXgc5xTfw77oApDYkPLTP0NXToCOLjqbVM
QvykzhEwpcJX4KqM7aIeYYs6pav7tjMvu/i3yVUEl1K6q5YRIdUDvQvLWo40
86l10DBcJkw2jOarNHhq7hdauFbwodcboze/aSt+eD33qY15Y/AmERucv69F
M4BOL+fQbyx3YfzWiaqtS47KZz242DGiyaZAbIXZcZ41a2paJ7KgV7cLWgA0
/eZx6WomC3qd2nXskcuHRMZRJc9CoS10+Pl3YPm0aLFw/RqneGYwsliZapWA
i8098RTpxCKb6u1OBrrZaTQVfEiyJ8PrqgGmRGHgiRKdd5fRuutGPb6ZJ7du
m+TbCZ0olIbEBQJbmiT4I/EHUQhIHyy5F1ElgosHzfEYxENQ2RkcD10UyPnB
yl9TzST2/fcNJd9DAxN0CNlolWUcyWUd3S+P/hoA2M1XkWN5rtIEK7qTuG/J
eK0sqxHAdNxnotf8t7+gQ2HimYpJ5gm47TDAOaeBeNm4cHPeUUPPgAMPUhUx
5gVpZrPDuHE2X49fWz7+Dyu73OyMkfwqXpk0/zT5U//6N44Xal2+YMt8h1zA
6RXSo/d7tjRbeZHvLLrMShGZuTxFmwQIhm99UF+kBtk+RiwJ8394n32GQTmM
NLb4QIii3809axz3MI1WnOpu2MNbIKba4Z0Fa2TRglqir0tHDs2vBK/G8g83
P+OWatifFxC0RQ2ZvZlmKsdgIk71xI6HduKMd7f1X++sy5NEnmwGmiP65p2X
70bFfkR5Lf94h+ijhgi41dZxIMtpqoFA2e6w7dtZ/Iv9R9kwuMVkn7tQyVwc
4eoQlaLAdUjVnP51hs+gqBgZOYeIfPNSO4DOHFfjHLSXkFvOCaS0vjlut9iN
PUk+3djD0FbxwVLsuOqLfNnpuU5h/lZ/efypFt37MvV/Y6jdhuBBjSGhUB5H
T4bdIYKgyLyg8oAsAtTNVKBfNatc8LohzdOWRBGPzWTGUeYzb4tNsaQheIwr
dmfg5skAwX/NjgbZketHGt/jihGB8ZBoDHW53Wq+WE/rCM7xVGCf/RfIIvfp
S/6qi+bc/QSrvsfeV6HXGBw70zCGsmaXsdcY26hrKdx0pifSG09fdIVnRVqo
Cx9RM88YRAyGMb+oFlRjt974ay9ePZd+0xziOeJfYi6W6+DEZerTUo5gL2Zq
rAXrnkeytgP34xnkwSzP91AG9ZSVRe7pt0ArD61tLfrxqT1q2wXm2aEXECGG
WzXtZ86Vk9oUossW6AxOFuaWut1niQbZKQbhnpnFn1UdqfqtsMc8X3bTKJ5w
Us1eZUiGrdB8eXfik2MauSeK2hqGQZgYJSZNrjESN9zSMjliKvCSzhfpxW6F
7T+h3YqrBsTxmgvNDe+l7NhKMdpzLe5xPmkyQRsXnee9WqkfjO+JzQXi44L0
nFK9YPejtUPFKGSd+Y7Ewyq2plVu5adtnCn2PRTwaB7b0VHczf30ub8ppf0X
5dB7wcoORfVQaIAwuu4j5PWbwyrmcjMXxchKwtMPevb5dFcGZrKoII0EUcH5
3ZP/ZzTOPtsMVmOUhJF1OqckV9p89u8byVf1cdCM/vrN/jLOU+RXEmVnn2Yh
+5pYtDdl+gH8QfYYfV3my2PdW+Z4JcnyXFJ3w3d2G1REB1J3P3WMGk6UNhH5
OVC2nvPyCcUlmojmM/lD0ELIWAjN1PFevlSGnVmYqsUKnzK4nJ8jUKrxan00
BXA035xawhQ4SZzegfklwsv/4yqPQh3JHbZX4EeZduErpjg6MhOMFmO0W3N9
De+U/6ddJR216ZmdRBkurY3WlMSWUnfPXGTerty2U6Y3HFFJSJ0sxUXmZM57
foxL6Cjrdtgk+5JursMFSpnkHAQ4pT91O3T9TrHuR5ntuI64S0gQcO5yIw+7
1nZNI+lc2U5DIQHyJRVPdJls+sEncNGHgbjSg2FmZ4427cUJc3UlLStsxeoh
xtL5uSWzgpZWVBttUN5Av8VVGpGxpbotpJj1qzL883EjJBq+vnCg42g7GyMr
sWwuLNrvF2HprU+n/HsaK2uBOzNwCH3NBHtx5tnbARJ9tK1d5KWzKhYRXwMg
XjNwOIsroUWghD91LPfwiciVyYAra9WS3uYuMpRoQ3DGaq0HwoAzpJBRlg7U
pCZTX7e+zJJ4mM6YLx7gt5usp79A5E8k1w82yLJEWuE3/y1a78cHERsqfv2A
TDRkmncC6K9qfctkvart4TSdQJZViCvLKfgJvjMY8CLnh7jLIAQEXJ7VX11D
Urzqz/9hrPO9sIH3st/30r13t8uGf/g66ZfXJNQ6MzWHHHun6dVitJXsulbw
2AI4X3gXn2z0Qi4JpPqtiqMfe16Q0vvHw6sMngLKQi4NzCDwNa7XyL5Ct2kk
bjkqo1cnqT+ZyrNdyewFkzBBZ6n7s7drOOgUehJ5k+K5rBA0+r46haP5R6aE
+qv2AreA4hr+nAX2iay+vbBTAy6KxCTFHBMHu6EKlB2zI9odaiBWPDO1AR8a
ytz8Mlt8wwhgupvHRMtOGDLEjy5adJ79dqULD1nBHpTsLSdQufhCykVVJAkJ
QQ9/OsekCaRYALAbpCbJuBsx6evi/Ta7/8hOayyatPTqKNrrArcSyq+X79mE
vmJVDkuolrQzFWIzlPUxNQywA7VG51ayzZSXys0bpjBH0D9LzpgXlXKi8f6u
3DqOBUK9nggMh5A1ymGOMBBb/bnEQUhlASzpTdcZWsCg3ZWkfgBq+RIB4u5W
C+KwGnidWBYypf1/g4nQkVoGrBySpy0K8xwjBtRjP0uNPA6h5G4Phg0KO4JF
o1e+2SIUxUAhvsmmsbadzxLfPxnXjNc0voAi9I+NlphHqy9q6hrSQy19ZHUe
cnbFPL4QhqZtLERArbEieRAyr+jOniNMDYwfmCYGvVSFCKu6RbEEk5aTftFk
UAci1IdcZ8gU01Wfgu5fmXaWpqG06F2FGHk7qRQd9guxZNY0N3NIwghEGl4a
xe03BOCPsCbi/3Gk/m5gHPgZdq7I/pP22ss52pTM2zzXLreo9mVmd/11d1pO
XRllsOr26lwx9FPN9EcEVZGh/Y4UZIiD7ltVXnawvtQDLzTd/G2U72kT3EYp
EeGgPEg22fBq06D5Sh0jaxTxQWfpjA3096lD4vq/sgjsHls57Mp7/oAYLO0A
jG9hQi1fJ5Su3s3yU98Tncy8y2u/WDrjgK9yHi2xq8z8C6BW0WfTM0hguwIP
YdjCoYin6AF8H5rDorbA1LLUsYzwXZNXRMqoEuRHy01c6Bju9XAQmBrOU8UA
9+eNdMA1tGhZ4Ldlnyi3DPJ6vk12fU8GQQVF+lYEWH+iwSuR9zQoF7kMJDim
T9yZ3WSpQ8X0nHyJq4CEd+B9L+2IcIiX2BUOgxDruHZm4mKq7KOtaSu1iXRI
HYSe4BIbGj+qAQAhsrjuWmEyXkdF0v2MlKKAeJHDMF5hFgyM4yuQxlxxmKsD
1/HYckePbDtgBqicyvbDf/z2M4HPkHd8kGsDRzMBoA41JyZGBmbEf1JflXNU
7/j09t4O9weMZfqyQafZk7kC07wNhut4QngzFNtWlPmn6hX8yFlxebOUwvy/
mdl7qDb2Bo0Tvx7fg3B8tlIYs8EV0ebhPvh0qqEs7r/fC4H4e8ZkxgoTg8Ht
Icd4iIVv5rAmruuq67VEFQNUz5/c7PT5pFEErS4WDOHrt/hL70PHmINSUneE
Og9JdWteU98gBx0gydUT0A7gzMiXD8RgQirGui2C508E3Z/eoRqmsxGVJz8p
AmeZY75PoaP/p4hhcp6wmTUq9i0aSmsnWCKTBzEqmNkf+sbQuPgQxYrMx0zR
UrJ4wo+/7tmJao8kwIUpxKpNuatKccaKyVGJTMuNfoPQZwZ1ikot6RpJL2IH
d1+/p6He+gB0GMc54BuqoxZsYggVaC3C2FEnBJElA49mdmKHnbMTYpmLDz8N
NixDug2DUZBpAgNt6t36gCYcmMdI5wDgYzGOvFI/dZHGF2qdzrW9f/rccEQ2
RyvjDlpKA+l+1LFUe0jYSgKoDsC9wrfvqQaUg6kZaGRyEel3KUf3nvCsx4nF
+Ofb3tvW+ASHXm+/DOzvX4CptlzkOgg3BGzWym9EO24G/EbJwoWu1C8h9sGh
1NUW8KkoiPpVULI0SSG7S288K/NZrWlwIC6aW22S+Ls54uBTVUSqILl3DiFA
IQ2iDrc9R7HFxBMwEQyZkLT8NnCkD6OG+aihAvyA3pX+BKBL51nmid68oW4+
6rV+bkX84kG2o6VPB9oNBWd2eCN5oz96B33kGqCIySr2x5p43JJvra4iggbS
ahNBx3RY2BZMCEQ2SgH0o81+bSq3o54uaYN9P6ZtJe+a/H2j//eLgKBk6tOf
KNQdog2X0A98xcIYbE0GCi8mr5pgEk0JzUnDzKghvxSeCyfNVdLWdmxtUqnZ
o1wM+QqqDH/nkl0QW2mw4BhwLp4eyDEZTKpfGb7ouCILSYRURpWAGoa4baaF
0yPjIEEseOqpvZ7il20W1pSOb/DkMCD2aZBHGFNKz4tTSyTuDRkId7RK95cE
U62YIIn76LdP1vpLwVWkPdaM5QS9qCN1nSt3+LP+jw4nlj3QypDrffbXX3B7
GT8/2gXWx+fjVepf4aKeT2HvrCynRDze6oOoA6SrntvAYESxVDA9TqzZvrgE
UAAi1PPWsoSfKs1Op2x7FGkfpFUMS4Z+XHt2Tln7whqVMX7EnbMhzhvKSckb
YDUxXNr6OLwj+yhNBGDzlQEwmCw9ehdzcIIvB9g/oZ+KGTCyURKdyhuoqnkQ
Hj1xRKvpieCCZNDbNmHpDjWm0iLvtxPm2hmAOX+OgS8ZIaBNfHEmzPSCsSsr
wANhS84MIWfmxeWFRGGzCknnlgHj3TRk2Ms6If3pQibzKPoG0YzbotDKi3FK
Zr98OdO2tzwUqKO5G8/dFP7+qSX89HZpQjVGhMEnkZsPNvBmXliXS9UCUB01
11kAS7yhD716NonnGkADYIQRP9YJvf1VU+IY5i0SzykqKOtAEZpwkNyID9TW
vLhmpAAaraZZ+itMXOG3gg+iPmPRDv7hLys+8X5HTyyptwWERP4onKQ1uqCn
E67y9KHsOtUFpyAHuNVg3FHuSJ/HeeVJJoAqzX/4ghB7cSvsGZ/Gn327+DSu
bsZ9vjbez9YQ6XYLUPrrTvxplBjLgahCVqfJ+FO33sfpwSZ57Ul6DxJeCEFw
kzQ4uTUr8fzjz6REHXCuOVEG1IV4rO7WZH/xtQxsPCODDgCSvyGNpxUAqaVY
Fzcnn7SGdxLo8Xo3eLDIQHCGXO75dPCSSe0SyuITV/GxuokDPU99mjh6kLn4
oSrDCM6wZXEbWlH5mgJCAtq5OZzo3RXY3tiqbDvjSeJHCE8V01yp6AR3pBpM
sp6OrE9P5wm4gkSKkEvDpOPDjiaPRhAMVr3sbAQV2FUTyEm45AaiobDs1BDx
M0QGM6OjOYLoCXI9qs1aSaahdR6yvz4MkbuNFt30OVWBi6CNhMnvRPE05d7p
7jtTPRPFSGMF2gm+UI0kK/+vvJTTQdaP04s1qIIWMz1lp6hDDUplNCko6RGo
jpTYbjigjdxOotTBJvfRcJY6rgX1qlsQAd/4Eow5VAiPVmPc/rEHRb72cHkN
83nTfmZkeOPqqRukn9IMIurUx07KsjhgUk7CB1urWq3+3yd/YfMgM1A1qXQ4
0/AMr61VmHx6eBJRFV61khOF9Js5CcTyDteE3Sotc9ap269AohjxHA6POPSu
IaZooVRnGGjNOWG+7CQmz8DNiQFu6wGi2EdSJsoFXN14A1QBDf0H2jUlref+
1hV3cvj/LJpGqe+yiiB6gw9Lw1jq8QgHXMEY7LY3e/SVh90DRHrdjYzNF+Il
SB3sct7oboM4Q9h5xYzL/aStBFUfn/dn3WN7Fe2+lxygHcT5vD+lZc9ZBqWo
a7FVM30ZsshtwSNoUvMrSzw5V+vcIcBqh0xHtOvmkvntxV/WrOYjUzpNYZBE
ggr0bhCl26cnBU0q//ufVSZGZoUJIBJ2QpE13yiMSHs7dkYsg6QujfQsxfFG
EHkvn7aVCxcmQ15mEByi8+0A6z2tPdJcEZhBTor140K79ybimmYJh2klEh+9
ainf/+cZz4OQH1BrtNQnzEY9NcjyZLe9GfgzRSnDz6ngxMPukzTLEiyy4TJi
T53QzrJyFx/YiEN6VDe/GLXgBMUUbDLvpI5HDR3dvgfiNBO1IR/iUR/kUDQU
M9IrFFixtfgSmT/eYW2+Wlgs6mdkLkXDgfkBiRYVI64nfoPAlK+yobQK1LbG
jsV/C015higChgt9o6heFZ7+dvwanZvIvWQhLvXFa8v8rKMnAOBCRYSMobV8
BqNVBT/MX8PJEEfty1OZ6gMpF1NHRg9u14echLPt/LHIzZziGO4rHpgua6iP
kuQjos9l4Qm/+KWVpupksIFi5+hgUxVouT50uyHOXVAGCR1wCJpz0s+EwQ9P
yGPvTpB2W54R6O/s4tP10Wr4hGptrj1cFRhbgjVMK8ISETknAltzTSON+KB9
VcnO4BFRIckHzUtclKD3ldE4BlzGIvyDSOJRhsOzEwOB/USf/Elc2HcGpmiF
15Rtawh4vco9chTjRVSBo6s24yuXFpznZsNIzUv0Cj281yq0Z8oRmvufcU1V
LJOrn04hOR+6mB1BphaL7vX2zcFW5VMkY88A8pmqU1L27Ebt0zIENmQ3XccO
AK9IFkmAfPC/d3b6/5lyINhfbwpLwXIzFjwKxFFQZt0VzanszltuUWS6FirE
aKKRlDiUVzcfsttGowT81wlsuMo4EkgnRbx+YPH2fhbRkoIvM+PwF7JkcteA
2/1l/KantDQj3EkExjVPMOhFo/WVOYdgT8HH5pFxRwkcltofJkzyhFyCF7Vb
nxV3EhrJIbEpDy/20hNjUyO8LxvQbKFn5vXiGtA5UwxJR1To3MmRNnxZkzzF
/sUIhFs7Ahvix6Aur+vd9avQZ8cMtZ1sMdFdy8vaIiSu/nx+sm+zSd2WsZkH
OF9r9iC25ozb5migWIVnzsONe1apJd7DgiPRxNrkH9r9gedfBm6Sd46sSOUv
vPMu9UmX02gl+wY6Lu1LVFmOrXFlYywHXvhSuUg6M2bBkQxE0a5nWQxFMmco
7vmB56hEx2LgOrD5CDjGc9FPT95GUMGwKseZZV8Ue+/SYNL3coZfYVOLFyae
j8Sw+AUbwUugjOJhMUgPpv6BjAtO58ddRjVcLnXyF+guzDzftbPYuZvBv//F
EXDqMi89k9PCuE9wssGdes09CHFHg+AQKa/d0QP4W2rXBivGAa7lP/6ACdwz
d4vKfTv5sYLCvSccOU84XJRxvsVI6ovRxZPTPBFEH8T6hDIumogzbox5WQUE
3BLQ9G6wydNQG5Myz5t9MP49PgfA/onj0nJQ2UwKd4+cQbC1X0gfB+hDdYMu
uKanof18XEYEMAccapdBlwvqRv1R+uJXHs7IfLYCLq1lJB23NQima0sGYwx2
iTnV8+AQKMTeNLz3StcIfuoDKQmVO+Fyk00ycqgRMD1rSHtpB0buGCTk2cBw
dysM/fq2nHtt2gJ4zLUsO48UnQZ9HSsbSBsFz3UeFI3cd2W8JLKUtsK2oCYs
ZyusxyagrKrhTm2EXVKGd0KcmJ+VMEurAQ5MpApP4VNkZa7qCwuoGnpX/iDs
3jIY12WiLsmeXL955PEZxg8B0quiGeHy3wLJTOMazdkVWEY9UQXypZAqx/5g
UfI5vv+1cNZrxyrpolbHTqt1bw50KeUNQTTVX2XXQ+aK671ohBjKpPDRTH3H
Q5PNZN59kVp3caaDv/VEKUSn9t2p4lltmJdpZFzs6qAcVZOeMZ6SmQXR7vJQ
27wjHFozHjqNSX2OQZjpEeAWBFbqMRUAzEfuSfwdUu/OehctnE7gk/xxcBPH
FTAW/dgydsiyBTxPurIccoEPVdAXxMhctfOFLl5fph79U6QLNtYS2B4MbGep
TmaKuiHiPomjv83fXjN7JI8xc3R1Ds49hNr7sk+/hLg5gbywo9EY9WZtMX/v
2EeZOSq9nMNyzDBs814tNVwGekGiOGAC9OeQxrmTJx3wY8GAfuubQ7Gj6CcH
4xkVbzCqPyOy1hgVZbi81OCqr5swAyd4XlVRcHXVBSZfC1O+BV9A31HSeGNm
VxY+mbRjqq9Nm3Erilp2Vbr8pKmJqjzv3daq5hvdT/K1HUzvLC4gLG8uHhSQ
1ZGqeoLkGLy99DsU1RghynwZ44eovfY4ZeeyS7WNrmMuPdasJvHbAcn8CDV2
LGqfOOD/ENYsvHKYby8F4ZzFdfdR0wATaFO65eQWVG01hgmXd/y5I0p2dzKq
prHu6wrmBtmF09scWoCWJKI8cJxsATmFxpeBmLzCWBE75yo4wOkR8TUroANN
xGR0s8dhbFKs3kE9tWYYiFBGLN+5wdekj3yKAelXAgeI27eEggMmWrwktWYA
qk3m3td/xzjfcvzepzYYrjztSnRWFsYxDlOLaK/WLtPcdu3qHlFLzjfTCqu/
L/SMjYHAKKuFk0a83tuPNSoUcenQ6dkmWqo9kNVbkZBY8XqdkNPv7ybB3q7I
jO8zbU1QdBCJkq14vGz+l1c7/zE9ePbjHif2Qr/n+pccQXAuw8MlHoO4pT5B
HZfV1xGPztOaokfvp9QQipjr0wBM0Frn9sN+fnMB3o/8L1IY0wGb+uda7f0Y
L/4+mWJncCfe8ItDSPDbGPAdAlgjbpeZKT/bJhJlWfQ15zA722ulNoxcHv12
GfWGbnpMnaIdeYI+xQMPuusb0zSaCP51jnPv/u4cpShkbfISYxl7322i6Bga
7gq2mZbI1X82PLHWfTsaEDDmb2fMXNlo3NSusctTc+3KNuBsxYhJpigC9ZvD
gnGuKN0lGZ4fYot1JZB5gNltmUdlieEBHtNkp+CMBsXkGW3M9S+4pj3IkmaT
PS6m5jlPPjyjxy63IYoOeisBPvCTl9tM7OT0lTjRld3KZ/ZaANfngDrCPnNC
TLWCd1f89MPTXWblo3u9XRxYwRKEjslJGtQuo510cN06qsSx15WIDZkLwNQT
e/4mjWgvYChCYKaJS4zSKEHbuwEHMZQvMoVhl6XeDNd0Dbsp/Kgm/U3+X4kY
23SUQamcHXKzwslkosFPMLRrt6GFlQCVtEsn/hcQIgv7uBEsq48ESFg1Sov5
9P2KZsVQWeitVKW40SyZaa4rwVq6/KjIDUz8JhErxBy5f+y0JoY0j1Lne61g
lFTzHgxjeZxLmsvo3onoeqIg6F/IgHH7qtvaBs2pRnezMxlWjAFe6g1pcpo2
B2UROs4Nwu4R7wkM457QnL0HU6AHCZSGmjuNcv2TlSN3EotbnQNxMJ/tqME7
8QG3C+GTqzB+vFmVdThWtEwtAwo9tIbXP8/eyJ9a6/3xtJPpR37lipXSf2vR
UH+2C6RFMPwWAgpeP06mbRr89stDiwAz+hqogN7K+9OLrLmHDvQSMBpkh08S
hjZv5E7eVSs0BjLz17O3j4NbN7iBTA/99DjPt8CxA7Z3Kjw0hcHG8SA1bCVR
B9w2Ysta69rieEuz5dsxZT4c9u6LVWKtSos3jcyeXDJvNlWP4dYYFIR5uR+F
Kp41KNiWJ3fog3QLpDCLfRSBicCMJB/ZnJuOoAhl7+AIYh2IHjAuuPRgCcy1
bP9IB8i8fs5rMrLI27n/CZw9S7VdycNV0X8dX6xIOL2i+IMiliVYAtsBHba9
U9mf9n3/GFsH9lfq15HbOiVbx/OYn67wqC4za4SiFSnuynrU8hy6n+li1UEq
qOu19OglGh/jUXl1zD5i9Si8N0jEVJTHTrwHz1yPyvvKHx+7lNpWWAbH3D0U
FmynvmmrPnU82TWsRgjI9c2yKPIWqmWanRxII5e5a64nLH2qQsp+q5Gg2PW0
XVJ/+g50mFbxOVBxVw4RLXpN2M6EBhSVtAPxnoGOpMVbkc0QKaoepqiImPKQ
aP3HFzTI34JOH1UwcjCk2DeYX9gqJ8XOBHGfuydO5p7ddZrk/n6EDpcvdfGE
QRGCdaJLDOqg2mCwwLbWfB36Bo2PthtZ5S25ua54f+HT1gc9qiHshD4uqrg8
azw3SQrnpUGApa9F/81fxxU9vOJMM28AuQWLtSkuZNZMNS5QvDaSbPCXo1u0
BL4s1iyQ4LM4FMdEG4IGoGD2mL3sRwJBAPSHPNeDG3NXUWT28lUdoUm/OoUb
qoyfDXd4mmgp80iiZg9vrtru8omTssbX/pjzTrxccoPxeIc1K40sMBKnfpQe
ncu4LRQgSnXQ2IHwx0hVlxpFm0fviNNhQ3lgQ3g2vMCnE3nu7XTvCIiDCGAG
vugqaGB0Uj/Xb6brdRuXhrs/56kpBjHZBU7x7jyZQt2ACFIyPdLTmyyJAmgL
LpzTvcuoeSjUgklxk/nnENfmk0zMWLdWiU3sfvPG6y2dhHeH9qgpgPZCeKTv
K/vbyQrC8M0Re8T6cxT3lCbhV7Fd/s2oixTTEDhWuXJmr6+rO21yOMULIy+O
NqRYZwm/p6xkrpO6rvzHI0fZQf1Q111y4jbMPneKGfDMq6rS3Jcz7wtvQiSx
Ud1eruo3vS87cBNFzQ0D7iRzVLHezPq9f2pjXvSkOVQ4ssuLgUQd5dLf3vsz
15N9DRhfHih9jG3MmBq2Hw6ap4BSR5V/cal4x+mfKExcDpihFqcDqDL9XGFC
dUHOiCRHE1X1ow07awEnbIW+EPk5jldweXrBpelUzuN303FMfcX6G7GtfmiL
EORLkgrwTzFJnoXr+mcs/jMakJs0BY6cXpnFycGbyQRNpwILW5F/kz3uSd9s
YyG/o5kTSciLk977h6mZ3XphxkNpAAS2mHA1LuxG5rUQufVdgEVMzpX8P353
XIxptcbis3SjclN0FAZYpSZwVlFS/7uXiX/3qM88b/OoiM73/TS0qROSHVt+
bUhcHuLMupHG3OP7yck4oUrv/AseVz6eMFLacJ9aVSmUOxRPO3KRD7CsuNwH
HRoyGJqHKwCbINSuRJngqAKvJxEUWMMWkx4FtJP6rh6WhuWfyXOzmNuYto8A
xmA9Z7jBrEkovOttRd/kd6vWCWsERQIhCvaAh5HBu6hzyXsnmio6JChF6ecx
syCZAlHb6avUvXr7sR+QBHGfqjGFul2v3np/aRWAqEoV/maAsr0lJonYKRxM
ZUMcCgGF/ZBNYkkNabowm13XHwSEqR/8HT+WQ3xBfmotM9QYSKkm3z0/i+Ih
7om4nNcYfcONxJ5dGozuwnBdMPAyq2PiM0xSl362MtZcEabvqGedH/Q2rG9e
4ESQW42/CaQm0gf3fRjDcECxGl7KUsFzGGCctvTLq2vSKeB78qr7ph+rMVq9
NOspplICyEwV4sEvw8rpF9PxpNAgCV+8/es6nLtUWEAt/MBnInvaFvLodpvA
qA8IvyfwKaR4szgtFKmwImfIOfnHrF0Sv7ksBRgzs/UVVV2p/WTXbUJ/ibWD
ap7TYw8JaJM06hLUI46r0piQYNbxHLmbeB4fH3RbP872ut+TdhqM+LTz9Qtj
tAIFInBReqEngCa2c12u9BTcpG9IUSexl0SyzGV5iNdm5JFMhSJpz7sYiAKq
24zYe0H2Q/qd3iWu5kv/P2vvMJx32qSQI/5FFa15RK5uGp8TY2c1+jfKT4rp
XbFYXe7OsjrWpqslYs+LmJpjdcqSpqESLD0LOuwfyKJt1AjChzGeLXz5aZdw
dOw8LwJjtw0boUBPfKCFp0bosByNZt7A/LRztVc3CpiRA8vFquEj0T6G+sVX
HAiZrFWpUvhJTZcGvw1r3QeEgufKBqvKKw9deB4K7LgBqSf3GxNPv6yS8gY+
bQM71+WjlU4r374UYPxNRHQIuOET7LcKObdfOxMTFXvCU8xliTibY22OE4kM
UbFrEF3IyIosbHnMRu8VGFQvedRKTtaaFfvG0nHtJhsGDHtPsyNIFzfyLfrf
+4gcMei+my627IX9HqGRPpnmBtrnIlyZLnF2BpgW1HC2nJGQckaNkYCJILPF
4bzv/eOb9KD/RqUnecDHvkZtlxZ+d7zq7V+HGBBbhqk7Uznnb+I0lfab+FAs
zfDnq1Hvv2OT/uZpefTCCD79wIaHxXXSlztgoUb5t89Wmh+8qhBgb67ypGDy
Ix2SRc19J2du51r1PNV3U2Ye1WP/sy2CQoummdLOeQXM3hMcHAvhbVawlqgU
MQsVdFYfRxK4SlNbshrfB6xhrpQ7zlc+2wfN9fZgZPkRgq1I+YzSKwEsyw3M
EIAcJLdYLGivwLTB2BFLy0WDX8X3u4jfih0UZaLa5oTMtrFfwKX2x1TXlNjn
pw68su3NafehuDXW/08j0u7zd2zxqmXOyxvSFs6f79oHxlzp8Yx79pHw2hiE
6uC2Tam4u16kVvsF3D06PFHU+3gKzl7CEXK7xt2dnghAdTVDFELvWlkLW7Cj
kAV3Uu+TBUrS003I8dOD+nwxScawrzTCaGW9MSJnSzbff9zIkQ5DEM3AHgyt
U88BH6EEagHq78polBu9AFLpGGyj1kbojlrCH4F7VupBnpl7SNUm4zSFBIW6
Mq7lHMmAQhTEzOd3yTgFcSznuE+tGpSyDh1eKIh/bMATo3ziiV9D+CDLqCrQ
lh01fxNkwB0E6RLXpnUTuet0MjLt8kRZaJOtnWFjmudLjIzO0wfTmHzWPuDr
RDodHaVkNVhItG9boF2o8FM1Aq2UIhmnbohULcQSfcqCr2t9QgrXxoRgwdd3
SpTyRuQwe2QUh0TkXQIiTSNmD5KUABR14XHW4pzbazwVyou5lUhi7x8Gavdy
w9APCeqEu0PxuBQo06Pc63rLT5O0yKBhRgjtTpW+eiHrWLDeaNiGxsqxdHDY
dW4ObVWPTRgd1yOJvVVAv1NBxXT3YIdAKejPPN6FTDW4zsMCPVDztemgSaYJ
HKNV+/HoIQpEpqrT+jy8U+HefJCSWu6/1c7sHFlX+C7GVQtcDkPq/k+OzEps
agYaNplFvCtatsyVbwFHiPWguA7qWw6yZI30ZJL0ESlaQQMfFlouPUeH3ley
CJBqQ4U3pAmQlHZVFaN53MNJg319+7R/DslNq6OlOJOj1NPjBjLBXYu0iRUQ
vQu5IpwlcCnKlQvTU/TbM+49qaqWbZYOb24omdUYO/CkTR+C0Rh2TvxYqc49
JsEgOnUhrfKNebgvhAJ7GWnOd142Dwof1mbho69ZLwNY/2UBzVyvXcrkeeUU
z1eutuS1fhyhNyuu8RzCMsnmB02BcGKvRxIm9T1uRwjNbq+vY2/ABUiwdO6m
c67GrTLBFLWStLmT4HHs1HrCmH+rGNKMtMzWB6rFwGekDcqM0uHCGLrXQoTe
imvoCZZ0p5uV4S6GBs1ZgWaqTpDe9J738vW2AgEqWktLRCStltkrOD5+akm0
STWjAXhL8+uqgwnlxRhbCvssZepj7FQjVEX2rGf3z0arO4Dhyi3TVCtyiVIy
sBqT0ANTdim7hyAc15Xe5dPyhWryoXmyS5YKL6sxrMQucXcI1dnWq9DKptWf
A6lA3ajoPGFdAOGKJBYK7C9iyGfREdpUKzLOyT0hnoclXniORkmFaQ6YC5GN
YXFgxGCtSVn+z3kVZxfgz3nXFU17O+bnF3Zs/CrYKirSzO3bOkPdA7sKvPL/
J76VWUErAnqtDDFe9yfDhor6+Irn3cO4zkTfP1GcKweYrHxyxG7y5ZLaJ+8D
fo8e6YMkjeMrFs4OXkBwu+mwHVMAQah9YyaskvUIxCvkpb+wFwai656XynUM
KgApR+R4Ed22E9sIps3XKtkd0beM4sbN91D6ZtZOsVBXS2uF4LH9dNKFJiRJ
i5+SaVPkl/S5ZnO9amZHZXOwgqDIH6ZtMuF/Qo1Scbmqadwgsiglqx2ct1o2
oh1VUu2k5guENrZn6OV91oDXHrFFSM+wFUWKB1WByh8QLT/ZTsDQKQzsk9U0
FEjfL4tK4ufT54TWk0eKfJTNogiLir5L1oqchNnI2t59SuLFugL7f/1xydOw
ZWDJ6cfdGvZmWAptTTfEJ38DUJGBDJK4JNJdTWW2OCmA9MdUfPycuQLp3za2
ukescyt175HoCqFsSdapPB8g3G5NgNGVp2HQkoomqxNQoOnmYJhZGdfNsaEC
CD8Eu9PI86unyeJV7lMDodn8F0JVYB9/mQ0X5BIFj+HcsIYp/5UazktxkJSU
BHg1NxxsU02eYbdQa1+3YoCEdepygqe9FlIJO/rM7s7NMi95UVHMEBgi5V5B
vVVcLTgLiIyZjlvncRpK3Y2Ie+cZCUTh4rPiYtRe4kUnxpfX0RZnpBN5oYoU
to5vopF/65jdKapWPC5mKAPScJgTeswhf1+m5WB+uJ9S4OI/AEKMpvUOU46H
7t+YATbcpjMC+8Xe1mLngiiwI3IH7QALtRVM1h9gTSiprECo2kC0xnhwvDqN
TZNjC/391ZKetGVRWyRNppLlE4sPzOa9Q7uqKo/BNYelhhTpnHhjs67DHJr1
/9g8RntQzsS8bPVWVdy5Bs6tuXnwdDGKpPeRJbhzhups+Bkiymjpue0nYoJt
8NpoJHbxo1P0prwYP2H6JC5gedoQXBFRTQiE+48AktE9zRV49Y2iqo7V/Kel
+gMWlXSBWk/BPWTq/YIsc25/+YvqXOF5cVyubnBjoN9Y3Lb6fL4Fq2YrceLb
dUhWaGmUOvGG0BoGjvzHKOsI70EA+VqYztZqYEkrJlQfBgwRCuiHkFiLb0sP
XznlORK8gSsH8Q74u4yiezmASCH/EGAJimwbWvtmWgE/2K+aNpWUBqKQnfKZ
RtWXg+Xyoh9AmkLoWyPlX8GI2wtaLdqQDlvSqg9VKr+9M5d1boOyVsRHDJGH
v741OqsM7XSfZDh93fwDFwoDIpMzqMjmtBcTnXLLL0iMguu//qz+Gkq0fUK1
WeLVJbOu73SPjIJPFxt+SZDeM4ilpU0qLOWx6zyjlREN/ECZYUvkJiXsrCio
ZCn4MNNvJr6wzKN2ffCchnt2CMmyxjmIUjoXwy8wlkmEZvqLxuw+dG+hXpGD
kJu0zJeRDE5F2Wn91wafXC7yDTxBCmH4AKPAmPKEnoQso/kK9pGHyTZeqjBa
rYaQx86o2cYI5sXafzVpSHPJl/kjm+wONztvblXpDYVyqZEn0w1lc8gJTSc8
tQExjDeVfFx6oGlE7eBI/8094Y+/euNCsJG5pbbWXqid4yysy+eD2ozM8E+i
xalh/1gEQRlFFNjSyG0XJQNCUxH9dAdhNlHI22M+Ogk2ybNuqMJJbyutivsX
2oSmjzBgdpj5uzJSNiT82Oj9iFNbwhz/LNvsRZzBlPz725qXEO6s4SCLoA6Q
fEE7Rn8QXY4uRrZ3GGBm8SK9/D1WhOt+DNs9LAVjK/poxS8ODO3sA1p1AeXB
xDy9i1I7SC22gXa1eYQeZn8Y9lmeoAOf/iiOVhuMXxn+YkWalE1lrUQriDIp
2ygkkmdsI702qg4Cabxp/y1pz7h93PRVnQV91TXS/MVmOq5xKfcgnkZ0JoDy
+TXz0s5HUqKlZjJHr1UECFyB9LLlWlOtoyqLn6SeQaoGqVqcUXIKNYyCTRUu
bIJJgb+cqk4mGJlCrmx5Wo28KSbi/gk7Jd9Xlx9FobplfI+mx6lkDNZDjFsg
ZeZTDTQOY885hWZH8KHjldaJLtP0zPkdjlmQ1s1jIPbQDuM/W2fwctHOJC+F
oh1E9heO1eWMLc6EQbuddVnOFv8P8HheQk5Ny9QFA9uiQ3H7txbbPvgwhOpJ
UKjQHN0vtb7s7LDbN3LmKxikDwmGdvAl78R6HMobaFFuDh5m86E0MhyGLFpa
k8RfNekAMEZht9vjayYQNfUVH4T57Ss00OlPIT+I7y/S70FqIM4Jo67FvPDr
+/fJ3rqIT1qdMjUiTQ0vs+kQUpI5HoPgCOha1ITo9jScCBRZH3D6iVJi79i2
7gf+HHICFbqYR+eOnZGKKQdQ9VfQRHpjCV86SHYtq7vbYfDTn9GQXtgbBgFZ
fkDsclrW5gjkLD6lNA1FqZ/xFRIyR/DP8WRpiivPeiDr2Tkd7SBcsvajPkTo
2BlsiARiWgFd2ynSEXva0sc2rzjio6u2Hc1LYIeDAlhXcFiuNy4XBG0frSfY
u+aovgpqrnCAYvRNqY+b4NixDQrHuX+ZvTTV9ElQ6dBbclTAr/O6mTjZXZl8
1uoTXFHfk2ijyjFEBCSu693ejE/gABAw2Vv/zmioEOJVsQ5XAFdojYcGQhkO
cixZClLApDfwLRxIMs6VAtWWYXWUbXf0GxAQ6DyV4m8Qzq9emCbuFhuyd8tV
ypHveIEVAYsyLuH0kKsiq6ySzaY3+NBeSEw6p/qhjKDI+IObpDb1wVWA5bQO
yxGMQOmDmv9MxBKu3OIJflUNh/ThpR2BOmKVvOjWbjDXe9i5q7Oz2i5KaoOa
8jHvpJrLUas0YiP0YwsjX6lT+iQwnDMBMqi22j8hVtbFnWmvrgYTXTPQDogy
k3JjJKqjN7EPCpsVOHys27aE95QQR2fx2yBTopiFffjPPRvMYsXsoCVOBrA6
5tmwrHmYGSFS2DtOGWezmNcV3JmMRdOjlC1OtGNAMdbHghMoGnBJ0LO5Lfkd
csXqBGMqCBG+2Gbf7KN99PL668yOEtED89SgpgvG3j2QE7sk0N7jt3WXKyB6
Wr0scLCgkoXyXUUfdCCJNJlEMHmoFccV6VaUksKQ8tMbCdeX2PhBynRWJ0j0
ZxwO5BLjZSsJutykFbQYdy/aSC0tJvuultXs5LwobfxWWriiGZivFvdFPJFS
BehTVg0Z0FhQAPOCaexV2amXu6L5LWbQJt7TwcjW397GVhFjhuBxV9ISIR7Q
cGf/QeRuYnWVSpAT4YALjOavIHD3rlSlRNIa580oGeAwew4Ulxa364C8nlir
PlYCE3oPxV2vcoyNzXCfcMCRyjOykKFaO9V41SYhO0zmTz8Dak/2peWNI9J2
I+NsrD8bSXRADBttyWtQFep+qUvWnHNEheLmEFSVR38OTr6bguUqSogtMljs
M/OEBa8TBWASR7K2LsajpLkhrXSOtfHk4PsIiMH6tqRP7QTLWHEIiTdnXNIA
jt0bm8lkve/BYtj+0GOJEhHzKLSiX6SZESw1akpuGgeFIUjKMLWFeiDqmnCJ
kfqHh+NA7C0iJ120Z4ME9keb/feWnhbyLlf0VLzSatmatO7vzYOOBYY21aU/
Xvi4dNC2GDF/vZBp2bDvB7WdtzLcZki1YWLFWwnE2bVQrxPTMJU1QC09Hjkt
CydFKXjWP3uZ5oWy+HPkblrdM0O8/aFnU3RaKEydXEuQJ4RDw+MsQhWhOYzB
ih1pP093gSQ9l4KX82Lhr4lGRxu8AN3D7EtrZ3pbyMLN9WTisQTR1AvbFLiM
Z/LnLuDva0X5M/Gj1rdooyHur+1Zof1Nyw7JvrEcSibkTgkSVYwCcapt0Ox8
0hiJqiUfVOjaaL2OtljDS9kOMizvFhR0VE5fffZMUHSEGW+609PkzUOu9iQu
ag5QJOJPn/DByMCZkP0B9lcW8PaB4anallQ/ayc9qukToZ4L1YomJvgoS3z2
FbaJP6Q7TxFbhsc2Vha5RftRk1lDxnlSsSXeyIbPNzOESlM4+UVWuC0FY6L9
Gj4nuOk2d83sNQLWbPaY5YhIMwTm9ZoKB6EERACKGQIsd/lCGRgJiR+2kcHX
5nxQUYhDFZNHA3l8fwYuE1gy4Q5gvfV2fYE/J3/rhcVNy0Dg2kxNzNH+M7wL
Oq9loKkbLspteKEzHeazBUv5BF8Ltau+02hZkrZn7BQUiXhiZtX9cFajUvl0
+l198KJmKtt8FqGj5KCRMMWbqFljxy0s4h/Yfl/MN6aIE8dhVOznalZP5pSv
qBqJXmR8P9pKfm5KihUgXN+mphMYqE0Mar9QuoQMoe0DtOBG4KS2tBlFo05v
7nclNn75qetmVPm+KeT0jt5010lKAyue7EZ+ewtGvZrAjUp9d+0qhQL4s8Wc
tEk1AzW8/8IXwVOCX+offiVO4yJ4d0xLWut61rYbqzmbyLpr1uemBabhthrc
T3UfgffNjoCv2FO+eMS9GYoLjp3LxColknmi+YMQhSi5oeAEZt5IMR6HYv8M
TbG9gQ3jVHmap2n6+mSNn0aix5BckoYyWgf6e2a3c21jFN5R7KgYX752CKXh
f4YZk76C33NVc6XdnkuZd46RwiSlm5Pf2Bl6kZAZnbN3wjyrKAA6OWrkBPkC
GAcLuZUHgpwoJxDV9IqGc5kECciIvR3EtuuKSl5lfLrhqlZBQ0kkxEwLZ8wq
veI4/HvB7jJHeVA7Gye3R8h2CX3VMQg46zR6JZmCY3BA3IfHntGpMRrYyTxS
tNaYXgeKuv2VMmxlpL67wTiRr5zYLAxd5kpM4gJlL48bBWAW6ps8hcJ3dqli
g4WLtlT41d09L/oPPZI83HhYpB3Qt0iHjT10xhrsVSHTn0FRIgi8cMZiqKSP
p5+1TaMXPpOWbcAxUmGFSpS0VqhiFoy6wNkk7rMqtSkIYP5y2Biyb7R46pbU
ksn1S6D0ISi6sVPHVg0TtSmMIqZNu9Wx8MkY+tdHsZopdeuhVV0CZ3ZrAnXE
6kU1n6D0hvHKzzV7q9BqaYtd+nZsZkPMIvB4UzBE2CyP8eFg9Ym/HAY26Vrb
vSncFrvH+c0Wclb/Mp4IeZJHAolWCx/OTkhnDTnLfvJQ9zL0NwBopo6Cym+9
N+Lk8BsLrDdZ0uFa2fUCJT7WqRFeilKFJJ/IHvt+8eibWe2fZU8BgBvIxezt
SOjcLsXS1YN3t2egmEe5xCqo4qvPNUwR1KnX2Jm72YBLaDw2Mp9drhIdoR2Q
3u/JuJlka/1C0kIwTw/eejgw/O/U3Rd3pwJ8AP4sRMR/qCX7AuCsxeTVyBJ4
fWQr42NKl+onaHj9siF+SJintINEB9Y2ZiJDAfhMNytciVIOXxFATLv1DN7f
SOYpvzN67CHVS6fwWVXZh0DDkBB5gn+vk0mpvaOYW0iqdULZhLYCJDOaYWqf
oBC05X/jWbyeQunSluOE6rzLkuUfgkdAEQWUEUYGURBfKxcNwOyVPKUNy+8P
5MNA6JKjbfI9HrMZ8hgdDx6NxdMQ3ciaMsnR/2qRrVGZtTkYdJrdzsUot5Ln
gqlFxTVNM6qg/OP7GfhUrhf06yK05/vOkfofaM/eAOjR3UGYA50x7TR/89Kl
AXpoUwn4++pfPpqZCx40jKyr5mBeRS0FvLp8PgCzZXAYNEARy/VCOlyV54B8
+m+nWT5AdEHO5Xems1yzIz8YgxkwfQN9AxOYbizaNb34ld8Id5AEN7QwAyob
6zsPnlYtZpNIO2Y8StalMbJkeVcBYLQuZNhdtHVY3olsoMuX+71EpZtVKkNJ
QW7gsFXCTGPZ/RLUmFGYaAnGzSzP8uzyA9CLGtJilV2x0fink/sSzgo6Rja3
3qIH3CkTBCU9vDJ1EctHZhkEmzAbgdZvezhxY6wHg4XEgk8NAdynNVFS809b
1ikmBlHQPuk/nduCb1obQaqs2FJJm2KvmbETrpmChyzYsgLkNIty15QrZkQb
DKnEE1SXONUTkNgQnSx7t+RowcUXRMPilmFoDMQTPwAaSbcfjI24YJ1aCcl6
IPnvELhWXtr+CF5iIRKErY1lz3SYg1qPstjamvY27HBn4PTspFxmpnO8KsiN
B85OauhScqw9u6wEqSz2O87v1gip1QytYzuKRFPQPAnmPchsTYSAuKN5Wqn9
0Pg29vGj5q9d7zjp7tBQbBmQK2HFTPjB8LN8x15uyVRLz2wd0431M3x2/gCU
0mJoA/ZJn4qUZp5TOIkcfNMfav8i+tjb7vDRUvfAmkyyzXPHVvvzFbaQ3oQA
r3uCEVVWbVVdNedIEwcbq5HFavpvDZvPC5lgWSLp/Ox+0qXsOxm/KxsniYaS
6q/o11jN9veGdS7015OC3eZVHwhR7zTPZk2RW+6bQpiVhkPbvTtqEGgmiezn
wCKw7R/skKfeIkLa5T9W5HyU+ptP1lGCGF3UK47xkRpU6OWfRPK2XmdBSKWZ
LmdGwFk1GdEHo6qJO5VLzrFrZTIVej7JPt0aNUgXnSdzeLPjzSxzniQFtb33
SjfZyNfO1DlXTyDTDxoRQ9sEG+DODYQ0rknJUaTXAHoSbVTzQ6V2vdETEBZ2
kQb6zmxSEVrKwJBvrZ85JBzgdctnzbT4vnrb7VUKbIz3UEDCcGRebIGULaPH
lSQKRkh8nC/oilYBMph0MU3P3zCpEagQdNLDVUi3ZO86FNzFat+0jXtNKaNh
P5IYNMX7Urkns3+R2p3zjVte8yMBLO3Q/vavcZh3YEnBX+zMpedV78MyhbBs
SBVKdr1UQoNfRW+PRt4i/YqVa/DVf5BlmI4RXa8foHa2CwxCGI9RCrAxyZeT
z6KO5SRnvblmR4GEbgHDXBX6eJb523qfvlH5IMlJs5MYjgPHOynt2k7EmDQL
odqbsD9StAmOUlRcHNBpEubNQ5S4T4KojF+G0ohgd79OC+nswx1o9bVdPk5r
QS9fWwnWNJ8IV3PcsBZMQeK1JVbIu+vCjentau6eCD6UhfDjiOsZiOwzVHoR
v2GL4h+yyzuMn2roTyJfNxidGLp7rdTrpG2YopDWHJf5pGkcTU3kU82/L7n3
YtAwC/3/m0aJieFH6nMUFSMhf3JIoMwkgtiIKdlq0NranTUoX0xeNq9kV7vu
CcdaLRxvgyMeptYH6/EMH7joUbRWAFg0mHi+EPihhsJELnOF2CmPHm9UUZF1
MiSyYKjpEfl7s7P+QdWOYf6DtrhcTusQb/AYyvFzRKXXs59mkPpdcjPmY2Xr
nBh756p5nSw7F/q2HcNcrGTFUmJwMtDQsozCOUGf9X3tY8on3p150GCWAdA7
4vkAfbe+ZpinYSZbH8Q62Vx9wI/qLhwf1zt1cLUNgfTG21rYNMckdPG6NhF7
DAUGv3DVfWPQkUJYAfamLVPNJ4fe17m5sg0ivXOtPL3pKjaOZ97AZtH18s8Y
BNjlz9bQQjbEjP4wNYUWxD+8J2HuWTlKz28g4vaQVcklOTtqr8RX+KsTBBqy
D+cGHghV1WCREq+jYRP7h6GkK7Acizfc4yLiaHy6wLdZOtykElJT5QZ+3Mtd
laOjPdy6ji3xxndcHONlRI1WJtiMIREhvG5sjMjSbi4p75kltGLtk9Mpc5LE
wyW5O5LcVNeGunVWa7WIXAVAHwRmipjva2kTr1aRbirzWsxtbrToIQDw5u84
cSvnd+0W6BuEjuB5az15Is2a+n+G5cPZXJi0o7AkNctRA3YE3tWUB9PQh+LF
MMZ+s21elmVnOMFlKEh6BeGtsGWalHdBcpMZqwbqJLkPrLOZycWPFAhnRimg
V2gPFpqoIUtqU73QGpZ2/qvilbkjowZSX3cZgyoMZHjNiAaX4U5lTAXd+PmS
Zn64ptDD9h7x+/5YsRCnBeGE2Sym8t161tuQbpzx/X88ggrTC7NrHETIVzdb
Ghq1nxfkxdz9N4/7niMr+xSVLJSJFswsW+Wwybhkmus09z3xddNJK93H6xsR
OnSdBHyNRrXaOfEZo/i6m7lBZSWx1xp3mYcQOx6x656XdwTZOgUaHSd3a/iW
L0J1ODm/QTJJ4CAbt3Y4pcLzafCwjiM4ONyntbDKsYt6tDS87vp1gYNchGCj
bO7+HIhZKwQp3yfGSAir1JNTmDNO/XiYI2hwi2+7LCftUUn1QWHb1r52BE0w
MdJMLtbn6Q5/S+s50p0rGsH1mqmLBwOcez85jyqx1vrvPEcUF+TUtd9Q/c2z
icNpCVRzSwjJYjdN7CdyKXWIOtGojl/9A9gL8Ec6hSSoS7m1ZxAZyk18gWaB
mWtnG20IRm5rY1MSJpuV9umnUFaC91KQHT9x+fEQZkM1RUpkSjeJJvL5PIEh
6LcqxrFIZNSe4JcLLYtOEBWN4z6i1VJL6LiOO+X2/iGUdsds5a96WXd05BX/
M95JCNRjaxsxzkLwIStW+yAec3XwZM8VZli0grnZj0v7aC3rqsbZauYBBTVi
n3gZif0VnSHnp1OGYdftjUPmYmO9fdpWaXKwFmT00xky8jtEe7Cp9cuwJqeJ
L2TTgqJKgZbKBxmZqv3NhamvpvgSBJSWFlB8rtEPqrAeHP7yDakAs/hEo0LN
A3YhTf50slq65XJVs/bH34pQhwGo7Hxax7Zh2c0mJGlOU3fyPWXhUVZO+Wxs
ZCfxJ0W63Z+JoQFUifJ7orgKaVIW/gBlFzRc21JRqHN8wWIHZvM0EhTJ8y5d
tNcTjO5K8PCcfhgYmiCSzNKqNXvkW6uO5AMUVE5UrCpGKKVE3puZyPYECles
0JVB8sZKcIDVEhqX7jN3nTAY+rSPm8gqihbRMqU23o2MRDmE/0Fy2HMjDV71
1OXYb5NkP1hb7msEcHwSOHdwD0EgPDOfAzWz2EV2ZmNl/c6mpz1FGdQu3sTB
OUddGpe+mSw3nRliUawg7A7dx17uY9jrPK487AzC/ehe/1otGdvieSGtEv6Z
Mj4Pt5a6e/xROoQZhbEPjeGFa2dNL6dtgnIQudrpJETYqcPdsImrn/sDbGAm
507ZWAR01zM2p3DxdsgAYxGoeJsLg9nYqmQnTg/8kveqc0d8d2hy7WWb9X93
HnzqizK6hozmu3+frXFLphu3k2HyLXPKGPTpBdIO2yA6vWyqgcQsWJwoumJb
DZ161uCQIOEN9R3pe2DaFwvR90wUVQ2DPTziNgb/9NmcduI6ldrNK8mf/G1p
ml97TcUjWocWUIjRYpMNvFD9ItD6AjobvqNXBRC8chxbxNrGE59yC6OeK8rr
wJzPR2NM7J4j6WhQIptSeoHX6XNi8IPgZu4GYTygyRLJbAHvm2M1xA2AhiKN
3KFJGc7bPOe+lBqC7eQYAq+i1zRsxqhmb93vAYP5bWsMcveaRfp2Sx8CaeEy
L6xOOQSy/xXO46ZpIF+2L0KxHhu4V84WUP4gZMfbyeMRcsfEc0yoP19DTmQu
rbe1OqwE6u95+G3KBrZjEQU/lkHOh3nmeuvBBO3V8Strqch23hSLctEOvXkW
mOBP/1sVOayLJkHxstpxydaw54JbJHQVVMSgFZ6mH0khIIAeBa5yTqug0W+r
Pyu46W+Bm74ML6bGUrAX1x0lOU3pSNISUznGRoFi5g7bftAd6D8erGba+vhI
iTEqPUTYSMyMZv2QMOLeVB3jLezjaRQKPpdw5ChGbMezHxL/Z2cVHzFHMv7v
exF9au1Ohj8nJQOoS75eIqXH3GpyrUsa+KA9ubVmJRlKI9LNFHmCTNWHJ/mT
IsL6rMnwMUgETXXX6r0+FQs3G2VKPb63H9/O8jdUcDWPSdKIxJrSuATqLvqd
6ZOpaXbN7YZ09MuaqscbNTReYz1Zx2raYxuZCSQR/Q4lLmt3LtxWiFlS7RWt
nbq7KMVyPLAlyKNbJexAnFOR7S53OMBsj6xMmPmSdWVHkImX1MtXqfeaDzhu
YyK6niya2cojcNfgv/lRbxWqtBQELk8RQU8GHx3Gh0Dut6q65k9rjtofNmt3
b7PvgtXgiCJuQAmqYd9kz6LPELW5gf+mEjyqj4ZnmrNXcUk3MjWu4+J4TUmt
y1IXQM8znBhobmWkhE1tvvhca1Obou+iZFohYviS//V97KM8JXFn8/D+2X3Y
IZNS1vLvjQCB9H5QbZswDoo/KBy13V7OK93UzpjnDuUOyr/NYzGJqDx9Ond5
RdlbbUm8MW9wzMe3oW1DvCMpMIcu1uDq03cxNizmnROK0b6tl2GDM6KB7HmB
HHtd7bq0J6LOgrLvITunBKhshDGe++ugbMnLiRy9veUg0H+DZKfT4C6IWQlr
1sI3f34a6wt+qAfQ+q8D3VixW4W88p+FPgNeKMcA6ANltAWsQasx17AhWF75
79smgLL4GjqIf72O1kj/ygn63M6AM3We5WMgXm1NPcRp+Qgp9iLyhJKRqkLF
XVkyIYO6X6NEAOOphC+FblL2fujH/js5UnCYBqsBDBcPrFshYXreyYuhlfm3
tBMfAf77YH5b9tck9Atgymz9QWuPTJElW2z4VBXD8nLHp2iZymioa8hNS0hN
8YUaZlE0eAesjpnx51OM0Bxiosmvchhh1ugdy0qRaPWmxmnObqsIwwUaBTzv
pyhyNb6q/PepP+9IUoBRG80A3TkrE1G1C5hvj7hMFSAAPs2mxdF/13FGkTmq
rQky2BVEqMSRNy6K8zMgMfvZxY1dGHI6MDawyzaF5ELdNCJmr8WuK3Ipykpc
pZEIJvbAOopyqAcksznIcbOcxcbs31vITmU+DJKOuegArIPvNwUhYqp9TgsX
o2++W8a3cq+GU7jHpYJr29vPhZ88T1Nb/myKUUeD5FWS7FOkPo1fO+CcRZsz
MD57whDE4I8JsDlBboaAJqzC5tZQwl+DS9eLyBhDJXZhJC8IfKlbGNG1k1t4
bcOCCwt3WaApLNnAI0nzB0vZqAtPrcABmv38zqIgEh7P9HCWzEzuoCmn/hRW
pcOzt00zbABzP8Icr4nwaWTV5whY9lu1FRnLwF6VN8G3XR3pzRk/ar15rRsX
SNmH9cq+nzyEDAK5BXK+9kD7rQ29e5krs6weRx+VTlsD5C8+jPsTfanIn7Mx
aaRGWlMliXFU45KMMmk7Jxm0l6DV9fS0u3iqyQVS6NqyIvjmrILaxZkOSKDz
owj4SU1qjYHvYMayMS4VxSivUIfrTaiH4I1Yoib3wOh5SNSAHTWxaAb1Cd6W
uczBjDYKSaelNESVBVG7gvmlqtgQL6DJQ81po/5UfpsJsoCRWcfAxxMEiWdp
6WeRuwSsd7G74hnl/42YywAk31w+KsgIlPfb07Do5g0azaLFH7C5vsm5vSFY
IOHYSKwwWiHzcCytZ6zueb8yWwJ/lo8ClqZVWh4ak1EJqmwcXc2i7XdGwQa+
GBB/AfpWalY/8KmI5vrYaZy4QQBUS+vGJ9gY8h+t5zhBIffwUlXNyXD6HB0G
3vrdH5EsNkIiYDJIvBJINkCywQQBZwC4AqFyh7J8oSavP2TdzYiRV0J6jWXL
km3XMNcJLi6eJdShYUb5A5KS+P4eqjPvliGSIQBOHhbSV1V7wKs/doGuxei+
cjV2t0Oa8WlXc7COQqkE2nU3/VU4Y/+agO2vn83pPK1KSKzLb2MSoFgfD9oC
JlwIgKNsRzd3fYdsKWmntUiB34nkz9o5u5RLas4Kfq4PefXA1mvOujJtvbFa
YRWiOOmQkeLhGiH9SRUjaIaxD4xyY4fiTZEXGMelSBgElwlXSWMxw0Ry6dwX
dxqHOGpLzv0Tph7W7u4f0M1W3Jo+FzoxQuUQBZCtEnJiAR7GVU7WNTm6Kpt/
CUpMC9LI+QN06px9o/rC06DmMZm6BRRSKcOkiFDmT1/gmcUcvWfL4+kUWZL6
OxqDUIXWl48KVTyORbwPWfzk32uM/dEsnD6JNz93RpRxaEnMkuKZYmCzEOyK
5xSx/lhsfk3p1ua1en3fip9vIZCzlvoQzyhX4G7hDco5fiZrTe8ygPKpKn9y
vFHbR16YO8ENRZb4lyHXdG54Lf+4GKhMBCGBORw3GUMYUs0ePlo/iEEuxRKu
QSDxEBCF6VHnf6GsydGER2VjfEr7W+20D5fB6urYb/ro3QuKDOwrSriwztk+
WlfmFAAAs+ZQcNWNF7OB/SQrGt7mhwiAHF11USqur8R993ofPbdRsmzJp3wT
1fboWX27wOna+vWrpeNLXcDl3XXTdNNeHXxmTfg8BJcKFVHh6EebfI9MR1k/
fKhGtOk6aSnewyTDcK7/L3NaUh5XWDrs0nmdSiD16cxgAHeJXO1+N7StmdHT
P4qr3buLPX3UsFrYIQd1kKbu0YG3tCoYuQ9X79c5jD+EMb09IozbrZILK6HN
5DlPFox/mAIlBJKSJ2hOYOmkNUFRv+crx+xRYrgyjFDSL4fub4XJxrHIQRFq
zFjXGN/5LMl5T2hU6Bm4aDQecXFaIAfLegm324i9A4E/edFHOiy+VNeQ4x85
TMIvBKJbhbhJTmIInYyAMKTPltL8vtE2BL2ZHgXSzOKzfsn8UvVrnLb9UGP1
ijEKzP3rId49BuhcO5DMnvnKe7kM96MTynkL+cC2w3k4ifGy8kL25jWid4ZI
xsQrKkq8ejLxcIMnqC5d5DryeIAV49yO2oZ4Sbho/ekvEMGsO4+2Id6u4fmu
6lBBRaX5D8YkF4Q/aY4FPXKmsQG/XwZw+flP3d9L3JdKZIGFzdybfxdYsgMZ
nkGpHCVTmIC14qQg/tg7ukoOxP8ku7vnw8vr3p6MztYPziB8gz3aO/f4jxXC
4emY0GsNOMEsf0xp++5QxojPSx/SZxyoX1wYNABQCh3bBb9LdzmUiBiYM6eW
G3I4haYqKU0iGj5S40nneiKDOebko+op05VvmAV16pvB5zjWMN4WH4AAWVmr
PSztoxTCOQWsqCyzSl6MU/5y9upXWheg61akiBcHuqPvDtHiK/ku1kQmhzP1
1B11hLf0hjnkHzF/Ia/O2+1PjKz3dF5GiubMZmV4k8HNLxZ5IP3qwpKXUju4
OeMvzxjqW5obtz3pS9qm7JOF8XtjEhIczszL2GTnHmMtnbH8p8i+L38DGrX5
x68OGkLkCVVDiTdRKy9hBvGcB0+clb89Mi9Nm2lJo8X/BFhgiRib4ipHJbyt
fRN0uCRADmV2iRxg+wlOpuX8fjP1cUAxIQjdgiBSad2/yczOQg9MD2/L5ySV
yOOAA0n1Y0WA7Vwph8jskuqKWVZIKiBwkCRmsldzQ8CbKsRZywWFbRSO76Qk
iUJ3VW9CKBsyxBkXRukI8vjh7wAlaqI8785LEiln3UbUUlXBMAC0KEfvwEvd
09q+AzIq5WMzk2WAZrDcQJAc4zcrnBRuJ3koXh5qzP0fBgM9KhwOAfhZ3V4r
j/J9eKlNv28Zv9jHPumAMd5PFpt1V6Moprj/mnvCRjTlF1iLeM0AOfUO+4De
xCFcs4NhebgiR1S9q30IAtYZnnu2ywJlw3cY8aLYuozxsu6EgYMGC3ISAiQM
ZRqxS0jxFlq9faPtEPdKC0elBEEcjFRQNwbutbnXSaYUmvUpjxZtOhUosnkj
Zv3C80V16UO7zEoUWFfpiicKRJ7YPT8adBuelzfA4+F2d3zLIWfeA2BV0klr
j+QKVmGSj+NYhWS4ZhQjDJkXx8Tqqf1Svyn23TS2987nEeUesi15RSnjiSU4
DpNAP3P3TzE9ruyyZ6hTMjv1YS1DfYv5Is99uNTx7juOQXkOySsYRxpSsAER
TimBlDH7uwQmhbBMC0dRVts4IuWSqGX4D2BGMuRdZnXCaQ4G2sbo+b74tnGv
FYEwLh+tFkJA8QNjKmfLxd4MbwrAub0TnsacQbPhMeAdh0n1YsddHEquEn3k
BCLbo067GqcrfMElfAEWbnXWhtMjybsjBv4gl3KZjSdUM6tGoFQvLi9Wmosk
4MCTvQdaZttFmPX9bzfjnoxc0dECiVzBeMYuAFkj1SEeVVc3o87W8wDka4HP
dgPloLp1sFdwWpvNRHFWi6Ng76v+V73YwgvbQ35vSoXI0kJMpIYQZnvOaTL2
S9aIywlXM4R4ObmMBaPPUqAQ0oU6cy1OO8/jiEtKR6sFzv7u9FjqKh2lSd8t
PGiodWGiVxt6snX1kx7ZKH6/RQxYRfNpIH79N9cILj2ZsOve72xGZbh3WiBV
QcZRvm4a3M+kwiSfbgKtvIiolIoU8HLPCQ2WeZNyp+h5ZO7ovVqEFCuIizHa
hUfJzxUs8ZOYLkQNXRiKHMLUPYriOaXd4RKupU/GbcqUFn50LgG5+lHvTXxT
RyK1NwgpfdJJH4cYNaI1Ti4q0kaMBQSbQY9M6hTpq5Fd/69VWDgcJFefvtL1
DTB9J7m929ABabN0dj2h5BC17DscqqhOWUccUuUXyefi+1EWkqklXb3/tJ4+
P8IdBWFEF00Ya1Mrzj3Z8Vu3PjfVh5klziPYry4mAMpcWdkG22Bltc1MJ/3U
z2Z35RyUPPJLilBkOnVCIfexHC6h7zQTACUexTcafjxSdamWhPE9zZ0J+aFc
gxMbly2TfYtudALfnSw+Otwc7/Bgk6rLIq/8+wdxULq4zvo7L5FK+G9ztlKY
ORJCPxODEONV/xB0Zpn16YmuwtoDp4E7RbHcL9WFnkfUF+/29Aqo8ixOhbJS
h7/YwjaWSG/UWsXhqWDzDL0epFX4UNfIbfetgqWT4ILSZJ6Oiv+OIvr2LVar
B790CcV6Be0OmkeOZ35pGdyC8gSPGZ/R3dY0LeKevud6igvMHIaYLLYXVEYN
WWNmBI22uYHwo4wc0kjKaejnLziidkyaPLSib8j+P3OwmXa0svNpMvqMUmX4
PBo1Z54DvUTtZ4R1+DX5WQwIP9+et/uOzN8DRFYcXg+lFgtWKba4M/mnwGxt
HNpFpCcAh8qprOd6ZyKGegfKDacVxtDC5kKEXxeGTHF86txisCrb5ewD+Ro7
gkHt4/Dqxzj2tMt1UgLRlTme2tvkjsGZmSy7O7QpfR2SLL9xgMUb2RMvJphK
DxXnX1I6Xaa17CNPOH1A57flf8bOXgttoNjcwSi4c/JBJIRY5AY6HQNPHSHC
ysS0qQk/XFiBWGcD0zkEA7fLEaNK0pLuWpYVhgh0TCL55TGhdVnEf1n0/0ej
oeuTPFUdAJilPbpiQSXRefUEX8txL+Nx5QS06W8Xe7UYmOqo/w8Yspqc5Uae
QWgAPPNMacs+tMZ5goYS0FC10PJ3ngRaV1YWgr4rGUxztMNBzhl3yPD64yyr
ltUqNmrZUt8K0n3JhIARrzBHB9Ta6i2CR1pvjV6MgsjxT79Rh5bwXxfamnql
4FM+nkUuR9S2raCIDePdeOHVfd3Azk8ZmgyFIzyHTbDA0c6TuNDYc/YiWUku
ii6R3+782NOzXjU/3E7Wbr/qu92ySEkLuhqsAbhJbRdGLj6nZ1MXyi3PdsDU
U6yO2BxDLllfln2FHmPJVQgU/NwBrrwWTfcNAGZVAHUqkkkKeiOfUcoTZHh2
yqfVp1ASk5y+gI8Ib/qmlNB1Zxoj9q9znwlRwBF0j8E+J/fXvSDklz6I7QrY
QEzjzGxwElssgmUuhxG9TzxCVwRUjXi16NfrrCqxlWe+MvLDEOauQUGkOfz9
Wtq7bRhcjSwZdBc5QFAIHJ+9oI4jVzIsE1c5jxzW/GdlVOp4AGQRAN6VMcMq
BEdEsnaX+naL++qV33vsdAdIK6PQ9wiqTIBP4ALq7kgQnNI+uqW5K/fm4o2L
ec8m7HYyPt9Ofh7Z5xVHRHkM+q0b0/dMMIfMR6g9SGyU7rvAnWFKXGOrFX52
u3eZTACix7TcTnYnClcxjvfwNgTayCL65NSh1KWMW1LsisJIGfJQt8QfdHPg
YB4bl/QaGD9ApyFYf6tiFgmThTW92csLK2rDPO6Dmn9y7vlH+qga5ho5GL3s
qA/ALWbX+oNt3eugYLQM5wLVY+sVToFlJtAquE+XwrY3sNLmfona1DAU4hOR
o/eXkx7q4S7RlOdpucYyNAXwvhjSpK0yjMveWXfz1zac3MW/HYz2J/6Sg+hF
WTKxRB/wqIZnsHjn9RhDStnfOHiceG+g1mKc3Szw/AKj8lhKXuR4wWoAvI7M
uyRmkhgMc4uJ+BvQY1iwPZveCNsU1nOGvoWNX+zzcrgl/IY/Za2Y/MtM/G8y
IFDPKqsIzDiX1YqenxT2N7ktMj55ZIvXCJYu4B954X813c+5go9+cY5fQYWc
XQM8hzkwR6RYI9Mv51TZap+ubDtkQ1Kl+sgBHNhfuAbqE5ur4hC3kC1+CJTi
dFmoSa2mJrmnrflgo63m26KVyrgdAxfM7X4Sajzx51itXYZPkZBpLGy1oinl
NsMXHw30/YXNwlKfnfxXKckeIEhb4ZxioNwIUArgxVVzFBasM7PhRZK4mOJE
rGFKL+jw0uBfjk17DE8OxPOeuYJd4ctCeCWOOhIx1PFtVIoptpezIERIGOB7
w4uRV70H8d80u9URSLMKaBzdZ1CIP+UwXU3D8JEoUAWsrSb1d9uLvluWZJ8F
wWxkEzlFRbun8xlmJ4JB0J/CdvvS0YKHxofdK0ATSOPLf8lW3hv7ji+ru7uS
mpN6NycVI6+f8xP2X/87jX32k8vmXZ8IVmrHGtGFWzwnjFjtVO8EFv6alM9U
BZ9BX1MZoclvO6Iok4RAkWHObeiWvhjtSSBnfNGT7qsT8j+PS8kd+4JYg3lb
qM6bMmv7U9PkEbh4IqYryRgcm9s/zjla6KLjRYU2HLLoobhLI5EpKSYKo2YR
TKABpCYGvzapo9sEF/oBGGj6PpNODrUjDSSvSXrNKIYhbRtFlTSiF5lWGC5O
FPSeuIyVdruITsyS9I++rPeN8fv1GCJgZAuafGUeCZWXg61WnDKu9I0iG5F0
fTumGEvUP4CGpqpwoedHwU+7X3+we+b43SIjFhFtMohNsM2pFe1UZsX4R0DX
7WUFKVoD/rAu5OTvr6a9Ucwsktg9jTAen9WbyH6R7O/JURrOEFLdqUBl+ebu
bzM3o/T5HvKE1TF9p07akWEuKzEHaXZ4rLOG6xAfc9ztMK6sLkqijzqfj8rf
p0OpLWdcsXjGjhwDRwAC1PLAIrBMvUZgA48Faqa0af60StVv1dVys+EzzVMt
/vRDNiUMp+KLprHKQsGwQEnBvfh4OZR3Wdr80MDRxucRBESavjsqYwUfYeF6
lccWuCYe+Q7sHUF6qVvAXEFzSgiV+OtONRkfMkNh6YIlJ39HFqT8NgzwtsO8
LX/FrH01/K8FJSIh6y7NVBRSSTRQbbz2mVYoyvq4IEG3OpwLMHrQ8iFahYOf
F8tTsWu8gMeYxwxdQRrR0ni33X/WBHALhKZB88l+YTpvKP/VnVSt84lk8s7m
mmY/9p4iN4WWQSMUPR4iyXANHG/7IgCeL8C+eCl7EVMcFQ/m64L4VMqSHHyM
KQis7M8EVOxrmiMOzOwSCqK8t+JHQjdQlo5bQifJ4sSV0BIezVTDgrOfo7Oe
iUM4ZLdPyvWSFZqQgNOxA5Mjz8CfK0Q5sEY3nF6cS421caCx9EUOUCnDdKgB
t2Mvjbw2xS8CwV8YoFp/kitI//Pvfiw0mMYkTnIqzZwODLijvE5WIY1E6ixY
sdbIz8bMYek9gqwvUfJRy0lHMWXDgYL+eh89SvNVwdFoxIMcJ2M124l51gVs
4HHEJxxvj0fSFVhmgzfVXdgU65zi7QIh8OJWl1JGIBnpgPud+6ApypotVKMs
UWKJvceFpT6QtssM+lauRaPYosoK3aIlE75smaGt3A64bvtLBCmxl3k6YV/7
OsiwlPWETbWtRBPL4Wlt6sxBg2F12pt7QL9uvBemrN+x5KxsAzGb/XyeKK/n
NdwN9AptnjcLXkQGFQZrvOKAB9fbJd5Xro0gDp86/d+Ua6HywrUghnYcEswS
yZ0v0eSkOUbOmledaf4S/o+lR7pBW3sMHX+F72PnhR5RH1+qtoc1poEhz6uX
KtX6i2eFAniBj5MO5R2zzkpERGQ/wvDpAu9P/zh39WFBKay5bAaclmt0dFGX
MOf2B7Tzvx4zv2rqMBbmOkckCkvqCmb/q/VA0kcgcqLmmHuv5puCNTfw2rzR
bj/SY89ZBZEq27cODkl5Wc1S6ADSqhzlyOILtd5puamVW4kzzkZAJQ391ddn
iaMAYjV9uccrTtvPgPwBAftaE2aG7z2+AuWOL0GwH5GJR/E/Tz2RhOlBlCR4
A1fkG75kwvWcx3s9D0wbxN0bcu36PXxsWsXtWwttcJoGEJQRHYYqIjatOjr8
K4RTBiOG8Gr8ZtEA5Egz1omCdT3E3XnXb3ZHqE9CqEaShDqc+CYCJ7oKE6B4
zpMhAItuDSnefH6Z8jwQlF/WqT0MrChftPZJh3aQe3sNdC7uahdKU8bW6V6m
YjQg7wXrz7IfZ70gP6CqhXIrVOAGIoN52uftjEAgbSnCFn/UTs71YM3v1kDH
Jfhb/pDCVVDgv98p8MuIjmi2CrHJN5G1KjVqKk0iitUwSGnWyUC53v7RIpgT
BPTii8SrGpZ2Yq+OfIH3ihNI2lWWtZn0s4YYwl9BFAN3qSxVTy/p4EEspx/b
H5BZm2SbPJqiyI8E2L4/Uzsfx/6hbfHaj+EZPd+K/5PRFH08zDAmTfqaqTcw
POzw5aNS+wSvdCDIdJiU5Jfj1Y6VY6UeZU8HgILbYUj+7Rzos/rH7Bh0Zq6n
1PE7CZa5tb4nvNzPfIwMTDRkgp3+V1LNXUG9p+gre2njr944LxmubHMxWnws
jKw/6hwEifzMxQkYkxupUbVGbRqQKNrve69bQW/Au74bYBAyzZsnLR9qE6fF
lJ242KERDQRW5FyWmAa9jTWcqog3JO6acqw/92kTFjf1rsCT7/DmOn1gb0W9
x4bfXdR68Sa3Qfxll1q/DUSu5/TtrpdyKPwZg4pYzQuDckf+cWc7vsMw2HVQ
6S/6mNSDxyiSuJw65v1wF68SU0xN0opyQJxRSv45PFBArwABMVRFWez/gcKP
+KoS4HHm3XB4D77xkdzx8tFYXET/iJVCa/lRc9F3KNoaetR8L9qSyPGC2CCq
m9lBVPqwG1mo4XgOkjUbKDKuTbswslIbsW7nBCX6uvNzCuwDyvOtpTrc6gc+
9GQideiticcDML99egPX4/MvTw2CPqCVKUnvzxfX7iGMHOtU+bYUEK2DBUPI
5WmyyqYACr9GnFrsrD9G8FFEaa+McAcmXPCzJv3nD/rudmizrOa6vEaVwDGk
qzS0BQJ9vjRdhyAQUb/5wRwfLJ2RcZAK5IFS5HMhYcJAGtmkzt0jEBvkzEaw
bSPbhySyjiAY42dGEJcmc0IGldlpsFU2Nbc6P+UA432LmIQuDPSoZBlskSSC
AJLMfBsXoeiSQsY0Q/7xhldXUQmMDYGQkqxszLIH2x0A8rnYYdbkpmD43Ijv
7bn+COtAy40HeARwJRfRt9jZPJiA0npLjkba8M6teD96FyP/Q9fSJpzQ7otJ
nQ2jFXwWX8N3Ld0Axlrqq9hVh3pkzoZnkAnhQ4PQQix8/BAiVwGxrqCvWfY0
KJt5scxu3iOiisIeByLQmYYzaYl139sLRpp2Zz1umrqpKdT7LOQDno+AnZ21
x8D5lIAIDcuzzrSCHvwDw7zZ7TQ4rfKREWl56+3M2GNeL8Qxv1dbrTAnHCkm
yC89W8tyPCDWtaAmxFYhzcpAFCKsudWytIKOYvBPJ2JRuLBlD+NsXix+UzFV
CyQqzQ+3SacxdEt03oWxa4tqKyMNyiPBkVw/BaI9ZoF4Uru+15NEd/NqXKkn
t1NB4sSAPCdYZLHUFmEk/hIATJdw/NnQ91N7KkSo742bAQRmieNhXH6+Mn/8
FdMpnHdevAGzQGeZ+pXASbYytH224MFAdWYB9aOyq9LaJEavGAo/sECkMBwI
LrLzY+VM0zfecfnOkbeIuRkeAYYobRkNys95yPUccEoLwiiphXOq3RJibI2B
gR7LT1tK6mdpgwczUjlmlVQ7SIeFgfEDppnU4Qicmd3GYGkrdA/DHEf/pJHQ
uAyFQAX0UydHhpKVwokUMbF08dk+CW675N0fT8RxflyXRujDjvjF9tsB+Z8L
SPCe5sjfoprAdERRLfqI8Vt9USL0e/3nw576eMk+Qxuwjbb3sNIOh/HRwO39
/K5DIRNWKDWw7oT3TwrFlq4vap/qZ+MS0WiTA51pW1I/n3cxxWfOqHBBdfc9
l0lF67m7n+4mfmYOjN7ZGq64b11Jbfah7gUG+llqcpDnQuFOZ8H0F2pn1eph
nJy4nvn6XSlqp7hZDPHt6mYUbI63l0ye0pL6os6WyBhI920IS5o5DkE5WD0D
VnonYdDmGA7jIsukg24GBIYIgcltCAuOwpH07ykcL+JzV1d6CQc8ksBWSr5E
iw+nOFtZE/Fc5yIQ4TVUzssIMdcMXiA4APW8cxDtjEauI0Nq3AJ+3v5ueUsk
WC4uA5n48dgWd4ykWWZjsxVsj2uJnxecbCUrnXFl827CzwzrrI3OkIQw9+Jb
9rw8XsMwmokVNdTKCKg+69So+l/8AwM/+p+7ZWsgpogwFi0Tjel7yH+Y/wyT
zQkK9JhedKV1HPuCydba0GUsU8clqzDhudE2NozHxfB7B2zua4AXMhICRjqj
WdjKhjGFMwZE7357APG+z9qIiRYrk5A2itQujwNRSpFEWiA4KEqRY0J87eHt
ujCb5XPDIO9/oj0SzWlvRQwhZ31yOKNjqBuKQviys7LlL0FhW2jvmsGwx7eP
N95MKKu+jcG4yWPQ9eQMEK4qlZ0OwqYwnFEE3WnJ6+Or2pCOw/L90d67yxCN
DuUUDPKiUeK3mnB6QHrC0OxRe2XBuMK2z7ZyNQXkLVO1rppVckLmg1ZZ4TAf
u/qAjsnO4olQiiioyRCYGWMKK8jXS1IYuACm6NtAA+Ie+nJ7pnYyEBY0DEtP
AJ4uHeK/Lp6yDrJsQOeL96hAqqBnHwEGis3AJIVJSmy3HRoIT2soOf9Ad3T7
mqiKfbOdTWhnj2S2KFe0LqCagYIBffCVOnyED9QKQ5QMCcP4tmSX9lM67gqb
SxkYnSd+A7F1DoAgBng72EoMswWAR//Zb28oYxovOxFSe8JZ+01cNMDiYQ38
G5myNdqSJ8d1bhqwkjROHS2uHZfpaIMh43b4jnRNyw9+WE6D6KBEBogIersP
dXobCNaVn0D+kWkymT+N4Zn1mqGC1fpuzVkPba6A2LgpnV1ZG2e3/wrErqkS
zB4SwwVDLvadhlaD4UXmHwiZdXVBpPd0A8svglwPH0P7wRgwaHFOvKDCDhae
9kiUDRUd+AcrPZoKqYGTHs/tVUvGxzxsdlj19uBRHPgfgFStU1Pg6mmSonWU
OpQ4uo3yPXofhNYcM8wsc3wtiwVQ2g/6P86rJgze10iKxO5HGikyQnMMN6iq
gHa2ddBo/vPyPosefUG5afDZOR/ehHPwWu10IAKuThIZU/94Xd2oexCybCHZ
bNEC2cvkMcXifk9PgXe4v3eLRDKc6DH6mf7je+7vS63KvmA7rnJ28H34fqni
H6SSK6RJt46Ng4jyghiq8LLSNzX3SjPu2chZxr7gB2aFPkdl4i9KMM7GJd2O
Nvrcu3hNpQQqd91g6Jc5oIe8H/RIN6NlKmvRmU67dnP/PvFUo2Jx31OCzrnt
byzE/QFv1FjG4a8YrZVQRfRtPX/TAYhdEK0wQpTjhowAnTbZSoFJoihcVTkv
gK+etCnSgrxUlIE55iRgbacvtjW18mFFov86e09s3kN/Z8PvljUhwqkrdW1Y
kGMHopFYBecMOrXehIFgsxb/HeN6hIFA64pvm9SV7DBkwkG4+8u4PbaV+UEW
J+cfKqjOrWwiscwoX0OTFX579dvJ2mT2Gxohs/F3SJV8O0rLQuromKj86B5b
F1dBlBqiGLC6GRD2qOxOAlKeK1Xs97M7ovdZW4zEO7PVEnFHty2/TFf7+O1z
5Az22QQTeU/uCVJd5jdku7DAXK1Xug2nhssejTOoZsc4bPyxMwLAbUmxAWcb
Ftj3Cpkm0HfWIu/q4zgYa53BPlZGuhKgKUp5YL+yWG1HRotLShBLNePA4XsD
TtnleA4s3R9xosc4JkgZMtktL1rtMlzp2UMOx9Jqb785zY17NA/hGaug1Bu5
PPe9xE2xiVPOyPzFPJaB6ielCGlIT6lnFgIaQ8VsVoK3u8beZBD41TYpVUk8
tdFGVwWVxBLF8mhNiJSysgB984tIOloeGzdymhBApWL8RshE8ukxU1o5MwiK
H2Bfdqz+EMPvk++GA/vyBUuUCvCmxCdWLYghuHA3ez56Ugj7sXEndaDqSrKR
fbZELvi6mqBUHmn91ZXZNw0SdJwyKy9nE4QViFnsQ5WFIVt06/riOwa5lbX7
pA5eVj/P9fu3J5paDZ2vD9oawqNbYjBbjdHTQOl4jL4w4SD70JJkZ1XkLeVr
skUs5hdnmBppBF7Jc+zUKxkxIHCVUuiV9Fjt/uvrlEug5Awn/BqL2oQdTUF4
yhxN2pGhf6GCWmQx5dgNMZaei10W2paFe1RVEwXzeWhxUqJYWjE9ipiG6IJm
E3APig5jUEBj1DecNnz1Z7mVmZ4unGIowECyB12imjkQGuyZP832Kmia7c7G
YkSm84+KkJMrNMG0Vm5xbpEpyxHJ5uyhS5BMpbuniHQtrZaQObXv0Fdcjr7D
QZX+zrQ10hva7qR12Vw4SM9fnElK78P0Z9Qwqau03dt+G+0293pX/Oc2+PQW
aT6JDKm7LCEBkHJks/izWtflWB2nIUhXez0tXazf8P/HjcLRc8uT1dr7n7Rs
Tnivd4QQjkSpmG+iCULA8Fd8ScKC/j+/o3uctbFwRK63wHH8QMRiLLeYYIwv
B/SAOMAIggi+zQExnFQ/20g/ItdSpYqLygTwgT0br25rXeQwvBLprKXznXjL
U5BL2t2+RovDojXIONETPPYf6FXkUPYwuxjUtrO9KmI3vKvn8NLa2mj9wmPV
0dnhUbmBW3kqVghvumXX+6iiYkDGsUrWbREFvyAesSBgyN6v8wm2GzrMGWdt
TPX6WaPtfAAQXBEmoMcVGDPO8EjWLJ1OhvYIyzMTJXx7zOoJc2PhSxVvtCf5
Zt8djd5t/g55p30YI2pCF0RCHeukhZdpfdEjxhV7mvJ8nNUY64lYh78D5byc
VLmKTgjaGqXGkQQeul56aYTkI4EinTdw67ShGxENChSmSEtMpDb6Jp9ewckW
hjkkWSdwqiYsPmwe8UwB0fay5CApcUYD5BANQuobuaYpMlcDMXZbGFZUUrHE
J6f0Ub5J2NQ3GWwN9Gbz/RtK36nRr10JRAq7P0IqvcoWHuxZkdZMoKS0NvcJ
xYVKT57tT77KzRlcqRQcrrO5/x9bQICylj8OJrfcxom0pumrUCifQurTXqM8
Rn4FM8Rjn4QpnxGEgH9e0cilk/AO5UXW9EKFCULssl0qTXXv7FbYlAidAlue
z8pjumhlkhGpFneZUUgIWPKHJ6UsGL7FlV954w/S+ym4WNMk5qZgZSbGnndV
oEdDj09g3tjIhjA9qrh19DihaPAv9y0GeHpXVIgLP2jz5VthYRynVRm86/0g
ANoldjlSxJnDyKpdsMTRZW4C6AWAg5bA/djun+fNtS5TqlXjmnU8JlGrVbL3
R5cEacpVFmap2LWkLL9B12f+dT5N1Fwrxdi51jByp5x+4tL3sR5wNXSFQLUd
7Dke7c0K+gBxtUGroXiVFbyU9BhhsAyzPC//nrAvXQrqvmtnFg8mCmIsC7Rq
+xtUj6IuK8EirFTO1iR4OGN150xFPLN75m8q7rxLkHbMoFY1mHzpx/xNKOZO
9+HguuPpCI4hxn36/OwloiYBYSf49tWBaCpyBWJWkKgi8uk2nGGxNSp1GkEQ
Liw/H2EtbUHzWxpopMB+1ay3Q+JCgK9yHmlvjUgnytx2o7NSMo3eyFlpofFD
GpGfUxalR21cLU7H1zMW5cC3dNNV2wp5JCz45w5dEOiC0NoLvhMlwIGJX3YT
BB1CJ9ikKa4vJX3rLN2wY05Dn+04lBOWwet/RpOSFFySYC5PAe7Txz07OC01
SkMZ71cm16GjBc7OzBeGA/1pnun3gTIqiwD0nuYaCCYTt5Ubew4j/yjWGyvS
PEkJuEX5Are+g86oZcTISFQfjKCVFokIJrzvZg/wEnCpyPwVogzX0i5jkgE9
cwBTc2DwxZLZ3kuyGITYXv3h+nQYGhwaAPNESwkIvbD4eygEK4V3UmSPN5kr
JVrd2ffvIjEFEYn5AkMc+vaLnKrqqvpK/V9SXFcUvwD/1wHcg37CgcA4/0p4
/53JitTDHcO1pazZ/pBt6RKsNjdu1HbN5la1azyo7/TOt8zcBhSpOuCQOOpt
ltysojcCRWDglFxOFdFWJX7aPKdIXmc9HrQYG94GUQhAkifacsI2EpRzs5eb
FcGKrNgZR1167JBxio7o3sxRI3vkQS20GyCUoqEWXseRql6uNzN5oUBivmxU
VgDCyXhYRY8i8w5dNZ1db6BUUYHhDDT8V7ZZpLaLBclgA1Ojg0wxlElQ6h0n
itPpVv0Wd0v7HAc9dizG9boab4Fm6Wz9EnqEqBLqkLktXR36ndU4cK2UEha8
bYEYQf/CrdP8Nz6ThsCXer9PBQ6NoVxXW/OVY0JYp0XV/ls/MCMyFGgy6EPL
w2p+8yswXbblUsLemPVgWsD9ga/SmLy5RS1UsSTrItNVJFQwEWEivGpEXzMQ
enolTw5o46ih3BjS3aB6XQ52waKQjZQBajUr9ZVuR1II5Pn5bCMd3Ox3Vs1h
c9NOYoKcvnP8Gyfvl2F5f4mPKYKsHJAyQQxlFazZcsBkEnWVDtqXHajpX2fZ
18c4/iyorxSRLMf8/0OfcX/i7Y5VU1JsiMQEn4uTc66dxeLhJGFmxId1tn/6
g8EqhDh/dm28dQvilHD7MGRKlWbiEyx/PSPQfjxLDH/LJUJYuIW2XwGJU6a0
cDhLGXhE7W0qnCNuhMDDCCwl//yeMmAHe19UNoYrX7ROknKs6b8mam3mx0iU
gynjHOgDzsHCUP+tyCFL0S2YxMbWjUPjYLA6biyVH2aBnqz6/oqPrhhY6qsk
ZnoFHf/Rlc4QMCcm9m0r5WXbeP8bUb65iUtD1M74iAAm2Ci71NOyTygmUsG4
JA2jkzidBHjKFZxn0SrjprLmeBO3WF2opfBt8IZQbZjRwRSR4d+8t12qTmuj
VYZlShI+gDj6Z9N/s0wc4qjgSQQ+yLF7aqbm3xzo/C8+qcQCtthlvtn4+3Aa
8MpCTHtR1HwFIwmv8JCecvxx9LqzcQ7M+BttyjQU6Q3itypXvNOBoS45v5Ym
aqR8MRt/tQG4st1BMXsNnDieInstZGswl+xK3zfcw8pt/bdLn/0X7twSjXgG
2eq7dH/tiyCdo94vfRvJp5QTOPw6kMpEBzjKtx3uvxE8hW43F0Wk66akjXn6
CwWQ/eYxbH7j1CM0z482BGWI+wh4D+YiycZk8TxQuGKjmP2Eg4qvH89YOzE9
5JML8SNq8W78uuIiRRnYjwl0t/eqvjKLXuKc01BUIa6LcKIgPyTZDUxtQ/Cg
fSXvZRW/RSEHOfZbM4Pw7wYLJ+se0KdGAbcBrBa/dWBZnaE2IvwCn3PGw19W
P6M24xIUcxoozDZCraW4VHXN8lO9qdfxeOAqZ8Zzj5gNcNiEZfajlPygCzdp
Adcc4ueiaGxCsQWUz4oOJDnlJC3POUMwttqzpcgHgtuykU5/xWliSm+wCW8n
UsjpVXlm6+YK7+3ZN5LVduq4nAdxIiJGZBAABa0ket9XiHhbwVV08+Lkmmmv
YRTvH5sKIBFyai5tQC4/UEseC5ojE3seqbBBUKulfl2AiOa0hNKKeIFhRasa
LJ9esCAadhubCxbCF11tREJrVe9W8CoYQRlhPQ7IVP2Cx3qkBePOz1eygpj+
2hcNIJUzHXQj96FP8ISVmrMx3w6puC4UdLL0NEbhCb5DKLdlK3qaUhOoZqCv
izpgmfCDNikOjm6JEGlzTFkShaR2l0vPigxDxcbHpgGr3qvOxqt7V9Y8w+FK
GTIL/TY8/xwNHgCbJoOr39NwLozhMqzSdnnMrAT6MkZ7fHMeE0x1zLmHzWsf
r/LAFu1hgr+pi0qTb7zWLlQxeVZOepksiE16yOAbukPEzsP74WKgx/iQvtxU
r0dX0Q19eiz6EPHkZGCDtpxQUbxCxfWLXGgwnd4KfaUymbUqgXktnnDo2/P0
8sLptX3fhU2EoHbqUWKfG/P6BZEeRPyOYG1gA6jhiZHHytosc5sLDL0Qi1UK
g2Gb/5kHP8kLz2sGY5Ax1Dut5mpfBHK7/BkXY2lnrJ4wrunukwu2d75817JO
rOJisc8YZmeqLV2Y8yKBz6dLIipZB2JgK9Pwje1+zh/PGyuVlmGIFDqqsIJ/
++F++kwOW+slVCK5MpaSpb32Rb6iiYOva5XqZEF7cdStDIT9oX17t4HhMAay
iBC79o3K5Y85PaPD+vNcmQ2fJU5OjcFzRLRBn1YQHXlFY9PhFpW7ZkSY67SP
VFTkbUUAr1Sidlt8BPRPTf2nW9D0QmeTz8Q8OOiAwNTCCZv2zNi4zBbKQ93D
5NkxwJkxUmDTkgATCsKmCV8fCxpfo37JwjGqm4zWeh+jFBpIZdEVjNfckC09
ipR5eGVj36YwJm/BjHbunjp1f+Xt2Q4OW+shLpF8M40MaWiPIL9dWSwaSUlG
TZnlxGALPqqfUO6YqV8M/7T7bXL03TFYWAZ+vQfjZzhj5beqZ4wlE8b9npS7
r4TkfjhkZxJgktqiWSFgsjKANZVLInflG9Xx3OOahYtNaBEsFMIjQhCWw7Md
rk+z5qBn2tjaeUGpfwmrtYhq8WthFhwqOCSSSgAEYLV5h+v9se9MaqRmFF39
t+cULHRlfgQ50PvAYd/QRHgJOF70dbu+RjOpgI6qG6cy7FahRJ2p6x9FNH8W
7SJtgOEld48rIH0QOXM23X7Sgsq7O+28OPI6n9nN5drQN7ZA5rn00kvEVfww
xp5/uOfEJKSZuLmhYMZmAteR1OIGLp4/dNNHQZ5YUqRmIvcK3qPd3rFaA7x0
lGslfngBKaxuk4k2XuMfONUFI45TB5m3LJiI/oXuvvyslL6zl2jtCqp/9FAj
DRlBxQE9lnGivftcsQ2lZ/6CmRNQ91+Go+msrS+CPPG6rRu/r7UtCGOfIqzF
Z6JhHSfxkOzZS/1o6jAjw+MYoC44wC5a003iBBrzGCUxWRh2cTxxRDszGy2N
cxPMhEGaRexH+zQJcikWiOTidVbxiflp3pTrTHxuGm13dl7oBceDOpW0Strg
Ozkt8XjPcZrsJqA6QdHhImK/AE9ha+6z56fLIKi/VxoILTLFnJbEiRY80UwP
NUkRebCH3sI8k4KGgyZWjapMjYxuvjSi3R0zONbequTCr0/uMTtxvbS+gBXe
AomuTTXNrI1NVYDHl6l/2RUK7m69SriOUgeMLon9NOVo45/hF3oSUCcs6B9S
pEnq26QDIuTLIgJS+DAPPEvbeNRFgxcruqdf/6d4R86W8elLW2wZoMVBA9Am
yGKunM0GyjazQwcHSXfLk7G0DHavR61EYkYwIOFHNWU8HGu3VDE1l9bQ1aBY
RNt8TIeL2dNTYMCvAdoiTeMYMIcLRHTi4UqqJV4vMDjA3/dGH52GW/Cmt5TT
4dtQPbEqDTYl2Kxi7KkywejJlULz4pLzoLPh2K25bf9q3PfCF7j2JjzXu83F
siNikhd8u1ONWfyzPMoX8mmc+PIu+Q/pqCQ+SS343bp+CoXPtHacTjQM1tIJ
zFFny2zNYGRKiJF914CdRQvqUmjEeuitI65HFIs2W0vs0c6U6lZJPwOek7ep
XzlP2n1oZJQdxAMj5dgEuArIKC4KnEl4+LI/AZ3uQedqTwh4lUaKK3+U6LF2
ldZqFcQ9S4XEaqx7e02A+j5+HSi7zfAg8IrWgJ01wfboBSw6iQABLr1pAb/8
UOd9ZiTc+fcXMC/7PSbN6WBQBpQixlzD0rUY/dq9mqCUTbypBeF8mMhD9G2K
vjCsBoK29SIMucDeo9JH3vVb8fX/96YWyqOhb667E/rRJKKx5S69qMufrIas
MZRgVyxMl/mF//aifRAGvbQ/1PFAiaiNffooB8FaV/1OplQK16sUwgq3fVkk
6gL9sVIqKSIbF+vVl+Q5H9eYoo3GCr2EQg4ZIF6ZVIP2M28k43n2lkaDDL/j
/suYDytNsoUzeL+TkoRJz6bSU3QqWo99nG3LE+IE4TZlNPrNGbi++lY+SPAm
I5Hcbv+GHgA+SMRy8Ag5y4M4fsnbbwvM6huScrJHEXqy+tyK7JesaKAAuM7p
WDYIBuLEkJa5uc1w3Q/DmwO7F282eptnGYK0sToJMV14bLuR4iCqdhnz+0LB
BMRfRSVv+HlA6Gmp0RORfZ3x+Fg1KZ2sxFCMmjNCbp+SlCQJxMDgfarfpKlC
TMd+W4Di4JnXdPYXQ5qn0LoDX2SSfiOThwFUHtZGad5JwfB2k6Rp/rXhSc7B
uzJ/M1+FHwlpKG+pnIqEMvK03gmS8cfCCnQL2s66Px55Z4MpOcUPQdLKgsYf
eYXFajMAAvuT2ADoZVTaULKw7AkP7JnnZeJgxnwrpSdKNqLvsdLGT2shkeIe
obV2N66IKuOr9iXrsG3rjbUVm9V4yVpPNh3a/nlgbkmwM1EPxVYlJN3cYHGT
QUh/OSovdlJnUOJ6ZXQu+L+umTp/tTVBz9yFVGsXkU3tzTSw+rPB2KDofMTS
+FiBNdvF5w4dESCoFjaf/rlMS5epntX6+hdMHmmfaoPxwUSbVdO9NNrflSUS
IjT5P92yg2uxsvp3oxIP/K4ZPJwlV96ae8FS149SubxCa6L/SeiR4cqW+Gzk
543ek7g3x2cusyKeliMy+7nZ2mHsDWWHW+pM8Dtbo6ibvSIXEASDS1FoamBo
qSIxTNKwjngv9hFNfZkksGCdSRU0pFuk1H9uH4sqARNcwIRZLFaNiNI6DfNq
Fxq9YBbZ5shkoT9sdP16GO05bK0XQKMbuhtGJh+6vrM9T6LquVAUc5wJ9HNW
FUyXRFhewhB0Ju0AeuxJee4daM0k9Mp4jPppszOXTrzz6EA8dJaAq/3WsfKw
Sn6M9cWpQWLgy4xgEuiIsa6tGXCRcdsba9LS35qSDUdaHWbnFC+7C1ZwuRkO
RrLqBSHC8myHLO9rA2h/6h3pIvdf2DdJ4FvV+RMf1KcQ78Zvh4kJjESoJLmj
4s96hdblZ9MKddyLHCTHdRqZGvuyfClQfsaPFjS8vUqvFeU2d0AND1/LCo4q
5R7jP6HvqjtOdc0nlmGCgeyMa/TGKm2Vj5c9s6ltYWTqO/ThLD0xXb7J3Qu1
7KgkLhuRNVxh+CDkSZPFM1UH5BgDOcBncya4zbK6wEiWhoMiSRWYNX2UMuD7
vLwh5pLJn3MlamV30jP3YDGxhdr6v0Pdu4ESCN7nfoeEDI8nA6ChKgGobarg
Hrw2GByfVmKJIfHo9WUaEEctpOp/lEHn3yfhPjFghxn9AYkMPuCCa4lpX+29
KgchGP+gqiuxXMrFV1bP/o+C+NF/saK2Kdz9x6sNciORQ0ZIH4QUOMKkrCHy
s1rib0mCYiw9cQG2Niikm2C4gFjk5yt+PQu2+7C6swLA8bVQz1JR6YgRqzd/
vvKEh3ZrQU3R4Cs7QbbYQ4wEvYSwSw9xaDh9bIK0yPQ2+M+J4o7fldRAb+IV
J18MtreZVViw2cdN4amwtQRAkZliXmHuyKVk+CKNvyVBYouufljK3UOONBNO
GC4XV9b/ttVS3cKqpK6xDhg8b8ks60t1olE/Tc9NmCvJTKUoolTjg/xb0uvk
v4SHfqyZc/L2BjgRLx6iJZ8VNk0+INJ3xDBXwVYnvgmavzPhWoOUIHb1iTIP
FVfltlFr5CKL20i0CUcMEpGGDuXvPPkEfMSVBSPH8XW6Z221hkte/+Q6DEii
sMGTmjkGY5rFFna+rMW3AU1+S1e16FE5+G0PU1cJBBTWLOz7yZJtpK4KTWSI
lT4TOKzhjcVv0OcY6AuLjbdWYwJmp03k986QDGUDXjatfgTi+6EtQi0oGTna
X6E0Aogzui9szEoBlpFJ2waphRuRDgf855jl6q4CzNuQ7q8YYDap0HxWkDum
/4GP1kGiMJdBPb8oyLzBghEY1p8hMBP5ZTxJnLKvFz6adxFFQz/8EJ/EhSTq
szTJgCVDwgePwHUmi/wPIPQz8rKQSHX/DXUl7jUfjX4HDa1CT8+VNuQ3GwIw
N20AbuB08gmUTSLpj0I6ZUeBBfSppIEnvD4RpbhiO+PpyIPN5TLGriK8JNw7
xYPPkk0FCHzQy/Y3t7nKALwP7ZI+El+J3WPv9k+9nLLnYiJ+v6IYxmHMuedO
ur6rsMZCdgSSYtwRBojrVkgRh/d4y8JQG/qHRgqX9VdjLkoZhb6PK/7m8BTq
VdV0lCGNnvABWiP5isGw41OUsTxNd+CStrY+3M9Ly1TgdQQqp3S9M8eUKTeh
bZFYkIg2YpVBo6bABopsN/wkE+ZxOht6kyTBBzgRuGQfczwUnw/0u4zWvzqG
V8Y5+EQkHvHrVhXVsFNaKU7F0EYrR/6e2MN76nlYqzZbGNsIiQr2LDrNQAwh
fekJ+YVAkIZoXgNm+1Pzh59Y4yWofqqDkK1GRTrjrrOWnpJmTRdXe5Js+x+E
fhEds6P4ZF70+ZkHrJ6gRVbmvde7SXmapmTixeSOe/5d8TfFWUirDXzZWCgF
AZ3dyjXg2fcYCuvz/rHo7m4aREaEYKARmtCqXxgPKn8llnk/876cH6zTXuAY
+ypVXkP+6xQDIiScuRHAA6n7WNAN/Rj/dWNjXMBawij2IZTyqLgBWjjTRv99
BCxTjUcnXvXcb9WZ9iYQ4y7kpVePzvDl5TcpOH9owhrbhMqq0YTAN7GkSmeZ
l7U3/cYmh1alHGIVdn0Pkroprz3kZZuYcQf1VxqDutFxeXNfrdl9gwvW2Hpx
3cXk44asV5jXNxJx+Z2p8JdUpHLVSx/xLYo4nGtKCtmf3gQlPapPHDXIUAXr
KrR3vv3IYkR8+tvxnvFQTA58AsNVqGzLxDhGqo0e08wBtHkccDPIKlwiqMaH
90xbyD6Q7fu6XtkjpPghdAb2C2K8n9WfVBpvtMpawCKZ5sSCJQf89jFCH9tG
YEzWjYnMF2R4keYQFoPOSFsbp1tCB5YnfMqjek0BsOs5PNWPjO28At5zydZ6
p4mK4e2tj3R1DdnCRy1FitCV79Bv5HR5RRu5avOQ4F2Q9mlwls8drB+gRy/8
gkCRVqesS2e0hJrKR6Jc6XY+GVMfpz5rSDczRRdWosNwN1vjYdtPwGgAvfe1
fS1IsXVI3WihGpBrSN3BlI+/vhPMe0Kcr6UnBpkefTIDloFhGDCAty7xvXWd
tNKSGpWaz0UhEkektP55ZcI8itVQ6BwlRRsTRzoZeXBeqHcdXuLQBBQeT0Kc
hxksbdu0WeojLmVjUX192mPvkS5OvF2NU7Vp1RD9FFL996+tPNu9p5V7hl1V
de8Lgw9dIMNZeZI0wuPxdZ6SPwXfFWiZfhn5JopYAwzptgxedB2BeTZc6uYS
e/uk4k8UKND1B8PmQEQTnhiGIFjDcOFQscxJ8gLLsrHN8h+LS4EYVXnTKuwW
T08uSOiNHPTZd780N6kVNY6He4dPM34vHZ60HBXQah7lQR6lPqDR8jagTfzV
tqQkPppOt5s6DSKJN2K7piAadMIklFKdBl1ZHRMujdNpBIvTijQYoeq7fi3I
vhT5fk9ATUx22oa7kxRggMoOg9u0+8IEzuQmCN8a5zBkX3kXRVCWTQoOKbV+
EVnyHvTwdw+fgvep0bcLlyxktJe1Jc74Wp5Sgi7S+JWwgjMORKpie0EW3LCF
Ibwjux2YcTFZP1nXFVk7R73TSMiB779zKzKdaBNdSvXieTn6Cm2/3i0xQ4WU
M4Q4xSx/oagioC+YWQoTIQJJ8Uc+X3d0PICUaLQGfPzbY9jsRd2Fddj0RZ10
5/GPyey9imdzILE7tKAxgb43Ob0suvbapau+kn/m1pD4qz2uf3gDi9AWdfTH
vdsKg1tLoGe9bN/iXS2sUFJ26YZi9UoXJ8b9kdbt0L9t1Kt6SE4rhtlJLSrv
S/nJtHY4/231lEhbFe8fxjDRqb4iSi32pukujc5zREohEZuUwsmeJvn4+E/j
hgx/MoZJ/SA0rCGqVP3UQa+LFsIm2+I+v079I9tF+vz0VZ+Qtruqg0sIev35
DEHSAHLUYPY9E6UWcTW1zV2RAL+SQB9XvNIftIZIslKWiZBFrqmUPPFVb/BR
what4hH7M4o7xQjTKy1GhFEJYXm1KT8bbpxyO/kYHVdldL6KMbCOhmLdPTkp
tFm7WRaSfyHAgbewoptMjOG7K2360KPHo+poYW3+EdBZ7WmyI8ZRkZi3jhuW
qNFdgejCiI+xjF5eMKiv2YAvSXUdSJJ9HPf+50bUu/nu1sPMYhqwBv34hmbB
d9brQoDNeZ8vk3ChlAEkI6uI1qr0QMIL8vXedHlIFxPo7AQL18b1uB0tnoKe
JwWvHjkdGUEJUnTa7KNMhKhJV3rtoubXoeaZdfpQFdkrkva/BcB8MkyrbnU4
wNdVVn4bYKjmA/amp2PEMugIUdaSQb0z9orPku+pYbcLH0DtHiT7DE6aQOf0
ifvKAtkxuo0t66Bc7tMdSs/ABfjEsvPxSD50Os7uEo++6F5N7S8tio8jEVFo
rjIIiwvZhEVI623kgI7HFy1+xIE5AjKy4riMfdixqJfrohmt30GSfInZIEqc
qwmYRSZIY8GSDlh8iy/jWpW8yiIXjOuFjL76+JVHV4XHT6qwAsT4AZHW/fHA
sbNNIyt8vkVExhtV59yxa+WF7hDsTt//Twn6Mt8mdbyviy48aGi3tBb0xtKs
b5V7RgLmwpnww/cIZ4dK3mOieGlRLXorgSPTiEnhdTM25keFftKJ0cSBnPA6
Dtj9UxRw9dMXcaJwYLb2GJ5RJPbRFcCE5wZOrhZFTU5Ez5fn2mBi3PsexndV
FsLSzOiI/K2KP7mZvyxA4MO2PBZHffb4YRdTtiide9EARBOVeTG/Rsj/ESx+
qwU4LRWrMLirIRAdkWuj9Ud2wr1x0lhfpAzu573LD0YunywOYq9mNK+La1CP
ysVSq2b5GwKTBYTiwgWju3r3A6yH0GDwE7GpE5jVmW9A7u+1lp7T7BmzT6ZG
IyQw3Ty2eIlfKm0tzvQ28Mu5doTe+ipImUFAOruqrlR2k8Mly346zpc1nqop
fvTolz6joSMaOn0KrDFjLU7g8H6gB3WOoC1z1r2XshSdZ/uvYRR76QKEagJx
YOoDq3K63zLdTXbmRKohKfQIbme4nMqWvzCxdj0WV5pSJru8ahKsxX9TuxYY
MbZBpdz7Ob3eW6d5PtbMHglM2CMl+3KpyV1g3XbPfxmxLTLvP7yDGI0vOLhW
1AQQncNxorj0WgjILdky73fGxW+2cvCMIVGBCSTKqiZFWsVXKmMuEwBSmI6/
+ohuIfEPSmRd8YvuUAEnwBGBmsOHqoKpFpgOLlrrPNjAKvqxAKkq/kOVZZQ+
mJofBVnVdmMVgnHER5Hx2gXpNsgM7ZgLTVNAz+GUUQNYCRXMt23hHQ8ptCvi
+rP/UHQqpn8D/ZE670tVru0UCk0LO5gj4hn8WAxu8aCOO+GrTnqRndkty2IP
jiETNN+pv1WH7S89NPiKsnd5fcyO3zoB/OS7MSIoNQ7mYL+EZKGCWuGM+4QT
TzQ2WkXLL+RQ6RaYQ7k7s5R1H60jJMg4C7yGwMwsI74uf22CQQLU095SW92J
QJfa4UxNmc9OH6iw2Djk6Cy7weXfLhGr0cBtFW63XaTXMZIK2TnynyZ7T8ER
TISAg6FA0766Hl1pV41b7Qb/0LUc1ONF/Y7zXGj2GhF2eEOw3zgMZVVyguZB
BFsxhmQbFtqEY4OIZU+GbNBA+xGRiJUimBtIDwz2vbh81yE0YV5I9KB/46uR
w1XHKc20kl+53p/VPaLkWstJ3jBiNtgulN/Avj1N4rvNGxCfgc1jy8GyqgAq
I3OIqPwV0NnC5/RiVHx5HaBPeDdq2jKHivlcehJVbjJABVRXdAHGgueRxL1a
+jyDvxEGLgCWPBV3i1VCfShE7sjZ0uJfPNK1hNV4qlCkZxZrcb/PpGo4AiPE
VfR3fcg+4Ig7vX5JLGtdpVtE9/PQu1V/0rDEhGfZ2rZCzCcqfM8qa1v3n171
oyrF4yXc2bSBzLFghqtfbBqY7h/3I2CrY+g4upka1obGAsiV6vHT/UwkP3pL
wt4jLzxTVRLsTMOKGbWsi6YGNGQ9Ang9iB/Ep3KI3RmEzjr6NbWp4h/IKcLt
7sJQ9Ct8iTZbolIWUp9kOkUuheuNjkpXWJBBvUCWHoH3RyB91jOVoKFuUqjW
cKnYUOnXMpaVAS9KM/m5kbWPA1u91yKLzTESgVef8jRTsw4eSL6Hc/5gJVjK
TidWDlLh+bl4WXNRqQJpYsPGyHomt0zuuuZ4sCO+dq6JWwalnOMSkEGGpI2L
ya4pVK/wdllksPoGoaVLgFAPVz91/kGUyQYkujUOG2oEcNeOFrYVALlfI90y
TwZgiHvul0R19E611JkUOoEivBFNjPKwXLagRoMgWnrYjLcoB+35Dgvhm8J1
WTIweWdmrJlki0MemavtYZHxYrLWBFEDY6/uJTCYU9JLfoa561CpqlW6jVZM
600oxYkSUWK9b2ndSKfw2u9YfOhy5OyNaf5zVVsJ5mJOSCtmSgeGJJF/1VoS
72IeB3CS1fTHxfJSc8lChGCW27MJ05dQNMLZfZcepN/ryiJW6oq29Ybm8i1u
ycJbT5nDBLdsIC2DyMhruT7NENKa8vjH0hxdBIjlz0q8ZaKxp65cSj7To9bR
9osS2DIG9uYf/S9kcS/NA/nt+74495YG536stVJtnE5dnAxBZrEsu5FKlICz
1l1XeIJ3yCF5znek4l9gn2Kq8kD9GOvZWTtSc6Sup7ysjUD0UDV2LwfEl4jv
16mp5UrFVWPQC06n/upcYv2mFxgCP5cKh0mXrpX5JoBGhPH78enRsJtHDNXa
vBEfhq4LQSIYUpWQGRPANCN2ShfxwbFQK9b/BEfTalxLmzZdlRmw0n1eKJTH
FnXbKEAXBB3ObysnboEw20IGAN/jbRgXhIp2OVWFvtLxXm7qEFtUy1y38q8w
CojZTnDzPTIGYjHFx8ehQ6BdE55LJoRzI4WqnF4FzSe0efqy2+ajTnoFcGMe
jK0yj/CPovcKx+Pwjgv9Q3QxPYJ2XA3U6fGF4/blS5hNIaY9To/Ej7OzmGTj
HXPJbvKwrH0yR7b35gXCMftC58eA3DCnBW5Dyl6OAogL/s4zzlFkxfxUpP78
0i6GUlBErY90a6L4aycFy8+FyOVw1Th0YIFIMHh0F4Y8CiyfiDwEPUbboYdd
IpC+sj19VmIjnPXCzn24GrjlJw2UvPGwcBLHuripBlrF22WYOlGN/EU2ecOT
FG9+qgX59rZicf7g6DFm1hGhEBb14y9z6NSZkffro+p/jZ/TbTmraL63Cnsi
ol2IiNhD7qqyTJgB+5mX3lMUG4IqOcL+DIJGqWhBIRyE1iZpnEPg+JbHvTx8
sbQrbWjHrOyXhokpeKRIaIjWiG1DhKbnkiMd8Kxf9rJnM32TuortcrqxphCu
5yUxCnmG0E5jdIWi0a4ekrrnEdykuVj7eEoNQxaachjNHx6O2iTNnXDe5Uhe
dA4m45iqQGhf/lQv7+8wCyVtgIYvEiaw4zkR/GDBNs2P6wlgL5BtjhRq7jc+
CMc3YMp+QPdmmndULZMrAWaW0P3viXL7mV16X8IGVmtOdmkgFvHH6KaD9zpF
C5U8vY6/XFCplbxxpGaHLuJcp1BjO6hjePllEGOyYJ6Wggu+wyuE1NBDK5DI
a5o9NnMHyxl6ORjQbXxJql2WQSeyx+s1shbkaooNWMtbxcVLH0xEoI8xQf4e
metHOduCaenqGnOB8szqq0EQIJRbHQfipcxG1Nm+nMqitIt2M+x8smSYd/Yf
0sNR5BvdAtADf3LJlg+fcxKbadxzMbzdw4asMHV0NXjyof38j5JUnSCCFbwq
tC1rnmYnWOeNWkZZ5weczn5yJrfCHxdpnS2+CosKHmqacMLr0YWsfSyzj7gG
8cDDmgwTxf1Qqt5KJ9NjwspErkbitB6ojFI8n9+YJVazNHA35+xlMDG8/GHA
1B19UOe9uJfiqJCfjWCBME4HAsf+gykwqnJ8cIFKPQbJoXdF6+ucx25EJaDp
qWLlfjqHB4H2ZnQpG8kmb5QD8Bj2mzLvbHMAzX2kQkkL8RBToMIHLtUqHKBy
hfZSgm8Qkn4oeTc6Wd8MfXNh1yPmCUcrV7J9C+tJAuCgam6aQd7jf9MrjiZU
2EuoiSVnIOUEUA16k6uY2a3vimKkemIaf7IVgWhZJP4y5SzqkPLaLtnVmN9N
jaqQ8tNE5HWpN8ZEc0nmnAQZhq7lgr3Q0hGLkSuNPofYeM9/t8QYODZ6AUDo
xehOxnMRRRQ5TwYdmUuwrp7ZmU2Ht2N8pwe7zVyW7XeqhFHKRfd9ytcjN4mx
GhgoNyzPL5pKrYmiOR6A4FFaZ+byQySaMtmfAW4G3nokHhgoZXm7JAEZ+tX/
/wo+H0b4W3cObQC7+jc6ZvmaQmXPZMBFZ00Wqr0mDUrJogXmnNgrpT89SD2u
vhNMxJWkrWP+EsBl7LxJoMIC54AAGNICnzkTw+bBbFReHtHnLJdzrOTxIl1d
ZBgHGX19iJ1ZP/j6SQDxHs5JGPqg6rzjszW6dSrkEJT9xh79ecyx0Y4D6ueE
L5L46k5DKqdtV7/TQu8SLPUu2z85pYt05FibqK22i0EpRsPp2dsg/W7BWHfO
oMy+IoBqyaGmh9NdIxh69wBZ8lWIxYONhHfj/k9soq9Ch6lUzDNfo2eaSvpU
IsmjMDj3I9pGIOYhJ37tXyFlEEaJmKB06yyVvvpO59Q4hgd+FALAmeGtgun0
pXOOJBLaFsPlWIc0iu/qvQsY5hG4Oh6m6pPnIwCRlGF40d4CxG7d7H8S38bd
4ZpYtmw9dfejClkaiQfK2cZ4OqxTxXN881DtekmJktgJd45rP1uvv41XA6mq
rLMxG1RuDtQxoVYJ2cI6j7tB/ibKPnwN5kIG+7gWo5cuE6cSDeXBCBA/v/DW
p1uYgrQ/nTpF0k1TSnnRT67X+wbLCDmVclf4TGWLLyYOuHjLCukQ98ijkp5p
dZHgJRypBwUrUPblDPI0FGYyPoxckAZMU4TbILyS9+X3t/ry6mQkOl8AGIyF
TOa5vW6NGZ8A81nyWko3CH8ylEAlQ2XNBOHmPfUawhgU62GW2HFgOvkeLrO5
pFpx5GrTJ1+u3pe2b/6xf98PH5byV5T4dG/1DoMTwGek9qmGdEuzojAtbcPx
qEaeI2x8lIZhx1MSJPcsmdd/UsXMlMgq2WS4jp7uUXtLLZcIzBqagNgcazOU
W2AvhvbzCWLxGyBlVFtnPCrOd2zc7LYjju545Mw7gBY8G4/gCHWd1Ob3UpWz
Ie1JVusbZqp5UeEuHB4bPV5c7H3v5FNOHQGFzuMSviP1sbd/2x38LjFbO3Ji
zuJGdIO7Clr08nSjkLQ0LFwEfI1tX7X6nqEHxi7DjIxLy3iSjrG3Ccywd51j
hjSYeyHZMzbKnnO4OVmkQTZkxpTjQfOM+t2x//8eWsBzFuXi/AgFvMZWYXJn
BNTkYCnZkAJAbrmZ4yFVFVurYg8cxX3ujVO+4o3przN9JcET/HP1jZ++rYdd
EiuS9PWUcR25gRIewjLFZr3QmEpHNpM2+zoUzeKuJ0iql6kduOD58kk+H9PN
aertx2Qryb+w+izSpc886bWWaGqcftQT7fC88manuv1JHKhrk9fXENRs8vT1
H2n5wiwvXBWmC5qxSrikpUKXELVSy3lexPgF5KHi2BagjfuNnI6FjRS8jAIH
0n97+jisnykyM0gERQEaHaF9wDqvBQqC3Fi0Qjxtu2+2nf8Aj6B7bd+PgbvN
+Yq+xRSSXn0xpmso/+yZau+qB97mLFPuHt/8as81xo2yobNIW+HciVqChqL2
OEBA6IyAMdvj1kldVttc68q7n9A+E/dQuP8XHg8prPoOrYxXL5q/+zBREGLH
jZv9e3du+Z2E6etCOjpyk1Sd0IAmC9QKjcWNkRpjoustEzMcDu0eoEV0K+ZQ
141jn+ZSPQa1AbhLBZs5DwGx6FDBbmu0jnjVRLCdgthDZktkXLvi6otBgTqN
L2F2hMhbT+gtL0ddZkciV086zlEVI1BLy8LwAGa8rQDWXiOy1D585otUYBRV
pK0+ApobmAN53/JBBtcm9qUeHmBhFJU/ObtkwRnVSC2ZQIeoHo1v8mYIWARR
XCrqG4MDpswik0mAS2PcMN9dTrooeoKc0zjd5Ei+LenJLzuxCw4iPfkKC2bV
rgCi4v3NKTY2iFUQ6zTLm1zYR6ifa+uAKtHXYyjY4eQomPSdcIf/LEeCDoKb
j2+KO262uL74/mxhhrheX3WTRyHZEOJdcaJ5QE1QPtUz5u2qinnZtEP4rx3S
/GnOx4oE9FtQRX6at999LQOmcZwQ5/+DN73p9CBcJyzpeGK9M2O7Z8DmH+Zv
O7xQTpR/6ss9zVoAahSMbvx8RcxTEfA+zCdR/490eSq1BXq1uYZ4IuC22HSV
RjrseYhmYNjyUWDSsESfQieJOfbMNSB6Zg/dpZWPnk+1anp8CH57eW11rpWI
gEf1stb7NGcd4Ulmn1JHkw4l+pd7zm8qgvoaPm/BWIf0PFo7ms3eQNGCC1AP
ZKHrmiD50s6IjwW3KGxB1fsfxpJhpG8foQCGVnzsRGTcs+tYnNaV9USL+VoF
fskdQaj3X3kSnBvKkCSRf7I++UF76xwO8I/jNHi7769bCXy0cASL3a/9Du+u
hJNce2EWHp2ObPUMGwyGhtmHgaEJoKP7uLn02wjcs53vF9ECSMTfIZBbOed1
u0MAJAs5A1hpAx4t2OVlJ+sPpYTohc6pKPrUp9PTtZHt7GkIjAciyJV0yy8m
dy6Pp2x0ZeX4cUcqNADVXoTyj02cgdUsoOKSSFGTBkMIRTWdVAzhbWYt1OKe
ixkXwZ4pvqq+rN0Fgbdk5nz1bzM+QeDxR4WNd6De5gvtUYMi6apXAGgMyDod
DPDkdH0tjS0+Jl8wZ5mYoNuq1ix6KaACbGQr16/l/FCQ7+soAU7VrAvDZPhE
RwIglq4rwQPCfoRBe2aTyO2nF7xC/zKfMVIiTcaShzY2dPmKfXFHIr6GRWQN
Vx0oOhYSPRrYh75Pz4rdj0j+9aCsdExkDHB+0Sl4tns5cA1d/mLZRxXsIZ+R
FzjLjNndWCbbV1lmqck2gEguAxrerrd0Y2EO6Rb/NV1zcW0KU9CVPFgEw0bl
POcb/Cn0vTb9/U3jovZkTx//kQRx8YZ9u4lwzQiTEkD+SblYF+Z3J3zQ0yN4
kLVEEBHV9h4RmlPeQ1kiaNejQ4rqtgsNEtTI8OCTXLyF3drEIPfJ7Sdsxj3y
AMq7/pGZgOSSvFbICxsiJgbSN5SdtahrV43ShZy2JpB9GWZowD/dnUOjVOSG
hOSypTwjYM50lDIBG8qTp0RnXS6zcoeZkUBpUlnLDBZ4un4n3sMZcY0MoZMx
Mh2nTalgMKlcFdPQ31CLg8KmBR/6qK8MLMWiu9AsLvoAFENvt7dNTpUwTItb
GGQCebKVLu9A5fLRETqxJZBCo44kDs1KiY3bNNTgLVBUGy942MW6aqV08Xl8
scWA35r37C8qZln/OwL/fDwICMHqOCpf0a0AMFkBjpDAbUfO01Ye+l9G9pVk
4EcmNu/V0LPcNEQAQCta8TYrLYmyIfNQdBLnxvgEdEfla5LzoTTnepOFCO36
r9XEz/uRysIaEFxpxHmWs8sEvGwZsLZjS2j5cmA69UVdJoxPTPT32PTRdqiu
LLSp/ulEXNzElLMxIsaigGPG/GtnX+VbuVTiJx3/y+MQ5rZLO0CNBx0IprvS
3hWf+vM8dB1HF3g7mzb146DrmDTielJYE9I4/YJMUiASEplmePhgiFEHuVU6
FO2vHKT5VdNkv8XYrNZdVN6lzxgbGfmyg4M6LR3bD1Ibz+DZblYnONkQmy6l
P5qqlEjbVmRaxnmJ/g+e3WsI6CtJQiI3O0115WR2lltNTXXSPwxp39yvwv2t
hI0kwr7LAYvezmMHtDIaNP/Ui2j1aTDb0YCyROBnZtoEXqeD5xIRpgiGjiYI
cJ+ZXnaReI+tzLaczystdenv72kM15ag+CeJWWDImXNC3w4yvUE4N4bWPiU7
geCKi/E94QPRgC0shH6+IE4nbTTcysE6NC7EMaLGWKsqsRr0DYdJ0EIUmXf9
6cdVouqQNIKksEYeiXWM9wFEQzgrSe2iexpk3NcZX9lxCp2i9giEAWk9DMjt
wPyqGJLakKM/2MXZuq6tpoIXK7rFCJy1piCjfEXYMdSvj5pmvAOCU8Xj9ZMT
zgx4ifvwK8Vg8Gcpaluq1M9aH5whFPe1CSgM39cqaz2WUnLj5QDQz3z2aM1e
9Jc137WUmiWVAy0C8OVjlHa9O3N5o4qq1QRSyUs88si7V3n5wma+munQBOQL
3qTH6L84v9bvXhQUxPmk1jjXy5UTbig/montNDmXxyVNHf/yc7HQ3DH5WQX8
MevuE0JHO/dZUEtm4cFJyeEuyPdG+cG9m3l0jkt7uO5guMD7hxe9PgXKKGoJ
EiwCpfCIvo/0y0trXSmb8LCHYtlyZ42D46kzDCXOiRY5JuNKynrq7O49CwzQ
115cymUOsRedayBn8cg/4BLZeKQ5u663di4qIRyw5rFL1j51+6DgnzNcrrnH
Fzwf9zBKGxWgq89WGnYm11zLrw5t5+BmZFcBrmgPdXC6khIi5fmUfYHGChaf
bfqqVdBOuDzwcjhdNslCSmCiHy0n+6G37bQr02JBBQul1VSCnJ311Lz/g4ns
BH++wrzPn6dypS91WZs8J6WaDrvGclRYX+0ntYkT1lbOKhxJQsGNjncSjRQB
5aOzZDbPW7f/sTtnUt/bpxMAU864ehalxP1/cPl0bxr/eaEko5jUHJLN3k0+
UXSNAiWd0gSnBjjEdXXldsfBWPQ+ma7MxSuG9vhIpAeN+NqTO71JaL4TKKmQ
knF13GSBwpYCyGAXsIVEdHsHLtBIR9owtrGDZXs4ZKsVCYdJcBTiusTSMd82
0pd2M8aAxqJtyp4u2jbhRpOazHrS6o0pny0trZ1WUaSnFPf4QX5C2mjbnwe0
Ammiq1hbASTxZZANI0OhE+qrDSwVVByAilld5uKDLV+VTyFiEvcK34C5adWX
zo+ux01siRkcQianEwLRsJlzsHgMmk42e2Rj7VHhjn3KOA33DJ4G+4ZONfuv
zT3CV4PXkvbehU6FEFS/MBbjBa/OvV/vpCfUk488tppCerPCqNrc46vOakbQ
2c+ufG4XoxQ9wMV2h1SVXOjtK2kveo/zQ9ELCXjLjQEuPNMV6/v1//0+bCr7
Cm2uy+ZDR5KkGmS5R+RkCwzXe5DF9M6rXX7FYG6O0s0fwovo5/KvB0/I38HV
eB1MC5T9X4LzGymBkl49VJCyYfBeYoTR53KTOR7Z8DfW/KJdzAlF8QLEpaGn
I2czK90DqbdVNJNX7tw1CikAQmp4OqqXIn08fX6BQgT8VR1KemwGV/9PLz8O
OtXvOuZ9+REdFpA/TFovcc4h6i4BQHf3BZZYT/HwmH/r5sa/YRpmi9XiiLJ5
udDKDPrtEksY5xfIz1Q7NryEhJDAt1X3OL4QB9ldlz2+81y9kofXnbpfBrny
oARCjpoyq6fkwpcAEqtI+W6YLMhJwks3TcUQrNzRlsz3Cco+CMAZJfsgQbDS
xTyDQSlJnFDzytEH0XIniPqrWnWKNzYrJCzGi5CYG+czUvWA0LkR5UakWysk
q2OKefy3z4utEIAswvkQt5r9GZFlsTweRhrS8IiXnX/X4U4QPDZJbGukEYqJ
yjYe7BMo/KHdt9mV5Czo8ZJZDw0oSpl9DnCMkVgHujU+OLzPioEB0lEngf7y
l2IGObxeri63eIRgiZRlXfm1Zktm/Fh/5YVoTFFISoKsoKWr1sgm68Zujt6W
NplnE+N6lzTx/eund0m/dEjG68IY3g2F3Xrtzw23ZV0WXS+8j9Nm8DoCftux
PFM1T2e1cDnr1kjNKmrGMWZbiFDfpvKVigwJmC6ptE+sJ11tTmP3Egb6f7fr
4bc06oNms2o//vVjAWY4o4ZZ0EyZNe1drxRe6077yuXM1jjy/2fOzhUCqtRU
cDPNJJviqmBQqzHiUufjXV+78sZiFDi2DCjQW+p2qUlEtosf9JwA3Y9ELRQt
t2iugyq/W5Ezen7HGBGXgeNYmx9IaT29tgW33Nuv8dc4liXtywz4KUxk71DR
fsKYBkjVbFalBGDFtR2k01YgFKMNSTTiS7AMjQL28WMQLLF4IT5mm1/vexm4
PaRi930qGubo2Hf7mpNybOgtDQ3dB4lKUjxw21a6z6dhl3ofp0gOXjRhOo+Z
JEDT7vNMO2ULU9x8wW2Rfjdeoljqbj1Y+rvrtqmGDZmUDEkQwSQCcytdQpRC
EinzD6P6S6mabYt9mdEdKUDBam03xR0OWY5bqiyt4ktHE7Kht0GVTIjXXedU
aI6YBHqL2dUZs/FjzoK5f7j0yO19u7uwkpPIhCI+xRBhWBloN2DMkIGwnfYM
98sjOLqJ3laLzEYnkJmryWEKTnlbLsJ1A0ljFPM8aM/SpZNIr45CEDUsn4gs
wT7vXjfSCGW1tZunAi6YhbbxELXoMdEC5PqeiMWMoknQfyZjH6vSw8b6hInQ
BAoZlThTCGs3nha38LO0W6M1Vsb43hmLgTsEg+j+ndIaL9W9H7B9XgC7ecr/
bD4fFrHKolc6izBqXvdxAMIbWItIf7etPca6/aGszqcRt1x84ILNbqbqfnPl
+gnNsByWpOtcdQ1OZ4BDObO1cO0egOdDtMYv4GtufRvsk+yWbD2O4QMKY8Is
Z8psHJnOa0tcOcwy/8lbTBe3whIdjSrw72X0GizhbOy5UsvtnsGtlJea5dH3
grSjoRrKTQ53ixdre6hpxhxmtizfjbe0KPbp9mW2/ag5ukSL5BfHTdaC7kEr
/Nh7nDXwVHPxECgUsdykJVrV68oxQuz5msGZTAHTELlRRChV7xVG78u92Lzd
pq4r2IryXqVQadrcRXOXIeYtqPpAsysZysp1UQ4ADWWK3BQT4UlNBzh8Ds9i
pJodrs0d6RRAM8RK/p8H7vbDvo2g03zKisqXjctCLGIbl5cHm7RSawz8EICk
h1B7uKEcWDvnkUb9ki5pnQLvQXHh3/JktlmPjLECgRXg4RN+ZM7/bb2dY1Yu
bgalkCwIo4+fmiflwgHUY5SqxNN/xLAxATgrSOxkL+S8jtmgS1X7tiSumLf9
aOoL28AVa28ixdYrIfKwVGyAqqojRnSw4WVtWFRDK9Ael3pUR55S+aUODzMT
FtcXyUVcGNouwrgnbPXaiD1X8Er5WCtVWXzFwLYsBwcXBjnK+3dIFCGtDLvg
JDh4m89h2OwOEXN2dGwbKZEmnvuec8bDZsUOBnzT7KnUkcbB+zi5badiA56d
4hf2aNTdNMH7I/9pIRf8931x0AVgDQBdYgWaI5bEaCqQMcHitmku2YcW3ox4
riJHQ+m8HifpYBJzBOiUXLiu7Oj3JuZK24oJhUBK7QedNHSN0fyw7LEiZWP2
xszeGqoMKjbpGoPpTJwT3/qBGtrsPal5yD7PWHx259mMSt3wZEBEwwE+nGXu
tKlQ6AspP3bPmqpUg+GyOYU8O/ttjGYOltjkDMaP2/1IkGj4OJpZW/e7mKN4
0W0IFRDmSbTAG6c6Sn3mLyGemadxzd2Z3aZsozpl4i8qnV3957ZJ5foT1C8F
vDHcISfK7fW6kZwre89jsMExnWTUBYbEcg0iInaODnLuqy2NoP8Ka1ZjW65C
Ofi9xSmp7rnduv+6Qzr/sP2YSVK49q1/4c0t2NwuyldG5QfdaLn7L2XfCdNa
NxaDFYFSziJkvnWz/nFIZ0thXK2qicHcBFfBquo1pd6d5oDhTnWWMKI4egdL
0UWBOefOzubSWztfJ6seeDrYZ9D2cASo3QMMhjQMcMW8M60XtnPUngZg/O2W
k389s9c84ljMT0IHHuTpcfUyC7JIagU3LSnTlPjdNLzg1Hcfyo5RDCJ0j0R7
o/mZg2dm7lqtRDqEYdRXqLyu3imaq032Szaz+QDMChoetuwiHZMHsLQBWVHo
u3ddSwZssWDKkUQVm7cCmLVWtB/RUV+/W0KA2Hg65FNinGpwuuEGA8wTxmPS
JfS/RQi9d6pGWQQYXVugGxZnHHJD/t6Twfd/ih4l/XnvE3WScAgDxHUhsBr3
L1Nv1QF5KhTJWbyvHwyIr3jOaXQYugo/eYFMYEV3bg7G/k8PW+zJ1RtIvTml
9S4oysNeD8i2D/k086lWNNMFpq5sZI6YSeoBGoQ6arU7z30YXcjILmWcTWaF
3PgTgDquNcz0nPAwqrdeMHjqAMrTJUaAn0bvydU8zOIxTErMl/qKnPZBboKK
EcsY0JnhtASugliGgEIbGoZlzqWCLnUThQU0J2NkC7f2jVSnG/GZaURnfwr1
5fPnwSOc/iEYqEs5AgIZEcWPzGqrlpcitQi0iRtNDqE55uvI90HnYJEQRFKR
KCQ0nZdDg72g15UZOQIOHnK2pad26g+pmiNwXDEBECxZDyLDyNqoFZr01If9
QxuFSAPmYuNQeAQp+r0UFb0l7+CT7zQHPr5U9Dm6w77pRh/Kf1Inn10G0B2u
zPycO2WJjruGNbAEuSNvK0r5zLYzh/SJXS2jW/QAp9xPKzQOJ4L4GxVqP5LI
NU9WvX4Tc6/HcR7ZIcrBdHk2oeKegyKsg2RhUAYdYMsw/N3vk4OVSZK9f8Ul
iMjqffq2pjO0YSVACeTyur3PVMRqMfP+z+aOoFLBFdZJ8J7TZ6y4cQW57V1y
Swxx/abDKSmKddPOH6p1UyFttGNE6zXAPb2nuNHKXlcvN9X+VDIjA8l8Cg2w
z4647IojO9iQy+yMNwl9vRRP23SwaAy8vKALEVxeAt6eogySdNLU98rR7dhy
izYXhso/WU4SD0jO1eFp85GssXicn5WhRBSEXWLogNg7Dcpcyj+tWMo6sf2/
QvO50e+YuH1H2qT7mgFqV3ronK1xSVQ//4aqTL3ZkfQxwrSlmNzzrMeZt8gf
Z7+sYKSU6X6hbVbEToXmDHhCOTXL/MAqtmw7wtwd/fVjsE5nR7qgVkVN8s1K
YWrdmop4iGOyEDKbfxKu3X0q8MK/5m89oiMe0aLePmYTvW5rWwe2mhYg48yd
tLbuhTekFrW440yl48OxZoD2jYgUpeNxBxEENcus6vptkOfZ78cNAHUpjN0M
W0HDinHr9RZB4XUYkVA8sMUQIK32YX4PkjOSLVva2tpOz39SXIo/7sxejE/P
P0DskJ8KKC+JNMlLZuF7sxA+UGhbLZ7DdjSUzpWXjE/0Cm4o4KB5vZMnoxO9
JUVjKBQtFZsn5WhEoHLg53o4A6uLSdHTo24W3UYUow5wcA4+TdlWuM+NDKMy
72rRCZGBtWKTPVNIagcURqMHu1kGImeSdrz31vinUPPP066b7DZu8Grb4dMW
c5ADpIROezcCIrFKvGI9+WT6NnYsllyqEdNnCqktdgPeGsXgFeDQKKma2E0x
Sfv2pBHOUhhOJqixuBcWvth5yijJHzwB32WFdsRO7ayDtDR2vTznAIR6QVAY
JSipEC3YFqiY/c9GzeKm/uag6tU31jNO2OxNA01pte2yqEZw2n0R3xLFBA7r
/wpHCG9U21Rhz6hkhQ6/+OCMhj1wYasHURhHKrimupnXf3FjFpdLLhXDksCb
EasfiprW3aFiK/UrZz7R0REvCddikK1d7jJpaAcs+COl8j8E/mMnNFR8Aqz8
xTShqg3YY+pBD7MppENJVSEs7OGeEWwDg5pwJwlb8ZE9PB9YuT622T4Fq9R8
MTF5jPinhQ+aHxtCCbC9GlAvDByZetiDH40uj6urWl1vUpALWinvpnDFkZYF
zZCDuEV6h3r1XDDWplSDi9mFt1xdGJ1qEl1dOov3KeQwtGBmjx3YKLci3zfa
qMbKsuv/c5Ldc09nOdTXgBUt5yFVTh0idj4BhuCP6lwFfNgPmuY22PNcHHY/
2pXvmadv5V8WB/twjScC0rfMgLJkGfI3UgJDC3+Kxi+KpeSgPY+Dtr+1yDY8
lunaFt6rFarMv6vAhfQMJ6Bo9ZRTKuvX4YU4SKi9t8YedKWTtQVUpvtUvDc0
D585SLAxz7p+Z3T+fs2i7WeJc50uG1TkCtO7ufnjPe8+m5//qunSPG3lAALq
H0eUXUUmi9+PPGGs1T7anklfyjnQVYN/NowcpiSxEWteCKjlY4ZQQFyJSTDg
31vK18BV92etQCVHBG8s5VKSKk+YwBThOsJ2jghyW41/3k95O5O2qZVXy1UF
t6GN5irkz1kgHDEx11cSNodWndIoWs15XCDdKlmi/4JzGjY4WbnzE/dn9/0y
v94aoaBcL05XKQ+bpA+aUf6t/YAIBJwzuLd3frbrJJFH87mFjfB5qLP7A1HS
CWbxJVFjyQnfjR9TiylWQb5+BlyM6NcMG191YH6cJ1Btkeo+fGm6NsQaqkHJ
7V81rsJx8neGpoPPjLz3yhLR0M5FYn3NGZ9z8bI+t0jJkFCrH5YEeZdLhews
0N8/PllomNAV3aHlk2FlpgwQvxt2gVmf+xwVd/KK7wlTDnSdMmv3NnOHEEyD
SftJcgsntwd1e7QRk+jP2XW43142iOR+RNWUQ8IRTcucfdPQnKNO7V7yOft4
XaRHfH7Zdm7eIgttCNsUjT2jO6/bC/XTXW9Rn61pVrLKEpibC0+0Cb1t7ZAv
Kvrg9c3KfapGjjmLOD/HOnrMk5VaroY2Y7PSxmUrYAoaqffIY0F87FWpqdYH
N92rBH3Eg6+K7TNEofhjXr6rsar7nvIKMC+jB8WbWknJZckO4jicJD1UXbDT
yDZdfTMaJDhTElEdBf0l6WoX8FlVsK7Oz/UW6a7JcIxO9+ZUYaV7LUc0Isyb
l+o1Tc0ELubiw7YohreciFe9pvqHiNDiLi3km5dIfT4x/zYULg+59UYFi237
6YhVB7Jb2p0+w0mcnNj/IpXbAZKgebvzm4DXeEi5gPZy21tySosjEvLkUNJS
vDpiEbuArhPmdbq0NAAZFxET0sOgiWoJhs2JvntEFnNbbwYPo4MWiIGQa/9h
hWcd4CwVaFDNeHbRD/2IW/yqa4kMPSEY8pZXCUxGrn2I1muZ164vgk2MKzHm
hhRyUfD7+SWoqX4wYDhi8u5uN8zGI6dXPtnLv0qVF76M2GMzjOLzSeh20krp
+q56RQ0S1N81GFLUPCxlwxx5vkcTwuY0J8kda9a//bD4HWhJdjig1cTTDxCz
IuZCv+A8RL24LBTpisbkmLo4GGchvww6mg2HbaoZxHocD52X493JY1+LptM3
pYAcTULYQlvcAPpyzfvrTVfMGxQolHeJaClsUnyZiJNGw82kyQfLykV7ncqP
MqsXPTKoLj1ps4oYh5Tp9ulmOs8vCN2GpBnNUgCKP5DkPLcd5Kx9+LCUNADf
dczhsy0lw9KMVHeY5uMf6hzNl49TKGHYP88Bn8lHwN9djgnmL4uuk3FFUp7v
fEmbfGVHOK+uUR+4bauUeuDHL4la6hk63K+3+fctvHIA+I1UQMhw7gqgDwsD
65s4VtLZ19kzkHtshLr+EVFPRiIyTUDPOoiufESG/0HhtqYNBe70P0UYC4TM
jLg8ndmDuWEf6yNp1WP9SsGFsdadv21DO0Z9PG8yD197hDn65YeKVMwcfMzL
jIhRJi/WBdtnay6mMXXdhNNGGGg2UxBcVGQvP/HhK+fPLVl3pth6E6QQrln4
0tPNlXnayZof1jggvWRLxHAS24gN0uaTWfwegXecfQjFZqew00zAYEtugXfR
5AwK8ywPSTqvhVu/awbAmcFoJ4Ag38ybhg2fh3ZQ27N3ywVrFhhoVWVyDXfJ
LNQWXMw4SNUjT0S+vXEJCuvbAg3yE8niBI9dJ2+/kihTugf/2dXXO/C3LbRw
fnvbGux0ygfcJnzuwsagM/da956qjF4pcSRQkFZ8kk+L7g7+S9pZoOsiq7Ze
Bp5eALaPkRy+5bW/2e0CKgOZQgDEzFamdqJ+WO3X7Xokdr8Y3KWc06cO4cJ7
587ujb+dH4kgSwrrPlG+JnqwFmf32AF6+1Lp0pZeCORKrWz/Ki9I78ocoF4u
IpIN+41fhfFy3gCQNYFTR/9ocLJ79Ea+p97tWR7yfSh7UmvDQV8IWzbj6zLm
jvbKKJA+8kXhkD9JcT61RDLwbeFYlHd4kFqFArIGb8WkeEltYEciJA6MVe+Y
pXipAT5+80F7rkfK3y7EcEEiY6OKfVlug2na/MS/9RNByEG6LeXhdMNNsC43
GzsjdfOLOjDxmPcdBLa9svS+1ZMf93Txy/4t28v6cjQ8S4Q+Ht13G2waqF1n
/M1yz7cJPrEh+kISB5jwV0LxPbOzSklZ9QLE7Bk960B70NLV5GHr+mStPsuJ
fPP+pxjS6G5QEis12lKZ/Q6bnnhBaSv2rxVwvkmXJo9DwOmDcRYxD06ca5/g
RzhvoO6hy/FgdpgDZbGSeCv1p7FSwpLVSx57VUxxSn8Z60qcctJm6dFC1XAx
kAd3ZSL8TK4jz+HXA8DDNu21hLVysNQgBDlGMz9hQvBjOYezcjHP4+dHJvw8
GIlZaVfUpXmtcSq/xMBxny9FWyGNnlS/lkjwle18JkE+Y2OrMY3LTzxcROjC
CJRAut+xr8mfYQFixfBMjwNsEYfMK2GZAMER3RO5LzMb+x/dCJbO07boQ+P0
maenh1XbUjR/BzEStfJ+o05OOM8/xtSUOr1a1EXMdo27EN53pVHZg5v4JpDM
nzg+jIMWy0GHQoLZIJ4fBgiE9BN6AOdfmohq/pxeUnx3NQFHRVeumoZnx+nB
RxueqZmeaPtOJDPveHVjN//FsI+hYskInxXX8scjnCcpEgBFokEP2thh9DqL
WnKCEDxKqVZlKPIN8eB7N0z3TAULiPIpEwX1os76UL0PTvtzpibuPoZxDXw/
lH5RhmuhQ96lWRYLJ/+Zjiv0Juj1IL6b2wLXNMYA+jaug640Z2hEkLAefEbI
S/p4fiMdrXuIMqjEK+cKv9FMt3ynQ7XQa6fYjP6GYwAEUzY7wdiq6wfqkyWS
qThz8DPG0KQDzB4BLgqxRRIkA0Y4dma3zBl9Q3WSqQ9kMa+TM2dx0Rp0ZE4O
sj3ggcJUqXgs3SFcrk1QrY7mPjAVG+j4aBvV8GlKWlTFrEbj80g8rfz8Fuey
zgwdZ/SzduFXKtyGrmrbsH411iJfz0u4z/OkuWBK0Ktc/y7ID9cZQE1rP8Jd
Kr3sXcha4gllHHkOH6fnx4vReoRosEpbQ3to9HGNlnaBPKV6v+bBvlKXKCiG
Cto5IFV2vE+fOlT2C0vnkIsDWDtpaxsw/LyDYYbd06Pv4xA05aXLFcn4oXDS
lA5tk0yNTLvf+OQ4vJ7e53Dxjwexsy6Bf68xfjlkE05vvLPbIVcu1J0VXpkC
G9o0lrg4aprucD+uw/PvebWxo7tHzYU/rm4TUxZ6ur+R35cQC9dLfWLYYPk+
bKNjL3VUMHL4pe5QOib6FR+X/h93GHgNqupfiWAQzOF4LGLL6Xvr+GBV5L5S
cUZn6v1VR3o2nD9Hoj35cSSScY7JyW8hOiTA6U627mh5+5bCyNDW5pn0Gpxf
aPeQGqjkMvWD2zcmWykhptCzpTzUSc33aFZYFsI6ZBKz+zWxp2PMKaiQZ7Wv
A0TtM5o9TdPFrVDeBse65wiJF3zWvRgyPlzM8Q6V6gPSno7gEtxU1TIGWfgM
aRRoeyV0uRMwQ5K8L6acG5TMl8POD4BwRnGzoB12t6irp4u6Mzeup0v75ajU
O3+zJzpIOLZFg7UcyW9JSvIfU1kXCqi/W31cFV7eQr+Zu2uSjp8gIu7IHqiy
MgDDiqPvIyH2uc1qxvQQwhzVDTlRS7fk4KMemSRV5y9egMqXzZvueuraf/US
Qn1/ZqkXRvsCKoBSD1ID/0XRa/9MwxPw34aQTSwKImbITqtpAmgMSUX3dWa+
CKo0qK8/CPpfhOD6Uv23jteqni1VMsXb44i6+XbezeGMgbJQCUe9LxcJQ4U1
qPwR1+g/4NLs/lZ0hz6qmhjxhwWhl33b6otNwGR9BEzchTy4UV4xrkv5r/zF
7U0o22qeoQ1wylLSA/QuLilikY7w1j/WkQ/AzLPt7vSVABuWvarlIIFyhnSK
G4LYE9nf+QSFBJNw9nQvJCm0DA0Li6FBxg3s3uEn1OqOQeODXFBAdaf6iBAg
lIQ0rXiq2tzyqw17Nw9JaNr+L3smQVYncyAhyPuv2Zglps3ReDAlHNjKVgAS
DQKZNiiJ7mn7aP5xrY72CIAIJg4alOHZ6dEwOdlzT5Qru7pC3Tb0RS9M3sbA
cjaQssIsFolVMPvLV/b0FyIE+y5VbrnJFEUwxxVsGNT3ceaLNrWeJb/PvpTP
+Gg71gKSTDvyIneLfphw7x9iP5Y36EfZhuEkafeTbNhkWzPIRAV+O5yzkM7u
gHf7CqzukQvGRG6fDJiXZ6OkQHR2qb14jRYafgrKUx4K0l7uARnbcE3TPYh0
DQ++DQM/v1IqaYVeriSOh2YULVZpWKqm728Twd1DdNYlpqaW/WT1K58aB+Jk
JFLygmD1M8wCb1rXupcmi4Z9Izq+4dgOjDW+p+Vb7k9x+0Dypuzp7sakcweY
BXp2buw2Yiv0nry5ZypEAYxEtwuvg49Jvd2tyjnOOirLvQZ4dAJJCjPlb29Z
yr8a0W9AwfkakN1QMIIv4kb4FwDPr3VS/Ez9UGunv6twbrSe2rl68fohrxEu
VtadoOX7eKe49kpNU4Oy2jMOF40KFjYkSusw4/+GqGbTodyqT1mgf5G/RP5t
5KxwJVqnA2rGrIbRqk8JhrB4XtWfOr2wlk3J4am5lRFAAyb14XwNNGiQxtud
AcLYMaRsmv+Ruh+poPLBeAjkkz9e7h7l78zeJtFAX596q9TufQ5dBLJSWV7u
6Jzw8K6Np3qqqZVsqyYtqvuLERDPndr6ohiKVyZDU7wAEurk4795CBZabEYn
02LS4nrXCiMjchHr2j0aWe6adJpj8XJdYrCkQZh3frn2HtbqUOekCWRUYk37
WOT4M2fGl3rMyieRtr8Z7rSEIiW1yytge6Z9F2gPCNFnBhOmf7dE8QUJgixd
fszwT0bfbD8OLFVsFAwRtSvUS2dlq04hyXmcTHMBdC5M8QhBkFQGX8oQaCa2
vAmgEr12pwTGAye0b/jumo3Z2P2EbP3SYErC8lZZsJv7IqUTIQsXCnBoTEEU
/NvX+NrLJjpoRLaB6G5Rx7Xi2jXp7rR/973jU6tb0++iK74oOIiQAq9o69XI
p2fi/jN8v+5RhwSvnl+NBAmMy62FsCcw/6y3JWZqmEuZayQbHAE8ppBLXmfU
sTKwkpnIbeVnctKyNEV+sjhV+cixhm9nn0kBrzmHufEYk8SoJSRpjs+rz+CQ
1K8LLfuENOmImEUPLTnu9aHqLbzxVEqu/7OBdx3q81aOmD8D7U+7a+/oBAox
HDTEIxIt6apXeTneXyL+zrJa6qdyLeanqnqjbMb2WlgR4mv7GeEW8BYeYKGv
lZagiolLwaXwienVa2IsDSadRGbjzGxyTIU3kpF06lSypE4tUc4lja/hM0k3
nkNMnaA2CYd/waw6NW74ObDu97OkqbvlTefI1Rq/HHTGIWPuXZweXgyOUM67
Bw/CFiJMmobkR0fkizo4520m8rYJRicXNxZFNfNfAVupVJdoExDXIvr9Xu1p
Z1cAVWn88B0gXz3mEyvrbLoym0GVJCs5bRvYO6wGMEX89hRox5zVs1N2VUwD
ynWXxzjSgW9RpQkM2Kazi2DaeC2w2Q5+PuvkS20yoFZcbPA6+0bs6ntjNhxH
YeErN11tFybLc0m6F2fl0cJJZ9ZsWN2aNYnipaJzYqofH/FzNKKq6U8ySFNY
DCW5fPowNTmEUIrzjNooDML5p8q/pJLU6ryNWH4kHvVP8/Q+qs39AMixazwk
th+dgBZBzPaDuW4kiX/EymdPkEWVAhMHM8Skd2KAm3d+MUYJ35Ena+CvCKjB
uuSe1FNGx+sZ3a7BscrM7v15ztndQ5p7WfZNBmmd4nNDn8dvtjunCv0hPj4f
pMn3Vi2KPzF81Qe9HKMwFSJC7DLrc4dZTOHq9VpZjSMrL5AsteoocwvXw98r
82IK49yadH/rhwJ3MjkMZzrlb5D9WeH3gLvqsiGBIwlqWMYoRyNbh8jyCNB5
9oK1sOppX/hSqjjiXv7sGJftrY6yq18n3ND/UdnCnAZqkLDRtrbkaQALo0M9
4W0DgbCLtTP/Gb0mCd6P2f+sUTfeNdIjqZpY/XTKLkiEAw2AOI1dPgqsoHgV
waHcGYsNmBswgHI3abd+rTH4tD97YRSNktgsMaxhJNa1IvGTefx1y0hJl3BG
4GXZq3nx/u3NWtPuGlNIOFxaRVt8AScZ2AEzOnt7MEQhiY2jWAArfG/g4E/H
//MBB2YUvNHTAX5ialVoi5w8FOjnMcQ1iGgx14pBcKlmoxLCBY0Hyd2g96JK
uEgkWLg/XK5XK5aWZ3wTZwb+BXmyINsZx2CSdMj0gMC+ti774QV9TZsB2uDB
hZbVG3H77Kgd27f/5fX3Zq5Z2ADQHkYsD+krMxjB4L1SLcGSSVaqdMt3CNxU
UyY94XI/I+RVguaheBhoSyYTEkqZqF04l+nicM6spW3QEgbaVUUl+Njy40qd
eSGL/8BfGZYTwgtNnBi1Kso+xBGMyGD70+bGaqCUrPbHDUt5xvNa2l3lN+9T
VmPCdgJPPTO3X9QgkEa4mV7dgA5OR0bUmsDWwQjIuDygfdz9WteQetXnshKf
0LwHsh7VZz5vdWvD+bZ74aRQiGHz07Q7oWDq5YSg3t8revAC+HJaPZKtonUv
bGz4kCXOY1Q+YsWxuK0cyj6xIYpxO3o0EwdGm1U/RgYEGSN4QzVp1VHm98PX
B8iWFAVHNy9+0GJCM8Vc37+jHyifnN/8EbbXrP9ZmBMngtLxp4xRUAyNENjg
6sCIFphPTBuFTogYOUPEbY6jvWn9cPOQjRVutDu/3BycqN7csEcuibdSAvOI
+34HD2AGXcXz3/faznq98rM+f3iX8Fu82w36FyQZxbv12YaMzAHXnb8+rR2H
kL556F0fkTxYCALol2NQpNUDd5CzVn3iSaxIV0E0nAcQE4whBkM9S8XtJopw
gVODDzf7ri0i7NC3kIvoc8HRIOYOuCB8SwFi0A2YMcY5N4H+pzXmez0e5mfs
1tvNNVOQNNj2qO0guy37ALMsVxDCq5zJWKXuxzFDdrdzyC8CS1vGX0h2cqSi
ab7D2H7mzCB7TSc+EL0z8gahRsMfmjebFPN1AZMjASTHw8C9uo4fZWDGpE8G
B6taDzt1l4abbeV8MYa8yad7WPqz2dlnU64mqV7TICzYWL7hp6z2eNxJ6lyT
C4iUfCO+gqWdfA4Do1fKJxmQjP3Ffwg7xcw+reR32m/8QqxoG+4Z8okWFoJe
IbLNHHqWj6Hp8hBhAYD2EuF7muF2FYfYfIDuqtN5Wa3+rA2uIi/deOVkwp0h
B3s46amh9XoU8Hvf2mT4gDkmX3jeiPQDLcPe7duOrGheUzsJNzxH1+YB4z0L
C5mNhcqrq/ptgcA42mjSQ+6blCIjWfhq3F77vu/suRupPw9+nqhAEzP1ybY7
lWbmr4u57Tif4yxttqboQkv+1w9ZQHzVAI/9jgpDw9taC57PfP6sRc7zUJiZ
dgHtJdeW60wKCF6gB6l4PKTo2z+ptABRBsSZA+hjc5DhyMB7Yf01G/V7tPQo
QrrA6KtBPj7RdWP+TdbxW5TNk/o6WBGxcilDS6yMWRFijH7MOPgCA3HfPkry
8bzenaLqoVej5L0apftVB1jx1hz4D7zHbBYjWpfWVsUj5Q2QxQ+hpt0IWLA6
GyFI03E8TjikIh6J1lI00mQwxsSnHgBywblj9N66hJzi0ITR/T94+OWj+8FH
9R7FSg6vmxLMm38lvGsOGZvwEWl7/F6TbmqA7iDubDtwBmApKv6MQMk7V+zZ
WhepcYJECPC+27ZNoh96JU5BYYT02iUXhliBLvxiO0NTE6wpt7tGNpWtJfBB
KMJWvlOadc7VKM9mIXqQ3VbmMFc8DKRGxi37UHl59RQ6s8DiYbjyr4e5LnJ/
4+tdUOFT72TYWxpJJULPjPlZIz8BKkb2/BM7GV5hGLp0RBk7Gs/OQRwqPcXS
RL1gtp/ynU4Kro0wPOc78GpNg18iZGEQjSwk3Qo51G2ITRdjR6RHxQvBdND4
tiBp2mj5Tgf8OJMm4piXylG9zCry+Fkaf2i4SIzEnbOO9mVo4X5jNVPhw3f4
buZG+8B9mu9MGRDSAqAo8iSq+aX9DrDCV7lhhdUhN5AJapDGg5x0IYTEmCzP
fwf5cFiWgvoF2qHfX2XJ+EaqE2TnuTU7fOIsIGmpC9K4gG9rjCf9ult51wwy
x73eRj59pQ+qBQYDBX3x5UNZ2bNoJ3iMGOg8ZE7DpB1MxIfauRhjWX4+POaq
TjEEpjedNc2HI4K2wmyVp6gOFtfSUfUDVc61TOurVJ9X8jYT9nq/2dkdrf8M
ezKCw/zOGU807iUsFV3DwvABJOK6KAu08wBsCfC2fJ8cOASsqZ1OXyYNL820
nlQSWawJhGEsZxOy0jfs1fZBUeq8AHdZ2DAqjnytG/aT5HPR61wPoyblphAD
UM/Lvds//xEQJDTDgs6wvMJWhasuSQ4WoPdAnUZkCkRmgADfovQ1U7CVy/IW
5965ZIT3M71m4yjw42vCxXnpkTmmBbpODYthak7wj78gqpxjxsvN9tqs/OsP
Zk2GNtQfhVDLXXCxDfSamd/4szAcoiaGlYIWKhNm2Qk8ZLFiyQyXs32e/4fs
w/ESNnRifGCftOcDL6cjNTJuVHrpSHoxyFifFivwMlQBEnlmz5qLPXqO9PPo
HeqpgjhXnerTs3LTi0vgdQFyViIY8vzDpyCjJVh9TUvglsBSWyf59Oi7byZZ
JtsD9fHYKYutWsvtYJgImoO7vurt7MqulSCHhiCJFhyTYKqxlzFQqmmeMPep
kpu3ZJxPwkSbWgcvjubecasZlx+sABzFR6v6AhtUbFkJWgfMMSzwE6DcwgqT
/nTmbvV/LswfVrscpDMeAukQKj9fgQBDUSf6bvmiKJDfflksjZt/lPaQ1F98
cLLedl/6GvAQQ+CSmt4NVg+t6B99RlLo8j5Kcad2ziSipy0+qXY16wO1dNYp
VZ6uE+fn19pQlcZ76XkHAF/mlpS2NSmgC1tqr2XXj2ZRtu040PqceI7laFHd
zwm4Nbriu7/j8dU3xQGpP64qLNIq5M756ofGmp87OY1y45oP41UbNMyKbkLk
TZaDRCJBheokKurxZmzKMRZWc9I6a7ITONKe6mO2VwvZZ4z0R1BtJh46LQcH
rDJ51SE7IbZ9jH1FpAohpcp+o032rGiOd/IhNQABwYEpN9TPa84zrGjbS2kb
l/xVi6JdZ0uVwJD7C+VvZiqEZHcFIh7H/SWx5GRSnS5C3dfh+4E8/UVVt0K5
/kdyB3b+iNxfFqIHSFO8xyqnh90aVnIYjqhJOrHwhSeJ2QoX/DnlwmaDJifo
iRcNreNwuEnuRdekgewpSMt+IP78ycbEAUc8dpIT/DguFm5qlkhATHs4DlW+
nLHgYghRTXM8vlK2k0XQdtaZyPNSzaQk9I+DEfQXHGYmirs1YJcmUK991BXu
b8xclEOsgTxd6biM2Ta72HuPtp17Ezy28/NCf2tpe6nHSFy7mipyFSSBAqp/
hHknGp1F2/OCF0x5x27lLEA7jcNPMJLWnH9qNtpkKip1AozSRzIuYzN4fTLu
6VI9/JhiEPdYW8NFaKlP7ORTQIIBsL8A7VEa6YFak88WVw4ME9FIDnP0xUOQ
PJsCgymDGDIAgy0Y5fnR2utEAvs/P2U2NOHfxnrwbyDptTs/ewPHAD2GWnNM
gxKGCoRghQ+SnNnI9S0smUNNYy/M1D9btJAZE649Pwz0i/s+Q0uaZCPkaRmg
nH4cvbbqudlULSOedS3igpEvzS0aF1vK/VMe8LY7BuDy7v5SfwTADZrEFOTA
EMZ7fDDDSTy8Kkoqf1MO6loqujF71D93nQ0mMhMkXRF6q/NkDTXXFpnzAVJy
qkYnAejWa4SZrxkwhp9S8UpwgK8AQ/NJOgTIpU32eSRes+WVNxV3N05vfmRk
ETXGnnDISPmzlNN2AEVVpaQc2OgTF6xrHwFez74srE84Hyams70dyp1/CVGt
vG6DUAEXfBio1SQrMB+2sJbYoTyGNu6/L9Oo3Jt1h5UxJs86GS5kF9dO1s+8
jY5L7ejFWjOWzcLmXUxkEH3Bez2BULgZl0vNm/dzuh6TtGp2wSL/M1SqCbe/
fnzdeeGCTnB+xsu3AgefR+C4RHAKPyhL0xLGiOSoXSn4c5BttoY+lteqe0yo
sOTJy7zGHNLEqA7EofhRsmf+WybkiMpYH4vUA9UZegCk02tK1iWa73iwPd61
w6s9jpfBxCFAGgOaUsoQJ+8LkS4QBb8YFzMKzyAWQxITAqPSgKf6NpTJEC2C
KLjM1rlpdg8q0Y0TRDPVtj8OUCAAps3kJfNA7wTvxIILs2ozctNf/J/kVuSe
9qpgZ0zKdJ24Ds8is0BKuzWqPD7mNRB0bRVLIvM0op2aYevfW1NABBT3SXn1
bKlPd0i5Tmp4oQXaP3QNHXk+8fqtjDjYc+YqiW+QBmYglGT8IoT0NR0h+MZw
6/vz+nKAcrNl3a2hpLWmsUFlKgeFzVPw5DsSWybJge/JDPChWt367sICYTb0
UuYqj3NdNOqG7KuLlQsJWiRbZ42UMWfLuhhCH10K50lhjRJgli4XU1M4w4sv
nLmHLPt0oxn75Yj9O68o6cTadsIm+h2vhF1yQ1If9H81buQWxTT/di7rk2aS
+B6TBbALtqlKs4x0lxEEurIsDbtYmOZ7Sb3ImOfHKgEk7PWnGFnmuELQC/jK
Emwv+20c1PrwdvxyvZGPjQ7gH4FFc8+VSaVIbFMGQXlVuzYBjYgXqPXz1vNg
PexmlQ9w9b7Tqgk//40JCCYNjj73Sce6dxmZA6O4A3A/A8bT17boElchLS/D
BPQT05p/TlA082UcsD5LIMICHKVhJ8Dg8iUxgDF4VifuDisrZnEhJDasO0ls
MKr1vAgoTAphlr1eXkNGF89OtZeS7CWtPjT8o1MdlhnT3Tc7QD590gPx5rNi
X6GCjZFiw3hNQbA9u4xAaLoiygSFm+Jh/BSvlmJFQey9Q0iybbX0J/Y8uLp+
DyJJ0tNR0G71nTF/WZlA50CIIzKLYC2/79R6zSlA1KLyQ4aiu1C/U319U834
dKX7+ivi92hspFLO/8On60A67bHXZhCGSbljaLvBg/cuY/RgXFii7HlVVyRT
QSVcVtlGeJqsuM7BlIu8nrFk4D2CBjvBqvWzuyM5kGTU+/vmdsa0fygCUd2S
qCLz/UvTcStyWMlHKk2RgOfB3iEnxKjG+3KNM3iQWEcICMbst7Wmp4XFO8J8
jYW9COhV1E34c/DhsSPcTjgc8hqLCv5ROrkSNdtLFLJKo2Pmlq//PB3m3cau
4TJb19c0bentdeL48Eshg/Ay7j+4K2Qb2kfer4zFrNOLHmVr+F09eaSUDJJk
Cd5wpELNwsD6fJIOOmerqNS4nCjdpyePVOd9Iopvqv7/5sMe0Y7bfG1rLhpt
0Gh/0kyeUqElkdy9j7yvHh85Y8DqXXEQvT+mMCkBJrIe7tU5IgDrndeYaxSL
t5L+d4D4NkeZd1I+pEaWZxmbHZBuYZcu16OsjZ4fLsfKUFFwC6dTAZVLFhPh
jwfrcb/whqAbQbEuSbUrIHe4gP8zniHdOF8icwk3Wr4bTbkfngCS2dvP/539
7D0dW3FywFlfefrn97veQkI6EYaiFBt9wAlv+Mjq66aMlwevLu6OJQ2g6ahr
Qj6OBIDzJFvLmJ99funDuK4Rkf8vnfrfT8jqDREwuv26QsY3vrOal2wRlyla
+0qy98F1QJS8qxxaXI3lPHpcICkgk94w1RI91bBN4vZ7h8Zg440QKUkmIh3C
JroEMQxXwh8WGpPmAYosiryCXytD5pUUPzF0VduQwftgflgZFtJDHmDYkTJv
HWFa/elxvwPcG5P4fuwd48B7B5Z0EBuhQZnx4ds4qprFoqhbr72wZ3I3EG09
EzgAdby7vsK9jrPqLkgYjeL1FWvdPvVnEP47zpKT556SfiMFeoYN9pqNwVlB
cF908ZgSwHayGex74QivxwYw452cvk2Oci3l9TQ3DXwkOdZQ648Raz0sMWdC
yAs/C2MXHtFr/pXIPPCoEp5pJwKiGESgoanNVczbIUGolruBi/FbqyM/XaxQ
Plq1OvPbrvvMZyK5duFXy4KKlwTCs4EJS6sqTHojR8snd1UEsuhy0aWu4LkF
WHkQqtgxqZCHhiXRONYaWNv9MZMSfEzq9IOHyKhc5Eswt5qHtzKltgJGTx0A
b4lDu39ywyMjG26ANcJdaiHVs8DvbhBwx9UvieG84rIDhr4KDj3bop3R35U5
gwMTflpJZc0hmXB52ULyYEG5KqL/AndudWn5Lw/kBYVb3ab+PrKWj7Xbtroh
twDWvLJmxz4jWQaRTgyPi+8ddiBGXg6ZpQIggcoSyIDYspKwGmFfPHXA+BcH
hn3vunnDQwN2z+8lKf7Lrj6vkNputdUyA4UYFy/lLLls6IwcMUpd38XzHbwl
FTf3kTfS/5uDpfO2SOdvRDS4pXA4Y8I6SHMNI0BVtHO9gchLyF4MIQO5N8Hj
okC1g2xxJJ1R8KZJL/DJ2PTa78UTnWNb6L/5YU9nczNpgN9byvXbAjZf9J2M
FbvpmL7YO8om8YG44wMql2hjlxHtWsaByQ/hwGSDcdYAl6ajLfZRRLQrmFID
1qUZcLvsQDDVm0BwV3V+49C5gieyrH5B3p6T21p1hH+R8/+gxk+LB4/HOpb+
zbAvwn4xHY4MbdOMdK5aXcUDJPPZJmSFeIjslbGPZjn7qST4DdEcubEBhNF7
iKAPMjHmDjHrgF7pcWFwi56SP71oPxqJeXuleNjRJnKThmUFv3f74gS7EhH5
68asyWPg4mbwgkjLSipjksMO4qiohfe2PbbSxnI91z7m+La3XRTCf6Ke26UW
CyyeLn+nM/77mXzQImtBMxhcybSit3Zra6u+xA4tXrFNxdA6dgzpmeZSa86h
eJQAwydG68Gscu73DAUABT//H5tsXrq03ZSxlp1g1DxKEI3ybqyUfpxaSfl5
GOVoA8BAVQMWuJ7/qJ9aRPqDERzg5xhxbp9B8A1OqSVfP8A8cS/3e2PSKiN4
XCPbaBpfqh6mMkzgBfH2RU6si8JytNT4cCNs1Ue32N9jsxhPaVs0I5xRUmA5
7f6zwsp1534t0a/BSWaWmGVtFkGiHrn/+w0syu3QNRjtl0QwaVt1Id/imLaz
6DtZ6vJeKU2HJ6RCVur9NOdPI2eA7+wqL6LMhvhafcwbe61pdzCzMISHm4sI
4JVNQe5hpw+0nW203Q9QjjhYnNGHumZ4cC86HMX4hRCpjs4CWUv6B3k1Z6c7
Rew8THKfFOFYgSiBZnTRZYtPzDZ5Erxs3nzWJsg80P4UOE0Sn6cAvZ7FXINz
aTDBEEZdRJ5E3pehE+I9Tt6+REBvPMjIa2vwQnXEPHsNPA3kYUs56uFsdf02
X8p4cmxlM6Wbpte85l8ILO/lejaS/W7tnG9d6sM/tyxqi/wdSrF8tXLFsD3v
S0BngPc0VcNCTO/KkmHiFh+ZzdeiovFA9J2sD6QwY9VywWleKd/0JJHsfnzZ
wBYeR+sSjlDXd3J19Tb3IY5wAFBfkOkvl98Oy8Oxzy+0UA/FkhAg9v76IHVM
3Cnyn64rwyXnXWQqRB7HXfDKD+etFWBtUBq2C7OxZGtC8VTJxfii4C8UgBPP
0jiirQPMTAmNZIX/8cersdOanqL6NDAjE25S+BnBBRedIvljYFd7znXM28NF
F9bg0+d4QnTLqvHxrDd9Gt5YKR9BjL+0gGN432xsHwBb82/RpOLbLa2rJ9vU
ZI5saKnjCOvZc12A7N9sNx4uHsmPhVHcRk9rulV5GxD9qUFbZkbJEwHZ4bti
9I2KCEZjIhshDsmVq79v0t0vzJLiwLfba1YXUrdVp0wLCLaObCbHhHCTjyRL
eLnRtw8hVWGcDoAMszK21HRHlckucp4Zw55VFmcIkdf/GE0pj7RULko3izXh
KQo2iaOfk0eyhoZM22Qp0P+tU8v4vZl2MO/P6NSDthHcD0wUXvijcgrfhBPg
x1qbWeZWbzBOwmfolLJkrH16VgikxbWyq3f42Aidx/67KoWEx/I66NpLcVIV
hcOLSkaqhv/ili19svFYKAkI+o2MXAmIemOmI0rTl8zya9Sqq/waWrxG3cyZ
SQMPRxHkscxD3U+Qki3+vxo0age+dmZSnZC1zoBJmGbaa8068fmIcIkJFNok
IAmbsE5QUaEl0JNPOIUBM5VwLmvctAsECrQqcYAMFukNtGnKo709rp+mgPP3
XcPlBjtRJO5lohJqE5+hJlpPPWRMT4w8fgkQZ3yPHHniR7LJn/tJIrlMMwZN
rNaQOfIfT+xEXMoRbXTOsLXtJNl1Y+kaNe5bZtkEygcgST8n708ZiiJhSner
DHM2MZ9voRYKD9L/NH+MbAGhEaCN+E+tJpnTx5pyVitS6JsgHvcF4o7RYgcH
90W12EJIe8eolEjxxs6td59ZguyvhzYhxnhJbZdtiMQ0th5O3C3/x55iJqdF
IQX4sSHKWLc6bEt7LudNa6NbQbo4Uvn/HnGQ3RInz/L+BMJnquCz0xXJjqJf
dL4LCU99GSs36YDRJl375p9TyuIAi+MgjyjfInB8M7VuWlq5vdbVIA0L2Tpn
YfUfg+++kv8s+JLDpbQ+rV8jntkkyq/KQEE3FVKFIaLHR7vAtkortSVvJGUk
OxbuszqeDkDD17K9hrVtbADxOGv/PiLoE5h4X5o975jGHS6SrXFhbrGFuRf0
r/YbHHnymXxgSwW8IrI6K2B7/3Kk7uEeBBSizx7Z8ixhN7E0ZNkpr6CNw205
PRiR2BDf8Y+7C/ZPUnHEZw8aOr6bwIu8DEN1hr0LRcR6Ty3JAWEtkWfhiNPc
xJsGmJ19scZbxpnvG5yqbMJ1zZ8aZ76HTFNKdLbjiqMpFz/O197bvcxZ9/Xv
L+mAk+FHI+SoBakdX/k5Zk0RcT+A8VACuOJGIpDiFexwt6sTFsLVYFTRgSc9
WW04vT8X2JPqHKlfdPkLV5g+O6YETLB6vzGBArDk0pBFmkMIiF9lLj/JdS3R
7Xuz4wRoEycCWzJWKAUgFCGJU6ISWHNlOjRuAg4uWNGf336k5JSu+IfhFIMK
ruEhHawUfGJFo/NcjmR2t+FS59hGduQzPglW9+3MeJj6MIDQF8PneZmp7r11
fq6uVgByohD1eDzADU6yBNNjZZ8NBaaX/ICWPLzXtBNSSdJRmUDs56/oamH4
/qr5jUdR2eXX1JmWmZuchIJkYsM41oEf1Q9spPvP6E9Kvq2Fqf2GtTt5g0/y
Y5y4b/CMwWTYemfWvxE4TgeQp6pqweUN/9hgyCnjGyFqlEscQrjnWMEQ/3NP
uyIqAOILY5iqRCwDX9h0GWLPpOtgbMf6TRyoU+PwGdXuckVBSuzWP7HhLg5R
7qC3eqagKfiSjW8Ec0EsDUw8BQHRsSxNCZ+Aoc1UlZlQdtmJQfU0766boPNz
5sNFVdcz/sySlyOCcD2A/kbrhpgBd97ypDMsBaK1xY59nDivbuE6D9CO75Hz
LA9TuZOFy+KWFKYpyOr9tTsUGHYAXWxvtul8WVx7rp48NnSt+5tQ5GOvlr+h
BMhxxmDpVGYEJMnJ0gIMiVHgnliZhs5uL+0ZWCgcG/Dadeo8XlYezUpMPFNf
ydpZXwZcCujQViilhtEFs5XG5bq1bE4nNGakjCE1tjYJkHAu/CP+89HKkVnF
kBx6b90XzxJO9MLgddohEhRm1xlwGMMRnLsecE28H4CWweUpPeDoKwvXX5Q5
mJgyWRU4qbx241P3tCPBL/BBFT9tStErf8nDp4IV3EKEkqMHjsvIBpNTmeJy
OhP6tKvSCpeWBkSH4F/M65GX1eyJgEVGi51U593CmLoxKGJBI3P5HG/9P3v3
q4AM5NKfDE0BXe6y7b6RkAjUUq5FXC8riODvLR2dYYCD+8IvPd8iGFyCU8I8
uA9Owm+60Q1VRzAizvXdIDw6bBirSx0TlfwhdFlc1uzoBp+WEjWVUM7F6D62
QBDNXFTTRXoxmvYQ4mtHg7hHMmJy7aHSJrjRzRU3hjCNaqAhmESv8NVDmNyU
X5YQqldo4NICsCW/LI6j7OvFb+C/KgBGgOM9LXuLbGSJZ6GhddWPDb7VzVSh
dtBfLqAuuxKx3odim4jD62m3pxuEdCui5dppwNS2n1bHTfJFqYioQq7mEOuV
yfmgIhajOASZTyMR0qSq/lnsmvplWuRo9z1tRZTEzUyM2MjtNaN9VLcRvMbc
R71mg1UAS8kUHeqpxA+un9FuaDsPdVQT7OfiUZyNy+HuSpYY1NTxjtcwAnm9
kJTqdTZAa92xqQJ0g6gBvWKo/H9R43dWDNbi8jlfx6mOl/AJbuTocqwcfiRg
uHg3CcJvX0mKV88cdxIeaqmJLmOe+VtKnQSFZiJ3CAiK5rHiFk8fGDExJ6XY
VYiWahb/v72HAfnPYnNVGO8PZepkCCmx+5cwNXSPlxdZHpdxc1u44H7tmThg
QuBS7jqpqzT/zwcHykZv96UVV7K31LbqxyzJxTsq0B5W+vSl507lOffnARIJ
vz/8uU7sE8ayA/ltSUrhT0aCaR/pS9T40ppKMUYbXYXsw0PURLf9XIN1Z6P4
1jMtLvRKfMwg6dOC8ml3zQYcPTlURsYdY0FQbC7iJyauFFrshrP8nc9+8KHB
ug5/7wGnB3Zj7YE2cBRTHYRRvllbEVtUo2iTH1y6lvWbVJBP1IsiIcwnpEIr
CUWYLfMy4XIv4jZJ55iTXdBdBfZ6gdJ1JxqxG9L6NkTvcRKRuK8a5nf/ikPO
8EHdAvyXbZtPCbTm6IoCQg9Fo3Znpi3g8oMBOYKhCxsSQCHjMwO1kN2o2lN4
Hs2Rr96JmMuQudJ8Es/q08RjQPR+TbA+OF1/krs5NrC63VIPuJ8Y73TUh+fb
ZqstVCyvE1e+OoTNdhQcQLa9A+G3wUAc2ZWgLYm+tWBzMb5Gr5Zi47OxaeVR
tkohqdjziyaSgqhLkCzcelI45IJTMfEyaiqE4nmE9CyB/3Sqb9G4SDB7X2Cz
rGcPhkCDaXZjXKkklTH7rJGwzZsbvHyh6v/12WV/q7hCNMYO1QG52nDlFDIo
asxuWBwhubA8yrbGUQH7ir7NRhqLxsLtpgMfPGKrngp6RcHY44H0aeLLv7xS
j++774CJZWFF9BAWxFp8IeLUek8sEDuBhzxNkJ99fbIA6Aa0U4ylTqxA/oVy
HPhcm12BR3aJvvpDsWusCXfAv6zgwsdNKj+sSKNWAFqpyydE2gxUKiHGlEvN
hnGSCJGc0ZYIbAxb/g5d4ayrynv7CTdH0bKYJoKjs+RXYUX9eR0lphLIbKsd
uUuMfXszhV184I3rfBhPymLUeICvj6w0K9rinW3Dx7go3na2k2SNrKg+4bP0
Lz8FjXxXuM555lujWYf6j44/4aFlCNwsFwUzGqbDVE3bSj9y1PYdDKdkiQ1B
Qr2QB5mRhO/zrFO1IqSqBh0iUsXh/vRsqz7/ntiePb5rk4C9KHZpfxgdP6C8
bCuC1Af8nlJyr1y+DpK7WQr+a0tQ9KzYbPToNxZKGnsJGbQXvSz94W/DsVT3
cpxYTnfT6PjYiZDNpl2kyC26+zsNo3YL08w9stZfwIhw1a9p2BGU8/Ce6UFN
8lab4N19YnJG2qxlWX/5lf6uwifs27TVKji+zr7Oa3YLPH11xqMvY53DtX6d
SUpddncpPPA1ybiUrvkKNUY6CqKiGTJ0eEmUH8bRuafkQUTUTg7uE1T/d46g
fNCE2NYtWwv8xXSrGIX0dmCuUkdZyv7aj0aZO3gSY0jruYS/Gmb9/cgFCfIu
6McC+dPJXJRQZR4SGZIgcJse0oatgJxbyY5Vl+ub8lNkD4w6+zlDNMnAgbPg
Lz9RM7frTw57+XpGi7qADmaiHw1ShGALrejkZhs82PyS1ihgR5m5+qhs8wdc
N4v7COCemdPvh7kefHMcL4aEUjylaugXqh+UV848SHPDr7gJrPFz4SkjT8iy
4NB/CDqFBN8rTsmdTWbEWIY099gZdu8yklUS58Qyz7w5CL81OSBaSiq4H8Ds
vIozqSZoWYi5ux6bKBNnROs2hBTSQXGFGWXLabiIhes/YuMpJHWAs9RpzTXH
oius0ttiZOv9tc1ceyVrJcRUtCPR/CxPgFyZeX6hLIJ3fbJ2y//ZnWnjbnbi
Lbew992TMfi+K4k2p7TJEDMkmKd14FtGC55xcpw/6p8duyVL8p/XP3JGFCqK
jND3BckMt1mBNkCgMtAg+KYGUwAtM0NQT5yIQwW8d3t1+tOBn/adVFOE+925
cWDGYYrfQLxPRtJEtCdiJcUMwnhOj9lkDI67g/rEcoxPNeH8ejVzG0YV9Sdf
zd1aam6ejPZtSH3PiZBVEfAY+F7D+i5RXVGhVuj1sPioZWlO3P84vHKwEJDd
WPfxFtrMbd16E7hb6BkjRIR5RJKjrYyaW8cEXLBKf3L0IZOt8muHmtzZ2HMz
7XfW3wKHEkbKNh4roDcBCQAdY1dWZ6Vw8yLiInLwaKrgmE1U2t+3kvkFyLxW
IQRrq9Q2TIjeeRZFXzb5RfElcBk4zAXwdviVRWBt4o9Wc42aIQvgn/VSn5lL
88dHMV9DXiaAJ6Tler8ucfnb8NahdwAyumLIeypTHRUH5pG3SIrVNLrpNW7T
9fiQl7YA8+zJLwPMOpLW0j/vtMAXxzYQkvh0NwzqYem8m0m7snCmAJfmzws1
0tB6zpcZqsfcnJ7JQ8llKWR8R/Gxrk2tVNPn2OzScIy+8iMbVZVCTugfsN/S
pJuVmyAhs6w+2p8q5Ews5zrOd8eVan1fhCLKBZz1iF9DQQmYCDrNxr3yFlWg
JdvhCcYzwfw5wEW3Z2uo1zJ1sCAA5Fris6Ekv/hJ8WiTxJLnPAzuNr8YijGo
J/v4bD2MdxcqKqP/ajqjfpReZe4Pzf5MqBWJOrKbtxZiasl7r/KUffZIzCoL
+ebTAcIOId6CeVezsYiTq5fu0VLizeUgQb3bMHc8rmyXTLcJny/6e0pOyyY3
I2sSV0aQlNA6nYJFmYm1UBen6AEauAMSYbiOXFI5QHeU5/9G9OzPdAkITD+n
2XzsRvyayBPayL2Umdb+ykpx8fofwwKsCMSAopFwvggbImv4ax9nqDHak7Ao
8ervHlzFh3iRoRJRKu9OFGaKSV6lCgF+v57nBgnL7Th3V3XvxEED5mo8blP9
4cBTcCbdvJjfkO5XDH4IjdGJOiXovnQifv3vjwUg9Q+x8x6o4G3K/0+8VDrn
g46UqIiEJEdVWXZ4KSdKKY9ljQaKzHQxsbndPu4jqPH+Q5Qz78D60ciIk64X
MOHfscd2vCjc0/EPMEss0g4r6/hQGsO8kbH4GSXqoBs8HFcWKWRuGx7rMJmW
TEglf7iEg8fQ3qVwggdKJ/StYODbWu4bmThDlExF7plrHsjYsn6QuJfLvHWP
xXl+l3bWvKoiHZ0PbIEcJC1Xo/uCoNvH451/WrVyFsqO6/9J1JdrE1wnfIFU
oLfuO1wed/vL0K4L09IFCyrKc5iNyDuoeauAtSgK3yyJDAUU1FdhB0cL2Ffi
TnYGb4/rNdnEoskMoFQCapZHoTQMqTOPini82W9WxOleeFSDF6KasR2AvxGF
Cpit6my0Cm0WQiBTSfU/Dedld0wK6/0NqnLtTiv7M/l3SbFvQglX/WzsWZzB
hLiVNWn4R00qonks08cRJdSSi4DEjabpTnKPQa4sxHb3vJLag/at5F7xM+HM
iUcSMgbztXhcfRVk6m7Q4M4K+bNP94wBtDPjDR7bT0JHIzMSz2Qn9QlRCR1M
vJKUtgFhm87S8MzQIyjvt8pZj5wnJc5Unwoq7KIsg0Zxoe8e9xUKKhQAphF+
pU1ErfA3pf3SI30GRlLtpoVq5Tbu+A9o9MMjCaAekIZB1D+gPtcPeyNDrvKe
/dGhhjg0m8wgtEGPqWWrbQN9joc3nh0+35ZRl5Pp26K7DiwjqspAMMkWrMdu
qfsvG3bEAQYug3QLkq8/gwnl06I7KPf6TSfUax4y9jHnD5qN6ogOP7tesGi4
OXmg6ObJi/k/fkoBcw08bSMCNskIqcczkZEdtKMqif8Rgxdo0d5bNyI5/ks9
Yb4hXvWLEbER7ei4ZFPsyuD9rz0r7Ds7pce8bpTWflHrCSu8NaurrFr9TkDd
uoBWc8pa1CGghUgnrP0Tk/1LNmQaSyaY/MRrNcTAi6NkLl1ieHeh0q4U/PbH
zIuCIEaqCAyXZz2pG0BP1mYc+HO6Ydl9C653U7D2GYRt2a1X8nprDaKw4MNG
59Rt0LmphoHs5rxp1NwGM0MO2dE5AvLJUQ+1OMr+BXmI+1Ds6brQDHIarf/+
5GeTJsHgQOvvqhujhOt0+rEzitf6ySwxzNPVBNJLUJ3gOunHATqaq/Nh7Jni
hKJ4CWemJJvsntGq9tAZVLYYlKvn4Qr+nCjLb+kNvxWEyvdGd8pW4nsxpF+1
VRqDEx35swmz1JlNYPNv5Df6HCiY5SOBFInRvXi9YSrBTvkh/5kYSW+ISX29
eTZxuO496GQVeyCRum7zZTYLR/NuPg07ASX9i/wBh0WTbb4pCTpFKnilYFti
It7heHYVzmF01NK8fruXc39Am29fCXRHJBCQSVm9llulVLFlXU5l1Z+9KoYG
DL4wyRF8MIwwirkfXvd56ZAZqi9lI/+SLp0WHvC1uOGxohSRFjzEPO2w7Tii
WAMPHGsCQd6vzl5i1N+CFdlAav82Qheqc3j/p5wmO+tkHSNegRNNwxzXZ6/B
g88960zXQSm8TZh4IRswiXLv9G/FDQhna2hpliz8/S+oUQPf83mvos1omBk4
FHwcfxhAADGylJVTsZ4KDioPHDU7BpxxBF8eGBuvYiE4KsWbnM7QQIXji3dM
5gPWSMcH8SOZptKDhkGMZYTKg7UFq8q1UbmjdaKi5MDfk1fKxufcVOUIefaX
kKA3zftnZL7JFkJCApf1Cy++35nGHjbxIvFKIrGPM3X5wr/uzCDF7fzFWcZY
aEVKtq/VtqI9ciSgUhlJKTNAJF/RyGqYxE9oMIFNW1C5av6SoVxA/i9DCPYv
3uyFZ1FoDXXoDcJ9crPte3z39TQn0tFdGP26jcdWaZakiqk5BItJfF1dfe4L
cl5Eyp9GDt0huFGgCZwVPnILou6m3ATSIfAqT3lrc8CObICPLf4PnF9Q0mRt
vf48gnqv3pPzquLsQmUq9xOi75+xDMgKWZnpJ/5te6SuLTbm4WLQdBaTbL0D
C6cn+ajGhn4jNkaebHrBYS+nYM2AOkXMonsi8DswYTuutV87gDN+o7mess5u
31V0XcSa4LZTsoeGL8rgR0MdQGytqJ9ekB1wGIxloWFHsowrKbQAnVNSmvXn
R/BPTCPfzaQ9FevblC4yH4YoGj5DCrYcoqvhFjkNuqEiqbSpSho5wMbQHz1I
Rt+wDdVVmLiU8I212b8sFxkCsSltpG7t954jSOHSs3o7wI2h5xKAeGHNKLYm
oqqaZl3T9/09pPna8Qnz1CcgW7q5Kvr90aNYuDr61CZm7jBZRBQDDbA2EpGm
4p/yzx8KxGW7nkJNDjxAfla/r1BJHnMoR1HFYRq+Tcc3NoSpIduMQQqzIzlF
d7W2mUDI3gBNXplLOlFxJoBXNoxH/NjBv0K6/+PcnJSBLTQZG9qRy4ieSJgA
ALubQx4dZnIoXJxT7zguL3w3Dv8bjElA7rBucPyUFi8fPKbj0PBc/BTrEDQ4
xXDKn0faV+Bc6D/jDBVewwUUCr83MQsBSP/qf3YUB3R+/XY16D2UqwG2WFJL
QY2lhc6ae4WYZPTwDUt5+LkK+QYCZYozDb/FHSVlsDnPnFr1+gWHDUw1YZ9i
PZOjAg2ksvIRzDlpUtVphowkJWWlUMCqVzt4d2Fq+FWANjUb/nD/J8JDd8dy
JP1yHBvPObt6lyjzAJkvZoFqjZ6VfEMybadpFJN/DKyIagQn8JWLjDDOflk+
LqgI/+h0MTUdXRE/H5l541P3gJZjSxt4dPFAOGc8wbXL4q5QXcVqA9L+xuk1
o5D+aVnKQ6jvwySQqRvCXXN6TReix0X0dEbPSC4kCa7Uu5LyUxKpq46TtsQH
MzyGwTbEkmbG6VMYwrd9Em7RKRELvDBObVkJKfynCOm1hPpOLDJVXWSfXxXe
BGkQAfh6PIGzuxSwEU2wwErKX+JJMl2HRXfJz5Hbs5lkTgwl/z6cyIyPdCL5
6IvWo9d3nUytr7Vo9/H6zfWcz8RXmAPTRmhStgfv/EYLT17wqJZBjXNoDStX
PoEfPi9SRr5WOI1PQBg9rGBYh6YRjMNc63c3UqrLwUDqaviOK/Vn0TsLXJ+F
yW2bU/Ik72s2symsL+JvsX2A35FIUWfNA4gH0VNeq0Pspn5XY0tmbKX5KZC+
Cze2h4j63WMFqg4+42C7RpYok5AY2VkEWwku4ev8EkajQ4zcDytQHpIF+ELk
h3oEOnmRAfF3DaoroCK2wTfc3eGBs7WV0rYLW9W1cfyv892uykBnCzZu5GQZ
OJBDZjT6BG6GeJc0wIbZS/AyWfd/VZEFcdi84Ql1bo0J9KM1u+VIxK5sSISW
5roZe3qj3G1gKox0HN0Y0tJUSgTL+yqhWR6552SmcuaDeeokW0JDYZuWdcWq
CmFox+sYzIYNWU32upU/lYKwtc2bWlzEsYi9iJONECW6sTdPyfANsoLjaM6L
I4dBqrHjaUffsnaCmIv+N3BQokrCNkxxSHxn9UlFZX6t8bjCa22Sy5W1WWht
RyAdQdUhNgC52T85wXgeompYjCnFTJAZDl0S+XhGk/YJbNQNo5F01hCOBg6S
3DjRQ7ouvqlkhxuygimp7KkWi8nbrnTlMeCWodPHXxI20KhmTFanhPQCBbe0
4GpNjOdijh33izbIdDjZAOx+/hOB1gBu/nqghZOOIQNETrWGlg8BLWG+8J3J
xo97hooLpb4pJ6f+I7thl+y1RcFMny2Nw3iNRqldxP5bQY1Cq3+q1KMnNWP2
Ea3sF8qq2+JqdduPaZ8ng03xTZ9EVxb4OEWX7StqCDSy8wX7WdF22qI7X9P2
eiX6GoFXV8PMH1nXZ9lZh1RikOCZlLgth0qXFxarpG+LAdpFEsg6AlEeQkL1
OXlakF/2LP5ohA/G0WPE247emvB+j7ImO6R68Lkscpn2dFKWcFjmXfI1D6R0
DtpQB/GKUqxuyvKR43I0HQGCuO/53XNpslfTuPxVdmM+lS90+4i+GRhyPU7i
VwgIcCdxPDGo/28bG/cW4Y+ZFNtmwGr5vVEZP0H1UBV3WyzjqB4yXXzMFzr0
OWoYc74WXCmOrgx5AzWmz1toY4o9fotDLRXvyppJ0nRervldfnmcW7TeN8/x
wGphgCbs143o4tkL07CMcYTzMyPIxyoCAu5OIkBuP1DqsNXq/hCYJMcIwc3X
8Hm1Wplzp/YiSeOrTUED9fSbM+1d9KHd8GV25pxlEhlyrcwCtGc3pi8dKPj9
wCUL7BkCK/R9lVP/HHhQ7IQerxzRaA3OqBkoYuIG0c5XCCC7TStipiMZInLe
YpGmSu+iGPUaSVNSqAuvkKTqXDf/hpYFtMMG0wt+8PQZvj8jPWYnBwMvjd0y
SojJLGQktqavYir9vp3LtsTW1VDyZzX6z8X1SmCnIjtTpLLhZMzZt9evUC47
CBEXOQdMxcI1mi0OVVryr/rLyROnAelxYy3m5dEJhZjPjwAhKxxYhBnl8umt
bJ8SeNK9oOR9cS/fBsywdyHM4Bh5kulXH82uSzyzRp1SgbeKTH3ru5K+4K6L
vy0vImN1QV2x5QvB13i/8HpQdF40EcJxHXC2Wi6eJiBNLaIsmHTGzHCI8VD3
kP1z6SvJ4LjSgebXGYXdEYAw5JOA6/JvHVYHzFtJCSqDel4fVxRXcvK6ybg1
CJKa3flmMoJN3YoGPi+w/QeY1Y7jypy8sBgYJ+YnxzcFSoybk/OnwcFHZo9F
EpvcsVBGDgcEqh6O/BJdzIYLLSbM1stlZBCupnEBIMSsuQEgNXgz9z4MPdp2
fmFkm43tLy4YKCLph/QZyIxkc4zd8ZqbRWUoV7Nw8EddBq4Qd15aX5QbZRIB
MI+cfMC8fybvgLZekLi83dxoV97feS2XGyTAvU1+8Sua6w0LrDZ1uslhxt3/
Sqk21DFQyL+yf9bUltEBxowBnvgOYQ30o2+bsfU133CMH0MkG195/pRKElvC
bRyPa/kY1NVbmMT5tX9CpCqRFQ21BUTyZmrBow6cdA4c9BpHUnmk3Nw4lwOO
QyvW069HIo0lxYvhf9ZdQuhM0NpB2VByfoQJ65P0S6/a2KUs02Z5OvOvuIJh
v8+RIdbuvLHkbDa+Jb8HtPWOADDEg7iNDDBXqTyidtoiEqUeEjznp3GQXlAS
duJJCW4ORo95zrxxISyDVCdhp+YeFWuVuO9ZxLQu0ULASCOIFlxJzM1UdFow
HPkrop8GP9Iiaskgge/Brwlq7VTazkRvMERDKh7A6WtXi4V3ynXZEuU7urJa
AYO+AXp36p0omEvx3TZhRnbd5LhpmIc5/d5rlEHjlnDhMrYbh3zD3qmwRMPz
bM2gNEQL1IwjMbG6OOqqwHFygMoztPPI0K5HCgP9QABWNXlhHnjSFcjL41SV
1GN5rv6Pyc4EoLI/ip96RtooVl3qARD5YVw1oWagu5WWGkRwwrR0jd4pocgS
HCNCbx6FhuLwynpVSpNZ5Ri1SWrayWzQ7UWB88eOtG8HOhZMvDI8pvWxf5xC
GtQXYn2Rqq+na7+CP71ykV1DXbRwkh1QKh9Qgp48bO2R1khjYKby8pvgG9np
N1FwIS0ns0IBFrBs/iStfQDpUQy+zyHPq/XpkVLthMVMF6rx2IA5HQcPBXdc
8n95d36GwmqbdlKMLonndMNsEPKcHX0IY6Nt4S2na3+bMBQk5+y8IRGWelUq
HYoSF9sKKctzMf1m1F/BisrxpTOM7mb/n+Wk9j07vv1PXnvdrX7to+oT7Sj0
VPXnDM3CO9ndw/jawLueRTLLhqIQ+y1yVF+/Sulfdp9TZRjWMG/uCddr7yKo
DsQ6ocfDus89f9cwnPBz6w0anoKhzxaqXqVTjNSKLOAPLZ7H/rEsMj3+H0j3
d6a5UGCzoPWZ6XTLCSvhZtBqokjPduxHPgYLf2ofMbMnpP2bZDT9YK01kdSH
xy4aAyiM8nM++8tHGObR3xFhfRceEyYAznJGMdPBEeND+k5/k2F2Z/ky0thE
H5tQwmCWebPfKaltUooWGVzE3Er5Qcis5vdBPJtheR3Sg/Gq8rNZ/kDS3g37
FATHi3jLCRmO1EhyrrFF3LLuzyDOECpiYkAoDzfrKkXVkbxYtKVq6p0X7hnN
O63Ki4gg0D+AR05yd/gvCd8qvF0qPTyHpmjXHQPjqNITM4gUApF/5SjlDCJ7
aRYXyybOqbYcqhfKhV539niEWzDPHRjkP0xurlR88anyEPjwl+ZPKF5bmtEb
ujn8XMtBnJkRw3F4INKsYHNCaiKmb2HTeWfS8VH5gCyPYrEJkBU6lyq4uDoq
hlTh+BWRXHZtlta3sAkrY/dQaVcJHvn4wlBEIIU3iY3YTwPJU2m9YKQKLc76
3GSqIyFhwRdtUlta3r+RbLuKxp8WBRKllPviscWRvZbQUWYm6gJ+pi1+R1uJ
htSblSetiptN9lT3ZpEpkZTme8iA5aTWegbsiLmU7KqJVhAebWZ40WdxeNx2
8cHW1pGNlul2HYwvObh5srO+3eKkQxaNUoO7KkfXJwYaUbakWvRrXFZvT5HL
ukaP1wibPTLZ3Ls47jPY54F7vR0+2X3LNELfatfCcw/01CrssZV92VLlUv4Y
KWOTeFScRNk3g4Bj/BVdUtqYw6Qb+hKqFj4val8G1+yyxFk5e2iWtBjBjl2c
/w1VYVOA2vBVZ5coNHAtr6ZAbkd8AVsjWWPia9usiIRUN/0745XistjhWQB8
LSHyoWfWE2L30SVG+tc6qCzR4jxkvldFm1cmjI6xAOUMM+2pcNjTQTtHhrg+
E1BwUugJg6YM9wcorqg9WoH45nSXQ/w1bqmZ3uC0eUDix+f9aUrIRMuT2tyX
r1wocXyikNlnNjmPWKpxStQ1nYs4DztJhmhcCCie+xE/D7MSQsh3B3QFVb/f
eAx7gZpzHUcRzhzR61eqX4FTl7rLFqTSoshQvbp3cP/cOdZF5oNhvW5DLepU
trhkvxpOqKAHQVLJx/xct83rog3fhozZrJdMXNLsIabcKfPdqN6tMYmkB9Q6
dGrCBMn5ztGYVdwQXFfRmgr5+go7H1wT37i/+eTIdO3yfVRGWsRmaic6QeAV
bUGoR1j5/gb+BDFf5LlAMlRynknU4kvBUzHmLj9gGCk4uidtZAGUWlwGPTEO
u7PkcEcXlFmLLDH96BVExHt1TfZ27Ow3tc9aP0OsIH7SVUbdQZcpDsnOu/Si
8cTP/6QdWS4J3tbeMdPSTepFMvGfb6w2i05KprrrSEAhDkhxViEv6kejbr2t
nHu98rlgJJI5fHaYue0jk2x0XZyK8YzaGp0tDfJ80XTPgnFWZX9GQ3KQEfi+
ecedVo/726e/M8scvDAluDbT2Be5334tTa5MyKGGwd28yr1fuLylZyJ45GSb
S8hqmue5MttDenLDSgRyerVR9SEHao4n3OGnMO6seJYaSAgNHb2+mbSrLKL0
Vl+Ghvp0mvhAW3V9TviGFWpHafVHhKlPT5sjcCh1HQnG0DfpySeuVuFlDfyc
RAdukYk/Xz830HiRJ0OVk1+WOVhPWOrPjekc8aBUT7hppXvmyeM7L8nRa3l8
pntKtZ9lHAeiFej12V5se/bRgbUf26HS6LEYMsOV3+RppMCPuka0hA7ADBsF
w40deZz4nQ5g8RcZPwppTmB6QZUkW4gyslWpG04+PQ+3UO9EOkpnrNTjLmaG
j0xBqb1EFfL66Dfhn8Bbb3ICPCiXI/9RAnWTzByVU+bFBpAvwRTrot9CgYSh
DK4U2xQEwERcWdThGtqLsVcf3ui1p+Jtk7xtsywMCoNK4zmV/KbpjBvvoWJr
eCDFOuepUWT3nQ9xHEJuGa9slcNnFzdmVlRHxTZVcHiygDVFQZjKCfHnnJAM
hTSZUYzctOtwWqTDx96nrLU/GeEzR6FOvXMZVVJ1VCXTAHYkRfmlAT3VsCY1
ssAOfJyq6fphKbhCSFHRv199iXYYIzA9sDsBQ/qEj02jncLL7OvyaWU6PcSs
xaLfxwJ6Kx+jrdKNrLDw1by3n5AX9/+MiiRZVbl27KGEE0M2KMiO3K6y5yoZ
9A6J5aSXvUNwt3kBXyIMT7nOQhJtPjQV6q8Es09x3oyVJ51gSl3yMCfs6uqr
MwzCvMSU9n389z3kq0FTqw/mzOhvd+jMnGPEeG1PitLwYCXA3k+87D3Tpv9d
OzQkBzFjViz/pEcErMaKcijzPDuOHLVUpE4RHXrZdGzFGgw37mwZ8FgPH0vL
179ETQECMCBRIyvUBtiSYgRLyZCm6YBwqv4HRSka9mpzbLHlkcWTNWESNKoK
gSs+ioqTGRw1Z+3zCdO6CFcnsQMX++34zD2pIhNhEJnUooTGiAb9Q/gmJ/nH
LGVDpCn8CuUKD7HJn6BnXASe3V0KY4q6XyLRRhuphwIxRR+hi3gfjb0b3Y5i
F+cz6Th1sTOZJZ/+0ya3rdchy8ve1/OfFc3AKLkLGdXb4TdAbrtfRyXQGi+6
msUSy2w4vxMQNKtzMObq3ZejKkdmIxwh12JDoynYD19zIwMOPX295RLlbTsk
0V8lEyqhixTX/rUN1Yilu4DueOyKERAXsJMhhTTsC3Alr5xHdpBfGMJ+hOEW
xRojUt6miZQTABJx3XYwbFgBs0T5LcQ6HESfnnDhmmSb7OPlAUvNEtIyV6uv
yiVU9dEO24VqKI0gZIf2pfhTSGyTP2KzYSa9oQ06k/uohi5Z/zymCG9vaGeS
PVYDUBw9uTfXCZ8FXZ+YMXjCV8ShSWYPzugbVr0zLTELJswEF/dgzaL6WOaM
2KgKM7f3MKSTJ9xsKdAdbITQEnVyddxY6/LLxJ9lQufhvKMFlyRvP1g1EZ/o
fe6AxlBHs9RjCsYZz/zP8+g5lCestHXYzVg5zr7wVbLtD9v916iyrC3xtrem
FTcI3jMmMMacFpT0oMNEivMpGe7OR1BpREIHeyNNTXIpUR9nS7P6+5rjmx6K
m7fw9iyxk9JKU3vUKz0IkFNsT1peBl5Sxkcg87KucYFKDG0lE2a+9vf8pWdO
7kUJ/NqlUak+FEMQop15v9RDYWhh++tnQRVoJkBJ1XEjf0iCAwhsn0EG8zt3
4rQS33iAmuDbCxvp2MjJ9xqqQp5SLZEdJ3i2LgGISFfqtbkO7GCh1VFSDIKF
/nXpig+xp1l3VVZqaqBpIwQKuVG+n3s5gOm9MwQYVijlYQoDFp/VmnqlgV5S
8LoJAfI4vf+J45dtq6nUMs8EclwWrYY6aAYmw2x5kxI/WxrUTigRkAp85sLd
xwGzpjO1EhgnoOohIYhcXJ/PdC4SJUoWSklxoRhCevXhDoPsrLQECklIKnTZ
iN9i91kc4VMAMZFHjfryJlxvwHI7HSKdrsCU0ZJ3yRshgcqQqwMSVAbvzDSx
HnhOdsbdZZX6wJ+1hIryGaINoIh6IhCHwhj6VcBjCTYUXk4lXJp+Op1I7A22
3BFPN9/QbySbUdpqrdv2KiQZ0h/r4Uo1reec00ENcTOpVrr08EXvyoI4CPYB
rYRhuKNkKYgI7BpMjjrzoKNLieLPLRJqyEuCFHI1ev33Kelq9yt6bo5dcEGt
jf4ppzRjVjKzfT4gg5upNFPf4o1e8kZxxULJPU7ZGSYj2AV1RA7Li0XW0Orr
AshaVl2LaxK5IHyFTzN8w4C7VC+BDMU3G4opfZ53gdYCJRiJGe9/5DFLvcfh
bw23ApBTDl2NwzbW+papasud4xWoVaBUW4Wh+70H2GF0y7IingyyOwVK2iEe
ivzH4ofbb7eWJRTc4HAPHH8lbw+XCtt2dAb4UtJpaI0W6ZbuOxDZWWEeLLul
msQCTSKhzyWosf4DEhhALJkABo44Qlccum9bZc00uo1FFmpRf5UqU7dgj2Dq
oggmVBmvuc9aSI/ytDi9S9jkcNhzC2RuQaZpECruB0FXhhJi2/SFGRWjXcUp
6+lBfXIDxphPNPque/t95prp3YYLleadnvI7l76pDs4UG+W7u0YVR5aAoWLN
Rk+9pxJguDsEkz8lTMnEm4jbfqic0/TJBRcl1vHgI2Xa9xyiL3Goy/OeqEpz
UTU4o9YLbqCEuwewBnsfCWB7QGwVNpO60+OsrYxrGGkzRXK9w+eqNd0U3HCO
044dzopSXiaNviWvwsUoommLflujTe8RnQFbP1xt6l29IaATed4ScC0THWhq
LVKApb5rd6Lr+UGsURJ9DWH/oEvdkTS46yF52+rQfIN0Nmp3nV6Y1juyNDi2
8SiFZ7BfYYISSKryaafwP0L4LI0hm4Uz1GtGAO6f+VM8zS8vrG+T4s/f68cM
knOiHm6hV+fVxcSyO3ItTb1sGKk1gJGTVsB53EOhLFSV9LQdSlhqdustbId1
F5IBOBIySrz8d+mCC1lMYRzEZq8t/WGL+mSnd6nT2sT+r2xsw+KHHyeR7XWh
T0H+FXhHkIMjcgWCafjlq5C8MF5VeO6ClxAmEXqDwT7/ns6OivMeOWqhH541
0F3dyvDntClq9tyEfblF9c+hkgGNaNQ8EM2HJQDA3fajfZwIey701FZeigAp
Vqw0I92iJYjAvu/SMGMqZpY1PyJT8BhR1vZsKU/yRK3cNKvxJ6cBt2vZuL3U
libhylDM3M3Sv0dBxtbS+sLiivZW2KEju5jvo3JBoIC3FrqycWpBcPECtmCi
1LkCHo61jP7XtuHPuI3yY9YcycvwR6/QdX56exzSMMo2yCUWFmGKX+YHKGWM
oHi7+Tu61+5Q+HXTn2EAmxne1GuVlPxL0SyGQlbuLilrk8A89YcLox7c2HoW
YYNLGSjj036Pjd5gd9MA3kUwLo2Uyd53LaKHnWbkCtlbeJdhLEFzwrmFyrJ/
e6CDJ03WVl3QsjnVGi5fDPFxV6tv6mfZ1bQ6inpPaKIbonYOxhXoxJQWge1L
s3fA4D8RzB+RZYGEm1WYO1W53en16t70tpLJbpcUVa7hezwTYfqZIHW8aQm/
mW6VP8R/sn0/urBIg0mmguBh7RQ9DJqs0X7enPcJeODk9z78bBjNmVFnHFUe
GV4n1YI6pBaiL08SCO3zppQemprIWzqSFNegVxJ6wbR1OwzG4VE3pA7xcHJ4
j/XpS+okgUgwzNgaKw+WD8v8obALnP2U818N3EHj3QQIOaxCTs2rpU3O1/On
Hu6/7rZGQQIJ/DTP3NP6XHNxE/rkjaWZZNkwAErixHE0VYBVAA207tmxyD+8
dkB/XZJS0LOkhrGFABzYsKAqYMf6HcuKuDjQs7HcMYnfcmgHT/mxDx+8t54p
RS4UyTnJUnOsup+BQvbHefIDQ/Ttm4t8lJupDeZris0wX4QFpijGCHpKMItm
3vsqp6igz8JiIqgS+Xd9Lg6YZqqQHN1MmW0dLQVpAcXbc89760NwYWw2TPMy
cr/tL8AAfYlFvyvWu9KFSIAJEgK80CRTlj+molZcFtd2j2B6ID9BDtkNGkRR
vAHu47nFOGb5tAaANwQ99Jod/m5qPO7+ExA8gl5OnBUxuT4ngppZ1389x/00
tx4EZxgfQimFKknfqp52KziX9RmtXTiZR/w1bckwHv78EsqNDDJvVgn/6rjL
GVdUVWEcn0ho20oPl0myhTQ0rHEjbMGH53+aZvIkwoRF9Og82YnYGh3611/N
Uf6bfNko3+FyF7AlcNJhRDiMwBp1GkePHUQ7KXYkPC/MHoaSaoaPfbAy3yam
hszE9L/gSqFtSI56tTXBwF16o/4v8Wm6dYyh5xj1skG+Cvs4rwdkQfJkinK/
pB341Um0mSK8Xw8FJ274G2F4/M7V4kVr9yt9/KDn0Rw3zMZWi90rMF1o6qlJ
3cn9Vy0cSSJHBjghZfhITdPxtn2Ar7U6OsDyWvmbXiSJWAoYPTuWLOCZuHbi
uxhH72FLeKFmbCMd9lkawhnMNtxg2NaEC7YDyq1mKFNQzb3x+HpklOS4b+xc
SH72IpGqF2DlYozmxf06MgYnz56ITNyuchAOzXj1l3RcjPgu5Qk3+xQBl8IV
daZyji5FLbi/vmBbL8W9b5VYIvSG+UExzTJhHt5YBh/jNe4N+YK9EcswlPo5
XdB4xUqqAdFXq1qIPR7PsX9RmvdOezgQ60G2zR+Iee6APbaM0tWcZ1fc98qq
ezEQ4BNwDx6bneYsI1nvPSle6eTDoDuMqg2XlP8CaCGCFQP6c8Y3x/+SgbpN
Gg8peLZrd2eKJFkJB1DJ6zudukEnha+RaJJisPhV6Nn91q01P0CQ1btcxlNf
yfqqbLTDAjLIHIrsu6vUQaZGtqRybs6lTulqtPJt9816rm82AbQHW8YtRdDN
+J3cZpuc0EpQ7tpoYcCiHbNXlcTZmmCmk64HPy7ifn1kBQAc044Ma1NdMk7l
30zQlZeCLsM6iaH8S7RNJnehFokfTFDsf9BYvItWvoq3NNzAbdxpm4rmWxFV
w+TyiAYSzlBabBLzxnDApJIAfPJter4NpB1JHJVO/TegW8jnQQ2SHDmjo0gj
qXi319JefVAGzIXsD0Yvixi9nzN6aH1q05van4zlmbSM4R9sX4H7qCFDe0k9
VQ0gcaHgG5iFNEm/JZ334LR519WrOIXy/iWKn7N5kTnmmTGSBSQbwKwxr7TQ
IKUM+TqscezkEbfp/rVRqgWxYYGGx43f41Cv51b3DV5e4qGrZLymhJoIi2Xy
e+9ALFUmomJ+TA9Zf+LMAxb/JLGM3f9E0SMAmEQHathrNRPBs3JqAOYQW5B1
Em/KH5VtUoaiX96/+MjsEzFmp0p+X0/yS+YbEwDxAfSfyZFmMhZmA/dj7N0Q
g2ph3gRfMwpJFX/TF9BmWjiJBmg16EZdCScK2Amelosfr9ZT5OA4mHINMsqK
XIflkjmeTN1ynEWa5KCqJJPCZYTYlbBRxpEJSFWoOzoVrjkk1BhBjb0rd7fz
aP3ajbKTcDQTy68kxVlKFIrM8KVLjckMHzBusGJ59fn2lbW+RxSdd3EeqO/P
lzaQ0An/d29/GbFnPGrQzji0nn8TyjSHe6v33GBRQNaSDIUJpxBvGCqnpxuz
RuGJ5KawkMwl9KSqfLRUVh5jEz4jvYfvB/3zjBa8MqsCEv+HIP6NoqF4jckf
CZEX96CvApObeB1x16iKxEhcAYzXux3QFl6L80DYm77Vz55izQvfwHOH/Kp1
vOJfg6OEVj1ODgqmdhM7wFgqGpEx2Sw7d9gkMAvf+T08vE6s0P5h4pZ8dL2U
ruWCDUqWP3ck2L/iXJTvYdfVcyCgANcM+uaD5uvPOCM/DMz/bHEtN/XEaY2p
lr57r6DD1tID/GgEcpS+duwMrzmkUszwbEw4jr5pU2Se9QHZklsyCfqFfTHk
hT8LCbjgIrlYDSELocutJYfrwQqpThNSsy6krgDEXGV4bTDRtoyO04Eqw2B3
k1sfPp9Tgix0Ccf6iTJqwCH+GvsgG0BBO1blNr5SVw1eukLh1uwnq6Ud4Sju
wAzySd4vqmuNavyQQfz1NfLdJjkT4Ly98TibY0nZwe1Tsf5QSu0TBKVGVFT5
JxCOFhS0Rh0nbxkZyQCKUFAxzSgRL73PL+lzn4IdYHwzRhKA0hRzTTnZLQ3W
zNVaDIQNNb/OxHmLMHHwPUXEYlGGBI7ErJ+QlP2f5o0SGgiOjh4x78R54VfR
PWdrgutHWdVddpDmZ3hHNE4k489RQQ/SSTcOD9UbutCkBqbRI/blElEaYRT9
R18FPRnruRl7lzllcl+vVsFWS0BvbxAcONSea31Q4BQewcAB7YaLFKZN0XzE
NrRsb7J0bXHdejkgW/bp7kzTAdcwt9r3EYUSU10KAZJOEdYApIK2u+3e4f76
sbmlRvnKOJBICux5fzC6SCN7aHONfm1OHcp36ozWhXv08PejdSzkDj/C48EA
gQM6D6ClsrclvKA+hZg4Juc05k/0uQ28gHytn6JK+5kaP2ZVXKDMJQKcbin4
RPxPopiGS0KLV6Yu2dLLyPZk1LaMiNOIffbSoyyoea7gH23OsOHEaKbESe2l
f6p6wlun863LhOzTGO9qBXv0GZOLExmE68lJEm0sQFZdtDgHv1iowrtTHLNF
JNd8lEyJhokj/Q0fFwDAXx0oF3Q49Em0T5rgzDI8JbC2X5/zCFFAZljTIybq
Ixpnsg+t04U1be080jBUWEQGRUonyVPEMJmHgHPcFyqPLGzjNGs3aJlFmPQh
ekRZtyFyaw15ZG3irIfR7a+K1ea8Qt+vgWvYkXggf5dd6IKwVFUDnyoZ6kho
Mq9MMiEyZ7+b26Qp4KDwH/EmY7oPIvzRR8G+G4vaanaWCvXmkLxRkYJ6Gcbl
UaXVCyAjIp16utOL/PkLX7AI2j1LC13OAPLdGbdJjKnHLcjEQyo5EfcBlMR/
BrZGMw5XmToZmxtimE1JaW7HY7mSegmgMIsp0zhRIxEKDWCmSoWtnS8CB5vd
YNy33S+IQ8jer302IkEFokx4YgG5POtcQBW72YGWtBl5jJttFKh2iC33Hfk1
J15GWoLbQYtR9xC+wmnD4l5tFg+o8aVwovDBalt9R/VJ12M7fw5OpFjgDa5j
Shr3pss5VhX792ZyhaHCYC0c9tZ3yAmaBtryxI9Ue7r9TusR/JW3Z3mYTu69
/w9gE1rz6zB35OU7mYZ2gNUXnHNtSDz1YgxZt9ZsrmLo1kynajPodXObq0qI
QXd0wJFoGhD8PJK9JZC3CMkLYCFV1lHiKuXe9MqpZJAUa2dKvW/cl1dJDUGP
T3spz3jlTJP/+OcZ05rF/ms/HhmogeEIw532qETwlu7TJmO/fQvWm//jDPQ2
ZGSwM2K9B1WHGgVUYvIuGNuWIKpaxVbkha9tKd39AS74+NTzAkyrEk7QuZEP
RIaSYl3fhscLktZDJiOfTgjvhiWFQTJc7brM2cFs2/okj46E5nVieskqMA3n
jDWOb9mRqsvrz0NOIC0cmPc3j/LKC/AkV/nkAZxGgxW/joN6d5Pi8NakomRg
VEGTfnr3VXXuPdaowSICdkvGIyza50riFxgc08hX+q49f1YOiFcuo2OZLV9Y
NYHSvHDkEc5Q5e+UPhiZeVYOJDTJlIKSuNOoC6b4OFL/E9Ub+O7heBQMJc1v
ylXUYuP/sMaP16AQyDjPD0/kyXoc9ivj0YH/KHjsrxMQUKbfwMQD16WYOYwZ
NQqTGTktG65GwokqkfJ7N7EnVO6CBe0ELr6S6Dam6V3/Byzh0wiHIiBLNKCQ
TsgXoPHLGoUglIQitb8WiaPjMk+xi2S3eG3n+pQ+93zJBUtDnMcb1dhwRobt
XQ6P8pwOCKx1g2DHWwaAOWLUUR5ithWD2p9+r+2Ii7D4e9Y9necAsvg1pc+S
vPzN3vVLSDP7f5jC2qys60t+NGXQ0N7rfMo2OFq47wI046V04B39ACw5BDru
xMY31w+iN01e+Pp8kIU0eT4XOIBdTkJYpr83kyHEwC73C0OIzVfTxXejYJ7W
9pRkE1u6XIXc3n4hntoNIuOC5Jo14az/Rm4UKIHmosQ5bvMv+lPsEhVv4zY4
pMTcwl1rzYNvS8EBH4sDrotLAJOWCxgVLoLyCaaxrLQhCBs+eY91cJVPcY9G
SuWB7wSd0+vMAml7X5pAM/RUtFVZ1G/t6I1YI2OY53D397xiqP0SqMHqEstC
FmzWIfZAB0CKL18Zzj3Pqp34met/kXQ9y50I2HRtetWx31qfKtTCv6LgcG/q
DUzoeNg35/Z3wMjRylzOiabB+DE+kweANo4g3ofWkEwqtfcB5GthJGj3CX4p
p7iF9nGY6gF2kJy5zTzkbO0ATPEefLn4gUswzXEx1H9UviLKnCUVk+vPeJAH
MyLgU26eokhJrEfdNqtu+MiOup3fZNVoRW/QUEnZHMmSx76isR05j+c3CspP
NsDK/S73rBn5Ty1Fb2FlTlws25CsEzl3uVeMMBwAQDKnknqeaI2+jQOz7CI7
JGxxd+mwk6E7rFA5b1GA2atVC4P2UGnE6GD1iKmP18fgXa0tDIVDnpYKj6Iz
Uw2D3hgMsiD2ZzbigHbaA+gwW5zD7CPmIzLRBbNFu9MqYrsC8lT46tnNj1jq
B/PNymKj0BwUuxlbev9d0OWe9uoMHj+eWZLyyBJKQQ+RoyvZvWp2N7gPERCJ
iekEFt02JbV6Rf49doEM+07iDc1w5QdKOn0CEOFUYfvZr6xr8alBg4CNwgmF
y8zaXCc5sjQiOPIvCIJpbUByZIT3H7yNczxD+Oub84+mr+HQ6QH2KP5cy2Zt
jY4feQS2yYHIOb5vo7zB03eOtWEYG2ELHRk+8w6zBa2rJOIrAWcLmKqEMusB
+ExdDAGRmSlVL1Y5zE4gJOYEtAlqbbTp+aRaOhCBSFXcTzru7flCvZ+clIIW
b/CWvJpMGJqjvDL7sldE5Q/M/qvyq4DWPKzej2zfWaf5/0uVOM7NI0s0l486
pFwf7hEHKZU0XvBeb0wFqCmAxed28+0tpPOW+ek90UZqFYS08mYyOAA1OR4w
maXaIRNxXmRIZ7GJGBbw8GQhd3YfDjUE/PigcdgWuQQb91InSFNiUP7MEefH
3yI7Dappbp1IajaS/BZZGpCFlf62yhjiADDhq00DURT5wH/1tXuvVAIr58BK
CONrsw8fwAmEqwZ32yCJ6DK84MP32L91Mdgt26zr5VCyZ3tEmncNWK/dmTU8
aNB/vPcSsFadEOjJscR9Ja3mrK/robA+IzB38stBP1yfEHCNXybr9H6NCaR+
OWeMhpwhMQ7koo1jpxq8rbXIUec8XgJI93ceFXPNEw/36Z8tn4+TZraIoMyh
+wbyDSawCDmFMvkW+LdqUlu1GRARXy1U4523iAMI18IUdWumWF6a05l+Z5l9
t0bSpcVROtioip0nUjzpPoxg6v9BiKZHPNWEyJ60bWEH4XJbKfhV+GQwy7DD
6ZiT47PK0qcCs9fgBNHTbbzOI48mGvus8zHxGXJpqajM5XaIhDfrhxpvKOw4
g8ABGibG/mZq5i0C5IzKWfSA4PJiT6rSAP4jTrLf09W9EEcuP0nsCAXGz5YD
+CTW8wDUfmSaucN82zmR99hz1qbotdKQoAJ8aGBFqddFCr2hE+G8J9cFV75t
ZYbGEfd5obYv4gu9IWVoQBiA032d+p2pJioj6gnLwuFX9boZB6C80qrT+xzd
hQfJRNAIXJPPDHN6SKNNreEOR2z54wMGWu8OoFJFXIEFi5Ue3wB+Nligzd1O
BqapCnDIjeVuybRm0GVmahebYn85MLmJIQuTD8HM+r3f/5JXK5sLB6KZ+aOJ
kfMnyxOd8UtKm6OAwLJklthtqd6N+FI9uaYRe1m9ZmbGLpieFibbGWILlO8D
04gvz6M6ZMbBiU7BOqj3QIJt6JOAUz/twY688twiT5q1UB/YXPBOjGTejqE6
G6vyAvun4CMRDTBLhT2nBOyoRsE2CxZdBrAramy19PsFaLiBw8ser4GI8/F9
LPMGeZp5C1FmdITBeBIKEvTOGS78WQlUlbRnusno6huByGy7lfZ+CBk2m+6a
v1OkKZO/OaSGQOBOMpv4WL/zVSMNMoFfLb2GZ/NXGbWePGfBGk5BNi4xp0s2
EeJ0/Q95XwGkz086LuYQm3l9sohqOR2+HKRJUO3MBEtMhSwVpNeT1B301LWf
Suh8AM1wcMPghGOCDS09hp2vSXeSkZGC3LDBBWzXBPzEa2dfHO0OETYyQD+A
BycV+e6r65Pn3P9aR/p8FXPzybi1yIm6Q2B2sOByhtMsfLaGG0ZMFiNo/YYc
xAmnZjs6tW3+H0QSHQp6eIArHbvZ4uNU0mpNDKV5hcKFDc5gEUgTDxI6VHFQ
quxlph5NY5WICKox1SQ8Ipx8IancLaix/5qoE2leGH2iePUYN0BZ5is39nYc
v4YuuwXp7UkezcQgF6/q4frK1G34fjuEDAmRiK/iJ9CKLTAKYLosqlbHaYq0
Bfe+Gdy6fUOneYbD19PGtFVFd6vGV1gtIXpXDx4qJTGYr6PMw9bnvozfiEDz
QC7xfPvJu9MOTWR+iMyUPMlBi93vej7+wVhCIoO8A57mBSnQYpeMLp4ZBOrH
JuS2l5RIqxz89J+KECY/vU78BdR6AWnfYltwxe9I25HYqQ0ItZZzFpXHuDu6
yeTHiUzsfIjcgOL7taZ8eDaBXUPaVWCq5bLS0cCcPqYRQBkirtxIOV8BCM7i
6KF0ZEsPv9h8y57tMvJdjINVMueWKbtvxFuz8RC54J4BFZCBPaTwdCkfXS13
/J2Y28BDDsBsyIWRATGONK0Xy7BqWJLgGXbEMpuKRzTeO8QIrttWeXtlMLi2
V3cvOFEbayeWYoZ0zidumrPyzy8OadEOlPIvegc2Cgih73gPsw7bxHH4eBm3
t01fBl401E6J2PrASDmpnRlTS9USRvbRDlVoNTq1HAyAnjKXFW0K3trfyM9z
2SGJETmy2SrLDZhPxLTMT/hXOJfaxMFrcoeRPrEnZMFkxmBEoP9trhCxDDEe
GJvxpf6eCDvIwxHBu0GYpZVAzDI21R1o3L/FCeHLFrxzyr50NI4SctepfTrj
JAocLn/J9NBZMUaufhbWM649roch/88pYyzpYllCkO8ZENKoThgSC/nhyZ1D
fcsj6XLypC64rtoNF2v913CL7WRqmyB7clIgzNp1gGwqFegdjgQJHPdPEPfr
s2PGtjjngIiCvglN3oT3gLxVGnLMEeJbwj2g7r0noEV6igUUVL5imz7jprgl
cYvasKW2X6qBFICo/TH9N9ly3V1R4nciSYB+m2erA4/Fmfwz+lMXe5JXj1RG
bjGvCSSatctIsNCBGc7jPV+cfIHcz7burnvad9PqVvK/WZ6kRQMgpUNDZNbr
eLLrGMqtgsRLGeeD3S2oxZK+dYdfy6RBYTnFPMyOLkG0xpqQwPt74GPMFRTE
/LQnY2CvZLhv+7TwymVbMJA4dCPEFP26gYya9hWjdBjXEREZ5IqlN9TDyRS3
qmqfC/9vNr1XHJ73Ww9ECFsW1JZa/E1T4t3S592JpR02Uc274I9W1VUN0S+/
q7sCO2XIh01PvW1mN929bHnGe5WCSo5lU1LjDWq7RTC7xVLiypPQyeWigCmn
nSeTSVlyww2WVEP0ksDhOu6G2Vj2xoJuVr9x1aB88w6KzOLMPiJ8rlv8Q/HJ
m95akpuj7QhLGXGgLtuKLCRYqbM9cVMEXNikpb432sAStpkyPFqr1NA/NsrJ
lOXhguU2Qbu9XPPELwFiwr1sM8+c1UVYcCDmT9fI4UGiURdWRfDlXr8QEBRt
KqSWEjJWqpHSroc5HeJhsVItUOIOeU1QRK1diGsS+6TMDObdn4cDx90JleyJ
5B8ofP4CtTVSLhkFSiF87UoDHXTx62039bsriX60nzMB3px7q2So9e33S9zF
5ifOI5JVEC0jpYM6KJr80OgDIt9EuHdNkDrc8eaFJIZjOrx7RlAii1ZPtW2W
cGQzBTss3KiajpopNEa5r06VGFL+F/XwtSfRE9OsXavSpJ02fY+3PACLw96Q
t2HQ/FayYUdpXA3KjTfVxgIGhtNzTzUdP7ugQRjMzHHntKDH7GM9RhbnMaZL
9O4wpTnBSfshDYwWPrjMqinTcqXvVaclWDfMs/ErhvCjOdsej857ES2XLFa5
jXZ9JkQHkcUmd9A6vURhF+KzA+f8vsRfvhhfQ5Xu38L6/tHHeqerSfA4hhJW
6q4EDv52MyYOWWIbHjwv8z3Uq9lFqrkAgZur4WgrwNi+0rHA2NafyHFEWmds
c7xJewsMzsWjb8PGTUXX7xRw6eYBZjJupB++RPKaeYtE6u3MNnvRj7KRt01L
CpXQl4r4HiCJDjODnrl5c7DaFq2KmkiETzOU+/LTZFPGJqBMkkt0XLlJXuO1
L9Hc69dfCLdN9zB+gkYXZMOUVtKHU8ASR6kCEisuJjBVbzMKitjCiWgWZKD7
K/IdBpffxEJdABeqYFPy0wWdMwoPG/icqNzUrSo0wg/FtJEYBmMTJ7WJw6bC
l1sE1XkIFh65R0JnU1TDU+j0YFawLUlmVtPcgh7AejdA0tgXbHjod1f00dL2
nK5tgbK6z19cxoXpWTc+PoKgJlSibQqCjRgvcuXgwz12NAnqBZyzvpXEd0vl
D+FkSvLQ3MXJK3HpOT34+bIMxwUJtv1bqc4svN/44qYgXEdWEWnytkx6whOE
J23NFfZl7xF3f1yYGKwEeRAdiGhiGsq6hQpAstXc/YtiIKqYxqlqBKTUFLwi
j7M/qAPvO8RCNrwn7wxkCxfgIni6heQD1C7xegLVJTV+LuKxJdZatd5uA+q3
Cc4y0WX5BMVJRzUf5kAWFt0UB8u3NfQZT1dgR2nObvU+fOWzbG2VIcf+n8qv
2Z1qxViJogpDqw6HXLUFSB1c9zp/w3/hsBOFh/nBsaWsUo6yHNjgaN/XLZNp
ITx2RnYd5LUh+J1sq8MOVBedgia0spghY7DgCO2Zgn8gqQZrMixsEDHIC6/v
3W/GhOhvXXk+BLvl3tt39/dooZiAzETYktvcgSdTRnCSuBX6i37xl0tcAqIb
sT95PqkxKNcfXwxhwYi6/Sg/lN3Fe987JRREyiIvTBsZ6Oobp+mADVBXE/eY
Ri+jtj9CQbgyrpBXZwiERp2TkdegC74ciiZzimTish7gurzfam9xwAL8BMBZ
UgXiK63lRkTQdmLf9ETwx5bhUjAxiRqbtkF47CagN2/hiGdyay0iGWgV8TqE
bnn1Xxa0LYgBxM4+AtbipAnxDjCLxePnryFk8yjADDHQXFBLqumILt/oSg0S
CF2hfZeP44nypn+uxjGrh3QI7/xr9AfxcEAmj3P/oD7FDRPdETM7BNtabzg0
IgvdnD0rm8B8T5l58eCLEx5xapdZemWk7k3u+yhNmCG5Egq5bLc9PzQCCUY6
/drMLLhfR82/dOy94tGy810ikvtewiaTsLWUwnr20NGmk0l0hU15cFdUmkh5
ezmSylwxtAj3rhD8PlzpbOZ8H/riHX+El4jFmDwoYOK6N9BSRCfPEmHfJQnv
JU+ACo0UMiL4+V4kQ4qIqbsrKuEGT3uN9a2x0rie68cbppfPYtB6e6QQXthz
6GyM8UfoVcXEyLHkyQ5vl/p5wVLCHhwqdoHmsUTryDBmRODtH2c48e16NK4F
web5lk3VZT7aEn8c4YxMnDTSghcfHHFZWSLaRm87u0UK1ErXpYLLZ3dmJRsM
btAecl67wWcLM4eVjdbDiTkK+iIVN14HwZkAzXitgQ736/rWUFydlFQH6qcb
7vnA6B/HidIKB+uIoauOQxim0WnLHF0lO9M50/eVDwXOtiMBB7VBcpqY2zPV
hJj/CJ+NZ4zFq9NYZoEWczXorrGdDAP0Lr08ZYVKzWpEPM7k1LhjEWl6OVTX
yIC/0CNTZFpf5Ut/dvxobm/q3++Te9cGl5kyO1gEUgqojEyOeo3+8lDHjxVT
KoZIQthxPn7+oyB/nVFUhnZFmDdYabkohsp3zYtGMAvnecMyS1A2DoFIB5hU
wNFtjgT4J+uwkoBSh01rKVLd2NOMWNGY2bIVGKtkA7y4eOSkPheJCGJaN6h/
jZCz2rV9X/9Z6hsJJWkRNGAVjG9ncqAIPRXUsXhSiXy6QLMej9A7aXgY2OB1
hDgWhkW8pBiEm/PAXijMkpUHbcw4PUsnhde5GbTXljvhLs8jLDz5E0puOFUf
PEuC4IWBnQAFO4TgBshE+keb+4NtAk9RZqr7GgbX4JpJ0jc1Tnpz4ynpvkR1
KG4PJLdEl4pmlyycsD3Sya9wD1mFTBZzF4PxwI9y7EEVhQpmqZ668PN7MOqC
8v8cZnt8kamLtSKToWe5XlgbNArT0/tHyQH7Ua+mvVOe1/m+lWd/odaluzfl
VcEun7DYPZxnhxGdVQ9IGqCqQ1bV37Uq92fahz3vLmX2i0XuuAZC7rms9I0d
NzZqsMn/FEaqlS7bhqdG4wy7PoBcovVL2UeHIRwq44R8KXA1udVXW/DEHnTR
fhECmx/LMSXpjFp/bUSYEzsRtYo6wbJMqV7qsvnA9CKx//szNkW9A4bCF8DI
ZlN0zmv+iR+6fG1Jgw8E7TyB1YneYn1vk9owONcVTQuWQEl8p5xNSsntiR5s
K5R+rmi0rNmw2fpyJmhRLfQJBXFZXOVxAiysPoPbRRI2B23B3kMQIkTk5B1R
tnBB49mmKCYerqFfGBQjcVAFj4ShW51q9U7jY3oxJp/kBq2dv5zqmfZDOd10
aeha3Zam7sY5bUdTQvsYjHmG7g+tq9zIUSpcmXufSS8h7LVPveYhS1evdplj
kGQywyB5svHXa830WNt8Pef3bsBCzlb9twqPm/A3EMwYpE6V9s/mZ63dieef
J6AMcd9xmgyzRg6fR3mfhu/YQoU7UDCLvWToQWlNL9ne3m9Y438zM+4almKq
oLdBE/4NE5SiWNqnNh7c3aSTk3+FR2w6xWzv+yrcwZugnaB3rHqFOTRKqPHy
EEcW5Im/4Mh4TuyMF1hPoWo4Lmvv/uR4Tm4D0beIaJ7iW6dQPiGJOYBASXTj
vex66rsZS5m00o2lkGmZEuw29alfVSLtK/nJSB9ricwkqvG/7Adu2FueokJa
eqaJaj/zRa0d44C4NY1ZnolvkYAqk2wufLEU17MaIP98UHuuoceEWGVf/Jr7
bAtH5WIxYoRUOEaERrDPeAr8/hIujUBYXE7TRANemZfVGjqohu/TrsE/YOBU
I4nOSsgh8Xw7oG3RjAdn6Tkpvwj5APtRyPihszMkhelQDnHqf/+p6UnF3Xj2
scPqOI2ni/4rJ6JtNq4I7bqg+2FLXzIA0abJE6eKLaN+zsd/ggaPn2M40xVC
CzRMoAaFT55VNtUPFRb5g2z6r8VJ9igyU2TkyI6yBdyQuGxiOv5EpukghrNh
Tjs9mXUIZd+lmbxS3aHvShvR8mgy+v+AHTkTZbmrqhFj+hL9QmwhVaJ/rF0z
rixIp6pxT/m4xHh6m+HH/ILQIgFMIlNr1A6lS3wzJaq+QPQP80+1HDJM0tXr
DfL4tiXQCCNADLBK59awERRtSNx+xkkRn7EaQzXABP83GHWmQ+1EdFkP2p36
Fszr7q42Nwg/XTiVYzlLkDrnqpzKiUqg104zNbRFQ9O4TGpRDz7kuTrwcnKT
ezHzwrRRI0GpGE5vyOonGyb6NUOvVrqavFnjN9U9saueySxOarF+mBuJcIlo
Pkij52SDqdAETprz7u5B5ZywGd9VfI5+B7SYiKTZfVNPbcc7GmtenYl5XdHF
ve0VUXt7e5JA5whzL/F9xOM3HmhUu/b8m8sAUDuBCGwtbA+EeNMtTm8U6/zZ
n0Ir5QMtHdutWoVzCumtSNulAceQYQLouGIAcx4OdxqGXr2MTASI1A/kPkeJ
s0FjJmIlFwqhjS5+co1Iq3QPwo36eShd+csUlGAxEltUUSrerFgpNz5Qjhs4
JpZ70SJTXgbUzU1WObqAaH2DekVQ7TQxSsV1v7gm9zFjBH1NmiePs6YHjzK/
4eEJT32zbfNY+QmeFwefd0NIix095zUPF+S1fNRZlZI7XK7WxsXvMbgfZokA
Q07OnNJVk+ykt1m8t050tGJgYzQLrrBzM2t4WSsorjgTXP5aaNR61XZuK3XR
sJuJjn9w9EvERRAk3kcvuHbrwDRr0K3vf7yMUmWx+Q+ekhFvNZ88A83eHeb6
aFibSby5uU8okbpHdBhBYi7f+/UXLsgcTw+jcyTFhYrMNY9EBTZfh/prmgLn
it9Sk6yjD/WhBACunA4TS+3RoTGx0z9+ARB+ObQ+Rwb7wiuNwmoahIqvhYvC
hUJYVzyW8zw4fKO9Diy09kNxx8il4XWRi82osmetxd72l32tMZSQhnMDQARs
BUHzETkHxObDI2bFrXfjPcRKgk1lj/HZ9BfX28Y4pnI8K9yOCUo69eVdSv2A
1ztoYWJh0s1zbYEFe4Pmzj/jlsp09noWh5efygSh/EhO6ygpmgyHJid5AKMu
/nD3rJCyyHui79bzFoTbR015yrYtxdy+dG+b9HzwREsOYDabNilCwGo9fmSv
ZcczYIynCBJhd++P3b3SfvAQATvkCP3xzUtlRlT4W4Ip5LOwnLcU+NrVUGDC
dD2Fu9bmFZ4igWpcd2cfnTlgf13DwamYaVOMYJHbAb4U8SWrV/an23Qeif3z
SSMnaEmqYGClYF39jNrErxo2qxpN4g7pOC9PD8g9Ee3S7vQHPPWnHZ74SnCR
pou+D4zGzrb9HDvVf2Tz0KgM8bDY6yE5FQZO5uV4DnkSu/iYBjFHZYJScLO7
4H7UGRwLnL6Ucn/x1O239eE1yUfW13+IeUIYMgz0F9gqPP99NLvKrZbr4mI1
rV2OkiGjWmFSfFmXlvY2cT/TGoesp6AG+ee6VAjZObkXXzcRDfwL/HQnxkYn
rgDTbybjjopIt3PFdtOFNMOVk/yBdDNBIj03WrcPSJ2KRBuAafvhxrL/T/CW
3giy+KsdX3liPP5Nlbx+HFYgguS+goNW48P2DyLQfOHyBT7gmYZr2+OuiHWk
wmBQ9ltvqxV7aFhbXUx/sNCgOgj0IffqiIYlH5bOPwRHvmG1o4nspBOXcPJJ
tbIgBI6C7Y3Gyep3eZoX085wY2ULdNUxEh40m0Zx7IqgGcSsP/nHgXZ2sSmU
2mX43vphI9PQRupRZK7LNY+XzcH/kSQiWtuaKTqIchhRdzSkaPW46yoL0amt
lIsr1dQewupHlr4YoeAY3R3Or2X1qcsnECsktz0Ey/lB9hoPrtboBqgpYdLv
2IrsWBT3nCAYcxyl++rMEzrK633KZQUizY0n7rSdnK28xiAPQVGsRttH3Fe3
AlhWZ4Nqmp+wWCorJ/Fpx3f/bSQqqT5IvHo0sdryOQRhZH55JQlTinBApa0R
c2rzgkvUcUyR6gVhIlEoa0IYIZqS4Ck7R+J2Q0BjCNcFVP15Ad8MOFMuzvI4
e4tlgT5mES5dAcoulUmsUnK8ggxXtTFhBeDFe1cZQq+zX4O94nr8r+LNJ6Ss
Mjzqb9WxbTYbzwB7nghFHBOTZdwMf8oGGvgvG3to0EQqLJPtTEbY6ZuaduKX
SzJb8Z2BHES2urylD0O84SGsRqTrNAeGrgnrZaNgiuJwX0lgSkJOlOne1qXd
Mh8LH6XKR5XIdyufXGltHzCeidSBmmtTuf8K6yz4p00baJzLT6j3QCTdtMd5
9GQox/f3g007obxZ+8QE20bHgrSIdhQwnCmANLJtp1NRPUfhaI4KH2yJ4U/U
REE3X3CjKl2zVHrbLwb7AREbxFyHumRkYC/6ueLezomNT4ApnO9wIdAPh4Tv
P9p3YgXBnRnJTT0FD+3KY7/jaJxcjrGM+2LquWLEU+K/iZ5hL/xedkMPPUCX
FfElGSZOXKz0Lef0sWm6Vh86v+fLmXSSxlVZq3a1lrjIu7xKlpD4VU+QefpO
dCJO+75KMkVoqVa2FxbGQo6qAFPr7KUoT6b6R9BkqgSPYmwHHX4GmMZ7hJsF
l1wnvzUqJJteZMUjODG7FhHYOZN9M2uCi3RGuUs9Eazv1P8Zg6uOsCJpu/md
ijn7xgqgukMyQZ19izEesQB4R/fpnEaxdIKz+IGtGKF1MAgKkz4lec7ifyeb
Mf/G4gT4bpj+yP9EBGX6HldijGO7D/C9Xi0VgxnremHffQCrXTzXbZK3X1FP
+aLclZi/80oPUvDt3Sf99wqXz+vQWxUUtnrUGh27YMq7HQ2Jz1bXAdn01E4G
8SX/NFsvQj2AVA7NsLYsar38Va1E28wr13kN4pvU5DsGLgKRWTbSf2b2ABE7
0WE6g8Q8cUzGO50qpvTM8NFAJcz/uKHAoDgbCR7UBKVzacjJALnovaIPf+Aq
a7bEJYGP/joZhsOi9olqP9t6jIzS3nbs2h6UixSwLY/qyaNQB8u/NEgfDDWL
VAHYELhqjWoD7IRFrStLpN91ZwBUpVtU+Y14hJNI3tk66y+NXJy4yLio9UTo
D/LhP4TnCFiO/m8mjZ+fhwFFelu5RcnLlIjeBGDmSQoszCaU9iwUXJ/EQ+5m
8Oq8S0ct2yADzuzuL4MMVkrUHX86BvRtTeMdZlS2t8E67vpxm6AZTPOi8PS+
vqvFGEGuNIK8amdBefjO/CNWNpZh9yh9KYWu1HPDsQtET04kVDzD7uoWvuAR
DYP2OCB6vldXKBV0P/KlnLvIwPptqqJM7zS/YpSkKP1H6tWZ/SosfpYRlG3R
scRj6nhxNoJoUQbpuBsm0o27s4FkReIInNgECPyCDuzqlNCKDonSjaxy5ZQU
gRReOFtdZetSwGwrJcqX3DZWEFc3M61HS7tZc2MB1smNlsI48wKWjwzBCkgC
Yk6uU1qmw30jjPwZTIlLpqNi38QblqOqUXcrCIvzxKejuL1MgrgQS3reS3Tc
nUXJmWEwmtuDoN3h8q4k5pMsBxCSxrhDr4jg8+H4kpnNSZel18cE2NaYF5+m
1Io7Mx3tlOPHKXkji24qBxwetq8n+XedN7rcaH5wpOj3WEfMsmuSqPItDI6z
j8MBR4fyOkIlpYqBxMnMRAeXFg44zyHj5SOVkbG1xclkeEtSS/RwrYf8hF8U
TkVmLiYHgoSSu4VjV3yyOUxxhGrOvyss0n8F5ikc0kQL5mIXDFmfqP3ek/Pa
CpHy9rJ6skWlNwfTlRUy9xQYbJ3Gukzjg5nCVkGeFkYUeUkDOzGLCHGuCR1U
3gPXIa0g2knvE5g2snCIGs/AoCqc8RDB7vUgVvQMq3QrKu1fnH4pVeLQTfpq
pRS6ijC5LRWHq1eLWcYsa4DSKulMP/j4qoC2g6ZUlWeHCg1jPFSMgvPTqdSj
sY9VwC544WMpsbVH+WSJPbv4uDyO/fsHpw4BUlT4gXXT+zGCiVAr48UoBqo+
0ZwksprInurAh5hMkG2TcVqJcJmfKAQ7u+/d4Y08IslxblfaEwOcnmIde92U
gueluzbf+GtMP5lmRWE/eYGBS5vqV7Bulnxo7OGWdy+Uo8K5q5Irkgqh0MrS
f/72zmWqZc/fMdPUV8MkhNSuNL6Tc2soCGr2emFIf7RQXrxKc81AWKYRxzrt
fjEUn9SeimqUh91k70mqnzPsT551rIPi4HVKztDlLPGOJVHVSpigxtGXRO2x
F3MJL/loH57BocP8WxBj/3ForTaeiaCgR//xj+4AsJUCDojhCqIUxy6kDUV0
a/0IaufvWfM+3spHYDDiOifKCw4Wxa7lEVPpXUVZwdow6VHsPBckvMywSEUg
0h35bhJRMJxPZCMfb+QVACr3zG3W1ihidJuYdoLeSN92KjQcGLBzBZ7XNcKP
QyNTCHtIPU9jb8EGAgEcUvBbg/Jv6/xNfQSAcBUxuIQ215kj50/TYtT9EMKh
2sIwkjzHv1iD7/Xv8MzHo8X2CBGRAlGXQt7p/XkfvolutQuYZf0RU5L5ES9v
6ACA02DcWNk3GQXjAASS9MmwRglNBx3sywwFKlNK4uSFOC0c1VCT9u7X3Hp/
XB1A13o0qjdp7IEVES9FwfSOKsbF2WleMYgC+k/4rcprFlMsyt3wtQvmBn11
WrhmUXUjvD99vn7w/2YhhRPlKlpCTugdfeRUSpnTpdwQFf7K2h8hsbQ/RO+c
oLF5T28qtyupjTTe+YBTF1RgKMXcWSWNGA4GG31aroRI1J2MWE6hZmT7y/g7
HTgoMjzBALZ/MV8tvUQRPYEum8Vkj7Hmshy6m1Hf8FDlAaBcZVRqE7CDvkqW
K1f2Rnx4J6gU2DI+zBYkU02XXHAM24NyNUfQ7qYX6TymY0wmoC7UEITPhNHj
bLnv1zjZrGIS55BI9pfsTMxLpbO6Zv6OjNVOmrtFYIIHzfqaTjsBBXCPaD81
OrqMLnTZZam4vhCWzlvGmoyGkltLJGlStWXHe6Or8w8QqslY2oCUl89kOm8m
2GSV/cZt2Vjf7OoQa/SXZJUdxQn5CFCFDg7y7wYdhQdvHMGP1G/dVqGxjvRs
fDdnZNen1r6qY54VLXIKZAzHLQP8wYrplvhu+RCRUWgAFioUzd+6aEN5Ck8P
XoNqhjUiB789cTK40l84X5/0rTjL1v9ygUHHYPdZurGxEZT+CQhkN+uoUrNc
a6cEh5O26QOH2uSZcn/kqcUALltPevzHfLAMJsfJ3P9ruTKf1QchAANL+gV2
/ppIS0PcFfERBSdjzUBlA/yye9reJqqkzfdTFTAR+oA/YI6i9pjnF3e5v0pA
6LWQjb3q9fhv8VgwJThDouWqCquGqxZodgHajr29YkkVQEZoA9YLFIZzqWnl
8pXWDT2T0i0GUMxgX9TqX4i0UuDZm2PKW2/2Q6rOL6vX3sis6jRGTcvmzO12
gDLB23E3iEei9Konmg2pnS6Xh2zW+vab/RF0J0lB4N42aN4HEx20ekl+c6Ht
fE1iPB3f1JALfaLv3cUDy4v7l4Sakpc0AEYpEnHUBSpWQAkWman8cuBBs2fL
PHXixS8ZGL1KC+42KH0jghykiYLpHITvstNzhVXEAh6yVM0tR5rylcAsYXEf
W7uKwT2pzGkSGjvhMGhG5LN0nkkfHbyFxJe9nLsZ8VXf5gn+5VC42eME1UWK
yq6qa5C4xizDP//iFCIIwwM/A3NbW8KupSSnC13mRHEiDi248NFYCW4Ds2wN
6KHPWN9qNTPST5PshsdwGqIAsF2L0c2nTaImR8KSe9uhHDO9rBcvFo/HzNs8
BEax3+ULHimE57PkB/19k09QBu9iKncmicTbjmdgBPnwqV++tilQ/mLcoqOV
y4KpYb4xD3Z8/AI3YFRwFXPbkW/sDXRCmMDjiQjixYYtThc5/oHtrodvReop
wQEWneWDD+pitCZOTb/RiWgWY73XuqGISAijC9XmnIqFrXCq1V0KMQUXow+4
2zn6kbKVWQSaYwLT4IYXIPNvxFGEcz0ZMpsk/hWVWB4/fDBvY4uUPxTV5eZD
lYV1+XnHXyfPkOo8AX97rSlnasMtkOeO1GUxJwM4TkEKy04K5+Zu+INedqYx
W5f8amr/UiRkyfpcz3t0whcu6mhjMIF9YXE3g3zD+GnUO7xRHxhfVh2bOetd
smiDHd4xJRrmivudscC72KxhC8vyEIAvQJ5mm/5Pb4brNr45d+Bh+J8CY0WM
JV6yJlRb8JGSqVfgKPN1Yg/VUxGBFmJtaYk14OjcR1/cd5nmCPwMee2JQFrT
JFXRsDLcWlLY4BLILgqeGc8oU1V8Uw2NSvXHNPJvnwTiI5N/Dwc2XOGB9cST
wY99jMsXnkW8p1IZLJHf27SxuDp+1pqIGOmYZgCu90OK9XX3e4OLI1kY6lud
wDVy8CaYrFRBijD3ezNPf40iwOu95EWOfYQomuha/war0LQOYvl6wShDrmus
3UJOPEKVV/FFBMdilj9OgdP75TfNefBYItB0TH6dSlfotctjs17x8ao+feB1
GaA9H2LoZ+dLTgraKvyX9OO5gUkYDvqsbnPXwegTpHVpXpg4RBH1/X8fK9Ab
HOnFHtZTpCN/XCnFKgYEAW4zcK3ge9cny1/6SWaRKWY1NXo04Kfq/mM/4wDT
ilJo55PUn1F0I+qV6DqwiMItuubgebJo7Vbc2X67/rdvhCtoV6CQB6N47X00
LKJiCN+rEeaiBGO4lRR8BYJWF4qAWuDhW8hRtVqj/BVahGRmhExmM6fsVPXi
02ywzL1HtYsgwmNqmaovtsOaU27m1n/xR0Dy2xiKZt8Kh6rYOAt/Q8S3pUUN
bdGu/EXM3j9pz9JSyuMVpJM80voYKQGx5Ot2WJL95wstQl/QTyiigJrnV9L6
qmF7roCnhQ3IqQya3Jd2NJobFBsOk5XHg3VEnxvMK+ndd2Ya1GnySAFvE7ny
JtbjRsfb47da7PEpdGVr3RqengnOzfO0x92GhNmmvUR/oohXW7mIW4MBzkNb
+oRqk4dgvYd2beePJ7BfQDmuVGSNDZGTgcg1Wi8kiWSCXq7klsO2LjtAO7Bo
/HFF4gsxyqwGQchhhbVo2msrwN0sZ8cphQ4Wc1y5LsooFWDLdLvFFkRcHRQf
gaa6aEvVLuWnQrfw8G56ht8bKdQ10pHt47a4Vju6+Fgp9bQxYzoqkJl8dSXx
+QI7RGg94MVXUwOD+mnin/XXbEKVpfTuGUNTuWMGKDHTXBb1sHKdP8o+K1Pc
71FzP4CRsFwZYqdCcyL/8hacvJMQEaOEA/RE5nYeo8eLwE1GG6l7TzpKAoXQ
DXZnima+/Rx9qUOxNZW3WciT8nzuQxVTmjLCgHOFGaEPwaCTJybSCvMLk8O7
AWoI3qnqlt0THMWpuDx5RET6RFEJ3+dnkMDt35OnLMMgSO00YY4dKa5OiteJ
RNBbYELjV3/1NVzt8Qm9Y/qWmSOL+oZOa8ws3yeZS+AORVfL1qQF39byqN7I
dk/zXjy1/UvKbE3CT7yVfX70Kx7fcHfwNdzn4Np0QUAW+e/LU6JrGBJgS379
00kpZlSOWedJZuSFEnD5hlGMOm1e6nt74lgo9ClhAFCprFmRIpW0i+XGOHTQ
AJrtREspvoTO1nBhgBdGbC61PcTbd4tA3SvuGKKqGIW2pL8vb11UvYHWd9u9
pqk8kOeol7j4a1kbqw2gfweKLdg8PvTXQpo/oWAhRjJE/VZ5OF1s6Oibp1QS
1XTDszEofbY4qD5lP1tlDTVIiwBq+biuXJsmM01pHghofzsG2RtL0AJ1nggP
ve7EwR/KW/MrMbW3Vwp73QR8MhdDCB/9xff1Nh1ijInjfh5jrnetFqwQP3IA
5aHnlcAMPt7YX3+lhIPYikA/tp3rzhFmNqzd19vPzsuatV+hlLuFXMZ5gsXb
UM8iMCkWpVsmBdY/vrzMwdq5g8iQaGS7lfUCIkmvICkV7A2wreE9okXGa1x3
sQ58SmHKu7GLUQ6Cf/QoPVDNJAhhJ7XMj+nhB9UORuXxzBGfc+jGfM3AemuR
Xf99SflIQ+C0x4C+Cmq0acpFLg7ecTxzv7LRUc5u0dlVzJtrEv2e0AQ3EAQB
+DWWvh3BgJrjXTTR7ikH+J5iS4dW+phFuG0UNofJChYzZjJin+XYJaFtE4gm
3hFXioaX2gpNZFcZscKUKRlcDzqFmOspnGHp9UUrG+wZXiD82UW3bCkY35yp
m04Nyb66xRlgH0696HyJkt7CqtoKLfnF5MLD1ZGGXICQtKsoLd1nEZcPoJTG
VOuGf2fwd6gpIWt1bUz+zdHQAlUt1EfWsdlDhfDQK/WcDzILFJHUv975Ky/y
4fy1vKAMjUZLBNP9QH+8Mjp40Xn+lPuq8GYBQdF/ytVMEzfXLvIUcjpqf3aT
iXY2MYrkLZTvrTRBDhJss4QewWgqH/bcDS6jqvgE+skihhhBxK5IN/AFXu5j
X9rbNJVjU6efeezmd+2exD7Wzb0YhBwmwifqFv/phWkrCY5y55xD00NQO8PA
+tFaMTwdHm9cgq1SIJbvV9n8pPDiAHpdmzzNUXIkDbnxeMS/ArZeR9ghPsnh
Jxm8ppQC5JhwIqScy8F88npCrmpTkpdKxF611UO65pjjRr/9L6yTKcO3wyQY
Dq6UzZi/s22quU7Qux5oQRGGqSNAVg0DbCg3sX29GJiyDV3ZuDRqE1GcijMK
uvVBCIwzGFeNf43lJpo106CXnvFK5G5ztE16WkFfrsCtYNMP0ACOYKPzXZUb
mhoQm7kqEZE96IL3l0ZwKANSk6HhuGmtEWpj0Ai/u5jqcsYZVUTstteU9E5E
fcJ/Hq4iNpVNvDYL5y+cE4A0juz4hWNkx0xiSiGKbiFwcb3rhhECz+p7BZJe
rIwLp3N4cp+5dCWoPxzPyTE7jUxEXanOvowmo/324TprtIyKZSY3130Io+I2
VQGO7ksSFNn/L8NSF9TfgU4c1QBsyBwph+ZyGQMG3d8FhGHyBCKRC5pQNXDe
u1ZzqvBthBokdrYTzxdVHmBrHVI9/7YLuvDVrYgxy8mxdpGmeDyNS+uEbWhC
4c7TiY3TNiqphQ9loSjEJ+Yt6/32/wYQHTP9JAd7RiYgk0I1Mayj5RJVYgG9
trANzsamdOazKw66LK03jmTWrBnR7UmzZP7kCDFy79xCeONTO0lzecXrIQ3H
jF0I8j0XhoD/poEs61U1CVlA23i800GjZLsaWWpBSee/iLVLX/zQIVgCmz8y
zOkwLlZFbkvoQatXnM4Mnwfn+pqp1EfoILJ2kwJD3GklvYBfL6qGjLTFavTG
7e/nIAMZ3IhjvV/Lfu/zl7KFTYAOjnoWEGZ6ZkSvse3VYm9drELQ7pUm4UfG
E6hjYmH9ndJ4/yNeV8OHcaPhdyL8inA1LVsPt3KQHlrrop3aqEOIyhsqbYb8
OQKohbXp2MnkXPh/VllSdIJGtdj/oUbFYH9r0ojRRX4ir0S0sJZKFFlNTOoc
5Ijsf3gvGuff3N9SgFPfzQqar8czj7SMgHdGo5ROW/wteRZrY9U0h7nqmfbF
ksmMf0fyOM1rtuAiyjrylZtkXop2VBEl0u5LqCfHyc/DS7p08Te6xtT4VjbR
AQ8Niyeqv2ZUkGCFdw2j3WTBIa66TQDvChCRLRGE37+mFVQqNVDolavJRJh9
yWg2Qb7e1O2JlWS9uOxalm4/peOKNcLxe+ekrzi9EutIvFj1Vn0rcRv8Ugjb
BM+nZwDwJPOzu5zpob5s1mb3YPMHsmSFV9xhzWQOKogaR0hxImVsBK/IhXGW
J/RYGI++KX0qrhDAzUHWJVkMJKn5isL2P6YhDwjOtuA5I8wJUbtjQhSWWis9
qhiyVzsQU8Dy+9wcgxMyhmFcOfPeDQzXDG36Zsl84o6B7zU+xehRSCwAyXLd
fZuyncaWBavui4781Hmay03DEnYMkQVV+p0HEh8nMGlwyK1jQ4nASs4Di5D9
69l6Wk+rV1z/aEDuOYw2pcbkDsMY4rU+VcwGXioAmc8qv1dqRf3vcT0YobEU
XqYMg6Qa3hiWptU/Y34/ZJ/DtVlbaUeC6Td/f5SXJeBgVgI8K6UrFs0Q6m7w
KK8ZFM5sU59kW5Li/GB3cv956FyV336MNeFZT56pV+q0Db0j2rZe9u9nrvzJ
Fpn3X4kunHry85MYFFFZMf/Cvc1dESOsbAuDrS+7ha9B/w7a1/EXW10jX3n6
Z9pJT6negBfh2cUK66isgdGEfSwPsujlvQSZoHKJ8dLCXlBavDbWKmcizfHJ
dau+7q4LqYIXV8/VYiUSbN+ZRQegjUaNOAfqw+6jx/T2GqOZPne05Caq8RMr
VjuBM7lRaFg1JPT0i+QbxenNej5e1AqjCqTv1/OqXDFz5j0oF7NIZ4GwHnvD
8YYhtILRzIRnyWjHaurInlphOSmHHkqYnvOVWFJTq4jS3sV9uHIrJBua1zEx
t15DvBho3haXwjeYBuNtQ9D1YGCK//ZiZeWtMMqwE/mg1STMIXFj5SJ6Fb55
kOCKTw4sDYH6v0my5GLeIB4t6eHcbeRZgHEAB2muBjd0Mtu/Zm+A1EbqxY9p
igeRe36NzHSnUdUC4Sc6uhtkKkwnGsfm60CfJ7P8HT5qaQ7l9TFlG1LNEvf1
XedRmnvtm1jGuA+8LS5HzlMWO9fCVbI96NVBv1621piJ3iNPm+oFJ/Q5oviF
nF8uWpNl+ljElF0xFoTY4YBPubb0dvTo71nnf3/HELjq5i/rghdrufm37Cma
7bwoWdMf48ze6YHqM7cXQFGkP4N6R0dIw6olhV6qv+1mvibAvsOpjnKuJFZw
mVcPjFCrjKR20GahyukHPIdxjGPn/7jzpUHzZjj/tLfCpEdPFs/3JfpIeXWi
Ux8n3l8wajIrOoLCxro/4y+A+mZYvi/cipH1MTm3gc6EvKOCCerpbvI5iMv4
jb55S2SmwQBC7Nt0Z4qPU4EQb7H8EI1TtiVLM/0Qv9ZxPdWDLiMzWtMD4IFS
v97SXWiQG2loyy3Y1moQLizQn/oGd78raHokkr8jK16nywr4GcGbSRIbwLfF
dr19m5Iomk/c4cTCTVjoMD4MamXQrCEDE6OQweiAeIcJBAPqFBCAE2Zn8hvm
f7pLBsEYEHajjggQPjrqT2cSHyI4fh7Ci+f5Pi1J3W0QT3lFUAcpe14s8qsB
NFpCTvhlxm8GumwEa/4UktGtJrT2SqaE/yKp91+QqaozjD7HX9rmQ8RI33Pm
wGvpqfKvwWmx94PQdQoj3Z954g4jSzQuZ7runOT7ICJooONYZ9Puc+kGzidx
n8QE7u/a7+XEU+OjHcQNRi3eEQOuOAocBoTcmRBdZ2VQ/C67tZOWPSMNt7i7
8YCpbo/tbncp0RSu/OAErkKnqnvxD4uoLjXdpYuePbsC6i0CSdpsirKEt/Ft
9IiEpMr1qn4/SsvQawFwcfyCP6hIT3TL18clSg3UmpDneNuQiIIk5tI3c/X1
9DSDrPzHEibFLE6/hplUH4JoEXqxN4275GYca5XhGnNQtG6GnAkjnuupdwgw
rhXYo8IMCtLHxeZNQiMY3ZcyB5lCvHsLOvX8AZn5ISa3EdHzWSAbB6eY0cg7
XJNTefO35V9uq+WQr8wCDNktnNNWhtLOLhyihUvhyW+Lv1kCCfMjaEItu7OS
cnzgyAKK9Eh74ODbHS4jEMXjFmZNeQ2xo5ESkwcewlXF2pj+7SlbHf3LkgeD
4Rn25AvvI3OBBjL9ILhsm8S7ks05BSJP5+on7yj+ur8jwZK9Nig2xmq7KkQZ
sxrn81pHBBQD6xMN+CigxZah4ACG2J5UWXO/o8Gd8bJEdQvXAljZ1ApkOtsq
lY1mcJhC5jyGvaiDd7yt0A15zT4Gd81ZQac5c40mri9xJaRwAx8obHcRD096
KeaFmARIbJIan2HwPbDET1GJGjR61VccT0MyeS/L+ZLCcompF76hckGP3vfZ
DctnWxE+TIYstDOOAO8qGKkV80CbzhXsgLaQ2wzJHAGwYBkIDfoxe0+hyLxG
sIsH6WRR3HK70ivm/6i0C49JWUWcf3A/SmgFS4XYoZoRmYhQN5alhGjSRc2W
EZupX2aXm/8NqQhdcibnmMbNutBln7IB6mC1U4REeQQLPsdiludDrlZwYwNT
a6jhhJU9gT5KXD7HCvVry+/0W42NtQtlcM0TUVhRiWSylNXo3Rw73L43o+J0
HWPvwLg7t9XVdXm7rL7EAB6jHM/xNcIaC0GZOmfzeQrsdnZonDCWgxTQPorF
k3X0LFz53cyhtNbG99IZ5CUUALx2+/ZS9dBPoDRym2IVflqXKGmZQ56ELFVr
FL/L8n/NIhnDoyMPDuYrRwhh6Lg0wFosevR5oC48N7BBbR+udx3SxOD+7024
zkcPv3Vw2aAL0GBglSCbSM4TTNrdA+6hVZMO0wdk3e0OeJOYMxhKuuw4A9TY
jcl7svs3bsaEj+pxSqXijOpar2CzHbj2y58CLAtPytehx9cqfrAp0yeFo6CR
aNX0z+LnHEDLpHClOrOmLh/KY930Htz1idpC7c8BI2zcDYUAJWSlZlv+wue9
3ybqy1EMfiZsnN1kHnvMWU10/fVL4lY4mi06qFLICTjEV2Caz5RqCyX38o/G
jLVXRdGYhhYZhxDm7yqUo7KBoNh0dxoYpxkHsREeZSv29B2IHqJyTB8MB9fz
XUE4dvlOx1dv/diHOqrBOCOyCx1p2drl5jSyADvITevULWz9b4Dh/TtwhFGo
El6yna/zXs3NF0Y5cHZMZuHXGW+3OR5VNfCjsDMAnGA/xgzDgMssmOdYGeyF
r2+tSHIUw80Gp1uzXud+s5vDnw3ORdFzEaiDrYoxHg8nWH2mCgz76HD2UyoC
Rdiq4dvHzU3VjOrMyyfkZra6tXzpWZ6WRJLE5imTbisT0lUJ6lJWC7ICHgMl
kgRWwZJ+V/67AIJQNcaCefFLFGZ+0X7837ldxwKNLnwmzRctGPIO2jxqSUTA
mwSgGH4SI8M9SJBjtZbb2VM3NKm5BN+gcZb+SAjpeUNnVmANGrXQOnjCAHt/
6A6LnAwVLZS8Z3n2rfrj7DET70xGiMvq68zY+k/QIfWmuDdRc8Db2oD9eRAZ
5fNnWr23B8bj6Lz1ywTFraMNeDsJGHK/cCyc7oMh7xn6jxY8763x4YClpZfv
EeyqQoc4sZCPwTjk7B6VQqb8KeDE2eOMXeO3QD6P9IXCpJslxp6k7yr6VtkD
wVL3g1d7TUB7G6Y2qe8BM1SybI1N/yzL0tdwa1yg4HXGpCDIrPNbzsg4lnVo
5N8/KnpWvKow6ts3RoESQREMaTXQBYe6tA8usgSA+avZNiRrvsazKW3JsAoq
Q1k/NwA5vBO3NmeM46g/HheDO/1a3zv5TQ5yILNB1X/k2uZzI1+CWs2AEuq0
CPl3zaO+IqfAmwlh5ivFcCStZ37cGZDptupN87EL6ewgWAfzrDTdQsp4vk5N
1bQoSThf28snmeLfFIfhwlBR+IO4LuWIg/nQJvh1MRfepsCNOprRzhsc9DaZ
gl3U2H0+GF1qRJbwNWVrnLut9/4ERT/qPDfsaowhezdpAu6dqPo+PUdqxFJi
Ww+3nL0A65C+OrzpjGEQtrriuivSwsx9Lgo/JeBV6R10AJO+pUV9Rbz4Ww4K
XVjsKS2oYn8gI4oYnbgda7Fffp/eyGYfvs6OoErLQPVl+nPgj7wAA35p3aoz
Xadlj7T537FaGqFULd0bh7D/OdPYW58t+vrfYyt+/pz6u48jeeYISirLuV9b
h323T4Z/BAN9JKjo5WMuvrLO02OO+h+fh0R5HCGazF5rUh5U5y7tvcttzAnM
MEQK/SltdX1dBSQ2GQXHqHZHbbxxym7ra/Wh0n2cEGkBdwlYDUeb4UO7O/O7
2QTLkOSfNO+IX2QiKZkpKLAY5C/GMz+h0rCXv1g2ktCrYV/w4ykdxRAp+C1e
ZBgUvF/z169nT3Jkgp58Ql5xMuZbYEjwckcBfEuyhHZGyQ46uDEiGkyV5USA
QtaHsgzUu/R7doGUfd1kSt5I3DEpczxwjjcu+rjBg0v72pbmHTf+blo+PjY3
Wn42N4eMEPaevEAjdJZHrZ3W9ssj1AdgkjDnqHWQpZrMJ/JdRA44Ol3XGc9h
Gy5pfNgjoE2mTbR89wD6pTEejCxrRAkeyG9WBjjPAemJCdRAAGu8hNbwH7x8
SR/HQxYgbMzQ1yLlojCcxNVZsmHSKGuxJE4X4ReBCEYdA78SIYxEadfI+b7/
6Lz0bBOtlBUKLF81dqADMEa3z17d1OuJjoXSbT8oYqn2uyboTzt1dmGLyaWd
mtyMVNd9FfAlfpAxvOpJJN/AXR3ipuaYD8yP5UY7CdGEwTtFPJBkln7a0jZF
RJOICptxvYnnoTZyOLXohPV6SPPVSiOh8hC80an2/3x/fJHh5tlNbIyplUf6
vmK9e2yFs0oSA2zF/QayBm9Em4jIm0BVQWaOUf/KRxnUCEY10OpBd43qOUC8
VIUm+eJW0HE7lvp6Sd11Aq4IwhrXiT9YWA62r6g+vdzdNMyMES7icNsgppQW
I0X/R1RtSGJTlmU3so/5qvALYSyy4VHf4oCew8sNBOjWstb6HEWnhyRObQNJ
TPS+i6glTc6mksb8wP5uOUF5AOZxKPX8RlcgZbwiRttKQF83XYQXW7+nsZtB
whbTAdSvV9U7lf8gPy1DgpACLcLarM54PQyfZ3whftM5BtgygV1+bZfCi0FD
LekTZxoFDKFcFahTgRxo8LR2kxlgBY8TO7xUVHLG32vpM7PWGuyy5QQIvXkp
wke0wvSyAUODiSfgEj9baO6aTE7h55vlrcp39zAK7VlPBMqgG02b22/BUuVA
zyLSabb2YnaKL8ViGc9qaSz1h6PUBs1Oav0rQNRs/kxcDXfae7IOBtJbAGQ5
GDYpl5VaaCoaWb1VFjoEctfwvtNOdb0O4gu/Kvw3njw6Lsl/I5iwmCnmr8VM
o1y/TVs4MseUEHTukae0GB0hJf24Lp9tTR/1j/naTwHzm7oMAGw9g4UwQGoA
uYUKE7ZUiryx/v0bIpBL5ydyc3Gr1gCuGlv6lu/gzAKZXJhOL/t6TB6hGTo4
9pkIdKK0Ol2epmta+OK723rc1y9P5txldbwMuzYHtYfzL9N5hlu5FIqj3VcD
kLUa4lHou1Jibb9ZSEj0MF8zaKWOKoGe9X7qmaFxxCx8HvKaRoXE8ZPCvTgb
xveEDBt5PntrRDreg9XgzlGXif2npWkUngiJhIuitBzAYfE9lABFsoc8HCiX
M6FjpN1mBPUPt+59hKdlgu9rfstujsC9xKwkPbaMItZXTCyQ4K1hAvg3fHTS
Y7QOYRX0z3kBjzYn/Xpjph8APCO+UxpkPJ5RHHNfl+OSiuXwrOEq9LgBq+uQ
MKKjMauivEERMFg7bEIbiFaig2NvCqi9YpRwHD+6U43bk1lI9X5m2+cCrjCQ
Z2MaOO8X95Cw/mJ6wCejQNbf06YNk6a8sZeop/e5ZYrB6HcMUivfA5gRMTzq
1DTXL9PirLtm2PqEgUc314kM70K2PZk+a0wB0jqwkkGppSSKcW0LjXF+n7it
/hfWCcVPfxERK+VzlC221gRKr6EuWJaZl4peuKutqAA0YuFdiPnfIxa8F6UM
hVf6qf0CZKlpCvqodq8JPNyU051jhwF1OBqgYjVFz9pHhEdGFCOwJaf1x7LJ
G6xsNIo4/aSiBaswVPJ/Xjk4NWOTZGbtGR6pJtFx4YjguI/mPECw+Q7L1wdv
kdXZpqCZacjJK349Mszefya7+Rq6ybkMeN6/KZbkoPLQvTRoFRa50w5wV5P3
yAFKQ0w6/4ZIZXuE4xBHa5mGGUlrr6C94qZRdz3PSZqIDW2P9i0/4WN5AxVi
zwpeHXcmfKmmqMM94wDlgLcnQ2TXfsxv4PNmaeI7N1jbhNFThLbsGnbvRNKo
KgzJQrsPLotWKP6CUz7Q+n3H6eVl2RAH5sy6m/Th1N6mJptqS/FRqhSnrWhM
9wFLBccH6Zp5szFqmKMPnLXh5xyxosnrthEJbzU2fxKFCbY52/qIbuc3Ab2n
2eUuqzwSV9WmAqbjbiAkXLeJEaypnLBqXdbkKaRNbfHalN9m66pFjUtiOvvb
Tt8ECM5eiUC9b9v4W1C/7R3XyUsgs5b7rSRc7Bu4FJor5wTI+INyKArA6wQn
2Gn3CDNszb1l9TBYaVpmeanZl1wdwyOYGr0IPWersX5QpDB1tXjI9lp5GIEV
tiTRT11I3b6vkGLg5769lUiTE1q4cOzuG59/e3xINOOStEf6kEAdWjN6gUWR
Madd1E4DIZ8UIX2oeodPjiwbj03s45xZtyxH3pYGCxZMHGdI5Jr7jj/26tgT
8W70d2HFP2pgbbt6m7aukDPVUNlQMhW7eTMZzIYMujn01f1lZNMbi2Gvy8c2
7O0iUwTMwVvaehhB9SrgBz98zYqIij35xcu4e8TsKrL5TQrHjzoOXb0ChFwe
BU8ahUF+411j6F+15OuhJmyVV67GLlOyhl3upbm9l7oYNeFjaV4Y47F1PTFK
ZnZiEH/pviZ2sIul4Eij3qVU3KSwHftWJR0zUhGt6Qs5ji0qYN01M4foq+RI
0taSngnaiaP+mSkvZxXN+f6htjlCuuqNPwY7fyyfHK5UhPjHAzUD+VERq5zR
0AyKDAAijd7ffADQyAz48Xqo5Aq7tlZm/qv8W/WiYoPriVtQdW5J/gg+DgEK
lv+9qf1sNLL8M+ZG0RGyf1utDWlE7zeBi+3tLcY4salyAstBPbfUk7c+bN4w
goA/SBh7OUBVl8CI5Tz0/a1HpzzgxqXdntVT3h5GuhQZX42qwe+3Gf8JQEXy
jih2Tgzj9bPQYiGA1qK6R5cct495C4Lio+cCDGS9961bICR44uE0/y7Ww+2R
PkRADm3F/syCImxqZ9PcKkTqJpNLNzL78dCBhOOy8DFPZvoYbI/8eOYbDumZ
UE1HOkVzNeMB0aTvtr+hPVpDvKUd/QsW08D+C7Ejvp0IMd3me2hYl7Tqhwoq
HjsyrHTsFlsexb7ko5TUxomCCjt/yrnuyLCp+FPafgRmSofQCbg9a5HqLdcL
G4cI4luaZbvqatbelB0XJLds9gFYqlkVISsxFfc9Ss6ytvXVlNPCKBKz9vPu
SKJBsXvT7dE8INTGVjn+ubNd2yJpeBOtpajpkrorKZnkThP2ECZj0aqYe3Mj
Trt6CNghIczIP0tx7onOFIq6n7iO8KzOuxo06L6ZToqguf8i/XWsxZB16U5g
ASiAHDTjoECjy/ZKYjSiEFr/9qoO9nWjVDF5aeDodGmZUrbxO7qRzeeiUO2E
Agx6/Hm4wd7LpijmEZM1wNO8r4XyWjICwbchx7zRKcfr/lxIze7PnAdZ2FAS
9Cv1SIvWxU2IXUdbwHi62KcsEssNfZmET9nBCZg2LeKqBm/Tk0+YZuYyIkg/
Kvdat+biwN7CZhrB9+Up7rP1d6byHpsM86ET60rAJxRy8zet8TBb4+mT3TCp
iCElGBZOKRNYTewYME7Vmr7736bPR6O1rFtkFDk+UQFPf5VuuPebGDARu0hR
QITD+ruoQLrl8pe3lUM7nR4jLeVL4fYiuPGHwPkA8Lc6bCZ4UKSk/eyr67CF
cy1GHt1sLQEfjpyZK+x6VfHkbT6gLXep/3DjXG986IMo5PYTJn5zYcTQc3iJ
ItqZQ6vsNeO5wKD/XUh4XR1A2BsuvMSBKrqeQCzVvKu66khniMzQxlSuRNNO
R3xx4xVwapZUv7vS7FJmASQuxSjwURQjPsWD0vLAQIUQCJ6ZNGPD0QxBhHXJ
JlbRplfkUzQhJVSR6sKc6o9A0uHN4b3PeZWysIm2dL2mQxXqRxgVq+fKKg2L
HxRTn7WE2J4zaPBdB9+9MGHsknyiifWbphJl0gVi1AhufWG/jCicL4BE13dv
yuep+xgBy8EvqZj2xSzB4r5EWQw/vbN4BzZiZgYuQuBqZb/lzui4Bowww1F8
Ugx3lPy4zGeX1rSWW7q2CyolngOdZqsP1GZdh2T6BFU+5t1iJBd7ai+2P7YJ
vRUPHTR1OMtPTG0wp3Jmrwl1Fi1ZMxAxpy34a+Pmt7I9plCnUZ4bqwSbjEXU
vfaXJp+2bAapmV83GeRHoqh2BnGnyGEGi8/Brjwhbc9oeGN43t9SjaV4VsNR
2FL4Di3gOlJd257LcdXygDz0wM2y0trvK4XWVScfvLppXfdlMWQmF1K3qJxC
EeJY6xZPJaxL9KyZ2szZX0mkzvhU/40gYUQT/45OxJq3vcVWfwQw7WsUklRp
tFIC29oO4ClJKHlrdJqhbZNFrRF8VFPl8iQ3GKaG0/GqdXCd/2qGVt5cgH05
PykhAM9wXF1JcTjtfQ13ZpmsUj4OE+wjnrt/b1pau/XerelM7XXuM0D8nsDW
bgYjiBPEanih0lFTzNSkT5WwRABV3fx19q/C7zC4bYA5KwkvMYJ23zSXpchv
kuWrMU2C79fhF19v0n8I0kZvDWwemd/r5Vq3eVScgzLvv8DGEy/K5egfe7cp
33+P3doynieh19pG6K3YLY4aNAnyDgZKfFIlRtyeTC1kYdae+tDFJ/xABGHv
rCyVJfw0zKjTrftz7LAf9yjscl3q9NsUGG7ZskrFIoLiRpRKYp+589vcWhr/
7GjdPBLnk+iV21BjCYceDrYqEi2RdV++BK5wz9T6NHb//DHjFbMaXTa8Tim6
9wwuTEhOWRVZyVodaDrs/HJAUehy9gHYXK+tCe9bRzVKUtWw2UcFWKDdN9kE
5j8xO+qRTzXigJpG02NWU3MXoL2+bEDXLh8tE/zOD+GySOQ3nuuma1i6gCb4
28Z/u/4xAQfhbhESZni1shjdw0nGC6zn8aEhn2QvNzgIk/bwFmndaKEGd0ub
DCQXhghYwUaq4PsaRoEUjEK//HLow1Gj4rK6GmMkzxnLt4jjkOlb35Ue7IN7
W+e93pXkUPeBDmc1ZQ/KPedler0mjd4HVoHiGnFv6Px1bo1y3D6GdpmLsqgH
4v8P3qMmUqMtxR6WgsgE4IfAuseelWClD+j032GMEGh6osPR1rD4ZQs2T+sf
LM8ndqHWjAsM4FEu1qTdeTeduD5MA66jRXhw3yq/LX7LE9hw0Ii+LmPZLCcV
DarYv7s1izeYwM1RcHcv1wTtB7csk/Zn3sVMu8DYFe3/UNWiXDg0Tb0vCrWp
FFAnsLC3v/kV1eD9YTvn2Jhx46NH8d3gdxzCXh7YpZml4zEqhAymJQ1dUY+t
9IGTNZ1Bo2uf6T2ESKY7xlD58GjIIPuHOfHE4eRxzOhPYZFPfMcaSwBfga9t
jkeB8dt+UyuYwMpG9w+XyJi7sTTMEuVh1ukce+HgNAtWIU49a7v1S0NmpWyv
1duSdukIFYKp1P5/IKUWVRwupSXmocV3QMXmLgIT+GXw7qHSCdDW3o7clgSn
aIGJAPqTQD7oIKEWcI0weJERDdX7lt4fuZBHrU9csaVq7x7PjSKAwVaowiPz
KitsNEr2fU+Kuf68o5MRw4uBYyRo+JYuWpZ6/MyNa/XedoozzB26f33AK4FM
dwV52Z/i71ou3mU2RgTn3uTbOrioL6o5+D4j6HjuMvEGDFCQPxK5QY5HzRpb
6MHHq3nxDjYYM1Tb4uSV5bqtK8SNWnKinWCthIIkbaX50MM1STafQUOGIk0q
Xm3kDPpv5UaSpXh0MWrgWYVoL76Je8t7MzkFmGKb4MI7pmQKb0QEvXSq5Xgt
iQszXEW4fnD9UPTzmR5x2XGpLom+hJ4+I9B/0KIfvGymEAN0V9kZ416ybz2N
A6uPw9ZaAuj/U5m4RL4ziOhBOJslQPKntPlhaP+EBdSx5XcP4VIdSgXcSsKQ
P02KrTZ/ZEzYYt+yaFVWhw2Gx3G9jdOR23/2OZ8bw1u397zGjiyBPu2B1Kq9
QxJvYN1pnObdAHBUMOHeUd6DZtDG6M2PFJwhJZEIKgjyAFMH4ElGwHBMQbWu
lrHxTPqr5YN0ae8sBVixeGQQR2eKdKGHFOlMVaT10Zuzk6z+nfASVZ5jcQ1g
6MOlvjq5w3D4w8GXR4MUjvmaJ9/5hhZORLsU9KItLP4NKbEHxX+XcQY8UUr6
qapGfDPfPgrOD5rCBObNaxV4XumCgEgst80nc+DP8yPUZHK2AKbIz3brldxi
qhP6BTmqHtoSYnR/26coFkhsOIvdbAT0ld17aqRPd37PQvuSCTlfQVDEfEtq
Nlb5MJjb0ishw6MGLiNfYSTRrCoq3rywNvehIfmJZNxPza5I/LsvV6aCztIf
6lCA1sDl/u0CTqkmGYTAW7iOnnpjTAmBBKB3xkvizXsHxYZo/Ko8JCn2uoVk
xB8vr/lwigUcaGpRWPqfSapwFliEn1lNoq4EG6EsWV2DWUAH6LSAn2WaDUTY
HD5FEOZCKCNMKQCSIz9BAztaSf57C0KgAIVLqBxJMcUfY1++aURdZk+UN3VI
Xh+ehd1lQe7aQzd4K8Y5brZVPX6Xi9sfC2neOb7sw1Ly1SR2xdMc5vygrREI
teDTzqYiGXboJLGvFCcrUTd5u/bUft7aX34qwALcC0BrfoIASL4ZjR6DLAzL
T0i/hHWrvCrdIrd/6vIkCiudDFKcFSRpMe59ulnxoXePPo3Cfip2kth0qTkw
VbhyDDxxHGn4W6DrvxS62BDC0QlIBv9mLut7Wg4Yk63pa0Z+M4Wp4xX5MnPy
bogmoUqGZRj/LEeq3d0W+3Yjlm3k9KNJIv+3QEFVQRZx1tFLHwjZ5oOuwS32
dB4nOWMFM/4upvYIFX8hfxJs1sMLgl9T9GalSWIxtsUsDyFmhPnAF7fCdc81
b8JJVRUJCJ+LcCS1rF4vepyEeXXpQyhNxpXMBRo3/CjtQujyRN9qkgZ2umqE
Cv9176MOdrKmMrHhxWS3D+G+xzVUKADtztqRUDrEFMNTDfUQPXFwZ8Ycfvgr
sUBpnxh0qYHeyQ2VMPomjv/zRRRw89zuOBQ7KDg20PHQuV4e1pDtJiEKMaGj
e58IiMQXiAHlP1yDWXjcyNshpQ/mmUmsczIhAvAA5oeKXGx2oL0AGWG3i9Pd
regxLL259aCwxNs3WaMcgHFgg9CasKU9mmNbRT6bhYxyuP6yMh/9kE41P36n
VVr4v9vE8lhx24cY7BgfsfjVhyk7PXGSp6/Ylh1NdsaIA3yOEd2m0LQyhuOj
rU5vfhwnJKMBJnKNIldADt6QPnuZyADNPYZGNMuLfxUyy4qj4PuBbJMDV278
XBJfDggb7TrT8x/Pb95CPe/rv1wEiMG1f/fmoFT1/95pnZ6FN34F8bas6u3l
BYUv6x+KorqhvzdEii8FGjAtozUpLEu0QMcOfj6dLSuiNholZg0zklCJOSgO
xKyNLoCKD65RFzMxXmlAUpNnTXEbNlvBZfQrIGorgYDx2rWU+WZvQizlR3zr
yxa6Uu7TXSlPQFPZiyIRfTytgbaQQkQMc9Fke8MXQ3pTbUXpxYSEIWJle8Dq
rnI7zXkShOJBVdQ06VBtedRPxWqYr0VDIbIu7Q51zB196TmAb8C6HemmKgH7
mWIvW2IcBMscswKNr0cJl4bF6lTCTwL2gFat0bnpWxhqpgvov8mjIRPndleC
G4GuBWGrAQ7Ar3Rf5/aIzhhzvX2mxwDZL45RYPA98LRdGQjpLTJ94jXJh/VH
b4dRXnIeyDkYVO2xZa9f4lBvdDTByzht4ZdsU08O3rF7mj097OzhCCmoT4jD
q6kp4xuTk7rsJVINMkaUtIZiNxg7g14oRVEH6nQ0Dqi3Nx+cffxsUntQrowZ
RS0oZ57/5xH2tRW+qgzTXZWETVZQMocdMhIvZggQJUNqOpXb9WGjtt5S7gtj
knaVJEBWCk6auomiIGOiGQ8PpyIKIqqGshLHKUNgB/uIN9GngJdmZpny/3iZ
q741lhPrZFoT2y0xKIyoZ/sANzuVK/FnaRm58DBndrePEG4Y0ub5cH9fdoax
2UpJ4TdZAnHKiz78QPkpE777oNnLxjnMKJdOq5hlxNyIRU+U09IMwouLV0O8
aoawvzcG1DJtlYl4esEX09SKo49bgMT3Vs2kDTp3UArBhyfRFvDFf0kZowsx
r5w7hV8PxlGyhgGbcMsn2B2F6BP/IAxCgC2OdG0i7JAAoqwZPwQmVGONC/7k
ru4PhKIuhCMM+DUGYzKHWi0fI8CD+erwmfWfcXaAPZu5bsuXrSJ3XWY/rL1Q
evOUdcv3Uo1iVqBntztPXi/pHkFGoNYBVTvaHiXtZEqUOrEFBM7F3VhJ3Czl
nXU4TnGsuAvYXu/BUaGsld99KWTopABVWimEPdmi9I2gNlp3ZfVwePD60OE5
TnnMkx0k+Cb9//1eP4H7JEWJnrbGScMlMbC7tq7MBA63JDtU8G+Fck9rDOHi
sshWyC2rKEQV87hsgBEFOImc80cMmCCQvfJmnnVP3+M4uiq/9FTcobOtmlh3
P5Ee7TKSEHFYcJtmLEzQ9QvmIOA09bvU4mht2fL3ztE6AAkV7GkD6zTO1L5k
NTPXOH72DQFKPt7vgwhaLzbXaNB0eSXDOY3mHp7tAtpfeNY5Z19PYACJiPFD
0+ow9EDbAtTBvJrDKUzB7m5gBfe5Apj4KYDLLq8lVqk4po5qey/YufV0/r27
EfMBbv0hO0MlHk7qWz9tEJDCKcroiHKzHvohcT852+SCxBh+hD+U787PetQa
CDFZcx/4wBtsK4Mx/pfbTOxNMkRyjfm5BDPEPwPrtLAPKrLONCSYaDavzzrJ
GB4ck516rf9nw8SxY1469FSuKahPpgt5DMbEEIFgz9SZDdGdWx76hwe7Hs7R
YcdjmtBl73klQJjF1ClehaJy5E4tcamjubCdKPvdNkmBjDfR8ZKrYUBzAhei
PGTByM5k7uNe9Qu0Qt8EVJfXwyVUW5fyFbDXpqmayJab2F5/7MAF42i5Ql0p
diZVhAP2VS4U63AAHLP80yessaKX2V7wog5ysAsxbx22X420ViqjUF+ppQGr
JCZ5YzZ4gE6eTgNtxksibg8XU93MC/LoNyjwaPLcome47gB9PEhe5mba4Jub
ayuZeaGd6HuBsdn4bsG1Z84SQFcZw/HnEGcbVbX91Rdc8N20jvhz71vmhEBY
gyvrQc7uPMQXpriFp5WJ4YzW6JDrhUBHdEawdu14y/bMKt7EXDyRnnQ0NRME
UxnT0EeMrlmmUNfZjoetM4EIUP6OZAk5RSTp0AjKCXQeuCt2v3Iof7Xlo7lM
o/R38vvliEhjnGhMkYNSG5qpeccVseAhCGmakVXkJg9num2D/WUlaEQFQYAy
e1qddS9XIiiofVrPGLuC60Spi6TlIxEQx5qRwTLYiHbTNCDgXKO0+EPuXAX/
HLZkAqc+DLLoSpapjUq4+omJwhcHfV9rULc7JBMwszoVyiKLQuXIw53YbwSy
7VXYMl4a8k9Y0Qk7hYxi2uh4lw36/ZeNrNv3rAkkSgEtSIy1i1Qlts/t4L9v
TTNS5f4Y3OTZvrXLdcK3z0xMWYkvSeIt5peGowsKIOBopIjJGEog4iMMaD+c
7CjG4jLHCchLhcol3AfXvC6ut7lgyVs6fbSKw6WCcREn0hkLzKle5DidOJBe
4HEsvx0nmVVDIckTCkf2HIr4jN37Az3DVAY/oyyVurnxfS43g+RclgUAxpYJ
HLd06ToQ2PmodaJ1Reg+iywQKj6o+1Z6TQ/L3tyYJ8/9gLT/FaX9yLe0iU1l
/T5SOwrtozvbPH/gESSGB2eT1RVI0N1wrk1J5GvPPu/9DaVLcRwZFu9uDZdy
xmgP0Enb9EOWIFhoRpp3iS6/O16EiSvY6NlzJ80EGdjPuwltbhpOUS9EZ1pm
t2aPti4nUFCLsrjmeoxpC0tEr+loArXvojZJ6oBfHJ1gJUhls/arqz7NGriL
hL7QzWC+XtOzTmULIitLHHePdPtH2/ALdXeymlGEvR6XQWJu/JDQgHe+c8cK
Y7RMILEcJ02CzgbLH66MghgfqrqCfPvnyX7UgQHENoa+06lL+69PpgEBnePm
RaWG8J4E1e0+b+ENGyPBVdcdjMQv89dRdau37Uh/O0Hz/va/wYf5bdQxnK+g
xZe2NeG8PkWogij6h/5P50EiVOgBSKE+71iaVNlr8chzf6EhvabpMX8NJnZ7
/hHtkfDD5SjwqCV3O6TRqL69zzvxQsnZbhR5zJNya++1fl7Yr54N508c9mxT
tmrGXhQyhW9rxFS3YFvcSbPyjpTso+LLqds1Ql8JmPhzYBgtytJ6egmhoHFA
xiKFOCnx2u31XT8uC8F8v+mLtnmEn4QvuzXMLxnuyIT5e8PoIAw1oE343+TY
Sxh9kd0NJEMK80B2SDDb/g7fEeqtsUxpwhCpYTMT6VW42MsV//sTPQFPwKRT
xPUHfJMYeidc5KJZXoWP50wVE+RxoMuFInry8NfKVxaqqtz/nj8W2UMP3yNp
m9vnko2Shjd4OqHIju5eJuER+1cIwaVP+YuVxDDvkg8qrMv+OyMttw0Zk8g/
YZKJmFoxEx1TEj55rcZ6i/0BkRMdJjBMOjk5tJ6Dp+3iir9nByBe6xpAoJfW
aDLWvzsYQ/YCgq6C2EhDCRkbGQVEcho/oZ/n2JPp+Kruyr7mhOdtKi08EOzq
1L3vPzrOGAQpMSJIvonBZ4nCib9yO52BcAFVAs6EaR524VfP145rASAm7cSX
kwV0WtrqA3WajttB/IhsuRoXsG5KnBJmUBG6vy+y9s6Lz2J1P5ipsLUj/Jy+
GHk6FN0zhhphy6bl+Uy3J3kOKjZ3J2tbGs7bRqUclYMxuE+PAbIgXU95UxU+
NLCxEGGWRLxyfI7K7nWXV9tNAQ/V8B0nGSvYtwiBWvIPOkKOlNhUlTJbM/59
pBYOBvPw32zOo8jeAXDiKCJvzIOaSPK8Th9Hb5r6Vk+E3Gooj3rOkzjnmVUi
QZdFTOF3SvFaBL0md+0zDcSyk9GF5AiSZMLfZnpMKz6I8YUBPa7ZxeImI9YO
KLKb3gXsYBx+Mf++I1y4RgpRrNCedY/phvM3E1RiwfWsN/hebhS4VSQP42Jq
BAupU6BrBC8SfGFe03GfAtr8UdEw5LT+h/VnnxaXN0W0fBMI9mi9AXX2Z2Pe
CVCz1b5cEgtWzIrqTwglINoT28/2bn6AdMh1Hp9eoHmDj5x1ISaRJ9L0+nVG
Gj6pxNOkaEbm81kG0f/oQeR9irlU1dMsIPL+DWZu7m8sVtL9IC+HmnPyC0we
76AOpgW8wf8Phk2mIEZHql9fIWfC1MabtG16XXCfg6E9nls8hLCaOfJouAed
bzx6SgdVj2ZRrIqP3RJO7dB/232S3dJdw4kSa3htfOKhDMktk+iTq1044c8G
SvFNe9Lh2yJYZLLR6LY+rUXfX6a/hzAHfSKFhB07v33Rj3rw63KeghL/WboJ
bkmwcOanDNGViOzVz2FZdp7NsUw9nyypY2vm6KC/X1P2P18Zew0txLJw2id4
uA/UA/wx7i8lf8imZTxuzvmxjSW7rBbgTHF4+IfZHJQ9+u5UVkiRY3WsrUH6
Q+XzUCHsnvAtUiRgiHJdsDDbkL8FN83BQh2ld+h1RdM44k0EmedYTQas5AfK
mRe8eyblBdY/tqNr0q4KbZIFVto57Ce2tMNSmL95eV+k5HJ21CyCSt1v9vas
9O8NfA6lI4dKZAXcPwg52jtWJ3P8zIzdpAEYsSFzZxgGZ6hTMx52R612nEkw
R0C70xvzBuo4UM4fyWCg/VEBTRm4S8xvZFGZ3AT08uxJv7QQAz/3yhrxQIRV
niJeTivLj/sZ9swkElDXRbTjuTI7mGrlpSMU/r480T+nSdp6blttjk2RnxC0
pIXbRhSowE5HQcjbc7gjwv6gwTccWfFCVhV7jSx50XODxzfOz9AVixBeh6eO
Le2jCoapDqWTfZYPpn/bLvGLWTvmTex88PvZ2LueQ0H4ufZUeR7UpTQryMSy
rH9PhlwPtT8iIW65rm+81uIDHoNwqrZdRhSQEOnsx5T3p0j6KZkvqkEPbGaE
nYJe2yvcTyfVcWMu/VcsEnVRALsGCzdv4Cb0uZdcwzpzFMDpTfuhfmEeveog
WPNbj5nru6SeXZJQoM3pIr3eqLbr+9g0EK6Bd5lFJ5ATE9SixbTDw4O5n6wT
uqBW1ZEVggwM/XWnmrM83N54fGaKutbbwE2YHz3O4exodaSxIjXPL2dBA1H/
a+m2xY/LgUX8u3QpQh7JSK9bTea3gayz+q3atVLoUegWtj6GsBUifilUuHbw
tBIJkjralZu5kUqbKu9nyrTGDPFBPJxrcZu4gwbPU2xetdIHtwI+VkuQYwwF
nAo6lrMzy2UngRvLafLuRQ6+0MpSHIO6RuvDHIt0RQGqXmu/w+QrE+PEC0rj
qo6u7gmU8ZCCTMHHNDuBaXVq9HutFVhSu8DQifQihJ3V+Uyii179nYC7LA6m
905GiFKszm5zYeWUhAiyyrdXOLLC3RuAObdPfcuJqaOEAoVGfgFH8zGNpE0o
hBsMzdaAQ3IYqs/w3MNnzb4e5UGh+WefFDXhzMUeA8rDh0SrRBDUX9cT4dIG
FqjzXBtcuzws7oDA6VxiiMO5yhlWTaz2LdWvktEX9bSFX+e051wHROi3vdZu
vZtk7QSndPTAjEUOl+MjDeHJrhvktVx7Eh8v/5VRrKADakzCgKINMi1nISeO
H/yRc1bxRFjoQoFS4wNtSMFjrgniDJ5YwlSNQhVEI0G44rWIAfab8SWr0MoQ
zAbpGu7QUjsorXD59wo6UqjNwRalKpXx6OAe2hVtOSInVIdek3awTuYOYFoP
o6rLnEXwlm0fElKAQsbv0bcO+bK6vpe/8/caj3319LZ/2o7KFozWnTpsd4lf
9UY4YxUzZ+MScKDB346q0dE0iIvBtSORjQ/2mNoEElCkzm71SUJZyjctZMmP
QnOYZb96l4oTXdvO8HzzVHJq6+ywG4hyTiAo6BngZk8v2qnGW+2648MOsxJr
JH+NcRJ5CYXl926kiUNpgHIzAe0kWZ5vEEDkBckYWfUC+68szZGo4hFYrtgf
VUtqfaDdZTOSuIqWnRb+hePHAXB4LeEmqO/E7Uqx3qW/GGsjF+9pG4qRqiLp
Lu6UB+3h8aGhbXF/wbqLZ5dod7nIDGuNyyXvPUPk1DQQ2PwC959nxa/cHD4R
ig9lkmltGjDzk1FprOrDyDVW3vD61p2QsQb8mnOj8bKzH86OqFZBY71y7nKY
yYfRp+KCHcQI604GgEGwGjkkNvt4eZI1CFCGA0gH1pAyWuZJvYN6yXOniVd5
peF8SNcXYDaj58l6DXtstGBuemiBCMPj6kLguZppxBQCxcCM1BxIIipWQa4g
DkCYiGjoayY/z4axfOKTNNWadeoTbXXMQMa9cJ0aQKufBDrtTrQ/v9UH7eIr
ZAy9r3HOmvormb3o/TG9CBYNWUO78fL7/5jLxeaIVlxYR9qvQA7pHRl+7jW7
/rhYqXLRjsDfA3bXJE6Nato+CIYSb5tUWvoZl6Z8z29gpPFwcFmxOi8wQdia
6rfXHQ4Mh9yeiL3yni0fqyqtoHLumWUA86y2eAahNPuhAyYfYsFV1FayIdiq
mhp/G0Shb2oF3t+6T0yxcKh8Efj0iaba+mfCz+RCkGC3gHg+wTm99R5D4qsM
LvXt7crA2K/2MdL+HbAkJ1bxSSBR6YF4vGLl3JG0WFdOfTyx49krU65AP+UE
yzLwQL1Hu0iP3oS4iWRGmhHvytLGpjxyf1H8gHOyUHcsktCZgv0SrClZ11cH
LLPyFLlv3cdzwBwcc8MCUqB+kK85kJrA2b0gflxp/KpAesJHZJkLV74L9/Vv
gd55Z2ATOTOekxM/4Cb/MwHPA1nHddwHJDP6OO+/CgjNpVKGwDeuGeK3ze/W
eMq/w7Y3U0ePzj75GuI7khbN1oWF2SNgaHXOcfGh0px5Hs2LVK784yPULXv/
Ote/oEPz4YWEePRiZQsLz6yiC3JIRPVt1wD/6NabkbQ5cDKv6fTbWiPqZzBK
P6BCztPePFL0UZBohTfmdq8HnxB+aKIRB5NDcJbNRfI/2X7RK6Z6xBWLBrTG
wAqM3opRBhPbtgdoYOPFEqrEUu4EFPn7l7RuNwiEVZFnRIQqjGhqldg4iIVx
XZ2SuQ0YCZ/G4LKC6XA0sQNOypvc1uE1UciLeW8s/vsyZey09MTWiiK7mr42
RO/q71DeYE2A6+wDfbtt+hMJCnb2oR//y99r1WEnxaSMp2S+AvsBjdqPbCjF
myGEWytbURSZQnG2/ciWdhq+tcWJbwgf/nPyRsMYsqqUMPcMi9P7bEVNbRz7
fJ6Zy3V5sU+zhz2d6u/3LL/OajzdkBNwlIbtG/5TOyb7UzZZqoZy4cToJ2+r
gb7KSJjTNZvV4VBLDUPm5Bd5rAt6DKzVPGY6XKb1BcpAfHCwOWMZoZh0WaKE
hL/HBzMU1k5Qj49m6WGIpFp/OKLBAXblMz4o/Z4sw+fZUv/10de/sACB2C8P
qcwdObJz/aUB2AqspwnrZJvbot+x2B/rTDyM3hHW+XqNK+eVv2+eamH9sqo4
tclEDP50EoENTT76//8cLk+dw00pc4rDMKnnNOUc3Gufz7jMSrf/GVkFHMlw
kGGOyYwXPeoCW57OnauKaRTKNJ0oG/3abBbwtECtOIt7jVp5hWktGiArweNs
bsNoamJ4HTyfcV9TmOzSLoq/0H2zzRthG9220Vdvqjo5r+0nKZ/Iu4obN34I
rfbGJBlcz2ichyc+tnPHW611M/NsVQdkmwwv9Tn3MpaSr175uC+bCmoYBB/z
4WCYp3JFYAtJZr51Z5kzeO0/w2/gJ5CZTSp6NIftMU1yiyGPviEs+I/4LHrS
iSyqtJCYzvTf8LVJWeNN5haNNgXY/PQtKHjwVPfH2yoE/ydSiac4uy6f+MS0
lO5q7T+7NQ8xlh+TU/p4CAGvcPPVZX8AeYHMU5Jrdyu4HxyYk7icI7qqO5f+
gU0XljdT0W8wykmzlsU3em4bayWpe0YKJtZz+iE96RnagRNwjIEi/5f+gNdO
rHpt/tSBngyZU/y9PjjXmgB3x88BhUEm/6dd8t2bHMlZeVTt5cqWqzJo8qGe
da4d7m4Vlbpxw/FSy22tnHSA2smfUqmaGr7RmYZcyYHr2WosivNckPH0JApC
BkmntbPy8rk6ZcwRypcDKNDton3AX+PBlcsZu4LDrFlDq6U45bfErMQyX227
icKfyprWyDe5SmqMfN+Pl/tEpSmH+p7yrzTuLbh9SLC7HnGWE57JxfpXeY1k
CHOI3n3V8z5GU6ZOzZTOSS+Jpa4cL6WgZFqgLAnFjPLiproPWxwHHIS85bFs
/5B4DqESWbRUbVzfCQQsElywxtcjf68E5pYwnRIVzJ6DwG/wwfNZejfbCOlY
FGiIPb/KFNsqZW6+NcRiXWL89ZUBus/48Wpo7bXdppFUNzU/4WND9WAIjbqL
5Si/dPMQTx+BJ7F+bXtHkj4sg0kBOKVYA4DS6xXz9ac110rWRP9Vf/NY7yk/
abV2r7yPloCFCtRFeaPG5p4OsuspPqK5agRM4XAB0zIINZzunlsIHrnk04la
Ha5aGVVGrBCrlB+ZpVXZs4WS/iI2QL4ghDrV+yXqMtU/fugNGI4pJqRS/itB
RRlU25zwm4CWES3jyaL8fGKcX6Rax08rEGQviJ0n5KhRfp7x+3BvyPUsXR7t
oKfsNQyTkFiqI5dkfve8T0ZuDWsFHspCY1ad3p82z3Q8vCeGM0quITfZQDSf
ZQ51Z724OGRQrPfENX/gZMBehDZ2HZvWvR53s9ZE+AoB2MoB9JlxXJV6iPU0
c2J1ZJgQNOLQxWQ6+Vw7bgpzcNCRBp3oEYdb/U8ffJQBe4FB5d/McLpj4ye9
dhMNJCRIUssMqy63o9zrOIDuGqH5pnUUNixU2285h8Xc5xySBwR6Oj7AVlXP
b0kez3sfxLYnchtdAqNksqq2t39k7JYLiof41z6+BnYhHRXAhNgnYOkSkz7Y
kb9ex5u8tZ1HCJXMUSkmy0sUmYRLft9zPzOeiq3rrBIdTFx+PrzmW2XYuPSc
R18cXUMLLSxmthNuawmSINP6/Y+bt/ddM3yH8+2KpvgVlS+eDhwlcDQXPLRh
DGQDmZlEcOfDFx5paZxP+orsKVns3vRDBcV3lMO6sBWxpbD9I3BRCAMJ4E+C
vljgZ4H7NEkJi/W05mTqY5xrls3mycOv3hlEOoteQRC7FJQl1gctmdnj7Ld0
8iwMtolIy4X4cAVFoyMVzfAm4rjfJR3NkAUVMd3iGwg3LmJMSMv1Qv4mHZ4d
0c63kuoZlrHCHg+FzquAd6HNmk2PiTwk+v+VON4SjrlRDCq0aK7Bz/EsVT+8
+HeJWHDODKyljlBpN5vdJnqrehOk4HhBiaMYbqtqAkUGIBGMUAiLeMPpkJww
YrqfJqITTQW5jmXJ1gwZhR52BHdYMP2gsq8gK5I4FA8UrA+4uN3WwrLsAvvX
uDeOf40ttRZAixiARVDwtCisi6T2ygHQ992Nz5efWtufT5EfPHWCu9PxCV7s
RuhYeKRcn0wnlZHPItyHVGxakC/pSywoyIGfl8kYxhCheyqup/U5sbLRtr0y
O/PpozZHaL2b1rerYz3jE9/hT2EywA6kdoGaE+Zj0qabjrDfubdaXTIiBeQV
P27Zxx5KV8sbti+wVVgFUUmnzDWKp9CK8pYqibtOiNn7zb0gBEdaeFSuMEHa
45gkzP6uJaMjm424x6Dj+5pHIqyAX0JON9mKau0XZTUjZJGJVxA72J161srz
Pm7ggdRL6RI2K0PRPri9Nsz6YoHjkT1gYdskqmcSggXm2zmy1R9iiiJVAATx
nLmM0DB3Oii7IX2IL2Ck1Lrbx3K4Uh10X1Anu5D1ltczkZmmjhbtCji48lt8
mYb5EnapFpT7IOGEeAXBujkPQ5eoNsrR3s5axGA+9Yzm/6VUEMgRm8ELuowi
5q3k+Yn36PEYKSISUjnju0ITLFyYtBRTo9/TqBCGYw9tna0ixkM8oKo1mMrb
ddAREc6uRNIYgaEd1qWJO1Lw3KlHUQa7aDd0TNk78qVLW9eSUHAsnt/f5Wp6
d0KBHAsTKEqaK9OM9T3kKXLgnzK4nBET4eDGLxyiBgxVYwPcEbZ889UTiCFk
SV5kJp5dhigNQvteU8tlhm+JL7t0CoLCWbuXk33UE0JJsmGN1MWH2wF67AY9
TV9+iFM0zp9eWUOrUKc2Wlzgsodafk+z9Cr3MPUT4ArEfOS5Rw6jNxqe3AqK
LTh8H9DMp+Av5FNgISXY02uz/fFAdanU6p8GOPZNsXVtZqzDsHWMb/RQCoru
NZt8H+rXNtVYxdAOeY03/rnJMNytI+hyIe/bcBHIH5j3chW97tEPTUbPxQWA
pxhZU4X7LUHy6Z75fxZcty1oitFctO9BLQIIbsWPo+uSiObqAuefmQRi89HK
oHsxW0NzCOInVmdSkAvTXU59WSHmyKb8x9r7MG9A3yA2DCRrcu/jPFK5QPsp
h0Vxc81lqS46d8JrsjDwR9Jk/asyM1aKuUxUu+9x1VlbYs+T7EHqxmA0fm+s
TzIKLrzb5s27rQrR13AfyQlEV07Vn8uXQwY2f+pW4fxMEzfONSBg3LxNGzHG
1lY24ei2nIYvzgPHNH7SND2ZZnuD3DWLsGUfvckIRFRqChq9C/qN3E0WMtWQ
TEWdKs9I8Kl99PMhZFpoMtVpDTDFJS2pQfqHHjahipAb9Vy6QfDFCK2YzBgN
yDV0ve01muHs1/mnfhA0nPkicaao9k3H/ZmPUCJ+EhEzYi1G4Kt0H2auUGn2
CIcgu11jh0N0mLRj7c1f8Fe+rkTlrMVi29yd2VaKF4alprYFuRxINFMagZeG
WDLvsfE02BMSTFNYBUoNYr5TghJvApXYVARPlb622/tyBB5iY+Hk0ggICkSV
rUFcC67McmTvnUwefzr97ax5YClrEYDIJYuPKPD4Rfrbr5g+4JVGgkIZyn2a
3lHhUpUK9ks9q1s099J9+8VESwmwFXaLaULizZmiftWtVW5Ca+5FZneXqYU5
LEs01kTRYd8qui5F6pih2zdv5s8N6sWcrQWEfMVbEr7kLn00hBsbbbGEkPeR
7+/N3phVfPHMHJZn1UrKcjixx8dgQeENZ9xkgUTDA9pi1AFbd+uNmFAGVp0h
fb1r95kTjIZtLc7baVhg///zphPmUI/L3jH613KtNl84IpW+6f5G4Et9PXdL
GBJf90lYhxYaSXPKUfL3I4OubIl4LI7x/k76+f/F2AJiQ4Gkeu+BNEX1LTA4
evWySf9m5ZHtFtsUq2BaY/zwGYoYDVOj/Oxu9fFjYlZ+zZ1helwCNwrhvhJO
o+lJg1Y4istG7ysblKUE4jHc+qv6MK6nUC0XmepFIzyq1ejiL1VJaVdWRh7f
1GEMvgMAaVjESYnXhUwKhuNtxxnUwk8ysKeqgfy06HO2dImlhj99qjM9W/Ii
EYBwXLhhe0+8VgaNUB8d8s8b+9v8y8P3fulaN5Yn8b07gVh84vSaTp2XqaHT
AxyJq3af/Ztdkh2aPHFtnWXaU3L4rsl+QV1UOUm9GAI/V3OJdsDhAEeC86uQ
qHvaOdYuOepXtoA43Mh5Qg+8W8fqmk6Us5LKnjLmO9xwP0GdGYjiJk5OsglZ
pgs+j7HWYc9Gp9vGJntzlwQChi3rgFNLXJijp2P/CgnOezWhS7sLxYsoz2aA
269dBxMi/NEyAHtPO+H/CLjh4eEy215NqM0cvUM1dutN+OcubnOlKEpE/Nvz
/g6aRkem4fjxA6CCfZtkjMzJKrt25E1hBiwq6LEKnYlHJ91H5sZxbAG3chWt
my1W/xkdXEsZ+11bf57g3IMM/z0AdqIR9pAfpEuLVQqXdYOW3ngwvNq2Qkcz
XsXZoByaD9sBaisnk2A7vglTFBrPOAGwhQey3YO6/K23D+GyKda+vrUFGh3m
Ogr09/i/cyxwHje5appNr8gWwZDoKkNfNBO+b9SU1X0C4IsWC8WMSBWAFNun
0n8ZUVFEIhSawViZnkGZnURIBbdF3vVy6/0WFgD8v5sf4NaLcQ6FAagDTTgJ
IDMnFncnAJFu8wUp+5t4JiC/b3f54nMZ2wkk4Z0FCvTZRMP10vFje1lLp33m
2aJcJg0o4sqsvxsCtyMVA/E3h8+5abpkxmnt3RAphdr3mjTvAJ4WqetN3Lzq
Y8Neno4xoh/Uja06SKPELstC2rn8mP94dT7Fs5hgMmjoxynSdmqKl1KwGrQ+
BrPtQnhqWnQeqn/fQ75xNgqCO6IS0jK3Ueunzh/G0tFN3mGSaWP+GZ6Rsw9n
SVRiHRAknHRJ09d4bYC/sfF/PmrOcNFAy7zs+5P+T86VeoQGUUokDWOou/NA
qy/rcZ5ywrpbDUxaafT62/GeG1ngcDER6CiLTtZRjkeOvwqr2uGw/s40aq+i
iO7Ym5ve9aKaGTLGyJqWBpyVYnTjV3L5WfnsqopDQolo5p2QBp0DxbHAl31M
b0HNc0WSvBvRrEo8MyYfky4GD/kUNNo3wqKKyG8MdGZaRbMVjDw0ew8me/lU
+A8XQjH/NMhgd4jZRJDEXgQfn0mlWz/3nicMjC6HI38TbYUqCfCRZ6Poh0gH
EoEmDoCMsx4PSmnN/f5wQLAbCyPmeViPlDKmz+HPkqmhVzSlC7TjFUcYAQnJ
zsi6P3UH0ZFNaa90+lKeafasQX9nMJ0JFLMuott8FsZPyvytucSPWihblEmA
sZ4/fS7iclfwoq6nYF1bTq2hX2mI6VW6B+v7qsmibUtL5mne8yNkF+Z+JaaJ
Fk621R+eM/WpzVadatL95EqZzLZkQz0LmqB6TgaRxuiH/NPSlHb8V9uygLRP
g+5OtWV1ecnBvicCf3KnkjaeoR/JgGapqIXFB3waqSMXV4UEuY8hGg4uSsrY
BMhcz2sKLbvUBxl+vhYqV+O4zSaXrPz6cUh6CXSLn51+RqLh5D9dsIctkmT/
atat5QMalxOJmc3m11oFLFwcDW+zYL7WO0swdwTcYdQaVKwbJo/Svx2bdciB
SY6MRJDyZLQp2k7L7sbpEBeJ7T/g0xrSveFPMf6w463zr7J+fXnw42bOfEGr
Oh70Smf6Ym0IOVWdoFK7OX7Ylqzk88WFz26+yeJSl8uOL7Ka1fwLDdQmms+N
uq3mQe3DODRJC9Xv/5vVWaUlXTO8cKcOxFoTPXznzjhXgzKojn0FlQUxWdiW
yc+YQc6B/yKfa2yhZsKvQIVa4pDa2kLOmj5+xqEksqpNp9Y5+VbnH/7g+Uhz
Cha3Gu/KQHN+qXUFuAdYQJnObK13hoR8bXKI19i9EHAj7qS8Nyw3OIFlGh8a
2qbCriMj9ucJdZTB8b4wc1S28tsQPXneGJpQqVV29QBUbBk3bL5z4D3RKr/u
GP4KfcpE/WO5QJDwV24BTjdy4Hy6k3n1USlaJKd19RFnYwEEmQJt5CdYuWF+
evHbLEoJl2GElEPqMPI0UNP+DrQEDjDaNlehwNymCTW2eea8yOJjAOAz/krK
s9sniqkEW6PIjDgDqxrbB0TPPtKaOkF0ZEIY9RAdHXmZ5pJh/XRoYA3fbkuw
ZyWcvX65x1CPC7nUYgTwn7XRKPyre00AmfmUzxqHgH7QuxjWQWOP32NcIAEE
TUpMbzxgtTZHAFWWFLtd8ZOAKt4LRAqGwtX2WOVSOJS+aDJ5TNB4cy6wezkk
6KjTXFx9+Rael0t5N9+3DrgCfOZBtAZBXwIrmNALoR6u18wsDF3W588foFA7
fe2rpuooztUUGFN764kpr6msWQ/wPXE1O/f8g/FDvS303JrTOeIETWiiG2vY
GuFPAtbSOqi6Rs9IW9xcur38MFhMYrnE9w7bcN/+avbtXjFdp0xEEk0CpQV8
8eL7aBcpJVcJQGnnsIMiqfA3BZ5wVdFFWx83M7U0lOfznl5oGOIDXQ8rv0lh
yCgFHBnRCAGkKf02E6uxSdAXdQl7tbFopUqI0b44CCo7dagHIA5C1P66pugR
OY6dlbDih+QJhxBSXraidQCiS0AuL0fzkIOwGYPLVM6s5e0P8IB1yp/pvwYO
vL9RAJPoB5rZnMjYPbMGqXbCAttvTJ+i4Y7MIsquzrA88hpINVoUlgmd83H3
D/cnN2ZJCY9bkRmoAqgG5Xrth9JyJqF3M9KFOUzaXoMxyxC1iNz9Cy5yZ94i
61j/A3KCAXIDQzGo9dDzk7MUz00sdwWCvgpEcCD6N8px4ffH/xVTlV7B9TSJ
khfc8I5WGDXBTuLgDW0og0ihb3grVecW/zlVkdPqb439mC58EOcDa+v3ihWO
XUIxn7Odb5XZiIgx6W63CzvzPbk1HKbPrPY6/z6dH8tcMmFjwmaJslhb5rTY
2a74q3ExPLx6wW0jVkCUUe2NeG7V7DE7GP1ppxXCud8NuTXTQHKwDDTc4IE8
qcZz+wuaX3rTRJZP5taVjF0gUmNY/JrWuAHkcY3Gvr6n7jRw9xlt3ZJ6hop9
N3IvCgL66kWen/r8zqKmiVDipLPgV8vLPTAM0JCziIpZMNkjpTYxv+6e8aSZ
1Rk3Tf56jTsN9/g1QbX7aSwVL9n4uHyMVfbaJi+AiPtVy4UFubaCqOgqcM1Q
SoxI4oPRpvO/I1VVMtuhXgovkRRHZT3wA7ByRswuh1+nDPo5PI2jndHslhh9
mcrqq1M0nlhud9y70dl8MLc+Yn/MW8PJhDl19kAsOVMxhqwelSV7jKwXbGag
LLZDF3Gi6vHqIt3b+RVP2sihXfZ5iBZnCR/BiEYCbch3EU4TuvXWnhnMErGF
EM1QgmM5Edcau8WyZEbWivvmPQXgjPVzA6hMr773cm6duxUh4Qjac/IkDqjH
zV1WE3CHix92/WUtmKxITnvzHlYoypBamirLBa/w+A1hm4zzgAXtGx0KYXs9
FHLLsnwb2O/e66Akx1CELnjhsU+GOs/qhQURKDs/rcr4fPnzRto6QjbaxL2m
y18Dmn71NtZahTnBIjAZeHai0gXAwcP86Jrpi6jf8tDMnLRIqpUtiZOBSRv+
Ww+Ef2TO1QJe5YL6iAiFdTGtEQzBtt9JX7nAmfttVubEnaXXt09heMsWtHWY
nSnqNqLBbZ+y90uuDpznyjBmEPnKUyUoN9ptPpHyNJdPhfIzn4RwF3ReEJXy
JsMsIdYTq9ypZVUvCZPNNo3w8DJJkm2W7NIgowNhBTolbHm2hjSibcNIcb6l
Y5Uh23Ej2Jre08BzT0x9Vkc3MsYTUKmwc82JW9NAETiggpMJ+zG44mggHxCI
20bZHG290WHRvNHBtMvNCz4+GT74OFzZdW+8GX0szJgU/pdkb3U3bkoHBViq
/D2LpBnsWeiV7qrlkLVFQ++Su98gXn5VZqVmSwe+YEPBPModQ+nv8xVu5rSi
VJmZD+DqnPUZNFxp2OJo1Hfle2DApQErPk/aBjj9OhB3pMlwtNX9wTCqBdwO
stZwTyxGvuiWgSHRxOBPgIDWqzaAvAKbsck6JKbffjR6sTt6d+KkOGsZSaMa
8GuEJ/C+M8XuyG7r1ly3/gIbugPzmiis+k8J/bCy9XsHphZsQvVB2h91HC/E
icAUjp4kPoB7xQZDPpRMej0pE8dQrDNWGT2DlR3wA/qgwRAgvdeg0IMiasDl
6XeLYdkwGQk5bfcy7+d/enCWHxlqBBFDalCqWVrBxZlY7eDnp0it4WrK09TN
/j9EavF71nGNgAR8gOuJm+EsKJk+NuuCM2t+iuOIvjrRtDDhEiNxeo0mD+7u
hmvqyR8CO3wzIsViu/LGNX4Jq029z8uTB6YPvZcjw0TeZ7GmFXYFZe9T09Zn
H7MnAiy/OAJ0cEH44icVnsUiDq+9vt9jm5r+fstfOY0g3RhucfXpuAvTEUCa
wxsmjeWOTEQq0kmfrhlBJX1V1lOGjXAgu5UM7Nm1xo8JxYU9UVZdGbggbboL
s1gKvdKzemcTqoFuc+HxHmcJZrLfHDzFVtApfZR1/UBSP5q4EVqelXrWbqNW
gV9aNCA6XuHiSi7nDh8QcXUCD6sfUGRmcK3wGbiqiseMFsvMPut4rHdKMlN9
HGvishJlDBlqRevwrwEB6To9EDTDKGRLAtyxP6Y3OjUd23Fs6r6/LTz5lXob
IohxIU+5S5NsjDZ+ES5O8yuWEt13LtKnuA6g2nnsghPydusvWc2DHX/lQMFU
/x/g9/JpII/VKJ2+qvPGCVqjaljG8hroleBhom4Nw545Xo2BsILYKImDrufZ
yVyH44qDj85hBzLbk2FNsPX1nsqfSygNo6fdQQaBTkEDAzmACnobnPSPqgGm
7KclU5+LONq4Qk2T3XnGSnuFWmEoD6opqZ+YBPq8mdrEjfZ+LKh+9A2yNAL3
v+nC1G3Us3L52Nok9UuJWL1g7F3HSDyixuchj3InRHGGP6j1TH7JYaYYFAJm
TtEx3fzFfZ5qb4m5z2d3w+Rqe1/dpmwGC9hKrzDyc0NXTafgyFG6/M7/E1pP
eraDiAWogi4vKdk8wtcls4tiW3SOw24wTtp87QWU/BzRJbmmEzmoRiXEAIk5
kMlKoZx62BOm9C3Vgn1R9bCijXD2ziY9YGShwgiKkuzuxKM5QlG2E85E5xUF
YlxxKWNG0xMtwsq5Xlm/C+T2m4bN13uSWbg6o0iClumuIjeA7EiIhDgqYNdr
RNTB9rPTdEVjSSQuR7qo3YZrUKoFsEXJmHMePkFc52x+l3MFiiLfOjGMMXnn
kJM5jRBiIgUkRXZTAMaRWbvi8wYYjpZ0HQ3Tj7q3cl0YlFDUfORmgC0Hwjfh
a67sCKk8RHTxP2wqRBtz/rwjJiFar/g4eKIFdX1Wi83hGEl2oaknWcMuwoic
hN/i4IbjGR16E1GjMt4YLWMl5XY0cfa0eXHIkdBxZOhGF9aYXQxkCZy5v92+
SM5rlxLBTkpMVEEMkvmV1PPd8a4vqUxNRP3O+Mfwgen7zQRnplIPggD2565f
JwtkmRGuy5OiOSDKMgj13uCboo5ZLSZrjhgVBJEA+WmHYKta5Sipd6WlJYGq
K+rJ9HMq1vRq2un7mrtPHziumyIpRX7OCP5M9OuwPcU9B2IZdJ9oO3WGAdsu
FBq6c2YbUm/W/s7v1UJyp3967lOfdSa3vBFy3wrswMTPhnfF0GTeMpDtY2Ks
RqPZ0zvjNQUxBS2z8eI8rKg50QwnNcdMn/BL2PQalKt6KVUN8TBciWbf1Y6z
4HfjkPw3e0SoFTkb2t6gZj9s7/5eeX05cZ4rBZYv+5M/cnt5bKGlpKJqFWEW
DSSJzAlaqrYcb1sJQAh9RPiYrqBjXjFQqMk6ehJQiA6Sbr2VFJcB3dwnLiNL
4DwSt2uSbxpAcuvZrOdJxZ1ZzfwG7OFGYaKglzWUm3YzugfKhMsk/2hV4+GN
MUnUzBKajtv9MGffioC6Qe0p3h4SdyfyfRFutR4OcdYcxPD4s34u0mxiLi1g
eBSSKIHaufxWPGYpeMJNspfWZGLzsM/b3gTOmNCwIgMeaNNYApDTUlJH1xdW
t6Y3gC7E+Qp3ekq1+AG+YCSohUTuD+FqC3RRiixB9eKeMWJfWHRAfxWBmt64
/OCvruVwymBpAxyA7xV7afAfvtRdwUv5TtVnA6299HvX0wshBrqlZYuLweu7
9PNHf3XTGypNDuI76A+k7UW9uPv7lVCTzrTJyJf0/MFrCUQSqx5CfqB1QaGp
New1EskaqDmkvJeKbA6zlpYPMw84Z+vIvPNlGndwm63E5C537Ig/uiikioOb
Im5wyryqSvsVhNgDFEPJrz9RdE78j1S3ji4G2+KQo1HezRgLZ2mEssoIa57L
B6N9K8S9tF5BknV043MbRN716w6pOmX8Phg79clLOjETj2GunOjay3T3sQZ+
jiCDqRApW2cO25eYMB9vxk2cJGE93QG2vhkhrDqWFu+oH23sM6rVGFFryr4J
mrtRY6QklwpRtrG+A88nXJi3BX+HFaXDGLnhHzZTwHq9PXxfdhwsKaP7YeD/
Ydx/lyTc1KAImdyfBzQ2MB2kchoxmYIEa6eJn/GKKzVWSJ1m7SWdg8pMWf7L
MFacM8PhtwW/FTegSYEgLgtp3Ny7NfR6e+pKEPr9Qnxl3PrsBDOOD514ni+Q
vRVn9hBQm0b6y/UbHOH9AyGOFX7z3McokdgUh8W7giFF7kHpyL4QoDPoPltO
9KfMqHxEO2MnJUXUPQsb9tkDPnuAUlDuakJ54xxE+sk2d5lZEb2jaywz7Oi4
WPNuxz5SuZ3OoyJj4EnfTKPzNynKj1kU8e2fCvng1TiszakJaJe+RWJk2CEj
dyHu3mZPVz2xDmj6x9L6BaAy3HNUVFw5TRVhTdAGbhwRiyRA4G/F8rOWCzU5
o6ksG2E12Edw1XSZR/599RF1R/7n7uXS5LcsqwmFI9ygOuXSrb5BmxzR+S2k
JsTAVwyegg08AJukPuc81STCiFAQj6C7btfTs4D24dJEcCXwwU2UdIBI6mmq
dwS2c8MIh4fhY6+eyaDJ8w1B5aE+iTEy6WkDI4mUS3Nu71HHZ1I9OFL/o37G
lYrBPKHxO1GKMz4gXpKUEG80eig8GLpKKJLtduVPv/hZykwsBEEMrCilnBHb
HWKmWBCmMBom/sVwqMFHx55WFdoVdi8Zi6PavSvjgc28wL1hftAJcc0avFba
2+AEgUW6d2/NbTJy/b7rSTLYWX2NQPl98IWnrEARmib6+N4gFiGdBbKq3BmQ
X+F3IWa9i0XzE1tJZhKz41UNFLJI7NXlrNS8eiHWcZVlUgw2roZ2tLLA2C0P
k865o2An1VvV41aP637itrpVh5qUrTM2spFLxZfF4165fYMRU3EEgDGDSDIk
IvN3aPaqxz1xL/i+/BW1mtsQQ5LkB9QTHxANdmTfwPwcXDfhl2jpM67em4/E
xlEu2cKcGiWv076L/DfKLV/GJW11wnitscjbJtJo/HNX/a0r4a31GBAXglKQ
EfYxvNOatBFDMkthdHEe0jBqBPykeTX54h4hrFF74upd1u/VZbNlUa1ya6fz
MW2oAfR0Mxdvs8LinnLHt+0fUYe+zwxTtuTp30vD0V64ntRyAthWarJn1aGd
Y+veKEnPUL6gyN248J/x1j+djNEjqEme2fErwombXyyw9MPGWrIEQlciD4TU
+FaU2n4YbZ//NuTi9+BBDQTI+VenQN4u1591zFpw1ostbAJYHJBa6T4Bpc8z
uQnBttwbqf3dTh+8STl9gfVZ6NHTc43aSeBJoz+AasZkHEBaRbbA6cRHISy5
9RvrNPsoV1sGWCAObr+GHPI0ypr7EuHbaSkal3EeIyVPhepBzEHJ+sd+MSoZ
hYGPyzOGZWp3IVm+CpgYwhxu5BNo7sYBxAdjWRHpOZ7IA1vA0p5T57gqwB8L
S3XXO4WXRz1YxlWtd6cETm2silDG6tIgYy4unvf/6dNtWq+YDCg0y4MRxYAr
e/nAkZho31qysUQfXfacI7wNCeDp0KDPemGz9mzK1/13EqAVX6jy3Gy7D/0e
R+ORNTVMNHeDR6U+WwqouiOMXZ6fXPNPzikEWKWBPhvfkM4JTtIHiWBxXAPH
rTPMIRktX+FDsivEMados1gM21LTN1fzFHVzYRHvbZKIJ0116hfDMeDzfJaR
Tg4epUYWO+nuet7ucdiGAvShUeglJ/D0qbFl79j54epZGXOCWSP4QuvnlaR6
6XReLogeGNkz4pi8C/wCBHO/OxYq4bsYKnIx+znmnCwRPm/hvL2V63TldJyw
T8WKYw0t0R000BuknlRQjRkv3pq/sREoRV+9fK6nJPUGw9Zkdu2/0PdNEn9D
RuFat6JBx/vcY8r/LzwgW6m56izkg8VaRhihb0OMe7U/0x+DKfb2EXps1ZXa
EtOw+nmz72jx5LBs+gk45mdX8PtC/3vUmoiyb1L+4coHt+PqnbCgdfP+QVua
gFdIe3GoVAJdSUE4tdIlWteM+ZaGFPBmU7DjKai0iUkMsdKVENLoGPMl1wan
OpGXkAhgnsRssr7StkeuP3UYfyo9NBVxmOKEthDnukEnAhTp1zhmX6CKbCGO
Co1bs5VK6qS9Oitpo6XR1fIdzp6tZ+y4o1vUXBDrrKGAlfp8a+g7qInVcfA9
vFwU/Z/gvG1PhAlgPqkwHSo1GmIIJjIjot7uuLbsUlQtN8QlvBMg4U+m9/Cz
12TT9RR2EecSU3EpbzkCxqCIO8l7XHNVHb1CXr6VKR18w8dMk6Uj+CpqtxV0
w4kwrhj8TUhN8QS7GaTZpjz5rOynO5sXdhVWS3Z+9G+jqvjBbkW0dGNhpmPb
yBAl6v+nTgpTZUlZ5jc3uSkjFKBp/mopAmmzmJYNO+kokqOtiAz8LI1fCXOc
RHEK5F8KmnpaeuT7x9sdPXdCk5C6Au8YJRccqraP7ak6+oc6h770KnUbtX9v
EcxWKq/buXORB/d4gEfPp1SJpDYlIDOnwCKzgx9Xk2EHPrGWRbAymXKCFNjr
GY7hrkqUjcyXxhHVQSECIEjt6mHkGnSprCLxXozXYtafIEkc1RY22+JipKwZ
NbkIp2daQSpWb4c89BpTSgxng1mrWewNmr9RiEUe0dGStJuFIYIeDyaWNkig
1Se8BNA7yuqPOiEo+AVVCgU/WEWuXtRdKMfdZ7aTwJ/E25x1fK2nxZcX/Ljv
u9dgdeZExKOfY3EoBKcOj4Wq8CKA9ZdSrVdcvEOSpYwjj+iAq2mWAcgw6WkP
3Jj3qyMv0LRJAg07/xkBys2KkZAjV4k8LtMZpsExj07NoR1P0BZrvwz1mFVi
9TMKUI0rPhE5CBN5EY/x/lDAexDteaGw1KisWIeJmglY4gmJMpEtb/OwXriP
Z4yeTQR/ElsAF6kD7VjH0EF0+59am0YJs1uW6B1XP3AFYoyZ8y63/ByeCbB8
Wg0Po2qXhzR9LKN7rhtl4jr8Rb+8V5BTJn7EOp/aUyenwIpQ2sXFK64iyzO5
FV0uijecdXTMf99xyD+EyVhqdRuehAlSOcHBy74GzHdwJkHdrZRM4Hlf3zqL
d88ohTTbOo3NZ47Z6253afBLxZyMXQ84e5shcns6KFWTpk13y4+ZOF5vqEJl
goZlK+mRWxRV4NEYnMl5eto6lY1z5lrqygUtOzJKrQymZQX3xPnOi3c87Mn8
LBqMf1/UhpFEV5FPhOyfAFXqI7FdDy+xbBMO2rC9kjUtAbpS50h4oGrZ6cIp
smRfrotXNPnOe42kgZhgq5781GXDkiZp5G7qXlFyAtKlsFEku1Qhpd8r1wEp
zoC8Vq1FYBcCO4j+0fY3SbjKOfAx5llCxkh422twwdRFhnpSMlc6zh+kBTnq
eeF6SjCd3QSwFQwSvwoRq7RtZoB7OS6AeIrsDr6zjDew/ykEey5r0C7lX9Zz
SN9cJp4PUNI3EI/l2TRQ1iW0wFFcNB/jioXJ/71NKr1ON3fN35DWov9XI3Bx
8v7YNIvZZyh/zP3HkgCaCfPFgNHMBhXIcRAuBH/byhJ+Iy2w86Yusvfy9yER
Iw9x0Zhv55gD86syxJf9hz6OvRjLfX75ueHZmO3LBb2nqm86UshBp6Lv4nHD
aF7TJong31/dm6MPFggE0bKcWQyfNAKpSdBw+9ObRD6o52Mo8eS2YXisOmOd
3nlRjZ3wmZIvleY4aptryyPp3EBy4P3tcqBFhFveR9DpiLxaIu30SsVQiX4C
MIunxBTRHX36JiIpv2RM6MY709pF4YPWKVma3JijHwhp8tiPmD8YkFPAjp8E
rjAyRZhhh7rlcAvBEvdldtBa9q2vmpBs9bZpARDkNEi21rjunhqOnhbMFhF4
VLzhWjEDbVh4gBx6M+/YQTszZQ1YC4U5eVWnx3PJ8xE/sH3xa5QS13ia/bK6
sDUSMQI8VXz/RuBLHUfMrbQvW84VK7cW/9P2c6rXCsvj17CedZJzI9sDT5dO
qwRCEU73R+1CWyRyM52NaYIRIsir0Zc9iiKocy3KVpBZLvW/Gx0qpf3LAac8
VHm4IyTIDG7t/rNTwlNDVGq2icyzRYxHp1cXEZRC1gM6TC6xGNU+J3dWpU+K
bm1SMtJov+Pzbsu4e0JLBjLNE3K9Ln8HlWktTRMO6Gvj6UAOPIxrBS4LStWZ
lOnnfJgK4PlfLFm+vhU4W1MVMjncICQyjxz3F8jqmR9MZ8DuNwe3993CUeyT
LhR74mADBuXeT5ZGkrbpS2/T2FlsfWYOHc9MbUYOfe19nX+LW8dAFWJCZLOm
gMQqcTH/rbXzd+6jCjQ7Vj08WwoSKzOvFUdpoquEaNo7g2/vWSNmZK2VPSVm
gKNjIcuBT7Bi8OqlEF8dFXi7TjdbwA/m6QmTuny5WjV+LVuO3r5nkpUPxs0w
AZ8Ut2cPSQGbVQ0rZB/1bG9FHiIhC4AOCsuVGzeQMpR3tqhIHz2oW57H68E7
B07h+sl90/w96DZ/9s0Z7BW0Cn+RzRlAUDwv1jp2I1PJ4LWVgu0sbLT3CbCt
tkuUdX9IUvFVrF9lGtcmFaBx5+/nalDry68On386afJWx8BSxeQ416a38UHd
F4Kg0UdLUMlTeUfdxcIFQxHLg+FzDQL7f1g/0gW43wA+QU31NrjxOvNfQhdo
MuzvsnGHNertcE+q/wLrJIh4v28HtU9/xuFIq3nWCkqO4aVHqzYen32wI4+R
N0jWNTndC9xXrzg2KhHMLkUOZedye08hf6eVKHBG3WsjVzmcLjf8S1cGjFyF
HczE4FC1HkZ7BmWsx0sIkneWrisl1Au5mnQR+LFYPwYz7iWx6j6Xc08vlbXf
2amtu8s/BLzK55ay0a7vyBQY42xjWT4QEJBLtxiYhq8OEP1lQjtINElBSRCx
FEhRsLffpHBDdWDErgB55L3DRMmKcG5VOkfcYZ0xgHAem39zG0v6rNppQoyQ
iMm7gJAfylEhZuynzPPaSC6quR8RGiTlsWCHOhN6pDo8ddRereEVRdGTPIs1
JOOLNjrTouusN1gsnhwxwyfoT4mvSaIj5sgla9vps5T7hwL9YisUAXxXfWJS
ScMRhcL5DpZb5LJKU9bv9BpDJNxmTPlZG2CxbPWILXurFE99LJ0pVcRku1NK
CBnGC1fqtgEbq3LzIOBXePd0TCT1CenPNegJWES5oQO7N12fdNqgATHF+DU4
gbyQw2aioikg1cqOVQP27QzA9sF7KsERDzsM0oJCUc5xGaVS6K8aHmYCiEwZ
MDoiDoF8yNzaW+cvqnUqIgXMTZkp8KtEjs8O3nxLZ8Us9CxpmLXoKwc19kkm
8DAwMCGaxdcHnc+FPzpaMSGMxZwMI9myRkeD2tzHyOyfHbe4vJmWEaLbgNa6
jf1ljOcaNW5yUBA9gKtl+iLUW6VUvYVseabDjwO+V5YLP+kYtmeCO/D8nkVT
h9SbXAHV+dPHrgI1mPs7+RGmaJc2BMb4uxDEsWprU3LaS8qetPPDPq3xFi5l
oubfrHetnpfrkWKTO3sgfTUbg+tY43d8gPSbvuwszw7NoKOSLgJSaZdw2VSe
ug9asv51l1rHE9ehMdvoGDKplg8rwnVnzBgkKjxNmzHPcR2/GQezoMdXhgGF
N8FUzdxiNsYOKcvmbQhBVJUL2Ijs8Vdb27/ZCzrh+2hp9t20H2zKo4R1LZKF
TS+fvf3Qdm1Sp0vHc3YmcQkI4NSkodAEWWNHTfg7jlubD+2KZgCMQAH+1J0+
3Uj2S0l06HA05C7e5kVkrWA1FeUc4fRvdBhyWJGRzckq6exIBh/cUVjU99Yz
K133cPsqGPPfqXs+RNJ+I/5V+pwYbrGITJjMj3o9aVKnQZBzQuhO5DhgPDSV
Tt6indzspp6jl/96y4pducgSRjE5/yoaO1edtcUxtJXNm/UXH1SYFJb/AHtJ
ESB9QB7Cb71HkwVsFdMLeMnL9p7AJPz5wVPv5nXvH59CX+HRtjsCGe45QC34
TfUFEj4uqxAruT6PstaT5c2BGNFEJDD6W9vEKmadgbXeSX9hv8fFxoIJVXoA
msrLnMoIYa3oiNGIL1JzmzDcr/9CfMB0TSXfpyKb0kyCI4pZKIQChKH7qPBq
HghT1y3T0O6ZEPl/8hlx/oMOhxeDgEj4DeP5ENRXdxQ7K5fMTFDWZXHbCI02
W4B78BLaPOMPcgf5SB8KxIWIIUpzM2jwGn+LGIBvKfIDxTozVe/uRFQIw7CL
IllC5QIemtT/UzEQqUlCfheFwfshjFQ8wPeMWZTfzl+HzfQTXSjuewTLV9FM
WKbd7gSC+I4VeB9J6a0BjzNbdSaoP8y5cz5myLe4b6KwEBY7lfkPmLINTfqI
Dj2wTKuopAjBvH0P/f39AbQysoR+2Ff19d8LFOuWhfcCInuEFC8TcR3Aai+z
wIvJH5UVw71o1dLfNx4UQ38H6YET/UIzkuFIzrkil0+M3ECHv+cf6ZRAARrK
ya0z25c53rtGpjmKSyPbn2feTefafNhchaReP/MBmKBxNRqZUWRHkmjNUH09
phnpXoEy6vQEDffDJO3oac3v2EFtzqgEHXblpkAHLr5xajSGxnpyx2roC6rC
IsBCdYNIQzLBhQi7T5Uvvph4qd54nDdX1dH8+oTAXgyXDuh6bpYVBeqERh2e
r5/gg5Y51ehlv9wzRnk4qJCo/xHtJY+B+VxGVFin4ewPvnO0haQZd8LKmvlA
xjM2FyfwMO5MsTPWg/Jxt4vbGdOAM8JDeRJ3viUwbM2U/byIStoW0q4Q7HYg
/mOC+7gvdxgjXEEPYqlb1r8ICRrB1jlC2vF9M3MH0WS37a4AdgmAIY48V4f1
W2qMvrORqx9KmiIvNXvLQDy+gxGeeQCN2Ji/IYLV83IQuMLwvx6JDJnprOR9
EA78y9zz3n+zMVlsidhCUj2rWf/YppohJMvg2m6FAGf5qJeBi1JLOaAKfjNq
WOta4BZLTaSwmXU1bxZGcAPYUofpRU4HdoEsXtvFq0Jp/A8WeYaqZdS+EfQY
FjTGuPtyre1YH7h4M16l+s8JQKuhCdaAjepZS4/Q0zNUs1ff7jJkwoyTX+9v
Xd9ZoAAsouu8K43VbZIAELTSTmBWQ0l3RzSy38AvTJHC81fkrHL2PrNi08l1
VFbSfLCaoj6jkNVnX4dV9p0SEq9DuUzZetwwSlcdoiHVe1esxNJESajztXcE
ZzVkr5WFAwB0Z7V9r6bLnfWwcktkO6z7K2Dxuhj/Nyg25OkP2vC+IS4/TaCM
r6tdi2fgZu48BKlMMI5WADzR1ltJgYNAMoJFviN8w0qgDOypJy0cdAs6GfM0
uCPFW6HfDz2C0tdg7Tcp+wtMJS4PR9Lsi3NyfNj9m6KwN7UjKnKF7OcsFI9n
gtCS2XRw8rbLZN9oTJUd/ibtRecOQHNAHY0rFZFCurCXW4+8XpD8CPj6ZaD3
IRhehmxSEHJrU0z07azq2ONHvK1Vk0RGqSuosR3VPD2EPb3uloKBlZqWbAVr
5LEsQmfjX+CWUvi6GCYAXNmYNrf20SOfjyh7PBMSsdA5H4lQgBvrxSicjp3U
O0Tmh4PbhHMMaqU4HtT51ch1Tykw71/JTZxC2AZZqISbqYN7cd8s6UVVOf/v
tCgaX5TLTGAzdPBqY32kgtQVlKtmySb2iqS/QNNSEEbXzMtAMuBNj91veooR
PKn75jdHkxZP2Fqa+j6p/wUGLgmkhVVX6n6L0bDj5RGQC31KQxXCgGURe5Ai
NxJ+6x4tOLiXfnKrwAJgFBT2hYoVo393KyvgLQWJrFndo8Ckt1fbeqzsqKqV
hiO91qm2fvGyuEfKqpamWu3AIoIAYv/lCBnHikI0UAAahCX5m0HbPvYPZsw3
pPjS6v+EcSJgSknx6/jAV8vQIbSrjbIIKK/ntGCXA2TTf8WWz3OzK/3EcCIZ
JgUY+lWcJOXpr43vDeuFfUWh8upNwZGqnrZmN1/U7bNyX8j3NsdL8tDtEwKQ
MBXgt1K73OtSjbv8W2YzbKTEvztWg3PnSOSPF8yQTKlJah0FTKx7yQ3oolmO
7CODt15jA6njb0fX2xpkUgc6pRFuFkfYolhGmKYZcTPwSrpZjipGhH8uN3yl
ouKMabtzxdmrcqu/x5v5QCYbm8DyM8TDbV5HodewYmsR1VqenPobbwHLs9Mc
vxQfBAfGLOqCNG3vj1EJKq16tYeY4rqxuyT2YjOyScC6HFmwoMJbaoEkOuyX
CfSqKZ44ncHon4cX689sEQsKBR2vQjFztm3Te+V8qqSuMnrULHPaor5T0RC4
3YBzO2lMTvRYbKY6kwlnriTDAQBpUdkJzEly7VOv+RpuUqylClfrr99T1YC5
W7xh2uLeNPveW8CB+6N0F1C/CSkRcyRGKq5waaSt/Eh0ai5SS1zMInryQ8h4
p3zxFuMVzGdSocUqLX+xg6rL9ww+7p4yPdXrkr81IhrLmsh2L2XYmuqoJMhK
vUyTCjVg2mCd6rVIsh97q3V7e/0IdxhtEtyqxUqZU3v2R2ScdSjGXP60Bp3j
JNhdWejDtQRlKyQFnn6M4t5K9CLmEfX4oRt70KMceVLx29a69kYrd8hdUwr/
63zC8cgBbM1PMePwURkk2BoANBwVQT/87X5vrPMbM+fF/a1fawngd4+LPTP1
matv3WpojCB6L4i/OJiGCTB6p0j+5BmAndlNYADR1O6yjt7hpRRx+r7V9XOx
UpteINu4V5oHgzWebDiIHn9dbKXDL44wu04UtRCbAvmJk3Xj4mvDY1e3ZMRT
6vV3icgkmqKVHH/lIQt4F7S7uT22lW5i+ePaI56KGDH0vBoIcD1jcz9k1qSP
7ANRFAKTVPczA4qtC6uaq3fjANPjRSuwanQP59aF8+FgxLtVpCUeZX22ksge
hdzId3XkJSVru2QW/aVGghFIYO4CMrNg3ueT1qQPOag4EyckrK2I+VyZlBxY
7W4kY77qhxpjMjEdKV2lN1N5Vft7mz/F6E+vC9FBZ4VuFBGLJ3l7oFaalXZp
oJXgqGFZrk3PEmKXRXjAWDDfbXWkOc64+QHTnrS2rVlOG2nDLTu26t0zKTiC
M4u9Gx6GAupjUijELmkPBhwfzzLR/Gd9KobJWoWR2c4Qvtm14oAvOk9IJJB+
8wOF46KBtaYdZaEhkcEwOEx+Tto9ZP0XpM7piecnvKhhWz0hjFo0QNzYFqgo
2pQkwa22PKIrQ6BYdVkGpusyeDDwE/rDEo7iwya6OHq68w7vOR9Svx+zhM/2
vY12JE+wo2aXZ9LD+p0A/rihFFheE4NubMPtM5J36W6f0ko83f8X8BDPr1f0
Gr6HWOT/B4wgJjZghDFUy+LlDMfD9mCo36klUYnyo4bw88PCwkkLPXyKlLmh
1db/YU3p9zBXXN99tEyNx3YNO7frGxeCOOl+yM0fqhnku8JpLXVItR3L0/Er
kPZpyHuifNWM0pxN2XCvPCqk5ElbUG4q+d6EIfSNk/190na0M6HhjSBgbnr7
TjopMqGxfS2kstzKljzBAHxa/smQ4Hk+UoCuH4yVC1AEARaWq3Eknv2MVpOn
u52o+IVjD70E0s1Mw3tE25yugPjSMY6wKwIE40fkfpNyg0+g2LBnRWlmJ3pZ
4OA4mKMIC/mWAyXDQPei+1VC+PSbQ0oQ8E7PpOUfWaI35Qid6ypeZF2N1Eia
J6NQShiqBLgErjQeDvJdUlJBDEO3U7/J2tQgCgsg3B1WbbV9oIjX4Xibi28M
QVQF8HDEJsI9qBpILJxnQJ43nvF748eWEYgQy5CYQpag1rdKRgdtLTmz6u4l
HSguDi1EHYlnzRGwtPHHSvizwq0Or5n0CIL+ofzhXR5cuaUfDJikPlyopg7g
IcdeUGRJD+LUSKwjxSicgT5umLKIVLDbu3h8WX2vYpRfg/Rp55J3cb3ee2fj
LaUWEFW1TTV6K+UO6MXv1G4Mhlg1BgOL0aBQ5+LQXyHte4+EHyqeMQZ0Bi6A
eJt4oYs0ZEp8yFkSe9zXW4ak0qR+YbSV7qSppmOalx0cg7ytai+DzJ7DKOmG
ldtHTpZEP/GKrdcBuO5dVQNl4CWmlQgn4Qpz2/KtwaqET5b7Y76Z0FstWt1B
OggtZOrPTcW8ULTVo2l8T8azdulFFdfaKm6czLY8Nc/2cnzHbuAnr4rTgXVW
glyfgPW8+NarbXJQ/O0yNbWrm7qS6w42/azAkA/aLIYyt0ojIFRUkCMMklce
LZbLgMzNA0KT0QcDASebGbzpfGqR34VASqFGfZUOyknEBxVXU59RehrOhqDW
a8Kd1FQ6bSPwZUy7kIMKwDSK9FtVf10DFu+KrLn5HNboUJfGo0GuxfkSPccz
/HKS29nAO4Aa9s3JTYkGnRlX1a5pfcd+1UxxCTHqAHj2uPgoo+kzk0sCCJ8v
YIT/P/Rw5u+qGq+Adl7CNq0hQblWN250afGOf2Z1gliphqf3SQECC45lUM5T
zLkEw4iuqt3BHHa9hophqtmdBtYxdUY8A23/COELP9xtB3wU+kwgROjp04AA
XfZyRhfjA1m9FSKRbrzWQL9lI/fnxtKKam+YkbzHpydgHD/M68n/P6zbeigI
WGncu/4gi6T05HOZnKU1CwBIPtt6clB9q8hUwHVb8QdrqAKXXr69+ZK9Zz8Z
Gg6EK1PQwEvyM7hjpOHcoJ4xt+jvCM+ljKVnkuaXFGiFiISggPWESiz0ckLt
QTIkKDjsEsSiuiSPzpQcrqquRxf7xnPqwwQYN78IO3J+EfYfc+962plscc1R
twE3ssCl9fl1/3MER4yx8748wB2aoioz1DviuMOmtqr//FJSmtj7CBqDJYQL
FXXIeAZLwI78oGZpaRdOE+JoLgpiUJDaRqf3xbEPtWdjt6Y1GtD6DJA6rwCP
Pr2LSkQgcZlb3ms+qRET1agiY5QcAJ/SXtik9BCPjA4F1MA1P7EH2wXPajRh
lCGMvRTi/SkPBQAu749yNBl0z4HxfZ+NKreO1W6z70ygyc3oSuy8yuBJb5iL
9QWgW/m5UDmIZBmKMwjHR56PUJda4echWJWe+C5oT9Wgygs6MH2K1Q9ZAEFc
x3QJ2hVjib07/jcqC3I8AsVKyGs1k8sXCThPvPlkGQTFjzBkC7uScZ2eGf/i
Q68bJr7rqDXeJo5xPbKydfzdHzDdxRwD28WJ8YdGmB6qC/YA3SxI8jAI+x/+
4TQbmrWwtRT5Yce98RnwpRvGV3oBFdE8KMVyRF3s4B6LYME4Odi35FeVkima
u+qZa0xMoV+Ceej+tPqho4uky7UkX9J22hfh5ddLDgn/0zm/SCai3kUrhD0K
gKR29kuNIHDzElgkyOYy0I33YOJG/8F27d/4bVd+XLGKjA2I6USC+Ie0JUoL
QK9zzwMAEnlWIftposVir3UjOxAt87XgqysJjjM7js9CLccrR2JfV46omSvQ
HxAX/K9ZxoJTNmOLWQXrtygK/XmfhgcWn0ie7kcXkS6zXWF+gKjxcI8EDwRw
UI2zNfhrQU1Dmn8DpWtKmBLN3sFA4W50BVNJHgFI/jfVaMN4FcxwZcOLpTGZ
soOfXj3VdcgXomXdhTWL6/20AUpMm6ktBiwkq9aAorFIa2BrFsSxau1GeFGz
Sh7PZATGd3zsaRSr83gFrwZCuDgN7PTh+VghHRKF96Q6BQ2xtsLf1JpJlwhT
5xA3Z9coLKUX4HqWJCxIyN0CdWBHnSDJt+lR2c3ATpUSmw2sYYkek9j08j3d
yKoPnImsf3qVXQ/44bqqWSFSb4ymPrba+0lZ5na0MN0BUnMzOvdDryg26khw
ufNKXarq+jCqeTRt+0IdNjs3OtmAJIThrNw5cVaOdKDEufi0qn5SL8iW7+PT
CE791jtmWxqEZqIdRAExp2QGy4v6sQMtCUxXyBQaIiylOOfnHyuMURZ4yyOJ
zxLthcebzz5t5gWIadpVrLeanZB56OT04x48TsyM9dP4QlpADP5r1n4GFUQ4
4VGDQ+lO/L4HcrK2P0swka5vS2MCQR+YvZHCxYrpRUsuIhsIKLhWtnl+fOwL
79NZQwlCqpQXMFow3aCZpgVi7ujyeF0wfnCltBLLvwX9EQcSITb2Nt4KcoHn
EyZcAUl+gGxmfu1X90/tBg4QI4nobjxEwO6a+8s82uXl+JqR2f5856ooS/1S
Bwo71IPkQeaAhF4Fjrp0MMA8B//PvFQYnL3C/1cgJWPY1wGKPEqjYjty+XGn
Y/+4zB7b5arENU9vpbUR4gbpKucO3esXS/rntvHef4ZNwSfbudwJ14OWzZp0
hP7ziFvxJqxeHlBzPQR/BBRJq0k80jhpR8wXaRJUy3PSLyL9FhobV0BzAUke
cTdsdIZ+8oOz1uGKBsyGS/8a9fUa8/v/249+8jmCAdHQ6Pa3uSnPOnZbf9C/
5yO4E9RpGScN1CS4QFAjxcfxKLwoPwlWwtxs6H6qixOWy8sZUjGK1irnSjwX
Y/5FOw6hGqsswoavlSDv1d0fMv11r62LiVKw1t+AQ+c4r5zna4BvYf4P8aHx
CYwKfvCFPmkLZSSfHrB5+bmlaVC0CBq5Fr7lfPs0LKEfdPNh6h0jXja4TGN1
M284JrLRVXx2E04SR9gdkG+8KZ+WBb7lUjF8sBYjRSX2/pt1aAcTjWMdodQq
N6CZKd4ouzslc+r4rjoM71yPQ4x5/AXLixhky1jQb1eU6PrWEYxN9LLXLTOC
cqTv1dxe4CIj671B8jzez7b32tWQRccBj1L93BQd0h17kdsrAERecMSc4+5K
JQN/iiWb0UT8JhotSRdR3q64WlcxBP0NkCeQzEBAIVq+a7JMUHboDiqXWoEP
ln6bE9YMwACokZNL4QHKjnGDobRzc07cgy6eoyERn6WKmwkt05MLZYhwAv2f
gJc0SgIkwBSTWC8+gvBy5seVTiZoLVHUeBMFcJUPvDj4Al8CzdHOLeT7EtHP
G5oTI+ddXNynh+nFsXJZD6GfkM0lYsgqDkI46/GS03FQml+O04BSoGpk/sRT
7ciomJL53cXaO5PtiH282eWFGjr0M92JIsNjKTsA3ONbRLFb7iwT3k4/jdC5
Q2rW9JeN7hl4vXxPy/myGbiNTXEyH6pQD2Bhg2tApcAKqpotgktN9RBfBTx4
CcsGmDmaS7g7wutHVdZTgIUJlMnUzHkQfkMOGOQIMsJHmVRX4aLhkH7bxF1S
z4cLWlmXGdCpxvrkYj2wzTKJurfIB3cDUG9nAPTbxJLd39Sa+5ov3NvO9Lkf
yTzJW1VIBPlLtEz0SlxLZEF/+LKRKCxKu1mZ+KXJ48wrTBBp3iFixMPTnlUu
3zULKB6htRXsgoAx7QOXptP2gz2j1lS1PH3UibKZ5/nK6wVg/rfIVlkufqvg
Asz/gxLIwYwxVLHrD52AQYumkH3ooE/3Hp97FA0nKNcFw29SOIZz3BXzpQ9T
3KJpREq0JH/50g7BU69Ysu2jQYYUWrLOe9RSHXxD2SRxkTD+bEmppcuX7O9X
flMckXJshcPb+FQfzJ7qbiiQ1/5Q0ztRBHHSVpVudjz+deDa6QDhHDcudaNt
qaIX2DU1R/JurzGUjpHjExTaobuKFL+266DCi2Em7Zj7yhyJjwFDCSf8b3h6
1Ic7A56bm09dvya7TZ7AbeIiRPvBBznLVXZn8OSUA4gZT5PyP+N/dfO6hWhN
27FFJ7wk9aiwvD8Y9uRUQLS1uhlQoeRAa+mfjCPCCrLOpJpZefeoXchJyMW0
GtsYjjeKjtEKTe6IXgMsmv6ctcV9+Stvba5sZJ6TbbPtmjgKx3+k6kgMMTtI
Q0tfiWSzcouXG8lMcIaWKFVzqUYec0fN06rw6YEMLV2IdtktZLWfj9wvgnLl
Axc8FKMHoIt7Cm7gWFTEmUWs2cXYkJRr0S0hXz5XzRBGhNrttNRO1y/XRorG
sE3ptcrZT2rTFRVf+Wvw+Axa6wp8Rrl3ECsdQzLjkbihYwP+dfr+QZCY+AUV
9wx+G+6unR7WTf6v6bCOMBBtliU3Wr4oWVSc+zX7ryNVD0mGgImnpDXdc3q8
aOm4G6dPlMc/zX9zRJ2iimdfQ0liFNTmghq+PkGuu5gaoxPnhrHicQwBQTB7
FJ5axm37JaYAryYkv9neY1Vk37QxES5zwLMmsiP6AjTzXpml2z7xS5xeH+km
cUb+6O6xHZ8hQo+DIlpgv2C2Zt08W6heJXYG/3g3TQexCA/T7CP92UKtQJte
5rKfX3dEptG/ThF8FkBduq4/HZKN9KwRQJ9TyprAH5O3FxW57myhZ5HyrDJd
5GPDYxQiW++5oENkLT6I2y9tQOLsFlgoUOTRTLJehmUkOEdmlT8PDhGBgbv9
dG5C4mi5Nj4E6UepTl4icf9oP0rWtpOH0cKTXqAlJyTnM1AA5O0simImr/u8
NYDoBdsDgrs4+cfVwPJLrrPrJDmLp2ftLNAkt5FyDL5xmlpsNq2k0osMwbsd
WTtuilVlNsRBq3PrGfIlyOifvsGZSAnU6jqLcuFaz2MEa2qpSBnq5NXhklrj
5+2jEy5ooe9nK/NQV2tYwOr3GM1z3JD0Pn6BDzHbMa88q0HUyuIuA/vUvk7z
ka1nsYwfVKO7CVAR9PiaT74N1irGb5FeRIbc8CWuEpHY+oM9GK6YXsEkA1yR
Sxo4GIKOwCM6XWjDKX0W8WCfVzbd2W+QhDTyDP+z9E8g23G5Zuh4SjTr39bf
i0BN3bs6FClXs73hAbzAWnCHc4QdHzc9rTGQKZtdhq93v3pVOQjf4aSnR2eQ
FPUROmngztb2Y1q1gCWk5mQW9OM9Sy7uLbM1vB3MVGgX9esMEYOkb/n5yeUA
RLdmCos3Jnbxe/gRrAkxLGuDYwO99JqdFFLC4iSYLP6EP9dRtDRDOW+g13w8
SIRA/mnMdbQv7IYMwj4d64dgA5PGTelxuAWWds5CyyCURKfVGgyasmTho28P
XY/pAjQlTAjqYW05fpxB2iXBvhJz6rOjeztA9ZxfRU/CL+z/oef3d9hH7yg/
NCT5RgtJAY8kmQObsyr9mVTohQTv4Qr2DPmut5rdk8+BkduR+YsN0QYQ6PIb
b2j6VE/j7/JZ4FwBNtnACaRZZI2kBFNav6GmT1uJeef4E8LQQVm6Xuav1vWf
NRenf5WFqVYletvRIUhv2IB2VVzEzEK79mFhythZZv6dE9gLhZqAhztcdoUr
p+RCXlKyQYnkhcg+hTbcW8mFYkNiCXXdc0/bbQafqzQD06U5ABazz2tGCUbI
tWEQjmPWBlAr6U7qjrrpt1ZmIZ25ODG6u6TQDiBjpB3NvUgt9fhhiYmlDmAg
yjAbr/VA9NA10QRdxWQPcjwP/yWXBO2wxb5jjZExRBVGuzI3YvgYky9scjNf
3yeMHqUB7aoUIupwmGJYDmZYlzBX3UW0iNzzj2+T9GCtNJI9SUOH3S7/IKrM
/9LEM8BJTGUZ4TaDAk3bjJjgRVEez6kXxYo8PGdkMMRFtjhCs38hQJ0mwBFo
MUH1692VFwGSeOzRjBPLMa6FnbdLQgSDXc/hQfnQoPa5gDc29egcMMhZEbkv
DNaUdY0bk3w84fJufEFNlgDa+4ssvUVQlZOM4fU4D0Wtmee4mYKiJ9SxDz5b
x2g0oOkYUZsPKEHHOIvWxBkJTVfhv0JJaNZbiLFUFOZVOHiHK8Iy2EbxO8Jf
WW/WGz/4hdyWCeFbQwNJFk9ZwlS01oSzV/Gfr+CYqEza2CPIN5gNF/7Lrf8N
65ve9e/nee5KxHzx7t9D+YNNoHiKWqtDvNbwketNtnlXW7zNZJoH5xzetUPl
QxyvbirSliQuQyaM+CUv33DfgnWWjSvtnigPnDbMIKsq0B9Q7XuBu3zrBiNU
H+4lr1b+Ue7fsD3WbSmJt/aHfVyF8jBw1SOxw+jXPRThl5pXiCpRtOCf5+bt
07t/qEfucvnrvClg8YS7aUsWS0nCueo20GUORcYC3R54nZmhl8qJGGxsqEXA
eLJqEYHKcSMseZURf42fpDIebyAXW11LUQqoqgu+Jf6a24Nt2R0tl+462RXx
oDizcQ9Xl+8pyDrf9fSrrBpYu/xosxsWpsNBv3h9WusPXys5Ct6lXj7f62cN
5n5KoSSdV55hJ8UFnzNHQuYbAE693rFoCCIQzInEsbAXpreXpLdD2UK03T9Q
AZ0970byn3AFqGvUlXFYMBJqc2B7BB2ukVyxqyhoRu66xU1aiNZxL8aLyLz5
3ZwDqAZuYhCQhJ8Zw6guTomS0V3iO/PSd3x6a40iw/L/DlFtMea14fIWIXwB
1KqDj3BgQQECiCR/d9UhESotMx08K5bKe5HZd+/AAb2vix17cTcuxGnyUZ5l
2q5Qvyu3WrUjvZrjRpw5LSgVCz9QI0rJxYExDE2okvJcxiiEUUOPi6VCw69k
Qp5E+CJdJQU6PT27rCCFmIm/CtQFUN2697F49VIAgJckvhtfiCwMvS97APM7
4FpCucUNO+OGJZS9BadfrI4w6g1TlETenRnVC9q6mD7XzksxiJTmOo3w4xNf
ZS3vQtvNy8HuwP7am7e/TL8hb7fbVOckLlenYVVPpT8gTtWQELPsNoqFZsS/
qNly9W19jRZusvweJkA8UB8hoZe71Cx2bl5iv91uDYKZYhYa78iYpCLH2Zt2
bNeuoDr79KCCoiS64+271cVVQbw7oNZs3R1sq7aDxcPYUlu/NCNOiMM+S9TB
VbFWT/PsTt+gVkkQaI++uKHaO4teB+7q4l7wFh+FhIeIa3jDEUFLB4CM1om+
/fM9NW7yLGz+jXZ/lENqtK/Ksmc06GildA/NTTRvtF6n+PIc63/A3vWdejuU
ToicGKKHmprx+hOy784GOWGe2b81kUurLTehPrnFdCpAi7UIc1pvBSoSGhuY
drNTNuQHBtHhvyZ+UVx5etum7qnzCErxQpNO/0JqF7oHBAqMCxok74u/85Up
CX++XrJD0h1Rjq81QEC+PAvKGA21RjjORWArerHOJyD4333X+W8NHjFYRv0c
MuG4pvZAkRXhm1Ky5vTgqPsdFF2lit7sqlFY/EJBXDpSVu2AKKE6CUBm+TTJ
ZUyL1irzHN2HpSoDaPkJwkcq3mcRRCZbkkdE4QKWJibt1+Gh99msL63qXFmj
HRnV6f9MHC5oU6RZbXLeJGkcW0Rccp3dvLPDYfFIqMipSVJRrn9apuQtvfAa
7FlnlfhKuE8nagIyRjJXpBq6ETaVtn0ZuT3Ery85ROg1mQhLESePes8Uea5w
86RhX5kOydWophl/zm+CLrvrAsfyAKKOl+vH4bGUqPff3Jt90fAc9/WCdd1k
8BJWRyo6uBMZCEhtgmUlm73Vp/OGZkrenYlf1ugSJ9na+8EHtv4Kcf2svGqD
xcRYMkvTASMcO0JlMkGrgPqdvDt54wUxQSpTL0230Fv0Kr16ia+Tyr3Vbjmh
+ONyfr6ECykDK1Ghgfv0Ahzwq2Kx4OPyna62iRUUxnY2+OJPSjVC3xm9KIFz
TdVUCAoBbqH9ixyOEbW6/ceWPDIMWPv/iYiCnd5DFqQHtwL94FXLQ/CQzmra
xscLVkk3sp2XRGTpVSW+dg7HG+LY1v0RBmw9Wx3J3maZC8zSAI3LhXYvRr2g
ySt0DaunxUzbCFYJKktX4eTFXN7ujXq2abxFvoeEBDAAH9UHmaeGr1Mm72R3
5BqGJPD+4mpAiCdsnW7GSm+y622Rieh1dqXtg351XEiTDXhy6rACYkQfg8gK
sBz6vRbDsunLVJYKFvbJW/cmTppLM90z08Dhq5c24DdwahfOWjhJwb4zKWnd
/MAYsor964jVkQI3AM4HHrQnZioFJD58EtdYiDYtbImveLdPaO6UaZTYYvIH
+y4nxlp6JTyMMStmmMGl3LxnZqpSetcSAYuKv3up/LVjT57TJG+YmB0Y617l
/sRA0pPkt79/y+s4DKkYyxxrbAGVjr2XObwdzLD445UZk/90Rk8MqvbOgT0t
fXKugfNPMzZUwZIkHjYqJ5oc7cXWZtcR5x1hDlgI+RUmh504HhI7o9x1BILp
U2kASsL/jvvIlkI4HpxRyc6itLiqSO0iGgOHtOR7wPSxiPdAv4qrlnRUT9Rm
gpBk4itkK4CWrrQiu7iLfyJ94NyzLZP5OKqBH5yC6AtGaDE9MRO2MyVgq5u/
KMUR2Lr+DF91m4l8hFC0tKX906qWzr/UuYTi9G1+y/WdD15Fr8UswPQqJxRP
HnzxaZ1jpDPmrQCK2MXKjrWIR8VyISULFofzx29l0ECI+OAUN/Y6OPtEIi+3
uPcSeJjTPlSgzg5X1W7ssPxwY37RLBT8dsg8w3gh3nDEueslcUXw5nB4cskc
SZIW8jK3JYEu6+2t8gYYTe5gg+lWkxLFeCba1D6Wvrq4Qk5EJW53WiHqxug1
6dm6zb3+7joZChbIU8PwuxBBjgxIbkOsjfkElHWV1B/P5aAnDn9QBZ+MM5HQ
RwyzAdVhBVvF8SnEqmfGDSjFEMC34M4AFEUzhbURN1u1bDCJrBjVOljzOBbF
Ccw9RSJzz9H37MVss+DPJEBJegdKBQ2QgaONB7+UU20I+ABKzfzhmeCkttap
jvwppf0pDO4cVN+6/vi5wAwfPjfNkp5HhoKqIUuLlCJ43uZhIZ0JC+LQS+CL
7RmHUjjE2JV/EA6LoChO/Ub1IOwP+ZFjfWZjQCqW00J/UYky+1qAeV7kHkxM
+1ZHyDcU6lkmbmrnC5guf09tsK5wYzkmON0wZYhikYA6jsrWSLD6cfZOS25l
uTmYv8nSHXDDVolq0eYvcQ2WZrI4+w/szig/yIu7Ft/mLuiGi+Rd2PmpqR49
WdFfyjSEBBi1TK2Jp1X6cnBkkHBiT193C9FKRqoaa02UxZWWvqphHlPuo+j0
BKd6EKGj7EqZL7Tr8i2zG+ETVYPQms+YEDZGv7SYEaRA/x0eZUX9lrjeqiYk
89N9RzwLehA/NPUee9S4KWMYH6N1kpHda7QVNtnIUQTExopAmg48xV5fBBkP
SMElK8gkhNd5mNcY8kbqKewq9vqNnNKpQ2PFv/ChT+IN9pZlGThkOTvN0piX
c8WTzNVM4cfkbZ4eSHvLRfcm9jWOgWpyV6t3cyT/L9nGLho0yogQ9q2fBSeo
lCE791Xq4P+Pj2KUZZ8+lNkwC1A5owO2nrcmdvrScPUx69zKGki6OPf53oKU
h8AAvDTq2Tklv+XC8iNeMqHQINUHwi/Qwkxv3INmE4od9iS6ZQ4vKI8N+STr
ascWzq5YAUdJC2/hb0i7C1l//gxTuWsfzJSU7XsP/G6/WMgVy1o0aBhrm3kL
wNH0HocXSoaEAo1IXffLr3vIGm41EuhHqExUp8DNXaU3BCQsUKWwPcUrzSQC
rLLUlWxnj6TzpfjEDvoVS3kbnMdm+UijOuQZiN91XNjaxb0Xf0sl60goiBXo
vbY0ZfgTBuzjQ1oaRkZw3FRtSOD2n13A6CIold0sqQmvqWqUaYXDelxI95zI
hWQha+SoMDTNOeTacMOM/MUvBiyO29rtgDJ4WQm5s5NRiFOJNpDwOZbcJWiY
ROelO42oOMP7ErBNV/ytCENzikH+umr60m9FBRA8VcJzb+tKDqTC6EM3cv3Y
jK40Wuf8HoCk4m1LPS1kWOYyRedk4T8Ek+/zqrsh2Qha783QKLkYQ2HuwqBO
pGz0enV4rJcAZd1gVIaQeJXxkFy/1oA7BcxOu4tPq7fUNcAnqVv83lKiFpn7
FxD7wsbtC3RirPVTJfl8Se6DZz9s3zzBDLwcbVxIz9HmuQ0p5e4QcqyOcR4b
4NsMaF5hkuZg0nZuRAMRV5fvUzlB0ZwyVk4/JKZ8qxGBzQ3p7rxKc8nDzR+w
woky9YIXU+WXxB+bq27xMx2Z73OIHI1tGzB/JNoPlstmhUp3lJetKx6hv3eD
weh2lycTHFrsRIlznQuC0je8Su1LUWLHQx65ZE0sovsTF5JO7HJjDsYOISrC
ELbRsLgBY+6K4kb+16u4nKZVaQZAKktE2CQLbOA5brso3U/kcFuyS9JEx91a
Ca4oEFb/h8AEds2hE3u+ESgYY0Njd+qarg5qJGnsL/BrRHASHEDBLK+0K+K9
8dss5kuQ4zZJFRw/p1Wku5ulAUgCuUXKa34knXZT7mNOZvcGKderkoLaoSAa
xDTfDeGnGHbHTxbbnzUSp7oLW21zquL17HOirBVSuz/3mfuguyDsnF770Ti4
4E58cNstg2EyV6Sr+SfmHZkw20ZSRU08jOw48sNHaa5w1CuLKsWIYCMJ3qRL
lh/4ou3PfZ/bf8vPnSFgtCjdev/Oibzt+QE1CVj1B0HowfV5zsZlck/EVuFC
PQBZzHvxpeT2DSNELsnedH+FQJy5Lt0q59RJyJyO35bngzBW/ZjrrbJIxFBf
J+mExQW5dNFwintZx0OcDV9H/2otWDrADv58f2+ejn+cxR45z9nz7DsAY1Zv
80yrNfwYkFwejyvfxqnv521waRn8XlBDZGRz9ttmGHfRVL4Hz3d42WdQG5nc
mnhCVpAq/RS3yASM8EbpeVzYv/cQuVSserz12MnUWyWqqOCuZoapg7iUSNcV
7SVEXAQ6Sb2FX0S4tlOR4C+tpJgO8kdaIyVsxkfzc5jg+NHWewZFkxgmVCod
bE9n3gOTAeP/ZP9FUTYChVhlDrzj3tXBtRSsHeKTI4KIqEdKF7avq4D+oAvJ
iEKYyt/PBYqya1al6zhfmLIhJ+42/B9apgAGVf/4F5p61oqhneR20wfTpHgp
y9Z0NzM/nPbGsq9CwVREMLa8n0r0b8LLIrcncQQfIIAM2rtNy62r3snOAoI4
Off5kCo2OjDPBtA2nDNAthzLaP7zI+OdQ0A9/R4lRNOTTGBayVOizlHP/cys
9/N3kFeL90ZH5qJ/fcb1OBJIwEVMbXPkQd7HcwJm2xTcuz/CIKkACkN+wtE8
E2HfLLSdrgB/AXhlUsyK6E0lFWuZ4vey7X93k7VYUcQBAp8QFJYIkRGVh+d5
hBm2upq38z/OEFIu4RfgbPJ0D1XVPmIjnAe8KAiy7rF0VgsCnf/5DwoeUgLN
f23E3odBMIXOX4inTN+mDXORHcbdBt3teihsYQcO+OBT18doNGfa/dWmSd7e
BJmNl/d1tohZiErl5RxpyWckRCheY0oxxfUcNumM59VzrVI4hhj59dUh9464
ifrcmCNuRnP/r1OxBT5zLsI9pfwpY/jfSfKuUcOu+HbBwxKSJVdL1P44kzCg
TyKgKqnMf8r+n2ppLZvivR6KhdM/wbfYcuA2O74kF0ZndITTreCl4N6vQWXG
niNuch943PHUmxxT1OrRJNHW7upr6vag9fbl5SNkFBudGsfWQxelKngYhbxi
P1M/Fqmf7iWXEBBSPtYRQkTPqxcoViqWv8NQgagmrp0XSuetvRReKrRSWLYz
FpZSKt3jPLf7BVOO6D1qCZDEWXsvaK1j1MnbuibuQW+RujHlAC8g6Lv8mdz2
0gccBxyBnn8jDMssmkqtDVyYCgliiDG5bnP4SQHA4XMjWtNFSkPYXAYLh6uv
BD+d5MpsjEkSIxQgudRvbRp17YJ7sSG+sDMdeJ8Py1Nrud5ZPg+cquFsvcS7
9lfSiGdXhbGF3chnOmMimk+qLNv7x6f46zhIIYrHPmwggE/eQ6RTYpG03B+a
mkI3hvVi7kMqeaxLVbe7Oys7X09TslrmZF+XjOTopWZc4bHKay7c59EN7r5F
0jQ/UmUCq8xKAHrfhwfr0H4fl8dpSebvJb1EpJqGUySBjzVwxbxsqabcro5D
rc30lwQ7YkPaGHkQlBYgP4F/RHu7Zy3xkLdhE00NndXeMUwtkrGgtuK6aRHi
kOTA3RzDkJ8hPUUaIs/coP337H8sBfMB8erjfbTHljOozJ3H6pWXOZI43bL0
TRyt821BBlqPcF7vo+eqMLRFxBfBJKoWzL8b6ZmEgN9Js5D5vHX6syXoKGqv
oa+9INHdgqKUFZJZt/emC3TciVuc+akcx7p1l5lRM9ok3kdE3nzNy16wguC7
fXELQnfM6omISkhimCoUIMEzZETab7iInekmDcFlonLdfZpRkTwsWzuolGiz
FfLn+6/cs2TYFWdTPci+XX/frnJdmY7/Dot6iXbcF/kCd+eGzIQvAYHiw0Mj
i5eTHfo9M+pmwxPKA7n6pgENytX21fVaFz16j8GvzLk23zcBjHjZk3TybBGg
cUVYtpoKKwamxDTEVEK839y0TH9ONNtdDGDeZvAKQKLUDYFP1Y5CPTho3U3U
VZ2fkxg608365ZpkPCEXol5cWztG5oS6nkdWpfhdkSZMd6BlytUgSz0iW7ew
YB2aNXIuZjEz6RZZAr2e7BuJ9ETYu4jPfg7+mo+vsigftlBnqQhiXpGY4LiL
fH86ORogs8WyUVt/BPLavxUN3Wthh+kj/WrNiQnzX1JuPxgw+oGkPgE9cN1L
HkyXGDvBUQwKU6uTE/kDAhCgu3FkOTzJyvU5fO7gn2NykN6osVt+ZAoqLqXG
3DxlUWcaQjLH0rU8anPI+6Ge3LnEP9gTGzbJp/Wt3Cn/yRwQmTi2hBJ/s6mp
/IQmxtDHNVLY9FKMan/JpE8we3bYutp2libo7g7WU+odzvYogs6GOJTXMrIJ
gjSl14/6eLJEGWWaUSOBiU2Ylvw8vrczTpagi6I6OSulda5LzINyO1MZ2Dsa
Vxe8myGRiSVFII4Xv1DRXRo/HBTl79jlnV22wWEgpmOl1FCVoTo7RBVBc64X
U6kSbKloWenhZog6oAOW6J5VpQ041gfdJJEHWV+tREzhY0Y2KLSIEdG3F1tR
gIgrYWBOBcoJf1YBK/+Kx3Zs3kc247GHv8yuvMrO9GeOiwo6MrmO9n3qhHz7
yyoGXFVjKCY7N1uzplrNCaK62y1g9t/nX61MMzXfx92nXiXtX5JfXpr/89xj
1XObVcI2Ta32f3QDCckzhIZXYz1Q5ebr03PVIe4yCtwWyhl2qGeMp9BVhC0z
LqRInP6TOWCSyWGwzCw9uZSOMkJurVxS8NP9gr67Rr/s9Fz4097lOQnhbHzJ
KECRkQp6OZufTe1ClOPiuZMJeHPWzzRJWMXQW2rUMQdIfwMzGYKMcYYQ9c0i
bQH8Hcy29P16a4yiWGWxFUVSKz3nWqpvbWxxYFmqbr50DDA1J8tTS9pHWFfM
sqKVBWpEWdBOqgRrw/fqfzUJYEo5YWAVwagGZ8WA7ixKOaYJtQEwaZHdkaBf
sF0LcXLXXgIvDfqnVNGcxWTbi5jmSxERb3iy65zgdMZ+qX9vbhH5i/Le907t
7tAIzj+XSiwbjxsfpaMIpaqPhL8bk58q9ER81JpdSzn7WpwdR9KQZfnoW9mL
hk4d9YMQlqQb90lC5a1fPYe5+Y83YfhTm9eEQihDf64FAGvQDWKw61WPMebS
OVSCcudor+rRODoqflhSgZlh16qO2fz9vEIt6czX3TmuU4sv3NjBwLl9rik1
SSojaRGhx/jswleYhmExp6d1pHcl3sUj8urM5RZlSUUcIM4UODTrwXer+VZx
dE037wqCGSuFUJbO1hYNYa0CkLsaEV9W4Ju1V7mJh4qlYUxrWwtTF1UTn7MF
mEs0svxy8x8yp44E6iP0ucGiFY/5eHdQqGPler3FGZ61OQx4Rq9XeOkdyiAZ
Nudf1AaehS7ZGUbKJByP3UirX9QcBdELxgyi5NkUATEtuAhDDX0zyeMSE56w
RsBJ+zQ98AHfuC8LnXBB48PT+6ZmAwuMJFH2580f2rfQ8BWxtZdNBPB+H7B0
t2Pul9jQwBzS7L928c53keyvdaS0glKCFq7BAF9+Bc35Jel6JtkXWbiI5l9/
0+x/sR4dr9gmqh2urSm6TP2MkebmFzTZAG5x605TK4tXQ2xhrL4Spg3ZvnXp
NITLqMnNh7uutkfBaENXk5h2mh+kXIy+gwp7mm9wWeIDyG7Ev9waFn8yH3QE
fkNkY7KOjsGHKCZe5g1/Tao9Vp9C5Npk3XvCAHt8bwIxMvDJIyGna0dOVDYY
OV9BaskjGb/W8almRuGC2q6NSnjEhnk23BzsAY5E571W0JK0GX1ozGtXagJs
incNA615dFG6uuOp7C3H18b6UsES7R6uL/XKOYfGsrk2EwFw3WuEKTGDC7KA
AaTM0Zjx9C6Bv6xISwqh7Nqzt+t3JYeLilGe8/jR8f6qYM6CETXwY4oTDwO+
v8UffZ0pRFEAnK/IU0xWoaKrTBWBIc1M9ffN8Y/hltyNM1Dui/YuEXswjBui
vuZQq5tHB8XCBSr5vwsTlDWHTCINBEiBfVeKiuKfpP9tldCsDpTu5VupMTh1
2wDS8Dn/U17Wml+0nkd6N6IdES3aC8xJZjJnrSEeMtbLPfd8todRkxS5OWNP
x7513pJ/8pDcHwZOCL92ty1ZuIBcX9A7TAbcVN+Yztbjy/1TOVkDuVCocaZt
b4lLYgre/I1Qh+i63xCys3PLeNLurMDoCPUtQ4GEpBuUNsrJdRs/26W8mhV8
YcaLDXLSnIrYpF74hGc0jY0EnL7g8emPwYwUSob6SNaFnBdEE8eUG7RDmDic
aU+el8I78zi8HBoXxBOgyedRLHGtB7AUuaVehtgDRs8fXOFR6ZUg8kC13/p0
2beAa+pJY8VmU4+kwNwgdX60lfxrBY/c6eZFRt+1aiU1k+QBoYqtWenij9f0
Lixm1dX64OwDoJz+3I4rlUeSVo5uFp+1Loxom5lC3zbrRErzndoc8pS3Y28b
vDnOvo94Dn+6X0nLM0/QD8zd8rPX9Og7CuMu16xh2a3KK5gt4oFuDInR3Y3X
DeeRHALS8pHPmJsdR+P46P1WAa3F3TgKZe7jVcqfCBxSGSZg97JRp/iivnwJ
JBLLM8dusWnuFI8aX8p+Ww81gEb/CrPp511WimGq3+nZ2g0xnJl4u0+gPReD
veLFdSkX0XNlsPDtAa6LgS3OxsKM5Z22DDWoeXy9f+0JiEaOYGuR5CuSX6xU
7wNpr8fSwtkwl3fKup2zgsMjZwaH9bP90E0dSMY527Cc2T1KtpR5KDu9iDYx
o7PSkfpY1L32bWw4im6+JrQgIan7UvmfhGNKnSwIkn5HLigZC+tnELbcooZZ
zuqs2Ig4h/1Fvswo1+LY0org5B33qmjD6GIO+HIIwXsD18WPG01RlmmWQrag
2SvsUyLK/GIjMPMGyYlkcwoEGpUrXDFJ0D1J8g4ntprFPbG+QkwC9TG0zQoO
OSr0IjU5N6tOHncrRT7ozBRWyX27qEDgpiv+YEwRzM13mS+VkvKL4vcQrZ4b
r+slONbS3HULfEsbSRQW/7Jg+F1hvTP7Cxo4x3ZAdFgxBobOud5bsVoe8bKe
aPbTa2X4N/qy7ANz9bdjm6FA4Y87dbrFtJyoloFGA6WQc01WKPnU1dvOQmQI
h+8A9butX1r+jizoN8lY59zD2sb9SR/LdhvSLLmf3BYveV81t0gW5FVBu4Wk
HpGRpfzVCWC1nUFK298T3Rfd979jdOhD5lzbGb3jICAK7+n8TmwyzTtTS/YJ
dtldH3cUXUF8pz78JOMzrEHWghz0oJMN5evhsDm9sNDgLRM9Ni088k9juxJf
8YaZmdPDcpXEcnPaFHsRofzRJXdrh6alljrTftA8JKzqIfym+JGi/sgT58bf
Y7yLArG53beAHhD6e7zp91vRyH1zipqr3BiPso/yF3u7H9qN7VisUMzud/eQ
7x5yUVuwCcrDsAtQteRnA3hoW7QKSJe7/a9Czk2ErZzeoOyugrWD5Cx+xYen
9UHeZCl9+qHPvGlAvkUds9AbcXrt+EsnF3gd3BNWwWn/7QBFzSfiicBsRdsv
yYi3r252oN1ockXVSB07e53goo6Muxkogicu35vSEMNMlaRmMzyoZlE8BYq6
fskkfA1kEl4aErbONbLBEx/YXhJC60EWanu2p+kJ1yiF65PITXGXKg+EZcJV
dAmortdKHqh1+uWN6Okgt88Ja95HihwHwYLq4TYtfDTvTDpa4jPTZ+6H542/
gADJIYTXhxln93TocxdMs9mTeB05CUKgGNSdyAsBMOLpCXLQP7cYpwnFZ7nJ
1c1r/cLpXcta/J+GxxY1mF5v/XD1PD3nhvaX7eIF/UY5q3hlUefcc7eOKpPa
QTFnuak5ztdnklQzQ71biHsCJ/NDJGdloz9lM4r1jgBBeka8s5wUmKafPJtX
7yzqgFceiBOohnMn8+hYqW9vFX75XyJg0Q0fWbUvwwp7DC1ab7msJwHr8HSl
Piv7qSIv5lEFpu+tDGmHZSjE5HmAqLiK6/cdVLMdlAHyZS0m/xKltx/Ep7DD
pHQWPdpe4MycaetaXjax59sTZ1WJuFRZrbo3VMjBz2cGMVCLIgG8xYCqGX/Q
gDJireDX3a+FCH+12rzfbRgZPpd8HJjsQH9f7vYzmU8yqXE8Zi6yRL0eHWu6
sM8OIEEYhmzZTR3JaH9fLmi/WKX52yqv7BbRb7tPJVdh1AFMNFtPOF9Q6XKE
OhhLZAfOYHLEEgIuLuOwPJMSSkjE8nUlSfTHr1WI0udiiDQFe0dbEpLeIUus
mCnrUqEVyMW+zdvs/thc5l6XM9GewdjgPojNUSIHsDOHlOYJYGc4X0I3CXH7
QDCik0mSZKp+AIjaYIMz4E7MpqQ7vUYAjy3R3C7e5H9B3H223dDPjZRRS/ok
ydTotLpTgYb/cGMJ9egwh/arYtx6rcK0R/9rn05UCgwRBkp8PHbnEDUt4kJ7
EQOAYxxMCHKWuJ3vhbA0P8VX013hret7TsJsfZTLPFNRLEtyly5z49PqEG5U
QG0Wr68Q2y9CVqoY4lJoCfUS4rCMnM0qeBuEwfdcHv26SlXe+d7LPuEljvsp
d/IbCWSPaNHm3T00v4dfVjKYkS3wqOFICyGKHlDbKOteMt7j/gSulAsIjGKx
+SP3YLZZrdm4t/N7s+mCb3bEyRJkEcLN9pemlM8ft1hYwpzz1BZqZqcnn9Nf
HkrehPpblWmGqJVVwkcVSxTNMtSnOWWYpfR89xYEN8YQLHxcNHxzLe1+fLrb
YbttRZKdPP7gbN0Cd7lh64ybQtbk+f6h0uslgejdn8WKcsq+cwWJZ/j/Pd69
40eVsuKT/2gu4VBT9B/vIqGv8vWGSag9odtCP3TOqj8l3CWT8XFraMMH6hWv
i3bIxQ12g0Rc7zXUT1HmpUi7wAfghnEp79If96uCK/29sFxebraqcFjRvBuK
dzqHgqowKnfCl2pnimzjOmHXOYogYDu48fuk8U+STCNz20kEhlVc+lmFY1YL
z4uBtf4Ot0nx6RknAtQjwF5ALn+CmAdRCaCPtwiOYXj6nkJ5gywOwzhFIzmV
6qd6BKJviGV6Id7b62zuBPOToMAmdr+KQXs1w5jIsNTXzT6coF7Be3B2LwAE
hMtutkRRaESsPiW+plBeT9CVRsKZ5/r+pHw7qTX63vHC2VpaSLl/UqyPqO5m
wWfVFkM5MfyYrmAf2b9nEj7G4krOUYEcWJHurVGW1KyJC78CyY+XB7GgJTRR
ETD/Zo2bKWY8QiUYqo5leHut+a4O6nBSqU/39h0EK0jK9XdS72MlN83vUzDc
Ma7fWoUqxZVoDld5dPR3oXtciAlITUW+sUNF8+qysop+pWUWGvvH0Dn8psc9
Fw0l4AO6CTZySeWIV7+iHG3cb9DFPczitqlWMFHLi9WB80kP+gstafjwq+wS
SgSkA9t619Q52XtU2yyzas/LqbWtGKfEhrKWPnYPCe7H1z7jJyPyZgy1OsKk
TzbawvIii72/XR/Hf9YVsRUVrnHQjnTsIoTsmUVvWs/7jWrdHt49A8ufFqay
PUWUs6d/L0gkXorALgXY7XJBlTkMMo5g7YWFK0np50Y6DBE3RP6swTuIHanI
26u81aQmVJgqsPIMf75ErnOyghCfRobE6ce/wX2kGjBIeDvpPT6hl3b9V4yG
MYAOyXluP2H7NdD4U7TH6BRr/oMJTGmpE6OFwtHEGwmMADEKuam2TDwOGnhn
6JjNoDNentUmz0x3kxQM+UcxwSc7aJTDl6SKIhavZLYC1I0jzMrpkRq/knBc
+7Dvmk9LolPplwMBFg2tfb5JQBLDHj/FS8FQZCTXIxby4V2Maf81ycOW7/Uh
r2qWEZBmlpGSuko0J5LD2SPejzeZx+E5I8FV4fWj4QKM8IRhN2OofycHcU9s
5SF+TWGmSd44DBF3XF1kb2d8oPGqbp45AldXBA6esOeRbMUafLsCnbBBAV2X
u0WxUpkGreN6e9nLzPfSnatPkyXq/i/jT8E+7kfq8lD3c0pJ1vKe7mkHLi+3
IKXgg/oHGnSjL+Q6Pz2hmUTlvXXPZ7TuWg9OG8T+TTbvJipi9tr3NV0ZICS1
bSuLDrNrnhMZ7iD9oeSf53UvD4ErTM0r2qEfef32rjv8r5lF5BMe58G1Wra9
8xMcvvHi5fYBIUe1HhGlIuVcgu2D6bANHuQ89r76l7xLgxX0svFocg1hOoHw
4+QRmn6Van42l7uJfBFMXRf3EENZ48TLbpr7m9eKh3u5fGxGWt3BepuEV3zO
m7dfKa/I6DA+j8o32AmgJmQ57qHc2ZQdng8jmMTGMI2X8vKN5ivC+z7MZ1Tx
5nX/RwHhKkwvH/wJeqKVmXNAYS6mXV2WPa/kDMpzNg/GbXb3Zr/m1RoeZcpk
3iY4quTJIQJvLI3Z5cOGJGVqV+pz4VjASbVG8sNi1hy5ITCPQGkK44B4jO/F
4NCidTfS7pEBexQAeDQbxkt0lYLHG2UAQwvMw2QDckR1cAiMYoalLOHfmlmk
fveW0GCIHimVvgczvUSPScvSQEhOd9IJrBQj3MdPI9K9r2sZhIkePdGWYi8B
OlwtQB72JqyLCgUR2Gcy2oSW3n4NLcSjAXeOx/ZpP/MObd5KQiAk/J4t4AZB
DUn6L7nbFG9fMn3lQmM+RMyTo6Gi0wOgO/eMi1Sg3q1ZJh81MKFk41jisxAN
J4F2E1fBOSG9Bj3YrofjFgB7GcopHLn5HXgZGUGa3k2g+/qgjLvPjPijWuLz
8oomFs/tVCByhJyq0WYIt3BUWKDxhw7UOO1nZH9qAOQK71sdk3KTKcr8roy9
SFFXrfP3XJliZcuAY/IKkKH+9I20FPD5DDZXevR9YpKYMz4Egt/KwWzHNH9y
Y45z/Hmhdh71uP6tlYRvBWCmnzvSrwUGzyvWP0tYoKt9E9RziUXYBbHeImqx
WO/Cz1QvSghyWEZ7E+bSvlh4zcfVwBolTxVMGD/U8sOMWaW+gsCqDcoZDxt2
SaNVuVoRcFShhazFDYrWwIY5Pf6pKD2+buXbNRWANqHwK6ANsL+SZAFxKtB0
Z9J/z1JhzYalMZmvEjPmtV+IfU6e6G9g3lghvnkJmcBtMLdEiNNWhPETbt+c
Mh6iTGVH1EPsxAJ/oZbnksmOITgIfce5/NEoZDV8N8lV5S8waU60prQhrPy9
cYMqTdd2M5RlnwgejvfB2wIr5Jr2l42xLmNK8ZnngxfL/NtUfW/kagxNIT1y
DE5R3DSEBmGClx9pRV80vq4rOfi+KPmP9is+Wo3kv+mJc+bjW5EjkwEsl3iB
XEHIgz1GTLTlrsXJn4dEVlMPFJoLUJnDWhhsKr+/lxtFrGif28/+6pv6Mi5x
MzibxO129vHLTKosUhCmt80v4KsgBofCK9ZUWzHtBtOptkRMazIDFB0TZELa
GCAuCAM/aL0APe+75zR55g71MxyLEMt5RKNlF2LIqrx3DPllaDBd2VmEst/F
zRPjhOZwV8UGLUFWv/6e+YbXgXV2SEb7y5IDHTl/EmiLlNk09PRNvpqrUlqK
cWppWv9uOXSw2tJTSJAxrZrEJKdXj4QdkO8vXhbhjT9JN0HYXfoUvy5ObgHt
l3hjsNk0wp3uL1umgpDX2govWSyU5zJryKv3vvbsKDLa0GLy9SPi4Vt1bnOk
Er2Hfmq/UJhgn9VN1cNGIAX8VfHO8/wcQRUtj6MMN3QWUXqgm7ErN16+3/DU
+7/6nTPfAoXpxT2I+jfk5AGAyYgRyNcYgqZM+nF9yLcBuE9rxq1Rp/s0XGrO
SsgdeYSf1t9Isux5mmjhyPys3ttoQH49ImHdPR9JnksecnFD9OPvRXIBEcbE
RebUsFtSTfLtXtE9Nugwz1nqE4DlcAcr4Flw/7+Yll7zgsI24ohAl8+Q0tfa
Cnw5nvqMOGjnz/n3cUBE7dG2srN6ObSOOX2Xpn0nhArglhOWK3REeY+vdS9P
0bvDg/QcnsDSjQKHwAbxnKp64XnXbNU35YBzHyPM/oPAYabzUEm/C49GMmCP
492FO8DsJn+uPoiWth5FBPcPbGQCHU/jEfaS8gL8sx7eGrUDZbaCaLu+Opv9
kIFq3oa0WN7ISQ8JZs/ERwdw/c/AlXEFGJMi+2sIXjbSyO1hZLUFJRsHgH52
mlAmuLLW2ZGN930uxZYz/jlf2Tvl5TmaU0zLrGa7HFtEZ0rp6rkD3R2YU7BJ
SGOZc9i+hj7ggJR898hhFYZ48rW8dnJ2HxA8vWAlnkR1gJSDnIYllLsMznwv
mmSr5QTnWVFMvcLXgO2KQPuW3SpLUkD+TfSmu28t6AIMoftVILyMSC6CFhAA
YNC7TuG5kVxmlhapAJhpegw05bhsoOlSe1GZDlE6W9ENV3sD7jaetB6xf8QN
xbGxyt7PzMwPDECcpDsw0yMlqhxI0AIzcYHnv0Q7UHlM5esm0PA8EweooR72
UbnG1W5S0ZIMOF7UCpr/2FuCXi6knLuEFvy4b7ofCDI3i2nI/FEzxLeGJqb4
pPwC00u8NF0bE6P/NFtyLRUF0Y1U+LH94YuFXVo59nEX4nsLnTd9xpEiJP0Y
9hrv5/1zgkM2lw6eaKmQy9Ifsr9zdduKLyz5F+xuedwzwRl0m9UK7sqyY29T
P/krOuvCKm9QCZq9ulsiEjvy9FboSoMNQINNmWLbs5glEW6IBleRURdY4r4Z
wLL4OI4poCINa20TvMTlcikMHmT6t6Y9FFJALbwtSHJqMzrT8TkeVeFoh/ev
5lvYq/l5hFWa/N+JLyr2AIVHfydrKfL+Pqw2i/QrN5ZU2L1cQ+cIE7Kz/Stc
WWaMt7BE6O74N1eWg2mIYD9jtVTEmPXn/Bke1dErMFU6UVydWrjjnyZMMfQx
FVARqlJoocUhlceuzPhpqmKhfULbkujb7fyG3PgkAmtJj2Sq0sL9RtZznWe7
ou8PIimiphTMMLx448+qCDxN+a2hg2LG0JNVcI4y2N9WBHJAYZiINYf+VcdH
80SP0Z4WbP2t+cp2WJxOZmpPt96v2lEzs3T3uQP3N8WpA3143Uh3TFktCsAj
W35NLbG6O2/9xOGuqJkeas0+x20+F09Feekh02Pi4ocOrbt9aZxjwzEnfcMo
bdRN5OjEBvkCaQGWIhtipCBXDLGgWrRxk9ZK9dXNaPEtsrBQh+/DD8ka6Df0
/X+YKFEz6CqxsQkySyvUlTVirJ/B+yKMdlSAk0fbGW03jOLcRC9jTP03KqVc
JyUXkpg3w/lNJpYnH9wYOwefqz0VyVKFOS5ACuCXg6GtBCyRqGZ563jMquCR
L2fA0yiAG6g/npG+Y0jKq89TEcnRu4iAKT2GYJJaM399XKVC+5jslH18rSXi
Rm1UEq1ZQmlctn4aI9hl5gwr9d85aZFhaVDEK/GoC/BRCi14Ii0jNfoPg9T3
uPJhpNFza867jDnw5tC45oncWws5vBNSdfnsi43ddyu0lbOdtC7AZaZ0q+sq
pF4wNLEFRBDy22kbfFS1iBve9PKw4eXUDsN4mg1uI7Lb6BoBLHp+mf7n6Tz2
wO7zANTzx0HCEaiWHUQ3is2MPwXFH0nm/wYg/bgpd/TAqyzFUPxHkCWsFA4C
28Ym2nnPHx0FBiVVAEXRpZ3kVYy8AYARMlq3Lu76/+2wb8UrLjvur8VkIm+n
Mva41DzEExogpno/MXGXeJ851zbP1quClsj0r0dLlVgaeJ4B9/d5wjEaCUui
7G6SXMCMyTC3DX4mArztU3Xhy82t24D0mRQlsZd/TdkK96ryM9nMZFZhmiDa
chokMKAg1EirqEL0VOE5tOHctePrG/HE/YpSTLoMEUy4QQ3In9MomUFA6paS
NkwY5Vj3Bh8rlDA/duS9kNs8aj8cz2OYHu+kf/FI4H9cxxUMTCDK2yb106qe
4w94rdXZvv0O2cltDzLnhReDrRpTavu2SbRMgTa34+w/QHWbOoHNL3oHFesh
3Z8lIdihSIWt/IKNBA1uJ8qiuwIqd/T2Mr7PdAL3r7O1yV21WvOb2Xte3tqk
a5AjQTiiAESyT5V2gbd7ZG4KaUGCvJb6EWexX1Tu1ZTv3sOfitWNiX36QHpd
KJrNAHboay2T5FiuYOSps7Z8QlVJ42KVzmUE7tTkqHY8R8Y2EzWGUGRRU+rx
seCsmZRAck1bAmk+WVA8TZMN3p+aEfy+SUe9HHcTLCelxBNLpDV7Fw9wO2DL
8Pjgs5Sgol9Np6ZYl2hOELnlc5engvTOUqdliWuhYUNH7IaKJ7U3ZABjbtet
DtE6o5jhhqtrzOs8VdUW9XrssK3jMdyhPQnARIFe5AmDBlrhldTc6fxhh2oZ
zUZT/x0Hcaq4B1/yWh15hZW7QS/kV46MpFSkh3LNl2399Myn6rca568XgJa4
ZJ59JnedEGUV3e2nCwl775craLK/cbmxgq2wRi3kl0lFfCtFdkF436Nvx8Cb
/kNwwoNN9BHv8HYKjWEv3DsCrED4Gmgzj+R6QzohV4g1d05LEToRAQ1xBE3u
LQsZsNOpwtpsBpnT0WfFkDDuWfYCgAEOA4ot475qTlaB9z+HOjpf+MF48K+q
sKyoexDqBLM8G3twD8llKEdWHql6CX7XzEy6XMr6JqfIEzM8gwPKlw/4XOD+
BOTDMfqkaphyIZDEm+WhHISwi6keu08otuTLdg1d6GUFVx2Budh7/nkvoUlB
EcbZlwaqznNW3swLK0U1xYLa1BQZVv/GoKNjDf61wqrr+hKNGFhzLasP6Yi0
Bno1M4udpEgESDKrEV26cpP2k9XomCYIBiVChXXcbqwxcfRzT37oz+TIKEgG
EUvVT6NhgedwTaTecCkQWbfQUAZfha0crwnudq9T1YPsJSInED/RbDsNpFVT
+hG+DebZjW+58zseyOpoqwUzT9g0QIb2vcfyBUxiU5KyxxNs7kcq+u7FHPXQ
L133tZdmDcIF5IuutoHalObwqw4dUO2t+pAH1zLWvjjLvJzE6xEuUOAX4WjH
Ei7Iacd1Fy9XNkd59vLVu3kHL4Ms8mUzIrvoD0SsdrXwwNDy/YR5mgk0Z8tN
uPaQMQvtyb/mvoeOXOYxgEXABSFOl2Df6Sjm5vFbiLMW8T1xFuu2IoIn0ZcD
rpf4TccxF0jAKOKJkiH+LmMeOUCOz/d/nXkAOItyJ3+A8zgMxiy9JTHsao3p
pTnZOTSTAgJ6ZIxMtZ1LwQ0zFL/PpnUzY4bErfBUnZlkhp+KNZFzwr228Ydv
x50V8JS0qskwaD//+F2DkO3VFQokELu8QJksn8MOw17gQqESv/cWHs7amqV6
rpvtRS/gFwuVmH3MGmAGjoEF676UU0cIFsM5U/MEC3QaH28OUAW8m1jHju4x
vbbuLU56BD59o3jk+eMMU8xFSelCHtz+fWwwjPhbfAVg2Jsg6KhMONGnhS9f
Ix8UVID/kGOufUsLmnaWefrpL/JUDekFsmKp1ldjqZPZEjMciJLRsX6ykDDE
ZrDBrxWNVGSQpBIkZGOELyLjK/2Qoa4wdgWq03TIHVIMnJUO3kQLGXy2iSY3
UBLmASZpRN/FUQLBZrY/PquGwAQbAYUDBuw2uaa2JIiFYECDh7Q1t+S+pvyr
aArzR6+vRkKYH5wUxh3DPN+k5QKTfOoLyO+te5FDAmGzqbSm6VpIiilnjjhR
2nRqvUuYaYryx9vEBqAouvQMEP2Nss2eIGLyTfbWYgbWtFPXPLWKqI15aazN
TnTZHPUF2kZ+am4Nipx+upXzrr5lUt9mMdNK27LZP+qqTkGq7jvP5fDWvsG6
vJErS9dXcgAOSOerFzkWN22y5VXg31XMB8uhHTqgjJJy21Cw9THAN88Ux4cw
QN1gXO+PbzjuHDuaD8JgkpZwcl7/MjfQ6Vd0Sc7oTppCLvAEMW2TwaB4F9n3
Wn9NKi7Fnk1QR/H21giDVYTTitQdOUOqrya9HHZjrVOxaG3wtf0MD2JX0lf2
YekmiBzRdOL4C0totvIR3DqzA1orVs9kEoJhbgIgdrI1+2FAW1Xy9MSnccLj
RQXyBi8EAQM7ghrj0FXG4S4lOq9mQJz5vUAJ/1WP8AMnzCc7ltYZGpp/qNNq
wzSRZ8ZiCYd7oscbz9u3dwE5EXaUrSOg05IGy4ctSkdL+PUZxKBXSrjaEU3f
6vqzFXvAA72dFR9ypTuepcut2glJslFniG/hnym6rsq3DakYjPUFpfrH+EzH
ivaOMLOL08Pg3+vdAP1JwZEDLG8wEyoMoglJFDGAr55Eq6PsPtVUPjfyLAVe
3cefSSDEiaHa+q2SGXRi9HMnszlqK/u0doJhXgmR7Ci6QlUtIGxe/eYs6Dsa
q510CsIVSnTY1Jcv6oKgxBWyFi5Rv4i6auTLyfD6mOiSVkjvrqGczDdY6akf
NJY+wOX9Rn3buVpk1bFHjMoq/lgXYTbSZymTARSfufn/9zdVuG0Okez5SXa1
lFnWRWQixvPZEDhL2mgJzfZI46gb+Bm76xYIhXVT5EbnpFmBvvWzpiCtvRaF
NIKuMC6ryPw5W3cv45xb6hJDztxcAUBtgi0G3wy6FPKVHZqhWx3UItwKXXTz
kSBaFY6ZD+QXeTlCx3n9pZLGKQwG0rVblz4DOsGNVPhH+ppGL4OMQMDX6nXp
n+5dPDUMJ2QKr+NOX7z+N3zQX3k1aXX6fD+hyw3lu+SCxM3OHfdQHE4DEl6k
D49eonMY4HzptbT8e0vH59/+stKVhomFvM65sMuszWxcar08+NxpTC7bEuPD
o6bFxWPP4aPny2Tm1WA1/tud723lpzZNwXCec5Cu5YPl3SzdG1dI9Mi3I0Wa
xNIw+yjtAD4YSblEwhtmuVuBVxvhHdUX9+66Ke+o3ol91thJKMzTBP+12yam
fOl7fGaVy0awBpys3xsX71+mEjsSuTyPQlKkGPO/BkpGQEnDA5rz5Ln20yQ6
PXIZ8sIJkg0xca7Oi/gM8gCJLUzvY61eh1UocpuRCbCg6g3h/btRXEEK8yhg
+QS8A8Ct+5rAhqlCpuPW17d96jBY/DPcAh5zmvD/opcViVHDFa0dRULf0YCS
q3yixxhW3D76cCwJZQzNwMoX+EIoN9Rz6yBNSoezBpNEI2hzE8NOlg/ewgkX
NwEc6uiiaUGEFn2mmVntH8ZcGzr13CraIrfXed6u2ghijHev+OWuEWljDJYZ
59irzQ4mGTVypffmBnN9ErnFuMISAM0SC8pnsGH89gPkr75nvN42jwHhW3yt
e0iGW+HMGGxyc7EDNsb1XkyxQ2PmRJ2prdCymFFC11Ofb25DZMPKhJag2bMJ
qNkSNdXgLE3gcl9bBd7ZNoq3OFh2m/NzPInqwCRbfVYXL5MmIDwc05QY2zQz
hrsbOVQwTG3FQ0G+WGrpTnf1qR0epZ7CBx7nZuHJ+FRiKsUom+xrAgXBnR8D
Vkz/Aku6oIDu1ggAWtAJdasI2LIWy+gix1Xpfov2uG3ECL0MTmT2/Csh1+bp
zk1Tnp+MdKDMJio3gvTjjinpn6JG52i79OsW7CLgO2OI0XaBnLJSW1Wwfd5q
KVBzMIj4MCFAaCDJeoGCrKg6+Czro5XgjAZKn0WDwi1jSZy6dtoAq5lB7HWR
byVYVNjPrVamQwxqB8QKIJe7BuSrZurjFa7eOa7cfzrvyft6BycVXG9nBrUz
o/sUTszdvSyYkkelsHnI4Rm6eRICY9hYATmxLp4B1jli51KsXjnzgsZMr0gj
0b2DPqBuk9P7GQQJ7fGmq18ZSPreSuTCM9JKp3JhdN4BdCbPNQk6W9B9Fnf7
lN6NXHWNN9cJqeqiJ8mDpiWoNQ6PI6GFD0+RnI4RqY3/QV6VaXAcyXe6tDgS
w+qoCBg+EdJMsKvQrh330hjvyf2jQkG+oeAAjJvcb+ppb39883IjBYB3oqib
U57Iv1r8zlGTGYz8PHuK0dN7uaFkCUQ81ZLNN8vbpDb29p3R9ikOLd5fjKUI
W9I8VP9KVMS4tPH5PhdnZR7Clz2kFwSiyRMSvhUu20ZUmaB589c969qja+KL
Z/0p13QAnjLxIO8gnnCvfUlr+Hw0svbpl2YWjdr8IbiXQQr6M0zY086XE6eV
vkXkamHHDPAd/SgP08kwcZpOcy/moVvTp6dn4L1EhbxH+P9MyExr2+jN4u2l
dFg+MExgwtCrYR4FdQjSR6yw7ox4njjowIvZJoS+XrJekA02os0dU413MCTJ
2IDFEVeWa7NpWf5d1yZg0ex18eUpQ2Kvu49fTO0fiQgk2a4bLWN0ewvF141A
r30fE1RE84Rgqx/6T9tS2YrOaZnoPZffb/hEMyrqUgcXZ0H+fSw936b2ZRJa
c42RArRWpCJrzUdtiVgRpHlSiYMKBA09TS5yO/Q0pZq/VRWuki0ynItXJSD7
rcSEAumIXNWgxruS14cXhtPqFVpvgXcArkx8UT1BwwZhHmpT2ILMj3YA2pes
meDDT+7poqZeMdr41+D5D1nXaepyoowE4ciAYba7aF4M0SBdpgQbX5x3yxq/
ijMM2lScPZ8Cy82mYILcuNLLL2kj0IlINvKPfHOc6ntxFj43DL/HvLBH1l1D
Rw7c9iVpIsL9fcu4KbDt5Nmcw4qDE3B2+1B87V/bF/upgqbAPtpAAf4EHGPB
bPC2VHFI1+x4x51wcsYHktvXEqVoNaf07WWRHIuibupGvz+u9Pgkp2TGA51r
GepE58owxykeutg3hexzW2orAyYAkqIuo1/bD2l25byuQIIXNbCzF6H0GpC3
jvxqsXZEnOitl9Oux0XceVD5yJMVemMVEcjN8J27Yiq1txhJJjxLW6BOVNBw
JyebBq/fKN+XnFO88R1/jbnuYdIJr9HfD5luNmzY2PvPfqAgvXAONoQqrKbx
B81eX3OpxsGp++HBaMkj9SkOATMcWf4jeD4mXnF1VDQjQrWBmFBVBe22Z89+
5ugfe3DPh5oFTtvJY7Nbb1gaqeqiHtjFQlAZFLZpTF+6lALZ9sWp20U/e9V0
cXAeRsPeAaReCcvWJEq782/xOAq4vCwrGFIpOKkmWQfTLav5cE+cqJbaI6CS
PYetCvJLLvOjTMoWOXSAs7I1FRGQaG0qnhZXAICit4KJukCKUpqear2gS+/2
m7B2B5g1KJGDupIJhuIJFL6pMPAMJx5KmTwDDBgFGsq4seDeGwsk2CwxW85H
dq99W+40NymtfTfPzDn7N/UZgFmIoF9Wq+fKSzH0IFJj2WjbeeWpX6odwPuJ
HYrVudG590GsH8hJngO+YndB7BTa+EanC0MFzfn6NMjwdB6fe1dpB5pKgSG8
GemZa2zweBKdCdu+145KPwuBTLvvsLGPFCJ9gizcTDFxjnZl82ART6J6n6AJ
/pheXCB/SUl6Dp3nXVVfMudmrIzoy2szWh4giso6SOHcPxtO6PnZkRCM/Av6
e6s/TbvWDx0dQUZlJnAGhYCxtjW4qol58CKF1xkuUZBLpRb5uAy23JpMEwES
7GQk8spxQ84K94I0oYuSPSKmY7anLsW7GHhEJ8zSW1AhiCfFAjCF4ZCib9UV
IJ3UdLIa9VRE3CSBbgQWb67zVSKdXgLNiOO7HtKlqHvLs6tYCciD/QQu2v4h
XYYbl0LL+BTbUq4fvA/wklKb9SgmXsk4r3nPeQGu6Rl9hx/TwmZsydUYhXxp
ThG+IF3yml5YBT+6nPhyBcMFtCGD2SI2ccnY41gN/3j3hvrH2bQZeHzSPW2D
mVQfjUngimw5HgVTkZrBkB5DLAEXsWMVTxv2wSQ5aMxiTn2TrtPzNt0oSr+F
NxQK7DN/IdqPTrK6aCntWKtx2BooiaoPJW5kVczMez2eb2KrrTOu9npUc07H
ZexVyxWOl5nUpSqnThCOrx5Qc2UYxczd5uIWqoQL0zQTJR2rs9iHSgih9NgI
D3+XsMc/ymLsM7rm+CjMiZjNEUYF5qCT8kqne9DLbgP0DweRY28bzYb/GPDi
ss5cRDl/69y100+ct52eQLe8MEtCx+HbBW0psM44jouvLIrZLGNAcS3004AD
Rj5GVB+uRu9JKiI7xFWM/lxKUuxZlAKBxvF+MeokGB9pBIQt6jTchhVxCT2I
j8RTexYDwi5HFqTQmW/YEtV7y0qUlFqHSuHnB4oANrvrr9MScZiNTK6eYOUT
zheW9gx2kFRNiMkhBI0n5N/AxFKI8S3Ay4T7FkbH7Ogq0ctQhecjmXNEur87
3OrW3HcZusc3et8i8SP4bzgmvMsAL/oNrnwKBrMuVgJ8REJmIoJmiO6f+UaI
7yXa5WQObNAZp+x+zhvxhZhwm4+38m1go+ob0x+eF1hIhfLRlkeVauo8Ar9q
1mS3exfnxF8xrq8ErHhJlqHx8JlYrc6EnsI3LGkp5Ls8vHYW/lOTny618XX2
KlTTSwUFkbT93k6sxcyEcZ8K61+bCKZy/mWl44wz/Q2aUG4CjSj8/VqrX927
A6ca1EkTTC5iOFQDajlILWdXpiNFJokw5q2RL1K+/DoBMbGRAAQv7R/fU2Et
4ZEvE3P1MF0igWkZlfwCujVgFnVx4z6duA9duebZ+Om4xR6A045cH/vYxWPk
Gjji9W6DfVHXeyVl8Qwhoityh4mnFCU0J3x+7dXhnT0LhQDUidaiK6Qcb026
fFZc9EZmE1YLlj57edVY8A+AzW/hc5/fpe20u6nEZRcO1YSEsxeTMSYQ6QqH
rXIx/Uv7npa4tTXSiXi7JkgbUthK0cjvDzsdIP4+DufeOjPY2JrRG0LKqids
JOJ/vIuWltCGJ4ELLRCd7EDhq6jDP2Iz5t8zoFmtIqC8FWpUqApVUx6G5QaR
oC2FKxDSjZqZcT5FLYJFik01jtN7khnz5wLA0BPSIhdJo5sVFcswHz+XGcZU
FZKJmU0qg1OfVM2yz3zbbJQcB78ZuTsDa2+oQSw1nTSPtqL/aCiaxT/fiX2Q
QGyK6Zp+bd6/ilk2v9xYDbT/2km8QwYWfLsUvSsTLsFSrGHs9Lf/fk29prCe
XYcOrc3Hq3NbZkcSQKdkWLG0Om+vyQrMPvgvsV+69NqY+UIi+dT39ja1tFMW
pMosazC52MA9SPwKP5Sew5eld+PqIDfTkL6mQhV0I3bmwVi/CH1eKlh8+lZ1
YCC6nfxM2Oq4vcs8BYW73KxH1MtpGsGWpk4fs86MENXarq+vgvAzkLZpRU4R
9P4GUBQvcq7yPJREZKsbtiyH9CS+mNRGbLAWfJo3X6wPgOIXEzQ+NLsaPuJR
4gzRB0WjS5lFvuFAUD76FFKMGS2lYW/Bo6c/5/NCgnmfMoLSfpOaXmAr/Vrv
YN4v3fp2GzEFkUJ/O58a5rHItu3mhbJVuVHukFmj0ZbZbJ1/5763quqdjy/g
7w2xzRDuCjhAUnk9zzwttbBVgMjpmQt4pqkaKsR4h15CU6eksVkAm8B/eoxF
oZo4nF8rYrvytKqYDB4FI9SBtXXqiAXQVyaODNxKZ1oqNPuH6ej+ZaUqCLT0
XoKlGgzYfL2PoaUXqtljx107ZWxZDseuRypfI8SA7zo7QwfLN0mETLbUe0Rv
mOUynZRjQ4JAd46bZLAy53njM+t4xHTQ1ZO9iL4OiGdlEAeGcYtWwct1OBih
DiObnjwbMTxLOWHBvWAkLjIOaBxPUHp/W43i04Dk1PF/lreGasigpSoHfsCs
nHAfx+Wxd6v4n5i3PBE3lj58qitkJKZ9DWNQ4dqhbnXPlgN1WVk9Rs2uZzop
QR5tXyfUxh73eejq0JAvq7oWeNb8NJ0cRd7z3pAr5bdBgROHDQ4ivSEQ8lG9
QEmR10d6Ui0t0XizPqLI+s9zm0eVgPDMt4LnMsu3IqJfmNXDgkn8F1v+9iEi
6cBDf+PwPT0js+V/7kWpXD6IgIIY2OFdsARgAPyCI1CAHspMjZoUywXwpbvF
U6cGEFc+DVpqEffgYO2Q53JA9kbwAuTfU8HLTDUBN2VT3KfUYOU2b7yasn9/
sy1+RmSTCfpnpjV5AWPxWNt287x4tLL8fH2pAeyL2o7tyNyhl+5yvLGGM6fk
wALlNs/H7FM35RHqFCPIcE8U64ZDTdAj+AVZRFaBw37qeG+tMCPR89HyHB2c
m6e8p1WL8vbuVjhMqsgOkdQmnINjob/nu5Wvhg7qWJoVt4zCIorL6HzdtaAr
0vNtqDPclzFY/H1NrFEgDDggC+/TjYKa2+dQ9MVfRn66WfXOfmcOpS8V2x5A
YaM0pQNjplk12iGNsICD++cgb5olcBeCjxJqzCJ5soML3n3wIqzfmulNjvEa
wsJbJhMQipnWg3jTumSHzBdLCjd/IZ7NYQlC1Je+bS5rx/RuS0sJv5tqxVWK
Xj34CetbT4w2V00yRCL3BoVxFLlg2MuZOki1q8PUU9F0uI6GNcoH6vp3TXcz
IwZOWDwTHcfhGJfahSU/dOiA3nG09xKN4gxvlD/AOm79iyGIgGVjXWzpO0zW
jDBI/a69NcEZgM5ZFcpg1T/Gb/sKN+dyYSG4NNwh8qFbVYaBs+uxwJGwFUxC
IxqIoe9rjAB3rwu0+/1QGwIkbWNBRQIBMnPlHn5hfnnJ0UmTixR+eLNp8I7A
SqmiNe5NY+eUyZNocb66Hm58i26q0Wqdxp8CchR3m4USJUWc1+Bj84ZfHlsI
As4pQ/nUMBixW5exv8cdS5XAfOy3U3vT0PFJY0Iva2mX5EJdcHdwXQ0pWABc
tIYpwAppRNO3dcFO4fs7p/JRK/1J1bxTk30ZwAU6oL9605DRxG++sQ33G+rq
2RXpNj3ZGebgua3cqPkQh9AsVCzjZ0dEk/lr32QutQneleb8uFQAdc7vHTpt
9tIGawMnaMoNbF86j7G3D7jlFG/p/vCl0b/oBYcVfIJZiiNk399B2rnMpfn1
iMjOMhsTsVJepMsmoY1HVoZdq6B4vcYtvvMuPRBWMf9IcYGh3IuJnBiQsdGz
L3eDc7/qoaSS+/2PdQcEb1JXCEp4rP2whDdXopd0G7VI36ZGy5K9MPgjjpDW
63vgDoHUueQEkErjxVE9lYZXvAXAzwdCMrnl6opdF/W70XYuSXCmOisQgVi5
KS3B3cUSPIzRhFb5iXPJfwRitJjifmyPmvje91O1l8FlMM7sAv7OHOHghv6U
OpnpyhQI3cz5zhGj1QkCAx0wZIEhKECUmuB4PywENvCBhx7lO9shRLHwrwpI
hkYopNKTY1YQwYAU13BPtWCHHEVTWdBrTdINEts8hNqgXMJ6gO6XW3gh56CB
0nR6mSEfOVfe07yG8U6UQwwkgYtF/HV0hooHFfeY/X/dS9a42jdh+exZNNaT
NjKByhWJKSyvxdo/ZMf4FBHM02EmuMUaKbQXmXxs0Ay2hIIxsWr5Y0nWkanI
7byJ0COv3Fee8SgPnSTT393Oom1t5AnalYOrX280YsVoM/3bSSgMY4+85o+t
sj+qawxRszny/gkmvxHpaeCrFBJ6/Kbp2VGXo/hXtCtgLP2oNFrzwKJR0KhI
YxDkmcqfRUhfJXO5uniGSSqus7NN+8d0+F1Bnf+LjQA0loRORLV5W83iMYne
ga3aE43AO3iGJKVL0hP1MzzOQj80A8sejJgS6KPAdqaC7y/GL3BvWRLkTYb7
OOk/u4Grdp6GePhGoQVYMLjszvewsLhYRfFevv1PDvRbMpSCzlAwYsAnENSw
O8q/ChN7ONpRRWfuiGhzeUl9CfIDQ4cR2qLIjZqg51p+hMwaDyegl8LFxxQp
Ye7yvf1apN1xD9vstV6T/E9UHPzP049ITXyMw6Snp6WC0LI5Vs0Ji7ttL+8L
rQMWAtBDmgHNNYzCTNl2glVQiMFV0rwUCD1SA4MmNW2c5YSQ5ZLfyWOZhtib
YmTV2nOUgm7qXf5Wp396SA1IO76cv/hPtokbqo5hkrLAoDuZ/v7456ro1EEM
ESh5kYakA39Iu7rgSxbL3xaseAe87GuNfMpnyzvDeWFJS8cKz7nUtZNS/XCJ
I+olw0N8myF5jXAb7mOyFvtNmZkkzEFirBNjbLeFg5BvI43vecG5sSu+t83c
HvPbTNty40ABaLz4eWNCktK7Wy7sR/pwHn0MD9NuRBjD8dwucY7SEUAbzPTg
jWhqOlz3JgYt1oUdEpLBMmLcsZUCu/2arvwFV3wF0HsSxY0XsP0RNCSuB4eA
u96xS+Tk0vPtWpy9cLo8yalBOcjlDlOV7j8CGoLahpg4Z5H20zckRreOdPdW
oL1Lcn4I0rDSkL9oYxRocQBeO3C5PNieTcMVwTOYHLEQ8Gq6F/xsu1QT9tzg
kQElH/JKeukveZPUTRh7zTBY3oTbLnNemmxHqAKkdX+joDCmsRWFxT4Tu9F2
XApF7gFK1j85raGAH8xhwPbU1pGtd2PpA0zpYFgOjh+rMTNtI7F27mDmQ/WU
BwNbSOAeVXz5kQlHSeu/xnL+qbgPX7xNcwGdJMVDdcVmiq1983m9c+3k78Dt
k2n7mKs5iTaQy5zb8LhfQpQFeTCutt6dl0h7TcyeiC8qSSPZGuE6PVbu/NWa
hsuKHZrur2xsLNbFLE4lApNNcZFgHD5NdhVUNAmi67CmvmLdMEE5zr5HHDec
qYTqi5Oz+T5QrPPMctEfW760RQUSUOgx03jelTcLvQk5QBziQE+EuifULXgE
fBAndmw3EF12/C9W5PgsCdK6INkX/FSIpKaKSt7Hg3IxjyZO9iU/nQRAJaRC
Qko3z+xrXJQswCyTJePmJkcCHikF2d1B5uVnkTbilbzoNHB2eJECOKCaBnaP
UZ441lvc8ZvHL4MhO25yj+wdWhuW6OtwHP82w5EJMc6KGuQVWkKrQXC1GZSw
WU/nKH6ZZ6tFjN7fob8O21G9OxjppxuEitfXRAuQNoAKVItaISPgJz7EL+3C
kcZhWTMcMfzNaG3+8gRzziQzgAejcGz9myXY6JViBZm2vDLAGtHz3kYIuE9G
9x6rXcsiGbOUOjFXumhcLdXnr3xsocS7rYACVo+ovN8KBU1pHgN3c/9lsAqT
Xeo0P2nNW2IXPfXmP6ebr8uEvbXz4b5VHOufpFcEow+Wg8L8xJTk952De0Tv
XGQ5yv6TFue7eSYQf3fXXemjnnNe6em5RX8SlCAKz8+YukvuRnBCFR3LL+Tx
6u1oA9QDZdm1p8waJJT1zRPjRKkRE0PPI4TZh0Z5mFolvEErUjmZ6qai31AD
4qasgUtaHid/bbSFQS6souqguNhg2GiXEETISoOKEyejkleqeHfHY+LBrc/u
/vtJKtZKHiuAucpTy2AivEpM5cWxxBkyNYT6DSW+K4iaKYY96ZRInuoNel9d
NHRUmdIYG+DsOdDs0ItfAp0cstZmocY6pCJD75qBkpFFLd3P41iQsoeoeaFr
2aWStu3uwiu9pCNbWp3GaeOLamjDSqfuQr4WZBOHnLT9GDj4dqjeuoxuaB26
QWA77O/Ujn1aCqfV8QaivSemLwiMxacHXN6d4uzCWonA0ZKTsjw1itXAi0l3
xyOegSwc86PcQZdOWiNvM1ar0wSvp05EO8cZ7R/TXUybA9+ld3XKokveyd+r
jMbfSj0oY8Nivgj4JlTwpZIR2s3E+pGc0YdeICt61azzhEI+QfN+NJ5SFIsi
fROyO61e9dqNv67apVR++B5CoXxQuAlYdfegWiMeAXax3e3iazF31zIpWKqK
JlX6GqAgflebF7RSH8JBtS1LGzfV6dGFTeEc6MR2XsZV59PG/pvLB0ylH5Tl
hfckXoDMfY78FyIfC9CigkY6w+CvcnCuvkYcbRS3Kao6PT1EZRN3HR2fc1gf
OX3eZbmdWBAT1QE/7t9Ls+kPKzmjqpVPAYgjSA/Ax6RBuhSMzjbSwBxiDFU+
2knFm+McWcn1eiW002m1czZr6sUxvT/No/4LB/tENGYNDlyzKgZPwz7E/cZL
CObRW5pxCVIxnQRDHnWUcyV4oSdep4Fv1XXImV2tY4lQUXiuqYpnjeNpmkUq
jVDpz1Ms3I5DbE42m9AbdcN/FLSyYy7X3RZG/xpylamY/oYHR6qlpeIm6Lrq
w3TpQWNre3dAWdhtXZBypAG5bKYS2OriYiAGGDC/TPZcvyVPqJRBegKs76TH
v2fYVqQfSDdRRDP/HxtrerOhDGdOYxZ1V2kQsWJAy38Cx6VJabXo94uTHM6p
G4AFAzx5SGuWnbwffucrkn6dSZpbRWbRCiF+s7/+T/G1gAIhxssS+d5YTMWf
BmcT0BrUGsL4PjnTj6dvRpDCbTOkikCdwdIgnXGm5aUUfSPnsIOfuYOiYdrS
leSBeX5shsBTDupJ6VQFF+wLW6/AfXdeeU336cEPZwqxUD1T7D+Gc9o5jp+l
+K7Hi/1c3VByk7QI2leKj4QQXtGG2w3JQRuH4kE1Cu0nj0tVlPMNtUqkCfaT
grHYbyQuL7NdQoXfXagCOS+3VVYnONt5+72jYynNmMo3T8jZ60jP6aJWYq7v
8+mlRCZxWwlJI/+ggkrELFREMOCdDsy7cTjpcSXRfhAQ/nPAj8H79YfUSohp
459/4Fcgs5W37k+0GhL7N2u1uS0UIRt0o/cD4OhyhdNiNczOhuJhgt58qTri
bzly09o7tkNjwwGCNlD8s86eQLUO2CgwxmeuA6QHwqkS0/Rzq7erakI6KLl6
D0SRbwNd6NlwGpb1uqOVw3i4BMDtkrxSi+o6S0Zoc8C2h0xQXM8XrkCfTZDp
MjHNqjqVgxOFsvKXMFdaB1VLpa4TXrNnP7IgAyWJ505DvHBM5ThIixL8IDtV
n7F6/ZqbIcoRATBXLPvVUZ9+RDZ2mW5JbjLECCdM1sYIlbxkpDbc6LLqxW4l
Hd98vyFJJnXGZ/+cGyPuioNFrpEL8wI6dEqoPBhTQDSO9xg82yff1D360xwY
EbEJ1K6xKGGwtCZG6B1OTY1mqOqhjzK80ovp5wKkeoFY+D0iHmHxbSVLOoXk
htGqXTvXEcOPGEtByRU90sWcSDgeaktIoGg31puRAKFaxj+KkGQ2pyTjMeTx
y7oCZH6Y4879M/TlhX8Ba7FsEObtvoZ2X/+XgSM67j7nnRihtNF6UiyiOiy5
xBuSCFZnS5AYgLrzObYzCHOWXTjRRipHQFC9vrL58HiicaRsGUlGZhlhdR4I
4YEgpAunZ/kOYTTeTjn4po5wU2dEruKAZ4mGrTqYvr+epzWAUi8R9JOHxCI/
sKZM7ErGEY0reNhv57lGuKlAx0pXBZxgGS2CoTx3xlnpn7OA6hJ2ifLkehfa
jDDZ/HOvEVjzrP7/K+P0Kku+mx8vPn0ca1+NtGADNOGpGzl0F/8cChE/vE+x
OKu0LVjOnK8sqwTkjXULsILP1VgQRUAdgy+n+oM8x17VZZw+0bOJVQbB6Y1a
GJZ5pGXSIU0DpVXIgwmqOZ8V9d1mqcrxe9XkTjyzGYslEPaQijWrWI55f7kn
8apegRPiCbyJHmfcS7N/VVdB0ajpnoHVtQPVTiSbSEw2xVxkKURFjVdDjEGL
RwC+8R58HOin/d8PcM4ORrFsNC4NbMRMixLBYNHbd/S4uCS0sPDjq5z2stHd
lvnBA7k3Hw8lh/ON0ZXx+x9J3UxyI/jiWmjyn02jdt5FNMtp5yOhSPfQ+Rwz
6kX57hoaC16XLHd+QBAeRgi7lJUfBsXHi7Q7IjAVJlBSlPaQd4fwYqw/Fmqk
5z5TciIILSljCOOqV7nHMQEljdoH6lVfSLLFbbmEsf9Fu/3EvNSlisinhZY3
bEBzHADQlSedCFCRD4fIj1LKrzAD9HQXJ1ATMya4OmiJfTnIX5ISp1KpwvEu
3BfmU1EzvghZNFBUMZ1S2jm09byzP2hn7QAM3w20r8Xyr9PCL9EYhKIi9D5s
AtAEY/wGmbh/I1Bd5GQebEonSe+1dajwI0m+Qlii+jZ3zNoilWKlTvY/b3ZW
Y83VkOZg7LfG7PQ6MtfrtNJIuDGF5CJ36VU1VeBR/6k//N42FiqOZB+nLcXh
60qaulOLQTYoRzEtL99RLp82DXb4PrniNI0zEM0YKMLCkcMc+Zjgu8if9b01
V1tdbw842lV78uAnbxogpOST9MRPTXgjEQgptJIl8RtIytKJQrtegYxckI5g
moaYKvrQ2krrZ+EcfbO+OanhBMDQJto7iN1WkgdTXz4/lCWxrID2FVt2S8ou
+TC+txJEbUH5Larf5RrZJBTMCUOkz9rzCb2AIiMe2fRav5FEDjHT0R2q7wRE
9dC+15eXQiSxAxy0lCxVTn0jbRW9QMxYDPLXiT43FZIkPHy5kD7C0v8POW6E
RAlt3YxI2R+9vNbUzsX58yV7ntZ9LNOUY4aVrRYonIV2cVmpBYJf/Rq0QdRx
J0tacGLx7s8n/RPSJdVTtjr2AJmRFG24o1dmlB4sUA0FEacqzli/Oawmgo6k
4hNrBn9ksJghZ4gc2uDah5HyUFXuupokYZFbGNm+WhVOiDL6Mn2pg0ZKpW3m
FbA+w4JLI0TJNc3mBnJAVXaLktPVX0ODiV3+gdO4S9zik9lrBh6JLsTGrpOZ
q+EFRchjaJN8xlI0nOrleToO6kUjK581SbCEWeNMSB6b0pXkMNAS/DdpRpD5
rqHIqwuAN/kGMaE2Vu2aRx5wMEuyndT8agRhwVz9zSk8UId9YtkOyFYr06Nv
52azoxASVuyLqX90IV5tPRNqVUuUp1vAym9CamKV6sFxdDGONsa8g70GZ75k
HHWWVsVYgyk4b9zBuijfgaforcOaVmdY0HRCkoCCiEelw/ITeeK2C7cQjBOr
TISk0FEyOqzQ+zAvwdG+2RnNWVhZ/ovWv1lT6XAzr6szEYBD4lFoDIuBBf4i
MKfOsTrUkt3kmBM1dbj/yMKohXq63ue/vKK+j5YlXk83730WGMRSoLu5m4Jb
KoqDdag4v7zGPQVOYJB0tFEQbV3YKw+dm9xXVTtUVsLQ+XvlMn/2G3MvbSbb
odHtb2e8W5i7BTvTuMKLuFbfp1Jevm104NH4ZlozpMiQPw9MCYrNAemejtZC
Wh5pt9lwbD8mfG8srpWeVMefkobH1Gis7nwJotl6uH90H9tBzyfAUbwWc52A
dtQjEd6gU6P3gFHBzhDvHbkwWyKgOSIdHSJYVEe7ex6fZrkzEXMpfkeYV4fV
oomvMymFB8j7uT8m9NxBqMJDcv7+rg6OO3kP0L2pFMNd9RWzZb3VGidolbRe
qOGrA9ZqdlocejzMb3t1ZWiUXa4bT14w5YzpKg4Q0XppMbwyeOKpSk0lKhSd
hns4/gC75GigF2HuMZYxtf4R90o2Dv379iIFG1o/uGdASvoIyBvXyTLk0eb2
OnH93+7DR9DyIlNYa/Y73HNV71jmLhfogzHqbYfKGnLpzpWarAIBeLxXOcDC
oYUmLfJum5tqc4HD4MtkdABsAoCDW+gnRvdICVsZ0kQ9fDD+s27EX6BTwvqf
Gfq1MHRazrSOtLjYtmU46+bsO5M9siSiPv3ve3uB5VDLGENqdCJ7hcFdhydX
vNLmnLCL+eVhdbhKhz8CcXN9QDtHuWF0dlHse47MkAIHu7CngMDHFcEIqNFT
Er99QT2rYiWHFLGog29IRrK/dC7qaee/a/roZCIeNg4Vg957/uZeNXhNfK/A
vwCZF65tOqQ1AhHzBRwohUid8ZscT6VBCadiE2U+jtvItcvsjzZNlxEYs54m
SYVkjrmFtKqv6Nv4IbMIHdcJKFil45wPX2QFxv1So6K7vUXKhXh8Ncac+232
l3zNNqobwz/r/cu78x5+ly3Gvzib8esp0Oip4HHJyNr8y1eFuyygSYllVd0v
QmlcuQ+yAlLTMWYpVfwGXblEel3tO8TOnx++9ZhPiw+k0guh93UTULQYCnI7
zgVHnYboff2LXhQth2MV+2V3vonwIiH7hoxfkF8khC2tlOWDwtzOkMjJ1rWW
T+NlTIP8WqrH0SCQqoMLW3TNG+lJyWZvdQCJvKCDf3JPKR83zntqceefvckN
aM5AeXllsU2bkUVH1EQWzqAaFJxINtgjML60lCqROelaCz43x4rAv7VPpqwW
JuVq/mDxo3+kULFvCNmvo3FAzAi7WUipc8aUOa7eBI/ezE4Ws722/ClbK0VN
6bn2aGSXGAwqgh24YJVexEU8RGMGcJL6KKdhn22iMVHqu1adqHygsJwg04GE
TSBTx+Gp1M8a2cBufmyjLJXiZYQ5Dd5T+qj6IvAv4taasyrnfL/LuAc0tCQX
cIzzFv9zsKSNHlSJOcsgZJTmkcktGgzfzWVNZWh+871hzEnz60d4McDJDDON
N/29MMyl7VSxAMBvEJqO3idHFMN1PXN/12fqYdviLwXVVWR2ptgP4+x9ZKFz
cXNiqusObhequw1lz3YGakrTf5HwU+5m+gteyhSC9YskErswll/+Z+1Xqr/V
LdkgcaH0PVEOyeGdL8J4lHUjtVGqsanChHyWutEIt6gK0KiVrlvSHpRJLTJp
oGbNQiIa0i0Uc+xjM3kKwqQ0u6c1bGyYjKg093LiSJV+XNrXLrF9eeLk7v2+
OkMHbB3FUnLlfJNEe3pDOvTGf2Am73cfFx9j7QcJ7aKOoAzk7rkdHVyYxx/E
7d3YMxoESiuQ76MtJy9bwVXXj1DnSr8JHUq/1foMiYJmS6fYyAFJzUIEHWy5
94TdRtP+97eXKBxql9yfEg9ahzEuScV1Vns2KduTwsk0+Jq2jyvhg7KsRjAM
k9Ojt46pptZWk0KoComhqjDP/ZF1F5L7i9jg9sGl2slT71bw3vv0CxccIffK
3BwbImoRspvV0n4b27UlJCp/dy+fOPYJ0QolF6RCRZmOXwWS3V65j78ShHIW
34+VFv4wjPlrFrbhfq7SDBSYvkZXv/BKZ5n7GWnu/dGpdk8CKwGPK1LgqxQH
/nzYShgR31GUpvaTOe8ATdgvB2gMMObpvLfTaGtCdNdwxUgBqYh1M246ZRdE
E4EjNbaDfBsiChWV1hChSKm51DZTfMKQc2Np5LizH6ExhmIVNvAUTgnd63zU
CcocFsc5LkO5W+h0cSDoWJRqfHUOqf7G6y9jgNnGmN9Dh1s9nzk8HBCWHJU+
eg1Kx34RyOED8KOfVHbhP+N7e/0DJUWLu05n4aSPpZME6KEgvmd0+/2ZUFtO
H1HAIZ3GsHsKiRJJW34SEDnJqB76GP2jOhTp5qUBMc8caADMMt6oBF5uqm16
7ue+ABRwnDnoDPv7458bddZpa+y9CDFMYmeavrnlbO5WhAPSDtSlw2jlXgKZ
AvPPRE/tPEl4O5D2nH7dw/ApHwPVo98H29Fi3UcSIW7qebeSauQbCe2EGsRi
PuwzMOVvRnJhpZLv7BorAM2YRnmkzWtavwdJsPMiXS3aXe1m3Kt8a4oCT4As
nPexy+k6b3hzb3ylN06V1uSxJI02pEe5zVAcRvA6AQdbju4qRYnr0q3zriv8
24HVE+rEidJl4AdnZm7yv9+g2/JJG2V7D8qWs0EbhKHyxU92bhQAdTMSXq4O
IZXwWRKz/Ds/yfE9d/TYieNoWimsiFiPfVDX7X7jMs+o2adF7CxklXG6Dtde
XGaa1tHSvShNR+QXTFNMywXlK2KzpiaGWzja2J4bd/6qO61Ogm3oKU7AkprN
fDRBp7DP/HasKGoE1DppuLmSQSc/v4rd6xCEubtu6naQkRD7svKD2S1FzMNh
y3TMARdAmJ2MxF901Zf/AuubbrwXzX3nqpkRaLKh7y6qtB4j5MGEEeuZoQNr
xJwoXC+oIM+avX1Zs49U5jv8P4ydja5JyCj5cA9bU6um56/67iYwUuJ0X3kZ
orPusySDtNWUBwpO6KvMtgI63r/N+weIpVH5DLHwLQ9QMJF9WfKgjBv3INVE
I/dyHthT5+NbMcIqkIkDkWIPKQWFKMOOYEYfab205Bs3vvIK6GE0qwb2/6PE
P6s5DO3AsUq9snjoW6MjkaXv2k2CsZolore7tMeSTsu2TjisbxxZEFR6unDe
Roel67RdUQ3GNqe6nd46zan+1q2lYkvmFeZJat4zhjykgB4xbOgVzrUfIGl+
EfSykh2QREhaXTZGiCcMocp+uFheRG5/saz8fXN8+wvHrehVqShXRWONAU9h
HGaQ+/d1Tg+TFUZOq8eI8mqUcx2jXWfkHpcNXCxX3907enbgfwdhqZzKpi1L
Q5syz2o1IM0Ojl+gWbh/hlOYMDGXnmWj7CW87KlRIVT+wro8fwXxt5pPTwld
xxc6CzSRX3EZqK0cLQQ7j0jYrlE9g75FqbUoJzaDI38qlykFclXFSPmtQqV8
sjdl4nblg/VR+5nFv2mbS8revFioLn/sCXC9ium06BWgdsSL0N9gWogx11Ou
+REAVuqhRogxNs6Cv6CHl9KHMJjl0/Lt+FUgvNR2cCW47Pgy24BlCS91lEvY
w6zl4HERbSaO28sbdoJuaaLCUnHq3YO45cAIKg38L70aAsgXV2vcDD/VzBIO
KpDucZySSr1Gt2NXdlV6t0ed1uoD9nd11SL0ITYO/4erF3l/9Rm7oCBNYs14
FWmRfKCOnj/cn4mx/ExW9ET7zbKYDzMfXlBNa0V6YYfVL3KhU9d6VD1LiIHx
vzdnrYBMMb6gFpZI2s+AuSt2YvgnVEay01e4ktNV9+/RdmVWCnsuIfa+5RO8
G13vGPX/FUpiNXV/gLZCf4m22t1TZVJ1FJYBZ2TDlxGSU/aes+bIxkz8s4h5
Y0/74rbDWA3qEpb/s1tMJpmBrQKxTPUFjOdMjXMyrzILVdfw0H8TtKvJa30O
M1ICZ/W8j2oK5JvJP43FeWuCayF6Y4IOEUKfQMOOMv4FSUkY0cXb7E5gsvrW
cYqbAZtNGkqH4LuGETsCwqHGsHgJUda4FVJNLPh5eqC7UD1dgs3MA6L96U6E
uSaWKaiyaDCm0A195F8EkwKVd/9OYvpcFdp1ofY9MQGwwljwAEoOjmkTog6o
uX/55e0Nm2p/TMoEnxrrnqJVHSI4xqhGFqXOxqJiMngxUngnXs8+96sF2F2V
3QF/SjLaAntPMn3z/D/u1hy7gNZrMUrsy53V4Rjjtjupo30SH269faeix7vx
cHK82pXdEvhPo5tQRk4g6z6mVPI3ZJ+g0hl8EWSYHs9ClVLFLA1jTgM0FmRD
HBUCYT6X4OkxaZbB2eOnRGpuQg2AbJXMI7jMh6z0R3WjQFyuqQoQ3NaIEVZz
fqGEWW0mtFd/C9OhlfXSxmW2Wtk3VhYo60wKrdLRjx/K33gGfKSXDkKRa+zP
rfPOrObtilRM+hGxizsCA8RTaGxIxKy97Gcu0AbEKBQntsQ7wePsm6Xv2vYt
ywX8QTU7MXtTZED4lbkHkEO/k82+usEcpvNxcj7D7g3AgE6GRiug25ktbhhi
DI6d7RilI1tqgLDmSbGTMRGO80tj+tt7+PMnPF7fsycLDDHy1LI0TbfTM0nN
wOyPmA0TRM8ImDjP21HqJAA0ESPThUkxsSawNiHIgUNfc+RD2zNfLuWAbalI
d/fXlizxSh24wAGGkWxWvLl2fQPi9oCRx8RzNidGWbs6L14BS2hc9ab8l5TB
APujPJ8OSa+m4mjEV6w9FThQQV9iXGD6wSz1Bjlo7kdn0Z8xQZTLl03wAjde
Av7E5DoxcbGI/Pv0k9+aW/hBbkBpOJzUKg13FB8k7NxjzWvjM+xMKfv+Juzf
1+xtifI8PlEPOqAUX/MYmCXqkvQUXN0VZARK01VdEpo0pLLcuNMVfzeaD8ia
8hMTrH5IX328oUI5eTx+uJ+JZ832HpQH1SDzpAuWhPHy+qK6B3/2An1GVGQu
qNtrq0QwXFhLx18kxb3KGEBRrvwjX/ScGafGJu0yQ4gyMDK9sIFYt4bBCCNe
b4DuN2oeC980gDhDJO1JHFvGPGYZuRQULChrJ/fsoWXhKeNVJYI+k+8N7KY5
xHt+tmThbG3FNXQi1cU1kXBHKkff5XgrmTWEx4WqVfMzo+qECIV+n7POB/fd
+XCcEgDhv6bF2+SvLD3pOqIk7R53UOjC+POumjJk4iq5o/Z8UIByriwFiWoG
Dafw13MOe46nAllVq10TwgfOVFFBbU4XMRMPUhYgcT9ym9Z2xogB7QeYkdjQ
A5PZ0FYtorUAYvr1hS+NI3CFSVWOXrXgpxH2LXT4a/p6c/M04/qJUIrq1An+
FkRZOLJT7wBLlVOhyQdT1+sKLduqc7gFDU0lDYiehLTFG2U8fSwGCfV2w+e9
U4fTUM3GmtlfMsVtJzfKKJXWKDTll20HgacinQVkBPnZMBWY3bxQ/7Zz/ShA
T8jUUhoYaZlij+3arrqgDgLfYhkFdA2ycWkxndMjv2ikTDl8WOx6aQzjMvjL
ufiKcryjsATWK08VnSW0cJVVHN/Yhxyk34L2wijM/SuXpEGBW8eSPZpXc63O
QEttjqyXFCxdywoPSOGZ9AKsidZiXDvPEHxxxDe56TDFeC8w1qiS/friV0SX
Lp/MN4Tmt3/conaFEsptqKTCnYEZ6tVmtKKkU1MxKlusrELSXbB2DHOZ5xYH
+0Z0xE8fXNBijHuMWZCJ0ZGRiapln7j841yxVtXUNBvS1IXIk8yL5fLvErCR
GhpW8AaqXgwdTakkm5vjGrubxEKeemOI4Rq0A4R9Nc4dwTqCqfl6XZnp0IRP
vPz73+tfJUBHc+QVVfIMrqiPMXxcm5c5GGnhXt3Y5FxIkzC7BB/9VRuNUjLP
cg5xQGPuZZROfKihHp2etVgcz0VUa6lOmqXfwzB6ER+M2IO8ReAtUWcYXa6f
yWBWUm4cBEQAAENyWDQWS0rxqEEzZisTRMf9G34PpBi6MAQu3uHawd0uYmX3
B2yn+IHN20Ri1N8x+xX4SCfxf7e0lHXtVTvwmYHgrHbz3eu6a/4kdVMRHFMO
HzeZDDzPNQbHq++NJ6DiuNK1XQxgX8dT44ar34MPuFTh1a1GSxTPcZ+/GwJh
YqPO7WBybd8TgxRy0gQpIxNjduWNsGKt1xIOAcRa6gB++SLJsanx15NrnaNI
gYDCX7s5+HmkTCnEftlHZ6rRvdOpCdCIvUaVp3mo7zVObHg76uFB99gSdEur
MEQO6o9EyzaLyDbtoViM00TDeTq27N5C9cG546u8Llzrf2xHFF5TFKgpdk06
SVPzjbz9zj/ZgU/7gs5a9MHBK7Bp2YxfFe8mNA46d+B8gFVgFC5Ax3UM5XUj
jk3lUA0XnCqMXZ1VUp3V4umEHdAxpNCGHRVZymcYfKqYcLUnRZ2ODNDisnoG
/tkdeQgUrY38GotY6RY5LnYxy5+mb1PMCHFfWVn2xOxEQjn6A0MCJxccLjYU
QJ6344hQTPzXbfUkaQJ7SX8mcPs+lHCeWNWB5zsiUNpz6Y/3UtNlLxRHRrRD
fpmzky2+JKGUZybhFM6Hrh3n076fLPp+TXdjJQ45n8pPup4bgd2LpTtL5/IY
u2qTNhFLQ3m5cPWNZjw1z8JMgCo2w2bDoRGkqV4Xfo7+zqXWaRozmlYPrs/O
rzMvClAwcAtoiumdbHBQpmnI+KI+IJ8y6opegYy4hRpvB1M3NfG3nSPCo13Z
Izt4FQP+Cwvr+OWJSZoTV7DMEahqzNdESV0N09cyMQPQ0E/sGir47uOSJxcd
55BY3yE63rj5aCq30V95PNx4I48VmlxecovmWAIz2mLmT5rzyROOml0jKaUo
xziwYFp+I8Jo8CTTZ6aWVS9W5UMbU1qr5WZ6Io1xDAUrPumVR+tLWrtGvF9w
b03ePZ6/WFL8QHCKjfO+IYAAMcFFMYDs1o6NkfUor4+Y8wEugyZAB6mkupAx
KYFkBeuG3RIMnT5MbdRYO5irXjMnA43/gwuEX7XplBq9P8Eq5ybQveEFPPL5
APLdUwCZz1WZIe7AMKtZYytkqCAKuCij8pMIbNmFRDtL1G+DdIurxlOW7j1D
o1M1+AZm6SrWc2sh+WVqg3eWjVigms3SEC/jbE0pyHASODIZRjgbqtSHlmtu
/ObLqdgh/oCPkgzX9ZVlxWmhNSfYrH9Z7Das9KpEBwfPF+PWSstZnpS9TG66
tqMnn+aJGPkl3XExSz3ma15WH8CYf7zyals57KY53kZx/HzuPUsLti/1IY7z
Ia7MmQRcwFoBMnGLay64RzZfJRfE6NVDC0pPp4ZJJjkxSGbR2YSvLOmbW7hR
WULWHzHRJwMjCuQIUCMGV6RZGay7xKqhLDYd7Zym165Lg3thOnSFCmqH0tK0
SjZ8HKQiVXg4hSoKffWhNC94kUnElh3BGhFodpX7zAjOv8HKzplJSHacP6+n
2VC0/1i+yLFz/Wt6FsFb5zLZHYdGF2fIsVCCgnWWoFuXOVu++5fgAEaB5C6I
mOe5S70jF4pZx1iZhZ7GFM87w7eLtfuvxIWm8Hjk51ZLW0XHJARkAtR/3fwJ
sG10sf5yM3UdFO+TU7zhYbzn6vkdq9dNSYoIFb1ZVOBFPRYCF0+7bqsoazBc
yQUgps1dpU3hADw2hccOHgzmLDbCWAeJ2m2UGfU3E+U3BkyhH5iuRZEq30Ot
QZ2ORih5gR0W6XgxS8zKgizYFJFMjjK3OEXKTSOsLC03t3MD34OKrnoOjHOw
etAxZeRwm5dXA0zCLeCAkFRm9TTl8qVxXo0KYzi6gBh0tmtEvm9BPSIuKdPp
wZDkVt5ouC7JoniELSan5bdgljQI1WQmpPHgl9MWO8F9dBvAX8tj8V4bRGfh
3ricyi68U7loXnYtW9ks61o10C3KWdmB2KHJ6cf7FmfYHGkvjxePV96n4Y1n
21AyIZK2gNOBleHE84qmVue5UOKYDiIWVXdW0M2zC9Kjw9hvP2VngF2XQPb6
pUzGnHZdgVxyKuYSJKgSJrel5Za28isUALCVWydV57DJIRMzccS7ckXd9qkL
vr+kbvNtNJQ4WyqMMUlQUkPhe5QZ3cv6nvYMIFSxk7XRErjK8uJ9MM6eu9kV
ZFoDrebB7xEh+0qoX0Vgrnk63BJD7z0B2ov1UD9I4BWUgi/0r3U6YHVxjwlk
VYH8DhlOJX21+bWuGEBN3BIXSrygl+JMXg4kM4qY5gVB/Vz38CGWvvscaVN7
6L8PPz18HPLI22NI2FsE/Tt9gBkTMdvX5T2ozKCqUlHPS46XpUFR7wehX23Z
mWJxhOt6Ctx/sWwHVMuzzg9Q5R7q/6O5Vmy1NSf+FdJcqFOOMD+lsc0v/6yn
tHfEhdXTOGugEnQty3GDP7b2SxhUXy4crB0O+ZmQIw5Ktv/t1xotj/VxIuvA
KOkrgQ8MnuKzbL8Miyg2AOalzZCtzn08ADQLO+PQsWgSNFh0L4mrsnHQDypo
8W4bLZtusprUROM8VGT+McYqXKUyb1pI4BaQFGmrfzftdmHk7iA0W4mndJHH
3AW98pzaafcEfgybjTxpN4qfQK92ZkBvr0trAHFYwI8WxBYN1dom9sUuVlXr
JgCBBz9KTpNf2E+ruoKrt7OM4iMM1Acs+r47cObmmHRDGmXRfmNmh1zsIJsf
xD3nuAELhbOlCron18b84oQ3UVRCYIGN2o7Yr/yYTWAmzVkrjjbuzcCTs+ht
xTlcoRau5+5CaCH0mUDL8WoC61RUsAGd7CBDN83/eGcnJQE6lucacBG9Ga/r
KpqbEPz6tYPHEKvSqPI7aVzr8Vl40Hl8KTyYtuwQaUOp6DJy77/xScLbW4vc
zBMQ44+/sTaJzPr4Qoy6iGaw3gItw078rxS86JNvIKEl0q+LPUZEGvJzVLWT
M6+H1voU1RTFlLR9vpobZD524i6f14ksO7UwOy5w8ZvdsLXWEoBYNb/dugA2
nhKeFkeQp+K08mPizkNbtxfkaxYX0lWWfxIN18UYLZ259oKEP8RpxZFlzUz0
vfE+e5rrQo1i2VA5d28cFtv8s1skCIasP8HkMKqt5m9B5B+wFvNzOPPVa8YG
QrxRVc5NqjH6hH5uQAwL/oBMNuxrtjmgVTIqimFFv/jtPInFoG7d0InUoWS/
Z0VMq5ojDpuicNNERIyJX0Uz75XVrK1I9UohtOrlGaAmXz/qQTFKYp7wnRT7
1z7YvSN/XdkaVkLx9HEttLSLjccYAyYUVtp7+AyW2J8/tHyIxzkjOa0qUa1k
gYjdZXq/hKlFEeXOaoGBO27iGbizLJJpONBo0m2a+Z6nVYA464K+WnnBTp+W
fmgebq4XrwFscdHHhVXIyOk9nq+fXFvyKb6fZ0SUv+M9PVAWgoCwIryvddkK
jIhxfd1QbMp1OUqQoFnBVt0epngCawXBVxvROBLMH2PGrBNJ+Uotm3vtmV6v
LPeZrTcEnhvfDyFGDo3vF36AFzzv0DPHOvedJXqQW4nn7kkUixBC5va5Fj6T
iIvj0jsJxHTuTDGA4t9K4hJvPb0X8ksFtgDSwJ3Hu31hFNPGoeP226qZBDuW
9ZWwKQK5UL5DYDvTwkRtTQsLN8AyX1eGKIOSBDDqmzZ8EilTAasKRZbqUkmj
pbKC+OhSqDIYdoFL3vTbu8FxH6olqSP74Z0ehU8szBL35kCmOkVo7Cjiheja
0ZAd15IOuJNy3TwAgoEmpMgBrZf2tu9rNjV/K3wtK58U44B4p2qgpHZA8S4D
PYjeQ5KSTRQIl9d1SaK9eXbvMoXLL5o4nSUYqBP8JTRX0TcbpLhcpE6U4o1L
ouJHX4Bk1bwKhMJCce9XkAPdiY64z9njeupJPKZS4iRi1uLIzxURfKocXrPy
0ygxDe0ysyV6gaStLgG+Dvno96OmXI0TT0/scwUaPjoSA7evnRCU3TUad7QO
59GaxO51XRA8FqvP7j8TlgyMrq09taU/FURwf7/yA6aVgBY96tdIXb8wVXOq
fhsaQncam3IjQfCc/vXtNmpLSydClk85CLKZRlOTQIZE7SrG99aCgla5cC3O
sFdWlbNkydIot75+Kn3/yMXQhhJ1n6uloJqW3nqd64oXXk/NmD0vSUO4wsJm
gk4RSzhvFw6XbcDAghE9pKcl+mI4YRZDaDv4ki0kWJwkXIwoJBWqEzMbYDCm
SkeA0f5eP+CK9ztL80kYNEGIMBPykNudc7M+x7s21oDHXG7g8gUITCiiQTJa
LlSO5fKf6XgUbHEwOozUeGCZIl6+eGz19DfC8Qjvwn5hL1DwChHn5Y99MxCb
HfNuS3bH8kdpOSPKPMXV4a0hxNhkHzgzwucGCPwEQCs0c0q8idVtP36MKE/O
/LHpWagoj/NiG7yh/QAj3MiFqu1iSStKx2IGFJXxGhQ7OTMPi8b//s7/WjD5
LLvDLv9VWXdQGb2raMpzgH9cmM7HiBx/I4T58MPsHV//AlYzuxNXmEY1GVge
S3cZbx7qtAURzCPkOt0JDbiKwvBp8SW7z3hWgUv5+zm82fajc7PSIJn6QcP0
/HB7jEvFGzUh5OblebOs9GZoBYbZpX6K8RsKn8RZcS6IFypq0nW729CxaUkz
OUGm8m1zE7wA0P2xOTBlkMBtLJ3WRcouF0fyGLyWeU/IepWwshJ2HQLT4Oml
PNT3s3yiO1vHH/d3eqUqE7rpyk2w/ZXv7ZM7iGP+33rJcHSwGlRZIDVI5FAR
JM/dzL43NI4/KKA8h+AhS3OYNnSuZYulV6pAPWsVMa03zN5omIcewG7QvW/Q
rb41VDsagTGHv38u0y8+Jo0l6r9Gjupq+RU7KZRWF8d5Xg6FpjeyhgEoFifK
Xayml1iCLxIlJCI9oYldbp48Rpe+60/jew6LA/93w/P6hze8r+3hljEKkF97
1ZxQAjF4MG+JX68KZKm5u34IArOD/CYYyi/MrLzCpcwf7oXSmg0PCE11vlPh
PcMa7wtf/0Cjdcg+KFhYBVLKxES+XC3bareGUz9rB9rTAX/M+2X6QaeoEfJ7
BQOuh44Fu1VSmxI2TglfVVg62n7KuPLCALxBJhQR8v6FQOW2Pa4lTq1tepym
AanjPedLpUGKQ2ujAaUYI1aN1oWQAlv0V5lBDHAG90Nw/wgdL0Tcgj+rxEYF
+CPcYGrcn9UUd7l7XKR9D9dvsy8lyUtqnMFx7M354pAb+yqm10rkgDVmcLMQ
9XBPxFo1mK5hPu4K7EHXX3jagb7HQTeRwgq3bgklRRoR87UBPXFCDvASTFER
i8EwUxDDZ44+H6l0GIiD0fpF/qapTI0FeFReMaQZwJEcABrmYaRYOaPXCz/0
IzRE3Yn8o+JjIskjeird/Zh9ZVU7B38CBAeOsL5j2LPOBRAp7g6dCn4EUuC8
V8NFMApcUjXBy3xuOhC+MqaQbLMx3C5GbVWxcmH35jUIMD5XW2MpLe5nVYUL
uz66IgTJDG4F6VEMsNmV5S+lpagFq8zEMySWDKZsbcrTlYjKJ4ZmhhjMWGvr
281hFKEaOx6tCmdA4V3f8FtTi/hk6lgeNx6brJMOKVrLAGsatFti3F5DjK1a
7yk5CD8asmTBmLF4kr9xbQnM0/L8b4LMW4gUE/ppqoQKdbbP+KY8FCLejHVw
jqFiFk+V32zE2bL9B2N4bt8CX7WLODbC6ov+cEPy0eOTCo89ANj0d1Onde23
mx5zAbOrxbHR6ND6sEo8byVXl/+FcSIhckXtz8iOwAYPbLnPAzAtv3vKkdTW
s/TtyNq8qz3hE5lubK1TbgEsj/4XVAKGVWVYPLgdeUdwYaXNhRpknXyjuUpj
PxYF54v4PG9AbVqln9K0pep5myvURlnzBQetxM6oKtS/4dTtiCvttOug9wMl
KUMdzsMVvem5qiDEFwb0PvLzHTZFLEKkuzvf222lO4cI7LX2fn3HYcPW8XrA
2PFJ37eXdQLFNHgsJRGWO10pmM+LasUghdD2aHXOp6ervGmNtlRkOQ4S5W7K
zfyAYcS++LsvjBblD0JN5R6jbUSqYqKY9EPUpsJyb0ADcgUva7jdyl+2oUwa
LOtR8rvct1B+e/Ktgn0THF5de6aAGjq1rePSn9YzetoXGYNWq72fIbFyrHYw
wS7o7mQ9a3siip/U06qVlUewmoCBHq3uBQkrVKF6/fkqYd2D3qY7EIKHmQ/M
y7NupZmRdkRdYW/m1PIMH+CF9mRKDKFP4C/iYJhtd0P3aGpATxQTmOpf8ogt
N40oM+eP6Y171HVi3qfw3eKvO/kRWRaN1UKXBtXCJn8IgqlMsfR6/7QSP3ls
iaJID5izyjTOrFilhTpdhenc5pIbCs1r303MtfLkeY1TZ50ub2sYWGqqoMHx
BM/MQi1erKwxy3wJ71sQE1ATRgtwftdoilGoppknvpQg62Rb/k2+TxnxN+B5
VvZlNVluZiFJVCmA0OTDTQYpNMFJWsqOy5VuHSKH6Z602tbOcTsE5UyDHfos
rJDxL9f57XCEnIGnGTbvE8ZnAtcFkP1Vo5NszZtW7AXcJUr3XxwlMGRE8Xx+
nPl37/8sQyHyKyPTeiSiyMQV1ZoBj4N4tSLpdT72eSaw7W4H636tmq/FSn7s
xfAmNqrmYEWb4VCWqTiR3oD2UURGwmrfnwemmU7dgj0toTxUTXMkeqe4U839
UEO3jDziDK8JWdo3lOTnThqMN7j19DZiWQIv2lwAlcBiXM/iXfr7zFbSSDNu
tLv+xUn2psYTTD9IPB60gOV0v2N9LIkimkWEiiHCT/CuKfxlFvDCy6mH0dbi
v+iT975518SostqCJzjjfZRkagRvIOv6Xp0VumSnK7JvFeh/lUpXX4959AHz
6mwiKUvKep+L/adYPZlDkXk69Wf1yizuq/cbBElK725hMHnrNZ8S354LNRn0
Ud7kBe4D486HSZgWpxlXiq99BdJRBi/z+LrFpXHKIUb5VhRSBOD54RIiZ4HG
M+7RLhb49oTg7eMJKYJKZa7c6rdCSLP7ObDSk3cQKi6uuXUEXD6ITeYHQB9/
WiwgC2eX5x3Q2KC8pIePtjmMARzL7dIrwzb7Cvf5htDxC6v964jLdWLQFYh/
GxGLBhUjSkE7nUy3ibcFyNorvQGuJj4gSUbZidZFsSl0nUYw5H6RTCUqP2Cs
goev/jXzVFell5flpqKFRkQnmM+t6QMrlfqX0FiZ+OBeeYd14ppyxfHLB6iq
Nb+fbK63ujtgR85r2IQETpluZ8xMclw5N5tLHTRQdztLm/rgxN38NwLuung8
6M8j8acjTAKiWbk8x0IkzraaP0/ULAcIkdWEZu9L+P1oPLat/6y6zm0mDAsh
ETKg2u++TFiiBm2+87TitPkj5XvqwMgrEJ2v5THfHwgKtwiDJkzo/5D6jYfS
PnYLIKKB+kD9/oJt0N2hmHt2Kfsd32xCiPa3wmYAPlpmiWMJhttxIvxmfgG8
EztyWq+2e5bdp26viriYXeNREiX8TMGqv4UDY3bdyKPPtCHeEVLcMAf7nN1K
btodD/Jx33RUtN1y2aSvCIIPCYbjQGQGrBBRfQ3Ez5+lwhaCs8tune2qrbw4
5Incw4oJAIWnJxcumomWouiJtcjieVw98x56XcQp8CpHrWS6qSpsbStAs1zk
wGO0ucA3xm/OzZpHM3XxUjHZWraxyogTE7c/BWF176TxMXWU1O1BgAIp12aA
JC+0cLS8SQVeZ5mbe3Lo2I7I37ZlBvyjjNIdPizM8WSLZBy2zHfzSWY/2rfB
GSrB6J4CfYMIPOMdYD/yU/ClZb8Wbc9fh/+MndO5qaSvVgp/cJ/eKVHoaGBy
Dv+yG6kWaPsnsBt67XszxXGCMU0YiiVA5oxvFkVTPtWF47G9DBVhgPSjseMd
FnElq3fcq2U74wOyjb2OPmhHIqJFqqZxfqNvcJPtYyMtPjs0/opZsHjQfqL1
Ry2quHhldAkqqfHdyD0PqaqRTFmdOP8c4tmn8UsELg2ZCpYdMgJJng3uC6zM
1WHjr66uw0/xwMGZ4Po4Lewo9Pb8k1r9673k6tvJnpzH038kf7swz/wnWd0o
pRuobXLSFEnmcDKt83yC0iSYM1krDvpQwGbGdnO1WOPllFcxERqrnn7LmEdA
cvyEPUDvDfQkBnP0a6f6Y1m8el5wg+jt8BJxGc1LFMSuMJ3d+US6hjrhhHCD
wXR8ZT1C4rHSjEMNEAiaYkVBOtPGYgI9fV0bY8v7K7SE1+zcQa1Sjt41ONad
Cud6jyJP2acPfO8hq84u1kFLyqUo0E5/SvY6PpoIZMmAT4WFVSWr2byYtE4z
1hDcN1bWTBAEWjuo93XHCneHCb07nwmGyHbjc9i7ZXqjBoRXG+51X2RKfcUN
bzIYdSJ97h2LGFISkq96iS/EVF6rb50bFXXKF+2nNZffLjx0RQ+hMmxHF99A
9aj6i8VifLh3kqJNdA0nvsDeeR+aGvl6FSuENYU0RZW6LRIcAWfdyT4i35Wf
VyTev/RG4W10hMgcscWBEuRaNqUBjDnU7iCxAq2WQMvImijUvKF05Lof+aP7
VwIoNssC1Y2m2GyqIy2NJQ6sVNwdZA14qEGubP1wnofN0thVF6pWBCcE2Mb6
rnFLIt1yqaIcpgS8tvdE9bNBFF33fJiiCD5k24KEKFrE24luI351wMQbvKg9
TmttEJbYBik7YurJDCFYjPf6ou//Igbxd0c3MLEhD2xM5qU7zqcOmzpe/J5P
HlCwSX1dbC36AIsK+MXpz+3aggB26gu46WUKkZ1RmAJU2I3/LJpdWabOx65B
+IgVeSQuHXPFPBsBya63G7Z0pUj2Tp85sEQ924bs6TQWDMTHoztKP3BMXD8o
7Y06/ZSCSeI4/biIwQo0DwOcNO703bzky78qwU5CA7GlepqfhWU05NImR4cD
uYO0SjnrONHJ3BEjSzvVSXO+CHhhIH7vSuSaURKpdBCClD0z+Ot+fW+W237t
ALNbD7jmvZFraEO5RqCk/T1HXo3+hyM3KVorBxJCc3kj5RRQwJ0CzPRT995N
Sg9SrIshjjZXViRVEaTU2+auSxLlA6I+DMlPy76J0P1LDeC3ILOsrN+V7PyD
tBN32ANMkieV3k+G64fnQ1qtLud3jejJJgWQ9QdFm0N9JoxGD7hk0lO7cmxC
QpW7yl3+1qXdKYFNtecwY1grJzyYTZh5q5gMf0Fr+ImWftM6cD1TSfSSk8Ap
SUxWLVFfOz55VqULYXhyiSCRKA7fhcE2FwzbS/N7AURA8HrF3uuuchbO7U7U
2ODu889FVyu7xkw0x6v02Sr/oeBxtQY+nxgfuzTM/HbTm86vfYku1/2Xw8KU
w/hdVk4sxLhhr/F1upurK3Qln6bXJIhYGUL2hXPIijVHf9aNsLBpHPi8KCPY
0wElNv8TnBu5pavBsxmNuATXF3715WG1SymbcYkPvjhHUE1aVPcMljTW1krU
85NfKZ+O/yjqRig2dEtz5JRSn3bNIlbhYMR7v5GrmmpT9bsKgWTwIdCLY5yd
0HPeDGrSlD8ZstCCp0yNgcQJkBsHc+ezWBO/qGEis91WtSbgJce1kS5ByXrn
fSSkv6Qr5WYcqieSs3BWtETxs1pgoWshZ9poOodLUGURdq7+qW6RrcjIjbAv
xV9r3h2fPdImGDtJ8RJ9MeTBdqSSqGhvdtXpkkKWakaBf6MPeQCTLIKi+qoU
xrQsEBzmVgWesVeMsJncOOPC1V1IIN7Zd6vuQ/aEI390nK1xMggH2qLbbtAJ
o2cr8AL5sFNZV++Z20x+CrwBQEDk1qIGiC9zeqYDkJInHZtvKwZizzfsjS9T
NsS9ZHnFqkEoZ5OLX/69TMIF4A0TM+uVQ5GyF75Cpn//UpFfoBk1tOhgbsMx
y2r0dauT9FDZoNLiZbW+95lIwO+3AJ/x2pnqHKlPcLR53xjapMvZtYY7gFlw
Uftm1DTUJj0zOm5/qLkzGrbbLmJN47RBC+YTx45vL2V+00Yu+GBZW1kGQF7/
ycNbUaQL1omv/suJLfwpTFNgg8FLfRwn6v65vpOFu1CCt3+I91G2ma81L/rA
Zxt9ltleYM/VKRp4kmZ1ZYrLOksB2E/VZTFsNOphZ4fdvZPHmF4nyEiid18a
JKa86tzbh9AyW0rcG1ykwkQxXq64VV19l0M1luAkAtljldK8N0kpW/vgoz3D
cPPL8AusOKF4e6QLjCC1FwrzI5Xxxm5zyXn9KPJ71iI+DtC4+uEU3C2ZSrD4
QcPWLkzTxJOcvyiPSyd4MUVoIr8h2gzUcEIspypGj8a7PD/dx2z2bVS6zWT3
F2NU9h/Qt/L59pUOf0NyuuEVhQDpOWeVLG5Ohxv/tL6e4wK180Ro34tIcoca
32CATMisXTrUOFwr+CsPpo/YTxBx9Gk1lLbt0NHryN2QZu1l+oWa4pUYvg3b
EzS/L8rKQyJ76BUhuj/fNtM9Dzjo7wJJHElKyWMUgJ4XsLtsi3Wzjbe1Nh68
ZYhvrbLL97ufqPziEkP/LxuNLNRBfPGpi6X28pyt+qFSWH4pRmHv6vd570YF
gtljZ0ia9E5aksdyrR9FVAc1UGNF/6o2LeITd3KGrDnBF4AC05jbaxKKv7QA
eVCRwvmw9UsieCKXtGK1+V+sevnMmvT0kBeXbfzRcWXK+ENcesYB0SBHuSWO
UIfxEvy5dgmH4drpTRVPQ0NEJWFwmDtvxkXGfuJ+XD7zXaJ7CRS+rQd8z1HL
r7A8ZMB3VkhuunyPvHPTMWQzJXABgskAM9osw/WcfiBae8ltX/kW1Xi8uH6o
+WaTmAeKo+mFxNymeV3TCHDH4e/X/Xr4uUdb/Z9nM1pnLX84svjwd5gOK525
OqCENzY3WPCjVkuIgC7XuEv/TsgPHVWQvMvKpvk0y1wNGUMl9CdWgse8IKVQ
PK+RyjuywzUjxu8lJ5MBzGvZHqpkDFmr8/eVIQnmzGyeH0Kq25W+UvL3Zfwg
9n4+VmxmhhxHgI+7SBpYwEzLbT+jk2q5iq33Fdnny+1didPR89eUnnulcOT6
7Xxy/8HGmSjsAULLKw1OXnOPc3RW+ciI0V201dXpDgdmbzmsuORpOfiBPiI4
iMKpP0T0EufbULFHh7BA3HFv7YFTtSW9e4kzjI6aM+Iqnimmwn8V476IxfcV
IqvPsyhDuT/csWxry+/EcXND29+DVgXbxuwi4sR2GLQqbpxcj23OIcn0CZ2W
Ch7RdVqXWoGbNxJxko+pIYj+7DzuV281dL3Hu22hoVPAaNxsl5uuiV99z6qq
Q8wTvlun4NR1JnXfImuQTdmWSyegKCG2y+EbFoQUvYmtsqfSiT4bXQQdFsgO
njorG5iTeIxyRjodZ9XcHjARXeTv2uhdVcOe6M9+nLkZgcR2KAdB8GhTbrts
+a7VQVIFEWoiR4i5J/eap7eA8mjjSHR7Qg/Cn4r8rsIgltTsq2HIiezbKjkI
q5S8MHE7R+I5Lzz7TJJICV049XAbdg44aPrXDwV379P1RuemxDKk9Z/B3nFF
KPT31UK776VoksSMstlGksanaGK32HKLJAD3Btf9bsFFp7jt9nkkyPy1cErv
G7meS11Nr+FyM/+2HG7+3Qw1rZA/iBWfSF3QGJxPmIPcR/+74x8fF7Y9Ltmb
FnvYj0INDXnQyGq0rOpFIwVjGJa7Q6MJx6r3RC9UgLJv6UEk2SvGAMgBVTfN
SiUqUqY6r2ffipHFFIaYVNbOtbOKExCriJUc+LkAiSudlL+Pqycm4+pl3PWP
HKka7Ihh6muBiNLq2iGz3cvncLFGhORx1QT/EKHa9MwiA4axLuC9/u541A5R
siDdqg5v6UqGeeGJ4c/PVYqcLgPBcpGpKyVSqIMtwwOu7RdjbDaiAtKiFa8H
NTOeTe/PvdagatWwyf5UaKz75A4tLwe1I4JhGM3m+g8oJn/F8w4BdCuF7+Am
5cALqaUK7OFsPo9TNw4ew+EdrNo5ktBioT2IkCm33tmrbxFvEQIVX9llmRVd
Nzj9Zpj0EUu4WzgprnCuUZrXOjgyCtYcROZX3pxXN9C4Gsr426wzYDIguVJQ
+KukNmQCJ898wbXtOfb7RCIQWMZgxe2TSYdv0f2I584ZdmgcIHG1OrilMEjU
7srVeGfJe8Uz0GS2yebpluP6dbMyK29VjrMAHhkut8hZhCWdWS6I3u1Giwop
qXWSfpm5jEIDVUxbbMbZ3q5qMOcVXFVO8UHyTR5Fk1WzYMOrTftSQJmUyts4
edxJaYGsjTL06UF0Aw1MPxw6Ns+W85B4nAXyseDQTmfFSLxNRoPlS+yngaVN
ASij27MVirVxdVwBK7lag2VZcRql+BNEVirZOvPGSvNbTYYO6jK8CDV8iTJr
vetf7vxZKsAsvrGqAkhyiL328H7vux7jnNN6Ucqfhz5f3/GCg0EOZv1pklLw
svAGAGFWtf+hi0Ej3qksp/uv2F/9x65vC+gt/yla0HIYSx2XIbA/dznpeCsc
zCxVkkSmQTC8nGmb0g9zO+RSd0yspwSgOa2yn3xjCLbSlYPyMaCn2t5DFDYn
1LznDoZREMmjeJr3+cnLWsCcBYFZL0h47aJiyzypAik8KLZ8li2YChg1n3Jn
/2BCogt2DQO3SBF3xi11YqsnYrmU49mbCJsK+wTJyA80hITGvo54gyyKLEBu
kvYjRalfjupi/6DZrNog1gxyeIbU9fbsKnyu/d0hZfHpNLWLfYQpmE/+A+uM
7zUV5IRGEE8UxI5KUrihuVJeDU0w+ROJQu5CiUvBhIppwF4W06xqgDYDeitY
vptI2DJ9TWzCJ0e5+I5LcGOj+Mj6LOTJ+b7L24vNDb5WwgYe+BQmCNm2SfUi
9pGATuvGR0LQPHzQ/Gue0U3v0xm37FWoYiIg4b6d5026+OqoOcVhVK8cB63O
VEuK00BO3an1tgT5v3DMtr1PHjmfeHSH8yKsdIJfr0Za/S+G7WJ9acv0hgWX
bN5grUoWhUFC+1gUCxcaQrFvLbWEXZmgPBefMe8au9+dDjo6AvvT6DbZwISt
EbBO+z0t+PiCmTiCfd6eiQWtL1nsuoy8gCsmTdARVEJNyBNav6tVMOv6Fvb2
cWBO4rb/yHv66BBGugpFcHNWE+ehlgE4IQI27ddSY4R2Q5H4jchf2LV2Equm
mfnbzEJWYHuCSEC04y1z2NqiCq2rTn7eY9A7qytx6uw1EgHQd9V/WYy5n+uE
yPo4jcJSWcMooB1EQqeDoAzjg/nynoVOVIIvuNwkX1T+/hl/uZ07nPZAiAAo
xSiA0wXfMRFLGk0nvDIhif78o0/z4AaTZdeQ69oSBFQ3HtNkmYaYLaC2K7zV
FG+ZQmpVaYpjZZ5QEMw11sU/6E9ADK5a/UNJ00rPXF6sb+tqwORjDelJlWwd
CnHkve3TH3AmGkAyJ+JQh3VP3hildnTGM4DMFfYgveTj3d+XBIautFmqmsG9
Siv5AsOCXpGy34G0CYL/0+ND6riQ+jtngx8RF2Z4Jml89EcC4fhZTj1WRk4V
GuEegDUTrCRLF/XFQlPZPdcFJk5UVwiDUzwcLuylukGtX3r9c1KYZQMaskmg
uV/SBZrxKkvniErRASw9cOdPiR5a1W5qnFpYzAE/BEZAs+123Fi21sGpeIku
gf3q/jBgnkV/ie/F3/tZGWG9RXuyN53XnCTXGhPx2yD+Lmov9vEiyoa5yWGv
8Eq+eveOaYRqX3xpvefueGVyjdGw7desKO4qGYzkz8h1ZY6CuWES8YB7qZtR
Bn6q1xZsWH7BPq6wy7oaZkNiLpUB45DzXI0PZNfHE/yHaCxMusmieiQY6ueU
zycmpW6AED4TwDSl5UHvUY0QbQ5/RwGxj6KHU7UcpQMKq4ArQR3JYWLBKLob
yW/nfP5f4GNE8872lQLTeLMYKYZe0bKPoGJQcCLjpV6moUKMMc0/KvQ8Zhkf
FFEOovIaDDIkivVOwEDbBqElK6VGz7KOB8VkfkGp6Enjjj8rnxVlgdvjj+68
GO00uCklHfZSrwPBropA0IGT6aw8Jo0OER1O1E6f45kduYXk4uzp21nGIQ1h
d9g34CLmP/vkqs+L/FGA/9DUgO5ag/BxKtwVVooq7HQpGqux4H/3jNk3EoKt
PT4sZZ3S7lCDapDPI1qFafCXjov1gLhRyvQZ/nqiFETIOq3Fowbk4J1myo44
rC9HOChc9wZGf0W1AYI4DTAB3kTULZarqroBu1+8ABeesDESrsB3YD2qQnv6
97OrCbdiMW+TrX/cR4Jo8ngiy3gdrRwJ6fS4TbU5yiuyWnYEGBwRJxUOe6wr
zSISKFy/HV81hxYJp0GZMEtmUFFUZBM26cdCQAqAGtbl8NXMjx9nRnnwh+ZJ
aS0mlWaPlBQ89ICSKEdSW2C+aQih4xYiTZo5pTCuxogRdAgNROW8u8If0JB6
DEQ2BOtT2dr7wAWNE4P+f1CYp6weNx8zUMf4vYiVwvNUm5wGMTn18a5y2M8S
J0E+JPuiW4D0WRyS0nPtKJjUlVmNNpHFvRhoJ8EnFgRnuqTNJA2//07cQm2A
IZFpyLBdvDKK/mrvOoagpS2el5ZgSEPm4CY9dFgbze6bA/PwL52cEqCbcoaD
5SSN0Gr/poTS/hRnDTI0jGjp6oWBZgE+P5ANZch/OtG34qtT5HmvQMQRaOv9
XpCSI2Ohjq1/QAv7pY3S1RZCE1imkqD+YGQEc82xyz3dLcjnINBm8zQGzUST
Hq7fhgEbjN+z7To8RH6c5isrDARyMYfTH0JRBiRYNJ3HXXRJlb2h1CTvM05m
bSjKzIUKYEYxtxc01JXc3CREJY28XghrDJP2fdcCZyiOb1BUizrW/UUK4FQf
9Uznq8r8mwZ0CzhSK1bT2MdPOqC8rF2NFWTORVyRHc4P/Dys4n4aYVwf2UZ6
V8TTMp2CTUChGmA0OMZQCmiAav62GpzGSzHAbpkL/wU4DIWQslYvwT1UELrL
cRorz7t0tWEFech5blchhMpVvcZ1f8zqa4t7gh3vesT5DckAbCMexXEly5sd
Jv/EPB3saZH6MrbFD/wfmBCqLpgZk70dx8nYRP+HoepLeG/pDvYgfr2Omw4J
qNSId36EMfCM6TY8u0SCfOAyFk3Np36fSUDYTbvydlg0poy24aqBreon82Lf
3aj0lQ+ThOiqkk8IdJy8YxfCzYUMyO8M2z7ozOrDzevXkaapGsz8cWkqoUlZ
+quRQZf9k/Yxc1aMzyuL1lDIeOCyPglPFdB7QbJJwxN9A4+VN3+sGDyqFR6m
lFUPiOvoUZSjF06asY3R0MeahjtqWeuwXLiailEGM4XPPQC7lMw3vngzl74A
wKyXqOFR94Fy0QDI09rPmUDkdpmXJHYTkohVRMLuVc2hoB2n9lgk2/Z/l/kD
FCrSZtiJN/GmLbDUefVa+E63ux3+Q6N3pJj9DBnnn02AqPHM/8KxBIhoEHqu
nZCu5b6qJAYAlHl/08a3YdMxOGroS6qbbDWwJaRqM+eEEM+IT4DxaiTBLx6k
uANSsLtFRBqgwWPqgx6rNoDb0NFbbUIlMXRu5a73Y28bTacISpk08iRfHo6F
d4YSDrBgn7ti37ZsMPxx8lFBXRh+IUi8+0Z282i/gbv080ooh2fwK7ZSOrcY
0rW6tkIki9zfnm8n525ktgjv5OVagiUKoKWB/5AKmJgt6AV3v+yZ4KxU8qhV
wjrlqAA3oiZJjTWfuWYHBYPYuv0aUWb8p64XZc4PdWzPiWWC7zxvkGQVMETS
g9xXp43wiz8RI+vXhjboWJL6ZRHw/gaYJBXtuDeRNFOzmJb01g3eARbRRhOx
Csi7aRvRoCaVjseV49g7h9IPTx9X8TW7xDQ5UhOBtIHFjPHuMdpzZRtztZVa
ftpvL/dlHHalFWJIyenIO/JqRv3IPVfIVu/IhwgWbDL5YDA/8cPjMap7FnC+
SkxY4to1DrZpDOKb6GLys4tOFCfqe49qlS5GzXL+SG7aK14K57HsTnjwgQUO
jEXYIXAQWTVImksLmh17a0a66RICoOcdxelvElMxRZMe8ZLv8Zpy6zvcr/gv
fOY7ba83x5ZANlus/KkXT3KvVo+MYpxXMcgZYCn5e/DgtHgEJahJhNwxvKAs
5ppOdCFx5PVJLbpy+r4AxiRvCcEkGlsDNArS7MULT0bJ8rmi0kGa67xgp1uj
FrRsV/ecLqF+rv6nSXG8zhWndMz3G+e4Jdh8VfVExJJeLj5XR7Hq8VAL0xNL
Rzps9G1RunB1ZuXK306LDoBtCR38ll1sPb14pH8JRVedlm4YMiSisB+/sF/J
ndtjaFMOQyRNwmhOB2tZJuV0tXC3LdGMpI+DDZpR97lDr8U4n6QPm8La4UP9
qUQSmaj153mVISbEKvaRiuQr9FhmElaP6Xcn5uhegof4EuCUDvwoui3UOIaK
Dj6rPWzMDftPcAydWe8W85aKRLVIFe00LJ5jD3PyJxOxBXuSYn0WgBZfV7GE
1B5fz/b7C3kEjAVR/tFXZTrXrNyUPasSJ4c3fwoHXtExMVkxBAJ4Bws87DJK
QgDZJlYcA10eWS2frSL9ZlHrl/pEMk4f7us8dflVla5PWb4DzAhPBi0cBAWA
X6eTPJNRk4EQNP5DGCcO3j68+XK/vXfVSuVS6U+ldUjekVpqf2vhsPeOYoWD
3qAJIKsvwkmSrWvkkfmW9wMXzhJk/0H18EtWgpmiSMjpaDrgtKDz2cBtMdfc
BXLctB9oVkC1mF/xP1rPPkSuh7D9L1ZKF1oOscaMBGjdNUKjNap5+4d8axAC
MYsmTXCQiVPKwdld0rPWWMfy3lT2ttma/fTiqb6BikUEnxk23Va5RotP4jdA
LNragQVoLyQo8iiGQeRJ/oDzh6jPk3RbgmDkXBmENYEbeB3hfn5Wc+EleVap
Jil3gW/rUV7n2UfEaRcrXWkcybIU6DBMYtuVqXQPm89TtVZz/PBN1387350R
pqql5qMiGxHjUJ4s1uLXIQq4bMq4RONeQk65akdRuSW7+fnDdwiABwpD2x43
RZfd2NEv1/WfSZSu3JBIl6rA3hlOLxKWxSlj4ACkYuhGira/2RQLsZa9uvud
XTSthbdXOw0n3xcGJnXLqWM85X8Ei1riU+vunJXCE01kzm4az+2LM+uf8BnZ
1pplOE71zUuFjX1q3rgWEo36OadjUy0XvqcJpDfME6uDnGUlCGtG4D/vrj9x
VYmhR2s0KDngbkHBPJWfQuSNqFpPbKmfHX5XJkiFTlFlwDkRiUma1CcVqMF/
hiPhXJejzEqK0o5EYw3MujA23xbGuvXeJbln+32V2wR6H9IoMhrGCx5X3ZFL
dvkdno2ah3U9J0muCYn8VA581K4thCdTmtvdT++M5JGJP28kS/bT8Rmbfc/s
kFPiOWVatEGmf9HMORtRUt+7lRWp4uNum+r6AGdgK89m1onD73zePOlG8r9i
aGM/xO6g+N7kasatW23GBeSsILZjuC+Jqk3j8tMh5/CwR6guZhycBar5InJA
hcJ0ZcVvnQ71S9HP7fyqxCICeh1rmsftBdigLborXFBP4aZZGGgVQkNEYpJf
vp8vUe7c00kH98W/q3GjZXqq1U1jWznWyOt44kXqzUGOUUHWPh99k65HETwG
aoPp9ML50usvY13CR7aVkGVVGhPTMmaNAFPAQ2im7BXItdiYSgYnL2QgGf12
BGMXeKHrQ+zUuF0wqE0t0HSAsAJSaxCQ6nsPlL6RiOUM9QvSEOCiMXM7M0MA
qVsKVrgbz45786CU9MlYdoU/eZEJhr2tObuVT69SuaXN3ZzrU4sbfWfgyG8c
8s+IcYp10SA1brUbt9+ndjeWdlEstQ/+7keVfFTY8annc2CCukx6CqD25XJD
2ZwtP2I+4DewbHjQRsy/HTXeshDq3Fwpw4NnMrEMIwt1Odizm6z7eD2P3eqf
SUDqKXTmS2CrE9ymXOtqfPXkO7tUz5M4fidANbSb+g64ncF2p0xeR8zlhq2z
U7UFw34ruU5HV7hYylqXgdSZFmOe9VlKTNEB8RwrRX/e6oV/jpdwXjqWLnK6
ffy7TLBEaYgMM3dDfa+fUtf50xRwj7RG75z6mb7ltC56XNnVGPBj303x7G84
84SaKczTG9JTKQsWk2dM7k3zVPLWJBtMnNiwHHEP01216Ih9Z4JUWnjKzqfD
3+/p8uOV46uio1XFMywvFKESq2IK/BXfOS0Hw5ewLXoPXFKCFv7QGhMSgAI8
71Vaui4+LhjeJx6dMcvwLCw5a/Lo/3Dj+EFZ1NV3wxM01GWDrXVYhMPw96h4
sEvgvzHe6h5qBPjBEvU+lV3+R1NArjGDCuCHimbWoiMQuyXqLi1U4or+e3Bh
RQ9AnlMUSAP5T3kK3I+pAiwLT6drZTIg+XO8dRpTulVXF3ENJn0ovMySXHpv
n/tkjXCVE/oP+3Xhi3o9DsoGQp4asQ6EQGKy5GIm+J+JdbUD6AzodWJ1HI44
SvHMIyP8WF/0S/iJKxU6cgPrkv3fJXlx+uRAcMWaSRE2rPwwm0lh7uw3ST/y
wMfSxLe45hHkWMHS/q9ZB0wJsiERL1Sfj/j33e+nQanj8EJbDruhpSp1fEcE
HGNERCRc4KqVARX/9TQ1kbysipEbPIXm+e9hLRnbeDwg4hLJSZ+bQzPc1rXr
+qkK/h39Jw/ENFKdO/PaoarOo6p/7fxN0jBu4cl8eY8LfQ9nLn0itENbew30
OxGulScmy7AUqQEUiUxBE08OjUG+45B5TRU3fSPxgY/ggiiOGM5+whJwb8e7
6r7NHzFI3NPIsLKdWOe1vkgYXc6N9pZ16YFKbdF0vk2cqBi8P6KWrzSwNPYs
EJoghHgp1GbFXWF6Qvsbs+DTW9NjhWb9NGTh/2F4jNiZc9N5YvZ+7SiLbkzY
wDReIG9QQ3NSWemC5bHx1MiZ5L11Ad9OTky6VXCqzBvv0xfX520BYGppjo73
N0+dMMS4lYSChtJRXBBK0uBC1EIw5wP5TZ9CwMsX5Vp7pcIwjGTLCU2L4gGF
zHnZF5qFEQn4R06qCvDQl40XGO9In6WQZG94f7ZVK9wi4hNsLLXOVIfuIcsu
wdqVEvokLH2/yQ53r88USvOfwB2M12mgl4+5C2hLx+Ywq3BNcRxaWJMZhHPz
0RS4AYUd9xFzVUpPyoADINQrfh6EwgbzEEMESNlHsH+3Cay4r7N2Ut9uk5/S
+L7Jz18eX7ogSHjWUrG/XkYfjBPq9GVh+PwJYXqvKapDSGWdfgWMf30HE7Vl
7PUZkLF9bzyBqZQmHRXcmTZ6Yalyqg82T1UM9adp/TZdaeWqZpHfT8o++t2j
zfXmmwKQXmXtfyrfMkDI2LFdVakiyRDGDuB++SEDVo3Z1OO9QP/ppDbgQ3bo
xeVT7ZZ4xg7xp04Mup6xXgWtKlBftclsVFdphKWgi389vS0dWKAni/gXFCcT
rXCLFK87Qy0GkTMMweNj8/HFqNPoj7jMYrw6YORkRC/FvKogOxv79/HM9FxV
JPvkApbUU8BknkHPr5VUe40u3N8VgzyTIPk+5Gujz+og+Vah8W5C/rDx+gV/
0ZEiF2KFKCQARNx6h+iDaA3KeBNcQwjp5fmZSN72hEKiVG8xLimrLJMGrC5J
FpIePSn/NOmS8WFIL55jBN4hv/VsCGyG29rEuFxJhQaYJfUkat8zNzcxK/3A
SZHa4a1N/G+Ng0G0WL31jqxwLVS9xRkhpXehL35p1orRtEEJ8FYB18XwH49O
O/fYyI9KJdkQWJDodo7dfo3wd58vIXRlk2npvgFZAV3F1KJ9TYgyEzjahwkP
OPBPzy0O6wg+JKQPRxO+uB6CVWyVhFpRQlmAG1h4a1mt6ZXKRhkXU2ZT28AZ
cYcg1SboZv+QCuq5FI0u3bnffVdFRACOpoLMyLFSA4X4ieM0W/gIgi+xs+J4
600t8O0aCubFCaOzhWVdyNynUl1kdyMaUmqzrd6sLJsQ7QxzMjA8EM2548tw
sI0OS9ptBWyaL4qEdjnv6TJfOS3roWfdwO7BCB8Oi+W6liXKSiY714bFvflU
weYy5B4OBeCNpitCTy6tv7sTytkE36C1uO62BLySDwb7kVa1QVywI8+bQAyB
RDzZLtF7S2zdqol/+8VJurHQAmcCLJndYC6TKMKz6EwBpS719/17r7rLlu4P
8jYJe8l3TW8afx1nqxDr7KKPuPiQFuIb0pLIxmfC2Gm0CE6GbYbc8hp3EWmY
LmUkdYbkO44WHe+cX1UKI1JdC4/Rf2XQfMUDwbnvSjO5oxG7RreAn8gDuPEi
2cl7wLxALMzBXtTduGBoZycsdjo96RLyJGwh/ZYCRaHJoHC1WJMK2Lnl7uRd
v0p8CtSWydkdNjBNAOOeq0RyEkEFX4ltlyMMk+aLKcCvL0S8rexUZTUCmvbq
Ci+RYLJmL6pta+BxJeqC35fYnz2FWP3d03f7cP2wsAne95120ftsgnZ9nNyD
5qjqnFPogXuKL2YQ4zLXzHm2Au+YckH+0eLXKaZ8YBc06pKCIzlfWAcxOarT
1NvaTfC4Gvny9nBKp7ouzZioO1o0S7XmQKTVUXBt/5RK7pm1MMTC+/CfyxHP
mQ+3GqET/gzr5Ct4baQvuyZkDIQgtpaF8GcbLgI65clDuTwfrEi7W9QxjPOw
oZkJKMH9ynhuHRBTaInQbLAIoJVDgb6nEgkcFPEMiQdNr/Md31MzYTCskgq8
uZChGa8ZNSHUUMS+oJn6IugsGtiQu4KwlggYN8sv4m18VZFaNW7IUmhM/nir
58XTP/9Ng3U4U6GoGbm3FOJtdfjVsUfBTwjU/2lE7sFjqUjqZ/mQdl+XgkxI
DzqaxLXeKCKwOr6MIQLfmMGmIU1i5EGb4tFlArg4j7rY924dSb+s1G6e1LMt
rjdv2oSRv+fjwCfUg7fnNvyDh63mZGAHujLZX3RJrYW8osrV3Pt4c9meC01c
VA6Z/Ly5VQeasSU4rZRqCnIqaodE0UkbnNtM0CsAefHHWrbctIsHLauo8rwT
Aq9y4JtvocVyj/u7i5mk/4PNNfnLvUW1l8BhPNfaLjll/kJQs2DiKi/SFASi
YJq7f+1UqyWzQ375g4SqkUVvplhT0DrDqy6GpMCox+p25XLAKI9OZJV5yYJU
kOim41NfRYiWE53BRnL/g/RYYK1GR1z7iFfsHF20D0dcvuV/OjsGJgJiorka
H+QPVSX9fw5eU6XJFnr4ysgXYd5Zq4nEFVUO9amcYQjtUWa+WuHk8BbYMEWu
dgqJKMt826Z7X6GzYIkje1r5TFGm+iJtoFSvneSxwWYplqdquVldn0AnagJb
zCWdR/joSKL54B8uIe3Di8wH2gp0q+p+EdH0kiZkUwN9JiEry334nnVRIUPF
ltO3f7yLkmHuB7Ot5OqbyJ3UlXTwlq7XstWzTWjH0wM+Cy7vL7B6sYqN32e5
VUUIdefQ/IG7iHQ+f1iHn0RXscD1W4/eYHXWFHm2O28UDH33+Dj39zH7KMoE
amtNf5IzV/MTn7jiTT3dVDCeX8AgXpQjRF53DcmurcLYBRhi338P3pe4Ts8h
msr+FSK9EKc9jJNdK75J4o38Y9qUIvd5GT7cxsdpTlic0+u22mRioPULnCUP
f2RTuBTtF2xMRgwmePmgw1CyYfsoi31B+sWqFdg5OCIv9Q9/yhWagl+VGwam
gJpe+EtpehaEq0AzTNwBpFYuhBqsjYG6c+AlZB3SmAfSP9qZMfjQoDpEzt7h
+s8rYdzL/g4mRorNM+Dldcd2xbcJ5q4vZ1Lh2V8CKvJkOt1eCVgU/hfQXv9z
2eeGhZ/jVpXM82NQdYZ8i6GymKinQ/bfldEBw8FJCM+HTqxgiBZJW2R+J5us
xmao54P0pbQReBrVJIGBvFmjOMGEk2H5bgdIZQqNoRTYdrMrxKsxNXBGpgq9
4PE/LyMx4v/Cn7E/p5v/drkBdS9c2uTbaNdJDsstmUvtm75JmnJPEG7lsjAG
mSDSIQQif1v1gYfdeYq+r7dlQ8AxT6LlSSBTO6u6W8SHDHrNJ9g8/1dxWeD4
zvTf5xnla9DdVOSQXttzUZUscN6+N8EDF68b348ZRT4ZRTZdlxsDLPzJKEQq
AglMxvsNAtLVPzICYvGz20ZXBJugGFNlk+DzRk+wH0FzGZozSYybaCXW+kJM
VLvk8XzUJJCTj8P+qyZVRw59qqY+pxblkyCeAj+OAg4ICL0GkmhAOJssMZth
SWKh6pb8aaQDNUdhfFBnUqWYq4V8/auuj567bTZpraUN3iHbsg295ggCqzyQ
R/dOqodYxPW8xRpXZ+m9V7edODO11fpOm/OX2hhlVU6X3luQvb+QZObK3MHR
Y01xjZ1J2OGcJlhCNuMLa/7IQpJu5BlDDSxephECKvedAghM7Qqqg4iiuKU4
jS/gnvla4BJaRJGfDnaj88Q0TbQZDNONRJydQESa1KZxHjgFVroQ430OJf/x
AY4vMCyIyftNaQpVzhw6d1Ffu1LLzeCFXwlK1Gxsow2W5hbNysQYm0fa30Ri
B4cycw/ykYHKQCWk47vHwv4VEEHmyclx3+Db7amr/wz3CQRpI2vrMLEGb6E+
AcJQXKhJLfBL0Gtkans28yUFouOll87wOfzH19p/oxNZaCDSAkw7acFqLuIr
ycgafQqXWkkT2J9O0XGq/7Dh5RVRx2dVYxRfwrC+ipVDe2kv/Ls6DN5itjg8
LPAYSwAeP9ogot2RSkoUtg43QycbEhDxVOVkELyOg6sTT4u+5to1fPhkfY7T
1p37+6ModORZPzszYCmPUDqK77nsJXErueqeFJuOfqCeZC2G7DhD+HSXuqwH
hnVyFvEfiDPxns+Vo21mdDhrmGaMytlL+u/LpC7yDUuGe6F+wtKArmBXbE+9
6ck1VBTpEQ9Wm5GN72B2VTMz/nXL3+zA5jrHpvSQrtR1mEhUIl4QA1r5UXFS
kV8AQretMVO2M/8fbRZJAa51BgVqjGfbMH/HatM+bZTGMsrpZX1H1kRwxa1E
l4hxp/kIIPoI11VodjCAMB7BTkF0V9nT1b6WMec03m+bjl7pzrijxcKO6sH9
23ZGayp4BmnYlI3TJRJQUjlwU6fHV7Tj5NTPuBvzf7Bh/WZ1pVy2ZrUT2utc
MsfzoFwywlcKJ33Ty/dKyFxaUoxXpBwAeig2mONbTFT9DtipZJvaG891scTe
//AuT2o38ToXKMxqiYf9Setecym2hcdfQ3vbPbpAFSnOl+BMSRJYmK7ea6Wf
Z5OtTYQ1P4j35XwSyYE59v7gfJc3Tn1RVMJixOmsU5JjZUIDhTkjEv7smmJP
4qH93YZa1/N06o3UccplMdODu9Ww6slhJaHSBalb+kSnw9CQZSGlbDLwAnzQ
kcp3lMeT2DMk7/uNZtLdV3tCIWUhj9QPpxCPVIUNeoWOVx7SpSUQ6+kwOUMf
hxIkSsaRET5pDf0Tdp+gVH5qSChF4gpogBcx/p8EGGo120O+eDFS8pZolu6o
HDNRFIYSMf0NfWgOXyFJ+N8OKC8yLOxSXTb2BqcWoSGWvr4yMZYDtEekDHlO
i+UgygXNFROdIjK3RLru+zrYQEMdZz2BN8Wsdy8mJvtpEGxsaUp449wcGzXo
qa2zn1AIeBLw356JHwEwFUsoerZ704uvMaHaJpHsFKr5NYl9z3Xk4LD49/wd
LrlGPkluRIGSYkoymwOKN5ednUUnOkAs25qIioOz8r++mpj69tB+w66Kf2dQ
YtTmMbfqBve/FEEpVP+6TBQymrSpcNMzUDlKyF4FOMw7gnokSnOIoxszVrzM
DH2sqWGaz1lrvPV/Wf7bUgHYzduIbCNb31wn4GN00J3/jjvrNNgsx3CSMq3+
kwEpwQq4uYc74AtSZgpdeTX6+FGIBeIJle21dshNbFnRxbQykhJrEWXPiVDb
fpSTPcEQMFe9MTLFe3uI98AiiQrQO9gTui49hjxiJT0VJ9BKRASR3lQJPyPj
dYOYAIJCLxl9qVHa2j0yoTLrUXsPt32c8k0Ea4NoWgZbHuOtX6PMbe+3PjIN
+tHP1eWJgzdNbL+SHSqxmM5Nph6uOg+cYE7UevCCEbOCCIgOdcC/K+D73TEj
Mz3jZ/YIaGm+UpC79Ib7L6/w9hkg8bTFUvbjR5iq2q2YY5oPWnfZXOZc7GTn
3LUH8il2LTX9hwoOU6QyeEFioVFoeF0tdrBsz7m6H2QwIGtbDhuLdYWfxDrG
XyVhxOQ2IOO7eByCunjPSdykfqTG17ugCcPYEt3wsljjyfC+CEMbaUKTk/b/
pH+UFb9b3umCLh/lGHgRHjhREERC+Ho5RER3aieNjbBJ+Rl7egtWoQjxIcYU
FRxRpiZ6ug2dOMRjMA5uPG84y4MlnsbFEKlDw6H2ZXD7hF76NW10g/W5PjSZ
evzeSBHErbCtuRXbklC9nq4Q19tCZSgf7Vi9yg17fMShsRdeH4aSIPRaFUaJ
tc0tu/+20zBTkq843RA+F+BW8+HYJ2gvzXDSOd2TbRoSGu80dF5SCWcBYzwZ
EzanQVUZFsYAEDeNrbXvv1UlV16alaSvRpFhDJ6qMLLpdvJnxHiT9cwslKhh
zM13b7QrBmpzuMQiNB6yazBpr0BaEY+wnUww5lJw3UP9mxk0GOoCliR500dh
RE33BvOXyorNZA8LaZ22IRClsBajX+13E1VJSutjRYYotZIhj+PMUJ6VX7aK
IclGiuhDfjnZcpQTRWRgF+wsf3qj4aR4BTs9peZPqmI7oR0o+3sA4T96otLc
xZ8jU2UgLnAodTyDOJR+xD6Hd6073GtZYO3llonsGdz6iJ3AnJxuyS5lZahI
oz+uZ1ghbeN2/gMRItZcD9ums9agR7hwC4RbBepvzV8l6K1O55GVBoXJyV0k
1CBwdZJ2404QFU+4r/7Ogxp9yyaBLEi+bTO/dG1DPO4t2S1BESIPIkR3vfuH
UbPKFcftXKxEOZ8+9VNezFn5JCiCtrunibO4Z8DRUhTVesqDbkkUSDsPJ37P
7Z40ZxSpy3YxJ1ETQ83lfHjTFl9YO7HdFtsuTbkok6Drplm9fVBtyiW5CfH6
nsXMpQnkTEpSZ6YOdRrKku0wyJkmUoMohHxPNl1EXwJ208bycEnbLKnvT8EC
wIZpaH9UYCz8o5h1V5pRGYWgWjard1uKdfF4K6YepvwZiofFaENt7Cex87Wi
t6KGfKJv1EvsOR1jvWz+HTK9cYW7rZCx/8YbElwVUNMDEywojEnx8k1qXHxx
+XfosfvcWjrgjtWx5Ixoo+AvZNm/CXFLXZby7jPkvuBqz6Gpqj9sntK7SVnN
YVR5dscPVbSbe0J8N6d3Y/FFgsCcodByUQHiX86YUgfLkG9BS5Hj3ncUBjvE
xfyDUZus0pHhA4SXz8QbazWPCcKHoC9DXkRrF+iLDko4sLyU5gaM3pNfGtOs
teOTVrGnXtZmuJYHdjA1jKs+AF5OJQQTRwOEyhkYKeoQSamrUtqTFPw2CDik
QdAez31TM8YjBsPsI2u5qi1tOAM4fzye2PjGNq8fvnlG8lk/9iGknDjOWcHM
NxrR3XRiJOWmWFQPIXmiL6IdEy4ocM++s4M5lMncH6K8bbeL6d+J5DQY9VXl
We2MJiITTyxrkPowUqA4urLzVzVpfs/Qq/t24g94O8+R5LtYFEoX8tZ9TC3s
oDaFlQcSgYzOn5wpJ7GZH54yjw7BOXIVCUj8rG7/kE8VrfQwc1+3QiQwyStl
7GJ9K/EmXBzSoPT6kyINqB00sATR013ZbJm8l3tNiimxcMDDkVaLf0NxXhz8
u8f09sw2LTMHXHuY4ogr2N9BaxdRvyuuH9nwfPJM+cURFanq8Yz5kgpUgqZ4
We5RfGYfKSa2OcHOQPObrReJxaNAr00ylMY8dnXrVPP28c94h5sgpCnmmy3P
KcH6a1d/vwjc5wxVU7Ci42+0bGCOsa/UcTdeWR2TwRkDc9dDO0y/COOAktZq
hsLlU2L3/Mhp200gkDNSFgLcHflfo8kUQpCb0yQJLhIGfWqZv6zR7NEuk57m
bnw83PN77CQPso7Fk935ajxbO37JGiAsv3IFTEmSWDtwYtEBECuORwCKdFFr
FDWg4MgGdzsxSHXRD/E8LEU/XsbXEN7Jpotf857GfzwIF4pM4tqHzxpsiTrP
59/xJGjeQ/I1RGtsOYHwSAd90VTxAOSyUE4ziFlripmyG3CuqOWoldLdUWQG
JgaZS0PqT89evYYE78ciMiC9pYXXnX8zvP/s1NFuCV02bR/ql0Dfyk6BBN8p
UgY5b8kr8hHbGysRPKjdQUtSygMyWturdynfJw7ewoLgNbWBpR/IX3ss2AQ4
QS7Tg1q4bNlK8iqpg+g5ns5oYCiZnGT1ZCCRc3MJQ93MzRCe5CmNzD60FKmS
w5XAYP+yhzj8MyGjHZhLrUVnJdR7GYBpbFA4FlRHGl47PUb1HI8C0/qY/eZq
AJfQiPQSCMfcrKLSAjbtPIuGQwtXEuy4oh2zsxCYq8TDmAUbMuMqkpYm8KEZ
vWUzMO5wIlviy1wSXzQdKwcRm1fX06jEj6I5L8Vvkjrv/cB+Q34YognEHR2A
RPLCzHII9QUZWvoVvACBRN2+nESJBMyvBGj4DITZwUAtjKfrL9l6DiWdntMY
wcSKaahkFLRUpQIq0rhhlC2e5UDrR97Ox4Du0DLYPbPmRsitF6BeI4YKkWEw
F0vj/X+mSDZUqNvoCX1D3/QtNt5OWxI9M6WmfBVDbbHcXi+a9zEJkfhv3cLt
fcvCjjUnyHOhMja+E8IxLYA45AFLo771WLLxoTQdoSsk+idA+Ctq5FTXXzOX
piZmtYcdlOvndcEpScFNu+Fhcqgmn6gPlSwpjh67T08jF3v32Cs71ubP2GuS
zQDavPExeUu6M1Dz/fEKGgiszRq6+CCQJPLHAlq6L+Ib+9DYndwSPZ7BEGsR
/nYTBjk3jbwb7QqsXYpXTfAzhf86cEP7q/6tvh2AWHMNMX9N5nXJ62U2dxwb
hLvSXLXiZjEJAuZRKz15TPX+DdiXgHSPU+5gf0ZwTxi87+2JAaxCtCK/q8Iu
Q+PCb+pvu0Lmk8HgNLttwGQH27VMbOWqCX7OurbdSItacb99At0bCGkuowaD
m67lIZBzeKVtQUo/Z6YQwqUJNjvgSnMirlJvOLRc1wsgkuYTzV2857WUO7fL
GPcpuJA1Pzfu4mzKb7YT1j5Xoj62P4CC3L/ggmiYGB38fIObOGukvErGjwMX
xPT+SqTHYaQijx1H2dClXmKDipreu6sGahMzJoaHXHm3dYm0yvENYkDChH4e
ddkRSgGOoMv69XkJXDgsNXLrolik5WK/90oMF1nKa1eDI6KIIcYYoe/7IWu9
cjYFOoPWUuhXT9L6xR2tHd+tJ8kWLW3dEKZHgD3rVaTxmlQS1ecmPGe6KT08
sqzVH8TwN/WTfx3QSH1mZLK/rbAswXBzuFQQedEF8S9x7PdpXzfHEmpp1rqq
mZjlAKbHzAEdgLLoi72lz47LFDeqeHrK2bAihRb462sdvNH6h8cdHQvPFZyZ
yorO6kEXtXDzKYhYXnOB9lfiIbbguqJSvqdeuSG623IjBvHCqFg6+2+UrVDo
OxaB/8o00nVpvG3IMr4iYxdX/GkOhL1eemiL5sP3oDJSUTjS574J7VdD2xRW
TGQz4QfyVacW3c7hJQj+oK5M4zlk/Q7mg5PKJbNlNc9elweMcdOXh5RRq+E0
JzAYVDzb87J1wpsBaqOZPR/Knj9GAItJclDB3/vTeflVHtfKERTKO8l+cayD
moCLrsKVZmKks/sgtVbVCtXee3n3m8GSWDQ5EcYSg83S9uDJ4KrrBIfiqtvU
gp9A405y6geaUELhepwnOR/urp4k+BAxrHnlpr0/MPxxn9N5bryEoaV4vrie
d/8/Fu1fHv+arsZPlAf05IYYXxjv0lP9ZoSzZ3gXmV2ToMES1DjVnkqM3eJK
NmSHjjrzMV/BKGxQaQgLiqouwjZpAM2ZlEizmIpv88jGwu8xtRzNEwm3SR67
jpW2NxcHFbtv1aQ8FHFRZ3J+B7bvB1XyVkFuJ/9IPTje/5N4Wyx8FySgwahf
zOXbsd3e1WEOsIT8hIiGyoI3WK3xz4aep2IRIT8HvIxlBR1umKbZVfAcp10k
bHfWHZqkbnlKDkYrWcpG+t9pYidr+RrgiwrgpTJudwZu4e7zDet0Vp8qq+da
20/+NU1v9Ckx4HbqC0TpDuwEXtM0S601FSbzw0Sv5SnNZJZUUTvQ9rWf9A0d
jE7KCYoX9Cl/ETG0HHhirwtmthMW39vPg/QNwPBQ8OrjESVIpAnxRO/ucz/p
qVZX4Hzzz2f1+GI5hlk3Qu7/BhE6xnkMpX3yDDyuVXSLbbI1anWpzM+qoka0
1jIv8P/x6f8Qbh2NTcvytEuVlPdGuDgveGAWHYmFJ+H2by6s3BrKy8RH4/7I
VguW5uq3STZnsmKYUZW6OFbS5OMAJaQ6AVfPXjxiu0ziKyCn2njNqChU0BT7
u8zNIvBZMpP2eyeNu3Kwa8QlTUjL08mX0sn+xIQWQxLSWIYoUoDgbMxhitoo
IYXf0IbYURrqsMe6N9kIuzmcyA7HDHcxTv9DjC4OWBu9xFLJTNpKGwhbGjSS
dK5bgfIigTPn8sKzL9VZ95l8VEGs3R4EungidNGn7ewyxdTVXlplOAtq3/Mn
2X2TnMuWUFl62G0SXthHkk5r914gWVGo6CImv4cHi4Ny7qq1j5KEp3acDqeZ
21Dcu2hJStR4Xijt83x8LD/gFxePD7TKXvqdlS9x8OecyIfURqlT7vqa95q7
qbiL/bHMYXWJ68KLCy4wFFzzUm7kCdTOi9ibxZ3+nXQiysuIgbBMcRTVoH2h
gccTCjU5hyjH64uRq5Xe/4cSA1R0k3l7Fukza7pQwmosUGrM+dViLmIPxzmg
TR3LnnZYwdwLnal6oKJU7mcZSCH2Fz7NGZW0cUpP8EZtStmIwN85S1Jg6EIi
stGetJYiasJ/ugwdX0uGsmWwNqJyrD7VOq/pUs52eal5R6PwzlrKK9rheuG4
9p0r+X06r4KVhwe4ZLIR2sBMC9/FSse5t6ZVwzOcsAp89T4mRcRpQsDBJdjr
o2N0aEgrU6euAI8maejJsoGnT7nc9UbKEhP6AYTNwziPmVqXF61L+85ewLIh
5YwZTdFPJ/x2FnhXA3ZqrBpYppr6EMabrfbJtGYXfljw2Sse5Ra+K0uHxoTU
L8KUo2txPI8L27V7xegTnZ6JEszJCUVpJ70KtDsutv/35gJjzhEqQ3zhGNla
gOX+iiy2D1uEWnPOuaF6elrVM4oZulAT2m+BOUxW6zH1FrRZjKIpsPA22Q6m
N9PZaq5mRULtVQ2zcFuQGU7BpRACDBgz06EosIdoO0TMWmB8AYh7lB0L/MDw
c1zBHUmYcM28QxoU83Z4MxwmKGGp/abJMzB73XEC3iyW7/7b0EXQbI+FdqKu
5kOkvoadEOzZX0l8Dn5ouFqCmFTn84CYs7xVl7zY4m/k5wLCdUTrYVx6PY1M
f6i1hGN2KK6VhEWRZuB+pz10ijpSPFBvwg+0dqLcWnIfX96bjb5N27D1QfRg
+k4sMCERf9468eP0B2iMG09UgcNa8ERzg2Xky6IKpTteNAPC37y21CMw9Nd8
rJBwcBe7IiOBUY8YEqA1jEhnpFy+J+OoYBRF9rtIxnCXbIn/zsoYypU6w9ZS
yWrGMYqIBRCRNh7/lDAqV+1b2h0x6KZVxGoiDT/TExB1HWdzaeD0GRfkRu3M
jq2ipOUPecjfherazzQzCqeQHwZrlVxNqwcX0cmwHqL4G3KiD94Ss0tYCtPm
4BWUEH7sBLJSGQiaYd56mDQYkP6o/vBFNFtnRyUZCmLbxdX/JV6qAGmYmBh9
PcTt895YbdTrbvzmSKhUFSERLa5aL44rCDDA8v/+1894chsmUVlCRBEyNeGQ
4vfuZlDrMHzcsjgAiTEnvMSVuRCkfgLSKMh9VAZZK4wVcU1li9Shb0f+x39N
umFq6ZQnjiQxSPxrT2wjW2awRw0ACU6qIDkSFpmxfzm9FG9/Pg7hHYNixl+F
o7TREiuwFfB3Y5YHsZIC3lczBqTi0FCkl0RfANNS56fQ33K5rfoHMYkHzO6e
UlH1cKovOn6tE1e+9FKS77ZUQJ2m9O4yc2eLtSvQcnJx/gmtlQnrEhpgo/gd
mD6lRGHPRkMdNOLq1pflObBpCeV7fz/4jBDmo7/RMV1jl1vQ/uA/shbCNW6l
1HJW2FDYoZpglqrodsinYwKUM5/IkMr91S4KylCMN0Zs5BlmuDJ9QTrrMHUN
iRK2olyrM+Ycex0QWKqQudBA7146NIbXLpjqHoV+F8MKK3WeB8z4dQFV6PjB
ktKxOqgD97+F3Ky+QA2vWfbPc1+zzjIdsjtaM8DCCZNHwOa4Q083vdTZkVgO
flKnQO4YwEp+Us5vKkPuxRuf6s9yV+Znuu/qa8lZBKFANCc0/dtGWvadPi7/
U9beXI9OjAy8tfmykWNVfu1G7ZSkwBlqT/P6oP42tfmd8Nwlwz37LAlJeiV7
AstCLFHA3wHUhoOIXFF315SVZHRC3GzI0jQ+ReXtJ+51tsPNCDZzp0SztreU
E7+gjCd/WinzpWldxh6ZhD+4mVuAcBknUT9bILsaJsvrQmb/ImIohoszlIBG
6MyhW4N4mW3X2vwntcZwnDXiZJNHRn+tg3+kJeemnGmk5YzqQPGqFRdCvBkz
XAX00f/J5L80EE6dcJ6bXnzU6iQKYwEcMz/49DhHA6dzunCAZ2GElzsdwKne
7bjtGvnxhRTCYN2jOdy/0myyPq6QxziObwYLkir7LiCeeT1Lauc8ZPRd+acN
BTCKNhEY00aiXFxnB6Yai2wsohFmUySshWIQOhfuBnr5vzouD2c3XYEmBMM6
jmrFESTVYDFIXx15fkFh/xiH5LJLHBM/q6MRBTKHtmvzWO1tBoyhpck+a80S
EcZ9sRxlNWGk2sgVbaJMBVIxRkVre1d2uOkTH/8Lu2aqbqTglPOGuXjn25Qv
ovqvEH+0SA3j30fAirXEDHMc5pG4A0g0JART1pnooQ0x5i9VyIGR8IeyIoLm
jDNNaqz9Q1j/lvFjB7XvViyM/5VfXIYxZnRRT5aDqCL9GGILuCBvu5zfIir1
zcr4kBXod/AKdJoJ6iy4HEEvRgg39MlhSaTjPs5M3nxA56LpdYv3/ptbx+oX
YVgcAYOJmiU+mHJvuS4MxSXKhS1pWce6lAgklzsK1KzT0F3g/w7ION9YVSbJ
OHsU4hv57U5G4jjhE0up4EW8akO+LvAQCGAVjlXQ8VPuSIXKSr1gAo1NH9sG
PNwNc6SWWlrw6kgcYKWXf/Pb8xMsl9/P5NCYOcgWn64OVUxLVmS98W1pDPCG
SCY4Eu6FJKZcyfO8joe0+1iMdJIuywT8bE48ZHSmoN6bgjkXg3Zp2dseb6qN
1337L6cc6VGJqebvow7a68SqmnuVFgNZFNEuOtnC86JCB8FmHqIwdGuYVgZv
6jT04eX8o1Nj4U1iL6pzejGyRiKq41sZ3NQsH2qbJl4KQOPCLR3nGFRf6DrN
bf53rxSLOLK1FMuinIyM50XvSkkrG70k/raDm5ApvlN6tiOgEE84NWuF9Ji1
qAQHIK1/KhC9OAmg7k8zIDZCbq0kpznl8n8cwEB4yvedCNYE6uRjS+dWadPI
ZhvAFE77xCrjpyTwESXUNOYabQt7iapOHZ2dt2q8ssn6mYToX7G4Pc5ki5JP
+nh8QXy0F8f26tuodiVdOzUoX7dwtIZJlwiQkFfu1Ei7b+GwgGFgoC9/zF1H
r8F7q+knJasqJaD+j93Ag19EakpzvGUfn16nZVIFzBYQW+LP4xZbbvDOn8AO
IkhhIDwoGTIYXELOoAHRBVexV+h17Z+m+XAhCvMqWvRnSK/mB3IyjIpkRYeC
Aq0sfq041M06em8JPRsi/V29ZG8rtKQV1qoPf5o4NStDs9P89WHtpuqF5gx5
ld4hcvIwrDOHBNXaEwkNWltbmPMH1Vc3HNOdDHfi21RFr+ufDfAdISPVkAl1
eisBJ5TuJID/IoJAR3n+M3IzlJMGyv2iiGCASbu77B0Fjg5zAV91wWUHX1Fq
+agX+ZSYCIHoywTagtJLP84xlmU174f8bGOpfy9xAjNqJ2ANE+17f2SD6ZME
LnpJgmOt+LHluDZeAx4z0DoNJBo1CaCaA2dL2TbXpnquAViB0gvdDmJDUtHc
7vZ02682QXgiBnu5L+vZk1xIcPSUDdIXbJYheI7cms43WM3qKfvZHZ76AAij
8F89pqsx+qXkW1A08ZCM/fPAA02VMaBFJhLsJghJz2FOfM+HseES7Plx445h
ml5gqDo2VslPEAMqTCx6VrnoFU9AMoFaH1z8Vff1u0sao7wW4uecw8jd3qOl
sZOfjHOJaq6sqbdPdBikVnOxOPfCQOmrHY9ivSTvVbxShh53eqBPckzu32yj
sFeALqk0uCrC9l4rSC2kXjnPbW2eO+U+4G4yZaGht/ZOvpzy4XpqjWP0OVQD
9o35rpEmxltlDYZDWgx0SQptCrhSjyg3aIRlVfCQkwDxLOC5fPTcqhLy7h9P
QiPPJbbTNnM/OVF0fKdtshmQ/77b5BWMF3UDug0iYxTV6xWJTl1+OnzoakcV
v/DMKIW2oTJFQF747BgVsb7eg2tCcVrqTS002RuQZ36YeWoGo/Zn6fUvuBK1
JEA/Rq/gIKuGbeZfMCH8Jiobrr8dwPnDmqhHTA9bWvF00fY6pfadiHkShwdO
gNo6w+xisAoPPBi1kVWfX6ky26XiSqlFb550aoYd/wKFOHPN5kiQ36OakyN/
nbBO/RxNsueq2Br8V8XfvgWIcZ/7K8LxRhVE2PBrtp8NI8y6wpArk62pi1cY
TdVGqay5o0vYGYcGibz4GBNW6m3KkLCcCvzYKO9qzwHk6b4DNgxcTls2uqky
+ah/IPPisP+0DorfwkyHVIzF20gYhhnK74dWd5NkjWyNd3Vey3PNvfDNjmid
81FMVQZGN4tTxyGJBErmQyJp7viDSC3UqUK20Sa66G80B3UBne62Ej79Mgq7
+GjsPEJxiZogw+HoeMegXwGBDcG+uhqKL2qngvfuqHByDi5QKBR4PunPvDk3
FKWmDOY/1Dxt6T8PcnXdAqOFG2amL4jkPnj18JlFnySnEqLYWe0i8jjlM9b8
n6AYaFt5pvEW+97e6wu3Mf9Fn0hY8PXjKCNmYVAG+id5HlXYS6D4x/C7qoiO
9WdXyievD53iqkcIEZdl4JLs9bWtWv13Oe2xPBbFqDgW/hUb740bE2jXP8aT
5Aa6+IBw2wV6igBnikt6uVA6ffKlU4U9RMh29BfYqEStU72bAyikaKj09Ead
W+SRI7dNPEW8bDs+ZzL6hqs1gA3YLDSXzlTAP/52B2aZuUg7XDjWhM0OIYgM
q2TTykQOYo+4bLGT32T8W1WeVmgMMGQ5JA5f1j18pV24Wgz7jPnJJ7dAFtxH
MG6PlGUSCGmRS4Rz3MInIaRLOipKHw5m7uVEUDHp0l25vph83LqD9I62nasG
EGgHUqAhgrKIkWOOZKhfH4BzWgoov5o0rQGxM/TKX9g7LXAtNK4sT0/TXc0Q
VQXVeKZ7ezndZWOqOsMsqrazZl1eDKFCEpdC8PsSeNu9C6cN61ovzoxpC/SZ
ed4uw3zQpzRIW/Q5L9llfjdsCWX1959nq5K5fBEkXPEgTXBdyz2Ry+krnsgz
vg05d6UxTKLmEMWcgBZItX6MlVX4M8i1tA5U839Ptcq9ynBJNugwHPCMPTW+
dBpTPX8AspHxNqi6MM07HufQY73GI+BvDgoR8aMB8XfK5nGDOmKu17Qhhbsv
tfcmCxqymEUmP9hb77hBCJX1vnB2AD83ets8jcvPg5whX8ka/kdf20/yvArG
/BKuozywAHcdUivQKeDpJm8GHdhHci/cNH2hoebCnYLgPvCDB/Ns0r7G2baN
gFJJyqq080OH4tnFcDSZWy4AdNbBdozDIkNclflijI+cwzEcNU4IIyrExNPT
oj+fXECCAmU7E6GcwXUOX8YbSun6+zaMB3wTPgiOj0EKH82KzgPcr5t5tcpC
M5F0KVVy07CPtiN4x0gDs04h8ZdQywiv+y9vX2v46Xm4wup8EGnUVJTBM7bW
b4rVuFcMzgin5LFo/+Mr2hy7FKNQEobG2xDnjTfPRX/WGW1wp4CynOaFK81O
FmjJk3ABvjJFlIj/f9XNEe6mZtqqo1fC2WPQ2sX5ajJIxkd3Rq/DBpPYVp/s
hoIcCM4Kk3tenV3kYyY71PzdT5oGyf03yupUbUc9NsYqfHWL6KuzRnRlPEHb
3xe5rsYw9tk0VZkNOWBMN3P3ektE77hEf9Wivil596flLsX7PXhR5lWDDjj5
eYtFItzOxTlwx0DtM43X014Xpzf/yX+wydm6t3WeTcDEOrHqNUQFhKbR6xiC
++LGF0PlBaErvo8KUvRv/lgUp9y/uLbeNhgqtnFZQenRx2ACjkhlb0+vtmIo
ZkAc8pS+vX/A6n416SC45wAbW6TU4w49GF4rmlTkWsQd6ofnfNvpfMATgHA2
WR5riX1UFYsVJU+adQaE4cNMfiNUSjjTKA4LEQigR+6jFIJ9uE20BaKkEOYW
bNXYN1XIZiHb5nn23Qy0Ju2reOdMW+EXN0hvlsEnWva/ay5sAbN5VEpLuve+
xPpRzFNguo7B4yUWx3+navMB1NZKD8H65MqKJ8qJNJc9dL74lhm0g4h31/LB
3YmRekLldlqpH7MdhYJGPPbMbU57Q2WCDNhauJ7LN2C7RpqFieJqakfCF9Y8
gViRZpwhKgJMTPdNyoSfKea7tYQGZLJiZzFFchDprnKvm5lJ9qrNQXqVBoxp
8cl30MWSCgzFPyE90diIYwtIXuGUcS4fczGij7FzNLzWPsjShwWPyYH4Ksde
mkpT1PFU5CVEojIhSNLM1E7yysORNAOswIEOk2T3XbjZVGGV7+9sMwQDQwJ8
OYT/Jee/Db7T4Kx9BhH6w7ZI9xkegZwJwXWTowL26eoy9jJkmJSHNNMpWRK3
kTxA71R9RrZOe4L6UQc399dFlxo1+4GIAUBqoLoQ7/cpNop2RqhC4L/9nANb
Yk8JuHJAdGOD3tFIm8i7VH/J2qK88EbiaTyBZqvXDs7A6qGlOhCmkj+FYLZ8
MY9FI+phtg21lMWHCTqoqLEzPkz/L0bMZxBE+HRrs2Xu+NRay6hanauQRDi/
41rAS2ZoJaB53Zk/rCah8C8Ycymj7ZBd/f+7PcDLMIqvCcwd2AvjEJdNr4Qo
zTGANr16GGsm9spD8hVbJ2fJWFrGn7iBxyo3gvnT/Xl5HX6H+ajXXcHqUh1r
mkGrhgrDdavkD1J1xlIBpgHEcq/E/1akIBuArJCpr14BeA+WeaJxB/r2/E4i
vAqT7zQzq0DybZIBkOOveLM1+4Whnbf2Wxl67KBAjTpwaWT6wP/sM2lsj8U4
HHB25j0Ux9+A5GitwD98VA9a74clNEUrVueqDT/BoEzZAOiM76rNLqM8m+Ei
bsVHjMs6Vn57jlYAkc/QPtiM42c+MWvBCqGo+bMhLqh08YemBRfTD8zlFR82
+zj9dS6t+YnEoI7EnmaXHyZ8bBpq3Qk2tbzfRunZ93yHyBCkZ/sY6s+ZiujM
fEdBGMMMrdcauSlSksjlHbmdCNd+6v6QPARmyDMybJ4eifqMtth5iXN7JwIt
UIhatVD1z4VvakLx2juG1Qinli8nRUz87A4MaJXum8VlbKQ2VevjuEiM1w7o
AH2ds5oPJ4VFHyEvbPjdsOFal5iZh+oVR91G6z/9MKikdaB8RGinNIahxYk9
soeDKP5NuzNVnbZQ/d2hlnSaLrViRHX+nxRdcpH4Cih5wk5Aih/1oeQKQqg/
L/Ivq6/b1FpKFI96mliJYZAJtBvFD4wZzlXoDv9Y0yYtMtskIgkhmIffsMZp
5PmVaN5diR/itLvLtxQAK85tNNiFFclf2JZ511W1geHxsPkiQG3KKdZMIpvZ
wcpOtuUDidGJY7EOvjGiBkwruxthVvMLdBJf8KZ7g2em6ThJkyZjS7bNUfdQ
eg8xv+MZb6XHSU32iKpSqFvLIQfzLIUjNT++5YGakvpDfnjttrebTRQBj1Yq
bTkhaakr8sLsdR0hmAqIQrqj34rWkkeD2weO/kz6fhGNdNR99bbJNVKQ1QFQ
Jw4Yc7FknKWRXxTAJOWykizAUpzzH1gorPdyfjKy64m7ktVjgwJHqeMO8mrc
SUfWzWzsNTU2LPUs/YX07zXmLSsgcG/rpF/C4Bb+kAoi83DoL/Q0hlkLG41a
ftYa9bAWFVbaU9VBt6apefZ+2Dzc+9MqHBaZRx8DwpvySR6shrEGp1yVqR7M
FVoICVtpXSjLnq/uA56saCqSTbnIWbadGhIk0/u0ke0c9ZwSHKHIAGODm1Th
f9Osc6TE6XIB8kP0nTOWJCZZoQ8WXGpgoe5B950ondnzleOGjxSj+z6W05/L
RcjA//z1fkstuiJsKsFQyfc6FJDg7nR8p/HETSYrarAmbRW2LdTWPYAtpCNA
8KcxTTdu6KyH8KZtva66OdPqgE7pjr1Tbiy0InRXTPrUzJYACahlem58C0bR
TSNCsOjo1tlbTFLsXSpUHNSFQQBgfhKyAKqI0YjAIRhLxbltOzGY3Td0tU9O
JcoPuampUf6k3/DQvgeYuOJYwKWQR5XMKtklL2xIoTvcewexQp1UyIYHcUUZ
BzmawXkWaOyeogxWFQwM2FDajGnzWbqPPYwE/qT1s/6WDHXMBfUuifaifSwn
iTqj6qptRVN1aXDjaDk7VLeMYOQMO0RTL5EHbltmA25s0va6DxsFazt4FPyd
uMeLsuP6m+EfXc2NTKgxS+CRYlkWGFskFkz/pHMDDQinwhShDCye72d6eBpQ
PVNFuH9GyJEhKlqVRabUmc0sldEpLVtTMDgVf8ivpFZnhtuwKq3adCs/E+Zr
yuNh+2n6IZ6NCScb/jCuHbbercEe/35WAPhiF0v6w1zM/nBOVAjhUr3cPyoZ
3PUrTHTbgetZzoDX8kf6kbw5xJp7DUSfoW1OrfbPB6J9R6eqythBp7Dxi1SA
S1YkUI7WzB1WWaUZpQRDKc7L5phN0R89DpWlQ3A2NWYRnh2yXEQz1YsMxksU
S3LHQNeb+ctMXK4uKEpdC5smi14dDELh/ilyUhYJLjbDt3VUPmP9mmxfZvIL
MeKmJUc4xOy7Nzb0h/3yLyNOwTrClC8od5bPOqHcxTZsas+otKJ3h/fFY2s+
of7LFr7IV9JdiZZK68HuYhde5vuMKN7GKPamPhLM/bbLKKyccOMmRiekJ/N/
8JbxP45Z2KyTiXf5Z/b+/r1sjaqV06fbUtn/sxeSE6xjqIFQ0Z1wUXIHN36w
KlY/y8WResv5AyPCxSG6D5DoQy1emoX47yRGSTdTXz8zy5MeGBzEiJDH6LFw
ZATVmsLHKls5urZ2Am+MKG1JbMCez9sHYxppaHZy/EPDgIkD29ofkF6gzl3x
ZSgpxKpakPwe/MHa+oEE71IzFpyRrRHdh+wWnjXmrWTfNPI5YgxyyjWg8xEM
GrK9q7EkEK8CdFGzp1z6ZDJb2aqhJNdZhOOmDDTi4LVwCR+yU5rrZiR/qCTh
tF32H+gbjaDW51SX3iENMgfWAFM/JC1eAvD7QKZYka0hT0Gqf/uaqR3t8PCl
FtKxR7K4qjU6Cufgbwfm7cuVG/9okhKmJW6r8/piu8aUPXzwW4G5x+kF4JgD
ZSTNqWhOOoItmUgyLthBuTZUVYLAx9s+s282UohB9yzKy9wnnusXjSeUre/d
Oe7n3kZIk5ot6qCv50K2DU5nCZV0zLDTFVnBR91HbY+po9DZ82GUXya5YQzJ
RC/txOdY8uPGAwyh3OiQAKOAMkhsX7fRsKJn6j4fvC5DA6v88xESconjh397
oyfxo5CfETk7LU0NC5G9cILIZhSp86ftyYL5wklW0DgBxcbWZE/8ROjip4Il
djARqgVaxbhUWjd+0tnqTAlGGjsuQs7xVVeIugFxhGGoNC8xFpy4dH4rN0e6
7AKzL6sKqq+qjQTRLli+DW9iFvHG0CClXP+kk/eVHKhJC58KGr4nrSkZ1MsX
hy020oyQZ7PODMHlOcxa/UrD7tUXUzIIXGPjSax7b+WLEq27bqmFngxWfxHs
H+SUhq2sIoObp3eH5Ls6vPKc4Mt/4rqFw28kuLG/nswhOvTqELy6/420oslJ
pZGrZ/kQ/OuhysQgl0WTDuvcACcv5EnhhiJLZsUxsFddk6cTx5zgd/ZDiud7
NYgPGh15mFF0uFKrYUFohQ/kAbD916M2JWcoOL3OCCf8/odnM2eSWrlmt80J
U17T7tHCI/oo4u4CZz+Urej8W3KRUY937oaWh9un6oNnydDGAtCeexBOEyWW
j0aT8kQ0VUl1Av5g0nQelSLKm/gly32Z5/VKP4sKSjtS9PJjJ4vOGC3Cjsr3
+gqjWyBhmGQ3XGCKnvovNp8UJA5OeNy81jvPejtw4Zz9v3wwFAdFr5hymRSc
g4WGukW1m013fnmQxpEXxYiGNJq7Xj+3HbTnbmfOClV/PyEBYAnKWWBYpfHN
bYuA4BbcCSSAvRVdr+5kUnZV5P9NRMuvMQwdqcAasDOQVu9KyNMdt29cGRJ3
qDdMTLTrnJD6ondFzlrG4CigiZRHlTYYecNuRUwzzbM6bSGQ07xKOJTEyHhd
DKIposr8ldizkuDiLIbyxdedIuB2qAhgcegKu0DVfXFwY4HwjXrmh2yRn0SN
lQWMgTOEnIbleDd1CemCpHP0lSmtSUW2gpQ6dhdYFR81oKas4Fw0MheoINsK
k4IZYbDked//NfU3dqcsCwEyut9GkohQdq8sm2cr6/UCth59m/olN5Nb/nG4
7Nz82/SPGVaMfkhBo92Fc5ueGsCpQsk2EKjS7T6K57+VNjJLkeaECNo4x1vb
UOZ6gjkULJHVYUzPI5vF/6rgF7fDKBpN8xZ4prMOKofCox9qxT1x7e2KcFns
ZSq5nOQGJNugzZA6Gzu3Flyqi7NKJFVW3DcCEvKvfjr/+UfS1DDhzHpe+lC3
gwa1w/IYxnjAjAmUjW9zuyzgX1JGvFJWm/oiHMjfZHMy8dqlVT0V1m+X3sAS
130fso5FNxQEq9LOox+8/fjRnD62wzlRGoI3Th4j/aCUBtq55Yjh658iMdD8
wdkwhRWdyN/+Emk47pQgqRCuP91qNTl23mX3JH9OT8jphmi+S652SBghtN2t
CANIbZdVNZ3rseOGaa+dbsFO8qTxcTj+uxGWm6SC9F4PzOYRLa0WaD+qFwSD
7WI/AEt8qiXtqB/taNef64Ml2E4+q7hTbCJ31DG2AOWTtuFDgKrpSIm/WGZn
HxTpIPOlLgjYxlAr/tRNH3CnpYs2rt0puTaqBA0Va1cI8mB/il/Z1wXxd0IL
fccvyIee9LQC4j3rAooBtFwdMThPkam0TBrI10WAqB62YHD2T0Ly8G0hc1bZ
ytJVRb0Y7K/i8wjGMBSawQZtR6T4WfcBiEaguwPWQTE0FBYSMFN9sbDP47C9
wyYMrpsxk2f/bJ1rRTyiMmODK3O6yidenYz6ox1xK1jOsN7esJxJXF1NQBJk
nwi4x1hnSwrwsj9EKu7vwtMkV0yGmjlVQIxDZETba/3A1kTBe+rTo+TvCP9E
ah2t3dZ1XWr2JP9Y9LWyWsRfMymAbToLBhydmzr+/GLtCYS1Rmx/slBHTo/1
dm74O27Ic5tESOvJqKQIUXXOSaMsS4DIwjxfnwQ6IijCCzK7RtKeznlQNJjL
u5xUo8MznUMgbOQnx9xP6Mxwj6aLt0L18FwBN0n+4lQoaHBeYpl5GzxeZH4v
GXwRDCPCop9A3Hjw69qoULr5n58jR408wOmi1HYG4SEy7Sp8OR44YtCr3nsN
kOGC9bnKAW1OvHfusSZS2D7lXEYQ4qtOPC+Elmn/M43LFgsjQJbkUogmVsmh
MvxHuz52eSFSgyn3pvyBei9ra7m/Y79hTa8CWMKWbZjuWFcQh0aavu3NWp+M
TQIpNJbsJP7/NTPtXuu/tGPvrS/lCFsAe+eO+0s0R41oa2YGQRq1Ta1CcRBS
p0YLcUxAv96snVYo4lQrA8M1zNldIeShGKbYP7qSl2cOt2pVFQcwvigFrdFC
YEC83UtPVvHMa4KG747Q8iCY9aEFBUisWmy/vlzNzC47GPWcpdAO0Zlh3Pbv
QM92H1uok1BjAUooKW6JRTCxj4eBvJheER4qDPWMIGJ34vS1MXjtPgyuarI0
NNHgYR/SCWwmJS2V7XTwI4hnvGU2+mgnWxGzqoPO1csQo32w5MdpwvhqRbtI
cxNk8m9+8UrOK7MlJtz+o+4OVgT0wG6c8sBU5nYNQeHo02jr+l2XB22v9ZxS
P/Ft1k93BsmKhB0nSt9vGELMEhGcvaZ4RoIhHWMNxHKvGteC+WABPqC+gCyw
5aPE4o5h6Yy4tW4L3fMVSm7JnH9X4+ybSVUFf6cBsvE6pZDPsGHXe3Qq18QX
gIO7UjS+trXA4hp2+Mgq9Cl6jR+YdiW1G+phj/1v3Up8qdROTu/TpG8aVUnv
tE32IpNI1/ZGVJfpSXOE3ZlArlCn8ILnZz2eEtzqaxDo4KjOzADHGXX9kQko
/Vm2X2YA2YySAtnAqha4nUfAZsnyWsNzSsVSicS1Jy86uHQ9Xvz0sbuCIu3u
nC7QDs6ID3VZX+lmulV6TPEPKmlJWC6MYhbrju7qzVo0j1y1GxnKfOSAeXhJ
xWS9JUtNXjcAbaFEsmX78wrL7bxPC2T9LaJ83EYM8INxJISG7TRZGUo5uHsH
3/69TKVC8XXY5LYc5ongrGpnnLr9ij9cLbhz9BsMKxQv1oZ+Siww16A8Fwm0
dGokH3nYUhWztg42EpHQrkBXXrcgQPg7XPKKUB0ovd0uD+0ESudkIaV2s15e
2+GjQGGU++rsQ+f0CnupSOA5TiFz9lgeVhjAHROxTM6R74/Q6T/lQS0fMgHj
IGMses2mIIdZqHa8nCiUM0ptflokl3vgwnZ8P5+Zetu5lmnvzIOMGd2lWblT
7TEUDRUDy4SFQNtliJSfv1ayEr2WATZHQRKWgUSuWHjS4+MAxkdSSo57VJTU
L1Jqej2mKsN2Tv4sJS4AfA2jJOREstuAED5m8o456HXOqeaHPZy7Bb+FY6CP
170VU2gN0K9HsHwaJDQfxMNh/j+2P1DooXVeX6feX53Y1ErdWSIgccdTZ2Yy
G9DBT8Pq71qtKnbSdLem596Lq0V7nr7tDU6uu5FSC+QBBHmI2PCMpLNqxiUz
dgHUI32gw35wuuClO0sApRf38zKgni58e/HGc804/bIPuXBINcyV6DwpvVOu
2XaE8E9yEGAwUdsZxmJpPwz29eW6yc/KywX2aCtY+V55/z1aT/ZM58fCtsdD
ArvEzOJOMwi6Jg67hO0AaIGlTYQEH2opDDRWyDkIP/sxzUdMeLDWqolUorNR
xUrTTCZSYEgNeEXcBqFpwZeTqmA/bLdWc5TTwJjEjbdgPk4jmKpzAkpzdxHc
MRDbdeHtkHB3of8IfdylPPIkehmR9gyUS0qT/PVH4tn9F3QR24rVV3gW21B+
PK2/zTGhx/B0Ij8T/3UM6aGmbrvpi3X1kTYsx8+FKhz2sX9PgF0//MG8Lb5W
N7LNaosgTI13GmaUusukWZa6ibmKtGAQ1iJ6RH56LjDzO1AfrNKmWUZ8JxHr
Ujs1AUvd9d8DT7Q0UFTGtc7zKDxh/5lYUDPBGiK+MzF/FDlJPTEtZo4zA3X7
so1/XNev8gnjrMkz5LzYw4pIZOgarJAqf4Vd5NVf63XyRVyFbLhFSXNcDCpT
5AkKyHlgolusbzsqvY/QkSeUZY0XSsFYtO6JBFGpwvJuvSmznfa7tqObwVFd
x//6iWjmlHD2L14aWxaWp6Gzz63zwuObgXzoZKVrgjCZFs10+BvqLpR/5rcY
suUSqvmIfCXRLBKdvnqvrIHIyPwIl7N3D1YH3Wmdo84jqTXvUosrUqSD5A0k
49Ccy8E3fk6nFLQEmFvGqSxqd9djXki2s3UIYb9HzUMYruN2RFhlD2/wSmAE
SRmKHhQCEPZWKDgzB/jttV98zFLR2wYw8MiGqKCnGgIMRux1FL54KwsHlOwn
pggwSmbXCFEn1pedzq/atmBGPaE0woefoKcdjQ83hMBgvoTEuC+GBfC/PjXW
6yeVJ+/KZcYyQSqfkDogVl1hYFzjD8dK8bP8km0l1BZmfe7uOHh4Cj7LLkJd
GH2LBwZQFrkkpx6x70Vof5cA20Bqct3m02rUYIEM6RddJEiutBFSMysGewSa
vE2itq0M1pxrB5BPAcvtMwMCk57eHp3nx5ub19TMpkKSfSAQHYL1cycgKKU3
wABDInPeNFedOdcaK9ve4eeW6cqbk1B0BLj5UZyJq6qgX/6HLt30Ze6X13fp
zOgs5uifWcQY/hpNABsclTuA2dULXTTSuBulxQbinly8mdH4JnW2YTR3yJDa
jDBsvaAIQDSlElTBR9OoRUqGbfKyTpxusF+PIGmYl+1Y1sQeAD5hdjwKSnQ6
SSy7SZneLWVJZR/4fFuI3XvzI2fZXuwG0MsVQDH4SOA14u91Htd/Xj1ZyNOC
lu2f8x5HfPwBAMsVBsbHJlshudgkpbamWvF4koeZtQXsI+uOQiHJ+hd5MMOa
ZuOIvvCcbtGENz1osGDU7kgVzGroId/Bf9jeJY1xv/ATVLUTwvgp52VDLcx9
d9r6eAwHqTphgCfrHdtHC9Y2QoqJ3RMBiGtpu+2Gx/8E6azaEWrVBnKnMQJV
igH9bzoTmxDD3XK0m3OC+RI/6xnfcHA/KwRs7KjTdbEnJuwEZRYzczmGEip1
HaevjFNSLCUzho5IzFraeevtrBXMWRfUeXN1D5WkI/zngkvFysEZuewmdFUr
+DXwYg6ojgXWm0hvcgWXPuXutCL2qrhYS73cbfkFYWLrWmqj/XckP2ItEM59
qlZvp53fLffsAQLQ3tEml4sLfyZ/JVogtmlrConLgFi4VuG/VsP9F4B3qyer
j5MVOzcZPGmhmRdJKtJDLOMWGBfUSlkEB/ndVNjI/1YvCm0Gda8VlJvopbZH
+f+2ZlihbHTrHcVeemsl445HUYbFlVrxaoB8arKiCiHzs+TdVSRgKTIZ6LWV
UXH3+0eDpnkF2iT7JP/U/1HcMD0RqenJI8A2So51uHB1jgMFCtPomaMHqyzu
dqUBp5kxXVcqgLiqOc6YbjG49dYM5CL159WZ5+goLLZCSi5iufjdDSsYioMH
5o58li2QYA6D6lIzYH/mosfKzu3xQnMyDet9qB4PhASssFuNeB3CwNUJhYWX
1AgbjHq2OgDPy38gAKRvyVoaiEpJaZ1dDje0yDO+shXW8W0yz7qzAlGyZw2o
NfblrThsDedRZ3e+t6waQ6lfyF4QhZP69lEmm3wipgMVXCXe1BMBBvsPTB6e
5wMs6OQT/ccfAs90twCeBjaPbrOWZIQXUbUY1ER+nm1oQILJeW9n3AX7qt3X
nmmeqG1F5DVHC12ElJVGHMAjDnI69RkE0akYTDx+iqEnQgXMxqB+mBla3FIB
xhxsC1ZISbFYkeQtgF+SIaKTcRL1qP3tSOfo6CRUzXspkWTHFBsdRikCY8+f
z7eQZkLLbS6PA+EMHwNmBPS7MKpy6j02THM/AIoEHc4ZfEHqacr1VzdpCdT5
W4zcMy4fxUm2aZ92fcDAGIEcYj6RTSwmvJNYl0i7JJa0/s8SYh3VWO7QIJDk
Kioaf4WHo3U68ka2kNPO2LjBQwFJh7On9SbiPdi+oE0f2GHt9sruvs4vN4ri
mXhwITxXF3XixGJ4QGP3TqOCxb1dbsbAKmviYiZnU02Zc8Q+8aCxte6Fs8Nj
x3JqrUbi5Cf3rpVyj+rwFYwGnahkPOwwc7AG1149KInMrvHiNCh07j2yQSyh
XZ8JZ8Z8K1na9FRMokzVPaGZ1mwp4n54hB1asLmffYIKaBDq2CW64T0DLQ+R
q0WDYZom2o8LeWSp6cPLhiBYMilwBFBV7J6Glkb8YxRYXA8hkreaVeErcX/V
/1NB9porwQLFCvOLulWR1PmNRTfFvSxR6yFaqWRR+cxqkFUts61QGA6E9gVE
0qd4A7bz63CNghQzPgSPO6aoIuz7KQMt9MPgRZtRZ++qZ6QGV/fcKzmmb3ZA
iLo3qSd62VfKbVGNMzLHus3KDVM3ceu0s9ah0b8mHHRElS5UhT3/m35GyzU3
4VdkMcy/D20e0mQ1ZABJ7jTjeoBQt4xTzoVJaqqC3pD38m4SQ8zRGNPIu5v/
Yhe4NxPLgfMU8l/W4y5FmtUY4dU4x6cEQRcrHRCNfA82pIK5pzwCmJtltKcm
pM2Y1ox4Gbo58IFI3MMlvEQFZ7/7xxGml9g+i5YWOPIDRizo0hahNon+6pr7
dFBk3Py2P4s2GdGFK8kpMVCYBwuDJRB2M1ROrB6S3sgG5kdjmtsiGz4ywaWT
QrH62HiT3qa2+2URwDI1DjPlM+avpkkwp0scs3C287X2lww8h0skyuWDSxNG
H4BJwRaOxcOOjpNgdMGnOHK3o59IP9fTjPfFUoW9Cu+8Y/UZ+Go28qwtrDL6
sU6poi9BVGx9pYdnitTrlAegRGSHoUSL6OSz3EoAKspHUED1aWpkuR8s1IeZ
aMHcX+nRrALz2YsMwmUQKg9Gjak1gxFGHCSm/Il75vKHT9anFaQP23NzHet8
dvB1qBbRYWCcfEUplvJDK9iy63g3WJJLm4UQ9Scz22FUm48Ogz7DAcnYQwR9
rToPIeW2GcywSFhevXJLwOpsZ5Pi9JiS/RJ0yRDRo5EIPYv403iyLRhkzZhm
bVSHVIJFxE8oKAKnsl6CNehNiO2IgQtjSN4ZtwG4ATkq3n963eY+W9zSsLER
xaIAYFWs6kuunLJywkDuXuJNYZRhUE6r+Vxt14AXFyrpQn3l64gLgtxnfD7s
QpjSV7mehgpJy8vw8CTOQG8mp4JQOs4mp3WaVwqDFwUQc9HTAb+o+CkQINB3
n7IOiuZ8R43aSXfCpk+nWAwibn65pnrEKXqmMDqy9my7nCIkCenOfWhDfFYT
5/5Jronf064xn3EGDviHWXOuCB8uNH4iSyitBqJbvyiQYuvb5eujFfwxArYn
LO7uL9r1AWrAibDE9Fctdusp922LJPt/fMPviiirDvyPvsI5wLo0qUJgiyF+
SUKfnRpTd3yCyAxe3bnQnpB6iX26XVpwtsRApgrIneSzm7yD3CKy08SQFu4k
wU2O3TPnEfsKJu2TZhV9yoQYENDbszL4jf+XH2iQsxrfdwM+QADtmJOqydBG
N1Hq7gYg0VP884P+Gznkd1EjrzC+UVNTr28/ezZRd5o6BrDH5jxQ1EA+YhVC
JS7fzk4TOnD7AYKzwyh3cKsS3wcSEmj8JhFMsraKOnD25TBvzvl/sKJqz9No
OLq9B26+wDBAi8GOpOqFn+V4pS5theF5XNoGqXDTe1Bvy/uzDWsfH580lwcU
MyCd18pSSfRrmWEJiU4+PcLKjmYne+c0PnfSZMBIeAh5crOdtnClF+L2B2vC
zbmZjr4DJ3lnLvArzOn6Pc+m4Y39adsgNj4p9DlDbiFkx74BQI4ava9N1qzg
v8NrOLgC0SYPl57bWRs8OUQtbEqba/wqG+qONxL7N1ge8P9Bm6EAGCXD8Cte
8qurpV6vyxuPiGw3Vd1x66hgtorIxenLuC3ekSWr7NBkcFI2mVJRyD5/jnMx
oZNrK+iBrrj4nRb17BFQKgdtmzRVrmf4J50/XYK6XFMky19uupLxirXfYsyS
vzq412k38MQuJpLPMIxCW/NIQ/FtBLz83g6c/GzLZJwjPVTdQTC9+zv+FeYM
s1q//KF32JvimVzOfFEi88KTbJuM8+319uOORsI+1MPU1uUG5C/amm3P1uKo
mq6RyKHNcMj5WW67cGAmhr117skfsh91jM8DHIhi0WVACUXKT0ZKwptx5sJO
djMzbFbwZbN95O79sDQtgPdQkhtTXKGazqc+ftQLU0xJ1yYkbjJksUlmQqj5
sv5gli33t+s99kKDdWnhhGr7ZtUaNNkt6kMPp19UPh4JiTMXMkCZUbn7LcXA
QD4/JH+uu/XhM5r0J5nlsm7uIfGbR24stYKqq/n0AJ5Qw//Qe4m7dOYARefQ
uK813SJOWS5x+9PDJSi/EQzO7YcS7EOvGTff8hK8QFGY3Olka8VG7ajdPqUE
1LlvOlf/tmflOyEV6QIhORohz+eXjzDdUCFapWPPnH5WHw8APC8A1ZaP6yp4
d1P8CF7TB7fnVf/6TDuF1PxNMhVcogZ2bBL0xouNFT6MvpGUmby1lLkmKquU
CHBggDsgy/7iv/LgZqMbzlPWkcWyMrXjuYGunAnsFo+BruRg3Noqt+sZtUzc
blSSaLTWQOs1YdQiJWIZ1Hi8wgfOruNCP7m8uFjBxhl1zn0BdM/kJ6H9nSHs
symH6Wr4PtHiw04JcMlGM/q4XoJJnbJlhnf2vy2x5bynvFzhyHefcKVhAkj5
hG/E6P+hNUABUt/ZXnP7KG2eXyYDBfLBWSNZgrgdasIA5JcT9P7gTtWl37Md
Bosl3G9mWKcqEHxfO4o3ubdI57OpHOYwSguUU57GXy2HLjn3nD/63ycig8dv
IdcqBNvCxpnQACzVMgQtdDCrwH6ciHcRa14VPY/x/hZ+wJ7cvpcV8YJd3zLl
vFBAlqStKs4stfKKSYz0gunusVsnei+qlxYRhSejdKWDrkd2cRtvnb+j3b8P
sj+VFwdT0/PJMdXMSLQCiuMulaVRHmAInpLL/W01J2M5l4rGo3ZVc+ziKRwt
8H8pBMGvMdZWECoTHyQGifGdCmJrUnTFyD/HdE7a9Eht8efrw7JcEod42wuM
gPquHc8kn8TQGXBzzFOnRHKkNXKO3L1tumivW/NC7UN7rHAfAzu4CrjjfbPK
KF9tVeaRj8BTV4DO3Jxb30T+qLszp1CZ2VXJt403zMaypIWVIRhpTD47JKf/
5HeUZ4aUl1EYl4EIFAgXLAJ0tOPfIJF+2sDcoUy7s8AEp9cXBgjZhIMdPBsB
FYj00TnGNgicP90QS9bqCqDdZIeHWzm913RmKDVzUnidQGbGrXzBO3EJX9KY
dSgUmR191B6/FWhN0dIXPS2nAGxlO7lEOrYEvjfKpJiNhmhHQFpXKRECTGh+
gGASjC2lfdHCczKvJoTI/CPo02GZq83NIy7+rsSeyStxe1phTNb8gpCA/A0G
zjncFWLqalOEV3UQk2SJ7oNMoPTFiavM/0RQmIpgvpaxljJifB7ZUnK7q3Vx
VF5fr3VlPEoXxlddCvRyfC56OFSLOhPkyAPz98821cr6JW6lHmqz+eE7bFak
7hqfgWAaYO43kvCfU9z8ZNdqxDt1Fot0msEgVM71OR9XyXusWlOjvzJGKjKw
IgFvXI+F0fpzr9DRUsp7mUGm9W5Wt0gCwUEFex7WRlkvHJqzp9bMAATEA3+D
J6ThiU90h8YkLCDZwC/mCL1jOrWyBoQt4ZJD5oW9QWiMCd8TFFCVDb0F8ksP
gnaXwJg+0MC0uwHo/TPqYyklUAPTaa+cykPBTUfX29LPtI9NvXWRiWI/Ffwb
SBmOW6zV7Rl5DIWtoqJBFLA6IPMksFhJe0sROS1+KMJBVFprXT+1hcxO2HJU
4fRk7PCiwFsl78WQ08TQytqTFt9ieVGezX53dxwOzQx3lLLktPp0CipuJZ/Q
LpZ7ZU1HBaq9dgZJoxGEKIZc2Kw4k2ozP8gk+54A66ubMYvS3Nx1upDEm7fe
Nmc8Pzx3+F1zKEbmOskTh9ZgxlBDHpUJX/YKKi6NwPnfeyxtQm1Le7gX2D57
WyuhjYaoT/cY7m/Q8jTUm9MA9dNYWZSjD3dyFIeukNvizketANVgOXhs/crz
mrdrkdqq25hRtcjAgufPcWWRj9pk/OhgP7Nd/x7C/q1HlGikUtGP87Yfra6k
wZafucTd6ShvAc5heIazIioF00ARIoL/ZaPl6SsrSYWpW3lSQxGwmMSJvAhD
K1WD/tg+rcZg6NrG63LAHHOFErxUfPISigP21f0He6vO9mJHfAyK7ug+agvz
UDUErNySrShVq0KUJoZdIull/TxqRSkfYCPQEiGohaZobkkgElfzv0+vte6P
Cj3jq+7ZNxyA6oKoIXh+3fTFGs+oQIsxtpReAawMKQTzhjtVZzpKhbmEmbdZ
TEhkpXZDWLOQ4VV/YIV+B5UukLXeARa8gFWlbRqQlTQ8F65mKMLfE1guQELu
ygZczvmvR84o+kpwndfIY33Ms5lUFT5JMVUg9NreAv1IoPweAcsN288ERd2G
LQ5RU9b5sUIQcDlY+TuKRF6HVLHWDjdwEacCe6g4hlY2pcjHfU3LuCMd0tVv
DIg0o1GnJ+gupO6LFNabi51MbQxIZ7Ve8nocx6MfgaPmCFSWtSG+o+J06Q8O
SCrSth323VJ34BlEGNLMnbvGrjAKO7LYqfsJPOCWlmuNzExBrJ8NAxasXCKy
wjcC5Q1Cyyix2R8gizcgxiiu2l2SjHPcubLjRVG9AawbUkGwyPSIdHbrURN0
zrYYPRqahdTvc/fIYcd1lc8q70tyRugLkDsoAVP2bSEwIGPb+mvPwsmj3RRF
oEV8JAHR6AOjy2bDVKLo1KpbCNkPk/jEz3KuhgXm+257BgFdXLf3JmOst1yQ
UQBR85hiKNf9Xu6BUuayuPqHhATl1XjTnNgIibxymUiMWXzuHwyStdT9O7pI
GN8LQ+N2vNWsaBvFhr8+o7w82Txnf7wRlPl67FlkZnzH6SpFt+XLz9MVOXUg
4LssKX9oTU+Nl2vh4k/Ymz8kNN2KzGXvPCGdn3Y2kYsH/bIQjkVOsgUuHtdi
3A+05BEMz2yBo9cLI7wPmL7cx1+tpwc45tptj9m2QbUveDnjhmMAk1jvMRkp
AapXEXwxTt1aq52IWa1rc5twSnaGrCdwox/LjWVJz/+podJvJv3OVTkbIdqH
nes0Ilt9DGtvs6RgqdRhS2GzThbuwwMaDp6R2Je4TVXpRgkv/KhVxJprgR5P
aMGZtXiwRdDLbAEjrFur3+D34ubuLZaNvwhWu889s0NuhxGxB3jCB4T8EWfj
Q6QwRSbIgSFP7p4x/oROFGTZqtPekl/RcDBaDl3Lz50hIGBlcx2Lk0lGWt9z
q03WslYt2IEQuBItRGYJgChWKS89so8O6Jx6i+egMuCqw05CKp84kfLsB52o
aZn55qvvRdP7QKc2MhysvlZvRF0g2+s0rP0U/tXp/FgTkrVsxZhqJCelVdtO
6YKovCPyFfm7oMvT1qe94MgPBscvnRHno0cUv+gqxvWZZgPNl19WToL45WJi
sqSQPDfGMK6wacoPtM5edzs/uagRi3oQHzG3ieN4kPyWy53pjbyDdh9L6mhw
ajJqMjct7OvbuzzlZuSAM9NMaplm9JPPQmRg5h4KYhyEsK4P04LR0vNJvPXb
j0hJjYPmViaZex6RhGbja7SwK/cJ9BSkyA/eDj75rYKs4qAB7OXgzLxyJLI+
kdr7fzVGUOPLnFESetGXSuaIqQhYB3v4WSw7+NeIrOgQf/cpamuqU0Hx4ASm
OCuOJA+4mv2Kmfdl/kf+0F5vfvnsbt9AQ9Pa3EtOtZC8jqFt58OZHqfpTeeZ
qMexgEMMU3FxoFz8HXLbNIonwCce4+IyqxHYE+hyH6I6QwJ78Wyo7G7wd5G4
OCwttVYc8R5q743YKqz46+O/+nQjbj8bVLqCCKQpLMzSDEHtK22h5ZpF1dxV
r+5cb5HVWOqatVzhmNNX/+d2vVupQ/uE2wzshQeqTkhEIAkFYAdZnWCqaO62
MSuNT4mjyvQT8ALQ8xDaj42aex26k6HxvhfAEpS6+ONBLfePlXEECN8SMwEu
LgKNYDA4wII3iDHw1gAQWuor0+TOSphTcYRpiAOih1bOULOAdhM7f2khURzU
Ozaxe1sVHi87cm3lymJZ88IYW8vzPXcOMexpjw3XpSWmIBbbxpf1A3NpWLiR
jOD8ndsLSIScazr9oQScZlz4rYxlBHHw42NqasDKyb4AJ4I7BTVxKVxSkUW3
tfu7EWZudd2ckjKblANkth4JRjbBCDto2Ef9zJvWuDFQ97/sqyNKayldOka0
fsc9dJqTnZ4SOzC8TiNU/hR2laJ+VIHFLIj0HY6+3h6fmmJI/oy1/LFQmfUo
fsegdGk1mnPeUJ/CGfowGqqOnUaTVycCM+G1GEBRMe6o9swz3Hbx4co8umnb
3O63modlpJHS01IODNNt6ZBQzMDhqVk5gp1LFB5z1fVXEyBzMKZ6RMNwKfFN
PtqWrcSy8O13v4kQAFgfqNiMet4yjKDzF6dZRhgVmIbGMIn+YsvlotI+TFYZ
m25GnCv67xYE5kK84GfDieKilh489OMDRPi+4L4Dygd6WJMYn0z1znmSFO+k
xudylJ/1TQriI4+uDp58iJHGMigDRZBSFnpdxQOKPG3XSCFzasI0irMpHAwl
3KxUiSqvu5bFQ0vp0O+Boam6SJxOr/sIxHp49fmdgDTY86Jj1KSZlPXELwk8
2NtiMYo1b2A7Y/9vikHSw2MXmER76T3Oq3EyRtjN7sKz4sqT2q4w1l8cAmuY
o0R6ZDZvqaOwTxOV6itVo8a5jM8lI89wMGigeHCy7Qqc/tbgFc7MCvnDE9Mg
dl3K73Ztc3N3+Ani7LEteVD9/XHDq4zsB0g68OMRdchuh2efiBl563agl4RC
9DGBxEIm78fDZ+/0cG9K+l7EyzgSgpK+Yf5uSPpEffsL2XGrwG3bDea3YYLN
fVz8w5nzrv98Rc4OfnbZjTvd5qsNdemq4+KjvQjohEmn3mEk+VMw0mmhMPhg
9MnTfrvzZrL0Thyb7vSyw3ygHmz9eEtrS/GD5jB72rdBtI6+STllR+c7k1aU
35gNdzTrdqM5FvV2wa9ZfsfhkEXNNNbA/0RsgL/IhZ9PJmvunCIe1meBSk/6
uYlfFCxakSmw6vP/aFpbunJeEuIdEWPX/SiZQdh3fLtMFAkdNwV5wE382Dm1
mzUrJH8OljHVvlvVeevDJQkmSkwnukSOVzN+tc2kJOz1aVM9kk9d+hkRPS8C
frKLRVnn+i723hGv3+q9EvfdW93QO4agB5lO3vTbTbnapWDLNKjmItXx3nRk
+cWrRrbSnuwlKLzuPISkWmV4lVnbJTX7PQVW7eGKSGGi2E87HZUmm/lso9ju
shEAWc3mDkchm4pvRF2M4nQ0G6xtWMajpOlsM5bmIGBqYwo+NkNodKj7VHOF
ueMOowPo32djpRUzJq5X4lRSVt2kwaXd8+AvpCZUtQ+6IbW0qSUZxV/brCyU
io4LXA44qxFH3qxLKRmEXhAYH8k/2L38tKgESUhA3EhqGsrQL02CHQqjTPUy
RXniPk4wMMy+g2SSBdmtqtpmYSXnMHjyAdl4eEHDxCQHZR2l3OQt4l/wnS1a
g9sjlTdOBvQzROhsSL1spJFWGV0zXhCxsIxuSk7t3sbt2bjR8kr6lHWrOp0F
7JyvYhW8WuyrqniFIaAcZIxz6pLZtAxpnoqDu+tnYlztgjFdXrGtmSx3fLVK
P5y/Z6AFfGldbyQnDoum1gKVSk19/O59eMGtfdqJIDUwP9IpRQF2QxGBNwHN
M+z7SJrwVynE9u4UuQQodJSBpq4ujsATQ3gFCekBtFIZYVVtXYBhUipTGo/t
fh7jutNLCWy31bmGvFdnMmOwzGHmnfukGNPsAXPxRqKZ1c/GsYmG1MlesBCH
F4YEpy0ItbLVcUR+DmAcY670U7ELOcvwIP9lX5UaU2HZCLWnB4HchHXLAVP+
HJziFZ1r6NH4MaPuHIaXhYIksLXAPFsRh7bpFWplE7dV6Zde5lmsK0gYwcgR
MiTpMI54c+42dAOPJirI5aQiXW496rZfOmJMGONw+Y09Xi6oET/UfDJzMD24
tQWaANoQNwF5nJW5GfqaVM9amJziz4jBPMGghWwAA6JLrl+uPEXIxqC3ynRi
EylDIlVtu4ciovy6nron8vovvcgMljay6PSWKOVi2nP2qDWTkDv4LYaBEJ6/
dAn7lenhLr2S+GktRpDRkKjZOIpBdPwojcQ0tzOXCxfFmQGvOUKPhoNsmcF+
WD8ZoZCov6cXEji8D8mW3Yo4/7exgUnhcnlL6ZyGw/lrG1MysjwKr5tbteji
on8Zifn6u0AVGs3rNsW2ODHJ8r51RLfFqc/CDhd0eZir7nAA5BgXju2kGV67
p+6IwbesYqoMKiSxHPm/b75hVqQUORxZXnNEIIKF9uOE38KdDs35P/Asw8BP
PHb/uCVsKkepdz7CEmF02QmHTE4TcHdVe9vjrUmiwyY/q0Kawmt2+3yZYZ7i
wAnInK+NfCqhfw209bt/JpkTqq/+mNTXvDmYs7NZCFIkt9BJJwzRod4VlThV
CanT1aFkK6UkgG0YMiJISW6gLRbBMp0lAf7rX9LdLUrQlrWfaGJoTgonp+Jj
424vId4p/zrfEognG58rMyci+GTfdX38UABbV6T+HmTnYFYISdMCVIr6uQ/o
T5Af57zZhviR4AgW1KPo2/5+oDbXRMFo/q4l523lYks5AhchY4oSJWeSTHXN
DLgXPQWg0jwhpImrVFNzT7V8fdZ9HmOb5hobZzD1w4TUzUhlCOuERf1hX7/V
ypoVTbHq9wcMq2YjeqFtO3Kwg9tQ1ceqKjOumnB2uVUDhuGkUHwYPPQHVp9W
YnKIrvPqR7f/KPm/ryqWcoVrUHK9teFMmkU02wYaN14Qv5u9wfLa9+m+1EaT
gQw3hEZjJQbG2racoTnQCo0K03EUG89oAXsl+/WxL61yMsyZZsrhb45ybOFi
aIIOJAp6/tnzxPYZxrfn0/LfS0Wd09m/sLauq59PajRZeE6QxvwBF4fYgC6l
A6WfKlrSMDa01KMAz9WtJVOB00c7MyohxGd+zWs+1Dz4ADnQ1k9kPPiWwNxH
9ohlKb34U9DV1JMJZz4h0ROwKv4sy1u/M0OXoMA/W4cHGfxq8N5JCOSUeGE/
Guky4hpFRO8Locz7OlALpTh3PiO2aFS+u/1BwvbzqjF21wKS63NDwV031b6g
twoZ2E9YRiwMRl9dwfLCm7PLcCUnao0f5bJlMe+QAthQUJ+jqcUb2ruViNCw
S/PDpITFkJPd1I+xZIyYz3NwxbV2jHOFCohVSD2V5w/BaQkkdxup4y/1w/wh
dRsjtvEyUUlJ9wCBkyQEhqEIVrYWlsyVFKNioQ3yil/kMPxJDQIFJTTL+oRB
vRb3yYHk1MuCzbbZ55y3S4JQhIDufl4KOPniuhNLykBHPbJY1UuDeYonCT9P
WNChMOVTNfNCkTc2Njjpy/TwwUMjYG1eEsEUR4wQ2OB3RjeGPMVZ/j1Zj2du
kaukgjfbB7Rl0SKKG4znBA+xmen8idON5yahQzVevZgJIBc4yd3XzO0XIDxU
vp1KC+c5lcatyENpc/Q0S4M95QwRaJVT3xMwr8rfPdwAkhEiVs6xWPrp1pni
pq8qsxwF5m+gAJI0M9vSkiPx+nMEuCibX9WAuyX+DEybCVNR93fip/G9z8Au
VhMjjCXUz9KVD2QyTjLMdbvrA4hDVvCypT2n/r6F8puxjPX/hG+j39x76rk6
RUqNMTBr45gi83IkqX+mpxI+FvAvjneR++UaHpfTGUNrir1LtyDowdas2szR
1jXz0DRTh61TH8qbW5iHxuOLBkBGr/cRTaVlwqx+DOq7lu9oTB0Oo1s6Kvnb
y0+I+E/mtI+aMKwm5VZwLwGhonuL4QGmWiFriekQG1gZdZCgdM8M87kIEewx
8oLW5FWfwf89q/vh+Qhu7Vdeh2HrIsC3RxUZ6qtlj/h5UIv5iS+pN+Mu7juh
NbmYhqqir6oqsaBugbGNic9H8ONWex0Ao06dx2/0j93eX17oaddkhnufGKiD
VJ9DypwYKPejJMjLLfRLO5WENQRfv5/D9Dl51Tx3t93KtiRaazXJak5yGBK8
9hU9fwMnrdd7vdIGx0t3IDF91g/wUFlN5EEJCxIesQTebnBiyOqwj/2P3K9V
HgNz1l3yqrAoiBUDL2jFpjb09qLY2ymWcEHWRP6GCsocb0xxbeNSOriQhXTY
5EWIEUkY2jrUaKxMhth7jP7LB8IISCjsMDVwsy3bX+J/rwXF3BiM5XPbIQwD
TGis/maJaUi132lA9x2fXcea6TNZr8+ZhwJSqm04RUsQQtO52K+ypLhZfGMB
fx8SjXNepSvDfbzXG8y0KCRLW8drAadRgA+jhdDivK/Dg4yuzCdf87yvhNFE
byfbdJUk+hIO2WWBYQ20fR5tjZQS4G50Xlsrh6GK/6K+x9uofHNPNE6hMmpX
IHOeapZjFAca+rxmE9CcHzkhFn6R2zULNeP0MctdO0Da451fnQc5/LJ3E/IY
CCtYWDt1aaWOcPUbUaYLT/dJBgdNrgFsHyO7JZjv1KLZAPNWD07IyrpRg17w
usntjuEZSZdmys2tYQaZtovRBl/g7XPCzvHzz3i2ZEQHrZQMWGH/UpfK/2WC
IUZ0HcgQTehYGO6GBL52dvpsi0zO2jughRiv4M68mgjCGlNCg8761HKKz0To
f0g4RiaI2vJXpCt9R2HVMndntt4f90I2XXCDCIp++PQQHeq/HJAKSuAsm4WS
rhmE7nPaqppGjXnMcBeYRDkNTlEqSYUwsnnOfaW7RnRU9ed+oJ1voUdgNMFz
YBBYwgwL5tP0ljSRVDHAAv84AfKMCSrbHPGJF3hdagyf8dZm1n5vy37DBk5T
SntKUF1UYR2v5oMzcIlw5lZWCsCXboa2zp+XvtG4vL7jID98Sufptwzw4SXo
xJquZF11s/OrlEnqW9rLScpKDuLEjTLshvjFrGn2iKnjaEGycr74oUAvE7Q5
1p1oqPMPgZlqIkcQhuvda2pdlPhIXRu2l3eCiLXMWNhLCdAIanB6AcrWRMie
n87AokvE8eEgwZP8GKhhdHf5B83p9pnAs7NiazbuKyPO7m2I+UbfYfitVl85
srKvzTezPy6tXbMJq4q3R2A0hsYxcruP6dqQLyvX2rU0y2emjqqQx3373ObX
Qnqx72uXPaqn9GkZ8ttYI6/hGBj7bgxoN3LTBNgbdDx7wLA4eLMTlKDLsohz
UTYbc9ofhxdq+er/EUUKJbn6iW+5/sLpx1vUJHJfnNIIL/yCdslKOoL1CxHC
FqEHLfXpUNpiNrtOXRlABmGtxEoNIw1G9fu0q7P07i0mByE186uMPfApJZxh
hsC/zSc/f4GAKItHAAugEkdyBENXYF89SSxMcTsZrnDIXzOPlUnHHuurzfPr
yyDb31wWU94GDSJi7RcDWsuYhWgJQlpYDNxfJ011gWnwdbpvntC3Bh+qJCrg
ep9/2FCT1TyUF+WD9erwnsYirXQIUXCuwrkQ9z7QxrZXNKxgOiL1q3fwaGJl
ZBmLnfJLOnRI88uQYxypwMamCLd6MKb5KqDzIP1FDgtw9qVAcj6aNsZGPvnb
W353sVpiVi6cwMZFHNnICeSnVdMxbK/RzALqG9e+jOuc2J419dkZsbzWFbWs
WUwNzHUhZkj39XfstIrktR+851PpcEtI0sNUuDgcdb6Crekfe7MRtFnT0xRL
1AIUt8G0J8v9Y0uhQAn7GL0ONjPquTACdE3Qt+MKIMLQKtCd6ckGCFeGejVh
Qm02RQZmTGu9WckAYt7sO53fHWQp6Wl7fV6iElCKziKeo8G+vKvJF0q3BrwK
Ieyqlb4Ey2atgwwgcEYknSBVR2jcvBFeQwb4tw96/PCO3k12diV+mnqUi+Ty
FDBPMq9n7C0FYGW1YS0YmOnfCp27pPUKaY7RKIZVdQxvBRvKbi83+pACfSeD
DUz4GvyjCaOJ60lPHGkDWr+YMDvXrk6VmfsqwUzzB5mRyJef1/IM+q5UwhV5
PHu6cCmBKv6ySc+ZV/FIuq8mri98tjFEIZpGQvcTF0EgDumw6cZLb4VFWPX0
JQ4i8VO54F9acfif3hjmAaWnZtvZ0daahnkTNxDjGCV9RMn6YP8NiLOzBhuk
KGzBm6OgdMSgMeZY1qVPQtvmCUctELjbLVBh4Yn+bYWrU9ebcw3X1lH2XmXX
53ns082KqEyusHljoizZ76yBC3e1s5KL4yMCJi9L1EDibB3y4JnegAsONrHp
TKzXATltlJy81OGhqOdTmwO2GxSGGEKxWQq3g3/NR5elHbdkcfTqYNlxSokW
xJGh1WA1M7tu7RiYXd9x5MoekK2rHvOOUadVNpmpMB5kmZehg6H6RfLAl6fz
OSqs5pOL7ZJsZkNTT8ird4UAzfKJ9rgAMQNBMTfGYAMU/Aa00iQ4s69hs3nW
bbeSBuV+Bm0Bf30aLQN14jZoKP3ingfjrPRsOLJG3ruPcXihW4mAVQm9ghgM
T3SnuiMpK2iChBidPvayp2DyzRrVq2c4EToDGLp028u9+Iljicb4p/tcwez5
jXdj6Z5eKSXBmv6RmfSw1AScu6X5limZwgY+SJPzqVAePPf8SvdXcGaMv77I
/TtyYZ3iI/M2O/P68/xGtS0fOWu5GKLFKP5RQ3IcXfuktXYCihCL9PuZ1VB3
//1pBwZYlf3MGs73L+iLCUSPzRllmAjLQN1Ebcy+82hPCZGan/vX8KvkHtU5
rD+4ZNtJ471WEp7AIPBf0yaw2bAQv0JA8Y5hyzLoJXvhdkOYWySHWeP1zVX+
MoCF+5Slz5FCrZTY8272GZrtADQpEnp1FlyKx9cYNjm7QY+x4BcCo33ZF8A8
HsKXIrq1JImUN+iTRuM0vYq0zJL933bvqfJXuJ3fD7mOK+zsVPYTOA6WkihB
roTZd6fVCOJ4lqlVB8YV40Zmw3VkFodbOCiyqUYX3vHP4W1R+wZrz2Yi5A1j
UKBLO6yfjTKT4lp4zRpEFFMt6geAWuTWS2z/4U0MS2AuJaw9DJlCiqm62nYX
7IEjw2ii09ugbm/55wiGGJf3u7OFEgWX8LEDl5CEtQum8zvElaCLVDs+Zrei
96+F1IT/kKwH87uDsNsFwZzqhoMg5UEHJJEvThqneBLLnaU5JdHSQQiL2ReD
SC/oE3CfcOoJSrIU2UiTaUcqeFhRjYNPie7H2XLoo6PTvnQ/3XpfoYS0vKnj
QBZ32zUCORxVA8nwyetEdDCcHvshxP9S6hKvYYbnQ6Kz/+Xy4DaUAJiAfbeS
7pVk5gyy8Af4Sh0PLO42KSOdtcbSutRkfhqOydO+AYEE9phSEELxsV650N4R
o1wLcUd1NgZDWvyevJCHo6YCU/rFruzUoIUuPctH+zrGn+gCLG+r1n2Vg13n
yEgduWF+qPv8aG5ViCknvndJoOEoLl8uawXZT6x12qASi6sFJJ2WYpy+S98f
QrOB9OJSB5m6w9J6leKLkWlSyV+FK/ox7P6rj2YNp5ETDd9G4iVj5d7wpn1c
NuT+VCZvNjPcWPNaKjNF1Y9LGhKi2ESH3RQ1UrmTpTrEAG/HiteJHMYB6+kN
+k+H6YcTa0/NMDnPg1B6SsfBBi5saiDf8cbOdGnQWGBb3umeeH4u+/mKEMx0
VYhu9q3ydyJHCiBnwCFqigtfbQ4shbOx8fp0pfkvcQ6Q+PxsydIzXF3t1NYK
C89iw167IElRf23LKfTgTVEA752Z3eNCjqrXaN1KDeoHHajNS32eDb4+aEdJ
KutPLwlYW8otCKYofBFYXigZajI9wSsvc3/NW88F7MQfkYMOm9eZOjJyaLcH
Qe/cP2VJ+Koq13UcmjOKtjAqheOuBWYo94yq3z2rFqXLApNnE26wkxYj4fEH
fx+cTXbY9PLJ1uG6Nw3WmO4+wMRwQlodg6+8YJ88FpRL5YNSxa2pqr1rpEv2
OMF+Bug458I8kuLU95bTidnJfo1cfkYewXek7vKu/HrydgIQxYZPtmwFexGn
4uAIF+vKcsByMv1lsIKUmZLvHfi3Xce3L164bLZ5MkGdMkgne9uHF5dx6ntZ
O53b/Pq7f9m747YstUeMaJkl8D4ca2kT6plTRlvZiKLQ2XbC/JsiTtRQIzEM
ybx9xseREZmuNuelKhvLfaW/MoRyf38Ua7PgY0GUTmvsCJywpPwA1jxCcZA9
MigQSZ5eCcH5MaMh7mvxS2CVs4FXHf0sF1EpO3B/0LNKpE5ML062xGL1KZWk
NOUrBzXwLocC1QEabOjH2N14S/vOj+sDcEpeXxpogarXXStaPlLiFWaOFcAK
P6nbcig0eyuCKECpmcu/u2x6g197bTtbBB+8IGA7/wJHGa50FctgXh0PeIbp
uYXIFuZphdNq416yyyB5KQ9X3kug2QcRIfwiinJkZjbQlAMY4iFdEQFCGAnT
CwRkwjy1zgkStG8+MgrM6wNsCTUjmVbFujKo2wIjugfyLKCTdOLQk82XdC0t
b0rXd3XlSKuM3l/T25ZUeORwdbLVFd0LPM6b96JZG22C0VcfmlV9DNGK8qBj
GJdWN8cIHJb0m/Q6AA8cW1TkqM+3Yo8ByU1DEYS1gzq0aDX+eCCT3ZsjiX4o
SPNZLHBLFrds5DaznUE4vUsnJgC6t3a6UA8ylZWjpS3dSVJb1XXw6BLAL5Fc
WZ4M42JgdPWYWYoT2X3S04vyJzU9eSWjaoGUkOoz15E/X8QndS1WvZfJHda1
vGu1moi758ErC3dswD1jrRqlLXFuocUug34I+cdPAEB+OiXLABIoCZd2EjrV
kDs7ON9Y4VYVhQHJ5uv6nFu75hMb9WNh9MztykqbUWWFJwNwFw4yqkEoFYdV
v/+oFNh17kWW104sAaiCwi3Td+2kANR13m54iCrtZHDjc15ZV257CO5yf0o0
upvEt8v+0za+P0oUWLhnpe+vnq0J1CthB9IaQ9cMawEqq+IeyFjnJCgdx3Ds
iMe/6U5AQDF49wUCHa15Dhh8VH5kLqWkqdyo2EO8WeM2dk1LR+3+yNxA1sfe
BdDqKNGT2IyifuL6AY8+j/syDTUXb3VA9AzEEVWGUBwePXGuZI7Ar+g5LKB6
nmQrwl05h3ALN6aVkHegwrWjNH3TFzmGehiR6cdAYaNJUA1BB6Jh2KRZLl7d
qT32nHtQynnYvSTxFVsiC+zy1qIrTPdvLEQ7a0sL95InLpA9cQQ74Q3fGYDz
gOasSJ5wOOcgU1BjNbgcfnGukc8q/eWgSWASllMNpAFbcCT2W/iJIhzVz+lt
JBasDQjQ/c5dlPS4PIj3yu/j04QvrSZTrO7oV5OqRNAE0ikjaBzTDopbpUSV
ilGYDUPo5EJaDUfj48cZIzch7jqWo2rtGh5o+vGPLstF1yj4OzcyJ0JgyYlq
/do24bbwR++2hjWVFQ9jA8JOeNeWQBwu8nsJj4XDIjODrurlon9oO1hHW1ja
sG4rNs+g2Oa9255oYO3FDvQYpI7LFoodj8PkMHq2FqF5ZVXm66M+Xyq25VZS
B3l+s5Db7d6GqNGUfen4dOAjVAQaBNO1gjX0uxqzJAXsKwWOXn6H1aj+gxx6
JkNAHPCj3634YUZVfEs9krjCjFeg5JYc0YaYSHOIoTvmAo3T6NTu3M4QvzmB
cXXe+inWEd+IBWgsCLh1jHAhNEDs4slkQjonm2swEDBxC+Wz0IUsrvvliGjP
7RCdmGN6gBQGIuyprcRLlGymITApQVL0l9PlVitzYCW4qOPWGQYZHAN6CaUE
QG37x80PiVVXD53OAxp2uMt9R437HjGa+A9LkyVITc7zD2pW/o2oCrHeTlJV
95zjy60mm147cjZRuy0BVuPqACDEl3tdrtkvXUyQUG9bsV3mTkiupL2Tj8ez
vu+spl6SR4SVFaUomAYlJAfHE/WoKQ6OxI7hi0Qm5sUIIsehCtQU02qWH2IS
wJC/Cd8WuXfxyHzSIK/orPG30ZGgArzNKfIbx3DeIohSyASz17kKplxGVPyP
bABY3v4OaRMTgN9rBXCGyzeGWoavbM2QTrhXSOj8WrKj0P9dOcujTCpINBMf
Q+Wv27USFo+WMqiof76bUZZvz8pjjy+Ip4SbB1tjksMAxVqoQKlSZ1bkg3cO
0xqf1Wv3+EL/oGT7noKoV1/v/4U9iMtHP8gkcebnupu6j785nXSytpQbEwKj
fSHyK5InJOd9G/qexDfFXlVIaQvn3IHhNUkzlJqvL+XA4ZD5R42p40nt/oPG
fD7wo+8dezrIed/+4DsaDTSp+0cuePNQm8Nm/HRMKLBP9WbDC+yZQYNHlOqb
4eTCtlRPdBGoWaiMOM90nDOYyvx19PXA/6F74OzvHgHKcl2wom05Z9XT65e8
o/8eFnAvDZlo/SvwptusFWi2WNJG9PvoSlflNqSA98uOCBk6hJmwA53O/5jg
z1qh8Q2x+ouDZOLELt1UG/SCropWkMQ2EuOHZzvWdgyZJeWSDEPZxaMpv/sU
YXdiE4M+KZ7lkPAobQvw2aK/2oIXRa+mN0LXFFBqdjzA9B2ujgfZ1JpEzTNy
nCoe4NPUUNXeuODza5yYzoB12Hu8Ay0zFOhCU9wGmq72ipISdpqMrOSdPWFl
hrtxTIaulvfuku3zsa9eUevylv+jH9XZSyyuJ5NB4IjVorBCqaLcUXKKLyue
xHrY00rJSUU6wZpv+eRaUDXfILC6xD7AxKX11VgSbOzr4W5w6+5pzVLIhJhm
HcfDUA1VmlLOXABsN27u21P2TwgWkIZmQswFv/aBOjP+UaAWWzQusv9Iqxkf
3ec7QSANC4S9cL67H1WxrcU8bmtsD5G6pu/rlG+4FRbeim30G90D0j2h2/iw
5Rs/TMB3bpLV3uRGE0bIFmIXY1Wb1DK7qHBi3TC5+4ttK8Frc39xaBr8lgsj
c8VuM7WiuRGoifpf0vECYY3IGbQa37rVD3k3Yf0zqzyzEw/TQrmePKRpCU7m
jt4A2ea9vQ3hfgQgPCU8jp9fRw/glQnfC9+XyUAGCgtGwmeIMZzbAxJge87p
UeORcj25rtLZFwQby3zrTTPuGG91wcf3sejTtJo2VVuvvowYk1Qj0xkfjJy8
wbw05vrCr4d2M5zHx8mB1mroaTxbF4ENmfm7bgxlkJlSYXKMkmq1dlK+AHLG
adTtoQA94xxXwmK+ZzOY+w78LPB1DoiELIceyHDnYzn/IciBuQJnblWdZfQU
/KcGi7hkZ+E8aaoDyOsrtns6SKwrlDZ4o+84Cl5Sc36RsPWhW7YADvFPRKO2
B4WlVHMpfp65tDX5bELOSKXhxxxT6itIpsgBlj77w02Jo909XUQO/9sPQNyv
jSOMJ/m84DJsZaE1tXmYRVbjWhlA8EK4YBOU/kTKTn5AzcNVEd5NP4ytqvJa
0/A9fIBuL2/0RhsH3zt2ArhaPGTz4cfCOPjDLMCiZAPq7P8w7eIsD1o9tsJY
31T7uk2Hpl9wtLpoCBlFrRhfmDmfleX/Fm4IiIWq+BDlFJk3oHI5GcVHqstN
HVZTm7NGDplHgO2rBD8nEjB0IZ+2xDsIy9Aid1nzW56oO2OpQuDXpGllITHT
uFE4WhgzMJG6SKffm6FNkLntGWSWdJrmXWZCZ6chm/+tkqFP9A+TL92+cz8k
ZSV6LqOTOYoi9E3EmlCVhqBdesEL+7ve4AvEKzltEFoRKRuyz76LXZ57A7rm
wbrZd3anRB/vxk7+W66YOYsEv1R1EYzRNdaHqVBVfcIy1a/oY9oZsSk110rA
b9y7Az8cVFhPeFYpmQ8ZYoAWq760zY2UIRUgTOaaPQMeeo818VZ1z32tKWpo
D0Pnnyr8kRHsvWH9cKr0R8rhAc+NKAIsW34WUldZa9Dgw0uUQm7IyOk9uVg+
rKw7xxCHzupqQ7xid1a//CQdpugUK7UPVlJabVKzvQ8JXqTxu2HPQ4ERQw0A
PCZIEN63NzIINcGwe4WGggwubsFfK1Lt5+n+iX+c1A/piQRNxbNPSKmPFF+m
ubdEQthGIU9wtN+hBdYeNfKTcfCfxUEGQofb+yVZlwI/z3RKtqli/jlehgE1
ulLn7TT4dIfuQqBCuBJiL+KIROQAoFwJDpnAhfETt+epk2ttJyDzEqYnSEwg
Kuz0I9JgKj1brxpX1DE+WVTI1DRv1GZGwZMFg1nDHR6BmKMnzx2yM8NEldUX
dan+DLpFPUJqsc0mXvajZfT7EUqzGOQjM/VNy2ydplnE6NR1B5nYRgDS8WnJ
LRQ9RtqWVSKBQsk6bt8VAFomghnPtvtztNTkbl4GmSEjSzoLUwMbKclIE2wY
bF0sS/jx7yZqaMJ27Cuh0Jd5mzYMP905mYtSZx9Ilst5qWGJWRRlmb8Q7Ro1
sB4VMkZePXEQWZaTIb8qB4BiiQl1bZ3qG4QQI885UhPoS1F4Ghz7vHMv5dRE
r9mRbnvx8KLh3HW2G9M6Xypc1+eFEk6Yg7Erx+cc/gGMKJVvRWg7fxXle5Fl
COyTWNMC1y1uld91YxWWoVjBk5MUuuf0NqoL+JYp2OzmdwDVvFYAilJUbhzs
UaiA56i4AGbbIHY1YwOum/cX0X1C1b1rCrGQUbn2sLU6eoE7rKO07m+m6RyL
LzSxrb7dyxVyqopHc4+c66i/iS08fKWQi86WEdTpnPMX2O7egF5lgE5IQveo
iIYJpD9BmRzuyZqQagmhG29+P23cCXZmmE36dZtugh7tWLI409Bz1sFQIV5L
s/EQOspjIUNtCUovehwF8ePXXPBZDOdDa3+G3PD3YIIfrZO3LW6IQR398hkZ
IZscqM1z2IDhmt4Ee4XJmsdUD69LjGOikniK+Yot5rijxnWAGJbO3USS/Qpt
re+tdS0hRZRbnuHlGiuZ9LnzDqnFtTLKTDBqd0Tzsk7B3ZOe0MXXdrhUE/7P
TTLflbtEq0sNtJGbMbdR+6Fbc00ea7Mjy4DDaUNt22smpSnQv+jDh8Z4eKrQ
q27JvLV9HJ8OXI/tb30V8Z785RLZOvDWYFLrshdJDkozCFfP9H5jbWfK0QUv
C+f1JgDDNIlKUvNRnLN8LOI7nCqPJveJ2F6rZt9p2ILRUG+QdT8gLeu2qKrQ
hf8To8DTNb+vrSLuL2sB4wCc+8izzpHvKpMcNHaM+HvAmS7SG5w2mqFDe6Zs
O+2dDH80aaREwFaPJbSeSHHHV2oSzo4eqpB6E3ZIqZCqHH7oQHJXCdw0ugnj
7S+V0tXy9i3Iwl4JMX3u57TzvmNX9LcMQfIPV6K5RNq6xHYHkHwazFwAiR7L
wrga9Gq1xmiePi5SArqwaD7vRx+q8GwQV35jyNQcci5XyNwkzGw+gerN7Af4
uh66n5ktYjk7bsXMwJmBGiOtfoY8czpUDOrcWHcs2Gbsy30Hx4/y8xSkmbeV
u+0N5ksZl9kk8rR10vuigmR/RZi+dQx19Uoq4km82IBPRAGXdordfgm5ZPp/
2ipJwYKCejxrXokuPBW20Mto5AlQRMhhvPF0muFa7lFdiOTV6GdQj8YUQndM
ryUhPV4aEto1o35EG6AqQOFFxTtV9Sg476NXV4M+GOWrBldn7rqwjAFubxxB
dtEkFDGpS7nr7VvJ0kjWmg0BrcvX/58Mnltf/X6D3AKADRU8IavHd0npISWH
dbjkdv5n6+HAhkJi1lBS9XE0vMDQPshpVhOQPeOPUsYqEGW4l7NzMq2rBxLy
Q8aWdaNS10iPlQcdUC/q7lKhlnaaKtCj1VlUpdzxk2EJuBN62Z+TuABqqbgt
TDQZe6r2vl/plavYHLeHHFjq/CifMl4hoVeq8XuAYxZWzCUKuo8wolbenuOl
LqK3Mwc/vDDpb8TGD+94CYDyInIXbGAB9kZ1P577j6mLBuMrY2T/iD5on6Ir
7jCUP0VV0UYrteWlIDLFqkG02cLzMRTGtvNnsr2A7Efjbpm3zBN6plSP4S3k
oBU1o1ViHCbSH2oF8xgZvWoo3ytQBWSGFwNGtduiKR9HYrVYWMw5+S7pLYv6
iVKhJR4dp5ekV8Y7e+JsgkuAzZTQiF6v8cClTorwcUHTfe5s01Y7nNoQRp28
kIYmVc2gKYmbkK97pgAd/qjaRzcHN6mZIsLDMttkkU5DNsqFf40xoLf/cnoE
Y0dsCqfMTqAJtq+kQE6N2DPRz8VPp0B+rFYIHazaXM2d8LZAEr3S4hMrb+2A
Q+RqFlbx66QibODT9Ne5N+bO8qrXsv8p/xWj/jjftPelmr9J+6XSf8AO+PeW
2AKSoAFVj0xGnzt1B1nyk0j/86bW3IX4L2k5+5G99gRFTmDHZX8j4AfiexOB
3+xUSkl//K9w5sd1akLCGKCLws/car36PAcGAwkIwUMcjc+AoPLrRAcpxbwa
5fsUl0tBc6yqKXhG9KKnArZhVA8wb85waLAbTcZrfK2d6ic32IudJyB676ho
CLkFWMn/zFgAGYl0iYKvgaXtWbr3f2hUdFVqtB0D1T9KZPUDkjE3PX6IIvav
SJT/35CtOuvNT6yHIlcAQsRiduwx0s9cffNtepNoCbIyPXhvkpk2jMGeU9Fa
eKt9O/cZnfPBGjfLl9N13xOtnS8OH7ColDkUC+S3upqw2rQ9sOB7nq/eTNq9
wIMFlOX+BLQ6j43V347z6s163oaQG+eYsE5F6Nbq2qhPNuFVLkBVjmeaNi0R
4U9rAP0eG3zCZkfjrBaLuS9QgyRVA3R7fGpyUAXiLmj/QjDrDX5afvBAQq2y
wjDN8qG7nQgIbpWZj3Up4LaE1Pm8OH7w6nzWFtD/Mngucg6FiUHNlOjWl1Yj
XQzE0pKHLr4MMOsOpf9tHhS2KwwpFBTX1lqDKgt7hNr9ihFZKsFpHjbCnsJX
l0G/vGdEcU3PpOWv2Sj1Rj+GmWkBtEgOYvteiGKwnBvLWz12dex4LZicsxHt
cE6cGpD+trKbhKSsZ6LbMZ7xGL9v3WBGiJJiaQdhMGTqwdlGcwJrp47VvhQm
5k6SKxtYBtTMqxmb3295+nlS+R7OMoRAE6pglxnhsrVBdWny1q68AuQpex8S
ZsKUm7xacFsCjcGkmbhJ3ego5/4NfkqA8vibRlQ9dB598jPCTlcNDC7FbAQv
2Qm5vwuvNSOYb1MOtFXsv0/Ulh4Hr7rgLKro3xDhTgaHp3LJHRaSeJ/fjTLH
YQXCjwDR2ClnnYl59BM2466M6pGkQhfF+It9TOSjqr0vcibl8bNF9aYo7eHN
1cbwB5BZqkEuCKuvbxpM/zwi8Bt2w6ipsJ9SSAIrthTx+ClRUUj3GgXW9I9m
9iiF612nELPaq/N11pHIsO01ioBNfUAKEhbgPJvAjPEMOXYulpuLfeGQkWv3
Oc/LoKr/hkac2JczcKHgPr6zyDR/Cr8+3fvS+ElVbLVEx5h5ybyeKBBB8lHG
2oa6Y/SFraPxoAX0d/HmANVoSTytpZPQ2sxeSom/zRF666qOccAdZf+x8P5m
KCOgFnCQg2W9W18rxwSuqsr8E0wJLUCvge/GkAkb2iASZIuhYjOefgOgmGF6
CIezscvwC65kZ9gHuS9uOTZXqixPsZpjTBrhV3gtYCGwNRonyAq8zL2xwNyu
Yp+zHrBWEsHfzmJ7iHXh7uI47wSh5xWY/P3IrA9MvHQJSzuBxNOtPtRPTTE7
WQlNdi9BvPCBiXcpi2+JVWlvyV44bHjRAxg3BL/aWzIXwrVrM75Qv3UX5nS+
3Hx+PJWNJqqitp+ItkgdFUHjXv9UHjgoklGdgjpKw1W5JAKGbSpcqZjrfU7W
M3laAg3PEQ0gwoemtD4CkwwWOZ17WLQ6QftdDu1hkvCs5clZo2kGIljYPTpo
NMwHPMTMGCfl64EfPVod1DjyyIfLHBFZUZRJOsiyT5z+Mn4sblFVNa/y7sAL
1GJmopm0d2yU4y0+hrev/DGH0pC7FwmtWY7C3UO5lbvA89bIOewuWNtRTybZ
tF2QfB0knxGo74heFHdKET+8e2KAyvnt/8kdviuuvnkZvqJZW5Ze5sfg93g/
Jw0Aa+R9I6zkzy0ezpj/2jupH5R5Hi3birvdy/zYOamYU07r1GYXACH03TR7
NG554j5XfSI1GpFEmkMXn/7fvRM+HLEtyXIoC43f7wXGQ3maoHsm5Ie4vCc3
ELOoTtkvYWZ7fLfJM74xUnYiRlr/8y4BBgpNafpdtrt6HRupou3tveOa8cJ2
pQwf6m1FesPOkvovNnWONX9YNEUC8LsJe3MhBz2AjDjTJcF5Fz1hOOEkjIBf
2YhvwQNrQKYuoR+umdCYkUigyK3NhTCvdn4v1tzJfPYXMek2LgSWWBVOuvMo
ft47DAJoQCbpdn8zyZHIJqH/C4e9+JdQrZMWxPk9roJ9e7yB0jdRvGhItjHJ
SteBU3y6bKSxUNpohqeEkuHaTGb26yCVqMxlYjhufMcersJhX98EtoOuFwQK
hunu/0pReIlKIS634QyNJWnp3i0I+sdTgVOOoFJVAqRx8p2XYq5ozAqrx+Rs
taxeIhm2KWM7tvfM5KOTk0W2+qVLScOE0k8kyjVnJPsr0VCXIvJQtVXWAgOh
/Om49Xu2SW/mPwDT4Oe4WIXg84edqyfrD+d7VjrDKo0w1kiTh8wuQaGNZi9+
aB3NE1qPMrmxJ1oCJYIa19kd/dWWb1LbWUL93MIIrwBMzTr/9plzxcjECUMc
RyQllZ7QG50wYcuxkDO64SYf1OlXGqcFMpHQpIopn887GR6qdNgEt0gexPD3
hEyN9bOtAqMGllnYs5bMdSMh9DZI6wqzM9+Uu3dGKr47ggji8P86B1oy6zyl
1wEaOl20b1qgMcCYYk5E5B+HWMLd2btEwLZgqHC5fSM9zXKpRSvfaq2WPwzV
I7PCU99vhkpc8HLuMfXaUKSMKgoxC6LM8+SQSafK2LYvTM5jwe296CdZXChM
JEY8FXrUO+x51LWzMZS/5au2tsokLRS8dSIeWg055fcjOx2WQ+qM0spj6PvI
jnd0ga2HK9rZ0j3cQpJb8VW8W686d01gAYPmMlcdZ+TmXFlSboZgXXhRBFuQ
LEv7PR+8l4FL+WfuvSmOnIBRVUpvDTAfz32UjuYJMGHgo52FTH0VvusEg7Ma
z20BbSRwpnXvIix65GkrQyjdC+b9YfplYZMXjkUow27rZ5x+TsLoivifX3Lr
h9D6ID7TaHu80jjLuzKbu3kEFoMTjeIBr6Vrp8IaJj/UbQS7qNr6feMGXZMG
SfBU8IWNeIt9j5IvkbZK/taDQLdXUxuJeL/VwOQHLUAP17qqsH+8duUjYZRl
mYyex6hcXKybvdqoRI8pHLkTZRqb4nFyYxBIHsNTvNQd9/IlACpfl2ASpmLj
O5gT9qjLHiMn2SdgY0Gz27bS+ZTM4hNsOFESgRGfOH69N2OrzydgLW23h88s
GTqZnsHMN/UEs4ByqF/TXmcF8AzX1/61eEpL2lFFssmT0IwjL4vCLPsl8+P1
52xQUDbV66wW0LSdUkgl0LGQJlTrnG90QimPOXqIFkt6rYOvhj8zapWX4Hrv
hyaZ12K27DsgXvT/ufZs4u+9wYdi9+mkrUvPa2zsNi4bFAhjmsOFoCNg9Kmv
yn6O37IaStjMXxOeb3ri7UgFs5PKt5zcsOz/Z9TGu2YAVwVMJWTEjpaCHynI
0D3K46jS9Dx3WMVHh8k2u6H4N4Mq4i3nIdnsVMQC0FmcOmn91+tbFFPbe/vf
pnym5jPjKy3xW4rIipD61NOsSDPTm8RuoFrclsrOi2ECqGOebP6k9n9ORAVs
d5IeCnvhAO7QnLY/WY+efV6tcHdAbDhXSVIEUBSllPigjkEKKzS8eQSihyWL
uKqQloaiFBrO3/t4bFdfQBQJR/5wOraXe2Df3AqsXn7MFgT+FeOBWeNX5IS7
F3IGo+7AhQ0jRJ/1RkJSL4YU49OgAnDh7otd8gUBWx0yx7vxX7YNJ4wMSowf
6Y0IyJhn9bUvGUcB2Qray7b4sv8PoE3jXm7919bY8Xpg+o+o3Q+edMSO+JQ1
CK1AXwqAy0iE3YCcFSr5Zce7Vl0HkFaEVB6sJqRMmVt2yQJSsCW5LzGVPmnx
CdVLGJoVK9nl6hiyrDPAPYWWLQ0wTcIXIGJTbj361CAO4nZgUJBut+h1ZFqP
Z5mHhvshBxtx06EPgVvSsSCJJyp61E7Miw5JyhrSsDS7O6W1srGPI0TMwE9p
dSluftHRfC0dtMu0KOcu7Qqp/Dz6Map+EJ7SwchQKCQVORFjyf13IIESiEwS
ZU0+6vkN2fWLe6YnosG9x2JCo8y5Z+hxiRjwblX39S1oSd1gpzwrobm167Hb
FIvrSfo/SmdGdzmZ1ODO9csSsBoj/L6moitQxIc2liBw35aDHwPJihQHbuBa
1jweFLlHp2eHMBkzUUw8WJUnfQxbIbrEVnOYB2thWJRW5ZScVXrNaB/PJU9+
/dkKg7VxFtMtUf6ffem+PNVdHcnxq5qjLMhpAtipvlN8TJG97vNLGNGSa+N7
eePSW/BAHxgwZ3/pSbxDfnc7uibPa5g94rIvMDrq9VRMY6BFcg8sDiCC9bAb
6XvlILg6lMGlXol7HuF/41nLnUeGysWeIlg9g2eY03Chv4cDmpn+WuDNzljv
2txZnxJI7h4eFv/+lvHzqJikdN6mn8NXQSNJKM27sTXkqINNBj4DIyIYqXIB
5upc5fy++n+Vh6L2S32EpTLZhqaF0+FZBe1xpTSbcqG4yR5S+nFIBBoV6vf0
D0YEGU96lSFRtaZWW1wL483Yi2irR4+61/Whe5rIt9mVhfXjcAhmWt/q9I8l
Cukw6pnG449/e2IufcyTT4tECQ761Oe3itY9wlpowbiSWhiXE5vLRlIObeNw
TMTb4kKuu1N8e+3L3+qCxWxpeMiBXzomq44BF8r0MdKo8DZNSmbRuMgmUKyf
0ZN1u0YxbGwDIFnWtBS95J2elDJq7yU9kGIdroRcXd7QPgcWL1LjhKEGwbXB
7gr8j7YUDkJ4p626yiytWvgU9XvnA+6w4SnNzXOgUGuPP3IvKcmFUil3AvWX
I//kea202XfdviwimiwouOxGXYW5dZXKd1ypboP5Tuxkq95JbomGQNpvFE3V
oo1uP4EUjxbZa7Upj5x2v11n8Q0DVhhGFd1oX8q9I1vyRtb3sVtccuC7WmCb
DFHZlkBhYJGwxPweLEy6Xn1+j/tyxcXD6UWwS80BE0kpZFsswPsVD12Hwe6H
8jLQgd2msz6FtUuvHgbn+LyN53WWyk39TysXzDuuuDuE3iIk0BDj8yNkRcWq
BenwgjbuYI1J1ZKA4z3OGmOjtuXfhMd2YebUKy72HQdZFtZtIuWO+MqPEpVq
q1N1wzQmLfI1q0fznRqA0VoVDBHy7CTFJjDu3fDNIx5NhgJ+aVuk6c88/C01
xRBUD8BOES2wy9dx/bhzh5EYlf6R6oz40D//RjEel0jG4N5/mAV853+KsDrz
cz7LPeX+izlr+RwhqhztslJZpm2RfjZaDq2qBTJTQXP7AwUNyN8YzSs6+2NS
TNjAsnkWSIVvef5aKME0a+4xolX5dMpVhIMbOfYBMvFEw6/IePas+AEtYJzl
u7lQ43PVYoJ4DhMpv/XmAfbVuaCYXcFnRBQwvSmWhm3tJSPwX35eU91gYzIQ
H4QNMOjqDIGWO39PWw35Hy18NnBd1b+BFQ1IO7W6nW5oL+BkvzbAsSWajOJr
gEfE045oLP5nc3fdvGx2erF3tWLVo7+AXbKHly04liIjwzk+c2fZaTVVB2eV
b7D7M/A4vbD2iXozFveb0hZORCzs46mAtnjhjg6R20+pCxRNYEeJPdNweiy+
k0R57YEIRQGNeRMoXKAbIscAZvFvONImlsJniYSALLReJnTu30bgbr4mYWES
pVTOJvBn3oJwxEXYk2D4xtUqVzML9GwoDT0zlLyL2y2X+8yepaNeWoHj7oxx
3JTLNARWumTao7C5wS8OuCZ3wWLGJ/fzP5TsiajPj6mjABNH4j7UicYb1Wp1
sILz2/CcNJ+55RpTFJUkZBwdm5XKhBYIDIIMBe8hcJQaTru7IbP44M++lO/z
Y0gSACoXcWVCVvTWp1Y4Nasm5Qc9N8TTd1Qvv3z+do4RjvlFgkgM4zZDdvHk
3AzeVOwGvceWGaJB8brZPATUcW4F43IJ2QfwxoXPUYY5DhNODSXcvoEqrVhN
MwWrUea+W4iCUYyhI2/iyqJ5Tj8rBEpr9ZeG34yqj9Q0/G5sjD7Un1anYjBe
g7CW2FBWQw/Q6WFqPHD8VAo6E3n1rcmpoir2Be4X1NGUmOpywDfGvpBwRZCc
ot1VfjwNqM19+A5A4JrrD/daNB5DKmhiPfUmlH9KsmKFFxZvlvBhX+uNH1Vf
Uu2hasDA+Vt9sxjedwTKJftG1qeV23oguv9QHvfzGMnBJV8bw+zPD187R4du
bRwlfGmmQfQDg8LokOHqUqliJaUlzx+VK3jD3PECnI3e7QYoDol8ys7fe2UI
QIsYFtIFxBs4OvbGZT7owwnkW+REXJkQ0mfcGG3ZC3QktRy9O60hl0Xs6abP
2uqYXpPhHpEl/W+ffObRUGvc5X/7i2lFeyyE/QNrEHsmAQ85mbSGi7ONlMGk
f96s+CXIh71kGWhqZxatizBT2E5Sw0M3KpdXxcfSzgMhXTz3HYde3+N8jjdc
USK160eLrecXKQTz0OjI2FHuJJKyOlXKmk4t9pN4zyCXygSpz7Kw3gPQpV8t
Rw6fnoieU3yXH3hkrrrc7mZlELEB1UI+EA8hSM7jS8zOlskZxOnKHdNp7/tV
XDM7+u/Rw0GkrRQw+LudwAJcUnSIbxad3AbwC4l2Evx01a8eb2BccekjIDUp
JQqWqoIXDfx2OsbQj+tbh8qqfFZn9cZO4nk3jWtsNNkxaFirIbVr3p48jNOZ
mjNLt5ek0mkSc22pmM1UbE+eqeG21lPLx5lREK2aOLlBc/ltbY6/thNPv0bY
M8UFFf0UCvCBWlA816Mm0RSf3tVdCu6gpPng8Q1U9rAA8zAJDHSLZnQOIihI
UnKsiIN4AejBsRmwIqMHi8kFg+5rv7tPuNR8uimI+HL0nfhUDYpCwmR8mTJW
tYkrwlzAj3tAenFygUkr5Njxpz+4d64LJzoWG6dvfEUWJv8jvXs3oH3vXpat
HD1uuiNkMziVCUbASr2Yhk6X7CgqUJsd2sEOXdsR1yIc20GgxPCvMGk5XoTk
RNB7/BcGJ1rSODj0Prq1rC0Kz5S3+8ItHKkHbaKJSjiKObcKz88vFwsOUU8z
mfnt9xcwJlhr5Whz9lIK0RIxaDLq+iUk77Ciu318g5U52bCHfHLkMzxlzGTs
1KEfB/dB3AMK9OvtuvjaInASiI8BN9wrWsPd0IiFixBahttzrM+7yDM0Iv6K
fJqoZrgPTrl42ipSsCop9kGcB09QXHwQMDJL7wNp5GUBrmQX4GIPxETkM8v2
LfoAr1bm13Gxf442gcmKIp/ZqLW5qTHihMpQJHytj+nbZDn17Fp72TN6CZe5
aekksknkvrNrgeqzo90caThZs0PzONWWg0fKHrYHgTYqq2iqCfE/XBcO22Mb
eqLYBGSU0APq3hFJoj2pBXAWsW4pLFxobNqsXIZ3XDaUGRq4fMOTmn15Aont
CLneEXsJT23El7zghHa/+peKM/jrCyWPkJQl6iBfAoGWh700k/12EYyG72Ig
uSFfKsw7Gm4ZU7/WuPgWhBWCRAhuRwtPwDrhOn/fXRTEvQon5S77+/FOcV8k
DmQcFdWkd796H1ZP5G+uCJc37sBw0P9t+fJKL64FI4rU/TWSU1N4zX70S94b
+Yu19qwI0yMG/L0ICcceBoBn9XIA5B6UQqPXANg9T/h9cMvpMqdAEZlNMqdw
rEoN5LGG/dcoqcszSHD6FJ/TjfWcAw9D754PGtYMbPRk9Ly+GXlzzfaY3MRC
kpZwo2Rbdo96UenOJRsGXpZsyPLJ56XLPWrp80YI+arCScTt5eskKnIyjkSL
mut9MSXmFuq8sOCyEFzFMiFTNxAzrWRiLk7QP+4n8QEkLFeNMD65uHcmJhMZ
s+PD6/3zzVy0cXjiH0yGAKfOMZ7AT73XmGXRnHz2XERNMpnPvIOfdvjh+QAr
AG72nNb3h+Z0Q5+K8b4Yp3oC/6uum3TF96u8gSmdX6wQhpMuGmZzKpQuYb2z
9LIWI0TWihC9lf7sFrzFrm7t+TLIB9fuglRQBCMAWPgCLeRRLD7DbkFSwwjR
uAQKx2CJWWJZQZCxWdIcI1nIhg3jJ4MZcoc+stfxTau9kEdQhEXE3DbwYZsZ
os3G5nTdRghMStUnWxCkur6FkwSDoB0+39sAEJhMjXXCtM7dQEhP22eqleZj
QT42V8oYR8DKDUWSNr8ogOy7CcdIg4Yp+YoasVSGQjYnsYyfAtcFp8Ls9YHZ
uBlMEKpBflCJq+j/FXS+BHNMGwp3TsfBAIuK5CY+mr5+c3qEJlyp/AV04Pxp
VgybolzzPYYRw0ya+g5bWA5SRT/2ojMRW1fXT27K7B1CjQTafyVZmWQjUbbN
VcsSNiXwcgoQAY15v997AYtNdNDRA+hAEG+PjFOld+SRnmr5blAtHMqVm3Zr
wqbYvnwx4O9TAwu4i2Sr94JweKFSmRLoMCWQOiicGBlfkRDEJzjtUMvlsgxd
8ffwl7SUm0n+7ngnDYgHF+2KeNsQqBLcURw1yiOvYpujiUQL/EFb+/zhWjjM
DwS/UjQfVnThAZRCQeNEyon2XpOl1jYXzIuVxkP5/Os/iUTgJDTPgjh7utwN
ND+8yL76nlo16mQHcArCdYzHGglg+Uconv0uwRIngjoOa8M5QndYoA719ewq
XaazBs6ck6f1MPgxWNg5G8UiGyfcPbPvX8dDbxVNNcTHMlTUGYNJc2bcg2/c
nQbioBjjB/CObEVUviwXxVlMyNpqaFHH6HBM8/w/8Eo6T4CnzoCSaeirIIAv
o6BbsNClBLwd0Q169z9azjs11tBwg8Ha7SA3hr7e/AoRsHqkZfeYyWyutPXN
8ndxk5Kagef19bIDYXlBvt/lX34e3iUHWIq/gJ1dAuku8vt/BmXGiTpFgfEA
EqrgQ9H4B/oQtvflqPGThj8Vk+hZFeuL1TypyK2RyC5UEvgPth8D8syWnWEy
XwQAGSUrUr5lWEL4s3hQQABYIopbdSG3OpStZgrDIsOG2RtUGJwjJ/UZptCD
o8auHQE1qfJYNRHBeOfG6wb7BOf2hOjPq/M7zH2iRgMhiI94Egy/Jvje968q
ZZdrakEu8KN2gkIJNzxJiNenFKBi4wzkhEh4TmlaDW3E2XdiFRUpGYKYIRji
HTd/bbBg0QrUzDcMt3sW2wkjI1la1Qx1i0bfsDEEQV8ZoHUHKVWxPrMAzms+
e0Aqf+VB2KlR2nfnQKEC2WRvLXFoy68uRHNO+uYFhPvm3+U5Z6JjCqzgvbkx
cULKU7nrIn/FsAVazYUFAQu3RnWboCqrnRv6f+CViwojxBZbioJ7skH/fRVY
anwacdeZbiJ5yHAzzz5HOEvS2DyLV2qi1aOdh0PEoaJZMj7nDrsk2hZbZs0v
d5Q+WkIM7bJDeuZYsumVwo2VanrD2K2QHZArCmhu2SDFVTu24Q9kd1UNMVpk
FHmIlOKEAxySx/SoHnHZkJtOr91wrjBFhkqDosgYgu30SkZWgqvxjwoR9YcU
ZsIOqnSzNZuWwH7AC6xWMo3Qx6VbE9C/e9xkDZbe6AvH/UjpKIwVYbkGu65Y
Imn03BXyhAWdbWYv2WBREGr0BmHEq8G5gpVJ4XAUjP7AperqWkGnjlCSBPjL
sCRap4EIkO7Zo8B7hF8L4Nx+Z2bk32cSdObU4I8DlhSrG+B+P3qYUHJc2ax2
Nje3irMGqq9YvvAXybfeNobERPaGWT2g2eL3egGb2SZc6DZ2guxhCf5FTFTb
z14FIG8wRtpi79H0rtsgsSUmhNp7unrmVwalRjAXuQlqOhkQiRccZSsnwTUu
vx0qam2jQxMONqQr+GP4JadVNsJbrag9sfXYth/HMpQg/zLc4gZkpLusz5Ij
L66vKOKfyZn6KHMMv76f8qo1cWWVmmRn+w7QyuUe5k1KXbAovwkn2UDEylyy
3/g50YAyrxA3CMneFm+2mjzdrznLOJ2FeIUDBowyeEJWlAnKIEGSdiy2JyaC
O/xnUl+4VrtCoI71VyMP6ZgALkwB4dhZLl4y66Oj+kQF9IHlQx5RJz8T78BC
fbcByWXVIycCEc/wcCymQ1rrsOa/UjkGEZ95xiIdt7WrWvUjxULENhQw0335
gZ37SGd5+flpzwKrzdipphkfL+COZrQF7vFy7XVdCHcAeuWqGcWppLJDegCD
nN2289i8WAHAy1pA4Jd8TILCBehW/4d3uU88LsFHvLUNhe7NeiuydkaVyEPy
dWC8TfFGcH2ACw8pTKT32KRe8FskQtrW9viswZw9LpBrczBgwyiIOajcKF2V
MzPIunFoAZCE9zr6kFjL7Gq2/LtahqJsKB/ZfGCzzbsQWtEFqXlopvRgrif3
6uZYDupGNQVSW3Xa5/dMehGFkgTgql6RxvJWCYYRdLFWCv/ASYddZZ2r6Yng
RmI5im4E6vYd9ralKAaQek3t+SYl15loCC5OerZ99hhMxrnsrR4RBtZ0fw0V
5jeU2g4Q69sCW6xuKNAnG+/IS+IQ6Q6ub+G4/uHRwtyTOFLMjyi3KcTcMf0e
1/Y3JW7vzv0bRX6zmpxOMLLt0ftCJkdea7q/PA+efPBgAAg7nPNkb+ZS+I9y
bcVC281RGBPCNU/k/Y5K3T15yjEYC5qs4hEiNBrhV1j/HdEqB/WjMxZOX1UG
7uwQVxhqJ212udUjQ6RgA+S6bH7KrfLHdE245SB7GMHh3P/4pgkdgvjBABPI
GJdeGMoc/w8BJwcC35dct7SkzPx52Ld90DVl8FCMY9Cdqbo7jC4Iu3Tl4CCj
yIKfOMmnZioXzCOuyVEIXtmiX7se77PUYYqwQvDflH0Yl2AGYAD7hbhpFBVs
MuDZbCMyzJBvUX4KFtfvU4NOOSUDgpI0PeJfvUT8GToKshWkOw/xCVwqcdUj
2WqjGXLrFsFommaXNcjCa4yQBZbufvy7pzNdvm5S2ztVOez1d8PEvIyr9Syn
0ZoMxU/IR4AbAfxRBPJvEc8jCJdFewYwITzg9ZGtNdoVBg+J7OapgBa8eLMs
uP0dmHeznuh4UhHD+MgbW5H/f9CmUiq0uZoUuP7uUMSo6aLKbZG+VwbCRGjX
IFM4aNRRyooYiUI5AZdpjXZVwegQBOemAUiYRTMf2VBKloSapLd1erWPdlW5
tkpsgvktFAXESTlrNV6U5Em/kk5u0a0J7VJFO8pgWS+vLz5BGm+Fq/UJPaTU
mtjiz1dTOIekSKKSqVMsmcB6fAyx3L7jfCdU5+biZf7tx2w7glRdHGxVKmKD
ybwOJzs+zJVMHcnfvuwzwDNshecvSk5qSNtN6gtBOA04MqUYtFrfB3ltNSQJ
OgBidJZZWq5SIljVL1cxW9OdgRcDCcxmJw1p/H77NVBOXooa+pp9GcgDAtrh
6DfbO/Hi4frViKtFPR+uQ2A9psqHpslEplXQRDDiqOhlDVy6k17iNc25OOZ2
bWWUbrjms7qSsEH3T5BmumDvxShOU8OfSXrLjrxMxfYwM02uN/TZ7sA4ZqQ1
w6PF/qPXeZlEm0gKMnFt9w+occqzk6U7iIXwoBDl1iJlNkmh43OGN8q2YAln
tLHzn91M6MXMgZucM6j3VKWH+38t+L3a1CKnnwJtzOiQFYEkwKwHPFoHBHj5
XCYiLfylp+b8RiI72Vvpt3UAvG1q7rR6zZqy8UozO56z/tVyyiM2OUw0gWKb
Kil4UH2OI9WbYhaqt4Mbn7O2oDD30hdScf4n+uON6264qk3OZR7CyJEep7zn
2G0vRQ28p1bfdhDryKvPnt7GLfnEK26GAwpMDz1FT4aoK28A7vGOC+m4uKEv
HcVx3J+sK5IC0Oedbut9EcDxqOnUvVrYV5roi5Lqavnv6ogDSKcen7c+9QC9
9fEuGSP74sGsYWvKNQ8jWPnQ5tGe9OoFMjiHLW2f12I0dP9J9NxQrIyw+dep
bHzzJ1VGymZXSPfrBLq0iTKLFv9gl3wVo+KxMuLKEZTSm/Uu+qGTKpYLdpP8
mHPHM3hr57q2A6x5AteGYVzKT+9KT/6JQ99w0EReS0MRGNAIz2hy6BZv/r0C
5XsxMyl8bPyWhRmFNeu7FjMbhRVb2U3jriMb9cDDyb+yDPkmaOA8CccfYAG/
lXR6+04CUgvRnhbBC8NO5q/1Ypu1wr/nBuQhPWmx5M7jkriBDT3Dh6NlD1/G
iSWME6GZl/B2Ezf5utj9FC+gamvW/UCrQ3pWad6zN58NE8A9gxLsrQYgYKvP
251BhutIfl9iDRyvhSGZDrlhXiLx6yvr5IpX/xDZY8+aPoK0Y2r6JAGwMNiV
NaJKXWr5WjCrzAJ3McxtDHQauBiFj+YJgD/m7wiNX8p0t875GzaxD42hr800
MWAfCt8jVlG297KdD6RVg8P4AhwHiiCMtkUp1y1R7pQuTuMmBdXPXq+X87Jy
n41cURtzlsHlHarZ/lVSmw9xOphdE+88LATp8lw4RZ7RgL0dR2lMtx2VgP4y
bVqXbiDIMT3OBCaCEJ7nAAwbc2KsbU1FBuHgSuLZ6600cLiNEoDJL7hzSi0a
nf47sf7IrMMQwOU3TXR81SzGiMJnzCnXLkiKzODO899jMgJNMBU2Ro2gJjyM
4877yYEU3FtCfMhIhP2Ovd5M/hD+j46bVo3cks5Wg1fFkmRziz7NKlAC/1NM
iv8ZZPMRqIZmbbM3TM1clNODmDf4vqoKz0uqpPncZVZJ5jPpF1IhS7f0bgPG
SPaiotgYSB1PNSB/DJy1VKD/CieJ3M6P/qA5ALuLJb68ka/zg5M54nnsiq7s
Dm5yaGJVls9gSTWWxl9MIz/rRvyHUTSlGJdbWmIcUB3ncECZzb1is+9DdNcb
DTlIsejwKxevbvizCKatqtiAa5CmJweaxZtloecf3ifkD4Q1RGMDsj4+I/7z
evVLcL5eH+f4rZ+LQqHZ60f8n3oIpxbwa18zzxlSnV1bmvYxrXYIacRdHLaE
dDiRP1D12JNryXDxk+oD0lbNwmHZNAyGPWrSsWZ5zsHeHLzJgSEJ07Aemm3w
ImOFFWhjESZkp/58OqB83bFQLEKiqYZDx7uLahnc//DBjDC9ZUfSzoMmNaj9
+h2ubfgswS09cpz975mLAYUMp2vaj1uFWCrKLWwtKd2H+U5xig2/ZgvQfWOc
OCfcL846w8IsvYkqEpLaBGmVP7RtmgGmb81ZGUtO3aUYmLWwiAQcIOsXWp/o
VtnRBBvGd6HC8U3lef5+S2fAlh5cbP7FW9/cvMVvD7EjpV1IMdS/WtSqWAYm
vv5ojnqeB9FlQbLj9U6qrOTiExLi3BYQMCBA41lPyXhJ+lt2FUxkXo73felz
oHP7Ephawp4JHUArImU0JL4DhXwex1Lw2K1gmbozLPhkDIu20FF4CeFV8Ca4
fcspHDvEeJWKSWd7ooy9fQQLe9h2p4lIcB4TZw/SrWreO2F0NzTk+QUV5y72
63vWV03DFkMKFOwv0Q3DRfwJ+gK6dNb/NcYqFgvJqS4qbTF3D7NLhcpQD7B5
Qr9aEzTNvCZFVtZI8jfQzLy6NqWn9EeG74nXP2MMzJipOibhsFxvZsdGR+/x
Wgv+cY0ZGwS2WkuyvcU7Vs2p7otVmDYDAicwihdWzDWUnO/H0uWyIxDI6P7S
dUlGl/K1rllKEJph/0SbH5HwOFdJIFqOhyrF6afHjPWWs+Jxpox94JP2qbyk
Q4q3dN/HTPhv0qHTGqXlAvFoh+kL26tUzt6GU0j44zwajJwi/BRZf+ugsnCg
uejRPYZFhdtGFV7KWkYAf+X2y42KPlw6WtDdj3cUwtHyeMEip2tUy9nDvaEX
MRaWjlPlx4bkGfNxUR0XxT9pY3M4DnFC+dkU5izwdm7WpzKZI5VxEW2mCSVv
S/wznCu1dApwGeiFmjufwpCBc0SM/OKRp0A0COZ78Y4i6iPugnd7izmHNWUu
DuBWf/NVSqj7W00lWgTNP4+7h2ErTDbXlG8WHxl7/8VO0MmQ0fyCV+Gpi9QB
MOuzWFTq6r1ffu9mEO8yFNObookcjCQAoppf4qJi/iATdx/8+X0+6iJ3GGox
MH1xBi4p28EDn1ccuiY5Y3+lOt9UOLD7YI9z2PLk9VG1RtE7AWdnpEIYVGsZ
HHfum+kY2sI055SD/43eRk0CeCSh6V7KhMnE9YCtGgvD137GFpM5zuMdk8B3
EcUiCvg4aXKk5LPvbDSqTq34dGwTTDeJ/CjgD7ICRQujaIa1/WPvw0InspPb
h/h2v1lGZgt3weYlW/+iYtgHDIuDvcg1BhRu5eimEMMwXrw5JOvr0E55H7CC
kGvsCdEFk/oefpt9XN/DBTECBjSIYoEl96yMzxxjT2IVM7gwp/zkfJfRucLz
CRbeG8wffSebDSwhPE2FlXATpL/4SM5AT+BkKq/SdOVN0mVKzsCS0yndTCKD
AzXi+1TC0mOkDk0e82kcBTe/AngLuJ6Om8soBqq5W0/43UBdRjmkEQnA7kB3
TKnlos029pXRqsbUlWRLRmMBs+rMD7hcvLbWdKYIvTPHEQ2J6v809Pnyt5K6
j1xWigEGKP/GV/o7q6CDAIk17XzYUcBu73F+Yq8IBVsyiw5xUjLPGleK1mJ0
UahUwl2krorObTYQYAX8Nch6igphX5PPldcvAnaIfZgWYTK88K+AtXwi7QDr
8LVoHK3Wb5cxu+3TmjUMHtQZ3VEnMHEjvzlf9yy6Sis6ss8kU2NIXH2DS2d9
FhSp+uQfAt2KbEB3UwhoYkPByTPsk10vZNHq7PdBzS0JNbcMhQEA2/FPGy6q
gZx0ZxPFTY5Is0VA3CMq+ug90hQL8T/AJ+pdjolDyk+QgrTli3sBiMtfPx/p
a4PVQXtJkHxZzLzeP0OD4ebostn/LoxkvHkmg2HNvicGFle2vqP4PBfLqSrP
O1H1SzK7Oi6gc15h+pBxmNh4oZ1qra7SvbcIrwxT0PXm/U+GOcSuTFPMAbOY
50b2HL0gI0zokPg88a9P060Yi7K8FW+bckonjkxVM3xAV7sxYWCqOaqvgg5C
fLd91oWaPmyws7oN64azsMuLqh2w6gitCRmvwgo8+U65Ab6LaVgrCeSwAyS8
7mgyzCT39vuuPipVNXoQSxynq3jfp7p7L8RnXtGrXs7/6gSQ0kaKpNMTaJM3
hzLEK1e/JzfDxKuhto49b20hVFRubOYhTniSr/M48ScF4FXUVaUAaCcLRg3W
YfZtJpot6iwkrxEWrOYtEnn/Y0b2R9H13aY0SvaLVAxOvMpFk97S/XPFdQdX
TOguvICWRtodL9tpLbPo4+awm89mquU8Kop1AXV+02KUHhlMkNpGVZNZS1Si
u3O9Q+NPrc85Ntxqr3yDxEcUIMxOo/scV1sHZqvcnG2HAI42jve7cBrqiYTh
xUgDAQvITdN39pbnDd/4jIovNxVeWFZe0rtRuCK4Zlnld/g0KTAaaCmpCUt8
c4nxMmM47bmdS9hfXI9LxfGZ1v/QnJ4/HUcYUJNNl28MxZqvRXjEmSvy30dU
A6jwczTnkHUzVAN2PzRqhtSI8J/pQ1i5q07XKjiIYNyDIINGND2uJhuZgpBU
WxMLhuCdh2hkMj+7qeR+crkTIvfUBAGrj7wjeR4lLZ9TpnfeiVg+AYsGS+K8
Dk9muER3rcjfEN97CNPW5HQLzDbpxmwCSGBErasx327vBud9QeuHrK7OQ7eU
5hcLcwLl7flgRmp437YgmfMFu/krdcMf5jDe75LCU4lX/KA4QJNk6L1InPkm
UKIJeRpSUhBG0SOSowE1Y/omLJdXF7weVCuDP524eAL6FhhMeOwTV5axcObq
3Jm/L6i7Bumf3iMGZxk5S5ZFiFuR+x+0inBFXisAwwl3ztCEUA06EAkP1abV
JNTKqjUDO8gYeKgOamb7KYIWV6jRXqR2KDL4lNJhhNXVqJRXIX0w9UKFwxlp
8PeuaW6OUQ6rjS+Qs/WRVDUg9t1FoJZqoCqCAXeHu7jrvdN/IT0OvIbagxFO
7cn1PWLoWC4iV2Xx2F/L8WPrH8LJrwQ27gJdgY9xwfbldeu6JfL51ipnVPiL
WOuwm8cHbFpoILmPD33VEbkArn7bfyY/2w4mzlCzBbkIfoUxNZM7gqGphDSm
NsNop9GKR+fOuDwOKR8zxXA+5CtuEy0aXJDlzw2a1J1CXV7xpX9MehlUe6U8
FbdCYT4eJtruW4aafKjqJ2fS+IKlmnopk4fxY1+0mhjIahRWI9P7E3pICZWD
1GJRKZD/sFGzI09+keH5nJw51tlpLdLymo9NrJxzrNyN0aGQVYYYHe3M/0F4
y9jE9GI0g/oNOCcNO3nhmq7mxcLW//JqgQb+T9GlkQsxvXzVHxbB0qL1n2bD
6f2Se2nlqF9f9lH7/P4N9ZVAscDF61e/6DtOd2wGEYQ10aqUUY+AIPId4bFQ
ZPoQoldBzK0nhhG/ypKSjF/332VPs087G/jhY+BrtiMYovwGStupwUWTxLyz
BVzgZxZ88Lup1PNzYdlbxBkCqw+v3jYaria2VL3+5I/NWLHMN2bEgOWXqxlV
oNXCc5KJQ7CPumvZDhp3I9sIVXwui4eKaJ9kRJXtwKivyn7wYAFdtgrUdSWa
KMiX0WHT85C5ZoZAsyrmn5qVvCL6TqoBzg2X/5v857/8Rzrqe7sFe7vdabWE
on0C9r2h4pAfukEBVkgasDALJ8GqeKZU5gqrb/wSNCbHxKrbgWYJAd6okbL7
FhTODZepys8G2vrHMdiy8QXus3nsFCbxskrXpuyX2bPHm85OIdWgebOjBme/
9m4ugpUq98uoO3VP7k21o654XXD3J/7BcEaKO5nEMs8hZ+R/y71hKgsugszM
jYxHWwIKqk82Xu6Iehqc6jmNTMqrAHP088wS6Zoh79RHVdLPH8ChVRclS9ww
DXnudurMScwH3u5/ljJa/77a5LX3aofJ5FmDBkveReqLt+dgynqTj7wI50qB
f4snc2JRaaSXzKXSuRrDBXsuTSM4RThbQbWWYApJ7CASyGweMaLVWM/f/6m0
ca+36bndtFHC5i9xMGwFt42awfNlZnfwOcQ0CYTz7CPzGVxv453g9z8vOco7
zKINfaSJYkAIjVSmznmEdm3yJiZ+HDATlzr444HLcRS7dhbfIJGin+ZvzWf7
3etPKQbRfca3tkzLXZS1BIogBgpBhyWCB6cfIn1h+W1e7U1D+iL6UGpqb9jy
NUp3IKPhfVrZHay+NywLmhp8izG/4xQ4xVU79lnB0KX2B1RYbe6FEyDOOm6Y
k6giIjj6cZMXbaP7Z6UB1NVGKX1kgDl7aMAth7dd2YWdIsaBbkN7cqj8iW3c
YqbXrnNJdHOx1oOOhbPMFKfyW7UDF2QDq3h1CR+bwvUoCsVrrZyUG4dwHizO
5ouqjcGO8nYtvnZygIA5bJDDjTodH5ev15JvntAL+esUDXJr/i7FIwv6ul0R
QDK5SxuUInc1KVQP8iTSUTB8YDh0wzlCf7yTajINUbcIXFMP0z2yOinqEqrt
HzFgXu7WQPZ9T2XInDNN3BKxb4CPowvB6hU9L3laSWDlVuRzGCds/XfHFkBe
VopaY5iO2TZAK2B3OZqi/dEQpOTzEb+/0zIrlKuEjb8cvxIO2BDN/GLybDXg
e1RGMm/CY336DI0SVaz/EKCiiXIwGmDdeJCt2qShgzTtnaoXlauFFdrYlnQC
JmeakhSP2FdvIOqAotWKFcowvVW1QnmaMQsEsy+7joDjOGDGlsdcsua2aOAs
xlXrs1kOHd6uPpig8DYxpscoY3hXyxQjnyXxlQUnBDUM5G4APzgXC7v4Hj62
O0v0MfI/SFoJBsp6dCIGozx9/TuptB7BmK2gWV/UvaijaJkPB1X1xhnBPxob
invrNGPjMV006Ga4DaXguatcje272uzW1+pMPUMEYb14i4EHQkGXR3AEjo/2
SEpOMR0cJsVaXDr2wNoF2UOmV4a4XPUglF8G0hmhiScuWrM9Vm1q4d0Eu+gv
aMZ+SWcO2tLEerxBE9a90OxZ+7LizAq0asHKvzhOAEKI8iUfZru5tENK6HY8
PVnAE0dP7oJu2n7T+55IZauJl20lz981UGaBW5LC9hP/08qsrFUKlu2x3MF3
6mhnjYHUmbyIGWriRwh+lk/KLaD/YVl82Q2SRnG/LoKOVRdXEwAjbBO0iqWN
8H0SnBoNGZ+dldit0INxBcH5P/G4a2Bh5P4b51WRJphVAZsRoLR2AYyo+ovH
9qnmTHfy19Y0LenQp3METd1MuqWleOJEX2Snp4P1MGut0uI1LO6DVNNzQWKL
UmLl6ky3kJkI7ObBnBQzcwdOOxdINgmiarsHebypWnPDndWp3DNKNEGHtm8X
q/4xY4gFggDNV0Y6PGh2zn/L4+bsgyJ6xjVRfVcCSqT/vqYQtDibqtoSl4EH
DlGzQ/fYqxHJa2pBd4aaqKZG9VBlUd7+dRr2pjkmITy+PJDSy1jDERVt0+gk
l8a0BxofunSxuglM/i3xLVL51Wni1riwvjSWb1uOMXIdKuCr7t2nGU0mpC0I
jpb09b32b5ScUdN2iHQQmvYycfQBbZRyeeDQwIxYTZ6lSl1FMdgRuImMSbsa
4Mj9jMXHsJZJD0noMqY0oM+86K+j6FcfrbBTaROW5H3DiIoDagCRMY8tXh6w
4wx+DymoQEJId6cHcTLXnuRhaTldHjf3ukD0wg88Opx4cyjBJb8SFjiARBk5
9Kykp74ffsdMxh1HwbQXyvCSTPWwrzHZxeGQJqY7DbWa5aj8G19nQDkaMsak
gw4gPWwU8RnkbpkkxRUuvdCEIJOEpykddJUpwJnn3uc5nWo0V5RjlHBBLef4
zNC9IGu61aA9B2VQ2cx9jgruwg+2QM2Qp4xaWkF3QXR/Zi3EraXGd+S6Qrp7
u7pEs3EFh3zGdESRmxYDqyADYLUFHCztJrUK/A3JOAyDQUIsYw5nmd1C2Da8
vbU3c3w99elXQf7LlpupLrZlCaOotU2R/mj/WQXQdcb+UwWvUqlZ9lseXFFq
lMBVSFf4xGI2RJrbziM8vhYmgXkHOws8JrbF0qdoRDOdBAWze+TvwdR1T+hz
G3nG+XjzAG0YiSH9Ti04a+kZUiQDnz4e33ZeW03VjjEjyZfTIobktnjB5vj0
xTo2X5raWOs8gn6iFcMpSeRT5tKA2rNku+Gsj7UHG9Hm7g0iS55rabL74n20
8Bm8fzEyJzmIrFhc3szrOpL236bwGu0n+Oup5YVxkLYkX/htatUGm/WFJ4mD
MQjURl5N74DM+JphYtNUd3zZPTt4ybcJT0dApOyztF3ZsLqVL8aN4eyXExfr
bZZfveZYRwsB9xcCgMg3zE/G29wHYHcnqEaEjMDMyWGiolWUcAXl0z2uEXH0
TYHn1Njc/DiSz0L1lo/6394HvizActwV2hagqQjnbv/vam49HCpAM4zMDz/x
zamcqzbU0fVxv9rXgMTwYGBHRFSMF59QL2XQ0cy7TXPrpVgEgzTaINgzASg9
tdct/BPdNU7VT7im+GLVetOz/bbXYPchjEDYrBq2QY0ihoKvD3XsF2M3O7gj
XTXf6kdMvmNqPnBSXmGgUe3w9PUPBNMjqOILWFtIHxJ2ETLBpq8HLrqhffOS
JK3krzwSFp0vkyWBatjW3nVLf6A8lbogIIOIZNNjxGLVd6Y9euWt+QEm+2qS
LfNxDqC4bNmQcmDf+VQOGOeIXl9ugXTGB8y6gm8xNZdQhk54mADB2BYlaGlo
fi//4Qf9kICY/0uJntYAM5XyPo2gjvHLzAKGyxxSvnuKG6/1gs+6spYazQoz
dYt4Qxc0LUgByIXHVu/cxX8c53o67KA/xo4qji5D2sM1FaurOrq136wr289P
eHvTrX058Ra3Qcp0UXpIZiu/wwJ3pSCo5TlzZ0hhx+uVe4cEVzEmYmoAejow
dllj/VMN9+nGWzSbhNCkdLnq55vZ8StkFEDdLGw5cWml7RrHrhsYS1DDHHeS
PIzDJge7VBLF308hofdmAOtFc8FtJNTtqAv2mgMEhbKIcZcHPM1AqXBqmGhn
rCiSXbU1upJ6jVPHmwnNNMCvAVu2ycCTm9KACyO6UhlPQVQmVD554M+JklPM
cB/M/tYem43IXRfG8OrOlbp/RvRVjV/SyeFpEh/TEr7CFPyt8PizE1hGD1fq
tK5P/lwvglBvsoKG9BxmaMlVOJKKLM47ReeZdUxXlzvDwu6p4uED3qVINWch
/HBg7BlSQPNzcwocB4S91qyy6Az4fJMitsvx4U6B4/dFUBLit3NYJ5U57fh/
LtETFVx7UVXD1popJDiiglKwj/EMR/rFzZdfQ0IWwntN+f3el7gCXx4WwOym
F3ArqPUlk6thMNpJkYrKSxEcurZsxrkhH6/ON6Cr4mnf69Gpc84nCGrwvRmT
BqPjNrrgIjidzM39T9vJ1Q3U/sUE76Dvy+ZyvyOEDHAzhzvJG6ebvnX6YaNT
J52CAaCEvbbBmibOveUxBcQe5tJA54FnjusNUy0ugf1fBC9KOBN6F7xWvVMg
Err4fzcZGZD9iuxsJVCZe0hurQEZbvJj0IEim75wCFCSASesKCu3LrYQkLsR
sA0cnQl3W21SmsvN47BXISIusipFAlLB8u4WzUYVFcEp/gZmzSQWTrck/BBL
+SYuGVxT6zFDrUL5Vas2LLCuJgGyKnD7FvioyMyEUwryaG/5uUJXZPUjgNRa
oegiKdPY1fC8veZYzC9z1nxjKZIwGh2SQ8QornTEHRT4CNdxxiycfZczQ5dT
ZZ1cVqS7g6dzAlskkobcjptdUglx2VQpGPFxxphUGqUsvdJKNyE8l9FIdBmG
9dmEA12lXtOhZxyo0wn4NBsQHMJ3xcGqWqbMaAuHgJbv/4FWbXyuHYKoOYRD
E1L2cMn9mbMTrjSLR+WflSWbId2OislLjuD5W3P8/cMKzRnhlj2Bqm45uEqP
DmhmpGymez/BpX3kCZaFBYZjfI9vapMHe0rwuLEIAzhL8kkgc5kqpOxMkCRS
jioUXaSmFXwH3vl6I65g3mkKXzZkRi4DZY4Cc3AnNYPxBssHQ4ujLE8kSM0e
GOWq866Kd6E5OanYBd0CC3GT0d2fziAMNZTLtZBAf4Rzh8Xd21KItpKsfk/2
zktR42KyJ9QCAdaiqcCi3idhFdPr7O+AzMM50iojrtW1/SIfvgGAyShQIt65
3pKxds43I/QGOGgCJC4IAzgrTJQ24Y6UibUOHilnPbQZBxQmhYXFcxEmyifp
iHnsXezvgmceiiKeMC3g/abCgNUUnFJloF735pNoTK5Vjo6YhGUHx/nZna5C
Y2sMZHLOoboz84KGt9DjatxSDEftRGGUkz2ukVC2ygGq2EIv9LP0rr5u85Zx
TUzIItF5C8L9uDcUzXVaj/axu6JwBSStU76CE+HD5uKFhnrnukfdfvm11k4W
9ZNhQoHOMcI1TM+0E9jS7Eff8aqEuubOigQ/BQ22l90+BckNlzGjf3SWR4T7
RSwEA/v46w1D6XrwBl4DJnJSB30fuLhmvridAgye/8feRbgXMiZZ2j59LShW
numTO/WwnnsYhMmbwSFG3O0dkLqe9JxVcyAnK3zCMXGxM0hkAtZ17E0JnQ6o
gMEXYnKy3+tGCzZiBr2wopSJgI644LFz3KRDxPLTE/90yXgkcx2j/wkK4l31
WAxea9OZCuZ1fhQlTn10cvp2Vk+Z1N0VNM2jZQcJQa9LPIm02cd+T+sxOrP2
+fH/RG3AQkFc3KyXUY/1NkfeDhl9e5i5RbCiQ7ehVvL9RwOGMNF7Wr8Du4F1
a/KQBpApEI0gg4LAzbCJFGJMVGHnoJHz6hAHpLuq9Cmal000YkD2XnzIuj2A
y0qQ3Sap61uVSV4U24pT2rpsDOm9KyaLfKVl8PGRElGz95h8cSbw+mE5h+tE
8b9k4lX9QCfBawBPrGBE5SgQXf8zVHkzIe8ln6V+hqOeRjs/RFRIx2i2ve4v
HyYKKIRoO+aiVwRrNrNr+sZtnD/Ci2oVH6QUzOZbm3sx7iVidpiujPgH05lQ
gYZG0aKUV/hEZqw180wfL8jgtyXXl3hTq2MwNJJjziIwPc9v8FR1ilBmtBRD
/N/Q3vXeH+YXUnifUGZal4EfAqCVd7sz5t1A3CNaUTaG/nJc257YovcZx0K4
a67CIG4/Ot4r/cu2dEsKlKZ1RAGufKMUez79E8jL2rEVaNWgYwi/6+8+P4LX
Tq7zhWnsQkqUa0JeXxkh/X+Ft1/7uLri+82HkZPcWFYsQN4w5xye7AWJeJ0W
J9/UpG7c3L4IuHq8DPKLLRkfv+4MTHEZJ0aiHzbD5myPPVpCK6+5fr2gK0UA
svu6O81rB8z66kDbU0bZZxWzqRAt7MHjTjC3xOCGhQi/KNFz93/u+B78gunS
bUGRdeHIilsrBqzhjnxWbCjA6GHNfEt6zhlzPChEWHqSD+qNXrSDYGLcnyb7
NzGiRWol/+GmSJYW7BTfJ1eK0w5g5jNTin4ZpxnifrxOc6XU9fwEf0oR213Z
B3gsWJly6VBc8N9XtADkhKGZx/5qXd5jBi6kAJAQvYo8r+KzT6NFlrWAvQAV
zoWIYSvpy9iB0KhZJXKS0yau7h41XOb28eRQqZPuk1+eaUJVbxN9dKqtpYVk
tPxRzduvZErvHUDgQmxdzKJ5IHvLLw1yrR66YQH1OZX7Srmm/ZwrHNvQL5FC
IMcHfOO8PagePgcWtieV0qXNul6tdUj6Jy03RgPOvVW/+HcNdhfEXw+dClv+
wYt68ADXlbdx1UReOU53Nfg6ACYflL491W0m7NZ2bF7gXdiYmqtd2XpCSRa2
aySAcICoBmG2frSVluBevcFXmh7p23a4JAKYOwgINL+BSC/EIQFXeWps5Gke
RYi1TBo3J4k+mle5ss4jLRtPXxMmmtROdXTBHZ55g8CRskTE4u1ZhaI6UXjP
o45xHnUBpYmiZ41Ub9db6X9kRAG0KGM8758naVKLT+naJdEqwaOUb4z638EF
1PnZLqMzyOi+oE/CIfCtmi3PGykAFpPM43aQ94Nwg77GL2H5f//axAIYPNVk
Ara6uE0DNgyXbg2MpFaSwlRI0O7qx9I9apw+lZSWXqXbzNOkug5J6CMqW5gT
c97tq7yand+/5yLpsECnuhlvKN6pwD9H0sOHY8sfkWfeEsHGECItP2y4RBic
wMkoQp8Cn6UeIfiWoi6fP8/gie5tw7Rg4ORtParqOgZbhicpRquiGFKPNeJy
PiiFYlokXYfiPRVcteWGHukOgWBJg10+tIYhMFVCL6YgvJHDWXxBImpyNf/B
1ODurIwzR3e9s0tzp2llKn+zdu3HazJvJrRfqtbwqNdWE5JA7nAAJpVGt6N0
kn8rzyaQfh4PEoGKBarfEVbqbZR7q+R0JQM0aoS73ApQFfWmOxlxDRTBclC2
l2vmXtGflk2e5tlgByt/yre9pu9SNOXPWeQ8JOYXiMBAhKrA/OK/SrEbjKcw
4h9+EoqinFdV9FQahOrO6OFkA6ZWRVh8PWlxben8KBZ0oUXhtTg8X6HSofqE
TP5E+h8DNjUXFCgdBhqqndB91nmuYa/Gbw38ltrCfq/zX1fI7//Y3bXxKxRv
bjBxoehr22HVjMQk/5ohKQNW89DGSZtSISpONiNhPLyyM22JE+YxEvNQihnW
g+FZKYYe7736NnPPMnHKVZ/R23l1hflkYkZDusRx+QjonfSu2hyOSEC9VjoZ
F0yiioPKOfcPtjjAFN3OzICjkYeAQ6cy25QxLHsuc9rqmXOSJoKSGkh5oFst
aU8itjTXlFizYY742cc4YEaq2vkn7IrhRA/ZLAUrfbjiuBRlzDW0JOOlnOPT
tkghMYAi10r9SmPDx7z5i64Fa8K4BwNVI7vNyQRKh5cIjbdxWspOV7sr8EUm
TAlMvK00eBko3k3vDl1R7QdpxawUUDzR58gyWSRIvFrqHAycOMYXFmwFUW6R
D3LqRmpRmiKV/uXDxqkafN0JIxcD2RY+ZRFIDVVH7IuYLHb/Xr7kUxPKulMn
TyYaxhoew4ujChAW8Jr5I/SJG2XiVgWL9+MNCOIvHooGjbld9aVxyxEHe5l/
/nTpMIbxVe5hRGvKSGrGL6PczfHchhgw6s9bhKHIYNbF1W7IfpgA+k3fLL/n
r425beqlmhlSZn9gARotGFl8iRUo5QaDP4V9PyU1dtS2ENrFJxEm7h9p9iuy
1FvOVbtkcGn+1d1Ozv6K9m4K+QpqBt0jbfCqcwuTWPW7d97FGfc3RZsKiJUi
hwy1LV5CLl+dZSKBIcf0PvpHGt/q51F6QFeKfWaZThtG3ONOjwP8IRZ5meez
uGohXsPFvBXs+7a5iEzFGKoNpsADkhHUSb/oOcLnhCkv6bzOIrBpTO78WyUS
ccZEAODB6PD2F8HgK9DLmKrfUc7OWr5NarrAy0lzyN7mEmb+PgkW6o1FhB0s
pLxIYkbM+STDk4/vpXf1eCgzQiRzz9uehGxnrieSyRAS4zGBiFX3Clu8GVg6
Npa/4Otofp0eirOun+pSBPjy7ITVXnDSCsViBAi5XoZ3p8LRRDMoqXzGKMGf
mJm6T8fHinob9UBfMIBa33W9L+uqY+0W322iSM0wzukEkFIBdMhvMf/TU6sn
xV5JGOANIkX1JwkyZ5c6eGtalJ6RFbV/F1nsSEhsALz+wNbkRBrSMpsAJ/oK
Iwn2nlkno+pt0RyxXA3vGyuaQvVSA58hNWfKe0QA1yd4TJR9vf4e9H+6s9cI
xEnBsevqOoWhMfWOrJ8nm8JIyeGZcAou26YxbZdSW7TyJyy2swaQHT1mgyVw
EPm+1QBv3oodzD4M2Jn1E8bktdiZrjOm5gPHcctWQ1Y1AnsoZ99WCjOGhJ9s
8HzsUjOvTvf5a3kRxy6YE1Vf+p6uRuk6UcBthtUmwwBJ0ZpVj9tWRwPThg6h
p1ssxW/Y3k8IjqSiRbi4AlJscsPZ3P2A2W/xSD8xWI4SrmwHhQn2B74aJm+m
tLTXgwqENtvzvUB0rqo7pfj+s2curjarTwwky3EiMzySko9slnHSSBf/dN3w
cXCgFk4zkFNOotl4wuD7JhHZ1mz1mwb6qHaV8O4vVsAdLMJIjCs/AzF+/48d
8NygbarF8ChybFTX7FGt2VRagWM2B34m9WgQ2OycMpJZGWgNzcp0hFye4FXX
yRnsmGGwwcJh9Py0Zb2hkmz4aXJyXk4FE9M2qAMOnefM44yAVXH+BOl925SA
qLGmsfFpo2n72214/e7iWVcv38FfF8epSbbJRVsJ479Jb7J+l1E5hk/rr9eJ
t0eZLqUiE2kBE8UwKRZVgnxQzLDymCTm8tIo15b08aENeQs2gMp063T9jyGc
pYEpvhQTd7TM1+P2RDs8MY8c0MIP+sapdg+pHNdqiWBvkRJfz2/nNRK3uKYW
a42d3YJUWAyYl3mwzrfB1o37+0hnV+6qIrLkMeyhBd7832bhW3SfBcxk1UeU
Wi5nazAClwAXP37nKBQNZJds5hJA+/fv6zVpCRihBXvI/cloB5vEYcthH3Vt
WCOEuaHXY+QmqflQMmI8igOieg8IsUvGIprmEy0oYjwQVLFg2vDFqO+fL1UW
testTNRrk60A7RAOOCjsTbGSGlY6ap27DBPF4CRXdvs5D8eXchQiJfHNS72c
sg75Q74Qbaw3q/I4UiaZtORm3I4c4HtBF05hAq5q+SakcFgOCiAcNjcYwkxu
qNXwg/xhWyRZ4+xF868qxva+PwmUJFfbgFyad1DSl0yfmrlvTmy67DCC3JE/
7yMw6QQIjgnxJ8FoaStx9ece8S2JNfJf0mJR5hMotZKh/kOOH8xxsxERZVhF
gPOZlPKR+ViN/1MYIur0NIuaRK/F7h2nzUVaKhouTIm+Hb/4Rit1/QKlA4YB
iTKre2FwMpP2WJoDWMshE6AVu4dB8N2QQ8MsZGHN0LR9KVadxGMYeCn7UjyV
e2T/ZWNCuI8J9SZmv+fro7xpuuYpwPhagJFTD4dhOJn2XLh5kY44hBqcgURX
/CSUKyipAT9IP/0ZQWM8TFtUEwDL7cv3jFyAi5H6J9ObKm53RiHFZ7eDT6Eh
INrSXRPxA0LXoXoaPcK7LuWO1w4cUqPNDwYv8R0M4XMelUEX4Gy814MXAkzG
bDuVBB7IgHsBA1YfwOrfG6sCsJaCLhzkKnee4ZkrCcY0xc3PlZgzAN0ts+no
vMmj5i2/62aPD4Q0M4LWjWTynw0+W04Z0I4fKFfx1RCHmdVElqiowAQq6lSq
46Bzfbv5oqOd/1rh9J5ChT/xCxXy4ZjqwS9tX+uQuXA5Tq7J7yz5HceJjjKi
shMOSoBWeYjadD1xxx5H5J0M53YmZ41KnAn9Cwrr/gFAhshhInPB6+7eN1lx
akr5YV88UIG3jcpI4iGToeS/KLYDnVfidChR6Uvb1d8iaktrEz691mu8gFIz
oOzOZgwI8hrPhXRVplFTAFV0Y7mv+WAJEHCPjNrfzi87ZRUwvbZzTTCsX2wB
TuqGA9SxA3c02N2BSOMNXijRGwc9nzOUlHiKd/2X7NHRf1qEGq0YRgJWF662
C8jUooEcc4JtEaw9JdUqR/BJeqNvdEYMTdIgLv26WFsFZ//AiB4owCNQ2U4r
tVb8+ar/Arx2v4IAmtWShGvOIX6SGAC0u7+AzDrvAR6dmouZxVFc83oRkEsB
gNwBz7gbLJ9051jn7pie2CQzBmHT2lab7Fn80FmDW/Ysv9dLdUZI2tWSxWOX
rO4oPYUWTNICpq5eQjLrfsZf259u1kS5Pwy4IwXSSDU75C+YHda4ZrDLQPeZ
eU8LfN1qa8TS+rpdzLDDI2tF9EX3orsRH3gkd4+OnX5IiFtTcSuESngc96cv
s1p/MBQmH2dkmIT6UcTHVol/dt47hrzgIJEPo03Lr2j6KeIvRCowFRNuceIp
yOvD5vwxjhrJmujnn2n3BI7TIzOviLAvsosyzPhxbfcXkNoTQP+gNg9UrOO3
iWsjYf36McTw+YQVG+2j+qd75xckyAiYsmBN8jVNZfvXrdJkRy+At6hZi4Mj
Y9iNMhP6RWkwz4LKjRSq7FLcN34htM7albjfa+N64ieiWcYE7aRTIOTglDZu
MCX6KLTEzYY/U2GJqup/bGCts1H/4zMzQmNpJBlnd8d4LW2u2bc0U6Hqhfwi
cv9GPGoyutnNAsQD1sv3tP+FdzpMBGGK9/MKB/Hg0HSB0rtrC9emUqJtf3jM
oGcgaGMzToQmHnAUv3EUAR6SEr7PizJrbznzOGsfJ4kNN/YJ77pdNvUbDoWa
qL6xbY0QMo9EsPzKuNdOHc1V7QQO/iu6Kx6zEKVINsjWnCCH4pUQaa2jnaSF
+mXwKQiihpD3nIaZcTDBdiRrJ1V9GDa+KbQiEKoyylD4ofegDj0ZYIVoNNFm
ZsjWCHhROJblC80t+p6qSHRmBqXXnu7g1CTm5ew8Xc8CxYIWqvZowhMD6tLf
8qA+nC9MGDBfW+i5Ab7BPLor7QdM1QbaHe5LTyPfiqffF1DjsR3R2Gi/mebF
37uyExElULy3y3GIVEQIuE6Da6stpqjHCPxL6s7jLldBn0/i7b9qbKs8fo3N
ENLRIT832clITYyloiGZAaZtlC71rUmqduLUpvOua2eMboEo8sPp35z6H+0T
vxYOGVaQmWXAxQEEm2chmAL4HVeDADaUJBbhoDtZ2jG+GUtAV3HNgbt0WMjy
j0oyi+eh4Th5lnLDbb676jVsqtheGU1+MLW2wHfZKxqem7BJkZWTV/B/VycF
LhdcJMoSscBpJSzbsR20+pqTgjcr6QlBtLVICURUw2hw/HAOju/M/jUvY+/p
PvTdsV8EHDQGbfMAIKOaaTHTh+mpchd3a4fwbVyRO56qHNfwlisPRYkkZHUl
/TA4ksvZgMGqAIniO9es6uHT+xzhOmY1V0A4Z0tB05+OhKH6XhAJ9CvVggcC
n5sY7/rxaAmVF+E08+OVfAvj2bkMM1pMqvyojmznDIDhYkL9CqysAwZ/l/EC
ieymCLYflMYp2CaGEB32h9CBLCBYoMPaVn3Z/EeicsexkEn3pWId3ur7zpJy
DclxjfunJl+bThkpYZGDewzm4izKQnQkzui9nBi/HKp/7ARsodRR/8BVyFdo
OrX+haJmfJuSxih4noJ3rqXazQihSs0g+9XL0vqzt2C1ywn8+ipV/2Po8+4J
CzIHkM7p//gUJZb9Fr3f58w3QEFgDO/fB1s6KENgJtRiygFMfvh6ddy3D64B
ZQQ9I1oC5DNJ+FvqCQxSyJxAQDFr57bmtxEYDnIBP2E0DStCd7N4bILf1mvY
+tXyrmIHaZ6k5aTFZyegTw+MMBGa7z5mhc89WP65bhOlgm8eEty25k42xJBT
m4VG1JTSl936h2VHJPqs3GLavLBtNqcV11FVxesIWq3XzfNMtG+RsCG8q+EJ
QVILQ2W9zp6EbLguwfaoHBkMYnSzZ8VrAa9RpVCPbwTEbwa4y0/GEQS3L1NY
ndAY6ZCjl7FoLCR6C+qfDDKyWrjJKVg0TzxiEl4+x/xkCLGThPyHK2CIyNRh
LaALZA1UeORFJJuJJNZpuUlGpUWGy6rzLcvImDpqE+SbF0nJTH+0SfsciVef
f9E5a1ytHUq+XUUmRNPNCjPAoB9MDNpayQygbk6oeFuQNcdhxI2vX7EQzR5N
k0+EoyoDSBaGaNil3fBgX/me6OaGo/umMwlaM2xe28EbRgAcaiQTk3C5ghI8
Mqwj+jAcYxB0a6kYURqHwNPEwaYD/6kMAmG2YwrO9Q8pMztCZ546/R2gRcWG
nQH78aSRvxaeHly/sNCqJ61vUKoczaDjUQlW4AvaLG7paU3W3gcPWyWykKBc
jklrszJHKworqNekjPen8tL0BN8X3DpDnHR1PaFqiO6LSJsVqR/GyzWWEiYK
OgWgv8BBL4VO8fJL76lbod5okXMtqCSs+TzStAcG7JQSM/6AvFVyiloOK2eF
EKv4aYiJGFWZPmPyBLEqYsHnc9anzKY3wTiTd/du069M6ByHl32crvDG1vGm
iUSFPlNT5vjEM22AVgyzB/4vFMRjwGsbD8H4yrQjKOJbbLRvVMLYqSQRH0xp
vQV8USsb/GYHrmvMkQ/yWb7Yzn7DwPJZwsvCb2uqeP2/uZFhZKsI7e+z0Jii
XF+++OSxwJdbb53k8L4LwVRQ+B0LpnLbiusfc5g+NJnnLI/Tjmjx0VoW7Dqs
2fmQQUYzf8mJf8HpF8GIyTU7mKvDU8v7alW42Dg4Jpo8GCWDI2GfPCVcFlaY
UJgRJqgYc+s0V/oq8O4sExuR44P8pDkudcUXwvgWjlvnhf0JpA2SUGaGSVUx
Kn45d+f1ZdbSoxTMxnascGraweo/z2II9/ylXLXDCiH+Rk0UDJ/xHNAQu4e+
cLHSVin/t1M2LMOgo27ymcba2I/pnzod9P0/e/ubUJQAiRaIO92gd/1xR2PJ
MXZ//dkOB6Pz2T9c4lzcfsrJIJyxtfVizKSd0LwQMlsUOTqw5ZZKYVC1BMDD
fcFUHMrlw+/iUt0Bt09J68IpnkEHnsMKiOQtp8D7GB2ZG1hJTaTBo7/+6ZL3
jJuJ99dchT/WEjA7fM9ppafmlyb9dQeYb5MsDfXyKusu87B1kEoM1SyU4MyC
R12LmMm6gUEzCi80r0IfaTZfbdFLPUqa32CKtqKZp4gXPgt7mjOqT1QTnreQ
/8pc9GIlR/ZscuNMr7QClYOH8eEXTJoRABRUyu76V2N1nZUT7wd2bAUGXbCd
FIHXQYjz2o82T5OZSRQGsVMumdxxkRCSwjwIRDeGj9urjNffeEIh2T0AM68U
cRTfNuVbdfu7LiT2U6pvzNIeKz105SWIQZWOYeDM2Qk8TK+CmQIGlOubT/p2
wSmIsRvJsfCjP+Yopvhg9RlVRm93bfTcA0KQCfcTXq6q875xdoFBHqsZO+g5
Nca7FilFu8q4g35ITUNcOpBYNCunumvmSq3ZeY6CbW9GpK4s/fYo+q11w1WI
tplPzFHU3BuHf6+mAEwyYnxcMU3BuQZBnSpL1+jcGGMhU/1U/k5z4SkILHDG
HGDRhxJR31CMTqqUvnmBcrE8t1RJn/Q6RuSudEqixmOMqkOQ/Q3awtcAO9/7
DuVEOAtVHrKfAGOCx5GEEdhBZWOsLFOcq7A1hF1UHXOM353NCaS8JQDC+P53
PHYAWN0ZXEv5OIMDupSOaFPfCW9hJ/UveJPxnx3Y8bRX88hNpH1rkA+rD8ht
jqtFPvLxWtdC8UeU48xqMMh9QV4/6x90/ecHFlRkgWv1T/dEdR1uONA2MynA
SdFJLaOlhH6CARX+Fp6pl78/2Mc5J/st5OMmy+1IMhFJEK8YDRlaDRB+NKj9
fTDkCcOLJxD0hY9k77kH7i/lCWQlVkGLx2fNJvA5FLisLqq0d2k8B04oyb/v
axbNLui7Se1J4zRrB77UNPW7K6oENUhInfaGNt1VPqR1D0WbzYOYN98xQiKm
RLx04Y/J1yAYbXWPezmIuJsQjreqoSaYLH3srtppYtOip9iDfiUKkeBgGhjz
vbNj4/Dg+1QiSw74wL/DxOf+cJj8yVxf3F6cJrVl7fTcTRkZ4O+eny78NhDg
Bw98URADRujtJdtsQEzt7j0RgPP8sgFXDhrs+oROpvft/KwvL9K7yJaN4y83
ptt8K0kx0s1a4t+WAefJriGH3R/XRjm/7qAeEB9IHe/ExB+BdTi0BIHzyavw
uz86PCeepRuiK6oQxbzfX0ZoNUM65KgrwsINBjMdq3bps3cl/Pwdx8cKsJLc
LjB4lW4x8PiFTapKwPJwxV2xOgXl9w/15lVYGY5CgxlAlJaQG+eslaWNnA0l
WsQUAnbawh12TAn/yTsjsWV9fBdeKmx/uip8864QdXnAXa/ahs5SgutgZikT
cKT76wUfR4S6q26iJYb1bMkqfhyi4oM6RjnU/WhV+Rq8wki3rnJVcvfbHjjd
Ol0yZhO4h3+GqM9/MdotvmoCq6fXGM2Vp/Jqv+afVO560WXkReKqsEIZXDSd
wyHySxUjyr4cZI30pUh87VlpZmJKF8gO22k4jOsTIC0JCDkQSmziQnHqpx8V
zhyHZrorzrdtZ7GEs0cmspiWEcLVV+K1Vm+hAcouq3WkcK8mYMytSgDSJsmR
Oy4I5TCyHr/Pf29d9sUZ0F1qLQXcF1TDr0Jy39+t3nfNDk8d33nhpvY9tgXy
uhXb8HlI2+z9QwjpaI9wCXuVPJgFdu6uCCl3DDtq1OQaQm7h4vJeeVd4lKIX
3C8dLAY1lA9U3vvptmwzSBhs56vSNfaGJVZyudU4t/OTfZ/clCcUVJEDhMB2
uPkEnoQx/m9VOQC1GVjEjqUq6Hl7sZ12f2wdbk5Bu7QmYPg4nUd1XPYGOpKI
WQ4wefbilqeSeQoY3YOifP/qHI/zT3KzfojRFWuhkoGUaC0QaOI5UGqC3exC
wCix5RRkwbij2qgrS2NsdhKZ+g3jJu18K+P0F6BS/srkakAEkERlpiVoEqu0
Da5R0FMCVMDryWrkYLn3HdtOZB0Pe0qj/6RT3pHBBv+3ZhmZA0d/PkRCC4cY
QQ5SbizORujO32onhbLQaslA4QSaC7re+ajHphMEaOD5s04INcHBqsthh7p/
/O5kYipGrDZCZfVjluxyyRrRWb0mVdUBc2Dh5rS86tm1ml3mZmuorgNkjpof
7zVe/ZRbu0wpzzNjcQRbx27ulLMYAb18plv/WHLVwbOUe1RAObMU8/D+8y3q
ngjJq1TcjAjCwJxceW27kN3VvZdy16rPsUoLwoRqM2rWuv1v/3hBLtWnyoLT
8iHn4odg9oTurOS/cK6TNhz/FccDzPJh5jblBBienZpoPm2xyjQ14hdS3drP
o5c13Vab2RrzqAgPTcB4Wr2Bb+tGNxjVwMQZvV3YmE8Qhf4ggNIz9yyzW9Dz
2+0+nZFLNKxApI57i7WVr5gwAGe2qM7iSQ1Cp3g14yaFHsSS8/KmE7YcNWQF
fx9Vz/cVs22zzd4VLLOdSEJV4AzUu2aLIiBVPg/Q+IjImSD6YbWIxWfo4avY
tCkUJkzF7WhfEocpGTWVPXG0eNjhNZEw8p1alZJq+ItvXnPUkDKUoKDVH5hE
XD6T6yVV0q/U7dq7vFtX1ogmyhsaoJFDYZhUmX4cvcg5P9o/mJvZ5QAXMwZJ
nxFLSbHJGXHQDeNydNigPFgTLM7nKZjt6Uyq+qPO/Fam7EiTm/KeNbBGDtup
LaaYPZlRHJxBZcO3cAEsdRc45Ut7AZjJO3M3vEUqdw6+nO84wOHdkyPXJs7a
bjaPWza8MJkvrTYd9U1SXeI7ne9VR4Rl3v2XvG1K3tp16R2dCtu8ncz1VIC4
RcE/lcRajtWHsJwzEy7w9vDPv5oj9phWK8UiW9/qP+M28F6gANAbTkQ0CDen
OS3EXlTx7ywez62a6t/s0sZ7KnOaMhDgUq2VY0TnIXaOt91WUrYSGFDQcYhN
NQ/rRL8aN7rivPh6jfq/MwqnMLqUv6oYA8Q39n7n6/TykDH382SHm0vfD5sq
RiKlytpci5od/cqj4V+Z//ZiFOeJ/d63pTuic6UQlshqUj//JIkCF4d6oLF6
VwTLxfjqxIQlhBGJ1ZxwXto9WrpZpT+0LAAHyXkC3cGTQ5gZC2TedBBiPhmV
6E3McaSfJRrRWsO90inHoYZ0/hlI8LEKJCqj44Yi8vX1uLkK1pvtCoJ9EFi8
f2ZbIMlLdHe7PWhl0g7mzTKQwNOu+xZqEi0PaMnrep8etw4V6ZCPMtECkgF7
2r095Px+x0x0Bq3Hl/g/r9bUZK8zoz3OE5tnS2O5emgdYO/neuULZKWaMO4b
3ttTEOOVvAYGrskBFI1XyCFa5SSPhcwjIBVJRtKxs29Wza897DfFN1B4RLs2
IPXInfWXQyrqwpGBlcbzIf5jTdiAY0kDZ0DW3GjV3jj4EE0dz/tBSM+pGSt7
wFeYPVCULsPhKjl7gCkdpcDNditCr1y45CMdY+5B4vqIZyHpT/RdC2oD1PRW
kl1OfPEv0p0hSITgwMIjhWscs70Ie0obOJZ2NDXDuqpWm0XwPsw2yHq8yAW/
WW9ocA9frfkdpU+EVSjE4F+B2VqcOkNCFhX9R7T3xLyu09oHwvnjMuGKyd3z
sHqw63vaJGpwDBkaexEYp08jFuZ5K0PJWZOFNm7ahh4fc7kBN1iw6NTVPsoA
5xJQGxI5PsuQRNLTaWKm/HZo3kfSa+3PvDycCDox53JaUBTcsmitwmUtiYSH
nVYSfx8uM31mwPvcZEBK0nqYMaqND3bVW2eqsAnMYV6zmAtZkCkvYbAwvjgq
XeZL55fQPcSe2oTsnh41tKuOVZi9TlewRc/sQey90wihyNQtKCweqGFKAsgT
scmo3jfAMDsFclbenNnCx+DOmNSQa5hzw300E71bg5l3vTwNDkp0oAxUSpBI
fHB2jD1t4AB6Y68mtllBYTJLPlbLNW6SzBaDEf/KYvebUqndLwjDjF0zSjCU
AZ1LbiWQZEHkNVCASMvPLShgegIJUbQ63V1E2EcVoZJrfeZdWyj4/j/jBrjQ
opE33R449eRUmlFJdUH79vuc0F26HhIIoqUDWhQnO1D217+QoJZ95zzDUnXz
jQbgg3FZQjdY1J8SG1dauSes83jwL4rNgSsevd/BdYXkHff5QWR20CTSQ8GP
WGRNkteMEsr4548Ck/61m4rWY3Of9WvxgEp2XzjcVxG+YhnLW/vrWONI3/QD
a4vrXt9OZJPuEkIfEWnwwj3k+wdaPmSrkJYpABdgPm3J0/KgsQMt51nQghfb
8GiUUXZUn0v6YHdGQ714kaOQBGo4I5mcDReatcHD2W2Zcj0yOObotDjZ00Tl
ekG3Tc9w9bWfWkVQrcQaxdRcifdQl9y15FuR2Ycml9+lCR0tGdZ5mhTMpB/S
5TTA5E4RPtRvfNHFCv0zArjU8w/jLkN1R7pVkAsHTOKQV98V0Y7ea9L97OrP
j+WzC6LnNQbuHeSCpOYSCeMun9ne7KQnRFh6ePtKK2XUvwWh5yv6pfBKiFUw
0pR+7gW446yimvAA5H3oSteBBaTxL/fbmdHQtVj+OZWdZPiQ9qVt4v5rkyle
CCJfW/gE8QF7d3n66uQiPWVgx4xy0eE+50oqImeDBB6nDnGlg2nQXaTlTRoz
Tds8M/SYRqGxUP3EPZyQ/xgh01hLs3NpUqYC2KCgyoMVXpdzvtfYwlzsQa3U
sjLSKp5M4J5fvUK//0w/idOcj0far1TDU//m1dgM05/L4PlUVE+4gzq/sIys
xoQdYCQKKUdMF3rSBiJGBCj7gvJt7f+uXvD1CUfR4VqTOzX59/DnNQEf+N4A
490uEiCTmT62t2wrgN12FyPYwB5e0ay+4eTKY2xAbc8Ed1gRR749zi5Ye+7w
1Jq1f0UHYvq0i5AS5JMotuTg/NKEbU3FWrXQBgKz7yY6AlVEG67ac7kG8lmg
ogGVwPECdjG9s69vg5mkJZydVpiXkRKjyLTWZOnbZGXG1UWN8ru/xXt0SKo3
jtmp1Zh914wW9VX8fhFUuv7BP1cCnxgMgPDhIjFwM0II8oTT7YWeYv/rk7Rt
0m+uaWXT2qNjrYkbOUlekiEo6s2fTOnIYhi9326hZJrmhoW59m4WieXnxSBo
ng+LEZYvSJnGO62SS218QMcX3vuoRJthf1CCnm+zjY8gs/YUTeSEu+X/rSgZ
YU3hm/Bv4bxvBpZWlxy2aDnO4aSgWu55gixHsNHr002NarjBFQrO1PyJmcQr
4gpIXE188GsX2unMdgZTJSnuP106iFO93u17uVcbs7KV9kWK4EqlioNFzTID
aw7Hpx+4yUgYCRbfvUnp740qDFARLsdfPq6dJIY/oiXqGvQU0NIyF6Ci0m/z
nWO0K6/jbKCL2ppNs2eJxVuMVYvJGKIf1k4LgG+TVoFyLtZHitgC4nXiwQ/u
Mt6JoMXT7skI/T7KSDhfx4EuuGIWZpNuT9M1YwRO9H/mlbIw0soHdjQpFpEp
LfnjLzyRihTRrfQTEqw1XN0DaGKSBBh7ZZVmEcrIyBtmY2p1xaQnO9094AVu
/ubWBO6XiuUCYc5ywLpTh7HXUUCEAdR8VIZVH3NtZ76pk+ESN5E8Yx9eob+9
r/alqf7KqgXQWoaQcXK8OmKVLdmT2uimujzh1WRlQQX9+zzdZodFYHlzeQX0
zm60nH92toMQysOJreiw3FLglPDm7I6ih5lmqlTx03vRqBRuhS6EzkvLoOU+
NPpTCbPGJRCA/SiJaKiiEDBtrBrEHjY3YCb8vk/32F4Q81KRc+wZk77Wc0iL
7L1HFOqRzV99wmcaRQN9eSJwwqX+YNk4DzMDgOQUQLd2Wfc584ugwax8PHbP
Zp594XxJZDMfyqZ+DMsLjz194EShT/T3RG+CbTXDtUw9rvUFxxAZTATiDvPC
10rP6TG6iUs/sJb0CRNgvTeOHoK1EwBvDQl0yGfgDfW1KDd99qyaZGrcx2uG
r4JcDSB4K565dbSJrS6RN3RuVLsVHSIcydv5zaNlhAQSpg5M7w4c50B9Q3iJ
LR43XKdIK0+gX7QmNDxFYYgzT5o7VnDz9TfnDPa+HOOQ9L7S0dqqHePrRJPn
q6PxRN9ZC6Tod2Dg1RZU0pNI5rVzAYKidJB2N/zoOg78S06fp6381NLsomq0
cjSOQrrOQtFBGbQmOVO9mFfYgmHv0bAEKs2d2gjHuN2u1lfscdVezpn8VNwy
2fG05T3MsagHJ/TC6YGB7sITwCWMqH5AKYID47MXcXReWJ/VKGeRX+tfvjyy
xNibs/08yjjpUp9M8s/SnVdE329etJZ0h5fbieu4Gk1NXwpr2L6FzAHWazX4
2pBZvbNfPWlvyFumsLfT9dSikW21EkGqnhO4ZQRzYeQn1qOJ8iqOg9TzASv7
Y5GD2IZhz7bIJFNv6JddN6nIdz/QSKnCzXTk3a2agRcX98t+UHzITt/HWU3R
rGYLbrgmIU++IiXSW/JDT3Pd0c0aPxZ2vRTg9UMNoQVvkATgWFiCTfwKv/4T
iSkEmZJ+PReiYDdGrn/JLdJonbIhcv4aeSXsUxa5QpqBckE0szJhAw9DQaDZ
hpvNBNy4+S4RPOHMTqrR5tvYUuwixOueRN0dUOKl5tYt0QJYbxp7HP5wIT8u
f18WV04cHV9COXj0mGsJ1pYGhaMpUBQqePd/bAxThwrCs+2zP9JibmSgFoM8
u+KQ8mUPdRU4LC2wF2kGRmWw6XveJLTvZd6uzaCEI6sGGo/ELEXCoP2CBQxM
qRbO9ys6/AusHHoAJkELSsIusftTyYqwE/LCIB9VlzPawt/Q4dR22tZygdck
8EtER8Gn+FqNgfSQHx31hreX4scTeS3kJZ3NV/8aMrgGTGf5x2OR6Yr0hE2E
5X8hhGu8LYJyzpogfN2hNpUMdQ3/xH9r9Fy7lULwn1sRfwjcA2agToTFuwQx
oF0Mxc2YyBcbUHxMlcTOcBEd89hW1zuKmMu+LXLXOaOojXetB5UA/msa8FT5
CeDWpkhwIPjzBqP4AVPdggjem5j7btCuREa9s4pfYl1JfSwWSmzgLxp43mv/
+WNZkPNW8Y1zpi0jRxzBeP/Xk1qTrmBO6iuPC1fmVQhympSzBeKXVRdrPEhM
P6RBYrocV0GWB15vtuWKAYpuZn3dHpFrKaLYiKANO6AceO7A63ZYqVmkRV4E
IgoukwT2loAMGdrllAes+AuIvujDpx92W/ZVk9HCrl0WX09y/TQt9rbGG0HT
RRRrJiPH/PTLx7jBwqTA+nUFg0t2bdF+zSMWD8SR3bfOtHqPCdsgpp1xQj9J
dAVpt6+o+m1BCb0xrjL6ln3wFV8wRBVMGiUUHVRxqPg9zFEHD4oIcv1SzB9o
GMtU8sVD+uRXhD6K5Q7D0gRJhrYE++/rmooUKWPxO8NaYJ8zb/fjklOkwXt1
KxmnuNLmgYwWAfgFbhjW/C9ViaKgNIc6SYfbw8huYTLv4Uut+xqPtGkbZIKI
0PnvWsFogg0fJLSPtJvc9g5nJMS46P3IUXMuc0DfHSYG67TAy//tP/O1b/Ck
QtFjSAuwBP4/rZuS3zyLrFmn4W50Bq1U8yO8qnFmasDaZn00kjYxshhzm5/j
A+W6qoBt4B1wgBe6WhVIH3rTm7wnCPmv2CYLrm0M30N0P6g1eq875soouZu4
lSTcc4Ql2pVFbTI2uqcOFdc+s9XFqQtpG3FUNqUsbyWYjMCK/Whxb3ZSxv2j
0CF9vGD3gGGV+IHI0qas5CeS2eTuqwfhsaDvOi9NzkW5AKvTcqumq3IMpCD2
DToWnV71YHc+DiH8f+Kui83XPVcdbkTCchS5VymtPXRCgFQA6Rb9snVbw3H2
DKDgwVymQ64THZi85XT6xa3/vhSxpo67IkIQCPtCo75vzYwxGV3eU3qa0tvg
Eha6nCvJIUM9iYaq4OBwgbrjVa5tqVGyx+7vychsWcn7Opf9Cz2VPftOvZBY
Jz2LG8QiIQRTKdOSvYZ7ScKuaOrJi1qKzXzhKLIepT0OW8Scal7I8pNjeHvn
a9zjDtVXTHqGCRKDTWisQ6Vtli8PCYDf/b8dBxBnW+iM0WxChz2PENVsJThp
/dMF3BjImh+xP6SEO++tIiUY02MNvD09yPJoOn74KM9aOaESqKPMhI/3sHX5
ahvSUDK6JotnwdHlKZ880Um6uEEfQAaPUTCC0PhXGZbJPr9jUY1dUs01w4Hy
BuwNwPFuIEv1vCl+3bbfp2f46B4VkHx03k9geMOd3Tx71iYFgCZuYB78R4IG
a7V/9LzFg3UiBLUeTo0E4xFf90uAzJVAdDpkN3RHXFTgUX0F3SAOJhta/y2s
d8UveTChDZd8iP9mAWch19O6YyGCvasEUnFIr8w24OBIi6SiCCUTpGQubt1U
4vwa+/G8c6pF6I3bg66Sg0D2RhAO9K8mb67liHTThNt5MVSeUgO1glzYQp3m
yFIrLdOfk3FOigrl2SmaCcQvs3kRfOitVfFOqAwjvTdt1jN30LXlIVqwxYwX
NNsNzPe+a4HN2/Xw4NN5+NMXCm4CzbnSIbd0djr4uK8/ihwhRd5OuK7WfkLe
SreBS/PaFgL5BT8qF8SebYu59LmjrhRnhw4p2EowHmHNslR2p6Y5EHWJmRdl
YUtWygH5kb/GyzT6eJX1zxV89kfqjq29Re5iOi6CJxVIjXvj4HQERnsBYnyp
UNc/7+t9PIa+nNyaIqvVUqd6ukeJD/ZYp4IY8NvGTKfvFtz98AxaY8z5l4Eo
5ZtztEeEcoHEQENWUMIBdfBsiq5Xr4Aj8ATbOmrg3lZGmNqxs4p+8rJrsNU2
4/8MbauJAbYkCGCeYVidBZY+ywZPAp/s6TrxIRkbhWjDuctHCBm4WuWOrv9x
uGZ66xcXR/GdIB97LyEm0j3NCpO4MQpaHicB7vs5k3J0TxArpoV6R+4DN+8N
6h10d9dKZ9PV6HeXCRy6QE4dP59gkDdDQmfbGHbJuk227Z0xnmowGN5GNRxQ
PURdarPkKrDjtTHMObrwVFKLETQ6LGXuHdcS11OVhTKXTuIjCQnUheRdTCZ4
ItOEbp+YpUflAX0SKFCp2+lSaaU7uC40xd3R+7ctgKVSevFI/IDODMxDEuHJ
SgBM3YURKP+ISfL63ECnw3BAp/+dA6zSD0XA4IrIjr5I3oUwNeXqs8uMGCoZ
B0YZBZe5BOrl5OAwP+0erbc6Zrw12Sbt+Hsjz2EpfEhOSGhhCrU6tjCjvG5K
uECJxfx1X4Q4rrKzH9yzvz+SY5gsrWmVAXHPEq+k6uZpLO0aWwszSl/R0lGj
33pG/+nQ9Hoa0ro9io/SVhKGHTzfWVxQz/nSUH0N24d7ILD2yNtnOzjX0muY
hrfZMIah2xEP78kehxE0VLUz/V8DVqts3wXGX62GAcTrNa7S1Mm6p8//eXLR
7ZRNu3U5PwV3Zm2gzRF5bNvfkgKn0ZK9rgTwz/tI5JzUn6fC04kRyiAa2AmG
xwULK9IwgrKQNmA2dW7mBuxtwGB56UgEXtFADXaD1AiqMpfBQJnQs+RmkogV
oq5jB4JPcET5lm82fLLfikQpRcIUTiM54rpLurbl/RO+DrBpQnOng8fv3ftZ
D71Q8Zae+gLsla52IVCqm96rQi7hHVSI+A5JIclZXqWx1ecuRdJ5eV1y+zbX
z2kA5yDs5pmlyDQ5HvLbXL3L7XEBsMsE8E5sC9f8FzDQel4C52RhxPBaefIH
yh/tIGHx/MdRlQlRHFEHw393jjYyP9vjqSF/s5f3zugMNrTpnyPquMmTfc12
5ymqfT/IarWfKH91q97BH4iyrBf0LEUVfYqZ4PpMFF3ukJuRVvFftRy16eKE
yNnQS3MstuQlSdLTOSD/stLyeDBxkZr7T6e3x5Sw1jhmoIYuIFAr1cOMSmS7
7T+KeTInuY1foJGbBB06W4QdCfotYlvvEYoUrTq4MCn1g1ikGzDYp+ibmM2W
vlFbdQmCAV/6auiMj4MOzVV54BhNiGvQ4dNo8XrEvlKS4bQRClFFn6G8CLXs
KTXI8tD74+aLRZ+1yuKUUlyqWcMESA/0+CK6UP0RPhZ89FV/Aae2K3LvbE3I
kJuTQSrJXpCZ8Uy8pJ6Z2kx0g0DslPZ7Kj9SqLS9euGj5LjC/Id/UM4ywSuF
9ByPtGfEeLdB7Gq18Opgp5Cj0y6agJphlUqAR1A/xb9uKrekUKmmdTQlTHgS
ImIkAjojaKWgCLRx/4nXv++THUPXXhoRq7PalI6oSlnCZQN45Aed9m7NcxTs
eTifUbprfRYTDC9uon19u8JAcaYAP0F3rsd4tx3PbcsJTud93KdEnTj9hI+v
VU0HnNUPvEAPPa7HOdFTEfKqkpJjlLmRNjeU/VueoYl2Vg/pToUIQaTmGv+k
jIWKEPp1LzvLavBmEaHfj//ujJ602cfbP2uZia/edeON5XhX7sA8IP7fbfRz
0u/UT2VLBAMDhB0ZAf2SfupQiqMvM9V5QNhwvQK+22xkGQrJDzAHU5Ml/T4L
5gSRi7/GUL21Upi47xOvMfBBJpMWUxQBseMEfVCuzm84kTJHF39V/dcAEkOF
f2Jcg00k5GJrT+MEcmcJe84swHYpFje5hAvjh7MRyT890sR36cpzCwGL/sNb
hhps6pVbEvaeI+fVjnbV+YsOS5Ki3TJQdHLvz8Fq4AFtHfcfPqtw1gGgu0lH
EwlFDaVlL3CJyQYUuIcHD2JS35MpvteKKzgwMkl4aXbKPoBzYf55ILFQ8F88
6pbL9y8pW3L5Z64hj5kud053VS5qJMJ3VtbJX6Gwyj+ZuOA/HyLXZTrkP4zb
hfHUXTxoKfY20PQpiKb6Qi3p+6XXKAaulDkIDHAktCrJKdvMdpJcGMMDqFnK
e6fP9VPZ9NYlmFZXNP0/I7qfhu80nLI6afwtoXBYXtVsNwm8feYbLAIztWFD
IacN8m6JwcsAu/ncjjFTMTqECycRS9zBG4wdaM32lwSwvmmd7wMOdkmu+pLq
GXkXad3pGqU5NlxR5jzgc6UOpwtkOCKvSltUYEyyhsV5SyRpHbKWH0Q0v+/T
SmLzL06MHkXhf9iQ6DHMbWJBPn+2uZ9tE5ftuYOppU0xotWSaj2fdBHFLTb9
8aVd/+9q04k3lhADR2jxXWK6pyw5ohjmFeVIxT2dq38dKNwQg3xkt2AaSL4a
CGwp7ENPUEiuia9s6ud7CGd+AiQESp0gRIxbF2fsVqT7J02esP+GSWO/imJ1
fqep8ZmvLCjsAjxO8YCBLF/TYkfOEfe/MPQHIBefoLkHwWG7MhGhoQEiFguA
6AHDKiKe+4DI1Kdj/MBC1fKqbLmtlqX8+UzpOKmRXbRw6jkIvKlIm7pZyroz
rZRpK5OkGuEzjayHZjUVwY6R7AMxAK6U8Md9KwtTaoRmGpQ0VsQqQIP2OtB+
DhxpI/G+vSpxePHFKC9pnxcSh+a4A45251bJhs/aAVo1J1btoPUIVAYe19OE
X60leqTS28M7hqkpItlOQvBr4ENBGqc5T422NEOZymqWcU2hIVlpJ6RBb7I5
DGg4rEpvMnZ53bDzosGBitQ5ojya0/hfkTbQSmmJuS0ncy8wWzBMYA9oVaHs
1UA83H2K8+oP88I7wrzdA+hh6oZfesihicditcKbFZNQhiX93QwLulJqSMf+
jEvLh4lHg+yadz7kjBaVDC51KxOBtPp3TUb2HN2LJLzpOU+ws9e9jlOofRLS
FJyHi8pSXwYmxRmA0A/nQlF0iPL0QYjN/QaNVAnG10Is138/KXBUv2fBGF8V
hxw6hJe9YdhTdX8Pria+G5KCFHER5hDJeViCwVYO8HUOwrDLDYCBIu3ssPP8
hO29zXKO6sshv09nnrpUK9dIAvkmM6dp9094QE/v2rz89UNcyHSAhQV0uK31
8ko89HvcdyyLlG+PLQbl5JBWk4aKcjs72dkNk+4gW7abrEwVm1kjbdYAhj0h
sGqA0YlvISCbcdKT86oKaUqkhux7PRcsrYZ4JhlFGKRDKIizCDYqUHfldW3O
jbK9fjOfz2PMaZx95n7exUisuvOK/d++kkBLKmBmH7tVj5djy7KpEWkWrjDZ
RWQqE1oXy+VrAF74Nf1U4rs97Cmd/aSQaa5zspjRn298R1OFtnr9H6ujJf0k
pKkpiZSmieTDf4R2Q8qc4mSiJRisGfNbDuKy7Afww3sb6IH8J+XKCaTjmq/e
/mH6fCqwdncH5Rll/B/ORdzdUeXYGFx+f0s70TB9B7/Axqvv+KxmgWfDd9ij
OcJiEwhXfCt5z9Xh1kTPgtKa3LB1v54+mxTYmp7ZDGt87egN/+JKl65b6NTW
kxW1scBcPsL2myTtjq42LOdZz3UQUxXJJYtAQaKxpcDLUi6956nWvy7031J4
Zn61xfTI6ZnGBnLezQgfMu9ZUvZVXipwcsvZZJ7iKJbKgSZDibc6EPPrG0Bw
pzbWVD97632K7Ox9+vUVCRe6JbSAEucM1n1TXhe5+xT7rx9swq/NqswngP5B
vbCmsd/3uM7CoTsayrMkmRmJFiGYzONsJmyJ+gFI3LuK2Mbe+6M08Y7Ff01g
hL4CTbAGQdPLZwHZPWAk6m2ABbq2hyWMIzC2BDA99a8PDdsarKpWsFV+rybA
bydWpmzEPyq1ksEOXoWY9dKrvYYNuHxnVbUPkGvrkrvr+whhPppx+fQzcxSu
DjEV/Ml1vs9JLd9HDlfdj0UPGMP63IOulrjw/CerDIn5yIowRxRk4S0K68Qj
FxgH/a11N59oZD30blDlNgZ3BQlqxrnIkJvJY/h+KMuoO8qsVZ753byn3VB9
emqzbTkbADTUwXZZ5TpRJsF98rCZ//ZU5Z0KsZCgpVtZAcoF9oNeon8dKFjH
fSGkTJ3Som30LJistZIdHtpSh6flqQc4FFaA0vK7TtjXJMxD8SV014tBouzt
GZD5obezq3En1akbXjcUiNj6RjVSoLc6lcQmm8eLffQxzgnYn3PWQBTlhSZT
6XYR/GYEfhfBena60HGzfHyLBHDk4wMtKAgwqtikHFIdvSrh0ooUpzLb6uRI
dEp2+ZJDCdT5f4R6RdVEae4uMISYOH/TuVnG4EoQ1S+OBYvCzJhETfd9D0JB
EUYml1qRnCWlA+Hvm99w/pcXaDdz0913s0EZ2JqkCjsOZazcoAPkrbciO+Xp
ruoFF5Hq4JUZGSq7fL58h1aXueXS4tqvxUeacTz1JEPuafoxLw9SBpmBo60T
+Huetb/pJ+ltO07VC5J1sXX584qIYQQv6Xhn0uAz7VlORynqxq8DIAZcgZjY
wCprvvOUs6I8/OKkHvGHfJ37sVDf92nRa2i+kfKQ8OHWuw+NVMrj0qw1rVNG
KVC895b6plZH6xSP9x+nBH6ZH8I9aioZCL7ZqOJXgAKl6Y1jr2cjZ18tftJI
2sgG2gyna5cdCBVYdjYj/er6bucKs+oe7ailJx4234IfHjiMlPoHzXjIcPdf
jrk9qFDmWU/bp2OrjSYjwaiSSkdh9U81beBaSn/6xGgeFo4AC/tftDjw+rIy
Phv1WG+uZBwytpdhY//baw0uqsCEZE2v6cBt2nyxaeD9KaJLluUFKFFPe/wf
L+ZmRMfQPDa4Goci6URGm8QatSqi2UIogmQfKJAY8BaHSW70rZEQr3GxAPfE
sRHQkpi2T6xHrTKANX1LsAAvCZ018aWjtVjxnhbAFO4k2hV81eKYnP6xTg5L
XtnXDHwwKKxhUGRfd4aAh49l+rEAiVqjF506rc0XfZE1b2VTow/jxOs5z3Uj
LvishLTN2ul18xRAhOJKXCc72qbCVqsyi8pUdpfU3jpQXI23M0pOtyYJt9W6
QziMq56TVxW65TR1wKpqCXz2C6C+F+G5LoERLmzkrDKaWY6ujNmD3pKoOkg/
sHOAN1u1STje/UFegcnjZ93RjUrNGxFZq/cSiFkbkku6KDF4iQjuW+z/FTOY
ldOjIeq1924x1YstS5o6MZaTf7p9wFcIcuNuaKm0IKJ7W8Auxkg1sbrQzhf2
dI1EXZQTzKKhttrLAQtBSLTFgwfxRtM4o1JC81oEJbYCuq9WhqLJQYcC3oNh
ts3YIi/AmFStYeAvhIJOiSBb2v24oGJ487DUfZmzsrlUIO6okBUGCt7yD+/f
q7YcCd1M3Vo7xoLdxcRty6dKHOiDy92GXJEsl76NOoGwDrcm8RmcCCa3AxOX
FiDWcmaumUgJbZKPnGPWBpnSiHxO1phbqDI/z9PY+Y+XtMPaxjvn7B/Mel5b
bAwKbqkfefa6I6Y5fPKyFzliAdEgUSOQAIeJany4LL0h/YYXL3LlgRtDzArH
KFZn4dcroSr8mdkLVfXwViG4k07AVYXI6iq73gFd2zCyq0S0jxQgIVz+0TSX
+MrRwPk8MmWozCc/2+hNHxU4E8WnuuZXzf98CddoGmrQ0/CcUGzJmBVs5SDq
sJlq26HNBTScfwngnXeIc05/9aqkRu1kmyY2Qj/ke8EXbyJNYq4W8+HQKcfe
jt+P/rm7apaL7zcCCIkKWx1v3v9+8XBKq2g9GmtUzN8nJ+SRRf3Yd70DTnCj
4Q/ZmZWKC1WVVEK2d6XGYuQBFgu/6pxQZhbamawr374aYFfYoNObyhrjjMTB
MoW67CWEKn+eNRsj5rqJ3NJPfKYdNcHguDwGYpD7d3qwV9PTAlYqShE6rz7p
5SRRWnzPP+7wcHHDh8doiky5CeklxgNa/Jl07TV5s0WrJxIYXY2/lE5n/pcc
baFrl8aDscQm8g8YFJJvelON0J/AhAAqi2JY9bNDkGF8Lek4gA2La/nGF6yI
aRhgaLZdYVje6qmadhD6c7DsAzxKH2fZEdMh4/HjB86daxZQIYS/w4JytLhF
XjtfC5H2sTNj7UcxLN0eQEUaPIDFqhjFw4NIGPjQgqhLqEd9M8GM3r25yieZ
EViLueh/31Bt9zVIEQCNXCNSHokVALtSQ/uhk/ZCWUlB3kMJdfblKIw5Tkm8
GpQTBfFglg9DY2WXwwQwLaR/j7gB2zKVR0BezOB1vQgdosGZMKH5L6QPNQrg
AzxK7GGDVcIDb/k1eJQsNAKDrA6vZBVEE+rf3fG6QFqKcYqmDF/azMZtEOsa
SOZlh5W63FxPcc3w9BMsaD8LKxKjukc73zCBsj/1YDLgBhHQcQlmSNmPh59h
lSMfnW8SCDydp+6CNE+acWWlQm3I6oNiY9lwQqnPlyAGOt5kqiY7jVHGCymW
qXqj76lQxXMe8CaiXgcQo2M8Vvgr4y5oU/gQdP67yf3/X5myzDx8L4YIqoAS
SKLfxcyKCmObhJ8B4Dm+kKUvEkpe9bl0/VE9gbY7fvbesmvRTQqQ2DpuN0zc
MsfIvx7emDEWjQRGLC+FreEEGqQfTDqeJ0PDEkKC0L/Jh74OhNBoKbEv99dR
UlL5NDum37OqZnDUYscynEU7oMHKdC2GuZQ8vzjFpJdyPbRAtgXw/PQhR3eD
kpdns+C4rLDjdSMBDREwVU6V06o8p4Zd3M6gInQj+7RaIfyGEpsVqAkxlZ/0
Y/qjvgNWJFND9D1FQbCNG4P9kCYuZCG2Mk3I3JUWya0wv3PVqFOTMHWg85AC
ZR+GOipKnaecBQBbF19o1vKAw76yzJPtpXFWZXEhi3OjMPnkKNZuaAnd6LV7
CgY8HfBivYn2svihAIMf2PhFoyXpD1QpaFGxdBmRKYDkCkARK3JAGEbPXVGS
kTlWgfwtVJvP7CA3nq9YZMTlLt4voOxq1MWBv06s2+n3I3lZdnYX7kZ+bACg
Ggf4cChJCg3ssP+ZsS3qN3rGhvllU0D7XyS9REXL4U7tZaGiXQ4X4omb6wsD
znbE/5jYKqKdES6rp/benEQG7xiGAgJHxVPCJmBkSjGKu0N9u2Z/q1l1yoKa
7ChqEOoGzh0LAHiEBa2d5jzOZq7qpgm93p6pNrRdGKadxcPYnwMxAUCNfXfe
W2r464OJIjyZ4Zf4mT0H0a9jRtbdmK6XG+3o2+8wyoTRRgNpcOy8a/6NvpIl
OB4plVUemZv2EJHbpasODekmvs0HbVSNe18XuzA5LzLtJ/l1W4QHy91+6N6j
y1556sRYxA3J62JCYW5xXBurZWvPhzemBxTDg6hs3VAFRehcW2K7DbSg0lD3
RI0L8gZ9nJWEPh5s8p6ng8rPY11oCImBDueQ+wbW/Qw5+VEjbsRlhQ9KGzdV
NkDXXSJGYaageVls4SLrty2XJNqzQgE4k36zQbgnswBctXBWiyG2gsLZy/7P
1oY1Vted5zJ5UUzYgdqDBgjD17GmkqFUeAtwTqGTxqhsQEco9+eETxhlj4AI
m/OEPdU8cxpO68UsBK86l4gbyQ2W/okC0jiu6SWVye7rAUqs1YbDgrECaNzF
TpiyZpR8MhkKwmVAQtyP/PE+tKHAJYUho2NbOy6dPIJxH1G5C/mLxrGsZww7
aZqgfBlqAeNvErfwl0j+hYB71Qj9o6YrP4FOSR0MFJWlaq3RmwOp7OUuJpS6
p+q1ebHxZsaJ+9ryhCcJJ6eXk0iE8GyCR6D7/Bo2MASDvZ/TsP/czxE+yywK
+r8FNlOeWZVzUbrslTwoXAug+wmr7B8Yz4nYaq22zI7A3rkwc0f+LVmGRf8C
8YGhxM5Xum/moHefK35KJHk+OibaD/ewsMSEroSKsPuggwPf5/gXeGwNDd3e
+x+Uvh71lhL1Fk/Np5FQXCMuh01CrLYQWJaodrDKLXsN4gMclAFg7crSyp8g
UEyaW+wYxYHLBC19NPzG2yCbx8MAYp/nDPzRHfskfSohiF8UzI3viSWpu3qZ
XtKCJSH8W4JHnsI8tR5RepHQSn8AwbA3lvVYlCqoI3cWhCD9x9RxT1l+AhaU
Z5QnAsLqID4SAmGaFmPMC8r49nc2skXhtUKPrEGu+6bks5FSsHXfAAKjqMaa
V+3bwJfkLv9ljWzA9Fdm/EvzCEsJh8JIl27H+M9so1KbRNEjZLhu++nFj1jl
dz5zKIIZ+QY1wDymKIrEt27VBWnFuZkDw9VAxzSCEwd1CqQMLdWiW+m0JDOj
iAE7J++D1RR4w1nY/DSGT5HIurJJOx8vGN9iWpbJ4z41FjwUBFU1MggdT+nu
2exDAntpckW6BH4lfSQBlu/vjOrt0QdKLc+7+DZAufxLf+su2zhPr9rY6taH
eTDzNbQvFuMYpVhOBOolZHNBN2d8CpQWsu95OnvRwaG0Y8kiyjp/MHpRJWvy
AquLGBipuOdFeCi0+9HUyle0bvDdgBklxq+poOOAJiTxy6i0aGSA+SAjJG1M
tb0qTR578apPpBLjugrkrajjhwxiswPDEyn/iB8z9ncBHTA/gFdc0ekM63bJ
/Tdkl9QlnV9D644rQR3tUTv4eMqmA5liWvK12GGb1etOFQQS2AAI7LGCsRpz
79LvBDvUFT502FUR6Wr+TYk6/pKRTj8ivFV79NvWvbXGCr+SsIYZbAIzDHNE
0pMf0km9neUI4cGEPSHYhgCLIa/vVwxrEklOUqJ4PzsDVoBgT3Wj2PUvKnc7
nyT+F+U/ACE/9wRCAZjRPc/0Tzu3rplnw0qp/XKgQIDtlWucHPa2raipCJOi
2H3VCOETh9cTGhkGv0bLpgx0f5rQtZO8udTSon+dckGDnUu0/dh/+akgiAT8
o+7BkjrunRY2DYEGb5Bg8PEQmKxHWJS6+7+kk/NGscynICRYRcm4QS6xPHdr
4DPaRS+CHMrPtqip8NkOb2Zj8DP0XhGoibPfGwc9Qt9X3owzThWji/g7tTky
vk988JYnU9VaRxYOtp+cwRZE2he5ixa2BxOgwXP3d//VgDTNWc93Ag4O0X8r
z34HrC0oa98Zu5fbohSSwqskqD0P6l+SQ/+L4tk2xwptzZGgeMIYBDi6VERP
+IG5eeL2OeORr2JD5vPB+4gg3MzBB4WFNY0hZM/5tdwRHhy6w0qR7+cbH3H9
y+uwKXJJaBHv6vvgdbqL9ti1vQR936SD7J9UChr5yR47eoHAlOtf17iPq6MN
bVhblfI0YNO+KVP+6RmjLsSU0Uc9dDTYzCT6uMmCYFy4MteQXxPn+JHx2xt1
KHThWgOcbW14sfQbhMk1sJkaxXzP83kzTTMWSTcWqTVq93bQyBoskntGa4iz
FX6uN5s89LZCqKOZ1sLzIZucO7MOe1TOP0AKTC6YoJ6ZUx6sWohr7EtosbFY
t55YORKWrMOoCSgZhxaCXZpggL8VBrMj6NwgZW108gtQyZzsyXErUkMMgOlx
qqC/Pe3I9UTr5suxbnGvRFvhEsJMllDDhSn5rOQtrSwK1U2qdM3LJbTEOUCa
verFoMsBZwpQBJWHfO7RbUGfhutvVeyE2MOZFKiiUacCbsRYMoG8lX9HTQ20
l9yJlfAPhrXLqR+LMtHCyT+R627JvfyTvHu6mVlLwcoYf7qKRKHYTzeaQtNj
S6ZkCNLVsYh7wQVwletG8u9xRaS8mLBdsCZQpfgLuZRZQWRDIdDeHCbvSFlA
zL9m68wVEg68eO5vbBn+j9kVJ6IycutezFDDuMPxwWeN1V2TGYX55V6cRDUB
Y0yZD1UVn5RW8g3Uh+75lRlYXF8qvtmMOm/bPfZygMTCdPlz8apOKCTSnJqo
gjMwn59v6JY0p7eUYo7pvpGkQvvqdoAI5s40MQVLeaPrqV3PxAacaAAPwS8u
mWep9EmFBxPTHCWeH5LUwXENIoC9dp6qmKZIl9ZrBB/txjs8p3XMM32u8Cbx
/n9q001QPq3lozKWpg2eJtqJtX9nhqdTOWlTILWh4KtGdvQYCPShAA6SjaI8
8iNDeIv0TTctCk9kIAM4p86+o9CW9qknGGMbpFuD5U3iKs0zyPd0SESxVd6a
JUlzC9GCD8MK0T/8njgiNDh8QzN9XiYFXKzvNPz9fQ/pN2k+BvHf8CngPScK
d5QInc1fP76pp1VJBcuUNnH/XJGr2pu02QD/oEjhUjN4cJ07HrOKmxC7lw3O
zH/0yyhde3I8KypU1awgzMGcwnhyU+Q9YBlZUIDGYvAyd5/ufmyYJ4FiuNUq
Pd7TXLbL1G+8eW3qaMpHq8WELHt/4jU/ffUaOT4RDylJdWBWVk4kfTyTmsnu
5VM6HqfwbhxmWhpF8cms2v5L0KSfsnf/u2TzzLqMCpzS3B9RvF/FfV2PCsmn
ZUlz/1QPtak1zfNtg82t4nFxBX9+MN1E/WKiqCH/hqUXImyvMkrvvXaANsvb
99YSSytv9YFf3sUuAwDhxIW0x1YGubgWXdF2A+nmiB5dZotCtc9w+/gdWaHh
BIlgcEGphHj78F/F8DcoTrjen071xb5gXF2ok54kTzuF16Qotzc5X8ayfB1H
qdNgjbf9sPsuenelnRgCLUwLo4QH4hlxHcDcdSwbnpjRSiSFniJT5++emRRl
nycLV5NwK+kxCPOIz1vYLjXUBkHqmLqrRsl4X6H9uawNOGKm8rgMeD9KI9ZQ
TzaoWhZ836kjr/7TPFzKITt8H/v8onxwNgu9QVWu5T1N/BaA0Bl3K1vIADEe
Alh/FK0waN4pV7MfDvgdJy42VahMNbl0l3KjFu++yignBwHTxoRxWKgjO9pf
P1ZfLRLfBbXsXiZbuY6YgU7xOhJVSRsOb7ErKGWmwcCXh6r5kmZ5mRRbj3MQ
nDVxFApLYhn7wT2M7cSlD71eZF1h5yH8JgAfC3n9bhdODa7v8r9b91U+gBU3
oZaLS+70P666BLriySjeSYCjXBynW6qGS/A9Q1ktZbhDtl5nkedIcJxeT988
B6oWO3fvuCCtYT3tAxtUuGmQBQp4kt/F/g+b7YqKZi2+KhEHCpdhkmgpDI6h
VfvQa0lfXvUYTXQcozVyShaPRzGU0+dVlIUqr8ubFEWY8Pz7dvCPbVsdKEt0
DKtHARxLy5+9y455dEPMo/DrXlwckQBrHxR2fYNFGMVejaRx9N9wixEy7BDH
g3orypz0AfKRQ4Y06x4VsRRSo3f9dCDW/TAedLdky2QvHECQxmUoJ0vxMnlC
OPn9ePyko6FTLTsi3jBEaEu0f8nRAcOq41PaWAUKSZsVx6V+lsyJDjW91mar
TO6/TEf9QDu0D1mxx4LD3V3pHXZrI8lEVBY9xqXYQ03Z2BzLY7JbZWP5Yd7A
n+GuOkO/xdovO+Ne1B6dbg38VSkc4N/WzosNJrtB5hnfKWlIbSgawXajKmP6
XqgsrO6ynL9F9/sCdz2uBSt/xrccHxsPGqm8SegDMfUypSRtwBnsIGDUUtDj
yrXn0744VHGDKsoOAsaafh+c4g8SV7JOIrmwKKUmXlSk2Fk8JBamDLDpOX47
QKN2Rxv/HNoinprsV3gOr0k0SqSVGCyzjkXcl/d/4BPBBElbeltVTbQvl6f/
hz91KfK9x0arxPDglu/YX6u7ZMf7IyzSywgitH5K5rF5Iqrw5+DrgDu0Wt9+
+viQCFOFQGmLqiw8pxGTlku7ic+71jSoxvE3/SCqL4pJVbq1Y//wDNKfVVlm
D3zS/OIWxoNoQh+5A55CXvngh3j88fyrmIkEqE9ZbvKbspzKB/0dcWzrjQYC
/EdIRArYk4GMJJ4WZYzKAPlGP8eNVDIbZat9JFQrk1sj56zmSgzUzHgKiiuF
tTIYbDZaq/MefjlW2+SfbAo53iRKVGXSh8bWnv8N/amF6HkrMl+H2cc+M/E1
zRrD0UoeEKrwfGo7n+6SXbJDh2DnAst5IPEtkZ8oHbJfVIGeGKr29chkch8c
bIlW7JMIckrN9uzfSjEAc+ntfOfG5YBNTUld7YZq/xCi78IpHPJKZgCCwdFK
8TkktAxqXSIflwcIdD2vX3OXru6n+54aY0Hs/aPV/6fSNvvxz9hpJrOFWCsh
jX5v4yXg8fpGlMbkpWW19DbvNRORLPZjXwoQSpWfXrEe2rQhBHh6tnaEI5Wt
xG8w5HBN5TfHEmhZ19qltv/qMBuUMomfNFm96dyScA2/1c+sk2kHJWbXgdDO
GXzhbxuDruvP5MZ+PlUl5SMjJtGLSXZCMlcVSSKrBQA/X/QKV5lNFMdLTzhz
ZFYQee35rNOu6OK9jB62RiTbqqktzyP9XyegDlE4Ovd8aaCuxkjXMP/vQtTL
ZvB1yEQK4WQGWmHxmQRfgslCYuTDETPiiQO79vaQT1w4GWtlgLbgJs/liaXD
dbGSeSGWfp5WzYEd97UePHgVGPjbDc9erqS71BF9/IcL/mxIUfBTAokblFRJ
b84gq2JGpMEbxCFE4ZZHiIh4w0OIirOw9DExWsbcLz5KsZT1/KGj3oIXY0x5
e2HHWzCb9mKA5urKRsiOcpli6cDA/A9nG/kPlSwV4byWMO9Mj7D9vsfGpvVT
kLK2Homu2uzY4VSQUCdYduZQRa3uQ2NbSNqOccfvSEUPGgFai2CScs4fKpXW
tzdZIKmyAmfMgDxPt+JIV/gqVJFUhOtAt3/7Qo3GqN/P0QHU7T+dXz6qgiag
h2f5zCxyTWLv5Ay8bn+FUXZkWteqK2Gt1mdTKAfZpPcv1bIso0Lwm9aF8pla
7b7muYO6Ft97pB44A2BvCtnAaIvAiJREj7pBbFgPntU28zFLRlAkX4nnYDdK
90DJm5EJ/8YdF8qHvVT929LtWTYVz03TPo3Ucq6Bes3tcLSUgxbDADz/KQ7E
D8ywgoRKLjhfigFY2KqIlduaM1xD4gXUxhbWEioNIDsEOXUy25I0iR/4EsDp
3Anj8OoxoQkY5GL4LF/r6VhzY4nOF9wNlTuPKdlO5/IJN17aw1jzpgCV1HZE
GeyvKbv7/bp5OcBPkMfVLamTzS/DHsBg0tccjPtS79XxBiVKcwytypDIwAnA
eyb3tEf19dowCwqnaOheLXOMmwlRwJsKbMZBgHv7MZPkuc/+VMEn7w5sEkzO
CtiRRJ0jdxSxKCi/UbqkCFrxU13N5wD71HDBvo8dtbNc3PhRrg2VPKDUwWhc
w2rU0AgZISZuBsUSPZ3YuNwLRS9VU+jHgKiblEV0X6iBp+nm1ALwfemSUrlf
O9Le/Tu80O/Mkl47bwOr+xrqC1SJ6Mb6gMozl6Z8M6rLbYLGu2TdHu6rC8b8
0WkhHDidI3xR0KPcRDmr4Hu+qNX/UEeCG/TiYT/S75Ozv5vQ3BY80GcvopLg
3lCrKdfAfj+CD6LNosH0ufgcdqJGLx19adr8IoenLNWR9tWtXLrHQQnWGc7K
CVqhavBs8joO3GtuJ6drtYOwLaAIoacYipDC+gktlOkVbXLpH0kwTLbnHtJx
Eux4u5z0mRiy0ZoAkZzvecKda1QKIqXOQ2t4KB94l7DI0u0P6b8/WAPS4vlj
PFgwnilQt20EqAs6VZxZtZV+gE4JmAVbzg6UXZx6+QvE0hmsE5Ya4owNeuww
ErPY36OdftSAaeA1FjIVYxlqRmmru2IhnwuCp+cqPvBKv2hWen/IE3Tl8dwR
OEPVWvGWcNx8YVqO/QnAerMeJC0csv06KTtq4++RZj1on6IWzeqVLVGnS2wo
ugDw6gIJ96D3h618TKEZBgjfBsJlCKtrvxAJTFz52bff92I4LSiGxWzbAJ8i
UN3VpRuzan222CXZr8aB8zO+964E1zEwdPZe6ncgv/AJ+/23GaCNJ5/QVaoU
1obrKHDI4Exb+Asb992dwGRrhmD3qNn5gI3Cr7P4Bz/HLvB2CrBQEs+2Yj6D
avHCFDdtR2iM06Tqi7D7Wvl47+3xyduLByJMsPG4MpXZlDxwJXPW1+gB+qrn
5vYXuYQuHzghyAfBkz1wR5rH5xGdsM1PBvEMVdkNb4NQ0ojt/BxI8J/E1kql
ID3y+WkvfGvVRVpmb2vq4N3A3LMGYySF1JETuZtnJ+rqjn4VOZItRSjzyefk
V05BcKuHyN1QGKp8E68IdndrYI+DwN0NFeihaKTb9cL4e00s21uhL8jE6XV4
zd0pT5VHqSzKjaF53dnGIsmCg1cd/VcgkKMAx9uZhVGXgbTuxTSVlbrI0aIG
e0ctiN7Pj7y3qjXpiu0/gz6muT+Z2mTPL7W4AWcXCqBB+/B9Ghj28onVSujj
kgpArf+CkP2qBuCc3OT67cuCfrp5IaGobfzn2DPr+1BX/8n7oPbOBqDaRCMF
+hZlvhrQz6hk0P4Isy3AkVBGzfCKwd0Q1kabnPGiGJVCUUNGpYrx3W4ua3Iu
w8Nw3pTowkxOFhHjsbecJL2ygSrgC4omUbGjCRksRlq6DyYF2uVoBxq8Gg98
SajvbF6diPhgc6qhEcpkrDd5/Dqa+HGZtgrAlJRift2qD7XuD+mCd9Y6Yogt
33GKFzt7ju77qs/S9I8vNPwKBf8aZGqW1nw5w0szAv8VoxCeqIjaV+T7rAfq
mEknwax/zIom1bHvtkT6cQS+hoq65uJG4dOApDxliBpLJXLuQAn4Hf43hvA0
bTRciUWY2t8Jv6oSmhPO40Zf2LIvR11xK52vGxnnhy9RDfGVgMlD+JyeDmxo
GwbwBAUWr1l2LMFHCixlLWcANof91VFk+/3uFkJ5b1ABcXh8fI3vzujwML4r
gNLhE1jFobazsyUmuQTtjTeZS6PxAzhAS9DgZshrA+D0OSpEFkYk+xJKKsqM
71c544ApDSxiZx8Pzsc36r1B8yG7TEkyfQ39u+Z7sjk13iFjwzcvSOVcnobt
ihUwCUoWjhPOAHZ1bVlVq3l3BwkhsqIww+rUjkkMlmR6AkVWkjAvwR0ZFNRy
OvknaXe2ScLFkE7fIscbXFLNUAIWNTu/uk26aat3Mw6tC+lI7sOyOH5u46eY
dBNtWgrktfxKeYUWuA3jjVVUZMhGvbXdDO5AlU2vuw5or+LsKchSi8Lcedvb
XGTgXaWML0qH06BgaRAaqJ02vlSQRHKIS0qwd6JSKpbF6YcvFsDJQQbhcuyi
0NSAaOqEBijQFQhyTS9FRHMrFwhAEoVZ7ErZ67ib0bjDzzuE+/EcMMosDCdx
Y7VRY9dx1eYg8NPu3PewCH2BwZRrHU7L6B/0VKmyueWfgSB+4tACwbt70/tz
8W1+gtb2GjLdNvA5sg/6s7HvSJLjb6+ipn4GmSDqZZXifPD8PyZT1e4EUdVU
667gwGTCUweaSaWbQFHoPItJvyqxtpT670+uI2SN3n9cQdp7PSJpTHzianxB
9oRuV2CpZ7LpHgZTh2RNJw/7+6xNxkOXopMaZBxCrHaR7lhB7qqUc8nIbc1x
cFLwvlAbhBsDMgjXy2XmkRnv9tT6FKPnvOukFR8+0z6Hz3qrlv5mtoiVpfqa
cmCZSQ+gCrNk8vdhixDZ0rgAvLZhP+k5YomQizRKxwC7iG5MzuCTNTedwJrL
VdE1XMdex9t1na5Ciiq34TD5cIChfJoJaNaJWKGGTiw0IB+Iwn+q1mN/XYxq
paqGrI30CVgsUKVosiujh4JpMZcpEyjTVjZfnLc91VvkT0HqE12iZybS4Je/
a6WgXHEZc9KsrBc+p7cU7iVhvSz0TpWicU6KTYeXk620AX/QPh1kOQMt1k+I
CQeKuzPo5oS5rtD3rgrOzKeg+MBu3VxZcBk8kz7+eluHSE/6PeB3Arc/L2wg
CZ6eew9SmqF4bgWxWHGsMYnC9O3slM0HWpc0ZgkkNTfz8sLOmkpKbD3XnsiV
kb34FzWT3qIC/VK+EDFsOzdanSDH46KV9o7koe8ENJykCPepbV1AHL1DmlFc
/fPQsykLLofxn3oMPMhgWzkcy3mtnQc4z8l0IgwfucN2nEe4DGNrQVuYjwku
bgbUmXNbffeWbHD2yYNtmB0nVykMc1j7+kJbaWlbB713yrG5C7Xk0hngtVl+
XCDP+TLi7Gsbd2AQZh+fp6NqmeoGBL9pr1/qwKkeX9rJFN9lNnPRU3q/qzPV
RLaEAAU3geRsac0jdaFw6/ZOAK6i7g2yXD8MtWMUJqNFfFjIhoL7xq9te9S0
aChQ6BKeyQSsYtVSXCSfbjc7+mRQ/o5QWVvXZKiDlo3fjU3mKxKw5rRSJaCP
E/pcs8KNfvgUyvTblehWxb9RejRhXoJQnEaohTYyB/RHLsBIfwGVQIYSsK6k
Uxiuwd7xk7PqpEDWRAmasNpAVFkqERGgJywzBPjHXtxNxPjMGtG90JWBl4YZ
fOb9DnTIMncXdW1zmN5eTfPdb0Cn5Dk+lknzQiC+a82LoOIA6NJmVqK7eSDi
pyzM39vJEGxNj93ic9+WhmKzXe6pWsc5VRbHJ2PFVlbhcwTd/++vyOImu/tF
r33Sw1jAgjGmmqKShbrGojp71xAjzrAbxZxtBYiHBDjvGuRgtneqHt1MMGnZ
e1U0XRIVZVIbgdQp1570t1cBiPlP29cwWCKT5I2dcWM43dibW6SEAvmtN0R1
IH0hriPRgTYIWlIbPHOBGLSB1z1NhgbR3TsOJt1DWK+DYsQmBZH0aqiR2bC/
l9HCdKGNnHFAoC2tVkVOAR4BeiDn+jutpi4gZVe3WW8kwkCbgDkPdTtEsj1b
cGq5GPF9tfUntHirBa6+A6052KXI8RYy/ZyF1wcAULHgEiMJTjY28TUe+82T
YEoeBMtubKxSkHuF7pT/kubETaxR0gKGBEZNAc4PZ+8ImXtb3OdWB7/x9odu
kgdv9OSK1G6LRouN3VAXU6bIJkUcg+58meDsozd8tvkoO+JmQCrMx0jHPVrh
b7wsFy7jBXa/N6Uf7RNIUZBu7RccXerAUibwufEeAqFZ1dnJiCy9C4PLXLaZ
Xha7iGF/xalfcniIKGO1gwlHgozCOS7A4/ls2BmosG3wF9YBHgqbccLEFNQC
ma0aSIsemgtKJ6DY+PLVeiMn3svIT5ydvWtSBphF8C9n68xQRk1Ok7nZvD4i
VlqNvHbGW4iX91D7b/Ek4ykMxYbpDVEh8of59DLk0aqbGkObuPezUtF8jfqv
Ji6/vhndWhDPW92n+9OdycnA7VqiIfOjuE6bSQajvCqZXPlI+Y3oKd2de0qv
4fLYDzDMTiMkI1LIEZp3Pjytt4amJdE+q+bUMcSgHE0lfmthj0cPqTUbMR55
QRspv7399GG2T/XLBjjwuFd7Ojgix5AcrZ3kR8vGE3GJisjcAbJl4Xp12jQA
ZbWtldNDqJ67L70S6jkhs3PCdfWmkO3mY3Uu7CcX5RnTv5bIG2ADJ98E3iHD
E/Uo1mHmDZo86HSzLEJgOmNlncF8WMCV64SzVTgZvqXCkFNKXqBJCYluaUPu
t68bCdHCNxyRkTb4EOOJhgotXi4LSXOW0p1vFnwzelLCXVYJdh5RzgzMQaj2
cxDqj/0LpAeWUU0cMWSxmX2cvYBW9KxntMfMnbzD5EAr8pdzccn1dHcIj8F/
L+qh5KVbS8QyFAy5jRHlVQ0InzNESlwyAtO8cSATgXNG/4ON89/+6om8mS0V
rAfr9oIrOvHlHVo2mjAhiJVoaAa2U8o6ubhOXnoLOpdmBvDyiT4utWtJIQo9
nJRkClPCHDrs7euDcH7yFb6DVvUHGmUPJ8hc8zzpw+14f/WcilvXS7+gvFrW
WLcQRv58iOyv+1mizePT9KRPnlHxw9lYk3R6PeJPUxnI3BRyLdz/kXZOoEsn
VpplvZqGtDaC8zwOx4LepvHZqT0lnCsYE850AOrXUo4IW/jGYjjMpAs/xLlb
H7ZkWlJWpkxpMIiOYQEeTApCn2+XiF6tEdqixR70g3/eqO1nmY8z4BqIb3Bg
6ppFpSdhk5njTJNVBvM+eXbN3MQ5n7Mxr2QHMh7SFrYykiJ0ruUlhKQcElde
V8sVJfmIgcdxfxPTFcxLW6Vh5I5i0ZryQ5vi8uuOZzSEocRkFVTDBi+Klvg7
8UtNXZ7vXFbWimfOtLoufslLiwRZ4S9ilRXTohrc8CaEqY3Cv+wd3YLd9Bkq
Tn2oUply9JjLdFrRuhS2GAtzpzwqEs0jpHB9B4tXG+faaO2QgDJWsW4aLatw
4TqoFjgZjKim/NNy1T6AszgRFYzFeaUkq6PQrwWWHfeoeyYvBBlEMIUj8jhq
vcoikrNfd1MZNkfcFvL9pjdeCxYPMdLKC2SLd1nXmmSDpga2MWjF2szG8Nzb
VXQ2dGmlKh7EQs5ZrbX22Og5My0p+Bmv2a1tjal+gWSCrrtUchWE2lYHqsJn
EQ5p68ar1THrvBH4meThbD7VIBxMftQyzTGo5OnoscJdPK5j5SzibVWWPDnZ
1Y+iqZT23k8IgLrM7PjR4dZ2MOxXfktpBUAvsSN6o1lf8eodkRQESfyOQSSu
wD3wvXA9/8nzKY6iHntItlMa0MwQEH1fsihBAlM46kNJ1YTwRlMAG7b4f3p/
a2I/mpwjIJR/dfByzf0+BhOhmZj+9WLFuwxK8OFDLQKwKdezg+51nxJL/j/B
Hlto8cKL8Sqv+G6btx0CPRlCzvTmjyW8x0CQ+CakBFPkMO1kF1KA+nJqY8YC
Dgm/j5x4lPb0/IaB8XAbqaRFWHRhWuTfJmL77u6fscUYunD5tsNw+kRI4bMU
6jYSubqdpgqS0Z8TgQwItDd8l38QrL3EkUyP3Kk8kl1gI9m/TshQDIyd9pOY
y/25+IXPhJ9Tyb8WMqqiN85M6Ox5sbQTZfyulJR1cablaGjtrg9ShE8yI0Q3
yLoWOwd0Pf06hoBCteyKEiQ0s7YyZxVY2mc2ag7MKH5ghuBtF10ogJgSjYsi
+LT61sPk/Q4T9R2aP0LYoAl8VcdFUMwZARWVH8nOaioHbad1UgM1K8xEFYoC
mNfusNPZwfUJJpDT+ClXgUHlQiu+Y0HL3Za1Q6YZd2/MCRYShq5S8yWIh9BX
yz+y7bMZ33W/DVBs0jjH7cOLY0e6cGrzWEwVS1taF7WTy7ROZWaQyCDtyU8o
BRRk3Hi8aZgLSIb7Njyn7sJRldq/EtSArw47lhTu3PVd70A9IrU1lIq9HOZf
8L6HmRi3uKzuAgFAuSm8xy3a469tzMGpiFY4BA0JaER/yFkIyj+15wENjFwV
Gt0kuuCXJzX1+ONgYq4xP7VCHjJ8ds+gANElcBvqgAb3GiPC/6G2tlaqGMmI
lI5TnHSQ+QCn3ZlVyeSlkuYKJRM9l4wJDRl75NnXmZnK90pRLFx6y7bIY5kr
ewAcviqKfL1m6BhoW0BjlI9rhrpHduwCnmnce7TouiElJH43FR+VtQboemtF
fIW1bSmMeRzxTwb5gCRUL6Oh8/NtUBSJ1WLs+UnIKz8c9WlIc8a9TR3eXspw
QEM+y+hUYIeE2SG4NfCj61MGMrRmDDqMx0x1mxilpHUzAJUIPEZZjArX0RPA
CTySVA/NrZWEaLJ4b7Pz4W06bR96WD2cwg0pxjfQJ89HLD39BY+U76gF93+t
jWguG4vb44AHFuPOyFHn+/Cfo3MJTo4wo6Tg7rLs1r2BnZ56ddr0TPNZkTj1
ZkErDVvbCTD1NUJUI3ksfK1ZpRZnDqKYrVEoxn/4NamPLkELtytY0gX8AX4A
dzV1YAdjzo5UA5gencylogHqIWy0fGzMn1yFGED17R7PZf3h1dlic0ib4YvR
nfKoBWrGpOMpAuSDMS+pN8FvqbgPQV4A+XuiPtJpzStAxZm+CTo4clscFC/N
Ly2VPHNSDPhkQ4ZiwLlUB1mTTVux8/Ko42UxGEWeOUFnk6QkppZEzs4OvGBb
tGfcqCEUG9rMXrApmySjE6PXtAwwCPIVQ0xqEKHb9BX+ROkl+dxQzOVJObo+
dHm5rk18UOYdrPnsbH7juLdco+uQQFnORSUDB1nLvmbJN92el1PeKiPyyYPN
TJlCf00Q5LthWP6k3gsvPaIG2a9u7eobccokBZLW2m/8EqQUOD77ckmWCTmS
6eK8Uiv8ZCjwf7ZoboYQw784YklSNqda8Uijqjcbsrm+C/OLp2cLYopBm1cW
I53QxNYxEpV7kP1mLciRyvB3H4A3XTWwNCwh4gR2AnTuce7781FeMU1pQFI5
Fc7S1YWvbC+/2EhcGamLAMe9Xi6JE4+m5uirniaICuzfQTURfoxlWTze6f0o
2ZjHIAkdMOAXY4Qm7dd+f3QXDPyTT4dYUaiSqcXj/fesrqb85NlXin40Vpbr
mUCzOCFoJHd9pBRVFwQOAxL6ixL4MHi8Xg8hWWI35NqIS+ngFb9/oStm4tys
3ebf6GFhoVYp93bqWJcqDsNOWIpgun7bvmgbsDyeG1Y6Eg7kqnRru+aUOW78
tu+LT0q0YmIrY17lCH0MmoPPG1rmy2fWqCt6tZeyEzursWuCDMUExhcgPpCg
Rp6HuDtsxIh4gpQPFlLreFY6scODsMnPcmtYz1M9vsNSpO+JipnnNzX3HIBr
sIYN+kxjlLbyc7Uc83Pk+h3UokaVc/Aziq2M7k8geT0iXvnxyfofOEwXHyDx
7qbjijrGKz7Pdgp2zIRXjxqv8C5TWh/0uxVNsSIhSfUnnRnJQUxop1cTZVvl
njDV0//484JwAGWu4xmiEYR7xf9Zk5hVEXC+r6FWP2ViaGU6obtE2DOxg1r6
Y/6n+uxsHvNRhqRyrDsMg+UBWSE5PA4DGujH46dvGq8J5mfCnANQbt3Rif4+
3mSWQgqXsGVUPgPSGEtGyiWS97Urw8AYAWodfrs1HGUeddIBbyV5Ull2CKxd
uZ9PCm1ldHaxeutgNsg97y95HxG0wmnvRh3yCpmhj/dmThkP8/+ySoLb3oMo
nm9hMmwwKQcW0SWTanC8j0JcZHkCbOYPn6CPR1/A+HP+0fGkZRqLYNt8bpGB
VZOLlV4VMJzxKmof+3w0o8XNbYHqIlqM605CxJXYYo/WK2ts+Cho/SZQzaSa
8PVRocDqnvTrtqwGdpQL4biohC1byQM4ma5vef0DUN67coKAjj5Yge9i3u7S
k72baXoJCQ4YADaAoYSx93cqoIZSvsAa9dlDyikVxHB+qX2ov2gAK0he37Jn
DeBwftKIJQETcgbR8B+J9CuV7Oq3vTcssr4Q0xjkZadyNV5DGg4Z8M0qvsZP
NGdKZfxoUqf/4yWsx7KV3/omJBtKcFGhbAokqOLQGV3vh5gnaO5zF6OHbozk
eENqCi6q0L2jFyAK3+7/9zIXi+0teqybVRmuQ6BITLrQ9QtXxA4kn6CURduk
p5o2usRDaDYEVTAbcEPdrgcKUVfImX3xm5GdvlIsHE9xiM/NaQcGaG46gYtu
5a4mkhzeE6ZdCtHz0vT03iRCHz4JIus/gziHYE6xHYBURH8+TPY7H/b4JROc
YQZBrRcQ/M9XHfmsrAyG4QMAILKP/Q0+jaMEr2rNyiD4KTw8rgu/aYd2EUbq
U4Na10xjy6dLLg8EVi89IDq4G3UeYp//8g8DgBrrLoRstJ7YA6/9IHz6zId8
NzQ2R+9c43uU3TqXfQIGNbPpvyhXVRtmKywXNHQGsdIOH2vYpM0nbwwyhtoW
I7Fb/UlRF8P7Ns09Xf6d+LtNhrwmmOVzG+bGz6oQ3oRjfNl/Sw/xaScwY8e5
0RPskHd+HQgenyehcgYxe4Ah231ZNfEXsjT4lXFg7J4sCPNGUfV7sCy7xy0E
lD91uwrWIYN3ZQlmWpwyrsvQSfWHrL/WCxFWpN7nty74wlAIUH9Dyk2r8sIz
tR+YEgYmAMNkttI1hEcarowAROigzxRcqSYN9GeVxFWWGICYNWozp9XgA/8S
XVXgKtC+qXYskZmT6mEKnxA1r9XbesXFOq2Azzr/9RfiLPzudKztFsxAqyFe
2QuPzYZuQ59Enj9blfsCSv1059GDmq75JtCun95OBi7aMphSf/NOla1iaUd8
XBZRPmDNlH8H9XVqEveJwm61tc+uV4Ec9TReXNHJA83g11Phas6v+ll5zGeo
lcXos0Vp16Lw3ICSdERC4fFaPtmQUBKsi/wyQEqf3VZpYiDvqKIXF9QGk14I
NcUtHlGCoF8hjDsM5tpzePXK1OV46G6kSPFo88vUplZXf9nDt/t6fIn9f/sA
rKZyRnhFL+v/nHFOf9vk+rXK1MjUCWsiMnM2fdiYTJE2bazK0pbeoulZjSJ3
7VNayiwWD37Na3jRyyhsTcpUsRGSBjNr9/BSDTEhTIiF2h04OguFqdVOSSzJ
r3cZFhErnkjiqkoc9mzjU8T+iXeA0gfX4vuk5gg3Wvb9R/oiYvzhpbqp0Hwf
M0llom2m7yXkPPYv4YrOvuspf8ZYIabaRg+XhX5gDeQz8Pl/r4KwxBK798rk
H4eQhPIfPj8FWucA2acXmj944HdKDpbrBvy+qIGzt9iBoIqLEU003K5TP6k2
tL4IXlEUDLOc0c2cNGcpwm2NXPeQqQwTM/FGRRxNKh0D/FzGzdVL6m7GOZwr
9xZ+7mh312ybnKaQWL6qLk7cUR1XBDsM9MbmoEKEkAhZlBM8tm5+5exGJrNC
MjaZHhyc/h7GOomFCiARmXfsBXiJKDrYHEIXBcSkinuQYWQuY7ta6P6/SmEF
ugvd1xX8d9TsCfOKfzjGdAKxeA6hp+2rLF/Fu1Qn8b9/Dsw23jLFTaq2VnQ4
bSb3JqzeJAxPBbpH2seDi4+o+QbXNfF1jwA14MLj2z1pPHlfqXxI6C8+hM8p
etqhfIgpcARMUla1T1T9FfkKttQraaKwRjnzQcq9ezbMztArNhMCzuJKBJyp
/leWcb68P3Q03XX3JteJU0RUCVL67i2IZ+1MvXAxEeAfOQsiGuwp/eXXnmxk
redtxsYLdgtKrJTNZWsHmC9icfTbtRMWnSP5zubwnTmhaqoJakLpEwUP9SXl
MA/IHrJcEpnSjFbP0jQvf7rAUiD4uPUUsMYQrbcH4lXk0nHurDL+CiKz7m+K
cKtLM8VOPmMCQC6EiW0WjaMDpxwKNQ1xnE/thLE83ceknD3oVsb1vSVfJdyA
0M9+PQ8ADv4E8Pa713l0IIp0KJD2qLFmoFLRzAhYFzlKmNUV4ZFoec7gceWI
ubTmUwRqttBnQISZ8J4X0aKztgx9f9hHa4IB/9/aNxMfl8HrqHhgpejukynh
vcdUELD8O0XpqVQzhNg7l60tDFEFWxy4odPLMR9MvoRYoGRPkD4AVjbBYlCH
uUE+fA3w0Z+Jb8thrpBasdKs/MpnFobhbAnDHyjLHZ08cWnPRNlX5zp4ImyA
uArhScF1NPl4su+gZ/YOrFBvO/w47LClEkzweHavqTHmTVyhSpmYGFSQ6BwS
5bqVLWVucroI6KRb1hf4gHP3PJuQe856DbhjJoYJQK1n9GiAPT++WDhW9aXt
a2Vj9ENJ16pCps16zaUKous9eB2WWcutVFx8htVg3pp7X+IvEiwsjnuDkjMr
rmpY3asvgIfrhym9HD+BNA/CbFwBjCrA04Yh0LkwNHOGsGFwVuACVq/++Gpv
tLxPoFwlFUhE5jmIB3LVi5rL1p36yMwlSc7pq6kWJllwUqMBcDm0ViaOKQaM
XSu+xT7ytahZnFPLvuDXmU5HSpUk5c23C7MScghChYZnx80WuRKm6oOXtVxM
yZ9yoRB3d66PLLGr5kwI+RUBXvf1aQ8eAKeIF4QUq4v28v5QNBy59Pdq+MgX
14MDEYfafHLuBUesw0fRbkGkpbFmi3aWRug7NX4c3roeEIYdvmm5WLmCIyN3
uEyOHEQUDCuO7feLxXAx0p6Udys6H+d+Wwm/m3okCefCRHtx7gZYo0Gp9kya
vdojV09/FY+HJhhx9Ucg3Px6HzyN5BHjJ8mNNMF7TXMYi5KbL8RM22nnJVvp
WlkGhoyxdcxzvf//6HaWRawYAL5x8Ldp7XTL4pL6QZe9THVS7FkHYoeBgPQZ
jni09oTr6e2R7qBMCJ5ZlJPYlSy000yjIHKCXk/tq7coZb+4j+9pEI0l+51F
cytfVeY7YXBybN74aeSAVM6Fz1CvkkfqmIwzsXsBDj7pkEP0HpKlncVuhNaJ
CL8j0L9NDqnvGBafYzUHxQwN2Qgo916EGhzjt+exBhIyQr15+CU3eVmhnFv8
kAvsYY9KOP7cyKcShz6jYVVQIny8pNJHe0cnI2lLM5n1SgYrprad0dQSuwd/
jtK4W4wvGfp8bWQXY/yUBaXNRn5xjVRL+2CeQYdm74GCzbb8FTGymOpNni6P
gmzOpFOnUCLz+tJ5kvzeps1ZS3pceg2TyadHFieZMXd9RsebbJBL103aWuxV
d5f6xZZs5m9fUhCrMr8zXD9TbmmQM7Ivj7cM4d7/GPj+adgFKRMHVJk3gbTm
SP4jyRKaedn+3LX9L0x2+DI/ZZ1u/bTxWzLMM7Aa46/zDfFteiFW/06afiEq
AEOoSqeP/baH0Iith+3g4Q9Cbl8HiDgrsKO8yNG7P9UU0s77lePbi7/xv0sw
bBb0xc2sorHFrmpmOr2BPifOH6DmOnS9OnsCBY+kqaWKMh6JQ8RXy/Gdk/Yg
nmeDXzPwOJDUGq8MLQ1/dD/zfNWwcDhpdV/ZOCcDqq4OKYB/+nN1CI5sxDGM
QAqBe+yFOCRDJGP0gtWeDbTCY6uv64EAG8DpRlb2NgJJtDBn1H8A5iy+76Ut
yzoN7SgJk3e2CrRJM2Myh7PSf5p+If5DuUeVvRNrzCM6d15Q/yYLhS0ktksQ
nWlcPpwQ6lojoQpe9a0FeC3CPOXZN0+LPXsue9ui7Vgy7rlH4bsFwyNl801+
ovAjQE58tAzfi1pE24naPF9QKugfl6yb6dC9JNfIbkqXYQ7C+6Re6hL1aNmb
Oz20I6GWIn9Ez3WXQs1i4NYtoW2AzZIyFNWLs8eS6s0+BvoPO7WlS5wFC4KM
YTcMYDNtYcm/Sb41UmaX8OHt/ALLh3uL4Y/nSoYdqpTJfHuKEra5xXooV5JX
oyoiHwcjV4YeHHjkF1oVYwWSsfVqr/4SdkOCWCmcuql3dgR1Q2tatjeuiB5f
rQ+5dJtc2f6thaDQRpDut+nMPostdtxxnVaPQISDhmTtyaB+UbUxGG5Bspt0
J+++vvRyKH/TMOaO/akRuNavDIQkR+JPnN3iw75bjp5h7kDhbS5impEZ508m
Gl+CDfDItax+yj4NI96K+yvpXr7axLMzWz1CcEBZUOqIiU2rG+fL/Zirmxqv
dEweKOWrXWUEy2N+qjcnQR9u3qG6z9RaL526qT7HAodGFe/kIltad8uXYdj5
Q4UtpxQs9fhtUunNuIkqAOeJDL4rKWhevrh+PqeCanULNndsD4p4UY4DEVpX
nr5MSX55COIpptRpbAjZ03PkDurA4jo/SDhC3cicPL0R9LlejTRMdE4vWHR9
WlRHD5u3AGgFskj/sImPiqWMN8hLsgni2rktXCXDkwzNwA0ZsHeAMZI5YBn7
pXwfsqZfC6QI4C0amAv+PYX2qAVC+2ltqtDwOM79MAnQHN3DJK7DOeeT+Zxo
Usz7eQc0JQ0/bY3nBLC6Udew/KE0TSub9E1TdrmMRAtNKsuz3WxOaYpkpceX
2z8IUcZQaf+vgCdq14jxh+kI5r7vJbuapYjmoGICDpMaTktYPbva6AW2QmLN
TM0quc3u7I6tjZU+bA/d7bTcaoG34f7nqBavEn7nZd5xN9aSTKdlohCdUkkn
2s87kOCir/KCVnNJM54Gt4/cIBpy/bTB0ZAPT9dT8aAhZ2YylPuYGl5OPZRS
EIVUJ7LcKEQO+ZQ7C6HyuadRMgFlbRuq3zhN4jbZsbQ8S6Ku5lpUnZQwWdw8
f2va3RRnlpX1kwLa56ovN59xjlSC7aBGwvQGeAi7zvPzwKVYcXDiuGu4msp2
vswVRhR4PYzizHQmJ35udE+bDkoCv0qxuOm1kvrtIsPqKPRSGUfI7HR503+4
CqWLFC4MeOnQPCxtJ05IA3iY1AT+W2R7YVb9nRstqG6Ky0qBgHbmNhJArR7b
Dnn4ddt0yN50cSFoTip8GpTVt+YLJiaz1XKc8sgZjlxyH5WSoHdA+34jAxqn
6QcIo6Re/EFlfUE1QqFAODTV3TDv39JlEC2GojRLcTlM3rAvn1MRCDNzVyzn
MrsgkILCfVX077sHp+a105g+jJLZ9HVHQHwBN2geV/AggZCX2onlI/mTvRFh
DhIimPGw7XYtBVafSSwMrOr3Qp7cmQSJEui4d94t7vLl7KCiXnLRQyUdDwRJ
fHo+eTL+tyi+3ur54G3HG1jvR+0EVyc0wYpuC8qITaTYPceeQwCdYqbHXRtG
dDb6m1ZnnThgMj0m8xyHpGUfjka1Q9vn829EZx9fzg8gMzXLCbJ0lwwY/yhK
fLl1/CdhJLJjGnpW9ClGs/5MSXl5UhZWfmexMTdLy4GMQ7dSNfNRezNQsuCc
AVEM1u8CIEcw/1Dm8GsIOIOGySMKXtzaCsuYKF8hpMK5eFp8phlNlkbrCndl
N3sNWkzo/WujfSO/w+3IJ2Zr82Y0cIutrCuDeRPoA1fphKOPf2wd5fnUUr4k
m4BZeDLNcXkpz3+49t/owocpOBW73hXASFjt9pltyMNhNTn4IpKWJ5JsCPJU
N4pdXIYZA6g65oh6VyjhEf69QETtOtVPtoT3j+v4IEyB4pHGUUrVjbgLzNfu
Bs95R6O0I25PptlwAh7AoSJw6PPNThhArniNviPf0q4rT85bq+8OzR5vTQ4v
mg22fwMYywFLOQ2xDsEADdxTr6AYJq+876fYK3SV51t4YgV6RBkQhDiMCF13
N8AQyf/f1HjIB+PA6I7ELoXRBgEitlKP2To57BXfinFpiEs/HPdl87Q1+5Ni
IDcekIxFgr6c9LfNpofUNvVE3wwC6XhSohuAAWHgF+cZn7qgn3difa60rBDY
ndIbPbyMAutsywUNS/mT6iyJ0ZYfj9VLSwMEfHgc8Twb05AROPO7EoaICgZV
tnKu73XBuDtvufxzTEs7BKZjSnAzeGEYjcI/pjr5Pv3XiIH1yoaOePHQ0iE/
KT9OsBWCmbPPo0Mfub5ShBQamu6ng6cfeluocx46bSsaDrXKlwgnPhTlrRVW
u/osku0qbHrGg70G0TgqBg7f5a6ypNVf5Rk89uNMXZwLhC80Nl6+yY3hM9No
9vjxYWkw3blSrSN4KWC71AaleKattFjnbgKkLKf9Vu8dXyRWc7TiTNNclugg
Is6VwF1z3ll1iiIdWthzt9O44zklB9uv7MlP2hTlqKVDCoP87mJ64kdCpFFd
+mQUbdj4cP2f3Xgrq969/MJKISUDRdJ96bzSOIdvC+kjpCfYhudSzr+vawgg
ASmy2cD+ZChNXbGS+POMYiOmxSC63sLBVaT1OHt0q8IK2lFe3ZFrPNGg+Obt
jRiuXFcfSShrmkEmKLPt6FYKNwffwphuQBRAujCr9RsCubpi8igSBePlCnga
zWjSedOsc3GUhpHS+gs4GjIXXXJGfo1HMwKCf8uWDvLidl4UOuD8gsNb64Xp
ElCzvJ9eHCUrX0xl2sQXzho+FKDtoUBKRiC9qkQgIyPDvg/K/hBWduwuIBWw
9rAw66VCJHbMNfJ+QWaIRUuHeEMFZBGTEC5olqyXP955c0e0K/7BwoDpzcdJ
ShLzg/YOWWWzgtXk405EyGBwrjI0B4G0km3uPDURrUGCS2LYeOEdXsBMriKb
9/gOe7DpWe4ZixTnLFGbfxTQ2SLrz63zVVIfMITefrSUzjZud/rRjGGAa1+o
kHDfJ4lkQSqYKqBOnsBdtNgbiRKKK/z42N7ZLxYBobXIEW2KsktvtqQGsWQT
+KQFRU2fgrNwZlSiVNuv600MzsAhYub0QYxUD/Jm+E/cE3ll9hvhV5UdJ2rb
t57pFW8W03/zwnK8jxgPFMfoJVdvu0W9L6z8nyaYRmZM4XGREssmovqjGOxJ
424v0WxQHp9IfjO1oJxrjl7q/qi3RGwO3lckvlxCVZXd7bHm40KYOqJzMxv5
v/bQwl9AX3SkJ4uanJR/D8XnN333qtES1f1pg2ntEvkjBXhHtzfjCmC46OQ0
35VXY5QapvolkAWFAcihzpXL/91sPLxL3zqIEkGuEsjhZZmRI2T4SfSPm1ZL
0q36TLljeZgXbmaoOqRuo7DuLBAqOm+KoAg/hdJ+NZCTlVw07059azvVU1iA
c+nRh6d1UHEPFSTJYxUKk27Glk9f7ZckaC746oAMdefkPTegrsZyU9hsQdW6
hFOxHkwLCzO7D9gCmlFO4oL8rfJhu4KFAVTvrX1zpX93fCqnbcxXdXLQx1VF
WUI+pgGKIprxwqO6BZWF932RWn7oGjDHGs3lBm8ZoqKjC30GDWtpmNEH2IoU
KwY+oYRG+qUuFQEw8upT3emvPrvxsSvD7jA7YFPjKL2cMQqXaDG4On9ctK4s
VxOdNYIOdKAZN2GmzAhfUq8ZbeqqCZKc/rwWga438PidvEUlfctcu3lMDkqu
KlIWq2DoDGB4FIir73E9Ng2mO+Om2wMIjX3cMtbAHjZ/JwDfg9k29jFiG3fl
C+38ZZ9/lYc7+X8KSXgRDoXEUT0zsg67NjXWOJdFpmeGehsprENnImW5B3A0
fPFUDSkY0Mp5DxSiiF+9EeLZau+fZ+Ei2EhtG6OL25Wo+crCziPhM/atLvkY
9o/qhjs/8N4NVYcrXyApOeT3j3kNNEkUouQMP2bjXxk97UmopHbSXlXUjWIg
kjdS4o550QhwuJsUTNhXeErAMHiVjnrnKgaYLKjrFLyZBcT3nU3nZvevcNhY
gYRQFjxdLoMCYSp0SK85RPc4O7plpwL5H/DbIUfS/DrdHafGiSuZRkeLHu7s
RqEMeb2dClgUG6IQ95YQnm6K4clDcMWx7rzNC41kuqXCtbXKJ8OK5zwoztBS
kBinlUHa8hhMeyoxzaw3ueGPeA4HiPAsOKekW69uFg5Kt4DB8TCbd4a/n2u5
TPXPnSe+h0tdLxOpRbBtY6JDzNgvMz8ftXu0i6WWGI8MZBdsJEvqvordPTZ0
bUY4Wp6E/rEHqg18olp/G7Tdscw+rgs9kS32Zap1NgaeC0uNuxEYVBw/MjB7
Pj2Ky1J8VD1feqVQA7MeOanHQHHFYA/KgSjDm4uKAMgMf981Eb7uqZ1x3lXo
O0cc31ePGF5HDvps4ybl/6tY0KEA801xjZGcOifOGdYC+IGFWYzxX0TQtbfN
Kqe0lsT0716ZudxW5JbDFewk2MunQ2mBmpZmkPvkjtN2hyTdjSp7/wXFn/bu
0OynQN0pp96KL80CvpWMkTnHYkzqX7ILVzwi/o0RNnOxhgDyvdLzeTqHY+1U
8c1Qn3tRiuCC2LhiFEj6yHKROHQqlXgaN8lXwcJ4REUJ+rVgupXEjb3/fYh8
lIHoZOYyxExgwDPJRP7tNDMTYhj69ORYxasKjZ5TdYUfTsoYCDtZT+6g5xPU
fEn9mkY43tthCkP090owP0qYXb4H4OWugdP77LzxCMYXmSuuYsToChQ58J3s
W3JHDBaGDrX0DRNF58CTywwZz3j82plq3nL+4NE2mdm1/jOSwOnpXPpj/aqv
D176NAMm6fz6tJUt0ksxBCPsYWHgayym77ioQ5Oz5r/RsqTEOu0/tKYSqzy+
xiPy2P7+1D5p0hvPtLU9mvVZ3vl/lyTBYGeNNMOMagZVHPrK74XUsjehtazz
0Feyqcl3FB6b38+hU+VZd/bLEB+D66AdJSyusysjqtqLrcOHHDzFjEK9Sq6A
bBOO8OcKpdC4j/F6M517nYZKBctzlpeZffzJZTDgXoXGUvrlvY3p8fyJ9oVx
0MUh6H2WsYBt5B4E22Ze1VQYK8esuzlf9cv29HUXzJTcOx0VstrZpK9GZUh7
OWYI0lfxVAbjix7QJTlAPtgYLu1eWp7sfIEYLKKqVzQbFnKzLL0yktVd3H+B
7oDVtvpv6LyvxkjJ7TtsX8Xw1IsnV+tzsOGY1P9DIUvfkNo3TambxKyAFaid
vAJKCctgVb2ReSV+hWP88RSF1+h+4+bGoUYoLnxdn8nUtQBkv/FTAwWuJ8rq
o3wlhLcTcVOUhEiogASTvAmMlXFKxJQqr0wM4LMIvjNWEPAV4/t8m6EQV8tK
WIQbFrMKJlNtJW4qYzPns5gy8gKcM3krdFFU4gxoEybfKhcR+UO06J2JDnTZ
i8gPJ9O42G1sv1IwvsBZBE8vtv8+Ru+zb8Z4ZMONkqAQMxdAzza/EGO5nswN
jTBi6GQixCMxE6M1sEohARwE5IRnPY3joDWBGxH2xYv2Lyh/0DNYs1VKyyzp
wY3DcgnTUzSv+KOJsGWf4pgJbYVqv46lt1oo9AwncScDjsQYySa0SSR6ukWX
MSSA0H1ZE0SW46LFxQqTVY2XeazBXEE9j3dljWem4aruUEOAd43wtrKwGTDN
aoIqxZuufXqDfjNKpVntnZ3EE8hgGmfRpJqS5OvKz264ujiqF+cmW5nHBD9G
r2FfAmme0urxM4Z5wuP8TxXLPHYpgtSj0/X3Z5iUIy+RUoJnhkfDl3imCYr1
kdrzJihvvFndiJklIIM0RqaJ/Mh+7cKlYcSwoAxMwQ/1V3tOh/D0a8xQZreZ
h6pN6Mn5ppoUSLBHKHEvEVyTtcgBo34DEoTi43TsIzAc66xF4qXlXg4Jeqz/
+sbz1Wsdzn+bcDIPxyMYC967Abr/EYQui0PSFFFCBRR5KnPIyso9PD7e1i53
qUZAoDdrcfvOA1L6Ki0eDc7Hx+a5CMPlMZWz3zrpcvQZwErcZBm4Vvp2Aske
rVHA5TMqKrKGHSr3yVFOjv4u21crve0b2lO1P+Ic2vDZhFbIwapYdlU0lmjW
p8bnnH9jtVe/UbyJTtKpdzks5AKlg6MPV0cXXLM1nFP8p67miold/D7dNXhr
1Q2AIaILMPEa2sCTXJFzpY9jAhMSdm6k3/wA1gSOrZj1+z3rfXcjJ2dOHDnB
WXaSilvZRxZP4JegEbDONET+BogK/aeXqu8mNLJd9TaG2P1N4NrvAOVfNsAP
tDLsI/92zJERr/aCwQ7ikx6TDwL8aZrk87RSmvssKLzqfoeFxuR68au1O97q
a7xeV7fTWCaGcLaCBJUoBFh5zbZfsUtaiptR1jWJFUnuO7ZgsJ1SSXiPA1O+
0nTAv0axZ7BuPegRMMsK1K/f71AqZBiaTHFnTprvbxMidFvvvdyqGO7mVNDd
7hxfyAQYkXki45MD/MRVulUX81dXARpZe69LIBDc7aVXNG8bsV068UmtdmyQ
axRVpXMA3IxzEZ3UaPDDzdHsieQEWPEuWr03AkcW1/Tci2jE/qI+wJS8iOyw
wcszGpHJgIaQ2t/BZIEnjhYegclkl47s09r3XnrWecXpBryO21O8zbUbGJ1V
6u6dqTBjmZYRgocZSgiVhlSLQ/WpyzHouZorZUxBQxVWNfmr6UrKgqj+rtq+
oecE38OmNog2lWOuweCQ5zu683IQUZdXwpuaENaGkBm8+ZL01OuS8t726DFY
zEuRadanERZXW5p56To+KdIaYK5fRvCSEfnj1RBq4onNvrFIU2KgrC3sFTMG
0Dzg/z54UR2iPOZcXtQw/xH8iMBrebq/lXZguYkP2SmiYA1n2mkaaQHrMsUj
9jxeUCmdZOU2OvnJDG8c6qxeOMhVlHOSretcUqmG0ZYYPmIVrrgZKAjZDvpz
3W2omrfM9/cPPaM3Id1zuMNmPRUUtfZZ1VVwHIrSm2jeLr2nZnR6OioKup0j
3igvQn+4xlPo4kkYcQtrkGhzd3+5ow49nf3NMZ/UOTdZjqnIPqb90F84GvHo
/wOlzh2g+v45/b/wJ5FGmzyetunRwm7afndA31Tro9HQsZC6siNbH/hD6zCJ
ADHnpptUFW8sN6YezZGrGFd9FV37GC00NV2XV3hqNMI08YYSpXUbWWjYnnGE
XdG6qshNt16W874RyxjbPqK05cUYxzPzhaMEU5/whfQGjISbgwoc8K1X9nUo
z5MhSUVPKlmnCLXEHCg2RXSNQgQXI65Rf58UD/jKrM2eDIsS4YYsvbS0WjiZ
Tr298pDv/hiIdSUTrBwz2pTO0Q3rcGLgUv05lnS97mJI28WRRMUxcBGdt9D9
+V4MqPbvLREFIxvQ3tN34smzZIzG43ugBpvfmn6kRmRTrAJ/HDcHMABPIfLZ
FgIaUJnwZIwJLPsesxIHlg9i2n8sJvclAmzuBrEhHkLxwo6YsGHTSggVv7Ym
Mij5imoK/iyTFwKC/je7PYfZHyUvsJyxx189ckabIvbNaLj1MVgSNhXu9Bik
oXMWNu6IJBaReAFJAqfrSCT9iWGnOyEJUuqdBNuSYLpX51/S8lcgCQEY1k0y
rIMC+9/NmxB3GWN60spfQ+QneoqStrSSdKE+/g+d+Z6iTzFdeowZyOtxqtGu
cXvJKkpu7VuE9ZwVoHRHuoEpMAxai2KXB+06xqSX7qBLiHmdbI88T4p/WKTo
4/1+otmJ3q2w9ToB7Iku/jqsNvTHz5nG8ZZsSy/Hs0bnV0x5WZU5VE0gq218
m4I5d1PB7DhckLiHeSdcGz8scSrT8PGMRVHuL9ewPY4sgsKsLPbCx5V6x1wg
NHWVYFBRhMPJsF4uP22dyKomsZLm071SCBtyW55Ew8LBtaZRP+bN0tNO84BA
65O3I3h59MAfqYOZbC6MlnyGTgJTrgl0yki45ZUoqha7JTufUXRQ9mQPgXpC
s1WuW4Z41Vpm4zYfSELnW62NCuX4yY7Y1f0qylPhmu6N35EKiVWQPFVxBNtz
KqCwAcPIkCsphXRhB+U8JwSL2opUwH4TJGGDoh176f8iFH5CLBRpxEw147By
VHDM1gVDwzRg60d0FpzDga4JkkkqiVGrDaMwd+sFF2X1SSHtWuwMZj+jAvsE
jpXs9c699lVhbGX+6tsAsmGhgeoEQHORQT5XeOTpPtkqKV4DY3TDanwyPBzk
ROaA0fyWo9bc1pRjefch5azcYxn1+LrEktu29NS+uLQ2D1BgPZH2AhReLdzn
Jpf/78X1lI0icpP8SjHHEG26oLUEu4HAiQpPew9Jwjg5vRvfrZblyuLKOylA
J87WdMWe2KpBN/gVCXPFXbPFi0++dCv0Sy55tJi/GsOl/i2qPq8o2brRhP2d
tEiWt+qdPhNIEJF6Dl5g9aq+vgUhQfoZJS+OcWct5M0fxjYbUPudiI0KTmf4
Zhgnr+rH2lIfwlPRA6dXuKDsoY8Kex1hAqAJ67miGlAcezQB3hD5GbrW7e62
k/Ethxmzvp4OV2hl5xr8kbmLH5blpQB+eWA+4qj5OWFDl0RM7997n3izKlMB
JKnf40DU3ROXuWGDKpWwhSiSDcyyWSuIPWWPoI8gpsfqNM/H+NmkJxvaQYWV
UJzb8FJEifYN7nSVeXPUplxQcTBY2wpZKxUyaxY5GcpN6lf/jMG2+n6Wajpy
MLivZyw7uCLLWifWbQ2V/xt9N90idmd/5kkMrahrDNSCH+nPsM05KuSpm0oT
E6uikHcTH0vuCn/HQZS0CMp6kcKWvB9nqF0pddJYOghzLHcU3WeiP+CuCDrg
ZYhJIBmvMQw4TdJdFKDb5aAeG/jqMa88Mqw4XTDef1RMRNMnDdRd8fZ1CXzI
G89nhPFFbJ/+1esLghM2PeQZSm448AByNjaC4aIubOybjG+lJEJsTrORrd2c
jcxTJmbxzYeWi8TCUfYdHaa2+Qkm0ZQ76fSbZz8OBgsI7VOrDHeJ+sWM/DtM
bErhe3WD7IhNmMy5ad7iQsbfaiQ36CJhEwDSdqUVUVOvI1icQ9Gdf62RunNo
jkvTaFyUcSFpARppWQBboblR4+ujos4UKdvCnDTq4uVWnilGl4eFK8XRCjH0
CP+9GbGKpdruszPyHfIM2JK5N2dRsBlRamVJadVX9aVCZMVnIHvI2ur8Od+r
LL/DAHegUY298OmkrG7agSdWR5fcZSAMA+osua98MmNPAoI03E6XNWmULP8Z
zW4jv8Evm+DgWx4cPEGnChf1jkCQKl1rpxPmbN7g5HeBXFv7eaVAgxRsmtw1
U+3gfGwJEPWIywYlRJkaQX7S5JcIUjftaKJ6WUuMi9Dxvh1wZJw4XIlYHpJI
iWYuDB+i91AANvSA5MmR3X8QavLYtSrq74W1DpMem+9S8ML6OHVmqOL1Dhd1
6F5t5aXaDFoz6kBidWa6pHpBLSa+mWMj9Bm1+pwyA46SzaCvlR7af2smcoN0
HjVwgp2e0KelFZlKWTpUhV5P3At341TXRrVug1EuqXL28q0jNPT3x485ZRMW
neV4jJAziQW3qtYikKqvqumz1NPYIONx/s0R0N5bAK5GCoI1bBDTsBeXgqeQ
Wy/DtOFfWxdMavulPlNh/XqXaiqvz9oUY6j3zxmB5pNh6/5w1TbDzBzgoHXL
q/9KPYv3mUlyLLbQzJrXOyqwSb4GYf4ObzYPwhrpsBNVIZaZruVkCTz7We5U
YJsboz9T+Ux6d6ouk96EgSo5bC/5BUd4gvbXLto1Csg1Qvbv+sgBGHV14CNw
kp0Rq1iJQyFAqdly+Zg0/frXXo9dc1dCk74VWpdMOCJHf5g3280RraJqunxu
sIynbBFNkQ374XFDA0hrrXouWPvfMXO+9Y34ZoC6F54/toxCQuEY/u7A0Lij
C0c/ye6kx4A7Vt3hxGBD42z8PqfH4K8Qsoin1icybwRe89WzwzwWPGoeA3zD
4yGE21r5g255Rs7BtbbvjPfss0MDpmOhLb36YOO7PxN3cZu9dFWE3E24FA66
od++5+cfkvTTCuJsWtVFeVJew3BB8O3BxdM07vBkhvIz6GTCIYzzKpF6LWUA
f0qpj1OWUm0WhUI9XD6SuiotGekEy3T2XnOD6iOs1USyYa3XaKopXpW9hvO3
JwGU+dxgP1jmpWBLBMIf9WmA0zD57u0gUW4vYgTRML+U+1E4LpgFtxgahTaq
z9SiUrtf7/hQ5fOwuOzaFkdzd6vL45J6fljhS+tv2MccXolZ/wsU8cpIoCIW
elzs8BvHxKWr6O4busCwsSWarPSJfQ1oCkJ7jGB5JUPmRn6YOXVcNtqz3RHQ
gIzfiuyKXvYbTtdumkVkcmDKmOqlR1l3RdoLSE/v8mn1UrNtn2WZ1vUVahmb
fR3HD2ma2nMuankobFfv3EgGocBf68Nd9Zf/nHmCY5UWNyq+/WyzsBTm8Hlu
rnHrBwrA5ZWhMQ67XSZRWEd0c/TTQTWN7WBV4I6vKTN71zhlJOPwIzURsliK
yDji9sb77EMCVcpwjK8RjvvA4yw7sKxVOYfifoNa85rtFsJsvcB3FyJ+Tmud
WUDtrAGD00ybHLLzO0cnpK1JbvDdkbCsSlxx194k1CLElXvimvso4UcidZTm
G+rtNdbgtITBArVGuZlhj+P8yAA1C+nw4d1f8DTV9LqNoyNmeyuUF1XAZkaR
4faBLGzzXpvIojYOMe+m6X2aDx0bP3pg3iXW+10kFQSTsuu4xKP/IFIoS02J
Yl34ynPk2SXSbOCzGQiEZB8NZ31xJqxCnBWBkHstS7kfsxWCsnWCfHF0AiTb
So6moC6krK1tSTxgvlMUdKv897+PFY+AYdlwGzrXirpSIUdNRM74NRB5b31F
U3ZCi3isVAENd76agxwR9v+cKphGOuoB225KQjHUxz62XaoBjVsy320qm5mX
+Zw+Qgv+KXJ/KgiOVEtig88L2oo6GyQkItBryopIYr/wstF8LFReh5NWTkID
cVTX+bVZPHPC6kH00Dj+jdJ0IBBVu3JDNPCJlRjHXRdvkCLVWzNBMHA/x4PR
OxfSYi9OYe4n0A0Nj1R1qPc84+5Vs5Fb0fMvW8l4OuN968Ag06HbX2kb6rHm
1dOOP246z1tgEsWlMjymzeb1OPcCOnrX2revDIeF2ES7LQOkllpl8f9OZlb6
mVZHtALVNXmXE5mLoqrDgwF1mGGJeczpdbW2t4cXFmU8SoTGf5dUkGUYsw0n
hFRJRaTahZ14je2Q7u+Y+W3mfBrDkw7BUzPMGmtASqxZlsWq55WlC2i06x3a
MkZy7TBbwrs5Fm9/ifh5cDTluWpE/vvNd5o6SvvT0is82YkDo82m3TZUbuZs
hOP39zWQ8D+YS3rL+lw2uBaObSDMLsEKKY+IKzMtr+lAl3g0LXL9LR7UNOfW
TvK7U900V15cvK7jNz6wM1YyttgqT8siIxVDvaS3Ip/bGxiTnhnOwMGzL/qD
ssXNWjFFDivyBTut5I4dRSaWBPl35PEkOuSuu30dec5zOh00AvbGlY+Idf+g
wERAUn6m1mUFPmUyCaHqy1XzlKq5cKvvkzFXB8LhDiSasmrmyS+90m5zVDMx
ovIhYKclAMuS0c9eomPd1TQJkiuvlJV/FycljL6Gj5sJo7e+GHDF+Vg7Xhas
GsmeZ/sfmaK/hvgscYMNb+Ks5NeDPLyBqqeTDkQODyOqn8hAGqVxns9BiakT
blzOoh5Bw84TvafXYDWrpNZF/eUK1pKHr7CE5DFR+DUQJWnnfm01M7W+ZyVa
GYsFg+8P8VIGYy7ITz4WIQS/4FuzIuv6uLvoSLzz8cf4s6CA56WdnfUDgDGc
PJ1L9Z0d7UyRzzJ7BT96tTqh0yK3ZgorGVUpnCP3VH+Xd324E3w/KifNNTZJ
UYkK711jDguAsXuEfebd2FloGZwiMnpFhCWIkZBjeWtLyHPplLHd0MWR23mq
hAkIQxqeplqum6mgkur9FKw8vQ6pF/rl1wR3r2Dwmk9vt8wSkY5YYk09Jcp1
LhLSKsmbpnaaWp83IDydOz7uPf+l6X+koF5mdiq6JxRFxbiXNROEApxIhrvj
IzJXat1BZdzNGasK4vwQUrFu/PhufeD1F9DDzKBwKKgaDWBtKFRK+Bxy2i7M
Cy/uzUK0DZ44VwRnKXLtPn/9En8Sw5YWvBdzRORBAcg+8+NnDBQf3J96kmTx
aZe7VncLRHsU6QY5bV/iv+tCtdJwypHEmvbtByLodKFMhonbuCXwqOtmOA6s
aotxSMHcL8OoXW3u/JGJsFSWXlFQfpuezl75w8s/JR2pw7KF9cFSNm2cqeH4
aXfsSIxE8vUbkYKSfZbdZmvAz+FlNd2Uvk1V6I1nhcDFGL+0mdWF+1xQfjyG
slrlB7LgMPX8IcLqocLU8segGlm10XhhJylYafwrT2R4uUuS5lN9jtQA4WAT
vQ1EjTXqWezkjQvVmoXdI5pSuTg7/ZgCJ8644YI3lfmVUb7V96QDHuW4Gm27
1dunC/2iiG2beDFMVS9o6qPxfdFa3pEPWncxhcYy3tPZEFvCi4H+kJAX9r9s
Z7SJgvYKq74vMtqm5edW+0L1kN/dan7hAaIDfu8Pk3kduL2Q9P81Pde1UVCB
zIZhg1MWkKeWphOWpZBHxg0d3MTSBl/fsw+dhLBvniPHotLaTcGNN+L/Ta9p
Ydlx7s/wUTYrFrTv6OpUPabligCkHoXad+9YwY/Us4Xr4ESeQ1m6Nzxa4TzC
HRcVOwgBpDwi3KJadXxra9yaLRjApW7/7PwfNZIhTOYKUwkxql9yvhETYUa7
X5o7dH3F9ioz01lRAcImXqx6GdceVJV534xJfDqrKmsPNmeUysgB4mUnrevC
wi4aEdiiEDIEH6DnIQtHMAHgDkKwFJ9NbA/HYZcVqT7PoYtAVKzQX9IxhdWD
h/12ciDcai39od3ZnURZD5JrSgcIID8SIoJFzoTDWf1jbfUqzJ4r92l+2MmN
i2QrHobvlazTLaCE9Ytfx56iK0lZGwqBT0TzTUgI6MJCRnJdsafSMoNVFmyR
n50yhZ1IaU/YY0sKzFZXbuZEkH+u5COCvABrV70NKWl3/Rm1eSQGlV0AauEg
sosL2i2Bt/woyViav62XOlH7iWSOXt1m3uwVA9UHSpamzL/ma2ZTDYOGyBEp
+hB+XSyUSEtdUT7+0s0Rt1muEHuzQTFYIEWJNXIn7vi5BRIhBFzHoMy1Hp6S
cGFrbnuRR4PdvjduHq5fRUbIMYduIA9Gvx3z0dNJ8RpAX1l6y4tW44clehKU
sevYvu0Q/4KhQA2nz13JaAxkwPOjpn+ls5+hcqfCKXeL2/iO9TGuMacYqWDN
+DoiV0qVNFTN7EjV/vAHqngEytZAwNK7675OajLKTD+S7zc+uwmuS9Kvf/vD
B0HFq8bbIUoBtuovxA2vLJtyrjvLu8/ls33Qgt92b6+aWigmsmYaoXaAofTd
BloREdxvUyOhPlgjR0hLi+Jj8WaSqvGXLvKm7PZh2FGCKMLuk61YFE9n/rd5
p1RGyr3raqCyXWtGZIYe77kEpoiKNNgBPyfv3BlrC9B9GwmMFz7VUPfDJR3Z
87nuJ0sia62+kwWcLSiB+ciVDg5jejyVw8g4hW9ChebButbRtfNsUq2Ylf6u
xALvEqqmkAuXxg/djjzfTpB3gvQWruSb4WaxbK1kt8m3k94HWS+wDWRJwlI/
pJ62q0jC+rc9I8JI5ifp9WyEu4idrq77Lpj+ibtg0uK8cfAwIRwlBr03Q1uc
ZUdXhsYuIhpI5995uH2f385v4mF3OZEBYsJoBCoYSwpJZmnE97zD2/yjp6Gl
QJ5raFLgFgnOMNWJMJRKI4vop8jJNAAgWmeCCHwcZG0tgLvOUuOuFGDdKCa9
x8peepwW83MDvfJuNhOA5K3fe5ETrwrg8MY/mzAv/bFYRbkBt0i2P7KAb6Sp
DnyVpyIUWLh1a+Vo55fny0qYJ2E3GGCNi8oKT2Ap2wf3PMgR6vNSEvUinM1m
TRMGc5NpRHBjgSwnhkKlFBsWVz13tiFM384NQ6sxgz9qQ7DLG0g4ikkX3lnU
RKtETmNm1kZ8y0v/25LIUANlEYXiiAt4RfSYSSPbdirShWrbGOgovvpttmUi
xlgsmsFQhwIYFuThx6GvN534J6F/bU5wA4MBW+SBUL4SW+Sk1pkTxio/N+SK
ZbXvnhyxEzyiIntVwcVoFdRqTRw32zxfAv3z9ZD/wZOCC+LbUM6EUpDBKm4S
aDCAViEPZXDRAqVebz4fftP2UDT+onC5jamS/7Jg6Tp9b+Fum2lya47MeFRw
NvyLn1uuZII9dMaootlc3KAA60z5TJoCzznjOb6kmXsYEe2OhxLEooHVxZ4q
+ZLSL7oPwu1WA+Ftzn73REQZnCTe4K1a8yikoitx5WSlGhOe5w0UC58smKZV
uRwsWhpdLcbjRU/qtc3qqLTnYPh9qgwSbxwfgRpIFtHW5l0xavPfCXjLeIlP
i/gqGXn2+rwlogeyTC0lLzcen0LDFdBrgT1zGeFAGspLseRC+niLPf9Et3WD
KP+sZ7WyIzgAFphm1z2sJ6aLVJ/NqErovWksryJ/wUwu3lzGhIaS/B5i0YLd
y5XSGL//Z03fHP3wK+RsKiqOlalHt92kgsZypLAr/tbCzArfwNzM0ASoR+QO
+oHZ+NpECo2278balPy/LMsP2qm0GbBXvCzNP5EmHN6us8L2aRom6aziU71e
CW5zjAjuXHG3TFjhINUEGx7dVf20isIOygwdQ/FVNuwoz/h1LpwEu24OFGBz
Mi0T3kUJdw1xjf1+QLG4ud38GUgI5fU4PahuGe0i9rNEXjKkDZRjM0zdcMu3
GwFEeqJhktTaYDt2M80q9T9QFQ5vK5YVW4SF0fsiJaGhi3DH2RtkBreXRyuy
DvcXvMQrZIJqzo4ZtEWVpuCykxOVkhgazSOKCAO7Kpnl+FbppNrEdpuF4V0Q
7f6jrL+z56xTNtnfqhq56XDzVXxgzNCwoOhxfv4jH74KtPlm7JagATDwAKtk
TLfXyOyEeD1bhXi29njGg/hTRCF0dVbRuOAdqS8NtxXKQGMoLkG8En6McsPf
WJz8vfOZh8ZaiT0Z2BbeR9ysGu0anppEz/qYLiia2kRsAc9r/CzdN6//sUsz
wONWBcyvInQFNe0k3aYoOsGQbY+lfszHU2LBS47CMWSdAj/QlOAEhsDAA8SE
wuqsmkTgCYPMpyOghrYjiwVblVU7UfW5FC3nGUngvDd+TfChUxLKNNH0Ih0K
FF6ffvHL7xsuOtkqJu7ZGe5d1P/LDfhejW3nluH45XKDx3/hkQLUTp8taegK
fpew8Uyk5hkDfgQqQLPQuCBLsEp1xpKqwTrhZ7qBsmThWhiJ5rA99vrzAKZC
zkEW8mXDDpnBCIVcWyne/V9ETrb5MtQpa1+04ZNKwyHMZUGzmrqqgNYd/QEJ
9yS+27aMQrm1JpAkVqWvv2gZfLNNpCZyWD8+o22i1EnAFPDQhfC/3BfYaKkd
0Rrr/e/co39ILNFXV5Roi/IlWB0UzG3U1gaAOZ6RsnL+tBl800EF30lxsYKk
nGckqiA1hbgKB0VaIOYrTf6n6i9cO8fk48zMKR3ysHnX9OcPd2KQfyx6eZK3
5GQJd6KKyEZ4DHKKIiNlvpan73qIjHlnqJdMk5Hlt5wGqAZNj6POs6S24wnO
SfJMJT9f4gn4Ocl8S5K7F938pFrobx8F/K+cBykdTlI46ndoBW6la1HMrcVL
AjmlGNOM1jhqDPJnju8AnAhp6kjDYqUrhaAGe9/hWkxmQeu4y3oEgbLOnueV
SzPDha3I8BPsImP0nxIaSeCv0uC7TuxxwUNJOw+i30AhxSQiI51gEy1a3Vgn
c9bu1AhCf/THYf7oI6uFyreUrqpePWeljR1MNRyn75HgsFCPonO06PLsE+C1
wj/xG28V31xKdjDZwhBcFAVHMriYCqbxRkPC470z4Yngy6zr1+k05ZSjs4jL
zhQStAFa8It8dgmSCZGIMpW4YcWeuz5SN0po3siecWkhOcnv6r+UyucOc0nQ
Dxm8ybPqQlWkoWbW/MOPdr1TfAU1n+QAhbILrwDLGDj0LhlNaFfNwV9w0/40
WDcG+rMOc2HuhbqosH3zQe7WP9ujzQzsGAlR+Bi4/vv/6MJ4MtCEmQM2ihYX
CnjFw/+NZMpRLhxJ/rhamyYBU/TlUqVdyKkO2q9sQipkaePdeGiBo7oXHLoF
ohr1nYYWqoOH/LDrM7toWnPxF9HChr0/frN5Ok2349KT3qz6JAAntO+oL7il
J4QD3K//JtBDjhqfxwNwUiquJEBJvq1ZD8vjbP0wqJ4Bl5ZZwZeucWqgqBy2
gISeyUrjs3Ka8BqWFgXy+X4sn3OHdE2mfayTBxDQQ2mJe4wGuLGSs7ey6iEZ
kzf01kEX9+yvP76hAeIkuX0pXRuDWgDaB++EXI4ERmr2wP4iruE0tsWxBAOz
b2ipm4w+GL3eqpzVqIHegeVLcFscgsKVWGKcZWqrkgbaGxXsnADEqnLC5tAu
6AV2AXxgGaGc/uGoQGZ0GMQdr0arQVGeuv4cXPHQa1m0nsoZciYDO9K7UcH/
Hi7Vq0xz3dgSU9Z7PP1a6sEkKV97SbG5RdFojUiFNMVBjSb4+sjOXWxicICc
ekDA2ZoXJSz3JUI4p0QH4lTgg0hqs01vP39ki087I1dRIBUJapHEoM2Vc72a
yHIMQ70aJLhgRlauS3tw1x8/B4gkeoe3V6P94bFxOR/jmHBse5yHv1J6waTg
72bRAKY03cOQu1gdA3CrGdA3E5IpQ1X4kT66YA9CMtdyuKlSuGpFQp2GXP0N
O+1tGR0XZhFtjf7lBahE0rv/1fBE2fbZRZIkEOL2+muudVC+DUxwLDIJrC0q
g0O6BtV7BaXqFCdvD8WoyPwYfP7u3pnL7ibBtFKIkV5Sc2EDUGNBBBBv2Fix
LE30/f4/Wcsm7JxSFFuhIIEdI8C0EUNP33AMlkz4wN43PRxGtHKC0TEIDBo2
nXEoGtFGEE8UXcgQ7ci4Tio1QGTQ0DQ5zUyOll9NPrlqT4l81iomegBtVBvL
XbLrXr0nexrNETiiZOV8qxQtJ3Xk0u4bCU6kwjh9o3wXKu3m+bZEBqbOq0ho
giZQ5Kh8NxQP2smp5QXxZXPa1AfA8/9DHV1XkAb7b+2MqRkoyFiqJSq1zoSx
SJ3jo5Al2lXSw9pm4IJ8xk+44SYecH3eds2u3M+Ak4nq7t585yksAvSoFw6W
nDUsKk65Rt8DMo42b7gBN8bGhE06bgBDSBM3TauSoJytBQX+aMCn3IlpI9/D
fjAkYll4MvYHflsIpBIcL5rq4VGCNPV+5CPX2hHAO4eJNT91ItpyTzFXReFF
x3dUaq+C8gOpVaSDCm/n8vw1pknl3xw1N5Fl7M7w4zPcqDasTq3TzruJRc0e
tNdN2Yf6bcncHbBZGEu7T3+bHcTGR54fcKQC6AyTwvsNiBGMJ3E82sTWBDpP
9Uc+zdZPAYWhgmABXf+d2bOU6iwJSwekzOTYS2b6hFWowgiJHPXE9f0U5yaU
hWtJOsbRffHBuHoXBlg/jM4S3yx2WKKswTV4eEAJ3QBPn3huy1W7RCoukydt
zZvSbBtvAr1Wfk9i6PO51z2B87q/LmW1bOYYFZ3jb45gIJ38MMdDpj5F93wJ
gKGlkQ2g4Z3VsfuOetebkcYbekW7AsUy6FQXWRXcKXO++D8e5kyttxOh12oQ
lY8dlnjnd7200aEoDOa42FFN8T77/YaWRcQgM7Hyhjiy0qafeZIrNbBl6GuD
UAZp+tKAPDh/CXmLUaKy7Iqa/qONMedraPo1D6Gm5roZJvZaHm2HYj/0X4RD
F5yCr+gtCxbTyAfVXvQFVkklUznXFFjItq1nJObJj5P4Wkj8jRUNZsp8hVb4
O6SsPfvnaYYVs+OY6oRZgU4udjLpx1KcUzqhBSlJzOs6KsvK9z5+2d8t5lvM
96j0+Ojkcmy4AosefADbO54y503/3usQ/Thaj/+HQVkHRJfyv3M0DJvwS3qJ
vMVoO0KGZFcc8Sg9SjBoulHs2JPt6d8uob+mmHlQV6zLwW6sLXdQqv6hOSaH
IKdnLyNs1HM0tUfVqzEk8t3vlbnBDQIUshaBe/iJLeWQ0d1CUOgeV/MTf2Oj
g4cbGmfX1r6eTPsgKhV2rNbKwiidN/IYYQaWng/YzQOBl7CLmoSNjolu91PJ
3ospSP++4Cdbtfr+k0OGtvGTMlbSRGIcuBZNVQn32IM3IGdLaZ1MKTFTTdKp
9DGPLZYiJwLSguZf52xa9lygfce34Zi7NirCTtocriJLIEFW/ZFlySQMah/X
BQvoWRXiwwjrBKVQXJJjJTaGD6cBzlOV0A0kqETO4kUZ8TXHnkdp9hGGJYpx
/W8C0XGHZrr2gN1wxuop/wT/n6ihrtGHuOkuKV61uD/I3oU9PNiHiEvBPVPB
4FWGBYC2pQrgnqsYEWE0hw6xM4uzGcwzCTVYJFSuWhY3tR09Y9NtUfQKstHZ
BQN8eGe+4DOxph8byYG/MQtE+2RlBNi+zjjKUkbwDUHdPjTM+9GYI3PmBOyp
VZ8SgiK6mOJoT6+MAnn5Qly6pyO4J7TcmLhEqg/qCX/GKC8ZiDYOm8G6Etbq
wqQscTu2vaJAcESBWmFXjLMc3Tn/4cIvf5fICrtkTUSSNDKhH4GMh7m+p5sG
8JpbZlnMT4DSeZR09sC2gZImiK+qR0DgP/JUzo1LS4BSdQZkREa+U48Ti5Rb
+/CYeTL/xElCAXv7po2eeavim2Xn4qVHLJq3w0eue6qW4IjuXzFyr2RcFkMg
1364GM4RhkTz4bRt4zgx7kStiLRXwu+xMdmZ1/Y+zyxeze26Y0ROxXglDGzM
TRxoX3xWo8eEMO9NT5R6OSjbKxy7FI6cqRQycuxBA4EFIRQN9ySBRIS7pV5g
4HUurkJzt0Z55h7/+Hv3W7OOkgoT0xhQ5S2Ad33amjQsLCZ8wshG9/W05geb
LxByp5JSK/AmRj0HHrWwZPLmZdGeC9oFq+44KqKHwg49mAtb0b2atkkJ1KmJ
qkgQje2YFj8Tgxhlz2fQgdzWuKSi6+rEiMxaGiW7URFYgb5uzUFv109UKgM4
OTOGARyES7M3yy1EDeG1DZqRYLNNT/U4KcGqfp3SLAPm99qvT7b0/GhAwfNa
GuWgI307DzGvYfHKxSa8csnBKUpxIKLHJE9XnmNVXzUCIpLloCXBWSLm/FdD
8A0L7FpCNE5wzJUbCbz+mU5Ov32GTs0hlwOE05dm6YSbmNmlRHcrShR1gtgP
OYL5uT54l4ug1C6hRQcYHoQobpQQD2ybvyyuLaO8644CVOEMjEO4SWAmMHlK
FMHNl2/mbUHnKFlCQvmgKlcgwdugwNyr6Nedxb8nLU1ve0aetSr42fU22Se8
8gmWOGyiGFz2NwJnb6ok6SbiNt+AR4NYcdONHxlTvW6Cr736EnCMaGb9zI53
T7tz1RQuOppZTx+omH7ryU7UfohGnfGuqbRHKI2Xs20psvIrTrLFNDWdekH4
s0KWtsMWPY7/iOtzmxVVTLUTRXRDsHIST4Y+zK4JwKAdNVSZ+/L+l3rqvsj7
I/+XZpNBL/MNS9ZTZJR502X02l5QIm6V+yrTAhWue/wisP7bqsJaoE9Cfq1x
KiiJylmg2KndQIZ5hkwzy5ii2s5uH6rGQzjuwMFL+Xm1tYIVe1VLMNEZ8p1J
JMqXcVV0NwW/EadOhg6/4SH2hMgLmWt5NVGdbS+ef77/eUrhsF7VJN2O00rD
ofUIozpVepuTWSNhC+jBCYd7ags4um/N1UQdm8G0WA3mDhHTrenzJAAKSW8d
N1UUn02HBfMv/Pxe0mOGnGcSlY8GUeG+Dt73kbpj04NcLcbOW001Bo4RiCfO
SMuUdyfe5M4lD46VvWQ8kZiFH2kNCD/40bHo+kKFQFZa9ZaV4hkceM0BCgGg
q/lQ6iLhOJW4icP94XQY+AuT2HO3+f9A5tlkf6zNaJ0ncsq2Cv24IuWRqKO/
E5JD0YCJlQcaSIV/LHQ4rzMIuT1iEgk50pvgiyUeeZTpbd5rlChxXbm9QbOT
KsvvHQOYFg1+ZrwSukm86QTk1BZAXOxevriwotmMMqp855U9HGebAg96ZHlf
OGHrrvYdu5iYtS1pCOvPalij6JorE7has59ElqaLDcIgvlIHOTG1ejXaAu4L
5rnarE2TdECtZU9bwwnoZp7RHIpKlDHLifL2J+3HZzeIcySS19B3LPHwPefj
Ik5X6KRnwtODO5W1IDwTBG40r7QpAQxnaPeqdCkd3TemwMmpdRs7zNO0JECf
29bxBuxbVdSxz259Q4eDbGe/oXR91ONI0c1XTKli3Sy6iwz4eYH51pYswEbP
X78qzZKMEPmnC9r/MUnMcI/US9ENnARlSkDUKCEzju/IPA9L8s9jw87Unflq
2vgune239akKBjnfmflWG85SJKI4fx3e1ug4LJREFvhB//OjbeiAJVzE3HE+
ajCgFQxljEkQyW75OMcx6XFu1TGMv7x/nt0Z1OfBUBiO+fyZOHVgjhOW3DNn
CFzMS1my/3RQJc5PFNKNukc/t864JWN4MmQAOQ43C9k/DgyCxVCZcI0hRuhh
Ud9FpYxDr1U8S/PUa8hfvTSyZMnytOKygBPOprfnmbZ1Pz079XYVB9ST/EQG
EKFEMqgOpqKBgT8355N3c73pprkBX7lV68u5Vb8xDYnkT6A3pEWIGi0Ten/Z
0qvqEivaLswl65u0mfTrk+9cWICaKuC5puRi/OnlXJRqpWxZJstA6FWCV81W
I5X027yyWzvXiAO5q7j8FOwNIcThbuJbivUiXeqnK8KpAIHW0/JVaRwtVNXI
AhYaaZMN9goJMPwVuJXx/hdq5UXW188G5soyYeSXLo4vpsEQkHsiDlLDnu2Q
3Jomne7JtVEPvpbroOXBKYVxHbNO1LokDq8qA3FqPtS6mtFBm7K39/Ru/s4e
eMPU/20vY8GdkIRelxOWR2D9gy538coZdAkKJcihvb6P3eUt6VX32eOKy2X1
qi2FN8l8/3x8HEz2xEDYnBzuGDZ6P1pvgUY/KQuD+bZjPNEWGi17jKZFkQ11
2lAuDuM+3o8bizn/DCSE6nWkg+XZDdC+amLFd8msE2YV5rIS8ticmOL/1Y/7
hrsozbIUUMcjqti8DLbxRgz/AuPCvmLjH56Kj8vZtF2+CkH2fLmyL1LS332I
FM5bp/mAyS1+JVi79JLS3kafJyi2LeuO+TMI87/nKuKgRKiDNaBBNO8AAZIa
SQRjFJ2qe81XKROlgibel12e3fC2Nct3hrzswSje398m4aTYEmbeA+HzYRfx
G+xKFXLlRP+g6q+jHnr76PjQdKY06y5+5/wnQUCdRYOQlIC6lWe7kpXusuhl
mocVZUdTFVdhyBp9a02J5Wmq3hM5iJVkv3UhJgFW5B4ccTr4KghJ2yVwRR1x
cKLNL0eLU4mD10eOmVk9e1ZIinz8TZ8dIEUkGzAoWBeV72+Qumj3BnwO2Ucf
3K/rWR4LKBXl++0JS0EkoTsN7fE+5KoITHyf6+bypk6BiUwAlTZUrCeVtzpi
DTZHHIGg5F335MSnTtolrLerTYZA0gc/h+ZlmAzz1D9GvD62eJMFLSqvLcP5
ouZhbjQrdZAv/83YyOdqczc208ZiygS+qVx68t811kty/M+5PecYSsOG4w3r
U4N/cLdUfSuK/K2BmqCLh9Uxb+jLCUSU9C4IHmdc4/+p+tbAyXN+pANCyvnR
lLK9rpkqNX09q2qbuLF/CT/vD/OaLr4UzGyjV26AVOMhu55kyCp/MFaDJUen
dia16E6rhmlzesX4UZolGbGyqnxQ/sgxd0/hItPmG7D8bdr2J70e3dwxND2f
oOcb97y8ehiuR1bBt5Veufb7h81XsW/qqh1Q9WbJyfSCADepsFWyBKHJPrZl
Uy1yh3Q/R7svlUogPCODa0yGt9E0XPf4HnhQRRQkts9CJ0E8kSnxJIyLkUDW
0PwYMhOIsBmGC5bNs78CLAMra/N0tgogtzCmE8TfwTr1W8jNRm2pI39528oI
lxFPJgfj0X8+rGTYz1jzKMpLSrmu7WGXseQlA/f/gGeqxIBbphnW9GfBy9IB
HpQNmiYSHjCiOugflFDAsvUwRzBnpy0qBiGWs+qsIiUrkNxCI4DsMN2HYdnA
OldQAprP/bHplP4EYRppzTMZCQbU2diEQb8VwC3tOr1O69AsHQsvp2VzFz9I
JLgGL0ZkcxuGpMc1qg5tP2B8wN7lR0UJffcSlyFTjjLPW8qEql9g4IaE+DQn
tmNzXJRGQTMQGbjijqplVq6MvS4tWM54rZ5MF3QPbynH0xIFuDDmcVg1H9do
4v7U/ZyoeehaUYKcblGys9uL5mrUtLFkSWXiZG2C7MtToeCZ/k1VO1vcoLvf
2a/kwRQsIhYtQHxhIp2uov7OKInFzaR5q6dLnbrWsiRSHCjexNvUty+shTF4
qRfzO7+V6zSD1IZNXYbqydDDO2nd+eAvFMZWDAjqeZwlQN5ORHKlYJCqRqog
9eN95WwdNJw5mfZMA/6ZSipBR7v9YDtyforY9WgxXFv1CdMOTT3IZANF04Sw
QnYXMLmN5965F/XkHBucjep2zsAjYEKQAfUXBHc8ht39NvC28m1TMSGOo1mL
XYh9FPOBLeiu0X2kbDi+Rf8eaFrESErJTr1BRVaEEgStKN7toRM7brslR3AT
cgpboQZzkPo3+fQKVGGi93o7tfHbj/VlB8fVXhR0C5fpXa2B4i/UhwamevBN
/pHgzXMQfqdjcApBOyfR4yrEZ4fRULfx1TT/atxsS5bQGT19WBgZ5DiPhMTh
s0IDIdWXf12F1iLQ1qgyDejjQ9qeQoeBMLb9sxAVYbYzbRVFOFmTEJACwvU8
hCK+xUH4zEEISQ9rY7mFchvV8dkgZ9Fw62FuDFPVwKRdTBbAt27r+UugzmEh
te8tsreSgs5SR9Cx7YfImtXHJCJZSLtYJV9xaaiUmIZ+UNun81iJwwpYgwnr
gkOhIfSsqp7Bt59AIO+lGSQrW1elbtNRoC1Rf41f29nUVBqF02kvAz5eUMb7
D3V7NdBwuZG4VYnTLfxHNIfazR382LkC7OJiutpDnom5ZMOjeDdzr4pnyS/M
oF7FETJZzxbIB6oaa9eSOPqOuC6uemuE1aHgQhxL1aTs4zMRyPHHSuEP0579
b2Qhbzg2pF1Os5JKV/4gmRFY3HInXjo+kai0phTMNx/5EUzmz/j+py0JwI5W
j8hV11E6nB0uZ02M2pkhs0JpOgh0HmJTTu/m5jBRkENiSjRALij5qioeOUHJ
o5g7MXy9pQSdTWS1WQJsE3aRPYtu2u4zjwetfZvTl8MzXfOWMNZsJeRgIbaf
NcMb9PoJgCmyDkOOI/wkHaOFlNjxIVzyObyIZoiWUbV449KPb24cvNISkA64
nS4ewGWeHyE44bua7Y+5+2QOtMx/3V58ys3U2Wk77rZYYzo4Myqo3fbLqH+P
jYP1PMrbm3Tl9rCqh89q5WYBAJJakTdf0I6sITYuXJ4Yk0GUXr/4FAr6ULmf
lRjuE5o51D2RUiTQB8yiJGu4NkBNO5HVvE2vMZzwXav7ulPLZdQwIIPtU9Mv
E9mcxGQhdm+5jQiaflajWYyaYsEqPx8hN3KiKkvw0hEmFH0VNbjRJnOMqA3q
3EyvW9oY/dLF8wdTG52jNewSeGPEdExnjb2gqjNSAme3cGKB5EBEFYH526cj
+tRftoYt8HE46oQ+PVSMi7ccA7zwJ1kgqKlJ4r7hevj/Hfc3f6EoclG3I9sK
fmObR7qxnsTZnQ7EhsImb4ay+9F1H470pGzyJNmRL4aqOlMPp4xXQhJdv6rY
TS6J8ks0aNpEI1VQ0igHxwaFITaayVqi2ws3rDteHva9XZnj23sKZ3WGqKN1
tgz69HQFmrroN31422Ba3qCupKaZeyRu3Lem8ltOglYXR/50hKqz4JyBVbus
2GrmWLZ5rUEOJZh/BfL9LKn2zobGaq11ywszSCEYtCcC8aW0JgQCnMqgctLH
VFAILtpxBnzSEBJVYD1rvLeRhCUH+vMJ1bl3y+LdkHEDogy/zCyY93jZItex
kyRUx2HTnwhn+IHShTfFHrBqtAuw+3EPl3xIKOb8w/bCh66WsuRw6U1O9UDq
CUKRTl8NPUCq+hzzwEhi5el6sbj1gIHAp5M+XR8jlMkxLyWf4/bpOiHWldzi
u7gAXlcjJ6KB3m+7LsirN+7VkyRtBCtwvmVROo216DKSCVjjPbg1Fz0nagdd
znFxnf8wmByHidPqTrnlFG+cMNTIQa/N9YQ5itSlopsXSTGjvHBEJ/FNWgW9
KWiZ7QbZSI5OnRGNzTVN0qHurCKXZaIS/lkfoBRE9SojHSB4hLFpRMQxLfcj
owtloT9/8a8JkfLOtGbN2SNW24OK1hvKj8D1ZVRf2sctrwGAoYnhC77k9UlR
RB6AF75fTH4+p+eNGPTf1+tNqjwvgLsbMQ+WbrUKZzYPAKVaBPuLynrRFc/D
dkXxZoyQrbbuHi4/GDLHsb0DgittQ+xb7ISXD9FqDWO44xeMlz/LLM+B299s
XkI2mGqJqRzwIGmggGRl8M2vpmzvjUw6piraVxcjPLdczxxPxYP6C8RC/MqR
WJOKUQKHNRnDmaPrrpapGKoKLLrKcVRIV0mb8uBL3ecCRroObHSLSChIZsOs
cOZqbttpyPYfKe8Z7mfiCJHjNDwzhoaCpZnDqaz73h1yEgr+xAF4/jnVo4kW
CdnLZPQF8PfCJMnGG2EFvP0LydcPxT97jhkeS7+Ocj3GymvbXPBMH6oM3ltB
PR7AYuM0/Zfghrqjmmy+6rU5H4kdMGUGuhw1o6YqlyDe/02cbHBSJpBldGSN
9ruBORgjYsKXpXyhtH3ZLzi1C1cOX1rJ6kaHlD8CJqGaHS5jpmP4HeWeRi3j
VTr5vzKjRXfE+5IrLUwKTbeO0Ia7qEpRcbFFiI/qG/pBc0yskUS1m2CsGFtW
/h0gCiZdb+QIZEny7V3bx8O88e8fBWHuQrK8Rk/ko5gH0Vh2mj2s+93NxPA1
q9IuI7bkPtXciPfW0s0FsiVOTKGjRjSRLEI96nOIr+GGig3NNqCHJnb6fQ5l
D1nj1Oaj919M/wk+4NUD/4KL0tRajxFK6xfFJ/vFVFLwo6XhTq85hZObKANP
6buC93wXoYw9GOn+/zRQ4/JF+xlEN+EWMOiZZqz+4lmeEZMGjfKZ37hhFupQ
hqluRSDqjLcP8gKWcwO2Fm+zfqv6OebbdGcDd46dALMu99xMe4kN0QzLAqBp
4z/8z5eZu5f9GNOWFnb5cYTBgInE4PA7duLdYPxyrbgn+qlulgtZmwJbHZ+o
sNT4832eNjTbyp+TFZ7GTysQPnc8mfObZMK+MldQup/Y5bjtK9J/SlFhqMNr
NfzBUah+MyfZq7PdVYR9GXXR8itfRt/1xEx+TOZkwfovm2nGNHU2am49rjyT
uws5kfyJfdmHe3oxbtBoPDNnVp+QaqMzXOwLAoWbCq5sPt6JfEXsiF52QCSc
Rc3n/Pjp6iNwdy9Cxlzhh8VvUmt89Q5/5cT3a4Fn5o430e+hei2uC/DfQYYW
NjbSuN1nlysImwWIHtKQf2X3L+WVZXNQxZ5WAA3Czw14PYhPRuSp3Ax69Fa5
gN1Tkz724ZUbXnIGVhlAj7PhvLLUUipKL7j/jmRNx8wn5ABTxD1d8br1GUx8
7mpnRlMv76rjI8tIkZa/7TsKGWrzi28Di2qqqPwAVEsEJjmQm2cSdyQwBwrj
TAWNP/ksNov5MwwEexArTFIj9Sl0txyN+tYXR2OIxq+bYAd7+FTGRkLcqjFa
M8R8fkQtDupyOWM0gM1yn9NSebO5fVTWqfoDOkkD6uPX8HgFDFBQzoc4MyJK
jcRjgWqqBnfFwlol6f+uznu6oILsXHkBXQSRTMIXfCjxFaXkxBtioV8tczCx
FWr2kQovLYnvWu+5G/6VBv9WdKCbAX9WXlmVuhcbfDkLRgiLpLUdCeB+iLQe
fXvj+yNsKgEdJ1JFL3VzIQN3PuqOG73dyqL+nLcWVHZqnQvCoJzjmmrxGqpj
jhpaB/uxW3Et1TLXw56PwU0ecV1yGqxXqyYoSn+FFGTqeM+hKi3fW3YWkSIw
Eofe7kM5cMp3BCDBfAG3UwTDhms6jnjpIYp1AgC8gHqRSBA1OSMWIgnUcHq6
4Ur5Z1xRBE+okXfBmANZCrl6hn0OVa8jjeLLP4gnVMFb/t1E0/tKnH7Cwuqn
i+hMIEWkk8BFB6IWdh4KiBw++ZMjaxGX4tR+vlNW53AIKUgvExcfLH6GNa1W
AreXF3Lub3E50WUY98TmVRtekQNURI68iV0zZtKTQIV16M7o3ZtnjSa0GUEZ
1fOw99dpC99lsEZ8htqUjwJYedFRfNyH/cQl0caVva6xAfpkZ6FISr2lgfMY
qxU96+H5OQoRRK3Uts/nZJTs54Mt6qbOo8Fl5owIkpWZMnQMB8//nz4cBrcJ
SJBX9E5nhDaGFc4GSjWePysrnwgv4N+J2RnMFAzpi6WVqVh3oPHluTuba7+r
0/C83eKYXbdCHjkqDRf5DbQ128irGZffojiUwQz64fAp8nY0ysINiGmnJg0Q
j83kjLdP399iZwguqkoEHwiRzSA6Y4ZJEVDc5pL52dT1iQnjU2uBSHNYuwlT
/kwzNfwhZM2P7DYK0/jjH2aYcFYO2Lf37Wv3TqxiXwn8N4PNSHBnpA7S7ApR
YpHpZTWlJLO2g+hvtLm5WuQSsHo/nPUrnmKws+NlR1lOw1iMUv/Z4X4tBo6A
nRvISH4FeBQ9uSQzdQ/eWVY8bsrM/glZZs4d+1z4QXSIPJirDp6RWjsE991h
UxpeFR9v0E9tsPTEInpHIUFahYS4Pax2CUsOZc6GfLvjN34CO7oz/f0P8a7S
ih9ld8QJSe5xHC3IvWxpSUx7+yvNo+pBSg48lQuamUxLokHMP3DjgbhLCiZ6
fvgOJgE9ZtjTuKAMVZJMfDcxW+HppBl432rbDnVOw166SdsPRpkDSYGQSgnk
lgWpb78E6a2VNp5Pk8E7X2xMSE84XDzkaOn7liLjnrS1SFfrtPCoV4CzhfQf
pptPSREAyTuJ6pG9w8HT7vqguSZByk7zg6go1I5ZoofvjiEgRoi++iKlMuns
cwTxfKtT+rifQcPJCachLFLLNh1cI3crw1s/Dct/+H7DZXjYuta0CaoeK+rV
MvfftZhrp5bPsVYoeb31Cz5GkfnvVOwtKuRefXC/1pViYJQYb/iDK6Q1PbA7
Y1OX3bs8SOh7I+psjhYSEbhVLqSHRZGlFIid/vxMTRtE08pUHyi0kg7nXBcN
poJnZubGY6lcbuiQG61gHZ61G+3X9WelW7tB9TxQgy1qB7r56gULU2t6ysGJ
x7n6WULjr+tsvWauVDe1ZW61pjRpcRfxKV9uIz/tS/LmV/LlThqfh8ODiT4k
4eAC2uX/TkPwQuKj7pDwZ6qeLqw8wF4fr+8FMfLwL/5EE56/MN42Kb4lvpQ0
qcxyVX8o2aw+y5RPut5Y1rQ1isiNlZeETm05ZOyVqOrRyXOdn10oOLkkTA8I
kX2IJB4UU/MP6nQAhc7RorU6CCrKIEQ40DGoFlcWioblAOtObc4P50AeDJzG
sCsFCVGtbfqP+AQv/iWpwAyGY1pM+wN9/utmCHtfppcA1KKlBnSs3CQcVQqP
KkT03sKYsWQU2pwRQYMjXvUgfqd35Br4KJVnIhxWk+RgnD8tZWBY147K5Q98
en8KZ4f0e15KTy6U08+ACNs14SJGAHh8zy0BV5voIWgUTz8fFUUx540jj7jS
dUJiVoFMUSntR4xQDLxXwVrh8YvCeuSTXaixVpq/YeX/akDRnMPMkl9UK8sJ
MGPV2xGDv0cpywTW4PhFtjr0eK0K49wRPdEikxy5Xru3q4IfgmvObcDiPwUU
pXo9I9D8qVAoM1t89WrLqGWrYwvpYTNrku2huJb307xtzBm4SoiPAxNITdK8
7G6JLdVXZfAnhyN6bOeb/uUkpXDRZ69/741UI9Uix2uDY8+otkPFPsfNV2X/
Sw7g3OMrtr2Hgr8/hHmQGwX8S024KqIr1vLADgr7RY6YdlidsPGqEbs7E3Lj
QCtIFxvjEPp0qb15TvozVBklz4j5lnlmx5fxZ86R6p58VW1briMgoN0xKBGi
rdbKHzxF0B1SBC5sKmv9H84HXxu/84XDb7URt8IdW+Z8WNMHn/R8931wAkQf
Pcj73ViDMDlbrvANbYFK4McDAja1DX3aGEWrT6LG3pCkf+2uVlrlGv6I4zoC
OGJRwqrD615hrPnzMbuBcuK8SgXha+uu0LJnAPfuAZXoJwI4fYvNn7NJzlUZ
MIoC/UEFVoJF+5j+xCOQGDUFJJXeMw9Q5s191C+JnIeLoy8BD++qD/sHmQ8n
0F7tvpZq0ac0SSC3u1Ap1UVev/WcX+E6+SBxUwcHh/3lCynCSmoKGSlM5FE1
vB5NFBm6CRpshbdUI2ZVTMPrAZyAinqb5ONw677Q/s1ZXn055BmCxfEdfB68
0y5ikEdcNBcFOjhQXz5wj4Ni33O3/WX2bUgi/ZUSrNE/BN51bDJmoojIf8Y9
gVNAeVMnZUOBPprr2E5WXgw9/OEZXrXqwLnfQ/UQwpK5Swzl3+EfVzowu7wf
O1tj2ZYs5TOg0/xvVhh3xXPe4TKzdkwqW1ePIgrO28Fdr0tiyr+L+yyKf4a4
tg6LfFtGLwsrqIZAARb6irVSOWPUMdboXDS7O5Yj1RaSatJ52VK7ySYqoBUO
tW/SJPAEEdc9EDAKg2IJecci9cdTUrPL6IHnXuNu0CFB+1ZlgVZXUr04+4ZS
P/BRxDRsYGIKsGowU1bNtAZb9Pnn926HjXXvHiIKY8lBoXOFa5z6D/9TPvVP
yGjGlNCRqPRf1uGLqsy+KManMmJzci4rIjWF7rl54XQYNrjJS117oIfXNAh5
6nF7EP4MT1EfzxGwIdXZFPqSmn0q+K9u0I+wplM4RBtjExaO2An8Gy5hSLb/
6culqp9s7m7Jyb5+4zBRajFdsfL133r3QHpWrduTISNetj/KYEkaiB3KZOP6
mk9tKvaALNS0T7HJT8ufinpdJyktB9eCcxrCdihEMW0dgdlQbafD0YNdGE6F
WywTazET5WWQK5jcyV8hehBsiFmF2auFaYVY23UTalrbCrQRbZjbjW2iwtJO
83Uj9PqDd1CqbgYYDM0f2xMzQV4/YdgrnhaWCIAbNN/RweqnkFkyn/iwBCmy
2Py3RxHo9RyBENtmxCkXYvPoP0sPBBsYBL5bcIjpKDIepPlTzig0djN4gIaF
axjcWVyg9rcDUjPBNcbRhXmW6QSFyK6A1gGuacAlH68dwWE2kLlEFdCq+IFq
T7nTfAopp/hqAfEgLm7D3hv8Zf9Vteddw5MK2AXNl6S5vdlcNd4YgkgE9CzY
UbL2sVuVPpdUUbVWfO2Qfq7A06kp4oBsXiBf80T4tB5oj9CEBm42BP7PxGWR
C54D6QdvrleZYXv1LwucdPKOnW3lbMxfmdvMO2Oeq8AWMTAb9gZNYCjPFtD4
tvggeKsOlpT+ehMaP+DORNFOjSKfK9d7NfAoRLKp/A8Wqoqb2ME50oeb0BF0
szLOmwx7OmkChJVkTW9MkMKQbxYkIXrMaoZHxXpGVts7ocf0LoiT5WWAG9zL
6dLV2sjjKO9XcliHGpOesjHrpFe6JJU/nff1VM5T1MAF43UVP0jtcjJThTs8
IOEpgnxojig70Z/OqDQMvERDvVMAoygP3wzye5jnIzOCMxlkH0n6lpB9p7st
Y29EprSX1hN3rb4EZsjo9Ww4frsmS/gAkOJEJ7GoXeDnD+2eCMt69bD+PkHb
LGdc8r+2D/dsla56zTJA+zyyNioK05lqdY/9K0LvWEw0l2E/toD7BM3ss634
VBI+dZxOyALQ/PVQNl2I9iVsassINjDpfQUBK8lr6XWi7sIgWI2Vt/lylP2v
GFhb9bZYXFb4XWSLrxkmx6yqKmGvg/b+JAdXalDt8UJD7P+Uj01hEZtl2xFd
mVIpmLOY4d/RBDx10cdOtnZRhuwfHo6VlASPhm6NjXquS7GEgT8FG4WiwpUu
s0jhlbkNJa1UxiT8EWKmqOvWZr1ZKZnZPzXm51xZqsrKMV8HzJo3HyISuyle
x/ycLCRveZ0oi8fLHddQwVmvbLQ/buQOXfW0nt9crZ4AqczqopikWtZFdn8j
uETkLaO1PLX7cMWxslSuXW0+HfTlyEgv+CQ4UkSU/61DsRYzAFQ8a0Qw11sS
j1AwqY5popBlhKHrtjxKuPQuMLzZE9tRjeWBNEZJDWVoXU7DFyQeaVQ2rLJ7
demOVWkrQsPVrXpKJ3WBhMb6SkKpLhfQhjKcXVDxvzD0tBifS94LI+ew7w6G
pZ0GidaiwT0VvMRrW95bmjdqET2ykCCf+t5wj0tOs1SJ5loX0mKiDYDX0ZDA
KDMDWoqWHWiSb0VnYIoyxYM3iyUbR8pbbVrjIckE7aTD4E51GsdquWfB+M39
B8PGFfHOoTmc4P6hAPn06F+JN2jK3Vr1buC7ZOyS85A+lhWG7IxOaYoz9Aoz
ZpO6DDuWsrWZg99heHLmzxGi+R6tLxGjc8EnImzItxTIYpiDi/5yDZRqcYZK
smUxEN/8Rt8nPReID+gAyiSW3gszhmWDZv4WZOVgOrl1Xt2cyrdo/UkH958W
yR8SD+z3bEGKGQnIRamwWxbH0o0iM7GzQNgSqaHjyXDQAIhfPAEL1qJ1+xCF
mn0Mg7u7yZkt0VAsx56VQO2uy1vs43qbwN+T6OTrvdsA3rmPd4x2h8N8u4F4
1jTTav00tQjQnTzrtdMMNjsT37FXDr02q29mIXrin3hcJM2X6IW7TnE94UpC
+npD4lg3SBzz31el5RxB2rD//uEQ0dHBcsbwcCPL5OOxoyuVPSXzuJGY6Ngp
c4yIb+8xvQNGrW8r/ZynnornowU4mOCjiztybMYFYRJg4+leyKIIUCDjeep7
n7ALQxSQlVH+Kn0cmP+ZDAmXGsX8AEfnM2txzjEf+yM0nnF2cgtetGypUQiI
iZeVmhDBq02PIwQVWZS6M0OED3LV03yUFUDh78IZbz/fQpsVGPbSVFtpwsR6
BjT+x+LV/VwOq0SrF7XA9ZHGUdMiYCzND7CPUvsFZNLMgq2GcDGvGhnOmwdr
tCRaF8sVOSQcKs3d5LZcRlmmPFX/7kATEs21tuc9xZkAaif1S64jPf+adl0W
mSNFvBEJETKPFWCAlE093dEtS8E3b8MRMxBnTdOGSfyPam2N7Xm0iYy/IlX1
xxVHmEKywLQwP8lJHTL8gN4JoigZ5R0KHiUKnq3vyULQKk3YV+TVMl3xdI16
3H4rtEKxXaBHFP0Y3uOUKiSUcYURn8yFz55LtMW9eTkcFyXnbxMJdSojuV1b
6jUIwazHfHEtOgdZuDsV7rDE/M1cCc4BuUWZnXuPPgxy0mLnNqJt5OSf2ju+
MIRIIyqugEyukcKk/jFwhzn+cl0h+9iHuUYpt40XAhehHAZuVGlBYZjFio/x
WlNyCIN2giGrB/r0LVFEwPv6y6m0FeDn1RxrtmXBUam2+kkX1iRQyRty9fuY
i1CEw4FgwH56mpBQ63pGjwAhW68UxHVxtDS3LMZx/N30j8j8d13eC+qdiABw
QFV+e/vL+3ZLfQXh2AChXtfqK54ZG9LGizbkiD2vbEKKluZAJ9rj0ymDRzdx
ToNTajOOItpxsZNV1fZmM7h541G5R02ouRjvMc9bm/x/CDZTuBNePpThvfyE
Lcecpr32a9YcuH9nWNAnxrY06m1xWa4stZmIuJFw8IwDgVTljnLUzfto6nkB
K4ZBBAstrVxKqvwkR7gKyRlBZS4t4tRjUNuZeVRxOCjQii72Dc7FE2yQoUqz
3bquB5yPBvFS+P4KmdYVSlYYUfBfRDU+xdx2df6khxUpEpGcxMcjpQh6Q+gW
FvnY1N6GkC4MLElyH9QwBkJJQtLPPlBL/nz52lfGy1TwMLwLM3rwnfXFafvK
LCNH+x49izP5MxCurPZmP+HL6qoKYPzv/2Uz9y32CbKcVTPgsNLL8f7Z2lrK
eHeSmIcXQFIuG11ZyFmeSZnsMUWjHYan1BSHy5aUlgcPatPgDqxk4xXfBhUf
Sd0EFjdXybRia1OMW+fTflCZZxX650BpyeI3VExyogEPdTzXgu6GfybC47PM
Ai3uD/05To1oFtTNBT28kH5ogfM2YgFQ07Dcfi/xA6KfNeq+uYjCOmEXKBi8
WfMeS7Q33vhlvsL/XaT9MjFm5w76Gc2xtC1H/ohEyH/93EnZIq/6hDaEXs3A
bS2jgKA8v8hNoJnocOj9i6Iwq7de7R7Wjgyk/TGtelJ7ptAFG5d0imYFlG8g
xF5k2SBaqeTxpDfdJ/fYdE9NcKdQUZLDf2k2A86CTqNUsomVHaBw1FrgXvB5
u3pZYvnjwefklL+W+c2I488vSHEIIKztWs1HJhlazWzqW1knu4QKhGoin4VY
3OejEmVBl+xWfgHwTxzdeoRPrVSIB4t617eqIBU4RFZ+u9uIk2OwvSA5Fm6S
FIjnlUtLLoj3V6XZ+wj3n9Rwh6yzpcsJ8XZ5FFKA1BRrnO03iwKGxckjzSBn
nYjWcFZ109DvYox55c2OF89MnBJvBiNHBYSuU9x4CLwFsSJTknS3bADzNnoM
rf+ZdO2snBM/zJ/XQv7t6otJybSF6/X2iDasG1LjiuW5GdGfgUmuGR8vtsQP
OY9Pgoad4ONFeELHF5CNhV9kN29dS3YuHZ1afG6G/cA8NebuKXy/QquEVVve
OBn3J6EqSzS0PAR21F66AFRliH+7F6VU+LZw9xAvZFUaT+kZ7KxCAqCv77j9
fWoLEmt+Eeh/rRsE1zuMTo5dFTUMzdMh54rL6t1/cGdY2ERBRbHI9nnbOm8P
9igDDpyrLdhy3DEpKOvDi5nvukJrT7sPl/jhBCLy7lnF6PqFLpvBr6kanr8h
yX9jXXyqj6Z268tQq18nh+EzTB1UklojwCsyh2nL5RhzqUAoSLo8ST4/1A9Z
bWURE/0OXR901UgWTA+IvBCin81bEB83kJdN6U4cqERddEfJ85oQeCS7nDt5
A/2uKwSnkVCWRR02Z4RP2t6uGXu2sFaXblrHU3PUS0MIE0+YP8oKd33Y6imf
cZuA+/lli6UA2jUwWTxfPtNktVlm8/S5eFRknawTo0hBsRPysrtsIW/kqyGw
6e1EafMkMW65m8IyKxlij4ft6JgUbcP8p5TevwANKGXvvmIARSly07vtsBsY
+f+D4VJ7zhavfU3KYuuKd/gI1GVEAzZqjKrb7TW31jluevrySNPdoxlG/jkw
qDCNzqNCba6BSr/pQCX/9gFO6hWtKsOzV6HSOO+ZKgViLUP1LtP/UyIthVvq
vV6YZhAcfN0DM0m3coYuxGF3GOW18z+O1LrI08k/cCpKT+UqhFyti3WQEMW0
JckgdWt3V9Z1B5JVQaRAPOnl0vyux5aHMAkDI3upZzVDD/dNFrcg+k0cCvlJ
nHMHdQcy8jzmj1PR0uPFcPgiio4qWHWD8sCEMJj2OavnIzwTAkSIP21BeF2p
Kld8TzCimsD+98iUSPG34hg475dDeVa+dDkB5daPhhi4bflcy0kRnVT/RRQM
TYNIRnzuIfpFMBxfsMYIRbyWTEA1EZm+yFDkk8xbGbw54XoivzhtmPjAQdVt
KJ4dl/boBkA0UpGRQcJFCPjuBBX6X9dMQmtc7GF7EN/JYtLxvWLlhswendFa
B+dAqj62cGnPUXaPItCZfTAMZXYt9fmcZgBtvECB3lPOKO0T1pBLOW4zVmMq
fXoSK6jgOankCagEaYNaDDC8kcf1hXy1IdvaeHEFLSuwPkYNBco2OqP24wwN
V02JdGgfgyNWKEMA2omIKidcMlOvQP8x1PZ7G7szQl2SnarKGZ2h8BdvCJdj
x48UbjA6h+rKnK1sfDRxJq/8P76Beu9++OE4tdF0E1pOBxj4oyobTV0g6oH5
cDp3q+LxmMYFwHhXBfW5VlALZIwxQx5HTACnmkzTU4+7OVnM0SD49Ok4U5di
b4kIiT52I92AqlELdKajjEoZfEN+PH8Ren9prRLsvKf+MoJ0AO7NcJPnXKNF
F53s96HcCyw4+V2wM/RIKR4GxxlSep4ENddm9xVbIAiK0JDBiuniRXbH05Dz
omeqonRbtDPapwIoXUouHNvhiqHV1QWyiDsUE/M96PjeVo8VipecN6vgcQNd
9qLUAN62HmZF7/2CiKfrDINMJIdYGz5CQhQNSp73HxIrCxLU/e96IrXAQVey
pNa/8lMyJbroUztw0m1WOGYjHwVSta9q7acLknGEFDFlzVK/Fqsnz0NS2hkQ
Tj3OMmU2VykLUwflr6RmbGfz0s66OYI2RmlQfMWHNEaVEOHuBj1Xn2Yj1gDN
dQ+0w54td9ccxPglUzWYPX8ATkrrPDAaTPHt5eNrgjim0BmeEWsrcfs9RxLb
DNA5GUoxDtGqirkz6I/DsnaFLLRowfpiSGXUQCTDu4IVGz5JRoeY4ji/ky5a
K7SVeNSYcLGCqHw98FU024Hvymgs6SuLrVyYym1RMDz1+eSzk6KdaNt+HNyw
gcgI0ph93tZ5xK+HahUFqp2VZPu7cWhUj5NH3kCkaAKZc2kbTahW3YM6tvix
slv5gJRbD8dnhhIqt4txoFzHSg9QVXg/JXhFv+7t6Frz525FN32XeJKPunsy
FZ5lW/1R/6lxFILbw9ksBHSOh/f5OWwwLHUiscAiJcNaO4iYx2/IOlXfJTdB
EJ0fpNCsiFOcj1ASFXucZLL+Z1Yg8VqL+IT1E+CsyErcY36TQI+bb/JWuGk8
t63OvlTJ+Ay2XmJA/w0/8EZg8CLE2jmfg3bSvlXDkWqlbATdUPM+xCstXasm
wUHgIXg3HhtmRHELWbT18uNvIB5Y2uzMAkc3q57HKqXEeoPaQwAiz1dOgcv4
+RNX+p6IT7bEWt14Xg4tsLS8JArqMhe58CrzzlRfzh358yGHGDKfb5a7tXA/
iGdNeXbN9Qne9Yn0R98VKVXHKNTG7xz5VleUtpKDDeI+HZ4imBcR3YtzEWFS
LS4nNxBW+pi0GHxgTIv7biiXdT7gLUR2Rkkr2xkz1vJvkGXCtSYMO+tresco
nQMsiPom6Z816KMAfy6zif+uiu9XUcdH5GZjrgtu8dxv6c5gEWrG6PWuvXU0
VnkmIg72UxlQViJ6s4aKPTrXC1jxPWH4jl0mtIVZWqDF7ahGFDZSv4aEcXBW
YocERcNVeJXnK23B9IMfSG6ySryGPZdWZGEb4Cy6HFdiV3+45Dj4sJs11NT5
5xSZvkKk503Pi0R10ex+xNv8hk5gmRcdC5le18AgOTBbvK7Oq7URjmKLQTim
ghRiBvkpIy5W/BTUKSb0JuXwrUvWM7mMuqXqu6EhGZtmX7BSTtFvtl/FJoTc
PgLPzWp2F3OZYfGFgcx95XPhB84iDzP8nzXvrdNWXhDc7HNHM/0njg4KrSCY
EvWyFUfuDhJP6pxRT/+KsET8cXccGBxBcVgcPXHG65nFdYbF6R1SIqF+E9Ep
gYJ9umZEkJH24/fuLjQlup3ZLJbNk3FRiSesiNU+kn4gl0zfpAvjT9bucm4H
o4yMlEApGBi6FvxEShHznecnsoul91SOytjOx6BdfG+WohlYdrlvywVxjVKQ
y3M//M4PLOhk0SNPlyz0a+9i1UXRYRqYrQHwWmT4jtpKUucPBbpRoKfPCnUL
8YEyk13h9X37vB0xUYx96q4BnRtHxtV3fkm833GaB+B/f2GrL2KYI0i9xMq5
Mo36pDSNorn9day7U1WQNHtmO/plO4LyrB6aeHf1nJypp2GnYTU++al1Axd9
uLgQx9oLrC3iG0OeaqV+qV44RvsiJNCpBAht6gOA2Yr/eO7OmNME/JnP6mAB
/+DBuM9pWybjucG9spZ1YeLJ+dSoQFE0T2IThyp26aRnkYA1AeRLivwXRG4b
Lpy9y1C9bJ+Pmt2hxTFj6Wr60EBeRikovJY8DpoGNkflN6Tz9rnO2U0pMzHH
40qcPyQRzdE7bdfhbK4oLthPgxl4SdkcC3e51MxTbIEWjhhkXrfEq4WbPRx8
tEc77EvYMCUORTgHt3+8IRLIPbh7Q+s0++2/UCvhYLXyjAiRsWE1bCszF+uO
8nFeYx9CxI76VdJQX1d3jQGWC94V24tA1Zfvtu+b8fJQ1UESZcDh89NeYQMh
rIf4TcAyuVJGuyj5yv4o1Xx4uJIVTtwIH0pgmwUMIsZFIoWf1niGzJVN1uOe
phi6veY2iXpONi3ytEVCnVdu4hHMVtnoNN7TD+jMtd9VbCKxAe6PpRnvcEgK
H096CZrX+L4uJ6yWkHEkhNXvYaah/riaYSYbIYsqjuYlOOKbMQJumZJ6P++H
/OgphC+enVM6Eg5jeuim1PZwH5BxCBRz52wwLX/XcThj36gzOe+TE+tfRGI6
ecfuAd7SRb5qpZkfwiUlt+WhgzD27X0RcuKeqUKG0Af59AOVqsnD3REjONl+
QSSkR0688GUJ7k3FBa9sOFOtf0EO1MgTzd9JxegIdrc8qjx9idh+mNFlS2uB
kDI4to+oL8AtOMIDGnrHx8yUI7IO3qC5LnFCyOkMe6SKJHNhDgBzTnZfee7o
nWBWSVxVtMcoF8B65jZW5E08IsWkN7jgISo8WjWOdUP99RJt+ykk6bFJDJF8
AdzqaGE1Ju21VhRrCVJlWNnkrMT9hJ0J5fnVK9WUGh2Bn8pGFnSGT0ifPt9G
u2KTTAkiAUmbXvNe5pPgC9PiQjWJyB/AzUnSslEdjOfTFlSubQD+F837PPVW
YKcxx3ZkHDCPHDQ22j6ArrI9oJFzftm3VF/sshPqG/2LcwK96EMW6T1m1qzb
MdwuAzP9u0XbILheatufuZ/p9xMrhVfZn2NpWrH4OylCT21zyCun7ONZaswk
8pLAtzeuy8p6PMyfOVYqGyDk2I44dQKacO11JGiT9Pf/uF8eN1l4+NSjNf3X
EFlE8txTL9KTzvKRyjp1EoeZvMIzWuLfYHGgfrq2thuPJIdCxyoWFS7ETblY
RBRd+Blg1lsXiw9NsqU8gpZOI0GflOf7Ry920rbTRFPsLt4Bd9PGXCZeJI2l
bH5ps2tjwmPOOUX0aVx6Y1wbP0b5p4lQiD7aCIppvRpCA5ch1Q0Q7JPfTiIt
VzV8SE0bVgZBEAQnhVZvvlgK4ChePJF0/UwqkNbGawbvq6Cbp/SsTltpNjdP
VqjL2lwHKhDmpVHHwzPxSD1oSJIoHWwVp0tZh8S8GF5f2iUs5GU6ZzDIsOz6
4BFHaWAacNR/nQzyPpj3onEgEnoq3Cic3H0ngiOTfVLYiRGTEeYl8nU+s/zL
V7HTayGaQqinlVXAHsmCpSHefX92VqUQOcQJ4RX1VZ6wt5p/3rL+6wPyr40w
pT936k0oBsYZTYItnqa1LctIXaDxxAF1nGCVh5DhJsWzZeUeL3NCa2XXvFFV
P4/CgKc9DeXkCEwQ+cl+UoCUwI+iT4qTfJ8MIm9vCB7Lu0uP78wEVGXzjcKS
7tmleBe67EOOB6k++sWOLMYJXtDXXVyOQkYhMf0NkGoc7IGSEnC4a9c7bBQK
mWA8AnGsR0BnYYSZ7X7Ew2uervHEfCwmytoNGCqn7bnWXCBO3u9JYgow0VWX
VcHMnSjikorXocIKSO8GVy9h+8k6vE2yX1c7Ns+f2kO4M//LSqYsZKtcs570
5iHTAMKFfYBqeqZ1JaehOAjaKkuL7t4vLku+5itB9bax39gbaQUrMepHJiep
UMYRdiWKSLyF62xFC2MAvKk8GeOnzoO+VTuc3DUosemaYih49xMJV0rty+A7
EY4WFdZopQPFOU8O5DSg8GVcupDSJoexDV0j8Xz3QqjtwbACbjcEfEBb7Jam
ESX0B31239NGuPyvi/EgpzQgkYVtIO2Ey59oUR3OIK3Xqv2Asl9lw1CQsfA8
Mkqkur3CPqNAu7EbgPXab3UMmgkh02UlgFgWsfu4tPGWaEP+ItqWOdjjAzo7
lNCQmzWnUzxOtHCICjZFrKU33iqTzIFAfKXsOkepPTRchC3HvtEF/8CKL1M2
PxZtPSxNMH5DBAlva99ze0WLKtLZWcI+aF2KTnpXzh9rAN/VjH098hoQrkVD
iadh7GqAEH0MptYohroPPwE8oK14PonJeB6kojhaj6cHcABcljJKn732GOGF
Yi5WnDOXmNS3wbyGeG3E9FKyqhHd1jFqy+IGYta7juh5si5vtI/gYLCJDboJ
kGBRVgbdmwbVGd/p3lYbbR/5dhnwZ9cHkyyUHPO4I85N0B8YXbY+BmrrABYU
UQLkUi9Hp8TSjWYepURpqObJ8oCBE+U6DITKBYJsSrrGGtOKQKaksC9aiGaB
ABrtlscZ+7meqPqFc+cVJ4v00ZDdaJL1hFuGmS3Z03ekc4XpOXxsGoax/JWE
oZ/RDY+Av7tFyFT+3wmFwf9yt40D4wuSyOOKuurhoLA3dUI4D6adFBvBOoPi
PlFJU0H1cRdy95yL2MIdD+ENhO+5La9wH8cpGARqde1GXMA+HA5WTptNI/bR
/o/dXZKLCapnQSz7lFa4WSurFsNvYkhUPqzEb8TsZRr6LJ3V6OcmJ/KU5/5q
PFPqrWUEcJFJw7EbSTlqy2W1O6L5asrPYqVFbeMzdFMUluhhQpkUvqrx83er
k9jWQHWCF0yRQeCzxh33OyY+7qtLLQwmus4ra58t5gzEZnpmPBCzuo/ccLYg
vX9NXWsivxri1dFun7sUnf97P3X8l02HQUj7V50rQPtovioQvL5wIbpd0n3y
94XqDL0lwBEiH2SugyYac08YToEVyF3TQTKTsvO7ShIlfTXUoARUq/nkAYUg
lwcEhFq71NeozjOh4OET5sI69z/rDh5rVxDchftFhRGV8bciD1lgKIx91CNa
zoKmmoZ9nlG+CUiHPYHte0JGcyR2EC+qBhvqBSSqEQKGfSvws4JndUheppN8
gZb9+TZLtxvLjleXda1epzk07giZsbuMEq+T+1Ume4gKq/EMSY7wHoZwu/W7
NY/VVJ+0lMKapWf4cg/esUSmrNsB5YGPBcKeFlq38LDEg70DEOyPIYLoPcn7
NMOgP3TzmCaGbcH8dxslfebn+x862Ij3T1KySJT0R1gYLOgaRdkQWcVA5wOX
BfyoTSJpjpzYvBJCSCdQifIYPrssMsN+Yk9dSaXTDyzJjXc3C55CAVSF67vg
aaq4GayaqqGYgMPZmNfI6sKDnKhoTfXNGz7K+duv6GMqkyx/Q0TBSDTMmV4o
ucGKZoWR19WGMjuOJ/GuiANRwPqIjXWQDIkPsRAhsXTnf9Wr4q0j8Od0BPf3
KhqhJ4uqvqFB+swO0BQYnLK2iXywPiSHTQJDenhvENFNk/qcZ/WIPm7P9MMK
FXwxDcQ1DT/MbLQoOuZXcY8q+BFWec4n8A1FqLXuocRxfgL+6qnUAtdkEXhy
bDhaeePwRukjUYyjcP9VxAHyReDMuZildC4Xarq8DklKMYZETdPKu5P4NBP/
NSLa2lP6wsQrqm74ZNw/4ShqLXHXRnxZviK47UxJz1qgsbsbKtPyuus4vLmM
da6yHMhQs1mxO2jOVwwrDv9gReIQ6/VEAeBluKQDoh3/eQqgCmIGMV3eDgZ+
5kL7M+WM7TYCqOT/j4Do22DfTuxXfaGMOydgQg/f5TaviBlAkqWckCfUebNf
dNSJfKCtsyfdChIVwLSVxxaLqqDTrLKXlzCB22cpgf17EvgFY49OZs7zJ0dZ
iNaz7QLIMeWONa7FFJ5M49EBSVvifmKDNekHpMHGy05ch2pDyJRUXbkSiZTP
8ljAKmh4ZSfRkGOI/qUSWiXHdMocW/EcrOGI+IcSwROROs3gzOslXJBmLlRH
/OPgi8tILyBH7VUH6Czt4l7Ad3obDFB0QH9i32EG3nEvcU3SZZ7mRKBYleNy
kj2GJBh9SGyUh3FVkWzRifR4qUnl8Rcysg3Lca0AaTSlJKKBS2LFL5VTaOEP
itG2yd6CrpotSSkjEpthraN5+ppKYm49AfYd/8b7DbdryWIujxARYk26fejz
TXs2ybMhRCFP3qrTvrOIzemWGX0QOERswLb3tTdeSc5MtJaEX9UtbcLu6TIm
7iSifaZbLHplVlUBTGTUeJz3OOoBdPdjYf13GCEBng87HLpq/4/WH8/QmPL9
AF5KHGJ330XGPWUL7sy5Zsgr6+5ypP3SKeVZe+AxQLVzBFIEmExMhlWRLpiU
J3XCnWm4VuxijZnvsK8DOlaq+VCB+OKTR0OLojXfMVrssqOrWO2iJK0hDr7l
sMjgK1HAe9f3CuoDfyu4oK+FaAagSMI9hggpuvmvIfI21U8jcJ7tzCegyVux
YfC5QvbwSoDY2t6yLTpaHx7rKOZV2QXePE4HHkgWf1Bt7P83n39jFVOV1fPJ
XdpasfTR11t0OpEqwhnTsgCTXjewvRFFlY8a9v1fcot0gfQIPYtty9teluwZ
evnOAW9uWbIik8Ids2Iidn4i5+8JTV8aOfK07yHN/xEdjAYMIHvdYrbgj+3A
FA/tzoWqAO5aMp3IRGL2ZoohEmcu9IsZ9Md2KUGc0uTwgOzS5mKIBbWRFGW5
AfrpLgeins2nt6w+A30e1Qs+bW/Hlo61eGIyYk3BwnsqzTx/qZwjkZf6+uL3
BrYjZN3u7FcKXmBEwzCzcw4pSwpJH6ijde4Vrs+LbPaDhfGZeUQPZJqe+H5d
J0fDbIzcYgewB3wxO6kCPKHXCk7OQkjhOMe8C2h6bC7bf1p+m1WPODnWcpt1
g2G8rxCy9Y02Z6yUhxP7xjKkvuz3nrrFzOVG2BMjegDvvFf7JOLJJljloHdG
kLVPsJOlENkFX1+Dt+ZHH35IHA3r1HV2fr4GrKWlj868+9H6poHHUI+ZFeT+
kLocQcif0XmBPv/y9/oM50nKDVkl4R3aeEBEwdb1RGvREg5zXFsgZBB112Gj
x5ShSbQvxDPUJD8EHNoid0vGduk3a6knRtt2p/LOtuFXyXqw80WIdDFmYGRg
LVKNEvVXVseHG+dM4Ni7epJuFq9kSJUNKu9u1x20dtt8KBDMUtAEdHjLCfYc
9URN0+aaF8OLQCYWuSy5bOCOmtJetsXAdM6rPmXzuo5c+f+M3lw9H7WYvyUq
sVtzc37a3J6RDNphL/2sMkUs1JhHBSPPvxYn9O8Yc+E0WC/uVTAC2MdKAMMY
Cbyl+C1j2C9vCJ79Zth5mezfn7moSML9jqk1HeoFEQUoncMuadxnglY2YjJz
D/u4+i7eJGs7XspZVffZq4jMGTvcLioPUttJ8t75B42/ooVZLyoj3eIVrZKN
4YdU235IetQWuKeNZ3UbcvinTy0f0qAg//9OLjGckalJKigszsAL3i2rUP/y
VKxkHuWZuVjwHIVmC489hipemevd0FMr2hrHPzs9VCbiUINYtp7mNsdTEyn6
DYFbo7MuPvgNwIhwdzqkqnBlIwRphkUB42g7B+8x37lREWFQsFfVeo9GdN0+
nSx4/PASXeU4moeDuGun7rWGvBKcCEJu6dawaxb0/YVFQ1a/ge6RUDUw823/
3LCs+TXVS9z90K4qmcuZdBzwq1zFhA6zPMs3W1nWps00lI+y4P9EyOunu7qU
5cJxkd2NMLEv192/7EMMpCkQwrjU/Y5JhXiXP6ZZA7BtORJcOGCfK5eVsCWx
ui+JaSgNZH9YtJpWlZF+1wtVUB9Y5Gwz0kgk/A6+ij11eCcK7GRBJcwmvjrY
5+H0H+HSdpBdS9mqjmHzylSGuaYNBRlWrdkdnSmsYz6dm2r+9MfFcsnr1THh
gWfK3VpBSlianOlwlN4PVrqXBX15woMgOcDVBExubcXUrP2w1rkThz4W8JEz
j8Jt8oajbLvmM/1bFxCV13YDOUjCaWQL0qEB2Wzb1Rxv90Clk0+r4bhMzWGj
q8EWajobaNcghraQKfAzz2jPJDHaOvYtXNTtEQkeKsfFnxs6bVIyVPukk44x
A7AORGvrM9bNVkrb+QDwxuUNM7ht39T/MJZElus/cyRBLmvA9Ml/vfBtxERj
7RwvZVodflvdYCi2CE+ttcVFT62dz817DJhlaPA32oxBJJhNyn8Nwhu1ZHqG
XgbpWOP/cx9ESpUHGkOLZUaeFQ2po8a3yvIcwXR/dvCyUWBbD5SOpqxJ3UbO
PBFwdcXkA1WOqZQLYFLueobOpDyNqJfUtztABP2oYO6+iBS+7AShxZhxSgCH
TxlxC9QG1gVslRYZZrBNKYcvYq8QKF3t1fgQpIFvZEGMF6oocrGAgTDk0w8F
5/pgaq6/wTSRJrfxW5+3MVbFTC3kZuPcgpXpymptK/R898QJX2nLY/pE08Pr
6Uw94gwGM96QMmn7et1b5+T2FKUzP33Nuf8C0gwDEjbmUCFTNYhtsZOfRc7t
dZFDhCFqKXhyQTKcF8cluw5BF9HpeV/rH/MWBIM2dXjYZco14VOHCLiVYzEG
zopAcstrU2hONWD/7EQjtJh6V3bMGGb8P+BNsZz1mbfzllMaFIvuqlZLzp8j
NCUVmHdesnvGF3Gb3v0cTq35VQDy+CDA7nHOToipTW/UkYSjmXb6VU5hw3Gu
uYIqb1q3EroJRG8rO2vWwgIezQ2Upq3qQ57y+mT3uTz6edvcROIqbH8LOn6l
H4b3JW4dPu9pfF7o0xssdE579U+a4fX1DyVudItfzGFn5uVzd7oX6eUS5ys+
e0hBY4OEUWHJM3QGDKT56wCVXv/1F4qCP5pfr5TBr1WWhJEKpoi7bWP6z0GC
Rd1zfN4/qbkB1Ya0cw/9OJahlBbW/GVYLhjIrnYhz/nGtZ3T1D8JxcYdtSRs
WHH4Y4DaxGiOjP4R5aKAcARnzYzv4ePw+w41kJ9MdCMf9A8qK5hxr+3NmLRF
IGr7y1v+Kz9JqkAlcxWSwGPEGMqc9K5fxgRqkXIWmDKQVpKj6vMdrfRwoF21
1+1htnkQqL35NkEQzA/j+W27VdPIgcKsgQJprBGep3r4j1Cjk/NQm0WMWvsM
UEZDpkey+/ZTzMfyWD/pL+D9VZAth3tgNE87uDjc2inOt/iFC+o/wZFkMzIQ
h8T1vSORiFLCEUjYfClY3vk64yhOl+vMvAqzHklEMkmxUksM8lqFuM4O6Atb
NdjcvGTEMnIZHg0+i96HY1Z01EB7Cq1RFtTpFbqsDKOMfd9djyFCQ2tTMMUK
EpA53h5NFebMrgJ9k3hVfSyrr+6/22HLBNrlr4Qx4QwTzbyTbSbumpShShFa
ll6DgFiF9ZtKXY9YBMJVJgZaG5vEbBO5D8uOncJnC02xP+/ibaQmfpjiXpDf
xRNatICV1XfjVZ2EujWEP+O9ffvhQKXlHeBUlN3ofSsMlFhbVYIKCB3bRMUx
Grx43PWPMYXYn9vrtiqmZQjj/s8qhBUqRlKBWD1fC8HDFSF34SsnDY5yU5XA
/yxnWBfMclmSIlb/VZh2lLUda64gsfwMPV830Nv3zyHZlvYAqYuSPgGUihGo
Eg5PxqBXYT+m4l6Dq9UkVePYCOj7pydbVJAcVHt3JmDtHIMuf3bw4YAc2en9
Gnf1dRgVbjkEJ1G8JFSyqkJFOQuovgzgoVM1epTgZIAKAW94i/sWINjXNE3o
BzS0eZG6t/fUGKST+FeBbmwqV72nxcJuFaJzZsDWUQGdsu/xDpsPeysVxNKn
qzCMg2HNSY3agxdqFLtLBSBDc/FoHFlJQv26OHqCPSLaNmSFL7sip3C11IsD
pOBN/IGwg0XyAUKDqwffcNyfH743tpmpMmgqFcDmbaZbdq8TXZDC/moIkEWe
/Nt6nGoBRG5xudtahrTZxW/g3pkat6Pbg4c5Knc56QHWH9XDVivr0ceGTwrj
mNet8JeRpHjGUqq39m3vzFMaM8MUtTf6/XM7AxxOrMzXbTm5kAZHY6KIK5kt
R9mD/HkzGsSiBqEwnL8an9Lsh7OwAwyw25wzy+ixisqrmc5T68+B+5awH1FF
cN5ZS8/GcrWwTSo0p0U5mSqcdRF/wfTrB27v5eQEnHFMLtUHuXmndWfo9bwV
wU0RUU5kOm1NFnl4errU9HT1FgeP+gdCf4CB3w3j5YVO9Fwr+GDThQiH3iGD
5DlRmyUzZcIFMRYXMfl/rYUkq19pCaS05S3G0UeDaaEXdAWi8nwclbkemh5v
RQVBFKpnKdfQzjE7v5lMPyD012IXkBMTAzhZ3hj2xdoh7IHQOJVS5ThM51CY
4A1K6cVjqhRvgPPjioudonYpd1daLyvUg8Y1VYQJjdVbuV/KijlpaxiUOI5q
ZEmLfx0Z0t6yq46MxTO29UYPqtqs3RzuXjKyx7oNj9WaKRcI9KhMPMGCSQY8
kfHS/T0T+9GGZGcRJ5gqzDmYZshOP2plDmAY/oiSjuowsLz897Rcgg4olNJW
NO/QRtY4NR7abnBcuDMmgM443/zvSaIcl5b4sArHFahzxa3vusgrAURDzRgq
iMTPNpGAM4Q315hth6xewkvgQtuIkD9OPof3vAqCkIOvJ3qe1nFINJDvYb/Y
0yTLREBAsdMU0gJhbACtlchAwRNS5Ssj6C7l3LCsk6twnGlIECGL4CiMtPtd
rYDBYd4oeM3+1jrMpzU/7iDuiqBoAtnQPZs2kj/UbIIVqYWll+HOojkJEcMK
t0ihxIJ/XeKFJo54jZyMBhwAT7b0yXnLUej2i8R1Y2TgR4e2gAOdMENoSxZg
AXoT6hU/vrGCvmlxUVWWFHk/J/qvKfalU52tp/whNu8TnDqqqg8lJLb0ta1D
EXmzE9pvPq3x7klehsr46EubUyuuVIb0LW7acPLBBMKTi8tvfMux44n0JDKM
DXKsqKohXHNChv4ruMmoW4WFQ0rO890hfGtMBXG62dsBZr5rfrB6ILep3szx
0jAEtJzVejtL2Diuq/PIqYbzajRV1cdDa+IL5aC/p1BvS2mJTCBRP5KGc/Z4
vmtQAHd9PWl66YGNTD3c8EJ/bffU3fO1NEVy7oLelFYyyTXagLobHmYETZg6
k6WgZZ8VTQXtY78jvnARLlHTG1C8g+yWnfMmt/+vXw224I/JFL5hMwe0/tDj
8iAI6qneqHbssY0ENE9Sts+U3Kt0+Li/W0EyFW+tDC4PVq5scjc/VPQyszOl
ZCYnhL2Mf0h/mAVv+TPh03ws1RsnxeN0O1M78D4iZggwnN+fKYMX2zCZGQqm
+5jFvVoK8+AF2X/LhhoLcJsQloMdE90GdWvazSGIqm99FJmCMQxg4rDhlw9d
Te79N0iXZDYW+7dcjtxYpZRVDXv4C4gPY4lOya32aSYJk9C/YSREL5WI88UY
sLRNahJGi8YufBLpd2BX+0j9UNiTRhPvF6j0I54sf5/xMprajlAK0ASwa/K9
wkKnl8XzbR8rEVScaaR5KC01DL49iZYiDWpi5duR2Lrx2AEdvYZ08AHIPtCz
QpEckGW6o2HclVvPY00xwPAuDgl3aCDr8uwyo7WvyQizz5/wH+IdBWJPnjYL
fXbJKOkk16WnZg3OfggZuJFMEnGalZJN43WbbkbaQf7yeTqEm4ufPWdV0px5
c/MdsI9yOCshQtWnM3T2ZbZZQ7XLJ3Akr5O4EkvXbi2BbMN32A1634eu5QVQ
8Jl3QG36g3PRYRHoxHWx4krt1LLJXiu177JAhjW2DydRHFLqlX9x1y88DzFi
ukQUaT8Zo5UezxIoif6BGJ7owa4hAGb6azZwrEGePwaJKWeDancHWAMEkHZE
AqIp9ZyfchL80Qsm7Djk30X4mp/IptKCNZETvCddKwWDzaB1YJP5t90j1zVv
i+coGbR2lExSPYFP36H9ChGlTGtjsqvZAFkCfYUICTWxgx+FfN1RroJiamkz
6eD6D5RljUb7cM6+q4C2m3j/PjVpy2JAMT1YpDFa1RD+MAczKM1b05XwQFG3
rjPUVOmdq6d+G1WmpAWRxEy4iDwAWEPHBlHvU3wwCNThD4QNhRDJ7RIMLBwY
ecgXz4/N6wS4A3mDGtZ6zqYCfhxxujLXH/UJ8Pfudig4nIJVnPoJnGIFAWZ4
zPp2iH4WuZ99ktfVGWCBdXDhehk36+pH6jXXb77fN7pj51PGWU8fffxwHUo9
j9dz3WBx4GDo5W+nmj/+enP/90XT7CBy1R33hMx4nxfM08A9qUx+XXv2TLYs
emDU+WcUPg+/1Q98Iafz4lTSlVTFWXkaHzM8fJWQDD4vLQyzF8sNPvtXFTQk
zITX2vatF5pB8A3gkVwBk2DY1cgfcGGMTofOOUV/5hQ+VsS6ved+qZ5cB6ep
9SFMcNMocFPU+7x6YfWhaXFcOQ6+q4kXbxTEZCDhqAQUugB9tE+8kexjeRJm
0tCYB7Gz+MmGT44SKnlcQ469m/fQZxxNOun1av5TnNwiAECt6uc9TlQ4qMTW
JvP8mUId8IiEs7lBJ+usM4WWAqwwOi/NHCUot1wvzLDs2YMy+jgSb5NjnWq9
XLbU0cBANFBFPMJXmrqlEmjiywaje8k4WR+nzoi52zCA/dglzkWw7wwgCtgU
9TpEyjtMaf9jEoLDaLrPE48wsFww2iT1oxBGinpSw7kekXBjAf6PpmJXSSsn
qRQawejBJ9RFFANs2ACmMV4TfCjoT2I92ZLY9UcQ7FQA82+UjdSiW4btAfDq
8nU63vdfv6u2Ow/Kmyg2bYZG/qEHY92OefqojCKOlC8WKPkaZS98NoKbXyOn
Xd/wSO2Cb6QBRh6btIJQtlpXWcCaC4nkyVYN+3aQTXi0ygz6VoAQmlsX8tCc
g8qPlAPxQmOwHV1JaYD2NXsxxYwTCPU6LnIv8k7QgSwpWcpsPZyGo3RODauV
Wnyr+elVzogRuoPBEs2hAo/9lkugzxTL9ITSZIHc4ATke7gfP67muv/a8nIW
QeTL47xA48+Q/gxPkZzmpCwvFE0ZsT7RTctNUW1f47O1mTB4QCZ5Awp1nc7b
Dva437zNLivMRYzs0GGyW1te2ATt+kibnhTm5a9HggJ8HPDj72leQznaB+pm
ZX2mI7TORYuHJrlK4T0DQVj4dhYgc5VKj5jE1V5IU/RSo8AuYwJWdsNfgtuo
zP6L21C8TUUmRIIisZJx5lZB08q5tChubOB0k4i3ilkmdru7T561TPe43UZT
qr6z3iIYOIX/WZZdDXQxwfG1qqrg+0WtxrZfBl69M8IqpboTwBtTZbJ2ZRYz
d4I6bp532jY/BfcwEKRU3CZs8b7Vk9n9NPaWDjUjm03pzd0MLS7tOawLEUgT
AHFXaQDj0ZPzBSyCElOK+16d/d/9zpvJOmj+ElVYNGbBS/Dg2P72c3w2CIOj
HdlR+Cgv3nHms+YTe/sOzyhy3nISdQ8cADAMN9F71fCkDDfYRcVXuhFSVyjC
HP7hUcKrfZQLoyNrr7d36Oh+j3kgMLaSY94OP29J9xXY/40UuivzouK98xkS
r36qslAYrQHBYpWKRvjLRC4nRtG3bluwUTDCxMzMJgVjXI777eVGGDt7Q8MX
ZIiOcapalb7Rk+oBlp1UbGslsYFPviu8Z+iMPue7emfYywhSwXL+pZ10qL7X
AxFgAiDFOiouTjxtiGDL4XaLc7IWdQCY4lIujgAnPGZ/S8cu8TXIm8GCSbdI
oA7KcMRe3YjeQgHz3uLp+OjighekVn4v1OMDibXI3EdZ2uj/63PyiU1De0P1
cQ1lETsd824xbhMnHvNMrvM5EQTBKcyiOKH9kOc94D4+7RkYzIZIxp1neXYO
7dcKaArX6brcmYS7Wq/lZGdAMUxIL5zrUF4ktnStc78dhddazbQTob/BA+5J
K8nc/sNdtzN2kGBs/zzmbB8tU2nkZoM0PRm3icnKu16hGA6Ztoxog56+4rQY
9dIa+6LwNGSWHCX5f8PW+rzYpfJYbH2AB9lvCZ+rVREC3gAbc5SAhajQHCJ7
UBquMY8zS9UyOHLSRAgj6mq3Nye37V/6iLZsiqNUTPn3nyfmFeRegiRcjDKU
c6eHsPoxa+4Su3BwubfPhTbjwvGFujNBOuXi+f9pT4YOLWA4MfjaiN3jNZ1i
T5AcDm9Gak8HAWa22Rop959BlpYihq8ENLSY1gwU4/aE1cCKB0ekliH0zBq9
SFty9ZCgWeZsrP5oRu3NyY4jhixeqjwuzmVUIXWEtJ+ocd1axOMT/IyGwA8c
NMaWW+kUR4DG7xYQKLusjk9ODDSzwyQ9MG4zq637AbHoC8c1PuCLpb/9Koa1
ddUuZ1vb3tv9XMARxxsxiHW4MWnznBP17LGdnNh55HHE66I+VCSRJDDF7dM+
OVsW8HgUgQedpq9Q3I0yqWJm3KOUePP+tkS2aWVkSPC/qZ22g9fntdIGcqQj
+1G5zAU2q/TDHShcC38vafQ9aMLacBDIPuDZVm4/xhRRHoACltQrWjYpgFcE
UAx488Rp8luRMOi4i41XdpQuh1+EhpIgLCnwwnUynNgRm4Mv8Npq1tnKgkdf
9tO2IolO2mpA9PIOizFoXGh47WM9xXsp+Pa5TSkhFN2bZT35T3iB+j61kcSt
YpPlDjkiMEa7OPZv1fJKRCqfHRU57SYAzBouSesWPY7xxegl+7fSqDSz9m8o
w7XVFRqb2023y+/gPHPKz1iO4Jn6CPcrIsVDFtZ4MDHOZvcAZRU33tlED96m
GWTFE9dgRCQ8Ne96LQCMiRHswwXuRX2U2ya7VcQyRdKgA9+4CxgGubck6sHI
WB6K+PNpOoZZ2Bv/4caokoBvD77uiGcbcCKa1tyxfyVjqqwA7R6I8knQ/8JX
rbhr+M+zSA263c+7hphpw0YjB8smXiADWwDi0vm2fBeMxlaAkNr6NRKaYW5s
AMlOBZehjRddgROoAgYgfxAyw0ACMb91IsOCsgPcXRRRKhS9Qwf4/JZWRiDm
jsw8ZjVkK9sv19VcdiEJ9H5RstehJlfxvoRQcmmAy0TLJGwtzCkLJv14jsjY
cnuPhYDRyEaNyTutaoLhYN3d/RoA1vrasViDFcePb2ViAFIJ1A1vypg40qIC
wjnZB1WK3/+oVVP0f1fWkXhtYfz+VxHu18FXp1AhKYRBpezFbaiuUB1gry9k
wJnke9feRIR8UOC9tnim9pS7P7hNVFelNjIh99hwHcLBOZeG6f/Rv/ycda/Z
nTM8RUBV9Zd9TAXslaZNFZwQHAp0LbX+6GxjIe0MezrHO68ouARdCipm73OL
bTsPyg9MwsyN+FfHVMPDItxwwYrwEtNADrpkTXCx1QkJnReoLup3UfmoT2Sy
ydozjwO1T95RX3knMOPS4uViT/dHL0joQbmLu6uFFzU5zNdEkM5MwXOhPq4d
lyBrQQbXo72q0gvCHY8fFf2B2pE6tVpcxoq25cvjuz+pUS685Qz/MBUiO4up
sxe8Vv0bYewZDjbZtyMKXjJ01jk6nu233GQjS99Vp66gPqaycA1cbnuiLp+h
lWr5TY3jXZ6HxfrvADjoD/7kgVPHb5+56dk2WGt+gr22+bEDNvgUxEcIbpt9
U5XZnloHvrmCNovD8Nbcdh4K3VC0PTRqyEcLVfpiYW6gakbIkz7uR/750i0T
tc+RKc48PmFjaZ0aeuFdsfLMaiapxGQ+IeEs0nasYFoDj6p72LEd200QHgS6
G+x86s8noq6xPnVZMgIMW+w8C4O87pdBmtHeEhJf0pGLMu0eQN7vDTAWDcY/
O/PFNH/eSZxl+slih63f//M/Hu9gBBERd5JfncyltUU8OmhbI1uGMsNxYAI/
eCaMFtC+mKH+zVpxY3GrYUXIwCajotdOdr+nF+r9+6Aq1Lc3Lkkj41ukj3Vo
NDcv1l1IaXcnuWHPx9uYlSFDJ9LiogOqqog2rAOF/qjLKhIYhyHCXvIuM0En
VbUcDe0CF2Ediff6XJ+xnx1e/QSMUgKVVGIMG9ljXDdO5510Iwf7P46STtAO
Oiy2BUeLVYonx2oUgcY+rgmihxwTmkhHKi+mX86DEW1hrbhtv4QKzUXfeFGO
wNSo1Hg3BqY3DSInNgdXDzsN0fiAlvnBWSKI6TtU95IwC+UMLAkaiwzj0r0p
OPQhmCUrs3nzbF8ABtdjkfrdpk0aIVr7s4OmvpcBwvmuPxlxQDLOHY24ppao
g77i/6E3xOazmf5rQfQ2MAd+wDDWL/k8tc77bZQZxT8aMi1ocVtPajEGTuAX
6z3rqkeoQd6w1tjBrZlKbXAhNeW68MRMqKbnlHwDi8SADLvjmszAytWHm6NJ
a7znVb0JTPPSZikoyRuTd8+IUgkgk0PHeS5UfEcxN20FumgBwbnY7lrees0+
bwyvYjlgnBRsHpmS4Z8cIYeZfZgojgaFn+oSsEei5HbR3QNT/keOdibAm2LJ
Xf8DdR1xENgn8mYZAxibrB2lVY6WwTj6/Djk5V03kFx4qdif7pmkE/Nec6OK
zvw5mADE8Zme8jIQpyHg8AtkAI4bRWgZXbHyrfApemwaJdxbXLDe9YLB1VAP
PSYGTzOPoGz1n1GDK67Pkr8ozf7sBJ9hJ28BjFB1Oz1wF+H/DLBB1OCL4Ru+
9X+BvIC06PZyoLDj09kUyJ3BkPCQ4BoG3vdVGTbtoq/FM4YBdRFz3Azdee80
BsvKhAWyS2dHD+NcVn5Be/p5X1s+xfTahdngP0k44NUm9dyg+SvRGbueSrG3
C7dEHoXYJC3yT/tRnigWjSqFa3kUpyr8qi5gWn/Bb97qwRPAGeJDawcyWE4h
Usza88MqwNQIFE0eYgJ5YCtigKzqJM+dBXSgvgxey1klmKUKUocP1qyDVq2Q
S0vTuhHiV7hWCaZv+am3aBOVF8vl1pJDKPlkKwtu3jmB0mImPz3eKoVOOXce
GvcXlRPVw+kY1Mpz+3ndheUyO5JBC+mJdrGfVYVU+SVDm4xUb0zEEZCCID5r
SbURtcoxjD7Od9gpWt6Vdn9m94K8CrcZZUBx2lArA95UEEG7hsyEhlTTucsY
XYf6KerpSc+dPcIJvRYDZzpDYpsCjVmNtbGYJj2No2PryiOz3WWax4mBMq44
5/TsyGPky2UIaODptFfFAKWWX7jyHnB56QFqPV4h72tQsf9BN/wnj1gRh69T
vaOQ+HU6x2qeTnLoVLBc/4QfNmFQOi9d0sUa768IvjJT143aaDYpQDd8VQEk
0AyYm5wPJdzuPCQZLiG53xb8LUXi+c+cdpZJlq60Xfh2aV4lZbMv7CEuPJCG
MatjQe6aryKDGDOoaf734D6nkeiV8deafhj8GM24JYKJX1u6dPTCdrbrsMX7
ih8Mcn7eZsu+AEgLoLObcjMUpgP0NQ5sHH0eggtj8FVWLOclA/4YMGQf1CRS
rDmrOOlh4PEfZi9v4RtTv+JvYqpGS5VgP0UVPHp4w0PjpU+Tv2odL7+ZoJzo
nhxyALx4Fx3QvDtARKf6zCtLHDNeX9YeCV8t84N9sKy+BEMpyZV0KDtIrTk7
/dIPQhHIbR504nLrYBxBrAeH9fUQcCRoyBZjBDQtNRASHC3Tcar59tPZg0fc
0St3Rd08A7aMI+Qpwgou1JEqYeOFvdJYB7mwBVCSfNPLadJRpaUBCFjKxLGJ
jYihz6N8Lqsa94MhITWLyT99OfkOY5uo16BOI8l/SnTRRWJDi+QGgrt7wCGZ
FWCqQ0QkazJzK6nbWqISP56zEQ/bNYRx++bDlNG4AufACCQV6g/USrqK4Zzh
QfGeOsBeDUlv55sZ0raLmwAYC7aIfDLuOUqvV3eef5nqDlsAKKAeImcAge7s
OdTl4OscdeMufy0UdRTfXo3ne2uyTURV8/bkYoOlzebg36/iVTcZDtdMPxy3
8DudB+gx3Jj2YBrU3rTP0ksRqHAhqGe/A5TJCFWU4F/x4fLIwLW1Pi1+ATnD
lWo5rUYGUuh/TCd595E4+TZ804zlkZaQJ+eQ61GCVM7l1DRjvnmjHZqSkKbF
L71K1juBPmm/nbrl04LWDA11EkJ1GnjIlBdjlJwo3TLvNS34b2JIu3Z/4Spl
7hp6H/xWxMnlXKh2bxjjvrbd/vHtACerwVnCAQuvWn2S0PiBP6hcLNNfhb5g
6WYD8C2f+ybBHDFo9alpyjgZq13h31r0hS8uZQvUbQ999DLVY+6uU/3g6RRS
bW6yqAY2zdbvkMTSGa+yVmItB8zIKAaWx+BiIwz/BgKTNR9QxJv/KaV978wS
/BvZLcUg4zKi5UUvZByVR/Ro4um136ItlEpDScVRuYKP6ukdSf956U+WL2H8
RWjXxP23ay386Hb61nomsPQ9Xyyhrs9oBHp8z6FMW8H4+8YR1HTXtKz8PEUC
m0ZrB0GgA60FqvAFmXM+zf7ptME3/umIC7Ul1DC239svqC70FiO4X9vg8gvN
J/3jhpll1IlaDSHO9ok3DT10fPbzQbcfRsqfwybzYgZr1n6jiV1tS1U4occB
diuVt/I+9wcuCfLYqlho1jrJb3XWWe3T0QgEgGaqgaMLqNGeGDyDGEusr2Ds
G/GXFyGrWF2kiXwbaHZAOt8C72zXHQ2ktzXHFr3U+uAIERf+i1ZXEET9hsGQ
zpPpX+3OnMBsGh2ZmUdhy3+/leq1LvQWF+lhIP6Ay8Tm2ORoFZrzoxeiBrzz
KxGGt+ThPr4Yi69DuNEVrWp0f/PzEjJiwtu0jKFZ+eBTpyP0JaDXPYnMyGHF
WMuyn8jMxzm2XRW/a3Vww6nTaG+jZxgy1z3b2MynhRO8foJS0cixQubQnIlO
mgSpLH2+WXQyW3vBlPkkENFmir/KcrYqA2//I6GPCgtB1vbHYPsc19hzrrNm
cdhlJnj4LFb/IihQtluJvTfX9c8n5gKIrfBUqS88kOQLQPcPVIMfue2ZbSl4
/hyBPwqz7KiIV6JNn8Z/Y3P5QhtMYv8dLM3sJYWi8YbrYutPf0gms/fqjzE/
1hoVD2gVQ7E9qw2Tnf/m5WkQxZzYVkP3CwrNcT+kvvQM8MdonMzb65DIbMTT
WYyBEOatm6OFjW/sQGH8et/tWhfbrq/BElgnzg4Mx6ytJqkknnCgndD99db7
LN/y6rdLqSDp/Fio3ZIGHVs3e59xM+5KIlzx5vrx2PFQj0AILwCglLtlGjVr
gz1k5+TdwyF4P/2meJq/AWKHOyCzGUL3diQstTigFpeHoCclse45Sz7fn0DK
7NgdUTIoL/u32hMuUnKXUZWXaJOa+ZBKB/yeC0dM2tz6rXxyJRiJhmrPouAK
RbpOmj2GkKZPTDWBUdbrtpknBylfFETgy1kxO4TqWVRyV4lj7W1oUITr1SN3
aJvRqDV/lzIpy9Vo16l4XrWn9DXUB9z5UfUvVvVzVkvofWkS+fEafHhd9ubZ
8oE+cTxegfH+xUWeAl471dGO383ohEHkyX/zf2pg+98A3atrw4d9t404BJ0y
CmU1MUNo6i0JvVVS6Zszk/zCtguj3+4HlOY5xf/mLzZeu/MZYiTB782ymM9A
afBtHyURVHXvBzJOr+KPAjAI1y0+pP/ys9DS8w2Mr+LnNc6ao75ytZmBJ62V
vkQsTTx8aCQbrsaOMb8z5rNm4EOYYKixC3z+cEjQ6vAH4P2h9mKvRNacBq9X
tsiVGDcnMPr1ojqfcexgUQmGDzMz543WEQgenoRWXQWtlTlK+y47O0/4bfrb
M9JcFLHQAcoDLhJCNqAWsQE85NQKlanlx0VE7dx8v2VqnkgpkvCtgozXGGI4
pJcurlnAm2IMPDREp5PrpICMrOKnCZR2UaZbCJkyZPAMiutfbuvLR6Ut3782
zUbinl2DgP17WawLYWJYFtBIK8CY7pNU9n6YBtuB31Cw0EAVsSj72NoqX4zM
KFNJilUgNwoE5e8xNfGrUUqfoCaIMYj6rqZz/5WYwQQbYffpUsYyYtbja8IG
YHFqsYinUY/+Job7nBSkZ6EpyjyDJarfg8V5i7Zr13GpZeaazzx3YEWhdlhR
KInYbkm+2RDiOhN4FpZHvJgHGriq3E1XZ6HQfI6v6T4/NuMGvjYVrCn2w04N
C2DxWoFwFobAAsGtQmHGX0JR9HUkuevUoncXntcUeVVbrcoVNDA95L6PA7I1
ILhf2qRyImHd739Z/3R1/foYp3vY3XYuZIOkxz2KB08isDm7+7bwptD8zLJ4
8A7Iv68d5XyM/GaVNmzfIGhDEMPacurdHfCNvQ3/XZGDCeZDQ/rNE3VaoXkH
L+z1tZBGdgK4wCRARBz2Jsk15TOV4d5Qr/pflO0j9fG0o6XCWx33+dqJk12u
aRDimXHonuHmoTZwTdF4KRAtRhmXlkxg40WZ+Gbc4BC5N/bxgbEsgSYNtXQB
JMTrIpB50jdKwJTVfad32zB7gN+jRXcb0+Pg4J/rAFM9GEqgGxaEozWbgQQb
+AuuCqAp6aWvcpCQ8WjFkJgkC+EMNeArm1N7mB4jiqB3uOV9KHWf34DSb13q
4eNjEKwj+6xlnPcL2hti5nDM5t8mnZDTtvnK1UPBlZ2/2rSlakPHvPnRm5c4
PfFgULGznOZqSDYKg/aOq8h/qgSWtt6nVqgvnt1JztJObhLZDToEP28aeGVe
cWHnzW9DAONSKuE3XlfcGD2BmXvm8dfCS57wUCLfnC4A9lGv4rtRcFYAuDjo
aEvOIsHPKa69pedAZhv2EW/aaXo7/crM0jRJ9zua9u04PTzHtchr19jN1ovc
Kb2shF/vPyxxCeljePx2WcFkpSLr/w+ATDs0pdbhXMMy6MJsa+V9tP/wYzTh
D6ebueb8CIvYCjjTo4xH2VJoaENbjP2bxk7rqtusq3r11xOa51XUegC4/0n/
Y6EYDsqKmqk14e4GnucUrgXpyNszrOjtpkCGTLk9FY7XkGFmmoORSZ7PUTJM
+XTP15R/QRRSdwGIANp7iXVdP6KhKLAaHINQx1m+WLxuA7wz1Ken75B5fTdu
gVpz5O4Bw8sCnbZAGTAOgvNEbf5mr5iII4bB0hg1x/cctNpLN4oXSFfZ1KbB
tmIquE9129xoWm1+HeteE+PGo36l+PhOG/Z9O2ycGuW4WTM88In3rMKcVuch
Tbn5KfCg7Na6oRFfnhRpnS4SYYPR0CwUwd3vXEAZJG/T2RsX7HeOOCn6QG2B
OQ9ukX24cMKj/jInurEQ/45q1Btc4M5HI67mlycPIodRXSrXxbzzvULv6ICX
wyjMRX2dv0PfxNNcDMaDYw0ayPl0IStmvmb0sLlRtrqh4MEWXhiH6CmDru7g
TLV8MWRaum0t6zWH96oonS578WN7zVsmfkur6PR/RLThTzUU4QQyt+7OfYvE
5Mis0YpldNREAtAdvZoHMVE68hCnyQRHSkNAPFOSznoHlyIdqdGVuUH2/0g9
GvfIMRhaVEELsoJgL7vgSnwzRederx+iBM7FDq4eYZ+Evn2G0INg9yvmc7lc
69+HqZcG6/yQvGafIlJMraR7V6M4teP5IGueXmXmX3XY05BuN+1yh+ky3Da5
2THB2GvHTt3IZ3vB4G5AQh6Ewzd8Uht13ZD8gRYt/qOp54F6qsiVNJrypkT6
1dNIHVbVGYkqJYmgV0ZSXEbHbFQp8ih3kuHcjNWFxZuxeDLme6Emuvs6eZ4t
ETIzO44mGINA5xTl1Q2njgpQDhclNZeEKi89W31ERIdGGP5aB7KI/mmflOxr
ao/INHK+Y4omMLgG4zRE0bCQysU6qURk4F34H4X/Pc/aHya4G3IbTle1i12K
BDs0NuAN7QIJPH1BkFiAnLYsDsjJEK9K7YK9rokqyxrpPRcH4DItrbt+D/xg
+A8AwQnmPPuCJCEAImTJoBa9ZPfTJFkLbo78fS5o46e2ubK6g9mDwt4lld2R
xy2fEVupxcJ5Ti+gJg1d2LdbvUX2gHTx/BCeRJhoqEpvjZuvegjrN1FoFRbQ
IXOj+4hlwry3xj74lf0ER5szI4fU3JRZWBJpiZhWktT2QZoP2vbPBWtpiH88
rlsfE2sAPKAr0zxIbVpZWDHEur5ApEakj8jN1syuVL9EwIZfqKNzcfmzGFV0
AFhJKAVAhCpInSikPaiHgrAGD7CmYynasymJJdVG4lwqgj9pzdJgX6WEyKoL
TBMOCDuYa1syqeGpWPVp27q7yRuTLTTgxE1pSNGovzdPIj5PKfluEFU5J+zy
D5MkDbQP7ZYdbVoQfSglsgKVgZnNzmQ6Um6hyn5Xcec1K0wvlZwKCR9g/3le
oAIzg0whJIhHhkpNtKxtBi82SjuNHdMbVKcVAOvSOnBTr01g0nttFSDYIuoN
ppTJldwzvUj9UdHr1pJp98c3tVSgjAzZnZTKVoAhXFKnGZTX/xbYQ/sviINR
rybUUJoR4wGJKlgJMGbzL+rJ036c6qNSPIfqi2Y4Szs1KQA2rf+UwzjKBntZ
dfWf5K2NHtyDbJCj1KwLLj/V3HWoPU/Etj4v4m8Q46Ij4txcO7CXlgx18sc5
dIDioLtkRjA8GMEcpnyOXMyAWneKLCjr3l0A2MeCIxo4eHJpZo3v3ff3EMCs
UvQdZkd0F4Se1bXKVRzKvjMN4N5Gp1dTcFaqmliqkxswziA2bExISPo7ashu
Rle2Iy5Zrstsu49tjipoQz/ZGmHXFJ/VJwmGUjXBR2QNeKLOP9wsiE0yuZp/
iQMVVh8of7sXp31MiRdVO7kx5S+W82x4t4iHZW/ouzbu5Hn3nNLFp7YgwwzC
mkESavpm24+/+qt/1uqn9VzUePNDwkdsjtmGvOHwhNf4+2zxuEC39T/csAIo
1z3MT1IGJoTrP1+TM7uHtJ753n3qxTWu1G0jRFMZ6kB/AY7jh8Kt9PRy3j9s
8Kt/oXETZFVSabNe93X7C52c/klwiARwhIGcuR6wWKu+IU3qiY230wBi41+b
D8D8DxHin1C4gF8snILHnFxDKUD3XdDj6uGVqF+uwyES/H5RasqIb23+Uk1o
DtzOZgVPo+ApN3pPCA3OBfPD4TY6D//jKSCfxrwcfPz3CNjv8rnCdBmjg51M
GtQ5wmC4dZ/J505de9Rd+N7AxGwF6Go5kvmczNSnBLM1gGdVhJa+tFpyoDsG
ON5OJQy1jDxjAkGJYRB/8SBbrdWfqMAzU+Pbxg5R0m1KCc7dpdUPpL3N4Arr
yeONxgwRGLT7qZEsFLIRTW0fKL7mUH6uknq5UiMUSi4rxKJklqjird7aFK7Z
rAjr7j53WUroCM46Wsz8+BvMcmumuMeqrPj3zJ3RT8WLywXGeFWnPoJSW3Ti
wKW3jbv4cNsdNrEorfscQY/MUDODQqMkxE+n/AcDW43acn03Z7Q3SvBGeQqy
0vSFzert9uK1Wdcymwyq11qZc3GG7TZ8lwXNHHJZppDnmeePRN2EHJDXwZN1
VThB76LZqn06NIKVEeQnsXzom0Y4K3DufxdHTUU94en+8OsRicY53BbnUjzA
b7BrEi/CM75/ZWWeqQUIjIA/rpVZM7OXT6ZPXnh6qnYONUaGjOmP5j6HExIM
AJemhZ84af0zquim7yNNa6P8lg1NTXLFlI3j4T66lxRKifzxB20kztwbRsyd
fIPKOfKpfATnjXzUsfS8y/rT1ePQfoN410js/2RqpI40xy1XYfX7X0MkNDlG
5aPIIkv5pbE/HR8otFIHfiZnJe7z3loTdl0bRWA4uLa2VjOenlFUCCqamyA/
FcgGlftjULNMAAi4H9Ugl5Z21SW9RnK1WLTgAww5KxrWz4CETnJT7+6b1vNZ
mgoNHADSocXA1m62nmBxAet5cm8N+dovauVvlJMLlklXejzQeifVQkfVdYzN
tL8WCHMXrNu2En9PT/5/hedyrNhXTta7nJWH0vj/wVSYsHSWKj6L9aaK+5cy
K8p1s85W7oHjiFLtErsNlWzVEhhGJvU5BHc9L77NFmA9C+O1vZlBL3iDwvWd
wwFtEk07gUx9lzKE9zvLmc9/w7IEuXz0MWZri7kDIGGRnLjbZdDa/jTDcWbL
ByqLKV5oWPV0c/div/LB9b/mVZ04myynda7LF1N42HlaQJgJomkssgNYgmoT
P8D3G3Wtq7WXF40q8LCOd8xoXuklt0yTiu7LQoG52B6HKRuubZsAOUG84SIY
hU2803T4dx1v2B613fkk9uq9tfZGSj9GEzsrRcGgGJsvhXjgtuvvMJUEEQXq
Wd8/vsBjI+FtSefwAncltaL0LTiPXnnfvxXagaifpGV9r4O5k347sru2XppK
Mu9ePNvb5ky4r6zdn8Oe64CgSDKDV+flqUUCzuB2KADhohEAHVIyfSGEljq8
UO+hB82/wz2T9G2n2g/rj3JOVKyiImW+t3UpPk/AAYzsi0/G5eyHzltT4uPU
be6RB44fvSQenLb66cYjglctXfp7Yak2pglzAXoyY4kN2Ag2UiWtm/GSjr0c
YVu6/jR41MP2ve+KVsGq6rZqg6ScXo0VbhrThnB2JlbhdWY5FkI8CCKBXHiC
Pn23rlVZUCNoAnlZn8aWwBL6eG9aARmP9SvUCxtrx2xNO1h1DI4rWH92lW6G
eo6S+yCO+2e/IIGRKBmQq1UnwPJapdc2pmyAKHrpetA3nCBlrtjW402FZp1J
Cxt/CHPsYLv199Omzq4w5ypAn++AiqTAbc8XtVuGh+A5eKtXD8oatUEyfu8W
j1wj6UppGoZh3HgG9B9ltgb3TUOCotGjPpwduCMCroGs7mpN0Vt9etGBSMzC
RQfsxXKwkmWyEm3jkKEO1oUGhuB1OAgcxa0C68HHSgpSrwotG/mDQ1PRRdeq
FUw47MDwx7Q3Ax3LtXFedGdfHirauFRX3Ivhe4w6bhLC2KkfG2F0fucuqaCY
c8T5pqOnvyt391wvANgWzLmzgRURDUZvrE9i4z9GZ+ebetreeKX0mopKIkcj
bfL1x322Z/A82+i4BpkV73Dwfyinzi0pqvkeEzhiIFyqevHwCnFYrDd1NsX7
7ikwRWBXYwJQot9hIVP+CZT9Acj621z5YjDzt0It9K+lCAYscEgfLTV++g1d
Pf1Au4EivN3mcYxwUc/ES08ShYV9UuIpepCzta26NI9+In+jcZsLydbjVyCw
a1TTzgAYuq0Vu79DL4FDTB7h6TAuv5drShvpFgYC37uxKyqembyZZVyp1Nt/
LXuu20Xo4znQvwMvfvG7MfvGmi43+8sa7xCeygdG9gYhNMXD0gXLkAlOQSp0
MQ0xCzYk3mWx+t3iQVNKF3DBZrrrc+hcd0NiqHSfi2ac1tKhMgWiYL4bA1Co
3yMKFnaKFPW5jqy/GQ1I1mr7EqVMx15zl6HgHDASm0y3lmi1Gr1brv2UPhfS
dzdoWwaNFavRi8CGldmkSdASIAt3RMjKrgshDB8Sf1iz2FigD0PuHV6CA7cy
LadXzkhjb1l9wb+7t5axKDKyOJMzXQZgYuT60HywOI5tDAQzutmc7pUAtYbI
J5xUTe9jdmPrCVYKJkLHZDKML//Xpu5GXo7/5eOUV3Xwfawe/Q/qiIfsRWLG
OSCIniLT5limfZLLXDbxSoBevARR2KaB+cSlvlNNdFItBbNbDMYUMMTYkMUs
aXy4p0wDNKxcEM5HLEBPoRdF5tdZG5J0zwisiKvvpCyS9zOPbBU45U5n3T08
Xo11+n6wFHULlrnjlntC8XlOYozzBCahyHbbEDQKNc3kXdfqEa4BwYztAO4y
wIxKkkFP5h2EOsQWIkPW0s5fakXkHWNDd7rw/pLoEnrrTVGe83Raw3YBqBph
QNSGB7upguPG0CFuBbgu/kN4FWDbfqfWT5qql59RDqULdP8Gws4krBlbsmOp
WOLK6W2U+M5v0IxDkn8vfCn7eOmGqN8bntVHHi+uyvbm05vU9jn2sWXqHk44
E36C+q8iSnvxPDv0IjSvVb4HHA4jL5X5FK52kMvRdkwj0GWjClgZDsrl4Qej
iG6K5zrLVE/Z9VH+yl398DVOGIw1oAjg3n/hT857vq8MRZ0zrDmpb9+Dbpxf
Vfy5kuyJn2uQFeML3v0hXsM+FnJ7/Jc2PJX9gGfPmp8LIUkWnyT9CuUa/H7j
xMY5tKTnqzKQOYXkmXyWULHSVcOhZQje9ZyrtQKHLeYtkU6dG9OndDhIH6b2
AMEevUcR9D8YfQjZAkGGaDveA90mDc6sxsb8DsP9667VaBz5AgU2J8upqwpw
eUgldwA3syc56TVs1p9UudIqkZ8Q8i4J70eTW3WIIh3u5CEjGOhsd/Kx+4lw
ez34hbwkHfXwNLV0SPPnLuHi/uTuFcaHk/mOiBpKqyc/uoWsRyHZEleWK/mF
egqWpJGAo5NxruPjSbK1DCr3wnfZdHjhStTcWui0PEQYCpirpGExVTCi4S3x
vNhfPcE/NPA/N4bX2peweqKOeA5EIPiwi0KDaZuuvvHhsTGMhwBR9g435slV
Aovw+OOSbNoOopgXVf9zllGQdi1DKzsmWDxxXLcAVhTjc20nul7wtRzwrfwL
ErbqkdDfIKC60D+FMOdos2KHxolfPep9EemrUN873OHU8SQuXIP64LsdfUxM
mP4B1G5eLiNqXIwOS7ynhlU5Kx5mvo2stnSkajjHy9+T8d4pE0B+r1hCbR8S
DARtunBrlJ5sj869FKJKbXlPVrBCYWIrHAgyi95Srjc+NZVbR2282kHInW5d
WerIELAIxeLMW4N2vc9Ek1KS3EYKZhKTKtYON0cZm66AgLrd/HHHC4KNvl7l
T1if+R909Ol1y78n3PMFh7QXzYvzhHSV8Jm144qd4SLqTOkKgcTH5XOg05Y/
PU8aeaTki6XyBG7GYkjpHxGEuLR+MuJSSyxBzsxBfS5oiDaPo8mqttiHKOqL
qFJOlD+6ZyZIEPDrzbCjiVeAnUYr6MO1KKQLtWzmfs2tJZEPWh7yvwOEu5Yl
X+Q4WL8jZ+TEfGjdFCbCJnB+B+sl8tDCZtfeS7h+JPeK8xzshlfidzgBWkac
5+df3ERWu/n/v4dHhmM/QkuGU1Ru+Sy8wkyKkceuBt42JqjqvBhcVSFQwqE1
ZstI5pnMrDAhU5J8pGfh6akANxUYKgfKP7ipZpCIT43buNbwgxBxyF9w6I18
KaRCutarxVqsQR33GGxbjhmeaWeCXgTPMcRjVx3+ZIyluZX00LfYMSJPqISw
iVLmobORGc6gUTqERSb7UbL+dO0uDE1l8tH3JOV2OMIwB+YHb0g5qyF9hBky
yrYyG50INfRuXE36obI/h7cks1PLTwvnDyEedEhkDJ3IbHCeGlAVy0SJUdTG
NpErnyXWxwhGCUHYXjFiW55aHqLJdH1sk+PJyi7zzw3eZfPT+GEYlNpCMAO/
px5GzvTlPIEf+BuapdnmyibT3wh6FClZRurB+A8HDSxZXD412pmjXi3/2yA9
llD3xgZRmBbyZCE0/1BHClzQXcM7u1nzSThF+7hPXEiMNl2K6ArBsVM6knUz
ELXghr/hEgL0odk/v3eO1GctpzKMtq0Z4FJNed0oWs2HSmsD/11I0E4h7VXE
CfdjAm3qUOJxmESu1sO376SIcHnXLf3Cksh/HXmYu9acLbX4uA4mcYRqA592
klpu+yZUEjx0mgMVfXFdT9W/K7EinO7uYjRbq+VYuKCV/pseQAMIyBw4tqvD
n+JpREsHohd0lhVyhqD1C6/hW42ktT7KIuRajchFy9bqSZBpiZnSShT8IAOV
fHM7RK+VZ/6OiClyyG9AfVg+s9fLz/mZh2woas90TCo9K5/7MjbhwBBplyQ5
Yb1gUV5rAVnRBgL4OozHNbVjsl3t1F4Xm0hsICJN5ov2X6/djVPhV890IbvW
uJN1UuhBwaRGIrQdYpGKtGE3sMBWGptc2K2NKW+EtKfapmEDTbmpQsN7WGNg
JGfoyfDvGW+3SUXnpj7YIq9WeOBMunaO7uD2SjrS1NwvANBnDSOuv4MhTDbT
0n+nMW/OxwiEN5sxzhENVJbBwOMjyOAkKHkNaUvNxDEMdLW+vpi1lFfuIwLx
ZfHlePfx4DItEBw06RZULabOHZkusT23NCbkVxJ2AjWJFSwvmRKyVTVuaa5E
8h7qTptTmfDGaMrlC1jJLF7yxVKdnnaucIq0MTQK6/3oW2Wi3sXLOrqgEHRg
IgzcipoYvvrpGS5gKsA5wifNSwWDeMJcu3H6eXSxbIGkOsoU1d2nBLPhdLcx
FFlTqFAQPwpGoWsU08qxFvp53gNQvIT43eWoVjopijctd1jAf7gZC1eKpXWW
Z80T1orDicyExWrCwwsihWeEIvxQ3rImSH6Xq54ZX2VW6w1Pp4WjEBDyUBaN
2Q83EzbtMOkUzlXGZkI8XGdsETD2FLTCtVwQRr4ebLR0rQznMXAXvSKnpqjj
tDiUjLulLXpQsMWFHJX9jMh2S+LltQlq7MHENnwIfDz/YCCMuw75+0cjVN/3
zrPNvhNAZFn9HlK4nOzB3Xwqk2J7YaIkpBV7+jlFWcWLbDuePTVYujc3LEAB
f+Xp+/jmd3178WwVa0fAFazj4dAffc0fPvWfyP1piXnEj7vRJiQZjuu+CU3R
rXTZfxncjdsF9iPFhvBLHh7HxaplPk4jS5dtn6tAtfiRhjdBecp32BCt2l1N
6EP1aBs5yo9WoBee2bajplkg1EVMX/jURCGeT3tIwV2FrE1jxiLssWnakWI/
24yAV9sEZbzUsVyYOD5JFZUvb2+s4Q7vvKFgSNowjbg3n++4+2LIM4Ce+4Ie
hpE/IYh80XuBAmx+Ne28P3+kCDld6DF+wvTZ9+IDFH0ZMEaMF38tkF++CJdB
MjeabZKx9vtKU8MMdUmlJH0lKsFPnbTthvVsY+Hb0OwQl9uRR1yjNSGNmwOc
fn4JncgOrI7oHT3Px+TeBSdUafh5WtT+NgucP/AI5c63228QxIwwcHMeYyKB
qouMF2BtK2Ohusw3zUPtDBvsz4Wwad74TOyvmqJrG6CtCqo9DCUvlIsC2EAK
Qgpd1I11AvK2C+ihmf2H8nE/USWQz9EA3V4KyrLzHUj9vAZk1GP9cCTeOYsn
Tk8/a2xTJMM6r5Oggu4kdxnOLHrxN8fYQQ/KPB8z1eOhL6H8f/XF1GNZ+S2b
1swgo1w3+4PiaIBk8EGDSLNQED+tk5uzTGu0U/iukluLIu4NfO/yNkF55n2y
21CV9YXF09qT2SQDECW6wR8mt3fRBcU7vUG+60C/L4IaQpBzFDO+vdJUK68T
xd5S4lc0gdjSb6w7UiwsPG+xUZza+wZJhF5z5hVKpLsTGUtZpErxUzuQxtEY
IQ6iyV3GXhTmEyTCj2TSNRqnvjoy+ZWNCnBnFEZ40zPIl/rEq23qwe08hnoX
6bKbrrC4yu7uIuTm2skqmxIlh/uDoIIEolMYM9eAlP+vIIXYCz3JIltzgibs
g3a0gvBVdnTlRj9r6Pqka1+yh1iHRwmqnSAcSofIR7nQLv+r/0Or6yXYl2rV
MRnpDV6gY5iHRv0Fn4hnhTT0weB7aRJz9zOg+PDZKniC/47eJI7KZF5VJ7JA
HeC1m5nbNFURJ4E/obuppm6X5GDngB0RVmjRQ/DssFG/OiVcOtm2c9u4pcv7
0gpoj3ARo7qYRUze3RF34MRvYvarz/AEP5s6+Guds5aONEEEGnvOMDA8LFTd
LFGF9xMQvzVPF0ckC5NYjeI8+QrXkSjOyXsqJTbSnV7VSX5O58BVul0RtQe5
Idpk4PnYOcVAKs+iZJQuPvbVpIIb0CkYRzOdXfo5v4XKY1XHd5oRk7eDJ209
Hpm+lOqi1VOCTUdDwsrAekze2aDvhelix92tl/mLF6KhxLQyCST4ox4eKrWv
5MZtoYWLTmeoXHNRbYwdoXimW2ZLzbqoxTv1BKiexZRCEMy45fQChCCMF90h
IptxxiMZkzDIA2Z1+ZKJaB013yW6U/rledoWx83aaMqB9vqJl1kov1V1ViLX
aawVhdoGl9KWKMQRyRcjRXqWjgOkKITKau8kXOBJFsH19rAruNVsZbpO/PSl
rYPux1W65pvTtODb3FVdqtOUl3UujAyzGnVoDqygW9v99SmChSlr5aSs+WWT
o707bsFTBXQq4CAgPdXzL4BaV6gSiWD1d2MqP7idYG/PEeURiSkgszpu0GVZ
gDEhYXo1gMTOVQPDNvX+cQ62C7/vOY49TJqI44als3uaJTl//YtFB9fgdE78
RUCGlQtaAYjVLeGi1kc9QM4It6eqqmveDyNVX0Cx0Rcqrm6RuYmEsNqUeThh
bcF5L6Kic1utiZWD4STd6DXHECrSM3p54+e+wl5jhjVRLr7vGar9sBydU7Xw
lZgAMwk0mja4RAtKu2qv0oXTgFLGN2tfCDeQhldklwOJpfHTu+14lW4T+D6+
tyFsQmxDaIh8EiYCoO2ja+PviODntBBQT1PREZ04oUgVt9w548zPH39tYt3P
fuef1MWotD5fZDF8bsXLvI5q1XExZbdX6YApAiBAvQEVsGhb2NNSc9x58kOo
7Mki/+qMtXJOClh8UAKoAFjyyAg1bsCJBtI+mK5X0WHf7BcnMXjGMmJMqJvl
mJDC6oy1c8rzo+s+0/0BX7QdBikTuCL7i136fLH/b6s6p66DMvlGA8zQknqB
yw/ckk3cV28WGe3OmXbJjdHDj1/5c9lqB1QNUjX1hTXEOkopp0f9MKp8kcOI
o0sQ4TRcQ0DdyW2RSqFPeUBiLKlHhP8mh0/8UbIy5f/ORWXk5n3IxtE/aHTC
aRQK5KF0M4/K8sA5V5cj18SuGnbibLiNBy3AbdXaDb7jdT32Zlc3jR+Vv7A1
4QTS9YDGDT3NnfSUzxtji7s/NMZMcleS6H8z5zcr68f3SiVDUbI+i+LWs/ht
l6UZtp9MLmuRfA7YkEpI4Cs6vgQsw3RTbH+ZUF5B3iOZJiV8T2ELIQZqOKTy
lIy9dXNDhlf5GQbhk6tuTJVbtK43MGqyIGHMiDA3Ieu1dsUOLtCGEgqZtBB6
mbQWxupyPXAk6wynN+NKLqxzDCfKUVkk0dgezXZll2tBdvHsPWRAJsaVV+VB
SxEeUw17P+PXSr4dVSppPqeaSXhVQhcl0PRxNXjS99jRa985evX534ZMiZL3
6/Sbg8lpAh3+k1EimhfYUzDPZQ/bUJxA04l4edc954uJDJ4XqcH5Qlnip31t
19ihNxGSxvnNGZx3GmTcrYASk79EGZKo05TYzrKOrJFMtX2/10/4nnwWjM7W
WMkRWGoP395sG+5XqOP+2WleQ1bTd4cFJ+1rCoxE5fV67YJI0OO5yHn3rcUp
2eEm9YTrW8Abq/rVD559QY92rVDbxGV0Oc62ZBLCvfLaOrZkjax6UPTqG0qN
qUZrev7njBMZF5xB5rLPRP+c/gKfG7xUWdkJBZrTAMnzEOGnrU5WVj4JfRWi
SzNqlEXISYOG4moGIwd26S/BQqmZUGPtyiGHNTeoy7nEbjHm1K6+vL4ufSvD
juvfCTbmxjCLD6mueRbolaG3J94q0DJCk9csyhOPzYe2oECvBT9yBMqANHoa
9wSRMW3A8656R8/Q4k6RUHqoyX3XRMZjeKGjJvEFK5YyDKC/g2dPk2VssPAU
SaHsNJYNMVFArPmxySouJAn5uUW4726r3UYaYbUbpMC6s9BqQETrLaJl1Gv3
xkeQsz0GdHWhYvsZbsmgQzzYqvdc+evj8aSiA34y2B3BPJLsTZgNNb006Q9j
hDQlfXDwPzlFfZvY0AolFM4PHM5MbteBffwvzO4UwzoCb3ObL2rDomEJUE4p
Hsd13mmTaAtxXLFtbQ/sOGR8hZ0GwMYOEEP62ti3W9oWfTqAEWuNp8Ek/im+
ykvAyXm16PQCTUwxnCMuwVFJi/nMN64iIqN+HL9z/+g4ho+BD7GCVlPc8KoK
+Qm8jxyDeRrqyro4UAS4mCJF9G3QTirTQmb3vlLVpnmkcH8THsV3yeW7mxXr
18Y9cMIwU7JcEGXa3RqRRijFrA+gFbXvpcP6EcfItG6FC+Js11GjojxxRXbb
W8+VsRUKvLRssjs+Fb/Y2HqYf1aKxzyblgmFS2fDb9KDh29CaTvcgxW20EUL
7BgyTc/Rt/nBhmJwUbmfGyIi7yLrIGgtfw/YsSpoBzYx1bUrlg8WJf5u0Zme
wVsOa6IjW/2nUIOEOvgGNE3+dH6Xh1tPIUyHsVk6YoayNatqHQaHXPnEkgaN
6gNBzbGgF+pwL5lBKBfi40w6SuJl8SnlNCsqpDAejdsHpRObN2yWLh9ob6Qe
Tl/ERjcoCzlaGQ5QVBN7Ik3ybHvV8GkoH+IHcDCODBS/CYGVQgiJW+P0UDte
QWui8FhH4KwmRF7lDSTMopHOJ5pWEElhcAx7qHW7mOsevV7Y786kkf0pdILo
mrw7M2ja0QQO8Z58dLQXX0gBv5s7Jge3hwlJwOqHIOvVLK8tLYn9hGgIeoA+
WGabjNc7/Wi+glmWBWmq740aBrZJu5Ckkbaml5zRY2ErPAZuBuSVy+iZfzG9
oFrvA+nMgrwfX6LnpX4VX+Wo4brdFVy/PtTgM4vGVZUj8F4vidx9yRkKqgIm
P65DFW6dujhhLi/KcYwSCEsI+ZyBlFzXUl5n99coBAijM1TslAGCKQ8R2yZS
CaDjT0fUyDIA6k2n4rJ4RsdST9vOj9QoiyGPM63v2TL83dn/dN/8fGQwbgna
Dhgu1GA7X6A9GqjFVBRpO+Vl2Wi4IdMU/eLE9XmIV3BqOpdN7icOiQYESKAh
7tLsJRmV8gCsV78v/BblE1dDOCbIvwFkXg4R2/EIW84+0fBgVJJCsUeCukFN
W+aJRzEjy2C6JSYw0jgv3UtevL313zDF3BYkaCqk5k2Q+Gl/bodOdxf+RK5+
swFGvrpwUYfZSv417q7c60DtFw3V64JY7AH9iCJJFC69mdeeKu1esDmk/WWq
kcRVsrbS7CtLETinPLr2b4UzhjxKaYOFTcf1fkUYrHDfrC/tEKrDFMLENgK/
yLH1NYFkmjLCQkftzf3w6PxT+eT/Aac53buwalP8gxp7nQN4P86HZG3WtvDP
o397d8oB4gZwFJzWydFitP25pp4qNsFFRuOT2Qn0pYQEZsn0z7Zp3Nnr37nk
GzO2ohyUAcRxeIpUsZo6e7GYhYZkLj2VchF9Gu8x0nWcuDpUdCvVlxAS3kJP
coXWUzc9cLCo9FXj8AWCuIj0j8uabeC3CJp4E5arBGu7LC/X6jZAUWHJHLGH
WgFmKn0iC4mNPlTgSwhviOg5ZVaj3Ocp8PSn3uCXGZvbcggui7SFKvzXHvPZ
IneUqBqxu24p07V6os6/0W3DSq6G4K9chJyGfNYW9AgH7PDbcnjik34Pdnsp
cL0SKt9Wm+rWfukqcPlmygB1xROvbYA8IgFb43377KashMUDuxcduWe9cBK3
h00xuQhCFM/0ivu7LZTRcdP+UiXrYsMj08eNt2z68decJFf/y1lAjTzeLzoK
H+8LLvnZ0Wgw407oWuyL/OkYleEvMU67rWQWE8AlfKz4x55F6hPvBzbJOx27
CuQO9CZHPF7TIdOXnDRbSDPNYWHjT80lOIR0575ru2uo2e7gcz+nxId/HR6U
iw3BfAvL6Mo208PLT04KftDMXqCFwx+MgOYfW9EQKfARfAyWGxqXsYLIIUdI
ImeC7v4GCRkueZ5JcG/FWQ7X6KzBir75Z79m+a0nzRozJGQfY/QIU+T4otQp
oKI0mtHve5KCFc+RhhgzJCuO7pUwX9/Hw0ikP8IMxvHaaw/sqnDgxYa2vsKf
lwHAezdLgmwLSuBdqf+zgYIc3rN6iv2XVDTnyoSExaIRH9pKiaS3MgIs0KAO
uHGNCuTCjMjH8u3HVDkCOaLlXKhDhzTqoh35X2KR2AdD5Z2H1c7tIvWFu8hP
MjlwDy+4WGF5SbeeFgPfyjKZE6mJ4ZSkBjq9GuC0CoUZk7+JGjuID0MpPVdl
nca1frad5bwATfT8UB8xiD545WO23XgI4NK6JWms4Mr7F4jCw90z87tlRV1T
Fc9Jov+1TCjFiqLbUagLWEDTMQM8b4fmS0Gc4e2zNu4YLtlL/fXVjzjPeRVF
F1zpa3t5JhoKgu3CbWIbuJKr7QYO5wp9gEN3G9IAOZEZz6dmx9vaokGBdNUY
MzLSM+d8hWmS3ZkUisZpSkoaV0JsXeZAOg4BIY2e62Db64PVU5NTsErno1iZ
WhWoTdFfMeDo4iKULKJTBT5+MzaqeuYXCUWGm4xvv/bpPBXlTZ+fSRXK8HBA
rOYJanJBxdMBgye9fJPwoRQw+iuZIYVXQSptXJv5IPE7hsvgcp00qHS8jAp3
ySy1Ooh/mHyPieDp83Y9mtcr5OuOAhYiuQBiXruxQ9FZNxE2Ak9WeGNu9yHE
PtgW9+JRMExsbxHPzJzqFW8HIK2LCJgkb9CZW74ifIzpcIdle77mlYLKtB0V
J1MsGwVO0pLpfT/Rgn4ko+tulCnBZt9PL+BIl7+d12RshPyitjlfEj+uCqTQ
jbZkmFbpbOSvSxdQwg8g+xZnSBgM/zSPJZhqcr+CAxqFaDO8sE3ds4LPEt+Q
7c6vPQKaaEUh38F4wdd0glgvB9qSk3FhR0P//4DB1NPaBgh2EvBPA0OXcEBb
CG19w7y2aYX0Nx+sQNLdxE08ZaR8Ksa8gkYg+nxvhNj94Uq0ndKCAu2YsIy7
ardIPrPSC3UsDmlktc3blZlW3j3I5YV/hdp72UYKWRpXU9VM8Q3pjNsTWoLn
j0kQdo5bRUPpLAzRpmDUbGH97DdPO0uS10OLPoLyDr+H1x3TmTWLkN7qx4dq
jsubxzp06luAZCs0OR35w/+jjer8cO0ICqyIR++O8RUxGNro5LqyB7IMfa5f
GWKXfx5OKdTnKgLX8jxSBAefU673Rvt3OrCrF8dTb8vOErccQHj1XT7vN2LT
MrE5G55ePyZ/MoU71ArRAhpftaQiUniGRm/tFfQQR+PSEgDeaABw6jbwOvio
nxbLUuRRAgrcx/Jf6FeudqJb+c5Y+QJkM4Dkwv+jB6aAeYDvIEF2gsWCchth
eyf4GpXhRUwKZi7GJX6oG88Xq9afZ/oeT2UPvBIFasBbFb4UDaNC1PDKqZ2I
7QlgH4Zb9ZNpKP7etIWi1CiiOqL8RtqyosgkcvtA6wFhiX9Ibefmx3+VbbkE
N/6vh+JnCYYiC9XRLfQ11xk7i8cBWLEwJ6kdImZAoJfsPLm4/ZW1S5HQ67lt
yQxVJY3aPzXdAWeow+V+ILhnWZWUVE0kveO3ZGDDFual4q7zaTZZN925SYME
3x39xKfsKbT+xT2zzd0wcoe+Of4ln5b1LuUjTPc0PTygJy4lsYGwtY0ilZZE
oka5KQuG5mjsAYH6rhwQ2sWcBUXtWb0McjoCZ5Gd9CURKpDP1sIqC7T501ED
59fPnppLbMLqqoRkPUb1ivJwJ8cwTXd0gVb7CDADAm3jmkCk9KnFdRyollZ3
VBwocRLq4hzQRDNkJm2HCWiOD0muaFzI6DoLWALohi4+C9wfjU+D8qlYW959
NV8LFi0TuOB95bngCB0Dir6Yo51/aHlJRYYRcXfHfZtcnxZWikpXaQzsT3rw
T8ajaPrgi1YzdZkGlsYWuGRXbR+IGPNn+CDiOM8jQTPXatA5Y+bM8xsmRDX2
fbpn570N9WS52Oi9pwwvw66aQ6L8P6JCxsZg7adgf3Dx0wI7Vgkvw1eFdat9
z+EvwC7v6VLNNs3R88I6+29P5bz+mNmJvYKVq6VJETo91u6Bm6Qa63G7FcRZ
VQyArNFASqYLhfY0u/qc0AHjEbiUqAPH6hIn0Z62OCNbJlMzOTh2d8KbU18W
bLIjsYRYD3Huc+jUGwMvOfyupF2w3JL73ga1y0CRYLtJBn1IWnRVgUApLByV
uODpI5Q6tyOWD4ax/XtTNcZXw5MyhUAwihVRaCCdNuuIuGa/P8UYvOb/VG4R
qUue80dnwuU9UsHwk0sCBAP3O8qdnuqIEXQeV+rlYlSsmlbxQh2AaJ+YRrod
K9WLAAHYvu1gCmRFhO7fnQ6bgNR3N4yaGHW3UzwZ/Al9IzLSlNdXdaSO2AWp
nfEcLNhS8GXF1wOfJfQl7lKUaYbyEqTMJS6ujWqD2Y1Z1q7veARX95/ozx4R
Zf+sk/BrCFj9OeuT/OATl3AvuF7Epx7zvTbriuu3jH9lxbOL0sMDoa0vKqSK
ztUgZ/7v/6JqFSDIlKf3nm95xUInBEhF7HalBjs+RfKjXEn76JY0m6BSHUP7
k08uSI/MIuL+Y+TAw7LX2aFlLMuBSjdeiSNNjeFS7OQjGyPEnrUmA0JFsEUV
qRDwmAk2saaVrDiUTH78WjTbCRQUPSsRYJWg6ZB3COeOA2nv2Ha+s/R3svUN
yPCzCpWRr9xVtZKVlu6XHt6EtXrk9GF7giJr51tKgDj04zaT8pKocV4U0+k7
/Pzu0Xm94axMWKkRtDrCelJQOKnmcpBif7jgneLGXrzKBdS6F4+kzzJr0D4r
2+iZ1/ccTy394aeB1jcKKK6xVHG5M+gbZ9W5z404kxFfBDjGcIhCComd5lgO
5/rn2IxY1VTYY6ddU2xE9optVYBQ7DTyNdeAjFJ6OAvKxIYi70u7tpjn8fWJ
kTqncKxKXOOLBqFoeE2soJHgcNQDaz/JEW7Sd/St53FI4WaADj7WYoguTq86
eOoYIKd37WVuLszsyBIW5DX04/ThqoiXzSo1FA9lUk69AhhbqiDXQxcFpk7k
t5Tcm0eau8pHyE74EIuIsxmg2JWX00IiHhOunE3SAPr2gDnUovDjWEq6Go6g
U6DYMu6Jv+W3hrjnii8GNND0cvtCezc3pgmjODR5SNNLT62mKZ4VC258Ttd6
XzlSzR7ULp6tIDcbyxWX6CozuX2VPFeK+uKrSByDar59p9xcHng0xRH/9ARJ
qfNhaZG2QarFO8H8PMW9+7P1rRPl2raiA67PDc75U82Nzbih1XbCNVekVPwM
MZ7VCwuZBjtqB48vdMI5y5nrc2B8KRjmCDZrGxK860k4ptWRA341GWall1SM
R2BfIst2+9LdUzBz7j0cDiFlnv5NmnwjjxC/vdzI0Ie5pc9bsNofbz7uVN97
zOBcFRH0HJOEUuus1M3kButIWvjBgm+3O2S/tQeTeBH5JOsIVElyCYm+tLyM
QsDr1dTnnM0iHvZBaU+uwkAiyDfUAexzn5PCnphtHGcEXzk3wL8M5dWizLqe
02wSxf5Nwi7H3B2auvQln5kBJm/+5P6/oVG/DGWX8kgoShSWG/LlNOjU8wTO
apZltIU2GbzqI2Qnhk6s+LxZxAMCY6Psgn871GOe1vUrJ4SvVA4kimrEAUEA
E50FukYRs/flPK1Rpth76lCsFO2g+1Sa9M45lRvJ0APbaKpyFmf8iJCJqkSN
EQmrRJEs6UZjNEO3o/sgMAGR/X7X6s2WylDoI3SWLfJL8CWIiPi6QfkXkepa
J4lXkTaLzSgAtRmUOXAqZUNE2a9LiYIwcHPTgOY/PnJGg53DFhiJeEnud7No
G4jMYrwuHrrVP20h9M3k7ytIEs7rg+uEvSvVheYPE8P43gvGohfpgv14Y6EW
DtUFG/g4rg8xmUba9n6dV3bFVieQaBNNCohRvFOc7Fr4uaDIggQ4I/bKBHEi
hT8YMP1qdorUnGJpwppcmKVol6UjVlFxy3iuw4oj0QmCF/WJABe5jFykZo58
2XbAH1dlTQUe5CDtFktToGxmRi3lYo9GH0vKPA6cDot3UmX8xuFOlceC1NMZ
GAMccUv1O3HjVxk8uRzSy6vBH1aFxiaEXfbI334NbC9WCjv0NZU78Yk4m6uh
ym0rriVVGwtl6xJwLLhPznH6KBYD2G2U4s9X2WzONL/VHXkJ4YTJ+j9qjmpW
BGILNJ+M9rAjP12BADauE5YGC/PBmjmfa/EscClCVjDh9RarFZcwt7IA+ek2
IROqaCgqNTJlUGKrrw689XYh5lAMCyHo5UkmqZGY45hBeVUxzxIEyhZW88QW
d1Ce/FoiOz4bsctrYx6B3kSUsFJZO2Ipq/g9cGd93+ZFlEZXGlkeZgwiJMoC
RGo8yo+GCE32XaO/yrTDip9mpQ479NlIU6LCZcwzilYmuWWTWrnFqtNFgikH
I/5IHYSvgzeOEWEnDtMko6OsWNOodphKmASfH74iyGfPjvoB7ifv4nAf3p9w
GX5CUZB5MXrPjExjxg3pPpnIHKpOdsn6oYbaN0hhlfMk6CVMZ4OJ1Akrjg+A
6SfTYd2frAPcY1o9txek7F8mqjAADof1W/8Bm14AeR5XNtE+O+9qmd/pjOEH
65SvaxCj9tPKm2LDghd13oK2VhbCtXM+3vfAK/rzkjSFGSfAUmQM68q5Iw1o
K16zFa16x0+q6iwDMpXDbzTQ2gmamy7XcYur/cLIiusPwosHo21xT4AvuGLs
TkgkW58n2qNBhZpkl/LBQeJrY+1bllI+AMgpDPCgBG3nzdAzMpgZTIdFi7Db
4C8K0tBNutQVa66GrocFRr+4pwfbEJoJv/fGU+O+Jp0Aw0rvXk+S6cJ1ogtD
c8iKFIbXTNjpVsa/xqFF0H5BcNjAIgUFruIbno9qagpojsA3ummXi/PJePgq
Uotz7qiP0alFPNr4o7lNihTw1JvjxfnKqgKhHS1jOgXCYDui9otYT7VcwEv0
yHz49nkRs1zprkIM20y2/H9CFJavrPLmDfhS0JxPQZ//Wl7ETPGjUP6aalh0
Yf5rsuLdArEkxbYPJbSGNmgrYRUBFBljA7xAWlCOdGgaOQA1+djGScViOeYb
gLxoWXR3ZyIq5zCHz+ibIzaQURJ1v1fDEHQqF0XIbl7/+0rOzFGqUsdDBEla
Umu9TDm8tM+hlsByU0Y5rDX7kbIYH3kDPTaQ2TVSfYblp01lUI2dOLmlLBwC
YZDXC94/hMgRMqF9n7jeI0np7VZbiBtuI2zJTk3MRm+KEi5CrGImPKRuDHvr
BiXUN5isAN1ML2VBXY+GF9Yn1Uq+YfuTJnSYPyYHQ+NhOr1Tr2YvL2qQUMNQ
221gnCN3BudscvotGC5+Z5bTS1/ihHymzRAJm59ZNA3zAHF4O1+afv495Roe
CZCx1OXZyLk7QeE9kVAc8DCgmRQ3c6tb/BHU7AiyUapDhQKrW2kzKrVe4nNO
peQZol06xwDXmA9aI6Xf4GakCZYlxqgT/QK5IlPmlA71DOFOWbhWHk44wiqR
QxUvTmwrwjXFl/2CiCiTFadZIh4VC3uwgf/0H/iSdOLSORyCeLP1H1knSlh+
dG7sSNnaaxlZ0me2dNs81sf2LH5dcqKvJfAIh3s/xnHW7Aekdp4iJYdCsgGi
q9NcWsicDWjvEiQXFnUZ19bD+t5w7olnzkQrYyB0TuXB+7ggf2OZbG6d7aYs
RoyWFEPeOIYKyH8ue6hdC6Pv7da3bExuMs05o99qnfQPPS60AETogIk6NrAh
mYINhmQUYoVJw3DRURNYkAOem7GGsWSPgShqnf/RPZ4iL1aZU57suHubp+xf
tEsXidGBca+skES8c3+Z3b1acwVnJyWMum8KuwVV5UdM2e0XS2edz1ud3peg
7RzZacEsI+VtPDOgmOj8pMQWBrlS3OPNMVAiG81fdYAZqlYUCgAStvqCG9Tv
raStPlW/JcSvwxJC3DRmhJ3lzK3E29KdY/cTCnyPrYGu7LfOugfb8zxFD8Cs
wREL/wKqrVA89Ck+TkAdpgA4QKijUpNKI85/AR+dakAvoaF1EAnsEJvJibzL
X3PUMCl8Ntqy3Ld1dCbvRZfjMB0Js/Nr1vEre8hkCDGtnl8Y8/nhc5A4ugW3
SazFR5DmB8d4Aqj82ycsddgoVRT6T6P5b63MP7ImgC+deOkGW6oRG+riteSl
BHaF5MGZt9lhanjdWvndZIDS3Q0NehGUwVsIyqrWwx+TBKYgGugddj3QK6yc
iDn7s/1m7TN37X9q1VBnn5dKPQYccvTOJ8BqYMFbRwEnfWIMhi5b83EaS6cr
x8UrExXo+qHIGipWQaM30sW3iBr9gdDlal/cB8sOK7AG+UlwNcHtR4IMUiQS
gFKU8ZEpaPUZl5WotTQZkfFssGUHmDgI/pE3foRo0UglpIAd6bsrMmwKLi82
PEALRRJgfZlruW2TVRdTLvjQPLluta/wGyDE8uNzBCeXOhS8gHoWVUSTVTp2
7WCd4P/UmU9XX9FySDptvZgCEnafqkXZgzhg+gUMb7CoiwnvtLIy1fTWPjpv
uOMKbnELxPdHo2nsnjw0zeX5hlMfK8zVAlTCHcIYsMjZXW3Sql/LZj5u4XVF
jw3WfRH59EyCMqyi+G1lbeMA6S/fPHWOhCuZ3QZdFye2BPFkaYSSiu/sikn3
2rmMvJdcJn8720fJ/PKE960FZOpTloG7QRYpT0x6qnukdSTEtuoTcgndvaEn
B5uZrVSM2TMYIMQVcN5HNH8y/+sUJ1YJwUZfxDDcNTM62wU6UtraGL8xvlh1
oW/wLkZFY3w7H6hCilWz3ehICbvN0FBAPgfddTzeQJhMcceOA2OtZC3Nm0WI
m5E7nfNOZwhY9VAiD7BScWaaJLMz8zmu0OptF/etxxu2pTJcSjhYRI2GpOv+
CBgGkcy9Sz/whwp0wfsl3EBEph67785MBkjWTW3MskzptfxinrC1dU2Vo4p6
VpV+aH7PBnD9LTZHnrOtOV6IMMT6Qxq6S240R74M0r0UJfOYlxwDBu07WRBO
pIJHJs5kAwb0e3fhn9Rlh0aOEDfISEC1OkV4ZR0sgVeoasrrm/XpPmy7bBTS
7Lp1KAM53SRYYnMWijCxPCvhPhBt3Owmwzk2Yv7rxtH8jhaheeLD56x4pshY
u4AkCzSI+Aicu96HYQk6h5Idpm3EcMzwo2sDNjBv1N6tGIUxyRHhplfp6Mi4
q3apAq1N4IdudRMaAnQses3QlsJOAGwEzbrOxe+Z1Rp/C4wz3U1iRAIaOLg8
mTAo9wE3D3W8yPCA6Gexvke3nj2DtRbcVoWTfvkRpfbKzbqkCJQ+Y8GYbtzW
zmKQJqlg2ag6M25aOuo58CgGsBgGxz9mpXbuhClYoHbqoVaNBYE6FkgbsV7t
ghnImSDZa/a1NJHRWhz+cXYgi5A23vTuixeZJwEfZUvUJe3mLOwXxB6Vccan
cEO1SXJoZggHBVf5MCPD6MRKIpD8Hs7xeJlqNJQa0t7lu74X5utHqQZjyQ6k
MWmlWXnA3DLwh/Hu5rFFYyzkAp0jZMJFtswSZAEWaWnaKkK9qdcEzK8KDSK7
qp6PS9yp+2XqefvYESnqwJ7by9ueTLVQC6VHVHJDqOGOlZZG2lToApBSYUsm
32Gs3slFEhZI4jQXfKxDKb9sCeEdmWeZSTWZf+8lCCTqHZd1op6ZJOKqAIiP
HqAfO9tSvou4taR/XaiBeuY7MJf4fu3AlAYC+Lflvr6ntgNVOvdWhPVndkZR
5C5mLzs0DszkVgmnv6/U4qvP1t9+uOFSwYeeU6wO6aLPkNDVYFHozZiWlzW4
3va1f6+S0My7ty1tmWGpfZlOMpBaOJR146TmYSB6EJ9N3oyDXddu2wN9mo7I
INtvgXZWPxhrWpJ7vstRWnI4rBm+H+rOYJrngdcZ1OfN6exsgCcPHpLRxcFu
ikASRuY1wF0R1zWdPNk7zBqJA6hx4o8nL6qqE5A2ZiP0dDs56eSdDaY+WmPR
M1cYqAdqkTdA8BcMnA6dC8LAFcvDd1gQR8f7TvRpJnYL4ix6Q+JW4q/px+Ar
XAZBFLrSiBa0YBzMkhWd2L7+du5K14ihzOAsTycyhmMHBASp0V0PpSWZOBvB
+Ql1LQFQp9/U6mZ8Y1oX7dnHDZfNER9bm5TYTOTYbJDYlQF1tbTvw+yi72z2
u7H9xHljZKhpb+I2FOCMUCif3f4QlF1D82Iwj7B/c1ko1md3gmOK7Q90GakQ
/0WLhwXUqDCiMvHv44UsoHMGqq8P3PjdAwyHXvg10CDfVHovUNjxH+J7KytX
/SrQuMCZFblUCd4lB25JYE/Zq889obvfk9MkTcEndgXWU+9Yuq7lNmpRAFoq
eRFDcBbTgq6yFvPAqA/8f1jNMNZuEIzRW1fMXinMpj0wmYVCf127G78Vb0BY
EW4DI4w61Fn//kyMUrGNpTBYwWqPvSDhS19z+QEZHRkVsIxZvS1leLhGMQLC
E3Zbrs6aBrRY4XeyD35shNnP1EmkqUDrSEJhRCh4vJcpZq8fJhP5Zkwlfcjv
wKUXpUx7Sx/hC6XIosV1zjs+0w9tEOMcv9lE+8+P7t8ATPkoioJ1d08IHqXx
IjIX1u/i/75w5SreKm4+44WnAzUmSVfobo8x6/Yjv/B16NH+RxHwh85Pe3pi
iib8VxVYPKJU7f+T1w4J+wsdqeUXr0eBrcwJs0YkpIXgxgHtyk+a1odPKwzm
sXU9WsTcUAax9XBnDTrTFQmok0wQ7lwXceXvBpy7I6eHNhkHXuDw6p3NDoTd
Vd/Q+wK48Qt44eqhjh8rJbkwsj2sh8arJ4TaClOqWu6QvGpJQLm0KZmzWS4u
90u8ph4oyJJrz6Yg7pIfk67KBYPdj5S6gv8KbDCSVGLnKLrZHiVk4lCmZdhp
4RIimPN2FnG5i2aFR5IpB1NlSnB9/14SSC2NBU+8aM+n7hHeIBUDUPH3PmXR
FCV+7X1+QzBGB8zZP+37LjOm1vVPXgtuJ0FdXQIfxuW9cJEMePIfo846//X2
JF0+W+6phvGFtR1+Ks3FoyWOo1m863ZiGv7FKZxg5QTUGTE67hPjtIYLah/c
MNTndOJMR0Z6UKmt7aeMJMGpl7+MYulhn8srOrd1on+JnPfguQh15x2uXPx8
hwBQiLCwUajn0Lfh7+g0BeCDGoKMBV7WilVqaAjQlfgDrYnshLIeWU9dc3RV
jJS6LiibJ/3Y5SZwKWLe9rjb2K+WypQ2nt9o/nRbp1fAB6nyCeb1LXRCg09S
LjKPHiN/iXnnDNQENu4C8qdzH3TL+KDVrgqkRO3Ns2Bw8C8ZhLIt1Qqe9vJR
Hqy8adnxSL/+jFLUOz+aFQXTGU7CZAkIuJE59bCvVNWOP/JyJ6jyOFDdDzcB
NzH98Rs17uh9+G1tZAGrDl3Jehh0JPgKHZoOkGiZkNmqwbwnRzjzEHZCO4tj
rJSbnn2m1BLQbRnAi3XnOqKNsMCedUWyHQ3aJbl26ZjmWYn9xd4bVgmDNJZ8
Y41XAbOF41My7eSyGyGVLt1nxhoLSI4AJ+JT2gTDkbwNNoEiNhh5PzGQDlo4
8UJ3/d00pbZCCtdsAdFwLKn160gk0cEd8f9h/cXoSBP5s7niheg5FPUMkcu+
gT1XCAvXluJeSu4kRfytYiSGPW/d1YlRkS/fFtIq2Q12QBo9E1blHvGV80dx
K9Q7g6F1SQFyY0jjEbe2ImPy8PQFHlOh8fDUz15zRD2y8nuShWbFkPVFS4HY
OlLN+T7C6nj1D5w5XMRTtCVJY07abZCb46RdsQ5tOCNhUXz7oO7Qb22J1Dux
gInBWS5hNU7aIzIe9YGs27BcN8KBkw17NoxaEVvXh7SG0zHlVBAtFcaQmioi
qbndKb487v5p6I/aXn6jkC12E+lLG+CY54J96cLUE/dS08E+YEVPiUxUSlAe
P6ZvJz2UCedl7AH3/enTK7CvJgVUl1+RJzdwN9r205z86NBrRZ61AEkYfVWu
nK8nFJwQ5lWVnxTItQvm3Fa8J3WR9Ed6NQ+Q+u0Oeq9mMwo5rldmKepylF42
sD8y3FqKDyAiFw8/OyRIad99PHSfHhgZqhbp8v0hQeaiboKbk7uVqIxQPUkI
64I0GvcIPIb+IvhmV/aWPOcmtnUSwoD59HK7jaxxzIKRuPXr7wkDvHCzBz96
I9CJk2cI+0pMfYL5WNiSoshuiQVIgaduODdnJpR8u0WdeqDolRAD408dwlnG
sNEPmgzLYPIULVcHZ++MwxgkLjYkB+gAUqMNV1Esxm6Ywt58eqiOkg540EHh
SM1rMhcRVj0FhJTZUGuK3EQVJ9mVORSrGfgjqIdNV1pXxaa3ZjTlCkHdWnJg
lBxs49kbYMVBhpii8WhO8ibFkiDAgWEOUX1bCDft+s0qYeo9DVJW0VV9w1OE
ofAiHzL92ddTv3VjJxxng92SM6pSgSDMEPJdxW3Wt53gMROcDnKKELKUBEYf
sKBJo+TZqjm1A5H8dFr0a/r73Z979NBIDvyJHFAaHEZXMljUkgFB2xFe8CHF
EBq2Vrz23OyVkfBorTqzFgxtY4DmKILDkaKVObtpJELPnR1wsGKzJv7QCgmH
L4J5s4R0QLRZrvR4mSIW6N3CCKyj0GNvwPoIABJxpnq3O3J9Kp80z4RlV2KM
ONgw+A9TnsXh3Yo6WnwLhH8psN0i4OHSjOqXaQ6mcF4Z0Hq2bwPrDJjAot5a
IGgcz6BEGcfMHUMaifrhFd1TazaoOzV3w3jmEKIvO7wN263LEtNu4dMTXfZR
YY6bB4P9uQpcm0bEb3xb8cTljteRHQeq+Tmb2fOhJEvDM0GQc2XH+D9wlJta
ZpXmEHo39rgVTICLsNhRU9Sd5R/wTTNyLiLcEYdNDKQBaEa0BDQs5cDqZJGD
soID8m59KSwMGRD1NEqTapoga0phylMeY0aeIceiBiLN3gGMFGlKd3Qam5lb
qkBybNR1L9xOcpc2cGxD/xJMw/TvDIuNxt9VEtcnXsujT0RLELtg9KH6Vl8e
NRuD2HVKuyUHeqJigmTr3J5ibhhSSmbBnU4bslLvVFqL4fUnmPOolv7DoGfy
kYugjSUo506R6j9LL1XJxeig7YJNoiYbMKCyuSBvQsHCjm/oIdqYV7ZBGZbp
AbOd9p0vg0gAJTZqQ4LsyJI6MfLhlh5xRObuZa27biz8dhtcSwO+ngWhp0Uw
k5mXsLtTOQ1ZgyFIdtNn5hMv3fsZMFTWaA2GOs8lQdWkHdSPP7qWUL2JfCYh
bZJmrHlfimbr0GsNnZqIi/nwKQMy8r/mdNRxma9Uw1foKDg3QVCuw1b7nAZg
RJLnObrYomcAjCkEZHV6kDqCPvNQhw2Vq2W46ZeOaIsqawsRszKNVg776hon
U7A53VLjwlGqp8bTTpjOBO9OO/V6McE0prnlEC5sI8aBEa7ZOFDBoLcIPKOa
h927/TP8pyTqvLctvjVvYtk2uDfquyYiNkYwsm8T7wyFl9LJQkut+rDXPV9x
4omirifrqGHHjVg1KAm3PIbs+CdtB7NevYZJPGUxxGgztQ4NUC/K8K+BzQNQ
or01y9fpCTKdms7IDNAdiBjI9+OWtizNssidGw3BpvP6rBWqFTQluTKWlRQ3
LZt2IYc5ssYmDd6UQLjZtm/d6AiQ5SCXR/X1aSTMOZeaC4F3A7klqnzpgopb
h1VTZ0h2HIX8/acgKD8KKSIobcxEmqGjb7avg9qpD9VSi5ZY94XMg2gHDDsA
uocbYIfTdDrnoWCDqysEMcAdT8tLhgkfuAxQAFY5ICS3PEgOEMwVX0j8cfAK
xvnrp6K/XGV5az++CdoRn1/+FQjupMjdIqmSYLkop7qPOkuQFVnyndTTwWou
ilrisaypVjrZza6uHHvFX4SVCfh44TrkgvJ6GmylkwGqhTjJ5p46iFmP+Ujv
pSE/Ryrj5ICU4soR1oVy03/PqNBnLHjWZb6ZcPwj1hmsKG9iucychfLEBmPb
SDScSnTkYI7HQzR501FIg9uE1coZI6ivQ20TsfiV6+eZSop5INFuLW/rGqMN
akjPQ2XU27EI9do8LwQjLNpn8uAX117+Refpv0j8h2gXALpreN8rWYZikc/7
YZaYmjKlGLGGrNOeqg1m3NnXaFkwQ//8Z5PERxXA6Kra4U+OsKh68pF9vJES
aGSodDbBqPXeK71CcjTaT2aOAUMvCgP6KtdK+ztCdj50xzkdqtQ9cZh1qcV2
PFsqPUfG6bJNsEIIQIjNYzErw/nQTCKd0+iGAv8wRytSF4T+kagn50qZy0Fw
go8Ic24fsK9+KRN6dcoK7AagQ55C9DSpuTfDWLu22SSuEQCKmhHqMVTOIUWu
2k6WCGWqnuP4rfzZCOePNg0ECBZrtLBtcbq48CACiP58Gbl/86fJ50NTKIhd
HhG+prUeeDskaew1Yu+dpubxyl4xEVMnpegvXrCP/Wn/5F82CXLtmRw7euSS
IibVa+EF7mnnbtZR4Jd5ZjZRXcdjfyjYIrXzXE2VuVprh/Lxl9ZJe9EIlZSB
ZSRaxVCILYpPEE7EmdoXMNOApWyTZmlAY3pe/KjAzfUYa7llOQhSllnfTRRJ
RLxVziqefMQ+MRknGiLB/xlCE6J+oewWL8p+5JBzdYdSotIqQiWICBiKnu+m
Mzw3ZYEi9ajcic2MN/X8oR0O2LK+/Q3UJRdnb8F6pOoJ6Ep+7kxvHOtOzHUb
3KdvZLmP5hVDXbARL4KPC2PATt/bqIuCM9IQmSyoKVRRhZLluY/EGV7GSzCC
dCr+eJUXwucJVdEin+Mc0P007uY48y269CDSH0qKtnki28PTRagL4AuYjawM
sheW5zC/YFKM1nGR1T9T9Q9Zds8HqYk2ZQSzTEDGlQwERAihuZqDHIiAFa+8
scQdMxvxbdfoEd8SX0ocSNsfBkoisV1rio1Vk+X9jID0ief3CGn2YKUL+F2t
EXxuqSl7NODvEFtJLEmqmU/cEa/JlaZAFehM8v3Ucvor4rc4BCz1CjEvnSF4
gbfkNvf5TYo+8IrEtTGEzU0BbiYf7N/lZMDRG/KN03V5T+rjj3Y1GNvzMfEl
aRbagDr5XkwYZRiX9v6zzk/Ih5J/Sc8tRNqhufnl1HVdZqTL5RLO7aj9YsPx
FPVt2qEKQXA1iidseWUJtyjZbhyWr/MVmOYpjQCE6qEIAFPxYN+vSzMIJE5Y
DfUPTj9Q6BaDiijyI19uw1Uf2SUpptVrhgJXmk3VrNm8cSkjoccyEkYJMaY7
bt1oLTWSrYj3aY4pHQdGuadQgYZr7lZYzEs/CpR3HFbGjldovReWR8t8gVVZ
j1+NV0iGg1OuSeR2zL5GeRRVOW8OrVgb01Pkra+NeV7gThHumZXsuns4y3JR
piP69hrZryMLm+42XpkysVd6jxb0yXRF/Kejb20SilaJcB8XWjAKeb4CNfVx
Pi3WFAU3rYRjaXVtsRWOtcdWiOqwG48D6OKqBVr4veeLvt74lPgwtMq/y0TW
QCmWroNI4jU2EnBi2K3eOB71ONWGFoCGiGrKOuo7F/IS9+RUgIwD7qFGgoIN
0kzFdVIHFMrRpX7APpkNjCKcxc8M7IrdMqVXOWZz2q5AKweB2p0hLZS4KB+p
w+q3K58IYJ+fThpxM8fgs8OWP1yBUrEtmsbqKaNSeddhh9Jgh3Mq66NjQmPD
MbqNcnmnydtxWIW1UaHX7y3Dm0zkBZqREn+R+g3KC1EPt65BLmWPZW2aW0h0
4W1QmB1XKhFm4CT1zZZdSOIW+Mu6RKzcEuiWQnzZ70Zxme8J+ujtqiP6mijv
YBoSBC2rKo/QxshBE2/qtL0YRL72ct7lFJAz9evzssTgQReXREnsEbYCGWA2
FX17D1KBfneKsrp5m1M1XyopuClxEfp+RzTBHp1LNbV+FXKxvJWQXNqFcQUA
YFJnB4lFua9PkHPLhwQJZRMEmo8zvZ3ipl5/8UhiNm3PksPQmwZzSX6SVAFG
gglUDM5GGbA0xwajvjb4pdLLxeCSD111f7r4iEoBXqI6Lf6OzKuTW4bxuZ9n
UKkPSjOelx/2nCUvUOovJdrp3OvPPOCzYOyAZFqOx1YzMUUIul6xdp1gi+cv
P2Z7LviEbdYwIIT8LT8imWifwqKRMnXmrboADdfQgMTMEwxb5/QSsw345uBS
5Di5nwTSc975YakKAi16+3W0+N/X0R7jzJtUX179HwcOi7m4nCWcRCyut1jx
WVZeeW7eXqlKipBAlPLr1Wz++hN72GS+tq4YX8Pfeqq5yq2kmk3n1SM+UH3K
S5Fopjqx1CJ5mQrgBDykMWjJif2vDTdiShEY7c1hteW6m+L94ETMxm+WbEIA
IoNzlfbgnjNNoDF9wjLIVDrG4cxNp8NJAsE7pgUnLR27Xr5itxaTdU66bv1U
FB83zPwetf5mAW6Ljkj/+tgGhJIdJwiFeoETuS2QFKP8FFPD4m8adblqmwp5
6X8u7KzpgvqXw8JbGxTSnX/eXBNaaRz5I0IjkWW+Xwo77FZiB/fdQBkTj0dj
A4pRqiVACoLz+g8LSlbvbnCJMOvW9EQdsx7w4w1/gXoRdGTTudRZ8SXEletW
V/MKCJx6PNHLiux6e9BCVPHGuv5FRL7JnP8nbzNkWo2OXsCenKtWrieyT+PB
K6kT++K1C6EmEm0bbqnFms3uf17n0wOePQez/gYWjAPzUBLpGr1q2ZpIppmn
YroOc4eRHJq8gj9kqZil4oLt3Cp1+t3xopfIcWdsTzkWqyeieyEsH455L9fW
4hmZWtGZveFZwlLKciSMTSHRpAKkgtq9b9fQvOzrv2xHKsqCGVfM2HfPIm18
RU1u53PIOXMbZU5L6QX71GvJ/OViUR+Kyx/FHLhqZjNgqYSOwC5SU5MmADq/
8s3sm7vJQUi7Qj3XGq8r0QuaBFNahTlKhMKXnmj+4CUmREwl8vk9U9sD0keS
FuMn8rr5AdM+DOWzwF+dg85iGFpfeYc9u2vxq5OqmTMD2auYnpA6D/75KxP3
CmHZOuWUp2vkeZDX8RklR1r61Ag+Tsw9EXLHDzKBbHuoicsafXqBzC93X5pb
tpmDPE4XVoIG9q2IT8Q+b8auh512cmgo88aubRe+aMnXoAneEcpam7WP0xRE
cWwcr+GL1xXRTwjE0fpp0oTii4DbWlXe3JCgTg1yu4apzRNKYdOA7ZIca7fH
4V/WFYvi+hxyoimHTORrHexNF2kw1OIl43ABI0e5cRrQ4lTeBv0WKCGXQFlO
hEoy5XxKV2KXoFoWsAC6HKmbsGHZz3nec+qkJmntXhpUYAzAHFAkiTJp8u8f
L8/Ho+XiSVOcC8g1cTjc2QHkVgOgmh/0fBIfZYq7pqtYAUErhkQ4RRmRpv2S
ETahosWXqEt+NIVLfBaeUz/0s7JRJiAnjFn7PbpMnymNocfXiEHjcXt3VNA4
igia1lY/vmIS7eq8DRXyaeTc3CNxkp7AwcznKyWihI+lw1tbApxnMAq8Ws9u
gxvGrjIEimBAKm1UssrOgfm3BgW57DxPomRTqQimQhoIdagNfGab504S3TzV
619JL1D36cMCqE8sKAJ/2ds5MVefrEID/RqJSvPDxnm6QniMNfMgUNuQbGg/
5u7oT3wDt9y+hR+h0DXZxLPuGDTYT9JpUYlbXN2N1SEspoFsL+c8Pc+qWELi
0hrpstZo8E4pW0HvlIJZu17suAGCaBzO1UFWJfOKlMteSeWKHaBOCJ+lmSxS
8n0KXVRwI7IrfOja9O89poibRCDgeRbx9H/ueIIo9IxR4VIBMwTWVjT45pZ/
YWd1u908FSpdOqMN9uidtkxtrbvvhM1acpwXsVIM+8ekdRQWS/pwDX1mrhpe
8h+/GYnwOAdR0q1Y/y5Fl9qA91eVZDqwJc7cqmojEj027GJUh37WGU6nBRGk
Coq317hmr5CEOtuxmh3PEV6Bdy9k/Iju4e0AB7JWvgqds1NzFBY194kCfz8X
LLsQJJlggei2eob4O0nnSJEumX0Ui8jlHBBiQsE1PbN8txmmQB8tkeLsbgXY
sMuZcZXdEgQMT1QC88ejpndtNVRbErmnT8Hi9bqcsafzMwv47ywtBemjNVP4
NaBbaN7j+H0gbl04FP/JuE6CA29bVXvR8EkkgR1bq1TYl+8JSgknH8tNMszT
6wp47sXiCg9R7HkuzDbh9qceUHdWbK4Oqvn/7GimaYpzXbJfl0T36UurvmuT
wuhtjpv/rK/09ZuA3VVP/hIz/ObXECK/M7DYjTs50ASqWG9hNIIwcNokXqK8
/jjpxCZywc3uCyv9nNY3IliwYT/LK3G46UVTEcEO2YTY5lIjrjk5P0wH5Wye
xAfQlHtBRirkenntlu+nPXAp/wZmxvX9AZY2kF/0op7Ya+4weo88QdZqXvy6
X9n/wJXaU64LSfqrCXkwh5T7J1DeK3XzckmOTVyFNnzJdN1ek5v7Kd5+qCoP
26+Gcl8Wdg118Lhna6sRXfoMElDZOzR2r12LwX9boAfxSwGXGQKb6RHC/9lj
0kiwTZzVHtfU0c7oK2Vs6/J6W2YAswYdoa+pcDwBoQ1owcH7FiQA1atZN0Hn
fGqP12GyfSLW2NeOtmB83Fl6cP/3eb0KspPSmGbDdA1nmTjR1Eshnz1gRSYM
S5XCfkrMBFNGNGmFBt6ficSnkHF6pavKfnv1T3yTcDNv/brVuKTFoVE4m6pj
TBV5JYP7uvjcVlRXxEJProQHWLYj47IE/aV7BGPy52R7ogoFAZ3Pdk4USPyS
plVEW2ohf1n164NHDJ124xYue3sIBGbrpCnb0toN91/VEhojOMLEJDHBwRY5
P91AWPTmBC2OgeGb9934CZjpRwSxzN4JAMFj/BDGZwhcCpbwWZkLa6FLNQI3
gkAgPfick8NIRvskMLtTMkpWrYggA8FTeisWMfldA9nkGW0NHP0+uitVCiRB
47326EYUY0yC9h6NusqzlD1NxiA751CPI2O0aFGVV8vBHx0qMI2MB/PcWiQK
JlhafJpA4jwcCUu/hrZ2VOkUYVzqXu/pjTXXGh6pxorhlehD0Q4h2QUEFlcE
ey8xEBG+vuC3u28M3hHHThiEMHYgQnb7nBIC5emaee+K2Xp5BVlCn5vgcnHl
Yxf8XMMmrwSf71m9t50ZC0NmuAAjGl5sUds/L7P8+1RSMmny4BS7LsLHRJ+C
c0CrP/T6/uWgmvjVHEKtiNZZPgQNhiq81GGunOYKJYwAghTjQHIDvQgWRkGJ
RqkSznKNA2ETDMBk52rosHbY6MHbpcgeTeWkYiOMPjkV591tB+780I26JOOd
B7Pzt44aXPZHm0VQ/gpZJ2ak1vp49QhuN/AxHB4RyXYU6h5UdRGDDEdlad7f
ISVXoKnHiirQO0RSz+fW9FrUfnF8y3Br/4vY9UH6CWlCe9+BjKUZQUGw4uh6
MlMvF7wPOjJA0Y5pVFTT9/6sGuKHKUBb5qIXudgpX0wVCjhFRToR7r3h66fN
kYBEsQ2s2h+am+hJ0nA5J82qm0OOKD7tO/koxpXp2pjfTrce5SHb20Og22WH
QqdRM2ZiI3eUwHK1gcs7tGWWSdgHMW/m9xCfXb5WIT4FM+VKTw0EUvlOXCz0
1Haf15IWr6rtenQLkYUvE55DkNY70G0/ioVoHULHfzT9HNKkfqI1V0jbZCVk
6n/+ZHWFNgShWtJjZ3ALQwmOa79zN3w9KWkQBk5oAIFy6sKo68o2nVfG4+PD
fO026EXPDIS1jC8RVTVBXg5BppbXVT9p2N/XoT5vnfDJ4D+6qGK8vm/4ydHB
gXjsn16xLhZM9uPGbsUeeqFN8jnThp71vKL/Id/9aueFLlXmM0UkF0OPeyFS
6DgW4eERc/lZBMkYmcpeYP+6WxtRWUS6KR1W6UMud8a9HRYbrkjxAfT5Pn0n
jmEntxqhDV40tMULjgbGtXFZLzBurdW38tu6YkmqXD/ksTHUFnbV8/UEXsxN
4xI5lGb6yJnLghmi6mW8pjR6G3mkJdWJSX/6Cbu3sPn75rmC6uaS/aPrf8Qp
ff8Px1E3MggZ638udsxYt/+mEC5CBkBc2xeEwx7mgTKX5jLH8asJQvcmKKEz
i8qw89QYwpCN93cVifJZh6yiNxfXn3WpgndPq86BZgOOiHYLk34jxr7591ic
T8tekOCFAOFx5GSWxPEpfKk6rOJJbdacnl9o/iQe5c3dfCSGuHk+4v+OpgtG
2xIIOJhx+AAPGJFl8ghYDLM8HGpW1m1Jt14v9vA+VdUE2I4wfLbrKojHYnff
vEB+sgUNNQ/Mp0OKnmJFsq7OlGcWMv59ZX1BGNO2w77+e08EvjEowmV7DLy/
Ua0ggBJa4i5hP16CRfRNMUF/S9KFv+4drPX/Y+MyLumO+Ccbb8UF3AFLem8R
cv+NKQDqRXzzvMn8XPqQsDexeqj9A8Uu+nP3jyKoExMvygYxBqQ9wmwBVncj
C9OyibWX33zsH/j/eJW4eB5bYFNiQY//VRBNeNFpxUeY/UUcrDysYPVZ33T4
6BAJ4iVFrzGn3XbjCxd0uLoerZREXNyobZLVf0h7F1QQmIsqFeqb9oRBWO+p
Wjfa6epXYNphhzoSJr+k7ZdqLnp+ixxbhS/dqMZFCOacQYO0TrAuCoYj7fZH
8pkceONbT2UqEB4FEAenaGVsJT5bQieSatq1yYuq7ZMcP5zmwRoA5X4sxPfz
ntuxALyBuzhw1YdL+4WQKBDqGeWDF63cVN9kx3bCM4Qbb0YiDYT6pVtE+9OE
SxDsLz7mr4zBiTP8ltXPUg/IQ8wyXS1uWQqVYxrK5fT3V3xiR76/dbunXL3K
4yFErgONDlZWv/cYjo5rX9aEjITCAFvdr//2Ke3fTAoL4IewLt2BSrXDgvrz
Rg5AMb9rwng1nxsXAxw2BAsbVMUMJURniGxogGWcTKdkG/59WK3P8hB/mMX+
BUaWidrpYNlyUAxX4sKtCrLNxuLPj/dfEI0FwjvJDxVn/YhTpl7OGp1Aac9i
RXc9vNgKi9VUdLpTvpMSy+NB4jnBUs/jiHiNhWFIHLWId8EjXh7YlqKl6vWO
IBoZdXK1lfanRpayLXMtjX6wtpcUJ7zfOa/wuAj3E+CQN7qj72nyM48JIOSO
p4rmrysP+rfsOkm3vGFsYEtKqo86JlZkte4kDin3Gj0efycRNBpZqqz7PKqa
ARaKmvRRYr7vL1caj4Up2LNaYLlvdyFD0u5pJ3Kr2i0aYdJ+WmU2vY1Ul9PU
/mZHe6u1+LdGKM+KX9OAgGo+xprO4eq+bAZZYA4HenbXl9UuVeaI9oL35LB1
6sI//pN7HSGFFWxIcZ+zpLmP41XyskUHc8eqHwFNS4g5tANf5nPErYWCvSc4
YLrnoRLnNf2gnf1db1cNbtRb2mRNpF9kZK3l3qbC98c0Gsrj/LrrQY0KKevr
/7RFFTp8fNvLXDeQGXduVIlvscE7GLGVe/i+FdSnokHFAktZybdi2KzIN7AS
KF70m2nWBU6fOv97YxUTcjfzW7DHiochxjQXqvNY9EESytNNgDYvGni5azSD
o5jZjvklUJom1mFXKQUJSWDO5Ui7tq4feIkmBU8ppr0NVFufl93LGyWW1KyM
Q9el+l+OMv2LH74BoJVCgxne+k8Qh5/lE+YBJzSMcVjxxBIZpVgx0gzb7FBB
EVIHc1UN+Jh9wLU8AXgdcSptRvkoBUtwvKCk578P/AljYwVnnu/BBvvnA2DY
5sEBzpeaZxrPwArAiM1SYX7oA1exQJxoAqXPQVWCwIQHXyrfZrLG3xB5JlAA
9lzAK5quyniC3cW3UMJqP0MCPOFQFrbYz57Ch6QG+gOBz/+ovE6Z/wPXU834
DXCPFQyslcVntDcE0wcbYE+wafD3tPVAV1jKoRvpDypQCSGebm5/6XvVKWq6
D3MwIO8xnaONnfTfL5EDFbAYd497oVq8gXLtc8eyJ8BSE8HFJWZRaWs6X1KC
+TMy3FdP6yx+ywETg08KzleDIBcRRc4x5byowh2w3bEmD4AtnT/snc7la8kN
kqhKO8V2q2oi7MrZwkt7fbVO9Z0FUHBAHBnoKGLR/tA2Hte6TSeQAyDxlTBx
rEzEbNLMwyGv3ROrd9eJbfoUvnGumjDQdFR3TbHg5Mzv3VdkQvxtzySftEh6
WRWQx6bSUYUJMRvJruwE1d9UFv3loJZ2f9Q1g7tVmsjeJ2i/V482t/HDGd9b
jtcmkd4JMFcQKYEAwwwBjlylmgefU4TQJZU4c4Usun3MrmRcQrMi/vGa51VJ
Q6+D/XVabVUB6aDx1xgtTqirXnF4cMLscOtgSGqDGgnx9JR+xJZTersjQ/YU
4EzCEX28aiL6LY9qTEw8PIOruJKgSn7R0DkNyQ7Jl4Q0zaiMthoEsxMNC6nV
7OeA/G3Bcdaly5f4r9tBOjQKv/gCTHli73PZemBE+5Ccb1ToI/N6QpJJ9huA
fgq32VMHrmWMZEHlPS7C/NW/l0PO1GlxQn88+NeFSi0Ykk9jcMW3lAHPQ1BL
7yZAdM0BDcQK0kxkVA4/+pbT5uTWQKsUAi9d8Sz2NNl4PvbbCXUAbxLELHGz
8ZxI6wjo9NamvCcbe2B8qps6YZz6XEwUykeofdU+OhZh9O1klPjnOE9rboYc
dn0HkjVuG1Y1rVag+Voz9B3XhmjgswREZVjthre4Q6qNooIjK6kb310xIl3N
ZjtP2noQfnqfmIL1zSsMjQLY9akaxOw+2uAc1MTTzzMiBb4P2AHet44qOfYY
LIUYYWFIsQP6hwKGGCpuoXlqD9k4n4xZFBlUIXomKMp+chki7Ql1PwY8O9NT
jR765CB34nRQvE644SBzBwoPD4D5Q9XAErFVtsK0AEXDbjvkEwCcsUUWFP59
6JSyHBOucjvC0d0QPq34WQlCBjFpD3meGMWQK6aPdNvHVTgHB6K+PFTIjlFA
3YBS1Wcwj1oIaEMc/cznGNJhAeeimQUgSkEUHo4JY+JKdXAA/74hClioyqyX
Lu2g+r+XBUkl0dEOXCzbRHgmDqosyAdMMG33AweQjVK7dVhrGlHJIukCjNpO
8U0YKWXkvwOLZkmpC6RFJdTiUbxl3ZjwHRcncNGrnvK324I87YY0kPW2KDb8
Gez3NxtrP4O5s1qa6nQ0L0gYGgq9+C37OlRfUMQQeATEBCDD8A3+8Zt4+HUt
IVkqyvA91Al+Ka3tGwCm/4m5ukqs5p6B8s+rRc53R2tusMpPHsLeDqTuRDv4
IRO95eyJhXJBwQrYwzCUsC3pJjhG1RQ2qkDEun+p/UrYPZypZ3r45VD9UsFB
7wrKEnp6Tf5Xy2Z/qrDiUNRHQQS7aG+jxCeTcdsElm2StGdY1d0We9WCy612
O3nYTt7YsFmpicIe6Ec16PcvKq9hKAhm6kV7+o2J1plmy/hUKiamX4IOWfQy
k6mnye1ePTZNtinH+RJdCv7UZysU7TNmxcmHwMuB9ppl+5oDHUOt/6NVRv9+
ktCc8cl3xJohu8wOfNmIipH2131fMzvKoo72w6lZ/KtJ/vulsavPcdvAEHLw
Q50Z3Dy+j3vx3U66uGVAefySRyO39CLM3tcaXyeb20bz/7rTHsvIS/IgzIef
5Z9Tb+iVPyy4msXwEE0ENO0gHqSQcdpztdzFVw9392BHyPuEah0pi2SZ4fml
8l2kmhO2zje/QaWg/s5P6pFbBJEoVXMmOPfuYFiKixwRWih0DVqF5khhywtc
xsYQy0ToT31dLq1sR/FJcu5Yd39tionOUOO+Tgus0uzejuTfoV3tJZ0UKQx/
cftlCAtBARNx/+23dfshso/GI+ZywETLsEpwNsInOsik/nErZr3FVj5kXWsK
u3EBRoUuvnkCh2KMPZ/KiOg8fhcGiXw2fCN0xboJcxKYiUGTe0pMv28pGSu3
FRU8G7j9ytwW5hK2UFNGEK7YINbpu64Yp5WL1659f+fxTuA3zz9RwBzf4dGz
va3Sljt31Pq+wBKeGsm8/MKsyYMlwvKN3x8fGKMEVM5QgGWr7dyruiL4Ecji
SIgfc+4Rgwo9mfg8peYKy1+9lA5QkWIqXhgWYiYjIQ/qntz0zIMYStXiVqud
tWF8ixe0gafbEpp5Xf0pO+1x17wtWm4X4B7KeLJQVGzMIHrSN6rkE9gAx04g
9b2L4OwcnA+qi19tyfxI5GzyKDp+oAqg6QsNWbp46HSxwy+zu0dUA+YaaUlS
+Ta0rm341Xqjeb9Ynfkl7EAWHoKKVJvT8mM+gM32egzJmsM17105u3JbvFLl
kqda3Ol95WapBknyN3BhEYDNk6eVZx8XKVzO1oR+p0viHWsTV3iHK1iQAWWl
Pyw0ZQFG4El/FH8W3Il3lXjyQb2kb0zXwyCAza5HqPQnsdVkk0CyUjtT7dAv
fg6qVR7XzaloQDWy5dAceuKB1XAYz+7FdMbkAugoZCNZ2axl/rG8RMLDDWTj
ptQniZ4UKzyaQujVvVVjqv4FojuFCcp+5KAg0uEOzYs1VlUTvsXKU/p+SZEC
Kd7qim/C9wnQ9piLTA8knK4xCO7DMrNtS4g5mzftMzvT61s+gMRz46PBm74G
ANEhe6iSgiiVuBpm/fLfHeBnQMAFpY4lHI5O+G1GmQli1vcEi/ojjDunUfWx
RlRDjp/AvrAKjtw6o2eCS72TIKjGTsxsPUmYPvxr/0G5braATemaowM4eH/S
hZWlYNwDs9e8MibxPiaktlxSRQ7BVm29gcSIIxRQbvGkis9WBj++7WsjvkPV
oGemftBDE/yutGpn6HzdOQFv97uT5594/C3j0AybvBk5lMSp0t0qFtT0DKWu
EOooPyLO4+5ujj3x3uDWtwdnYju7cY5cDSJ9sfsSN4g61vuHcEguTRlYFjeC
4f/eT4KHln54ufodnxJibT91qOJwNorfAzIH2j7vOzMHfA1rjNbVs2K7Ts0z
8YsbUKcN4ksK5nlqKtdhElgCUoKm515s3840dHoo3nFyU8EMeLpmN+0T1tpS
AFJmNVswhNLl2RdYiphFDbVBaTPmPvUane68JH0i61+tOTSjyu/0Fc4iniAw
BvVQNEX5sI76OAJnyeMLPPcnbhY4dt6IgXdTFXJlLunLbZ8AZeLQAkTRpcKt
n73yahWsY6EP41qfqWwJsJyYpjVSChaDa7G+OrRoh2q7cQtxPyfzIjt7X1kr
rGc8XFRKU5EMl7jcIX4U+BN7Rakt20dE/dJB/oy/NWEMqCJVekOgcV4ozq4s
c6oNsBEc6dNHavwM0J76eF5WQINg8I0C0/USgorIOniOs1+6QVPJ5Xd4NCI6
03RmSMLCqvgoC3pJYvoiESITATauT4Odo6+n0VkImj3BcxT5UKwrAk1Elme6
N4LqJ5GQrvwLE/X1kmFq320OdQdqx1M74nC+FgNOOXopnz2dbg5UdhIsgd+A
r66eus7iOG9U1NaMlbioaOHyl9vVu9XWEi3rpkYcpKGXjcVZLEZBr7AOaE9o
rjXWte39r/GJC5UcnOkf9CO/mneAlzCsTSs/ZOlngJvOO3k39rvqJB+Q1mLz
uuHlT0KvWQKwKGuLaAI6Q1cpRwIjyJcVo82HtnNsprr0mV5ujNvkR0QLJW7/
8dIOqQxXx29Psaolvh2tRrT181QrJM6e4CRgOQ/p6ZC6zA4LRlDUEOC3GE6y
4MTmke65LfNoF4rZtytCYCT3QPejdjATCrdlg5DTr0PSXAHZEWraoKAo4gfj
UqhuBh552k0X/HG1W8wDvC9RoiVL+KFDtGkLxR9Mwwz+FSOD4eH6+8h9YQdc
knCKy318V/fYboF5zJbq+D3RJdhuOO660gld9CyH2g0Vxa+GAXQKrG4uoapG
vZmCrfQLvV8HOqjoUfE2ha+WhJ3iPtjQ7xR01YSR5cuE2qQZQ6pwPMWb/npU
0pgfUf5Ln7RBD82cQVcwz9QCLscsoPwyJkkIIlwPqGmzd/LwDY/LNkOz29p2
GE7Fw8b7zGfyZq5Rm0qWGs+1lutgKsRhfhQZAVQ9GQ8J/XBPvC4RBodRrEUU
fNxkTPOqk9xsf9ARNd6tlQIZ39iyQ3FdajEv+Qwwj1bJUawZhjsrqewu/yuR
q6ewznAwc7zEXZTOf3h6fcPAPJ4dtR1nxnuaT+dzs/i4PAYssa5Y3ABjUg5D
hOuTSbzoATFQOIMlO0Lpdy2JQIqKlEn0kT2A6eYfSfaZ2Jt4NNZZkGMGOz+3
/gwWka5Noha5N1bE9iT2gVXmCTiRFjQFKKowldkHGImRJhJgqt6st4pV03Jy
kiUCnMVg/IOSIJzBROsodnvNU+yi9DvlAWRH/A6xV0QOGiMLLEM0HlKr5Nn+
dYhsWSGSAiMpoSKG+9zEEnIdQQTsPnLEHGdgZcP62hrrQz1ozLH+2+akt/3X
eokGHFwRFy3L5led33hNVefAACtfhHMJ1SCwVN+5AspjtCw99ch3yB1io2N4
xCXCWIDGph6xQ1WBNoBEThGD9Cf6ZhuKv0zlcI3wcA9roOJQuUKXfuBKWlJk
B+cnPM2gzwSQNAJ3nnnW9Ns5Tbo1V+N/+NVAz05paHzm66otrfB73+j9fVUe
BRpmyt0Re6Il2VTnGvFhX27cJOiOr8CVdQT7XLTvi86VKQCnpRya0wggtdl2
sO/l9TSIn80wb8iGFKq51mKNKgQtntVIgrinAh7GHU2qgfom7+DawNc+Y0pg
CnsadEMnkvSwzsouhxUf9W9e0xH3/ydajraiS+KRzF7dDg6zP6fXVAbUOP/h
F39d9YMlbSeXJm0UmZvsXkvRe9xW7nW2YGj4jhkGzYWoKHnKbo8hJXqbpgIM
kTtndUs9N1yJmPJtKnZpuj5zNuV4cJwMvxt8cv90uFCS4RWO9Eqmyg5kLT7d
9wKmv+2uqhMwzeO9Qwb4huRzHciza7W4YAL0PX1roRzGLq+74LuTE+uAoyR6
pXJFM5KeKIQwvdudPmF2RHc8jP0ssMiPoLYXYnq5KcnsJsMEtWcD0Hc3R+eM
OcJ8IXuXJSkbkYzoTY9v4ZyeDED0sIfmGFW4Tf5cSv6IkGF20Z4LeGhsqqG9
eOtBuUjq7nQvLV0pOtOvE+YT6Nw55/ndbV4m1XdJ8u3kvJA+mSvcVqHd9dEg
RjVgIC33QSPAaOObhU8GenZ+qCNFvfn7zM8Xm0tKKyAGopQ/5KrGFXpACSb8
mxtairIO/qmJBz4PCUmiD2yc9K+ZUjpF0R/eQYL/mKm8IGvTYQmYeXkxh41x
AMK8hzCJMPYOMACupGk83CSsHpeh40ujahQhKosaWpLKfxxg1K3atDRclxaI
dyjkK8XPP35FCpJTzB61wzd/WeLPsNyRm3XRs2WFxBB/19fLuX6XIC1AduY+
nuby914StyRRtlq9pG3LEw86Y+zlrC2kszwB9DRQgD/TwCBHEzQ6ir2rzgC5
uqg8C27S2YH3M5StJBZ56E/Yk01s19UYjC3J1Ymb5K047LeVgANpAxjxA0Mk
Th/i59Dy7pnqywJ2xSudvDBmWxUnzxW/UlBiTEoA+uluTZMjgUUy3WXiZwh/
+TX1ovrMpnEnuMITntiAucK7JVr1HuDVhDLiZVmsOXlyALriMVezES4Jlh4Y
U/qhGMc7A8A6di63kmJDg76oqbuDVE8cTwxSy62lxWgyOMxzGzqQjwpZkYx/
4pCbz7w95WX5XzwBSVb/EKVf9eD2HldUzDFxZzsHzVBYANNME5DzE5WPQ8SB
1xa83AXyq8yEJTIfpv4u6adGBlrgWbrxYrPUhdPZGuRO3fJBq1uDMC1Y8tya
dON9fWb/8x078Yol0D2Nw0MkJc9ywqG7zO0BVHNYw2B9lvgNIr4R6ReZ/xBw
27yx8RFH+Fpa7j8cUG44JVJsqp9nF9XcDIJDOAy77YGj1ubs76rwGq8u8GlN
67lEcbbpInwUtrTXwJTnPqAJqGjBkPWve4uxC/n69DhQ+wPKnJRS1b2Jrc3j
ZEHjTlohXlIgOR+pZ3o9bKLcMbs3F3OI5YAMstn2JJ2eFQDYDu9/J8f8bNNT
GWpUgNejbZ+Y+1yn4tVqV6Lw6giviA65t32JjfB4XOM3uqYqunl3Eo0og8Gb
l+SlsJaymZpBIJC5XRAKAFteM2XeC+a4SL4VlipOK481qcNwj+XxYsMOTuQw
lI3NfGh/dyYY7PmdRW2FEXcecFgL7B6dv/HJ5Z952SK2uwfKfD5Z+TKB8X8X
DK3Z/LCEBVnlZ/vnBP93MNztJiALqSx2YLpZCP0Wun4XsK5QW+3iMOtoBlpn
LmdWvDOhGxDuVwLqbFjXZuqBxdJkiqP2oOR+MZWM9vLo89rZAmrHQtmIf2d/
hC+SM4c3XSsYpVyQlCm78r9e7fYrVimLLLm8twAo+WqmVEuH598qFQrMx11z
kvP2yKyCopIZdzEJHf439I5MdmxG6Ml52Frsw/nR0GXiSmSbFyvfVlU7ynvg
x7WMPrCWDhQ6c4A/pFpVDDO8FawUOYy6tLF8BdQbVrg2vmEp8hn9QqErMYPK
pmRhaKxRXoL9BdRjOsizdUWTPv4wuKcab7cH+mJDs8EnRBXsei4rwOU394By
BJ1Oo1jMwl3L40a7gMCnzwm58+6mQ555AywIblz+HlzWNmKv4mzKq/q+qp0y
cTtiO7Vq5bgZQdLwTJkours/46N4t9U2lGBH5NU9HFiUuLE5Dh3GPHVAwPgW
imgpq9VsaVfhUYJzYabt/OfEDp+RH/io/6whaSrh8XY9/oXL/1NJmAy4vU4O
rX11z6jQsU+tnFQZIsYu+dYpi7L+DSF7Z7Laf7habpL2OQD1/O/TedA7cYFu
4opP7M0sXk84/hXZ5e+2wOrEl6AQCndhcKoWsdR/iP43N/gB5cXomc+9tDWj
qRioJYZa08rWHK4KNNkjgnyhEnNafyyjYpWzQwqJNcVQyd9mZR9g6XbddFFc
sHP7JAi/WZj6IzCKjh4UqX7zf9PKzzwkKsStpLaKyOtQS0u747LDetGdeksz
uKK0fpghmYMcIPGd+PwNzlJqJx9mPDRQzDmZDdYpQ95YtJLpaSsDGZTXI1px
TVKAPknlThjVmR3yQzOVDJuJAeQkIDe/zWH6cC3zWYgYq90uzsaOpI4evduw
VS7w/XaVbj1uFueZw/WWj2UYQFl30Z5486nWnOE1ytP6XqM0aB7ElLrh4tqq
/JkqiXmGSMfKNPgq90imwvOtmpdGtWkk73243JW3W07/walrnDsiGjK7EX8A
o3JPWYRVf4SQ9ZNchoIBDbdgncowwCnVGCH2miWX97EkMDZFuEyKA7+8EPXw
tav9ewIASxBtGWxBfL9mbml/QivUHeBvV6XfooxbKY77Vi/OXSsKi/lpBPc7
aSO+NLTNlxN3cp4XQ6kh3R8VpDuRpFfUSUBvlzXCb5aNkAnpOYaDGScQuIEH
uJdsEKtcR0lwr1A6uw7I8vSwJlm22vemxl1BW4icMTycQ3O+VUaD5zyREIRN
fCcjxXLTAA3W0c3HxjYE67foJwbZH2FoT4L9oBTyj6i3NpzXkqoTQEiKmpJk
22TsPDCRiHlJMAkLSLBfELGKFwwU0oZmz/zMIspnTi6ROb5Plpxoy/xyu3YI
n8oca/ydxGMshtr9tPtbigJIwm1l/WIePkUIMqb0kxg2q9vOFyjU9k4tL4at
hiWb1/seO6jq5YRZ9oAPqoAb8JKt2ybngnTRml6JtYWfH5cL5bMlQ3l06z1P
10Ce7sUVz7Aw++91JOT24dbUGaN6LZsmlyt6iywctb0s9juiBDkzGKco5gvH
mur30eVov1ojamf7g53+iXNlVNBX45cQKZi5yoDVoR8BtlwcVcGZyxm1kEFh
0QZgjARmObNNb8M+qcO9cq+eUX92FHhYyu8XxTSjm1s1jqigVMuZW4O842Cl
HLUKcQl6QrFPm4bcdLfmkDzkca6dBH+AgeSRRSam8/cs0tBm5IO3HpDOh2mA
gGHAiXtf5VW3/mjVask65BDjPGVslgDV3IV8DSAHWuOSRwUKe+GYzo7bBG1a
IuDJXoyUMXfg6+prQVLxHr3hrRVz1Y1kJx3kq45QvyAX7boMiM5lErt79kyY
SXN6btxpr51oAkYvSIc1Mtn0wbe3HOzS6oDH2tu6QFrXonXKCLTwSiEiaj75
UaCOgyf358C7jftfxOFA0Q4pUwzTSXzeqDmAwMb4mjInWEHjhUyDmy+HBXRu
IPdlOy4fPjY0wq9iHdYxMpuwThC9UgSEbevpP0NPZD9l9bKLYkRNuknz/7Wy
41yZGVana3nyYFM/UfK/pdpwRWF9f/jJ+12xNN8si1qgN94CprQLPwgQvJsj
q4LBSK3csTtbqsa1G+ROUcLpJEZWg9ZmCYaZ16nvyyU4WQDJ3vdsfHWgfXEb
QJJM4Q2TrIluNk+yRySIR3JAFwJHkJxyWeItcymK8jYCVvuqai495+ppciac
rhM21G/jQzzi5RTqP7RmrOrd9MQK5/GRh1YXnCzqdQ+q8WlKmVIuXAIvmpbg
Mlg3eseI8J6y7PpIJiMWPYlAgBsDzFbIblYZknfO8M7CIv3IlpCjxyN1ioNh
daUTlQnFI5coKcFHWq6DtlFXdzg5I7YoRkFucKI4L6mBGCbKJrLJ6DGRFeJl
TOD6NtmlJx7bfWn6gXHf7XnnthjpUJ3pVg3xPqXMAx6SKPUtFm9HnBE8ogSL
QQnpdqUoxNzVH6JTWeCK6zw3WVnTZudJK4IWDEiWYvkNRu0i3PjM0wOTADK+
WgdfGjEd8K5o2jm3EiWYwWu0saJQI+8TooRBElCsyE/wTuOIwuVsxhFdmg+o
ZIfAFLlatQoqLzT6YU7/4MLZ4+4UWQKEQRrp/dGGHPDbcXQysjHZf6vYy0e8
6u1KH2sk9EOs6cKCO/l/zHLp7zg4amdkPInhF81YnzlRx90EGmWnT/VJ+dgW
39ldZlkmECfkieWTaQkVOmjdfkwrrpbClNyiTODL/P7JECDilgfl0oK1D8jW
AjKNsqp5C0uyt8zJju8s50Y9IJjEIBAsKEa9Cnu6XpElxu6ZqU3PxPGX0apO
e8ji5gbInZKFzGEUle9jWcGIXo+v5P2UWthG727Tu90E9i/5UzUySiZe9Prk
Ejc2SgI8ym1WIV317tfPOl0BLQxcu9FGI4RonbwOOFR5elIHTOrffOl7Bce2
y8h9mqSM1SzPgbCfVQvEnRe9i6AOQbFo6+MLQec16YpJWqQ+23IayFS8M869
ZDahLZ9uNqRCYwU1qkBHZzp6asMqX9N3HuH/ojjxzSbHSBQ/D9N86zHJ1aAv
edQqw1WXR+JNc9rJZ/xKH/m4eVxF9D5SF0h++lH8goA1910YSJLF2Q39/lB4
dhK1Z89L8eytC7mATmEuhzOO4hs0DFP2WnBvxVZKiNl8CmV50KL2UT8Gpg2w
/8f96sXbb9LEOiPCO0wvaZRMeAj9aoqs7XIebKFPkTGT1IkoUWL2cn0vXZZU
QRbI/397s5BrCrVX2FjAFmUXefpmw6u98T0cPHZirUqVtGjL+f/vdGY8eyIT
q2ibP+kH9F1FKTdWcnHUeGH6ER4GRJzmiiaJPhViAZzB/fA2rBEWNDtOkHGA
m1/S9aLkEeGuA88wDU1tWmJBmBQrIrBXg3DssmOEUul7/LHNXRJOyPVI15IB
unSU2BACddxv6edx/nquLqxSgcOquavmheSd/rd20IXEIeCQFFSpnc3H9H5o
9w73mV9HiGkDJJXPZnlxk0bmroXSJOu8HAkdybZc9RfmeST05k3nVnsuBEyx
JuTPvTjJEnrdufL7GoAaUxbHLN7YobZoliOJWnDphbXw0oSbPaXIHIKwbss4
qu7RF9duJo0P5g29ajjkKxmoGomA7fFz4NXgJSg2f3nibhu6qkYgTF25veZQ
CMh+yBL38YOTkUAVt6oIDWbKs9hj+JGEhOz9F4d3J5cJaG1wrl92SpchbCqq
Sis3plyL9yb6q8IFVvRywXqwpg3iJCUaHvOBUX4+pT5jUjZSJe7NddmW6YEe
lEbxJktra/k6Oljb6+bh4yDhH8CaoeW01E1H2CYOD9Wnwh7+DcJwsRS2Gf0I
b2jH2iPx0ro2yYjngu/WoXIGSxhzCLj8RlFFevS6ahrZaL7Httrc7iQa1WUp
DaPGllKio7KyqAOLUxEuBGjQmOR99TZntaiKGy++3DF749nyFSZd/eAZXlif
oUaL9pqYrVeBcYkgFBSSzFD8KKw8TuJEdcaA+n/NcCFfzgEHrE0SJRwg99zY
ub/pdnPuGSswmxIQBC1BrlnCG6KHuBu6mV+P/0QbX6Pz2hcxDKImZMzB0WHG
JqViK68ZmugiZ7t5wzNgnwaGLdJDbQ/DfHvtCT/xaCscmG5cdmFID13wVqZw
PHAEFUOGY0MwuEkdoKrpSjX6Rz4J1kn+m2p4l9bz6GuiiW++zr6ZAAKXE/7d
9WtWARI8jjMeAyjw1RLa6GFro0QXr8wKQFbjhF0wB6t+pm9xsDHLl9LxiGxB
qDDCYcDV6M2TOiFJuP5aCXculqvg5tohSvnNPs50bb3NnR5KOJRHtvvqUNI5
pvWVq1sk4ZnvTJYptoreiifoIk4WJVGp+7jm8dUfVOIKMDQ5JQ0bD9oKvIax
YrofOxpOEUtr7y084g8vqizcafYy2k7FO5rkzF4839keuKriM2ZiL4vrihfC
VHXCIGGJwUnG0tFqufB1+EsHeYFzk/o2Xve7kxLF74ILtKSMuzyHBxCIDUs5
OAVjsXLZEYPcuC6D8KSxtpl2SLSk5shoG8r9Mrs04VhGyNe3R32p5SXYpeLk
A5ldJWIkgoYppv3EtSgfv6p+Lys2SmcPlpWRho1qMRvDXg6KcBjey5qaV9Q3
4ooDdah+yI0c9Wk5rWXXJvIpcC4nQZHK06w8EVYty5tTCepxkznZBmbGmKc+
Z6OxemmCM6ILuF0S7l9NcfpmeBs3tR3JsJFiaVzoHTT6iM9tePd9nIoxx001
OtFD0LiB9j5xCBQloRDWwKKqRiPRLvqnNwpZ0okIIuDUAw6zAI7w1HApcEk9
UsRVS9gG8oe7Ogwi6CrOEJcV2AU/pGoFm1FOZKMDXWzdKlpEYGyBLhO6Or8P
4CRsG0QueldcMCEcpvMVVwIKu6MsviSBtRZ4MIYyczM7Xohl57Po5dKnmJBF
1Q7XcH7QLjoK3EOU+pvxaUmeQ6jDyKnFvV+XsMd5j9dfkFx1+NJRcjzqC/9y
1cgGSSPfpj18nbqfCyKpgK0DtJtMXhz9gQ4yCsmTekhiOpNpsiP8qqBFyCmy
/vJG8jRacOHYLWaUKXDs5iCAjbCz6f44pMuuwKRPPKq2se/uhCDymPqWioAr
au22izoRIT4GNf2OwdfMlOz6qt2FQz0GKMFPirXzYW5/2Fv9MLqMhLLEOyCV
AdMucaTy3OW+aR3AB1G1BBzgiX5R15O0U5TpsTMc7tLpOlZ2Vu2A8+fjzSja
oDmQ4FtYBlHmvwzb2eeCNDepblduMllUNL669tXl3+VYHsTlWwR4Y5u0TbyU
UPnEM9nRxCk95eSFTpgdxyfCRTYggjHlC+uSWF1uiNUJPzidd+ds7lbkJhqv
TeC+TAc5G9jmReMmxgaGqC0tqLar1izgA/cYauSeM8nj64E6Qh5cE/QO/pu1
ubCtHDTUOjs8vyGoz9vsVu882UZAaJLRfmWM83vwmtC7W8wwFle1Fhy+oD5/
y7gHO8Sos2gEKpGLHDP4aA2IIGLjRrRMqMVasUr9a5YN7jXONAxtn8EDqvxG
QJIxqogk4bNk5xj8ac+LUFLqRP6ZrOOBKmaCSz8olLBv3gMeuQ/DvwCTAseL
MheM90gyb5X7UIb0pKKs8GJ1KNE8sGyP/nwEpsDgD4CX50RG0Lqy/pGvbGDK
7j+cVy0pvT3So0PaD12Jbo3qB1MLdkVXIirvIMwHA2VM8KpTwZO7anRDrrkj
peJ4JybUD5DxGV9s/RAlMNH3xjHFmvk8R8vKtVR5+N7YOHmDmQAw7s4UIA3w
xgN3txYprk4TaDJ+zt1L1/o5hlnqsBvE0c2izxWAizjjvV6wCw9qDjmWS7Vv
pwUiMFxGUJvdyqWQti6PkwJRoWJqSJfO8QueaEjKY1p+U8cgzEc5+Nfd808n
kl12nCae5bmlfwGlGDDExFvQ7XggPdmgVTu+5BWAEXJJ5NSjBOAdE3qB+x8s
FCSLCdNUpuFXOtOZPfAmv0n5byv4ME7e6jtnNtOazYshTttXpgHdZ3ah/0dh
tHQ93WGAqiBPYnVQj5Z797I0WmHJlAUqENxDHaEO9DmdWhlTCvyIRwoeYlv8
erUC+ESFsDvSeMGs3Z5/pHF3OEh7MMErAgT2T3AT1SJyjUYrWR2IJo6BmZGu
ehmacPgUQbUtCSa+l5CtyDZ9MHbmD0GszNzOj+grUFLMm9Ls/UFH/cZSfehl
5P/1DO3YYMuMBuWlwBYgcFAeJgZMgKfhCy+h4aRQblDIW+viC+L58u0csSfP
N0LHME4Q7PVHu1KJFm0jpNxQayRajbu7u1cnrFtTSC6bX/KUuh/U8KAgq+3z
SN0eu4pnm68klRzKf5HZMkmR6pKfbxgyR1uVvB2VY5tNkeOepCQMl1GJ94Gm
YRa/IPId/dOjWKgBs9VKTfDaTexAQ/y32pdcmMZs4QCicEZsxVfcdSN9CzmU
UxNzk0s53rN4PLTjz55DRkLHkqTinNgfR7EoilQGoQXMPZCeNbqnRk9dmV4K
WC7y0bpLyXHeQONDwUThBBs/WKPlaPMisAUmIjGRiq3LlHdUW0vcpLLDxnTo
FG2vMzixOHB66cXxb3NDaz7LkyVk0prAG5ou26JaczMxfEjIGWpFqrb9G5Vy
i2mu60QK1UKbLuD/LAtYXuHMzXFmqBC+IO0LOWQqQ06xarOH1pguU37ZqzlT
Ns7fMtuFU4Efww2IvrXLTnAom4knqi8iQt8DFbWYjaAVNFRUYVQmqzYxaV/E
dwc3UkwcA7HKLN6qdJYIVSnZCzqmpPParYhp6T+GQGm5G4AIQVvRtaSTHV2W
NJQGLx5S5A3vm6emxE/BwzJ3C0YdrqFiDBNiI75HpeqRrPhxxc3owTAJerwE
MsmVSPygtcwSBT1MY7aCSza2EhmQs8Aw6k9Mwh4fqqmHcKd4SQVqlWIyegbf
MX6GjRR7yBV/vqqSvVy9OmTKGjHlVQcGZuOREv3AZNZfXlGO9q7EqmV0z6JD
wp3JdsVWIsEPHmfwH5EITB4zQZ02aMgDDyIVZUpQRWZrW0cX8PuWG1Rp8vV+
J5oUZY/pUrheENUpyjFPuPFjDeaiOz2hNNlz6ygBsLM6+LE1A2+9PnjJzxap
rGrxnXoLuDLcY5C5eHx5Asoq+uy0Gdni0IkwfFSYFK1ZF1TmT3Yx/uDAs+9+
kXSGZhm1s0gNgO2H6xzIbecuZkeaGTACv0/qqLRgU5ZFkt3zqmqnun55w0I8
IaJ9soRvaIe2jICy7GV8DgVdNge6QCB5m5F78uJ0DWW+NomffquhkWI8IcvT
l0/CAE1uNEK1Es4GwNGCtj0ae5W0QH38Nq9uQu0eQK5Rw30A4egW7QoGJXOy
s9QgIt3xAhIsFWqEX8K0DFyx6R+rzCBoth8QFTsPif3sVQhiGVQSi9LZY8uM
8QoKMVfD8Jg8Gp6F8KpF6LX1IA3vxDS0pyTs31YeJlQMU0h1glzuOv45hrcd
K4c6NJpyJmU7F+OOQw0yriehMX4+snkTTubeLT24IkzHXVdAv284QZ3I+Jpt
4cX96d5/58Rbv1po7ItvnjUeucOYyZRqsxKjkwgyR3+rA232lI4qMeebRiEU
GcTX3V89O1MoplW4PhA+0kg3MlJQ6Y8+7J1THiW05f4Q+65sbIM9cZJBxQNs
NpFsbh1D2cpz8cos+HDi4ukQZXvdEvBzCVRTIhYkpdFHBsLcqS2osiUApWM0
+GHiKdkqsr1OwuiVEX8Wsar/rInAQtVWw0erHv6o3Q92lfHGFxLN6Gpicn9h
02bkeWEswC7bXQLGCSt8Yo0MLUPmgigCB4o9ydq9uCC7xNWq5Fl3vgFiRVvs
rkqsuNC0mAYuKHZhNwRvD0EkHQBd9EW4II+irJGD9lQPQ6+U8VdJib5m+jlC
Murm/B+23un0JtirnVmnz+7GaSSTeM4k8xJ+HUgpoK82ler8vmR2eCxe5AzM
EhQejnDQCVt9ANl4JiV/Jiy0BZhjOs395TzrUMWPzWXKcBCJScvpugV2lNF4
dxPb4WLyKNTNn+g7nCOc/Lib3qebo+Vh4xRP5VH567C6Pa65/wzQFVpZrRhF
DH8o05aE1/bGzggOkDBEC9Ll+3TZIwDD7IZg/jTQRZQtOls78x4OWCoQWjQn
98TVucLk/qrSa3TT/BokFJGtSykXVLWy57zJYqO4uDos/eHG6x1PdpvmUQQJ
wbRFPzI5+WGK5r/e/ww5hA1YAYBFgLj59pzT8q/NfITInlazMh+lslh/fX/H
s4+rkbXDFD7f147Asir/bDl8W96WU1syrpYGlEcV5BZZOys7OHVcnNanHwkL
08TM1yjIsT/olQQnOvusXj4G36W/EG7TGVo/pMQ/mE6BBy3CF7g5vAOme0d1
56ay12YZKhyejZVgdX5A6JS98ReGa2gL2HFXnUAtYxzbkAzSTgOsiSYENKcP
KyLjzdJ1natnPT5VsPfDT7peNWrsLg3wVi5EH3baBMZokvm5nbgYaXWj9cmd
67wztkBCLUsA56DgnXwjhHnrNvMhDZC1phzg+pxEVcm46wdV9iKX/jdkUb0M
SIMvbVRx8abmAPAN0hJ/7hky0+SYj+ea3TDI4ZGrPBYM8ZGBB4gVZWceh2Bg
3PCuorGXamWPf4BormwhbWBOxVX4OlAzssleUZiBmys7DQeqWkyq3wj3l8I6
TAAeeyH7sqUOVI57NUT0XEjPn2vnINY7NMHYZsq9kgZAN8Rq3A3uKArrGlLv
vnWWj01VtBiWUGPGwbd4aX+AmOb0CwestY/J78fiaZPeOK0ntg/3XSCKczhM
ed10BjHrAW6mgI+UyG0T4SHXWITU+9kPL0fAtKUKT2ftEKlwNyERahko7Fs0
LqvsYvxZzT/Ep5/y0Lyg1Fkd2+xpQBjIlACuV7yEeG0hBCHK4y7fcGI37Cec
PL9Uyy2gGcdaRjMxsidSdkp6gdjKfr13w4HfWkt1ibrUu5mhjPkMQXtsmfok
8f22hhYsNHebsOdNbocKzluQftkTBYqgBb587M7lZYHqDAmP74kwvYQtw0Vh
OYsKXU/JtSJcZtVmeHLlvljnfvQddWJyHOG6pKLeUldTGQGy5oIKmZbxS66/
VJxd985KGOYW91E4PbnnhZbGcFM8GD7VteW9uuXCdShDO6diuOn9U427Br0L
bBpI0k2GXyaAIBsvu9EDo0SAf0m1EXleg/qfV+1Xr9lUoCrxCv1IhMZddKU6
WlRKkeLFgcMBYl5xp8NOg553q0y9dpdqAVxn/6Q/as+YC+FTBJHF3AxShYKQ
SzWo+mNSqMfBwLUVaYVxkMbg/YrpsX7M+n/j/7RjBtHFYUgKwHevtZV5P31p
6CBkezaLfinqEMlkyySS3/xjKJqgamTwJp6WylFjRKMZkILXj/MfCSntxO3l
o8zdKnoY8dKua0Kv+Q3mkNhyh5ieOukwqIX/VKVPuK0JtXh80//SINJAVgHn
BzqPqI4o0MSik1baum0kpp87CG3fKaj6E4cOglVsBwbf8UPKAWAh3kKvx+Q7
TBUqQqZf7NDEXn064mCjPl/jLNRSw0RNRXp0VEkpyiDo9lRfMDsmSWDDDI+R
DqQKe4tt/RPIQ7iBfegbgPqZtXKBUDNrLfExX+WohF7X5mw6Qyi7SGj74Niv
+GzdC68DEtK80J/ED15hWk55T4L8hcInUOwdawa9PxLhbgrDyES8Yh18syQt
woXJS6IbcLh71+39QQI2ari8gyzFYzgE84G6XpZaDk5+nWQeh6tV2Kf0ooFq
6VGr8m4y9RNLEaSJn9aEv5+mypM7TNLvXjPSRpchfeU6XJkNZ38wmUFNaUmr
kNlQItWJljAZBvKLHsKpGasBQKlS1qovOkgXT3ocRGnSOPiZHUdrbHzrjzkU
Uz3ZVA/CSyxqVnTPd/B1vvyLYRgZIue4YhgKFoNwzsdYm7Q+L5zbT5BPZBwt
2Cx9jbnTbpMQrV8YDqgMjCojAAnVfp4WA9YciIOjIElZoz4NZM554Ygg3q0u
HwSbCG13XHdHZrzQKXhNNcv0eVVfEaM+dDVqlBVSMSa28Ez4DxvM+PfHT+xB
M0wQbf4Tv+xG0nw6WKtXd9NY6DtvdyUTaGZVCmk0G9wR0fvM65ePBz3kL07p
xuSQZt4yPsjkgrL1J0JGHE9D8ND/Q2hTAIvnD6c6gcrrVIBl+c673XgYTKpt
2W+t6plI/BAQ5QQNiE6ErodkTjSOtUAD9fAbvxniMP+j/Lshcrd/Mrlu3GMg
A5ruD1FaaHBOSCMsgAKOBV5YzOoxxTlGeGh+SPi6w1YAbQF9Vs7smQhKP9rR
S/Ggm/y6LAMwAwUoc8LBc/SdIMCOV+US0oS5f7IcIcEyJAiePaIAqCDopzTn
nq6EIzsv2U5W5sjCz7UIKWwPHe2vfov8OknFmxPNMAZfPxZfkYJ4HrrHV11M
kLD2bwYmEsUcaxVSxR68hwseAYIHW9hfeVAoEXW2TFn7mtjs83shBT3DTxAr
jKnPkuDg7rbmDYMiAM6C9JNoYEkQTJuJl5xlHagrSe0veJVs1KpKR39UH5O/
hQ5lBQyiL1KMA2+SSYuf/xBHwyCwS5uoNhtfvO0DOATbqzX9qj8xp88EhR/9
bv2/3A6XNGBvoM9e+NKB98ejwFuNz7odrjj7JVl0cwZurNmsn7zhzbDh02r3
emeXi9QBKADH9Xr3WhLeJ+vgkDL5xYetYVjfx6zW8ywm0lSRRSH5vw5lmDO+
hJa6hiA6DCWX2bfS3oftxWVCiVfvG1jBEzcYt2x1A9S0GTNLpvLVyuR5fYR9
3sU3dnOsvwxMty8O0M2P9F5CamDO/JxSw9oLp6oVhMKmdO/EM29eanYnuTQn
JueaOGD/kMkffX9ftQWMhb/ZdISyHGrjx+hV/kUph/nVUwxPgp5esNu4MZcJ
HSMgDnIu5+/QS+LC4FD+Z4YRnOlkJVdhlkr3z57yyeu9gQLEKz2SfpKvN+L+
oC6fLtOuIx4XxS4ze4GVPRdbOqwBgFe6qGtBLIhENvOBzP1Jqub9Js6bMcqA
8nFVvHFlTTUfESY9isFmajTcI9/sVtchw+4SI96twhjK3aG5wEf0H6o8QJ2O
Q5UCeA3m8qL0WZPh/1ClBdhLFVtLMaCbJmcTJD3VZIEji9eqQ4w15BbKEw1r
gC3vVOdnuMiN6e8moNlC8lHftxncjEkjgPbNEfHhKeGpgmdryLyJNxuGfzsj
DUTZMLjHWLsd3MZCsI4zlNyDDM5YXyj9Gd3pdqrJQOLRZQtQs82zX/LNooUe
7c9RqWAQr7n+v9E65ycMMA7rna1K2vybxYLsFS1tR8aKv9fgqb0FVAPB4JNo
wYL2/xY+xczykbRe7kwaNWn0rxOW+821VVbRonzTmYSV0xAJcabPPbtuua35
injKLyB7Gf/sUjw71ZmC/mOzejDW9+mKnQpVn2FHuecMGPsKUTs+V52mN+t1
0CqPuh2Lfcxu2YcCFh3cYvy40w1whfv4LvOBEvOTKSlXu7GVJ2ral0zmhomp
nggOFGNsfO/Wt65HTjXC0G7U/xODdhOe7gSjlFzU6ycHVwC5TV3s3V10mScR
pyBvcLICYdfvNXwdP32Ogdo+jbEY2/Yia/Hp2SglZDkzDhciiK6lzHW9qlXo
P3BBmJFdluCyLCG2OxYGH2p/OvN6WEqAYpU3aSVluoqdncXUIjXu3D0dDOPk
KcanCNu730s8aEBmuMAMhGy/LS7xL5gC+3WRB3PBWDA1GSvTRLjqoSKi6Yxs
q2Sek6qDewB0Lj0/b20t/GvLTdTfbVY4Sh/YvGjnZm3T33ezrHv3x8OciQG8
MZWUDAHeOGGYJQhPVWaJMuKouUCp0PsDGIcC7aZkMaeP+/gUr9NiDNDeUUQl
GNhhE4wnOn8A6h9shebWRnZFIvTZlpQ4+z0TmADT7xuoa1K/brZUOc/8ZyGC
xCyd5aHoy9QMFHKW5/04a7As+DTPdEpgJ8omyxk0YRjhetrNzAIBqSteqAdq
m9WMa8NjUA2Ek/6yRcVdYGv5RMIaGCsLxAQn3Ieq8gbo/x+w4d6yjB449mnf
Xh9CJvaeDZ4MyyqXOKCAsu+f5RQj2BuEXqv8HhNTd9dyl2ejy83u9PiVoF9M
F3UJL5iPwidDj/oTZrtfUuZGvTeViRfp+GzvqM5cYERHqJOzRvMMW+x0Cje7
drgNokPyFHHDlXpqOxOzhcsNR0Y1xVIxkiln/xfnuxdqsnbHdGmB/QXTxJXS
XM61ogWlxVhxd9HkiXDTOJ9nWR1Y7DY/Po5Bc+obRSItSfbs0XO4IHlWy8bl
76E8vB2NcC9lmyiHIXeyMQEtMPhpZHarAItFAJCSssM+LJ0DgZiSNfLOdfET
ERNo/WGiyP94S5HyxRprNX6SZANSunYKAMOcEUzYsNKWwe1VO4gpdZJ9+xUl
Yiqdd8jX+Is7l/Lkyq/9pWnPejtsTagZ1ktNWgSKQ+KVO4xgnyXLFoToB821
P8jQuzPaO6wniSaGexFMFt33j4a53utjhWU3b5YUlNZ1a9ijcVRMEoWncMhh
3LjWiSKG+aBJLHxUAD8OcGDFc0U/CLiX4PZxu/FPsvc0FivBWDN2d1GsrpIo
puzgPnkndZMJq90L5HWoUsf/2waw8yap1ROoQDhGaa63UTnSi51+XJYbSBiH
3RrWkJ1hBpIqyBQoMeidSeyIhiPp67UcK4/tN9ziLxaKRB6uQCCC018zn/fG
4eJFOKlz/lRNIRuLZPx4k1/5pOn5xAoEP/VtlF1OrMpI1X4XDsAtE/ONEe5l
2Ei7PTyukkRtpUI2s4+LijUyBhvWO6uSybxBHmbefPz0NWpsHhur7Gyt8vNa
WQC4DLcBxxo4h0QvDQ/7DeFNm9eYgV26HDR/vpOynhUHvzu72zyBNoFoIut3
IsXI+MAuyOVnqGONrke4Y3h8IHw2NX2w51yNjL9gSFSI/6tZ/pLjthQMmOZ+
ZanXluGFm3Mumk0mW2ndbsQPhigeOqdlkq4Mvlbgx+fVSwDBhbKsJbuENrBK
KScNzdBWrzcJlnXT6r91bBEBHwR7Kyez4a5iSwOqMwjaskY93ZXruuxMu9xI
ib8iy9eQLC/rzGYYdUPBBdMWiXw0s/aOluf6RJkWsUz8Bb8xfMLwcRQEY9Fn
a0svOxLXL7AHIf4HWPNHtBBSRcKv/iztDJgrI8S4JmK57yRTw2UgxU+5qAsT
42CQT/p1BLTwwW39YSTw2t2iyrnw51Bjw4OvClTNg/7fY7OQwFUOtXoEqqwh
7M/eiErA8hO0HO4V3e8cqhWe/50BwJmaUA5M/Fa4BLJYdBP8jczIM+hAy9Cz
SRxIpr/2F+QjUcuzrBCX/HMqwKbdXWCelrLJwBlEPSY/25UjBeFoZBv7OBTE
+aNdc1wJc/OFGTigJIziLJGDv9Dq/FMyGwRDAw+8RbphW+LCD4X0SB9UZ/mX
CPXkh7lIo5+KEgLTuDHJs7nK/D3iGqo1lm4tDulDrtSSmWa1SKKmKpi1RzdQ
2v5awWzO7jGafyiSWz41kAxHVRMLJzTeCBktOQKl3s4XWXjLtB+bephd7GYY
24UUKRzFX3i5d4Vc578Ux8bRvhzrbhToi+3UtHNQoNOzICD52PHLIVgEgoKr
GH2S0C9Amxt7rYN8R8Y2uWes0szbgkvKaFAal6IPg+lgOMRuq3eKsLXDVGeS
/ZAuNFwLbbZPqwX0qJ7BTDf7S3uIgPdjnbvPuZCikje+FLcjYMwdZh/YAqE0
U93Fp59+oWQsxd5RX7D4MhKajv14bWO8KUUbl2B/JcJg1xPH7/BA4OnbXHw5
f91EXP4lICtCv4Lf78Irt0DicdPoGzdf7GucZ8WcZGq9c4JFHHSHX2SolkLb
7NEJq90BDbuPxyZiNyvJfboNSSPjkl9W9II9C6DuXXVbkcymsZGSmJP/uM7H
Sw0+3DZHt830ndfNdfkzkEmpBkzjDLi9RvA/nYFRPHSAJ2wkHAdsEA1y1aVP
BoqImITBOZ/wgwde0q+HC0WzVBibFC4T5YP1rCjoXykrFknepWQv8VBm72J8
PsToZAvAIn8IG499xsUKZd7pf/2SmeSC3JAaAunP22FZEXuXDaOL64e1bs1e
Op3P0UI41wQnpoR/2otOUzwn1HRf93pOSET3cA61iOg9UwgFOUlnAC836vae
yKWTDlPbuTwQgg80AzO34I1nxNh7wM0HhnRcGGVe8X4EFC3JEsuw1JBANGc7
1S8vBrLRUWaCVKIDe0KRZhjibbuGhCFKdbtQSd5uTzcsvC8HtZ2UEDPKEosk
noL40jqpBFtA5qYsSfylQrY5DtXWRChqBsZZHIEDf1ynLB1q5yckXfHXQCFG
KFHDMVYw/vZ23myLuAtZryPpYHcn0ucH//a23iY4+2NKo3lAM4wOC+/F8QQJ
0qFm9zUKj4tx1/D6zaJ7lhnPEOhsxvir6DcUSiDAzawfdvvkS/H1Ance+Pju
7l4P54VwN2/Ia3cS0uX2INaidICCWjgBdB+tyFdu2Hl71Zmm8ODWefzgmC4D
ckrTZOc4iJoFD98ze0sgusGZQuOOUdSBvqH+u/m0237T0ElNXKoNEEVPzb/b
cMe6mYV9IAlEyRssisSszcJzoRNOUl5xI9UeAXZtibMpDEpXU2iGdvxJLp9G
adWrReIdb9vJdutw31lEjtvqyR0/0fHNSVrE4+uFb42VHWPiihkUe2netU7U
exjOVHZbg3iYzh3CocrJeU5SoqKPHf+8elGArWRe6Thh5w7irnuxiXTVeFQA
kUb9e4+I7mezDBTq/8hWC6lhFQE+NdBdRn2CHoxngPsnFZZUaqVMLWFkBu0D
VN+FWhtuNuS4WElubRi8PyflyRQ5d2j3r1zoajayjuwdhJE9LL/fzU/rmgBf
ckoZpIgVm1NHcOn6Q0zQXAQRGeb3NumBMEgO24OWN8+ZgEg3AYj460pP8Ir2
VUjwBJxIOi12xANQRf11wb4SMj7NBj2Ok24v4jtUI7260V/NDskKoBAtIuD2
OH4U/BoJXTXh7GhZkgZwKO80gsY70Aut9KjCizqi4hfz93OHdzL8OXwZte5G
HjPSwgK2jLXighGKykBuVgpB8xxMKjaHa1B/12WA1v7QNru9Bi4pErXtcMbv
+NC+TDYvPJsCecj9Kd4BOvsrprERMgDU7yJ+/oEZYbHJvbb6fYbtVqJMGoG9
zM5qeLWICHMfTwFKMo9TkMSlPvEmjXE92rLsUPvyQQDRXt1/4NwdUlmvj9P6
p/w7z4MDEjKyYUxmke4e+wyTdTAbh+q14GkbElhd7kTFsRoY3MVmGkt7UlnQ
TZckP/+JI0IQOBx3R17uDCNDrSiMyHws55WM6LibXFzbPEdWdYLB7tbFhEgr
EAqL3UP98KpWjTv5FXCSnV00oTEZj04qVi/YU0PNmMg7/In1lhu1k//ASIZM
mWcY7qU8sOsD9t3hqCAzVTmEckr2s+KXFSg+c50JWyYQB3UZVgmusLbE18yS
PebW/kBpu5A1iAifV+dyCYJXO+if0JEj+N2hSSJTS1eFqoD4bmTJ1eWxNOjD
ubQmykMXLZ1nJIpQAsSVht4MmOPXg74HwinguAvEQcIGR1/mE7SwXlKDuRn8
OoIv3Z61TXm3RUqC24heJLD6KzgxT3Mcmi4+xVaXv+RfPW/7/45gNfemmvuJ
5bI1fLgxU4UbsgEMipD8NyLdrz7wFGA/P2XKLAfYr3toHW6pndAtPkcS211Y
lIdKFTDjP4x+W8JsVziCx2ASUKY3bKl4Tg07Ge5omEDb0gMh8yYRA2U1SLL1
tG9XSFqD0eVExPD8Vj0R5McdrZNjJMbDWgFt4j4zNnVSuOcarzQGYyYmI9Ou
Kvo37/PDtsRZD4LfmO0XJ8FMeY6Bcxo7SLHv6agNkLo90918EOnMACIOOC0W
FrbGGmNvEcJ9WxFJrqxbEEHeLTbKpyit3/EHe7HJWicnLhcGaIEC0PHtjYWA
n+Knyc5MjYREFHRy0+Z4Zxwqyg2k+0srrgI0DNSZchJkOo1QtPHkAE5h0pa/
2rHbw0z6DbJGLKOfiPjhvdhDd/6xLyws7KE6+qvpzRYD84hyLPik4IDwTcFC
wKxGx9CKCA6zY2BQt4sFy1p4Qj6brCzMWqbQmaZJvJWFocwwzQrlt64DTsI4
kiKQPPEy7MbfAP0bdOKtsseJIjyWDiS3qFa0dESfTn0FkBbY4lzp36BWopeM
5wPWnWJwFGQO4Pu3+4UDX8PaX2WCKXmOaKuB9dwKkerKh2kkTnxSFFl513K3
aseObQ6usAKGsuQc7u0Nssdxw+E7QAQurRZ9CNBe7FUaibukRmjQESRusIBC
GtGySsXwNOA8SJxMdZ9IlyYhS9dkRl4eKqmju0o8NdSkvSbj42Vnljxaw6SS
gpSAPYs1S6MVeB1TDdGLH9lKKSMm0N5yLDu3ZiICu8RTo4As+9zFWFPVYia4
JverVCozFwfOPpAgzwBpt2XSOEouNL2yp3jNWKrRbs5klhCXQgo6wdrrSCZP
xAPPUPMvv1iL0GOpzP/badRxO/ob2aMJVrEGkssMAZPDzTFwOt5ieNftCjAX
m8nmzyDP8gGXi/K+kxNHTto2xIMwe6jK8qVLVixQhOpHeyKovTq9zI6BaItu
A7e6nLaPgOr/4jVOTi+lqkYVwaDNsQQBABqT/cDO1LDwXI51JYKdtKZhzlae
gg3jcW5w8QAZZOpMlM8COnN27IOP0ubdVTLCPyMbF3pm2BHxKsc7LJDOf7aV
qSxedxcYbYOTvGRMhNg1W9Ee/OQhFA+QpWJpT/P2kzpVIPvvf7gQbRbeRYlh
EVt8QXVFyCyv8QYc5WyOOJDg0D3AharscyfZXe03c8urDJQLlTxJycicbRwI
xIDRYXqZupdRe44EsBV47CmDxXYndSdEoFE0MSO093qPI7UOrxTSMfJlC+ve
DAj+g/Ll6d9apmGwcxB4pAyHR6vOADpokuntwCCAPrhw68x7mUExvqwk0fZg
Bw9/NuwznNx11ks/FfosQNz6AYF6y0/W/VqwTL/mnMd5Xj/B9FMoOPw7um1z
o81lMu7OH0/o9Hwj5WhNw6XvtK63LMggw+JovzjSVj84zVC6D0zw1bv9B/jL
XueTerPc1B04xI5pIOxQZzjoOvuAce64jduznjTMuzU8bTS6Koe4ckDxih4k
9UwC9hbU8PoDu0SOuFrz0osTd6mSK+pWZhc2rqxBOdZtxnDv2rVCdWLSoIoY
LZKD9Cy3l0kX9Sqy9STnwiDybWUFbuK4eTG01f3g1o1h+PqzsXJW9rnD0VbD
dAkIZZFg2USQbpHZf+2EUXMiuwOE3R6clloEe2zCrELqGO1Ok6mrr2MPwIq7
AheQBlKC2vo3mcg7P4VpdewOpIV7TTxK3yfKW1W6tSKKsJ6qkxRu91dGUkx9
OORp+p6IgMizCIyI1eZ2qVxxn9ic7LXoY7WdJEjtfEuXFmbbVtS2AMDjRYpt
caOvok1c2cKkNoWrdFoCZJkJCB8A8WVXN3nY4OFY9ZqOYgBeHe+ptREblpMt
f8LZo9zQ1+Xzzf6FxiAb590vWiqpPb553TW/wYq09NQC8OiC7O8M4fUW9i05
mn71eKUkqGTCuhg6xFqnTQbDAIgnH8oAmFenHPWF/h0a126Gx0Cv7IDv28+z
ornHXd3Efcp5hHF9KGcxfTbAXgfM34IoMSOYT3JbGsg/imHmDZSJBghfY+R6
DVQC1CjmAX8SojSDoPDHJDfBYEU01hZ3G2nJ4okAZU+yKUXztAmguZzV223b
Q63ELv9l9GZh+VZYdOazkv3edwBLGv6mRfTda8uKNGC3ViWhW0YCGPo5fm30
NFpQe6/avphUehcKePE0VhmPPA7HeJKuZ9I7Hk7xdxnbCjvVkL4/QHq5lLDX
MD3E0IWRoiOdDHi7aRa4iThk3xNwEy1xGiCsP41gLk2k/ypOmPnkca0KBF0t
3P/fn3J294UQmgWyZdqHqrWJw9p8ORXhE6e50oK4DXWfpAALXdVArCDDanKy
5LkLt8mMHFD02h7oTWcpmbYT5NAALPOHnFokOWuUs8OZWppe7xiZEPnklj5R
pqdEzo+FG1bupJAFEAqhOMlnoSx18+kfddAjgGw73s+q0VfrfiT1tYn8QGPq
qScLAPxteamGwTq8jMc+ivMMOLAP5gPVmEN6oWmDWj/NCMZpd8Itn1YOqIzX
gSNxKyl8raT3gJchuHbLJqjp6Sl6XGVuNf5l1yhHEeYtqMB8l2Okncekp2JH
BgHazYcBRrXtsg7viDzjSmlQIgS95nsyUIF6z261wackdZ/ebYv73YCZTos5
/d5iPvQ8IXUOTwUoz1PEkxEa3NjASKsHAkxxTQ59xoANLulDuLcT7mMYAmHq
RXiV2/m80nSvIiMAzUbGuYw3m1/a/Y4JES8YARZcDXxjpsFCZk8D6Oe+lv8l
IfOon1IoBKOYhy5ZAfAGSyY42kUyBGr9RW6hzh0GhMvScnCsZHJy73VcPReK
jtobJGSM0cRbq57B6cI0nmbrAYzKAbzoUZ1nmdf3iX0z7SiUPrTg9pJzcS0f
ZFRKCHtKJpYOtV4IxbabboydEqMa06bqfsdwqqr7jm0o6jwFhMqsZOy+b1hR
VAicMsdiYjkDouUSw2OituHj5JDVv1O69J6QEsLUna4RiYmX5VGyFNk3IUsd
NjZ0RIIZC97PDwEH//qqk7W7kxYO+nli9dLrKQk9kVuR0s5v6mWPcxJscDfa
6KbSuEauHsotdapXdLsJza044o7hPwiPcXb912DTkMLnL/iEQtXyFoNGqQNU
ag7J6V519rRe44WEJrDU5HDS9MfVeCvwzSHnc/14UkKUioFZSKHSNi4ReQ1x
mVVnIIdFf2IO4wSjZ2HnPT8nlKvywH0vcMP07IHJPEGzviA/eS0HxMUvZxNQ
H6WGG460PiOxboBdXXTWRJUVHsIbQQnZPU3l95s1C6uDl+SvT1njLFg8nH/Y
tmZ8YFO1kSEQo0S8EZ7CYuk8KEkxqmOScl3NAG7HIKPNMf+LEFTeAUubq0T/
OU6CLT3Ag94r3Xv2I02S3hu3gNgaEaaVPvjF+AdvP09VHve7lo4dvVYNHfA8
AcvamNREORm+iF/DbB9/M7Q/Ypcuns5xjdqq4cyw64xxXy8Mble62ospSEcf
9EQayAy6w75r4eP0ShxDvxoHRVioWyHB+6a0c0aD+e6H8HmLaUZWr5h4OY6J
eaWaKk3oXydhy7hgDqdSdbe6kio/h2CgQ9lt9ctYqWGo4tFSICvlvlm0TiOs
3L9govp+RlWVVn2q/5TPz+J61IKpsoLZbn7Zia/t3941TcWHjNhvatHb0tmD
ReHa/tqQoAr2P8FjitrcXqjyqdP+H3fyZOfDIuDQrOHx9Pf8cnxZZqXtRHta
+UlYjG5XZoXx+GHw+Y0h6QPGcq8wg4g+6IKkeAuEqdMrmdMU11tW8U9BXj3V
SFEtsvTSfAEzHz8CCZKRFNQcH0hGc5uNrNLZmpDEBk2Xjs435kFFjrYAvaja
Er9fAIwiEp78nHRB54LHWhNcFfiVU2pUVlkGLKlqHUtqI3ODh7JDr425MJTc
y6odTCoHS040amwQFXnKtj6CDG8k/mTWp0/oBCfkVSF4B7pvP3omTaCWrZhb
gBmtv91j/n/poDmppzEgXDh1gq6FzyogmAcWn2ARlK2TGuYPpfkfucPSyT7j
g6wQn2HHeGRgRVq5/gxHxirS3thCSiF+DjdpvfMAwb7F9AyIwTFcKs71CPU2
Q3kQFITdLwwxOv6KzwOIKvDWud7ha6T7bWrvHkKVSggdt5RXEKbxRCpIwnzQ
rDu/adh3lvwdXRYcfUQQW2alNQb4au9YRQXQddJG2/mW5qTcTG6lGdI8UxKa
3LyagHJjSCkYxCeqwmiqOZ4ta3BNdCd8fZtYKs1l9jBhdO8m267nnKhr4ZHz
zaiWyH5I6kxZs0EtkHchjgrISN9/MMKD6175tsfi7pqhWJBYNpGJAOfEYZ4r
aswii16+F2aj/1wG7eyMVaYAD4XnC3rgoEly5sqkusOKqdFt/ohOxskYn0II
SYQ+4ItfABHvpkPRNBMs06rDQMgwtybymp7Ffp6EcAUpZ7fcpd5kQNE9lxhj
qafeKPBB8PRMTU/Hqv5w7+wx4qnZB19NqqupNwxAareMeigl+qWE5rOcYjd/
8oY1PS+gBA+Sj9y1rVlz0wb7wRsG/Lh4AhPcCZaCdIvBxlzyFtASdxADJipA
rtABRWTKLcUKhifGMp8BHLMgTvU3LtPQ0bVbMRfD1lUC6zuowpYQl2wSw3TJ
HNoca2ngh3mS+ZShyG2SAyfzoN3Q0BpzrQKBvh7v23zCtqj6hUEJGTtieB6j
UVmIyINZ3GE7ffcxX02tHt4NYS6VDjiPUBcKExCt62DCFoiIi6T7cKKzQq63
WG5X2WxB9xrY+BIqRHuRRVARnehu4KDfivAD1LzygPfz+kaJEmBdxm4ivTLn
t/cNPOLQOMar+kOTBChfIpxU8IEJmonrrSA4bbr8rS3NwxoYwPQESL23zDw8
Zmn2gwDl0le9fcQIyiQ2qHXAVtx9OZ8H2M3dgNvuUrpXiwATSHIa4m/mIn6j
StNqah2hYSuAQWbaMKylziEWVn5eqtTONlNFmJhc61VUhfErZqeN+bIg9P9d
ohHaeuB1XfHCms1ROr3kwlIeqBdtkc6ACo4AucIBUq02JGpjxZlAqc3JN94m
2+VGUwT2HI94c8FzHpWY0U7uOJO1cQSLA7e0Czi3c7B9XWbtt1zhGysDNknz
WtI6iu0N+zNlktupRzieIKDldlzCH7e2caueWwAb7GR2z5eng71gbQdD9ign
ENycBH6wKrTlbYhVUiZeiHvm3fr+D0eZbijcOJjSpxN/a+gFdcZJnKfZ0DR1
32nOW0iklKPQJkRUO4/2e6pE12VtSAwr6Zo0GfypKcgmu9huDNWhWF8MU5IK
3OMI0V3OiT6TGxqZ26zZNHdHNxp6fQ69/d8uyxBW/MGGH4DCo6ZRYJMFXuIH
CZnMI8w/kkOcriGtEnO1ismUiZIGI/OoJci29IEhrNyD06/yOU+qe6l/CoJI
yvpF9DDQY/7Pq/R7iryrKfoBw9WqO5V+349IpmO7Y6hag4/WQ3Zs36boMlk4
vpsMdFNlFHzbiai6myqi2VhUOjoSN1i33Jgc4B/zHqupn27PsWqTW+0nRZhu
cXeTcU+9zk2GTVnNbf96xd4wDrHvjYIScrgTzujhFTYTdNSceEHUIyEOXvPB
I1gspJ0JbuM33gfzf74xAdMDzErdUcGaZA9DB9GYLYlv96AEHbXEmQnTG7Sx
iN6da0MxLb5BUEPTyyZZDJspq6CwwC6rdatCCOxLgKIl3O+r1j3eN3wa9/Nw
+mInVEIx8CiwYrPrWwxCY6gtkqZfD+tx62b/csp7vN6BJG6+g0tmHjkxmlxa
EeJj+CvEA/dwWx0wo3PGkx95xRW+t5N86gZBrJcOCyzO9IKh3XaIbHUuuizy
3avXjJhbuHQn12jGIcRZv8sFrU3fxXTitBpbA8+OfMIF+7ER6cAGPHcmKGNi
LSYUhzGSW42d+B+1SgJLAJYGqDTUmmb+0AouSKVR6gYRB0m0aAhkvBcqJYfv
L4oU9B8DxacEkRfoC5NbJJTEFiaeRY2sW6Wjaj5Ng9K+1X8/yMfqn3KtPxKp
kknh0MxzAkM8Iqw7HRrSLkLzigpGBn90nU5wscfKN/j0xsnAR9nZJANjrZow
6CnZLKq7QqzeuSWyjTsjcRCKM2D+98YDiSEGEyfYZLb4ItMyYDuGCjSqvB2k
xZzKW5g3gPh8h2ZjHc/C9Vm9JHfex6a3Kgu+qM4spJ4x44w9Wuc4uPv/UM5c
uA6aopYur/Qs3iwWGBeeSrL+9wZh9nbXLBCGh1Y+oS+V42kFJnEVqb65/rBk
rWLbZNhepcwDmg4YUlKP5uncuAuBxuN35zr8SnDJg+rv/gjmiHsGwLQoTVa4
2pyRNlt968yGTyhTneFwPu/AdsrC+oJ5dKohZn5OuoUh699YczSOGpyErENG
b6rA5gIO/AePpw5bPegIegasV6pYChE03PxmM9tLxlwBE2m5eZwxeAIimS3n
BXMoeNntCjZ0sKX5JN8TZWXUCbptx2U8rFvO9+mc3YTAhUK+yMTv32MUM3by
ANs7RIVP89DkCnXVZjAU2AAPdrfDSfyOE/MBm1jpBuCZBt4udnCycZMMjRn0
sF/+lZntEAfIGJcM7b2zE2Njts6y4BB2d/fv+m7KyKmtFXk7TYwOn7y5qkSu
/mW4piHTUeBByDH90G4B3OHyp6YJsCU7wVkb6gRLv3rF7eB0+PuS44rBzmas
lp80KHNF3TKRZnmigXUYkVj+N7/2SD5OsiobhqnR2E6cEagpUOrjppbTsdeE
xYMhAJZK6OqoKFWJXsLLwXdfYbuL/Z8jWnAFN6/lCllSHs+Bth2TEmj4c9xP
8Vdq83sxmPLTKtuO88Rnh8ebo0TK8+zXC/wE8QybNFR59hxa58gqQzpS4sHh
lks3/rha+SMK6rXin/EWEWeQlezx6SVg4MYEKB6yE5WzNwYoOov1jE4T+vRH
aX2SpD2o3ftEJuJjk/PzzKem1MdxlXolQiJ/3kyspSuGg6CMCFuGZPksfc/1
e9tO7XLN0yBhFS1grcWMy0uimEnAAf4Yc9XZJHoHG+2G1ZV4MLQJtRv0brtt
zIJFmuRsGlQmm4i3uhln/s6VaEdwhUglfxYVJ4BpPIGmpuKfyR/mAuVncMRs
Rcdws+gExEuzYfhJBI/o/s024SK5YiLeTrl5e8FWTRZ12tODhm+xXwpADe/s
cdXkFUIBRrPKvBedAMXOLeo06z6YaAbNjkRP4duocpICPL2qT0myHEdrnwPS
tDoheTWKiPH4A9FwdqWprwAaq2Wvt04ck9hKIarQLFkgJHIhZzAD+bcEz02x
BWcCSbmisjU0dEyA77W8p5+YRxJNMeV+5myrC5dZxrdUnEc/0NDr8tZ8+LJ0
JtOdHsEBCWEPr9LI4jBzomUOapT3cSsprVANxjLz23mMMV8s9FrwFvxphWDy
XTmNC61pQWqjkTenO0SXh8KnUYyMK6Pxpyge87JYvrrrewkMgjb0DbDOoEr+
FuzOHR9wRcBTLEmR2CGMIMcYytTDao5cCaSzzrQ1CQu6QJ0UL5oT+tfG9SMb
Zlu1L13rB6quOwOGBRHswduE5vsSvzsxE1KQZ5NB6Dg4tVahegD2EkLbHWtp
eg/NWRxgHxVeV88cASbgUcQZvcE3gVSPnS0qu6NQkNVoCYR2+SGoravVCSuE
iOVqWu6WAEnU8KyfdyOIlK4KbvvizkewmIeaHDh6QdVPLZ/OKfD0X9D3RucK
MINmjNEmtWjvqOCa3SC2nxoyKiDG95JU9Ea5wy2lvyU5i/FyXAiqOEq1qWJI
Z4jBlRxeISNR0AwGAy3OQYbh8rVJFlvxsepGyZfysqDPAvR34gHTZxonuUFD
AMkApilo0OpBSYuvAywStm0rLqFltY0+eKCTdrxTZaIDuJ2S1PTejKTNaynv
zxcZL5SbpXnzRFVfTmT+8cFrYhOs9OqS0FShVQkZHElaycd2tFeks9LJgoCo
gqxjF2Oy/KUibmbTKP2BNnQ8x3x4iUYQ6FAZT4vKKqkDaG2p9euOouowvz5i
uGSvKF9MLzvpN+ZH11o3YdTVtp2Qb9Ftb67f/upoIGLAUtORJXLxqDzzXgfu
4AWJ8LDnfzwEFzEKd4PrDJw8MhwJSDnOEowo48KGI2GVmTxLNboTUPWNCjLT
5pyZL5W051FZpBwBTHO3SpgMXIADzIj7gjzs/TyTP88rdJ+JgBDdaWW8p7Vs
h/j7dyBO6nv/zDgxQjC0/JrlXZ8aHwElVGzAtDHj5QaEoUe0OS/0TRa+UP1z
4Gq1ZLy231YY/p0ncisK68HVSIyFC8PWe7o/P7tcPiYITvAM1cO/JGHqqrRS
KuSWitVTgBZlGcMH364Psw6U3V+3WtHXGhfGxnKBxOzS64XB8C+tY5TV/uFi
czgI/+SnohyoVC/KY5YO7vQRqGjGCPnpGQgftVAxm1+qr3KJQtMU+xR1mpWL
8jcDkqpA6P0b2OI3sWt3QwLyL6LEL+hoCoF1QUafPnFqlWUru01Zmbd1N1ts
bkplqbx4M/cjaLBpNHaxIgf1Obu6GO1ZItMouheh8fQPkVhJpKfGjjE7JvEF
CV3U8fr0efakHCcnMjB01VUGnaXUvmMESUGU+X4BKfxtezOtPsLtFLY6cQbf
JSKYGgzo0DWJi08rI6KEDEI554qDbg7nOhB2gXYr5EGFRND8dHJfSPtDKYUb
KQYRnoNvSS7WBMO/KdE/Tsm/8zT/ELBdfE7UV/gCcK8u3mxacaTRYzzg2Qg9
dR8FSO601fyin7uXs5zIoXtXdCcSt1p7bW+wS0rnqXdNDnUYRBIZuveuniT2
ScT6Bvtxk+k1zkyFdZ2KHRfw8vFS3gq2iYxFr+tw5k9lkFVuJZKem9LedSbg
wc2lSMMfEkQF6WQNUBU7l32G7oUGLYaE/nTpeM3Rp/J7uV+FBtBnBw5ynWiM
SxVS81yLSQGis2HSXW6RvSYL70E1Iu/q1PfSzt6MzhEtqKwA3M0ETaRryBNh
9mmqnroa1yTDpcJKKqHiCMFRKrOnIh7Vpwudjy7jdnsoVt/4XhYZQw18wwvx
q7GlCpoa+9XpOBkNyiGuJuxyTan5k/Oah5vVXb8vX2GnXy+czLUbLRaiJ4zo
ZXVgE2mOPvdtZpqxsn9CXvoh/XcglPp1D2iw26PW63Bh9k6g+Rk8iE229gPp
2Kzi6a46L1USTdF3hLhslHQY32wrRwg6UtbSz5zFyOOd5c2Z/I7lWIPhQsZZ
5WUcGYkO7Rbae3ctZpEiGXoHmG2WjZXYWCZyECgtf2HRmTrDXjvlMSQ0ZlLX
TMvAXNuCXPt34W7AmJ7QX7wryxZTN7gIGzfqYSCG1czIzKHlqcfyFu4Zj8mx
j7/3Dv2A98HNPZFTBTDoSQY/2LiTZDyFPXiLDbgG7864awrY/2zJyhLVE6PV
/gVTeGMB+dxCGC1iY1CWVZWUWF96Hef4ZTzKUH3RxuFFn92AGYIRs6F6euXy
hr3vg243zNGqR6ZlbBoiiBhU2pZRPU13rdUvMouF+ZE82t/SNX1i3G4kqMtr
EfPbdpx+CPxahQWa9EKjaV5ZGpv7T2M3lCTeNaHy2nm3JL7mm18i6A+RjxCX
4/CWz5paOgTbU1GGhUFaAMFUSjuYdF5Jq1+r371CmvIBAAjdAsPVx9KTkuV5
7KqEUs5xri/5DzLOXgU+XabAwaQXlpIB0j+C9bCCs6AxthYuGzDa/XUNF669
3tgkQz/UjCro+NYifuDLVG8eEjC9NtcD46VkNlSGaV6W6for8MIVgNNx/XJk
WB+Kc5Re4mKYC0Y4DTF7dMgONiqxMaLMp6if4IsYTSgvS0TBuZXSq9GtxBK5
rfHEVIGMdLcdM8bRyQEQmPJGrFGT+qo33rR4PWLJ9q4VxU3Q1qRXiJH6YYS7
9LAP3mUcZuEksQ1+ToEGIPyKgQ6vJEUQNNqZJfShfVyu6zgFbzbNMDynEfYz
kx1dEBoubS02nlWF8ErGd1ASj80gc9Jt6MUkE0/XUfLRvQed71j4VWQOf31J
2YE9wRnD9h+asBEAvH7fenBp7hPNh2LgqTug4c7fyjDTDVW/VTb2JycKM4S+
lOAmcq1yhWz24cSXtWXCPIKEuFpmYMbQ/oLpX6jJ08cpY30VB2Q6/eI9/k+G
fd/6OuNmHLssttY+Mo0pRXqyXGwbPMBWkxMrbabAuVCPkqpTqfVxJF1QxWOY
zNQfixwxAE3nCTKOFWE0M++06ujnrZPMCzBTBWJtedk5uCSpbLdKZ3v48cUt
6hdBftDYH7dB2U51iKVe74m3Vo9esO0JpTxULebP09FSqS5/+JGD9nFk+R+H
JKYlauqqnhgBcelzgKBaWFuKsoLipK4A1xnAEr5w6Qndr1Zat30lKUhaKgzn
Gmpby4T8sCie5IxEGY6FvJPpbxIoOABLGW7jD1eJyA9KwTdMnS4RFkQapcyj
i+OWVxxPkDUwCmqcB5jlm3Yqp6bfJuCsfmvpbrb1Xxj7ZWSV3eLTvczYO/+E
g/YJTRo6TemwmKaWZbWADnnuSTzto1THGnkjwiKY5WdD8MOg7OxZFtZ1WpSG
tVGHpptY7o/BAEBcI6c9GH3VJnzWCvDMfACTq1nBYO5LRLS0FHtyXL4AARao
PZytQW0ruebphbhI/h85WMQjOylhR7+fsbXIkTJUmtqdZIrp5Jonk8bNAaoK
2pKfrXSw9eAgjByJgKgchiNFIJYaBmJIf8kWLQu5v/o65g1fOKK1dyTEUsIh
WTObGOOjANp1EkwQEG81Gtx3nS5v1MH5CrFb1uvBeBOx+jxmrRL3N7L2cYJ+
K1WhbiqUzBBolCWzrr4EqEQlviDlJW5HkUtcIsGQRTPYy5uMLYMe0YYKNatM
+uvs+xOlLdnx0p1wM95lgvKDmvB3kH0GVAbxbTVuTJmBXNsBGpwYm4oNuYQX
ig03Gd7RFRgPu5Rfj8shkMbjCB9tTxllAZp2JD/3732QT28A1kvgPY8c9ng6
gq4n3m6SF9i38asA4LQzJwMAfx86lEwHkE0Yi2gp7A+6oH+NWk7Y8Igcl5Sb
PzMyzK4GyHK4JIwwWTrMQxRmmT5a8LPG2cs2+fYF9n2jypVQvsVMS3nlI2ZD
f5RGEB8atFotZE/r42DzUEyStxHpr0bq8Wd8V4h9FiRydIzlgKOExTPwjHhS
whT9OGWF1Z5Zj0XEAl/BIcOkC+0HN3fLh/AYxNCk/styq3zYHO+Gkdne12Dw
MADTEwfwwCqimqxUln3bPvvFYfK+3CXn1DICbfn2Ej4fpxtViqJB8hc8R3wN
E3HGYNCHuAjkIOikcpTDslkOcFIGhvhnaQc8fFIRHzh8lmRPAonNhJNHzipc
dOlpsqVm05ssCH/lvS71hIrS/jVMG2fOxTHILLJ+0XdtCVeKAYi4gidVbIpz
73nCzVU8tIwto/oKGNyUDF+s8YTW9JePt/RacUkdlxfMUbxKND8wkbkNgsli
QUAvQegQlkoZMepKTp2j3ohQjDb2ZsJ7jBVwT4+XdiMup17tzCw2lO2imW1v
hhxt3Xbn7f3gP1gqBlFIbo6wsCfV1wUiR3YYas9cCL2GPKu10aqCosjAjIzx
smuejjHrPA/ud8hFQA2EGs79eqjA6wMoR5E/NNZNeqQ4gYcPxGt7SJUyjiKK
SpOAuKbgx5k9Qeiuf5RPeMDYnBK9HnmB59mkUf9pCGLNGnS3+SkkBmUqnBJ3
dbxANWnx3KTzJ/HVyHuH4TMMgdqipg3leveDqb+2bz5I3EGq0Ki5NCDBDq0N
QrDJQw1ay96F+m2k3h0YXJ38UYvfaxknSA9DsgQhY/jW1De08kwt2hCjhcND
eSfB3bvPwwfjfGV/e+fCDFjoKangXar9wc1TT56/p2cw/MCmeqVKsSJ/4jTm
RDHHmg1LMt6pAp5fYAZVwEpugudDvLyRXZUG4ewDp9Q4tRWmUuMt2HREuNiJ
8euXxxgQygikx9QnavtdSyfRIVLAZWPCRS7ucG/yVO79hFq4tiIfXZmlRzZy
0rhqioEuHgKNLDw6kHb2/6pbXwwVwGtkPYiHdODG6B9X4Rn9bWBq0kcLP2Tr
Wi1tZlw6S2jcGPh/9KZyBfFCF4J7N5gpp1YgybAF38hzjNx7VuqWr/BfJjm2
EElKGRhjBshGunO3Tb8WFPMZR8yfafHOe0Xcvd8UrTLNAs2kcyl0QU80wo51
o1wosSl90hoxcLkMXt0eK9ZUDdW9tIgNqDXO2tpoWpCQxgbGGUCNrppcsopW
l8vkpnHLcR84HiqrTKmvvBo1f2taq28uBzwX5EAmylDhxzZomqvqYWi1aFwA
IBZvmjnUBx9eRihv6HKJsikuxbxgIoHAqV6Y1m3UZjOcR3454+8D0iHTUowv
BWTzJn6TlqaohCm/a01jSzMS5WkxZX1hVtxKNtAmfhJYIGESNGl61phgiF9m
cOakBNlxpBiIzHKgEYBUw8Wa4Ji7p3moaw22vIdOEGUmbZPkvEagosYHzxR+
Zy8yYkA3QsyHmu0Drz58RTsSwzy2dO1AKYXSa12IM5fIv5XGYmMJjMfXWU62
Lpskg55KsVZ2lXWgTo3zTFHGQTclpCDJSPXKLhbbvpmmeBQXf+M7Y7AvoMyN
RlGDC77H8B+QkIdnOtaWrUmkaUNDbLrNjW1pAptkGpJ/B0YNGU+XxSWSbvst
9t6222JCkn/rau/5bcqRpKJnjVQjgL81mh5VcN88PnK6325O73kQdvThri3c
0oQuyDorY9K4hBNL53WjxCGixDh0p8fNSqDuWaAeU4En2iM+PSKdNy+4Jl9E
lT9JNqXZjtXWwVIUu7xnH+xSQlpcOrpxPq+EkEI7+MOU3Vez1axjA3NDwihP
3P44QWlz1q0eweOMrf+e30ETL/D539FuqQpE1Dc2D9FZUy9zdD7j7PPbp2HW
+gHPg6nHeguYVab3brYpbk0yMwN9Pn9oidMAJvCufdKj55GdUkKWY/zQ67Hl
8UOtCsCKxLox87Gm+HaMjkSui8Agk7eXi08rl8d4BuOUUSIDRC+HjeMtijTq
jzA4dz45UJ8/lTgtaMCb6WRNv4qPV6G32nTFqrR1n4LXsKT9A5J7LA7oz4fG
I/7vQQ07+srJEjZMquJKkEGqiY3nxhARcTH8kzHtITM98JYFHkqm1nrFV0l4
/3m2r7NAPzYUgIjpHkC0kuH9tK6VBDtKezcXUFAoAGOI3rlxFKTZnFiwX4pF
tt0BXWlx3jkqKeyNXQt9cy33d7x9wQFrLKoWiPShx5/A6YL+OLrAthZIIBSu
gwejZVmDwRicwKOyFhgCShSDOpTOLPAA7lgxApBwMW+FJauAw+/lLYuBxoTr
iRQLNZ/6J8cGeSTg1nqndff2nrfjSALGTjb6MQe8vgk9s4cI6GBeVYaH6CQS
Cfgb/pe6fIuAUwnmyAMf2AEZ9buXUVY0lDfLJEfjI8fEiVbNWX7hwx9GamqD
gzXdye+z7IrAaeOAyBr8+tvDPQo9QaQ9uJCLO2V7XJLleSz3SMm5Jha972W6
WP9nOSnDcPQ1NO3heI9a4zRC2uGG5wUVQqaip1ZInpYcjRYbEy7ocaw001K8
+kiIdlCFKz2MGhXmSTeUOglFSSkWNVj93GgkRax5sq6e2F/A4HfItkXj/ZkY
YngYsYypPKvVfvh97AR06lVHoD8RC7pld62FzebrsB8Sa0zsmZraw6/T3esL
pGuT9NisuZ3ysVaUStbCHuB898fI+Z6uSPjU/oIwkn8wHsc88Q23LcCaCRTA
0oQR8P6fJp6IbJlEJyFZLA3zcfLdvkwZ4p2NwNorGCFkQVkdSvqP/btD87sp
WmNQ9r7vkN7hjZJum/HAcg/rYW4Mv80NBYFjp9hEaQ/2zymiU+B+LL/ddSWh
iyXhAr0jFdunMvoe695RtrjA5KzuGD3UBuTNEQHHUAOxvyXjtDwqvU51Gxkp
ER63s8EKC5ztzOMLgM3x0Kkg5r+vrKVUraFe15iOvikTGoUseBXH2nJe0hb0
MJ+fybE5/6j4UZVOuFTnY+774gkU2sUT2AW/RuPQ/Lmwkxo3Dciw/A50EgTK
OzuOQzj7D8u1NyJTuLXWfFNT36zB+JSBmxLW5+BPfVxlkpgXFMN3EUmgFU2e
UG5BcjjalFmqjazDDZ29WrlHAJG6QdKFDY3cODCD1jXZSpjcvX47+iFHKJGq
c9/m/AUAICf96onag+TZVKWjGzdPqWkKAZGHXHufdqBRtQdUsvM3lTgH9oIM
4GOzpEpuxikNawWJsMNnoJ3PuTiqUaojkl8sDk8uAzba9j3MSasnKo/0I6mN
NF3wP3oltGJrd4nibEErLpJ8AJ1ARawCDCyDJLRKkHO4qtp1NADXbJH14mZ1
Ssu9PQNYejOxO4PnZpdM9tMlM+6ODVBdodfstfg/RNrypqwZ61kyvBJroYsV
D+TCS6+V1FE1V0YgMtoakL+BKbxJXv8zbOvdc2megVXG/xCfrBTILDBrj2BS
bm4N8nkGsbidKxJRtQeaRRD3yJmWtVwKinWPeoKrFMnlOa8AxWjgyQQx5z/d
lCq0I0eG0HlrahIsp6Ql769BBzPIf6/5Ek+VHWdp1oyq4Vs+lZuKkwLgjzfO
5w0sYdxdxa6+xhESrCVPdB9+UWtXzCWU4gO2EJlJigAoYb6XzVk7kQ1SBc2p
8a/TgptLEc6fqDCEHM4Pwq8is8VuG/wyjGneBhndDZF2rSwu3f7NJZnq1bvs
+jGPkAW8aX/2B05sxNdVG8jROb/eS00EjZtPgt/WstmsvxkVPaaOLYyM+m2+
sCNcXEhd2Jnwsf9mIXXBqZJ+lQvKxmgtgrcJA3usVBvlONYAT3cNee2Lo3qX
aQ/99sPGSzf425097RQTPTWyB62QU0+zuUuMXlN8vFISJGrni5N4FPsETlvj
kjaN3giZK11gqlz1a3TpE3x1Y+J0nEdmVB77+3/OotXksEY4WbUZ1uA05iXq
epgxAaniDhTqDOzKo9wzXx8JFIWXfPV8WFIRGmB97+EinOiyb2FtirOux6Le
i3wI4M5+3a7YQe0H+kneWDkmLTLvqX6vhfRfSlJiMetk4alw4U7z3P0898nH
I869KJDwIaGWb2O9IJYvn8c/6HL7fWlYhrbKPHraAylPBm5gDJHBRTJ3cL+Q
MJ586alPh9+D4AK3rpnSh9StlmORvz2RlZWJ1bKoYLwvGamRkk+vIX5zielZ
UiaPs6lCcX6WkIIpq1tyPMCvhIwkSkmEBP4Xq8TgPx+hUJbwBZGlSsq8YIdr
AeHoQ+3b7GvlSdrp+nqxGPm+T9i6v96UrzQpXFYPpQpRR8DybElOyxkIcObg
VObYUB+WDGCIbVKGcUb7SsDRwIsxymRhw85AcUq5pIGXSRn5AJScWtW+ZW4x
wGtkr/Cz7E5H0VjzJv61JGBJju8BLdvoUkcv02YrQcNiNX/U1b3jqFlu+vwQ
Mayj15gYg2kK3XQXxUGSxqGKpFuwMlsykwrzKEYHoTSnBgP4j1g/NfoNshat
l03o1soGMLoypBqQQwLH7eHNGEZWhA1QFp14ENsc04fXmPiawJfJt/3sLKFx
bQNnKQnhbB4fQGor8jY11irdeTux1XodLX6y8wuxxNQYKRbN3uhpUOXCveDz
ws/zIV2YyFHVocK+OLp4KubkOoPJHjQT83oHxLoGjVlT89MK5M2RFAddXw4K
omHzMxvQefqTfP8oK84QnncpnYYpaUnNHVL0B6S8ji4yTE1OFPXTbVnJlPhF
t2g1akciP4mBhMwHnHozGcRAKPdeOInYIt9+jJ0Yj7mGN7okZIHO98j3dJK5
of363Pxel1vfk0gZwb0H/Wj0C/xkZ4yryQ7SLfWuD0s7ITc7ese/SnY8W01R
AVoMBzv0zA8WnuZMutXNOZrSV4t4zQF1D0b3tfu+ESPlTt5iiMk/4GXhPiHq
7bTB8Aar9KrtxrM5kL8NYbPaC+9dzHt6RGbf4A+1WXBUCucDvfTOKD4qagZj
Po5pao2JZ5idnNBm2p4aQTmEwK9agmZpLd7UGjAxGQ4Ggl8xU2Gx4zSG8HRp
tr/fzDLB1Qpn1qTpRFf6Z2uC1esmGeHeW9gbA/IcUUvd7NwOtjC5ed9/ePqK
33iYBXSJyAvG48evLXRrsQLVP1scwX3cdHJPDSpZ8Mjake+5pSFYGycTo6Ju
kv9kh4dEm3odXMiq9w6Dl3z5IKfOn53lqFjy+qrdhpJMYnlhHU6Jk5aFa9oP
uUhkVuwfHY0r7PymaYH24khz/xq5PRm/Fn78qNGsylztpOnG1/K9o6v/3mX7
pnATUVMZ4nzedww2wNfVpK3lJQRe1FwgaZhvXLYS8Qn8BKQdQoqX2EDWlDFy
lSIWcNgfzB6dl7V5JO4axnutRAddmMh3FJuNraRHjpxtUdIEji59s5d+uurP
Cf3kZDu4qyqg+zdmP6V3UZIPe8r0zRF0okCTY5EWr6WxZexvsqj1r+E33Ydf
dYBF6BJYvk9+KuyEXaREy/UlPPaFEA6QFY7+Q1g6wlh6c6iIQIt1Cf77jvLI
bSTgFL49+/eLn7rvFp/g5PC3Ci3Wy3oUfdfbTiGsXypK6WGC2cRnE2InJC2H
4b1PI1nI/J9XwwPssijy36a6bq4mTR8qmCxtw1KBNgIXmDtQ/pywrOyqqjUh
nuSDoVbtZWT08BzTxE5r7zTp9VcxLbotFYCJoOgwWNojU31h29PNm1r97G7y
B/rCH8R5k4yzFNFbqeMKAR+urzP+fvpMwmydrrn+4rjA0IqCKkUZFD1vEaMS
bof+xYzvFIuCdyXO+hTICQGFBtlo1gIX56dPHe+U/R0vIcZiY4STpXZYJ0IR
wjRzsx/FDPh5d9MT0NvE4jlDHlggzhsHmZ/0NFNCG6QlOouFK/KJcTwuOExz
UE9nheeKuRnRryUCvbZz1Wq5us/mR3f84aS6+VX2zUCzd3RVd6lnjWziEGJs
xOlUoWN5lA7f8zXpmcNBfGrmTvxeFrrU5gWFAFLRQ4BJ/6qcgCFJs7kWyrC1
eaykYkNqN9sfhJithFSrj4J7cuEVvVDTDhRPB1hjLFKrJtTZ0mXNszxdKAAJ
GoTThpRGQN+b1mpT6feICJeQwJwffv2fIzmZC8lJ2geRjT6fgKtp471QyB/E
6bBVL01w5tF3lVkRvdGJFsd1bizVDKjQwfdNQhIAVQLvRUBxk8WoBuN2FN2Y
1ICerDS+39cBoEPaHe6h4zgvvHqyQvMVXDpuHkaihEtaEMvgxu85dohBYCHB
9WSXGolB1/eJOo8uK7PT+sHYsMGX/w+R2isy3k7tYiW8Ku2Y099r/pCbLrLl
Cds+LIVRV0dpa5QkPw7I98dURVELlde6MhuXuZU4iZ5kyYZpdobiZOvo5408
SayJpwroanvbF3J7XHF3wsOj/E1eS4KU1rJjrqJ4aWAhQyZLabz+WJViaqwg
n9rJoG2vJqJUsiuQBX3+IbkV2/e1nt0k291WcPdXfbBfHO4W3IrdWthLVxv6
c4oei4MZg6vYZT/zJgKzFVdSAJxnSbsnLGACcWI4Rpn1THFAZiPJ1aMpKSOg
86R3xQxmsvW3y+vjCwoiLcnGKWpqUn+PhvHxdzJ3XMfuKzYpRbWGSm/20AFV
+CH60uuDu20B5K9ZCm4NuT6bqHibPwp5QEbTniY4VH2r75PmVeSnY2JLgHpk
Kpn4XwIrwqljcUv0B70PI7BEpUEOM5n8UBCOlHtI6Ehr4UOVQstwU9SK+f1s
NQ3f8QZA4NPNEcYeSq9Xzvo7lmhtInxVwPshs25eK672TW7ZCiFCRkFIn3oA
EnLuoTC1/AjnpC698bvjA3nK39Ix/f28XIAJE9i9hdqgcu6edrjNpYZWycVK
lEBVa7vUJZg80BTc0rtE3kVUTM6D2G1tnFKxKZFqynD6uOlE0F9ZKsHKlgp1
Wo3rOzMuOEXWvabM1tciCj8cPKT0WJW+xovnFF6unE6DrxaDvs7sWAFEIKGE
9a6QFlx5J+wkEUJfCX6SKJ8mtSna4u0wAKHEFizuir7+ZO93czvX2k7SQdSz
903JTV6K6rdvDc9ydK2D7f5R5EAtz5ZTajdGDkhxvhdiPAL0QL8CTg5W2/qG
8GQUzqxI6ja30tNXn+96/tj4WwgCYr6btuXQpP1vjcdSl1VqEOyPY5b2wt+q
s2CaAgy8sqLIlWTHUoyGnrG9bkoox7fiDVtmiMyIJoz8B18p/HDmLe/Dk6G/
eWqVAK0hf1xdLtY9532lxtMNgUjGHaY8Q8YgGp2sd7vKtG32A6Wt2/iHJpLT
eTmAq9RjGL3Roi5XLYnqsbCTpz9JlXkR9kaom2fk2Wb5euagDV/PXLrRZfXb
wh0exnnDgspnmK/OYv5CAfrzkLG5Glj0Tdnf9VApURHTG8vxLwhETj+8/J+I
fj2+i2inBOQNrIFLx7i+wTqQTFspucO36oJ8WLiO1odUlq+f9W82PG+LVmgs
LLz5iWOWau1WR4K9MV71thotgttm1D1SuNormNMCqnvfZ74YpoOEaibmn08s
NJz2IzQ4T+/WGAV35w2tTwDUWlDJS9Daw2SshOW0zETruGcSHvmlqLlRFE+z
zQknSQkdk9vcxGkUJogZAQTvXOvNFXwRQDKlPPzGSCuUrnokne9dGG25IZhl
FJ0BDGQbPY+fcXvsY6PKfYxEbVvMMYyhOGaXjRJvBD08rDlTSh5uZMKSdhvn
JNohgPxFCJv9JiV6Ia9Acs72HNsRNzpqjC1ZaCosKxXHh21Ap4e0oX7IyOGt
k607l1XiXgqe4DOJp4VcgHDkF0qbaYaBLb+fzt1eZpfYb9M0wVljOFnVXedt
Xus94TuMPhv9U5BNQE+DZgyedhO9Fgbc6ubPf45/SEzJx+LJebeKOHB/fZMr
t0q1jL5kaRCxMol4ynRfS8I9ReCv1OtYJb/41ZdEKTRrbMqsyBJLevrbsIXV
4Lqn6pygf1ozUeFgbaE0f0HmvW8LCt5G7TPb6Dnmi1GtNeKbvRxzSvSXGVSO
Kagc0IrMmvRDTw5TBIr0o9W9RDJwFJrSlGzRlRDZjXjdMyi8HYYGGFvqxZLE
my7qKKRXB6MYoTtT7NWDMV4AffQZunmxkWYx78Pq55masVe+WdprUpWHJYJt
u7CObWhgoad+ABx3h2AzOdg5uJCiLN3ovW7J7vzJquoj/NQvM2bS/xrtU8kV
cTbl9AKujHXGtZysTv3c48L23G/hW+NY//Hexvyf1tmDZoCpKGI1zNwTflRD
yxniczcMkmTmiFw8D8BsxLS8JeVtDuHRzIEVX+LuVhoAZbc9asp4HP46s0lK
OQW8zlDxEJ2vPTcB/KrnL+Y9u3OYpjgp+/YevDCZKLk2KITmebh+S2xp6sKw
y1IzDsPHDZZ2e40gV0ezgGkW8+212+iZtmhycF959rUf3SGnfAB1cf+DDOey
TMGbNxn2nGTjbxvHq5/F3OR4uVeS/ATRLl454dwTV4lRSSUBoNnDNom0pNb6
bB10F/v8aT//NXbBJESn+Zg5d4fPrqCkokOtETSzI+QcS+Am42HjlqeEDbvE
5hxt02EPduOGENmFfrFMstpgdRMPfuPX8OcBIdHUOQtQRENJr8KT6NIGt6LR
X7GG1fVF9x1OSM8zaCU7WnZ8+TZ4tx2/OPuRHw6NhL7UZsqC5dOcRDpOykAc
ZMCjA5VPyvlmzZz7cHYayV90P8QXaOVYsZTcNo3F94/vbl35R0eEjItGJSC0
jimdTbfk6q8sRFnW9ezjnlkKQYkPpWe/To2hVQH38thEzNIzQ5NidyPmZ/gv
yqldp4nivAHWP2+6kRqRVe5qeBDW8SbrR7PQ38d3KDVsmA0gp2dwFiEuOg8G
644NqV6BdIzYa5m863ixhSflFwHy9yLfy5SG1EyxTC774P7qmWqFfbcNArOB
wEBktNTT1shV6ZZHrpgZEphqMdcoxEIaPbKYg1Rd7sJh1uQLBlP2Mc/2ChlG
x/35k70x68z27kOh5WQfLNfLI7059ACi9Tedj7521JWtOjdvPfr/lGuu4B/0
glwf74ly5cH9KyMavTeKBVjfci7uOOw8wRCdtE5cI9LHJbiEoCNouJVXHSmj
IWwgw9kJKENW7DeZGUyyQOvPYRLfZVFcSVF2Bm4Z4lUAhu802UIDcS7VVu4O
eunejmqHonVC3dZyzNfGgPfDGhrlnX2bnA9wcPOyuXtgkjpnaUTpv7UVyGhC
YlCCEEp+2X/1yJX9OM/Or7L7+Zztullov4Qg6RyyO6ivkcjC2jzUJ6Pr5OxQ
Oq1ws4/LkS3eSTs0dMCmwhU2/HRSdWmudA4g3yxuZ8iSeAIvjUSSi5HmFzl3
SDF2rzC8a1+AqE8wnTX401RCVjzMmhQ48MCDiNypabh0tpnp4h6l1EKAb7Is
UPWgMC/e0GQtibMMlGyEvXSo+yj4p60m9MKG2Jezf42J1s1RnjA7XPR3Wy7o
TlVW5jaE8wdh2mzQfREaV0LlID/7Rioups8n4ZptEH2AMo07gqdasWIpLXq4
aXAoFAMrYeLEG8zsKmWxU2RJWnfgAgVa6hZw2L1+K9CqzYKBn8U7PDn4mZFP
kTgw56rHgFYWkyzx6c72iWr9S9s0dfdrqVXhdaQt2Xrdy/FgM3v19saEktYV
C5eQ5l0BV2hzJMzw7XqlHoa/t9D97DeA0J/6oX2vHoThlOZ8zuWGfYnoGT4M
mroUDtfVbDMnpBuoY2CaDFAMBDVqJnSsB7MQBiC8nblGJsC9F8kn9dIEzOQL
LjhhLiRQGjhQ5PnGcERKBBYHGZP23N1Qx1tK/e3Tmc1ykqw/Fh4C3dnbn+bH
IeD/Fso36tDK+utp1Y7+XSyV7NEP4j/fFB/U/u64xA+RfX8f6TPpbSDHgybE
7hOiF3ghPF6jOU64koCPI/nSLC7tx+urJRsNAcix+8yDWhuYIcTOhxWFqQn3
hh4AwHLXSR2sygZjoI9Hip12Rt2+JEAw+xWB6ZFHYiS9P6ASodMwGdVKvtup
idxg3Fxj0R2VpqwWncFIgbmVlN6frg/tIatr87ML+7CSBLtmlS7+qiJJNY48
SpVplajrHIVZvOxl6xviZkKdoQJHUFEasdDt5PHxHP7cAcKwKn2R/VVW8dGB
cvO8zWUK//dlhA7BGl4w3gGggug+kaJo8jjS7sKLVlfVWZ13GUp9Yomo8uvT
IGOPM5KBye2KV57c34bp+s/3JmIdSyr/3osDdYf7g5mWr5gGlxNxKFX6kSMO
lIg2pM5kMyHvymbkgoU4v7va3OLhALn6sbe0UdyW9YLh1rQ6A48zeeDIIM4D
yqApsnve/0p/wBBCsjUYzCGeXXLndU/LZDH9x/SFPIpbQxkitUGdWkH8ySgB
eGTHE9o/YK4QaSIjmnPP3zvJJvat9ABdKGxyMq15al2czpPjBo/4Mq9UXLJS
Sl97hXHJomRVVjbT8eXowQFmfMk77HJW3KLPM1R4moEcFy9XLkRPKV+U+Aks
k9dRdeVYb/87iHRFHnyjkwWOwzsvLuTDI3nfTdAtgN9wi7pPIZOqrDquKliJ
CAQ+pMCIuSALV9DZPrRcakkkBZoygojDe6uS6cqDQvf9Zlup1RrCHLo9mx2t
Y7/RFxp1Delsz3VuqP+dKZmTx9DROeczayVzia/etnBz6A+k7exx2s/xDTaq
49p4K0t/5U42xXmtWIiQswplClNM0msgnzhsSSVcr2YiPadhb+ZnsjSrWZHL
kxrQi7WJUOAk8mpJtxxfXRGqGGrZz7U2fTUxTsNGz+opEdPzCVfkGbSq0T2F
Mup3ML4ibfCZr4MUCzHKMamDtDFpPB5J8IC1FBZZ18Lz0zcpFi3i5j81SooH
+L6Y7GSnWOutCkGUQhs0LPOpspoI4zZ2JoMQJ+w957ntHykBrnShB7aUtTI9
yE88d/hulfejVYjR6PGY66moQ1dcTSnJPHZBclIrbmmyrkvVCzklKsZNhcfa
vW8A4ZHlH+pCqcchUuOkmwj30eBBg81T8trX6bIdRF9wCyKovNFyRZ45RV+Z
NTm1cp/oTtP6qPDbYX3vI5wVVAFX8zM38dznhJ/jhlhYiswaI9pI7Ij5N9OU
iaiqBFd6OzbzNr94Rmv64p1xHm9kdN0wfISwl9+yXMUyptGEyUwrEVECXaN5
+9a96eOpHjc1hAT5h0mDZIHOdXpoDuFNfSoxpW7HyxCIaaKUmWivfGQ+wOrp
3iNyw+2PqBAV8q0UvHiuV/kcuKVH6UODhQuYwKc+vDjsg3X3096G7yP80+aJ
PS4RlbHOQHtXWqphHVJzhHsBqInxYlgy2X2oEa5k1ZVpkA0QwEqcWy4kG5NE
CZ4Ta2RguS40NPC+ySySkRuwcsUN77NPmP/781o9OQ/yIWogwsEbS43+ZPXu
37GyV6Fh7LM8drV6XmkBaC+YrdisbtmA1QYGWqMl9UFjAmb069a3ph5CYPz+
iYDjytb0kOgZUKUhDDETYYturkY8fDDUGVq7XjwxoIwk/uLvZcyUOJGxbApM
25bYvqRm9zf07iguSPKpWbVajJV2U27Kt33CE90r2FrbcHQbG7bfi7ZFGMQL
+ffKNJY6crFaivVbhcrrMldIB79qalTyFbQ37D8I1Fqr7toFJcee3rU/rqx5
rPPtU90wEOdkCZtRKbAIRmLvWotkQkwTu3oO5hT2AA/8HxUWJQt3ItOf64SC
7HzM7yB6ecEmmN9KTo1tEcCDeXWw3rbwecJsJjbVQr96+B0laCEAMlbkEYEg
rpdigsDLNnYZaDMWqjSpb2iikRhRZ9Nytgv8gyyruNW4/0JQsu7siqI+zVDZ
MlickkDBZxv/Y9b73WsnNF0qW+rOBBEZMKqp/WNNudbz87gq7EAWkOMYb6IT
dseyvinBafjkJ9a/j84fIhQGGd2eOU9OLJS2DDP3DCGSwCzB3W1LZFonOsQj
P+e1KcT8FqwGt2yXKfn0AYwNkdt4nRB5UYZY2YMu9yIuepKTvPpccAX5eQ5/
f74uP409fOFXOoFrlR5hF5J76gUo/uwB4bd+au/wJXupVOtZhhZlaDo6Qfwt
MaZGruof7N0K7JQIYGdh4NK+D1PZMnEgX7GEPZ0vRE5g5nfSO521oCCPMsn5
Vrk6H3CeZRNYdimQIeNdWlaSYbRwk0v0ztgt74mU5Yxs3nR7cQQs/4W1qZOu
bbYHcyVgqSorHPvnkgEjhOv3lGUcxX+obKspNkJG//BvDiJsCIiNUfNXohNh
yJ0BJFIrfRX4hvqW5aV2lu2czO1u8RlMANtNyn5uvJG4VMekHFfK3dYtfmKP
o91WiQXc6uNf9sc/jbPKqSqHrYbQ5ptIjrAWcZmBvMqeRvFuwFLAhh34Z5ww
zw5KJCjP9ZHUNy8p3tneBRn8UaGgyPyg74ePZkW7bujnMn8MsvgQc6/XRnp2
vTrZDSX3LtCAseYaLKKlxFcNOcPoTIM7Az6B2t2e9A1LAxoQrU2YajUNq2Qv
iV0nVdtV4mvCDIDQBll+hrQcrsVjKzJUxxq1UGtBNap74tP0w23jBZAD8VMk
UypJZyBFIZhWAqmeCuACvzkgwwVG/8GxzI8+RgzDiHNNdYX7x0S7iYeQPbs7
l6THYc8X1YqqMaREiBv/F4ZGX3YErvjjnYa9B399eeLTMmP20R7I3YTXF9T6
glxXY8aw7xFbrWp7daDg62VhZDl0JpbaOwJ3R45CUpThDVMoAdyxJut+4Er5
yAVz1+tgnjthYNuSSdjeTGumswz5M5VFRm/Z7NONN2jUbsl/2jUB8zozzQdn
7HFKAzKDWafQG+/Rjb5GHPumk6ZNqXTPQl/Aa035Ocy4OWxDLYWelzo6d9Ys
zPAZkxl0igIp8Ygw9rdGe/NBmOEhuwz/sKjvBgtZA4SJRe9LYZ/EUnE+DuUK
fspAAwlrqiZ1AVJ9CNdbaQsnaP74SaCN7poxUPung6GwE29/Y48JJqgmoi5p
B9OK1gP6rd5ZUF2LsLWG6DnB09VIKF/XYoiJ0LNfHx1A8H+MFNj7WvceJVVt
Ooku9CpE05b6+YElznAxe9y8dbbWsN0mODPexc/nlwXddcqSJCPsUwWpQad6
kZQf7DBKL8/w3cXq1MDX0BC0e540MjRXYkSqMIhY3GA4a2nMCruzcKOod6jb
e8L+OiDiuD5t5i8AbTkCisnJe/LrKJ37mbWtdvJy3dT6dWg5I50fkcf13lX4
2B2BVNQu4SNV0LMyTNF/9QNfYCYwnlJTgB5tfYUmAUT4TW/P1SqMtDQjhxE+
XKjhNvDzqEOKmlSr2VKM0pwsp9GB0yvQlRO9/HZbVFhZbuAL0zTXBIXR/cTk
D5MAKOuoJZ9uAbDfI7M3DZWqQ+l7br9TJU3MPAGPB5Lcd6Va42jGdCIA3ifa
PvtwIfA1Ct6i4TmN/ybO3FTjbTgQCJjFMewLJpDfl+lcNK01LmcPbA4/wWCp
tgf0dsoSC84r4bzwgVoHIjr6b14Rw2/rdxJNNIOCnOFe3Y1glKnv0t9+wuMH
t35W4IIawCa6XC6mi+WXztGjZFpS2CHC4TmYBWhnc9Vc0uAizyOa8z56+2qT
xWom0JalwzwNdyTyP+jA4GseCEOqgAucL1v2QfCIfnPZ+grs2lzsDXDj67Cm
Vmcef3s8Y1G6JdDJ2foSkLJVQkAhIWvVQMrAbDLIPM7GTIzkiSST0pcR7/oF
tdkXlSOE88+w+4imMJ/rqLZs2H4I7sxEKYM3MmCyPL90+a5FHiOzrf9MRAYY
1br09ez7Hj50SY6JjDxOPfoiJZqnqdmEne5un9bTAH8Z0W53ROuMrbl2lVkN
Kxfg/4EDygsPUaxruSo0/YfHDCQIKfJNbpEHWggE2HhUvYzEHk6U4dJuayEJ
U3lo3OtRgBpLN3pji1DGVV23afMnLFsvU82n7R7FSvt+BgUGOd2+Qg27Ux0m
f0+jcT9VIhAmxP83M/dMNRZFeuoTFkTnqj4K1Pc09fVTdnJFWJnsuGpoWOAe
cW9TcxvOIQF8j+Xgt8U5b6meUgSVfTE1o9L1N9tco/3rp1P2VRXi/aGVwsjx
eizUSyJSVYstOuFAE4aUq1F0uHBlW06z8bsxTHn469iDCOLKaOqiJrP88WyB
r9IuGlCfK9pKYzd806n6coHIOjKjV/NTzA+Gfk33wv4KpGcJyMU7ANUUNMGf
3iEH+vMFb74XAg9TA4/FXUA1A9P+dJQWJnyXzzyVVyruf6yUAhjEYsT9l5W2
HCq6cV5GAl7x1JW9qpuEIwnKd++RZWpNXgXlmjFzWw+flnyqQiG6EZQEl4RI
tUIgaq+NE+Fehi/PA10XVjzNnplBGzrqLdsoeDZUFRyh8vUGByx44Y6KMM+T
E8qg6bF+BP/+MtC22AVXuFu4lLR+P6Zo2G6hrCnYDmrOc9vK3TL8qUYkkFD5
7x05g6FL9lxDrK5SKg6WQIVLZ4swjO3XZW2CHHkLjAXw3aPMzNm8IGnQ3Sm3
PhGy8fFm6wlqsCc21ewvObH7rpVA6NVk32oXTcq61NF+Ktmz5/wsC5aDgTJ0
tZZZ08WW0Ld7b1zB0SbX00GFoDpMB+DmSB//VI5yaN04G9C4hc/mnVZkGB6d
a2P32NC6VFgGagauwMuYmUKfVCzRKZHzEh+n6zxzj3tsp6koF8SeSz9DvREz
/Tc0CuQ2cLsPAYTF+1IFi2oXPc7efAdbXybn6OSGfMotblbjkNNJ/1OAl6Om
RGt6QfEQhhrTgOy/2448XgIXwNSVl1dKP/CXSWBcEWTLfv2Cl11cqTwuYc8k
XGf8UYSPaXe/oUP0t6BhNDOb6FtXsM9j8BJmj7ZqB/TUZWmU1V32+tbW6C46
QdAfDqEm4GodmtkEhQ8tToizKw5EoSfx6ejUO4xONrhW32f26KKKbguowTMp
5iRetXtdzN+phuwJ0i/qpGv+ZR/PfGIXgS3AWjIp12zTyzAUdrbQOocz4K8U
hQSzUAVfVCS0A2ck3+Bz3Z//euWC6Lg0mWSqNRViG1EZjVVVZTbYwU2QujNm
36+lJaMoufyJNQogwueocXdsrX4GOUGE2f8cRYma2CGMzrPLxhTnpdsHGoEA
IN1b+c/+cRmqez0nOeKjyp8IAKeDjwiMRS5YaQBdVUtM2yhTQM9m1Gfrby9q
QyGgVC3XcVjUpxKaO6NXIv5knMdeYaD3LGA9GirR3/mTWzXFZvc5XwZZMKTt
NeRN7GKyP6cOEob/jaT0Ev241xSsB+H4b3s1dTE3IoXyStugSKAXiRMQQZHP
mq7+tuQXe0jfefhDqTBGGjo7bVan8OTNOa/ffSmmddIdJ1ev+Uo8uW6KPIn3
HmM/eIZFwzlylCK9BdTQkIoPWmln2Kx2BV+CV1oEIWvlvL9SI2PjuH1sI1jg
nnbl9eRMVbslFUqXE3iigbtB9rPPjNRgxbams9hxidLdXittazeaSAQ5aZGg
zkd3qht8MfSBQiHNUdFHmcCH23wx3M8dTjVhsfQIhMEUfKYsIK/jBuS5GLlN
o1GUEzQu0z/3l+kem/OjqS5HRzIKXkGH+nBvseAfE3vfZpu0SoGzNy4avDfI
U39Syj9r9/PV5bK0E7p35cEGaqKHDUuDBjfJtJ/Sx2R3h/kXn9IaSxPxCZ/1
3lfsrDtuC1NUgH0+j2SzG1A61TB/yAPMZWx+I5YysgOvgqnznZ8C5GAMx+az
XGYv28j3gQ9pEk5MJqUV9TzOfXMn+VoK5yUs+WXCm4R118bC4rOfsc5V4sgU
8ua7zC8KwxqyZnJQL5XufWZFvEgScku4Xp3Sh69bfbmUg0WUILWLffGUaSUj
r8mtXD1DMPwOzLEM2kDBD7ArOQ146Ga/0P0SNe1sB/rFWO8hOJuLIxVNc4mc
LcpuJozg2NNYWNMeLMdK3yIkbA4AKaPaia+RoA2DsLrYOHPOdmIm+DBqduw/
tFpBQUtMyUCbx1Dn/pbl3i6aALsTYbXDyDviUgEAQPAugtcIxkcblMu4DRzN
Bg4TuE3Mg880Bm6oBFpkL4Gtd6dnw9AnPVKJJ8npmTZQQWrAobtd1MbNbVPV
9UCHqmj6kh5xNOZF7wn5qjr1pluBmPYXSUa9BDiGu2czYapaTyN/ANIP+97a
02/8gPZjG0T0aJvA7m/Dfez/J00Oi9nj9jkmq+k7K8QKbn4XnG+oQMMRfzrF
5iwUF3E4zeYq1dGIq3hCR2FEMShSbbj5wyl56tc6St8+u7bp3ulTf9EzGJGR
YZuUeHNhPEFAabavReQS1K5J/h4jTVmLClSzbyBDGtBo3w3D2UwC4a6Dhi/7
DX3pIlNl8DrAWHGHNrsJAeGJjixfBLErP1QLO1rLwUPP9Fy0oA+OEyKZowjn
FI/oZSZuwjoAX6juV/hyCEACvyl41ileAwGuUniVfuP99f7HIxWQk4dAUuwD
x01r+/GBSuves7/K6Z5+KAz9go2bearpj4y4R8ZddGTkbORvLqaceDK8/IIR
JVVQOjPfPRnzft7IgJf8MtHchal5SOYGqT3GDter59UyWrD4nFlFN8zIZygB
vdbcgD+k2S4AMba3CZX5HGNAC+3tu5XheNG3qA2j+UQ1zQ1Vc2yHdSl5K2bR
vQ0MGoVf+nX96Gwfvg6OYg2YLoJ3rUfyL/h78dmVvNBB5EsZjAbF/S0fAS/J
mqUIgHhu2LZcBR1l3ySKHgyz54DE2/kPFTEUQkZxivlnJ1SSmyAd/ey3l5jM
LguGDJGhFqxflGoiMVy4yjmxVg4WAD6+e4cKmBSJf9BSp4ZML4v3uaLM0vsr
jDlfHVv/olI2MgZsle20JKhQOvAbNp0LpcqvJTjScXYeDlBvYYjNnFoC0iCL
vrezvA5YHzlg6RxKBXHj2/ixIPDN+6bOCl+QObtD8nNZPoat5XTSKonszpGM
S6XSxiAsZspeqqF46yqPziLK5g7tBGNlCz32i/VnSVDRHefbjXgxz5F0kfld
INrFK0IL8kEdClvpsouBvd0KRr5lJORVfzoWWpn+ZZiRhuyZptrk1MHNSLFm
v+3XpuisoH7evHJzBQmZMUwqVniSNKudzlI6jaCDRYT7m2M0N4etO+0iVMbL
IkwNAbZXN8Np7JSEv0Ie8mUzBLmb5vnPGjd+Uk6ADLScivv4txi8pQFRyuEM
r4Pof6NaZgGDTRDsBIb4Qqr3USahJZerPtNIwWP7cdx0QmOWkhrBe6oNujXU
Sz2Jbj93n7pRJ7QOgNfJXJrRxMhk78nzaGV0wrss/6M2vwGuePUIpLjdS9ar
N5oxCE5x6SzoDgeFubYPq0l5tND1TIUCiAp6gfXEZJUb5CnPrOWDX7uWnSha
XP9LCNTW7cxXMRkNdpU+wq8nVg+Z3pRfE8YtN5aG4q7B7R8uplC8VOZSBWKc
g/AyIpTF9dFGQ2TCy1wTQV8YK7IyWJzC5Vj6dc52TNQ4d53R+7xAOWR2Vi0I
GU1qj5Ph28nsz478rm/vyJwozWuL2XbTeRn9FBgtZwfExmZ6T5XtNTOtLXMP
I8/7S16XFF0Lo94h/T3TPy/sLPpDIR1LKYVmZh/FQ4QGRFb7VSFtRYXLYCVW
GhQuAwoerLAvptYEDIucRhZ+t+BlecoJu7S+/0380rpL54a++MU6uiiLzQaF
x5mr6bUXH85KQmmwOEm/oPB63QYicDJJ6A57V0jkwcwEFAGcnArTIOApjMZ7
01ZT+KUfGnRrcSN2CPvHV/ATZ32njkin9YQ6/Ja2X80mjzc82oaP7oJn+OLX
x22xiAsKMd/OkO9Kfpj2Zke4znOFq7/r4HW+akUp3dakOB/sQW+UkLSBGyJB
pJIGQ94il85/eIfdHQ0Sst3D93vSLRVLeUldaA3YMHTozl9Gp32hhXZ1zM3O
6F33adGb/5WIOTM0bMtoDuNXgmmmvBGQPh+v93uRoA4k/h9m+g7emYj/yLPg
fMWOqazSkv8eMRc7lXw/7cYOXJQjZ0dMg1If963/6+eF5EVhcjPxDjiQqE7n
RCfYeb0vpW7eoiQgP+LzIKXZrRSt/FKdNozZkwyIpvCL/RpZY7wwYHKLVzoA
DhfrWwBBvwplYiUIrIUjxwDlPJhCFpkYPN0rvafCLfWrZ0S7ld28FHuexcoL
3NaR529iVfrkrNdrSvXCEFDOixGRtG6UdyRsZUnYVbttlY8FU3PszFnB4oBp
1hoAkQ+ZOMW5i9+/1gzlIebp+ab04zxxkdDwflT8n3ggUoTDLOu5PRQhX30O
2gExsAKkNmOz8k2neRA2yUVNJvyvu85X+nvsdzOR02jCKQpZDCcW72B4Xg+1
Z5IT4WvyxexACatE8JbRkhzGvsv+M9sKqZpUPxpNyE0/EmMKtuwCcy6SoC/s
YMQx/AkwlYTjtJYhrDu9uQ0ErDCl1hPX2/gqn2M50NcV3LXr27/xG1m+SL9V
AKwT3ElS24lk6YswT88qX3jLHvZ6VpWzniEYzjlKaCPFafrQYu1aqybYhM3k
O7+0Kf5ZfsJSHFXV6MUea7kS4GVg5SGDTj3YP2tWF+cVibvMdQI3d4+gsDTF
u4oJDW6lL5V84cSGZVrYcgbpq2umVwDFGfEK4pXOWdkMzjbg1xTTIql1V5FP
J9ecRLJat8v6hjLyCHI5mCc4d5zBNjNI/yVkYX0Zg8y+5n8/BXAE7ilrjTdV
CHPxNed8FA5SgkZnf/JJ8kc9OdscV8GMqo4Tx48icuSvpwNnhDUFWyL1xUfY
7XN2cxA/ouXX4johN78T+Y2xnJiCyt2sSdIOOPd4YnJ9CT3mtbvwj/wG+00f
g7ga+zgBiw4qHew5m3t5kmD7Fmz6Kex9B/OjvKvmMlB6ym9fwVSlY5HZgT0b
GRPVw5zWwcs+jYuJSDcoBwn7EMi4jLB7ztTX8fy6SPTKH1g49XU2SkZmak6x
ZBMutPv4ppcNrlpAc19HU/cFw11oh/kd6hsMRPLruQN4219ogWiM8m32Bad/
NR4+F6s3GmRh0r5esTE3oS1kv35mUco4c/fFtpEU2w8lJr2rFOX/5Pi1Xjxn
pR7dtFulJeKxrDQlRMyBTEk9DoJqcp2YRHJgcyhrbZjSxYwEVij1Q83IKjvx
O641VDbMvcdBqzZZgYIR/VUL9p+pE6RS3epj7/qV5a814Os/k7/ouChxGvUk
1R/Wh8gNta5NsIl871Et2JKBP/8QPnOs3nmsP5nZoTJbtkvMeFDyaqzCKuOM
Zxb62q5V11Ra5FeoFRxFKknocF2euM1z51oMbMTz5KwuZYahtYsU9PPM8r1L
PrjwoFleoUALFxIOgiXVjMPaChHz6hN16yAKub02X64fG5y6xh5JDQSUPGfj
trrFJKmVVHOk0EcA+mswyhBbqdUexTm0XxGb9H+6jAAOBJwCppqq+Y8pvEys
oOla8jeKVFtrbakiTm3X5tQKzngxhCZfSn/orjAW4AnmiWxESkef5GPDHLaa
5ppzNGTSXN9HeNOJhaI0/CLLpJkvFTbU8sUrVW7ZgIWed6pbsz7pfkjx/Yrq
ba3RAQU/Or+fPq9crrrdoCF3bt382IHxgkoNXC6a3RRhMILmuh+bzL3C/1OU
65LFyhCDLU4m1KhQpA3To8K7Bt9iToNdkjWcIyVKlFWpLKn+nvLscqNQQX7e
aVMrTspKomBOVlWiv886x2Wh8JrlqieVF6Ekfz6E6VK9o2Oq0RaWhQfTtgSB
YyV0VIxDSCpWfgHhBLHlHhG3PskTely9ffoQD2nriVR2M2Pxrw27qkjYbL6K
7nGd9950tSR6ymFfWDaUc6mPYD7JyOLTgYxJ5ZGNIRXHrUZMMwklfZ7LVOmR
Ob5swst51+gko2ZAaDcIw+4Tbqh0+jOFjy37S1rFMCOaw7a3n17oDAn1mQ1L
QNWmTFslQhLtxs3Q5o88ihijFLGZMfL6+vR2IrZIsH5kLi/bhy1nlpNUE/3K
rm8Mz4oN+mU/QA72h70lUKtaCb2F/HV7c15A6uLIo4/VJn684Z4Dt48juoBM
MDTfxqKp6fETjqi//FOc65OOrSKd5JIkIsFRCZwBaZB6yXFxTsEV0BhWkvhN
zhqUYIuNbeyo/Qkk7AQ0P2RKOY4aHcO7dsrET7a7V4rbIhNoSEJ1hPh9iSuf
+7Xj836CRaay9O9hi/RXeXiE9dcXsDUOUFxs/Lo099F+x3aLTCsYGfrrMOwX
imm46UR97VufKIHZIp8C1XN5S9Q44GuN9NXgCFPZR+VVK4+lE2jypy9ldura
JEaFuof4uv0yc6EEoGe++OG2lfywFgMfKklpJhhqsqmnXMsQC5ZXCFGJAvX/
uDha9dvw+oSFZcn1USmBR4A93PR0OWTBveJhmnMEWwltYC2hP9Qs2VMJDTEl
8I3et81kNCoHpsoIUHAjSFRV8SPbp4ft5rXTrjlqoibuP97kkKod3s5PI3JS
2c38qJmOfgg9ZVKheV4NBAPMda1BmZUkvveHlnFUlDmsRoALEAe+fvFwr19O
Nmv/kdDaBh6lvhA9HbdNtas91dLkajyHiRvHFwdiaqUzrTi1GEie8NYTw2gL
sWUugMbVnRqRtvGljrj0I+CkLl9RCKEOfXo+of3ONcrXCZsxo/lfs5gw75+j
UoiQOoKd/wqnyq7ahloVd3cySOP6rUF1Et9yevxbNhBYy6UiEBgWhhCx+s8P
zj958888tVs5ew3MDFMBMXUhV184CwgyJI8cskKfBpZeGTbKqQ59wbMFw7u+
gRycOEqxBxyU2kQXAKEVb/aN8ZGPctYbJSFuBQCZ21R39mfBd5F0WQiU52Rk
SgkgOuQssDysY4kN/+fjuJ6yjeW480yZGsedjIT2ugsYFyk6/czGYoeF0Bc/
Io+KeKfILzG+29M0qqqua0XXyP9TPdYFQ5kmyYC+iub8VabySj6DlayoUvXT
BDKxhtHtCm4vDfLafnhdykrPSMG04pvosAmY/YId/k9HA7qDeDckQKPG1cjN
ds5qzthlX48fHemhL9jMud8ioc0LojJbLKhtxbJ03GDyKguKVLIZm91XetaU
FfaNw6musG0Frml/ep1l8DbijgIiqeNpEEmcvv8J4tHGzbQejOjICMCpP4M4
au2tiBt+WeVyKyZ4Thv9/DKVz2O6tQKcEolum11Hd5ivkZMz2oeNvkSNeyPz
7omAyTJuxrQCE/n1wfeuiimMGY1U8gNoehhtT0qIUhku69WZlJcVHjop76xj
T/Gs2JTk7t4SdJ5TbzyYjjlC35VplxT3hVOxY52Kd5q1PpswsCiMNA+fjc77
wzY427B2mRVTbUKQvnZmMYgZBunIvbjNRfORfpjby+TPdmUgoreAc/r99J2F
wWLsueszXfthg3cumLCbXUncMhpMOmNW7DmOmGQIVu0Zzuci5YF06VpJ43rn
WtjAag+KCNtG4DrMno3gYZ7AzkJ+HMlzNoGD/O17V0MML5+zYzhiUKdUkOg+
43o8RxgQPph31Wky6y3PIrDfmB//FlWuyMSTSaqxmhebP6rt4OffCMhwCyFU
L3GBw2Xv+8ISNP1dw4F9Hc/nkC8qApYk6nTlxBqaazo8NobUsXtdz0ABprm2
y8ioOzZMpVPmaagH1q14sGFUFibCsubym+kxle6krLPLl8oWHRAB6HPFNnAn
6DBwkV+GwNub7uG0Yd7yO5T7umjV7r8/8O2F3CcnRgYhLRYuK96ibRdbyqLY
y35JZfGgzi593KC3SG1H4FC7ANsusfNoIpfI+aFtqai8vU20JFroTN0CYFny
pstf4JRaer5AHGpnZM8mzaY/Wm86bJq2TH/OwYkMdlveDGobETKq7os9NUlj
ehEzkru4uBPvV/TkWKYjb/5pHvn65E51rTaRRlqGG0IzvzqibtTRPlMj0F/L
damirZFoqD2WehfnFDkfdaEkjBc5IBO3SriXPlYxFC+DA8PnsETI63809rEf
Y3nTQpMmh3pRo1xRDWMuVKPaCFEjltoaNxr/VLCcu4LIiFriBnkzXjDZ1Ok6
BJ3tGmDDUmo8QMkXw5/+S9NQbvLWGlXZgShgFYjC/wBKvXhvOnzox0TDt0IQ
l4V2ZhP0kTkITDu0bn22UqGuUnLIkHuouxiWSGfdWKdcJioRg5JThkEVbZPp
9RW1Od3N780LfqRXCk20Qu/m4IbF4JHGvIFdjxkng7KeJN0NdeLnuYhtdi2A
Q6l6NAPd/2xbkpGGVbnsdERz4wcY/PhPxtO8dnfnmzM2Q3qFkf9qQKAt/ksM
nSq1l2CLbS5+ps0fSsQACJQDSDmtwkNxwX0lAY/joroxq2hcIIRfNtlK6ljB
69LuqMJokVhOA59EeRDuKYH9dKeo/3Uj8fRpjFiYZCLCrpQc4DF8rprkQ9dK
jq56XMNh6jlDygGWERohUiL5/FcXUYlsB11ZNenFhWIbpTEVE8TpKNq+f1Ti
diEB8CILNHl6qSEB+Q+BEP79WqJWJCUmeUGo/ts+j8bhrqJn8/isNNua6VBI
x2xhKS4xie7V0hn5WACPDg1ccSPgOKWIyhtB6ioatufiU5XRhCih7euWgz+u
yG6Wc9kWsH7je7knvaE9R2ccjkOfn7Cel3j1VDPaEraBYtzXWuinO8Dyt1OX
IMjzxtctq2O56f4OBKWyykxs7m9KhmUnn3605M+1BPKuL///OV48kcy/FlZx
kRWz4RzbNj4gUDEeE9ZJ3H5iR8vlCDnn/N4/ltzFokLmB7Rf3Yxaypm9fZvT
yQpxRZjcg/DlNRXQ5EGQNzIwh2G6DWsWkjpRvmTH7GhOxjhhkVkMPHPDMNch
HbBRvUBODJxSATI65tuJSdY5sZHF/firADQ3sZJKJ+jsUOl0dOhUeeZctJYS
2bLedyUX2Tg1ysQMO4Ofl7gVWY5yge0GlfzLDmUXPHoVrzxOMef1G+mpGcyZ
/CfWomQCHk/uW6FlARk5N7A6908dxUuguLfT2UYjeVdxeIWnp32qwcnwYQAn
EUC5O9x84kk5dYBJ9k2gwg5Q1ooiB3vN9cs/XSTdpft4c9Qhjey122pWNVUy
XuDWVVglRAkRePr6iODleKlL4FwUFHnylJtkwubw/G5L0oqMcMJ21duhp52l
QtKNWMldPOtbulYPi3obTSip4TqpmZ0IJIUTrMBDFSetx/d3IuwF1duF5Dcw
QgNQ76wRqWcJ37RDjL6b189CzC1z97FScm+MK2imF9R2cgTGXvPcI3y33YIV
UPQwjXZx0pzgTFM5FpVcanLLvfqlHMWEJHVxn9E53+7mPpe/khewjTb2oV9q
l2eQl2Ip4sePtxrJUAR5KUPH5Tt35Qyhj/YThybLwAL8V8oY3uhasCyZjTKL
OBV9wXdjzvMN4YYOTUEIJdk08JmdO5yYG5Dwbrl7OEgneXVP/49N/TvbMw0x
tCYXX++cmMGbLo3/qd13/e/6B/TUs/xIAgDk2Y+LdPmIiiA81vzAZdwmR0u1
ktuFvJ8Ig9DCIiCTZHFxuOwdvRAXtW7FCP52Mtd0moabc/rCarGHoPJiL3lG
hRcyLhI7OitQGrVHJT7hX0Hopwe4x0JvJy6ysApgiSmN2IyjtdC1pQJtb+hc
2WxG51tlQ6BvHwu7J+dgY/jAd79sH9fPMriYEDr6ogqwVZaQHLEbdNw94U51
nugHpYfG/6uBrUYIbal6H1201cyi+QPcn21inzVUgjP7AMFMsxEcZBpOlVFx
J+H+kF/zS1KVmn6WirjO0z2vUWY8CYwTH+XU3LMRq7WfxJ3sRC7mOSf8F6i5
YQ/MIXipUHg+AQUrg3QW9PJ5McRn8KnecQZTfIhVj0kkhaS8+GLzbHSvFKjS
aMiOXNSlvZikP91TDDvTIruJiDxd44HxQaGCs+k1dV1oBs2T+fL9RNKwv9vu
0k+VkTDG6lJEL17VO/VGKjRM4N+E45o/34Uxf/V8VXOkOUJ3vKrZErUffjVM
UfhJc20w2UR5ZPxUGIjXbABP+WnSbF41jnI2LTs7lazsARolq2wsJHZQKpCm
h4fmgrtUgRx03Fn+1XqQQAJSs7UjaQ6a6FxtGcZb/dMCFaIJmPBvS5fgWyiN
Ey/tr08N0X5VozWTblrgPg0aXTgShYfI65Lw+8M50TDGUDan4qoItp7nvyah
skzXjOGijW+WK9gIRqxK5iA+T2IOXW6g5APFKaJiomS86KNndlcyzYZzGPZO
DOmNDAEJGlQYc0DdPKAoRDB3oFSTc44HZkCAKBghaDhQhFEU6a+7f4xQ3Fz+
F8N9hSpDBl2/eyJ0SqDzufxEwZRnADFEenp++UMWaCTpMZtqSWVhEAw11KXO
TzHgCQzD5DU+N2Z2nqV49rOMMYlfUN0gbG6fhUnZMxJ6Dj69OMo0Q15kH2fo
eemrXNuQtvE05tc/JwWkypQbV7hwKSoax6qgqV0aGuyXLsZyXyeQJMFv7X+b
qjiiVo482O4kJ4SmD4zN+FsdamSEbklmNALG8ZCy+/9wsjRzLxT/tKGQ1eza
XJDxMr4De91QX2wux4yapPW5/3SzcDNkKJhlSJOZvawBJiaYXAlZR5/DUFMt
2mVSzs9I83d6YGIq+XTYIh5K3A8npTK9xjqs3p0zZ7YTQkFAwhJPryI3+XXQ
l59attO2WgFATEjw9eQ1Bw62QauFbBsBztWBUuNDGG4JqCaQGw0nlXvIYD6q
yGQ+gcBTT/l+d2riFsF+dOE8svQ8SBj2jDSAUPZPHW+bswM3FY5rOIOArqDP
lbxG4O2cU9nwp5EhuhF+i9iJlwabBP6Uf84VGsjMa8lmoBV8ysLKzk/6eGMb
c865txe0QlcTemtcWIfJjWXVhg+SoqIhV9UvRAcsr3xEuZek4wL/1Tv8oq+I
Mzhw5P64LX3QVFEiIzmJXdGgNvGQGVozmtVpiqHgJupEuvEza6eDe+GX/Bny
n3s/Qs7WF4NKtMiqCGbXyyJkM+tkOSlJnuKJsQB3YqYyEYyenGKQfbVU8j7+
QmVfC6EtKlyJjqxFCgF8tb9S+c51lFXsPsszPnJ4iWRtWbKORpvFze8/fNov
IG7NIKBIJKJKIJ/fss5KAhc0iCEOrztUqjpDJwxNMXsi39BMHZiCpNY7xLhe
u17apeT/PiMiYkAL+0x5IVlmTJvpQah81NSepkrux/fU3+x2blERN8JD0g4r
IGLc+SC8W1aS3cZbgKj3UaihE6Zd9UpkyBptbd3bhopZ0BPUBRO0yw9044+W
UxDhMF25Trtp+oim6Da3zxTt+EFqou3My2RdPmPo8B8SRTnJoNhhZs9UOh/7
eDyxYAF2biBoChSfruagrp7cdXgivVza6jbxyQe/xPnTVYYFKI5oLjkFf6wX
txxr12b22Dvf73phnf/x5A6tvZC7NqfCXC1fQ3luY1vaeYVzG7lYHIh80vC0
cN1J0qm620cB4vOW7tdfONNSjtF/a4qvPNl44zlKPW9N1Gy6WECwMz/esYuA
ofx20t36Q+dJ2U1OK0OOxiNaKdm4NwGl3pe+QzGdddbV5qlWQHh3UUdaFezO
8ypLEebj5UQRanHxmLJk5vUQGD9HfQoA93OTwAervnt28T957VavSyv8dSXW
JAg0W2EzzhHOXYRuefrBASZ04ZvhSGAJdA+DmAqPbnExnuMQSfrjgTiuHmiP
iQej4Hpi46xh7rbj5QE7HennO8jQku2ZaUPJ0XgDSbIGb3ATrqt3nddqIWCF
prGsV4PpmRdHLoPmYUBTH9VH4tNK3saun3t4M22dfAK2WR53nPjLs/eaG5X7
guEKbX5Jl9e26Q3X623UiSht5xlNjBpDorqP4hNOoeAvrMepf1zdiggFxAfx
qfFh5E0k+CQ+anynW/yt6HIKpslrW3AskDagXAjL8PT8Z+xKTd+qk1LXDUBg
dbFWzC7d7n+OzkTqapFfy3w5XyLn329ayz1XL6bbvfdtMj10xtKttA5aWZ7u
Kp9L1uhL7tIF8ZywF53jVDDQCL6+zNcTApMRVa0p3WBLMhxXEYSIt+W64h96
8cOdof/M3O0me6TVggYg/3clWycNd61nkpejkvktHb5SWRLaE2/1THA8eIVB
nEBy3Y5Ofr1BHw9A4nS1JXL4fvAgwMYON2NthIx1Dz3eRmSpwtt3Xuuc4lp9
KUo4lAd94g7R8cMIPc4K2xYPbp/xsNs6sqOZ7d7NSfGPBkHwrjZ8ISyP1ECy
jZfa/TxYgF+/IjhO2IH+v1UCuQA+56sbpx3HPRqcoNgiKHZggrkpfZDbRh7E
bXdK366Tdw4buiFCEZebj41k83fa00faK3sglYKDvdXeea12ix1bxClGn+1a
J1scOdA5WVUM6hiKRaEUiG399SJB2pQjsjo5kQPFU94YkZEobf1HyL/urTAj
o+WpO7oh5fjZRFH25yu04JPRNAVaTuRPsvgBZl8wg/QTDfk7tzvCJ0LmmQcP
t+wNVt8xZsYKgB+dl0lq/5+8P/RtA3EJKEjuGZkgE4aYrPdNyblQUGcolUJG
puYQJwtKh55ZarBpyHKY4DEMlt4uG4So+ti/8lEHzBk+1FnPdv94Mz5Gdzsd
RQQJ35CIKC34aYLO8d3GUP18OV+WLlaKfdNDXxPeHiqcdsx+p+wZN7L35Xxg
jEcszGpaaucLTUSAwRvknNOpXXa4LvLRwNxzvUgjOzY+xM5mDhGEaHn10aKg
uPhfbXr0NNp5k1EfwnXV+jMqkfPMIIxL5HrXKBX070GP2CuZj31FY97Hb/QZ
uBehClzZmbOpMhB7hjVUsnkLQzuOMPLSaDm8luox6RkZZbTJLwFogDRq3TTQ
I2zB/Y+tDNZxAAfE3h/c7kOVIi12h8V2zvg/uaTHahtCh1lfjOMCA4/OloMt
YPyBU2824u+97p6A3lndyI4hJtonR6kXXj6bsSQKwveTavyRWlmCAYOOYRAD
/zyHm7q0NcdZl39Vj6mIOIPI7B4Ib6z59zXM8vv/gTCWc8zZ7LwdL7nL7xAF
YHAZkoOKWR1jk6lRlP8f4J0E+iM7HR+OeTNF2uGTOSGSVtKomWwcPudGgjCP
IGpNA8Zu+8sZUe24LEfgaqL655gZuvUYC0R0Mfe5vv6LAQsNsC/pkWNbnK08
IOkVBvieon50DGHgwXHoLCUJfuVKuHz1KAb8Cs+F1Lai/pxHO6jMOULRXDgO
l0wNpmkNu0a5Y3yVjyKJvScwcVQK5XdUIgYNmIBc2fZp1AI3cTYyyS7+v9PF
lpq80SAmnD1JUsDKvbdfCqpaH8JdByKLdd+Eiij8YUWEj5EK204VFo+yhqss
2xG3bf0kAqUgQIbkWkaKYPgDsc5ttqFuiiTE6SJAm4o3JfaTtn/CGl5W5iNM
hT7J+hHAv5TrFZWVQeOeOWZoR1+Z2kC27/hGxpLeF544xYRGsYeFSS+19+DO
F2wxxykD31pSBXEjXBhBmt712TB7EpEcrFODEJZChkwyQkzKGXUMaM9hrL7t
NdWN5UukSt2tQPfBocOxcjLl1WRKDtO6erRfhIoFmlxtrHmCwYQAsUmEXZH/
BhziDhP5M9IHoKCEeBp5pWrqiU5EDQ0GFX+i0ZIm9Ae8Fsvz4lTaCEhABQlJ
OoNg9YXM30hI7qQ2oV0182oIqDlh5dkr1NHdftHYzhIOFE+EFD+IUeMVXbce
RkIKqqEuFMh+rrkY0IByduM+3srtYscLscuTsaLF8kxX9proyjG3LOrBZIlU
7kRHB4KekzhoFGx7PlvnrgqgdEHVVhtpBNE+g13IUwzosuHCbFNTiIX2Me6u
oWDQaFYFFQP2crzdhoru/PMhSxm1Y04v1CF467OtH40Bv6WDMf3u1PBBsBwV
Ey37Lx/nCruMt2OXqlZR1pwCyZrizNe7s4/rkDP7CI/vgB06OebyvYb7qPDF
KiKT2+fy2EFK9KOwjtqJDNOicht+sM6pWqJ+vMgyXFkZl3oizaclhOkDP+L9
zaCdIbwV/+V1kFhtzZtQ/ffnCW0BQJTbAgk2zAbkwl6r6pPK/ND9bPleceWZ
Bcd6fwTppxINxajqW2giX1QKL7mnwlqXLnAtgPEwF4usS3Rb9U6NUR3Yc6hN
ZE0yEPDb6Zf0UAgXo11ppHZJqGpr1/SrPahyuUBHnFpzcXyHXctvABfAIPi6
upf2YbjQ0yCFTWfurR20ZoLYu0Exoqt5wi/boEdx0T+kicDbx8oHCLUpjJte
F69RzmaX37Q8Y+X9qRrignPuxcXuj9VraCFNKPqDFXWWoSuqNFalF63sRE7I
zAMmQxBqC7OE+xEBQCrH7VHAd2Q4AqejoeFsaVPGOofjlz525Onpop0BWhgJ
sC3By/zlJQJZRWlShhe8VWgl1WqcCBWJwwGy5UsO2s8APNVF82SXHmsEw7Ij
EcAO18LGlGuICWGkh6ndwH2oIb4dd+kdzuUWlCJ1TbkVJNXH+7g48vFXRsRP
QzLOd7BPsLtQ+bwHLYCraggPzB7PJ9Rw7HZ/POk0zFbNmahwH6li1LvyQsab
i2Hilb9ucavuLuiPXGNdIEziX9FqZiBDlAsUKk9L47WWtsGhKSOujpomtIdb
cyGlqJAOk195xanrzLT6hXqp5qa3+lseFyiXnRRdykCy6QRwM4NIMIvcezXy
uDENjxb9wTqdrWrOs/pYEFyrcsCdHzrTNcNg3MkjUCgRFlrpUJCTtGU06FRG
E6B6v31vUSwd6OklRuGKVkY908ol5wuCrXS2V1Ege2gpsAnCE05/VdBm43i1
b2YF77F/36OVPmGL3Nn+XkAakngRs4SnewfcVFawzZuDjv+MiVe/CzpAQM52
v2ul7sXFaKOecZ0DoOWz2JL/oiOJAeIPgmsC/lP9Kw2K/zmQBa8k7KTxm3S2
bhNl/O1x4NRQkoRavpC3MWrifQ7KxMWyngs5T/nh1SJE/ly+Lg/chxL9EG/j
NRRUh5PEUTR5Xt1xe2Krkw2aaz3v64D5ShOw/83/fnDsvQMPTA84+grHRmAp
kQuYt/BjGNTzBJvOhaBdkiaXhpO5OFIRf2Obb9of1RP+D1W/qdF1LoEg5Z7N
aGMtbqzEw+a+4Kb1FaUVqoZr+tFS/8A2IeIS0AuOJi9c+gcwvWxE9/Iq7pi2
PqGWcZYIAQlRcSHdx5AAQXabTUrqyrxKwLBT2jHzhqVDuvP47nP3V1Q3WHHO
w0+71b0MLm7hP+eap6edq1sPca2SqtpyFDSrKEJaXor+JK7IUC803/xFY9+1
CM98H0SNoJXs60wQymqh5a0zkgGzpECRvK6F+TEGytKsrk6ptYD3liTrkYw2
gCu4Ekpk+Rxw1og5TS3HoFKnfxN/maB2Qmxb1ID2xV1sCge8Ft5PRBhy+Hza
G1v+qtTB2Qy1KOe7930ZkN/7u1WN0/CiqQDKu7DukuWZnNzYZSjeElOj//zc
T3mPswq4M7aIdJr4pwLH7H4aa4pc6d0GzI4nmSApVYszWLyNIPvPr/goB3En
6Cx3QFNVYrnS8k5yN+8THp6kzFnH4mGB4Fea2Qtjm2O86MbCn4D3e7qWDdtU
jlp4daxZCpCP0W70RKk8TAWQGhDqtVIrE2U+vCuCnF+HHWwo+Fa854qf6e4E
IMiCujYAs70rrJZaYU3b7Mqf34xbosf+z7gYH4YY+T7R0HU+MNaqz7yVUnNj
N85WKnYegZNhiPlFD//q+m/wNvDHefRI+iByLk3LMjmAWlgUwG3ddtFTYca/
tn+MKw0fIzF+8vk7fequnzqoWHBZ0TwDZcLzCQRl34HDYhVVP/DNPkGbvIAR
ajlE1gA5xnFUH/uKxszXcZlMV42333dVnBZS30V19dfUSJGhJahc4S64iXN0
2/SmWVy1sUptKfAq0ZpnOeqbbERONNHG97660Lq93ho2KvwTN6WXVw78pH3O
9RCBs83X1/IrvTg4WKg7C6KsYK79ksKvqwP1R/JlHfY7PsVOmFHdXictwY6j
kIQqEkb/i2zHQ9Q6hKKJjHrLqsGZqIDIrz+80wIzlTFI1xs3ySHvVrnNZu9N
VpPbswiVeF23Vr7XdWJh5rqx4erLRWpB1s9ho0tS9q74f73COjOH+i65XQo8
GU+HCB0C2BngecjeRLNJQRCCve9e5tBZmeFfIHgSHp5a5dmFQuOFMmm75PGH
/kQlJaPw75zikqot5kUyUze37mgT2Qnz/m97gqWs9Ju6ZKny9J6Gl+gzqBmm
FrIA+n1aVbQesxGPxE/fYkDAoSXDiDTh8R+aAbkk7a0VsAjz1VcCVPh9nitD
9cdm3OJSIHEYt3P4snmaItz6uatBdH6aGz2DaLjH3XAaqq+FFptpcP0wZcHg
0TsaMee5RjDLEB6dwCLY++XB5qHp83j5oEygbr6KU6GuTsdFwfVDWa/Eaz/c
rHLXjcLNDCfOkbdHWjggICGwEf7U3VLfskFCSzraMI8E66RKUX85qyQsCwGN
43QNWGac7ywxfAm+tQIv1wRH+j//qh7SqsFVu3Uu1a6KArHpwC5b15Ray+12
04YX51bsLDg5RnZ6kvRY7l2p+Vggbwf2ZiHAExI2F0m4KfUNDHEMUpx5NMW0
X1FuMnp3001R8uEyp78TbjyuCx1+uobcRyFMt0qoOtT/TaqWXRHh4oyZs70I
CqToT8kgQtj4m1YT2DsHvtbdHv2OvGhLzQVQ03rwTjYSpDmOiGqiqQp4ZGgI
szrmWGoINlLG2xwQIkrQ5OjXwkje7k0EvKN3U7zUzBsMeZZc2fP/kNkQ7qFW
jcMIZ2hSCY1j30UzWjk+to7CxJ+62xk+r3EUavME4dOODxjtuH3KV0RjjZhG
RYm0grA5ac/cYxb8mWd2YJtv31ufFHyFOIzIdVASMcIF/ZeWPzZBi3FFR22p
F6l9FTswoy9mrmMy1o0xmGF/iNV/5P4tXarByPH5Gcpb8XxdeeXkep5GsLIq
yBFm/ZjVTdKND9D9doD0PpvBxmYwSx6DZ7hJH8KDtsu9Xg8no+ThLdZ+1tgm
elQaPmzlpTAbzU7junTlOJjWq7T59nTZZHUKVLB+nJBFPMYmnp0C6QnqDKhN
/JtLSqjRXtFPkyHsCgGm0xitnMxJCvquzElvAJHAPrWCBMPHJ3xNc0cW7gVt
JYwYJy68eoRAlH03jBJqoyjisY+2g3uc0loSNmoqRQjrTGskEQjtFT4zJe8I
jfhy/pR+JP2Scge7A/P0at+Hx4x5DzFXs/63SBjctM3QZwTcbuLNiYz6BKr8
AwJfO/O97ymSBMqtqdr0d9hQEChPrHj5pAUmWEyivCMAdHNWNspybE6szWLk
F+LX2Fk9Vk/FWtCPV97Y/2kiRd4VWkGkxDli3CTUHpPbtjKjECJdEEGyKCP/
Aa22B0dc9anTkrIe5A9YfX8lEwEyWZBHfu/xZpXpS/Quh3xJQ2yGhCWMflXD
ROMKU9JGC1imh34F1Ss2HFFsITvv7aVv1NB5Ud9K0Duie7DE+J8aF2amzQdn
GZQcliXaECMJSkPEPEzccTu1VKFCglPN8QnODR1wD0MWTR+Z7Cv/+nSSGK7E
Hi0hGrVGV9DAazbIbxEwSJpQnwhzHWWTAZXB6nkon6umqe2GrSJ9fCRc5Gsj
CUXg+ysxKQ/OdFvFoXZXJNVFAMSSUwiU7fXFihRnwLeioUmPX/R63GbfSe9q
FdaYoIEPSi3yDFzyTX+9SFth2cZ7P0/AK7hdZEQtjbn0T/RCK5GWtXx0X6Vg
SABio2vsZA2IjUzyVPXZ7p2liIBk2+nzZ9UVjxWnTEzUS/AgFB6JJO3+bVg6
Xm6lqKnd9B6KU+xCVxp/GOcfDJT0DsNNZiEEfXzdhA/G38M65zw1+LER2JL0
kJNvcb8t7EEXC3C+aRcXtYCN4u/i7G/v730uvZufB89j4WxHMKZE+VgzH69/
ERk0/G6V1xHzLpmIemdXRs1TQWLiiAEuHOQYcrOTwHQ37fUf3d53e3V6XcSO
ku5KmHOG7gV7T5HcS+4s2mWrzUZ23RnOyzfI8XFgXWb9Z2BgqxnPa+iAti87
cKhYlgwlpXZZGAscqr6ZicX0dFayXWk6q/Axx6x8wD781u4tGr5OH8lU/4Ta
RDOxEO0g40pDXKWJW/R5Bw9dKLf746TXyFIxgPNdKvcpWS5xS8wjFJ29mDgZ
nS0j26Zbq5H+KOzogU/PXZYrWlTezCLNcfabnvUzZzWdWQf/WYAKsldWTn/2
TQleubr+FFdOCUvhmMSvROFpJmUMRKmYUiyCtz414paIOvr9hAs6Zv3JLtKj
RRJeITGsVAS5I01ewXzxrMamdap61R2Up82iiYyJ8Cm3bU6q1MebdMX48uiI
H9VdIgx77Hw/t1t9lykVBHo1A8WOgvjSGzDIJFl5x2232LBtFHoKMd4OzBuy
2uR0MLKWRgPNM+6YjbkOiUopY+3rCW5yBr6Vt+m5mpVwjEpwwWKg4Y6Hmlar
4MgVvoV0jX7k4gPczSGSwgd8ef9XeoLOAlNHZcoR2CzSbmP3m2mHu+/mO8Ij
cs3Eb+w+uGZC4ff1xEQCVvKpEr04rNUL11j7cCKi6hc+tiNBYl1U6DDIFu3+
jQyY4J/UIKCSc+AoNmpnBuMxHg/tRAIFgn2VkXdGPlvdf7dFOOWjQQIZrWci
vz3tk7dYPGxj20k5fzf0103LR/zFsCF8w32zSDBeWQXjvVCbHHg0dCkJRpWL
R1oSf8v4CWpXFuFnhIdunaugCtbBy9VNboFYc7e40CufJTtxTF6COLg0/s5q
cPCV4dAA1NZbkrvXV0lmrNXwnGmkDwBJIaVFwyvfUfAZp56uHDPHlrMarSsr
Ef30K8TECBo7pVcOJrQmYny2APB899YxZf2Z7G/GlSCUQT4omoFugcVWh19D
chHWTryC2MG/DJsDL3cBmLJq6wYnVHiuIFkyITgMEGHi5P/whFa41cXf36op
asA5leuk6cwuxXgZbtKlltOVGX0NLvnx3wev8OxhlYTEnUsF78fP8r/NDkkl
2JWK2SB6cb1Z6Ts9xL3DyCvLa2+vz1CHTLw0G7IfMlJUYZ3CpgEQRpBdmTkD
lbX866AR1aBcfILbu2S5A+FYiCKR0gaGtIk994Rgi/ae4omNBhLVlTmS7+b5
00QxyjijNCoh+ECN+2F1uhe13iGDF5FAQIjss07GtLUIHVlWjIQFRhL9e9Tr
5om0wLfoEXm5X5oe8fLp75ut4gaBWOqHafDrHUdrXbWqMJXwu8Y6zRjcUnG8
i6k1O06NOdb29YxdqdmyS8/v4KpUOEfT2X0oLcgFkgACHMd30Wjbs3MIgpUW
7OpH3K2i/ZVbJUfhgDxFDwx2YivyCwPocKIKwIIuHBZpXj1BT8wm/sBdEpES
wy13BNBbmZ4W7UrAerzaRIm1VhGRhy8ovMN65fJp3V14/AvnV7Bker+ferbY
z1awYvKD/bRyDP7Vau//EPTlLCK8lO2K2uyMHVJBfRrKRHHnuLZCefet+uBQ
7XtVYC3kSyFd2nLup+MWvwjhivdAK/MAt8FDoxXRb0fby49BLuhWa2q/OYeN
J68lS5mnmyicMAevzEVXlAJEpKeQjp0cjioC3rqn3H3vaKGinRpuNmB0giTf
QDOIUP5CXh6+WUjIM1NfqoXWlgNOA9EJ5kH7sCAao0raWXPYHcR8tlWzDp6k
TPdEqvqW/yeT19MxaqxLQl/D78rqQjZMR0BbVbdpi929kW2ZSptAg8vMw91F
g55/r9edAKu6srMFNyG0QI9j4kxc6pB+LfofRwd9y0/YjsDaEF/nKD1N1Xkv
6hjsVTkw53eNwAxVqhn2G2BiA0cSocFyfnIHGAdFXEZ0Sx3te+T+oQqn8Fxo
qkDjaL0fTyX7UeuI+/PGLQb+RD13NypnwtjLjPjDgjpk9C9YGP+kBjSbiWJj
pPaLmXUSGkw9CQGpfhnQXYPoHh+YVk9M60OvFvvDV3u/4k4sNeQEQ0o+PC5R
U8850d2m7gl72l6RF4D/53BNgtJOwO2DWI9IgUiE1WaAAuuXn1Q3OcGx/kKM
AidUYqZ9nQlpptBKN0v6L2NhN/Ts+MGHYueodGzXdYdSq1Nm6ODaIaC3qcNP
b+yvGLrYeDwprgNzvqfJNrw1tkyukEmk9scX88UjX3um2Ty9dtSrlE2orQbL
SnqjbB+2Yq7y+v0dYIiNtBa/NBNhZwewfRS9G4cOTeAVxuDUE1PJfnl/osDw
mpLsQefmaQUH+092KfBEHG69Sq9bQ1nbWvynwe0Q8dEqwdg6QcdEztNfdAqr
iZ9eXb3rhSWtYRIM3QLFgYNXSp0ER2geg4J05KOK78jKMax7tzl7ZyOLeGJX
Zq1bvGyUQMaM+/cl+aT5s6UscokOgz5wr/nAQisbXgFt+w8rgKr7CisIdWpq
xgxfYhvJeuR37HVThaTr8b7lfio20GsrbZR2uhBRaMU7WHOWceYxsJimaosM
Y/M/2eCU8Wb9th11/qugnJjenX6b2T0oghcVu6du/yzU12cJ/GYPKmYkgy8I
BI+X28vC2bTHTJqdOa0d7/5A4hw2d3Q0759EzTr7MHttC9DNbuFfwZdIF5pp
Uubp7GcrIJlU0RKlHs6NuLzoWQDJ0mwZZISaOe9sqf86Oq9qCtZGbv5c/wNF
n6JQ3ooaVIXV32bThxq8zyTnTXHlm1siG6s4udoIAtgsx7eap/Hif+mZq/T8
I6WbyE1YXLH1Luwi69B9dMYeZXhpNMDdbWa4Poowhc34QCemVk1Jn1W4NHht
SejatB+YcO3+H9Be976RqdSSoE4rGdN/YYpYBu10sYAN9xQYmvEKQX59+hBV
ejf5frPtsjmU6uOELAj30XIz56uYVmATocjpD4Zeyf0n95fEaRG2z30fQmOi
+P5sjkk1NPY/jL74SLQbLM9MZchMtr74vKQOm8am+C7upXnptR/c4XTpKL6c
p8dXEDFdFeHzP5ucCeZc/FuqYsqqrNPh22xDDdi6wHsyzCo3yZNCqGouuyms
2ClVmHGOvPpSAmj9kW/usU79wmJORZuF7GxWW1lF22HfrE+LFB/JFAIftuYC
irNFftF8fYNg/Bzmz3nxnXN+JQ0CuWL/Sg8RtqTJQXWJflq2nJyaUKt8F+CZ
oVxprVQ+QYx6ya3x8Dy1B8LcJ9Tish4mX/7l97Y0CZ0h52V8tD3a/m3F64fM
s/tIlgqzws6ccCw9hIxgmUnagcuqZ6+lqFzIGThMfBHnWXq9SIv1oElKWF9H
KZ2LiQA8om2niDRGjurP3eiXIKqmws1IJFfvJk9ouWGvs8KLVZLQlkx3xvY8
dLH5ygy1r51+hqSQHQfmd1AxIdHgY/TtUz1niPX8qFt2MIunDnP3F/p4wcs7
gZBgX10v6GNyYmXw/5jndvekBS9vM0Qriv+L7oO3TQefRTmBw42OIOlXr25R
olk9lfah5+e8nzsagw2ObAgZ5+PNLYj/4SlGRqmwtySWRCuoSitU0uXwUwDh
SN8zKev0qdxdafgVD0vpTmtxhufRMsY9xtVQUdEp9luZhf9SCIOhkByz1xSs
wXp2YuT9CO0Hgbx5A4tOe51GnLPfR+ew2RIgWxQPGWPg0cJOELJNUAq0j5p3
lJAA8knG5bEwz75cjHTt4YBZ047vqZlW8mIaVz+/O5fUJNBa6HEkmJ6couEn
Lhz7mNdbiUa9TtVpNuII7PUpZyQ06931nycVenwkJoXQEC1UddqncVC5goz/
s/ofdjR1nPkD3+f8BFhy+tmPd0kCQfPW7Ybkbtzyrp6TKPpagR6VnhFuisJF
ERLxD2j+0/uwBUlmhBrlZUD6t9UKvy2A5GLhnN+9VDukk3s9tLVafIAMADwo
8vMgWiGJZKUqov17Gzws2zcR9rQd4Dpp75Kb4xegcCV8PdDTlXBgczLvMTkS
q/KwF6pk+hR36jeiLdoHGrbJyXoBf5loZbOMNK69rbXMjbQ52fTSApRfKzLQ
FEV6OtQnmOZf2QxmMcf6PFAyxTeMkcARmNPvi5ABmNozI0POyMtjFhHoWEt4
C1gm2GKGhNIEIbKE67lW+Co85YvZrd5dD0j/B3+aE+QzVQU9SV7DhlMSG41T
R7Vba2GCCAEtw9+fYstDk+shzNIQ+BDR2y4PDDnK0TF5tsLDtgc5zqIvyshI
OCF7F/cDEarwrL5+bnq/Weo1jB8bEOD+oc/9iZbyKGyr0bM1HrDiE7MZMhe4
sgI2JG3HtyU+KENhF79RIkY73lVl3r5YLNjKWjh5p+T1Hm4Kfmf2JqZch9jv
utghpBaLdeAhgBYtNS+xwFf/EKkHcmGuKDWiWnAW2mSyIigTEP5ng8Sxb6Bi
D54rl0GfoXfpRXx9+V0o2H7sJqe9ccfrV+HKXNk5TtvqStD9xSm08iTPU6/k
lAp42TlvTAr4GnJG9L4nOa9sQHlyQ4RVmRb5MzCk0PPQWf75a3BcT8v+m1Jb
JWdYrRZWY8CUykV8r+kep+7GBOXhD7JIQO5eLZvjg63TIYmGEhRqoNR/5xfy
WpSAlmTl5wm3/rM+0EGxtHPS4Wu1EDPlMIOVUe1e25Zlu2XnLd50MQNDViR4
FLWC3jcurNjBLqT2BUJmYV1I2ggKGqpErZHUG6vQulpLXGg0kGSAGNK3Qawy
Q0yMERcykmqEB4TIILlRDKqj+6n3jQgZl4c6g3QGJobJ6CaKniB9WKAK5gCm
RivuL/D7jSU8SA14+VmpmkkKmxb2/ORMgVR1INVWcQZe5eiAsI/k6uHsrX/b
eg1bKORjtWgs51b3noDoOLIgiV1kk3nDqYHBmQTLZ0ERtB0ueS7y6oRbFvMd
HY2/ZVFO8llD3FCb1d2XLT+DRby1UQlG8nTtRMhT7aIj3YJg00fYOoHv8s5M
Aqq9oT9USfLfvCQfopHm2kuWpXpo41pEjqEqLwKVLNIKZpD82EnzIT0hkhpE
NrROY/gb47sST+LFYWajwwptu6l7TMnOHhwi1LuwAzYIszCw0zrTP+ggZ79x
PuzkxZTZavs3+U+xLbcy9bxamrWfKF1gOAsIe7cAEzr3+oXDIyd0R7nFgHMO
snHtRzQjtgdCQ5IfL7n1P3vXtGjw9UaWI+eNrzEswnI/oV4yRetyqhAAgWFV
4pJdiEIuWJUSA3L1u7VBWPxiZalyhHfznTiv84l8IF9nXfa/0JKPp49fFD4P
Y6zgYperTVwWTUDi0/d6Ko7drh/xRPEzI8xuif5GeC0HVZaIDt22cWBOBl+8
k4iEAkTSu5XEBaFXBkUA4vhQJVikjdP8nIyUwEbJASicycwKIR45Tvrmb8m1
fiibtvbZi120mPjBhc//8cnUW4jszRa9Mu1EO8A79wCq57LKwGswNnGjDMcV
lKVUZHtXF/jyksKwUtRQdPlkvSMJq4E8HG5HCLNBvWIFK+KEqfJ7I3W8D5s8
Rs5lZaZcVEqyEPBP/CJVL775SA3bUz9aQkSuYomrdPYoe5bZHg3Y2ZPG8pb4
XX224I6El/o1umOmqdOfTD6Jp/EMLhbMrGmMGCpBmpxsb/7FJhE5JBgWaIUj
rI+9Mn93XOrlFq29AjW/hz8Vm4HRz4WetNwaUPYuLyI5wrQ3mwMD7Wiadafq
1YyMBxnhRzUQehY6opnrwhNsbc/rgX59CpNaJ8m5mco6Yy4b35hHCyMLvpmI
Q9CvXotKCWCchCjRxfAoTXdQT/aSCIz5McrcQm5WT3inb76PBI3QrXdEMHRk
tE0QhEjHVvlgp3FZLbtaBFP20DHXiYnLYMh9i55ICkR0dY94cFnkPRahmBXr
R6Y7ZsQYhh7fXnsXvUYwkGXSPHRIfdzxGi2Df2PMKXxMJphWx871gwAjUF9O
0l47efOAH82sU0S7VOSlpgaSQzdqbwgwfKbaosxy+lUdTfQZfyz3V6eYzaMW
acfcLE3VZDaV8jKDl0N924GH+WEtYyOVIDaPxg0rS2f6BzYkFUy8JmWuWWOi
sEyzxQKNRhn2xqHQWOSIpcPazbss8qTOe667gDrGqMJ7h8cszXFJbQA/O8Vb
zokYIfAwCYAlsIsOQZeX922ilYMbar69ZtYalnz+i2YXwx5uxG8pV2kgqxeM
9vgIAGpjdpEhXC/vuD47vlKIx/NzKq2wPvJHiBbFxneGq9EOC7fvBnmL2u8g
9sq5qO0GqisQsjlggd4v1IBo2UuEWR9mvqGU/Hs/koE+zBDO2/tliQHdaDGu
bO4HDiNxImZrONTdMIUzdtrTnxff3INkoosrsgAGIAr80JFcmPJc+2hz2XdQ
6OAbQthhw+ffeCCX5iOrO58nIFS0h1HZTmyoQIIoi5hG8CqVNwUNqk5uUZW8
+5aR7mH2QC9O99Bz6Fz5+kuGWolwnvMB5qf87IojeIcMyrxjBQuAWXm9B/kI
HQN7ZGkxOS7dHgV9/fR+xLZGEsJW19a0gE28EWZQaRLHbLFMfNgJ1BqK2+PF
xUzLSZWBGDkG415ePTlNValwVVVt45YcNibNJub+UBaxjYePx2lItGLC60N7
bWPxjBcea86gH0EKLTpgEGBnLK8jAyFQUsn+aReWV6ZlwsUyHmlZ/0BAgHbm
wuZaQ9Jh7hjVj2rJ35biset8jwWEnzr41ptor3qOsmbmw2FE4tZu3GkY6V2q
oDF05NCHeGRgyJEnC+XMR0uu97O/LzRJS3tsGaTtgT+DRCZDMEaKyj8jMcgN
R6ckvmvrVqzZ8JP428JO7iqsfGy45ERtxO7yGNL4YPflEa+MDqMhFBg47DgN
X81O+A6tz3uWmGpDE/9quWKxHG3rWPac22iOdSSljnklcJ/pMBEVUymJYqpA
aIAmecoXqTSBhRBi3en7WviHTqBiAt5NUOfAnmdFT6C99Rvxc3scfjQO5gJ/
7Ay9mtl1qdWZiYFf40jY8Br8srlcOosV3Vg46A6OP0rp0qXnuKBsYcwNMrYi
hqlA2nZb2bn6dFqKJib4h+TRzJL0U3HJ9q7KzbEQ8ePNXpl0GlI1Qex+GmMu
c3e6cXel0C7gEySotDobCrJiyZ6yP3dq6vTxduaqBLZTlZ4W4+hFc3208NcJ
RtMb9YQnoqVTWw1zvfcIkwO49qWWo+aTkHkGbWt/12dEbOg5cLFyGrADHK02
yJybxgbnj8iYSJHRMQqDSRIvPSRpERXnng9XJ7CAimz0z2PjAxXQGfOEaj1e
ESqJFdDNDmZ932JuRTpxT9MqRfdjMYOS8tgwsd3HvGRHuSl8Pnh5nxm0/U1u
yB8OJirThg45wLsviMQdYcuwQd6e300uyIF+eOYjNMSNsw8zaDNVtndJMNXb
InY1G+5uIlolx+OJJYZGuudorZ4GCQmGGAemc84nWNv7aRyvuK4hqoH8CqRx
HuvWSeq14r6xe79/7lftx/bQ3lgUQziZlklHyGOrF3NME1Ee9/ZBpTSrM82n
TGPB3d2cgSQFaT4qGhM3BmWZJq9HMKJmm+Yglse41YwG88hK+v41P+/NNFGB
xcIRz+j3NT2vW6dcGUpPj0IsulrAyaPj9SAA1XKtBDtUKwO2nlrrYPTWKyZ8
Snxi71pI6ShC4dMDpWt1LXbnLzSrQ+fazkmW6zX95ht9bAbFNv7CTxL5PfKz
T2cLcIeS4n3E76qPK9uF2++U45CFNYPhmAJJsWRCI6NwY5k4UBURXBhoohDC
Ez8w2tAKdnGLqdqnkJsxX1ZRFF9opRl85xyYvPNl+CbQbGR2PVuC/LC8GGqA
bRs2/PWECKWhDajWzWEIQCNx0IkFhwgp5/CmxXTtsM+42X0RPkeUeU5xUF+d
pu1fyl16X/QeWSqSyNtBxhiEZplZTpF9GRm+gtpClRCTRZr1d1LZRCESN8AO
3cnsMVfoNh1pzZkmCZ6hg5zpRAMmfvrTgBDviK5PJdseRFtKXbrOAEims2cx
ei3vbVi5pbwYkGlX05uwIwLG0vdktMt426Zo7pGN9zommx3TDrgeofHHxFsM
lS7J70KRSjRPbo8PFuxtpc2zOrbzOq9DtfvPFgthmDTwVF9Pwex+FgLxk+k3
UlGCSAbpen0fypBeqp+J7xjTXEYpL8/cVYOYVcN1YTjVS7uerv41k7LL66f4
HKfY6G5Fs4dodpHWIXkSSTVajEbvE/Y8BfWsOBAHreKVvr8UqhkqOYX5lzoC
beQqL3uO1Obc4DGRl4QYzpZyFFe/k9AKCe6Rh5kTJoIyOk1mY1uVwVG36rNA
Zkzz7ow5k4byvHxMDc6nCQHg3YFBl+lCjamEMEs1/xAkuU4oRJ2XS4FsIu1w
tqJgWyGk6roBmsdOwpXUfQcgUROXAOGgZ88z+jg4m6qHHXoZTYHB3msezS5w
A+S3O1lK70U0OHiAPgNPpwIxtDGBO1VHfe+pyxr+u8HkmRCkkS43Y3D1UDnf
Tq7bgoCDPkHcm0s65fEuu+WHvt4Rg9wszrCpR4EBvJ0lguVB3khBDEZP4xMv
KTo/jsIECPGevj8CLjC0yWnfOxQELEOpYsa4ragTGLf9T0jQt1cgP+iAs7t7
UqqJd8dRzyJWEcLFshS5345/et9UEFpUncieXkZHSKtsIgMHeMg/bZMRZEkW
kMIclqHgRA+7msys5iStqX+TD6E8/PgPgJAXNL7b2lrqP65x7dqOaxh8MA0b
gB+keECtcv+Kk2tTElzTnRpPMfoWRce+E5czMvRL6I6Uc6KVthS3RCj+7Q41
TdYdGM3/zDUZAGoyxxvvPSen/+/ibRYH60967VI01JACuK2hX5xah9UiP/Ay
5/5iJ4uwIY5r36GSIClX+E8QsP1QgG05wL+fpHaQqHK9FkNVZnLhCBsEAsFi
8TtQfNSVQO/G1JLQI8OrfET8/BHM7sW59UUYnI+imFLn1NpMH6oaNQmttZ5C
ZfAaSocRTw1J2pP98YbB6DF7qIOBVmc8ydsWLKXBpkxrCCcf8teffy0raRj7
ktWFfQXdkBVLs4EwmvQqUqLIT/xH7p6f4PV94gj6cojqbKzmd99WaOMQLud6
nYCXP4xrk5rQdDv0v5kaSkLqqrecVFLr4Oy+ks7OlAVttK9Lejnncp5UsTt8
TzzoAcs3cX6cEAoHFtJ+vTsJK1Q2gV34tEfZQKA5loB5QXElMk4g8m8axEuC
USylEWlgwNsdYUDUcnuvMcoiqB+6S5/uyDbUTzBIdWZLBsDo9m2DGzkBejYW
kgVm3ei/KYBz1vywl/68cpN+1EU7cnQqvvGnwk2q/ds3AWRJvs8wbMNXP7tz
MHLAilfjTOCjYKPXmpwT32fIBaU6+jc1xE+ElIydrJznEnwdpciqpoEu1QZp
ReM2oMAnCm6R4XRdi7nFYCCUkxZXFaeiRohk5RHeFE0RR9G86Dx5b9KJzYbF
5gGx30oBOwl1zam6K6mzrAcXWR3DHkjbKqiCAIYAtn19CHI1O8roG3UzpUOD
o5Pj0Opx39h0QDT4bpHe6Klko2MWN3InqZM80bygoNRZfwZh0U+yXXL9taGN
ykYqppjlajGCLxEmxBhsjJtlVGaBO7E5/IeHy4Lioi728pSJMGKFGa3xSDjJ
xufu3dxi6s61EuIhOGcCotHHHN5iCwfIShrVyPxgn6I9HbpsSyzkk3qV5kVG
bj6DYWyNA1+TZ901Vgpcf/dNLLTF6Z+cuLr1YtD5oIWNVxus2CVYQ/mKcm2S
99OdfKXCtgqRFZ/my1uG2miM08SoZXgnPKyHPmnGGW08AZ8DNG8atnk0x92r
sHOudY81qOzIV1F1yLV2bb0DgkRDwuFamr8B/W/nGFBZVkaqCFrjKQblgESo
6hQZn1uW5L6YQWLTZsko6hihHZUnQgszi8l8QoPDVZuxfTMI/Sm6AnCSSgWz
RSAHsDJ1BT+y7Oq7Mfl0KOxe0ePD8Fif5iuATQobc7HUs25IjMEbAMX2Cw7d
jWuwzC1Yc0qQAAD1B1L93lGsXmPjJhF8b4ajJ65tcvwU/nwAyao5bIgyrfR+
Jfti18ZSh20KCXZl3mSf4u8J3ZTg6mDcdC3EMKCPZ5YkCam14FfpMzumF3vF
uvfSavvC/ov2ENrZbsuNvcmQp01J2mJIq2cl+zGscKYwKTZs0HjEZ6dvH5cO
70eMttlOy0z5+ZNf/ZHNkFXl8SDp+im1Mo/7+mJgBjhKDkg7Po1OojuQWSM/
ktXwikG8FYY+fd3XBmiXY6cDmHOqApqcL/4jdutWtGyXbWukFn3gI8HjknLP
Q/Tu1UByvyi74ZmmAC0C++/0ktE49WrlMhLfPSOiBJuNSibWvWS5rzH8+2jm
XXxhrUUiulUVN7k11op6aNzpixqCwuZT9ASBc/FdW4mAilZbhiYQTm4Yp/uK
yc6IP6ghpZEbxE8KWMtpOJtj5q5xPmmtWG8K8VISrKTtvWzvBlwK/wfEfCSv
MrydKVX/hQKseMsSE2Nj6I+IcwVgGOxAQojiLreaFDXjn+iIgZtiVMbe2NIv
fr/eYjeH+570pbUhfz/kT7vw0p1k3iVHkatdX27sKLv7VoBTkCtFTJ+TZa/T
a69oH2Qt603iJEDwPuFvPP/K5fOX5RhHGVDNTfwH0o33Y9I4GvSiHAH8P386
3ZYvj6NpW0CE7rZBC6CJV1c2R8r8JgBIV8L4KbPdYuO/R5I4d+md4NjoWfZh
MoLbSo7XykLC7UJdFDg8eI9e9X57/WJUwIM2m/wxDkYZEaHxqCGpMZUcL0a7
csE6YYGcz4gkNbr0U7PTvtpwj8Lar0Td/85rDguiLglJ+8F6Vdlax/gQ78tW
Dmt0FXjYupIPWikOmSbLvhzCifZKoAdgllLAph9e0XewBUzMh6KMuB+2r2a3
xBn39bNsmUkyniCIxadRsndd9W/zIbZ+1ujOCvZoVRoCMU/2brEZwV1SCWak
QH0o1KCHv0LtLNw9v/nbld0JdqOsJPwI3kQdgmMxqL9F3ySEWx8Oxq4bwcV+
Xt2joI2u5vP/vIYGAQt7URwI8/0fAMlZccwKVTfZyBxva7FTU+FWpMPSHobS
SATd8mMqNvUfQxHCQ5HRiLc6BiEryVrNtGOuDxwKPvcOp+JYccDoL8wZVq4+
5ukCCfCpEsK5REvlSXgPG2nvRzubMNzS8Sol854RJK8XYFnwc+4fRCqy75hI
gMnMqJrjO98xyC/LCqW3yD+9G3sbA0apyaA6OUOq67ih7A+c90e9rYHZ/8CC
hAuwiAueZTX2LOihbVXvkAKCl7zHCRNynVheWogt8t3QeU8Gce3brNAht2Sr
ZQr+E4nRY5pXuGXVP5tHtKaxCn63g+dAKo/gLmtn5o/M+y5SiTaBmozwBVZf
zFtNJbABnSRjvQEt3Uv3Eosw6uPg9wshb7eMQMAKieWvUyrcDnPYpm24hsYX
D98aAS8ps/pumKacYElVWn8gGxPSsftOsBcB0Cp9wK4RHPIXgF9AVft1AdgJ
y0XKn8/k6XZwTAVoalxL7APe1/O3spUz+X143hV+9UL7wp53JbXICF2MuxmE
kRUQDVT+jomeoMGtWJsSdM+/OzZABrmqkFA1NZLfw4tuoimikU/y/LBTYeWK
XzBG151vltBB6+pjOTJRvu5oBhf5p0/mZf9Z6UmjiLjWXvPs4LTbZ1kUyZ5m
fCYlIUGF1aAQNMxzHWBOcIalauHU7cxvUYmiALqLS9FkYc/awlnPfr+XLbdL
qMMaL6CX4R32H6P0mSsu8jm0YsylaMWGHHchOw15KXVkoxjTInNPLmGksBrf
bvaMU2QgBRy22xMpAkVt7kp/zReSCrxBVe9WZGaYphHfNby33v9JXC2FYg99
trwFjkSo+R46enRFDhuoVzK0g5e7gQVqbH8/vOo0zrcL6x92ghX+f71BXmDm
CyPYQgu9yNvfKHdhdPENt03QNK27o9t+OGpbOF8Dw0ggcbvhLmDZ6egsLy5V
yeD3u6dplX+E/XKqL06oBzD9v21N5/mor3resk0cazzPX0uhN6cWRX7rNeWt
Hks8hBCbiZ9D7uw/LUoux0zMwC2Cq1pFAGwnPe+kR1tc+BEyzz30ARwmZtdW
7tMEt5vk6rl4km32LfRF2dzsWUyu7NqnuHEDBpLJHK3JUFcFKEGutVhthSDp
uCTi4eo1TuHLJBsxh3cTVbsLQSINSWEQct/e62TYip1pUbZYKWoRbHh4JrBX
dpfbGkw2CuvipWWhTAdPUNfDabXx2qppWJdZ2qacExmqgjgevqdk0UcjNwOa
sg/pmW1R1F8f5MrTagnv22U0sDSaiCKi5ETwILlSejop+bWHIR3e3PifFntQ
Og0oe9pGhtV4NFAL+5j+CqlEcIJFb5oRmZev05agfoFajthT9TRxEBG/piwN
Zdgc597V7rkT4e3rB5yU+xbbHae6+EHvJqZXcZAKQ4SWO79RkcF5qn7YkL/N
O1Pq6CXchQeO5HpIGPbNQJiND9zzJX09EqftqT5ODYKRZlXvLi7zfXs22trq
d88na24h39y986bIGUBFYW9kpbpN3Z7CJYBI6TZMWc9rL6bgoncjaX3n8RmS
t1w4KnQ9chtTDCdcyv41c0zwSRF8LtIRt2ckWnfQ0+JkiN86XZpFvph0VyYx
IAoNlUGSv4pSW925d16zRDa/isGGwrEAuWsUxprJ4nOh/WJa6BLIYunfSYa+
V5lw0c76j16/CYMpusHz8MKlByZAyyGzMzeyQDt2297GO05hcAC1PjSgXzPJ
cd3Bxa3yob6nMM/p/KSL6bGHX2zLRebASR8sMhNdh16WLq9eJqR14fc6goI6
t+OFSICfu3TpqpQcrKjJhipQ8c5jSPVTnzc+xlcnt9uOEcRh9DnONKmdgQHn
rCPCJNdEwhAfv/CvAF7gdKp8aYe10+Oxoj2YVGtCRjOwQ8z4TDkVJ4Eht4Ug
T98QkziOu+YpAkrQMiT+TzZIHHKKLGdaLYTjehnhFPA8LQqr3Ynh2eM5M4pQ
oksP97NQhKCoSlBfOx0t3V0nq4S7nl9zjF6Owq8ExhGQHleNqN0pimEKK5c7
ZNjyFD2EV98NamNqOlRuOtKkk5bciBmaQ22hZT3SJ0ruk3K9Lc/mjCnRY3qI
kujTwyvAtrIfWOCu7i1EiUVPOoQQk5RsLe/3P1ZMwaUf4wYdxup1qCv0xs6e
SLtggPvjcRZkongH9hS2g5+6gdYic8o7gp6jU0J66zBL5pDa0eer/3th2ykI
E9TmTzwl5uqlg7YPtgV+yV2+ard2nOw4eTFw/+WBTB7RxvGg9b72aHW7Xfo4
Cp1DiPRlQCT7XwLJTzX9eVwMO0hkGWkbMQ4DDLdKfEi+TQ3Q+C6W+7o6xItK
fEaTR/kPPwYdwdFuDvlURoanuBVxYsOfZCS2VdQd4PJ+BXdZPrLicps/p9KR
Xc+H7qG23mr2KVip6i22TLPcm+rVwZ1I6NTKMwRJTQOLGdPfxYuMW4Vs7+Wn
xN7njwsTIVFsWHoFL5L90FRLUY6gnjjKH7yhFHuSrRJQ97UcCAW+npvxehmj
DMr9UqgaBs+IBY9Jdw0PRvUe4amgrtgEJPwX0xvypHgxtrfos12Aza6Vm2Zr
g5thlhNJC9zclj5S4HsC+qPLUQLseIVGSFwTTgjyxP5bU2YMmXXj6EaO6YyH
OpEkqkz+5hCs6uJBW9dKQmc8mDWV84fMjiFnyij3Kdd24rZi5DHJyHaOd2uQ
E5MGa9bPA1TCGzY3TP3aJyFWr3hhXWo1VWbrT8PR6HpCMFqyEtMi2dUPEvDP
VcxOy/4mbYlofts//j03U1tsicTwPujpnFzs31uZr2RFAVPLXqoMAZ4VPOsx
6w8t/T+YleyTLSTGM9YBKH7mCcWdRsXRbSkTLqJTpRukK1fgjt3aaLLqZZpK
pCRf3MKKwxMXueRccbaN2n6BqfFg5xOTnu3wCQ2DQXig//JFGL8YaAmS0I9m
6Trmvat1bpo8nmBvXB6Aq0of4wG3+gqXUXFXSDy6zKZ4uALPK2hjLrTertNX
MFPYSWLNyl1hIBLz5dsdM+m6Af4ZgKKCZ2SvHnlQZ30OFUEPwXVaWkdGKNLT
igVH2UwhoS4DMmojxM5BNrTJY5GEbYy3lJlt7hKtGeQlgIyK8aJO0ungSCHi
xzcyG/VAujW4xoRHYXDUdIG7ZBwb/J6TtYOAmGZS0wOAOFOrzuVkpxMJoJP8
TXKzFaLhdDjfNxjPpAaLx9deQUE6Us1qYKdmOYLk3KaYnjAOI6Qc8u6MVXwR
xM6D6R74kgQI4UkNtOdjfGCCMcBh9rc54XTBoUj48vw4BCGrm+qrAHx2X7vV
JbM72eLRpecoPr5nk3jFm2VzTE0CP5BX9P3E2MWOVawk9EfL4ExEJ9BO3eJN
jfQ2VnzXlQTZDSfxchcAiJOTsLLTbw09Ii6wVrhBb2O3Sl+U3o88IwkQu4fe
OohsZ6DfwXSAiAFY1Ee060/ACjOsJ8ibNp98QDsJh0CHutB3tzUsTsqxok2z
xw0L93gmHrb0ns/TWh1/abcDkO4AWdzcC/SHDizwxk/JQ378RmX0G6/C1vaT
QpjL53jzpNzGDwBdegcdqScNHFw1s3zAlUOuRqqTh/p7p7pKC+66SeudU5of
4VMgNXZaZNEamMRbpry/EE/ZwXQSYE1eRruIazFKnFiQ6ClanErC+5q1OIML
1/QfWEw1V1MtWkJVpTIU1JyP1TkqF8cWJexdF//q1tIbIY284OCVyUCJtWkS
hG8Si3oxEQ1fu73dbkFlTXRKr9hgvqnhyGHkZL0n+vQgpYfaDvYfGbPKn/dY
q8wjVqajk3U+aBiR5Ul1x2bdYMYXUSle4Seyr92hHmWW11NNOSeSMMRJrWN2
R0Z7jO3cNQCm9XvDC8AqwFhaVmPE2Hp7LMT0mopKQbGGqQKo3eBdnECMNNjL
eVf6erpMM2OXnkd9iVf+GI33zfuTYu0/XzKLzx0nlvEWi9xlOpEGo9S/LTJQ
CLhroP7nese0Sb5Qs2dkDO8nTSD8abBCp8wdh97Ls4bZU0ZzWpn3fSpzM5/A
iovRGdPxh7QcLnMk4OG4z0VMlXQfstHmLygm6ePzODnYAAeUowJvHKlcqWLY
ozB9+N23JP05Wr7oyFRm/G3AqpjItU4L9AkBHp3ae+6uzLwXzwchXfo+eyl3
znfKhuNHTq7bRyR69/igWzC8S7JCqFwB0UMBsKaTIQVTGeNIR9USdqCOg+BF
3GlxOtJBSYDBfQ5jkCSFBQFdmhjbFy+uYjKfcNJY75TN1wpMofObZgTXjnof
5H+shV5jQqG1IXeKyEu+HUZiqtLLbOc4VzrwU8Eo5vHdfz5QGeYqBoGSHVhQ
iByhHDMXKBq0JUx+7KJTMnBAbwZgfNBzs+NUdEvPfXLgLGQM7ghq67GwRPUG
DO1hgXakc4JCs80tSozedXIrts6QZDtkA6xxcPV0YbQQ4dYjKgb23bpVUAaq
y6k5R5H+b8PGTZRJUwQEUMqpxfkONdT6BY7mX5qYZsjdjH1nTXr2t72qPmfn
WqhbFLhil7VLzTlJFRKMQWjqDBLCATv6viFgnHvokAZEGufwQzGnbaBATv90
QSiTC9vzEaultq/9kpSrefRvjmOHsu5E2tcgOVp1ufwr3+4xdQNgYVIvf5v8
6b3epHp7ikIzyy4SuaLC1wS8bxDhCGYHCOwKa8GLBs/O+x5j/goL031t47H4
H5YXGtV3QYj4EqbHEmw3RMVxfm9qGY02JOtuZPkI3QSXmRUOEJrhNUcR3O9w
CbOG+s0IFySBjLcOXH86AX7LkabpAXFVezVoEZz2fEq4jbQLuIr5cZGhe7sn
ngYrt0xHlXTn0xjr7QBLrLk7MDwsU6DNPP9/qTogvpgstyhLFrUvtBHEzt4V
HEZQjWZBsl1CW2OX6XKa8y68EL7Ht6ZwvXc+FOgXpP53RHt/6czDOCiQ+Dx3
tT1+HYdFH39fWbq+2a3QHR08PkeIl43U2KRoI1oJB140stNZ8LjMoEfpjwPR
lcEm1y093lTQDQ3s+/1c7oAyDKLtmo6X/SvNaLV2QW1i7tM7Gbo0pqpQIDbX
v/7d8ivD7gFTql6FZYh18wDiVVx2oHbV9v+Iprlku2ACv0t6kVxDYsQg5nJQ
sbeBh2EONX3RisGIl1sD6BP96+VXOOol8kqCJwBE/K5vZGxuNG/SbZj4RAa9
XPARd5pq+GOO7rHEq0WcB8EMv9RGRv/sh1HZulzVAsVaYp9UJz6NofyoRJPg
vHgrywVzP0rdaQ070C8eWQ085ChVBpjyhq0uPeyMy89jABsvWpw41ZJoX2Aq
+k8vEv/OaTrZD5Ym1FjjmxL5jX46xlStuPamQwchNXLzcIGDLHTQA6PEnKKx
rkPx6xqbtohlvhMGnnnmXAwNZWqIBdAq48WExWRFthZa3dud82KXcXIWJt2M
oAKUcjiaZ7QBAYQUGYivK9g2o6BconBY7ioTNbVfDf5pfcZ1Xa54XRSUl986
r/2hSbKDKzZlfXEqq9RVHASeUl1pz3dFa2k5ccLKr/uUBebs+CKGQsFM2AOd
1zHfAQyBU2XqfZeOarQ7G10jGL5cqXSJjQQhM02HzsZbgu2xdSFX3/cIaUS/
0Cjx8ET/iuPW3S6i4PZDh0lTNPAOZaUwBbhMp/Jn0gOlvXxq0uMPAEeY87qM
C+j8DNXnrbgnLiTjG7baFsgMJPEgMR3NBCBpl5V35hTM4zTl5iXowwEsRIMS
uk1aKTgZa/I7o4dDCbEPeUxmd3s5UgGftH2N+RxfWjzfl5hze/4ZRM+y5k1H
itZFDP1LF7gY2/ehBaHtHw5oQgQcLpBzv43jqO6Iy427U1x5vOkU0bV5gxhm
zFpkhcNBeuEavd2gTHDkjg0raQvwkBJhr/eiG3eGEmmLSW21Ij6Oz9fqVmma
setn76UjMT/3SZagrJdaOvZ6lDmuKvE/95rBLeYoQ0s1DG+zI2qtAiVYihkN
jmbUUJfqqFapbGbDmaKyL1RU3kCThDUggpBdOD+SZVMecU5Nf5jAr00UXKJc
mFOSdFXHoNyt6lyZiQevGZb97hPGiqJYgxzRpcQRAWnXbiOxwuZ912ZDVXW9
2UlYNei9UcKYpA++bI+y2kkd8HkQyahkxspxM0jkcnFzsfbKDCuXdcBD3rw/
DNZEIIwryWssyi0KaTyG4D2lZXO9q0kKhw+htOC4nlF6QiPttsEkKiM5emDw
Kfy9jfYjj9NWRTkAKAvwlcfV4Q3Aqw1PN4cdwiOxeAjHD0XRJtuW8kCVTQZ0
/LpC5UmldDkf2aUFp1/J6lzDcHBsoY1XlCUB3joixj2Xcd1yShCH1juBmBf0
YqcjBjYWFKRyNBnAuW4bxtPb7X5ABMKcu05ahNhmq3YuoNEjnrrZhyIdEBJa
yDZFNeUBpbUzMRHYrlUZFhua2/bQViGRO4VEmHf8lVeeE4UOapFlbE9lu13f
uRaipnL8CPtAZBRkFj611ORhbHcIXyUySSCmO995VGJAPl4pYYX0JtPcda7n
pNNZDUM/Im5rvAjQX28aDxlzqnWDUobw7tXJj/g4XHCfntx5OrGH5VYQ4Dab
HQoyI5o+GXxrQzaOkTVgBaEEFDwUg5e1Onrul9+ckwfxE/iB/9OydgGaUdrs
0giagWUb6ZMVq62xp1iBKcJrxh7ubU/f6vxie+xWjLLSULFjYox5Mf7dwyzM
zNO/b3hHAaugcimYZyp2yOY+jwsTfClpHjDgKMUt5ZsNzVSUE87PvCdPftCX
UwfUF7x1B8Rvp994fNYqYV5wlw4PLpgJBKVPxkvgjU1/Eh8XA5QhcW9a0H79
YmF2l3kbEW/Ijn6ghfp6RNp6DlPLUvWBT/FgKo4yOFy7HaGDuRNSKl3IonQm
Tr+sNfUuO7vrku2+E/sy5yjAk/jdZ2wO+DEeWWY3UWWYcZuukbV96sV+f9bV
SDERCZa3pV+vMJRNl9Y2S0sT92J7Y9N31hpt0UKqP5HgjX9m2DDowJ9eM88q
JI6sp5gj75U6oH0ZX5qXEzSfpVF00BMltudpH3tg7FOgarKV4KRKuMez9iun
9vAbkSkReD+G05mvh7LBR8DT7UojAe31RgBrPF2E4o52JxG6WNrTrAzgEUwI
7eLp1GLXQ72iFzs7bd+UhIF7QDwZiq5MWib3yHeI5SQPcAUwQ2ZAEHpFUi+6
KE5bHoM52sHELATMrnNrxVRfvTRztrB14MW66pvo+nJpBOykFBGvNgLQivBr
TrR0cGD23u6p7+JGLdkGCQyfkkjW6TeDlqBLCHLjQtO+9YmndugzbQvBjch9
Xu30AaCcEz54dit1whK2oD8haAuJkJ1mnhDj/qDcqNRq1FAiJQXpV4OXhjH5
NHG4CAwXSWUwX9YIR+jhVmdqEzM3MJxO3zeveUXjkPi4XZYryI5mAEufTBcf
N+I3A/yQI1cqlWBwlZTZTocVDymAl6sXq3wVRK4Lqx/87+hU26moGxrsJf3b
X9Hngjg8/9QqvBDTq/T2ZlcUvfI83w2+2T1CZ8TXeosXvRS1wyCDAUr/QmOq
97V0qEkTPTgNFsN/TVP6u044e7aiUo67IRxGlHV4MNVCzO0s1j4xDnyy3pPv
I/aLvmC9kG/eCHEFXzIGvQ2sdy6ZZWHd9dr1/EFURhIjw+AQ4ym8x4aQDGN+
nTLI590GeKxDTSfJc8fAk5SB79WBeZqpjHHN8Vi3BzcxA+MK0tDvdc70o9WV
vS4lcLoKAlgx/BHhsguiL4nQfnyVfmJy9vm9hnT4qNHI+kbh9HZtsh8xzeGP
ZF1AAxjGSQmKaE71VYo8rvcvw9ic+/E4SO+CDeJJL9vGYfjoYVQku3y/Ng9q
H/KIoIjq4xbctwL5z3e6tnCU1+vqqlbeVYu3l4L6W+SWL55p2LwChCMXzMrL
9+WKR4ahEYJvuhhQzgK7QWZxa2Q9WjafFPn0vnkHpH41FSK8dTZKe0PiyEyc
V61gv6Cwna2hWVqSUWXaNyEZxEj9FaPcA6YHizthMm+NdvXQ6MaoNm1nHi96
XjCZE/mLTDJVJ6JATaKzZQZ0rljmZMVeQN+5SLh74ytOlNGCICGF4Y2QInwn
bC8t2Af1d45JVwUeClksAACZChrXhOc8tU1s95tHdHgWb+O8SAMpbl62zBpJ
4uSpehM7ipFzKIQ0odzPQI7MPdCHMmlDnYjPWXPN4hPtYUa2i8tef9ShxqHC
aLCSHpprXP3GQGTOFrWbo2kf3hbD0v46f/vi62RIyIf4VfmTs+7qGI+HC6wy
ZtNOWM90EMkQ1j489RjAObtpZ1BeHSem8JXjviFDZLbpORir9euHOe7noR+D
upSJh/HeE2YfbKW94zTv+3JNbq46qyfPkld/9yFIZAMIqomMECZs6oFlBlSB
QyRVji9wYYK0E01QPNxruELSGq4hEy7IMIVSa0oSt9SJH+duoi8jwFx/0w1j
JSYpRpDkCwfP//qwJUDYvEOcqRC6x2puplkVed/yz3KJYQKbX5k2JzZBUS+3
+Iwxus+1RjUYVTuygMX5YvZHs8qz0e6jdDMTcdkwaDe53GuFSo4Z4MTtoBsu
uwW7DFdpamsf1SqsKosOv1NjFGrROkQ4ZZwvgRcyRv7wS9qMvVNip18TTDWj
5NYSV4hSxpEf/ex8bV9HCNRB3C1ZjTcMEQMj9vz+VdupN3eoS+xhLc3h3TpD
83RtV/KlMAlBvAUtkrN9PcGlxAH7q54x0MqvKtffLlMrCi5KoM8By1COZyuc
RYrgwboCn3ht1RqsdE++19BcEinJ0kPXAGPY10NwwDGWP/7/BVaki+NQp674
g3evXIrG/HAYU/BA6ZBP8sh0qDYKUiMvMB7br0EoDZNV7vKm6DKZah6T+rRN
R8q+0Wt7EEBTN1F4Th6xFTZo6T7vk6egcjKL/H1ezG/DZOJc5BRViSuatqlG
URMr/8X2h/DwPEDdkoq1J3BjSYbbZnvXkOLstuVdUCHcffDthXRJk7nKmk0N
lspAG/19cNDmRQjaSEToGoXBHJ5ILBozfAPCAU+6Z3QnVWTaDI44HOeZ4U5l
0M3XKtf9D8tOTaf+LzSnHsl+m3qg2Exl6rQG3nC2FKTd5T4rSp7NFb6nZ4a6
D1CGVLNuAuTHJKWIlZkBYk1es0mDsHNcCsvzhEVPsqOIK3nSCZ/3pA29BIe7
SQQVtPY8WLDXSd5mgdEsCDUrTdepVoziM374e7VbGGePii7YR9EGCskkYzr7
vkHDKQdjgkTgL0mMrdQIQG+1veQzjHNBy3uimb3E0+y0SkzFj3kH/kvAT8JC
4NqWnTvVPGtF7vrx6vJ9fQa94iwze4z0jSTMZ5AtxFlrQPrsHjCJldOXw9WP
whOD0UHAEPV+b2Edu9uW1fQBNU4FY2bHplxaRZBaPyGxml1Re4hKlxRWrAP2
AVr/3smiDHQxZmDAg+vBmrvwtdxy0iry+pRhs5G8r17EaD6Ta9iGlpuVhPaA
Q6EjS2xbWb493lB8WNxL0n5vNJJOmjNZDbvoaAEmZFkIzsdxIrTK/Ra1g8Zp
eSVn29Ectyz5TUlOiCQpCYY++fM0AoLW6agAONLSaF2AHhtfxuFuJW8b6JwN
tjPKJtvF6a+4AoN8BU3Gw8Wvbi3yjFPW3Sg915r5oK/NNbcTInUsPIbMXX53
CkpAb9AV8vaLk0wYEEzDCFgvUORe+OqJNkSuHGVXrwSn+mhZM34q35KfKXDJ
J2gIayxAfNiUofSdx7Br5fV+YSiJagSOR4RtqkV4igsFAt97UjPQZKRtCC/7
0+pD/A9a+fhTus/uzwXYZ5uIVejMz13WqqKGUVBh8baNlJZ2J3QWtUN1H6p5
ZZ5ruNjFi8PCkbY1bNBCby7isrL9S2LQY5TK062GdoDKRORBYLMVYeqUc+Ai
AxzWmprNEGSJ6ldp0vDb5+KMRK1bu86bR5BWbs1xTwa1VA8V1uIhhBJD+Qc9
OtkJUDOntoWkX+BemvZ1PaXa1eub12tGOMKFuU+hc2UA02As4Et33ZXo26E9
0tgNzv8B9chId3iZqUskzD/LdEb2rE3jIrMIG+Q09TO9jUy12EGXh0+t+MD6
HJ/WSEEiysjoB+t3ous4MKL1h3xMhFderpMvUSBtgxe/XcQCfWRINdtxJFvJ
mOLsJMn3/ZTtSFWd5lz2RuJay4y38ybBn/GEBRLaJmKqaHURkMl8StSRe2t3
45tWeQyf5alWgH62uzcXRlpMmU97Kwu+8yHPNimNZk0AoSSOGxNZR2Yx6MLr
3jGj9zO9qH4kbCgeHBlNxrEN3HCzyJvaJWc/1xX3l/WEmdJfRwqOUg2kVPVs
yjvSFtrQqSYQ4DDjB0GWyf7rsEhsJYCgEq3F7zkqtxhq2Cre8njrs7uBH/Np
5TVviWI9psOi27r9Ki9Oy8aDkcIOUu0dZoVXtQppyNeTtNkDVLqs59lsQaYk
ULx7+cHw6fxtEnjGbnbXs1Tr7wZnGscqW6k3q6eRIV/BTDYDOafF/UGUtWCc
ItoQgkcaFSd5LOSZE2F4s7CY4DSQyM38IcYRbacmABA18UwY3DRvbTTscazR
lp6gm4Bvs5wI8vCuXykI6JvONkLo/iiOsuouE2OVKT1vXQJzbgWB3zWW7S4e
8Gmf+xvPkGS5oUNJF2Cb//uKFSpwG64ls9K9ml9cFBme2Hst/hZYeKzLwAMV
T2K+PPl4Fc9EUpRFZ0GPrdCb9c72X4WOF0iwDCjvOQdXw1xsFti9rAV1beNG
NYHc41Ew9I8ZOw90Ylt90B3GnjlcVaeItvzDLGz0oPGG44FFfAOKHfcuWooG
cblnBOAdUpC4atHxXEJ8BHcPkff3dI1/Qc7I2afofJpJyQ1T6aYv5bf3oOb7
7OjFqNYI9TjpwCwf32hR+ZDEM6BrWvJzo/4m5SquMAAONeRHODLC1yMARDx0
/WdLo+u+xyuWGCkzi7f9UHbBnxqoLeg/6409j9EM5G3ZmfcuiKS6VaSN44bJ
2144zNboz/K0WfmndRu0K0jCTeFHFtKmjbYW7sf0ReW5jipijZWvKWhdelVz
VVBwx/+hlg6GTDYFgGjmmkg1P1Kx697f2Eye8S1JTaUUiHcdWbWLJLGg9KJI
Yhll1mdEZG7uJRb/rvtQY6+OrTTSTR4CcpuMmKSUn2LDZpAbg6rCWYl2Z4c9
w8RVstpMRSVu2BCyNBX6mfxYw4ciDKuw1P2DrMFi5xTc4l9ITrTsKyyT0MZh
qoscEV3iEnfxezex69PYEa8PjKg1cxqZ65BHvfrUKFPMjnLFSQKvNqNLaBYK
AczIJ24+2XuN7w49tDRoOmGMojRGOeXqqZiXJRGhukikROnaFK7eeqLrzFdL
s6JwGT28fFlbEGVG9wpOUwv29FkbinLggjhKXNW5GBVaT0Ee4/wErskUjOnX
g40oWRbbq1Rg19xy5QdkGDYd2m/6Sm//VyX/51J8oKuwylyaXyyW8au6am4x
O1BQx5PXpkla7vxM16tTX9Rtem5KndpbTComLoxpRyEfoLtaWa5HuH92jkEl
xZPzhqrWj12hOmVr3YRiaaPowvQBw12t/HmXjSeD0m5Sv7VNRpApDsNbk1vr
hdzsLYeXLbhFtVK9PDRSYD4JpsnKAbhvBQaBk6WuL9UQwa/EmudTEm76KZLx
6R+OLmrEZDov2MoCLKQPkt36ChQ3+9EDfwe6Rt6EYrYf9K/Aaah1akrxCJ0o
vPDAa5LoztoikOn1oyDMj1SOB44wN4Zvdnlq+DCy+mLHC5qBFm30Pb803xgf
MuRgWNg9bLibJmTK9tW2r1VsP7xLX36zl6Ul2D8Bb23wGemLH2Lwn8hF8lIm
oc42Sw6knQ1/E0uU1G1xFa6f670mSW0v4IrVPNhlLLJdDJv98JYbWVnG4+rJ
OMA6vKKxvpOPGoQo/RG+Yvd0vekDM+nlc/QCDx+oOhDhzC3T6qO8B06v/btK
xCaHmfofJNVLGsWnvzvze2aROx0mkwNU5lm5sTZD3v600miZ6CdBNULlxya9
zoES+M+eLbYQ6xij2x8xhc5PQ4cMlcWCRhV11noYtmTv4JEC5EysCB9D03kk
UKR4Utc+VwM6d5sKFxrv6wdD2wVSCMjSG9sqXVMwQPsQYSne8Ljh+AE948sm
oU5+4MEGr1Z6KP/obuRbSxhPCLbn+vPUyrHkQsLlJltrApJW+0/8GCjUrI5l
PSRdd8awJBMvuFkCctjSo0JVI6npnVQJlY7+0PZVHiQizqtg85OHymnk91+h
9BNIFz0KdM6wsREx2c5u/vwXzYL+SnV5d1FBHnk14CiL4grj93EORPMCQjGC
z+vGC2BX6qy6samJeFjGURZFjapVBrMQHS6MmKNUy0mmDPUFX0TLwkPk249W
nhLrXmXgeEznfGtqbuOJHF/GIjeN3i4ZBaGiLTjXfrNPyeu4u/aUc8sWsx3i
hkPF8tcThR8Uu47Y7dwFE3hfQ+M7RpVHUg3BVYyq8y8t3XnVX66CZyuZl7cx
Ndn//YwRm05zmO1L0rRsZh9oHssR6skbk4FCXlMhk+bagwsKWd4n8LwwWSgL
O7acgXMBYphg+BSqIwvWEiY1v2Vjn9EVtUPHAev2DT4p5hHod5FQ6MYo6DSU
MFeklObC9FSR1czyHf1YyCvZkx0AVKVN7HbsGPmYs3coztHshMfxrrWSe75r
vZVJbGVYAd+ZpAyV+UazXS3lEbw8xcXuoSeXm4fAE1+o9wnHRiY/UOquoO6P
grwi3jYT/M78vxhh2nhM/OjVnJeUNeNWcBBGe3+uveAWIhMDGPJ5pWKDNKpf
yoKpVagWnhJ/FtU/T6RZvBtWsGjSpfC51rqYXODqNbim2pQnmXEPVfAocZ+i
kSE2C1PNfAVvAonXY6bKg5Njm6FJL+qO51+YghHV6nk2t7NEtkPalNJkuTaa
7TJ98jcSQFOs4DlfuX3YZ0Tro4xvNdRWnw9v6VLNkQLFL5uWtFmg3PiLzVVm
5Ypc02cGNHp8M3V86csRAdtXkJrdHBdvWI/Nmu8MT8epiHu3ofWiJX0VMNWa
LZKIl1JSWTnZTGZXKzhlu9Os3UfP6Lb1Zbw7Fo8cZvJBNtnZ9Y9MKTkZF9vs
t5umsnM1L8fa4VuEcGtzv6qgrru8HMXrXoXmJDzl0fzzHGZeG+3dP01mPbV9
LpATkGzSb8ZF1Y2kzalDMLJQMWQRjf4pjPT7c8HKdo53DQooxX3OqKeYlf+4
yfVU/xohm89S1fpmhOtepj50QSxElakL7Cx0ezMiFuOViEouZ3qznlKoF2r6
Ie3K6DkXksMp4tn0FBuiyBrilda8gjRd6JFA9J6++McZVRjlfcDFDs8XjSIg
l+g68aZAJgNd45APwmmUW0QXq4TUw5dTlplGgTggkyAKnolLsXbmx5MGT16L
JiCbiiupzJMU3tAh/Dyo4Em4ZJrz+Lw2uuuY2rJ3G5JlJQ7BLcDhkPQVvA92
QNkN3NqbYUHd9u5DZa7pVjc5TLLU9Jh/5n1WRMac4PIuz6gcWQMCZV4RMC+7
JDtunc+ZLrzQ8WVXaaczg+Z3LEcV71Jkk3QBqWcN4s/Dh9Emy5j9xQ6JnNnU
p/I+dJKjeY/eK5gXnbMpDXcqKrdiui3tFsZPKF5i4Nu54FlZGdbygYlwhOM+
GT9zDdMOoTwLIpcn8Z/4e9y4HZGYTBHqsIvzHjc45JS8JZCQ827JGeW4BwG1
5o8xMw7urx2Y3mMcDsALwmzk7lsHveTO2Gp9Cb4vIqA7ETTElES4UnqoQIio
EvBU9fTec15S6HsIRb2hL4YZxuPzfDJIWkE4sEqlmDjwbqJBU+2GAvsgh25y
0/wgrn3bULwnAPe4wnymHmYJXxC6Hs1Gr4nKr6mS1iI88Who8iM+Zb6nzFke
eQnT5xDt55SFuhZLABccLGrQ5eARSBAJB9VHM888uKkq4RWtV3Vo6LBMoFS2
NlAfI7muJWWFWAWY3qZkxxOfJL1ZyXEaEnSihMpBFSF543wsi86Z66+mm+vP
2Ko4xkAQ2D2EZ7A7hlNwO7Yag9Dh43ol7cgBvyBQ7yq4wa16WD0AhqsQaLQH
VWV+ysSFzXvWpe/Ff0tbljiIx2VfQy5XATaydgYVP2dsRqo34uUEyA1kAkyo
lP8jdt9Q5oQ83I1OUnmWYatIrkfcqzg9vLz1qcHTUvX4e6OqJmoeEsQBw9Uz
+e2uMh0L35nRIiyhCAAtKNSrgpZXDIAeiyv8j84p7zTdu0f9X+KVkBXZaElS
1cuwCGMr53tJ/uzRHfHTK3iNBBmknCG1njytscVtChFAq8DeRW96ZDj8uVFM
vm1J65nQpUm135QDoKyJt8eKZPUogVO1aVC/ylt2AfcsWr7sS2RPBai7M/mv
6Kh7osm6R79d0CkMYM3au2K3Nqw7CvaTyNhGb+180LFsnRxwr02J4Cj8oA72
B2OSx8kNTUAyGwqpAuvQw914xgagAGLyZNR7yaOuL/iUnipXWfSkrhyjP7UM
ZA49J7whoKIJ7hs3NTtWN09JIM9VZonHkFs1jfiMIROH4KepE6Z1zhjUhL1m
fr7PPLjDEt70Ll98ZpK7QJOZzEB6PWfhT8bcXyeEeYJ12oc21V6NfR88yN7d
bFXNxp2XB3+K9P+TzGCN1CRW6e4oup7IFes/sUnKoOLDkrYdnGBZF/98KhfO
dcut5TzplnM1ff6gYJEze5bpHfqGuXnBW7pemVVXWC504RQzlG6aI9Ue1QqH
C6nkFpHmhUIDgQgl9ulEYox5gH894t6Mg+9nt0g7V8IV5FZbY95orPaD0CZO
JeDjOviDL5yVZ4ENPyf7oVwI6Gc9NQxj0tqOK07wH3kfRKLOhf1UutxG76D0
oAowi7gVULd7lRDX9kt2jmclqt7cZljsaCA9BqsUYM6KvqzCngArQm44sf8F
4/EiXMJz17UI0rh5waF/njMp+iM/Qd7OlFuLhkgJvG7eNTlm6i0DnXyeqkbW
K7kD3sH9xpXtLVJI5kker5330+wv2qZF8MO+EubjVs/orJN1bsFZFz5Zvo6N
wBCtfCj2MauTtCt/zr6ht5513HQX3DiOurp9HwYCrB+x1rIpHbqH8mSw/0dF
ejGCxWF/ZciWRtf37N/c5RqD8MFITIu5k9JjFO6OzqHgDhwYpoCoyOUUKnRj
dahbaqg9NSSkHLVbGhXsb2SGJyZJSy+YQmrTjFuiprZt+sVZGNaHLGrbDUZT
OPzhlNgz84dc5YVwOJV2hTHWBRq5DljFSCGuHVTLeGGZxCwAlYEbUpX5c6eo
8O8AK3cCzQdtUsWYQe42LHHIGnDLvtx2GIoFmyYiKmZwMfHotBLiP7IJyprB
r3DOZMvt7rQ4NRUj4N2o6mZWmDGy085D63PLs/OGIQa5sVh8BICY1PtVNXDN
6N2Zpi0ZY1fXAAA4LqD2xVkQAyUJWqZoNoKpGCSTweCBe0IBtxv39FRyaSNy
ydAg/35Pj9lAMynMxqYeJVTRydCahDrNAxEzMd7Njzp0PB5sftMKq9ONQFB+
UwhpLiuo278iEY5/aV9AUkJ6jpneLO8O76l/T5QhzZ/eDLDKi4f5rKnoU5Go
tHkszfqQWMbdOLkfVeM6xSJlPDe7exvZW/32m8Reor8gJzQcUO2IUCWkc3gZ
DcMrUX9FrT7ureY4rR9tlSQXPFzLWAtL3J2NV9O9KY0OjJqO41woqqG6r3ms
vlDD3d05/Knog1qMIF0taNfR2BwQNil56BEwiMiBAWE4eFjqYqIp1SMpdkzI
PzuhnzdcPFwC1BWSRuTrsT9/yg9oM6wrE8MFRUqx8x+nG25/AqVy3i41tOfs
HO5Us5mwE9ItDvm0GsvyJRV+d9ZRxF3vH6uy7w31T/FIRLX0G/Bnezq9RFrk
+h2EOW6WXPCGkDac+P8wA/B8yyUj65uCFbqrr73XUuxBXdSndnzbVuPwKEuU
Fz5G2jV36pyvnvDCMXAWJH2eHJ39VK/eb5KT1DOdjNAdJHHNaRZBDF+dtiTR
xCbofrp/quanrvEOeRwhluG5OYziReM2PFl6G5GYbNLsPVqcXmRPoFOza5KQ
V6fAhA7GXtv8Q64sYBolRvOsqfm87p6fgUslhGoHn3mwISVsSIl7rxN22ALI
k6AjqsSh6b9S7unU2jZlLG2kiHdy7o2t+RbeZS8kjixCVCgO4QUO++XC6+Lj
ENAomvfp3ZOGQPHggxBHGu7qMytT1+wexRqyDOMXE763RcWR1VDFPjmuM6Pr
pI52+VIHKmnMMg3/z1Z6fAX7c8WtcGg/5ud9to2wVKRUjsZO/ZulWT4OQrbU
C91oV7M+y8b0jq5x+hPKMTF4HBH2IuLWju7VBLv49b9OEhrgfene+w6PVlnY
S2oyLEgkIl4AWsVJ38lXdbtiSINm21ImUfT2P94i+8xIJd2OeNaBKmbvyWBz
myeEMTpmn5ch5KT9ysYHeKswQ6nUWgw2T7a+itNrKvRV7U00pdblH9+FF5do
02p8ThQZojh8LyVjD561ZYlvCeujX2YlCzHZLuJGfZV1IDsfln15Rh8tleLf
/gvdhG44SuvNDui+g4+nPsieQWhbMpcfz5it0aXc79W/anaBpcQu8PIRYwi2
cWoGCnfl4ru9PR9NlcEQ81ztP+hbg+I96zV/cJX/64d3JFGpce5a/PC1d1TZ
8hs+yRxMOTixaSl3o1DsELrZRS8c1vfUyV+50TcHO20MFMKtb9eqEFOntWlO
GxBzEdVif1V2k0qI+es8z0DevvGd7aYosSCigBQn0v9lhbG/f3U3uOCGk+pl
XU6Oq8kKykT6YvZpc8AgzxsJkjl3PCIAZsCu4FNqXV8ao+XtWINAA79Gd/8p
ryHLlzvvh9AhuBMb7jDOv12Yk5YYV3xBpvilpyI+3Re3ySGI2GP4f4Jbnset
K6iySYx3DKLD2S6GLVv3LhlxxEq238kG/rHu1Cmc5K90z4SDH7JEGg8lajXa
OFA0eBMXr4M+zK2EPNsphQj4dCRujpoOr2l46osJAjFHcPUPNGnsY4d3fQjX
HD5J9Lrqir5PFPIyxab64kTUTeDnFlOsiARFhdTgtF7RpHF0TxBybO5NP+8S
HBJrtTEvI7cVzz6tweIt9GXDloIzLQkjXBe2faC+lYWMx6Yb4NE5mE0aY4Ph
XagBj4a29KZaJnYnYm/jUIzoFJbEPA5+0tmDi4Nprpr5PAs1FVKpKrHS2ZjN
SxEcu7I4WFZXj/my6QTOkl44i/v98q9s4xMAwAH6yxahYQ0D7d9PLng/5P5a
z9hQn985axsaylzqiWdzWHoxUKg2UQq/Jljk8vs2tfCO9q2JyoIcjK/eX7g3
m0BOfiPDzNMvnu667eOuqACIbm6ddy9PWLfj0qJlxZsuf+YULzYZhTePWsej
eX0djRDf+PKiDs1QFSubeTXUpIE8kwsPLLCEA5ToTmBccgPu4oaQkC42RftP
/bMDGUw0lGNwOoQU8kQSVEyMmWM81SBgORd2pogt3ZzqNfVSO+Pr1mwjxRug
nhM5m70D7nZcAri6xd1ffuIZOTewyh5gvyIfqFpJYsjGpxDo8LaXo1+li/a9
beUhPxxcNIL2O/DgHPo4RQMrYdwCQ5KyaBF+qG8G1c9M6kz4celNW698Y+iI
T5iMYQQJAQYJOX1EAs0qTATp0IuzNPCL4IcC8WFDyP4lE/eHjM3VGogeq08e
YbSfxWSdNDzSQI0tMvt775Xobh8j4Dc4qWH/hGnHHxbSGAujyCxyQMJkZzRj
c8UMmlLm1RrRZgH1BsKWIMr4mOjMXJ5x+iR5VtVJYPdTe9IMBqRkL+RFgWwX
ffTFjiV7mi07Ozr2pWXW+CZkFgshjNC+JJwH3kfOFFKK3sm/w4Vx3m/d04it
HINrSTuUZykt51xjPvY4ZO43Y8AcLu6caW711aDSj9icNcHdV29Nfbyv1iSi
qjykNct19Ew5i/fa8Ip+aJbZhXTz6iRK6aUVe8KEVUIpmLORQT6f58avBNlL
V7ozPy4rh0qptNg02NvgO8nFNCGY2fNgKsrIRXMBlXeudIHfgbThmu/Y0leT
gXI5OzF0rgbd0599SloBf6q8lG8h/UuLW2rYYuDBmHKIOsYzUyoCa/W56+45
dQLg0r+Yd4eioeq1HWt3VvA9NJAa6+U0dAGkWPWn5LPlS9veLx1FjJ16s2rv
/Sw6XlR61KqopgUzltio5p+fk3acyxYvdiuHGiBBJqE/wq4A51omgKyfADd4
F6nFbEcTzBJfptHJBI7CdaA2X6uKi3xQvu3DWHhSabV3Rqu7UxJde5v8cTzd
mbS8SqZSyMwog/pcSBYjg5gdRGaP8svF3iUKxssH8YRjl0Owt1JFUhlOg2OV
n7ngzztFFD5ABe8JHwij9Nom+hd1G9RljJjILr1D+lKMLYnV/97do3sXj4Ir
OqpWaO8YtjEPdeOyciFTq0uNTysrWv+rJNsDsNErmvEsI11cEymEd7hVa2N2
TfgaOxJCZMpxKEARYw7iDUDoKtvIG0usJGV+7jy7Fg+Q7ho9NTM0CCnlxf72
lFdl6EGIxnVfHtsin20mW/1PFlWzG1TKcpw2T4yD9jyJXAEtEg6p4gb+ZnXS
+XYsgHsLM3LQGRzdgpWm3lHs07uRnWKJY/QREZTyMRiWrGydWwwS2iVAAWzC
6Pkn4rxd6BTFE0NErTQ0bjtyY4vqkt0rSODWu2zKNCWPNukFhxfmFcCKaN9D
1TfTyTxT5XVgf0Q5FDSS7ijWTZhwVgiuKVto1Uib90EW4ofYYdKgd1W7W8bs
8hsLZnjlnTmhCQYp44uTjg8pEnyiea/Ss1gWMkVS4f7dfbEi6CGzcPLoQJ7w
0BGrq+kMjqhiONC39Xi174DdMPicCSNG1klF2gQQyrWa101o32QFeysawsT5
ya6cRXJTpPzVQ9fbxr4rNoc49XEXJpjX1G8aYF8iSfdp7qOJS6JHgFPrZ+sO
YjcKJONcRnvnyzNU0OGZmU2Vb8WLOLrcWYXvKURqkb9X/Kk/5HnGbDpNYVwl
3Hcq0AgPjkBRxLStHuqNvk+2uA6Xa8Wdu5EuD4r5tAnosibWKz1jnRXDt+s+
xvM/ePQ1I6i2hAQ2FCfI7uwQ/xper/3uxybzLF4FrhwwkWu3W7y1XobGX3Oh
musQDmSdvGoNAvhQSBKxzWlxreET98XOmqSSTKKtqKE18/Q5Zm1uCupvbHCH
wnUof0E4aHE/4hdEYWlFXEt7tF4EFfpX5Uy+xnFmHPPsmxP0noqSyhz3+M5y
sQ7Z2XZNaRid3yGepmzimpvLl4YEVeTP4k0hHEs4zMizJiO210yYc2Fw8uiL
UH9p9JEC8ykcEvS2xAMxhx9fxr9o5L5WSerta73WZgLmq2ylGXSIytw99fxj
/o69talhuq3W6E/Nyn3iWJ7CIYUb0TYxTsI60tEfdjcpn7Gq3jhhGvw8FWw+
CHLlXSFZyUH2yubBJD8QQexrOjYBvfu88Uihexp1jLOAqw35N9kWEm2kQu3s
UN4XtYtxNyMI+0n4lVSwGwbsTnXda+9BQ46AJCJtkxmru1mFqyk4bR8ojvUD
7b6nO1zYhI/pzjfCJ1ODzwPqyYrn+gv7UCFUv4rIthHcgkLqZs7QAXQAKwBh
iIk6YCfYpdUziGpg8bqjQBO1EyN3GZPeU9jIpzQTou/lgIDIBTMq1t9rVloF
nr6J0/rg80ifmIWpn4BCAjk8CtVvKuZiX4yulFB9UKkF9QgDcjiaT5c2f4ye
sRn+cacV+W/6RUFcanLzb9NqpC4hhutdhybeaGFS4Q21sG3bXp2bGZT5IrJF
Ti0gDnO8Ymmo934pCNyB28ViKGWJIYSphhjiCyI2aRrXcJeMQn+A0uOU5XEW
bQ54k+BECoreylbWMRFgIoXW12qEOepT7W1+tkkTdycX+GJSu785g2WJSoBp
Tfluv40D5OSYBDzf6/EO3l9YEsmNbjOPOP8HarIVNbHjpUZcpnh/o/8QQlDG
XD4Z0wuxWcD4kylIqjCJxP4xxJuAeeUHKdKCd3ho47EPYY60lzczuPN3WOM/
atTbHAYgHkWH0zrTkz86FaDoZMaRZSuhUurU/2CcXd0iUeXDpWBCmyQyxffh
3NayjHfPoyBPcYpoRyPtxVJ6iMvZAggH70/HbVXeStL5Wp+cFHnteMXTyf/K
Dd86LgeubGCj2v7uR8U34h23YQ2Eh8S35lkrROrr5FvY/tAK/MNWBsow7/YS
SjC0KHr3yrF/yznFOTpm/TIc++6H42CuIbewALvyyF+kJqXiLv/NshQdbw2F
Yug5aqEwNxXaCqxsPm9GWh7ea/n73Mb1JfSYqaBfnNURvsE8wrIpg/MinMMb
Z7OvgXQqWxti4ffh5Shq+G0rWiKEOxUoIDa8CW/cqh+xj2OVq/yMOSfEq8Q1
lZNvz6Yd4YIYH2SLemfrrBWi40CWhYhMKEgQnraOD3tpzxllLq2nJU14m0fc
vqucnla7xAgmNX+e5w+ykj+6ekS9P06ljqsoBrMEgsnY9eqS7UgwBt+tsUKa
luN6iQyickiMztG3ZqJQP30W6PCco7OzqY4NrsoRl2vnSbcOC5UGEqN5nZWi
DKACo0FThjeRqERMQUAAfA2TJdfzzkhI8ByRB2kKNgiPyH/jxYKhyiM1tC2p
2cjh8Moe7ulGh2vyTtXqsMe5rgAZuBnAXDpZvtAgIPto/4oz8D/fCSWBa5R7
EaOB/DCy2XNdn4vrJ4qxj2GzvyFOJb1zK5VbWkvO1m93FbKAOSAfYPWIvEQa
w/SGVRXxUBQ3qm9f6RttZdpvFVmixCMA0RLPAAq8/vaD29VbUnIk/ld9t0u5
BUHXWtMfRt3cyBHXZEqngXGxAItqhno2QQ0CaLRAwtRP7LXrGZ7B2oCsYOVd
szXRAnjeNzeRpA4DkKt0Sq1CmHRfEnQXyzsPWawsn6Kqv10ZC4wHdrAehsjU
sec7kaCdaBBJD1oV1co2DxLXlI/mAWjuRIM5SPrfxCHT7AWFv5ystF9rrV4N
F9RHYOynNKz5PSkTfExxyF3FRGarl2X4Qib1d6pkl63LMvAsMMlCs1GmYsAO
af/hPEA+sTIbG7brHRHaTLTz1M2QB7/CtWSebE+zMP+FCi2VLnuQNxj0olfM
E4+OMRsFkPTCPEuhjLkumTZtOiKYcIvsJ/cj9v8GPdXky2wNt3eUV2rJslGz
nJOgBpj7U3zOE0X3SJS0/G9I4qq///BI6UlpIZUrhn+soucUc9mB5cUf1KF7
Qje2hejuchlMlpI7TE/u/TeaIsuablN5/Y2BQgMbCBRnJlveoP/IFSl4AbOs
MV8rROMGXD0I4AzopICjv45wFGBoph4SEBvIQSFQHvRiOUnw1LYLFyd+fzVH
QBTfpu6SnLeYWdsIYNtI+ecJv8XaUro7giQrvGsf7CiqD7SMF6pDZ8sTkBBH
B//aXfzGCs9VqbWc1sea0vpp5DHN2rEeAh9R9AsOLLzUROz+0YSc3jkGjJch
aIRBT+Y799q+hAu9TlpDYgYmKJcRbIf2a/TpnKUHdxINeUbga5MTbDgWPstT
GCznFzS8mGtt9X4wLY/QQTGBGL0lepIFYARFDaARqYRsFyAvtyVr8NDuLZsy
6TNNE5eYKm16gAzVSOSDMuGlzW8K/QCSF1ZmvpflkiBvbcnig6NifXq0/KpC
z83NL5C5BVTeoSLisHrF2ZHIr9lPi8vPjORf1NyI68BtcItQ+ZVaFtRGS1hd
W/XsdikCZtLIquy+jkHpa60gZ2gEqFAV1m92zpO1M4jRJpnrAT2Kzq4OnFO2
Son5XJhDS5+Dw/2MXvsghX+3tu0SHugk7TmIal2mSOkyArRpSCFM03zLQWw2
GarDT1qr+MJiNS7FGk2IR6HonUaMT3KkRsTIIQDVQFPnRjQ1jl5SoM4HAzJc
RXFgiq+Le15rd94aO8Fgg7vahhLTLiyK09MNbOS2YX6Z4VJ0PhQeXx6bEM1l
QBvEsekzGh0RZZWJaAB5PW3e3GtBq1u83UuFPvvjLz/QAwRLLwJW5DuFUNWx
TdIxZbDHWPl3oJfvJG1iyawRjrrx8zeKyWtCYwo+sz3yyq/ZXNAOJY1FSFSW
cqjd6J1qTLXSAIEirLdcEv0lsRUiJp+xddDbzWgexk3MXsou8vMenDQDfgC2
RPx0K6/8naYpEV0IHo/TaqA834eVQmckNoAG2aUXO69xhnBW+lJKayUpjJZm
VakB2Uo3Zdob7rycutvTlpc3uMEajkYQ3lMjFhHmVoy5d3eK7h8AWKZztM+3
Ez8adziaernNQzZc6Btk3ymMFS3Op76SHOwfKL/9itd3rvwru58oGRK7gTsG
8IEvC8lSY4RPy6k0PfNNDTU0J0utL2+p+crPfknl0cLUd1f/9q0lNId/8Uur
Kz0kErtnT4b+zK7tk+PR5+OsTPHRiQ/TY7kPYyTHOB+7KsY0zlew/7ogKtsx
oaeEPNHu4i9R6zcb2in8HdBoBJsSEghSpcw8tnj9WLzY/HhmR3eLGoyXjrbr
+ou/po1SmqshLi8kBrNKaF3lF/srfVDnDdI3VC4JPreiTX83ww6f6EbjjsUC
GCN0bB49eSWSuKZU9PwWEhD5C/zB8/aL5kxJt4XdcInGbl7J+wV4Rhyt9JWT
qkzZem4rJDlVTjI3s9POyXmkS91ZDz+vEep8nlZGVzvo3plKChYEgiDeQRuY
XHRBa9nU/lu34zcBdyjdGW06gL4DR3vipgCSTlFCslavdHlyEZp/GnxUr6EP
utBN/SCoW8xCsN5MUPF74i+95NSefvoFW0etUial02SOCtKHzfoEhX0FUKuE
iOrS0TXGM+99tdlh9yGrB6J1Bwh79e06Cy0ohRXvxNNjnzPQ16Znc0uqx149
eompwYQXBzjCIsOVzHTDlgtWdafvBIEY3zzEysy5Brq1UppwzIeotz0SZdAg
kx2w7DoIFG5Qy9xND2byLIqWHFg9dSqWb2gpQUGIiURrxkSrtyEmRAtiagsB
P5RLk2IWSXHGR4lMIZSBcYYq5nkg2jzI5ryw0Y5g/p7XS+xzbpHfCtXuOdmD
am2CXh4QEaPnHaTMFmGxSfbbg1R7CBhi146WM+Svo2Y31Dx4TucxX3Bk8hEd
97HEVI+lQC681YPyj8cp9VtoD8JYowCv9KOski1YWUOO9GDDb5SyE3jFLjwU
QBoGT5yDy9DujoQX1LhErv0cJts6c8Pq4Wn9XIsl3EFGYgiS6qfvPlve7VB7
zVKoOijv8V/Q7g3r21kggvDXlza8zQzfbU0fGmXeozchvd3++aTTjsq8gAx9
qRXHJ401gGgZnrbOXsa7EePVXhpoVn0gYKrwD1+pcZRX4DCe2b3pl1KFdAM0
LJtoUeK/NXi6rigMGijjiA63FmI2oO8Rb6pRMRuIuh6CGKoXcnkFfrkkfaHe
jQ1jULqQGGLI3exr1S74A2r2DdYoTtAiQlFVmLz9sdKK6uZNmt5H2gsN+qKT
9W/w4NesxmM1+l++2RfbZLZel/qlw/DWGbdblpLMfznmLihDbQ3E27OblNzL
0MhgNUxeNpoSvuqrncE2pmzd9kt5LHxDKYeJ/FyMoyZdpad9/rOCWpek7zBR
AnJ/0s2lrjY4Yw2bOoRv7EG6wUywUbnAzIFcv6uDiTi6OZHgDrJBf3J8sDCT
M6iCchy3S85ln+r3ZWxEa3MiVZ550J8EhD7hTeGqoKAUBr/EZjxHJay0wXCB
7bbX+apuUhR15v8GmAV6uAOg34WT4elsj6rhtJx+985N2rFzMFKd1tPBBzXy
AqVkIlU/ozIYnu905FvU7b0cufm3Gkk7PCt/FXDZMEbaW9kxrHG1wvOXlxw9
fKYkHZhIOozqOn7oAIYTHX/07wSTyA4KCnkfbbEzNTYtmS6zFCKbJkaGEhIJ
oqPtVYh1YI5LfP2Xki71t1zkrmywIKF06aWXiiemQmwLYF7WK8s1D5QVhG2j
Gg50Jy4I6Y0rr0jXdVN+EvF4e3k+zqME7O6vJFVJ6aummVYxISvCBi2Q9EQy
YF1r49o2puoj0QWEsdvVPKLFIRbQM7A0Clr1UJvAPlFn+Pv7dHGyA2x1D5bT
6wUlYA1pYjVxR8ZuACk0gycY2pg59DrA4c2SUtLXhzgva1wqSwS3uKYEpddf
rZiZ/Uzh+oI0zgkOsQbuDVmM71bNVyJloSSb+aW6n6vpUMn5A4B+1IReoXso
NPuTKzTqcPKAVJnnITeIHIYiRbVBqkxwved/Pltdc8ocxHxQeN22TkMERawo
uLrySR2s21RNw3r2lEd0yTKg0kiLxv2QVAncondj7LVakO0Vlu6qpmeaQwQn
Mx7/DMIQ5WWKaTTYh31dc4lQcEo1DVmh/AJWOvN5wy/qlzIDvdatE7Zho07O
omTOwgbkBYBhvozoqYx/MYTQPWJ2Mr7jHDhFkOMaM+Hi5Ez/dtTwFk3BHj/u
5252ewF5TtaLr9oq0qXHKKpT1D3LsCj5BvCUtP6wiOWuf3R1dte6cpK5YHV6
p2J65+P5QE+0NZJ46fkQFEe98cJn6YCsDGF/jauUKICq/idRKKt8Ciy5cSqe
AK/9Tm/qzoVUJEQtim3nfuIehAxu2yDFFpKwsJUJ3w1ee8adW4oMC0hrZKwV
lHnmAg8Z9zABnFeEBuXNP08yF1gZH+x2pExbojexerte//HG9fiNBmklPSAc
T04MxXZsiaXeRE1zV4Iu4x8Vx+rfihItOgelzVVMDV/0PoT6IQ/xTUrHdi+l
TvYV5wJEhyXknGUM54hPMBjhfXRkC7Rf9yK/P87W3yMf+6PWMJSMg7N66JUF
LBjV06UP5r3HXMz3DX+uK90pV/mt7VttxAL73/c0hN8b/HEsgDxcR3ryBz7O
xQ7EVstWGmoxCe6Kp80XlscpLZAjoeslPb+1N0cvA9mlSoU2olR9dWuoUP7A
VNYp3taEBsN48fxKnHI5ysUg2wdQCdxBLW4Yya5kogDwEq6cY98db0vOQFLg
fky6R/ds3tlrKKiB2RRAosdugsBK2HrkPY+WKqZzA89H0ZfLqcBxEQC8s7BY
jzpa/3w3gYGajPtKyQmNbJ6PIXVRpHjFhrUvcu+mx/92rb7YpefnhfUAOo1+
hTj024D5Syt7TjXoVZ8nw3gln76ESnoDi3Z85/CD3ehG0S1VU7nzuFijONHk
EnN16kSAtOSAlwVxokUD1ZUyQLNMGCfsweS/ch44qcXDfztCJjoG9Bpcv+Un
DPzooqZOMYp8/pqQr3o7h6pz3KfXGfK2w5pi42B4WsQA3RTXTCuNFhC52Zye
T6dE512FUqcRA2bnAbaOcMYHCTjzlDo9HssG217QRUuOZHnkhjKL5zo0039F
k/YOm3tKOyiYdtUEQj9etrjgFsvkbFGv4fIKNqRWign8+FnB2qEKePCCEUen
KoDhFTC/gGEukN8Bzk7GMRpDeZUblGgNsnuImuOSWNM6IyCo0TLk2eBl/c8M
mFX3pk5utfvFfrR6YXkLzhIMxplldrGpUqnL2ZqBl/Kv56i8XS9uF2WSP2ve
2+3Ih3G4E2yy6W5qdtgRId3jMipiNAH9lTmkiAdZMpGHHIT9eg03ubzPBBbV
A1s8Y/NZ1QvBk9EmRt48NHxcsRonFNM19H7RF69AZfj2D6uJW2i8vFUi5+ec
l9DIUICfMF5dtgZpCxMQzNpsjj6nBy4UHJeFxfawf8kIT9i9/Vh9tBETtFqx
RYTP4gK2vp0CbCtvQmDO4JYYqc+I2C9dd9VWodKt9jMIfJ2B0cazB/U4p3kd
seYigUpjCVEGOS6BJMq9kVQEsGbOi3YH5oNS3la/Ek5bvqDauB7WkYbmqq4/
iVZIzDesqQp+w5ReOJpnxMEcLW4tY8BZCOpDLSPMSSz2a2PMlNBu6c0i6N1g
dEiVuy0A4Cu6Hii4Tu6fUk3Zt3zfNUDAlwIvWC9nuMH8WvZPJXXFlfx/tQBV
AuKYpBS0bgkW55S1JObj3fKBAhdr2KPwj3WTndyHAlBrBMFNRXckPqPbu9od
FISVAeztw34ZfqFiJ5wH/WRv4nw0zmEv/Hzh7zTqJZmAKXzhJKO4KUS+UhFo
0XtzdRtHQk7SFZskTRaciNl69gYivwida2lPD5ZqvKflpRpkfwweq2+myPKJ
0nkhUAtV1pZt9kvmM6kxiMBRflpPdye+0ZLo7lXJHVmUrAKOi7zxFUcWuuT0
r1tMaIQ5nCYULyd0ixtNHiS9a/o+EQy44bvIZTvWWIv5N5Tx14SKKFzZB/cA
pWY3/XhP8CBa8//uF/YiEbfd53s3/0Zq5e1TeLlxxCqFQogZkrSqJkb6yCIr
gPdNrmK/HxEjJErBaCIV3Ja7FpAXziFKAhoY3G2Wpvv0WfPWsCuD+PWFn/Bg
8QXhwPPjKLuZlDGS79EroTSZi69Lgeb0ipN3lLfoPcLjiak3BuU6+y65gW2B
npsKhfmOoJuV9fkUMxfGDWgpB2huJNoFQuQBeY+rwkVJUFDQspzLKAAdzrFc
md3JmjIv8mBUjBs8AAblKi4/a1+8Rhf+8ERYjwTsI+YG6OfK0sQbhy5vp5yz
s01TSMM6kvY0DtxzLoJGZA9hOqbSx3rQhhaNgfD6EO4v6lVb++02WMVj8pRa
uzDohHd8YwBfJDHaMAwyJE/wloiCEXjBiZy+iSVsx6l2Y9SZsrIbOb/yeypx
Khwe5gD4qpGMP/OJSgVjgcj/A9u/UtoYOU8nsCfVmVmPlSbdtfmD0WtBzS9Y
dRVTyfIVjAl5BOgZzBOxzNseEuOKmD6l7cuYyct3WVg+zvHuAYVABzjYNcb/
OqsozWFmW4e61mDChKF7MoADjTDt5P8Es56+CEJ0miPWqYEYCLCxT1sZEMPV
g4wdcAcVEX4As5mrVijt4JJWU6+7d3Ia5RluK+Z6pouHcuzkg5q6XcIeAkN2
JeGotFqjm88/yh0G7fqgW5IWXXlwRUHjnXbAjT6vQTtxIFP47KIpxKvYUXyF
2t9LRjcEkBk4TryRJ6SntHVe1E3F0ycgolIjqOHAB5xSSmQtJI2HtwPWb2fu
2WoJp1bZP9usAYcjzsI0oxUPLKbe9/+mH16TPkkxOvEniqHzFHC0iPRW/DK5
ATcyerbn3YqqNECwQNqrWOGFbJFtXBO4Ny6TcWqFme7DinT8CL6D7mXfjEJX
fL2BeLCmY25YzRnZiyO3YMcWO63y7Y5zT3DMGvcaWGeHkov1Dn8hbpUV2MpQ
QF46uKFHX142Mw13RYro+cJG4wf34TwgOWfKQFJM6ZJzLjC+PkXBhkAv2aRz
2yeqVb3aUdeWZ09vKz3eb6z1JLTrLGmDJ39bLX5B2WsDKLLwUNwW2CLP1o3x
HSgqyR4x0naUHseMn/YrFmudr5b6wJr3Gaq5sGWziNkZWl7AZ6jfu5qL32Ia
ig/J8HyuMvpY42a6Z6iUm5I0yEi3LMAaMVQd5SdMBA47mUoBx+OKyaRwfhmm
MGU1OvgCU/bRUjK++eE3tseKLb8MAMFDRJTfLtHwO0SW5b0WHc4XLWt0jFVJ
6q4n91SCkEIAl9198sPg7D2hhWTZ/3+it0T76kOd96ixUko2c0Nk//bYROcH
f3owEBR76XZ9CLijqJf3/kjkKkKMT3kDaBqhTexoZ4HaUsnvp8SZbpGz4XW5
1TapgBBSp3TdH5ewj9zrr3JxhVk15nHdYS6DDPxi/oGs/xOreUf/mQggarHP
a3XhK2poGiwpmDaD8alj0Lkf59bau5oG9lC5G3qTRz32dbMXusqEw3WIFu38
JzvCKU2CPraD5KIun8JuKJFQTahXZgCn0nX9BK0u0XTJlxaKYJHCU6Dkm9Lp
iB/ibb92MdQfMhYAcObtjTGlsxmJuiUy4Z26Z8rRmHkX8RLj8zUJwmta9MX4
t4z0ju3FdpbwJI5fyA4ix9YbCL6yadsIMoFaGEcdD/Bj2+thtSCNDyI0jNqG
HpblRQYwSbbX/jBOSryHs0Rk0geglZFB5xEnrCYbz5LpKeFF5kvzke298Uxy
RbjeCWAuAEPB3wwXWoVPY9TlcirH5TRcejWjuE/XBWP/ZR+rmZxp/zKKaSgm
SPIIppuVIhW/l9ORsyO+aWe677P8KbEPdsOifeU/wkHi/ESg8mPGHfI1Intr
crWefS9HcesaEJFWRR/9ZMF4pm+eS1UhQPB+FsYDlyWbrspLWXPJA1HqPwTS
wjms8n6faFRzUUlA+Zs3Fq1rZq0rMp+zVd0fajvyVFQDgGuKHwP/JF2IOd1X
zNPFgk7q9t/D81AB7yU0OHCmyRd2k74R4R0Uvh8Fvsl/tOZtBy1d4HSInZ8M
Z79QZpLX6OUTfzeEYxru1UzFnYBW7tMqNxWMb9ohLKby6MX7j/SlkyI1yLwL
bTwppdP7E6qxCXcWs3HC5qk1NtimcC9CLzto1I/4TQQV96VxyjTZwQlu2WuC
vmmcIsEDlbSzOB/SNe+X+xZcJzkEtS/cjP8G58wkiFvi4FOFnD9dfLy17CvT
12Tve52PAv02382sZBvzwRW3ZmD91R3EQIiagaeYN8nfr5tKTvgv7xvxVmGu
ABuXZQIbbp3krXXqYRQ7Ms2/NLsjsgipOjz5ZL6kFTV4wFm33RTUFAF7j93z
nLesBnPwNQvM39hsFpXrDKt3s0TMGUtR0fgrsnCwhbfJ6fATES45uc+c0fJE
AGt1npIA0ZTU6SY3iOEQCn46XXi6W20qvV+DfdahfjlnwhP/p1Wz+mYMNlRp
+JeMCoAWrPIfcYJCxbH8UvPM7Gz6qFTYrpyaRxA+3bIebNUwgS1egZpvY1HQ
0/bHNLvP2e4P56reBJ/kHuSx4D6nJOcwa1HNPOViKPDwJ5+OVFDMPPY81U8k
nwuFOQvKwwm6crGDh778cmWZIkg9Hi+0c7ES4NV6EcGFtrQyMptUmEAmiO2v
LNt/e3n3Bhh6hMUA7MSLxbISW0UQd0fYokniXPap+IAUbUx8crDjzVGN5hlZ
jCWCUZkBzgc3hUyJBem4plRk0bEWap0jsWzXYIMWWBQCCPWwmtLq8dMotVeB
I106/07WX6a0KH4NwI6eZZbjXXESeNWvgWvU/3FIXH9EFzgI5jBwHBlyds4D
cviQYudBJ0TvbdXYzP8gJ7bZ3Ym/pcvRdvTL7cfkTcdK0yDaCovjLwIG0vt3
CQnUjOW5F5HhKcmk+PQPHqPS1POy/l6Qp/7wJvWHsO1Kt6cYnJEpes27uRYi
3wPv8wFXnWmbjSV8k61o4B3f8j2/uGkwTTwwWC0wWUnND8NuMfvo1t1keDuZ
n0r7k9EENgJ9rlH0ud+/iLijsuE/J/6IlGhMjGTUTdrqTCGozPVG7Q5GKJ7n
p4fzIV+J/rE1gO9tvjR71wSfVlAvuLVGi87udIz7lL6V6il77O4zY3ti4V0d
baqVCMU00ppALTS8Lod0cm+P9SJ8WBjpZIurYzEICUmrwauqRHKDHFBC8IRZ
sjQ6D3bw5HqsEdPoEcfX5XQ5XQ4XRIstKKiBRabakj6OvLvXb279IuuY+PHz
QGbE33AJ+VEGP8d3DHB2WENbWWLJxOrBlm1Q23UJ/NbtpSNV4ENovQ/FzCcz
ooWCneaQP0NoX7/ncpGdGO+mXaX2Ytwu/q2pQzz6/n7pagQESSbLPf/SsEJD
PoIOAk51bIZT6oIpnE0r69Zd0v3mIu10ydeDG5XpaGt4Bup34WYlXzoClNWS
jmkSHv6GQPZCXDmVAhM/JnFE5o+IK8H8zwpwTacIR+PajzVfLmDHljdhC2is
K4EVnivwalkrpYqe33puSdM6fnkEEfbtsLzSkWf4cN6bd3CSZ7C4LM6fov+5
tlDHeqQHU8hkXzkBQrjmEaZx2i6Kt9tZlvdAwhsjMq42MjaKRQcKDSjoolS1
OIk/huCmOo154v6CD4t3VHygtIaSsmLPpo/HhqywfO2CcvSRmjh8EFBXUfcz
VUGsleo9Oc+NCPo4yP/8LBxTAlVbNkvGs3nKXGxj5z7NhLsuBOyUZfINXG5I
vHArSOynIicHvJyBJXp8G2zOv75WS4lbmqlgUkcmfsLN2z780pWuhXJ44Ayk
iu3uzbuHQiVospShw56iX+BfmjYd47n82AY/w9YtvzK+it8v21La3AQcnUZv
FxTgPR8Nq3nmwQqChuAxnponlIz6qOJTSaCywY40LndKpOdJK15MP1bmFA7S
JuOb5IoJ/yXz8KcoFTQQFjOXk8bOdIbhXLPaMU77cx5fCzm1Mi/xuBWA+zwK
Z3y7cxOZVju0xvsuCwNMsDUPZs/S+zzAo2BH1Do90DfxttPJOAmVqjIOsczX
Txe5fSoQMfgMvO47ymVCl3c+i/500CPCMrwIglb6m3FAVIzlMypVjcDGM/3s
2nBLo8wLLWP5Ac5FE5v2Obk22VjUGaT3tLGDcDHf6XEJHFgj5WSbajg/VQqQ
Rv/wPRopFVpmtpTplgLrt7x25cfk8gtezkZ9ec/CSaoiaKXORlvOeGC+mBa1
DVYq1uVcb5ApaptYfP8J84V5Nw9BABwDh0wCpZOFhLQsp+tkoJbS7EoqJe9N
iGOBDeOSmnY6+GAU0CZV8CHrFH/akOcn1SL3g8ABMeVK9FCgqA/8yv6+Fmb3
fQcqfRSnPEpeqhr+TWRjGbRfM0AcGjyYXg4bUo+Fh3dC/th8eBYMEXuxaCW9
+ptjkwk9PO0jatKf+KQRLpH2zJ2Y53x+8TYmC89Bkw+P0i+BsEpzDlto9tM5
1CbzNvuitN3OvIakHBWKNxpUlsiNYYhDGkcvU9gTIDX+GfVZYz7tAv/vwfVB
96xUCQhtiv6CnL8lrc3KJHxPwAnVEeotTfhBgUOTMFk8WZlWarpyifClzkKa
19MRC5wlpPuW5OxZOQML24bpGUA4W/A+1XqW+kJz7P8gcQBI/AyXB/pVa3uV
stzTpUYtZprj6bqhIugBG+yP7LsmgpZRBhm1j4tqWRbWUMaYBZc9O/vj16Kt
NrlXmQI6VgaYbb0g2OVhDiZq6xZhyRiVQAf5u16THY943RNfgiDehVoQrbpg
lTit6r6KI2Yowx9Ephyewz4FXKOXdbUU5AOaVvJ+fRZh/zx6izAJhRjLREYB
7yFDC2LB3NMQRa8J00NbcWN1daadByFROH8ynMqBI1PmAw5SZaVLh0aauoKO
qOp/L1PS2xUL+XJaMoTm6XYCsF4eymE/p8k/benfQxOYRpzVXWmEQbO2kyZn
wDKCR4Tbrnb1RPvL9RwT61ptUcJGzkZRjsulsgC9VccrkSKPmwAUsv0ERcbo
ivUHRHfHxlCVvZ5R/QG+U7GjRkJX6cEaL4oNzGuj5xlSFJYEqtAAXB4w3YEe
viVnQBgDb5Iv5s5YSshZYpdDUB6XJHFp4XoYsoSuIpRmA4UZoJXvuCE29kC3
z3xB52+T+b1CzQLqBXkMw3fX79CtSCy4KBjhA5gXbiEEKjxC7/4PjwCS7eiZ
ZoZ9strNMlP0F5E8GfLlCflbA5ChosuM/6mcT4esGinXZnmq40WxQ50YqosZ
WQjqCuL5ACGY5+v43l70rn2DSOQWQT4vF8rmfv/+mK5QLYivawf/ox2R+7TZ
e2dxwndexJLmelj2XVJDqyaVhz9ho1WTd4cdj9hpDri7pRaDCq1+29SOraJ2
zerbX7nfMkRtEuDmSp8lVdP4IBBRhdyAzFWs8bKSNOhu4AoAhAZd+/E85Bs+
fZMnbAAUMB5P3lRrZGvccpMQou7wW1sxtAbQVGhE8nK6xnKmMB/XdMbHyNFc
WcR4wHBlaqlmIckHUDW7R27cxLA3uh6eaLj0CKnpJ+B5YbrICAlQHw2RZKfq
KQAZSYlPLiZzy/eDDOn3MfOwdtsTl02kbm4rcn0RpDTWpwIOr0OmjWdmaz0T
ZU+H8ZTBaOknl8ZkBWc9qWaAgsBQDiZhQor6CRZQtoTsJMx/Do997p4K1Pd1
XZH25Tlc6BYpxb//x3pw+pa+SaLNMCK9l2TTTSXHAzeyEPyi8ipurJVcdPKJ
WTp/yuKJnjtexwFxfGcN0XgschkfUB86hNSqh0mCfzAAf78tYOSb2q+IO28Y
kvmri/T8GKeQBU3vTcw6tfhvUpGe7PMvhJf57GoKHjjqF9P8c1mOnp3SNpmr
oVGmM51lcRpxaeNqD1NCT1QpQmgALJCBrRLm/b09BulO0Z0mHezTS1cLPzLK
2gTeLXN+GvHci3w6G5VaxgCmt3spEkgZqHYQ9oFTKXXpatNvSnkVIFUa7QQt
J1IPYIeC4qyaOY11fJcp2Pt16W8utqImZuw4NagqwynHM5t5+2+rMrpXNZpc
LbPO2Oln2v6KgsqWfjJu85otYSHRx0tkXBBV//h+kOvAiOV7pSOjWSaeh1dp
b1dRFMG3Cv4Fe2qTLQNIguZMy4Hcuci6xNNke1+4zYjnmJvkP/dUtwXjf3Am
zJymlEZkc5+A9Xik+SJTDaswov+xaImrHoev5jpsm+i9ZkN+WdHODJxCA54R
/kvI4k5H1Tb05MCxR1IPMBjeEgo5Z5Pld6HmtRrma+DSvNVI0vawDqhkz2pb
JAsYvI64wnKmFU0ju69LgPblmlVVmeO+/QDaRzmoNvoIwTi6ruBKaLn+Tojw
ewbV7mo6qIFDlqmmhGFfSkt72VDtWEa5ki4DoIEebT7y+1kJrzJmJ+5AjrZ7
h4FnM418772KwoJyps4HYQIx8T/NuSYeEu2wNWf32OV2JwkuSCf9TXJYJrTX
5Vc+VehixRa4bPtdqAqneh8mSL6K2xwLS+rsFM9YHLeEu3qbftEGI8owIuan
GN47YIeIrfrpcZnRrnzYhLUh6cqopAH8uyHTQ46il+XpFT7kjOnfbrs6kcz/
k4liCnAHWnfVuBd7vIESzh1vZ6s2WoSa2CmkwNt7AVmU9k7HU/WbqpuudnUq
a4e1ZnCodq3Xfq9QksPr5ReQ1BCkZvMFVhYrDlgNiKROVImSZBevMDBo3BGR
pvu0wqs3UWb7GUOTciODLiwge9feZ0zFQStyjQJnEpBaHy8sZaBO2d6U0hc/
aZHAvcBSUHI0ausWjOb86mg9Z96pzT3eHQ358gCax2BzhjTQp9OKqtLK2ezG
epw4aY75ijjyWu2cleqrNaA7qi8WpRDy3k+zkCcjZ2op0lIMQuPfEnX1XK+i
PbcDivLDPxzsXKxuVXgm2QQjYcrI0DZEZwBbGSPdi1T1LWCJE+Sr6jaAW2Xy
FNmDA2Lnxl6X+KlGj/cqcr1dZZv7ehECfDRhBrc0qykWH5vPv8SIegTnUkwW
120dCmkpMRutuAkbEPUqW6wu/iCTyBFN4blwYbOKxP1tmDcECcwZh5gltok2
h4wbOkUlAQjS1n7ZYzGLg4LHCcdycng01gVOT5F969sYUBtMbysTLk/BfZmT
yFe0VSOI9k7KPBev8MD4iV8N5z2sN23ceJZPOv3qFSQKvjdBQ7+0T0iCaYEv
JPXej8AyE1RO8r9Wz/K4XPOzLpltcqPMHZ3BGV5UUuMPwc3m4FXKxu+YB3nA
oHzDZqLfCwJSQ8BZugDOTZRY63UylMl04wqR7rMwAbHMR68gso2h3bYsdWhv
bk1IVIMPd14AKlOlM3Ep1hY5ydQF2k2KWzyLdshtto95AQm9rSHgxtJrGWH3
HA6DIkC/mgTctyTyKiKbpwSF9wxXXz0Gm0d0NrFIXCTPVmooN5+kCYgB1jGZ
l1DBhMACLkhSiW3EMZHm6q1qGTrxhok91X8JElkDtDGUu0DwcfxCwujfX3SG
d1LLIL3WmvU0oLusu8Z0OGb7tnqMW6fjKhjC0U4IQ7GtUb6ZFdW6wdkRKod+
Oir9Hv9BAHR3PQ1gXuNY/Urx4Bpd5JFbu7rmues0KGCtjA/9a8JsEVm1GwHO
dKfzcbzoy3g2FkJpKzrbIKzSDBjMKbxO10rLqfhbpEi8WLHzYvwIUAeni79T
839dHdqGL/YPlniQKZxv3uTI/t2lqFIKEJ7/ESueQC7hYk6kVqRTY9LZfVG5
8T9IS6AQouJ25uHToUATBm6fRY6uIZLm0WCE7LXYbI9hcbPc8ORxSX8ONLWA
z+OZuwJyT2NnNUUAEaZiuQ7GvJg4oNbtwhKAGlerUHOpmO2wXX19Q8x+aJu6
h7m55ge6Ntwz3It/krkuukyb5DnstOWXSMWjHeoh1qcFWK1/rbY5Al+Gd7Xd
S6ZEIxOx1VGU91Kp25yXDgKh6AjOqCd6zIBhBECMyS0DpmX458aCK+LwYTul
UXV2jBXmdHvIYuCWkpRd6/Ps/7suWFI/FL9zC5XwttNpFyckQGg38YqtdDO8
Y8cYIUDMD/mwURPX55FeeYrU6h3eOAVobShDTlK6u7mdhUIlpZZO90XFnYHn
+sbk99KCPl2t9l5ijCsnx4whdlCJTSPZ0L8s4VHPchQpM/qxwwih0QAnSVke
MELBxmWNODZCRrqMNLtP4qPxS0g9ehQK1wCxAElQ4XDypDX5hcGOor1ZMJ6t
8Byvwp8JpPRc9vj4Ut2rcjq4AbOLHx7XUJI/hQlf8nd4D++c91IEI1+z7odq
hT05YFCQeBpsvO4mFu8lvaIx19i5nZY57InXLsUJyiX/GG65euURLm7bpv8R
7FEpKYp7Hik9gKo6r+C361EOu+Q/fkKMvrOpJTG024qqz7cVr8M/rZhIg+OD
nmekELc7F7xx47lJkxWG63u8PGJQfanc6Din94a1XYsZkjbIcHkOcHO6WaQ6
czn5CoMiBI6vcz3Au+qVNq1RdrNaH5jccGDaJTsOPP8FSUUM2f4pLsfr2dhe
AwyYIVRdpaViuFQ+IyLxqhxZ1pbQcG8B0DrE95QKrmeN3BxkYT1QH9mWqNx9
cIU/623pYyC+JDOFd/nTcYtUEnY1lYBN+PTT1C242WBRUDpOYNLQT0YRENIc
J3ocftpj74Hrcq4dH9foMXXUI28RRzDMzXd6O+2F9rOnut785dRdDuZbe2c6
+T3LnG0h1dRJ+vvUZImMo+vcuDA8574gEn1nwbmbcr6I/gtZMhluIV8udVqb
L0fkaMbJRX2MIt2IJJmX2o1VEX4gvX0D89UyCJ6PG5LjGAcQs8NxlJUAO66w
VAEnL+C9ZN/kvqMAGzikqtYFykVDdMNgdNYHNCGM2B5q4MumJDyaD3hwWBrQ
eLpD2gDPJWBNdUkmBNETWtWikN9jPFoU112xlNEY75gBftGvEBdJ2wT0lGTW
WnbwI035mv7WxZzNQwdQFkPb73aXJZ7B19Mr/LO4nuIccbi2e2YLsU6jo0LW
WBfEfbH9i4/fpGhDeeBygQjseKgObZ0QapR5y3YzP805dwCge04UiVN9YR0C
9s/FhtierQrKmzfoWFJMgh+j0T60fjPsvCFHDMZwQUkt7qXM5/wy/SC4iMio
QTQ1ki5C0FNwq6C0zQrjp1hHYuq19D2OUVcBN9eDNxKqiKJdGeTbGDwPnA7K
LhaYB2JVV1qn1bHhEnZHJm03KVxMl8+OVD98spCXq/qDygg0f7OcHCVLBONE
bMToMXThl+bJNHIp0JPNi1IctmIRUdrGa0bnkOnbGlxptPE7figMIlVObR6q
Lg2UNnMv7JKGPZPzuYWti8sreHVsqUek57V7Z9QTijTFgRKhbdPOLMl2NfYa
wymudMNhRj4bMxooHvkR7k+F3oPvE5Jm2qtQ+d5zzBeXThRx+cDB1glE7GS+
zpZQ3Y3joI/53gegEO/rBPPsMBSHmtc3pwvgAYU6q7Qi/cKHwGnLdmBxNRpc
dQ8cdofA9PPJMmNiSkwLM3mW2SC//VLFYX8SkJpsF4e5f/REAV5c9cKmv6ok
uBJRXmLCHVupQSyquXsRgniqEwCNXtH4CPEIBJS6rBeX8diy/1pbalMeXTm1
KCwtWVSeGiNRnPkRjYOSDOJwG9AkV4CuHs+fnvJyY5wT1eDW7d3Zd4z7azKT
3Q0lmOjSZiH2XYLMxoSbdB+D8Rnb2xAfnUzL4msVzlDWK+fd4j6v4Snf+MK3
SDtCh8PGtLxddtW3zGbGFYxqfXkZBsT1ci+lLCVgxMw9kUHz/axys6Dmnsfi
t2DU6mBeL/563VZPpCc2DlZgp8f8ht0ihFxUgO5snCH0euNQFo0USN6ZPJr3
pt4q+RWSg0Antfg8GgWyrlavLXwnHpOZQ0qij/r6H8Otft1Bc7VIJeX1wkLa
v+gLtV9d7f9KOUxnU3ECXCYWxs5jrtRtSsGIl1LN1X+vHG2NciQ/z68yTksA
vmiV4k/o70sspCJ+d2iwduV2D4xN4KZb67xJXbm8X9tAflUrcjzv0yqyL7vw
UwCEDRjN7TQsyJYY8GFz0bNsPZ7y242qMMJ4zLM6FHZQuTZJgAsog+6JRviR
hD2dL6cINp3G0ONvVrL4GbWMYnXurteAUB/RXhlJDCrRvAIzOznZDj65VJf0
GQW/tody1EgUQJvmezk2musKV//umKRom/jZ/o4INzVUMrA+ZUpGriX39sOP
iXA8rDff2+oNN9l3AJlIWeG2vcQdPlJhf9Gu7uLriHSwEoCX/x1Zw0C6XgYr
6XwUd2jcCRiXjWmurPkWGamZ0aErudPpiIpUe/JA+kBMe1Uak7vAdRLq+89A
U2e7lspIis88uicwqm92UC8acHhR5KrvSF60bHKdDq7eMgtehNz8fYR+E1nH
ymLtBRD9ZCSy0AnB6Z/9Nx5Ap1n9nyuFSgw3qjslmrGZa9DeSPhUsFM6F7Pf
PExSDmYpkilQ+xIGOe4he0AtMn1vOSkE/GuRbP2x42HJQkTYM6xtWGSMceEW
DNnl5BJJh6B2/WRkp7nbfv5pPDliSTYX6AN8PL/GTvNUkSFtpEvJ1d77ylzj
uLCUkdCJbv+KDKLCqI3VAsCxfzoVoPi7KBkegA3B4I+scRK/YO5OWdPklu5F
2duB8/MaVbiT3kbAvTsP+nT5jzMD/d2yx3fWAZfLrWW4Fan2htldbc7tY/NP
rbPYWytAA3APjuevnZ7yeGjP8PlHB90diBgTCG/aGwwiZpNIgBeLTdjLXbhg
H/W4J1C5S/hMez/0BraHTqR534XBL/q7WAGppT4nEAuha/iNHNoTG5ev3qeB
pEQE3zeoUn2Ytet0NJfpdrCIaVDiV/HiSDALvMg3IYcVjvTgDAgpnnTVqtsK
xNJPthnUCNSuhesx4AgFw2mWh4SrFPfIOi3Xu0zd5GYdmtPX9a69gmOqXPxQ
vl24BkiGJbGdEiENg03atrXa7/WOmjAfg+5PrHZM/XL8NXvzIrbm32qTZ3kG
P7OF4nXyEcFPlY82/9c1we6W5WnzN7BlMY7+PyknEfwWqIy38dd3FnC/XjAU
VCQGTdEbbYwrGD+eDmsXLt0YEdm27zT5QnbKNJr87sZv1cTH8iyZHWbeUVVC
FexDkpQ3aqCrfrWADFFrBeDDrxIt1YPewZyauZH0SAYxjD3fQWis34vQaS8O
AEyLGCOT48ML1l9qYRfFomxoJVMvvEl3hnUfXhEst41n30rarsNJlsS6Rh83
1c1NUdgelTUSmiFCcVhg5UHDmEkrLRsRX6rH4cnLXlw6YMfUQNQJo/66U7dI
h2dQslc770cIosP6/+8fmNMtTe8WtYiHjat/QirPfA1DkerbCSWWW8HSr1m0
rCo41d4p8YzvrnGVNQubSUNaWier+iWDGCy4OUG6m7FSayP0x7+xs79n8iap
+bADD79PIZXBrLMqa/WnEgM3V3jg0odkidTaJ5Upy5YBjJEKxxj+oEre1GvU
BR5+gkPo2FuDtotmVTtdPpWPuq7QFngqS/OEZ+APg9YmP5nbIW5LQXb1Z7Ze
+vFS/8++9AZvb4hqMOoF7fFk5mL+rVHips9HGiBVqXeyiwf/Py3qXtZKJyhm
XZqagDq3xGNK6Xxsi+pg0DmB5QJF8d2psYeTqQ2r141Mrz+RggzwOAnQNtwJ
6ZM45bSKsci8cD8yKzas3y+hdALiMSHh2ZSmqZYumlt5vG3QyRP2sHWCCEfL
bxw08R32o774VfsirgsbarBW9zH6AgyocSojvjNzYIZFAZnCS3Y8tBF3e9IL
4AbZD90eS6wj58gD+yWbcFCNy1GTJUAdCE6V3goU+mxfSZkPqVImqfX+jLwU
t5p1RZYTTwEuM2heKQrmw/1WycIz0/PlbLGn+IyPwnYliJjtewct/xiMM4as
IJZ5fwXRsd37/c113yy1frW3ULQYSIkStQ+zh0sSdN/NUUdXwlySAbilJNqA
4v7sPXbMjAfNNJJkgTFhtKFPxsKem/EBRdCa6H4aWaTSFrI773Y/qdsUbiGJ
0m93aomuakMntzg8QoqsEV/q9sXQ2OrKU1pFoVUm2tdjFraf64H/pBYydohR
gu1JWiARfiy+hw7+1wWAp+LWb45lXG949dlQGE/7E+E2d7DxMtiErd4zgfKO
B+b1R8v4hHDO3pGdVzen94Guun6cF8K4H+0oIejrNWYUDxqtJWlr9NPeL/Z2
DnOn9Bh1x7qk3q1sWc2jEeaokq8UrtW3NPn1aqNRpisTloxLlrARdA3fUGJr
sDNvOZGk1yzI12Gwj8ul24FfqGEZ8Zr9AzxHMhaFhNIt4pE11OCtjB3GoHnH
ecplMlvn7Oqtx672C/fNwq3iXT6jALuCJbCDOBjLwkTvsVf8YjalvePY9bok
3bZ7za8gih2nthmliwZ2Dk2Dk+v5pd5K4ydWfFitU/qjfWkGPV0MPmpcmPWx
OwOg8fBN832elimbBIr5aTMCPgi8yKqULKmwD13H71uLo3P2EM+VlSH5ATze
8f0Q6NW8gnJP9DnyRcmyI5D0nTQCTKZ3Zlt+ToS/cioLRkSLiD5+h6ja+c3Z
AlFsH3kGjzO4PJkfIK3oAcrXl9l48lRBvBf+ExcIRO8bgvhjtKbJ+0fRTFBt
xMkzpEBd6nthbaStP7K8q14zbjvgqwCNl67fKMCDYxy0XNOThHrceSI3I+D/
53Fvqbzi5Pj6cz6lvA+64McWaAS67o8eLfVLknXcJms1DKvEU7rQ9JCXHk7t
5SjkXzf/naa6vUCUW4et12S6by/wikBaS19trK80gLNVDKBd7kbK31/nXU/U
A64jwRr6hpWZJWJnPXPuNrLN3IppeTeWiQdrEWXfLOuqdPymEdYckgyiuAZ7
ugBvMD6KdvjP+SiYMnXecwQscNW+RME0BEkotkuTUKdJ59Tg3oc3lSZv43kI
c2rnidUNcCzqqFixCDipJqQK6200oxPIqR6mODjo5Oim35lNww0btS2WQEv+
Ue8JybMuejm/g/VYbD0PleNMhZ/X4SBAJiyVg5GD2X+a+W7hnr1p0wLRIvt1
Ae0jiu6HwOzdyXnLXBXW3ANOLAtAFJbfQOYHzxZGW7EU/CoHsr1ueTazFGH0
toGHLeaJWSCZxvxS0hsap/+C+5HM/5//bpgf/YjkHB+lLVZVsGPPf//lfHCR
pP7m7+gw1H58+YnfjPXzd0DAiO0Cn6Ef8DuiQeJuUXtDOBoFkHd5TsQWw+U7
LMBWnm70NWppEgwV9025HJlyy+ifd6n0QSkduB0v6JMB4Y+6g8M9FMA37jcO
VL09z9COLWGiMUQJkrEzEiugmypB5dt0aMGGCR1QTTutO418c32wzZyPszzN
yOXzMePngOHkRIp9HRUp8tNH4eCwL0LBFTfTAaiMN1Yn4apMvhbRmHZRop5c
rMuVhDD2r0ZpWbLmsVLnjxhfWxXIVwJvE2sbrd8Xn/AfuscPnRMJKopRvbVL
ZpDxM/LzkcXWuWDvBRj5ByvGPyZpDtR6PmcWBxvEfHSvQvtwDw9Tv68YwvJa
LuN5MX9Cg+bNX3nXJqDZexQ8vkatWKyhuiRd6F7Iwjl3fGYjhYdyNd2nG1Wu
V0RW5QTdqUs2hO5ppDW9cdmAvTBSDDnFkUoNGEfW+U0yPAbydC4EOOPHqRB4
nic/Ti7cME2gn942fgP8L5Od8cLURQTdAgJAAtniwf+/2ABnCbXpJTA8QR5f
Sttt6kQzYzWeJNZiGrEUTdsvoJjnxy/C8rmO/7Ajb159KQGgA6nJZMGlsujQ
FpvYRSUMkW/GOKXbkUZHrh+mtdDlng88+0otbyW/0ABaPHCtHhYoFf/k1Mc0
dXSTlyV+fYT4AUEqrIFiDeDLMQplu+ROOlMOzr7D8ShVAi/yVRvExM3/u18X
hNkZhmx3mExWWWH0a8fy749q8WufA5ufMRJXkvW2SppyNtbyaWOVSL7Prb8i
zxN99MUxC7ZTmvujKp2jI5qDiybRG9YBRvHPdmFHUvHirMkYy/aAqTW3CM5s
3dq9h5w9lCgmIq4uvG/TyikWi5Gj14QUzdcVUuV29wWz1UZW9SuBVNxEcY7R
xlxKLYAqHct+wCj/qG/E29b2nAQshjjh4Hjix8ZlxW1r8JXCij1Rcfip7yKc
Anwy/PnL0kce2YdKA5z77FJbNHE4/7OozrsmOXLN5VL5Li4X3LfY9xNsGTEq
BqlOVqS5l9GYwnsxmo5Vf3cRfXXrrxcTkM2jgeMvMOND+Lspq4C52/+YtCMZ
uOCOKmoNFnhyldAt9ic4pzevh1aqTxL72/6YAR10EsgkugULt5oJjZE4wL/u
yH1AsIQKi1CQyofAI5oicg0KduDGKAY2YkOTKPDgleOKyfkDZ78Y/aL6ydnQ
hbu9F954jDewzBT6R6djRGMK7GmKCAaJ7f8WOKebDnI5coCXaQaZiBvMwTH4
ZaamZ3wOVakN2ssErsgf5NTgyTpIKg+k5f7gy7GJwEUXjSJ78RCGZTTgZtq9
HivSpfgOxNtvOgf93/264mN3CarUQt+DbZ8g40epoekc0w2830RcnakQKfAO
V2Zan6sw+W2LDLWslfcoQcNyGG1xy0rmNvlc0thTCiAE8B+tvL+aYsvTb0Ls
E7QtvgTDCbJbBfcpsotIBdDdp4zIen6INwDZaGS07vj5eHRZX8AfZPQviffw
SEF1Z0Smxn2lDeGqde/5yYiRjtwnLe5cNd/A4UYjVZ2oGJYdOmjEoFuZjUwS
iaDRmGs3zpj4R1AL70RflbiaVPqnHI+iXEOmT5h7zxbg1PX1kYR745RRYnn3
bn/dLD1DuToVXegdEG9MJ+llyJKhnyi8F4JI+wv+YuNQe8TNK4grRQwKwB0f
QNtegRUR+XwzPLDJ6C7Ik5avL5MQnYJ7W02cb9gOdcmfWx8zyCSudNUKFr28
/YDd65JKBm1GmidO2GuNsUqmAKLBjJPKe/V10I+Zx4te5lx7Bf6WxUX4eQgv
hO1iT2Vy1e0gshAmvPQkoLewyPkLruxAZbWjjgvqlv4gG+ReeXw62zD0c4FM
z/E8a/bKcwQ6EqBCeCzkhOccMsUfGQkDs0C6C6k5L6SWh3omN5ydi4ijexpi
iY9RV9szjTTvdjpuDjXDWTK3HYta8Hw1w7+1OtKBWIKt1OP2a2Puc6ScMHgT
D0OyR9H2/PqG3vVmaGchZEI2QCjP/oNNGn7z3bRAHrdXwQYvHBASSlqe3ZLH
PwOpjThJZIlnZzIVLG/1LFcj8c26CPqZsbVTMciwVkJ06BeqbHPF7qF9mQTW
U8Xat/rC8eZcRrq6FP1cC3Seew23UCauJoYjY0HIBNzkexc1NH+bEl1g52SJ
IEK2Pi2OhAySIRQ+pbWB/FehudWq1MHH0kKpSYbzmwm4oX0KgsOIW/7bKKx5
oWNKPGz2tesXVW+ZefUcHZrSw7W6Pc/dSnLPThtHwrBIKH6MWFmu3SRjx2j5
ODp5lLKRc0V7qUYBXH41Z02Er7ab36sLlMtOCkAf6GV1dveO/Fylq8c1XQxI
iOKjOTsPVNLdrgoVwgvpBbTJ6CUHmEjNww5wNRQpateae2p1u6fPbAcxRdqs
miie54NeIjXRouylv0b8cKa+qufyS8Tn4PbH3Afls0Ud8j66SOsXVM1En+FW
itF+mzfWSCrMx5Hy4NOJafGbilZuetfLkuiUsbNOo6k4NZWhU9EqZa+yWdFG
QuXKe07fOjNZtHp/M1Lmo1NxHwCtkSgd0F0Q+bYOI7Ztpsyh1sDGMvLVXR6O
6zsjZmkQbBybPNUL9SbnXMgVPdzT66fmEbh/wyclvHp45Of07BLOgmZ0y/jr
RuAvCB2Elocvgil9n2hBj2eDrhmohKEw7YiLv3D6HYaEHz20l5a1osKOc2RS
+c+e130LBfzOLOgTr623TBGaIRhcAhCU06XYvxNSeJpctS2WsxpGLf+4JLcz
MhYR/2MIviLgo6TyPjmIteHnm7g2L0F71+9F2kvG70LPsWxZ/hSf12CfjKrE
bDxFQvcZZKc2FNzEPMZs7/ejGjrnyhLfH/OBO/ggEy6fD12VrdfB3BnRkdvG
wmD8FPaPa0rMPHbE/I6fY0IXl4J2Wj08M0h++EJPjKBHiIWm4866yMp5tu71
iLOkaE9pxjaJoVrAh6ks5T4ZPgFkKLOifqxSnXfVMTqzHYque4hS9N0VnX3p
2oxdg6/YK1YfyrMwQorzHExcoTKwAaalhyAWU13jmkID8ScqOr7eoXOfPyQ0
m1cdzyl9NtDWzkFsq/Wn0QSjPhstjkn+PcA63nMlt02IY7ecWj2E+kKGyXHo
nuLKDhPNq9kUi2F7lHzKPm/gJa451MIY7F67EETgFILTpTcE9grchNSzTYiN
2DEx5W0AR62WDjqFBr4zgEIrfAZyvQkpjfrmO/Q0zPC/20XzCzUHZiUaoI1N
q9ZeQ1Y9Ab6Zolfb7CDDNtKDwCpQBv/CsGHrBO99EDzNwkhS3YEKJ+F0HjKz
vSmZwcX2HkYeezaaSvMKmq6ec5vbk5BSX4azyR4xBRNhALLks1sAMjdL2tKk
sQsix0UWK4KV3ABflOg5vo/b3J6WZtbMSBG4eFVO7qTFaVaEpGBpFmCHeQde
Ip52V9fs84Yh1Zp0egr8ZRK1CY4+kFBXj6fzp3J+g1yjvVB1di108rAXp+h1
MRxU/mElPgFbEwMk2AIBI14dSVd9mYYnJRO6FwBYgmqQtiUQzS9MB8Pwm4V9
SAPgAbMD0Owmqbiw2OlMza1O9LlAaEWgQPfbmFiJjvdxb6hHTcNXv+tAGZJx
/n72H/e2leFVW7XTB/cGOT0sMiItOfWAXJNUqahrvGD8IcWGbYziMUQE1VT1
qboVa1Irt6iMASOAXd8nZp7cAhK5lPfpotE5pKdETRg8G+OtpdHeykwQA321
N5G5ncFlDm8Eg7IClYDt/dQZj31tuyHBKldyVz17iR+x/k7JFwe3k0G5Dqjp
5kOGphvjyWIo9Uj847Ay/SBXV4+ljdwcplJY74/MkT+cGwQyJw8Y3Mz95Nvd
1nIpFfLDK4OoGcXZwELVzRtO/2WCsCZ3ng2VSz9ZznWiQw5+mMR2DF+mumRR
/FcltdAG5SQmTtuVtrxJRhJK2xnw6rXC6qBBlueyQE1TA+MamSk34Nw/8Tx/
QfOWnB5wLJafYK5W/1yfr+P46r6WHWwpX3RJ1RhwBqAu1IhVU84bprlglM8V
KArOHifi8tg00BRZS2hNO0HH/9oZRHgg+yhYOyoe8/PKk30/u5mTy0RyzE6a
dGMCZOXHsw7wTGGDVZtk9l3OIsMbUDfYlU/zSbGX1GuSVuAbD+jSZgKbuYLa
zPSo7i9uptmuS0v1iITbUyfHEBWok4vVHRQSWJiZ9TzIGif1zmIBwp0JN4Qm
qSOtPjWVxnuITaUcoKxYNrUq/R/rHTiZkH1JQdYmy6fLF16lB2c8kq4D5lr0
r/jqFrl8NgCHwu6LaMoQW2FvlcIiEBhGOjYV6Cjew3lS38udgUGkYFuIuGxD
va9XbtvWcNHZzUCz9GU/swiMhv9K+tq2fWRehC8QSHb3P1BuVMOfb2d72dye
V09Fe4lUBW2i8HdMiWJG7WV8YIF6jA4EBMfx5meZoh8q5+zrvANk4VhcMdwW
yVc6neRAO9s9y1D/8um/A5aYPFq5x5P1k8nXifbkLlV0tBdGgEJiWKOd/tca
n6L+QM5qhbKmkLkyFYeQxIg6aP/E/dS57Ih6ziUyK9lVDfpyfqMyT1W/W3DL
oIRfgmAFV13od2b435SyE3E7D0SvbmWLJraTo3vn6/S0qBgqQGIy7TmcWZ2B
ZYOtXZExsWoE/usADF13DpsFU2+rKTtuFH5YflwzqnTVlsL8pBDb0XRar+WP
9zBWwnlRKA3bA5nCKYySzEM5IyYXbz0sF4EiEbnvbcbyEmmXZfdeOmIb4qAb
3xGatNJO0oV/cGLvIp+uSKupY99CFkGTFOtEu1+ND5kj82+RisMxc2sSyz5x
GkTUn77kYwPL1FQb/NOO2W2ypdXZIt/wTIRzypocLAlVv1Z0IPLVoTh06qcg
s0i8lQtDFrPLDaoqLPwVHio0yrjkaheEpkw8l+vqkhIB/pGTFTSOXNWlF6y7
wr2HySy+FeoUi9u2+kmAr03H7Rm/kGrig+PicVEh8u8AuJAhAETNVdJ9pC+w
2+LhTZIqHRTxBTjXQ2ertn3vdXwPQgn7UEIrt6QvqNfYuKjn6hCuszXMxGaV
JhicYxEjHG+RKBAII6wiC6wg5Wtrx9vArpAVAP0njqIlvWmNO2GlEFgyD2o7
0rvHgggjImEbtUgx2Nn36rkDpv4Mrcfq4nIAgOcmPz8SFZKrLwS6TVC+bd9P
vMDpEZrAivvVfFl70Xrx/ytBdxHBfu20m0Drt4XTCajBaf8fjJlC02Q8GF40
SQaJvDwjr3jrqKKmaTXUHMlcXYbQ8hHL2ERIyU5KGQkUzBKao26m1amqJL2O
9ZHrOz/hBQUdOwWBMMyGGr+21Hr1BR3rLeIe7iCU5LgbZHW5Fx9u8ppCyUDB
ejL9y5GBm8b8gDN/ZRl04gnNyTrpotOX/aRJCVs131mdnxcMSbbsWj1r2y/j
wi5Z8ZdnmGM2jdsotsDGcoo2ZWBvf2BSHBAZVs95cDozczn1/OM7QJ2rfO4h
5er9QIRUvCYdCz0M97qFOwlsCJs/XtmArqs8o0HNgBHLFCyxG/UbIDjsBKBq
lbAxRG+ngwRAl1tB+Jtrz/gcbyDrg1++kacgKaIl9o4rkXK4y0nRNGFh/N3w
94ZGdI4EUeBH9/ImtHfGbj/AroZ80NHUn32GPUbHhyQXYfMdNZIwNcWCtqBZ
gvB78Szs7Lu0f4CaXyJeCprtw0RL6gMMDWo0YcdXkISMzhbeq1LjlKy2w4Br
8GD4rOuBTe5zDRpBArVobqizvM9bwtecPABt5AsI2mVfaQyjRkgE4rMGIpIT
VuCGc3Q/W2dUkQIcP9uojjQIf76CInjNKXziefNbKuJ0kPqUgLUQZuR2gJz2
Xi/+aW0O/7yUyeAbu3L65SgmvqEuXlZEvy1QIXEa7l1NZbf9ncCLpTQh8dLl
4QZU8ltsUhgVzv/us8PvjqCiXCoT2Dr4JWqVtLdZVoV2vZwl2yWNNPDntHWY
2iW5ru5mYjBUMsP1VIZc+RJTAATsK8P5xOIYCz1j5Tb4MS0et8Zy7cQAWgOD
6UHDte+zO5BR8PoaU6Hez1MSw1XWEEZBVBkCuQcXaXNDGjP9pN/dPaRnO9rx
Vrvzatg/tqf+mtouxBDJjB3WETHl+27+B3H0B0qziT93YpiHpXE+fCAq5szk
HXfChIk0I9/xIl5tn2MSUkouJtCQvizOPNbRoXQArbEFBsQwnfqy1rwn7NAQ
03ewhVDUBUVf6nx2ZCZObijgPm9f29LXoQPH9/Lbh/xqv/XNHrwh17OBJstG
wDBIpeLu4ygRgIFr9QPb7TlpkFe2x72N5hH+XUEfAKd2EEoMOD1qaWKKBgXR
p9CVa7w9uc2u8sMv8ZfChcAhOLPpNvcrbZSnfQWl8CDj6byLdtpmM3QqhUl3
RmSDn4BZSluVN3bkuRB7cSyzxo0Ol1BWGrCcYeg8GAg/RRiMDccY0TaijgsS
Db/HIQJ4WaofWXknlf0USe8+lX2EMAd84pHhZu7cj5pvdOjO2+8naS9z40j5
Nk64Jnj+o3/1YJKekBSd4eV2Yak/p5TvWTo+EES3Fb5lTYiGCEGPpqLXeFDr
Pb4s9XIyA67Tveyu7ubxps2ANZ4tjOjUogBuiKFPKCQi1hLKmL9Apdt4MWd+
ATZCEMJFoRiVkccTcUMBdCBxPEo6x56R8dtrpbLcpZPfb7x4H/u/do4Ec3mp
NuRr8IZGbbkcSiPvzRu8RUwjbpQy59JPssq5ZiKgAADDULS8/RAp+mLg0+HS
nOAYE7JM+QhPUwDuxsvbY+cVJAt5O2rvc0A7R0x6VV7MXmCgWjsm0tJvx1iX
EAodcOvMPnOuQVmRTjHeFEQ54zSOZjKvSvCqRihwzZYBUEUWu915QfXWMvkQ
+LglJWOhcIkrn4jbYJf7AFvJvOl45ph3QRwZGdC0q5lJC6Pvv0rYoWIJPdAg
KLHmo9OFOJQ3pxB5gee5+gIs4GX5MrzJGfYNPUnpTQCaLXrJ+t8ttw6b0824
RSYZdkOg8M7HrbSjTvTpoP6khklJ9Y4x3ML5ewhVAvxrFi7UqiNEe3RYwIeR
dixn+gLpEobDiC4rjIlTPx/DIN/BABCJHy1sLWKx2VX9kWJ9QmALa1v34Zge
BumKZZYHCAup3NBy+ydoQsmP24smrPet6InR9e8ZjhLwpvBM7cIgQmwEcdd4
GQg0L6WW7+KoY585r/CGlgwbXcQ0rAN6zlpVOYROu4Me0luDOir4Pe0rIUcj
Gca3x6VSpyMNy1qo2NU/9NNHw91VLlEk7YcjjPrF3/N/U6wODq2ogfZ0vaaG
J21dYU/g3RJUYGH5r3eAF5++vO+sosJ+KkvxLK6W4UMCPm5+6VZzgGueB0+p
Yst5syM6SIlbKRq2fx/Wyo30witkM7e8LlqXu8MLO+TsFw1DvK4wkLIAk4xX
8HzYIIcoiuCGvPqWKKiDRlVv0RvSwoGNkKZeQUQZZleRvDJhwYwvzUN5HuZX
jUDPUeszo6uaOS/empuO09gyzmWkz2dRg3ni+dDen5Vu8qzjV7OG5p5m/CY4
idHiil2eKdwZmRczZqbEtcetYIJfio5kg/6qo3PBIcOFV+opo61aJVi/QRBb
TTngS1cEtzLrSO0z/frbswIziIiz1MJFsV1MM5BYUYM+cATbr9jf93axzrTn
1D9cWzldx6XQV0BM4EOZlSI2+XWOujVFrgkRyI4ZIjSsWxQQiDQiceNdeIUT
BEEbzbInQkt0Y9l4BNtF3ez26j2N4KYmDnr4j9mhxc1ptO5753N2p1P7zH//
S+7kZG7R8wJRscZrj9MJwIIzIbFdWz1a4gLsoB1FOWrKjRttUXV0IlJZafPC
67CP6nrfqgokG3lHhYTKS+V4BCnwRGSCKvVhhHyiE1f2edQySQKKOT/vLKCp
8dJMFqfUGY7lt8pD/DO79h3m9fr3c40R+n5Pj9eweaBm1l/bn/UB2tGYTyQg
jo51Xn1YyLeBS3Qd3Z+H5YBxcC1KNMtw2EEpDLzW8QfJqsBInoU+ow9zfR6b
dfLAMqTv6AjnSxJXaR3f+363Q3OJOuim7FDPv/qHzHRlj4v+REomg0743KdE
oJ8oTX49jIGabb6j9JNMYfgj8uCSpR5R5AADDPIPxaFAWH3d33ZtByJRdw1M
hSyVC2Nh/d6SfVgGXf433DPEZTy7bFdKbYyX2KXqTRAP/mBi6CLTGlsw+UJb
rvvoHZWGDqXWsO1AuYsZ5kUSI+hln2mOzDlzZNnot3pjDGdG9LNVmQuRRb2s
TnZaabtQsqQYVO1STrlMkJ/OFvvF910jg5LQSs2nZ82mcZKQa5Oqo4o3y66T
ZUpi5QZsMSzd5zNnSqQBU78oZd5jKqz4sHgk7ZNpRUoqLVX9XcbmWkfxIBMn
s+YSnkPyjnZnUuzXuL5BI7OOhtVxBxsprxPqQ6oEP40+0V3jrS8B6+WZ5FvQ
LmnVgso3FwFag7i8yQz4XK+C37N22lkpVTqOoJnFrCdf8jK/ukfCKSk8+iva
gTjwVPmJ2haggtvJZyaFbLby30eUscAe7wwstpseGBqYdHARUrOwz6uT92ZR
DIOyqh66qFp28y7HKMhKPl4+afBtViJF3IVoHLS8s3cPChBbcY2xH2aY3e/Q
dAIIIWAwNRtbhQjtuDummdAdzUQOaHVwKbTCdTQSg52qCz7+bHigcE1y+Tj1
LTqkysWX+tNEKr1OSD7SnUq4ct0s9hwpKStx0KAkjS506+e6L7chkDSJ6Iaf
ioCQmd0v/o/3ANeVqKmAYscQEvAMqhG6aBOmew28mujqUrdJJ/INbEB5viq8
APCXRztkhdLcLTpKJ/RS6thq31vfK53kQecYsDTIRkjJ8jHMhvxYUM9rTkSz
4JdopQAMCi6h1BCnTUyLd4Lqboz/04DuyW5bWDZgmagSMYg3LwY4G/cn6DId
8ruVLwHtplu1PewrsbGlLb95K7H6q1DtU04YCyXksR6wW0tBXJ87diBZGB78
4OuBMcvUp2Nmd+JC9J0ggVUsYeUE+0QXk8ixpPPLwSjmvjr86B/cNVcQV8vn
SLhg7cluR3VFIrnArrP7V8EehpzQUirAm3z+xXhlclUMnkSkL/OLBOHsSn5a
GULPxqdFVPIdd37074mhCqjevr41ICXNXtmErz0ZhQMmHwfbmHW6sMGLFZrW
7aqtIJ5h626dsdEiCHISwdk13Z9avQA1U6w3e5EgXfN1oAIsEMP1+TJ3DxpX
iEJIZUZZW0ZHL/sUL+14wP1IJ3pJFKFTRODB51aeBNkg1dbqId0kTCO60sot
2dfXi363jvllODNwcFYDA0vLTxteGpG8EzN4wY3/2iBe3W6GcNcMLZurb1RG
iToMmFfXNKpd5NnqtkOPwFb5vRpL0w7XB4Mo9jPreD/6cuz0C07gKAXtHXan
WcOyh9yQ8rfQucYNYrHgzdrduxQRRozkCIMRqrUNJfUSGGnuVO1klRucAKqG
SLT+SF0HaTCovcMd2bvSPjB/S4apuLwMbUQ5sXIZYP43Vh4pPGVfOO+buaMQ
4p0xGB4EeXzBvPo+rP+N0rjqMXE+scKIBLANEb55fCJIBRZLf3vjK5HwFe8z
lVM+OFNqq8ZdVdKWnCdYcVhEFacjIVjLu0a4qusptFzzz/R5Uf7spDm25qea
QqPFSkn1f4Px4045m85UJHtO/iki8FNrgskPaYqdN3y/F1W8sFZsGwaw+kVa
q7srZS13XJCmUTbAwfArNTL1Pti7Qf8bPKIto1VVCBHyecvfILSP0pHI5Jpk
AWg8h2lHzt9P3jzhXIzgEiDAoEXqU/P7gt17FsX9mvJKJn1xzA4RS4sCrD17
1EHxpgxm/IySjNjr4P2e8VdKffjgcjNEnOl/bvvaS4A9ikeTdYzoO/ZCFcEi
xzIXE8QwvNji6UDDClbj+7mDggxxBCP7XCKcumoCPbv6q/1MbCiypTTfx4bn
LKqkhlsa/onQLNaVKab0nKevcBDL1fAY0f8ikccdnFSIK3Rl+QHV8fwlXYj1
LzxL4AtPlmxHn8+68dnDdbrigVegXX4P7nwc4pJVKzRGWNOWCMQrBjM0Ijeh
atbTcdqDkhyzCO6No5Glm1mro0BtogdQtKn7DlENhc0qQ3WVdSWd2x5ePfER
O4pr/0vZOxch4tqDOoVowuLc6Gci2++HC7emBDAZp+f7yaUMsRgRNQozHSJ0
XNgbRIc3nETnJXK9Mt12JypRoZi56xECmVZLpHi5vLL6IxFTz4F/fhDvPFaM
KzUXHC62GZ+rV+jqN7G5QzkwZkT8I8F6vdBbmyGjAjk5tqK+7B/2j/uzFNai
A5TemRSocs6tYQzoKok1yqn+N3oxy7jh3UvAi78wp0YmOaEAOidSgStpT3kv
/914Tbnm+ByLpquDXqiXc28nkm3P6zMprVILUu0C0qRJrxOltFBJsnBkFGFk
zSWshj6goCUR42NazXi+scAnQQF0HWcx+sKR2tuggWj+yINyhN0Pwn2H/WVx
xKQNDSYep6V+UfUxKihjoO1w4Qqbf6g7CNkr5zlGgmqeOL19xIJHxGkcJ80c
QL5xlPQuv7jldczSP4APLNIA095qj8Krbsbru8SB/a4sUV6xqnKPFgWluefZ
6NBTu2P1UcWHB6MlupJ6SRqHa0ZHGedHEPQpm9bjJWVTShixjdZtTD/prkUX
OGHYn2/Ih2CHw+Mgcca2hbcWrj4TPyIb0TD1NvtCESDO+Rp7LHui/D3P4aY2
UzouzMpULc7KQlGR+OzIxCIiVoabXUvt3XbkRkmtIE7+MRQzyzJtG06Oo/id
x3Gb+tpBnKuVaYo12m2tKratdXvEfGQKcV+z02mFk7UVhVc9u1indt7N7kNi
m0evq27uYGrtm+lhDmx9OnzuuxE0ualpfT+aKCy1PO4iGOIavnY13GRnaCjB
6gZ1eaQv9RPUcrHRLl14d6V4OmknhfuaJj7ONhbMHGh0ua/oluq7sG8qztcj
yNyPs198jy7wrjATZDYkinLrd87eJgx0Es5rTqlUVZ9QP7XivldIJx31iE/S
llM1QhXV4x2nEVeAvDW72pIRshXh7m/LG1OG9xGKtZ9hSoJiMd0gCumduGET
qoPcCgOJlu+iJ8GtghhL5mlWU2oV2jQSJfmrBxpDdVfuIXCWX5Q3pFtLsu1x
L7UoEurrV3yKTG/zUD8nP9j6Rcd1ml70y+2dHU34c4rlPwwhrAKe3OZlU1O+
h3xOVSDRUoTx/x67a1S8qBgguQKXP7+WawHKAfdQujJD7s80MBf5Sg8z8Kkx
m6djCmW8UH3PceApEpZEVS3OoeQbxcgUINdMlDcc4s+Ld/YCuFRZ5Jdyf/Ea
gpDQWNXEVL/DYHZxScE3zCyiR8XFgFJOrEGbx0/qVAG+qyCkoISj65DZQFFU
0piuG87aN5rRKl7BJ1LtMGoPwnVB2Dqm3oTuBRvpTSwHByYx9e7uU+AnR13s
R6PQDFJzXUOgrn0lhqzOJcwlFyVShOYjSElkC3Rzw2q9F9hRExg7PyaXYabG
VzkL6nQzJ0ftuMslvW+O8zLlXJJ2Ft4fedkfNRE1HrPcndbPrLWw5UZBo3Fm
MoLeOZjh+24lN3mbYXMOVmzbfKL7xIqcCfJSyl92MGDyFuiGAxUVXkZB7IJk
Ah8xBlDMLx9xd4kVoViP1922bOsMyq7LH+IRGHippooVtAdCGcMeqCt/8Eeg
yOOX/WnLMffJQegUCGV0EkRFhPrLWrPgGBNgX9WzT2LorXyaSKAP1yaImpO1
LHFc8J/w4k3pIZqWW1if3ZZKDQq8Yqt6A7R58xrOBmmRxhIVpZ9ab6ymouW7
kKCt71eaLuGkT6VTKAsxKi6i3MikVCfCZxVC/gLJF/fnCHYg1f9Io67JEBmz
WsfveWf3AV6FrE7BssvF3yezoDk9EHDQ5zTw3HI1Igrhu6+CCSLUoDdg3VzP
vgIundw3FUoa/qIXGVCCbK4CALePFaIjPz2WXzeamIRggQ0B/K9DIxMYAvx0
oYlg98mqKaNxcKF/h09E59IxW9RcWKvlt4ieo/w3oF1iuMiSil7Q0a0ybk8x
Dvy3R2NntIA9SkugtfY6Q/aca5WIoPW2WBK4Vgu+Qd8gz1tGS/mt5pRfKle/
PcyLBjMeR/9Se3VKFRYZZ4YE6jmu8LsXM0RKTZZc4U0MUKCLKtIpIZ4Xy5I0
IWOAe0rolDWI1ieRqzq/eOEOJrBVlOPt7dAal4pTCEpGpVXoUYOvou1J8IxJ
uXcA5SIzHCuKgxhgfdTBvh2qLrTS1oe+W9QEFlSy59Kdw2CrlYJ/iJJxGDkN
Pf9nBpsooEGfKNDyogayCZ3jrvWzV59IIz4u39rsM9H4ccR/cCoDGszzM4sK
uIFob3J14evijRnyV5Dr7APt4BvdFgBncgjjlKYe6bq93XYGSZVG1KU0cvl2
kwVYwDTMU1DroytzRlYYe6BGI7zhxepcGCHGhDV2OqpMW9iHDMa4LlmSF3gE
D6MiDfhX6yLlM9AECSiY4veISL9cECSHuEf+2hO8f1aLyOlvHNT9Qv3AE3hi
EhiN52BU/dJp9Myc8rcV3CRG41cBzED9o3b3qFaRfWZVzjiFoDbLV/FUng9d
iNaOg/onrqcKJu8iB/5SwGYxmR/ewaBE+5ox6zrS9OpvvAvl21ixlKe8JyE4
bmZOY2ao8FBcQ/qJM7DLjWJMQrp/CYK4ejzns2c2QqrmwjGWIPAn9yKWTd2n
ZlwwQtpKvI35humRqu7mubKid1vUn71maQCXYfvoU8JDv0G77D0rVkRQGU0i
U5Z7c7eOeTnGt0vO2ZgRXZ9iA9dOAC+GuiAbWI36oA3WZtih1Xqyy6UbJ9aP
wfcpu6LFEuJM6ujVUNPavF1wNBV09zC9NcmkhhLLghw+KtRXJMQSIz86wxaj
W6PfRMS6NeKUMplwFEdu9QnmVeWLQKp6vI/Ys1Zuw8xRaQpeF0nHKi7/rgMg
5b1pbvnM+9A6E2pkdXlV6LIW8PekFc44TaLwWwhqkZHlVC0kUm8jjqcZdyaS
HAnsDXq+v+yyCdaSbbYDc94sNWTyWunrW5avbp2mg7aFU4usdPo8jzWsMSjo
Ep34AHdnIrl+II0tqHscjKOFMUfVZ9sQmtIJAi9ZeAE5oEXfKblYYdf6mC9z
KlOYefjiPl6/iOqjum5uOGLYxFGfjzaR1aU+YXecuFkcCDXljChvOLMJ1S8Z
1gDIXD34WsJ1Te4hZa5OoHuur+ci4QWUogwi4Vfts7WZXP4CHq3MuF4cl2DV
lQLRaKI3yUzGl/urIrJzXHKiemdzudq9K5CYvJxH3Q4GBPC0bE3KFg/IJOVe
ZeeIsblYZ5j3v1AgVo7k+mWYQaMX3RS34NRnT2cuKGzQVzkdKd3Jub9jyt26
wyT7intsLt37rUv7hoD/mtskj5Q5JLfYWGqss25FiQQNBXkosiSNAfCZMnpr
VR3UPaQD2TCcim7khNwCog4O8GOvLvvxR2pDgDXO5u+psd0UOY2BfAisEjHp
hoybqfaCtvPvuZU6X5llc92oizcCBESSPRqZnnKt2NKrM91ZRn8MKcc2h3YN
fnCB+FXh5jltUaJXAitTrTRCUOXRkbfnsjJy5Kjja3C6F2Pgr5h81oQ2uqIt
iE7LMurhbr/ulEBTOWppx8UjXOplUT+E0GUCItdfnbfutTq3mD8EYihM51QK
uHhguTHHpJage+B4mR7wySKLLnucUjZ4nNV122ah1j2wWTyPzer/pOxF31AF
b/Ev8lAvY5Ajf8JpOTfsKzbcJkYnMYZUZesSG+LJreyCq8hP9FxXQPyiJqsw
MeEYyU2xeOTNDjO0tbamqdS3PerhZZBDuPQZtvehJneItpSFE3hF7EIheihS
0/7znd64UFtfBXXaO8BLGeSYUd0KGTN08YsynAErNYltptQCcv/VtZBk6hfV
B3DUm3B1YdEePqUPSfepbTCgADbFvmeZIIDm/bKLV300LIQ6lpQJYE48dDrm
dFFEv1jS45y8RPFsOx4bMckA5qiAPDOmq0DKwgDVI9/oV76Xizh4sEyq80Ls
PW26R8ts02aEQxIPfobdwDItWfyeJe4v+fa4Zm7Daj9TacefWO5YoBVw0UvL
/+UalT1LbxC8M9NgAQAiMCxcGjQf4yRF5ji3b3eVhVAoJjBz6LSsKpArTNVH
KwlFpkBQcKBq2sUpDMCcmArTYnWp1TtP+ElRN3nwA8i2yhWb6lDnqAMv045t
3hZ/ACKnhU/lOIpblgc41g06PrvJIwN74Q/doQHiA7qRc0zTT1qBHLAz3aum
mZFvhVFmx8yG342cYfbX1TMtv6gYl70mrjY7WauaD+WtQs9tC8w8jT8owdUL
EuHSSXPCeLuPKttytbmciBlYWhuMce5qBrow6FvzbtYstMznMR8/Riy3M1gB
8lkbzzNioL2REcI95I5EUCHrR1XvVcaWyMnn50tuiVHAxcmR2vipKHla1qqI
QBUd+O7gv4BjL/ClUstnQes3crOA1L/kBwchSWE7DwWf6KWLexLoPyoiMgHT
xLw4r8oJWfjexdMZ2wrT6Ex//TvA5rLbYpp/FndCNSEBWhgxIurCGDS61ZT7
l8OafXO2gEmiKwSc0rQ1aldipG/wMGlFv4cnb+nyyedjc0T6j1GPaWRVYRY7
NfxdAqDqnWJxf3NBSTGuQJY4r2rDSKhg3odzr0om51afO4ZSOjgUyA2IhPgg
Zf4Sq/uYbf8wP+cXEJFyYF7dcN2gAUvV8y6F3oRi/21Rj7yovs+fCEBnCwtb
ALT/oswX9HcnyYtwuTmPnDK0A5+S8yyE9bed8ImfTkZWDMXz8oE68N0JqIuS
X6aQ2KeqJczYv+Qyw0ctOOaHtQnAOQhiiZgWDGvayOUxcelzx3tQtgDqrjq3
gDk1NPJ405muHbCqzJFhvQYfK41mFAWDD0GfdrrJVM9LOaSCQpBDf/qM9C+v
M/x1f6YgROHVKj98QzE6oSCTVHYijPI6R+cQYvjG0gD1EgRA5RYX91nuQjSB
+LKV5IERnfQ19A2MKHW3EcSfpKpA7MZtcuLbeKWcj1WpDoZNnslX4vICTaC0
P/3Nji42kXeBnB2XuKL/CISs1Go0bRPs7gg5uNOvDTemYhCAkt5wKE2PASuY
T0XuwrizV9fti9k7P4Y/Ae96xeeaN8CeWIvBT5aYX71ueNCPVp+Eu7udirzu
sO8GotgYhygnuRfRf79UggQvpui+ws73iyzJd80YE2eVOT/iviwAyFWh65Q+
fttL7CNsfrZ3OAzTQ5xkofXsub9qFm7KysfC2VVj7WiR3CkQHXBvNRNkJzwF
BylO/7QFp2gR3gfCAmaHFJXaEtqjK7399vHR6qBUMnz/6+HyAyr1Y6BgfupX
6w17nwxDRJiLBNYU9LjSQWltudbbu++pS4v1yRmj+/pNyrWzsHDZe0xKbtpK
FRH0BanR0QaoYdM3+NqeBcqzzTCFbEoqv/HhBlIsWoqPSDUSxeOkAPcU3Cu/
ZeG0qPgVnC7AmA1D10oLJvy5u79ekNfKlUtyjSYE9+48JrodLsEJqoaMyxdt
uaRYZUOgtLKehtdCbm7fkUsIrDPHCnL+dut1f718dv+gNMPahkZIF5ORlYuV
vlYOGFwG/K9m24K2Qf2l/P7y0yLUpDxqmM+fRYG/0KhadS0/tFSUq40I7hKG
A2kPWURatA94nZCcqdexfsnTlnqw80Ve11owLb8HsI9OkG2xyh8bO/KQDyGx
tBediaH5iCwYXozvGL7UJwgLFwQLih0HRk/wEAqQwqiI3F6v919diO/EWsD8
JRO0J3vS0Cri0T7YPRN7I/SD2O5IoF2NGw6bT1QhWI4QUz48mrtBXGVKCeJC
UneZDPOb0tovp/eqaNDI6zz5JjlSNKDpcJcgwg+MMUgGLLexr9QGsV48u9Rt
sBgPSTqensJJ+l1JpDYIgzW1y8r5yVvmYya52NuXQ90VRTpLDGXgHWhRRhAV
BawqYURwe16C+dP8/aGeYk10nEUaeyC6UHCHU/LGJZpf0wmtXPnRfbt083cY
Xebn0C5zrvGUSMxD+h8km+cycflwa/g1oAV9k2wAvAo45UKILObmuOn4yeWS
xgHy9CRh2ccjbYztkw9nieS8pEmoMelaRG2ONYTaT3UArirbVY7OKrQDIiaO
gxccgE/YMdVwnB1h+Jrv4JKQexVijtB9l6pPNgvdZvGeyimaRa4OlcNmOQi2
SGqG8iWPYkaGD3ik2ppHOhrags0gCxStHA3piwCQ2T9v8Ldr9qHF9ibI29Dg
O6yIesFThQDyjOT7UK8nA1/kDyI11MS6Cco7nYViXlCUtIrHl1h+SG1sInhj
SGdNC5YakZYyU+c60/+IteFKD4NeGQsXzwEptQSu7FJGZvUJmu0EKacqmJ+b
GI1KgyBZaZip1DwCx51RFTFhQekJKo7mWX6ZJuHtRYaamSBS7ZVKpArq65wR
9tH0JvjrKuhMkbCydAqlvjgJZuSS5mz4cvHjiO3Vp8VsUhumJMI7lYTml7Qb
qLzL5EnTcOn6SqPidZXwegXWgqctFa+/GHP1SjKv7m6ADfs9fiDU8SSj9D35
ZglvYB9aX8Jt+rHABLNf9ct2tkwOpBtEMJlot2NnwKji4n4WPkE0vhFJDpyp
7KJ/r9ZrdHYNBoeMs+L1r1Je9M+n1FX0LAJP8zu7uJvwPv7N/LCZPjwLs9tn
/lxq3/5c3+X/DX5evA7rCIfEDpBAoo0d+pjqMXipOtl97SunDY7JNDKTfy1F
g9VgOEHkiTfkRoyM4fqNKJhk9bIcI2idme52hPnCbQ4tPe6c9M3qzwx0xqxm
I66zFMd9kkrbV/qsPWSGoii6F4d4th0QzdU1W76Dc736KlSUtFNwiX3H2iNe
MOZt3OF2YGSo/zAPHES0x5cfQPIn64XQDmATq2KYkYQJsDhWidBM7Y0Z0mfd
xdFXRudOxjarqZRN6vo01+VpbpehjS0IJ/pZDV+5L6HYuJpe9EcR9zEvSWHP
wPiGkOjR3KchK9cJ1tZrHYUrAMZ1pEHStsa4bIIsYzrYtsTljQ9c2CM0MxhQ
1PcJWMLBrIPCT4fQgMZ/ed1BlU9shxkBTuXCHyBRQdKTCkkuZDbT2jS1ApR+
Jas1xnwwmbPmstcJ4BaALjg2NDptIUzLxE/7RFwodlO2ctttAMxNznWxUbcO
Otf4qRXd5oC9zzaB5c2ww7rqErtTDGG+isYsp6+ag6dW9Ad7qAwN9oqaCh65
WyiCdZJiTREcPf7PyeEvy+LqrkTW9Ahay8WPRaMqHfVBZsPcRd5NR2VDCS/h
N1R9qu1L0xeQx/7GzDVo1u7SBtgHqu6fhSbbcTTFAHgl6oiDiXsxZMG8ZblY
dgP86gsHoiU2mZe431D7NkelXNs4iWhE4tNVrlT4ilfeavJVau46Zw/s/Juj
2FMn5uo3rudjU89t3yGOr7D6q48MsIeWM+gdIeNBpXZrlSYlj4z2Nxo7CXS1
paXc0Wn1DoylAoO2ycUfLnUTCpzKDqb6a7MnYWhVuIRAdK2So5OpGcxer96I
CL9YVxfl0bJHsytCZ0n9RmSO8G6FLB6lteVBZHvDLTl1XB5gSVAl2TWG6pau
GamqRMGzAvsunw7hA5+7y4ECbvWUCVbhh+4OI7lO6mqlHf+55ssYiUiFM+dt
7vCo1+RBHTg/c2qapbW4cESSgFFjT5W7v0cTdGkxAbu4nsHYSaC9GF0eTGUt
AF17SoXJ6IYjkSjBRIRRVvNm6pubFSlRtJM8cp/rEo85K9qj4VV8QsKzHXVw
EBEvgiwd1quReeiI580L2QvAiQflUPCmdM6Ohh+AVdpWVShjHzLRwErCdTJg
Xe4DA/nzb7I/A2rB2Kl0gg2+W6o6XZHpXgrTf9UXK0eQ12gkjeQ5huBn1ar4
bumdiOFMDwd0KYTS2TdVW7h/1VtPLEc1ZxQeaDkeP6eC+QC71aTtF31W17k8
luxcvIrbXWyEImfByiVAij3uykmCFEyqIRFNDVU3KsW8o6WV2GbqcWe+tRuo
KRRatjUpvZpKtlxzvHp+EiDtE4TTsmeNCz6/EifcRaiMefeyCAF0ZM53Hump
/2w0CTsbGDXHlxHP3iilK3PVukRl6TFkmhHEUz/bwKhNkXaptevF1or0y19Z
YD+lJ4FMPVar332cVF5MZLjKuu727rK+g3/HPB7QhWrtoFWQ/c8N+ZFXFqNO
J7Y+dV6Hi7Q0HEiwfRGwVlAD73lGmZhZTm6SertpA+iNS3pdr0JhWc+aUfVB
vBYspgBmr6e0pe8yFDRZuEEnUP2Qm4xj3qsDb866C2jvBAQN79bOQXaBEORC
BW7RdYxTPeVTvq2C726JAa0SOuXVOJvTXSydLWfXcrFLDAmXDJcqis1s9wtA
gkIE7Qzh4KoZXqcLX7qbL9F2j+Ey0Qq6dwwag4OAzb4u96iTBP86iEVCjEzX
Wa3xSErxo4IlYu8Rt1rzRC3mrClpRX51Hla7VFofnTmO+ExOTmSF6ggVGcdy
C4ZcWM8QhE0XOOkh4xFUoxYOnoxo0zmIR/WI1HdKzdi3BAXnkWNEPaWH4zf/
i/5QLFFIH53DJPEa+m9eMUjqcf2Wff/aUM56vEtf9ShRspniIyGYqt8ctg6a
RkW3bNS6UFBjI/57mb6VsnLIIV9ARD7uSPfdjoKKbKwyqlJ73LSpgywDBYsr
17koU1LRd0rgjwjAr9sfuL49cPp82uFx+NmvRrmN+VxXtmjMrCnIEaKk4RkP
FMg6F3ybRd8HyoVj0fY/Cu8IQOiqq+0XBuCHeyys73zqT/ZC0qJAsC6sjfwY
TjQ9Luf2foyHZXxaH4MeTeUK5uQp3UEp9C/4mtr/tkxM5k7ObAPYfbakv4h+
nONIMURLGNH1xzIXfoqfNx89xIZlJ6TflddLQfpPsRowuTszC0sMQ4skN4hJ
vMVgOc7hcc4wC1iqxn9P3O0SL9nxGepkSmgPkUT7Eo3PHt592u5apdWynkgE
9bWbk2OaVO8IVDEH+Pqq0IBxrMP9KURixTqBxDmmA6v07CFCeuCnZ4BAvTot
aEuthj9gTijttBL6atIxeibBEZnIDd+mZyS0mFTgeRMI3bIwAqVEps1c23XX
91o0qO7ERJPNeLPdhnRX0westaOmpt6ucVAoFD+dNLjv6+7b9CGumtUvAdn6
AZ7CTuPJ8BGGC319YfsiawFEwBaIisv20wDZVbvS/rKp/oPPYDHj4qMpbrgB
3Pu7f82fLVw69qo2fo28wTDThrrQc1L+BAJGSupmVic0vjtcJ4x/FiaMao0P
YZL+orAMZu+1NooFwj43RY58AE/YrbMAr2AclzWl9XmIhKTxTZMm+HDsoz0L
TqWCzZsmx8mhxGBnCHwy1VqswJqs1nmZ+NI9p2lqo1eCNpOHzNhNg04Y0fIT
iwaV/cHH55Ki96GIIQXRGTW/nrwBjL1LzsVdJXeTEaNSsZtWjh0RFBLkFZOW
EQUs9B9lWvCCuSLhKTe/xYZCcNVzM4ki8GZJZWqTlBK7gOGk47LslklZtSqq
f05/pzosNqV3Fae+idkSRr6LjIxwEWcTl5hAtgr/YknSju2lLbOOBVy5Z7OJ
6jCSSyjK7IR2zWIvuT0L9rJU6AoetzuvTRjjHKwkpA06nGvHQ1IUPVwmasEI
tj8jewAoaCD/Hai3ZTolx+fxWKklMS/1SPD7u8+tzV3I0YRBGcBP/HTvBHWy
Kozuxao+wUfDKNkM0wVARa1/f6ESLgE4VoToJBd8mK1RCAYIvPQP6kW41s/R
hmoRAcL8H73FdsTkPF3QgjMIEYFIdFnS1O1AWhcUJH9Vo5/maA2UzGaIMUSa
LgcOs9vSpKhiJPXG0upN7VkPvmlXa+bkjuy9i7wIS16R8s+0kyJZQmTsIVpF
QasvpaUCA3Ube0lta2TQvHskYx9fqcSnyenHFJTeaM9BBRmbTkHMC+wyoo4C
C01Tk+nMiGZxpx4rMy3GfcVqItvKwETgEwlm5E7e7mbW4X+mq9TXC3IG64HY
judZZ6TKdW7ojkhSIdY1L9ETLOFS5tZ7ZKBkjIoORkNLseLuexhh4hSuiXWW
o9l7L6sIYqIfPxL1FbemR5cH0vnozUrS5e3KLTefGyECVxvDMlG+W+S+30OX
R1mcmnq6yYny1n/IW6lhhsXmv9l2q+f26nzzA6MbjuVj37VSREdb/MTLSmiZ
7NF27dAfRCnj9TMX4KBHdRJ6QxB++zuPIsHVRChGRSQ4R1n26rjrc5T6A0h7
paLb1s9ugy7RiSB6XYnLA34SdYoGiwVwoxMHCYyDU/n8+D2PjhlAwrhU/9uD
85/hl5Cl24iOOfctr7dNT5hbtvbdbu/E/Xah3ClLBTrPdaaA2cQs0QZTA2DT
5HE3iDqZLgdCmGPwLWK3m4+o02PR5c55XkxJMb79kE+2FMHoD+sodswBFk2e
O3vnDYMWT9k4qjU0saAw2AWfk3Im8tIuuyn76ThMSIstCsQ6ggpn0KMt1kSQ
Bapztp9kfL0IpiI4nAMHtAHrDq+BJnm4BiHQMX5dYFisFgKanz7iOiD+wh71
Q4tQa0SO4cF3yHi/z5FZrPZp4ZTls9Ur7t3y8rp6piHb0siUE88zeJ9EtrPk
HwtRuiiwsdi5ZXWXLHoqYp1jV2Uy+xkMu1Ijjo0DNhDy9sxP8em/NZfyfbG9
OW1hrPCtRlmvjp3VdUWLkfcjJFa4/4U5GMDtrXNrmpE4hAY1oxvSiaJez1Oz
TBxdz7Lxl4bYFfc6URSEaZd7LBLbmSCQETlbqQtLf6qN0tItjAy2fmzauivo
OuAS9s5xcj/IstZiFO7F5hPhWQTljWa+t5vP660lvKl9QkPd8d3bl2lVN7vA
ut4qCOuX9OEVCJWp/a3q5y+rzzmuNqTFY9jBAtyXpjsXgI9GY5mo0EQGFkjV
b8YU71d5UJ8sSYjkwseK/HwFpK1aj/iBtjFf0YLzJt/MaSlRq9Tp90YHK8Rw
NfQ9HJzIOXGt2bVcTCN3DSsbpbRRlNo1kEChZYFMVK063TjIuuypOm4RNf6u
itQeLMfKor6kYYUoBFhp2O0SiMFnk+khwBlDQm8XZusbB3ba++nN65rPze4H
46Dmg5guFkdxNLz4tH9nvgWrdEgqid1TBquO1u1PKigdX0UeQlG0cxx7l8CS
L13pDMyF3F8cWsG0DgrahBrieFLjTQySiTbg1nT4pa4kX5Nwjn0MEy7Dtn9h
ym7kdOZw+kJJRPBtJRfCky6qHSwkuA7ZRUcGCp0SbsN4FyTo909fxZl0l8uI
a4k/tE9w2jN36z6UELqn9m7pSTX3Uhrn4TL90lPl/u/3UcWscHdhzoNM5A4J
smY7TR01wr+cUT9EbivqTSSo0NIytBKh8rxtiBqLdadXChKQ04H6QLktr4Ow
pFxNqJ4pBWMPIWmmuzOOPuedYPHiC6EbKirYZocTtAGI0xkv8AybosNmMXWe
CcJh0lnyC1w4HYHmEGDe//YljhspZ0K/EWELMVWrYXStNCxX3yO2Hurs13Nf
jPe+nHgJWl10WiP4lB0DswRaAGxEL5J+AskB7xdLAp0RkWPo56QoqlvxxbvN
hZLS7owh/r00dI8Sr7DMGCkyYnFC5CH3d4OO5wrAZtAvPXR8EmRSXjW8lijd
31rKcWLCHKX1AeGGzJD6/5g9WjZJhAuhFbgLq9446o8ThqxmUfuEUhZAz5yF
VNnjg0gV7SrcCSWlg1SU5CqXlffj7HOQ4nD1hnT8a8bCeaohPbErLZopma83
YPnqRimOCqSPQ7xxsYx0S5M+NxTa/wrIENa5BdtYCf02UdMIVd/0YT9Rjdig
cJy4E7VvWvukKuM7D6enO1y8NHRU0RAzvvHdJN8N/Zce4FfF+fsmHF2pviWV
wFNOlDYFeRUZIrPeZq7XxhH9f4C3yx0nNdXC9PR5pcvUHtaO/kOe5zLpBlgO
qNn4dR9soIOKUq4p0PGoIJCCcyQUik6bIv2jNrkRB/9VyMCAFROTkxbb0Dko
SOYfH9o9+IujaToffTToh0t7GWyuixqEn6buTpsWDT2QODdmbTW6R1qYEYa8
7FG6VbHwLLEbHU/g/sgVVEpVJbFNucyne9aG+tbH7FyWu+G6MMPCZ/1Se3i5
P6OcSm+8om5HuZXK6zxAI1Ne0+nsfB1heSZudKKKIeMM2V4c3OnP3t141/c8
rHxsI729Djli++MyO9F8y3QwSnG3bKZht8+9eH80xRevj8xPd1PdqzJFE9pq
yFoJfhZbDxNvb7G+nQ8oMC6Ls474DqOs1v5oF1a9EpioiKkJXiqw0H8OavI5
3DQ/vxnX/JudNzsqley7XeFocaKtmUDeICLzLJ3Y4xrDrkDX1cBiNbG/HOTh
mXHAfYzT6MgquH8Wk6DSBdiQ5v6B4KQtBhwqhvLoFsvjciYM8h82FrGeTywC
A2Jcviq595oxPbw+pQZKVrJvZ8SyGvXBnpSKV5ep2OPF6YZ3FNzck1uSEHp6
i9gX3ije9rqF0CHvHwhQdhYARKepn94x3O9NzMddgI10rBH1+rzzlgl82gAH
58reJStBl24ngDDVEb5ZsWRr735YaoiwG2P4TzKUZssYYW6LqyMcvBZvJ5zR
ceefecKv8itgS6gpxB23CYQR8hmjbS95X3Naey8sjFJOqRVOU0l9ebAMwCot
EVv+onx5H8T+COkVQw/YNhy0jg7RaqvyuDZHA1UAHaunpfCRovX+rXKMCk2T
Tl5TAju/axUfoxWBd5/nyyQtfCksMr6x0k31ez29S3avRDSzWUTeYCWXnHsX
heVpc3tajiks2BYvTFbBB2YGSANB55RjO53yHPEotYvdfORYyBGteWqQCcma
2mDeuD9d8AGmina+CdGzc/OVpo15Z3XO+j4inpRqgrkmftX4EcjpOMqA3I5Q
MRWdvsQb/EoR5gruAA5GNkODgDTqrP8r8T7HHBR+nR+tYYyTrbofwL6yo9nw
mYzx8rYuTjV9Y09761uTu16LCR+T/SPVrZJoMseeFUqp3yCumUDd5+h8EWPm
2ko/xWBmFx1MEtPp3+i9qS28aFmo4e5bNsgXiI290jfaw+lVINJ8Xyf15FJG
1V4yNb/OhZb7dID1Fd+ZwzVWubxAZp866IemBxXNRDa9zhU1y5CT3zgf0Ggf
MU+OwdpNoleTm2ht8msFjLE7QATxYVTof2nneshu6xHpwfsfBxV0AJbFJK5H
ljLDJFWehMpH4RD6G6cMyL4hmqXcR5/caXwtjGUBzdN+rBEf4xX7EdqxOwcM
3M+3vEHZHLv87rhGDdfrxyimx7IeE+MhmU6ROcGcy97AWuSE3k9aYH6UlevG
sjgLk1K4mNaHaiiwk3I1o1N0GxXnTkmbAePA+65wtp+acLPn94LyWbc8pP42
TLNFqLSe6Uy4EqeJRodOtCr4mkPtS+IWIbvgEJX/lwHlAsNUlRXTmzN6nWcv
OsFdyKR/LsUKt7hGM+2dxR5dGhEZQegmNT1kgABtxFE0Y8ILT5wZrUVVK5KS
uOFlKjDP9kHmmfbX0o82Vjf97YrRTG2DBiAGIdH9a5tUHnViI5E2FBMxqzZq
U+NQ8grAKz8FV+B8NVHPApa8At7JO5d5FSroOqbUSMInOKWVTfjO+HNkA05O
2xVuaP/IjLhJRZ6XaspgEXa9xXCra37cNBchPn5cD5eCBxqryZLYC4eDZE3b
CgsOXa+r7kblP0WK2CnHeDqk1WYbI0UHKHDElAOnCBp7bZSu7sYO3ogJ9p7e
P0tap7CLvFvbQK47WqhpetpsPp+/WtUcflVI/xLXkLQtVzBx0K0oS6bx2sm6
gNRIz65icAeWd35/0sip4MqxVlv7jsi3XYiVB2hKLmIMLNqR8tlqTtCDU8i/
Ji/xQH0heNHeiw/zW2wNB/VDVAVVhN4uVAnnNni7dlvU3V2Sibch/wxYTNjf
ITuZnKBh8M+lqvdkA9JFyygXOHHm6ehNVcuUWklo9XRgeI9zamo0aZzhAptE
AwLz2uqaZ+qBbPZ3NfyeJMwIkEx8+tULORusPnhr6f0v8+UmeJ4PwGLbWNGI
FdPvVnCx+gIQEN5vOD0IkDRbVkLAFx/g2wgofCjn8ZmDJtZSq2EExVD39kwq
9Sre9olhD2OB/7jqhwZeTANMqYVVcQgm0b825n0txkkb1XDDINlTrgFElDO9
NLwj0Aq6IrmALAtQPkR89EIXihYQkgPm7AgYs8PRMt+Lk9dzPmJywFB/Br9J
ySnKotWIVcDBUMfmHlqkTIwr99tTTlJYzu8JooXpN9USkLcbLEOngmqHgvPr
nLZiZgAkWGwCOqYre/Ijc4KRGLqTG/pdkx6TH+jlozJskEmTmXgDCe/THJlz
Z2hxHjsnZ6scdFgnW5p3PU9TpJ4yxirDwBpHbvvLc1yDqi+NmEOYShnEru3W
Eb4b/FxYvGtwbsHWdwJ47358gMW9LgqoRLPVYVucbIqbkLKFV194F7V3NR3l
rmXxlhRjRa/wYA8tl8s2JHdBt6zf4/whT5Rphirr5Rxm0mffLsFPqSLeb+dK
NzDSZuF/jebOSPgc+yuVKqqJV7gEJdSdmJ08YZJ/pMiNnDnmR9mSrcRr4LZt
gG9fBjJ/k/y04pkHYTd/ApC6cSVlCU2CPUMPjIKSBvOX00egBAdCEWcOqEkq
G27wVMjEpMqZiilFZYPHG5dp7pmV3jngiR4QgKr98S/zAPP4Feg9hsdl7KE1
0hgZIDKMUPobKYH64Dho2ktWPnMVMsgcbQVNgQTiX+/Dhh6otivrYtJfU6hu
dji+eoXn/dtyaLf9LSb2MkqexZudpmmahinp+E1rguX3ybuaKDIed4QwiTJL
uluPEGZ4XhrZuLuqwNKWuCG8iHshiOLvmTGkunsZvO2diPlDnFF1sVSlZ4VN
92EEhpP8Oq3r1p1ePt8f1vFT9wTCvVh/xGeOcaZBMM31ySvvi39Qid6twc88
1rV+hjGpmFTvCPKEag9I7236fYAmWe17Nw5UH5ki1I5ZH+KTNSeoXPofKM7Z
ntwuz/lH23G0EW70aW83IeXbkfbb4JsNH7RWNVTbQIhIkrCuWeKKN80eWBpP
/2jhzdfS0uA6asNJokl4Shxq/IP/vQcULnNhdtRwFH3IDGSAhJli9DCAED3g
IUBMqSYlmG7rzobkdpZrihedXj5mL9FsQYKgjdZqPhf6vLVmU7OoujwkOt0c
bsVsOc0ls3Zdv7ilJbFwQzVpYLnir0WfyBH8T3wQemTJt3+97aR/uakPRqF5
CzWtqz7aR5Zc8XO7CVW5ALRAVpZ8PLAKGk807Fu73NqI8feVF2fMpUK+1g4t
jf35RtK8TJXX/tgxJaHNxAaE5QIlNKz8FzMYPM8vzJiGsKBlao13U24jPjLs
8r8JAt/rd36Pup8oaEZANjyrhrqRHLYnq+0dsMznt9m4Ee5+wGjeMd9r3zHn
FN711ORTdhK4kGxKJ9Ug1/GvSInqG7XnILhQxmMeWnyfy6TKhgUTM7s3vUxw
NRqguo0IhAgTSBHnYMYq9O2fOQaK1zOQZhy45CTtt7VDWmaCRnDCJWtbNJkU
NciUx6XwvURetqnHcOw3DdwJ2QUupj9PIBs7SMtcTLo7akzWyNCMSGG7L5U/
G5M4tGW11AAPkqkmjLhLUR5zagrvky4bhOf8HB2na+5ZPm6PFeMZx38Y1/5N
WSLpZvUKE+gOuXPSkMgAxWz1xpBCww65cDwGY51EnWhIuC7y4xI/maMW56hL
3v59Lm1RQTGdPF0QC+xt86SAh1cRsVndXvBr0iPHQ2AXaHwXp6bOPj+OEgsa
IR1CC/F5JaGqSmpgplL0TJrjUxJCdRE+jefZr4KqL46VX8tDQh9I+GAGityr
S4aNYxd+3i2FmKh7LBjjOJpQ5S8UyJz6SqL/ndwatJ6IdJz41Cb4jvjh1aJk
vLcymEVpseyJQhYFDpyF5u/2hk7XHbCH8KQPutYUsjabLVdirdN5xR11VsbG
ybVgWnjopyhnP5Rg2ubS3lHwi3iTY0cp1LAh9/1e8lS4EnpRM2IxIc9ut8gT
d6hrGmMhWrIvL/Z8lY3jZaw/IKKdIQjcPe/5P2CPd2ZsVHCdtiZOtTVSJSlw
2xPId1RyOv3lFFBTSkpwA137SaZXPH+V9TD803fw65KLk/B2koadas5GK5Tq
STfsA8lohou870XenaUFJFJcpm1lGuVhOL0UuDzgl6V0d6cCGL8WZu/v0Pcc
/NYPeWrkiMFtKlEL/q0P0C1HE2wj8E8ySjohGVUJA0dYGRwjcX+6H5JNp7kq
1hu7AaiAB7XN3MCpFV4MyO6oWH8e2QqJfcYrZlfUTitJlD9m6/qZxabO7uZ8
aopJ6cn+tJWz9eaIvJIxJ8yfVEXENtusfNfDY/nmvv7jI6wYm5M83uotRwih
xf+uNUEpJprokiwbmVc3haGGFOKNrulvicK2OEkEHw0ebmaScN/cr6++KLCK
jEm10YQayWx4bKjjZV2mNoa5fMA08xnydUyF/YB7Yp3aAqBabfA+mcbsn3w0
6c6KBy9XS2v06P7GzEo433vILy8AefExQ+sCVpoNfLYFPC63Nwu5Lv0KEAhg
M8Ipsv/mQQoHm2XNjIJ6wPXx3IzSppIQdQoj0WNYe25UBXt51Kz3nDoVyXjZ
n/32GkQpviODeJkRDaXkH+csyUtWn0qep5O5ydri57QDNAuwbaFefUpTFw5O
OICpUXLZOWBSx0GjMhjGwu+WNq69Wo3t25L98UfxKe3P5kQaZ+bd98eIJYHJ
0v5nS3AUN/0MsjKvtrRvfX902TlHascet0iA2sN6EuVMcutZqYHawB8oQ6Ny
kYyGhXjMFkYsqcMjYbYnLct3mvSlSVZ+mEU0YIvPrT+HYm3La/XCKd6jdlSm
jBmjFwGLQyyjNZTWIR45lIb0h8sK8hkJAxNBvbqVNHXJPgDyGGRePrvRnjuc
K7eHQKA1XQ2KEGq7p5ISTybF7os5tSOZkib2d13YE8WHcK7POsLZJaE8zBQW
kYQQimVOFN/ppD5fGLnjAUkodrefTTwkdwGTnWeiLF5fh+4OlaSz9ZJszmCZ
EBDEAJZhBQ431yDU5XyKgVm+IR63G1xWo0WkIuhujB09x68TEGG8cXSPjmOm
i6GIUOf2kfcjc+e5XgCkMjf5L51WM0eQBXFqKmSckppvKLMM9WZsFoVhfef9
r7hr8gm361KfTisQPwct2dY8fFlwTrzqpU1+qLHmOc2zrCoXsFRNBzPfKdSx
tGtidC+ob4dMTHyyVgjiHXczMDzwMWKYx44QbFN2bYSH28SwVrym4TXvSsK8
eL92Fdb60JHwa1hpUn8ekdh2XEVmVlsZywDVtfCnde2HjDTp3pRHwNpf3xsB
nC+/6XUQa8nys4N0o633fv42tG5gW4kyBQbU3Ib6OHMo0nEkuOUMeq03ZHdc
0S97poNJbDtxOWQEffNmMPD3RgpoeMZfdkq3rZmvZPUhWiuewUAQZyl7MO/b
xBfEwBKmg1kICcqpA17+LUe2wABqLniMbGvEccwQluYEICFp7ZU6ccRZs7lF
PMy01EtSgDEGKGLskOWAS48j7CgTFYl4r0hv+P4/1Bobtbx8PbIXoLDixglG
uXeSC00sV2Wjm6GbO6HopwdPfdR+RhcRFVYTA4V9GrjEpH9NhB9JSaL+4a6D
vwO0dvaEsiOAq/SpT/LwIvr5S01mZ4Hi0FAV1YCPF2Rt2Op410mqfEFZDC9Q
9YWDcdGfxuteVsTwZvH/o5akFtg1o2SoYRMZA8JkuyxSCmfd/G93fasYeG3S
sLUgFkcpKvWwSVLnBHk7mci6+ZYXxsRvZpSfn3HIjaFdbSY8vDotJFTuGCVL
SSrSmy6hVnaPlgthZWvOff7WX2/VI0dhXT4Pdc8Y/T1eUIA/hczdq0e+LjZo
K8a3I9KPeGh7u4gb8EJziPGn1txsjCwet7FAX5quYr6aGl15CnyfKNgMAouC
5cjPaB6W1q4to1lX7F3NBr+2VajtEqRbMman6RloiaqH9S/SOJhJFbqKJBRG
tdX1JN8W+akoQxsakxFb1FLkB/Vn82T0ZU61W4dCnzSNphlN+tiJNSi5Zcyi
Vh2YP56S2I5PiWlZKFzpG9ajMjl2tYNXmjlvmyprJnZTdhWkLBZBaffXFvvq
w98qSBX0Tu2oAamUkMdSUAkO02no/sLQ3T0xxye30YZbRi+SaF9u7XH0YaxS
F0OvhDfrj/UHU+o7FH99afGPQ1spxED6zXyZ2KJaX1VImkJc9PwYeRQtgK1g
Fu0/eo61qRxOabf30v4kSJjahuNHWrkID7ZkEuKPok6ID8bQUn1DA6qiAVUO
jHES6/WIGn1z3aRs/ownVnL1OsCFSR2XTndNXtRpAgxQvyOIdsBfliKSgysc
944h6nxqj1iLvAQDdrThWqpCO6VVWmeS5RMSe2YcMsKiYg0SxBqNnz6KhApv
YPOHzIn1aludcXNkVdI6ldgw9UDifZl0cfbxQj/UVnKn0dRFhpWNEszU3ANT
cjTVLcn5m2FqHxUQ7fGxtOXSZ40ijWnxTHl6sWtUybshLI7ev++9j47crP3A
4fPUzdAqXPZM2T+/RwE6glFXWnSDa6h5FfkvYVQa3eYzsMi8P7Ux2fIOfCyK
QSDJ0SGzqs4kQi1m0caeZVLVvc9YmmKn5p8OE9vpg52Pyz/hNDG0pb3oQfMp
unxRV4thaS0sq+QO5ma3nWO1AajZEnfSS2wtxob1ks6n9DlZL/e2nddCKLXU
UTMeNDUDdEH+6Ec2mHyhv0qGg+9IBDzJTi0qbvJ1fysYlJhy5wL8NUJQRBCM
X1oV2f0IfYUU7Eg+uplit52d7Z3OnEZwqWaXWjpz/jq1sY0JdPHcBiFsOpAg
Ig+gnto4OUHAqa4BUO318mCgQMigjzLBq2cHRvQ0gUxgFImePJSKP07ICD+0
mGeDFffr74mZP69r7CMljH9LCRmyuXjxklxVAMOrf2VCgvZtdoCJxB0xuQ2V
uvForrzDQdjiHnT1bTDKpSWQq/Wg9PHaExVpKb7qF5ipaYTdCDRceK+oCyGX
zeXExGhT2Esoe5yR/VLbdV8ZkfzPbhF1LRW6OqcU1k0O9Mswy4z7StZiqfnD
ZfI7zUJUqZLIhuMTgSfQjZLUjn4kQ90lllrs2xl6faL0YL+1SlUCBkE0bJVN
FR/8HrwqHXsfC41sqJ2OeoPOzvM24ZGwzakFAEJ2RI5RoIYb4FSb3/Gv++eK
bpvLQuy999yjCwCiUoHfsi07Mo8bo3iieV0GTgmwTL2006JO8tw2jZ8LGGWp
vVTnHTpwB/y9qL1WvUuOFuzYrBbzmfL2vh8JyU2rP1sZYR6IuQxQz6o6BodV
vaJC4xE8y5nbt7en+g3qtJON1jvd1Sfw6OZReAHJC6Cr0oV3+nCgU+SPK2YF
XZ9GhL4rmWbZ2EpYM7PJu6MdcaWXQ0RGP709xMTun0mlQuY4c93k3QL/dy74
eacLAsgjflJSolANKZQ88t7vBFo6zSp28clxND7EYrcdyQXntyoPzvcZei2s
B1X1BOL4dJN2PZJSG1iscUqgIbal9J7IBI5mku1jRM56WMu/CdHu9Y7SJnQ1
CdkgYlCMXYsG1NIALIuhE8P7GTfKJAx0IDskr2LSDUyvTsiSrT0X+voieyDu
6CbqcJ+J89m91yJp7N+7Lh7OpjoSyuBTYI/Gx/LDc11+tKI8yKO9rHICU8eJ
C78O0Dpi2Xxk6MwEk4W/UFEVkd+/5635O48GojohF4cjg7Ke5UBVbH1qhRyx
jbOqgmmJUqf+F3Tmi4WFPNpEmukvvOQyry+e2pVIaHXxfQP59dIH4gyripBx
/e+P5p2qGKssJRWwXVNWDHHFF7QxSA4JYBITGHc1p/ivv+m6Q09JOWLLlBH3
aa7i2xBmosp7Ipyn7FEXOiXeDHMQMDSU1TaHNoK54Rbcrbl7Is1/THnNNmzb
CISlmbyauZVaObBxwOFQO+BwgCIMUWoYafv/ZBnOU6WdUxXSTxHUGBJ3BsJj
58UsVHjkXE81Xy8M4C7RL4upDW2BXo7I6FQrVMD5W8f95J7+aafiAbpNpezX
95Y4LRbS6f8coOZ8zEJDAmMK95VpvRiABgQ3EdyJY/gFlH0JQgzskFGJtGzu
t9EQWetQTb8Ge1CvAzJavhMIr8pTGwunlY4ZeZeZivTc9XejJifoBosj/dEa
iS9dem+N4TJHl9IvXG1biOudOY/xfXCPoohGmHI8J5xMSd74K+CnmlDlFQGd
ec5cjiz/SOJx8cDmx7wdbIcAZVhsw074CnoKfRShFZfem8Vf5tPegNNCPRlA
G3vsG6wdKA8H05+kBLN7R1xGnPXXT9ws6XOUcv5OBoF3FAlv3FW+OX9q8em4
dWjtFcbQaz5k1K3gluUALKn5LZIW7PoFJ7pj4Qdr9NwgIpVbHWiulY6JQTQk
UE/Jwtbhsi1JLPZLdhfDF3EsjLHSKSzwnEFyHB+xZ8UNfXqZPKZDubq+/+ZM
m8f9Tl9oQlFhTL4jLS9LrKJrbjgaUd3trK7eNT/BePF66718pf7uIOMJDujZ
wM0k6P4z4ROIXz8mpeATA32iHo2vpNbG4Jp6JMSC/ALfvAqCnCUq19ExbGIj
NPUuJ9MVIBwbX96K/7bQOy/R3xw7WZHoZABdxpnWGa/TQrtaVzN88t44YaRk
7RCrsTgTjvlHxCpDOJHzZiKDLLqhg4yHYl2b2g83b/G1Ev3GfLv0UJzveKeY
w4NbRHQyaWNockhO1w3ith26QSzLH2wNme0PJ0bfagV58YDOl1wfhf6ZbUJI
JH5GrKIUIE1J9zjK4afN1GyeOjtBIQsWaSy9Zji8Fb10rj0eXyYNjaRsoNp3
d/m7M9ve46dbD+V5uu2Mjk5+wnzAk2Tc8kLkRNAmmZ3tFCuXmphGoqKTTotI
Ms0qkBawyFEyDddje+yfj0DQiX3NYaBBnZbHKOHerN4g9ZfHqheWknS6hWV4
jelhXz8j+NFCqMrh0jhB4L11D3lGcNc2wnkA5pKoiuQh5AvhgrNuLBbjLDSH
J/tc7VdHa86BVbezLxbobD0zlMAxEZIqm8g9dbC5TIq87vI7xwXto/nB6nRK
6xqF5BU0kC2liUUZqqOyupRTuQLIsooa+Jd9+a+spxa4BoFnXMJfNb5bRKJy
KSr16dpWYgLbPjy/sKGBVjwxyU+SZt1ItwG/qTsVBUUT3nF3GLUoapX7do22
9b/cHKVzRevOUJOBOQ2He1XZEQsEKy2xT5oa1Zsg8tZgcKivmf9QiQs1J60V
9ipzn+aK7FHPHsTZqJvyzvQRajWhQ0D9bcndRSbwhzW7ZaMjJmCnYvJoEIg6
IElw5d2exWg9i7+s8hf0CpNajVHM5RqBCwi1PfNEYdvYHvm0NVANdpTeRfx9
72wk2P/p0ClxhVJK/D4FQH+LlsmdR0r+sydRhGLXis3alkV8WyqTFMLK3QtF
leSX9fYzdAi0D+5cYvC5zL96+IH285wU53bdIq0rFV5HWZjwT5IbdRZRhkgz
XjV2V4hacub6bnUetp8/ntvdKpJRLTnrBQmxlmBZae1cFZHQZkwCDLYN/oma
lUGJLQO4DtIL3DoQK7uI0wkgVfcKsZCITADJGhVvz8RiMjaw9+C3mRUYmOjD
sfe6/nmptI9WIrCp69dvu5eXxmKP9qr0k76ab5CiH2CnyObi1qV3xQJPW5Yr
s3d/kW9dVgS2xs5q1ZU8z2WiByjKxmctU4wt6FhhIyZrV3YneCAXZt9jvYEY
KknDWse5sn9czhbLFb6uLaeg3TXf09tYAgwEgKTNjX+rAJvqNhRMl9UcBu5T
fUCbCoFD4It1PHH8LClWlmKFEj7T9isR84w6GusZ2jEB6s5N4439foP2oSKI
8rUaw0u+6OPlowu9JU9ljQJF7KGJxPM+R4Mw6d1NLZDdEbENl6EGR02gRWY9
LSmjjLNmRsIQW1eFkxD4LXfmmqma5qeD2GZCyG3obew4zIvMqKdFb4HoplsM
fnF/fuX+7HPTLmUFAlhCNU0+PENCEsNwcrt7hy9RMm2XI8BlbTyTXf6FyJ03
SJTvbkhZWqBMa1TWTHDxHLysgDxyknYB6sGgs7KjrtULjoUAwK1gI1WFAfl3
g+knnZozxsAsJw7FWB77zGrlt0J6/JFtuQTq64MoOlAXBMpwNiuLy9OKIxl6
qqLDhBxf5F18nTNk5MMTlQmQXn+dI4x1JQMNvlYN7l+KEHh8SKijxMR5KSNg
LwtRMyjUjBjV6ZqrLOWT21OT4sJg2u4nGmpVLlJjFrCFVB9+oOyTd75zAvKh
2w3B+ZN/DnWWexZiBDxN4wmLyacYzHxiz76kMpu1fzwVvAQlUAkH/rOGBbFo
5DnS2HJgkoKBNQ3fOwL6lnegHGLDyplI+/qgtnn90UZMWkwGZL9Bhnz6mpQR
XP4+EWvHifwM6EL0hsmKF5r2Kw88/da5gSVroZE4UBR03DSu6SJBLuMvcWbo
nFSXL3Lt69yAf4rfcwYkVTGKcdjhDYF/z7mlU8iY3xRpSUpRfZo2D1BnlBFj
rrA7gtAuM7fG76yWKvf7+n1B1uFAUIHOcCPj0kg37kkOpHrmXQaFQcnP5jCw
3Wt6i+/Lhh8x0yMqy6GvokWcUsHQHC8fc0vdOy+1tVSwqrA7w9ZBv/uxlA08
8H4nWYqd6Ru52dBSgjDMW5EK7ixwzY9dI73kyzMhE7DmiBL3w67zgqKfYAkN
Am1zV4HikIvasMDfyCImOsWKutozoVkevWDYnxVGSOQNAB7CrgaBd8GLZ6xk
2RXav+tr5XIk6AZdPrvGr0eXYW5GTj6Wvgs6sCvmpmksgRFKvhDKmDlmY0x/
Eu1EgXCDKWKwaLEqKAH+h72oS554d+JvK4b0evlRnaUM/d7PErPicnlm4Yfq
Hzf8hywr7YreXXzfjWKCbn95iYWZUZ1XBbdwYgfwpbJF/qcYd2CfRya0wJHc
y2fI068AZFXFq8ig3iXpNnt60LeoOMwxG5V8t2FbrhrDYhr9FV+fFwUjFjKd
HCxpNGgFAAsfSQrJc3YWDf6kxZVOdfIuKrymepmW7ZfGCoecUBfTmJ4/srJV
6cwUDSNG0k7v/UWnzWooeAn/4QDvJ4FmgbsXLbvKWme8VxXeX9TCP+ywRMUJ
Vjj9YTPtsRsKAWBSpjUHt+5lNLk2+hWboDPub3i9EkmiHcbBafQruD5jEy3o
eCjTAJbw8J9bsM8o9YkuZjot6qp8mcoji0SxqjHUzZxaVb6KqL1puAxpJSCZ
rMSv+5jCvQSpN9wvCPzeNTlIVUaFZ6Ed9JPdYMBwud5H32R0lXjvoodQ3Jeg
jjoI8Pi2cDGQeg1qHtLeUV2H0ErIUK/m/ftvb0Q/JSw2j1Nc9AlzOqQGqgZj
iiJTBYx8pviVghzNyrTh/a3zCQS20IRNXWpFcz1OBgTzJgwky8g2cptpNO7f
ixVFwrzEiVuLa4B1O0yArBNByk8MOPaUO7u+7TmDO9hefRfUauNhRe7hy6hy
CJdcEeXP/KN10Fbo5AzwFsLmLZoHxaaLu98vYrzc5Mf1h/Tl2mgKqUB+N7gk
pNmrlTH1Zu6XPhNOKRBlmHEZPB72BQTM/DZfvoGynDEZ8L75M/l+od6RbrCC
ftu2B3WeMjH6nY3YpvJBE+5axxcW+NuVDgV0PyHn0nIf6+6kNVxIMbeVucc7
DvkGSY40HhuBXYwZ8xnmHxejphtEfusKlmrHySsnxRnBnAYL++9SWMXCC/Os
+XkgTRouUgerldNMq7nFRNZ1RcUCGo/ZcNE7MuxhXeqzR0YgMTqDSiI9O6s1
MMHjm8AQXWZ4+PxAJxNPxPB3sLfUWfvRSCdw3WbsjVedkDyGtm7cvj40QEPr
DTNw03Vk2Vfpp1XTSEei27To+7UnkuGM0XcWHKgLhKx5qoYthBKnhPh77ZbB
s0AMp5CP/7sg7WSDj8BmIFtfmKG5tEj4U1CcsLM+RqpJIO6zqEqw+IVqZdYB
VPDxbFaRySGhQQeKeMbLZhQkRS6J7xgruvNQt67LLai0Dg5F83N5JpI7khte
CHF6bPMgV3ihXuQ40h97+Qd8Ej/Dt/OrtCd1KKNw7hJhJ3JzaFWqnkIM6SsP
B4mf28m66M7gYdcXUWBMDdSBAx7M7MqWKF1R/LK+sA067G/UHbrRoAVk7dTe
RPG8LUr2i0O0CxcCzTdtWCcHMNZsmTKADZKA6+KU00uYn4baRt8YcD6rGLrU
iS3bfyfRPGfXk5SfCaaUDmpy9JFp6+gDR/FmWowDLlA6IL2QHiIBJbSIwg5j
V+2W3wa1K83OgcIoeyr/I1Ea8uc9+4wSgLLTTnSwsCqA1gvfdlJ9Mv6f7Kvt
vcNNMDHJ54C3TvPmiphXR1A+PDj9zb53RgWMNzu0fyNDcA35livcuugC6dfF
32pIVzKRY5EyUYZbOOpNUDYKH9tfBSunP1SliRGmpP8fGlE6DMC8llKVFWH5
+hKFy7eFsW3YfaWaWBdIrTheAMfmrgVIJuJZ0NbLk6FmU0SJ3KuPybGGJJo5
mV0Nu4q34Sq2GbM07CgzjndsyfWHplourLDxdB1y3N7t/BbgExoRcUlFDXTc
K9/lH+a7PS+ce/4Zwot2rrEv6B5RGjf9vXLrDxcdltNQ0GHRRTHqKKGn3Xip
JQH1XJI02ktrN6yUPbGvfvzCzS8/mXESscGvRsaO6/sfhm6KJaRhrDC6wVwc
sSc6HVutfEY/GlyNf0Hd4QWQNmS6KePWcXBpgIxFhoriGTNwuoOyH4g1ugfY
bNJVap+SUDlg6oXe11tq4LoubH+0m66d6ajZJrPwRuRYrZ/+JXAogUZ5tvie
LfcAabeVwfooQ2Uf5xyibiCS16VCGJNuhQQ6rwnvqdV0O86h/16JTtmFodiT
8xDlaa/U4R23z4vVlURywBA5Jyw+WlndDHkUNF7JLKxE2VK/yTooIVg2yiMu
CCNmClSDbFhZdAy+nKslKnb9uoOKdp4khWCL1bPm+0HfhOXn4BgRdllO0CT5
S8UGFGS83RnSFuzrjHYQCTtaGjTtTUfqA/wjvmBSXhLdHmQh/UscE7QZR8SE
NfnUIgaYL4XV+eJHrXZhguyEbjHXq96QUcRqfalcMC91trsLg1BTfcJ/zteD
et3CHE3XImja8/nCnKIM/YZJ1AHSbqd6I7si/7hT93UNAMeSuHy7uepdV/S3
TmYJi+PPJUihnUsBzkWwen4YeyHff+sjMClAgSdsqnpxE7ejOE6gDmyNkwzx
gpLABsT9tcF36osrrTmU0EmX2LEh+TCkgDj1/Hx/Uo3OIshDE8vxmBU8Gg/T
hL/mc9/FGtxaQsWCY7jl+ABBgTshTJrdPsuZJunkygZYyEhGUv3D8EUtddsR
d3cbFeOVx4Q1c60AuKQ+rhXBvBSRlrtoYNp//CesrZPNJnkK0ooIMI+jDuaB
JtEIu73NxpMSp87e8U4RSlP9r/4XX2QBlP3szSXvKGFzE8KwUcCmVjOkWsVp
H1lUteSpZdy7ojAV8mjltiMDM2ozy1On/qIpY/2bjrlP39VIYNFsExbQ99gB
3U0n4Z+5BYnUJiSdC/K9XOUGnDPiZppZN50QAEw+BE6jPonbSc5RNvzvphqc
Mtr42YKL/pO0SZOZP1Iy+qy9D0Xx6R2jGz2y056rkwECjvExxwaHzoabgFqX
ARTiWDuBN+17vTm3WHLhiiSQDAw6afdYAqTB2M/XFXDebROXkDxZ4MB/sxWp
X2JbglcCMfNwaaYRUlzwbrnBLWfXqwiTvKB3gfYgSzHf52YhYCdJX6FsX6LF
ch5L2lvMnqetJT+uJ8hHAiMMCq0S5TBoPcPosMnp7gKUzL/jzssXcw8zx+/j
gVR6KZBf+grYcDSMfFplQIXEiCDpEKpi6Rz3begiFusrgYVJSOOu8J6pbeN1
E1iaWWLtDhG7+IMTckGAeV6SPdxZUph0NjDxouDHGxOZeEQmPz5G/Aw529qk
jLicjvqORdqpHmVp9U3aqxVbKlk4WEh3KErj0gUXqkPvU9wafYr8B1zrIVV8
TmFPTRGSeElFj0wWA+fROeaNHFCBa4nfkEw17Ox3VwFhQR5jMOnedMuYTd5e
7xfHYNnBDY58WDdLPyByqjHzw1Z/BQeaIOIyXLqmokuVo2A+1BiA7q+2bPJP
zwbEJrLINB0q6CxA/AQfMt/QFekhylGh4MGzYvH7zQ7Z+tscOJPckQmHrxZU
ctuHI44XvzhucdKQ3WD2pBYz16PrWtm16LvrcPsMSZM0NeCfryt9ZZ9RDKnd
hL9Hsq3PoV4TYTJf78IPzMR5PdU5EzXGBxlIjPcqF+gvtTuQSxVfOWAdplcH
Rz0K0r6gKih0Wx2uFoLG/PmBIipYBDLTvVbRhkA6sCgmSbUqhIKJD4WM6l/u
Sc25nefvMI8mNuZ6J5NvGDvABGWWoFmtL8hUbRTH41mch827blqK97JOG7YF
WpV5X/huj0EWZbrfxGUz2bL4X8EcCjaPneTXninRR3zd6ggM9JnCrIIOb6Ki
KUR50Ztaw4+bNZFU0c0fo+RYGrqwNq6naPcTfRS8RvNT7cWmGjcz2Wt+Tyb/
12ymASN6fYlGoLohavykbnqJwT0qd2NWdzUO0TP8niTObpnpvthOnDDSMRLQ
7i1LPW1lcICvL+aCokzZ/5eXo27z9BFIuSfpKTpOQrgxiXeykebp04R1vYF0
gFwGQDUZ2meysxUUQw4i1bcfPY6qP+bZwMRjlHtAjj3Gx9slm9faYL4A+0Sl
ie8ptg6ROGuXB4S1sCKK6vypO+3trjfxEmyS8PGMqmH1UDAZFoNVxiX8PUlk
tQHieLq1VtdHTSNLuza9d/l4gKCen26UTrclo70/KGFC1ej/S/Ih4Ro4yyJQ
URjeoY6B9CCuBEk361M6B3Hxuyw9jF06SxDslxvprGMrwfXKTOjjCadJZOen
q/77pl7stLUicJS3yJrRTbxqgQ3hJ0O/eDs5ahrlhr/ALlU3MALUr0xrPe7m
1yoqSfsAFgQreMM34+1cLXC5lg0LjJWHMATg15JXfp8tIzYmcicKVLwmH+IB
OBl1LoG9K/jJZx5gL2+eai9zmITELETTan6JmIwRHXIYjqeXkxXkD44yuWiI
h0uUgWY94aKAxTx2C6cHGtQmKqwNQDkDz7gUjXPNrxTsj3ErGEb/ZA0CYIlq
N7qh5vw4FDzWeiQ7yV8v9YaShOT7rWhMxbeNicQaCXzNXJjVuT0+7/ngWtUn
ghxXWEVFVNkE2RlaRbOhh6zzKH9MxCq8MN33IctYwOxH7AaiksU37W64Yc7R
Hu6MzyKsb2Epn9BfG6n5WapTKrpYU1ou38ATXRlXhAJu/pDjRQ5qFORZE8i5
Fa2iMq/YlDljlqvWTItzLsaZuww85chKFeFmhxPHx7Xyu+eie2/QieXlMiKH
U8UZECjn8lBtr/r8qoNLrD6kPO5Vn/pgBYYeRzntsd/Xsw+b+oDO+pUM8T73
+WusFngN8l0ofGUdn2u3eM3TtNc+FfI1OQPlUQG2v0Ev5IxnKhiNFyAc2RD8
E8rkJNHWthBErgyHdB4IXDerLeY6lHac6xZ2w2atWIantWPefNSkro6LiFmY
hH0Qp8f4oUeCLppJw3Kv8dYluBhuhe1ZWZFWWbPXmouC3yLCoCTdaM7j6RRU
VHLJqQ9u8BUfwsFdpCW5Eoun94WE4f5tqNlgWl/bvAvk+aFdy0LLUwyMNMmA
gWi0Iha229EeKAF4DlD9D3/Uoyv4IQ5a8qJ+WSMwtvd6YtkxcY3lNcKkj/V7
3f2Bz9ZmVz/g4eahwQ8C+F9xuYHKUCotJjBXF1CfwH3sXEa20hdPJXdqBg53
+qZ5qLZZIv58W9zqe2bi/eOzj8SGRIblFYW+UVrt6BixUGvT8xlfUFEAFqNr
/jKtu7Ez/60toT7UTgEMzmyUt75k6kxuVm2xGMEDDCXdx+BeSknFp4aXiICB
ZklGvQ1x+des59mczNPT1aib/NOyyTUtG8VyUVTfC54U88wM8slcHskWD0PW
IlTe6KhHKwU+A9SdUCbRHzEJRHl4EOJQT+pdiBJwpyLA7HXoLDiry8zb64qS
BlNBAwlg/GcIrRbyAccIvd3T1vBU8mmDwEnh5vV83VNO+VkWhx3n7mLwJF2K
UFuTDD2r49AYO+bxKxw9YmGt3SPQjgl/c06uFJvDH1J9Vxm0+RqIUUO0Em95
/3d0XCU50rRuti6hOONBTlxE4ziSceDGAMM0UUUryh9AC2nALHCBCvvFqiR+
ORZu9fHkyiLX0RXoCczt3FXyIjO1clHLIpguetqkNcaU9lKJ+l5bBYXujrf0
BE0/P9ifIu0m53USl9fo9FspZayqx/F9qC/vz73kfWIrkzV6yTEKzbmBXXAs
Met/8NNfAMIYgmiJlE3akNdFS0FSXU5mH5YxKpzaVoFwZUGmdM3kBW1s25Ft
gIbzi2LEXyINrJrDE+1ZIcVjVACAY7N2zt7uga/XLIxB6iHkxd/hJiGpO+ta
jlwxL4T2xxe810waJGR87u1s/78OYtzAhc01I7gebvHjsc+fOsyQMIu6GXzk
UX4WzJp7zKXsTlrflswmJr6jw992NHFA4REo5znRXwt6zvESLBFTMQHFZazp
M8FY8DIkqGBnCLwxTYce3qaQRNVbfmaqixoG5KyjUQ9OQRX804iRnreBXjGL
zfYT/q+NoKiWA9+OuLN15yH3bwL8H0tDZp4JGRhwphMG/LZ3CpjgIhUdasjt
auOB97O16WUCJDXlkruTY70hfJnp5xn7MznQsVPIK0H+VmKkKXqvFLUESUuQ
9J9dgmL57tXozDKTEqOoZ7rUKXBF+i3wsPjrKkLtx/FDpmlEv+zop5kNHJ7M
TI5+uhab28v1qRX1TaHAeT4ZH1OtVfuLkJq8M3gxuQxG1y3j11qKmZfIH+Zn
vqVSosmrB3NOsv77sTBBSoSltGMNiNz6io98kzopXbVbkiQn1jSWqIpJWotx
uYXVALvPvngRIxRU7HN2nK701/9qPOZm+QtUlqZAxsGju5ZzEgG9Uaus/Ztg
RQlqvv59YMnUm7OIEmcBsgD5aTlwJhO7RPd6z3QbyOz8ceZ79z1HJ5v13aNP
C6wFtEjQYmvxrdeVGt3riX8AM3gYEeztz3MLLOOqYMnsAgV0LTPb8TSY+WEr
0QutDx4SKSG3PSxtcwFTeVaAvdEViiYOWZbNuYcbRSZL8MJdF2IALlzo8vWq
HMS+u+4aZZUl2jRWdAdLiTFWUzB+yGvYawO1q5wS2pAHI7CSYas1TCNfOHaE
TBYBM0Ye3axdrWx2m2ZRWUe3wzLrdcorP/d9Jq7+1fKMPd5Qd4YjSdZwnKYz
LfG+kPZbbLQI0c4IAW9mJIbAJSuhrWq4jYVXD9quQIr5YkPvNxpqQ+Ojdh7X
Di7f6HuRNJtnTKMC1YWh5d0NyqJ3djoActs7V2ZYJzxr1n6r5lCojI5uEGcc
Hc0xZywt+e0inRby6hKQtd54DxWSxl0DoxHrBInUzZQjsRXu9qyIXzBe/0HV
/CBNMYn+S/qwkA3lf4fcjbT90+QKUc/MjP6fdX3/ud97/aH6i1XYjmEr/8RW
DJeK1FXjbJ2m26GoC09rTeOnm+wm0BHLgmt8j2subkq/Myp1NSEXi/x+8LL3
7V3x2sQY3/wTTZf5DIyZAQeUeFQ56h5+0b6+WBHBGv7jWwyorfItQTR1ucno
Qhrlmg5pSVxbJ/zHDR5+aofxE1A9ocRdrk5yVn+wALlPgtyMc4wxlzSgR6rF
WvVR5eBeAUoERbuqxIx9y1t6ERacKxSx3pTy0xXzOhfkfmAnYeGkmoKnDzMu
9o8+pGlxGC30jt12GAjyUyYltOPuUrEYfiWhOcyFI1RMPKgTgRv3zGfQUJtU
US1UKf6i7T9Mn6TQHLjjNwwIQYo973yw7FcG9yXAW24ViZ4swv/RinUaSaXg
wzNCoIHvsg+rtDnNYk+C+wxP7BTWddmIru4cEXSLPo1NF5YjKWdZ5+v6k4jL
+EYh0+WN5aq5LBqhEGy6j7/Pzb7z6CYvDZmeYhvVvQ0+s0WXvb9H4pdAtWF1
bf/+S60bSP/ssGzJ92iussHo20CVGESSOGEd4lWtz3wslcBK9VXcvzb7rTpI
kUKYVMLMXeOlHAMcghkwQIrN8oVxcSgRNqSAsaNJPNK7QNrZtsXxlYLWsFr5
rxLHEiwAEccSRJ88CeQeGDvHkd6HTvEMWI1S4cTaFphkCAV1YgRc7f1gwScF
/fbb6/BPcvUhdYGlZ4O5hKNmzQ+tIc470lUW2UH8j4MaUZ3ZTxdzS3Y5vOv6
o4/YLbWmebMSl1jCAF6BPnAq34QZ8Aqez8m/tjH6I4nQlEd2Mgs2/7kq4cGh
bk5LlzhOyv31tNDEvagxY0zXlS/FAnJzTgIXXp9ZPpBsz1GMVsNhkemZwaBk
HizB5NpcwNoy7QYSjn1DK9RkDaMft+WMJXRG1l/hLaSbAJyqlXHq8RhnrEpI
M8rHkpctdj2cgxQ8uY8dDp8M2+LpfHC+I7SnP+hZpemPNPi0OrJJTeRm2cfL
KQzxHL0g7ouGTu3hcyQjwdLW5Tx5hvrFvsaTuPtuCPulLYTIpUgT4XlxAeKY
j+Q8NM7TtphTtW67tViTEy/2j+GmYr6rHII6YY6gqGnRnIZX5S1Gfj5nr9+B
cXG0WkGElpgCGjr9GuZ1rOqEQwvl11GM87pzhamh46HMmziDCumBuFeW8El3
NLy0LjlEdhfeTVrkJm8oYFR4tCcYt2QsHdOyZ+5VMhLawqD57/fHB6OC7mi8
lKhGuzRH9iih2lDShKmbJUuy3cQMmYgsqvtPHOVYMQfGFiV9cycfMRVjjzys
dQEyb1v6faIfiinMSGRnQdfsbe/sVvmHbRz0z15DQ7HX1fxA3FBWirAS9eI2
+ho4oTSR2jEkfiLwynvJW1f6gQs6uFPF9xbgqP40GGrha3fpzUcKV4y9Vv4X
BbyyMfrIpiSIl4+0fxCxxfW3ID0bk+gV+mS+ikq/ipY8t2ELeFlRhont3gU8
j5jdjyr/07HNG3Qh7lu9IzbPMIthWFQw2Mu40dFOvce9DvEOXWfMfxUeTHht
5XUODfgUPZxHpSfuFxL5v3WoHo7rg81yStb/yBne6xYysqemLTy9q9xMLbUa
6lYgm0oVVtdHUJ1LstgIah1I4lC4vMu/Tgt0rXNqttRPVdtkHv03TF0zUFIz
7J+KI0NQs+okaeJSChhNNUlZrMZYq4z9/xOe8tador5bwaHtiE4yw9sLBB6d
QvrNsdP+nj/O/C/ifWuvVfR9bYfBk+h8xgik2SLNhrxDt2Tegy2k2C6ffyDu
QP3e9gYHKGfGMjHohnUoqNfZYI+zW2++3QXWYt3fKEzHpu+8AvxQ7ubPgpAW
T/3uXKKxIGwzg15fbkzEwW7wI9XkfQHZAeFJM4I/yxeP2JG6Ck89Y5acDPmr
j23sACo3n3UB2LiOkiHryWzC6wD5pLjp2N8M1UkOugws5zQ2Qr/U4toqgyEh
wHnLPEruo7vKUKqMBkxVjmkcQeI9yEILPZ0/q0KqPYYW3Ec5G2X/OYmdFhcU
Opi/85ReHprb7u4gZlBPCA2sxBdMa87uzi4vbFh+o3k2cP0P+LKyuQ+p6rqH
/rUyNaJ0b98H41goi8uumckFWPZIgVXtldA2KKntMrVuVKR9A5GofNFYMuIc
54HiufDzshu74Tt/xcBG5B9S+b4044moi12TDWkdJXwyUW3FUO1IvpDFaURe
6bFUbmtvsm4jwJbgQNS8t5zWd8TEGeyMkIt/hr9vawymfA6d5FLwugsV+z5O
rS41t0lmez/OLStPxi27vfw61SweE+lJC/4st+JgyYt2b1NGNcpyf7U2ndDb
HimaIbFoDg3Wgpz1piljW2h8tEL1KcSBKV+N+46SkSaj+dnIglNmkTcdwNV9
KKtR+4U4BsmWe+IS7HusootsH2d8y7Pku+4g5zMEKrYi92FW+meJCsFAsHAH
z0oNagBJP+SJK0wWrwymqwLRUtILcuZiuBcS+sn3VfA7VArRJDm91XM7eoI6
AyKd05+nIEPB75MlH0vrdmJD8ax/uEnw63JQGEAUPG9Y19ZTapm7F8Yoedir
inISDPXnFiNQV5w3qCBjPaG+1ggTcYO0kHn5Bq/n03w42Gs0G+44zNO/Uyqy
cdogPm1cP2SYjl/OpdTdRmUoY/WMNap93o3BDQKkmUKKB4+QXYQ1iI1AcCfq
vi8TOmqHS5TBgRyv+6iEm2WEXWQNGzhXjL7XwbY98IeTfIlIghFKq8b3IU0u
TUKowtQOpylXL7V+c22kphyma9lxx4K5bRUbw+vtX+KKgDeFeQ49zqoL/RGh
65eJvaKkV3vKFz9Qh97wOdQE/azeaFzmHJo9iuC/hr1l/oKRbLc4yJzlDz1b
G9x78iw81Kg8tx7QIvqTuR/KMAWBJZe6htvu0k9WTBwwkb78L3CPko46stNi
/yzhgpEeX2+zak0nQZagFxgl4OuO6u1SLB0/r1xlinI8PQWqiY4Gt9prH8sm
dOm9zJiUbmynjtlEgujSWwtJilmcY/XJ38QBt4Eyd5a7wtMsWWIpvleoaY03
nX62NW2E4jR0bomVAK4mMYvvEsy5TywkNP041TrL3CgNw6g6n+WJcD96nU8y
gcMVLAKqyd1k6ioTnARrEvLHVEtv/5a2Re8954kNwyHfp7aCWNijBSdSRZxp
VkWBOG2/uifwAnNlCGDjgdGMv6rDn1PMrzU13Y6c9TIm9ol0n6lO1MMOys1w
P9y8HBXjp6ToJYlWpSqay45kXxazhdiui9VFFiXOi62AA+dHRZQiyofxr562
pxoyGytEAXLmAe2waFskgxoimtQNMrnARLa7nLwFSLQt3QT2jI7xq8nAGd3T
zWEmB0/SSvNhVRBac645d+ey1gi2d7XsyNLfVCELjeKVzs82kcx9CCwzMMYi
aJbLEw==

`pragma protect end_protected
