// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NgDDpZoTPuZZyi4HH7h5zH6vVoXgktwKnlc9Qji57q9WV/+aURUMEorspjWJ
VZUINpFVSI9nGCfPMvmQS8r4HFBmIQQFojD0XF4GsY49dgkGc+P4UbPfdIVx
QZRJEMkat6kZ/5HMBDAi2OY6PN3kewa7rbUpH6LrdRyNB3ySKY2IGiz2w1F6
UixxmO3cQYrLC9TEtY/Rjf5D+kjGGTRYYO3yx5xG4JTq29FsB7pbz3vamU3r
8B49ZheaCJ4QnUFDQJBX86Two3VB78yIjtifTrWj/11NdEyfo9/1oIcY+tsg
4CWM1EVZUXq0LPl195vwA1ocOBZI2Nj7oF9aZhXirQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kFeWHUZcFAGU2ROOscmPCu/bDIGtU4a70QaxgL32D7h1dRhbK6OmKKrweyLw
XRnz+cdUiAKsvEKaHuFO9WWa/cQLy085g8F0ern7FDZuCA9k+DFc0Y1eVcNv
U4afHCqRTHtLEmB86IWxkP+53dSDM1cUOKDgQsLOKX+RqTKwbyGpYSZYAg3r
krHWcddGxsSHEdjhwMVapGxOfT9bBnJ5/6zjbej59MzzjuctOhcVXE7eKHT/
k6ziwljmG7Vwr8LPpoj6Wc5mXylQ3dHap1kBW+NrNM1yF9KGlkr8jXjzy+aw
MXraUu5FFO9qx/MKxgG8IzvHjl05yLiW9VmuvlynjA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ejqx8Y+T0RrLMbHP1YKknWmVfyGlZ80BN6Zqepbqr3E1CASnFctqXwBcrLbF
PKGQUVeiVckT8BvksycQLrl0FM/WK9GUoRFDaksYaFrjjSL4Ds2CDcyqyabi
7+V0V5VTdj2frKN22ZFsuoEk8qpJxo8f42EypyVckkYSr69v9sfz12D9HHTP
vpuEfPGMwwSYQoQXGzQtxf9XtQU7964z4xGqeya8QOnkk37NRqISZ0qFlgE+
dp9rMoJAbefQ7eWVeE1ycCgsi0+dVeZk1ZDNK70vyzfjyvN6D+E6f3MFh69n
vzBrzBOr4ecTWzVVk0q/0sSzXgonT7AcIXuw8+ghXg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YGt6886B6QQ2kszC3I5YoN8QqIYGw1gJXPD2XGyxpadt0IGPvvvjYErj4xn5
Ce4cqaOt4GMGGvM30K2CG+lzvpGnXdtas90gTae0+KJlgmtM222O11cEUEUQ
TmcTJQ1oPMVCp+B/Id5BYG7Jev8vOHgDgvoAfEFZ2fob9WFxcjU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yH84hz1TS1NSHfAuUYpEOeU8rWGS6dQQDBUSZDes4Ms1e4tgWSjlbjfwh2/w
rzknpvAiZeCShBf6PJ1Fxhmmlld4FxS2QDUz0sIgItpyj2RvlAdU3XtjBNy6
YnFhomulsAMAJb/2dO64mqb0PteoSQ9ov4wqqWkWRe6JTUCreeQGUOpYPdgn
B3KrAMTa4QniyaXWBM/oEnKrdcL/7r1SKktOrDFsEeiwW3CKVIus0q+Sh5Cb
1VLij4PR9N30RZjwDMHE1uALKUH/mmaF/+69Ahj5GJ39Q949xXIIKMQujSX9
DgWhUqY0NGSvKA+0fNQMTIsIdJgd48KUEl/7WO5+Tw+bxvq8uOTxjWst5vHX
pA1Cja72ORaNSc8t36thCup0HwnkFqvhlONYWasJGvYlLAgFQ4qLmIHb6qJN
ygFK6PKn9mdh6Uh7l+XPhxRl7Ckpk7EwhyOzM7hE/xHHjDa/w0z1JdDNhiiW
4hiqoU4kExUNlzrGfc9ZWeN7intUWj3g


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sFJGmZMo8fdYBaW53xjA5T4q+3fTB/TbpObFm84l9P5KOha1zLuKpV00NG6n
KDdvVXZ4KFpEYqSjiX+bBuKV8s5rQObeGoWlKdKD5E1OhAHWfp4IEfzHBGhC
yt/Xv3MgYCNloEU816sBkxg3pO8ttO8Ni36e7M1FOnuaK0Vq+YU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aRCDHiQrfDbHct6VJlkH+ru1O8EBb7ZLTHJE87RztTbvQp9RPu3oGIF5wyUg
ZBJbxjrmdd8x388UegKOS7RQllcpE/md5blmVyDodExnP8I8AiU6i9HsrMAZ
SluiuAWWOhZADADARcbBYxD9EU3SL9KWQ4VJKWsb3nWjQ+fvlFM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2576)
`pragma protect data_block
EBZabHXnMueoupHVQ8xyMXdU0sc8Mk+qH38nGmcne9ewr36v6+cM4L8FBJQH
LTQPezdGAbplGPaxOv/U22R5dVbonWKER9o3gCj5wzKsOjaX/eHOK9RqPJNZ
p367Uq5FjbMUfhjz0EvqhTn7eASTrQfJfsLXidvZc9Q9a5sHZxfhtLpJC63V
uqTVug5NPGZtd/u4ybAKOTHGkMu4N4yK/P3SnrTV4fTiV9yu8QPYBLKoQ+9K
l0xPXf97cIOBGFXkD1nSRdFwoVAfy19JTzjEBSLhMuxWtanRpnEtImErf/Qs
iowxzaAm17l0fMj8BzhthzZhODBxfBjY5xMu+dWOOiWKA1fgBR+b9LC/BJQl
WhAfzrL1JNjOhiDFsUJH67ZbjH9e1LPiWEdeiGFNzoyPLEKmvPtrgk+MC47H
IKcJqYYA6ckaPSbFPYyKTfobcib4Fbd0ETMUyxgaPSSB/Xk/4eDFARbwljeI
UhKzanQddN+4lrbbt8Mu1m1mbe57QvDiuYbFW3y/o0jD62z/ppoth/bvxxj0
g3iyQXgO9YgrjXOWSKpGCbDyjVdt6eug8g7jIIS7vVV683cC4X9NRxJFgkck
d1aK3jiWUP+mVH6K+mKvtuOdRPieQXmnPXwOPifRV8aJcEmBLy3FzJaPWAcl
ioVya57Y2zr0AKY1hY2fs1ynAV9oH/huHmAuUghglYhZUwYmo6ec6+ewgmRl
1Ndc7UW/VBBUkbCUhODQjhj5UTkZPX3adx5uaQ0K/GLGIilmtrQqpcxQU7JB
akYmtzEPUQM5UqdjvoZ0yfg/hc33RdcZ+8TGF8x4GCDN3tbZ/qD7yAomgTrc
Ny9jzTDX6VY60UfHNf8bKgdjAnt+yB7gIvxk155cUVev1QLWJVy3AlMyUrc3
Sn1qRGaPxzPsrdtrB7uPz77IAdt1gXkDFoXsHrQItif20DqtiFo7y73v8YNe
CUaE2HK9d/GNqFSt4TBK5FQ4zY6NaoU3BY1lqMOOrKisVLRbcCFVOFKcvb4I
+//LLMRKZ0omE9n5BfvWun1kbOUWmPkW4j96vYrxSZLFdHfZc8FadWZAobF7
OSv1Pvs/2Uk0/8kmOHO2EqHTf3pljsoWDLWwaE1ollVHRkT5m2OL9KztQyVW
Q5xmPyCHO4/PQBFivqnLva7uccr5UbZ7og8yyGycKd9ebSpzniIDETWMTtfO
HFYjGpWiBlSk2sY5Onjj5hxqKIPX/6TXsNlCC1ddsd39lE8isqHeer7vC7cq
LVH4ijwEsMZQVBQPneeqTLAFzJEtfg9B1CGr8YotYTSQaVO9zly4cZrLUkRG
zLEkw6+Oz/nx3coXUARlyNDIpV5GMN/72wO2jeAV6bPPXS4GHUEj8ePOb2ZX
5N4hJIOI3jTwzd+re8tTRIvZFpxRxzNqTgItTdGNtodci0TSIfxBi8qbmI1r
0VmRawgleCKZFIyQxYkfiQuSdslEr/q/F1Gh8PjxqZOJ4EIY3Aaefjs9CPPF
01iWHUUX+z5bH6ZQHe+njxKehcNgZYnubfJzUbcS0p0RFFI4Wa+XosTpTKiS
ckXrhrHtLz5Y2VCXJuzdvzPtZvNZ4N00kNX90Bq1uQyUKfvviqMvAOGhqXez
rB1zWo8Dx9ZwhripPNJCpLWYTnqUFV06NIk+sX/lMr1DuSc6eIiacBuN4nHv
2Gf5cFhmPMeF6GxkC5elBIQPnr+mYtQUfQVMjHXm8cM5Ty6B9qFcYIfOPJ/0
R0EbYHJ/xEHyNIGxKdto0J3Xp0x8n2tiZ845oV9VY5efJ0B/qVav+TInjTUm
ZCAvtu9PVJswoHybEDCUVQ9lG219Dmpv3QAxVHsYifYdGQU830oSdzFP5U2F
xexq7sP0V4ucfmRCVokQ9cMBaZaKqPvai9hUB2xDe5vNnSUv52Y6ry4xqzF9
UGImS0vsQwtkROi+dGpCtVNLVt8o6FuPuHw9y1T+3wH64d2Cp1TTzSqQEMvH
ApFyZocHcH522tXih0WD2hTOKx3IP67C9dfEc2IOUCiAckZo+BrgMFxP3bwF
ElZ6KAeDTvEsKrxKi5MV6Upu4Tu4qduKYuRb1ry/mNKXL13snMGsbL5znOUJ
vAVJ7TyVAsFv/M/uY5hnW7WxWp0SGx1RTYq4cOSPNHFE1DwVsm8A7OL7z6J4
evMuMT4P5ZVGlzfsqfZfFDcxKOoUp/o4MxtJ/XTGuFMXQSGuxLIykGCj4bG7
73l3bYRQqlY+7cEyQkWFDZoTx6BltKsJ5K4PTJMSs1Y2Ew+mpxlHVw/0HAnJ
mJ7yZ/uEg6bdueczj7MMB0oJdnBWUuWLEhBhiyzfyqOwgvQdwr3i8kDzkrj3
YBOGR/SuZaoDtLaZCQSNRYKhVF09eTf60M1tO6e9nfwSLm50nm/OgT5RNLKM
3FzrOe9nSDoXCNajvOZbTmKnrViuK9szXCEyD1Xo9/JZp+GUUEJxQh3/BK/U
GoUXj9mq5C0KCEacWnVmrAgWlbPMaSPQO+p31f9TKWcAwodumvIer3H+D6JZ
mifWtsbmSMpVkkaD/aV/RW2cAPxqiHjKRlD+DBu1nbS9mulqNeksHXX1rVlD
YZOaEQboSEozt2A4epWmlhwyQI71eYsaUU44AIA8HRtGK3oi2lt60IIpnFMP
werOjLtOp2xBLgcBNx8Z/py6cIHslYj5D4X90QG6wxPay/EZgaCARs0eymcC
NARHqtPUrAClx+R8HttEVdq/85r6bSqcF4ifRDhrCE5BEQTk9ehoj3WURti6
EQsj220o7pjOdcVJ9sapaVf3GKrHEJ6P44x903MfkX8i+uQNcfGoHXZVDkOl
anyp1AIdSyajEZAh8ZD6HwCTVge1qKQXGRpEzM3sNEy5XU/+hfuJVscf47zG
asRihLCz6e0kZwIYZcPMpNMq1Bz5seGQr30aWXv+cLc3n0TmG+MEdn7CqQse
Fuqb5DMlmkdY5IWXdc3bsElygrZEsoMK0xSXukTZIGhuuTxWwRwjfqLgEsm4
x18zmcMLZ2ObRTyE3dwOmex3qsXeOpnFKWJ0R2O8h6sqH9fP13NhHcZpPRld
KcndsQ8JsrleUjxPSUHDoAfgnwLozABXfEgo/LF8wfQM61C/oTcBrhQJtRWw
hEo24neFiKrA5YMN5iYkbfeqLvYNUlulFONOuiiqBqx/MeyYnLvOAijim8B8
mR26IptqmHNsXDGjQURoBAJ0BU0oMRaTipR8W0yWO3xImxil+al5nJP/Srlw
NHRlnyA6l/5+pYt5aB7x4yDPQi/69iOyIw0X6vo8W4pVzh2sDOwQFo3G3Bep
Dj/Jk1Soh0J9J3lANk7C6yHADbdAUQcEFia/sACVUAAUlWyNmUyfbwwieEcc
Qd12g4fRzCsn2DXZGBaR0X1d9+uj87wR1IR4z1drrDAgCtLOUTOdcex8w8LH
PMjlUNbznf5ilfU=

`pragma protect end_protected
