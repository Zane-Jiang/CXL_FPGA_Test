// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tnhLUH5so+42XQbNj8BnLFKCuAIUbq8NNA9e5dhdEcXt39hlxWZ83Rly7fEq
wbkp6JuzYrv82iPbkGSDNKCkF7uAOLjDnPNmi2FHzDYA/k6dNlNMu8DoBn/A
DKr5gX31hZCdBfpT5twsHHRHa1zt83siEAyJSeefCelqlxixmRECm2XRxjF/
EyGMu2WHLARn/QMGeQ8X6zXP07y7XQDlHgw67PNPh53byLcbbQdDbiD3zpXb
ey6csgJpciVBkqdjxxPj3QjVsjUTZ5YxmM+66Et5/ZxyxA8sg6d/v4bMvV9P
yrhl7gf06DsSr4FtnR1/M5TrsFDtq33CYj9lx3p+ZQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R/LE0rSAf7CdEbs2oWCN5FeUJFLB3GPhKeintQfoHgxaTVkZtB0SYinH5d7r
SvolFrvaWEgjZdYuxzcAoBohseaE04cWJCgdjxMfs36tIgeBAMkoXuaENMqR
YM/VSLvOUMNydGBS5VWWiJz9+9KwpOto6t2SmJfuO1rjaJtHqfOa88WYhWxY
8hg6UikeoNkg/0SnFSydLwFO+AEcc0cqr+eAohPOozJQHe/MIOq5qEMNMiIy
veh32WOAhndopnj1ODpgigI9tNsnuad741rhym1zk9W1M5EduzAGcg2aVLvr
tWKS+2q5J88Mz8WX30m7Vqn+2dmEaq6FJtjTKuqZsg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VojjAmsdCUMu1qgxaXt5+6zy1yd5jtNYqvDK7gMnbB3PC+24tMPJ3p5Wx8mj
m5OtAWBaLY8J5lDUhsvPb3LvPG0hMvXuRASMfhjNkIIX36xYPVdyCaA+44qC
J4m52v8/dFiW2GlmzSZ/GqzLrM3GzSL2wLKKZSS4VahV9XEeDd0xkbP7NjoR
vrQa1el6/2Fg4S4Z8QNsZlwZswD7yMt3coCsULxos5bB5xLrDdwjkeyEaZn2
vzsGcaj4RLJ7GoZwFN1u76r79LDxM/x9JIxHhEm2q49BwNBt5bc0hRRL3C/S
x/kibL51UDhnt0d49i4cLxMTsqMhanagI12hmkoOOA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GoVI1Yb9gpGhbXOtDK0wHFZNSNPk8i2rRvdwY2ilZknh+xoA+0H3KOemrATV
X+Gy4bt1+mx7NXu5LcbT/Qj+90CZpqphqPNV94HDnGAD3R1bXP/c+N0KjOIo
og4EY8NeoKR9rgZ0f8G2IsVaBbsefnkWyO5GmpKG09167FJmwdM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
slXwpXcKN7Z2Kf/dj3gKxKecInN4sq+rrslnszmzgogsG1+JDgz503iJivHv
2tkBOLa0Z3c59c+a3jC/5q3EdoaXrkZFzhtUdT61vpgakWCv4jQU3OEr6o0V
AyrLbg+b6Rm9iS7b6kd/sZ2Zs+di6BzjwjxmbSH/iPLcrhQM5teBMueHBe4M
VQl829KNDiK0fsArOiLQuLB6aA21mEK+azDut/UXWpkZ1fFNf1M4v4vg5bLI
s6gO8yAceTgnl1Q+lS9II/pHycX9StB9Hm/Tx5Vwg7U3JiPmVLOxj7osqI4d
418QBKJ+3IFWmShkND2vryVOgu15qBwOrrgv8QDg3VTJjjyvN9QALHYNRwYq
5OmmDigmenj/zMjhauEBDlIGE4dEPaajNay5dzEd9oFXUihq4acIT9bygKLM
k+lChuNZ/BXl/lMa2J7zREYV3OJcprxBC4o++Za7VKRepFA4sPfuxENS2Ds7
F05DpGU6wWlaAeZRlok5klWm9EMCuS//


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PhSLwHcTOvT+P4AQf3wMxxN8IkzU16aQ72Ui6OVPA835ks3BGSw3z9mDNwMu
zjrn+BaCRhPzF2HcQW0SflQJ7AcwqsVzOmxEq1FxIdIalk/63LAa/QQhFO+w
vvf4EPE6g2nykxH9OV2hQbr+LmQEn09hOHz1Y148T9a6hk05gNQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H9PPYghusYM+4qPnsq2y6mBK1fviJr1xrg3zyYaG+wjovt0uVI0U+jNI0EUX
huP4fBw1xwJkX90mLFRfc5y2moHeFmjCm5GqJMHI0YwUofezgZyXg7kiaT+g
99Pi3DPnwl05zP6xSPrqCbYwURmf5PZoYXvqGYIv0ACWMhXmpGM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 992)
`pragma protect data_block
bXAvsrWtqCMnY2XYLQAGVN63yW6GhCYikqL0PfcOgNYXNfogz5K6lJvQyIlk
UX4VDsmcmFHAzMpcOKj2UmhIVsilmhk9bidx/yuSfGmBkkIavRiyK1Q0vv++
ZZl8SEcitqVsTIf5SZFuh1r/QTcn8bAwRr8wNXYO9qGoGaPWptl/uqnnac+l
ROK/Up9fFj1GggVkv+1zw00k4+fTwAq+uRbomFLLv4H1ghWUbBdO7gY32yMt
CyTG4raIYDhoP+vl/Q3Gt4GtJH54UlUbQbA2RVeT4sBCB50uCVle0SMT6qbu
QXzuJeAEqn6cffnZZgvvybT4OM/hRup5uAi4IMKCDrXbNlfiH3iNbe+OQs/b
dPgkjHcafpKPqS2F1ZyIs6sL2LLoaZttW6isGdM7pUs4mVay42kg4lVwuyQy
I6WnwAer6E2J8Rmgt3onjySfqeUzP2Gltxzve19jt4WaEUaPlHBgCNSLEN94
/rUr1rTt1e6bKrmyjFWoNVg3vqqIKET2UCfAgw42Usd3XUuu2CSUrA9/3leW
hWZXpRtGKo9NOxMWVAZiyYyem9VcmdFtuiVZQQ2m9D3ffwpJHNUWUcDEfv1W
cM78bewcely5vgvHvZaop1tiY8TDE2P/bG6WyO1JKrJV0UzHeygU/roddq8s
6CTaJHOAYxuU3HFNTP2GXv3ONinCdA4HIq7OCm4m5sFSEPefeTiCRvPy+nJ3
HznHeOuuie3XFxN2L4JoJIRYmsU8wuFsQpUpd21+8QvX2EFmw2F5AV01EDDs
6IkXlu76CuDCiSegHo9U7qu7O/Z+J8kxfS0ESFslV/fhNb7/2ja4etHh5U3b
N2Y4/+pk3Ua9Q0ZSNNq1V8wTV/mbQcWaIPfs1IVu4g5rpYIHOVW3L85JdExK
RGxJgNgsW4WyrqheMSx0CHUPx+2FT4LkIFvxsmzmbhRPF+o0Lh/4XNYY4jkS
6LRWaDlEQTl2RFK+zheby6Le7rDPDRuOhuaC6FYBP6HBuCOj8+jV+7muGe7V
YNUy4A1VBO7id72BWYXck8XpSUv5bmFEVmKlWWMpOzOZyGxzSQsmpTc7VScS
T234yl5o8NVCQ0BBMBM4vYjf8+5qZZewoFwSo4Usxttvaw6wCTT8M9tqLmu/
xplc0dGEGhRnzjp2P5LCyu1UWFlJtjM1lmAjOzlo3RpUCe6FldtFwH89jL88
BcvrnYA2GXmbFMYmDcraSmw4ckDx+bTcg9h03ZD59O7QmP2Uq3IZ8mVT2Zly
nvcmTjfK4Skzf5lAZl+gqdV2ORomSLrUZQnsj6CPprFpdf5juCfiiYNsRLgg
q3c=

`pragma protect end_protected
