// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
poP5tc/HmBXrxxphG6VH2NGJ9TXZdaipfLZMsvxUK5pgH3xWGc7oEaHigrkbhRbk+DgeJF8vxFMW
8Je9X/l0zQhJq6z4yn8faCX+yhX3Q/0/FRboTjmjFyDf81uhgq20H6Uw2IzjTfVFV3hC/5NxO7of
F1i2zLPASwRcen0YAJZcfGwi407jkyJC92KzurX4bfTPbfw7l4OqP5cvFcB42+VjplbFYE+0jHQb
Q6kfsBQ9wR9Gh+wo0f+xZRZ4yrVm1Qzy0O4cXot2jHNptm+d/XOY1v5DzrFUVAwwjDqwmbPEQT5e
+7UgGKRmtO9wYW7Qx1fIhfL7hkjFtzC9BkyBmA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2160)
VKrEqDP5fVhmBajDTvsndVg6RpOidUvs2ZLd8sJwE9ZhvY8o5QSxXn3DwS+sc+fqQTEBzuGfNhRx
dZxOK2F6GfjFnoblb77ZPXRFZWjdqcsbzs5U8dvFTTlbimWdQsIG20efGHzAksu6ky1sxWE3whpJ
BcxDmeNZJMjuVqOZ5twJGM2khW5X5B1VyIP0ngq7ZBxwYbD4UD//79D1Q6+4D133AHDq44sMCC1a
Iiqkcly15Pt6fhz0qSnZLSe4vYWTSBnXAOFrqs18VsDROr0yqLWy6IBoWLJCZscGzrdt6AkiMCbX
ba71jKzbqND/I2SThjEX9EY5XcEPVd7MvkircYWyBy+o5sodUhfRUcsR+vC/YKg/5qdSnt0n0l6T
dmmEJcvlB4z7ds42aGAPByMkX3fDCMuN3k9x/4XbVYYh7E2FAkoSG2aaEqIZh+n1LBp5wZXamTeV
/r5jUr5KcBFZEzOgcFtcVoVpkF+qObW8fu6LqLUgBX0a+yQFjrWzMnJ0jrIyKw752Z1mtck/0bFI
UYsKS3IQOqETfmpeWhPRJ6z0n4Os76NM04xMdnfRb45mMaOKwUkMBFJ0MQWX8oSYng1t+bOL6BQN
2GUp+1eMZGEqUzjeShyqZDFvJTXun9hvFg4dZvDKiukEfM0pwz73Ug8H9TbD9aijQRAVdEnu7EIo
v6dtgJZ7qAeCPLtsuAjfQ29utZGKozFmDPpF979zAfXRKeUzjjEW97E/2mv1ivhI/wq0whF+ZDlH
QgfHY9ODJrItdvy0IkuvRTnHFj0zovAGKw1CLVw5Wv29twSuC7Z6EWNnX3ZwwwEkqF3PXqyuTCXy
Qif88hchpturvG+/FCjic2iv7SSPMVIU2fGcCh7Iulfd9a+qxfB/Z2wA1Q3GZ4HnBmmo/9V+oYMW
8hjr1mMmej/9s0EtyGd31J1Fp5n9p0x5yJ4TY40c/z1qlod8haAjE3wVj51qikgVDM0DdhRCDCLP
EbTItxZbirUqCVDxDFV42na8QKRcf9MHeMtFvB9DjmATh/bL4+bU0m1aKhd57ci877gnylC3OVE8
nNB/NTw9l3T0rHV5H579CvKYCxjAiD9RuNQg6psYmhdy4adqA9skZiPTRxmMLMxcBROFbOCXYHdq
Gm93FqEicb/d3TZcRXLa4/EaM0ak2reE7lLJzJvWMOt+DfLRbAac3ku7hZjMCV3QZPxTlXkKdq9V
VlV84B+zmDVa7JI7Ax+D8Utwjxm+5G0qyPqZCLbEc2oAQbyBeZ2mZzjdhErGcLm2+g5IBh2c0YIn
5Qwk/ZrX34WDDtPzcIz/KoJNDPwd3y5O2CPS7qvZOn9KZB0zrQcn03w9/Nlrg991b7xrlpUV70uT
Wl/uw2YEyhs45fpy9MmF+IoN1+dqF9tSdXWWdPw2MRKfD0tjW3NJ9Afv7wrKuZCbzqgOHCc5/9Df
8GDUEflI/azfGoLYu1Pbyn+WNIxeWgdaZu7pzNNWWy+3GM9XjNdWU090qXI0IlBLwmdXGYbwnEzu
PQpEOqbtBl5L8om68DbbQPfSn9TxcK/REOHsEDNhAaX/vD+L6Fz6dOFj52gZ73r8bcT8yHKL41SF
HxtYn/mMUXpgP18Wasdq/p511bO/kcXS/GSlUuOpo1vwCiCiPCOELLU5oH6t+FnRrRe9F423fknK
BX3d2rJ9a9Gh607lq46SM8ijQa0cV74nbUWIzGo7FtPi3novGFXnz1eQt8h2Cn31DAFt+d3miQWk
BYxojGZUFGZG9Oz6K3odHjbTGFhRwbB53bLJ7CPkwqLzh6oU0b+W7DtLPVCIgHWopEc6PnKr5tHT
831BnI14h0n6FMGc8vQUmlB/5/m61yO3RE92iCq0pueNbapvwiDeV5XVEoZjUGM60saPlr/x76B5
8rG/zAIoiLhSN/St+etE/y+AUZh5Wkc8bVcGksgbeYefm9GUjgdK4A1uRnKueGhJc98cwARAbwRR
i5lBXCwm9NENpuKFXLygYXa1Ka9LbVTcvEcb6XrHiDNTQ/ARXYZWZb4fDdULMtH6uIyaDYoX8UOl
lky7l/X0UdiOBt9MV1cWVf5T/+BFaQ+NHpxb449kF88NB8eQAq8mwqYtJoidLVTIjA7uN2QsO2W7
k9XQJ43H7RNHuoRtP70MlJTVPSawlSRW/8HR/1/NIHjI33kGsSeTZLTXgNpoPF7QiKvgIVna0wll
m05Riy7a49mzOY7Rj3RokG/mv9jRb3aMhvG5p0aVMP3wXyhJNWQC3j8hAfDOBC32k5XLqscGzlEK
FauZwCPCAtNte7XKK2qcnGVOuJtoK3u+s00LgomfZONYzUt/iiy/Jf3N490wZCyMtP05+ZBXjggn
3L5iatt4VtB7kcvuot/lSbFPJJ76KNqXkMz7xzKFdQEsllu1nmXdTmKqg41sQeaLDAyCtsUzS9Cj
IcfcDEjo37Q2fUolsDHYOS2V4KXxZ78c1TVScfJ6Sk56LJNj+fGvwYc3jYNTFpatQfEZvFNIOR+K
Ke7i3lNC5L/KGSF1G9snnay4Ag10zNohfyMlgdZlfUn9uViYGIer/Uv3eMG329pqjsJcX1iCdzKH
YLRT9p8s2R4dGCxJSwMDoW+iiuqxunwvz5TomWoX4+j4rjuUzcthhgyXr5D+emHwrmjU9Ir9bdCx
qGK0Au+oxACji9Ol6d8m+ENjkAegTdGhB4lztCi4OYX+wjuefkyhayJ5Y2/CfQZ0mYH9hUWFEeGo
o/sWjgejoNOIe40NzpXTn0BSfU+tY7AJujhZJC5JnwChP9rjmOQirzCNcm+be3jrx6cxOtiAWHiP
fNlGG1nxZ+ygtYRs/L0O3ZZecgjbj7q8PN2X0gMs7jcPoiCCMkUQbkVrJ5tHO9wz12rT
`pragma protect end_protected
