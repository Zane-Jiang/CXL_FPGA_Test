// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rIoBPHGAtqQVbcdI9pJINMAz+mmixahZPM3v+WplPmuvBGuTk6Ab+SJ4grNC73uEyBJu4Xpe4GT8
Uzmca197fQ+mfgXKhbuizVllwYMe+wdM8fiQ1Vsx5iig+0078vT06yHxtN/2m2jfH6eJxyvEIksk
uE0ZBKpxWojbS6ouf6ZW//dCPhgG2FfASRMSzpX2XvIYDQ2s30FVTRBmyJ/j7E1gi90Ku375WM8m
YifVJes2BlkMP1gD7e7BNKj0oO1IpRYh4QBbTr7w8Ezie0kraQ40j5BRzamfykwRo0BhJSF25PP1
eF7TlsTLEGUpghpJDzobGmqXz/vMWZO1Et4b5A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
+FXbS29fHtKa13RZ6QQglfmWuxqfNrANdX2fgwo4kXzb0go7BLNdW0K7YKfOLxRuezyS1MsJRyD9
kB4vCpaBg8fCwF0UqP5uz7eXK2k7HQZWJAOtd9ZbaUFLjFvQvhL0hjYD14gpR/2RrBDbr4oV6aw+
px8y2MG+9362vijJsh7DeaXTZvDsMcsPdG1VFs4mfQXmz9J8yFDNsygV68cWlNqrvpJCGFdpsQea
+Xdydcw91k7RqyCPBqQjgr0SQiNBocLgHPx0SHQ85S3j3In4i2T35ylfJRdGTntGCAtoFzxorBfL
Giup1CskdwGm08wE2PDdzc0Uo0NSKxsvOemiydspJbvhjqTw/WU6Z0VkFZtakQ6LKDmriJTBQXlU
tVDxjJv7SXL67davHi56F9/ZPP0HuwF8BZJ30opSiU6gIPmhlLxvBRIIYGJViIurzw86ra7ExTml
tXpRGaE2M/bruGvONz4iPjvu/a3MB4jGVf+BO/2dVSNUUWrENjbDs3Zok/0Z3Lk4/Ratno/Z8JkX
0siOM2BNeFCu7hb7RX7Uq0KZfaJiIu+YJX6TB7qIo9jLRHEXaLIj7FBCtwWoV0z2GZq7791hIfF2
W+MdLfqFBJTgWkm9dlTj7IQ279khn0JwIddA/hVaw4VCY/W+XHDoHxUfYs5RC6Rc7BTC5F6FgLjZ
eMFzhSYpnMpJWPSYvvST/LoASBunfEjI/ksvNBmI8e/FCwaBb+BdyukdyfACDcVdioSwP8z28yGF
PsKQs7wksEh27Utjrgn6n2ByoqWwjLMcSRooCZZWLjZ1MQgehkOXQRRRfx2XclX7z0puf8fITB5/
jlVOCfoNSOGzdHR4+FUj5rAGtDoqpniZka8Bx6DduRri1i/wiOz9TLD+6jhaGuU3UNCg2VY9x5B7
/dAEw+yjzwEABJcZreO5G6q4lCzh7ckYog5SCpveqFGs//Eexi5VE38bREdk6iVkpKBYF621dBZO
9Luk140//NJteiHlWDw3fS5Ktfhu6NpR1CTTtyTrQu/1lFKaEuEXoSNAV7Q1UO26qAaR603PISMA
Pcs56HDhfCU4DyZh+zRQMGTnipLdPHnoBHO1KkxI8mU+nAUV7jSEbSXktXRukd/ZP+AcxcfD4HOq
6Zyr2+Cgcy1vYAY9vOotkR4QHNZQp0o0tRQuvtOwoAdLnNYlzZPcf1XSTri8K4k131cnHg5NzrJZ
cOZf1IHcXIGINPqG8Xrbf6Rg+kXo2z+FNEmzhT48OyVIpT6ff5TOqVm4ICumm4DClPCnKgSksxC0
hbQMU0evI/sR6XRJOVySwm8kzZgvq+ahfRIysQW9HPHBHd58gExd5VimGP62rtsvLnzFc4DHtJ7+
S4swTmPaFvIC9e25FG8K/anlSTkcOoQE8ltaI77OdSxBc/NkZBoRGNkkOdvXxnksWFTkqzokTikf
DGDNBLU5LsYgTqAbFbdMkl9zR/JFiS1nTKSNWh6CrKHCD5rAJtF9WFyqH0vSLBKvHuMU8IExlQky
EU8U2pnLp9efVt3XF//o5kmEFppWwibwF1MkPL/wMdsT177JEG0JOuwBeSkAM7XOV0R/xSRC+1aU
jVLCuP6tahqgj/ROtjo2Euin8yeCWEORJ8mkZ4CzQQUk1q9wGVMVfo506BTrMroly5DPTV3c7d6/
6cgw2/4CVFz+fndx4jROuWDEvAaAHo80pg6by2JBzarS+KbojaqNd0n90uyjxFZ29+ThxHUCycR9
uq0E6xWsRVuO8QwNFCYHSJbi3eop4Kw2Jclx4AwqDtbDNsDIMk8pzeFpyYcNlQ7m+znP9jillAWa
Z/8eMXKagXPh7vtk74XsQ8Qb5Ew6frxrXWhWi+J1O78MYLda45xREwPzuJVRCyXVuYaiDYN0jM1q
jmCSpshsJIHCzK5gCbfsqHQrLgwgub3jcTW+liiXKIVz/dQ7ByUjP2qk34v+QPxD1eUVMmlZlxcn
CPfOvILd/XiJpsx9ckwQZhoV9KlCTPCXHN42yXDvaS8p1D4KH9dS6ei1b6QWeDuHKsOF0ysYtbD8
k5E2euhMyXVTRl0ppYr38+A6AndhxPi+4gXlxNSt/FN9eE25WcjPA+RVrVipmp9H4nHudDYadgQi
FSza1xX30/LoVAwup6fD/IWeopPdEDZNgBpOZHHVq6A2Qh8z57P0nCk44PkZqoNLBXodfIUIQn91
E5q20ENVRu3OFhABZVis2M85kIMuNVP+B20+tBacBgl+99np0WpxuzZQ4pPQWRku2AKwNl/THEQE
CFTbF5/GSIcI7asqvlDYs9BqdDLRLaXJirIjJJVeBM33gisfp/gysTZErWYHrDsLvD0Kuv/aLQX5
7FJosexdmHYKtfCNA+YjkIypfIjcGH6P2aG114SKSu7k3G5u1tdsYzKVfOXmBsSkAH8upA54SBXp
Wn8cIytTEXYb8tspr1NEsKUDLAie3VyNmNHWDy2bKmRDccaPEntvrDcUU3OOLdVVQHqfzkgJSewT
G8Q5Ypdr3jTgPMsvfq4R6fCO4GOw72xupp7axb1ePhh4PnT7cFOQTfU3Jzg4ipiKhtME/e87c11f
eHxV0gjMddLBHxLCa+B/cyYff8nyTuVYcxHJCk5tVkXmrMiogFx4nVzG8SeQLr+vFIGRBrLMLEb7
gSYWn4mqdMDIQoH1ayCUu2uDmr4PXi0+He970PrxfrIrF4CtuapPEnOVYcQeWTYKssD1Q24S6QXk
j44j/rFi7FiP2ECXe1IVgQoD6/F4xSJcFz/jBgUFVJUqzsDVlBJYx1uv8nakladE+QEB0nUJrSMO
Nc8BNR5YnxTzLuGlRtyPDxeJi8YWFEYZnAsIgPUZqx0vjvDRKOyNyQk1uScDWdJNiv5H7UFKZYWu
ZvbHIch3Q+FV/W0M7UDuoRzLyyBgDQHKEpO8VxCb7dgQFETVN0nAw7PhR7v6mCin9B+7KDqaIcup
8oJEp81IwcOCKqYLiQtvvVME6mSaygIyG3CpAFuJ2+7qXBp1frcJC+Eo7G3jOTPbjEl5m6WQpMsD
GYi03xKVvB2ATQM7IgJ+YntkS+ZsfnJnXDsmeis1p4MJh807zVT8FL5q61l5iYgRc8UFIwkDQuSV
+JzObreYBVMWS7gvla9envIMqtzeQdMJbn5N6Pqc/34i5xtUs3mwc18l50L6sk53yFGMcaSTlFtd
2tdOASfCL9apSCHetmc4iMCXNEQDOukqZGH9fwxktV6YW9rZjCIWPDR2ykI2zj6b1If6VTRtgS/K
Hc/FyK8tfsY88jHc9rM/At525kFIcAQhvag/I5VMex9JEw6c79Hn91yV8hmnq77Wjixs8VZ6l7TG
QR6vgA9vzH41MQEbHYSzITXLCtTfR4iwCOUZxrPov6B2mH2syJ5IEMfACPSsF2bitkj2cDL55XBS
zAne/retV6Bg3z2UUD3soz1WCvxL19r2PFcZje3HNWlxryte11+mAffjHHKPINRrrgoYo1HmEh0j
NqvrGyJF5eZxRL1Eue8S+/41hyw7xafytIfNDAPWkKDmZ8WrNcy7Cz21XO+omtQVfzNYrxGtCQXN
o1M8z9gKKDOcwJj+WpymDMLgOqVZwdNk8mKqAfY5GZkt9NDK2TgpiT1iGd7E0QoLPUO8zGKK8V5g
GxipiW4YWgSyPHqGtut2Wjt9Sse2N2cRsPLssbp6GSgBVd1u85tq86Ha/8Qi8UDIo2In+06c8ucr
QEIBv+uJO15Odz7LKXwqjNfkuntI3YXZYOASiYiHV4ysOatX5j0xGK1bI9ul0U73yQ0xNp/GocCJ
VQMF72FU04ofoLB8JXs/U9HaHIaya4i0l7jF8gaL13ka3/Kk5uTz/+oodT9jw50dUiTio3O/GZ3N
jwhXAj4XL+SbhgsF30eAY4CEFABzZ1uFAngTQ3Bv+Gxmcg2sm3FIrJaatIu6Iq4FG+WXgTZfrxfp
N2HZkUXfpxoRp8aSnFIH80PRdj2aI6jUeBfEjkl9s29mKe1FQpgZ9phpvV6RKjY+XnFSmon+rWSO
vzYbBMHnfb2LulmZEESfhKMS91rQnps0NySFZYPYxdTGELq76HjWJHVsLID7QOynVCq5JCU5qww2
yosGClswGJIK185rC1IQk4f4ehYIoy97U4vFRcQTnBAZqvOO3+z1bZcC5uH19LOI2+2BmOysdUOn
0GU+ehq7c0USXr7lQwPXM2eAA+UPDUUy/4qUI9fToKeDALm2YqrALGeS/AY7UoxwMpdq7P3oe3Oy
u+PZdwiyw+mvy05Q7BLI2tZsrojRuF7vo/6+nfiPBrJZTq6kCIRvers+ab0IyTnJIrip73tOSOFj
8ZIrehIWL8zbYsvGc8oWv+YRcp1jMZQ3KxJriYQbecPcktoW+oqk48uXwPompN3Udc5D11hZDXPK
b5RZ/T4y6zf8umbNEXU7rwzfy75/CRSnLL8SBTYfZgP3ze/9DPYI1uXOu4GHAY3VumJahHnk40H6
hdfP07tGiaYlfsrSVoQuhc+iSR6ez1caBd9+xuT8iH/ZqX5LsILMrcRmnhB3Al7yudeODjpe9ynv
3L+uG2KGdNmB9yijeHfM/NoXmEkftkApj9/fewGEXkR4VwwK+E/89Blxn/hS9Hw4WP22ZqeQIRT+
D+pXZPQz/OGGTrEEj0j2GQluqpKprzQGuLcr0NHf3cQ2dwJI/mQPFZ9Mgc7l5YBwq+rSPgW9P0bM
2FwTSvG1gjcPW/1C/ES/pobHF4VXjZe+O2a+9B66wvt5OnvhMnChq6WeX3O1l1CawAt0+eANPJdv
F7+orn7g9nnWGestcNR0pvTvZrysxJDyjxHcm2a5356tL36kwgF6y2jeB24k1WVt+8zy3KCS580N
igde/OR8KBfbXPWGSwqf0/dkAZG0yrzObF89yLSW1j8A2fvM0Iys6sW/+Y7i8V07siYGYQz8PtxF
5DQDPKwC4DN5oDb6kZCl20lblstVnDTm0TsGtQ96Ifra1Ka95HV3tDIM3U5ugD8yvwgts3wEcJ5x
3Ac7y8gHgC/cLzGgGCoguw+hMlMhCZ/LxjIM0xECTGFWXPvVZr8LonPj7vUOwWCARSUwstYQFHCs
bCGOOo2p0c4nS41LrWNUNeweMhgDd8nFA+Rm7gTipnCfMd1DlzlqNckWc/OWN0aUhfNBAqY2eIrH
TCbD+heJmTIRxMhGolHOrLnewCIoIrLFBW7VMbhvEAA9Zb4PmGTVrH2e5KMGhX1ad9IdebAE5PGr
xG/N5VMsCwX+Ez7S9rcJTp/xa/NoScg7QprmWUDsVxSYxDS+fuSbRK4KEHPjIAXIaSzACmKAiqDu
ApTXnPw5ojcGevgDWe047ZTQa6xHYcMTs5RB01EyRIqjpQMFmn0pGVaI26MTaU4APDliQ0JRMQq3
btQkVowMwfybGRW1zKlRAAYEXoGaux8owWEwiM7+wSyLY0Efm4ugJf9wHvr8Mrp7dZncq39T+lS6
KqE189HKXLSdnHE+wfj2KsjxrJgnIMXEGC++DRdeh4t0hEWDkjILKFXi/jx3ICF5qQ+aZ6ShJgBm
AhTmri3+5k8dPxdQHbSl4ixlZ21lkuxChsm5pVPH2LjmM57Dm2YSLHZDFEEl8AC0Y44mwWw0fKDQ
GIoEpQ1QGJFYRehbgGLXfouRmKZHJLeis4s7rZw+m4zbhXg2loL6FwkzmHnsB5XXyTm80A0Xiogk
pkeJzp5+9ZRtuR8UtSQSV6wt9+eCeV2+BqZsIcBJ3phixe91+Iv5fWsKHHl7N2oMd6nLvSU1gRpn
bqcIE7MhJYsii9HhItpCEn5rTykNTCtXfym3VDMSUQ37MMRrebxPVPWYHHqQj/tyh/32QuI1gcOQ
kbQWjnTtxRY9ADuFMamVuNimJ+uvx+eWZFJPqhd6sWfD9d3GGB6Pdwn58hHu/D8C2nnq177L5ptz
LSF5rXF4LLWfEdkLuyKgi+U32HioxPAJXzadH5C5GLV+OUFSlK/YzKjTIh5fiqHgR3BdcyfkudJm
Cj22kyeMLm3CBql6gO57ox7gEDe4W/Y6iLIGYLX3n0VhxvVwvhXfeIjCTG5qjlqD4le+wZ+DYpaD
x35lJyEmw0Nda8BXHSxkf3iraJgFLpRpHr/j1CudECF+Tb0gGOshgZ4VUjAv2QDgu3HhZvzmxGEO
tt9tuzhsbG3bsEYkQbg/Axk9l7YnPuQUzi5MdgQ9XRGFtd2qmAP8CztFkCw5kUB0IC9QJrxS0ynG
I0+QbB/hgnvq5qcvYzLF9P7w88R/jC2uHCIZS085nuJTPq6hcQyapYP43F6E5KuCfhwOhfiPcNE5
0bczT0PvCsRCAAHLsfIRffzoH/a/GVdWYxqaqPrFP25f4a4bI3QcqCfPtCFjdgN4C6gscZYNR4ZF
lFJyqjAhfjueBbOOTXnp6gliU9iX4iyszKoqV9X0CQv/9taC0L8NKhSHrX3yDtRY59KRmjoFF7iD
0N6qWOrCvXy2avOXoK3PwB6h4KylmCzCO/i20iEwbULMrSkH8sOw8k/7OzuW8LyJ0Ak9tQ3pbZdi
PHQbE/2+G3uIRWrgGBfwuLIg7PmBNzzN+hxX8u+SiiLBWFuSvUetEX7Tv+2jJFElLrQPBtE2kEc/
wybFTXd0RzS+b6o/m5hthO/wdi1J9h6QzME/Qy8Wo5Rrxat7lUd85qwnlUQxLXkIdKC6UuI967s7
W/jzV/T6yfB0V/0HKonzPBmGayrYp7BJnu0ku4cSQwNjrb6GJbksCrujq1v4w7aASkRTOZIkzsZO
bamM7r36TFq5ikmCwfFwRLo/yPD2OIA4PMhbR03bxixVhdfDwzB25D+fj4XHDN/qu6rILOQaBN0m
+jVUui4sQDbReN9KFV5brC41qOXwPFGRWkmH87q7yUfMXrZf/rMd8c782yeYiMjMyDTLXKN3TV8A
6fzy82Es+2puxK2csoYCC+IAMElafcuCA87dN2X1itz4taoZVipNsb4apvOZ1ZayZzTnB2VDbjMB
hhyveTs308apS5zimLYXBs2B6AVU2DprADOZY2jb+OwGTsiAzBIheqfKL+sEK6PJX15b0ioLTnSr
Ci2O5y9J1Z3jrRSEggECdRmjV4kD7cNPG/fpaR2SZlHd4Dj73iXR8dT62lmcedySArPGcW8xPrwc
McaGhD5/211NXe1qC1jGwtfik6Yux0Gb7DATDifLWJ1t5aNNsz/cgc+k/941bxBdbSe15scDdc0Q
WKkhhrOC2VJEmP2mT/Fl4caVb7S3ZMfXnyh6YnTavPA7wyAfdEm/FAVIA4AQxF8W9TUBoBCn+BSu
ppTssTxK5t7mZ+Mr2F+PHmUM4HRfgIJ1QeF1zv5NrSmMOzuPm15Ltwt7R+Ju/rejni0OP0GcXAeX
qtSwQhI1dXXsS2Pjs3MhBGqQbRqhIASBL8VHth/d9wWjWqHhAH04IS19dtk/gU684v8upI1CpPuP
brSdh8CUxz4RcbDBYkWIM3lVu/G+ecKqsXc+1TwwkKEma4V+m+y7rpwD3Zu8gz209vo+BgByeO/v
xel0kPSG/nhDxKsCaXG72iPTHKgc0j2lMUKsFrU5xtDnF6erMZlG70TRHYbmch08LMtwOttN0IHI
Cegs/4dWpnX/IzKm60rNm8D0zJ0H7fVbsmIbycOklZN0A1jS7lReJhOY3F4IcN7lBVkCEjJPx/28
WIdfvN0WWy3XXG8hhGc5mdtBETzLsNkhIlY0O/yHgxVBeio80Juhh+W9cOI74mhDrPCoS2E3Anfm
aBFomGPY345M96bjr+1uum39IKHRkyPQdtQcsPAXx53rdcs9CZxrO7GBDnWeuVd5SZmZLbs3oduv
LpbTQM3avA5+uHKHALicVmTbSG8GQD5SfwaadAYGPczhJgAzPCHpr9CWYG6ZEW1KsPpX+nE7JwUB
DUVW+LR0lA98+Y4sj+ABtNkbJOjMbqZAkqcIzFvhqN6zBZ/HKfqELYNDXzYgMQ6fc4jWyQW3Zc0a
QsfoAowOJbeCFNQONwKsLhwiDY8GZb8hBkvDSrXpvRsWzeDaZ98ss3Cx74U3278K4lAX4Po/0cm3
+kuWL/V8qmar25ZP9kQI81O+HUMipRUac3TZ+9CHCO9qHyxSZG69iPCsRukJFQz/f7/ncFs/InRK
AFJ/1/3hneHZecQa83q8M2yZz7LjJfk5dY+b3IwT8DnfuxuloKuXP4jCh8o/UxGAb7R/kGXH3k3+
FlqYOf8/6GdXMNxT4iNgEKtuHh09FKmsyUEJY1myEcRHQChRsSWtkFCGrImGj/NgjqsYvDbxxZDS
TQCUlDFsd41lKR60QL5s/O1/lhfHzPKm5W03tJM45tUJfo3jhOdZ0yAwgqzShuFcCAmdzmNVHTIB
PsFDaLGFH7mJbLg4ioIP/L5mcWjdnIIiHjA26y2plz+slzBa/kSsj/Yy1S3nT8EwaLAxkNQlTXXP
iE2fxbDu5zgPvhO0bJDwD1tpEqdMLlz7OtZJfT1sbeAVJyIXt1BhmfjYRNroVC7ChgEbCuN+bLGD
15jB3/rHZ6JJ462GPMdR4QEqust4ZqxoZWyoY0EeObw1cbEZKzBCVk2dkLYu6dC9A9lpm5PliIzM
F31HJMCDxRXx2sAN6j86fFbQIYRkhmkPPCealtsSeJZGrECwW3FyNs/YKwuXeWCOkX6DBcANLXRJ
jg2jh7NSr2TKGUqC4egsFW/SON45uUkHfZziEKC+DwtY9pEAgHUKNYioZ3K32UDobwamnVyDnE3a
HYGVeb+VxN35o7yJvG7QVIZr+Qcq3+/SlLveWL8NuwECtdN+xmnkSTyULg+2J5U1AHxknRFgHoBO
zuu9E31Z0v5oa87wNSYeQxXripCj6+l589ts5E0Roj2iN/VnRU1LbRVtQSiUYQmwP5s+USjzGrUl
MF0TodI6+/FJNXVikbU+4aGNENylovF1Bxg2dLo45zR+yNZ4MafEEtFByzMdam/VwQY3ZGL2N9Gv
h01JhE86SvTz9AiV6f80yXD/xknbnwjGbHoBD+DIaQbITEJCCJcAQC5CCvxFsvC5p2eOXIQZGj8D
Vr3om5FxQwAdrU/+1m1Zbn8Vg/GndKims6Ml4enkuZwDEwVIEePyBZ3ZniTc5xR10kjFa0X8hPvq
XGd4QOIQkJYZ4S9CgEkIQJor8vWPfW1mxKNFVLJNKCB8iDM/+7mHiZGn2y4FtaVJ5he1Wl5PUyfk
vas02eJeJ41soSDIevTJLWFimPehJPkEzNT2UUKrbdBeTjMLYdtVWFygIJIHctQ3WEudMTzDN6If
ngxi3uc7/rWvHkTYjV3wtDQuha/wMRZsUR+abznVcWClSxoo6muyWHOw0ekgfOtNC+MmCZinpKEW
3la6swDEz1+ldRIwEW9Mn+54WeU7HCJ8lvSz9WZKIJkIgjrow0gUIA0lEDA1YHc8yGLVLBEGuZ5u
V+bn2aXXoSUxRi5XUDTegZWl/ijS5IBmQc9zYJGeVVVFuCUrbtOYWfjS8xumGX4hL1fOW/7GawYu
N9VDvCsbiyGyFd8VYXVBzWSVN3tnwyu9hpLEDDFqEJknJMqwjwMcX87OjIwrD5xfV7oINLoG2AF+
cEYDQQlCaDoOMo5xm92Ck1RLTX6FbT/zaT7IM9hCDbujgPYdXKpMA+bGVht26g5ue/4T519/hvV8
0gYwhYrDd1XuuqY7NfQ3V2hPorPQO1IIpnOs4MwcvgZ0k6jHW3dY6R5LDQZfSTJujEdHaT3X1KpC
x3ZMKm4yisYsIdDxFkjZqOI2KS/5/yTLhXLjewZWiL/EmAbQ3mgGIKl3TflBKFL901quG4zMUVe5
WBCi6mqZw27tiTDEcPZoheaZPSJ2Bon2LD2XiY4M44mCBtWpdct9q+hRze8KaxJjNwpXBM/1Hg8Y
VarcNu6fDKEY02ofPNMWwUzh0hzzg5HdvBv6oRF+5cfU+SKBj2GdB1OKsxh75XFjS1Vfct+FJPPH
qRERKlYMkYgbyi3EMAlxwOqqzWhzHrCaw/7SpxU3pB4Cur+DYkA33Hk8x+RTQKBjbyvWFIfXrQ0W
pfuh/464BsgQM5+wMA3wYA5xl7nWOv+4C4mj9XgcsIB5BsT7muo/FiQCRaa5pw3M9QRs+bCr348p
DUFgGpf1e6FYr+kWrEQdX9+llSALcEEiTfO6m96iMWV6Kmub7T37u7m56Tz1mwUQD6gH/mVxQyFt
llaBwPQ/vE65QTpj/23PeQptGGYfWtyqGC4e4YOo4kl+XKPESz8SGQr9H9F2zYlQM7NMR+RMVfKa
VZK5cDXV4B/VPf3xiz4GtICPnJel/QMQLASaJBeYR+MWA0KxTWB5mrKlM/KMgXbdawreWuwEpjLb
aiVB5kxO6r8d2057amHFDXCXrSImI7XlrDeE9M5KXgWhKqM+euTW1Ytp1222LAHnA+xXA6HRRrGe
Y/bMCOMxpvIWU1ZyiU5G3LbkvtROsstYzGLu0yhzyO8/LrUn+MvDkd/xvelWzI2988YPFc5i5XSa
bgsvLc/Zqhigxol/WogFZiLVtnjB3Wv8aYhaOGGMz0YNl5X+PmB1PnWyQBaveeq9Ne1iZMPm0fcq
Cu3L9h/2tdux9cfn6RSs7fZHQjDikltv20sac0H37cS7yyERQL+ZMpuLk43dSAjKfyfywrQI/xbU
Y0BAT7Wjgbzbe4KWyyHahmk/cSnLtgv5e7XRkmncncxN0ySQ88ZidcC6ZVDk/8Gfpy1j+4udj092
psuuOo55jjmtyB/BWbkc3ps9X/bWMbu/RaP+FMy7f2nByKB9TgUS+kb49PDvBXlxinp2cpoHaCAp
UEQVwWYSYSEeD9770i1eYRkbzALjTM5tQ+FxTue+7u3dOJtId/RSTBCifvL3pkXfhr8L/AFE0Zn0
1gWqJu9Wqxij/ZPJE5vhYhpMxQ7piyTD5/yd1eZnjDb1Q8R1vm2UXr/xNMsUevjE1I92HAz4Luic
qw9aYO2qjNkJ7WdXUQeG5i4BHfL+I2UOK9aG63KjAtr6e25gyNpo9Yzvnmh4b/0cPs/LpPuM7MEL
9hyn9lHcSM7ESVuWoZz9t7Eo6aesK/YZo5TZCeNWGrLuzSJlK4gzQGSOr6UYHwPcJcfPHE7szAbg
muxzIxXQMxK82Skcc1kRp3xuWX0PmLz2tm/gs+WyqgfPB+W6x6j96jfvYt6nqHFzJ45j+nV85je2
XHnC8hMCVcbBQKr68oSHFNJI9++TjBcVM3rExGGt5snaeAV24HVpx9GkKZdFdTlTWeX7KkYyoGTa
R+C2gVaYA9mBj2HuTRRXjhgZ6Hqlxa/54PWOsYZ0EoooHWWR9fFchQcTjtnyAxr/ffQH4X09iXG0
Ew058T/tDcbAEStgGhJYmyiB/j+c2E4LCZqHhpLD3fET059ywUC+saJVG8L7ECSkuo43gQYB8vDA
/droIEde4r2rntSTvmrJQJs2K5e30sW8K4TrFQ4OAwejIiztIi196AFyvLFl/gJG/tuHWGSjcKzC
dYV+869qqiMTUuhk0NuuxZ6Eqm9EWhhjZHgwLUYDzVbFDF/Hy250Y20hB7CYY6xb4Bt7dpLoQT6r
EZOBMXS9WzPcyAZPFSC4K7DJRn74TM2L16Sbn42B/YASpe7xiSHJWezZlxA7qGt069oZ0AD3It0k
hKY7dOLJNvhKdxaNkrAwZeFcvsxeYq2ZY0VyIYcCk3j/0/E7FqABAqnP21RTCJRKJ6nQRURFWMrF
iEzDhDTVUMebIN0hnU2cpqiLgdP7fwld2I3/zpSX/YhtXs49flUQd+DTQjE1nWwpZdGbV0N5xGsE
nkHz1pl+2FIDTzDiwXMNvqRQPkBU1lmMM6ecHg06ZJl5G/KxYtrU4W0RrnK3UZXaRikMj8WV3eNn
0UZEL37ifIZbufJ1Q2RbzrHvTCAEes+x8ZW4uDY16Ya8VZiTExoMAgqeZ0y5AGJKbqjUu5/GWIHc
9HN80Ng1Zo1Wveti/g355TfgMIU+CCCkV6h3je4vhuGwSMfsax2wAlYePSlDGtN6YeWeIIlqkWOm
ANs4xpV07x06BKotHvi5aDTgPT7JCwuyAbZyRTLxch7OCzi2JFGC2d1J7y0TPKta+xjKWxYd4yR3
ZjEsBWF9krKkNzimpuK29LqJl/mNh1IyjM6o3DRuXF4fGVvvakXlXrlG/GIrrEpwx91qc/M+cjea
FTfV5lpoMtA/zkUYvsOcW/uEUaA9WWb707WLuQPcnYfX8OLl474OBHcvlktnrUtGfXepdJ+cTaQA
hXEiJlDBkkokwGGZlqM2aEYohR/5JMo7aF3ukIJAMrEy+zL0A/2SUj2Tncz35xS2fuw/UwuYqfXN
3sBBtFR63n4it07+U41KgoV4U0xyXqtKqSfYGSMG6Mq6zwG6Y5MMvLS54pCsZUQ/H0DCG5d1soTs
OcXk6yh9vxKVW1kKT34H03t63cpZabriIRZwkzq+GGF+KhGbuzchEYaCpxCIAqje7Mj4BbI6j7qy
3jUywq97+dvmJyRnpYJDT+8gqDfx9aaAwHTwQMzuyI763tKZXtlBaQXEHNZKAofG9Q5oYvyxXOfl
NhD2fVVNGgy0B2yjeLw3BOMRrwYRRDQaRrEfn1p9oToMlsT4Xm36uKgnVjbuce9xs7LBySZGJd9T
fSXM6OOg+VVjKsgaP9iVH2c7FSSnJHBscE9HwT7787rzS54pi59lVf0F4JROB35CI4lXJNt8AoOh
ULyiIRvRDoHFHVGin71a4TPml52PJzgC0BXBw7zsc7mdAsuvMNIO+G+OYpOiz6Kab6UisZKfciUj
zborVjHguC38aZkTtkJn30DWgMeUOr5dXsGhyyVRGYcrRf8Geq5hEsM+yNh3HEnOPiEw9V1ghMVg
NL9G83fhA2gYDJqKry0faZk2sxK0XCfmJtpIel4DaHzZGg9Utq9DkyJxmX5GA+//MwnfhP4Rr9iT
S3mwIRrV2pRPOzF+3Vx81EbKU0w6yV8BaXNKW4glyfIrJmLSHgbCExzajnQY0NBlBkyXeDy+Ps5K
u+kxL97987n9l0oBueLxBURr/zz58St10ChbfQtWgr5vsqhg445xImdZ/ZIBp8paIogYR/U15Q7H
19II54HhSmle8/pojvACFXLXlOpj/gp91H+g6+E8njPhFSEEIw/FUZyf+kFY+TmoHOv+p7a5bGyv
2UmUfVnCSeLmAA5vBO9xB0fKSA26AOrINpbsvI4cc34XYo9j6JIChr3qjMYbEnqRLIM6r8DxOEP+
vuMGPBVc04ay7KjAqlKK/mmySZPg8/iEyfw2YqvxvYA6HI8Yo/1sk5Ga4meYm3r3au/pW0xbs17i
JGGH9qUVaxysbf/o7kpm76B7nr4ELL9Owkw8QhKk5391+ziY1/C3iyjrcHDGo+aCS/CPqtkqaPtH
Z61aLWDaiB5AzjJE1ZSvWolF3IUxKKclOBrNHAzoMiGPWgf1kCfq7rqE+Ft6LklyipG3a5/6ohBt
cWJ9inK3Gn4j6znuBPiEZmArilNst+NIX2w/EIB0tJv+uMxa5KRnOKxFlGePPj2bOK5iKgM4TSBu
Q4nseH54KWX0bsychCz8jR0c2LCGHOr2/Zs6XZTEK8HdtRO42aRpVoNKzkPaoQqpladjf4+axHl3
Bf5sCabQOPRIgfboIhFiYCRHenQJUorM4/zBgvtDmD6WJs46BBNHTBl5PqWlULSQhi/NsCe3164x
5sbdUPoJeG3UgqiPs3Qg3ihntBLIRPu/fj4kfqvoISCfcuAS2i2YaxYB0EbUC5SLa6e4RjE3r28O
9QnvErUVfvN79HDQjNfio3EKU1Xo5+QNBrBHxof4PzQ7uX5K3SB0sKhjhjG6n/+mmYOwFvnzyRYB
+ttmJI8v7BmH/35kLfZRkbzrM1cg3Wo2wHvQxb9JYfCSnTfvUV1pRQTRMhgXpjMsDwTrW5GnfED9
7tZxzRFTa8WA7+5RpM9swRUcVKiFDfYk/iLbKOxMzk+2Sg539FUBA4Tqv+MXBFM4ravmKWxvMjm0
WGoRzf4r9Jws9/URqS8pUn0RZV6Ps/CXy/pl8auSEZOjNVfFknwdD2gRltI2GhqakV87T1UOAizA
B26P0pmUAO2vc/9H3OrinyGPvUI4tzWURAM8ynycxPWXz8mUJTVimlk7A/PkCG2N1ZrO31zvV96y
E6/KKTWFIDh+pzRjp94UIqIfTVBN2gc9rGU58XyvXmrc8hXZjJTS3lW5FiegTFbkWWnuORIlL7Od
f59qW8rfLA2t3qBnFnuTYkpnxbkHVe5Bi7YDiNuSBe0U1F1EPJbrq44Rb2qDjpRnBgPyuAxNE/jr
N8WSAfSetFAQ4PxtEfaZ7m8jcWijkLYbNu9Bo830OXDVJTb7XDFIvarL5vMWpQSDGX0/kak9atyo
Lchqiv0TmRkgcIit9bkLuUp8d/L3YPut7qr7ABggUpn9T78S80CC6oYiOBPxdZzKKDqTRc24oIVl
8CxSInvymKEzkDNv+Niakbf1KKlpwkekZgIDCI3E+LdULe3bsd/oAIwq8g56qgnaaRzRQzgnQ72i
P8X0yrcQfrDIaXJBlhKHeEP7jSs+ALM8A16wuh/Yd3z9+0vbQk3Qa6Xg/kMupWYaw6MOA/g70so7
YMJy0xMHigRAFERbWr+anrsxxTzOTOWAEXYYUvsrIXCnbvRoxqeok/nF4QdzlxqUAmvhlVDYKCGW
BmWjhIhR2nz/qcCvE1moC+12AkvbBiv3D8YUZofTpdg2PSzk0vHNXmcil0G+7Nkbv0vgf56dwK+j
2T3/eJplkxGsiT5TGNTdc9jQewSRY8a66I7NELjqUGKyULkqg9JRo9mVdFdR8MEDyrguTuQ9C07W
DF4nXNM=
`pragma protect end_protected
