// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
agWGzBljJxbhBbGkhWNfdQJkLaSpcwrYa0wjlhrc/uCwJw3jrj8PcOfjdu8j1BrY
ouP1gzlZ1n1ILaeYuPX+9V/oO1zhIPCxUihojrnJCXnrRCG1feHccj/f8oDNicRZ
XGDnTFjWUQRYDbzAk7Ns93kScmggwpdyo7hh16l6yjo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 32288 )
`pragma protect data_block
zo2SKrikS1uwjiXdEmScyGGVR6tByg8QtJXUKoG7182dedwfQpvJ6vLk43vUY1jr
ZG0LGOTra9nXqQQ7UocabfdlS79eSkx/GYWF8PXJS7E2sbeaXSaudWlRLuv8bgRp
mD/pUDyDnSezhOndlj99fmm9gxFoJoQXDB/kxt6RW6Re6I9W7DTjugIG7CM12+2d
B0ZTsCxwIPmFhUJ20JG2uXdWQuYO5OB/u0iI5xV7WEFQJKY8soILx0R2vAyC/oNV
Lwx5728kyD7v8118CWUz8YDgZBrHyaMRT7WMnVTcoM7Y5wB4rdokvtvmDs/HNNeM
PvbwPldPkTEu0qBCNxmW8astEWPTMCFnGMLbzMSEzXCLeVc7Fyh1PeNmxz2/OK7d
EUUeX/6MW6GKJ05ybHv5J4L7NZ9qQIRK87Y/7yxOjmmhCSNE/Qzd1wNi4NpBmSvV
8HSszHQ13sK/RSz4qGKEsGyAek1tMJ2j9N2VMPpb6ZvXT43weknKD874RJI1bdMw
bJaOtAl0LAufAt2cTYwAAMnkYBYDx65PcxkqfzqscoSrj7GI08yR1eiii+f2lh+K
9szOM6Rmmh+l5Yo6Vrk2jBhRzAXMT343NAQi9uZrhcsgNjhO1O2WGM56765LcVAm
fBpEeW8ZzDBr8PGBmiB+OPyeDeXgx549cX2N67aQHZ4HvptXckfs2es0D2kGnI4z
UNL66qv+yQfLMNYQvGYEu9XzvL+0JjNqiLl4G2EPXjat9yXFq+qhC2nDWScq21Z8
OuwoNEPgfhHN96jyAEeTOcIJ0ZSE+gKcRShmLRbzvA7YX7BK2En0JxwBXDDA4w93
ZvdgEOWnN0IBMQQKAlXmG/7t4aFzjiCUV2anpGRfYIKObQqNO93aGNDC4Q7hm380
XdR/0AUHoTZlM2ZySidEEobUVRZUKURqs7DzaRKemAL+puPGTDPm0TLtJRm9v/qs
5W14QxpJQnaeB2Q5VcUQOYcoHV84tR6UsllBzyJPXum7mGYYrka5r4/zdelNgwRW
w301DsNBrFyzyubDtkvWUx56b92B9ICZ0U9ZFNOWdpTw0Qcb1ByfT42KXk7EXb0O
1zes9T//R9uhOOnrJ9T4XJMoDID1QHvcaI+3X70z14VQH2OnORuabp2O1sMAvwYV
GFmPD5qdRDtGTCGECLeMdf87Gx0K+hU8mBAjigJdrbxw0t5EgfZ7OVcsO9C8pdI7
mEXS2MwBeykksp53PKL5T23cenn8lPv5aricAhcqLwNlas32riskIbYwhJIrybiu
Cd/bYhdcTFr5mpdavQg9jQa4oYwaUxj2YgSQOpui8eqxs7nMOl3NXJeXQU2ZiAlY
JXVrDukwIvMaSMufukT0CkfIqaMANuK6dQ5Y/8J9KZm90BAlAxkL2tTHsrIS6TT5
I8McvU7yUIMAj27oewRPKisY4AESb8FPrJoO8kSMIWZCMWW4YYk19O72X4wW0k40
MXsPxOxZ6CzRNASF/KHpdJIiGSJyfXzAyhudOG40uCu2DwL2/y4orpFO7EMrvVwH
mrEr/5q5htK6OxEcemLJ2yAKYECGp3DuVnzWL3YuuIxpSyocx+5fYCMcftAX28RQ
OywpBkZOpAqlR2ebuoALK0Ired9SxOZxMZVjG6xStjiu0qGyjPasE1LyuGe/5qpe
vIi9Q3Rb5525VqE4OuWhzOCOLLAE+o72nU1+JZSoHE7conafpVU+inu/lJ0xzXn7
L3NA+9pY7hZoSQ1glefE2n8za485kb6RJqXukmOSMXVJw7jkjTpSrzI99JXkgH9A
xyNVj1iPrVLElxuvNJ3IvRdoCcSVFwThQcNOFzMkTW9lbta7Qt63YC0WkLDXNmgL
DKElf0h0wzZ4RUJ8Ku2HOauGSZmTgIuXbohSWyOAGNFWJ72kqxgd4tGYac5to8v1
qbxl4xr6+UTwpRNUSiWay22BQ2+AX7VoVMgjQmy28znTmUXrjqm9MKZh4upaHCQz
DlVOox93wvLoIcknwEY20cShN/AECw6aLlUIk31+HWn0a7Qro74d5B9rEVyNPgq3
gin4RGTCMxI0Oy+FvQKW+umXpqzA3I6yFePSaHbex2nIRbN0Llm846MrD/rGOWnQ
qM/8Vj1mcEXGWumcOZMb87tAOPn9tEWjW1i7lRG3SakYw09YyEIntd26mMo+no+I
pmSYVwtIZMf9rvAbOKOg76GNPo2LO0Z6wFy+P69heC0qHpOQHfGjj5PX5g6h4Xrb
DEUzo3kN+WNDqagBD/+R3BotgKH3+h7h4YxC65I/f+4M8Eucy21Kv9rkS1RZS3ct
16h4oxiCDCB+mwMguC9WJ2Z69qiIJMguLbuZ4vEzDNeRH8q9Fw/bhHBSuJoKip3t
T4e4vCShPMCbZLkCOIVqAGgIlkeMqb8mWmIjZnq2S6E0YRiL6JbvGREcTRku3jSb
MhPitoBe4sZa3a8eueFwMYvm9sGnfbq1qDdUh9AK4DRrNYccWC6dp+nnzbFE3SvT
PvbCQQTQ3UomsK1Ip2rf7aQJFt/qStYjpvf/uxGIOqkpxMuEXqo+64d+eXWXGBHU
Kxt8LYPHjCxMNaMiNn0Vszl4lB7rnOwGINDVn1al5xmM9e7vKq6C/GVO3dH4SDnr
jGkysEUy72ci9t8GGqmE5sYYkSk2S9sj4VinL2/gEIlxRKuz7kS9jGUds8DThq99
N/tomPh8dlDusjVoU2vhntQAcKlZ1NptQnzfp7wD7XK/SEH/f/MCR2BAjv5MG0u3
sfKXvGcJIf/GRK7/+adAMgdQAxReKFdn7izAu1JVDk0EY+HxrRT5gBoOsAgFlYN5
0HmnMfKLDarbiKu6oKBa7z6yX1UC010wgdZBhl/s1d+PR6NTXpnI7BT8DozGfuTp
jzE9NprkvChw8MytbyjaikRyoiU7kAxf/Xi9FxAG3wgbjgoWZjHZ8RUcZVS8cDJx
sjMLE+4lkCX9C9U3NJxQhQkAotEpTWsWNWRyKY+w6DAvRW5inYwPyigd6wU3Sau/
FSHbm50k8qKrNIxagJ3PTdsIKi878WPSl2MicORDwBgna0WAsmL2TEzTl8JzKjHq
x2P+51dPt8OjRTDAj4olDpDqe7TO5igH0Nj8HGa7uUqviZEDzjTagb0dyoSarF/E
CnLyV6/fzPptEtbBsWWzJYDh+yBc9s9Yg9VHQFnuYQBx+T02YiVAHvrRsKttomYs
s6x1+WKJyJkU8GFgVUj6iFjhkXqgfnsDuJ0NTVyi0SKZcQTjBN2QOoSiw1XVeqFy
9HAsdKdpqpvRfXvrZ5xVpRr6LRhCQvbWlZ8qoHKN+UNHzmmMOYpGjkjgJpA0QmiR
3LByorLPZPYORfcmHYYRKPDSpQTsqXseNxcxvNK8abBes/YI+xgN90petm1mjOhN
mgfmeEckDMP0QL97rq3ezmuzssOsoNBKH4XOEOlXuRSjUJ+ZqwuZLrxW4xt7TqHl
dBpi+rKCD+x1vIFjE7CpqmZBzqc4ncanEqsvIF7myXWMYS5kWJfRr9+5GvkV4DS4
LZG1VZjicoN/kP5J6EIxY79mMbEZgynfmdzWoGloHvtTavg0ASsthPJOS0PuTuAq
pwdfz1h7oGGW4oLSs12heNf9GE315Vd89tnJm13L9J1aXia3S0yc6wkNOHWVIdJv
G27d9Mp4uODLJ44M4zlPce29x0mCCXBqGdaE9aXdac72Xh2v8mH4nbvqcimE2HHV
aDBg7a7ASdh+MdIWBLLEXqB1C+UDO1tYhh1bfVaoklPlp8SEvyMF52iPe/DzsidI
IkQ0UE1he1eA2aS0kaunEZm5fM3pIXv1h9+ZWpRJRcDnhAe8CPjrY8+wZks5keko
ljlMEKjS1dow5XcB9jSVWDSaQ+cKDFA5eBtnyJwiOpmlB+SIRzmWleAMX05DDw0e
hnnCnz1axBSJ6zV1WV3vWTfbMfvhMUaa6rCdSJZeDYHGiAMjJ7MYkRXZPeOPfePG
vbhWHYLACdA2OCy2SlytUGIhWCYVNGH3abVTqQZxknbrcEvsRU3jVfeDy1FYpjCD
p4/OXbivRamqhA0ifXrWHJ+S5uuJT2MU4TM2UIDEnMfy6brocau9vfuAguiLGJvO
HENkNOZk7ujDKYov52yY04XYEQcmkjxRUaHVy6/yTPIKXFVHMDlXIdf2DBY8Qe6I
gqNUwfEwsYC4K4rlcXOib8pALHwXdsn6sTT1DUTADiTWE602mLSNrorzGr0ffcCV
zn1aJz35L3qKTeVRkg2lKlQ4pBuVsTP+kCvOYpft9qt4GyKyqSa53PViakxQZon9
76l1qZkuNB9Y39/dY0dalTXShPSA0jdhQOzNGVBXpW7svT/CKtwasO3ZJmiIZB92
dchuvz9GtMzjETLVpz9ACrTOXrYhVR4TifqadzdGfkvTNj0d2pmr/GXhXPha2fQR
rqfgKd6aqt8K2tt1B4MdQkBIy4WjEraYVnBNanP4WcBO9Ver4SW2ZHFd4N8QXHeM
d+uz+986eqEVP6AD05vsQFT9JAk5dTjo/nnAfnqC1bfJ23tENqvjifNcL46V5eOE
JK+5KVEC2X1/sWOLua0KuXGRYOQOC36eCJXev+7ECVFdhb6skV5YAgtqbqf12ffp
MYaVysjij/N9kewMEnrlT0ibUJbFd+741GAVAhv6IXBmMTs54Jf9DkN6DHiaJDoA
bXHSgkXbK+t4Qft27Eo0BalZ1hPxx1W1jeVsmiS72Y8xKULhvqwqFSLGEFC/wTBL
Z6PIUUru+DevIH+V26YizcuUXa5MMC1HNq1/t3uLsDn2GgMjKOSqNhFTESLJD8u6
8rlluTRQJuavde/s/cbUrQ2/7hitGBTlSnGLbO/U5atdP15nZHPpBeQIT+Xsx40H
LgVhht64BPBTaZFVbmJCPQT+WEZXdTa9VPeEcOkw71TB3AaKbGp4vhbCNpGFseDK
RBhSjpzKDfOJx6OeI26Fg33BHJMpdzU/dqm8mNWm49Njh4oJaKY/+mS4auOLAP1c
UEMlUMh9b5cXmmPPtMAHYooeUa79pdqZxTMVmdkKemp9nB9I6kzz006XDTfNH8Y9
7bULplpe5srxJpa5jLtsdYywO5kPphvuAIDCEwXjF2E+cyYi3oCdvm6rQjyhgqgM
DcfyGubM9DoxfKAP7YPKA79OvOufo7XlfE2DzQFRATdn86YVUFcsL2NxMxvX8xKp
mg+AwAVD5zIhddVfvuR/hyfs76Eie2P1TvXtXXjrAZSuf15S2kk0fz8GPI6JuOYC
bUBcnW5XhSps7PIAsedQ0hhdBfMUsPhRP2WirAv88N1m8zsjgOqEXeAgAl8+ZGZH
504vt9d2JidZlRKUQt3x+7wH70hlwDFqrh/NQvk9OvOIyDEEolQtLFgDeWeJ+Zl7
r+Jc6fg87XkK8PYFwI7EXxiW4nLOYtCaHoCD1wRNk4Pfj/7ECrpa64ZqPD1CnpK7
XdUtsikqAs9tnjEGh9Zhw94nd7TsMrWnxT/ohKhgxM+UISAzeeUM/dmCI0Y3zUaX
0ADXvN6XMY0FPElRxWXwlskDzK4ODgmPrHUIkoPUKO1Mxl8wIBAtB6k7F0M/mtvv
/YwklTZt5+vG1VgryJ/iXoL/J9Ok1kD579TCsrIuXLdDo5NT5oQyqXoVYwpxQRTd
XKl/VrH2F0BYs5P9j4bkuweN6lcshCMCTKmszoi8L/ynCwRfGJrHETSP/Xykvw+f
XuPKX8WQYssa1nV4K6LFapbTccVe8UPvYTZScuowF6Hvg+AvQpQFibZM7nsSLp8V
HylHB1llYKoWe5kEiVHbTH5fp6TbIthAyyCnstEqhoto9DHZg4dP1Rk8ZOmnVAb9
ZsxTOaU/ZYFbpihUcwnP6JmYoDKZIXNT5lmMNBAVzxhUmQJ4Egz4xMdDWmJnfXsW
H3l+B+JhSWmCvA/6b/YswxoLuRzn01plUsqDqr05G5kbiym0/0251yMtTNAf5T2G
mZGOJX41K8JOEGQjhVk2PFwmKOawsuawofmdXuAmjAX+tL+kALggHntkCrUGhEXF
ySDA4cezGq89Zi20EXOiy7dMx4LiLn7RzPzUCf5jG+4DPcA9OtrwMdWXfA9Wf7DL
lI7+4twSXkPPeTCjuG3PlrCpd6HPukpE+EnCmE4tUW/3qHc2I+VdrQnnPxHVTJ9V
SvGVFGUMfPewINYIS6aUA4LRmuYs9vnw+HD/NjZnXrD86tk/5CKXunQe4xCyurUK
UUxC3ddDQX53fu4IsW8W8MVq8YS8PQjyLcf6qbKyxoStV49TL9EDVgX/TpP8Xc+c
lZNtJwKwGx6Md1fqCU9ChEUznnl6P9UAAwu2qz71pvEn/t3X5QNGO+xS+xEh1tKv
9SXAzkZz4QOnydom8XeDtKq/0DWaLpIN8qB74+y55Ny2EZnE04E7xxBf+G6WW3Ds
Tn4/IpyIt203OssKAXpdTddaXS9Dmdxo93mzSHYDA6EVWMCvmjrCc/A8jOmGaCv+
v+B45cQ2IlnWVf/WdEu/jJj3CqfpD6JdpgzNJ58sM6azLFN0eFFmORoZvs1myuWl
LM8RqiWO8wjjcwFvxF3nCD3vL0B4j+SaKHoFMkbHhUHp4X/TgN4T80DV/C+fyPmv
8Iwe0EW4C6DQLOWU5kcMNTv2NPrVOin1oI1qIWbiZl1Z8dS/IRJxDuDFHBJ7WMyU
D4ZZ5vo4o9LSL/7yCOTBM5/2J3aYk84liHQ71lPsJPaMm/woKiC/8d+G3Qgl94Zk
h/zelHG+0TAISLkbZ/9p/DqFDqYOIZC3hx3Feub7/u3o/H/cDEHQlqalRcEBxOv8
VS1fCuJEBp/aHoAR6u/tlOzvw2fgMv2ykfpVBdcocXlgxWr9tc2u4bcAJuSIDkbP
0ezDH8N5vYehZ+T1APzFlgaUa1SHNxg9OvIaiTLsye4nBJz65UNkSupQDQK2nKsz
PDuB0Q9iJZcZStJCW+LTErgJrZoGkxQmIwd97p7cahWn+WxVObVWFp7RidCqs6kA
FsqHqzBUi0b7HD9X+V0XygL/D34DRIuqMWTDkSaFb02FkvkJAEmZYXrLm/u/xs6X
DMQ6cQUu9CAAS72EF1iu59bjDt0481FIoMmINp3BqcvRwDuavN1rXu0iOFAjc7BM
bw06NM8eVa/XfbQfS5D8kSYOynihG5WwEcWI4LW7g5l3lFC6zM0S9rCo5GviC6io
2NI0Z3dGklgoH1CRD9+AFzqQUuLc0/6eaw/KGCZPEueiJGru4M7urnvhlTKMlvgt
e0gwqPMuQ5TCzZuZ90rrr5CZvBItdbLXpyypOWCrSXDRMQYUTQ+XPNAEkjovJKSv
gwgfhtDyCs+HMoeEtezXZOZBqdw25bdGIfylpxFgpkoBzvjw4q4TAppB8FKpTuCJ
CsSN4FYoISdNL2hw3v1O6umKSqCOfA+ktcLvV2VmMiDk7r/sOz/kqLqEkz7TeuYP
MNOuBMt5TGCRdPEKB90j/viwmzZsxFMD7iw00iHwb8Us9D70GuTcRbcT/1Bv/JwV
OfnhUySzS416U9n+ZlC8CvArrwDACPfR8IgSJVl9GJMmn0GkNGXMzUk3Gm1ml+sT
9cTFa28pISXcXVimMfRxmU2H5L8w1dZfYhc0YjvH8TXLtThaTEJ3rrVk3facOGNR
xkBrHCBnCJD2Mv2hYUXDek2r1z6VgUViLitIRG8gLHppDB5RE2LAmHMX2qPhUvR8
DppLUydOkmRQc1xfUXCmU/vYc8Tg5E6wN4soI5zek58ScAVBm1Xyh/Rrvd1ojIXz
tgN7wnmf/5CyKxATODVqmhsVInTsVoEyGX7q/Mgs9KtoHGC+nE4ZiKvAlRhN+zfr
YfC3j0/nIly/eqQVJGLGn25eUbuN/HxDl4/7uyOfaViMeOWRR+jnsUEBBo6mg5KS
kGON03BIKCgdJZzVFheTyWlhCBB7YybA233s6c9XsW5jlBSeBdA4Z4hPfcHTLpSv
UrbI6Bf3DzthsyvUoPAxnX7kYzcscyg1DNyZSTFe2XbhxcWsy6lgphAfZBcqyw5h
JdOcQcRccBbQaBo529F1Kkk51GVbd9hvnCVn1zKeCDchFAimkRTDuV7Gn/p+7YLm
kXmHqc15oMIXe5nTIORJh4lPW+92tGzGKPdGGIXV0u3QPqgbn5dcljnyYdcTCLwJ
5o16piuq81HzXMnH34uzWBfhupHKb0De0vh7Jyv2RCKqE2V6DidtCQ4saVnVPzw5
amIRrO+/oUyYLd/uN15CU6xIh9vrQYQeTguYh5mvwjY0w3EUm6yMMhjNvuhDVXRZ
q9tseWOIn6uaxvPoEvR8p75PXIOVRGt0AQ8yJB+2J/ClIzAR+ZI07sPlcVhf9c9N
tR4eKOMVsN0WqQJWCNsqXtnWhLpiBLwnzHxGAFBaKvLfDsWheeM2Ctqa0bRygHj8
NBaKMnPoG8CtHKlDgFlNy9bvC821grXjebUABb7YPc5DFIRHz7Bfbglv8+YIJPLA
7ODHr0iFHxx2BcIioYFpDXVTNt1bHnm7JG7T4OOpfex+VMPdgQl6ZtwBSLfTdf8j
kbevfmnVV/uOVgYPK6Ly2Qkn0Z8/H8QdEhxcykdyXCQgKceanI70WaK91ygUJTJu
GnFtyFUnWKU7o6JKqY703vbUEUPlxnjPhU4zaBiuzpLM9GQ4QLhppNRzmtc9rLlw
Drj5ZYs6mY8fXlHpbln5qXCwMGDeS7NSRzzm3dqZweQJF8wuChhIiokYUhCrhbmu
ZjDqL3Xd4CP+iSKy3b4kjTC0ncfrcWcVOPrDH3AR4xLMCEezlWSUoQ9DzPtFg52q
gTRc9dVgajCFoiDugSTa+2rZTmxyF3C/SPL6lNaZ1enaIrDMz51LGw7Ei7qoZ4Tt
ujV4/ZARMjdZ6YaI8iZaTQtxEHS4eu7Btf0z08dHEGRX/5I5J4ovQHQqXl1hEw9p
akdzee0I93srS4HXV6BFHk1m7M3hgDNESvhonC99bWZS4yBq0VeK6hIjpQVxyXuI
29sqxO0k4uvdkVH011NrOTGHvYyBwKsevNnCj3FGnw2NUt3YvllTKgpVwQ9EAFF6
/Qw4x5jo34KolliXlfpHIxTWuOiLlSith1fvkav0CZOTRfnhqQ9e5I3jew14+u1A
2swwxSgvTylZG8dKdjgCTVRTuyORmRp/YD1e8UzgKLUl+eP6hNgwQmcbL+EEORc4
NVRFoo9yhWR/oTv+T51Wz1QPy4PQm+OOhriunYT8+5fbEfkgVMtHMDpkogRT7LFh
sZVRjYJ5TvY/MO3ewUzu1a+FLcQJjXNj2U9aoAl1HMvltJDmVdsgpXg1PQbX2lPT
IC9o9rWlfWVNfbraQC7M+DoRX2gJIthdD/umzuDcv9uK591YYNp7KRWIjQQ80Ayf
1vk9eW0WgeCL+wgp6txf6Zo8hXyuHcxHHkhF8viia0R0pVLHcKykcYCzxXo0h3WU
d5wdwvCaVDOGvF+lv25Um71CgbTwESYvxY+D3POHbOAeHY5ZnzlalzlNTlFs7Rfe
FAVNASET2uFugYezAzx+vGF/XEZutVLbCpSmGjDTH2ILZNgHQyonBOUQd1YFRlL+
p9BCe8SnyJgpJHmUFuQR8s4/xoaAJ+G50g3bN3IOMfQt0vklw3hepTj3bV3VR+1e
WF40hXAh2aWybSqLGmPJnY1ComziITCcEcgJuexQ4zPkj+uffn8YjmFxRhe3Ao5J
HY8ZiuCZUO4miC6oeJoOQddU1mqqwYbehM4IYN0/zgWWT0Q0Qwc25Kbwz2dxWUWy
kQTlaow2P2IMr8RO6l8RNyEr/4yZjMxsOkDOCm8iC5Rho+9f66v9rDUqehELqRvN
J1czDCA3lOojrSlIfsFq0YIfvHAQzqC90shcRgpm3GBZy3QxrqL2p9a2a6MUbN2U
dhpP/Glh6SqwKPRI8agCZEVLdi43F+DP3ur+y44S0CJcPbXe0dOJLEUduGxIW1f5
4sOn2dyJgpyuxtalu9C9MfYKcQuAirDWmN9BrduxP2fDIA5k5ho43548ugLcS+8M
DfSmaKiSUtIjw0gqo0FlgND3/xyzI4wpN4yvNaEudaclCExpQYImbI/FygtQb7AY
D3ZEdzEGrxl4/UUosZjBG1njsVEdXVZ4y/uarimMwa1CtF4sqSqKbp9fqnc8OM82
sPdLMMB+1k0KPdxbi5oOkTdewZIKCzzlEN3ovvnQuq+MAaF133lJI04CrM70B68n
GygqhAyZsFY+dFUbeuVUNHrjA3EQEC28XkuQyr42D3GAb5e2CBOaop54Hu6eF92P
WGesChlJnp8zJCkM6nzvByR/F9QdHhd1Dy0pEibZilZXSpkWC5pI5JAJRC8KOF6M
FA5of8cdGKdlfcAewQdxzJ8lXv/EUpgdsLqKtr7geO477V5VCvoMRLviVPo13Z/x
08uS8HqYB/zQx7fMpt4oZSBnEqugGqT5nKWkUCPyvG7bv6XUb1qCdBVjoP7LsFYI
xj2/+cbl8qCPUHlAlVLKTViogdESFAESiHY4ShSEZ49iUVuU+hSExPBKKEICKJeO
sYYo0BcsrsCK7LExs8HyuY7M/6sKPAoblfrc2sZFJ026N4uOSCPKmidFRcEpEaMf
IUOes0Psrhi5PL8at+PhTbXWQeGuAzkbfGUWk+kbJR9KBDlgwruiiR7oApa97AVG
LuB6mhurvezJw7DDoK7g0p105ZgW17TSH7FCUMNT57jQtmP3JaqDpHX1lYtLnCl1
9sChoH/vkwthcl6Ge6oQqACmzI1vCtn5zsK0+I5hzY2PM5ZIS6ZWQ85YulDhnlMp
KybD/iLcAU9iLetMNK0t4DALw+Dmi/VbjcRzVL5piiXg09aZkgovDn7V4jUsNcvJ
YmjZGn+ZX9iTxffR5CSRXBLDx1fDOL12DQq9O6FDVykpj6k2eRjJcvZYWCC2ifNW
uyS0n0uvbNy2Q3YDozbuUUzo/JJpbNqjthUgR7RIT7Ci9cppU6KAztshWxVs2JaM
whvO9xh4z06e3qTQtiLz5UM89tGn+0A5JI3TG6SxyTn0O0kAN9YCm8IwbPZlO8rv
zgzOtsQQzo0s6hdQ4GlhPABPvknfJpJhxIr2FOFyAJflmPUiMxZxgBxEKbczqiYa
0u3Vqe9iGAEAcXDbfyqy/V0ozqqzNwizeRwOvmHny74N2M9oJ0/NHEPkErWNDq3z
AMAOCloxzEVUNNswDIlQfTHxgZTt/C79oklFH5V8KoIGjJMTSrC6IW5nr5dOJWHC
yK/hBE7jD1tcsMZRhQjoMmNEBPebZvhczZAKZ7FNV43lzezw1XEujjGriFqBX4I+
RH9i4PR2AZQjWdDODQCQb/ABKXoVNnlQVA9oEdyeI3HO2DlbQJCrW4UGw2Alv8ot
PkwebgcvNlA6VU6OtFBSRiv2is5kH+3QMjxpAc3bUczRo8fEqw7r+fJ9+dnkVL8g
L8y5zoPZGyVEzUtTJmRh/wYa+q7vOhfN5IK+fIBI+EewRo+FMRpdw1KQdiSOJC3T
x4oRoyKbE822/eYsfaugt29W9ZaRe66+wCWksB8Tgi+h5ag64TPnOx8HmBtUt2/m
dWaCZurPBQWdW+vv3I0CCnIOvQ8fC6jfeLarX1I2KGhi3i4EAhczu8VR3Qg9jPtA
2+DSqnCTcWVP8/+tc6bsIfXaaimR63l9joZOzBkInojnsWA0j8Gk3hhTzkeEmxV1
wL1eBpgV6xUTvi4tqB/g6eG/S86kZViH836qrtdFLeyiSPhmLoVlYEFEHkvjKeDd
NAB6CrI13uJcTUy4iE/44Mma3NTGojyPhyBCjwdBMFc2GwQxy5n31L8735qT7JQH
xYiJYxQrGV5uQOIgiQBlC3CIUjdqzZagI/RBc4q18aoHQbNi0/u9h9lCj9MdU/Li
IiwKNr1oteuLppZcxDrq27Ig2GXKDasoo2QtBCBPxanGcipoyuxhLnYcF/LEUl9y
d9ajTvdsLiX2+e97+7Ku0J7R+Z3PMr8Kk+sQVLGXZCgjpqqiA2usAsGkAyDfczTx
dhzTrzvwKhoUgIfhw0BMKye923nsVGnCwKzzcF2FdnEA4xURvYeTxjNJdBO1FIxS
Jy2J2+2A9UXu3/1hJlPo3Mk5HrehdHU0u1YF7Eoiik6/FhS4nVoQhdDTaU5AkLHE
E7fZTRUjMkv2XV4pOPs7w6YVqeaUGXnFRhL2yx+xHO/MdDv++NieIeblfKa9WgkX
Xdrt7HMjvvfzdlM9Q+MUfvdrI25oZ+xKkn6EF9SXz/9wWghG2kXYhim/SYj7Wwu9
SoOB5b30iBAGC2dMeJIlFBH+jBxwCZ4XKbTDhjhyUujoyLo+XCYNkNh3nEGSEyuq
SkrgmGv8tEwvr0qWRace4gI7ihwmVNwH0vYa/2VVyCGfWgekT1xcW02fp/s1+YuV
GQ1jU8aYkyjqdw8hxJd7PQaP3ypw/fBMLby6qd1X/azChNDYLqnLaQtifZTB1khY
3eNeGLdCBm70nqNE5nklnw9aeUDWcjVFiGs2R//38e1Fz3DYN8W++Ig9bLFEEWbl
7lENHVNvNeITTKe7Lb1iaUf/VldEbHxK3JA9Xwp961SXZPbqc9DqS3L2ymVf1bZA
KhRibObbW5XDUWnBHGVQ47IUKFGQq7Ocqx3k8+IPJLyQjIGFd7FCpqQwR3n+3ZAk
7DmMoB+M6q1kJAg5gtURj11oZeUCIb9QZyXxCoRNj1uxi0U/SdDOBMfC2StqyBig
dNZ6J8vDa8Zis80lS7a2iCDKXY1O/ES4/TBM7hkWsll6q56Q1n3FFuJ7cGk8KWK3
s41hDsOx2euX4y92w2ZdgOzXm/gwM9G+uA3wBJ6Ys6Simu5juWSG0dlN0KSWa117
SFW2+N6wVmvTOyjL+HWWm+EB5vvfpz5pFWNEkHeKIosL9xDAsqcF2mPMJKj3KVLY
89o3D29+4PtAyC25IC4miRYG5DPhT79wnyKX95XN9qQHqnbeBWWjEorz2gW/bfQ5
HxBc7wkIFkfcHF1keAckVvVe+MjZizC/x+QamA5076b/NWusKxbqMh2vnFWeQlo/
KD/5SuEe7yb8C7KDi+/mr3em9aIdJ/mMplAMtMr+mJGDt/QWIbJW2gtKtZXLFM87
//4WnhRJcv/wwFTqtUKvEXMkqnimZ0qd4+XhK/De3P9Fw8XfCge954mBPGloQY7i
DR+0fu82LIdtjnJ1eUbzYiUB/FTrPhBkp+3q4o7A4ITQXFjoOHyTHuor/w1pYT2m
qfDuHJ2s0AqF3JZKn8+uyXMpcnYJo3s1+uFqyF6B+Ibrt5MPPbi2GqwsYwkuufVV
3Lryh7m27mBn1Pzyo0cTObtySDcjFCCZM30PHHKddPgGbxdgN0cIRykP+DB3P6ir
tNtZuox0+sxd2wF8EceckPpfjNZ0KESaTac3aDIy/SqYZhggpW4LywBK+qt1bLmP
au3OX9WnE+O+B2xBWxnhnbmD9FVXF6UE2T7Wzv97fVjDeuEmu9ZwLqWvwiwLBRlI
f4sXm3Pq2Br/4pwOXUlLRErIkGn6b8ynMzwTGkzYMkRT+a41LSb6MFhxBy5BXP6T
2E/HsYyaHhZm8N2ZeOuX0BQdNlWHL1rQCiL78dVLuAMHGjRkW26oRhQ2QCdEYS9D
YFwhqM3yErAZRUt5UMIk6SnsdEceGe4ZaaqokAJevlvDYHvAvWWoNRq3/KTKr7XG
CGFEeirvk9N7SovAmSDkGaAEcvmc3XpoGmgbDZeAYEzIJqxO47586i2eamFDHSc8
cf2R30uQFvG8uRLG19Z4yHHQxGyWEovHRYna6fVcvoTFUANrQnQbi6R9mZpDC2Cp
02mhtBsy7YlRu052fOHfAvAN3bsMFkuY1R/AtaIxz5DLVqqYw1b0dRiRAV1oVcBv
rCHxL8rZhPkO+adf/YH4zMgMozcABsjG+KxF6D4XcRZ+WKpwiyU+lvn4MPXdSLYw
/x8fsZfIu1FWgwNzdvirGBeDcniHbEuv61juOrL70tXvSycA2IaH8a8+aC2rmuUy
I4TU4uDEyPYCK682DGUUBQ0qwk8hFzFyX60/M4loB3XgakKGqwuh1PGbcF+qUJAj
Gv4r1aOkQllXLy8KHU6dnHaYn979j+RtBTjXieVK8eR9HeVr5IU2WpUbV3G6idNG
zhwShSbBQ24JsPiDPZSRcBJUSPtCB58ytVHByW0rQMC0rfAiYpzmfaopmE5iYVcc
NnTfKMlJ/p3/QHukWkqDhLqDPKlnUO9hBWG3Sv6wvD9w4tui0M2p1IVnraO7xCGM
osgNX5Xl17sG7aGRMxpeODThdbehUgeTnQyC7Ngpsk5Yx6D8FwysdJ/YW1iC31sK
iCH6F/j2QYkLvzhFcP3LSS1dyf+AzczLUSm5RyRykPbYK3GPse4Tq4ajNR16W/pT
zVN9X8WoTV2ePt8ujfGo8fzJFVvKG0Vj/1fnUoNFZsSaTu9ofIUX4kitU6vxcAH3
PeH4aCu/gdeOvfi3+0si08yzBuwuy/tGBy0UfA0bPndFAQPM5ij13zbe8NsBuMoW
2iDiUrWojJgTQJwX5K4mU+01YV8+J/7FYAJXf1ZvEorlw7MnxKQ1uqxBO8lVzqQA
Da+INR91btmmKwA7ZihdQ9hw1Qin2LAjXYDwg4QDLSaGTNx4Sy7BHG+IBeQjVcPi
vYnAZV73meufj/hysNg+XCdvAkpkrPUbSy9IAXkS79ZzsEEfZC2f1RLp1cyp4AL9
gs+YtZ73zQBNffLvkPf31UllqBf7o7ZEInFXM7FQe5jpFSA5yjeMWwZk4jXTmLeA
3NEk0YoHYs/LLiMSrTZuC5xLFSEiOs/FpjQJknn0CClgsM9cL006hAPDfE3nZZyZ
yal0oPI/6bqv147DAi9X3Ed7qLPXHSZjkEXcqeS2tQLQjbXeGSiTxwc8paFHs+Pl
Wl//g6VQlh1vKSIXtmd7w0UDmv/cE8YqpaVkHCadtswGTEYA9xJCgk/Oh8RBl3wG
eCTwT4KJo/8evTt1iVQqBGMQ1g/QuiT4amgdl6cDQwg7JOOp3GgNs4Kd/CgFGX+Z
T4sdYscQxmzn30rtj2B2Dv6k1h0G+YGEdpcls0z1URhxQxOToGkHFa3VwBAuuzeA
a3oVk2Y+CTzu4schpMMnzaCf4ILAC6pf+PuZhjTpKBtnXDpMg/75FMxdet3qT9+j
oJ8WOqVbltWPXw4lx3lyFw3S756ECeByhjMexSp/5oJ7tLgrivib1URLLXDHm0IU
D/ZbKKnxQKemHZlxAwsyM+nl+kXlC7S7rPnj4tLJXg5IFp4ZU5E/FA3GE2EcQoeg
pifS2dJ+fqd9w4tSaiKLkKndRbMQC+2om5rfIYiPnPtEi+5SKg2z01HQbrbFfAjs
4kqEccuhGKHHSkAVRCkJkfEnmikQjitKyOCLE2i8aun1ipxjT3O6eGMJ1yOUCwWl
PNhKTlCcWA44ACvn+0dB9csIWuL2804AIhgF+yOXk/aisUP13n8Ez+1rUyGV0mA/
oUqa/h1tt9bDlk145qKEtwIv1Df0NkBjIhztIZ9OQvrHUBiGyOmt7OiZuDt30d4O
4kbIAfeXcfn7lDpw6jE9f1InYPSyqoGREsYcrgSTaLNB2fdt+J6Cl+4DF9sOiYjH
hz2SHk1YUh83g6GWLRVsLQq8vYSlnRyETse7YpamKzsZskazunWHWpl8C+qVc0Eu
QqIeSCB0kbl27OGgJVlJYMKKIUHXbHNTBJ5dwnkw6YxWrNkR7e/7DP1lr+QAyCht
Hbuk57A1YUs8VwEHOPBV5b3N27xspDCt+Etq71MoVfo18Uizk2ofv4vn9kSa7ag2
k11p4qCH+KCf7xdDOgGTIz9CKcMENqZ7oe80hmDH0Wfm/E3Kzj0cpTZGr2H3rJXN
qC6rL9VESScUsCW9d75EKSYE7HVQpyVlaBDvm7A2ILLoQ3Axk/O7z8aygBwLZBDF
Jn3NaBiXIWP2k1JPfgm2y1Cf8M4SUSQa/Ek8QU9GBjv7MMImtKJDkz6ou6jcNCSE
mJXJhzk4TYSK+strjh3mA8Wi9KalAJ7oUQXoubHe/sEwe6HRvXl72oCblYQDEYjd
wGheYP5jYaKm67ur1iO/TxY9/SVQluYxTzGSZh+IdpjIc4VPlmoOFj2EByW8KQX1
k5MAcfzsCB3popNNDdFElo5F19AS8BjyOMCAso30X+tycpepFMlq8u9ahwXyR45P
Q8ZlQpBreWBv1U3mSL+XL7X84W8G21PXcv5iuIG5X0oU2UX2WUYurt7KYiSBta/T
1EqVnhKNnF2DJMZp7lyoK7q9nfgp1/KoHQUg8ygumQStL9olW9vOOwjfbJCk4J6W
oOBNamhKBXOvPCw9fqKmO4wFVwa9kZTXe2Xxj9yzlY6ju+vuts10FBPIpiR5Efxx
p00vaez0/yycRUDzqiurUda4/xqaJw/+8CLe1vJRsppMGOitFwMxMLVFLu7jwPxd
Luc/musokg233G1xzbOXImBQOsLqW6iiJ4zItdKxkEaQRxKJ/mDtmRsFb653YuIw
xXyGHD563tVbhvdqfeu2NxgSwGDcm8rJMNzn8NJ7H6tQWzG2whi3P1lXPe10IUly
NvhF/xzJpU7DmIJINIjyo3MEZCXk5vCQY0BZyUXcWRvCxFBEmUizqrbsroV6RDjN
vQ8rwkvSymIuwt+JbiGvE/3sXSPZxVbYbkkmeMQa+HmDYFPnUuW9Ta8cDiw6gxS7
qxP1ItCo7HNcjb4pRb0v1pQPkgO9U4ryVTyqTdvAl8J6dENu7k1RvSa+lScZdUfo
xu7jZl1hIj/sRsZZ3DU2q4FqiZxjN7co1jWg907291qQZwmHvb9hdTkZV4fC5NEy
SVldQ3A85eY/nAFAGrlqt6M2F/7KEGTkh/yF7B4rCpjkfwfO1faZaUbLmD9kJyD8
FH6LUYs7USn2Ogn5UrolC33lhuOzrQZZS+bDtt1FL6xbLUVSNoN/vffuG+tbJ2Lr
PY2rGw8TCXpAEfosGkkXI2mA0VOc/cJhcOei6L/AgGNRllzThEeGZ3+aXg4/NSNy
lN10EKBrQ+rru/FYfSTmfYMLIXEMz4hJOX8jzMRAuXntKc+ZqU/Oj590DQJ+Fijr
TNt3nN7Fhsh9tThSdIWUwaAX1HJz6yaj/UchRtP/AsQbJDFgbQ7mdqa3BIV/3qLu
wwUDYqoAjTgrvxane0Cb7fnLWuVRRz2QTaY0Pg/v8oUezqiz/Ejrvkae74BP+0ft
oi2bwyzBTSGID+NFI4aqHef0Ikcsjqv1X7kcUTbrfTalEGCVsgI/kdsH7qFbc9tF
LgG26yokMaB+U8pZMtHch0Uz+fI7awf3A9L8Lcc5EUuHmIDTIvBIzRuj4H7gPSc9
d03w+g0486f/cK7GILyJY3/GUGkjtnJmlzZm9Zdx/AMfL6DFRoQXvW0t9Wd/BGfo
MOO/Y5y2lXRn4GfXmgbdt2WbEsQl5S3GxzK3lBpZPqOnYgNba72YvDFkRBqcaMS3
Lj5HTpL0lujNyqKgcEPrrNxqKI6Z7XuCfhXV9fxcjJukKOktYPCTJsKhEFH6+EmL
4Q1PWLSEEpf6JCcw+gGS7lsDJ78DjdpXc4URXMMobAwHN2AI4G/oMKubWnQvLg3g
yVKPd3kuv+jQThdg0ovXQBjQVcI1mm63Ujj6rNfRj8a3gfP5u9pPD0WrZ32mIh/K
yeljKFUqg1OAgJGhDuE1fey4VrO+Ufrl2k/PSJhq/2i17iWSM5T+14rF4DrqIZdQ
Z8QDP8s/pxKy1St8n8vPBLJLDLiI50PYsDUMocWZcN/g/A/CR/CEnvyeYxprDNOj
fxGb/wdbeEstyIty4K2wjubDhk3fWxRawE8FLIlcMjXVPPv3o4PZcxlzYaEZuaIS
zES/+F1CmJZWr85GeQazpcAvAXuVRRolhqlmPbV3iWRUhVo86+9XGF/MhZLpCKx8
4DAsX0GicGXgkAT3X46dfUEjACtYTwNIbgMxb4Mv5i16ZvsHYRsYhfqX9rbrPbE5
TNFYVWRYtCsYwawSQKZ5PgmovHtzI3FgElk2DECYHzxr655G0dY4Bu2dQY4OYM61
OCOo3w8O2U6DWTDlQGDS2iF7BVESGjdhCHeQKi1mc6lyAB2KRS5zrf/vPEKvzrHP
bKg/FIPudg77QS3FDwQGcaTQSU1BIZCFqjUoZFOXCYRahFLAzpk4/KNqr7YUHyfJ
q7njmKVthX+GsjKNC6SKhFMANV+Etn1jKqmsYcmcBfZwSOFtWuhGLqsktOPOZqbv
jMNfzqdEezwacv5Fx5isE7ASd7se341DVn8dwD9b61W34aRl6lTqG1Djdr8IlacY
93X+6o4+REjuN3GPdKN59inKDP1ZKzPqldvr4uJxVfG5JK5sW6iQvy3ssLA+rsEo
/HXMNa+w1Kc2e0ZBVWFKFDAb00cne1tOFHBSGhULWst6Jxtr3Xkp86o5VxG6VT3p
30np1tVqnKjna/Ef3DveX5Gwgwjwt+IVY0MKtRRD1oP1Z+lK5OjQokqvDJUwwcMF
1vjmTzUxTQlGdmYS/lRQKTidMKQzbOBXvnR//TMSTAWfAqEqMHv4VtE67lpybCIt
+IWbO72D2Bfx/5m6cT4vFDWBEm7LOPzEMy1FskDdJjRf9brTK25nCuNYxScd64yj
bjskqIlvLS8ITrltR3lq3eP3EhTPwLu9YCnekIpwOMqsOewd++/ZNzmHdiXfsCxQ
mLGlsyB3CN3ljhhT4HdXNWRCaDvWgpHqpWeJgTklw3S0vpDEF2yUf7sd4npf7Es4
YTRelL8Gj88ueGmc53Ght9elTQ64DsPTt7qeEK1lQI2oC9C8ksJ2u21yKVn7UAJL
h2cBkmAo/wrqgH2iplDCfKZhsMLo3NhRjzFtzaoacgtHTObeDtBv1WIv2gDxbz9+
ElpTLU+DPZEPpdWmS22pbIWCf5jB1NmN+ntFFZDxWTyO7rL4DgN1Dxy3TYd4yHm+
Dx705chqJ/3rgMPMeSkD/uaLwF2SnnFaPsC/ka3/nUYY59DgRpET13nNfTiHT4tS
BOm/nCbT05xPjZbc0HVkDIIOCIsXjddjbA2JGhImMlG/PbwKkBQypojxPsR5smYW
PvnSj5G9HQ/Grdcjx++ObhNRiFhAkuHDqmb5WCius34nQS7eX1MxRe4tHHGP/HgN
I5n5uPsCoPTru1qptWeB/FlT+zVxtVlSNyOKFhBwb4+o4PiYNkoNiYy332swXv+E
gNUBQE2Jn40rW0oTKEb7/9NWVF2gI3T6gHvxtER/IAjzWUa/otzlQ8TOVO/hj809
XczB+zcrubFaURnVCfNW0uRhOIhogtTueVRmXSsP2Ov5U6tWNadcRimWQ34PTZtq
pr79VjlfNOcblZV08UlPEQTCgqhnhN3STVql+TG0PjBIPXCiCYEhFq1kK3+Xno51
Gt/mci1AhVpiTod28TgA4HiuLkSIjaNz+kAzMZSCGruDi9KdBLnR+FeMQyYyhCwZ
2hXimwSzb8QdiwQCYQcDvjjmWU17Z7ybRFccSM8My3YQfn3ip5lnso4UZZhPDxxz
0m1mVrPW7C6rbyOlDdL7QvQrisPUjAf9+ANtWwDHsdYlZ7MkhGVMLC1s1WHN1LOw
FyL3X5TUNlMphQwoOFl1XaQOGe4IYhupPP6LgxOLV1/cnU2lMO8wzyh9KJCIj0xx
54u+Q+OOPu5qkqkDQdMXkbVHHBy3PtjvQ73O2O7D1gzfPSL31yNcgm/5Rxkl0cd+
cr4FgpeMa1QpZQPTrj8ByU2EInAoR7fdwGCfBrl3u/r53SR5+MBVefXTVw5O3GJX
9tKAY/Ie0/ophA+ml5CDWFL6Y/oOO/iCTk9QcnKbxH/P6aVbO3xz9YP0KabdXTZ7
LLoNHjw3hl6aJv7bjg4y7raXAfccBg5cU+b/GIB/LWRRGX0DlVGbFVPaHv8wzofi
JyBTGPHN1T96JWCy/2+wjnpzpIBoUojdnQRgiIP4O3VSxr2HXWeUsfCBEhFZRuYD
ld1tPxR9rgksOrYpAta9bdyJ/TQjuw/c1cFzwjxvMQOG9qIck1QdfQtGicQu0Slt
ZP8YGjtRR1tJLUtHyOug6/mHGeCoR5if0wFU0mxrg97BxB7+z9z/cuQgsDInFawU
94BxXRtnYmAh4e2yyufTVk/SHwcO9J321nMCNZizP5PPbHONVGBFkJjzx+mx9W8a
IMGTron0Sd8w7WQlowykKT+PXI2DnmX+kvrZ40GBBcHomYMPgKa9KvfXtWm/WNyN
U4nCqW2+zP1hHUJVfpYc9kE7StBrA0KLdol4mOlq8ZPABjpG132UVNNgmJ8iGCY7
PehAbp8QRNufn0gZsIIiWRE4aCwhU1ceaboJzeSvEWyl/nDWLhnj7V6eQJvAUAq9
t3NsK/zQxuL5c4iETILxoe7P8HApk3i4xfDZ/0FzWmAm2mXtRX+ty4tcYLlAyk5H
KLcwV8uM9SCVxXaGu3CsLdHBLZLfOVZt6gIcOs9UBexpCpcW1fY3pWQYRK/DqvIJ
PKFRDA4FST+PTI0ur48H1Npokp/B2ZUG8Eo6sGpA6TZOk0LsrIpObkX21MgvN/76
p3cFLWxZbKjDKy0U7eYk1bvnjhxhr+jTy3qzhLPZHH6pdHZ5nonE0/iBlVL5wy/u
YwpzJY6SlwJuRCginpqYIQFRRdh0ihuLGpgZfe1gB4dvz7X0Vz/nWmMgOtIbK1W7
reeOJBmcDq9NnZtoRAUv5h+Tt/43QJ+5q1SdpQsPIN02OVyvNQvalnZIRRTioeQ+
hMamPsMKkWnxl1NzZCkyyq+p3EEgNF7yaLtyKsvE0i6ZjfBujaaIRtJty/WcO1Eg
QkeFmsnUrl3KhqNkWoahMLOtSe7Z3ssF8rvaBpoXfHqESvR4N231jQicClIW2mV4
/BhjkYyYZde2KjDaY8zf5ZJkT/Z2flODxNe37YS7CQ6VUsZ6VueGaPkDRFf/QW4O
VEcB/9CORHVJtoOBeozJTnZz2VpcnEiLH2vv5PmHqPs3cz0oc3Xe64D6Bqdqzh8q
+ae4n3HoyYMc/4CilDa42eSj5w4yP9bNCsOYXly2V9Wn0YBDkc9jGoq96ZGGf8sH
0cU+HIdEiOQ/ibcRxdrI5zqv9qyE5M6irx4f4vMVOp8dQztiLTyFthxfUcF3Aj/k
w24Th6IKZXyAie7IMVR0TDnZ+cFfSMLt/2iq2CtaUSWz3JDg+RnDU5gU+JAY5pwt
qswPYWhVDkPY8usC23q+K1Xc0aPIPsMhkW/4bEIVVfTPOi0Kj9SiJuaXj2jn67ex
ciZHLQ9wmkyLk7LK6xUxK8YIfHVSrEmJr859Lry2ZaWVeQSdTH3XlHollTKImevc
lW/SZgJw2D2YrvXX1i6o5uN8SPUByVZnsJ3DbFpg78H12T/nj+VxuwreHBPFvR7g
CtR0wFoRPOboncDJPU1PM5/SsgTcDKBXEeLZ+B2F3ahuuqAIQQugP+2fWvMyWbOT
ArXiTJ54xanwHO3y1LKLaluRrRw5aEfyV4uvAH14wcU7vGlFjNzFZVYCGjX4Pwyz
k4ldzsGM3EI7VPLbFh8petpKexDdIU+9TPhLxxOoB/bBYpyt5TR4vocnUl0mIlOK
riiuX07GfALUAw+BaX7f2TCi1kDGkpTG/5om8mZDTTz4QSrRkTxV+i0DSHgs4pEc
kxpOEREELf7Tu+4Q9w7Jf4obwEtHBbGI6vzfJ45DKdpRVh1HqLI3mli14SiY3jI4
f2JCFMnBbhfo/i5YNK5AMM0NLbgK3mJmz0CDNAF03saD+D5qaYO1lSzRfU2rBGse
ZljqCu6kKoW28I3NV5JydveIwpmhpQpeh558XP1YWP63wf5t3GIygUT0/5QmSsBC
AjIKxfrYc3yIzFBUX+2UZ2YU4DiCfE8ukD9IkTl/4AbeQVnKAhgUaW/zpx5eAzec
z/55xS1fREOFoMFP/kmilv8ZDT1s+kupS8oqm87U3h0+K3uXYzstj0Zbr+weCfy/
mHXexzJKYvwQm5u1HHWv56dKHRmIpTEGT7i36/gRW9vkXClQZ9VoU5CZeGrihV0M
p7G2WdwCY+IkbN7Kx8MnqsqELFCHEOtyo5MEFiI8VWF86HoVj+t811u8dzyemylR
fSmPwelv42TF/mX9867sG6W1inlIzTgxQr8CoddTV/jFrxyIonXouCBTGxQfW60k
W5uONR07f4oms9EvQ7UB8N2KOEbpa4QbjCf7Ms/zvwrf42nR9iphuJTRwTGNWasA
QtNYl7CSSL0YW6UWJlsud4KcrRcbqRDZ2D71v8rYT5QryqZUmBsJfhPI4pfrbGps
ci0pfbzaBMhxsSHT5yj632yyFvyRwmIXhnmKT5z1Nde1/Y2D2z/EzvtCxML0PeVH
RGY38AnHL8fFQpjH7eVZEtUcQ9M5PChvPJ8XXMFErqucNAOvn65yLiaOiLckBVBx
h7VRDaP6eRQVPUor3MlzUX5ir3V//cXjMiZMDe9L3vvIb02LsqiygMIYXXVCeY7I
PuVSupyZy1pv9vAARNhD73lRLmY73PUoFOP4/z3vXkrJ8qKb8/YDVwwweeWpHemC
J8XBytao8vGlsRjYyQo2Z88lNb464WdjZZMteO/7XXl5qy/3qIr1V6gpDdHT1ACG
se4eCGJNwDsCtdnlFKQJJ6Ppq5Ndm/1jlHwjl1mJATWmQLPZKCF9NLI2aKJgApE3
29AfJsIZ6yQvIeqq6hc7azJ794WbwVIzV7WE0WfqH4FFLcgNSUd2hib5wmO3JukQ
7RvqEcLXZznvx3mJcuHzPBnBoEO5r0e2rEz/U8oqftZ0swyGFOP6B3OAtFJiBiV8
U6choV8ypz7QOphoKoLP0qG3v9ejoFpobfyTRuD3oYlnePPmLSp8U78mOpH2qoSa
d7OucmZWhDsKkgCOb6VrTAt6Q90KayKgZOi1VCuL0YaCnH4NGh6KJPN/56qoHQ53
CHsvOIAmjTUcMAU7WSIIzuJ1sHz6jXO0lcL5mgvyxYm5AQAr+k6uos8oUK3RLoqf
eZwJCJDjpsiPP46u2/IB6mOWTxI62yvRNMMu4vGZDnv3CWLI77cbtaxQZjtpDP/u
Gyxi1ZVGFNexhISSEvnv1d6GrCZmbjJd1MsrjvDbpsNTLm+GbnLyfzar6CTyOr4y
f37JVrxsnttFUZsWRKV6a7kgiT9rHVc4pCQUVmY8vMf1sEHhIQBAlnKMiSUSkQAq
Ve3wgB74LEEMwbNmN3qEgsjsw6esU5pP+X6J4C/ebu7BwkgPcjU62oByCu2RoJI9
ROY8xInCHAOrfvRNuJDLX11wZk2ap9nIW7lj7rhgyIxu3uss2FnZwUY7riscn4RD
ZWaU6CZ/YKM1FV3XjGhQuyKw3Xsj1gdiAQpGdxJcOvBWPu37og/Xh55jogbAyp9J
ZeoUoETlDAjvieV6Qn++az93bEOb7hpMDC17HA0L05UP33c/Z0ac80gAQQMggpj/
4Ch4z5fyXJcPozHSeJbE2v2HLV4iusWr8oJm+B87jTQb+UtR6gwLo6ofLp35ZIJ0
UOjlqHL7R1A2hiZAGpn/MXbkrbN+5Zrdak4wV2NX+7X5jA67jZLf3r58FjoDZakT
mzL02a18Prp1UDigyTESBc1SEB2BobS9pMc4L3cElS9isQzOGDfZsN8ESgf1S710
gzwjl/JW6KIs1lezTyauLES80uB7MX81p2D8irNnxA41bv/0eQrnRY78SgLeGCfb
vOwD9FHxp+3f26QEv4LXqlFvfhypMQUtTAFjefJy2+NAC27DHVpR7qL658iwEwzG
uLoWWQ5x9YHRxFnqKN9+HdxIzTV7/Rbwgxce2w14Z/X7r+upebQJS6CqFqQPGi8e
0POecaZU6FePEC2fOIlivqjg915O4tTcNwwLbEKQe87L/g8PyX9efUljnGv07amE
14+QjMpg0+uqz3GmOY2PAbEdoA55yf9K7QlVf7ckX1BkH3NywfBHtkgUdY86O2Ox
kbaRxwcI8IrspmEnYcSBwTPmq+VPY7VzTw/atGSgf/GdOSDfoEYKWSWEvAhXTRX2
iFYjm1+1MucfXwuX2PDm9ba1C4j9fK6KurkxdaD3GYSDijBXvNG7BtTNe4ZxQRdS
r1sKLyZHm/vq0X6xEVuxEVCm62aNI/tvr8n9/OtyPgzSMFeD8k/+gYQK6typThgz
/jBs2b6dG8hDqH55IX9FfDeHkK/drDLugWS0dqjOPjvWi/hEqtJ5x8sDBxq3VKaU
3272S/iBD0gejcnlGkn1W6sbNr2k8X5753IjYXyMACLbsvRD301CzEhv1u/vsmAa
Ol//T/Wu3L47pfhHHYaGxv8+A6OVzyrBay0UPs/j66zJBCGd6yS9Kd8QMW0W4Aaz
jw7rzOM0o7WKrBqNb8vXSSm17rs7aH4DCOJSZ5QvZbpbVa8hFQ4KmmPjw5eialVj
ss4H4MWhWESFQa+hOavPYpAJwBbN8oGlSHUdCRVD3FFquUHvyZVlBs06uaVW5XUw
Cphqb3Qv1G6Nl8N3995IKaxw64hzskK1VeZle/zXVrNxstUeQXwLtg8KY30iVFIk
IhiBr61fNDN4HOREfASviqvlt2+sRCDQl5VUwBkCnvTpROTzTE8XTzIziyWuJO+n
6bC/ZUbkC8btit3WkbQyR+XWdkJ/hkf1lD9f12YmbY1XZ6krQJWVwD7zVumOnjIe
OHj+RcEY+KlVbRuk6sW4ELkDRlNuXZKepuLU2NozHE8PY1A+sPPxpioXgXma/VyL
+V/i1GhNAOASUgCqkR/Gv6/NVqBYM808iYOGAijRjQjIYIhs4Ic4GiRBFXuDQchr
b5894nC0oFZlm+ipgngTE83ASY9yyw92qNq1Xy7s/e85E3fyb4n0xvLM41s8CQpo
CxighrWZZ3hoTTisDHRWQWr9u346HI7xQ91tf0vQscTtweg/NALi5F9Gi5C9RzhU
PTyTzc0prwqDs3OO733DW2bBCQ0/Txger/cJj9E9CtP24JXwFDzt9wOtjoAT0rKX
a67PstW28V/UXqXtHhpIRtiErfT00iMaASORhn+mUI5EAJqLpR2iGcPL3IfjHyOY
DVd5zH6Hf+N+m1slq/H2J+86bpoHJxEnthAbI/9tztmC71+X0S/PA7/uOTZpuzd0
B63BwVeYkaqIVMIQtrKgxyNuRS6dbbvcWZtJuYbRgiF74clDvA55Sf1nP3Nttr4r
jKDNO0ENWVOLCV6tCPEO3nbgiHDr2Wue3pEDaC5Gs8NxNj15D7OljJceKauOiavi
kd6frEFzjNjw6j2gFBR/q9m2zw2R1v5UVmuxAiWF/hbQ1DWkI8+SHy8yo5HAcK8s
E64T3bRCBOF2gpHwjGyjbNMGhU4tBP3RWlB5Ogrr1TGuFVYCCOWBVHyP+FryPax+
RzgG+b7skJxWcGDE92DU4+HG6nH/MJtkgQvSPmXGpLfwzixF2f13u7ZmWvF8dyll
3079J34+8kaKT1o0fWd1QmHD04anTfF8iHnQajMO1zfwV6ZgFrIHoVI55huA7jiT
1H+mqAoTN5NOIQio07NDdHBDFH5d44MaL3CLOt3M38PANgZ+SLy+eyI5U9bdJeVN
+Z2f7sVoHeGBdMmydRN588bbhB5SK5yEYgaAdlbShJHcz0YEzhBH5KxqeHh8JyGT
/DEOSZ8G2blrybPlBz1tqzCXL2RevF/f+vQgeqjzE02qTmIQ0r30HxVBttN2oINE
pCiuQNP6hZKpmf97z0AizKk1MXfR7sFa9wn8FYwGqPgbbBdKRBmnfs+oS67cVBPC
ogs4Sw1x4/o0WJRpSEaGlbDGQqTsEvPczKFV3X75mlGi3KMfYJW8K+v31WTwABh/
ZlqHTTFoWBgL9uraSvHSP8RskQPYM/HR6S6EBW2BaCFmeHd1iPto+Ik9ANTzelcn
y5uciNKIVgKDtnPVTCc/fqZgd2NA3H45wvWZxkf2SA+z6S0LEUjA0XPxAV0Jcfpb
xHT98EIGLVCK7HJEwnkwyZnKVoav3KAPwfI0PzO/FabdezHz9tt9EaF1Tfvzs9AA
jGtgKOXbmOYSOE8dxmNhL1wtXeCTIWuB67bQAgqjpXbvsXFWTCURpGJITPNxC2yr
40lrdisW5W9EFdQkWn9T2cdgJDzB5I7aUyCDcscED//QzpdDObnTqFFpS3EmOjfq
GDhP3SS1SHZeCxcAsp98CJU7MKTuM6vR9hdxuNpNJbzPiCsG4Zu0Sx1hLu88JWSQ
r+A2qfneSiaQjBg7r2l9qwACG7Y/bTJPStfgzoIDxZLNn3VuzTzqm2TBHTdnC7cf
GfFrU1EKL9gY3/84AFcbi3F/u9wvDAq7xhLRP0q9p39kTsexO6niCbnI2gvGqo1M
8UghO4Q64ti9DH7XEuTsmTmIq2zwhfsjiM8UX6X5Sm56J6n2EpK4Gg4ERLOQi2tH
MfEYVg/BbD3yNsmd4mn2fascLS6W0ameVHMsuhNQBgbwR3D7Z1kyq6hOYKCvwLB7
ahG4+3SH7IJ/xZT35SzJmJCnMKAhPz/PlRSW1Nw9+LCqR+BJngT59ZIHwsOgZS62
aCoVOYDPa1qQQaFQJ2stdCTEGZ8Ox6LOF8hZNojMXEj0I/rmjNX3KQmV9nx8vhd1
UmwhExdR8sJXlyN3dKH231HcymU7v96vIKOO0Pl7sT2/dY2W8WqTl/mcKIYJhgj7
RKOFN7ljimn6fqbH6aCHaPlJtzmNiYvl/3SxprftBS1y/QPKFVnHtz7F5q7Nd3Cs
6TIq4H9/QIR91t44iMV+fseE3DWNDy0erF7faDn8Q5PV0dfqhcM+RwD1u18DDZ8F
uTnB2g31A090rZqkATmBP15x4XKRieDVBqH3KORHSil1OXBy+Oshf5q4ewM4vd/W
uMOGFlt7MhQXz+aVZlv7ajigbh/EsfKlTKcauetSLI6BrzPK3RJaYTWRIfwzxAmU
cAKk6wO85qwUo8wA4izFgSNPgSHsoEhEg3+G7J61R05fY84jcE+PzzDB8vZFqH5w
kNA49layt6QnHDCTc90/cC7izyNOqjYjy48Tr/CwdL7sq6c18EfFIVKU+z1iRjqL
f1R5+AVbSCjM0C6XutZKZn7SSdjU6E5NPC0Z5K4U8nCsKJkVXFdQQzFi0j5nJZoV
F8OslJMIfnMdmyqfc7d6yXWPcV55FzithNM29nfjbsel5j5xDsETMFNW/CetrM86
q2lYyIF6AFxHddi/87ITY/Noa8guaqNLmC/SViAwkLhRLbYZs7J5vLr4+/TxcbGW
dF6L30XbvovpUwcNXtAf7e0PUk7z1KTiJDLfP3oyBO4DRyua3pHZNE7MXDPXZQwY
1eenT+AEoook67QJETEp2/ybHbJ7wnmwJRBjVJ/zXpx/IkGTT78ySTAkZ+gJAZD1
6IWEBE9x0yzipTP4n0U6FVF0C4MmzBjGYT8txk9Auo/e0DI2+48jNjta6cc7fiRo
MS+SyCc18Zwp/8MAKwgy3YDglJ/ZPXxktm7s/Omup61VZrdXbCKwQUfohmuWT289
k7xlgG71fDw5/xlFztDqaeaG/EapEjmfUDBQiBuomLzJEpdBEB1ksbQgVPg3apQ4
V1wkDOLwa2nV6Mf1IdojUdV0Luz7zeq8DaEzJy34JH/VMYJTKxt+S1yK2EAsTNP/
2R9l5b/zn/5lqnAFpzrWDqDnjL+fpOzKjLc+bqbJ8qYfc6gqm3SD2zYxckN9GPuQ
WnRO6jqEkADVhY29OD980ZyUXeVmb3KelFR3XyheC8gcIND4H5kpGHeKhlMTU69i
T4fSNsHUV8NwgiobJpCbdejbjT2iqdjE6xys2pj8qKa93PTl9yD5/+OqgG47oLlr
fiAJ3d5s39XVY+Yd2QqvyGd0sRfPkifk/RxVFqsGqSUWib5z934EzeEaQxJqjBZV
6bExw8grou5i3MRrJIgi+ZMiDy8y96uQ2+y+8M02EhNiaufVF9fz5/vtFTpjkn6T
BfggijJ4I7+0HOxJH9vKD5nrXimEu7rvvmH5ZYWwgZZlK4oOKW8wT1LfAAbG54gY
Naqrvl7b9axdS+5hRXmTuTDNnHXDCUP4WeBfxMfq1ifNkpkXy/UR7LadaqDhk7kv
MSnoI7Pl/ekwcZACij4xJ+xNhd0NOb9nN5lct1wD3Xt0zQGVgQPuYEMeX9MHOol9
a+BFTUtium6RpgAkURdOahNaW/NHuEyG3pAITqLyqCrMG7f+6sSj3chXdrxeoLvf
cgUo7QYoUzzwDki6gB+GpabmMvIUR66CSalfRtJ51iVZy9NFhn46p3Q0bd94SEGH
CePMKGfJCpgkoIx4rVh9Na0fKr3FmR6/Ln+ZuzSnP0KRBMHdZ172+lMXxEQWPjCG
Y0hq3QUDFjrCQgm4HHwVzq9FQH9l+Xm6hbW6JQBogeDLZuU78YMdRpI+67MSPSNs
z3T2RA4puzOJUMpMvcfkp0roW9X7yQ9VzptPFmoJ04n3WRDn/5xs7/PPUEZkvmEe
RKD2pPmtOdisGFpyJPnPIL4GgwFf3sVxKHGifOOfQyZrcQto5wgDc1vmdMB7Zc95
Cuudn67DxPQPAXqpujCqXxwE995pjztSdTJTfKQA8YOzUvwzd2GoCQt+dGcIZDou
5G+ueM5wiLsHM/b5+8QeT2Gr70BIWbQUGkSnzSyHa2zKf7yDTmePUeELdFk5r3QT
RzMmcAFwMSwU3M/YNicvGrFRAZcNlwDDibP/xZO809djlxftHWZuF6fbswEcY+A9
5RViKTWB7GPT4eOAbNOd4RCQlwYf4qs2Q/5OCLJdXDidpQM4/sAzhA3EaWEvK++Q
uopOUNK0nC7Ojp8B7LsQOlHBpmBcL4GhxHqLRpho8G6mv+0dcs3ORf8DfWleXEUV
7yQPdZXAjqZUIPlCJeGnhODeKMn0WbAuq4FlJEXQoHIVbpwUZQ/VoE1hLJTtFCbT
qgg8ptSiRxrmoBhoFro1nVenirlhY6lNxUeOLd/2wutyKLguLvjnYr6BWdFvUgeE
fKVQvRl0qnxVxrbJLq/PeejRVwe9I8qZ7SmH88pRTMHtZfxx2gOc2sUOt2Q8BJWW
41WPAPieNYsJps+wrKUp3X5KqEdfgEgEJo+URo87P9PxwlzWL7/qWcnKRtsd0e8u
eNri/XTMsI6p3bN6o1oB6TPhTicqe8dDckuOMLUnxVaMMdiyLEu59X4UGEJScZwd
bx8Lgz5GrmdNjtdb37QZETeXY7LqdKMiz+EhFVNVbrQdRj5CTr3ibYNy7J0s/fgy
PGzPxl8k4wDYhgF+SHmPS8arEVzdnyfV6OlFR6A40bBNz7LEWVXyReuY2N1in+Ku
VmGn4P7WUQ9iBS6n3HJLHH6enN77NX5OD8a14yCKTH5pNRclBqkfmB0fWAR7O1fE
Dwdc8S/b/Nvn0oPIcXDsvtoakGW4rvo0MBsheyUwmt8UYBIvuWMLQkPRaIgJkEGr
B4Q4ZkyXUGYriWMGebIfLndTRnioZ61GWTRDHVEl4jGyb8N3m1eD20hJFipjSSrb
3xcR9/DPZUfCaFZHQFPhX5iqi8KWHXMkaFWwktr7tkTeKPHQRgHB8DM5ut4d41XK
QrupXtyLwBZJfDe18xW3BPnaPukFy4QJdWXaci9fEoFY2tzFj9CtJS/M06YMLABe
S665F98HnlOdVnnVEjSGwnQ25jiK9/NaiLDMnNF0UF+rlLb4/VYGbauQmkjoYWvi
f7pCDRHVJ0pBkIHty2r8HDiBSr3oBhC2LGVoseS1UXF3TCu8Zb5CiuZeLDR7VyhR
rjrLTujS4bxc5rpndKM1JwDWVKnh7oJTcmwX6+8YENRU/dP5hS/eCyXYKWO8yrWE
EBOsylkJdr+NGtbZevEc/43XYR407CDE7gFb6Wo3y7aAvBP70pp/lujA+Autz9fM
8zjBV/Le9pMarwUY3c7PWtkb2FuZfGQo1eme8IiQdPI59aX5aor27arAgphaBcUw
HJJLXqhuCGq2onE7ISIfHWUD67XG4frhq8JKdRYlAMbK1T43F1L+XjdDri2A/p2C
BoGXu5wHSKV5ExhpEWwSQXSAEI3pb1Zmjx/Ch6Ew103fIo1O+UtDWNqkCqaCnOpy
saTy/APtv4EnW5CjsPL6hpa3f4zued4ixXdHyEDzBZLoIKGMkEL0eZSI7CTNM2I0
tjqMkNrgvk/3z3uV5Urx2visEo4uFPf13rnW5sdWRg2tum9PzXg3q8AygsUsAeed
gCAJG94aE3S7CJUbhz5unR2DYy8l6Sr5O5mf87zmE6bzzZgt9fZi2A93ACr1DdEg
kWTSNVL+XQEvordoPcqv8pI9oKKnq+5Fd7iMSG1MRVM96IaPIqAfWIaHGlhR7zOH
Nn+V+C6Abwn3w9Yxs6bp2OUeFhmddRsOfgs0PFDyO2jtUAxVHAVkBvt6Wpa8cPkx
qAQaxea+0Rg0LgbwPNo1JyXysvaaronnMVbuR+alXIBbBXwen9xGIBw3XZdV4GnD
xqCZEjwl0DpHjOChPbGcizApjcT1IG+0JVAdOgjtIQ3ghjNHqUmroBTZJmC1sXI/
ngrthPFroWWVLkHW2zKQRTcia9QyIxw9VsHpG7NcEMiY1Cxvre0OYC5ILhF5REpT
175s3wRw/Hchl68JFyg2s8q1FXuow2T/AEE16N/i/6oqhrB5a90LXa8foSZhDY4G
AYtsZ6nLfjlxa4Cje9cqoGoX31BSNh9mw+9v3vPKme5USr7wEfS7GcBzgSJv8Gvg
ACSfDpEXfeqJ0TA4viZ8hS9vjeKzo+mMeWxAwRuE0eX+AZQA1EULHHyYIld/rgwy
DyLsE74P77K5PBySgay0tth0Kf02cRr1dk9jopVsH+wf0RAw+/+q6OE+EYoTuAsz
jPdp1r/BwLF1VpYPL8BB1ok8f1U++PLxES3ceSxYw8zBJA6khMnGmOiBGj2eYeDw
J8gA+BRnNZX7QQQ/2Aza4169aMyLTYDGWhuATyuSSpFjD14j7Dzu9P+Bkurf2uGf
XP6KS2Ugj/qtnhmVnawX8mXzaVj0D1u3UBIlCFYBHiA8MVqiisX+iDUt490lADEg
DMU1bEWP+I/mSP4HNq9NEHErPKD920VEa6RbGsztWcUNU4yUILGAZP/CutK4N3v3
YD4zvb1HBW4xiM/CCEVTkFomPCpFjWK8wclWKdJg1ABFGPFu+V5XCdTDLnkh3Uy4
qYNnIYgI/r/pKdEW31r2MkRkU1Edu0qmMEgKsAmX1LRy1uP5YGspS7SEF4Ci6amW
tQwXV9b7cxUraUjTfJMgbHudomr9p1UoZIGb0y3KMNLsKMBXGFCF3pDsyR9IWX9A
rYBGJVFMhS+mvVKQZdW2AtmA14r46zx1FGES9JPE7eP7/JyYYfkBcxJkkrOvK2P2
cfYXdjuu7MOuylhn8fEx/3sGBl60lziEQh7+EcemTa8ty6B4+Z37RLSMr+Bg6h9q
eyG4UvRDoiqgMqptfqikLy3m8kCb9vJVU/70t2B9lpL9f0RfQSVx7JaWJnS1+gvF
jNGvZOCL5y6NjOnHeUAERZ9UiWLH6pBeE/gO6Iu0tKMEEg7m0A7BAlh5G0DWfEUs
hy9ZDuBzapMY0eUMpXeEbzjUvakkl9hpx0yqLeyo44yzimtPL1ZFkxIBKdWkrKIe
lZPPzxd21dpvX1R9erEEr28k5Zss+kBNUeifc5nLJJg6/EpcyTanjXuKJS8MmaFW
h828IBjdpokAcSZdKh8Wj87atoxDwxOB+9aSvQxD5ZCFnst3JKbENdOocxAtTRP8
dUWmg/d+N/TEdPWxNZ+W8NBaof6sCW2flfxvIpq8PS3jbcwmJOrrn0GmUXhh1q4a
ubMK/G+qyA3XWxJP5+giikljygA1A6Y5cKdIRF/ACinvX/AE4qMYfZWykD0OT8sY
HFcDS1R+CdfdRjH/SDIRX1kTGIZ2IQFV1UCclR5qN3E2KN5Av0OzZ2K2uBMoRvs6
M/8v/gIbApEdldi3VxLoVnXRwHDlFto9PSJjbDod1tTUgH3ANwdeFpboUilz3cke
JdO3KsBby7yq834yWMlfXE+djGBcpqu7FR6aEopcqfUzHmLlXkJz/eCT1IXVnkfV
ice+xAagv2cu7F3neio16C0XdPVqL2Cmfpr97hocYrQXndjdtVCJwZIn4qq67SqF
ZgFrCHuavDAV8IUqANHZ800xSkMf9+B0auNmH52Y3w/vXUl7d+eJ8KsjEU6qPv/U
RnwoMEdYKtwbHzwS2+R1eJhfHvU2USL/3wGvsdSOwGR/6sb6DibyDYLyQC2CFsVn
EsSZ0FurEuQL9GcsWVm82jQL3w/lUoixTelj+2nNheLAGfBXMcxKgadrJwbtwwXx
kcEDCuhqmiD9acRXwjkDlckn/LFMNzYaR/EDXZa5lHasa9w+If0GpTqExRkoNrEE
Y48Wf04EynCKxVv4dZ/pVQbI6Jy0nRgv5dfPJSTthWhnGb35w5N1pGEgXN9L/mhO
/GNLAa3kjCVRLvI7WHyS39Gy83G3CT5LGXAg+XYvNwUj1CYfyOw4m9vL43GUPYb2
F6zdtv6mXmG8xLbYpJi5tEkZkUFeHZerIGtPh1QY2Bw2gJzMP1EucXxpbqpmtVnx
A0TLyKvve1Xqky0K8VR4FwWefhnwux8M3W4Jii/dtMINKIwVGOoH9OhlrwoPsZDl
0HgnQY+JpqZZ1rV1WtjKCXg9MU2BAnMlnvNmm6OxOimoy+dqEdzQYzp1F8WzUrr3
ZNASnM1dVOMyfaA9jTOQaFQ9emH5oOCXxaAGq8uUOSvF6TcEMK1mhNHLLpg9i1Ai
Jq661HDJmxTe9EHOBC54FbwC90CDeU7XFVsktSUNfbr5LTGOPWXzbaSXop+EeQ6v
b43TktsAqvli8b+roeipe6YdOct2jPb8B/11ZOKF3/O01fPqWWKV4IeGAYRfaioY
FMHVyb0NRpsrwKxGgIXqxOCcpsFwC7pmKE4BA26rSVEl48phstt+JDWsFMMCtSO0
4aXZqYRadDY+N7b8xwGJTMwyMVsrON7f2EBcQLuLp1Dq7SZVUSCiGdZdwNoHtL8y
APc+TUApaWVcd+5RomzzZ4ANSghs4/dl4UZa3RcP9inm9RZX9ZH7KiuLUUbZLtlR
diFyt9+tv1QY6UapHYgcoEx8btmHUzLq2wigM+3o67DzxMgknhE5QmtPhU24w9vs
axkwo9zx811cXDWwaX9O+pCw+2aZ775Dzysei4Sfo03iHmfRQmx8naBT/ppN2bGg
AC4kyNdcwFwA85krTRn0q3B+4xwIYUDkLfXz6N7SEymZ1cBf2ULdNAN3/hOMLCR/
LZCHdSIJxScvlbBlvQ4mhrWscs8J+vEkiFPA1oytwSuC9sHhw7PcxCADiccBDg8K
NIvvHeO5FjGTEE8o4sJKyLg2QOPj4CdEp40eC1NqCS2LSf4HAMAM1PBvs1NL7947
qRCJGn0mqpxNhpAGdzLgWY0RCSlKIi1IVxfM2prkP2jO9BM9l0YWTHSbSFfmKXCk
tAD0nSLvfitsveOPXW7KuVqwZBVJqpHkxdwY8L7tolvIxd5XFe9fxH2kpKo8Ab09
4YMgxtBJqIAfRMth4PfL8e6D70bzSqC8gONlkvbg/WrnDMPZRhd9e1kqs5Gh5QOD
TP1awT6dmGF+88xCeWlXgaq6eP+0Gg/MxMbkoZxaLkgSfKIt58u3fsykF8MuyO7F
ragunduqJUDDKwhoanTHlezQduGuiZ7mE5/eqwu7HGToRUrXeTObiGLOkzSfQYwD
u0cMtHk1afXEZb3QGsi3otph1cVeRpsLOjt1PChNRozw98Tu9FmE75stgbEyw3Jr
MAfSTe5+xr9+WF5HLQ3pJspkCA1rBi2MbF//qbG41EGpELVTM7TUar5lmOZFAQyE
ptFrfYNyBV++GmpWwIGn45zVhO9Jm2ax++oLh9nxyyKrFXBlNPfOMI0uEsC5vzLe
xrgeCE2Tbwy0oJlJ9N5b51KDK42nWBYT3evkPoedgQ5bmv/YwprNjWUqZIP2+Pfz
04rl8spwxEHmE38mFmCpVoXrHTgSAfvFDybGIago5RvYe8lCCIYdjig7ha6kHorT
dwc8M3gm9nz1b2F2pW5tuP3RZ505mYakUoJb11sFP1jMlWFCthigrb3AzGKdz2M7
HaWbl2eFztYvA66obMCt0dECnQWrklytVxmC/u5VfwN84bw8wa8XRTfbr5L74Pxq
vb41zrdSmrW2az9Rhm8UuoYUthNwvFsvwIY1j0+mhJKrE1CKGySjZdrpjuzpLPFA
aLsYaki24b8tVJaE7/WHrAEpBQHApjTt/y2/MguDZutO/jFrzNf3gRGNqJlbkYlE
E4SiTQLEGDD+FTvjK00A+ga8tZUSz6TqUGjOSzcIADCYiJ527h6+Zn6Bd8tjeq9W
hj1K5ivBxL5VvIZ0dACDkTScli/CMVISLJBiWgdrhKHxv1+Tf0AfVxARSZEgA6C6
VyfVk4H0b1lHbo5IGVF4Pq8fva3MLff8/pUaXPTwaTdkt6E3/woO+NKLAxl2lnb6
rjBOmND8lvYZhc8Labrq4vpUfAhml51DZ3z9hIL23eM9aw1T29NrwNvAzv1xMF4M
xNn2kCivtVns+FE0JD8BU6zn0zO+WzdnJ9NByGy7i8HrkI2a77f6qBCRcWi0t3Uo
ATc1LSu0AxwGTdHAa0bcrt0/0ugf4nQKFMUdK3bg8wvw0AWrDoVd4JjYx3ggPAe4
5lWZ58Vg3vbeBmbUBSzrP50G0gOoegMzvWS7vYf3peQGzRfda9ExjDfd27+Ln5ko
/kciV85LqfZ7Ga+2ai3DO2AKKjszSatlXnVr8utivEREfKoWPRkKeodZKC3O2aBg
DF43Y9dHnqwXenCLyhr5CRJXgQYTkNMbEZKBpP4ajCMKpvHa+8nVZXiPZ6TWTF2c
g6Jm93/wkc1PXI4nr+ez3hbUMcwHM4Z8BiZtvGfaEyCMil5zXRUzmgpWTpLINn1I
mQMjM8/fp5/mMOvmcWwOdYLFMrmZXwodOBr5LUhpx3rY2DZiN6xtQpo38NJKblXA
Ks70DsoAffa6Ru9O6o38ksymigYX7v1soTjHy6Z+p7gK2HSNw+otcxiMq6aHjBde
+Y47HVOabenVqTHDlPFBOTuSA3esXwcv4HlVCp8N/tSHJZ62U3pKLZ1zT1shlAsl
isVofGTu2AKiGsBoVxAHrJPxjoFLFl1H47w6h9dxhWZNwfW5qZWslmPpcoDkLNSz
TCOURi12T9nE4RlsAago0Tn8nWbpKdOQ1fhm8RhshKLlP1dqszBlnnHy3hoWFBio
0jgM6XiCzs8pCHyv7BcUz0R+Sc7enToliR5Ni5li+4P3gFrf8v0UgN/KyVcmURJW
C5SvS4zoPnWykiKpjtTQZknfgXs0jzTi8gljst/F6jmaBq5SoGwhxScNqP96BNMh
gwIemGVgkqZXVpSsso8294c04hxPbHSQEfNL8x2lK7lYIoCZL92wDTprbibdf+dN
LadJomlfFGn6CZCA6S2jL2gM3Sjz5aV6sxwLIUagk1OffFfAhTf6LTAsCM7ZVpI9
FuP/qvE902UafuLgtBI/QNWIvsvAIeC0qiD0LfR3eODvQi/yjp2Mtk5SMjf10vm1
XhZ1JzDXJ5MVlJXLA/45Ygb6/b2HDuCXm85cp6rfcOjEHBpOe/lbmEJoyi4z8NE3
uf0SMmorA/UtlUofh55Qipt2Bn9X8vKYCjOdpvJPtSy+sQPJU5XmK3lWm8WSZzVj
3fhwl0LsZZohrDiqwBS7I+Wri7asJusfIW3XJZlY/hAVqNHDBxhlIYQ83Eh3B+mA
RBBcvoXCjE4ZFiohgUk4x3JWRZaeZotS0JvEhniOP1anAj+o5OgbGzsIi1n4YFo/
dccjQtDrscdQKNuqA72ce2WR0yIamHiQMPHraG2Uv0ULvosn0g5d8cjDcaDKe3vS
f1K6pcV8tXOg0KbQSSmxjXYdwGsC+a6HYtvIhhWr8e7IycqNnYgOVofSvgbP0tj9
6kzc8J+hQGJKmlb7O0WZLwWOsuoYn0GfrT1zKRk/zoGFgR0LLbmyyJx4IyuFK2sp
qxRHAGqMf2ywvC1hldM5lqGCpaRFlaEbSXHVMrf4iXIVTi3j5C9qN/nR9t0Uwyp5
LdKMNrctCrRb3ZTTQfCRSkt8YULrrk80TCU67gb+vnu9qYpplRdWvQidia0tSXGh
b5qLW0gJUA1DvR6Iea/M5YXlydwalRGSiQP3CMoPTl9Yjxx4QlQJ8IpG/r1Te92L
Jz0CYXSdHvffZDq7WR/z+/5IQ4egqtFNt0t8XKQiJqBUwdevZPqZpP8Jgo295K+I
kXD7/a8tYFHUniLt10Mw367bIbDHprSuZyDPc2s4myEqnlK55LwdiMVB2BZ2Rr9T
omptMtqc7tBb6K8RwrG0vKgIVq3IE7sWxB6ny7mhBWcZnyXqnhBqnu3r/Emdlrge
fzwvhzko6ezgiVjw/bqm8Ayux2R2xxP++C0kxiF3fnnuoCYlKj7OOymXWYAsJrtC
0CXqHMnTEjnobVRXYubgsc16cyxs1gYrTMvtWi1ByMhCC7VOLV7jEagSArrA8je9
WNi3lLd742WMJJzrakBXJr0XddbOEuAi3LnsgHy/NSSFF60Im7QF46xBR2EPojBS
K+9M+zz+saFFBTTJ4g9ha0hXlnZfTAlFELD7uZxJlwjegn5th2hBARXYVaAXRCf6
XiqQUJsaefDLeeZZZWTnFZb+UpD8fx8xjy0On8/9w7OKWz/PFjXoSm20C0snCZpV
rpoujDG306rG26+FBO8Wam/fp5gCeSdJK7EiBVfV1stM3+tyXi/hNihNXy4Hpq3a
7EGUoBO3LC3kExwG2juZJ0Sd8OX4kntbK3CZAkDv5RUZkyLzY4seYMesPTO/5lx8
GEzU04veCLQz4rMjb/mznlaEa5XSZxaBHGk/E7Z9X5TeZEfKO0+ztkoZb2Uszldy
vk4rqsZbGNdlwYDvK0bWyD8SSjMGJtxxKnGlYR0OXJ8LwWgjfszyH/h8XT20yePH
HX0Zt3TdKuh9CqWYnygZgqw5HUjBK33JxvAvBRJVcTeL8L4PArBTs315Keotb8ie
jP8hk20NxaIiNoyIxc8pvOFUlfd0gwZvT4nTi/ZoxlgG91dVPs7GzIJ7oCslamXi
7Cnql1xYqKJHcolKY+bqv0ZILuPBG85Rs6IEin9xxqxGFSkx4L8RagMZSLqU+Vt+
WmAqUbV5WyPzXSAXWi0Zow6CTxLP9pSjot4VKA+zP+K/bwyxAzUzA2XX4p84k3Zn
Ie58E9lMqWx9lI/8NOQGlHEAZkhMRxrXZOkAzfcD1OiGKMKdVI/sBpJes37pkhB/
LNzQLB76HlEQJvWCryRYxr93+Y4zXfDIimCPTxqqklOjklhZyuv1MHu1YqfWDENy
dgYl219bjccEGGELseug3BRegJbIfD2m/hGGguu06sa98c1TUv1g4zsIf4lrzTEq
W2uBDl12gjJxcegIUfH9N3y1JhrHlvqZsyZUmDgTu7WLYDU+7s+h3TgFlC92JH5i
13raHN7hgFDXsr5K7Sc6ZP6ROiPBP0OT2tFUa2nb29RYoLajlspQJvKB3nrcvKYz
4El0ZK87WPZ43IvxZul3wSSxW0qIo1mUwNZwqn2bHCobVfviXhS560hdKGeKreJ1
NMd20SA+gY6ErFzUgagASJK75E+9lN4o4Mh412kMcz5H+daqHPhmuqkYdyoYYJQ7
pXvRTeseewZjUyNnw//w/NQJ2l4rvZriFmFrm8FuZtxJW8FARV5RvleNsTynmnuB
szP+X/4cpjPkn4TttWnoF18n0r5DOQq3qhrKdcmMoZXQ6MlRCXwICXtE/KTZOGsz
q6DroWoxInjWWODsw9TWUY7hBLLDLMQE5++HrJKe8bEWwam7QlO+bQfSUdQTdyvM
bXJtanosO1daFK+VSZFAi3U8DfrQqDApd2vUCcxvGSzPCwMp12/RaKGduUBfn0F/
fF0sr8jqb+rL40Ff/JWnjN/5pzsuG/rKELVF+FZ0MyKmaCGjol47z/BI3ru3YmBk
Jvucm7Z8NxMeJoVeWlQ9/DYblWkhGJ+u0fB8s7QG0syo9BEu0NlX3YC2esUPEEOA
rV9siH57C1COtKQZaKkU5oMzw0uIpiJnL03ZsuSsx8JfZ6HOsJVWWVQFJV0TJna6
ed1zeFDzIfIGKD3WgXpcMXqYXSRdk8ENVep+66wMGmqzAMPSm2p6X0Ho2ObB4Cg4
3t1nytzh7mQI+n8Lf3pV8LOUCXdNn5rFNDOe930dRFNZbR+r1ZZlqsr/GvHf1hfr
hs0mgpEhF9MwNlE7/A7c+i6+OuRf3u/NPMR2bBPJfQsn6XtwzSCjUmsxXEs5VeIU
3kfEN+uO5F5IlHRJPrqrZdUpep0rlpfw+hVukK3R667UDTBAGu1PI4XdWYngXPbf
d8Hk7czW4VQfIu6mg5JhL6PTOj04f4W5JzFL2WOAkrpn+4p49XsXwj9Qey8/pLYq
cyStqLcnfqb+HmbhwDMCmAf3+3/vQeO9VBYjq7/uaXSx0XshwIpbzmAYcbZV9Iwv
dh/VXFhFHKwoRons76dFwU+tRVErKSBFTXfaacB/6AiAKx1m3oqkzsod1nY2OvhJ
CMDpA18LDDho+rde1+BYGepGh8lsXMguqO5oR0kdWUuSJ0+dHRQGJsjhOa2zlH+j
pJ7teNUdNgnCR7oQwzClCL/pNVMgeKDL4At68mJ89sufKwdqbxSmfI9h/TubEkKE
O+V86642grRTCv7deqepngPzotgwFlZgXH/qh3dgelI/Qs5IDmwHWnWWzKAFU1h7
tBvRNZ0MSPTnOjF73d4F98kcUY8XDMSdHK4Ufvohog/XanM+0wJJEbXXghXNV+ur
FFS0cwsyoCffCQ5ro/E5BzRIPxI8FCuE2GXi8VAwMGA20GTLN0OaDyN8Utx6pYLH
hb9rskuXXZ1x/a2f8IonX8aibiNPDH/qYSgE72dF6CceAyvFbx4eW/QTx3I/qZKz
aJJ0hKnKOkRqs17pKhTw5E9Vw8uIGBsFyBjblETuzGesQan//+RkfNWruY7S4yI8
6i/u+0Efx1AwDOukLhgPvI8d4OLzfcnbK7hoJrfG1SpYr7EFidbjofozolEtBI4Q
ZpETXdhXVd/UTSrVRMWgReQykEKxLmhVE+4BKCGKLtm4hj59yRkKWvuRXe7lY0QE
51IN0JWe4mcNUW8jsEwgeOt2Q/jleshAlhwJJEu3alTNNdpqJPR66YKevKEEmtlc
wexe8bekQsv5bPAeueiQgKWOyTmrBJAncM6csOEOfDpF5WT6FbOLHcE32bgPbpwa
eeOC/NNdP/6ecsVX/gzoZ8swHQSZCRNsmgOdIdsH154M7S4Ad7D+DIbDYfZwjc4Q
SbM3gVwImoZEuGh3DnbHHaSwwXzhGauA51nkfLQXuA0vOU85VEmlCt8uYE1GjgOh
zTDhD0X0QhLLh/0dZR7QvubKBLCIbSTXWgNk5uOuXw6XSJDS9+QTu7XnUb0sc+s6
Kl4PpHoMyyPJgKuz0MiGVaMBMLBOuZSZMhYEpZO33irnK73hkkJ8dNLP4HZJgVfc
BEPjoNkeG7I+9nmQWNZ3Tzb+AK/StBE+iKQWOwPM++quzUCnxYcw0YhKfc3TB1QI
OofMNIz5TswMRXacftGzwoIVjANq+xJDo2d001gtZY9vBQiRooWxJDsqc0NLHMzN
DuiNkCIVCL5fxacQ2/nbCGg/60XmklhuuIlOz/Z7oUVnSQHStgtgeHL3BUdbjZTp
T1/AnmfdEoX6Y5xbj/oVDdlQ0XuYVvgP2z8W24KxEfIvvx03/IWc0xA1eXCDjcN+
7djECo2cEV52564V3UNGb1+95t3EJ2s4SPrf2b/9EomylRtV8DShVCvgQOjms5RQ
6CfVY9hDMo2Vba4bZvcrNzsIz8cnEN6NklZr2wVQDvEoe8BQ8uZz5PMSNaaSVLwC
c3HSKk6wckkFU93naVJrNbp0FNwDgqWOTA4mluvL6lE5gcPa+Xgiji/qUdQaHzrA
GmtSIQdj9PxhaAGPzzIz4lg/2OdEhDRo6c9v4EqJciPH1lN9Qtuwiel+gBEdJAsH
jl4KTNUYdYcApTen/rsEma08zrx/MJ6QdWjLahlMLNro45Gtj0WGkx2jNaUnI2OA
KNpbM/lJp/fNUbP/baC7Y+n1I1S3SszpvMQvBnq6efdp99X/V/FlE6GpGw3IOPYp
tsRafxvCDyuid1H50Jo+ASrVkW38xU0uhgN05cTW66b6fyHBfDgK0XaVuFWzI2m3
q+j6ZH9VnQ7pjt18x1OM1BiNPM0sxdERU1wsSYXg66U3U3/xBDB6//XDSNGCPd7r
k9m7+dBMtb0wlc9WTBI6SGAgpq9tWCG+cRqY2TsflldwB9t0nT6d1YynICOPj+6J
J/ysYPTXf94VBiaFVa+1inZx47ed37pEJ5mtb79J+BF47rOPYEs/+SAOosOAVvNc
URew79hUg1jCBJY3dw5Bx0wjkZp6Y6DbU7jMkL7XFJaCngz/tcZy9XSZFOUJtbPs
LTHP5tDg+5L0hSvw2DhDBB794xLvOabygfUE/GdXvJ8jhULscyOzlznV/FM07ZbT
5Fhjbk5LMAyZUmaxaafdrV2JX2HckxPNsiuaQVb5BAV12TToMBQ0wsdiRbpbbWNE
gcv2Inr0iIq3EtTwfX3vO8ksrYaBKyUiQjz8/tdw9/+P5Gwzw4vK07d0n0bn8O4g
o1d3IcmSZrLDDHrlnMDTvWYF0iT1uGD7nJgbvYbYaZPg7QLAce2OW7O/+ibVA4Ra
qA8T8LcDvRhvIJ9jRIDUfhKfgtRb/U4LKndpMismKaJI3QHxi3Zg0q5f9E+Y/RBJ
ESaoOz5SD5bPq41F4vc2hmOcB6LYknxKKRn9IzS9w1pWSgpdsFHfLap06w4Iqk9i
7GmscTKhfNH7Mr1BUN2i3lk4kSZs606VXroWcP8AyOUG47xGWpnfyuMt+MonmhR3
U45fQi1qsfR/Qr1yKKI76cgjF7EfIEPpd7iYZXbI6+LLQNDpT3a/QKM7zDz1ascn
Gy9ZQEvfkSN4rwl5r9PUGhObJC5fmh/HDEwqO0v27gprbafmWvVSbFj0XIJIBhib
tEiL9cuZ+bVvfWALVdg9qolCN30GY3MNNGjOB/gfrx3hK9vw9Y+OP0kXvCt/IVpp
7/db8Ptb/PA5sw8eI9a8ESlQnzYhcvAGa2ordG/XigQ+l9NEMiGOQen4qVqfx/O8
hGhA9+LkQ6YrhsfgIQG5yMSTjO7/j5+d18tI4ivgBe1mHGp4EaXXSKW5hHxv02MV
wdhOZ73gJAHGA06Atmmqu80smelGWz33J6bgx9oxyceA1d7F70ZJtyA9Brtl4Cqy
ksLCXFJARa4VeLch9peAR3/u+A6jyH505hfuensDDbDVGNuqnfYiL9F7QK3G2Bk9
j64/nkztbkf7gTKqcjf+OxiqPyj72k2R4R/Yis6KGzrAMjzkOzcwpzfvLQxNHfc3
udYdYQP3QoF4MhKJ9lxSmBK36UT0tPHgifSA+eG0/7VDNuuM+avZFR4kkS+8GQHY
EgAQmRtDlyk3iMB2nbi/fQ9MTImNisob61jh0otT2Eu7oHu7HxY+d9mJPgO6pXJI
gaQTl6IfcaW0WARKzqU7hLnzi/fBmnfLnI9fjehneSW9TagVL2Og0NHCretuJPWf
YEC+bGWZrv11XcM0h4KD9MjcFjjJJbOvDnXo6CnQrxDFIW2IQz5TXw182wwwYFP0
XeYokKLZm/toyKfymvKwB5nJu3rn812TysTz9TEq6qckztKXXJtzWeXaGoDEB9Sh
iPBPtEXsz6wXs2Tu1Q2tu0Kz+7OCvQzIXtw2C0xBjcB8eXx2p9jQwdXzBOLaRR3+
xLHhzuTNEN2g5LzvaaM6dLUfIcVKIsXIyjNaft8mDqsMyvVJcDthjusqN+vbk9/C
Q2OQ9IS+/mQ5cFa00XjhaMmFNsIRg0H9N8OqB/GF8+sNr4wb0ERIsRtYMdbSHtBi
rB4zzFruz2W0ON+b1JLT56CRb30mihGwDYN5hu6t4fYBBkHUh2cVRY0tDkyY5B7L
9aeXwnCjMPZY1i+YHorcLgytlM6I0F/S84oOyWjqNCE5kjOge8mFVdDGB0iKUIc8
AMXpB4Oua6+Gu+/Vgn3SoUD7s/6jSM5VOAQKi4p8zxNuFqYNJXZZTpLA6WhGitx5
5kOd30MXjgag3eZUwMnN2a/HG383QPhRqEBMjPiMR9//jFvsiiWyCMjw83l4qzBF
SZOXqG8IlOpIbuIu+QiX/UyFusAyuyuh8IEA3l2Hp7bolNgeoDvJzUbnTZbctOum
lW/x1a6vBBIAb4NfN5HvnY+wvwEA4JISxND+sUhj8Ycf/mVYJHhJO/tgiwGm2Iib
sotPIR/6xX9PwpERh+Izk1vfrmk4CMWSr0oAErH4lUbcWRimzu2kjsqWKRaCV52/
dyfeEtPb2SWqT/nwulgACwDpev0quse+HQbUVivy30sKnGPzQ5Yljdj228zjut4d
Zch2Tp0LT0kJl74bhxHA+Cm0D5zCJPTKApR/wDD9IU4YKHPnDwyU8S2wrKCtLIwe
U2DL/yXugLb/hzi6pgwtw2K8Z9WE4Y/1JJsdJ8neKF5czY2Aom84/6QDQQIH2Jft
xUlumV8HXFOmFHCEqRg4Op0Sc4cRNe6Pt9FuuFOzhaQtXOcvG9ivVe485CBBte5O
OF++SQOhYR1csfxtTRHrqYPhWSKsoXHzfzUNDphYxAtLTmFV7fpwzk/R8qNCRkjj
EUxygeb+1iAKcz4tmHmuIduxuHxAk9OglNM3uI9cx0cPZSZljAwDHL+EIDYaOlHl
Rjn4x6qutfoH5jWY8ru2BMsxwPPtsZVUFU1BeB7ByuOP/XpqCi6ECd2VwfabW9qM
V8MFucIgicmhbZ8tRtLQS8sLzknwNRNKJBRY5QYBMNn8K2a6HXd3O5ydQh8Yiz+p
Zvc7Clvu/qdgq3n5mR4BKfWXNKxVzhZNizTu5CQ57CcXCnzJ39BaDMBS8fgvKsA7
RFTbr4p1147dU5f4kDvE22WZHRfIHl8JXhSEDI2RyRY/pE/y3jrOVM4MMnIggjKL
yGwXTiap5OWMiUdKuZICzJnA6f677LQoCb7qNHy/9d1bkJAuPYGypDfywFYhNqUR
S6JALbLmC66NgAQ1wlROJ4dUxJy3Jbc33aqPL8oDRfo=

`pragma protect end_protected
