// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
tUf/GElvlm2hE6NT/KCduBxoUNQFpaupvLgg1+n4F0rwDCsCkWDzN3pAeg/Tqmid
+ha3WxVJ4fqjMTuLsD1UVCvh8SN3jmCusGAdIxOIJfLlVXHTvI7v7b1HgmUJT2hj
vUmdm5hY8L2gaVA7DBVoL6sHLW5ghppd1ZmUZZ5h9cE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10848 )
`pragma protect data_block
wA1w+4U6ppUuZJ1RdGJKR+gc64q1PUyILbJkCnF63hlW49e4G3G3Q7OuI/w039VQ
As1ZC6fyg8qZHwgqq+PMqnRREINQz366TDK1iYlv0YgxhpTjpzTc1EUoHScl0sq9
EfLYV5suSn8gSJ3OsUT6siAzL/TcNaEtCAimC69EKPbVnDqrJiuKKPaEpWW8GzfH
2AqlngfSvUUgNvZBtYGKjxqzwTGTIjTJslCswFXrxHOq3Wt7+PaSMJ82ehPgyQSM
SJvPsbnNaDbyHNo+rS0AEeeGDN2RYWvD8N94E9h1TxwMn2/EVSt1RTwgY/S4jVXs
3e4GEyIdTzL+EMlDI2ZfrsI0D3QyPlt4cmDZ1ZK4CU5by0BGrGmoUQxdda1a2VIo
Tb4rFf0CbkiZKNDkdOLgHYNOgSFmA7jz50CKOmH6DDLloTqxZ6v3dSh7oD6dkQ6x
QAVucJWx5e/m2ZfiwBiQbuCqGQ0bAJj11VX/CmeVsc2CvfQemUcZXzZ6odK93qna
oZm2I6NPv/JKKcpm1qItORYYvHUfI1MTGYHSsvuQX0GPgt/Hp/R4ETLNmTOAYF1e
Obu9/++ElVsCytkwH5JWRFZAIoSmnn4Ouwh5aAI+SXbv+lfhuM25vZ6nuN6twtI+
tdWtZOjhZ30o5+SZ+GXGnBgmeH0o1BukRFUG6IXwXZpmBUBeVguPwYn/muDYYGXl
CzKnAmNozl+uRQEuQ4OaF7J8urjJRe1jov7/27rkFkffoDMUQmpn9rvoNIZzMlgf
eCapv6Ek9XrZlSdROFJhHato5wF/EVp5HYTiOnWvS+dsAKFkI2H4kmuDYIe6dLvq
mq4bjgwKZ92gcKkL8uSoH/SnsaBmUGZtQQwbzuDPVvLMIOsV98KtQBVVLt1ATLhX
ghTKMjPVrQL6c5j5OtfonYgGU9TjhSQsZroRgTqJOS8gUsg8wjL/Pt0hl6TXw/UV
LCQvF7OWqypxeSJMLkv4dAWLYRHlDd0n4JSmXzByy/yBUDZSsr6j/lZt6njHQMIO
GFyfc93EYmzL2G0tN8XlvDkpnO3OHJ8IftKrFTu+e6pYwDxFTo96ZY7KnBtkFm0E
u3mr+NHszWbdYkbg1O+2V7wA7LD/JYajccVfnYWwdjgKu7IsCGjkNOsIEFS+JhkJ
GfJKCNBQYrFK8DPY0Lks9SIN715IyHbeeU38enVD8ZNUIT2r1I9ZTBaTwGy9wWLE
20s4x5rC22mHDaOHeFMl+NJ7SVPBVAfaw3QCWiSpxMlSihUmq/UuCUXr++1l+UQb
wH0axHV4j3foaE1B5zs9yS3nvNbSwrEgyQUUeAQLhLV4/ojNREuhU7jkJM69QxkY
JZcrSZnzivrCRVh6i4nhBqmilR089D4bbabivZaJMnhvHlYDhFZW8Jg7/wmGXbNb
XMpNRayx+bQ3/uDlMNF8ePnZYZAJq46Hf/xTLWZLbRV8WA+k0w5juidp1KgWaZcj
yWHPcZ2OR+RHodC/X57zCdBRH8r9WbR6L3oRqn6uScbamwuaHadjS0cpyo2Vm2FV
IWCh9Ndp7dC8GsFCWAVugK2/fQv6GWur1QyCl/3uZucoTldfCv4IUHoLRHcesV/V
XU1SDkcfdAHktJJjUCQ/dRA7xFhUFRkl1p6P8xUHB2CY/khtFs/CBBzPSeWzOHht
/FpY7xmBUJYwZ8RX9V/A09MfYkOrr09L6HW1uc0WKET5A4GZe/6dINYpn3OPrKbn
5nRPo9e4sHytkCbJxWrTvQgMz/zfG42G06+3gTVGkN+y9sXbszKNWNulsNfEcIrR
4wQNwA5r/BpApIRiyBuNFe/aTer/lkflIdmPBySIq+qQ3JehCbj6QdYCbaLdnPUd
2shWasKtfQp0cCxIChfaU3t84kcs7Yd5fPV+b4rlNgGr/7P9saK6ojOnqnL2aaNs
0vUerXH1vj/9GiBj4M0hdL7lyojNv4dJJn9S9Nlh+fzvbY6XIEDiSoso1a/1lGgL
pc7BP+5BafozbuEfq0klN6/xcHKDGiI3utzRnzhB4OYLQwDsPfAYYtZf5iDEcJ3i
HQN3mlpC+6fRXjFvdCmF2+E1fM74mMqKhApgI93n48zA/gt+HSnE51QzCrCcRD++
QNNjZdnYxVT2K1zUxQUHKOnaItW27eYp8ZxTK/5A8l75ytImNGDRhFzila+3z/mb
k6SiLBDqLUr6IjAT+G/KY6z2Pipsqecxl0ls4CvfbKUllTGau7s0P0pRybUaQd5+
uzFSg1qKe1tA/oxKh78/xJ2a5goLaAFfoZqYPBhUbu8q8wRSb0YaUjzM7SzmoR8s
SUK/3rtbaJ3xo5RbZavUx915T3Ynq73mm6xsAK0D6iIjkdxY9bU/ZZQzw5NVK720
WCv+rsnPv9Zi5wYSVL1eeS5yzqxTEvTu/aCVgfJzaKCdGm4fr+zLhkJIoc9iLtur
PqidmrSFSYmXTS3f7F+O7+lo9QngoSkJpuewUcG6mKjyWRVoR6TSCfRlK5GvrOL1
4VQcdZIhVaZFrC+V2emE1qnM6/mTH+ksUUi9dYTyZMIGNUVhOv+/EdTTQQKW2zo5
HyG8Tdenhbf4/zf7ULuxh9bvZgot+Jxd5dcLUUQ8GxzlK55LwIzdDHVBnUnUGl+j
97VW9WQXcW5skzKZNpKIQZV/aN0bXo7DYcJjQ8ht7pLGCvAOsU9NkDDsc2RSnl91
FYIsWdInmZkd6zjdgRrmQL/9Gen3kZnGuSwUyXsS3OKwmFZxAWVXDAHKGUwfA+PP
bOSwgGqeQDXN518hkMAwrQ40cqRfKSm8XpF2Vnfpk8F/AO51QuHvixhybyGFfw3+
tz14vZ1fthoouF8XShqz8rd0GBuD60zSdhe5LKhnbgFKnM2IoT82FbGXx2r4L6xT
vgC+87VsU9c3TMIuIg9oEOjsL34GE2wFGRVg61X4Gi8GsFt6lyckpnxRt7l2RtF6
w5z+wVx5O1MiWb3IUZFyElf96xBAUmTiT2pll6zRQ6PliWu927NsWZzfMlNw6MYL
8yNGOIJ22OaBSxiylQgM6CianycEK1bn7Txmt6BqJ/uFSkBxWvPO7c2v5f2siak4
ZjSF6+lE3lkd/XzQDRF575ipzwU10KQEYH4jlm33tNtAPsYQGKY3A5ZQmeJG+/ss
cvDilJFQW6gcOLXmYSkMJUOIXZ7eFozKSzHs+wrHZrxo1LaA+xhOrSfhwSAzkJ3J
qcaqeU/bgwsg/KQQp/9ZU8mkF/1QPZkD/+fD3/CxtSB6b19xxR+MR4Y0oiHBDS/b
G2+b73A+JosUa2tFw8/+X95zP3LTIG6rseGC3Onw45GegUtFwOrIBHCgdrIVCiH7
a6+/9EqPdTSW85G0G0/m1+vXkxjDRlvxMrw4lj2MrKfh0xU9RwmHBn/OfJNdqaYJ
QCzymiR2jcBx4Vak7NZ6gGXyqgbvKH/bdECKM7UHkGJxRPhCqqhkqDbSEM3ZpgXv
5ZhXUmJvkNXrjDP2qlDHMRpe/QT4oln/zqXKuX4pZ13bfELnjr2+WZfAMDA87hLv
CKpXGqX8cccnme+LNX8raNPR1Htn6/PrPLqetBw/3UQCa6fTr9htQJ9CKkgk8bzS
yMcBh8NFcHjzSx2Yp89X2xTWUnYpdVqU2ZIO1+n07c50TXdCqNJjq+niRLjk6SIp
L3Cm/D6+ddcfOI63K9OSbQE1wpxAg47JOQPe83Eaf9H9l+Q/4DKncZjFh5pYvK2Y
obZsqakihMFGYfa/6UphtKNrR7uIdvQ1VLhlWyo4Z/CBSdJjU3lwzq2BD2WMRz4K
ec1dIqzZYGIE94vZq7y3wkCFaXBhjkHiOd3mIhkeLfUb3YPCt1LXb8ow5i3EEpw3
E550qmTwPlRDBenOMzuzj+CFC2balSJgKM9S3rYq+f7dILY2nI594miCH77M9Ofv
kgCbGZuoJV99wGEV+hukE22Wj/z9h2Uh4rZ695NQhMNQICdHYZ9NY9nMRfzgAihx
nex3ddVT/Aav4QWFTFgqPN/OdvlmQQ0a5Yp8aJVi3M0FEZ7bVQQ5d06WhhFraxCR
y8r9ArrNYa69FFZ5uamLZIhSgAVnNmU5aKgXuSUgA/L2LrihSTLsfeO5DoJ2VCsN
glPY9oX05Upnx68NMjzbNpH0C1RQDXsjySGoSgKNm0lqd0v/WBv6cHHkP65HAzk1
kc0C3vsTtS40wk4HRw2cO8daZJxe/+nTPj2/7kDpZM2HnNm347+0ETmpTKc3to6N
rMdRBlyKeYoSKiWTBMW7a5KDmK+nWdQYEwrxLJgk9EcLYITXrqMuVXWZg3MugPoL
aBxj09y8ltHRS08QW07rZ0IMdyCIYfkL/34fxm93sElQ7ChTy+V3/SocAu1k6S9e
ytps44QJaOSHLPmTkbxjx4csSY4KsS8Qanbi8Mn3C0rBLOOC/x1rvy4HhWdkUw4n
8g5irsSACbFccBxXhTkKpNYVS8qGqjzdidc+oeixfqVowRXLFcFKO4hQVtWh77i7
PG9vXBe+T9WT9qV4+0m2yRzkEAkQIv1qT+WtbPo4tUVydzPucSdENm7XdCOP3Fv9
vgD96qsMGL7D9YINPDx3u/UEfKedwdlRKHQ11zmklYqrUCvXkbpJo6JUGG53Mqmh
KfNVprzDo1ylVvunTHNayhcoYZgLlf8EGGK2dP7feTPfO99Nxdo9cduzBUOoJ4xF
ivZB0zKS0npUDhuJ2Ayhzn5hAn2NXpjfSHlF/vt33qFoIbqzoM+/TeuLPnvwNabf
1nq5iBa5IrP6ViUHOI0PGuNloyHehJagNRhOY5QcXj1hcH2LV0gKUGB2zGLEqy/d
n/treUdyxfA0K6IhCsPmwWdLNM4d5IVKTk1YifFmcz7fL86lexe+mDxcEIvwzXpc
BkrcW/Fy2uQEXG3wPGAvLCX6GDW20ez3H1Ywp/6eRDdTGpSVgZgCpNI/GqhZs7j8
tvtpbH5SKwN1sNDdofQ6VsDilwrF9X5dwDrOzG2ciijZMQloeoyvZ318wTAsiV2Q
JsBFodSIEsqnBO18ypLB/upEyraKp865J0o+FccZMpABITp/yQitOi7/Io20b+k0
3PUu0+VmU+FHyVgikdHzN9AU4n72zkUcK5Lnchq8nhILuDY18Knllogh9GDhTsl7
A/aYT0lz0YHsC5rzOU4xAPIT9otLEwzAv2EJTN5PNKsxY3ZV2kY2pFy8JffgWduy
MIEpTXIx/U7ynP5qs9LFh8YzMpAlbBhbSthjnSZzGqOX0DKU7EGnP3OyIQ4Fq4ER
IG0PDrd6PH7irP1Q9bMx21sCgAIYRVtEQdkaSA3YyTlWYmAPgdU1smxTGXfdgEnB
LCpxfyrLROdNM6tYp3Od26WvnSFcJ9LNevZttgbU6QD2XPNi0Ux37yHKjgXQfUVk
dtaLkYB1imGSbJu/2xm6LDZKrWNVCqdRbGlW+WbG+W1BbYM6aZp7HOQt7COLMJW5
Av5ugBBDfs7JKM4ibFIVRdQ5XLeAK52Ji7XG9FR+Wl82ztAuXVwEPurQeStqXhIk
A89XrBcY6x+egcHbV8cluGNVPj4RhVLVUv0HBKzVNeNwNq/rmZ3UdUgqImBLxZ+o
VJfpM9sXwV74x+afcNtaVV7oR5peM5FQiny5e3wx3jn6MHaHvljTbOZOo42PQMa2
GzG/kpSfxHBYUIfbSUE+8eyKeSjERc14/zOOsTGCkYbXOGXXrhUw8MxqWrpGt4I1
S9eEA5IjOBbzgkKjZa/4FeoFo5hpDR4G5u/zSuLmFI1kajqHO7QiRG2Bpxd286OB
Gdk81yR89hBdfp6ROoe7hP76eyKI1Bkp8jao/j5hIxP39ypxxQLdPcXk6iqU0kEl
+fnWJRCjucjkGqfWatvJylpZ5W3rTeyv0QfqsMXRu9tdyzGPPs7T0Uc404eI0zWD
ABN7hDdOQ86M4tIqntAiOJbIaPk+xH8JpBDpCBwRQAGo9NrF9CQbgAyoQ/YSFusv
9ubO1YoTuP4DVmi/BzvOQXNIk/UI+2WrTPO/PyI50d7pT4FQHaP/E2pTsdlWAV/M
9LsyAHuN9ZTk36+0rq2aRn4dXjq5cWAYVxjw+QJnMz/VE19Fzktu3Zybveh73ccY
x1B+Bsp3cHguAZY5C2xAg6slSoh8i4GsudksOXW6H4QBkjqgAZU7oNvXXfE2lJDf
X+dQGKuouDq6IQfry14Qh9S/yKTv3/VJtugJiG0g72ByvSblIePkxgh84r1f/PFk
ExyvYgBspTCkg0a+VAn96K/SeqHru20YgfB7ypGCzqHB+5N2Z8fZJIrDNMXf6NDk
9iNneYqysE/WngnI/HbuWWHBQFnA+ArJah+PaujOvRYPU91U0Jx1l45y3uyZASrs
ZBYyHDEl9TBCZPolgTFIpDG1HxT5+UI3rF6ebJ7U4jOMFJxSPI4nbzevjeRmls+9
uVC84zFDUG534nnPJdKoJQq5yyWzgQEoc2DgTiDlrymv3HiEqDecSf/gbr2ySqX1
ZQujmTh/IdWfs16VoTGQI9oT0yT9jjiNf/iwWv2qpwwW520JiGHY0t3QEz9c/Jde
u8EiAtmQMopG2ffuDiVjk1pXVfTT2kHlSlOZmdi6r9U4tY8TAOVPLDP94yl+b31Q
xY8vfAPb8oI+ddbtB4/vyRPtkd0beQfZNSL4tlXB3sfHbgHV7RFIvJDfaOhFuUrw
qWcHSwQrnC/wdaj0rGOAHLXJp44lnAQWXeUXIQJu01Pijf5dcdICa51UIwqz3afK
zO+O01B49mFDSB+UxQ++TMRM8+7W/baCbsQw9SbwxWQFFW2DuL6yaEoogLeyDQRW
yS4RXyQlxuFcxtCFe+ghGj59wi0jM2mUdjAUW0NCDzbIrnQgKMNZFxWHSPCjU5fT
nIMXP4bp+Id11dDHa8EKae9g+5g6j7RETZPAUDs5HavbCihXlkQp+Ao+EVa0JGz+
Lrpcw+4CBCiRPcaWHQ2pUA3k+4k6euw5I8H0cBm+JApj4K8tw+PdrzBQJLTbc4ci
AmfZHeNyanZKzvB4BrDmRtmtX3MCcLyVnq9XgS/w33cllvbONg/jtt6k62YYy0RI
QfZZo8MdzHfGjrIfBbxRoWSDrYAdWdAWA1ovI1MFLjzB8zFBQsUepkQim1UawWcX
uPTIy4e3zRRfoqnjrRvJdmetF8Lta9i1dFP749I/5AbthW2DVmeWkhI+122bZyf+
YnG0/JgFBTvWo31yjeJstSEMIfyDMTASQRoRG2Q6qTSjtoakndzvAgWJ2MeHYm0K
erx5Y3Ej9B0MnzgCalZWThemq1AQpW69OVLq8S213C4IQFKP6BXb5njxP35vBt00
kdka/V1GAgv+7hVg5sW176i3QcqewyHlvQ4l0ge5yQYvp90DeCG874E5fQxmu7NQ
PTpk+BnhWvzqvakpjhJ2csHrT2m2S5qMk7t1zO345Ac5SOO07TiR01clllWJyom2
3urTywhnK9P7UtFJVwQ4dnNlCAhlqMEPB8AnKkV0PMzldWdSQZ0LjunxD75ZTdL7
xxP3nxC+DAg0o75XjWLbTt/9jm8bAuJTodGDnxKmgAr0d5j7IzAFfjibQmLo3xsB
7F/kX4e6/jhJukPfKwyeWwlLBxULc2FIPsggaPP+yp44PELA+qxioiVhpkFCytsd
ihF+/s8P9kXs+uyc1sXg/W0ykwevfjrDGIbqZ97IT44+JrBjDJImdKppcLWnAiQv
0laXqXL/Jp34IcGD9HGIbAkeXUf3rM6LMXDBSs+PMe/xlc7JAAy7NPexT6UTcW0c
CDP4sFqFckR5+NTS6Ti9halfg3Z+/FLMQjXre6WOH7RpI5PejKh4f3Dh23AGlMbv
XXkuYjLP7c22FfLApV/iv9SaKbXPxPON8jcBS5NtWrInKEcJdPmQ1UXc95mJf1y+
Y/kupo0rMK7RN90/clsw5nSc+szYA2P/EXskF7g+NPhIGAaE6VPT81K/2JjBhSr5
iB2jqzy6x7jAqepEcp7R6QbTl2NiYy189LchZ0pTYJMk13eZBvCSMykJE+xzsDmB
j2otzpVPir2JRuiJf1JCyaBxPzwaKE16B0+m1RlIXipt+NjHIgCiHXwmgGPX6x/O
DTgnr6JW89ICCuynRbeQ2BW48IPWmj3EhkBqWKKU14ufXhTIJ5GfQNPv5dK3jPzs
wcHv2kgXjtxMinrVRr0qvrdz3uEkXTJC5DwhjNbUOfgRakq354jNHR9zaQKUG8mc
+usei4uDPuv80SqybgAPn+I0CvItc1+DPFdXh2vwIsjOQl0zGQ7H8eYQb3rQav6p
+azTlzYMwbf/nZs0vIkcFGAM/9Delt4UOebg5N0o3R6HskLsTdUx6zxjWIU/PA9s
xMjv3ofSjh8+BA5dSo9Y1RHe+iNM6bRo4gpwzCChhNxzsCJE4iTx/GYotpd6fWo3
8WqQyh+Ed+4/jHf4oDlu/VEEkd1IbSSVrkrjxvRRCUwX186EgYAAPFtlHTA7KIDW
uOd6WAiDd5aLWw+SnnS561bPuH1ifry5g1JBPe3qa7bz0MzvWCfohs/YjpesR+MW
9W9yoAbwFb6hLEMCzACLVNPd+nc65Dgk8rgF6gGLT5+M5ogr/oSoktxeU3Q0DosV
gtttUDr4OluvOSdyj0RV4+C6+As+9gsuAPNMvLHTYR49dZLAeXl3J2VO8yXItOJD
p608iV6BUAKW57SRHU3NxM7TAYgHFsb4uZU4A8Edijlb+jfHv/cwY9+OVq6iNTMA
J1RuSGkEY9FcLOhMtOil4QixCcFLOgI4bQ2T6iuLYBlCegFDCiXfn8MtLIBiSHAV
4pEM6yZlkxHee7zcWa2474+hNeYIo78wS1qY3oHkwbMVl9qPcLvpgFNUmtAxWrIt
ZMHld1x8FXUvMruvKjm9IDneHPfoj0kabPfmtUP/q45B6EHFeqCr4MyLOnL+cWxg
Evq+NnuisP2snuB3PuSghBWbV8B4gioktgtr/vKAYdDPzxOvWzaObeKw2BAGxEYE
AcsHAG3P8jW2lRfleFqminz8VBqKkujgS9scHSL6uAjxF2Q1iOsHOgmulAk56cQy
XIB1WQMbPiTMeLR6tdBgFu+u+QWn4ZgwtY6uRAWUcthFu/ihmXMpotcc852xpLTN
dLGWorsOpl1BIV/gIEtu2/+a1oc/yqxFO7PAEDoz91Zbv9DKJJ07TPJ9j3z6QRl/
SZmZQ4u0QC5uvZ7n+itcAv023XzEcNDOkmJs5MeUhBaRsBfnzcpWDVlotxkON41j
anpqB0hMlYNf2nAEes6nCXfaRm19XFyYvFLJSzpTczx1biH/bAZZvHddr2exE/h9
05wIlKIO2bFfnlqO20wdRgwvQ4gN9BrLV7S63z7BqptYXk7snY0YnmKt4zo5do4r
FzbXzmiyco4kRJonmxIsfxqmcB+DkVK7RqwEPR5MGhoJMeajYQuxlNn+bGMd4PXY
KIWOhg7gSakWlzZ0+N51pVyLmya5qtrvQFLi5/7JLh5akPI3zhUBK4qzgMw9T0mK
uu/Cy+oeoW+ywIPttSvIAV+XpmeZT7xyztuZqM/cfSS4cm3keUckn1YNJvkUQFZM
NxUOp0f7zKyCOCKIfqPRiQeZx0/ogXTCegLFM9Jn7Nw7Y0YufOuQgGmLcqJIGRwK
4ssRaA1krodNvrj8jEodKr8fv96IQgxhYvRYobutNcWpDhEZcvSJ+CNkV0RlqEnJ
lEijBtaYtDHLcFYdqTEetd/CF1XuQnPRsSSsM2Wu9yhEK3YR6+B5mcjIY3TXsJ4J
ZJx3N9NxmyHNIfJxt8JqgpobUHjMsVWwVTlnJBBohdBPaHvRlkwSKRN+74o//BCP
x4u7tIIZlN8d1uAcZDfQ0NnNwFfDk/QRIWr2vXd8igrWnJivjonpLLJiS1qWORF5
HyMPJd7gm97+b9hkuoIPCoR8P53sIN5YsAWBdKTrcVV5WClQH1iFtiIOhxh4VwzS
jx25TlxReDpQApavBnoyLLmEDIOdhNm10+eilOavHLZ/6UAvlXK3Mv8invvDXnOe
PnkdTSUTJ2WQbvJ9iOGoxlcQzaaeLfMf/9FSFbQ3IZMWbj3xNjFSsEf7YRmj3Ftv
jcSDAxjTc5is7v83g7C2tKyjhI9+o+zy6ZCm/XZItjeI8j/dz+jcyzCUIT8mvV1y
m8tG9AGC/OaoSBaVo3DnXiyDFYzwd/Lg/W/nxHMHLmmhMq4V6t5C4K4b7XYkl4zq
9a3ljdq/k+/TQlOIDIx3nKKsWRqo6j56KzxN8mOLiYt15fTiQJjViPtJNynGKQG3
Juc0pksJvH+rJktUXtOyJdQ5+tOsSWHinGAiq9iF0ZbV/sNLTO0LgIIuC3NX6cvY
ozdtt/bxjzR6AuKvyItO5PZCeNZCHNOYz6YdgjDqEB7Os+obmUDP6+yTIuOWQqZM
URRr9KzHCRPFtVfooAMcORifZKvDp4Xa1LDnshuzNOido62Hf6dkSYquY1gippko
89mUcYVN6HjlOmka3cM182VrGiEqceWvu/K0ePO7RDwV3nmfbjcK+D3/C9KSbLjx
8UcGfHVvwPWf5okXGK6nxJ6jTZ0aoptXz8MqIM2cOjas4JKnhpd3tJyIjb20EHj+
LLtvBErhTdL4nXTTgf1dGZkO7nisQgoQaPoGx2qiMmg53MbWqL5IcRdXBygQj95E
JAEIggSBpGLxgF7ZU0nRI/pR2Kg/CBWTejscIlYoXUx5i2oWeb0qiLef8zpgotlx
/Q+1DeWvTsXBAC2+B5kgb64y/abYJzGc5zVpIvz2zEWG9otTVOB/lP7OnfxuS7NQ
cj7IRShgLUPd40ZR/UndZ/AEfM/WqvsljkbiUP1234MqgjtrxRQYIFrOdkfCSZBN
3rru7rHTI+ldkJMlLCfhWTLDoKQR8XO2CiGDgXY2SFC5/gKJ9BGYxeoIXa+nHXrH
50K+xI6hIuZwLrYjiTyYy++dA+bxzNULKxFag9CwMWVObEuSMfqO0/eBMvcpVmfM
HSx8jfBNJkNOHxhT2PAwi00JxuVSpsrgpGRko7DHfHATuDksBa/crHx7VxD4GahY
p+9f23IT/RFju8izDOwnkv0EJ6V5p6T8tLpk7oZD0ai7mJhBlHPwUQiAGHAjapW1
UMDx2yFVJebKuuMBcRjvcJUjXcB8htiqNi7TERyziLVM6VqozaPOrHBoVTetWFwo
jXHqhshtUIFD+02hF1fKsuC+7TW5BsEN/D9H5nYUXWY1Dohx9TI+uTr8zFcsUMIP
GgNQqU/qYFZqE9zrYyBh5C4D0qLei6wLjyJ/OecFftXA+JztG31kpWi2oh7x6GPl
VMpZ//DWrv5O8JK1GQvO+gXBt62G5lvNH42IWCJo6TUGcx44NpfbwRRU0ZrO9IeB
1jJa4KB656aJo6nI/dFpUQVCnqHnr8mvPz3bqDs/v+VhAyoTZVjzWse7zlW1akMe
YomCBlAAuYB4PuEytBgLEAtNexK3l2yiF44c5aLmPFT1egXaVfv3CB0iHbAWPElZ
uSHGzLuRcrUOz4cLyg7EC7F5DBRZX5yY0TdL1iCgqGhD+8Ide+WKEPIarljUENrn
Qzk+BCeZauQg9vn/Vj+Zli7nJ/nIabAOHOd7u0aDfjkw95NJznqSo9hno+4S9zGS
7Igakbg3ve9/7LdWtDE4Y52jCXx616QnXgqTpk7jAZfKdqOS3eAmQrm8+OJYzdW+
jbYSDjfVaOU4UiDu51WaKV+6hI+EG5w2Xxd3EVo29wUUgYzHTJy1d+ujEh1HCGRg
e1PjuhyxjdIFAzB4icxESetlWTRg1/S4QLK9pq7hZCVXFi+vlE6lRn8h6qmj5h56
dLt9ibuxK6UeamnchG8/j529MEU7/Y3glXtpReOmbS2XO/IZ8xgnWZ29r//hPe8U
RXwxCllpd2EgTuNy8U8j5Oz1nYHjJf+SXEWqCR9fM0ruLRRjlQl5uNQzlbVVrU7a
e6gfEwQz1iZK9+0GR03Tof0VnP+yTwlz+XeYNJTNP+093N6cxT+HnaRWjD4CbWvE
3cNUkgOujRxjUd4++I7oxyvGXC3F0eEn9kucGEG3h/p+RFb9JIaGM4MqSYhMj1mi
pp7mnIcs9jK9PGXAl5l6uddpMHip1aO6GaFncxoq1iwkLA3RV4dJB4yNKfFR2Ykk
CWGXilKWJXdcWcLUluGbmZwNUcR7qfG7ehigEKra3s7LmILIbP3joy/3OtIBFpIP
JYq04y8/oyHzehNGDjU3aTTGsQ5Bo99FWmPbeFgJn0jrFcTNimP5FiXCbI/my6dD
tjdjgY6S7MkEZCE0zXbireyF0z3htaoDlmwP5C/RM9/FSgLvL5hOIdxeM5mASzCg
EW6G99S/OY1/O3LMH8bMaNpI4N8IHRv3g34qL+1QdSpsB6h8uPHpFX3Ti7qIlWwK
kj2k5/fhXBU4jWnLobAUBRL9v0dwMRhjqvcYiJC9yEvBT62jfCFbdNjoViHwv8Uf
6btseyhXpdCqHJgHKIgSmLVwU/AKbceDlT/EmJHgBh7lDUsQ/ufGjQorIzhS0evj
nPYZWSzYhBTcEnrweAMGVrNagIopG2JawGxwggPN+9YVjSPa6f+EMc4ktkKfWO2W
nW0uIrQAipGuws3hW8Q0Z50OLiUhW8lS9mefkC3ZCxFRepowVTnY1ZpXN+DJRhWB
6BtcgJgxG1wxWzHXsxJJpp2cpKWifiTGO6gvliO1c7b7tGkhKcaSlMA40gVy/6rt
N7gHluQguboHABMGceT6r5eCCSpC3u1ymt9TouvA/ilLw9XZtg53G5aKdWBWDEeW
cc3+vZivtiWhi1ScfiydBc9V59pu0I4hzvnHslqndEH33Df7eMUf6dzWhgZ3nArD
5PGvvEzZ1kA3mxDhFugLFim/yDx+r8u+OFDJkM1+n5Pg07kCy54pPNbmCnJK5uZA
u1gLXxy1Se/hXDbQPGarLv1c15o6xPm2wpIu9F36sWwNRYFfx+0/z81vxuhkzwCC
EtkKxsJ2JV2InhY7f0oSv86Vs3UT+a3lP3BNv1FdcuNqw/rbHIkJLDeV1xoTd9Ca
b5z6r4qckaAfD9qAAMR0A7TW4fuKXi8NKmtxkj4D3xkGO8y6O7nWGNlfX6xBoTK3
SdYF3k8tQS3uTTcCBE8EL5dnEAbxkl5Sc9MoBQ+IdKa6e5zi669//jNpY6y3d5dx
l48ZrfgrO5NKxnM3s7bx9TJkLldyJm26EkUlXIaBLb2POzzbswjmHkWAWJdIKecN
HHMUCZsO8qF9gLc/dgyPQkrRgQfwSRE8N4Xhr2kGCKk6bvTo21fECpb0voH2Mv9f
DynNpSlwy+bVfLs1vmaarl1r8JszT89nqjCmQaRSFboIKAPv8RlS3uzo0YcD4IWS
bSKjzL2IOi16AX1N0S1Z2xOMH82ddBCvQMFTd6JeMgBt92yg3q5QeGwuaJ0QH8uU
QqCiPFCIL/0r8mpctLhlwLH8d6iNKr7ZR917KThqqTAAB4gDwbtObORO5H7AJ8wZ
RJsxkjLda56otMSouycKfXlJ4eKQQuOn3iGguWUrN56Tqz8JdliLKgq8vMp9OPb6
FfhyTp7m8oPohMVbhVNHP00RVXEkRm9NRYyAVoF5XOEZZhO17CWlXi1oPpBegxoW
wB1XhIi+Stwe/UoYX+WEBMC8Amwl25b505R6Rg/Kk8hJ2SEkGvYQ+RFzqdHZTehL
+xZOvoO0xhJHfJF46m/iDosWj/3EHbtN4obDEo0cJCqJky20t1twWtav7yWcG8We
su8Mfdo7MP+S6GdGYkvKdqhET9jVz3TKLd9iCkDR+s+w+JbG/EfnbJF8zkwbClCG
RP6/rJHKLIu4O7lNmFcmz8OqKfjpHT57/Ou0wGlWmarAfe3x3opQwU5NncKffk+L
DtJFRcjLI+uvefNKDSBncxIOTQR2yNgdbG3OFyh9FTdMR/tlgjp35gvvt2TS7KR4
OW4geYhp/SuHF7P+lONgGlUKh7+Q56GejOir/CQljF2JB8PjRXlDD14y+lvWh3dL
5PYcChKYAO6GwJ+srScoILfbM4jkVpqd6hAnKCW8K+55UoZAUwrzv7FHdYhr1NPs
kH07PazebFcFDSNEoUZ8lVStPsAfe6l+6f2JvwpcUY8aDxYwARpRLnO0E0owrhy9
P2pu3Izj3TwUnkNyWGTa1+Y269qZB9BmGm9uVg/UTUPrflUr96FtRYhSmJyroXaO
fEkFz+bxYMB5ArC6dkXBeqaFXlM8/Z1sp/79iQ/WoKm3F1mdd+T68KFlxpXjEcO1
aZ6rcAhhnq441sxMpaLqx/3QIYCet4dzNPuU0gdHUy3MSw33L6cl3bZIJ33+04tq
3BGGt9IkW4Z2FymWDHxQu3is0QlaZnzHPAdVX9xejNdz2KOSX8coIPkV796CkSQq
BVnTMqyTlOc2ZD0lD+7JKF84lq1i+w36aEnpqx2oCSKwb4WBoIY6NV4fbEf1GNmH
6rIn4RigKL21QHN9MKeUXjJh+8Ww7J7/I3zhOcYnAejZRjalY5+ukl1ZNkfGUabi

`pragma protect end_protected
