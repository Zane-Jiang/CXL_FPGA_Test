// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
w16/KtHbvbLjqeF31MY7n3K3dM2Ge8MIbFn4XNcXuO+4OCZ4xuWzJ4YjLRVi
AYkxvk1l5IvwexFpgEEmwjTaE+Cm9eXlU9pZsHFiUrLdEEhEawF1g3LyUfeL
hHlTHaC3HvF6cj+EzWATRb0O7fSOK8PEQUOuQRmfbuc8xekgl52xUY0q4qTX
L13tZVlbSpI6Cq+xzzOPthR3r69F9YAw8WieWJZv54eCUeKpvf6OEWT+JGpx
1edh7MuhLbEz9OqvHmqW1Mld7SPhLtoRuBnSahZ5wJlyoxxf0Whhc8jjZmX7
KoqPM2vudaiiVETrVMV4x2qmMafHdPkpPa1tedFsYw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ErQDQKcX83JSMD3HAObR1tV4En67qCi4Rm5bjJQWBivN4qADSl1EPlYvOT9t
dUW2MfkD4grHlaM7ujrwhwd8Y0SdhR227PhnUu/AfSF12ChY3pWdQeh3cI5E
iUSYCe1AyYvPWnEtIaC4ZTqCrElClDeTIOwct2o4RfUGjjFPIujt+42uxpJk
qIWHxsu7tLacgAEUkPONbSRBcY7vLmdvHe/XbAbiKIeP2PIgS+hnT1IS7SPo
0Nrqcv4hLAGFkNofNs8GywHiJ0MLvEhVD9lM/k5jJfMAZBIB1qashln6hui/
qrO0y+yy7nBteKrLyUlYoZOSOi6TndLC4+1G6UNFmg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b+tgm0qiMdbtbJr27lRmjoX9cincCMclL6zYAkr93d7nz5btcjF7xK/zZJOs
WnZtBN1JzbF90miqMu0If0NHgE1VvUEQLIb5mMZhK3LEsVJdI5rErZJ1xHEd
UxZGR5gkDRtO80p6q+upxZPQs/7n+9OF552lL3vREhpYU4GlnGcaOrtfzoKC
kc3jHI3VpK0mdHLYo7YNwIPLcp81L/jSQ09pt6iYbGDyACPmoZqz06AJOg/H
qtxWRdRieF/mKyDXAmXrRmE7s0GD8sbC46ZwFZS2PXmWLRIaa/FqPdbXTvRu
MjtAVKu5MeajIpZklLZHqYhmSuQwlImc20McbWxABQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ic3CFHT/aWXeCj9ArfaVdThBhp1G2VYp1TTaUk/+8KYYN5Ggpq2qhXSNViHy
ZKdeX9mCN1djWdjco4sObJNwlMcuyvz8Ztte58T5iH6NeyVrRk4Jq76VDVTZ
HO3ljZJQ5WFJFm/nhQPauUrduKmvh2B4PC/Jzo/1vUYUOhCkE2k=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
p8UunnSgl9WUBCqN0HP2fAnjy3XuhoCCgKdoCt/NqEIiRf+YJecrPm9SEc4g
9RkW540E5dcy1bRHeDMF4j2INui+o3ehakzBVvOz+GHkskxeWftLYC6zg0et
EVCUMUZUAQJn4kzMYHE167VvrsckW5GPyeRmOEjrSX9+R2tunTah1M7oHCtB
vQM3/GtHaICWpuKFlMxSm4iPW1RU7cUF2fk9ndMztPY2NE5c1ZZOZCEGFyPy
gvRUOGEcINlBKegUWH4/Y3NziforiSvvQ7HIslx6AxRhDb1njEMyc4Glq+hB
nU7y9LkwprS+N+jvkb+DmWeFPHvQ/+GWjeq6QSZc0JbiiC3mzlM/YVcSxbBN
YznhxLxFLSgGiehAIvP0h0sI2VVQeeEUGTv07ukQjGu3xwHSIBv4kU7G3xjI
DMw31GiBuzJUHP/xTSYOCcW3UrLZQtt/1t9wONR13WChJ2gG4cJTVKRfAF8K
v8wFHKqfDSRheRGNsJiTYZSahzQJzbB2


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TWZO6gZp2AUKD4eNbKpNyo62WzVC5+1vcVwh69EzsfXvh0sHoj2YzZVmYS3x
hiJVndOi+u4OBplSiFHbKIU0Zebn0Ppbw0abHjnE8FgwlyE8nVLtA6YqRl0T
Mz/jbEO+6kPjNYXi/fJ1xF1HmtWBUGnRDKDcWBsl20n8jKMa1yk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p1fGaWE4QaPfjhQm9b2mkBSX7v2pffxkL1vSWt9svS+eI1kKGmdfmkGME5ed
kIISdIcLSUXmrNDMEJpj1y/LdpCAjuouwIBC9T1oyI15p6025SfpxPMYsg22
Nc6XU7gw4DzjKsJSXvMD7aHBs6qDhyUATs2VbxEcEFtz/7zpZoU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2464)
`pragma protect data_block
CcJlb0NjOGTb2B+Flea/up8+WkLoLq3pyO2jN28uniySV9AwRwkqnrbrDbpF
LXaYGLP52/sJUDdAOTNCqQqM8Upiu7NZQzHSehvs12vvyFgb7uNW8z6KA4jV
1Jx+CkFq+1NhtjuuxfOJli/iQZWT+PAPt8UtEvx+aYLqzoKEcFneF9eTn1CM
ar1s5uIdTGfMe0+WgemtAyh9RUYiIfbrJ7VI+SRycebk6iY7LtBuuqZ6lXKQ
NWswIcPH2XKoOZ4kjWCJeL/4+XgYMKuJFuK1lhOtidtD8MgDOnSd68cYgtaN
rbpHd+MtkGh/bITUxobPdXtgYJ76hz07tPd0NXfssxGYhacw7fe3wQ1jr1SC
1ys/rG9JK5a+u8HNHIs+9wweyl/ytho8ORIsc9Imbl0f5vA7QXNLrrKRCAjb
oUugQShAFxLxVMoKsEHs6JxSylT7pUobJcp2Cn8annOkAoZrLpFmR9SAzTEX
JfpA7pjfsTo3etL3BJN+PhnawLwB3Qg0cbNmRiH1BgieoT6vDRjSF003Svt4
JV54jY3UhzjrDEgYVFz6AO8LnVtpbdCvxlmh7xejTdp0YOJSq5YLh3H/H8oS
geo4oUaOFxhTakai0a/N86zjAuFj1G2VSQXsu4CsVmPrJ9NS7D3NlX99eYzn
1UQkDlqJ5xlU8xpta4W/ha9vtDJVKSaSg1im7sAuk1rbXcIWZhz8e9fUMFeO
FDZUsVcRaOMm0ZKKsRl0itqr37Lr4sVAvqpWBkik2TJbIMv/wIsMaGZQfJSF
ABD47tObFab3M54+0YMnis6/E6aX6j2PoZ/0ofF0gunF8epJVyA8nIs8FS+V
gP7cHcZpDNIfAABfvNclOgDmfMm34ZrRST4oxgONYG4mrn8KY1nwt5do5Mlw
vG5yQolDTSSSdzWJBwcPpaFNkU1pHLuvdBj/pINrIWL5mM0FvOBYm/biPY+C
g7YtAvyIaEhTP+c62P+CnSZwdC/BkA8/szvxy7yA9KJE+2Yjz3cGXZOstOFO
/iUStn/aTz9fexbWwTBAzodHJe6f+wNFscjMdJbizcYstzgVcwdTGeJ+xeb6
LC2SLvyR7FS5pcnz58MFAORyUsUB4oAeR8Umz6vOJVLDxRzF+Y1eNjaDCYF+
jLwauGw/XB0Q7JUaUwfHBghWn6+kZX5/3MuLnVodGib7U3eMPVU3NQvCottQ
SgbgZk/DhmGpd3MpKUpSzeUti6HPtf+2UUgytUpAbJhwpnX2vGyvq5/spnko
xK+tog8oWf3Vp+9z4r+icbxOvn3GqEIsvLvQjzZvNfc5IgwILjhnJqRnaYn6
WpG5/buoQg2DIwVQiyiKgv3zGyqXoyBzAPZqzcZw3Om1i7JUoc7/zef4QsO0
sjYUhk3T/q+1X4cGEut2cZ74R2aSb+Dyz2zqcH0STMapwVPhaWW71rVgB/aG
RhltiCe4+wAO4TzJdr9Hj43vkrqxhMVp0ibg1V0+h8vBlr39i02g5biXjNZ9
BzA6e7Li6igdfMvroBdca1YmgwhhfcocIIv320YjuCntzzrouT6pUZBr3H7C
JtIdzCZo26yAKFrmuaTC6IEoGOX2ej+syL/sfV9tAnxKUPME/njDUbxW5u3S
31eGSvyksILBj+oTuiLxe65I7l49wNilsUTTIo3h9uTx2sZp6o3ptlKmoBrw
yB4ECmIZ0m+F8J6WDv67/0JDp5lnk5RX8Q30XaNychJQ/eASbWhastsdtI8j
e3z+k7crl/uxG4u4kOm72r5Jk36bdMJ4zkqtAKISam9vnZO/kYZF+ynzm3bk
ngV/DMlubyOShPcE1JJtBFq9UqkcuuUpWYQu1xEw2b4N7C1T5/rOs56U0l97
wPcRyKD3muvQFH1k0s5oM32T1g9JXLbxMs7DOCbfohn0KqdndNOYaj3iwTUx
vcJyIxGuGB6+LG+pYnWfrt3T9SSOzGzSVeNZiN1LApHTdxzMGEnR6fwAL8EL
/JZRPkyjeYLfWU8JEaKnI+HpJAY2M9A1x5KVFDcRTwQB30CXqlg7ST6uNU7p
y5eedZLISkgQ3vBNVcOZerhV7pq7tOewITGjBtH6s7Kl5159Z2F3hgAncZgo
Kz1q6zmDiK3WkrWTXHuP+G0U3mENbhZZB8PEhiUpLyJ+ciMMvymjjHuiCc0X
GioEqLGRZTwfb4GO3TiKPwo4W64Cw8pGopp/xaThQVvacYh0QG7fHOLn/HDX
5Ph9AfrqKRejArf5JmpNQK1k5j8qxgE2q06imXPBlvnWI8gyvupH7CZsgTwA
7kOH1IdeHCPfqVk2UGR1AytoFGsa9WCYuUdK7RXBISr71CkrLhZQFNVLTBJO
FWyS4Cl+7Uvbno0dm9XMyVcCK7gF7OVjQe08E1PWaQy/zXIijm8U9IeIuDO7
hLrWeeGdDbj8gw0Ixc6sZ8CAeY9V0BwU6O5lmdMRK3tGgMkms+qS1GGyB3rk
0j3Bqa3b8AKIT/YCwN3dtYx29YUOGRxia29HIz91deNPJgQiZp1KnwcZGwKs
65tOjos2rk7yLXVkrQVVjHPgUMYB+XPHepeGO5pcQem7r5aSBi2bb+GcBpgN
iwUlASVKMBJcC4P7gnHH7fihK9TKF8WbsFMX1a4vW6ioLuGAJLwJtZBJ2enh
cFoVXen4U6D1ZtdxZrkvs/fnd2nF7g1tsNmaeLH+52SNGeQpEC5wx/E1Huyz
fptBFO9O/N+lJGakBdyU3KEgnAIxo1MR7BxWgJe8ZbhicvSb3LacJyA4sBJ8
6nQqQv9UqCXTMo2+kB1d8RanvSfcl1j3z5N51/COHwNrbi7ovt0aEPFua7Y2
94rneNglpKf5pNBPZ/4fDDA5L190wq47gfXBXwyvU7vavL0uxWxV+9GSTtwl
DYa19I/M1tZbgbVbz7EQICkyaLLKuk4O3qQi0W3T6PvJuSYA8WK12Kji1Oxs
kcujGx5Sne00fsl85O7ygX14DllznLd8V1ObnSaD9h4OvAbgZv1XpW9+Wuvc
DqzMsmfKJr+6sGMrBCDuKmHEdJK1HEH2qL1xWUn/81Wv7xdtVjBDaG82RiNM
ldvv3n/LTmB/ML7c4Ct4i6GIa3QkcuEPoSpUSuXRUmvOwFgL9Uw6JgaPrM7R
3t/IwmfNGAgT4btHGO9URp0CXJDggZX9PmVhzSXDW0hY1ueA2vIep3WQlABj
Nh3spjeSWPagk62WyLBInkGZJ/qStBjWkT7zNzHA6f/V540fdACaPCvBHLAT
5IYlCRW7jQ4Ir/Qj/M3iyoqNmbPTuq6IfSo6RVXgRwofrw==

`pragma protect end_protected
