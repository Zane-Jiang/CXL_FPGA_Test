// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
jDuhdtSZuurLJl3Mz7Xi4xCxE1BZaHv3BiAtgH1GvmosRGN1ihlvbT7TyRDjLjw0
dlb5U/Bi32CKaPhmd0MCiYcaBHwyAw8OYdRnBy2eNoGe0711qNk/0JAST6HCtbO2
HUy/pcKN6vpaGdTarmxUl4Thm4/gLSxdixICcdOtTkM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 91088 )
`pragma protect data_block
5Wv3x7M0mYq9nKEUkGkqnJnoTRPCbVMWz/dRsj0ra17TNG5x9hqr5ulKDBll5m+r
Jmtrmu4OU+MGgsKvdfhumIxBMT+Vf2saCiO1+5DxM0eMPG+63BQ/aSDSpStoCyd7
aHmlAXGxC+AYmYjvmsAKke36QphxCoIOtF2b+i2/pAFYBxrCFOMoqjP59Kh2OIN+
KAWPyapZh01izjaUf0DKJ5DYDzVgdOTIPlJnn0BW5gMS1aQck44PRER2/S/+3MYO
bWL8HpymwPZ1Q6c0VVp6cUweBSp17pCntCAtj0si4BijSdUvlmGNXPTd20mmp++h
XIwxA3+QLewmyQkpV0vFvDOcAAEoF2M6k/9Rw6YwUPwEwgrDs/i3Y5rXl4YDqImA
GIQxJ6tsrKPWUnoT6bFJKwd0cK+4q+C3GBvTTJtBdAisAvrhWzLNukNIaf1GBiB9
R6vioeusbDhmA+oSSFXWrdMrLmlMl6uGnrKrb5LE2Ty1mLX8qdLZCAeXn+nIce7e
nXvKlN1k0j5cfRab6Hm0j40doRqnGr/m4fIPB3kpxlLMj7VmkO/3doSeEF6VlQS9
ZXZVUgIaif9bnNOWM/1XWreYTBLDBCP56kTjfuVSXx5Uj0YbrfK6c9ka8O70xjL3
j2V0G49UpyrxIgHLglv1j5gTFp21o/CGmgGhMgA6V4K7yIDCtmUh9wTs2gYqCV4t
IagQboYICmmhD7k5zSSSExsu+Llmpq1a+MwsbSTcwYzxXjAafaehPvP+9WZRdtSz
rRe3MN2M9PYEP1GuM19BUSOOg6FSUc8cp1QH4hq7z1jNr4D2IG1LOTUh16ClK3kP
QZqIbAc8uznptXofCCWiSderY/56o9p24fKslNzKoWkGEg6cCw49aVYAdVdtL5Gj
mddWWGrExoFKl4cJBm2nGBDnrij9lwPHBzItdQDKN7nvtGsl5nJP5qjnttzS8gns
vP+voSc4H+LWcX0Ip9zYVIc1UEtfEBZebL/YlIHiAu32hE1RVw1k/tipi6k6kCId
uKmf48hsCHpdaDYAkScGV3yxzM6caeM6h8XLti0jer22GD5MeGQ3/SOIu/Ju5s3K
TdX09/0YEFJalAYh4rBLJA4g83TFa8y5+bF+hb32SPVsg6wS++XmQwpJof/UNEsV
2x5/LZnL6L0Sh85ogE9PtiaUzgU5R5rDFpGp1qIBhnCuOZYEvMHXHgu6CtmCPxJE
Yo52QFLynFFuY6FgoHg+JFptzXze1DC45Qni1Q2DSKYOroMlk3w77ElwdTVv1peq
VDZaP++8+m5vi2uAcyM064J0F5Ga8sO0L9BjALmwUkbA15IE5y92QdqXPDinQGNZ
lNQYI4FU7fFJwmXZI0MjQx4v3twjluZAFVlqMeWt0xmgZdbEqgQLbDRT1VY8rOAe
JLCnaqTdeOSQWahEd5Ranu69xY+pXWjVLBGGAeJffg03T5lcmsbX59fZ707lrGNs
oZvEIEqNVxpt5rsDzzg5VU7jNnkmF+/Z3M7+BE/BjsptfF3iMp+CAi2ZweBmdPX6
SeSe+gaYOGaZjjGnZsB+yo4Pb1tXWvjzILXB2RBFukUmgknwAgMoYghID41iwHYn
15iNYulPOLGI/+hknNVScMwIjDRNFq97/oTueQPIIXWWhhMc4qp4Qr5auywgWyGX
a+iWCJecFEcXVxm+khd8xi0F/z/3kjsFB5+Lp8h3awUXjblJ9p+4ctmdAKHzHDz3
6uVORjR1FJ7J8uUbXA2a5etalDJ7y2thaOM9xHM7ylt2h4UyPOpodLJxK8QJi2qD
tGoVA42LONPjOuGK94OZFvlGovjKEFdFEH5ElORWVpg4V/EkXUlsAIe8tUMG5Vp0
BEAam8ZUZsNOzdm8tMtMwLYIENmCuZGgy/6I9V09YDxEBU1PZDH8e+5iwRsfn9hr
49vtCbC0M1bZe9naJOoKGRVG+NOXbBp01sV4p3FKIqqVUCPDd1DXFkcAftsuDer+
3OlBArUXis8Ib6X3YlR3HAukLThE5nJWICjPAPhMXjhTxY2ExdkiXnsGgFuwC9He
5x7lN7/siO0NRjCxNE2la5y83uJrRGt4WN97iaDiWBt4nFMglQkgzw6ZwsNEhdaw
ou2VqQk2+mPBZ5cCCQfh5iwnaVy0SaL/6tOBN6G9EhMY5/UZyo6zY11dbprnSf7P
m2gkQyfRTPRWljO0EQ9ndxtOpva5DDBcj8GwoorTOeq5twJJgGCBVcoSHMZ6DlZy
e6+/OdSg3xtJOwF95H+wVhP003yaV4zOxJAStI86hSZAbRRKfO/7DXrMnmB+JRik
dWcB89ABVHpd+j2QFuCD4Ap7PBmK1WeP5K8GDtj2gploRZJOIetMLzH1raVTnawN
w45vBmyMWM3XLs/tpe7qdmzRir5gqi8GOCeV6rialpcQJuZj3O2PMTJzFtI9IaLC
GJucNxlgeyBqg5QimSdyQFZjDUTdbV4UpDNS7pojL5D09W6P/jNkIQTgtSMLsMj+
FvsCBRCr9QHW/ZXN9shnZ/WRzC4MWjTCH6ovNvACV7quwcnAm582TXeEYLUCvu7O
vrsdZEhSgS7g4UZr2r5HV8Obf5aY2JK9O9NSJT+D0UWkX0g6zjWaH1CP/s82vqxa
5NWOu+zduzMkyA3kGQoym7JCWTjtYtUEWMbosA6HrJIfdjDAX/Vg+lV3++0VtEvS
14tm5tNNCHnQZot9bqPy3L2NzNOePEj3QJJcuIaQCM1kZ/VwOfmmf/BUW3360Bsw
UL4Pw3xtg/dAtX4zq+aVxlX8pT9Xyfu5gLkQNSTD37tZWvX/5qRSLrkccCH1gHlk
7fevm/a0qEfUni8asdGFFarXjpN9LK8LPX6IB3F7PB3TEgH7NQDM+KSZD9TSsCHy
iyKhgqZNEa8oa+hp7HdUkt4Gj7/RtcOLBHKUq7gyOy1rQE+0hhNnlT5Mb1QyStn7
/33s/ym74TANwyl5tLXD+GcdHXuTWi2Loung8XGDTdP7EHVncoN15Fie5Qsz5e4E
aPlOKeX2Po/dq9GpLCtVygsfrA56QWOl+tdV7yheJrRRoXjxzPKisDonL4BaeF/E
t22CV+YJ+RxlJCKU1WjD6n/Zbbi1VgP4hYECDpvSf4YBNlbDHZwwan3qnCnC0PEo
uP2x7srO9DfBX2OWBNPyfjuPu8KEj9PtdTS7nLAIfvH172p3ot5Lp4mEN8y7mRW0
W1B1Dz39kxl9n4P2v9fm6d9B0eS0mA4kugwcXwcfrDONsJopcGOHDHS5j9fZrV+K
vVWFjy9xJlMsk09pz6rXkPd3irx83KMRgXQUYnBm/fWwax9QyHgzY+B7rcfGMlyo
F47soS/Bs0llSqvI5I9nkujG4QUj9Llrb/CJUwg93d/zM12oFi3WoyqzHxtusUJD
l3wwmNLrMCtvlPk7JzvHahBGV8qJ5j+XVJQtkzKB9TMRXWEBPj/wljWf2+gEuYjC
CBx6DHfaJCU8CGU9lBSYw3H///4W6xExGTCTEkX9C5EIvDvgfAHhAueBhh7YzxNY
rwtpQtB0X3Uc/uGHktJh3iGgSlOtiZ5vnzTV9XqnphwyG61rQsspEMegA4YiFiMr
3alnIz/eUYSStTEedp2AR9Bxx7gh+6FtJM+y+UDOZuoiRClKajND0q9rxhBrQpmQ
yI2UvTr0ZVyOmuyy6x1PTsNSoey+P2zPoykf2fOcrK9yYAaMOi51+96RmqJAcJKO
F7TrgzYzwrV14GRkxynk6ZYjiBTtVZAxvdhh8A7Y6GNMMqS4/BUJVZCilnLj7W4Y
lEzHFV1uSg9ZtrZ/9mk5QadF6ghsvnqCW62fXX/CaT5bo+FFsU2Ui3bkt0hXopou
vkxKucfZ2Ze9Lc3vqwCKyF3GE8noXKEIbNsVw6DJEO8Cte5SiwTwNwtx2BC6KjF4
H9FYZMA7DrBgWamvgPGF/00BkEJg6ytgvs18xXk+abZDJD6BMRvWEgdyvIZ6UdaV
5X6x3rh1exnhIEa4KGjkKDgujp1N69F0IwmcmaL+CRjhKqUMReVes+Xhn9tF5bYU
PCccsftSUFYvxVswmLhKyWXxxx/THgwoG/cTqsTan9zUhKeDAgufgXCnSFfM0G+P
OQwajoU4s/sVhPkjDoStvIBzVocC+uflADZlUi7IZEGFAmz8MB9tDV6QFwqZnDdY
N5Hsacwxleavh4yl6JisHStF9E4qSz1SCb09NoFslqIEpVRdTsXAJ5GTdHwbIkff
yp+L8bRbcWD4SY/f1jUHo9Z0p2Xk6q/BpniC7jZVQJvi/XDR6Jv+VBvYqxFRtKD/
nI9AhZ/Wn71rQ8rpX7uWJ1w/9DzYtfEHfGWr/9uJBOi+sjAQz8GGWk4suC+qDHKB
2aX0nGLrcf2ajHIGmd+PmcwgXABH7nsMQkHD+gcoLLDZrYPH22DZjXzEHLR+2iLd
BDqDGbnFxa8lkVdsaoWD9+pNBg1ltpQJ6z6NtMqeqxLs9mwwFaJ5GWfqkkeRWE0S
F5DvsZ+Qer196qQiE3PxNlMlNWqhd2mljq4VePEFJnuioap5K5efWUy/vYIuePfm
5CK41in9JtsF4C6fe100tNlwK53Zmou6mLEe2d9AuQ6h7SSz0+hKv6LCWbH29aWW
O++eek9SjDbz4ZhmeNvV8DIROPgyyX2u6B2F7FvS1pnuhzPXebPxTT6SeRHodbBv
MdpUQxsIwe8+9v+R0UrEkG+jIx/eiNjOtfN65qf2xSNLESR86wxfk1EOxHRCG0S6
4Y5oohowOqdemsTUSCZiAn3Gmqig2L0Ab+/GiQFnZTfgLJeUwT/h06Q8aJ5F0Icx
3iY8vFnJ1TbuaM46VHvC5anxIeesrM/K6H2NcT3lj1pNIndOuptOiBKFlwjBUIyQ
lucCyJuAa0khV+MHLpdNbPENmeaDCNo8Xc/OjKHT6ZBKAuiQGAZhHxMLXSSkhA+r
CiXw25n/3tfOY4NT6kr4UcGsQdRk/s0/eDXMUJc6Wj637PnAC/Fe7dtdXQvP5KuW
7bWhoKkHReq8JZHbH1pG8iS2xra7lgW3SveCHLRe3QkIK9iDLXNdw8PqRWBZHnXu
VmBLRJPHAHmP/8ADxK1FEpkCK6FPY53fTA4yaGkWVJPVpF9Eg7a2NIzu5OtVIM26
ISgXuNPUOHrS9UvrZsqzLJY46AIA8Ph86o0CUL3p1Mvg83Ec1nZtIxqtiTceIkPs
JspOawwICk1FTSmCtkEm4Icrf7cqzQcKC1WpVOZxdlT1v9fuWRfLi64Cs0n1Rpi7
waejkfR6rHWPPGlaqNs5/XaLz516nTsPMbQNmsx2GY/RuHdFjYI4DdEymIk/ThUT
cwhVnud4+ysBaRmG0nXkajtooDYHdY12sdm+yjLPWiycnSdxFZtGMyC48njVFG9t
NTSGE2nIYdMliGneJIJ2fS6G5ZpCuNlonzCGxJpO9MPx7PdVQIY6xBjNtg/yvztd
l0xcNSdckqRh/5Nur+Ow5dOL2+djEksHZzBCUD2b4wsySqqJmm1u2mEfnJSgMk/X
USfIsJd9QVdQRDsVqgu4P3rE9iIu4kGoXz9fDebxhPgOQ4s1ErAD6UX9m+SPNwer
yy5joJwwkBJhz4v5B7TfCUGiMjoraIBg3tutvw7bl5wfGmmWcprHr7S2Z4oNYVMC
QUAjgBe9wdSWtziy3Sct3A1W5idN19UJTjBmRo/AZ2d2C6u9v3Wdz34EJVETV2cl
Sgh+7H42j8N9PnbS6RSyBBNLOFHE0kV7BM3Grhnn4P1YMWhiPE8zsytuePSGeMqQ
IT18gB9zDu5wylAYfD1/ZLXp4DelQ5XjRzdxcRse9K5J+4cUPgUgsaOkONzEGtAS
PUPCF3Nu3eTCl9A1NJoaAz3Zn2GSCnnsaCb53274g8MI2fh/uDJrjIxet+Nhe4fp
z3qegm+B7E6ieley3gF9cQG2o8fEe0zKz5jR+syTfK7CpaBN/BouaxE7JbwIKK4r
INFnFg7XfqNA24dnfGebo1Fe8Y/dPTGtXo3KPi4STq+B9am4U0i23iMldXPtJDBy
x/LpIiOj+JOXFsE0vF6J3F8tmPUCvGxrU2s4ZEyg+Djz0F43+Q+aKFXqq88MfK0k
J9ltqFGHubx9aRcA54EGfujclRNXvaraQ2dW/heQ2C+GS4ayIWjNi9vwHSAe6peb
70HTLk4tXHGTJiMVAOfEdDoOV/vFoQBm+cBZyjiaVqs4mD7cljj4xsF72LtgHLRb
8FUO2bxw3hwAymWc1jtc4YleFKm/q6kwhI1jvIoVl1VUxgtbR1Lrq81ripsMARzY
UaecwVcdBY0Sf7Lmshx0sl1jwvGjU4Fp6YoSemI0hbat9iqSi+DFuyd6WXigLvAL
mPZAMBHjZZKSfnuB060p6XPBPZod1+A1KnLMxkELbyAu8pvcx6CSsvbuvABo4s7R
zRhNsaACCwL3G0cAqvIEg8Apd8QD1NToy7qEAHxi5nkhT4lKCPybVTEeysU33mU8
rkNUOdNAMKYbURbFskWaG+rIFfaNUyqExW42sujS7DJIa2ocjmK9pJRxuX8rDV87
fcqBFOsF33paHgo3Y2qSHjJGtMC49niZcJq6r9UAFmnWFh9ADX6XVuajARw9K+Jc
1kvQ+uQOSV+oNWz9ZiX6gPu+p6oSH/cUTF0N2VdFEw0a9TmMDca73fecNsI3V+z+
GFN70Wbs1bFXQG+t5YdpVhKlXsEujeTuAYpwt6SqC0iyF5XrN2bGuXCZJKf3iV36
+cS7GqPFALx+8z4oRov/wvWrljS08eeoum/OLBgpQTsgj6U9w6Qo/f2l8OSjBSH/
HvNRZcuZb1YK8qlHuprwbxtTZNodBIdel5cHxA0g4A0v+tb32GlUIb4PEdz1otU7
l5F0+b6CfkBXpmYQ9ikgmMsb8HC0fNIlZ34R8CIiK9XUMREzi1y0C+30+MAlnnvG
zhiIRck+AG8zPLLQtoUFYn1phcvfmMXzPrucnrC6At5c2Ekh+h8I88X8kuuvV874
w8Tl41/w+tHrRWX+DU2jDNOXBRtXr8NOd7YDAxjOExhiKCGjs1BSskg0yj+KGdLt
JEbxzv5tc0UQGhDFqPIJllGqFkOr6KGu5FycrrxfcjqFStVERtvH8ZBoG11kKidv
MvAqs5ZwqHXTx39nerU/tvyzdCyWleFw/VfFGaBLVdALWZgJE4w0rcFigs6ixvaa
K3Ff1K84nBeklqkBod36T2yoO+KBq2S7jCPtDC2Wx1OfBI45Ro66yI0LtPU5fPIb
lhNBEVdMlhKYFEaWYMt7/oAdRF/ipcj/KvGoui2lYabLDSkoULvdQbsSdGOn8ZYx
yozyO9pKOtirRi53jARNNQL4djHFMRzhoeTX01Xr+u/NoVSW/yJFfnG3VoBYUsfq
cwJhBH8RE5qdO0s41W8lB921ShrY7cmDgn/q3w+hL4s5CkUL7Gyt+LdbA3iQiTLr
F+yUG8Vh/Gk+7NfrGjEmSmX0IKBuROCwZYAZahZNYoDGtClYaig7pYtYzqiLbwR6
b0IwhQpV1NAEZVV2Dw9C5HaW94p8SQtcGkW+TtqJrbIJLNWk5QI4LRvlgad6yc3+
5R5LYkmmeDL9Vu4xqc7F/l3TCgF2UguX8CJVyEKBPdPIDppLukXHoo+4U/lQXMKO
TjGXlBvvO/rcs+33oMTV9zT1cbY/1BbUUXVlhQ4Xi7TUFKDdj6fuCrd0b70gmlbL
V8Lx0zwXOGvpZzOtgbKDYJho2EJv7RRF4BMQDM6hBi8Kleb8TSxbRctpRGqh+yJr
EkhpcW51gRLpsq8LPvV9UuatU5UhK7L2PwFvxqmW6VuYW5rpfVKyCrowuYflm6rW
mBQBl5PUcwWAK1KGO+kworfTvW4cLqJtDBaJzl/Cee2dxl4sUJtq/1g74VlxOYqb
6hb9LGkXUFnpGeIVf8fixDAqYGNUyub5LgUU8630ei0Jfl48WhqTQKdBA+zY+ELp
5QG7Csto2yfNS5NmtUmFGbt7atPfjI3RKk9vd3OGxDTsmGoF5Q4v6+5uUTSHcKc5
QJOI8NRyQQUAB6RCo4whdsHrfF5QsKld7j38st8CjULWhrDBxiDTxz08mOaVcv7e
UVuYfbChvpD5aNGNBmIBGuHyh143rQd+kx0V9QS5SSJOiJaTRbDdgAHCejTp/Kqp
8UwEcJqcfoCUVkumRCxcVGuojVVAnmp9+2aT03KGIX6hhmI6rjux+rN+W83+3o8A
F3sX1t5DLkFZTevqjSg8iFAhueQW2XMbThzDRSZnbziq/FV62UCs8oKKnlMfmg9T
ywxheto+uPgq/exxXg4PBDZu2yykF1ug2P6Fk/quEc/L4b1BZvJcU5dI8OiiKyw9
mO3xFG93amqWh4Kkd4m/NRHcuM4e857d90jGoU9YnkdJOnrPSkMNx83+SrSCR4Ml
QtN4cixMI+aW1T2CshBsYYy4Fox+kjCifoyj6jbqiZv6DWSc2fUIfxbHvyKmJF1k
W7I18HtyVD170iUqFAfm4HD+fC6Wk1FzKwji7/0NOpC84iAod9eg1zl2Qmccoqdt
wRFCQtY19Jxn0dxr7QrE97oiVk6ZG0E4oM/jyqaOEyQSTJp2kD7dr1If5z8xgmaM
uzM1SWl7ncH6nu1XAenTq5GGocB3xPnab2mdCz6O97WPTcpFeU7lxvKOgz4Vo6fs
o2PakZiLF24UgPJBbyNAecSodMJrB/nqzek20LKnbA01c8Jl3ergu4hopm7TP4HE
dLTDITXnPVhX2BOeJud4VCgL+pu/6Jt950LHPZk+kUekG4SSglyGBYKfs3eQrnjq
niWYoBjy6vclFReXc0oyq8rngKaYkVmc43HaTjEwZ0Dqck89ZrJRZe5RtKO7X+tF
JXGx5b+bWRwZzrE6XPxG/rq2l5G6OsofrWtBWE4a18vXJWBX+DT9Wu7q+/guzXpU
wPvu+pcNMYry7pFoFEG4rrctxUfd4qQ2gic4zXrjQBKjHVOgoIAf4Zhd+zu3lMco
tR+PFg1hs9sgOzUVkQ6qrrJRfqnQzh9EpDh65OOgjMdbWdB8aqNMEmxfwUIfZPFh
UswE4ZoaW+PXscCsY5nblO+LPPnEfPhbMWXtFl4eHvt6cqVbDKDKPwbajj0hca0r
aUcdygRV/p3cnpqzWYPaROTHnhEtrEzRQcqLz8kdZ9pK5afMJA4aCKl5QdkfNGhk
GzlAC8bv7X8Ww1LQDZ/5EgUAAPc4Fc+l0IJzWNEwX+IUeUGXkxVJ5wybv0aofcet
6yb/irArh6CsP1EXemfWXiC4ODDHQ0qeSJDapW7o/Tr4iOq6tyJhKoFFjLTcX1cd
T82G3SyrFwnyGFkuxE91U2Cu8IObFfar4XNp2QtY0LBvcOw7B0vdqfC+qVPfKWUw
leNNpVtLzm+e9MPQqcj0ei1rpVjCpLJwTG6wdsb4q1VcYJwSzRuiVZop238Gki1X
kwkwMaA7Kl6guMmyGrxa98qfmVjkwPXzDp5lICnedoebq55jCe+fdkC1hOqlX4OW
iiJQYYMfwtmtysk2VH3P1ZOEsVyS09EUEDHD4hkwqKUVesX1C8UW/v2nkJ3TrBvb
BtY09z/c5qDzNby4h1UkzRgMiXrJSD3woHb7xPRESbKRUmHEhEVq8SdBXPA6RyYO
l50tgTkeH8FVY3Nd5/rkcDxqGWKB62h8Wr53ZbutQrwULIrQl1aG2YPOr3mtxzCN
QNHWhpQXcGx1/jxA+K/ampuW9ld9tnd7cU4Xqz5HO8jh3ZXQmBOv20mDNPZdcd8x
pgTzopufmdKTo7B9NDO3E2PvB/FZiZ74DOXX/ChVjD/y62bZVbq/AaEFfOdGwKEE
4251XwCYTvh5lZDUzLHHb4yQjgET8/w8uMLeHbzImKZ6Whdm4AtPeJWbj2Oz5kLL
W5vYqIgtpb9aPEzd3qs/wvjTc2SRtenXEDbCzoaW2HpBDZG9SS9kvM1OKNp10jHO
e8uygTQJUBD6xYKFUFnDkZUIwxMHiBHO9TFoWzYcKPZMgmbv1AImOTAZHGUibtIw
ojPiKqz2ligzXnA0LgcinyZls4TwDrxu0hlvzqmeGLv9+zV8d+4de8xjrBXe1tfZ
8ZlvRKjmo46Cls680emaxueK78/hxijBPFY5e89gYodAyRrbK8kSGfIEyFPP5bZJ
YnxgE2fWRUqoXr+ASTgYqPgNS0UdQB8RMMdNOrtsfOWsa0fwRo8wkFFOaYkWPrBd
tCOBhWEwvG798dML6ZHdZhCf8A6EqWmjaAUYPrrrwgb6r7ceF10Bcz/ls8WLtqqI
db7rnAhZDoUKKN/SQVxwDGHUzR8XkNrQq8sKAdOSnF7xFzVfN9p3OwPPM/r4lJjo
OjfKoPsDHoK6I+IB5gyH58FL2wgz8Apapy1Ggf3S64rvOHZSZy1LfLmCGcKgqIiy
fGlUgryZ6Xho2hMqnCLA/4aRpbni0ZkKT2Ke749FfowwgQ04w7F2+0mndDztLAcA
EEZLadRa0H66YH0DLWS0lPaF/X5GLHWzlt8tcFr6DL8bChbMV3NTPi/LPUqkDuHe
71ZzD4FYFf5eTg+BrQA49PTcDsF2wDJ5wB1iK6xJP0C5nRLS6Ja3636Fu9TKjPFL
1SHb87UOsMqpdasY7c3/vHDiMJlNDDe9ottCq7coZD1pBIEz9knsSGxes4LHIqs8
TdAAzvt46x9+bP3Ba3nLqLh+5j0jiJibovh0e6+mYaCP1twosdTzhjl2rHyB/3ka
aPh8deXeOeqzsafjJ2EUuHrEtvxKGFuS7HHCTeFndIJuX3773zy+Lnu8L/Baeu8C
rDevjoEnZCCZMfgcNtDFxyOWVVU2FzbjJWwXeHbMM617uLugK4YsJRiRoxuJyqSE
R7nWY+97jPTA/QaV1VSQnyLZyfrLEQoT8QBXVJMcagt35v9AeMavjZY/fFdwgGZO
U6JmQQLURvWVcgVAYolbJ6Pw7iIOjoqgneVPX8AlP9JicOgB++1qCBw5vz5J/rKV
mfEMjEp/xNrZ0phvA171LzJjOPUg//S86Ui4zvQFlBnW55gjoAREF/8PLSZttiD4
FisrzvOPShcFY8Skg7Xp134Tai87DMGjq75DO17I8lt2+zSAd8mY9zkgQxbr+G98
DYVfBGtuySIdO5DrQIk6/p1VNfucsQxXsjlgJ7wNB02uAsKQjlqxNzzCOU7sb1YC
YYMJJFzDORo4DKJJhuXYTg7yMn000bOF7N4pjZsA/it+yFHLO3irVCQhhnJOh1nc
974FYNRSVOYKf0gKI6m/XjcBpJxzodijy22GuMd82kFEFFhu11FQaL+eNaVHxbyi
3VqYw4nS7Z6d+fSSigsXn/j5gKLcMahQJt078ooEAGlSG4nbVXvdNJzpCXT43aan
cFPZMgD3ICaI1H6ubRExs9RQ6uEOHengdk295A0A2Zh1uX3OmU0luNSZ/e/3/eKZ
UN8PpcUTa3yaRSO9/aZv9yoWG2NZSmu7hphwWsynDoQg96UTaWrSZwxrrvP+i9rC
CzkxNOSvCHWpKBLFzJemD+QRkRquKZxl68hqHpNplcB8j135M6sgzbY+slEqOWJl
Mb/bZWjpF1A3ptxVTLaKENPuSD8H2JtATLVWmNek0DglhnMvdf3lT1QKApIJ7CrJ
n3nIGnwMTZtRnm2Cz5DN1UwMtvh+I3nNyoRnOI0vOUlRXmSkNxlFD8XU+ZoYE72a
wRpoERW4wde/75Y6fvnxMMYnCbpguDLrcmpd8H31kW2mxNcHgzZtHR9ATtMKTfdv
FJvdiM8ZssEZZZzv7FoPfZ0b/nkyOezDlfeu4zL7LYorCLMUVlRIWHnQAs+nn6JS
/DgtL+yaw1Bo8U8q+y2bGL9Fv8w5woHWN63GKk+1uTmLIeTUU181qbqKkiuP0OVF
5fy0ONLjRcVdnh4NP7Pndh6XPbAmGkLV8SvaKkkzvpWA7N4UM9hmUuYUsVwzIBgh
U4qGkxa7v8kAePjXTzjRPr46D2iXX2s54NwRpa30Kf19J2iDngFEmBJVtcqGtGIe
I6sn24pxzMsGfkxQx8E+ILzFzKi5nqSdRwu6FJV9sRpbKsZ2jJLw8XQxX114SvSx
08x/vyk11WUVzOFnVyDPnE0lBib/d6JJvJ/qB9vGiujKn7ZchMeqGyrQBGP/5FiY
mW6rpNBfu3zOASJCuEHca91tv6xirGB0+tf9mbOtAiWyWGNeDEd0fVg0RAZl5dLJ
zwlOvBqXKYvtIoGnfvauvSmOa0HZlI2kFLPXcHOXCazUojH4m/t+XKnkUbWXFkTk
0ifdwSFNCmeMbNYHMYHuVGP4K/tGe1moZ8RqGE603KYoFGpS4cMJUkcKVhlASJTy
llVbrCNqVUHbhxwENWndGu24UWJxIm9UsN9FqDQKcgDvHDM7/ErbT/HwOvXp7omD
dnuZlWQkVzS4EhQ0hAOpPALQAdMuaY+OwxxXUqS4G/5IAceoLa+H85k7Sr601GsA
vZnOBh1HXmnhMWoTnaRRuPqhSURo++jBNE59pWee0nscAhPqwz848sspUzEa4eEG
IKbep3S/C+ui3yfGAgC04WE3tMiAUNUPFfkHhOWNT9yiAtgiOZY/WWgkK2c2Pp+z
udoU1bELgTwldPzUglqMxd3pDriL+cWQGfVSI31v4RBrubKuQbJG7Dq3CGU8oAIT
aqa4TWOT4HXk4eQpVs+1ZJMzEKr+xqDhuZZgWDoadZNuZf20cy6NK4h1lJBdagE1
+XXIDnE2ctXqAqR53e2oJh40vZFy/Vzln/muiY+E5aWAz6YufIorR5pCsE0/DKeD
mucjws5xa9BNWvb70ZfwlHRE5Jk2pxnviMSXJGYeHAb11dxKxqpvTLlxO+GZ2ifw
yHruKBCXBe0ImG9V9Z7HnYFc4XtDeUK46aYQV71Mx5yOc4QoO88tsXvviA98yrRH
2/pxSy+3zfRL373I5yh3oeQzYrTS+5z5mfxCyUnObxKcuggE+ZpBWYYrxTSdq1nM
AGfrP7nSZBBn/h9TxFCazu4uEDnQ+aXhvwxAlfo5BwJFYG/0CV1XDHhkL6fGVaBf
SHRGLvbd6zbnZ1i2ysCB+n2mZX/riySo3+C/3twmaVoAXqZRhQVlekTB6B6J2oK4
s+2x3iAmBlU/FL2lPmSrBpHZd+fmzYoJRU8jJ7jORNU6Bd2VnU2RrZiSaH7T5opm
2yJc0oAmKNTaLUr1tFBXQyklGDZU39eplQTRME8ZAkZw8ljdhlBhnF2AEC4xc2SH
IvhKoZiMB8XEjc4rBLj9XZvBXOd2NBpun09xt4PXhucSj0Ld6UVKcXftPOT7k8qX
e4jRMpCfPYuy278MZNmlYbPPO33UIf28arX5OzOQiwmyV5606OLpanMvas18LDoA
iLdi3Gg0H6nUKF3/PIJgKsPXszFdlceOJMjBmW8bQZ0/TD0eXWLDd1HcJJy0Obhu
XRTvomoMJQFlD5lFTv2t0WdH8iLjnI2O1TKonqQLWfQ/spZxIlImfu0tuZU9+3o0
YQe2MWeq9rMyIihFuFUJnFbqohjODR1K6iiUaEyC1QZyApXj43VVRzBahKJEw/4k
QI7BHGSJa2knehHzGOutmaOGbpBdqaie2clD1pZLDQcM4QP2Y1zmf8PdYTf6nYzh
dAZbGPOu2k21pzGL/Sdfa++1fLpyoTAp3cNsagOiRmMDAHkEb7ldTyqnX5bBfg1Q
efIPxTikgaAm9GwUC7SlY8jHITUPCaq7FRqlk+Nb6poOujO98PVO64mWSAD+hpAH
dUle4/PmcMzjsOjgIinNy7EwB3mJhaMTC6xgw3/cJHGQoXGUrk8El+FH21uSUD/6
DDZDRAgB7/58iNHYkSO6p9ZuSGutNlF6RcZCdTKRRJlK9tDEh51E5hDlAVIzWNgG
vEFijwloBejrTFOdTtdRY3LrcBlGIKiMknWo4t3jl1ShJA/cIX82SxDQOUaRzsZN
GwKtl/R5fTbenlzE4d5hBgFk8I7LL4OFAByp/Bnf/pW6BMrCU5YHsKkyAv3PglGn
OAQSM8HO+6FCTttFtrBLEzocBsIRA8puRrkfW4uWC+mNeK5PSg0xV8+blkAKVl67
Vd4U6Q7PTqxa4dvv4VKn5JUOKCFkrIDGKrZnPhfaH+Wo5hREoCPGTZX40GJYzovp
J9M3yFAzm7/zNl5H90FJhJGfHBM/oNRPSjwMKFVQyekZ4P6RDh9mN+0WZ4Gbu+AJ
7JjT2qZLFqTz07HVI+wY6XkezXW7fdRMKV2BiqWdoo4D3jSZ0J1VQ5PXwq6qlYt5
A6tAf8/yYnBlqYapQ1Y1G30iqOiJOLZ1vULpaijZJfISllE8QQvnb2on01yEzC8k
/JBVGXlvNMkxFc2VPimpuqqtPSX/0eWRQ5wjVvIt1UZa/ZA8Vb/qZ7Ajt+Swk2eQ
aoSNIP72K48NsrLURYvhi3+EPmMC46ajgLELEu4QvosH9plUPpiJK2heFMSBkppM
YfLO6tAW3evfreJEotYnMVKmEs4/4/JUwYMaONL2JCyQ44P5X+soVYw3dz/Iwaog
H+jY5PpHqX+nesi5ldM7v3QKFehsUBsaOr5jeboPhwgwKpX+8l5/k98GY1dgD9GI
kiEpaMxKOTgRtlUVytxYorsVT/eI0K/odHPbE/IFtXC906qG7UTcjERAyDxEaU8e
yndDNALAbYPFPhbzsBB3aibskZCloUtKCRDg0K+PQCiv71mLs9Sibyhaui9IcIrw
u6NWcjF/me4uNkjC0DQIuQcFqkwHEC3xBLtgMty96xelWqn8ARmSJoxotY9TzpYY
f2FuwjkQePgUHkL5Xvm43kCowtXFiUjlZkfvrC98XX7bzph1CxsZl5z1jj2aHX+F
l3qkmHjyu1wkmxpnOe2hk6/Xs7ODlNiqCXxmne+AcvpqQmX8Z+oR7ZNnW7O3Lj23
acgXhkkMIRTCpCHIqcVQVa3cozMESO+e6JJBu1ogb/Y4o/qstRwU4grA5FRPGezn
9Lq/pRi5/aQYTB2htAaGVdbRuASyYowIOR2Pbu0wCBU58YMD2JOJIEjgGXhjlTIp
DTBPziXo+Sn9z8qGxmmCnETB4Ny96Msyh6XsArC0urEKEz4ZMMpSfuAfeLpc0i5o
tvtWG+QNWFo19hwepgQ+ecXj1Kgx92YoAqlrBJtZotj2Ams1y32LFETD+E2Ch2MU
3YIF3/YP+OqrJJq5zIYp6ummViskyjoiMPtJEVJnTfjDHvGhBkgi6IKOv4dhyEUB
HAgMj/YDMgvhS0W/N9eQtmZOKUWGwHnOeIrFyP4C7RW8ux3dkMlh9ddO1FKNVdE8
SMpmhH4NaBrRDQ0fiM7tevnQ31sz39q/sm2TC7bYaSGGBprAkiPXAghbcV9Q7o2B
xy8iqXDR8/pd1P1nRxByUnL+ClpNoQx+kLIipJ+Djivs5daLGSygh/lQ0WpR7V7F
1jXINJc5tWeKnLEBYz03+5njoTOHTtVqhCCQqxNvJBJ5lW3LeTj+ZFPbrafuP9PU
ZFoJd7RfmxBYWHX6e+iv5gJ/psqxrjQ8EulIQ0Wkn/1rkit1ZsCrj5PxziEHbTve
VZcNE9ZDKLiwP/kVlJGpDacV0XphrVqEG8NQy4QgOXazcI5ZhMjDkd1aSr8GPWqL
wHxH8vFBNgxgoFtpnduDcfsFyZqrq343RgnxbEF3FcGk74ARhiMmt2WjQwx3+Lt/
OirK7MbgqfGo1IlWzKQTIz+dPOJ5vIzB/qsah087IHtE8IGHzOP+6eGbloSthq52
6+hekk3j4vmHlkYh7g9c2QfkYrrN3WczEy+f7F2QExHn+mRUUXP8r+6loo9kDu2N
StT7i4dRCAnkcKkMOKysJTPV54YRQcHJzDba+8GV1jXqyTM9kreXl2tWT+MKsTHQ
nYxjGc7JEV+E+GKtMEKQ3QmZvqu/MoDOajnJRHDL/FvLyn7eEq+rBTR/AyRkkqCl
V84onIddhDTDIm+R6aLjzt+zL4ma/R84NjT//SAtqOBc4HNwCERe+YySWQuampGp
e6PbBYbDrdxdEG9aERmFipfV/Hoc5owKx7NAYXPGRxHIcXWEMy76bwb3U07NXMOL
OexSVWubZigNdWX6KAOjS7JuXHOxX8sg2qWwKdzdCzIekak/eq5vir4Roj+VvzAL
CSD5xUrNEkJ/CIp6P9XCjPQRNmR604mfh5ZlnUOYrWm0PpgfyMKUzB5Yxk8+MyvS
BIZV3C5UmFfBpFarinn/hNlkf4kWmzV1dRu42pZgx0P4ODw8XMby+H+XxKBeupSX
UQFxTROnGf/MxGcrqSbpCrpNRvPLQisaGdqPrSo4sOmSnosnDyQTpXzzkwewTEfw
CMAWuVzoT/KX64sFpzHlCVN+Xg7iUFnJWTWrU8xCI2kEHB4sDPqkWx5pwjGH7vOc
ukEhazfzmhIXtW27XDQAJmrh5Z9KGnRbnTQYxTqn7rqBH1ECA8LHh8KVXuvodLs3
V2d6Ia1a8N0aXYREiA/StmUA9bG15xLgQekG7WV6e+JlE8ve343rGnLtJz4tIfEW
paxh4eOJeTgSsbcdJI8g7/ceN2jkZ2Q8ArLUHLx0df/Y91NQGft+qs1W5xVggkAn
EBFOGJhLzW/dXeCr/8Rd0hg0AZhYl/OhdPFt6Y/K1tfaVMQMuUdiN3V/Bz1+GCNu
Czrnxxce8Ima/NjEMClJpHUs6T8A2KVXQfYLcBMMWTg3kpisPqx6qaHI1qxHqOpr
osZh2OfP4jK0aG/NvobqHM4S8OIQOuYBtUFI//HLVhaCN2rG3ECOUXBQ7qS8EKkh
PORpnANINedN5LZEW2Rce+5v1sWtfHQTpAxdHZzCGc7vbcn7GP0LyASzy4tMnINX
WI84GJC2TMgzB5zqy6MYWl+hd2qlejrzBJoFE7CHaxR/2bbqp4Uah7rLHuNVYGce
uiWRftqYsHov+Hlizb8hVQYx728Fegjd6n+MyW8HSPbJLgWMNJxcozmCteluWsWt
Zr3HBAJAknj8NMcTuKdosQ1wQMmiPR15JO721QMULfC2mC5B/fywg4FM/84n2PwB
zPxSial0yQcwVSq281RCYKMcF+DllrYj3In1YZW0PpYiMD1dfc7ka5FY0MQ2etLH
0eZ1Bwo0AJGnQFo96EIfwZmXwtqhNCozxuNqKeLMs86EUR1yJLCzzmZhv+R3xe9V
zY9j5ldBMJQvaME8IcLaG/036cTtKeADFn5l8+lB12HrH04oFq/JoiBIOEbZ7eqv
22oBcEO9nbPWqsuUAlEQSR8z04YnpSswNvsYkBHO1utoBdRrdTSKQp1rRTNvoox8
/R7/V7YkpKhRYsBSWXsZRUTLGRhyaxe9dI5VsVd84DflHmXtzMB5OHTXwg2TKTQ5
9BIARcKwd6wddYFFEXxdK/rt8vJPZquLBDOz2C2T96RA32HA8+7dHM0K3LrvtUTn
9kQyTOmQ7vV+Gcs+X5njTN3rus+jB7cvMBabPeJWOVecQaAzIOLMxfyuy9sLJ23o
GzBCUf7Z5Y3PpGY87hI7VApuLmzSfMBUlHgawcTCyVA5ko4rVGKVMo+4EMHmvNnu
IKrUQSxbYV8XFCLBsvyGjOJBo4MfI6OGrGZNYp6SmCxE1kr7aYf3K3ftKG8oX0tj
80NEgVHAzt1qMyYNqBdo/cWnWQtl2Q8U+VOr9+/+cEPL7PMBOWO+BNgKEhLIPdgr
0not+zSzIv/lv7QRk4VnEpVrrMHZvkaeZAUgDyYDQ+p1kayhhCa8IWrxpROMcMi+
tEkxnjRrzf3rClFts7vcBQV7TlovtSFIiIJ76rOKz1FlznPO815HRiix5uElCp5b
+C6VYS1DdE4cXRqFlbFBXjBT3lDttlSpv6lUgbjeObux3epP/VvyV98jlkYpZYJR
QqgOu5VZOoKbzmViOLycR5vj+rTcNPt/OPon5kwgT5EoXlP7IEPnjZgpqfe0CMky
563h1oLZc7ntZKEqmR84YooBSdtOb9uqXgY7PCprfhkHiUx0xBtcQXb9FeY1P/n4
EwV7dBojbgiAodISI1jVnT1xMBaWqIAukCJepr6u2j3tl30CpyOSCzje/us9wq6g
1ml0hZxcv6rWWnddSQCLUxNSu6Ln/KptuZ8VKIvZ+rIoZwXJmgvZgOXw0CI2Yqjp
LuuZG76GWSqCTjRMQYLQy/4Ma8byUcG97V37yDo1dyrrkJSmYEMhqw7oobvrutJX
c40058I/uyNBd1haq3yWnQCI4fzMd6SbxfG6TdOIPyfOrCdeKN89wxXLhxRXWK6f
J83e5D29N2aDRLIlX0yehKYgRgz9ihtcO57fSOc28N2+v1KD9YHXgobejw2XDpgl
BPpzjvHHMOW1Xnh/7CtFt4KE+yCdO3saBgKvkCBPeLGqaeN3U6iY8Sg2UildNZXI
7w1LgNR3jc6SZKO12lnfXkpRd+mex2OfDsy/ytRPelA4RwvdbWGFHIlvlSCuFgvb
8SG7euHYdGjuRz+3altvp2VOhvwcVbBLNXMsgsXS7bGkNqpyHoELmX/+ogYlI3Of
3CJ7rAZnWs246ogPrBq8gLTvfw2jzkfQi4rz1HUkpecdtIYpbOBWOzKstL9p0ny9
3/aLwcVqzlVBiJDtgpkNcIRtSQVyi1ALDrn5cy8Srs+OhfqG8qCiB8JS/fQKo+LG
gzPEIqrXJlBR0asJ94zmaN8q76GrXtEGR/TaHEP6PJkx++lt+rT4hJi5mgU7EjwH
6fji5VZRPMdrdUoxxsQjEFLdCocXgZ9HEo6lXPDh70+XmzNkHbtuhxPxeV+02RBf
qxLbJJUXYY40JBda5N2FLvw24qUSYIKetGr9HyBCoxZxkQ4z/KrK37/HvpAq6zFe
gvfHNpskgDINXiJ1x74DmgM2si2Vip0IXO9d+tElBTSLYCcJGpXfaerdYz3EGjfa
HA3XTplC0arY/Z9ui90kc3FObIteHgw/qK1PY8KQKYa8aXCWQ/voXdud0ommyppJ
9AIL/S6iPO+yeiEc0q6IzCR0oN1HEDDYQqW9Lt0kV6XJys/ezge6cIg4PVFj9a45
LfUPpF9PA30Zg2J+RlluQ9cBw3d75S8bGJmxMPTyBxsGfQ/FaU/l3KtsAMRODR8v
OWs8k5ESm0uYGNo0WeMiiT3vLRIO1BmWNvetrhZPTo0Dbxnf9XZX61F8PHNGalLD
Mk5E989+QIsYteKxGqGhgA0iZZjoGNg4pqWkmearWFzVyYtN/WzHwV4K3a+MS9d2
0AjnVfmyZHfU9KS23Po7VsKMVNAzlVSHF+2wgc4lGa/EPDQ8/T7hIuuz3EBOY+3r
CVdOLGApZhNUK8TdhyK/TumVXrJdTxEukHHmL5gO19B8FjMaUfIy7W3fN4LXgchM
kMSZrxjgVSI89SSumc/9VmyGChe+xTb2SuOL+qMWrcwfs6cKjLGgsZAWA6ln0L54
oQPaySjLC2qf7LkhQx6oSOPKhmxjyQvEJ3KpdWrAhbZ4Neueo3JQPauQIbTAMcfi
jl9G6x49T+yTvk9/Wc1vfpAIDoBVDORjiNlO1XdC7Hn8z1na4e3Usd4bHx43K5he
wKDKs3Nm0RAji/JYCSJUXqGVsbgvb5L64wQzmcm6CX0lYFdLTHXpkzE7roGHmW/X
IaaxxedHmh7tOUv6l24LPoBQBb+z/L+tiknaPxQ8Oz3NhhOEqXNqtuy5L8cUHHfP
VESHzwSitjyp0C8oD3Nyal8X/M45ZuMetLWyOBrqgd4htOS3qMsUBmTHYMXWbq5J
9kOD5NnnLS5aHXN5IfhjuPjvYbYbyuf3AnUadx3b29xZ+HIV2XUw7z+tkz2rfGgb
/W/TYX20usDbNyA9ObtNuqvQD2nDWGGb2GDm+oAiwW2dYSMvju6pKLd4fKt5dDhD
gCYOPkEuz9TnsX4aLsBH/K6Wy90+/9SiuHHAHsJcBwO9++q5HI2ST6SMQRUwKLZp
qwbG/GFlRp0ghSLPNGvd0WEbCQjb1kysh7cxUaGX92XUGfHr9R8xwXamKsLJhIY2
wEkrXsg5ZXZyf4LdUFPPdellR2UoPDwsIMujbj9wUOB8jwA5fmqJ58zy/hAh1Lz4
Yw9c64DOlqePQ2vm04HZ8dXV2ltTt60Wk2x0Hs8ZupYxjHEMb6A6XUes/DAIiPTz
XMfdkOd0D996wxFmsZJAE9ESJbTK079bRv7rnwIn7qRCC1esVOmyil1DPGJcIoOJ
Q0VefgXRUfCaZTf17Vl317fhLEskissUP1G08PIope/ebpvwxVNAQK0H8kgBjIDv
2VguVKjSxgaDEcpbzQD/WwhB+IaMHxjnZXS9yWjx8yuEeXSnU11MQnjf8VevHMvu
BV4ZcNv0LO3Zgz5byjnzsLGGaLGRjCiVbUNVsjd93nGLg745IRloaQIpNE0svSlL
syiqqFjJfecmFyZaBnVa+4FYiwZqI6J6MDRaS6/c5zYEBdcXOG8Q0Mc3Vp3D+DNl
V4PFSW1WCZN+AG/3b2F2Dv+Bdg7rQlbo+tArxkTnmate8cpAxj0DIDdUKhv2uiI0
qMqDiuMoiTcivmA98rfYgBxMFfRX6S9up9OxSRMktLMTVo3UVgfGvfvSY4LTBSC7
ZTsERKbFmprSczBRCosk4CiV1G8yhguQZBsolF4QmL1QE21VgVo7BzEooBTp0e55
zrh8kL2pL2oVHPQTMnZ5w+whxUXuPBWgfqWs0YoNuGfUGAJkmmLmO1ARneP3RTva
Bqp0FPHJIBGQv/yzQJM6mGHyawP9ZHClgpHEMWYk4/ccnIhVQztLFaJsUQ0mNE8l
aQfWUJPS71ajqElEyFy6dLf3kPsg6XDyl5PRSXepugD6bKGpgz+R234VbuqpXJ9a
NkvksAXEQlff1RTb7YcSEv3kSbjV3DTAl8nm22EabT4zUxnbMJO9rg51dHgTJwov
98RDqv0dlOLOwQ9krKlWkErEpUqaIFsJkTamdD4zknK032UKjfsx2FHFVbvv/nMp
9wpUuQ5wDqcow2PlTiM+l5Z5MrpxwpljpQGu5AVdp9HEBSdI2oWEZJ9dmsTcURfP
X9PQv+0Vr5SG3HPvEy4n+ox1CUQgHvi9vATTs2+cXnmbm+MwZ/CwoY97TTmYXlV0
sb2WsFpc7J8DT6ePLQb5G2y29qXJ9laAvFkPB2gRp3VABlU5ezEjd+o343O/B2gg
qVK5l5a/2tNWBQbGhlLjm/xP/9aF11Pw52G2fsv06B2C37TN5pIIxuUAYzLGATCH
Kk5CK40tyi7OGsYgIetkMp+NZf+ti5hAIc94XgL7SQ0aHW5H9zsL1/X0Q/E5Kw6n
7zPo1maxd02DwlFZa665mLMAcjpconGN7xJe/cjkQP8MTeDdo43qhiMIXlYyDIKS
1ZRdz6iDdESg6OwKXhyg9oiI0/SbH+kDVYCAEo3dUWZRDYJlmN143VEwpsnVxAaX
z3OgP56eYDbckDO9LY69rHPWCXLZHPEkPIz4DoyzTQ2uHxta/mLwXC8gc7uFy2Nv
JJtzUEsQHp8JnvKaGk3RivlEwZDxdfJ97VdhxXjPz5h6dq1T64ZJPE9OKo3nv2aY
tYzc6pZZcfu+Z6/rlLaUmhxxd6k7cGOPasfEba/SWzRlsaP0+fgYhC0LL4g0ZqQT
uRAdAvRZgujZIIwKjqpw5S/vd5+7C0wHDnyUrrKAw59dzJyKEcT48L3mitHcFcrW
rNci2pzBo0R5tYdq1PLfwOQ+GVM4tzdjeKLKj6uj1SY8ImEaPFhAEuNrAUVbvlk0
4S7gxaS7l8seeOouxjRX5+dgkvNSIDgyuDc6If8rIHEf3kB7qIOgSB1Fw1L/V5i0
tMMu6fkYqSDQnM3IeSERd83kRJQaYY4GCdg5Pyn9LP0oL9LTHpSbwYVHrBnFFpBF
xPMqPM/Yc3zJYuHIg0CeKQJZamteqDnh9lxMrK5EK+zrbzW4kqw1SVnepVA3AJRH
lHPX7LIPRAecMWddjo4vsu9q1iatWqbAQFPlR5+LNuBPvvW+2Bs72lk8Kkper4wn
cCI1wp8jhiLiJkNLPkWiDNfxxKuegahrB0OpgT4HhXj1eNL2Fq+VfaFclVxaVRQP
wPYG825ZjHZrBI0+OOzNrg6Hkeq+hOtsEB2yVy+fu/pqStS+dZhDIN30avPZM7zN
IywLbEsYvsiowQg9zbETMP1ETCXdwDV+bc+vsa7zBRghJeS6ZSsaAG/PgrhTKDqZ
dYPvsxErt2oGDdVt2cCGKL2XjVKw/ACE/zqhD/LIle4C/SbDgM00UpBTGUSRGaPB
JqItwr/a46WwkXxO7MlM4TH+ep+9QtDeV0BMbgwp/MxE5p8VWddplnCTksgjrQtH
MqJH97a/hpI3sMksbyc+1lDz5YVK7bxbAETWIOzs7ieS9j6ACWAnYJZeAw0eooEk
ZIdaaUx/A19RMQxI90xfTLCk6DSQa+kWDo8HP13Ibz/q9uFsa02VyE/8fI7x1DoA
bCTWxy6ZkQLlfKbDZTBi9cHO+TfGKJuXNpuUeV7i/qXWLlJIOMjIyDcVAV48EIJw
+FxToUjbOJDjpCYSoWqMWHB442deM9k57/90q43Eskug8K+uvgGDgZMUeCdflpyU
ut5HcHA+9isdgEG3PgAlDmmkEvHIGhjx2GPM6uqWI8OapjUCTvGZJUE3kyACmVo8
l4rIJy6ivEgLX7n+ChSCcJCX1BndnrhoDjcLdGi4Piy6qwx9rQ+0V9G0eTj9puQF
fH8R/4fPRB2+MV9rdSW44dqBFSLf6QuTR/0Ui+gmGkXJ5aAhNxydIF0n1/JzOSOp
vacPS4dfYpP+OSe0q52p/smLYZDJxcUCrC5GRTSsxZI8YKiFRK6f602Nac0M7j8g
89bqHNgDWeLRWtKudXYrxDs57MNay0J4yyXR7hdNb7r+ePHnNbrwxhGY/B71DVk3
upm0Q6mRcKybKdYwIW4pQL5rgOhpUnFtMZDcP+TtN+NE8zJ1ToXpfV8vHZkfWcPK
pSe2iiTahICJmo5TSCWnGclUocb7oapEC0N0cWSO2r7T9z3Rpcn5ClwIJy9/Wpgh
1/msQ5NdY38H6Q8TTkVG823eC/1krBTxOFfHR9uTquj77RuVsN+YWSWLedHc5LRh
8CEEQx4H0qLdsW9RwmiWyNdIYOzHKamIiFsGXTsGZLpjudCDOB21Yxd55xsjLlAs
pDZe4MNzgPn86UO+SlrXp4N4sM91Krd0Z50ErDC4loFJtsm7rrEsr87pdtkXNuse
Xt9DnX7CN4yZIIeBtfpmgWhMEzFhA21Rc/EYeNJ+6IHtY4EkGxvikng4/rTzPbOY
PlBlUqbkmtEr0mNnAAnxb+oK1EKEbKwrQjPlYtX/3OluY3+uGmJ1E6CBuErq1fNs
eytJRhjJNqfBGxv3mS17om16qpgyPphZcIq5RPbkLdm8qvHUvX16wrUgrpNZHMac
oFaeI+QDBSgVY6tSd4/7+nfCP+jGuxjheeEoyduKzbkYPbdvSblUtr/zbLG7e+R6
GUoyJ/qADTkxbcWq3e02HxPLy9w6WqwyTsQhzinJyNU5wsLtmBiyfn/4TaTI6w2/
l6w7OP7ZkJ3H8F1lHWGKSMUJsZL/SRFG/D4joRAncrHN9cHBgIEYEK66fCS+07j8
f9JdNGOG3mSnaSxuPaXwrDiY3gah8ENHr4bhG2/w1aOZa1U/lDy5Kxd8w6R0YgSm
SjxAaB+HmxTYrKTtqJ7EoTSTpocu7zPZ5lOQY6kcjIuHp4k5LgbMaRRdctE0xUCV
/+w9r8cvokG7xd4/OASEK6iDzPjsCCCYE4dOBZgcSRJBVr5bu2FW+Ke3JHnDuV0D
qsRLrjRNMlxfVcifqIOMMhVLE+pwSqgMsXFRUitHu/cMljY+oElNGP4X+kxlwOnJ
/mH+daBLetMdjVzVo/G4aBT2VMRnJTRdH3bCZLu/ECEaJe5Hs7aT34x+STTnrxY0
of7kWdUhv29uL8WlchBf2O6Ki8uD6iyO28iLyH1QMkHr8MNMllj83KY6r3eR5mAt
HhQZZrdmof14fJ+d7e2M7dQIFsndawmFkCHqmrI0l8S7W8u2f5FEDEOTxeA7jxN4
0t+Qn+fmSd+WZFOCQO8iRWy+q3qTkZOrLR+YhZ/ZC9tXLGTSAIs5xeA2aI+qjZdX
XKTBgoPZ+twn9d21ViPTYbPaRQF8UGFHu+iVQjFZ5KrSGrHB0facEy9bs6xaxXHJ
MlPGCAgUBvkxaGOrjr6/8n/IjAgDmLe0YKt6n2gJd3H+bsOUNMPLYMGQMT3aJ/7G
agZZVDvIqxRr8nXdJrhv9U2Mt0XCT5uK4uq0xgU4uOgx7JYpvSg5JtTOBlC+Qh3x
GhRB+NEdS3sk1BX+a0ZOccH5CXvO0P6uOZZ/eDe22c1EHRAwDm4W9AaNmrKBqyTN
BRPpHu3VdJSDfBRPO07qtZ1VoYGUh1Ilkc/CZr7DDRVcVqXAgrGti5jNG5meViCO
8hwCbb+zw45ZolIy7ewEui+EuiIPV/vkEAx+s/r8BX7Xg9m6ZPIZOgB2FpO5ktHZ
+hHRFED+sZekM+MJX4zQPFZVaH4f6i6W7Ew1C3pEpf61GxMs1P6OIJrObqNhM6hb
tFV5wDj0atrSJ05pDB3fJbQGuDRsUtTiOnIJ8t0qy1IWSh5YaUv9u27BYL+IIcTU
ddOuwIQVaZQZVrEq6WUiH/cCzVS3aYfZpR+LGOwy87sSofALTwuu2wD4PqiPXwDj
Keg35ebCi/Ed7HFTXc5xW7bUFB1puOuaWBtCfIMNzVOAll7/ur11DWD2PMQSjbjA
I1ITiGygTLpe/nZNeEaJlLBrUiV7gl4qyXVeij3rQkFZzI9gwBNu3JQpm3z2SDon
WhMVSpd3Tdn4CtGjGqxmGw7uac449U6L75XquTI+mMi9+7x9N2m/vLdWHC38Q+qQ
YQdalzaC8HF2Lmq4I8QoEd1Wquso0we5V2WqEtq7VwfjOhYNNTCY2xISW5ICyPv1
UlOcNuFkAusopg3NcFQCZutE2IDHGg+0q661BLhov/2vB1aOZqGugzKRtn2UiJaX
lFmNdq942vbv4lxsUrXccjQ7m9XZQV9JB2x8DjcqrRP546ylwMe2iAOPqVTASsFH
NlLh59yoBpIXDEC9cPAqmiYRsEI3j5eH0+0BR+/XOIaL0M1GR3DIK3BrHNIq3AN5
1EsKsjEY837qNRzUzEg8qs2NkMwqgjQDNdwRtpUxAfD8rnltTvoddKvtWW6Ib7aA
IdOT33+gA08TR7+fy0uaNkfO46Oz3gU7QBnSevTMHQiB/r3TlppiUz9S0TswmK3B
kprJfW8iSZxTyLy4WGVrksy+i6U4N4S10Dnz0urV7Fmc48iourzq/27mxPqnCPvp
p/dGXBEdrtqWtbi7ABKCAoZUkSldTr4rh19CfUGt37uqTGVnxa9l8tHEAtxB0X/u
/KTWQVOBmsJNft9WiYETaQJeiGZ66ksKIzI6oO2jbtKl/Mp4XW8B8FqzDoLssCN3
4xvcAp55gS9kDMbuqI+uKwNXlpRPtLGywXHmPB1HdySmzwbxO6UQLFYf+V9GbulE
AYbPPfQIHztkTfIvkf1pOhm2GvHAn5mz/FdLqqtFqoUy55BCriCOfNOgwG/Ty67W
SrmPCaG3Q8ZBdpBFRRohELX4BrkBYSmtQ8Dp3dwD5kWYJT0S61c8XQ46zH3Wudcp
8NLxi6S4zznA706fdGCVxrUy+0J4REkppYGyJonozQ2+bZ4TqZQlS0UhxaTrZgYB
s/Ip8lgO7knMGq9Xo8y5j8mEw8Q9Yc9vPEVDgM26rMCtowott2eJ4IGDyHJ7217H
PxyPXsG2z0tYovFMx1/X00RerUYhU9j9daJEPBEufQPqnE52+opnquzjqjLS3VuM
K/TMbzO8paVOGdUQX35Jd80FDedbo2KAk/TKPqFFl4aDlqq28MlBN+P66a0tgCBW
G4iLvp80nO1skjnrikVkjWnGwAwB7tq1oKVml4c5Xnh9KRqjjkYxUQV7TlLgxWVk
LX2hPa5qAcKOOOQDhgN2o4zdqr/V7vLpt5WshNwULEM0zPCTnm4sApRs3zhr+2gS
X/oy8a6sH+5zjFvxmXqJi0y+ZrXSIhGpSPnTMv0OynMgv33HntYJidyWxEdBYNQ+
+mzt6DZWHFzrdrmij8MuTjodplH2s7MW3NlGavTyNnWuwWKZGbzYHq65gJ/r9/3h
00veXCvaE9NsIbq8MIyUdYNOEJm+ceZfzbOmfRnGqGJIMTEoqoH+Jk7NkZQWMlT1
YEM0RdgWPOx7bwpFzyRk4PSo0b49AeUfUa4HMBBC7MFgKSDQC6ZwoU0j7hvMNFQp
XqmLLC8ztmk8ekXjP4UEF45sDy4IVyG7I36TKqSYGi4oijEQhTNNgQmvVh3xpDGh
ikn70eUHq/PpaiXMcfxHvwbZh2+Tx2hc7w2Ii9XXH0SxETZ06hyc6XqcLTVfGt6h
WeDx6fW+wJM9GzDyANUfISPHKGW7QQE+/mHaSbMUhPjkAAFbfo7TaEdHl8iNStzD
dqrojzy/cVGqPTFnEM6tSBEXHgzb176vkgtHbI5p2qN09m//5onuGzWUhnvfpdfs
Rql9F5FleZdMdfl0aphchcLce0R+tsNNKq4CHGp/Fdp1CJTHXjx5DPntOyUd51Zl
AucbdpvPzd0pmbfDq4bqnoOyeHvuzbNrgZHBATpfiVQM454ALg8BngAMdbo23KzF
Lo0+IvpqWcj39cWppUONt7cG5yM8PRXBB71Wpu7p1of8Rs+zEqja8JwcA4wvK2xy
S3klbS/p2lWtzDlAeHnw8IXEl1rHL7OHqI0OcTj+vQ/GpU2gU7QPPhglgI2iENt2
Gi3e3C6bDGa/iGItdx6xiNlLZ2rpiCP0fzFLY6i4cdLKk5xgta7vPi6KAp4h5zIL
YkI5XqT4MBl+fSX8NTNOTngIxQys8Z2iOJ5Qc6APgUMMSdHD12gOzZufIuv4PkSE
bdBLMyXoX8B2WFJ5kWXP5o7ekrmcAqyaat9vWAPYmjltyVaO+dhSopdsmB1nT3pA
125u3JRKdl2P0DQZv6wBG7HU6JfkeFkpHT4jIQv2U1ej89URI4T+OFm2MVojRog4
DDlYy2M0fFQhWSi9f1Gx269XqLS5uohhtfVaUWmvPEfBJBpjbYMtZldrjskNdn2U
gnwqAGqLyq8PFkwCrRZNoQVxqPEX6/YU/4ZLfnrpDJfU9FWNNuokvoV7Abd1QBuy
ouwmTzI3Ip3vDr/JMw0uHon59WQxa1TcOJD+ZUkRJPEXA8XB4JmVef4zgZ8Vn8VC
xPF3hzV6qqW/lwW9p3s8IuGz+I60+iaLxWyxXddgHJNTK2g1AWs7ynmlE/X6PK0U
gZeow8/wTQ6v+JWMOPPmLxIy8ltVb3pddXKyfj0Z1LQwxrMU3EoZaCi0WKmVwF7G
GqqZc2bX/5vwDMEnWZiupQgYJzy1NyCK0JN5xuVD7NOUKB8Qe3BC0X12p94/jaMC
MrVwSSKM0RZJ0ikg217FBKv0otG5frihEcmS8mlA0gEPPZ4Mcjp4pKO00MXvXTE3
DEPonUuAsYjEay0Ld8tBaDRG1pYfOIsBRLSZTdW6v1P3q7hW/OBzNopUQII3AHnS
HrfzpcVNEZzQ6L2pWMKr7OEHYTzP6831SDrBVkkGFzjE4McBV4nZGbRyNPCTy3KQ
Ty6DVaCzaRVNhUuOpTWSoLZX0GJh2m1jYo82OSOK69pIsXpUw2raincPm0Gaoy8A
3x2GiKqejaxkp6GZBdbM9cghBbzfXcE/cR7TJZ7u+Bsqv4D5Fzq5S5ZCs063wL/X
3Bji/Sl44GRK/gcqeBYFxB8imx7Ps7Gwj6wWRY5fnVa8jd6QUfioA4x8rdRTWcPw
IKs1D7cOl4EZuZ1uuQxslIjKk+lBEJsCUQwSDKe4qmWF7UXydVEZwmuFy3yIS2pG
nbEMSSW6/+z6KGH/VxLU11XqMVXs2IeWb2dtvhsBY6JOuMDIK+vCqxhmU3xBtv8E
39EdTDY/NNeoXC+YdotvrXvjB8F+dg7Jr7SlnnWBYGmxYlznc4pKFYkI96RXlvfL
0Bsv4zkDSHppXHWsqorZDSzNgnvpPYlA6Mst3efHoHF273KmsGu3kUsVr3dApOTG
gq7+4ja0VEaJC04H6pBEZE5TIhPKMOPWO+LEKYIvCcS4cH1YSCgaNZXaa03+iYkE
9nCLhBV8vCMdPzk40buHNYPjJJHF98s1WozJEFPXBHYOpGsSy02/kzWzitpsqb2S
16Z5R6IP/KjRHpHtWl9pk++n/ZuJ2Fv0ceU5cTD3U4PxlgfMnG6/lmY8gwNHWGR4
WuMqTPxy1z4FT8maAPStScHzM1P6JWJOY+mMOUgDBdoWHXwz38WkuLuETAes20U2
pqOp0jS1L54D+WW67QMVFczIwrLov7mtKm1IjdpMhKYIUkYBmhno7QWq1oQqGYXF
KMH/gnVU7Z1bnAPliYKB2WWlPjGGpUmjjW1M1SzRiQezf1prYrYcdsDa+pBYdqqB
M5cLITYaMgl6UQSlLJwg3QHyR4Z8FSe/mXocJ6uA07Ae9E8LHImOEPddUJdZgZec
gjKZakgQtSLB05XRwfjsgFMBIFmVxV8E8I9mdTaKbbHcPi/6/+RT2iTrGgo3rzIK
11yXaZNlVrnGq1Gz+LpUf/TmdIixZpkAZ+qFQTnm7/7qKV8IAVwEULEbIeR3lV8q
sTg18AlFZiAcAm2mJtP0QoDosg/qyn2ITnyW/9I5r4TT8g3u7ok2HxRilPDtcN+I
P9+ETczIY4/y7D0T9tO9NnHqMHgfFVk/MzLeorJoGBn1r0wBITzgpDoAv2BwCZHY
hgo60lnkQ0WPM7GIuKfDH4bJrWbl7GreJoY0WEn+qJk9crD5+fsAAkOiBCnq7GWY
USSZRWNWCE6C4IEVaOSgoS0R/qRpvMKRgxbRLnXGoxe7IVY9F+BV3OyPC/zzVKzu
/pfDSdhTipSw0LoO2RdQxHuB40HR71oXHofRnguTq04tc7PufmiotrQxsJG8J4r+
2zcE6qSvkhPtweQfHUdviJOdu2AOQqGwJvYkNQGZcQIOsbajaanvOdMpcvr4XHvE
HcyEfOhXNiL5oxHSv1XRNUU6VcBolMlf9AU49RXJcva103AIubG0OVBqT66CY36V
Rn4XAIUPZdTKSozCmG4C7lZDqbOHdc/mkMVJiiC2UKwMNaUC9trjoHC0v9Xw3Yw0
oTEdv98/NZB3/sT6sGAvx6RwFlwf9+lF/kNPakrU5LOIY8xZ9wiHtimkad9tvUfZ
voFSy47iygbO0WH5XB1FfjhD2Fe1cEizSuq1N0lHgy+StkNB9OM3iZmp0dBp0VpN
Zt+gTegXOe+IxIhvHcp2io6mSldCT26dlcegibQXrize9e0X/6R7+FNdzCQHwV+a
sigc8i/yyBqzhXFHNR0iudAqZFx16YG2TPPSKjvXFuUEddzcfHV73AoM6qYAgrSN
8XFnLPWOXJta3VU2OzoYmvhI2e2+32z85m3DLHdQY3CYQiArsmzpZ8tHJGYAK2ym
Y1KYtTAFy7niGH3Avhh2CYSZ2NKZrX5nmMqtxYXvqPerCaz+VBugEdT52z9C4XYS
IyROIVHgIhrOJNxjREhMa/ICVS/ZbCqper4ixZ7htcnP9bKJvuDzz2XsGhTRe7x9
E55WADtfh0lACS9dGWhDUyHcLu0Q1xoX3bElCXYEeFaUaKEFOZwOL/RY3YEIVNq1
9lHW7g9Pwb9Ib1eU1T0RMzdmWQ9h3GWAo96zoHLgtRksx1FhuGHqMPUeZ9oJLy2v
/KLvPiBK6dKQDYoC8xg4ionRSDQlaLkIj8vNis0dLcVSBCopIN31m9KhDidp6uiz
SiEH8GGcN2aH6Y5IwcxX49UEiEGb0+o7erQT1PS3okssGy/iiKL1tu3hRQY1h0SZ
98n4u+yIg25mcGXweCpcrBhwuFslPXAlFDcj2ojbavZyqzd2GOXlazlHJfmAcUQD
3elVQEbMu9N2TkgMUfs1G/PeoBZO/LqRLB5z/oGRrc13y/b4c4AV5E5xCJmOi5Jb
A0m3KjWGIh3nUIFzubrihVpFifRrKN+f/VY8J0JXQ80u7uSfIJvNsVHZQM8Dzxqd
GQPSniJiwrVyNMxrgsk3ZPtFwWOcJ2a4vKbO2ftYnz0F02nSRmcMs/27gJy/MaC7
yskNCHRahCpk2newuZXqWTlD3YpmKHsQovFPw2zFz0s/nnGc8dPUCNaKHIG3mEMy
boeHvUzdoqGbACrylWT3k5RksdihmRwhjwXeSoYrhFDBt/mhmiqFYIMOZppVitDq
85iFYonPdSwBpJSuC2Oc5EJI7RL6FFZgO1zQyeKQC9U5Z8r1fHQc7E3Em+AhYpRk
LREx+boSZyI8HqxEeOMO73QUACEIAxT7c70T+O7eT9CqaINcHDV6hmbSdcp+ivTT
q2v0xSDdtu0GLwMFGuGyIEwBTT+4FNfBZ7jXXubUJAXsPSK7E25gpLXQJCiYUS0x
IUUEGAb3lBmAmUbdgvpkgiKJ+bJrs4wXNk0RB3TRTOEh2Lx30LQr0oF4dy6bqJRY
6A4KeeXRkv0/3iGN23h350Qz2xqbMNBKFMjcpCyCYlViUKPDhldabrihZkYV+ID8
ZuXtmQJXTKa1Oe42/59RNB42CXVqn1/yn2NF6prRsb4YPXY47LpwPLdV939S77Rw
D/iA27CxHmIr2f37cN6qhqs0qkg5Gavg25xVWgnHBIOLMmSlKc5tlAj8v6s/cr1Y
5itlAaBOCoJ+5rmPwYcfGPy8H3F3kyBsVN44Au850/m69u9q/4W46yLFKWpS3ct1
UBTssTV4WRx3gGvHaaqnSB4IkvAia1bjIR3iJPdQu52KkmkuQJlKdMEq7IoOhh8L
fQMbyZdbtet0dqq7QSaUD29emTD++LN/ORThNY9b15IHRbcvbKmragvyDm1crdVi
9C7k0TmVTGEot1Rn2IfdoArsO/4AYHUedZUkFiAanT9Sts2zQqN043chz7e3Fao9
AFRmESZQBWXgrkwBVVDMUh4KjkFDqkAeA9NGvW4ew2TX0TcYYNe0sRXbtdo2jpN5
p0sCppM8F8EoiV38wOZxP2y24dTisKO/VeZSxSkFeCGzLjdBBCkx/YU+IGFOHnnP
TaZ56AwqO+DTOJ7xzJIyxzT5OPg3T8gTbQjnAzrUj6WkbtV0lTWx5j92bNO34A5t
DnSI0inYb67bSHn/+2ofxHRcMbYGfBJqa0A1wPnt0hSHKGmW0/rfjf/ZaYaQZuN1
MKrYOTR7ObTsd3HRlWkc45x6aItoZ5d7QL0guJ2VYJfEheKJBlgqFVS8MVgIFA0D
ScskHed8MfGb3dDKWA3B9AvNHTjWz2w+/ghfSpB3jPsSEHmiZRIx2PWq1onZAjwK
vy7bZqiKJSyTzKetu3JaXhWnJnEdlgvcXNG3YlnslqCzVG1oEeup7CbAzm5Fxdly
EXRqGIG1/qOVhNWeVkUCUydBZeq4OODDqBOWWk/hzMIo7QXIDSf1gLg2RWu3U0Yg
fYdJ2cNCuuYmohmUW2Pn5lf+dE+9CWIFGwABBg8Y6zhvKlfYFrn50d4WHirpI2bd
FJgR5n2HIuDk5fGhnz/tTkQD+VAMSybEBxry64LoVvLc9i790XmlFZnXrmZebLpm
onTr1xgCeWYIP/k5Oja1N9kH6YwAvPnskpt9yUl7KuNpY6VRR9X7v7O3NfogXjAM
ofEC0p56RbTeYTUyshmT8cv5GZ4DzWLeg8Y/o3FQVQv0dU2LmcOnKZ68EcUrlBMb
X4YUXlIPNUzC25GX+vtb/IDeRplecSaU4eeXkKL0wtMok5gHN18aUfTrnLLu73Et
QQv4GCsuTzzVe+LbFPFsAJyv3ko3z6pLbkSxalYqwKhfjkhNKM8u8Oh8pnwBuRPo
pcvMA/PzeztEjGaufa2uCMJK/DJMVwyJiG23NzN4PUhpu8obbrjAu9QPwFzhY84S
JOyfjGa4ltYQWTAun6sUlIuE7Xh7PBdnI7wVt+peDcCWSVtuDzLXuwq8VIi2P9Cy
bq7y/LZqL+ho1UgB9wA7vEyV4kq1WsDd4GSioiaNMuFfjeV5qijDef7eQwZoZF+Q
Oug38N0iVuDS+agJXM/WcWZ77oOUSVhY6LAeiIZjIAXsvQAgLVfywFY8VXa3XbZ0
tk8Hfjfk5pWlWW32EewYBRwIxvgAl1faeEdl/KA5w0fR9Xjy4LLQ+ujIH+X7JX1s
SJvQv6wfF4zhDtRgz5AV8MwjlZd17FqXTad4ZNgyDNTl2BBHhNetydCc0W/ccqMV
VP60vl0spmCjOYb353Gt2gEbfp7okqZeLv3zD1d0PV3R4xxHrAv0FqOBofxaJ/+G
tZCzQnTBN11QrqJqqXLed8ssigKiOycIylu62Tb6xsKEg2YV/WKtwndepkmyAZWj
/VEmk9rxTTgl1prVuPC/bnnWUu6T0NltD+n3G8QDlgcYqtwPlHrx3wMjFvwhD72t
uTwx1K/K6bTMcqMkH+JMc3WmJfdo1e5NnADRO2fewv+caqPUt+Yj/7lUuVsGX+uQ
7ugwzaBGt3HGAhO0dwx0T0YSDuwJe0f1GlhH3M82QqCc3jxJHo766u9thFVe9Ykx
rYA5/Cj3MvEnkWS79QZ45auOok0BZtq3GpBRO2VxnOgiYnJQxVgEkvwqJ4atN2PL
UZXUyekTCzDUBkbudFhNajzQsIGiPPTKy/VKWR9wR0hd6/X+deWnBOX0j+qFC8a9
EFry91CA9eWwv/Nq+Ql/9NO2i+VPheDrgaPLQ0jojhNp7KyI4sD9B+DKg8wGZ5g4
PE61zQfmCZdp3bhNTaFecZXO4Hfsi7mJGn6xh3V68hzRX1aM+KMF3EPVNEveqYQJ
oLSOihZiYhgRbt6u7cG+6rpH8UHSQaO5NGG0KjY1ckS39Du596CUMaHSY72eN9YT
xIPUWZsOP26ToOhZCTkGw1mgPEjB8AEMGGmEH8p1oEed55vqzuh2HqXo28F+jqLm
G/oLvhAY5FT0NeZ2rag1BdG7z4AWmg3H77jx8FLXnawfPKAs+wvJ0zccKpO0EWs5
fuhch5inZExXWWYSIYfFcE6DEeCHEJObAa7i2oCuy2yBSkzdZKvWjWQZkFCyzOt8
yI59dwM4EEqhHy4rU43IgvWcovmmaC8poEv1mJp1BAuVyRTpXGzkmoxbN1eR3r+p
VrbsIZvv/TdN45H/AyFK3iwBH1SAJrvN8kdZgqqpowauVtiUhoYKJ+8aquxN0WUd
3c1JrfRMxW9Ud6nfMbR3REsG2H48mh+Lh/77vhdG0q27ejxXCEbLkMGFsjs0/UuV
ngzCrXnx9YxDnBu2SwykDA9HtPUQ2lwr7ra5fJcWxdj4ZRucYlUJGBuZH1RFyech
K+SP8NW+ooz+sYyjXwUVEae+TwneI5Lz99gP1FNzlXrRdOtcg/YOSumvCJ2sAvsi
5FT6I6W4VA6LoM1qm8vyeBwI9N1JkKQdczL5IL+ozuGJd/GP8ZJiPg3MVZcLbbtW
J7eLbKsxhb9QjoSPt8rmRkGlaidhoDCL1OK4Xs5xEt49BBOMHW8hbhu6d94nDgRi
PZd29FuquLhMs6sCzXwE2JiRWIxAESaKCeXaRa27rdu06AeVkcbo1M7fo5hVaTSD
3bRnSANPpR345QoKOGPTDRJ7bkND4WCn1r+kSzHRhmEagllyygBWwqzz1TleCLZE
B3P8IFfN0AB+9LG4psLYOGlW72b1asX3ijEkquqWbnXUHARdllODJsE5fbOXKBux
5SxCw2vBPtS5mY2ddepG/FmwrDvjlEEUhim2TsU82BKTsZHUxxB23Bs761jkADR/
n7YV7eC1VKsxQhkpOU6sEusOaekINGU8PApcmhj0mpReIxTIHkLaqzUk2CX++Bzd
TTNwcFNg3Dr6hLHuU86Kpfnr/U1HLBJDLX/XNs9MptniY0GafQim6cUlcO7RDIz+
V/BMI+CUNVYXyxOvFZgyQmSR//X02wl5xZ4JyIqRxHz3G+x+xMqv3gvcoqzvDPxv
O/inCAGer89dnTYHKknjDkw/RfRLdd8Tv+w7Mp5EinegERzsltJvsBWIT6yoTbbs
Xw38SF5crfgtAAp/Oxhote4rnAgzxcWKi/rSGKtJI+WFB0gNFg4Cke6ejsJ0tjKm
paUeG2zO4OaM5ey70xdStZpg3m8JPUUoe9CwDloK5XJnxau9ZQoH6o5eFdpc49eU
6XBRVq15038uEBNmNg9Ia9ysbtbvVNyMXgV5fSVAa+DRS/Gk3I4kMj5g3wj7TE+f
Tzk01v1Dp68oWD2Ow65Wz/EklvKly+78ZeqVIkovvZ6c7FYY3Mm7cJA4ZVhv7nkQ
//wiOEdmsGcaXWDf8UWurcfqByo1r9OyRECMTTf0ZPSZuQ46KUIe71CDDRJtQODF
SQvBdL7cENpNABuE0qwnYXY3QKuRM+IlXN3DZRHXhNBr1r7O5zpx7f+5NPQ+TX3x
QWUUclKUpHvcRfi6juESjW8aAvYhtN4vjdbFfTDs7al7T2kLSe7jaONE6DL9N2rA
W+6m+O2iamGeLDmlJQVSZWWUzBdFT1YOKjsWNVP6KxJMmpH+OMad7E824dtxgtGw
wT4uCaUD4HpdxHbBWnOzvB8OsNS9PWnP21aUL/gy//escfvri04NpBCfSKOAT6hc
IMGN9BKpMNAqTdoKYdplmwiHvpniKDlfIOuMoAkJYTO4FpRIUj7zze1KPid+ZQHO
2uUZcxjLoACrXoaL0YPhng88/Fj5W34bpgZBA+ip7pnqdnOHQdaB7Rv0FoBvgWzc
CZWvaYgCpg5bpNJ/UbIWfPFcmGTwavU3gmxt1FqYql1ZOAImG5GSQxpJLcqYo0rW
bySOFPqfkl8l2lrNiSKFBi29BXiX4qxiIXyt4izn7vmExLX0ybL8eESLXg61WHn4
YbI5R/ydciv2cHZCBb23AESrsjhBuzVoCHHUdsYC4+khmzZU5z75j2DOjShe71q7
mPTfVhLhKTR0G/Ac1UuDBH56+4zqvw47m39FrvYQxFMSdEzGtEkbnt0LDu0PJv5G
pM6R+Ic7nZ3NF30oZPcbowj+i6ZNXrH8E9WriPH+eWPToLmkzoh9NkFc8kfXSipW
FItXFe1ggrSSZ6Hzw5XPXaS6YPF3rSASl8o6z+2qspX71t5SwSGcJbg/C5b8fPd1
k3cKkhYTxTKDLTvJIyEwfY/yQiWp9s5QAB3M+OukgJROOCZQy5L2eQHBrrP8frlx
+w+S3wQd/PgIpWcxcwMhLlPXOXBoxByGneOjXCm3daFvaV4vBjc04Q1BJxOz+zse
YR8Vo/IYb93OdXMPwxtHTIvFemzqhBzZph++LWGZsqDMUcBUItzG1L6na/vtRhr5
6ILksIBECOuXdH57jFiqwBt3QyhzB8cmV2A57BqWwzoQf1tfe80/n/B2bzKuchHh
CMzRbW1TfpoQZFRm28ntFtdabRR8DBuyKVTSi9cdDdOjYpO9iCCiQwWsC5vyRowb
hiCxV5B1u22oJmt9OmyzfnUGPvsR0YFQ2j65lrevMgOZRBQyJIZPULeTvf1rBEmT
Em7N5uNvce/XKXtaGimwQ+w7vtqHXUVd0U8vupqGZ0DCslDFkcCbK9GWTHTVxY8/
dJaV4ZDoBxBkw0KYRWU0YROC+CFOVlhxkMHDPL0fq3Onr6Pnl28NyPSq2aX4Zi7b
f+ZDuzpHJmJxduCyMIH2P+4YtSgfYCtNVSmktqvCEiImu0GZfOPCeO4UrrTAZmva
B92GmHjv6YnaHRFjcwg+ocUjHa79wfW4XcEmNu91PB+3TwrcOWMHbHAhAIIISTzq
B7rXhgxaVM50mMfOGVjf68WkJdiq7+fhXgRjsIyd84GyYY8jad+j0af5XKMpa1e1
T16Ze8HYL8hT3wHwzL813yyhm2xiGmFm9vReltwwRikswxYOeIgHfLYULIjnXXo5
6Jx2ulMok7WWvIkrtDC2QekuoUVY8+V6toxH7n9yPjbB5p3A9qIRLcR1A0Pxe7Vs
UpLSiptoz7yb8NGBPOCnJ/Cp0vmjyJtkdf793wbSqTxpzD9xRKfttH8Drh4H81xC
VzNxdFd7ocBcohSMGxtbz8BexS42AnaSQ4pksREkt1pMBKZS0OHFoYei8JPYwvsn
/VNnouvtJee2PjIIVab3/gyiaIB1ruhojYurQLYRPTrGIqXzmTcSr/cnnHhHgn2Z
uOKk5IyU91XbaJfz5iZOO5OG39WoHX+Ujue+Xquzc9wCsjMf3WNA3d7cjSV71fWh
jukECzrN2YEw2wglP4grk4PUI7L+F8VwboS523Xu8k7UA/agkd9eO/UZgzmljtnm
p/K4odMQFUS8s3RyNm7gCRuJ+M74BYu+tPK0U1IfXVsYT90mSIl816g3ohePztAv
eAY4BFfHkKiHarknyFPltlm0FbmgIHoF9nYsGSuNqthQtQJxT7Vc7GCCYo9HJJNR
RJqiaIERZ7+2OpXpw0gIpKQFF67NHKvBuLggKx7fWVG6V5y4gFWzjpnm1ql0BuL2
wNjmTp6dfdEaP8HO3+TEW7vNO8lXIkfwEC+kNUkifmYh2bCSVH7qS+EAdOpYFGU7
N89N4+2M1gZxP8idfD+GF/I770xBQ2zGn/qQiItiPQE27CMUVrLr5HSGFJiQw0rY
OD00bcULyq84XeDzVvtJAhxCdY+cJSa6nftH6StPo3ooAWDYDhQJDHCf62CatQUd
bPXtuIsS/sC/1DKAbFA8cerDtWNzSKa7pNxMQYV3xl3kv2EuBI5NkWoD2IdyMJH9
JGulrHw8AjhzAKP1Kb8vzhAowFT4Nk252w9Vxrzx8m95Y0Sdff19/c0rtsH+L08F
ME+7eiq+S8zTM+hia0ktX1aFCU8kwJ/d0BuoFVS3qymn3r/MY9KASH28/lxB7xTz
/oAbtBcZSDvaM2BtrWjj6mzUSDvMSEb8+SjH1bcDf38WO1ktKvoRc3S+rtWED1B/
S/4Pp1FOgWW+UAB7U8Rc1nsV0AhbOQu2ScJFrzQvLekTdRhDbckYxID80lX5tcN3
Q4kUFZDaR7NzhTAAVpYuVDQKioZA1xIQcXnk0sNX/11UlIYj0REtNNoHnvczFZEv
T4Q/JLOu2xwzGOxdmAehAM1xdOfTpcxJXh4UC2cV5xHeA/A22T8259Y3iIOfmoJF
6dPKOFBrCuwu/7M9W72Icr/Hz2o9ViBTr2K8PAE2xxg77fVx2WMDmjqldChrg6oI
PIqsOgsyuF709w96i61xGxTRk/D3wKWs95jeZU/PZCx462NYBm9HWbc3ykpZnHXg
sjUBhanPtfMaIXH8T7AM0OEAf87tuWlSx6uva4y6nbqDOEZdxtouMvZRh0+JYrUf
ya9qALmO69Mtb6px2D7B4o78WFo/Zb5sUdeFNDZTSFMQbkmZXuyfoUEoks1CyjMz
jouWQPsCapOdYzuHF/a2M18M7MyhijEDvi24h0iBuB45vtrFY2vnVae7nsZ++vUZ
4ZQIOMqzyWHNM3TXTPtzHUxu+cyqiSa8ryNz1CE8zxzggY2xC0TS0cZB6qdQCgnP
0DK+2Lcd7jDTfXuc+P6GIUJ0v/TL3eEcWpvlS1ut1LjQ4Xn0fwiyBCw2qbMhPt+j
cV7NTMzJb7FOAHCB9MlMh0nB3+BnFizbg8oHCPqzjbIuT+IqohruC2hBRhGxUYFg
DHTcSq42v2xDkyZOHk34+BDW6aILrHsMUBurywC5R3ThyZr9RLWFofIU4wZncuhh
YFusuTWVNym5lTjKGtHEct73bLVnS5/AFjIuPcyu7wr3msrwNKJozGynDdd2H6ya
eEV459GgNurcHTuRFAl4kqRUzfqDgztONwuWTvTMo0bsAcTXXNsLtCfBIDLrjsrH
LejYOfhJTCi488NYcq8e/MRhKuhOP/YWCNea1dsOQe2hrw/b2qHDg3soefDFQqnm
pHEQWtIgYcYb8zQcK88abQv5ZQdsmajBQS+lm0818opWNZWRHiibSmkH3OPSgxED
eBHb/hAAbg8y3pxzk229dcCf18nNOn1hJ/i57UHAXpmOy+5bz6PjgFUQagbSPeCZ
P4pRvwDI/i54XRyCvJTeOY+qc1YVbRHSalOD3kzDrVxzquOveuRcQb3Cov96oiKA
XCGg12J3/yug9wo3iF7A/7eobqEA83MJSlHj7sRYOLLzpAh1W07FMLydD9mUCIt4
rSRisIyYlVzNVMynxiUAhsXmHJwMMSOQRAcx7SNaz45ZCCkGtaePz4rbhmdKkN74
vYMZHDFNWz4jvtUNr7x5ki7IFUGGQvK1VIe7nSGdT/0It4JKuf/8Cl1V2qGZtj1m
vxoP3sKsPnbq4PafjZOhncb3jP+J5pqtCc6ThGMwHtQeVeMzApXjAbSRUDdKE4PL
Hx87Xa/dzDFYDxQs47amWt69BrinUdpIQ8th2MTuDjJakRPauZhwLa3glEoXNcfL
tXpnxD0ZvYyfI+1QJv92+I/XDyH1BnK44ifx10aJ75HZEskFcMF77+PFLSvNGJ+K
vV0F1Hrpeid7w4fyiQf5RJWtd0fxc6ndaTWHY9zw75lJCVR6b1NcrdCqS4csTtNG
ln28Y0LaaCg1GLkaRVdZDdI+km9DpBewx6Bs5qlqnImE3ulKXCzlzBl4tdidoHLC
D8P1IkhKAh0WHezP/x8AX9frUFv91RYJHI8KXTrNwt7w4SUMv/meKeJtdkoTcUyG
bTLtuidtciNIJaNHtYcrsme7cuphNmEBnnVVK7KWjYGlrvmj9QtNfDJR+PFTOASN
0jtSNnAIvFhfn4Fh/yNrjc6204cUZVo8dLaYbY6BJvQOtDiEqHFY03w6aHeQXE4X
sGvYvYFK2/R/FYJaTcEMeEVJ6WJIhDB1gx8UAx6orvCynThTHifYkqh3TFtvoI7d
Ys8iecgDSg5LVHKO2hLWXqcLVHIwgQrWt2YsSjfAf9KseNDXchcyISni1vOcI9N7
XbfTwL135K0qY4999Dx8NXfyviVcl5ipjU2Fnb4TqrZUaFx3VWrusYS15ql4sodY
2E/rb45dbo8zkL17+HlnTGmiQrhlsEYPVhKCZi40xxRXJza/MtvqCLUgDAvz9Rpo
3yl2sjWg103ylj2E237Pc7bTm93SQYyxl7ZbIyxZSueqL7LX7ssQT7LmW/vi+ekN
qoQauLsMmRGOshbocTfx9aJZZWC4WaDKhPeyiueyrfKG4XSkkbqfzqynZxm8Bznr
W0vVrtl2SM0GMlL/udlwS1M5e8EjH6lO1Aod1rrcGpVJHSFS+jKLLz8VnSog9nIl
GMr0zBMGTWaKq2L30G6g/eQqNB5H1kYZZmAeCiw1ZeS2zZIYM9YsUDa/9+fmxSgZ
YVswg1kfZn/BroSdy5sf/0ux1DWDucQ+rHozbtnyYrM0n89QpNvrxc5XmngmkYjO
ZodK1JHkAeqJMwzWqTD97XezLYA+ld3PH7lM9lYZ7fA9jWZP2NaBFn6VWoB0mMZg
EQ/Ywt1z6JRB4MlzSZZSgdpomDkHnY/ZptpYTOGddpHHVKdQ8Gsrt7o69i2iLzVy
iP8rJam3rJVdJSV5v134lch3clmAgVdJ1mRgL1GiYwKpmlaw6oOtAX65w4g6y/xL
eBxBarR2yHfhx5ylMR5+L6FPAmvd+V4u+3gbV9X+3uSe8WnuHfzW9Gv6tFNdOzSZ
6k0rH/PmHZeR6nJAemKQPthN9IyG8NLPCDVf88aTG2Y98pArKjHH/Uz51MqQ90Es
lH/SNqTnCe/u+2jK74Psv8JHDmgSGaHM3yYXhXgCUYuH4/ji6sCyNsnBeNa1Hk2q
l8ZfA1Zj/tL5cHrAGmkt5jsGcaAP3qJlo/BIJtRlYneQ3c5fXcyJMZoXzYZOE64P
Wa6XsLG/35GYdNYIp90JV7NjVOaZ05GoORlIdZ8b5tVa48COtV9tFILGFBGkGSr6
CukXxbxvwj8oeUcx86Rt6UbNtGCmA0of9fkdxCqqNE5rF3sNUfbXrB2BIFcTDecr
pTzKekEnsFMmplBuGkeMCjAoEVXrpH10j0GdU+gF1hkjrIIo9iAs/WswacI4NVPL
Grj+pSQkJlF9agupAYABDglycmAkEJyvH3ObSc92MN6IqGsdboZEfyQ0cS1JCub+
bxGeABTEpx8ULdW/TAjG+XPYWTqBh61DRzjuhe2neR5ziSnqukL0winRlNqE1zIr
dnEr3PeiD9d2/BOK5Qsp3ZBzP9ObaiuTjqHRGar+bbkOgyNtpmALcyp1poPo+9EM
C7BqKfFANt8UdsHwcWzBAKMSskTYYyeNye82c/0LPNfLsyKs7txusLGEqyquTzVb
LwQOK5AQDLcgniEwqrJu+slH9zP3cWtvHNmx6ph6hNHtaQGGRQ19wZ5MiK/Q0dND
pzAPw0DUtWRZRKB8iqxOe3PekrZyZ3gNECzVtEE/5OoBGgIbisiEsqX5us0CUIh2
AQPU+itQQNuKa7ZFPMEl2/d3bP3fbdk72gOngN/4f6LIg8nwdaz44KU6bSbpKna9
8PUOM40COzNRpy6cAt6jS0bIJR8OQnve5pjxlsCXpNtibDOR+puDfn0BNc2UAlhV
iSsttOvJ/qmAvsmqODTqlTucLUJZrKCpe6UKktLEo7IAmQwUBxQvxuS3ElpWHRwi
q2FKfgrZiKPqIRQ15yXSr3Wq45S7dWy0YgIH2NJfdfK/+QlfVr37Sr5+UQaW4hd7
9bBKGnuVQCEK2DOBWXI/PFxruINNQnfs5LAmalK7yQphFowE1PaR6FVgwrDBh4dX
sRzCh2zUbkUnRjq7E7dN10v3oh2mSpPKHtnuQ5VwtELu0P3Pcy9UbCsgzSywd9lD
vgV04+EOjcr8FMwSbQp4Fam4Nx9jtXZ+36TNxFBWGx8ob1hmcxa4kDVHKqZ8L+6V
7K6wnPFcthmtc3rXPd1B/tWXbMfUCRLrAK2aEJgTRn5Q1TTk1ncb3eqhXW6cn/Mx
S9CYBpP5wNUQquYKuMt2OB7cfJ0nVUf9rq6VXDwHXCobNEBlLIdKGdWRUffOQHVv
Gp6TwXP4cdrItnOXQ/aHsgaRl3rfe8AoxK9UFqoJgyLg7mWe+JjiLdByAhzrXpC4
aX2ogfyK++SP014aAR88exA8+B/Bd7IldD/R8TXeUm0kW++YB+PgGhb5/jRvMU5E
gP0hlVHxeT7LAtcppc0lObtG2YkEtVyMeYYLmS0H/zzTlOHh5Uxph9GHdgh32FDm
SEwiyBqvEQdcOBInp836rZAOKOEoHIi1lqgf1f730trs4JkvFUmnLwjPyGp6Ms3X
1ca0QccJdZKcEWHNeY0rHF6hNk8SBGS8gOI3zPBUsMMhszIpPJh96nj2CYlFfrHq
VMSQLvRGKXz3RfdmehPmSfFYOhIjYX54ziX+zKSjWOZMZYcWtWuU1HxBC15c/c65
FOCwAhuXX+5LRivJ88OZ2fPWCPSDZGX7KX4X0fAjYHHMRHzy/JWpAKG3/A26E82T
zFSDbxmKpfezva/tKBHduQdKpQTFnQpTaXKI/FZhnUOC3yM5u5m4bFu/+UqJCcp7
mdCY+ANukrjrmfaXZGDHiDA8l7CqKt9lYAbEMWYTZzJoZQwihq1w53i2p0FaQdcq
R5oQuBv6JhFzFS1fHKlcDMU1mo54nZzsbQHZNRN+BvTN4Z+X0yvqMRCSJ7LWCHFX
uVYKtWV+c7oKqXoKAHpds1fGDT7Ny3bbQn7p43eZtEp+Vfun8gDWU6yJSTJ0OKJl
pwJPvZu8Jf1vVbHitQE+gN2qhBM9kUVmY8ZgKrOg/ngZfgrx6NBnj801P/4FDXd6
86rpHOXNJPU+zhTSCNZxtpV1kcqBGhNU2kqWunUtIDbTmL8y4+GhTgQkX3RzJnGz
sC1z/kRlmSpHOQirgc98x/GYjhH+NSZVaB0xPiOYkH1W6BM8OVubGlx8CYgJAGL7
EAwTmG7ZTZ2fNjvFglDb9DWvSySTtrmRJYCEGDcWr9bZsCVrhn+gNZguwBCz8ykF
EY2n/00twM2ueMB9MM8BMzcGbBfoKcBz6qw2UkXwn2p9zdR1hk63Fni0yZEUoywM
trsje/h1fbTn09JpNlGCPE+tB26e1HiOtkaQ/u2xWA5uIM95Ah00otBgMVmo6TnU
Qlcqmlg8AZVW9+GxmPRsf82rAkDOM6J48fzSzGGEau6UdthtTEs4KytMXRbutqdz
Dh7kfj08zC826r0SVnXJrZeaH8Nje0R3zDsG1ahyQEHDo0vrVukjUUvpRYhIJR5X
hj8KNGw4q8MvpOy9Dbfgblh4F7XWqx1YjVxKIGTvlLccpup2vV6gOPc56SYLi/CW
hVEcZMfSWYzuqgid7gg722SzF9gffcpyTo+FX84xn6X9//XhX3/WDEnMlNW31pCV
5uIXwNocBUokko7HmyPOPqaV/9mWmapaZfak/skFQ4An5nGRAEBCFtQW3fxq8syr
c0sZTpoPMwsuKgILWN7jtBb5JVsNm745CsjvJhTse5wmZw3Q3+TUmCHLVGNs91qe
bRDzXIvxB6H+usG57A1iStjcpjSvSWQdnR0ORDEqnzywI3wxIksl2doLlps09h7l
wxKzY6EnVb3VNARo4ziBp1Ra8o1GaW6QKG7ABq1ODOhJykhotm01UNXrv6ZSrkkV
N9RueiCBwNIpabVCZLdxHRVnRjTGe7YwACXxfhjVzRPWIos/AN0SXkfVNXDL4RHG
8xvmFOWgQ5uamFsl9TGGQNKDzN8aEB6ENGyn2wVrkN1mCQObZLjiP7BC/FnkyBCs
T/tug+/3UyB7cnxudSJBqP+LQ9F4DzOu1j7jDyXLj1l4lTqOdXf8gaYB8oTBotwx
/rPEudGXHj9MvCrqaruyskaCU8YNCOt0jYWyuBxpflWgQnZI6w6VQ2CS3x/zmsKx
H+4zljAgbqDus/wLiC8KXu97kd/hxnaiqGvNe+PpAaAHuaw3jtZBB6Sw+DA+7tID
ylYVxEdkBIaJQ75AvDA3yR6Gyb9y6D1AokgVOVnYbBCwpzBcOwWigY2yVbGfaMXT
2K1KdSSbN/rLz3EMTMSLmszZ3J3Cq1BCBIonOFqvFyg91IMVkDFY5HP3UADe7CzY
4nSSYp+NVQcD71wsBetZkaIl0B7USOlHYThCu+BqyWC6FE3xUdQhHaoxGNlnIYes
9rRTI5Qb/okJDXR3GFK+wjvMldc8PveeS12hRIu+G/PcGdoQ/EMnjduSgwJ0ZBU2
QODKXGKnrQ/Z9PvUGE7P+I6CofsviuEJqu2eoub/D7idUgg/CCb5p7ebFaWjcWBa
sqmftD6Pyk21hRGIfnBpSKCPCJSO2lPBhTAm0I5NI/4tI5V7E8oU/+uJa7+jAnqB
irWnZWvJeR0XR/UEJLDV0wVyVO+sPA7zrB94Gl4ev/JRjUMFsvT5t8IZS3pfgg2I
uLI4SXjOymwE6u7kHbNcXaKaL5jnF9oxQ9cp35bKbweJCmgKWHwe+kwdvA43gHMP
+CxSCZuhUx23vyoZYl5RLNqyMk0e8PMdG++xTWP/rOB8++AED6wGAtn+Ar1JFTLf
RytkZIB00G4aBSjO+mZ6fstQJ/eLgvUx0XC1Ev395+YXjp9ZUYeqdqMmNYQexZmc
kRaDZG/znBcuhOe59Z7qOUTP+K4IfTiy8IyZP/qYPwDVadJgk/SHUe8IMLKASh9G
W09xdEFPUnFBYpK9wRdGqGPBuHID+8loqAI/9qXnCakaafywIsCqAtRY5k7zk8QI
VLQwo5HdCDKUusne1y2QL8rKY787ZssRd+wZMuVem2udPGVdrkWUAyI7tv7k3sfU
5dcyTIc+1PSUXQzK2eqheCarlsClc7pkZICd1mvFBBPnp23eXo4ky1I5Rq9dY/zu
sLwbmuaOxU8bS4GPhLnxWVs8HtuJ+IkfoonOsYW8WBo38RzzImtK9lyqAPfqi3SR
zvg3iH1DM0fU9RNvIsX2/i0XeMChe0k5Wb4eHSB6hLG3gAAirqby1sks23flaRPl
aFMehcGgqOormGaBnMDs4GD/cW6mNeLqe4oJ4e7B4zaFe5ZBvvdqqkQu3+H/llIL
XxwW+4edBbUOfJfLStlkKHj05kBcpL2b8Gv7w4NXt/T/LEpgnopfEps+l7sulqEB
qVYtP1oTbYzREEFS0T6tksVAlxmCvLkzn9d/8ssotd/yQCRoRlrFVvJswI2o1QA7
msOnLxigkbN3CooG+feP7NCuta0rpShlsdxPwZDZVqnT3doRG2EnwS+AFyAsOMnf
5r7gvyHIA+IEj4c37G03UHENu2oe2ymKyHQj8kFqbT/UTK5hHGXBKc87Qz4Ad8Df
ic/He7GnJOWc4dS+N/qKEapSlcFBUzoqwYLnoHB8/KFPlLlJSiCG8Yv00cwU5eF9
ViM/cyj7JVhNgeq2rkVepBmkX2Pgj1NGjufokPBzh0WUVLIjngdVDOjpPGtOfeuF
XVh90KjcacnKd0H6TxXC+vBoswuY7gmhHlGTW08YRMXVfqewsKkQC/1tUJ9Y0fAa
PgjsIZsAjLOFusWuyIRvQLprxd4NZFhV9eobDCTiHOjPdxdmQdGREpKKauhwwK2c
BKUqfxksZcY0Al5m4bEa3dn2OMnfUQ60xJQuP+nrci6dwsZn3pyJvml0nvjyv1l3
j3wlLhfdjHcvh7aF9i95QhyOyyTcZoL7T/MW1r4BXv8rym4tQo1Saqqoy6MBf2HH
q7DSOy1EegXWkS2FAk5SgHzN6z+QVbqOJGNsaYGP4EJSI2knFi+8fatX7GTBaIJ/
GgIUdGQyYXOfmrxjrcNvfF2mfdw4xSI8OSTwCc0GheEUWrGWeT7ernlI7Z+KUf9u
uuiWPOO6aEtT6BSzjoRs513BtQ28s7UhX5Jp+XZUeYKtFprAe68EEMdCL1bulcLm
OVnIhlTcE/wndLfHLjcbQUHYZoRwp0p2sUT/Il2NBXUCQDvLifZ+35b+1Sa8EYKp
RTr8sjljAvMCMSDZX/50rJoWn4KNoCacYYXhFviI8ffelgD5vO44Oj4YXyB0vY13
wdYWhKe9E1LL+UGlPzxWzD+cv/1/gCT3FHpYMp461JSqB04ZIJWuIMRk+elFR5I9
dJULIgxvJ3fRnubZO55gw+1OTiPgHbcU1gYlffHNjpS+KuDhokDDXFv+PrzQqqwv
IwuNBYUMynVttJn6Ue4rm6YbIGERYtEL44ulIonIxlDxK6MEJltXnypqQQBmsThl
sZjTVMz7ad0MQrA1I3KulXmleH7PczO+wtHQ+kVG7CUDvsfGzzO3eL8rBQzmWTtP
nx4A3fYjHLo5chi6umW1ppeAYfKBAYE3PqI2jClK7mjY7DZg3a02ZEfc+oj9+n50
hoSFZyCMPnFtKPV5txsnjZQdn/n5/2SScZAJaU9WEugoVTW7Ybib3bf41cRIw2gA
UxhyjGT3gWIv8WPnOSEjP4kRX7ojPSF/D1VFlXW9OQOAUkx0s4p1fCIocb7AD6Ew
n0m9UmaQk4OoGFI9IPLuaSbe8EM90Y3Cn4jqd2LJQvjaYiqgKcl2MkkTnUwW+6Xt
cWcXEVX4WdN7mPQDxM9Wb6oQ0qNtoLzAmV2K0N3NesSOiO0tk5fUPQaFforujFhw
Hw79pnxsCvUCakL9Hak9J+SfIHs5Rqg1urW0XqlrZ32ySXa22IwKHwWze0tMdZje
WnYmYjCx2u942U3jlMC0C9sl3iVsZ9DKxRT1ocLYiQ5XBO9mf/TtfJVTrTfWM8hB
SFo7pu5y0FdzwReKboEQE5LaqD/Fn5tg0uHIJC6uWLoUgk9FwBbZW/xSiIZCno3/
Kcw8E2+WJ4zmupsiqlua7yCuCjCr2BrZOvd8silQSKGgBwHe2YZr8TRrH87cc8oG
tkxJQfdf42xSnsFyxulvnoipYqM+cK5T+4KF9Abnjc11jCidyCR9imwMoutrlVw2
PrUMv5QP9S52SgCwMgUspyXOtmDGXpYoPoTzDjNwtlU1tp7eWwbZHWU5K2FOFlWp
AhULKxjJCE3hoVtcvtpHrhZ4S25H9IDG2D4YUAlVWXnvpcMOstIjR8C6puqN5+tC
O6Wof+tJARI1HXVJKJGWp2DIkTIfnT+hIE/nnXC4+In9cR97dMT7tSaAQNut70Ef
wtLYMHapQ9LZpbrGPZv0H4T4F1cu/gVTmbsZv6W9K2RP4FgH6zRFqyMNfJQ5fdgX
Joi1B7Q8l/hGBqYkXRZGjITzdyebQhig8kNbpj2OD4C0AOIKXHgAAOQeZpsQ/RLt
zvT0Hi9+Ci8exHVKd5NvqdY5rJPo2YdoVIPtMjvbX+QiPiFejijASmuWcuzZj0vs
q+01JB+k9ebnCNjAaevIqUAlNEWdr0f6YZA319CcjAyhPNAoik627OTCKsD0ilZt
qP0JXkKr43vNSEFGWVCD/fEyQ9Z5eXpAjh9MNCvJt/KRaruDAe7U8zJrAtWH0zhV
j8bLV5C3FspCSalerLY5+MZLslyZ1Emmj2lcZl/T/xjJRioiN301BaMEVTLkpPnm
6PXXODsRN5LDSt9zed2ipoUS6Bq7pniFVJBdJCRHlDVOQmMdJqx9bYmZ80iva9qo
xl0pWHzQYcw/HmsAjYshOx7gqOeTKXjBlmmN0hJQdP/NQK1AnwckMNWou6tsnzli
+uvhZFUP2crv4pgetPEbNy4EE7Vz94DPRCYAxhvdCjp07KvqJhNxNY40HLMGrOlQ
GaImKkCLGcgPD7YhzRbsfMh/MSkDUlsnds6WEoh5E1QXC4j/jvrFYUSCux+vZn7L
1fNVDjpX5C8cQ+tR8+6EysUTTvBVOgEsHx2d/9HJj0fJxRkTGBaI6WHqkRiMqGlA
TlmD3bFp7mFqNqnI0oE/NibAVAKLHt3GnOdR2kRLQ646rh3GBtJmj/UTY8VUyXcI
E34/25CzfYNkqyvPvT+KZfRR+qf35M1t6BB3g16U8D7FMXFvXj8FX4NC4IYsVlrM
//hgXDKebU1SAUG0k+0gvVVgaD6JYxFGKQxTmXtHjQk/6X7UKp8HW1pjGQzfy0OH
EDuklJ32yCPxDzHTd3HFmMrmqTQj3YKJ98+aMXBaJfkltXMB7//Ny7ztz3zrabBI
lncqOmfIMF2p5OGw1pXOpewXFtctiTquHUVs1lDc8mjNPoyuHrWYSO3gGiKV3qOR
vhpeAI9Rl6C5Nde5jzC8daagV6DO0esNpzgVFdkbOl54GoLrkBpIU5GrzIWuPu1o
iciFu4q7pbdnKG9NZsrqjRryTJSxTFIjoa8eftArgEZomb06c7iKGSLrbHfknB3e
+/AJbUEn/vAg/4Vkobh8dLNh2smMrui9qrDMnSIdMMWH7SCgJJDN2wM+gWKBX620
IgCHF3JP/o3Y0H+vgRU94mTKRpmaL4JiWJcclni9j6DcqOpz3vClvCVDj7cbxFfG
ATDJlIR/XYkgINuOaK9Ty5JbLg9pBBoctaUGjKqLwVyTkXcjj2kYGbDjsFqXaJV9
GxIUtv2kViKBugVwcy+ijpUqsG7WsIjW/Qa1cjhj+zbcEAIfyiMQdSCBEQE483Sl
VXn3RyHhuHgEN/LLoaFslmkNHE7L+TUXpcSWOcEuT5efDa1KTsuHlwhyEkamCSki
GTpNECGMhFQdpoGLqrWFamNRNgTmyPWaGs3a1krAtnq5zP9NyALp/SWwlEbjbgPB
N2U5XwU8PgeZ+NSjuIiiKZvSt9x1UBY6Aqf4VYibasnLC0HNYCUIM4OKINMfh+u4
lkWk5Xxasc+qt+Y6x6GqcznqF2CLxeHaW3THTdp70bnYNzGqqVYUKJtFw2nJNDSN
rAyJ9XVHE5jzBfDtpz/DXqvrM6VhnlRK1DIPqW5ltxioMrYlJQaqYpCVHM86s7sW
9Vvo1i9f82+c51vmHWVQO9ghy81+W1rTDxbaWq7YwXzTgr3oZoWAM6YzoSLfbxAg
jF02IozZIMs7TWSVW9L1N3jmwAHvvgAHxA5xYmn6CQmHOdAHqCUU04yhmVe+OugB
uCIKgW38M2hpaEAcccV6XXF4zVDJHcIVEpUuVbW+ZNE1JybxKBm7zHkOERkTducI
17QvwTImiOepxGpdmnzP/FG07kHQ/646IcCkQcNehR8HgVNX3ZFaAXXywlXOQtQR
EyuQRDxzACZEZTQL+6HT6ufuIFQKY/8x0ySKBkTDKNNPpoi7lrp11uZ43zskLTSH
a9LdFMADtqyCGfufNCGRtCoQTz6New1Kt7y2uNgvxRqYryILxxWWTX1fpRg1GEOY
DqDSRbicF7S00d33w+tIGRwDcGcrgWttCbH8lEp5kd112EZiJjTaCrPhrCmV9ugT
+lh08ceOGQqIXaxeQY26oYkgBF9f6oKJr7jLeq8XWND+UfZvUvUFDg3GJcER6dbx
JYIdrrdCYwvLuALSMy5nPyKvZ/OY3Qcvaq/aYVQ0b3Voch726v1hYqjUoOb8zKyV
6KkOfsbUzuXCaPw9ncCuVlyGC+SHBsqtMqpVJy8XM4L96phcZx2ZqFq7OHrq+zxM
XMoz+DnelrUScx8SDFRgqdf+hcpnQKmtdmnP+wcxMIq8bSb+m/SziO3Ty1jtzIb9
E9MagXAy/sgvFlTeOJdPbCcz18F9uqXCP99F0TnGhI6ZHZr9llqoCLwqYob07Vtc
OCZGkO80bKxZ6YbAj1AKSPomjAKt5Bo4jJDd5Yc2EStBXmNAr7Z/Splcxeme5lJc
A4XxXZLSOMbFdonKNcVvUyRxkuaY0r/TE70rtJ3jQM5s36/b37OGmK4qr3Uy95Xg
zlr5GUYBXwHdHruDa+/DHtouATHSxrjGyCLwVkuujptsJG68/xbdfo7mlFEa+/ZU
GUSyBhf9oK4BCdXHfwV7gV416gCE5kijOvWfBJ8npBiYjE8Ypc/rFOUFo4pon86b
21dP8mmQFKRsdXqh8zqu7k9m+qHGCQrkvUN3rny6T8D/9t7o+rJzLJGgdQRhE8WY
rzLU1lSrp+GpqBvTEbzvak1dGMRsATr1cWC5R0dv5qbbwCD3x06gvmUcrBpXSRvU
/F1WfTbpHVpoOApaRU+M/hHSeaKFa+hD9aDi8VJa3EI19I3b2WAqUUy5rB4OnxTj
ayAD1QYZfnkRGBwAjc2badLURFC/8/aTrZeCmzBtSOCGc2vrd7/iDRzfcIwMzQRI
02/pLp0BI2X/nJC7gl5y9oWi7sAq2Uqa7c/bIhDfuCavsbW8Cpu5kFsnfPI0Qk1p
cSQR6UCrLbvOI/KITYZ2NShzJjqTsTmrqwddcfHtpMO/C6vgsmrQpOEHwmH1KK1/
cVzSzQTbAHEF0rWHCpgT306cmD9ldZOMFnPR2Fo3gxuEafq/seh6CchRAAHM1Loh
ozhAEKk7Yd9bNXEnJDe53hgDe+3cHhAmLGz8k2qjs4B7TEAUduJSnktGYz9H9R+K
92y7lX/h4/w54Vkg78Z6KsYPVOFk3lhJHEiUAFDGAcXX30BnZ+eKq4vHDA1nltqI
yi1xNuzXYhObK5ZjEX3aUa20dsTVTld8DgrQmQd3XSqFzTrcKvfc/mGbPyJwoDfr
RcEhXCG4jm6TmHe8kaoY5rwjlMlpdzW54fSBUOA/+D2oxzXOev+3Z2EnrIDOY/X9
mUw39Pptknav+3DK4MtlSlJyL57sYOtt9dEAzAl3gglg6I/RZykdeZuM7StnjuYs
evTR0K7/AjEsp/eliUi1IaAz1efUpc3jZHOyZhXrq82uAGmg2Q1pK5LH8Z8uoSK0
7BINZZ75FjzztfnNN7HJan+/XSq08MvFlNED+BXYgwrXSW4+84K74CzONAHG/E34
DvfOUFRyWb8evsJtrlprRXD8YUeWbWaW1uSmlAfk0n+ZIojE7JVlWUqCQRkML1b4
fxUooh/U+BoSGUXaQqLERYimpDERkMEy7txKkRtAQkfQLz/l/43NJEJ/8xarajHY
V2BGVfTRmWRUH31tKv6fLdxd5Kwy8mYB/d0a4ggS9fIAXI+ZjCVakS5IiPxfgSzG
vBjWKjGKUg+BO2C4Ht/QopmuY+cW7elqSDWa+lC2Y6BrqFsAG6tJtd6W7AM1Z1Jc
jju1OUZ4ewHpUvZeWduMlmLlLD+682H4nZo91olh5rtSPKbQbCP652734oMnfjDd
/fbXNv0UUgL9azFjQY2jzSeqAzl52us6jT86+e0GQsFdJMGgxEod5AYO9oEUWGYP
X2ASKs4730dWhFGyI2F+Uovv3020nPILBD77Z/QOB32ziCNSsSq1DOovPrOl9zOH
SsOOgfL0d54MZpLRAZxQlhowmMD4ripUv/A6pQCyuWwdYH8V1SH/ZMhm7frzcL6M
vYTQaJLZqqnJWXl7Hfuah3CRkWidsWSrTv3OZbktPr2zLLS31QwLjxGuO7EH6/Cu
mNMQAuGA3guYJaXZznhO3yNxwqy+k/2P5sVlgjhxSKELUt7MPnqTk23gt7x5RmQV
dqsywPlTYJr4NEzzF3ukzj52t77cVm/NshSR62GpDHW+IKoCzjPRBXf6tdeVAI02
RtCcpIiS4zXQhxEFb9AIRFpqeSqB+GGx+Ako3GVVjDvH1wcuTOuF/Rc2B1BVRM8y
jY363YmC3wLM62GKQKaMngAbuFaIBBDOQuXPpD3VZGsqnPXonUUZAPR7SZh0GfXG
PiX63zyNSYSK1PuCvq5RJcvXxkb9ZD7FRrCRC9fMDf8eHHhcMRCNECWDWTYh6/Xm
1uHjuuMYisNBiiVhvGGAVTyKRsP1xeY+Rjk4nQ7feslSYkEVjkyMJVjTjejM6hvE
lsZSr7VXdT5yZ6W25oI5yIFkmvMEL3VxhYPIT03dY9e2e5jlfIAisnla2eCpAKWM
EPrhKh724wZmisUdGe/a0Aw03j9JyZD8c8D2yo5eC2xIzgeAMJkL7DNTCIhTnS9N
Vh5AzJpYWVBlvYIDAxehZHdGKgtLNDhEtXIk/SqoiucZCgA50JJKCsnSkmt0aaqs
/2zuuD8hxhHGy6b6jC9vMxrW6l7KGWvISbuFoLixO/ff+DOF/2tLLG8DfzHi5dCe
3IlretmcMkcMtwjiEVA6/VT3mD6GFSZsRYzbLdaQYuqLICQywawS5h1oACFE6YJC
fvFyMOhPGHSO4YHcNT8IVn4RsnL4LRfGR4XKrudLO9Xzvd0JLa3qx9pjgtF/i+Z0
0YzmUvxzQunHujF7VXsnt1rPI4qH4u7iNKpa2qwzIJtga6iCbSo6jsx0Em9S8lZk
3WcF28wU3pSgO3pa1E5IfKwA0X0vYp3XPewDKwg2BdXpNcKMjefRDQUBA7PFIIMI
HjYDsaIwFDnXqFUxs3rBIgndX+jetm7+FFn2Yaoyj6wXJW7btMkLs9QuPo7FEHX8
LHpfuPhMwjgmWUWOETfuM6+v9j6P4G3/A01xNB2S6Pd6TwRACBqJjQcrpD3mvPbB
BG5HhTWzzEi6pbn8/vwqeT2w9RfyuGUkdhj+qDKw9fswndq6yKe0m/aGkb9ENA8t
EL54VFnC+ulPH7DqSchYhVPJaFzKU9DNCzH5lIlZksDiwv1t6bDvyeVwyjkdvg9L
gKQGb2bk25F38DsTTLIhe7Gf+ahwxuZxccllHV0hc64O/avO48z8PvWg5YnildrG
b4E3t8+xJTD6geuinwKCp7j9Lzx2q9CWMUs9CQgrbrBxbwBb1FmYtI78ZjJxBnnz
nBnTvJJYDtg1gvutRou7yTALHgvzJBkMHwysk8XBenD32s+z+O0qaPechh+QwD4J
KjaZ5bsYlRg0zENetWGiTA+viQEmQK7sC83ttoQO4yhR8J5tg13OanoNooEmbouY
QfoxEC0tE0IyIE6HIgbYIlGG/iHMVVujPbT9mNFeQsSFlHMH0y1yUifaF6DG3NvM
AQTRFhHlKFvxz+VuEWnrmpGZwwFOCL/dFtj4fk32Y7pFwi6Ldb0Ui1/iuQRQ/p73
LgFHzU31L165jYujB4WtkiZkmmvCPd8Wmnv8fwU9id+m3Q67OOJCke9e75FWejXK
pJ9cqOiehe7eIifzAXVFpP5Mgu8cPb7rJkjK9H2mR+nSg/KfgmhsTLo9aUWbQtxx
FL6Xt2WuITkJrxN7Ks0QA5sPmB8dtWXedrofLVxaxmz0+MDM+b65E2DWeMkut9I9
Db9I/2hJR+aFmfHjYN01J35KhnxWIJEVXuBH9Qg8BRgs3Z7uRSUF4WsgPt/X5f2V
FLvuigUtGh9fU0sTL4HomhZfkEf9no/4Vw5AELzvVgJ8bEt/pr3iQXOKwAY4R38/
kxy831I4BUxmrroud1JhcNbJDR/z9IbckzsWsHgqmYXE/zD4WbokD8RRdq2HI1en
kTtp2vamzdb8VocFTcRS1kl+VuqeQp04OQG6jXzc5OKMjKbnbGXM+eJazr/vtGnN
QKy42rEksVUweyxuX5vpNkyzzbz81NYsYJDRJiANLvTMID+AXw13TedaZwajZ2/v
FExEWX1enJhtaoudDb/KWUv0MaminoLoUwinbdewBi9K1NMiArGAWcFdzzWOZV8A
9WCVJJhquTq09DavPAczBWV5BbBY2MnHT4xeNbzqHXfXTe+gk/HeU3vess8QC3qu
k9S+PIBVRyfDz7YrlTkDHOc/O5ILiVZiite6lrMT0SE3b5vUWbkqe2aNy3bW+NX3
TmX8UVBCohy8vaICgMn5z4p4MyHWPaICP+MTkZupQxusZJCKwHVqgQAl5/txk1nF
6suU70EHLCi0IFbauRiEKdQDAof4ymBZtRll2hVbOi5oM5iApURLZJZG46j6dQ8a
1Ip5ehhNYloCPhNBgowLCnUc8XfOc3cWTITDp2D5lTjNjcehoYRQTyU35iTnQpKZ
jP2kgYzo+XSuRUFYjfWQm30X5cjG3oCjORlqcIwXJ/nhgZaAKk2QM5TEQR0K5R39
jK/v0YaXNYnp217ps/A/FWjsxzPwWp1Pj8mO/BROzM7nnlethuj7zWEqb5euSxDl
h40ZwRTWV91fG5aIXNLgewz0HP55XnTOV/gpMekYDeNtkOKbdB99iyMu5nvZIkxg
agF6YXjkHrBPk6FZ2qdLvClPc71JnPrOU1Njlu0QRO2oM9+IqdKcRZ7mD38Nde+o
Dy3C8VJJV6KGjpjf2klbOm3IKjIXSoq2ivhUQ7vfaa9sScUIygrsX8khrmYGbfSA
fqdmvkSA00372kWzmbC2Vh6uYn5ofddblq4FwEflIpCeuhC77/StQJbwbi1kAuxz
0nQP0FoWfXH4UL2b5swlBheR4XEGHA6hmc/lEAJA5g7NT/VJqbq2wj9Cy4/8f1rK
FH6UyQI4YyyeKKvmneJ7deJhXRoM04IyQ9cbE7e3dxGDu5MB/lXj5JDM1bpp3LeR
Wgk7L7irBapbyYZhSVmTwlGdP+Gm8kSjXR8PBPZ0xzMH+mRRxKy18KW+QG0R6lBO
kfvVtwyJ9RK/5puxVeZJH8m2vkEZMP64jv7yA5Dk4d4XeVQkjgB2hohxq4YvtcJh
XMsM2nq08J4M0DP8SnXM0KIKWethWy3OYIaIbPP4xJ+iRXIk0M1ur4OFJi/ILizI
u5xP4la3ts3Xp9vCD3g+hxoav1KmKpOXM8Tj3Ha85ajDwpyhW1bTD7Ne6+AaHTHC
SwNG7tVfbpjzqanSGNrEyJvGHOx5JYPV1DFGkJezuVZSxOaDPJrl3tOvU83z6Swn
1AkNCi4yKcww7K3h663NqNcTD3P37wr+iH7yPlPB9KgzpEZOVA4geMzJ9xfiaWmv
n8nUhibSBLX8u7/HvjvqckUEPIkgjPV5g6zTgxda/X0p3vObecapgEFpxKGHbqbe
bqvBqJxbUYm3FKDtDSCLADzWhyPhGZIoxrGPlysO6cUmFOJ99EsKSeB5TkPAl0y9
WKJo+CI9jMQbu5up/H8ED+bjucYuFSfQ6H95olRXf6fHzB7Lh8ZXBgqovPLWV0JO
QnFpI9inkv8b9vrXNS/snOfozMqk2l6cAxeQTOhnQRRqqngCz2y9CeEqvBfaTjHk
MLpBBmjCBIvPZR9tlpdIzH5xYjWIhONhoE/SeXi1YGl6HWA3NW2WHp733bkqNQMf
DglVbv5vqbv0jRiLfrayWNlJEGFf9LZmyeJuXD206gig4H+2/pnLT3q00Ee/WpGE
vOH1tbnM84dmrb+Mp7fCd09A+xhMUMBQshKLp3HDI0FMagWm6VXSIjqkErzULPLt
DdJqXylSUx1kQm4dLpgFbjnjqIVpWXhW3VB2Y/0MVOkPNQjCj9TNZnFgnxfP8WQs
UdFx8fvKMEJjyq6kK2dHAUihEV1Hb7wwW2lUTWpDyNS8GebEjfV83X5BiupcUbIr
8KsZWI7rjn9YvhEyytjujpHiZ7YNSVtLYh6dmTAs7pVN6nS1JvaCjK1N4KT5p6Mf
J62+kwiagOR0HDInd66EQ9JCmX0BzL4/Cb/1UMirwAKjKXQ75O8a+S53VoWYdynw
IR4IJuCbkIbjXpMuqCtOpHe01E7Ulps82q6uBecZBMv6P8gx0MnCru9VXGDbIhcc
iFuR3SMocrBFsGAB07HBMuO4EfnxxsUw4TnvqTC94W80xiR4wa9yqJVPxAfzwUpe
K+qnQbbW8DIzNyLtVTU7exOxhhYlfyRcy2yY0jF0kgUjZeW6LaaTC5a8cYaLT7we
UKMy9TERpnOPLesiZOTB3Etn5Zh4Xpg3FdnK+/Q2cKlpvFCLwDIoMh+V/FmYR4gd
oLn6M0bHJqMiz6bqZ6S85LHltXWOatVWiUiX6FPXLuqX0yp+AiIzHbvdF9tA5zsO
3LcjEBmfhUVUxypyl3p76HlJfeZf5UOVLqHbxmoiJo4iTpiyT5xPpvumAH9knVKK
rf866UUK20n8ICzhOFgfxvcrtWBz/lIRQOtgtIebHFJpS1+2BcOzFLUGcMEiHfJH
1ZICPzvs0ZXl4gWIHxex2rTdJDcmOj1GiQ5qFS3l+cMrdHoo+NBS7/KdvJ5zn5d+
kmNiRPF1e7+yCpFcQZI/ppsHWjQoO5F8keazYuu7+UWKZjoxvqHuLRDXm/YbGJIp
qMj0ipnjiqbTPoHIxJPngdh+uPykrH+PXo5i1LCWe8R6Pcg1y8ar+m8xAGuATlp3
bQbJeq8OMtxnRqyk/E0iNzuZddFg4Z2lE0+JJXr4tzSYu73SEmxTIYV9yw88KMe2
YAHol/9CaMmmjLHOn2GpXVWPVxrGiWN4tn2FsYk/eUNkYaR2JoiBS1otf9NtVquV
qBxRQ3bJfbLsWLIr0UrvadJkdQd2aIFAXToxoMrK0xGtLEYmPfoIGOCwKPUYTbxe
zHLZxkluZ9CKRX6CKrL0xUx3qSRXh5X6HTTWXqTYjjY8BvDtCPbl05fiuiOSduij
38G6IDI9EQfQfa5kjYfruF8xJBQbXdC11ls+Fe9w0ihafAo8QXidNXTISMgXe/jJ
H8LTRTDyhoc1l021yKgqm8NUrMhszSKPxRq3kBbLBjFRw13Wzol+Kw9ovgYuQ7fG
10jiebkTTodmIdLh65Z5iNq7ZfEG58gKdfmQK0hTtwJC27Oc/JjoAlRBXT+cjHu/
usojOsJhqfnRCrDR/984ODqzi1A3uH18LK2ZbMh0cbwU2epJ1qOJNjTR98tyySNJ
zEB6wGjtoVz3Tud8Dq2u+vwfvTEM/WEeTyInPj7qyqQiJzh9Kuw/ErX4QMcjoiWv
40zq1D+jdHHgBcRxikweVzdFycVtlxv1fX7BF9dbyF+rzJJNAV/pkY7NhcvYFjub
Ci4TRAIflg+khRJgVXCBLEgapOEzpz4JJqZIP7NWaLDvrs9R2eyg1e5w0/SVkMfs
5fwJGOH9WsJ6wTyV4lfLB+feRwtB/Y+3SpLohS57OyeG9rc50F77Inx5J0CrUiXI
MzQs5TQegc3oxunp43ttfGHiK1Qs2ULgyHzhYDHAzDw1tov90NgIcK6gagG772cI
h8sa/RSim9mVz+DS5tWeD2pJsIZ5bNA7AzL7O6FsvfHr591xtxP9kARgPgKtH1Zo
0DAXYwuWM24wuSbj7wkP7SL1kv/e0GfU3WNZ2XSDtaGD4jYo5nfdT5sZscglr2k3
Vu+DHTy31L5fWuOxGWPxkOBJJm6V2XiO43w8TzaJMV4+4fpucfSeZEo+JeDiTlzw
ve3VFt2385VnY+DSo/GQXBi/Wmf8TwjAS2zAaZOmpcK3JfcpuARa8PLMfpTEv61b
C2aDZp05MX+vOT/whzeijjitTZAIwwVuI1JH0utdgrpE9Cb0/rN7GfTQeV+175j9
wvRsgPwVyrqbdombwbam9zZJSSlTAmkQpIC7bCR6GtsITT+eZlIzKWt4F0JXQdlN
iH1VscyGl09HYWZkSNK37zY9Zgu7gmNRRDsdBPHZyxC4wQ/m6L2iw/X78kDF2Aon
rrLwj+HtsDQllzxUCnlb9zwbLjDlwLI0th0MTxrsf/vKapgp49qoX8bNeQuuwJlv
hKNtEWpet4BO3nAvlq8VXTK0zaB37+QYLImSpmTqkUIHSyx+LSIcv+I78wEa6HgO
rWXKPzPz/KmMX9S3vACuP7AEhylTfyggL5tV5wpL4BhaAMteCbxnwDsdgMfR9pye
JbnnfK0khO4NM4MX8PYuFg1yPP8IkxRs4zDjMvP2df6jZuZLvwuJsBJcM6NtF9T1
/ixDd8cLBg87RP9zf5/bjPMnc8+7O2UOANcijMMC+nLe/43xF+iO+bRfd4anGN0s
gwNOEDoyGUw3KeVIuUrcKDGioP4tVzBFj2qAJGx738EsQb77iIN99Sw/NSSXSBZf
apHW4LlVjViLgDvx3GLbv5hyU/0a6JZ/EUgdH2ZubMnT6zXE5nUAC2Tk11jYSqBN
0HuxRtRsVOkZgcQONr+D8UYSC3EPQIDs6b3LkR7b/go0MzzU1ThMkzujcftv8KB9
DcQTL7UoUUsbLexXDhiDNior0KbP++YhFlcv98fFKUTmA9yYKG8Jajj0EDE+9Z3W
FzWCzKuexmMzD2/LakaOSVxknegQZtDn7HV0j//moDRBFgSC/Lr9OlR+j06W+BZo
gvHW9e4HcngBO1mT0xNTGIhfwivg4ecoiSIKm9zTU0rVoBx5mNAIR7F23iExXpLy
rbrdw0RBK8SaHx3ErgsTwG55CbE2qSMisvqLESJukE3yKgIgtL3zeiKT5Ar3R/b2
Kc1KLdi0lAeSTDfqR0HIa1DkI2NoxFmwYvAJHaoNlsJEV5NinTFeSpiT9bFxkTf9
IFTiOrd2w02pH1Prd4exj+n9qm9RLcgOMkMv4lK0WXOwvhAK6jkjlXBzb7XIedzc
23XEm9soFaG+L6YStZJNAl1ia5ALfwiE2IDPGkpemcEgexiM+a4NEn4aIUfNMc/f
kePdVo3rGYVQqvL1q/ysn8ARm9VMGNDUWan0GUiFpY5PTSAclz3Y+xRZDQFUcwXi
8dOWvFwLmWx1Gms+sH4yFiRZVX0P8dOTkOEKKyPir9be+1k8QqSfl4IFlWaC1yd3
Uz7DqZxiROX3F5ITtqb1V1b7WuBDhGgol7JKvlC8TjozJzKURPBuNRFlLmWT4Kjt
G9266+NDftMMGSpdJ1+ot0deQ+xbNAm7MkvveNwpojsiF5S3n77MMTlujkwQKWa6
S+cnawXqQIoqB2RdRgIXARIiPG5ryC/uJKN7IV36OJ85pejuaBta21tOakfL7I3i
2UdNF9UA8JCh9pRUNBgXLQAp4UQosFgSN/gwEvYMf40gTxF+6LxZaEFHLr5WYoO8
uHpo2jj/KjeDtl+scr6XsdJquwfvRt/CIKJsoAyAa6q/Qvq9+TLoxqG4t8LpfzeJ
WDJqC5o8AFHlH2l9xHN6BpC2HQmt8HEbuF8nTXmWkaL2Ecb2mtK3krxgJryJXhEo
XOm+s17gYdTarmYEyDZM3KdHw33TiOuuu1FYrpmr5H1HZ0HL/9+zoKA6eVXTtvHP
nmHNWAAbO8gm2n9Bks9MhgoUFF3w+ibPCC7aTWmepTC12DJo1NlCWZAJZ8hJT03P
ijj/PdC751ahU8Njini+pgnU+B2jHYIcc79rVwjkY5/CRawWVDw74Ai9NAPdg4Ph
+UwTAWVNfRcok6uxlX2Z4kpS6WB/RkH8VgnLqmpgrdNmw86hlXyFL8VsIABf91Ux
PN5jA448zojsNuY9GYcARkIQT1TulN8Ak716T2WQYiwCgbpbQr3pK4Xjw2DKE2Vm
ZHu3v/akHXrCFEIMDDnxTdnVAnZtT+/NRSNINA/+6TTYEk6iBUFpuN+5/xgMs01T
tvlk8CEZRpfH0eN5v1vUBbCVPrhLSP6pp9p8LXCVM+8JOA3iR45CKCu+Px1WByzI
hwaECY1MsapFEGUMg/NysWDffMqVTwJZ6F1nmj3M4C4ybCpwLGKxzgYtl613qKF4
qXYr56MQ4tYRvD7A0XEO96nyYHG8fMgSfpd1KDCpMHJV9b72k7tifBeqJRU2uu+/
YV1ip6O2PqhaFIaIDsQheD6b4zsOPEW0is9mWLscrN6QWOSqdxSx8pLmvbl/oHjO
XByqT3kKPWT+2H0QMDv9b+UpI4O0k1ZskHYj+HCV/goADNkfUDmp6PaHEJYx2g9s
dUhHgxrr2lT7NHVouRw2Mzq9jA7Mm7mGCzHVzavNBYOczovUkRKxVfijoTb2xztL
hQWp/GBsBy9G1iutDHoT+LUO8sw0JPa2eX/NEnZr84tBLDm8szrvtY3QWV9Pqw7X
8lEHnn2IksmbTyH8eCqD52oecZEIFbzJEmwDNy1xHma9iFGfbx7fbcB8Pz5BfE3k
fM+WvOsHgIokEyTsnkqPe98KAKq+p8DsQ1GK9GA92w/y0fC3vf0udENQ9TtqB9/R
/W6rdZWNGrlY13vRLTjcChJ0I9LEAZT7oXDclmyiBVnObHdnoCvBgF8ZL7bs+7gM
cLp5pzPx0ihRMrkVmPEKCbWs5w6Sl96uDSX6Mq++JNYUorGKcv5ZgIJyT7QBIQlk
DI6MUDn7H4w9Nrm9r7Pj1igViz+R2vHmbIH3JzhyyQ71Ksuc5XTkA4JXY0vuUBDR
8O6ehowTL6BYdT9vvo0Dtk5m+3AkvnegjjhE7xs4vLwpPecZKtU0tSM6qMntYbEF
fXtJvhIFKG5u3RBVgrwVESruEziRHnQPfazZNCvW4xMe6/+t8mH61LweLvzFX2mL
acZ3TPGSR8vIawhpMSAs2haH7cLTX1QnIg800F8l0QuOuG/3OrmAiw4U41naaVeP
vvZorshrwYPaOEs1ChH3OEXNGqulGejBCfWm+uWrJkh5HkV//JUx10YPovjgBQJ6
OHrGbgHqXbaTi+oNqOTrQPqTepTxgiqZRjjPTMi27AWW3gBCU+5iBYhhfsGajr5n
93t4J3xr+lFHbZjf3wypbpCLLg5HQUKAxghhE0pFrJF9i6F8PjYln1GLN2hIA1vL
GFZtaY8PopKVLI1dVqrpFtsro3RX817Nrvy8BdGjHCqnvJcyURq50EhjWywmF2KP
p7/qmSc6VxgnFqPeeQaxR2Wy9u35fiQdhCi2zRm2i3eN1jWMoxxdnH6U8Lbd6teT
qXt4kz2oY88suApNwNuTxrQy1FMD+hEktrcTKqkNVC0Zt6RptxvP44Ine63BRss+
f4sssSYIRE2344r71nxzCNl9HDsSufxVLVh3itvPMGo9tYTdV+biGFsGmGoMn078
AcCU46tQQnGmtGSutdMK16jX6Pa4XOT8Y6O2cl06qTwrBqbL+5x1aSpITI5o+2uO
DP7qax8m6CMizDDKwi3s/e/rEUTpI7MnzlC+Bba0isSZ61Yah6lr+Y898XXHzo2/
o1neoPWL2qCUbxTxPxmNTeUvtItWzc5yPSuifRhyfItSgeuF0WMm5avDK8ATquDc
1Cpd0icjvDBV+ygMZiEHT+wgvvj4kqRpKLKxchLarQa/LNxDwnrAcvKKESFhxE01
VJeMJnZaI+Ztns0hld40/S6l8cp5ZyOvQXoOnleF86z8vq5iPv2Jbu4bb4rcGNGb
4GPCyvuUSkfzXCuu9Rcx8M6DdZXD47UtM00WqO+o2UbgtqPPa7itfCMG57lRQnyD
zKab9ZTnlqoE2dljzQ/Gvfq4gA9syl4SYgG7Q4HVnQVQ7uEdWofdCWzd1Vf8uZmX
8Nu5o/cDqv42BbGgwSEtgoK6TPmif7l73v3r9IAF8j/OmBFXP5O/pFKWNQXAO2nn
yiKs0mQ7K6gq68dkivfHtcfPOjl4ZVCwQzifdo7qCpdoFiciQiEBZqGKyDfnKnm6
UREI4Du3+ALyZhQMkpJnndhInnM3VCanRCEgOzl3fZ97NMwSkkahjuexi1u+JBEP
ZqYBAZwU0861bpWOLDJNvKjHgRaSTU0x+89EgUO04zzWwbwgtcL5tdV8ZfspjXDd
DLA+Jf9+1job/uG2oin738+3LJFVj5+rr1Y2lnGVOyTT6bfcf9b4SG4sEEDiuZEx
X0EIHAJ4dlm55e7+aTtspNSjfDJYriqTvu2vBFqL8pkwGhFVsvnpkrGwvJDGgPxH
LukolBE8GSMydRNQ+b9rjBh7DMmCcO2Fr9fRp6frfR5HFwDpEsE6kjmz47qT8uxf
IaPAeyzo8znSOdEN0pKzudMWf84XfSg2abSbeu9JA454VehGe1PuGNunD147zhnw
Z5ZjkojxWJM66cF2W5ifoMXCOGHRNF/mfvCmX7RZ9MJw5jIBNgtpwFJXr1iO53Cr
o8hYFZm/CogrHEaahhT/495N6L2BGgN8kc0lASOG2tTScOqZpwkGTFgypZ63Eg71
HsPp5OszPcEq/ZYlDqDkxAu7pvTN888s/Q0D+qQ/KJe3Zx3uOd8+hSYJ7QRbNfy9
gcPEYmdOQJzyjeW6vFoQdlXfNFeDqH4PCTZ0A8QUyxBIhjMaEoH0BLdfpRT9q5uf
NHkhcZA8bgqIlZ6T8GJOZn73AHNbqpTM58Sej4/06Vv5WiJAt32t2BB3c1uGkioX
jMNuh4k7v5SC2oHNhtqD9pvk80vmPoAzHAPeIvIF7dPZ+qcfcrp9PCDMKhjRwiuf
UckojwPFXtnVairzidj7vUIWt4f0ZW8QXE4XXyXYQwqgUFlUtR/lY8A0Ht6BJ5qL
y2y+e8xUG4tuZzBYEtVkWdPw1ZdYD6mYJP3+Xq1/ZyIHQhaaqDeWJIKR2tSR6nqR
ysfpoxgcLaie0y59Bo8k8scdJNe6PQHm1mG8hpOKUGP/Ta7Uz84hTPyUBdm+uPd5
XQ7xiKd4mffEmGMSv2wSN/928yIQxmqOlPa0nM7tEDYlFRHfA6NJD4WDUPJqjksE
qRXEq9DdnCNaGxfu+gZx4YP1q8sq6zR4CfeCjuD3+pq4JSnkhGS7yXx4CiJzeTX6
B0oMgLzDUhHH8VdkxPbuNqnitylN37g48OATYPO7Adg9FJWiTqPa8Zy/f7uAU0Do
wH4ZA/IfPm60J75ay4/WBFH3RVc6JEUSx5TAOxoUEn9+rwN8DF3gxh6mimOClwD6
M9l6RYkQ1gc3+G3Pe3TyMEFNxHbuPnEp17/7v+qIAxSa2Rsuat+8XflFYpkVfipL
VrZb7vT5QX3lwkZUAYjMORNnlsb7DvIMe6fFJEZrIChzYQdr3aJo7xM+Z/NE/IFc
hw2CMGtIN1GzHwpj+wJVtE1FsloJNOOSWYKAkCEdNsJ0xgAEyCXbEhsWPbry2RQt
xB+oYF9NwURHizG3DRApipp2iVneuqB+0A+w4+s2BWOPaJN+RAvjWBquYHpiPc1A
a1tKVxyNv7EZp/fhQp7WOpMyKyGjweIQXK7OtxFCu9dFOLjVkpvJ3W/kGiRfMzXP
oXxxu78CcwE6i7Zx48HwN3hrXi3m1UMKAJ0Txz5lXodPxXUHuApO4iDXiagy4vNe
xvICS+OT/R6NqYLQcHMvjs272kFjHsG2YfhymAp5sZvPDEtjoFKwUZDmHkbUKDuf
ZoTRgf6EbHXmCVfY+q1mgr4f5/VcpypUtYLw2zHbkSdFMry/epfk3Y3IEXvkmaRr
pB46E9wymm35hCzLqse6bESysM1mjk0pB/5Pjtm8yvYw6dEhaGTqXb7a3Ftc5GJf
uv1S45e6sgGx9KNM/yI0LmuzpJ1DW/nPGie0J+B75113ZCaPxSzUGsNYea+AYq07
PD3um5HHoscAW0I9Gw115F1pP+vi/kFXfGOwEEGNzaUue1jObTSVohHTtPuu+A5l
LfG0Wk6NWRSmaRHmnD5HVnyqPGFSSLqepECFIs8VLWn+WqF+/N59eBzuZ4tD4o8I
viZ40gBfRXuQxd0XRD4rtKVuE+vcAH8yityk8qaFO7XBQ0mk/My/J+Vi6k1WliB0
LTgicPcaLxY/C8GSpU2KLB7PyBvKJm8vuxGQkIac7TmdopdluWuBPxAFHz6pm5Ps
GPx7uXV3Bh6Ji/Rh6nQh46tGRDyxqQpAu1Rdyp41Kr1qmvaZaT7e5ulj8HhvDKun
KRyVCwsSeMqNt5KGLIkwG/vuxTsFWSqyR4oGOguoYLh4KA0tQ7HZxK80aUySzy2h
xmRv5WL6Skb2U7oxtCb2al6IvagZ8dIybKW0CEqhYZ/BYlV2ROtvAC8+Z+dKuOkz
wCnxmN/RLzKtV26QaqPJgSIECGAzHMiKADeyIFQq4TgwtlTqiuP1uTSNa7l0cDy4
lcricVo+Ylq4nlJ5DF7zMzkETmlJpnx8lNRF/dltPafwPsWh/wsMBUbLC3oAyJ6Y
N7StoOZUusjcCBENPZ7RZT6B5phFrSM1v6r5g4aSej6fHNdhmmeWM+c69saKly3f
MxdxX05ZbVAN0oM0IW2LL16LEVchgw2P9kUDqhnzZyQToz+K873WRhRnG8Ehc5XV
GGZCRfZmVBrFPab9gfkDw5yqkkjWlTzl8i9IYt8UUCGJxyYSvIXS8EY+LFb84Xd1
I3mYTlQywFAKfldFsNV90dLtH3iQuECOP7V8TO81l3m0XNCA3zuEBaSOEj2AX21z
eb47iC61YO34DEhHwN0fZWZW2DYCmB2slm64flPJFgx3LnuRBJZ9k8iHFJ/jaxwZ
dnIZNlxhYBy962VF/Pi9aV2Vdc1gt1aCTW6d+kiOIdxY5ySximf0MzIS0e/gmJyW
E0j+w70rG/l4RXylfwvpKAr8ZM/be1U0QSTNPM9Qxz1LSpTS0APfsSkt53DiiITF
+p4QSDo6tu3kBJUZwsfLf5W9e9VShzuV9fl/lGu1jx0tBNef4GOpVr9RTdk4DMT8
aUqQKiFpCWznWiFRt7K9GPAcmQnLaD+pIILG5SShWgd1ubYlVab5DElXLcbRTZqC
I0bBYoj0AoWyTKnandARgMt+glGIoVXJiQOfpXdxJ2EilwISqU7KNNO2fqd1doHH
BNQFLJ1Y98vl9GlaWiJ6VwAR0EfoWnM9vqXcMO8wUq3KQA45MERQdisE4auG+oOv
irzvPRtU49XiLhDyH6OPVVrJA34bqsm935l2ejNO1H3SPe8KiCNuC5MXvw6aYVKh
yUT+f0gDd3GrGdTQZEa5Xqkki2j3EzZj1Le7Zlq3Hd1HLBj719oFr4jVuhm/I9eS
ohntoGwCTcE+/HDoNHsEU7Qri6HCt7+iFGOxfqwQQF8mk3ONC2bziICrIK7lPr3y
yR8ZKkBr/byWvzpEXS58OnaOfcbKtA6MzatjZJLG2aLcjO3aDguG2zPrtVTqGvyN
Kuv050i2Cmcy2v4iHzOoXY3FBddmDyHiXTunReWbIzX/tQekE2jiEODQQ1tG+VvI
Rk0RAz349K/mgcXDCLi7dVgq5CxInQSSq+pdEz3CxDrStBbm3SE/pc/KyYNSKPm+
z/k5O4pUx6IdiZ6DC6O4w6mHEKD/6+1eP10FkH+xPxzg42DbltTl/tvokhAcIOKs
2avwQZ9mMrnf0uvH0Z02SkkscURUgy8nOpfD5KHuokfU+pXFzJWgg0La5vWkJPkN
HrdyRxNFxY3YfDTs9QZDV5bUwInKoZCvlcKiTbT7b7HAja/SopAygFztKgP5Cpgl
04El+EX3HBsEHJ84b7eQvIaOdewDTIPhhdB+/TW4krXNMO8aAx+uwy/Lrm5CokWt
88RRady1Wu3Tm0xKOvb4hJAlIn3drY7aPpSzIg5fU0giTDr036oQibPnXHcMYgkO
R6Zmjjl2OpilKXnFaHYTZn1qcJPZVRohVCHSobjszy1fNSB7WMshvQmVs+gDPRDY
VS8LulKPaiZLRvVY828krUmfY3dUKALBNDziKBJqclpazQH2UkBXJGfJEhuw/tSS
RqXpnBzb2fj+bTZXUkuMyrcWF55lQ0SG3N7vvqaNClkdMKM5uT0ZTIIC51e+JNMz
AS3w7oYFyYreoTcv9FAIICuVWcVYvn/TKTFr51509J55qB+Ccvte3KapRN4sawEm
KEmrXpYyMlJ2fdKhGRfbeViFmC3EOucY3vPwldHWVVmrYzRRclufYyfHpo33RRCi
UfO2lZnr9PwwXinb5tWyL3SBOxw0NTRUYe75IybSWHYTVngSp9NMMymAmkeXb0KL
yhVpvdQcrd7cSxBzlKSEKTkPObj4Kc3zvwxaimLq95OEBZ3HH3ADmR6JuFkTRPUr
wiVOPUSyibNomGWmKJrh1zaMXABTjVNaD9tUB7vqx4cEe/1Cb3Ej628IahqNi0E3
cTAKYgytNtcHj5SY6lSeGN7WreJKW38Mxr4zyncku+mq0uVvKRndqPErpnd6QYlw
qaX2j+qY1IKt//4Ngj/HpF1sG1vZN+KZ63VRRSCUBq1/7N/7GEpK+98OIYv8Apx2
f6+1KWQbO7l6bft79f1bL66ox/AjqV+vu9585U1gf1OpjwhKGW7sIrXT8Yg+QhOU
ejYJ7nA96WmLHH+sBN8nJdPXp4BvxlF8ttpS299O7i1Y6ZW6ehgJ62sMZ0QEaDZL
jtW+aVhPNFRBAhEz+G2RSftLKIcrrAqq4B3+eSeHrGR7ZupT+jZwyRdzo/PT5cbl
vvvIFC8PdnJg/jvPu2NODFdtF1UlcalLyohuvH6grXLji5fbosYYFXA9KoFDuTF7
AajfnpP+aTL7Aj4ARhhcLn93ulzP1u9covHXgjr9W42URkfiIh9U9pwO6W1GDZ5G
qIsSBZ670lpzZTKjWvGg2HxG8NYPVLI1QK9+fGH/laagyWDBpDO0r1TMWGp4Q7a5
qFc6R23XjhNUf3uDC3Bpz/xX2uFlWY7f2EmZ84VXQfRlOnxs9E8yzm/waMx2NkIH
vspNrd2jygDHo/WIuao719Uckt+xsMYBcp5hPV9h9Taf3ZBPjQvu3NtBhAgw84nc
RC5kJfQmmTjoIzIUXl/R3hhNi7Cw9mtZsdcNcl7hceDGuSMnEW+UuM0gq+1jCrOk
oQZtyWfPe4fMUxto5eAtRKuHjmT5nyY4xlkpqCIesbii1tF8ceFpNlP/8sd8SfXQ
nSx43lkaB/Lh0W8bfReq9wNcM5kUGkZopfiu4DxBaYtGdn3BVhX71p3zTyj1IwMq
S58cELf6m7a917eEuWgaoYnc0SRQmnFdHmW6TKDr1RVSpSwRIdvw3TB82lCCLJOK
OPW6qx7oRQdIikX1FHSE3D/3TK3Pth4HkupHRn1wkxYJsRCwbiLJuFnHnyAwNmKA
KK4lpYissgWKXV4B8giQO2KcdJDK80YCJfuFDYpOkiaO+v/xUAmjwM7LzHYSsFS+
VSfIxvrdHyrVhrv4zk/Ttxfi6c0Kcy1RylNb/MG97ufOKJqpIu8hZWjvQnozOCAl
Mas/WKPQYUan3gDcdnJeJ/4RWLpPfFLufrPKiXjVW1TfEj6F2lj4oTbC7P77BmvX
DSQEteYjoRuPAGADv17mNAHR6OO2nOzT9Ag66VpLpodazCcHyj7AtO4eLV7oyzN6
S43MSWaE0xuhwngt0jlrgwPKQYhuaGThH6aFh6l45jUAjN8frkkGDOIzVxT3y2Qv
L+DOhVksjRP4WW7dxhsLTmtgYidY+KubEO8C5bv8lU2ym8aVyl4x+E6aygN8RJZ5
N7g8B1o4omVbwc6UhTp1C8L2qCSTg0CLzomaQT2xOLG4kq4sM/70C6GUwl8NX+dC
VuKLcFooLGOtDoTaGf/4SO2clu0Ac6iK9MF8iOmReZpDVW1tw53OlFkrY8JmQGwN
NB5xlUTElplZiQfMqmk/MV/4EizXBQWggBEkQxRkfQUnmIy/uQYPuDUbAYiUZoHB
c5icp5pij/ic0nL46JuIcyNlNZYMeN7CZJr7CLdGhdijfzK/iCwo1gOgmr4v9Sla
L6wVsTkF14JOpHpsU5IB3D2zZBeNohyCSJmNMyUE27sVhsC1mXmh+Lvg2AK0QNH1
qhNXXDpqFztHaXWrCnDcd0Y/UHhEouG6K6HvBmqBTPaFvaE5UkSZ22YlAxc/G1Cm
miVGJP78oWPjSktmTO+7q7QpAk8+2O7C8jgrwzbC2+kTgf6xwyYfZXSWoHA62f2n
nGEIU5ohSX8UnH1BCQEAq8cZeIhcxyx5ahLsFe+NpcUGPB4z5K2FviXYQuG+gbsa
KeeqMQDkjQD1sI83nGQVGwEOcFCYV640GCsLVNPV8tYvF9kp5A2493k8uCcxRK63
/zbeCyiD4WYd6Uo1GNszIB3Lc9vm3jJRoQsyU4FRU8G6PWo391gKW0mmHx0512NG
gQvi/TzzY3o8Gt4hZbyJB9JnjxTQ5EttiM8+PTz+ujHE1Ox8wzEx2fR5fJ7tTXXW
EZQLTwHPmeDmSV1Oev7WmcKvY1a/lNTZCy3pcTQVI0XoaxRMD3Oh16+tOo8g3K9X
UErJIvq2LsGRL57lguaDLPtAr1u7caPEyKLIsB3qaITiT4qTss/WaogZnolnX8uJ
lHWvfs53eauGJIf1ky7x2nL1GD3jGH2wMSCGbt3R1mbHFyhUP+hXm6Tj8m++vA7Y
IGsG6/1dzug6usLVPbDX1AJjONiar+KzDwTBitLXpmXZtQ3L0Bc3w6VNf0OoiAMC
148hctdzXHwK4CW4/oYmzayqdjQKcOa6FLujisk4s9s7zu7rzXuAvl5RwWRa6GWx
EuQX/CtOGbgxWZxWpXVe8VQNrLYuz38KFSYz3umMVk6jSZx3Ztq4m1B3+fizMDYJ
WjidgaM5C8k4dbY14G/1yaos+vwAnv8VbHd1O4XQfqdsCkxbQ7Flf7l3hnVvdeZi
yeDTs+QNLTnXbzd8drR1C5c/k+wJvUrL7M86q3MP7lHtmSh8xQpxbxWOxGQq4w4h
bdSleUThTaS9ogIseJiYNxbf1+uUBg11tVgY9/fDh/sFbixmf9rg2FbHpPg6+dgz
in3YmzmFgJu23Cxj+DygyEJrsvioRFr0GPtqIfYLelJCJBv2Q+HFGNX7DOtijB6T
Q3p6/FTt3wyS1YeJ0NKb9xwEYhVv6PpG+U5VHLu+yvHOTN3OvY4I8o6PaYBTuiFi
DAxkjFNB4yHHuPqcqsyE+Og9dvrVzbR6u6iEPJMVMCpZ/UqpiWfCobZ2diYAzqUv
kSm3ACDjbOiikYUU3C1npEiWjjD1bOyl3zZKZOT7MyfQb/Eqr+877aTG79GZgfXx
PIES3crTZkpyh+CNS7+6NgztIR+WXocdTKaPSr0ItKBiboxyZhsq4qYqxyN4nCQS
wOhnFhWDvDqyQrZCv/uZCsQaw9Awm1x2A5O4GYxNBQXJB0M5D9/B7YO+PzqpjfmV
9Aacfz3585d+83roLC0nCROlXDlSMSwmFPzB+XOJGUP3ih3EcREAXBn0kjbnsUrg
q72AUVYBjiFVKQIraoVblMyTceZaQtTbHZr7/9ThLqJW8lF3jJ/WQgBp2VfibEFN
szQvbB0s3VnFo0ASPb6iMjS90SsixS3X/8eECDYCmqCFtHc9jAyfW4tAjDMiwfXF
bHpHOabd87mAEGYpBBzsQcV+Ydo4hcXIxPb8RQ87CF8VygvbrGXcaA86vkmMgfXX
mk1qwDu8I67fDMi84KydbSs179KYvPrshISTQqL7u33HupmJcbtzqGKurf1Ed+UR
9z3mHcowWHZNoSFLJHis6HaeyzJkWVGKyl8qowMMrtwBx944uJgrZSrHubaGRzyx
7DnlBGndVvgR+D9BYSIrjGTqiw57j0zGbjGL/Bd45J5874DB+AnmQSkipA/w+BID
mXzBFSxiZCfMoApWCbIEgXcjVScIUPtSBhhzxgH3MR4u2LkEudYJ9fOe79tJt4bO
AZ/FRwBdM3tIfvtfu75/TpBdX8PZkCnwTXQr1HGeVgD8H30mjWk9AWSZByU5fL0c
oLXJWmu8fBPQWQb+TlK+vDFsNXXKTbozOlCRYPPC68LAgO7ugAppTc3PQRzxj/hi
G4Umz20xw5C6u6tl4IL8PqoWNLiqVCVTYcC1mKFgkbCV9kYrfIO0dhnHR6FHE+VJ
VlonWIS8CZxMsFSZlcVcRgHrxRzNQ7rvO15JraCo+YkIy5Uf2IFYTNAY3dbusvSi
lPNrgdmf2EyGwRT3ERk2pQlt+Gp87gYCRrJkzF6FELTeNaEyJpsEjWJ6vGIQ1D6L
45dnpUwnCjFYM7i2QPK1fvMmoBJQo+QVFNs7OhhVX08DxCTucXh+VefkNqASOpCm
H7MMlQajCKO+Hh8UvRbz3H9elB6a5jywu9DT5uQuOa2Iw2se3fVRfnwKAI96V1Sm
WZh2j1q9QVj9GaF1Q5f0tHbjQkByhCAq8NijaAwYGV3KpGZfiYKynKSVf2QZClZu
fc91GwZkXs+6d72czOVViRBarX4wCxocKw1XfllXOrpuQ0OUY1ijZwY3a83XxinT
SXhXD9a7WirWzMdvkxNbFaomCZspqLp//OxVn6/8g463jCjD3WryhsfkPF+y0agx
WLzkU8WAW3KuYCtv9GhdRV8XBxjwhXRArobdMr/ESX51YCiHiBNwGAuTAn0Tl94K
HnLdw89nAi3IL7qm8vPBbc6puG3a+doA1xUUBWX38xjmwD0O6qI5bM6OUiK2+8//
cMGaoTyEu83TUD1xquldM/QXcEiqY/TdyLvRQKtipN1sudFQukTJc/+Je5hGG6kf
VxxJmSHZiGOgnO/D6AzMDVvJm6sOx20Xvr55AzQqsQdYaiskQ6w8KCyO020ZwqWO
C0W416nFXVwz37r1VyjyKvgcHMKi3uRSvS4koapRlUVgsMX0ovqItwEzh1DdF5mq
gGG8fts8vU3e3PPLqUvKK7BfUY76YUxDm0SW9L7jVcixOl4rVu4CbTYBqNwesDVo
9d+kGsfpA3faKDFbsyTUDzW3O9D921BVMUMEwdC6nlOeyDOhMCRWH3s9dgn67JKn
9SB9zgRfkPfAMODYjLtzYGAkZm1PVwvnT8HURnOzfNoh+6Fz9rKtMtZDShgsjGjh
MfVywskiErJxaO8Q+YStJJ6UJ2Y7ICucIhe5kIggscc+yUX5aaOMgj4t3aLatnDh
VQVAawPqyQBD0bxOjvOvHgoLo6qGJg+EEfeFZ0mXf1kW0IeWHtXIuripTkKu3mr9
dF4/DY6kM1zhYrASEab0aZRT/uLb+37Vp5jcY5pqt1ryiEDab9Z8bQF3Z76v6Ya+
iJZYqEprNlpeG9OAfyLFNE0n6GPRERd4ecOFkEER172uTGJF3St/8Ba5SQ2m41fz
qGwnHZ6aVOlJmBIO43m7w0Pis8Qi+CuubqtIYOqZGYvpfflUUGhP1YO/CvXZFXJf
10XLJ9Pqi6pyUyVEirr3AhPnHngKKLrvzguqq8f+Ld5WyacEtBLQW+xy6jK9pmQX
19bY0eva+ty2S6+zF11KG6mXst3heD6GVvvu73zvbxC+RzuadPuURF0Uz/Y/nD47
aeLykSYt+XMwn9Ckx18DNGdKUHinXuWNwKHG2bKnwzckN+Cv8ZhnftQFTZerM6jd
EGCk2OotZt53rn8RecjoTEVoKL5OKrVZaTtGC+Kq7k2CAaraKr2wuLeinkuUgRuu
obxCk5eM75kDoFaOIhV0SuubN8vAg+WvJGABdiC0N6tZnC9PKN/LX3rBvmmLTf1K
RQeT5Xa3ckaVV5JH1Bn3depy1Q67jQJ62XI+XEJlAAo+9xaoM/zYXIcw+v9b8J6f
oe5FxS2/Fd0XTkUXYh0e7UkFvt/VYSZBL9GXazWR1H05xlDPmr5H1p7JAPnpLR0n
1AH6fhPgKl3npshgwSvKH7H8BiKSuPECubBE3Piwu/TTJ2QpjsXvZpxYGCE363oR
zvEpKxA7BCmMwuCPAQoATrx1tjHuUHaO7DD1b6ZPH/AsCjfXqyvlrgnEL2Sb4kGV
VYJwNo+Jx+FacwY1VRx2d3eVuTrZ/oUDpzvVxEpAK1cbIcVmebRP8d4JwFj7IciL
CIdqxdQI2yKw6SztPhWCiG8eJWO4Es1Pwk2zc/DflcsjLuMSHpUbYLbkeoBHVAnm
Vk4Y+6TmFeVQ6BnSc9UirYkPQMul1b+u1dwYRWz2G4PLDFRhwwbpOFR9AMGTbkAn
JviJcq+AM8KZQip87XdWN19ckt3RrwzwnRaMN+lPmtQaIyX2jodqIsOV5tbKgHGK
tyCRGRJrSZC+EJXtgFVqKss2Qm6ZUmSEKE7EgtowFITwAGWegNbecP50T/KeWvfH
55gOmXwbIjsY1itbkhk/0UQImY2isX+tpVLlA5bbg/zE04WUCpfzFmdaYbxXWGSb
+gEL995tikpmNPJxB6zc3QKCPTdo8cUN1QINwu+9fhnGWVHl5zWmZNfi1DbYzMQb
+76g4TdDfaJ69Dmdds4Jfsnf+gPJTfP1Uerf3Yp6DaeK7YlEf1eplF60ZXJOgxun
pI9SzR/YfgPpCalOnv8cBQ92tPn2VEizx98fzSeMx57IOdzZOJiCC7//wF93+H5X
wf3tjzeVo7O4++IclTthYsa5TiXbXp7QQ4Am9fsEFx2MMhOwD/jsnTNBMILA3S5m
++GVRYC0UhO3jmtDsP1fmEuc3bAJ9/WpK4nUNRXjjGxv8dBAGQgEMzQv2/cD/w9O
9A1Bh/w+s3kwn/pJRIkKAWtg1Yp0x8XXWrGLFFFGo5SbbayMPqWsWxOMg3lH8oiO
6Goa0ZkmPgPchrM1Txle3/JnfKAhkNS39O4tUqzLZxP7tafFxaQQXkbeYo0jZoI+
iDmWC536e+TLb46zz7/idmd1+vQhGNscYabN7SW1o3465VuttYlLeLH1Gzl6U/eY
8sfJs3lGZplhfLSeQGa4LOTSUZvmN/aomSwqFiNaF0Etwli1rUVs7VgG4xroaeRt
Pvqi1aLzj8GUrK1J1eMxEH8mMNEjEZrgTS1L6g2GjNgwzn9pehf46+9SqhddWk5l
TxvCfdCGP7m0VNS+u/tpwOL3IxE+5g/uKhzkfwV2C2EOtv+aeXcV7zkdQ1/IHZN1
AlDVP2OiKhpn7WIMe+npYgQgmehDc6i7nTCDhvGm+Qr9wb+BB42GRDbWyZdU0wrV
Lhz/I4wZqz2IZRxiMOGwEpQWqEFBF6nloPJOukAnHfXneFrO8e268gAVJMBaCHTO
wgLzwUgUabBIHMz2YTs2u9azsl1IDDHLiGW9pIbm2h4L8plLs+sVa1DQ3K+Vpt00
Fv3xn+ngMm5u0A+yKvHa5KL9vwCp+7fFIC2aSILUK9w5Vvb5y/M/NKM7TpgiLWMz
DzXj81fro1webMxaXbOwMXyuxaS+OOF65Wh+ZhR0T/eEivSr+VQpxWyyx+bY8HZ/
hdf8YZPgqTzrgMBcro+W9sE8/PER7P74i2MD8P2Jsx8YjACEFAap9w/CQyFA5V1f
9lsEFrkqPvkUSi/r7+dGcqNZa15N5zR0TqaFV22OFdzWw87/VTF5q+sRhRXe99Gj
6gD7fBZIVqCtbe0A0j0sSHJ5oAM9Jvb6vErGOQfGNm++VRoyEwuulD1KE5y3BgGr
gyG/icXzrZpQrC9VU3lt8B3EZTV0019ZVZDUp/WoxrAa5t43Hibu3WCwmIVXLVp/
LO9v8ZLEjzxASC4GlAN2uB3nASZAT87ebBRyvBePWg8bch3PpdRcEMTGFBigXHO3
2EbeIbH4pZ17ZNZ4ghdmrcUVUkrI2/+URbLdB07cJLV4W1qqaMz0WL92kKWCBR00
aBvtuR633jKRK0Mo9e0oMKk1spu6nlL8+r8zK5472KMTmcCyJHeYyEIJ06aO4sFi
hzVFHBaLjDr75a/Unn0XnuTdB3crkQkFBQ9M/vfTAXH3+tI4F/pvjFpzTXqrbcaX
RBFE9wj3FJtJrGcFT5ApuUI1LBzwTwi4YSiIcY5LDhd0WzQzYeUabNQPEurU9ZGN
f6dKdLm8z6OlOlM6d8yQ1oBUfZ4jcJq+I4zuuFS2z6eFpE5abDYJ4eLQjke/7+xM
AZ30v5NZbu7Dh49PS/VMlAs8R37nQ2Oq2fC38bTqKyrnEOu1dOoxrhKq+TMML0Hb
4b1kWoYsRMeu6L6dcsuFejDD93S0haA5mv5fD65l9kK+2i57vJUOPXk1vzqA8tm8
AFUF/kCXlLeKjinD3wWxRth75hWZcqRfDhB9BmUX38z+Hv4J/OTvNmRtjtrq3Q45
WviA1OFPiCFoHQtBJgR+n1GqlpXSOxlJ6oPJA8dGGZJasKDbSBZ51N+m91xGTKah
RV62kfa+tC6/w0UBvZXY+y6yQtBzhGI0StGFhttAMNQzKJpwKZ2kR18NtSIVhFvd
g8/gHxkc9HL7qLUTI9qOA2Ca/eqHPvHBF05C68HCQYwnvb6Egf74JrKTxaz3WBQ+
c9gZky/WQa0iy7GiNCsBWoq/fl5MdpDrcY8QjSQ4p2p2DNcjZSeehnsSnxbKqqdK
pfKGpzgbRNLje8gqMuhj2HtoAxxQAQdVbZ+Aj9sZOM9IHDZt+SDlBWAjSnEhAxsK
ZhGmkt/nD1h0CfvCXr/2z2cgJZuIzAaCgceuqfUP24sOkKWghRb4bYRV5VZMyGnN
5rpt3rioU7QN4GMZuPe8ggReSmwYaA59Zv4e5CJlFLFXgmd2OZEON/CVIRHC6b5/
Nrguv3ri6048vTqXoWgDHeXru5sE342jA/b8Um5tQTJUigRvn8lAqjw08i6ZZBWq
tG++RA6WOZHUFmKAFKvj0CWdYDgohTyLp0fOJOcQPtwd3hkuKD3cRDzV4secc0vX
R7R15ixJZ64RsGuF5i6/UJu0WKFnfVgFx9jh/ZI08NhBno5f85f+DcIFcN5wXfiF
SQhYSlUBV0UVeMjcDcPGj0mC8pBx4ej/pfq082iWoaxK/lNE+ZH5zvacui683VcO
+WroN47pKw+Pk6F3qBbXydSFDhcmG5xwNuJfQqElh8TGgzK4DUSn6sj/mTAHKxfk
wx0d9GHYM0N95JHUIJYuMlNsl31hZvAuwEtWT5ZeOZpgxOdUHV4eUw6aAB+GdZcc
W5ci21kWzWgvxEbJqZ9V0TBXGcKWP9vRnAfjT+g9EPguoEGjnlvvNlOHQerW1/aZ
nVtOFNg1yOW7JWObJGjrOF68ncRczZAFo/2cC6PI9LdOK+CxoofW0hqmPTb/TAs6
3wX2qYCDCM1pFWiqpLyeQ3AS2TCoG/rxxUkiy9r0mMYwILPnQd67A8zbR7xHXnWa
OsVRBzhk+uWGRKsUAkCknNObZ175ndNz1TJiiv9C4Spx/D8MEJbZPlhC730qFP7S
col0tmSzOwbCnNQNjgn/v0qD6AJct5IB6M0TmjtOycnhpJTPx0IMTtrBmu0Hud9g
kXwwBiJ+0Yb/AnA6J6FcI0R+iSqaRAQPk8uubX64sXSRMhFZY51AZutCoAUu4OPj
MmLWfQz+7H2QAU/Dks8Uc8BW1di2gMKKC+TIomY2bSXXQ0nDAlgdi6HQ65LDrd8W
15K4CSCnHiLO08+O4vm5sKQWseK9IYHoXDz001jFa+ReQUBcra561HvoQoXNkt1a
KzVbQ+l/3l7yvYlSRgfB3ue4p4H/mSrhJX/cvh4sSNLDdaoTBmtjQj8BWp+Ioa8G
mudb75ypl9NIoM89HU77xKfp4fnv4r+gtly5XM1kIk/mIv4VQWQUMZs4WSl1jMQ+
kwsdW9dulPVEsNbWlEdIub9Pia894ipvaDArqFZ5wYDyifqnS+q8KL/JgeBvRtz1
g8dSGPz1McD9rz0gigKtY01XhZV3T5LFD0tRD4/VuNywmX2+osabqX28C8d7zaEb
MnySCTA+bOv5Ysvhv05Hmfhch6vk1VlH83zDR4HyZrqRnPAa9mwx2cQ/srkmLiRD
PB4TkxdYJpSTOPAf1aBWOA6phgD2LGJqEFYJSAMD9ao/jkgHjf2kNvtVelRU73X4
HbOxkCxQfXbkt11nV/ql/DJUiyZzg7Y6wH3mMBgmEfOkBmYB5cS77bAoIHqMwIWr
v5BPnBTv82D3QQUounrBOrRG7ZcR11JbNx4HpBJVmzXi1VYOWyhsz0Zlunzu+kyX
VcEp8e3jwMdCSbLzbCTYbh+dpV/+QEo5JzVAr6jQjyYjC19Z5p5/u0IO8AH/f1x1
HOnNufEyPAmWY5jqkQGSSrFCamJu5ywoeNX6/rCB7rIIx3kD9YCngD+W3Cn0edeg
uJktSESA6wuA3QFYhJ5mDoyubyV/3YUNJ+AJbpAuPKYIL+de9UEgTJsIaWIH7Zfb
eXot3cXE5zI69C/e/YsSqOobDanrDsJAleeVo6fuvSoUSWdVlxx8e3WYD7JYWtMN
dDi9ttQIbhhyVQzQROkO/ihijqcHVma0yQVRRQVugfEoVDjD4shFRD9TiQ1Fvf9Y
ji5FUuJ6bx/Z61XaDfzlhRux6Kj0h9Mdx+RGlIvFYpuu1IoFc2lExKW98vBANPK+
+v0LZkUfN5TQUQLE++LqioK+J33+a1bRomza/FpztKtWbzlmsdFPxB2VXQL0U94S
D84NNz29/k/hqimKd2C3dWhhD3/pyvKmES0p9klET0H9eheEPFV81LA5kRMracLW
SoRMgVxOk77wctV2GFfCcwI346mLLiA3Y4+5Ea6Wr0bR4jIxh9Udusu2PkWOcaVk
BNDkNZTn5/I0W88X3c0gJZYzQd32XvetU0MeybhMlWVfyg5HHgkLyi2+x2gJBEHu
CY4RNLTiZCx1+oTgiSt7GTm+o/UGyV7qL1e4U7tyoFJOvksBH7m37vx+b5+LVgY3
hLVmeub7dxlUbKZnUA3pQ30v1+wGjs4t8HXPCkiJEXS9EHNlIITFxO8KHWVvlyKP
GpbueW2oSiL9M33xCUEhvaecm9DCNx0YWbqDzOGmuU7dXV9Fl9PUGGzF5hG2uu/A
k1zJ6w3CJFi8mgnJWfU3XuC+tx35o7vBX3Dkp5/SvUkMt0u4YKToEeDVWw/TsElk
nUgTV4o4OS9ZFcy++xrpjoT6Z+xwkFJh74t/w6BKq3d1XpIEUbI6uBlZmM5O5zBt
xSWucvzt7xMqBgrNA+k2i1lvjGcMJIgVeIp17yWgkvCxwlYkLMxNcDlNkq+enLRN
PkE7xeneNdROaDZxL5M1Sn7Yv5dfMA+O4sknklTRjCW5jGYcvqkz+G79Qpg4IWEU
gIR3FRjwzGliCFoEAeYV4yjPBwAsTIb70dkbnf36LC980cg8ZCx0yXt9omIfd8Q1
uAdJ8PYbgLmkmpJJCxnCcgHMS7+koi+KdCcqPS4u6J+Qub8pnjVPTKgdyRqx09mP
PGyZI4EAgTaonrEMQkMFztf9sJVBok1KvfklxLprm1NqhB78DfKKgzXvQPm0cION
VQSj0EVF0r6T0pmYxyv/pKkWvVBn1WkUrkgy8zNtdTPIvEJf2bpQmX7DV/DksN7T
L6QrbQhyJi+E9sSXxIi5otU5vYjPCH4FcWPSqyjt28CMkShqDMY2oHYc65we4eVO
KxP8CVRJpjjbCYAIQ7CGw4VPa+7AW1s8r+4oPkfx0+YWHoY4pK0NDKnnkGcyvYTG
HEUqmFAIN9LC4YTSntetyPA83gGdcYpbzBZ5IhF0W0wku2ofPaFmiD1L0dCXZ2MQ
nUcbCwdQC2pfXwuOc4bRo8kqAXZdVzWBBotj4WwM7KPzihurcavNUFyCeQvzn/Vw
XmHzSJcgBZkUY76IfoYxd1na9O+uR+TecnWh2fyYnq19vJ1UbXfHVZ6lhBJsZRHd
0jtbcPDvsY9DNlRAfyNaFWtrrqdsbQDELaEpqo5W8F5gVhzhY/OoUxXt9Tzqk/Lu
/Tws8sr723O0y8EweLI7BHHwxa3rIYYQlItQ6oCQ4bdnhzd9GMdt8sXCwlAifmxf
wctc+jiG8tfKOvC738W8rnQ1+9brUvqA4ibyUfTspUWbfAavuVK106DUJMKONVe6
NFi1QSOR35dscCMPiJGHgUHFWKBw+YsAMXeZZNqH2pNJ1OkMWWdsTr6ufppg1wu2
0I4jxu8194bS9dFcW+5mMq4eLAkuOU5UjdNF69Jsf8xnr2wmbU8g2PyKR/L+hGuj
rI/LE402QnRcfn0v19qLfbL+oYmufqmcb2xFSkqPMpeWr3PyWDXjHoAwySn3wQPV
2mgjbzb8pIA4OGJG8DcwrRdCav1vHJSscxdoy3oHzuTt+SUPJP0Tyks/BgE4QcUt
Em3nDy7vgU3irVSrqatNrQSCuujki3033Bd7YTkLgk9pLD2mqDQeEwNAj03tmY+W
FRrOxZLTbQHYmNj3UClyFE0fZS2wsaRtonLjEmxjt87/4Djly4iGpZZvkF0SBAPY
4g2UhkXeY0dwzA0z8d1BKupRm+uVznE6fhUUiduYib3pfNcywH6f7cKct35YRU6b
3Vr299GRZ586gW8uPol/pL1MVtWUG/Ea4fS1E8HoZ8Kj44sxmp4GvXDeS6IxwckJ
JKApgqKaTdZKolYmt01iaFZ3hmN1vdr2InRtYKlAacuqOMRRP3U2eNgghQYdpwTh
9GDHaALmP6rqG3GyT6if5FbY2uiBTkgyEiLOMtU4JnxhqNemF6MfaBKqkhk3acZv
ilSqFIVjylFzpRicxJdhDOanMSnZaPB05w5+EVk+9VZhDyhHuYgwAArKYjZ8kyOe
jLJDU48qPM0mVUDSMweXYuvV+iacJIvzu1WfH3/5XmkT4ws6g7t6SaWa7Ck8QCS2
KR2kyF4acwYM8OoBsNUrb/97MM6KZpJ45DPDNtgLK72p52RKVuus6kAI39jSI08L
HITXcB2ViwrAE8IcgKbsCgKKb3YL73h4f2Dg8gHmPqKP+WV/YWtU7P6wCWOAdlo/
TrdGBxXY8XVDuXbXAqFiNyn1fcgNg9Iy32Z7jhiQyLVV49hQebsy+pDAhWZqLsab
an1R4/QDzhsDhtnHcbCiRXbk4EXrC0ILRvwiSNFGl8eibdkDjQWypz5d3/vJp18q
vOk0gBPrRTB8F1QaIEsjel5yMqBTkv/KWHFmOIhQM7mDQfreZQcjp+FymoDe3Tg1
/Hg8fATtO5X9qAIfwWIsKYju7GutEwgXf9tTjiOu133ji66NnYE0i3F8SF6h/T3u
SxZ+6buHaqh+FaOwS+zMdsParamEO9BCXsSHPMBX+ayW4rDI9Wt94QtEs658BjEj
ABShhr1c5puS546LobEKldTrt6qjfuVb9GdmOCl32TzAy4SXkbAc4T+ivUCT03Hf
UmMQmltFp4TBbKU7LnlzLAYGiKchO17FTEVzrbtOhAJDUc/ABQgZfqGSmCfWQ7o2
YyxIIW2tD8Vm1oPlUkPP70lkQokw/CUQQdK/gosugGGTREUoC7GewxFDYFZogsai
pDTnOGWOky+C023yLsZ54ymwkEr9cfqMClebzYUpcoO9ysyvxIhWhkNYr/8GmNq7
WkT5m6pFoIH451MIqYBi/Z3zadmgKJPa6Z9818+Y/GEUoEWh090ThAiQSGcefWxv
rC5tFlQgzLWf/ehvfN9CrCslij9QEtGovIObYDrIByL2B508lCkyt3vnpYA3ZG+7
yypwsv4XgqngQt6Pc+nyOiqFdQj9192Oza/owsDvOnJ7dD/LGbLYqFFyCH2SeTaU
0XPfZXQHZx0ZlfwsJXlercz/373YnDUfLASGcdcyuTXLtQF3z1bwfkACcV4NCKeM
rV6H5gUfv/OpoNrpb+lW7Twu+MctSkKx1e2/7l8fHzWP0YxliEgnmZzmByT23tKb
6RrfltvJBzSY5hHbM5RVveqWuHV4r3O0rQer5D6YScZ67iWrTl201p6s9Crtet4j
h5sMJieRoKfWZ5RNKXARBVcq1VxTqo43FleDEbv9XIho4oTEYY4iG6DbsGuzbqf/
nYusaYHvgqzYXv1FAw2z+TXXR8GUxDaa9J1/Fie+5kWdCi8oRL+8ya4r/16DJpfi
VhWibtdgZ+qG00icMofQTZkfNhbCMxOAk495NksyLBCGCgSRUCM5jRJeZvISlBgk
bP76D9MpJsmMikDa82DYGXaAdm2LqG9RVGO35vL04thnKtcmgGjeX2AjgvJT5rPZ
fihX9s09V/4PuG7mrWu/njJWZ3YN1jFcVYO0J/l+bMcRghuDlrxYLCdklbjTgJs7
L/RQ5Xvpa5jR9n2vYnFchr1vQQrfAccWynFX/ho3HKiXe9gvwM2TkG0towgw+aRI
J3IvkT57EwyztcDykHKAYKy3IkpGxio0SLEV5lBi+s9FpYXxsmkWJmRuW+89P3qe
Rio5/XnFt3evFH0FAln3a9bqALw5de9PKsQo7wTyASkM3wNqPaEtZEabASUsvxZ7
YbwYu6uTrzE5XPKeSua31JWKddn4cmf2cb+3Eko1Lw9wq/jA4aMTnZ4Ze0V3ivHR
v1vGDjMzbYNLNDu3opmVW8MYZu+tzDXvkH5XSbMTy9P4VpzjPk17ZCZzT8uEZPf5
XN+MKY5jbtClnmaI7sG+NZ4TZ4yHK5Ua5XQCArB6fceaJDE0WUioQ2TwH5t0CrqK
Ny0/O78gpBNpPbg2VxYafOt0d2HVZNJO2cAq9maAsfFViIfsbKiVYrhh/D5RlHl6
sMPjHuA7HWp0QybHURF5/Ndw/QVLcqL76DgO4KXRmp0vJamy3dxFti+NKOVtRpyx
HYTx2xQUhm13h3Z0S/ilTTwqhcRfbV8ECV0Vxsf4RScfnuYQmn7XvujaTk5bI4Gx
9Bq9RiX0eYX60vSOvtN8f9ifsWp3ADx/Rc14VVU0BdC35FXkXtCGcEhfyMme2202
1A0+ZSMr/zL/C5szwoJviwshgeRmlyh+l1skcbejM3mPiuriJfJZkvIVk7sj/cjB
tfLxPRkb53UvepHMYVGGs1yigRqpyHTG11Kqc85835MIgP0K5Zfr6N2QixfQSujo
3+gvhiqSxqIalhev4rwsyzQhqdpQP+K5j3V8m6driI6rCYqeOrrGyx+ECm501KkI
cEa125JAiG9/8uNmR8j03nsoc4Zx4v1h0MPe4l8DohK1OwEp2BFqsN7Xe86pu+2U
T7oOyS26z1v0nAU14dfZK2/xwOJ02lgDvOW0cgZmdDVulysgW9NrHdwPdcMGrgyJ
VIEfb2oQA7SAOXB0pdMhlvPt/fO2vzPuJcsJPf2qgvNDdOPjw76BscCcywCurovO
Vly/nZIDBZimp9ylZeVkolHVhdSId4kcXVMeNQjgv9obA4TDd8K+nMUwW58i1QsK
97IrNtR69HWqhU2uLJ2lQlao5gCm8ST/R3cyBcZONlJiRNjvZMkkQtGn0FaevjHV
R3tsDzjKm3zbQhfO279NzXuvqbgW1XqYXJMmjDEb8QUKQXzO0fXBtxVOYt/PX/hU
J6c5l3Nu6WyEAWKYcVXNHne28QCgcTH9VcVihwJQqhH96srS3al7L7EaG4PaBXep
G7vK7Cz4T0nCLufcClG1/afNOdvNT+VsIK0J6BYUz0WNxp55MTgSlrqeS73n4lL9
G5q6JGAXhcUVpRlrKNtxFcP6IZg0JyQ6p1krA+pOkxtFUP0mIofnh0AY4dBiWxPN
vk5rPR3wtDJ/GG2zKcNKlQNqQCiXQ4ZypAVtcm1wngyEjeWtQD/0IuZpqI3bcTE/
UKvLtFst5JWXU15+jNwTRLUwHnF5oxiphby3wHaNJoofN+C6w3tpEFj+UDlMTnfr
5gC4T00S3o7kXtnEBOHzKpeToV2Bk9j+pIGCzTg12jpfBN4vFlfacccx1L9EOAHt
WM4OqdIQvQDEzVoFaDdXjiQrVKM/HQBio84jyVDGhs539WHlHBEsDB6WKxe1gFte
fhkoZ11ceUxd5RQgDg+B0rKcHVdVzbRBVxgEqZp2pG07/NXQJjw3h/KDoB8LAQaR
mUvs90a39QoeTQWh9zSIr5Z7OezrlvmwTLGSMIN3ssMPjFzbQxeGrbOxwzRIbvHs
EmtfaiYORBnkjkkY7eO9o3OTfNnDUOqUW4rbQc5td8gWoE/AqJitthqSbjeCquPm
I1RhyJiQKBFHbQ7mKTqgPiicfc4l/lOhU6+jODptTfCV0rJ84EfzIJKaRZyij5lq
B6UtSZRN1NUispKE6QMfL6UZtFMi7ZyL/uMXJjHNGaURF7kSk8lEPTqds11OdvUm
zz0lsGgaEO2IPpuOS7PjAX/RaAnvsqDeSHmKikS4XLVPbE/0JqBaJCRA9osF1nR5
qSUGBMjfLOmcTzbQFV6YTe4dURiObGwg9JZ1jDBBEYri5A/Dlhph7XtqtfPG+vo8
oR3JzkCIPkIT2JntAec6sGVmqWMut1uynIrUIWYZnfxSmPDVzajPN9AA56cFupSo
h0F7+0JHwbeDVQCBoCsqAaP2K6GwIQy4td7FNur7LECkt25cAmszijWk/cgJ9blx
9jI7GpJy6piocfIAMEvLcGBN7c90OLSjfaZUbi5bwutPjviuL0PjEkmCzlB7sbbe
fSq7T6nuARfTIUs0Sdw/4wAdr9sfm9wt7Ls5HdzlaN2pSj2Il76Axtgvuaxk8GU5
VC+490lbDvM4CC8PSPvvpdx3Kkdm37yHdaEdPG/xW+qb0eAmaFanDjyJVZmW0T0g
DF3PALBS4m6sYyav/v7ZeDCZwymmAeb4j08BogD5Tgg/IxzwMUWRvXpqnARoeoWt
2dmmcfEjUoATAUvTx8YZ4XcQNJ5vs7BQSpltg9kqvrd/O03H0fXuQ1bdqkXypv1s
QFw/UBi7x7CIu5qUU/0LdQCIddoTmAq8+dFmlSxglg57UYqpYx5dkzWn9B4iH6GX
ml+ckmP7Kv8DoAU1keiXtS7dT0/K18jZRJS2tbYIhd4qd9ZnoccstJjgLaUMwpBv
YPYIzEAEPr1Lkocwbq1Hioj6ja0K7RV+h/yiXyT31cOVEk93DCDbptEEB6PwIVd6
7YmyvKVhEJKUVJlHGwbWLmpQVGyDAiDByRjcv/wng2gjj6TsadeRAUXedAcK/nDy
iyBgbvejor9JDZy0lcIm3/teEHYd5iSRcafLkP3rmL4KJol023ZfuFxfm6JbtmNl
lLpM9c/NgQOrDLuAmJWtLyHXfDOVmlThbI9cLBt7bKh4U275VXU1YX6Uzham1YLc
+xpdS3cMxYLIAAN8Fsqpy67gMYj056/DNi0GTGy0zukCJWJOGkh7jOnKYzek1Wxv
HlhxpbXGRejQ3VeNmFXwSUE1A+oBs4a+cn38tq7j4cUq0ROvcuVCQ14b67jZEnE4
GrqIA5UEl4e7lVC9izfJeHb0lqtx2jXpizdn/pR7S9WFvdKH4VclGV1/IVhoPNec
rIVkjdIjYrNJQ8SwTNNmVbwhbl5fmVi49MZnA4d74KNXvQrUEzPfMkeye0XvknUa
HatC2EK/08R8z27c6sJbYYITsuhmmEYQ9P5X2MJlomlhftjWvMviY+2L/5mcJBvi
0s3m+9lGCJW1pwiTIC08ZhEPH/q0gU4udzOVVYbHxL+C9CDVMPO7htZ5vhHcgr2s
l9n+j1KF/hVB8B2vnD5pAFTAxGWbooTyOGhzA6jELRHRRXCTn8W6eDUTuyQz17K1
SZT2yeUcMQqcxryw8jfz6euz56YLv9sMvmWrwgcv4nWFQBNrDDumE/iEYft4rMNv
pQEmeVyVIWI7gQTkIVAKgEGzSPJsj7CGDKnIWs/lQl2eQc90cACsF/LDO1AYEcqj
CD3XGwvD907cDdGfOi8cBC+jysjBll/fPU2q8oh/9tBXP69SCJmJtbc+SGKSCvCI
enjAWMzT1XhJnCtysnpRhufJRw/HtixLs9nKljwHX9ffSSzsh/YxpYhEZrLRBdh5
6F27EIu8Gay/keA3YGZm8lxJt6AzAAfABBGFR9VnC1O42I079n4U/IP5ZZc61FIU
uu1uXGC/tXPlEcGkIFSybtWqDDrAEVFHk8pknd+1PS3UL//ZWlctN8m1yPSnMS7i
IiS3vnDzUVKtvpDhAxMcnafcJkQTCxB8wB5Cm7Xhfajf0McV+8OPhhffX/PMZQUG
jlPJN2E7T3HAvLx+4zyVPN8NCcwGt2kqVHes4qk01mnC0rv0MEW9m8zNTWYQ5/Wf
m1/Iyr9AoRyw1mwGOHztbvMMkk0O1I73BJVK/1UbcsdDf9V1Ubam+jLq+Lrm/r2x
mrx0MtZzyIFueefYLS8gw1ntYJIdSP8VRKMtfGWXDoo/WYAKtvQLVXduqHVxEqNA
EMqxDeZgSRZ86+86ib2K5EZFypUGDyL+jnkxs8C2eNWm2wkfMpGWZhVl8ZrGctnL
KxqoBkkMm6BDfvWBJeJKZspORTRtGkW+AWnSqET0iiUC2JARKmsBEJLpkzw4EhGm
6TPI/4OnXSVwmgVxZrLnjYU64GP4iiGTIG6G6CqlkA+IFrFlaj+Drwl6qOjjYBNJ
W5pxP5bUm+NLkHX3yWGev6RyP9+4syG/wzvd4OOhqQV3/hqLrKMdNklKjTzQe680
SkRR/KMXW99dwWiJ0FTIASyVSUdHUPah5LNqSZteGGC/Kx9kDkiLxtpJO6F95OKT
Ndi8ATsHw4FCjKc47FB+VbypFZwt+Qe+zh2duq0yW4StRjz11aMwFKCo461sWtgQ
Up79IXDlp1YCMYL6a6G22imbxphBJFOMzy//y1FhcKtlrQ/9Qx6gnzJOzrF/kFIZ
Av+H8LRrUv8MWSpJTjwZ+VGfMRZCSkY+VEGROpjKxPDk2Qp7WX137jz6qC44M2bd
aMyDEmab7HPyL/ntroy4h4gurDrl1Xf62KVZy6qs/Yv1O3AjLzCLQ4Rv3i//ooV7
c/0Ygarv1lUKyVjAAA+WfcEJ3y8S3fh6Jat6ieghGQ+h5V54nGp7P4qqogSr2ejt
sSHzGqdUlc0qA9vy9pPUPMihCvXeJccxQKjMcLSGbwwmLsc3f8PL5YY+TDCNW2SP
dW5dD3Cv59qGn+RgvVE3BLTaNIRHweBNUQ+KnIwiBXXbSY/GT8GQ+Z3aya6tec89
pYclupjxckQHUyajKg2wQ0VrNynY1WDzmDREqGUd8yC6h8cM8B/laQ++mxkeSNhK
2/vGRInhKSzwCj3FjXCsR5LtqzewUYeCYX6Cu+cDa9OzBE80INQF/QtI0amgXlTS
NN1ltGSdC9fqMzpe0KfnTkvCABuo0aMxpxbZSGIPiwWQLNXcP/uIdWWA9YLG7QfO
bvuIk+wVevMAlij3uvoFZd0R9vKgrPaZyNyU85WGZt6HJKpv6/c6A25BnHDVKHF8
5dC4jrV+u6SWw2yaKCT5Z53TIIL1c+fP5NnGXiutRNluKlyRh8EyzUaiocARMD10
+HSSADRWCp2T3lgLrJ71E6HTdDCao0llyBmvpY9BM7WU7xduLV2HjAb69CCUIpbp
r8RIYkjxqns9nJxQTgWlt5EXKktzbO2Cu5J7dDoI2YuL2O9a8XMciTQu39z3pPe+
GqBsZrr8RrywpxpUuNuH32+5C4vwr96ul+46hWyo6eUTQpovKpsIOY7p5OD4AYcX
BoHFk7QjWVVdaI0gc0RBWePIE/7geTkHnf6izUQTBafdw8+Ldo7qtUSMxNKl/uin
vAfS4VijlntLS26vUWczTMcuqolMYHtsyKyS5ELCMAB0wtyLH5J0CqMNUXvFxWAZ
Fk8MPT+MnOMNXDwVQnBPvrxaP9LqWUZQCdT4gdJd68BETYpAFcmsgSAsJJSod0Ho
lw2Oi6Ww40OE4kKnN0MmTuqtKlEc3tjpg3lhjLJdRleUK/xvxgy4ZbdcGFK32p9M
DXgwg8fg1JjDgwVgBKT3RcOl1uqsBUAqv6p2gh8HToJMJ7AsCYYgTDJmJnIMPxo3
I1Tc0Kz4ru1uFx9xe40pppD0qQbMwbuzpYY66RR7QvlUojS1MXrJXsHCZ/qADAKO
DZlQFRX8MffXkCBwBKgoTo3mf+WqMmc0EZbcA3G2k5oZ098U9ryUhhmdyEq4hIDP
5GvVFoiP26TNfkx10ZzJ4PmnmUv8yJ1KpZUWisHp9PIShIbdFp+Sjk7fWC954N3K
yXGY84am/cUM5wZ1nqbBkvmSfy2oqYNE/H6hY7gSlspBpwNGjFFl0B2MrFDGxvQP
qNyboVlWEUair6Y3zIfwX8Y81wvE0jo/yZWrcZRU6SnesHx45l7pj9dYCMx5y+aM
43jtbBoLae0eXjB2lorYp4ZZsfroHDUnHwvuojOCN2+w5xJ1OiEISW1nnzh9+lSO
RlMb5PwUTn0w+LR26LFg3EE5mwzRl/pcPVeNpX2JKXVNo7XVOiHZnFe+6qN01hnV
OGFtZEGuK9+ydRLAWBQ/gK8YGgVGukw8xsKc7TC4FgJP+3IP1YMQTh1H6q1ilxLU
x9lduRSqwDiNDuyySOhmLoOTKvVF3LwmP+negxrwbIFyvNASD7a4Y10GlJiocU0k
QvAG2Fha82corIPjt6QuGJj0203+cRT0ashgnKSKvlRSZ/LYwEgpISEWwF2MwpGY
r2FQgzG9GULuCuiJaIkeEjHVstaazo77Hlcen2cikDYki0Wlh6E0YQqcnXDcCyzc
fhEVUAcdl8iH8bOrAyx3HsyEvk71Fv75t31GHPvQhwhaf7mWQZrAYrxbWzac6NVU
ML86hxV2Q1d0UBpUa+Ib06eH9KkF8FfpmpOLwmZ+Ffo+G7p1NgVd17FGXDypqzmx
YNAaTut2pc5PPIHYbYARQiVzNbX7QiUyE2BVBtbS9JBzLNWC3Z2uFgN6eBetP2/O
iHUfSUhTjW2rT7FC5pZZqLm3sMvWK2UG+z4zhppZb5aRddu5kkmlhihlUP+f9jEq
MzOBCe8sinDinucoLDgg3p/vKZzNK2ayHPzu2GzVuNy/juQchQtqaWB5NdIJgM5s
hrg+cq9+B1UsDtwfohJpIKHuFrB9rwKf1kM9pj76B/lJXq2ePagmIkD9C8BA38dN
SVuQM2M0Vez6IpQ+z28xUwGeAfnOvjBEFBptOc/8YhCpO00qoLAKYmMpp2Tkd0rZ
/hfyPd8Kg8VMRP9ZfmOh8l+slMaulVohrh434F5eeup2Dltfo5aHU/ygjr7HopfK
4T75CgPy6wA9gKNl3qZnJMQJ7GAvh/7DtI8ZZpjDn4DgytOxo+BaVhANgVTnEezw
9beCiGNh6bPOnwEOTUzB6VetMKJ8Gzc9mylVtE+z4QSGcDGzwzIv3pwZfjbwNlVB
SpuE7TqrJ0kZyT7jFqP5eXcIHzXhv1JBx7Lj6GbCyT7u+TyWxWTl5VKZVrf3CC9L
IUggRADHKoi6TvEmvDNABHTnVMskRksbVFUXEvZ5h2qBQyfakI97FwOlv8a0ij8h
H+YtAbi72SNctG28Ag4EgDR71S8FQshNao8fcqCSu4ZSQsChFVDtvzNCGSDfOQ5H
TWO2bWvRER/bKJ1GAJKhmjbeIYLvmHqK0dQZ9mqVAUSzr3Jl4Gnb2ZkPkNNZZkon
RmJJXlWoDBQzpdoNTfkHdLOE4GgrHGQXWF3/ucj0nFacNHMGZE95ds+OrM+Elzu1
6wPd4qOy2UEHm2jlrhx0dBdfEcjoxUFFKN2u7QF36o/dxNScmIrDrkcSFagkCIZC
Hv/7//ASGQ0XArP4mgrBWYL1KZ/X/bskIjCiCvawSDdgboM3DN/xRDFbiaxX5SwM
sswPl4V5xbZBSmH4b9IH1P8eFzJz/86X28I9rCV53L+ZwfWZk3iEqeHhoJKyEetz
MQzuNLODNTdrfFIeMuC/O4N7UDIl9Sck4tSgfziHsV7n1xM7CpO+Utw6NIfAWxh1
t2pRBDQD5uX/mk9u/AhtwNmz00gUDGc2NE2LvH/6r4qx3lTtMvKjxPsKcteuXuB/
BWVwJpT0iyva1vKE4HfO1/9IAm2IIDELIEFkHtH7Kv8UcPL+s0OPq37UcFAf/iKD
SQfuBjlcui/lB55zcmqKHfxP9qdPpGV51V9NnFYNaQHuIHWCE4vlwyAa1eydCfSf
ZpdfQBt2AiK2hhWYTUhFiMllLPGcWFiMR5mKb4sH6thaijA2QCZJlCkxHK+VJABg
13JuJhfJSKPyCkYgQUXF3cSlVQi43av8j+FmVJ62W2VYPQHiarlQvaf1X9I8Twbs
aGrSJqopRlvmG4dW9MkvlKJNmtPoOmgFczt0GJJdP5u8IYkvGNEO77I6RxxquEfb
5AtZmOYnpvO5Y/atr2ZTxcYcKGMpWNKTYwCWNA4PbB+tEaiq/nbJ6GGs6Riarat4
hLFboETcTftzYJiEWa1QubqrDEwpF5v3r3CD1o926m18n9hKWKJhZl4H0sDMxEkm
Kmq7CiXwNdizXBJef7xRGCTiPgTJJ8wdABqbbhEDId8hbh1mCoWq5o9VmI1T7CwG
ip97/WPWw3lPhgd7WxBozhAjRulyoyAgOIv7ustGKFfXBd7fmPKSeXTCzepF2ZGQ
HGUK7apXTgWLJxTqr2CR8rG9Z5PTcAWdEnK73EVlZGKgU+tPJhozlc2FdBFQpBj7
K943izCp01gXQiCDUSIjNkPugsGggPkqWcyBStdnquECWHaczjQxw+u3UmRU2r3e
h/dUjXQkYY0+1t53S2ItwxCDOZrQ2vxxkC0UujkcKPow5RQjTIsN2Rl/ll3sMLPl
TVS/7MEl4vh1rwP57bp4WcglW2Ftr41swCNwiKIy2fK1KAxSaPNe3oRZrWBdiIfs
9o+mXA7iN68U2PBmHnrSpHYdKttjf8lCiR34xRZr9IPcAGeVvVF2mWpDRphueJAt
DQhAvrpKUZYCDfXIpAcdeeKHrveb+SkK2/qfqncaeCXk48uPoYX1onSVF8RGn5ze
oXNd7EkvQ+3mF1DiezptXk03ecBwq9qIxvF4O72hGS9idKgWSPEEBnoRJol7qiZV
IQe44eDmQ3W1Q5YuYJGeu2nA7fZk2COp5V54gmWQ5PskyMjCNCh+W2ZR89ogSQC6
/3EGG+mnj3fVT2TfbFGFNXPN4abLAtOhX+2Ruu2Teue1+awgeRB/Kvf2gSqIj3XK
FnefyCZ8Lcm3XoUfhwBYKaa2ldiiCh6p23aNvzrUxeyvfGCmkyZbJkfwd1ebZz7T
5ebWOHh67q8f01lCes7OGTYICBu+xezZzukQ5gtEZSn66uc8ax+aLg0m3SCo+usm
biWgMh/4Xn9wNBXHE99c6KI55knhzpkNnh0Do37BUqtVsdE5o1qwN6Iu+n+auZ85
TUyMd2Icq1UpZNptcnsF37AfmLHHvneDY0nxRPyGkTrxRMQjXRlYPA9Ag28JJ1DU
A6TW8QFte4k1QwWTmxY4OGjUENKmzUDInusfrKIhKJF1SHAPHjHiztVhK/lvwCi6
Zt+LtY/iASBbi40lvod71A5yqm6PwmWe5dGmAhDLvMOqyqmUSH93aI+cv05ez0e/
fz6alS6OCHKm+v1GX/5jG73EtWfkAPeOfYtRBVyWS1kb1Vycl/eEWXnKWWn68DnU
ZZlInPH6WGNk+NUZwcEyQpzPDMHOQj4D5hDr0DbDZZ11meTTnJkSKcXUwLs58r9a
DPES6wXxy6VAyMtrwgZqWLnRWy9S9HawuJQDgM2Fu5GhVdIIN4c/J4M/yKairg9F
yOPAz+2NOwNpdqYgczNQU8kNdQeSsTnsibY192OOMf0lEfB87Uqq36CuD8vW80PM
CH6yorTkqZ3XVkneR1vVK3NM86FHcE/Pqf2C98uA6QGf0kzOW6Hkx6pWhhvo6nVr
3BpvoPdVcu3LZRL8jqfyJaUHNVE66yxGFnNzXET/8iQG78M7x+5hj3PG3XgYkfJu
MW+qXqCdCxTmg/nYLNKAXS3BroCWuFWRksbUF5+iv6vFatA5VSLRvdvYTCANeokB
z/6ug7I1QZh+6IpFPcqVjtk4BKCrotKEDra3NBgmdU844wYVKb9lnmfCiM2dGrqN
6/+dbMohWbhbZs0xu93TCxNU+iO0Hg2NXePBAcYhJQ6mtF2n7V3bbXPw+jMy/yWS
Z9imqGhDGIVMZRY9uB3rbst357/DpDwVjIADZdRW8+udHZjbn+Qjg50Sjd/P7hu8
07I/ERduD5wClwU+EVXOuw/I7dbA8ig5FIQvT/vQjOlLNo7lC2iCbpxyih6S4XP0
v9qtPA0vf8TEgo2NxxOXtgGEOcsTn5pBA/hC7aJhjFWzfuLjBOzpEV1pLrzGrbLN
yyhWmFt0ci7l345MFPfYLTYN+5EZM3EzuAURrnx2vk/FX+0EXLpZw9Phgpjc7HNu
zMkgfFKbVA8rOoCSUxQpl9UFPL2WeT60O4TvmAwu+7Xk5NEShw53QjFSYA2Aga5m
7fO/9LprG4DQonv83WTbkjBD9/jDoSp1PKj1S4kPRY56KRCoGF57kcrPjBiyJFlE
yrV4imSyBTIDpzMXOiXxFqv4WM3lOkfjsxHNB1WRnjh9k98wncrCD60/Jr00m/9L
zKfqKE/jgEle6z+fJJLBck87Ed9hkuTkCCZfKYrAPQNBf3ITRj3rCgjyv8crmxwQ
/0SlXioTjIrefW6WeaYL5Fi/w4l5/kcETtTdZI6wLHhFGKk71v/7DVGToCHdQ6UD
3mVQKvTzSnbxiz3EjcnlYtNOiipx6PhqVrAj8MOqlNdSQ/r4sTN3c3yhoXoz3Lec
2VqP7iJi2AaGNzqVPIbnxf2pFoLhGRDlVHfaK7NLoOI1PBYklVSPyGQSLy6BxhZt
Fb/sOi0RVH8E7mQZka7SUaMmom0HL1sBBLKMm6pSrb/CW3Ez0snBK7ngeQ1xAHBf
oGDoZTj/qn/nlgIu+iJ5uaXocekirAHpL8cg4DPoLOaOqdk/ov6DRdITuSjbogY7
kpovw/VASaQ74aK3BKEtm/i4PJK2zozrcr8/lIrvO09q8LT4tOYZU5uEDxDf+ZLg
kuJmVtNDykEXyym0IgYH4uhdRbomyrYbC52ZK6/m4WjohWHBwvoXmXpIcdSLkKxF
QmCpm7JMlf56muw6B+QhtZsK5pejXMDVTMSWaSwaoa17RSJ6D8qCs5kHODGcyezu
FTbg24aktq2qkAYigfJ4oUqhlnFvKuw3QxwRhGHmmZizSiyu5bgjODJnpeSKLHmg
40XceUXHRqOKpGlV2gw9w0+6+FQGJmBN/oPNjzeIBYJl3RiRSABMCNEabh/Vt2a7
C9DgAee21z3cKyl1PH8jzXzq+B7NrgvzV16aiZue42bcC5yesowFpZd7lsZOY9KS
QKg1HSbzzvUP9kznSBRAsRfHoWmffHIRoHLWx+WhVwultZPkRlrBTn4mZuwKVg6C
LW5lV9GS4EjBN4+0stMIs/Bir86RbVVIAmUU1g6NUAo0Tt49scvkAX10aZhVnXBv
svuEy9ucyIext2E5vr6ZXqKvUHy6HX4yt6KDlP1biHOnMvYpBe+1rs9Pg/AimPIo
rH3Q8WtmTMmA6mzNeQbAX1iV7RuVZShJYirRFo9d8c9b2d+9ti5PETU1/+0DVfE4
/nlkvUpPItcYuvJ+YCK9wKH6DzyPTA1V97O4pxS8eHDmd8nnNFcQlI/DiWFI7GfB
VTBVsSS+7P5HmkaV5oUY7KwKAQDinzSnQZbik6SPVkvpQoy9p0fOSciM9VmVMIcV
0hAGDB+nf/JsUKUoh27Z2frCm6nGEZG67tkUoyvva8GlquqCMbKpTjepIedWZ7ST
rkjuyw/ZDI9bwiWtJ4+Bv+RxO138EU1QCd3SZGyh1uUQmBRGnqdCqwCKnF8KTo9S
P3qO5YCKGNh9JNMVChvzNbX2JrefdqOeTozBtLwz1vbPyqmfHADetUzsxaJJuSTi
ywDLXzu1klXTQ3RXHUj0Qf/CQ6Z52DvWqkumMMjZfmO/pX7imxpdZch5VhvbfVhp
8CqVdgTz+mPyJmkCVHBLIMTVP+25nLpX8EXt1U1KNFmUpbx06wZp1fkO9MTrST/5
VtBNp0kxDx9llPDTJgEHjoCwLzJ83tNQ4XHpOGCAAu1MKpJrP7lZbU+bbZAawzH/
aLaPWnyjMQWxGqTJ1BvQGg7Xx6JMef2tC3wPTatx6oMNgIbKv7w+XVoADtUUHKDP
xbk8lKx6x5tAKdbr/52FXcPAWOVqV91QReWs+P3oLkyEcsmieThouH5cdzbhHEBt
tAy75QEorqqsZWHuCck0/UqJmxdxAZ0oB5u4NDkfy4Wx0U7Wj1RLbsnh4W8UZtPh
CHxeBHLvAIGKIdDRxXZ4Im0+TIv7jjUpOo1Oqc3Lrse5BWDhiCshRxo12MUFclO/
wi0iUPbeACksjYXDJ0Ph8q24Q/+BTYUjzUiZ7afqDV7p8umPmzqKvAWERwJboLAz
CUY/Vb4L4GRrGXDNRaLUUZRWiyYek39CvriCNDhjB/Y0RqFARCuCD4xOg4LSIbgJ
ZpKzBW8xDtBCxWwRAYMO+SjjZTr4BfyGhtsXtsgz8Go65pTE1LwIJRhXwR+yWqWZ
DTRt8ZBizeNF455CNtAJA4F0TPikt9gK5fDazFibgcwk+8bE3ol+rOck45SJL+x6
CmbrnCoDj8w2ASEX0/W7NVf6dhm7uE8wJfJ9TeiftDgfGohuI3BjG50PDR3CMilX
dhSpmKzT/Ek0DfE1wCXgihJpRTnA3DUKT7vU7cpruwsn+FEgYfekvJ8U55Y507dv
tAo4fCqIFL8DlUQA22kXxno+9OBKUrnGKgmRoBgIoCtIdtUUy8w14HC29U6GwNDP
DoHOZKMQkwMMxFE3a2Yr+R/ehu8EZot+dYx5Rl1p0CzwBLD83Hoj1ss77zoImILb
oI/SkrlKeGfkq62aPJqhW2RbSpLOh4BWfghH6aWM2sFZ+DtKYJ7Sf8V2zkRuV9M1
oMcfWKACfed37XJ94ITRPrOhQfb7kh89Oxdspj3d65mKI+wjJPynvIam5LNDesiY
hWlet3ZKh+SxEFTLP9KElDhvOoyqlWLfta2BzX8f8g5srEPw7lZ/eVGJcRQUxBid
ce/arTstZteCc+C9pChUo5mshLfMjKueUnBUwfhGb9KbJTCxppZcpXw/Xbr5Dofc
g09X/PBoWP9qY1qG9RHoCgnyRbqsbNMQbOuLXnT49hC4NuP3va4m7T82YvKY9s1V
T+1ZV/UpjgUHqU6qbniimtf+iMWrd2KiJihuz4HN5pr2iwKJ2rW9jvxO9qnQHNsb
v9033f0BhTDETI/NTzqD4+QtT/2JYA0BB+nbmrNQWsPze1tW1ECdJ9PlwzcxCnEC
jgr2tUkJfVDXSm+LY+G++vsUA6Lc2KKutjGDxhHIDRGWvZr2Ae6En28PbG0XYCxV
EPwlkMl8Zvb0PIp2N8Zn2SmcJ5kSLhZ6C7XMP8Uo93BOxEBno+qoKZzNMVYzD6QF
kweLAehMMETjljyob2Chzd2+JKwzVMrZxly+0NZZ/i9iLvvgcoUNZJw1hx6+kMs8
DrB5NWI1KpYrprgjw89fJYAbecljdQWb8oCXXbEQU7AOUPknjrVE23ldDYtMvHX+
FX3g+TXtbIuPsxWh7DIhELNdjVr70U7xGUk8sQyk6y8jtHqZHOYHP75eyXyLUyCM
nkMO3tpmw48FLeIFAWattO6oFtzKf4vKbdm3qlj5CZ9rp0ozR3WYpUiG+7Zi2xq3
snggQGHveGCM0w8u5cWeTq2zdX3TAxUVWsJpS7vFj0mvGdNRWFzR+kVLWv/Y3wzQ
61HqK4v6IbN9wBWEUXaA25sq1/lenr3PP3YXlkbdpwERoS5riDz4mqdGhO0AkWPN
321DzL5S7PpwTutInDTMaOtFbJVyLgk+aPm5QdGEPcD90dVmj5KPVGmb8KmvoN7x
+gT+JksEGKcmKUbxfyOjninR9taDEvf9lzvbhjK9RTjWVMgIWC2tSEgvServiNIF
fF/MvBp9UzkbfWIPYwTa76F7b3KgQtwJXMDE2sXMwlpRge4mA5wkaot/9fAGydIZ
zs1/+rkSp6lgM1Bm+XthFRYNSbwEb16max/kz8Xo7MFdHSQIYa5B395iZdeG33eu
RNXbEGmz3YUsxtdTkx094Oik+tmNBSwH7/lV+52sbC2D8+L1oJ9UV6KZ2FfRXjHi
uwMiF3EyNpqpBKJ7ZTTnzC2cIRzniQBeSovDwOo7Nyob6EWibKDw3kcKiMDFA7zg
hgaT2OlbHYtcdTGGak5BltzOhCLUz0+mVP0zAyomHgIMtJzGmQdUZi4SgHNj1I39
zEFN1UIqub1tXx+7FdTBqvkJOWwAZHtKn4H42s5mndRLUfxqoOb6br6XZebSmPGF
aZgxNHt3xIHuQConcM3ZQeUBQOo8XCCUfVvRvQu+ixUo27laokFeUUqkLEIcMZ9c
5iHmjNFcURFlJlGArhsKHoF3pdvOy5yfNUQcjw15K5WxToSyeHpK53YWL6w/XV9Z
adBGdos7WedNMu3xBIBfc2oQVbYSXkmfViGqQ4F3RNpVia10hXT6dCwXavv/Pq6V
RDANNVJrHZguR0RgCK3G52UYLx0AMAlJCTQbgdm+K3age9FYWyhtD1bYPVA+A+Fy
skYHvMCPwJeZ/JpRzrsobjY0sEoB2RmoJ5WDi74487rgtA8FHo0Ngcgf+FTqysnG
KdJorScXBhT51Q8nWHJCySIkHy42IpzP3CHRmMPqiDKzGNVZM5XWw8gXsOVmumww
Va+/4/T7BnzZc9EoVGGqSdfW+Em9A0/XSDqObYOX1lw2XzN5FPIDRsBSRfcwvR03
aSffjWGHNGZ9qstNiNLt394w1OsAE2K25C7PHCHBxOH3pzdQHtKnlFvj+bspw7dQ
9QOXzUWd2iIIXDR33mFOxJEbxoTMm7+X9gj5979s/7dZ1Az8KR6nVfLRv8pStldt
aWARRZWtD6dAp6nMyEt/Patqyz6hg8j1xFRsrAcIVhE/sODIJmO/hG44J/tjClBi
OqDHqnLj9yDYA7/LQaRf+2SBdxbwvA5RxLK4UMLS/0PKhwKraMuFRGpXT9XGMcWH
N515lBNFYherbtd6yrZ3qJV/E7OO6YlyeC5/bUb/DYPz/hv6be13K4v1DRWTaFNV
TWigFaCCQiZytT3fJw36ZSmLU3N3YC9RFsiRereosqopc4jNH6d5Qbc+lcDfNUF7
gh2JvYMrMJscNUAAnC9M8RuPrmzo1hAybG1y86/FRCqBKDHGQ5lOhkZRw20n8OR2
SYCrFWEmwsqI36wXqEjp7io3YBKhTu4z2uQ6o2Mr63kC9rcqo2kmkaPOvs4+i5w7
zxPM6xevLtIQrCi3aQRwJU2gV+AkWYYimmdeunU3hSdWIpSqX02hUccGuLIjKrUr
VZgmuYphYc2sejiHyZeUCyPZjInIwxvSb+9bg7zM/Au6N9F3ZY2rXpk08DXDK1GA
1SiPjdifZHePYYGrawnI8NO9vqhZPs/n3a8ISSm3nK63ha2ugnqs1kMWpthoukNI
QU3c0wjXLaIYReEaS1Zodg9bFahsOhqFz6L/rIGB5DEd46i3kZA+7AkKp/lYhPiZ
zrltrtaATWGZ8NXh2AzVJonHmuZ1KJfVi+ZMqFC0P/AnW3QmbMC6dGVgkr4tt2fF
QPwNGEnFsPvWZLuQFDyZiWZbvnHZQYLXe//HXtodY/vucAjscPb/nCmjQjoEHgLJ
GUr+O7lfERtrPE5U2F+LTB1A8z/NRf7MP+XdrLzHgrXKBvJf8mzE8R/+3eMPi8wt
9L3O3PLtS0RtkZHBAcuk2Br6F1Ig+ojoxVhmyeSO1dKtyjYNLPSuSajyL+0otw3V
H4tFdoCLvIOQKJKnS9Hw9gZ1Lzmf+qT+muoxC42lUy0ezMKEpny/EE15lfajQ5hl
oo9EWuae5m0Y+iJfZ5q2VkpRPgoeswhDin5kDbOvuQYnplClqq0dMH12xc2gg/Yo
KieqrNz+gXqP92QwDPpN2hLgWTp89XT+c3cmTuJpq4uRpybZhVfZLRkuemCQhglR
YbIqKdHPi4hJ+7FU+xXyJ7AvLdV6uEaDR8EneXfNACQmDRjtu7OEbqPm0LEbLJBA
ICsqNK2B6GNGp/67RtYHJaN/W/0DlAcjOLYvZBH0WOJtBnJFsMPdpVD1iRQuInan
njYeSzfBcfJyxT4yZ88+RSEymYSTKvegDHckf7OE+RfZBCs0i5SwNyQ/bb2ZpQxc
iBnBmcRKy3IJw4NUZZyc5J9VC8rF1aj0OfYGKwkVe4NHvhQ55mkdo1fyIJ1bm1nf
TmrlbTR/94VhgBPCpXRJR+DtfhKwUHH2qaLBjrCu7og4oLIl6rC8OUY6KQZ68S1R
icM1Sm8uisO/8AjDpGfA14DU4S9imohtmNCto/54aMBOCvfcgXRxIzzAuipvcigj
S28G7BvBZI/0+Wsyq5DeQ8jX41iEwi0Ww8ubHAPnKX95qG2uMHZYkbpsFID6vNf/
7KHGIpbS6YBTe5HY8/KEwHIf5kVpW/S916IDRgOgTuqcF1mTpPVymAYZJBjt5qbj
YTBm2AXmiDjCho1poopo6+wIxU2rY0k46CtA0Q1++RDGgdDssxqpY7rShMsw4cjI
w6zsZS3AhNhsVWEoErDRozwsWWYGGdrdGVbDTzZPZvqjVwy1oikf7h7YrtOi1d46
Kty9UtU6cjFJzCB/F0WscyvxdXnMIurcqW6U8rKkT09eIJuLDDofkgvsbQq2rg9p
1v8gibbm8Fw/zPZ3FVg9TfxBcfi+/5J1U9yePuhZFVScUZbRuJlJIazDsL94H+33
Ta+i9XtBm4rScrPdOi+Xt0hZSZALKrCqpGyTsYJmB3fEtxv0p1QkL5aG1uSswzAR
Mj24A4Zl+HVM2oYEKRuJEu3g078jQHZxfiADtLR1uj2/9KuKStY6yZY3U9WYkwBt
yaqx48W0eJA6+KKpkI9sKJta14tdHIkiB25kdXttaU8r9RTqRArD0mwpFCzS+ZTg
nXzO0JeeCxb6wkBLxQZCU6d5kiA9ne3QSWc2db/zYKnYm2o2IiqmiGFFVF8kyLOp
Wi1EfKaOST000hI3jH6E+fUZIx60xr/lHmXtv78+TiGjSi/DYGjunFHqb7wSaoAq
m2Gn0rjDsQsGb/mPp2haTZr9ejpMxFboyUH7ouxEgA+vuZO/eWPQkmQDVFV+OIxm
QXhqgDRqYkVTiK8FzuVWpz/6iRbwln860140Uw2Z0xBS23IBJeSdcblCVSlEdAs8
EMfwu6k7xYpwXx5M55NjEzccZe/8qZ/oOgIT1doH8IPavhjWIMMm4fPnCIugKBMX
x9kNHO6CILSvaoKQzoLPhVq6w4gNl181PRCV70RQRAJ2QQYdNtmB5ymvNWFy9GQq
lj3Po5vm8kfXKFXtRj/cFCY3bcIBYhR7loXd553X38DN5wqy7kl4pwX3N4Tg1EDE
XHr7E5mQovl5HCiB2LdK5QdrByHobd86Hk/ihVS1FJwRcXhZsDbKEwtxtytD/6/2
O4yzHUCszFHKrDGRRgewwV70Tcd73edeNJ/pbxEXkUGTTw28GINEjK82qT0SXHdV
MkwG6REyFoUhCyhsR1LUYM+4irUKED6VpcN/W9QQO5Uxu1+BxoPyRzlaxONEQFdb
cVsVHwQIUwzlos3AhSIG46lnay+Tyb3BBgX9+8XGIn++VRseqSJfePozt53kxXi3
z60M4dgmjxOxpYTwR54+UK7tmYdQrNzE4wLS741rL8Qw2VoVf/0YXvG9k3TlUhQp
Cimhu8CErqRVOInXKPdkBIu/i9Rqsh91vb6Qd5WDtd9+EDeub7SBEKXn8ntGEhbd
VVdKLgSw3vHLIwoutmdwwNYK8Yj4Drpvp3fVwdV/2E53pxqjyvt1DTMR02WRe8m7
Qloj2UmgAuV86Fm0IvOkb0gDEnJx/Mc/orFATGTwdXkj70t/Dk2YUIl8/dasqMLB
vfgHzwG0EGo1dTz1KOtmciwkIG92IeJcwJfzbrJnrB6j6gcoCWbaxvJX+yGmIUIw
GWI9qjytb4c0cI1i0AoZ35dqxMdavqtLGun5INZXeIPDs2ALe5/SXDbAoJNVC/WG
uU16rI75cr/F20bCJSBZqY68D2N+9AWdbOB+5epBXcOT35KvOh7LghzHdjzXl3Lv
8pUpLHgTA76CYhoG/jHGPI82ctfTQu/z34Cx1lIItQ1W8C3aQ148YlAJLsrDOs8w
e+E1Z7Nu6wq2FH6AbtQHaKhh/fuibTpNIyatTAxM+n34JThx6jNf56g+BJCbpEmG
aY3NRn88FEExxo+mihz3Rlhi2MatnH794rckGIMLk+9l7CThEjW3QlCMhIB0bT07
2UjFa1hdXGXJ6U/a0IgLEPsN4dUsr8b2w7849i3kgzyswQiDQMC2TUp00rLauuPY
UFpxndhU1jkPBEijWG6eLqcJLxlxL6p5T1Sw2YnoeZ691RsbHkAC8sHkUi+smwcJ
8EiSFZjsSemjGZUzwVRm91AckX3zMHZfz4og/wIZXaoZPl3neS+93El8PEuH8SyJ
lRGqRFhPuL0n+nhCYXLytQlDsz7wP3f4GKX2DvMacc4X1e8mf0atjdkQ3m+fK44/
IhzSqv82MBiBor0g0+ynbvruxMKKDTAbtZBuUVkEcvWcJEa7YQ0fNihnFcgYgKKI
bPe4vzojkAQ4qmtZHcu9ztG7in5vqC1FL3d9O3NyWvxG7TT9JUHF0fJtbmd1+I2w
ZlnFJ3c21J9Uja8EJ5kkbHTgp3eOYaE+TZSHzTHJDqg9gaGEOoj/j0MDvY6lv2/8
mSgtHveQvC9hs3FUBCKRlyVN2Mq6feET50YoX5KE+QssFaMKHJAkNkDwiTHcyUG6
e7mdzajxGIxPZ1ePZ5GJBrRdcwrvp+DlOTjW0W3wL6aXsrCb4/YgBnUNBuc8m9W6
u/BXJ+Wn5/uO3fWw9A5/I04D7qM0PVUpjut1GnGrkXTYqw8X3qyFmH5UwfT0Nin4
+ceA0nKUiVWWfZq9lcNyzZORRqS0hcLUgYZZXF3BBLj/OfiTJ8qMI/tBmPYbKr7Z
VY71LH3fqoTIt6o9/pujQ6GHWkfph3JHgx8EwsBaIQlejociPg4eFbShKz2J+Jci
i6b7hIJOlf3QIZ66HowBJ6wmfNAUsQUpe4kKfWbyPSRPvyLEC/v+jtqAmyBnRDF2
rSjqOoeLTdYWjh5pMIXSmu/3TTuUunLaO5mKYUjEL9KJ04cYUVygJCZqlyrvQeMo
DNkg6q0OiFXqlcYdBO4yK6oJZy3p5uMgtp7cxsS99eXvVJ0scgzQHQjJ0Dm6OFtI
sAjxX4xTHDr5wTFl6NkPF+pdsOfAjfymdWmLpRGm3KFl0A6YMdjGaEWoSx3I2nHj
v6wF//oEjIp1l6jtzvBjYpm/zPtEIm+FMesM39m5D4SIw22dOo7Uto7gxvHkOrMe
cmTpDa11A0RJt0eJIiUkHXSLie/aHd+7jxQ/tN5LnJ8kOHTzAFbrEA6T4uV+K+2s
vDnenJqr9Czkm5c/rhtKoVoyQbR+NAcWtqJUVxARWvPJBeq4QHJAgVyAk8teUeXi
CA0y4pXvtc5JHoWDAKhr4/qPpDRDwGRGtXHqbdUBwvtOrrjxHTGCoWWrXy3EZtad
g5sfMoZacq1HGAVlV1HDm/XtWP8CFHuHAJQWDYVLSKTTz8/QILGZgB7qdHyfACdh
Ubv1+l1/v0DajmUx3UI+z+LnzspnEhsDHmViXMdATJbJXyfbeGPfxsaQMU0SKwCI
C6CaXeNHXa2rMNhgj4ht42V4zktaTFIps5BY3NqWpYVOSh+AUhygIvHTMa5iIfj8
KCrQQvgLLoUzBLecMsHQ0Hmp7XJwCCpm3fBwqAN5YqSp5u0wwCNQmevDbgOHabSQ
zIlRkf2wP9CzMTVEs4IRFEvx7hAkUM8s7TE9Ihy1Gv4kWGIpWldPJrmSwSHCsS3K
yMKlhV005My/PTOxa56oOR+SN5GvywAz0lb+OEWt6L8XW+7B8AKqECJbnJ6c/qXd
v+/FW6YONNtlIZPUZAciykRdQ1eiICc/JeimiCHyaZrxsvE0gxk49gheQLJ9IpgQ
CPqtr0SPG9+ab7MQYDSAk3UbXTMp1mKmc5TV8A4qyJV3mBkmJlI+LEq7tNTsxKfj
JTe9AzwAJ9lVKq/rlAwHTHu3yHQWeXPSrZ3BE45998D4BS4L4yO7dDYAYT84Fh/O
TxUBEw9zDes7gxkzEYjojgsbYTyROvqlz9d2XrU/ZNI7M4AvupfjZEGF0Sfqo7G7
r96WuUxrJjirNlmJxksiJlhAtiKd/VxYp6ELW0po9RYX9+c3DoDqYkzGUW6r54xL
4VPoliuGdUMyNK3TjfqSqoCOaY+EhQQ7nJ7n5fktwVVU7mXo+XazsmNK0VNPHOWW
4AqlsnMATopYebwahAFxxmaT/d49dJjkgFoATMWuzipJofO+Gzb+8k4hMthsscdH
1LOv180sGh5gm9VUR0pz6ND8n1r8qIGiy0t8x9OnhqH9NJJ3iI0BWJC0HTTExbCB
3iZM+3oHCn9HR9wh/MD434xZMBpymyNhDy6ml+LqqndMeFYmfMvWGz74EuUlgGT0
WrsYe1PItKkrckHb5u1V9qu9DyKj4zvOyI8wN6UbcczF3DJIl8CBeo3qMfvd6ma4
nBFxaIyEDaDP1JDuKBCtsoJsNJ88AWUiIg7FfXjsY3ymq7YsseLVrqWroTCywtnc
6EA+oLRTWeL8S+GmatnW0xJFXeJuTdp3kWk9MuoTLNZGDh6UuT40TL/lpzxj++F9
D2892nhixD0QHYQMWS4qxynC8d4Wt95gbOT3o3G52Lr/W9tQCxfh6DcevaNBa/db
riF2CWIAqnqJT8QDKPM3dB8YHYRnYtRsUUo1dcfvZRnS1aKN0cfpk+fBCqd19bKY
XzRfPDgTgMkNAl6OKpuYbotNdxcgSDmRCXBaqnPfqkswoRs+c6oWF4JWHArR3c1X
JavDrvrkz8mQkX1Le0dijuDy4gRN8gpkOH8dI1VPPF8QWbVDVmMQVWVF9oB0am6s
rBFnF2n1tlc637iG8/4yNqWRFVf2owQGAdZ47yp2EmkIQFfU3bWgRMd4KkGQTIM+
dBezojHrH6J/pk8aKJkOOygVMPabhS7yGGpiNKaEB3l0d7BAl4J8+BUOENE7tiQ7
YLCvB3lVl5JrzgHOUUJ9s1VkCsiOpReDBD2IWIL07hZBt1JoYoN/pdGi/jY+GQRx
3sFoJQrCdYQJ60X8bqjuszA6D97IVcJUyOTrmeYg4RsHQTH4hU/EnMCBxuNu7Gaz
hHXVdXvO13bwFLtqxs0OnWFnCNXiBMXCwwb5YwqwiM+7Ib0hSMcpeqaSJd0us5Yf
j+N0DKioK4WJxAnags7l3Pj4fc80KbqOmC9XUpzUrfCCSIKRtHsC4chtPckXnFbe
tBZ4xiFFeKRbdKfm/L2dm/yeL5DyygOHAfkdERgvHqFYQSkMYcjRTH/Mtcr/Lalg
ExcCUXWbgJ51PYmMs0Q+s72IoWgnl8tQtAWIzuy9tKp7iE+hstZNiNxFkizonDoi
2F7VTbGBxlJ8xKNolntRf8N6nBlXzTa2gshuGFkb63eoe+/PxfbDlcm4PDE1+Uuv
8zEC7DxJS5cyiKm00yyQC7l2E4IInKxEjZEjX9BiD5r5BJoACmSN0vBkaMyk0/fX
3IqA/UmsVYvELXbSf/5cudKWbycNNCU3SOgzJmFlYEQzr1OshhxA08KhXdl2CECL
rYRlqLM7yURtdJ047NLbIslQZWcsWYBMli3lfFjNg+D05TrrFeXe4Q1lnXaygZvw
JTLvs4mWaIQexrL1gT/rUHsckibQ9nLINWAWDqmI/BtKxGmwWypJbqSTuRkatEtO
Ddg+ktXfZvwvb7iDOCTqQshXhCk1ALdE1AYlin/uLPV7kinuEfpep0V6FJGh+NO+
sI8yvSNj6b8Jop8UzY9SpkSqZ/wj0ANR85E2715j7+rBTwuIVHBfT5XzR26xJL+U
QalE5fWO/PoUE08FfzDsWq4/fuwW+OVwnyqPc/avtuHNNQytaxtz+fo/Uh/Xzcmp
YtoBugcmJkSW6K3uP91LvoLtjR0TfW8DKRvlBhdt1vckcbsoDldTp/98EfIe/BWM
qhv+GEU98GgLuNepv8afnhJssJk7qC3KOWn2x38mH/XgDba6oWAvZQb9uXT3Asti
Q7LIU51Db/AC1sMS3dNg86Pm+vI7t4DOCgYnDpSZZpLa8doi8M8b/NnHiHDbDclx
Wv6R2yVSahwhrBESoPtg0t8BN6XFcZePL1hHbHzgDH0XNPilJ+pjFe+WGqINlxPf
RrfWW/jLafkd++LZ+DfZzkOf9MO3OEZVvgAyjKAAOiSNL5qDRy+I3qDx24ZI/YRK
lA57et/giBs6xQCmpANYcHbTbzvRGPpOQ3lWvUsE+uuKH6MFmMwurz7TNeice/cd
7/3z4K8VaUb3UfS2gTgocTWlZdflKEaMtAO+SLqDhItHWhZbczmXXTgFWfHnsRr4
I5ANqd/tslc5gzsmp/ZFyxfWpoN3HOf3xD6sCHTAPDdDUZm4iw6kDMeajCVSUVF2
IBSA1OaAiwTQV2+2sR7A5Vc3Z+p0HurnlcusZEotyOh3ffmwC8J2LNw6QtheU+R/
+1Wkz5M0caKsvRZU9r0YBQMZCuzjAVUcfZ2qpOOxFGwGmqW2UJD/e+eASF6R8bZJ
V8xGMp/ziRCmqtVLwMJoGcuThFgap/USbGs1recLNqe3BxXvA+IHxHINtG+OBX+9
t9e9UMlk8HYLDJ0xp+LZifXxKaBRGyUessyhdr7fvSu7Aw4deM4cTIh0cuBNMuRA
iNVNXpxQoT2fhuA2BI4m/VSNealUvSH6Jx+lvQfgmUuHbcQxcWE0tntAEFit+jDV
5yAtUrYdxaHw8n1aIZJK2TkA/A04QWxqF0BZ2ZVf5P/mBUEKwULVd4E3TuZQYjJO
L7MmPkkI4VtVLlZMT+uPaXdRe/Ak2NQBiBFadp4RXBXx3/MXYx9VpXT+M8nZ9hYN
Vujhe/hi926aclh//1S8bLl+A79uJ7xF3p6CHyhOyr30yc/wjW6nVl+8rS/p/MRT
WSs3vASkih6gvObQwaqYGnI4kIUrBHhhUy9AUPXLmgTJda7M+rfm8iCwrKMfzdOB
F9euLYztWeth8f54T54lH1DhHxBA/5GXybmxRBB0N1Tuk7JYQzdlFKme8FnJA0Dy
lBNSQ7tb7NZj/AOUyq7/bDfyQpZAAstVnePEQinbVbsEY7G/jZe5bzTSG7ZdidBt
E3H6/fQbRyEXS6rof5AkDdcEVfz+ZK4qMnr9ATYlEjoD7+Cms2D3eeTnRGhlxak8
m4hfu8Y0tSCw91RCcvnHZoQJui/VZ2tgaizrOmd7ETWmh9eaMiOXf8HxvJ94uyHM
LKcNK46LwI1vuWI5qkhhx2PuW/6EjZsmwKZjYh3RkYMXdtfb2/QN3UdauEu3WIpd
idlBhLvc5msCGhB2KwAwx7580APSIYdEdYGl9Dj7nUzaa2Bn0jWqTzczVvSC5QQV
wSAh1xY1bS3zXGIwrVjEHiqfcMy9oTGmNkohULcoHMxTQ6sYrW3VShC90TJqNT+r
+AN9h0Z3X2KK1jACN0Ux0FZgIMdfjSpKz9SH5CB3b1SNcWqXuqYb61DQP7lbn/KR
PBxJcdTbS8ZC+K9uK2SLMgFZwPteu8RqSM3nX5IhmoYno1F8PvAZfOAFmjj//LMj
4MJGxDv/0pw5KkJh4ZypoFXiTuJijiFXbJ2QSBnoCxONZmwEp/2sSo59zkJAeaVe
GcX0IPmERcQ0XEPwJXEgPSBQrvo5TnvZVoFDe9gbUngY+pLwE+hLgVlFIllT0KaQ
tg3UhkUmRAZ19nu6iman2PR5xhAHYBN2Cot8iGMYzjSXa8BXYpxb3lzzttnJ1tcD
dV+tjG9BpsU7nnyVM2f2rRtlhN0iNTOFrynAxjd7t8aSafDVW5jqwnyp7dQu3sTP
wsA41jrb6pdYdWs16Oqds0+4ClLvNXyegql6zfnITQzhTitEM+lZRCcH/1bww2DY
NI8jXVdbbfUby8P/9r9O7KOjeWPX1kg/ha5gNV4H4WQyLtqlBr88FspCXc815Vhb
H20vvluQYorvs7WZ6B5pousyTH6FWmWoRrFwNF4YMbymzBJnxXUpMtOtdHgEtfHd
lsKBfCUeHf5VrY7T3lK7+PWfNKCAcGH6X3MVnwfnZpzPBLUtB33uUcQjdwR6aqcJ
H1KuZxfTA78hoE5iuNKH0xr5LvhpM+G9qQEWkm357FhL/d4G1dGwMqF8uO8/2FUZ
1b0i413dfusE+UeM7gcdTc2/tUMIokOjmJG3U7vdq1xbAKeqEc487k5HypX39QKS
HQLuMHnhhk0ZgLL4zv7HOC+F14fHb//Pjn9TONSR+PiOanHq5jHw86LUcVjA+bG+
kGjwve7wFaTLMGU0ssYCgEEGCgV+2fAVI/VKCZ0WfL/DceZ5IteFX0VnFLQR/+bH
HfqIXo1jRnjqJ+pX8TLNFJBgRPwqB6Vk82aqmJlRpJ5Vfb2CYySUVhRsxNPsRjCA
bsmCaHhYi/5Oeyyfit4cLxAmRuiuwLS1LYu69yUz73YRGgod4er8KNGsvn6Pnrdh
/28Bgn4Tu/zT4PinVTEbMvJS4ucnjbd5kMJ5t78B2FZ5HVHPl+Nu6EiXoRcxXMcf
ntuy7TWWcbwE1PAer1LhPKf61mwNmMtVIJPyg8zsVWQQCA1vAzI+ePbyOkeSwpYb
v1j16/6MlU6ERNy5C3VpD3/oglk7pAH+CWlciUQrn2hxd1mdWzJtpj5L/pqgo1Az
GOKy2fpEsKztljO9Q6r5TFGXyovWI7y2NCpQdjngnIPYRGg/nTgLtCM3EHOjcmtB
I/JI3ETkEC9Z32RjxrAcniWxex+xQz28ZVeZoIrI5lidBzrePtV0/mUbtZz+K4Zb
qKDsH7Pu/dM6GssTCSYmViRCTUS0zdyUR302+XcZFG62l5rlIJjGM9+4HN8nXLuh
Z6/V22GIQND80jOetT6o0bdYANfofMFfEd6u3HoK5gT2UuUeYXfopqGRIgCP/jB7
YEDSz6Rjo0lSEyghCxMgkcaHNIKIXaTcn92mUrYVvs9fSfuWc8pnINkjMnf0zrvd
oFqHakBHQ2TqtRDan9upKWm9CFcbqjjYJqVzry0rC8yXTVH+8DejwUaNElvcBG/l
sOcGWpLuAfNigoTtIMZQKteNVN6Kff19LC2kcr4OMRFS8rGKhF+OO1Gx937nMwl4
bSm9qUMO29pcbN725u1tDh78vUbnbO99MowSFNBkUWrb8EAGZMEZJRIPPXMWi3yl
XEL5ylEj8wD7lzI5C+sIhLSnf4q974yh/gOGhmQKdfAAJ5r9OE6UsMM+q2+a+FaU
QuAkJ9yHbfaJMnM9VDhy8IRU5ZNQqx5ytxp0eNxH147f7oRTfui2F2TcuNuIlimp
2OrHo9Q/wnuCyV8/0HvujlrvwI+sZqQhS1AcVewnmjr2068lwI/Ve+C/Mg8pUd3k
xL3pYDO+PAo7ZUxtjqQjmB8wfDrmK35H7yrRF1pgKP2XIHRHEOVsQ3azlBaLOx7E
7J6iqiou/apb8e8l7hvhVG+nWklPlIMjDV5JduH4knaYeGhBJCaxjDuSVpNmrnjh
eWQYgA8ItLP2ZyhlXjUcHPzrka0sgdk/U19/xMbCk7fIzeRsd3jPp+PNQ/8VnFZ3
X5qrGX+1t03Yrf3fYFmziIsOkRYghw/MBeB0CzoCpYainH1Rcq/j7O65IWZ17fWm
zCXkMZc+24hX9Gx0xStiTDwv9qbBJCq8TWZUYHGExSGdj/ytprkTkDRUgaFumFFU
RMzAvTS4hfXGzhzsxH1tUZ6oKl/8QReyxfn4xtcMZVXpi+If140WEouc1gKztKiD
DKk1Eo3NQr6UaQMu9jc0gjL15OmM6A/kWDmB2k8dltDy6FHXk+GSHCEEzr0ztV8f
bCslk5QErHgjF6eMFWoN3VARpJeTC5HdtZjScg0yQq0F4D5OQx577LT3O6pcYvyu
o1PWF8MctVNLgxWyjEgXtjBiFTcwkM1NhXQPPDIJ/9FQMCo7gSjOLnxWKVraI7Og
BcH+J+nNXcgInK10tuhmrK6E6NhihYPyrRQJ0pk0ULjFX7k2oOwnhi3NoqMcJ9LB
WL2ZaWCdepYnMiuu2vDmIYYO+d0H+KtXBoCvNYTv7+6/WfNhMQOLneJBhyjddVgd
x8loSKwqs5XeLVE6BfEy5Od8uPucG19uO8UMmuebgfHlo1B5kejJEVgHCV+TnLxv
97MmTdrawNvodZ3AhENLFZuvhc7HMiz5urewbFrraL4/6xDFqn+AbDZ1vzKGed4j
xd7Lida0J7cnsXEODKzbwObKBmdQOa/JKsSbXwayprFIuGHL7UsDa+EX5pWgatQz
f7B/jewjN1fBdmqR1DldKlWQhpysCbeaxKUAhhL2bDptXFpMbwsurcv+u6634r6I
+w0NaqwjURdz4DT9TDokih6lBbQFas3vfhBTxdMIVot9N1Ky6RLjxOXjf2jswZc8
+DKTpkuMZwxgiy8jLHVkByzqhOlmuM4mj5TdsoCFAy4WfMhPEIvIWNH/hD+PJCLf
kI9BSPdJ7crcSKoBQECLqrSX7BCBbCSzIfHITPrWGeYXt/Jz+u+YBxAZPIIf1vzQ
K7Sdb4Z2192PrcD0YeojXECbU0bkDOw1FSwBDciOmsOrjJdurFSwg9gB5x7OGJ+u
JSK2UHMiY19OX2G8q48CtNdprlZIJEXYtwa0/Kg0giOEmCjtH4O0rzbv0SJGV5SP
LS+iFwXjgi7ELDzxaWdH9HBzSRoEJnJRdkft9G2K6wdsyL7T1AbjVnPvdkD739Tb
7yzTuZMwLatxVDXH9Se8kSJW3TU3Alya5XqLTAlkYzGwJtGzwnpWEObSy2m0APKX
mZDHQBx0DG4MD+f3eyMCYbwsNcXC6W7XfjPuqRIlq/Y3kXjs2EKoyFznUcNSQ+de
UlrxSqoEpIyIRqnkPk+1mLwEDwiO2TD3H5H4bxkBcpAjTHJTNX/TQ6LmVJKMMx0g
OVeqhkobCievP/3pk5cHB+8HC82tQdTt6Cz3r8PP226JpeCxgT4sQqTa57tY4bj1
alQPRnhfCtT5imN04wUBbfpl10IQn9Wn575S5ncDhHHDhkw1NoUhZz82c7HCuY4t
Z45b1nITLRY+x0GtXJr9UnyDvTLHt4iP293+owcd/rq+jy1oENJBZsSnj4LXUA3o
fE0YuHyunDUcasurG5RbB9sUUBQ8yYQKLJ1qwtfhKERklBCcoWzffAmKhsLTR21P
ENXuEwE+kUPC3+qKMmVsCnw1Ivs2WS1UesXbcY0YN4xjwKHPclEwm2+C1qbU54ng
oz/MCMsGLQOgHftW9Dl6PwuhcHPml1tn6CsHcfYjkr1zwqQeWxfMvsYxepJ61Uc1
+VacdlEWj3b/h0dtC9c/Qo/n4pbhT7K3a+svY6+2fwxEg1SIuEu4sARFS2W6a4kv
9dz0oGDwp78r1AkGHe3/q5onKW2Ds6xW7GjQXWUlZcjWMCHFqCXoMGj7JRMudcJH
k1BFD7jc+ZJwM5pqTqbW072ksOAL4bGGI4bvKTwZW4+gk9r1wEXl9cHsXRcpevcP
cD9oegNKRsfYAFQQ8HyADovOj0juYznfnGCOQkxPsfoVxO70itfaPB/c36iEA8rx
zzZDB85Ahv7Q0FgQNOlmw77+q6YHZQpKvTwleFZjvqMS7B258UWf60pjbMtsbDcY
VJ3MpB559vA+obUPUGH26TXPn4gznSFpvz7IQzKLRMTtBcHPDWv/8+b6k71VMhGu
BaPpkxJnzbEnRbVe/0QqqHmRO+v0WgjbJjo5uRk+TlmzkKbKWwE3BGoGIwZQAXPM
E5AQuY2A93b6r9ddhruTsd3SLU6M2xJ8BMOuJUYxXJqXRNPvROojHkf1SI1n1fVY
mmQZMB1h38IRr+eIy5LYWDE1SsIXKfLoDVxE2cT2VC0K+Bl2fae/H0x8zv8z4cHM
OJwrXGpy+uG2PMn6gCleNZHi3EQIzgjoc+Uw9JpJVPIoTpN3vduwsNzSuw4StrMq
8mNLt9QU8lIxdU2o7LVoQ+h3Y18DBBT4P/BpRBTly4dTXf+XdzSMDEbTLwMYNQCi
DzS4+Ep9oY+N1Bzqg5tYKkFHKb28VAoAAxOW6Z1n5GgtQ7+8teXD/3+TRz6bS3KX
EJ1gFD/sEnQhEX6lhnrK4wwNCgZZppu1KgTBW/LvDSBksiIjkgvZwy5ypMM9EGfA
n/2mM/v+abyUy/q53rt4G0mKVE7hnhlMTVhgNrM3xfSmMqR8KuXv1RB3pDbCBDT1
zl5yQADzNuPGwRp2obTXiMvvj06ymHMapZzcfDCIJQSw9Yss9f6m2wlgWt6gTCiU
1aHha22zsN8OQblPtZRwU9ekvY5JyfMKIG0tC9JWh10e/yv3mg1DvQf4buIiFWAq
HfRpuhC3zgy8yBL13JP0Z2fZzD0oo/feUtuLGb+jU1VP3lgzV7v9ffEzanY9vQ1u
py7Pn3zS27xdaxDfRxWWW/AafNTlfCPMEX/GoYIjCrkexmuqAoWlII+fI1hGuGwf
XyemwjEPijyTbW3Uzl9MUNAoPFL32X3EvcRxXxGqmgumEPnamBCDEoeHzeJsSz05
DcvdF8ACkCj3vt4odm4KyvBT/67TCLYKZwYhfjfOl0XjTLa3FYsycYD2OML5fli3
w0NOdGb7aIfeV7GhVxMMOMDxxqyE4vR3t/WKN5VqgIoMTRfDmDJWXLWVLpF4V5Aj
uPNrIgyBYzd6fIOGP4GwNYeBVls4aDWKWU8f8DtO3VLau8d3y431L+g4ReOZX/mF
gu1WUVdyLdHIKTbXIE1biPkczC6rqdq4Gj89hBumS42ngxpbmMOtIL1y55TsNNwa
3bliWMFg+F7tjwiY40KZp9xh+mW8YbrRDz7BvWjKFax7Kd5FbHVWdcpHuKquwYvw
W2p7fqQEx3EsAeW2H+bbCwrO5Ok6+OKfo6jRJOIrRcoFHajXVkQY0l3QigPI6P+L
jEQSCt+UcvdrfWhUbyfjQRlvBvgw3yleNqIlOx3D+KXLphBzzsFGgy+tEKWN01VG
j8fV04vTvXM4NR/NEy8E7tVbqLS8/VeBvfAwLjgCTvG9asmSgdAfFyBDZGsOvIov
no3x9gFlfsiXWiLXLVk8gPqOFSmEhZxRu2v69fREfmfSLjCur+WmOn1DCGbRLfnp
u3Y9mGtEsAC8+TMx1Cx5jmDoqHVwzjKQCY6xA2pzMTe4leMPSr9GVeBu4EY+8p/C
n5eksaBK5Nn984036r3KwkoMuFwwL+R4kIMWF0+lJVHWkGCFyrfCYU2qIGcZRVvS
6y1yE/SCcvM8EeIH0aPqXWGsT2gxKQkW5jsOvjta3kGF990ZRF2ccS6wpskNlYvm
/35GoS81zGjx5RBH/24LrY9ENhn71un2ZanggQpso019XBApNjCLBAKBiYdObi8I
6xl4yq0hgEi5+emQTvyeRghZMO0JXv+qsze3KzedZUt3b7vh8E5lYE2WDV5fS/2p
jY+Ia3Dfh4HTXkoV0ShkBvqBmD7AYHS7WlDxAGshz8H+48ilS81fd9s0kYfBdHDE
i4rP7hwv6HSnj4bFhx4+G+5StcZfNNC/JdcY1bUoHvDYXbQ6wnPYyT09nKyFG3ug
B/MC7pUeVyM33AGyUQRw8NGQeP2aqXpwPkiIwy5ODjdTe4Aqd1psLBYKNBWWwQ2T
wz67lgRjYkYlEcfk7OEkkDYikeZcAxn0CUC2QXFhq9dTcOPc2qT2URXms+gsMm9G
oiWf8YSjyotA8D/mrC5qukTdXo9HTxUkjjarBpnWnRZi7S1ktb/W+4VcyGkMzytW
G3Y9NQx+1UjUlHjUYBCk1HtwxsAZCfwuUHBOsLA3fcr/QO/RDy/uiLx8gTiO/4bK
aFUPrVBS2d6/cpFbjiHynoCDf/5j7w71dZcVKYarApLwvi38qLP9XFcPyImA9OOp
w4I1EE52N4saDLOHmx4JR10W10lqhRHZ/817qIooK45+IQYtvrzXHk1v4nzhWLvp
0Es2KMT4flW656qs3vi/8MYBIc5C4uPCAeLi7MF1dp6ru509qk2+Y8qP8KWmy+cN
GT4YVejUWzmYPKWXf7ztRrYYqTjkm5UjP9LU9xQtWmUoH3cKI4ogqZJJBws/jgot
6qmFzlBESD0H1VAezRKuHLHN8OvhpVKKZyACOXCYgLD11JI8/y6YKDgzT6XkyK1h
TH+QnE00QUvhcrNzIPgF/0Tw5l8cjnmia6GWkmMPyHF0gm6ibdpueZ3qR8enUjmJ
yHVnlgEiIIjfpEHSGtfTgTt/P93GIwcmQ5cMvUD8wpqbE6HAP/iCCdZ7VWmIHrAT
ECtwDoPx5S5DTNNnlp1FOZKHmkecUH4zQphD+nynKaEb9wkgWTa51KBYquR5u1Nj
9jVYLnZGvozj480DyOxJQOHgnwkvzUIwvX6psQQumtnUvIyIHTsZ7ixiHVyLHgws
t8agdwrCXEYFQkKC1reODX9GJmgxPz4doTyKubiah8sR5zDRbrPklYbGoZMpu9/U
5LKnpWroeW8atdSCDuc78cy29t7pyeE3llK9S2ajIiy5Cp/k0Bm81eZGpqQnuBg1
82TENt0EjmQkyjMGfpbn195yFquLVLXzyUVamZ2Hoozff8xhJnJZNi63CjkGzwaj
MQVFzKhksAiPjYnyp/+xl1fA7BE59Qlzvw4Us0KGZTozGpdwBNW1eVndN0RLHj22
c4h4oEZuJCVW4UAu5D5mwRXW6al7WNxGVHRWUXR4tY5p8gxzZFerwg4ObTaKhZtO
fMgSmkQLYO9Pv+HDf70qhNkMm4OtdRB/83tS2nygz2QVG4yQGSob6lDjbXIFgqjc
Sa2pVKQ3up8K5QbTLg1KLAmxuHKQ22Y/sSYuyw480yAM6RWKYMydD+DW5G5F53QB
Zin1DKlKFZFMHDybBjkHlrW//1fRwz+RYm2XNkiLXzm+mMbx2tjJityXSDmn5Mkb
biL6EXSqKm9Z1V2DjjtTm9J+FgUFEZf6BUY//XTsranFFk05l8mDZW0eeoHtLXGb
ipuSwozJxQ7vRZaPWwPijm2a5XHfvyEl8OIp1N26b5Jt0hH6DkKwDm09QrLCpH2I
keZedvKwksZKHnaKyxVTFxAlOP7Oa8YwpzDSd/IXaKY8s9GhwC+lW4LvdxyP6xKN
Nvmoq3Mojf09CLfzAlivtC28Dho6a9SYXHYQJiiyuh+4pn6HNHXc0JOR7lUjxCp9
xJMN3I1L0eSeHxC+oCDUDzo4TMnNUAW05h/9e304JEZlJ13Xvtea8ZuTgzXp+yyf
tE9AIJzZc6Xt+ab/5yofKOstbVXfXuWBjIqdSkrfijln88o3w8c90AnVcFeopJLz
TfvuGDJPEUDQIzZTpivmckKyuT4JLcQeqLUILCedABFKG99S+WHh/0DwshpC6hHJ
a3VMWwuuM0H2Y2Z/VkitWayrBzsaFwXYNQCi2GNlED7nqR6qU1Rw5Bce4h3I3az3
5jClf9V0iWrn8aPZRco28DcqdnKap4Ub/69tWYZHePX06AKBussgNDbCVHswyurW
0Te7YQdOueJ96RCXoPkCMyGtKiOFuhDGYI+gjnfY7GyFWs71DnymnaVoaAVq9sJi
XuWU7i/JHQdzQ/+8LBJ7izeCvOQBwXElhcl7g1GWPjeaeoTTdCSBjPEhOaiy/09k
SqUEFBpF93OoxdQ67cCAb+LDe4IuGSR4bNyt2QvcXaMe4MXt0H8emLTeU9aOcvn4
wp4Luo5LDXTf2ijOs9RfnMp7UTSe+uftEIzFCMbI4Iv0T5rcdde3rv90FeZiNlE2
l+ob/AS3I/v17AgVAaNJP7/8vSpSYEtXTCDk4+l0eX5AOlGwgSIMU1t15D7mv3vi
eC5Ev+yHeB4Fu58ZEqnrkr35oRa3qptwxWgV4ro63MK5EmDiSwZf6kyXozDjMV6i
xCnZiO3vCRquYLEQ7fXqtADZRo1KLdlg6c7IEfogz+cf7TuCbUjXGsAx+rUZS722
lS+49gRkgfyToemejpkUcV5SSSdLxMHeOPuRddNU1Wk0r1APnl6o4Et6g8GDYi2B
13Mu4Fb7GkmhMDRXRqlT9LN/I8QW8f2H4eBkYfga+8nwqiaaAi0vU3MNyjEMAp5L
KUlzkenQV1ZzP9xDN9mhhyLuMuSfQDMz7bMwJUi4ZuqgTeKehjL7UMmjDo/9io/8
/zcuHdYS5r5rFMXfR5/QtA+d8SRpHS/d7MYQbKXzer0+okIULEg+p8GtO+9TYgDu
3DHqtL2AKy79ijs9Ehn3VY3yegdwrWvU+YSAGbxOn0KGVMqhR7WfX7xDoZ2nmWJ4
CvvTLAuehXcsc585S5ZsexzQOp7OWxVwcVrUYQ7BUuXYJY54h5lhfjT1d6JH5l3x
5hyQX/lgrkziNsGOjiK9KNyZ9Q+ePB+kPzgWK7w93ck1D9jdJbqdJH+KU8sDLJtC
I87j6widITwL5ZCgRFKdDdY32AlkrTx9Xpw36RiDUVkKEvjRnd1RVX7Wh1HahhRN
xAAclr+e2klUzELjH9jPQV+R4iLLk5zqeeVUXfMxT+4hXUYlNQ8xRbvTSE+FORq6
/Mi0uBn5IruyEM+AD/5qYJ6SXo4dkmSbKTfoG2/E3qgkzq3+JHDnnfb4yp7qgRmR
yfVnYY9S2mHLYJt/MyW5zgqHX6b3spTdODy58VLEy4dv8TS7GSB4Pd9UigxY8ErH
2iz+6axopbbNyGy2w02kUtBharIKstj297SQDWnf2FdC3KIEs6qPuYkkbW+otzic
/65PrzhzITdRtb7TFZmRHK4DiHmv6NsBnZ23h246hBCLrbrCAHpSXMOHZTFkLNgB
hBvwhkFqWEL6Ps/8VdTuF0G3RZnRh1A3CTYRDurHTfWlr8i5uU4mD5QS9HFZwY5D
8vlqrCd8vtgKSfuPhkqDpoP5SZv4jKG6fgLJsxEcSm6XCbNHVDim0KtAKQ/ga5V+
94Igmfi6muOtVTT/xyJ0FkHI7AoPibCkLlj1xQa1eE+/v0Es+eV/s6j3NjFJcpEo
B99g0HK9UHVzH733TF0AmAFF3JM+BbrAUfw4ERhwe9Svh0Jo623f+dGaIF/CJMe0
CbonQ2ZRjSpc+IC9aT/GA0OPUwoOvIGWthGJ5mAQHbmIrRGGx7YH9I0yC2o6onyg
Te+ELNipCqzHTdla0hDJ4iipYqNG+ek9+Vp7YXDmWzdPiGP49rB0LgAessouM0BD
oTHN8C5kHthIqu/z96LC2yBvzFjMsHNbkdfdzSQYMnFPdGvqIkegt/XSwuU0jHnP
nP5hHKG9QKAO6JihofgJzgVCVONhejn2rsjDCaD6ItJByDWVqdycdT+1oXp9aPAe
M+7vLyGdnVEflhaFBvIdT4wHq1aTVhczCxldpnX0jqbVoMVrMK6D5XJ+7zvkdaA8
TCZgr0Rpu54DYoEOBU/5/03e41IlgfxrHIP+Wpo6o6KsayC4qz5I4AOUj7raiaa9
I4RyAlgclmJI32TYEQnKCbncEeRChx5xGTauI6Pw0cEq0R4df4Keppu318E+QE5z
CciZvDb2m+9O+VafnyT9CdM74jluekc9MjWl3vLf7iUJTfa6v9BZFw3rMzK053pJ
9N7syD1GziTWV8+2ka8K8HtXGzSphejJNQ4Y8P2qUCQicpIYFafjtqb4hT3X3Ds0
BbXJ5b/JCodHfUNlmukvbbz9Y5Ipb6G6lgxmwk+qDD/0cmghxh6K6pqEU8405jHX
1J7pWlOnZa/8p67QBTsFaubmmVY/0AmKHafr1xT5b/Gxc0xX4VVYD5oBjwR/wEVU
j4s0ZM0jA+iAl3Mu4ySpPQKEWP6bv9O7m7ygmEADCdL9IQHUS/wnuzpbEOsL82bk
aK0o19WRKenqJXEa8YvPxRY0chpV1KveD9Wjf1ixD2g3aIYe1afMpMyHzmz5KMoK
1PiruWe2vVBXamqy/alq2fo+vVdrFqre6r5IU/DgzDyZJaoiB25jy+r1NCc/duKP
M/1YWgOhbBd+oOVk8bulswHf54O4EMMfKaaLbNTLU8TGzMZw6UbdOcQ/FHAllDml
ecZVJj1EtR09tl4tzxH5+aAhFo3RJUfRl8nIq6+FLFX+tdF8dasRD0rXuqyW+B25
43gwzKS6wJfDTvF3GGUqYod1whUcYJrRumPe/ArIkdkiSTfUvJEtdfsJ7hOPvoBE
/X8XLkeAukvY3SM88VXRAQlMd4iPeBz1ytULHr4Vp4CXEu1FA+hmisK+wymZY8pC
g5pRQFxrlRR45wsxHPxxwZiPVc+D/RfCVZgZRcPuLUCjrrvrNnaxl8bt1XtDZS7j
aVdjLNnFEMYf69MXwezZe67O1cRPvY0WeQt5wGrHZmRLuIogZfgBcgoqXSZxBjFf
qyPuZYDLygTLbh4qcTNrKV4jD/MRvGNPgBodXXsUEMUENcQ785BMs+dSVbHlN6AX
Swj6c3FIt4R//UgsTqHQmdUgFN8DRKCamcQvxX+t8anOfyfxEx86WP5tEUftXASC
1PN0njG4w5iIbJrhiB8XLNJO39nY6dscv9vg9IzWOA+O8IVjOz/FUUtLSgTerV49
4RA3MPGKI418ywcAGZukAx1OU6G8T4J5j6Wope2IaWY+u8ZfRUPVqx+N8kIpmeVw
zuMB/hNW7Qv4VC4M9nWJ7hsGenFCnJBwrwhrfCKebUbIWsOe1uHctWh0MA6kLciZ
HJTOOyw9CYeIhPzzplb1Jo5SNFhpmgUHMy2CWUigaHUE6Tne4wX3h/OKMU6G96pb
GloI5ueK7F5i/YMSDeCrBh2PWshT2Xb54lCwFnOaWfj6FZdYyRTTxyTxH3oOhDa6
u48RUzursbuPluv8tgsJ1P/jIXB6+RB77o4z4xoj/r77+snuh6I6EOKA1gpUfM5p
hR588alEZWZhZ9b/00JLfktMkJeUG0x8tWZ5XCer3E268nnYUVC747JtAYZcnnTf
9rGdAwB/dtj/drEK/i694jdp/nBdpx8ae3JUu+tFXsL2aBk/ytLWojxutm3ls9dD
AEJCJ6H+FradHB8ySmnorCZEUgQGQfWsAIK5mwyM+oc8Nz60AXyoB1xEMePq8zyd
EJpaZPQpXmJUmp97i+VWREn7HEPdJ7vF8JWkd3b5r8597oTq5hSCmw+I0kvHdhOF
yJN2OcfoiJ6bxow+/W7VW/mlAhhIJfVo+E1PAbiFxbLuEWiNZPaXLBwvcRnOEmEx
8k5bDYoCBQl4zm4iABhL41EvGOAOtJdPftbgpc/Utyo98ZFHwvClspDdux0BbptB
pV6d/THzi4b1rxAyDfK5oduCmZRAgT44XZ3NE2/DtfEh8bXwUbQ5GH6ceQ2h1Epi
pRgkhiwEVjNAsg3MXA1/RVnUd1Vn/BehQia+L0RtRagFb9BQvcg8FXj2iLVH9HF4
PnjY4avMOYts8GKV3uga6Kee26l5EkpAWSPnoOxVd2Mhc/hEY/ylvkVpIpDwS0yb
KHyV5DvTueyVfzYgV86TV6XB+q7Mnckn7H66ElLwjFdz7OJcHAN3PXoINbZO2g+i
8x3vnU3PK5C7Dyp0eqZC8qPQdI9rLB8MstCeR1TMb4ToPy5zL4wB1K2iXnFHRCpj
MhtYh1oGqX7k1zI7OmyEt43qTR+SJp4kr34jLik5nm6F4u/NFcjcbgiNcCmtzNsv
zlB6r3r45VTdrk4HU5qKe/dCF1fueAhMk0QPVC/ByTwfCmdzUmNScDWeVuElh6lo
yOWkdoLJrB6fZToQuaSiiUL40WXXGR2VHeJeL7m/v03nOGLFgDGS4DtrlJYUXqnj
5YGa9jd0L0HcwEKvueJoHtK7Bfw6GeTF5mWmniZIl1Z2V01vMoQKpNmLc8IpL53a
ePBgvALvjEz4WDnj8NTmTFkmW+TD7vg2JYALOrk2fmrIeX8Fmhznm8YGLhP6WdIP
T4g6lQjjyWQXxTIr5vJnDnL+y6OPO3Yg33wMLNSnYpHzSFLKF0HEnr1donjzP9qM
i3qX0CtiwWXz+jsfYCxYr6MWDov5IQgY1ii4oFj+pMs3wbVzLP3/JPF+prtuHbwH
YjRV4k6//tD9bPCa8/XyXY7yhrF03LuIiDEGheME8DwOKeKg/ksIvVfz/03nXoQc
lJX/Z5B5qrCtQfmwVvEhOKfX3TAzOANZnDvaeoP0b5Kx4jMyt5VEhQIkZLRPmjUr
MFG4Aa2T53AZ2L5Lzt1vXm4mlp8COKcX7Y3WpNovaOGdpXj/f6YrynrNTBuVk8Fs
pT/2MnwB7EZaheGgyB7DtFXnRvOt2KMm1LXLOEzXTyckv3kesdnTTU9gIDJ9dxQs
VMSkrHn3aCrw9OC7kAsLUsWFxn2xVWuiSwpq0WxArj4w4L6KcIKAZ0O1gGwP3ogn
gbyVNkrIzhJ7vY710wkzYD6NTFns7OkL3MVN5WZZNaPVmCp0taeLbMjGYiMf5j4I
TGRJ7fm94Bl+dB90JYDwz5fTM0xkDLptHcMpisZWkxosRlAKW4YtVUuCN6pAHPyV
0eCiiSqEmMXFRK7Raq+U1HTdA7PhI5PgHGi99CZBfFjyGkUV2O4ESBBupN0d1zF+
ew4TjhvAFaLevHBkSlwv3Q7akGK/8oafmQjJiLtMwdGirja066hyMHr0xVjtjQeX
E9xnHLi8bD+Mr961ilh4PGNqkUdlFetVDh1NPDBFEoKYhPHxJquXN7DLb85SQck9
ljGYK9IjJP/25zamfX9u35p3QJuZXGHRbc2Br8wfPuPK2CiUrD/NVctlYdGKYMh1
kz2ah39rcJGJ+1Etr9IO1IbEap+/WVB+OGajNIyPvK9DTqY6S0jZVqzV1PuTiuAo
gZ6mWs8hqqJSRBNev+GgKY07Is0JsWxcNwbhVcf/TZOFvXQIYxzqCP0PjGYREP0F
VRm6X+PlV1if89AQKL6WCoqs9AgKgaX0hY9OOIqOnPVfa+eJWCyXoD++6EoUd185
pT+ZQW5ZoyXnbA/Hs532+vUFfkH/jbrY+TyRwEdwhanBFWq1H7bA3QSVQE7Sr8ky
weoZ3wRYfXL6S3Fe0AYsVmazrSJQX9YbsmFEIjR9h2TCKinneC5OR2vrGyCtYCvs
aOoN/3qwzxNxYR9LlqwoU6feTPFmGPo9M9dz6eMrQg4x3qDExzNRQyumknL+nG1+
f5ISEAMSOiqwlWp4vy7hLuo1g+fxkJKnclR+xY3f8EOJ/tfdsAJIvofqx+ivrh4x
e/dOCUH/m5dg53mrnq4tNUs1pmUhZQzMstifi2NVFrzqaK0xyjL5TZHbNMgP5nnq
CtLRq0x388EuowCgkwOTBX1OGxqNXb5vTRLIaERNF/hi+eOwg7wqjforkBIJS6Ya
jNLz3/1m6nCNiOhiHlwjLctdi3R8tsRek3dp995O1rqUKtL2R5VUofwh3s6ScLmR
dr/o3F65pA3567O2Qbsa0JsAkcWvIfom+7rM/W06V7ZKRscQ9JESFzovr8gz1sxw
xyX1QrwFAMz6JrgK3WzHSmxFTLT4r2wyaRvEZsUdSJs2RXQ1xW6Fn6YnAEKZTJFo
cfDbC1rWL6q6u5aVwUJjJcRqZXXUUPXjfQ7dspIB28gBtrehCZu85oa1ga5AF+NS
CBfvQ+R5PFkGboSRTpc10uWVx89fwlcvMViZwc5xxTYRtjhyfFzKtxo0UX1nvlPV
7CQ/lf/T5Pryu2FxHQaMmzfqgwkMv+rNgWatZCL5EVpatRE0ckKJoWMWqpT13XG6
tikeHxC51CE3ND6W2vK4Wyw8G7OngWNl0n6jvDsrhLyNglStOQwtgajpZoLiHWO/
JRYEYTTEXd2cm2HMs5E326hsZQCxItRthxKZ72DQCKj4fXdQ0A/o6M9wn93BIuk2
Dcnootqr5PNnqcWFn03FbTkTiaV41HwAEmbrjEh2lzm2r+Dcmy9aF/zpJ+a+RmoK
Lwl/GWumLMcBlhjREnwCJqBG5WEARaJKWQ2wnatck8fCMIj8jH8QvOjXK+NWIm0G
uQNlz1cVUfJL4dDftEQ3vnP6QxqrwrAE/TKcVguWhv26JXtvMmw/NmCkj8AzGj3E
oV5zBLWRcLXM8OPaszFgV+pPghl6pNToDN8p1GkoOoLVb/T2LWZB01ItHD3edIwy
Q+7u5ZuK87vjp92vWjfk5JljOlo0luVG2QfXdNXytatIDyz7q2YZF+iQbsEsfZJj
V0s9AOwWajouwRU/PU2Ds6o84B3TEyxpzrSFsguv+1cfN0e14RDUBbcRADrtflDI
/bloFq9nVtgCc3lO2qMcgUIQ7aeJmV3kW9zWqim3oyBrsX2JuQYykYNuF4HKGGVw
A+Ajd+tLIWLxeFr4+yOqT5dRePWaBow2MvddCiYLjRoafmRrLZSbsKLoXBUH1As/
XcpZ/NL5bjIQUYYEyd7IGhBSghdEMaeG/ReVQ0kDVC/T6EanWfCEnAsjRMUB6nvd
5o+lRr9l2ZbPrlL2Xrf1tOJvt22yR1EPZui/++EceLffh/hoNAOt7BIC+/7xSxH9
2Xa2Tq7QaB2mUE0lQcAGwsbm8KJpAVVGzMSbBXWWN7wjOBLMa1y2BPdZE7XHfKCi
41pb88ErCiKaNYsztbMrqXPyZf4H+JOSR6RgwlPj2MziVXRH7uYJhbFiyQWLcK4A
r1zvy9k/sI1u5+AZsDPrMGeBNucilOmh/J0EXYU6RGCLAuPMW9l2ublkZdbL7fpp
o/Yi0NlzT6TpdawCVBRft7A7curm3wpNq6rVnKEvkLWba43jFoRntD9roggWF+aK
abuzxfZMWIlG86RTSn4UWYU29fd+FGwofur192WJB8Hk5Pf1VxZCI1uJ9j8Ap/cb
VRY1HnYQ95fFLWrhHYFJpaVXWR6OlvUPbZN4GwpWKsawwrtZaZI4QCo8NzQOjKqf
7vH0Ue6R2OxJZSIMRL1ujQb8pABucUWhZjBtCVxf6810HxVDpJo9vQDhT1D8p89j
k20kRJDFNnWIKULL2WOeYbf+rnqbLCyCCeHYjltgejjVujn7axf0hR4ncoiBaY1w
JlrVje7A11H47C3pxZ05rpxwRtjyLqhzkPXIMoDR9oFB6ufKI14tQioz2Q0SI1xn
3YBK4pgqduWUBi7IPwksDWJ8KmNTqLttAEOssXcjM2iOb1Y5lge1aeuExouPtZDd
mo/Pw7btHSJs7at6XLD1b4jWGayhuUX9ZW95TW6a9sPw1KzDm4GkTnHo0P5Mk9/z
3Uu69t3xffdR8bAznDO2CaAaPMPmqEAcJxeLAIg+ouloomegaupjr3jcxdphaN0v
BgxmIUHsvXnRCMmjQ0YFnyKqh5tzZjaM3E+J1KFU1OHMbC87b1Y76CA7QIyoE9HT
c/h7eiKYxJ22PQQuI7s4rag9YPLHM2BvnMuANgvS9K0G170ZKEBsah8Eb+jnTNz2
2Y2RNuGzUrk0jHfnQdicEh77UtEufwLTRMhnf1PLFArOjFWfPvyJ2/ifdoc81kw6
eMQj3TefSy6sLRhAQxA9RflGCMSPoCPSbBCKZXgkp/auyFpu2wirZ8MvjNeqBpFC
Qe8R5mwHXrR2EadmR7vD98D/mPD2N/L4vc+RQzndFJLE1gzj79lu/Wl2l923fwV2
5lVh6No5XHMOyimSAXe3odxhm7xsBoWLtH1EHCkQGNqd17trlzeXZYiJa+abGEde
O/iNRqo1rDDedBM34Cteriyr0L99XsvSI4LxrbSes0acpFv8VysitH4hz/teU4Bg
fVrZnk/jeqv1n5sSRjbR83VQmuDoJCwhpdfSDG9j/eHFUwqszyfLLYllPv/CLXj5
2m0B3PNVHvO2rfIKpc0T3iTPISrCWgFkshQ5igi9MKRaWcfnNtYiDeY12CR1rvUU
P3mmyJ1707e0Dm2tKJXlX+k7/7BMeJVTFFXdveiAnthd8CxJD05c2epDEupCzJqw
H2sBXJMu0u6O2wNMKTfRZC+PpX49fIcXUWGQMhz5yPIgDzm70QSkrT8gin5FsoVa
oxnFCLHgbxuJu+YFIe6mrjveNOQzGher2qYLCdW6IwbfvGqirGHO+4cEQbg4gxpQ
mDoU6ryDhRS7NPmzHOdOQIgm0osGfY5cGw1FJ0KFP3Yvjd7AbhN0oxPKcNm+B1ET
qza4hqtabCwKAUPlCv6S3zicXL3POWScsn408/kasa3GfevnMLNl/VDTtCrGItkp
St5jYZio/ilfeMWAbyyE2BTE4Tj91DCPqCna7xhUpSyH8ZO5/ggrVYJm+kxo2ACA
kJIXBI7SXYH7qyZ+fSSqJmjxwxqqBZAtrZQPdBXFh2sAUX5zpbVso1KFDdUkQdPq
kJMuwJ5UDCZ2xduQfBV+4wFwYgpm1/8cMR65zpcE1pht8APQ2ha29ga+utukbrgA
gOmwMufozzgiAnfTOD6vlWD1ewrxcYxoMOSIfV1S9Im+PkSHDn6vdDj8j9Qj9Kql
JJivyJD1f82WJ07X8+ENOg6sQ28PEVkOfBIn4GB4r6zjB8LKUyF8+fIKkOtTrUsJ
HgHP56hkSEqQsTATMPG8GrqwvibyjSy0/qBn3NDHBHL1Jv01U9PztP4hz0EfwXnU
pwIpBAplS784oPSXYp8ULQXWTURhhqkEEbUjHviLODaXJ8ISwBmvYEu6Fw03fEUG
8cSUglos+heouQs21/WDW469oEEMuIhsWRyisAFBH+0MjBY+xf5zcxAXQ7J/BqMG
3JBq+ZL2Ts14YKVUQMa00UAs+brA8yqDm2SY0RvNdChI8KdE+YX16o0rh7h0sIgh
4PuEuZMkVGmaSDk8l7pMRNWy+E3mlHAuE/prODy+LCcuRDpRsQN7u4kUP3O4Fnma
pWNf4OIyVTbugaWtpTtDSt4ew+KsVw+kZTe+I/L97j7bLfZDaIaEmHAdFjVFZydz
kzWtKu0r802EPoKP6O6xdZiWy0l2byoW+oz824zbGVnXAi8J/7eSADNpwcQgxzbA
y4Tijyyv3S1cpJnlLbxF2uxqRyEwAXRNUNry2IAcJaIVJMEma8r9eWvS32ccC9IM
OpWvxENmOhSSRzC1K0u/QElbvOxqMTzA/x+BcicssH5UTgMuV4KhC+hjMNxmtHLD
79e1ydZtovPHdyeX7wnYID1mv9X0znI5pFTfeVU6XxIDq6ZMzJd3yXAc5q40dqFI
CMrSMC9Pzw06VkTjGJbZosHZ4+fKjqVCsxR0pR+1iBsUWYo53bjYPhFRR7X/IMBr
+Y7gFhytgVM7xzbj5Uu/iG6dPY9DUhA7GSNCtmcqAo02zP1PDX2Sc3QJu4ohjyqv
fUXIHrQDas34kjSQVSJIHXzP+Si6f0uMCCJf7NcdVGB8U87TNJXS1Gzg3GAVOab3
anOjkxQaXLWaGl4EWucZfvey8IUkcBnFjvhGdObQsFzn34BXpvwEvYyRcv7VlvFy
BtBB+VwAxweckNrk9me+TvoSJ6D8KPo3XExd8g1zYJmKwTjy6dMMApQdigVW7E9t
A4skX+yedv7T5USazU08l37nPvUjDzuJatUw0fiFFric6Qs/xkRHsiIRGIaq/qxz
KgQuovihrZNOpjrKQ1DIVnsD77d1R8uIiZTaK4XBwu9Xpt1U702viT/XMZoAMe9I
kJMZadLwSjPyPaGOymXhjf9aRE1W39inARDzRLA87+asmB0IH3mXVWjhZn05WeBI
j1oYA8k3E10uhTl/ZijvJc0PCfPkcdVmM3Tzc484GaJlzJf1vt9+wbc2Z8YNvSWB
kcCI4BLqPC5fRi4XZ+gnkhpyOHiViqsnAkQGYjRwAk6IQRrU7zgcCBWR0sdvNGD9
mJU9pP+IUzwkjrNBGRB0H7pzPaT9nCVnuBJl8usJG2KqgX1uUAH4ZwjW4dsVwYyq
nG3+Rb6fN9SuyxAvSPXx6aP910TGIWJHloI4zQmu2dLjJL34ObRgayIyGEKF7vH3
WjO2OV5IsauSmU6pZUHmZ2NN+jscsKD3EDbRjTdqZyzg5yuBkc+n3wHrDk33sjT2
pN/gDEKkFuP7NMcixZZcEBn/YYXHR+L1ltKC+9MQ+qVF/QpIaRByAt4+uDDwIzTd
C7i0F4WkIAe/s0pxF5c80ScrTmZhpejxwOUI/NfMnMVkHdbHg8EOqVUJhNytXPj8
nArYdH8I6oOfKJeQjrizem1N7R2OtPJMX2IR80ACVdmaUKzNaj35PrVcVUr2d+7u
ilbOpIVySxE1Dhl8zV12elABAbfwZRI9UjVCq8RTBsME+bHtvWhHWkrmkunP+PV8
ZXgxx3nMeBJU5EGjYLo9ghdY6QmRnzjvsZMnXQsgO0NuEDq3n7vzhxRnDUs38RA7
jLQzREZYr9YGj/Y95tfteP/onALHbZi+cCTVj1QRsHzob0tTdhYGO6kYl3dBsaPo
7HDcLUuCcdB17B74rU90LzxPT4V7EZUX5IhMxS11jhAvQJubmdKQ0YM+3mZKSsXM
kOT+fq+kHPgdz73zG8YZXhtLtK8JZzQCiFjqN/L1eaUSBUg3Pa2aMWE5dReJyupL
sLj+H9hiLf+hduj/RySP15UdeFJyCKywcZwyt9TKX59du3svifKxAX6dnB5FerQ8
jJR+Sm8jU/cPu5+4mPrtXfheLsmHjbMPR8S29qO9igVZ5q3pbb/u/JUp5lhtadSJ
T+QZAiXbscSvgysfxpPz0s8XzZdisLd2Y4Io3XLSWIq7MZ7+6GRBjTR08rgjyepY
k5KY3pt4CpgxJ+Y3TGJXWaTmKoIdbCBdUaOU/xW/y4CTkHN/GwYt/+rU4Knk/itY
fUA6Wa5n9taZIJO0mSjcr17EIOPglsPhUl2aIBCJimqD/TyE5r+pGuGFTR3gAZmt
Flus+FrTU1Zb4ZgurZ/gp+0hgCN6KYpBowpNhhh0Xl6qvnF9T1GS0tI630ABzb3k
EU7cWU//gCiZMrXI3BoIovPKF5wqS7T/pW9gFEYfG3BbrcZz4pBJw/4XlVgI+e0l
T/n/KSlvEv11iCdg1cpYzOaF9+FYdJWbp+r5enYFdkDIWePHGT7B98tZmhCWQcfK
YUAWwSdULR/fSeldEMOtVqwGFAUibqxeQZw+06KCQJWfdg8COVXNQWLnw6x8N3VA
8V64RAJBc/IB5LchGAGl7sJwp7GcXHw4ZElhZBngoWx45ML7Vv5tHNuX69YrqcnO
rKBSIRci+2yt9aah8fU9IZl+E5jX+hiyo3XIUEDSi+YWlBmMhfkyzMgBZA+a59SL
HVTpWyR3WbPtDPw1iDU9LN85ME8mwzAXG2NjtdD3OPv8oEXr8oaFedthudCZbbtI
GT7lU2utXxtgFiZ7cZMYPHrzsZnWJnbrKNMzmoWEmXMH/MWdzzdk7cdLBJFPyhMT
bT6SRkxiqbkI1j2Q4grMgIkYflN7wdq9qNcIRSoT8TR3q8S+kVRcLIiTyMGoyYss
XTmUqTL8NTKIXODBHp0WS6PvOYAAkhoP75V3VfLtMB2i02CrNje/RvrtzDySQjUq
CyAzF1jqagb5BISBjqA1bOJblGrVWVpB3rLNyWxFj2WdpZwVSDICu10YqcDH3xK8
b8cMEIlpLKDCA0e+17nNVgjKSnwYfdIgcaJNowC/4gal1LfKuAiPQI40plnZtf0a
ZGkQIifjNE8YMIT1dtL3fJKO0XJ5uZVkTHDPSTqUYF7g9NRhPHhmqC1R9mHkp9+X
0LBifda0pnahyCLhrfZm/VbV+kdTo3aGFAyMZbOpH9CVfpGyKoMWKZayM0HwdRGl
4qwoieORNnKppt/UK8mMr4lA/A22F1NO0Ixv93SlAoAy9h41WUsabd8v0C5/GayV
Qv361eu6RBw5AGDLC9qaD3m+ZWXWoLKSXftZuUivY8X7YCvc6z7awGfuvHaRILgV
pJNJDyqH088alrBKS1DCa0y6UTVHVaRLZGjdga/09feMwzrg5v3NuXW7ug6Yr2Bi
6PfHgaSba4HAh8fjhaFpFbJzX7/R70hVM/OVwmwXjYg=

`pragma protect end_protected
