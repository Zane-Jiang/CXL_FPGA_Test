// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oKYOQ3ueDnivJcsn/2f2a0A7LlXtg7j3Cgys4lyrHSamcO2ICkMl7e8nYS7r
K7DcNmtoaOP6rkW73MKL9pPLbHUclPfzkifx7hr/fje30+PEEVfjQMabs4PQ
ZmHDJPfE8fOi9LzpIL16C+AcQ9joEj1TPX8S0AC8ifhK1Xw/eoAkGUvcGMDY
ZGoYIEU6XsHN1ZXh3Qt2UP0DAzqN+nNjHaxlDpf/JijyvQ+xHwhMckbijZBb
/qALxsOgSVHseugXXPptZqLX/lrNBOVzxeg9jl/JUrJvu2TctMVWlQFdGV+f
riPkl5GmbN93ChoZwAlACn4vkhThbXBAtDwHedchYQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CHi8V/bZOSdj43k2QmMo1sOoampbZCBliU95fcQodRv0mHL1RSG6R6fblr7X
7tviLhXb6XHsp73tyeMZblnisbGUCuj7RkgRi+FwNi+/qHlsraIq+tmYaovV
ZiAu4pWv/RJu21G1twbwLfcmGYgqsOjS1q93B6TRUCV57S/Zb381SblXND60
wpReSVVFOpy6ycZD9kYLtFZ6c+R65OIvI1Ui8t1mUzTuemlBPIQnwvut0pDi
+G5geYvlvSxp9bbR2s4ksZH28ncHqwgcZ0LvZo+dNvv0KNDu4z0rZqnZhYZD
64O+Oi30TkSi0twboGDYhxUFxzhq2J5v7/BY45OKJA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C9E+169fkob0f/j5fXQq+jYbeRyb/uW/cDLz5gE4j5D3p2tQczZ/EoHThqKs
4kRh9OL8sKyy3tYP+5mbPoEFz8CaS+RS1lxkFPoMOnfdYgBWftTj0AJWrXRq
fw4jm/yqISZW0fg8GbBmwVSe4gdF7t7rvsn33Bg2+kU/kLqrzK3CwVkeDYDB
t+Q9SHwI16WelDO3ZB5O41uxZnuWnKma1bk5ZYkqYYpp4W9eT7UqVqwLQ9it
IeWUOvylLrQ72wihuSN6x016YbKqsKXlqmv1/3kpJqHFVtzCVDPepD2EnBN6
0kQQohoOUFOVMROOjIjHW15tSDnbI6riHmfoQcTlsw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YtIWzyepv9pSOrqKx9R2lFF5Usf0bwnYf/R6h123QwMVihWtkq6MnhHuk6Sn
h+7IS1V3U4LzhGP8l5VuMrR5S5RYxGLkbcIB2pCJSozb1m8nTJHCfP3YbpyX
18I638NbPKJNDSlb+KL1u+/6NMupBcTmJo1T4y207PB/SLH34oo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
U6YBa3QIlBc0++XfAjlIAe0BJA5Ih4qDzEK2EQvtiNgJCgHDO/0mFlpH8Vo+
fG5OPiV8XhumgGCGsk/yme+rO7tXjYsU8uq45F++QTMdzmSnwSyPouu2b1a6
469jjClvEYYYBpIICVUzr+iGRDXKJxyYRqm3QR0UUo3WcpZ7vqzCcCR0NosP
e/vRM3sNY2BYTaxX0xzQEj06GA17QDg2xOkkFr1T615vMlUCvZJ0DjdcvOzw
1moymglO9PN0AZKZS5lVa2E4RSm6RXnPxkbvgnUOcjZV7O7DuI/8xMItl9kh
7rlsufgVtOlg4wuiyZYcWB6kY/2jnwwvFBnYmjELmBHGA8j7bSEeTuf+23zv
gK5/9qV3YoYEdlHntJcTbnX0sUihtfmLAoZBA955PrNRqbWWxBE4Y+NPC3Jz
tf1RyKX4pMa16+OffqMtS9h3svFjuP2YLK9gdy1pIKfd1wjA4z7gxElosIYb
ioCr84oDxsVvun3hmAYMYgdqNi3cJl0b


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nLSCKSdEl6FJaXjmTnzrEZ3ZWBtBTWBdn/Ph0pLzgg9DoW+K8sCfz7T593NX
EHYbPod517DL7W3OuzAHOZ1+e+OozAroIiGBQbU1M1t9xj17G1xm+AQLsszE
1ffJO2g2/v6m7PuVo0ASheRTJ9Tent1whP/Jw9lKkq9VCYi6rU0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Zc6mk+7oepwTePmRhl+3Ozitt8B8HWVIvO/AdXouXqAhyX3etbfeOn78JADj
VJcZhWS8h9NxmDK+ByUAcqMoEzgN5xxKHrW1SDXcvRUzRCYg+maORl4NfV8+
ARG+lLnURYRoXu6DptwoV4hvz+pKJPgN8Ra49UuuLeSdGuwUp2s=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28720)
`pragma protect data_block
2rPwCaN/EiGSe5ly8yvhwsSqElM0QWo5pwEcfmkPbkYxDhJtwB65mk166TAR
8psEM19PNCqOB6R65nGajtkb1Npwhr94tMop5BQXABB56sdA6ClVpDZDy28e
DQcd2co+2AlHT+OOzrUQlwFxQZzjg2DnEpDNoeHeaqYeCHa2mK5oDYqPSyMl
pdkK0uYvDNxOkKv/vuEG3UnPPgeC3sPbHv/2J9gaFngEDV4rqPU0YvjFer43
dtYL2cV9vSbRg98GQtQSf65YllOvX883RAGjAH9nHsfsCfhfrcPlvAh9EeED
ytvIWd4M5nbqUY6h1VaCupA+9viqbcx1mLvkv2mymAuhtNd0NhO/SDvTq3Mp
ex4QlsMZl1euUmSUFY3gCbrShU6avRWE6yPtESfa2ZOK1qqzc85q3hsg4LSx
xHbwWvmPe0ScgBTgGxtyKcR/aE9fquqHuxK3K88T8jQPHeGe1ee1lFryjVaC
nZQtyOdTR09UKKs+Zf85ndpSKAfvhcguDe8kT7a7+SFD74xRTL3z18wswmPa
KgbcVzKTN5tic2ztd3nOXcL0SFfeqzjWmx1fsOKm6sWLM96PnDaC9RrgwxPr
23jWZ83seGbFfeq9xgNvVVgUbwS+SQH4fIh6l1Jpmxt0ohq4WCUbAUVrcEA9
y2y53ByXsPWikX3U7xBKiw0cqx63GkpAF2y1I7Ola0mQvsESrHjleAZN13Wq
ZOe8XXhPeJjwkt9aI2ce6/vgfYSOxU+KgghX9vZj79nd4ySpY2sIreelPYBO
7r4h8zeWAYiMrn0nr2FIldbasi9W+HFvOq0DucLTWBSVzveepQZfH6UGHemI
aYrQK7jKO+5GW2BXrctOobCyXoja9H7LbVLj7P5Dp3xFEqri/in0z9Kns/YW
yFwYE3a+p6vvpr0KQRWKi0VCgxl3H+ZsVLYfKQ11AUamy5FyQVzJqpH8KlWa
QjjLOGT613cfDEmJh6esEyCIxy16wdyyz3Gk5Vj1Ai0wvF8j8U54Q2J/g5PL
b0CJ9BmyOl2MQP1hWFU69vX3NmJbLxvZiNR0MPKAwx80zUqJxjg/WzPlgURc
2WHO/vuOCf2KugwTHanEdx5VzZRe9DEbLBodcFxH2gdRUTb7pLLu6zjZAKFm
8wGVUIHn29VPR7xy7yODbyRelIH7agPTHYuilC+zb7Oo8YFSsvQjohRCV2IQ
RVBsQ/f6uRxeHxVRkU1V6lV2t4gdWJlvj0OhtUWCrnMVt/pJLQK62rLh1FRC
TKvhbnNnYekcfeWUhwTSwTKJqXi2LEhSenTkXzJe9WqVRCPiS9pGeD7OUSyI
3VacNWm7MEJk0KKlKLT4sjJcjbejzzXigo4Hob/RB/1m1t/t5uh99wMlWEpV
rXxk4AZqfcR1SuLQdFEsL+gPiJ5gEh2J2AH1DcMUHwGE/jurOC4AV09JFqHH
YW11GY9J2u5Ugu1A6kb6lFreRwhIyORJ96wHcE6N0ZsqrY/NTq0HZeA+Z1nT
eoUwPIpEMscnPFAjjQ+STwStr8Vl54Gia+myCRzcUHE+idtcvYOI9PUyID4+
jAMjw2WiPm4q05D+CsN+b88/0tjVVpmdlEQW7YvOkPuvv+yQcJyYKSxU1Ega
9KLKWrUkr8WSPkGLJhWveZw3TdUUjHTx1Mlr3CwB322xvG1fGKJ3XM2wDu9T
/RgUVyTYsB0HAtoQNx9vYb5VrqVg2G1A6WPi6bla2gm7n2Wputl9+FmpQ7y8
4B7YKr2sHjzc0YQf7Rwtw9YN0wbV/0/ctu+0S51UH86y1KtaKlgCLpOZMgBm
MomzvQKwyzYibHDYxn9DCD49SOGthACnhQjzpvxXDvxTKVl5dn158cv0nzVT
iLRxEqR3hSY3deabxThUxcI/lHtcgiMibxKNiBhJ3LaE+uTghFAuxqXCJCaW
P0DVWqreNm62PXnvtDIs6+WtuJyH5WvhJ8BbioB/o3Y1g/hSJuxRdmij6qCJ
rEJ8rnIZS+qOt3DalIRRV9qCCjYA0RJvx3JOc3PlTnepjF3Zd5zgVGM6OFzI
0ihG8QdW4ZRska3tZbtY9eVnT4/ulKuOdsRhJY+HHIgtra1MFIcksh88kNAJ
XDwxaaHWwquJ0kJe5POPkfsC+CP9ikRhZEJmwjx54gF+uf3SDkBSsYFyZi0X
Cu5RFfGAXgK/jvTU34FbNGIhsRsLD9Wt+1ZtBZYwbm/IaTzu8tTUldQOcopb
NV4OWIwKnRzG/BdgH/fQGBWzZI0XnUHNIQmR1oHE0pf82NOS2VvQwAx2xvEF
gzkk+79TG+jFQOfXm6vtIDtPBnsWF9cyGpKyWvxtKNevrVJaqETx09xvtKGr
MSdT68lqGoURSTphQlenZR90SAfehucgT2Im9gsMjJxq2Tfi3RiyzPmhdC1z
2D5rXhDeVOYYjx0WqAkb5KgLKYnXdHNYw/J/hvCKDB+fP8BXNx66CLugyGs7
LMdupqgtTZ1/z3TQ7+XdHCfjkaP3TGV9HGSEX5Oq0a+UOej4Xf0N7hJfmUWZ
v6kGhhqEw7SVzVRh9zWZOnZdLFrB9rULpJUsZbP0SrVrx/Y+7Y2AWWHUCeuW
ZL5PJfVfXdWw/ifEWQEbLldln3FrbpwvlhDYn4DAQsPxQwBAQew4BBeE/2U1
f6eFV00vkzd9zjy2fvdgTcVP0tq2u2svdOByKpUulezH230a2/olO2jkrV+g
ZvDjXUIExXr/LAPETJKfjOReOqlcfBdBSAizNDgNGdJdzAWcgxHJrrAwnMYw
a9B1ybBRbWFR2iA0AbVFLDobpLBp2fiki/hSgwdv42NNBvBdU/ICPTZJEwce
YWRq7jOy5mfZsOw3X38tVrY8ToB6T5J/JZrLRz8JJlU86ljTj1RRfjldRz1K
FcqgJa0YBdPR25Cr0O2NWx/KUxFACGEH0mlhSup/RIzHwRIhUMkpW2LQpNpk
5Zxm8N7FhNVshHuUznSy4KomffFmSTXx7Ua5LMLpoQVsWPaKXk5Q/vU7CQ5d
xdk2+I5YUGr88GC9wZz4Y0dE/ttTyuBN331Ibm4RfUIvtV6FbQ3s+KwSReGc
ljcBniRiM9tU33yBk840ylv0XwKdZN31U1rSUcU+K0LkfYvRR5eW3sQwQr4S
wp0EFJH544NkGlQdVnS4p/Y35+MS4utmltAt/cQLLRNAhutBoascuYkAaUmT
hNchpRzmBjmMmXK+5t6BS00xXopQdI3t9c+FXfBMM3TA6uSkKWPeLKNmgVdr
ojHwCzf9OnZ3k0MMNqOthAXq/ke+X+KZ26XNoMJ2RKmnkGI+afN1RjT3W/C7
LE6h0glAirhCLSW7cq8ycrjYSz34QVak2apWlBkulNNdg50072NE8jKeQppE
nMU6u4e7AN+Dgwbx8uC9nkWHaJuN0hfe2hUnRWSnuSsDwmpDe+AL1LIvbqsD
3hpuyUvE0roSxEAAr49gFDvH0h9pVOL8INox6ilxYXzQtpA6Dfb+pMw+6B1y
dTvEpSMWyg6dYR2tOjQKpf4GXTLL1kwthxB+bae1VG1IYu4XFeq0NTF3QaDv
FxfPmDMEmsJ+p2zkqZ9IcmR4O5P30WS4uUOOFTnO/JiWfN+CmqfMEs8wmvi8
oBetz6fw/GjavsFXGqWaTddeZzWrXzaAZUW9r4O4i9PfGPxovpO8eb4/ql6H
VqWJ3w2mHKhCe5MJ1N52FfdV4GGwIubL6of7XX/f7AL6XnD0c/pI4gZ130lO
GokKgJxMBiLtwHzW3SVlWdeqiLze1Ywd3JCs9AhWxn363iNDS3laXCLcwuN9
ZiDR8qqHckCheC/9ddTQ5AgHB5Z1S6SXz6Pm9zael9iPmWDUwF5ZAAJyQaO7
n2jRwikqERbdFzdvZwCatTefbo0g/cfDVGpwhVQiJU8uH2xHLEiDYMsXGDj3
AkVJPlBtdjFobVqbvzO11Lj95ciXs9b2d1fzHxeH3v2ewzft43AfLq8RWp9z
w9/ZWdUZnfk2Poj7oEEngI1KykV9cXEe2/ET65W+wgVajty8Ak8TAH+qM2Za
8a81BiE4wBMHuL8mGy7UJvzzKCv8kJjv0XXggyz2vT5qeJn69XV5IPufgCA5
PaFqSQ0COW+9eMUnMiwS4OsFBekFEyWgc+aGqWgEaDTKKf9X2GDpRO35zx3d
opICH+8dIztzU8bJV04ynLS18C4mzfR9Z59M1Rr0AKexljm2McHI/sb6nkbf
7JnRzl412oMWfXVWqEOYcdfjbrpmZcM9UCz5eRu3o082pDfkI5xWCbTpis0Q
tekrB88Z5M8Y5+v091eTgjTOxFiJ3PLbcCnnxHpQQZAl1c6+hW3kpYgTi9l4
G2DLUu21aeZZ4e6yMnjHOjlokBPbC0NGlQ5qbW0ZJuoF94l9k26esonhboGh
+sHnEskZ/fllG9QAWYpbneD3YS051CIDQUKWFUr18l/XB4MhLuasxX5/N/TV
n7IhCFHSaX5Ae9WsiPLtSR1UqCW0VH3VpjoRmeW90I+6f0bAlWh78pEyyjep
rlN6yGFBMLdQADwgZavM7fRKs1n3FiC3KJ0JR+ouDXXqgNgPxI/kIrfUVh1s
AUPm+FzKhV/g6Gr9tLa31MmCPbQp2T276+FJPLsRRo0PobZJH5CwyTAPTnG2
VAaZfCVVOPgPnYK27Qs6rAe9fr/F3ivzQny70MqDbiPexx1vvlvbf2d1b+DB
qTRACJQPv83EnXBohOZOrw5Mt2DirzqZdMLqUyoKvtS9pFaidlyn2Ay2M54k
9kgMlUf/ddKcshca5eRG22cRVMAR5NyzKEaiYxDjXzsaBH6IjhFgp19z30jQ
yKLZ9WQBt0ANUMLKmeB/TAD8H1uel4+kZCnNsdNCuAy19hTKNWlEjXUF+e7c
UZXvbiWpyt8uvdOMJv6yUXAx6rbQ09Sh7EJ5iKsratj8GwyIpvkuWhcTuusQ
cHnNiKjPqEYaVDQt3VOVxfJ8sUF9x363+dAngc65l9BbEx8jTx/MvdSxa4ZF
rLKmcGKuoH24gpzlObTMjEFKxgv8mj/GVGaj9gg03voa2RVGRku1s/Uxv+i6
hcwxh3QIZH+VeclBDvGqfQQZR9QZv9nhBhiJHOgiEywHFGzaP71yLHVubNaa
3gcpAatFH14yEBIkVarjSJy+If6l3JCRY/QgjkhBf59zZVzlFD1wRzm8j5Ly
wSHfGsCtxDvnWwdFV5GqWgbt08lvS+WyyYxG/Hmt76F/A24bawfXGQ0/ozMr
TEjdMv8MHTla3f+N6pYeLnGqQEaMvAjRZJB220sBXuZlK8MFnp07/pVNZF4B
fARfblFL3uqGyrliH/58Ro/Cbyj+8tuyJh8L1ORS86bdNswJrMzvwGp/gU2o
hTWdisZBF71Gph7UKJWoI4wxrNGr5rhMphw5FvLkEz2Hh7SMdl8t2x7zcUM4
PqaZFbNZzs1LQ1nh61tP4KTz3VbtaLaRgqfOoZUJsTcSpUc+4YDR4b+dJ1ee
4V2DwKYKFRbeGy/NuYeNL+OLAEqBEPsFIj6Ro2COMcLxkrPEZQ6hxP1KXVjV
LgJ3qyNwkkMy9A5Q76jvfPIEix8Dvh4Ctz/+HONYHkMHLetQaW5L0QQ/xhpH
IRKq1JdoYuNJLG2OHMnD17NpMAcIDUIH9hCMunuvZ2yYQ83PbsBB0AlkjQkd
PxBykrk2Ph9R5Ufp1NL6nrZbEXnlXLD9/NIxneFJYqabmzpfu7+csU3e7U+z
FmYm2MqWFMWl4fH3a8ypTC0PorPH01GwoB1tfpBDDb7vwZ2af6sEJUiV/A2k
9CavaLcvxLuFIAYt1Fdt4aBBN3EqMPtWEBetZoauyAqflhcgjCqDYkD3/A2j
QrauWhfg9+lzcpaVAqOUlCcQh8uLNVz36aysb5G+Tf7IYDXK86oQVdN/EJ0G
MRTkCFGRzZPtfuRamAambp1NuZjTxe4OLYvZsxZ1oFzyyuAtv8LNiat19yTQ
71xZzfgJnkNIBP75Giz6+MecGpmZTz5RrfsgHEflv7Qwx0annDCEU9Lmt3Bj
Jp1t+MgHFUXoSXK9l8LshSx3kOuRpn+5GYY80qxrfYI1XkxKLCI/CPtwlPy0
Sf0EsTy70rFcDFRzIJ4BcJ4p8rKKCrTAR8/5rT2gYta59LvmH7HcwanciEOj
U/9aqCw4BDJDFnaYbdfLrDIFkW1ADNzKuWNUGUFsqVbEDLhuJ69sycwx4Tgc
Mu1T9lUvccBZMOO9ALynDIfp/s/Z5/rmwGemxUmdS8NnWZK6qbF4/DMUr42X
4s8agZbUSc287vRySdlUaxDVlvShBzJjE5qNi6BMGc7X7RiKZ3U6+UaqUUA2
H/viVto7pFKJQUU17v4sGYwGqQWv4zMxzvkrfZggJTdf4ps3nJkmtlGR13nc
0iOoBkEfx+iennpmAU7o8fZRwg4BtXF6Us7hCT3I0ecmX0Ys+AKzHQkhplYw
pcx9rsC7BbvCNIj/WhyzHJPIQwOysVIdJulkc2jRi4KYGGnXZykA79gTPfzk
SIcIa0T6FPX6/JN6v1Ah/VaF1kjLPmaYA1kpII/vnXuwqvxwFMvcybC4jUtc
je4shyQtAEfIN8Qn+oRo2ZNssYIQM0tXvkeSG7At3uUK3W40B8I2TfyZIjxO
9igQOj0ROslcfp5j+oBIpqd5TRhLugcp2aHk1HUlMPQ9KczFL1EYV9McbzSW
dW6lgaUK5PZ5pievBDKRQkZUeI3GJyJAYAQrtsPZl8xDgrtyrEMYhND+OK0E
TE0fS2njNBBBKlomVZmTmyU4cB6Xs/5BgauoFZaydz0F95blveKN2AwWuVFu
VPGM5qmGkhibLJMGBhF9xU8ZhBxIZMpaxS0btVhvfbmZEqiihclfpIIz85ua
QIWppzTx+cJvd9A8zo+awPhgidoH8JFdpyrqs8JSuZpmM1+pwDiZO97RMvz0
fn9PkdX01CLMw9j6lHW/5x4VcD7SVXMdYujtS4j4HHPLFNhIzl/qgOEUg7Nv
+AhiIFfjBGNegqbcaP3kIplh4yL4UD9GGY2l1jA73VdnIA9q9FOsAZwmtnQ7
uDFcrBfUZs0xQSMMvkOPDK15GASIX5I4sPZTUjPEWH+vBGl/LQ/F7vIZOsgq
b6xv49soLp6KFVDOV0UDtFI1VQpx7GOl6xuGsVhsUNPzsqdib72iKtDmvXdY
siY1dQyeKFZf7MmXw0qqeXrnpBSu5d6mpDLm7F9jNfkEkIKRsgfjfXlyZl2n
Py2t60FG00R8tUgaERD3zO0yTitEDSAGSPPxLlmNcMQiwnajpypTKarycWqO
NS7KKwm1/811WJcAdiiEes5CSf+uNfGGPPnLGYPnyWcWd9FGQjcZqmsopoud
uWQmwn2CYFMcKBx73+Yx1v6+uelq847H8VAlHbpIEd3lah/nlGsvBAcIwUR0
GfkJtY5aj0++qQFfA5NxuYMTTOd8MzUwYpWLnLYmF4e8Ljl5JtiI9/gWuWod
1BEWHUDy+lxC6u15UhcX6U5b428BgOgXJbMC9xf2wi1ZfI/MirifPf7ZJhWC
b6B2zNxBrA18BlIbve08q6Jp+76c0gfsiFgvxShMJaSA3MUKiIr8rCW99AYv
SiiHW0S/E3PaSNxRPp3JCgcau+B38B07HsOnrLlrN9HbGx64ujdFnMWeke8P
A7nDV0tlx05gfvcvibXkKwQc/gH/W0w/wB05nki/XO8R0h4dQ/c/GDmzFYkP
zLdIfCvBl6a7/qRFMhWF2Q/+rOsLo12MdpTeOIIqNOA3G+SGIk1nIGeiKKDn
bEO7hZgW15f71YiQ03Gl4rnLfI9WAN3/A5fX3DD8hEzmetjfKRlQhAQz6y7p
0tvwWHWdmkXhjg8F8VUhB1TDr3AQKkNbtqYTAxlA3y9IPJEFsbU5ZsbMmkLU
U8viThH5Oj316apWBRTCk9ojuBTRD8XkUBdd0AiemvI1mFHv8Bb2L/VgdWyJ
9sRtM4AFW7m+3XjkgTImN8wkeDp32fe6ivCsetkoBCq+vDI8UxuNO71VOUc1
z3heqQVC7sRuFrv6PrA9ST5nSZtCcoXXKRdtj6Ovwkn63pLP96UgCegsrYlT
zW7NEzenzJi8OAgk15MypZMgfvskRhj9b+nSfV4GhT4dUulTgA+B/IU2bhYf
sDMzQrQQBCSgBOMxMeyJowmgZVAxWUs8T3srKA1mXpj+/UI3ilaDj8BvIqxf
kjmGqBITid9d8ahs5tVK2QT/hoFUeCnB0EWZfxqlzhazrc5avCnDVDyoWzHJ
9ZOSzBDCNPgBAv3sRSrfno3qiHAKGQyp4R4zf0aUgHYxxgfmrTAuBPpYbYw+
H2bI3DPZVKelRZNn3hmCKooU3sEwU1m7EEJfKvnOF80sTKE9wbrLC0tvn5Q7
v9fJntJNw9wZtr0zr9hiVSg7qDk4TpqBLIYM0NCV57UAS5cLoLdIVv9X4lP4
F74i8ljSfQ2SGGcpgepBvh5Qomi30tIRjZZXZ9c2QJ0YYI3iYRqdTsJ2Cku1
KF1CawOH2nAYBzp/rqQnhSnudfPwOJyW7v0UZwHGqJR0DOWTDncYaA2/3X+V
OlDUHUwwQBwEHeepzUj5mcLKYOrJ67SAxG40jZBLNheIMeFF2ObkfnkJ5SWb
vJDHEraKwNkGNbPDTvKA9ajosF8fO5suEoTAd6fpWV2ExOSF7IeAPUlWRZoX
rSeAv4Z1intiSDaysD9QHqGAfRg889vpu75dyVaCeug6MCB1Vk2rHSF6Wip+
Kse3/02nPMJfvXcvCyqO+sfnyCN4YGU3g94Sk5/nh1xngrkhu+DNvR3z6NzG
b1rpMEAmVnsHiqL0E0zDB+GEBz9W+BjasA/ybtv2KdSyCGypnpxQytj8Rg7Z
uE5QFjnNWjVTDDXvvmhWHgBTqTJzUG5Weo7e7lV4s+tGQKd7T9Ef7HFeXIcD
ryRpe4oUuUBBLadSesq/loeZl3nfy2gKTn5V6oj7WVgHw7tGlP9u4qJLjM+L
crKt3CvwRXNNGQd2+F0f7okm6hzU4MhGPQ84dEwoQi4qZQn8PUvAyX7f5oAB
meZA93mv/tkDekbGuHESoZRcdhgOu75cmw4zlSdMQDsUyes8i0OFvN0OWtcb
lyhRlZzzACszfqdDiwYWIb+9JZYf2+PA6RSh9f/syelsxqY6NmB3w3HZb0an
tHTlvhqY5X0TGCFR9nuob9ZCG9/8luNEf6ziv2KlUezG13kZnHRMsokkJp8l
iZRAzF3TR8Hmevz5emUIvX6uNm6NKImsz0rZqzwFcxazh1WUUXwv+YFlcymd
0bFzt4KtwzRCJOPbz8Zk+QY8kWOpdJySPTUbc6cA+fw2puNRBd7fxeLWqbHr
CHz/GKvNv8y6lbBHp8Yg0tfYddGtTU8473CgSM0qrAKqYzdt6m7pdALQbZX/
sWsHazW+qqquHA1zEs2HRcs3+4S5SXIXGPKXwjG/IZwq2CBMQl9V1EZ6pMEO
JhaxhLhr0MBwaVACaNz8Y5EHVpuOoTOXesWS2MPsAi41N6KEmtplf39x70sE
0nv0cOig+XhnKKrGF2IE2S0MN49CDQWhvLH0sN14WBrRIwz3Pf76sr3JdpVu
mdeSgpDCMroHgW92/HWPpFYFZaZUDbGHEqSaayzpmHVHOlH6oowagBfnjhUs
ZEdnSJsEwHiP94PlGCcVscYqFEGEhzXl47kpFthwIQxFotZBDvO/2OynwxFj
bIFeoUZds2AKODtHtjXjJ11B/VqSUIyZFRmv1QItyRy2/Bk4/fPQcIE8oFaT
mfKyJfx0/Ro9PAGzS8FgcMib41HKAyTWjwIZ+U96QFD4W2PCiK6h7c4Z+FH5
/ZnnUiF6Ir3uEy1jaMs3uG0ivsTcpt7mY7JOZPzhtAX6AnqB+OYUwcrg68I8
yfwFtFgvJSWV5S5soP+zGQe4mnElsZcm1GsNWKre4cFQJh1gth8YvvU2JRYK
b0aNp1BlEOH0IbDjU5PrXzAhqPwnDxNsDASbQcxEd02Yv/8oKIPtsfxnXBql
kVfOUwf/2LfvRKsk16leeUz/v2+K2W7p3qKGIL6s10FKABIgOJSjvIQyMeBR
eB2Pl0xHax6Nl4JKWA2VCzAdnQ55Fj3qeVx0uc1YiSbmOvXwWR8S0UopBsh5
O3a9mVcGdt2riF2IyI4Q8hVAdx/0Ao1TayVqV+UzmuyU+Rj/XyB4Ek2Qu4q2
qmrQFu4kLTbsJmhTOC9jTmYfjqu7jI5X6ku1tTxeZdLf7loFf/HrfvDaWMgD
z0fa+utzSbq7fwsm0mcyyAH1Ilospsg/OtDRx+bBYxjfy3L3EDFitF/dnhBf
Ej0iJc9OgR1z9Nvr7DM1GPzVtNIGfdwdsGpZgnRo9y1NhmXbnCTMsZT0r4gA
IpwHs4kHg7GdRbJNXolMx3n974IMYCm4j3BZUf8bYRnKlruh7J7X1LfIJMi3
nnCewpYAKi6uhVAyG/WcD7qfe6Rsr4WTyLb//tuaX0iSVGk/ilM91DcamgNy
eC5rxfUrT2qADrARZ6JEXvpeHeL7ktZldRVBhrYHlJpj6AP74DdCoFu4854S
2211Mslx+x0CWM30f/cW8lmit69zUxAr20c/OoqdOQMuyfHBLSESiibe6BtE
IHlvFnicSC/UDAVo9vwtdT24qfqsk/Rlm73q4OL9d1iAc1cZ6ZXiokY6GXLm
PaD9BMx3Gcuvo82uhwzNmJ+C7zjf9x2eu6l5eLE2BZkx3zeRnDEFDx9dsTjB
7C4hE594u14x32Ah2SaJ2pW1ZlrAjCa9Azc2zoLujApwB72yEQLfQZ87s7vZ
7H/qqH/zhDlNxq8u/HgILzxgHjVCx9oO59sznS0hk7PxUxvKbICBlimn36f8
I5bBBc1H1QONDtvB2zra5Jr+X9mpCmo8aNTW+ogk7ZfNsEiT8xkk9ONWBNYd
epkq3Ore5zyDhxImnr1UNvD6fwzjQqmfUgXUCCc/LLTVopb/7lsfndN8hGyM
wCki9oBuZ11c2hCaTI8HXYrkN0lbMhDTOijY2RDGTULP4ELqnFU+xJvdVM4Y
HrBrNg6MN1uTpEFIUa1fVOOgBID7+ZQGeEF9aCbciaMlPzgJKc/Ie+hkN5NZ
FYK4ATzxHpdsAhKiuVApp/fX1CHWpoCHyA30Ga16NyKBdJnb+hbsjWm8MdKg
hl7kneZQSvsrN7mgtfLpakbcbM+OBHlT4cgIcLmI4rEqh1a2AGk0slcd8rnx
dPN83MKsWlr52iJXkt2o6XE8Yg0srACgW+EFeGSDZnpXcYmGAXYOA30gMQZA
o0pW60N8oaQvWjYVgW9oAGwWPr3r0GT6AHvEyfbgKEjbXJU3nAnZFK6UR0CY
FoVKf+Q68128OKiI4mz0KdjBqRmJkhx2Hb08tgumzUiidryxN3ZaxYxalpEk
BEYXLRnqv+kPYw2BGLXBTU6mvWu1Bvzxpfozj9WkpANbF7A8p1YOahqggp4H
h6Ho2Tcj9XPC4G1ZUTCEx5sLZ1x+WcWhXh+wk/uw2Lj5koRqIuwmy6ZN+wTI
G/B9YSXGyrLegieBA0qd+ddPDItlmu9tfNps/h3llYBM9UWsGMlCE6EXNcB/
ghgA3RBELWlNrBZdAa/sYQM5N4OR2NxdkpA1sOepaoiiOzJhTxbTKdG7erK/
7+Bp9bvhgiQSSEsyYdMB6XtHPIKbFx/NjSoR2hZqV5OapvL4QJfKQtQkQcNh
z7+dW/0DHwLgaAeoLu780/WeGhFwk9LGVipy7pqJOcxMdrlkTm4/S8cbIwNn
UmmW0JduO+kSSeGIsqwiGfdpaxM06gCc9Q2ySrnRUQ44gq7opIJfazLf6NQ9
iYwm2GV8bJwMhtNUWS6ThP+stQN8dQhEThMW8Gsl65CUkBCIPQoXAp4Euedg
25Kho7Cf+xJQr24Tz5tLB7d0QzFxrT1/ZsNI2a5LVv84PYU0F0zTsSCaqD4A
woryrgN6mMiQ8bYOnyi/S6+PTmg0zbkD/mh+IqbyebIllfwqdB8xfLXVXLsz
cGTHHX8BPFfS0Tg6dGZo7wFtVmN1MIWa5FWAGmACmt2ihI4r5PbXxm6qEjTz
INiMKom0PNYEOUXPHd/dp4GESi0ESWr23SnpPvxInXzPYh+/rGQrnDkvk84c
0jVTzSDDoACo+QvEfPEj+3AZN0yf40UBEvVVJtDLDrzNK+IV5XgANcHgbokt
NS29PuaLcD/URFPz5Z83FoOppr1AAsOxR/eIcgaMwI4STZ3adEBAp/erHgSm
k7Vx8AhluGZnGlDCJF0KYsnkglGF9bSaG5QqeILEl/gVLb9/3cERSqCM1Qpo
hFJQvKgoSWxOgbnni+/JWl0JxQ24LfuCXgQr+88EVg7wQgFol4kpz+j1kdR3
qArHTZdZfsKr1K6O19q1mMTR1zdZ3xo0LTZu27+Gx9/GC7MEMoA1EdBvetzR
62JKFDPaTnuZwsChrDsHFMyCNXAni39Hx+iVGcJcgBFBPEaJe6Rz+MUeaT9X
/azk0wzZvN86luImnxLSOC4tCc8tXnUbs1EhD2ncp7SKMtvMfYm6TkisIDk/
ngrqPcFrQq3wTIli+tivBgbCci3IgcFoVqtQWr6pNkwTL3MdJUId9mDYliU0
qtZLqXFvOqEKXA1Da9R0mKIBQBflpJs8VbmpKZIV7SEIi2vS4PRE3gyNKhWG
mrunjv073/BVZdsR/WoL1gGagdh5mqgZ97mSQyvMsGvvhMWSkdhIp/9+YQFz
irY6oeED3HaPEdJqddbqeh66i5e7QZ7ZsqvWfPRkHlohkNei9S48HngbNHCE
ShKDtaD1rsIV/GYp9HOIjYqjVUSwlzzPNgUSWHZ+y4AEhHKhIdBcaQMvwVaL
vjHgmma3YuxI8GCsZtfISxiAJhCUS2uUrnDIBZe5tLNzvHvyd3O9Np9iqUBz
3G8a5smDPEqctw/R3FrtLjF/UAALu/MH7M70MU4NWxFniG90k1c40JpoWFZ/
kN0gp4QcuriQxQ1CLEAIJT7XWY8iaGYFrjGxPTnIm814tysvo564BMGLqKni
s4wi9z1OJsNvvafxeE/6IIYLJVcggetcNo614CoqllHC4nvSOlFFFVqlO+3w
FYX6pUM/klMUYBNF1dC0dJN0tYTUbqio7shTliZ0O4jaxXvcRygNq/RnFPah
MxcIYiLBgCK17oIq5w2WShkapWniwJQkAc/ZUM27UGMgnveTwKq6UQfJZSoe
TUQIQZGGDHU3hTyDw/xWFc2J7X0vRT9KF1TdX2LcyYcW2eTxMYjfhMvb0DsN
OFvBIhUOCA/bu7VC5Gb644xUSvMJuZV4LW0FxRY0s3e6eTkp1BHLXMVprPNw
QJEXEe+uq+uHQ5zpeIe72dN/J+L2f+fg8FSw1sLECQb37pV5W+TtZwqVTQ7s
QDo4KHngiEe7cnl6mi3u8AZvCiLTbeb5yBwPznLbpbTrdQdaXp2rQFrmlzXV
+UMBlNGGBiBAwT0FUuKAYqhHCKi7yhP+iUQFksnlAWRuSmNkCjRcOhRo5vRc
oTYeE+1M4MCqwolspElxlThAyHORVjGhkfL6MY4eyvTi3Qv3pK6vpCnhnvtY
vxILCLP4Ok34BRSDWrangZa2lgMUf3gXL1pcyoaY8m/fNAloqnjFVJF4mgD1
5AL/TSMB7wD5K+jZhr7r/UJ+DGMWUqx1Rzek1jhvyLCe2YrNjue+oLMAnzQl
QrvX7SIdQoVey5wqKa8rTaOKkBC5wWMA0ApSLxESnWCA05vRVfcIyxpAHnIN
7lJ0gVxH6oe/F6urohzowxwZhrkPCsDTn6H1bVm/k7BVtmEltscQ3OHZqVFT
8yjREPFu4Ttmzl+b6B1UqsS0k/6w5BfAHYeQDlXXkFq7ecq84M/YLvInOqsa
x8vhWSRWvRFWPQl1ptnFWkPXILfbVgapHMRMogWx+DP3UGhMEa21xJmRkuvr
gQd8Q6vcCNKdPrIZJD7KH3FH3CtooD24SjqXsd/IcSq4RZQX+d67vgKu7z1j
xMkW1dM6vd3BPjK/YdYhOFO9wtgjil6v0ouwD0kLBIiqqmdgq7mbaZSXfdFY
p2VlzdhLaFCb1+y9f8ABUgmTNkYNE0K3xRODRlvJtp72Cq1EkMtOqY3wzSFq
wQX2WJXTiKknKzicBlcETqBU5XLga371+hQtvLmfcTcMQW5n9hHI5TowLDgC
dm5/PUUciw2TNtc6KXa4tstQGC7VkCoqY9cT6hVo6Lc3rSdJppPnFYDP0e0b
sdaHLlxWS7nSL4gUiebL39zIXocHKvvwmbJw9alB13l75Pf5rPCkhedaLbid
mD/aHaUtnh1ucn/qbpw5EBVRwuAG4y3Jv3B1k/RVSgyvmmusfnES0ocGKgWc
GST7uayiSJk53SVAB4tSDpehXuZ4zdKVD/QD+MjhzvyH8M5PGE2qy5iB+TSE
EuTxv4IMJslCRHJLKnqFuQhZWHpFYqgSg3xYADRIKJx8laC4Y1QTmlBhnKwY
UUY5ClUVk96rdGVGP6AZvUWAVOq6B9ayce9jJdc4Caq61kyrxjtB6+iV354m
TDpeUDnN1dzm7Zp3K7bvduxf7Sge6YL0nHp8EawTkJMyjk+SK5Q1zNZSVu50
p6mmxWKhaRXpd4RIHDEZk6wBVCwrgkrgEbP9VfH/BoXplpwbYHvZyh2fssAz
wsD/PHCs0KQHIane4MZzw19bVOIbur6zadwo8lf+7vwsrCBk7zUP1KrVwRTF
40nGAR55cZ81d5wU5FnAVTWp8k/1L1AYznBwRL/2FIy91oPLpMjsIuW60S9j
uZ61aWkSkGf2bYZmg3e1mDVgY2tyyqI8QzLurqxla/XG6zEEx/jFS+KLb4P6
T2oYA1aY/fUkNH823hTZhPLEbp35iU06g5wjYmo9uuIrvZbWvA0qsWDZQrEv
UY7RegIy25CYWMh0MRHLHrYxH6SpgkleaFXnJYpcVPM+tV5FL59zkJ6fYDCb
xvHfURkWDIrihnKHJwwpDSCDQVGPz9DLY1I5HVOFO8dvcRDO8qiuKLXtUGf6
B9gatR9khZ7aKaL0eYy7GBQRr6CqDc7BBR6ZXYeUXKR6I+yFB6Xp4kdhmSdn
15mvyWF64vPTdY/cLvjXgiY9YE6Gk46xNBm/Z+8slVfPBUNiY43EEppoWRju
4ZP0JccuabIxtpOF7BvpknALJNnBDjZ5azQeIpQOre3k0u7J+XnaNM6tRnBp
d713GamGIlYlUu01Z7MtY8YKn83ffoBRrGHTjTxpkcoPo4QXL8cgvPIcRA7r
k36NjH+p0WLv15HbZhPW5MMhPYWm9lvII6r7AK1kS+ONviQegd4u3lkVNPKx
0uhOiusbahCroVBGDb1Gl/N16C2tIakD3qnrP9n6HHus3gN2gTkrUPUPsW4i
E+pUcYmLO9ieRT8EvhgkHJ2B3nXm4IfTcYKcKGt6OY+rhmHmDz4gIPoZKYD9
vlc9jr+e7GsZ+0Q7lBv2P5DzeYAR702TY0EiZK2Dy9r++15i/xZvc9PM57M3
dtyP/ygMgIIx6JcTqD5QhTwhx765nPj0nw46Igfr8y+KN/iLzGHr3TrG4Z9G
Jdaa6/sWzQi9fRCU2dgpbUe7IyWsExZtRzpPZpIP3iI9RqTogdINsLyd4wwW
9nPwpo9kNYaNnTWflS+x5kZdOB7s7XHPp1+UDLW18qpUQYdD3yWZTqSYQ6un
u6h79yq8xrBE4yZP9uQ1jcn1yw9bt7mGJe1VNkWGvHryHVeJ687HoUCSpzHV
QQ922GrIF9X8UM3JIttwPt+UgI7qzgHPYu3EjClqUEAnODPjNDHcKqPljXmL
z5a+6X4b7BneadqGgMJI4caGQmGqYHEcNxH77YwN81vAQFT+vOQvGg0oViCU
D8CZDAxwvC7ttxz0h24szdoit6cSl3Fz3ueJZygUbIGd7cz4XSjyeIYumy2j
4PKlTlLEwQ/gDtEz8Qei3DCNGvx4ku2JDKEL2UjS7ALah2AHap4P5WeFLN4I
UTwFPfg4FscTAsiWrHK8y2tKHG/pUkASpTS8AtFyjfOTctyOCTKAci5iYQT8
DCpEFHRIoCur7QlFYXtl5zLD2To5K7w3LDYeGO2hD1Uq2igbQlRUoYKn3iYU
XWh9AMTlxy7TmqtvzXm535I7cyMJWksANqCntMhoVmI9ZfTl1xQAAODyQWnc
I7EY0Sl9xX0lYh+DnG1oX1zzceTYc7xKfqTq8pp6Ir1rfqIvCVUv1Uj2KqJY
V3IjvpGCoEKlttzIJSf5M7crhh2zeeValdid7tm3NzaqI3Ork0lls0WsX9X+
FBsSnCpD+bFyt0g0THTM/VsTkQwD1TJDfHvqOpeUOGKDGpMdU65iy1MJtL+p
yKOXNkSMINuKFo8Rp8Mp0ILcc6ORnpTRIrdMqiYzQC2VsnXOgzWmJ3ieN6dP
bNwLWZfgmB3WmLhNeOrSg+26K0KspbNEKgCyDRoJci8MdEsPM935qaNZLyNd
ZwggZLIVKxPy/nn63T2KvR/JFHnZPM/wQAY7pe7rBOKGQNeCoP5UqF7DqSF0
il+bDoLCyVObJJcC3NyU2ZF5dSDZgfWobBmky8tTY1qv2bonfD6DttjDWD/R
JcogM0ubTFULgBu78xe15wwb50hneUTIAa5QRJg2BAOESQPQvjzzShY/2zVB
I0fVM73sq+pjZgGW/cVwAwsSUsaigu4YJ6I00tETII/cDhMY6B9i+xFQZ9w3
jlBsU92XaInTAWPUd7FSZmXPzU1fmEqL4TGt6l1GwNOQI1v1S7oz3zH1sp7B
VOlsYgQo/OgFxzO8aLZrp2qSpBIWbJbAactaWDPFYZx0Yf2b/+mzydO2ZaXy
N8IdUzVV4rkpng2ZO2mDHUCh9IYL5+WVe2KqVBW2rBj2WkhVMo8o9i8wdxPP
iFSNPICB9qwTbsdXKSi1zekq+BQ7D24969kBNQBbI5ix8+/Sk2HysU9+ZKT2
y14FxUjXByQhS1SWKqwnXcyOWD9th0Nr0FIf6huNB3q59tErD3Q6OD+xEVrt
rusObdc4MDcpqwKP3GYfnx0jikG4rkWMGm8iVuk2+Y3sl3mUwA9w7+qdECah
1tDoxvA1YLbXi5eY4WUm8xP/MUwiMm+DbkTHp2zAOznk43PE2MTsKEF2YzYg
PzxKANJEIAWmnF6EzGyc/QIm0TSnv2NdOKCSOzvBbxDeukTAkfpg0S6KIbCL
2JTFgkmLScSz24ARvRHX+/fu8LZNn+jGg/rAvhC+dfrN0KmyMt3Cno7RS2zw
lT+gZxnZFBgmDIFL0wzELSQW5YNYleKwcbAIGzR044MjrZTMF7CJRhN4USAY
nzD6b0EZVD19Z5MQ/6Curb/lK678KgpI1JWLA7LQWKORwECofPdcaZn+6dmy
2ELDQKIMPo3fKI4xls1/Pt3tkKshcoezC4jWsQ6tcHJrpJ9tGbFMg85/midb
e0IKtxzvl/peAHhLs4+FZ/VNeoO629gXeqpArzSQKdWWN7K0kaFXVzk2MRvj
Mez7eg7tg+z6F6Fl7tDa5XQM1YstrFYvkAvgvaNfPZUu9VEWqNecK36evQJ0
9zn3mLRAbjXL0mQHXtFtIITmb9i598aR8aZIXx6EEox/wBiwrJ3ATaNr12Gb
pARiWfDOzLLhkj5R7rxOVkuI4q3t2UlBZfm6pzeEHM3ZJPQFEa7VDDVrvGeo
HDfquBcsOFeGotigJTRRP1giDg5BKweBfq6/B+LVNSY3FqGw90nhLcYuA7LM
aNMr61pRwB3iB2o4N54+c/J0UyngA4yZYyqMKr8SCane1TeESHsXbpCaG5jH
JI8ur4RKu+7RaYrreehg9Qw1BLTUaQ78ef8sBMefwTsDGpijcqcCbxmcB6ur
win5F5wFhYdkuf4MoUkAe1HLUTmWKNU7I5CYIZ+TVAfkFLFxO/6HrvlFBcUb
+jZ/ahtnGTSy/SP6Bsf2kL2p15bku9r2Ff06EYIo7g/hzNpiUuaUifqg+2iU
CXdlxpMNK3CYH2NsditNKf+QVTpmDoFcy3vqItYJRQAyF3+m/1Vtx+Uye0P5
KJdpDlBpqyKF3RVbYtrVP3LCQXIkeDq2j3Bz2lppAjo3j2O9sAo3inw38EvM
jNwaiI0UuonKJdbRHUfBB+LvtoXGoHbfxXdA18iezN2nogiQ5ftLtnyOio4W
gUSKcO5BfJ8MHTMqNhdTEl/dtH+ohY/y1mtemKxGyzbJ0cCQnZOyllV/J74o
QU43cpHHiXYmcqT9n92IT7f0VCDxGoUAx4p4QsCxnTKPH1wHO/h2QJV/JCt3
5WlXaUzuWOY8QqHNgaZ+P1IgstcwUeiXGXxvqvgyXTcz0Sh+o4N/5YoZcDZ+
krXpQtJwLn4am9wsQb7TdJXY9Kyh8Jh6ZpnHJb553lLCWKU6xHq8uJcsDdFo
0Vo3dFihWtFYj3jS3vBxJMfIRqMxkfZCpNdOE46uLcXEcmrarY1QnVP4n6WE
0WZcKKUgmM8QDsXyIA4T61aqHKCVMq26aBbsPfNfNWNGZ4kLT17vqXR1uSc/
hn5rKo1Wl8CRXruWn9nHinW0x2226s4OckmCYDky910XJKZS0ZMlcQq7u9cP
wpSjBi89tX3YUJT18OhseQ5UCB+cwBB/q0W3Dtp9oxCRs24Tr8o0Wr9i3elP
+QvxJrUnkiSYz/sPAdE8Gssa+EMrsASZHFEPo2EyjK8IwBG65bL053KWaslB
ZvcF1XY309Mk+Ql7zXWohPCIt0oY6JOHdjtFanpQwcqQiUJxEnHfakb7gx5M
dnqVOncrznrhGosXZ/FXjlwvVIeSSbrj0tV9SLQPag+PAKJblb4blmD0LbR4
eeqZ1cTq+7fUydwjTwGNCyqYJmGp5vHORB7BRgjb9xNtED4CbPJWLNenBGB8
A2YnbAgfz3YlRtD1yNzttfPvb1eBNEpp8+RmxFLQbTnKGAL3/Wvxj42Cg2IM
MpdvF+K3ldgS0uZEZDfeRhGlfeCXvEDIy+mgCyMRB9b6YJ0rYEKXPKyyTNa6
rrFfagAz/ZwjXqKwqT0xAGy66bY4SQ4dl6HfYhS4RyfrY6fmn7RfYe6eYPx5
kfo8HWgPaU7H+rTCpad21RMuNvYkv2yJHvzNXi1Akcf1g2Hw+RkyrxEU49IC
J7UhLnZb/M0BXwK0t63hGQ4JXNEUjfHWAwgTYzXd+pAxTt14KtHTEzCYlhlR
/fS3dxZeG+pOQm+vCUfiWADQRwTeEHAlQtckrl1h2G5WSYPdsbTsXV/hkL0U
d7LK5AJxcNJ2W9RdWFuh+qtPwFnL9EXYJaAuB3F5Bb+B+Q8oUPfxI5nxgem5
Z8ahXhKZK//fH3waQr6nOLarg0S1IiUsPLQ8vnop9CwjbAjFreT4s50Taay0
G4LIoy51LOgQXWm7G0vPDnDU+iWc7naLwvbcNd+lUt3G5nVd3z5b8mthuYyC
QUrwXMt/k885Szt5vSi1FD+m//6T6I4vqQiJzSsNPL3BYQpE6LHb4GjzdP9p
FwqH9YKzQhnPiD2ovRHoPT38LmbP3LtsHwOho/NWVuRQSsjWnLBhOne9MIJZ
mEBJ6BQxoNzsf9GvVIlMAZjt1nmseOxr7yI8aSG93QzYjmjFPSPmauaMpCs/
jYP+FOxNkLG5tulL59Ff7hIgSI8K64jDHgwcWo0Mo6go8SWR6jCoijrBnOXf
svxMtPX+zzNstN57b7M2tIVX0V2nEmFcqA5e0pSJjdsg7Lt8fIO46FtovBN5
bVma4ocQY4cMObQ+wnL3heOySEcKokW7t8E7tXTyTFd7/tEHhEo4u5XgCJhR
bWtf7T7dp4oagra+8Rz54ukxaYlDQvo7jxIanyDF9Hq3gBDnu0dW33dwcIf2
XrYCwvA3vN1O7ZXHgeZRFBwefCUjiKlkm3lmv4b5y4uewlcSmb+e9hNfjns7
Y2VBv1/CEtZB0STIdKkc3kqTZsMl75A0Pw5LHkIzXG5gZRS4Gla7+NJQJoKS
WIfKa7fYHsy54G/36UZqIXSi95elR9+lkINDs1CtGxjSV8RwRR+ay8MY85v9
NqIcPUFR5YQ7Pqg5fncJSdiaQaKulC1oCq9GKx5KA9fOe00heclGz4qGQ+RT
aM+2gl754DIlaOE5cUTmvlcait+XTY+rHGku9JYLvN2HHM8rIy+dvd8NyzRr
iAW89qFj9SEfVHwqrJzGSJrHVHGZ0o6JiyxTJE431eOWPNRxF3PZHqgsG8UQ
qbrYVDaYQqz0BCH7oJkTggam6y6FJhqC0+1Kc9ot5dDm2hg9GBkONwc3xr5X
Ort0mFJUZyZ4Sx9AN/IirtNbn7vLDBakNOpJrLzuCqwdn9kvt1kYVxqhvUWn
db5AogAsLxUz827CjeebwnwWhKEsu6ZrFcmehr6Cvq4N50hiXVLPXG2SRUOg
ctdDG0gyaGgt/oJ2e7w130xEZl8q0YuwTCPu4p+pSkMvNLVPKsKnw9mZrTDN
lPXKpVJFcOKyova84G+ryHQM0nWMyPZyG/JxkQZwu2a9j6NGhVk/i7m3Dihe
vycSb+FYKMNGe5huXm6YP4y/mp5yMPd1ACOue2CXO7xKZGGEa0p3JmNUiy1E
Mi4jzzFYpFD5aZESjmB4XgPTpjPIlGqb563D3jytfLGEeD3LKVLFCNSxqn14
Ppp+T0usO2BQVkL5lQUmGBkBTWOMODfGi1p8CNRdTGyAbtJiHuWAc3Jgqe+R
smRs27/pqwl7i26ayJgMghZWMhzSShzWor9HBtZ1/EbQdbviBhWM/xvJvtEm
VcWHfSozBHjpW6B5bQZdZmj+wIHfZupHBWYMZ1kVCvMHYvud30CylIhTkCfc
q+Aba+KvqXFGF7wcKx8jE8lEoHpNV/60PRFUbjyGUZkepcyo7KWt6tsjzqpX
vvzEdKFMbmCwtuB0qJi7LYAT3jamyePSPo870p4i2qI+xEIyJt4x5VDL2JGV
zWCYw3KiZPXTJzR1iTfb7VOOLQ98fEFl3ZH4hVDNYb4w9FBFjLzomaZWRzbr
IBfq7+hH4AkRZi+G3MddwzyUAE3NjAVzrYLnXYPqa9QHwWnclm6IyujYqmXb
+0itgWu9DvV5Rg+4Bp0aPCDml6Yv3uDfe8Kg+AHYbKyMP7Vy6wodwXkBV8io
W1R4diP5/9jL6NYgGP1jK8c1Fupa0xqAeoD+lkfk9qDjoEOskGsdY/alOa7y
N36mf9Wm0QqAzWwBItUW+knQwH/HbmcqJo9/gjFnGt+zhEFLXRgLS4ja8pe7
kG+zHQch9+fAAsVuNMh9xXZ1YGM59nw8qAYaWmwGB89q0KLqyjGNet96D1/x
5Kxk+0C7vY4PM8Pv4WWJuCWKDb2IAIeOAKIwY6eLFMysdVSAkXZb48t9gq8+
P3/qFTZx/FSbbJGW5U/GnKLPs8ifm+Lb8SjZv1Hipp8qHiWDzEsUu+043yO2
ppAok7wGijDdRkNinEgb5HDSssgixMUQ7LRboBDHUR8pU5IVCljjQJS5jxc2
2AefGhG2KGxuNFjrW1H9c3EvR7TH1MN2tLUcZoZUF5hRfwqx2CDP3uFnHEGK
vCvE6JBnmo5LpXdjr7Nr9bcKUFxa94lp0kdqf7EesgeXD/hfBEPHkrpxvo3Q
OtiYbj3/EXOQ4+LwDDk6Elr78Jtjrm2041l3cbKMHqEi6shDwOrR+nge9g7L
T50ACq7WANTjdLbbAulUEKWyRd6WWyuQviKfpvkJbw8pPI+QWook1fR7dHil
TC8pEUUTbi79omW7dnaRuI4uJYkxI5Fudwhndd+3K8u/W1sLq5XfT78uj5VZ
xv3ZhtTHPN6OqnZ0F6jS9Z5MtOttjwHeqf7JTj6ufKrniM678F12zV++YGwX
Kj0A/Fo2nd/7b5oi7Kh7Xe28tslZhzW8NOrtgiunytuPgPynbRpAOMOXiz2l
DqqCd6SlNVKbFGHBtzFSRs+tnCB8fFHbh1MUDOA5MqCmtMm7BTcmjnLO0KBn
vGf57tt3pbBFw34qI4Vv6UjDXl68QdM9zS/REPplq8MJ//ObRwjZm5ZYUz8X
Ujo65aKF5epJVsfStFQ/YYusbDkW9+uXuWIf03xYlIhsokms7Agb0YBzZIru
RLdfsaI9w4YxC5jCRcokU75v7AxHhkRafnfwCzcRZVhnjEqD+ECTPXadSKa8
kpqKxsUO6G1TfM52FtcdQtzkwDoFCQIgn9J+zFKx1Wpe9Kk7zYWLEHLaNPC6
SRDuVhpzekOLXTJwxajV40KI8/T0l0dxSPfzwZpK7R5lUcWn9BHUSMK6/CeF
BWxx+fSgjB9ubokcFl9BSJROHRnD9jc+lxTGvCN0qO+z2peA/JJ3Wehh7Eka
sXz3XdAdawr9D5eFPjGwfsNGucB77vjbo3jw20Wt0ZvYy43bpgQl45VF92cq
IYV/aB8Dy0z0HQ5Ak82bv8riSX3y0fGMJJR5eHLElKCOyxXtM4+3naPsz0Fl
ja1YQnzfDfpFHhvDD7kNDJQrj2nPzw2tnTs5yvbz1tIEuBoH11/qRFXKGCrP
k8uaB83B7WGAUpW02J8Ik9BAZiq3T7FQC+RjA0RXxwyqduMrz9yVUqdVx2WA
T0CQSGs/yIOPkklL/5k792Kyy6CcS8ArolHorEzwM6nh6FXBjsCL3fw1IsLO
iIc1FfyEJHDLu4MVPHDgTTVq4iTE3Q4p5VuE2cnctKIOEPRlm4tKov0d0PYB
PEhlNBKlp1SMjK5+phHhcngffZGaFBOdxlYaMyPHcgeqAnXo9sAl2SlQb0NE
hEMPttqSIos14r5qyNJ/MHrVSGhb0xW7dpFHBQXeZoYOWaxQOuERD+GyU3L+
6ajJYSySYz6jC22xDgpRx8M/e33qZjJkvpTk8dm9LILZya6xSKnOHB7gTHI9
ZtiBeG/0iQPSWi+Gvvz/pRQYGi7veZYgoP+MH362WysJSj5HS6Ed4GZGAvzo
5VJCk+XWvh3oCFq+lRZu4IJptH+JUXXPhcIj7T51jxVDVkqe3+l1IscPKXHx
KvjOGv4wyog/pJB3hzIc/9Flso3kl58LJDdn5GUaK2SXhRM6/hI3PCiKVN7N
aGxvvLRtyqeA36TN4K8gHA3BkfmkJimC1mPXgAsC/fVJu8wgoF1vGbgeFQRD
49BGhb4DcUG0sXblkfw4TeCtMjj5Dd+Qk5QFBNpibP3O+zUI0qPmDSYxRX2Y
nTGTVFD3fewQxsoKTu2yWmhc0+4txrXDTywNOtXdlm6Dtx9djuBqTRYjp9ak
KeK6R5JGX0HKqfAZQGhBDXAHNm1lBQpE9tq9p/C7iXsNeJi9IQ9q37080O6T
IhHzeHyWLO77JJ4ytluY2iRcEaRYoN9TeblWro/jMnXNsBirXqVdhFs6XUxa
XVjXwU4d1QMddNgjZ1e0hQK2NtAUsuIvB4QdGqyKIvFqhE66l+P9Ik6JoirJ
3o7Gg5Pl6JMN8bevMyfBkFp/wkfgvoB6ckGcbXKZSW190UVR3wImw6ca2RHM
hQnSOwieDLoGbdO/sBSoua4SwIsPmo/+df6Bfs8X/6OxhTZeFz2EXAh/Nvws
NFjAn8eYlFvOkp8b+cd6SdoZfEaarcb+HXei06vGZECR/BbIxJe5y3YjjOnJ
9YVxOfLiYdMx/SPFbkYld4c/yU1hvNXPQpC5x/9YkzJ6IVW+QZfbNg4Ey3QD
y/+iThtbQ33/1nO8dDPugd2Mxktze1SX6S4hk2++lCYP+LQ85+nyT6sJ/nCI
rzmidssAYlBd7v8TGYCAgKY22FHnU4OCnq9z4EvtrfIiAMFM+ecr6ITNnBA7
F1zeh6V2FWK9nhZxIm0cvEAAh+3KJ4YrXqdd/mcZic2clO5NEQPn5CF+sW00
MZcJYhaIw0BlIk+Gp2Y5TzTZ/jYz7gM9d+O8TBvtrIjXpy1qAwDIjorMngSf
7LrdUNN2YuZsGa89aEEN4qh+8VPwgHTky5/NhqkKiux0JydmH5tHVstYXsZS
ddD8FazoeIILoDtUhTM28Zjhc0Rm9Z8NLPxS+NtiMetZ6yJoKAf98uBB4xem
t6mxCXeUcyXxvqjRTk/83/kzT6zITOOkUPbcRZL9L4vokgdgQCOv2Vsno9XG
Ol1uoCT5JKoZdDN5eJn+eyUtzSfa14vPi4b2ryoTSS4dE+7n9ChTGllo3mFB
LwX904nYR/d//R09G/mT2jnrXBz5C7R/YgzbLMsKfqAsQOM8qwaHzzS2ThwM
9EA8cUhbzvgcoOYYLE5F3YmDVF9xJ/E6S9m8Eco94uJPaQLF09TBDc/FO1xL
l4HFMX2JuVmh/auQ/rKaZK6PNoJKEFSDq0UAdARUwTiUKdkETDmzAd3iSVVJ
ETXTsnAQ/USjo1urxyCRVlUe+El4aAjZXcLDDy5EbAUzzPjcJTS8yJ8C9AxU
QceFrPrHW9Rov3BG4C50DjlujDLc7q8nwnF8ycnUVVyjq2DHTnycYOVflV8a
uLQF8cLwooN6fhB0bPdGkWeZxNC/REnbrZh+A72HnI9erkuDmsuUY7e3Qceh
vsQ4UB1aBHimEx3sTFreFH/6k4D5q0yLlgYP7+0WiSTIAbpHnzMOQAhhSXbB
PkqwrumWmAwrFm/jENVrqtdOG0X9iURB/jRJqbHtWe+7q1NJ72H7Tp9TczyK
iXMIhHUkMI6aD3IkGC3VC0yXnKKOnoAWxQSynp27njwUubXwpvYRHUPa1pRV
T0en4lVgPU+wLKZHBtEq0IG+8Z2fcOWOSX4X1nzpX7rKP3roJ5rHZNHzUOsW
1TkGJY5WmQNG5uA9Z7/PMefgfbMyydgHhRuGWMI5eb+PU8dk4CvrlBz5x9Z8
7WHOA+LySTMJ5n5LKoHOrpCIO+i5LMgQC4lqtFRU9xsAPNd93Z7fq3DkWwv3
zncR1r/Ne68MI/v62HgHD0vHw4z/mjhZlpxkM7JUH/fJxJ8ZB7NF4XgAlEgY
uAVTquxzJ43VQMVDGvROITdOiVYArw87aKhqTm79s2/T58WauIOFaqVyktZX
zaB5DBgOeQ8x1vgCVwx3HvgDpHwIyQ2dhtljoN1DMHCqYlaYf0Pyc3gC6g6c
OjYRnDfxRTPSBxPl8Nz5C9IxrArS5Kzu25uZLFJVDonP8GTNKTXqcb5qj0gU
gm1jUvsr91XAqTvSP7k3QEwXsLdj0q2iXoO5GjcXiqK3P2zz3VvNLmSkKRHH
oae6IHBgV8neTc8zsj0H7XzX/2NX5hTG5zy09iahca/CKqlYle+S124KF2Jy
xJXOrBx0hFdX/Sr1YUdfZdyP5zR5vzk9LDOb+HtpwypUNa/+xmJmrfIfxf7M
dzcMqk32BDDV3wRV8edujx2daBYhkLN0rsdP1+r6ynLEOyncF38e76PZR7GJ
GqoAYvpyBwvxHTowLr+a3D6ZCt6QY2hzRpaJPpe1twDr5X1IomDY1yDcpFSo
C7ooC+IzfdShHKnI+D2/85RsrE+f2cJbm1VrUcKIXH+pxjBNkszp1P46bHr8
OS7lTOE71kwQv1BEisJGLpZAKfMMX+nIhNhOM4eXs+s6xgDcB6riydOPFMDa
I1jatAGJvUFPPghJC9uWKL4Wx5rPqOEzIQVJGlxrUFiVbWx8OnlscmiP8Cre
2W7Czm8VrLpgiHLjf5m5WzykMTtL2Wqz5m6J/rkEnR5zwLLsyS8FyzaoGnhI
OAxPHdhZaYlIL+H6GUNHpeggffwAeNCDgi41urUrq5wJcELjGG3Y/KZhrGJP
YJh/4eWZMHTN18+wMIdwqZhfAp90xCExOLdY6K6jHeYYNOTNpXxNQHrnznOA
BAYouOpWaI2m6Gf1DT6y/PKaipkUDSFY+xeu2K5L3SmUWwaRcXQaPsP53WpV
H8/uEK0+2ZGvyQWXwuZRPnCKqVKL3ame5vhSGgjmFe8Ad6ap+yBB4Lk9jVWq
jP6bgI7E90imMiXS0Xu+u6AOPjYkir2rO/NLK0aggmH97PAveBH5EWZB/Xvx
KY3WPR5aYQk7wjEuWh2r/SFf1j2j0KusHUCzSlDARqAyDIc7PeA0qwjx6Fvy
6/TIauNLO8wqjZKbqRnvUnq237R8CUBfSLRdwJVWPmNgTN9txAvqOICL33yk
xlTNy0q6zje7KYLsE2uqrzzgZK2B2UIKaYIxDs/SmpRI9vuBv4Qg4uGubjXd
07MrqpE6UX1oDZW8ZAGXAKcTQfzwMKipApG4UlnAPc5RXrunKuBbwCZ+6LVx
GRopjkXHYo3JL/MXHK7zI/3edqhLW4Kf24NkXy1r+HQY5KBZBIqOTtCxdgnP
5F8b0XYDMxM4l55KNzbyErHpvszaMizJrCSJa9QrJ59BRkYA8b6kzM1aCKn1
UaSUpwxXf/JZwMx1Q9SdkzV1+HdqDFtyJeJBjJjoQwTQflmt0r4gQxivV7DN
kE1qP95CyClUl2gmYisionIWfftxHVT4z5NAjw6zzc1dEv92tgebvvDmRnE4
AC+a2xkQqt02yiMwyAA54Igb5jSYllGasT6QWtMIi5Djx3ka4F2vstDenUgK
fxgh+6mSY8ck9LeD5Y4+GQ7/n6fRHRaKcb1D53Vi8O+k+eR04EnOqzyEGwQU
Buj1jKcUAJuB3Eo08BLBgSmTqqGdbfigugskzJ5g1T3EbXpTPGRbz+TBHHcg
22hQhjrV8KG8yTXLLwZ5fk4EaLAmQlqe5gtsF/i0biNc+BLRC1AO4OcCTDB0
scHU8cVmMnhGkqwwDldw/rK/4Ckw+5hNWWBbmq9xOUc0FbLQoFcpTuGumY/q
qPJIgjh30lUPAsP500QYbbFDKyrCk+zAlRIPciAM9j2c8dwEgZg4nT2uRCXB
S8ITCsmDKqz9BNFZ4qHf2bvKEkxEkw9qX+269ELcvlhO8H7nuLeoGMJLaL81
L17KJLw2e7lSgpPVJ+ZzoaBObATRK9Gus6O68geZSzmRr9nV1vOQ5HEtoY8S
NMQtIuOc1dtCeOwB8E3UuffzsQzQK5fBTx3J2dpDgqIPV67IYVTP885EzNLu
9glcPwO8aXcD+xzYTrYOMIaEQKaEsqH1XaXi+fqS/gKpdz8kKUrYWur2E7H6
FE2+if6cuWaJHv23jpLIgKwCyTM14hyq84qqBnJKow/C2vDFFn46XL65JI6T
G8PGQAgqSziQVHJJ8Hx2IDZMmmWZNYzRnWKcsRbSImUPPs+0BCvp67lKK1iQ
VqxTayvk4nfl+rP9u0PibBUPWTq71xusNUtasGdnCTp3eNvIrhRczjJnm3dY
Ki8qMRF35re1WQAn4fpXPJzk/NbRP4vbEC8EcNwSHTBcZYkdyGkDqINlllch
ojoxlU2GrUVUZVxnlv5wMkxT+Zm9BXYiFOOpI0AhUKw6clYbwWpTUESC7ubX
Gu2yThYtTNvxm4+m+mE57XSC91ijO/k7iOZD0mY9s0NVjDvPOBSHJdPB9Me+
skqGf/LTXGMEaHZGWp0p+B/quUDWzajDsmlEIQF2FG4CFIL5tFpEIpn+k2l3
ZClxpADMjln8hCFkj1d27ANoJLIV6zfSowmRl1oGM16IHQ6cg2dlEKEa70oC
jbvDgZLfzo4sk9hx7SnS2hAIysHnFyokX55Xay21QC/1J6YtbG4yujB+ZXR7
3nFJpIKiJys/c6OG7ZV0S6cf9FOf7cJavM+K5orRrK1Q1V7uJNtewrVMz7Hu
xUQXiL5FoKztTFfCmu6g1oCGUFVM6JNF0QDqpHM+ICtQZcysIkyTx6qmriL5
8qBoV05dtT3MtelWsSTwr7G5wnDSfRqE3c7THtRHXqViMoFzx3kSzUy0/3xb
zP7lsZIt1aBP5ziWqkdjfY6Mu7Kav6UmRq+X0mO32hq130a0CvvHS/I1wAw2
uuk3syyjkoRDlDtsL3CBGI2fqIJCJZ0xYw+QvWppDRN8XEC7UUccVOBrncgw
PBVa8en4JSDnvEy+qS/egYRHmiHVuyETXt2A5J+WIBhkl4xHagFe0bXrTA/A
H6ejwK45I6LpbtaYQmHBKpgnnxqHBF/WFUhZ1cV1LSrkwBb93yiSCA77TBaN
UaGKwl9W8D8ffZto/v6qAx9Tb+OFgSQ0wvRigZh2+RzYItD13F2dXnT/7bR3
oBzrNNJO/t4DwnpbpxmI0RGEMpF+w7YG+/o1M11fc5WovcDGszBXNv2eAnrY
mIkDjFaXzmIWV7hStNvKbj4/vpxU2f55wmMPMvKeCwQlHRePOHbKQKzM7MDd
Pcoun+NqlBpngrzQ1MCNLEJcZ1clEtCNfXd68WBNbi5xXNiZkSjevSHlK4ee
+Jm9dCAg8uUX4EkS+06amE8mqch6PDWb+mUbuktrDN4/kMaNnIzb871pf6Df
ADy/qv60vQirRXagyj3lzLMtvyFIy7yjaqBLR8NSpiUd0Ze+Y+Axgm9XvBjh
EoFrtDACtP2sWjanTM5CDVaOBu0xAQZNX5/EJkqINTWb2w9FhcMSQlJEVYAx
zqHrd5MiaYnMHK2AEVPVLTloAI1QkhAy2VTzmdhCVw1DW/QMPlIk/wBlvx2H
33Akp57nVV2WkJSsGp0fta8Ya79TarAAVoLMlRnHMthl/KSmsf9o7zHMF2Z1
3eWPGUk5ogDZq9pjt/iFZu7bwjv7nNxVvvWpOFF8hbWikY7SI127A0ybjlu2
kvQgI8sP0B2VHP/m49Oh9psh7d5h+RByTZW+OEJ5zYIg4DiYcd54LGUo8hBS
ZSi1gOvmy2a7aFz2eLF9niZ3QPu6Od2KLaUfJh/MO7+k6JxL/Wcn9+ggI1Bg
0FZq7OSm9L8auLPLCVxQ6maCTtgr8obDjaivbaArXq3Vh/Mq6MODoc3TL32X
OJ79ps0BBFGdUm2acE+s1LoZvRBsJOf/W9tezBgJuhSP80fXA0YrefCVzkxE
yjrGjHEXlsBgBGdk4iCPxLfBD9M0LhKTIPdGB9trXKxRnXe/0+DlxVZNTRhq
D6kiIguABzWJFRrVjpe0gZtxp6rauhJiBDV6TuCn5o0rkVyvYTLwnKtGtk7L
fnXjNB9eO4hYPI7Kl9emb/n7Ib2FKNoMurh+CP0fSF2J1TeqYjFdOSBgOWma
UKvAp/sJ+vtKojaKraTVJke9OhQKShYaEXC0Y8VV3dKJwUPIKlrM9Mq/vdP5
aHcIb1RLEr2Bqiyar5cMqT4sIK8j575zTLQBaLffe4FJkvMiy8r2Mph81OBg
cl2wNcNE2SKf1BmD3S0ffaup2WfxoFFcwY3LO8uDWh8ceBinX1wabAM4bLsI
g+Zyn2DZbofFs4cJS791qMo9THHE4IYFtgkgPuOA+RHi30ZUMp0kj1AHcYd+
brTR1pqSh6m+wt4TBIXX02Rounr18mQD6Zkv0/+Q6/a7pYxpK2UEQmE2NgA6
Ar/GCau5uae5UYqjqDE6AsrzSgbNb26TKtZx7Mg93qcxSuYyTvYL1IVw3iUw
oPvGkGocvXyk+/xA2VnDqTRpYLyg9FF4FjipRRFnU011kFDp0EYgpzhvmXSo
CMxJON6rJGm3dNFImDEGx6HEIOWFmC1li/LwCUwnKKL0E2HUDXxE5VF8iKLb
COqXdG8Pd2WWaL4bK37kuHZaYdGS40xQHUnuF4Pc1hW9+TQm+pNLz0DO2glR
UC7BpeAvSBf69BXHfKn23sY7Sfjn7xI332lzZjLlgm6RXPg/wmuMeq043Rtk
iSjY7NpSA0zsz498Ej4fa2Roc372tqYL9gitIfHXXRSQzCgb50EQh9bocyYm
qIlfLjPHJjgV+bb2ulDopY5LDWwGBRvK7grxjJ3rE1LjOTj4rWw5Vdc8efDB
yDmv4cPc0qq21kTY8tjCMA/03TZJ1pQ2+/OSZ1rnLnSj/Hy57ReY+sYXtJgQ
8JAwJGSWGdr9zng/MtQARDTH+4DilRdI+NC4PgVxlyI7YFNVpa2FJ9uvgXpo
mKfzVGQu9sxVp1np0QSg9ki7RftE2k/0XxOIyXTN+jw5511KLQhT9w4sTYHz
feCfohJRCOOp/jpe6jvF1sYnipbdIeMEHPpsdHpx8BwimRM6psas3G0n5vCZ
p9dHOnm3FW9TMkEUS2kTgcI0mLs+nMfH5gFcgPKsufGm0z8D6qwgpJzaffgj
S15HZggX/DMroW2trsmrgw1PZkJkkGS0lk0h/4heU8nvvB0tMoGKDLTwbVZa
yJE9xO3n4rQL7HTra+0udLJoY08OxVQGRLvSClqSRnGHkw+WIaSYbZ2J1GwI
8dw5f6Z1pnMdyOKDCLcTwa0ad9IBczAkKMd0ZEDeJjTYNpNrDagGUGIy3wpa
qXizIf/PxzDijSF1tYx9DJP+J1Nfxtq4XhmHThPsTOYAfUBMPDICiPV3OdHu
KPeJnFIwM9NkJmMOaWIWyb69LsRVtDk8M/MCd9XzgPjKaiFMGlb0IeTnz+iN
oZMYeE2Wqx56X2TvdUjqhSuVoVcL8FFWASbRlRHunCzL5I3Bk9jaqE9xus5+
Bis1H2h8IbuZfQJRYuxFXB7nAHfAzpUL1bVwvJXsMDtD49cmakocg9hZLXTl
UMX5sCausPBBDyhX6JPr2RCy20zv35EFk7pOTyL7xDsVGnXOXMMO+l4qQfjJ
qxz/X4tRG+nlcPo6UdoqtpN1/d18iDryWCb68OQfa50z6TFwY+FRb7fOYqhL
bMXwJNisg7LbbUlsRq94JDToAHrjTKoPZjNsedaZilgaRwehmytXtpTtstI3
ozowOkrJkKsMAWKCxQew1EVqm+lZHN01M2DRNPGlMYVEFbEEKa2fDhhFw/h2
btlRWjnixkDE7rssIEV9WEkmYIHXGUcAt9bxILjiT00vcJdbftNQTcA5Cnet
VpTu2Ag7lSNXsqdW1lqMS4JXyNBmhSOjjL1JvSpvf0jo/1qXnL7Dag5BO6EA
EYGVNSg5ttb0x4lE4UQPfJVhTqJ+ASR1na8ALCr2oRTQ3I4S+TK0m7Gi5Cvb
glroAfzrFp1GEAksOz0YCK+H6HNBtisLQcDPgNwx6VXQrUBMAGb4quMIWjKz
ZSpEzeUrEi9eMlDTNBOwZWAJrEd+zqAalSOngPqPtj813Ijtcf8Z8w46KcLW
b8zkjBDtp76zdOTohnsWy+Smj9Ez7ciNsAGzTHx4AyXf1jU97Sz1B+DNEo1T
Zn5x09w9nsBQLFHY1InZ633oC8IKk9dMHCRwm1j8ksV1096DSqrcSRyIoRSI
l2yeMR1GrHgNYBNCw6Cs2daz0JZhD3+X/PoUDBDXMqkdOthHtQNvatn+Fj2D
AxEXSKw6VEetgLeTPed7CI+YxVoU0Z+WS9oGpS8CEsJl96oDIrcWJibcqQSL
QbVXYY1D+Q3jpUXddyCs7XuZlb3dKTzuo6FdeOiu34ch9up5RQ1m4FbNykWn
zAmPvThRa0rfM2nNGqOSiVQ6IZX0K4pYIarFH/Qzilx+WK87tNuRfbxMOijD
IxjfhmX1cOBR3jhP9U7mUSu/zB13KlzsfvvncqFTVT9vMJNHQ3vWBlhDEuwe
o7mRyah/epa2vsf1rSB+rknT2Fdm/uislXf2Gp6JMiHBAd8CVxFhMLbJ+UR+
WDIXcj8PQwTVceP1tK5L3koSVfnePwigF86H7p44MV+CKsc5123CfJph4RBC
TXtoteAls8Y1lseq+8WlXKEhKsTOK7LaF8S8nWXTXpH/MitUmbZuUpkpsQMQ
kUXLapIUdzxxy0mSG0n/lc0l6kNosoc5XZsNG63cI8hviGx9dIidGhoFczT5
mkhSgo3u46DQ8aPouZHqgX5jJ6OnmoJ6yra7eZST1PcfhMFgsOUQ/nLxmD2M
KdJ2l9cpqHFhT/VM3bfwQXIyyYIkRJG6+KjUZxEDo3WPAUitHYx2ry8KnaHI
yj4JgLtIMHZq+Uu/76onM0MystF9xou0vLROx2Td0nIGI+kxUf0PBawFqjTV
nPfM6dHJRR98lURZM+s40BsY3ik4zhOv0kN+DIRBwvF6qe7RjnNDvuq/GCh5
uuCFwr3a4X9QpmBDUDTAF2uZ4LYzc84ighyRD7mBa7NFK0bYlXbOeKde3VE7
46OWCzI5+TGuoARc+YrHft0iAQPRkbSpKi5XM3VwbZBP4cYmP9wPQqkn20kN
vlVhEtvnTUA9zDm71oiH9L5jdxtVSoOOTqimJSyGVHLndVkjsY8mp0IVPbl5
WExf6X6oF8JUCOjYTGhTz5inN3C3NcsGu/3G+Nq7Bfv4j55iaUIBu2aoSrER
KGjXEVCnWuIEYXxPlDuAIa0bJpsh7ZM8KKtd9o3dbbDuHTWsWAGHOFuAcO5K
D1Q81MFqwBOrrfYOxXeiA4M/SXRwCekgNBaayOkarJTKeZ6vvFyemA9+alQ+
X4j8KgHMqjVJrBkQZeGIMLz+CfOUEPjecVeZ4CIbBln9y8zMHhCraT1HEGkg
JqWq7ppnDOrpdA/S5GyVXhEsTQnuZ4zSeXqwUS0qTV/+lxbY4PTVGE7teG6J
dQ3luP+opohSFEirNtwFCn6vel0s4iELTzQCjbX8BJC3KKX8xUntBTxCHl5U
alj5MPapNOtnE1j6iA/R827BPIpZjaIB60dmKC+IckA3gfvRP16GVYIuH3qE
hM3MGpf+K8Rv1aFZMX6Urg4LPu6YqO+YAEeLac1HLZPIIrznyOeH0B3cc1+E
qHs+AnN8b63DCbBShCNpUac0cGZKgIdJYQKFAdPThHv6T8fYOiTay0tma5DK
HXf5Kov0VqDj97n9DeDXKpgajcSAMhO6w9UxhCoxMGNpamwdiazbfHkB0pNS
oQw+VDXqU7pw6KpY2QRgq93xM3Dz7TXZ+++qKZYywo7WlkNwBG4oN+lOoiVn
yNJs6J8PCLbB/LO6aPghlzNfMN1m0ygxjvdI1MTy6YVFlX02XwvAs12uvh7C
lf6Ni3rhmfmM2fz8ACXAfny6vmGQmw5DgIauinAYumGiKkyKWnaWGN+gW+ZY
5wxboDB1i33yyfHBOM+PWFlvcCaB67EPnVfWGoesb75JN4h7uCSG/khfSOxf
bOQlZ9Fls+Zy3XCMNy3P2nbui0lLFdlyDmbr1khYq94HYazapPRmGRBLisct
FqYbHKvPPk6uJfZCaVen3zskzbUzvmzGkCurYJ08xNs8OxSa1fa/ONvyCOII
UlbZqdrlvRDNVdw7yhAg3ydXvNvYteAmOc6KdEkskVQvPoOKz4bQcVVjFOFK
pquFAB7NlysXWYxFC0e+aX5f9zyY6QXLysRX94ClOh4AonazbPgV1eTGyAua
E7NUBNdTrAUM7E5N+Jng871eMjLBn+yKSKeVrRdF0NhSlPIO/ZvF46tyJO4Q
Gm2slVIgWOZiEztSY8l//U5pLfs+oN4EK09s/3ElfiGbrtXdukVmLRQow629
J7OXG5AP287eC706jN0v5wsxQVPnia7qyEkQ7jrAKZkl4liZaU/DD+RPywQz
0sb4T840ZGydix285mABbEqn8ZnKhXLKhb4ESbu6EFeI1tG21pZswkaWlWaM
aboWTEO2dTexn2SS3AOvZXrUc/D30R5jtowlkBlz/3oI5cz40z8dxzXphPx8
WPDCfswQR1+qyODm4IPORKJK36c/HpSrlNZw01to/rpR1oPR+f1ngkAQyICC
MPtAslZTibFhL1QEkLA2SA7gfgijwfE3osivFe5xL23PhKtSMqgDdrBUekse
vwWZ3Ch9nc8m9a55P051QiUQWp2ANDka0Ch8VtOkJe5kJX/snjim5Nizsa2Q
oNOpkHgK08y30SdkEssyL7XvNX14wHassP0q4NLmVZJ+6IcEm29ipKXQxc9P
ChNFEivAGJry4T7QTaUmYo8OqfIc8vvZQRUq1hb7SXm6DIZjaekf1GzbHsdT
oGSFUrGx1aFkXpbpIwj6Gl6jqoDioftN0pgjiLBBqhMd+jz3Cu8QMU1uFGGz
52vprcOTdnjinFSM6KElk1J82gykWdVeYVtTp+oy/Xwq8HJSPeSQgQumW61U
GFO40SUlcd0iJDZqzp9/7cXLYi1cHYKSDVervW4v36V+4XCGoZyZkxFa46UN
5hhZiY3lnJGI3eSEpNXRalJi9OgZoNuGwy1NmpF9pXzK0Vm1i/3UzxGcE632
mVsKbwTNFMFfIwlL2VF17MdXOKCeZgfu7GM3CgRCwP/vozdX8UMdSO6ZDaa2
O989/ZJuKls6gv4lSIYaWRzuTFra2lHjLEiL9TZPjeYF/+h/BCsin+bnRuE8
17LOIBEhOumpiWdQvj2tXTcLIJ0gPfxraTp3OfpHlg22WFe1iMOdnCqM7EkQ
nDGx6Dc0kp9ZGw0fz7IaEtgaPf23KLvgMsEPjU+2mnYAJ8hfCsiNUigczcRb
U+0QKtXrMHkWn/xls2/c9R1DcW9SR4Six98e2K8tUNp1t6gTyJYoWKpoIr1K
HE7OctWKVOENw7zCfdFW6RyZXH6U6uLprBl9WY66JYlB24rc3hNs7O/6mm7Z
46B36IUMRIVsYYY0fnHbYwEkPWPmRfHupK8LKDriUzWQAlNVusfQ62EBm1h3
MQevCeti21awAb4TmBEqxeDtni2+JxSJHG7m1R915qfaASLtbJFJCRafbpa8
72Xwc3lyhXxTnF1Q1mgEc3J6ryp0HrTMoajOOG3RtDiBb1UC6fGtnUh18qUF
e+CNzxPksADm0OsiZ9AaGFjhjNcZRJQe5p/BEyNYasAw7sq6OdYDazNQKvf4
5/6bj+aD3x1O/314WvYW3RtDLNyjFchepVuffObqV5bPJpmkrN66u8ZMu169
5LiGQN/9IstnLNCFrIEPxkrvO5ze6z45jitLxEsmegHSiGxaBPfedI/7Qo/t
HOPWXZW9FWyIvrS1VeOAeFazvXvW4wMJAwzl3RFgz0TqKwXo3GOSH/4fQZI0
cjrkG14mCWYXxcn5XuXE7nQuUYMXsQmC98UXXe6nHCsAhUrKPvsqdZ5GGVJ3
5oBoPAcSQTLnZWk0C/2JmDUJ63XGj9XwfO2Y9hga3njviakbIYtikZ0Qm4L9
YnKiUjIPlSZcxoJd6NWMd8HSnQS1QkzIwwCu1jCeo79RX8P7/DFBgrgXo7Yv
T445BZjC550aoTht+FnLub13TlXL+HChkIIkCuKcfsRJaGErHRL34RXNlnP1
Wbi1hK4zcc/AlduDUTBT9RpQhrLyaJjrNdpOsF1GqXvGjOMLivw0MOkBiGNN
124IEDQHSseczcGhCderuZQSH7kk8as+QZrew4SQarIkrjeSt5vsng35m2Xe
AKawfUpIa+PmVN1eEtx56c5gvD4Z/gv25WnEUITkPoto5phXnThPF0GRaJEg
AswPOhNNYwsOJv4S1WWmXxWjcp9zDbeocawp+5WLbiR0sC+0NU5qOd6kHdx4
940+eiOjr202GfheTaz1vdNBK2cueju1ZGFVVAY6jdFMQE1x/TjS3qjk9gnp
CLb0o86x1i/YzpbPYoyC25ejxcykoKRdpMHRgeJxr9A3dmog4KGO7Y8K/u0j
No/uYU0TqRLlyDaRgMXatkqAj008MOs1s3megM0dODPSY69qCKaZp4ZUYVe8
aclQaG2R6/4R7gHkfWo3VinDYe8Vg9FxKE9ao5cY/Ip4MUY9cinNz6nvQJsc
k0la+VTomYPJtLddsZCkBy+y88N3uSukBKNZf/7KqE+zzXlDmIw44tYmRtmP
PB2y6bPJk4+CrDNE9aJzH++eMy8IVmJ+OEXCzgb8q1KR4qImvGn8pOb5dgz/
LaML1BesQ4yWj6Bj/AJBD8cIdz9xsF9e/Sw1djDlpppFqoQRNJAiXP3iyyTw
fGNzS//q4CeAkpyAknN28uHImzKx0LQeKgjchMoaOz+/d5/zMB7a0eDpufHx
Nj9895/snmWwVMoBqzRKhF7SYdO9Kw0241bixTCFcJXXyRABqbA1HdD9Ly2X
h7QfutD6XLxhIxaYoXjzVjhOR1BJhlhoQH8+M4wG+dcwhGfGwFkR8a3kGVMx
oSZh1cxD0VHU50vyU3JbdfUichKReoD3BKE8/21klzyGLfXIrC+C98btBFxg
KaGplhiCgLuR8VY4OUWILOF1F5NZhfbAi+L16oh9rFo9p6oJSWVwRNyODT59
o0+4F2QJrTIai4Ai+2/SqyvlZeiYZUbhb5XrbXkTKKc6VlsU1fqeYJy8+wbI
P0N0Kzs90duUCDxAMQVvYp1Iga0Pzt2y3xRbw/CixxpN6/zHufmjE2T4wATm
lWnfT+ZMToSHja96N67jqgjmyNpdSIz4av9jndwmxfFlY4Z2AqgG6rpJw2A6
LTK7cCHmoXzpuo930fLDguZG3dB7gr0BjqVHnuzVgvBqliQYiQJUYHJ5xuwu
gMI2p1NwUrU9/EDM9rkAs9EnXDlGR2PvkLM+XtfsnxMtz8MsvHHaRLL7pR5u
LO+ZpMVjIRY2+urVckZpDORqEPCNNIO3JEiFzt0Bm+pLRvLprH+FovBAktvZ
gIDMJ1e51D0MjLOV4K99hgM0Bf/nyMS41ojDG5F/2IOPoDqTDgsBk4imYQGM
7J5jd+0hJeXMT2M/VZLjDrR/Wx3vzZLHga0nOSD9E1OXt/1Wmhff8ynKr0/l
4EWoJxzOhBFIf1T6pvJ8kgwjJnW7bn9Aq+FwRfg4lFny+FRa4J7rSxyzH2BT
dgoR4eF8RlWqYSvm8OM28TJyreU77qgqcqbwyoH38N0QUXW1v5rTBRv8ziH7
fxCHkX/X76uR3eaj9MiqL1qldzq6r31bMYt/aNmFzwlRPRXyw5EqU46vA9A9
q5BI+FB8xZDYnM8ZU4GwdE8CR48DrZnmYg/ne1wakcSgchgQOrceH5oYd+HI
Y29JbSDlvxuMow5szF0TmWddvlsWNp8pcSaw1QXq3dAGXDmJGM+XJfgK50L1
X0V/0hE2ldydAwaxe9pJSeb7RVIYvQ0VvFKnfyq4t7cnUtMGO+hVWBJFCOEy
cXhDVSRY5g8yRpAs053DSmE4wbEF5Wa2kZRkqTUXqy9+Mou+4LX91ppaDh8I
nC7WlsMaXwC36qXnKsMerETX3Y4AzVZIntIPaA6u25AR832k8p6B1AwVSEwx
1gMONrXuFvYNplc1l/YqpoWeCk6Ccu5+SdkWXQWYC4RGh46wz0jcqzUlFgms
xu2IZCccP9Y6+v0fONEgjgGophGKgdB2beICNchB63krRn6rWxG7qxBAvAji
Ztzf1/4UYisut9GX4UhIjODTnn9f5eFUXRBFz6YbeBaOeYbGumZKzZbwmYHE
ZDagRZQWEZq8Fb8wPYaIHb31+EqhYoFMvMjo8qPOVXSGzNJZmbq3cHzjqOJm
fT5NUNlpWMtBuyU7EsORoDx1rMXa+2LtstJmXDJinnfvnri8utFLYD7hXWtX
7ICKcRD3JlhC/5aMpPIxSRsWuILSTOiVOQUynmORBj3t6MbzSOxDnsXvWWc3
L5KCYGbTpc1TFgGNiuw6fsEgzPidM8F/TuUafLD4zthiGdpg6kYtZGJPCYkj
I5PXwlPF8mVvurzk7j45fxgnJPrbJQL4QVCfY16Sreh+gTg/KB3ehM8Dl2tQ
mdKFvdK/kNFXQS1pk6TmjFjF22Oso3143YAy6UP+YBawGgq9XGmlMDWnpYEH
DAYn2d77glX9yN0GqTE+EyeTWDMnajp1HMhNV8nHT1pIho7YG2rBb/JE+z6Z
jrygqctL0wr2a7XpzcekW77s7mIDUvrI7/LkB01rwu6w+c4opKnmFbZrqtez
RzIYi9+zgGQxQ+YE7OhpEgTxeizWEfDOwP6b7qS15CQ5U1xoV+5lkhSrNZEb
TKH+bPU+NZ0igzOH+9lT8Qr/YtnxnyFAurussuQAss7/jcjwEHN5dnE46ua4
D+A5YsbS3LrIr9YmNBgfZx519QaGPwCOFm1IeLGTpycBbiTN9uFGb3c44ifZ
+SXGJZJUEhTV+a5XmGdHiPpBGQjgQ6sxrJuJVeceRk47VJEty5rlTT6P15mJ
VRYah1/H5ZFVEklhcblnxJoxdhzHyk5d65DvdQifF5NUG3bEuBnORISbmnxc
7KH9MhMwP/4MF6F7RgrNkVv0xjkwZ4KEkfw88Tgp75RTWQQ8h5WHrpBTGMJP
78C7Y30L4IQfux36jPm1fUsjg0nf3i0e76+JIRbb735jlsxXNsr5Oc39XZ+2
Pa3C4fmAIJlf6hSqQfL7tDwfj0rjB7Q0g/YIhM5JQ2um94aoaXOogyV7fwws
Jj+x4JwMGdKHIzPI0bh9IvIZLjcL3UDSMJdVSWC4Xj4JI89H/gV+NKMVGgSn
TVK1t5RxT4oSkALsLVMIE3ZWTXFAAyBwtHN6wbh1DMwbTxlvKXsqW4BFWJfr
dfDS5nPZiNw+DlgEUEdGYS4fxKbTosr95ATFTk6CVftzo5zCWiWvtNb+zMkV
GSLkcs6yLd2Gq5uRDlnb6x7nZHVPSezmXzhyJg1RIJx7dc1so9JoFDVv9ADi
FkPfe1kVrfb2nttnhI+y5hfp/CMyZy2XPyXUWShDyP8eb4o0WwhwevkTZ1Cs
WANaAvW23u2dzny/4AfJoNbRZYSRsULlIrv5ZAavKrE/kiR8DBYnO7lN/d8y
mQ1vMxUPKR50bw==

`pragma protect end_protected
