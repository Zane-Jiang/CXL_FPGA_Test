// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I+mVFV8mcF7k9HI+xQrWv4rJDxMTMIox9wzUWEQT6ZncTdWJTn1mTgzTL1UT
iRFU4FKQVLQN6b5KwecziY3pmjG5K5UAE+CutlPWcmbayCsh1B7NPrcoRLie
ZoAIJk6o4gYhKsQ+gFdnQ56C2Le/TXGaLc0clvqus42XtTo6wOJc5qLBQVAX
dt3pkw+v2HLQXan/vTfsqacN3n3s7a8a6hdmfCqBh8E4OAD58Zc3lXA6d//z
XINiZxH1GVHZfCd7Pr12UJpN8sCD+HqfFn0qgcEW9SER4hOYsvSFYeHH0uKq
+ayfl42fhTNdgbihe0O4I7lpeUuFTDVv40qczA3GYA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pvK4Wckd/cfpD4yEQ4cHY1PkXgSEHLmzVpWK0c3mdSx4ybK1IpS0HeeTn+DC
qw0VFR/TLCwolxdNgSu7d5cX0uDo4syIU4wz7/8xRqGxkiWTQFbhoBDgCX4r
DF8tF36m43mZpdnZJy4aq1IrQ5f0ihkuGN09Q7UNF9CcivJAtnOB2Fjigrq1
sLIQKlKq/fuFxPazneopaUu5jlrGbTpdyFircLHSEXK+h40BD1fm5hM+/8/G
FHJ9iniKYp5ByrWRa/Dnrg/9yHGr9KQJeXBYZYfYFDUlS44GS0gUvP8VOstc
GhK+rZTRbq6gDd5r1Yc3fOOkJFql8jhJrCbQM88/hA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l9O63AcZtynl5/FFgegCxRIuZ0l9bdsnnG9yH1/ScBDdOZr95Fj9cEHK3jNj
u+6Q6OG7NM18NyPWA5R59mrzdTWiTMan7aEQUw/ydk3rN9E6Rjax4dktqWIG
7OakivUXVgxUMSD5AXhOQDjcF9EXE4WE09yQiAb+fwu+3KbQ8buZJ4S3/pJh
9kYr7ZF4viU246omFCAVv8O2e6Z1xWFr4XDHO2NsGRPg0avHZsmwbr5NhzyT
es1gJf3JTqs6LQUpHcZbdxnX9tciKYoInzdncDbRkOWstEWxMgy/qgiDG09i
yCrrP22ZgsAUoyyGz0m2+BsdpclYJ5/Ds/BGDMJ/aw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h5CzN13BzyJUW0IIp9KtR7Ub1gVu4CCsYyhDG3HG3iyQqyGHvoh9c8/dYo9R
gHAehawr95IbKLPQKq11nHz6/aEzsFnB+h0XubLOBal2lBk0heANCOD8gWtk
IWGSq0TxM/nWoLaLeV34ePLf1zae0axX9T+pMoYJ2UqH9iCbdsg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OMGtQuQXSdPokxo1emscbZvBQNEE38oMTMplYnqrCA4iX5tlLe2n/6JHv4XQ
JA1gezYHBmRXYWv0T5hSUWDgSxmo7Csa313cQGCk9bidQYtcqbQj2lCDoQmU
jgI3y6S0XAFtGR6ITY5uvYqsBlM/aE/mSHEb0Fw2MYyjMkRblV/1fMm/zTpg
Dyu1l3oI/9sRDGsFLZMD6RBNiIVcFICyzGpxObK5RAnSeGLII+TlmWv8FrsJ
A35cZQvVMEfuF6NpUORLex7L1gSMuLGbJaHPP0Sm1THdYWJaDTRQ/npA6bss
EzLvKYqT3NQ50UcsERxeIhkibdEPcejmOREdnzfPh+7mp+NZRsyplfUfVoko
4Uxp/VzaXeb62nraeSLt3hzGDju2fHmFzIvmXTynRdgeAlisMVoorsBA+8EM
0CN60DqpwReDJquCUJUALp8hMS2JSfKjwHtVuEV/SSqCWmwOOVLQ3jygCbTQ
Eq1psEh/mjPh2e/JvZvRjqWYiwKsVFYB


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EBg+KuJaTm6kqkaUHrLO1U8j399YrwnDzE8CH0p7KYGbesk2GQcuy1JFJG8m
OEL7ZVgzQGHuhUCKNubshyel7vAyG3qKXxJLCMjUP3G1KsztxgixO9pBmwv4
KpdD9kT4HIefTvTy5rfW0GAv6b9u5K9luhPvi8ruGGXwdx6732w=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fjtqZ7bnfoT+e6U5O/swcI4En3wONYlj9RvMxVotu7netiokDQ6mj/7hsk++
vmM1GVWdbdrcx5Glt5ncqvPO4/ipHeaB246Kdi380KU5Yxulnuy/A3x1wLQQ
HEr6vShtvUJgkVQ/GNm7XPIK0/qNP2q2tUUoSwCpS6uW5LC/giE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1008)
`pragma protect data_block
mCwcwr6n2p7wBqzO96ZIdCPAOgGHmFfvcFD1Ll8x0g6Bzf2qpnu1Mkg2XT34
Q+e5LzBTRd7jrz78BXb2rZ03pj1m6TU2aSpKwuKdfbD0cdfqz41uxRSyhGsx
cvj3NyBo4a8GF3xufyPh8rxL11dX53zgmqW9J/+vizUUIa3uz752bqo7WA14
vi+/2oorQEJGsXQNBNq+FC8J1YddOya9AB+v2wpl+qoQykL58XHMcbqeeGMI
daR+6cEskeim6Y42eAxXVRSpYbXBIyOAObcQ7jP1vbuGWmt7u5NkpY/ACozN
hWWIFNv8IHgrP92hfXQjQNwcLCiCKd9RSx++ZFly3O600j/kN9Ha+pwZYYyL
1YE/8HU53MfDdINf9G0eIZRsVVNqTh/f/b6HJV0GyQMAAWtmlxMiJyxnS1xD
/NbkQoi+Ul1cZnfPWKb8pnot/Vvydnc6x5TPDFKyuelaEIapDnKVzRkyPyU8
E3dei1TYnvOQbgzXA2nqq3z3Dx+KzrOM5fGGRDkWU1sJ9ufjzyhILWinJYkz
aEfZsSkJyWmHk+V/G9Hx/0Iw+mmY9qx1yc/oaYKY/iQxjPXx1eBIGNiY7NDf
9ML6lTKXpYf4Og0G8hcoY7WWpF3NAwIcayNntQfrgJuR2LcN1Oj8rgZ1iuoo
aNXEN4IMd28HzShpXr0j8pSS86b5tJdcyFKrX9TfhGSqu0QUyH/86V6SAffP
2jngV8xD8om84xWkUyE/Neh9BZ9P0Hf2vkJUTA3rCE0cHDieZrdzWSWQpM1h
ZVTG5EzG63evCYAB8GYbhUqjgMGAp3WW+LxhS3keNyRFVSYMcRRuea746Qb2
rzMkfqw4Umzv9xhseFCIY6xJsr7+yPvkvMxf/JD2LfuSIJmhT0p2WTZuL6Ej
pm3hP/87DZKQtVmsNLB0fj98MkcJDfv2RkSnc1rNgFOkRw6uGg1jjL3pucXh
gSqtSTvFyF/DkzC+FU4BC5SL2j3ps7TQRH7PAi1lmblqscxtrMl+1mj8ylp5
NdZg6LtB1WWSvkeAgF8e4F0+wTenEv1y8jNcINmX475JUFYv6zJXspRhXGu+
5ccHD8P9Ec2wofPuxC6lFU5hCtgn7oelTyUemldRaBW9m8lWdnKAe6FbiibE
yDOec5C5SbbfD5+KL+hlzaO1Qg7sWMR9pkBgG1y/s6O+LuFbcLABrhHIG2Lv
oxb4yBOPPikAzIkwpcONz0ZbLOV6xU4K7Rf/GI26Q2+Zc2LLC/jVtPVvBC7B
bL1lkWFFGuZRhDmg9i1075mVcbDvMxRuQ9zJvYWiVOwoZkTe7/6vbIBr2uuC
e/Qz8dMFEsgME2lJMv+ZsHfF

`pragma protect end_protected
