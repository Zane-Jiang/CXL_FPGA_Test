// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
SYjzIAPmlM87eMOWffXDy69fofOjCDN3JvRElBYDcJl8JRHaSjW4iFHYw4SvhYi6rjXGQ7iz45wJ
bJa95b/v+ngb5YJvPD6MaF4zIJYBBq1sCgCRWsZRRJtFAChHOq3tdgk7KSpfVCg80Lt5qvJGcMui
aJvDp35u8MXmIb6JsU64niiaHJIubITZSRlIOcwT+Kwfuzc4Xv1G6xBOWC1CjnjPp642NPIfdErK
jnbt/iV8VHbtUthfYD3pdDNvfpBT67DbX/2FWJu42fVvNTYOIcFV6+VfFAy3pX8gZosowlTOb1kr
OcS9jCVcO8x/ZzgnGYpHeo9xQ5SGWXg1EGDs5Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4736)
Alai3MnSo4yztr7vqKomIF6Iito8MhSFfCRsaZ/4pRAGv0wz269D6kpw0VOyfmAQl8Bt+q4OXsVX
HTQuSP8ebDj1vSGcUFW8i2npJSea82O2igWdbcw1L4S5YoHowi8YSsc4lriNfVOTlEl5Obf6ftuP
Yg50QmnUEYdZSGl0e21vl713XScR5IOus3Hw5L+9ZVJMb+gm2Fjq0QM+kbd6+4JMmfPJRiwGkirk
lLv2eX4ATFx2dawF8Z0V2Zn9KkQRnF4ui6qhBudDIdMeN8hi2koKZIleOQ0ZmxjdGxKrAbdbM1QO
mHtvS7mmMxghXT2B89ap56NQuXDHphMOuWPcIE8NaMyl6hrQHwStvgMHocXhgrO9lIWosdK3a/Ez
aoJWoeuRBY0w6ftt37/gVyVqK+3GYN34kF1Nf25L/3uw45zQ9F6+jY4qEjgt8v6H33cygHnHaA2O
hhZcOzIwlavOIgaV8ywBxlXEVjTQjlUlDe0GjIg/A65Oj2rRN9UQ1TJcSJJd5IsaexlXwGlVuNCo
2UZeD96HmQmbVqiJ4BCM1RwGSOVoogi63MePxMOcToJejPa+z8aPyIqywCTe8Yr6LRi1sDGQcKNC
0w9PPHyZV1meXZ6QTuBK5a4ghJH5Dzck6r59ST02jt5ZisX2MO8kiV91zP6Br2KxEeKaw4rS38K/
N/PuvzUwrZgqWM+ZXPx51pZuS1fzPcNPm7ZJIepgUuMlOeR6XKpVmbJRhma0Bfj9RmDaAhmaGJLl
e5Hn/b3kAuiPnqlZzRpJUyjUX69gncqhPHffqIAKjwgQgK5InHE/5MR+TZuiTbLYNDyNpAIhnqHk
dSgY0QPsaMR/csCZV4P3ofEl+xG8Is/y3NKUPU82uAEQw7aX/rHmGrI4PucazVkNCRX6x/VsIb0U
vHLzNRvbIvfaEjyX3/RLm4WGsLvCfg+4hBl7CQXJDOXbuF14yAO3Fs65tBey8eMkExfToCEZljqE
jT8piu0Lu/c93ZfW0TCZtO+zIG4DL7MrEFZNAzm6sgpmJ54SCWBfWlbrKFNtoTzRgiOMJPObZA1B
HehQBXEajfFbZdvteirHz0SzmANvANAlycZwklxfm+/FWhubSgLasUKwDJEhLDvcwjmK5EX2WazL
3IdPQLyBQIpt+mYpMcSVMNg0lDbigbuK5m5UYRN5t4ncDid7rzyjPdxIslBhootUO+6xdYtSxmUT
YINXW7DD6pyLT+iyE0VxG/WMuHe2ZSV4vbp7FgkxsYj+bgT34PEdk0oo6lBuecnIu5H0jXF9iDCU
zyUbeiXfoxEx3q9qNi9CDtDEv/bdEyrl99VeUqrXi3y0FBvltZf4qwTFCu3/5FGeij68PTQeoDp3
DJyN2FFItiLOfbbkUmYNZEoM8wO7uWFJatDFPHp6OhXewYUvrHHhMU8ylihmZKSfy/0RNYmOvqeX
LP07ELCk+SGv4WAMJW9v2+mhthLNWTn4c3Qo/va4d0gn2wFq4Wgo8iR3fP9Ku2dfubSauGYhyz9u
Aun5+jUM/9QmfjF/O/bntNLe3FZHX8hKF1CSmZma9APAzvPuMljP0RCu04J5DVAp5a+d2mvbCjRS
P606dbA9u67iHjU+9Wi5nj5ilGyrhRrv7OQF8FEWfGklErzm5xH+BV0a9FQmZ5fIJruRuzKqf3X9
vQQzuknpSNsJvx5bKauxOe/yjileTtdTw9vHC9cSHI+vq92je7n/RzsqGpLyO19RxhLAJ/59tfkU
caGFlBHnMMEnjHNKq36d+JcVrSFbrBuk6WDGzB4obzlDHGeikYywb4oQ1i2so7hpotlJrIrD9y4j
LfyTo1DKSmvNUhNZAed746jA/kBy/RS5niRFsmOOl8VdpLclxNxWAdjxD1az7yifUuic2eerMiw6
xaOe20cz/qLwEjDQIWB3iPlPYBavnZXSBiDiLdxgGNMrLJkbVF7k90sQ6ThImgWlJ+KV9sqImb2o
GFA+7ht6fjvb4DhFRQkCK2rVK6g1wjaqbn1DWfJcEO/NrxyjjLCYjLfQ427IkVcF4IcGcbFT39cU
/r5zUu2ux5zGu313hZJLAtEgBVOq//iccKox+ifKIJdhowNlJnlhFJwiseYtiXbxuzCcjZ/YHCx5
zzZp53jSIN/sq/27pVj6v46xabn6oC+fqXVNUe4kBw0kEscxrIazSSYUmTTvfz1j7jutAkI8sOID
ZneA2q7tAVfQ6zs05r2gz3x17jcyWIdPx701QjluE4H3gUVy4C9elCiZtxg+lHOqr3ITb6Hy3rKx
RNare4GhiExxlzFhnTWOrCw12jkwop+fNpUZjITZNx7XDZY3+ZAQ1kChdEU4H7rrn4u3RH3abIgx
d90ofoki+o3I+YNn9/2qj9l+MgVe+qu0rQO3TnzQ0QKstJiP2KLflUFsBQEl+7WG+gz2srp/ypT8
NBnLwRI4l2SjMjjQtPs+SwNUrL+YB5Re3nGA5lwc4haNzp2PxXsD57Sh01B3RQupY6vJ98fEBrME
cWs3IvQHCgmx9kbGSBfsH8IsorW42Q7imCKKYHTH/3IU+uNDn3CusKSbuydswddu7incEKKKpJ+U
Nf7Uf/YiNguyXHWp7F2SX1JeYpXu6p9b2V71b0N6LeqGvRmhIikWZTusdx8RVboxc5SPy4phg3e7
ERnwjvxfU3QYZqDiy91oRf4XGWDLIrtCJ7iwGWsguuoBgzjeDfVGEKUq/opQSDCVeqJDMvh3z5Zx
5dwB9GT8qOfX45PZ4a4kzjfjuHHGX0lpcjCVSQ/IdhHvmvbL3AT3QgwR1tA3H78bLKznIMOyuiGS
4GZqueUYoXyglZGgk+pjOwnn89bsMTKJACshO+a29HChaooZHXt/zWrfmcivHqSkNUzyY5mnWACz
cnp4n6oVkHrOsiaScsq2V61Wj/Cis3sY70WOaQIsGJkhBnevCTyN/XjasC6mSIKNdDEpKJXdAS0n
+Xng3jmBUtHqCTBe1RHXCanEUwkuevxprgQuqDmsixqeZ++BSWO8pKrieHi3Z+CwOvNXEdu5ifqS
rKqS7If0Fbholr/XFzxO3+Tu9FREq0KCa7LA+/b8O9bGHVaPArzn/OwWkZLiYYI3Ae4o8h6b1rHJ
2HEUVnlQPSAPmLGLnaT6MLYxbZoWiG/nzQKdzTMflD+lXBgYmELUdY9XddW+OpZXQI/As+25MrOm
8x4mfyx6WUc7txB5EkyVOcqQh4ZSSoPLK29l4T5CMx62pSka8DkYcFcAl/BX6+Doe7y1j9QVxQVI
a6btV4yuwDdnJka3r+dKcDqn2y8qo1G8DcdN1lSrs4gUylx8U8rEsRPmKc8tmirTF1uiB8+Gq3jr
kgl/Kp2DGXvDBjNWsEZrMFtH+z/Gghi4FrHBDx5Y5LRpICtH5mxfKaaEjI4dDj/8nV+6rO9J5jmI
2UHpfzWAnqHTzoTFhP2ekmP3INvBkDsaa+EMDQ0eSjQHhXb7UHREvLxxZblbjFV5aYxF8t+mAhNT
ltnN8QRKG6K9Vio+6RvWpBrZFkIkvOdVLvh0PTpMqdTNMnavhqDOfKoy3UU0G0ZYGdLQQm2CuT8m
mbV7OgsEOXV08pW49iGh9SztruXzRJ9UDYSeo54B07nTLv6q+zwjZMljE+NzmbOT5MIomf+W6P39
EfkVXaFl+jfk0YBqmwLTu0nAMOUJFClCcEd4fQYGaLaMvzjf5TfAAPq3HjHWIMZV37h9RrIxxjlt
rRrIA0wUi6QlkZcKdeSCMKW+JlX3iFBjUaofzrahlHEYt8n1olgD6qNMazLDCf8vr+As5+/Lkele
ZixfTdzOQHZteRx/qv9wrHy35Iar9rghko2LTTG16WaVHnlFDz+8GKeVUmFmwk0qFyQOVN8Th85K
5ZVI0PSTe703g8/fdEJljABuVCqWRzJ2RNsxCeCTsVC8S8XikugTufh+ugKHvBfk1tZyVSrNf40u
AliDLkoAntg3ODHyF1TCJkN8k7OUM6mHoOP5Rrax3PIJKXjtiGKoYNJTsbuRxdpe5JM7y3OoEpci
vHO6SgclgYMJ14KWy/up2Td28RjOy8HV6R8E6Eg87tATRg5fwXyLjvenThODEzuj3i/lwxm0UMdD
m5FeorL52O/XdqHWKVB85Sr+0dxetBHIGslSKYxX1MJyueDyhQ6dlY2JY8a5O2CkXPMIgU4e874e
meVMzC/qp5kUrIWHOLRnGq6ijYMgwOBPMp2E1ZBdih4iL1RiPKAT/TaP4flQ4Ckyopxj0mukmqhz
fdzQ0vhl1yaice0jE3HGLdhSyX1f7U9W9ex8nbGNoJH8y9qjjODUcyzlm9ux0FZveEOjFxMZvIwd
cLKQ4on/H5O8nYMKdnDNceq6ZF2k/OSSsaE8eeu9s9DhpTZiG3WIHJk4GozVEIBQmj/e2/O8/Uc8
MR9YpKzZ/kxTCYfutXx5fYrmQgPvg1HIcbs90L6152W6nXFtSuW1vmsm/7LfEf3N4f2sH6MdZHjA
M7f/W/oWGEQJZsJAfaHInAEb74SP5wa67Jhv5Lu7zTnaR7rTRAD53D4/XrccI3O1iNkSWZghce8o
CHu8QREtKTf559/PIZbpoHNKGe/DrsVSbVLr3ylnraN9yYPts8p5rELyETt2UQY0Kckkn0N8QblI
3LHSqONIEudhJuqcoPEV+pdFyvz7CAWrgEjgXPYnvkJkVKmcftOmrZLUd9eW7xKEos55u9mAirQm
FALSfpfZN3/3UnjA92sHb+8e+DHxBpKe4dhSfExvm7RzZcW5DAC6gEU60bHDZlUO/q7+Jn8rC94y
E3XtH//8sKzgOSe3If6LKTKSKZAWN85OVlgaz9Gcj3We/bPIPhYKz0qANhxQ5DsqnnZZ08Ncdx5F
HSpUwyAaicyD2xS2WY6g99eHYODkhjGQ2YvN7lBCiSe2942iarlJZuQUTHOOdTDOSh2cEsJTh3HN
kClqh4izPQpkVr7g+kCiWQktZrMUdho6Od2E6PXdt/N6ny6AoA5qTE/5Cz8JfijA0LYECeSiZTwQ
rsPjuBSvIMJA9uoceC+qqKKYim2ndxD9eHdVhlbfgwIZeE6FYlGeEoGHJe9vgAVU1vTaTv5j39dp
0MkfHH0jbMJbvnKpDOYm8yL9csTPQcCmYcAOEXIerVPZ1OWAryllR/EUV/m6tL43orMAJKOrn9Xl
VCH2JhufPpg+Hv7Ys2aKqT0BRbZc7UXOBZk+TFaJafxHfspO2Tq+sVsBtDl086DWP7vLrPvyaQRm
tU+6JVs8Gn04m4HVIGIkzNANDt5iQ8c7cry43RdUWOti2VnEjzE0lKusHkQDYxxtda/I2xlDqp7B
a2MkRkE8znBpbgdV1ywYd5hNBorbG6HeoPGyEUvFp0B5mmyP+8Nmk2GsihImkzTMV9olZzI1I4Wy
kx1A3mdp8eDCiS1n/B4EuqVN5fVs7lmtY1Kmf+Ibkq3czy6HgODN6ugfge3JE1YIcxmH/n88SiVD
bP0AkUkI27ParFotIVDf/QcSWqm7GVxUKP4bWLnaTeZos2PwsrGJajAfTpoDCMCGt5ivL15risWa
ld2EnsE3vkDb06EsnBepDubqjtHGLFCob1lRSC0qN6RoRJuGqdSzNgimY6+aCBdPTnr4J5KjgieO
h/ilkCSi00WpOTLuUS5S+1S+GjItESk9qQFRm6+DEbAsDXu1wkcWhEDyLlz1M9uUQT5rh6O5p6/J
P8BxvPAsNwUgAENuNBEDuz1NRCyL1B3TDRPOwNFY/qQpWXi+g/tVkXDY+QtrCXWEd9LSvjc/pxy6
LrgEBspCsUlvTpQO8WrOjSHQ4rNBQdWqLbpZbbr3Mq6HtBhx0QaT3rwQpuFsfv9yBr8P7eR5gk8a
uHFdi6ZrKRBnhivd9wnX9ys0uJBIWYd0QshcuJplUjPLFtB6eSEtgTioMqzm3ywuZas18Y7MBBRm
5PXqiQE8jYq5lJQHQ4upA1vmm/gZU3Yqtepr9STKxLTQSshzU8u4ChKUkHSB4KT5kmrFz/ZGziSG
JXnLLG6mT0uGG8OyIUo6OlBt6vkknCbxUi9OrRtS0cygDEnozz8vvtF0ub171rvTV2sMpusvOWXD
4UZk73awpMjwaPT9Sc1lLIuf1ksqn9JpLE0B+q6YMAT5XYzX2F3PHCEeoroOC70qSPt7l6ymlezW
ve3TonMFJc0N7PicMfdNyk4NTj7ufjn9VTdbrTfZawioYf++lWICF5lNumEg6kMhWPuJr5JQKK0z
6tQHFU2gfxaIw44ZAIz4ovbvjkNS00C0Er69xzz93MZkF+E1BTbtm3ir1f3hKiSQI4ULZi8IFyYv
6SqRQZo=
`pragma protect end_protected
