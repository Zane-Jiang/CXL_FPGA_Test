// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
VhRba1HeWIGK0ZQ05gd0txpGgvYDARd3OihvroMSuH3bdVgwh5m+g0u+TXk/JwTB
yksyPbWWogJWl1c6t4wwbZ2zy0VhczVr4H2boqmuNYVDHR1MGAV4rfnq6RIspuV4
+ynIwV4N0fNgM7sP/YgAmwsWepaOMim2ku3QH09QYXA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7040 )
`pragma protect data_block
QBMrY/nfR1zZvIzC29XMiraAxkHhAv3FTePwAsSmKGNZ9M8YwhPtxsKUi57KIYFE
P6g0MwtPDCZjl/friUrL1n1t4gRUZeuFksxy5qF7If1feCOAINFz4xzmceRwh/ts
vNrltBgYHbfQmmL3D5MmDHyH1kKVZJbvxt4jD/l7xr1NUP3NecdmXvetSrwp5Yx1
1p13bNDSkigae6wNJyynufn/tir1JKdV8HWwB5se/BnI0818dlQthwxD/3CGFCEK
JjPppCrYy69p7sg0rhVFQKB2+7bI8LpzQCIqbqDhgIgca5NyF7AxopSiElRf4LtQ
YZpyZXKNSK76Gxl8pNd2RUGSTrKhM4Mv1zSdZL9ObXgCWQ/E3wnqYgSY/Bl3WrzY
7TzVvyw1F6ejozrr7mLfm9NiPUjcye2xlqYfAmoJ/L4fIDXSextlu0PxAXgiiUUH
VdwfsRlyTU5doULs87wYO2b5INS1/cuI1PG3faaMBFD9cmDU2dpqkdK83MXMP10A
mj94UxLGYXaieZDKsfD5WfGBPKw9M/sB/fA999p1hfYPmAiURGKlerfLpjp1IXfl
+3BagsFzq085O4rrKJq8RAPf2zlsSLwK7Bfe5EXIPpcjwkjfjD2nbZMF8LPqpW5u
IFS3HVgFaIvTvv3SWWTW2Mxryy1+nWVchfy34Cp0Z5BLNSoXGmAfKXDnYIBMTv/6
huYNQruf+s+/d9ffiqS3uwgpOC7eU2hT2jqFwww+X+Xcko71e/1ExsMknOF14gBh
2BfANoFqJqaZy2v7qJ0a+6qFNeDM8UXFpK6eobG9OQONu86rS+tmF0Vo6l8R70DM
52PhSirPDvqxJMpeggsYAPAckDeh4G+IfXHmRpb5c+SBElgb+fZTz8/Af9MABDkF
aq+6x1a2KuiJuYHJ2VdKjt3CoQunNjy7kzUenIfF4xUux17y62HEWEiG3a1FJJHi
FvNWJOD3i3jJK4IOG7eB40DdPkQITl3DEzrXj3pqAXb6oVXJJLOZL6gfhcrCt6fQ
evTaZn8H8CtwJye/CSy5dE5jw4LC2HL6B+3ai3I+RgrTjzXxx3aRBgG/4cvIZaBA
uCg/RvfwGjPnnEhcWdYAnW7hIXWE52to5UE5h7mAbPPY2y50rCOLbWxi3L5CgUoO
Hq7lFY42h1UOgtO/0faebOrS98qszumgLhUxKpjlcVCgv2+SzpnHYeREz9yRDgbt
5EFmenOrTP4GIWG9laqDCoViq/QFSEF450945+SHi3FjuGX50eco+exkIgvenNAA
FbEmTkQGZ2fZf8RhhoucpBp/LTOvEhR9FVzeLr9AmJdiMdKqBxmQt36dn0g0LOas
C81PB2IubR2ALFHA4YztQZMG68CtVVdVI/pIDMRImBguI2DwBl+CEW8xfVz1Hokz
0Tlr0b1LI1cQxhibd2FwOCBUViPh/QKHAHnds2Bs0Dv40pm4t19dNVOIdAQtJk+S
sT7RwgOGq0do5BshaJvjHKCrOxEMcTD1PUQ8SAQCxM67/2M3DVXMxOLA3XAuMcwJ
m7MB/m3OdhWdgdOkua/0Bj0q7tR5P/i7kex9Q3+v2rpMJxoo5K6+mT3KL/8B6GH2
LW301tx+oy3ZwialTLfno62F9tW2nzLrSGXm9kD4NhtDSEVOrifUK0C0HeZcewfl
t0us9pNyL5MjimGVXCujIXUvDghrAD3y2uQSCcSTdR5N3MRdWHOYXVMxDkqoMk2G
PfuoYNso+SpeHlIxQcnE9zW+vklHRSNN1V0Pc4Y3oZ1ftu9yxzb+6MsyL11GqJP2
E92UIjWzmzgxHGKhn9srKzc4aToPd6Izt2Ydih4S97qWNGOU7zF5qzUIf16xur7L
gmIv8nCTTg4zMpE0mRZh5Xpt6ISLpzPXrEuUmN+1ThwhLT+XiQHDtpv3fqW5TsOb
pnKhC/YVSOErdXe2y7TXU68Ttd/AUuEHmljuNj+M6ThhnHpug8BInYJOc1KIvZjH
ZpJODVx5yhiQkXxc/l13aB/uk5FoqcyqeDJVe1u3UcRR7AvV3bJJVsRsX6GHATh2
gBeMaMJFUIG5rJ2iodtNjCmq1dZbA2JFIRvUruWFhNaH+J2JJNDekpYDu/pbeatY
z6syG5TYt/c4aXn2EJjpg9qNLmFJAsTvasPmedGthj0mjn3sOJDOLf0ss9E9oWa+
yhBEWz0yg1f0j4pAEmanrmQKJKrHJItP5+0/6pntSr27F/+junRCoDUTM5dGXu10
nwlGe0ZQ9VGMzRDCKDrC8Bcig05gvgcj6IBsQ7ziRGt06vigKp87kPlKGWzDE/Dt
jTvBiKn1XNvNdeSf1yXka/6gTrQq+/Ro8ucIpRY66B5r/2Ldu9T8iGiRKn3EXEHg
TO8bcurXLhSGRphzyaLuMH64NVoH1jjZT/1V0YC1tdMd1Kaxe4mQ92pA+EW2DSDJ
Om4z4/il+9GXHD0uqBCPLbUQKj2OmquFLRYsIX5LOi41oXTmmwWWpA00TeYCIPeJ
E7s+yfRwLkvd+R++sg6fOg2Rf++7Wi+M9kD21pk8v1aUO+nXtjiN7SDNfigGuSmk
KKz2oQAFMGDCOa3aHD3rCv1upRN1JRYL7P1KRExP5w2u2xsNkrDxfpR7i5xLaaoZ
AvFv5pkqFjtiqF8OCJVAKlSiDW9OrCNcbFDO9/o8k7MMi1g318axfhv+zvKUoNj3
ZhMxXmkiw+zagn47YzfHlOfFy6xQRUSUzdKMJFYWrFs8IgakHLMa4+orIHz+aXRw
DIqhGK4oWDSc8X4h5mrBJhWhhQrnGmGjFWfjkTVqkIapwa35kv4LRABRZ1xy/i4G
tDbfdBWPLiuj/mJ3EFRzDzUYAf9pYRA7dchRP4hENR2Ki1TVEqlE6IY++236sGgC
E/l6iIHQJv91OR969QAB0vU8FENCPgxNwm9haVukClEbLrzb4JdRjZeEVcyWDBRk
N7dgY8i7dP/0okcK54Qpj8Kn4lvPp96ja2oyBH1m04xt50sbQ5dkTwpXzo3/PJzt
K2n7zyfY4VVy3Iv8E7MhhqaGQ5d8yb8aiF3thdQdKzD1bkNse0HLhcDo1ywjUBOK
xQOfjCQpz6ov6v/MNoPX3iFuAP6gF1ZpH8csJtYTcg3rHHGzpRWTTzUaeUUaea7/
tVnPj9Uv10c2tfVxClATSQv7HaQLZ1OKe7Zi5wbwSFWW9qAJvRzvNXkYszZLqEEi
fOGtuK0KkqzbWCopzZpLNdx9+yOQhZbtN4K2sBW3kUtzl58pck9ciKn2HJuOSUN2
PR/OetFbuEwzHPNrgwq0w4GOSkamrGCHg2A0Qrc2B2ePCQfA972EYXg3IvPX6cQm
50WBGsZgtG8Ysby4To7obBrlTsH2AQXarBrz5FX0ZOZHqtNiQBRgiAG+L1FyYGBs
++qtc8tgYmZ7sB4Lg8JZPi68NuqcSbMCd//AHa3xAw8U93QDHY3empa8S7yhavfM
hJ4lLla88Wamu+b2MpoCaGsMsJBcm9Ykg/wyo4hr3IK7qguxdVuKlQyAVdSkoOa1
8phcfZ/FTDEUXGBnFx5J5/Utr4cVAFdeV9iaw9X9geKGPfjRtS0u2KW1oTvXyKZ9
hqmyHL+Gh93oJS1zdWavldYKfBNHS8GPKfGaRuwY5ltUz3y2gQkXLZ8WStGGxBVI
KiTjUNn1aKhO59dqSKsPr7amVO5OmSvkqqU5g16fu+wBoDrAYRelsBgE3VYeZA51
3srm4AbFE5nGQ0VdEF7N/C+wix/K78TCjiwXAd2ep+g1xtXJQqTMR35NpRPd3lXg
/w0sfmYmpMUAxoRj7MbYPlugX14F3oY1LER8m4YZ+qeK7GOl76EbzUrcfhtwoO6w
TVX8HHihW3ZcPxCzeFNL6+qaDsFH878UcHKxxdOWKa0BA0EkhKCziOf7bGSPtyc0
zvXQL0jx4paidWNw38XOf9M0kW1e5SSjdI3BgrJpS4Fc7sRNYgD5s8ZpK54SrxJz
L+0bJVbpODZg18HxOD8YWHVW5LTAhXMt0/dppw3HEry/E2+TRgP2v6ApuysortZL
9+L75GPVqC2oA2DOXb3/h5b6jHui13si5VwH1DLxw4MYaZS/zakBxRHOIwCsQQr7
TZLB+D0LLfjnOX++uib9xyghW6lzIfsBBhcT5CumqGbypQdLPJL43HGxa1MIehi6
NraP7Wrytj5hmd4zlixM3aeCPCNVZ4OxkEBCzG6dL26/KmP3KByEbYeMAv2ZwjU9
9yvWjZeJPJDYucgdUufYkJ0jzZF7L9TQyD69M9OOZeOfUNowQ87+yM1WuqFS5pSK
kU3ZwZI8ahxWAlabfp1QyOudpXFzOkAQxqX5wsD8A+8pmKrdq/hw7cua1QmCswhO
g9XpgYrLEMX0msdujzMVZ/kZbHJNb9OtWRBqBWJPFBQiAyqBV7lQxVfwyOGUXfpk
m6D0o7VJVFelcfGXM2y2T2JlRGlbOnNqy4Wn93yT9ykh8ToamFQh4mw5ZMPKt56E
faEkR83TrHQWzSfTQD7cGFulXpE194LcfeE1nDEet8qwOB/hBiNisu+zMxq+S/q2
TaLPHy6NtJVC7PC7609jRQeHsN84nQVG5qvPEIFHX+zvLLeGPytuFazfPILnBFI6
ts5a2R3giMf76i1Urz3Yt1FiQi36654iJDxk5TKgjF1svWl4YL2N4DAehoVX3K3N
MQprUEfANOJH7FfKv7HDs740GzJK6Iw0B5/TB4bSEDqoZo1LJoho6CFl1a8XRck3
/BNboqD6byCNLH+uPrjEUGyHhWoP5+9cytDf3SLL0vh03jSEVAgo9oq5ncgZcLJf
0QxEcpMW/a3abUuoT4/NYxEkfae9rXpjunxyf2fJFlaABD5yxZMC409rwxHOf1XL
Hmt8/QzbwpXQMbvj8Uq5/tUMcXFErvfiZ37BNQmN/pXDA863dBvMJvZ+xpQRkWGm
H1WN6hu25dcrt/DYFq8CYx7S10S++pOtzDz0iM8LFtjeh2nr3DcrSJnD5kTYukK8
ONOShVszXRb9bH1NlsVJJUm5PrJ5v9gQsejPyrpcblWFj0XOiUfso7LAjK44r2ae
y8XimhnNCz7E/zmN412o7PhanXAcrHnE8lpzlp9yeeXtc29TAfyRkLuBC3OPSYVH
EBsgJZKJsnXfe0U5LTVhdP7dO+IZvD0t2/fpBu5t61nKANMBeKbyAYFwxA6KheTP
CKFxNvltQmaYUnFBFBilAychpSmWMuzTCm6XPa+6whpwsMgltn+mLdqNufYK/sve
8N17VyARqyeyoeWagp+aewtYHoqGsk/hO9Eyw8Zzja4T7tUz7nwIg41TdkHx213v
xeY7eJ0RwmtGSenUKGJsr7vJE1qbnNEZaGG/dnanqZqbvkGXighcnOP5ONjr77Fz
JhrRDY9ZWJqlRQpI4AyQIkcB8+LKxM/2Heyatgg1YmmgTH2GMUJTqjJuGxYG/E2i
szk/V+VvCrXubJ2Pvx/vibbFKsUIAXf+bqRNMvmpPHuuCFUdWPSlYRNbmvK6tXqC
SlzQRCh13lZmYllidXLk6C1Pb04qicyRXlh+oz7O/BPpZJmDITHIl0af0JJmxdrx
xHUMgu6GNUT7Y1KOFkfCO14hYNWjsHzzSbT/pJlrMM95OBnBWcuQtC9tIk7PMGFS
KbaUEHD4qXrTzKVieNN5VqrYLnB3bii62ERzNQZa0RRMU20QrmVKA8ghOdhC8bO1
hXA5yYtq4oJTt4gcTkFAH4abilDUbA/Ch5H0kwTk6kCugbP1fF+Q9wvixWM2gv1S
/uSh7V9j5Wo0Sn+NGQ6+LcYIdJXjsFWOs3n9ZBOH6Ovpt4V751e+CHe+rBlwG7Se
RnReFbKHBZdg7CapC3HyZtGZRyZbqTa6btO8lixrfhfFAwFSwPai3CG1UHgz/R13
VsuVEJfriCeuhqxml8SqXmYFycUhZv7ggfqv3rL1GiRvuzjcHM8P1UwLhIF0PTRB
BP2MAVJ8bzhjgDPv7o2pzBmkCsPQ43WognGy1SlYsrH60eDpBg75LeYN93eiChtV
ynCYG4IQlfEDNlrhTXixAzWHe0xEJ7BwZWJzwfH9JHProvKqi/lSUm/ckJFPZVF2
AUtsoz64EBPc/BIqcSbQoQeR286tFkq0c6no/52xM0UNEC2Uo0doJtPR9fJkPscD
mXWrPMtpuYxiD9tFczgsfOT8k7vuOaAQKBdu718rO44Mf5tXVSOxweuwA0Y1u5Jy
6DakcM8+Z/Zread8xwYwVYWniuGD2H2nJwZP63XqbGNQLZf/B7Qtu3N0cdaVBnP+
pWENw78ZL0PUNX4FaTcdbnDdlAKfkqmKOXKVVMaZi003twalY+RXJz5PFQBHTfdN
xi3tAq9M4biWJFggGLH3xNz8yAbFaRgl3ysgGSuWqYCRvdFaqWHWkDPt+M2sWt/w
nVrYsH40HQ9xjZE9lK/f/K4LPFiWdA3Lmdm/T4MDOYKbTm/VgFf3IT8PGo3A1c82
SmAJwh+pNxDFyRIxgRNfYtGjCXxWlDGqqJ7agiolR6zAyHU1+wXtf+BdpUupZvzc
WkA27pRAv8LE+d51hA4QtN0oFbNl0SOsYXgKMecDnTdOyxrpdpWCB6AUqKaagdTG
WI8ejjX0l8l1MoVANl8UJBquOviZj4Rg7GO9WT3yElFpQ2Wcwv1s6E88b8OmLnKZ
VlSNnWGEAvqG1GRzS3Hgn60y0Eth/qOqiZ1r+qGbIASIzSZ0VsSwW2qmRoDT9Vu4
FVynsR5lzSh4ieco3dgQt7DcjC0DfcTvm+fG7sgdnLDQZC0xlWkki6HtCY33AIUK
TN+KCwibIFV+ADiXhWjjg7fSx3+PbFBRtSa3bwUvPiOZu2R1bHpQDMXHZi2nqD4m
iVGvYIRloJOQ12U+kRrypwWwzrj1IzmWZB/P+gAa55X9DYsMymIuCXNLP8j0jHCs
isUtRprvSq3i1PDz6A51+RtljtUcFEdJVi2peWjL5pbVFp1UzlxeM30wJnTbRrbh
ZV81i/szU8We7AhNeJXkCtWA/R/vUDF533Njy5+0pil7pSm50AUuv27ErTgHKV8t
1Qs0wNVg4WE+Pp+JDogT2R7wbaQwBiszJbS+9bdrJ7HXIMpEHxCp6isBf3VzEeg1
Pb96qbMTjoaUId+elAF4QCSj1JnQtUaXxxGqe2uDr7BYUiHc4Ivsko3fucCAGdw2
xb4DQ6hzKTc8oOe/UGs2PRAmBRwMavFhaIcehlhC6dWOX3KOO5hvfg1svutwzACx
W3ETsSkUgZncdssjYbJA/U0ezwW+SzO5KqordAC0/Bki5+n9xpMMf7mxqYwdq6WH
FvYqLsc0QPeHEyfwcep6n89qgQCbD1V58rlpuiHXG/PUVr0WZzD5ImzKsc5Xc9h3
7YxkvBCErPA37kvTIOmUkPD2gdNQ+x5rZ+nVBGWyxEQRtKb0edOec/u8jG+QQuak
msbwh2dn0WLWYkgoZwUnujjyKETDhbCZ1PUNtBPbELBwKVYS01RVpKNJrNUParG0
V4N+3AhyklcKK0Sjcu7Jrlsj70aqje8nanOtfQSnC85kyPX2Kqylp3pJ6gTB4NHj
/UE2cGg2oo9Vd9yDpae8eYKWN0MH3vFBOe+JF3AahdAwBlPfUHliSmN+mA3x8BP+
24aJ546Vuf4WcJNjvpaOuWtxHlE2RLO+jrJdpewKYuLbaJ+SMlWn3GRbzJiw0rNS
vzoY0cuEzZye2NiDlkNwjbABGBznoEtOA0pZDETmbo3tGFDEGYRHscso4I30XghY
DvtoF/HESsHYBHKHr/3CfbAzl4zTk7VO4kPlXqdEMYlelujuYo+zzebsPa3c+7hx
XZO0GWAQyydDBMqhjH0SHYCnI9dkGrnjfk8GkfA9KyKi9kvsHMXhZ0sLUCK/k3ne
VIDzvdvqdzSLjuhFUFlF2WsXuvrjc3kwtLWWUlbF64GQIQvzSpFWnDNOPLZeVu+s
1M0ipfZFzfBME6fj0Usm2+u3+aXlxCi6l30jRVpi3wh+b4gfnn3p2TOrpeRV+wxK
KGQj5BGe+o+MdS/ZuPEwadNi8abzPYnRuxN2XDry/IgWd84f9TkZvmlxPso27tRh
zcZDXvE8Z2j81lWO4S2lky3FXBz9H5m16LgBKYSbCRBQ6SEQZSUPnohJqayiWp0s
1Cx2m0uyDmcSHolilSDj1mbb1NmXOsaT7Rbb+qVcuRps9a0W+kXV1X5UTwbwN+Bp
ki9eaF4nYxBfkvUDSOmpE6hcqcFAR7p6pVvSBDIJ3NoYnBU75N57WQxTwZSXFKB7
esFKZB03wVJd91GiQOuolyJDHavOJMuKNfa68QVAJJjLCwUrvI4A/CFDT+jP6hLX
FkFW4YQ6DAiKpmYmMVUIKMwXDX13qjyvgi35tr77IBhTP3vG5d+cKMg7Lr4HckdT
i5y7qXQXXrn09PezygMpdcvNuDX+k495yBXjZeGZ+Tpml1ft2Tf1FTbN00FMXgFY
6lNWEsqLtRAZFW9I9HLYkX2V7hQO2lFRKfoAsv1Owj3a66LWwpBJ5WmtQU1enFqG
AeA3ASKJ2uZWD3bN9CLpHf0erIDH5LtHlAM3YVj5/MhNv9gVZx5wOhvly4wQxy6w
9QyOgMCMe7MdlnIRU/CwHcVtHp72dwJ4dp+AS4EyVg/FkNwmoZRD0i95nTi1rFdT
w92q8KszV7RvxV+wpFCuU9khd03l4JIl5kCMc3t8H+ECPk2DRff/H+/lMl5J6NoD
YInj+XkNfTWjcj0zfl9R4b+GhZo+zCXMY+/XAj9BII3pshoXg53bQhJjRbwzTXjq
P7JK+U8+RunEu1CgMtiktECVfjTMMEzPWFiLkwq9imcMHD0Cw1O4TRbn9WP4LEmg
gxEkEXQ5kKOc+4uN5W51NSmGRhvsRKCDAKgMVKhrQPzUHZmf1r3DggOknDdm2JET
uX8P8ELLzS6YMLFMo/Z7EdgsQk8K4eR5PSGTy2AvgozV7gc8VzI7iZ4o0CjVNMuM
wAj7Hg66RakKBmRuV5XenMUpa3nDB6macb2Kl/tHkueOCZdmh6GBMXZkrThUZ1Q6
UUn4Fsx49FQcF8b9Lq95WAgDOR0EDH9CX6Az68Qy9znVorlmshv5IiA/5C7DT4c6
gwbCuOLpSXyEKDmQDoTxwEt5Uvq9loo9zzdlDAu2XHb3rwQvgxS7RtYbazlYk0Xt
W6Cvb+3aCBQdETHab7+sw9mGrrCwQQdw0HxJ8VNH/JKC6LgWntZlp4q4mHzyw26k
z1IGO4ZzRt6P8BGlOXygDVJhe04K2B96+GzibZtJUv1asM572uu4wBnP3MybY+wP
bo5wMkEKv0RgGqLD+7Huvyk+fyN7yRszvAEshEwodDpTLZqLG7AUbQAbM+05l/Me
nTHUgnWQRJbjezpA+j7GPcgmM/Ny/5fw6xiagJq70mw=

`pragma protect end_protected
