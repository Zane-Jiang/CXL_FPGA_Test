// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
XoFuXd2MRdzYoWLFJbEebYQV1Jk3L4eH+sYrLlmq6gf3AvgUzIvof+Ety1Uh0S7u
B7XthtViCjufq1vGvlzH45axZhnVd5F11rPmmpwl8b75IaGJV7rG3vv7ZSAVt2LP
kYrCMw0bGECJ0iC4PLrKt1EYr5zDLLGBPkV3QbN+6k0GXC5VllzMDw==
//pragma protect end_key_block
//pragma protect digest_block
R2iFOFLiWJAtqXtxw/bR5e+oqj0=
//pragma protect end_digest_block
//pragma protect data_block
il+FHR9YTu/oDwhP1/crKqRUUPgHmPZqy9BeCEdwjOz+l+1TvLDgeDStT3OtpIWM
oVUIv++Jc6Gpmg4DdvHkaRRJm9+WotascmCQa6oJK3i3eOk7m1ShuqFeIZe33UtW
KTrE9Js6KPhRpkA5+muXFvnZkvZoBLqxgQNlC5MCmkLe1rJhHPjy7hu0WU8aTHDo
ymkn4Hf7t6JRnfoV4k9rR6j48FgP3X2tZjISiLyyW5FdLATQawvWBEKrrhSFWiU4
8XEHDnhu+GqfXYjnDy58YS8DigD4hFN+B76JOMYNGGGOFAuXU5SNQloJgZmDOR6j
Djmr1RvBRWmHphgnTeTjlBl8Mu6YL0ZsZ66Kw+IpuqeQ/Rzv37f3SxxoDTZLWb3/
97AaYSOoJemPAFsH9or+fFVe89x3EeLWoNMUyHGMLhpSLABSMJrCcMZpxxZyQf4g
vQCrUCV5Lv9p1fzPdVlc4H9aZ87EbuFRzrcaEBE3LmdBk7ypjOx2WoBwX9NMI0is
e1Qt9qvUOM0m1VTbuin/+AzF9yWvrdYabElMwsuUo6kgxbBqPowgVjxAb4WCZesE
5HDwNxTt1t4gW80pzmGoahVxMKdVVXiwtDByPFrwSEZHwxwPhHD6IbYOO3w5jHkY
EYtpZdIO4t9DPF3a3l+rxVMhoVg9mscCVHfkcUASGrUb+ins/2U/vcUFbUs9BzWv
vO0blHW8O9PvcCUz5Es6hBEjzjuB/kGCCprk8wKrdaKCUEWjJ3GWDKl3tatDoBMS
u8dp1SG+DxLrljF7E/kJrTv6p4OhKTuHTrkv9wii5FD/fpcwbjvt8n7m+DUcXkfe
n+1SNdZlc8B5rq+J4O0DUb5J+VCLDPEnRRPC9GgqPXtLpLtsdF5AtjP/eV1aiHS0
YBej95XN/9Z3TFLJgVVooLIO45D9jucO4q9wGPKL1ryYVU/pkuUrE3S+tMzFpGOA
ufAOvTd/J26TfB4ocVelDZzaQdvqJqDrf4S3bNSUxh3I0syfm7ewkNtxi1LRVeWS
hoCyoJ1wxZN9Aj43FTnhZYqr8Y53E8VYlythl7FGz3TCKROVbZotvFz+tUodnHOK
sLYjbysSvgc/+cE1uEMzn2M2ML5NQcWLRmfY2yRbAdPHhp5t5fqtvAgWEszrJ2CY
xs9Z2HyGF52vMBdKV9F8u+5CdHzxf3IeVjR7BIr0hAEuPRG3CFBBnHP/oHVuP8oc
TgmGxVF3+Lr5s+i0x+wE1BMgfK2/pGtktGd6kM9kIIdltCGUjfv+bajb3e2CPLUg
MGEfoOg+f0zeAiBD5jOJ2UbEh5KYItvfbRLiZZaE3jBQETEhegMpBLAIB2gkAyKU
89aWKBbO2Bx4RJ6UZPr7uGryQpyRQEEKoDhMDxCxDRd1ERKRqpPanZztes6Evmzl
TtmLlW4JSl6pU6GP4K3nLMMCFXRd7qID0ZwcpogxCBLzsdA+0h2sVsJyCgXxAm6I
ZnYjQ4fOpntjupX4I5BjO1IBX20B5gQ0Ve3nwO7tEUTjmWfSOjJuH6IZPQ4w9mmH
mGJ1TKV6GO0lEtO6z1YAhJc7C7ylcknyqDS6BBwR3cgtfTn/EgZwaqq6pCS3QHNP
qErhxXdp3hFEH5w3/aOM37u7MHx3Wt6EhutnzomgNjknzaFxLIo0WirmdTnSiiIU
HZjD9RqfYScQpdOJkrWu441OUNByeUURENkV/ucKpu04Ss7/Zu9pmeVwST/Y0BXJ
XHZh91YRozOjHtJo7UvuHFSAageXMCZqPlMNbUU96Fx6jr2tkGBuDw2S1TIh6NK6
tLTl/JkzEt9zjIQrtCqRf0Hq9RSzhQ2M7ZVlYPzk5VRwQ8qAwL5OAYSu2T9UW9On
oue8Okc7Qu7yhMwe+YdD/icIsMju1wVEmY2pbR9NPzWfc/vTsUS8ioYmC/RPBkvR
A2XfXs2SSEJtPBtMn2gSHUOggnh3EgeK5KJMenTCbmfAXaZKvM2fTJp5ZSu4n675
0aR8MoKwZjDDDcNbc3+LTIPYnY4p6/NEwza4DcgBaEp3lidfsZ1Ao7addGOsgh7x
rpSy6lNR0kHJbRYbwc/DyrGjmGBUkeC5l2aSMfGrfL+Ru7YXf5AK/5Jt7DtITvsL
YzLQ6Ru5gvUmWvFfD/9s9X4Q8Y3Pca5qwEZOobqT3yD+UH+CxyK1Z3IHPQgD6l1b
SejBXhSGiprSvIofZ59rYMDznWexe2bWP8tX8ub6ZvXSzKrx8HKbUaTDyo/5bdhH
C0X2UJa0A+gx4dPIF7uRskCykhBt4z3khmHAJRB0yoAF/6RH1azHqWdtPAizyXti
cr/ljMCEVEOk5h944cSC/PgWWvgisvJf3tOwNdUJu8xctU2NP/SI9WEI5W5IDgwk
kVLBjeWNqFyNTkuE1Y9aHBaSid3wAww7OSfX3w7JIOsXjGmmrB1J9IMTOxGIAct6
fSCqBc7c/AQDA/xa8YlG8Xq+Yf6e0HEzWLxIEElcmG3fP+zVqeXdTcyp7cyfYdw2
QtDdnpttWvz17L50CQe7UHD3tRkLqSKZYp4VNC7l/x5iZm+iV95/yMYOC4blmj8D
Q8EVUUbnJjUIpMLA97ITTk5FM4OoCYbaag/ElsaB/1pFZ7W7KUzhZ8C3z4yRHzrC
qu9izejMKmoJsDw0+4MN4m7MquPx6g5PPHpoBy/DA3Uuviya6jcUPaVRn5U6xr2b
RQr1dM7Gq9eVsNKELspjhe3HnNmziBrwNFErKx8JF0YrbA9BK7YtcD/DGSRgDyi2
OXnLkgw0jE5d5WEzKH7YIhPA2VQKIEIk+YKmhA7pDuL2iNSe8WdE26b1H+Bp6JzJ
K6t4dpuIrMRRnPNioOuncsE3jszEKyROP0nSTjdlhw8hkQCuCSaTVnGvvK1kkgzq
P5y/kT/yWpug5VNCw+2sJzFX9tJXBghJQSUvcD/7f7+Y/jDLAcWqdqKNbRInhPDl
eYHXhMUl1NHcZiG7C+192PeJLJVBKRBQ4mRDsYHB3qBLV9KdwYsOAl2JtAHw2c1P
9R+wwgjA5vTlDcGYtFVGbcpVP6daIlZOto9zDRWAVK56dumtG81gqrnv4NZarUyT
zVzymbBWGDftpvHHyogZNu0eErHkKyC9EXd+gk5lfELMl7PFvorfX/SYI20dCWFv
1cXLH3UUqSbPHZta33iG27cA27dGP1RnwwmcptTYe0cGRCqN1gfmqxSLbIGYHrXk
E83RiqhW4SiLkVDcoNAvtk9GGpejwWcPbE/Aj4ms9dl1qmnak3UOS7uYDZqIP0QK
0mEw9PUea1/isJSEKkIIoFyccUyuShBJN3zRmRMuJNqL6LN5KNETPcCIcW365lWS
cOPTVlP7/GTrNyfDEDUKVrFjsgL7eQIRxMjxUs9BH8rZfP9z6ASEvEIUvbuUkRz9
AetFHogFZeIzW1YZqVLG/Uc7ruquG3rnGwSvN/nYmVxhZkQLl4N1bf4uYeh6ni7Z
K0YvdQE8PGYVzg1jYHQL7h3ZGABWCPHuzedSG21QjaQCFXdOGpPcYMPlb32CaTAB
gBWImCmX689YhnUZBS99Z2ecY18SIXMT7CtFb5QuTaGL5Blnbju6TI3vj0qTRvoN
TNzFVCnIcAg5+NcJWQvGGpYTGQ8DNKJYq+yRu0x63xwDdzqRwA7cuwLIz6d4/jl4
utGvfgYWMNridn9hQPiFeNZ+1bBQ4UCOZ2lonN/BUzqt4du+p2GWvS33CSvMXNO/
ntroyLCTvpmTuVfZ60JXTXGoaImIERdWS1+aU9lecrXistPeL6hP9Iudylex4PrQ
DWyX+6xUXEd8IfrHn+54H/Yi6V8N0zZ4YpayOcD/uqdcztGWmSSnFPes9tQcT9mY
Lc0NVevDoZ9E48UeDLX+P4DR2lIgbCLF2dengP1vgG1B4TwSRml0+JAZQcSvaHQz
dVeQCHWN/pSkgnoMoHis5dLBB4pju1RNIziN08Z5peddFpWiNQZME1b78My3AFQ5
v/swHyUR0TZqEKw2wGNwph3oyJ7x5Ph24s87fxyLGT2zJHDilHofAtc/KlBs+gOC
r2Q1ReAdynNYV8rAgvK7RG2o6ceUNAsquDDX4hS4Uzn7vKNd+haM2pr9AGGTZ6Sk
5/OMWF3uH+0pDiysuN/PPRlI6bUFiktGZMM0mFsRo01a7ohbHGg3eI4mjOoELPwl
GizLjccNjK9xicyw6Ch6pSfeLCIPtbLPxRtbUbD86fpHvCNKRMqBQo/U3NFUS5sD
cmEyQIevkmQFbO8FOND4/ijpFlQKGxKaknF/dt4priMYq99hlf/QQ20lbVJohtkU
vFD4yx6h0LQZOsLm/lrjKXlNJe3kU4X/Zj0kPckoFElKmxpkmNKOtr70ARpZwW8z
VvU9oxhOjVpu5IBkebjYaG2hZMdsuI5OMUxhBZl6gwD4BQufiSfLnuCERjahXdIC
yEFZ9hlUt/eOIsTI0w5CP91ffZtzjrVslkODWBuFr3n4b18xWPPwHsVxrgzXAyI/
qec5n1ZdLjXE8tvoFRxlAD0pvqIC0bsSxzv1FgD1C/nmT9EHvZYhLxaN7omrIjeL
CDGykbH3gYaZBP1buc5UiZKlA5FxewcAVxXAPU5qtll9xb+Bbl0Lev5i7isXTuUH
KGGbRM1e9LT8qBtKSJCDx0QyTgY1LAad0uScxrTgPm/RGVYTEX4LbBzs1U/+qULe
erx9pJ0J8kYPfJfXHeQOTE9ePHCNaYPeu0LVMRnC3OOA1ETaCyZCVJ20FDYwSPL3
HGpdcqyLPBxlW6h6ER/TLHfeqL9Ff9M/OqjVfZTzaM9Kzl3xZa8oreIaFp2g9AYj
LP5a094yHHiArxRWYVSbMU8YS8XexDmmE3w2Ble/xJejlwt32iaqoId4cydJq+Mg
GVk0OTKv5mDBR0vOGiB7zAfcEIgzJnqE0bWnvyeOw5e7SejO15xU6wsY8pNVoSEi
7nAQjchfumJG7gPSFOqNtY4GMX5VAP4uvsuH55K0kzRNwsIPFydEcyjw/qGbFO1t
056Xn8lAyDAbDb3IAGyLKSx+5AFyyLNAMC9e/2HhPEPUoECDi6LgfMYBAWni9jFp
aolL/Vtx6xP6nKav18K1GQ9uGNNaYVbF81maTo+tm1nJidQluxfZbZNHJfBpUauB
wD0HOl6Qpcuo9DaIngZUj/y7lwASc6KGGBZUuGTxeuEB41Z0fuO5ZsUF95mg1Jfj
XhfMnP/wUUh/8uKe++GrKrvSHT4LChnmibeiWAE1P4+HxN2IVFo3QmFiSQrjQ9lN
yPku6grMgfRp3k/EvKwc7fSoVctwvt1VpyWy5BKnXoUHbMwztFb5Atoy0l2hZV4Y
8RMp0Gaq3fCYQM64e+Y89KWc/BYvvb5jfkimV9/0EPrIf2C5fdKmsHejmvPXGuqT
Bq9AiHm/adWSx/zzoCjBJVOdr3mTGHXrXlBTspi9cujSXjVgtVSJ07b+UQ98sQey
faQZnPN6Nw8BEiT5aIfszEUfg6Sj0ekxl3X3kr44vlJrmN0kNdn5cFaUdXKls/EP
cHByS4iiONhhvqkH2AKgIjk64ViY67gaUjObi96EFI4LUjm3qaesvSU+bvKyCBEe
cFRA7waEtvgbqlQ8UhZnl+cyyzbAAC44Q4IBdv5HNcAIuNWI4A7css5ghU+yynbB
9dZtgwmAZGffIp5A9O8S9O2y/2OJ2YMfliWBPmRDdIz8/GaHVpp6zGThpiKGB/9x
ABEsZ0dguKXlFQRa+rUqHpvd70HRQyXgm/bVOveKgTyGXZLPyVIqNq9c/DqgKVWw
iSbxt5vRPBGG8b71CPwk4pLCZyh/svDDz8PChxvaXvCkhIBT8b7QFrmRPCeRDcEL
M7xI2ODTBdXwi6nnuoDPsrlavrXhs24hJmHZv+c2MCOpyyYlPDiBygno933edAJ0
/u8dE7m8tG9Ziz+AQqHaau1zUMgP7D3yJiIljOmYr5j1dR71fwQ+2qHP3mfWrQKs
BcokeGS/Xyo6y3uIF/6qwurLGK50RvbwCP2eUP7II1xyz2YuKEeHiyrFfDKcB251
Dv7Vc5kM/mh3W1GQf1ZItK12BWkXCTRatzcYf7kh3aVCqx6vUH2Ivv1U1gXbatF2
Efl48XWfonQ89CM56CYws2EcOmOw0H7aAwoUR/dOT4DeElmMtnZz6ped4vQHLN4u
fbC0kSZuuGuVm0R5QG7Zhof0mONFx//GBQDWiN8+ffOeLXHByTvXxBKVofYxioLz
Jh+IcPqtt97AYXbE4ds4AFFwOtc3FTU7V9vz5zabQW+j87Q+NrnbBpHo0wIkdbWQ
NFDSRtoEK9zUBjz+wnYrpGs5vJK6zFwkcihLajHvu7vZ+wUSmwSMpm3/uPxZQ03i
GlFvFfLIAf45BYHWO2mpFT8kSXKryIN8FEod2Uy6Fl0uVf6p9RXR7Vc63h+pD8Rc
XEJhzcTixIkWcPjF25XprUwKndNmPdakWJ7xmYky+auvOoACpu28qFWSYNlpgIfJ
YY8CbIui5zpQhPcdPRhN/D6SmcQDZLnQZ+4wbXHUUpXhrnDJZrWXuuvAVkQdiuhy
JDMfo48mRVyeQELoqF/Xpz861dV3WwYCuE9pWXFOJI3aqm48dhEKw/wwNlTUrJhZ
0eg/MCiNk1+AyXGZD2pLUlCy9anCs7CbyZ109xv1Tk5Xsm+OAC4cP6sUMqN4X/Z4
kI1Az6B60vZD41dZWZzllWa6qEqje7Txen/WC4L515BIlxQdpSW2L4rz/u+52Chn
zy53B8YndHslht1cLacQVEP9ugTPt8s02hXusFL03In+R1+iC0ooJCGez7pR9DP7
ughCPcfUewLFRJlOMr5DKvcu5faPgOu5PM1gqDlHqIluxsNQF4OpTCg+bZGV317i
9GqnumYxgITkL4/2KzZSzqxaenXEZGNEieJNeueQC33YSQ+pJuGe3gSi90i775el
On0Sv7KdSj9jyQvmwobDMWr0G3tzC5z5bTR63I9HFLZZBqmyIewqGpbaEIErlu0w
TPzdonOcBkUU0+o5LSh58bv2DDcLK7sLj0rCShrtTzfEbvhcOi081yCmTilGtCIE
+l+FvBzQFAXiZqeOhI+gxN4gvJX3DsjmU80pC7Yc0ICOem14aIo7h42e3SrpIh47
+JJlVdxkP6V49DyzXedd5nQu2iisrBDgqb6cHLUlPGYiy6QrUtbc/YjZVFlfEu8j
YiY414+ZNIQfCFZ8iKDo/3YTVVT/g2ZzyKJPkC1QaJyjVXTf5oqA5S6DUJ0nXKFb
XltFBEGw73LdZzbZCNKDmRn9jEPaEjHLZAFw75NUiURqMqpkOChprJqJk/ql4GSP
wMPIVNQ2OfZbt+yD1+s4j9W3QNBJd9KaiGcxNhGAtk7kCTbMNnAIbMSMx2kVLWhp
eRM3whJgArz0mVct1rma8VSTLCioD7K6+LLI3GYh1y8JHLTBG3v76jpZ4YdTAsj8
W9tP8DRMwZXNTRXoye3fc3NTWUG8mUobSsMPi75yDBNpDHpWsTd9+CP3sM8kIzuS
ycDl2ZzSJ6UZxKL2MC7w3JM2rFeF/u/gVolTxccjUXLMnBioYmQhQQ7Y/KdlcVAS
SyVutT62QOopTDeuaSh8k8juttQ3x2Nn4v6/VL3xBV+tOGTuf9+Fggp6kHyWwBSM
sV4Llz0FlsPqmi/Z4ZNuZQwnTpeKGWYmJ8DRteYAOzW2PJ+pZeUqQ7gKXG6hwULz
CRvP+u8gj9BsYFFKwMAGYPnMMoSkUpUkTQe7a/aLNY69xmscKPfKtlS8uk3T8GZN
dNEevpN/psCmEbQrEPQogUc+1URyjEcSF1rX0+Sb4Xkokr6cXRmYQ0L6sG64jvBt
DufoLU9/s679OPv4OJUD8YMut02blu1JpEN4nsA/dj6OPIfrD9Kl6bA5jaopfP2b
EL2R/nQ2ZfLal8gZfUyFmsw+KRn5bb5Up6byZTJhBT/Zsl+CFr392pAG6QNmbhgc
rafuALJVy4KiWHkI2BEj/+PT7EbXC9TAOiimO0iPMNSY/kUPRWtK7mcoreTpC3oL
/iezoKrYIwVNgMfkXhkcFuE5KC676xv4CJHNQTYWOmw9N7iGDoOzyH0Uk6/wJ0Jl
+aY7GPj52BtG32Yx/YvZBB2UOy/pCv0AwmLxSuULZyP9QHLCqOyRW/lb9zPawwm9
PIXSDg3ywgJ3KQxbg56wTgcz6IyvDgH5cuYePyRmKAXuO8l3hUePI4LSmVOQ95HV
L1AbE5HEwRigQJB0eWCR06jRg3cTkYWFSfDxOVOPbgoZMHy0XDIyky78y1WqHQ7K
XlmCCbuZlIr1hylmwvYrtplXXWL+PDGJj6O0h3Z12Skrrg5sTCQFNgBmymJs1zDA
Cn1N3cNIwr4dX0NwX46DiUGeb4pdelU+aTPn5NnwF27WIQfaPJrP+6n1X4ioudGQ
28lYr1L0HJWILJC9AdClWLsph7m2Y4YGxpiZFq7Am9JPAt/G9K+znVus/gd7t7aX
hHkvj6PJYEnIY6f3QOiUl7MvHcUE03texkyx0nwCrgSs5dgyrPnUmUBdKOq/CApa
UOEfx4gidhbP51wYF9Z32cx45YmL7sb6tSj7wnJN5lj85hlCh4zi1Mjws+0q+zTI
8Nd0KMzuxZ3iLCH/pyTxpT9oFOcznSOIhUg1dOBw+4xHjh7Fv8DM0KciFOn8fzv2
gmT9PRaHsg0mg0P9j6Bb+/5uu5/dmROQJmV+RSV5CF7bsEiUvwI0ogBurjLx+b8f
t+r3G8fJoFsGJaz+v9yFD6yKsNMs1SANWKrZrwK4If2CteMaP372Sx9WppDLrPU5
16EJni7yhUjn+9viGt41aQIdZaJbGwYFlPFwEP73+XO0LxuD25zSND7jFHRNZgJD
CZ2Laq8lhJbVQJGGAdsCa8yw8oMeVCaGKjSCjRB4Pn9lJ6T9xwM+W6Wtuq/CIU7J
iD/VSy9YI2m4Db5Yvym65gPWoExhkx/KK72SlwafX/Ad1+dF5QEuegcrEd+wKzRH
DcweQjPcp0beeKojVknUK3XUWScGsS28soB9HzWz8gLpjvcbii4Bxyfdf7kG8Jj9
otkebBqUL1wpIWXbP7n1DniBALS6jRXx+Exvz6w+JiPUfn1zmz1g2+RKLICBmoKt
R0z1lP3uxKdTKRYADxZ7dZ7iTIO4tgw8SizvVzRLh+X4ZIwV/NIb69UiIZbuMqMk
glyGm0D9VxdWV3sCF6nQLmK9gO6f35Mqkslsd/zKEwzqBAHBFmHrjLWG5fAYWyMy
RU07BgqT0QQgRmiSfMPqcL0FGiOgsZ58RtCK6PcjTVUOYkAJcatHUQ0UrrI1y6nv
oe73qPWyVIH2/nGjbSlUBayI1h1LUPaCKVG45pJ01MEKsy1QF+MBn9RCr1iYDxGZ
kWntv9yq1fPQD/S6z1Ap7AAf5X4CfTXSHA+P4rLGvV5zdL1JPlPBydjh7A7u4SXI
auNgJnbKjQahhSxEDcKk3SyfoY9Kj9dksK1YVUF/Ws8PySbWemNaF5Isrj+8IELd
ddT8GRkp3QD+W3kIiTCxlDysGC9N9dN8Dj/0Ksbe6SWoVpJl+HRsiIG9lcF9xHu4
c8J/mTda1I4W3fSWVIVHEF2d2yG4wU6USWZ1Cd4qE+oEGVSa/q7U+F98oYwxcf9C
pMbRcBQUtsBDFBynCJB62GDPN3c5ts9Ga2RtlePbP9BPO/Ov3gwoBRWRPWwZzMxD
Xl9wKCciTYboV2qC9zmN71eIcyUCxijJ3kOu42JO+6mjCWD8pLPZ0YDwlrM0X2pE
1qR4rf5yfmmms6iTh2+LT+nKWT6AAIubbXiVLcwu5k5sRtPYhhXGsMNrRxHPPWAZ
Ob8W3S+7wyNeJQV6WitZFDv2JkWaqVCGveKxvIGiP1HfeyTuXSqAfYDig7vG5mKn
IUgtYyItKJctnqdhpGO+imMl0SmzHH1Q7xxJuLBDJk90sUzfSQrwHNbFACLLl15Q
JWbMmFl2QcfCA2b6zfoTu5VBznNK4L20D5qCNNDpQGM9+b+Jipv2xv0DdnxBTfND
zUq2pcYv624fMBFsxjGwWEh0jEbcpJEzdCI6084B/Xhfx/IeS7ZYjjnYhUVM21Ya
jmS5WYD3PAlEroY6/3o5M6sDgUe7QoRjiH5uZk7iFk1dV9b3Yv6Ve2TkE0TYQ8tL
2Pr4mxDYWliGx25IyYAWEjgxBiVKCr5ul1+HxRAcIbxtBVzaCaldJUUMWlPWtH6I
GTmXZODjSOlBPqHm+IBEyvTXJMWCGeytKx+Kq1FM+khEnu86JrSoDFfmV2vjzoKR
eviw9YTaFYSfT2ikxMf6MPX9BUcJcsVP4sw7UVZY5fA/B02CT97O5YrtXpk7h0YM
sHdEDS1fVcdYNltHQaMbdv+paWF6+ZlSGMRD62q9R1cRKPydNBWl6idqqaDiNes5
hpsYYOSK0Tgxr4/BCqxJNRmZZJrZL19kZIuxNXltiSZNBAsPpwCIpTQk4sh0JHaG
9WOTnJ5dIIC0u73YkkE/5olDReR9qZsBSXYzt5TQTEJXQWR96WCZtLTEI1YTm/aB
jUzTuTZn6vH9G9qL0hm8/bfPf+K4yh20rxuc6CZxTzglr41e05CQfofYNHuMLupn
k3WAJ7DNEHfvzK/STaLC2c9GQRD0M775dRDocxlRuMML+5CSsgCsglHmg2SvwtT1
xcIp1ddnvMmVAEEIlvd9UCl5zNRGhAXv0m6H+GERbHtnrGn2fdizNz4HaZBuD3iA
7E2uDaUe437Fu6CpHOQ2aZPqrzJ4FkH4UVgNrzAyRM78fxOQn7YoahdCJFt7zin7
h1DjszuZgGlENMZdWB3NrV9BbB1lMJLhg4VVuY4zFiNcEf/S3DSY6QaMOfBOk194
8IPnWSanmJW+7hOABDYKT28Uky5b5ON80uCea0jWnlHbKaezMvxZ5bY/JlTKmYor
J2c+t/ol7UF2iG5ih7cLwFHEYPRuxyiqZziCa5jOm1OrDJe4krkoWsEO32e3j5m+
S5nUvKHG6dO+Z/8CSWrB7TgbhUpkNET5ZDJRCt8OA0e/ZADjBA0IMVuKgMlSl0GP
xIhNfagUPBBtfQF109DNSaMaseW0LPqPbuFpUDY8P0b2bnwacEwle7jGUtcTHX7P
fd0Aa0aOxJ7BrmUjM/SKUysnYwYuLTlW0ATxbMlJWZSS1oe9cvETogR8wfSCU3xL
o6ecSPk9/Uwb8ufKQTgUQfN2ZzGmHBnP29OXsAFIs4U2/kSPZ5rg9TkQj2BEpv2L
TByhOfi7u5mqKm2+YiYly6ahrRgmY4A/5e5TmfAIXTBifFXbgdhM/wVTEWxj3Pcj
bOCVXi1NWxWZauKOyoUZzZE2thhw2eVYa+J7cc84nhSUdob44aGQgOGiMdIcXL3I
EpEKOiRkJsUYyEyqaXIF3VXq0sDYrjzfkW70ulcEQ2Kp/gd1scawaOI6vHGuCTTz
lHzLmh32gNME0mgx5EdF3Q97L9iPJvP0f3tA8xWa2QXBVE9wFDORr2mo87OV9rKm
i5ZnMj43uE129N17VsEoseCEYw0nKWuIdsldiopoP4ET9gwyNoSPrzog0uipVERj
FPOf5HuarzlGpL9qkZKD/VHs4QYd2xb1tBpHXrf6OFtJ/7cQPg0CCFNHC2Kkwj4W
VQk+0TeJeETHjlr+ZrJeos0ojkfu+KExshbUS3qnQYrhYFAKfxfJ8+MiXTH8ECpK
b87zHpGtWZt1ZL4R100scgljVWOHOYP+Xs4r+PFvGsKcExPCNEeykA4LmdA1vXy8
AsTxicWfkgGvjHt/oJ6qUWZevoys5Nf1KIjBfdzk7dNYDgkzaVE9qfCXL1I1uPXZ
kGHq8BS8kxtmytEGywhStiyUhNeanu21YI+miM9YQHubnGF+OW4MlJhE8JQMsWJc
d4IHbt19hdIcXj/VED60wDZNLgArAUG0aBJQCP6zFy2k4KFKPodkMqdsZzFFGy9l
b64MTKKUoOzYZElyXhyq1utLB0GHrt/v+q19zHbPOQMOJybgGBPjrqg7cUp5EwN0
Tq4jO9YVCNxcwXmmGTSj9S5hFfsaZ7malBH7YkTSaFXWo1uJ6Gpj4F7YoLkB6fqT
RQJztchcyRBo9XT60LrVErMeMA9kga03XJoQJRoJAOme+dLe6TwUKxGWMhZYO0fg
CCTEn3jaj8eiFhZQ3qh/gtE34hgLd62l3p9ApRWqmy7ktfHi4yOM1U1NtP10Ivnx
strMFPJLgbdXrnATqc1m8JRQaVoBttko5TMcniZPPMc5NgQOfW+gpJS+F45CB4lG
iI48joGb5i8nvfbksYTTFbpPRXzhVUGtK4wd3Wj1qZhXRWOZBmZPyCWrC7YmdI63
mx7CxRkD07A5OwuRxCz8eGnyjtNYHoTqjxkJ28gYtnAj64CSrpr12xdzDDLOx8hU
5Q0HdqluBXzC+M45fA+lDRQ+R/Wfo4PwZvUy3qR1e6I/rfaCimOed6M/RMHBP0cb
EQH1nwEti6ZHZKJez594G5XC6bAoXaTLJZqbYDckNV228ouo6166QhacYGvdNEOG
7Y0taJZZHKjixIDpaHkLigwG5og8j7F+5NjaJmWxaCgRiU/ZwjzSsPcaaMqg3Rb1
ZVVl1qZrLPedDcLXoSNuMhAZeie8XtC+qGpRk21LDrXj5EmKz3Tve9c17HJbBZ55
z+hiURQvUUyGgbYgxicv7T7r7+S2DYc/gPpEhcH/9j508Nj5IdvPOuc/k2UCywSW
OFrzIm5nAKtt1NhI2eU5Q3Qlfv4+8KiMitGr8Hz9GMNmQN5NeI2IGbB8YoMevssj
sD0cUNRTo4ZZvugP8r1t/ISNsrs/Gf2WWCkZ6/kCc8+V5voJf/MnythMrlkbKHpd
KqSCk7UMef5LbYo00p+tC7UhtHnE8Feeew2icn714bkvXoTTq+45t3FNzKNSabAG
IMMgO1kPM2/bdG2FLXG4hLybp6d3IFJ//8GYEfd0caLe3pidR2Xn+enMwBwlpFnP
kN5qkIEq2d+2aHj7gBH7JauBqR7DEJoYR+twPofYa9YeVJLhZAJRV+sGPJ+/mdUv
922BvXGE41+JZ24rphbPMRYNGYce2SJAZB3+O+Lq4B6oCyyJ7xR2wb2CYrrLAKxE
AH6uqbCU/+K0SYN8AyYVLl4tCupwe98gIttk6wfTzCz7eA84p1lqa5FXdGBlHJjD
+aSZyQbyCdh0tjB/SIpvd3MMeIiFyBrnRq7bzn8rUn0cAWAnMi+rZ0xZe2xmeLsf
OTvdk+PQUATDqMFuh0mv/n7kJ0WOAuDI4JPEoZKC6x2YpESXYMih5u8Cj1nCp01U
ufiHtGIxe+LwAr2HXzsKYDt78+MNK9ZcIgWICGvfY22NnnM8OxtUC9j048/LPGV3
3sVpMB14O1t0+vY/y8JKPYE/Ojmj2xphyuqiAb+JLubMhS95uwr0aa8JQXYswjZM
ZJea5XC+8Xc7+XpEnMhugdxMDp9NdaMgLNwoB0iT9j20D9No12KJshNz8wimI+XL
wOMIenX8Ir8ESkYnAOqVkHYgIeVTy4346xBw91pLmS6z6FeCAZZsb//n7O0sE9Sq
JyTeLnFVkANx6oRuXUhZ+ZiWYaCms5r63R2ZpmTd1yUwer3+TkLzeqcaeUnIIUK5
hV9Fr1Vfy7JhQVWm52N07cHFJAzbbrnLnEL7JFXwKNzJjAkSY2ujWlhFmqZTPJ98
9XF46h4NdM1beJJnXN7pC14dwyiUGOXiW3QCdeJTX8Ex/K8Spd8DbHKzt8MZD3pG
FW4NhiWL+Cxj5JbXZ/pEJDYfKdZi75FA6cc45k0VOpLhyVNjWmvbVTKTvqjKUkUI
uhHTvKyqDkQzVT0Z/4HxR5wnZRUo2xeoxYDNpBUlBxAwLmw+gtuHD823AB/7NCHh
i3EvAG7J0fsEM3MyoWsWeASzsx3A7VrXf8WthcEf6fLzA6paf+51RrLzJDNASfpW
itbFnV3yE8CdiBmp+yxWoAofB2Vkt5kZ7uH23RHptCGnSSKauLDcg03pSh9XkkGV
Tjq9qjJtwl+yc6MRHUNvnXaFXfUBfHTkN2eryvPgp8tbcGlR1ynya73+9xl/3kmc
0QlXCG3PUTRIEer6NXF6kjEIkvR/VkmEB88L+N6ghhOfudQteLueAQmq5bPV8ONA
b790pBnTi8yx1U50/GHj6dpy7Oloe7fjmzUnqJgS037fmFnvs5a92HfWbN13U2Sw
uh/iTEUaeznTRZ095+fDCrDMpW4nc5GdMdCe0J49q2R3Ntb3sre/P3yRKhyPsL5T
fN0KeZX3n8L4ThLbt+3D+HM4C3p34IA9FSjYTCIl2GXXzeO8dlN0QSac91j56WLX
5k02f7Z884oRXZ/Ad/goBDG6N3vHUoVQOrlOdHUvUcW10f1UHDbosvLPPwJYbZ6v
5YCinfVOtfAL4humyJcI1noNzFGAd5pdHXyuTPeM+IV4BDG8e930JvzlG6RPgt8y

//pragma protect end_data_block
//pragma protect digest_block
vLAsnrxUKbDjXe6b1F3x9KbrLBU=
//pragma protect end_digest_block
//pragma protect end_protected
