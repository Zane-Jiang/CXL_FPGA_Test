// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
QCDlrkj/JB++hZb7BJewZuJPSp1bXD5GLRHl17kFE3VdoglLs4s2eAodmlWOMMcd
AmXSJzSsNP0+Wrt9cR3Pcwqwb98pAzsuXeVrcRSL0I3Ac1k2bf7LytN4+VreL6BI
mqEYF9iUCPrjUma725yYeZJxjXDFLBWd9UjwhmhTyTXFtCmL7qoy7g==
//pragma protect end_key_block
//pragma protect digest_block
RRfdROgR3OBwekqkXDOpjcBFwaM=
//pragma protect end_digest_block
//pragma protect data_block
Xn53M916347aHTz6+BesutQRZNeTfOYwNE48zr41QA21zJQf7LapSSjI0yilSKZq
/31ckEGJ9wIJWLgPb8LxpWyC/Z9pZ+rHgseXow/4uA/7ne2e/btouCVVC0smUUWI
o95LZsbe9+YVlZRdE9ewr2fG2G2YNzwweZ0D7ekIL9GYgv6eGEmLIE7lPE5gjHun
m9msTe8pzRCEZdKUWm9xoR2tgvC2eupqOFhFT1T9AynKTU8LTpVFgmAje0/IEV4v
HrzJH5fKttIYrhredLj2oWuqryOXLc/plqDE17dc1e18mCdu1bqMfw+vrzMPBB96
eBL3fMdE6m3eYz80Nt/4jvGWPgz56u5C6UjVHXLTrxDa/H87Zfo6eAaoWK4sHSz8
gnUrrbHnIqJrXctSz/dVJLknu3i5btP9TY+YEl0liFJ7XprWNMIebK+Z9PKk3e9r
/e4gJnSJ+Y2zaql187O7XAxQnjWYri1TBRZifZmWDAx2GYcMa09Xu0+JpPnz6KpZ
waYGtQS3dYH+jn+ZI1ruhNdq114PKFb8kwMtjqmmuVWIlfQv4FE5tPr1qSvonAwU
tuAjBpDCTboEOEKNt9K2zn+XI3X/dBxtXQHcVIaZf5KVMkYs2UGJGNkLCdwbnjUh
ReW+0e0beYXYCTBkBK50upJ4xtpZZyNsh8FeElKkLXuuge68+GYJq1snUPg//zyO
zylOC5zi9WncravRgIa+T4FbX14xzZBGgLQ4sJkWZpxxpJxnYQ1I20oJXsBouh/E
3u8MpN4yC0n7wq/WZiMKGhhYSFWTR9VvWVvvxCziENvg5lNn5k4YnyEs6HGfV052
xyqzTujLpJjmbp6ng5Z+2TWvllemzhsQ7pOoF1cwp+BhNtBE6/j04Kxq4mzp0PTx
qsHD9/n3UOVX/fJ//o22lL4DOkMxGsgKpOZiYbA17heUZ9AT7A1IMGrKvN3KCZNq
jF5fyyPSFFlhxmLIiJFLgIuQlJPOa0h17EmZanDi8856q433kW0XX2suvEVKOwmc
uHI/DVdA6Re6k5l6UaVAlZhI9wo57YDddBPU0Q2cP/IxHhzOwleJzoVolQ+XxoW3
4iCKGX7mXcZRFTtdiRzT7Nn4l4PdawwXYoJpprOAVj0Zx4gy+K87M1MXCDMzFLqN
acSCdUoIt7B/VIgnzqYCaZuCBVXwZkjlkNQ5uvoU0cudkGpAXu7zVhw6/DcK0zgW
8u1r1iM/bcejnT9pYAVVwRf+sTDf9qiOLnacU1D3gVyouRjV71WiORTw/jSOxUNU
U6YO8PuykRwYfcNtCYRRF91QPQ4fCkFuj394vqbnDVbwpSBwcJy6myou3okng+iM
zA9MM560VmaIp/C5TIoXK1sCN2cVu3brYzfJi8SH02CfZ3FNmInCCE30gduinYO4
UNTlm1F0HEd/FRfiKubhGjJ7vf9O1NfNUtUceEMO4TEI4eHgIAJrm4/jUCz/cAoR
i++0mzGoW27rl3uXMGoe3qEwYpTNylSFsvYyV7rRCW9cv+4hKHrtVVJso0Eqmqua
KfETEDnPE6Ryuk/bVaTq5MKQeY9jVOzLSsXir72Fg8NKrrJz37WpilOW7D2UyU+S
i/Csbc21LaSWOTKwC4wFh21ns5OVpfJXGK9vFCj5fCC5bDRtrCfAqXgsd6AvdpF4
wenUf2G6U88d+fXpjhdBvMMgOmKYl/nGLEUI+btFnjLxixrNoK6VbwLkqiL4NB7W
1BzCSxUmKgDGTgXxg7ut/eFbAw0J3UkYb7cg98O5rMH44XQJm3JSnoeQ6a32+wfZ
47Avaah3/2Ki+TerMerJEcpIQK8OQZTMYAUTJsYghAWwEB6NH/rtDwjD6PjxgCrP
wJobvb0TaTgdzLSFe5NKX4bDpIWybpEvQh2L6zc0AoAvNgwlTGhOYxcS2uwagHUS
iG3LOPeZHG72pT+4k+qw6oqpary8YMRFiULnuXqV4ga71jkcrdENNhcLX02498vz
0BgRR9bGoSmFcDCN5/44UeWaWxGxu/ECwqaVTXQdkjnL4VBTgKqv7jslxCF0h+QZ
crp/+h+29YJ5ZdawwK/rVzZeYbk+0XtSbg/PD8YZZDRTW8UoWDdE/1WmnrNTwyRJ
HkNsCriz68SUykqDpr/ysKvPhq/wfu20lzZCmRH9JYUpwSijQY6j3WpodPl7B7hD
hVHsPzQKl9F+2k7kw0abhVL38aKa+58XuM75HQ/0UGj2wHKl0avI6CYxGal6xMPH
dctecNYW9cgJis9ClXYmL18W4/IEWKCNwXzTVFQ+SygkV/+h/Z8rZI8gDK3EM3Lg
P6SwuOq14br3I3itXaSv0wT0YQnP10DGkkChi4PKMMm7ctS0zepz+8xPDqh7xahE
eSTvzOgkPApGVmSguLmYi5cVyvbP7bJ9ajrOcSZoaVc5mToRxTgizMS2NYc5ak/V
zHwU8KnMdTR28porxK0VDuTC6+iZ6GOi6KFlgPy2bF/OPnI30phZqL1CqX9JYEaE
pPJIji+NPMlnZyvwAZwqgRBlxr21TXd7l3ngpPYOtLKqKuc6r2snfbk+Rx2AQKsv
GUvpQZMY8L1NxOIT2po88Z1Q9tKSm0dx5Pa5V5/vF7v4UVob9AixooQUqRFoXZgm
mr9v9XQIAwlqMvBLO6jNilxBgIs68pBbsCaRuU0IqEeKLXyKcrC6PhGqfj8/5Ysf
V8ZKxNyeEA9BxZVRbZq0J4QBWQnDvHSIV6/ShbZCHtJ71/gbb7kj7FaqWBm6MxRS
VnDdkdKtpZ54yTjYcDgTLSO0/wyMiMYmK0lBNGrRM90czlyPv1+FJBV+FsDBna/L
IKIZEJRbd9XF+RJ7kCbAawmg1x3aoske0INZZSbd5Z2pqPsLWW9focfSCZ2YqWkV
rxeT6CR3IDb8BOK2fxfnWgXuuRWesPmgDOow6txlV3Pcnj9oKU2LSX+cMFARLhMG
WP940yNAmpp4MYdl4EB8gNILxjTCUzSSDOA3ilyI29+STqCdH7nODYsc8+fpPMwI
3jczOjL+3zp7YtKEX4zF9TCWwe1W2A1nfyzkHEqysUhva1fs168ztNgbwXQMWvne
yn3ixV8amMsb6lkEyFF7+egO7r+yjyEz/g/8d0gxkndxk6VuIS8mja2n9h9GExdP
6RI5wIp5TyMQCSw2mzZ7xG1jCDFb0cEbq9wr3AmGKe25pXzJd21cvIuq914tB5zg
+QyXL1RjfPvu4A3VlgODdTiPnTWoCGA0cjE73bSQHjdsxNhrIKyhs+gXmD278lC4
mJeEeEuX5QlFQtqZmM7dXlmxjhsahdzxcXvH0/fQC9/79/+9xf7uQDchx3DUm+9R
+hbz0xmBO3FkgPKpdPSwmNWdI4TNImhGZ+jd5LNyFRI6lHGbNZUXbVBRS12BbaU+
63xtLsuQ4yj8abz+zbVxvHIBL7wciBKH97MUFR21Idcm3wFMEQniSjbwoPfBx0jB
3PzzPfVZ+r1kV0PHkuJYiewU4mgwz0BbF7zoBCjF05/emwcprvmuAImYPD6sZyQb
AN/8CRE64zk56tXwjPTf7Znv13kqI+nxz5JmwkwfuMhuXlWyJPEDcO9lgv2VwBxQ
496gS2kbKtZUfevIMJA+Lj1eUfsrnJsSfz10G8BqNtsZ1dQR5TeLX44hCN8AtW/m
A0aU8G/aca89bcoHbNGXADrOldkR+IZMRI4akq5AMrcHnGMwUT0pD7JKBBOJvi5r
Z1ytOmfT8+yFNdnK0alYbz53DEwLn1tkWIaYz6AK4eJ44+tJZkiXpMLTyYrt8Lwe
RY0UWn9j1qrUxzXo5sHv/gFepvE2uC/AtMVon1qoKh07wUjfGFMKbNUhBZ8QkCs0
JN6wagfCpB3LEDdLoIwFAbmTpN7kS7U+4wCDOOBdEhBwnAs6uwxP0W8r4O5twQ1u
/WJkPrR/X9CZFcfpDJ1/DRRiLFU2UG1omZUqsb9SK8d3AWO6gCT7UR55JaGvOctH
XSBT8ZAFd+EWk6lc/6WbDxjNbdesV6yuPqRk7v/ctcR2+QCndOsnPNxTkcCbDqsY
KCO2DjN0BItX9i3LE5Pg+yVn4FiazFkVzMaxRFhHLhqHZJDtDnLy5CChJbGNdsiF
9R+pi1ACCgKtVZMJpU6ic4KYXACQllDWTSnIzq5ulu8YJwiB2DQI/yjpxjh4EdcE
q/R95315ubWPWSE7uMjEkQDoN+A5TdI9bPtsND6vCeR0Hc36ScI402B9M5dqsGFA
BmsnsLqJrwakL60fPyXBeRKejlMiYlQY7b7/FozYaGvpDN/UBhIuY1pyaUqjE5np
Hqty1DkRS40382TEdIMmMHFaHBr3SfJ/TK4Qo4lpv0UkgtcBcar0wo4eKxdpjJBw
5cNTq5ghlMSSKVx6ZSoZEZA9g4YgjSJ48cF/ufVfozN9oCsRgaESFQyRtVUXoMg4
Tt7z1dq8GL0yAuUfYBhY5NPM6Q4q5LPnbhCuF8tHr2NgSJybuLxtTHVmzfS8WRdt
QU4nnu1y6K5LPvIhqv3lMQ56Lm7bJw+NgyOCpjMY7CrMosnsHjs1lzKhZ8xLyKdK
84DiNShDTruvEMzS7wnRVeMLF3Sj78iyaDMxrcQKEPQBrgWMFPqN0bAYHug8p7BM
EgnkaicQtpZr+wx5RyXwrSrxO2RtaiT4ER5ISqyk4EMhxeMq5R+f5dSyFNjobtMq
2uAQac5FFNIHRatzimdEvk+oVPy855R2Vmrbe31eJ2JuWXisEKdSzoZffCmMEfJ1
wzZK0msBtJ/aNWWl7qTqBiqBPtSbPDBlXVueJ9Sf8a3EBiaPw209KTbUxhl2LMqk
dD4Fj8vVVRz3/ot8lCb6+BrY1kkitq3eoMltq8BEmJyZ3q5j5HPeeXi4OlKYwmwt
sVBvUz49l7JBK1x60YfZt8/mAwAwELeOsn/Rxnx+EUN9ZtXhLvo6VTMI4q0a9xN8
SbxJs8S7Az7CrbGhNPqErobsdY3WSiJmTrz27nxPIk2X+P3zJfrwDdBZXeqQ/xRK
4YnBsQ2rBPjJPWUQVCmf/F2sYbCziCCn4Pb/1pVTX2Q+YqJwov8d0fL2dBjoxc4k
bkyUAr0mEYlq6hGv9KQYcphXKCmgQwx54399L4OjoyzeKaL8EEbGWBgdVSmJd/wL
zMFbLESEoENgHN/LQVW7qPlQ0Cou0tfHzXje6pfrGVCzZ3ua86ro7NAuonrdoHk3
5t3tg+qqNHA2aycMotcP7H5EeV57LeqwWRVy+HWWGbl+mecsO2gEIfLmcuXoHt6f
WFDnsI2oE06F9n2AWmNqvqmFhKGsl/z9zaULLp0sCqF6LjzavIAXC8g/LTGVcRAb
mlOeH4CinUzrHUA/C4EcIQvll04tvYubwCi9r8/1z/izRNHqQdfnMVc10FBvrgVk
0LOVgsOfqlyNjVYptG6yhnbIU4uG47peNjGKTABE9rXPfZEvhjP6I5gYA6rpZ5b3
ZFGsSO5HWawS6uqrssckzdXrth8UzWvjY71eclYUaufXU8K2INKViuARJ29AM/Mv
VZwTt3ondFL4kMy+Pi/aQ9f0/dzlFPgy2ZcwDwKPrHxDtFYaVO4tk1v/xJjBUqD/
fof/s1r72L7ZGwD1zdvBqv5rJJauaavOz96T07RzK23SHM+iPCu7CtUHIOcKm69U
B5GyC2S7JyIpX/yLWFPlo2ySC20ORhpKPGm8IbpmS/2+8++QO2N47QNo9YIIxFSU
+ajpbmovcHI8oULiSNTxb14hch6+1rU54lkR9sWMdhYIWCymdyR9jHzoeQ8l50fV
RMZ+VgKLdLH5ntwvOGxzIR8CMOumMVN+KdjLcgePMNLR8xTMz+f/GX6MqdWPNZ8U
UvXcYJdN588PHZPoS6Kdy2AluqAHzOfrbQdvSSRwQXz9Zt2Fgruty/LoIHjKNUTx
Zq5MKoXZjXOz9Pf6KDOQtOXmsCvI5TXzobICXoqAU+vNBjYo9tUa/cMTVWlfi8gm
hAX5s8Czi91lIA/mWifu/U7jZpW0MJ6bD0sSIVxvyRGqB6bdpbnu0NtxiHFVjC2O
ay8ksYXS8t7P13PjreJl+jqgJc48GfPhPiO0PPSZyfIoOGhVWyFNacRsjUwWfwqS
qyYQY+L7utl+T3DOprz8KqmBqrT3E2zZiIkj5768Lx75FKlGuxqkk/NW1JAPfRYZ
H4IsmNehPFJyTJebEnUVXLkHsgqerHiHVI6/uWQRTBo0MTwYeoKVlgfhdI1uEr4E
8Q/zgJGlAXO2QOsshgdS2pvr+56VP5prl8bbhmPAMKTVxZOs9Mwn3sLQh2OZBcyz
OiCzBlOrJGuBLyubgnjUR3JSkqsC5snqaYY7GmCo2c6thFXEVSr1spvhBAUEzQOl
pyvCF+u7CP0A6Os0TVASX8+ZUQawnjij/jYq8Gxp4Brvxb6K9Zo2EcKUSB33HuZ4
O3G0BMpr9v1J/ysJ/HMLl9mW/i2Wctxp7wc5D8Adx+XngF4t9RajzXUXulx7tvhD
VaU/o6Enl549yPh4SRm/DGlLsXTnBUBJDFRDBy6JtfAfHHGF3aRgS+svElgCt2Qv
k8MHYHubLRXl6MPFEBpuZZqcIlVWzfXZhIlkgKqUDim95fWavaMVUdkY2ZbtxohC
f39nTH/STW4VFKtptZXS+6WPaVfo/7yTIWGplGwRIvL4U0dUZfQCVENk1i+kkEFT
jqHD1v3r+A0liE+nOdM4X8OOwTvMZAfPEvd1p15yUA6jSjQfgrKAKbt+8qZ84ke0
ZdEy+80LLkytwTIXcHMqV6nGQbey214SjLYjSCusfw5txwFH2bxu0//kam4XubDo
8PdhkCPB6qwDrPKOfgSzjctevhOVhk9g1KyQwsUrj8bsty68OMxT1Ojb5mVr4+MD
9oLkRn4s+PzFMi6CRCNCAvnxORWG+KWKhQYgNAjET4u0rNmx+zg2mMcvTO8e1Yeh
P1/lJDzWB3zIfVh812Ioq0RKXG3P6Qi9Up46Yx4McWdYh897tSVDY5Z3rhkl/KlI
FWkKFJc44KVKtS5BC7uJUW6yZm1GmysaaUnSd1Gdw0saDkj4/sY66WmRpxRf2H2s
g4UzxwOnI7I3iRnL3dSx+E33DK8Cbs/rfMqUxoOxriHmP3K8SZhPaALrXczk2bsO
39F/x+XPsWS4RcCDGRNUfeQbd1mou28chLy33VxbBRfXX9mCtFCJt+ao66XP49az
BmGKG1MeidCDG3htwfxj+JQBuzbMmUZDvq6hMAYi4IOEy3yaQRatl68Icgcw3kxS
kSHBmdKz2zrUnvvwnLtDtW/KTkVgyro3YdBrwA9aYN0MkJSP/NOO0qxddN9AWYiA
09/RZhYR7yHg6tlA1SpgYER/JCGNlaX/ABLLV/05JzNAJkdBKcXybDFZDJaob2M2
QpevlptyqJb2iTsvwjMxies/uW76D28vOPPU/8nWY4jVVi+TaLcEWWbZ0Ruj1TKd
WCIaPqS7vF5s+ncEYIDgsLccN9wMpYWe/QkUw4EVG2m7UBPmAJSkErE+Vo9RGWFe
LNvA2vYEq4zYgB4qx2VBy13kaYhMKk4AoSwLxvo1uG5wbgRyZWlJupyrTb3iqr8P
oESyfsmysu3/BPL5OcjRgFchXN+TMI21ONpVKdkropBdG3a2wPe29WAlyiwS3gmF
jg9g1F27CwesmIb/6TeJxvfYnb9YYA9FT3UsOKE5QPAivh/GjvyOtiyRCtL6AwVv
u31eLqPPKzl3DVxeUygp2cEL3yaGJDhkWbUOcAal6KWPj/fFAb5STokZUkWkXCRu
ygwHgnWkv5RvOnqmIYq6Pn5u5JFZzqi79nQGU4R/2nCtFZtUJL5xo0SH8deG8G31
hRA8u2XZG91BOdxKZs1wNNUBLy+Cgp3QxACTF62hvSvTQE6LIgEQW94xrNTmAqOx
TVqidJ2jRFDPsY3JdEMzGxDuA3+5npTbRLkBCv/FDVzUEwuj3cAHejMDLR+S/K5A
19XAOU0KTghuigjKjwqWsETDSLs1DkrPTKUgAK+u9ZYx/6Tw05l9CJN/gKhcNym9
jjvxmw1x+cgWt+kIELYIoIJbrSUJdmW01+pSM7IfKiFMEUy9SLx2LJCIufPRCcZP
lIAxu/spBfuAZhri65d6WP0sC5zqghpJtqZcykxod1OlrRIwPscCeyr2wHQa7gjV
XYcwowiGlXziLlHW5iVHzuArWZNZhBYNSZFkBo+4CbXdhCz9+CLtmd+/NIKMR8xp
JjPNJN3ZxB8H87qPVyYOynhTowP3h5QLfYSOVN5v+bZnnQpUhMH9IGMECSPvzSh8
rjH5kAj9+YqHhJWXwt2F6mBHShF4iq43mD1J1QcBqck57s/XwyOG53Bitoz2pW+g
Lr5cpw3KNt37OnH+VwRCI8IN1AI3roIpjsqbjNYZpqvcQL9fiomiJmFkoDwmFdSW
LMuoYs7bBQXPg8Vv+Y5Pn8/FOEo4c55drmANJ2Pf6NfHTQhTR/CoaNPVh7gT0q/6
HJTGiRXzz8g1baXI/osoNuAwZiNpuhCcyDQS5clVLZZqiKZ3LX/aKOyN8i7lOpvR
5KkF40hdfhQcFFrBmIWcXHXn/O+e05Geu/fZk5zWbhzghu/squzsiSAirOtgz8Lv
o4w5XoPfS2E1Wck25d9kqczzp4CgAuGZ8+bomsR4yyKc8ta5dQxJx9wPzytlgDuR
eimpILprrXS1dJcd8f0znqY+u4nCQN5t0Tk0JcnVZ4ERL/MAiGCOxJD7vTSrzrwx
z6tO35bQm0TnVyT22LIakgmZZ22TFpvej44FPHuDaEISfDVqethJlfX1yf6SOQ4a
19lCdfjNKe4Q2vuLj8FEnzdp/RksaDFK+ENngxuOWxlPDM8/JcOWgeOlcmCNltux
Ey05gsQzbVOpu2pPIOk9itSUqXY3LWYWZ6/Zukt7dniLgl+KHp1XWBYuykyw3GOg
JF72oCeRWBbvaFYmAIZ34Lp51E2UmstFaqY8ryTTTx9zrog2F0cS7dQBkf1gjgP3
9t9YdzHNZtQViy1cQfhjfKk/f8EbfWZCfgfGsV4TaxG+5mbl+yW4E2HAiMaU+NUE
acdBI4Jxanz8L4wCxdOVxudIaaXVSyat2uuItiXywlhQJi7wnKvjViVgU4m+PBWC
fYXuMizkbnIu8FCxMt4kcR05fA3b6J0/codnj3hysDXnSZ/oKcZkRadsiLTY33H0
djeANZpGrft1R2HQIlVyBHGuCqqHi/NaUAaCuDixf+G+R1qMNUvbhph4No8s9Tkz
OOf7OMul7Ap1+1htlJKX0Rzf7Ibn355gGwWjZJG+KYzDiQ/2Ign7BL5nDS1pfEKS
v5VpiIs3CaGJJUSR4XZNDdFJH0zukjS+hR1XVHkFPXS/vCfUP2xZzeZ3R35c5Sbr
M2LZ+kHnrp3711cbzgpHFvWHUbpjDrpqMsMGiZDUPY3D8pdi7JUSRSEiFEyKnAB/
m223Tt8R2EpyND66nHfO5zHxfjBZ7o0yBUw6Lp1IRL/yld3Pmc5suUC8gyeqVF6Q
vYpXvenGXE+QfHJpJ2rMTnNSd0dIeiOQb3bU8oSEnTLsIEluAiQJBnBjjv2Kyz/I
Nbf4m4/ipufjJRWOsJZFg7WwqQAGLZF5WDMQFRPDQBDFl6sfSvN8aGxTM9XxITbL
/vXnzwQ/Vnt0l3dGqjDOH5EE8Z8wy56ro5p8ZTVs4yA3SN5REBuX73cj2TKQsIPr
5dyDVqiVSq4Y4gZzNVqpGtlTk8bAr0avalrBb6Gy3xpgSWyQpsx9v0glyrhrIQZ9
aGJ+dWi+QoShME7AkNxofV2tgQ/JC19gXkS+4zTxjJDbZzBL3fDnaTSF+F7KVBiq
KjyaewVmSOrcSU1yelztBtbJLFb+bFof111RhdYwteExlv6ZQioA93BLcRZ51NRt
ui5KctS8cI9Jkly1y7yXhzlJHHJ06Haw874lFOiNSU/ocnCmdcHXPSG+wGozb+NT
ZnaRW/0hMGn6PS8VLdM4tLHDcpBMEFQwN/WfzAye8rPFbAjz/UW9RAl2t38p4K0x
Q59MfecwLHmTyF+MRamzCv2NkWK5B84oAagSakq+HaVU5L36amTxPLmZffrUZQop
lCZHCU71SMh8p6SLhVT+hk2W3/gywQqBov2DVlbVkY2MnHMZYJKgSVVkfEJxAqy+
K/h2n0VlTGcxaNVZO5Ch247Rwo4Xjp/Vt/VTwKZMXHfYSdULRNIdIyUNP9V6UuRH
gN9jPpUpZRF5ym8UNzt5S9stT6NwY9MbJT6f9bjnv78rj0DVqh2Rz/wL3dy+aITt
bDLY4uDZUYp+E2w0qHkKPzZo2VDQo1TnRkDnIjefpSbBcFH7FYDpEzawhV0QUb5r
iOuVX2DpecLNZggM25/ZcFKYLB3B7+DtuanNuHvdvcFPrSaSfr2J+dzC4cu2uiTs
7g1RfxyB+7AJ44hdYcUJRRvdK9WBQ5dAgfasgSWrlVdYqkwFvTMhQynOn6eXzPew
YA3pu9bFcIs7VIz2dFfwsYlGNnjyZw2pJ+Q/Hg5jsjR6PGq7vVbs7jGDJkF2P0Ja
+1y/iAA5sKHISBGY73VkQyPlcobO9QVexXihzpQqfECKmiYlFnzNtWXFXRPBfubv
FPzFq746iVvS/Rwy9vJfv2tyTp2Bnij3+/yUB+ULQshWFafwSIcu7lMKVD24fsDI
meeZn8x4Adt5WFVyY6HKQti9NgFi001z2dHIb2UPDZS+h8RlhIddpTc8eRUIQQW6
HAsJxV9AA3tv+WQqcI6aB7y/RHQVbS9QBvFOgRKC+LN/HBEV81taSQnYBy46Vrst
AtlpGZMlOwHPll7en7yqcn/7WthCr7fWU9e1sXDDQ12LgOWIV4X1C6qRfSRnuwhn
QNIdV/AnRumtDh4OTUeDrA3JSUOSSBPhWcdJSOxvBQaMLTMUmicy/x7sE0u4qg9N
JcUAyu+axvAm/wmZ4emRQuLtlzdJ5ecHIBWwglqW3gOwXndyq5JXhD160npgOx4V
netrgH2wXiKR8J1/bHzM/WJ0NSemQIB4VXFWbJybol/XRs6JVtizG8ok1gEyzq21
p2AgK7Xf88E89DnFbzkk1HxHqoiDOTXP1SkkKfDZH4f61idjyE/CKX1z9Y8RztwV
3OT8tE4GbslUmvZOpMgJK2e3ewiIVdWL810VfaUKdQH9uwvfz8DAYPkCivGrOY7A
xhM9VKpQGpY3ho4tA5+vVJhp4cs2P7jC12C14LC5Dy1+IcJAv7tzxO9Lw6TxGcvq
YwVVlp4IT+72QA8F2aV3ky4FMKfSO8+qMWOl3zmm65UPPXEPm3BcSRpMh3coa3M7
IEhYBVmUVm+9UTWjHst8QBBTL7gBQjEtMuS07z7H4oTo4HRJP3EWNLOpLu7+XqQO
RpsBXeQi5/ZlhLBpRG26Rj+fQlkK64QnjEhvs9RF9B9qcEOhvHqvPx23DvD6hYA9
JvkETuNM0aEhHbTvUh2lLrdHIKT1mkK7XUc7EofTIeUf3GR6yWXR06qxBrMqTE3I
qcgy9JEzo0GjDwUh5DErurma22a/rIJUkAuF8fzBondZkHvg+0N2ZSRuQLbK9YWQ
Z8njoqVLYdBVxKf5q9Y4gmUaEL/dCDbq5jkxK4l2q6ttu6QuURbvE9SJJxTpc9in
5SmkmKcklVSPQ89jWryofieNFgZwtJ7Nda4CthtbMpAK0q+9/1SCsg88HtYy/af1
rNbojGP0dcE+c8rY5SsnKgqHVWBAZmBfb9WTWzT0zrE0GZBkrlCaLMIILNEEgg9x
H9ZK1ACkoQ/M4Kj/v+MG5vVT1rZIvJC51PD1sv9h/sHTNy9j65pOYCH4kEH8SEjU
a9QTxh8nDUvlCygxpiJf6ediUf/OCpBTzragQQRGXLdDvqSBS/EPeEpUdC6kEp++
dfs5Ig3D5JdEf7Egjydbhhz5LtUy4aZqM4K+hCqqc/VH2dMAmuVk1WelmmPH9H1T
hPblY+kJbmfk6d7BKJ2+GcPHDvYqynqPdwXSqlU7WmHbz9g25rE8r63Oi7gezR+E
e985uYHLDb2/hpvCIJnI5kNEephf5cmJagt9ireHzi0/jtoGzomrYevrgUeyNZC9
tOdv0RHSBLdrMSC9SbLELDqWTkVLidM05HAiXf+JLr1rjawnEzm47iFG8HeiV3pA
+ulrhemaOUgNoh+hGHY+g845IVbF90Ep+pfwMMBpSDuzD+aIUDww916KCXz8xubv
C+tVUGeVccVOiRCLoHd5O368+WPE6FoIjKitCyP+2weiboRALkIAb3A/8OkONuAN
FO6/JnfM7JEJPWYMAvGncoRcoxGPgzusQaFtNl/rC6bwlvolPIaksGZ9DWBNRNGM
cKa03eejVg/mhB2BoWAaYwIqO9o6b3+Nf0k3XyYEcDqrgQM3H37XS7T7X+Jkdp8h
dZxrUSEDfXNv7zgC17BbIHpbo888dUp4zjfE0tTkgqts/hN/DpUTRR3Zf0TpgfnM
JSYbKUYtDJMYBO/gyZbzs18U6tNvu1VZaBohVeJaANh4/8Wm3rX3Yy/7bQkr4zlZ
XJM0ImCAJb0XxyWLfy2Vh3/KKj78XtXrFEzYsZCNsBpTuRr8QmuBbv8tyeT9pA2O
OhHqMs3sj1gwoCCPJyeI4YK/uZxRHcZwwWgSTypuRNWVlNVnvh/8vKe+SR5wdCGM
D7jlr504TJ4xTJXkVO9gcoucN67JBkg2VHapU2Sgum4SDqgVoEXCKoN+iwH+5BDX
YbVq+uyhRJvwb8mufPwfAAMowjHIoncPMkaJ2/+qz1PE23AZTr4X6ee/BUlrsWux
OZ/YdK2TNPNB9zLKtCFB8gNZUsCGNv1QuOue8b797Rm7Mu1YS1yUlDfC7qi17H14
j235exgyII7T0mqqIH4ZZ63WuyMuIYDBRPCvyua1aM8paQh7jEEsZ9WSPzXK5esZ
jxc0H0TGMWP4hk0fHz/nDMKin+UuddoO5TkrGCAPloeY7l+OboQrj/48wIveGk+a
4ACS1nLSfwiHuRjs3N+3y0p0adL69VAYnZxOxd2NPJIqObWLiMGeolLrmRbuEYXP
U4C4RYCxwop9j/opy4KLaPpxgBmNvJ7C/YLijfrIqOLtqN/n+40wKOx8uD8b6HSy
D/YnU1tIngG0zJjm58RdoDJNi5B7XSOT4yZhVUCP0bE5SoFg3gbo2xAtdBeE6cZa
JJrzYiOARR91ZRL+U1L1SPMqGd9/AyiAmWz9iHVi9Oa6VCdiImjdJ/RfhxEEfAqX
5LLTsapa4T8SvQr5IphrhZWSu4i3sUYVrTSvhQeOOvQSs8e4u6rgxto1+NcUkmNP
tlLQ8JkSIy5lUcjQJ5bWB8cXBzG70hNOLLc2W6jPIeae62iOUYY52HiN2aLmcDIb
G7U/WopGFJY1pQmoFAUyJyYGU3dQbKqgtmuBYH3PLgLVPL+axmVwNfdWxvd1e7eq
u9tPeGesQbQqP/ukpG+imG0Al9UFIcZmmObS/PoICKCz4b5Hr4hcC42JEIOFvBYE
iGc/CkYioTRfgJnLkvqXNEIx654bqBKPRo61O2hddrtqlD9FUxgyyhLUuRwnqk5Z
7k2xeQ87KeB8Arl6Gi/WA1ApDnsCSW8ZE9VKzNGc6m9ujkYrkwAwrAVyrTIIHd51
BD3emQSUv7IA0AzSebYqAJnlEgWuP93PVGpn+7lC8vxw6nNwZ1CZhROIMy3GWYOi
/ZO73q0YCZ2MJss+rxBoQ7Og2WNviQe980FBrP1DHtX0N9HYeyR66fPop2GH0N5f
UTWDBN+ng2mm2bSlEx3mLeQ29FO2pviZnQoaKHjB1Ui1TsKj6WIXw7PJfqL3WwC6
zzhueFSoHTyCSyk0iBiSEUkDiGF4IUMzbjmEACKuMbXJcNhVj8Fqhk6Z1QsNf5wE
8yujK8EvfJGSCkev03gpI1Zu9/w6nucrH5xqRO+dcouJAdvempZTWzyyQnC+HsvH
+8nBykj81MZb+nqwOXYNps/bcbrNQOy3kXxf5iRrgv9fXxeLEcUA7uQL0CSVGsiM
aPwarzRdZnPXfvUI+L4JY7ohlLJpp5aVwpJVdmJbQt1XAgcODLhTVjm/zkbklHFU
lv+optrfDE8fFJlAYb0e8MkI8x3qnpTh/KOS/40m2D9POnCH52YuuKXB4wosoqdc
LI0Nhv5sGlr6dSg4XQm4/S2H66dXiCaXXkKYPYgChmZIFp0eAUPPxn70Kj0aKPE7
xeAC9kOI73guKjLLEKeRk7wm32SEbMVzKJ7dCpVt7bNSX2b+5pjFhgYkJ1BIaoHb
Bd1H2TJZ2Sk/MS2HVh/gJ+rrBGuEoG9ubVNPejKexj+CoQ43Ll2m/qtiDzsxCTrL
lhnXGs0DtHJ06fLur1y5tPApmtgE1jn3+u65KRaKmzrYH9P7b3UbKX8/LsFceMMk
7qboCqpI9ABfSDjV+wJdp0uyNnDzemoxn3Ftg8fl8iiEis96z4yIVLXIPU6x3pYl
oImMu2uof8Jt5GAu4DrS/FywKe55NVDUgto6KRtAuGUWqRTbw0lkUseL89rL673X
NbBg19L0fPBIqlDV2+W0YycvXMp0D/jA5g0O8GPH0gQGwQAXXhCyopvPIuCPQIPz
VS3Z3fAzJ05h9ymx4AzC6E/y3Xvcjd3nv7Ub3921TWjdoXeBQA8hm/XKSxVxwwlo
auYv1cCULu76pFuHThMHPWsNI/FTXjqu0tpJyhIWLGJQhink8CTigM7ac7FbElNS
fvU7zf/KL/WEwqd0DiLaHOh4f3KEv0sInaK0QqmUwPeB5XHg1jAKofbTH0W1mR42
VrERUbmTul++EoRj3riEiueGM3HC5doFm0Q5vK6D27r490yXxKb3LxXOZmADhPx2
offX4FNkV9oTP40az5BIjXf/KzDjuUYr1X04/UYmMxgnKZZvxugu4tgMSYpBS99R
FsORAmjLy2bThUf3pg2zjZWjY5Al4PpoOPPDyLvWPENQ7cwwRwYiVTqeXrx6ovK3
gWrTgiv9VdAfLg2Rm9DnAUZjvBJbcBuitfZ/mRHEuo0y9AhWamq5l+jS6tQvVDS5
r6qM1Z2oiXK5DNFx+X9ZDxGTmLUxnG91ShJ0gxqYT2znHrrMoF4ELcX42C+QiMYR
DYI1klefcomOPr35c63nFZaNv5m7s/vQE52wJ1dVGCIZLqVBXMMPP/I3EJpYpZOK
5nYOieWh86qWy8g3YSMgs+QKj/MsI1detvtBGn4/O6UvH3fDVOYvggvFxm+xLxMz
oRcst+YFE5J8/otKOZlJRaF5VcVIoudB5PDvcgGPqkX777XHmLjce8WX4/pGVzId
sISxcx8po64Rz/kBsgAm4yCGi4BIkw/uJTKQGKVOGvyDf5/odR/L+YXj76FGci4X
bAlKmsXhouqdFUpFi+9sRTlEiqzpmaSOmna+r9rN2I84LzCL77QanARVUTthrS6m
HCrVf45PWhX9mqAyJM/Bq+F02lGFeSc8mZmc3S3wwyqm15PmfrMpSMM7KfCSwZZI
bIL+jn6fqdfgwnOWm7ybG4WPIBoosx5OG6pZ/2lrLL7CTUHd3EmvogTYDz8DgEUh
kkadjIZHRIxM6suhvfdiJ5YKSOJowFzHLXHVVJ2S6WKvgskACksMAVrAcAP4EaHu
RVL9LKjH+oWo+/T/FgNaJF/73syORKb70Rxh0+uJz31pyLnFqFbUmg80SavvXjgi
vz1+6y05pWJlg6809MP1hG2n1CNLiJKZg+j/XAL/ZzYGjrDXVc/TJFtKeSs3mzDx
B/GRl8zg+S+cZPtxxQD37AOi6wGEY0NEreQkjMNNaHvriLjghoyUoNmWei9tDlHq
anyskrmA34/EjQqA5ROVP2ZJr/gIxUWMx2athetaYcEJrCJSeM06XweKhcs0Af+v
5aUGjwr3CmhSOzM1Cl7ppbshxgyPWSwPtk//blFDVUSQc2QB3KoOo9g4TmJp/tS0
upJDSF2SV0T1MmsNK85OvTjHhdCNjwCXUuxYUVp9iMBZYjryz0G+jo1/4mMdCBgO
Lb/Ukgu5N8E7iUEXDkR1hvRs9Z5KVbJNRpTLlBXXqtsv3OEovTlIR2JA/ZkbcGHV
FNPtspT0ImEtlwyO/niECgS0Adg496XJfSVZYk3rL6WCtmi1YbZpTdwDrsN1Z9Z6
2fGl3ukDUxXzBnd4cQTztpoFZwEU3YaxF1wK4ipvB8n8taWzxgVC3rhKK0kVY8hj
cJnbuZZc5Af4r0LmocCwj9n6xd/kYemRxKNY2xqJKH05SmBpLAJmYhVmQIfX3UY1
5pDnCOJiSBTaiRGv6B+hmI7PXD4CqBtBow2Ge0m49rP+QlPW9aAwZtPAcXxirDHx
eDW3e8dk2nyOmuAe7upencRPUYiYAaY3nZBpaIUyM5GDJv4U2xjcxoCnji7GkV3f
1omhGKIQyfbtSNGx67LKqACiVgwIavLk5/PiXtowaYlpfZ+sbt7Rx7Ex2JOIpDyN
jFcjTwt3zp8Y/CBIjiRNIkfNSshQ5GHqdd80NQ8nbXUyp8ZG7hS2E83PxS+FAbGS
iIGj/Myht+rBVB2GrBd5vkBpZIXxQmVg2/jyNu0Ti4Ok7hDmohjl5P6RWoplX6t3
VxSoqBimS9OocsPTJkH2M5daEgNmDvK82gJ5yLysrFau2ErAZLfworHTe+njXbbE
paXi2PssHPEWry0A7fVOZV9nHgzmt97Rz2bJmBc6C3zCgf5eTuxkhrlNZzmwYD+g
xfJaESAL6GJxBr/tFZ3VQx7NELQDz91w4xSS+7SDoKScTuJG4OiTNvFsHxKEJsz4
BeXLLg7NqmlYi6aFzAYFt5K3Nq0bqLXdkNZJLHhe7UhTtuYxHjxzcO5owqtaXsgg
VrJMNjHcjJFIZUaSCiUz35Gtc3nK4R4AzU+WCcCogl+1DQD+iRlLLXR/Bk5soF7N
NzFuS1tAMxszeAWKMTwHKBIG7yDZWOLQQR/4k68BUgrPsyyYxORvGb2BYaT9mFMH
MI3NphrFhKNsxALj6Eqa0NmyWmxZBZDmijzY/AkgC4NGQC66TFH27Jx0AJbn5jnR
7HCH2h7lSLimeaG2act0ZymgZ9qa7josoymuVfTkmRy7rmZIRTRoiUnQk0alOz/M
i27fjdeinVBOYUPLBnHkHI8TSffhuDDpSiukJRqzIE4iJ5VS75T85x5nkDW2O9rF
xqLxUDBohkz9iy3aTWXM29N8xKYkPbvjidUx6LdoxHmXsfeIWW0L292d7VhP4EGg
ki23lefghYbzbToGaD4BHquy+Hv0s7xfxY6SUgHM28GG5vr9Rvjb4GIbToyaPtx2
W9hhp4FYKFLX17ksBI0gWRyhdOZ4Ar3INc/V/P3SkqIKKIepyfUh9PdfHF+z/Wkw
HVSXRY+pL5RV9+hRD0VCFxCwUP9c91g9WGh8qqlsMukYKxTkRtrw54vSsOYEb7VS
kBMw61RLrh0TjVgcN/gxN4Y14w3wBEnv+2P55EKDz54Belrk6Y7lkO2BJgy9dpM6
ydCw0IDVr8SA5oBamvIPV6UJeNYjLCfKWt4ssAlVe7RCrUPz11iZrUB8qAvLDvh0
oQxC1kT++SQ3AB6MLBbdBFbG7ZU0yGWihXpnVGpZrXTliHrEu5pjhKUKorm8h5tz
021Ss9kxgfdK1N8ED2MtcED0UIHojcr7D0DUCtjedGm3hSkceb5YCcHVayT+NgKi
HhfiDXQOH2BQugGscXcRFKWCpTotot5n/i9oQ1QPgKs=
//pragma protect end_data_block
//pragma protect digest_block
uaQEHeFxFHz/oYAxpLsQKAzQA1U=
//pragma protect end_digest_block
//pragma protect end_protected
