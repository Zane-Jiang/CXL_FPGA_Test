// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
QHRucSGLx6zijxEuDkSqqa4Ra7wtFCPqTcJBqAQZsf1NtcrLQAwDmAUnJxnOZRe7
unNUga5qIYSU0N9UDp7GYPdZLyCmZSizUVaZ2it3aEBMD6gUhOp/4fMAIH1NzFun
7WWAGAUA4KPFXoi0+x3UKM87adKe4lf7J4Y56RKG8hJwKtsjJs+DRw==
//pragma protect end_key_block
//pragma protect digest_block
W5mwW2BdLiyVZoXLw/POVaa0ooQ=
//pragma protect end_digest_block
//pragma protect data_block
pKtUaBRgEJtg8DcNNeLYgOKk3juWxRl/CWBQQM8TZTIaBFem1Ip/qH5vtxeY272u
QBjMbckw0j1sUf+5zlgxq639hi8ZpTnw8eOCyjCtSpPkUZNnEfmv/IuHPIwHBe7S
OLN/6bBLUfSpOxOhDnlda0dF4KTQ7uOzvf4IMyZuxzYGF9/QP4esUYnXanqUL5c9
404baABxuJkfM9KVmK3IkD9XPFZsQLJqmJGWG3lJqnXLPnep+YXgSoP4RP71NbJ/
tn2Ejuqoz0QgHtXd7F9eU8xfBv+raCLySL9j/BYQoXF0bmE60SGxA8ZcoN4+BSKo
iszQgfmAXbS1acFtNtkn7DcEBEaqHOA1IkP5cSOhLgh6Dn9OzjbzoCRwsW71vF52
CNMXxUOHxHl7KWa3DJOdhDoMM7K+BmLqdh3LiWagqitw6fAUMd7Hx6yaI0BqzIG1
7IniMhZ1ByLVA/oAJPg5b62nkiESkPcqHkAvWPXVLKuZyC2f4faUPUhe3018JkWF
TQwfp0+f8UnNNF9Tob4aLNGXQdQ534oo+qjvNMwL0MA/KBx7zrAVOwKa3rt37gh0
VWRDZpOIYuUen9Ec4hZpXMKWhA6bC3M6+P4p/I5f5nwaSN0zO5bpUwBn2VQN6jfL
gUK91sMm/ZOJhPhEmXGJyVn43+ry+kA/SYrsYGoD+u85yuBp17wCOEyDt7kIRgtN
5WeUsU/GBCeuy18RQlg6Q4FlXCyuzgf0Var3reijukxeFYogHv0Mu9oRcKocm74Y
GMiIwbkZf7togNXBCRhYR7Ki/CT7LOJCXvOKf6Fuz/fdvBvBp7FS155STC7aSBrM
2Ia9F9hA/qVaYD3fJNHwqsAG5T4l0j+jZT9ghNLQWmjXVhXYbozJsPENbOPtbBG6
M/cIbRgLcuwaJYCDdaa4aWLPsPDFEiBsY0NEClCeKeblJA8Ek8ylgKnQ8tR4xNRP
YPo8sp36+lenuxD8sBt1ZdxBDDQAMmvM0ciubrR9N39frhoQBAeuMw0LGpP7gr3Q
0PvnddThv+UWCAZKKlzlL6zsoDhY+EmPH37vANyPgqrU4ypuUbpx5OHqrqi5eQaF
Mzk9CE69kK1wDX4y/vSTHZJd2OavYf+kdkQFNr4XkUnX9C4VKlj+3qJAwMn9HQZT
D9fEa6RHSuTsEjcMTNQMJP9TQtmxk/JXYvHApzf6Meb/Bq9aL/h/H4x0g7x/8OwR
hVFzk/uxdiM4ohbcvpzz0UtBNIwOnHCrmFqLiK+KxIaTIWgU8DIdIcMCamJnoxm5
kYb5BLrVNMywycGjMOepp1pE3aLJrEPNv7gllFFGB7r+8mtY7PppV2uank9mxSid
ZHU+Ii6OfOooGBjxxJT7XG0kk6MHMMtaTdMxI/CHvPHj9E0T3jkKSg38UprnWLJq
gPGPAKGmtEojaSNdAGFzjOGHv0IQAr8l5lVa7wfKBGJWWPvk52JGGXhVMaiCmtI9
v7iSD7WOahicf4VKZogCJvkhZuaoLGZxLUJ5+hcj6LHvgl66074D9LOP3kj6SYQI
ShPBOJRtDmS3Nr5btwHrxrIw0BhylWJu5KunR4SVzjiVfaeuRPEKOJEzdZSyYzGy
xvxbD/7dDJssQDiT3uRjJ1h+tkKhWQ6mLCyWl0UpBbrXnYuhMKXtBcA8tYYEQCZA
mwjDXdt2Q3wbC9RsIyZwmqcOYFqRJSsPscbbvnfaXbhWCXhqVgLx4yOSSZBHYMOK
x/2eELTDfb6qQtMS1E2wQfCy7tPch3SvL+LtjpQKkfzhI/wcr9mQ/K4wUfBEzVuh
qjLniOYF8xcxdUB52hy+T4/Ov/EWs7jSBZDHiXHLp9eCZGt25MAWVPRL5nJKD73K
xnBzlIMLCbzGh42aLWhhzuUifyfqYr6nGojOTxJc7hTJEd/eJ1R67ZL/kJ5GSKv1
UTn2zbuuVvZ1lQnB+ZQBUdi2DkN+MAvIWWHxc1Qg+gzHQ85SEPF/1IOcIWoN6O03
nydqgIGkfPlpOmHd0w92MDXUC+p3NfV3M9SKRG6OoIuxPNXSQYPBRdHbsi86Y2f0
sDw78KWIkfmPY95qJ/Qu6OS+HW/QlqTyzJdiwcyBv7RyhoYndap86821By0wJbck
owFBIcTuBPXSR0nLYNWk2CCwX1sgblGu9SE+5+eBLXs5vHKsd3hDbqGHcsUzppWp
1rIyWDTR0ZwuZbY3slfDkPYDVntucF4UdtIvm3wggEfSUxPwBdeymZzaSZTlwMce
YiJVPeYG064Cljy7k1o49f6fEd7ooOPaFd17wNufkmomlC9FllQOu57IkhU4LH98
EpUQ4E97ZjCMC6H09//wc4hLMZDCz14xcTmCp1dmy7KxvdqFl8Ufz9i3ZwnELJwJ
/KUhPvXus0A0iHm8kAb6TXSZ5sxl+zHRgDsBywS1weA92lPkeqSzCT2aKs8uoRy0
WTdtQTL28l6ViJxiELivRm3s3jcy2Yv17fKpOHdrAyDNNel7FZjuPUJqqCPcUoh+
kGlh+3nx6lgNMM+QE5QGu2X70YlYh7rYs4K0o/7md1Tf0/yUg1/fPrOpXm0TZ44+
ESbuDJNTBIRVGWNhTODBHKO0iwmysf0Ncnw10v3+M8E5mXmySWUeDTl0ZpGyGXju
YhsVnYqxv/YGXCTXNQUn+VZrTbZ9mb581VmxzW3V6XWOBstcos2tHoNwwiijs0Me
F6ZkzIEfqUVialMLXqCOOxeNK+ayZ3ZXpgh4auGT4RHfjOdNVTqZUoxOEj56Rpgm
uppkbcAE0LTtHkmkpoIooDc8slN5m9ScSuYotDxOpd6w6P535V2uuVO05kRC2JAd
a+AY9XabS/ZilfCaNk5L/uCrm6cpkhxuYX4si3zzKIPt5RCQ/6QDI5P2JtRGwoTi
kSP5upRHHRnOdxslYKzPy4viQrl5FW5twKOrNxtK5KhCpyGKJgWZmuFQ/sccPirB
S1T2HH58UMx5e10Dqlf021e7wpyaRAXIf6w73n2WQ751Ks3S7X+1AYG5j+h0PesG
WIkIvzrd6b4DJdAtPCK9CbyiUt8sVHGpnbnA9I6pno6fwUTQPflqdVCoXBZdFYkM
d3XlOsxhv+KM52B2RD0VBPSgGDVVM2eQtjhk+eTPvmft/dEpeiHexoBoC6EXh5cO
DtiqHsCo8exP4LlMrOEFV5W0oDR/1Uu/YVLRDtmJeOTMfUUTUiAboTCQ72Y/vsH/
68plLUn3m1/UXbyI00uAo4NVk7Hz1bIzZ0PPI2WPTyenXPORMBgB5EKw2XFPK8q8
brIO2WalEUf36US/3fqrvs6FeqHUYGq0v4nmING0LM0IPdVbSBgBRvzyq9SozU9P
74WbvML5Rli482Ro55b7i1G0V7QvrMC+EQ0o5B+GPdoAYqf+nBna3ycZj8ndovU0
FUbVXhqZJxvjb6bmzFXYh9INSKsuzotpvRcQaoMQqP2Ks+6dLwPhXGWYHnrJRvp+
pRt7N9r9HjXqRj6Dx49tPcqd9vWfy8f+e656fax9Nin2b8oEN03SaIyjVigxukGL
JGvxRzHnRaAddW7ZOXuLpaYV6sFCFp2QfNrEEMf4QYeal6MP/9YRl6GsuGcuVQIn
ouRfJCd/hDLO8IiV9BP5rULJHMNsRoHeADn5q6dnGLFQDlBzoNsSulNCOwaYM8pb
B4oUgkhd4gtWEG5bby7CHrYwX1mHGKFjrWTlz6igPglh2Ta/FtdWDIhuiJetDcRx
1xAB9DhVoomDHXtdXwTL1FjTYmPPCDA5rhwby72LP7o68at2WBxS9nMhs96Wdg6r
NUYSo5Zb0VfS9gvZ0RhP7DIeX+cfwY+8AN8vZULN2QKrVpdeWewHBsmyZ3KFyQKP
wvZ00Tz8b0XBl0jQY4tMzDzNAwGN9aRlfLeE9I8BRgBh8rwgp4bzWl8vcf2uPkV+
682M2m4iGv/cRNZk9EUFOL8F0Z8KOp2sRi2Fn9+bS7rzkzpkwhbwoDo29Swxlqkn
GXGec4tQIPozzVDRdNgd/2Zsf14ZWhg+SK9HD3jJ65Cj3PC8Sns1YGwclV9LPpP7
/V32AALRg4CRztEXyDet2aftBpRXw/oFplgUFwPeOZqWMEIgAmp7KhJVbrSLNMoH
pX+pr72ojeSGwIskWzCPnbs+n/Mb/W73KDH0wrFRRm92WHj8AQ/kgQZB7rqunD+8
SxwXTgCi3G6jTAEjdfMzDsISLPFC0R1FxdTMlgq4OsgQvMldwAdmQvshMn2oI4AW
JPS6KvbcsxAWCxUnIFlnlpEy/pM6SUvlkfzkz45qEkwXwqshHC9DddM171tPIMQO
gWaX7IUDL5PggxBVdZ7rnuZ0cLqtzpwEX9JlGDLsJX5xUI8QrtwjOw5qwy8+igf8
1lI3CPP8uDbPlq7Kq/I201dGyzMZtK9if/Tqsbdol7BZVIRYN0fvj6Uq7axEg3sK
sg0ZBClkS6MVJrYMBrZ5Hy2OnfZFo1hEJeOQm8/D5hUVVK1iwrErG4BYlYeyErre
I+LsRdjMzxYFu0siuDF6kGBCeoIRhtuMz0vTEePUpHvFAEuOpVOQb8L4NEpCsuME
w3PU04WwN0Tu5l5iRmvpLwrLaze2rkafsCYFn9J9PRVu4rc7mILxh4y74n1Ac++N
BGZ1i536Y8TJIP/zd51N0A28DtDKcyeIhMhTTi5yFjfJWNfvAlCir796iveMcVws
+uNtO7j9AFNmlba9RCYa3mcg+tIvoFjMVtVETjRbHYQ06EJ1jevXy8RcVfgCYL85
m25KYX9g8KLeTe9bf4sLzMUO6RBp0abywg8jpT1jWu14F9yXHnLsy1DSLZ0vBPSG
C0T+RkqZnIWCWjJouXLlAOPtrgzWcWoqIKY7fz7cm2syM9ZBjZaQLfxpxT8ywZez
92hwVm1p85asc/VE6C080FpTq5Q0l92HoxnfhxPUi+sRUoNYQozAqpytAUli0j4x
zRQg55DcLjEtodVqPVfLsn3rpoJmI/0mAqeHaj+zxIOXB7l+zs5fInOUsFmPGqk0
h+xtOfdBH5KqEJVLONd6/fjCrB23HQJI9hmYWXCYGRF9eolK7QpSOYZ/VlD8KRAL
ZoVW6dOB0JbuxxbOjkHiTeqrQivuKbkIIRm/Q1Qcnxd2j01UDf/xflD9qyw5FYTb
GWJuUfY0CTA69v7oxSUenvUwr8HMHYD0/lat241jwEon+btqk+T4K7QwEaPFKuoS
1vdQ4gZTqHcHgIoEhIr0B/JTGt9TVbjkX70eW/rzkiF9pETf/8bp725o4wXzfsto
k8fPusooqV0fNg1T+kL/NtldbHQ4PNWUkmJul/qvP1ov69xkg3LNPURwmy0+Opxn
iGA5I39ExIBcWS9H0QjM6K0GYbvfT3xBHVLmYvKr+NvXIdGKy20HNqqI+cBHyQ/9
K2rVNgTmu2yk2Lvgy9HYzBe5+ZUjx09HLkipkvxDfabK7gklk9cogZDBAnEEKEpF
ebGpGAFLMZYCONkWFmufnHyEoWlHsczba7fZeWfo8sHYS+wFgemvXGpIGtH+jExN
fgd03rzw6MwghHHMBHrt43jrWfHSMYw5hcjxb+ykXsVNSoXxpRw1sLjuiWjI28Ff
H30QkvGawJ5orkikUUMn8B0/tjStcVMh2XtluVNvQCt7SiDeKuamaJQ4BxGq2fQ/
HyZIcgwV7GwaMmFFzOXa+o1OtF4+KUXXJ2GtqQC1NHL3dHxN6r3hayIpA+IqgTp1
n08AFAqjfU447tk5a0z7d+ssWA1M+H1PEoFNyOWktFlSg3KMgzosFVhjAjQNVqnM
5uysUuukABqSoIC5wXE2F8d0Wc1Gijiq6S+C1QSH4AQg+i5liKzc4zCLGtg1kyGr
dhOnEJaN2lReOkwzZCeAcMT/vCWyUYgcQuzgWB4Olenj+DVHXNiREqnO5OvDkC22
XrOxGl021oibjHFhjgZAmAfphGlsQcxeQaVzNhxl9stYj5604zqpUEdRqFvnOhLZ
7850qW0WZoGeDxFUb/7Ag4a1oW71+e6nrslPtchAJWQKC5FqV4NIf9oJwQ2ZC1Iq
auYBnQuw+LbDKCiJn6vhpyWz3D4qRsT87hjMo9itGfM+KV32XZ7bn295smmTUFIL
13BCkoZyJ9mAAqOfMH0vV7NY26Js1j60odtJ0/cFaBxZxrTh70hYAgUTcwmOfDdD
xqnqQ3fBcDkS9MCzUqH9SvPG33DSqGaJiL3Jrrgk1eS3wntyOqXTilA7o+eMe8S5
/SeJZvmAOrbvK5br089v3g88Oe20I2cDdq9Vqskb+AyGoLDRhuYLJ7xAr2XmgjFq
an5LiNMe6f/2wEGm3SotBUTJIJwkqOJfOdWuxhiEsADaxBpfcTkGyd5980vzd3sM
uBOCF3OauXSXxFkzDyT5A2q80QLLIS+kCQDdNtJ5/Ou4nxh5Do3us/gM/YRboN0V
bSDqx0It1smLXk2RiWoqESMurv4knD/4hAOS3fVVxUyy7zqmXnCYQkGi80eOBX6k
5EXyfD5JO614bY5w9N3F4w/pCX9AQS9wvy3g9lMnJY7NsF+iXB6gTTr4HWuMG5NQ
APt91sT/Fbc6sCP7LFpLV192y339IJNf5CbUbrrlDmX6/JfwiCMjRo9xF6avnXBu
CPmB7tcUCemW/0l8NfNsIUlkt0BFJaMsPvvAID08T4E/3qFElpnQteyZwM1wSk+S
NEaZ+AX13RIgEtXo8GTDwDfsAJ9hVMp+lojxKb8zDxQwesY6ZN7AJohNGPYkk0mU
3l4GfRSH83Sii00Uu7PbmFhE7veRQ4olRzLHuOqIA+WNDZM2EBJga7jqplxg6gGd
3Zt0DI27EMAKOwTasg1FxNh5cR/Oo0QYkIzQ9CixUYfE2xbvVUT2q1YM1KPgVOZT
x5ezOUHmHzYR299Yu6rMQHbjI8XAmrDunbid1rXpatckaVDAFlctQCMENXlPlHgI
D8V5ChrpsLkkyCXJ7+H9ce5PH7HYGubHX5u62DYEOYGyPezOf5qqmsBVCMvTC5xX
wfZN0mhIwGqJXAesq5nkFllJGM0s3VNBdf6eNJeW55Mkw3BcFek250k2RnXBb63U
Z+FRN9GfhzNK50LODuVWEgF5kla6xmu0T7LKo1aS8KdnQ5yX7v5IoeLp2V8gBWzr
Ud40JXZpyV+xIfcsiviTgBUEi4lpsKHEnYoSRSu0tNky7vO4Nwe8K7cizu2cIWTG
3ppzy3NYz2kYe6WkSXwthKFu286fX/wl9NrvgJ7n/2+SpKQa3TsS0agbb1F+r43q
rfWQvvhxC4Cw7jVEESfTwO6Cj56s6QrVzY2Q0GDwbK5I7hdRxIsDxn9eeJZHkf99
QYZ/XnbTLdbuvnhnGnJV1l/FKht3FTlw9CHTGBDPL0z7xUJStVtvkWtmY3HIGet5
T383KA6SFPbyuH0ms9eoPJkvdXFZgZk2Scker6MTaodJOJUoefW2S19qHuG+Huvn
dBxHH9VfPMea2aREwpHG/OvRJ7JLJ58mnnlKt0m4ojTMdFZXYfDpVkh/uaNYqD6a
8VenXn+bgrSBC4UkwTUGBEboBfF8HM61gLEJFdY66sKtjkJPmK+plDcy6UOOEiDF
FOzoS1IMi/EC7D/WiEhZ7OlvdYpUxtA8Uv75VNTuFtHc5UC3vdNvvy/l0knwoxSU
bpjKF2dUY/Vl5mQ47SXTCsGKOubWUxmdyJ4MXVuROTepwzoISboHC5jXFAEpKHxJ
+K76lzMysGRV4Xg0KVozf67zUPMx4FXLDgRmIKYDkq9Bisinoklbo+q1Sr9rrBb4
bY3gt9NV588rW29NRagWeU1Chx45jMZ8SZDhbEkmlo+OUJ9Ndih7mijPUWjd99PV
sBp4BnpakLSyfSr0mS1tf4VxgUORUlZxHPuTWbyJGGExdxXbxezDWIL5AdSOSIAO
6HlGJ61ZLWjhIKRGwvvnqPe0rw1cjH4ioaT7mgzaFU/4mto1LaRdC0UL5Y35kiUD
7z/pEjZQDxWBqp0AOhP7bBK//oCBFHZWwpEMuT1xQGUMbw/RmDRK+9VMyzvABOPX
T1MDFGwJOfKQ0a1GOVGANHEfnJO2bd2K3gO/MyW+Rz3pQRAemHSivfKLKa8pPxKc
9XXF93Sk5R2WdbJxp0W2+M0mVoiNyDRMbUsAzNwfKMPC/DaKfm3d5UZa5GtezrA6
sXTWDY0zzakwoe8oKSceVaAesXYdGvV9WgAiiut45hVsMRC6Y0pdZWRgfxTDP2vz
NcfT984LlhBe1Q/KAvDDQZJ611op4W2v9uaS5KNOl7Fas7iLSKhng5Q1tE4haFQp
+2EMi4EiKDPWh93xTpiSqFxV17Ekk11cKGKs/QWm+bpB6xwEejIOZgeqx81e32Q1
bx57cJZLpCgs7bhsgJZfq0e93YKdoTtx7Ioj0yfgN41VIY3kGuORikNdvLXORbjE
Zn9ksTifNOAr7Y64kpQN3TEvqsCSJuhLmz/lMXyzd9KFwHxGhZAvuTenRPjlRBT0
iH+T0zs221vqroSocK3SznlPexJxprpMXY4GpDgxLqtNHykoSgz9KNTO88n/nToZ
WUfXTJgmiQQNd8/x3LZAOSqMtUXR6ROXu2MAt/SjGQ6J+va2fkWCYNMA51XJgo7s
/E32islTZFFOeRMyekiMxlZMARrDIWEjMJRJ61CGu1BbSS+KHWuNS67HHNXDiCmE
2gL95NKzQwE8bsI3M3mPxDOypwa8IyTo/o/BX3wL2TLDEn+DgZ/9xmvFIWFOSkKt
BmF/R43s9gLlN1bFmU5gV3uILarBXM6/NUbG0fYNwdphfIc6fm0dX/5KX4K4MSh4
JN4pf2rJUykVbnqUQzjNuC9WjNAeiLO4fZBqq7CQ+vIBXLh0j4LKjy7X9+bQfzqj
AnXjkF5KjAGKJWW0ocKTwVEe2GF1223+1tSYzYtmWHB8CYhvsDUO6uLPqfzzHEhz
R+lwSR9UHWGjAUn0lKAZoOFsz9smsZvVdwwlcVy5OJF5Gbi6QUtINqZ/2QvHpQ+3
DVDjhUDtUjccoVd7/nxqFJYSL6MVR5rjs91kod7AULyMOxyq08iaaRGDgqFiL7eQ
yO23w59AS/jQIRQi1qv6147ZgbxUmMrm3no6FcbQ9nfXhZnMHj6gc10JXj9pyj/r
/o5a0uil7gU7UG8e4KU1HRtuLo964XG6tGcXHt/pfy6Xxdtl4GsYSVu5WfbYaBDl
2decQ6Msx6jmE2iM6Qtj+Ec+mLNk4iGqSWAQ+hqvr3dLrizndCYAZVsPRS06qr/9
EFppoBqIECFAuDXWei95RV3V+qOOZsIAcS4rDTVJf2qN17T2zv+6ao1ZKHU4+vzv
vY/aRYCykYSaLngCFp8r24RfLjGvm5atjLDfx9S1JM2IWFYZcozcvX1Jt66qKr9I
atnwhL9BtdIRHvJYzqZqpv3kGML2xS3cSZn+bVZ+HXiywMivZZE2AalMj06bbODM
yRlapbygshd0JEzBwoou+BpNoxeHt3RBXZtXT6x2FAlKiplH/hHrcGwEXiOW7IV7
ekUDFqHcr0gBrZE8SGvKNtfdxBon7IA5XBFi33WpmfYfSEX5bNr3ywHScr4b5gws
Uyniwc6x8GrJTHoNHqWWtgJ9cFOaWuKtf070VNtLinGhfPCf4VG0qrX4aUCS6tvj
qd7nERiyNftU9cs3jNrxDYq8hWgvxQnZgRT7SSJIAlJ9MvVqEAA6alF2uw9VA1IY
RPeXGfkU2JEUzhhOn2U7xtEs9Xtasth3ELTydjY1p/P+06RMwFH27uZ3w1+8eUPA
Ktie0Z58OHSDQVGR58sAa5K+2h91iXIOZ2qwfR0uJMmDB1dny8FxR8m6J9b12jIo
ZBdZ0m/xJHC2AbETkptNeUg/ONFILj9SNRmyYTkyE9cSmu+QjbhROWCD7xVWtmDr
oo8zLNEWW2Fx6nKW7SwsNk9N4ECjDmW7HYYM1j8pJyqipcT5YKV/wWFYZo3y/OxB
JV6PR+1fEa8Ulai10WV8BslGfPUVr8a1FSldvGWGgBMtmt7wF03cSoaeq0gYvTOG
iH8ThImhAqYF+C+hpxE7yyBSWnX0nIEB/hvZB2awHCzkqIItvbICAsgZvELgzYRJ
KXIhW0smb+8QC/L86t5CkuFgNltxGE6TnZePTesV7DrlL58K6kdUimFW5xkpjzll
72WkpwgUB2juGaQUFCftM2cUQLy11H5VGlSpMWdrzHNtgAqY3P5SHciwJiMPQBW2
p0gx3kO7u7SKKAyDOVFEgq3umirYNJKsjVzUkgx6VPQCxXqvjk2jQVLAc1IAGULR
OEAoSKH5A3I009F37HUJgJmqGvg0Kgor1TtcnSLhBGJcgUf2es1RbYChBxvRcZhO
oP4ykOyivhHuoIBIz7hhiAfgtmAs2UYV7yeM0My7dmrI9FVFJDSXdDkGmLHLuUSm
puRcRJhY7M99BezZpoMZDoC9onRx8C+8irEqVZtUHZBV0SucBn3dl5iCcx7TAolc
m7bgQC/redzQZsBH6tcOU9rz75zhFhVM3jay79NPzi40flMJTiIizU7GjyjaSlOq
fUmQi22uROMntOpOPzFSOIDia25A88suBX7TBjP2wi4CWUWhc9GDxB/P1hufJtla
Jyu4p/Hl/RS3I2I8ByhyDmFihDzrm275Nlt/HWn8ShWmAVwq+1DyFwhhlNJt/Gou
Zp0nV1vGD1H0Qwv2uDDWgb0sT7D8obFa5/d+uSSyQvKO9zjVCqAW8E1jgPPuhLIX
HvBs+blH+c02HxYJVVpp8/6wMm5Lyl8wB0drXfdnUBan1+hnTbwp0xsILpR0TqAf
qYPAB+qUjv+4YQKUAcbO6uAlLM9jOyBS3eDk3VEpyyqKWW7lS9HNbvnevDQBV4Ty
3D8zz6G/8hPn2NMS9V76zQKFPpmy39e24coGhRAGYcuYHejcGoY57bS/dIIAjPvM
9I5Czweha6RTNxm9Stgo8It/D90ATGGjwRVXDc6oyOpu3xjMOClL2Jw9aabg8qhF
mfUoFjCHLI+awcTzjFqB5XpVjQuv+gM2Jk7UewFHfuSMjhB3cZVVBckAW2+8VP64
3l1RLZBEI7wdn5cdATUOIXfPCbsnwecMt7PDHr+9pfgmW5NA2rEE/GHKnsjafwGs
gVFpA/L4rIUEWwKBp7FkT9JWppv0GLy1FYV08Rv0kxLBslGdpTAsISR7fYVmcQLb
37RmzhkiLzTg+LAlvalrpiMQDafIt3GzqQOH/j73h9q1thxAVbisSBUPWGKMRysQ
GlSSOlPq9mI+dKBteRKSAmg6+z0+XbKKgzCg0l35T/EmK99nC9M2Ezzv0HkPul1C
QABamFsmEN3bBcj2M/MVEk81+Xj7HtQ6flKOc577AncWzI2MuKUbdmOh9aX2dcRA
YhTmDhQBbABwXIbFiR1G+BndefwwuowGtLiL6mkgRQT5erNpJLtMnoiuZrvsOWCM
x7YEYgP1pql4pH6BlEC5p8HgJTiXKRmOpQxjdoPBzr8pn7r1IdkcS+9sEGDomnuc
SqNevbktZ8pDYRjzotOozab7M0FdbJjzSt2wQy6Ud9a2j6uDHTREOmmcU7ukYSOE
E0GHus2j5/ypjsBIbQRitl4fqvHp17xCyvV/Sy7Ihn0c5O6zm1A1gyiYbThZB6rj
TRVT51WbCTBrqorMdTxTa9hRTQEA0c7p0bc66/Ioth+B9BNiOEloAx4ZdVry4O+o

//pragma protect end_data_block
//pragma protect digest_block
/YzhxRr95x8BkuEqJ0Sk2Q6K0Q8=
//pragma protect end_digest_block
//pragma protect end_protected
