// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
OhGtXNF4Qpn+n4UtRk0zRnn1L9tuDyQEh/bXvc9SRGvpupvzFtWSwMQQp9RaxvP0JZ0tun0Q41Lp
SsNqcqEPmuGB2FzRTKRtKW7jdk3dw3RBUsx3FIOPEMbs6AplYgH3TsKHT/KrgXv35w5fqYQ107Kt
QRaZIREHrVm0q6RucqiZ5idDIe9xHqSnD+Ras03NEXnCXYpr9Zut7edGS7sScAkb4esPsbD4NJp+
j07qt1OB1rDx8lTKj3y3RTEWIn0CwCJq5SQI/bXiWILQHZhchT+U9rp8RjC8ckSgpiKxdQiKIy2J
ZL7bkuJDgxW/L8NnBltbEXeALol9Tq9lqod9NA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 32288)
Rm7ydQZwfBwfgzFzh1GKKA0hgqzud+EED4Mg/b9Dp2GepzEjFv6INaP1mm4ec/D03vRXVlDvoqe+
Eox5gRynCJM6+OhsR65QaGgSxg2aRMkJLUQI1A6h9d2rP+0xrRrhwiJSZC9m5WR6hTilCZMXsrpG
re25B8oLG9j65p5Gddg0Q/j0pP36FMx0zpkJu4vh/ddP5GzkmQbpodPQwiD3MiOwWC7PCIpMHmjE
0k9Vf4d1c6WyRbO5Z6RNIn64wg2gk/9jq+GKWpL1LY9pBxnkBiBHYLXjDpBRkB4/YIHxCCm3O5O8
8oj+kuKbv1juLKjN2PuDy4JRHNE4X4yAQ81kkZ8HA83eCFXoCpySKZUkz6x2GpAmBQ2n0vCbfNXn
DNpjaqMXp5qiaOvGRp1EaMX6sik2FAcnul+LXKesmkRe3MxcUpCze2EYBxVEujGfqC+r/tt3rnxs
haFEy2sKrNXsaUq+VhJZ/k7bc0cOA5Aj3eXu4+uLbhQXxAEFvHbcgxpp9YEYfHFyoUYuOXIVqhcZ
eN7K6N/7V+A0BlmRd0OETn7dQ6pfJabwqDZ5iSeugUsYC246Ve2v8Xd4RriOj10+RBJcG8wx3ri3
JDf1VUEy+TckXT8OeSEHwkvsMY6akEv4ybohDQeowTuZH5jH7xcb/MmyZSCuWKud2dE9JLxpf8kG
vVVNUHPmORCP2QqhlC2XOx6i+Ckaf5qvm84EzqXdzPHETRCrl9XZivlKiZPv0kGJp8LllLVa34yD
9IYhU/oM/8X7fAZ7GrFiX5KGG9Tda9c0EoKB1M7tKmRwptDOmSOd2W4uTobC3g6TBoWx1WCW2bcI
F/9oqWMqIHs+7eIohBVYOhOsz159rgSrHVQJPRaM86YMNBsAchkJ1YheFRpPH3DZV8yth5qsXyFj
mKrzbM8w0u8Eql8QYF+8Gga2NWkJiCPlANuA+H39K8ZkxYjR34LX3Ar90MyQchxv8gpGuBWCLCSu
tOJZt4URlFKk81Mkyi0c7fbHC0Y5tRjwHZ2Jlo59xMa1JkQwEoP2IQtuhlw3CgmPt7KCYcsCplpi
MMhuuuTlc+J/pfTDsZqObMSqqo3Tn846ckg7tZz1ZqNZPx4/Py43nDGyxpCL0s7awslWKY/Gntur
jb3C4yEMP+lfW30BKsKf1n2xdvcl/9kQODQGfOx7ZTJerlip8htiIOnU6Xs1LJbGjxptWWGlB2/b
KfZEAGQtzdSbMZqVw4aokf8BzOMp0sfwf6elkrFS68TZq3N8PiM8gZSVfLgPqvkZLdM5u/nwiNDb
ffGZwInVCKPrUISYlJQTUIeRnfvtJPzKSRLrr0R6yh/uptXIzydg6Msr0tKT2vLUnlwvm8GpM5aO
EV6XR0YFx7Aw6h+m9KPYNQw0L6x+QaW0xNL04HBE2Wfdz4N3UPGYAdpltRo4Ea2QdH8WAVeaDxPM
5r+ky+qRZlTykk5hxSju8IRL5O/rZAqdGk9lzkGrXtviC4al/0t7NVyMNqojikAX6dszf3gqeorY
iTmldpA/sc/pykdPXRTpsiT2ZgDN7cKcrRyCTUbY3OK6sZ1nMj1V16hOp8U4PvBRvT4SZUd0C7Vs
Jv8TfWvB73lFQdUXdy/sVElUmUM4NxvWtNL9WDmEhslF1Dm0WE8IaCd9GHOw/jKyKQ9X/C3LkY0G
WPcD3bRa7T9Fa98gJF1x95AANnvzCSFyatnWkjPmEerl/+3l9I9WDOSSOurBS8O8jQoO6rP9lzQj
D6nLtwjGzSyoQO4lCSziCRCjeHWwY8o0peY0O+9o5ldG+fLHySMrozhu7Ko3AHDp5+G241ZihxIU
bYyXIH4E70ScLkM18mByvYgdsABcDgDOAidtSmQzJgjjBjWOX8PB8U0BxdRWhVMVFw/VE02a+H6S
Qmsgb72vyk5R+SvyoMxiTP7FfnpyeLJ3pJJYyl3kulGpncQIIsiTGwVq5eeyRa3Scz5PfN0xGCN4
jAsDOvu2KBk69JsAJ3yj9UJmHXNh5byH+adIeDY7/V0nxv1UAuZwRBMlL7hc0K3Ew+P3PqzTVvqg
LOZCyI10+vxFg6BqWC/AgvXiKIvQq4CS57Fk9l0bH4FH9Ja7BihrkF4WMWqZI0NA5ovEnu/37+kr
lWcfLyrqw7OkGyBfNim2Lrr7KH6S88e7zoeHrzOxQiT2/O0Xqn7NETJkR9Bq8bIpT1r5OKZ8yd0x
Gqt+0Uun7dHQTn8vI9butLw+1W/A5Rak1+WBvUjEKjqTZ6vuGoButJ0GSACm5klV434+ez8UmKHk
IXgbc3zVVOjep8BEII4c+y5+ckggSaBFTLmtBD+VSsXwD8lFvA9Dupysp7zzH8rXtJqohT4DjigU
DlNeZoLqmbUceTdLPRrkCmc1rHXhN98gdeLExweN744Q3HDzzpiLRcsdjuuTsZwtTsoTgH7kAr+h
Y6IsqNffzLXiyOo1+NZkkA8GTc88d3OeQvRnfPjvMrWfb6rtysJIkZAxmUPbMKQ9Emk+ln4ExsKQ
h2HkXqAeBJu2QdSOM80ewlAE7gRxkw1Id8tCHK0ucRQWazCfcZcDJBSEPYmybYU2Y0iOP41UoeNH
zIQy5h/xobZwSvNlooUDC9rjjMuJmoEad041WbQ8eN5xQ86rHPu4ShprhOnSdA7VTBvB4at0hUp+
M1Cy86GvNc+Qj3hqPZEcvA3PhHQOSsp8qzqaqcevsdnQvFEclaR0A9hQHr6Nelrqu8Hlhueez8+N
dDeuX1yWIF8XTaPHQp26WWco9NoIVqi8XmQwKta+FaYNF6ahZdrm+vYFgvfVHJq855hY1F58Ziz9
wDl4dFwopyeJUuXPTYv8stBhXKmicxxXkVb0Xm0zqAQusxfIDN3/2qjVE4CP8n6bLRUFj7XJRo4f
4okq9O0Dj7hbJBfvVUSW+fETfidYv/VymqwX+ZNuPXqoAbLklHVMOyT6jS1X0071b7KvoljXloLj
F2wrwAMk7VpG6BVMnRRXkHXGiSMR6oBPvkGLo0NpBo/Y6xuOEWJUWdGT2WqyGMU8Ot4docnUP3zq
a11c3zPMx4pQ9gLHWFWloB/5M5TIDCdG7egLofJXd4I5b+UOm+qsNFAuUyyw8VYsoVNMMmD8rLXh
UzpakUpW7Iq3BLmAIkSBqMDUQEkJyeQ9rOrYHRa7hFzfxzFgSrJDzuj3TIciVXpqv7mRSuFGSPjL
9k+JfcrLl88bpL6QT65T2M7glFGZf9Aa30Qsqb6r/4CNWfdkoYwwJzu5iwK0Vz5VuH1tpOMiZGF/
J1ifkitqehb0BXZqaOeMWJ1bQlenDldrNGIjrDxuEpEqyK/V7iWMLXZ3XK3jBZd9NiDV/hTs5M0V
plv4+PtyemlUAOIbCSQBwSaj7twKrhKNDyi34hx1jdu59EZTw5RYf9E+GBh1kXSz74aPV5QZCJfE
N1Aj5J5Ez+nElOAOludV4O7UhqhVS1Q1h0XMHfAFF1U5F6plqCad3F+7jhlJLbBm8IHBfKGKAewl
zYJeicHdZNacwQlDfyuOVvJlCgZWmycgdu9FzbmRkQnUUjfhCS22uxSv+ny6URJ37nm69shO0I5J
AsoEWCLoEtOtHzsRmMqmRzvdVf/Fve58Au0IkvoHNjexA5YOcUKHxZ6hsmqwA8yKQmSwSeprPvBE
KwNGc1X8sLA8j5UcDn/fxlKqqXZadwgxsRHkZvNdOC6EHF+6MVgQ0kxf9IEGrKPClfLEGzZBB/Ll
93ekAqldE7MiSt35n/wKene5bT6G82pu7uBANLfJVyDuTuNyCBHJssRuhBKvM7V9tWjhu2v9rPXh
Kc3CVw5MXX1dCIrOd+U5om32I/52lb1HapSMzeLbOqxvyKON5fLPiPBikOKK0GLqos0pPl72aSmB
RnEoG1OOvSeQMxzA6wvxyPZEqIbzWLy4Vi/PhaCHFhJD70zwbaKxDsrOt5kvxCf9LwAhQI0Yrnyz
ta31VfMJE8cU2rOwH1VcAJwzXPWfDDQC6HvWQds77QOfkXK7tRi0KBD+GWK/iXBtnTGSEFSu4Qqy
Ypx0pKQnPrDaTpDZxWZ9Pzlh5K2fj/i6Yc73/kwc9s+0v13zMXE9ZcMteWTFMQfYTpUFn4AfRvJ4
njPGTSidtORMtwVVaStvsbOIgTywQMKvU+C16Ge6PVscWmfOn4//WyU2+hdgdmcdgrenA30Nui0S
NWlZwQcl6blpTExd0oMraMXfQLlL2GdE0gN7GchsFmLLlLKzdZNxX+AsOf9C7hLhQDDN9zsgu0e3
TlJXFygo33ATRMcCyfnEwnuGHHRDpk6v4Qh3/DBNeCKN9vEH+diuY61ScQW+JA9vSjjFjpE72CkY
iKYhOo8Pvcy4PM/Sn/4zxsVkGrBI0uSdgA6PJtY7JtW3LT3TBQtczDhG9arar6DIr6DyofVktObQ
gWv0Ux0jC29iLtU/a//23ZnvxqWWIiZvywclilcAiyKhJ1xHtxGtPeIrHvMbng6Lqe4TKuaXMaQ8
GdjxI1jGSggI7P/JgpW9f45POH8JmG4pl47Bt3QMM/el2EWKYfIx9JNyv4Xp4a2SenqjetDpEwad
UCNjWi0GRJXIxD6O6uOSDvYfmBafkcXUIPWWzWpo+B0/pLJh3aLsUyAAr0GFhilLvxRnowLadO2b
ivSSuTTjNfWgOhfk6jqhHt0j8ayr1RRQHRnC7aF47U/6Gi0twDN47cAth9LH2Ce/IiIbuRYFQExA
pjFxLzyJH1sAYSGSSCy+13TWSX1dF3OaHVDnXYbNo1jXweHD9Dxz5gxEkjtQkN87F09dOgiT37A5
h+gmH7lb2Nmz+ZI/ZK0+pvhZRvHEp/2eQq6k8DbmpfLAZ04feq/JEYXuGg+e5+4FBlyScLEtbZj/
gbpcKsaXnaYSp9aRp/sp5zkAdWLjH15OmjI2NZPzvne9nbiJhOgWaO7XfSyXEpDk1D5Miy1FnOCB
JTxvzTC+I4vV5KWp1ym0PkUyRS5WPpWJRo+1XmSlo9l+vA57VZC5d4SiPFgUDHxNJdbPRU2/FCsl
6aDyvXEL4Zp3ToMcoJo+aGYShPtMrUHgY3UzVF2irGQb8pUO6Ntdygvge29HefhWyTJgTRvCXyE6
Rg6A3Dcssz1KiAcXm849+SrzUjfYworbegtObF7zGERuVAL1wYFfJILIW4GSqfi4xtTHkV+/4RDy
oenZ+SftFA14PLXqPOVvysBo+Bw1EILp86yUuVX4+4gdekVqy87P96Bvg/GeKoMPCkGfNs4mlTCx
uCxCujt0FZsNf7CIRMnrg8YOJ4XOwerxg+KNvfkorNCqDY2srEC0ICUL+46hjlusTGZN2WkALD7X
H24B2NxwWoLW82nJdUx2s+VIQXMeNOy2PlX5h0OZlygoNMkaGxEU7q4Q4DRX+VsLqVP1ynqrdNVG
TWkhEUH8Wq7p3k8Hi6v/cGDIuBhu4o+q1fTWRabaRHca8qdVlAeYLo3w6f85niIaaJMzHcclR6OJ
0m+hlBDwZbsEMSG4jjpw21r3J6vzzOKoBJ9ctTpiRE50REGprJNisuRspDbtUdU5Jm0gNKF0p9io
Fa4tByyo10zjuinvUrA1eTpdtB8NDv4H7vWkBpYVs1lJixofTl2TX9eKibJyrxc70V93ats8njHc
VYPEa5cdjj+TXpb3jA2+8ago3VgjtHZO1LIkPNQfU+JZvNdNHZjZjA1kJ/dT+OihX8dU/PhO0zff
hbr1TkcdmYuhz9Y4gABBIJc0NTmhmmO4JKwvaTHaT388/+SaLCboTKZLUjXYcxJb1+hjvGerhXpy
dMjA4RZptLHdQsA0htAUJd3rfID+ZjVtUJASHVw+8uglInHxYstTOZfxhaCLJfb71rWMW/EY5Y86
uTictVM0NHI1CL3hzlIle9f+iXAB5UvcRNIxFW4KmyD4bigQlbIiWwJ8x7XUT2+xhRX7SXkLKyjl
hdQK1fH1NAQXrW11LRc51+0NOcZ5X/oWC0+YMHY7F0n74G9xdHJEgooPxLriKqpeu0aFXyxKsstm
0Sc2/ByCcHr/EiuzUeDls5LII3RMZgb5VcalQ/iPBF8fxLeVDIyhqOgG8NNhX+OAO1Uf/lxxmbMO
zrLPCq8wCWkbcF+Dm2YG7xprdnB5jgWoX9ywabrL41hXg39wPfKETbqChrIPX/8c5YjaUv29egTZ
IV/AlaoHoLyAF3qU2TSx26ntEeubpRqt0nT/ZzsdtKLliTjLKI307yTJqYEiaHoJi4pMCWtopseh
kRsO9JKjYBb5mI4ehuadk9Y3x6CsxBc8Tpj6f/fCRFzO/i+UkH46UAMMJRWzEt5w9kEL+o0IW08x
Q6bDSgi0V712oe29HRO4nUhir9KRWhGJL4Kp2EY0oHJ1kV2rWWSf33FFQvH0grLnL2i4pewKEt3n
oladvRlBqsd15dGxaxIKB6qUgXYf043Q3LoMNwTx8geStn/SUejXUWqm6kNc5aOvLaoeYHe9pPK9
YQxIGspF8ulGKuUrgEW5qgh2pMNvE2bvPQBFCZhrNWC6CuijHxhSTl7Icf+3rKKlakuDZC1D0niQ
YlKpygx0KQ7r2MpQ6GoqtnbsJie1Ls7zcCL3f96dpB19dCz2wzj1YZyu5LtqqOfyqlv7/r0uRbc4
rY34mKoZYsBBLoMp8wOnec6b3xeNg57FbO6Q/ACHE9KI+54EMLlBzavfM4A4EuPrlcXnXwwx2vM0
mky05VdTdZ4txAyJQfrXMYs3aZopEXHzjxVr88VmaJTygeaFQ/HHNjS/zyIUa3XXL1Dif4fhMXUR
ofFX5fWBSYaJCt4mwXwwQUgmRbTwokJoGQ5yajbx+EynfrgtOQc4X++XB+hR7yIQG86oXVeNawOQ
b2FHCBsmb/8p4cXQQEtaSde8J7GUeAp+wq4sfX35kH1d1H9TllkXtYyXCc9gHMODitW0kxok0y8/
wieLzWJSOVGcnZwS/oYccyhCWxBHg7NKCTmuFPAXZ/vsZTxZksjT9d+ShPJhjfHhb65rRH8sc/VQ
t6P4MuZqhLNk2lHyKiAjgHdkncZT+Q+6qbdHCsHKDleiozZE/RUD/WNw9iAtsYXqhoiQnwgr/F1B
Wb3lcwYLeeuGmrgxYAC+qy8WtFR+qy5mxGTIbtECfkExwJrKIKapVXCbai0eIQmwU0o2orQDB2BS
QEbTgOiB+54Q9r/egyY4H0eDPF/mjOXhGZzGlKuwuAc0pUKb5mNuhVuoUnRnmWDfVtnJschX+ENC
U4nBLyDjky0nsVbNicT05+nQREVYPR6ePjdOUUD3IXt2q+B4u8+D0BUDWv+NzBNw3swXsEwwgeYQ
H1Ioa54ip1DFBWhAoGH0sb013j26/52jW5yMw+YDuMoTY6phRf1pfjwo2rTIL7ESuYEXeWXEMITO
lHvLgU+88xaeZl6O6OHhc8kFHMXAgoM42rRRcIoNKPGEGm47eSg5+IiKmspRIhMp6e0cvXlV44y+
pLAruzgioaWnPpRShwhMjhxTPfRihfH+D9aVZRJxj2ML9ath60S8xuE+1X/p+w9pDcwHtNQbO1DC
mkC6KqPJvNdDvIs7om2Jeybvx5XDJ9OQ696tiz51ySS9NU895DJzZCDui65AvIl6YDK2vTu0lvAF
RNKv0xqPa2JenQbWHh5CJsc1Ja9liSF4/5LAZiv4sI3MTVIGkYNXXaQLjEbuh+QPloYbzavruuQz
1YOBmsGP8JqUq3ggdqvxnnqhFhf1dxOVt8rZBQezTlPZnBKq7/UmAAgOCfk5/mnb5c3UFzxRlVsT
5L81YdGCKk5+CRaQN8cbVI7Jm3fWuAhEmLuBS0L3HAdi+3oiSu5Tx+fqQajKp8JKF7vH6O/JsnGq
QTgg9Um2ch6lYoBUdEYu1koPDFlEuYusuCyexVFV6VOMxGshv5qylH2j0Zy0nasHEZFxcmT6DuDv
1F3uhjNEEcn3Yd97EgRiIjeNTCqQ023zU2Jd456oIjsUTrSi5SLprzIp4q84uJFDlCGCfNn1dNSy
iGHqiqE9A4WfefKaksDm4L7hk2dYsn+V2e3mh+Q7bbpnmwbHkwrO2P9g1y4d5zEFnKj+xiqfP1yB
v8sMeYlZUCDwTzphNpN/5ikSUgQz+4o6sNUUhlXUn1fQBvqgQ6pu/F9dfsrVDP1gJK4Pt2SDDxge
hYJOKtfZ7+FeScd+cwJPVedjkge2MLC3p3sAEyAjLAAQwPxIxUDPQXO3zdRzVkFKu2ZvXwLG4K6S
8GmlGQhHxAxkmXyIKtPuxMEYMUgBbvS2oLBryBYAiRNU5mek84OR9XLmuUjWO0AvPJ14bs2y1aCw
wQjWfqusbDERXF+3mIHMBL0tSHT120TiX9CPNCGAG93naYJJWShwgFb2aOzCyj7gDhnxrIwzB8P+
BcVRLcR067VuDzM0sb2bhNtVOkZ2ETe08WySNkfBbMfbiMP7d5qHvqEgILhsI8V+HmJ5PuIRfZx4
XQIx9t80FAE/WcM2nQdxqusnYfRxQU8mv3UpL8VdAxMybG1wz5cYdgCL8qwisY/8aC2k5tlBOY7m
g8OftOl0eyppr0zP5iMiOcaWGo2EpwlxrcVTQDclVY2DBuDjc6riLQpuKIIwmIw+QeFfa+A3MQL7
W+3tyS3itV70oUTdMG5RuuvB3Re5xRM4LbnCQ/s/a+wGpk43zqjY9KGo9eAU3D7UP174HloaBlD7
EcDamCrfEkjt3Rwz3y4NK7ogSqG7fIcYCwyrz9DndH0QOjwOOBwkVlhzTa+8m6iDxECWZeARAHlo
e4ZdN5xTMiQnSntzNz/PihgB5ogmVh67SVcaw6/Xn5bEqP42dhn3JX5YNDAoBm0KbAIzILFPJ9Ff
3PZXO6bR8GlBTb69aRRQsvJXjouHYEH6D9lVTulrVBwGsaOa85FG3Nvy7KT9KtMLZkFnZa0EBSXg
rBj0XoYC84v/lsiwBnVc4gW2QCP+Dubqse4mUwgQW0tbPUCA3okc3o6vSz06lfzk9hIWZALD+r4M
WryV/iNsJyddJ8FYpV4zTV6no/FJdfvHAb3jMmpkI6AgFlTtw+n3tKwCrFBr4DnIle7+RMrUoleV
gF8Yk7gOsRvf2tLFmssO8kxDPiBqs3N4JA2IEVr7QqTS4IILPYFA9rgv/gEnaYbFsh0Bn8IeJ3TD
UBc0jVE3rQCis7b1yo0GiUg6k/amtAQv70zq7zJdvSeNXcwWCnFegmzes602rIyG6gkItJap5yXv
Uxu7zoFwOVIN6fjT2zJzP3eCprLPm72oEEbICmbSfhqddnYq1y03RCwI28nVWqpIE8D2uNHmcmZH
BlT90YL9Vp515aX935bRbLxOpg7fc7ZndSI80B5w2htGga9LYUti8E56LKZA16n35yvFLT7qDb9B
oUnuy8F+9QO2rVRGIFS4sTrRgE7bWT+0fXHDD+sn2fm3VtrkqCeQUbHF2eWcsrr1Mq1DNeX8f6bU
5gmIozRBXio5/SI55j4xbyOLBd1PwF+5J/BMxRSqDyoNUWqNtmyaxvFxencuEsxVS8YUQmKRqr/f
nLQwzSt7y9tUHs41aG5nkNxsNocdmi4PieCJSnFcm/B9joGwUaoe4zEBzcGXxw1tllkuBmQpB1bH
i3bXavGgZF6GpKBVLEftsjStPzVTt3BcJ5pZCzxHc2PLlLqjXESg19y8gdtpkh+cDdDiVoZMB0up
MrUmCkI9WdKiQlfUFtmcQCUcwu3Q7Mn/OkSlX85mVrbiaslkgHy+X/MwQx6a96PrxpzNzBuDYNIx
rFODKsh/WlQHu9K7+93L9AIWQLGXOqjhfpJV9lg8MpTx5+kLl51zTPpHb4dhSme1HpdjvnIxKWrn
xTnI5yvpToTKOYrg9UOy5F2UpL1R5/Z3LeFmyCMabb9Dd+oIeF82t3eLM5zJGBV0D2rcqQ6pDh8X
Db6AQuum/qWGVphiQIuRyrt0aHz5qBQsYMmQTO5BexcNzgqEaH0XvRs6dnMhlIyczMbmc7HGDDz0
xo7kRlr9GchVMTnYZXNAistveuaUNGgTE2/k9O8fh+VvXnWamy3w8wj1MnoLNlWfQgpGJPVgVOm6
CdrjV8y/06O9JB7jUlZmYkyKlilmjltB26YLYWxbvTvNXEeafFZ8dK5PubYg392/ulY5U2NfUu8m
SQoPiVnph2BBdY0v92VI88pNvWBX71nWXWm2UY/UlnVuwGue+OMyDiBNbEOC7Y7v/tg9xyd6ey8d
A09V98BGWMxYOmPNAkGymVHK6RWn8VsTzrhTmFbCivlYNw1b/PwBgz+XpfjrZKqfgsb4e5BhcW3j
LrMIRB89g1Bb1AzViJNelDXe/BiZfxEdqn0orR/r/9XOpOteDNwOGu7qP8qSBbAf++crs89pkEtW
rr/xJRLKqWvuqUiyvpEJ50MR2tRb6rO8wY75SJY2HAHUas/k0g5yGDw7p0a0rrwXHX3IHqfHQi4W
a0roAxsgUZM5f1BcLqK5DJh4fuX0+E5EH613JmJAJegMjRlvRX8fhZB5B+/UiEcXLiT5wtBLFK2Z
kAmDMxSW/qLhtmZ88M+so7s0Kuz9DGnzF+NV9EXZ2drHLeNLBcGbnTUw+d6jBWgKUnZXxzaFuu2P
Uec2wDpWh6AeK3pkcLxb1pQCGFVCjp4Am7kJAojRyvQL0QqKySfDMbPWUjeEASIVGPMX0s3nhvXr
VU8EI81tcyayFdCPiyqkVNdeTHT9KXR+eWhcG/NVjCf2JkxYBhuqK+bn3HpI7kkXlblhEDjwneef
4M2z452lxEgj5KdwaivaYkLxU3IxeTTOBPNgcPpZjol/69Pbj1c2WeaXtlw4yas97EseOiYZpiP1
zuxGWyVZ89xzS9aqLJxl3DfbZP1YuK9WhuobRYSKnl818w9byzFXFGinZ0URCAo2moGSxCT13uv2
FxkE4+KOWDeWi8BScH31ZG55seyfHKB68PFXpE41Y0pfYhi+RcPJabrCm7Lm+05Zjux+thzLgElm
16GBbyN16GMsdUY9p8yt/8Dr2lJLTgMzeL/TcxDvWMXK8Uaqf4cBRxwuhLiNzrUEkedIM6prj2N8
d7Ne54XG23p474pXiDw2u48YY1d+PP+zkSGQ+eBHKscaRqMOztUeXrahsrC7TRaJG/40LKPUbiJq
S85XRJc+HpSSHH1YumXHpF4rMb8vCiud+yTct5vk8VjP4r59odXsWk7lsANjLgWTJE2MaxrbW2sF
Gmc48B/g7r42atDRfdhpEMRElEoy7gmgGjbZ1kzkqxZB1gAVOivVxYbF1X4nLWJQ9WoZhi7xFOOb
Mpk45sMtrmzypc+xLJYNqEriqpvNKleuL/nA2U04+mXuAC5PBnpSjOOBpu3c3ZdD1r/uMUevkxBV
9XSqHiZ4aA3XcRVSqCQlLjFpqjfwrj57Puii3RmIjwkFmz5/TfjMZw13duP5apA4N8csgqM7EAln
fV6ab+ytcMSnIC/NMX9V++qQwon5lgsfT63mA1frpoDKdqecVBEh/UoDmnMZkvM+hFGbo0m8T62p
Oe3RObO4gK9h0Qj7DfnmjWCnAhVUoPz10lgLhPkj7IbVsc0svXX6eDiepYkqGsy0m9qM2mz1uBzk
3a4ikismxP9qzHVprce33rzE2hzjzQwq+Zm2WaURwsZrEv0bUlgkeYIaeEDRRHtcE7Qzcu4U6wC2
aB5hFZgQx94wubMAG2dH6xbEy41qwn5igdeTXZVSdwIawrpoNOCYFD7C47SrD0mSjJyuVLdW7vxr
2wenlUtRAFlKoXIMkNs74HUp+dbUexUzUSjZS7YDo6rmRI5noaTBxpjxiPBJgKhXLTXDwDtZPunn
wLi8uXcg4yVPt4b5pwhpf2bODpp2WEgp2ApmZwPbOuubVT3oISAaWKHDUYS7Nl8ViEfFKrPV+L5y
zmyFkcrBwWKXa5XRctQFNXO+Kb50xMDcldhDs6CbbvEuYTB/2AsQDqIucw3+XE3udHnlns6Nwqb1
3PxK0IprSctT0KPnwgK6ADG1c8MYM2pCQh80JGoeZ4Crzaja6gkOvHtX89do5UhdZv28SuZ316TH
9kxU0U+zNqtFLHTGQTmUczh6SyXzSkgJ7Y9kqYT/Fyr7wchdQ5dLfadWuKluxRE7VCwny6NpMaC+
WVnEQnFtymgq+8/kegdsNWfKMDjdIKvBEd/ArE0ckvnQYIEzvahW9QHtCBPu8Mt0BEcdCTtKSQA1
EXsP+3fg+gO/8721447Ylqhd1kw2f1x/9PejUBPzD1oUgCzqWEFrfS8dg32aN6m/XQXB7aAb7V0b
uc1jt3qtGv8GBS5gtDrhrww5tNX8RBOFURH8b+1tKh4meL7ka/pzc6BnS1C0Jh8D2NqvCvRyz1xV
xYhmt6sFkNxcMKzWqiJWgcSA6Fb0gkValXPbYT5yAMAWaQoYeNGCNib7I8PAnSDF+F9F8cfAJfOk
SMV3wzhZQ2XKuMDBxg5QXZqSmUPPXrNprqimo8lvgHBLQXkzIagZgbOIgZQ7+D06Z+aK9ndBhd+8
LDns8zCCBAXqrA8+oKaM92MRrAkbflwldIZKES62XUq3kBBpKJ22lPldSN7It1nHnQ6/0sRLJqeS
V54gaoZwQHI/CNU/houfNFMHn5Nc8trAn8q55V3CmjyKH1hvcfxD3nKHZp7S8bEX8trYf/rcocXi
UCGMVPzyzvV+PdVx2xxpqUTUMVagbDkCpy4sDe2CsMvs4ZUAQd94FKMXAaC2skuXenUwiYNsVHtt
t+Zm8QinQGjeMmRnAyaZ4URDr+vg74tVYVHqs042LWVZn+NAhG+bpQ49fWHfSDnQ/rvkKRJ84b4c
VfTrsNgZm9ld9kUnSHS9TJhQwxQgJYM2zZCK04D5DevGRzGODE/LRF2Ldc3u8B/2Cpjhw3E+0W5j
UYFALH7uGa5YwDxkFv78fOT7FCZeCyaC7tlcWp8N2i2uCjMKmkXwa9T5KgaiB+Wn/+i7T2ixumRV
mR63mv8jsVyM3bVWM8my/DzXAwrHfg3q2iaQyn+3R7hNrKqHuhvYjNRshVOraodeOecNOURWWREa
kkhXRMNn3VX9pyRFZhMrbIbq/1W1vIb0McgJARM8Rh+eO0CPXVHttANOeDqyNTkR/+vJpp4D3bCZ
kq+o9woPq18tZqiJt6ABa7Ngckcr/UhvJPDV4L9EJ4wAJMvoZIKJmcKpDhn5eDO9ynrF5wbsoVwR
6HMieXxLyM9lOwOxIyum4b9jPkjP3HWxGYK6g1YHVHdAwotN8rLDzjinkI3q9eFQ/ccR3etqqtgq
BanN6w2a+dzbd+epnETVPRsuaNizqRu69jLxGRhbN2tQoZxxEhicCeDn04KLqsfTWSvceAH0JdsW
06FNZZ0VKLjUkZuRSDcszKcFYx5n77LI/faMpGEa2Tu1jroQQefMICItNl7x/AkT/koFDVJeAEGD
P2ctaaZ7kzGS7091s2RoOZgQNvHwZBrPopE2Wot8IplXv4f9CkLrNOdr3bwqOeVe2QRu4Zf3dH5r
0vzSdAtxjyI5xSU4pvRuqKwjibLEoHUDeU4+wcpKNRbk+bVjAfQnmXb3jU8B9KmUVgHa8/ZDPz1V
eWIL273PxXTTvv3UsUBglLU2wOguJFsORUi3nAMUIK1kVls0PmGUc+25uGIrgEmYvdS6gYXHOwtI
57S+H7wNKNPOva0IiQMv4al/8YKdyQLscmD8PMcTdhBzDGuobfZkwZIwSr8h/Bfnstv+dl4x8wlv
oDOFkwTQHV9qckcq/eaVynyCEcYpVgUbXODQAeJXcdpbwFpLY3GbJLUNw4YUg2PJzoxjHlVjeJ4M
HjdwfAHHkgqQSPXjtBJQ1Y2jL8RikOk1UxZaQmTAgGKOq2XDO2GqeVc1eRqiZKLtZRUk5++dtHtP
PeEibVg6b3mU+/C5kuQkCr6AIvGdI0fmboLtMzje7tRT9VNwAaX+Rf28CVSmwjcW/dUiDxq+P1fG
g9++Q0/yB9SdJlJBKrSxTI7RLPv7iWI9CFLOy+VReFEwS8xjllV5kbKp7/O7+cKdWLspfAdXxH8h
OfImat210yxXDv8R+f5YZS/hanQXl57Z+vfwraXVm+L6VUtT11ZpI3ZZ3ZAtO3C11k/c50mmOGSR
g7jIh1LWwh0Mf9UoarvyuNzNZ+2TrivTwSXgv9NTu0aBZqvAPFdl+HPEcc5kPxW7sT+ipPyCDRvu
9DZjyLNlkuOXK/b0KvsHCSsmtW27RZDUfStZm5AhkZ59l2Ty0TZ2JT+efc4hU+xK2314bewJWvdG
60Nn2s100xVrIDyp25F5v1do9oMCXlmJ0vyWgdH77P7WG0bhJVOSLmI7ECFSDZYvAKsVi7PbXZkf
W4+U4x2wsm5voyW8LdK+5aUqPgh90KApW7fpt07FFqs7ugsgc+fPK46PsIa10/GPHfYfGWwSjN4t
/06eXzcdGefKjG7mOA4/TsYPCgtuWxDj4+NG+53o17flkIlA6272N110GCNHbSmxRLfU/syJPrk8
lrdnA1OeU/9uUBlK+MZNsg6ppEo+gF5lBKuEzEWBMAy0uS+GPRtIqrE0lDGcl+ObUb7RlR+ZNxJ5
YkGBJdu+HBAV6kH4f9kCf7cfDnF6qfEyXUCie3iCA5RFXyUFET0nPS57QlHO0dKyt9W8k9QC5mgn
jKJQD/50c9KecPIKLCZMHTUqgM2xzRW52YmBe5bT2uUb3m44Ff5f8EHLNmcejAiT+0ZsmYeqi8gC
2t1zH1TiqCOIGeb9vFE99I5Ag74NHqetfEhgPCRLPrCWDxLEQtGYU4IgQqIVw4v5Jh5R7NT23L+h
trDUlg/bBmS/h8040YE7L3rgvGn4j4CyFGiQNnqt+Uxh6nO8vhuOT/kq2tHmQNtPW+3NHhCtqtFw
zbPr/4ukurkWTmv0HJ7fT1ybVQiVHwA+uH7/lPkfFPAILkPAjGxC39JOnOgCmydh8r2B4w5as3TA
01cGOzme+TTvp4DaXYeTKLDVTQC/qR4fXEQVjQxEfhNvoFE3Drq08D00eWXviVK3WPX+U3DGrvv0
8+wl6JuqBmNlbiu/S8OPyb3R3Qvam9uR9gY8sonMA16Rr/ryvrv3OeeElzXqNg9hT6O/vBQjXV+z
XoGh3umiGqR3FbbCPO93XdL+pTBC7vT56+J+Ef6qsI7kl07Sre0Fi5SyTJi38q2v+tn0Xdd3iLzM
xG3O75MlS0sV2sbEWc+ZlMTyipZxrENCO2N9IlGBeQMlcQAym56wIvx32cSn5fRoOpyL4Usa9tKU
fiB06Bc9dR/mQdS883gbVPd/lbyCBeoYtPtv1S575G0RPdLefRTri+b+BhKzWjbCgfWqd7dpWVrj
4O/BsYttVcmfsTToi7JYhX1xPVglWwpPEscpFWXSCtOcKTfFC73HNWHIrZPwkaFk2PUpaVZ//6ul
M5A69/BFgKJyR2OLKydwoPZYOgEQTnu/rgxaTPqCBIdFtGeoe5ZEvYTosY7Km/2uJuLvx7x02s9g
iAoOD1UoNJ/5933j93Ts5BUGroTaoydzwFVYDts9CHF0ayGu2P8qnBeMsMHTJyKfrTQyMAbZr/0l
ONU0hBYUzxI1wm9oGGv1AmzJUiGfm/GnoIUtUFmVQn1HiUHLnROyyVgH8TBEpMbIDoHooSYKFUdN
3uUHPWbpbgUlGmgd0NMOGLoFyCqdvSwCqEuWJx5WACMqE06rLo/OVMzt1ApVVA0YoMQhc9s1X2o3
UheaDhvNKH3MrPUwcv58NGjZnOwgyQBTmdphSFIQuAnHNyrC6m+8Tln48gZaM1vQrTC19kv+jUON
UPYnpSDDbh9FJawgGpviY9r5xsrRKkl2SAUfxdBcHrYS+nIkDfY/f6EcrTzEf7GTd39RvY1+dmfJ
6n3FMLHTD9CdhQ1KtxQ+WmtL0pFh3dRzGMBUcRCmCcMQAGdhXQMUPwbPq94Ni7RZWkvg52SL0z8y
9N3IleJpUZktFV0COVTjmg9DdCWG9rBppxhOVQ+B1T/UfeEnDc6TkqZbG7t25RIoGOYEvV5Ts8S7
bemlH5SmyAcApMet4TWfLjdbY6TytNMx/Pv3+OYRX9jAb7feiKLjC218SdqDEqVjeRY7IwUppPAu
Q6BIBShRpUSkMLmvQuMc1DN7F2JCsTh/k76avEZekLHrcTzeBfeKfFNQtixU308b7UftTE9FPzUu
bAnVu9doyGeSL5iZUcFzjwGW7UHJmeFP18QPn5136ZdJNGAkQqL+Rsd34NWFY8TyJuvcZwtvAPnS
HMYemrV23sx2QhtANSYn1LQKxkEmHZ/36ZmQpRdpaDr5Yk/C1PbvsWquFtigUHg66QMhOXtK9UYI
pKm6qehwh+0oui2jH7YMVFor/vj/RxPrpM7/ZwsKOQneYdTdBxaariFNzMcnMSBbtf54nszy4m47
JEV3bmU3onBmW4nD+uAjkqmf0HzygDijMMa4HzhLdUQGTqZDFthECFk/bdgEmZkxxnnFEeUCYz80
JMTzVUI9IgPyNsuivLeNqxHa3uQweeaAG4IqBkPGwVbuss3JzRZNhKgKup4aE8VCZw4T9BkfWIWr
tG8AkfODVQOx8x+cAkXh+sqruGfVCXxytNFIWKGRLUB/UR4a/JiHFgy5l7P8DX0BFvoGT2vtd2Ij
uM1YfdboumvhbRyt3xSYvywZ59fCsBKRFxy2d2arJKe8iTSg8usGUEeldAnCkfZutjLnAfzyr9xT
WtiSniiLfwNqj0o+ILKAe57ygdmwP2NqouzxqBGWVhm1rq4wUY7/8vt6Dg9YzaIwu3VQar4JbCBg
VAM96dLuE9EGrRNAx4//+f2KZnhyjSXA1wFNnHNPAMdwdQ/DQcagTBhGavnyBPNmL6ZfvCe7ieXq
zoH9N6EUrKOHA6NxHzvgCPeBSScD7HSfoRPluHo3HxIRwg04O+rZ4suuwS0hVToucbd9SVi1QP6h
HOAq//WzuWcYGNOspcpj8GtVqdxQn4h8ziUvExq/3rzC1196Jn2RUjg2/1yyFbs8LtxXRTBmOl8R
i5UwYfFFXVGht0VY2PZPjYSpbRn91/0oX36tbqqTZtov6tZn/9m7g2gRPmOKBzluE1sAEv3+DRX3
dxZBImnNYakK4cgOqxvVTlJKbCxc8G0F1QFrK2jrqJPBaMvpIoJbgEqAiZoSDGw0AKibfbOMh1zL
2+lQqn6e70ZWENVV2hhf2oGs5tuwIsK9abvXhmNKSkKy7XVplyG+P+Ig6+EbqX/9THsSi5BkvKAB
zFMwc9BdfKVY2xkNbEv9isYW+w09gI+2FPVeCO0ILdABvK2BADK1vuJDKhE8ATLjMVWVrnDzeovt
YWiqMFwaAvFHNfMWc6+1BMSyc1nhdVBROGpL+f1/Vy2S6lp0JH0Um+mjxm34bV8y9XyfR4C6NVvL
zeYxAoAdReYgxHRTM56asUy8QAKZWA/Tp6DtkuPWYDp7f/Gy4HAIc+PHl5PE3GeM3HEZV5gGpi4Y
L0xzzUzLD8QK7m4QHTc7rmrRVld8TsO5nrE4wWJV+poz8qDbZdaUZIk/07JqyUcXMBHtiz1ieL6K
o5aGstj6iZ1vTcg/8Cjur98q1naiVZ9+HFnoPrboXHb9MUqAuqBOFf+N0oOApjjF1DUyh/Ci4DRG
dqkPXej/oj7DkVfqm14MM4IA12ThJ7mRrwF/hMec9kgsindA1dLz1dPpQ6krbXs87VL8en16YiSu
f7vwot+f92VlR+aS/7pY1dPqr/DbomQxBZ0V0iAETGoJJ2ejlkXM4a6pPH8neNS8uIhjuDB6E7sQ
4FFcug1Obv2UAUmAzXs2yjHm9kM0GrfPEauu4pqIBq3CABsE5UfBxN1yeqMDJmVt6ph9j+FLxPIu
dV5AM4s4LdjPyK3td3ziIjvgJQ6TbUTAz1w1rL/gSiLPiMLP1vBiufoIdjXqjPj9B8timca1+P7z
Ze+dVEndOsKFYLPsbWy1R0n2QDJ9IEZWjcsZy0mWzfSKAFJsM+9dMIXGS5LfQqmBGwsNdatWHgei
3peePZSvsvoMXcPURAyE5YmAc0XBNWcwFm7Wn+2Fn7Q0ltoCA5dO3/fjjLOoD9X08J5fzYI6eV2B
zW+GDgEkGkOHY1vKSq7S273Fv/HbKEqqmyV0L5Xf00zVyLwdPUxOZhI1pllXZAseHsrDkgnNJctw
0t/HKhe2sxNw3nTMfdqKywM2XgLzn30+GbO2EU17jeydT2tw4XXIEvMDDAsaebBDrjjXiYKeWgHK
rn31l4ARFJl+sbjJGqvlfiAJ87pimFpmFZUWNAyz75iPzKHALloirsi4d9pvKL1jAkIacm+K4GKp
QjEdm9k53ffeMLFHZFLrKQIZRkfbWPI9s1OMHV7ENxfFJrDVAvrlGEtlg3VGqQI+LdHJArJzivBM
JLNarHK4pRQ9pJZtNMvT9U7/ve/mmanG62dxVkWvVbTjiNV6Ujvj6z1/FAvYYNVnaJElOTLP6SrD
0MigiJPW1uh3p2Xc/ziLk9mwxLyEUn4tLD4vJW5rKsoZRar1496XA3Xzqrif19qKd433uNEvnNZl
MhGXkwgas+1uJaiW7jE97lkle/YEzuSAuRU/Th8sbusVy8nz0rKEqR1g0IGh9wduJdxKgDgYJ9zP
aHluL9SP5j/GSiMA3GkQVixT0wU8wfC2OX9IaBo00GG9gERcEgm2Ly0jbn1PLdGz+BQ/tv3M3FeH
+iRykir0xdmH8nQnAIIX0okOpiwJOT0Ims+o+vPVjrOXdSG+Pb5UlLuch6hLPppR1aIAztzRZLMy
lXkiCgxRa591CgXyUVlPyUDaY/a2xmnNWhG9yGGsmeLejnTHy8p9SbDQ0j40KCvk7PGdP0yZN+TP
rIIHliHlVlPi3kuQOryVTtHy6jGjMLEpcJDb5z0+v5etB9izJ2u2Jm2T1H/VireeXKvX/Nsh+KZc
x3Pja8oiDsaMogtmammTNbwrNcoDHrumJFVujPQPQFxr45y6+bFWdaX3n8NYABtWt6b6ArO+euCO
xrSynLAr0cYwqjaWYYxcrIrv+2QXpYV6cLYTWWB/zDQCxLc0oTVA050npoiebGviwhCn74IsnnIU
KKb+M8pdBJrSZIyr8+CAakLQV9y7gGsS92dTsZgqGGM/NGeLz2nB4SQPdroXedEgEp8/LwaeoIvo
0esYr8X73VGho/XRsGsalSj/KgcHmzfPXsXDyH9vHOvuEsQKjtIu8gJFMBKVQAQxn/IR2KPStvX+
6m/00PX3WpqpTJZio/gC/VILErOKkRQC8TOwVf3KSBMompUWni/wVyCiILR++yNYfuM8JqGnCc2E
bGbnpnm1/rquMTDnsACpsjL9PODOOy6af78ponaZaSyFdCNvVgg+dwcR+M62XTTTBmLcSMaetnDA
SRmkxm2WN87K+/DoMN0L/+EMpXaf0gN2BlXa4a+seB5OtyykPJkZFy5DMEYWn9dnUyB5MWdkwkVt
uG+KU7JxybqM1tv+jatJnpzhBB9BIPaOm7grfim02p3qfnR6t6AbeAgN8hOa0aNbxI/PxMR2yKHY
OpPcHdmgWI07kJ2qcVoK+4oR/j9SVRYtnnm5SkztywlhKWHg2zt4u7lNKhiyhO6DwHEMv/ddvIkM
5fpoVJHu+XMe1hPYZJ5CjL1s893ozEIYwuBefodlzJLchyytUZaiauzUh2bXYbvqzCO3oFUkh1jx
2j5++d3wG4qTPbPQ0BoU5tqexypjhXnfOy07HJhdXPpp5Ta2gEAjnz5ehqyDuCiCFn7rTmqDeiN2
kScb1426gpSFdoqN45AlV2TDqfXG16uAiQdTuK8g739j15S1WKCFsSCYTpfzjWVfE5Xv4b8OlaHY
6OXTG7Hkibwamvhq0A/oiCHxaY14UggcbvuINWo5c8xMTDo/h99Y/qpCcN9AHXYkuA/CkE7XNJtp
T+c/HmOP3e3w3uWompApb/hL7zBE3DKvizNd40pVayupxV+0O2/zKNQXQfHzORPV2QqiJRmlsAZa
BV/FLM3x06aXhpjOgr1c1WJbiQfY9IscOVfnOe+roKt1T+KF242JphPhzDfiBgtlOgsFRUp/m/Uh
K9JwL1AD87IPGCBdlk2Zx+sX90Amzbbn+4MlLCzW0QkCem/kHe1JwHbA5h6q3vK9sQyKFFfRm0eE
Bb99CkBMyxXEkgMK0JaCYIUkzH+0AonIllGmeSbH3DilLWC9mgyHWDib2Puyx8OMj7sf6jK7U18o
Rw1ikgetkG8pHis/N2pPYk/Em4wS7J4VFL1iwTfd0btY/qTEZJR7u//2c/9Jq0fU8W2pu5sD861e
5iEqAZPOqSXKHxPjfjQOW+DHihQIl4yddBg8EYT1yDTa00DAF7Jfja8CGorPWHUEZTDzuwCFDKwK
ek8R1lAywm7vn4y3rEF7oniKG3kwS+CD3sTdpcnjFtK7t2sReUK7KdJldcjAPdAJwur554wrhDNK
4BF1XnupYr5CPofdcj/Fj7zn1sF8Pag1xem56MYrPRd8skeVyplqnCtkA23xscGUC1VOXHO93IrO
vW+tvaQfodhm2y/6rzOmdfDUAYXxkjjyHEQt19tyfXTuuH3nellpXc+znbgnoVZDV4c6xxZVwuvx
JL1O85BamHmwOyoFaNQHWbgsSiSB2z/sCzdH4i3qULHmSHEOo6hVbmZTfNBkr38lLDyQlT8enL36
aEcll6iNXMJxiQLZI78Vh9fWT9vuJj9vmg0tjF1Udcl2qPO6Tbfg8lP8VtDK7IQZzTgOpS3AyCcY
BxAozK4inLS3pKNw/FMyDWf7LYiQZUp49cLP/1VPMyNERbMRCKyiMXMJTJG+gjDxI03l6c248OHh
JmPj1wVyTD/25T1vcpTsdYINlqT+SNPCQdyQRKhcvXcuvsXAL1UTarxg0UxqQ0FEntZ/4whWyzqG
QqaHt0qAbNG8bQ2V3+6HOvoJW2NrrZoQonLRvuzn4uarSbnHfci3jn4Iy+vWvGxEJeGOxcD+rwIk
+MqmRG16GNfBzkVP8/ulW95xPNvXm3xgyzX6lFvF5aPHGtA84se5ryu4edNxrEKmW6JS3lpTnY9f
8KWJ+RXUjlq25C6vp1u2nueNinRTCDEdbK4BRUJx0XCn0LNpB9Ghb+gjxLDRBeMglVB9eIXmG7EM
WoCqE+3BHjFa8lMg44fDzHRyYKw7qFoCYfL02XRiViZWbiNY7A76Zn/hnSA6za7s/IZOTrOlEG35
c4lSuoYjZHq2630/NHLwD/A7Og73xuleStI2FPS5gpjUBwzXwjwGKrQ1WGy0rceVaOyCqruAKMCY
wL2LFtvTB1PCa7l1MTIHUSwbDUaQwscxvXm71IoiMJaAjlCgNK9IYkr63TnjzE8XCRSSd9c3JErD
PJYIo7UywTzjU0LSzyP9+X6t/Nwt4s3sVtKyUh3eLTsj7zFCj1nmAzUyuTiB1eT51amr00a3Z4qb
aB5hFqC5OgOXAavkiLPcmyYijK7RECcqCTWYqTxOFVH92lWYd09nI5yxAUmdg4sDSBtiL1+2dlNT
vb6KdIOT+6T3HtDngonYmZcWfMAI6YoTOjO65Y2nGsIIVt9nr2ipITQD/7Ogeqkl2gVEb1/YkjcE
spw0xTbForkfNX7YDb/81ZxcQ+PxN6Vh5AUl/qtdfDPuMco23dYjjzBD+RyCcin8C7QOplnJhvQJ
JQ7eukNeYJ85vVgpLgeKfDp/+jvkh+tVYz4d3s1KFDLm8e30aOGaZG2ZWjUuMrUuN9j/aUx8fial
FHu0swwdWqxqhqlANJgcqH8yLNEbD09hX3niMTcoiYEw2UI3UO3K6kdCvixm2RuIOirwhT3DdfhB
SI7dpv8QzsIQ9imdYQyrBKUYgCpMdexCNepZf398Lz0wqe/n+vdwIITsf0OTv/lxQIj7Qx8T200+
OslUqnCJOQ4XHo+ic0Rpu24N/RFzhJEQ4D48l9Zcfi2niRUfxnQhCLvTO/DEddW3z4UAa4QhAt76
LDJt2wBCs/UNSHcZqBsf/2NdNeZICEMqspWHpoNRGOTZihKLbf2tGVJWPvZ/UUpptZTW6bnUswpM
GrhipgckQ6DIfmaYhSjLHVjh8Bg9gdS0/vrxGlBfJOD5f3dch0s//FQoczDLWEXJuE8wcfAW0kB8
wSfYjMk2HXGf7M3qZDY/jlRRgquz6stEKeFfGn3pRsE6Rml1mXsiLO8WiDpECYRkVQzxhhKc4QLq
zjwIppix99pkQrHx1xUCVrqnn0gjK+P7CLjD6sxFlQhHf58oEmcstBHr92Dn7MR/YyA4507KtUc9
tLVQgXsDbMuyOIXGMc+FirbtrHtjgpA842lNPIXN+abHkh3Ut9ltvNovPYobo7XjQhdEOQZW1RV8
Vdly1FS75BlyOo8eq+rt6WVchHAlCdiwmgSOCy9FQIgxSmPKTknb5TVp5iOQ9OF8u3rMXk0y+4ef
aiuqvRB4fU6PDfsOzmi2oc3bY4K6sSn/lfNM+6b+AnLfDdxJmITF2V/Gtkun7CfaKy4rhBJM9Ffg
6EBrXhRaJ1e1WXzLDjTosvsKOHcwD0RcjCL2Tt+yMftlZrvdyYUVxni5P3/HNJLvhk7oy3xmYHmp
BNIKpGbivPO4CU0Y9bw0LXlayeyHZTcE/2JmLpK13I9BTZFDfXeRbJpCklRqeRZd2SiLmkzvD5Lf
9h9+b75Gd/1Udp2rQl16x348qla2B5LsjboTqKcoWFWyvbLlg7mmxaJ/TBF9RJ3sDtjO2yPEYXZ2
Ufrv15mi2qfndpWMJMJ04yJQ1Vd/UUNAuqV8Wrf39zjc8Ft6u2Wk+l2K6B2b7Hz3jLk8XMK2wUxT
QXV3f47GBIzrHQIMzkHyETegd8XX6+3VPmlk6rYIxNOUgPvLYAeGMzT2BbiXJiWpC50062PDBnkX
UUSy+HBSfNBZGEyktpd9zZumChrw7HavuXBu1LHLw123atpKM2McmtzOc7Edtbmsk5UMl88G0x2i
jRy0cPON4IL/dIdyrEI85vx/G/Fa8lJ0pb8DzGEJ2EpsUTXhowhaiY9IA7SRCYmCJOl1I/HyDULi
bb9482e3c8Tep7mMlurGR8KyU9rSUCAiyeOnqLyu8tMe5QogSzXl21yTSN9A1rmJl3ceXa4419pd
cGJgFs+slHqzvZ57rZlD9mI5lSBLeJosKUip9F+DUhomSi1+kHJsq9ePdZCc7GV/yiuAwphGwR0H
xwnrc2kZuJutLs1h+5TJ2andiLvaGNkBqYrlN48zErHk2EjRt1RzjcWQ5vUD8GoC1eoYxHfdenC+
lmxteY1B54CCjOOU/8NQujs0ArRFfI3hll7AuUcWGzzG2rL8PqyyweiAmxwJOgCmTUUhq83+oo+H
7T5Bk8LLs2YY4MbtmYSdPCrw7gqVjslv2q6nVkxOqfCDNG9N/ZFYV3BDx2ZlqtxqYUcEeO3FDfKd
kaamsthHskIyBedb+JE6w6kN03m1/F/ZIQxMEU64GkxsuJ2cIOXu/PQgHYJYcdiLayJumPXkcx3j
2Jw8enlxJ9+CW2h11N3bzmDRxwa5suY0vGtvyq7jlXj+6VlkrOHpbsr/qszNyHAS9cwkUQNGjMbD
ukJyJcXwE4jDHsnzVdN0VQZY1Vf8CqXuMucshV9xFTtvSwR+8vZimrVrTWutgsUCHzmGPO0hBy/i
byqZWOVH0TwElC7wKSixOMgQRquyn7hex6qo+eWQczdSO8onrL3HrO//BT1DRdxAlQrN+zTh3u4D
2gPdX/t4jtEiQEPP5q2vNmUdTf9AzDVbAkHAsA5Js7t9qe/BT8tk6Rp99zA8A9bJcGpvfIHDuak+
n4U/56EBZrIoFj2JhfMKmjATj76ncOynuPLVDLK/Xku0D6mY5Z3MpursVgdHntXYQNeaSQ13WmlR
pXdTKCYR+t8Y0NMm9YWUyH/8u1QryCWPkWZ61Yb9RkiWC2Qe/QAU0p5WNLD2vtCMHKl71h7Ihzrc
uSvJ/vXXQhoSDSJYNmjlvxRIHmbNuvgaRh44pCKrY/4QNg47hzf5hadoJ/hAiAPE7J7OiAIP2BhJ
t6bCxPwWQYGw7+A0vuBx5pzCJOzNkCs+tNZbrJ7ODHifH8/ugKI985h51qL5UlHDtHh5Quhp2Z1c
ykPzG5ngI9Z5a93VI+j/N/FzMqEeibWz40091KzGbX5TQqD4cXawhhyc6xp26IfXF1K8a/kSdh+I
lXwq4IPLPg79NDKJCV1IiDRwHKI+MD+6FJqpygHV8h9mc/1c3XsvS5OE4P7/dge+IpIRhLrHuAlY
2kcV0FIKE+S70DMtmq2WmWs8CphGHSJ3Gs6ldQ8De9k83WY6D1jrVsnUMDqfuyFtKS9PsSWXDVP9
zV/xdX1OpJWyDVVYOkAYMpik5ump+AUEQ9fT2NWnDFyyTg0DtUBhMDm88MtfJRaNPTqH9dupNZMK
9GK1OCVtwV6Cerpe8FKjWQqpgMaIZEKPNDujjzRz3PTk/EivyPSxAc47xa+Z6y2ulEXyWt5pM86h
c4nHezX7FKYhGAHFGg2pHa8w8YJhnL00M9tO3poZuQjkND5s/q4T2ScXyEYRDEWh+0LdB+ZLbxuj
v4h2ju0vckfzcz+kMfKZ8zT3CKES5YyeMtdqkNTokyWZruYlJIQ7nBSpMvv11VrbxmO3lfGqs7RW
qUBMSkff4i/3Btaa0rRxaOJWVI9rbkQDFhflyIyas8c3aT27UkF7uxoNeHuDJrTZG8hZOYu+P5sN
aktwn7eViDwWnqFNQzO+8wBKb1Vnba4AcmVnGh7IP3b1gzH2XfglNJDqjtZY+q6zKfJbHaaUSH6K
XZy/lTdxUkL/Wkn+l8yg2JbRiPl1N0E8Y7bjfEjaFg2XCemv4DY96FaxAmL5gHSgGRXJIqBQlLWI
u0OTZyIzRi/2DjH9U6fNAKnMuIL//rcJcDhQ3xpXqmQT5jYdk23KhcgWV99R3blc3wXcGSENt76M
frNKyjAXFSUgeLajUPDPj5SMM3hi2/vwh6C20QHjrNlvhVz6TGgqKthsyIB/FKujbviI+ByVNEH+
VYHABcjT/tvy6aV4Fa3Q5WCjq2sfkljGpVR67VOzSVBBtE3Nevu0Kaa3Y8d6tkPn8K96QUKDLHVe
usAfMgPg6WLi6pS6DzjCr8zkatAnHFV4ujXQnEv9L+r0EyyUbPoGW4scTaJJzsNjPQLwHc9A2BYs
DxNdgnspEc6PtCQcQiDjfzFv24cuMYjHH+tvsRvJf9aN55NvY8RMbWTjh5fuVvmwUtz1S++dhVrB
DQz5XsFv7Vvm7AqWLHBXyVwSfDe64df92oQPotaGKxbZctHkadWlsjNbkBA0EYrikiXttpUsAmLo
BiEjfaaG4mBxtUXPm19jBlhTLcpWzykrDpA6TYnGghIo1CUjaezytIr1EtaaC84IM/MOhIVHzl96
zqra+2kuN/MV0c19AZd3lSkrCHxtrV7XlD8LOHL/sH+/K/0XxEEpxNzqFlLNJV8VBe91fs1GytHw
Vsk4KCtQdX+UkkXBq0AF7Xl6ZS+tLpvoOPIfGmjhPV4GyoKGOTOStg7Z4mNypp3ndj1P7F6qwWW/
SaVLhdB4p+GokWUq85qRSPBvlPujZi+Gm1WSVhwqzIVVgmz+TMgv4w/3rCCO10orR6Y3uwydNk1f
aVELDZQ1P5Z4Zx9L1OH2O0JuuOa9Xsvz9n/P7vzqpVpOxy18x0aQf3mL8ZZykIagUSsaE0tdOhPq
s4LYn1jUoK3oD7e5X5pjE60kn0O8/ulwlqMu4gNaUv1QsPjL9mpCaCw3eb8sb6OQwdX9DtJbTXR9
66y6JaGfFTVlNkHYvYuifFk4mYhOJLpnht3ehcTZV47a+azq3gb7/4rcEdfA09UrbuorXSUasf4x
eZiL4Hb0dapAnkyLI1oJk+zBWTvURtNpHru90ZtgWSXMYLbvmPJcjBfVz4TDyS9luZoIJbKUOsg/
y7mwpHU3WWzVvNPx3NXCMcM2aySCZYk2BkvUDHSiNrx6QRot37R45trlIy5cp6H4tDz/BgpQFHOW
1FJLeF/yoQJglvg4GvaJMz2u7xt95b3MNYNEfs22J3SXhvbZWS55CjwvneEO5bwPoaf79VZ6tD5k
4+WQJ9OBeQUA2CwTFK7lyzoN3dEg5vJ1CZaQI5jNKK1J/VtnRNqmvW+sdivBxRPWqMK4UIWVKqTe
0muHxqfRBspfMLbsaTiQ73GhoFXzwOTRzsHefHfBoGKRgkb/NiVuJVe/albKFES80OeFOZO7Rwam
LF+xxhQ4ijj2BrmFHQzi4uf20DgX+MmnN2P1srbbUh8ep3A97VtyGYEnGimld3NMavcNfQ1hMMtm
HKIr8uF0dnFTcx71Lpf4n1bdAR1Xaa/PdQV0Ixosv5tID2zLeACjNJeMUKwEUTVMxo1vgj1MxgUB
hz1RYfVjbeAElPrXQDspMzviTEsGGktMW2ds6EdRr5xhVtGeJ45uohcwrToVDcWQser7hhNlAgd1
D7uRW4QKPo4G+kLxAccq9sAPk7dGJHdG4v4kDOHP42bENbA/EmxDsOSJfLVet95YrxYTApFVx1ib
FmKYdyMxRITtciq132CHc7N4CYNLk0GR5JaNDgril6oMX5naYpkoVOwnmZ7eTwazcVsB4Jdu5bnE
HZgQ09SjxBMKNtULhjWFvI6+rAF2OZDJgokNWczaoGAutM2bptXfxjfgsLQ+zZNE10yRBKHAVpVL
rl/AuSFvX39w93B8F3PtdJPWFIJlH117GgJ446jc3HV7YNAFiC3g0sYIszEDFK9xyjPa/mkT9t60
gnFAi4J5gb4KlgXFQoL3DloCUNFwxKcf44KATtzexgN2fgHezlIc0ZoR/YZvWyQq82SPtbBQ0dXh
eLvbMcnFi4hHICyVBwNs6xytKfUXpsXeLJv0sThULfLAz25cV9MXVWyzIYta04Gk75e3KviMjegk
TBqC4mqROFjxb3BEWTm5PshYXe6SYGGIvCNmvL2tMwikjsxCe8qw7kf16RhKxp69n8MIEsAfcoJ9
DPk5isRu1j2hvx8l3ZNa/TmLhSDwRoKiy4fa0StFK10/h/Buba9Frp/+AYtKxvosTxEviiH/6M5+
qYgCyCFl0JVLvtjEJzytpdA8S5KrMyciDbwtNNZ69vqF3dlbL9C9mYZ6EQ5Iwb2DPuOrWZeKR9PF
rKMABOsJJC/ImT/soGG4ZxRrB0MraqsGTphcnAcLlwm+drlqxgQvYK1vtJp5pBA22XDwrf8ffOz8
l1o2XmiTPPpU6GVGDXgfKj6y4+4Hj0fEMt9rV/H4O2nHBldHJ5eqe9+R4KZJMzgO231pnFAYWQe4
kgZhTnK7eBfO0xFdYAssB3+PU+1MTOvaU5ehySVk/FvqSHoXI3uoxM071P+ohOBBodDt0f5YMPR9
kPm7NN1XFRJD3Z5TIcC4G8L2hFvEH6k19urlcARy0PXlZeGlmN3Hfm60I0qEoMsvJgIUeRUguwam
pnaIqJO23iXbt177EwPq4pCUTSJkSMmAQDCcJlXnwqg7nVaz8d/kebxaRET9eB/99Crl72A4sprc
f+R43Pu5eXaiDHwV3afm7/YoJWRbUAlfSyJPr3YE2W7X1eHtG9KWOwxa2fYAg+ASuTud4rWGTEt6
5Of2U8gcTkziGCfFnbNYe4Mkium4sUKzI4lgfv2CN7RgXgdxUkDrEVzf72P1ehtai1jDFuI8jOW9
FZPTGN8g28Vc7lpqCTMCutv/3mkABRfqRGeJKvtMOBSmGhOBgDqo6KIQ/1Tpc5ih4ntHZKj+b3nq
OMinEim8Go9DRMHufQTJtFR3iRz0NuVZ5GGe3XrHf5cqdHVhipALAHrYdKjMy9mV+kvg+q+l6N3l
CYwyUJ/WvO1S0ggJ6WY6UQJP2C6GMRgy7nd9ctgAAR/NloiN9XI1xOWy0rmja/3UO54GWbWNrQGf
t1aLmc/UhoRxaTuU3Jf+ZipESl4j5tg9oJg3j9loKXpbYfyonGFYgvOjun3HEOqbK7aI4VjZ+BgS
ZH2NuWWafMsbDinhYFW5jzCQd6c5L3pk2DdKsFpanEUEuNUmkew1qf8t8JGUp9Bdwmm+mmBuz65l
bWf+lDu3dmmcMmzORiKg65L2HY3A2aP5cNxHjqk9B/cOJR7QXBeahImbgARGbLn14MPZjNfIrBQE
/m6jhmR66aKhYtQKkAEdzIe7y8Y6bb8mAjAtSDQVp+5D1303iScOmCgirLO9rpqcY1287LmFSM7Y
0kkCxoqy7W+x7zjFCduv6eHdazsInEOqyfReUk6RlGn9GQzGOwm7cFVnW9V/9QYR2vOJvrZL9KyC
TipnQXLO1GA2+nH7Iomr9cwJal/37bC04fFwZHNoVdFl3fS1+vmf6VuaG2R+L2rSs6fv2N3oO9rh
zdLNA8zFHv3ZA2GRpCZiUp7nPs8cM61SytbQpMv2CYS8pDTjiztTj6RDRxL2AVcfgzvoL6/+Zd5k
CYMyxWW4SqiFcZTW4kJiZyQCKOwJs4L+vYSMFeEbii0QyC715LCFLIucj7/wW8Mx230InRXjmiV0
g255sR3PpxrEIJVjFxjD9DPE3ltPv0IEW5qRGqZARl6uF/3zaveeNJurl/RQOtcEE8roXl9QeGeq
d3P+9VxtEQGss+ud6RTrSFj4M5lZ53Ju+4NoxNudaVX919MgZENKv2L/F2QU4vSAklDD2no1zRgc
IumIzxRSFxSREj+4frv2uzlFJ4Cf7chUwDFG7BRicyXdAbjp3NaIzoToQAZHUZDna1fbVfNSBVQg
bfHkuoG69zW9jyPNEPiAGYv8z6TjNci9R52LsITtllgO8w2dXaNv+UH5hxBnbIUpK/T0k+5pOH6I
jrkBHDcm0KajGtbyKT+Hj81aSsFrh251iibiQldSHQW53t7G30j+xTCBUJ8HiX2MHTCUNZLx0fFx
79MUeIPwYwQUP5+oSi2jYb9D1cteysrHWysGN596yQHIbq05PGGSMW882ppkJnxsipUpi1P7NFBB
kovgp+ub5r6SW0ILS24LAXwhtK6XdQtJucvnftGLqBkwWhj1et6UUKTAB/FUEFgesIQ9vJbTnict
jvfpfc2ulzSAVZoe7BTRUKL91GiNEpPRH/w/twE7LWogScaxy+5iv07ixkjzd91Y6E2aZ10RGZYp
5mBDrqJYtKwOylWM5i6eoo9SXYGOOFq4zmIhDkHxY9aCtkp493IdZsUI0UiAg8luSYoOpnNxrIzK
CDIr97ptyk9XSdtmZSiZizTybpIFW6M7EFSmxthUgX5zu668HJQcdmht0Gj9/1lTF3mMCtyvyrMU
gKEHwmU7nzscY1RBfr2MicGKF5k/K89B0I/7SljWQtZuhzuXtwIkVE7IbvJfXvTTpMowXmCTSAvx
j/DmsCTHU/vEAQndaHmPC23PwCdjgame35sVbWlCPbmFFS9zXouYGqTzsisg8jAnwiFii8b53NeR
ekq2mfmYA1pG538eQ/NVfoTYIvqtuQSv5WRxUxf450jstSDyXfnRtxPMk2Sgqcd+nGq+6GGwW4p5
DCiqQBTeRMs8JlMeN+dI+bQYAhiZtkk6iparh03qbQN0KacXgij09e1itH081tNPm1pDv+vxcSfH
4P8Rr+xiL049pKbi07Zbu5CO5JLyZ7DgexqCfaDovjgA1Pue5U2LuSChY3aeFh3mHg3bVmQbb2Gx
1Jo2dBus/36wpl64a0JBrtzLqUlpM10NkcwSHypgvR6/KP4WzmJjifhrq/HeDgBZtTTOrq1B5z9o
i0S9vvbivTgrSqNHCid7t8vpo4hJ6bORPSjTjVeuc4UKFOpyf79Ix77xZ2o63IC9FXKovOXMzd0n
OglkLf/2N8tACeMiKwwxhoRT/+5tLJZ3iluJ77dfDUjgsDjHBjCoqr9c7mIk861XlS5hA0rUrGQK
c/KrUaFgY05W5mjURkJa8TtUBXgq8BLeqgWVaHFpOzA1Vdx1wRc6y6a03nzOFiASe3XJdEorSBeB
QVmnpK9dVEW0bFwLWomifPwD+KhGT4SUFdjCQl7haePUnc+ppYU2xCorHufbRTLnko2fJBpCnJ2/
dkoyTylPIo/7aVLMQAaQU3VzdDcUrYZ0ZuHxn8OluVwix+9/12v9F3X7QieXBuYJPK09FHQgl1O9
leTRdQb3HyoAzUEb7eh5smVlp7RHogz71oNIn0+vQK1rS8qvp9S7qCSpDDM3+jB35nLlA2tnyGe9
CcwJIq+wRKxSRI1ZaWcHJYG6NhDbm2vQ2Whk508LL/7U8hPJUi8SAcNgBhdLUKv7v9fSTx7EdYih
nkPulDsIdVbo6f2fIHSUImwNZWZQkWew2LXXstvawLSPL4yBFbldzjM75Oukq4LsI/7TDyg6Oenh
k0xXaKRXO794bF6qUXqw7PgtDaGvN6sNZ2lqxDRynwOXRmfIYeV0sVYnaKPyhHBrMiWxKiMbE4Bx
ggTwaU8diBiVcYQvk3FhiRRUSW/VJCnsn/RpdOEICqZpmok2lQet05NjhMW/8mfmqvZepWJoB6g7
/uhVxMBiC1X833F2sFcFOi9TasKW7PzipF/RC/PU+Qz4XMuQ2Zjsg39WurZSiwFgHhLJ/BQMYwSK
cffWg4JpCltbyFBazY/rqw8fUlt6A3h1dZRlvjFK0I/tk0+33Y0fHtHqecm+5SXY2pRo2TBoQMy9
zVJQWaaPCbAOZw4Y03uPxmA4KIhpeukyAhREsVbW4OX1LGRYZEimSiR711QiiReDqN3SdkZDJa7Z
6P1mX+x1BTC3d7ZD7eZ5lUmFvlFhYzvhrNhqlVyvNNW1vzZoVtZ5anyn2B7KD82t/fzyVNJB3p2N
T5Uj5kAMfqOWpXeRicJCAas8JAN0APZsaP1XQ9K/tE7V02GR43BB3uu0sRUXD81Cb+0p4CxBxEou
NPxucKt+PpwW6Mv06LTo0B9sb/pjx+BQx1gZ4x75hfXWhE6D73SLEMFV/IGw2a9dMfXEAooZdJfh
NN7lOoAujEM4SS23LJwT1Ait3kNgmBhr6A8LYsLsujBvi8zfzPx7F4AGaDj+IETm6JV9yevcT9Sy
th4v4N/LZPDYm/xxiS13lPYKDh8M0xb47hX3ww86wXvOx55G0WKyDS4ptgd78AMrIVCU8E6Z9v59
zkShX0BI8Io4lYaHX6mdEPuadvF8S9+4zRsWugF45zqHWM9p1Bk8+f1cn9bObavCvEDVLrlHiP9A
Mnow8nPNdpuTneMZ5TK0q38daaSgmHWiqucfDYnRHBE1vIlyGMHZ6V3Vnt3LXPzBm4tIoWKldg14
YwZDW+PM9cykCsi5nC5qYAUxzICcZLz4C3deRqc4ilYl70qlVqegPIfaDkz0H7KVX1ozvoolMrz6
dO2igr4sdL0LEDGZEksqKhrKsr5+pVjMoXWD8vau42//HJoY5mFcnNFm46d1bph5paYReGEXCsU5
CRhckI0NDuYdp1SBRuKZtFS/cuTTroXpyNoF4sGclTahGDivafTxZTkGU4OxSld0fX0WT87ejnOH
xP7NPXfqFDWM2sA8lCYqUIhfKYaM88SkWAKQuDkkFstOhdXVJqhlP/CL1VjIAgQMfC2FTUP33fkz
clYpOQh9UkArH7EeMwUsdfMaqgf3ubemFL67xZTvoF/EixaflfFMxSuVaeqN+0MzYJP0RFVzuHY9
CwHBXbvc1fqQWHskEnsiVP4LYhYDG4rU170I3qevR+KyMB1AnjkcI1ju9EM8zYq/JQ9V66OCSn+s
HCnkw1pgppesBRPT42GvKmXrWkhuR9NDb0DRBFaEW0Y2LFDRb0BZ7wYY0DsoaWrl1dJBHlh+8PbY
B00UlMKpySpF7BAYah/7jVtfeRF7QBdqHcSCU3p1yueKUejvIjuEVtRwUAz2/18Djd7cN79BIrhH
j0TwcaXaWYmRv1se/tF5TB67NbbvJKLhTEjfpLFoi7WRRbK0M3dfS/yY9LSmFB3JfpdmSIHR6r1F
SeJgFy8ycZ7De+sY/uuO/rb0nObgIl2RfbcECr7NiuW3X8aqQntT6gv7HUmBLqK/KVz2fBuDoeGj
/rR2DkQs8oXl8BykZOVOS81OGdOZRs3LExWyMMoexINoNjlwtGN2sZROtL1jewFwFWpjsXdqL2sq
O/R2J4inUTp9C/zV8FXDneaTA2e89jBgzg0qXfOd9itHDFcxzI3P5nrXQLhZJ1NHrgtw2rQZ4KSV
MtF2Qr8yrVPB+eHtBJyPFbJd/Uh04uGUjk5GpvgL7qK+T4zJvsNwWRB7/7jVEhONnWUiIkQXbmm6
DAj0r0aZdZx5PyZeL5LqRcWZX6Nl4qhpN8R2hEBIScJWSek9Ed+C212d6Vvb415Q1rHwt/eXKhu9
2f6L6tv9Jw2CkvV8tVU/yT96cZ+tXb6vLoW50TSI0+bV6b4q45qUtNIFaXCgyPdecA8BP7W73kGN
UYf4QCzEDYFfuEK7DrNzmbuiXt6htlZGia3iVZV7kIxtVpXqmyWrKE1D00lR6Z+sk9mBeP6S0njT
DU+RUJWAEde7S04/yHGtxbZ8k4oRSA2/EYius4xGBp5v3yT79PlReLMz3xJ0lJGdkM5eKKvcGo99
xXYtpgPXudgq4TYMJPBvOBpQtRN++RGSwr3lOdXnK3Uy+4YLORKYwlPhgZzc7af2JJysJGpmN0/a
S+9GWCf4S0xfwEFTF4gaE8DBXEN3cOFQWcyxA7BR+1RZEuwOZQNfNnJc7O1GUIzAD0jZ3f3JwErq
sd/B359pAzpKE1cy5IgdnkWxhQznj+E+Z2mzhsYAzyhCqx/SD6kQSR8v9XHnAXKPkzyrW43BBR0K
x9U/4IM5DQycQ8nk+4H64jaSUsuksOFr17dVnWqF4M9WX5yjMF7Q6oUVxJRS78+j+OutpGiUBIC+
59xO8uNlVzoYDjO74CMTDsVdquoyv3K7xpOvASHow6nHOFHxM0ltfpfIQswEpY8l3pjIxclg/3vS
ERkQczu/M9S4fSErXt4y2eetETMpU15NfqIF5zvQ8HUCdcVIADOo8oNu+Lx5G92+GvtY/KZjkAUa
esUMjPSmiqZdBYW/lYR7hb/oRAZzkz0vU14gjA5Kqh+ZXTpDGu5AfBp+Q4faiYRkUKgguTYIPkND
AJYdE3n3n9vkeoO/zip3HNomyycwa1wfuzME0k+rA1MnprHtisv9XfomS4fIXSr3Ig2dbcdSDrUZ
EsYnBivhz8dA8BeJaTLZwk6oQ4PvIJ5uF8aj6xgaaAXwqgbEWHc/lM06tB5DrFeBPUDMkRzpRTfD
9z5pmtgGkvNcOfz3DPE5y5+qHA/gfQ/GLV+wAWskh0bZf3PACKIWrfqYL2N5GtoEwLIkweJiWvns
C4akkaYKFh9GkhMpwE6Yg7p86ZzUXR2ixN1kyBqeHlt+UczBb1ffsBUWRYF9z6GMF1kvqjVaTgsN
CACm1LaQRJNgHv3NsL5QgYuXog3CXJ1z52IhOcglPemFRj5j3xr14+uGpI8GaQ1314DoNkYFcPec
H8UW/WkhEBb//hTeqh5XZkZHu/wlrqAMsEtAAzhXzTHWoGi/u87Kiz8fn5lkCDVdxiRxN3KC3cmq
IbQ/MgQGHuYm4BuVyD32NlsrI8KkvRFhQVg2Bca2TBrp/4sjI+KD/Ocgbtb1ikMga2KFFkuOeZwe
cQd+33TzgnL84xFC+jbeJ8eRUevgeUDkoI/KuLQ767W0Iu+Mv1v2Gy/YOB/g6E3vveaYHjJUSJLJ
PDOuUUPSaQmiTvr5+wrApI/iCZIkPEK9Cf5wp0nY1hDhXMDT5MKpTSEd8Ix2sUeIAsyKNJSL+kEb
1v5jfdECob3q4bxagUAT1552RfQ4LCEEcPRN2lmmjgcJZh+R1LtMEyu4l0hpna28cNEeq8tEq3VH
t6LbyQOK7WBk7SuvEE2u+09ydQEFUspPVey4xaI6BivIjjw2Nkxuvkw9HAnqmQux0gdjFFLiPrBd
6C4Pw2sGuo7ue10gLOkpJTHlc76b2TP82sLyf/IjdOfd5/XxFGuEQgjeeUdMfr4/0jzgYZN4G4CT
bXjNMNVxR8qINTiTVWqo5H0fXuU6I9Vy3Jf7Nu80SEf8FccgIuEE9zcyNesBWZl+ndHgh4pJjY8z
hcftVBlh/nmbjB3jfaeWRrCC5XI4H9attaJmffx/a6CJyBBYmrXy3KPsoIsQWYUlQzLtV0+iFkIn
KQAjJPxVuz7/4bLkownH7DZ1C8vIGNgcexcL50Tmd65M6hLzfvBJlDwSHG7vd3AFaRPOT3gRFiXc
hofMp39ENIspchktMXeT7QJvy9qMFn4Ir9aGxOI9/1vXp+wUGMp9QaEQbKttXbF6jsOecDihLbhr
2CZgAaok0dmaXlH3mni6ZXK2IBPfyctwmf1hSbIFMIe2Adm59R9jm1C8whElq4elwaPpfy4Cmc+e
JX6fSSkFUH9DzPFTMrKqIx76tfRWzcLnJzj/5PQIFmBBbFFbRvFi/8A7VzYFnYGrJAro7XIe864L
84ZL6GlIYsIBENrKCt3+FR+5vLXy5HB6aK0sW6p8m6CO6dRqdtqPw4DffHJDMWTy7Lq/qYcwm2V8
92hWB6cCd7xhdy2uYawZwpvI843tv308ubym+2ITgauN3psK/rC+oFb7jvxRSqOGQ1nTe0F3GcNJ
AG2QXH/RhTLsnCo2+12QtCMAx6x2v0Qi4PrX1VtKoQjngRZcEogROZ82MjJnFFgKRer8QhLoBgS/
DHrzjRDUK25aB2rHv8DjRl4zgb7UZvN8XgncELp8cI49smJa7hjSI19KGh7rRWORuTAzKXNPaR/L
O+IuVineHWwfcaNDi8tRvOmZpDazSYK4hJH+dwrajAy3gmbTYWfzA04qIhXo52Wkx32rAPH3N5+x
OB2SIpw9SlZe2oBmLmn4YwDQuDVPLt0Q2VPc1iC7wU2QW6SsXfP+oSGMHdO1wc7mbwLiohINHHjx
mp0hU43emEMu+Zk6iel0gm3mFAqBBsN30hDbmXx2IP06yt1XExBRc756S5KEM1MI8p9n24e/PGS+
zp0c0CQpJmd1mFHU6PdIzlFfv8wV0ZO13SdxqgVLmPmr2ys7d5UGxQ88YwoxeSmvOhYi0YzbDmKS
bB3z5b3/0VhCFt4mh4hYXW4k4BpGKKgCctY+e078K3CKm4xP0kapRdFfZ91DKyaow+gbsBYSMv3N
AVipD63soHRdckET2pAdfHaNBEJE1FBmHBIyKvbs0+9RkPL+J1C5jEmQu8RaxUmG4PAVHqE/CgJn
vfp0iIDupPjUCoI+MTB1C42mk5TLVao9sZwXCzrWPHIDYRO2uRe88Y+4f9/SlkMH1disgITZfcB+
wInQyzh5O2FaRCTpBXuTc8twftkPK0LhqXsN78QIdrD+rFBVR7avNG5nHoJLtiipIubPuqFH98sF
XmVgEc/vvMYFq5tM3rYuNE3UynwPe9ec66w0NJ8oyh1kyAdGZCvhuSJA5pjCvHv/MtumGapl/7ZF
qYr8yEQXsHLoegSFy/a51jwK/y2Zb+tPCyF4iYR2/LIbeKYUbIbZSuBc0iqHtPHOgFcCNKlgD90v
W6nweYwvsK5LK6sPsZm1zaFk8NqQZ6ma4M6PS4eVupfWAaqxYDB3q9GHyUSvvRSd0GeoOUE5ovZE
OHmA9qcVo7ve4QUj0uCUydOxbO/yzlmY/dmwoCR85E1vnDDCj7EyjFJeQ3GcoZXiTSe68AZcJzK3
VVlEG/SFXp/1KwmQp2uUi9A/3SN9lZG/tVINyC7PZ5ecq85WQAexF5nsC5aCU5HpzbQdGmcXlrb4
+zMRNajz+YnYPja9HYuKFIUGHgNlNXlKwfrcqjBE+6+n5QfIOlV/byBdVW2n9+vLiKetCDws4Cqo
fN0SYTjQfU1uoTcVxJ6BhEwike0TrU6nZC14ISleH0N3aDcFWs/bIdULFTJ+VS6S7O1zWqZG5db0
+ZUJDMfviAhx4Ka6oA/O98fquW4IvjXM0eZp5UUZGs164TKHCNlaxJVYkVorW4GmWA5n29Zdf+z3
K/xbptGE8zMY6kNwdfBLsTDxnbVQy8ep9txrlRpRlj00wOWI1/o7YduM/UjZb9ALiPcbT8vw4pWl
17OryQ4w3i/mGIHXgDIIQo+kMsvZEPHuYCNd6i9JOyFsO9z3G1GY6/0rsH8Ps/7v1ZQ2sF3brBwj
fu4YdbBRKheIt8UZvx3rr+Yp0FxuiMcqW1USNOxvI2Xz6Rizj7tI2J3Er0ah0Jgz6SAU4XMRQdmG
JzVyBc2ccQhsYDHQ/QDG5tm78GxlJsoFofHOErg8xTwyZ3rVCo5PKOdY7Jln3ykjWH94hDzKuaOV
G91NsUWt6PuQ7e1OOuM5BvLGxKNga617+gD6kykFUfH+ZvHdJ/2b5xQcKj357f29gnUqO13TPviY
OKoDAU5CPu0f+HkajXHjqlDImU4ENbzIAGuhID8Gkg+mzTG7UKX06Yj3sFQynwO78SCkzfeSIDKj
o7x+TC35vdXPARDONcdNRyii8tXaZ5Wk73wYvJ1YLFWxXzL79eZB4/M6sgd1QAmitNMxhiQKiIUe
77ZIOml8BM2+u1AUWnxfl7ng8dXcPNFdpa/ONvixsQBc4iB15Xr7nxe0C0YeYs83K2tic0RxyIx6
yXXGVtMiYcECvZpqY7TE1dGDET9v4AQ8o4wmv73r/T8OQ/doeqSxq44ycV2mFmfkx4YNcSqGrHnW
ijAJ0N0pCvEkXCy9bMrPEMSH7pXMDFPAoF+VZvOazbV+KONWnHB56RUm+vh7jAl/CC1w4QCAsNl9
k+awXajUQfR2wP48uHoSpXbwwJncbYEAi3vPXkVdWcQsPFLyqxFZYraSt27gjR+mb4crYc0rRE7f
hiDK0mPbEINwtH1hCjKXd07c3+PTkx+Xw9or4P7dDEwEsD0B+QJK4koS1gKSYaKmbYiJbwQCr0u9
+Gb/UqtddZIXJ+gSx/UN9RPKappuWVJr0tB1IH0cQouLP6TQyXcBSbfzoQC4YbbT/zJaoaBKzPWu
qrJSTN2ZQ1s1HpjaD3WLIvvQPa50kdKF0k/+R7NUhNB3VWSjNHRXEIHS7Hj+Opbtm5FmejnvVZy9
NJ9VKyhQxI6xN+q72Imw0u9jTy5vf8vHLTuj32FeYnenmbdKgVvjvBCPjw0uisV+17H/LHtAGccK
pU2hkkidkph2fS1/jr8QzIKCVHYgNMFd2szv07eDXVkCH4992mn+NPV1zT33b5JgizYA1jpa4QJX
EZR3sCorkOz9FWzWB3s6WKUKUOQkAULHD4KpQdrFOGs1PMBblH76IYzmSx9hYZr0m9WWG+9PTSky
LewMvXELahmiUBLg9sIxZsUmEOV52eG4jxZpIB5Rx+YGkHt3xdW5TdhNde6Nq9C59NNU50QDMdAx
p+BUy5Mqq1c9Q1aLw5A39BWLGy849cHpGr/S8mCxFIUAz01OKRk3+JBnokJSDrUFfPq0pMBa6AaO
3wG1Y2K0AvivDDDLjzlbpPpLBQI8J84FgxxZHvFBi2xvgrcF6B9y1vsFS5198Jqg13oL71BcEova
vEqmdMTeQ4qDR6M7znBhynjj7moe2GGFMQt/pOzg+llPHQOrHtHJBp6isL1R9FhKQ35zs9gs7Io4
UlQd9msn/25eSfRqJ51Vr+UF8jJgb7fZNI51jqn/EfXR9INB6Vzt0/0HfxpHrUsviqMzKqn6cH4p
wJdnj1DicwQN4dLvGpvY5rU7rVgvtxewJM4/uZR80vYGPMgvoGstT++K/kq0i5oHDUavZPmNie6e
BTq4xvUfwPucqyEakYwt3PISvjTfILc9A4Nx7ZRnydL1ks4Ia+7t2zxyGonYDpXe5/pNdgcNlfsV
hUSgmkUdmmIuw5hqAR4DRH4NBzdTjUV1pWFNBxkzPIeu0lSC4qGe6H5XCBOSj9E5wjfHUm0CYgIa
ZyJr0XjdIYeyUizfeLayjndHxiYjEAn05Vjsr9A5yzu3v9oylGqHG4mbBCyCu0AReeczeoOo90dS
8X6p5uKk3ePdoc/xCWcSnDjDcp6Z9nglub9LSkTr+qgCj//YA7ja7gV9+JVQdrsdxKHdijPhZV4U
nYf1kMC6S/t1NMMH3q/PAowzDsMY3WTcS0s0VjN2OFAp++tUpypVxONaQ3m8FKC7gjmGsRPKY8gT
tY6wHkiOuY/bYmn7Ap0HnFqCwlpxFrLxCaB0306HDY87PYfC9okVH33gF2nZqwDoBWhquJqNiJJp
nDOJJR0GDEeLPhOgx5nrPYYBwIpMDtY0YX0mgOLHvFFLUAQKEMsLZatOV1YU6Y1Q7bzgkMjHZNOH
QoZhHUAnnYdTJAhhm4mOXG3xATtyMoZgGqXatMzs48ehJx8rGP7Do8PLP4PeXgP2pLnfvYulpnXh
v11kPEVVsK4VELlcrwGVChaYwwmlOCzt4s9bd/sMLuJlm+hyAz4oSxpjwTjyAcRj5Q8uHMjCb6pp
NZc+3G1AKGrdEWI+amF3ck6ydonlVI3uawsKJ1JM82xXQiAM28M7hPxzfcvVezCvm83dTnsOg/qa
Y4oL8F54nE6nLnknIbKa7VCfqbu2ewlnN06MSY96U/qNOtBdQhK89U46zs4RazNM6LNEsVX5AOjd
C6UAShWqv0FvXEENax1VqqFNdlPPbYTvVVHu1oHFzyP7yJEuEYZAA+uMrsO26+hbTrjKV5C4xoCw
rWocsMXhcihc9zNClVohaXLk7B0XeEWVc98dyIwBHitRhKWlhTrZs/eCH2NzZNzHvk3yZSElXe3f
YjzCvgcLC6VHI4aruB38rTaUD9oT98yyjqASAN4Gdyf16m7jXJpOMMJ8J7gQbyf7nmN4yzajSPib
h3YfRSWrRmajnPdR2+85mPGluABrO/DnwwYGi7Zg1l8EH/swyxGxNlML4sb7XcJwNF0+LAmcUeEf
No5+fxVyJU0M4MAELjmJr+h09UFx8FyNi6lknrQuHTmWjo/KSv9RlbhEGFjG4TnY6PA4o9XeEyWF
ENFoBVh1cj0ufb0HzaXnSHaGPKcQAKCUktQWWh4wKFHiHrCwq9O7BjvONVEmmkHSh6CRwAhW7E8/
TvsMvzIKnGvUeMpPFW6tucFa5sSSLwVPHuzAhK0GquREzl2hxCOS5suCyD+v8LS/dhccUa3zt8dJ
8amNuRQv26zJrpFXhdoqL+IzYSJJ83ScHAN5rS8Flzyozu6LZFoAPpReYim6muVobgwOPdlhM8n4
v5Et14ybxFNJXyEvruzyeH6PKyccDCnpIKTz3zmcHmHqX+PJ5YHJ+rlj4/5B/J3dYNubTLz0zd1K
/Qm8at9ZtqNdiWin/UXl4XDZ6Ed4TrhooyyAPqwj4cAWIrJGvPFTYvgigxjziKhgMDhqyIOwP8uD
mWGBhwiMNa9xXB8yYf3ZBDOS8wtA3JDhc9sim04EZXnDBCE7K03FAeIw4UXGNjRTjDoIT8W8tSUf
WcvEwoUQGFeoWu274jgjOfwr1B7YAoNKxENO1WbjhBP2tM1lk0kGK8x8Xg6SEYFlGnupOpQhhEqt
rdQxncUOVc1hkUd3WyK/BoyEo4ShUVuV+WdZC9el+t5+YS379WfVcd5g+zKzSpt2RLg32AROgF3M
imUDP+nBigrfRxE5VfOUzRWcpT/Ovgx5+9tJZQGwRMBoxHfJPUZJBuN36ye4kDMQRm4r6NRCLWlU
HZLI2RKWSmI0Si+BDbxo4GwKmIOlygYrYAQRCMhZzqtszW4ruwkms6CeoKAlPVFAE20bBK2rZJJB
2Nk4st2j53TYqu7xIcyPdzfq55irrH+b0iS6/BUlOzdY8gakGBnu+T/rGdMLkSGL4miaZr20CdNZ
GfOccb4/9wSaTa0AMkeIPCYcOR1I7bh1EMiYbEaS0xcDHAnYkF+RylVtwLI1226+cM0a4aLO1ZKo
FpSFqzLRSdsd9E/TbgJHGipnSXTpLp4/WctfHIOGiQezRafX61JfMs7r+v4yCQH5m3DXpUpJDESK
tGC4v5DhOHRvpaZZMgG6HqQLXmrFMbosKKukqnjKXmut3m+7fx9VwVlE+PjkA3Rrwz0zX64FIX30
O62DwRMQYPpuyIv6gxg7UBDGcKdD1V0Hs56c4vyozN8+80V9Po6APL6fCH3tBH7wAqLLkLWjdfTn
wRdLCIEMYmaeXC0bzo+MoQd6ClkRT+3MrTPI4tySCaLWmCfXc3vi0/KyaD2dnmD4Bq+TWB/R6veQ
ghDk+PhK4T7v1vEEGJbntDl6PSA3zMxibpbnsBgJvc7m/m2f8CAK0BlAh2zbUEtGheFCg3+yHx24
EBOWXNkJ7LQSPSlL/esIUermOEl5RNq/7lgcp9Vvrnu4xosIJs0TR9RhQhEay568IPVALH000sAq
6HVJCiL2dVL1vIyyJRxANHfncQH9hPuK1Pl32CIqh39tEUIWIzpE0m13dT1B1F7sBN114z0hRGjz
HPdxwNRZ+m3g2/L2lyMymXUAGPGjjfHbd3PwH/YVH32k7r6XKnr5spqjcDLhwmFA64zbSdNdNpZa
sEPVi7mbZPm/0oGktmqEQpEUM5nTAPeRfXrp/XktwbNjh2ODi8zO9xPU78GrsDbOIiE6wtpsz0v0
IySKa2Qyc/UVbX7/4tt6gMtWpbOksudl4EPeRZJc9FRIbpTviV+gkNIL/mbj401vM/5aatYQbL3N
dT3gNbLp9bViT6zj6A/a6lG0qqtRhVpgoG0b4evxZvRXCbYeamm2w5QfXjyXR+yLmhvAQcTT91O9
PWW9ie0tsWzLfb83bVWKgji5nWZ3vI1+Msnap9FwZVRZj6T1eLIBMzacnzfnGBZ/+p9BNKciDwFb
Ythf4npeqgRRPypcTNNSFUc4XnTuRIgvJgmCu/9bHiYtgnhZFU3QZsSOJkYEzL8RobL898nQzE2o
IGSW2vEHKVOtY8kh6Uq2xtiYLiOsXPHKc6PvTIX1Ls8wVpxoNh5hISeHlld5rio8s2IxH91XxaAJ
MX4BFhm4fbhxfSJMOYLQmCNj3jPcHXdTvIp7Db2sgUXe7KbfKb5Ro3FXIZenxI6G5hgBn0j/DvTU
9L0bnANyG96SL8UtxXjgFi7BXISuuI9TXtuldpNOWJVYPB4ugveYAGFDOqKHssrTSeHJa2UIPS/k
VBQLgDEmHl6576kAgwgJe6RV1eKyyKL8EnKmIhLrxIAon8o3rQ9InuuBzeY6f/hgjS1J9N42Y2aP
H7/wld2hEjeUdOC9S7GpdKLA21LJ07fYUAs4tn6zBUCZhqnVU0DgVt83JOf6nVW61tVu+K9UqAeJ
MSI7RgnsYmjXOKjR3io7XmvcIPpnt7gSDx//kRsTSxiz8dJ2kwYI9jC+gruBxA0X07BQ18RbIJx7
GjjaNjJpmymXn8cdi1dXQzpGzf7GKAT/tWmwKcfwHnsOttKE6WSKVX6fgktbOo37Jm9YyOTAn3Nl
UZsPtl7RSR/UbbCedeSut3yegu6e5Cll/zOIcaYzso68e2aFGUtxFASbD9QPPHsHAvsVMONyHTa2
vNJlEEv7f7qmaHjFCbPE+bL60xU2XYGzF96jQCatp25X4wTDy2L1dkIWeediCZCyVdxk/zxTZb3F
rk1jMwUPy+W8jSyd7BX12J299V3DxbE6K6S0ZGgLu2ws43Oo3dnn96ciRZSdVkEi0KbYCCn6qhVo
DySnDpaodDu10ZuQLrk4yshGul5ckXYZgKxzKjWzpBnYJlUSiKN43Sv762jNyxLx7VXq1S+Br/RT
J+QkuH0VPDo0vPuTvH5UN2qboV340HQaQRESdkVAZykGTnAfMHP78WOjQN3XcIH8ZnzYjcDIDmcE
/VQC2V8zh3GlNuJIkX4QsgdoUc8dKV6svyotOZlb8JXN1t8DAkqf3g4t8mVK4QOVWgGqvmbM86mM
StcCEuiyJQ0dbh18MLJIHSZ8sUJkzVY+TKeOfGV4ATe49+kgeLbVPSA6zwtXbiSom3lAgZG0h6tY
VFndpsqCzZwB/bi4JvWcEizraBcPoz/uWnIXD0ZfM/KzzOe8ooCd4+oHz+9E0Q1RVC4niChl59B7
9CRHzzdIB0XYYnR0QPxrF8HNcjCauyMG/kpZ9VtGKfBTqJ3PYBE3v3a2w46MT/Kq6F6FkRTmxtN6
A5c1N2JnafOGb4s+CdvfqcQmFR+yun3PjJgnsyccaOFQT37OPcO2lVeqlVIrGQgZ3zn5crpcHDB1
q6Mc8IxLPpDTJ6CzTQV0lknG0zY40b7D3vjK3GbqEZCYU+DhOJ00NdF+MC4O7PRzOaJ80necn8Qr
PYA55xr71tw3YDNqA5F6bpTTJU52t3zuxLvBxwV1yKgqV42T+lpEE0ZkguRUhScgfqsydIphs2YQ
EVUKZ55l6M90Z+yJdlkT01zBehd8QJe+m7K5vm+yrfU6QosXpirfDTQgVogP3T3LcgmW84ZuNcHg
3ZlUfo8Ik7nJhFjqDmLidd6F5022AHhaw+O9XW5S6ZsKuvpQ2rEMIhbaIkdYUx7aeOeJAnNKTwMg
K6urbc/8+pKDY6NgXlkegjrmUpria585YymE9V5ioLm11Zk8kPmW9B2BY6/REtfw7pvS5d1/V4Ii
WECzYcxM7XKkV3FoCDMFuUBRwa6afWpflmdJoUBt7DbogfABI0uTetbXoeCoXyK/j5OLwvZDmo8u
vgKrX33D3acm+n1lynrZ3d7Ld99Ht1Rs+xjvw6+BDcoHZhhVtn2tZmopQcDSy8+srds1YY4/fN/v
++ty5VtD7yxbUTjbEQj7ev7iE5sd7/tIsS7Oh2lAEAsdoUUyo1nxYlMmu6toMUsYld19Db3oOMxx
qPVM7GZTI8vSsg4BPNuy7cUlhVd0UJVpeQVtiRjXF/pDnm1vUxgp7jCXPWkkAFG01G8PrwhNUUH8
MeuHxlxBxpU461JpNqbInk1UVFMnylDil2ogCdlBPsr1LrWv/yvNrZKUib4RWkKeNtx6R56TxAZq
Bzt92l5QTGfgcN6Ypj6/256um+SAAfcDhltjgkssqG/9ftPhInyDwrDGotc/hIW8jV5F9scdMf2E
8HYWioo6sJBHi75aC0LqAfcQfBj/vPf++/OzidD07+bZAXq8mOPuQXkwUHX0eHmfyGBuWPn1P+5h
h2vUfbIewD7HyUaDTeZD4ZnCQLvlGtOa32niUopUwWBtTzrYPC03oDvKk50pJE/D3B7sRHTn0/4y
MuUPZUWwIvw6BvWoJ+tYlxeunkAQMw8DMPY=
`pragma protect end_protected
