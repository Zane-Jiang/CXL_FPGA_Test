// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
QFmILsoYSCBqPpr90vsuKHgdyYw7wLXldok0zdTZGgZ8Wb8DaccII3iIJDGIcpJIMF2PnQCUcFE1
kzBIce6lZpJOOCJ3Ry1LIojnql2IzRNVPvJGSmo5nC+xSDy7mTPFacY9i0g8IeZD6D6sGqnk02Ff
+IJWUGPG7IWpZtTM1i94Ve3yGVZeh/SFVWP4TbAzla/T/qh5isNIEr567Tac1itrUYBmcMajIUkj
yXQdFZVe6/pvs8P6J/u3rssZe70PKCVptP7yNA+iTbEl5TaiDCG5xNMoR6zS5/zcyTH9kBL54BI5
wnJTTO/DGAW91BOGloaY3kPwffHt7bS3BqQRXQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10560)
Wb4Bb4Dq48gyfWMNKgHyoo54OgyvVzS+3nxuD3TTyUyK5ln+11tNHsZFumBO1mdlZPGrLjXU5Itr
Owq6bb8tL/XNAf6df/z5TMjXq4gCJeZoS7QLbjZK7cNmPetyTB73RgX3F6zHeO/bQqg2fUxbRgv0
V840gPv9q5HPBXF5TXeGNpOtBOELUzccznq4ZYL51K4KAMq7k2Z00xv2I8P7TLNaKIv11nJMbsS2
+h7Tt/4mo1ZBrHJeSlYAaczBM/LeO9nL/SFOhDxhmJFicOsnJdbaWCBLRX5waZ+MLaW9wpObMFa2
VrynSsUWaszLKXAY1Fms9RkkyBt0UxdU2hPV5pTUli11YywbsNvDs/DqupjNNDgbRq8Q1i0k8B6a
9+teqqF2z762mfVOb5M+jvWN5LvK9w6eAeXuRNAGSMlGeu+Uf76GRZ86XQLe1v+XEz1u0+YhW7bM
Bn6SYjPBc5K+hkS+8aXtM0K2AmhUqHNDIDbZ+cnX6KsBi5M5TVTEDOeHCk4SrHV3aj7xcFbo9Ln9
3XBJQseVL4XpypTFxuX4eYN9qoZ+fi7jf4notJclrFeRLnP5ngb6hJsmE/WqEflD0/Ug8KM8oo3W
DUYjyyEVjPjULoGtWpZRxk174KsbLji7zzxVyu4vilsEaEbYN0stu0o9oqsoyA7t5L+zduHe0tCi
lMbRmNLzCy4OSlUTsuwhWrD5oi4Us99MwV3IPQAZmqEmLkq0xPd/n7ksi0MabZruqrJ+3VuIVNFJ
SqPMHTA8O8ioM13yDmnOn1KwaDsWNV3EVI9XABjtqDcRaKOYL0qWhdpWdCTnGiEe/BVoH0N634ye
Ysfo4Lx7Xl8c4MeZpO2aoqsjYjdrfR8EDMM5VCNKphLtJEIL0ZVBki6Ag323FxgTcBg5dop5/A57
IEy4MwClEdpzTE1gA6Mu/6I+j5f+lMbLd2EbuZlYeWZHbFFHgvWgf7jwr94qNZJPyAMQA4oIRs8G
HMTE27ZJOQqEITV25/IMjADBUDBD//gtDPA7omszvnidiFAUerHO6Ban7NPKKaepC8zNoy5Ymqjn
yW5fltIDIwZLo1+c4bnVKKxtad+J1D3P+j4/c1zT33BKyYca1njLNgIABwCHH3UWkLNYMfD7ipul
eHIeqh/caogd3DY2LWCNmwrmyRRP83clLq7owgA/Wt6kBvzyCB46mOu8FfWDBl+UO9zB/ZkTRbtg
K/l1GDErG+2D30nYhratpltoMpozI1X4OcsXIkI/1mA/GTLXbxtAjUrHvX+DwtF4XGYAePM7OxiB
AGNYjUNiSUpoBlNf8Luwx/3XEsO5QPf8SNg6iwOkaEMhj8zajlmPUacK2gMX0vYLJdtj2agdJix6
zIxomdKgYXwfpuJyYMTwDl9Wdr9MFBVeNRQ7yb56IVTRDQm6OKtCC9v4EoeIwdmp7oTtguaml+6X
vW5N4b5CHMxfXOsapDM3k4c+PKX/f9ZzycFt5KPf9OWlexAIEuXWnm/OsEDh9soIKKFEg9RCgtnm
F0ciDCuc8sEkvUxBQ67KwnlAbFjT3l4vIJ26eFwroLsLBPz1HUrazmbDtQO0wqmAXmXm7Yxvgzp9
eWTtPgI4npfraF5goYWNtm5AECMqZxWf6UxeFnVx6QFQYXU96FS9PA/+W3SZDfokAyDCM2eFaMxv
ItUqk9DFfS6H1zcTx3SJoCcGM54AtKnj9Q2mudRfo0Oqgi9oUddV+BKwPZeKJtkYVXiDi6Jmfjd4
wMME5XAarPoCnTzQUB+sgOw88gmpoUPfEPYGL3UZIYwksG3abnAdvmxOACoCcTojEBiJ/Ua+6Ms3
aLpg2WoBw93nDuBC2K2bV2ftpGyP3bRqF/oVh3Yp+Uk2w6tdoD8UevBsaq+sklRsswNSgUkkp3iZ
+oelqdJMkoGdIvBsP1e5oI7yLB12899uFtsCcAZCBColY+sYSo6FGqtDSZRy4F7s3CfnBSIGxheP
ZPqqb+b3itbAEmMIspRfSXI1UXLsOqpUuDYoOx5XAYDW78VMkVdHtA23l96O/mfQfOFBBIlmI8hI
GMMA1oaKcEQLQ3pzW1bDaxesktyIu487GtIEedGV9BQofIhMSwRGp/Tp/pBfXNqvZAB8qEhjWWFQ
UDHs5BOkBhzDpOkLE6to6UflnmhW1pWO5ZHurTAn1FaUbM7m+z9WDyRwB3+56ABkwpdf7CsBfQNd
Cj2pQYoAgr1/64F6tf5NVUecOLnSDCu8iLCnMSV564NxC1Hi+OH6EJMyPqlK6FN/TqC2KV9LQR4R
Wg+QFrL1t5t2L8yIgadhq6Ejc6wpQw3eKIKDr8j1HX+IIVyUTr2bcGjdgH+MvNAT/eqnYKIqJB8i
+HR+4Yy9ubQo4Xe7JdRnNamFa/lJJfRMLTGMnhlC/rvG0TIOH8+JMJMgzxDJXmWfe18iw+72veDR
3FHqmUbhj4pbgIpLJlzPOaAM/1tEdz1tNCzzGh45EqvcEo6SOjunVx9PaNqUpsbhRD6YEqRetGON
iWN5pMgz8jccilMyhNEW6yX1gyZPQRPSRcbdqx2F50JofwAmvYm1Ysg33OI/fg521vLJ0c9GP7gF
3JAjtE7dR7BPfGiHossat7G212rbaS3baC70+uRuk7ZWOEv4mbJBKoNjJHJz5WLbu+9mvbfSW8+e
ynd4B56wKbHzxDCzsTTKoe2OSe+DhJ4B/a3Os8Bt2XVpivdmRHYMXtppT4RR5LUKI8vq6Bs0ZeVP
CwmmHwNQxYFpa2S49TFuyKxrKIK2WMyNFYDUZ4VqT05TnZ9/NKU/rFbcYrY7DRcFJGQtNLoQA5Re
9XKk6+K8nexBeokRfk18oNk21HXzZ2VGEhNl+p7N4DpgYrk5UMZwfciMBxNeVqesViJeWAxmKrsM
M6mMlYTVF8cdxlYkhQvyrRmY7Vy7gJb5aLxt/Ap+gGfyeFSlicFRtXq64s8CvFGf7+c4c6m3SkG0
XFl7mISsEuDLGTAoGWhSqSCZLoYqbAV6eUeWN39dDO+3M5HY71y/AluVdSWlyMCQbJDQvX0GD+GC
/zeGNiWFMhYI4CLgZXBrsO4gUxalcaBEz6IkVropSsQXJVRxM/A1HhECc7IZBD5L7qrl0DUiDOjr
KBNBsimKWtDi4l29GoyIvgoVU2LDhaY6B6R2zpQAFp4ORVawy4WVZ6rvJm4+SL6CWgS+GhL5l2r/
dXZFeunjz/mHmmYJ28E8ngemneUhC61KwSeYfxdDDH0TtyGXGoipyKup+5WR7FfrV35MyDBugQLr
qCL6at7e8SkvNU7xL68SGXErZbTNNHFuIKE+cW48GXSYSpIazb+9EaSJnR4vrkT+trq6/LKvtmj0
CPOL7umXcDThs6VZc7ejdI8o3KH0hoGz7N4LQFyrjba6JOlrE7vtoSyMAj9Fg7qx9AMaveV2U5vz
M/jP+EnqqnL6IUsfTTp/AKySsC7UEC+04bMrzBrsWK19JGzJo9amwgavvEtROWB9hCjlvFE3Setl
+A7nJiyZAW63B8IOlXlCPNDbpAhOfyA/YQYeaZB3bNFKADnj5wWmmciEZFlwjiyqzb/ZR2j+gbap
GDsCCU+Q1SvbAO7g09oOhtTUkn0x180y+oxy/TwCBzf6JYnuaDacerpAo0i8Jomylo7mIgywHFOu
Ru+Su4SUoIJxj36jBZBFhbVDDIjlhNttqp72bs2wf3Pxk34LE1zmdj9LGdBCk0EsZyU2Y+LyGx9Y
E0SGeuBwHvP2E/ku2w+ODxaEqzn1jwFhT7OW27zWx/dhQ0zUA0S0dhV2pCxw+jVIzEmACV1AenBg
HrSs/ubfHdDc3jUN6d27fkf7DnZygh1BCToXszR2DQq7eI5JryBLylFDl835y3/LclGapT9mr032
8WVqhfQE6IFv+jGHqnDqARmwJUEsDM44HMNfsvRtf6FXrA6hgx4eM4UIP8jq26THsb5QcfQ6fQol
lFpVBn8qpP/pR4IEkxj9hg6bu2e7WFxRTkd+pgwor8XFVqCinm0SuS2PO3L4RUX1G17z/Esq+u++
rF2AnjtWxTM90/cU9IB+Yja8wUsCSH9HdetK1kAp2nHdwLWQmPgR5p1WO0abDGRYXqiXCAvMZsn+
NnOkvL9vuWsJZhxeavbzEOGBKfPV4uYOsKonKkZ14HolHDTcju+1w6Nkmrv0YZd1zo1FajMfZ2AH
hRp1k2uCkKm4+mVUHT3sRwuv7CWnxYjWXW5WTEyVXeZQGv20w4RHGSGjeapU4H2NIAZRL9GMq+6v
k8ZC2bByp+indUqmvQ6iseBihTIwzO8jNTXQOtFRj47oiNbyclEtNlW8VnrjwUNHPe3Y3AW1RPfc
ByO/w5RDdgcv+sRe1DOhhsMIGBLYriSdnVm5zA0QiydKDqjPs4q6mH1dJu763PAxKG5dzbC6HMjk
QXq//wk9/Sk0SHE3Nik8FnM7rcPJ1byv7zrI6i/pYnZ1yJ1QXXMvnT8cbeKOoBIC4tNLBZd0zr1R
VN/8vgaKLp0M6YoyXQTHdsEHQUb4foYcyvMcr8xM42UUqsMJoBzGVuGomNAkVoQ5lz2KD/eJk1LB
MkgKHBctxv8u0kGBYE4HxGqMI4tJD+a80wX+X+AhK6uJfV95iyCdxVIIE4wmX16IJmQ6iv4LUIxN
c8SBJ6IGatfTyu3itmuDnL2/CMFNP3L/LVS/g22H5DGkGiwux1+Zt4LI9zVD+HUrUA/7wnDPrf5b
UWeBAumyriwoeq6JsiBYbR7wmP1dZcpdsadKhUjE6lJWCSr3xmgHj5EN3y70eWi5B7SWPr8sflS6
VLm7Tr9f3CjIe9aoKc42BU4FGXODFLHcI1Wz6+eFaZfg7WYNlrM+m1GgRkaJcQjM4QRFiRyvpVK6
52LYmnyOdxKJTctHZr9pIJT0QmDSDt4Nd5LJoECEm5G8lZs6qXkMERlOc3imuhXyivlerjLSZGGZ
+/bYvbT+bwBj9WAmtnOGc9kFN2vG9lV66FEkMjftzwvs6sjxA7qL0q91KAGHtkL+Gqf298Vt2aZN
yHQ77rB48X3fAyBYb7hy/3BOlHGLIBgjY3EO118UbPnFGbPNaYMUNkWKhyLH0JvouUTew12qKUja
MbeGtN1m9txnL4tX8cs0KvsdJ+vdOerpLMx4UbCNVBxGYIkv8Y4JGpUPYnPKW3QlkwFsQ28cDGh3
Ge6QkKvgr0n81iLI+Kq2vP/vR+L/sDAioLziQnI4o8NWovYgXLwWJWQX4s52NeTfvG/XmKQmNshM
31wVG0IybVUFPHKWvQbn5dM3TxvBGqWT6ZZeP/Le0v+8YR7JAgPmzRVAMsSfcpMbX0m3wUBmsFkO
DfYsEJ3D6oTOYtcNep2hGgpNJlT5kM+LpzmxioZR5gY+dTfcDM6cvO6zEIPc4Kyju2MK0W+gbzk0
vp5G6SAmz8VkhSxK398JKshD2bIF7vYaNTQ05YAC3tw2VMJZ6IFbSwxM9Q0wok1hMkcjsoe5c0Y6
fEZoVKOG7ulaJredmxd553QLTKMf4qRAeCY6Hf1a5hkxw2CsLAJ23ac7UOGOcUr1jEJdgthwwQyE
9+cynqZyWE96hdrG9DGpleXpQEV6M1RiosIHr3QpBNskpUsaSv6dSVz7z0/QcfgSQHGxcinEYgPF
tbTaxTwhjgt9Gstj6PMGx5TsyT8BMZHIfGeVuddIkzckMubrSVY45ECYgDQSVVs7v+8xCL8ZCvUl
b+RycwKwSQdBOqrVgIsAYkG/0MrHHJK+us+v/J7Z3qW1u2BkFNEbEZO7catWWCy0hfwg8jEcmnQj
1uqzrXpY+jFYAq5efMHJFE6j8Q20Pf9d/qmOxFMJDFRVCAPTozhMVAcZLhVI21BndvUPRP81eX+g
BK9ysin0BhvQT3fwGD4CnzUsNqxdNgpIRpcDd3l/aqPZznwaoyqB3BAGXoWhXhfkLPe+IEChX+YH
2GbWdg6GJ4uP3reSE+RzBQPnRhkqcY2S+sbQCgyuL0OOVHH2tszTcECGNuvIF97KK0lJCTL5sE9p
NqbNIRw0edyX8R2heKeYiMtULAaR+ifGDuI5R5sHC1ZknOjMlfMQSifT8R0HoMwv8yH9IYEoR5t5
QbDxq9NY92e3qwGJVU6wdOffE1dHjK8/L1aXmOv3pU+n0hP/9y6hkU1NOB+E4K3gINdIexSd9N5O
CU8cX/JBie9xhXwOV2LjuUXcMXEQAO6C2znJUnJvqhi2QBJd05e4YPaLHLqOcm39KF0CaUuxyMn/
xCbFvIjOcJgJeeoCgxcEylYyEW673tGG6lFsU+d7MagpHIndE0CUyiHeC52e88PzGMvSfZ8imdQk
11ZE7VJmLCr3CcOLmWpUgi5c6YrN+XebIYvtqm8PFzWa0BharAB78cJ7HYThhw1fQAFh2pODj3Ke
ec9mDFCOUX9Wv6PsfmFXFVg64XN5OcqfKfJLxCoIua6mk9e21SgXcn6Yl75jEjkNFAROJaG3sD5M
PjMk2ZQoaDasQv5z6zZJtWAL2dxD7JjcQF5GO9xX0oE3aHCL3tf3oi3zRqCayecP43j7sGVGTNUH
9frWXaJN8IfU+kk0PTA5Rp9jE9d79ioppGEb/WF1LegUyuylqoLbwTfjGpx0hMxl/vsNJQ7N2zVM
z7Vq2d87cnGrzbM0dZtT++6CWE3qd/463NPsluv2q5AeE2XmMsBHF8/3Z0Zvd+KJNWerv6NzJ/qn
5HruT7SGKbR4Dj5JKlYSlLEiDBEc+Xq4tvGLKAIXiYebDU0fzc/T1j5mUX2heebL5TYmzZcSUC6x
z74oSoGMW7nHjq8NjrozKNq828wCBgpkTjmX5rLTsSkpLwwX+2zI6xLsltT2eO8Pwb7KfJLmYnnF
FS/HSgltsIdE40hgcLYElbvCUOatQjmdla2nVs6BYeoKjb2UIv7QAVDgdKSEIezrb/ADqliNzEHV
AXrfc0+8g8SwhUIevAQryQ0GUR166+ypsG1/RFaxsPKdDWrKn/ktC84K96gIy1q4NGAbkI5VxY8/
iBeNmIZKMCQrm2KYtx7q4rLg5oxLgJjilip0W5nVPyK9xlMYMNqi6X+JxbkYag+90dui/GLjBAG9
zWJa3NluCe1N3aqSupdT7Dh17haeAOU72MbsMO6YpDWyi1R++ooTRLM7gcwdRzu+NA1U8M2EYbNX
sgLSmb3GTN5FodnG3yK1J6DS83mFk1j+2od5NIUzgL9kQcB9SqmlnXqWctPLk2hK4C0mZln+bWa2
M9bjOU2FznYOmeFK4/qEo907akXBzCURjBesBtUny5OtsFucVwiPfBpMwz/nK9RHNiPbNPcoj9Q8
NPeVXgHIxIvguYsatJQ+JlCpbjDLsEQi5nSh2ZDuixL6IZVmbSVbMCiNsQV4i8hHDmBbav0OiqVk
s47oESsoRlkF0O/zmFexfIkLYWwsHHVihiWkoxR4VRimZ2RsIbJEj6950sHlVG3qEch9yazXvEVr
owY6HZsxs7DYK98iRnK7VF1WkGUa5vs95wO9HViVEoJytokRn00AJCrfPrVpYRwzOUQhkULsojYS
fsK7oI/rLLz5qFpcRPAKunPUmJrk29f3GXtG1TlXqFZXgrcCldbGAbDF1Cn266/2zyfZ0Zjo1kNQ
gQRstjD/tLeKpDankmj74baWgxC6vEE598OaiCrPgC896oGuLVsoyFsOOhn082cM9aV9cuoLMTTG
5FMyUzxgaXb540bxklIg+78nTnFCo2MS0kv/PVtKL2S/MIV08t2LVktTMFNIzgXRGTIjaJBp57ST
1MxPzwPLEZlzWodA8iOG3P2bPT3ncMgDN94qgihrMyXzKNlEsOHpYwoKZhhOT//WyX6iwfX0FgL4
KCXTN0INEKgk47iUPRqehmz5ZPqptwmaF38jUtjY8drckfHlCwMdhzMXUevdPORbzrWr1qfp2Hlr
9dofVdtW6oty1cEVLokhaMkxdmvg4mzBaBagE+U1AqPHd016o4HwXPSF9h4DK+sitiOny+JgnWFQ
iw0hxzdvm8cdcoanEgbVpVsOe/Ee43jMQcz7r1nRTjCdOc3ge+CBWFdC4NNQtKKspr2t7M7d26ij
DzczLAup0tKwuAiIuOB38mc3ibHKDqFOCqwSMYro5c+3FtRWZKkBdDNi6LLcXCOLjAaXxd2dWLYY
arjnBm0Vpbdzt/B0icdwh6qBMODthHNEm+gjFlVMzs2dp2c9GZN/z8gke/CxxvS0/MbJnA37eOGT
A75YHGUAPGi5vEjLWEEDw3McF5HDP47NhmL3xqoVFRhJsuqRtEakSWXwW7Van8zYWwWo63JKyjUF
5nGGjWmMAJB+xtR2H4axNpFQbBb5KnN/32NqRZeHz0CZU//hrsKR1JDq4vRAasHL7lzJ0jWPB1UC
/OMMDRgZz4wyl8MfvRGyiceHXKTr32VFOTUgUarBQfmTsFH7w2YthH9JN2I7+8zXa4MBEiNyHSWL
dckEaoQMbd+Ly3GZ+BVOcLBFYVS5SW+F5Ze9HcymJ7Gg2xq6hfVBYrYXvgs5Dkt3qqI/x3s/OWG3
4ZlpYfyzU/RatGILJMVw5eZs/sNei7qfEYYbDh4gQIH3lVXgX6a+q/tnfOoxHcG4qi7nTedIlJhB
C6tAozirtD6BaRZQupujEklf/q/0FbG/h09lk1PTEuwpVNuOj3YZKHAdfLBuzvAY9o1LFi3xX91s
Z6YffowI0EY9YSDob3lCivp83z0KPKb05jmkW5VwfWjX4pPl6S0AhpnMcwU6azy2c46CPjT2tLe9
xmPsc0KwS8jf9JlC/cxqrTvNYICqvvdKsO+eCgj/bsAdR3YD71uwOLz0wInNP/tx9UKzH/byWpED
jU0ahWzHFUnc0ozYaHDXn3/oABNZwbX3sJZgeFDKRSs47I2ZTWFt0x2MhQHgq+bhOMCuXRTrp1IZ
axUSfZGIArFyN/Uzya7guHFe/afNJ3PVKLRVQxKHxK+qRW4hdnKTKYSOoDj6/ZcsPEJfTFewD1Y3
QMA9iw4C1K0KzJDM+Hn8BCCu94jEeNIToTCxP9tq6bAd0eTKSkCoxYwR5l7QlZgkc8gbQqqcczDG
VNqZKntrVnZLFthSuri0WFjy/8KbHNqg9nqP17IfphQ2MmUKjlyZgsTd2JwXdZJKRtFNMaVNzPAz
ZK6OPTSS/sW1iVjQSeoR37vFcnElLeDMWwlfXeQOnP3UPSW9ktmRJYdHAnp0G8+3d0hxOCF5wqIk
CNle/cb25x3to64oyVpdP2fsPPl40mv6oNg8EZOr0FFy74YHYxDLcXoGoUYPajeEODqGCT2uRy+o
29IlBOt7y2BZp5/6n7aHY4xAHhM6g+JvqhWoDPeiSpF25sKvjqvpnpUr7cpu4M+HJ8WUFSMTMnhZ
rZkGmn4mdfl6byLjS5isTjIhh6yocNsvUSAv+sTMVnVws4qOs8t7cELC3y130+uZwmL/vNaFr1Nk
mrLmWBwtXXsqB23/cXKO2s+FCu/eznUTKuf33WGhUBtCAvN16AUfas+zDsFxzbaisl9/B2lqrOWw
H+LOqA8PabXdkso/bKCQS7KI7MmW7dfsSKivrH3cS2IUyj454Qfto2aW5HrK1L3fl2vNhaVRiiPP
RQ0x8K3kWpwtESpPhDxW3aCT0Bbzc/Axq8fDK3WRKEKx3uArY6w9vkOZpLATaGeJETlyFUgdoy/3
2lA1rOfO9+YR4dVHF+RsVueMW+Sjq13xZ7X3iA0jJw3q3oq0AL+ecy0udqZutXdh8y/W9BFySBb5
b1qNS4z6UEsNPqfqJyCSTP2yKZfVVIvvR4oXy3UXV8sCRYNG/SGq5iWzOfOcl2jvKgptWbw3cq5L
N3tZNUYl8cmMvQzWtJW51sNLblWql9BFxMmwcPFzT9qNtG/dppkbse/9ldNSN8L/02ruymWfk2+j
2VBz/QmrLAoC5bSX5L2Yp3qiUk7U7NiA5KOXgGslwg8H1HLZicgF0kIJZFojYke61eBu5KpSR2HA
RhUTgqz5HP9Cgd9eArcrbIoWWNAQf7YjMN8gWja/0pgNW+r3LSOfW415TyD+yzgci7eXGu8rT1Fz
8Zd2xjUtGgPcou5b1blddokpEV1QCyGL4MIedMXU4cUBeFAFYmyngMhWrXNM0o0PkRJJubOYljWZ
w23Ug7GjZ4IuMpwNulWRfBvhAyMh/ktxGcKIuh7D93b7VwP7XTyOqgy1vqXiRwXrnOfNRCUUuXwS
MXJjlXytBVQqWJj7ydM7bTMjDeRFeE3jiFixvWFabRctNkfyWvklp18T10LNvBQ4usSkP/VZJxNA
fmmVDZOC+v+brtQiIWA4oPnOZyVRCBCiC2isEJP5oRbKuekvZEMHxn+Hebxz9CtNGmM3qbFs2YJm
w5qbtK7mZweJFAwvO/X50SvJtMCA1G0mXRN6JEtRXa4hgY42XsukzdWgq0slgcT6N69mt6CnYl80
EhxLoDZqkhvycuun2gykYdc6wOIEm1OEtG+E55ZjDTbykJjEZLp21q9uKjzGUbHq6ac9cpFriLPa
7rd+QCh0PkOmsngCdnuZ52ARlYq8ETRt/h2e718sgkRJVxBZSLH3l8jBAW8efLU7KAViUlMfIWzg
qhDpEubMy7Odgkvx+i9o43ucdHz8O3JUJvywn2l+WPAcoNIoopdSOqbq7TbuPuI+kFlgLaj7RYGc
E4q5th51rGjMSkOt82oeJdzGt+niSfrbyWuqfRc3WRPmMzLrIoXNtxXhyVKrnDyf4Xz5oYJnxuY3
W7qBSQMxpwPbrlITBm3c+A7RkMMgp6ueVlpiryZ2KlCT4EeO+Ulr1WnFTuPC4idNeB6UnaQ1S5ZY
8raAzFW2U4cJtt2qLPoG7wEWGmkDAgW1GJPJkVuUNyUR109igIZ9fo7YDREsOdFLEX35ujy8H63w
Gsi4l/hiM6Q25irgjSz47ZAmu0ZfJQRUy03sdmOUMYAN5SSj5ASk2QwjAQ7tb7434rF1MWgBLzzJ
gW/lTzd3Cred7Pcecq/1FC1eplrm59yMMc2zHlfxBB4RjX/qrkW0nbb7zAGMZoHqtvY04q/FyvMd
trBpSyZcynqHeMuq/F/NrYifd5fGpI3rSWmYEIg5VL1ae1koB4AmjvZUkvkWH4dW4Kdd+IKcTqW1
8GCUN4sSyh7EhHzeIiIYqi4uEZ55tZUYmxhrO3l9nSa3Z6GEPeOa/vv9gYTVRnpwbeynJLgyCqRe
251tFNRHv113A1l8gth+UQHWVrCn0P2PU70ztMvXPUXUHy82GPO8G5KVtasWKmjQPb96eeaU5WNw
BKj0fZYXVHb1rrGwbLESysRQZrWiirQ3SxVFmawre25C0pCA2ClYfSbOqGhvZPcA0awWT8cD0WSZ
XyBpvcwBAx0G5JSpdXNGBw4ZBqNTU6JNxYhRb4blaEnpdP1GXk4rBSY3IFV/kk2D//HfsWmQDEI7
ql4TcI19VhG6HBzPv2CBxppbl0QrKoYE0+TspFczjqBQIvxM772aZ+FkBEaPIP8pdbiqKm0VGKQo
e1947Oa8loL0B+FXdR2nVC2Oj79xb/eLAspCImBaw8qR5o0PE4QcD3I25RfwUc557jFt9GFzVak7
hTVlF1TKjsK9LXkP/KUQr1qJ7HpbkUaVHXop/1U/hDuhBSMVuOeHtGYdk0Tk/PenI2Pdst8LhEcb
1RaxzKEmp6GUEAGvPTb9eU5amipwZevXg2caSVyCltYy+QkTym71FjbfwmImEJZpn3g5HUwMCXSg
q1TW/aYS0kc4Yr5erHchsHdE8Z/A5YN0iXk3u8g7llc2nElCt8J5ysYxuGuwjj0Jma7tqmpUTfrc
LVCJco4ivFjUd1qt5l8RcNmShYY29xb8Q7Gdf1kJtpDOVG0AOa0iLwCNZFDH6ThRDoC15ESBHWMd
RtR+qBI1AKlPOYjXjyyHipMvqHufRtcgltHKMgyIqKzP5xJRw71LllP3AwLGBTUcBIUACxuRcJuQ
2t6PIIojFF1ZSGw7UcW0jh/Cp36BjJoqtEyfetIQAlYUFFJnaMLm1dPfqI2Dx+0jOcxJQg9t2lHL
mESLHIsYlASQOgLyNpr/CyCeD1CRc//EoNLb2gj7Ai8ClhFmHQfDMX/Q4XEpHun5vqy0SRox0FDA
0U+XTmJ4qG4LL623H7SFe3C/1Jtjcz0TMmeYm4dlIxp2i1e/X6rG0SKtHONSI5FwAIii963LyaWy
dMmTGMpMmTDBQd8jE1JSOEiJ8aAjr2ANYyObxW8jNc6AwsLc93KXgGk8afzjibnB8wCFT0s1K4CU
7Gly2Me2iSIoqXSESdVIMopgCurbb3ZSaFHXSbO0Rld/qjOcVdXAyLMi2LqgkRLmJ27e9Hq4JLh3
gEauGJ548rj5M5ScsdPz1bRv9ra/7wG85zMBOGazrAxNZqTnNBcbvEtTdgn6exnz9w7fGsh/0TbY
rCP9uhGQb0tq0qt53rINrZ/y/rM10CigNSJ27enDFZWdkqiH2Lfr8mePlpIzgWTu96tGspCM/Ouq
/oFw2pFXIoZYa7fPZcR7UPRc5fAZszfLhylLLRxH88BaqhKlJ8MgAYiXrkHV8Yy4bbQ7F43AwqkM
HXSUnZjz5Kew6xhe6X9Dof+6K6RR2MZQoSS7+i9iPpg2beoK/+8K2NkgqAayZ+BmGoYx9yUqCQET
Xk7Hl3qOkdFmT7bkFXv608KX6uTzPX7GkVn72ABne+vbGQ8na8ROZeQL6nT3ys9Khyg72kj24lP+
8JrmNxkz5GQxZPZTqd8d3PkNdk8vtoqD7EKGwLu3oOT0rAbFHeiR59/af1etQJdHlIBlP/6vJGVh
TbW3eSc3T0L60uFVx79MY72X1K969eBsrboFVVOAbSqlN7a6nuWpnuCsa7Qp9CF9KlYxsnijJTJU
tMV3IYXDOUkeNNTC1DLFh7ONAfjfxMJBVYxhv+OC5oXTK1A0YCrLa+Xj6mo+QMmiBm6TuI+s7Fwa
zezXINevGHtWZeQZR4LajAKwzlnky0Q/zy5x5Nzkj3yPUFluvmd6g9CVou5fOxOkFeb+mbaAaZ1g
1r90PkSyjzLoZ2DYNVPkEiPn0QAPFlW13JCLLRet7MsgDg+UdW0KlGPQh2KOFEH3KpTUNiAvir0X
I8fK3FxHF9HgBOKRfasfKPF3IiorRuUDctDoJujSgTpxXdJjCBACmVba6K4yffFb736X3zo9Pksj
ZoarzpqxDtWOCc4/Fn1c3thqVoIyR7lB6O8IUOQPnH/BfbWEed0j2PHGEn4RBpl5BIQ8obzC7U6B
Z8jnWFukjW21prYdgvwm3NE/668pOm3mj+ApwQl+tl3m4tfBU0lsgFLo3BE+E4uKZ5W7W2FvC61Z
EyTxhLkZKUjP/PvMlv8SZuKoB/TWqVtSvmhUi/O+9x1GC/hCD5FYoG5iRxSuvzd1UM11vTn7O4XM
9dwk4fFFLvW3UcombTKz7xWbipj8f2Nf4Hh5AAQ1J22E3UoG6Gxln69KietKz2abqcQC/j0hNa1m
hRvaqnOebaNfj1lhZO8xUFIq/F14FL8uKYfBs0v9bBGUaGGCdyzNqlPILcqkcM3v3R5IAiIUKyYR
tECLvytbNN+A1PYxXXmgS76TEvNatw6O2WE6nf9z0qnXclMRopGAY+PPTzw4oyQFFw4ieySXo9/F
Tbq04Nn52o0LniiJk4ZDMaklP/27rvA3YjMp1Rlf+Jxo6EjT7uRYZ9cT5khLudjakDWPkFpE5v90
0Fo2gby8OmBIH+xr+TaiuME5nzHWRfXYDGti8mLd4hldubGySmLI33OLUDGAbzM1DiDoy3Bl7vG2
0hxrv4K7joumDj2UeUwfbVBhkj1c6AbI6fHUDR6S2AU01QANgsFxf0TAT8bMF/p8/C5TCyyaysj0
oBeq/wYkA1bdW0XqeQ4HHAPddHYB9HIi1B54UBShvtpHOfjHy9wQrYjvOLIL6uPIFXZhMGnoDTLB
o9qmKlId9gzuSwgcAUlNjBbE4Imj9+P4V6BPC/zu7zsAMqTxxq7fFZxhSCLBKdusHNv+QWTYsGBr
LCFUMD05Qioib3NzXDRHYCuyKr1vCnMen1LKNPkndwGsD5zOLYwEAHR3VrI7Rk3N4Bt1It//RBLj
w3yCT71JkBJKH4uTIuPm
`pragma protect end_protected
