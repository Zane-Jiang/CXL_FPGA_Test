`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
EAn20iKQ5um2jZDzcsZmpjDqASTa2mpGlFgch3NVxyr7tpFXSX8XmidWV2epi/SL
V0naQFhQ/oIlaihnBkSVWmduCf+3xBGyiq7mCoGxzlG8tcelf7DCaelnmcBhb10R
rLPcM8Foaw1bPSgfRwFA477MC1aYkxsvNrwUyw1YUwE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8592), data_block
wUrvC+kEGXhsZuOfIaKk7IX0gBqCSHvkS08bl5QxHGpwUB/x9ii2lB2op0o/64+L
WzGdEJoMSUEnBBb0GNbJ3tfr9RQUBdH59nVPk4P6COkerJZveEvpsnN1o9yEdyrJ
YfH3mbUCC+3f35AL/7ZyDJHklE2Fs4tD1CcAqsexMH5QT3WNFNQzZ5yIdQVAvzPH
XrO57XHsX6mG8P1TQV+RjkpppHFchFoA5M1qVZ5rbqBO1SkXqTm46SVoyHL2haBd
wNnPHqix3aLdgekRBx2/qns0IHJFNtBgZ3D3r08BzKFOp3K8IJgU9Dzjx7r96PAY
PYvJdAuJO4JQzYrwXXaMpjaZyEMp1/tbMgUvotKacJ/55aiRin2GZMJ0l+xY/uOJ
QC0EwuLhFHUsz7tJuBfwcJBBuNP5Jn3VdyJv106qokLtJIOvmXBWywNz5lrWlPoV
7cngALpbhtTbC0rYKL8rey3uMYmX4ucEF1II0SfUqhCc57KW2VoEdx3NMRrq5/iW
2idkkvEgS+46bR6GqbQQxR4mKQaViITX7wrAIW8+pB+ghfHynWMkOyFlSBqmehYW
tmM3uFKeQ93vzKbRWnxPb1YqIkjHFGWNAPs+XdWLp9TXlEChW4FgygC1sdH8M5VN
zHmlZc/Fowe7TqjOV9E0zE+1FpsBHOrQQjDvWqG/t9u5jVwGRoQYdv3Jori8iqJ7
7qXVukMl1xoE6chOZ1xmcm7Z4mDPcVfSlDcAu1SlXys+EAswsv6K+738X3niY8X4
RG7DHb3kommu4Up8G9Dfo4p5VsVd5ULSVOfT/f5gZ02MeaoNXYfxBkSuf0FRupiZ
Pj7DOv8ZnOl81sHgdWmp4EFUK4hLEfFU7a8Lm0Fz90nQLsNnItKuGeoTTdZXLlhF
hkbbMzEfxATrB70L8BdooM+leNWuLD4Z69G57MFDIZKwj1zPFwMrKPHCVC3xYvBZ
CRKMMOneRkrRDE9zBSAP30PjtTuhJDrJa6vc8l8wQfZO2II8DAeMF2lw6knwuM8b
kr8FBUcIz0EUZBg8sO0C9mnaXEEP50EeNERYVG0GrANlqGKZ2AQTl9gyTFtZFfxJ
C9ROCIlSWHAg+5jRMR+rN6EVl9B3D0kztGtvQmP68XYDOIEtBp7HOXXOoSBAjZU6
H285Ny8JExg16TC6IM0nLUGS5Ff4jtvXqa93efUMViI3elAESr2Y70hYf9qKtOQb
GBycIHPlUFEfrHW0FLegDw26bEeoeZmFGSMfzUezeDIL9xogGrA7lvo8C3QtAgwb
NVFniwqnL3jp8Tg3kXPZtEIwIVinYO7gRqqIp5CHUDgKuyzd3+StqcbzgqHp63cU
Bqasvew70Yr17P+Y5jTU1enoxN8EbEgq7p0fYq0EnQIkm4ZXHC8x5HqQC6SwG5/d
7OuYmUjDdW87jDGFurmFm+FrWE6SSdw7nUoO7Jww+/cknH1QE5S+7RM2gwtjumnh
hbQ0I8/bGm/q2xNKH1d14EUye8OeaBazsxQ312AVX9CCetF+hHbA8PLI0JMp4qpG
mfUp9OrmvLUmIQ1ge22JsQNmpb3U4DSNhvdS1SVynflD+xlPyyDNDWHEuPfuGZe+
nQ9iKGD+wdWbySVn7b3CRQqGZ1Yg2Dw5KQiK3wpVBzGhRso4hj53sQPfn7oFalKC
Je91KH3JsXUhGpyt3JYn9UBgvGrbNOMARhOtFEJdbtD/pcTVh3ROnwGXN35mNzbQ
Bu1UCe282xiPmp+hcroyZwe05ExnAUTzMNLvo7ttsk1wVhpHg5e8+yVDWsYyiuh0
fcKCvROCNHH+5DyZc6yLM/iFWxGjgPP5UWndNJ9qnNKQ/oijzm80ZwqERI58ZvsF
xiU0PF3v02CKeGucpY70sGkfu6z+dUG8vFC9EllZCz1cvU8nZbXN7nKTZcsGqMBE
1R2OhkYHp73eqlNe9dqNPAgS/QupAYej8rtLjNS6r1AMgQ8rLuhMRm1yIqS/1fso
L4Rb0mUxwHIe82HkX3Y/D3RlmAVFR5hGDKRV099a9xBGmVk76a06iz2U7y2XSGmb
X1kuEDY1gt/GxSYVDluuAK9f9OvsIHaxw28E/YkrL9m6AILRWywG/pgXs8kNXSXO
MW9+8p7J+7yKT4uPp/S6nXVjt9lzX4yCnc0SbU/01V/5NZvQS2f91NDmIDB1Ad/4
NJDFpmQQwF5/okV4sXpmw8/EgQDpd2fSTB42tGMCcIvD4Gm3nlNJ5Bh3WNwiNHfh
VVPiOu8PmPfcxF+eEXbOOYjAv094EdmBaVnKR5Mb+BYGHD5TybchC5CmizjBIF91
julwBVddjIWQzRLDPxsyodzr0ufL6jS21MQ6ZyYu33bjASrRBfKMuinRt2BppokA
v3JsVSMXE1JW6nKW5FnyXJ4RQtC3FH/ChHOh/hI2MfQpVsUOhDiHDSw7bAAnOTgJ
FhJTB8RC8NfNb1WgrABdTiYyjY+LkSlqBnHix4P6xugC6eoM1xOBCyv7qo8jU6ZX
qW1HLe+NriX2zO/zxdBI9faZCBAyHEMeu402TWm7INxx2sJGv1+jrdbwj6cAk6jj
5kbhHKuhoNZgFtSLbOhTGIMNcbGGy8Hvnyj9n7PlXHFjw5lfj83eZJokZ9cEd+iV
b8vF7XXuKePS0hWfLwGMlvzprqPSrTMW1fcOVTpDJ2aGZFfPaTJFrHpTjgCH7FNh
jYoG9hSxTL4GiTIejQavTb/xgEar6tFAsvXRARufWN1KKR66zESrl/xax4H8TjwU
OGkIw3yF2k9T6QjpPiHMUYkQ5fQQqCYU2ak9qJoYDvJeZaOx8H3LErtvlUeyBWF2
NACv1GKTh2+TFKJP0pqS7OFsA0e3Iq9XaN3mqeiksrcA44ablQQDYvp16NlzZ1gv
cBYNStgABl8uB01uapEIxevRU1mFzB3yC4lhFgy8JXN/OKuPTW1MTxCh+dxNjW43
ylL6xFV4TodEJJUERdH8tTSPyOpTgSCKyfg8skjk+Ya4j4WosarlKpa/sTqp/AtH
A8aX4TZfzJMkjLorrMbcLPiGaE8F4dimZuFoU3JEO1Kf3+3VHolMS8vOKbnlXKHT
HYvwXrWDmZ0LH7BuZfNpbdbcmw3IuERHVgvLRit3zYr4TGakrEQfBJHt2uXkTVK9
wPy/VVT7ZTHVStFl9n1KXgWVxqmY+0YxtsYJ9WT3BUUXaNgw0GG5Js+pBykF91KT
STGgiw0a7nlW2oilB4hrZkf7qfwRh2erBWITs5iyfWCvc5gH8/TKPROCfGQPEDEC
mOxiae0FTB3StZ8SNReDtbXkssx+OH15G8op673oNK+ujIPsC30vvEWxijU2OZXZ
X2wisZToyyXofaxvLrJjS239mp7GpJAqyynN2Mv65eMVOCcASqdKT49Gu6kkY38n
jlnnOvCwO1hh39CGPFG+aXbIa8Z5Hdbg+CYRCbCf3iT2cpdFaKFFt40vIUWkcJRn
MYw/cuFnHOPtczE7+xqpMKiiE3S3W7wdJhcWVEE/sRJhIeHTi/iJE4qokE2F3+1a
7eu7xdCYAfHNAUaZiaZeaKHiBUAbR3C8NF73NQqWE5pX0E8adD3DcBylf3qpzR9R
2NbbxPDPZ8eMuYGobUfc4vJZ9VFfkcxrWDTD2oZWquTO/gzqBdvq/W3ynxM6TO20
rLN96l5HxALqJAqu4gQIpmByTeKvqgQNSEofFM+shvoXbDxpEb3R0H6jksFOm6ej
3ECuwjqiC8AhtNR16fIt/JHctMfstfBnjdbjTjpB0R7RoNf/cwK7IiQtWOpUA9E+
/NLG6ff4rLpCbqd++dJHvPLgxB/kc3v3QAN00vuwXdZwCFBx2QS/xpga3lCRYGwU
igLqGQ3MODmK6/uO7Anvma2xwrVc1ljFWFfUpe4SZzO4kQKikKzrZhCnpli4469L
ClAxUG70eEUOCNf7z9gz/4Yj+LiV0MlIllXYq8nMDcOCFYo/JM5hFcRzSq2bTEDj
4zX86iW0UVcxfksC4I4JpwWKhLgJAvDY3b+zP5LhLF0Rtp0+sAf2nYMVYeNsgHn9
w/RYIIWsTgywuGATEU54yDDFQjbPFESDXyCGY2aV+G8TiGh3D1XbsQV4QLfI7JHl
/yMBoMgG333C7AjLIanCwL2S/TvDSmjWmnCZu0OxDZDlBWka31FrxFCGo+3fMPe3
gC9/mSKfQnvmf8mr2B4OX8KfYYARyYWtgR2LBUmzvemQb8C3gAfxt3ei1LdJOp2g
qbWVIaFyJ0phTJouwH9D9btaA3nGSI/X+HOkkbwFAd1iD7RLZyhQRkUFyN04HleT
xvyseJnY33pi+GFj+mU7jCQPv/wye6x+6p+tZIgXzUfBh7uJvbEiSZJKyiH/KxSD
TNAGGrg3MXk0s4wZw5A1BSpiRNrQVufNt7OXlkNhcWe5UgSTKlzhcC7Xob/WXVwa
K5XAhsiLA9tzYq8BvzMZ6DdkxRJ43FhXe3/i/r5h63rtdqy4BpLyUChbIMBoH8yb
6PzF/6ItWHPLmmTqoYd1V8MNCdDSTl2txzwQRIQGzq7aNYYuq0JYnCy4z5Fp8jzT
vR8SApRQ9o70MrXa9IlSxJBelj+V9Cl0ddVU9S63ss0YVF3JMmFyh2sxG9rzdBgz
nqTkJ9xlxRnd4WMR6bylBNt1c+jXI9l2lcY/UX1g0STgPNU58H/KksxOqrmX7P46
uOyedbjK+f3b6qz0LUgGaQiAUiVGV8k56KGgqtky422REYpjNzDzOmUhy/unQzXT
BNqWvT7uhyhyIhDcgb1c9F5CFmCl1jqOf1c+JeUEYmugTQUsmh78hh/PD9Y2zyld
5HN0yLfhhMYt0gTY0phaCuQficBkuw2jwp2l0zngY03jJ5SYWfiQ4vWWYtTo8WW+
ZQm7rB3tlV3XD8gWu0N5W79SuMGEFJsbFWZKVWZkqGeE6vu7kwCaeb7Kv6SXe7sC
6tiluIS5LdXzCR8RSiutTN0Hu/3nlnIBQ6dtICR5uT2EShRQBqpO0RRRuplqiDOy
I1QYmT5SLbjxHaCkZ1TAm2ln5LWOCE70hDJl9qDfos8CltifzDpxKg0dotftGg/F
CdDb0tUwU+v/L19o0k7BdO/yVZLj8d9BUjvJjrwUoeNNgJHLcTgEjMI5yRK6ufw4
9wS3a+lDJwjTvPoZ7eGtkyx3rzSyQIWBnKRBxc8U5DgmFEndsjTa5GPqB5C0cekF
vy88SUwT66+a6f15DTriuG5ga2m42v4l75ncG2rXjXVhbVv4W4LsCXiC2F/PDWKk
xOJuq6MgA6VuWPxsWowLEaffoQrFamzb2zVVyBalh8tGq+HOdq3mV37KohKTneFa
ej2qYJbTgEKa23yludW63nmlRM1iHuMyXxbyj8PTr4PsA2ZEqVdbG2usheLDt/nC
TKVL3uhTYYYtzF5qcmp0POFAqoyE94NHYq4LjIFeJ3eGQRl8SNTyqMo3TYJy/OEY
wcKl4AWvPGI/Le/wDMIjZuCEzTPTrVzMQzgG5ryQXQoJJOkSKM6Yb19vYl9IEq+T
eXiOKiyalCqgzh41cN7Koy7ZwJdfVG+zZfRBeOSRUOCHARly2LDbp9fn1toezjMh
4jZUvLYFaVtySvLXCvBg/H6DHOfSohTrZyYzz5alrTESeWe4wG2i1lM99VBk4St5
GUm5CzRFCzNAA+Vp/xcIf3r6Ixebry3QmaK0eUlsXsFMgQkt/SchMHxrUNaYHQqy
Pd+Tem4BKG03KnUzalcVzIujiw1i3LRCipwRWCqkAtL1QucME9PRdycZOm2ip9nX
7NCWy9Lo5RPtSrX4Fv297Jq/UXVSd85v7YSbz/FLQx4slUGnxtumCAO9PeG1eoZb
+R1ciLVoJEI1z6Q54qAQFQHFWI2ts4vuhfkf5o4RbXOXdz5r+1bf7s+ks90y2B8G
M/uKmUSqg9cVOjRX6yJl6e3yr6p5b+UZ0j/HvEKyt0bsSna5eKOL9t96vO3G7/Lo
iYPX+Nubv4lcrCNlxEEtepsBffXJSiktbytXnAU5WltpLjPrYd9Y6SVjLiCouYI9
dBqMHvRAQrf7mscQlb9xQwRRBAPMdkHPSiwL0pNWUN9shtYHiKS1ElQ2qSizTAmu
ud0ybwjxtw0W9bHUjaqypVOU/yr6crqogir76zzqBrcWkiwOZgSeMOyfZD19IIbn
q39CPA1oQfTQyh0fJi5hMOWm5w2BmekbhSoLGrlCc5BXHn8tpXUhHB0pjbYjzm2g
0JfN4TeyLnQd0QhASsgwkysFHDbkZ66KK9Fe6Nlh8W2wmeaCoITAdjEOsiI1JpeG
9/3vDN5C0HjcQ1lXOwPxvjE9MYLGMlSDa/a/RHPIDEk6LzEWyoPe5QIVK54z+8MO
LeSoxkztVTiR8GT4ZfJlx/qgb/c195P/cb/ThofVX9stySuN6k3j8OYmjffisVFD
AXc2BEQ8dmmjyDhJ9ZBKb8vYZ1iK6uJ/0Aa2c4lw+GMRWNWz+SPebeCh3Qd6lBb7
OQYsiq7wIqq1aidmrpX9HwkujXtAJskQXNFMJmRBsGGU0LbUdY3Sa321GX0YiYu9
dco0+/Iv68hF4KnLmOmG04Kvk9B3Z623RG14KdaGcjYx0XSDoqc9V2MMrRxN/EMF
CZc1IOENeqCMh2Y6Fu88s0z/cjDNakQSS/6oRkusBOvsUpPydV6Hatad0SISULJ2
vAg+H7hdDkfEyV4o8wV4McWI1PnSLhDtKakPyFg/yGUSXpDEuZJhyG30SBIuj8VZ
i57wdx0nJbT6dXob0XfV1daA7A7jyW7gbYwg2VfR6M7PfD3UeMLs7jKxnar4hnsB
rmpEqsEgo+kgbnD0bDzw+d1WyPGyKk44U09mJE7G7Exigg9C5Lj3w6V8ctm+lGeD
As1SKrVxVtD4W/WvbD5RlroJYP2mAJIJX2Tz0gqTkn7SNem14P8rsdev0pTEpHq4
tT+RNc9QeOag4Dn5QqIyjlb/pck7epwcw6FEDvlaLDa/EneG2wm0zQR2yCT1fe2N
gYibBJqIIsgmGfCAQzQ7fDeToPNzDDsUEBNuzoN2aF1eVUXkYCpLdluOzUlX8xDo
/QxRYn8lZ1nhZlkby7M7ZRbSoDm0rWnRM4wwtaJOHfZzrsU4iXujazTfPjshxcB1
7jw/5u7vxzHOcyay1/FY98cVvOQpjt97+iE6kFG68LkKEDxa+ErkJqGNR+mbenDM
6HShnDyHtuTO34sirAeqxBM7sL/k2jsDLYasYnFFRmc9Y8vLoQ9s59PQlru8HqGj
ahZmlW/S0/2jw46ZQBjjcgqBPOMN2C9xvsYMjinN3dwFqBikHYujGoar68q5NB4q
EFdjSxOxkECN9MaRWxGbsGBCaHnqyo0OTmZIqmGR9P5y2ChoOloXfWJIYCsMWZNM
jXvBxvx4OBc+tn2xYjxz/z/TWCafWFOi47PmSjOuAmgHSLW/2SUFCFm5vSvODFOS
QS8QYoCqxBG/F2qR0oDE/qJGEUhU6zqpC7X+UMIZFflp94phrjR5JrlEk0RoBYIS
Q36imsVJEbmzrtKc7k7VmGdXiLfktBE11MXtFekRFfL4ZAXVL+LO5UdfkCPhBSg5
vTy1r9m3g9sf1uNv4uW6olVNzOKkBcLhhdeZ3MCb49hMaigdnGFNuXQBgc18i8zo
F98ZfwzUqnCWtHnDJkdY4DO5Os3JqiL2m2Y/XpgIdphtinA2cTw8hN6q9IqTh0O5
wyaSMpCgeVQNYgWJTAzlAxVevAqeOrdwW1Q93lfMe2Ryyg/U7V/qS9607EagmhO0
T5P4TACZqj2zGbDhW3qwLMNogZjU1AzcwTsxbry1l7xyraPCuNjiy/tnceJb7prg
Cn6cwimRNDY8iAbbUfk3SKI0Hi25PujteUb17nS/cgFkCPN8NOko9YScz1dwKLvJ
mIqApW4srLT34LLxUoHe2NV04pDdSapHT+CICES2sstbJiMc4MtSWyFVM9wSdoYL
WXEzVuL2h6+mgfnnKqL571UdBUDIcOurlBHDaGGckm/OMBN+7vw7PrBfHUnH4XXd
qfEjmIS+iPiSNNuLclOa9uyicfTPqOFp575LuKD303cD/APXJeiyOXEYGyTG3Sq3
FgKIqP85wxEx5OjyHNxeZ+qNCKKnyVYshQkdMXR/D/DQdvUl3GarASlAP/k8oLVB
eNtnEWTfBl8xAhDkVpy4bBjdDuUr5VaCnMB2/o9XNcgUXjWFsR5yzPw3xLPdDxJA
3gKkoMCiVPGtGU5fKbVJBloCNcjECGf8eHC6twcJU/VyE8xYLackKihTIPxZGFgQ
K/hK7FQqIIkMCL6YqFh+Ve7XzqCeROsTmDmhZRdNAAjYhAkkqONRvP73gV17M5G1
R8gueJtOxGccJkdgbdgErZD2WZikfv7x1WSJI+OEQtuPRRXnw/aEqF19a046Fh9C
JwkKv8Z0fWLi6w1EGpgTa/HmruqfQZ533b3lZCnpXOcU1gRqbLzXG7guP/1vy7JF
wWrliHeedYA+dn3yi/1dkyhXl1Nvqv1kGT1g9538XqvjVe2Avb+7iKqzO4JQvzgO
5lEGyxfymhhrR8jSQ4TBEUJ/zA8UpEIbiw+lzFO+lloa19Cuwk25PXHrGJ9XgEO5
sISurlqKrDLVy4owuBngxkeNkCj30taS235OlbCeRt6WpzbINWC/8MLHbr3Y5sbu
Lw4aExj6hZ3k6xtPDGX8ebKQXrRSI3M571rHWaPnL5iWBEXrVpUOZRjSOKIv4Sug
j4Tky5NMy1H4+8hw+/T7I78hsgY0MJbt0tNTTvzt+wsK9z7iEaGkYnxj5asXBcrx
rL+tLMmvzvoj7iwwNPE1MlHV3qLdceDSG83LZTeVG0G1kCKmUZwwv0SUoPqMdSnr
veKXPr4LjGrP+HZz87m71pNsV1BGsrA/UAG4wtuW+n/UuBstTWgD3cJPFxdxTjeJ
JJq+i921apFOt+f3Gpq/xMMIivAaD+ZRC20wd/BiwivLvjk+Jffk2+HxvUnLNkg7
RWPeEixHtuqAn06byidpq3amG1SXmWOicqRJKgYif6UB6vrhSNauxUZLpDv0Wao0
6OG6MZ0abPwpMZQTt9vmmdtA/Ec8kCmRFakrhJRp4IC9nhgeRifKDc6dvnJfwQdZ
+afHIeEPBHrPgpkMv1npBtzfPBsrsQVWxyblzJYkAIaQMMLr3ltJBMSlSLSFPx8e
Y918gJQQVU5E3rLx/XicYGMc7Q1iGwF/JfRGyqedV/SAHzbepAomjtkNxYU7zwjx
lrTmIh/Oe5+VQ/8RscSpACnZEoZxBzTvG2YePwBcfj5l07tfhopPFJ40aXvAaurO
hDxSz8scadIo4iL/Ua7hBgokBwxXV5q+JW2sBn0qMC50RxaPTfRef1k9BxXox+2k
gp3ITMSBhipyq7r2iv6qVxdsaLFUr2E2+gDKXhNIMAPXAOF1BqP1J1RZfaWT0wjF
ri+R3aBwtvmLaIoUNNw9DU1GHh8jUlfQiIlOM69FesMPetfqmFa8rWsD33wJV75R
gA9l2tDgRdpKe3mkwHFhP67vOZVh+kO+FNnQAMIUG5V2M6C1WKsb7dMFlFP4WRUa
1M+uMYafZNvhayHlqbj+3/vmFaxSK3nG896YasuaUcewFc60Erwf8a4N8akE5VLk
kXnutZGnK+K9icnTfpsExY9rW3c6nqfUsnAT7KwnKUSohByLGhKiiDo8SuWbaw/m
wZv6gbHOXtfJ1rRMZgSmSvPi1tkgXGbCPLv1EDQFjlTvvJxoe/UrLLaQvrAN60UA
8lGjYGCJW4aNG4oD0qKXc9bblgeCuPKPg/TFQB+8RrPdL4ZN2oU482yslRGrDwml
oE9LZ04yN0zMimqKn5NFb6/2h2zopnoblW27euv7bYqZCrI+eCxwKOYkcij21/wl
ziNoNbyz1z3CPyJPm1Tj/DIwkA5x8D0AYJTJqw7QflVJPAZRidsKcuz6c/oEqFyy
Omj+Sf1O4nGo9l7DmGjAXUYcBsbBUOBfF5sHKnq3kZ0sJxvaK1qAuS6PpcYZ/93t
7ZGeDeyNGjaSV48XcrUTB3Rri6OWQzY+I7xZ8peztHluT+CacVBz7Qo4BtPpflA3
t28VAIBarHTvarkANOZ+Ir5rrHVsDL8hUxiyIu0/toujs5bnVwHUa9WeVdngS+7D
TfWusbSeJSwF8OTErsFq4tzT2a2H/8hu0L6x1vzDeeI7EJaGEGqhfJ/Wc7QenNy0
DSV4BnYvGHhf0UbFDKyv5iwJMhEtWnawFcKYXKs1I2/nJyC7bc3V3XpPOYKOP1l3
4gEBUfkFnXsRTKJzavmr7hA9N/U3hmhk+qaITRlXKaiJUlWex8JRMA8rlhjXTK59
ScRD5trunmVkKefYa8lv/rLar8AaXHD6x/E67SLQG1HU0kZSeJvm+5t3BZsSvpI5
qM6UDrmUoZbktQWiyPa8oTN2JYe3xlcb80QY/bNDj8PYtmKUPUBpwHoFgqMNiLM+
vicuu8U5rmAWApae5wleBoa18bMoTLmUQRvHaI2DOMY5IXrVqjlgCZL8lphXKxhU
hqEHDyJufaF4ZsoMjPdq0e1zEaFnxZEqMAe7hPZgDyahaNgWfq1ZeH9Vc9AHDLM4
7wJAzf4lFA4AXj3Yw1cYgvWWykv1jr33LgaN3LH4FKQV1IsJ3PfXLmcsS1tKhu/8
r4RPi8WwN0yMTL9Vcu/h9Fk+v6LUFqzCeq2dUq1JkN5aCDaxN6gCCqEZMuGK1hUx
2g6/MovvjoocVQnDbqkPBbH6fmrQv20WzP59HdI9f89M992rHgZ18+ejxWJc2G8/
f9UgLcjNk9PTaIdwpGjhMsliF5uRQ+FGCkYtHkSSxiho9UuXSNDqpJsIfZtJsBlj
KhI0g9LgF8Eq5C51NMb62wFCdKCMKFqKxuoCZtJcF7+KHhqiGJqr8ofqKxuStNRG
QoCAzBS6J3OU2UnjgU5JQ5rQLc1o8M/yZm2kE1GWA8FwXXkvMfVE7sjLchnHhk+y
2rIMGUNyEmIhfXmDHKGYyMUC6DeFMMmIwNmIl6dnTyIKc/O72XKFYBgQ96clO+V9
m7ewB40i8N0DtRuH4ynjQAwT4f36XGv/XAVe/Kpf1qM7golrQ3Fy/cgDd0lc3q+/
rwBbcrtHmka1rK16CaEt0BK64NxDnIE662G6igRSiF4q5NQ7ZrgFYu5Nv2OCgFmN
Ol24RDTOqf4l1zKLQ2c6Thc+2vjuAkU0qA5fm8Yh2OwkBOiBWDhHrtHWI4gd7lmF
vOU6MAEoYkN1AhTzerhOMAgP4+wBpoTBtzbOmwN3CCpnMqTAR9pmE9RkOGDc+wZn
3aXaLJoDoxQYG0aQ73//UofRrhxQ8SPnsKANjLl7kx9taWkAnSTKcWMHk17LO5lU
Xs8V80p+ilsRFNH3+S1zoeYXh88Zv4cgVL6O6alpxD8Z+jjxOKir0D6OsIGQ9Ldp
ZEotEF4IZ4sArp2dO460i4fPC7pzfyV8mqVKnk1jc7lqzvY/x1D5PKiorSSoAifT
`pragma protect end_protected
