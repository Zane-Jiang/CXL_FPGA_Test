// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FMGq+L3kid8lZCnf9uX2aoAP9aEKN2WdlWJyI08ADkPHiWlnIeIbLJNhbP8y
6PdQKaObTLSC6KjC9SrMhtHF7XrSy7VROdpimZZ0crRquTOVWK/VxVnT+hta
2CdyKEXRo/uUMGJ6HEZD7YrOHixaDIO9b0E6TqhBSr3+YLN0u4K/gk/kWCrC
xkVfSZ2KPWZ8iUPpgoqiQCvMA6X1SVrrFCUaX+bEifpftJZP9BUdxF0R3G0e
FgicIe2vLcTOQNcjXL4DlD3Gm0x8hrRFgivu6uqREruOdgIfNJBazs6XT0ad
pt7pwSJ5MtwZF+K/P1zqPQyivlzJBkSbNIBPe6UAhw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TYtjoKCcpd7Evj2UDkIzTZC0fCWos18nZJ7GxiXFinuf8qGYRP272MFWrVEm
dMWrrle4FPydtLnMOqyJCAtU/Uow4WJ3OfWRZ7uZyjxkLK/GMbLntznpmRzt
tOoJt/stCMmIt78u94BTJwiI8a2u6ZK4VfwgIuIiUCzXPAvYI5d34qGGpxG+
BoFa+AMUs4QkUPULdei4XfPR9jr3O+jMjC/0AhBZnfEAmzJAeBHnhbiAgZLa
8sgP4J1Am3pa/pDw9RUYD5AIAjiZjQi5ZeuURCyudoYMOHISuftOBBUFGj0i
xgP4U9J+7xXJ1LaoWkCpYNKKtwpX096coKQWzJbYyw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V18gImo9Dr5aiMBviJAlM0wqqdaHK4J7u27KiWJP5XSmkqSlpHYToXFmnqNY
uB/j1d/iHjxPP/h5tglyvr87LOxC7L0ZZpa1v8Ku9PnhBbD3ClQjiy8SVJIN
iV0KZ4kDuSq1cCajcnQFdE9b6LNJHcVxBSdnjXSfKsblVeQO1GH+KgThJD7M
syl4vaG0JioTNBvBA6xPY+mvbjeFDq59ziCcHHbsvy1RmsQ1JgiXXwEeA9rj
vfHsBka5BjWnzsxp9JNR57hbr4YJEg7lpfVktw8ZqFGpqOwHbxk6CO+KvdNN
GgkGoXb6ppGLn7CiKsexPdP0X5U2OrF7FGFOCseAvg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ilesC1si2dsgaqf3m2LB+4KMakBj4ERziepukxG5zF2EU/jmXqTDX8p5RrzW
AGpWf+3pgLZsfdeu4fQx81LrFFDQmxFiPJLQalXCkK0damHnvjj785bej4vy
n3vBe5glhstNSrFPtBAlBSZPR9j8bDxI7I5vi4ZZax18j+7aOW4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Se2QY2GuHUXPRrlEtYDyszo4xBa9oEBwc7BbbMfPPwuC0vNhkRWn/+pvm1YL
JHZxvJmis/9M1VPdlt9xMhPisAMr7idWhZ7E+UkXJ241Gd3FGXQafrsSpvOR
3YJQBGosr9PBGXiuguXH9VPMv/6COb0s/HQknOlpNiEUJrTDscIL/mOkdX/q
DlRDO2Ejy/77638g2YuGPbV/tKDPtyvya9xcQlFA4Uf63ipbNoiR+HabefXD
oPEtl79NO5pOPZjlP39vMmDv30GEeKfeijCZ0pdS3daZqzcj4L5ULs+lDufr
/8si+prTjKvPZs6Mxv8NO37iLmJu58CPl5UzUSDT+cSJeF7F10sq1stR0hBM
ij6YBLc9s58JWNgybqJiiyD+bNH2TrFtxUSZlvM9ekY0DU3nTgyMprwKhhOS
tAyXcso3RqzmN865+5A72rwNpyJVItsaqmKnyt9U1Tlnqjo0YeA/YfYVUB6k
8/o5PKAsX56qYxSJgIpQhD8KiikRTLoN


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
neH0IjWbAh6l23FMEO0/H8X9lDrhjuO2XD3MFidzD7PtzKlML5ECGeUkXLPP
sjJMvlV3MUN/xSb196X9yhrIQDeX7kZtgnRtLj1Lxf18pB2vZjRmvmIZwJ9X
U2YnIvlyKQkLpC/bCk/9i4b+XL6L4a3yTKR0LahwK7aqnOtvEAY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gwU7tQqioUiaPFKAcV+/mGkeeIJKOemLFgyeaYO+bptXH4y8ZI9Xl+c0go8h
/gB76jiTsZ6xm/ihy8IxmdNLeZOtPbywsyaVsehEH/RjcRoh+gxR9GcxiboT
g3bWFRG1NHTDQt49OETHebTkhq395oKz3/kp8eItBQvEK2vX+M4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1072)
`pragma protect data_block
/PtP83+qNbGif8cwQfr+v4XwQsTtp15IzZDaWfdvCZROhPd7v5gjlkp4PaAx
urH3FUwvD/uIaOrLCLkoCXBps05LduMgGgGQfyk/OSZq0X2u+91+IfIB6+us
ta/93btdBwGxcanMHVWxaguSVyh5BElhaQVoZT33oCe/g8M+yZcRBw7u8BQt
2Gv+hcEjHsmTFJ26wPvu3z90HJ+UG8Q2Z584pi1CQKbSaCwf+V1mq7Ui9vR7
XvdkDB74f9EAYTS8QH0ytKzL5F5FW2yk1RKPVSWxeRH4KzbQIvl6l/NbGp2u
BTXd9a8ZJxKKsRlpWMZth6GZtWnD0gypbFJ94DUwOM7jiyZYPRRkwmLM/Z+u
DkG0nL2ex/OldOPKGPR4UXJRI4C8kpTaohzxRgFEgUOp17CPxuYVLJ7UAwV9
kosgn/UvP4To72jdXs8HSVVwsPmmhz1w73Xb1OSDLU59TockFTOhjg+l6296
nYVlcaO5xW8anIeLHLYiyRHY8os3E48g3PbRSKV4fazOz0I0fRHmPiDPyG33
IfHuzQHm/sXQTQtjckLpqwknMYTCM7gsohpiTcgqdF9xgDTj1ls90RpxEzb/
reLVxophVc0mr//DMgbWExDMy8qZXXbfVzh+qyS4tPIPOqdVhgvZxW8EhvgJ
Cbs3VwulsAhkMu8ml2E9G8HRx1esj4AQcR84d2ohOw1osXbjtV/V+oTlFMXr
wVPXZI0y1xqZdU7AhNpB3Urk054nZ05rUU+ch3bS9NU9zbRoH6vZAgRdRMTv
oCnes/IlQK5mCKk3/ichaWgAtLevYFi3XHM4Sxsdwrs1AdPl8jZ96QVFe9hU
yExoQvdRw+RBZBatvGas6PxJWM4CdZ3BOlW7JmobxauQnwUCHy5xXKJ9sE07
1h5XtPylM14e+Vzt8pL6yTsO/O39QAFIX5kdFrl6IQElPh8YP9d9dILxj8Ra
eGPH4rmRM1FwwFzzcFVf2+Rlw9hz5HOIRl7x1E1eB6RzVhrcBmOWvDRVg08M
rzQK8iiKNuqsAtJ28dyKaQaiq013qOcCDee2hdnyU7tDWMK/mXQl/IQebARe
UXObyyrX7StNdCdemYzVxWkg6+b6KC7XpFZ5r4XZsGvDlJgQhC99Kr7pmCp/
HtViSk9hi8uPkBLviwmUVcdZOguIIaKf/d3bqmP93i5T96663Z8Vx4XVw5KA
EXFUIsUY+GSkzwQAHrRvV5zJ6TYAPdB0NxtOh6HU/pirU2kphDe+y9o2ipPx
NqbuFIVaVELM+xa8XHzJW48gQlm5jJ/LsRXOpcZNgCRVEFZd8NxrWgvMMrfx
ePpcDLjzvbYr2dgs/MepS18T6i0G3rhMqtcNhK/7lXtqZiR896uVe6eqhEIy
FqhCVhEva9jQFqCkMx/KssnOYZ/uJp6fn+AjqB5mDT2PDFl92w==

`pragma protect end_protected
