// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W6AxSY+jVQF8AXQFR4zHE5WYlexiv//ZR+S7cMCVohdS78ggfsuJFkAVGFyu
/tMNky7L+GuBbmyYY6uxO9GifNZcUQRtB/Pw0XAHWwQuL2YmSdozA9rQ7Yz6
vbfl7BQlUNQMhaDCK2UUKvaWRHeML7aT4pmcW+lzfAyJ2fK2jdA4ISmK/yhN
Ffj6GoFtwi9cZm4lYHjx/IipY/JtM+TBeEYjU4YuyUkCZNb0G87IYCIFq1Ti
hyrGp2SlKXzBx0RLqPCEGk4e0BD2IOiZ99sZXxflFYZBoEqzl3BO4MWrQ1zM
D/n9SX85VT2wZCoMbWvBFHpgsasjy8XXNM5m3kYSzg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nGy7qEkZd6uW5mNmEG9e+gojZQESu5unY/YrirfxcwMnLMIP7q4UqSXZ1Hbr
4sy5oIAKtuvmaXRNCJUWULS+YlOwrI2lWHD67QC10GJRbEYJvvQ2bHFBf0Vr
B4R3G4l7YP0TsG7GKoTcsHovG12sJDaNOzPTYOlBY2hJ/VVhsvEAQ4Bp1yxU
nIur+NBchQ8EKb4+gFd/lbTu4tJUeKSZP8c4YCrw2bq6oRXhozHL3c0m8UUi
od3Bmp86VkEJQjlFCBib4HB+/dQvYQbzFLknSkxmS1E5iugQj08xG8a++kWZ
cZH0GspsWxroNVRPn3r6wipLhDpxZ3CnFjPPMHsPHw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gM1cc3aeBi7U/usUcU9twz9whjQWtsaiB5McvGU79ibmLpOm5BVBlRBCCVgI
/T6xF6ss9wVQ9/17JOthKE8Rc1IoB31E8VOPiL44QldDSFfEXzXe3NvFEasS
i90tatD0ZuYcnY7gdzYqaI9YyzyjGL9gFjR0x5aJb3XUvi0cW2X/sLhLKM9j
XASJ4YIRS3EYTmzsO2TD0jcIw7vSaRi/SLKccr6XFah0+nStYTJkzNWz9GYy
9VWKllzfWfCJaAjXr4eJ/g1oHPQ+/CFMe3IzmLQrdYounvSlk/1O8GE0jNoh
P770EYBI7hce2utHQKu8+HexYRuoMQxZ6C729PcxrA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R1rNCblHuUudXfPU9Le6TEIqW2MCcUnhmkdrQdkfhg0jUluPjhDXsvycuWWU
kcE99iDaKGdxvVLiLg73LFU5x31Tl0Vttoc3igAllXXuCi/TLOE14G9yuSmE
BGfIIfeepXU8J4GJ0uhdIC3cA+TOR5CG5IEq424zWCBFKEcsldc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NKZb5wMtI4Bkc/gaj8LUtKA1NTFM+YPxdFOJYoUo9Q6uk9wicA/EFvbqC/iq
nJUInz4Bom70n3ZKpK2CopW2SMDIezl0+2UrUC3H6EvbWkiKEB3ebCu0qOJ/
v/16bf4M/1qoWbDQlZKBrT2zdAQ4zfgV9RsCgoB7/Oa399AliN2hp7yYeiMn
6phWBIRmXw7rDNtwzG9DU2bJJMnaPX4KuWVXgftJecwjMUgUN0bf14/Xki3C
VBb7SI+Ae+mD7eYjU2fJ1KJZMfbHaaGzRrxIO1JbiDPR38wjr2b17W31QXF/
a6LufZ1nZQdmA1Nzgrv9gF3Tq1G1/GrQy0b8AQUSdUjTbt4/xSxbbkmb8VYq
u0OPy4gmLqWvFY+vAWvlYfwX7JwslvFqJhwhWGuqHR5M/UC9svLyl5t2uFbk
cKziSYAxE1AKikGw8sMc61mRbq4eCtjL4aB5r2hwFPjZVETHAk1uh4JRKwSL
2qBDimL5PSjBKpeCUcFivXkZiX3jx/aM


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FZuPnA8BmaZEOWRahpHdDao+oFv0hIssSTA+HtKFtMWcjlaAzha8XL3mivEu
93UoPTmhII1PPZ4J54wZ22ujeWB+oxokXqVzUa3mAJuT5nnkK4FOEudQFGck
g5iOlGSNeuuFc8QrUE/UtxdgusxgAv2YSFK1wQuuTGFPT1FJ+Lo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jVJcsXOeSsTIfv6S53h1wM9l20mNoAgnfL9QfK3Ichv6Eny1kfscgGwYp0Nz
GWW8mKy+oeQ2v6OvKMOnhpahs/Uwl7X1GCTIUSDZKl9U9XbneFJJylVGMy+X
EZ98/h9lDMzV0NhbVuGXLwZkH4zz0eEXvp17ts56zcj1HchgaIw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 84400)
`pragma protect data_block
ylz3Fl0GcXVrwV2XrNMZYsLFm3mbGtt1/8/SJEfyE2swPz8U2Dc+13uPF+1z
9Ii6nL+WpcM5nz+7vHvdYkTu/WY2DWXQHp5xgkVFJ+mDP1gW8SQVnC82vLB7
zT5rotr6+8DumV4U7z2eeAWN4yqqs0OR74G/gXbFYWSQH4OZX0ySCdT7c2kx
NhmAaTMi9XKQsb+FYS78sTa5/iUNytsvdd9m3GnXJBynnMvq6xIp2pn8hSg7
737nlUCgAoeUmirvEiKD54lG4PLw2rPKp7Gh/vAdEdoxesV8anxs96uHscLe
WUfOooXPgopgtLIOBRorPVZLKQgxeNb+AaLkpCD4lVmYyCWBFD7ygRx4dipW
NHxfxtxfCaEyB+aE7F7yufhNpGCcsaGiyNDQGxddJOlJ2r+czajkFCaH8uFx
eydopXD3MRUW3Y5rFbr+AamblPVMJUodQqR7fmU1N+2BDPbA3KwrTvYbzSiH
STWH+IXL/neYInYKGzwWewPN1QQFpWFDiS9WATw8BV/RgcZi7nAEU/PPY0Ru
pEvqihLKrDHrT9bhTSzfvmZai8LBj2wMW/COdwmh0aETNhWbJdQ3q7JfBENj
bpLcStHBqCmlr+oL7Ed3sh/0gD1KjSBf9lKsUorKTo+WbQmW1eCyHxdN3H8j
/4NdG3GcWbIMQ5mgmte3tFo0lUoC36ra/wupdxrv1P5g0JB/zXS4f4zXONBY
ZNXosMZFrvDknA5YlIG+n/Av8IBAB9k+UnG3snALmNxch7nvxUi8F14q5lRZ
qWuQIsgNYondW3cBRtAajhkzTae+pffmtWt5cH+p9wholaM6wSdzZnGlH2h1
raB3CTWxUjGrjJlBpeQlCyDMjppXuFYKYb7kk2vdV1XsWSCe/WF8DRiSaxwe
RoTIx7cM56je7meLReRjj6BTEZ7m47KCmvv5GpSDBIIG0556FflbRhD+bIW1
9rebQO8YWyjsrvxRwJKAP0ZC7vCA6yafengdSOBIGtbItUZ5u4OU332OSOM3
6Ail1k4S6gL0g5lCG3WuFFj3Px3sSHZ6/lz/Cu5C6sH8mQ2m+2e/ocdlbghZ
/QjyVsjYb56RyM1WA9XGuZqqfNhx7Lk9Y9qnvCf950HgrjbRifA8IgyntfDV
n3xUYiKiTMuzs0FgO8rOWZ/6Rt1Q+FxAUTdZgClT1WNr3Y/l4NFTpRh9Nw97
hbJm3RxKyxExEOvAeCmuanOU2Dsf9pFirj5rvyr2Zu074maWQbqTfA9SCEAT
ZGS0BxZHrxpC9g2EVPoiZnk9H2d0vW57D6b66emOIO7HOSzKYUd5inXa9Yww
SO+vPOAlp9fQ+1VxzEGjA+YeNFl1Z8ZftyK3aUJyVDb11Y90o2ix+4yIfXEV
54ItTlirGCRW27TvIl8XMmT0trZIM12v6w3Iqj0HudcCzmR0H0hRiLTZWMLO
HcncoqZd7OFOaHfAen13mRXPpiibPO4d+OQa4f8AYsUxjQgiPsLVlacoGM2T
ulDeSyP/rmpb1Vbaw4hCg5Ed6Jz0rkesNdTwRTJdZCTnTUaCqKNupaARAAvK
nROlDicfs+6dtfBuTr1XMbx1VXnUezPmqsrDRUBQpK9NfyVLqJyvzWIOaIUj
QVt/JOs1hBERP80wKRdrxu136RTa+EP6f77FNX7HZXiRouLzruzLFY5RMcPY
/S6Gcs+BinMLefl6TDCkiMbcCsH5pSa5BRN27Y3KLJGMHfwiLuFzF/D2vxtq
htu+cNmdP3+X9slyA4XjGwPU1Va5UxRahmezB6I4Kh4tzqk72zLc3G//Dt8E
I/K5NsQX+EOFkBvuYyyxO3Y8jCQPqGReRCAxnFxv0auwgCAWB4p9qqVy37yX
XQeqj9OOCDiPuv+M4LNGdkcHGCe5ezFJM1P2l+jNqsjTHTaLPh3md8jJWINC
fmkRfciWrR35yBEXMqUtO63sYQr/kdxU8j22bw4WQoBY+VmcIHKda0biX1x9
JM46z4xHfYcN83HO9Nitf2jqAooPJ5MYM3r8kQgnY3Tjo7raNwl5EhgP9zb7
UuUFAaXVfVBdtae33THGEfrCMhvBTcnUHWsZ3RWcBg59EEMn1EYo3VakdfB6
k5B9naZL4i/br/a/b8OefLVSI6CWWSF04D33InfSfYeAWchR39k9dzaG4UUG
Rexc9MTDwVs1e0DSLrgB6+wNQW7ECDCAhO+x2DZRvyDKqGMQoCYuGDNzY4zG
FEHQLHsaYALDPmHdCy3cDF0OPJ0ChGjUzcyhk99BiPEOttqgKQioiSpdDnKQ
PTPPhhTAJobR//JsGpTWlPDFTJkc8bkq8F8evgXYLXs3QV0y8fT2BHzqvs5c
chciIN4l7xh7r+6icOMGYHkze7PS/nOC1e7Q/C4KSeiyqJbp38fnS1C0L7CP
V7OVrFHyEliJv2dlweW3GDH4NsVH9F3BD/ZqEbZdQYLvBXec/OHDM6WmbLa6
IU3e68DzbIZNDOk+Es4hlcHhollRG0b/NC1atwggyiGVPjAd1b08wjYVayZ4
pecFfFUGetci+J5KBouHGDrH1T42wUxlenvMp6jwZDj6itDJFTrmMOw7cmqv
9H2HCZ6TkrqW6INcD0WulaSaZ4JlTyjl79Hl8eCpf/5yb6nNYPcA/T3MIEk5
2Es0TMcxR5y6XvLKXxGqUDLTjpFsRUiMnz4qC1yb/qYxfX4WXH9ba2C1I3vf
6qTeCNFTDvke2nPi2FNyof3uxpv1sHF1EWbMpsdUwb5wYgDYnJye2OtSPL0+
N9SNgkCrmjnOixIvzTfsKVHgl4Qhi/fzay6mb8WsaCcfF7claqrJi0I+i9uD
W8HhSspCqm5m+OrG6YDoXAlyt/GmR3p2lHU7TEKF6SdYKToJHbT4OXk96YFk
DiYUbpgKtSgklgrbwNOQRmEqOc70vglVPF/NPW62LPzjJWFR8LYalNPS+FPZ
7KbWiQlVgVmWDT94lJF0knBmDCaOwfWraR+DiSEmORNDEBpjtvGwGmU0c1YL
M/1UEo0j9+mSjITlDM0OaltWmZdHUyBMM57eu7PNmNKSNx3M4GluLcEOlho6
PUDPPGxWe45wT4lC4p8mEnxJ0YnsCOKCbcoi/f1KIIjIy+hCtVoKEN/KEsYN
7lNmKEIbsaYUPIgP3zW3XVE84Q60gk42InlX9LNGR0aDKa7DNqU0DgSaJrMI
/qOL6AvMHhWlvud4F8ahztNuNsTdFfGfEdHnohSFK8rkJbzQnvwjJIPFH4bI
R4BFSssFpgTjBQ6Agb2zCW0mVdVNkpoUq6GIIaGPmhxi7QXQWpT8hNpA89uz
cm5CIUbVXarkTRAwI84+tcWDegDbst/incMF8riLa4g6UbGI4s3Jz9QRW5g6
TBL+2nMqUowW5PvAJBkDarZ6OapIMyQv9ZUoqYFNUPIUOONxBSbi6PpsA8wO
SZRx2Kw73ZuIQarE/GE6Sa4Jc/VWj4ViDo8huIiewEPho/q+4QtL3V2QvLLc
B+HPZ7O8ryb2rgIgh50XKO0U0bC6w7zqNor0HLAoOHjb8ukPYf3/amWT2csv
iVQvOexd+w4uS+ItBAkAsoeY3HTR7+26bsj9qN18UeG0ViBsxqPAG0rtJ08q
WHbQWBM8xKHFLgmGHowLpNOJeM303vblpZamgYyo+Sx2FRbxe/RZ8k3pB69+
zoWPnScFREQYZEmseU1m6Z1NTlnn/GnsSI0tZU+sJm7Gvuq1QeclowsgvXu6
TgvKZtoSDNyP+YEeCDGNUGa3jDDzLerClDfZcyAx8uPD76b2Zmn89M1MgvM3
KbFYHJ1BwC9WJVG+zkI1I229/RVDxIxDbaro0AODnoulxSJHQEzRjbhpvrnN
DfUuT0wRwMZmu9I8c4+C5e+BoX+lwtfqpAITK8TuGSUgJn/adU2GxgErfUpw
agt5pppfGx5zGP1GCP2ct61iiMHsNu9mdQIhmV7NrOVQnXg8nnpI4v4ez7oj
2Hl4O9PjhsZ2MMOa2PHhiZvpuZOuVXiBLVaVEy+QGWYbdiUoIFZs4hSJ5ol2
VRwRRybqI8RINbedd12fkd8n2PYTBnVF/AtdICDt72Y3OaTdX9mnpeKJbLsm
Sty4G9YCU6hAI6XBHq1h9XnJNQ5g66hIncN34/r7PowyAJudfeRietergxyV
vcug9UXoA1S65SNRHIf3tPr61KDGHNML0A1UQJxS9SWwz8OiRRuCIj0pW6Ru
07mkpDczh6BbOz97s7eTmM6M3z3c0IzS5tRiKHETVNDtqeS41kOlajtYiVns
hJI+HAKYGgO3SVzePtauD8V1SQDdRlE/zXMkj+qdvp2qQ1uKpC8r2olvnB79
waZg6eP+HB5av2zdCGwW6lFf1yaNgN9n+atQenvA69x6PvDYEvDyRTC6h0l+
VjLapi+lB6DCEzCo1h3wwiWotshBxuQTILT+zKnEiLQWKidh0X2iMbh2d7v6
0nyBmb4rVZLi740TprAalMacELOci2eRHCn6MmhEyKH03cRgt9tcvMgMgHuZ
BamJyoqtr08ZeWBPuJy5cuPax4BO7ehh0dUHohx8fpx0lI8PTMSqMWGk2js9
wwzqZqtzh+PIATofHfW3QG/K7XbCwSvnk+av98CVl2sZjesXcTksJSkvlz8B
A+EkxxamhGP5KwgBE6zTjSCgt0Y0QnYvfjk2eZLeAjXTpXmRIU5irkhRDXEX
gXm1yAjA9cKAAaZK6L92TCbz9Gt8Dlt1A0az9GfbTMqIEjefdgShYRpL7I/0
zT9rmI6hHgpJ+yflXTivV77T62CRBtiUDamjiiXZ+Sk2E/lqAj+ZTwMm4RAZ
hFtXtQ7S32/F8tQCoZUBODAvV2KwiUJ6W0DVOcrprxcVCHl9y21lJaRXa2ug
IZja3qGLuDuGtX/A7tnXojKIa+CFm25K/GjM47dOTVgV3eleaoBwlnaaR2QU
WauJh8aZ7f/bHWFiu8Yl7zu20EPXsfbtQvX8MZj4caIeEjINZgxV3RqyiVll
vGG9T6q00VBQKpwPkuN4eU1jSlVo5UHuKxjOx/FLXGvSsLlsElpj4WnQQc2n
leMUApmDXt7tbbgnI8K2RuO86PiWk/QW5j/13urBknE3tNr9MMrXVd5KK0X0
AIdETpq1/JIxyQC3uu3iZ1DTiPf/jp+VxHrBFEulcX8vk+tbB1xlN9qmkL00
siCWZcKV4fwK7538fg2BdoCac9QDi1SKJWM2+eG9SGLPtRO+ahosb7Ed8ZdZ
UINGyXzpwcc/TVNo3ucFbrR0MQBdhsnCFrizpjnLv6mdtlXLXKgLhsDcAhcu
91oEthp7pUt+hUq95Moi48vT5rh7j6Q6u7vM5Rkqj5+3OhvfkizXM7MGrvIo
BQZXRBu6ntWTXqFnkJ3nHcwKUr/rXwRneDOjFbDoLM+cObwyDuk1iw+6MQWn
0BbqC3FwMYoL8Nb1dqMApges3DT1qAGbOm3ZIu/qYUw5HUXCrctV75udS9Jf
M2vQ4/nHhdEU/cszL/v9j5w3cu0OgSv4UAZkP8wxndM7naheDqBa1vJ2XlJX
/x4LuVRDLdBvjRLDJcSiUR4IMiD7bN59Z1nk+vvutQnm/cK/8ivRo51qwguN
8hugObwHCDzKRoy10C5aCf1EegPnC77OMQPOLHkw9fFe++7eXwQi3qOHG8OM
4UUOxHCeQd+KySxK9yxzHjz7fR3E/OYd/leWrvFjrnEi0gjCnR2SuQzJMcvr
cOP8fka0WZ+iGt6W9cC1JtF+DVW0FuJa2Evr68A6RXxp3wYX8ptNvzLjH7qE
D3Hy1F9NO2KtlVST3z3F8PQjkPXoJ5OSq/ymJjI6mJEzRNYPNz3Cr8+Erzq+
FOn0SHTeM5tiQ+6emEpvZw109QNxc5EaE93YnA6ffgbRn0Xcps88QFIWowHh
we76YA/u0aElQjFQnwjgfgIvnQJM8ZXEZW+5/UrtSZOQegmHcCWk4/Jd7knR
dM7Hdzeky38JaJv5gGgZu2MPuUtK3US4GneGDUKzJrf2R3SYDl2mI5lGumc0
nez9FdhkV+qTLaArSi31BsOOW/DVK5wanZ8raLegoogYgeoj2DLx3Zzb9OgJ
ANN9cMuQMAkFJ4U5GJh4gyIs+xObsPEIBE/K66k3xGG3JoYlm11vcHPQK1M+
ei69iPpuJWIps28Q5Av4eENtDmiNpOhXkeOfPTpjIzDfTID25Bo9UJJFLLS2
mK3UUDKeLWDLutPjuAVjvxfDwAL0433YGBKIyuth1RL3gg2d+qghU0WZVf8q
IvMxuJVVNyNtt6Of+x2vnfO2asLSffglUI4DC2u6Z0ZQ2YobKFoTY814cDgb
4vVIqGSSOd7/4i4P9cSxhaRGgnE1f068WkQDr/mHgy4o7WdnY+kefSQaLWYv
spxAGX2iGON8NelezuZVfk8wOvwGK2BGiwesyk4kZ+2kRT9qdhd6WfVcKOrL
C8ESCtWnknA58/6J+9MVyKuCpXXGWNsSLXgvxJdFTzSjeZWnM7ZQj02tvOu9
SHFSVOUyPhvZjU0gbKz6+J1kTS8UdbGMfcCs9xpBKqNbXspChcnz43NtQLd4
5XYEbOPgT9L4FQWnT8r3FJ/XLWJnHKSxIzrc14GYV1ieWtH9jAsAdcGhUKlh
Q36gszx6fgbjBKFvw79+HSHn1xX9QHRD31Q1pUrcY57ztz98HxIy1SsHs005
wpwi+VGYOtcnhJMSJe3ELpctdMiOpFj9CwqzLh9kBCFhFqJmlct7DCbYVKDy
ON3Qp8aDg+aRCMY5b8PryIP9UqiieSO+bD3sqaH5pwoVx8OvAttSqKJwIWVA
AlCzf/0YaAfgQA1CZnPVZG64fStn579CLwKfiMF/2VLsOMgb4HE5cexbcg0w
ZRZivyuqYao8XzwFZu5ruZxWIUqZ65RNc/eDC3i0rnyJgezT2TJFpqiTsbrU
3YkYha4M/WwJrLghuO7AFWebcrM8K1S4B0uTqoPzeuTJkAuyVCNXqk6UW/qW
OOvQjyq6UCzwn9XVZj+UMLtnKgd6lYVMRCzVcG7xnfoC/aUQ4oJqFQ7gE31y
935B0it9nMtQoWZzEmnbKNHEDsAJswfzIAsLC9kOVgcbtqbJD3mi+PTtoAKm
QGceEv9FAxyv/TZUdbMPSIClwnYKu6c6bLLeBinJIblhk0HyeVjFRS4Vv8m9
4vqb9hysZW8hR4lFypomGkmn04hLQ4e2n+a7JUbwagQvlJafwhjVlIrGepAz
1VBl5KZO57GYKC0PLysDdletpxNNvYOcAwnu6uedbageyuh3qiOXwaajPnYJ
H3jigHlvZqWtZRuauet3U2TqGCAOUG6HRt9X0YEy02jF/fdMzqYgqglZ7bVR
CqCTOMkEjtkye71cjJxTJ6WouOZUgwpsYmKep+ABDIg5wS1Y+Z1xNp9Y2I6/
fOGPN0uLw2hJ4iFKa89x/UQvB8rpinPYremeYYzU0x3tbeWYn+K7l0tUC+PV
mhxDBc+B4M5x2QcjINI2q7QXOTwkzy6ZbhBZEECowPQOcw5J76au4iSQZrX0
dbC4AazWUj0DlWBPx6wk+myEhmQDqid3GbUhaHutsFoVmdXNnBekZ9/eEWtP
/3VgADZb3BNqz3dYNBYgrE509blS6V4mBUF5+o8/5HIaFYOq5bmhqsytv4AD
DXZDxVHQ/bExHTVJci1X6gmp2VS9GONWVgNrcPOB9f3FCS3ihR9uGCd+7vWd
zRJudagEIbhcJmKkIwXPpAQ3MQ5O2wIl/EoGDt6dkmTFFFzLmbTaOQ7IU0NU
6WiYbvjfF6Jylv/Maf4ml2Ir3kHr/QswUcVLig1ql47YW7IrrBuZZx4kLdxd
D48qDnpSlL2i7nFsbRnNZOLFS5mcDgVV8QXVxZqkD8Au+usSvmdOUlgCUfAK
dq2hkKvSsBbIISOSVRAR6Yh+iepsG/X36AiqHD5w/WIf+JqDoN1IOTMB4GKA
Q1la2IPQ5Nd8joCbuvIUnZzQim1+gdLCI6rLdjSMuwfd1iZr5cANk21Kuev8
ziFk58mjij3LY9JMkHH+wSCUdJuG1AO9YHdADZ/pZb8HD6j7WoaM9PJErfLM
m3Vyqkj8SlmRNnLKHSDv9w2W9Jt6PIdPvVpy3BTP3JKJ8MHH/PULHcbsRbjK
w+KEwHbEBGaBF2COYm38xX+JfRmfpE2sOqo3L/D53gHvRbTmacRDUG9A0jBc
10LEcBFTqquLklwy0fnnhNytREyK+vzQ7XGqoS9h2Q5NdACBsS3aWU3JOqe0
0839l89VR1xbfcMpfHYQ1JnSYbY8r4L9ilFMN5UMjdXKqgMPeiPgVntWOptI
riEBaTcH3Fh1M11lCkgfzBQxWTUbA2Xcbalp0GTjghWIhO8tGMmjVDd9UHJ8
4kElsOdyjW6oHpE5JmVMfh1S4ZB7C3l9HwW2NbspSgpMlPT3JHxHW3eVcTQ1
wmAr+2SjXjEOPjoJnBRJQMPIctpIeepdetzUwnSZ9o7AjC55ykQowrN2fxzT
mMoYhN7DUVbr0iAnhjniYh5YrI5yXlX/hyFw8Uq/s1/+WERd93MWYQLHW15d
oA61UymH9jON0d9zrZn1uc1ZsWiemVGt+DGU92ZxuRYVhZ0icFFEFVBxP344
W3W4jiQK8zG7r+6DFD3Q8aomNO2uPGRSzhn5B7HJbXPnsUzdeS39a6BUlEVe
hDxrA9N+gYlHmpybZDsPstDpPPKGBhNCt98dzsf1O1E7RQKADAnWmCQcbZEV
mNrd8PneuPxue3Mgh8T4DVYnP2RFH9u+v7VQu82FDNsVOfZWCawhcAwMqnOi
1eW384EGBEMpDZJh1ZPhxSYgNrQ48917SQI3mplUAz8xmFIGcx+FLTACAaC4
NhHYn5LlaugAhjmwkO76/satO8GkeVo2V30cWXEuZ+7NsWqmDJu4GblneQnk
RaejljgfzIXFL4nGkacibmgWuEUO2Zom34uMMz4eVEiuljS73E3EzBGDafgu
1Zq5uT3z/nWULsIr2kPXrFusEFMdhBjcTqhdX4R4/zqrakDkdnm/Rc6OSM1r
h2dgRypU/UREP7GtVIqxp6ZnAexJtQhuk8SOU2rSluZB1ibrpIg5+KbSx1CE
px8t4qUGZ8F3qk/Jr2D2g2xucLlwJjxL4jczDzkCfy7Lhn5acn8rmtJGAyQW
cxxDwpTunbMXKO8T3A1843giQVi8jAf9AplKCO0JYxU4LrpU+Gsa+onC6r9V
tWDdzlRl3DPjIVXXdTHkTA/iXgLg26R9kPhKcjSDiDveTqgTNXhvVOwZnW0T
0ezacN+FUGE58ZfHsFQxCLwxP/JxwGLlebsC1HB+JxD2kn343lYicej2uLyf
VmSBB4qEcZgtEJTXxUIpQe/oq6b0zOncCqwTBIWHE0uL57hWHvXYhWA0jcM0
HYW3kdKVowq6oraM1JtNqhHtQ6d5l/MymklUpq/Sl1BZqDNTl9mTUWQjW1fA
SC1i2ZCQHdnj7Kv8RwYGQH0o/5SnfsPNtoM/iSE/nf+qsfkLGNIkYl+EDIYH
t5At2vuvEdgiEuhQTX+OjPaG79bHYLKBLAleyX2hrD3TFPZ01bgDZu8jun0X
Hk+nbefweIivm+16LcUpjXo4HX9wxuPuQZ6r6qwCEyZLiOvPMl4UrmYsilKn
IqHk7zbADpAqidtXO8LwRpv8A7R+MVyYnK8zp8Vzghrf5nvjQtZzvZ3QiXnI
q9pmGMrctvgePo8iO97mAHbWVwwvH92YGn8axZu47M/AiTp0Trugp1QeRzxX
PqW3lRjP4DfFdf8355wkYwErxv6f+PLn/4KyQiF9rZWuMI95ap2dbYcMLSbX
WRhNos6VczkBouLrjKHjlDOyJhAikca5nWJD0Qi4XAi8TWasUbCWoZTibyOA
D+06eh88quaIHkvEp4nBo+gt//D77sqhO/Ip08yLQtHRwMcEZnHYzlZ6Bv5u
qdRElezheiX4AA9rjxuPJhYX/nB80VUzGWVPYr8NGbImIoBshBW3HuIjupJg
k4skBPqtRIhPQHV8j9tRoD7QrlHAjx8Tn4uOwvd9C67Noou1oKP6gjVrGgVk
xUxjNrqjcTZ4z9YL+H/vXeVdE5lkyXnjtIsCYX7fS0LyuI9XJfLuhw7m17aa
pXenxiov/CDd5AORP4X8q9Ad1D/Dz5Qh8OuTqXGORxuuhSEvL+SrFce6UVKt
WZxDyP/8UMvonkOB9YcBaqSlz6wRtPO5lFaFDGsBKqrV/yni1My9tpxhAzoX
w3KYuAA9mRVc6J/8vKipFTMHXWoME7Rucw05qZxa2a+hO0KlR0loDAYVz9pM
bhybUS0K4qrh4mYnA77rlhhz9abcguj/+l/inuUHlGFmnlTeGWcIuJyHJrha
Imdt1rzfWbOqHtz3kCrpBqCbR/k7hvFVvizLPUIn3QPnvGGZMeEp70+gQwFl
T75ttZ5FxMM4VxevLKlqoXpZGAF/IxIah/IyEUJoGsdhIO9SAl0APr1MfZOO
MDiCOyxfwPaVdHE4V7G12JLq0chrragwbtw/0OJi4JkYfnwFgDTpeyL6I0jj
eXJcpWgt9ZFduqztBNO74ImDHgqaVjid9ElN0E5GrUI8M4wRLpXkHo1+9gDh
7qvyFRHHKvJmG3V9x90i+IEK3Nk81v+peaJsi2SFpVHZkawU8FMyk3GxH+Uk
R1h+8RUTted81e8Fh+2qdCoijuWWqk6LIblQ4byA54a5UPKznpEH9s9XFMwx
92gub99n9WeVLGWbYYLXU4ST1krzzLuBHppjp+ZVacD+O3EDYepTs+s8Bprr
9MR1HUd2NsXo7ujHa7zuGFd7vwLOMjEBegRm7B5OYmLrGrBOIEMRgGouQUT/
t8ELMchooZK6fQ86pvhOlRkhs+oytN8RZJox419ZEiV84FDfyr2ze2ZalMhd
pYcXqeHC/iD/+27OG1WUJcR+54C5wtBAZk5j5k9hSpEagK/x8u1FmKSHP6W3
R3AbZUgZexLETC9sQNvgImvPv0ovXoj+cf/bwbWeGfUUvmi7ATQAzfFuaV6A
2s4n5RLdHxGaoFEj2jxSShTay18OQT/Ff/iKQ6psg6XvVBKuSo5OSCl8IlY/
jO+NA3dFrerpz7U/MkjkpIrKayj+8sKL3FD/hgstXV40N8CD2NcUMNKGY65M
5BK3yQzbrf/GOINYKxQEHD5hAOey/H/mAw/wAvA+CjKlLrt7mzhXFdASZPB5
514CnyWr6tYvznGiBfHgIxxKmI6SVwgVe2FKIUYVkVUmpffo6N3S7N3CGrYM
SRx52T+yTa4+rDEkdTCmVp/tuOBz3CQrAIdqcwQ4fnVOkyvppqJddtzGaA0n
BS92ehYRqMPdRWcBTtutBa7artQdLtlWaEz/IYEoC2+satZnvFVwi+BaHNf1
b6zWuuOlJcrf/W4pvEzbbEo7FfiIh4UkXgb0ERliIvsDMzApjGrP2z6ia8IP
JxfkN1nAWQNd1ns8Gf4N96Z+VDfJ2ZA/nKMZeMp0JNVgRRgdQ1papvmh3EMI
Cm8XyZG+zbvhrKDBkwc2mh6P7qB9oK9YlK6Cf4I6zByOuyYqj9xYE75OecIA
gZAQ2oBjJyCn25xo3N+U9AFGwJNvngdUK/1+dFKfqwY92sPYqDjdFCIax3PF
+b7rqXbDtDsNzLbxn+ua6ZfYRefjVnncqsvUgS8PB3gtppv2PBN5Nty2a8Rz
mDPo/cpa35oLCATWTEj1LD5+nbbnYNNGLq/J1k3b3dhonuMoGSAawnMfer3u
87YqJQ7Is9eZXBZsZVcCx49zmd2D38Hy83lyOQlPzJn4dyWJr0V1NtN6XHAW
+m3urmHMaFmFjNxAvvwdzJps6DyUvLl4Ex2qESVS2N1d3VVDyFraOWye2SNg
vWk5YOBX5QdGYH4GyU+BDtanvoAB1qBx59d7j4GjqoG3vMXYYt/A7LMnkQXs
nINCuhqIiKHla30/d/IOsj0c1UmNHc2CotWVonOAbkD/JXcevZU3vxdfIZqY
zVnq2R3T3Iv9EQUSSuLKdBIDKaIbKGWMJPjpCXIUHG2Pbh0zi/l20iv5vGU3
awboWGqJ3C3YxLc78egYE6t2H2Hil+Mgonai+0sXogla6AC/VukSUFLHvPMO
++gC1x3byAyg9mvD/CPZXL28pRwg+krRjbtYeBf3jMacuAvno/DVualOOwIx
qo8cWR0c0jQvQ6EIiWEpSd/tB0d8qAqpb9Cxa33IQiwnYP/6PCy7+XJk8sEG
Gny6wZzjJRHsytpnq3jPmgmClotsl2V7/SyFKtjFl40UHvM3PokpK8MY9EqO
TruPS8Xnz044oFwv7LryFiLKbr5BrV5VLna3SdbylQRfZ5/C/zagaIMGR9oh
+bNRQMAJLllhSRTa2B1EnRdQrfR8R7Q1lpYi5R0lCJTKTS5gx7hsf7d9usUt
045IoKKmJryhNcGP41MPkqCpjdaJrRFV8EA8sQX2X9lygBkbpxNXZt6J1qTH
4+bl3YDQWnD7/a11FxSww0EipMRqPqd7zKqCidzTc2JEmlL2t28VCNey/put
Je7FjBwJY2v7UzS/OIcwDBt8MWgezcfaH9qYpnDaRNHNfcEAXxzbOWsNlEIT
H+ckb1vTxO18ay0Eia3im0w5KNqBd7AUSwr2EeZWBU+/ppVw1StMWUj/m5TU
/Z65HH1oBA/9qIMyayHsjdEAOJBGGADxQWDN0o8cPJaizdA2zVnDO7xKxUGY
PDPMGxMClt7FKEa1Q/+cdN62NOLFMLeOMCsHVv8bERztDqEnj0E7KtLVUMSV
Ot9FJ+rlR52dL7Vcah5ESW4xwdupSsq88eHtAV7CJabXI2Sk/3xC1xgdwra5
g3NQ5f1PNR/dNWdGxQvEImbWDZ2yMogK+VlgFIMZS00rrzXEL/tKSufoTTC1
B3pcSo4f+u30hB4T3l0PC0wkB3gh75HERVgmhJNlmuI4OOiGnB73MU061f4u
n0J/4cSFawkJTYyvPvPXBq0qVjr3hjRJZWGghi6eLLVYcWtQDZGMo0rAZvl2
6Y1if9fV66Th0Hy+56az6NqoCk748uDYgUIRgPHd5wTIQKOuiZNGtT7d+YUj
6RQ1jRuQws8RMxU4wZH3HGbXVAtaOP9VWIcxdrNKASkvzhBR1yutIBYX1+fC
IwsOGW62zw9y2nv45HJ8UvB6CLqUcyoQjpV3vjKhIMJW6WvLTdZ9MmoljqzF
pQ0+SJHgLJRjwU/A4gLJmnXPwUn+HOWOnitNtGIwBuOOOtTvRA+XaQ8xDihN
mHtMd5rQ+2PBdQ59OBfqkPBdZcmZxAVvqwXhQq9EBTHhNH4T0ZgNQWPnwcsw
3uOQVk/XA5sxkLpQqYIdXfJDBh2wxwRt48zE76+X5DXexNmJ7kAmRFutqBpy
OkYK6WzCzdfkgEwfxdPTTN3Zudk3r6wZBY/TCHZf3GvdCMRClQNHjVAmtf+R
tB731RfHhKDvbSo6zO6THuSPbgvDf7jCHO1moCO/odTedOdmqtsfHez6UBMa
dWNyYga7qEkALgHu2Y+pKz8q6UFokvYQgUoOnezcOdibcysgjKViZyqTERLs
qYp6CFTEKgzL4DlWn1XDW+tRGJTRDT6CK/cRoX4laWPUQEE82XSSGT7u0htc
6a3K9X8ji5SZ3kEVp/8BAG3EnSzTPUv2a2ww/ou1KaKRBk2tSxWBy2xtv/mx
4fZDTjoJWEYd5xsBVWpcDLcb7fbwRKfQ5X3u5rQsURn+jNro3XxCM27GBBhK
Knhc8vfWkH5ujO+4qy7C0m4Q8AdRJjyCogJxa3ZzT8Jf+yiJWDi2D7/5nuoq
HfBmt4wytu/20Dn9kBJ/BIVei3Xwo0JjXp7q3Z4+htV/wsO2ra+Vzoq+k8ge
nXeHB5Pz8Z3nUCHQf+FUHCILzR2+AajlcmWIEKaIDp2fZ21LX0T6Ys9rMmso
BXrnHSbYTVGakXNjd7qGk7QDpm8flwFh9ZBtsucAlQTlUtysY9riHHVPfBz4
ZWLEJT1gfzovfGCwbfYdvDuMDm3P/0vsaoMC1pB/SdaF/1kIEWK+p8hTXyx4
4Umt3r+yBR+OBI/fpemAtO9ccsi1UfKLavCqi04eBsI85+u9MZcr+0WMUkGQ
THFnK/fv+pKWwRoDGqlsPbkZ1K1TE7GACC4BhKMQAymYw7AZELuDMSjt7bIS
V983L50GigTRcHP8o6glY+AZm4jLp3/cSLMlf74XPNUcebbIRHxWDz8DHDqY
sliHRlA+hTGbl+QFiARSUqA0BToBU/xaCe0VWGR4OJvY3OomTQmLreIDQZ5C
4PEst83WrBgIGH9SdP0+WS//Pqm0l3vup5PsgFEBQZuEFPGil7382g1miPlU
zXgE7H5KcRBGuNQ8jzPEirgyuqBFRCXeqK1bjoPfJCeUT4aMhRwkZCVsTqAj
JoSTxFpc9AiM/m9J3OEsTgbIN9AKWoGjcPQ4aaMWAgkXJL4imB5bD2XOWLln
3Bdg0a8kfW+vAh6CpvjYSIRjkVr/JSjdozwiDILhuTO98FBNXjx1v+TlLG2W
F3w/pe/JShHPWCtMmg6oCqTCw6Bm1lsKlF1pCtMylPIjj9D71aQOcxqLYJPy
Imnu0j79I7dnmnq7zp2emTCMIY0P/vOdW1NrHgjJbLsscB1LvKdc5MtAPrIN
5KXrbTkdDafJd6L+i7ddNwJvuTvGBmoXdRsEn9MKk8HrNqVdEH2ptlfG/0IC
slh0VT+010wbamTW38VdWP+kU9ZmK7ee1MYm0JeYdrWgaNW9gIk1bNcPQ2I5
KcE7E6cX/9Vldm8Fcy5PmjU2UBPD0W7vgWU/th+3znxf6pofmWrwoVObRBsi
CwL/UoLXw9SPwQCPMTlbh+u9ifRnx/S5eenNhr/k7MQ+7PfNj162myuFudoL
iKPIfIMq+OlK50mSx6FFvSSxHisYNUIMUishBAZzFlOFaShqo13m+zaZZecp
8e5sovRxLq2pDuNfhJ8QPzbXaUxjoMz0D3vr77OptUAf+9FMOIRxL9diQ7U5
5NDT4q10Yg23OpaxZ2HANEGwxMq6uZZehRwLlogbFd7iyZkYn8Z519d9IEcC
BixPwT+neDtAPSPkgQrE8hLbfC2Wg8TW/vdPHR7TS4oDkacwPQJTFLkhvjse
NTn8/aoaulwVC5YA/ju+urvm0xJyMgYtxt34BSHfP4elL4egMWDO+ig/aQBk
Ou7E3so5D5wAS3J7xS8Goj6wKKLd96ldNPXS0QH+Buwea3QJCyw+CLD/B9xV
Q+T9RYTuMCAx9V2UvD9yirrC6hdiRTd/yWYlt1ys6pJdGlsaq+NnSbFR0kCh
nsSii6GE2c3TsmyPW9mcwVO4W6VA8o5bEWzMGSGqYF5q+JqU5Rv5KHLdJuIx
neAax61drHkRyfPBiwZqJWqnAepXREdMqCrT1VPLE/wc4ouOfgFOU6JKUDLc
IlnzlD3gH8EHfm0F+58ETLC28Cq66vrdiP68+j4mWMwEhLGyRcz5ux9WCzp7
+YrsfMJioE1zOB0WfwQHposT8IH4r57Mr7/xaD8/jMsBvii4ZyRwHFYBLQui
PjBJmC69QiiUV08O/ioQqkBY2IjDluMVDLL4UYbQ9BLeoTgvfhyv9t6VIyHo
SUmEaPxGBJhs8HMylj1FQiL69U5sd1pKC1YI1izW2IRaOIXMBwlgnhJP/cBd
/LbGBPi16IQeL+/CHNoyI9emfRVgxKg1u0gD0Mye3PWwTA7thV3Dv/FKYGzy
Pte5gFvKIY6xP6o0mFTWQtSEljY3yRy0mCmUD17gjaAhY0oTYEdKUZumzBML
JT1HFoI655f7OpYLE/yjlKPdB0wj2ILMjWuc9EV9RYOkCf+sFLjv8fv07CAE
3akhPyq13xobRm7grShYEG255ZnEuvhKwOUnFah9I1hGlQXZzKKeJ1/JVHbR
us3oJVjmmoJoEiK/JnfL74lIibzA5RFq8rMsELL8K1z1YbeenyLv7NW4gLSa
xb5KCK7xBexEo/bqAzeYZwyFrSZ5WrGGwSRSF74YKceKDAdnosOkwHJjGuGU
8/xgoLekg+61Uxxsl0KQokcZoYTm7IbV1go54yl2J1mcuR9aSJ4obGuu1qfd
H+kQ1p4m8ZCJRVgcaxYFfiAbO+XKp+2Ex1SaMFf8sOb9CEbv+M+yWdAwWSab
Isnzc58F+7WmSEfiUeZtnNAhzH6QTfQeCY+Sje5JmbqQHyJJxfpS/xQttY2O
9V6baAgeZkkB1C3BlarzYIGEmxGG8pe/seO2jxhPIoN4NJazphppyhsGhVHl
BGi0EKE4dxsPOLUvEW2kXPsOlpYzLUAtZrwV2WPvUU/yTkNYV7VdWoYRJmyF
+Lq1En+FDDz8x4gObovI3fFnoFj1iHS5QVhb4IPl8I7lxyPjiIPxL2iLEnGJ
14yZOZpIfIx2pOf5dFTz6lx4gkZQ2+nDe4k8lL7pz/tDtP+05WIB+ySMCkdy
ggYV7zxmF3yS3M4/V46xBKkNd6AKH2SgpYoNSfIaG3CJ0PM5jkx+g3Mg8Zga
eZk9BJyBW9QjXBAScCV6qwXU5+j0XTcTxov//xAY/njykDGguSb80zyDAMUS
FOPXNWWO96W4N56MnSmsvTKnqMX48rpDc1lJQ7cz26KsTqMr79wSFHAv80hK
w7ornVGjrXLADmExnwz4P+npIh8cvTdaLZJtNzpgnP1pYoub2NMjU/G3IdaH
i9FHsCk7aM6zRoAU7B5ZKQ3vAkr/Ltl+ZnMIiBhGpnsELxOAvYfzrX98wZwU
qb8VxrGTvAzXIa1PkKoTM/lzkVp5sWH4J1nCHh/mNGPdihm5SsnORnHptMjE
GWM9lVpKoBaHAG1AefnES/3D9c/Xhg8A9g0rgLXmAT6zomqrzQ9hWKXaYQK/
88CPpo29O34Ab9H9L3o7fWDo+qkQR1OHy8otiGLCtQGkiZ7RJyzZrqaHp3Sy
jvGgpveHx4g4m0X+SzT6g1OZLuR7E7P9OPrYGBcJrHTY0GJXenNqTEkHVv/F
sMO4OJ2GtFNkhqUUCOpysCtXnKW0ufj6L+9rQxfnj1SRNwxRD+d3S/Qggcat
OnG4Ed0+fusyREDidA/kRKzjm2lvO3p6iRyH1j3D3ltGCYio0dbOwFWLP8RC
2Qqd4GO591bcBFzZ73/D2kWgUm7HjPjEKM8KJ6z+oBRGeiBzhKAx7m8fLc2X
UJoBCyjgWedy9ipJdRXxA3ocDlO0b4hgrtzoYYZbg/ro+Pc78gGP1WZzu58g
foBWndMqoFbRBuvOPwy0x45ABVQaQgp21n0NSV/08O15yQZ/TmLGgptkSyPn
uCIreYqQlR9zIuysOsyr7pQE+d5SOhBI/UqzOtR5nGmZIPFnQB4gT4t8YOW1
oAK4coTQDdIhOkjd9km7ZNxIle+WD6Pk87Pn3GVFL7W3gj1vftZzzjg+tkrE
Gj5wVYiRHzexfi+nD5rKuFZj+vsyNYriXaRHe+VXsyyn79NjU2UYPqpp8ZEw
q7ibxUNnCy/S2mQfWmtphtN365BNHAt/l4e/I9RyWZ2HabJxD7CQ3TntiXh2
DUQ4kFCTXVHrRej1SclCiPbt5X3SD89WFcMM9g69QmkupSgyZCTB8yV78rmv
+22TEIkHz+mtfUFA9KIbohufQ+pmKraNaR9rqEI0TPeo56C3Kx2vRSzoUWPq
fvallGx5Asy5YnDnk89eqBI756JqT8WgWPCm2FDjfwlGY0DTkEBkKcO4Ucnq
DNrIMDBTzNR9P6mXG5cLxSVqmaegd+B7pacK/HgaFvWCrY8nit2uLsx2tY6w
x3ljwZYkfQxzL92si++JxDHe6n5m14LXhYTI6PMBDT+80PtN9iHDyRpqQaz+
kovQKNCOFRtys9aQwWuh271FOAntdRB8+M/ztYD2U+949nycETzVrIAlLqhI
WpXtWsYjALCKO5gfN/7SAbDTrHijb+sKQUXYyHTcYspgToHRifBJ42udqHIg
jafU5VZdXiyHy991+wrssDgn33hGNgmBTyPKoeZsaFaZ39UwO7MSMeMd07C7
Z6q95AY689kFqbrYdajb3RYCWuEaVNrBBg7+geVZ7wfAGAZ9i6P1X+GuNFEw
5WkFNOQWW2SE2LbEyomWXqRmruyJKef62aobPRgEc8pyHEpgYgnypofLteJu
BeDwV8waxrJVOnTclvPoysum8h5hVwiJmvgi6qKYtmdHUEkllGacUnYbjCB2
DtIV14Wuv9hP8U3cNVxpJ23GCeOfsIEBDp1T4IMPnBVzSAFj7wmoJuki+MMN
tR5Ojlp+GxuWJL+JI9bsi9902UxzvCXwFRs0M3wThS+LYEc/42h3YsfDUTQx
Nze7vmPUZS5xEt/a4lzxDtpPxunA8taFAgNq6zLKG+LqTFZmleGkYyuuh1tR
nOsgEJqUHSVUSdcNDnHqXlMGv7vyUsNH+Q380lsHyP9avwQkNpMJyL2EHV+r
lZ9CAKkqF9loo11bSgjvKT3AnTstn4FGga8pStjrf5M9gDTWbqgD4duUB03L
NKdcf8QXKZlPggo9eyxpORLd4sF2ZlxlaSAL2SKmmafeElmjjCKViHtfVrEa
9qZCEjT6ucLUezh1Y7lGIcIdAgnXg2bRETJ54p57BgILSX9tAXnMq1frcoIa
UBkH6OMF7+tt5BrOAv+7by1NujvwiRtYcZRjhHK5cVGiD7hnpWXUbQD0aoKs
/8rQgWL1TvMrxzOw5zYmGt+O8aLNylxnlANHAKHbJt4SIbu6DtfupMSwSrLb
65YutyeiGsgVYSfIBZnJB6tSbS+XEP0aJbV/jLoU5TnQ4dLh7YfPRSSAPJiZ
xBQ8F/DUSyzPPeTUNtpkVUSU51JmbTHHkMoZG9K3yxvKeaEC/dzpBMsYzf+Y
znouodjEcxiBDWjUnq2/19Jfce8AhK1ssljTU/zyCP0PJ6TgrucXZQOWnJ/K
QDcfhLp6PjwVqLw6Wpod0JqGGCYWBnDmgjxOkaoinK1zdNl6B72OK8Uj9HTm
7l/FU/rcqEbTZEEbU66gpYRRN58nIfovcx6/tCXj/VkkVw/DQaLjtCcKRvVY
Zjnzlmwn0Ma3IFcc8WG1KRioLigebcthzdXCeuJoSVdr46rIPGo8/nvCFw4T
brdwj4GSysi8XoW5w5hp1qU+Nby0qnEn7vhVHDERo7gnkBRd5r11W36YiAYI
DO+Gydw0ZvN9E5wdWNFIFtIasXuIQzd4okQ7qy1xSwXsiHME8S8SY9DqbK2Z
pkFiqZh4fJ1SvFQuAs0TVO5BAZ+4AEhsVnZDPszamjYaKOena4Odq9irBlBV
Sm9XUMWujKeHWNze9KomEXdqCoa/t5T4xIKLD+Fyax9AWRg8y6+MFI3P+6am
UQPpUsqTNOAKZJ8vigVPLDgI0GQrDz+gyPdyKDlbx0yCKf2cHRCku+bgidyp
QW/dbJpVl7Yms+X0LkPd1Hv1CFi7xfLiZxONBkAN4IGEX2qpO2/XemDuYuj1
xXduT0KUtNg4Yq2ElVadP8TDUs+agTX48QqML3E4oupr7UV2M/R3CB9i9YwZ
OzGDjRSTgPR7NnPpF4WzKzQDVoxDiUVxKUpMXndS6NK2FzAzlWJqMzoyNRHc
ca0WdmuTbm0NC/DaYuhU49/M3YRuzNwj3dNR5bb9Xl65icX86FXKbpJn19Vj
j5zWBR4ITVcuNA5GLc/Fu874n80DgsjqcgJm9hTdi5EpUcexRdEV1pjhdDLB
sSYpGKTNqDBhThuCDHtpZK1P7W3t/ZeP24972d9VZWrDjqy+ZanM0jjh3HX/
eItGRFhLdGnqPFonR2NunIhFXXvxGJeW5vOGZ6bn1IZHam98vojOrT5evE1N
bb0Ckh4aO1KNpnH3M6kdeU/gK5fTCQ1ODfFuIzQRL2dhD5s3mYTwjckGnV0z
dmsIzL9W3PKCK8VUixelK3XN3LYhaN6gcdMVGEJC+/wmFynA0uIZSljfJ6ZT
IuCCvxOanNv80gjlbWlBjh+PYSe6cXmvDvW5VQg2DRKpKkoRLEcBdONftrDL
zjimhFEOOHKm3FhyRQvxZnJSPga/lysV7+MhAZlg3KMfmGNVATVjgu4sjNni
Xq1N0tuk/ZiTxomodb/q5OYIti/wO0Y8qwh6a5CI9UsrGlQcKmEF56SnhoB9
ZSiGKb0pSSg8J36rWO0DQQxLAmcEH77hTJWmBFqv4xv8/QaXh62XKf8L53Yr
PN+RAg1738UfLndY6hxq+Kbq7pZCWI7Gjvujpl98EdRlpVsC6YWflbvHWyDX
bsERIlHJ/KyfUIeATls20NJwfTtcSaRIYKVkrHNeeJQqMENCIr0AvjzNoF7V
xKiKULi0mpic9aEcePG+stcUdQvCxAuhAHYCt6OjOMWZ80PqblKadBROZvZa
9FA4qEbqE72t7R6d5yToMvU4K1Al5/IfxS4+4x3EEfQmdY0Baq2oKfbyz9x4
GRSzPdSvKkPVmDwyLR9pxDuNRW8NwmATYUxG69g4KoBEKDKeYV1hfnKF0b+7
jsKCuphLl1FZEWkHwbSF3sQE++AwVy/Czz9qc5RhRkApTnWPU3fgVHaqYQ5E
T4DQy3qtN0f2LEPYuhkMUFqZdRlQIgzE/s4hslLJakU+93P4y8wu2D6hiVRA
QWopiZrXdColQa1D95w8KgpnXb9r+vsALKWFApM2tezt3DfxKi1GQB772QLV
ccG1ZGb70E0wiue56AMvQ/MTODYYhRSsHbp+3QGls6XbsC0l1fzI68cxdaYu
WynSKbjJyMkK2Zqh6+3arVH37himsox6VzbgUWkxT++IvMJU0MY9xbMeOXnJ
SLCG0PUCWdLNUo3sRWvSfF13wuhONSe7HUREWTA+ZC+M1TxRbZMtyfNYngFm
mgKmgT0G0qrGuLz9e1qagJ6uScLyMWKp9Yxk/Qns7fovqHB/+BrsUfhZBbdK
5YS71LBcNlvJA3DRW5WRl3qgEHeKLJjd5NNhBIecRLOZDBVRfdxYwVql/smo
+KcRKBo8Uu0M94Il+S2uFNuBJwZYPyWam0Xm66d/mwxrhXhm0xnn44DYAZSk
XJ3AvhGs5pQIT4KoPysOfoQQyvFqZuXYPIBkNkHR+fM9AnpAufyRz9+oq89c
iL2rjxkHUIVZjhv3MR3d7PHglnWHnXYHTPHFdY84g+L5Tb9BcXMWlBNFMeiR
m/tb5qAfigr390e9QBEnZnMDHndYxW0I7SCE7Ipd33UrkenKFYfEciSg5P4+
WdMLS1biButXmg+JS9jhGaE6zfBuGBDreSMJmDq3XSD61GoT+6pwM55KPlE3
hJOIX1DqlWVFS7tWAWOE9v+EVsPlXDVVCJ+FXwxY/B7ORhYF9E2Iak6GUY/f
Dhj3UTe+YLgAbYjI7/o2Bq8yx3LdAm7z92zrxbUrhXhgvtnqIoSSBlqxx1eh
x2o1elcvqNmfEPJCNnT1griRx3THVsa66eG0un0pX1u8VpDCWkOzCbssh/Xu
EoUroSnj57uy4LjCGOr4ql5emdOVHFk5IuY+A5O4YYHY7VbGbT5WQsfzNYl4
r6CVlokn6vc8vMNnllnzuUXrU2ruaDD0WCHmt8R9ApE2ieuqKeuPpms99Q5p
Om7E6MLpNmUl++1hVuOIPJHIvVX8ZYIeeRM1Fl15Aj97pl1PBhpQsTzn1/y3
eTM7jOs8fWU4HdOH7pY1pf7uKzHmfV+QiOVARvlcW9xcJAR8EsZA5BjrTcEt
TZZIqQM5EnUHkN2f0+YvSoSij3dV4+RQFabo9WX1foKFtkCi6BrOr446Z7dW
BSMZXmblQdbtyIFOIUxC/4ewYl5xKaj2frdmvVbLaO4qCidkAA3UUVmhcP7x
5TBUJ6wbfKuGh86P66KfVcrwBg8Tc2WIHplyrg19y8/AMRxa1/X69iffxmmQ
FDx3usgLGjJTP9N7Deg9NQnwu3eNHhvCOj1MnkP6vFTX+BTVL82F47NRanpl
CF+IzqXpZjrLUqua1of/UDJNlHDyV5tOnbE/ocs4qGUB+oCPdnlpWfdKydRQ
kXsizlWNJib9djKA+ImyKYCp4QciBzH1tf8qIL0G7IOrb0Hx8g/l+eyyNLYJ
hSItIkXhVUtVmmC9lmav+IPi6Q5tvDcbFNXHzUH3O6kVgVm6nmZHwHFgyWR9
jtNCAvW9T7U/a8vfgoj9AMHHuSjoTMAS9cjEwtC2VZJWWXiPgXqI1NCk2GSc
PGoKzDn8MX86MNUV2FqK+x2k//zsot1RLEK+C0szzGcvaCD96ZDKWEDzEcsD
QkhvQneTF+iWCOhf1P3t59KJAtGUZy0l2DFoadYePmXJGVOtqjhTS6g2dwzd
2wiWO6hdXBM+hfLxp1BcXqOxyGIXnV++lU7XPs/7/IMZeldSoq0sABGvHf3u
JtFHlG3w85gvQpf/sKitOibXKzSAsubRve5t0rYHP7DHUFrKEBNY85Vgxi5N
LPkyPU7uYx0UlzJ+W+Qpj0J6YKV3acr2nF7kE7NEpSDsDKkXfzF4202SsIPj
2alrqZJQTCdX8SErvXQgolEUo7x8Et3fZwglWn6I8CczRB7Mjh1ahXB4vAtm
5ue1caz3lmoohsviUmeegApGM8bacE4Fus2PV0gDkiCVL73VBVzxluY3ZKeS
NWGVm+3h4+kKh9loz84Zv6R7ExemtykGHKLNxu5OojUM6V3tLBHBqpwj52bo
HuAiXdDkP4YMoenXBrcM8I6j8rqjFWlGdX4BkyRz9m8oK7W1cnRS9u61WULf
968xBf4TMyCLT/oE9CdBup6x8FOudXXQrHzlixqYnfSW4Who/27BAydESbQw
VItkxsUzGpGmv5+E/YmLl9VUBZqcPD41ceQ7JjqKdCKW+hyVuJpU5IHjuyJb
WvskOaMospoCwMol33rcSdcA6bTQKL2Rrge2+5ikzYmD5vGiLCRpflR39bc7
UutAY3iRHh50G/GYhe0AxcH2tXFPj8/7HRZTvCOc/sim3MZMy/+7Hy60Re6D
JKM/3m98YZJBeN1WX/8I1X6goxfaRC2JGx40xFtQkeuHSJ+ewJL92DctbZVH
Rl3ws0YSWVbZf7zPl6Mcw5AiLlmIrPXkYlbwsqLC+bLGTchSyYCF5ozN+i/Y
oPBujBhhHtTO3RYz96TR0fmADiu0/UoGguE9tjnBm51aF5XSPDmC6T2jhv3e
24SZaqFGHT8SNv6GTaPedSEq6WURMJTsicW+Izq519I21cVe2EoHnBcf86HI
dEx2fD5Bq6HWYE+uMaVF+TG0Z5IEyH3F8eJ7cIWztEVc1kVXAN5qMvoxeLl1
cUvDJzVtNq3DNcpVghQ9Q2HXjO1g5ih4dlG3TgzLLjQYsrK3TCSRa/PfLrkU
Rg+sK2tTYjRHNhW81/ElCf4Tpe/LGJkhlEYduwVPU4LFdsLWJjQ1cLaYNCeS
sRcY9F0H3HUHSR6KAgawlON2hWNDCtQAENG0340H9bdVmIpGFncVZpgvKL3r
jUAd/xi5K6u3g3J7YN8MTEYJIAHGLzkTWc8twXygBUR72CMSU1785zFjv1e8
yidxlal5KDER2t+UiLiZrL8XJKd/lnhQ0DUnUpRllujvOMgWGeiN/QD628x3
nfwO86p1eJY4fuXctq2XRzwHsQWIL5McchBlpo9jrJpS2qgSp4IJb6Ha9TOD
kn8U1rS/WxQvf1Ffi9rTdnFx8Ud8RVsh74xIGBPliMvFLolPhRHJoHtGqGGd
QYAypyT4in2sLd92M41IgXnboJC8QMW0rrBSes88scWmglqxXZ2ypDROBIqX
1bUILOLUylO75QCPoKD3zigNj6CI9PJSDFjbk95oBdoGer3Qzdl1L8kP0/fX
H+CZdCT/6dTSWU4/FGZ+3eKgOTZsicbQOQtHoWECLu1WtFvXAjTf2YDEBJUi
6jHKu/+UV2K74WHWcUOXI/QIqLZyNTbT2cPg5+edGaLqkBaV+JvONh3u3DU+
0BeiWn2fRsqZi7XD72Hgsg+sKjN3WAx0jgTK7ZUCKPWXOPpFsEou+TS6Iw70
xuKqwzgP3QuQJfM1TTq1+cXQV9eoYk0aOOKK8mEBHhrHWtKlJElFkPKoGxo5
eVRQBH0vOoLk3YsR459vBzqrOIlFDJHgjBqhioK7l+vAE+eyYw6hCHCx06ec
5Vyry62cmmYRY3fAMRreDSus1jfM7Zwrh25ZiG4zbEeWgr6aZKZtTGCoB2pK
mcx6X9I1S4BY4aAAORubOSp3z+brvgelD9+WWCY4d/dQ41FQ0bKwqyczY/yY
7Fi+Zwsn6zWpmpfQmRTYqnrziGnGkgF33boSgUasc45feqsWv2YkH3oHZShX
QwbNqHRAnG1i6sMLBtZIfPC6poXiOBpGO/f0oKNclNv/YpUQWfxNper3FSG2
nTQ0PgyvslGk1mxs3yc5QRekAm3ctK2kh+YYXlZKnn5zScR4thpoVR3Tra/j
n1ucx83+tUQ78BmSdPtztC+Ssm6PuxMSZZEv4v4RuYpJVsZJGDi9jPN87rG2
AdCfDCCVFFU/phlE3j7dL9NUXZJgC0GBs2u9Lg8vpjI3LMzJLkoNXgm1AgS+
GmvCTM6lOGroamtooXgHjbD2K/ZiTyrlQRkNfTDhoG/jexMSbykZObQVuzjO
x5UI484Fq3lYvwo14Xw8h4dZRxszQ5RNCRE2WRf3T7eB+41CxY4f3TEtGnMW
cBBZRJULlPutNqt2/BOs8dw+rxLoAoxESjEMtexgUSh3ijWXGAAQMe9qB2Iq
aTRGhTAjGCFzxET8r8YmU4Y3aTfI2/m/lAfQ2uNxaifUKXjqkx61tbs63T0Q
jhQsiOXTqQbJ8KNxt2T8sOP5TwGLGI9fsRQ4ORBwWYrJjuXdbEkFEYL1nTiW
jJA3BTeYnOFJaeeKSvuIgJWMQ8c8nS2DuIZwTUDy5Gfr2hGt+JHvCfNfR6Qa
Z17AhcPH+UdrtxPDjTNFE4WkWbR/EIIblTVmvEZV9GDfla17cxjI9jdAOMDg
eS0B4h0JI4U+meauzcnjBmvWfEw7KgJ1OR2edM8uuZ6fV3C9TSW8e4NYrBtV
ddTwWcH0mW+LtZwNfTJvvL1AxAymlH3ZKLYDgC64Mynna3VWpTv43iZ63WzS
RVYRXwBHFFFMbqH2SXABWPDVrnu1j0BuqudiwnX+98UF8ouqTlvAQpO6EOed
7DlAFS3WWCMCVlvnzVF4YjSXgbFXao1tH7GQJh/suUzBv4xH9aHUpc0MBzFC
esavd5Z6OSxW60P4n7ZYr/W60YkudBnkRyfJZduqN/hKXvICDPL8/Qf+zszp
/Km+Bpkj63tpViZDNjEWIfs+30w9qVaPRdtDDYSEK+WjZnlrZkNNBuhWZvdL
t4WcqXPYyz9bmq01uDi02U4LVMmqQN7k10Iu8x1tCiQu3zqDeGx6oiu49sMy
yU9rHvIIL2Q4P30ks3HKoWb3UIgCQVqipfxLokqTRXEj9Dqsmvb9RfA3oCIn
bAitIrFNy8F7tJGzlS3VW9f67ai0DIGvHCrs9n+MNFgIQRm+rrI+ybmw2l0/
nwmTeKsgeJoHGf0dIgz8V4bJfvnL4WblwiZMvCwROjO7h9nyUOnwbRMFcDGr
hzRmk1gf7/IJXJjlCDWxzwCIznUwCa6H14eWHlOCjyTLVhaaXnWsFYPt6Fd2
gByV1XlrhZTLHGlapSeRi5fseZE5jIpsJ4LQ4facdVo0kKmu4a/eq1MlgW7X
cGWLfGQWEjDg8q14eQ1bAMgHyXJnU6hZd3yVPvHjN8Lfw2G9Owuqg82YLhQS
si2057CAaOWDFPf/AkAT+n+Qxn5DGJ2V2HgtiE5ZdpEELnG+9Bz2cRIoagkY
uzmvnpZHD15m05SK0ng/8qUdapUYTGf8n25rUZsihXlwziy2bHCs7l5BkY0k
/Mu2wBTDjapzLgYJsW2dmAT0nasIqcCoVywqdmRTrO/M56QCyO3nI02tzwC9
JBokxVY5tV34W9pTZpxeKNgX5iCayYgYXNLPMe9I/2z9ZuMhhv9C7OdlNrPX
MvwSo75w6Ek1mAMWDqDIFXCURQhcNdafvIrcOqxDQl92mBz7KnXAG/VUrOu9
xJPSRXrOcL6u1lfK/Aa2EaLUAmeDFmsHy1D04/G6ljOHTaJeMACrTL5qVRIs
95ogxNySGxYTHkRKsjxVPV0Fcq97af/ZkXyRrJPQ/+T63XiyPWVlIY0eRC8D
1vq//8dmfgSS03lTauId4JQ+PnjOylr5afyHBXbY7DW/IoTuqtuWNFvaOPd1
nX20aEMlhwiu36QXMCGZNxwvYenMq8nhq5KPFgdEZde0PqvuVXmtj9wT57xQ
FmK5trOIoYPLzJg0HaPWZlFfMUuk2KRRpqoEtnzx2b1pPNU1Qliag3/kTmTO
xoyhHLk9SlE4S38nESos/68CxEE3o9iSh9kTxHfCMnLRl1PLyQGVfMpVfeFB
4Dqu2s2I3eG9XHcfIQ/cP6ubHj22xE7Nrp45L1q5uIjLrcJbol+tQOboDvD+
DXuMmNoUNceUDB6HsO+qu6XTpR58fhhZ30zNiCwsUdFjo6le64k+ztetqCLo
jPPlV9B04bJRSdZN5jtHGSr3rUKsIzzWyTfmSIuq0/IF//mvZ6VxUvEyWS1+
ycIaH0R+JDYtxWqwo2o+pVqCwzRf09dns70iyt5h/sVnknx7oAWIw75DOPCC
ioCFmoBFLxKSgqw27Xr2neYKStb5nPVwp2sl60gfDK8MsaxAI8cqu02cb6zp
LQGZ9xdzvuo+EMXKxDjySBM7ptdygKYU8Zxj6J2Ot+8RUMaBMOObwrj+ipyw
yDrlAQ5j4YXiB2wWrf/jy7tBLB4JxZQATP5AoAs3zs7l1Ml6fCpIhTr+WxvO
phqtW4mtHgERWyolpdvtZhImpBtwYNVco7WDBSmnoO1eC0xy44QWGPwWvpjY
O8huXcU5ZQQiRHwmYlJdwsgsRR4N8GsrCwOb5KD6mOwLYGNcums0o0UE95z9
0Kz89uGvp5UhSAX805BV9zLwT0PEwiYpMNA5/NICqROMb2P5a0l80nrYNGsI
LyCQ3E90HIC9+e5BhCWiNcD0iBZTs948FrdPBiypB3S2wiF8gFGocj/4plRi
chC8Tyh7y+9WDvuOn9OQTmxymLPOkZgCAWo1Oa3Kw7aTgsKGhFABbo1CuTF0
fniF1yxCZhlqVe9rb1ULGjeiiv8KOyaCmxDuSLRXnVfHzIe1PYg5ZY/ZF8qr
lhmdsjRQIuWe86Aj0vSq9j3UiWW5cltTVzQmyJPXtFffEcxGDHZPBbZvgzv7
sTn6n/n3KZLNxmtoJA+BOImG4JTBjkRJq0xwHZy26D4tMiprySMXNOyrt8Iv
7fmNTTMQpT3TDON/rvEAkPEC8Ao16Ku5fvDYsjzSVbzU4oS/JWBtk/erzn7J
BQIXix5B5KfzG9inbqf+1jWA7ILyzFKH/Kvjz2cKmLgMAnqyurrQEaSgz5cb
Hnc/XdZYNwOJhSrBemLx1X+oUNjpFmfoZMrgASiAivtOc2aIMFUcDvUr/dTg
gMvzuCkfjqV67ned/SNHV2s2gHdShS9aqaYFGqY8VbIq0pqIvSNJ4shjiyLr
ehl4yD0XEhauNypE8wYwsA/JcUitTJJEgI2nB2k40pDrcboiVGGcr1E22BT4
etal1MpPQ4bpwW0CLFg+V5ShWyyenFfJ0BRKf+b4oMDWZ2u2y9YitwseNDuO
LY5qseK3UcWIChtdTcFS2enS7ThbPRIFOHCUlZMUCyvTl7lFVRELbiSDtvk8
rV3+/fMfgIwgE3QtN/rO4XyxcdoU0R043vE8Ukt/0jX6RjxO1ob2DLeqoUxn
dUHnTw1NsaDSkURAkv4Sxm8lYl0kbVmsmr/sr2W8vOQ+80VxRm2/7435Bs5i
dW56Z011K952zd+U9o34PQqcc7RIFmlRe53FHzBvhdy7HtAT0NcEd3kEPO/8
481q5TGGMSCbJfyA/pjwEx9BumJHRWlxdYZYQ3+q0J5Fev9SzRM7ECmyLubI
e+8woYRHgyyTV7DeiaNvQm5v9DpIsLvYbWGMMNNHRhVZqan48mBwhrigkqJv
jXjvAgOoAfHfjmftY4cAwV9EqI6XmUWwdlIx+9u9Ud6MaGJ13C2veQU721p3
yNlEjTlE+49zM1SEvP3IYLxUy3TuMPaFrtuCVGyMa63wkiwTe7nRB6uGmIbb
O33tbJRbzOHfg2KFiVSmFiClMQITbbwjyn5iIEnR6mjn9OOFQO8td4VedLtW
aM0ya/VF5QwwtdrdE5VQ5ogzFzl751kJOO3+e/RYqGFFJMtMiF0f6JIHWg4i
GWEZQ2gJzE1j7NywKGY887/aCxuJvpd5AVxEjceNmuakgJLtK1vtByDasqzX
fsa3O0Kuu++7OPUP9h0bRd2U6Dm04lNXNayWlvTIaYQSICgCvN/apeyNG2Mt
fag9V2Z77LEjHTS4X71aGmuj4MUAjPxWi5dhdScKNms8dTY7CFiFSp63dkRf
RfajVRQJGPrLKRkCuxwc7EL3S4wg9Edbzs0EOW5kaxxnjE3hAKdVNOnACtZO
k594GBc5Hp1h7U0WSVcIH+4OyX+NIo5fDlx2FlRprZdqqZUly4mOZYu4QqdZ
vQ+j/xhcR8AE9EW888O2ioFBvE38WykTtiXkcF/ytrM4RQajMNvzz/04rCHJ
Z6wiQofeU5PLfmiqbl01nMi9wo5dvUtXBH3pjPtFvzSEm2/GctVZjUdkfQL9
3pjZ9jYuJWQ1JtSeW9YdwdsrSrCm/ZNVi6419vXBPOJfPgeoWNgl/cjb1Dub
D60iCFhCx+AYXaU3H0QifLerKUWOFBruqWQ2VId6KlxcNoHir9ah1zHSmHES
J6IWKXSsXhUnb6ftJ36z7MfxmQfy/lVFN84QjH7TbQnT74SanCmKyNmfPm0T
syjh4AqFksNqNu1+LQI7aOYoq4DDiby3zV/HZta+RLMrYN0b0f6N/H0ZNtuV
+BPJNnExhd3aLUf32u47C0T/xShsJJiNFxzk2QcDivvOs9v0zueSCc0raZxl
eDDNrQpO0/2Dt9VLk6OCw5PhMDuNuPLkV8J4J9lX7M5i23cU50DpWXJHqp9d
TIWwxBqLyuhVHft3mjx8kHIEgLzVrupwjsnY7FkUlVaH0I0NHuiiZhl0DHhp
DgBr9Z3LTdfXLNP5UqvEAj3kP0lKhK64mulHQkOdkBFL7lKYviDYBXSgN5G/
uYiXPZmgMv+weX8qUDC4mQugQNEHBw9eXUPQJMzReZ5lO9YO7yJces0PsBuW
zFVC3InfhNA+4dIPN2TtM6D27k3D7qtLOtbj2MmQ12bIDtebYWtKyLnVBUrz
qybHUkAZtMTBPLXSf3DhzWcLPWZZnVXDn3bkFRe1rxaxtPE6PFVzhESUloUI
qKXmrROgXIikq/cpqQDLRGVVm8jsKokcV7286+9tNBqjXHuUG+ou7vdeSWpj
2lQGpaENEgvUSbtKaMkrn3hIvu8cSLcuaCPatgD2PZ8KVOWF1ijYHe5fD4X+
vT2YWe6zvN4WfgDTbQzWGxuoSGx/+K115ni9wldP6RTJU1CLqjs/wUUsWKTZ
f55jIjt8et3SUKU9fGgcI74548ApkDCBIksDFm7m0Giy3wkd3/Hs2CA//FDZ
7AVNknhXmLhXuoDDEOVmBhNI24egkFEj3GSiogFE4BkbyRowvMrnfMC+DnCE
BtIa/4tQ1FwhIa/ECQCRycY06lNCFMpEcRFVcs1WAqafc2msyp3RUmWPLFwf
jOV2oDsaDmwHNf2p/8ugq5BWoefvIWLhB5KQgGWuO52UCSHEd4RLh/YRFKkB
Z0PdehAMmCMAxpEhY0T+oRBzD21Cy1w6xJOjxisgSKalTu4yFskJWSmhA+ak
+6GlL0Pur9UTXCBRTwSY2D9fwpFumbiY0gaDrahLoiJwIWJgoZ2OcOMFxN/W
/SY7dzhFAu2rp1hDcp6BEi76+vfDjXvRfic608/Np9PfTNkiBMcyxIE+nccZ
qJH3C1McgGhmOZP6sHoXnJBBVv6cNSu/cnw1KUj919EeIklhCeZsDSeIetiE
JJig2CVzCMGDZvxh3Qy+f07gtsNM/P/tsJHeP9zICNOOoL/7v0XdxtHzBhSO
XO15c+7uHosDkrFhfkTONAMLh1foj82R1sIAjKReeEtKjs3pxtzObsj6XcvZ
n4XahjtCrkpwWOZm1A3dp2NSFowA3FK0ejVnyUB4IstJjZArTn2IYCoYBXZe
8xXx4XwmQx77uwSOuzGvJkrmppUh1rnF2emjFf9DyXleF0ANuMHQWXv9mVhG
MTLzDmEmFayhmeb7rbKvnmZUff8PIT+qhXYPFM02bAUEkLRLmetwLeaAK71N
cScbRy/ekDs5MGy9OpUlRTz1PB8awbDpfU8SPlIUVDV0QQnaQyESUORLWFvz
/fDn/580KVBYiSQotLqpHEjQp6ms+cIomVn7/qRMe9URvZOn4y7eiIehlZqo
kRZu9YPcZs04KqMqdDk4oNt/lv25OCdhj6pIqHbxRB48YDLvIF8kymgjZsk2
aOr3WhD15UeVJCQ/wwcYH+W8JA6d36SPmDybVECTE1+liBlhiozka6QDFeY0
dwuwGgqvGtrmN16y67IPsoJeaIaAtEjOs4B4k1p2LWhyCNAXBEqVD953gT9T
jWz5OVhZKoXdx5igxp3QeLh1aUdOVksaSX/geiwfEVO970QQEn/KzT+GKleY
mGpt0Pny+q9yLRU4+bLF/g85DLLQosTDaVv9dY89VcRudZC4U1rie5qdua90
rwDBgZm5A8swqo506iuHEOgb61qOgz9HQ7H2cwTbzcuYulVqZu2oIm/Gd5Sb
ix90vO358oncQOiXo+wQOLnWqrk050MWwNLKoQc2yX4lb/f9BckvFFyPLbWy
Uj0IWGdVpCOD6l8epWIXr6Y1HsknCmOC/7mmj2J5VK3iD4dv4Al2X1zqIjaH
RfE8o8kX5c8mulevSHqpfZm4m0fcql6bLqbqiR2i0P1TNJzr7MV17KzGU2Mu
z5ZZSh2impNt6/ft5MWRe60TKiT8XkTKAY0uWyinYa66o3ZmcFIcrD2195Dq
fZO5SouXIo9FIhEMqt83ooBSJ8smjtadjbBMH/azPAgAGIUee+U4somDfmRR
3is9ojCA7c8kAwlEwvPWe0RS8xY2KaddwiplkfkSsuHdGmG0gSQAOKb5igN+
xR2u7EMr0QyQQhwDSVF8FGzOYhPE5GQccqw/s/8H5wKyCl6g88GS55PzhpWA
wyZcbfRGNEtlGs0eAv6trLmmCro0x3kGwxngd7sqIDqSJRkwWQWIFz2WqcWI
SDgvOG566AjRBXF77XU8VvYBKQZX0ieTynSt8QFl67Qz6L7HxMUPBrKe+K93
+UV1BAjS57XEptriwlpyZHAA5hHtBCgej+T/VUDh8mDCxQihPlQWptShnCXa
/+OKPta0GYBuFLIJXcmIXfUVE14bOr4OEhEWTqspz7dMnUBUl1UOSc8BlJUl
Kr31cLtGa/nalGBuTwg8BISJ+0/hKisTVc4xJAQxvDmG8EcuHLeX7YZc1bP/
uYqVcDF0vvA1xVLBAEigDPoB/JwQbNkQPrcFtZRtneoPD0480WDZqp9HDVDD
OBMhiZo6LZdcLm2kyrJ8kxdEUPEZoQ83ItEe0k7doYvaur0A4PWqUfzZ+qte
CrWUrhqV9H7v+NRcku73UqAeA/obSHHgWnLunpey2cP2YzWcXaQc6pP52Otq
nTjg2D1xze5nC6hPujn0vj+TEjL0BC3EjBr6zqyAUH9VytHMo5vJuzEg6omZ
i++VCRIZVNiEBNpuct/NzcINioFUrlV2NnRFpMP7WXon4a25mFY3OuMLbWj+
SsyxJoG/2i81GNGtRykAVkMyLEaIZMMd1EPtan0XJ/9ciJ64S1g3d5E/og43
t05DXkcRrpMqHgPlXtE5eS/Ukjwv2MDPMR0Y9yOnB7nPwL+K1xNYuhhnG05Y
cxPuODJ2l06xasKzXitC4/VZ1L7FMg9qesHp1dZx4Bpfr2Zqc7+JZ/PDy/dK
9CxRksHsUoJ+crF0Hl5+6RB2ogn9+WecmL1EeXL4u/NePNAa2SjHm5H1gGdM
hWTH5wdRF0Xw9iKKnZnIKK4WZ6FJ9UZhk5aRjOZfXrsTvhtZujbPsQP1p2pe
15E7Km2toc/WI2eZm9b216ZM47/nWvGPKZ57YWuTWajvNnKCdqI7675Ta1Ov
EUCs9aYLMo3mmsIhT44chzwNvF8cs14PcUB3ImV6jb1CnfoQ0FIBDJSHKUYV
V6W3s1767c0/3zcJd5yboyrD2GlGdlzSrimL8Uw/ifUbY5HKfuKlvVKvBDep
p+Ejoiw5hsD/mbW6GpXqQEtBbc9KpXi/bDjGEYmIy2fFBkDZ5IW7XIIt8rE9
aIdgWrYMhDqXVQkhDFe2GE17snnDQzlhXCYl1Eoec8DtJot7W9FethprAdUe
1ieyuanNTM5oIe4Zd6SU7XddsR8+Q4WQHSf08rG+w5soAgsZequrWR6ysUu9
MxVPlvjrpzyUpkP1dF7UYH9RIw1XXsEIWv9JpJ7lCC+zlDTdCpmPfj80grT2
aEvrm41QkCuZRV7USv/cQFs/GUPYOVV0lSfYGSgHXqGrWJGIM+i3CwaMnxls
l3T7ePTlwOhYTZYhiP6DJBOPifxLQf07gJxtFTNaltXLWS8oYH83EZ6ZqBep
2Fo1t3Bp/zgvaUBxGkoEn0qIT5DeaNk/DTtDDiushmdu23apD+15Z2n5s42n
+fxWmpBQwop0I8edAVMvZa03p9JS+W94eGdcav65XMb61+h0rxoegnpedaTK
/TGvuoV72m51CJwjAcdWHjKnRk/a20HWpNE855xX7tJ5sA4yfYLP8EvzxCSx
pgQiVg3ZX797mWIALBpI69vGWxN2mmueJc/7124EWbfEWvYpT0Dcmixax7wp
Qi0mDIHdLmJgRr2f0uECLOTK8LqVif0S0FZYFVHqG7c9qAjN4GTykKnmZKnN
1g36Wgoz/BRRk6L8IUq4JWgkSVBOMvb3F1a0I5tkBfBBNyXoz4QD8hjy02/z
2Sk5G+5uLFlVP6gvaaMyiIS6II7737yee+5Zxzc8Rjn3Yl/gFENpw+5jsJTY
2IXNt2z/wwNijkAxOKYxKmBSViT4/KXbh/wWjgsJFcXK2n3hf4V2w0s3jSkF
4XgpNF/BSLfc7kRrIZTHYXM7fXqVtI9jkRHiJQAu5KNenSh9ZGaLiHipRDUD
XwxaekOErSGaZWT3tsQ/emhcl32zGNmJ+en/pB9Isbc9Akll5hqXr79d+T4M
JpToT+dNrRY787PZsrdGRp4HB887qs3qQeUXDClVNCJhEM4LtPVS2Ofn7ycm
1HRHd6MnBfYYgM9JLfZObmUJ9FMT1zRN7o2Wyt86DsPHkII8zBd0CrgtQC+k
7Q8cXoJQJRxsb3YlaaKKRUzjMfuuaAru+2t/LJSkD6c4r3yjVuYHzBhcq8pL
C2qUubHE3+WogihfjpSaHHRM6CYFfU+QnqhNwsF6LVIBS91Dj6Nx4ZiR0siA
Ys/D/XxyC8QtwsXRwoVtL2eyoA58B30s/YyRAQq3HzKIuMssjepeD2mIqBZG
VI10cZ1G/FSyQg2oj74pgXpCYv0+Ca0uikH+BZsF3oIP1dOGdB946bEWJA28
Ong7LqykHFiyleWJpdZ3gwBBs4czKwQlKNFATGuWxKLIwkJPi6pVujEN3Bm/
Aj9n6EjE8Yr1fTweYzPUz4M+2VudciIFJu2IeIJhjvhSvQbCPwCfN+MBHSV0
PBGqctLn5Fsp2RFr4IVMW9iuVnTTOqkucxFqK8JDtSjXxi9nkyVnOolimaX+
g6jjE/kFAfhLnkBKoY5vQ6ScmjjKz+PQV+GPrNsZj9RcwAZjBwdlwiaMFaPB
MAxyd/B4amjIZPGgq/zTOCdHH7CRxutsR7OAqGa6RaIRlczb0ZcazDnDTqM2
KN0lbM5PrAgqoBl77HxZrv4riU89RhhHrDZI5bfiYhB20vHLQr8AY+UAFIAh
AgIcUwkUwCKfw9CTCt2ql9CWI9N0RmzlBDN2tz7uRqtSArEpxJhF5mOdmQW7
vz60tKOrJpZ/Hya6zPckTEzZQvNsxe4XQ7l8pBUkDSL2zJOCE+pIILcdc/uC
v3JdqB7IHb96CenSh8MMvsNLH3X8p2cQbu9MHMrX5g89xPv5AB9JAYMA18sb
gZuOnRYAM7RVdizrmXDp8SnCEGSRJXYVR23ElEjnyTqFS1yCWvLtksFf1Lui
coaF1/KDDQKZjfljEKDVeBJU+hMmyLS/YMdb22r3pzv/M62OoWMUFcgbUFDh
paGJPCHKhrNy0dLJbSowPISPN8IrnZ7w0vUSu40wPgmyrTN1ydSukWsbOL/r
GpRPxE+p0l/2qe2QtSlvYnRzh5/vIW8JgEcwTBjKO7QWycYEGDlXyVDgJ2VG
dX+K7znSx9AZr3yWkfAJ2EVaPaMEAra9qsllAyjkaznSyoL12JF360THLyZG
ORmFwQhQ37yBtRu1/q0H3LA4hC0OGvzhfNexJ6Y9ugFRX5aIQZpohgKscD5K
fxw9oFIMrhUQMg2XCphpsnjbZzPHD8SzBSS0mbmC67/eaNwNjbP6F/nEuz27
VB/IX+6VwcF8IPnmNmSA+Y6916mK4kOFKluA8qQxMj6Dan/DAJAVA/MjVGg5
FvTt2CnpYmD9dqmM89Owvzvbcv2E4qdBvjBfGZQ8FWrY/PH8tY6YATgMA7Dp
U5eJgwEBih7zZFQiM1jj2BNHOYJT5x20IfDpyJ3Yz6K3nEMrwYlrqDIOEOMc
H3fwoZ5023VhSz9307ln9+j5UWhhbRZoxQMBuiSsNHBLsz9xlpPqaUPw8krD
frjVXk0uQeD2+yiNqUTRrTS2hCeW1zu73CO774iF9pvOZso0JqxUOCudevyi
GwcqOzCis7xdev2cKJWCCMJ57WLYVz5Xsp+GexIocKdrbMXahd2TeTthytD0
bVfaDxN7bBIqWVbtJmJ/iS3Oj7d16MgnGOvGOZuJItWHeOwZpv1nK6Pwpeho
iC5SujO4yGx9d2QZBM+rm6VsAnvpppqLr+hqbW0qLSqQDUg0u+ohV4537H5A
hQYRpfcnPzcBLhBHvLii/w+xWj3eojxVt63ADU0+TPzuwYz8RznvcPAfxlmw
ZrtYQLBRcH6KxO58chTSDu0DXNa1RZVzK72sZ9/UaBqzKqM1pDqaInVRaoCh
gdHFCkbSA1c2I1orVlK12nSmfnQ0tpj4hf2oBRso/cysM4VzzgEzVlMi48kS
Nuh0PPjrq7rgCw0XtUozyZD5kRXjyB7JtYfWJYsrjtS2PMscTuxs+73aSTBA
BUgozLXaIKYwMkXv++9KlQDdRKwIrW3VgfRiGAJmE4d3+e1Ak7bK3CDE/2BE
JLUP91FpIhsWivdIL1UUD4KNDJSsyeDz0JkuRR4/OTaw4sv7ljGOrf+ZNTRK
ZbK72F0LjT3f45AvyMfbgxiSlGtZsGgcg0RQ1rknAiwq1w9nFtlSB0fjpe3B
cwrj0mSAjB8suX4GCmF9BhkF4jiOGVq953yLOZFtNa9WZ/ZWCMXn4Pa5pr1N
K8xJ2qtx7Ul1+f4dxnoc34mu8h+b9MO31qjc9S3shD7z0trEGXV4Vzh6zqeb
ZJN9/x7H4r+E/wxt1PEvv9KDq8qGZKW01ndJg11RnkdenoggCR2fAJKzJDlh
6131OVT/5+sky4Y9gyCLDN7Fk2QSjDg1H3khvoZ23IPY2xrr/q3GVJbcuTsP
7nhXwNlsEsO+r9i/DW498G6BqS6d7pnUKCXzK8AMAjVwJLWcJgqhS28a9RrR
cUYfk4DtoMGFymtMB1O9g/uIma9UQcpcnpX2TRCa8zkjo8H9ttL724C4Qgnc
it/DR50WEjsPPYxy/GobInx/5knOU3iEBRrtnQucB2aYeiMQI5F8XaDJUlFN
vH34I/d4oYcxW8gABvjeRNulmHRh+dqXYjzlDxllJHulBjULuzMUMKktrxne
VEZ+G4bVN1iCBnGKkHGFP8QDXmAvVZ34AYUxeOiogXnab0QIKw30XenjDLoa
9Llp4MOEUGLTR12UdgkW6feEkdIAnRUF1JvKUxxGZHlua1H1C7TMW8lw4Ho1
z9kdIq8h3HN6fDmDJuSglfWFyrTyK7CLPBaW9QlBjsQK1tQLit+ngAuuSw3F
ECedVP14iTS6vfnjz+JNHexbw2ewHMN2RML5N96GVAmoI+RwO2rZTA24Z1lK
eCLwnIF3QFFiE+oOKJDn+VFbJDr+JIZLwFinv61xeK1zGUxgvuBCQiXLdZym
SdRTIMhjxTvTSW9h1hZhTHx+qzlPv7JQ2RhDk7q7AE8TNDcHzPHUr2lto2SE
zf03RgljQGDczvzudvD8AMznQbQRy7w9Df2riRHPeW27cn9lpQ/fx6+5Xbl/
OrLaXV0TFMGHgabRq8VMJUz3dzGrFftuPtSLc/1Kc3cnWi6zJfJo8vaMPKNm
buN3mkGuUzff6+JyZjz82i8jBftc8y26P/Y2k/JJxurA89obBwJY3HnCR3ww
pJAZLBV/KJmp3Ph6E2lp8g12TPDYwQS51z0hf+Lx85XkiIk5MaR7Oa3ZVokn
20WBP7MNRVRzmMRStPJldGlIxaW4Md8gqCZ1CeI5/pkc4nV5rGTSeC8Jikph
mvIel3eZfPYAOUF6e4hMuUfaYUvv8sO9Ywk+iRu5y+0g92xn2McmTNkrtCsb
vbgD464iQJ4ipm3/7datjGCxdo/CWGPGswacOIH4+AUmcN3asfA+VRg5ae+E
e31mJkPGh2sjQ/aWIundtXav5pmuje412k3CTLkrCgsqPyA6Xzke2tjGkeGR
sDC+3uP7SHKA2yn3MYfFxI0pcrjExi9Hp1u3SEMIpZDiU13kORczuQ+ztvi7
oYWhuPT5PKNchar/PQzmPF6+4wxYaazktiV3kRKepl6/FEUzYKB3anykwZAs
Vr2cwUAJ+1tpYEE52tFr3JwWxJ9SKl3Xn7Jtx1ZXGGzQDcfWMFnYaUu4tclB
5NbTxq8yKd4w7bj6/AEYv1BekuRZbH6UNOmL6VIYRXbH/T2V2lCkLgYZHBkD
go9pLNAGvgd9nx0QidWP/SMrsrCHQhkSblm3Bc81St8Sotnaddgldzp/v1te
Ri3mvmWr8m19bUnUhakHjN4WDdtQVgzJ9PmJCmiBTzNJ2JlSuPNmprf6L/Ge
4pFX5BMXvKpV9piEDNEfx7O/UNcjcZYppU09Mqw1P/zsogifKfAqGKra79dK
e8r0oGMUZ45uVIOjR79qc+Vvdj3FAL8vHlUPM21AzxeqP5euY9s61MNWRe39
dC3DOpL3TZtl247iziK3lMj9uQHYiKJ3yIdzR0RhrraKoArxOuL1dx10c587
MUvmz5hSi8kATy2xjmbyZ1Jqq0KEe+lr+GM7luofcxD88Xgwlx3oUC06H+Ex
tw1VkgNHQ2fxDKnSN1aZ63quSb6VIB0iT2pwAREjSP2g5npcQEDgUpU32PO1
gVTXtBV/cdA6driSqTJsVCekRO1Sr5Sx7Bbs+2AwqeQPceFY3bdeX8dHz/iS
1cofQTdDCIZ7+C85MhPKF8MTiGU/PJBtTUyAa99b/fC7IOX3vzsbr6p7kBx9
1EGy5IgKAGtQzPIlSGGneBmHIaOWZo4uAfjZ2C4MV5d7OoVG0KQmZLBVwsrY
lk58bmoygofGd5w1tyS8JttlycXUiZr2PofRsdmwOVMu2TvV3YPP3zstcY4B
TBliIYSJ6L/hqOzP1oEgdF3FVq2iZKAKB0ThBUTajNdZfki4iVnEZmNO31hJ
iUvkrbS+mqCovCvUpuXmkPWGk6YzSDn/PiO8McQDaTgRgkZIKoZKxzB18Rm8
2E0US3q2w9fODDa2IObtfljAhE+i7KZMHNfPiAKNe92OasK9eseWpw+LeBmp
/kcB/PwU5Nc3hTmONXnqW2CXJf0ZWFmeuDu3BhzMh32P6K/jyVOBFEEkXi3w
Uljkq8oNy8bmWmWJmWz0GA9R++OQXmtirHsxe8pzHHdeV6EoWTB+ujLqRb/8
AOGLO2eaNm5jru4GvpsBtCIByIaNWeOeYN0fQHv+9I3jUlE1Oc0ZVBEdX8tX
luCuAvV/68kO47f/eXZvluZyID7FUnfgJgbreuxYFfjMMFtGnXIKLt3OohIL
mCLmq8qBwK+BGoBfq/Ek2l49DTfJNWtmVHw+5pqoiMPtxnOQKuSeEwolCJnk
u2JieRhpxZYfjNEHcF6fDA93WMTNiozaflH8v/HhCzrMYgPpomyleBXg0NGK
UdjsgWDH5oKfmUmwCOAqzANi7MDbU8R314oz6ps4ofMnvJoOaDYxSijQhmIr
YDbmgmD4v/gfO/QorsC/WEIi5nrsC1pZ1Z50+wcNxhIqARFUq2TrE0r7W8N9
xWnE/DfaeETeVNDfqWeS/z+7lUdLFem+QtcAhgQ1J4CPTHLnHIjrF0BqXtw8
WE/1YWfKAbrmWSyOKXe1xnbbnHNSuEiyImVPmFI7yqWZ7w/s6NWA6ENBq7aO
RcN1L7lqMCgpGW9gnriIy8gLCRJh6uMDSbI/fvIwB1UOcv0Mk29L3OgM4nVf
SjT8frsQmRstmhgQ79gvealt1vYQXYZWpE31KCLCzGzU8sHwVWbz/LMZ2dcz
FZxV1A4gkGbVSwsR/LG2Cs4bLpFaG7uRRa9q3P/h6oON6zajC/GsydCsckVQ
ppmgs+dVeLx719DDqaVUnXD3xQvogo1RHG5MEMyW6/1LASjAe0v8CMsR48Y1
FyfHfVShKnJvN2rRc2R3LZtXVKjJp2JSgevm6L2bR8dKrB4kUrG+5Y/hGHlO
z8ulAzjwruIW/qIMcbUxKqSHrhub23PEbW5r9/9AZX8TfwG51rKUpdegESGB
Zj47r+zgKEJUIoQt+BsajtSd2FvRz5RUZdwEyQ1cKwBf0XG9hVYPnct7rWJR
2LPi8oWaZ9GuEV2e0ZNItRTTdX17ySuxSVGsYoYTj4ShR/UQ/iS1b/VSm2MX
D9aRxIzrK99e+7FZJNNODvo+KIrEBKvcZJKzIG+FhyJCIShFSILm3xjF77wj
P+4YUbIxT/c8BIS7bRwEuHSABOjgiPU8Zo3fT9qQvuPhpHI33P9FnqOeGOll
KqnGNbeielGX+OwpoRJ3yjP9EsLr/yG8YekmXB5sd0ZOWOGbLVR76SA9qduW
wcdKQVU7t1BvEsA5psCtodNPJR6Xg4tECwsJarCWtQLsfowrNA8yXmJsAM/W
H2CH3TdM5HUvyFyuIV95kFLPCt+v0JiLPxyLaiYynXAeLIHQcrPKr+8uUx7B
FozYbwXNJ3Qs+GkpCs1Hktq6NBtiCQmv+DzqC9xSyYeQcKPe8RtEzv4PiRxv
Q8fcehaRbpFza3GWjN7fVbkO22LRQ74wJred8X9fIxps72QCiZKNtnbzQKG4
0FDu/Zx9EcVlphhsmHv6K3sSbcqIh0vhY6XNBdap+vpiiAcvaF0H39cpOb03
OBlBDxMNaOka6BeZwke4jE2rZHjSdgh2eseo6B5M8DkHIRKnx4wYsOh2TLHD
kLNq55lEMWd+jSrNlYvB1RuTkG4QdIZFZmkHZZh6qTCLvmF4k3SGOreBnro6
JOgj4H2r9SoiCQarEj9KBTb4SxcnD2y8y8Ixd1b9EflsoWWtN2JrNbxp6a9r
XpSVvVYjN6EXhxdGcEQTMB20LkH6R1BijbyoJFUtJi8oDBsCkXyh/BZLv86O
FdfbXwOg1ybf5WZrPjnNsQqVUEZWQJgEOWPYA8daGP5Ey1bYuMafaSnlfTNG
jNN3kXez/gvoYt8rgx1ZoAr1mmVmiGBoeO9O+QOvdUovVLbk2kmt3tjzbpN9
TzT8gvryWhxB4lFGbPnDyqPEr3IFWeqx6iV0ddy9MmUM6QVpec126Amn+CQI
gnPOdKcJlxrjKnxg8TYIymIK7p7Ve4wJWJHVT/B6/SNsMZxnOfq57MEqoXuD
Yg3s+7GeSVtB4D1hFawcuZHe0KWw+k4ctmsFbY4pGUS/qwHe33gKf3mnNcZz
vajG1P3vZLqqx21NSaHmm0sOoMl4AbQKcAZKPA5J/LaUOSu2IDrC2cw3V6jh
FTCFYI+Wf+knH2xj6UbnHCUSn1xVrj/cusBM+W0IaC8+H55EXKW2QmmD0J5E
wI7cZtBGnGaeEi0PjTx1KnslB7Uxr6bwJtUfb+IM/RcMu/IzbaS8D4IGcd4F
LX0Xx9m1Hk4KqcpndXeFlHxUV8eTR9jC7JTaGwjmJWADRdrZI8AkTNGBetwF
hx7cOrpAEtmLa8Vv70/3qVI8NkG6ePyZoh+AIteNkyNNpg0tPf93f5UI4I+r
GFoX+P9N6dvQmvZOIF3Pj0jEHLbmnBONcFC9CdTARjIQ7+/8Oq+KtuLTlW1B
Ymqr4lJobtFTYpB/TrmVki8IMiqakekScwyuBIMfosAZ9DpDecW9VFlKA/17
12MTpbhyvtXF5qeYP4i/mo0TfbQCPqDSOXe7FYxNAUZpCvC2HDEJunih9Xcu
TEpOEvmLg4lxUnurNbrI3Ix6OAcYuvuCDZ4eBuPZWz2W9eLk+yfyrNb+4Nwd
LeN/n959Nw9+7ybamupypom0G1wAbakYb8BGtz283arm85pBPCgZhptuem8j
9TWtGWjR1nbgO3E+yDpbEuAqz9YbqalBwaIQpkFPL3CIrHK81jTYrQqG8xdR
Tm7fAIItGAcl/cEVJmNEC+XdiFAZhqfn7J4ijutBa8BzfulEyc8ImQEZahlb
ICSEQUTg7gpc4Mf1kYdcCu5wM/S1Zw9M+np2qZmIzJAwFzm/PgJsibEmq/di
IFd9jbKFOY9LHG8AauFohBFcalnT6q73XaaOSpsQkb6FNxhLlpehr2glhUnr
VWgBofImGF4wZt4W9o5k0Mnv3QWHQydgUD+Pn2Q2erFZkFCMeEAb+pf17gvi
IKdZUN1jMHao5ZS+XAPqbx8Gaq6o/iIin7KsUlHpMdRURTFsBGpBvfNF6ml2
IsK/VFAXPTJS/wtk/kEMHakSOK1BC5pEuQb95Tnoj2Fl9Jzc3pfOXfPWqLcn
GAq5UBBw8glIdaIwuk6uLHjiTCkCDJdX+3LyBg0xDln5q5vII1BsYmm2hgWC
uqFnTOopCG1ySZwx2zTKGf4xmw0sKYbA0+gtR6di6xRP9X4ZY7laC2oq7ZOm
QMu47AIWizoeKUPDC1njy9o4uscfKTNWgRBRXJxOhLgMYxA7NQJG8PcaaR1j
mgQA5mP8ydar9bexDSurRNF6WYZX0i2dTvSJiCLmnA3JS8AHwYI1lTjlM7H4
r+iZtr2asII6sQT5HTV7jjhc/TlbISyxFkVzoiXjRDkGTlpbWscf+PPVsCWV
YYGPWdaub76e9idFcfWjoTUCRCj9YD6feLF/kyKIs7T6IIj8FfZd81GIZ9L+
vstHPbLXOLwa99t4MxtkryR1sv4/SQQK44HW0HReyW9W9VTmPdnYJ8lVua18
R0HuOb6aT91MJFa/ZacI+GWj8GbY9rGkLfF8GIthqcuITbJ05QvfQakP4nkT
AatHPV+YS1VQNQcuaiksjm45eb9sHsapa0Ga6DjxObl2gn4F1oLpAJGMwW/w
MNqkwVmdINLQOfNK9VK2pqsN4CpoRYzGPT2feGXVEYSj0AeTFXc/IP3CudbU
bWZig0X0wvSyjYk5jqovcal4Z0l6F/0okvc5gHlgg/AfVwiUdONzmt4fhnLr
6lVCKnGz1c3Y9UEPsV2Gtrxz8Zd6cPpYjI2obRypjUeY6Yxh8MDfLoTUkxIM
CcezFNwKPMhG253+N7usC+x5cjI+bMYl0FzVL4d1Ist5G8vG9oloYaRom0nD
IthR748HTjsxw3ibPfKMiM8A7JMlPy+I/TBf+0PgA4oEXQ94AxrcUVfLyIGB
7uXc4es3PHjLPEAxk7Pl2R+voKRAbndFq+qTB/LthK+6veA07ZRIhkong3vH
OtTQgC3II1gbmirqbjwhRv489RF4Wvz34/rLW8bpJAcfZBGD4cLTnnU3XoxR
3C7ekB8mb0EkVMpY9HJA8c0y8+xRIuKAvfevVvQpgOFZeV6C39vZxszs2zWo
mzyy/MjG4LEU9oBys6qRw0rcfBgssMiS6pGJ3cTiouG5ha1J9mtPayJaIvwe
poyUn8EvVs7L0CH+tWoyvV/5Sm4wnGm/bh/K8607GzsQVFs7JCiUHxMYx9A1
BDBAMvcp1qSVHkRhzMiRP8XuZQU6lBad3LWFmB+U5BhpYfFnjZpsc58+zL3A
slYGhXc07byUH0U+s64XYTmVr5CCdnDKsz60cszUnvgUQV8L8UFbuE0v4fAp
yOePfwJCtKfJA3TV20oLXgsAHCfN/v+Vep3o9DpTwiYAqqL8lI7jzBL/Wzdt
X9OdTwmP5p9wntV886hnodEvknU/v2hlQtkC14zsmbapuEPoEMxRFyu60QoQ
6vJngA2R+mS7IreWZdO4VzKTQlNqGnltHT9SEk6HpRcndT2ISJhawj+bWgPM
+GrWnZUNyN/WmwmEM2mDfsge7XMiTnPLrRL7tTFZAcneiYBVD9PKXfKspdzn
H3tDkVVy3nXRy4R7nuEWl6eYVojqrGgvXysieUS6Z0NVaTrRGSJivAG7pD8+
urFWjtMHrE8EkJcYOXB5IukVvpI0craNxmNQVITWdUGvUthd60nWIx1xyUuP
hLrGf+fHLIX1BdX8Mb9s4ZJO1y4dPMGZ95XUPRTtyqSjwjyQqXpc3W6aXRM8
0x/oSTDwlg90C6tEljT7rPN38qvk/Ops/QVKz4WPwUpOGu104/JyFIYe877W
u5yyK/fCZ/u0q8L9WvpZv5c7UgZ0g7zP94SHb+p0x+DlwW8SJ47Z7OWuA54w
nvOv88AqhKTN2PStaQHKjHYID4/nWL7XdUkzzk0bw7NaZRBaCCtVkfYMEc58
J6Wfa/iF/YB/H2NZQrnM8y2Nwyd8i04vgR+fKFZ1KZnptOvJeferHJWRg/P5
FOVOOVYfqZy3qvnoPMizUTDn0MZGHY4HCL7dStpPS2hp/Ij+88zWAc6qic5b
RHhY8UtUYHcPGH1djsaK0e3yonGkPYRYQ43dRt0hJAtt7kMZUkZ+XVZXicuY
y5LcCwneQr0k61GbEN3RW/AqHoxMcQfR6DqVvN0FnQUdYTLaMSbPlYMd+1vw
d0mCQ15eHKu6TRVZsIMqU/btiFO2R1MC6Jvy02gTF2AO3rzGSbYSg0XbI0lt
d4BVJFRQ6+aqRLh6FuJKYHCjPRJ4PObYr9BFXXB+XXotH2/hZo29N/8teHRv
xfmhM2YlL6poKcHPIaXCgPvTcM7WM4Cj3On1TWSV4LXGWhXS+FXRKKMzX5rT
4nlbaYTYHmh1VCkOyoZrw/F1Hckyd640KFkJ2eO3pthsdsEKPK7HuXWA38fd
45/WIvirImp57g8hr0cwcUpArWmhQmBfxC2LNU7CAD8dxnCFX2zob6T8LlOp
G4uuVNp6DNhsWj8onywTst5IdTQ8cs0fR1GS6+BJLG9gQKVm2HEDOk84dwFO
3igzI3VXJUFS45KxfCTRd9fv5zpkj5ZFjVa0w14clz/MblH7cZS+qBgCbfNo
y2kHsro6veSXrtzCwV6GYoRLAffDC9s2+3BDeNmQhRraT1Q9S64LbXdjcazQ
KTnuol2NMVGi+IcWW/4Xc8oLtrJCIKcqxbNTrWhEFBCUSPoQIfaxzYdKgsL1
S7VNrJIYnRT0HBEhGxBHIpm81qFnqRl7fMUI6g6N7YaIKmcyVX7J0Xo4YIz2
ELtYg/4d1VxFrdzppjL7SOdZkM1svjm7XbPrT4Of5waohHjLDhLj7JRJUCow
lKekTo9XolNDngeLIjzcNtAPpa567EzFUu6qSlLnZqRNEGSY4fBZdz9wpW6Z
8vKMyqnldnmfO2yzyhQaogt+Q0cmsgEDZztpvrQSFSKr2PstVmYveKJqKH7V
ov3njv67E1rzBHVvOWHf6z5PqLZ9FCfyO/EDX00nHZ75LUpiuxBoxpjFNTkG
nBrkRxWiFwkmNey5WX5prCk5kTl0NWAhIDp9Dv6wiYG10ZysXxykVGg6iGal
5zQnwlZ5/YxJ7QOI6Jgdk9IPpAKBMvvHOs/Zpt6HW1tQBNADK+9QNHmRxpi9
bMUtJKBAB6iSuKXGVPK6lAMso0vALVEUbCp9RBq4PnZMAVqVcs77/5xyz/NJ
OCrnks6mLVNALBJC7zNQEiNbpiHztcN/yHQNM9KWBV68MmkEJB3q4DgYvuTw
DnBqqa1Ir69sh6gO5pDbV31N/3avWotGTzMJ9EPGrf62UxasjbG01wYTK9ye
qS/uvKPL2wsrH+Y66ObsKya0+CG+BinZNqq/fU9KtVLTdt4m2alw+gpIaANq
AlDim/kD1I3BOCVUUyxUzmlMgOKKBOl40IZvCjd42LgbCZsXwXGysXzn/7HY
z7XYA8wzEKmUkNRXau0AE0TGO3CObkIhDqQkAD6YF1Wb4czpm/Z4dRNwMTdT
RkyimdLoQFj+/X/b0IEQT1t5/CSygKERLF4LYJp0PveNU1VE/zac7BG109AC
2rXji6sKiHutXuhI6EMBjlIjXoLE54rsJAmcjs294br1m4dtkeHaXVjCBebM
NWD5+Xu+6x3eNGv/oMjyIAFRNq8+Kxme+MPZqk0nc7eZ2sKm5b0HarQF8OK6
/vv89XMfXMGBRSKxDY1k1AWr+IezOZ3BzrsuQ7A1eMwUjDZkarbwH6paAy5r
a58t62eVhjr9XabVysM/0OOVFzK237bTqtKzSss3Bh/aZlcYFWX15BBhbPn0
gKKVCyeqSknnDTgLRGJcFFclGNgtPYPsJC6hJg+HtfxoubYzzVSq/B5cT2Ji
m2PwHDrNr4rg7mcr8dJk+WNNiUgdXcia3g1LK591ZujfbU5OmEqS8gLvGGF1
zh57GmXZQDWIpfEXAlf9n3Zq/SC2/tFjDVzpvQOMLOItCX44LRvaC5YpxPtY
gHlESD6KdzMtRpJ2DePcG9TRKM4vEGyIS4xrHIwDrQ7uaGv3boMNssMJuAwq
YQo/MlnlTKkg5rnHpCwd4nEcoB2OLlIQ/W0P+7jHPOYVt6sb3j61BMaZhRWO
50fst7mpeY5V01J5172JQL9MGJDkrq/snzFaKG30qSF0H67VWE7S80ic00mG
G6Ff8vsF4YMsdLEG3umc1JEI7M1PktGJPshXIjfiL3dtDwmiRqn+6tEX3MUP
pFoabqsI9txf8sds8zzTLBdQicKuK+76MZod5LuURN0+oBPz+MQOcObp7LPY
IzwHLMtPskma8PEBtwAnTqUttm0/MRbw2ufgl+297CiFrp6Kpf8kp76QpOlP
toMp9NCyaHJMlkrC8ljW7uPtn6wSoCDbSwY0esVUgpUkHrvof7V2pOHcDJD2
0QBebVfXx6RqRwAjE9UpS781MilEwS69kAYZwxcaI6V4gt/dA8zpoAR4hw6P
3Z3BF6zJWy5Ungmc6lVsuGpxtM9OIO4hggkJ736OxER9f0HsNkc0Z3PWRzyq
eHjA8hjjhTi0n5w5vEX+MvRqrrqqBYtCcWHmt/u6PFfsVrd0/U6o5fWAiFnQ
D7KCHEYu6bPRW8weIEI7vY8AgtFG0ELHAOvtpWnO6+gWevtyXXZTlJqWHopC
c/nf/UXjIqmbSC3vJNuiMZRzmIKNu4tMvNsxDOiASw0bTVnNBB0BLCCLi1Sj
2sRCPoEk6hAC36NJ8QzL0CjJkmrDb8sBDrGtoW+6ypWDuWWhqinMx5fbcT2f
QkzJhg6QKka6h+HPYZdo9+bW/3EUJJ27ffm/6GHVYDZs46ZLpscE+f9iJQ7e
RO46FxP4BREvko1lCZDNyDO2zf7Mqud7dHxqQbFnjcUOE+068KdCNwE6H8/Y
Xf3ow4CmjnS/z1WscSppYyQLWIbiQ+rtpiKOLd1qI8P1SiehpoyeZQtuZY6F
Gp4uefBQks0cXWiawsfsOjYNflhthRk0bchZ/ty2vmPtvMIUQa2zfJ9l5ZBR
TyDYInbdcZMZsf7fitVTAboO+czGe5lhzUTZb0QNETV/6JDt8PviD/YYH03p
alamBFuabDk8arYjTkdN2KLqhpY1Dk9qZ6XY2KSo0UI+pHXABoXh1ErgXGdP
7og9pnSM3wQuGtzrnbfzMvo/hSXEDSWElWmn182Oh/ZxjHD/BUbY3BkmkQfU
cV716y9AyuCyStHAyrA+AmlG7OMQgsDSeSL3ppienWzPCCGcZW03LRdeZaDq
boxyUhrPdLPycqt+n6ZCAo50bj0CDZR7lRzHEcv9Am14YVRChRAWFYDjnl34
YmsC2IWwWM1vxlk80s+OsGQFCA1w91FSvNftyxCYXgP7WUiCBOW/r4s7swNk
/BwErIXNZ4dscK/5X5PFMCCkPzOWj9UMTo9NSkYBcXQAWCZlO1xgt4Gpyv0F
o0/cu9CAB6BlOsyDv7bhCwGanwaJKLavaq1/r29igzi9gAy7SRtpevVW1dng
XUYaOrweB0pL5dWxJCQNUP7pmv8Gy5wkyyxNX10RaaQql7a1JkyHGKlZk8fv
QKBIzoO4QJgOoPqPj9qozhuKz1KsyUug9+cGNMKCszXL7jMbm/pwLbIsDsX4
gWTBKnxudPxDna+/CmUC5MQlo3eOujWMztedlk3fzb0rKPqXb9vPMgQ1p4mI
hbSxOaVUhAYPUXcA81Kt7sWMWSWPCtAIsOB8uaZW9fu3/blO/rru2/e/DJPK
LscO0Blyw1xl2ufK/GPtpDXLk9VTJ+vRkSYsSaCYOpwLtcQnq4kas7FqyBqC
nulUNU1iMvB80HMtsyG/1J2WfLy2mME3lp1WyGsRYtFBQ33mbMRcTBmqIBFm
n7EGJ27q/XO7/4vxYSopC1jIg8V3u1az8tYaI30G7akuSqn2eoTx2XqBJokd
tJyKiiQYU6doGsJXqxUGPmOV9Ec0PTOcEuLQDdKL+QFjzqSmxUFs+Lc3ob+h
21XxLUZRviAiFt0TFossdpNcQEnpavWUSALR5Fpl+yOWPHrBN3UrPVDH/IRa
kJ4b174FxjebFDii33eveyQPUhbldZe7A2tzym2t6jx3ihfie2yTFzqopN+d
cwQeAuXsyllpFdkbAG37YIH8UKK73erIAY2UmJVujQk0bEvYExI57rVsSFhS
zeYZ6otSKiG/FDkUJBY8uAJ812k5A3dR73GjJpyR75l/zS0p15EMdfOdviQv
ZxjOYj8QlIO0oxy539L2af7gFfQX526cgpmxX5fsBlvsuWgRNUVGs7WDnl9U
Xpp0r9xshEL/0IBhKRJ3Fdzn61za/DR6vBl8h0wDHoGmf2+xThKh6LqPo4xq
QWcawUQnShXoP2nynvc7yLuvPJkzf3vIANKzAagQNUR8fbrnBkFfVDXv6Q0o
m92D2e1dV2/VzrmP7EZEc5KifmaYcgDRRALN6dk+ZHbxJHMIK8gzjJCxSJhn
0fJJZDhAdzpYy8aTqMqoN0R4OeZ6BFznCcoxg/u/Ov/irGM5uymGo9TilTy0
NtxAnbOzryW+PtEce/Pqx3B67HBBWLrrQm06tLzFR0wDBMYSKWfSWMRLWMwk
TUpvKSt3a20mM6xpg8VKlRAlXn6qzX3xzXrUdiaNBQlkcEkUDgqtnJPl2FhY
51fRgpcWDsfxnICwpUUcNIQChpQsFYXq+9no4rBmXbYXrs8/TZFfay9iQhCp
sxZa28+JlSDXkmKk73PV8gqLwZropxxqK3rIBDO9eiSI4J+fJrtFMv9lcPZX
zYFnwaipdupHSx1LcvvnyNkYWGbpHs0z4xYuO8fwP9yRYTpJXWz7MmlYhnZS
hH2ePc+hoGJDMkFUWp+DEKOgMFwHsPPbHX77xE/eIu/GrbdtnE2qpfiXtux3
nmphb+3qpvSr5FakeSoPLFvj0zgVu+9f7C82ex5UawqeSkb44ucmgdzK4C0w
yEkOj+M2CYEHHjSicMxXSt7WzMzSjKc4m4JRxTAdkJmc4Y0faKav4BDL+7+H
HjOxR6Bk9XmIcz7UywDnoyB8N5C/YiEkgUO6JKVBTwNHb71hCa4/1G3hO4Zn
wh4MaHVkP0DaSous0+ESPnTvAIwoS6KaGtRaLXqG0g+KCD4yr8w9AVUNKxeR
qKoAt3E4Sc0yl/NV56Fw0dVSSVlca3g9jlBx3E0xTa6rIoZMlFes9EPLUqcP
tu+jhzkNPfafFpaHkZqKGfim6hjVheqMt5YX4TtpL56bnaBfqanhwix4JvkJ
HL4SO88FGmdkbD1BgWab3ys7v+FWutyE0vA470lR2Q81pFrXfF3CuhZ3ZOL0
9j+l7SilU3x4/YfqCaGhFYIi8RUVxjyfJSX80uKjIsOXf3IzcYNFGftrJtsO
Se2HrHKyz/dgL6j7aqRltflfBthwKhpnQtlHhW/YuxGnPW4n1z5iAw3kivoj
Pzh/WTt9WrhKSk82IGZ+6l3CowBnz7mE0J5jcLwbnV+FKNmvVLztfSSqwbO7
3MW1gbYd5fuKtZVQjugLB/8gQfqD47Um6B/+1EgdpZs4V7WZhJIrpP2BC6hs
zZLshCWtnuQ91rl1p7d47eXwfm2sHhXC+dbNQ8NZyQ7HHz6g5ZoQnZATw/7J
wl1C/I1HOGSBOL8BF1BcMGwXXzkhQhCZ3YTPrJnS6mjImyp+5aehjRgHMsmc
+bMnHxY6DWtCOKz8WrM8UBdkkc3vePKdcEDTPdfz+Nkxhb6EIZ4YkIRs2hjr
ef2SPn6zSgACrKyrmFV+Y3uZRLilNyvyVoldFCOVbA7TSuil5ErUClTACv9H
cZAz/AiFvIi1Pd5OYcNSzgA83s0UZovX6Itrh4We5thZo+8TDgeHL4dg7A+A
EJOPteH5udyCALgC4B0uNuUjJELBz85MJ3mXis5lC1zbWeoo4SqwbAMD0SFi
Sr3SZuX9VdCXH0Ifp65kqiwunAcT70TIlVdFIgEUmpgkEHcQKcHYlfLp5YUY
Pper6xzy+qPlN1MAwTKqw/4ziqs0bXb7EqnWVsqXmZpcni6sHqJ09oayvvue
+2NgqNnmsEKtm13pgh1+mim38I/TxPSpqFpdAbQsz24K96Ko7eY0tLszIos2
vsmuPhze884qcCtRNX0cFNZCMCw2ngcooSEHzQ3abCl9tt378gT2GxfQXO2j
GpElR5q87XsvGyEVIYBspOgC9bSvubdEMEc1mrujPxoiS15iVYELPzmkarwS
3D3JxRRY3W28Ibn7g4zgBwVQLhdagErQ3eIcKNWhRjv7ukipfRBmTZ4hSXrc
GoG+2a+NAeNkqRmKQPnjADnEfYVTEgaf3NmYCjT/7sV9jNbMvyNcDRw2lbkF
mzcFDnn2qVW9JsBMJfJEjoKICZvGxaDStST01L7AELiUSA7HAzjS6zinZd1/
hwboWF9GzL0BR5undzBJx+IWucxY2iUR3SlTMu54ZBaSMG2rn3pyfObguS4L
DEvoGZY7PUIH/FyNi8OzGIxQSX1iC89fEd6rhG4PgithqtFwfD/YnqwabqxT
royXp1ISXoLVvqDzW9Q5uRdkJEZ4XJHYG4JKd8nrAd+lkfYUhwdP7+GjF1+X
F07nikI6RLTZsTACPpKIo6Czo9lXLxskQx6xlzFhqgiTbIB5IApRhxR0F+Je
q1BNMABc+DJo4bI2kEnZ0T9NYg5sXM7rknMVobA8JNEimnQmYO5MUNqgTOlD
sQGWeyPF3SuLUePwlkrkwRaDxtOG3jHhtYIHaHXIBitS4sXf9lpvHREkJZ/S
8POU6K701tvHXi4HuhsYIZ0jJ6PxTsvIl7Vgo/mBd2wO4TnvKtt6n2d8Q+E7
9X/HsfnQT8uGtEdJpXtAx1OdghEldFEx77JE/TfTni4cIfUaPC94SkXjU0PX
QGqUKutAYEY+YNGU6QwAULEeUlVupDzOCF2EL1VuN1u/QApEIKviTIL/SdyA
JGPCbuEyh088orXM043x1wMDoa1nHIaMJy7ZR/3XnfAOX9VpTsAafHfbmQ3/
Z+svcWhVaw1mlM7Gv73u+h6k/bY35suzEnFMakOPJAqmCD59C6AXQrmcWezU
qmymN7kq8tnSHvJMHqq07HSP5a0klaD1p/yk5qQQXvGjPkzbm2pQU43U/go/
soWMqzW+Lkui5aD0liTmVWB5s0nOWQ2siFIEWs6KVqXZwPh03f19SAzcMxsM
DY1uemJswIh94x3/dB4eMjYL1gF/rcSAsmJw96ujOrlx6mxGPdIsxQf5ONQ6
TXYq0Q2XKAFXCxh70dusiQDhLnhaKCt+boaGPJige7oHNPzpdsDu2C3RMsii
kRqNHoy4Ou1KHIuyEE5Mc3WP2J1swIFas3GQM+dSjf7e7lTaG1epEylzddAl
HwgjNp5Y3bseOtVI70ctENIZ3g4vHbNtWasTz1+5q2Cau1FfftXgnWKYsR5y
N473uO/HD9irBwtjVj5aDM5TW/GV3oZKMttUUQCtERB2mc2bH+ojEcb6gJEz
eKfABEHM5AfakwR657wyWOIfUPR2TuKdURi6Dokb6E0MrT1fARj1MBXkYAhJ
WCIz0gT6vJHKf7x52CkUUcr9UuaKahe7/2/yjXZvBc+P25qhTig/kJwkAyEY
7EF3TpEn0La2o3Imtw5uC4xUWJyPl6SPICu6e3BNV0zramNJlfdF1NjSHCf6
NszMnPwnMFnqE68jUK23tWAyzvok5QeTZgAuTFrFloR4g26+XvLkKgQWCEzT
7EhSnGs5Y+HvQfiMd7+W/dHdxBFihKZOIuefj+CG3QONmy8QdYx4y5GFlvyE
fO5Hwh9QZj63NHr5wuLtl584Rzb2oQPXa6iHuq00dDFcY2lyOBrRbvqSYSoL
UsbF+nmqb+N6//cP6/RW1Y1FNvTpf36AP7KOAM8ZcCisOBx2h0hq8FjnlFEz
TIHqo+rF+iyrgR6m0NmYH6Bg/mUatohej4mJKlRMKVAc7eTtB/FYJuihywJr
AIhLORUCyVN2F5vey6DA7Ws6IELGecpK33RgF2wNkERvHRgFQ34hi6Ku3MWz
2UD0dfSbd9RzIe1qK0SRsQYnCgeMPZ5yxGpBvI0b8A1ScpXE8lQTR5ulbLrQ
GeDQ1IE1FYAo2HaFseZ+RmyRX4sddo0j7fSjj6Jsj0UVvPXAsbPJSfiXNaYe
r+Gzvn/ykglpgJ84siYTZERIbh42j9cp1wZT2mMaN50HnzVpRG/3TvjKq2A0
xd66LXKQrfYfHVM/5/cexvSwJa8iXfZRgLuZQVbxl2ruchZ3hyxhslmNodtK
mbju0KvXheWAEjMgU2PwA0GHwDEnMA/WCaBWpJrmte/ppSnV7a6+L+zc8Ljg
RDmXqyikBf5C5teHr1uJ6PA6SPquY1RpXglrGkNRsu+d0mXgxi5HDjji3dr1
fgiFZ22G4deIJHFvMfluRzkfQr/lE8UIkLKV5KVKCHKgB2RK27TEUUFaDb54
1rlFcIyQ16p4ueYZQumD4Ug7Q+LOWLym5PhA2q0eUkZOWwqdPxbLkaqw0hQy
a0p0Mn9xoH7MLSah6K2vOQ5jQEUyVNYSC4oWR0JFnKvA7rX12ug3+qFu4UWM
9cekgqMd2lQwlnPITUznC07T/8LXbfdgxkqpD/3zMUJB8Bgw2AoE82VdgKje
Jlf8u6dJ0iW85KOn+DpGiDoDAHSQ450OB8oK9YGFJAZzNHIjiyfV54QIISlu
4KViU6nau96Pfhxbio1peH4TIaDOlv2RRxHcSoLwkwv3T7GXImfUIdJLaHhG
QIjsNFHNg8pNJvA8iBZ2PwaYBIIVnvDa+HfJx7//+Dr0xlOF2pfBLLQ5hkem
fzBBtR82frH6qBM0g6/6HCiDitOQhzQFIStxazfaPvkefJ2axEQEdlu6kJ7l
vOKxzyBADF76kaq5ucY/jRwrmi0Jpgyz2wWOrVvZyLNgdXZqWgR+KOF1SASZ
DCxU7bfx3SNk7qs06fFuQP3EMy+LTc21XFURyQYn2yNP98aEgaTl+FdlNI2L
z13KuJP3v8eVYGtcVi/snAuZMJYNn2d2sF1rsz8HMt8oWXT5/3bzDEyRdBUC
g4qXVX5nDSXEIwL6sruwhUWbvIC5meCDFU5Tm5tTORsa9dWFDIqtENmJ1AM/
j7uF+MUP7cbioequAw1MArmWpdrdBlcDtmbVBecwYlClG/hGoaZ5QcZX4nFO
JiI/3Nc3N7oTl/NEBVBxZVnFwE0gbLCrrOXsG3CZjrouD0jF7zaYUCxIj4LR
Dh2yMCpqGzhOFkijetzXhpU1KI9B7dLt2fk2AjQF2CDec/5W7pscIh/BMLvY
gqzV8upcBWOQD/bgTjZ5x2m7T535yIbSaGgJFs3AkCAGLUeNq+ESwuia+4IE
EMLhaGR3myqGk/jLenAwsbc9EM/w5ImyrJtuZP/oMXW1XcaRJWLV1+cO5ic8
K8WKXTcQTY7bsIkXv68qfcU7l+g9Saa0af/E0WATeXgGgS/T7ugskSXhlSwR
YTlfE2KGiAoIxIyDUjip/SgAYpm9AqqepHwwVn0C1Bgf+r1uDXKwU6HVm4JI
CvwddCesZP+ebWXw1YMiu2mS7kPtsdjGcWD5AcQKFE07nlKeeHcB2y6C++9x
RUTt7ipQ8KP5WFO+4joMZGfTqyKEnHCimjFspq+Od8jJisspji0aFcCbO+0n
+QPKcb3fenSaad+LXUmNSplL8jeV7wFVI/C5Gg35lSaKJEFSgmU+VanZhI8g
963iM/xG1lfH4oUFv/UVLkYipJ+XKHjyfL9L4E2SIfeBL5KAP/mwjUxiBlvD
sUdx+6TTpH1FQ7qiVkyp+C2XeUNMTCO4rjYBWipb9/DxKOZm3UAcsYaArOnH
xwJNTqQnM8pvxX7XW3DqGcCvOn1x6FIrJSkPyxxxiQI71/S7hQHROSD7ZT7v
qsrgjoSLfAm+9sfcEzQoVe+/Xk+7T0X0dZ+cTkCUscanc67i+73G5q6+NZXH
fzScZOW5jmb9amd9HzZ3ku+R3CHs03mOMnrgc3Qz8Jt5p6f1WnWX4x0X7ESv
Wen24GxN0Qs1+QkfLaPE+KGKgvYmhuXjxecLb9GVeWFiWX1w4ZbdgJP/U13z
CqWrjkCsVm0JBJaZn1oR3oSn/l2F0D/IXgplyR+Q5Mo2qgBNqqP6wV3YKHN9
5RoPbfkf5B0ueXaPIRs0ojm1EXOQyiYoyIMG8cNaEmvBizm9ZmSFy93zmKLR
ZVwPC+yTMgKvdgek+xhELdBZA/yFBEzcKkMgZ/ycZyg/MoOhMAufJpc3zdGN
WcdQmc6mQ6shpkHHhlV02twMwVnutII1aVxA45pAMq9mIJRnoJlaJB6e9NaS
rDUlRzrGIrmftPQ//4LEgkAca0q1tc5hMwSQ3OVYYFGUVP/EgTxhovsxTsn2
TEklyQpIPmLt+xFVPBcH/mdChGOKYFRLAbiWycnaP39LKGBPWxGln1REmRNB
XeCE0yZ6Y2ROawyS34pJBSuv/1WkxFJXtmqcRpyEdA2vWasufeU0/xHdTxTR
yFU7msBtr3kgk1tSCZtD2b9K8sn25nKgw5kBAPeRTTwu5xGV5KiBUBSvq/mw
Fl5AE97SEbjelzlZjtJivFHcGgp6KNdb4XvJ5MazhOBO6tskc9P0rLUCvFA9
PHr3PaE1p5CulMOT41lmktHRNSSt1EfYun02Lz8B7d046S1eCzyf4zyvnH/Z
P/WmGp63XSlujlqFAvJC1zdoFMMoDhJ274iTp7vRFx4PNh4egV9knbd0JH8z
ZzTxHjKYoBl1zTJBthagp33dfzbf6aRBF3duL/lgBGpWdeNfUIobRsXiPVr4
AW4AqPzyD1Xc9vaMTGPaUf3ogntjSKm5RM67oXBVlF5UopSX60oYIF0KIAHk
AbDbB9hk1EdCrFrGmEhD5D+NV2l3MsNAuudZfIJj9Xk1bDPZrykc6/mK+Hm4
B9vmJcz5acUbY4IQXs2rXxum3sxkbKGfT7jcEC44mc0c8kd1frpAOXEZFkoI
1t1J51BmeAjqBJnjQXzv4H0vVXgKQ+UnblpiIsAGUadiItFOQ67dZLSVUS2D
j+D40wGiKjYGvQH6DzMJqVldBeM3c9Q13AvQSFxAEB8NMG2AjtTHWV0j6LwF
IJ2u/5gsinzXbONcWmxYYqVggCM1tOZLWOZnY9XUu3Gdm1whGcwAXIIBZgr8
np5gMXsmu1wy7BwhUKXAHWrkgfel5R41dc6rJ/Yzf8PgwSaLQNpp3Wf4WMhA
HiPV7tjUxK4f/xcDDaa9ySCCSzy2ky6CRCFxaGvXT6VK+6GaszDseBAYS6fI
vLtQSS8eYTLXsaxH5ys0JeqtLsfcnxhd0ISfE9tpFdCOLxzGYsRwLMQucw0j
lwHzgp7inItyRYdqVtj7syRfc+NKAOix3MqHaz3X7hueYFcQPBn1LjWQ+EXQ
e1ykOQbypUFjogvVZZZCKttFKIwDV2AGqxMw+20QUMUbBAhcgaLCStkIb1mq
aTfqSwIxGPHzgKjB3SdWicLTsEsmTanfwZEkxkbhWNAZB7S1Q8gTc+fT0VcA
kzeBH/zCRQsaWjsv0dMqkVXqnn4lE0kopJt/LDos+IxZwxWLWFrQSlu/V3Zh
NZSdsOSnBKZBVh1u/JlXkMTXQTjy9PPsmE8ZPWvrn5yG5wuZbsRzKF+YMF5z
2EHcMB8hNDVssxARGPwWAyCocsRKdg41+z6goQq491J/tXfRRFOVM8OraajW
gCDn3MYS342WdcT46EdI4XzPfxakgepuvPjjHqRJ/2KP2qmwfjj+hgEpacQO
IW8A21MOvilbFIIPT5BQeCGe+TPKzqz4riEgUQN9381lYEQbDGQh6P2H9qpk
7uQfs+YDAPlpKAcZ8gyt6mTPjeGWoSbn/F5gvoKV0h3hslAAA/kBbn2I1cIK
pd9dRwuQQWof+M/SAotFq7Wk1XWSpDIIP5UpjTNAfu6QRZbITdmFhYMBx6XM
WdMEKVw6RSu36RcgPQl+whS4AVEcG6DYE4PlDTrKGM0byPvnUOa1Qwf398n5
DVkr7DimJpFgSK5L0EE+fkpRSMTZV4nFG9EISv3SAjreoikXIAUFW4Afsky0
Ch9HC1+nrGpLghOJLRPoiUrHjSPDVqhA2R19xMr05t+9Fa5eh1+B2wjYyvYS
1sw8to3GGhHyV7Qhl65mNWsKAU6CsGRHL941S3WPVE0nrpO6B+t0LX1m0fy+
Vev5Wv98ytUbMtKtysRgUxP5A4JKIoa+JxcYoVr5BDAfFfdG7DEyDrxBsos5
B+C12PrEyqIVm+qDFOpGiUHarCh+ZbM1oIZoqHwqZh0hbBmbQt14I3Bk474d
eJwTmr8H10B/RAG8Q98/gW5p5lF5R1MDziEz6daTm2/bGrJ3JZbh3wz+N6Jd
xmYlBp79A9QcLR9/JXVGMMzUmuO2ZPrwwahFyjAHZAt676RHOhOnd6lU1blR
zCr3pvMB1owJbnk/GM1i1eknevuuOVR+C5B+5kVc+JPMtoq2rO3gayaKxa+A
2yw02eWamt6g0iGVRq0IKY5er+uRB+S9EfhpoOqrZpcNT8/xy7Mba1mQ+OIs
DNXffc9R4b7McAl6sm9SOyJcIkF+f/td03Zq3wRzwRS7yjUHTrIvPQgHDZQg
xbzunlym3i0MGxnGPVIn4BmCSUvuU5z9HjJaYmNb4uA2BjX4CHf53vykfJII
bdNZ0+MJBHQSmfNlX5Cb77hRp568eTVJGFAmVsUuphuyRj/A2WerOrIbWUeY
jJ+QZNrnsLMbyHeF/ZlbcnnZ75wvsop+12aGYnv0jHB8R/Iq6p+3HuGzw4yi
YdzPvtbNH0J9iLukERKhbZXlx02WQwKB5u9yIZhdAs0H4wM5z7UvCJPVb+qX
FEru2L+ss5vB1sbFDu8oe7+fetCTHFGZV+s+kaEZAOCT3Jkx20Nhvo6Rhrq1
4JX+xq8QVuO6YevX2PBo3FyCdrzAE0JhnAvYzFS8TyQwL7qnCbN05CZkhyKn
KoDBnFBF5sZKpsJoyXYUPfbRhSr5VzstkwJvVyZNv/GJJFEQp2x45nC4kv2o
jHaE5sUMejU9/VhT3XZ3Zlm0R0CJvaIXzmidWB059ABI15pLGoyDS80by8yU
x4ZFZPcCZeMv004e4UVKeXMkWAMfAb5owwZye7rouFBFsE11CUR9y3UKk3rJ
aSmJxB5L3JcYvwXF7WUFu8GhB8yzPJq+9CTgvBY9Dbz0BuR1d/IbGpfBhsHo
wTtcS6oLTqraJDOrtYiMnmFFN8APbKVFAe5HE0ni8wIlU4zOTpBps9U3P0aj
+MjUrsLFRDv2gBRT6a1FdSx7Z7IxSx5jOJhMxr5EBpgepujOqcZx7Mh+6QF6
Bv05Bpq43okbKDWINlIsqMEcogOWZxN+DV0ngiAvhQhf7HGocekvqe1ifLBv
2l6WJAdtvHlJ4OqI/hLkSakJZdPhXj1JZYfeHdLFn5Pfv4wrH+z02Wy52tyE
NUu36Yw8O+exFIcV+/T0YCe6trSrr6ul3g5BpjDpwsIuNAeP3yR7eUba1GAq
kjKvBCH40RQ5Iww+KQ/NqOQarYipyk5A02MCwDSZ02XLmUC31jf3y5+EJCaZ
ttwm6pGAWLjXgC22Oqjg/KYsTMC6VP9a6UorYxyR9+Ih5x8CGjF9mb+I3ytL
V4lqp3ZuuINraOc9d9ejHv9CeaDvgqbALEAB7dvYSNa4S+2t8IRpIS6H4gS2
YfPwbywag+Ti9rYdveuRY2JYV1sdaAjntnuopmSiKmsG8zLMExh2PfkzmyEp
dlS4oBbUH2drQ8weQT7T9wmfyROD7ICAJqXTSNhq3gzrFarGnGOUe2AtCQhd
82rLI/7fViDiCjwxsnqRBDRCs7ARhdxr7dYp99JKi/L14U6J0bXUhXONwx7k
l3BjB389dfIx/laI4zi2IQ4DYCGor87+Nw8pQVK0hKk2THsBSLhWZEwhqq+L
Gar6jc7X0cu0iZP5gMBWsUjzpVzfmtc6s6GiIimEJgozRl0s9gyE3ruBVs7u
YuU6b5WCM80OZ+9/SIO+id6eRltr9DJcjtZo7AwkZap1lP9OG4l2vbJaGbOD
VT/jxl8N/sZ7pFKpDQbLNlzel4Zz1OGWlmhVKZXcjqQHhr1Q2q6qodVaxb6U
avDyi9TRicItF/84217uF6twJSqqW/wgGgsYZIpCptIs6yqE5fnQt8xiZsTJ
0uRYJZ3dgZGL270sQNQfdkCUVJeHV7xG/wn95Q1NzbH8CM2Kmw8RP+zs2s7D
RgHbxoJvxwaeoFH8nTjKXxnw3h8hXJcewxVMW6p4bv28sq9V/HDKnkERlaVd
Kxx6J6ILXMPf5rcP3klCPCvpg4etDajRW/4NY4/YryPSPHMGzXWxO93+BsWt
DDH4Z5eQfx2V3l+NAwA8+RKvR9fcQEThKQ6F6IzBi7gtjij5WFKTDOcKMPIP
UQgYwDSTPxGog7nPH0DMH4YnHvXDPzPJxair9OF9vjctWBpGSd3V/2UzBYDx
dZPgXkOHiV0HM1vcvC79hP7l+wqkgM6LlLeXNdy2lv2BSmrRsZn85yd7QoW0
ohdE8QYFopQBCiThmzR16GuHFlV2UpgRA62ZBTUluT6BuEOhqPkAG8qquXTw
2tRSE4lLb09VaUWJiLG7ugNanJFjnmb2GJQ3CPwPXbfIDBOKTZkxEuO+8Lg9
Boo29k/mUa4rmIY/iVNwKUNKgtNRUMXFJtpzSvkwR4d3Vkng8kmhO55xwPDH
bsuhlBPV9gEIlS9SfuYJhblzt8A1HTRcaHhH5eUspiOe72Ol+IOdMLzMsi4J
SafDY7YM2uVx24dpYegZz3VFkQ0mK9n+ezESG0Zo2/I8osqs4J1x72+Ovxxq
0LPBBZtThBO0TUmvMSP+c4Fk3eMsSza8f5szbZu+cb4Lir7e3NBIqTPBjN+B
RquCQLQ8mdcLCX+iF7fGnwBcomsK2L9wXpSN93vI2U4eA916b3nt+CbP8QHr
rTsY8WZNpNr5usALp261sRf0VmOsV5QzAR7q9o+Q6raVvQPV1etgEMkhWQBH
g9cDRmYZMyfsULgzrvP4u0NYOvrreOXVkJhXqjB0a9IEhV4tdkmTWpCNp4YW
GYAtJQypg5Wm5H3H5GaeuuEQnMJEoe+4phdDlBDKtjICEDrm3Og715CnL0bQ
kfa3UBhVE7CNtwehHieG5kvU34wuQeLaBeEtsBChdYN6wIQwv5vki8OVMxF4
tCuubHsNCNwDqAtbAGXbB044mzNG7n0j53tmPDMNJdfcD2dUEmlnW17vyycS
MEAEWpfR7hkKIoiR+vcNhvqOvScVe8n7Vsgl6i1+IhQgE9NrFilCV6+t5qZM
GosOikdgU3SjMo8wUpe26ubNTu34HqojzU+pXT9SUR6aQS4CYAhk1QaI5iVj
PhP46dtRqsNG5vle19hjOQfvg1qlecysqMF5l4uZQ+1Dokw453Zx+kDHttMC
E+VXcgyPRFhxnyzdhugh1S6cW9FWvf9FmdMLQ9Cm1eS48rPL+eqAuLtwmYGW
xnmxgghfFjILe13Kj1qyUVYlq37unUUUiqvEp54N0Jb5OT8fsJgV+F3ejbqy
sR7VVz3A2TAt591FqMoc7Bo1A16QDPU/6DxdCTm+oNQraPHlWVQmx+1JSbFY
W3nL7cC9sxwXTye2gBHMUiGJL/p9DlC3bXTU0BWCWij2IYlknv9XnyhrYInn
7lBYQsAvPWA+gjU9ca7znt121T3tJxxx831c0phb1a4sbgtOklzB2x/5MBYn
p/7dqnACcf0UlpRxn2rLqV2DD91dEHFG/rnTny+C+8q3Kx/L83SoPQzOQ6XP
ru3iL0IXSEWb3bsdzx2GgTxr4rXdsbknmvQmQ7VUMp/poMcS0+KXVJF+2cgA
MWFttv2266IQ2r66OZVBdnDrJTDvEb036W9m0p4Rbr0wktogGShvfuDQ+uls
pnFWqVgfY+Pl2YUk2msihFfQAmtC31uOkAjTy7JtFNlY1xNsCB5lt3tEozpy
BeQq3k7XqY95taRsKIBdSSuYO1ESEPoi2KL8rTI0P/behKgsmHfx9uIP0H83
lCXbd6arcEPXHnlvx6c+Tjb55nAi+pZW/CHDOeBcknRBxi8uBLj3+YQp4Tn2
dAEwFjxta8Kh+nLqTlbIA92UsQ6qrnF5B3tqAZs6+FWwxK/WjwEzn4wnU+Gp
sVj177FN/k5v9JVm8w5AKhRZEpAx8f0nPvzwQda3qFgeww/2RWV3qj69p188
hmzw+JM3cryrjq5u1ob5nUD1b5CMea+u+UleK9mxIwiHFxNvhwUY8QKESZPP
BAAiqIVjZL5/8ByXpDMqdZ/+pEN7VfRlDj9aZqQ8qSQmxhvwWWLRVcJCuX1r
h3l/9H9SS7YPb98Uu6YMR5hZCQpn8NTRAhW79jOcH5rHemjBWtJRfatEBgRi
g7dORrE1UEIwZY34cAB2XF/3pbiJkO4KAPQuE4aoPTGQ9T+G+NCpnT+yXlz4
LsggsTC9d9o14l+2q0vgpDdVOpkcW/gzp73YPPq+qzNz2oqZp0NyWoHZp8Pc
sI80xn3qyT7vCI8e1JBnrC00dsFrPrD3EkUftbsqzbrfxw3ulCnUm3guDBNS
MI+AcrvjH6HAdJxog9e1pbMleI4AGam6qtN3dkD+SPZFVAUxWuov+oGLPEV4
GBqFVddjjMbGmCFLGIEcdqTKFPFoaVE/OUmAA6WXkHEsJWczQhPY55LIwKzx
QtC2sW0N+00DLSKXHnbbJQ3vJ8iMGVk/L040lH6ZDsa2Y4m2Ng2thOkXxTmu
hlboyBj3PTsfz+WBf3iZlMZv0/yFauRDtwZyt9opVyst23N8drBeKBvWtk5X
O2kPYf6uzGHI2pqJP2sHGLjnxRYr0mTM7s6whjv4ppUOzKo7ys4sI402BImt
BX+SC1UKRVni4lGAR0OLJI4Ar6XxBB0KA3V1r2sJVR9f1Bybs0XFHJuET8Kl
vQI3XORw2zN8ZK6aFU0oTZ2bogjdFMGswOW1ptf1VfdU4Os7QJbv5eLQnH3d
MMDauY9sBo7BIRkMT82tP/ohWM52/yMpYKQGeXjKeT3+yjqrwuSJtz+0frtW
duzmuqfEvipZlAcVT4RmsMnfWXaa5oTILw41T43mHIypaYFHON+rWdJjWR5A
puAZOySw5x9sXL8my66AXuzOCxAC1n7YT9KW4Xv8LMLnGicLfMEUFuIWhDif
ri2LPU/isJjt2+I5+O2Yvrs7Z1E8cxpDRnM0DQSr/QmwCPQbgxelZ50thcSp
tQfY2WnO0NQtmqvEw/Y5P9AWdUd3ML71wBEjCpp80LNSpmKEFLQM6Wp3lei5
D38rluPw434BethSPgS4rxUg5L3uoPRKkfckfxmsEhL0lwwXKG2mwOdknD1/
pXBIOXOj8TzXU+D5EiezibCXMiDMY10K3U4arm82lTq730kia5P/MxcPT8zZ
Abbi/ciCUOcEgHgo0R6+cbgjSolDhoPeQjweQz0hNet2ZIH8Z6k1TbpvizwL
mUkme2qa3DfFb/sUduSio6ABam8y9BHQLj8362tKKID6h8uiYwVVo4xjCCgf
c8hcphv2WMhEpi132vhQJfXzQbedjD2TM8ADy4zxYToWlaG9iDo7kI8dg/bG
ESOuiHheLeWW+KUvZbcyE9oEs3yzLW1uF2tKvBiNMQZ4wjhyJEi5mhFmRsfu
Bs5Wl93GfSbEUozR4SNB+Y8JGPzts6zGb9R8/b6bYKL2iDdzYvQomdqyaCmr
yRhQdkgHNnuqxuZetCeh+pmAECXkM4GXVMcsmetsn7495tWs6k7nqCd/MlAd
MpANrIbSb6RdPWT420Qf7rkWad0RIKs+TvZ2opd+mPJ8jq69+JqbQTus6p8w
DUY0G3wFhw78erjPmnNCjyJGpPygiN7V/9uNGsA0DcYl31boqNfjgvsjDf8d
3Tw5jxOrEd6wgobI3hnh+CoErKeN4YKXRC++V7vwDcFYEf7lFfG+EOlFuxzE
Gxxe3YAVNZSlz57eG+L6+/+CDzweAt8iEnB49280wXOjbBMj+Ty4F0RVS6sK
qkMTT+US5NTsxueu/LWSWCNviaCAGA+1mcNrmdS/U7X5MsVvR/HlxJUErcOz
oJm3yWmznga2Q19Nroz7EzuCwoOdC0KxL2Bdkq+20XJo50F5WnT20B+7AtHJ
M4bBr8KyFl7gHie7U9TQngExGnbuMtk3tztKC9Jw5EzRz18ydkXbZYSt8Qb3
pDgvahHJAYAPqZzup/wgjdlTJYRxEJTVNcuYckXh2maaecWjHqQd/EdEWjc+
lxSgpkTMBxKV+0PluHWBf2V4q8+zAf03OdQeV2XEB6jZu/scfdCl240gv/4W
mR1FoVfZK8c9GRcqyqfGf469KT4zIVR6bw3zz7xfvHZ6BJUt7wJOOUgxqots
/rogefJGyMUoeuxRahAe4hyKcFBEovCvFyy7rX1I6umacaohnRLSLhtwKUEE
ypFnKn9HIDaIUHTzTOdxTLPO61vw0FgxRrLwwQSOzLtEjd5NVRo7NwjWXaXs
62i7T2QxYvsoz7xVXtaGS71133VXltV/cPOdaFWWQTLeGO4avMmTkffsAUDU
XWgul0v+41iyiofgS3e6jpH3u5hKOsOZbQxReVh3szSfHVgZUjOl79WPUp9R
6Uff5e+F4rpJnEqrJDjRWXAaO1kYfLMPdGbYIz0cnxFQiRDLg0wtCq0mZTM4
vS0/OpHSjqd9ulqxxI3XHXusjFFqWInEsdf7SbYqiXuPInKZ+4xBXgMB9sB2
bpndSxrNL8oA3dv8Jp/lUslOUMrgnqk/CRV1tgRDUBXIgcUzBpjeqW7kg2Gv
UHiPPI1VlV1yyg7ylPWMUndGNrlUHyWAhQr+0tKx01wsxiEtn6rp3Of2++kI
aPHpCnxE29OfJO6CNFZRV14pvEA6+O9wix9UMjvgALlSoq5tQkQ4twK2ovbL
DdKGZeOYq1ATlL63I/jjcJld1ELXaDDI2Y2lKugmDa9+u1c0iDPxz5iIGU3k
MO7d0xMfDtu0FZSckkrWYJF0XZJZ3+RDppf4K8pyRJTiW70MwztEPipLiGQA
hCHV38VUcMsFvq0487cmrM2PCXPu0UK46Iy/kF0XNPunfT0j9I5nJ65vSMW0
j13N7kVWqZjgbSkE7G5Z5HhlI7R2WT8Lf2n3VMAVxOcHauj8hKJ4HC84iX5r
cEZXM1QY75V6cGkZtChA4iMQUy+KOlXj0Ph61omq9xuPzYCivjVIoNyhQArU
BAC6w0+DT8vlupjfl8Ya2OtJmCy2HqHEKCqQqFjYY7oaLfO4kA5A+TUqIud9
935NR1byZP3+Fzy7tjX6olS8dGVup36YlGwHMfecz/gUEIV9Hgqx3bnqTkAI
1EYpejnQ4HmrxoCBIAB/wF/KAvvX6doy1zdQ4MkdMgYY4rMFkZts3fTvGGh0
Y7rJOyD/bPt7mWp7FIRevveljC+ltMnpPWE32W5ygX3Owj02qQ/GCpcQu8hG
sqHiJA9f1Gv0MuIdNkqHm3a9U1r302SidXTKg8plky4czkQIzjbUA5dY9pBq
ksxk/gN1J/eouUgFtZE2YJlyHv8A+hYJ1qLLb4VJElXVZ7O0lxrSmFvVUawC
822xRt6jEY8XWPUUGEBnpRsZAjFBh6zEYlOcW6lNyJhZy+2yw3XvuAXwLfsF
pFKvv/vqKbUhhReWX+R5XwRTMmjlr0qwj2c4xK0qDw4PuYjg+mb+w7TuuYrG
M7Z3kQ9w+yuuhEiCtxVV7dWZx5jbVsevOCd+NE151pi66TIkzaXsvR6CQfYA
VDRld7blRXntMgD7AJOEOxuNCX1Eg3SyE/O0x+kEbusd9QBZPZnjYT/BDi0a
mF5vCPiWUsyzp4SnDSGDpIsNrbAd1bAO4/unyzY7Rx6Zk3u+jE+UvD2ddgI/
fqHON1IqPxThP6iIm1QaczbibXCZFK7LRK+da2ZFVgqqRYz1IUK877BMuD+u
rOkjuK2SXy7ULQ3CFqvzB3PfAxR3l1WrdvN58OY22tzjWEu2sceN/DQmuglY
Jq1RlgDwBZTjqlOml7YCcTamR972BxtfyudbLZLnkcTyZVsnR6jYCeA5NATA
HX2AEqD3LHP6MqVvINzfoTaPJatyvGUjnjcYKi82oCJs215/lzI+oM/B+YO/
c4661/rwL7/jR5zHD9ugXljekqCnTrOJRU9pmgMOnqPxWDN/kBW00vjl/8UP
xFzIj5u8oVPydrj21uAh1ArZtDQ8vpgxAzaqYA5uEgZXu2AauyJ+qsIpjLm7
ZifWOkiH4+S38J0UL8dQYJvxmz7c3khsQqBA0l/b/gsQti/K4DsFVpyd97iG
AFH951IagES1s+bp1mfPYR6QNCF243qyrJl8j0Li8yLOKhfqpmPrCrWQEqBB
0+LXNHnJbVYFwHa1LNtZhvMh64oexQjv+Uw4zdHeY4JMkYGfLlMfTtEKixkm
rkxCHgFIvZNQUShJsLNivl/I1SlV/ujrpbThd5qUgWZQWuNQP4qLcUMRJNsq
ySZ6dT6mygakjEnTtgnaEuULFSS1o2yjT3Hpb8mGdWTaKfFa7p9Jlxx/OBUG
zQEY4kK8rqMurlbT/xGv/1ABJN/bwk7hKa0G5cwUAJimeh2l8PnB4l6UTsPw
PRi8yHvUjuzfCbjqkmfoZWGILfGujQ1elOEg0G231keLK7FqWgBVpV2VQlpC
Kx0GBCcAEXi0eu1fCmllLvzdjyQMKEeC43R9U53kbqYa3BGvXkRV7FRcUhVL
C/e/eDAg0QYfrFhg40pbiWPxbKCiL9kCe13q4aPxfcj8Xyj1mkweJQ5sPBaZ
6xo66P5b2TQbZCLk65ode+0CLY4VZwt8iIBAybJKsEvPsmfeC1GqKo1K3jY1
jYbPAVaGVY18PTDXIVlbF+stklUi+lo5KJto2lAhBBCTORBpfLtLg7fWLwqL
jTYAqgf1/+TfETEZtdaYdsmiWWrXKDL83nWSxIWNIQxcdQv5FDgBSs9axBM+
+b95lPfZ16a2Mxzm872ySj03RLYYhblo9vfhmBg7j+A2lKKWqpXu/4wuMFIG
OlQGEax77gVf5YkI/48nLEgV9r1GuLljeL5F4tzhuwAULw41+KYfiASjzQVG
3fmxqN3qI2/JRDyf1raE49qc2SuOiU4v8rkRLsTXUZDIY9g9REienMUJoEML
Bh/9dhyoQm2HqPhpnrLxBVja44pjQqAVPl3iPFwzYggkxlVWy2iNqvaMYsCT
UnUf3MnMzDATNyoQ+ic2hy59kjRqLncN9GVaCxJX4ZzvupS7weB7fnxRvD2e
8jsToIMIgIgQ3AkvLkHCw2ay2nroKgWY81D5b6c8d0g1c2gUpr4+286fVlOM
qC6bD2eSz0dg8Z7GU2P33HcotvisNxP7CYwr+nBLMY2Yo61zoBqOCYv4Vgse
WLKqbY3MBZXVPtLcF31CpqcsyrRPzWKq99h0A/RAdujEaAK6lkwj9MLvgQlD
Km/C4CaCCquSu2SlKZQgzSr0HXnTDGh59S4VrNj4KvhnA7adE+ib5ppsaW/+
vX4Cqtyoe+TRLxsoTXb9gmR0VWeECqfgPHAb4DIlYxGwHuykBMQI29L8Vu7t
2xYNBEbR6ty1/IYF0xtQ6vePtZ1bnZouiHvztKWKFMANmHbiAucUJebY/u5I
ebGQJdc6kA1MSFqmahZBVGBo4vyR9VVqZgJUvX0Op/IDUt2SpOks9OMTYrtr
AliXFXMrEqKIimuhXwxstR7f6TzjwQp5W+lviPAiOIKfPkUZWkFEHtdwEuo1
bTmHwRqaxEJkQL1F5h84/2lEvEFa8T8yqbLtSFFRn42vmwLkoRzzRVZJAHNY
26JdrOb9np1g52/Xg/3b8S6+BLxUSnw9mA0maRki2kzocDQ0+TamWKWUk6Ao
5qLBS15iVrnnxXmhPEGPMuO1wpLzG6O9OutKDY6eb86E7hhcyiCRml6aYTcT
q7bkp8pnAf0OTq39aOka/S7evEPfB6tZGvt4n+PrpyqYVBJcxP7dmBMezftJ
d+V/rWobsiDIIZQ0bC2wkqe/kDHo50ITbpWqzH4Srxwtl74ELwFMfFD8JMXo
yI48tCh8xIlVOGd6ZcZY/DVCpPabUzBOeu3E7a6TOvLKFXcJNr3eZum3UtHl
BuHPjmz5t0QRMgWs5t+OYnrWya3voyFwF0Og0NjwAvydLOWRtS/xJ8J0GwIT
8bxmMTxPPHsltgelq02l5DAmuAXZJPEgUzBRGjvpn9lUyKN5Nsf9P4Sc/SaH
frWYopq6RsMgHrMxhTWo3tXtwEHV68En0LsBnrWUs1H3G0E5F7n9vEXNXkza
suvFnYEgu9z5oBE7v/YXM1fuoTcjQacFEQHn0dKyiS9UEfQImbe1dBmWWo2V
mXocZ3Vl1T9YOM8fTaessBfmnLyFyK9XrPhovpXIGdmGk3FkqZqz4wnwnv6p
RcDyBh/+3EHADrTS0Q8erWIJNVO32aaHqQ03MDAd36abFbwhE0+x6Zd4vm+a
7HQz9mZ1kPOuNYM1HKo7mlkckC0RYB2yZjrsR+XAJkJ2Nc+LXopM10PcNkdN
MUqwh2U99FuJQKChURbNxaAlPeFdo/2pb9klLGyyb5G7B9sUXfNga1YRQmE1
FFNX+y7k7p6m+ppjiFZnEAYualrkZXsNbIe/K5Ei3/ZkHwD6kRd2fykmMHJh
J+RNxUkVDsnu0JoAN9wZwoUqqXQ7TFUhHWQ2+YgpJ9E4BmYMrgfQySK7WjnU
OfamoMPLrcQfCObeTYzLZ38VCnwjiEafXYYMCY/lQmWaCB+KkRa5DM8ZlpYe
4oSBcaHtSTchGhz9l00N8BqsWKEL5LcAG4Pp69D4nApfX61wWMQL3VT9HH74
eJw7FHNVriLmtaIuw/QkUnD4W9KvFDef/xsuYKsBGHjEyCKQi16bf3Lk6aYx
6J3fWaZ0or9cGAAZ4LgZEdTbyFwLUPl1cb08uemEQzzCHKZ589az2DIljHd4
OVTehr7Cr/wvnUkAyUk35X3Y9+1z4kI3+tr2B1mfJTg7oyJ/ES6DWmfQV3Up
ca/zeRxzHKHJCLNesNCvQI+4os8Ijk3N/PMUR9uGRYUZ7rv/IYNNK7Keo8DU
bXBZas9DVH1kDxyBw5np6RhEuHLKIdGYuQn7d6QHpchiJ60WIDc/EFgIIz1g
6YvbIFpeA6pLn/n+HEphD1JCk5YIggeRQSOdWGtoycDvsNI6DMOSVyPwiXZt
NB6BQ9pygdoxPw/ZpsrSq5VL5hOJBuxn1u/HwoJd9vxuO8bMQMNTfGZy3t6B
Iyw0TwHWeo94ztEGRIxjrATg4ewYIKpI58hUC4zXacfjw0396RsVMmGQ6+sx
UFzqCWM6OiqsHzG4vZxz4IcENLOAy0D48wFTjQ84HYexgQ1mj4zcolwP7T6o
YqlaSA1ohF3cwXCt/aPtBdmCkuNCnnuqn2ujvGseAL2q814UrFHtoZeylHJ/
BHBDbfyS41eued03jWLnfRsReDqWTuR5IkndhBkFuRtMwd85vRIF1K5i/P8u
ds1PVH6i4fjfO7VZ+yxKL1jCllLhrZm5kwdRNM0RXCSA/GQA4OwdoKrSUM4H
PkA9fmyWRc5Wc97DP1mBiPSFrLkxVNP6NM5XC5WV1vKgE1glxNV1FDUynoBr
GL8ul4UFJZROdRrcxc8pxZmVlqjO8or7XewYdzFyFgTpdx2DIHTPhtcK7Fr9
8lf/ZVTeUnngLjeqpbVckwzeBcla6hIIPlEcV6060FV2evSNn/1ew3ntAE4E
sNJK8o6LeeYdI7F3KfeJ5Y0ipsok7G355uWrhtpjbns4taLlYCmC+rC7Yu1I
adFZeilg1g8DHQ2D1kn84BM+33nHwxuc7y0bzTF0+k51ok0Rs6z4OxExUvtg
nA27o8xcENz5EhMj35DfYppapw4lGyyof+G1w9HwnW8XvECNPYLCGoSeW1YK
nj8H7jiMIloPQ0CEPLeKKF85vAqqDp4xjJ5ImhPCWoPsZz3aRsYAR3aW2Tr7
Fu2d7XVdGJiiZ1jvkMziDtEDV5fQrMZJOYRdRMFUIPw+qtwhZDw7HRAuOtsV
qQEiHr7aevwk7wYj2G4JdZjNM9vbg3nk+xGiYan5WDEX2xt1RgFtDLVmuEKR
fvS9nSQ6yJVOa+z+2OQ4VYwRrRNRygUqACYs1KI2UY7T0CaEQKjLaEkTrZeN
JeENDkUHYVgJn7pP3vhov9xUe/CGCo3DMmh8+NcwnaAnH+lmZQJ2Gh9F885q
kmHxXizFrQfDDm80/MJw8qWtBXulfMuHNCMs29Lg5IBYzOissNFoW6gv5PzI
v7ucBPOgBl8+C3CcTxXECFvPsjPbjwGAMBsiJAKRB/gGmRchd9NbDjwxH7fQ
Fjyg+IZWZWlG9O694Z6FaiJhRetrQTYsk+ZKPsyu2zmsX2WGMuE08xwuN8Lf
6k0+4jkFIJKPh1Ryy1xT3kd2dZOcGNB3jtWPoQBNV4lkJIZSJ6+As19RFKcJ
2mI6QqaU6qpELTQMRKmwdYmqZOSxjS7kHeL8LzlxlypTNcaBeMSYwW5+hO1I
+a3/uOaMh0rEmUOqRicVN0ZxmCmDsegco+PaW3g4rY9Mp0blV40G0bhGWrQX
TLjXh71g4DFFmKP19C0HK4/MdkfkKW5YeIt037/nlPlzU7vLvl/Wms2QtFQR
zMH3RGBvQPJ91BdhmHolwTRCNfO0W8Nu1BcZ6ukepPRiJu0R6I5hFtibarmX
tSZ0dFj/Z2P6iyxut+QiY3/LfhpAgFJ+ucG9vc/EyUBahFoCaQIobeZS/oof
+lPbc0OrW0sbCSpNbrSMcw59C4Gd5+5/mtifPjtcT3hMCZifTOqiC8WPhy2x
mSVooKdg0jLYfdevQ2W0oXXRMGM4QdOeCvvIsFVNkamEdmINBjiykdwTtNdN
+un+HbZdOorO3dhLgtRmDiqLe0g4cNq9+veFXtBfImdHcji7iDOBQeiHbXXp
gx4KEhClpVGDOJhacSlmOZlLHY290wJBCNddLCCV8kO2JK3N6MzSH72JNyaC
PgOIrg6QLXMmhpnWH89VLjUihO256aVIYfMIfWnImC+g+QTR0ACnzywnvKtK
zA2Fq56thuJhiDI4JD1Y5sxjuS+cr+KGzwNh9HHl1ULyXY6sArIGs+q6gvoB
lE/DVsPPl+ZLDr27CHgft5eUP0tUhLk3hYiq/vr3kLppPobRmi8NQNpTVW1c
VI7NXhoan6WM56MBi5mhu4arm3yZIn5hgurBjz53qZBl5CxryFXFTFNLaZVp
K4NdH0yLQjZP5TxSZsh0l9AwlgUGRz6Ye/FNhBMu1fUT0Qw8O3ouxXYmIy6u
kqUd0+jbW0EMm+2oSvOB+azGq7928K1tRyGegRHvi4rd/rc+B9nwYxr7sI98
T08opABsGuZuu+/DC4wsIv/KW7Saio6KbSa46QGY7POO+LiQmqrRnKLLF9f7
iOM2D/ac+HQqXVGvE4QIGnBsXe024xLLssDVE+wRrDEKUlemut04cFcoSk9r
8QTUpr/WSGHfFqjKvj4YR3LJTPRe+vXO5WeC0QhEObPLUCQiJQccf1lcUkGY
5XomCXvUInh1fTvGWF87W3gN9IUY2uTN/9yAhn2WFJgcUtDqVXuoqC8bYNMN
LtnlsvSMqNv5OKp3ECaNDodRzNKSDn/5FC0K8IyZfLE053DwP/VBaiaIimEd
4NzOMdDGm48f5RQID14OxoQsqcz7KWv0tkAQnS6Ew2Wyi74G+s2oNXD4y8Th
FhbsJjOZfQlMZfCXCT7syI1ZToN5VXzfPpXlV3hi2F7LH0xhHJx+jSZKTci/
NUeH0++NnYtfGfcTsg42WFP3x/3Rx6DOs7ypWkffz7Xe3cCe9D0RRrx7toih
msRapAR/j/QNntBjQzIyB2J/toTFWiB0K2cXk3ZN2kLCXMsg86Bxhq/8CfXQ
iVbSqsIAMNbcitzZSc46qp4g6/ouXIEigvAjWSSKFI10DpIOCaXelmeRmpad
7uhK/30pvZIl6xwKT5C+/TRjAD22d7qhwCGUuRtgWHVdYLYsngN1awJWySYN
8u8mQYjvHAg8ANVTxLViFi619mcQIbkklwZRnHpXZh/fUT8BVniv/mfYeJc/
rNw1/EHO9v207+rjdzwmn73LF262lGJNYIVJEoCfjYbLN/fZXqw4RxNPROeh
bmknvJyaFeYmUtIJfXdG76C+kmQxM75dFeMMytKRyg8MTZWQsWF9XdUApDIh
Iwr0UAuH4wLLrFkUyzjJwx3udNrQmguUU7O41gSf52kdUEag/2ZC/uQ5FK3+
raRTTTDJs7iEKpwswUYd4+HUH84CntiHKYf84VWxHeyRB4DwWFcASYMv1Fmm
mOOBKRiFRcdUpHxL4KMOTJ92lOiGfYGEQJUnAx4Xu+N3JwEMNHEYsZeV6eN1
la8lPj1K5Opq3grcd8Lxt2/jWQ7UAw0tydTwVv5/rpVTlGkb35B/wnJk+4KE
RdDOONmzFW9m1IKK46Yxk9zimUuXdi2/EGy9uZqkSTRtZw5MuvcxpntQSd3v
pcR1fMxeIC48EP/6OOYEJrUFfPVujwWdu1l/TfHy3ZqXfOV7/sZlvSGuJsaV
5XpFuqv/iug1/uPFGvfmaZzxnV8f8o5lZClBPNxbWsSaFRnuTHy0zqJ9J+Fg
MRQ6IGWvHKYboSvOyz+/ej+CKWAFzd5JrHarOsWUBMQwpIa3k6yGDM9kpXMy
+9uzTWSLvB4jY7vDn2d2slojKyOsG0Y0rsewzqZcWOXAW75UQs+pFtZSvx7n
ZF6x7VhtEVBH6mSkql+E52aJQjHXnVoMQicqW2m2qAu2eOoOU+qxwW9SqgC+
4o2u1ziqt6l44VpWPhzJMpx2i566GbN3U1IelsI5qIqgZ/plmX7Pmb/nHGsh
G3m2bgs/wVD7cl1mE1wfvR/NnahUBvkkBRL6JJiscreIed25n2ZYaaGZf/yr
BYbDNy0yp7N+iqg8jsg11qb4lZC5l2zaAssW/eUp35AKUqn7uov38BBkRCeu
OCDtAS8KDWa7ojV+CAJ5hJsgSSG1bltglYc1NCmb1S2T9hqhSWCvR4v+6cc0
RdnpXzrR85O21UtrBTA4zVYYd+1t9BjB6A76eRksVNvU5kof/8Cyx5r1lcJu
t5BaMg264RGqkJ1K+2UFFCOJ9bAuH/p0i6fEUDxLphNOUdZkufaL7hpQZz6/
SzOoJ8ozUjCV44SG0dM7zUIjrUU2097yWZ5XOgRh4lRJbJhbBPM5LFDU7N+/
0hi/iZubu2W/YgsgHJRK/6cK2PVwQGOqlcSC/CpoiqoUZzGjoSr+u47FqcxI
7JilUKwHaxq/LF3kU0XepQ3BZD5A23+fabUcAq3OjxRgqfDpWS72ssNniHbe
YihnrPkJkQkMxmBmEECMRk/2Qq7TzPDppewBNIvsNqwPdHbXUsBEhY6JdFEm
CZJYTsf84ooOx0vlCykAvmSzwihvja72NmM/VQwvB57JQzC7rMTYSlVLnbkL
TYYJs3EQff2fjEFUSk0x+hZdFxuyFwFxmaRpCIX7QOV54MnREc4iqa8nxDTQ
XfyLIx04CAgF3hUMUX2ArfVsVWWQhQadVxdPyI6nBc3Ny+o2H+esMnJm0BRB
DkAdUoo9PkKCkwBTeBdLi1aJjjo2qLdf6HiOWciKjCBWWrXfkFGq1sj7aeVl
Ymn+7u9j9Bs7WVr7+fmCQWGQ06p+9YjGRP/e5xfbYTVs+cgo0S11iG9xIK4r
BLiihQn97eiPHP3hNIsPmEX+v8cIJw9Lb//+qC8Um3DlYY/j/7xG6XvCmw7v
heeQ/UO0wdFEfY8FoQSQhszo8DVbDumm2VLnXRKU7JlRLZmfjvLO9RFB7RMC
pB0j3ND4FFpu4mjIcO8bAIZipD/OKRD/3rFONqyrC/FU5Hm2T+4oKAaaSyXa
7DY+gb/nsEdZ/KFtpNKI41Jua6z9UxTJqor9ZuNEhwGkiukrtlaBv8i43lRo
iRsqsArTzf4Nppkxno2A9uPJt5QPQDbxL85jhOoblmXPq37o5UZxtHqj65QS
SQSTFGsQMYyKVpuae61Rfr2JiJ6+Zv8es1cE3QbERj1FQdlJyZALVvNGVlxw
mPwRSBQ6KLvrdvE2lAu5tyK9650F0UvVVHfQmODjYxcXO8zhFjniK+3xA7PX
rv0uCQ1HY2RsPauVKwYW+MZIaoRn1ixrwJ9Fma7LM8gKivA/mWIoF6yoATgA
Ma6ReAl1g+3OXr/lYXRc7OvI2uYdqgJhxEqcsGmI/1hT6tdJtNeh6jBeVsKI
1ziYhi37mKz9vYLEcWtaHAddHiQyGZhnoxhK4hOjzTpewd5z46btJ9wUkgXo
BloOsBULgrYAhIThR+7Qjwczwm9lPX4mpak8C5obdYsKzv5YtoDr7OlF43FC
V2HIaq9+6lGfxQDfW4dbpjS44dZnPACm1E/2WbiQ6nUrGm9p0urfb7gnKOSS
swUysU8grQlS8ytQBJinfzniTdhAa4j7+A03bpU7MhM7Z4HKqDQDajl98Wny
FzuDCwpPk60E8RIaPT5wmIx8PlJ8LB5zgwUjHUOFK3TuW5QpozBpylpNZ9c9
KBvYUgY8W95dSichLf3uQLTH6rsPQTTINNmi17X443TA7XURrlh437dmo0tn
gxhqPHIqa5Ptv9k9WqueRKtI6EougztuH6C97Qtz4CPFNCrAzdpYX7PV5nyv
BdA6dTzmesidEmZH2aqnyTav8D7ryt2R4mdJk2AJMTAyA746ASlellghmb0L
x7litTBouVwKTSm7+xftsFW0mHf4zubhV+9bgkpO2gAoT72xU90e3t3IFR6u
OF3sOStV4R0sf3yPrnYU8Cpo69eCuJRDZQHGSrsPfghDkpqDO7p0JNuZTVFO
Sm/J8EQYWzfbrPGSzkZKKdnyNbGMyy64pHRTvQVXHYCe6fZt34ZSIg2LIbAD
twffGTzgp+nleP1IL+Ot90YkA/QHRKfWA9QlIqNbkv9S1/bJ3aelFqzxIAyu
XbR9PAAEnVjJuFv/sELBLctbERL33rak+In6M5ZRuNs4ewxoDkg18wRqgNsc
YcjN4m+z2CzDlfJ0f4d4zM7/xHB6fUYYUlpQRd5t6PTwEcXHDrYUY4X3tmW0
pnPnECuwK5DP03JRt1NM5i1QFUwfGa4bkqVZe2Gg9wjMuS5Oa53Yud8q1x1Y
6UWOEgd4yKedw5o4I8XLS1KI9s6L2rJFqca5XJKB6TqIDtjH4fgXM4uO0OdL
94sFMi4/UFzxcz6Gzn0qEU6EENoSmygAWvg1C/jbReOHVC46k5FiorizMq1B
jnBAOhWD+I+/nftNI5uV/WQ5whWrt1vpNSUvPB1Af9m40eNxCNAe6aeMKKSa
n4V5WgcWyYhN0Ueqj6+ULWGPbZUSNgEvxvN0S0KZGz0dym+wV4vDRtI6BLBA
bXIYLKVImCntucFCDuJGxVTS5f6U3gemLyaMR5B7oHYTNgYRFBw0pNRLoWUb
l9Qm4kzq3wd1mF3PUV9LMTXqgqHnlz8stOYOH6nhvScSX9VXwwf60cpaYH1C
8pm9ol+BSWGTuR5oBKqEcUkFoyB4G7VKhctxHtnAedrdR4cjST6pFyzvcwFa
0ZDLecqy8t2CWu4FW0LxKCrlll+MW93uBhM4G58i8XePlR4aT91s7x7tGwCu
+3Rtl2robjH+Pl7WJCq5DWAfP/xG4Lj1Dnfj2wSXwMRLi+po11N9RDaIDQYB
IBmMq7upc6OrOz5wzpHQTEj0Lr7ECO4ZAHOocSZCGrHSPIiyjQdh+H4zBmI1
vigashvXRRgYV/8YquM/Vc5cy5A2fu2XuUdPRXAXg/bAEBwev2KWU9KLkjOf
S9w6bMr/UmPuEH5MBf+It3XEDVjf98VJAvZJHos+eazNW7m7JVMXTD5/Y2n+
wW/rtAVOYF5yKjJovrKTnXYP1Ndr6qBWQEhC/pj6LuKNaF+BBDwL09eruyTz
8u57ttvDRrWKWqbPaO7DW6U23VQu8jCtW4YY2n0Pa+2C0ZKRtlowqzTUuiKT
BFAt11TRRZyM4abVazWoWcY15w8CLWKY+3/Mbj1AAZlEmNqLh96Wo11l96NM
0tQcBg7WhgSG1xLWafjHblASjSzKsNKcW7e8ea4COQ+n4g8twlplIAihDaaN
EYniOuI54knDErfd8H/LEU7e4TyR91L/2mX/PQ5lv0JvkUp9QarS/v+V61NY
/hMGb6IpZiw0Hdc2H8SaloGYkpbr/RXBAfArU8WjeJQv05mLd5m9/8ONNJeW
gc+vv3bWVQCbIRiPWjlfZvPnVSdo5Q5P4AYHFPww0QZjVdYrF6IfNFzHOBak
fZ6JR/g41jmcVelpd1PuYHvTHjVlFwUE6gkCFTYT5r35rzps1T66lyNndiNc
EOGmXBCvgYHDDNSGn6Yaj++sPcksUOqD8cPplSGH3xStcDf7SUYNjS68EIo6
PHlF80lY4XupcRlPxkcrqOw4Kkrn4hJ15Dr3QUB9L6RLdRK4JHYSi44gmQ/e
pcHuWedDS8FpqJS+26rRPQMmZNX5WQ4T5wXB+nvs59MeJH4ziRnEb2UXPBfv
9IVl1NX+1wSwCAD2x+929VaVP5c14qp2HLegIxyMPEcIlZYs8Tm0TqWnPufK
IeMxzopoVgCGtJD9yjxBES23xLVf2xhZxvJG0hv+exCa1ew500ns6x41oOB0
5B1uAfCA0C9gtXB7mFaFE00imTnWSqlWckx5UOQTwJlfwkRD5EsphLV0dsIv
XVeegDRlAtFvygPwqlPyE+zkPYzsUT0SUa3npBcD4s0Chr94YBdV+nS4ckF+
Dbgd6+GxC+dFRzBKAvxYW1YIFBHcUR9jg0K52dFy4qGrPvanJ/UonGS+rcBO
t0VXiv7Z8Vy9I3JC7e6xt9uOMlQF1tgRmA7JkvAkgxVMOe9+iP4gohYLtmn4
0gywzd6VrQBq3/RrmpYjdgackCnWkR4khPZxWxTFvZ+8dq2UaKAeYME4Gu/T
Mxu+jtruUs/TnvZlzq9mQfcViW9y/ZBwIEeET/QPcjzIZLp/rVhdyU3qPeAF
f0OQiCHYT0RVV1zIDhRWOsF+VOFbUS0ry5OP1KN07c48GzbUl+lwdY7c1NU9
KY9RTTFCtnamzDTu9BPqkUvwzZaFyMCHlkl1pqPm45IVHlcnTuLp3mjYJK18
TMdcYrJTgqKOfxdf7TWn6L12sQwa3aIhnYJjnESKZAYl4fVmHYYK/KvrH8sm
2EdoFoWdS9i73lSTcgHHX3hWNt2jEdi44v+aq6jI03dMhFCMi1d01nzVNiV/
Blad/DcUTqVmVRRpwZTx/0hB++IRYXdPFbfiR1OiXA9jcJ0tshbEdC4cEoJE
ze4ujEviOAg09dAv8xcFAtBqGkDdXbIOxTUGzELkA43Eng8ln8msFSC/OKm5
dKijz7BGfjrV1di6IZit9L/j0rOiQ64RXHTs/MVnfVl9w50luGqQoI9VBnc2
HFqjNUKOYzwnahQJRtoASzU02cqA92luukaRZO85/QjIfsQg927bLZbCLV11
zDaTFjZIaY7RjfTH68eogyMlDr+Xz5UutaJZkDVCJZopEW/y5Pg+rFcIh7w8
dmjgXafAwqqPI5obnuFRt/w/4rzH9I6IXjCceu1hUXusq/NrlbKjbdF5AB/G
8S4opde3oK1+KL9sM1gy4fnkRKSClBPab/HVtCLxAQoWIkeu1whsw/KgFcNd
Uhji6LaZt9KSEVagvkd0ILxRy/poG4FiaKqmsSoefyrV15fbIXsuWrBAwvzm
/oAcqd6AJv8aybHugfCuQU5tCJGBZbWIDjQRagi0/foAHuX+ClpwJturPh9f
iy1V2QwS3u9Ik4O5HH2wzgOmcijNAfErshZJd4oJ61m2a7DHTz83xXaI/7Cc
F8rTLMhD3w4fw3hQMuKbr1IUf3ig0u9zfblB5boXAfJNGZyhnrH3TAWs7oxj
nSnyo4CEUeGsT4JY5D2jkTJlSKhbuNO/iyGbUM1TQvxj/yBeUecl7CVU5EXp
e9oUbxDsTexUTrXSszZJETwfqcv9lOLqKOLQJdfgvH+f3X9lkSJPA4bHmgME
fantkfI2If94RVh+iRbrzgQf4eBablDqJuEEU/IllhcE0gWszBRby26Juk9O
zppOB92ZBV6vAD6ONfZCXb07QIeDwWpZT0O5Lri9gQ3+ZZc7GHPUDEJNVNIM
4lboA3iqOSZpEEYIqCpaM+KZP/MUoA9O6lwTYorWxI8PnzzbF39ZhU5sv/t1
/yDXqATzXK7HA5w8BDW5QqkGMXsdUVZ1Een4LHoh65EqGhdm+Sn2FiFLr2/X
BOpz/McISM2R0zYWUR4nlQlU1u73aX2Fdl8f8MWFgsserTAoVAF2JuG2QM9s
CnyX5gRSHuIPPqhDMto1vjSvQJDhZ3JDUSJkRQzetgwoJaVbnqrYqITcyOD0
1Mwc6eOH7jg4id7/yhopBL+7QGrTXP3JT6GqCtbgYBRef/EgdyWQc+Zpt9XE
5hhjWkU9VuhE1Rt1uEMaF3Z4aZqYTqSWm4qlTc1ZnCogbRM+2/D/rkOqFm1g
5TWzHnNUcosS3DdYt+7p+GwsJzmkBEhfn5ipcI2sMkAGqrvuIrSIwvIIs6gJ
lMyvItnPHmZ+HmxL2wDFdHnxyO5om0DxPWa3nNKSZO5dQEvd61+/SgUnTtXp
MttC1eDXz5paaaI/2YxOjFYwVlAmdXODYHxVnE6WL9eI9BqucT/HC9QiZldq
JAB4FY3MrZ0sKunqzu3AfkZdAC1c0gN7YbHzsT346ZGPL/PRkAFcbeweG9oN
hPRMYU5k+wEDK67PVS7waM9gOasZISSNvxUOUplO6PfxDm4DJIXd687gqITD
L9kGsBsGVVymV+oLwGIAhNjYIl/hbPZ4IThFvSJhswj+5XKsyvXim9ccyr07
PINW5NEyAJZBK0uBDYwmZ4QTls9YhlPwcbShsSdoBpTkjvyDVA2/F7DIRZIe
d/mGMVm0+Szf3lw7FtgbUb0Wneo67DHsxc/SLRP8u/i4PLt6OrKIR5hFI156
v9LFo3tRfjGca08fHpCTgJ1pk/r60d9Ewp3Q+Gz45eKIFQHp0VzKhy+sUmXQ
4t9wgMeM6lbqrGLOD5ofSVJ4Q1jliw/r0claVEX3wOdZmICAA5lpNZy8hmVa
EBuWfeP3qmdgB7kdN5BOhbo8LCqODnir7RkqLsdoD6QFkHHXjx9GnN9Pbv/K
VYmOn9S7ofqw9/mxmXxD6zMuAbT3bwQPiS0H2lMJYdyvyLRBjA9m5E5BiiKV
kcxbUpMto3hUyKnqF766FzjX3OEJbKMmjVIIrKHO51t8ZopJGw47mwDiWoFR
gUwsgJMp7NagvyejhAipVdJQYsSo6GpYjMcXQw2Harp3bIiIW4IPe19YRMMk
ZViStzSNOFq1jyfp2c3m6Zt3r2rCtsqeMVbLPDrHWqqQdfvBduMqcI0PUAK5
MjrvaOUdTpDPzy166eBdoiR0iKZ5MEzjlFM50LZRny9sCy4iAOLELdfAMd+8
9sUmW0DjFI91VYOYeoJM1PtSEAuMHpGQi0tFnFpyBlx/QHV85XsBTw4gzeQj
Rh/U09vSL6skLtJhhbt/G73iTC5SxpiRaH/gT4aVNRzuEOEoBwtryq+D758o
oLOm4IXf50g5qWqfySidxxw/AffuzqYmgTY002HfMwsFEm3AGZfaqekfxpq6
PhmKiWkZAj1ZTKiu2/uZwvjFCKdQkK4fTrt2VVrBFUa10dBpnBIMgihQIxCf
q48UQQ0u+N65uep5xOu/emsZf7trrdSCgZcUx00rDwusyXTOKSBX9yF/vaie
biUGRzSeIZY+rXmKx4fDDiRET53MU5Ku+VZPY3+IjGcVrB5jqO9p1u0hF4bK
1Yoz/hAAN4w6NZ41ITXJyCIwzv/Adnv9h7Bb4lXzeoyNLE2yYgdmLwBQOeKr
urtoYLutjdX86AZWJfqLFpAtPKH/bIQ3rwOUHZwquPRM8xHVEnJool4i48Ld
i+P6nPfuQaSosr0H6kAVDKq7X2QyYF4NodB81E1QFU4QubG5yt1a35tIIHen
3IXZB3mQpYu2+W1x8JRp0qcIEcUvtuVQvJii83OabdH8OFNOJOA5XTny2yPS
gou9OFNMd8jFOMi7gJHA+yNy5zMNlXNn5cuTJgh/SGhpf5YqqBIsU1BW7LT5
DPhBxasA1MJwy+PEV20XiQWuFotfDI7fJOwByUO79xoY1GCtCSI/3OUBzp3k
nSDWKZlotlNdS8G62N1jc7BPe0v2gocIlXzQuVWTRIUOMJsUKjY0grnZybnD
Sm0ifTERo9JHQZd9vDaDfqEYY8/Jy0/3bAmq4QxzYc85QUikiIpf3mt+csp2
MDZlGyO6JH2kbuXNGEn9cqZoN9ZduUVlfk8/WUHFkIeSJzrd7vJhXNB1PnbY
SUCbnUIc3MQqY0MO3fbeZFj/6jqc+b6tg3CnoPioXmWfgLxMF8xyyV4xyZEx
Dete+BeMqV1my438o28kth5kMDYEWSnQuIU2TWtP7Pa3Q4u3PNweN09KG9Ws
Wn+dWDWOz8I063072tjqx27YUkkKGGYBtkSUSguWIwZim8xrPMEWJfiAY3Bx
lXJ5tLE31qO2uF4El1CIIwwVHUzcYO7Cz4INJFJOcpmrS1kvgoi7dylHKT3l
fW9dXsdstW13gV7J95D5gxGiNgqFOJHaqhaWWbPuOV72FnDCSZN2dd89HyfM
NOkjh0cbM7TM9efwoJJ8nAgZmXALACf2FwUK50TwRo3c4GGtuq4rzdEXdTYP
RbGX9vsIiGaGtl+dHYLa0mnxKOEBD6/w/flTcV1daOyzJd4EnPqxtwu7k+rP
1IjtI2ySWlOYNjSMiqhAVnr9SOf9tIhijMSMkXGqhUq2QiYw1G/HhCzBkVZJ
Uwjp1K3ix2pBJTaFUqQyahxQtP42GFHwe9bPuADprgqPNg+XqwI4E/GOMLGr
rq2wUlKgS1YS1TzjhD8UO5TrbbdsEcmTNaFlI8qoJD9lXzR72LioPyZozrax
4qRFZFAQqodv5qNrbdd6KTkI+iz7mxtzT35KRL3hMkYldk12gKa5UEFvd6bw
wEyv4W/YwtUXLnW1Uec5NtSdOHAbez1t+bcM4F3QWL9IzmvZR7r9lmzagVTD
fw1neSEe4WbElo878GuVAftTcFuzL9F4XTQjozHVDpogvBeuFiNQHHeY49mx
g1xJLimyeGpWTW+zfTtI71zvWaWuyJsB1eO2vckdvn9+o4jMEwUPKIUDjjZ/
fAMeMJqbnu8igQniw32PMW+VoHbOwpEdPcUWFER6/4JE0AAXK5HhYr1IZB+S
o7Xd4AqgSQtjTfBJQ35z0rmknBVqXI+y4rFQKTUiO9vCBpj60RAEt5qwqlgD
BErf5YzUIRcMEh3GrlAbkI3ZPVunA95bZD5MQE7rIwHmZuOIbGWlo952mMnN
9Z1mOTdp4R+3oM7yp/aJeRc4Kk8JMXqm74y9r06Gm78P6z6BUapaXvsQUugR
qY/yU+Ka/MnBMK8c5x1OnoCWtIwLAIV9BqlNfVo/Y6/zTjestsa0n1MFkkkf
Pg6Mk25NbeghqOiVR1x68/ISeP5mes79DCCYovZuSmfECFsLdiXk/FXrbZ4G
obpccxSu+edhcr1pwwowGf5ChrjyGXQy6iErpVNIJVWs6JQbllJgNaVmH0Bu
KAjPJNY1XUzTgdSj9uWQpuquvOoNbUHroHvonAuin23O1SliS+ImUh8PZ7Gj
EpnpjgXUBAZAaHg6+WsAlFMrh2KW0BCtOzBZcb1Xq2C7miyWj3hdijNhw3yA
TC38/mDr0Q8PwX4Di1qmolJpdYzVZrkBDiAnq5rlwD94Zm5pu2C+97VEU0nC
1gfzke3jk2XDoz1wSoV+2dKGW3ScbkEjQNjOZ6seAgv1RKoZ+CeBzz3aQatQ
ykRADCc0c/hk47IBKAIxahEj1EcMEqIcVXzRgalC+fm9+X39UqKAOixpkvV1
t7sFE+NQLab8QKgKy/jYzId7DZjUMaloQ/kBlVTyW9YhLEsS5zVFufxNpW5m
G4NRn++U5anuIBhdDJAkjcP0AKIPy3le1Pd46WxdrADjmc0m/VpYVz5uefVJ
6kwWorb0d5vGH3AmBioTlATvTXz881VDLQ/jIESCgM563jux+9EpCtegndhw
ycTM893bk1JFc5nSAPYiyZz88hWlLVFXpjcDI5aKX8NWn9MjiOQErqFl1jec
wQB3DHbRFYVgTjHT8fhbFNVg1VcoZPiPtROqJ3Ci58V/Dvr2PffIhTSHGC5R
SvvhdmKDckI8GkifCmTBtMZk6Wd99sEZxcUbpH4qkUPh+5VMXXyzSSHDRn1G
qnd/beghUZsp7RxVy2FIfVRO8qTI6y/Y1JMAnnYCcz172AX4aGLHGbQdXn9n
XyVjx60ugxIletOq9xfZtpNfsbwVaK9gTrw7xxnP1j7A2IN9iGfumvBVgyKH
Qmt5w4AJiBNBOgXmPDxWHc+G6g97p8sLonISgHlqTsAnoAZK3GwlKy2L8nia
otUL28K5KPQn3aPtQi2tuA+gi0ueuS9seuLwluezk5Zm9u8th4HAxxgZMG+c
wew/njKbs6hP8FHyaRSZE9w9g/tq2W1L/yf2YtKUTFYpGCTbyvskLvhIObN7
d1k/bnfMv1lK2db2rmon9mN1CtBKu3pV6QTYCEUO02rQh36ityJMLDsGqZhN
/ruudq4GaaaSBgvpYmd+v2uJ4xoCpgyh/GfUnyBV8e2XehqBogn2ABVexskY
8bb4hz6OgTfjkcHJ3zWRUcnN1ywEXcL1rY0cdka6f+TvaM9yMSVef5juZk6q
VDPeUm4OmQSsTVhBYLcnt4lqJaM5NUq/7GcVTZBoKLJWOPYoPSaAoqhWcTIx
3wtV4Qh4hdfp5rAXojobbftpYX65YSsPJl77WpY88GquARxMkktr2WBcqZ/x
TqQ4UvVEjIE8/zgPTp5nwSXD8MSsfYU/iC0yKylTyyS2VWa6VUrplmU6bmPW
MK1oQ1uqhlHU8C9abrRtYeIl9qhd0jeqagaO1f0q19ncnhL3stRAXGuGwh3d
B6F/9T70ALBkrBNqFY4vP+bPuRmTKExz3iXsuF8bsiDWZfZyuNlGw2bL0wFI
fiHrLalTLoW2I6Sdd3kccp5VCeh4MRAiRjB/rWlMY3l7iIrODEDH36sST6W/
225ZGJ76QTfD7T6GVVS2vioO3Ha+fywLds8c7AvJbv+XXfMFcHSQTmxe+o9U
lgcfn3JJscTzFFslSNRh0T7b/+utaiI1w1rZue1d1+iXPkEqpOF7sY43Pjgg
9XMGFdwB8tIPKZFIRgXXrzqkIO725xcll4wDDKWVSzmUXbt1IV6d+q29TdUT
+On6rrA8sayHBj+jU0u/spALNtWuzTpPHiu+lve4yo6o/nbOWNj/6vJ9WTWk
uGCOdd0xSJyvcdLsfJxpm5jpuP/0I43e0wJedNRJr2IxCTfwlinl+ZVn7akz
QK3+rKdm4bziHHIsNHeUC1o1GtEiuf1xmLCDaZmgtHm0B9e1tQpDhlkOFiLZ
3YPP69Vin9mDz1VhNQ+r7VtVfUCS8Yy1+yUUwuCpMeAD9oYsjLZzH6NN4HMM
xc/lWMkYK+Fi21IPTQ8ppN7oLSyKUm77YXEe0usOK9p4Z2xMmoKPDLBL+GTQ
7ux/g65eGVBr1db+Wgb19in3ciwoFyO4lcfS5JRa2JtTCnE7yzDkR4XOOT9J
T6s1er4SGfMXguX7ZX8i2DYIosUutSNiwn5Z7gM0s1UpmfiNKPGdHOz6aCgL
ruzeEEWGz5YVkiWF4TdApXfIryHqWAr7baYXWJEJcfuDsG6IX3S5Wii7D/Y6
fD1B7B0eIEE8iPCrVx5ygzWXM1OknUtCVgglGcEMPtY6LNhTJZSzkn0+gF1o
RrnTHVHe0aOBWwuTKOxVRwZvQIDYL04cOC3me/vbRMtdwmqQewt6m7ZtbQXX
3jSm3NcNWL8faMaalmz2PLpRJzi6rokA5l5tu4z0glZaqCEjAsJaI85+CsHJ
WCz3RCcRNLVvv7GEJVOYyREOXJB7U8zN7dpFiB5myfk8Nwb9T+TZ3d3mPw9m
XabWAe/J08Mvuvt4nHhHVXiYMBVIBpkWouZeSUSI+7zOxLBXV+5vZLKInqDd
PKPgu6kMVbZ+yZtO/upMGhCYXlDxhUMdpj7rz+DNOdkBPCQg1TRnh0V7822j
D1TIbjl59k1qHZupNjlLoaXBEcgrQl5hTaUJi4t0Id/D8k0zT6EAYiTfAT7h
gl9sTJBJ01RuzAXU3wpcgRFbie3mA3ZUYb0iDejQtI4SDtVNdzcyNSd4SSnv
cmtk40k3rfkHfwH6vaTGW5W1ct+18nTMmFGUZg/y7KSjN8f7CoH8aHVeAlWG
bA1+uQrTUL4k7n9n40l53ka4dDcM4He4Qj8PP611BnZpEwBQ8PkDwdwVkdGE
Hh8kJZMDGdeLURfCTeoJ8ssmw/lfiYyOe+YnIPQ3jLQ2krE0+LJdIsPfUFqG
OZB4udIa/P23j0Pl9SFRxUQb7vAptHctqYQHDWn77DQgVUnMyR44LGV+sq4b
iUP0N8JKeb3vyjK734YLCA1rsAea8bzgWsXwUO7uf7z0FLiqUWItvdxW/eAe
9oZYEpU6j6UNkuZd1X6tV+stvukskkklRLcQGnkab7QL8T8W08hDn75iieEh
/aBV44ijJh19lxoTVxmMNsxRon6mImamyU9cj2QQZuPQKz8uXFzA3ovAkYe1
Udd3ucZ/SI9/gOE9zvg4ln+ZSmJ3O5RDHzeTiZxJoz2xk1SJ7UODfdnJmVSr
G6vwcWn/EYwgzSjJKmnx0Iwo0qkl92NtD0+8V8EF31/NekWXVWGy6jrMStmv
AixD60f40+fLZzkwc4dcQWBG1zBk89DEEaHRqwtQNzGmTsdNPL4ZkvMmfD7S
xVFy7rV5SqAJloP1K2Bl9XmjCwefb66dNlY6P8t8deFaeTTV8gdPEH62JDH0
v3a9fotFrDYvhhzbyGOjLwD1S/nR1Qs/YHAw6NbsW6Xs8jqc1Ilau6f3Q4Lr
BNxpJF8JKIx4lkMMxf4TnjhvrJeoJXBT5ADgCE9SR4vfBapZQrRuaifdCYah
KqfK2yqcP9UNz9FINuP5haEsrluHAoSdqgKXs0EYYPQ9T+oZreS27byCUEip
VMpbujx/UOKHaY3W+Yqt86/p407bx1rHi3/Z+/Qq2F5zyNWCRH+QdLnhrst8
TtHEo1G5xIfj/mvnD35HbSdaVcgVFKYTNthkJ0S59qWuxEcYasyWFporMLE+
Ipe9J2FBaMfEtZQgeOJHQK61TysOw2QwkIvRqDlkTdJgTQkL8uEZcNaj8wz/
BySJol3gR8ysHoIlkHcXcW0u7sE3tzOyx6Zadl/H97WhCNkMnsDukUaTAfGy
k/L0FCcFydGMkibJvHOTXZKD3lVc3zyOClLjmzeDsmZi/yOzSC7+WAWgUmOf
3+pb/y1HE+LRkzbCnLS2a+UzxylLSoGglBzeCwX4sPXNJhjC09h/6hZulBuI
vkoxido9nA/aTjd9WyxtI5s9lBCV4GCNkgRBzx7MmeIxQXsW8EGrDNFAeBVT
Y1GQwHHCaf1KxaCwFcs2q0J0Lz7q+8LaRTkJxWl4typbdkfbfZbjPj9mha9J
r7svpO+e/W26Wi6MmyRRKHgtOxo1LhEABZEJr2vcWniuABEOd8zVI8ilhaqX
jQps/7XR/3Z77QemWFBwxMsRZeERIrrgt4KriUQ3SB2EP59lraSHVlx5L9ss
RQXaNFSG+Uz1SzgFeY//ZT/4r3Bk247nUI2458QlspREzOKZKQIrEEpx5ptf
f+I8KtZoLhcJLzgBfXi2vMMgg5o9lp0G1qjCfiEWVYTBOtzIVaLax92RzjXU
vnDf1hxqqrFITNezG1Vlhe17abwSLnnfk3CvuM72LqN9adW8bR8UPapWF4F5
/v3bXVmu/CE/EF3eZbMKUKtH1ftEmXVa/gjAdqW1wrSckMPGPHbFugpwbqOY
xz7n2BYaobtXMeiVdUn/0qNswjovxoSoLdkwsYuc06NVn69axe6K+bxiFldZ
TYEG/NixUCS8+XWFG0hPGKDGWAI1m0oYsKI7ZUDMkvkfaa/RVcu3z4iwvct9
1HJnF6i7g9a4aAoz8WhVbwTdWPgJvrMCKqQ+eS+1w5WYUmylRgwv57KhP4Qp
O1tirv6K8TeFXTMegUKWl+zrLOchDJi9VoeoDzrtcgnaGjVHicmTpNk92YYJ
x3H+U59WqEp+hrdd/GK0DHWW5yLWG66JHNxssWVsfdX0FGZ/Yo+1CJSRRv5p
jFfOZhsG+PSTQ0Sk63KYsloe9D1bwG+PwQ8IlKaFkygGHvZuZzlcv2E41GYs
0g1NSDr/hWRryEDAsfG2fM3s9Hc5bklpfe7w8KnaJQ3rpMc5VlfkfH/zlNjF
DLNktlOZzwc1p7zCxNdyap/G23Ndb+9NrqZPlA4bN5FEJtoV4a6jrmxdH7tt
jANom0lSkQJ5vbIRqLDASVHmMCQdF3GC5L68rs5RluFxpKf5TIFcWyOLvTq6
EuUjlj8/ZX8p9kdrQNdlQ7Nuo+Ngb85Sx7hrF173Q1uiGl2SuPf3qyeos2l9
M1Uw0h+PwcdWrB+q4LIluomrZpu9FY7c3THgGqCVnk3ZhHGFt0b7qTmKMHv4
1ncRNfCB2W1b1kOYdPyhaMGWElFslEpi2UuEAB0XnpEJ/VxuX+teElPXX3U5
chKLbrDgK0NEppTqBIfbjWz1s+bnbUHiPGJCAwfNeeaxSa4EoUaRHhMWgs/D
0Co5IzJ5wiGWwhZMO36DO4NWk8NbILV9mvSzHdV8FrDoFw0ywgoPu9BX19HJ
oKArco0ZFM2keTyX53qKtV81iKApfaGk5YfB5PJXM8DtlqAHBOqLn8WnxlAG
yCoDhfYPODxZ8Iu7QhN3z0WWjTpk+7ymh0bGeSFMdzNhDNHonHZZ+XqSAUTx
8xVNdD/YhbKUkWsL3yHkLJpacOvypTWVvRmZdydMfMlrXAgnJoStdJaHlEGR
3Zsd6TsWacePBPbY5UBeKcHf4Ih4ViRfRxHAn1qFmv/9Bq6OYVmMubNQ4DOi
dMkXsXaNjHmrEDm4z1bCEy/TRQQn3Ysqym8xISXb1ht/6pQqyYQiY/W7Md02
r2rfFlwHT52Bs7nlF705hdl/I7sHkxwjM7phj0jYuaIihKInMFjgS7WGEVXn
xD7Bb4pf8u80JI26MtkwUAHdIioax9CW9+Kbc1TaovZycJsVBW5CiMGD7f6L
EPkH7X33wQBDbrUMdL/qekwRrrEFtbdfqWMg/rNjtz0TUcdKD9l6JUdqikAv
77gKHFRl6MARaA/4tOo8RhuNKh4obkZAefWjxwWxnmV1RDrtzCzTC3IWA++F
salszl9YrNSKAyFW0LEXIYE4uKDPEdsl0XiSAYcjctm+EoHqdrWeiyBqOqbY
gthZuGU0Ay7EneJ0Zz+A/uSTppCfhJHXbtzYakUcjwY4qb/uli8wHbWBQTLn
qEi3nj6oYOQ6kS8TYg5V95e0ZDbfRXeNJ9oicYOK4/ALuBhVkuwPV/N/bqjJ
7dAuVKA9s9IjoOZnIhjNlNw+lbLEqVXtI8l0Z98Y1gBZwoHaHxRTYHTsm1mg
usLtwV3SNc1YAZ3aCLsqya0zg8rWKZWhbywx5yrWlr7PYatjTrq4etJj2RlO
oyC2hsPxKMQaD470qp1uSpCoZqR6FOrQIbh8Dg3Tg1/UiAkiXn+hm1ME/Gdo
OtCjuItvjF7rWUoj4eNI1hMUAIZaXSyivUz/AiBAJ+XGSRHxFtzbFapJc0dq
73uLB2+AYNuQVG7CVXuKUI6002nZIuMs5+JYO2Q4V/uu2VLz131wQO4FQ02N
jWfmBYGAFuBgJMVJmntVvqn0qrDXggNFcacCp6/HKY8yEdtMiUzQeXbdAzC0
GV/rR7qz5KgjQ2gfJPRg6YN1lHypSRfR0dhg37PNYDgTD6tHI9TjM0DDZVKO
1ILsRIG6/Sua9B7bOWeSAfvzjcXRPt4tE1ziL5WsEJVC+UTg+c6l5Io3JQMF
j9ygwydpNQTWK5HrPVnXlcOTgRhmnruTpx0KAmovzct3s+jEe7Zy2iUbTOv3
gzQM8o4kAZmD13QXoOfHAiloXJVDokaP6yGJLe0GrZX6dMSR7RfgtECh8v4A
5layWYGQFCcH+ywCd15tSrBZOla3oI3tzg6NqmM88TDycl/lflyZQ98SzP/C
EyVjiCKyrattWLPXUhPtpC6h2SKsYqu/wV/1g+lETP9eLRRV1wzBNfyc5YXJ
VpmTBTOU7CRjZ7PCp6ull94xn8gFB3BAZj1YHoid+3gfXsDoEuZyMMCWElh7
dFONhi/NbKFf8xSoKi3KoArMX8ncvsSszZ5l3XidEOx3SMju1oC63gBtQur/
K1Z8DEABu4B6LcLQwp56gvq530AYz4bG42VJhrNiq1qgAyw2rs25fGC2KzMF
YkQQ40WS8UTa2kpV5XTtAvohsgmPnm+p3LBVf/PXEtcOvT6YbHLh9JB26l+v
9q844CVpklmYFoaJ+BjGkUSrcjGM7vrQDGutTDLHuqLIyWi1LDAGy6AaZAdB
2xT7jgT6I7NOvy7hWIpxmNYSenBq856jFgCnKotu1RLrh2/FhI/dXNulff8e
kUNkSkeYAi9QaBFa/GX1SAjzZuJPht4PFr/xh+KuA7cYlpYKO+6uIWGvvrtX
rD/wnv2ljV65dFIJLUw7suO9rA4QCbA0yldKhulyudJZ8VBgHBJiTluh0QYH
0YlWOh7WRPDJrk6I5Jsl2SpHrOCwQG3Y130Qd5op905KuHwR4z/HD2t9xx/p
5uO6aCMSgH3/FjpT+9IHZ5qADqGdeimeGIA2dCh+SyJR+mgvTK1Vt3QOmq8v
b+0PXvyXyw6fkEriT1KN7AUlUPe+6w+VtqJZrBgodYEwIvNkut8RFSy/iF1M
cxvAcsyB7bpsRXEkpFdLScIUxDsFZ0DV0OOjf2F7C0BNhizEXlD4XthQTghP
sEgDOtEF0S4ld2TGOUEx/Z7EvJ2sXZQ/fIRHL1ADc4kOj6V4gKSf76Q76tJc
TPN8zEMPD7D3rPWOdHcG5yQ8bVlBwg0OoIN37rYlyz1shVLR3jm0kJZHuVBx
AcoyZLuSHdFk8XukK0V6zTE5ozUt9vJUpl884aX55jU1mIrI6i80lPA2+Msp
VzBi/FZ+KWQwgJIPbb0w40gfImme1Az9lQ4ncFyxDMaOsie8djEjqrixiGXO
gaaO1DMLWHHq5j2qIEolXN0qKdpgNqcdm1f/UEUeGYPPltseJw3SsVUjEbQf
cn/U3sq0I5d/xWL1c2fc2z3KA+a2AUZYCy5UqR1ZlxMPcEFVGuZwfKBg/eh1
h8EGlIMphbMzc14CfzzLzZUFZxMXzs14FszGz9VtWwYZkbNqLJpCpNSOjGqN
QKBUnTTIArmo1vz0gvoeHrJpkpXlbvZ5vPpvxo6v+FaQVQDDA5RO4Ouybd6d
I00SXeeYcHdZlDqLwaSgrc2okupFq/n1xF5xD9Ab2uDQH5VGMH5kVI386fLg
LXJjOlrjLJqXH6cddLUQeOuRS4n9VBZuUoSo5N7TkNtN+itSDD3QbbIh0896
rB+0ijU6SmMTcAylUl0daQc1UlFHiiR/tG7pi5Sl+TCz6wpZF833Q8BmWmkc
vBVeP7wEYbaLhNvex8Uo9XixzJnROA4duYJgib3nLRy+42eaEYIN3+Nywert
ogmxPuZcvRrZyTuFO+Np2eVWdzGSIZUqrMhiZJh7i4sWSioomOQMyPzpEBaZ
1LYyzDpB529S2mCHNPZdYpkLOOpVHDzxszdePWt5KjqKf2sfIcMvlvBmR961
SnRx6B57tzqvrHTudgonIHq0O/CYwfOyEMfEnFgIkxq+Ymt1i5wpkWh4OjjY
xm6Rmc9Q3H3k8SQWIx4aVnRuG/2tJAkOzxlrBBYCzdd3OvDYG1kziXvtfLmk
oxYF8/ihKFOOIlYUBbDMizW3LJ0K30sDVGC9yIac+546dJkHTmqpAMnCNfAg
1DKc9HmGZKbRoV3SOx3vkxrNDhMHoJu/dmT1gR0kCFwuYFxZzOUqzW0ROXs2
Qqdz3pTp224oePwI2vy16c5vV5G1vAoP4LNZad5BJQw+1mVNLtbFdor0K0hQ
JZJTOYLfM3dlJqotIvkGgLXisHsNTjYnrLXW6rhzrwBW4S3MgcGWTblFZIeC
oNIm4VH985+isVs8BdAhvxMKuOx5e4dpaSeFUDhGqn5DD71gSS84iliVJICK
8kJFELQamONQr0dj1Z4AITk9bEhDNCeu8r1hsgkcgeB7kzepSD3BeGrFG/Q8
eHdrmqOFe/DITnC/6D/o8MehZAbRWosxW/t+67Hs+k0rPPLF+GCPmVcauGii
GD5BvJ7AYryIVo9ejxtScVvS4W8gZZg77FTJsajeJ+/rO5fOVFb+BlsdDpvG
d4pN2moDPyp9iBadcrzhrwSSs8VH/sJHkJcfCEjJWj6FLyXJErPQ4wB91s98
UtHuUBEYcKoHyczAtCTGL05NbD4JbmxSwOT9c7rD/2MyYMtw5Uyxz78neU3Z
cuxAvxI5i2MmptqpnhpObvYbpks1IdiRM30cz38gtfc6+kpaNn/u1eR3pNJp
ziuZ30KNjQXabOekyFHgRPLQkBfIm793wZp0xmzwUJCcplQJ1tAK4Ik0JrGs
L/Y/JMQJMmAZF4wS+Q1f4qKWkAptBfSAZ2WycfjkiMQWVVFbCvjdBjX4b1uF
VneohglIWyhHUYzjeYO9ZTt9pL6y0AZ2B3Hz0Tb+F309p/T+BkuQQSkXpr+f
LSSO5wXip4x8ikymoum3NxRYFTq4HYZaMQbAJS4PEWNMxu65VPMkdzaojigQ
ioIl1IWczO9qCfkZ2fgK93IiftJTabxNWxI7kwSaV77dUpZqXNtfAwSfXHWF
T3hDWn/hS6pNTw3/NN08oSmApai6+u90hgID/AQnJwETCIMTtON1eFt3opuZ
RP6+oKLUV1IW3tIgZg+Rctnh/5JzlpHR7A2AOtCl48BD/I8DyWwmdREwNR/u
DZ1vP0GO5WALZQRGjMz6ZabOPyxmc6IHBUt9/2rYqdPSHPwT2S1sTS4W6C9b
/lVCdYVFb5kVs5C2cM+l3ZFvOM5+lFdMLd/M9Pm5SEe2VYOAxauiHwv8cMTn
zVSypoHuMXYh8PCyTsjp8uOUiu0SrBM92wrvE9gH5uxP8fx9fOryUt/xtBNU
uNAKUCANVyAj2oHzy6tMoKEuFMJL/uuQUC16IRt1nNRFfnTLger1ZYm6ZmLR
kM/970VLVGJwLhZ0XhtUACikOEw3/mrTOZ6hH7H/oweNumjKzjb6w9d7IJuM
qg8INwxJ3H5WuHsq5AZUCtlfTYory30yZpkGSMXxb8+55ro/X6SYYFbRqq+V
0FF+rzqnpap1L429ko6SZdyMwRdKQXIqCT993718kBu/ro1nPfGqVGMVsLZi
w0XqHaEo1wNPrVZnIojPmYgDCD0rBKM4dQ+zZS39i2PSSFTNMNxBrU4GtBdW
YPug0sNlLHhHB1Dqil/QnJufX7T9K5+9mIYPbgBrp3ZqNHK1gZd9vThQ0Qw4
htdP91kgH/egQzteBd4LUyiZ9JmgwOrdbaYXd5sPf+hPTxKbDn8XkVYCW3lj
g8U1lKng7BxWcdXSesz/PQNpMY9lCV89h4aiukSTK3gQEw4B0q7UadOgHTdf
h2uYYPSyrTVmGSa1u5/zixcdJ8Fu+8ir5i6I+tdjdMykS4rY7rt5/KKRePIV
/TgcGgpOdU8JbzR9RweHL/gxtAdg1uQXlUP7JwvVQVYvF2AA9jonaHj1Uoml
Py78X9XJgXgS4zwn4+ahs2ZQDEhvYmgIc+szuIjBVUy9tXfEuvyNpZgKC8D8
RhTx5lRZoCuJRq4Rh2RuTkZ7QMQkhIxfy6DGBHRg9KSd/d1yAMPwWmY+/Qkg
NbbjWCY0u70PmBe0e8ClR6kRVYcchBHauSSTTlcQ7d1qf1FMrBXStBnP2Fqd
Nm9FJJP7evMpbI4+1etWvMY7OjdGzFTfniGI3QrzJfjTh2wkKUKvJq/qQk3l
IOEy0BO4UJ+yAAau8lIlI+hZr5z6Evfmhg/UQtFC9k9VYCT2fAS4lM2dMJUk
ikFYcbfVMpMTuu8FIxQrdrb+3pC0oR0GF3Y80te0R4sIyQe/ITYrVEhMtyle
8i7pCmZ3g5rCSVLWYAV5NxdxnHDm1v4vVxqKolKvh+ad24z8kqcxvxHLdzyf
AREU4Cv2uNm6Uq4jC2JcsN2g0gJ0+np7CFSqRg8nX2BSNB7fiJhxhVvQSxLc
DmfiBlSL1QdftOj+x8MlqD8p1DUBl0H9kH+EFAQeR0uSJ24F+53ZxBNts3tz
N+9VqCoV78cL02aZhIbc5BVgZfFhNaJfajBoDmjHsuWQln1o5kJgWCqQrqRm
pqThjkptLMo05glScf2WrwXzNugomtMqZi7Rz7irpvo36Vpbya6IL7uTbhhF
oPItSM72OTCcmJxUJnchDEP3weRXfwY1sU0kkI2V6NQoLaOEUaooOtuMV1HS
eey+eeMdSJ8Qql2K01eMpitz2FjkGMnfC0j9RuzuZFYzLyCngY3hSWNX6I2D
c0N5M4zKGx1NVvIpl3/g3bDaMnigokg64hubS4FBYanmu9WHtLOGAq2KUabJ
TNI3txzTeX4G/Wnmj+qJEW9WYUp3sMU5h8SHju1FCUaDHf6H69AF98spUSaI
dymbIJRrX2USyTh24gthn2zUV0Jp+1DIRuYLnITkqrDMGXpaQ26u9EpyKLeW
GqNBqFWYTQrHeAljzft+8fg+yPTMvhRnJqJ81Wf9lZEZQ9gIHSkgFQ3IoRkV
6zEhBKqHRyfr5tsuoWhPZAWRpHlR6ym78rJr6ErUTRV317OfEywIU379w6o7
JQQ2SJpRw1Hp5M3mT9sDeQn9+fXPs9C1n4jbq4SuRhfK0bNh1X31FBiuFno4
84OaUwo3aJpdvn4lSb3qFzexdfJ7VeB0ufYu3C6P+b2g1qR99SCcRzWGy2t1
aXKrq1eJFHhscp1SjzpuglWRKYAgCegMtVQZ4mdcWrrV+uTJSg+1C6P3mehg
0p9qpe4llAk2ahusCyepQ0VrLKf5ASdMWSdqlI17C94dpapUT/jbcc4lv/B6
kThcPOl/nXINXJQq/bkvx9dz8IuMRhIqm4nGPJyUplN2M5wFvfdin2/LhytL
Q08YlqeZlLPqzUpYbRa2YQR33aCEJRn4JKlTvYegpPgcRL0TDtPiDxVYgGID
HNOCBOXSQQHGCD0QK1dJN60ktFaFQN0orSCil6/3pgDXEi2M3yWPyODEB/oG
Mt38+pOYsmmDZgck7S/peZobOMw86s/zf3e8YNg2NrLatz7IaYGg8+Jl2Xf0
QPXKuEamWwM8oWKVwDSzjtacesse6i7gZEQZsSW5GYp1Om1VkrSkO2xy8S58
2EmR+rImkwr/tnOoGoL46Br0drJ7qQUrA5VlCvNesbtJQ5aY/KKbbGufCRRy
Y+dzJACKDULlIj8LEBzjVzivhAuatWJH3QNSi/Ei5Aue+T62C/ZneCoUlzAA
Bub7orNtmBV0LWhyWELyqi4tBHPPES/eNfRiDz7kAXygbTBA6R3nBK8J395T
IP7hFLnxEjIEoieHCIj11z+kosWIRj4p4nw7A5D+bvifBxGeSqP9nsWy//ZO
ub8sqL35x7sN89U7mlWVHkkunQK6qWKU1yRtnsiBSdJrw7P8Mns/KFN0Gs9E
vMNFKV/X3pz1fd1+ymJYmjVq6TAHnPM4H5FJumdTjUkED4J9UTnZqJ++30Km
bD0Iz9gOuJuZipaaa5aF/7+FYd/jgZ661f5BjxD6mI8VaR3Xn6RRL498S7Bl
6likFHHkwWCkEqxyo7Bfmn4W1awkcGl8eCgUmn5IQthgaLve/wTBiPxaKZjC
0X0aaZ0RMIuvNWquRUgQUPK5+Kk8ppQRYjH9BrKi9WVijijOM54TrxeN0Gkb
cqbgNfENaD/E7c8KidCFZbBCPKTfPYNKr1N5Z33mWKbSTf0DOi4NNLa+VMxY
HEmSe2zenweVMVDhyaWPsqgCO2+czMUWPZJMNpZV64RHnX68QiLtELM/csTl
N7Ot3QHgUYIl7nzBG7XweTNjOK6D/7Oe5xR46yvyemM4oqwQj166v2VrSO2E
py9ztLVSEAob+dMXxUiVXeJ78AEXAIesES2dBRt2eluc7y3uQtUfBvlG70w7
IJB7t9EVOzgmghzoiVGb7zxaZEEXD8LBHoNxzbBSDyHM3b+LUCvEWgs3CwvT
mtRxR63tBA4g4nnoEWrQ6SVLestJpORH8XGqK9cqIWMelnmYL2I5sh7T5F1M
qhpfyRofm+/PRDAZgvI/fYTMfgQ8EYfvuvcjPpoW7dGUP39+P6eQR1hlmLcd
7M/EZbpB/FFFRj593fYwq1b6KtjTcHKydNdOuNtS9GjgJXg5mCTB3TUeCq8/
GYhHU9VLYTRYoTl//qH/80W1sAz5l9xYmYM5ofnlvApnYIbjb1Leapod12kq
VnCgaU831BWC7L+RWvm1u4ngKud3KWtl4Arm16oEFFo2zKUCH9VB5bUKKkb0
MO6kWUj9CEr/ekXPj5LPh79yJ3rFVsZGbLxaxVDeOH7h1M6mj88i63YLD9+4
EGcYuhvX85S62pJNIv3lCRWN55YszlGMIj6nG2/VNq9wOgnnQF4kJ/aWyOF7
AWGbB5n22LoxqH7snh2O6QGXEvAgarXSccfHnq9Ac/WskfVL48MH8hL3kB1o
i6+4scNdpqrxPgLyH9NhcpOfkQXDTUoFw9WULU85LnvLRjeJRM1NCVgC8Dga
nJLGe2gYn3UQUGwrS+pllonYeZm1v8XtPO090FwkPEFduIt7dls8ME3aEv2c
iKanoA8rJbrqrQAcNVWz86CHhqxGvTwWinZoLmrKKRv88wkFzVkhfyiO+SEX
o77kMx50Zz1usz+Sxz1ItrqlONYpNQ3L8R/8faEPlcJLcRc73l8LvvJYdP34
e8Sy1RfaM/dtEopA9wUBYg5fudXDL9Cuf3Efdz5Zj32JPOIVwb0E6Syprt9m
kneJmEjCGN42wdIji4san5YUloM44DOlccR/7AJKQyvX9MqsUqz5HfCEqX/m
Ba7Y9sso+5ofQU5ZDfNy9C5nu+a/980SmLJHV9UB9zjlCwmzl42T51Bia34U
G93bcuBN6PuZyGy4RHwGXdgx96GFxqLdQQtDCZKhgAd2I8AncdAfvRe+yD/d
vzVS5auSoaKovWx0CiFEzVaQ+0NM5nV4UO6m0CHZq43t6dABMv341kHjD+gO
UJIsfabQOe8FdN8P/S3Hv7aToqRgtt1EgaxrNW41r9JNgQ+RPvudNPJ3fjPU
6/3xvS9ang//6pnPq63f5ocmJCqaYcQrUJbPZmwsjFYwEW5GCxepfvXn+fgz
ALUKByLuaPZMfyBeQsuGPztQ+a+pRWb6rQWQo0UHNS9BZTbAg5p0n5WOc/9J
LCFXpTEmbu27lTJB4hUzsXfA2oQNVh9iGdm2/BQ5ifCmddPFQ/JtM7ojId64
AsN3uj//GVSADeKZgv66DXg+3Oa0VgPdPBAqVIOrBRGyweeTaz2XXlcX3DDU
t6Cb0ALfJtuEieaW08sR3vpxpa0VheLhWcwNR6K20O1oAAfOUafdpNQuFQbL
UF4KuYXOAXyyvhLy+CM2Zh/nt7OwmG/xelSDRYHtVyZdLKbF88ovD3TQvalV
Ti13lE4543qYPhyRAdKrhKH3Fxu3vQyFZmd5TTBwO0wrkDPlSnn/nR91jaQJ
MAcQt4aABpV4BX3BZh8uleIOT0SR+ABdz8wiZZF20zOsULkIhTpYY85Cgw9A
2IO+f6HHh8jN3jZO6ntDvAG/Gj+z8COlUIL/UPlxJ2f4jYIfNQxW96rGvaUY
kvD1iqIoeUYRe1oO2/nE1rzVrW832bOgB7qQcAoJMs9UO74mJJ6yqJ2uV2ts
JuBBxLv7Z604KCAYr8FIF3Oh7Jkm+R5fAr65Eu1s3SBK48jrkMC0OFXH5PXe
4PwOIPd2pB520bkHSagj8h2tzzMCNioo77PawxjhZukCuqhd2XiqCt+MBmzI
n2Npzxajhdb7UhyRhXdDOXSkoV1hA7X5JVvAZ7RqNfSmpERnxrtJ8TmJJ4wa
MEd8T7Mix2ySa2STbxYLrMwnop3rq/O4NaQcgSe8Q3t/frUO68kNd+n2L8By
ARWJMIXEdSaNis6UtDVTc8yWpJhnpX1Tm7fYXBOe2lkTCnacd4eWiYCwU16P
/l1jDjsgRr1boyza+fPvL7cJad61dvCLJeYy9pXlhzqsolpvrRJP2n+nNAlg
5f/pFbXbovsX0AjXSEFLLlIqz8n54vbmzPMaw9NZ2m6/yNQtJrwlK1Hses1t
ycK1QFOeiEeIpUlkCoLm0f6p3/NIsenuiJpiiXZZ7uzC1pbMVMWDuP2x7gxB
zjnlnhJmE01lrFYbVPH0W/vK0jOjkaW+J85ZLPtKW+fwMj+y+FCpLY1rxyWP
QbPRGKO0dYRRqMgBnUYqizDhdtZisL8hLk9ORmyCO9AUk5y9fljCkVaVCqK6
OP6gx6JKt45oPdChBoUIm48tg/pOwBZewn9uKEvXsoRWwrEB/obTY5pHV1lD
OL6805iPXTaWT2ABH06unEAl1djJsQhPeNnkeGN8KOnXGu2wdtcJvwD8C0+c
RI0ZLNyhkJsokvKHbGXY2dcSJL3g1pMywp36YIwVV5k4dl6mVytVRrrkqKmC
A7zmhIxj7L+Po51apMCSft+E4JMW0I8lWYgec3CeE64WR0YY4eb/sTJedxU+
EHliw8Y7ikXfK2qofQOSs8uIcSmEwpqv4PkQzSN5nibi9ayXGi3l1YaOYI7J
XU6Isi6KN+YMxXTNzGQ4JxgDsYOHadsxEyfJir4hakM4xi3bZgxIE2HUNnRd
Qp06j+ufDNyFhVKoQgFxxVANB4ItPXXBFr0EZsYpK6L+0XP4wrmwkAY8CQR0
flDAnu9Tj2WhUvmxxV5inYSMJ+6lOt1AlrQdub9Sa57kfor8ocssKGBeZfyv
G5+c9YSf+oJmezg7zqO/ujbv39BKvBZN2gXiHivqzcl+D5splYSF3WKROHZe
iAql66zvAd7DM9MgZUm5QxmJ2mbKxoG4ton+bW1JtixPqPcIVMa6MBFKyRBW
y80MCUePbIBt//yBZXO+q86N6fnRQWmxnjOvsjhgZSFVy2PERajPJiS0790v
jQFP5BbByFP8QHTUVHHyRUWG6fEIvB2HQhof1q5UAM3VCxqf+cJDWePxFIa7
sJXLzQ+ljRfotp8c2O6rAA12xOWqElQQQXblopQWqAfvyQvJkti4aOs+sHFO
H2yIvHeQezxAU9RTKXRsmTA5oTwUfP8c0yhpCPK2CWWGeBM6tn+Mj05h3vNq
xuFrcLLHlniJ4ORywgOynQQCt8whgoM8kF0LP59OJmBmKCcnNP9I2vhV4FIo
DZX3KVV1R2UrIg0J3/sKauazWdPCaGL77p+3OgUxCG+60Sfpy9C/YlZ0+N+L
yFaVEl1MOYUAAefYJrqIdY56/YepIh5hqG9NfgKBbkQnwqHoGOVx8eMzl79L
pbwmR9ZDo7HhbYUAwkOEs6h6yy8kgUtK3m1cMXwtWThm/drg4hX6W4/I/rNm
I+ntom+zgVSAt0BTngHD52YcJPJP69ssSqoHLDAWEf4qWXSxQ+qvBr0O2r43
WxLRNx2jbDJTp/CemGCgwkAqTwrbh/Op19NcytIt9wmrOErAmxz+Caw3kkCR
tcIgdu59qJhKfjm6890Aqz1HQfl6zYtJbiYy5dHfsX2+D9R6v+DmHCZpeNcl
5oAgSU5QxCDq4IkawyM/sjByF3P6nXRA3zMPYUlUHh/LUmFCXpAdquGw/yFV
Gh7tt0bfBJA/O2FBuqxsM1+ILPQdoxOEGvcBxRJ2iWcHMZyDs3LLu0u8l3kZ
OecW+wDD12VRtUP+NKuGa7NzkTkFjsZ72F1M3s8+cxI3arDb6Y843MEZn+ko
ccbpUDvFqp9ZPOBF72LFimthEG+f/Wkjfw2NWbZs/61z1yy/5wr3Rch96Oj1
0QkDmpNyzK7njUvIh2rG5JW1t6aaL52gMlIb4jhoGftn4GJLWgWf9GQH1LQc
IwDvRSlb2OyTRrhIFDoOAvqzI32yxOzegWZbsBsv26tH9mk6psBYwymvOP5n
SMu6uQ9o+B7oMPwQl0labpWrysNg1ha1VKyo0DXYVxb6iiJhYevLHECqZwCe
09qPp93tfuYjelJ7+vxhRip6Wq9abJQCfY9D7WVRd185zagi0H3QZkTr1xWg
Vq2S6AwPF/zE1eXLVLgECZZieUy9RmZXsdF89fGuuGi2k29voQP2W76glJEc
0m67Id1FyqCYIWbsn5hnb+FPuXbqsFgLMSpMCu+mrU9BIPohxV/hhAJB3QQK
egJVm2BazkWZMHmQnaEwatpupMxKSps/kh79L5t9al46K4nX7VHHOSKT2Htm
hrp7/CLA6MqmxglgobA3i+Ss0If+yBWzfsrX7g/nRBykOMiRtTxWTU3og/7J
I/Y8WZFtq7LlhCHU4FyCeIkHCJkG/U6Ud2v30hYfHBqSolYEb/Pa5FvwE5qo
PSVrzk+SmmKnIghHTO7hr3dd5zfYmEqng75IwCiHSEfh9Ta1LjZEgBCFsceD
ttDvWwxPdwHehdQZyiFYVkaeRql/f57bIBG0HqeZycyet+Kr4sRov7YC/Hbc
GzA2TZaHguEPRRnan/Y1093hjyN9L9P24FbgiR2LRgu571HpqaC4O2r+RP8H
+9bpgnqh1GJlTlvA6KMBESMtEr51zPZSnqqiaYYfJyI6/JJXCi9nEgdP/VIv
WSg0OQNL8LQEMChgXNwCEtN9cdFOyuYOrkaNaCipyIYnw8543heYLankThmb
yLT+5c/I8uwxRBIgNtO+ay+eSjI9aWbBPZMA7DFcgxkCbZr7k5DqgXMVhNIH
/wVudoiV+RL4h0cd1pfACw/WvKIYW2bHC2InrZ5F9s3SEFcGz0i9pX4Njhy3
B3x8BvBhCvDS/WglH6woz469OSyFzpZ8lR3Wh9i9YmOGChe1OMUQ3aGrATTb
7ccD7VpZcsUyJ8+1CMxCVUD4NVxUxDb+opmryYUySbcHMoTWYHglJIANRhA4
miJkWkHTZJxHOrUxI+dYTj/p/DAgnZ8G0BGY8Zth3vOUUibYRzgsJbAH4BEJ
7QEUjgWJRjlwusVzyIISdorhnUUWKZPNnYe8muMYGntB8LdQBn/WRVDdSD6m
g6E25AgSr/chTO+vk0IdlbUMqMAzWYtK3tPYhLh+NZTkHAGls5h1fziQXWK9
MGhH0wDuylp9xASiFrdJZkfm/vV+5vJwylsCVRxxCcawO6MZrkx/+7BqO7x3
WpqEx/+oNiyokdKjQtvLkTHGZtil5vLCRTvte0b7/cIMSvXLRo4QPKdNNZwZ
MISUmLAbz7qTg6ezhQVROs9XGlOkzcIeTxDySOeT/eehLiCTooKgHWMhyW9d
zkaPSRB8gSu+9HQKsdpfAS0K6taKSR1E7W2LBfzZqi6OE2alSGG6qnBFGV3U
llxTgwYareiKHS5cfA1IpNJvdsvSIFOfb4kLyV34zEZafC3Za6Rla9pgxz7z
67JxqCz+rruyUUfxs/cGpZqc75mgHFZs1yAK+hDkOgzTucqn9W8KcrKVg2PF
slsshImULIDJwy2tu9uoUxy3Di2RqjT+veQ9rYL4UXrM5B9hzV69TxxRzycS
mq+GcUYN/4clc965BJ/P2/1yCbMIOg2DTW03dRHglTrWPoVLJZ8ES4axyFb2
9ml/mfRbfJl8eXdm/CTTsbZtrrTRgckFBQ/5E/WcSp5mt/wWSIeyaQzeKRRs
MKfaykXLluAQ824Z3TYwxygovoCN6OM4o5xo5TBhFJOf4ma0vJ06X6QD8zFF
eY7htxHl0AtieUpbVIZy4gnHc29nuzzzoQkdUIfqRcmWYF7g37VyIwnRENVh
z0mcSpXqRyWKpix2LuLAwjuW1G3dedzZGvtD8OfKQWiJwzgb5HGcLi9lpLf/
rjKd8X9HWLJuiYtH7H7b8AVkL63d1jHTAT48jrCxuo5NLP6MyVYkuzC87YMw
T2Tudh5GVeWUbkQUUOqeiIq9KrUDLvfnA5L5byuDJCYxF5q2BDvXKKA005sy
3JSDKA0IESNSjGRdiHnpoWUEiHQw+R1JB9pou63kXzF8Tlr3ig13lK1eUcJS
KftyYFHnXL6dd99d0IJvu+8nRw0+LiphxjlrDSdE4nrvKQ9+bkD3Gh3aqkZT
N92CWLlU2267ZA/Xb57qn4Kr+Tx5H14uwUQWmC36ISnxcEGZH57d72oGP0kH
Q5dLxEK9u0vGlecu4wt5k78RQun7Z7cF94Ef0s7KQP5NSBTkrRipN0Z4cJwy
QuTeD3/ISkwA/7vCYkbrur84/X4mSqVZsZYW7KwbjIH86tTtQQP9cxpjE0un
syitZIG0CyHcyaeHGWjl852Eyn7qPdEuzVnwhXFNIc49oAhVMh7sogGUPXSt
v284MzMq36y13tc8ht7jFM9sBt9l9tzjILHL8Kpou7xtzbvRzhbfmNFZYE2+
SGr7P8pveRZ1MgDq5L1xgOk1hJh8a/Oo23CBigL12Oyj/GqeRfZtXOCRh7Qz
UagOfanGWMvCH6yi4MWxm7lPe9+D/mEqgX6ZVUvqinp02yqyFltD3XB3nvHr
9LAGt1Nlcikf+ce9esFJX56HXg60NNC7Cuz1f76CCSfZ09kndns0tQjXVIrG
EKQUk20ED3jRmRs1VfbL7j3VObNKAiU1bfgRzY4yBTYLFf5ShO/SHqPQqPwl
VnioOehtiEajCmzb/Q+6sy+zii5vNCPujesVDYnPgT5302O2sEX5X/b65xMv
0hsh9JzMGJX0mV6rKmHcTYYR25Ixbx4x/mknwwqlYJ/k04y4uWzfEkPePNVf
OSrvcV2gJ8T4udYyKTGsRXXqdH3SMh3NjDNnXoXpEKycT67T1zg54HmAwYyR
2N04INGId0ujqjG+ho8ShEXqEadRzGVpy6rO34rOBaTCzKKsUu/0X86S9F0q
fChSRtDDwk8X9cd6z3dp08wPY8Oc7a2QFsfuhF84l9pLN42A8UAsLMYbG1sn
tLMfpkvbYbYIsfdWlEsLpFwgo2vvWjTbHPoZ+hk/Act7j5FR6VLC0v54Oem7
PHPdADd3ANw3kN7I4qqi3yn4/rG8Q97LzuW9DcZ/ah9bWFjVDRP3uS0tvA4B
Ew55xTQUZUQVOjappZuWI1E36su87NdRPUa9jILVBL1c4zdJ1E05DjIozrim
hrschEpCYt+QLghO17bztxYsUxz+MENxyHCIN2gRGb0+XlUfObarp1pqgdb5
0Sam2cD4Z3LEKzE42om1BxkuZ+1SHEwoR4WKz6UYq66N3zcjqNZp0mcVUTwN
yoiTt2aG6U4nJG6tNsF5nJO55or05+ugo3Vwh3/YF1sAoZRdkSEa8ZadoaYh
cgGvXp1Fhktwnmt9oMYNE8C7tL6B4RSktIiyKjfDlDXR1r6GH/Nuk+cOcVeh
IU1k2x32M2v51cSsMjfnAwTCKU7VFlQjHxXQEx3TL5eds4naD/oRqddUy7UM
Sy/UFDZgfDnZye1/Qv1NiCAdJO+/pSkBsY4wUNJ6oH39S7ySxWw6oM8qmv0v
aOSF9nnQraW1Z/3JreMSoIIn/fLRflfXmjZyIZ3gGMnuR8Q2ewu8aFaK36Mj
kfTAYYbpNpjLRvIvfZ/IEeDJuf+Mc0BLdaAWlbp8hTbIjj1a56wPT8RcL9m/
0m0lCKQgcFpxN1YNAnrYSzJtgyXHhArIa+osMiDwt5y+COnXDREQjAn8isY/
UofLkK3VacbRSB7WP5qEK/NAJcgUFzrmkxJ8oyNS3M1BiMWG5o3qhY5LcuoJ
10mJPMoT4gTUZBjN4YpQ2xI5v+11OAyPigOx5+HY2nAOOZFx+y033VCMbI4M
svPMJgxq46EJGlrUg9GS8aDNT0AjSqdHSQv4P6Mu+ni66fk7QheVNrtpCcpo
tDhTNI53ovnL3uH5KYDzARkqJhe8fQnueiV+IkCMD3mSiLG38qda/IT8F3MR
Qq1M/09zhqoWcF+GQAdZAtrE9CrFhPo6CR66v5xqmKbGf930/kf0B2Qn+S8Y
TUsmAGoKr0nanmoYOOwY829fPcZuR3WVVAhnHHFwxDd0JZbBGbKgPAekCo8M
smx9K+okISWECfdjYaDRiDHCVuAdmav0aspmHQDYQB4/Sl16XNiGgrjIBjut
T53b3bcpiwhkYK05KRikSx2OU08bx0Tr4yFY4Nr4bZHQV7OeJosI2gh5vfB5
04QnGuDJRONz2UzDLNujoVWjGnVBH9AvpxUSOliaq2z2y7zF8BLu0rqnLAgi
Wkb9PEoMorFfCipoy4+XG58ekFGgYwfO88rfq+cbw8gd8rQguItUH1SMNt9K
th944wwFkswBZVtGAvKth9/DM7vFUpfn6+DkCWs45LapwNGBkRIRlbTATITx
3ZdFOYeTu4nV86WoG9tZEosld1UJgr1YtG5eUNW4pMGCIgAHfWEHNP9cWwp6
OnqnDk04va72Fd8Sk2QMTUrqoI1xkeLNphbBmfEpi/jzq0KAZCYL2E22Lcje
eLaaYn+fH89onyE7WT4UaeyP+nzLJd2tBBJsp8nBy1vOGHDEthvT2rGl1pIR
bzGnH2g/TUsB9K0mtmZ9b8GF7+//KnpBAe2fC70NduYI7kSfi7jrpfPF0ZnQ
hf3tvxibPQ5335Lrh8yC+CjjTC4fZow8HNW97G477uW3b8DeSzlCsSlI9eYs
8InFEFp6ifpD7tmWElINRBBm8FQmZwpeks0ropJ3+DeIPHGfpDJyVsZXj0Nl
b6FNh1iHx0pPlA0LShQ+nU0mqQJXY+b9GkNPb21V3OaH7yb/lGimRen1FP2Y
gUggtM60gKrJOz4pW9214bac7CrDdhcBso5v8uhc05xvRpgc8vqgTWmiZ1+A
QlwRluh1AuQmBaQBCfAO4s+lpUffgJlZk9Sstd4f2wcRHSbTuToc8A4etFQf
vZQzWBxbT89rLwxDmsurWFkSOhmq1vjRsSomt2GcA5MPLqJmtW46V/uHsn6s
o1MLOw/O8Lgno+xdnx/EjSgdAs8Sz1lRDMtimo02tW5tWyKnRjKERevVRQgp
83j7K+zR3JSiTuhycTIrfBsNxzK3cbOICQVjtNwjemDQVkbPK2bBJ26r3ivu
9DlnaUV3I0hRRnisppQ1yy0OerzwEVH0cxoGHakkoMcF5e3vQbOtDPdEhYTe
3Y4vzQnoNfICul/VJragzpzk1mBHjFanW3mFEX4cUN8rLunlFAoMcM6emiXb
MxsjZKCL3B1GYr+bn7XQ9x/URNIzDbZwrgdwevARzBcgohIJlY/TD+0EKjSS
MLo2gM/HKXfH3u5HYrt4piO3a36yFZsehvgrvLB0wIeftTXCPnFAY/StmR8D
ZMrHLlKr0I0DVBd7UM3rSu1X2amL4FNW5BBcDp9/1AAwulUn3J8udnSe61vG
Qr23lj4taXbYHc701xXUxx2/bcJKzUyQgAKej3GthRpzK1FL+eKSAgBz+oLL
cMXZYPKjot/P23nVoUJAJdjZL4sGwxqCAsKxR/kNO/AsGSs/R8hl1k2nLUGn
2/d9fD+LZWWPXeCeTlqtsTr7TDs0Lo6dZyv+TCAjxixIXGCrriBpyLK0sg8U
OeMuGnklh2SMIlaJ7KfVgGP7+jGFrEos3krHDbbMfleT6bcLqz0+16C09Q8k
VxIlI5NY5/vmcE2hwZuVKZfU/xhK+gOekj6uT0KJ3ErSVDpua8dOLzjSzhqN
nS3q8uDW1hgbr5Y/9NGGt/CsGAAxceEZre44B6ExC8HwkahcMW6ggewe9dV5
aMyY4KxkWhlSXiAs0mpqR615gE1Eab53VQ7F1744/f9O9nIkQ/2N60OS1o5G
JpmCz/bo05NVGowBoO1xl/yR9H2HuLWXDtS+Ou6vHuq1g9oO/57NL9C6krC3
c9uXOtd0wUaLhdKxCNv2GXmvKgckrecM1e49IGDqfz27r+KscaqVkpdxkruc
05zlAvZ16qIebO/mO0GLKUuf6sB3FsN+ryHGe07dnoJ/v6nNh9sL7oaMeAfh
ea8JbdmySq0WNV6OJ8uCH8mPoi4oBu1M1PxiNi3ymaZ8gyVQ4orhjN8dqIqV
+QlphKXLqozGWyQwQf/WbkQkI9PXDbIvvGlrRQ22bGz1B0D3KOZkazynojxN
1VW7PzwIsZQ67RN2EvaZ5PfeFGua19lHTdz2zPlRpY9mOdLGRAfG1f+b/LHN
XU+IwFc6PTHdlNQnqteuxxeMDBz7GBVd0C3T5hHsprYWjVISXMYc4ilboh1K
ujRlQbDbaxBKbO6hFyWU18KUUj5nhoXLcfMUJY3mHfBFeAGrwrk0tys3PX4I
gFWAY6lppRLxLjzLWFCgG2twb+6umdBrAO0hBu3+bnYn7IaWRLFIhO2WRL3F
KLX6F3gg+ACeybQIlf36fUOHNLUY9qQGRFa4aQpDIePLzzVI5ue3ox51omed
V+24WxZ4o3UyB4U2WOnYShCgK0qIUgMgL7RtRCToncFt7JyJToiItw0veMDz
ihp7AptEb8G6ytimHY1iOK53S1Cj552h1ZR3edHTqGrJC94N+QkKhxi2ejlX
kNGcb1IfO49KRBbpPphimMnOkFg6jfKAr8Yjt9+ZaaGjr+3U38/huOIIjkdm
W1VaLE/Q/D5Cquu8MHJPAe9Y1E2edvdloFPoxodteJKlxOOWOhZOkqdfq1IH
gOCJxqef1FnaV2FysQ21YAmiVWWslyz7YXmRvey1+TEAAxhUNCTJV9VWaWry
9GwLbRCV1Qgevr4YtPC99XftuG4vfqn/GZWnd1Ca1V+zeLgvW5fvjBQsFL4Q
u49WFUfZ3u3Es2ziCmQ3isUqFmJkQ6NAPXvENI7XOugKfECyQoJSos97jcvJ
pEnw5QEKTZHGezbANhKcFFtVbG6/fAksG04HKLa2wr28BzwJWS0mmBkS50cA
b38CbifcH0j9IyvrH2nlLJQ+QYtnixtNj9hEK279RmWqKjzcuJaXT7OnTEcF
Pkqx/DbT3YZDCKG3ibU5kexS59hP0QvkFVOBZc8kco6J319a149D04jENmW7
jtmMpX2Q6rTdf+tnmlEJUDLqBIBYct4RwxEJ8osWQ7cEk5MbVxqcxC4Kzj0e
xSHK5Dq98RPgE9T4jozopWx3Qqx2hJRzU03jNkT//ew3GcriBJ6+iFExFstW
27JbFk0Oi+eAFhiNVNaW5kxabBTLN6UWsDXvEsnjidHRWQJXgOPMlq+VxWAe
CBtCzoTUgeKP5CNSmzx3GNdPUv3NU2hNzim36xiu1toweqRf1/x6Ynwd8gvI
GfddkVogP6/VCHAJs71FgUnBPPS+mKxj5z7QHhg1hUCEByq5t/mlp2LYFy70
w7h9/GRIvDHjTlTOKmzmOsntwCfU40wTxtTQIvrTwag46w/cUmiAkrX8TAHn
bhLRynFpkooZRisjcTB1JlF8vEFWqWjYmnNEeIx7sUJM7bVxRa1SmwdpToaR
NFRwo4I+Knzuc+q4WuW0c5oFFE/Hmc98aH3qQ1Anw54XCifccLiXuoZnRg4z
eFOy4M2S3Xxcva0VNiF+lvCPUFjm5eFfwK8cktVSCcZgPFqilbi+54SeGbR3
Rqo7nv2q9UbfNA5bKRiec56UWbjTrPK9B+EFQiusN9/jTNdvZEmKIn2WjaEm
l8gDITNSPVobfB//b3TF0/plV0hFJG+nDqMhBlgTbGd7R9cgVdp9ao/9XQ4Y
Cr1uFYC3jAPpTLaKza1VLi5hWFj2vzuaJdcp//igGOfAWB+rofz5QJtxboX4
vzSvzss3qoVDCAUuztFGFoUsxyozVCKwh1h4vtNXcfkmrTXdpxYtfcgYNxDe
lwuIGFvEs+d4CA4UOdbBqu3zBb+ruN1CeoRFLFkbvIwqlgNpIDnd/uewMuIp
Z2LhMM2PJn/wHiCFHULnC2+0fxYenScpdx3RMoZEv9/PyotDtpRmYvb59FMA
TLy8P4CIi96Ugnz6x0dhgBHfGMWN79iJ0wYjCM2zNn7VxKaZjPtxhYzP8/n/
uQkHpqnKhgGuAgIlmieDkh0ZvR9nE9mbfeiXS5OLZwdR5BQBZPoby6Hp6tc8
CLec0VQV6JnamVB5WtIDsdjWX890cTwO0oT7HA6KLnFc5gjQ33/RkRGLfgIJ
gs1dYqHHR7UwfXOaFgUQQTQDLeVWtYIllpZoNSWRmYgNNwsSGgE0AJfFpmik
lh4oYQIU5bJ6P4bVw6haM8HYhaY9GDVT6/W0MyhnP8VbahbgATTrpSSQTlv7
irqERF/KBP+oPqgsAGmICI8XohTjHE1EJQv3v6v11toKpoZ4xfTCYRBcVjPB
YhfsbOoVsSce+gGxKuDSYuN/k+nubn14oZzka3Wex58BkHFrHHsGUynMHGgv
ziY8FDLCDLvjqU5AW6dSFObdup6pzHwRDnA4+nsI2LZaaxYY12ilwSLYXodu
7uOx+CA7XXhuzNpaUPaNkhEbX+Z1rCxEW+5xgwcG4b+qlzMKzs1JDMh893tY
6PkZE8pTmZfJRkQVa+6VaK8s/MmmXUr/Jm0rZv24XT8u0moeyabTX9Pqrkyx
7V5WZNz8d3zrJZtaRSp0O4Gi2eTFfmhjPn8c1ZSz4VnS1jICRWs8YGeNBi5K
nPbSBA8Xfl5bKUl5DlRmFrgb0dmrTgCxpy0Mm/m//IAzGvUkxTGMWKogkWeX
MgsAlNCS6AZnSLDE9m5suXaxXeNnYqPkgkAiJczindIUFZ4SKxtCuTXecx8J
n/M08AufoloOPEY81qzGDlF6Du+N7/BQqZjHT0fr0wKVkiFy9EfpRPz0qxQC
XesxTbs8kIamRXJEBV9/pH+x53gsfmCCQ8a4XizvXd5eym/XDPghrAqUEQnX
FtlKGUG9plxTPAbB4P+gJcO4Fo3Zt4d49T0XaVDRdOYdfbO2A97Pd6YzHJOE
+iXeYPcQJ3tepCLri+axX2COwa23XhiH230TTy8ghgrcObowT3HzYWjqmLKJ
/ce4Y+88/szOOgZFsI2nkedm2vRg4V7iZZmeGnodFt0uW6rMFmiuWusYVcQq
+VgEsbPJjXnEv0mw0tRzSOP8xTrCG7iz8ReERPFmP+Ua196PrXwYmx6LycMh
b4+zt/N82cp0mo4qwtAstOfzIY6HMWK36qxRtYICvXw4PdTIVl6ULdBVFmCc
h0YkF4LnSjhz3XbL2tfeQDm0U7zcTH6WyqsLu6Zcy9S0QeJWQvzu/VUxbyd1
UybC6cje6pomvyuuC7LOocOpyN7H28ezZ9jh6DD/fRO/aNQzA8+jAqIWrqCG
bqXYFA87ylh56+JcZj2IIElojOeXj5imMNnyYAeXYSE7+vRs4C5l6D/BpTZt
0DKSqjJMoQ30Z4kYCBwFfi8lEAQ0+9EgMYc2Vy9IdHQZTAN56k+YCXu6VTYP
FmUO6AaRRHwZzhg2j1SzDTC58orn+El9M8XAXn6zeNoU2RUld2pnywcn1SPa
k4QElIWGJaCx8hfng5q6DE64iGx6K24UgbOt5f4b6tYL5xu8dhl4yhpiDg3n
SZzVqmtkiUPTx9bfBfE7fl12mB2A6zy20e13sYeYVKWLgiR8FmtQYPcowSUq
2IBPrV4fG/oXO4VpxMwcOgiECeGfZIi+ygLZFJVH97Gfu2Hi9pgSnGXGIJy6
eA3TjQ6P+9wJU1wAVIhQuuYn7dYF5cNoZurIri+wl4q1akVvdJZy4OGaqLw7
ILBTw9H2QFzCfrdaWKbM5UzP+kI2dBAvPruYtHhIc+A0kGMNLebogcfOXrT5
8WtWuNkCByRuFWvJMiqPd83CZfE7XZmyumNuhHIAJkurFRQSNP7AU2lhS5yU
LGKb7thL2Xl2AQAW0R/aJ6CebkoQa+inaYSsAGc6vxVxcMEBhYFcjKnaNuho
m93BQL0ozswfdEBK4UNsP0A8rEva34NCmJy7lCt0EpcZs5u+JMw5ajloUGtO
tob60rK4MfWD9ugumApD00OXr8tn5Luggazw3firYJdYBqoGbNn34I5SMGX8
z3FNpZKYg/c0KhdJwUMksvy9TYfGGrvi+t7+gyDV4ogmXFORsrAJHC6irUcO
g782wFVHb6nHWZHo4JLMmotgU2jl9zqfSruzF42+jcJTwVM3b6OW1Ic8L87F
CKswsZWUsyfZYHXJxof97BAtZeLrO7FXYREgI4Vh+T3PtIbd6fHMqqnPIIOs
XRaLehtb3RiUC/fpP9BgH5BMRXjH4+xPxgzvKYb77Rl6QfAsTokiDr1+2ikB
KOerD7OLPHxMSaRhdQPBxkKk+6LBh8pNLI1EsuaHwmEtR8ECqydopF5mv2RA
ONBItwgoWXYvGyzCRQ/B9dK9UC5oVHiihmteI7t8m4t95OKRre38ZlqMWgvo
8Qjm1ZYNmzVy3SdYF928DQ4LatrJOqKlYXz+9t+DfCmMjhHD6lZf6l27Pxzq
8MfX9ZpFruu6SjsrfUfAX0NbvDz06O5l9qM7PfTZ7zi5uh546Ar0eHYEx0te
QfPjvsByFyzqD4ZHgqheE/l+tfAOE1pmuEAbVfIsSAoX8ub+4dXhe4b5/Upm
Fdj9k7VdTExKv1gtKDH2/oF+6S63P5Ovnl6eD2hc2GNMfCfXjv+xynvZaioa
znq7Iw/wYj0KlSMcOKp1iu3Cf/ogrvA4AltxKjcqn3z42eguTuEnge86TfLx
gb9CbxdcAPBh+qHbFJDKHtsyEmwN97JFwIEjCZNpp1dqYEKwQnTfVC52rxXK
8pmb3u6NUhsGmZx8aoadZPAy2rgO0QJvMiQ4cprhu1GfXosBmwtR8ftKQ+pn
FsKiJHurbS++J2fN3hNXR4Uy4L8VlNftob0pG7agYWAeXYe5fSXoKbvxT4K1
xA1hdfB0Pv+4fgpA3Zm+rQFU54rpyqHp8xjPvg3ioAx/sZJbtWAKk5yv6Ibk
Gcd3OaLT0AoatfvvPMVxpdciACMR1iZJS69W8bzbVCFBTtO9MTUpwCvkG9IP
MFCinpXcVBr802GY7anx996RFDkojMOa9cAcd3p6o4YkMugrFqp7kJu5wQuJ
s62Q9wLmShb8njtJAj5UdoeKoH9LWiq/m4Z+8e9PjAjbkl9sOUzC5MKF4I+a
ZpBLSsfwQs1jnB9LjUTo2IAIWLuw3c4Jop3C0xH64ELJxr7IBQe0G3LakOP0
rdYEm4jbImMvxxiCnEp5m6dKFh6hsTzZGgAyyXyAdMWxo6igDsAzp52Myqa+
WDlEfDrx73FFwmBWOeET+OcObNCjy5S9JGBwXvB3HZJjdgyF8+GcVDMdJvrN
XHtOrnhpiiSrH8ws+w4cepolk5pMh+xijBIN+KKcBOgL44pZua+hppODNNet
GfwFoQwoFA4SyGiuh5xFyrpzyw9PGtb6qczT5/2g2zZ4kYrHWeBjMCOdIhhd
CnkvkI5CVnkv3XAM2pPFYKyXHfLG6hVLKgCGH0/CZjreNPfUj/pJbNmUZ2oz
vQbcRipGu3Zx/xehQqbUijSNtsyxlnFUhjyoXf5LKEKKEbgLr8bPEdLCBrH3
5JKM61XfVLWrh8O7fq6rU7LTagF/SvkPrl55WFLR2SORBLqPgmvnCL2ma4+E
R/GeAuATxB+p0Inm9UkKaYHsZ1q7LyBMmeIUE69v1+gGYHwCUeOVOYv6qKyY
R0BmXNXVQHc8fgDq12DweOTVifwUtRdj9ODO41Ssv3hbWxHR+7j+vl39zH8A
Jc7+BqfUZLbVX11OGPftWJDecGgAWgbH6V+eMQUgvL9SsR7lWl0Q8zmrtIQl
lRXAei4n33ibZBEViBS7+qAYhI8B5w7VgwmXUBAC7171Mm+QttmtH+tcHPS1
0uZZ7ObABnu7Fbwp/y7AwBD/u0j3V74fUNlQ4UhQVXvsy+zwDl7AsMigFJS3
w7WXHprlSR094HbpCtiyB2SyzD81/FXjpfiiRsgT2LKdLhN/LVqbL5a+Evs3
RzSEXr3PAi/DoF+s2gAMt7nxzpaBSu/f8UYgf2ztjOT7vphfgo6ERD5k0njF
0xTsbz+r2aqIMEYdjL8WtSpJVHyJpovBS06Sr2IP+kRCYJWSSi48fKBfHski
n1xZbrY5mAzw9/7w3+wKyLFvB2kpR+reyR+gqGDUUL2aq4HO2ni1MqNo9KOr
8CK03cJCLzsbewvtmWydvbdyxJEy6Du1O4y6TxXCSagG2l9qFvbur6BeKUt3
SFVyzL7KqajYaWvBIgSKYdIOPOfLLQ3XW5PnHJoFyQT7dYVapMyTM2CLM0gR
RgP9+zATUuq/Wrp4ZvP/OMaGlquUHo3GgPib1qF2T9Za3AZFFUOUJ15vebgX
kGRZqlPnQTsyzluXuxZHcisbMllCIKIUtQI386FGHcmc2A0B+QAkvdy07hQD
8xAFcoUCK3+ly3yN0COsZnU6ZY8Esq+LrUaylgFyUrUCZ2W0nhDd8om9BulK
FqE2gF/brW0EuhUCuTmEOe/ki+dmmZDxuUxlUzMU3WmlI/lHx5DX2vpv3vt/
SRZL2q4WuVVb0sdWeTz0pAnji4ZPYtxnfZ2uHEtWt9gxabT88vh/+I4Z9ITw
F0//Gen1hk+ec4hjTHIFl8Drgwwu93zcLDtWD9rcGNAOTLafaYp7JGGWIczU
pbynHk+uGPU+oC4DmCo3S/QMPYjDRiUKmVaY7yWDQDWqr4qyLjlhDqv3sD9l
pQD5SYKdhNQMFCrthhP405wp3DOX1Uiaa4vGOszenFEL/eYaLdmbMFyLtGoO
F41BOyVi4CYHOFyjycRuNL4KA22k5EolwaAIMXUyw+Tx8HbK+73q5SbRiwjY
/4Lr0eP27DdGzVzyDpgt+aSn8Qgrg0yQdzXM+vqWo6z6Ek2uP7DcQ3VgJhqa
L25h/hU06LTRwhHiuv36NUAjYOWStdqgAa8PRXNUY0lzRutyc2RsmMOUedr8
N9lfWlliK/QYaMWVdrcXdc55f9DxzBXnDaUY+45vd5tB+bjgJzLbCSAPCODD
AC6N0kps5gnNeqQHNVy8QEOWscimMpX9wCB/T9e0Kfkt9x1Uvb7M/cTXWPzo
aKw+RmHrJ2Yz5Q8k/NAYFyjtjbM/aluhMjOTCZC4T0orNGktwhSxDPm42fRc
stR99uWF1AU4R7T9uTL7MofPKGokMp1gMmxrrraJGPNoayTe4V0oXWItsvUH
g6rnzKjH4paVzRDCdwEYiyIUp5mkndAaqu/NIlPhoNvQLPCemdZdhBBHqv9H
A2/0qITZMUyQ10suqyEigM2FA26EPQdGmjxda5As1noyumqTnOpyBJEs+yn0
otFwAtx/SBXBO8zYw+vC4Ud26aJZ0tEGnjWnpqs05mJZ4FU+FSpd+wca9waV
wqrzWjl9HVu9qSeZ085Wf+BzzcXUKDjtndalhwO/AXWKuldUOrQObjY+u+5y
VaAeEXvZJ3XHl01cDSo8/XXctZvqvV2vtWnt1pUKT2qib2IwZu84D+aKKJrs
I/3aqs8A8HTVcEsb9bI/kjX8uT1IUsn+6LpxjArQSQX282H+eo8nCFmgn/nO
vvhykszJ9bcVQ3ScS0M8k5KikefWQdRBlKIZdmMKNu/PLjhRO2Tv0+Jcb27Y
lQkj10WqBFx1oSo0rJGaoobzbf7fCK8ovNj4amY8I8YMsIxVAVShdTWQH5Pv
8yHEhWmfOcY6Rmdrc/xQJavGAtkCRvtueObnvfAZ8owsPfyEH6MzIUL7O6ru
9105wFzg0IvUMksrnYEjnwyyIfeQkjBBTtuuc65weeYjGjaVwhlpxmfZa0LA
WlsjgOIbPxJqj7ZwnM//B9gKiL9wxtQIS5neV8/vc/5Xss/JXd9/7Ysq4jKM
DDny+bHmB8nJ64ROumtoK60VZz4z1ZTtah71+TeIbNn5IBldM90yhMK2PnHo
ivzn3e8gzjGaM+/TXGnfOx+MsIHyfSHHO8MU1IK6v1jFIC+liglyjQaYYZ55
ZNIZ5ohKyxMyLxzoDuvueKi1oxupPziVtWhFRbu1dLXKqY9zKVzwBWcNc8XV
PuTnE/F3TixLsiKLsyunEFQ/gl8T3AWFPrO/BSX6ZnbAZIIKBWIAviTLYHNC
B9QNFPqnGkS5ejR4jzIBvpM0PUCvLsSh3Eilt3mwpPGkewtn0vOoczPsInLI
XizKVQdPAiEZHgDPfUrNnzFgOICKBRBIhICL3QI/fAspFDQrejNmtYj474yr
dC9DgFP4XTSJ3jOPme/XcBUEXDJObcxlghlGYP0h15UqNX1Q0RKVFL2Ipk7L
uU0cNF+O33vJDXLwaKIO8MGHlt0nkZ+vJ6af1zJVtxvXqQVhYoKKptWiFK75
vWLsaE3e6VwZuvfLtCU+x3mDbZLG4H2VyrwEw0riR14XU3beikZA7J2Zvgxi
6DHd2sPB8GKRjh4WDWCxgwQv5cM1eYPynPhDZuenfxHxqhxT07xQ5kCdYoUo
NTsdFFdrraGR9MclvbTkgQqyD/PaSEO70I9SahQ7RVbGj7JK8xkvCkJNnFRj
dc3884vBD8+Ok4ZsRg+bB3kXFeg600gfkMDpqm3IbMbtfxsDPrnibXc6yiun
Umx2/m5jYAfav4WttlvV4ppT2NM0Tqk1M33VmoP8+z3Im1rIl3HgscBuIzkr
lDXuYwVsytVZUDC43z3GKd+bD3dB81VO6AoOLEG1pvGQuKzM6K9rpx6XplP1
JyU2Fl/cO6BZEQMSdQ7h87OYffRqe1cqKpUgcdyqcPNoFX9gds/2XBre2Gr2
VWvQKPxyu4Xlsxaa8FUBqd0+tH6SSF2UDGGIhpNl+OfE6dGI9RDwbzbkOq5F
VvOr/G7DSBnGkdvu/W6qy9xraOhT3zVXt0BeR8VVrFHt2FbLXGxDGx71xzie
WDQ4IHkadjTnzyecnkDuqfGdxjqFuzVzhb+YdhkYeLnBdKBdQs1Di0kHW3ZL
+FZ1v8yEVuuPjl9GnhwGS2Cwz6LgxFwcR+xUDNtZpIusJoVCdEuECZqPhkNQ
m1dUBNVXVrAXPkf/l/8pNT1k8e49MvH4GEqzcB4P3oIGFzLhhfS/vj1C+IxB
D8ogaTGylL9Be4yZK63yX8jIeSHW5vggQ6mEevpoOsJ4WvuPpYFr6GixQCbr
NoK3x/kSSeUe2qiHGuOvoedcv6gz0I6JXBw5aol4hKFnhpBxfxO90a1w6gp5
IDaIuzek/FllJ8WLKZ7itEvMhmQ4CFAMC/5ReR72jA2LVePp9FcU3wqz7LVE
ASaaC4He4DdGf/YKNx3D5rcvhURy5tXk7mHlV9HPWLEd+tt845g963KriCQ0
bNa5dZ5axht9uglOPz9BhrWBDvmBf59VKnXM7JER/wxmClBBKnAyEovCGedN
XoachfBgJQB9ben4LJwucMCrKw0YC4tuYYkzPGtnjXY8IKEkmUOTwkJDqlZ5
1Ya4NKufFSSQNWS05eY8Ov6rLaVg8gethBrzqi3gTGSdY8utXAyycrS4m0Jg
OfUa1u/CVyemHBGPvQrS5Izk+2jvXZhPvxFI/2b/3qz7ttNs0c8nuZ/fErSK
eMeFUQEEvX7G3JJZyBeS0194ohxx4DjwHxGbttQ+nVjHLeN8OTjZnFjbSyX6
un6zEzKWrSHKZiSNUAfGtvqpQcepanHMKxH4XIxTB2rGDiPOtQgXryeR6VlM
ZsTdZpAT81pCx8SOVLZ7/ZhQRyPBT7uQnFXZxzlR7Cirir9edA7NjYqPgKCM
hYnFZTYWqU6QjFktPF3/L1e0ivSdsF4XqHJ5K+NH33TQQvO8UyoByRFHs2yP
JpnGuwzMsnUCqW1tYsQikmEOcHUgOCaQ5290ke3Hd2FBYviEvGDytakIT4+0
zf1zLChKWMA05G4QZlfo6bEMX2t/KRG+SbsCbs/Oyd3Gqar+egsTSVaMCteI
VJ/ku55zRq38uiFtjwtcrPqxvt2UPMf7eYpg2+RKmN6XLlJfbsGG7KGsKvpS
MJ1//GldtjE92Qb83KkifQ6EjAPZMXG5ANYGrmxJ6/cuum+Ml8T0u5Nef+O/
CiHj5HTfzmEQtGKPb6myxNJYXTCJgMWU7f5DK+FpJq35nxyjrpbQoO/kGezz
XQxHt+5Nw1/5i6B+Sk9GHskXCB1QUXa73iHXylQ68XxWAkdz7TvjxSoU3jjv
zsiGbZJ9X3Hfj9sqg6vNTbfwje1dgw5q2PE3KIGZc6u87xEy0/BaoYh+TQpJ
5/Rin0gCUvoV39y3YwDti+36IqryRexhLDH/ZuKy1TiQmHyKHaYKAGZ7f0N5
Kt5D2FbdCdx7ABVDTkKpeZtvtK7gl+wtlBQrI7hIkUiYF64xAuo5T0jwPvNg
zek1ttRAVdtCOOoFB4LCX7co+RTvDHE/v0p33MEyaNXC1RRvcOiNrYkiFFhh
WWNX8VfyYkwJjq3JGWE4NL/2Hi/3fC2XoQLD8Wl8vCAIf0ZyTkGBqMhKmyls
PXpjGMLTYNTjOir5k/fEU9A+T/fdDRsIxE0GEmzLDy7fO4eVRBEe6DaM3ib7
D31J3E+zoD3i5cdoI8w24W7cWK8xajPHjDsLT666T2y4xNeHidJl9JeEpgYL
uJgHIzHJgCrNm6MwQS4Yt3FIyb5XSHGpmjBNrg1zD1nzCF1Idbwuh1Aua7Lm
/c4C7A8vQ19aat/KnYdASgjIDc4+CCX3inAXKbIradUbnOm0uFA52xSynhL6
I88UYxiGbfh2hkNsb/+8PMAK+2lK6FFyj9M4E2fOkg2EOoJnDx35m9kfZvBs
1psUTr6ooGye6ToIVlDeGM6YxoA+NdiM/+Stb0BXvONYAmukEUI4pgiu5eMn
idFfqbOr+jVrSJl95KDtL0MVP5nx3DndmR+rbmp470TNn7IB9UCkCDGiZiO7
B4sfrA2pAVVepgFsmq5UKDFa899GUzJahutkMVzJjZ6Y5OrJdEApHWc0HHRJ
tgSI2aUFt+XDLpIaCeYcC401/lEuNP83MLNO2VFGdm1Z6e2M1YdJGMAEbK8f
pHUMvoix/qwuzd3Npc/4p71VNUJkoJ1t3bLysBDR8h+v6cAB98PRtor3TAXl
AaEYAsgcF2yzITxvw7jMIVDWs63aejMAMXdO9vCaEEiAlXCnTafTQODWdrwO
tzEzCypZbFSrE96dLbMhsbKa4W/HeRQuyiPYZsO/Z/S9Q/NJFvC4vQQ9k82c
aacgacexUn4EY9wycXdMhhhkZPT14hPrjmtotLzg4yysQWLyX81l9cQjsIcV
shoBgyWj+lifYYl6OWxKr0XoJRTtKF6iRT5k39rj/sEFpiQFrLJKiwAuczxc
04Mkdo8hB5vI92X/967vRe+x3dFQOhVECUcclsbHgJEcOUDwY+lS4LQcMSUw
CqbDu8Fq9K3+s+/7pmCLzSMfQk9e30iBMNmYDTqt5nV82J+G43uLxJekBc3t
gxt8Po0+vv5XgifawEUuBVBXate3as/ekGYWUyTn64Sp7+4WA57WpG0zZxzY
melVOIRzEN07QQTp82AKJgjbxpww2EYorx9YqWuA1whMbxr7VQeqqgYexfzj
X8bqzg9Y+bxdHq7vw0Ovd4PycFrtL/xAWGpYHnttgWM75P2DTo/cMTv1VOIv
LNXnUf70QCWbyV4gKG8h3QZN4rif93bQV5+mM8bHmnTuyiwUb0Jxer+fr3gD
0m1wT6uNzij0c6ki3/4Qr4K0kpgeJn9VwTq6fdp+w+oftzCcjMHBw2ksYMBO
4wbMm9ldsjenzQNqvExuYarGS3bdCy2fTtcRPfiLePKCYNlCuHilNR/Vo3GV
ld7ogUSQG5pkDgfpihdJtLUTKxabTUhuL9o6NaplpVDOMFBoZf72ADI13paL
YYisosiupQUjqC2PGvhF+j4pX5YbzhIL0K7KE9aW5YzXnp2o9+QLJGUft8ha
ey2HTivo0Ya5uzTp8p1q52J/4poOkZuRdw==

`pragma protect end_protected
