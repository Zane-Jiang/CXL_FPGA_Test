// intel_rtile_cxl_top_cxltyp3_ed.v

// Generated using ACDS version 22.4 94

`timescale 1 ps / 1 ps
module intel_rtile_cxl_top_cxltyp3_ed (
		input  wire         refclk4,                           //             refclk.clk
		input  wire         refclk0,                           //            refclk0.clk
		input  wire         refclk1,                           //            refclk1.clk
		input  wire         resetn,                            //             resetn.reset_n
		input  wire         nInit_done,                        //         ninit_done.ninit_done
		output wire         sip_warm_rstn_o,                   //      sip_warm_rstn.reset_n
		output wire         cxl_warm_rst_n,                    //          warm_rstn.reset_n
		output wire         cxl_cold_rst_n,                    //          cold_rstn.reset_n
		input  wire [15:0]  cxl_rx_n,                          //                cxl.rx_n
		input  wire [15:0]  cxl_rx_p,                          //                   .rx_p
		output wire [15:0]  cxl_tx_n,                          //                   .tx_n
		output wire [15:0]  cxl_tx_p,                          //                   .tx_p
		input  wire [35:0]  hdm_size_256mb,                    //            memsize.hdm_size
		input  wire [63:0]  mc2ip_memsize,                     //                   .mem_size
		output wire         ip2hdm_clk,                        //         ip2hdm_clk.clk
		output wire         ip2hdm_reset_n,                    //     ip2hdm_reset_n.reset
		input  wire [4:0]   mc2ip_0_sr_status,                 //            mc2ip_0.sr_status
		input  wire         mc2ip_0_rspfifo_full,              //                   .rspfifo_full
		input  wire         mc2ip_0_rspfifo_empty,             //                   .rspfifo_empty
		input  wire [5:0]   mc2ip_0_rspfifo_fill_level,        //                   .rspfifo_fill_level
		input  wire         mc2ip_0_reqfifo_full,              //                   .reqfifo_full
		input  wire         mc2ip_0_reqfifo_empty,             //                   .reqfifo_empty
		input  wire [5:0]   mc2ip_0_reqfifo_fill_level,        //                   .reqfifo_fill_level
		input  wire         hdm2ip_avmm0_ready,                //       hdm2ip_avmm0.ready
		input  wire         hdm2ip_avmm0_cxlmem_ready,         //                   .cxlmem_ready
		input  wire [511:0] hdm2ip_avmm0_readdata,             //                   .readdata
		input  wire [13:0]  hdm2ip_avmm0_rsp_mdata,            //                   .rsp_mdata
		input  wire         hdm2ip_avmm0_read_poison,          //                   .read_poison
		input  wire         hdm2ip_avmm0_readdatavalid,        //                   .readdatavalid
		input  wire [7:0]   hdm2ip_avmm0_ecc_err_corrected,    //                   .ecc_err_corrected
		input  wire [7:0]   hdm2ip_avmm0_ecc_err_detected,     //                   .ecc_err_detected
		input  wire [7:0]   hdm2ip_avmm0_ecc_err_fatal,        //                   .ecc_err_fatal
		input  wire [7:0]   hdm2ip_avmm0_ecc_err_syn_e,        //                   .ecc_err_syn_e
		input  wire         hdm2ip_avmm0_ecc_err_valid,        //                   .ecc_err_valid
		output wire         ip2hdm_avmm0_read,                 //       ip2hdm_avmm0.read
		output wire         ip2hdm_avmm0_write,                //                   .write
		output wire         ip2hdm_avmm0_write_poison,         //                   .write_poison
		output wire         ip2hdm_avmm0_write_ras_sbe,        //                   .write_ras_sbe
		output wire         ip2hdm_avmm0_write_ras_dbe,        //                   .write_ras_dbe
		output wire [511:0] ip2hdm_avmm0_writedata,            //                   .writedata
		output wire [63:0]  ip2hdm_avmm0_byteenable,           //                   .byteenable
		output wire [45:0]  ip2hdm_avmm0_address,              //                   .address
		output wire [13:0]  ip2hdm_avmm0_req_mdata,            //                   .req_mdata
		input  wire [4:0]   mc2ip_1_sr_status,                 //            mc2ip_1.sr_status
		input  wire         mc2ip_1_rspfifo_full,              //                   .rspfifo_full
		input  wire         mc2ip_1_rspfifo_empty,             //                   .rspfifo_empty
		input  wire [5:0]   mc2ip_1_rspfifo_fill_level,        //                   .rspfifo_fill_level
		input  wire         mc2ip_1_reqfifo_full,              //                   .reqfifo_full
		input  wire         mc2ip_1_reqfifo_empty,             //                   .reqfifo_empty
		input  wire [5:0]   mc2ip_1_reqfifo_fill_level,        //                   .reqfifo_fill_level
		input  wire         hdm2ip_avmm1_ready,                //       hdm2ip_avmm1.ready
		input  wire         hdm2ip_avmm1_cxlmem_ready,         //                   .cxlmem_ready
		input  wire [511:0] hdm2ip_avmm1_readdata,             //                   .readdata
		input  wire [13:0]  hdm2ip_avmm1_rsp_mdata,            //                   .rsp_mdata
		input  wire         hdm2ip_avmm1_read_poison,          //                   .read_poison
		input  wire         hdm2ip_avmm1_readdatavalid,        //                   .readdatavalid
		input  wire [7:0]   hdm2ip_avmm1_ecc_err_corrected,    //                   .ecc_err_corrected
		input  wire [7:0]   hdm2ip_avmm1_ecc_err_detected,     //                   .ecc_err_detected
		input  wire [7:0]   hdm2ip_avmm1_ecc_err_fatal,        //                   .ecc_err_fatal
		input  wire [7:0]   hdm2ip_avmm1_ecc_err_syn_e,        //                   .ecc_err_syn_e
		input  wire         hdm2ip_avmm1_ecc_err_valid,        //                   .ecc_err_valid
		output wire         ip2hdm_avmm1_read,                 //       ip2hdm_avmm1.read
		output wire         ip2hdm_avmm1_write,                //                   .write
		output wire         ip2hdm_avmm1_write_poison,         //                   .write_poison
		output wire         ip2hdm_avmm1_write_ras_sbe,        //                   .write_ras_sbe
		output wire         ip2hdm_avmm1_write_ras_dbe,        //                   .write_ras_dbe
		output wire [511:0] ip2hdm_avmm1_writedata,            //                   .writedata
		output wire [63:0]  ip2hdm_avmm1_byteenable,           //                   .byteenable
		output wire [45:0]  ip2hdm_avmm1_address,              //                   .address
		output wire [13:0]  ip2hdm_avmm1_req_mdata,            //                   .req_mdata
		output wire         ip2csr_avmm_clk,                   //             ip2csr.clock
		output wire         ip2csr_avmm_rstn,                  //                   .reset_n
		input  wire         csr2ip_avmm_waitrequest,           //                   .waitrequest
		input  wire [31:0]  csr2ip_avmm_readdata,              //                   .readdata
		input  wire         csr2ip_avmm_readdatavalid,         //                   .readdatavalid
		output wire [31:0]  ip2csr_avmm_writedata,             //                   .writedata
		output wire [21:0]  ip2csr_avmm_address,               //                   .address
		output wire         ip2csr_avmm_write,                 //                   .write
		output wire         ip2csr_avmm_read,                  //                   .read
		output wire [3:0]   ip2csr_avmm_byteenable,            //                   .byteenable
		output wire         ip2uio_tx_ready,                   //         usr_tx_st0.ready
		input  wire         uio2ip_tx_st0_dvalid,              //                   .dvalid
		input  wire         uio2ip_tx_st0_sop,                 //                   .sop
		input  wire         uio2ip_tx_st0_eop,                 //                   .eop
		input  wire         uio2ip_tx_st0_passthrough,         //                   .passthrough
		input  wire [255:0] uio2ip_tx_st0_data,                //                   .data
		input  wire [7:0]   uio2ip_tx_st0_data_parity,         //                   .data_parity
		input  wire [127:0] uio2ip_tx_st0_hdr,                 //                   .hdr
		input  wire [3:0]   uio2ip_tx_st0_hdr_parity,          //                   .hdr_parity
		input  wire         uio2ip_tx_st0_hvalid,              //                   .hvalid
		input  wire [31:0]  uio2ip_tx_st0_prefix,              //                   .prefix
		input  wire [0:0]   uio2ip_tx_st0_prefix_parity,       //                   .prefix_parity
		input  wire [11:0]  uio2ip_tx_st0_RSSAI_prefix,        //                   .RSSAI_prefix
		input  wire         uio2ip_tx_st0_RSSAI_prefix_parity, //                   .RSSAI_prefix_parity
		input  wire [1:0]   uio2ip_tx_st0_pvalid,              //                   .pvalid
		input  wire         uio2ip_tx_st0_vfactive,            //                   .vfactive
		input  wire [10:0]  uio2ip_tx_st0_vfnum,               //                   .vfnum
		input  wire [2:0]   uio2ip_tx_st0_pfnum,               //                   .pfnum
		input  wire [0:0]   uio2ip_tx_st0_chnum,               //                   .chnum
		input  wire [2:0]   uio2ip_tx_st0_empty,               //                   .empty
		input  wire         uio2ip_tx_st0_misc_parity,         //                   .misc_parity
		input  wire         uio2ip_tx_st1_dvalid,              //         usr_tx_st1.dvalid
		input  wire         uio2ip_tx_st1_sop,                 //                   .sop
		input  wire         uio2ip_tx_st1_eop,                 //                   .eop
		input  wire         uio2ip_tx_st1_passthrough,         //                   .passthrough
		input  wire [255:0] uio2ip_tx_st1_data,                //                   .data
		input  wire [7:0]   uio2ip_tx_st1_data_parity,         //                   .data_parity
		input  wire [127:0] uio2ip_tx_st1_hdr,                 //                   .hdr
		input  wire [3:0]   uio2ip_tx_st1_hdr_parity,          //                   .hdr_parity
		input  wire         uio2ip_tx_st1_hvalid,              //                   .hvalid
		input  wire [31:0]  uio2ip_tx_st1_prefix,              //                   .prefix
		input  wire [0:0]   uio2ip_tx_st1_prefix_parity,       //                   .prefix_parity
		input  wire [11:0]  uio2ip_tx_st1_RSSAI_prefix,        //                   .RSSAI_prefix
		input  wire         uio2ip_tx_st1_RSSAI_prefix_parity, //                   .RSSAI_prefix_parity
		input  wire [1:0]   uio2ip_tx_st1_pvalid,              //                   .pvalid
		input  wire         uio2ip_tx_st1_vfactive,            //                   .vfactive
		input  wire [10:0]  uio2ip_tx_st1_vfnum,               //                   .vfnum
		input  wire [2:0]   uio2ip_tx_st1_pfnum,               //                   .pfnum
		input  wire [0:0]   uio2ip_tx_st1_chnum,               //                   .chnum
		input  wire [2:0]   uio2ip_tx_st1_empty,               //                   .empty
		input  wire         uio2ip_tx_st1_misc_parity,         //                   .misc_parity
		input  wire         uio2ip_tx_st2_dvalid,              //         usr_tx_st2.dvalid
		input  wire         uio2ip_tx_st2_sop,                 //                   .sop
		input  wire         uio2ip_tx_st2_eop,                 //                   .eop
		input  wire         uio2ip_tx_st2_passthrough,         //                   .passthrough
		input  wire [255:0] uio2ip_tx_st2_data,                //                   .data
		input  wire [7:0]   uio2ip_tx_st2_data_parity,         //                   .data_parity
		input  wire [127:0] uio2ip_tx_st2_hdr,                 //                   .hdr
		input  wire [3:0]   uio2ip_tx_st2_hdr_parity,          //                   .hdr_parity
		input  wire         uio2ip_tx_st2_hvalid,              //                   .hvalid
		input  wire [31:0]  uio2ip_tx_st2_prefix,              //                   .prefix
		input  wire [0:0]   uio2ip_tx_st2_prefix_parity,       //                   .prefix_parity
		input  wire [11:0]  uio2ip_tx_st2_RSSAI_prefix,        //                   .RSSAI_prefix
		input  wire         uio2ip_tx_st2_RSSAI_prefix_parity, //                   .RSSAI_prefix_parity
		input  wire [1:0]   uio2ip_tx_st2_pvalid,              //                   .pvalid
		input  wire         uio2ip_tx_st2_vfactive,            //                   .vfactive
		input  wire [10:0]  uio2ip_tx_st2_vfnum,               //                   .vfnum
		input  wire [2:0]   uio2ip_tx_st2_pfnum,               //                   .pfnum
		input  wire [0:0]   uio2ip_tx_st2_chnum,               //                   .chnum
		input  wire [2:0]   uio2ip_tx_st2_empty,               //                   .empty
		input  wire         uio2ip_tx_st2_misc_parity,         //                   .misc_parity
		input  wire         uio2ip_tx_st3_dvalid,              //         usr_tx_st3.dvalid
		input  wire         uio2ip_tx_st3_sop,                 //                   .sop
		input  wire         uio2ip_tx_st3_eop,                 //                   .eop
		input  wire         uio2ip_tx_st3_passthrough,         //                   .passthrough
		input  wire [255:0] uio2ip_tx_st3_data,                //                   .data
		input  wire [7:0]   uio2ip_tx_st3_data_parity,         //                   .data_parity
		input  wire [127:0] uio2ip_tx_st3_hdr,                 //                   .hdr
		input  wire [3:0]   uio2ip_tx_st3_hdr_parity,          //                   .hdr_parity
		input  wire         uio2ip_tx_st3_hvalid,              //                   .hvalid
		input  wire [31:0]  uio2ip_tx_st3_prefix,              //                   .prefix
		input  wire [0:0]   uio2ip_tx_st3_prefix_parity,       //                   .prefix_parity
		input  wire [11:0]  uio2ip_tx_st3_RSSAI_prefix,        //                   .RSSAI_prefix
		input  wire         uio2ip_tx_st3_RSSAI_prefix_parity, //                   .RSSAI_prefix_parity
		input  wire [1:0]   uio2ip_tx_st3_pvalid,              //                   .pvalid
		input  wire         uio2ip_tx_st3_vfactive,            //                   .vfactive
		input  wire [10:0]  uio2ip_tx_st3_vfnum,               //                   .vfnum
		input  wire [2:0]   uio2ip_tx_st3_pfnum,               //                   .pfnum
		input  wire [0:0]   uio2ip_tx_st3_chnum,               //                   .chnum
		input  wire [2:0]   uio2ip_tx_st3_empty,               //                   .empty
		input  wire         uio2ip_tx_st3_misc_parity,         //                   .misc_parity
		output wire [2:0]   ip2uio_tx_st_Hcrdt_update,         //          usr_tx_st.Hcrdt_update
		output wire [0:0]   ip2uio_tx_st_Hcrdt_ch,             //                   .Hcrdt_ch
		output wire [5:0]   ip2uio_tx_st_Hcrdt_update_cnt,     //                   .Hcrdt_update_cnt
		output wire [2:0]   ip2uio_tx_st_Hcrdt_init,           //                   .Hcrdt_init
		input  wire [2:0]   uio2ip_tx_st_Hcrdt_init_ack,       //                   .Hcrdt_init_ack
		output wire [2:0]   ip2uio_tx_st_Dcrdt_update,         //                   .Dcrdt_update
		output wire [0:0]   ip2uio_tx_st_Dcrdt_ch,             //                   .Dcrdt_ch
		output wire [11:0]  ip2uio_tx_st_Dcrdt_update_cnt,     //                   .Dcrdt_update_cnt
		output wire [2:0]   ip2uio_tx_st_Dcrdt_init,           //                   .Dcrdt_init
		input  wire [2:0]   uio2ip_tx_st_Dcrdt_init_ack,       //                   .Dcrdt_init_ack
		output wire         ip2uio_rx_st0_dvalid,              //        usr_rx_st_0.dvalid
		output wire         ip2uio_rx_st0_sop,                 //                   .sop
		output wire         ip2uio_rx_st0_eop,                 //                   .eop
		output wire         ip2uio_rx_st0_passthrough,         //                   .passthrough
		output wire [255:0] ip2uio_rx_st0_data,                //                   .data
		output wire [7:0]   ip2uio_rx_st0_data_parity,         //                   .data_parity
		output wire [127:0] ip2uio_rx_st0_hdr,                 //                   .hdr
		output wire [3:0]   ip2uio_rx_st0_hdr_parity,          //                   .hdr_parity
		output wire         ip2uio_rx_st0_hvalid,              //                   .hvalid
		output wire [31:0]  ip2uio_rx_st0_prefix,              //                   .prefix
		output wire [0:0]   ip2uio_rx_st0_prefix_parity,       //                   .prefix_parity
		output wire [11:0]  ip2uio_rx_st0_RSSAI_prefix,        //                   .RSSAI_prefix
		output wire         ip2uio_rx_st0_RSSAI_prefix_parity, //                   .RSSAI_prefix_parity
		output wire [1:0]   ip2uio_rx_st0_pvalid,              //                   .pvalid
		output wire [2:0]   ip2uio_rx_st0_bar,                 //                   .bar
		output wire         ip2uio_rx_st0_vfactive,            //                   .vfactive
		output wire [10:0]  ip2uio_rx_st0_vfnum,               //                   .vfnum
		output wire [2:0]   ip2uio_rx_st0_pfnum,               //                   .pfnum
		output wire [0:0]   ip2uio_rx_st0_chnum,               //                   .chnum
		output wire         ip2uio_rx_st0_misc_parity,         //                   .misc_parity
		output wire [2:0]   ip2uio_rx_st0_empty,               //                   .empty
		output wire         ip2uio_rx_st1_dvalid,              //        usr_rx_st_1.dvalid
		output wire         ip2uio_rx_st1_sop,                 //                   .sop
		output wire         ip2uio_rx_st1_eop,                 //                   .eop
		output wire         ip2uio_rx_st1_passthrough,         //                   .passthrough
		output wire [255:0] ip2uio_rx_st1_data,                //                   .data
		output wire [7:0]   ip2uio_rx_st1_data_parity,         //                   .data_parity
		output wire [127:0] ip2uio_rx_st1_hdr,                 //                   .hdr
		output wire [3:0]   ip2uio_rx_st1_hdr_parity,          //                   .hdr_parity
		output wire         ip2uio_rx_st1_hvalid,              //                   .hvalid
		output wire [31:0]  ip2uio_rx_st1_prefix,              //                   .prefix
		output wire [0:0]   ip2uio_rx_st1_prefix_parity,       //                   .prefix_parity
		output wire [11:0]  ip2uio_rx_st1_RSSAI_prefix,        //                   .RSSAI_prefix
		output wire         ip2uio_rx_st1_RSSAI_prefix_parity, //                   .RSSAI_prefix_parity
		output wire [1:0]   ip2uio_rx_st1_pvalid,              //                   .pvalid
		output wire [2:0]   ip2uio_rx_st1_bar,                 //                   .bar
		output wire         ip2uio_rx_st1_vfactive,            //                   .vfactive
		output wire [10:0]  ip2uio_rx_st1_vfnum,               //                   .vfnum
		output wire [2:0]   ip2uio_rx_st1_pfnum,               //                   .pfnum
		output wire [0:0]   ip2uio_rx_st1_chnum,               //                   .chnum
		output wire         ip2uio_rx_st1_misc_parity,         //                   .misc_parity
		output wire [2:0]   ip2uio_rx_st1_empty,               //                   .empty
		output wire         ip2uio_rx_st2_dvalid,              //        usr_rx_st_2.dvalid
		output wire         ip2uio_rx_st2_sop,                 //                   .sop
		output wire         ip2uio_rx_st2_eop,                 //                   .eop
		output wire         ip2uio_rx_st2_passthrough,         //                   .passthrough
		output wire [255:0] ip2uio_rx_st2_data,                //                   .data
		output wire [7:0]   ip2uio_rx_st2_data_parity,         //                   .data_parity
		output wire [127:0] ip2uio_rx_st2_hdr,                 //                   .hdr
		output wire [3:0]   ip2uio_rx_st2_hdr_parity,          //                   .hdr_parity
		output wire         ip2uio_rx_st2_hvalid,              //                   .hvalid
		output wire [31:0]  ip2uio_rx_st2_prefix,              //                   .prefix
		output wire [0:0]   ip2uio_rx_st2_prefix_parity,       //                   .prefix_parity
		output wire [11:0]  ip2uio_rx_st2_RSSAI_prefix,        //                   .RSSAI_prefix
		output wire         ip2uio_rx_st2_RSSAI_prefix_parity, //                   .RSSAI_prefix_parity
		output wire [1:0]   ip2uio_rx_st2_pvalid,              //                   .pvalid
		output wire [2:0]   ip2uio_rx_st2_bar,                 //                   .bar
		output wire         ip2uio_rx_st2_vfactive,            //                   .vfactive
		output wire [10:0]  ip2uio_rx_st2_vfnum,               //                   .vfnum
		output wire [2:0]   ip2uio_rx_st2_pfnum,               //                   .pfnum
		output wire [0:0]   ip2uio_rx_st2_chnum,               //                   .chnum
		output wire         ip2uio_rx_st2_misc_parity,         //                   .misc_parity
		output wire [2:0]   ip2uio_rx_st2_empty,               //                   .empty
		output wire         ip2uio_rx_st3_dvalid,              //        usr_rx_st_3.dvalid
		output wire         ip2uio_rx_st3_sop,                 //                   .sop
		output wire         ip2uio_rx_st3_eop,                 //                   .eop
		output wire         ip2uio_rx_st3_passthrough,         //                   .passthrough
		output wire [255:0] ip2uio_rx_st3_data,                //                   .data
		output wire [7:0]   ip2uio_rx_st3_data_parity,         //                   .data_parity
		output wire [127:0] ip2uio_rx_st3_hdr,                 //                   .hdr
		output wire [3:0]   ip2uio_rx_st3_hdr_parity,          //                   .hdr_parity
		output wire         ip2uio_rx_st3_hvalid,              //                   .hvalid
		output wire [31:0]  ip2uio_rx_st3_prefix,              //                   .prefix
		output wire [0:0]   ip2uio_rx_st3_prefix_parity,       //                   .prefix_parity
		output wire [11:0]  ip2uio_rx_st3_RSSAI_prefix,        //                   .RSSAI_prefix
		output wire         ip2uio_rx_st3_RSSAI_prefix_parity, //                   .RSSAI_prefix_parity
		output wire [1:0]   ip2uio_rx_st3_pvalid,              //                   .pvalid
		output wire [2:0]   ip2uio_rx_st3_bar,                 //                   .bar
		output wire         ip2uio_rx_st3_vfactive,            //                   .vfactive
		output wire [10:0]  ip2uio_rx_st3_vfnum,               //                   .vfnum
		output wire [2:0]   ip2uio_rx_st3_pfnum,               //                   .pfnum
		output wire [0:0]   ip2uio_rx_st3_chnum,               //                   .chnum
		output wire         ip2uio_rx_st3_misc_parity,         //                   .misc_parity
		output wire [2:0]   ip2uio_rx_st3_empty,               //                   .empty
		input  wire [2:0]   uio2ip_rx_st_Hcrdt_update,         //          usr_rx_st.Hcrdt_update
		input  wire [0:0]   uio2ip_rx_st_Hcrdt_ch,             //                   .Hcrdt_ch
		input  wire [5:0]   uio2ip_rx_st_Hcrdt_update_cnt,     //                   .Hcrdt_update_cnt
		input  wire [2:0]   uio2ip_rx_st_Hcrdt_init,           //                   .Hcrdt_init
		output wire [2:0]   ip2uio_rx_st_Hcrdt_init_ack,       //                   .Hcrdt_init_ack
		input  wire [2:0]   uio2ip_rx_st_Dcrdt_update,         //                   .Dcrdt_update
		input  wire [0:0]   uio2ip_rx_st_Dcrdt_ch,             //                   .Dcrdt_ch
		input  wire [11:0]  uio2ip_rx_st_Dcrdt_update_cnt,     //                   .Dcrdt_update_cnt
		input  wire [2:0]   uio2ip_rx_st_Dcrdt_init,           //                   .Dcrdt_init
		output wire [2:0]   ip2uio_rx_st_Dcrdt_init_ack,       //                   .Dcrdt_init_ack
		output wire [7:0]   ip2uio_bus_number,                 //                uio.usr_bus_number
		output wire [4:0]   ip2uio_device_number,              //                   .usr_device_number
		output wire         pf0_msix_enable,                   // pf0_msix_interface.msix_enable
		output wire         pf0_msix_fn_mask,                  //                   .msix_fn_mask
		output wire         pf1_msix_enable,                   // pf1_msix_interface.msix_enable
		output wire         pf1_msix_fn_mask                   //                   .msix_fn_mask
	);

	cxl_ip_top #(
		.ADME_ENABLE         (1),
		.PF0_MSIX_CAP_EN     (0),
		.PF0_MSIX_TABLE_SIZE (0),
		.PF0_MSIX_TABLE_MAO  (0),
		.PF0_MSIX_TABLE_BIR  (0),
		.PF0_MSIX_PBA_MAO    (0),
		.PF0_MSIX_PBA_BIR    (0),
		.PF1_MSIX_CAP_EN     (0),
		.PF1_MSIX_TABLE_SIZE (0),
		.PF1_MSIX_TABLE_MAO  (0),
		.PF1_MSIX_TABLE_BIR  (0),
		.PF1_MSIX_PBA_MAO    (0),
		.PF1_MSIX_PBA_BIR    (0)
	) intel_rtile_cxl_top_0 (
		.refclk4                           (refclk4),                           //   input,    width = 1,             refclk.clk
		.refclk0                           (refclk0),                           //   input,    width = 1,            refclk0.clk
		.refclk1                           (refclk1),                           //   input,    width = 1,            refclk1.clk
		.resetn                            (resetn),                            //   input,    width = 1,             resetn.reset_n
		.nInit_done                        (nInit_done),                        //   input,    width = 1,         ninit_done.ninit_done
		.sip_warm_rstn_o                   (sip_warm_rstn_o),                   //  output,    width = 1,      sip_warm_rstn.reset_n
		.cxl_warm_rst_n                    (cxl_warm_rst_n),                    //  output,    width = 1,          warm_rstn.reset_n
		.cxl_cold_rst_n                    (cxl_cold_rst_n),                    //  output,    width = 1,          cold_rstn.reset_n
		.cxl_rx_n                          (cxl_rx_n),                          //   input,   width = 16,                cxl.rx_n
		.cxl_rx_p                          (cxl_rx_p),                          //   input,   width = 16,                   .rx_p
		.cxl_tx_n                          (cxl_tx_n),                          //  output,   width = 16,                   .tx_n
		.cxl_tx_p                          (cxl_tx_p),                          //  output,   width = 16,                   .tx_p
		.hdm_size_256mb                    (hdm_size_256mb),                    //   input,   width = 36,            memsize.hdm_size
		.mc2ip_memsize                     (mc2ip_memsize),                     //   input,   width = 64,                   .mem_size
		.ip2hdm_clk                        (ip2hdm_clk),                        //  output,    width = 1,         ip2hdm_clk.clk
		.ip2hdm_reset_n                    (ip2hdm_reset_n),                    //  output,    width = 1,     ip2hdm_reset_n.reset
		.mc2ip_0_sr_status                 (mc2ip_0_sr_status),                 //   input,    width = 5,            mc2ip_0.sr_status
		.mc2ip_0_rspfifo_full              (mc2ip_0_rspfifo_full),              //   input,    width = 1,                   .rspfifo_full
		.mc2ip_0_rspfifo_empty             (mc2ip_0_rspfifo_empty),             //   input,    width = 1,                   .rspfifo_empty
		.mc2ip_0_rspfifo_fill_level        (mc2ip_0_rspfifo_fill_level),        //   input,    width = 6,                   .rspfifo_fill_level
		.mc2ip_0_reqfifo_full              (mc2ip_0_reqfifo_full),              //   input,    width = 1,                   .reqfifo_full
		.mc2ip_0_reqfifo_empty             (mc2ip_0_reqfifo_empty),             //   input,    width = 1,                   .reqfifo_empty
		.mc2ip_0_reqfifo_fill_level        (mc2ip_0_reqfifo_fill_level),        //   input,    width = 6,                   .reqfifo_fill_level
		.hdm2ip_avmm0_ready                (hdm2ip_avmm0_ready),                //   input,    width = 1,       hdm2ip_avmm0.ready
		.hdm2ip_avmm0_cxlmem_ready         (hdm2ip_avmm0_cxlmem_ready),         //   input,    width = 1,                   .cxlmem_ready
		.hdm2ip_avmm0_readdata             (hdm2ip_avmm0_readdata),             //   input,  width = 512,                   .readdata
		.hdm2ip_avmm0_rsp_mdata            (hdm2ip_avmm0_rsp_mdata),            //   input,   width = 14,                   .rsp_mdata
		.hdm2ip_avmm0_read_poison          (hdm2ip_avmm0_read_poison),          //   input,    width = 1,                   .read_poison
		.hdm2ip_avmm0_readdatavalid        (hdm2ip_avmm0_readdatavalid),        //   input,    width = 1,                   .readdatavalid
		.hdm2ip_avmm0_ecc_err_corrected    (hdm2ip_avmm0_ecc_err_corrected),    //   input,    width = 8,                   .ecc_err_corrected
		.hdm2ip_avmm0_ecc_err_detected     (hdm2ip_avmm0_ecc_err_detected),     //   input,    width = 8,                   .ecc_err_detected
		.hdm2ip_avmm0_ecc_err_fatal        (hdm2ip_avmm0_ecc_err_fatal),        //   input,    width = 8,                   .ecc_err_fatal
		.hdm2ip_avmm0_ecc_err_syn_e        (hdm2ip_avmm0_ecc_err_syn_e),        //   input,    width = 8,                   .ecc_err_syn_e
		.hdm2ip_avmm0_ecc_err_valid        (hdm2ip_avmm0_ecc_err_valid),        //   input,    width = 1,                   .ecc_err_valid
		.ip2hdm_avmm0_read                 (ip2hdm_avmm0_read),                 //  output,    width = 1,       ip2hdm_avmm0.read
		.ip2hdm_avmm0_write                (ip2hdm_avmm0_write),                //  output,    width = 1,                   .write
		.ip2hdm_avmm0_write_poison         (ip2hdm_avmm0_write_poison),         //  output,    width = 1,                   .write_poison
		.ip2hdm_avmm0_write_ras_sbe        (ip2hdm_avmm0_write_ras_sbe),        //  output,    width = 1,                   .write_ras_sbe
		.ip2hdm_avmm0_write_ras_dbe        (ip2hdm_avmm0_write_ras_dbe),        //  output,    width = 1,                   .write_ras_dbe
		.ip2hdm_avmm0_writedata            (ip2hdm_avmm0_writedata),            //  output,  width = 512,                   .writedata
		.ip2hdm_avmm0_byteenable           (ip2hdm_avmm0_byteenable),           //  output,   width = 64,                   .byteenable
		.ip2hdm_avmm0_address              (ip2hdm_avmm0_address),              //  output,   width = 46,                   .address
		.ip2hdm_avmm0_req_mdata            (ip2hdm_avmm0_req_mdata),            //  output,   width = 14,                   .req_mdata
		.mc2ip_1_sr_status                 (mc2ip_1_sr_status),                 //   input,    width = 5,            mc2ip_1.sr_status
		.mc2ip_1_rspfifo_full              (mc2ip_1_rspfifo_full),              //   input,    width = 1,                   .rspfifo_full
		.mc2ip_1_rspfifo_empty             (mc2ip_1_rspfifo_empty),             //   input,    width = 1,                   .rspfifo_empty
		.mc2ip_1_rspfifo_fill_level        (mc2ip_1_rspfifo_fill_level),        //   input,    width = 6,                   .rspfifo_fill_level
		.mc2ip_1_reqfifo_full              (mc2ip_1_reqfifo_full),              //   input,    width = 1,                   .reqfifo_full
		.mc2ip_1_reqfifo_empty             (mc2ip_1_reqfifo_empty),             //   input,    width = 1,                   .reqfifo_empty
		.mc2ip_1_reqfifo_fill_level        (mc2ip_1_reqfifo_fill_level),        //   input,    width = 6,                   .reqfifo_fill_level
		.hdm2ip_avmm1_ready                (hdm2ip_avmm1_ready),                //   input,    width = 1,       hdm2ip_avmm1.ready
		.hdm2ip_avmm1_cxlmem_ready         (hdm2ip_avmm1_cxlmem_ready),         //   input,    width = 1,                   .cxlmem_ready
		.hdm2ip_avmm1_readdata             (hdm2ip_avmm1_readdata),             //   input,  width = 512,                   .readdata
		.hdm2ip_avmm1_rsp_mdata            (hdm2ip_avmm1_rsp_mdata),            //   input,   width = 14,                   .rsp_mdata
		.hdm2ip_avmm1_read_poison          (hdm2ip_avmm1_read_poison),          //   input,    width = 1,                   .read_poison
		.hdm2ip_avmm1_readdatavalid        (hdm2ip_avmm1_readdatavalid),        //   input,    width = 1,                   .readdatavalid
		.hdm2ip_avmm1_ecc_err_corrected    (hdm2ip_avmm1_ecc_err_corrected),    //   input,    width = 8,                   .ecc_err_corrected
		.hdm2ip_avmm1_ecc_err_detected     (hdm2ip_avmm1_ecc_err_detected),     //   input,    width = 8,                   .ecc_err_detected
		.hdm2ip_avmm1_ecc_err_fatal        (hdm2ip_avmm1_ecc_err_fatal),        //   input,    width = 8,                   .ecc_err_fatal
		.hdm2ip_avmm1_ecc_err_syn_e        (hdm2ip_avmm1_ecc_err_syn_e),        //   input,    width = 8,                   .ecc_err_syn_e
		.hdm2ip_avmm1_ecc_err_valid        (hdm2ip_avmm1_ecc_err_valid),        //   input,    width = 1,                   .ecc_err_valid
		.ip2hdm_avmm1_read                 (ip2hdm_avmm1_read),                 //  output,    width = 1,       ip2hdm_avmm1.read
		.ip2hdm_avmm1_write                (ip2hdm_avmm1_write),                //  output,    width = 1,                   .write
		.ip2hdm_avmm1_write_poison         (ip2hdm_avmm1_write_poison),         //  output,    width = 1,                   .write_poison
		.ip2hdm_avmm1_write_ras_sbe        (ip2hdm_avmm1_write_ras_sbe),        //  output,    width = 1,                   .write_ras_sbe
		.ip2hdm_avmm1_write_ras_dbe        (ip2hdm_avmm1_write_ras_dbe),        //  output,    width = 1,                   .write_ras_dbe
		.ip2hdm_avmm1_writedata            (ip2hdm_avmm1_writedata),            //  output,  width = 512,                   .writedata
		.ip2hdm_avmm1_byteenable           (ip2hdm_avmm1_byteenable),           //  output,   width = 64,                   .byteenable
		.ip2hdm_avmm1_address              (ip2hdm_avmm1_address),              //  output,   width = 46,                   .address
		.ip2hdm_avmm1_req_mdata            (ip2hdm_avmm1_req_mdata),            //  output,   width = 14,                   .req_mdata
		.ip2csr_avmm_clk                   (ip2csr_avmm_clk),                   //  output,    width = 1,             ip2csr.clock
		.ip2csr_avmm_rstn                  (ip2csr_avmm_rstn),                  //  output,    width = 1,                   .reset_n
		.csr2ip_avmm_waitrequest           (csr2ip_avmm_waitrequest),           //   input,    width = 1,                   .waitrequest
		.csr2ip_avmm_readdata              (csr2ip_avmm_readdata),              //   input,   width = 32,                   .readdata
		.csr2ip_avmm_readdatavalid         (csr2ip_avmm_readdatavalid),         //   input,    width = 1,                   .readdatavalid
		.ip2csr_avmm_writedata             (ip2csr_avmm_writedata),             //  output,   width = 32,                   .writedata
		.ip2csr_avmm_address               (ip2csr_avmm_address),               //  output,   width = 22,                   .address
		.ip2csr_avmm_write                 (ip2csr_avmm_write),                 //  output,    width = 1,                   .write
		.ip2csr_avmm_read                  (ip2csr_avmm_read),                  //  output,    width = 1,                   .read
		.ip2csr_avmm_byteenable            (ip2csr_avmm_byteenable),            //  output,    width = 4,                   .byteenable
		.ip2uio_tx_ready                   (ip2uio_tx_ready),                   //  output,    width = 1,         usr_tx_st0.ready
		.uio2ip_tx_st0_dvalid              (uio2ip_tx_st0_dvalid),              //   input,    width = 1,                   .dvalid
		.uio2ip_tx_st0_sop                 (uio2ip_tx_st0_sop),                 //   input,    width = 1,                   .sop
		.uio2ip_tx_st0_eop                 (uio2ip_tx_st0_eop),                 //   input,    width = 1,                   .eop
		.uio2ip_tx_st0_passthrough         (uio2ip_tx_st0_passthrough),         //   input,    width = 1,                   .passthrough
		.uio2ip_tx_st0_data                (uio2ip_tx_st0_data),                //   input,  width = 256,                   .data
		.uio2ip_tx_st0_data_parity         (uio2ip_tx_st0_data_parity),         //   input,    width = 8,                   .data_parity
		.uio2ip_tx_st0_hdr                 (uio2ip_tx_st0_hdr),                 //   input,  width = 128,                   .hdr
		.uio2ip_tx_st0_hdr_parity          (uio2ip_tx_st0_hdr_parity),          //   input,    width = 4,                   .hdr_parity
		.uio2ip_tx_st0_hvalid              (uio2ip_tx_st0_hvalid),              //   input,    width = 1,                   .hvalid
		.uio2ip_tx_st0_prefix              (uio2ip_tx_st0_prefix),              //   input,   width = 32,                   .prefix
		.uio2ip_tx_st0_prefix_parity       (uio2ip_tx_st0_prefix_parity),       //   input,    width = 1,                   .prefix_parity
		.uio2ip_tx_st0_RSSAI_prefix        (uio2ip_tx_st0_RSSAI_prefix),        //   input,   width = 12,                   .RSSAI_prefix
		.uio2ip_tx_st0_RSSAI_prefix_parity (uio2ip_tx_st0_RSSAI_prefix_parity), //   input,    width = 1,                   .RSSAI_prefix_parity
		.uio2ip_tx_st0_pvalid              (uio2ip_tx_st0_pvalid),              //   input,    width = 2,                   .pvalid
		.uio2ip_tx_st0_vfactive            (uio2ip_tx_st0_vfactive),            //   input,    width = 1,                   .vfactive
		.uio2ip_tx_st0_vfnum               (uio2ip_tx_st0_vfnum),               //   input,   width = 11,                   .vfnum
		.uio2ip_tx_st0_pfnum               (uio2ip_tx_st0_pfnum),               //   input,    width = 3,                   .pfnum
		.uio2ip_tx_st0_chnum               (uio2ip_tx_st0_chnum),               //   input,    width = 1,                   .chnum
		.uio2ip_tx_st0_empty               (uio2ip_tx_st0_empty),               //   input,    width = 3,                   .empty
		.uio2ip_tx_st0_misc_parity         (uio2ip_tx_st0_misc_parity),         //   input,    width = 1,                   .misc_parity
		.uio2ip_tx_st1_dvalid              (uio2ip_tx_st1_dvalid),              //   input,    width = 1,         usr_tx_st1.dvalid
		.uio2ip_tx_st1_sop                 (uio2ip_tx_st1_sop),                 //   input,    width = 1,                   .sop
		.uio2ip_tx_st1_eop                 (uio2ip_tx_st1_eop),                 //   input,    width = 1,                   .eop
		.uio2ip_tx_st1_passthrough         (uio2ip_tx_st1_passthrough),         //   input,    width = 1,                   .passthrough
		.uio2ip_tx_st1_data                (uio2ip_tx_st1_data),                //   input,  width = 256,                   .data
		.uio2ip_tx_st1_data_parity         (uio2ip_tx_st1_data_parity),         //   input,    width = 8,                   .data_parity
		.uio2ip_tx_st1_hdr                 (uio2ip_tx_st1_hdr),                 //   input,  width = 128,                   .hdr
		.uio2ip_tx_st1_hdr_parity          (uio2ip_tx_st1_hdr_parity),          //   input,    width = 4,                   .hdr_parity
		.uio2ip_tx_st1_hvalid              (uio2ip_tx_st1_hvalid),              //   input,    width = 1,                   .hvalid
		.uio2ip_tx_st1_prefix              (uio2ip_tx_st1_prefix),              //   input,   width = 32,                   .prefix
		.uio2ip_tx_st1_prefix_parity       (uio2ip_tx_st1_prefix_parity),       //   input,    width = 1,                   .prefix_parity
		.uio2ip_tx_st1_RSSAI_prefix        (uio2ip_tx_st1_RSSAI_prefix),        //   input,   width = 12,                   .RSSAI_prefix
		.uio2ip_tx_st1_RSSAI_prefix_parity (uio2ip_tx_st1_RSSAI_prefix_parity), //   input,    width = 1,                   .RSSAI_prefix_parity
		.uio2ip_tx_st1_pvalid              (uio2ip_tx_st1_pvalid),              //   input,    width = 2,                   .pvalid
		.uio2ip_tx_st1_vfactive            (uio2ip_tx_st1_vfactive),            //   input,    width = 1,                   .vfactive
		.uio2ip_tx_st1_vfnum               (uio2ip_tx_st1_vfnum),               //   input,   width = 11,                   .vfnum
		.uio2ip_tx_st1_pfnum               (uio2ip_tx_st1_pfnum),               //   input,    width = 3,                   .pfnum
		.uio2ip_tx_st1_chnum               (uio2ip_tx_st1_chnum),               //   input,    width = 1,                   .chnum
		.uio2ip_tx_st1_empty               (uio2ip_tx_st1_empty),               //   input,    width = 3,                   .empty
		.uio2ip_tx_st1_misc_parity         (uio2ip_tx_st1_misc_parity),         //   input,    width = 1,                   .misc_parity
		.uio2ip_tx_st2_dvalid              (uio2ip_tx_st2_dvalid),              //   input,    width = 1,         usr_tx_st2.dvalid
		.uio2ip_tx_st2_sop                 (uio2ip_tx_st2_sop),                 //   input,    width = 1,                   .sop
		.uio2ip_tx_st2_eop                 (uio2ip_tx_st2_eop),                 //   input,    width = 1,                   .eop
		.uio2ip_tx_st2_passthrough         (uio2ip_tx_st2_passthrough),         //   input,    width = 1,                   .passthrough
		.uio2ip_tx_st2_data                (uio2ip_tx_st2_data),                //   input,  width = 256,                   .data
		.uio2ip_tx_st2_data_parity         (uio2ip_tx_st2_data_parity),         //   input,    width = 8,                   .data_parity
		.uio2ip_tx_st2_hdr                 (uio2ip_tx_st2_hdr),                 //   input,  width = 128,                   .hdr
		.uio2ip_tx_st2_hdr_parity          (uio2ip_tx_st2_hdr_parity),          //   input,    width = 4,                   .hdr_parity
		.uio2ip_tx_st2_hvalid              (uio2ip_tx_st2_hvalid),              //   input,    width = 1,                   .hvalid
		.uio2ip_tx_st2_prefix              (uio2ip_tx_st2_prefix),              //   input,   width = 32,                   .prefix
		.uio2ip_tx_st2_prefix_parity       (uio2ip_tx_st2_prefix_parity),       //   input,    width = 1,                   .prefix_parity
		.uio2ip_tx_st2_RSSAI_prefix        (uio2ip_tx_st2_RSSAI_prefix),        //   input,   width = 12,                   .RSSAI_prefix
		.uio2ip_tx_st2_RSSAI_prefix_parity (uio2ip_tx_st2_RSSAI_prefix_parity), //   input,    width = 1,                   .RSSAI_prefix_parity
		.uio2ip_tx_st2_pvalid              (uio2ip_tx_st2_pvalid),              //   input,    width = 2,                   .pvalid
		.uio2ip_tx_st2_vfactive            (uio2ip_tx_st2_vfactive),            //   input,    width = 1,                   .vfactive
		.uio2ip_tx_st2_vfnum               (uio2ip_tx_st2_vfnum),               //   input,   width = 11,                   .vfnum
		.uio2ip_tx_st2_pfnum               (uio2ip_tx_st2_pfnum),               //   input,    width = 3,                   .pfnum
		.uio2ip_tx_st2_chnum               (uio2ip_tx_st2_chnum),               //   input,    width = 1,                   .chnum
		.uio2ip_tx_st2_empty               (uio2ip_tx_st2_empty),               //   input,    width = 3,                   .empty
		.uio2ip_tx_st2_misc_parity         (uio2ip_tx_st2_misc_parity),         //   input,    width = 1,                   .misc_parity
		.uio2ip_tx_st3_dvalid              (uio2ip_tx_st3_dvalid),              //   input,    width = 1,         usr_tx_st3.dvalid
		.uio2ip_tx_st3_sop                 (uio2ip_tx_st3_sop),                 //   input,    width = 1,                   .sop
		.uio2ip_tx_st3_eop                 (uio2ip_tx_st3_eop),                 //   input,    width = 1,                   .eop
		.uio2ip_tx_st3_passthrough         (uio2ip_tx_st3_passthrough),         //   input,    width = 1,                   .passthrough
		.uio2ip_tx_st3_data                (uio2ip_tx_st3_data),                //   input,  width = 256,                   .data
		.uio2ip_tx_st3_data_parity         (uio2ip_tx_st3_data_parity),         //   input,    width = 8,                   .data_parity
		.uio2ip_tx_st3_hdr                 (uio2ip_tx_st3_hdr),                 //   input,  width = 128,                   .hdr
		.uio2ip_tx_st3_hdr_parity          (uio2ip_tx_st3_hdr_parity),          //   input,    width = 4,                   .hdr_parity
		.uio2ip_tx_st3_hvalid              (uio2ip_tx_st3_hvalid),              //   input,    width = 1,                   .hvalid
		.uio2ip_tx_st3_prefix              (uio2ip_tx_st3_prefix),              //   input,   width = 32,                   .prefix
		.uio2ip_tx_st3_prefix_parity       (uio2ip_tx_st3_prefix_parity),       //   input,    width = 1,                   .prefix_parity
		.uio2ip_tx_st3_RSSAI_prefix        (uio2ip_tx_st3_RSSAI_prefix),        //   input,   width = 12,                   .RSSAI_prefix
		.uio2ip_tx_st3_RSSAI_prefix_parity (uio2ip_tx_st3_RSSAI_prefix_parity), //   input,    width = 1,                   .RSSAI_prefix_parity
		.uio2ip_tx_st3_pvalid              (uio2ip_tx_st3_pvalid),              //   input,    width = 2,                   .pvalid
		.uio2ip_tx_st3_vfactive            (uio2ip_tx_st3_vfactive),            //   input,    width = 1,                   .vfactive
		.uio2ip_tx_st3_vfnum               (uio2ip_tx_st3_vfnum),               //   input,   width = 11,                   .vfnum
		.uio2ip_tx_st3_pfnum               (uio2ip_tx_st3_pfnum),               //   input,    width = 3,                   .pfnum
		.uio2ip_tx_st3_chnum               (uio2ip_tx_st3_chnum),               //   input,    width = 1,                   .chnum
		.uio2ip_tx_st3_empty               (uio2ip_tx_st3_empty),               //   input,    width = 3,                   .empty
		.uio2ip_tx_st3_misc_parity         (uio2ip_tx_st3_misc_parity),         //   input,    width = 1,                   .misc_parity
		.ip2uio_tx_st_Hcrdt_update         (ip2uio_tx_st_Hcrdt_update),         //  output,    width = 3,          usr_tx_st.Hcrdt_update
		.ip2uio_tx_st_Hcrdt_ch             (ip2uio_tx_st_Hcrdt_ch),             //  output,    width = 1,                   .Hcrdt_ch
		.ip2uio_tx_st_Hcrdt_update_cnt     (ip2uio_tx_st_Hcrdt_update_cnt),     //  output,    width = 6,                   .Hcrdt_update_cnt
		.ip2uio_tx_st_Hcrdt_init           (ip2uio_tx_st_Hcrdt_init),           //  output,    width = 3,                   .Hcrdt_init
		.uio2ip_tx_st_Hcrdt_init_ack       (uio2ip_tx_st_Hcrdt_init_ack),       //   input,    width = 3,                   .Hcrdt_init_ack
		.ip2uio_tx_st_Dcrdt_update         (ip2uio_tx_st_Dcrdt_update),         //  output,    width = 3,                   .Dcrdt_update
		.ip2uio_tx_st_Dcrdt_ch             (ip2uio_tx_st_Dcrdt_ch),             //  output,    width = 1,                   .Dcrdt_ch
		.ip2uio_tx_st_Dcrdt_update_cnt     (ip2uio_tx_st_Dcrdt_update_cnt),     //  output,   width = 12,                   .Dcrdt_update_cnt
		.ip2uio_tx_st_Dcrdt_init           (ip2uio_tx_st_Dcrdt_init),           //  output,    width = 3,                   .Dcrdt_init
		.uio2ip_tx_st_Dcrdt_init_ack       (uio2ip_tx_st_Dcrdt_init_ack),       //   input,    width = 3,                   .Dcrdt_init_ack
		.ip2uio_rx_st0_dvalid              (ip2uio_rx_st0_dvalid),              //  output,    width = 1,        usr_rx_st_0.dvalid
		.ip2uio_rx_st0_sop                 (ip2uio_rx_st0_sop),                 //  output,    width = 1,                   .sop
		.ip2uio_rx_st0_eop                 (ip2uio_rx_st0_eop),                 //  output,    width = 1,                   .eop
		.ip2uio_rx_st0_passthrough         (ip2uio_rx_st0_passthrough),         //  output,    width = 1,                   .passthrough
		.ip2uio_rx_st0_data                (ip2uio_rx_st0_data),                //  output,  width = 256,                   .data
		.ip2uio_rx_st0_data_parity         (ip2uio_rx_st0_data_parity),         //  output,    width = 8,                   .data_parity
		.ip2uio_rx_st0_hdr                 (ip2uio_rx_st0_hdr),                 //  output,  width = 128,                   .hdr
		.ip2uio_rx_st0_hdr_parity          (ip2uio_rx_st0_hdr_parity),          //  output,    width = 4,                   .hdr_parity
		.ip2uio_rx_st0_hvalid              (ip2uio_rx_st0_hvalid),              //  output,    width = 1,                   .hvalid
		.ip2uio_rx_st0_prefix              (ip2uio_rx_st0_prefix),              //  output,   width = 32,                   .prefix
		.ip2uio_rx_st0_prefix_parity       (ip2uio_rx_st0_prefix_parity),       //  output,    width = 1,                   .prefix_parity
		.ip2uio_rx_st0_RSSAI_prefix        (ip2uio_rx_st0_RSSAI_prefix),        //  output,   width = 12,                   .RSSAI_prefix
		.ip2uio_rx_st0_RSSAI_prefix_parity (ip2uio_rx_st0_RSSAI_prefix_parity), //  output,    width = 1,                   .RSSAI_prefix_parity
		.ip2uio_rx_st0_pvalid              (ip2uio_rx_st0_pvalid),              //  output,    width = 2,                   .pvalid
		.ip2uio_rx_st0_bar                 (ip2uio_rx_st0_bar),                 //  output,    width = 3,                   .bar
		.ip2uio_rx_st0_vfactive            (ip2uio_rx_st0_vfactive),            //  output,    width = 1,                   .vfactive
		.ip2uio_rx_st0_vfnum               (ip2uio_rx_st0_vfnum),               //  output,   width = 11,                   .vfnum
		.ip2uio_rx_st0_pfnum               (ip2uio_rx_st0_pfnum),               //  output,    width = 3,                   .pfnum
		.ip2uio_rx_st0_chnum               (ip2uio_rx_st0_chnum),               //  output,    width = 1,                   .chnum
		.ip2uio_rx_st0_misc_parity         (ip2uio_rx_st0_misc_parity),         //  output,    width = 1,                   .misc_parity
		.ip2uio_rx_st0_empty               (ip2uio_rx_st0_empty),               //  output,    width = 3,                   .empty
		.ip2uio_rx_st1_dvalid              (ip2uio_rx_st1_dvalid),              //  output,    width = 1,        usr_rx_st_1.dvalid
		.ip2uio_rx_st1_sop                 (ip2uio_rx_st1_sop),                 //  output,    width = 1,                   .sop
		.ip2uio_rx_st1_eop                 (ip2uio_rx_st1_eop),                 //  output,    width = 1,                   .eop
		.ip2uio_rx_st1_passthrough         (ip2uio_rx_st1_passthrough),         //  output,    width = 1,                   .passthrough
		.ip2uio_rx_st1_data                (ip2uio_rx_st1_data),                //  output,  width = 256,                   .data
		.ip2uio_rx_st1_data_parity         (ip2uio_rx_st1_data_parity),         //  output,    width = 8,                   .data_parity
		.ip2uio_rx_st1_hdr                 (ip2uio_rx_st1_hdr),                 //  output,  width = 128,                   .hdr
		.ip2uio_rx_st1_hdr_parity          (ip2uio_rx_st1_hdr_parity),          //  output,    width = 4,                   .hdr_parity
		.ip2uio_rx_st1_hvalid              (ip2uio_rx_st1_hvalid),              //  output,    width = 1,                   .hvalid
		.ip2uio_rx_st1_prefix              (ip2uio_rx_st1_prefix),              //  output,   width = 32,                   .prefix
		.ip2uio_rx_st1_prefix_parity       (ip2uio_rx_st1_prefix_parity),       //  output,    width = 1,                   .prefix_parity
		.ip2uio_rx_st1_RSSAI_prefix        (ip2uio_rx_st1_RSSAI_prefix),        //  output,   width = 12,                   .RSSAI_prefix
		.ip2uio_rx_st1_RSSAI_prefix_parity (ip2uio_rx_st1_RSSAI_prefix_parity), //  output,    width = 1,                   .RSSAI_prefix_parity
		.ip2uio_rx_st1_pvalid              (ip2uio_rx_st1_pvalid),              //  output,    width = 2,                   .pvalid
		.ip2uio_rx_st1_bar                 (ip2uio_rx_st1_bar),                 //  output,    width = 3,                   .bar
		.ip2uio_rx_st1_vfactive            (ip2uio_rx_st1_vfactive),            //  output,    width = 1,                   .vfactive
		.ip2uio_rx_st1_vfnum               (ip2uio_rx_st1_vfnum),               //  output,   width = 11,                   .vfnum
		.ip2uio_rx_st1_pfnum               (ip2uio_rx_st1_pfnum),               //  output,    width = 3,                   .pfnum
		.ip2uio_rx_st1_chnum               (ip2uio_rx_st1_chnum),               //  output,    width = 1,                   .chnum
		.ip2uio_rx_st1_misc_parity         (ip2uio_rx_st1_misc_parity),         //  output,    width = 1,                   .misc_parity
		.ip2uio_rx_st1_empty               (ip2uio_rx_st1_empty),               //  output,    width = 3,                   .empty
		.ip2uio_rx_st2_dvalid              (ip2uio_rx_st2_dvalid),              //  output,    width = 1,        usr_rx_st_2.dvalid
		.ip2uio_rx_st2_sop                 (ip2uio_rx_st2_sop),                 //  output,    width = 1,                   .sop
		.ip2uio_rx_st2_eop                 (ip2uio_rx_st2_eop),                 //  output,    width = 1,                   .eop
		.ip2uio_rx_st2_passthrough         (ip2uio_rx_st2_passthrough),         //  output,    width = 1,                   .passthrough
		.ip2uio_rx_st2_data                (ip2uio_rx_st2_data),                //  output,  width = 256,                   .data
		.ip2uio_rx_st2_data_parity         (ip2uio_rx_st2_data_parity),         //  output,    width = 8,                   .data_parity
		.ip2uio_rx_st2_hdr                 (ip2uio_rx_st2_hdr),                 //  output,  width = 128,                   .hdr
		.ip2uio_rx_st2_hdr_parity          (ip2uio_rx_st2_hdr_parity),          //  output,    width = 4,                   .hdr_parity
		.ip2uio_rx_st2_hvalid              (ip2uio_rx_st2_hvalid),              //  output,    width = 1,                   .hvalid
		.ip2uio_rx_st2_prefix              (ip2uio_rx_st2_prefix),              //  output,   width = 32,                   .prefix
		.ip2uio_rx_st2_prefix_parity       (ip2uio_rx_st2_prefix_parity),       //  output,    width = 1,                   .prefix_parity
		.ip2uio_rx_st2_RSSAI_prefix        (ip2uio_rx_st2_RSSAI_prefix),        //  output,   width = 12,                   .RSSAI_prefix
		.ip2uio_rx_st2_RSSAI_prefix_parity (ip2uio_rx_st2_RSSAI_prefix_parity), //  output,    width = 1,                   .RSSAI_prefix_parity
		.ip2uio_rx_st2_pvalid              (ip2uio_rx_st2_pvalid),              //  output,    width = 2,                   .pvalid
		.ip2uio_rx_st2_bar                 (ip2uio_rx_st2_bar),                 //  output,    width = 3,                   .bar
		.ip2uio_rx_st2_vfactive            (ip2uio_rx_st2_vfactive),            //  output,    width = 1,                   .vfactive
		.ip2uio_rx_st2_vfnum               (ip2uio_rx_st2_vfnum),               //  output,   width = 11,                   .vfnum
		.ip2uio_rx_st2_pfnum               (ip2uio_rx_st2_pfnum),               //  output,    width = 3,                   .pfnum
		.ip2uio_rx_st2_chnum               (ip2uio_rx_st2_chnum),               //  output,    width = 1,                   .chnum
		.ip2uio_rx_st2_misc_parity         (ip2uio_rx_st2_misc_parity),         //  output,    width = 1,                   .misc_parity
		.ip2uio_rx_st2_empty               (ip2uio_rx_st2_empty),               //  output,    width = 3,                   .empty
		.ip2uio_rx_st3_dvalid              (ip2uio_rx_st3_dvalid),              //  output,    width = 1,        usr_rx_st_3.dvalid
		.ip2uio_rx_st3_sop                 (ip2uio_rx_st3_sop),                 //  output,    width = 1,                   .sop
		.ip2uio_rx_st3_eop                 (ip2uio_rx_st3_eop),                 //  output,    width = 1,                   .eop
		.ip2uio_rx_st3_passthrough         (ip2uio_rx_st3_passthrough),         //  output,    width = 1,                   .passthrough
		.ip2uio_rx_st3_data                (ip2uio_rx_st3_data),                //  output,  width = 256,                   .data
		.ip2uio_rx_st3_data_parity         (ip2uio_rx_st3_data_parity),         //  output,    width = 8,                   .data_parity
		.ip2uio_rx_st3_hdr                 (ip2uio_rx_st3_hdr),                 //  output,  width = 128,                   .hdr
		.ip2uio_rx_st3_hdr_parity          (ip2uio_rx_st3_hdr_parity),          //  output,    width = 4,                   .hdr_parity
		.ip2uio_rx_st3_hvalid              (ip2uio_rx_st3_hvalid),              //  output,    width = 1,                   .hvalid
		.ip2uio_rx_st3_prefix              (ip2uio_rx_st3_prefix),              //  output,   width = 32,                   .prefix
		.ip2uio_rx_st3_prefix_parity       (ip2uio_rx_st3_prefix_parity),       //  output,    width = 1,                   .prefix_parity
		.ip2uio_rx_st3_RSSAI_prefix        (ip2uio_rx_st3_RSSAI_prefix),        //  output,   width = 12,                   .RSSAI_prefix
		.ip2uio_rx_st3_RSSAI_prefix_parity (ip2uio_rx_st3_RSSAI_prefix_parity), //  output,    width = 1,                   .RSSAI_prefix_parity
		.ip2uio_rx_st3_pvalid              (ip2uio_rx_st3_pvalid),              //  output,    width = 2,                   .pvalid
		.ip2uio_rx_st3_bar                 (ip2uio_rx_st3_bar),                 //  output,    width = 3,                   .bar
		.ip2uio_rx_st3_vfactive            (ip2uio_rx_st3_vfactive),            //  output,    width = 1,                   .vfactive
		.ip2uio_rx_st3_vfnum               (ip2uio_rx_st3_vfnum),               //  output,   width = 11,                   .vfnum
		.ip2uio_rx_st3_pfnum               (ip2uio_rx_st3_pfnum),               //  output,    width = 3,                   .pfnum
		.ip2uio_rx_st3_chnum               (ip2uio_rx_st3_chnum),               //  output,    width = 1,                   .chnum
		.ip2uio_rx_st3_misc_parity         (ip2uio_rx_st3_misc_parity),         //  output,    width = 1,                   .misc_parity
		.ip2uio_rx_st3_empty               (ip2uio_rx_st3_empty),               //  output,    width = 3,                   .empty
		.uio2ip_rx_st_Hcrdt_update         (uio2ip_rx_st_Hcrdt_update),         //   input,    width = 3,          usr_rx_st.Hcrdt_update
		.uio2ip_rx_st_Hcrdt_ch             (uio2ip_rx_st_Hcrdt_ch),             //   input,    width = 1,                   .Hcrdt_ch
		.uio2ip_rx_st_Hcrdt_update_cnt     (uio2ip_rx_st_Hcrdt_update_cnt),     //   input,    width = 6,                   .Hcrdt_update_cnt
		.uio2ip_rx_st_Hcrdt_init           (uio2ip_rx_st_Hcrdt_init),           //   input,    width = 3,                   .Hcrdt_init
		.ip2uio_rx_st_Hcrdt_init_ack       (ip2uio_rx_st_Hcrdt_init_ack),       //  output,    width = 3,                   .Hcrdt_init_ack
		.uio2ip_rx_st_Dcrdt_update         (uio2ip_rx_st_Dcrdt_update),         //   input,    width = 3,                   .Dcrdt_update
		.uio2ip_rx_st_Dcrdt_ch             (uio2ip_rx_st_Dcrdt_ch),             //   input,    width = 1,                   .Dcrdt_ch
		.uio2ip_rx_st_Dcrdt_update_cnt     (uio2ip_rx_st_Dcrdt_update_cnt),     //   input,   width = 12,                   .Dcrdt_update_cnt
		.uio2ip_rx_st_Dcrdt_init           (uio2ip_rx_st_Dcrdt_init),           //   input,    width = 3,                   .Dcrdt_init
		.ip2uio_rx_st_Dcrdt_init_ack       (ip2uio_rx_st_Dcrdt_init_ack),       //  output,    width = 3,                   .Dcrdt_init_ack
		.ip2uio_bus_number                 (ip2uio_bus_number),                 //  output,    width = 8,                uio.usr_bus_number
		.ip2uio_device_number              (ip2uio_device_number),              //  output,    width = 5,                   .usr_device_number
		.pf0_msix_enable                   (pf0_msix_enable),                   //  output,    width = 1, pf0_msix_interface.msix_enable
		.pf0_msix_fn_mask                  (pf0_msix_fn_mask),                  //  output,    width = 1,                   .msix_fn_mask
		.pf1_msix_enable                   (pf1_msix_enable),                   //  output,    width = 1, pf1_msix_interface.msix_enable
		.pf1_msix_fn_mask                  (pf1_msix_fn_mask)                   //  output,    width = 1,                   .msix_fn_mask
	);

endmodule
