// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
DHYyFcPzyNyhDJL+2oyzMz+qmeX/82ds3tHyVMTpui6qFdm4yOwwiP3Cq7sABYeW
xveijyajqhV/TASTW4wu7XhfnWOhSEB4XyVJZUVm9BHiXl0q+Me7Qya2moad0lhV
cG/cfrK86RROSCQCpUMFI7PHGf61SNsEg0yA6v0kSIs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 27536 )
`pragma protect data_block
Lj+3BhrZMxMv4HNV5JUiQBICsCK7HvtcSwRrPg6AQZT/e0oJ8EG0vj3uMs+/PDin
Rh/U4jWxhjFCmJ0pzJXAN9C8VZ1+cHMbrQJLEt0WwuV1lYuvICLPfzLacnd+ZlGj
GNM7PEX1iJ4nm7v5zZCMzNTaOk6tJE+3hctJLqgcLivQOMnOd5T5/imtDNdRZvjI
YT4RDEmb55oSSX29zA5CNjLpQ8tFPGjf9KO6WyQUPalEdFdr4synSO4FWz57puQw
vgBEQd5lN5PMSEONNvYeoSsE2aAiwwJ26JJ/PZXF3u0oKEOv4nPv0WrPFfFS+etK
utvLGUSUQ0mMCuoTCudRlO6T43+YQC9pxAOHnRbPNNbu6+FjEqCEgvhs3fhTp8eD
8cFvyvTDbO4TEi/eHHQOIdXs4j+wWRGeAsDI/2/BGn/1g+1xqn0tFPp/DiVtbQ5I
ioM127NqWUu+lMVoje4LaB8IswjhvqFShTN0bjI4O4f9Ui0RzDzYgB3s5M/6RGm4
iQ9XaxEgJPaYCyp9x1oTj7Bo9d2Wxry9ZihBdyBs0Gn+lZZ1Ag21t2oceOlvBnV3
3E8ixYUG+WV/qbZGELySWxSL0IifLVoFl/+BOiHHBLdTYahassN0wHQSAnwGmLqG
NQEsiiBNiPV71apc8n9rvGNX/JUXGWoaIoRDJubHU0SEZKdWUWwhKUX0WsVwUrr9
GSJymmVUoz6JSfk4+v0cgE4x2oTAKVSzl96zC1VjDqQLbhVmwBMHftZmDKGu2cOM
uZQWcj/3jEmD2OTPZTEwduCkyjt3u7lzGRifNJPIRcYNLfxfZYieGfg7Ma9UhZZm
/ggcu/bVNX0ApT98Y9Pi68Ll1G6sX0xSzPMRUI5Q7TmHp60CdSe7fV4u7fGqdPyM
TCINYrL7eh0y9HVNGc2Ez6oS3rIM6zipwDhgXWYnuxp3Tagqb5BFTwJV6aDtkA3y
pmfXRokIrFrJJstJVtAkyZZkGH1xikqWWfa87KsjysaXMD1didRRo5Y30KgNnXcL
RzU8jwvjKzZV/hxaK+JvN3dj2s7Tjid+EsaADmXr2NoJmTOMTmUVZMdoA/4Byw5u
f5e7j02GQ+vilJx+HGzwPOgYAo72r+P96g1TZEq9khHZKn2i96nJoc38YfXr9erj
MubXDbyu40O/CV+kMaGT+csMPy4VqRME4v0CZ2F51omKpFY3Kz1NJLKxeOLDHT7F
kzybHi/SOMDOPNJ2VfqH9cFNr5vwnP8ItxDv2WOrAY0MzamhjwrPlp6016bCHT71
U4shfgJjgnN6HjR4Bh62Rs0WC9gg40kq73OJMwRLsxlVNF36SirA4NtbNUCFqCTo
RKDLHTxX7KOPZM8J9H+44MLrKRhkweHWPr6LN3k6xti+MEM/EHSmtgyWazO++qS7
eTqUOJlHOj5sa902iQHY1j59GvMrGW6JBzFrbwSKptKl3YvtY0Q72Q9dGxYe3UE4
xs8Lp8pAO/adsqiccXQGK1kFt624ou0tLQ3ciqM2YxtetpnsKvLFwxiz9Xm26f7a
lptrf+p/sW5mJoPOaZanZgdGDSpYJUjBeW3O0IJIAk1pj8UCYJokPbCR+TMLxupP
2QWYPuuOtAf6vLd7k1GDsnLWjV+6Z7JsEtOJrgOOcv7n66pLfLrC2g1J/0EJmspr
ZtDWQatbWv2xuI3VBU3wAG19yFy2LD/NYZoB1EV02rl+EhjIAaISILOPOwJ9kncG
m1yQdG4c3nXz0S2k2Z/ZfJEB1cBJJhh+veyk1zqWySpiDNfNYNGtZJ2uox71E84G
oH5655XcFenJXuTRQ1C3lzv34brayStetSzHV4IZORSvw1j9qOAyC+qf9/1Z1eSd
d32hfj1m10qgFQgIKsY8CwSzHMPoTJsevprlILoBpD+BCaSa0RqSBuh2ZExArHWr
xKu4ZBBJnPRFuqG2b+pU5BM4+TvHNLy4FQKlWCN0ZfA4k+qYZTV6kyuvQe6F10CA
dQlRqA3FRCqU/5pcWpu4XM4lyZbUPp34/qd2GtS8dpgZNaqxrQwXap2eYAVS0Uby
+1Bmbsktv/GcvsRiRMGQEs165Niny9TVouV2drbgs2aoitDbc77qyzmfLRFzLiHL
bp5VGWzUnAD10jbzQogtCYC7PiZBn7iJAAX45esO5/o6dpcHs8mQhfRNeDVIB0Sv
vP8wgnZGwBvdsBg8Rg1XZvYwC8Z87Nc3qtcYWcZjqKEQqUZUBuIIleGRUgaV0BVR
Vd14hB3s+6dRYwMTdm2ME7mPCegbFrcH9Y++cv41KvM4VU9AZDfueG+3sA0HUsF7
g/2uz4yFWTDbOxe0+zLnWsWiZ8StN8ZjCtoeOpXXvW+dq7qqQDS3uZoNF5uQq8y3
rnXQIevJ0YXp8uhNNWEQId82JcfPHB742lQwoJafZGmjt7fBbNSi+DZROfNZ7i+I
u+NPJlJKN43NxNBzFLnbG3QI7maZRml4UVTRnQdcO5yw0kDVTnSCVqEjxD/nQ37B
zimTlVBl2oKaI/xbN4SeQ+2b6AnVQnWnHdlNCjNEniRqz1Opr8Qn3pu/duwiIkq9
ZBV0ILR+74ucaCk0OWD9kZtdS6yfBE4IOrBlOQgclbv67DqOsMKuvQPhCGy280+4
wKYEsTXZa3hbG04ImWLuxJma5sc9tGAjTUkYVdEDLMzvk9kaWB7i1GkvX6+Z9tsl
h8xYbkOEOAUkA52srPTZbD50lRrlCaPjROGcWOtGb/IrqCKNR24d7FLqfuAhTvBh
Z1QlQOtxfggkzAYHSSsKFRRLWzYGoaur38KBJZzvROSG5BeCjKDGOToy+PGnbBOs
DfUYfT6ZwD8dERsS+M/2BtYBXePGa7gMMS7bjbGkytuC5JifPylRbBJdeiADX3uL
F1kiu1tFwtTLmr/l3UYJCc9n6Ka3FhOe9ICtaYTNgzLd2lTMMZPBmGYnNeB4QDlI
aYmszIOr75W0kjpmv/ioDmETScx8fjQseXZhfijBJTbsCUaZIvv4y5otJ/wAbWEa
GKW7A8G53cuzUF/cH7CnliSypXDMFEhQUvOPtPz9rriX3AVROvjg+6iHKM9WKQIl
vzA4QXXE9UBob0LN3S86nr9ervrCGqpISysn6e8OBjOa5Eb6HEz04M5+NpfQhHCL
Qcn5alCOM4NxBmVEphnxPQg2/9BHB9P3++aPnsCcUkhfoP3F1Z7tamuq5BQHm5Al
P9M7rqNowRE3KBd1pTe5TwLQn+bbyqPfDI7ZLDFrvMjgng90cXJnyrm8XYy/0EIB
hp2ig1Kd6z1q58TcGpEVVAxOgyn/7c4waqsd7i1Bc6eVDxqONuSu18iCuJ3ETmlx
t5QcZMhyBe742ernvjMouJhgJNlZIrr9iDYiKvh6EzN0bNDScyz0fcMMZD88YvVd
YBcDt/R64o+wHWzK7v1Ain/Gd3zjIIeUH+56P3b1kSd5rsSb7mL+EPWkjCPL2CXo
J9O/x/88IVQwmbO3xP6fVcFSKpGnk8moJxfm3kriPuTnhCedRptkLn1IK/kKlT7R
0Ou3czEoLkVfGingNUMLPFypi9rUDcR7l+pvXSpt/yuRj00Y8ZoAF8v6vvruswyF
7wj3iFGJhm/+Wf8BNKAoMTnups73J7WGjgWEbLJLinBqYYpWPV4fAECivh+w+U34
X7KHF6ZVjQeClcjuklXrC+zm72gZmc+e3ZlI96Ame8D2dDOe95yUSnTxE18tvNFY
IAx2ZCTpw/UpubU4xHWVqOC9n2hk4XKV1UCXchfrDqlyZq5sIWbS2QyVjJug4QrL
0z8kjQvRSxvzJTyiwcRILyPpJRTOVvIA+fFWPVovEG0OGP+ceCvLc+GNle5/GXr6
EhdnkNScPpYXivv1soyxMvUcFzBUeFWIoPOtreQRgDGBSb40PNpUJiLSomkFL++5
DdH3o4/RgiiR0G0ncmurXWp5mW35gnwl9NT7D9w9FX90ntjPK1ERuKZdz5nhPai1
K6epdjW0kne79bNtVG/yAHtBMnwgN7xA+kNL8gY1YEPe7r62g+YuKVeTYtzP7UBY
o/wCnKXYO2ToEgFkIyRwEtxq+WEgCnhK6HvXMX8+nsGqVS80UOhuBnNFyoFFVHtn
EE9ak3/iHvq0tScgrGQF8wmzRHZqK2WaT4kBKTA1w1sX21LdhrJFA6noA1Fy71wA
YukvmFP9CSoF6jIkRB0TKBjp8ZthhmF40i/JxT7EszCGWI45qNfT6toaLjS8ejNY
iF8Bsj2IX7ZBRpca1dQOB2RP3BYH4YQ5g589Z3CU+FnRywaef2OmlPQENcuWZ3TY
ii9UbinNvfqUiPV8KkeOdUkcirdJwZlVI3NSG+fZX1tz5DGE2u3SYDFsxgOpfdr/
Id6izzg4DvlqhOLSh1Rs3Bq4smZT5VzWJ3648PjSkCw8G7xp4dXSGCtAySyrURrw
DB451Cft/4WYHr1/8tXtN8gecx3mVAkXOq3mqIUlYdN/P9RYsGuS8tN75HkKsYB5
9fC4v97dHhAT8fcOu3m/3KhK/I+cqMXokILsT+7wbrVh2LE+FoV8DSAoONBg1f3z
qa0CILDS7yz6KPfgzcwEO4075KIPOqkJXc+ryqg2+PB2906JiUt8FomGZ++2ZbB9
4Bdq3ZPKzhwnyHBmKyiWVSszOc3tFr+Kkp0CsyzjXrnCn27rn+er17JYvY87ZH7Q
WDXANS/mspWOGD+mWvrf0cmLdp84SbuAwtTkziznIdDkbC+uUqLDwCKpiTgHfkKE
2c43PvZhX542fux5gAe0ixWuAtWSnSHNJc7PC3N1AyRXjDkXkEGOKkgUsP930yfs
FG8YaB3iP/WWhmfgnUBVKQlZQEVE9c4mHINmKB6XAtuC6BfSIo0egTrOuEYDL1Bl
VXbEiYXTE9JiYPhIWPTRZqs0YQiM4RnX0crRv1BEFC2wo8AM8U1Iiyw9PF5dXwfj
+l2lV+x2CNBE4vEBaKxSPZLjNLRgzxrfCYoWu26DER9jvAjNxewExc8uBlyTsLNl
p3IvVhHW4vACS5QaLjsNFugfiJApLOc+ubfOn4pOUiS+ysT9JeqF7KAF7AHIbrcK
wKEFQ8flH6J1Y+rPKBiUz8dWrRrUF1fG21+VmIrBjWc9wGASE3W8phk7YGb8lSXU
5ZEM0gWN5jURPXrXEcG9TlxXc3/S9kEbUTS9bUTUBecl0lxMRE0pLOdDR+pXmjxD
UjxZIijwIvW9+dXwMGKHg9Q8ehBXoNLb7vgq2ZDb18g7mqR5Sa+/6hekxrb6bxOJ
hD1U2KH0jKCNaTFc0x5N6c6vcQecXl5rvOfYlj6GA3eIhFiqEhAOauUOj1Dw3Ipr
M+QpOEJg8PvFH+u5s7G51hqJfUnqyqG7ixtYXpdragqz1jJM/MhUOak7uEa2FUJ+
mmNICGrmWcxNG0vEAMgG2fUBhlM7w0k2n/C0AraPjiKK3KCKG31SLr3Rfg9rrBXM
eQe7DI0B2q2tjhzt+IDqBOBmmwCelJ6bUVsKtPrtMXL5N2OyKDHH4NmUVSU1aQeA
i6OV+VGX6qYL1ZAwbE/sRrJTyZnosP7C8leqRZPKDYl0b2R4S362Js47pYvArWZq
jZvRia9B1D6hy0lK7fqzjCXHOuKwi0sZ1SkIS/l8J+nRJVTUYo9AzqHuX3JB5Wl9
HQnJaDd9OLb/MMT8p5nj/mVLwgPL3tIHv9sFRUCQ0vYv+aDf+KfVqRuAlajY4TVG
jSBfJoKRGrBee8wHUj2hO8WZbrS9AAA3E0qorVgzeSEBPE3zx2sI2sgHs9f3uLRu
2lDMKgCqYV6usE7I/g2R2BtGmRbEMPt8kUvaOAucuSXv3AHjZI7uzOamRWjx62bo
s3IBPwnnIPWBkYss0uuzuPCI62UBO+01/QdcdKjaIFx9T6l0UuolvFZ6ZuovkdFa
lMPS+sw/sp6H/Luk8rWaGE/yqQgolJhyDgD/FT3ETIckkkWDi5Llv+W2lpiytQCH
SXPtSmzBSXe/4b47mQh0ZkHo07Z5+A6So6kAlXRPjo6+eXetkRafZS2zZsD8FQtV
2nowv5Nn9ncR44z8GMzIIIs7SPN7WQu19Gy4BNzKntJE4CXLO00GvhF2MsaWKGKn
IBeDLL+tzObiWVbdFRv2i+FeTorHIXTHPOhpOER3ebBG2SLo+03VxvYFHBt8cZj2
THXNcr9XLCGeykoHNnYDWYQLRGjqgg0TWWA/WH+TvmWvawxTkBD3RIh7iKJlMOdv
rLodbDCRGH3mtBSGnd82FJ2nZjJmZ/5h+6c3UDm9dzFXD5p7PDCLcbS+qH2EDYuk
O6RCanMYJkjWMzhYorc2k4mS4RcvIemVE7RvqGOYc3RgLbzAAtz2BilCd6LVnlw9
s8fIFi5bu2sm3oULJ51lfbkHXHlIkPYsuZXSkSSV0NmC9LqQEjDsXEmF0CREViza
MeBfRLfCavigF3U2ENc3s0FtFAImT4o7I4nO1RlHNWdTXfpw8MiLAx7+VcnACfTs
/pdIJnk8yK79UvxfpXRPgrWYzvLsuC54vibo3+ZTvPeVkzAHFkrAGaPZV7RpqlOL
2fkUAnne1UOtwFYm0KagRQfr9UZRt0uo5pcwB6HVBl3OdyjlvncfR8Ao+lO/tF4O
iirzrsBknGlhBshyfZbYaQQb/SaIBPqeMCBNQ42yjUg/nv+jajWUCBlR2QQ9HiuJ
X+HTyQ5TJNZDVus+orsubgJO/MiHPPOzs/VX4GobUl4//q3mZs86tQGHI4R1ng6P
TbKKwF8W3c3LXtq9L7idcNlT/VNnOdi5o2SbP8Rda0vq1cJzNQlJF8KZUmqb7xSI
B9lfUHt1qwUv8mBfHQf9V2OthHg3+ZEP0Tj4/AWZUN7AEh2rygEBTUiZNYZIHg+e
mJLU/qbUOX1Be8VZrS4BwpPbUzi45ypm43AGz8Hou4OaA7sVMu5V5yR2OGoQcCs/
e7/tVwg+ODrwYdWaXkxISvL8klnCpykZhRYJKPsIyqTDm8avgOYDAqXfX1PkLOjm
RCUS+Rgf3XJV12naAheSmpOsL0l6BcRQs7JOw/5trvYxJIYXhT54EmFfP5f1e3Z3
ztQC6EPJKGHH2FgDaE000xGqba3IWY9x4F8lQp8vydr2RICHkxvEZTdHQmzfJyU4
YEOW/6riI85kF5oIUyQOcY/APrEm8aoRmTKJqBL4EH8g1jccYAwthGNGoZPGe2aA
R0a6HJWbFMmokVBlRXuHRTQh0Dy21PqwDOXW9stCnLi/Px8duSxrYhkgD4//oZxN
G93uRQlU+tWEJmCggtsPehdDU7VUOoiK9Ff4RgFcemOydDovMwF5Tqh2Klaga9BM
qlNLDXowYKz+NFUm2jSwltZ2TOfNjC6jK1grbEsUGNBn4NZriShlmxyCX3ajpzFT
W17vUjbLRF0WYf08DAsSk4JCZL/icOLK2EVM4TOi8PFhH2UlpJ1lMPdYKk04QoBG
oXFp0x3TPLes36kP5tWsi5+SQDW60yfdpL0pzqX93RffsKoj+CbPdXZ+FZg4eVB2
BI/dSL0bI35hm9/gNZX3dKRn6EGcOVwqhcKgHQUOMHjuUAfKZFvglchTF+hNZGki
0HjoLLVMQB2uAI23fdgvSXOgLpyTlKkcSDxF8ygCJp7pgAFxl2AQczDgFZpZxH0T
PDGEW92YnExoY1wMXD2VNxgnOIVByes2h8UV34OJkWhzbSsYjJHU4W5aqo7bDp1R
IIieGpanbugjgQX0AAJ5aRr0he1a1VVFcwI315Ig4sNmoAwrjgup3xsHVvTOjsne
Aq0MlzEVSRDla2XuAtLNspaIixxIL8itbKmqfIUYFaBnxJy55moGdN7i6ipNCAVn
Ggr2l6UAjn0DVZf1QKj+Kf7gwza8spefdA9J6wF8ZyfsocQ5fk7gMslYNxwqZkGE
PtngLr1IbbaBhgR7wAUoS/0wGC67xVF7E+Jm0UBzbRlz93maPhiZCCUbTBX3jNgJ
RpW3ORd0cgZGhlXdCBW2jc4ge54CTEvm+OW5F4mdvQTtOA+Hv1iIGeQPgX2q7Oa9
U1Vl97moE2KVwjOfyo07FYm94y5I6sytQCIEr2P9NsjQZGEovIunVX/eiC0lTeHX
2TBLV3FmzC7+MYx/7pAsdxu0RVCI0zj9+FSO6Jvm3Edhxc6BMSI+Aqq5oySRPDeB
pnvwEHYpbxQiKqTCp2EQ4GZAL+KdkciRdV2UH1F2YeUfCk2m2REU/Xu6sInxox7f
mWArS8rM6DlrCEQMmzRQ9tqmnNiPQ5T9zOFzv9kMtAsAHqaF51ijM4bWATzRDUM0
BP0B+41pu2um0gX56IKNHC73aSu7HI+3rHORSeVQDe54Fgprvhkjl1pUPMtenea3
dYwM3QA4ZMczMIEGtCMDjrdeJCxJRq3tFOaIeEe1LxCdrP8DvQxR+f1gewUy1SU1
2TsajPG9cH44whiJuGuAYZ75YyP2xnTNbb/D85tF6AyEKKRfjmPcmapFoAtUEG7f
g9+U29w3uaFqr30vJ2a25HtDnVXJ4H94nZ9jlew/3SgUnU+xjdejxxNOXPJTExRj
dFs/NE8i/akRs9sDscyT5ZxSJ/o2crbKuGHR3XtDkNivZjlHEmMpShTJu8Oe4acm
ZU5jTBAqI5ceP0D2CCcZzSmDXK9CtlwcnRYXDsoZd/mkrG76S29uCxPVMkYlsleq
wq9TAIDxiON0L1yocHyRLWoInVIdo2fAipLUVD1xENHw70A3JRtihOwrIuoQipD9
YFxwriatYM4qUQN0ux9gfpr0N/hQar8Eb1i5ESHtzpAYfEQPr2eiHA9qPFO0Uyyl
Slyh6L+XsXOCkmVuG9ohN/XcTlx3I3hzDXxKGqG1YMoLUL8wDr2Ut4cF6HQ9BWQU
Lni37wIlDWOgB6r+V9MWaFEeeTVXSscO4dH6hnkFYYoena9yJXTAMKRkFVYe99/f
Frbsh4/xz/s5Jf8UCQP45tmRKfwUe9SWgt0AO0EiVxR6xrLIPfQXDbfC2/+XXvR4
PJHLX9NidVDfnkxXO6cp2k3Ziou6ysozDGtL/W2B4C7/EHhOZleWCzf53m3RPcCP
LjT9rSCVq0KGm+s9KsUCv88oKNSGxu/zcV8zspkgJ6A+SHJ6Kvvmu71hR+7yg50h
2S/SaWxmCI6Gg0TIBA0hkNxmkRLelp3kc4rk6lte3LkFBBh7Vs3Ppr8/l7M424JI
JbDi20T23gQHtQtUlAMmTaguKTR2GK894OyZp1irrtJuOhpxEOX/LbUOZw4AD2Op
54AI7ulOoNZkHjXxSRBZOAYNrlrThcgEjBJ5345NbVnh3Lh5g8MSM6WONrgvgLc0
lShYG8rYlLAhD6YIZP1doxXlYzKKv/yO/YmAG6cRQbSP2Kxusfk98NkhdO3tSDrb
/jAx/B/HftucnJQQ7vPHeIAHxcxHibtKnStM36Dbts4pJGruOTFHzbjKM8uwgpoX
ZkKIpHYy/7juoQgnFoXEmYUi7hz2svXosmQcte8vW450BZTSQOIX3kucWBz0GBxa
AKRluK0sFyNbDpPfrKtCRQyMLPQZSS9tZcUfhZyCvVu+JSxIVXHRY60fcplsgn8K
ibrUtP9kvcQlOWebJGFFYsuaafiRcENOny5Eiz9mhJ8K4SdphMhEYlTUWwfW0XAf
+JcrXuT6Fj2OKl5pcShMADx8v4kINrqjO5johZz/hb8aDp7I1JQ9p9/I5iHL9BLx
pK4x1YY9GpIDr+t0utH8GQAU0FsJUD2c2jNGCxo9LGw5uKW6+P/MhF9py+prR+87
P+bOzmuKo7hQG3KJ3MHtZCzNhI+7rA4Cg+YsyimAeQ14lmAh8frC4LhTla/1Gjpw
3n5cL+jFBkScGZNhsZ6c/GoSF2HwSrp/tP1Hu0gyL/s64e54GbUxlx4Jy+Q82AR2
9pm8UCbH/yT6T+tqgta4ASQh6N3jh9NiiWD9Ju+8v3FRHSyssEN4th+OHBFVRX6T
hX4UNoYsnf8KCN6jIteef26I6ae8JjxDzKOcYGaqAYsXglSnECgq9Budfbh+xE20
C8e+WypD6+nheSHs36Q9nuoVOKBfEy3e74PluKlV8B/Pt5/luey1vp7DlkNmkZ7I
A9ae4U0UJKzTFnvR4S3FiOdsd1dpUHNEtga8uOllzgwKM5fzWSmJ3qJDRAjDwCAH
nq5/QoLXUHNm7rPrsCvAu49/OfBUhvT68NSVjWYqRdsCQ8xSQPI+iV+8042vJSzI
Del8/jICatYkWrO8KXy7Gd8fg2uJbDC7mL8XV/bQQVBbhyeg0jb5pVNqUYSYbpKA
f3VkaL9jTJMtMscfHka79XvuAI+cqeve5xQ0n1Mdu4/hAcOJACSeWmJ+ot0o6/rF
Gd2YvBmXOYW15wGCmURMQjCue4ipfn7xDSLQ4Zn6WrHoWxgiSKd1FuZa9uytm2KR
atjnESeSoXlHGQtMenGq2sBo2ZIM2wP6R2rOqIgDPiiS5qx+8B1OzN7PehOc+Vw3
ql4lZaRVuzAB1yAPPs9JjyvAJsh1tuibXIXfNb82HImSr3sVaiM3JT3mxK1uON0Z
+McLTn4ZWI0HqbMBKY4C/eUTk6s8V68wVvlV1wz2Ar/xdAdVNDnjQQfYX/Pd9n7Q
AvkMSb2XYU7zI+313uNcupupxqhmuYmQztkIvfmGz+FiRQ3b6g/URBMiVXaRcgTJ
fevvgOgbF6Uj4dxYgdIse9FKOmS64govX7vHDRpPuNAmH6Ra241JiOd5lmTK68qb
DWb5ZsUaLgfMxDMJy8L6kuNhnYwHQO1pzp0BtLLwOeo9Gx5dVzuVx188qRt594Sj
iKjrc2D3g/g+8C4jKSoQ9E7S01hRvGWU5I25VvJ4eS+PDPjN8n1LhhM7EOIjLh/D
Ecwy4oTsFMoSLjj+BONMqvy3rPFjdox8hPCqd06No7qBzwB2QAA8WDjdf8dhV8bU
l0HxiGJGpvV6VJrfviALuOYSg7qdWEgl66aMex0A6CAsTZ7+8NsHsSSMFnFyCXjY
+pLmx8Y+ymhPBEca644TwIoZA8xl20QucY6CdOHq1Kftaomol5vdRwQSeQoVyx6o
BLS0YvReezSIzx01wqjvTkWfGTBYqdPSww/C4vpD6x246VdqoJq6S3+2VCVgrid2
m9OLzpQEWfpAhVcRc2tBl76twwHH3ehLoADM/kZhYD6gyddDcMO1ylSsrg5rLRpo
WQ1M7mdPVE2UxxWOm7p6MYWNqKh+avZhfj8H9KAo9vT1/RvoUY7KVpv6axqEwP3v
AUj9l2mEjcS/KbegWjFis0c6FTKry7WhtrkHmozLK7w0Wg8X9oyP3cBbPbzwN35Y
Nu9B1gFlkYJJQ64/vAXdUNE+gcRN6FH1Ms0Ffc4TwTRM19ZedVoEf3LZFZcv341U
ibs5kwCArA7tsB3cg5GpFTLiwqPuRoPE8VBAW/SM2OkHwzeKgiysP3zzSuqCUUbB
b8GpHeXw30He0JbPHqV5GdA+4YtPND2ecZU/2ChGhRwYFg4CM1BUrtzG/CbSrtSA
y5JpYO2uWS7d9utCGE3VJRazmXcjzGSzo7FTNPcxUot1lQM9w1T5cTvppTT2xYge
yQUdCF5kob01YkcPxLtp77ijAh/ttngroOc2T9ndanfEJdu9mgXtMlHqrMW+cb1D
qhjd5M8aqwN7t4RqYap8fhLDRmAtOiboIfl4vEqKF7cS3iJ/8r865EFtqvCskQTI
0+FaCCaH6UWRuKa4qAkc1Au5OHLK4eIKgYNY+lHCYy5F1zyjUdBapFexcOe7GIQ6
qu+VYDYmmFoXl4LmmBHCP37FBcxYsAekpe4ohjk5YwtfIA0omw4S2MhXKNgtRpHU
PH+Hpya9nIu6rrsIOwE+5Gkw4Z1TzU/EezQytsgc2Lx1f5Wz6R8uK4EaIJ7KDgoo
VqoTTUI2rjIWoA59sY5HhC2yPvipnfnjBTqgskkhWSpf42xrhfCslTrchAgrVtdu
qCUIN/Hd/1uQfYBX6SlXCdQIQrHcWmYpiPpc7GcP2aUy/csxJU8LvcGEQbrp/ytA
9TOfrBzmMrLR1ZXi/19zU4/Ju0Q8ZVTHsKRtEwDNGmvsizPaLI5R8TNl+ZkAq6p+
agm3g8sU/SqGXTyh0+R1KTUM54e8/6NtJ5CWhJrVLkjw1GNxWYweNsVTh/Aq4CgX
Md1A/38bJmA/f0hOwakEDo+sgVoN/QamFCPCuGIGA7SAzUnm86qFGTOcZukTfD8U
PmqmLahQx0901lCubZM0c7avMjqDVOPABn1Ds/IInS0QaADnpkqWYlcEb7Bcjdar
BqsVn2Dw7mdr6Ks6H75VQndyVbgX4Q5uVInIXXtewNRhPpxCNWOxFZSTDd3dxcQq
eZZ3rAx4k+Kd0TckAPdwiCdWw6n3va0gNbX2+iFHgxIArZhhN9qnBvK1LqtLocbG
okLQmUCXYWUK9vXfdAH7IoBiunA61UhZnc2W2gAzXn7j2pdRNHqdG2N2IMLD+SX4
9cOxzrbRLVawv4UXIFQF6r5tYhW2FfQsR9LNAigvftz6bISRrr5NHmJc8DA8byj0
LL40FWzTuyaUQWslYKX8th5Ia9rGdfekphqtZ+4YpcIp0ToHQg1wQweFPvC5OS8A
8QjbMPtI7ru8UfZShoEna0GqXeHl+fyOxwDKCiSwqhpsQuCG/2QRtvhuFR11iCXw
nYMq6WAsgoLtdfBW7OxRR1To8Zh0MUxpCxOIBHV8M2vIzDbKP+bJXQqlEay+V7bo
odtHArPzb42u2FP17U4coCqIX0FgMqhegnM6d0DdWtHOQFrKhQmg+0a0MrTPYoCQ
m+QAAV/CccAfJZfPmMO3e6LNJKd7bDMYHef4hU/EROYrUnejtc4J21W4HxZF8ZGI
/gz2O0C4Sk5qaHljtRZh9H+0EsOTTWafBRJEX22J55pyM+hF7ADa6sJiOk63URrA
i94ylacuF6QLYVB8tIIpxieQ2v6n37Q1kONyJBjtZ9IikLJGVQN7ucjHU35OQKgY
Zh4pfreFXHdl5KX7ulpXewbo2b+/4xQuOdTcFpYmRGIKChwDNkbbY+dJJ7hWfTqW
lLBHzfvs0JOcI8lsuC9BKv7pNf2gs18pNlHxE5Uc4dt1RWi54A6/yV5RrGIxy5/t
TOWykIJddUXoDuiF+y/XzD52MOsidqDoR8MbqmNc4fKKr1rYMI5Mt0r2URW72JiK
cEGr8/zownh+K1Ebtp5tRNUqvLSbYkpqK1GDXQKa9TzFf3CkSzdQgLIH8D8aYhq9
Dh2XBLtgEd7TLM7C4nmMlroTL+eLWfZIUuUKSCqqJnjG1tomSPTYjU+9iM1LPgVU
GQjakoyplzeSDVSPTYKEHSUtx5OgzadZaNjKRZI02HVdrF9+Mak0VufgTuVKNxGz
lCtBTqNwJrjYItoqnJ9cQ+vURvKRxiSbOeYMIF992Zc+ijSr4ScIXV0k6prjgy+E
Ml4QuhTEm2Lxp9MV8RAE7wPy/BkCj62K3xYoVyiDq8wmuftUxm74cxqoxkWfZMei
tEbuj+ooJqKCAsq6hsRW6uZRrB10+x/1hBFhEuM+io/9cAQnLD2/t4EftbzhTbxP
Z5pL7EXPfI5l2GzU+QUKMR1BsWoyWH+lmPhpBjEcqqHpV81rvQSU7Ax6alObUa2E
lLLCCNRKb52YFyysZfx1NHWdp0+/NEUXpJjkpSSegupyPYN5Y1T/xikqajpvbYco
/BofcoGp5pyqVTK2z+mSTUcMZiyowl1Ij/6qWvbijf15T5IriTKTBSw3UXY9nPfz
t2YGQNg5jw6RztqzwiKKigNGo/C7vPqCagmWT/J3Ev1oeULhmAg8nndlk6kT1Dvn
6Ki5vToAwgmrkYEIPyaFufe6cbHWbi/fjDYBYYV2rl/tawWt5mszabT0k/kcm/NL
OCorCGb/vHZ+OHlW0mzwcfO+9GChkkuhvwSymsCk8gvtUoL73T5iYdEIIKgpQL46
wGQXtCZ4T9R2COu+OyKDTphbCT0s8qYl1VuCIYWmf2CL0ZPinkHq/iBUIqo4QkEu
abFBVOceHrLBSZCCoEJasYRRJvGm3hFSy+xjBn9WqFiZ19ifyBjq9dRmDfZV45gz
PCkgS5hJRVdSOoyvgnC1B/t6CBsNh25KjV2pGiUJCxVCeVHTo5Pcw49xj1c6iRe2
RbUwBmYiWQzT6COmtwfH1IdJnT6XTc6GI39GLd0TLMt9S4J+D4tOmprbwznQbpK+
xu93NpU6ADvRhRe6ePKnyeUHmCR4jJJw3v0plyYSVfzH+qrnfaT9vyoXdIWYlAiZ
DhLWidFWM7vtOx1gM4OG92RZAhN8278OIK5YSsxhj9iuHThBeA5ZzjFdfMvy2yFq
j2y2NZYcAQny/fDXF4x8usTzt6U70hW1OqumYJP+RKyZqZ7XL13j+ZKYCh1RNkxP
AbXU/vZ+YBBdX4mwSqgGd0iMxSwHOI6IeeOIPHq1kNX4etlVS2gpqmhAVUvqa7jB
ncuLO+oV6j11doxtkBanITaPQVBE48zAeji+pxHby7FTCNv02tOTxdGrVFnNAHoK
oLsHEF6P72IefIpeQR3IqSRNbdWPjQjBMrKtW3FpVfUG3rqOXhb85H8vvfmum7xv
k/SrOr1k2RXGHGuoXvpya3w8x4HCaCmXMFumlVVj+GmuxxfQDtFmAXwh06tzIh65
F7TXnlNm/58orqfAtQ5+HXPI5Xa+8+YoXDhdZBEIxG9KYzUyo1LZnhuxVlzFTXG5
Jdvlkrkkjz8mBtq9zUSdmcYE6WpYmrBgDWL9wwoYyfOwoExtgKPm4edT6Mdrf6aO
aEsDEmKCfV+yHjAAs187tdqFmA2WmOiiyCXQMOTGqHWcmYaX7QTLQKMmpSm7i4h9
c3hDq14/cGM28tUPNd6rVn28zpUWoxWPL7o5e4NoZCwcaPbCPeHJeqnud4yZpQHA
VSoJh/TF+MQbRnIdReccGz+JmCNZ6Hcr8X/2I43T5yIQ3V9PdTM+NfMjWKstwDmY
HtSz0vdVU4yYw46gvBGN5L0dfJEMes8tKGzYdt102pR9oLaMfkAeXrcDRu7NnOrs
urSr649xbPQHJnJOyhI4yrVDAkDKcCqdjG333wKpPupo7q7blYKQGTRsz1SF39jh
eUd+SsoXjFYlm3C7qEUs0xOFWRCQ4iDe4UNGunRyNQjdVcsTd1jDDYyvNiDq9xll
7kD4/CU0j0zN5gDDnq76aC+62BVS7NBs85imaVG/WnihHNQ2zr3x3FCHn3xv3V/S
+qm/NJ2pgbUOJsd7LRAABVq/AIAtkBEsvzwUZk8xE+jW7qdmW40MlyrjXn1BpVZf
ssQjNRgR8VWAOZ+tBhgdPwDi9OZ05Hnd8c5XXxCvbZUDA3QIt1Vv4snEGXvecR+V
pTIibNZijC5EyBUehoH/bKY9RQ8rp+kAMeDdcDxsOke2kQ4asnmuVp0F6RZ0QPBs
uEV+2rfClgKAtWVRna3jlyrsAz+kEiWBXMbIKFmMRiVnhQ29kyb/VfNUVGhYq/hx
wDUDvgxVhXSoArotfSYq96iLW+/k0WjkrFw4VS2dKXm6WblkYyFYLQPM053oAv4v
Euj+BtAMjfhTuvUh/dM8/rsIgaRNgShEJ6gQUUQtE9Ssppa9VqvytMv2a6zF25lO
DHnh06N+ZkJHf8XmZGnBleKs2s2swzv++7V2lmzox5oWftf4UND/3UWCSvjuihU2
qMh7x3wXweyvMX6TGsbPuRvmxxDgnoN+QovH39/mL0vPVhnuUiZNho0DEGe3r20H
KqTaBKZgS/iVbcO8s5uNEFo46luAxADcfHaavvf8i+I3xvfnwhMeX764J1ucQK5V
jyDsV0ALJrsaNNkqqgBPjqg2gFBTaw3UbZHvaeofo6je78rWO5NjShULMHKQVLh9
kCqOnbBaTkLZWF9pb+/Rnb9nCj++AxmGHf2YoX4EsCNbVv/nqTha5j6ZpOG2dyk9
ksUKEDqDs7Osw0xypfZ+Hf0A1cB+y6hM5NksOmlHkNYhmbc1HdWaRu1pexQ7EtJG
nYagxeOEU4ndjne8rUa0A4aE3SjP4he5SyWmah4cY1q2SPtAjy5HszYSaMZZS1+4
tES03I9zY/amtu3a4t8mmTiT6iRUtKsAztXh8iqNDiAQx/gAbQzCaiI05fbD2HRQ
PAVaRYu9XoqQwvUMaYL6tQLjhEwHC2OpCSdn7lWhHJxzrkeIdsWev9yoiEXikiGQ
Yq7N6wIg4OublFNoNzTlHFohueYK32RvKkJJ7BMg91qjgdnrW2y0zl0mxS/qRrpZ
+9/6uZzjIMci8iUnw+/Kt7ofSHEbiShst7k/7VB11jm8c8Tu/HIm8dS8loQxi8Op
mEXKg82rojnhIDibnylkugNZw20g6P4AEYij9BS6nrrIFz8TFhNyqeBr9WbSY+eD
gk6CNgjk03OwlcqQZWwDKJQuZ0IGDrolq/9V0/qXQrWF6LmsVX9RWRam9wFQeCeT
pXMPKLJxp/dgD/i/OQCfEmhZsCS375up9NSFErAgcXKoYJYDDGyrH22l8bTgmeGv
EN+7LnHfaN6CUCNzZ8cIKyg/lTaT0A/Jc5JNFM2SOVjgW5v2hkwSRypiUYW5vrG5
3r+JFZkuAB3+a6W7k72tZ3aqDrcknHF9rLiJJPLbTOexQ0L1hXHJZGmm/KMvSnxj
Dv6AuUjtkN+WP4HbhrVHBnPSKN5s5Kwb7c8jvcfRZWns/UJZ6QUKgcPzHPJEPApT
zi+4v3qYaK8VKUStWyoNIE9OUbXh58WJVwBltfIaTxlgOJSh4MOKwAdaSJmgXQk9
8pqhys7cJ1vcoky6OhwMGRgocRZQ5yxeqMlZO+tLLIPqHmeqHW7GolTz/x4q6fJk
7wx0abFQhCI06tUtDZrxerwrzor5FcS2fFnoz7n1MGka9HjBk8fuhRg9KxewS4Lm
hJXxsB3r4SrHNVx1Efn2yfRINl2uQFZYiQzU9cfAa8fwDxj6x0Odigy6dZrmMdA0
lSqPVAjBkx9WgNgbnEt/kil7OznSlC2SJAIiuPFDPXs1Efv7MlxfS0XJl+DtcDmo
1UQxLTJXT7f98kcJubfPw98VnXBqJx5GON+xyeDZviW6xp/jS7IT5iOWUKE9exlQ
PUS+CRULp8+lJ1zqX67ZOJnqijbJ8pa3omJsuVy0zQ4Sco/OMFOGsNX6nyWiPf9Q
u/db6LQoN0N9t5VsW6FpLkHnc5Yf6jlhIpGKoE6a6s0CC79jmcwYooeBQ0/RLkpr
viTRqYY0nH8ixpiwfoweXpW6n2SlC9zddQGaSJXFHipSnxg7DUp+IXs3H98Bincs
Js3iHvB6gMA1KQ1o1HIK5j5NWbmu10sBTtj8wUUZP9eVg6HWJHCl599GgTzDY/QA
iJDiUJHiWmqA9MlP7qCVpYvB4yWPd3GrrDTGW8GvEV9cykU7BbqMCjRUYkBKnGb4
3j5Hnjw6UaUMuitx0oaa+su3zWaynJ1t4WLlPwBZTIsrmi7f5Gu5x+Gdyxt+tDZH
oMenPkCsqhAsFotpK1tHtvtPJXfq9/Ix54a+OTnyLq6ns3rsL57Yg5VmGGLb7D5c
PgA10g7TJbisx/30SXDHjkLlxDGZqcLjL7Hw4u0cTO6N0RuvFWtvGXRJRUPDyeQv
AmLX93PQ92D1jUnkfHqYDXY+NkevqxlrgbF3On5nKO91hqiZy6bu/xsSsPyeaJ8n
3jv1ukBQoUK6dCxU/uNFjynTvnbjCXb3sTUoVVBVMvG7mAnb+5/YKITljXdztJJ9
xaUTBtsdQjpfoJOYQM8eibEcStCKqTwbg04deb74gX63KiJ47OVNJaHJsm7PdZpt
BBaAM7nENf4w7PNF+o3vaDSG8Aln3EHwFg20Cs8NAe+gKMDIk4+LcStSt37f4/7G
3ZXuGocvjc3X4DnHBIhiMyEwCW+94POiULa7JHC52o2HY49E1iYOyBCoeVCBQmsD
3ujO016cq07Gkbiqmm3I5Eba48dIdblE7rGm1C65HONw2nsUF9vVZOimy9+4hLp5
7uEPIhYNr/nh2jUTrebrb4hHDsTkzHaHxb6ufjikhyGYuSdBrENg1wFLRRQHVjB4
txKKkmHCEbt9dM+nQG2ZaVpgAqVnlpztAXcVaShacWvxoO1baVsaGsdKvJprMJCu
LsXGHzVBW2YHHn+3FmBR7s3T423ZQG8hFdqo4hl8D92RLSIBjI6UwWdikkdRcT16
oXsSLkCQ9wwL1gkGL+5A0JVRckMYM5n6AhjF4t4FCUkrlWF2uyGiZDjcsB8kbtxx
dXt8+FcJ0YEZbYlPL1XQHTc4dUMMvQOGt01B+a6G6q1+KcNh10IxG4ariu5kMhK0
LzqrVg30XvNyDqFY4R9gmvsYCsLZ7PviZqv6pMbEzEZ3SOewrz/bz3dHSE/pqD5G
WelKsC+u0nJIsv+mC0/dUGt6DAJevjrR1Slap8Ifkt1ntx2F4u675jG9UK4oL8nt
QOD0sqMWWhAnVMld417fkAznwRhvSQK5SRgDT1ZR1dsOlbcCKA/hyrshge9MOj2R
HKvqHy4Q/6rXgiQEu0N0SddNTZligaz3oV+Qy1NLTlQ9Ccsp1Co60NTLlj9HJRMq
7UFdecTw++dZ3HsPG80cJhretW5c3vxTpeVdjd3Ed2kFZ7fmfyDzh8XwuoNAKac4
uUxK3XVCJjsnte8mtmiNDrhrc+0YVdYoBvrJgSWZEhUFjFErarCalkJfgjAmo+GN
7aODBrQVjJEJ9i2sd/yGR/HH6ENfdbhlExMvLXtqaIYQ9mQ+tnfjibKEBlNC4zGP
VTCAsDKMNWnqQHLGJz/XY83xo8YRS2j0JGoqGVhIYl6OGo0xCG4dKOwedQ4w3DOb
BBQ8/EPYxXmLXUy5GZZwclVW92HiqqFTT1LG4Vugx9QBh+BQLc8d/XMJCa5kOOmi
vaffrNROEPIkYebL1qQou53v9nfh+BLXj4tH8erv+/b3sThcwPLfxhXA1LvGnmGz
U1f37qHw4/k+55AAQXOapBkU36HZHWv5kYOIvhOyrk3zngI+3oZ3+yBysnHDirtZ
tWQ/DtRfcKrmdTmyki0NVys9h3ao6sv7P4NjbGWP5UmXuP7JpfUeAb4viXidTH3H
DMp+9J+KKJDt8aruOHROyRMkU+7w7z3yjxw7tlz8FrY7+9Eyt0I6wSLxK61u25cF
MWV6LV1AzTj9mYCFjUj5xYNynecyrgzOzcnxEH5K5KaY4G9vFjHIeynBjS1fzK2u
C5zn1q09mnJIEQ1sh6OEtrOxVtPqZ4X6KFuWeHpE+oUuqDXe9T0MMqvoNdK+tQUB
41J4X38DKOByrKTwZLc1OfWQvy1rThL313elceJsxENfXi5eybvmq976Njl9pqxj
MsX52VAY/cS1pi6kiI+4LRpkHrJbfqSrrWJzIeX8fE9brnUETalD5rRvKLZEKsvu
CMuB7iIvagvaVsxyJrYlqPKAos2uFdXOaj3jLNbzxWCmGdKRn4paXpTHoAkkAii1
VNGjdWZ0VCVqWudojC0IMFi90csBz8NcnNxXetE3d5B/z5LpSKWCRAclxjXtGhuu
34p9wjbh+97pQ1NA0SKgt9rc3aD+CXueAWK9guZPTfWHxEka/wIvtOusZRm0BZfv
HVhkQQLe6sjvPFD7RGPZCHS2dndk6dUYlrbhvW15cjUgTyDjIYttkQ8C3W0By5jJ
VFNhPN9sQjlSg5Xvj19nAI4jdCF5fWrRH+JJKuPuoO7C1B97fogG66E/06fJaA6q
I+wDuIeNivcSwnIfPKEXBy7a1GKwbWMFiwYMM1/A5Hl/QU9/Ze0aVtMh13AX+ldp
6Ps/pSGuhKqRFQJFpAQb9OmeTpMjR8zqGsDs882ktIp56Q2K77IdImlrY/znR5MA
2DHcdRo6034mrANJinfekWCTU+bU31WYvwHjPF6pxG5+/u+QPacu2wcXhymixgX5
pt/h2OqfIT6EaOic7h2i218PKdJN/bS5rG2ayVh+PqEd3M4nAZnbsOnxMaCLYxqR
ON75GF69w/3o+GOYztEfKxVbfY7n0LzzNNGypr4fuhp+/KIzhxJxpRyBDFMVLbSE
8EZcuRPYi5ge4Capwp7+jtCJQIH6GseLFC+EdrrVlkbk7UCuxkGp4AtRtEO5dDQV
GOTc6zPU4op/NLg6pvaJxdueq67MtqFgzqEIzZFxTPtBL3LlnXFWpcOP37NUPNQK
FV2y3Bu4+edel5k42Xk3BawiulDpDbzRuxA/u/X+P9Rq4/vDna9vzqGYRTzBo6lp
i3GQMf+2cWl3env56Au+vHOSGy/fU6a+rgVKA/LadFiO2O0/5b3t6tOg8i7NcpTj
ST+fQRgCT52SMjp9SxuV7xbC4g8DkHMk7ZnI8Hz+kR9vESNE0HDDUGrQxtjfpuJJ
KjSMOgn21sMnsyAVSUFPPFIDb3QRPmfSMF9zVZ3yu4iBMT3yrcBMCFaJTNTm64k/
HNudQRXGOvCDWOMbSJJ76ns+Hc8n66WCXI9MNhuY1uisO3wsNd+AjnyRET4L2SVt
6/1Ekn1HvOP/vq2qtNomQw50OqbOE94iX7Y/fSwbsT5Zlb0V9jcGf69L8vi4Y4+g
b5I3jKvSroV19pZGHFhFl1eow/BpWLL1ygWAJGzvFauGj1l6ucjYjcB9vqi2DUKJ
nk9lQvi4+BI30vuz/nmYLH1AgbHjs6YGnUvbc0aIeOq/nbMSuoY7JoFXYOQtA0I4
jK/TDU7PaGLYs0HzsJaAo44Dnl2d9uSPaR+MJJxtUAxtKn+jEG2UhU81kTCVj3Z9
06eTiSixpn9lQt/2oNU2zZLZA0iyy8dQRVapko55dmGzMCSeUYTONiDDuvTqqi0c
LHs23o1Q3f0YLkVE1Q5EOaGooaNkMum7w84oWIPm8ttMrRt1Pg+Dt6x1YMflDT9M
A6f/ZWgodcAlK7RuO/4XaZFbORV4scR9Bp4rmYzA/NP/ZSvlE5r8pOeXSZIyrVir
x+XxinOZI4D1dFPMylY/mD5C9LhrZ/gg0pAhNlIbu9jBHdQcFq/bAjJN6G310A/M
z3BiN+wfDjw1zqSsDasYpkXtsYyS076D4HIfBSnCk9K9je42JDRBZow7kSwJJj1G
BA/+mMXG6vjPoOifOlm/zpjMad3MV2SebZazB0d6JQ1qtYZA866qh4o3WZwAh0bs
ItoM4o/DEVUAm/2AzZ9T0Z4DM6DcxcFrc2Op4kLEb0V+YLtHMNAmfD56HWI0K2Tu
Rzpxjqvs9ZB6FZkISixsHMPxR3rPRJy6oDJZndamQUri6MzlQA/FprqR6RaN8Ay+
MpF4YEtaCLz+CzwxKCrLN7TYOsgs66oH8+i/VKIUuHWP3EPe6lC42F2I8gjsIGGz
cYBd24RtzBQApAoWRHgSUhCkq0aX/vunrrmInYzItmFUe+j+7xMPgDZEZ+Po1v5X
5G3MXirWJ7xH+nEET8nUtnLI4TMdJDErMMq7pdZQE5p7khVlaxF+Imy4yj43F2n2
182oz+qqPlfi+wecG/XqFGervKtkvFKBGAcCZLjz46OdsxmwE+qQscYrMA8c8Two
pzutzSeVRZvGyKcUk88iRBNjBP+LqJWu2StrQtLTecWAakAmOPzEDc9Sgt32qAMP
hU8frtZDLoF+JTQLF5VS07E4skpgJ6V7e9Bnocmd8FXqJxjyvAop/FsOhmXE5gyc
1FDdogewUfZUu/l9doinV5HOi2pNMxdrfIA81LubkerhSr5wQGQwPqvUcb6T9DWk
dd1Pcw8DN7bXt2nzXeRPJfBNhLtmHF0Ex7fgmq1gNAlV6TC3G4BZutiAbyQdFa9Q
G+nvBlui6emPon1SOaPzxVGtCH2TsdR/ERnjme2GuN+mixIMNFRVqOrqfoHzYXKZ
8Fu+oRcO5yI5sM1Z8C1HsyLSQklCY5L31Jvr4OE7gdhuLkhPhnJVGW/arOV3MyO1
AFJvTPXqHGPJWLOgViN8Qw+enfnBj3rpqr3tYX13hNxVqzpyIvS9wf8qhKXHMFFI
3+i8RzdUK61wF7pc670Jb9puTvvkXwEjjLdx3gN9P6dxZOLgYm42o7q21asZl4h2
Z7fUeSA5QYFp472EVHUf+ZNk4ieGKAWM7xMzC6Yd+fjZ0F4vUqNf6Rwgh23yJ/of
LWh5IEzPNC+I13Ox7zMovDjrTOrmHMoiIfK34/0JXGBJooa0dTvle+1rRNpl49zL
02rCzYCWRBrO9HSxpC5xnKVPVA5moBS12SUASnaSVZWO1gcyHeN5rJNjnaPp7JaX
AM7MFN4zA6HhPaFmk0QX6KLEKJrMAmD4j10xmCOO9nRVi7PoHEnBdcLTZWvlEPtC
mh+Myl7gSfufz1WntpeExamirn8mtFH/4eXwwMjeWQE9wNyrtFXYucNrjJuvCldp
glF59KtUUQfoA5O3jEALx0XXKSK6aSEbeeugU3PCZ0H98mRtyf0x7criSHiTz1US
dGkEd9v/tCJEvAn5DVCSq3qJ7rKsgrYNRV2ddivQTDjt1Ck0wGG/M7aQpbR/mvEs
rnJv7XaNCWgMLuwG2Uc0JhUXSmmyoEFo/JvMpkBl34d0nqAoetG3PMvcKv0jvSPi
3HPB+TXbpgAYOEO5DwDibPnzGxlFkd88mjwbj3DtFFIFetoe9Tm/Ub6TfXhrw2JA
e1Jav+MbzZgofjjMDlKcfpH5Jn8+HEFocYAcxDdebrwwaz18leS0UFoyNcv8BNtD
5OJfeaYp7n16Wlpcug6EQHRTDp/fkehYHAPV1fn7xPaZNLtNZTS7AAAwJ/9CXxgw
rlHoLyAuhh16aLOJB7HtUv+vZuFd34Q+9Wyq+kLnZjVKPtgO+PlGxoZzlaDd88XF
Nq2dEO0xKyVzxob7v7+W5YAPSR1T9Djq/bJG6L7rcHrMGuNIYThMPqkbD6wfghOp
2oVfVCwInmzVU7de2C/eV78oG0I/CBu1yySDfAu/0gbu6D9WU5NX+m1sKtYzvUJv
mIsLdhzcwkUDMbhXN57gCTZsHB9b8jw9hlFKgmvKzjMc8zob2ci0dLWVbHARIxfi
cFUhO2SHtBrvNsd7z4CQniDbbqjKdIRyOoho0cAX323VIUMXY55dYglSl9EbH8Hz
sjckUE9GI2EWbEdVToxx3gu/BBPD4rHG0un6vyN3bkU1+333o4vTY/gt9THrcYQI
JwuQVpaF3vm/we9KmPXONbtIBuE2i1qo07G3/8U2KmMy+mXCWjaVPTG3yAVkc67X
zkl4H2M2U0MAETKUO9t1PosKr+ekueLpyCZrJrNOu1NfE9fkN656g4H6w4ZMxA1E
dA08V1m+XLYSCGd4Em0ndNtmqom/H0/0GkA0m75y1kLm8O3DBaa9+QiLXsK1tvyW
i/DkXQrC8hHOE9PF6yG0TOagpA6ED4vewYEEKEHO+/fi7eGXPi6Eh05K+452y23w
NytdKUezud8/U5gdrnUx2tgzcWlowUpew5fhalKmo/pPbF8czc1MSoYhLw8MxmqS
C1UEQOtYjuRJV9BTVb6eogA+h+dnjuGR18gTnL0+NwBR03hohMicyAAn8WOoiWRi
iYipE4GdbpXEV8owkWmkV0RSCnBy10WKfI/kanQrMh7Sa8VlgIQMcaSURgBovVGb
nHPRY5MzuGDLXqOVWyhk6THwvPCMt6xo2GBbmpC7SNA28JWHdeQ8jK1VCcQggwRV
UPahvs8PdGv/fRGBulDCwBCuBj0j67gA8oiu7OZ8gB+I0PpK2iQd0BRWAZEebh54
WqeK1vlgL+3DcDYMQ2UckodaIZOdYEP4RNdBzPhal8NQiieyyTxo0sGIVDVfJzO3
YtdxS9JiZ4iuNnyWm2NhlnyQ2CpiKwfUAkGLN/boTT7AQn3YgQxfZcFRRaBxi/2t
iWqjkSvAlvpauuQK+V3IxyxPu9Hxv2L3+M0ZN4WLJ5Oy9rTIUQ8ri8o/3dqJgi5s
u40qW6ULZvwC393Ye51nwJVLX3rm+h1xrXKQrw45hj28/damgpX+Fsc+22I0gz31
Vol7QPSER9OanbfdSuxzw0s/qsElxCoSm07DGpVcwGwnWLKlt1lHm3jEPj/lc+tG
i83jY2R19JON7zTrJNxcgcwdO3kf5d/tUz9n5PydeUViDJTIUIX/dShL8F1ZkRur
bQcQy770HwIM+OYlmAoxP1o8t80CZZxzpEu0XifIeFsHJ+6B41A9Ilf84ArJNRBw
bXV2onYIONvOh+0NEDQtouay5ORLZAjrD0nfCrC8z3TszqsptUtfVUUm5R5UWsvQ
3oACVjWyt4SNXkqhV2Wgjfzr7xbMwsbwa4WINKSmbybpB5aR1N6DLfexwKFJ4d54
uhKs/GU8Vo54o4J6Be7K3qi+hYVRdi7bJ44wc3GLhQbTZPCGbwfI2n8gGAAdGZb5
E3rrEcJXyFcZ4EbQWylqSfUHRbmI+ZtzTTBQcf7P1GPm+U9j15sIAhbZiUTdlwX0
eKwwjlBZ6dLU6FVOokItWKW6syn2T+a/O6gnHDcJDvv5ZadWKG1d46TTHPVl7mr2
m+xnv93JiRhy1xlBoehoVDWuS8nlMoQe3Bqb5BM7E7zbRrMV5pl+VbtoDgc/IZyJ
ILv46N8mVcHD/WHVP8tJpeV3m9Syz+METUDXvcAno8wb5rNOYg4bcTAoKc4twK8T
eXs7NvdR1cJYUC6pduj8LTuM3RW5rwsVNh0dD6TYsV2nKW9s2gy2wEKlpE+4Xp3l
mx9rMSkTR6biLJ9BFzEJ2z0Fi7m9XKbXb1ZsG3Dn4unIN5UjkWFvkP4OzEjShgFG
xkfb2ZVI7K+RYKg0uY5n8Toe5aTnwkJPLuAjCTIA3cq9dSTQcjGWyJD54Zamx5im
sasOl9sZrsWZ61q5P4/fRpCgx0KeaJlFkNEuvulsJzfDWLd0t8ayx5tfwPJn8mL4
/nLm9MeQaf7cqklcdPfi6ss/1HuRH9SFMxG1E/WN9uNrCr3ZyhkYXXgE0JG4Y3M7
8Jph7ewY47bZMRemj+M9f8LTZU81YXsy40pnS+t3Ff5b6zuliceAcdNiKwPj1D5p
LsGB4oX20r92U7aTdQPyLz7qzuklGnm/AYmytafdpcIQBeQL6VmEqAUmukXmk543
Bi5VtO++QxgqPldgHiR1WwsqIpADPoaMbRFkof0fD1ndG1oCfIaEGExBj2TOZup7
6YCgXFMeNIeooPF8AOz1spaFgbeyls53HzQdr6TH22NSJwRa4UKlDFlsgJsJ9LgV
0T8ukByNxLtUKz3jUrsjlnnpU9C11RqvNAlgdqGpkco7pm8U5Z0JMcwb8kbVAIk8
ZAkA5GoSN5qGUkPXjJ6xsagkeEOswCAjPwUhJ8v9oOEuy12fo4Tef/CX4BJaQv1q
+ZdWU0kYpRwXWdVHWO13zy7ZIMtjNXDC0ZECExoO52P1XGS7rj8FTBixo3YJ9q1u
k9eHqJGZZJXMnk+UvUu9xzFvMUJfdVsxUVyWMdZXF8edqs8xDzrEq0dJ2AMBfWWy
5ZQNtZheYOgoi9H1Rbd1Vg6GJaHcUNWWZE7B9jaL3gqfbRtMUL+aMSVi+m4ecYqa
3L8Oe1Cz/l/RXMmTGo+zdHmrlKrEFOsqO3qIGHn6fY3YKlhAlg9Q0O0wVgTqabUY
gqwfB/a9keuVaLr+oNwVViJ4vULGEFcDOxB9cTiVx0QkBFUgW5mDMtY2dOXmRZgO
AFa1KHLKmlnN4dG+5Jtn5JuUojx3eNmEys9qN54hPVu9GUHZdXYtxSoHTyG9AcNo
COajPlbohnRkYLVQZXNIon2y1prnyh0+DGw5+C/v02DXeON4fEY9Eg8C31Kx4KlI
LKm/HqAORYqV8k/rUM9Z76ki/6UuWaPhQw5NvzakxTOp63gKgbeEW4ZxpYBOeqrB
hNHAoH8LOvRdpz2CHJhTynlqNuVQHyw4CjrgZccHNizIxhcrztA472V7CCnGdxWH
1TxNMa3hl6qxYqtZammjXD8Kux+LOMCK20TL6n/ssLPTTsTv4sIvy7mTUrGRHXXB
vJBn3R61oBPRZ0YR8ePGLyMYs4Ol6GOVIyrAyF/O4mJbsV+nCnjFwKGJIqHfoc0S
xVflSy+LCYDao3RoeF513xAw2nwcEpfJc9UMwsMrUzkFEvLt3QR0SB6ywp0d3Aaw
DMFAS+ePioct9wzgF/468j/tRw5AZnOx41Z3Gx4bX+w8XDwnR0RsB1tJIiFMC2Wy
ysF7xNIhbtJEqAsHXw3xRD+UCQ7940GYXpANZBWMYyVkDzXzoav3jPaJu0RqCxde
XxjIl2BvmoAbM4rf8JJ3APCs3qwVjfzuYGzR+pmf/G1oRSZNBUbvwek2WpWzXzPI
jv0Dse/4YDHlpqBlRBZGdgee+eOBnsfdYzIXLWKYqJTcvD1S/OkIMk8ti3ciPkVg
kYj/2SSOfbWHcGjm84eIPH4JiKumdFig6SXWICm/lBv9fNeypzPJP6mMsRVPyGiJ
ysVf5Zag5YOzHV5T0RRsMRJn+TnHj37ncDvaph3qnbKXOdggDZDj1d6xc8ZwHFzg
xjPNwvjObBR0Prkkz9e7exFsit6sVjWKnnq2+a2xt+knVyCDmplXT4NqUPPP9m2z
LyGxGPnWG5Gjxdv6HtppIiGBROJUr30hA8LvvqRICJvQ6qZzr4b233sL/sk5R8gF
gBRZjNvBmvf9g/IguxBSbSQHrzJ/L0v1tvGg0w+ozvvaIbP5R3Q5XkZGwdoPj1g4
q4y7dK76wyxtmCJJcBPdFqZTn5qiqTJMIaI6EaVDUBMZ9RrZoYLXty4nPweOgK/K
pHZcN31iwGVTVch92Lpliw9CRVDL4auhp414tDAFwLETF4AIj2aVZivfjrRI2k2D
U9jxJUayrksgaaZJao2+8dAs4qeLY80orFhRVGKiwG6NoIPVdVOrSO8b1VIXkyYE
JN1dd0XLYDyuCbuRjIw3KtiJ4zqcRPGDGy6+0P+ysPO0PThKl0nNDuaORZSKx8Tg
cc/ZCnYRHv41g8rJqjE/7gJ3LI+lN7eKLXh8sMfNCbJMu8hHbImqS8QLLLSikWsp
LgnC4Jp3FhUDhJ6x2OfcBvOd5+ryQEOp7pBZ5F+OrgZA/8o3yo+NlbW+4b1Lw23F
13Uw7lI0ZOE9KA/mu9F0NJGWBsDg/cpu0HtsEwwnor1B81s4GTyNsOnTsKDuSq2H
YQMytHMGAgSKHqgUzWUFRdPdPubz9/7wZuZFowAF7MsqgbeSnpvd/+WK2hOriw4M
DX1/0uff91Cy4Uhq8uRn0Seqzgfj72geoPSTN5N2lt/DVHy/NggLkgGNtQhHY37H
x92Jl+1XFQSd7Y5bDQnj+YyDw9YLA6zlWu+q3kQlP5QBxtuT80OsIzRSi314kmw0
gx3l7K3u6Tsab03HYpQL2efFB8T0mBb/vjcAqU3jEEiJXLu6DUKMCzFtBepVRGCt
BVbnnhXNBlxyotN9rVTB7zvcQFFh4UycRY9v6xrLcRTVS8DoFA8dUHb1jUpQlG8c
lx/GHY4aKbBieddtbeVb6bOcSvYrTJDHPTEMYMtHjZ8onjiV/oa0uggEniqGv1Vn
BDUrmKNg2EDzR7OapmT4/4U2nKLQV5+8deVPQDtSbjtUp0d2qRWblljpToaQr/do
XkGBclMbpA8ui/DBnKK/xhApjWgP5aWKS+lCdAShHOiZpO2ZQS+L/gP0Dmu1RuE6
4fLpKruZgfDkpD5XpSh6JHx1cIc79vEPGywCimmcNTm8NgOy96Bt0tv3S25Ks8+i
y8itID/RnjH1dYup7GfmWLfy5UUH71+3YmRNW76EVP3wF9uaYFexx+5IEcJ4e8S7
RrAejnPNgpErpoyAk0UHs2LKRUrg2UBe48gzCJsisdtsIt+r39v9GhToCn3WZXPQ
mrQ133NtfHJLouezltjNMLaIBf4L4TfbNc5tjL/8xaHUQFIfJGTXTxmPqf8//yD4
uMSA3Z2ZGB0ERWMHpdPYpRhzfTemGZ2gaYll/e+R/dqKHaVFqKY1YWxiHJs/rGts
kcRI0seVb8fz9In6+4Sb2NFTHZyhwZn3Hlo9ZFhU1c//ONvrxEPgaPJ2k7Heb2aw
enLipKJWUlLNMv3WrJSxR9qua9SxIMWdOoPf1Jc3XgTeY4mkNE4+uJkM4A3/hSPb
SlIZ3Hw3CxDylEO1Yyh0X4rMjdsJSi0Q6jjemBoc8rK1ViH80SsBamSOyouEx+zg
Q7ej6eGefFokh+AH0fKtqm18RIxSly05/zhh6xpxrampqJjnJcHILBXHQE7tHy25
92LpiPYFsZWc6UnJfcVAfG5JUUvm42XEz2zOay0h6YUdgBVta2N04iNBd/EQp0Ys
QeTmN89rmCryRxxKhjO5Pf/8E9AjDF1TA46xLaou4OL1dCNZpCWjH+UuWKgBL1Bh
hcE4+l3DU2T5ak7QmeUKcuJrmgn0Ak2dV7145VeBDxGfrogrQRm5SzyK1m6U2fJC
YdIIc30ZdGKyP4ZY1gbgNxbmSm1Tyqg75QleCUIqkA60nOPQGdC37DTyXKUmnieB
MEOz7GuZvI6YV3OnWCSa9wN3GItOgYm2XaTqZwLymCI+Fm67x1PLbb4SMViKvf/M
jD34IA4Yw18L8HJSw7UkiFOF2Vnjz5OVfTmCRZUmuhZz0rMjp7fOiiQPjDAylVzV
8maiXfxnCRD941bR3/mOLWkoEIlmfFgym3WZMUtPEMGMEd7dja+uB2w79Mr2ifBS
2/n1CtLnDC19uDSuOOb49q6C8ViMuZVXmMpWB1jtKhw7QQdFP3Zunow6EnnFi9BA
b/WtxdnOVfUOALwK8y/zwQ2K3MDqpH5Dc4eBZTf7kjxxC3oCUJrczyr/TuScHxyl
0M4R7v60joDxGtqigNHoeS4BY8Ot2Qjeb/dMJ/7ymN+2pHQCVCH85OqOmGGhWLLF
KcljCqsQ9zG7ZTVxm2Gufdq3OYhlVcp9azXpXHzkpXoPQxeKluqEEFUzVQlsNuw2
AoUwAhruDpL2XKx3MzwFT1fKv0u0NcSJEn84pGijTESXA4D68CiSRyqfaEUMd5BS
ri4mxXWNy49LM2k+fxff6u+Ajde+mCD0Dnro9xc2HmwWP18amLotyrbB7R5gl56G
+GY0UExfRD0edaIbIL78h520u95QW0uQB0s+KkeczntrWDm1G7vaw3nxPOSjcSk/
L8tTZp5/GSymRE0Cfl7UqY6fM/V8x3oM5j0y7vq/I2lU8TlU6TeQt4qhwMHvR/h6
HMPwA4Mqji+0EmCGRYRbIeDH0K0R8f0mGVlgSEkGPss3XIuXqZpJK2S/u2EF2MLz
0CBr4SS9mhkVEHOk4P0FFOK9rY6IaC/lzTkVPd+vxO2MjBDKELnSCpvER7FN9YHs
07sPeyg3xodXxgkxg1yvHlj+DFBI7AoSY8pUchfHu80+mMQ+76DKBIgzaxciiVpr
Xr5Nyd4HYxDx7oX9nf5/kiZLjGIVrr8Q0ixzQI0yH5MR0X4E7WL6nkVh3MffJRn1
GkjE5SnKbdaBjUjhG+C07RE/B3nk4HZdJy0ZCqUxLIu7a7L+cTAYAE6GwBM3kcAs
LBgbhj5HzsYsL8cPlYzeGga/claDIR1HODcshY+0svwLnLMNvyxDq+mEnXkFG4EU
9Pjvzb9XsEA1CXsy+mlE4+44APNZ3kaPgsOuJ6Qnh/jbFT2XjOR1pjik4xNmQiVs
Cu7R1SYrC3NC+3al3oJ8n+JJvdDB4uJnRtRk16E+eG/mI1naoqDvfhuxTx5Nx0ZJ
8kzjgY13LeONRRkW066VdXVPUaJNyX/LfkaXTbSij3kVzgSZLq54On00HsUk0nG7
vDzClAMRl2Ao4tdkDhMqpauZn3zPjEUjC9Fy0ig9CleydNmS7jD7a3RVjKZcnDsZ
dwvbGOUOBtiyf5UOO1hFd0iT7GEzYCMqrccANJbyk0SQi8lwE/xvTt8/vw4wnkCk
BuKJYpSvRVHgLsQyNQPqTGf+ixZ5N1w1IkPo7qynonz7Ju1hzBmaoNJprgLhER3b
L8r5M48BlqMLRUutM16aCulCyUmQpGJA4NlNSA1Nm0JubGdYr/6r+RpnED6cE+Vb
JrJvLsgg2rTzQEvAyhoOxxYB2Yp7i+NRo8AvNeJtuHgUF9TI2vIOkX7oLt2O2lhb
jUaPDllZ7rutl1oRHVa6SVkjbNV1Rkfg8YXRTZQX6MvdsTRrHjKop5P9+Is405sh
n3BiOCBhDCJkxrB62tlC+uteesUZ2BqntsKYHla+GL+YqogcwLGhZ5n1awZ+gDF+
8AVsGfIJsq8F+C1r40HtulFeghWfOW6t4eFF70l1QCkeXD0b5cfxv69e1F0tjVdT
u7h5tWqHMwXrRmrLXJMLshq6FBWMavgMaZH5Pf+pqkE1OP5Opl7RMALzQ2SwQgJf
+3PHU0gNJ6QZnFj5mMBaV0wfnpPkDAHpYV0VVOXXw/jDYa9keEkwFFeHEXQF1WWq
zhU0947OtzFgQ02tSZsUDnsUA0iN+QrfeDxkyjciTJC3O+qleH7mcggcM7XtIONx
wHT5JZhTPbvfLkYJdMTPqgqjGdau4RugKXLJOf+CV4G9/xNw8fiUgDdzu3OBp8/j
kD2OTIU4s78IzJuvrs1E+oqe3SBs1jbm5cfig/dG2GRWkuhIy9eznfHseZ1XsYMs
eACZ05MECw54t9UywthGj/IMpuavW04lbUtVzvgQe3da/kCoqEa2QakKj2DOvvXk
Gk5aQDkNKbFG/h8TnkrpcjVal4RElxa5S5NSMI90IbIrP0opPOnL5pwXtb7hVTNZ
2Lljh6vfW9WErYQEXVNzi9GmLBp/KpUEkPM6bi8RZeRo5vEwjF5M7gUFugIokS++
bjFhQmRUYGhJlfOhscLh29ncAY06TL6T+zgXtFXYnRwIAIRREiBjO6t5QlxPM5su
60pMYxO2hY4BBsVN3GGINMgyEqwu4M9FC7QE3QHM5qX0ao+NdkPGWqQVhsN9OSy1
EF0zF5N0whN6INkYgSo93QkIgUGM/P/8GgaR2iwMXv0DXTwcAoLtKl1nuQGMR4Kj
S5GOrIXhkvzJNRjEBl5J/cgOCIQ+uzfIKXCof5pu89Od8YNkuYDHdCl4WBshnBKV
oEoTM058EkWYoEEr96HLpJHGHVb35CF9D8+6ks8k+aPu/85OE1A8QQRkBKFkgZhT
WFDFJeXQR4yKWuj2sFLdwG6Mn5arUAhmTKIaZM+CF/8c+ihOMwCWaKYPDGHJ5Dw7
0H3knfpR5B3wn6yVlo0nMtoVW5Njv846lR9PedouVR4DYdKLentgTvtISor6BhGs
eMWBNQLoCOOa9tj+tPNu3lVYWSBkglDqc/nFtEgu8BeNwI5ipbw+PoVA70o42vQr
vBG79JM4LiYyjUlBokwwjcXWwysAStGRi18O4DY+A9EFSL1nfpXZzkuyxuSi1na/
ctEnPGoNKVubHLa7ENmsrwXR2nv5tM1ylCRs9TJYKgvLc0ED42VKqr465VBLtWCL
Ri3v736mFxfSg/jniHfqd0lChZVrcQNwqJaVC5758pKpfawrKy49AGydapiy1PzT
xy7H1BrQgC5ACtq1TI+FeSLe7e4zajfmmh+gSB5T7/cCn9pDdDCs5eeRuxumx4Iz
02nj544thSpQIkiiGnb4Vp8jVbB8WiOTTY28dqzOck6Jxmmb0ct4DoD+2ptLcAv2
2j/fRPC3xGtdV5OGAT7mkvQUqgIDyYMkpqJsr11QHU7pSDePMPEiJ38QM1bWJcnE
PNrpW9DsRV6U6wy6qnbMqdG+H/evJ8DhTqNp2t6kOTIpWsMQJBBvBaNjtxc86GNP
YinTi9R5JFPVjYmGas9rXYmIM8PmeflFUzhXsCeshBM9Wnr7lHJpRyPM+vujDkDz
EvD6S8yvI0GSO+3lVbk30srDJOQUq6NvtoZbYPxM2jZPY60DMTTZE7VZ69PiD2S6
5K7WDCWtVQCN6chyun9wcB+ISvpiVDpP4sRUFLvXyzecfKyh1KNl1oxuFOteTNhD
5ijCKsLOn/AbNbBlSVOeS3D/2QqoU/0qiKG4uzpQhbxACXjRNF1MrJkHafb9Yavd
NK+qM4MNWboDRlt9/LgNDiL9WEXNrvj3xY8rYiMJ00wPG6FOA51pMYuCvZNhTsPS
m9l9VuCoTA+IhBUX6yczTq2bgzXU+rZ8kOGPHvRzhPOFymMw86OqP1cmZFduYYJI
H3db6nXrxMAxqQTwafEaoATNTxGyHjOiq8A97Y6m5y0h28clT287Be2WAWDpUBRX
XHF8lgVCtjwMZ4MAcWCnKjnwf+OXzLae1CkqnsR719t9Ogb/5kON+GFwaK0g8iXD
7pUCRXRIUubTXP1sewbXBAmv1jK4R4o1iSXriti06a+GW0JvJClK4CzFOPYPRW9A
MjMAfgGGdTRQZRHnj/x3qGb95kHvU0Dkfdp/K6wwhSOkkMIL9no3ZOJHxorXqIPS
+hEFYVuFyai57t9dg3ZCQmWiblIUsslTwQ0xE+muNzygYT8IwhCxNQQyfDT0/Wmy
+n+QbgnmVnBK2sIE0eUxKjVPJgBDYwulIFrCFLm1YWF+zW/z+ZLhMiYPWNd4drGu
UKqm6n1WVLF13YbW9MBx5IbmGwZrTEBUHUgf+cvj9bnybMwJ6qEe8JdsiTmjcOaJ
g9SjYZhANB6CskgzlaPn+S7wQ+U366fpe+zGLDWYWmvjOQ8P+d8US1KTpvggo2lM
4pw0/ZnrkIrLzFY+NMa6vMCNCd2sqe/ZH/U7IZazwzdfBdw9tNMz2i5Sjhvpya+C
oz+1Y/QZJdCRiTtxxXPDk1IWhXSkDm60jKv0b8GtPNCCYSQ/daehAQGF0qG4W3dq
vuAsVGHD5Y9g2C0G8OI7nVP5dcawfqSjAhwdBymuvt+YXI9RQ3PsMghmNquZzIyd
1Plcbcc14sp1JGSqfXC7Xbg07vc5bHUn7IrCpco6KAh8eH9dvWU1QErFsXZicmvy
YzperIc/0I4MA0SoVA/+FZjO+PONEi467yTkeQ2sYX6CAONGMjBdQOia4FGK1YjB
V/wnQhsSSEmCJjzmsRY2NQfStddqhgpr9ZdRZbWR/TYN6clzNSo7rb+KyU8sgoob
rghOoeQ3iQCRGWpxVfRfsfT+8Q+jfb9bN/Zi9UZP+K+2Vo4I5yqOteei621lcMIp
TACV8R4WN8VojgzqcskSTloDc/r5QaPLjt5q5LjT53i/MRXubjEChfLe9zo7Ziul
WbmXvDvVO6y0+SjbpyLUA9gaqtaxLeL+rCOhmrj4E8wOSsi1o5rEYrLaZwhEU4VL
VuL+ZM4v+HMXol7yib8aK/CofEcwC0x4qDbxytI1QYf8etVlqhWo4/khVj2Zfsm5
HNugWq0Ygo1uuYFw6bSDVtU9TwIBHYUwwCrLHFzF7xFZoScoSwQ/y9UF5ByxtcfE
UmA+HHZuURqpGpD59JKy7J1lyoudlUnraCr9Vxgke0OtuQd1/Tb3vqaWrJd5vjKd
TnrESzY3KPX0rh5CF8G82qBeLLnjuMP0CXkJpAWLRClkwXNosTcJThXfK5HgLdmS
aJFgvhjzlHUuZxG1NhEpiPE51QUcbCMmYs6iLU22SHnr34YKN5zvqIbKfuPVOJfj
39a3WQ0ryFlPhobfRvbElZOH1qcQQnQcpyXZaPaKqae6+PvgRwNYAJuSvaaLSIn0
6GCYK2c9wLPLRCzkpK04pcSSuWC7cLW++49oRfZxFBWqNXeGwW5AJ9fg4BRB2ToM
NggqjqXWFGnKenGYWs8DFXNOzE2BjSrCGypWCk8EnlE7ChvJQZiTH8dHQYYcaSlO
rUyZHwYc06Kvb1ibbZ5HGLgmPz2/iXRrj++Lr1k7TJozWFMKNWTLurjqD3VAuMxY
E/qjcN+cn/CGCzoTFMvQCS7cHygXFbn6+1HqellJQaB9I8zk3CqENgjIkuoTvmuv
IWYuLJZgA6EQLgTqsLKlwXi20p8MYIetNMxNuG0ZorlI0YTQcGQ/+QdGyja9Zy8m
WamUeOjVtVBfVEqhpi4W4Mu68CU/iLVnn74Rha/o3wMP9Lh6VXAzlVAlX8W96S4V
cQ6qfGqFDYWoaYIlhVnVowFDTWsqZhjmgJpEiuVMUfNgzTQZdFV84jjm0iA7wIBs
AL4xwSqP4fQqI4AvUTDS7whYycb9YfVQ+A3ZHuRLrc4AsWKbXyl6gWkSqg23lKVM
8K2O3BwlloFYvJsziTeAE74gs9egowUbIWNIk99PImxM/IXjixNCBPQr5FwPzsUz
eqZyvNE2mMO7JxuHG/VqLlKeDPBUzV28UZR5b8w012lM+xLM9gmxjkbuVnQ1uRKM
6Th50py6EezE0JqrZDdo2UfFdCO8fWOj6dQkS+BI6KqGgb0RKcwSrWbVjof7dr27
9Fb/ZejZz8Nnvq0isx4fkppJZ6mh+6DIg/3odTT3dECTWeGQd62pZ3lkCSAx+y0E
o3UYBiZvN9tYCD7DKxgRIx6L/v7W5ZjzYpvzjBGCW5F2FNd2pxClwCF3wCu/Ev8x
hMRAyod9LZ3xlb9I/+yZMbiGw+dONByTmUh118hH6cE8dCDFpC7Knld4Qajea5/y
CTnINfFWjBTPO2BYlNceGvMhUjoKYloIFPzQS0JShnxkGfl+iRZqDgvJBljte2rE
6twAXGvJl9FHpwggVIeuQ6drSsZZegqnP/Ky/H4V/zwACpGXP3jlfcoTIicV8tmE
mQxLkP/OApLYgg2eO1khKaRjb/rysV/Z38bBd/L8SUaj1wT61HSAZu5bly2OjXlm
BIEeSHOEMz8NLsVeF7SguxeMDBDbrC9/oaf2B5JX0o/1d4PSkcNPWZq+sm+Ef6B+
6pdmkKDco6WfY0mud1dKuBjx1QsloE0xbT11MtkRC6+1plA4CaPkKJXDm2n9cjyq
KROiSPE17I4rnjDgvrBzkTMwVFi6jV4DNk1JOly56PBUSuX9gbUGUN8ot4XMufv8
ix5fYuYuxs1YB4xil0PyUiCXFCJtqDwrlG6f2jyj5BbMLO9pxnhcK1925IGCt7o2
HcNKttTwkSYcwR+JZ2gS7L/jJidz5advXnD6p8dRNf8o+ziiXR2fStXX1HBvz4UJ
p9VjNZkDu/YO1Emmxa9Sd6Mh2o0tqibZSHL8rPe8OGudWC6EuyetKd9l41Ht3u6T
LLsB32T9FleJRQCxljXITXDqHa0Zymqo97JCa0RGqNa76dqBKQMjyINlaaOjqAel
aT6lUZouKmPpRRClN0gaoMV8ygjH1gw+uSkq2izL5o0Ur8+SAR99Kwnb8RfgEou5
4h2brMiDEcTr/PntECURulelg5ZDcEoDb0WuV81poLC0dZdvRMWJNUNZstr6thWV
xdf4ibFHzEcPOwRGImI1Y47rrQjSlz92LPrp0/XS5TxnkPpIu3d88yWA63XpCGlz
kCgKKXs96Oo1XcCAUSwXnmRCcUsTzwUpD93xFf/7Dp0RxTsjV42IOWIZI+7frejY
nrdC/CFjl8bwEHz/7f4irDXfUoUxpM3UhF/a6FAkKTS1RTKPNRbMsRRB4gIrW8Cr
1QOppB8Be2VZzMXcgkib0I1X+DbSCtz3kFk/PB3xZWIbiwy7FREfUjURYE4WWRna
gIAw4MxnxZhBqif9O+h9xsfM7K8QFe/XjHXiGl87Cdw14uibnpum6QuVoMsXh7Gm
IgacaPMMzQHCm2VBi+GQZ8fwxK8Zh41mC3gK9lf2wS1ZtEpVl7Mki63Zmnq75vSJ
xaj8Z7kltB6igd0L2H3VRULzprYES0/5cI79ecCHxZ+yWxCrmtopgk0NQ5+Oa/DE
apdU8LulQeHu+H8SxCuXLqwzYDQ+AjiS07uZ5hUu1JHL7apCmaJ9xEo5SZCyQwzG
pnQaSSMEXJIGJlvSmvIX/o0vOjyhfdxje/UNm7OR7iOAlGe6uyi1Q4TDf/N4UoNI
1lyK+4CGPwlWdgYsBs7q4GKM3Fgk29f1BTMXpaZC33oC3IsBar73Rp/FvXkpGA7B
PcvcoOdc9C7WdBvN84nltlLJeltHvQu+SlaJ2iTGDph9zBUpDIRU84YZItMJCLkI
cCLXEOLBBSHtSpip3725L/PIsQiYhbf14oeTkgMMkU/1m8GzMneviJ9OZwxAjLOe
XhlQ2/Cdt/INdCmcejlmILFXpMeKxSklpmg9tBwuGEF8roxmxNa/eLviR4nd5ADd
epl+tJh3MDIZgdbpRIwfId7goBpInuGPgANSo/sWZeuh5NP/lw3ufn9EHXkg0q04
POsX0J6rQRnDB2e0UtHqmWSI2S3mMjvAsP5GZN0hK6Pp8Xj7sRafulS5f4tsRa0n
/vwnOVdLd6bf6/k3o2TT2y5Y7w7BwzUUpIXyhBBsj6zM186qtNgR2Oz7p8ciV3jr
nmCsG0a2VDZQtYfOt/C0Yqc90+IofMl2++PtF+UYXYE12ZT5A7ikcfaiaiUm+tau
r9/HRbIe4HBFISsUA1VwuhP1O/dLZHxpbPTUYwyTgiQZj6lvTh21yfbmJszUpF0i
FqWaM9iZqdUlo8xsaQsdbjNPmDoFHbZCuh1C/YUpXH2wMrh5m46xk1SPQRpW9rDh
Kpyj1sX0m/d/xPUtGDxB1cQK3a1+czTFfSS2Ke414Rk5gsixuT7wiliegt8Batw7
Nt/5ml9JuGEdGttC1yrQjSMHeukozElOB8BOjqtKS4g+azxm0Yie8fNcAYOjzeIl
hgE+c2gEUv1PiN6USuyz+TW/lijSrh59ZgtGTicWwIGrArbhowQYZbbOBjQUPN0N
DGXFIdw6Sf4qr3CYnlfTPEmhoQDIJHYG/RBZWbRpV5HXna9ETZGXxwg8CekYr8JN
nNPtth/wmb/WTmryhYpygfYMkWbtALKFflzQ9X8uuTji27+P6riK/J3yHbIjfuHp
kL56boEOWzQXXDputGNr4+epj5/yY4oKelDat8ehJEc=

`pragma protect end_protected
