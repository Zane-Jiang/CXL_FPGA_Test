// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eaodEnH0rlD4oTLPeXLOx3zBmZi7tRNmspKRWFvA728IoouqJCVny5pSoFNm
y4swQ8YLkWp1yunTevwqfgo7iXhTggO6nj4npNtE8FrDy5YdXwGGJWKznzco
6d07DYeNvjBxdfE9gsyJQTegP5Y65ozqRmaBfQrW0MZ5dilfRWhVxt9RhZlX
gYZkA2PQ2Gz6BnYTqq4m2PxuUPpsQdP+MeF9RWnHS8bcqiqgSYtMBM8Js/R/
EV1DciIdl0BzVo3MTq8N5CJyrdPN1aLlp+cTrM8Zo+sq6pm6fwgIV0ksdNzs
Ufs8RjsLrDZrs0mYuMjfokF+A9FtANzOoEd1sAjgrw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FKT2lEQkwS/YDQSYl3KyINfKghZgIpjV/dbmS7gJLNAHxHPq1vGK5YZNND5s
K4pBePgpjjB7H9CE1MWR6zzP4hokYACe4+ocD5HGrTY8Ye8Tnv1B89/Qq+b1
GUKO0mKG+TOTpLOds8HqkNp3XmHJtACpZvmir0g36JRvkIJ2wHyxgHnJzDgJ
EfuVUof3MLgPAWzxX1ENNotsbpsxIL4XS8h37ynEYYfW2IUoexVQia+0VYIR
ctsoFt3iUKHSTuxUANjDXMIrHraxKX4f0+riFRpTjQX5tvzU8WZi+a34A1zx
3jDqTLfisP36R/803AAAKXctjHbe5Lnjv13LaiJ9oA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kyvdthcwq3Z+9pHeUm6Hjp0qQPngpDR+C9JiZGHzXgXfNgi5hzpDRsLbVi54
HejGkRjv9Md6c8dd0wOew3IZfB8aYVxl+zyFdnIibUUo5IBn1lsxvrx0BQAf
+kDYXefAyWjznqpZQ8sWYzryjUyZmzOyB3+Vz/2sVpN4Zd/5o+fSJbLtDGhu
C2//MxupyWIIKtpHrkpeWON6QrMzOlMlQUFV+Diez+HOm3FIUgiD+hxrZu4z
AyYHDzliaa0r1m91hnPvTddvwKqdPZuLf4ghNdoBqG/Re01DIpafIOEC9T+g
Yb9PuLHtOlh8L6UX8gQ2coc8bNIXgl8ytdW7E4LNbQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Dh27XLBAPn1KY2EIEQQ/Adajl7WKGXP0moSgU/wE7/aTi6QHD0pb8uStpQQP
H9oGgXmLYeUKUBk3hE91RmCJ5TVaEvVLyP9MFbX4iL89ZUSW7C6pBC47vDyh
edn2iDlgwJ44YhFYBmtE8+N85ALM87VUJ9sF6w5f8HX2Y2uPv6U=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
BdZ+ePnHGG+yksCfpNArtvwamifydZoGVGta2i+EFW5h/wIyKjNQ14qIQ4nx
W+vnF18W/C7ZNawtXKB5z720JSM8ptvHlMMlBYAroVorS0OwRfFLOpL3ZK0g
2f0riz6a2DaO+4Cyc807oGO6xRb4g7nxVIRPRBBYRehOx1FvldLztAzf0woC
v4NdAouyHBJCiyTgCE44Ai+PJXpaWswn1nQu+O9oJ/8xYhTOXsSqr1zYkwfr
F7t41+0X2bRmAbeCzg371r8v8q4+8f2YGMZ4OXNC5y+YyAzK+mfrVEYhLyKz
lFixo9gP5pImWG+gQVcCv/0BrClgw1I4Iv5fOiMHok8U1NNmuUhAtVss1D1z
4BkUqRLrhBQWvAy7TtQjeyOiuyZPgjb5JucieC5x2LJDPjj/N80Vs2IUsT/J
Zv4rz/pzTG4zk/FBedtSt+cfjkwxGs6SDDaGfyXY6W5oCxmNi7lD2TjDhyJ4
43zAj3jXFpQWFUzmxGEMfycyJoz4ElXz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mGnDuolv+1yfOimu6/Nz09Lu6aP93+bpfmr06WhrLBHRSpm8VVyNssDSIzRp
+CTTylOFan+0GJbpOua9OG5mld5JKtvMzH8QAezLOwJWpPtmhqnF2r5cBXqj
LQJlfi3qBqENAgFA0wlt2yTAN39vP/UdBn7BVZis4PpgmW5z0+0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CSB9htmPkAO++cmfPKggjlX2c6Z8WUGQwNLfswOuD572G/ow0+ayzKRPBEW2
bqT2HLTf8+BqZ+piHO2t1ruysrVbR70yOCbY8+ONX9nGhAc1ePgulpuMuuTs
P1ffmMX4V8wOudtwSlgQ3VUX8t1FvzksVEzmqClMIhW/paNV4MU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 992)
`pragma protect data_block
wTHCkwkiBCZn/NrqDDT4nWKNzEWM0NNrHJtA/8EmeeIv1KbfWeMh2ifbmLVW
05pIssSmNPlfE4mEDBv7MCZQ1HV8kYu+Dh0VDIdMnmeDUizKWzKituxatYea
ZE8LIcijZ+/xCq/yeUTsOT1B4ShFYXxO4gCjiGuRNrwgvDT5Wn7UdDoQwrjo
UVL1p/ns9tuDrTspp32yG6+sKvHUtBmE9wxGWoT2tiesTvOqkjEnOFLUauIp
oSz+y4o+x7uV+dxWjHhHRy1NaxjHUaugOwToaED2Rxs8EqniQACb6uiVQM6z
BUicGQJwTmIbIBYeoNv/ZG3UdancA7gzk9BCGXgp6d+81tvgp53sA8ujGfyG
LEEjmwbx8xkvKaC0YwEW7/K/BlHGqrm3UDt6+Uc7qFqX/D19a792nXyfPy+d
KOyXWsIMNRp/1nnTfmifTqC6jukrqup3e6ITJnfQXcmCABnXUSjrOSzrfxzV
keX52TxawUtxxS1UgW3kMgBLUyN/T79yscxWC0zY6B5LVLKjhBOjagGeYSYH
+tUB2sPUFSYSRNI4cNbJLD5XHTwWwSoE5qW3knhbovo4Pn1uXvtQVuTz+ad0
4+EVZ3nmzZjtG/OBHO6MBkJSUxadCQ/gYU/U2N0x/ASBhxXcR3MEK9rKilTk
7MUxLD8oCBQYbMTJB1byrFdis6Qr6yRWGMldL3GYb0dRER3TulYmD/W0nuPl
4/dPwQy72LSm4Vm5gbG+fxQlEG69k2gehw5Ry7fO9granL1IrH6SbtRIW52i
EoZxrml10JUkN1bwunum5k719XGEekS+zhbMbjMvcipm+NM5rsL8/rZBKRzN
C6CvqI0T6VGZKcrel8EMrXBy3pSUVO86H6Lc7D62DmBH8KRjv1lg5aNW1htG
P11xJUEPr3qD/nbFYTnDZqFpTUCNxWgCAchMQpyh0nI1Ag3zd6MlF6BtIv+x
rU65TBei0eSageHsgbz3VK4r/L+wmbGEt4rAzXoOul5ZRQczJF9RfGzKi5U3
11VeN9hKqfacFB9M8oLWu6scPHV6B/92Herfnxsnu5inRXoqUpEohFMHs4Jq
455C9Boav+blXX8qBLB1xBvjbH787o6P5UneFN7BYk7NdXCSh5wyTcuSYbBS
J1w8T7qCY/e9oz865V1iVuTBjPi7+BSv7L5G1aHvfLXCH8eaVpZt3FbOVd/u
/i/UOsCoRCt+uy9WLAVqsbUChIA+BB83vl1RxdY6pNRc33Xaxc/IbufuZAsc
k/VLm6aTeB06OEed5Gm6vDqb7lfiSYsCB81deeIs2EgRpc1gkNDTqEndcyWw
2AU=

`pragma protect end_protected
