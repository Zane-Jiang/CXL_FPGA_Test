// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GrF8ex2/t3zBUy1mA0FZXFfFD2BpDaYYNkVqoEP6Tg406cl4Kxh46tU4PReA
dqjQAGZeowUmCM+iD+4ba0owEqerdcBUlVBrq9P9L7dqDtPSYvOBHi3oePW5
9b7m5cmGakEwX6qbep5BF9LuUpZg5rPV0Fjd5eKI0Ujff9V3NSLqlK6oUli0
m41CK+KeZMilDhlevxQUj+xQ+pqr4oSDhJL5zRB23tIxqbKtzSvHkeSWVIGR
ufH5UtTPUJwAhAiR5UGXJMav0MoAqklrf+8u56FNniCckXAQHpo5omS22iQH
ywTr5Whwl9Px5WYHp/xxfFhmoxOsArZItIJnTY76Tw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n3/dbTVZYHMvylrk+MVy9bWHxSRq760ypH6p9pevJVGnJeZPLcK7UOew0DxF
b54TwJmqIvCVuCbDT64Pt8VgFv1TA/WwNdEcrN+StjB/i/i3eG7bTKUWJFIt
nwCw+0bjLfLrClGX9TX/QLwihKpgd12X+s9Gj12uOIb/c2luF5N3eGV3CxQG
vABVprT+VZgyedpFfW5w2X8gEQwqn/Y2PM2nbJk9iWAdWVgYaPQcP7rCg/gr
A5+X33Fhg0VVcIs4bYs8H6xZR2eRkaJCjXC0oRDK0FwRUg83pmToPZ/Jusvp
bsLQ2+z0NcrDSDnXpAVvgOYsYRhh4+aT87bRjv2c7A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NCdXwFXQjlDiFgiHuPVFGed9TXiiEEv5k6bPRMMqElwaohqvK+JRKC4yjzot
FF5dqxXsDwdd1rSVY0L3u3fdJF5GDDqs1Ji+e7ACggPBaRy76fgXVUvhnyQR
DFo54+Phr2EWYCw30cSjOaDjRVSOQyzQRFTfcEmyWqciqcCPJjASxW+CRQPT
1iuJZppxJ5ey7hAXSobLkTAygLL2qQ15dpBHMHob6CRgSp47COUS1dGOfe9Y
r0tPGu7keTlTCe7Py2v5K1rNPjlhKVhHvW2GsEjFKUxcTEpa/y6ewxehoDZK
PasE2vTLhOGpJdXlfei+m45EPkcFSS2Gg2XLe3jvnQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cONe09v00OAI00D4ZGL50BNgM5adNfV5M71xG0ASAEj+/d32Z3KjEY5vgh4P
m91Fq7LhALdyr6sQGmiEPBk8nm4p4CN5DLtZjSCRC2jun+a/x17XN9L6O5Xt
WbYaP1CkurDY5e8iEEtcGNsKJpnhBaLO3V7CU3P0tmzzs0+2KMo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XLQc1/CJD+wONGa7vyU1yF6zYebHh4yYZEbppmJ4ABe4oeB/tNOY+xdMIo+j
ts01MCISTjbICkcMnvH50tXqn0EwW5BDF/VIhoKEbjBArHDl0R0J9G96a4Lm
4ErI+9jhYYbASK29Qw8XoToDACoMz7+dh3B6JhnvlWuHfYRTURm17ws+wQ6S
CRWYNEJfNyV0lKN6wyuv+refLEg/bS+/BCPynz8mHc4lRh/q6EY8Jmvpj7R+
KixYQQZ7fEK39y2Z5OivM+G+wW4AuZymESfxkgaTJVqWNyPEQtYmBDeIQ0d2
qJvDBbzy3mJluNVFDtVIGF9lEVGEPugISdSRcRBRB1j9Ab0iJpogAn72kNI2
35U0m2ohlVmcnW//6Vi0ijqC07pXew13JbFQHd2AKMxZSmR/NfkJ52yg39Vi
CiVv5dW7EsHMqJ7T/4aXWMbP6HQaCXJg2REUwLRUhzKshmK3XzB/GHq0QviG
rIVZ6i7qz+KSTjRFwyZOcApYpicwHFEi


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W2WpQggDel4CTGzTpay2dg4YwWXLD0xI21X/DpVF0E5+3snIeUiHGoUBEUp6
vQeR29c7OmAz7MU3NT8BpkvxyCZG8wGEnZSOCevJjHMv8rMkuMc5xL8f9tzQ
EdcJ+/RqESaVDYU5/xh7+XxWRbaLaqBVccIoLjHZEtIAEvqjuS8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eXeUahl7YHeWmy/svAjXHRTUtghKU2skEDs8KNhuRqNxdk7WZxkFniwuZWBu
kdjZv4ddGjhHzp9p8Bwa21pbCpJvj+NYBFrNryw+NqOnqVii6DJzumn3/h6l
Dt/hzjCKh1BIA6ydvSCbXmrmqjH/Fm7WL+UVuxWQ5NZtUtI6E1k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 622848)
`pragma protect data_block
BFzW2s/N9V7T8yUoztWzqgji/Z9Petv09FjKgPCH98Q1CZupizbLEeYDlTQH
SKQ8EuQTgR7xRCFtcHFA1e7hBVMveQM20CAAfCBT1fyRdghusr41QpWJD3Na
rx3C04RW4rjODqdV+kFBcqvox7oOehGV4yXkJrNQwPuvjp5LMjk2Y5l9PCpi
Vr3sGP86FNYNVHaSicCSH/HHbl2zcDQNjlNuk1QjyONhfjwjl214MtC+Gmp0
AhhNmQ7v7uS7Gmb6cq/M5sp9IHCqt5IYS91FYUNbKkNTuyfcM5TrB6bOMEMR
mho+MMXi1NM9tGF640zqVWd2lIR2joUz0C5kwS69nJTdPtkj/lQVjbLpsEgM
gSbepz4SC9tAZok0fYkwX3pXdL7KNuqUpIx4+lLcOPbfXAE/CYh9wMuPTdHv
310S4VQEi6o0kE9XYPA2aHUNLGrtzs0thinxO0Ay2Zo+9viW7q+RGjfNmppI
S3tFFS0pX92cWOGHX9DcCIxBdKrJvefPp5KCun5gEzPj3DXii9TDedn/EcOd
2Aqao76cPR/lnFzb6pzzJPhSvbtdaclyzpqvYAjKGc7k9fi5EgEgXOQnE0m+
Vbn3QwAoakeAZsn7B7z27mPB4O7h0Oqhiywj/PoPyuLlbRhFGosEuGeHP3SG
T00GvetVUf/rfTAWYkW1SDl1080NtDtC/Qm2q+YNpE8+vt9VNRqe8/nra1Gy
Hk15Rl2bzu0JEMRIHir2YbEeg/1eHFarY22OSdXS/hjP+NTha6hdfT5bWg3G
CkbAcQPgB1CJhJe2scofEb+iwdX69Q8eMg09PLMgDO+66vu6IFu3qA+EHshu
ngX8Oimc6crkWEI8aMIIY+/FG5rm79Gx0xdHg0ZxtmZECnk2KT0fyVZE7XWr
dSur5ZDJnJiCErc8mBAi7MFP9Ax9r/jHnEDXbR/tSP1MWtRHkVq3i9CXGDCL
G9tOS1D17qG6LeBz0DVL33NSbT9zxbGyOj+nSBBO00rMVBNQAfSGClcTB/Ft
ERLes+gzQ10wbq4S3vvPvai7hgSn54Ztc4N75XloWhV5QS33sjJeSEEQxU4B
SojZ0XhqofHeFO+tnFhQk0OKBP/h8JtTtLYUz/zzPpJ9H2l6gpywr4uN8tqs
cs0nQMHfuLh0GrFruppSllH9ww9FnpO0MaguK5J1qaqS2FHX+jAWEHPkwqAS
8WT4x4S3jkfw2fxjmpI5+aiKtL+jYiYTliu/gFhKhDPeUlqXBjcHxyb02Grp
jzqXmfqgoW+La2iCyNGmDG/tID/rMzvfYodK6ZjtDzlUqzBa3evfB7/2Ar6a
R2MfN1ft5FKcjNAfhTHbtvK9ZXzl+UUlHrfEoc3EJArTyTzdN+/58eAVL8au
LUGbW+35cxhtbXhySP6cCrAb/ylHM3EDcPYhNeX8RdctcjKdeoMjOmqxoOFT
mHxTmvDfw6GQSbTE2Qo7ey5zHNOhLGz2EPQteXc3FjH3GgLvXjWwYjadB/NV
fOi9Nt2lUnf8g3KyXR52MfzMbw6y6W+65bJgBHK6qxqg6/EqD9pSJSyxcdCP
EO6tIKNWmuY4ONISivh0Ch2ZiUstdyv4SNiWhbg3+e0hLfq3cRMl+yMYSEJd
j8zXP1cwAnaCru9i5bKY+0NxJMqTV0eGHX4UVQZ+QpN86CEOkYNXMXcyqRQg
CFg672BeU0iIC9K0AsM0irXiNeLWFAHXBYfHHuuUv17qmumj6yHomcN4FHAk
wpOZj7kycHdOCAh9XvuM6WkX3hHXI0gN3KLAcTVbaLpAn1tjtgIaxhXn7c3j
LfTjQHxWba8Sj919J3AY81soikY72fzOC/rpUGonNGDsHlqgqJk0CfQP6J79
WsOMdWd6wuQyQ+qbfvPF5McAywZotQoiSyeflaQZbk0lcknyO3Lxsme2IN1/
MQN3YzmiZwYGNQXno4RFSHhwgJUxle3E9WVAaaEjtwJMQwc8ac43dmETpzE+
dwCgdKfCacriw97BRPzaVe6lDQo9MM/Jtw4HH8+JYqKHntraQ0+xVbLPZuUr
EkMfPP2BVUi6ppoxEiUj5rigkX69AEZkmpzi0E5ejpEK25mf5F/DqS9IAsEW
1wBGWsAiw/Nk7dgwt5jwqtz1uUkAo99/1wNFotNS5JtqWV1lxrUYoHWRMgbO
I5gi+AXQGqwWEYJLVYQRybV7RV7gHm38TQcbRzRT1SOtyExJ8XqTTBUwyo8R
MgsVT7FZ2IhVBF6JdAmzLYMfEwAVOaKuVH5NBRTLmrtm9nxNhpNHJPrJ+8e6
Fgp8bGgjAx6mWiQWkDVkntDfMvcZ0b/+zN/tUdHEf+n0H1phs2iWVBoKC+Hv
pmFRpZ1+k9buicJa3VHrBckpQqrcfZfGp/6NEAFUeRrbliSSUdy4L8UuUqMy
T+HmPIuHpr3t18lkflwOSvqRudsSVeGOtWhJSoQlYrU9CwXUcu1XLhyOviNk
4DHwRPH59ELcG4OG+SRpJwcOuJbp/WjypM9SRBDsL8AcGIP7C+OdenrTD2K0
H5W52onZUfPRN/yT7GHB3R20SmaEO4tVOLWB0z/4VW5KrtDbwdSghqxhshmU
eX6sz6BP1hBl8Mau8W9zu6APksRrEsHg2Z31N2jdG6MCDzB/oYKmwCfoHh7A
x8BIj2bgrWT1E+U7qX9mkPzjeucdxFsUmE0nNRnuLJFsuFNcZXcYZ/LMYrIs
Inao/GkF7FCUJHHBRn2VioF7cE5O/IhYtoyxbJ9/4KgCSHnnk13oAECw9Jld
dGRu9FG6p0eHQui3Sb4qqRQt/uExdK2OZUIMJ0jH/wKjiMm6PkkqKCY/YV8n
LZlo1qNNr/09q9zClCZDr9W/l/DWdPEnqkEUkHMeEWWPdUdgsm6v3Q65V+mR
I/oDjBwEzhZVJRZd6f2nAcNndaR8aQOEtNJNRXIAjUXxyN1dRZR8D0k8ibWS
K/n0h68GgLOZ3BDSgr7/pHueWTrkFxobD7PgU9oSRE+eTPeMPYBNZ2xcR4U0
wG4Vzqnxxwu0WHYxtdcqb2JYOrc6XagwZYsCeCN8+HbyCJHxR3L2T+PASp1m
7sUTt7ZL1/KOw5zo3H+4tWWkde2mG1a5RtLhxNRU9bwFGMYO8ER+yvk35UNt
K1JKqkmt9opCeGmZ6+bgoYXSL1LpBkn1+grBcVPyMGDYRDwOS/iWljmsZciw
/PHIkTl0qowCshFkuedHFBxmmTYmYr+ejA203+iZ6RhEh4bTUVgV7rEaUBmN
3kskIZl3S+bGAaFU6OUl3uuCDyW/ao2tCZzjohO1JFi15UbvdKWqHCVk4veR
SFh72f3zjCvmRCEukIEgS2296NdCd8pBAbwJlethtPFOJxUMdl5MPcY6ws8w
37O1Us5oDEcugvcJSetsKNvSNvgrOWd2j1cw/KyiwJ5q1rFN+KaIh9kmabH9
WICdUJGwsxdZZZ7Ghnf058pQfa90LYziwP6nWvcd8Z5C/1V6uoaaXCH/Fq0y
DEV17jmFcc97PRIteMxnt077KBy4OST4d6RaQDmvGibUGWhxsmNW62JQQBwT
MH3UYkjEHXODoGO/cXHF/x5fEhfRXJNHOhiX0FWN7DcFU0Of7loEsSyryh64
eax6MtYgUL/wCfaKCoREdfuCsXpusgqEtQABYcC/JDfrvCSlclJfBIpEVLsO
NrLlhb3yaw04fbMcAHb1c2U4r/s/xBY+k/jaUTIN90OfcJvpAKlkrXaKuR3e
xs4wg2S3TTVCnI/V8z9QbLHWz/IR8UKa5EWtlNc0tdcqETdFoRY2zhwKbNm+
l1a6AOKI9b0T3ez3cbblSoY0n4nQxXKwlK73ZrMLB8Pa+lvZVDU6IGmE1Dy9
8sn8r4B0XSyqUEdeBGGZEBWB9sg4yfE8CR9BYP4vOy/MnEQCdlIurCBTTrYy
CnEtQLXLdEIe9d1OmfM0EiDO2fr5LzjGT9sO3ucDHhiqkvolao01qTjxM3av
n+dVctNB1Ksf537ZXVFc6olt/M6Pf0tTgCHHP+cTaL2stjPrl9iHeqfYkM8i
rfrUqHNfNThk7F1mMAsx/cFj3RsYtlB50AmG0S9WQMY6QjkT7qKjW9At1rFZ
L2iuU/e5DnuDCyiswcvTWcSWwgd3YmPqf67f31pdFP3YYmE2KO4PgGRMFqBR
x/iOyohIenP+KSowz2kqfkQkHpTswXp5nSa+YrRPqGRiSY1twi6UwdoKA1jE
YnSWspUHIkdAvrnsGVUqv6KsaHLX7X4Nyrx2OwFowhOoqU/K6btojce+7uoP
m91xfGdejv8e4M2uHGj2to7zpWXOwFYWZ49uYmkjivAiwAo5e00VC/YziZAi
HXZ/osagvTfqj1DxrAnw4ZeudkGjgCMBE1CxxtYR8T0DSB7Bzvvnd7l2Abxu
CEN7hxczo2nUxaZDxX17fD5ogJfI/NwXzVQs33tYHEP/Kj1K+Dvgcz3HgYEE
GnJdTDpucsBq8FIyiKZWBmzHCLGbrGLfZS69nOiawf3qIBNJpj+457YnK/1z
pL+1mMA19dsgleCICMYhXxT4W1qsHABLxXTqk6K0FUYrDSccNXuQkTwyLjjx
AQr9BeKh0kZZ1DbZauigHzfVL4n7nk7OT984Ieoo8LM52qCC1580ZwR5D2aO
IPKbwIcFWpa8+pleSgitTnAvMTNVU5RQYskxxx7mqkpUzQN1aTn86AjnnQec
OnO56GUDPTTFoQX41ZJARxtNCSKuID31I9gjQFez/7DhVYCS2EJdWAwy65A2
VJQ4qVBJ5iNBaW+3z7Kea18zjo7rXNLTs9Qr18FdgqsjoEFCnJC52i/yhuT4
5HnRV8bR8yuJoeMzpUQASuO/X3gDsLmyDnbSVXi69LBjLZEXeQ2s+2C1p9IC
Fu/SEo1k0ivO5vYrM+4QoR82HV9W0OzS3FBkL70ZeSat6myauYJfjAZzdSZg
mdkF+rbVIzkzCvNWh2AbknSUi3FPNln8zp6ct6FYIarA3doAWy+Qd79nuyh3
yZzwNZQg9hNHMi6kY0HE5xl/hgm801FVV2/L5c19NYhi7VqvLH4S3j+DLHkZ
g1xNMiffBSkxSvfC08W0GnElOAhRTN1+0wDv2n1zm10HCnJtGT9uzwCmkPYu
5boVZR/kSneDCfCGeS/uykiAKzlp20Mm7x+zdK4Xn7JMZw590cGMNHDXf/jB
1/yhNosbulNzWMz8LWg2tc1xCetNmdbruWFG585pSDXSzyGIsBO7gzzfYfbc
WGH2HaV2oV7mMFRlVftmj0ZLOcTfmKN16logPorP5e/i5v13D648pD4a9QZ+
o8FaqVUEp5GE641Mt0ws1zwo2YKltSreAepx8I22QPTp2INUTx5GMD19tXOt
WkX+3c7Q8Zu4Vf3My/DCsa7vaBgLKi2Jng2vtp8EVJ8rThjmrAxosAA2dcuF
xU+Xj+E7GQfyP9+LRxeomWdO+t0pcItf2Ut5+Yt02WeqnlpReaSlfv0d4RL6
MBPlgc3HrLwfPh3wpSs7GYnRCp1utCl+f32uEmetmeXLHJrCUynxSdX7ftbO
zjKh+fCihPNCtShgmWhY487uC2hwtAtd+yqWqsNTNn14KKMIirS3N9bRYF0T
oEHCrzwSGZ2TbX8kF9hrsPuQSHpBMVYWf7aV0gr62AYbr0t7yB49ycqiEW1q
9kCaz6cfY9XuNIhF9XM/ODTxv2IwdrvGaQ2eRC5cN0ffXg4vqLmfo/+EFtco
fRUSgFbBljpACA3iZWMnmB1UDTYXw4yuJIKUux823EwdPZ0Mz8Tn4k0Qe2A1
YT5DE6gEegHrqpB5hcsvFV/KYosKXqCbPcs4LSC5CH1durHOCLdGnKhpMvzS
ZybBQCPke3SZ9aeSH9s9tdQUaQV6eEHwsPZE9Vw905cjao5bGzS4TLPK6cnO
EaKa4pCytcSscRKHyeDRUjQiAAcBn1DM/r6njQNgrtaNxOXYmm4wZWRj5JOt
nCTmlZX4S8myJ3ECvLSQO5vQXJSuOOy5ZncqW6kXIIcMnWivCwgL/t8bFPoF
qNPjuc8ycyyREwnBGnGb4No/r9tSEZiSDT4+xnayqRoNWjU+xS5anoy9fxB0
s46seeNII0gg0Htenq4Y5judTxUHxkxFMY+Zp5KRa+lB1tQpLPUnVsPQaj4k
qJIpHWCNsDg3kRPyrfrjfCuYsggREokSCaRxdh3a+dEojEYxmyXOKyV6Ft5i
PBlvnxUGTEv40wbChy3huBK2/yc4ekAF9cIM+6g9BajdQT7TzE77sKafFo2L
xKeN+L+SDYBK9fu/1NfhC4QgtAmOy92juFiTroxGmxXAlwGZfAQn1DY/UvYl
cny7UQYvcjmW1Dvxfx+kUzWNceErnT/pO8bSB8WdIa186V8o1IG7l9z8LnFO
QACs4Mu5CC7nLF2SGoTRYlzu8cLr9ahMA4bILPgjbO4ER3jQeaGzM199Q8Ax
qP6ApHDwniNEd+v54T0l9lCytu0WkEAPagX9XyfFD/jRgiy9BB0eqK58jfRN
9Ekcm2rs3XUaU29ROTF9oDJx5eVoaB0BGfZRxToKnSNoQNhh+1//4N6EtAjg
rKf07L2AHV+/0Iia6uYInljjzQHF2XLWa+QY0Z2s98x0jaFE2j30uS65bism
tcay4BNgLgkXB49Yv0qp/gSgwj5kvHrnrBVEgvmpPuA4IWoRrktvKHDJTje+
Pn2IFZSZX2FdJgC0rlyhUChIfyr1d6oh+U2L2WnUfrDL5/oZk42EFZRssikT
9vTv93yexm/rq3k+sMbt6uTPLQQ2y2Z7SpiaVNVlDPn612CECb3tZ76S5p+e
7+XufHm40icDKTBS+5a5WQlY+5bsZZCJkp96i60QD+zYGRJr3vIWzeSdXU95
U9lghLoqKWnV5zO+MQwHp0QfN7zu0d5+nu7gjvRh4B6s9GmqEkl3Bp8xDx/A
S7j9uMUhAZbvuvctE2tsEx7Vbq8vinEbooh21Oa9rOBhPXvOHJaeFae2tiVC
si5tQYanlnPWVvzf2Btte2OJP6RBBzc/pvFm+K/iY9WJojB3YpBNbSemQoU/
r1G0TpcBfBxNEqXCQNhQhmEFBhs029QCQwiJU0/2zyQw+92o4bL6lu3VNPSA
fSBJMIJmTGgsUQgAV4Wu0eR/15x3SsRnNi8FCG3wOsmJrPVRmwYWMoH1zEsx
4IT9HRKKU0pDcUHYfAK099TOm17uY2BVAHRI3hM9vL1TfkInBmiXLcPV50ka
afkRFz0Zj1BDkc0yWvA4Kp2sVEefwbf8SWFsjMcLNZ8IlBc9ZkOXdZEH6L7Q
VSzz+5IFkc4CVjedRXjbpQ/oYb2TawcMwvZ/1U37ZGADEeVMYckCUBC4vZVg
K+i2uKWYbm5rTjnf3+Q+da3kv3jB7w1kop8V5Vr04tPMvPT97X0qaJLvTiTK
cwrScEq4dyVuUzhNve+tyrPMG36w+e5ySwB6BZiihBNsudNGHOKcryVsw8kI
kCaP/hL92YFz2ycn8bsgcCoExrrLsHYYDM17o7C86klqhFdrUctEks8X2Tjn
pMEb8wtbulAE2rNgZylEKdmAWr+ehxip4GOrsgDClvxu6D1yDcWe4TePlDRM
ZLXMRNJdmHOiR7B+pqVPD2T7hICyBXiAgiFPM0XLM8D3rjo6WE5noQtXe+cB
6c4HH5dSPvIMBpiAcHtqvYYSu/1bxQ8nNqgqbkUH+IIVKufL4z0Fs1qQJ9jZ
9LXH2DvwyRbhgPtLwW9CbymUvdiQz6hScMBtC6P0CrIcWTWdlA/S7i8pswR5
J7SzQZtJyKOa7yyhXyc7LeoYxlpPlofnkVEvA//A2NuA25QxruDqQ4dm1/se
ScW1Gv1NkWpDBV91pi5PyT1xivLSpnE7m792KnW9Gq1OjWWaMuVxK8AI3eNp
/i4SJfxV7aQuxYLdV4BZbvbz0lpw2l39jcw7Qwuv1yNPMNk21RJ5+DnyIh1g
bfHdNkL4jz73znDGfxYqPvHX5o9fni2nYaNhHPRbh6wup2iemfSaRgcMukEU
qJHkSBVHnFtJpAHIcjwtViW3pHesTPZ7zqscuPTi+6VJdDzOyw983Y7dLLIe
orKGz5WbSUs/wn2X6jLigym5dO3KEeQUrQq2kLRyXgTeqnjvbiOP0XccysNZ
3JuSKK2xNrTAzOuoK/CEc+A3NSvpu5eNooD/Xu/KDcp0c1GROcIeGw6QpQKv
Sb9QF+aFyxScoJ10uNDVkpu5QyAcsNOeDcTZaDM5Z1hukeK3a2vcNLRYKadq
d/TInjZQUm4lkjC7MMWt/czwhbz5tVfqjDMPfzYunn95+Hr5nmwxNL9AxaJD
Te8D+KzUxrsujS1KwH77+1fJSh0Ho8wnGdV9xuNN6kFjurPSXbB+X6rwNXoi
JU+a8BZ/LnC598alVm6c3yDCQ3VcBp2dfaL/pIGXhB3psAzJVPrviVqC8vrW
bmzV3sIxW1yAoNYtptH2zlYHwv0aLnbg66jOjzN67n3c53F9RkMk6hcBeI+C
mwsDZR/bLvIGhsaX7YVoGtrdibt1BNtJ/s0uORJxjrIhfRoKM+Lhp92vHsoP
pBNSHxvN5OPy61lkryqaO0lQIB1/KroWKIml//KyqyijwT9dbZ1aWkaylfAj
DWSfRoNaAX3+AD8OH2spomfTg+SeX+i0T2KsgSl1+gVUYuJjRVqVYciflLg8
4LGdabxDbuYz4pvLKq7rXon7psqIPGE45+xC3eIjDR6JWG25py1JWPbP5iY0
ML0WH0CSZHpdrTyDfAn5gBPzAcWYLqQWLj/9KQ0rzVZtUXg3Idn8R0oveGHe
4Q92uhWnHizYYR2K+/7SjJPG0z7A8vPWehYBreqchpjt0MYX8wzUnaURRG3S
wefh4chuHNpZEF9i1faG7w/8AEVaYYtAQoiv1ZOzb8WYHU8gw9jpaqbA6rMv
kZRKRAy26iRVc9fuAFQ92iCacLDiHAw0/r67u3+5L9zNwEedeM/hZnU80Inu
VQomEfJBfJ3uuzTWP4NPcA9VvDeNX3xtRJ/LNpGGcgUJhUWycYD3EUhYSOxK
4Wvbeaf6r+rVMbBRjwa0no0xDoL0iMcZ4gps+wswCpdXyKS2IAxQcsO+iRFB
SlQRDKcZZVCCXTIM8k84xnGjYtUcoOxZJ5nKgbz9vkqVouOuy9G4OWmS9BrL
LwURpC4pmNqETCGW0OOTmjxQgZN8whpf5Vh6E5keDb601aCRforFunve1414
HJ1wSwvaCs0FOCauhi1gaSMu4bOw3DJQahLELNqwEvUblbYqzN9vAbVJoaKX
bFB94AhnjHgd61KUgz/TsQpoXNUKPDNpbyefZ3lFRE9YqDEf+TrqjVlfG2Uf
I+7h87T5Y4wJhssW78mBpT7UQqX34igQBIj66Wk4E00z2FpM/gyzB31N7ZWx
EEa1va6rGFLjs/YGZuVgEFSgXRMWd8lomOm4YdEdpQB5ZwSrpaKbXbzf20Nr
qFoRbVannlIsRDn7IMTU3e6lWVYEmdHG9ErwSUk9VFV7Z6n1E7E0RynSW+4K
mmy/FBWcWNnMm1GeR/ipxNxB4ANACcKEawdNlkueSGn/qdfvwmXDa7x3hOvT
tGvnKgpkEsgGMCu+MjSBA2RKLsmz7KXYF4I36AopGq9qiIjJv9OzpbO3sN+P
uLD1+dLj2cEQbbGjW4ykd7FzXUfjlUaa5aluyd/8d60AsNFVum9RtQtVc6aK
sowdE+FpZvquyvr4Ni4BbdAB1Ck9WXnsFgTnVZqBJ2oVsXp9vmKt1pB868pD
JEZ3ccMw98keIbP+A4KP3mNJ6aOoPt6SMV/23AnZc5Sye9atV84108AVQ4W6
9bSgEsh6C2i/rYG+23UQHMmXrEBPRC0GDiKx/7PbO51KZjRDLtwG57/kcnoO
FAZ1t6FLpK/EDBnEanhA7t5rkqstk8TVtDThvPJt+J6H97EtFMx6WZ9ho2iX
hnIm8FIEqTezrhDuBvdoHwR09wuZWSZ7aDE2sep/hiW1WdgFcroQyN80GgHf
e3jrQY905R1SsabJ+YhO7aFmvsqIeUMW2KalEAXBthCkoZwoTE8J6nzC8FUa
kZVAQbJ2WbOfXcnl9+WvzwrVNDXmkydN0l0s7T/VZdyKRonexPmb0JRtc6kv
OwoIS5IH/6vPSPHL6+/Qpvn9qqoNDA39fLCeWctWdknqrIjKrX7X2ZrGlGTZ
BiafcfpY4kkk4FqvvFss2VzO33CaCrWIVWorlha5HfceW+f5VPzyK8j0BpMJ
ftwdC7to93beGE9prNM/nxKsx9YYMaz3xmUa+NPLDdRRPQGzhxst/pXfSBXK
3Vc3H6Ln55A4f0+dYACAB9TKtBUf3sXa/C88Atw4EjwEanqMoEondX2635AW
pXk7cKhTYiQJYtZJde1IpWd2tVA3TgF/QETi5CceusID60DF2Cbmkc6THVz5
LI84GOGC21Jq9jvWRcSQq1FcdbRY/ZHcno1rMkQBhIzZEDnUvuCEonGptpKt
8ghdkJqZ8vTdjKQvUHLM0DXy80+q1HAbnH46J0wg+kNgcyPHWSPxd8Duj3Ya
8cpDu9sxkEaYXKnL3Jw2RNNBT3CEGdxTufVKDupEAQSToi0L9u+rf2tpD2ej
q47KIdvkYf4/yKAVOCaeGTyQfndUd6X90HfFwY6qBIBWUrSIp5EmNpaV1qIF
paQ+uJfI3tLXS5p5G2J1zVqSeuEmJK1FbUnMScRfGt3VAzonjYACLTPyuy2Q
6iQed0RQwp8shBXFli148vlUX7XnIxbUEhfcSMVyx5CbXGLyaaiZ8DoulTac
MsE0W1ijOmOqqDXY9TnVDDq3J6/fPNYQ/ode9/OF0xAbSELXFfHM3P13sUij
LrKNEgYSQevgv9Bb/rf3hhHqP1BfA1wJ6dLHRWzUqgO8JP34cXFcfX6VZfJW
rlkJuYu6g6vZiyirNzh88JWA8nfcQAtErXPRdilTfFK94uFLe5rOTXvt1Muq
8oq2C56NRE9emyy6GsuZnFxHU+cOJtqybU6bECj2DUGbw1mR2SVtStKydTRf
KeAvCv/Xtl49s8KEg4jKNDVUyzkNjq2uynZmvDTobUsXo24caOx0xABuPxaM
syNv6iDzRDm3iWf+v8/7RgrP/PH9ZXDuozrWzTEtgEuD5v2XB+l7o9S2fWxt
Nc7KLzg2lQghqhf9b1zyAs8g9JISO+5HmBMiJTYwuxBECJqWhG+mmPmjlHJh
XDv5mejwK3mrWR0mBevOSACsP5JczXMSDvzfuSUMOx6hGjgvhYRIAHSKhk/5
5CpD+spNk3bv+8tH3fWZ6OlzeDuXihI8GsO2co22HvdQMvAJUWvJYmgF2hnv
bcqjvKLFUm3nB2JQpEfE6A5p4joeJJT+pLtx48ECBY/8ZlrcD55GuGdWZ91t
EXQ6TJVCoXo9cgxSs4wxQQJbkPXlAkzxkncmZ19wDQlZTxYHos6I4wvsbfhU
a6deMZWu1/diLwYA7tfsA+jq8oVcsnaeH++n4quYkGR+ItuZ+OTHmFklK8Ez
KQnSU5aJ1q+Em3481OPx1Rw3epR6hEquSXniY8sYvMTxP+33uOcE+2sqx71z
+vFVfozGooM+bAuRIg8AlVT7y19DjtJLOKhNLDhAMFQmjAkr+q8apPNkYjeb
cY1mwAnHXRjPT7Q7YkdDwpFO7I53g+R9dZkXAo7DUMPENs33bcXVvznVS/72
9E1PdUyBNIByo8saQ2Ngk+DeTa2JGIh9AC9JR51Ey9zA7PW3I5GsU24p/r6J
SGhiUtgcueln3YAyKMG7iyOrPZByts2kUylEgwn+BxCzWdbEmwqZY9QoQO7v
pFdkFi7no0/1khWuN9wS/D8SlW45Kh7RWCxu65U/9aaCQtw7JiBw7vcddQ4t
mvkV/r5emhJt7xHAHhmYswEzKWLML/l6kIHMPddQPVHNDnXGo+UENYnVWeYa
6Klxk0B+pcbO2AoTxMlQlQ9lj6+MkFhz/85wJG6WX8uYhImszLD5xFRj43A5
AlpjEQriiDJjsNEIlwDaGO9iIG5L+fn3lzbFCT6PCXUWvRKR545RB0+rqYJM
mJP6pfAbTz5WQaVQcQyvvFWjm5lllrmU4QwyrzeBIIP0OnUDUnAdLekC8o8D
tURWHSSgAdIlZTo2pSAYFTLZ9Cc3Z7eY40W60oxFZgY+z2kZ7Avky+sWVxKl
HhmHaDlp8VteMudOMoT4raLciRxcVowV/yfubOG6r0PUfMLD3ZLK+mVGKQ2o
puOsHEpcohEGyOsCNUWq4H8FRofhCG3W7kS+Wgm8l/9ffPALcplx/A8KcFge
E2AZUcMTPfm2PZ/P0lCWtAuaATivl+sljqKd9yNsp/oFzhydzRSQ+MsOw6oS
6uX/IYZSnPuVFLRpQgywbRVD2QyqI6wsH1y4iYxYrXyxqouaRxwT+IkIG8sy
CkQIfP0WHGcMYCSTh4SYqkQIYAvq8UDVJzUkgO/7VTa0lq+LiVM6xRSWdSSR
9ik88QNIt94DLAK5sqa32DGt4UtSO0WMv03GXkUwa/AwLsaruIN+6XZSjzOM
T4zy1o3ZBXDkyRLO3lHBq7DhjZ08BpxG5bbs6gG6GeCwrcfqRFvWUFUIoc8Y
1OKGuXFBeZ3uyLYN8hV1MZcXhy22wDMF4GpgwdA8l3Mety+UCSdZpv2ryIn6
htQcmJ9Hd/sdGa0l1+BRbzpKwXe9BYynza5TS8C0w81iDgC+3BimFU4t0Dft
oH9EaLXlsCESEta8ZHA35iay0XTNLjM3USJhRvhXu+XoRvksUrh6kBOLqNVL
JCFepvxuyqRyaziWAoEvC2TbSli9DMG52GuQGQRPgxfm+4+5EjK4+kDx0fv+
j+5kkuZcZps1Qy+R6VPi9HkMOeqIM8hWXU8XW5WrJMGD/4LBViGF6fmxn67Q
pNLWdK207qJfGRdJNvjANJBK5EM7qhfne+4yxRZBIXeot33abbOYAw3fkO4E
b6QKUIjmHt4jHEU8UffI/A65uGbJWf6j+yybbwUvjt4pmlBIb1tLok9vNPi5
6o7TinL5WnlXbAErhg6qJre28pqVY09AJXJkujRdK9b3VUVHm9xhGn7HgCSq
Wz4OaOGVRsVODSJLoikM8DwWlZduDoNp5GVhsmzPYQJhVv5VFiKrjdsmCotb
0QBZVEC7Z+3yT0IDn0BmsmbnIo3XvrqUoyiYgM7NPINjsa0p5uRT4dCtTADp
SqbFKEQevIFtSuErBAoewKKceUrw1iSSEDwdv1ZpvuQwqDPg+qOLqjp2Gmvo
5WsCTAQMTFneH3F5PA8keWcp2PDQAUat4dhKkzu1Nx7lJ6LZaFMNdGEnGYlR
lN0EPPFkMZg84vhP66C22YrHBR8ZGhvEXBkaM3FkDGjmsZirw0tQbqMin+oR
8BIxgIJdGVqU3jdD/G0tROjL67FknyTnd4JqI0P9IfsMm/S+Bm/TxZhElUpQ
TX3zMJZfllup4Vmv+JdqZPrNLpoDgobT7e7URotqLv4gAIWHgsFIqin1czpB
b8HjgNXTE0itz1EFMKNfbrLvgvmEjGPOT3lot5RcNhinCOtt/zus5I7fNXiA
zfIzzh/ni0mxJYk1MZVgvCIeh6dfKp7wjLjiVA+kIWzpwYRSNygoz0JrRlZi
Qb37LQjJZJ1CupQ6PK2wdNpRuyk/1TVUtvADJR++cEZIFrFFOPmGEk2GMaRs
XhOXnza28WQb8E20OoPu/zoaCTKM2HnrFDgUuHZwrj8/DLMI5xukpH5I/IqR
0OM/G2FGVw231ipWtHphoyHHUyb5Ljt30sYmgwN3QLikQOIV4+NEggUxBYhk
zsaaCu/01+si/SderwjOni5ZXaWDYnof/6QlXcq+YA22IBhcMXRC6pBYPpsd
nX0p8b4zXprygX0v9aDNiamc4xh91nebrygr3vLxMDaOHQL7V8XxbFu1iPyE
lOToVKYJl2m2MtOIAxnWdJEtugQ1ca96liqWCquR+ZsJE+cIHYD/cSIr0D13
lfvgmGPv4/LKu/y9B59+NZ8VI8kELlLcx0eUMz2xk9JlllyZDqcaGN1qIz9O
Ejfx6FDlvetdZ+vEa7lZA9rqSL3+Ild3mBPwXHhSh6vXcyijBb6/bWHYmsVO
M4kWci2Bl1pvRSI0Rf05BaEmDdK7L3JehI16PPUNHDKaEy3qHrwkuDInEn9t
RZr/FffUsjQUAwSnIAbc0WYGyrjMfJpFOMflb5iYGrsm+TcQrzaSB+bLZ6X5
5x/v1xekEzfILjT8OldN8EMg7cf647vMIDZUHpDeAr6PiZhRLyJd7HPnco3C
h0+POkctF0FQdvn+Sy+NuNfTmYSqup6b1utgkvDU+fJBM/76kh1tdSPyddmD
0ynGFMW7rZ5acvtn3P/lz89LbG5Ie+O6DJIs0kIh3tyEdmbn/5M4UjywJrE5
GkV4RMCM9uNb4X4f2bhfXF1+hkG31TvQzaIgaKnrfz13gf3Wa6OE/r9WfvM/
BKP7xH+sagif+IvhLtg1HLEPJNHPWAWaFvuqA1nT8lIIcI1NKjXDP3KFVzHg
6FwbGyD2uGMxMWc5vrOTqaSpPL0j0dqDI+YH6oCn3oettlTl/mEtNzqEZwk2
tM5s0RwBInvTys0LpRI8r9va5ptLY8P9UOLKHsPVwZsOmD9uaKXZ+Z+vy8fj
B4hixjjmJNCzhQob6ZI33TF2bLhTG/UC6TIwWh7vL0PIqXkGdNoe9OoqAbZO
8P2EsLCsAwSAg/kMnrcW4z1CGCfoXnQ7YC4rHjf0ujZzaBH0xPtCLKOKKXsy
pHFjKZBDqBwUf6atnRsFjUAbJOlR+eFZsZPfiuvDmy1zFMGYfZUpNBUYqJIv
Q2660D1t3diDxPzfUPhYCA9hHQDZl8Z5pucbbEKCihcrpHHcrO3wqJI2cODD
6v5LDQopSmveJ32U3VHXBOyj4g3h3+ueysFmqNqa9wCA+Ae0ZouY8XJDNT24
XJWzuv35CHT+Li7adqXR3u90F1qlqn4LRsSHzRxuD6b30a4czfa0ARSGJcXg
2BDvUnC5IUTNSC+S3M1rHm+YETbfEl0h61SqrG78RwJYYIsXhHr4oz39rEJe
PIBaZkW9V69rGukp/AURq9f1TS7rWmIKt1lKmhr9sMP4hPVppCFcCz5RBeZP
LT0m54bkvG8GimfSgMynBrXZ8604HqwmnondY+Q/zfXbpuTjPMG+kox75rog
4wZ6/8ADemswAbV4EwjBpThyIk9EiaEFQKLQMXCL2JCY+5mbSqpRjQSBM0WL
Wq13cA/yB9hrLB56zA8CHFOQGT6bU+5Fe4hpvgwKq9yIQ8biCotOAghN3JIb
R5RiK6kon0KplwhiKsEfMK+EwxyoULD72zYEhzSwhEBMryHHtJR76ZfQgrGZ
apnvbFAuMuA9bFtBDZHti/KUQmJMBt67snPVqbnY38U99g6s3nqXJiw7xLaU
Q4gLx2VZHWOZZ6IEDkyCMqCw6+cGo/O5WTFtX1UyVcw3VdpWLcmzG3lnwM/Y
i3p11RdJD6e+xQCpDk46au40HMVSlU0NkrIn4kfVLAtdYkPOJf21KZOheflI
iHm3JcgMFVd/SpZ6ca7Bo2oM+WSxxcM7f8jK6sKSVSpRq7m/5cBb5axnLCiU
C0lZTwxs03jyAGvfj2qy31KC3J0yw+W20+dkcN3B8MPs6i4IaSw+Bvu6v5dO
vudvO5y0YT1bILmLxgocX2zDXV5rfKCoBvpYuQ3w0ZdN8BkZBtoOCTSs6UFo
5IyTVqrxbTdLm50hntuxp90aGJr6//1POrTZmgkGS7pZ9MUbgFyFXwwXJXir
9fgy/qbI3929kBY03PSBbcO0BZtVkQ0gqAmv0HHWesf7pCxXFinmzK3ctSlN
jlB4Z+QcYUYF0YpJj1uWrjMwFPDmeSleV23Ib3xMTF9fSO6kH7a8wk25HvHD
AZFhOnswabXBRODX18184WN8PSOggAzRxngFG4hwiLPCrT3DjZU8Dyn9r1Hx
c0ovRFuFcONrbhgj9MV14A5IFeuvwQR1TPwFs+uw1Fg6DONg6FMNk4rEQMt1
ipFN3LE2kQtNDa/Flq5evqcZOdWyGCdWy68R20GjUxwpUK0088SuUAlkC+2a
11AYSSTewCzxjxJLf11WYBl02NoNdZNYPVLqNtJHWqaKYV1GoHnqe6wWXpl2
oVVGoXG9B13zgU9kMTo4h2QqMY0RnWZcJtoCUdNkyj5GJkvhuiTj61l6El3e
YkiDp9qX9Y0oFOWKgreD3q6M9U8vU1bs4g66W7aPIaPBmj/wusGiM4jZAnr3
HYEopA/JbrBYrf9kSobcYm4/L2+VJ69hv6x36cOU6GPQtdTvw3kOlE6/LLUh
/WmNcWMbTd1hxl+mQ31kONLKf8kwPGTXF7up5affDNpn3y5oLWBPA8zr5sbw
DbkDxg731tou4DkOxr4WeyPeUDp1wdmFMSH8u5nwcae8wZKiMDu0ERl0pV2D
aa00rBppOKSfeVQ3zOboYRv/syp0m93ptnLOEwCO+h6njh6gi/oUlJ8EOxSI
5xBVl93geUCD2UGdVH0cGQsEMyrgx2iZJ1okHmHxYZ7wt38Ycw/dR5HmBJA7
5JIOwxrUMVNMYpFKLq05hhqNL+kCw/q0s7iMwT967opvhRUT6ujUexuoso5P
JC+1qE9ls+zJ13BpQmeS7tPrPksmbE+bbOx69H0nwSyYH8/5sVn0UHTtiiOU
sQDZeWgIFA7i4P8S/h/5KULpV5AZ5/xKVnGJrpfDLyFK1qMPJawbOi5K2ka9
NtGhD8B1Qmp5zbs1352dSk47amiQuq6iRnetGdY44zVGIOnqS1IbAeZaZ1GE
isJq5l8x6Cf1GEEDuEdvv682FdUaKl1FekofNfbVchFFFV8UrfEFMR2U+cBx
HRPSHt6vWqgifb0ZM+uXR+5+wl4s98Hq/+/9hB7owDdkNv89ms+WDgVPPusK
VBFeC13JQbT26EvGvq/+/w1dGkQ4L14exom91SDR+WIB8az+4+FdXwDAiLrr
5S6uLspYrBp0aU1AgzJsgEEFgACgv2ev2xkIiJ8TBxDSfakZ8BCbfmkmgiGF
bR3/wgqOMGgPF9qeE2IXZk1hRuUGK0zNOE9BN7+t8yJcMouPKJkmCBf2F5ID
8kO07NClUMOEm0DMpiacXBNmPejI9oHpEMlOF4It2TZb35FRVm1EQ81/pOVR
Zg5jirLdTHk5ItZxvpT9d9kLpU1a7129Rod0lGfUfCZ+bOnR5Wfg+8nfFrJ8
sd9V7BkF2NzAbRWE5o5L5qTMGZAwcZhTADbjhpWLJuZFMuy0fxnh4BbbkQP5
XO5gaSBlLQ2+oHnNNe0i8PMHDy1N2syAag1FmEUp91fjxkLBD5Tc2Ovnv7AA
Etrs48pPpVedCASHvob+IeUw09FehLnhhyLCjDm2+YhclxSlAnsEWuHBDMZ6
mktCKqY75iHafHJ2lVwjvkQLjlTNLWfO+CMRoLWjD9c8DsILvVcX4vzDU3jn
YNSqFB4Kvw1r6AlU3won1p1NvU6CyzV337mVS3RltWupl3LQmQ4peD9Rmool
VYQOa5o9ZbrV7/oeflEL91rcVeeR6KdIQTm3jxUI+S8kUVEp2shP/mPUM9ri
73la0jyW3QbeuTmt2eDxnuMfGNrsOxIf2cLD14q4URjHpQ4v8Y3swANnoppm
hXYO0FyS26SL74h5Hima/ZlDN/w1mfR+M2aGVxPt4PZ4aN/Dh1IcuI6+ypdD
bDXMvc5PHmZ5P3GOJDRgXvCfFpPiJaBwB8dDyzWcR/ZsAE9nCraji73zFDhT
2EIyjemPe4W9JApkzLoOIaY5/sIWGAuFk/OawiDYBIe4yTQlbdckIbMAfSSt
IYxYWBMonE4e+OxPmmArKq/JwT19jCa7kib4g85W4LAU3L3rHJwb5Ml/x3Cj
I5yPo0wEsyI8Vg3OLpRFMnpphu4yrBfYVT4O8tPVRP3+rtCwSwH/X7k8BuwW
n44Ts1f7YtmfgNl7oS2j7YUpsZF9GQ2LlQMAcXaICRZrJp8cjJ5oTRBtNUlM
4WvsGaplLdVr3fWs4txgX9SicuaYQ/0L321wGMhx5D5bp6u3X7PYQeF6heax
PSCbwqauZ1x0V64OHRlrTACu5s8DlyHj9SzTjcTKr1mBAXdNRDuCElDmIlG0
ecKS6n3MWITSqdeuHRW8E3E3c+1XQqxHYiYbY1MfQSrFH0gzXKFKTbd74rqF
Nrx1l9dZoOSFFRLo/KOhWMnbg5Nq1otiUrw/FiCLkXq/t53pNAbSiV673rmm
nrPPhXVEwAlwzZZrFgvYGfaFVqdKQ04lBtQVUsmnZHztCXBZXWGjbbyPAFOJ
gQmyQsZrqhos53g+V3PcoomJKqVbRBFxz1ik0LZDGcbqVNZ8nU7NAgUFHbPk
KKxdUdBgJZ4tyik0sAZ37YOTG+8NE2RD+N/QUXcomSj9ff9qsH+GdY+DgToH
a/HOCwunKVM29RHWnSTNHewKFbr3JLG0jv3C7GE+l977ZkP3dCoX8LDMp+Vl
zZWESIxmeWDdsYj1v5FaXhorl9pavowjwJQB1SMgyCDAkDrjUEVz6KIKUxBU
2lgs5cZaVKO9ph0BfN+WhwoKgfIgv6WX/h7K/wlycWlURi2n+H40pNhny9ne
RWLaAYi5lLoCYllGk0DD/38fg34Cg76A4JhiZeCfStNpoCuF4zdIOsvG1Lms
t2qgOeuNxim7weyJEZXYPhc7DlA7GhNcBk8dA8lYGD4uRnVOi8LXPxsuW8yy
a63hYMlUv9Qlb4UKWca4Me6PMIEzg73JsFbhaFodtvVc1RmzhVFXpUVH/koW
wp1HfmzVvGCnLE/F28C/Z7/D40bZ7x79fmmw5pWJUrqULt7ukIiUz9sfhnJ1
Vbc1XDuvrgygGMycysI0YREn88FlbSCSreKnLZ11ArMFd6VPLSiKmxVfZ6zF
hCubzQHiL9LoD9ROC+/YGuFWzw9juWOm+paFatn6sPmykcPdrI2U3lQcs1KQ
GZXww2K++RCh1V8oSarsllnsBjxRSxZwI/k9GyXZS6sY2VgqMaPuxzOBOCgT
U9eZ3uMGLWuPZIc0iQFq9FlQbCU8NKHp56aR4LX/oIYpErL3XuGXPa/X3GGW
VtlJmI6JzPV5QQ/HCM4XcQV3efVts1EDhBaq5akaS9U11frZ2AE1EXlCfdrR
CXLfAe3Yn9C6N0k3RBtciqD2ktG/EDpHuHNbN/jitFeU3Qu3pC3prEABLFhq
MkzZSIfS7qXkDLl+mC1yBOsUb4V9Ad48jCRq4LoBIZJYBIHVTtDOH2ZHkXOa
Ykp7CP6DUMp5XGLxJfeGzFlVOuYVbu/Yoep3phkdNE/VopJZI0Et4f270Waw
HxlMkawf0sE1qrjw1WbNnQ43bIqQajBGQA7Wub/HFjvZKMSyHCP3KSHDVVbT
JKEZ+rZLFQ3hE7RzEmmBrTTSQIerKnOFC+dmozO7+E7q4PIeV5Qf/DsDD2ny
PAhkxypon79H4btXYcs9Okoig0PjS3ttmrZ4VrDlIu0swWTYj8tMQy2e/X1G
qWIcgLjKceidnE6ZkvDLgrQzNdahl7pwlabIZNt3dx81jByI5LOLq/Nimhq9
4FOG8GA3EUQX521Xjfoxwwh4uJ3Pc+I5qK03r6svyAtlfpRl+PbZfoKhMHRp
OgW1AZFD/afMstdHqLdVuA/O6HB81rLpr0uePe5GoJcZpq+sdUM/DjJKDmxx
MgM+9fo4m15vrTq6PX5n/3708aBH4vuaJJaDNMCPpq6+59eVBodg02tIlt2Z
/LSu1F48AAN9DHUZQkk7GH/vjcKous2vyRAsvzWwx5FcEZG+H6zGnCJDRUp5
32Ewr6qe3gHPszLdkPSF9pVIGvN+xntbQZlCggHLCC4HfzEu7Cn0pFL1X0L8
Y108lA/xs5mt7/FVYAM583JP083OCNO1Yt02DMBGPtTAfAh9NbwcODy6c4Je
mFzXR0RAxuoqhBDqll8tIZipHb2D5EUXUGhGsSmC6oXzcxOmcKUGlmPIEXMF
eQ3DzMnVxA1qenI+XAd0VWm9nDMap+L1B9eDsshsv/qBlwJMKDfqA/vJISan
U27OOfHaBGJOxHxSnjfG+utd0XkA6PHl4ZuRzMhoMc3tQmsj3pEiZmYz/QK+
ODDbT50LZi7icBtoN8PMP9fvUNUSk5kzg60imw1CHR9KZDy6DiBXF927ycEr
kPlm+aJ99tGBooZ8FG/2EHPjrvgaHqgbtg0AlWAPfu5H8aQuu3y5mISreWSl
KIM7kT+rVERM0HwU+91sGqvM3QKX6Eltuq9r2s/bbvNO5dQxw4TZq9q3LyEV
XYzLfiC5iK0zucCIxieZrvikiMqWmmi4xHOa/q0K1tD5uZIysXCR07ZntGYF
PUSWygX5G2UIHTcD2L5n4VIcis+jypMriZsQFzpJ2DcRfzMTLEFOspVxytKK
x5zHRDlG+ITctSbwyDfH9EXh7xxArzPkc0NWCqv3WfxJHBmBYYrqoMn1LXTt
ee2mhQj02hN9q+aTsKotfNp3cYxw7WJjtRvxdmeRQhrX9e6+AMVzJlE4H8b9
GaHVLDGLYWfVy5hbR0/wc7g7YFBR60sAsOG9z0SdEZ0YAvVTfbCgpJMCA33L
VHOV4rg7P8EEuNWekbcOZiXvEf9b+bFPC6krn6Ry6c5YLpozyVda4H/isHAU
aDmJpAg1LC7Vn37Nd4qfUF2x1Eu7gzCNDQgkt4Y9vicZioE0vqIyysDqjUHD
IXZDHBqwdjZZk9MeV7hKpYMBCG0CfphyCRwNd/Uhg+2+YKGFmTgYskc+MneK
aFc/DOut9Y9Aj/3f383wdx3yZ5ZGQCzDtmeA//8v7Z8pdCnpnM25PrPM0wss
2dmR4G671Wj3HtzvZdxeRZMlcrxycVuPhxXD/NTf3cYB3e41povtvhN21m+z
aoKGFq95M53FQ8froHHqIi8IahBVKTHd8WJo7z4YbprMIBNViEadO8QBjLsx
7u2nEt4cOg8+loUvpqe3gjTtBfrhM7ozMLNr330lecgc/XRtoEZyZKXts65g
XQMuw+NOsJDuNmq2jnR31KRMBWr0mEKCw8ntwSTyn6SgksLim0MZoKqulC+X
mb98LM2V6u/2AamBQ77LA/T3UqhYkHewR2AGYcU2jgEGh20fpcmwTn+E7c9P
QR1cqJOexqFI7Wm5nJyClTcBunWsVOiLi3D27JHzNek4khayTa2Bi5waQ6yG
YCelpiLKL9yRLX6Tq5aWsQGjDuT0RXUvLGmr5t7kb2aRc/BaGFt4ezVK7xXX
OdVjDYGjIl7dC3VizavFo/O1gAIcs07P3FqzZ0g2UBHlIs686k4QIRkcHpTd
M9UjpOV90cT/RmZqB0KiM9aCSQwJbXud3XsArOg6KKgl+aD8JAcJDStnwDsN
8/7h3cApNiVb8Waicncjx09cJ6JIXSGIGRaIAy7HhnRwngApV7PNuP+NmsMb
YBZOTFqayJoiZEGVSVNLl1n6XB9JV2dOg+0u0VQic9JR8CByJAZNndyBBnbX
XOBhHZbIHZBPGDbM4R171GT+nv5kOBM7BNaE2yX1RpcLsUQCJ92Zrk/Hu4im
J21qBONxtLpBJP5Efjc2LpOzBfSCLLoIwzeQBVBISiGtZ2vsCrQUV7Oyi65M
CyzGvrwgvDeZz+8QN6JQLc8IZg/K8DnOUm72fGcnpc3FywkSceVGbQJk+Wm8
swQ9zsK58Ayf1cYd/BGi0gRPgEvFuELiFF5jlHrQea+V4yBlqAwwzJLYur9d
HyOOYJetFSz9a/q2MC5XyR17T5Rib3vPw/r3RqdcHUURG6YTwEmaqz/Z0zlU
uL+06hnaFOtdj6o72IVRLyxGxSCdOS9UKZP7cQ3Cy/rVZ0tIWsweZF+u0WeH
9IAgxaB2XMX3qbvlB7M/JV1y0TZAPfw3GUncZq9ijsJnAntuRYecqjWUJLiS
vghKR9dgqay4Lds7YsYggyOzW0/sg0BfsazTqnT+FEguwT4l5WphkoBFSc95
hCOrFCqtC1WEpUnRUoJjNKWgfa4qJp7mLPe4zdYqOxHSGfjmNYG/RdFrngCk
cXq+l7w4Figr0zGlGh/vSyhVO+WZP4nXkt6sbJAcLgp+w/hdpAB7O06LpqUB
ZlsXBpxWkpq3EVDkz9YlE53YD6DGu8t0qPSFswIfz+lA41P3YZpj/Pl0HSxt
Dw4IcOMT6kYWvMuDoDacHDuhsU5xo363gMFx/nNdMEycUJgh0L8u8Jxx+qaC
2Z0iES/oflIFmWiYlmGlDZAK08nrHMXxWA8gv3M0uBLJEFCZrYjV0w+uNKpL
ymfpBurRZsHbQNBetJzGLYM7UV0aSB0snHkKuEYR+8IZ5Nnup34QtFUC1KTL
S9ogGWKcdE/hESn2n6NkwzmGy9ljWtnmBTGcmeyVxTTlJK/dCjM542+3zPqp
9e4+TIUhcylDodmRNeX6HiIVtoBe4r3SEh0UiKEscDDRfl2csCN6RXRBTimT
ibvdRtz3tIywpbQ/uDLbtEHaJ6zpZUOxWCwLEbIJtAeXQdYLIoDmAltJfJwU
CGu1+r+Ij/b2EAiBAJ+2LkjlwS1yJUWyZUHCqQ6JhraJvKvXmO1K1yQlAVrg
656JLTiOqjc61Z3wm1PjLw5q5KnBk2/17bQahWBoCmC1KSUmLgNZHrQZi2z5
Ii50Oubn3OxtOo765Gpto0fjVXtX+3OvAaCBHdAljOR5CtVfgHglZzcjkobx
rM+i2aZhE0gZ2tJDY5sDWCOum8C+wNK/O6ParZI6+LmPk6wbzGWtqod6g+RN
JR1qURP7waxvflwHBcI42WoWW0RXNvHdFjWMPQDmf99vceoUYZhxnqAdBAsp
9a9p9xjrBGVttmiDUoJQVd/IaRHj9MaIdsnffSTBRdiwSPBQ7PZa+vJxHEJu
9+fhPP45k2rSv40hQz2Rh5cBZFr1tzF0Bk0yvZCIfTT2dH1iolH8ERGv4615
Wt9QUu1YPXEalYx/i5wxgytmPxS5bbiKjNBBm3MKs5VhBuF1tBfsSw1p4ea/
fpekJMFWaWPwioQtqOCvsW5Eh6mlC1q5koqW8uT6tv+q8MWKPub8c3Y2ef5o
KuFZxU3KYvB37t7P0lvS6ksWZulxyWf2KOVvHA0S0CZWM4pelgXgED9E6Dzq
7IzvXUsB8pesyzCfd7C+THb1zeVFONql+eCIpsRcqNv9AcfZeMloaoHwe7wS
qkcWzd7kJEMmxhcx2R+SYbUZNNuKwJE1JhMW6igN71zN8LOHgW7L//iCquUM
B+m/jHUR9W1JyagqKW8plIWjYni4jJsjemPuypUZ3tjH+HwfejN6ZVwiWS3j
9uESQOPpYijL5jYOzzAjhB+KvZ97e//vuVs7zlBFO9U6KTKum946k+pnqGRH
oO6wRkNdZE0fE0tLOrOPY4UtnCJfDokTBTJgXwNhRMq1Mx/qoqB1pBaRvLue
Ot8lQjy32iH/5ZeReLCvGejfRHK0TBl3w+zBOziCBmRSq7wqkWtuliy0ncBo
tbVEMU5tXoPmfVIpY5ghnrKDKg/JcvzEaqFxtR5PvsU0+ZPyvnsz2cg4zORE
rY55acaC3y23di0C76a+QjpeJCv7eXXdYjRNeshB2nzsMrCV9pXk8gbYzVA/
v0NWNZXZNd0pufuxpJt0U5gC5L34KB5d10By1j9Ch1gl8GTA5rF607OqONcZ
Yp5EZ4NqZ5APcgfE2v/MRHZn6djPGu7MJP+vvDCRxMG2KjsBDgOac2LLNfIQ
5P4Q9pCEkx9dsK1SBKQmxWmQi9Vu9vDczGXPl66Zg8e1Wzh1r52KH2bdeO8d
A30H3Z/xlzTTCHCrmw9KYeZGfaryune1C2oyHOe5WUc59id4vQenRnlEHxAc
6qvq9tyEmurqaVR2uR++YkMBin3/ypeDi7mjDYe9NKD5YqGyktp+NdSB/kNd
Ro8DeBqblFC2gP9bs6kEeG5CO6/JjenEHgnu8PYb4Zq3gs2rM7uiTpzjwXAR
ADanAxAAbWgjCTRym8pNE0oKUdSoPxyz8+O5QyJzoKgVkr+aDSiqlQW5rYmf
YNNpIhlUf+GMr54zR+9wJUEqB4CEQvPL8agFYbJNU2hfk5ZS4niCru4j/rGK
5aj2q5Y0J5U/sFOKxZfQDbkoGDxb2BItYgsB7yQYRpQCL7Aqh9UO1MUdHi7I
3cOz5W1u8IWrmYH53ENFBV7accJN4t46fLthEAUsx7QLzvUOJVQer/EkI4Ih
TZjWlZ0T2HptD6q5+cMMbo6YJj7cEhA+U8qNP/Bsi2nfSv0tExQKEFevvaI0
mGMjCwyxSgZnHtlmFiknnu4+WhW8eV9tS1p+RzNTrcnjsMLB4U3U4kRuTQZS
zSFWise45eGHcH5yT6raLDiiKtRrpxeyzs9G/Y2e23EfMbrU4eTb0a4/o39+
tXy3ur5J0lyvt4KHNbXjbVnPhYWQalgEOxSiIA+sUyDVaCH3jMFlauRaBHHq
O6a9z+X6hY9j6Kk81vK7P7H0pC+C4WhOZCeh+7GzZjKNM6u5WVY9/gz+9tUI
lFc23gLImDLHaIqfu/ID3pDcC+YoJWx+cd0NRMR3dJucz2FQ6cKP5LTwxRan
Z8cDq+QqSBqaHCI3w34TNePGtqMYADUH2NrB+trmcde+7+PaWlOfScCE1CoH
KKqVMINulyXCUz5H0g1KmLjLdjAYK7I86WVGITRBjq3bIjX7oXDe6vIppv01
l2PY0vt8z/vCmPHrACY0nOiuc/fz4E7qqnW/8U0zs3TUG7F/pZlYj5zft0R+
F/bZlff/0beJIf/PGhGoZ3TMPAOv3D7a5DzYByYdo6POQkd3jab+ramlWCjE
zSBpy5DsmbE1p1jErLg7gsrfbrfa5SYkhV2wbYnkMRv+WXEgdsgrWeAFb22d
sFSLa9D+NctfPEamZH03LQPjxYK4aTXPuELVz+BVMWJVV8neOGvIKX3iJOUr
M/cBp+Cq1ZMk6z9u97xdbF6YWti8JHyk/fD/ARg2K758ts+R4TELALj0hmun
v2qCLE17vteEsN5bTZGd1VssOavBGyK7URVDvJeMdRxS/8ivsXMGnRT7JkRH
3D8hx3mRDCGNFX2R0G204Q3XsACJtW+Caxd73Pfm7fJh1juEfDd1yQb4IzV1
JJ9YiQBxzGkhzz+TU92VzL7vkcULWo6RS4v3EwRZDmOifAC/wHljC77o06/P
U4RNGe6Aqtmy13qfPFAcFVVh7tOhGm3AMyI6y0+XO/Kcd0vCUgrXXLwcgCyf
yC+/SCoKck6WWYu5PkuuubWGxT5mstnsZ1zC7o7eNB/x3c7rX1nZzkzev65k
HsJJ+8rh8lUPOqt4EnscJUP+EulCRxg3fxSg9Q2pGEHhOAVh8br4R4kegRZR
gsBSvPU4dcQ6cFMg85ig6OKO/DOs50PSU8UyNKpuRENF5dJY3iTtbi0Qp24l
F42Fh4Cd/D113YR0xBkY3g5bk9qP6Secq48yScHgKL4awPbVGfq97XCZ3Slf
vI2UKziLm5uzfDBsIHssdU6lAuXcKW/D1Uft4tJjy/NeMG8OCHr8LPe6uKtf
xXtAsXHvpzm87Hjuo+Zy92XWlArTt4u0XpoMCKzC40vtm8PDeOtOWGSHN3HC
qgpXlERWfotMrf8VdvsOZVx/1r3wG4icv6GcCEStcQjFlOT6+1ecgH7eBzSq
Jw+4hTINxsF8N8S4NSp2lDYNqSQZ0PG0j3Mm56ZphiBOE5wlnIljOGCRgc80
u4r5AzTcb3z8FA5WIzE2UsNI6fWyTKw6v7Ch6nmKK8q61ja+/ID21bcTcLQq
4hlb00TulM94w1bkfoT5jH+Z3lOF/a0Yj0MAjU2NufQhSuVn6e2VYna3K1Rs
4wjhSd+vqlqLphic45dZCe1fpzbdOJt+OQ+cok9GKLIsWZoQdiBqLq/WMR1F
RNFJ1gGE0m3qfE3BibreVOdWvYwbtAYAB3UIJMQ20KR5NGKehJ/d/EOO5MvH
j2/FZbcqtVHXfen8/jkHjULwX7r39SURrnm3eKvZMUPgfcv4vltRx/IPCKAX
B4jJ6yBSFNvUJPrJQL+AIXwShjVMScFeUHK+qMtaFhisP62Grt56j84dy+4X
3f6T8MC1XxRZkbGFLoz2m9KqRmIZJ4nz/gUXtwlVn+osU1woqZFS/fRaJVDV
zBDZRsodHdOOAR3HGCksRAWb2DEk+IHKm427h9JIR87+PyZDvhLErgpnY30z
neRTSObEodtGFx1dpIfB0EhYe0B4hsoDxcfgVmT1m8hGqlrck49wugvUw/Gk
5OIFozn4hY9xxlWs05ffUx31rp1BiTtf7zN0D7fvJT/NeLEeBbzmVUyj5v4l
C4gU997xReSxpZhpBPqRUh9yg0LeQvUH753IN/msZWcALJLggprPFBTyBJ46
7mBCrbLsgM9+JgGLCc4wMlCbbZ0/hRrB7cN9CYMdqyVhLAEQ4Vc9Ytw+4ptW
sdHs97YvuN41veriXZTfaCK1PJmlBX6dA4WgX7S+SRt4jdcEwlj8G20R31vT
dB/GsLgZAUKo9x1Ps6jr9m/11dY5h/uxjQ8lo3zEDEigaah4nX7SPtf+3su7
dUj/Z8e5daZd3bB9Dq9MUQtCCaqGOys92qZ7OIYwMS6kSBF2MskqcV9hSuys
5BROAJgZXsZgrk8MoZifjdTBeVE6vL1108ExsW23v3jMK775JS3D8pJPSmtq
6rWjxHQ1E0ofUeypbjDGQnIZYp9jPY1QakOgGQsreerYFiFMHNsxEzUu8khC
GDtSBw/ScKpDfL69RXxSS/73RJxA/C/AmEZoQAv41bZF+P1Q6X6lGRIROUpp
Io3fpck4AjeyalnArgNOyX+E4yeRQx4T0KJbW/qYbl9sLFUTP4XPSdV5RnDw
h2Sb2vg74HefShABpUFG2+5SM+l14jp0gPPPH5VlqaIoEsT81NxXoErhVG4o
eSiZFQFa5v3SL27m3RDLp6KWiWP34loF256DYlm60KAhN4JsB8NVleC1p58W
XFDLtN6w1XBwuulSTJQvYR2HyJ3Md7ZD21zWXsl7EWPw0fFL/1t1EErhf9+f
oWKf1+yR1tf+6bUVlEX7oGn0blvIjCbChXRiR5fug+0O6slPR4to/9mfAgXK
KiVu5Udzcxh6NGoszYnjx/wQjHhTLa5uvqvgndIvdgimDJKyf7eAM7w8vf87
ThbUk+J+OmaRdr0Mv/cCgoD6Haj9kGSqof57opnhdoDJgUlZ814NX3V7ccpA
D9cH+B9SZ39CVjKSwUa+rRNk3z+EACtRBYEsTAlHkbtr6+AWaoEWrkEpPUKQ
pDWkJ+PgPwsjnxKiZN4Y2D+W/VcOGVtR/q5qtWsQ1wXwAcXQ5yqV+iPVxplF
O7yqLhaXHeV2X9WtdGxhVe/IUQiFM7v7ynuuQAEoGkV0EIHRQpal5i6YiI7r
UcHY9jRxc9lzBsbHdZsGNGe9tgKjDfgCo66jZQjHdMSOdjeb6pOWBo9doXCu
dT+SLPJqjgnoo6w9IEJdsCEUuwTAbEg3skAlz7hp4JCxJjiEPfIi56GJ6Pv9
y4TMyvqffaoXg7FAZPJdI6AVQeoHaWtf9OT2ZMYFmphQgWDSR1q5DD1Shu0R
L4UMmZahdgap2kjFXULSigLxMsjMkY1LHfVU4bVNRjss32c5raOBYM6vEo1b
JjtgKMjCXOpIljCvKztoGQuofWHEQuyi8uX1xopYzKalsamA6h+SpuC8Qot5
rJ7c3hMGX7z4/GothFN+JOzzdiNFyzWxhP6L1uU9f+n/eZhXTBmcD+3842Pb
tOfJI8eVN2kT63fDRhArtm0cOrcIy+ug9VsqHT8AiXOMJszQagwy+9dq8/4b
FcKc1AVv9d8bExIId2En5f4g3K+R5vSSCghS74YHG6utApqzFOCDnjdcEO9y
BvJU/FbgwXM7n7I1JYSS+/4GxtrLCnlbCs6uxhMcm+hUKTEEhk+rlYhTHZ7W
u9HZkkkKWAPiVme+mhrsXaw63yv9DAJMQ5MZmLlPCGd1GLk+x9AkyzBYwjFg
zSmQikc7lihUpuHFKUeeD9mXFqqRmPsHTJ3r+lybX9xtIoKf2ljkSnwykVJR
gRLqP0OE2sKqtN0cIdmsVj1eY2i1A5cSICUX2PTr/XsmySVfCDYHbAIOQdU7
6Ap8prhepI3RwXIAPj4iBuDnanuteFa3hqOIUIaOp1UwKulxx2EpZH0bUKi6
Ve/iWFmlCN5YS5Cb3PAehiu+Jv6zdJA9e7eEeDj2OWoh1MEVvks2OSU0RBFe
6dXpP+FNyEOCSKbnDRENrrsN7v4ZBmkiO6rSHIvfN2XwDt94eiOIAtIC3Ywp
xK1u96b6924gc7Fd6t46lYhJp1+MLB+/knf++YdW0ATS0hT2Rn1k00FA3KQV
cxy2kp3QnB93Ze8t/faIMBcPCACq+Dv9SXB8d12X2/qZ6Y4gj9VVeyFa+P9J
wa8coVpt5X2a8dnx13j1RJTzV50X7fgoYAivhq3+Wq1anBDI+fKqPiUoReHL
T5DyEq0k+vPGyC1a25zXPI7NUyW/mA5iUUT3pFSI8eEyxLPlqIgplmO0AThf
VHzGzRuU0mC4XCM9L/TVYdN7d6qgamm8po46+0zspqkOp9L889QqHCK7gULp
h8rBhfPwlZRq+MMVifclEP8WhSsPV0+35MXP0RA9o+blnx+ptPbOwXcSRvuP
G5KnNARG3JOFVBfWp73s5a8kSUUTLhw3RQYTqlKNwrL7MVnLwDK5evkX3XUz
Z7zZPoRKgTcSMXYJTjhpCmrnKU0VBemyRTpTY5DXNXB0bDL8aK7VaG8TiLPh
+ewiiHNukVDAU0cbQrsLW/PVHgJvHiEpFMP+vhSgVXo/BG2lM0Mb63X67eB3
SWTwt+/m1DBk7Ie/IIZvHfIUYBpogYo7llu4wvCFvEjMXTW+e80xRHWK+qzX
kzioKe0ZRp3xNPUpk1vHivcunhcg24X2pWeIlm7AEgTUyTtYKyQo4vINduyg
0RnIIS/s+UbjxFBeZZndLk63VCQRhJT1TYRNJeHKyrv2jr8VEE0NRnqiNaYY
h1grPb+4ibs7UO+Qj3uX2H8pylqe6pyJgoaUHub4ZXlInUWByHpNSgt9rCUJ
DcICZQIpVBfc07oLBDWYrIHw/kiNzoED1Pb81eZuNxl72YlnG35vnyjzwXZm
FBaYrGK4zsxo4oM705Gw3fXc7c01C4fY6Ep+yUkJDVTfJUZ18QMYYhuITYmQ
bNgpqLDTXssNKynp3R+KnBv4s8KJakD9nTTvq/oOFAE1ZavS1xV34qRB1oL9
Ykt58FTsu678KcTXlKHcpAA90SELLd8W1KTEmICgK4E7u3XP6GpPg4NbuGCW
0zNBJ8WLTyN53XU6qlCPPmjXm4KlOCAMtDKdlSD2TM0Mbp9kmC1wPpkh1Kjo
Z5IqOXDzU0W5GZIrwG49OIjhbcdh1zit20PS/LstnhgcGYuJ/U5w2DNafo5B
pRl3JG2Mf8eU80FUs7+0llJ/Ym9v8HSvi/VcShyjRcfbMMXvvGiqoNcSytx1
V7NOgRDUwhBiaNPjR21Z7kIVn21kPVQMJGZKTk+TIKk1e3N0MkOuowaQOEQF
8bbhJTTkkD20rBXQYC5xhVzb9iPAdIAclumQ6HdHEdAWkHTXQ+To3mPTYXR5
k9TgI5hA5HPK1QtIutxquN2No1LpQoDqRsS9cUeTTy1pS12eYJ/Y+rMzOWg1
FS61aakKZdo29i+6z6BzWzQLF7Cp+vD26FXqgqfCvG+v74iV2p8UvTcZJu20
koAHJMstEcwUxnJ59FqDuSUe0pbaxvktHbCd1R4PA4T6tqMvpi4gMHmXudHL
tGvvpt7fTkUhSM4Z1czp+N9aE2jDZdOPrybm8VNaDCEzzBO+gHkg1Cewvx7C
2RN39Kbfq0nU+ROURmpJAppqiK53x6TM/OhIP0h5c3tRYAGhanzY+wr3uY6t
NpvfQRUUDm1N/uBb9aFirdAieIxzjMky1VXymcUqKpmuKzO88vpX4Ll94Njn
T0pO52HbgNXmasjcoJqSfvzgL59fKjZYFgcOAqOflegM85wMJeovBkP8G04O
i2pVsBkYH3eBRcbX5iZpS+5EnsjLknRx2FHyXON/3dLt5giMHK2OHpZtRoZu
VnQ6UzwARgot2Om3HD0HviAcpAm4+jbhKK2s2ZXjOkh96P6BIYUwCqNUk6b2
ZHXYKjZFCcVTNDGnKgVRIhdbHJvsh7lPmy9ONTJoafOzBduRExx+5nJg3T+T
tiFkwi4xok1zVGcDkhySWVvDusC0xJbsNpqDat5uf3V82n3frMfd/SWmZRhd
R1jWJPj6gILlckNsuTGgZLs+IN5dWGQezLQWVqRkPkHnx4QIMBE1Bnhi3yCC
YuNujC0XF0mHCW9Ra5HyPp9qvjacJFeYBLAmmdl3ymjY2RNTs+pArW7HWoKG
W2XGXZhdX06rCOKaC94qaKavxu3EHAj9NvNUuw+jsvZ9RSIAYIjkpy5CXFs3
1OJuxE1xK8ZSMZM1Vl2z+NVnB63qC+EL5UgyYUDKnOhaIVLrvFcLV0dEIEdg
UrwmWxgbgmOHCvl4qyLKQcN3lx2ZznluMrHSL6eQePjSLVUsod1FuVl6S6aS
AOgvcJ5DLOewd9LunolI7QpcLkqv1nho0rqLgbfB0GgqpDsT8m+HKCKXMOcu
Z91GLLT38lYmZ0bN3peCZHZ/sJoRzOiBwvBBFIrSljqBS7v8XWO4FAYSEArj
VR3TNnO/hPe4qsA+HmwfeYfl0G/C98+2LNmoj5LK/S+V57Z5fRUbzGC6MUQ3
pqMkF4CKXCFYoQXvqxHPuuoN/xpKuOq6SR4MBkVPTw56gGXcwhqVZfqhv/IV
wUsRotIvYvTG6i63O1OKzEwJLPhoVIHc8SQxuKb4+zSGjcCAOjHD6Dy2UXp0
h1XKh7lie6OVHh4uIc/7X/s0XWp4lceevu5VvieJ5+dJc9ZCW0DdnfaduSDA
wMY+LeCJIoTXSn4WLHVZFgfVtRmHaf1lQ5pRv6TzKneleql/nJQn9V+EcyIt
N+uTIGNChxVmcx3VIMvlf2LIUjmo42lRqVM7I+Hvk4g1/rOYWa4QxMR8e21P
mc1Qsy5qXkyMjWgmRHbtT4AkBCgNp5XYBR4XyyAxmlppfIn4uw74LftucUaH
gwYDrGoIOWWJmB5oyeqb4cWyAQAEapEcnk4Fq9GeT9CBPOZIXNeQ0KAGo3Wq
v11GV+TJFJOcPpPvWxdw1SGDo11E8iI9GQNs7PA7xvjJuEVI/PxwIDkLhyrv
3k/eM+28Fu1ShvNW5uH5O3kXGC6P5acT3t4LZ1CtYa5t5+vRL03PG7v7SVII
oYQLQW0cw+0nPl3MZNjzbdfYLC2L+k1yPwnfIy0DfMemPXGziaagfKqG9+jv
8FEzME+hT/Iny1aKtTEocyzPZfom99d1/WjVkGvdJyYQOIYbWYXsupooCFbE
GF9EFs6Tur/cxbUBEUw5vLBnyOw6Cr4pT3TF2Cvvq6lDLpWuEzW/1+b0ip+x
gIgDVAW7mYghiWTeRMRAqNcngsECj+wltMVylg58LFekcedCaMPzSVBJahq+
IuG+/pj941tIe/YZCl7ErWYJ2MDyjnmJEOb9AloOhJGiAGnrOXSkMzF3q3I4
9SVCuOQi1SMjYkaoLv1KLEiulNt+c7hDjvmXwjX/LpjPqSeDj1bYp5VG7aR7
5SHJnXv0KCcbFaiL8FhHeeANCtnYai/Y3o2tA7EfKgUGddnzfWPqnYmyn+9W
MGJbvuBUZJxgr9FefpHKR8USRwCFJo3xCTO8RC0U+DdmgmWbblmouvXJYPWe
pcb1lRRQV+KXccj/+qZpj5zmm367YfqI0J6ucn6gkTEk/hf5ORziAt4MDSq+
ZuPH2bgLxdB8Ee6AhXnwX9Lr32/7QqcEEqlbwbFNZ9A/AWQ1knr6G2eL9s3y
XB9llzmRtd3KZmcZJEgyD7Zfo30cGBanWqMwrQUy6QF0U8sw1iB6mDfgwMCD
kyFmehgrhh9LVEJNMMlmkqbTfXejF2yu6s5dGA2479F4p4QCF0W785UYLFb9
7Qfc5g2xrBwKrhQtqghrcVL5/HjYigeKlynmPPrEIZ50/n+oCmFg5DRo0c6e
azL/XXbvkUZajIPtR16JNZcHzqjeHjaQXBUsHCq8ieW8X1Y/HYbRASUxP3vI
2zzJdLomTAlU7LYASyjCq+KBicY+upXz6GZY0EqvKBAHDTvXnZELjqwNg15k
NH1+OICcxSjOywf36Cl+0NfjBePAH24v8I+d6J+dnef9F2/ymL6oNojtIWzF
QaIWDmus4AV1xA50Z3M+CdJ4sxos9Hk5H56dCAy54WcoAfCjjTu0FXEEc7SL
cMHZvcoYYgSUMoUIENkCc4l962W7PLbdVXrUrztDwMA6BTxuVEG3EIV/o5pd
sfjwSp5eVAI9iWpcU1naSEBcfilBGZznpanJaVcS3hxo+gKM30w6ZvWfZWTf
mIht5dPzJUmTdkUGaiofjxOM9p5DgVvseEbp1T0yA4twQS2cFCwm1aXv6P5A
NmG69FwDVfJvVAF7KZzZog17j2Tb8txPZSNLosBKFvu6lw0UQ6kdg5QJHe91
i4CzRAjf6PWFt49BViYlg53O4KDW/UmlGUfyKHd0CvQfDajacUMeEUKhDQct
LyX7/SkprWzms32eil6r50M5v7U9OjA2oyzciXS91uOYptVTszonT4faFfT1
Bf2OIlHY8d1/tD49K+l7GqaMK+ehTW8TQkRzrar1+HLtBnAx1jvUUYa1X7gs
8nTjZjDcbbLYyYbYGtCOF36YCe2CcfsLSIYRCZBJBS9c8LQvXVtz8ZummgLz
VBROZFVDMA+WmYhUBwThXX0pZSGUg0mDf8xeSTcCM+boT0eMed6W8k0akdgX
6fvdZ1VfjfgdwgeQ0tWW2yIEMk9JoJ7UXl1hvn/ks1ArVPYX67anSTQRrFcl
ddpCV+vpjoMpDx6U1L06OBGwww7uUEH6PItovtEjjptIK188lOCEWsAyudqG
bJ5mjmZHI3aVENooiwsQ/zrLv9h0khPXumhN6VP9TgklZ/KfK1JNHsurkGW0
CXg2JonbgKBQgWKKcQyLoELkPLskXnvwREGMX78g9b3nvi1o0n/8Wd/l8yCH
5WUat6pSo1VqJ+5HDD1eiXB+6KjoWSwS+9R2qW0W/YvX1Im74XzZaT1nWw9a
xJdSIK3McTuVsYhZeyPukAu2MzRhcIoDlY/4yoh9dNWffGkQjr4/VmDUMPIf
u3SKlbvanxTmoZ/W2DDv4WiZUdwlYF60aoogXggc0Xj5uy9LV0IDYgZ2ip2E
cFxvgKeInsvGfcwzEh7QU4ySCYveogPWgupJ17MYTaR9ojOcJ3oBzxkDvIj8
/Cdp8dYPhtEjUvZGpr5IRYOlq8pkqUIfXbMZDsfZIQiJ17TilpjzesokAZmw
R+7f5SGBEj9XVDvyyo5WNMaBdXLjX+ogzJZq2dUeD1bRXUDXPVthGqCXarKO
2C+F/7uVXq5aFGrDBuALfpSJANY8rSrSpS9xGSKTT+yw9zCBr/93DAagMO9u
/6rDnMylnNqVsEgk+2JGZEgLkoAyuwR5sSEBKgFp42PvdLU0Vj2PUEOUjkuq
gYCBVyKTPqBYr8/G1XE/qt3TnGQVnBZxTDJri8Nw5tqVj2ab8wRr1ncEDJLd
YalvvY0JGzffky789wRXONGg8QpVxmK+uy4qNgk6E7doOc/UevJXtz5bqkzM
PjNWblXB4P5Y8eskul0GDxpu/9lgcaEITyPrcSHjqCppg1olv8gKgINXmD2n
M2ipjhgRIjHapOmU9jsg6c2llKSUPwFLogMrrdeMkVoTVpmy3hXeFclZ9wkb
BnWBEQJY4wMxUDqGqnIZFif0H6CfN4bNuh5QNp298LtHgiFvGidwUouJBHUj
I7A0nyTh9vpeHddU7Po8ecQO4+a0VDnPxf4y0bT3fueVh4Q63wNCoBDYyWzS
P3jFv9evSC2sjdkrhi19F8707uxpeMDLD0pikygLKPVEH2DpBqMQRd4CFhIR
vWwPL1/ME9SySX1qrviL7FLuMttjOmjYznkXd+Jpx9K3feNUd3GkXRDLrHe6
C1UjwBTNTK/59fORbHe5hOU7zluG/LdWB3L2NrxO4JhZX3siRl9rsMpabDbZ
RB0MQ31lvi3B4g2rEWzSh21LkZIIEhn5uSI1/ptpFbtBCFsjvywGJwvTtL/G
hwQc22lDnRb8ydtbi/3sHqxgweIyeQm8+nF1RR06q7LvMGrFjukoMeFuJNbz
RYKeJZMUAEP47vdslY8I2hZkMVH33XcwNkhiZaf/iPZ0hwnUDosdc1ihZPCB
Z5Bh47ynO32ReRFa32Zj5MQhcmBUoxVfs0i/TavDZGtIUY+KHD2L387oSmBc
F5b4TZrg/v7ywB3zCht/IQl4lrKAZ7JWfAmDV3KU9ieA602KEfzPGznckdww
/gj0u6uoZl2ZtCLU2eL5XmbOhZ9Q9p6/kDlmN3so3/acVC5r8lduW9cK2sCC
AlabqIYqkKoYzbt2gSwzL7l7cKJ4p/KKt47ejjRHOJFwNXVzXej7i75+wy9W
dlMkPm1IMuLjF/OxobhgLCbHtjBH2NZWmANr7Rqx7CooilDRmY4RKhbt/cFU
uDnwDOUvXc55xqSTE6k0F8/WV51VboO+0LjKmZjpu1vE087GDEGOod3w6d+G
FFqYhfkh1RC3nLYfo0OUrHXR+bDqjs4xZH6tA+/S7naBJkUwLlN+LcBx5oZX
yJnJqhMDnUGSrOtWtuwV9NHsfo7CggziSVA10yjE3lJZ3elYsIHPgA03Ez2t
cush1ydCdCFGq135Ovx46/JzjOjHZpf0rPmNn4MQZb6BlkPf9eBbEcuaj0w2
8sYMRGwNZrYiSoCsi9b0vYtpd3T50b/FLfFI2uO7KeL20gLKww3GiMWQY9zX
xXPpy+xIhILNHCdfKOpY/6dlpm+GFOqz11NW2dn+yB70K/LRehgJXhVJxgqB
G1v7jdkFA3a8k89dBFCsRA5CKP38/EOdJq/MMaU4fgaWKnyb63KQwRrZHtWE
LQ6U7GXv7dk22jk20+PJbknX8urrB4mdz+2NgBNUZTtwZTo2m6wB5TTq+tQ0
Gr//vtSKwJc0byuthj58TX4gdQpuk1Ct7ru9gkzw9FcwuDPftNhMIPKswAXk
AzXsWN7XGLgP9yy0NgSug61uNf1TLMrfJikG2AYF5eaWaJ/4leA1R2gCjF2W
u8gWWznOv9lm/cEKiwnXn8v5hCrPfvxHWceRJC/yAH5eScXonh3Pb6N6T8SP
KSqcqtI14OD4XfyfpVz/1tooQl9Z88YXm2ZKG7YNyy7LgXrOUmC3demWhyRv
mGU3fcmxmAvKyXnLTB5f6aLt7q9ADnAvoltPP2L/DI2Nqz8F9+zOroksuUzj
AdZXHplfVpbF5g6Wkye5+nY40WF3IjLTiZtdiqJtXEaUtD6YTx/45nJDkCnW
W65abXNs7Jz+bzmqZ5KFXYnBiSRl6Xk6Nj+hu9W+AfOY1N8WjCoARGcOSi6W
7+b3npQ2Kz+ILTfWIwHwTWESwM01Teoh9VTIf0tfUgLxhcx8n7/+PUQme09s
DIpMdEBz0qXk4MVq8px3mSMZNg5fdV0LkKQS/hwVomXSSe/ZLvY70iejs3IF
X4M0Db9Q0uyqS/JjdlxKKBDICh8NmnbV7EhnlMa1ywuoVz7N6zr0BPYwqRD+
DHegEH4kjotG+grBlEvYKBA3l8ByHAEG99CmcFlE30qcMA/odMJIpMgSSkKO
GQ0EGvV+7dTG3G3d3Kzfltgxo7xUO72kXT5PXl+sWhkj1gHSXGySEtfi9/3K
dFskQKT5bGUuH3cLDN6hgEDqy4IEa/JaUUhX+SmY66gVqeYe8ZZn5A468FDG
OnfIXwRfXCjBEdTBDg3nac62oa5rjzhlHrjTGcUzXgXV6bH4a+xQux57+MWv
1xmppFw2ncinsu2IC3BDacpjZo2rsON9bTuwYzNlsdArmCfU7legxkMg3UEC
odjHHJnuareAfK2YurddJH6cbHprpb0Y2RKPI3LpRQRhtR8j8aNAmhki0DMw
yYptUPpURhqAahCOo0yZjVpc/kDgCOEjK7FUIeaxBot+nXS7399sLOFPVsOn
7UZkZgE4X3Rm8rXjNGXZ9F1mySs/sw2uSShEVF9hhYvx9jMiHw2yjVc67iBI
HkMSkGag8T0dx5unPK398X7nd7rpFyVj6DKl2bbEFodJeHR+C7lNXoE3mFbA
HO/IVC2fvPWwvoJxg2CM0lfuzZEGrYhBrhGYiA7uzqW+6vuDTjpvemp/zMTp
LL7sIFIj/C7rkrYWtlzFqyHY4f629W7oNxnR6pjySAwjAKjL8v27XFNVQDiX
uVs/8KaOi+IGV0I3jO6m5z4iShGk8l4ArSXtUZRoWFaonGLHuNJC9hGS90At
2hm7CJJse2EITSlLqbRWkF1gvM0OHH/KAnpCGt8+12amTPaxikLPsPNRlMOV
wsQYdrddw434aMDOofE0JXgG2TbWhrQgsNsC991rLMVGUwxwW/2iyJghDK09
g8Prd0v/cdDmjoxtkx/KbUPhGlI2dkaw00dv/oOidWEUalxDSbjc8bjz1slD
Q00NXPOBWTvAOUF4vBzPV1gmgfkz3eoNhieIKGMAZXS38B4y3siXegrtIN8A
psIaXbtFYXfoiEFGzqutF8wz46Bi5A/IuOT4gysUHiv4Z5IucVsPX7vDTmeD
lW6/t1K63hG9b6eZ0WuH2cpPxz6bQtOiMLlHD54sUYBVbuz4cYqmtERfjNI+
194gU3+tXD71AfZbKSjYXX0hHawhLpRboNmM13Mm0ulxSQv/3n1kxN3g6V00
xhgdEfHiQvGYJnDh/PHntrOK1Bkv4gsoWI1pSGNXHAkEIXM1tGpSrj13Q0L1
uiCI4goR6+22BV88asKcEuWZHz9CP3RI7QEk92kZPspQ5fkX3W7Uw0QQMw/i
Rtrdrkp4eiUje6xh9hg+nzdRCsopMdIT255Ax/AO1D1kYpMWR0dowS//WAPG
KhirP9a3twrs+7B6k/XshHVjAlmk7ZXvmTJvp9yBTicrkXRX2Eb0JJ5RKr6j
sLTHKVVIRXBVlf8uhke3zzXLw1Vdw4pyDbXT+L6v2MfZnUbaaUc6TW5QcUwd
M75PkpEqEloapIyZjTZQ7LbVZv53skDpOzrNZ+/iPD6OD2t4hBQ+Wa3KMrGV
0i59a6aYYKibn9NKKKdCNMosIvJ5g0b4zgoSz171Nix8C7FWq/0LwuiBqEB3
CJENhUCyOnV9n+StIOVIAhdi0HE1RIoorPx2nhZLGUU6GRul2UALt+hbJ9+8
05WzGesnYztbpHFspgB4aqT+e0p4wDMgxlkU2ldEevt90/xmAblzNU+0fNZ+
1EZEGkctpMId0GvH0zCYr3jY2SX1JYY2xTGrxkfOHv6pmTc+/tgRhyLx7V9u
2e+SusyZSaNQfvDKHjJtVocB5O/8NsWjhdxovnpmgZhHSGRvye5F5HKVYk0m
W32ZnjymUmZTpLK9FtwVdu1uU/UdokXZfPSZ3PkFCk+59KqsAkTkcfcuqS6/
hN8zAs00fWUV1KE7lhCMRnPbmGeB/We2/20B54PHg1jGRa8YpZRy4WyLZ3WC
dGYzXBw+tqAgWITDpxoqj05MrzExRk9BrZPc4qkGHsbbhywFeJgu3wq/3bmq
b/pkhyJB9xUMOpyOtS8wc3dT3FMxnwmqB1KAEC/xrdu7eIrtkL2vv/8eFNKJ
5hel2mOlFoCqNftIyOXiq3+lE8mznzyatt6ydlCcRPf8JtpgeaEf0vkifKxn
st2b4oyRZHF9chKAq75R+svkr/MROETdi9+GYvMKMT+jJf1w9m/DWBqV3tDe
Ltvce2Jp4gNiXv5DnSXHCZMWyC3zBvbYBo5zNClLUXGF+9cE7FbZ87UEec5h
WPSTRMQXVeMQdsvTrQo2Px8HO/xdRojiA1fuK41elIuXXLavz2/3WHPDUI3l
ykv7IMyN7b06wW2LX6XhsndrpJRIJRqOXG91o5WImvwF9tNn8SxE+3q2COYH
hk5skyUksLvmFpezxY1oenQyC2Aj9tqimKZl6h0H/Eekg1bbMJE5kFD5h2Ti
Gjyd2nYyD+zwrfrDVpZfYs/LGR+6DvZm6c0rhCDzV97uRGeZmApQI7IDtEip
XhIy1idwDMr59zE41HVh/zJxnb/SiaqwCupdeqfePl98fwQ6VUoIzVKv7BKx
XWc0Robr/KEctu4VYh6kP/sTizBV5vYWn1bCoFk4K9RH6TIiEZPPlLshA4gZ
GlZUFFm3rln5diUCg2P6Jb0jgJ1D7hOGyMpcO7ez6nPtwuWh9f+qD9YuBM83
gYdtskpi1F3Tp0fVFKXdanIM6uNuhCscwv5km/6Pq+BAqtpNfanz/l+KGWhY
oJHZ9HHYEsqflVJRlzjCByPqcHfkDhL92Etm4Y5nJkOJW3YQVR81ESXZzmc+
EVdy1vIvd4iGHD2he7Bn/HWJAtUmDnDLkce0KFewu5v2YCeJfzyR+WYFcL6y
cH9hW44XvIUHRnnLJwf9Jbrwv3SIKPqzkwEgQ4AHoELYYAW2Trsx6AH2rBJo
yDo3vWRQaWvNUg5iPga0OQieX2ddhJICSVxcAEbYhIroof/jxnDQQFRufuu/
gEHQlLHUQQB+WPsbApWDCeH0KZGUBqWiUit1/cBRItT7qurm2oPnHT0WtFS6
r0lc6UkbpZNmzRuBHwr+s0YAX9LQigQuWrJZC5E6LN8JAKtZ3E5H8USsmo/G
N+SDt/lQ+3N+irijBzN2tvDh5zo+ry2GQiDE7fvSByVFEtYJIyTPr/TuSy0T
m3T9nJnFnTJGAdiUbtgMyMcnT7C+OXk61lnHJD5iMYiO+dwj/sUNEu8erxPY
NMa9x0Ej615wXSGBA6uuPbc9XT5umykXRVj+wzkz3sCcFNqOFHC7ikKigv0C
Cpvq+QI7BirUTokF+mgs6Qs1/mMBLU9Am+OHL0RjHsjRDi6nMBde9IoABUHY
VQfmG3A3lVh0cuU+PGEbWscHVZiYzndEiASpcOm9CXDSYkk9GNwTHvCGDG66
X6Ee+RrmO91JA/DF0Nm55rTMjyskU22IBj+mL/ZTH+KV2DvZbxppfzc7MV7c
GjsydM31FpcSstWJeO9Zz5TlYeX93j6hiTHQ1OMspphZfP0/61vSfoU0VMLB
GrvJHoTiib+av1uBtVV8hmL5lnJd8NmlmkBfZlV33pvxxeDSDDruptsqNANW
TwDos6SVRHZi+08PdMyi/CSPQz0X8ZSA49GGUE1pb8KWnvigM/cyv+7pNXxU
Um8xCclyQA77+qIFCGhxYx4kljKGgfsZ7rNO07nnXtMxPdy5XzS/ukxhGTDT
fakaxLVpOKMAgLkLQ2bBVpanprlAf+EG9gJZgur4vwLh6B32IB437z4YwTka
Pf2r7kvVaAIXIm2r3S4llj+3yrINcQ91C371BL2XUVbyqHHGqbFBPe4Lg3Ga
lz4ZPhEWtMT2hX1xK8pf57qd2aWSzOq9I5mmwkTtMW1uUs52uKwinAhnoiLY
vgv7gAh5iOp2a5tY56ACbdlR4hf0byApp33IGgusnpkILdz1+l3zZUtwrAyI
GjVrjPp9QKw7TjA4CBfT5+99dcFMn00ny7tV7/+iuu7mVwvO2T8YO7dkSsLx
2Baij8MoRKual/B07ZFUlmIp2rZ9MszojOuD2kOittkRAfjgedf7NnFrs12Y
6fqaSCg8CGCPeWXZ4Gpe/JseCWcMruVhfe9t/Vtc2NnPJm268Vool3HfoloM
iQmEjyU/11Dtx0a/YdZb3jciYj14YtYu73q/apN9Im3Q8tsjcT1f+des0iNx
OqXiCr60XqeezF/jM8PCE90lRhqPdf/ZPghRpS1eMQnm/2odIP1D9L9T9smx
fWYRwiT6JCFVGomuVNl9kovE4g9250esEZJ7ezccQSk8AiWaDRR74rRog9HQ
I4iYVJWbsBypJVI7H1tzedHWm92xy6dZJMU0qjrXOX6rlEy+nxVgvW2zQugd
ol7yl9J9B4NFzZiCBmEfvGk1ccdYOvh4MaOp4U6L117/SDxrD0NIQ2n5xFOL
FE2eCzCthZHw1H1EIf7jm1vuHHFbCWN8sK0M2y0EE23drjwSkuJShq/wxRi7
os+q2vhcru6JfQAFFdNgKiZ+t9w0XbkLZmtXAyC94huDc8DOGGxFoE3na7N+
r9NygVp7JlYLkvlFb64whUXrDsDBo2QqHg6uWkQv8/YVRwkyD/9gvjD74yik
Vb/MEVKYGG1nA7NB45lbMuyuwmdrf0Gz7u886x7D7fq/TnCGGHfNuYD+qk9a
pjHUsoHr5iw+ShpfvZR11SjQ0olG7MaZ9KBb1+Jq7EXXnKZfdgHeMnCiWhw4
nZmkIm/IlLj/Mrbj+j6Z7cRA5MRtWm/LheHbgQ4tG50QPLLnyWcEBcndlBiE
SoL9mMagBka9za91ARmC+McTtINoX+HAyzACje/rhbFlECSJzvovJfRWL6EH
L/phiTrDk7MzyqIbk2hgQ1wnPuYe5skEf6C8C9Hzu8flv2a2y+cWWEKDABEL
hlJofMlfruT3d48v6qx50uJBDTLA+U1uEBRJNhw4bGqqeGUfe8oxMV4RgGR8
sfrMUcEQS14B1kIUbY+lid7Qj6A0QCg/d/cRCM7hScecbD7WCPhYK5KuKwl1
jVKOciylw4ZQ0o8JPn0r0EOmrwM2kfgZc5PZMe3ziFGlNR7kcqoh290lO/AO
MOexw6qPOXxi7M3Kp3FyYVVj0fUkCpI4cuO7i2hXzu2fu1E2CgJb08WoTRg9
F7RN5nxJeSOQcFXr5niygJ70KMRr4QpOLpP97byrsqgjMjm+c5RSRs4GdNbs
XYcd9vMsO1zCjEHiYP75xggPLz6n+iRNVGWJs8DKQ9dzU2zJZI4UiHh5CYDC
ErvFi8aZKwOOkmnAXTduWhK78ikhRSujqrbXMfiYP49L2KuGoJqgUYm1IatB
2V46AO4MRzFlowYZU6Usp4J1Z8jMwoerlC0C8MSTNi4Gi4uf8UjzpeVr331H
ekT6OiYy2Rfp11/R/4E6v+6RWMVY5J7vdtT7x4Cg0/2ihDlpp63bj2eMRZun
NRyRIGOvGc53nlpmtl1s5OzqFifL5q0hXWkHSU30M1Y9r9yZVXmmTC9TALCG
exfXGKl/rnAYLx0kSGcqXP7oN3HDA/XVJz5y7f5Rh/UFXYnOcZkrjbm9b/Dr
5EpbTt9g33cHY3jxvZouvUx77F39PZVm1pONoMEbejg8rdLX4AFv0ZigokEu
CzYAaI++36rgJwsQOpJN16rCu68hqK5K7v46eJOPSOjh2y0188APBW2l7WcM
dNayb8TSgrVx+xGRYa7JmDY7ucSpMh+5mgi2FbcNxPDthEk1WS//nYNLcS8d
ewBJXQ4K19lBgmOkcF/C/q6rOtK00OOIb9S52j4QlCIvpXYXU9u9XHqQwQPs
lygpmOGDwu9SzUTcCdmE8XLzfbVz2AKAzuC1dz6h4xvbuAQpuE4BEBWX6cE0
0lf0tI7Pf3vDRs/bwjeF5ug0JaeNZ8UYUv61LptfpV+LAobUGqLC2O7dJbf5
KXqtAoIlWa2WbaBeSMpKtX7f9m602SeoFu2DLzLzCFIkReC2Pzqb4/bPpMrg
4eqXQv9AmjDbxx+HVpqNTvinPWUDlqKkqzBiYwRrNAvmncmyyHlv2lL6pT/T
FHrrZnTZgm6ZtmifbUALbmJopwC+gLXHTaOBX3jK9uH1d3JNNKsGqlJbIFyE
gY1H4hXx5vk9iTROecKM11f6JyPwOgnoMCov83xU0oFHSGE1XJGPuUx+9p2W
7nbfLgt8hWPahB5XcFwCAsNnxXkENjHrmG9peOaHc/IM8MVqCzTWsL6e6xcd
pwav8QJhCymPl/NhgLwDXo/No+O6erUQEdfcbPo4Gp3wkCDJp1sP+SZq/GIg
4owY+J552cHGGgYk8FVppx9b9UChjLnftUG/qWNcczpPz/r/xpDzot7S2s6K
7xJY6PQsLJGFhAPsdttOZmRzQ6PApVIQrukhZmYH2kAsA5Zjj6Fl8OtMFy3H
62VQ1lsnX2Ur6ZnSJNf/gxOO3cYDtVOXAKhYj2xdJcnVPP+fxvLVa5WvUs4Q
mPqpzdGfseX5H/OzZv+Bk9XEJYBHnpr2sbN5/SAspmIZ/uyyDVEtGNLM+0eZ
ZOQDWVmEeDkFghEyyRSNQFgKMji2XHw22LzkcxpNbxxvWWO2QMlOX72dTbvk
SAFMu/hFIgKszoYZZ4V5yU7HyMcVyMZjgn3vfh2LlFFsz/Gmacy3F5nj5Klo
pr/DAdd0hAdhxQSSPDDCFLtmuzJJbNICmtAKK0/C2B6xHjzsxo/Wz0gH8dnG
3QmSWeA3L11ESfDyH0JGDMyl2g1oprz0U2GSffRHzNIFm3HRv8obUlTMYCpN
D1yxRL+BO1lU+BGpl4KmjsVLYQ9vw0N+xxArFpgaivMhvRGEfA0HttF1b4YI
uh+LDq5PJ43LgzBj8/tCw17RdfGbOEXKcDBavrSCXwXrvCtGvhPWGUEs6e8C
mn6/9uCoYi3kQXujtNPMORM6PQIBneu73WF4sgfxVQJv8P9FYrLa0s9Hy0Ti
oOtNafe6nyGXZdwg14nNbQgb9gQrsCzCx5oJwlDEMzLKkgycNsrKbQ04Z8Dp
3kbpZnoJs15FEiVA9OzZgwNxUCyqYBh5v/gK65RIaTCmb/Rz5nG4D5JiRMFC
fokrNpF45QhWJyj22ZuW+QQRRxhOMJN1UQBBdeq6i9e22ix4kfHNcnC8AF63
Ub28ICL8TCiyTUqipeS8kupnUQysN3VgCOx94Q0OoLkI0WGgrXuXjjj85MkB
gpuGmpXHQL2yw1oH8mWr3YJX08Az1YNjyHPP2Fi+zMRzyrorIjQse8kKW5oS
HDx3zxDRrEgTA2Y9nT1MWs6pjd5TYVU08Sr2CLCyqKXc7uJGcsAwn5l9GHZI
XlCKh6gNvQxWd3iUdRr2fEe7LDMrYd3tPZQ/m0ON4wUT67kmzKNfcQIXxG8o
7rVRIZ+Ru6MElnyuDiAJ5gQaEovV+sVutHcf/y0HKSIdG/L6IHX4pcYBZc7V
O3tWlXvW9BlCjkH0m0RjbVfQYTEdni4ZsRTJPdeT2Psveod5DDxhmid6OAj2
KQdzlSYu1vuGGAxj0ctMZWG9GPyMdWT2Z4YnYyw1eJSnR/giZ73DjjBLNSwW
kAT08XDW8VI7/jjxhv7Uz8+iO/S2hFQG5jw4vAYfYwvd8LvK708f4qylOUw2
69ZSsEUKmjeukBhvWidIRkEGQykB64uIsdj907hkczEXRY2bkaCtxI7YfJ5V
GdtGdzULeW7TWba537aVyLU30Eq8pKz+oKC+fqT89A+ytQfugDZbEDj89sEi
ckEaH9+CrAiBY1rw7wVAVCy2B6pN/VD022P2CQkTJ9iAQBNBdZYJgR+xqBm0
z7WgJxp0PutpSrIthP67aeNIG/hIUN9+qAeF2v7r3E/rffOoPC6ChGW1UAhF
G96hKLBbyZNLEohd3tBBrzteWU46G53wMS3gnHCJ5PdESenkzRw2goeiL5lz
2o44tMj/UWA11WHrDE/GDfuB3btoBd97CzYYIFycYjdKlz/ZDCjpb5N1MJm/
/tPqLdDfsh5xM+GaE6+EsAB9rw77I9XATBmqdDdWWkDwq1jvSIr8LkTzb8go
yo/KqK8C8Z3wPATjvzyYnpeEKQQ/mtoO0JfllJN/rsEW1dTPEK92V9eiCO2t
OZokweQulyPCU+iIg8uTVbqIgkKvMpbTCWgTk4e4saPxjo8qwT4iMJPPzJl6
OqBvnJodMQhx9oJ0AhRJna+kOj32z2nuLtYAt04tufkzawZkRZjkjhB2Mkyv
ezflb4yu8CYPFPvk4Kwbn1Orx6UQOV/dPG51ZPCxbZg43RITspuAABW8oody
1T6WI8Ny0Vh5b0+KQDgrg3qhiulcQWwpNJR4TUkq25zQ82gARHzutP/BY51S
kuUCKCSc7S3I83/IHdTSy6U1HAqpYUqbPaFTKYtO+J/7C+NSFDO7ib8/DxAt
aylCkhFQc7gkbVspzUr7Dy5JKzqGWsxVn3EcgQ+pxo3rIh30AD7CyM94Y0IT
ZfhB3XRiVK0qLOdvmp0bQ19dIWr/p9ECx4neQJ3+uJj3FFb6BlcMox6Pmeza
8ua4rmK63OSjLS8Kq35+heYYtezT0J2wR1LHLZ39h4iQjtVNhdRH/+AFuchJ
jCHgCXlcBq8piXT7jLn4bMmQ91jlsICvtGZP9ctprCfa6Q2Y72164sECo/QO
dcohbBiF7UU/077VfB5ALvT0IORjccRo0zsdAEzX8pjbAjzp/MeBzRJqc4qS
cCqn5owujRbWoTaR+aF5f4zot7Gzw1Pd3KMMz2VoypGuQq4Pdfsirxkc56w1
aBDj2vhsSmYUYeJrzRswkBNzcJp7uZmS+cEzgRUyW9sEB+pK8fn7CfJXQAiq
FB0zm7Gjiau7nxLAa9oeIuX6ifzSd/SiT2zoaU5nrh8OxDl8euDeXo+k4qXP
OgHmv1IclriPYkngIge1zY/v+ZoTNKIHvRJgoiqnBmam/2cJqFgDJ/jkiaFr
et93266mkr3uk/L4AHDT6NoVoIqMyE3H5aQyGAUeU6ZDwzPbLpe2cgVIJNgq
bB59BLc6WqjvZGqo6pXGeOenNteAniN+zvkBxs3roItVU955mhTTU9rc1nB+
kx5mylF7DEhZAo1XT7kjaXldFN7DaUMXQ9nNooPFjwl6RXGEVskMnfOo6Gvj
XMPsAFkYGsHoHNpP2/f/J0aRB4cosxBUxqkk40hvpmVL4yXoaomWSbiuTQNI
Ven/sRIi8Im8EOfWw770zFrtdwZG89yrz4ScDht/RfbEOMl2Ytm9JORxKRdE
pPQGPI5EOEFJs37Az9Suak0FcolJPw4GL2keJhOadSgMMI2ajSjF4TAp+B0d
IzhaZk5WbXIjb0lTZ4emE8oD1u/oJsqAcOAghxSsLNAMzdlRWCUKSnUKfPa+
YRr/XH1+PYfPES/buBjqUGr1VwdO4aNXSrEgHso9PMcjejwSfv5FoHo2ldUT
Zsfm/BJOIXYIeQtSZ1rv2SNkD6zLUdaaWotZafxAKcS6szMmJrR2vBeTlXm0
N/u6n3PNS8+ypOMZ03XHB9FkatMLlx1eEmoFFB/1DWlpHrXjmbsCdfqwNmed
G4GN+Vt6j4McRLQRRB4pGJFMxd24Ztjg+Hu9reImVMhqP1q99t1qZW6C0bN7
5lseF+9xPRcP3lORcEsM48JC/3ioeCatINCKe1+hlpANjzp6McnLbsWyr2Mn
e/V04WiLkoFV5R2yBbXhytKdkmeyvmAolF1hc/NSrXUef3zy+13H2aM6zr8k
5+3JmLVTnfRYJisK23phMvTh3f7gcdroHTcSKlw0szKJsUtHKFO04DwC6RX0
E42PgPhkXISdWfjtoxvG7Z97PVRXRwhRhBa0sjJZubLUwnjfn+l7qOsazOdp
GTXTNRG+sbww+br5YjMze9MsX8ahAp6Ayy2s7FuM1z1THE+BxEsd/qsBbJbZ
7jW8HhPgR0gI+/in0HyM8rDsamN8ELC4n2V94qgHZkbKrknQcdTAYgYgyZPt
e7r+N1FMIl8+RTUL8KbFpkLU9mrz1s+zC9lpTCXlj9QkzhKN2B84cPY4RHwB
u7fel8WU/2lvhiwM/HgBrocOTz4HZGH+cOj2AhvzdPTXnF6N1+j+7+4FYkBr
7kfoiZ2Yn+IWxulMpmyTZJyfLPStKgDMsj6Sez1FdyzXCMidJIJ+7sSmDsAM
LCH3MloThOQWo/c/g7BFjLNj0S3ZujK/kGwPK5snK3xOrSS06sHvDg7NuWN7
L7RYKeaFiYW8J7HzXMoU8QnMfrEsC9k05jUZndnAsVFN9I2EFHGs7k7thb/E
QZeIl4eD+EgSB8FOQsjsAsZymK1rlWKq+XGXtjBhJ+NYCbNanAuOudtm3Oi8
r8j2dVHOK4bIG1o7c+5uibK32Dhkis7MvJ+Xrl4AgU4Oj6+mwnFhifmfc/3K
ZYLzfjqHVjZ0MhzL18G3ZD6mq7pl9MwSa+31oExYKj7H5k5KMnSVW0odgwP+
QmPfdGKFcQbIl5XI3quD9MIgxLUKIFakvt/FSWwF5SHryqTC53WgYRZJpeta
9145Fqigk9PEbpgIR8otPmDWAARrSWm3586sDBipRSHxkgZlLuk2okKCntDg
6XOvfQ2xo1benzLey1GKTMI9E92v2JIfxiG+GC+eVS5jvD+Fpy1+dujAM8oL
kQ3NIDcbMFe6dOsDNuxp0XZ7kmcFZIqbLS6UmMT8SsMSTPG0JZyOrWu0c8y/
sA1/RK7kyncp3eK2f7OgUBknS63UTa86nvtv0dkCdxsWJ4xuj+ehLiAxIIod
sfk6MGa112FdqM/NhFuo9JvDyKUXh+Sjh4EenFnImzFRjq/Bg0VEs39g6W9U
XI6LNmNlvxcOu3UfGpqckzaD6bGr19zvxcId29QqWaKlWD/dkZGKT4veNGJz
6OEkrgXTZt2QcbCTPWok3K4TIHc9usLTgOcxrOuaH1erMbojGc26CPEddF7z
GCBal22lTdbLmRicuyVMkNiJTda2XLADaH427F5Ii14aeGDpZxc/9dfupepv
sO7h3YshdCBS1+02ZX9zwxaarO9On0NjDvMMT4YNuGpWfGOrKXGeF4TqdsL2
LkOIlxNmELRWnpk1gSqrDdm4I3Q8iOX7tsp/GDy4ug1hccGBP9UndUVOL+t8
IwI1YL6PjfDeVu356he3mSFPKDpog+YqlIzCBsrkDa8zq4olFZE0/kLR9XqB
hoCxo9noekXPvkii+l+iifo71R2oNzetklOY4DT9HrbiJzmWYCJj8bYOem9G
bMsbQcuf99KeRfTSfc9tqoKV7I+CjuUUSVsCD4+YE8rrosQabEkiy+Qp8W0s
Cd0fyEy116r8GI8gxN3GyoAprHg+3gb5fQEnYBb44oLHovGmzBjD3Vx0EGbr
Z4Bmpv4fhzHpcR/i0g1K41pz/bD4DFWEP5qUn6PxUiJkiYayWMmg4G5DwieN
Bl+97rdaNGgblza1LGinG1utWONQEnsrAzQTxDMeSt2EBDDtdKv/vxqrk6LW
DT2SbZKiWeDWsbEPkWURyuDbX5eW83q8N1Mp6YIIke0shFOjUhSWJIYm4vj+
UpjWPdS6dGhbmLgLb0BDENEEKeN8YeC364eT9+byAr8+LojjqNcBF4eCAnMk
6EwKnHEnQSBYNILezJ0qBTChVIGqK83kuBY0302s79ar2ZBl9URt9iirtJVK
Q6y2pfiqvFTz+e4hzBPIDj6uVRPMlidPxWxZNnW33WtowAi3PRH6p73+5piV
CFoeDHDFjfCRaYsApAZsahjywrebO68rM+t3gIeWXIAoj5jBRqdCmB4dKFzz
BGCkx34oQu6GXswT9t0e7ENTnqJY7vCzkmpnvQABgHYIxRAksFGqqjaKd+OM
LyxYHTWzsHD3EM2c6D1u1mHZknz1mY19uhrltS3K76liMe2wuxDatPyGFlA/
+cXPpzreGk7e5mfuGZ2j8dsjpCRKdZNamhbR+chRtiuB3QeTDGFc0CThv9W3
V3zIn71/kEmLxzgpW5GSLWaz6VnGDWqyb2T70+cZbCWH8iY5wOxTz5Ek3FBn
W1vn1e5t6u8BzD+gclJ0d/wUqAIu3lC6kEzsYUbkW9s0c02HLiykkIT1eMRg
cNdzp8kvp3xT1W5c4Dp8Uqdc5sdJRoSwvntXJ5f/4DjBc3BzEisffDbMszUr
lz2UEOlqo/XorcQaQSmtBOh+Zy5k6ygfmeDtqH2yHiwDYWEpSngvcyXx+e2/
M/JA4GnUkn0eygZ9Yq+i7PedqPGu6EFj4lwk7Rt3CKUofDgUvDquxYNdqbuA
4VMKBeCYuD+TWPNuXsN3jUlj5cpDDww6KKSFFVychYtU82pSwzxKHKL3eFcZ
qwd9dQk8hqAN+3rC0Ej0HMfuuR3Op8pOemVl5oIuzHpkcOHlYBaFcnEZa7BK
r/AI6nDWSuDkI6WggLD8T+lQvgR4hIb4e7LKUK/Gjdskq2GSAXNJ37pMR55l
1c3C79kACVu+kGduWmLdNGKrcvETS6B+7bN0q+3Zbo954OutlsHCygLJ4s3S
iCkBfcgxSEDQmEJPugofv5oAAR60yHkbVRCptQEXmGaIMM4YDDZN+1qc4oEB
sLxsRGo0hvQ9ihvxJvuELNG31nLbSH+9+JP6Xvbgd9/4KhQaBIqt3voRJrYx
HE2zR7YAObkd6PXrMfSmwJnbpyuVPItnNGCOpdB6yQJw0YmprittLMxH1kmU
cgfRuvRVjitxAEQY+SMJmnMqUbSy3AnduoZhwygneIHlw0hOeslscGppy3W0
6um/y0lmIK/L3ovBuqYhszfbgQTXbs1ZHFtYpjh7yZqv4NEWm8pLUtaUATwu
QIySVJMhG/mamDe9rY5gQoZaBN8sN2vAfL7Plo3NBz4MkkLlvR6vfhRpN5HH
5xADG8xs6y0O37wWYkm/aVeMtVlHqePkdvaxIXJWAO4cVs6NneAgMYTsEDLu
APwwVdjR1hoqpdPtYo/Zh81n3HoeueVLUgbDtJXEcmSSMZg82O8NDvAjeLpy
HjOyHRfUuRK3clJe57zlI75wNM5DwEx3OWqPgde0X8LnwW5UsvytXZGQVQL1
3UHpIyge4qU/fyvbiC8E6M/brf2LdnYD56/TAFDuD1tmJwGzRHLcDWhgZKu2
V7Dt8Mnd7QrraLFj8yNBU/kl9wGfqEE0jFlc0D9gdfMaVdxocvuTgSgzV5+8
TcD4n9lhq3XskNGfOww+np/KNVMJrWtJbXvNcPsJtwkvw4G2M3PCu0frXu0e
z8htd2lw8ZCTDY4/11habwNpqTrn2OwAZkpheobvQvKxZ0f68ofI0Yh368FB
zvvrCGkLUyWRzC2p/qIs8qWh4DlDKecL+rWsUqk4wGOkdc4xnbFO9LMFIJgm
urGfYEJK+1z7bs2vimqhTNCnjfTggIlWMXG08xpD/R9L63uenfVvva+GdGGq
hFewY3FJ2tw8TZVZgQRdVpHMw8ldLRrOUA5BOHn0XP7PTPOps3WS1gV3ICbx
BBIdkKpYD+S58XbkQurjLuYeW1AyFOCm9L7ZyZDpk7yl5dw5R7AZ1wdAGJY0
tC6Ep3LBsneRBWMUKk8GZ6eoFpfhNTjsUEEeXNG8WhMTVmGFBIP/iaLZbt7Y
KT8KR120UjnqwFdFWpQmBJ/+x1dRCEBQRPJgTaB7T7Tba3wlPuKW9eY8DtOa
So+l4G92RLYrSIEZ8PeJq7XrU7BDnb7X2/X/d85jtkp2e6HL0mzyFmTFopCB
CINocfBor9ax4ehnGDSeocKLW8MRBCw1WpkZoRYO1CrtoRWZVNKGudVkhYjH
rzhvf47zi5b8iLxlNo3lKarRIIzw4o0wSBQJ+NvwijEHKNIsGgzy55isd1QP
E8nv8AWP9H7z2lk08W6+Kq0409bfbQ46hC7DrxI84TiCiDAE/hnxvudrHai4
67KaVFXSQ3Oo73MbX4vtRlKxBPrZtkapu5eMSKqd+fJIelgRgnu8DxFeL2yR
gNOPXjaIf6WFb2HWlLqGPKMKJrxWJeh2rcbCZkJfC3qOzX3QtXJZfswZyt/V
Cwo7oXG6DU5nX/xSaJjXHpI1ip68dF1wJcOKUYiTiWGqORSo77HtruH/LEiC
JOvHNuE60LmzaKApaBSSQzuqQ4ctOxu5z2uNwg6zpYoFWel3gRRAaSM02SYF
kd0nTQUEFXD9N3lnjMgwFlngZuTNZmS0ZNaytkeg91TrwOgFUzmCR/rPj3Ox
/o4X7HbI5EHrleXzxiJVzppIEdgWtuxzqEdpV93hBo41AKKdcDO9irmwAHZf
9bN+3SSqQrY4MZHrRI/5TvCg6Sx/SNhHHrsL47Q0EoO7BwI/3npukPQ1cfB4
7VaMOCdjlsdcEs4iUlFYW7qgdwmNuRZH4q7MmoCn5CLTQ4zvPwJlqK+xEln0
NyoULXC6MOIOnOMF+fYxZRHs+4vrCkDeknr67p25Jt2VUxLOD3XK89IkIgzY
VRNQzHjKYRT5gdws4JJBhUqMNN+QU9PV/dQ35qADm9svUscRPpxjBArSQbqm
1vHewcp1buxE+hU17I9lxCuhqldlw/K8WHwy6vn/tiPD6y0DNnGjm707FQyz
1r8BOe3McbGPFLZPc2n49vpGtQ+1o+FFr+aaQ/x+eA0IbaCwAPwoIXLFiAmH
vex+foy/D5BZMFt33NzoDSN3fCY77+yXh2MENb0H4fFrdp00Onmn/fLFZAaO
Bjp4Gjke51H+lYjLk6XwoEAGeDXaLnCUmtwp/opJZGr/PB1t+Jg3HO7DUs1T
RJqWVBfKxjoMTSiGngcu9w/yGUwHjk0OGKeW66TBs9zlulYRM5Dj19oYnMF6
mhbdCElTb26UkivLosRxWyg/CYzFTjVxMh3OmrMpHKPAOUJwBS3223Q3nUP1
LNQEiVSxhdx/Iurl4oBzniLN37nL83aCVYkwgEJPx0cCMs1NWRg6mFe2imju
hlz5SlliDMWzJWyk8aXZJgq9LpYQQzxU5pmLdmqJ10vcTLCsSpYtNs5HitVx
Eqcmaj2tNbzIhzrHoq/cvBcHGduSdCA/0gPhtOTTvKIf3PaqKQ/FWxElw7ye
/RapjFYESnpXM2bvPxt+Jb5fGOPMH5rHAaWwLfpZj2GRdwTHOHgp9DYCN/iM
a0C9Kbcg1nKX8FYiA0Zhg4OtBZ0+4ewyv/2nwdsDX/MCWcL1EDWTNAIjflpC
1hmMbeySYtuUSnroHniJwPGDKJrk2rQnOBdvg/C+iFCv0UvukZssJRtmLigm
Xeim5YofiOL7BuwIZMCozxRy9yOq+sGGP+43critheMFX89EdiBboTgpowVG
Z4uF6sD3Sv5Z07akUY0/hZSgAqUMtjFMwwkoE2NojhZximDzsohNgzzo6BBa
ULeDn0E+03N51hILbcZ6krI28tQaoumiyhUQHakKf3Sy2YC1WJhC8eS7yfNo
/YLOXwR/BuVQgfzQx1iHXFSgE3jAg9x1NErfNudtz5IWWvPpH9KDQMLi3zYT
K4oc/Rjnf07XFpLaMg5R8ox4ZsGfpgo0QCcCmlte2cN+LLE+3vYf9lbpDcuf
t4WOYwuhyzjwCRtTIzV4opVQZT1+EVF24nSzR/cRzi8UgjcWnLxBFmrBH6d5
Z4RwRLllYOQN7FtYJj3iNPtmh08gbgmxJQwnZT5HwqhRHdNnm0ZrFNWANmlX
bsE7VknrEIopXqtDWYgxZ3iF9trE/dvyG+NCovRG5C65XERx6KknbWoghzuf
AvKeNAmA/JG4S7gH3wCkGMtqbl+4VIXnydlde3ynadia8rItD3jw9isWEYWk
Z1x/7e3NdS2FKlYLuEURF/SVm/5EA/SNN3dFwcdYQf2w1cdmxJCxy1SO0wX2
bPTuy/rCALpMUPgsjTAGpi7V6iWHs5y9bpt4rJL6GmzlLI6ajn3iGooWVvo1
0I4DyFJpHI1XQQRDhN/Kw66Tk8AvQ2EZFC7sS1I7J12UGgGcHFBt+dXoyfdb
SGno2rmtRqYhkGlyh6m8ErElBkhcGW6JnnZGhXilXKP5229fcK85s8lJI8Ou
ZflW3n1Y1vXCEc6cYPFlDthbwjVPuAuN5lo7oHgEnQuONBDDiTp0s8VM5P6x
xFEoT9hAgA7LUUd4m7E2Qw6WAGj321zGlTYSmmg5PbcAvbpe/SVuk5f4jTNj
BRJl0kQkwqW+Y+Ogg+Hm1KYSnis0TBd65+Os91rsreRY5VHDMtXjvJlEgVIm
+gFYzyZK93D/77DSwiHLts0+FqRPEQQT19pNRFIVenpgQuVR0IeCbEkqGYQ2
Xf2l2HgxNS+MbXjNHBdH+h2SE+mKvISSF1P+1v7h4jFTSO8zbrMgoToHZzwX
x1X74xOCoBLArbDW0E9IjLpYb7BzgtObuyplMx+OT4GXikkbVybYCDszFt4A
fWKb57JaNP1Kv9n50nAxnLdoMoPhXRoafZeFDy5Keluf5FLorwHOlmxJg9ov
SmYV6vSxa/i2xceOZ6Y++f5OeJ0aKDucWTj7U9donMSJkPRk8P4M2Ui2NPGm
VdeMWWUTtV9vbdCB2C3t3Zv0OxmQprCBZHfHK6B6I6ifnIhOu9geeTQkqAyW
uNBhZ8DG1Jq0IUIL/xqx4g50Dz9TuyvJ4jqEjgEcmGtUNAsnH+/vJvLq6xwA
ZLotV6EcSwegtUmDffvhIFcYkU4z3PRkYf0Kv48K+zTR8DgLzWeQPAuB/Mzb
vRBbKwetHmRXMy5zo5c6UuF/zZGgSSUEIZDvzNnlb9Eo5/vanejI50Uu5gTc
q1tgajCweyA8KCjWS9n/A97LYdlBFuI3hVeZu+vqOee3vQp1jmdpS0FPGXqP
Kq0VZBO95wpjzovc9Claah0Cq7uhrI//ZZFcS76Pp2edjnKfYXXlrGZQ5s0R
hibvy6FXW0iCSq5u95Imk6avBKfJ5bi1wvXRS65iOHmMcfq/1LPvpnVV6oKa
8DykGi4fcWSguU5RxMNtSfovRKu/l8kuaATjc4Cb2Ga1HHh27IsZLbgWPB28
gClRJ+8Ld3+hGQPQ2xh/ZuFtzTKssSFjwHeXAhSEPWNJx8/qQjwCGcY5zx3N
ctVmRw4L+ZYGkQs2RJFqIXN1blIQFHPvl/xvMQbQvkQH6jiFS09KYCvU/4vP
V2hSFW3lGwnFRsEssyPXoa4hoWfNSTpjM3EXlfPMJpCVpzLS9BevnYM3Qjdu
S4jS0xyA8bgVmDbGovhWwQGVfpw0dFyTiW1M3r3rvgAI0sJbmlfuZllIzhzR
FfMTwbhz/3Bc6Xof09Qicogl1hgimz/s4tf8H8IpDSDC7J7ePTxlmaerZX1C
lyMxl26Uq0dPsi+1b0EiQt3gqWSw0bWA/qst9FSbW91TgunPHw3VVeYC25xZ
UsIx7SWHO5u7oSzHVO16EKXon9wDxwk/4obw/Nqwi1OUXdTVqkty+qZLQ4rQ
U+8nA+4CZZZEF1+IjfeKhWEHtvqn2D5NK281cIHWWFFBwzdANAQMKYaIueF9
sEIMLZLpz47V/RMRT/4/z3uTDB64Qz479FIlsIFu5NXbPDm//yZXT8JYJ6uP
qD0zVJuiUdrVLDZJ/KbVA9UPUXbSTm9OWskwPYQ1eiOKOaJkDmf3TP71cqSc
AGBsxtHjPjIMOU5nUzKn+gTrPuDzL09i8+SA2k6OT7VkxP4wFAcc2b1WfRMY
ZLoEXFgSEU2bVzj9/WGUUYfeL6DA4ipzgGsyEI+9ZxkjwDV7ug0ncj1jij9u
zA7MoknJ9OjT4Dp4VJVx19INExqrgnMbWHjsi6y7ngRqmReHYT9eEOl2+pPM
qDsqbGDJrE3pApn5q/Wi5iKt9VcJJmvS0jr17s/I60ueNzikvluzOjX1vZHa
xbrrEKKqoc+RZl1DBNtsxBAT0byzvx8ByvIN++a2wwpWXuq+MvO2ItFmxmcX
3lUN76+joaOH9dgGV4kXY5JiwnT5IxuTWLiUislePui8B9d87I3wg1/O7aEv
GIwnQH2RtP1RU7IloLHPP1xPy3UV7pvfeuIPrjuHt9RskCc7FM3Yxgg/wcRW
FNWBw50j7BzBO2p52dtq4fCdjWu8NBVPtL5eBVAhed1ajfgOAYi0eDGCTuaz
++xpuus4ErI9XyxKq2G+lv8ZG4Uv4czz40fXpb6NA5HMVt7bsWOCaAdB4Cnq
v2EfvqvT+7dIRcSiUkqFB0nht6tkNXf/Wm1QBXJpxa5SNE3i9K3G8ioUZNKr
9lCAMMx304hBnnReuXVCKFWB5lxd0E8lTDHW3gXJHm3dOgb2leNtoMbISmgx
EXYeVDRJ2FxCUL759a1/Bc4xxGpoxe4pBRj8myhg2RhRb6BEi01Y6h9RtUKe
YGgGib0Xim5nyKbnJQ51ERoAGPZeR2bA9nj3nclkJOxElqZv64pzRTPnOC6j
OX0FVyUcU0M6LQwS/QmWbFTkKrBJaS/iU3trVLd7FfkQh/8cgoRpx1fF+lf9
qSl02ZoXcwea3FqpO4nbT8dejso+ON3bsqTqQHipdA74DpCund4X5bUSAWM6
lzBLwfXIoOxBjmG/ot6WQcrbT1hHYmH6O+WfX3KRJxMP46/S1eq/HX/Yendl
oevJDcigsQIlOqVMDCBdJY0g9xGK/iNL8yx4sy3zqR0uXU+NoJh8IfuGcySO
jRpDnvq9CsLzFX79QL4ZM3YPXEwOieR8nOJsvgU5MNkVjbRVCuUWo6Wa8KkK
TCofg+78Z0PfsEUKFMznMEctKd9FOmI1nHAvm+ydqQKMzsqHAJ4VU/YZMGpi
VzHv/OOdrH+9X0fW5DSpu+QLXhCBQev2eCivUh+MFhPtNua3VOxByhl44Dyb
VjnnZZc5kHB+9BAVTkBnkixIsx7aRYyB9cNZHrw4Ql2ApOsQtyodohBTSIpl
IxggZ3UCJg5jVKel6+txToojp3f6N4UQcW4FheExL0BKf+eu6zO79IqwIIPJ
CwcfwzL0DwqhUGceqGNFCq1PtD86VLgPLYql9W6pIfOZ6IRf043b0x5HCMm1
fjWIitUYkcTZPyOlFfunHHoPT1zOaFuuv0LUWiaV5yTi+dADArKGA4+fKEem
MrNlmAhRF1GbszT/K6xDy5Jkso1ulhcdy2pCnGF4ot+HKxZDfWUXUQsQYT4h
ErkomPa94vYT3Q5kbeqnzBKwE4Ut2T6h914tk+1CAQdw27mO5Dt0h8rn9GpV
+fwBi0ctpv46sF1RwGLy4VCLtGnAYxpnkBCyvqgBEyZ2p9EL0ynjMmcaDw0b
Bif3LdHjDDDBaqr8V/QOBuUdPwNio6JRcqXhMyyDLBT7wi+lu7qD8eTMWS4E
2kM1fcBYtaGxXwBVCPmDLndwBhGt4HM7cYNIRHRSLe02iXAG2ObZMfviLODC
ha64vdJfhUjhZ68OEG5woHF6JQpw3DwqZhZWUcKHDx/0WTv2tDaRQpdPendt
NtG1P20HYB/cFF8gqAQdaWx/V812Iu84bQt8pQ7EZf+btjjGP4QEJ1lhmP5d
j3RK6oq2MWdrrIjPpa2/pa6ibQNsOq27luPGF3a1pxjd0gmjL5tn5oM2L/cv
qhrC7XZ1u2H9ORELwR0Hsd6Rl+Z8r7llhycQHVkS/Wxtk2k2iorKcijpC11P
M+LPEgXpqLcWk0g5PlwNd9NI5y0b4BpgHQHcsZ9+onBREnCwjfKPoxO0a635
WJ5iBHQ+qkJalUTCpfzlL5slCU4/e9cVDGLLoAZtyazSC7ZY0jFcDaCdXm4u
OOumMMSgdKdqqb1epkbb+6O5mB88ex1ske7jPi94vk45S9m5xB0BJ2GR7XjE
m3Ij0u/yHKxcmAyvpNlVpnIyy3Q4msvxdtVcUjXqou/ERyfHMIp/v4H4inTj
ejkDd+81Z7kUuNvedZ/rqAnDFoFuEmaRo/XRanBlqvjGWGVE1E5iOe2Q4Sxy
JPNtdFt1cqfx1ylHwyQgYtXXSo3h6RPN+Y1IzzEtrtIMmETjPtv8eKKQtNaU
GB+dypVHojfnVLHayyATuN4JJR7B+ZGj+fcRJU+0GEF2f65QiyWghysOMcfa
b6/ZN6+WC2xMTyQz8EdKEgLy0vo/SHERWDxSSVnTyAwDJiz51wOevVYW/8D0
oMyKKTNTk5mvvL62nLJAzUriaA/yKOv01SGO+7MxjoknRDfTBQev/A+zjn3f
skOIPEZRSUR6P8orP31Ulkk6RU5CyifpbOPFEx9wLcaErCyB78bdEOc3EJcV
UR4kfgXfudOlfra5mPNVoXi5435gwWePNTvgs4rFSZzzdnOFLXbcEJgkCFxo
aJ8PivAz4Zvd5VGUHLKzT9RUeldqwa2zNEAHDv3QzIYHulLyWT8zVxkgqF3m
zi8JiVoO/WIU/hqgG1wB9LLjoypxgBaq7Dlf3WrBA+vNyGQPBIlhRjm3dSc8
HBkNjEJVQSMFBdlx53VXZgLgeKnkBk1rKHO7jCrlsjl4HNK0Gc/j5dZV+VVv
4ElnM28NIfH+v9lfE47/hEkDF13b/F7t/l6o49mWLMw/ZHBblygnQIUyBLbv
VxnoABmMy210tKZWZqzQ5LN+o71FLA8V9Itqs9ZHaYd/So5UCJsUjdVOUUCU
XbOA3bp9NmCbuC9oPODZywFgN3QyEdEsItIzvQdrXnniM9LpCUB1v5ZYKFZd
8bw8THJZHiKhRb0IQfHIs8IloNB0WvKGTqwOgZOeP4wLITBVX7mhZ081vX4g
N5g42v1fvIaTO8uwWGmZlUoYkiZ9XT9wiKdEmiydCVln1SB/1JGuSB6tR2P1
HJMZDCEeumd48YN0Kr9GMYmyPLrOU6iriW6FhGwavs1q2/MUJFf1ktoOnLt3
HlYlvHCKSTFwUbyFmhwsHjJkcPSBvue6vGLJzNV7oHYwD/6DC3/6Rtr0DZ0I
mxH4JQiPhDh2FwluhLzNleF9iJFK3vbyGXo0E+ukz3aHWPqX4bO68qx8Ma9X
YyuPPc7eVcv968PF0py6qSe+f6xhp65Xp1OQ9D9h/khYXjtI4dPQufxHx12o
srLzTV8TLL5j+EOEjCKNmkL1QpVDucJJV3Nr9jnivSt/SgPhnkLc7Yuc9nPh
u1oTqgUW/3R0odoiT5d5WXX9JeLkXeCXinZvQxPZpD5mnSBU7ipMuOhT558S
4hYKInr3seHZd+HJRcFAtXDicqDzkfhvrPDp6ejvx+LY2ZNxiDEDJVKlKI96
iKW0jErxFGl3PPYeovl/OH6wSlFRNorq0tdiA2ZOhgplBVyALYBzgg7FJEu8
GicipcmlOd3ciYGs1WDl6d7iY1VSSlqhLxuxKDK9DjvyFi5qcpiau2NcL6aq
SslUhoVYT7YhwbE278S3ioUF1ZW7nESfEevfp9koYHtbu8N++o2808arwbY9
YIJHRsRLTYdeeVKgI53ViDjjyKAdMmqIi1wGZ5sQXeSr9dobqxi3j4jUl2hb
C5rnuCA1fYoCZXc761Wlg6nm/Tzm8yBx5oQ5Fq4xxpJqkoY0OBjWoU7iuQdz
s9rVL0yJ+MOUGOcLDXtHaYcTDbytYIUSZgZi7LSwAM14gVHN7aCNghFLs+kQ
BHkwnfZwh8UK1i5m/XZyT7xXA0T8wtOazsx+puLdS97MZUyWevxM4KoE2CN/
iFe4/U9l0PjtvlLJ45MeR2ZvJ5EhgwvdzC4NtsnfRaWPtWnRwN86ak5h3LLA
EXc2Am4G9X6WdgPzraiAfjeliXf5+1jnau5DqJlUuYe7K/kHRD1g2YB+bzAL
f+3JgOtWKgALa16Z9RUFyHmxaGzgPYYymx4W6tVCczFt1ewDML3nM5J3n3c8
tubuGyfjcs1wkdpzWKFEFAHOPaq/+GWZasDUMgHBTkgdV4dVSiwvJyC4C3aq
HfnP2k2qJOqhGg/sg0kKW3UTSrMiMCIwkpYdCz7mG5aa9WsQQ5OfLiBdLfpR
6zsf/Ii7y5B3gMJjS1FI1fJ5uTrEhaPZ5lx4JWgg7nnh7WQzJVjkOP9gbUN7
3vii3dVtwxr3jbiliVgBhIoUc4aC1cx48LnWkcAZiqbyis6lLN2KCBSc1hPJ
sZTFWr7RoGPvoV4JVFZDwjihhoIbHA2d6mWQ3DAo0P+XA/G0cMkWzenhZQxt
KK0ck/v0lcgXI/Bot54WxYHyL4xo7VaFH5Bi7P87r/JSsdBm1pg8vGIqDabv
fxF2Xa12UTWxkfW+6tvDmNqOK65yVm1RitTHNBg56TQswdTVlQ+Yz5/poNfR
+QT6tZbfY2XfhKVGVyy45mNll0rrTLqBOMPStlj6o7UOvDUFUy2hLvs/iTt2
H1ne3CYId1q1YS46Aeft5BZD9M9HeAmFndTi0JDbQPd1qbkCKFtokPxiBKKx
CRtcIMdXerHMI5tQxGGWw2yDyCy1LsqIVv/aalHWhGd3HQKrqk6YkXI336q/
T0FKM+y4GCSbXuBFAQw/rBiovrV4oBradZ6mIFWpZNIUo41hOC/2L7feZxZZ
PN1Hgo07x9Voda/CZi+B+dtSyJQhbewAkUYs4xyB6871nS95MiMcEUoTcv8p
udRQLb/VhHRKyOgVsDwl0eaESfeoXcUPRBktVzSyzaSU82uCQGaeFCGNp8WX
+nbhggUaXWPBYKFu8NsKawSD0M50vyZQKwFlCaGez4oH3zK8JGVJvotb8DMK
jOx6KA31Kgv+vX8WnGVni474xT+iygDDCKT+W2oAYKTUPxLUrcbymlKRbQ5s
76RMUUmYWgov452djTK67lW88QVNHMvCCJFciJOydtPDCTvv+LKHn0mWugTm
k1/tdNfANTqqMyEDUK0Kt4X99xGa8JaqykmQ11aH540H+o9CWC87rWyMBp1f
oC6skpHUDcG2XzslEc9AB9C8ex2s/jeNmyzzWmVYRCxuNrS3jT07/bEn7X/R
5pPzqL/6+EeFeUxouo7frG5dSpamRHcxuQ0RzJvnQGcKNj+HoCBcJ23nhjB3
KRMu/GaFOwZ/F9u90OusD/+DjS4xta9JVzQbJBRNVsIfqyT0OlVDR+RW+3un
Gq098R6+Lconj1GXXNqMaZbmK+gD05l024gDFtM//l9ejRHyqvVcQXi8I8tU
tV4KoXOywbMFgTUUZjIWdDECFQXtwjPT6aFJhMH5YopT0YTmx3C41VYoJKfi
NsNuTfhoQlgSDlZXU6wjLpXGznV8cI7U0s9r3sHyBqchzhPUQ2YLtV4G54ZJ
cyO1oDRJ86pEKzQDAsrBMgeYW3fzvpNDi2eqh/FEmahh1aQNM/5JWRf7uif3
JuBhypYBZx3IGNmNvH+nzAs/XvL1IOjom1tUXZKRrotPK5smOfqKc+hMf7ru
6a89wJRulK2s3JsP7K2TflpJ9uS/YoKN55I6kSKX1rU46FM3TKuWrVsZSKWq
lVwdMjz+cZgu4FKSu+4NVMtf1wLpZ7sEo8uzs+xulp9NLv7KpG9QckH5JOYJ
o4sX0L2K0wAc0hPvg935MzsqGcrzwzJUJO1wvZspwvGLe4MBNAHzRpO9iTbE
MorfObyuQjlb2G/IuOcLcfwpuitoZZi4RuP+HfkDPC0cpL92wbh1s5N26qUK
BDeCGX2WsCdwhhhTAAbWIwFLN/GSyUeYr20MrNUWB5CGuthlNpuuk7C32odX
nuQKdTe6IzjOlJF22MURLohN4Ceu/Ug8G5y7T+n0CTG5jAlN/UyxfHdg/O0w
0b/7XaLNGcITdMN0rKztcqhWFpj5n2PxsiH5oK2c0i2VKXrJjSAqakWyHoMZ
2muFKegodzeSONhZ2fIK377RBN41rzXShIzSD3ub6kTwgOn/SfaXUOD6GX3H
C2aMAu6q74JqRxLvmQcphMW7AJS6kvxdnz244j2OpCLm6teBU/QCs/1XdeZw
nYxDfTOsF7kv6iQpfHyLetblRtlOVOmKq0wHT3/DL/ZgndN+9rt1H+RtiDD+
DtoGu3qomL4d0uGEnG1E8b5+P+JtsMz/rgoSg32pOLfVgogUvFvoN119xMPD
h0Mn6o9Yfhzy6mIu14PArmQDd78F6n88y6lq7dwITUQ5IeGDTlNp9r48IXah
FNxLQ/SEaa5neQO1MFcDp291SK0EgHkvFMFukqrw6iZvS3ZalXkquX1TXYGp
dpZYSgZR9xhyHh3IwO6LWhrC2jA/ZIZNv1vJmdNQsWdnrjizFEiJMxunksqS
QF4xEgNP2/7aE0hnP3p5lhRR7rcgeimVDPsehcXHRneRk7xIZOiLbQ/Uu/VV
bFZrwU0k8+XehYw5MJgdjtLsBhsinDC5vawiXch9OhhCfRxpxAlrW+d7OvYK
Qg19QO0nriTtXXbIamVR2YifSVO5K+mNfQVYi86ru/nBkOcKQUTv6q3Gr8YT
TFGRuEPnjfY2C7DEbQ52ZWkwEyAd2yGD03VC0H8KyeQMHqMOBzjzh40S+CM+
+TzocB7R4dgxFGrEB2YxbTM21TthO6HDxAmsrpWNLD+4b8vbzkZgI3gDGRmP
oJpn9C8UqTXt8a7mJnvWylfIT4KaaGRSBuXJbueozfeZUrG+qUtfp/auQnCh
Ya3vxWbBDZJU3Zsj3i+4BgB88LFhto6Rr0E3RLQH2WQdLk1MJUJ2Jjvf7JEf
BAw0lh0EmFLRDiOKRDPsUGl5DL+Wy+/vXnePMHtUAlJ25OZ9Q+0u8rvTeupl
OhnYnc08E8GD7r1IOJUAshYIIPm1Di8FoFbdTorAywn2K/6dfqCL0hh+R7JV
a3GDr9No/zyu99WvDaidjjFf++wztjZ8L4USxUbwJs4UMj7xLf8L8FiSfWBT
Auwch00whwVGCD3592Ju7ylYCi4jaJs5kVoJOlaIjXKbN+PKYdGe1jQQnp6f
eh4SbAYTKxOE1tX0L+IPvztWLT51Cl2ua2BxXVEcTv/AEGMkNFcs5Bjfishi
arF7VK9Oe1ybNEh+FQPJZOJ+vulufwTOz/qqIaGXBHkGqBC3W6LytiSTmcVO
S5sPnTX3v0PmbihIYWD3mI7iZJd5Xjr0Zv1Y7sinD7DQm+rl8VgOClVZ6Dzn
cpvJVWdizeFnNYs1b0EilF9gDBWXUb6oD08CdU/j74a96XNtYwmHIPgh19Sx
0pnDui7d740SpEqH0eP/DLKQLhRLzI4y1k6PGLy3K4/F+hTALEiCt/UvVCbR
EYXcvqStt2rXyIHOV1TzWaMcyfpI5EmZGafHF7Tbf9pbdWXRqgzAgWx71I9y
F7R8y7ImhN/+wF7A0D/i4bXe9+ZSHAaxmX3ckq8k8NjmCfcET/C+BFP9skN4
6VBmMxC8b3FQ3oX9nVM70jyf6PgClGRNaVK9m1VAIh4yVAiZqaHomRnIl3Nt
R7GTc8bCfwYkp1FYgRTyTfn9gcVMUMvw+ppfd/rA2V2SoZ6y3mKefr5DrcHf
fzPH/hpDERjMSlIYhTynwTNsaMtKpjni0D6XEcsVDrbMOsmN1/P9NCxwyUVd
TvY9jxAvj4AcR7I3mIizqdPY+bF37MPj0YCDarT6dsgNpKbywGX2rbs8FmUe
bcxujxxBg6501OBAE99ivv0UF4dHPqkiTd+usbuxCDhRaZQjdjQbDPSCA3/7
UCsl0pGoBsay2aaGjE1L3gar6Sd1GcdK/T4QkGXpNUx2uAQy2Lr10p/lbiRC
1V5V5f7xOKEjBBncVzib9orEOFlulafonkhbwlXi+jWbduD1KQAbMeFPoATo
IYOupwn9isldzQj6JdOW4Hni7FyDobhsqsUK8dTL1aZ1agy5WbEU2rvzu7GB
7dKeig+BYuc6CtRGVP461EMoW63TSDISv0y89ROYKLXp9MM0aVeP4u+oLIBE
FBM/d+AE+ulcFZ4GB7RnLGish4iaJhkqr0G6ccVLdzyfA9E85g96K2GvSZBW
VEZYozMqB3t2T1kOIq4DtaNp3MjHbaqvUnoT2qSZhdhxgf/9AIwZH9PfReah
zt3wKYjtxbKrLpMfJE4H2pN+LJMV1EArU4SX04GLuQ4LT8mh3fiDUALF6wUk
AVRGMNU5Sfj7uZ8iWWNzaBSs3+sIhPE3cu8/ixyuOb4J5omiEQNTKyGAcs5P
V0A88H35ciWnBoMCNW4eUcMXPlmr+mXUyG0rwtsICZo0NWCdRxUQIbUaM1Iu
SieXFjWOQm0ZwwyeVQMXuRqy3TF412geUuzL2uQMX+OEoiWDEN2yzED+waA1
i8ikhZCF3a3vMWTr/fPgBAOrBG1i476hW1X2TW8Iw3tRgflubkoJXTR4b2bS
Tf61VdqGfwuUebQgWLct+x/ZMcxv+B5AayznrQlFnzzcOjgD+SKbzvgjLiH7
6tF4umt5UcA0PM4XOks0Z615sK9oy0v7AlCX7EXZnB3wWN3XvfzCsT0ehF4K
hZ8rjUMCbofxS1FI61jSwf2tC09bsU41M6Bwpye91pS/xVGbOlo6ONsBDrcn
OZoES0v2bjsiyPsMyrXjShpy+lsgBWd6v9QuqroCJvE8YSR9shTJG20ij7dc
cKOudH4YhCZAYZ1Dy8y9nPMUGhEbVW4qLNW/rYVL/SoTwswmVk5b36GPbdRo
xTBPcnvVYbnPoaOG/30VI2Cdl+CMDNRdOK8vdQJmjf4BLjwK6e9L1y5/ariI
/CUvyoycm9ELK31YfOt6fpnWVcGCojaHl+JJ4G8mBy2LjF9edH2n0w/1g9vN
LAhJuzqtV4jFMdb1xlkczwEZZ7m8mGacvftEUTaI2sidfVsM2so6/1w3uCU/
AHjFN1sbJb7G3o89MePS4uzd5Mzk+7dyKRkLmhHHYFRykHQwsDasflcQ/eYw
PX4qb5vCuHjtnaDjD07I3kGL770rkxr7D1bHdjTGnE1hzn9n6UNwa4lg7Dh3
V8UXXcYBAkvUNCPWGza7TdjwixrGYXVrtCQiugWluyhY1XTYKssqpE5OvafN
FzmSRD9p4TiMkNPQa3cYqlBwFydQs9z14aPgFwHE17tY+34nFe+Le6TJ2eP2
MORjIgr4AwRz8l1PZpXFToFK0l/3sLGhjVWPwsCUxJZf+oUO3FfBAVfzYAeN
2EbkTiouiYUlPPsaTc9OfVxfZMjZqo7poqobSCR4kVFkNoZSzBwvf3tRL9vN
Gw632MHzM6TO9Z+zed5sutmOXjEMI9kua28tVeHBclKorYcIOxzJkVg6w6Fw
lESIL4eMQFR4s1nTO/5hsTXELSCO0BGZ/QUgUcYS9NmIghQWo3NEaaBVTlX1
GSIJ0uB0+5d3nz9JaQNW0moODAyiMybkYXaswNMSyP+IrIIeEGQ77swgANB3
C23EZu/uL2Vv0stsEJ6V+luvSXAPYB+AQLI/sdhRGoj/aOm6wuC6VQNIUqga
m9WoU4YdvFCnUrA1KqcWustz03inq7onoq8rdG8eL0lMcqCHo8EysDIEzcMG
pXHYby4dJClUcnJiPOE2CkabDPZD0mek0cNFFGjp8Sw0jMs8PVEQ9EpaB5A2
A7ouuGZrACInjXW97mgDUA6PMDz8oaORArlmOwZpKfNL43G+Ralai6frzbGB
lY3IFhkgpwvhBrGVzzkBtj7egvAeZUEAXPn9e7Mv2j/Xx/hrJUda/yKfwI3w
9OD5ujcY2/A8mWUPtHvw7MjUhXL1ea/x3NJgrKq/HlVG64R99Za6kmtyh8DU
YfqjZuS1MAR5wBvsQqhqFmAG1n7Oy4kV1YktLT3A8Fl95dQX/7lsCgxmrw0t
NrWWBVmkoBdr8u/JqM5magJM08NOC+TmdUg+hu5OJ0eJHxKCG3zqEsKec2T3
NlyBlUrDOIPcXfKE/mHNd+9lJq890L+7Nwcx3GuA+Zypq5m0b1Gmxru4vI+A
5XgZOjYGB+CJvJE/Sc93oFMbLcL7HAJ4p5qtFUdk6fyLM/jhrdUdOWjKuS8F
sZD19gBH+oHTARB2PAY4GyG8y+I1ZLhdRKmKhx5OY/gNsff05v+v/4scl1TE
Tlk7uuwC/BKvGm99VdhoBiHyXC35YDfG1Oc8sEX4P3oyVwy8qfIJyC0HMK9j
B/EJaP4cHMFdsgrm+HGQdPnF+jRDy/fYQOKZnrEdqjvjwhfn2IpCAkMtl0j+
qNWfs4Nr/AwkN7VX6FkCXRPtAMzrc7wHrD8WO9cS54RKgYNm4oea72tGQ5DF
jyjNKwvDqXiARh+JiAkw6vIhS3tqsxdBq9P/4V9Dka0Byf7FJSfHF0eHVXhG
zkHiHrJjT6Y3zx90jgwesGrxuakrODq1t4cOaE1O8hziXwxfnEs5bIBKrl/P
xAq194IYYrw0WdZs+uJR4YquSLDWk90+1Z2aa3UTCQSZ7W8xEPewykqPf+0U
7aqt1sBDCEK/0Lz5yPrXDN9DDdLx8PYCki6BMAPgtGsPJLHGcRTLueaVShr1
9tXgxGerq1qm0sy7+3qTCNIsq6RuA9AUd5kXLadxCpyk8REy/Jed0iaFRVBt
QlfPZYfKEQQx6CX2oCQClvdvmbfTnRPUoUvIy7oWHeyQNXJ7YX93dZ07eCE3
BlIn4aJ52wG8zGbyi30r7lS7TSlkd94B0kRweBP46DKmo9BNDUhY5ycO/pSZ
7pm/2jzgDD4qcqp/dIbC4MqpKkY+nwoAhG1MVFjUfeP/HE+NcM7RNmxi6lSz
m0T9Ca6b5tYc4s2sIKZX1FGQp5x6ZcCRl2kR0AU7Ww2cpESnLdQCqikpEgST
tMGxk7THI01Vn77ZGX1U13MBGdy6cJevCQgGmPVQyGn3KsUaU7YosDEOyvTV
mZmzVtOXkGosXWSSADBSGLns54+bhnR6r9YNr/BDruk+MlW+Jdlg47lK2mLn
rTqF2/ax64D0LTTjZY4FrpPuQutGS2pU6gp+HNBgIYmCcavETEDjsGRaKton
VAP6/VNmWUFDzj8dtJwPwTlEc8ufHLX7plzZjv4mK0wPeWf2iDmvnX046UDo
eklWJl7xLdi/scOr4rfLDDx0B2NT7CEe/cgP9Hatbg9+e+EvnzfQ94dZckxK
PpjTNO+YPin4iejp74/GlAyHoyEtLM7OX+o9+bW4MniWL59CMo6q0zNOHA0N
qqLY9k/mWUQjtJQ3nvqeKci796DCkKg9549NEPDRePOAh7oOTRn+gaEddKQ3
NXdeoCSzWFr7PPv0zFfe0MD0fKhBZrz5nPsYodC/5s7INdttwRqu+DTa4+vg
jPfrAdWlsuKFpjrm8jwXm1YYfl4PhTLsnsEQy8YU2j2Hjdk61HwhDzmvlBdU
Jh2i4/SLXBq6v06fObn7xZyVPLfjUH/2qA67Sfe/ctcQ9kZbUGY3aoFxnqCd
DGGGtmcrGZMNNWyKXaq/MDLYAS7At7EoF1gp45IWPFkwDyHOslFoilCFFES6
0JvQmP7Vw+6aDCQB9KLFmwdebzeIIjns7bFx3oisrizQzp22ywBHpYUuUx1g
sDJvIC5NsqHIQxFzaXUX2SWfa9Exauj/9O98iYNpSPPRBOsCZuQuBpqODV0s
2GDD/xwgZD6UockQVshfxNTjZODSQ0V5EldwXHmgFk7cHhcJAOUuoES07nYM
eBAE+9A+JYpSrmRlXnPhMe9qsDhaPebLMQCZ07r4g2OAeqgTSWEmMbqkbcga
gdZjLeXqaqhAHwrsJqno9TQ2wqgrQjg+HywxoeBAc5C+AHdTi/HtzzRm83x0
a9Y5AxxI1o/wByV5vghsWNRHw87E5poIr4sDXf59etHqL81Wyk32mJlo2Ol8
5BnJU63BLiBe6kI/29Tix4ycG8KKgDhOJUV277mV7Pfk44O5vBpk4l73rWS1
isFrNvDoR9ZJn8FbhsLDO2GiPqqES2L33vqLVk1KKQUPQSwublWQRdNcWrws
O6PrwffdYryAnICHA+/b7CiJ98mUEdcpfgIVRE0XSsMDZDSOkRpb9BHk5+xy
3Udjf7R6QVLxjMmgrprU87eAptM26YUvTSVy9JbrONgLyubEPpJVOikGS+Rf
9FkcCogVeeqHOZy6EZodR9J/iY2lh/hlKJG6rao2gVSLwcoV1GM4Ry1bpzII
s1OIzaYtfpF3EzB5pxnSFgo4wZZRfLwH3xtbvUxZeNOxGiv+uP+owyxoMsWA
/jdmuzKPzVMaCceCYVavTsEhk4HkCUoCy0NxFHhfoyZ4dJEAWCOkELetUCqf
0xQhqN8aYmmL5VAwySR/OkUdjAUwPxXAVjZkczw8hSg/COmF9e84lYYgirjX
V5yBwD7iz74fOXVwCr5kU4WGddidKT7SQnnGXO0RJSkGRn5olNm4V7jfgOsk
EZqTHPGwDm6lgLu1GtH4Kw+SiXOJUmRDfsJQBb6EGcntXuxCoHWNKq2TMazv
qgQ+7FV4biUGneLH9xwCaU+HQqeCCA/Aai8khDjuuVpqKo5xsPuUVDWl06AS
QpkHGO6nqZ/boGp4dXVtBtUZECnnw6ckgVBObTPQVdJmdMnLOYdxdLjwun6T
l2B2xSxBc7sMmPbt2oP+mqj+2m/+y0kr5pUE0ybkLRnJ43kJ98fqL3CBvkxO
nATPAEfTG2qct/LRsBI1n/hxRXpzWrjhJrhrqbpufmLeqN3MEd4aUW7rTp6B
fmp1u8kfUFqaWtrrfaacQELao4U2ZA2g+qh5NRBGjPxQqYoxMEllkO9j3yop
8EZnlV2pUQbJ7bb12evfuXSauGCXrt0sv5WtZINdUSGAoUuUxHzsjg3xcdXf
a+0wrUqpCdOEBcbeb6SLfS2dHttjh4XhkNkWjhu7QVPNKXMYp4dCSJSaUZ0d
ZEWmVTCcCYvnwfvkcrx+xHDuH2oYJaIkk2mzBESKUyJsC1kyn3QcsvYp16We
eDj0G5QeGBHym2dzWgw9DlGFt6L2mp9XqqOebQVnD4uIf0pIV6FpLVWtRBKs
/MUT6OIv3rRwS1xu0ELlzCclYA9XenNARU46yMDUYRUjqPddc3LiIf0/ax0J
7DFdFDEJmLz01N3W84gi2w1bU4C7uwwRYz05EYHvlZAUuxR3jcpS1id22JJS
WTqJM7e/Oa/HaCiSoengnlpbpOF/YcaWxYLS5xZ+NchqRBhka9uTMuIzYbgH
PWOLw/khIk9hc/tSq3MOd2tUc/IvTvrANkjnpWk0/7+Zw+cbxCyHpNtorsif
/IdhHPdGmIKNLPjuY0i4hvHiGM2ILbDi1VkcGJMTaehS+jy0Ckg1bYudbuak
d+mt1lij7tFcqYKXN5FdgDAadJOY1SfqZoi9B7GRUxQtERiHuBb6bTtJ16wF
jCVg3AT0RR2SeO/Df72bj+M2Iy5+oi/TUVVAbJJbFZ52YZB2d2D+RZhaQADg
k04DtvsKrcnTlYfEG3x1F6yXlXvB43ofysCZGQCsHeBZCJBlzUlK8zpOKcCG
O3Y2YyyleLiRfLs41DJG5sLDD8/8Bii/s+g761s+nOG27XCDa1+sk4/D/LME
nLfzSKDFU/vRCWHDgXwNms0A9HpanIUmHip1qeKm4+2bkNUq6u88KtXMIXAU
n5uK2BYIqi7rPN/Z1hkPC/HDxa2ppBHrcW+oe27JrLHnzUIuYIY1ffDjGcW7
LUF2Htuc15XqZL5SJJdGMN3sAXkBcrYFZ73U74qja8Axy6gWeyxCbdAP192C
Tm4uxnU4rC34A/R9EqMAJNUIRfmGwpWAUJhyqjr92Z9mlyZOrEp/6e+LkvVH
RBp9i2TrY0coLxwHQh36bbG6gCRV3R+elnIsZXDJC9O5pMO6yRmDcsP8qkMH
1NT3U2Q4iwPKe7IKOMUS/yNcz7Fc1RyISTvmh37O3NQPSthgCQAuwdyZU32b
BbBuTboWxv+ew4L3/H1IRy4BgzBDsNGyUuEhfX2AX4xF+aWHmb4lzEtbtvMQ
pETe199pnARshZ5JobJlbrTBZIQS9tIO5TIDYnm/SblE6I0OwoPayxkzzTN1
V6NDPRAk4rpW6xpEWptsJJDwkBj8BQa+mmw5kcUif7DXY2HL0785R9dlu3LM
SV4WdzhT2pKMAEHxfd2K+hQ7Dzjf8j30SQOyKfzc4zJqUnll/+7tJqhBBFTt
OG8TaTuTLxk+nDMloe7cYMQf/sIylRj4sXE2gYCDLWPNwoeqBclV/HRGtI2u
ceQ7visfM34Q9iVo0TDtD1a0llqu+VuranYdAb9kXw8Se+NI3koUMFzow9tm
Rc7syOb91Y0WNXhNiO9SuGCQGCcKedQ1wCwVv08ZO8FJ1yF42rtotViBxZyV
gBTl0gvB4ThNGU/avtfdJnLMH7ICqcZymDh5UYmrVD9klzYCR+dZ3E9eg5lL
pJUKKmkvy+nOqY/DL2eZAAL7Oz6wAmyzSIIiY3EmRbSfApJ9L7MtQA+fUJLV
oSXVwf0nwGAsqoqcEsDh+A3pCKtwi6EkiLrg80gybfIgItRqIWlNAQSPZ+9k
+cyLS2r37TaJKbpccdL2v3q/fQthAK7NW5hfa064ud12frY2YUC8qacfdXhh
BTmp0Li/3Vlb5x4eCEZX78r4cMZ4JAsKPGGn860CDJCBllk41YlGWqSny5m6
qEogia8OJAS9ESXe4ssn6MccMvmyEN1JhXCPuuhM7lqc2m3z9V3bdWIlYRkH
VArwEnLyYOM05nshf2vNkoPqMlu6rCJO+7JuOwr+0I4w5jQ27cc+bFHYrZ2h
OFdqaJPxox6O+Bg4WadXfBH0IMuVCfTGEaPMbGzSgJmWQPhOSsGsQ6Cysjl8
0R7DggeHLvjUQfmm9SYhC3wY7hWMMIWKmj5bYdwA92jUIpmHajmXuFEml3b+
DfdG026CHyrkxuXrJ1ayqpDgjWWOAZxX2aYIXvQC5Da5O1oCMweRfC59pOTy
i8omVJZO2wyE3p4p6DSLAhHLXa6CkuWG/XU/jhl3txEWleQwllKwQnu6zejL
PpZ18N+WfBBnnLpUdAdpkP0cy+2nIxJgbzgbJnpIrkbUTZT33u3Nv3ZoOhBS
R9MTDQrDsRRhzU53empg392VL0PbDg/usD3yqXJiMbGRFz/m+7qvQTsJmjF+
vlrjk1FqECZXDEn5taTH2LCKT9THaX931fXvbywtqeX0NYr3O6Hag2dZcaFw
/8oljVZKDVGgb6sK4Tmgl/10pB747rD8d3YRujoYs6Y5HFaiQrqaVC5rS1aN
yoRWagmlzUBdoatVQ54o1DsjR7GjwXtHsjV0pqx1So3mUjjwwjRus9kcZicE
gpuWznhpsgD/y8FI2pEc9p4DUWreQ23+5e9doPep87E9dx6RuUadOhJ7OmWo
LyRU/+Udbq/Pdmag5XLWdk+1wW/c0LOZWjLfk+w4aMt4reIJipvZaWYpJbC+
voY+w7B1EGxpUvbnUSQ3KhN2tk7QPzVgGfixM/aDI5IHq/5pbS5stjLyE0gK
z+9jugGMb4GCYtHOdiACkPYB4lYsYbwPLmL6BmYjoV1s40HwMeyIiWpqSL6I
FSwYexaP8FE5DU+7M5loGmqAqQElDixPQ4PWUIaBOCHN36uVnMscc5L0NSeh
IVQcXEL8DcB8iM1LnwAS3gXpOGJhvho0v5XnLfdtSzvybgfDlmtAIfpofDsd
37szd18t5TbxU8GiywyYb/ABupCBHofLACPVhZFlRVxSlH2kDviQn81gmV+D
C2JqmOsNjy9uLwvfmdZIl0UBTymjQ7p1usD2j3nSfM/02zbJ0fHg/fV7LN7u
enp5QaWhre3TpFG6rz7OQFnfXoeZ3hzD9DBqs0jbgezoulqn6ou3iC/k/lqZ
qQj7+FT0TG1fkqvuCbizYfAOPv0XqQPHQ/SNKju2wexpSxdGfc13OSBkuxNl
ZCQdSUl567PI4oIO+6DPt6YlhpLrNLM7TnIRafbukV6KZuPykwQv76idOddp
XISmGTR5ajqhI9j1njbordApIJErn6IREmchixE4REXtQGCRBTgZ+xyDipmI
xq1CNfU7x4m3JYCjtxnaNUVwD5RxQP9estWaeRwKe/pYQij52wtPhJxJcGWZ
/YRARVQvxwNJS1bHc2WM+26YCf+1UUkZcHlstk3yTIbZPZIppJlNcd/jE91A
XdHkYivsvMY5b0BPVj9q1N4Tbjeavv1/xu3O3vhHPU9IhZ/CqnWsabAIkQFl
/ksc1iUBGgrNFGksDUlnvGF8xhx5Tf7+WeMRTncVeT+MV/mTs6sQoZx9EbXk
tvV9+GZZo0aldgIVj9Ru3sOSa2kQrgnJWlsh5307LEj24Hgy2UW/trY/sFRW
w9s/IkUnYwNY7dk7zUG3mhW92i+UbjgoslqJ/gPlNfBFDBJ1xmTSKtUw/aqV
Zj4yOEoYLF2vtCt82Ctac5AHE5kXZwh3liHB2vMX93SbVJouwbKpkRMHjVvv
jUtojOO+dAHD4U5CMe9rPmqJ7JtrbQpyL2Xpal2FVV44QgmN0JDNsNoJF6Fp
K6KHLRgvzLIq47PubfThmV29s61dMjfiUw/UAHmtJ0MBFQgDCjK8+mQdxOh9
+kVvpGybUgf/wqHGqFZXt+D+gvS957puNqluOQZLdyFRfJUw2P0/v3/WZVCc
zmf/JQcz7YYG4SzknFmwjwy5pXBTmCZ4R1/lsUcoQJHtJJ5vc0hGc2k3xSv/
za5OrQMvVXNq4X4l885jZ5bCJ6oTMuWg9QLBUqDb5pZGOZdtrkdgldGReO0Q
UgUroxWIY5C5tpQv9s1yiOpf9WDhqP890AguBCrtrkxCEfMRH62gpN3aHhm6
zh1f3uOdCwXhxA154+aGnLaCE44XpOQpiDDsaSHWLNa7ygC0uzG9K6UiGiXa
vP4dEjvyxr+71cGUwfCWvUtjD+roMAJdjyaFGbPcIKPq0LbSWSGpFvYSKMff
GdbJk/kkulrS/rbMPrP42lcZVeiKRtca3ewAl9gN21bMB5nKMR2Om1V8xbma
aKjQj9psRV7zSbNp5CkQ35nJWvh0nvy5gmhj8qXjdeTELX9p+k1ZzdUVAJlE
Te9E7XyREHeBnf5eX2P8mK4rboPHSy+dmrFEWCGfXi31OHEkAK+2OTW9pz6E
ec5hvP3J6NPKdCJz9N4rtnFSa1zkB9iLZgo8CNYEEXGsCwCS4HDjkkNuy+fQ
rmjuS/pURjfnErQ47caewn9MFmWER128uWCLzy8/Q6fSM/znNk/i53Tb8z5w
XzcKME2hFaUPq+1pa35M/TjxvecqPyKdf5zSBxzKOTwOJmdZTjoVRnYsox5X
kKDbRwk6nssya8NEckWUEtUPOUMOG7mp56YBDPxu+J4TElCSKIPf6+FOrrA+
PT+so88iqk+9lfOgr669P8u9WSX5UFPAjIivyAR05ZwW6Y3BFlh397Bd5l13
iI0Kb+DM0Yfw+4FFtMTXFurNZvUxOyyLTNW3Hfx37CpwWAh9HBarXsU8lxkI
I2vRxujEo63Pf9fnjiu5fEKKUspl4hSAd5eXeb6jVyFM70t8PIJViZJ4KbfG
LFSVQEFTSfhPJX5mHdpbopNuamJqWfKZW9t0h23a9DLps+BmLQM5Ctdy+woe
stSA5v192y21nyKdK+n6LcgP61dlv1/3h+P3bN8xAgVqfepZXnO8OFwQKmpY
RiD9GS+qdOdAXD/nG+24lGXXeRHaDZOalvcd9FDLLkp0QgaTpGCVQYUZQ4aw
in48h8WTbpJU69jZA6C12x+yKxdI2LNCp1xoVheLQKWKvbh2IfytDbjU6frZ
oRA4vjZ1qXGpDvsnmSS4sFhyvULAbrnTMsuqOyrWaTBBpq1D0aUKbumtwu1f
o9TXEdKGe+3IXXof5Sx1PlzZnC+2zYcGbTj6cb91HQ+pTEWtzzkCAhaQP2j2
SLsflP6GV0VAhR8ETW+qnATNrNrsP1XZKe6iSW32EPcgel3P7/NxnCrl7rZt
G48zBGx8i6OXGRI9++WUqzbfBoVQmUb2sUIpb+ttKXDnb28VJIT0fQaD5DcQ
bxcdkKD+kfXG8nN5Az3yAJ3VnzXJqj+3HVu7+MmrDsF6ylyFFDUqBIpgO5fV
pM099r7WPwitvelW1APY3j1FL9kkk93RQJ0AzbnO7IrByVVZI/PvMoa8Tb2v
slESvPyNTkOdm3spu+IH3gUoyyZtpDgK2pvcd+pz14Ejh7X+qBKfnpWANKz1
8j8TJ/bpaefoIaUMmMbwMuH+YC2KND2fT7zSL3bwcmY3F0akAVIDMeOO+QdC
v5qjTDuIGeLkq7s/pQ0/zk7f3sPCeajC7VR6tAz3MPVEWUgKonoCyc84NDhP
skkgy2t7dtEs2IVwGPHQ4UYVXlXIB8ak9ry9S2SPsHohQemDHgLu4/JI/VgM
j5rUM5Z4cTqZ6IGnaLSj3MMgh1C/NvDyBxfQiYGVHdBYmoHHhIBtcSeDFIox
nSMJ87FjHZRo9NQ9iGndZeM/a1E7y36RPzoYBUFYiAZXhJbR4FDWOi9fWo19
X4YzzgYcWyPkBRQyPPEWDFawFsQ+C60ZlVBdHo/+nnpAOZxDS6qPIjZ7On6d
GU9Ghnq+5PpHMnyJ0VKry29xLbi2q3ngnAtYwMDbjBazJR18E2uPuEIZt0Dr
KS4AJHznCYQ3oh8Q8tGkkb3DmMoXeGTOJJHsr5JzWUCyOFrPEpRmbmi+Gwb8
bH4aHZIxDXHu9kxHN0oRqUSsUiNTaep8ggeIciLK2YcstJ18mczGo06R4AZk
hz2qm9+6EGQhFaqFITT67JFpziMccDm3n8ifmeGLAy4y7j+Mxc1+la6Q8MFu
4ACnwEiDJGRLEuNsHVqcz5K0RioUTUwbKDExtCsO3pkajiHAy7uNSydjsXPM
N8c+ySTGetd0sn+bEH8Z2WVmnssksIMJmCCistUj8lD9wF6C5+uf/TVRoUww
QfN28UqDs+Ue+JGcdyNgXF2xqcruQm5azoKMTCE7jphARdKqcVk7ZvvGN8Jr
1pA6KBg4/yWlupuBvaFP3755VlX0XCjQy9f1y+E9nTaJaMQhJagWE6Mmqjro
Ynu0XIXJf8rd10qmT8TXI4bCJD5WNh58zOvG2x5XvTbp8Sthk42qNIrfRAme
nwI4Jn0kc1vN7kQZIyBnmAjNx1mP/mJYTRLUdjS5za9DCYvscXAgPSQtcTqU
fVL9xyjhG/cIxHD6kl9Tpva/5280ILrmonRc3wy/vLeTAn5hRMVY0ssJ8AgF
mnOdABZRT7B9BQcGNIkwJ53VICI8QLkxw7cTkCcqwi6w/YiavX8TufcGI/Pi
B9QuoLtcO/3ilgXIV5V+hEchFS1Rnzkf506QgljBlua4gRIbPwbqLywWOVbo
wqCrbRZT+nIhH305or1f2CnS4mnDVWe7TSXNZI4cAqqhm4UoQyn3Nj/XcXFs
FlcD9CGVFS+Lk3Daoj55t41q6uDanvYifse5vG72Q40+h2AgDD5uGIllTtya
tsUIiQ3Qu0q/+l4h5LKxy0+j5Zu5+pSoPL5NButzj/wxF948SuFLJJRWdmW+
4kY1uY1ejZm1ybYQd9Er+AtRUAovTgxPN1OsAJHzMXavyOf3y9GGmDPUKDGX
EwIRZJ1Pf917Xp+iqHev6/BNhfaNyYJV7nQ5oA2gJpO8vz68RspMUYk4kOHS
OKIClrjNCp4fT61/e5IZpQ7rQHA3hVHlAYMZeMnYBvf9yJQX6ksnn+CqtT3J
iPR49gXxcWk7+aKwX1TES0qboOYUSbr2IwpZuRcBxRLxcJNlUftieYfY/lAf
5ES1Dx104dFBW0IUf1Se9FGSrwQN+Ym06TmPhnPzbzylt2ncb2cArJzxyn8s
hSGLVZ1gkaAwrC8Tq3xm2v0CbZqMLOoUih1i+q4DqJHtXGICze8nDAHQLiJB
2Awg76Pf+fTeSlYcKZQdS1dZ93iXS3ymMKk6Q95tRFOT71CMQCyWzSC3ZmgG
A52BY3mHvZnwKi3+12auQHhtIDdlP+xhFzM5cg3vmHP5Van6cPNacJXWc8o1
XHwW6pWRI6uRURWCNBIfjvIooXkc9vxpYFYu6H2I2UpoZuPwUZGf8JsDbH4K
9E/dvczU+hbHs2bOajl6Q7Ya/WYBRdXUvknPOFVXZ3u61oxfgZatM2WHYudT
QxXr6CbSMF4Nkjw2GVsKW6wAEVdyFFDcFvscRIUgUiRLC6fZIiwzXKkyRayx
asgF0uWEtzPksRoGTTaBDc9Ixys9nrRbgSlolNZdNv11tOgJdyDhjN//ZKWA
JAElIvc8ysQXrHQLnNbyDjm+kmM/adGq8J0Zrzd1sOo8B8jFpDem5ws0DU2k
mCS36VKBwSky0E2iBYIgAvCxxwW9WWBZ0t/5ihbLCtRLY6k/J5z1pfuO5X4K
gdUkIHI/7v44murfoWOgh9/8Mlehp1a3HHRGO9DlThz2jZyIOkUT+we27IFC
Dkkw9WpmygX+XvMt9G+Y1lrYqmcWgUQXTM3lEM95xZIwoMauzQNoabYzunj4
MnJ2nf+ZqtRtU0tpmnsfn4CkqDMwJO7pNxqgQFx5ryWZrOlrGMkhDjsXejzT
xVPvKvIIQXsq4+gg3AbdWyDtQip+kBZvTMV8+zO7qz+jkwjA2ZpfOOPxni3q
6ePDFfNqnUxY9XSoLVtWCnhBgA/cQaDTGR1fpJ21bDg2qgoCLUxUHu61fyWj
Ca26kWmcqJqVGuDVpXG2rdeBJFKlvOlkwtkcsoMScaZwfgdPivn9dvsdwrY+
xGiNnXUGCceYXzCjngrpC2uo6slyXYrUV2fUu/BT6UhCEQCoTg0C0H9ZkrJd
JyF2EXGgpW/Li6qXPFGnF67uOnseYnXsCXfq0XgYJcWcGuLAU7tNreAmEH4d
4qcm3WgP43lyp2BInPb+kIq5oLJB+0WEV0Evc+Cy7Q6JpcXPsfIc2PzLORan
yL2D97en84dKCzS3Xp+fisMH310k5rvhZZAkKu9wCORQBlQwkWBijAe85bFe
htfKAaVnD9HiXnXCzzj3BSKbAxpKhD++tyg2+NOzU3MgWLeKWYL1PcYZ0Omy
gWP+jEvbJtu//M3h82UxKlg69NqtuCjsEgbx3F39oJZbUg4qW9CIGhxXR83t
3ShMrA9p77z2Ht4+LjldRw2ezs1NCtgvXVerXqluEMrynEoAEF9TYw4Q3dZ7
7PI0ata8D6U1hQUjRKryUzV+kD0sEcYU8OcqE1pzrlEO3B8l6VryjxlzscKK
SL206hrbLgdE4serk/DNkkhBFbPpLXuDepA064G34t1SLERwqLjOZF5npJQk
lT246/98PTNzpVYQ00NqjWqN14tWY8LOISQ6nhRB9teFe4HusnHY3Dnw4K/b
szRww36L+QpzWtV7vcewTTCx2ZDpXRg7MMHFt3B4sp5Y+tlMZoyroLSvZm5j
LnFjrUvB47MzfpalUwmWcpWOjzsufonPAm7RZbk2aV/8YXSrpgy9ZAXHDbgK
Vjqcpg6fLPAvDypjO9qW4ud9q8gJhNNRkH2CutA9E7C2m9A2IotYo7/eiwiE
mFV6ulcYp+KgSNRRk7EpUSocqG7YZ1RQgpon7Sp09m5gpwr4nj5GpCSgBURf
3x+8vXmnNVkn8VwCGEe6gpcxCWWwz2fZfoiIlQSh6TMDVoDo2NGMNY7K8KSG
GFFP0MmPTWeUIYN+8fBvZKP/YpXZnFm10BGqG3D6nDjlCUh0onlM7vXLoPk+
sGBC63rOcblCI5JhveipAZVV8QjX02wJelyr0NTaNDC001w/0Za45dqIHJp3
rAF2eoK1m6dfzyNcFKZyD2ZGpr30pU9e2rBNalt+5CEG8gTKSN7+Y2PyccT1
AMBZskSNJgvc4BGzkZsJQrLF9Iq3z6xnXUsxO/KpoQJI4XajstPurn0N/hyF
1zcjFc70knhogtiPt9uGQRhlw4hms9calL+d3RQVrZYalTCmUlLgTAH9ouYr
fS/v8Qm5pEY+p0zx+FNRRpO5D7VISBeCBN54+Ko8i0LOBxIxda159Kknp7Hd
9jEh8RBq8OKv+c/WbeZQlMfh/V/plonO6KvwW3qR4/Xmlt5TiL6nv4O7xT2y
EHozuKgDYLIX67sY8cNZlZsFClguNF35SWf1BSHdY5i4GQzbLZYS4LupmsAu
QUa+ku+ypC6SgbdqPx/ZJug7ejHBLiYTcAuT0bp46RlKZdWf9x0Wm+hPGMdm
diglJ8z7JxgYMOx/JOuV/v/1tWtyEiwNxbmbSBsPtt8jfOfy0PoZI0iqJn+I
A7S4BIxvYMMgog0lgy/wiSCHYLsrypLzP4fndifiY5F4R2XqGbURgh9ttlru
vHbIiWFmPOwi06BFW7taPg1F1Y24WQZrbccxd1twvZVjJTqAWaPmO/Y2lM/z
Cg0/IKNq05wZK5Io6jT7vnbjJ2y0lYvyFydjXs3gZCsE1vEpxfc6hu/N/Z4e
H1ALjqneyuLoDyV/rcI9vD6jaznFYOFAXGyMWCITk2LEen31ts7Pi2QE0feX
fnFe1nf7uxHuLixOjjcS1d2HEvaFrgv3LNqe8rimDMo9e6Vb+t2lneqUPoKh
M8nLRcsQATyQr1cnPZk6Ee7rjLieJuitJro0b4u2DtOQZ81/wT68Nmfvn/Kn
PnrlNmSUcCqjcfDk5iINj0agQhECgCXKQWu4y5BS0uU88iKkQxx/hKG+Jvdj
IdLBcn4mQOieAE8ho8K1BfgaejgX0/g+ecGvF57deibR64kQ5u29N4nGrtrc
siABdZC1FAP3f7mRjCHznxjOWrSgs961aI23DUpBSEyUHS3mKXWBZyReyUeM
uG7xbaGUvDppRGRd97TPKYRxjDTFWoOTOinkT14fsZnpH7b9KNkagaiK92fY
z/RG5bNULH4LIwJ7CMVf9nOS5431xWfEhplPZKR3/ZZjqqdcFz0q3s7Xo6dq
3bGmM1ocLEJWSvmSyx8CQ2ozkoJdnFpYeVX9vYzqcasetCRp06yMjfQk1+dM
a+T4n4bEOVaWRWg1GFr33CmPVE8FwC5JM9pBSzX/LQ32pTac2FQECI27ZscM
u1dS0yIuXt0DP5fL15krt9dV8H63MDOuJNTDMzUhOCz7AohMSThnXe6FI99i
Yc+c8HDiZY+UYA8o1itzOuNpTi/d8sdAmZ/AkQT7j76aSxSEYIeITVVBIOed
QD8YQhqvyAxTExWHRsSW/7A9DjNz3qFpYsDOGyvfmJqm/0/qSe4XcZwFm/4C
G1ERmEDXvVCPC5biQSgDcqBCcNSaINhOlUuCdpLP8GyS/vi7mL40fAeaNs4Y
Tq6tFbwH1yRc3uuSmgwbcynRG29AoYx7SDL5piT5bXh0jRSA7ET9/o/JDSos
QVQEKKr8FYTFSpuqOCOuGlbKeipgI1PTTTUY2I+TPisFMJMGFaUev3HjWBW5
fEKsYHmqURsYmjYzYh0HFFb9XMUwmM7rEtSN2HtvJucBxFElgpf8J4T8eOiC
T3Jvp8flRV1X3MzhNKndcycYS/Wkr38PbwPR/y1CS0ftAw4+KqEBB7HOwhkg
DcVkoXVu2ULGVfBO0aJhrV6saqE4glcq+q1tPOBKrV5eESGdh+U6SHtgEls1
schZXX+gzc7GYyKGmc4qeHiy+c+5X51MWKZo9DZNCUyUdaB+PQcV7u3Lv74T
SUfNc3JAI/LgD6ILWufjBB+OzMdZLONpxXNMVQlWUZDvXFLNwaLk02d/iSyM
NGc5nb9h79O/0+O4RzUDHk51VOIU7HV2SEqOTK0zoAFXsWpCaSkMm+ju5mKl
5VmKWYkQI97M+QNk9SMnF6jWGguEeC5cJnu70vGCBkSNrIVIsCox1ianxYA+
7O1fAKbThUZ2n2YAJfwJeRfnqhMtm7r+l0qb63+U4HUkdEfFSyS5Xffm8MEJ
TmN1V6hs2v8uVOFKERUHKi0V2wDQxi+227V3omuwGmBXrmt0Ft8ks8KQfGXw
ZUyJMcKsBYydQ+GgKDTLdYesrPL/+agpYcptlvSnfvXVJJwOpjmMzBnhZfsx
4O14CZDmr+vF5pjjqJKYvx7Tn4DxgPeS4j5BqHkeo5o6OassjYfnbeEeCxhi
YcZihSXmZKOr4IeMkxCsV1PgtW4ixzO7XL1cN1aSIKjnsh7Gz6uJb+2PZI61
eO8kOaKnUqrGGZTBkOFVwVp3gyv4HquyFjrVW4JhNwcuNg6q074J25Zw1BXF
YRGD6mRCdQIY0HjjEMuljA7xJZU7dSWuvz9wN9B461qqOGa+QZgfoa7+CLRA
DXSIvkfrbKs+LT7JOh1KUHc/5YvmJBU9yhD0B/texBTDnCDOtD8jeMygKnNl
oltXFnu8RJjcPmr+Ykx5iBwXJ1eSeS42yhmKJVNBwaq3X1jfjMxusbpyZ/h4
KYLT32h+rZabNnbbGeKehZ8t+SmXCaN3ewmqdtz9OEaO+AUBt2QXHXn0j0f2
r6P+Hw0AyYGNzh+BhGaPHFrc7uWjWC8VfzcbAz4ZHPbXST0jLNR+UtrkcDRy
g+CcVdVxpx7lyBwqINkCo10sz1TItAtIDzBlbPp0IfUxd+3Flgy5Tgg7ehUC
OPk/yuI1ZiEFCJ35BqxZZucIy3ewwn5m0mwSL7YNkMHdeRICesmC4yvewS3x
EFvnsCilSqamgZiR8XbX3C0IjnWoDzn1dUMcjyHRp85AyUpdPA5ZzBgKpgxN
TsGT6jaUn3sf2gU3cq0lKdDiJ8xZV5NbM2HcjWTkzP3fUEKG+9aKYOxkbXFM
fv/QYy3cMv9RsJtYfabtK+TvA8MpZ4s+99ys6lyaTWKT+b67yYnPi9vCS7jY
tMR/U+1/fWLhvXZUWhZ1gK6RFcaTcwNMrQ+UVcSBaup1ko+AMgOOkM1Pel6z
HAaKwCgoncHsAFjqugdbu+GWFPFT6wszMc1Icmpb17fxRJbD3Ps6bvuUmMc0
qEQxgDuwPphF8keEXenK0RkndibZ4LNo2WLSb/aEG5TN4O/0VPcPhZwxt06S
tDxGSIN1WDpWZtlpZH8hviQEXi8rfZY81K2HpJROHILeIzX9wLyYgmh9XD+h
sKRW5S4hpiG4WDSHTIu+BV8wzNIegngz2Nqa0xp+XcXEnwNcgUUpbxPqLfC0
LwGcD5O5VbNSgZYiTFEUcCF7C0fMTWANiEMGaPj/imQeh1tXfLUXK2SiNgTd
i7rexc5K9PxAbhICct6G+DPCeZ3tCUurdc9aQOtIPtKtMc8kxBJ3hpasxEMw
CMbDoE/3Ml5AHm+7INcAMrvaWPsDlY/erG+S98OQx8AylcgP48tyxQbfkAC5
iKP+uQr+YgVUVHAiEUZ/W9UL2j5KM5x3LGPTLuesp54J/CLPWy+hxHahJJY1
IVadyB55iAhw4lYRonByvF+wIuFtU9VK80b/X/GxpxlAg76cGGWlCjCshrct
zcOH9qK8Np7OCyHxEOMj2SWyvHhBWLmuaHSpX0VqUbX5mU8O83zBRxdvkz94
UkUCTWJFSPRCvvHsgo1KB2y3FdF3nQxEut4unNcSljWj/25Zdrc10hVPL5UL
hML7lbxsPqcPz6MoBduihejIEAp2z/BUQT3H++TBKHpfMRMa153JceNtFWUo
XcRvxVm3GMIAL4c+qDxWg94X7qqQzMgvFaU0ngNi0nydzLMmrOU2TXw4Efd7
DA+8Yp5G8a1DWlle4wLI9y2aezOr70Vj4gS4ruLkcle/IDnbrbn5GCV96rDr
jOMEoZSBhYFijFe3rYhCwAA8vQpa80E/Usb53BUgwqO8Mj4QNngXFZE4I96c
VLX227GAgYtaTJsYD7EeYQZEbKS8Qvy5552HtPSIbSQlf1ptmehj7grN1EBc
tQqjLmF0Pw2wLRRs2eVzOcmwrc4hRW1iST04QgnFiSLknSzd0JTH8F9B+7Ed
6bSEbFovHZOFquyd4MmnKZbcsFjTkwBrVAOQos+Wb3PRQpO5A09Ea2dWi5JX
LUi/msGhVkkdKcyHl9qk8g5V9TnZ5SXvMQyKrGncwj5upk3+Lt0niCqwMIej
E99NFCUhKShN9LYZFTF0ds9EuoKs2wn2gZio2JZqOWxNDBY39KZV5VAvC0+8
tQ2m4R5ptKnmlDAiw3iKO05wfzYQbmNNdPD9KgugF2f7Iujdnzwjj28bc9Kk
3wDdQNzwewHfNf1iQX+VxYxGQnmVl4cRC941aAe0kaTOUdYgTShtZ8nGXN0n
TN/09xfzRbsG3WzqF2cxV55umAKNiJB47MOfG/80esGr7kKvI/01+aWlUIBv
y7JTVWbFeE5F8dcfcjQYOw3xSqkyA78iC7Zf3vEpzNcbwIoBvsaBKrKYFHv7
F8XxhrO4KevBViQRw3/R6LxH5LQlbQdAkqGMLsSEvT0b68uupSIKADyu4Hph
4p/Gvq4dTQzDOgw+ffuMazquqBKiusICNCuYsygEXZnk+YQJJDoXddcEun8c
3fUajyJmHSjyROZbqfr/QSVeERT67U4mkmyNYKg2W623KErdRQknMKGKC8Ub
3aVW1IXro9n0k7RvsQSgOqTbRQn7Vu+aKxGCfs27w1jnQazz48PoEfG6bwNZ
BGIT0bFkUWaVSdh/yGPGPcwtcY/Db9IVUJwpWStUg6IubELtPT0oVC3Cwb1O
ZLrsAp8pB5ZKVPnglBUf3IwTaZ+3QEJGZogCItBmSLzm+oDZIPLFVP4QJvT5
7nXX4rlEI7Y3+xxf9JuEZSUa9nc71fLDX0w8Zvr1KiaeS/afMxwJmSLFOBt3
z4b3p1ieOa+EJTOA5LelGhSpzMdHN48eDDqrF0jsc7Vl8qUjUVeVszIABkmh
M/b6PPUtpReolIFbWWVErc7vmh9+5eHqvgCRkGRzYLEbwDnUIStN4188gntZ
bamjUECs5v+35//iRyqOl+ZouqiiaD/giqh7zXxGOrpI0pbX7VseK9irR/qU
XswdU80EAxDMgBFbf7aTeh08K4LAITF3gfICqk8Vl0eMDm1kf1ZI5UocPOKj
7mV61dtT/CI8kxVdvuIGc2ICA0Z6q2TrBPnmJlxVgJXtFf5qD1PGd5wMekTb
yXzHhjOMMFT2GgOcvxU8Rd6dAsE3is9Ki2TirlQTX7MLhE9b0G8+UmMYuHnd
5TRbomQLpKWdzo0CV55KYyJvQ3GkNrecrr+da8b035z+YIVYnL9jidCgENTW
WPgutPTeNjHGSgrY6p/EtY4//ed2s3BBXrYGhUcbiq3oCC2iTutEFRjNt2kF
CwTvupN+WtTkhUOYsnYARPXGXGqEMWnwpgpZb0tM4j9NKzQE1gIV6Q0lS8Cd
67kZaep7aQbNoyRLTL5G2BM/v0sSA796bS8nYq32CGMU2r7fRzfkw36Tw581
GZTcAnMYB63KDFC9vp6491KxtEdrWoG0I2H3ZKcFA0y4jMTprliRjYGTsbWK
9TfnkGUM49PYUfy6zVszONlFRxzndvl/WjotqawHaJPWh3zxV7Uig499NLGq
eMXGyC1ByHyaSiq9aa2uOCKGHb8DUbIrXUb3pdDkrx75c62F3M/HM+kuWpCG
ieL7ZiEHZquIBcLteaMu+0blFKMvQXmaFVCMZgf7lGRuI6PSv0NdmVBLyCAH
hY1wwqpb0LZ6TPhw5g/s18MJiKx1xE1r0WKC4PdXwSfZBASYKuUOn2mt/g4R
bauUXh0Taid4CRAvWyoY5lC3cneWHepN6m/2jzGli8FuBOl9MC/nxY6856ca
V75WV8cCs0slUvKjTX+0SyQH0T9+6yqaTa7ISCOeCSQgC+bVnk2lkRCw5xx9
Y3Xm8/IFcnGg5c9q/0vOx+S2CJBMvA5zBn9U3hS9R5PrEz9RTOZJcb+xrEJn
h2j5o+iQf5X3u33CHp9BKGtoiJk5fyImcCgnk//NY8lGKnCXYNz+TfMrj/eG
Lm01ladORcYpJcfQ8b2mU94tz9+TX4SgjGbYPTVVRWDVe7N3EI/kQQ0wYSLd
4UVqdw7oMGbh2YlVwnU5nxFfDLlFDbyQOK4uVxHp1GVXUJjAhKrfrBPMkVMF
MTj5K11A0kxuOh4JveEAl2Ld89S+RWqiD0f5vZ/7MO+1dME9WoP3tuiva235
B3FEbB2V6LSHru9d++X4xTH0Gtp3VU+o3wbFTMaETSkGNMrrIClgcfSWxPST
iKB0y4Rz89UvRcpLX8L/obKYpHZkKZaTGScDkgbAjAAFx/fShxcJzpZo2ERs
JzhpdOQdJ1YuWgbGGcSdVutS3ROBvKn/hC6dQ6pM2hhUkRApDzSxlLYKUVvx
FCNlOG/Noas71rQTEBOrOIaIzUhNOv3eohiS7vS75S+/bzwkuZpVlbsInecC
CyiriwVN3Ow/o0R7ZdeyM3+ZAZo8bvMowmHNodwTa56icdWpk9erS1Mj4iWO
Ba0yM0CzPJPORP4T7Zj18EQoCOiq+jbMJZYoxZJ+Ds+YT6jPpfWaS0SVjDTB
2JSKSHBXhc6scYk9Uvu2irOBBF8W7ACWJJWaecIGGgtrQcRrgXPPL7Aa5uGa
+aHvLWMRuRQygQuhBA/LmtFlGL/UF1VS6VxpsGH+EWg/D8cKqQGIBDdNtt05
tkEuljMXm7RS/FqeFADc6JbDKUztQcy09lE2kYierf/HEehh0X/vdRDHBGrp
9MjBhpgJFt5cgORmyML+XR3IfkCSyMkF08DIfKeIyyx5Ht8yPcfgPLGcwyyq
y5psHZR378lPLt8K6XP5ZL7IctwdT9aAbp4MfBX64YhOLjMBrySHa6rV4UlH
JfDAGFQZY47OWUOwZGBWrq51+DwinFphPHqGP7sYYittSPblpBN9zEWGmFBT
kYX4Ks8zvp4qPt+UGc/xCLc+g+15d0ICjsmy3mdg4EKix5LIiJ0yFy1IV3Un
mUuYDMUwMhNd+QWVvGpH3p8ilcm0oVQUf8H01lqWjLA1R/O9cBBILLzHi8nk
Q83S1Adiy4y4kztKGQ7QK0Bw29a0P+lFbBjmODCgSu9yUg99+2HWaiGLAkd7
/HroBQVtZdvvP8ujIH5uTRhVEnJK3Gn9/zM3keBAJxuxR51TIGedG6kq/ioP
t5WXoekJFy1SnLCHXP7aTlkoTCjlmmFkvV1rD3I5eFyVHm0Nc4eauoiOhsda
LtqoG9NxLO+Qdem3mtB1nQzfs/72xQ5WLWgiXTby+uDzK/0OoeXmDl/F4vYq
MPnTbYDOyOeScQOBWw1J8cofjojBmmn6DHzXg/L55+BwiEU7mDJREQUdnvKb
GlmhxJIZC3rGcqCPj+e6u46bMA05lmvf0lidvbOgrZhcnWgiiArPlMl6o1Da
Dk8kB1H0w09H6cp8FaNPzEti0mEFeiRTN6iDu3eNO5MXFdaBsl/k4N7EmutO
qSEC6GmMjTmA3pAQ3c3NJkTbG8dg9g3Au+mED3FS0PF9z9iwLXmb1JJ8bp2m
tCxFPHLbJu5Xmso2cgmgQRMbwBUNibG0ijlNBaEG01LzmpPVvsiuBVHs1Esu
gWLf+h53iyIiYHeSoZX64r6EOiSwe4WcPF7GR7ThZIRdzgsBlq/Z0ZEMKsE0
5+wEqx6qKFJcod+EWMzO/bvy24+zSW1D4B1f4e2zFWRU3kIeu2ELTAEriBTo
Gde+fmvZkEEexUfN94uLZ6UpTxfN5oXCSB6PIGuBPc8Qp8yVRbKfD6I9IgKO
eQTRYe9RK2jLIH3aubAekjffD2+9ZtiBzBaqIadfatvk+PGE/lv3d8MdvPIj
HUVgjyeX7rXxxGzEh945qq0qJ0rGvFlapyuKbt+WzQp1n6yCLUvtBafK7EdU
Ois3WJF+t9i5wG626AqwBBwGkyrhUXhBo2U7P89ORJ0IUQJ6y8UBXgqxNmbC
Cb9eXhs22I3dLX1WsldXQZ9bcwFGG64ETKXCeK/QtZV0SI/w0Zd3qjoSLTsm
HauUXJbRnI8yCwnT13qIggLce1/hceteu0sEfVgr4fU7B6NUzs/xTJjhYX2l
odsGo7oaOuoH5Jyp3iGN+UH3bffzseV/FnxPEopuvVKu39XfJTPRJ1bHV8wZ
AoziZSxHclnvRz8jKFFOJp+ZVAmvaRPs/w+B+eKqvdxt8fdO3m3leR1DJq8s
CSWJ0MzMl9mJcfiWbg92XUPfUPj5b0sJVoiXRLPZ5t/3UlE2qmR5tmtayZBD
Yg4jCeevzi3HKL2Qz9lbAwpH6B7d3Lr5Eo2DAFRnU+cXFmdpi52+IAaOYqkT
GLy4r42jvH2F/vkxaPTLuK/X/uGHfdljry8nSJ9vCaoooWiGnpQabP6Au+6o
XvyFf8OH/vRgNR57KLO0Dnsu2oXQPQ9k8i2uVSvdjBxN20eKNUEAvWuivIDU
tXBZjEkXgPHzuhNIL885sXwN3pm33uYGCKQSganYOuEoiK9gUzX/KvgwxDwh
wNeXGCVQauKmd1bI/HGgp0CfPurnJI9khEwhLCGFhkV+ejx75bJPiau+0Hdp
IVb3+/VbSOJetLt50sze0lkG9YQ+jN5SQd7D9XEl/JzsTPqmm4t0ybqAmARV
LpcvIujj+NZRhbCanl2E+gT/uTtsXrjxTGu9+H5pfDybGZMJg1zzgPJG/PWj
C1fwaUh6jx4Y4GfZiTHlq5KWEdByCaVMVaA8Hb0yEo8Qtc1H4Qf/vRo6gDTb
2vD73vYk+Qu7LbFVHyB89p9C26iwr9iIMj4xO4mz39zYxHapqqizg37US6hK
Jlk+yduH9WwMtPdOH7q3V5o3atRgcId3gr9JfglVUxLWC6Yhna+FEe1UDq9j
90DxSf+cIQgsvrC5d9kdPfn0uakNXwB/lsnidd3troHa6dcprX29IOjpd/Od
jZzFNWEOt1dEf+G9Q4e4aiMdIU7NL2SATHFOBaTHGUtC7VUCgO4D1KAv0wBF
r88lOqNyULRzcsWIKzL2kzsYH2cYkDiI19pchJUGqFrnkTEy4GJGe8d3Eq+A
E9ZvWOVW2oXG/hPk1iFkMFiStvGFRnbMTT7LMtiAa2pk24DlEueIoy08Q27w
+fmdAwfqBM+s3t3d1mGBII+0BRo6hlQky4rOJb/sDKerG6LK/pL8kc06Wq8n
ksyoQEI6/wu+j/QVF3sOvXmdqYD1HB4YkRFLTe1DkM+WZXF89K0JiwrgpJ8B
5M0LEqGsvaGf+m9xfQO/C5jxXezii1HdnXxbMIUCXYazWYExantkLpfZxUSQ
ihFQ93OgbBpXgtb3TINrVLrWWziEF3UbClE2PoLEUnP20RdkSnW4QGekvH00
Fps2tdvlIjiHRN+UCf95bZUVnOw/GbBugiUdY5n7h76Kq1oCwwIaF1eKXDzF
F33gyyZFo+QHecx1SlnfcmheXRqexZdoZtqIFmhq2bckM5e57yG1hH0eMZ1K
L1ygO+EKisqvX3UQoDAGxMDFx42wIb2AcpydKhKyP5gJoa1wRNM9vv4r7ohW
hWhGqbknzDPSbDodT4KlQLGeUY3OcP4RkZ+6oy4Ncl1AeMlOdzsit7xiRPii
yeSg2Iz1FYWMeoQyBXnjvhuOUDzXQLyzbXmwELUaj7rarPie249M1drd+ZPd
q0BdNXBf9YVXQ8G4/RoGshcn5MwVXQJkdaSwmiQO2JDyZa2GpuQ5EkCV5ToM
KREalh381R1+Fz7pA0fKfGzZKlwrRVB/sKSlMFA61AoSJrfwVJAMvOMQRZ4X
XlAHP16lJqNwXWZDd2fWeD6Pl5aEOxsaiPFjhCIfy3rJxGSC5Kf2jt8UZ7ap
MHr2QlNFxevXEEfGK6tgLBtNecX3x7qohgxX6UkjvyntPNw4yEb1r5df4wfh
ZaT5qScMbHp+s2UZVBazARFqDAdo1kfp0AhHKdN0t429RxZ8AofJWn9fulXG
FLwqtWKWE8HReEYQbZ5nmw+v/wi5hu6/75rgmi4kjaWqF3Vp+Lq+N38NYCq5
8y18MYyKFPkWC9Y723wVc8HuGCB5AQMrt/7vuJi932nkXcAizZaeXxXcotWP
RzRMEWqK45tm2B2CVgeNZ2ElrVxOeGpL2gERoZX0DoxpMS3ligpcuhh+SjRD
ducws5ZBmgp/fcBvhyhXy/31ZZnx6wWFushWipMfYxNmtNDFVA3tMJf3A3JF
MaYyKDB7DtjvND7j/TZtuqfjWkSjd/t1sAME1E6d4k37duXGIRMQcjS3k+v5
xK/q7rwvVaiDkKVV9pzPzj1afpdGdN3lYsN14paU+Rdoi8+i0VPcWEbSUp2+
8g8VqZ0UYWjqHtT7yZamNZFvNp1E4I89tPYCx6wiZjjNykexWR4F5NW+fgpX
/Uq0YCpvnCBiW1b4AhBYaTDhVQgws/+mzHw+G9SdCppNj/QbldRQbdaOd6Ml
Q2eZLtKx9aK3SbuPJwB+/GBPipSWbbv9LJiVyITn1Nl7hgRVud4LORnhG1WL
6v9MlWx41+ncJnA64Qzb1gxfBUdj0guLJFcSP+MIeN9KyVrS8lgyk/LVp7vh
Si0jJPynAc+vl8uBYDT+MsTtB83d/Ce1FImHgCV5eFjMMxmomhd2WoYnziR7
736fIBG6C7OrF1Kn2kKfiGg15Rx1Eq3IZfjWLwcs2LJ1FKBQR4PafNkCt0mW
5zCNgCPgtQSkpJhTVLb9ghZLsCV+lsLeITgpYUdYSayCS7yeRePLRPNndRbv
2tFc9oFxEwVF3lhDk8MMp5iq0P/RlRp5CfzonygCQOD5RvO9C5g/8heHU1jM
4aEDTybCCqTanm/xmyzo9c/0JxvssmBCj2N0eKyvbRcboFr+ZmRB9oY28/4Y
bS+7w9whfPYpeuJK+jBkkc6Oj7GDsL46CrsSAOLYdNETss2nmNLkhJLuf/z8
OkHsE9iRNtXM/nDt4Y7C92sjJHDMFVZ1jsNCPVqwg7XIAf6wtB7p8p6WzRWZ
Jon1PsZXWNdBskm6BBW2xxeHp/L1EmOO4KAtx58BHkOVLR/UZbgoZL/Sj2Mp
as7SgIkciSjX5e19sls3Du21KOOC+ZBGx36xpGAkDAxP3eH2EnPETvO+sy6z
O3InlxN0Te38hRS/7nLKu18oM7wbDHw0GFaBnu+f4IvJhqpCPFNAky9FxGLP
mXRS9PA+b+nmPvW1ERKaTwOBAoS+VTX+eWpzqmF9csX3sEGYCyWGcl2SBTEd
eGOSdIJM5zWJ25BltisH5WJYANnaWp23/4la33/ZPqSIbpd/mQKmIFkEL2mU
kDEaPtk4W/pCHcYRUPEQ7p4syJhlCaSyK3U0tzYVpsENJOY/x+ssa40P0zcZ
sgyQGUu1yS7PHO/NCX4VXMdYwvZmREe1DolhZzEj9oGQ+ev14gbvW77UeT6b
G+ibeCsU4vjPXmRqd9C0iB9mw9JlZ2QMPNgiHf08t6TS/R1T2LsovcyUZ+aD
XJAjYPfkQ0w+KsYoEcYLWhd3CyMP+DdydELZdWCaxfjlMUe6958ax+ckMGji
khCQedPPqHkASzRImyagltbTPRkKCI28jkOrBwOY8JQai0+/S++SrEcWc8L2
5RKN7eF4Tkjn5JH2A2Ik1iYI0demRGwDHvka+zHnObL8SdctUjMLZIGtdLzh
sqwKHpfYtUP68uqJii5oWbzc5MKBoWIVMt0hNFmyJ7mXXtylsXLqSiQzRrkH
4Xkeo1y9Qcgeq6L4/cB4FCEGW8mL/oyC97HbiemdwaA15YOGgNTvcBWva/Xl
k8NOUX7MVgoTeOaJYMAwV1sfBHpWcMG5PhkWtfHqm4ZbOKy1mkUr67d9lBVP
s+wh7+UpBSwMkXE7+VmN76LeH0iWU+OZ2tcavQMEsLnLPD5GUR3WVJtNj/O0
/dqGZGlCW9OVdQws7FTCh7r3RUMH/qxJrUQdUuuFcZf7rSExmLSfz51NeNr5
Jya0BKD4jqO0ZuYdw6NvxzmWsXtnGU67LBYRquP7b688QqgNTUyp69SGKEze
oBcO5HsEeahcfr/xiwdqNH5Lg/F6c1i6/EkYxCNPZOgoWYHMHrQCzPs6l4Ck
Egq45CDjm0jWlI1hJOguvCBVq1Td7kXC6lBUx96Akdx3mXChH3jQySrQpPSM
LGEOjPiFHWYSgZ3zdxcetsbOlU8qLZ5ssOcDgC0mjm9e+NIITwqjm8GAMi1j
nHwOLlPNBUATTbupHKAy49mQjvnmKu1dtUFDUqEpFfC61DR2zaJGU2gNl15W
Vl/RAXkA8/vneq6NdY5YVH1f7RyFFvkmUtlGinfs3vHOTpZFouTXUn4NNxL9
vwH0fatLUuCwky0OJkShUEVFTiHgjCmboLx/vzGqLZMOVPQz30OMCdzePaEZ
z46jFQ8HSJoleBp9Scu4Zs41H2Fit777gQq+diFgrOijz7NA2DxGKi0DovMk
XU8ev3AFJMHRSxAkEMHANar/kgk9rNg6BmEy7pl/FS1sHaK1RDhBznO3OW7c
ItiBszF1hvK29LQCRIHKYBsjCgQsBXpvpUjse+tX4/eVlk7QZjGNpR3wwTPq
/73g3DIocIp/ZMt+AuLRlSV4K23OEBtt9BHTrc8wmO2YI9yxn4H8zPrUSRYg
/+jTD39XVN1gsX5VWDsLzUjDs9q+QQTkE07etLsHQAq1E52VyXKISgUT2U9P
7juxQwPZJJzCbYE1qX9pBVXtMJpZQvJL5gYtenM9UVwUPSwaFo1QDOn4smsR
WagaIEni2TK1wtZqRKHGNx5cgxQJ2CmYitnCVwcufSCO8wnbojxZm83dqYEf
agWZ0IoSGf6s3UJ7LHBsiMMgCixyOR0Szq//3IhO4s7CbkjxR9k/yhrgHhle
Jtq9YfbcltgX5YwDveE/E3iq5sqdpdSrmJHnWZ2Ky/5iSdGzBD2/NZKk4zmy
83YBnUpOu97AfRV642AxDmMSNV06enuGq2Asa7cVFHyH3j9M6hNZnZ+tLAER
Ns79jo2k67GEXqS05YVZWAL096L/4Z/mkyp+D5VSTtZ7vzzk9T59TJD71Rhp
5KzWtKzO7obtWIvW/WvkU5+4jyow2z7V2NV6/VIm7E/oAde3r/X2tsYhGSlw
6z9P401rGNSCsS8odZ0W9+SOYNWTAO5DQQFRQ7VooWMzrRvjoaltGrIxQxKA
gtNSoPv+IG/MB+CieNr1Jc0Jt9mqzh2Ack2EVtMTyfZY+C/DiIozqNmbbqLO
J/PDHSUmSMnVf2WWVeFNJ+rRLxZxmAJGIJgDfB2uVNoPCkMs0FCHC94qB0qL
+TZZjU1KFSTe5ZaUcYSVKA+8GYzyTTI7YPX6xDgYkZ7peLhliHiojBOFTYKL
8ofs2EXvLlM/5l5z/n+5vGhyYHZZua5wI8czvjI1u/PRD5e+4v5GMsPJa3Fp
lxPcE8vJivaGnBJpKxHtBa/xHIG6DbWj4YGyFPQZsnXcEIsEsiXMMs8w8eAa
nEmqZcJZrTHJ7fe8uVVhrOe58ZQLMYn5X9hmDDYQoky5nY/rBN2Kp7Smx0FV
Y7Fv4bucyO7Xef9bfhxjaX5jLGpb+Cgq/EHytWuJqUPg/vXmEYL58z18DsYL
o+8P4+gvLcotYXVTkEYau9XfDKhrXTaQiWs7fRQmQjzhf3/u2codMB7zlM1U
7MmfZ3dXPAnt+GwqKZgTK4IPjOFMTSGMZh+35m7V9g2rF+KGCUoZtNHmd1A6
EsENBdWUp93bi2B7M+/z0jmYcoC9bXivAqgM0tQoQL+83QUr1l7MbxpHPHBK
Prl5brsQoXtoMxKLlbJI/1Khaf6v0ZkbJJWEsbomlqihJSv0mxMt9t1ESMoo
7RYnH9qCWHKlBGOqWttVarZTxZZFCt9Bd/fQ/MTMCr8N6wPO5iUUxEiDE3js
GweqPshyPXbePdJ2Vq5ipD+B/Ej6RmujS8Gy1fJDLlpbyi1Lv/CS+xTkSwKX
3rOhtCno9ABSvvlRUh2N6RibiOVV92qpBnIoI+nrevldxWgfAIrsePqoObuA
L73GtxMJ3AWLNN0mXAJUwe8eUqv2mcTBPp2xailsmeo1aAfzO9cJLZ/lrCB3
+C7fwJH3zFlHXieLZhMOmKR1nP6cZ0nOQobmz+s6uFh1B7INvnzW4lL7fJys
0p9fEgBoq6Pf2X4H9HkShAQqd971EmwjseWu5gxx28OHefHXFXNWAvgCpyNk
cPG4UX8u1Z2tzBYierEGqBYzRcfT1FjEcs7xu2k5T3TuTlfNfhj9kx8u/pg+
uCFP1VG1u3zyLvmObLrdWBCrfGkMrec4rNK6N4Xf2QP+JBm0mvlBu0VrXefV
bVKHbAmrdtDbPcIibittJ9SScZ637qTNd3/IQc/AxKsbSrCn+b1Dnm8BMVEp
awSmYbfA/wJIkX7MQrI+dksynq1tvGHC5raZ7Vq9ZJlKRQtXaD4VIkH0cC23
V4xEEjakKWESGRf9Phmjre0ulk6M+AEqOD2UrzsO9Ot9t/N0nVmc6B8aDU9d
aa3+ssWrAdvsSmiP4wgPs6p3Rzc+QCWNfrVurcOYRJGDucjnyvFomt21EzX1
NsAGbxd3EGwU/6yXiQnxJFg9j6j72GGPEgCf5QvISM/ivKFRqVPn29nx4v9n
vfB+EvCoGIdNjf0J75jCZfJjLJgYt4t7R2BFUsOu3zFZOyG0FADKlT83i6cZ
XZX3PwuJmjzNAbuoAuqPQB66q6EoS9IbbQ/sZoT9yKJmhpcnwe1DgcP8Sw9O
oc7BHW50qXFenQjDFFupHLvaP0oAIZerOwdzlTnPKwi2CvL/qX2TwHDRMGUS
rz2fl+MCY1rUnpVdFFO9L4LpBzKOtCUTvbtxPzDN1DNml2d6EOa59KZNIAec
Ecnl5ZBFKB8Y9D32YfOUbV99h2CP2TVTtWnrr5TKJBBa7lZavtwpFK+yce1E
NGlHLeS/1117wTl4Evq6i7t9CCvCxYwcGIxMD34xE0TgmUEd2t1T5TuhDyFJ
cKujAbhxXtCLRRvi1fXGQvky/1m6uWjAeihn/64K/DyGBfQ6g6FA4TZ/MNtj
E4gzYE5IWjehs/Oqc5KDsR8ZLJW+rQbYVFSAfm03IfbKC186Sb4wS+dUxl5Z
xYIEizhNFF6w6YeH8F0XAqKttyGMiuiCHaurmNULZgrpAiMjzxZSOyaFQ5Nn
J1lrxrKBGQUoj1Z/gJ4ErxtR2mqAcd0eWuUKe4pnXQBFLNKH957ghzzPYWx6
IDuIRKlD93JyKaL8X33u39i8RQ6kd4SUYOEjWJLKbEVWAHAovQ2PA6IbGKJw
bIfSb351Xf3noF16ReY528nr+9auJH8F+VJYFdXsdWxpEJHnmKiwZ0ebBRfS
mjSHb8/MWe0aXg9fS3kd7Kdzl/CWaf0m9wKjzMU4UXc0XYxRNMC7s9X9gRhg
4SmDKyqk3s6a61h+HYYb/UbyTe5qmAORkib6Ih1y1vIz1UgCtTTzloLPW7tq
QMGegsJMuXpsHfG0auS+2LEToftfZWfroWzbgdSEpht8OuYhqvO1T9rym0Sz
nOtmymWUDo/GkfINBprMRLK7zmhDVHUzI7TZzmI5J97sgsxykw4RmeVRPeQL
9vKB+8KTIdLfTXQPZFprHddXwQ5i0hLgcQGsOQEryXvLdkeqlYDKECz85Uyd
/+MdGyyf5SN8JbLJJpNogZOMjpcyCand/QsGqvEsj2wpsQ2H7H9Rhja7dN7P
olcMPOUWvB5TCpKiSHJksFnS4Xv6jBJTLFYDd9YG7AhunX2sEbvNHIw+pAhv
zA1CXFUfWjOidrgHL/W/1lYb8jrFDJJKfQ8fsOxPF94d4qdmy9lXdxXayu0t
OipRJ3st6BP3dZ9YRCZgqdT509z3p93KAHfeVcdYn8hCSTq30uR5rB1zytWs
PYSbTYOhaiyx+R7CyuS3ZLVg6ugl4FKMZrmWt0Ex7L8PI2vNzpJGc+XpHAsj
2y3Frf9uSd9JDb6iAECeuoSgEfpqrIDgUMqHtAH4PaNg/15oRME9jHAgMDrV
6bLDJOdSKmbNpyV9kaos5keS0ISVgAgV1r6nn/mKMoVgbkEknTrubT/c3TtA
EsxnxzmhXLlZkIzlbCPvij3VXj4US308S7fD3eAFpnwwLIIbgx0rscLFfzx8
B4TXFH1JJJwUqKr7ufK8TQBZVucz2tM6iAnyQuVKM+WXs7S5DdbF/PKGK7Kd
bjxVGUpqe6Ikcuko4+d/xkCmQzPdQwL7+iAWEsT6L04Cgh9kWt+SGWSRmGLg
/G9JiA/N403dWjmcxnx2RAvFUlG2pOeYIaHmOrW+IGWdBFTSW+sbnFHGeJgW
0DKfImISJTxvVLR8XIquQHH9xDevKpqXUVlRvsh1khqIkoXBf2NquaFV8jZO
PicKJNJpmipHGrglz04LU+oNPIePIoerpdK+G7vEOEAqCHIcBDyW6lWhQyqt
x6AUfuPPaszEeYQsTUswnyj6A8wR9M/w9o2g/UaV7588QIKJpbCctX+3X4Hh
ssmfL5Oc8eglFoJHRxHOvDsg5C1382uEqZ21IH1qvSr4MHaU0iZd0VUxBbJY
O/ULabpn3v6SUkthsvtfa0VGwcbQpNho/fgAuZzsY7cLU48caNooMUmvwbbD
8uPK8/YLLzaQVIfaObe2uOfCxWmJNDvF66/tDFW6sSBy336TB+pSDAkituwz
MQFpabuzaeAsMDd4GkNi0Gi5PMIam1qCNnSknynbBG5Xt+guIs1QzrkNt4ad
CStai5AAVZ4RXsdwW1T+8TtMRbhhGCE3sdbrWnjNsXnCu/aNTdz/wmIvE8vb
BGe7/k9y/dICXEoi7COsSkQ1/QIBoBlObnv3H+NNsROAZQXN6ULKUTOI/XC7
OaW4HlKmQUS6Gl5XmE6j6NUJPkQjtXwpJB/eaBLTPiQ0CSS0US5Owi+hYzFo
oFCsQuhXigvV1HoXYqRuw+b8v8pIPF7xK1Jh5OIuGrpw34A5pwTeGu6Thbot
30amBQ6qEx4u9S8Nr6GH24hmnVjssfw87151kbbAufxkdgzPc7bMkC+mkDrU
SU4bRUmLHnVWTiU+h5scc+RvrUoEumgJt+OaLqvnao0DSY1bCrw84/rp/Is5
IIqXpJyj9ikfApWOX3Hlw9Y6YALtCAvTAGFXlMpqli7q9JBP4lxOTVylHOhb
2+FJlO7v9pC1d3ZmUVMzaRMYgmPVzCmeuNYiKTcFgeXdmTDjkkcIoGdFrgS4
XVHlmW7UyCDm8S7CMaToDVCahz7X3Sv630QXs61SZuUdWq3Ib5LbZnwlLh5n
hFnF+vjLM6w5GGo16I1FOS2RBZy0KiKHVsJKbuS6OkyU7TI5T1IS8fXzGDTO
xWKzFTEQ5VOsRrAiI7z4bW7japn3lE6N4oacaggl+cSaVyB9j6EBZvRZKYuF
c4J5Z3auwHm0ZNbiR+oBefZpgApMyzUh0xtxwlO3YUNwIX7Mj235vb9z/sHU
efZ1LfY+ljp7Y2VT8Zqmc37ur9oKht5wELH+tooz1uhNnLCX306ljZFJCFji
fnAUkPxkjsTOh0eMBthgRNKw2fNypULI5A8kKEvKCCL5tub6uiXsQ9lBj04J
nSAEysAAEY+XXch9csZ/d7y0ZNKzM83Xlr5rokTBj3C2jfHX+cLUsB4Ymvd4
xi7uMB++l2aNX1VGVU5u0z1K7AP9qbIErcgFRDOmjl17CStYPjme/+nSXCZM
lq3H32sFflTOsvsO9Hq/plG4PWHE505rn334L4QE02v0mqFetetgy73vFyj0
GGulv5ynEVgszE/kI7ql7tGrY8D86epxJc3lsMdwc1P++ThKgRVnw6HFMfn4
OsDKltNkT62JwZ9xmbeZuxpI8vLS9gv9beQ+O6JlwA7XAv2YuJ951pC2ItNz
92iFA2/UKPLQdwV6OCO+kaT0iegUpT+82sExY+sfBiSBJIYuI+2JNu9NDQWi
Cyd2KyOyKR6R3rYYwWXOVOo5GXyYyB/GPY/lDtcIpBze/KSl9ovl84fu9lMw
UOlM/OwyP2Q7N/Cij5YoLXRrciDIP5LojN2fN9MiC+lEKxeG2LpaGnhowsAJ
yIGhG8nhDyIbxaVw6Q0vVMuTp/1clTqNNiXe0piAi/n1ZVRYH81Ilh3EJ4yJ
K7ae5U0/6a7HuhWM616lYf3a3RJze2hKaL3qFhN6CdHM0MvX4HeQUt+ees02
Xaalq9AQfgfYf+IKTZouizQgbTIvq/+fv15Io5Ukr4M8AvWkO9XYDeV2HYAX
uoFJ2lJeBqIjb/jWv4Z6lR2NVx0Pk9cS0ChO7gS5zJvXbZK2d78xtgZFx8Vv
JK3g2IqIOBdi+7S3TFYHqX8pU0/NwfzxXzWZEKqz6rECJTW/5H80P7hcqLT4
/NX3KHHDesppQLpsk84yDhERf6fvdnv6I6+2XHANo/tWpiwRxC73py0HHFFL
+W18Ld9Fy35vcxMF8Z2KBmxbIOPiJvHyRJIWU8kvtNArw6qpPiTDPvMIAO9y
5AFZm9jb4XGPcTRSk6P+G1aLzAfAiRYyEZQDbIzZdIyX0ScSNYbtbftMxSd0
ZY6cyx4fRDz0VI0spt4j7rRQo8ovNCYKCFrE6YqXpuhKIpAkVL2fERSufQEZ
BpQ6QSdgOq+NIamXhGFr+A/GExRBgUV8hge8YFx7tP8NM+jjb0QeSjhe96ge
qCZkYj46Y00RD7jhyo5Fz8vfcwSUsRE8PA6prljtfSoKIrtzQDoyb5R9pTRl
+Znd/VwqLBdpc3Kp4cBOTA947UEWDJilId0k68CoGW7EmLWerIVbbt9ycB5K
OgkilwgVfAEGcsrqalPZiw9jZp9ow3yoVvhyZFeGrjzeDP+QsaSzOel+q6ng
lHW7oCmil+unr69QZrxvDKmnboDEW3q59Nl5gMEdjwbdm7tSepcwde0zBkJG
3FvoBM9x1SGxGtd/kTWZ/fNJuh1Ck160/WgjU9Rb9g93Dm2qjR263wMR8+H7
/90bZsa3rHf5X4D6kraSBlZOJJDeUl224Q6r+PMI6BPKWA1o31oc/V3iGJnm
iP473pWHz3gAgn1ZUe5JSaj5Zom5t6nrUhabV+x7IjKt3kJpJzQWZUTCMGbl
2Bl95mAuzVBR3x6fRZVmv1WbhKAdfkHmqnKPLOmfCFvX5EObj8+3rjOLUFAt
cXrykvr4b2B+Ylxz7z+9QD41voUcCxAIKAXopaHTHmMgrUH0CBkQgs89gE9C
8LD/gkfWpAJtbPRf2hvcZmneSf0FJOWTaHy9ps9/U6xYcmsCqnFI8IgMFzhp
3J/lDaneqypZZ2ZkoH4K9a07+dAIhQe+UaWKG0ps69lA8QPsrtC2XIarXzB7
84IYSyKjzlyRTpvHQgtluDcWUvusLNGrl1YGvEYcVctN/P+vim3pVHMit/Cu
K0cqo9Z1v0v7KaKFMbZPc+KK6molNfk9+i23s/L08r0WUFW3dpUsDQ0mxmGp
cCMKBKzz/8bXa+9TC2UqGMxvA8lFUzL8GWXOpi/NWICFekbfjTPMNNypirbX
/SdLcsZcJjE48RRUCdRE77y3cQEk7wAAYrJpdPLRnEjZlmH646Q4vy+4laAm
hYJsHY7/fFQKixpju67AkyCmvlmVoEY41sHD26248KFVxFTEKK+Hqab6NNYC
iBBMjVO9zDwuleb0ggbZLBDwK4m2zg238y4EeTsMC5gUx7KAYuJN9CsYRmzG
BX7nQWVSYR3DYrqbqmHqo7x8BHbXE37Ui8Hw3BHj707aOCzWNQDISJlWdRYH
aO4XPprH5pv481pHkXHzjA+8Mces+gkuP13uW0mtNbUFIIus8Xp7g9pAapxM
iUTfYAWtdPVf2H1wSj4T7VJ4l8P5lqC6RrsEDDdCRyDzMHx5sCJqbhrfN48W
mTc5Ce6pB2jkV2boLRWOfFPVhtFtjP1tY0M22gva5oyvDtIWKvnGs/upmM8F
Q0CKlgeZyiuJ04eSoT311Nn8TCZAFA6knpo11OLOiEkCaKoj2XfSdKt3z+SR
qMY1g8zBW054JTNrfw7IQjeKNtPbZb/QtiUKJV9XcDky9J3wqC1HmQRQ/EfE
WXVBqVRM4N2RTqU51Ff32gAWiNZickmLGoz8imQgftjmJtNlmlTa1SzdBxZl
zjQWXaFBogqKFGALqm1NyUj4E5N04xU12pvlK1zZGlEvWsUC4BitNL5rZgzY
PatdObuuZTCuc+SgqlDhT/KqpRCqHnzQ7JjDPY14P5iLlzalgX+0RkjP2h4P
DsVAg1gnTLivNo8sIqUz/OXmAxWmRbXh2078bR15mZ6dHfUPiOKE2KApk6R2
UbLNia2ipep/ns4kQAgEjMx3x5lP5TWav/XsVmChrQdvO7gwevRLXYLgjkVW
tlQ7YskS2nKSFYniW9Vc7KoycMzFwYat9dtDtBoUTgOIQmI7Hz3l8NnhcQOx
AlZRft1Uzd7HcU3rdX+yhoggLNaG+l1ROgTzhcx6kIgbBgMZx5EFlN7KbFZW
jxW8kWNrkmWD9vW+A2tjLsQofDuDD+Qrc4MDQCMa+8h0V30u2REe2rEV/V80
Yi9+WfhZuFhAel2mAC0BFRxEB1GFlDmidHxSz0inedDQ8czzTH0n4+W6mD1R
sKr9dkOfOS1bVO//ZW/PGNED8OQ0nzUSPpWqcYP5M7aG0CzhlCBl/HQfsGoU
k93hG96c7v1FCCY+u2MS+NvsfTmyvOfzyE87GuLVTgW4xzXYzoCAkK/d6LZC
X0S6w+8XG3LrUPjozdR/hTj61DxfB50ft9asO3C0DhnvHD1+qgOCN1bvxTkX
kmp0gmTBY9685oreqoryDbBXxCzM+xl1CUKjgV0aLTHeqh2rsqmt2FnCRY3S
kfP0YS5TCKEGIvFMzPbW8Sx28vbutSnQCuuzsff+Ux551dxhQEeOLiEuksb6
EV6mAXFaFC0KD535x7/7zjTEyCAgnUiCWO/s8RiZssJp4jnHFcSNGASagvV0
PhjZctxhKhZBgWCjUmxuWtcT6YfcDwwvDYUwddujwhP6NFhkXzTSXdKbO6vI
/k3llgUIPqM2vUOxChkXBhVCTpBZ7F1IhiTHbnJxZiFJmbI6TcYlUwzi7PFw
zSd8IfkzdGlCAmXoBMBEIw1ysPMYy2+HxwnPe9oqhS1oSlE9+9Hqkc6AtZwO
fmAgVtSaL3grgjxHsaN/kcwMIWzDrL7CuyAeg60DbLHMQmHDP8FEiwpQvRQ5
WgDQl/O2ZUdqeBnS+nrGF6+Ffu+L5Xiyr02F/5Yk4FEcZ06EizxpD3N2k3bf
UIXAZ6u7bJwjRh06/BUmGc2hMSxNQ7J11C8GM84L4w7CPYEvsQZRPatHJnhP
2/nrTmLQPdIiQmfdTDV91c1r1i4dre11UcfERDPLWC/P6AielisIxlEKHLPO
6+kgoveIJGTd6HghI+x9yMvb2mS150jY4TO7rhxcSZsCCq4M5ZXHdfu4kabI
09KEe0b2mQC6YrRUZdyzRiEXFUCaguYkGBbpXh2/Uwn09VZC6HCj6f1Yxzrg
3umoW1+tKp/8acAcn7+tBVGiFftnJwgB9eRxZF2WLZwUV4rWH75YWJZ+rID0
KoHA7cGGmc0oqm/EtabOZLNPL+4epcN2j1Iz3QOvLodcMel/KYcWEQetjlKM
aL+R8IwIOo25oD1EfUZnzF3I9Uk2u6bWQH5IaiEQWcRKAIcSBZBg/qSQ5Oah
P4zFuddfoaUgbmn9Hu+ZXcZkxjv6qLUYkTLv1ldInXlp+bbZQOhpyLHPtFUJ
t339dgoq4vWWcGDQHmLqrkIh5IDIesvnFdMYTaw+Q7cM/OlOmf/WLmqzhXln
486UqcosbZovKJQRpR3syqYXpQdES8o7t5WcbopUN3m2Gh86OWK+lE7K8lON
j/hK9P0b70BZMzvNkbYKEaVHKIdGyG1QAA6gEJnthW1LjrN8l3i3FLj8niq+
QfEDWcC+uUzImYv4aEuMDZnUVbpcMh9WD8VKjR+ZxsYioU73f3TavaUyiEVy
OCSPyCTYf7PMvf/SyjkYBzBm5H4wPTPTWzfGQh6mX/MbnXlYNkaF03QDe2h0
Mot0uATgyBoJ3/fYk+lKiUJuy4O5VpJAT4w3GzmOH7kFwYTvOMNSkomHBip/
M8R6lQADSuj+/K2GX5k+j7LBKK8ok8O6ErtiJG99uAFLW5VCqQYr9LMV492c
4Xy2cn+NC2ztYJsSbFHhF9KIhONuL0kH6xABqXyGa0YVNYWP/LO1w6ON4eQQ
53BbdJyYbdjoFPn+QHZ+e6sD0q8EJ3jBNCWmIq4wuKQwr2NFXDNMCsMP3+/b
4SKHoxACB9iLJ+UmVOYe7teB1U5AvTqiwY+oJ2SMLucpOc3Y+JB48eJKVJ0V
nrodrmvqLc//VoCkpiGcPmif8E35ugFKHkIop/Aduisow1zONqL+jKF/foWR
mXdKsxLjiDrAvJhpxxpQtlKM8GxDKqFMKR5XvtJJNDQ79OJ2GXtcY3A9aD98
qYfMsm+NNGCIhtvmEwA3OU+K4fCi9r1CvzrRNuQ1GTI1mXiqUME9E5vnsVnp
BKGzdCediIfCCWFSrj4DlyE/mS0c9uhsenwIpRjqteKvkLWcQXjIDuTn1qBm
m+WWd2odeHk/f4VKYtI9JvUl/RpC0xaHzfEEIXmuYCxMQbtmAo2/r56Wqc1Z
l20F7Npwq5nyMnTU+GkUXki33Uq8NPB/T+V6nT7ixgY7paHY5v1TXvDcVn8C
pHLbWAFpzksoO3MLHKYsoooc+tpZL4639AB9N9uu0o65pb5ay3qn/9OuUUFX
zJjWLb887DNNRixOxzcNmCaecCzhUb88hWqvrmH1B2UyrKkfa/NzlnVcQSZD
5CejxZ6hToBB+thjTE7RNWPE1YQO0eKYpNaqAmR+LQqFYA9jRVHZzsziPi5/
ZWpDI5pHTTziIrXczK0KyZ20K9p7Sxo84mPcAtqgS72AalBVy5X2g7jAj+pe
4gexUrJbPMIsgh5cHudWah0Dl7AagEL8K2i67ed56+lMN/fEhp3K+Td+kimy
fGso7UqKIyxDSGIhjE52mD3P+rM3ozhw89EMYjoLYXlMxDQyK5z5pZCpYNgu
weFbCxhpHWLc/xGOHfCSJJYKMug8W8pfnVNJZIXxaM+SUSn//SbxvmzfZXAr
Uhn53enljG28vpgpmjvgZZkvFQpTKorJl6QTypCwwRqgf6nVlQIFRsUFWPls
qSA6qVI6xtSPG5Cb9ZBxvnvxUQDnIgzEpvwunKaVpZWDWxGQDtvvTX2+pSHi
gnqOlaaPkr3rc907VRRC1mo1qiTCPZZmUYfCi64q9+rEy+KbalZodgDgVART
na70wt33PeI9PocNCO5FuR6TBkVAPhv5bLSPjw95psJQ+JvjkddzFjeV7wMK
zo9v0t6Nx/C0G35jbeNDLII30if+lStkAOZlyeA7IqB6mmxgP5PlsmklZH5d
IYUcf1Z/i87LFZZsLm0f3ZBx0q3jsbdn6ZaLWkYvb0ZoNwpRph9MAA+Cxqf0
qI8jEew0xvnxoGTWuq5Mw5X4spfPofFtJlC5Abb2ni7xsf/RDupbTQthxMsv
eHU/Al+qv8E8OBAqN3bdUKeJfcbN+BQO828WDlm+x6yUqivgjdMXBEyli4Y2
tCVxyqDtm7xD6ek8N9cM7mdz4aqE321ONL5tuEN7pfiLR/kXvzzqBL175CfA
cZmhoRthrTz/pHhXeNWFEMyMZTvq7ZN2TjgVT2SzyyZpsfluPXvpT7RUQip0
kQ+Pp7EHZ7wOnKSYTmkm4kKc1OoxhsDuKdnFP7OIcQwC1W5JhE12zX2Uih2c
GQvu/hQcIYYNimc24DDVyomhM0jN3HnvKzlB1UzqUINP16+NDVbePucUBunh
Gr1lvFtsGSXNbNqP2qelor5XlrO5bw2rkr48PYwBQP4259PKaV8Ex5qiA3JH
OwBODYbbSVnHiOnYjhNsVKvBfKPYjUpQt5OY+/lRoKM8JRIMvDbPIPjdaStg
b6skQoUb95lNKE4xzpyukgesW6bO4MF7IJQAY2uX4RL1OvLw//uxp8WFLO3n
dz/78bR3t8+OfZe+iDLVwMwnYezkF0kc/7kbO+/FP5TSFtm/Hc3uhz5JKoTj
87f+RP/1vRJ+e7cEh8XzRgJlKhsRHNRZyU51YNsU7QcIJuBrMJwPYfyqqcZ1
w28iizMfvJfdDl6hvsmKfdx+b92JGiST1Apv2/Le1+HcTmVH1jKih9tJu/Zc
qd+QO2OOF3R/f5L8k82Mifv0RQYU0KYbijDmvus6ujxdvvQw+filwekLXtWr
2schjCThAMSaB9mpZwKQRIRqoc8vzIIRRsiZz3IWn9wrzJMS+ReVllbk30z0
fmtiiEnVM9BoKqPSEFTU4z1U8WhRcRCFr5GfM85J73NT4k9XiZsjE3AOTuh9
kYYxonkz7qLSFrO21fLhjVRoKot2RYfop3DtX34/Innzt9mW8L+g7q4xiBBL
TWgMl7jl8tJaXEAJo0y50oi529lV0YDilcXnBX7hGP0VbpXqu4nme4znMm6f
KvctwetAsJQ4vbz0JYTIN/bSvadQZN65730NtSlQLYSzvoeddOyZCyRK7U9v
BqEcvK4zY08blj2IZSGNe330FqY9AZSJ0CJ478bA5EQcjT0mQ3nqHYvYzCMS
HUjv0OPGeL/ddTsokWXIOY2b3q7coi77gbS9mfNSA/WuLVMt2V808dFn06mk
jYJqT8vNWbGce3BwIrh9N7QkPLSN7P4ZonJ1epAT95IpP2pLwy9ke7kMFnos
NbltLlarM4VunXpdTAS9mhaVLXwa1AkH2/xKE0OsW17S1MwU6cP55UIzHbTz
nVfcry6AIIY0W4ZRujsmz05NxYOJABSRRN7zfgXFHE916PW8o7xBmErWTKkZ
XcNSOyVnCSIdNET750eQOBci/tSgrQG4AJbJVLnbW1wTGyRHLA4RV0o5KGbm
Mn5MnsGsOMPrX0anci85eR2ipUGxcc+9XHA0ImRAFcehubHOk3tN5I4AJWQL
R7JQOpmA0oc3NSLjzlUgKDwKY54QOdqoR8rQI8Qqa4/cSHtLBnwtfYMUAixI
cDfFPH+H7j7xz14u0UG/9RaKYVi12nKlByfP9qHPfhtee0TvI0O2AHHmYzYN
NaAq+6z3iltvvB912VIcqMJ9xDKK45s/JmD13ZcGmBO4VWHsEg4Mkh7ZF9GA
ZQAqwTeiD0M4XArkgYSLNzcvPkkR//9mvaqM8RqhPA6yfWzuLgmZzwuEaoQt
3vQjoILd8tGCfOv59Nvm0umaBSrfiQuOSEPWdgQrhOVWUv01PbXKdxKzYl3I
3d4Wh8EVoplVubyBzR72BjQapF1UQm3Gn46RUXdIDnOZD8cFDHBCZAQKojyO
O9jpgQjYNLrNqtriMcKyxmeWs/t2/4MuFNRwjB5+SV557ye0WKCtc1q6bHgN
Jq58LI/DHLYM4fWHfaypNEdf63JFF511mf919rwzRqZ2qy+mjlWWpYzInIPU
ue6nHWMkWgNdsUFWDKq3X8WfkarpjMpFCxuC4UkqG7VmJIlDTioOudRotqhE
LoBsHITvS01uYLzNW3xNX8okX8Qp9yrdf+jCDa0zjIh95GPeNO5/kBfkV115
kxNVuSIVi0nlppc7wcEfH6fcNUBf8quMOIWael+QQ+/dWRJqasKN1tUEcCBj
ghMkLnJ/ohGlJTC5wXLT1ig5dyCHZvBNIGHXY+AYOd+T/Wi9epYf+2fIynt0
G2DzQ5WZ1xU7DDt2neOVXLXLdQ692TVSKeG+Rjh2o5328K76Ny+KSoQnsRKG
Sn2IecibravphWp+4QtRLZWnHUc1gzw3dhp4Aph2Ip9UL9EKMLgvX36/Sid4
s/+/5AmAE8UeIGsy8ruc1lP93T7bW9imU1NQ8Qljb/cZEqryQskCYo4pziGW
qSnJKJI+qsuT0AlGee7eg4c+bW7uyUTj0gQH7HMWDlsIPlJVfR1DiaTgo8DX
EOI3foMfjwpgw05NrXyxOkpBNgShqQJvp3y06wzNGn7/D2GiKBNqu0CxZbqa
VLKlE9Xbpedj/rU74ihaqb/k//6ov5Bb3lQdLwY5P9682RRJWPxQuhgYHuU3
lVHomRshikH8qhmpa9rTJPyHOWc+VQdhV6WJyHEdyu6ge55G+Sk772z0ZWFE
Xmgn7UD2n2xoiAFXRurM0RtLO0+vU2zmugYHnt+MiXXCf733X+bFhDaoO6Bl
cUu1uKdKfxOcrfz7WeXTOMh+Gq1mtTN2byKtQkZPmGB/ljHZ7rF/JrF6ipr5
pJBA4M/XH9xEmNKlvAgH+B5/u1MKgFHcPZniC2i7sq+17vzYDvqLoS/JGF1o
IlcnOP3BQETcPx4h+13H1xrDC/KRh2pV1II1jYluMFByXk2qOFHwhWV8gL7j
b0dmI+XuBkQaYpFCbXUMNoHjD4tw383rhqosJBWklVgj50y9zCjRGnJkumgB
t6qDRT6z+st/9p57hUi2lqpWCoBFchkY4nVm9XymPRp5qDlf12s6lPEGgl72
r9A1PbRlk36+162Ijc2WAqY1RXLy8K/6po9tUU1Jko53YAy+exDuMUd0R+LT
T//uCxYgyuZ1RGteJaue9f5Dgc2a3pmJ1t1d9KewL/KfSdz/j36SomxMMvs+
xalyjYkCq6Uj9hGC9twG/uILrkgt7YUh0FviHI9SgD2t0i4vO4MIkvY34ghU
H1IEK9KpJkbsHycxAn1/Coo8E5LSI5AQjxD0/PVEofvkSLq9cQnUmY5+GM0J
9eRine5ZDFeyLWHA19ZOWDtwKu3JoT3OT9NiquaGPQOoaE93QvjVIDY6Tztg
fzFxXqtqJMz52e7jTwA8JnUdRNtG+ELO9zXngXXAalZ3SfutUgX6YL6YcUnH
Lf6xfMg/eiHWUGCinNLeudBW+zeyuqqooM30eH87XHTYBjuDG0B3I/hn8WBw
/ra8eKqfcT06f/8u0J80I4TCeViqbMIWwVrtlqITqRzi1XZ8wRqAhhJzH8hZ
jqfaw1Gcd1Rk0D6skFneTcxNxW/PcTEVf8Mxe9XluzBKq1FP62YUZrfdneNg
02ZUKtygZUDqBgMuq/f4gtZ+LFSQSzhbNGPkr+SDrxqgeZMC7pAKVvgjEw1N
6MDo2GttPc+VCzlD3rEjqqAo3o81qLSp/LmC3lWY8dq85YgaMvIAMrate1jE
n9cOJTPnVrJ5WzpUVVSaY7DcmC3DpisFabxgwYvsxcwBZKorb/cNrF+7WOGQ
IMGyCpuAM41aYCpuFoS79/BtyJ0ogne/TjQ6usAz9QC57GNPAXk1JOVnPA6k
Zuw+BAPaQyntVEPoyO9dNlh44lZVai+pHHboK1XXBqT0gAfaCl2K/v7sVLio
lQMtHHT+/zM+KzyX64OXJzMHodewTVcSjmLTECaFSCllX4aXyqzKDzLYkLBE
5YZt4PfqEOwQDkH4ISgRtbpy1ihqyJRxzkBU8QQctygWS/qTifo/RvXhZ489
S/imGqLpIntM7tzl5Pc8VKFaaoXOPB8IQnhoBVjelEdx/nlk4gF6OhyCOtdJ
QyQMNc99LtTHeQkUMoztOspvF8FMaMtA+GlzNkMolu0+/hqESHSuT0OaOmay
yT3uYBxyhLDSj2Y0S0exagw1qBN9oUL4+XNB4kWz4aJI2Ryz1Td/Lx7icpVE
yGNW43z0sSfSGRqo0WGeXS28qM3nb1p3HeVa3ajiZevYLgYrPmNxGFmMqt2l
o1FYsvhoXmRUqrahQxKrVhYkKNnJ6i1i8MWBuFDv+vntvoY0FQWF4WfsEn5g
sRRciUd7cTtcOUOgBZKaWA2FrSEMa658h/tZT2wNqRYwW3EieuDE7b4CkA+y
/mgq10f8Ae0BJoDfsbnGvwg83g0xOKuAnAj7en4uIeBfu2RERnw9mU52kgCa
fHpacktEHV1NII90J5VMyvFk9NdnMW5oGEjDd/8Ko88Sm931T7fn0SI78lhi
rqh/0MUtWJvrHQseb0Gn7LX9WT+IQNdzHO5jl6oLYQO/RX1fRjL55nr4kt2B
u4gHXdoi3AS2GwI9LuFw1KLv1KDNKxZskDCzmgTl8fKySG1GiGWlFVpbscKO
X7mfShR/weSyZcYak+7BXqk+uLdqqp9/39apterKA7vZzdHtTRM/+cl/rABO
2sOv841joHtKcu6jkoNhwbJeJFDixVVrdNpMP5dCSI1H8lpQubJ+agEegbad
hHw6ybNgraFvsRtAyweKghCtUkHE1OB/+zZ4dFn+BLi2vcskJ9utIxjEijpQ
JeEre5iNWr4EhG2yvzpZtl0FM92RCIvLr2nHAV+eLMc0cAjPMTG1hNpiYEj7
othGYOm3tLVPXpiFggFt2McsxG6Rl3PX4M8ulFOAdS7zC0pE+rpvEBkdvU8S
FPkgROR9MfvrdLTTraqcRn5P5ayuZIVWZ3jLuB8dhtRY4Y1hwNVm7HfMfDG4
txQh67tcojfrtqbM3jr1x+OnpgkYx70/ucGFZdNpBSmtO5UI+zV5gghdttUS
VnkC9KDEYdQNnQB6fZrcvWFs2aqZVxc9OogacurFOgAnGlcCGy0PiwxtvvZF
s3QuTo9egHiAdjecqqWN6yi32UFGV9Ingqf0V8PGY6741OT3KcewWQjjCndB
A6FnP9bjOgY55MdZvfj9vu7Yfp0145Aoamu1hw+kTHHbLoE+g+Kk1d94qTGP
GaW/+IT4o2Z1AcxQ/5jXDFlcovef386giZ7OIBC3COZapcEmyTdZl5AxseKJ
kpYMvp1FLarJlD4foPH6U0EE6pxLJ87GKdfkIaz1nmDyAQ9/7etF5qjZbbvw
8AROJqPlmVG3UGP6x/bEiQ3Ib1DxKG/fwsxf/PrafsFx9N8kuzFhGZnRVYjP
5oTdT4/AN6Rh63R7iF0ieihOtMw9KYfDUykOstsxd836Xhqr4ArZpBO9Bamo
SFg0rOkJDsXB75l2ekPCg/nTXtpfiC2Pw8G3zq0/u6grli7GRG1fzph5jCBu
tS2BCHlULcqhflm6ne3nG8NPLQrIkjiWQaQLQhAW3SbTmSlwFhsjjKZXA/ss
ugdBgymfUie3lv8cIVQhyBu+0Wdvr1EgI7qWRg9QotDHliw2b38B18Taxz2c
2ba9mjknpxofjMs9+bZTt+W6zJeLn73FFR9HL856gG01FLBmL5Sxjc0v7HDQ
j6ngemvJrktaY2kwtCpr2NHjaTe/pwQ7EgUELuw18Bdw31Nt0QFWc7Qu3XSj
TudPNq1kN/a1FGkEo1sltTDsTvRwg+aYgYJP2K4Sx1dexgrH+u8R4GZ2lkoa
4uKkjJPfGHkFhCf5xEkUlmVndYqnQV5Be2HZiuREzECn2M1lnXzX0yZI/7zL
LWo/oIYckJOQFZnXvW2RIMebhJF9iRSIQPdBsyYkpNWFO/25NaxbFJ0Poi4I
RdwMA6KcC1QHwGgpXXC/BIcQpSne6/kSm9jJfjnKkKz3oBA4EtRGTRi9XAhz
2hjMU6xRv6sOfyoQSbdPhdR8D38T5JH/NX9MW1g5WbxDZAa+Dfw/1H8kIz51
TiH70BX//2xnRZkWVnI4mVXyYjMTAhSANh8MV8OPt4H+9VPRiRmasiTzZp+B
X/pDH9ssaOWeMhlpjRCMIqJKJR7sCXgsMrmU56y+DmDNVnCI3vUMzm6icqcO
XcJ+bv7nWmTebkTXKSEwaP7lW/vnbz7CTM09P99ia8pAM/ASTIMy2cIUCwBg
zRqF/riq2nqrVOiCkCmEcgm3R1bF/PEQLltBDqZ+hpZuRzND02jp1Uui2Yez
9GANhWGCOCBRucf9s5zZfM9DjIC8sJVDT1QYv1J2wNf90RqPek+lzgDneJWb
6FZqrIUXmpkbis+ZMjCHSSZG/gKpKU+G1nEFRrJ+1dWiEnOLMaPih5mkBiCy
PaiRv3QTlNpCktHH0BWQKtl+FR74hKd+NQOl4Ql5sN63/NQVsDBy8yZUHkkt
ojUuyzRz4aiwJRV7LbDrm5VFJAuMEEx2xZji8unx5DjZnEOKIguEWz8dSnHC
KMPe1BQeHpPeeTkqLo41aQLEM3HQ5pSwsVFQ4AM+ZoOkllk7Cl+6H/coUM9B
lAKLwGO+1lGICPS/nDykkgRgX6pxL/ueSLeg69yW+JvLv8JBCf0uZYiRSTKc
KOvswCzPvnWK2Ehwl5b84AsXXWM5l7B87ueSE4GFRoSRhJMtCTakGYMDTr8t
/ubb0fIDCWgHFWZegqMIywMX1ihWbEvSVIuv/FId8MIQGP5zEBxMnlC8B4Is
9MibBJFsu1lULN7f4MznLteUmRLIcckL1fDWi6D4m6k8Y4d0XciO+8n6Ujdw
nNEkAzTMVCa673megazQVm+R+5mRnGJMAzdOs1qqOBJuvU4DETC90sZ5onsl
YtMJ3w+wu0wyYU60unMjDXnATplxPD7YLHYkvX7KfeB2LVK2vTO4Zrf6DstZ
MFRa8HqRCIxiqi/4jit+9czClD1kDollHnntvlbQdoYVs2iTB+euOwr1gl7Z
TSuvWs95E2CkjnFFrrahPU6y7ShoFnov2oiEmQlU5YX3/56GS39C1lOnhB2R
OYfinLHye+YpKuh6+Zn0ZN+TDz5DxjlyKQXgdqvIE2b5gIOEI+e/MNs5NOg1
LTjUmItVfVfx6J3HWHp1irO6ShHY3JNQK1W3j4G+Lxp2Oj58BdORSQh14KZL
Etsc8q6JbgLFByz3puV2DFl5ZENC3sTxYOluPo23xggvIQmsFvLGh67wyg9Y
5zjkDcDcKrsXsCnibckUsBWBDjfPVbJrpsRzVQBk8f0Q0wVYFfm8SwsHFXEj
QqebhV1r5YarN6nNuh+322z+XtNWK2JaLpomfA7gWllY3WVKPb/w2j2c2t5C
ToBcXv7wL81jTeBJBTMJD1Hfb5iaS+Q9sqbhFNkN1uzCJKJXejbnZyYiJTAw
2YEmMQPLRKF1nNInrM0Xz7EivUIBktocrfHkH2YLCCU0hikAfIFqat2JPRE6
TK+MAnY/QH2+fVDzZysnOg4vQoSu8IvcYAJxgma46Qvqh1+lsu0avb0cfCYe
LUMJ1dPETYBs5+zEv1af8g0EBRjJmEYHxUfWDcIfSJYklqi2B4/k1nVvUAqv
IIJRFNM/dagYfRVDutyc3Hy1mAghI50GRAOZKDzoel1fIzLebqo931+/RHv/
mOWABMSLgIjuBxF0uIVUO7xYOsd06yGfYxD35O8UgvVhVzo4DtW/14nOP0LH
9Yj27tj0Sn8Xrvn8Syme2D/D0fqFwOK6UTvNUIDBvmbNqPMnRGFi3b/GAc+8
AzStFeq0AlGCc3O8MbbvIvq03+/ZlK7SEYTe1y/dy7866Lju8HA4dLqUv1PS
6nC4EaN5trr3bxa7I3hq0TAiza7ivBUmb1m90mAt+DUW337G3n9jLnSuTHlr
ow6yScJPJiYmbqYw3k0Xr4D+su/4Ek3kTZPxn72LQnA/lj/7PAQxLv06L1hX
Q+Sqm0ZNl2lQbCb8Xedok18VvzC4m/PxjTjHvOzx69UDB8b7yYbOpTXTEmgv
3C2sVKTOy0ksuyMNB7MuDHmmQGZ9tpgUsgt18CD4tXJ7k6WyR3RSUPjm90A1
SGBpV5nmFwso9Ewpg1dt6hNTrw/06ib7pV9amk1sqxHL5K9EWVPqkuwg9+bP
ExfmWpk9Q9Z2zjEwDL3bL62cCv9hBVMVnlpZo0RSXmlOw8EYeZFWyKFDoePH
UgVKGmUGRjKfZw6Tcd3xu1l2TbLLn3FCWa9ccD1ohhEhvTJTSJDQzO5o5Rhb
p3s8HRCYD7MSnve9qvUDi3ROvK651DGp+14+msHOSOGDwbw1D8PLSZGwnEpC
EA7a+up+glk3GYKEN8C4PBI8KR37YMFwsKKWdNTWf+4Ci6w5wuCidDlvCnAs
RQlEqe9dkGWTWusfUvbZs1Y4E3yMEicOMfY6z8kDukwbS+1MG2EfY2vryaxM
9lgF4gong9ufNQA03+ET4uPnfBBVXhAtLUtrq7mHnxfbvShJLAG+1e5TFZ16
l+f4qwOwt+Knr98NKxMS2kLN+2bFJeofrySEf8BEXKtQVAYkMCbkpNs5PP8t
Q8l0+at349ehihDtaUyuuM9b+fWnvQ2+jA9/rfS8+4bqZzkvS5PTnNBLEqIp
RyvfSOay/IHYv6gwCAe6zTB1umecauCufEba5EHbdNEc7gQi9AXf9UO6unnE
qHrQ03gnHwZnv4nc7Qmr4uajk1zuoPydSJWxw+Kbn8u7SYbDsjU4XE4LEh3h
PHZSbpF1IDkMW8TbJN4/JEFrld9vjKRNPcQf/jUAtTQBLSN7QRm03bGFVz/s
2KrI8Ix5JjNESWwYY7BI4E4WNURVhN2wPxwL7RmI1bwA9Szi8ND0hWZ6Ar3p
gZdhFEMcKqQS8Gu0towHU7iRkoubrS6tDvFHucZItOy3XQ633MwegTzstuq9
YA9tLCw1AA6tzkceaqNLP6cTC1JJ7WoiYXPBQ1oZ2g1a8NwSJKXe0C1HUn6Y
WOJyYMHDwJLTDOTThM9Cjh+z87s2+wZ/1Qhuv4zR54qnLCEMu0DmXCLFp36n
Z4SROT0eBMnjuiAz+KssTDhAe35J8Ezyy4eeeMIilDZaPTBdY/MIN1lDz3h/
cwoy24IekC0zvTGwWgiOEZF9YvM7ZDz2Nrl423+q9/JHZBh91Pk01twVoTya
nkKWtCDK2C8roSwV4/5CPjybsYjUZW71e4s1FHsi2bQqidY4GLKkM2KwPlGI
LyjnTBIFd2D4/v/o+RcvU2RqeADvQt+w13xAc9PAySjgf9aEu7N0W5v/Y6J+
hIFEgiqftoEg3jigvpzBc16htQ3Gkt8MJwoVKD+YRj7IBJAXXeEFc3P4pItN
hF+xOkWrtJG4GanyT91iR5Dvzv+YZvX+xbHTCI0ia+6tSRZrUV4rMlEnGHVO
HBCGPwt4gxp99KVERj92hPr50Hcu2GWQDOHyuu/jBGyk3c53PuQ3bkhaJS6Y
GAZIjtrgYlt8lbMhGtF7IknQW9qmcjip6rAW9i8T4dGmDWdsah1lOuEAwv+t
Xb1OYdw/nN16fXOgpc9TsiD7fpweysL0k3NISVkrKc/lAN4tZ0Zq0DnzYA1g
9tG/1nzxubk+oeLCYU86Kw89se1Zho8bQhdOk7pvrBo5++/AXvwm6FCtrR8A
FIgg+3+w+73v3Uw5KNA2UQANmNYNGWHssKxYzhwM0XKmwrnbcxvbXmwne/5G
mH1kX5EtoxvTs9YK91xOS8nM0l62w0GqbYS89chhfdiNBGmDJqx9YOEdM8jq
RT8i4bn0kRqEIs86DDhoIQXUzC3mVwQmDKUv7koEtqFjSeJtFc+XHPdXr1r6
j/51Qa4tRIUAPxtYxHCcH5eoH65klBjvQzeVOB5plo6sqfPRxTQZDNv7fBfy
2z++2nTsW+qznp1IImx+bHSyzSrKpbWWRpjaeChiybC80inlsGy9NXVTauGU
j6iCm0N3lZs9MJtUawh9Qz8YakWG6C0v7pwi79VBOZNZLbX9aFwfhpES9BGv
IBaDbSamyrB/1CdoEiVYX6fg4yuYommu3vTtkPjTVE1wNttlq2CutCOeIxdG
Oh2CeNk0iOJwTa+SfgioYHeI2ABNeSwqlVRP8NamD+7qHN5GXbh0lRrfECRX
BdKEfQH5zWo93wTjh4ygcigSnM2GBg/oTN3S+EcSyqdVri+mQq6QfAKRwgZ7
tiirAh+yuo/5ejPDwlFkwsatcheXweL5I55SwC9KnoxQ5/y46Ya/Zu0cov9P
vG+S+vA8svHu7v0HAL9Xd5vYYDm3KsW2We3nkAME25P4hLvsSgjIkDNXUsty
BBmpMg0+Oa8FVhmwSQklLdwbSByfs1XaOrEGnnWpw8m78StzMxZdVQn/eVCb
q/I25gya+MLAgkxWM1VtzRWSNSvC8IuYV2a77ej7x3UmrV0JPNP59bQxMcJ7
3QdFkKIb9zOkuABO/gLr8kD4CYt1fQ8mC7pBtvHm0FnGjSSsd2hj0pLSLHzu
mOyPSx92JTGlxW8rE4sNsmdbzi2Nr+qTerqVFqhiQ7AQF+BRGkTApD6XAcR+
lq5oTl9qGMM3Z28isdPqfBQrhJvX0TDV38inHtTomrccSPdx/iMmID7ptinM
HjPkrWmy86O8iZqwNsM2pDwvH4bAZxFyU7cxms6WSLLKAWFNUfQxOlDXElcE
F5SgZKnfVb1vLkJ+YMDEdpYJ508E2r6nitCTVIQB8hhIk3lbK2cNgmRfM0ZA
+qnAaDC2ysXytXI6B0I1gTtygZbo0ydAvWK6LrYzCbxODhLWJTxJVV494oSv
9Kb+qEdwJOChgfcPvzC+PG7nvo2PyqeyRlCZXsfLcDasdsK6swWHE5eBKZZW
dApcUMaxHyroH03bSgRipcjWU/wS97ODi5KOKVMrUHVPANeU/CFb/uru3FJA
KuevEthYY/n6WoB1JraiUdfUkvYgQRhM7p7ujWg7yDt0g3OGRQwZB5bkYmd8
cjmOyjOdm6/XTpEiXjnaxwD0a08yvLwSVuQr8Z49Ibyo4k1k8ml17PE2PId5
lZAMzQ3lGlm6MuXJK4xsqO2Z4FgssOaekzfQdIxxM6GBtCKOK+LybnIl8UqT
1FdvfjuWooNjBJQ31lSzGuPzPBMh2mfcn+cCI2y3383O/Pwn1a8RtzvqXR4A
dE+dbzQGJAXNiSMwffdx6u6NWeTf0ylBUKqIoYa9ixi9uWAvJ3qQssEbEaXT
CQWgo3q5XU/py7ACrN09BUz0IYeeIAtZhk6NJTyCGv+TK/u5EMk5d4bvskh5
eBhimUs8zxRzQ94F0L3MQVyaiRnZah37W8Ppp5FrB0BEUWbhZwNwJEfkw2FP
n8vvr6JnNTEHOsFwr+W/f9+RAg8cKtY7D18R/rODdWBv67EPE2GezHiQrBYT
Bh7nBWcJCw6T3ERUBo3ivv/UqQymyp6jJvkulGvHzbu1/96kTbEIowsGwYG+
tda6gk6+phUkPl8XgrXcdluY4lpUU1MtmZ3w3+xv2dcL0LeLZ2MgDZcvU1Fy
p9JbDf/jneS8i3rejMtkwltG3oEZzxDxNwSsM6XxrcHpxq3+eg6gH+zvtez5
z78xfYHvzVT3Dd8s4LHtWIlGhrX+fgiBmWvE2W0kVUygT8/cBA55QrlUVgH3
z3XAWW5/rQAQa2x8OVhSwSjh7h/mfWeTlzkZEAVKB26pXVQne3410nfWxwV/
d912jlusW3BxkJFv2VhnSrDYSCmY9e1hT7Lhc7bbh8BbzYYnuJjrUZuAkXHd
Iv35WVn7YtkIVwgmhYcGnUdmswLyrVNcX7uEOmrju6UJOk4tFuwztZl92Y3Q
UjDt2Jo2T9Q16s9v9q8ykSolkyQjkLYsQBxd7zYebbrtuOUDdHNb99HWeGOY
79IFYKxFyBKTEvOwv8271FbmWYGZbvnfuJkMli8Xfumg4LhkOHM89Ee4EsfI
eUiVM+5qUX/RbNCOS/LEIJ3miyWzi6LbIcEq/yhTENcAD5r0rH/t7n2lRnuX
dOCEfwVWPGTBisCTTeCB21a2AJ8NONR3I6KjfiGVDauZGpBELwxEHaL0K54O
rAME03v6fjrek/q4slqTi/oZiCwoqG0N3FP55TBNqYgIZWo0GZpZbSR6itbO
oEzp+0IE1UqX2MUs4ffi+fArHdq+XWpwFQbOSkw2jVr2C8FJlQk2H19im2Td
ptrIJOLyLK/8crC+so2/8LULEyaT/0HlqLmuqWsZunUEp3MqZNuKFHpM1kSI
dNrEReS7eJH33GR963+QEV5hv3QLvGgjyTKLAHj2SHwj7gzfxuXuzDl4NTmW
RJ4aC9TgeNNAk9qyAyurSbKSHWP4Gj6ApkThBq5B0FT+27i5cJ7lc/wBUaBE
FYYe1TGudqk6WvdUcXVR38R0HM5MK6cSoXtLd9miftcn6nbKFycE9wpOGocQ
DqapiLY6sTmH85LKCt08/TWHO/o87ki0n0Y/DhDuWqs4F5dJkpPtlvFM8n/r
L//4P/txIVX34ItwkMQxbAbDtKqr+UKVhGCsNjYJ115xJ0Bg7OQCFjHDTSRR
ncRC0bydB0Qw+PsHT1f4J9VP1n+zx1AGPHvN+eYmzT0Qjdp5wBPFcPg46txi
3u85t2wKP15yex4F4syfN1J2DAuKon2uwS3mFsAUHWdgbQFO4G9/b8dYQ3rk
Kcksyescj8ZbeqG2gJzCIqf9+jhqykCQx4pMwk3r4F+wFxlT/WykPEvAT3+E
o0c9QTmb03dRtURP/utNSLMVaO6c2MIvKpeB8uLZSir+30bJAaFiOcS5Ck6r
l18hLFGb36mA01JoemcQJmLhkkY6yYbTp3biSss/Xrqoz+XcGMCc6Gjci27W
w1LXasKPhNdD22HQEIXw6w0yRMwaLW8J5Wbb+2SQfhCY2rkPdgq435d5vn2j
H54UnucdXpvXSsms/KiJgGKMiDxsnq4Xm2n+/zw38cqYg3f7ubLdjvVzF/hO
xEDg3kE5kq7119jpPTsDS/I8ADpGmuhATPNucAmi7831Zp5c3a3nckFlYlTx
nQ0qxOk2FDlaj07nHVpMELzTKlPDXCAbq7fdCN/P1T3aYAFMAmmEgAyYKX1A
MHkPlwYI4WpLRn0e5Rqd7GFzuyZapFT/QDTjUGdPsdsGh6QOguBNtf8X8o5t
cuhKH4ebPwnr1nDpgA8PoVmLU+syqCesM6KGC7IdDYUuxRzgLZvJD0J7irj7
iJBfl0uR2Ux+ck7qTjW1iGGbySrGFOMpOYWqtF45oHzWe5ecj59WtIKXUfPo
/uhX8R19tmd6txtpKeBZnesGChrwabl+XyhS80fP9B9sBX9mOwblbgQcTsuk
rdccKZh6byiS90jzMioMu824wI84mM9jDiwTH1SKzG+coVs6bdQDhLeU71EA
1y7go1Z+mWdLn5W6xo0+Iamn9lLZtaKgIL1cqJzeo+Iih1OscZ1Fuc94FCv6
2in0+IyH7tavRX1YbRxLkTcj+6aMw6QPWbewGmmi2UsDrQg9EYK9jXyxeun9
zDprLrhHhyXlhTLceEca0aBrtY5LDElJ7Xi6HvEYxWuUaf7wp+uO7j99lW63
BFNrn/gnwhKp8YMrgxs2iKsMsZr7U3WCfdlkxXpwQfrM1eAxgcQ6GrlGwVmA
KzKFn+Kca16iA7x0Iku1Z4pO6992nh3MMxs5ccGwUbwDlQyTIgyYZkv08PkR
XBsdzCk5IHvzNm03+2uK8HF1kaJ67aNcEroaaqN+/UXfXXOX6QWcIvimKabh
WYrKaX4mAUYeLBllvp5DyH2yKsHz3iRbgi4aRQpCJ7D6lVxRAXVjgqBifqoA
iIfXJQSYy8IniuYqwNnZwgKiS26AVWncxUzfmyjdq6zRJkXgsmvzVdjmdXvU
me41EfDfZEmK1T+6uNAxMUTxvoyYF7ASgs3rrgyQqNDX7laJcc42hmXG4EPw
4L8QiHhS+zraqsTVTePXSsmETlOJ2Jr8jtLqfEPCfHs+PzQj1gNFK256Gc3s
11g09c45y/wieqZfLdsrbHdqeSYBHTTnfB0PT+1kjj2jdrRCOCyd5bR/tCIY
brVsCr16O62vSC7PH9OILc99KQ5ajy8ws8l+3+cYz3ZHpsBDdCqlZegiXh1X
Tv6qSLILQ1V6whQeG4Slaqyx5103JLbLZ4JATJ5g4Ql4C0cNq79xYL+VmcSE
MKsLIU19fnPs8sYrzktYNKPmYNhblENqmQymrpcnyAwpIVwmjsqgE+ZXRDeD
M1Vux/f6uQ4uIgWP5wO0/iSmvLWKPdHGD+bNBUohU2KkiYxKjYba5Is1gvNr
7QLaKTRZZRxM8fi6L7sLdnDtvGEFzi6VD/qi8GglAUvJ3Fn0xe5udGt8rCnQ
3N0Fc3QbV4/7FQlTtECYaCiFa97D66b+ZCnlHpv3bkLDW90D7b3GJMduup04
zVA4Dgkcv1e2mKbisFwktciBl08JKSsLLYTNO5J1mgEjSn98XNy/MleOfI+i
m6AzCQqaE2cMFjbFDgSEmfUCPdvzOyV2xsFNPQQYa8SNWWSz8qUDQMX1D810
TMxaYuxp5FQGbDkvR/6Twqy8Ww0O2j9L2Ex57qutkfXo1DwVBntUJNMQWn+k
KoQ1iA/56f6rYo+jUAQbbQq29RMlI9SG5Wua76i8hBixlDsPwIcNcJjadalJ
CdrzHF8U8TJu88I3nrbjLc2JuoFadUJDhdX7rY0aMujX6irRbLBRMxDsN5EP
hRudOzZeXuAX/qho/Q5ey5pMUSyTccb90Mw09+L5U3ggRCr4mxkVN/7jg41C
gVaiR1VUEB8pMOzulTyfOGxnwjFedcvnzq8r0IqeriemLdaWBlfwbgT/xXRp
MgmcC9wsPMgDgsqC1eTrzGjy6FC9NC1WUNWOR1fwXXnzPNjY9tN1TEmiv2g5
w+vDi6jmxC25d3UTJlNeHNG4cp2Z6jc+KHo0uWYbwawwVbyb3A7zEoNQfQyE
m3RXRrcbNN3t8+mxYERMKRm+j8AYEMYXKJu0nM06I8F/pJhaY0NrfZqv4wdQ
RZOwZCkpvNtqVNNtKCG+QakBcmpU7eLUpmHpjh9IRCvgTkkkqB0QUaXXsg63
oKsKosOXlrBgZeXH28mhQ0OUjDCtn6Q+owvXvQPspQHTUeBz+yUgJpCHFV5j
3ctAqK6pjd+XZqmSyFpwQHRQ3LAy/+7i1HpLieJZ7//fuyKa+Nb0Xwi/NpjY
6HoaGsKl6iCQ6nP38Z7xRcnjjUptAaxewQDSRBMH4IXLp87byly7cRHF9Tuf
NsuB93/z3xz7wLtTt5RmZzkV5Ye1d8FRiLMDw4gFgalKmiFgtsgMBB8dre7q
6WZ6VtzBP93M82yB4gX92F5BhUXD/ualccpY4yYUuMr5RWCGR9yTjFx+CN1g
dGyySwIbmXLoo20ycoJhq2ozhn/kM3ydvA+zu70G+le0tg2aY/2vmoItjXRF
HCRBQA9MrPHpFjijn3pZ5mCV3u/q3N5i3Fyo6Jp3LOKM5vuur0rWeNGivkCi
h7ROXlujx/7f0qbcw0rNml3Szojnn6anPAXYET6FRTi+HS7+QEPgIUM/fc3X
9kqUIlgq0Wj5EShjiZmoSGAp5fcuHyRfnnou8lV3lgibkGnkzp/J+mtBrvt7
JKkLjhUPgJlZLjvZ3bL95zXDjWh4QwoA8IzVygzxbgYkFIeyT16DGOyBfFM/
piUH9u1/bWdKoKC40cPbRe2jlprCHIHdcnD3uXDIZbTkvxkAQQ0x/vSLJ7tu
Ij+Ni7R8SeFfwWnwsFae7fFv9ZSw5/EKzf81f4VSbFaSVcFk8ZDiQd2qweFK
S0xy0avqv6oVy6+zb5Dw/UbAG3ulrEwMdsj/a5oTLq2fNqdnVYbUJNHTIBno
oHXjmEflhaPrWGm4vt4b4JTfpV9/w0QcEJcR2MPKcmDOvXzoHFi3c3ct8TQk
H8LcMt9EpW6FvxTo8uFB9ZkengeL3eAwor5V3CKVkQXUe/aUkN6ys49PaouG
81q/03RySuQh6SeqweDoswYmOZxt0gPZrPf6cPld1PB4HFV559FZ0XMvQjtQ
OmVk80Cp1/4xK7DllO/q/vsPJoLN1AtSW4F8QFZuB5YPmq2fsVpxapvaIdp6
5vy5zPLw1I1CWFEIqPSNAq0cOefFhl49J4nluDCNCkwf7VDO42uO6/R3dh3f
5qQjDlGsPZ46HoswgUiN5Ba31jLGYPiN3pJCx4UDEfUhkK8cFQFLe31WqId2
draKAro7hxumMEd5cyGbT3PBmCt60k8N6HiCozmqHdL9ua1r4CXogupXj34D
UDQs73dUJtsyp6HyjbUWkPPFgoiKiqHJH2FLsEgiEukGkHQ7FC1J2e05Qm3q
O/rPxu1FUKRPQQdfLv2VzqdI/UnJHeqULlMtc3sENfGtnSIyXGMG2EjH/n8N
GNZhhu8SsDObak0RbotHrD5nDzkYi78eho3vsGtQxOrH6wJ/HeJKLoVbOuXF
N1yJR3uIgj3nFe608WGn3fcvEmMcjBrs09hktEv0lnE8zoXiIHvvhNcr2wF6
qMxvwwodlKkNkSHEZSQJdFBzgfnbpGEfmKnNR7raHvAUhT72/6rSeF5GV34A
s+Vw4dRSluaDVx2PYcF+POlHVny7NlzVBFwe5ZluO1JxanthOstwHnPN5M0T
Y0QRCmA1uRIUOLllibjYGppAe5GKftVHRWPbIM+srQPrlvv1DQTm0phfnQc+
kj0RZhehh497Uprb+0IXLWdKune8Ee9txaoHWK+BcdoN/HWakUy8bY91yQE4
kQkxGc6sATwUyIXW+X55qlgXPpWTCBVYFDlr2vSNhZyfvfc5qnJk5xsTDHI5
u63HmgQ53+Y0mqQbkMRSiBlZ6E/avzfuoAM9rmKSEzKjj51kywqN4s90skGL
5QeXRLZjzyp9c7sDSz9MhgFAcCEf571TKEc//DFF0AgrCn5ChK4k+fg7Qh1j
X1XXQuETXaR1lWxspxgVxKR//CizPPe3GvTLqmda/6fpC8983mUP//cxKxl8
py3DHqVf9u2nmy4lTT9xVxmQ9EXQ1bPhs0H1MTeSssJV5c9boRWcmAV7bEYr
rwIOX/OVFGIg2NRLK9hAuwcbogUwt6TfkTqPkfxCLeccU9Cz/D82L6kSWxvR
PhGpSHP7kBPbjTBLFV1vOoY/Kk5dB/P9W+xGHBdI0lql41oW+vT7JxqBEvUT
MWuW+03aiKh9AItpcnvWVNs+t3gPvzhaqeTRcwgd1mbexMNWmstIHpFZAZCp
cl/c3weLj+TMtudALDhKEZ6h4Sxlcxvb0uk34Lqw1lbQGwvoXIgi3cd1ekx5
pq8VP9aB78tZO/MNMcyEWo8bazE3Sz2WfoDsfOPYHZWVZR/HfnscWI69FpDF
+fRdN2Z7nL0rkQOp4vXDxjql5gJbT+4NACs+XmLqjCEcOfKuzS9/NDmA2gmy
6jiFGBxz979uJyPRdJSC0J6unruTRrPdWXMAVSdOaenVkWRkRYPdoQD+XqJp
y2Y6A7VQLxj4OYSCFhg75E8WvQMe7RD4xELAg2qLEE/uoLHx9eSexeJJheGI
PQcHA1OPpTlXlzpDoU/D3TmaIsvRCh659pMP0e0iZGo0m5vKfeyPZtoNKDW6
nLC0KpiuDISFMRvjoUBgjYvw08tZQIqaAVMy3DRThp1ZoYRj2c+elw7ZNvSi
GweUJ0NNTNbMCg6nT/K/Cfwz579IGM8gNPRdEIhl0M6X5ZP/MJ9Bdm1o6zpe
6LEcRznihi+SD+v+A7zXPKDWvNIQZz9sOxo/FI3jl5hqkbuf3/4RzUNIxC6l
mj1KW6ezx8RoGkpflDM3QakVQUJEClhkcoyvlyv1iM2vxhkwKBpvfLaTMhGh
s1b83wJDr9Ci6YSGuUuwGTH4YGGOjcHktWY722OXAEl7mkdoSHDYY0yJ9UvO
QLXMvIiulSiANpfyhh2qzWymxJ403NEAX3t0wjJ6F7/2UaG6bGCHqyhX42M3
sMpsU0sBTtU7gFkz6h6zu/NepyorathXBcR+1VH2KZIzF3FVBclgcOtMLoyZ
DefOrgFo/XluNaCdKzSkqyqNrbKRQ6GsPhJiyivQdiQTOK+u//yNMzyELD6b
//T4WV/LEuYmi7DSswn8V25GcQPToxqc5Qih8k71yxCoC2/EP5vKpPZm6OlR
CLU14qajPcbKjNd0OEyaxPCSll8ZyCOmnQgV41HrF6ikBj0NHUCmrunKMpgy
YmudRL4HXRcL7cteclaYWjrGIij22GsJUDZBm6aJfIHdy/srzJ0Ko1QJRjub
hH5xvdZAmyNv1hfovpS1xHMWm6LVq8MJrtPxfgqz0O1vH1zYqSFNfJ426Pr9
HEfW/21Gq7V4vcsLHB5Hv/rdH+QcKFdR1qoPoFT/MAGXMjG6iCes5KcUuH2w
GjqMJwGGX9cXiHmVcdGpVuaBX/lvTKH3DkglN+Xfjm5TFlE62CBn0rFLk+fV
u/f58i2sXIti8LxuWz9rozRn6obvkjAnkXSfgzmyEFaknAXtaVR0jiCx52Gs
uINo9FTlaSlQUKi2QDgppB4a+pYAEZAMhaKaotc7PVHqBN1jNmrBjxGhHEgC
w9hR+qhJEoXwfe1QcL4j7fQiGmb/fK3cAudavJf0W/qMMuD1jqSO86f2Kls8
VuqaU5u9rod2uPY8W47gmZWStTac3o6aSB+KA0UvN6QYV089uXicW2bvFaIX
1W3sVWlXiDX79ybXVYeBZaqpMHYnRZLJeUAPQwcpRJ9Wo0BFg6GfdcAPej7U
xe00Try3dAm1fu1bpwSEP125UqfKXFiTWzAJCBges7JYXfq+hjkypXlwEaF6
Do2P/83ejVVKn92uSUpByQ1jUqCYg9zPORDz758uVsVKYWsucEQrHCtHwsH1
c/oMgdY4+cwspeUMY/+Vjd0hiHPPejrdflfn5QgJIQedYDtdByPHOUHwwF9F
rP2VodqZkPpW5FIcAqzMGh+Dtzo7mPmfDvCBsAcpfaoUDvG6Lz1Eb8Wv5sAD
EMMjDQFK+GJnQccF+Yhs6QVqD9Vo6iUhWBkFqLeYNA3dl5SnPqdWmYIQ9qrp
sxAALlkKmfpxzJcnTrqkUtDwupOkqyEWvrBJ+6XXBFfE9tZ4E1HkXCdJQE9F
+2Y6qOtprpCNpvezENWdx+k1na1DZQsH8QlRXOyRYSMvnNJ8+VPou+oF1haG
sH2OqmAge5kC1Beix1O17CipnyjbulERMajrCLvLgGCMPKI88HWEVtpdkxhD
+UurpdrD1c9CeaTwxo6Cx4VzHriZOeNyyOyP3VBn1a7ASItLKLG+266EweLg
llkB8MDzzmMe50mTDs6ubj6qVfQbZ1q5D8viMVTEG9VBIwUog/Bzp2+CZ3Hv
4jy1z7ADByh3Z+dVxbV1bl92ygtfVO3gm0Flmh9FAly7UiQM2WT4nCgMYsLt
XFyz8YHiQ+4jfUW0UapCpUtAgqx+7FfeOALt5+xivf95Ap7B0ehiZK2O/VXk
Qr4vWsyPrJaBpiY6PM21HE5h6lxMNIOIjHLJmYsZ3XvUkUrEJv+QU4+BQj6L
50B+tA1Ik4aAmqC9gY3XcVBlqpEfIXgFkiw7P0kvth23hK3BwVWRqSfBF1mS
iLhJPGimt8nzUa2L0V4j2XcH17kBA8Ns4DYd1UkEvebdveKmReN4gxJn6LlH
F/xuxBbO/3EkNyllTaCSUB4fk5Adr5lvytbIah4UdH84hZmiCxUyBTyx/pB0
gRYKBWReKQU4GnLPDZXm+RdSXbWhOKIEZnp6SwEXpXRb2+OXcS1xgUE+4Kl/
NYdEhv/yKD/th8ptD9IB8oc1dSQbyJ41L8NpNJM1HgcDdtGSSih2RU4vrcAJ
BQOE3T3ymiLQC00Hi2+WsWPt3vFoJKbe4ekULico7R7fXECIaK2Oeky3M2Th
UE2oN+wEwP+ob8g3aq7R7jvVCW5b6/h20SKzWgRBXvl7b7cGYCIgVXx2UaWa
gyIf70V8ExelstkgLa8R4pThJNby2zl/FjYdwfvjO+Slx/GpTDMAPQnTqtEF
HtMAh19Kqw4Q7RU2orE44WY76maShilgDAi2ULCreSayiUK90WNa+Ah1NQdD
9ttasQESNjC2PWHGWA7QwX10X2vp4iMhX69zAtRuwYY5NTxzG9l9zl+woPJX
DmHqTdzrmpttg1eg+21BP7yfMdQiTM+1IAHgNpzQr6BKph+INDojLyHKbWpT
BOzhQVGYErkVhyRprug/lguwYNSHLZ/BG313A2M/TNoCdupva2PDdbIZMqj/
8FciEa4y0HKvqqNLTLFD/u92hzI6FIWIwuS9X5u0+gXFO8hlfz/R05/cAJ9/
JWJxcVhxOAJLzNQW+jP7AO6pRBVfeGVu3HyDXEzWZVtKaG0LK9PyAYnEMxjk
dBPHSomJSsf68c0zut4RrpC/Jr3KweUZUJNLORnc8/lV5Hre73+4Hy5iP2EH
Wqps95nOA2dyzNqZk39tsY/W9bIxh0WLL9qjzemWC+8wGWrkHN/3GRZ/ZMCs
tOkxVukuXVGNE3N4LyI5im/amC8ZcDGUnWbuezPZZ+R3PRVvDZKLqOA0nd5a
qIL42hmmvCIGGBKYdsJ7aRMxk9d7FGY0DF8JV5bwcDPFxg0kLASw3JNX3zNm
YXBhbEtXAGwQh3+0PfXZz+kyCLHM6PJvW8zkv8U80uLTFW7nNOb0+Cv49pMj
6GF3lHjx1qSzXAqYBPPG5+xsWbMKYOkpc4sL2MWDy5G+8dC+1wk4MUQ8Zp1r
50+41+KBUmDKc8qYEIpftQ9iKzjjXGrTjyk0/z3f7SRwCMBiAD+ngxvbriEn
MDRks/aoUUwVQj7IEhe9zyvNjDyjJ4xZ1s2EGgqkyLoASrthyNCFsCBV8QTX
BuU0v5ybaGwUIcYoMh4UuthfOwuW4lIRRM8pvsmuXGduCTyH7KsFg2HAj35M
guFm+oP9L4tqwePQshxxQQqzirdeVNN3oMWQQqwK7hnOZaILVAmPiS/Er1bJ
4x2+Pt4YDEuI+ruqe+fadQZO3bFjDcnFzWLJiKhk6JYu/4aobqmiJjDDgZhC
9QtNr2VRX4VYvH6R+SxhQd3JdwFIcCPyCqn+fXzZmqM7kaTHJJlquMjHzUwA
TTBzfKnQ81idVup+D5kGtX6GeFxebN5CImceHAYxXPn0lpUQXAybmZS7RRaR
EoMSh1v8nNxKyVw/ixnEg6kuhtfKgmD4Smfifm99uaNGn+wYmL84Mlk94fQ8
sAh+ugG3cLuBChH2z8auBhgDJv+mQFNiqmR3IMHP+T1Vlq5D6ePAcZiLjRzX
6yglZB16TCoBwLX7/lKEk363mLbPSsug+BwzuDGzspB2s43suk/pDbqp6Uxf
MVxvJTeAp3EKqOzAg9eL9uSm8YgOA9z8ovmJWPeuHYOuWRuotQ/zyKKK8W63
2tXdJe4uAPK4G964gA/DEt2/BPUFU3c1vATopMhlYXkNLgA1Fy6RMXhOSzhs
KfitxPE5Htu+mFvtYMqOPeOqmflNGcewtSiiUpkQVHz0dq/uZXWs+D6DmbAu
mp9LMtqUngYrGay8W4OVc/H57pQhBRKho8rJPd+XAT0f65WNIqjvgV/lXb10
8EIjLNxXFUwa7USTmjgL7zTzkxyx6AFd8joQNo/jtywFA0w7sFtkIfT/AiZV
V9vhdhqSofkAg7oC9Wqiiiqw04Lq/4fu3ZZSIGshOJ7UssWROwjnOh1aOGEB
L4XSnoVxm4gzxer8auS3ubnEVAek96/XX7K30TgqKUr3POzw0dPy6r9XFKUD
SkqiOOwS37RZ1wWV0Fg9kW2EcLK58Ic22lAVEqDbuzPTx8amBeBE3sPFhphB
Ezkg1HyWSI1Dqqb8m5kKKO1Clz6ewW7o6RlaElPD+x3x7x/qYPff0+d99aoU
AeskFP/28kiwguvtyBpdfbRRB+s0PRqamOEly6/pEp2KXM5fzEFAscV8FFaG
bh3hoNiTFtotdGlQi6NOHDUg71qOlvg8FAhYyh/mBB7Q9I6/2sKJgy6oeWjA
ZlRo//tbaGNNb6On8Xeb08HnvIuIlxyPLfkrQotUHXngfNx9wFtRXnfm1enV
HXSLkUU4VAuU38XX7KsNT8b9OGw8ppCknS+34yLAmeruxZf2RC+nOclSBU9j
mPwWDzBYyPB4bF8UxcgVjJhNpj6MXxIxGmrfQpEpYerNfhlLX9WNre6et5+7
0Q/z5eNNVcOViqXMZeT6lnJtigao5NSzD84ziDtZ3MGKoDiXgUB9eLiTIWE2
iHa7iYrm5s6fXjj89IOf3v4UrzT3Bk4vjd1oeXEUN/CzKKef0o46ARKJR8gV
TGoySbbZ24duJ43F0o6QyIAaViD0bFBIJBXdyDgs4o9iB+9GDTDa95QdmoaF
MjxMImmM3mwUJ4doX9XewT2tuoNoNU/aAQLP4hEgd51viNcc2QUAed5QlPGk
VbBCItJLFI3E2ptQYWSFioVVB/wVwqCW0nxVxCRSlTX4lcjdozRNGI6AjF8M
IEqiRISL4btSJNwSMuvZ2dz/kUknp348JMvQHzXJiIzqYZ1UudGQiuCIw2D9
ZG08B5hNotIqX9XiAQKnvzbBK82/L06jVqyUbw7EwNSbvcRH4+r3bJvKNma/
/fKIRVeuB1TpbzrkkJrCAqI2DNe3J3a78axbg04uXDfkmvl03BShXqFRtsRT
CbLsRze50f2l6ozSKoX+mMOrMZilMPoOybQlXcDK9G80CNOZnNjOZr5HYy7N
dH16ktUFLCfm3ipynJAS1pj3uo8HVAcqyqv5ED2jjSBYkSBev+M33Mm4/8IS
9362E3EHiphq2QLRk8/BQcQ1WHnEc3NJKuLyjUfhMKqEdfvwdYK8O3ov26/r
ny6EFWtS90er+fkJ7y+K2ieMYmlfdkQIwYZxMhYxzR1OKw2j4tHw/TEKktho
3iZHyiQc/hAhFxTYewSr2MSP7h009qGZGfTHyvbRbvpmbM28XsLWDF13ovyk
cwpnLGOdhQ/Zoc1zdrs563NynmMaI+lQA8oRtwuteXNUGzGwARAarsHsMwnE
iTPomUmGttmoQ5o01TPCaXRO2c+mxKVcPdpY8VSHc0QK3R9C9+3zBSuWJQ0V
hpmvviyWu4yM3MsqxHZ011/IpXTVYyqNk/QUriYBQJnAc/KoY5g+ZkIZwfe8
u7Ob0kmFmbHNFRhNdnX6tv8hDUSrIoEhObMdNivLQnGLeaoD9uxSiDqWbuBt
QhGuhOxeVc2pBFoOQ5bl0RzQequyKo6iDqyb1ib7fxNH1OTf7eKZxb3L19DI
j7MOd1PqHJf9RwX8qbMXRs+O9IX26GnycYsMlBF7v2ig+/DlZxuPfwxUpPXP
KWVg7zxum43+8SBMavFWEelatDZHZ4Arwm4QKit0nubFziCZ55bsq806RGqz
nMMsb/DSgQnHJmU7k1/l+/XAquXv15re+3vOjqS6WYdKu7YgdwRrfl5a643u
cpHLGPHdAqRAB0waGRXdzwn6flVJe4TkEyjAqP+V1H8N/qbIqK/YG3bvEiR5
xS4VjjGEkL6uV9kkUiyBQHhHg5DQDULIMkgZCl6EcLEtbWsLiCbWkj3PG97r
/MrNl6RCKaBUFVOkz88pOIkwW5Gc8pYBH/EDvnq3Hw4CXmjAfl1SSXvWEbAW
nDYNAwJnpg+RgD/OjxrDtj302sJnpPi/FDPgyno5DtYkmaBX4JbX/JSZAkoP
wuuPxXEDAJr5pYhgjZ1KGyNW4RlYZQUk59/z19fDZIFALfYuH884lr3zuN21
WB8LYFsRdlNwm15VTfmyb3+367UtLHK3uaMmvDmhmA+3YDtV2RHxUSRgsr25
H/+FsvVUPWRDHwGEpPF2kHnr9/0Hcp9lT7wzqXaTV3aTQhdASzXXHpF8iJYx
zE0qmJ8GPdVgVF6263KhzYqL0kC2ndHKwuF++4jQOk/Xg5kdysRekm7BU25U
ec7kG6b2nktr7OwpuO93u1uFpgljMb3cUJ785swRFuF7oGWAYnd1Kc+lNf+f
UKn3WBQ72oLbafEm34HAUb7NQOSJGVhUzyLgnnOt9uyzStaQ2mVAjed4dgbn
2XWse0TjmYBuq2VoUHS2sSxgvSFUPSTDcNogZNB4kGkbTbNEbxIi75xlsIU/
7hy3VuO9/thdPKDfEy6hf1kGG8hdv8hC/RH4+8l62DOf1ypo3Psof+RYITU6
CjedCcwaCYfFV1Nslj135J6pLDyJ763Sdfmcdy9t0z1fvWKdN1e6JelbcbTb
tO1ou/41UaM2s1A4fvwUstPuL1cJdNaiWMQUjKKBXrT3CaHtp61Egu6Qg18U
wVs12hmY5zp/dwqRVOe0vJTAsAst75Hl6TzWpSHt1Xyn5XJv8i+hWOpMM/TE
V4YNkd+OZ/gCIak255AwQ8xno/VoiGt0D/5X31GKN4OAk7yf6U94ehBakRqJ
BZD/SwI1dDk7HFJ4JHdLnFa6ZccFwG3srLsrXehj6/3lSO8P6n6CDN5wVgcX
+a2jssEBEhamWwiCn7X/9dRmfecdw2yIeT89X94risNqkj1LD+Wg/traKpBY
BbfYuRgrn4HGyFsCop0J4aiXws3D/Oc2eVlTVx0Dt+u2dKLmDO5zBzLdNolb
jN64NVhMoGiHODAkqbVoOvEdqNRmSRlvvfj9mnnSnBnQ9HOH/7rHdKEmSvxN
h43gpBb/nSlWKWzIhZhTfpksKC2X0CTI5MM2oQpAZsYy9j57TJaXNHzcBpwM
dAWGMH7OqJnmkTKY6vks/DBQ4qXf9rhS08HYS+vIom+Il6kpVCWsyTBAPr+R
DmHaT+QWZ0jMHeCJ9UHYgMpPNQTJ6hOrZsXB0e3XuNXEU6MZD7z64vET6tHb
zCnK/0GUO5ykMLxWVtY1wk2wk/JUetTtTd6Ff06IlYdO8+e70Hg+0HQ23x7P
HyklZzZFRvxBbPPXVMBsI82XcV6/sjOwFzTY1tCcc/KRePTKhT3SGGLdC1MD
lV/fbGoPplIav+b+TMsFVXTPhTp8yoThcZSuZlp/mG9np+WTf3mP55xF/AAK
ItWsdKXjKjZsQCB4C7gfBDF7l+2ysYhBHppeVgGvvJirEsDOdl+d/2hYFZZA
5O6LNqpTiIis8TD6/Hvx63RC9eoRTaZfX0am4XcOx2rppzMWiIWM1/TlDYQq
RAms+G6SDzmNEwkMorxF+TytNrHduItO7BLSeT3fIOQL6Gtl8ThMIk+SOHFL
d3nnGcptyodlSSF82zKncbRiFtt6dp1AN+9jKkFD2vqHKDjq4XEXAonGb7et
4FiHSjHtHLSc6w1wVdZe6KPl9JTRPwqZMIU7MJmMrEyLATZIiC2Zn/87Wn+E
0I+b9QsxpwHfNAzy9zQPSI1pl28N7m5OyzAIbUh0fr+4PFiAfsShIxW6einT
2JbVmmQKRogO3NY1eDLbvqo2WKO0GFUK2GI7LlfaQVwdsH+0NDzI+NxAk9G/
NCQHuXNRHHGIICe7F1PL//ikgXr1kIgLjVLQcRpPTkSuSyW8YrUaLWQwPQKL
aycXadyAg87Qd83jhC5mm5jHan0nLs3FYp8QDpGTULY8bZLWzxAoR1zvWvt2
FE3uMEAyX3IBy+46P4HsLgMA1lFet5TXJvBMVxaHTFINm3XwlO+5YpY3/yeN
kMbV6OUBZjFeVt02VUX1Kbt1HSkavCTk7f9j7KYc+Vo5XquTxlp+47LnfnDa
o7vkttrKYKJOh57+zgg1s7Zb3v8x1Bd7VuIqTHXfCwE/q5kTMBFVD2a7YAaD
bQrUXkmiqqBsq8WURPW7ODQfhh2+IJ3HhrIHXwqvtHbFpn8ujwqxaI/ztKrm
93ATptIjnOLXBu46E6oYlrSo+vnyzZh4ymak0HLkCeyt/DBXvmLelsv7aMoB
Ua66xvQM11rkY9ExQOplQwm6S/auwKZRwElIQMPJ4bA/S4W7IqmTCrHlBvQh
4K5nkPx7nGY2eXVN5Jn/TzCxT+kdI8t7uUGmS3isezUaA7nDJuht3typvHKD
ATUzGBJu/G9XTtC2usEm5uEpKENuEwcYIUXW0YpY9juiNwAf9axeDAU45kuS
piUE5PL5qa/ZQ6QeSMzBytLrAUfaSFO8MfjtIV1J9h5znfmebmrGgrttAe7g
AVWq2Hdo7xSJk2sr+rvC1/kT2wz9MuM3sw2p+3ALH5OyqwqxsbzMkEUWfInt
quFnbMiTnriT9k2HEzHWLgmyr9yn5EmtB/DkJ6GO11e/fVO0n/Bio9CGm+9e
ANXqQtmF60kcLVnWw4VvTZOuQ4U/vjBtjGEji6/WrRqoiwk0xDhOaqAtKvvD
1tPvKeIKJxqyw332JjOI2yx3mlghU30zTSlb7xH1AtCtPYZC2vbyl+UWH2FE
nQCmYJT6Yf2FpLJk9RdUcoX1T8j0KyerZ2qbkZkxNauY7RNJdze6vs7Lcb2Z
0+DQIQ35K684UzamJrFmtdiJzs4rbKooiH/OVKz7i4WZXIMabInO/uC1JcuE
Ix4F0f83wVDcRDwm0ZNGGE5EgfK9LO7hwr0+GzqqJkM98y+NdclvdQ9byOfH
98pTZfr6wPE3RzLT38aCogJb4mQ27P394l3kGGqPnPU6pfhF6UOL9zLStMQM
4g9DUgSx5CQUo4y+iUcncsk+8Y8+rFHwoqkKVFDBvUYqedVB+Aaa12UBv5q7
B0yIaCzjkOJHeKrI67h5Lg8rqLJDzLTzD05VekkmYVFgWzUD9dVhbYtrwMNk
mw7oRJcyTE7wK1iS4PzNOVUPhsNgU1fkr98nKYzgRVnljOOnbRZu3EXe1nXA
duiD3cq3+11igPx4eEGbh/hTgamW24vTpQDCkqHFFD5+9YmjRfwq9QlvJz1Z
IUeC3bhZCKPr6amqEH1qKka6aPtObgvNR31BN1axhuNBY95imY3CzzuRvlZY
4fI/OWQCaKVJ6HkKiYpUxHw/ueQHvrN4zmb9HDJrQQtW+bEz+XX9sm8LFHEq
bxmCn9RYSst2iTWSph9IjR7fuS6SN6qztdxSHq3B3cdhTkuNhk7LSz7tijK0
vBRf6RewF3ZUbcXH4T4SGTWWJ7lnFmO+BLp5ODPufqEsbN2UjSWHYpYEZCso
WhvjzoWPPHWqwEHIr72ZT5uhEddlyOxxrEHPZaCMiUa7e3+D0zCVZ4xVhy7E
qkOKPtocpau0u2MUciinhH67cZ8/blZyxoRq277+T06dByJDx4G/EzQNABN2
/RpdW8PG2Tw/Ot9YTVIfCHBnHWU2mU585tm0s3JmN3sdWwCpeC0iY9N0UczZ
RgFOtrAN0h9MCMiTkPpjXgQyi5MKdXk0LcCYDNP3sckBp+qgsNet7w/RJMRj
/rMEcqr3lmfzt95cN91f0FdbcOjOfZzCFJvk2s3iNVx4EjpxENCLzowv6CZ0
lkJDmCYa7WokFRSOB2Me7mB8r8htsBv/nwBoNbL4lETbYiml6yV44SE+9kr9
XZL3Sipad6XPSb8UR/rC5M/0sFBY5lHCKH5eD63KVulqXweF4A5i8VA0yJeq
PFpVeeOq8qF9Oh9nMVWNd0qWENfE8FjyCCBoXK0TbpmUW4wiUQMkoTC6nqxt
f05ASfo6Jx0FEFn7Lg+48VGN0WaHY6iyxoZHtASsMFqKb1Cm/lInUYeqiUcZ
eL3bzzVJOUD1PlMF0T4B/GVKpuj0+2LSoNeTqwg3sYiN61zHZBynIvpWJoVP
wI/LZu4eRNcuHYqiQ1gpYltzf9HJM6nxCtiX7XHq1iTNl8OUrZ7i2IGfrISo
F7FujENyC90L0DbD6/NlAWw+kLb+FPe7MqHIWXethju04vAF1gY2XXi8uzaN
3EO2tlLvuNgkZR7sru+QMQq9gB6ijtPQIrCBsp+qFhD26B391X2KdNqcJpqa
5LT1xSpzmTro5p3ifptiauLt/gwvt32rweJBOw2pXfTCevrGjkCATj9KUPkw
vUwrUuqMzp617mdXvvOW5wpxFu0HSGdjBIeJ4Lff7jtj9fAw3pR7Te1bCkvC
zu6HWiAaTPZIMTk20MUduW6xgkk+Pz5goPPvOjnvin/7Kx5NQ6aupG9vP+jm
xtHVg/TFOBtDqpa4Farjky/DcJZsU9b5DjVrf4LsIReoBlpb3VPoUGDcRdi8
31Ae+Twt4aLKk2SmHrIytjhhg3W0f38Vs+VOt910YX+xaiAMHTtbIvcr7Ee3
vvlcp0kowdMYo6qPDzGFGwplhmM76/5JJHY0pR+Ff+vkKnBk0xQuB/6C44v1
2iizvj8rLXnvlNBSiYMRmXXQOnFGxShpwsJRH+7lK8OrppRATg6nPLtR02zx
pz/7KtmioQadVaL4w2tWAsvDp30mqqTLfrfdrR0EiyuN2nAwnqk1Bwh1Oj08
nvO8Yfmg8B3brhLKJXQN3I0J9l5SLGceVEL1pYOqYYKu3ql1mAlnnrKsMW+c
IU68CkqWaFOn0JqVxUH9AKGsmW5/qKOWus65yCaVi3ykzsTX7sbQ9O+m9SA4
sXOH4Z4ViTvAKiHr841s5WN3HWfsTTOhwCVnL1EN8c72LKub2mKr4ESPEdCe
Y91RskmbZxfIzGEfPmD8hMTl+PWL7Vlbn2q/n2gTP+JWXixRQDXoCJcbg44G
rXEKcGBo76jqlUF78WYQZtp/QSr1RNVOqWedDhiQ8lsfF+vGJhS6x9BnW1nl
lAjxLZ2DbkzNQ0YIFWdnBImil4lLuseMi4lx+wd32CMRIOgDLcBCapiLURc6
lxOvRhVBbGrAN/wiZXbBIzkdikM1NOU6sCxyPu0VTpBiafuRpt+nkDJL56wJ
LRDa7aegLWE/4DPj4AbfBZn1dZwrTsFnHaMQJ6NILuKBBowOlet4dJAK2Uzk
pZEo09fdg3EQ5zj5e0Eb7LcP7iTZlWmO2cdIeZVo7iMUZ4y50sBzeeD4aYn6
RKdgHvB9Tm+3DgXWHes3qmLp8gQjzjgUCLDq6cHhsOm+i9kppvMxuV4hdJLG
BDRqWdPG0+tfoYsg3irp0AHBy4aeJbJNJGlgdf8MM+mTjnQxFFhSPAhyOrIM
R9/d1Rar0JJSHTcw0aN90z9sC8/2Wzw7itHRLki0IwZkDt1g/Hpz9SZxaUI6
zaM1HzbB4lb0/dJmX2A8Juoqix+RF6srD1jowulUcAcG+P6N+m4PMiDSfZSd
8KjQXlN2Akg3RXQ3Xn4bWSMmdt69xEwOlk0VXYqGZuk1mxK8eOVETLoX9ITD
yVgnCOsKhDMrIpmIL9fNyuFBoGHmo62S0bdU6LBKYVHqaWT0VW8eomKcfg6j
G+E78T98cgGEfZTuPIQ1Co2mFmb0MRmxahWshMx4TwdF/SBRzR0PXjgouved
gV8nf/t9baGugDurqXvXydQhZq+z4YR7uXLnvTqhCF6DdSGFmqt8vmhoFglk
/TmtHzJlwTxYaTywO5OVvg0J1SzqVln4FivYAB6idRLcFNsD8t6IUErbTeWa
YWiST2gT2EJQHh84gCITTvIdFzZTvfKlmJ4cXp9kYOIQwfarZ+DiaeDwsxaI
b5lhkyyPKEz0vGd7Q+/9Ij1mwp4B0DaLMhjLqWGSRMzz8aiFAuoS1ABq3yAl
BNjPSl6dnn3UvIxvVBtld7BtqCO5FIT/ig7BWxu6ZjUAENtRcFH1d41MKyA8
e0jIqSk5pg/sFTxytuOVv4A7JGaFPS9mWxkzYjKHCUW4QfmmnMvHurqR1MGD
X9UDba6nTM/8XGVX9C2KV/LsD0R9xSeXsvwqLTtWkQXJe47NuVTfgz8UVrlY
ZeA8/1yox/knZpJBTA5v62VlhTols6Dkc7Q5CQI7CZhMhGZ28Fbq/qjrsR35
TfEsoyON6v2dRXjMSHE+TfauNNrZBfRQahseTSLlmGFSmMFIeeBN17QsI0q6
A1LPuLk416SdEzAVSd7f0GXdeT6Lm/v65V+qO18JeekYYi26gb0HIHy2GsWX
d0DmApcI8GBnlJmlezFki9LV2QGeAKwnYL1IDAJbODsvmyMq6JxOg5jDdDzn
BJOKgUIDHP19YjhLlmB3BZrjneOHwaiLcPrTQWphBjLiayrpzfuv1Q8AmaWe
gI17mtbKG92HphD2rIcEZcRKfAOc2dhU4vh/iP7eSkTKYZqzwZdLVCwiR8lD
MJG3EFX+UAfXwP/15EcdVpt7u59WszopTecuMFyg+5z6oifH6ZlGbYZxiFqS
GJYXpuTubfqyrfTP+WG36o99itlb7C29X1r9wV/gnK+ezj+zF8LsVm8BvbVw
BlazCbym8nkOYCfAH7keJ9U/cZR2pJI8B03GlmCPo9jmNLTQ2qPdDfEqiOT6
QkUqWrGqqmCASH6du5qoR1vv4Njk3a/SIM234wT5F8yCp1749nPYmFzR6vdr
WB/IGIGhiYYWNa6vI8eng325gWDTkMorFArkQ5HaKDojM20SwW0f9CFb+clX
aGPP/xMmoSmYZY+5NK0S2m6M93gaPvaqvWA3UIuHEASS5gfyCXvdjAgQ/hhp
tYuaBANDLWjekwZ0xJUPGquZ7+HZsJrOZ9gZ9YHc+tMFqksZlxqYLRUksCjR
RiwEjczbHIUmh3qg95F4XHcpRWXJOCfgiuBHLNx459GuKpjD/3QW9KCkZnmy
TCPZwyIpZNR46J9jNsE+al+9Tx1R+EUObVNLicS//fMMsB/KmWw4MEyjhoRM
azyCHBeiE+cGwUuMuJI5N5k42HDKZyjqG37DGEKCWKa3aaxFP5/yn9QN5s3e
NgxzUg8BeAWUZuIu6JOvdfSKr+OvB18aXUTbONmDzQWcDskDRZpp0GsjVLaM
ppzFpRsxltYnnhRuNumO3IMFFdRPiwosh3HrrnWGFq5jNY0csLPhRy6IhWTa
Zd+srLMQWBrdYMEkJMAAbF+EMFR5gtG01kTWhPewYL5rvTuqiJabNEBYHEyY
FZDiEgOpmeZqnWPcZpsHDg7s5qR3Z+H74UV9qj1lozfARbJahmD3YsOiou2l
deL/zOy/ytLlfB9bLYsTD61GJXVmonlCUd3Fcgk2JDsypaXdI2a8tJJsr7il
fLIG22dPpK1mznNSYIK3SjY50QKNhcQ71LjKa7ju/OuiUDNKYdYN19U3zupI
cT10pMS+cF8ILTcNXrfMdkxpiYC6u9B1atJMyt2486oPL5dJuZCNQz3o1XIZ
hh4/qSQsb92pq9GJvQLFWkEtXEni/O8IFXIOWPwFThoNf3nz18zQAdWIze/p
hlXz0Mw2zttLVzumpbRFq17ICxrAogbnmtEQB88sdpZLqBF9Ytma8vhOrJ0B
9N9BhXgvbKgyQytg/QrR3jjrBiVNphSIYMnWPy4UD3B5/gSoV4IWCc3k3WjF
P7EhP8LgRgSnFrPit1c5L0m6bINgNwr0bKivmj1K0YthRmpwIv0lP6wSwFpZ
tx4QcEWptmo7hEl5t257IdcrAddX2ThAk6HrFN3HEwkBlerc1+Wr711R7K/r
HzxFoCeASpxCu/GYO8GAWhDLhEAjCU1XCeC35s4v/Az9ymGlrZUQ81cik/5m
AGzRNvmiRJqUfW4hTHo7I61iAP5Fe3lE0bWaV9SIG1VowCXH64BCQ0qvo/YH
+lUBD5UBA3dTLdG7wB+W+Hn+i206qranP6o3xZX7K0XFRWhcByJWpt5gYgtn
vqXzb+LwNGIv0bWOwH8B61IF+ONj1vMsOEDy0vVmrWEWV4bSZkDKbzHkVlVZ
pqHd0z5T638wo2DOIhAe7NNQbtTWVBonttAEKuGb34aJpVdEQmjkKMVf6ZAQ
AWGV8wJyJX0VK+dE/l5LBCXD6zBFWD7ZaJCnrUGNbqj8Y13Mhec/INShNdMQ
4LahP19FZfXBprff2yjzMHpH3yt5q5EYN6A26V9gqMCtj0//s0gIUJ6qTE32
eOPHZ90k4FS6vpYp2XN82PvH+ZjUyzJqlSu5yJxv0OIAnFpXhMz/eEXTjsYX
XEG1Nc9rD/K/qHWznsetKx6D/6uc2seIB8oiOzs674bU83T+0Kbsn0gvRPJM
DLmrOhQhausetDJ2oAxULtOWorbPDpWEX2pTYKKunNzHNqtUIqQcq1y6xk6l
j4xje7MFdGv4cVQGuGPIvwdtf6ITJvi1etovfvUXl54/zeBWucu9hzbBVPQn
fAsdWm5uEdZIwcBHHBxeUmVx66I+uylSCgMQg/B+Zb1q2ymXe+ZgAyORkRBF
gM+RYsUjjIrnVpSD2YLz71x2ePxaXm7sGxd8ctaEqyxh1MwZTwvPkkr2gwY3
fq94XdCC5wGEVvVONMbJovRCa9qEXpEtV3N14MzQiVf78NjnP6hlY506/p+o
Kw/9P4+R31D8i6LqmPr+jeWpVlEbL+Q6xADPdEw3E86dLQFJQ347usBnklOz
ZoVRDeTsdul8Z/S06zevwUWvq+otx0FwvMi8mWlTzC+Ub1RudL2t+t/Lr4Ga
r5ak3d4kz0a9R0/S4Py7DdUi25xEZuAnId3hBASk96DQWJjujN+04H6hcuHv
VzigAeLXNO/TjWrW4PiKG63fcEcIN1HhSwTCWfjMEKMH7p1KqHW+rtw/9IvM
AZvzya3r5ieMUc/abduF+DR7FKWROHvWDVdOotXPKamC/NgPCDqu8RGEsJ1p
njHldVh3RSd7F2UFUgO8bXl2vtLTkrNy0cr3ViaUql5GG12u6MsRSeo/8S+v
kyBadDo/j5Hd/yukUaNoFT0GeNtohAtEjh9HnyP/RUKUHzR6pjdPv9xQPEAA
LtifrebR+vnJQrYf9dpP7cAyUDGAKEc+U64Vi+E9BzeZ4KYNFb10cQhQuacF
hEvRvXMsOsKSjj1oAqYz0x67jMlwwew3+Y3SdNLHj/kmGPDmPTCtG3K5/xsZ
6zy3Ov0BCDKbR7cDMYb8lfMihqmKgRq0bvDSunfpVzhLXvLdO2D6hRqs7tdv
0bb8N331FZP/bcRzTroU6SxtHC7z5kqFzmOJsFFWbzjBV2t0JBuSA8ycTrCt
LWiC9HGjqmds+NFdVV7oX5tiAYQsadQ3eoFtNqWnOkDsysZfYhTsBf/Zw2I4
hPqj75uTtU7UPQskeCDSgLW+hQ4GrjvQKRVM3kP4BJXjpr6yfqUEJnSmUC0Z
3LABBhltBjlsY4Jy9Ri05UsEmHRuw0J+0XAsKyX8P2wnuESIc1to79UjzHC/
ydVLhcuq4ZXWmmQnhjYHh6yNNReTNeAdzd4oWtJGOU2VxdvI6dnmQhiqK0js
cDzM6a4Wk188Aq671h4K3ouZhvlvGW8Z1+OQBceL/US9gcPEyKbRP8HOhgId
iJbzgrMV4K/jqmqh8I5vCtwb+GBtq8dNgWUjY+YpmVCQu4ny/XJtXH4hjFyE
ds0cUqzMK3B3LcqvHaQgTo9K3JtO/dQhI+tS6QDArrdziVZDNMqjZJxwLEJO
n5FzVxnQNNEHFGDa6P5+7IbYE7avHwyouK8sqgd6INPin40WKV/a2lPX59oq
+4fplk4HNmxWM2CFpb2Ebepe6UvklZ6LS5nwSHSyyIdgD3NF2RndKrLYEwdB
3AVhl5JsRRQRNurN/BEpR2zBToKjSnYLI4duU+EaA4L+xzlUcamMFLtYN223
DPK9tNB8xQOdRe383FrlkcjT370Aj8R5aLCloIYmV2qjCDeBVqHwpIPyfBWV
VyQiVkwS5+gxNx9Rgrm00lA++VHMAAEzLsbXeZ4A0XiKoRzlh8c1erkTIPTj
LsPnYpbQupiGpEN4iyyT/E5ez4yNuQdvk8qYsw7tgmUOL4GKmromPcgJkGzw
i2f3eHUlqQFbFjZj0KlZgwkrY/vcxrEJS1nVuzOZLHlCGv6yQCIM16p0d4QP
HvJEe6PVT9l8Ti463dossXxLcBE/KsIKEqInhza7UxlSW7aFOw+h0YxvSWOq
ehU3qJ4B7wAPjG+XK2ag14eQLabzTVydvIpb0G7TvTVEpT1ueMKJH9GxDIB8
xNV6XJFLXS85wmfIsRax7fBkd5pQTexyUBktCUMMWmwlCdNeCvxs959a/PoW
19VBK+B3Pywpo5JtsWfrTktfoFjJalCqUxArMhdWzBz2GY6EX4UM7X0VR8xm
j8LIBCsrwX+56V3MjBRENCkExtOo0ZvtXE+5nPv0EmrXqNmUUjZ2NKlpOSTu
pU9CgCFtm3uP0KMJLapc7azLo6BrQo61SYAQUKSWE4GlfaXhAokZMu8ZcpGA
CM9fSMqsbSByrzyC39Hb1ek4hSvnAF/zxiPxS0HMqd//a4c7Emn2s/CwrQCB
9vFtiLxTwilaq7DkEkATi9j/PDmxp2SUEjIUwVoltfsypFM0BL1q3VK0mcPe
LSe8E9p1TCMMdClWDNoXYbsvtCeXNlNO8D0tiRYAvtCOwtkmJOxluVncGO9w
8ae9VQ//bZUnsRGFuWlznJ+aXQq1IEF6C94VxD15bqpgtrNC9gmlRXfVrZNs
pBRd/g4jfKsb2ifgL58wPAQvk+4yOGNZfPmgLYX6758vjpSgMznb+xz2eEjD
tgbsaqGHccFYDl4T8KZyYk9kPPvRe+JRf19dXbKdsQ92xjRnOxTabtX3TZSo
yoqAoB6TfPxR14REKFLyMiKPEUv7/2hU+Zm9UzJy31PQ8ceaedtlKR8R1HZ4
S56LiHSM0iIxqIdoEjTc9WoGD6GMkkSFUm2rRiWBORrBKd5GdnCO0/7LyQtw
7c81ZbyNyI+pBzMHz7daOFUSHUkYoCqr+wvlY2j1YxG9mlBFzkftssOVw10L
QdmZtTm1d9Xnc7a/F/yZPxUPf9j+WsNzliFJ/kvHhiftnAAi4ts5h8gqe5BQ
gtW9TJp8+hVa19w2jYUGDB5fuRZiXocfzDZtfqD9sVluZR553FN0Ak/qZJJO
/P17sO6PaeBMLITg6n/+YLM34CiDZPjrKPp4+hHgi/rUTz7s3v7ohRIc+7KE
Hb4DMpay1myHNfMs/WFoe0OPiFLYmpKiKbEPfn6ZHB63/Yz+RFFIhdo4ono9
reMz/NQ3Su/S0KbNJb+WNZ675/sdNAXHZGoFEiFJFdI9g8skGwaE8MDBuqgO
vHOlf/ef3cLmUCHPEKjRSuxHGie8965JVwI9LLlSTtvbDdnNa2bIgS1lP6Zg
alW1zNT0cipAc0S6a2X5mlV3Hy8szvp3LGcuSzDf3vCJaFl9Sr2COHBjHwfs
xK5zjjL8X52LWO1A3QmLH4l93NL0J2XaQBxbPdu4QX5DMJ6Sd0kdAD1aUHZM
ZwyjibzdyLzYO8ZaIWtCX3SfTh0bM7li+AAVJ4I4rksWtKILNEi7Kx7KHbrD
qZZf74xcBCnxqvE1W8CItkhYXyFJiVZh47hRWtfGNAc/ZCntyS3Q8bzqldXx
5hKXGMuU3teWmh2p2hbUMwNx9qw5AYtJvZFom2R4/a40CMZAO59Z8kTyMeT/
+a9MNas/NfvzvLB1bUo8hOtffup02JP2VJVL4Ab4yqJvF77Y3YUrHOvq8fPD
32FEEqBFGxSbx8wD3gr3n5ZDSecP5rft1BKApUiVaCiy3jKBf3Ds1iYqo0i6
i8ZoQI+pFpSdQ43P32jn2HdBDUfEM7OOuS7kvooJA+3O3u11XCRmVZmbIY6l
wRgpvXsAH3RRrV8P3cFwnQw6n4rjcuxJTv3aidOJ3hqd28p7kVnxGDEYfuh/
+yj/H/fOoVix8+sCE20bHdneURD0V8AzzMQBctLVKfFPPvp9h94yh4p2oOxH
8Bke7p5l/4ZeS1kHKDN95Tlfz7ESGA1b3CwSn63ijEUInGWKL2cfi5NQxun5
Kj9NNIL7HF8IXTDPXtB0MOOkSWcsxWamFgD+xQi+x3wtuKt2i3fnwkqCLc/+
XNhQ0/3rQxTjGveIs95eGQlsILS/c9Reac8/Zc+w8woRyfimNrP5Ekh7wRW1
ffP6UPt7nP9fU5xUMczpgB8J6eYFV0ZauTRz1VlnBFWatP//GtO0HX73E9zL
ei2xbo+1DHeGfse7lNwDJF6WQ1k7aHWNS236vJmiQT2CqUT09ElYQDTyGQB9
/iIAXVALaGcOQqniN9xU0Th7ArBEKq68xDxusyqkIdWupP7kXDck0oa36Nzv
r/xMpMQ5YiRb40aEqy0dcGlhZ7VQJLoEPO/0MAzy6xU2j92V5RnP9pfbsf92
SDsJ+Opp9o2Mijx5JgDG/QKwIAD/izhsmNlHzCo1hEEdaJuFg1ZXJFnsOeSh
NbuxIsRfBvb83C3uFjlvdltk+PhZcl56pOxdxe4PSZzj8rq0blUZr4uo2qsZ
r/ex9ag1xKcwRYQoE7z+pbpXjePSq7POiZEmQ3YkmwUe1pqk1lWZaU8D7cS1
sihvVrpHHqWRoj0VnjH+32syHDsBJtxEOVW8C1K+jAiuxh2wPR/gv1RbgTD6
zO2rhQzrrPTJzVyedHYyBR4eJmQ7NG5817TEsRpPmHqn1javIcQRVBUTZipi
LYIuo0b31zKW4Leg/GAu8hZURfH5Evknr86g1ka09uwoVXuqluFbRRaLMqT8
6STpe85ncdX1zOkzexhy8quC5EyE3mBzDIyIRpwHul2ipmzIYaKTndbR0JlT
Y6N6+IXOsdTEsUE99LAfSXwN0/zuVlJ3LnmtKBq9MOwNuLhyUPzX3Ja72MOQ
NQDb5UFABDtoD7X73iSZtNkW/59OIovqUTs8zoOi92fl+4gqWwpr+fgvFyAr
TEDSQIGVizqnI25XSdqnXKdsc2bn+bB4QWZr3bI/yjgQBqE2FqdfNKwYDbh2
eujkvfFHExDDatmnxHYNlH8OYy9HdRQDCxm+Dub98WPpo3zx85f/d1LDPY4I
n7QUXn1D99CKY1GUV8G0w09aG1ZdbVYPCioNq7O+wQEJ/uDBTTCdSdCbHYPv
h9kjs0sA2oj9CeHwk0teNMrD2Hi9i7D2gdcSlpDJz1yzlV0mMWILqgRwp136
KxyV8CK4hT0e6XeeXmhuEwsJKUt7QqI3rV9CHVJ6KGa88CjEvrJxiEvINzNj
i4uDtWdWpsrjWdzNpxSfONceqVT/nsdgooeWxRnJGPYxr0ddPxZgcDMPhOLb
nAurFCstIQRdVEaHGrRcwzXu2pdVLCl0eruxWNADo/3rE0kABj+iUb7Xxgu5
lDmtB+FfvRWFlxWXjTptJf1+258BsexuNaIAHWc2JD4HXHEuoQTuQG7Nqhwm
U1g7fglTxLxJnjBjYv6Y+bASEpvnG9P7UtOCaKdQ2wiGh04AXH/rE/fWd2EY
AjSTIXw+oTBnVQ6+pUgHvR4QP/T6Io7EWveP+SJsz1+5yszomnQ2BzVgb/6r
1sfKg8mMouhq9quF9mjD4MYXW/R9AE5y6V573A72ZzTE6A4d6oEM/vZm7Q5a
wVsDeFtm0FsFZKYD/K/AjL7JNNixDrgjAn+k0PlPHZMkVSWI+/GtG5HKHSNY
U0TJGvyLAu+U1cFh7/0U/4nABpLLsnNtHv9+zv15vK3fyQvX1zdfwa1JIb1o
uCS83fSItF3rAai4Z6KBrNsyEnfPBOVKiigSOzFO0Tzf6CAZHtcW5nMVyji5
gxuX12oqc1zZd7RfQSs6rB2/hBAt5rar8fmPjYd3VVF6hJK8hYJEQfOW45X5
bxOqTbC4ZKZOojBNKIqHAXZDz2YHvr6K6v0yhWI3mp7bFKQ0nbHF0BO1fCnC
YdhIbgLDxHhRGB//aIhFu5Wvq7d49g95cyfFvU1XO+Ke3aAAU/CB8pYvGfol
DLDZuJAB3yZOQ4wTyLF47JME5Wsi1ORP8S4cdz5W+shIT0IguQJ27Qjxm6mi
wCjYgeiEiv8mTNpu5EYNKdvdQWanpIbqPGSTPH79VQWsy0HNSTnRIwgbYYtv
XN7jHWLSKvm5Owa01YdyhWEfifLg6AUlbKTImLEi36lwGZKA/H86/iOZhB+9
A1MKjfi3d1PNnlQyFDVtWskVa3tNZ1NMGQoCWGQ9gXPThao+Oga0iDRNb8ei
ikOEhHedKbyvj3oGn7l2W6b4iRoTw+I9jOtjVcTnXbVGEqLS2QOnSnM7a/91
DfssRazFPS4zIYId6xp/TbibiqRqHEnX6uliOw9hjH3Za3oDyurSAYt1M8s2
+jXiOyPI7nWgepqNv99MRGxVMHFcCRvSm5nDfWSx7dsOGbp4nEKFJbXoQ3SI
RmJ5/FrAySoZx75FFZDvwqVGW57MhbgSDAR9JtL9lgxrVs4FT8vUMXD1qXzr
jRItg12lLRrgSBMqpnmXrdLXb6nNkv60+0S9g8PvwGTB1LOzjQS78kjcuWph
xYLBehq5JH6O1cajMfgOl1Wkgc/IJ2cFegatpKTrxY4d8/fBtwN5IKj8hjQg
sf0ZsjiaJUDA2HwqyusxaMLccXMyje56KqneyVsYg+d+qeQZPVUB0uvV/Pgz
K7CpuPu1WLc28HoKTBmtTd8mq3VKif0GzYttTo/ddn1PoC2mjJwfQbt5HMI0
WBpYOPqbno87DYRXCbAbV3dDmagRSfZ5IkK2VMAYouo+BfZBe9ZalmzjG7MW
l0Ac03ji8iRtML70bNn7t0VZ0VXwvJIcNJkjUWGYpegqIHVLPHoqV4q6jdDt
/cSnk3W2BTzL2vja6DTCD3Yr9VfJyttuNJO33rJRGUTbFL3zA8ed7gm0umyI
zROv3Y3vUy2/RFigZpObdAMtLV+KvKmV/j9Hkkuc2jzK/shRGlYc1vRdiBAN
vOZQZnmCzzDI7WEcwadFmQTL53J/VLCMDfBMJdjovyPodKHLgRKoEiXMpYDf
lKFsYbROloCfURyG5kL2bEGKBwCHbjlwYS4jM5hXQOph6o3omI4lcHMoKAa6
LegcI/MAjN6LI2/rqCApdp64VbfLWaNBcsjwgIp5a4xs1L6T8RPYjCs4OQ4r
bpKbLZ3WhuqL6cybzRVQc8iT70b2lhCkpZvxyN1fOfAz+UXjPbZ4tha0/KH6
qp3ekje5n28RqrRQTug5lsZq4cWU+RfT1ns+m8zoyctUpaqQIFtRItLGsudO
dMkTkekVYh2jR6PJ/Oe5Xml3hEV5oKhQ6132F0nYjSeGXF5uLEGeN0/VyJqw
o2/8/gz4pNX4Gwwcsc9RL+SJ5rjKNp8R6KMZmy4y2BfLD+zsoUiUY/K/3bff
DBa//PQaVdddzTPRtICduFqLETbZKY6NvNz9Qlwmw7BpOjOj22/df7+rbIGR
1ttgINakpYE/uUf+z4AcibISrwT+ODABRnGIJPU8qnUeWsn7cnK55zar2mx2
ZLi7wkT3wtuDGfeNP5csZLNSQ6fKhfWzuDazLlG3rczMtu93YphifMPwRDrq
2Z6QsZTeKtElHk7pTrQUA4VZ7CINA2DcJAVoTVeOICgHuq1jvp0ECj5B+GP0
kEQOTI+hFBHnOXgX+2gceSpsV/oqTvjj1mzKuYJeQTDiQC9ciSjh2hF07GXc
YmWJ+03CmbzHeLEB+bhcpVmmyoBJlmEbh6NY1vsJGWRG9X8RbIHXd+OmC5SF
dkRdqWLGfLkO+HmMoqglutZZ3CIaqivolz9t1oVevkWwNu5w2T4KOaMP1rQH
4sKXRwyKe4kUzRU2LjJDg8mAwrKBskBctjJuPk3vv1JXyolAjnxaJEueCIvA
viedpP5UQQgSTP6QTh8WdqFyQn+DoN2py/OtvxqQ3mAZ4ioLiagr8RCxxLMU
ToSmnYsqlRFXzJv34JKPHII4TQL4t/3di6C6UsagG7o5YNOm/hYYakTrdR+o
D1dcu1P4YAExExHjqaPczi5rMTo+MpKKPdLUncT6lCD5ZElA7PSvMb9WoRfK
hLfa7IinSPclcw/YPJUG0nfBPVpdarTQsI0FTrQSd5e33u0N3Bm/g+Gg3mSK
FqF+0krGDBwzsbdEYa0EReNBpWK+9k5+VUmUKggvDaSHIWE+oW7DR87Cm289
lyPLSuMc9/U4yEPANFBNQNRJUaieOI7joHNapcA4sSyGobRzqsvyx2mt6hDo
baK9iOO6CIovVmWhy+IOwz7QI26lSZiPTpJ9SluYLuRl7/p+qMP6S1rU4hYk
OD+Nu97F/M3K/uh+oIai5Z+WjS2gtEXOd28fiydG8d37QzArEyTff/Y5lTnB
nAm33H25NpXK2g1LQFvvXNt3Au1Sxr9BJQnpOVmLiS5Uda3Ydx6usKe5BnGG
/VRaXfknku6/tPCZwmn/OKuLDk2FwGHNQzcGY6i4YwnLBLzPAOiuRxz24977
C4jOym88rhbMQ62VOou/YU5NQ4oeanz28bbntDxPS8AMlfLSW47eCZRFPcbj
88voN+WAf3zQ0Bj7cV/r+8B8PQchooL5O0EFD9XiK0HvB48gfPQv62WJJmOT
ohEc54JjwbaIZ1a7G2tnWPzDTSeK3uKb/bCSyCKzTnqJFpMj0xUAa5o07Fn4
rBcVpjtB0DWh8Z5PexiGB+Xtx8Krsct0gQP2Z4Ev3lxlZ0CWf1kJjGD5wuMY
hCCQCFYvZax1spG7Zd3rsTQx6oni+b+yy3stS42coOM1Xe7GrDuPx751we1w
llJqFnwSyizxLsZkQ9IMtjersJp4mllWkl7EKopWuQYDjCmlLxMIqyZ1txdS
cuMIEOH+NErsgn4Vbhkb7+ASUNX8p7cd6dFjnA4anj9pK6L/ljC1Y9T1OuUA
wigUaQc61MZdI4EGqL3jCfmIV0drvUqhXWFetP83h2J+2c4x7AMlvBFN6v5F
nVxnFWYSg4UT/7DwLU3EBpypOH/PS9rdfPQI1/JuWdmSySgfqp/LeVbKqc1D
Q9fJJJbkvNJNvkp9C6y4sAjUCSRxAoi+x+FJzW8vf/M/5txhoF0L50CTPEDe
bIbMymqYdrlY1FNUW5OO4IXnWBGtAIwhSI6oJB0ET/O1wdusG/I58/eL0spt
uFacbYEznjMW7FeWGlzmqHet/EjqdQwflMwBUSQB+WMmAnj00AausNWHeLDG
ISUejnkkc+QVXo7SnwfmKjod8owZ6x5lOFAj5Bc7cyvGgS/7uwoE1yIkGWdZ
bUFkv2UB08sdfUs/uenj6jXx3+i6qcHnzo5hoGdjfvxbU1YOl3ohgxvjvTd8
ayuNHSXzj5X09eW2o+NjvWmF9BDCrfyuxbfdZAT2V0szt7KjJHhKixwu1BqZ
Wfk9bPjszWLvBkmJkzKEBlsV4E7o4pH3QHBcnAVHZDGEriNfDEc84onxYbkc
p3f0utxb8bc1fTWTsg5gfhtl+gwxsS+1bzPB/RxhcZsFGE3bbg4yCNlL36es
SFwL7cbMprfOnqbDNBddOvWfv/EHaJYlS7M1ttExxyO6fgu5CbPUcMoXmyMt
c5nLvbTChjP5C9BkvrTP3ADKV22e0ltP/5Pzj1WzeusAPWjVgI1M+lon0sJs
sLYsHfQ7qI3BddvkBol5ZSzh9XiQJ9dXQPd5ZJlg4hHOjIouZHf0M7kobG5b
N1Vbkj1samhncytgA/srLUYh+YDsYvYnCn2p82qWVwceOJfLLmkliwz3iXCk
1QoZdgX/URQK4Dpe4iK1LPhLPkrzDIWnFsT9Ofu4OBjSMGcJXBhZxnzK6kcO
Y3kX3V+r7KXyaN8AWV34gO6mj2ekbOpVrsX3qgydNqo/61kcDbA7V2z47dBs
8tTNjvOeN1eQywFQ3joX/f8QZ275nP8CskKEr8pkf3Dnj6CH6epreZrUmAPq
mDfVgVnIk+KuMuQeXYQsCeN2CB893UJASYhY12jrsnKrQrpNGECOTjlw4PXN
cgV2iQWwJ+dNX3M/0gRzUl3UNyNJcXkz9WrZ173GRnW6iT5KVxKJHQn1W9et
GkaeTidph4/01xEDxUb8GNJsjcsYQItjUvOWEpF34Q6Ict+Dev6qkxATPCga
Jvtjctr5/Oz1OAIAH/8Ij8qn7PEphJu2nRijYYYLQ9d9UejZtgToFKfEdcI2
2VXJA/u45BhSOEB27fighuVzuaWEHnheXHEKve49o+amYIPWcfIbk3DHkaiE
JRctngNqHot+FNrRqmMQHDHMsRjADKwb8VJSl1At2DlV1T4QYJ67JANez1BI
Hfxfhrt5n1lL744HOLeQ9vXvmVH54h+xoPuqN/JaLSIcUUrh4AjHHo/Iv3hy
PV4QB4U22kYWYmLq21JLAvvOr9JpI/FWhRZJITwvxAWLrINmAKfHDZPLapA6
yldizm2YH/3dGMamSbhWeyVKYMXnKan2ghbSXken09nMfdInbYT5vp4ulilv
ibb7wDZKFNhRzrej7JLOEvXJ4rRRXPH3upRVc9qA7uXsRXWmk44q35pMJCax
pGYLATEcUgMD+Hr06tVC+o1xMN/kNZ0pnfWqzTWM0h2h9HgLVVL9iB9qDPSU
nYJj2rTaJtirbkEoPattUAYXUR9/qADJFDFi+JkW2z6C7P+Em84S12PocvE9
0uO6gqAGMEAVKpWOCBIUP3zO6HeA26FGcq0jsXNApd9KFtsaQY4oQ11j8qqO
nUzlfO0v4vX7QGu8QD1P58xZ1Fl+X2U8Qu/iDJdHtku98PuC937iJ9hsaD4d
vos0v7AJyk6m+aCfMadlNGSXOs7z4t7801ctFnEAF4lgZukIZIUiSVb8Rwma
/pYx2mZVlLXtsLmjX1Itqi59r3ie8Cm1lw3mWSe0EuF9VmtdaWAmUjlnfilh
AyiPkniBd8agFbHxX2QepIoGfgOZZlA1a9Vdww0pJE6t2VQPu3a6C7D2ofN7
YUmPIPFiAjDIvEDnxvdrC2WQIx2LkzmWJlcru60eZ6jVkzQyGTxLaY5cxaXt
Wro1f1aomj8SSNNH50AT/VzXy0cJwvULL8lqcuIvfC6iZmS7rbsP0f/Pqa2q
zwzWrtNtspVwdnp/Ugn3UOYl/96OjIAZxkUoM0ZzenqzzBKOA8s3fa6lvCC3
JfDCfnNGk8hCVCZPHKoXcdpB/IkByThxn0IDR8SrTE7stGmgFLJUyzD5knrK
M9fnPpZbmyamdWoRlX2KL7Q/s55LgBuQHBYLNhEw48whwdJ1MikGjyTM+BKF
P+UyeRLEnUXQblklCkS7Byx7BD2tA7zUk9omOzT3tbbtjYV1sDBHrAY/RS1r
sTAf1e5c2Vc1ucesEEKgj4ZLUf8wS7/Ag2bBssJt61RgNAwBzZZsDIEeDXT8
dxCuvBMrQRJaQanlHo4DA7ctfHTPjoyeS3GQGSo1kjovt8rbo5OLyfzaU6OT
wsOj2iQvRWKdyY9flmslftBQPql1x1S8NoUxbzbD6tcscQdzWBvMxV2bVUec
/tgMc6gLfpJvwtyYHwofo0Su/PruYgfxPCqjAo2PBx0qEgal5gnL3d8S32Ph
B49J9b9gKK1vIY2QvFUtQle2fmMRfqZKe933UI+1lmfUmcZmlutgs6WYfAqZ
BGgOmnBc68sv/FVhnqDZFv7OHn5I8gKYA/VBxaB1WZmNI+Q+3jfLvQFkguGi
podbyykB8eFLAN8oYlgYVF7ZNOhzEFc36dt32LyZr/rhXY5NnJD7818syvyz
4dUI8rL1VfcW3WTt8u57wMExGs5qplU9MhcQzsI9ftpuq8XoQf0Et1Ba9tOe
STppeJ3MaEHExrdGxlYCbKKL74IkWYTPCj2agpCyodgSY0FWqXlZ/D5Suwy0
m1dArBPtvZyHaqoEviMubA7XxP3DfGrL9Ygu6aH2jL8wwtqIqhPrlcqXkVph
4zZpYoyAnTDd0puUfOse+CBcOyN5b9zF8+HFIsMNloBU25d8rxZicuyDTwkf
9ufmE/izn4mt/cepshyhu5WlG1BRe2+KaaxMuBNXwDYoP/cQzn9ADHbXDq4Q
Tec3gsXjwWVsyHwSfY5EWQlDrLsRyP6QhahQGSD+RoPNjtX93mCTeSsKXxoD
Ne890uLW/GA74rpBnixktngMUcceeutt7fCZuC3mp1PAx2j+9KnyVRbcWjRd
95LG2rrEmiAZgL1GI9Is5u/V3wQFx5KFl+YK7cnmkKp7P28K+is0VxIl8ywF
8r7PA2LKn7T1AllhE0WzMRO4kBmPOxo0xWCysnf8mL+ghu5n7GpqwTqAJ5tB
Q5zQyr1JhA2ZrTic3Z6Xqp1a2VFzLYbumMFD0fcJYCS++hmCF/4DjGEWP7L1
k1/dO5GXIU+ruRurF45l5y6SL74QOJN9DPnkjG6L/JCwF0ZzsGuC8gERwFI1
AsLzhwfzU2ZXUWoLeGzr0L/A8HkxKiA/OE+8flbowlN3UxQ4sCODPv/fT96j
HgH+xKJ/6KqA6yi0ZGvToscqMJwozRyJ9me61J1Pr3m/RIobIL8ExDG0dNYQ
dK76c5qOSxeP63e2Zh0tfVu4wMcNpfs3hYWMW3hXRvghKCt16Kshql9X/U7V
w5oVx9JwtGlP2SzjTzX8vQSP3BEg4Z+rwhZgRbQ0hPwo0Z7qL0oPjLhkhhlH
X3AQOZEzQEUYtldZo1FcSbwxBdW0X7mHPmsjW05do+Ks9kvSTSsziHf/1dj0
7PSk4hkmgmZORM5ql0ORDi8y0ANmr9oSy/1S29PvVQh34yZdKikDYeEzZtkY
21D3aHh1O1pII8Lo3elEAx/seTkTXDnkaDszQm7/h5eYibsLBqSVpIpR6QLG
hbyfbD9wF3VQOPgK1+VKzNDCZlN2x7zP+Gjff/GEr+mAX435gO59C5GnL2HI
42XyDHwM9UE5RzuNc5isIiIhuPjqrHCoJauKJCLQ/sYx8MLVPiKCouyi6qp7
Jj8s/syohGS96950sCl+W14JvbZdx2k5q2qwELXr2q2tZxxsjNB1vzbm+yzZ
HR5S/9FbpcgQlGr4vPRblLKFQ7BYMnBtlzRMw8S2B8kPjwOkhRFlDiC+yOD3
Z4H5tvckZfG+6iPhRDTzO6qAfchk5U5ZAXa7SwfPwDseuZ2s8jY7yRkfucqO
J6BEyhNjYak+wBPqowcpk9ClJ1+7IxoNTy/nwnT1HhB96XAdqV1chie/sL+4
AxkHrYtrW1NzHpSzUkmeYIaICvca66uef3+gbuPEB7FLNeVo/4R4Wg71GA7s
tsIIcrPMIx7xc4YqwArg0gUzt+GRV5MRbgZEuiW0shcslxiQYdIr1YbXtX9p
nDj8BzKtGeuVyW/bX90dcG2n4GK9BrFHcR6T35O59WcpdeED/OzL/71ikAno
1/b2qePutXXVKOSWWUgFcy5nmUWp5XxuFE7bfIBfxryLR94TikQbDkzGq/ue
KwTkP4g+Go41hzUQ/DJ90K37nQ0QnDH9N+fDeyTvSB8SoRyOLLDarNHH/zBx
GY1LQ0XLrjerDdzehdVObEf6y9FA741vP70sKabcvm9gWue1tgMB+ZWM2fbG
NKDnxIaqcU/1Oz3DyYE3g+Enlu/QKR+tULUr2ehXdkh76PtOhoZBQnkh8lpj
aDXkn6ECrbc72mHivz+UA0m6QQj+xrHOQJaxOSijIa7fV8e5UWjuV+DD1MH7
saqYzaUPsAmZ+Y56JgVNJsu+SWwyha7ef7Uh52a9/gb+y9R4nRKfJqJeffgY
HZ2SLLQzRDEwvwvnoqXx7VhQkmzgRhQBJFwV1xoUXijhr7JHRoW0h0Vumncd
/+gKIyUrq5ucHba1YsHrLljYto8jO+H9/GiCtfSzJnxWw8/VcTfJeFJJBaH5
6SQwDDlSBoR1/uh/WjIul3gmY/MhwDfzrgn6ACEbloOHy7MuEnyHhlGyoRRC
5dhZ3kZODwWzyH9ewhu3KDkpYxnmyfW6MqI+gNCfuDNEwumzDrt+BmEorS6c
VnNThtzqY7u5IZ1vqr5paraQHb9DBxF4wCON4DRKwYgc0GgT783j5QQ+fqYO
9G9iqVM0Y4zD4QWMhITq17YZj8xW9d9r5M5lXSLr11Bo26CeCJEuEGY7eq1Y
YcyAGPCWUCX1TTbV4KpW5YuqKlHQnJLpET3yIUSZdq8UPf9FPOl5C+CbTOdC
HbM+rDgW7b9Ob27whZ7rbz6NsLLmWvTVJvIyQkrkRrj6aj0QebVeTNg6tPQJ
CE8ARH23Oi5ZjjWZ/wqGxJkp7VtF82SmcXBTlg3D+tiJZj7Zxv2DHMrrAndE
nvTRGIhzocWEkbCO/VDducf3BK6IyI++74/Huo1QKrDH3w5MGcClsZuABvOm
tjVA6ZQ+kl/nNnBJioFbDo5s3Qea/Sx2PQBiQOXa95baeXkOsPfP8/XEopII
d8VhWuFiX5SeBu40JUiCmz0rGyGO4AmUi4LS87yxQJy/XbQ8LIViR7PKgaIO
WpHI4mGEJRKfMrVUScB+vYann2RnK/Z7vRovZK/jrnFqP5R+f7wws6qz+sJo
HOVzV0mslpbuoZESQQ7pqZFF8viFXi2l/T1nJbWuWDiGrTyzbptiuyXqQhcf
wxXkzlos+i/2PizCO0YFzYBJ9quPoEU2JAJ//UV9jkvWRqrHZpqf5EGbLDVt
jLgXv7S+YsGkgYVAOGokvVQKCjdXEVceYMjT80AxaBNoAeZ7HhxM9KsPOfuD
/GKU75vZ8IvIFwbpILxgvPeL389yGBCXA5RXEWYhtDQX/reJVhBKNgIlpzl+
q4qYh9TbMg/3d0D07z4FoFkKNbgmlcJk6SFwmioTg0KwBqZE9TRYfFqxQRaq
QX31rKWbFQP4dYSF3uYJdb1PKU8ZxqLhNfN70p1/khM9sQgz8ZqAinPmH/DT
Q7XZ/YrhHcjBl5GSCWsYMR/dR+vHxMDEwwbdy1oz+MD5pQDYA9t75MMCV+bD
1xQVayl/uHfuPiEfiCEgOfqUKleKc/A5jEhFINxKV8fimO36NOAFqv6OIQth
lMoP+gwUEZ0X/UuNI947EPVxImfjWgLnVndx+HsEBeu7gy3XsE0IDfzK/q2i
U4y5q/kf4kCgN2yxf42eiXz1NttkNys4Y+/zcMPkPkhnlqp6eFd44kcikfdu
JwqRw2Ku+Qq12togXbB6FU/VZy7DLBQoZUAtg8gAaV96Dw9dQ8SnHxJIufa1
IE0ubFB3Lcl/QvxmTFMyS/Pg5svwcoZG7znomxVkPBbDv7GRFJ/TC7egBYpt
jixadWEtz2bGQ14mq9FLigsNbTlB8mtaNiv9QBuKhMpp4rgYNsFAF0AoCtWP
4JyS+Bq4OgbuwcDpTZNYk6eleZ11Was8kts6iZB+7BEqQx8dLpDYUjTTiqru
PVqoM6Opkr09qTHoHz47vBwPMeRANpUiRfuPAQYFnicJ+SrhF2xI1qHgrPnQ
uZjBbatitCYkGbAnSs47iORjEkQWtSo7E3VKD5HKVcQ/ZWO1sditunboYVAU
vAOmnfe83SftKeov7aa4a2Zz+t8p3I/Rz+Kdxj8aXYSmPgn4iEJRHy6CMnjf
LuIv+7zuMVTwQRjoyZKygNrAOE9c0HxiIj1QwoYXEoSF2fJPQAjdrZ5qlzdi
ib7DFrAYWvfUT59E0o9R5yFrGlMxYJZXSUHsoh0Kuz1vSZYulb5z1sd3cb4u
SHmRd76hFAn5B//hriUmBWr8NOQWhjj8Qsu5JmcHwe9brRNn780qHK05I/H4
6XBnRor8HxPf9MmId85GQxIM0HiBDgLvsicYfGT6E8lEWei5tROZ5CnHUhsX
KYHrATFNAvHQNzS0/MOApxcxbqZgGAhcaaAwRR+9d7d2Itb/ZGkG/E0fRLGv
MRvJuDa5dlVm8Pvlyvd7iU2AOFub8WYF0Q/16M25/Vio9/h/HfP8A19NX1dS
D8JSUKO/brdGLV1rmoVl2xSMjJm1NqB2x8iQfVOVXYs66CcSAlzwhXQXtNH2
GFr4Jza3//J1qecS/nsV3P5zV7JIZ4N/KiSWBNnIFmXQ7iQPkDI3IROPVRhA
g8ToS181iP2VkUZeIjICcmeT0r1PC8OQAEm4hiBoPyMKUirugg59qzjvGiIA
CpBhJtwCTAuV8rVRGt6sg+HKQTiYLndIKTeLFGFfHft/IwZR6TfL5oMSzucW
+nyLfqCVUeHrz3yupPyTq0W21TCntpB98llhEBg893nIi9je4BqG4a17yX1F
UjvMcqofR3s9jptPkH7h1lmu60XhTRyk5mvtv9Lx4LhsMwskZfAdNRXHuzon
uGqiOR/M+ek0dylbVnZWInTI8PVoXbQ6E+bTGxmknAfWXsgQ24QN61u3D6Eu
2uU3TIa++ocVSc+Ldb4RRKTN2fvKyCclRinmgP2g7bLcnFI0VS5cPwstc4I4
2Dc+wLYo1PB07d4mOvo+J/kMfwJ+VggI4zWV9jFZLzqDOnWBJjPmGBI+Jhya
wUCc+oGsZgdW6jk2qCAmqmWFmSv/qFvivndSg+ADwsbrI3RsLN1gFbqWEvr6
MddNrI+2Z04BBHX8MmF8acljTDisMRcR7dZ+5BrhvptRLF0ibD7ZVcTZGoC9
mXdkYzJHHVrM+uTV95XwS2BUB3Q7KsbB5iXit2NfH96toAfJRHG9OY/56tSE
fsFIZn75MfPx/6t7GsTYnrbA1ey1Dv7WV8W+8iz2sO0rozk5KlazJ++j2NGD
gmyQyWy9XccSi3fY81f7lNXjrXiebdlM6mU0Gp5zQqN1ynS1dPv7AJCd7wm+
12BNICTL7dQMkCsIZ5QbJiBLB+y4v2lmPp2q70FbP55WOE/zK1di1yMQWwpO
tYDr8+dQbi59g7y8sz+LffLXEOu5tFw08zsgkYEt24Mwj2x4dZ2hyJIP24PE
TCPiQLF8hEUzVQwH06y+mvMFFb9Jh0t8Hm6ICAq4yZlaFtbe7439enAKX3cM
v0eqTJ/erPRqIkYGt/Jfak2YsoVEHa+44nfLGHxsllrixTEcZubnc8scMPEB
1Pa/5/UyHSXs3OtQLZxXRbCVWfvyceiVaJ8OKS6SOGOmCF26LEYPfBBBxEel
6mW+HUeIfSzIlD6uQBFpuSVV0MV54oITJxawtkFSEeHku9WCu0mhFl7EKaZV
9b4xusoQTZ6PBQJ6kljdPBpmD8bk4LuAEzegx4bdUpXk/CdcYG5ZyCKkSSZz
aqMfKVfRp7ja41N7F6Vawg6vqaQdNcrhBOayy7rWnKt9M9v89M2woMEopkFE
f0FqYEMVYSTe/VjUAXW0S5IDPm8fDWuzV0mrsFqC1zJiWr8IDVQykV641EWu
p0sAYDZNQqI6L2gG6JCm/ui6Kx3GdQa8ziUFUKHEFqlkuZ2O91CvjaL8qHr+
HCZIV0DcVimHfhmO1CKQuYPapeK3PNagIJKpHgmuQhoOSea2RUK9SjlZs3Xj
3XxtaD4e+Ik6evucEOHbsgKCHY/9DjiNv+s/0RaiPQeazxR4E1es1hmCxBTu
jG+LWS10Mbxt3Iptyh5aVZQWbjkq4h+cFyJ0zWWtEHAEgLiIG1YOAXjBaFrY
I08hZftapJT8Bkzhrg8rwj9EeYGmlp/5wTsp4DlIXMKcjP2SPUkXWQCk76f+
HFxyDo5ugP8hDwCn79jRUcosID52CKP6XVjlNcR/hpNVTS18A/Hq7Y5e2nc0
KXK8ILPvLCFbL36VZ7VjrF0wn4iVVNWICYenaIgpy3ApLBhPGoVdH/XFeXtx
nqe3c6/TREEPc0cZxzAiCqpiJoS7DQ4DkSeWVvfREfvVUaEOcTv0HDIlHiN0
zQFt467+kGoBsNvkls0KIA96MLD+3yRiFPi/xONbl4l9kpRH+DZiKP3FRBWW
b7O7C2pUDGB86zJ82MWM/TVYZVQkIqgkOBrYAPK3F6oMBGHpunMopKn8Zckj
wVotA+1HXw6ru7uvJ5akTcLXGcM+UttYx7P6gMHp18KhSrsvCjaOxOVdaveL
TYvvliWEJBx2ypkmTEzZi9EukUHe6CPCVKW2cAqXSW9Unc6hO+8h+jy3r9ow
fEijFAjHFWf9zHO9fASmUxGtaJv128DfQ9Vrut+NFa7ekhG6yjQ415Jza/vt
OiXTWTXpiDWmgOP6dZNeuw2/w/FecqW9msp2oWB4zudPNPyAeAXGcEN34MVa
FczworiQdNmQVEic1q4V8yGUD9mbGPPXjxRUNb9TzzWZhf/Ng8cx53Sh6kYy
p3/hsBTD8yUC79J5vZa75wIBIsp+YqdLgABvoXp5435B4edO4X9FPDMMi88r
e0DyTDr2MzVPRyoxQslEr+vTCIU5EBVhsoThbrwFBaCMy7FT+tPVK0VmczGI
J/zyvELFGjgD5nxX/ZcsEOeaATd4QDTqG/0ymMhPETt/WZNOtnZjZB/lHMJF
PIMnM1EOWtH3ViPfduEQk8LEFZ+q9G8k/XDsR1AtM8xjYUKIq2NBlEs9x2PE
IZaeeX7GP14aOnxk6OCQDk+B5PhvziwogpWfVR072Ch4dOchDawObcTsUKCm
96CnRXWaLJTgj3kiiqbyxsaDajXZHdMFp4jnv0nAcYGKJVTsZ0HZv3so5w3a
+tR0BVrlS47fjoigvmSGL1bEpsL3uXt9q727UuuP3f/cZ2pc3nRwnaHOZDJe
zH/BNLkiceh3ZT2eN08tMZ4lOv97srRLs2QlWyH9dEiwlfqn/S3s9HgtxLFD
SzEGDnMbgA8hUEL7UjqURbIxkTus4JFLsLc8gHPImXcvov9QoOBX21w8huXf
0539ZZhKBaXDvB/reBZXC5zKy8GRxicmywt0RP4Q0KEm99zLL2b0OT810U6K
ZTLu8v2uER0AGEGIr5X/RcEF9+8nw/HGyxXlAYD9R2025ZJhRHgvD+dseS19
v2AjUlwI/iDJrM9+WGPcAV/f+0KG6K74bRiY+QyMcIRDCyt0SlLNTgmHwiEa
uCRWByyp2HBAazcv2BXApc6Ha8b4hu3/0C3rvlL66LafuU4JgNCIZUWV07Uv
GxWyx5uPFCLpVmUWu8ngj1c4Xc7iMpIzL580npIlV5iR3dmlnlhDB20jspit
Yq9MZBjtuCkS2ZfPHwEYsutuU4Sj1GT0XS4z6laemDM+aNOPPTMIL7IneA2V
F7f2a5COg+kmWycoev1b4foAbul7EK+9xoGlCceEjmpRQKeJfGF7Y9SSAxiG
iI/NIwfg5bI2L/znKKKinJLnVMfh0pZs0TMdUtQI/8wujS/wvjebusJTig9F
m7dIRO/1J05mD3zlfct29VCy6H8D0SNXKlbnpkNXTPNYEo4dB/r7yKC4cZLu
LaUJZ+4E1XJm3qi6P/gAswmAIGDh6EGBsZjS6/ATCJ/OD5FrbfI9+RvgDGp6
tEGjQDA8zMuaZzeB6A0uDH8qWjSmzfgAyaoK3IL1hfXAP9m9fkPs/ypqT3ts
O20Othv/sgs62eAVCZ39kH/uwxZ+cGRkPFNKAeydQELzrxR9yANfsubz0cL7
FLplBEvQ8ZdTNTX3Ak0Jv7DjDQHL2Syhd2dypslZoE+lBqt28IbBck+K5nNS
dGNoBwK4sL+GPfXbQOGqNMJdMn4sU4w0xq3xl079Va7kuhLsrENQDsc8sln2
Bt65/AXOwKgvpCyPiniQIMfEH/QKF6Ziq594tu9Fyq1IuOos9SXN9+hECL6P
vtapwqm5R22liPdjxt2Jjgn/ntBhW7/yk8co5JbtTb0NQXpUEQoNyWI85/mn
4C/gQosKBPW0osDaIEwnIPTSXZ/5BcOWSgLPn2DowRCcUlt7jibdsSScDDAx
RLehuF+AOR3S+aOK8Z8rYFzMSaGhh5tCxZh4io52VHiOz8HYEFQk2K11Qhp6
pcwyGicXjjEQnpdbOFE7ZAz5a6kJ7RBlhAYZSWcW1q4QgHf+4W/+NMBrdsRX
9KiYwMbgb7RLZZUsowZufFRwxhqaPKTVge2+yxTDUhFUt40kUFNbKim1iEB3
dNzFav25pXxRzWQlGATCK+nx62PWcDriZdscbe6Yqbr1kIaED9Taq5USanPr
ufmo795owk4pCBXoukpnCGKEcOYk66idww+si9adl0Sn2t148/Yfi1HoaIWj
UqnErRkTGpcDJaAVVf4t22iZO+smLJSC3erw0V1p9xchRYZbFdyBR7HZ3Sbc
oPNv9xJcF7vDW+wJHKiKeWv6vjyKBe7KwPvuT/ZoLGPUvRuuKWFOSGKGSwp2
KxC4+vFRF7ToSxK75RB8IXmJNIx4JAn5rHs4G7tShZa6ok/q0cQ7JeP9x48Z
s3EnbaL/Y0SswJ7Ch9QC8UPgthNMLeUS3/KabdMvWPDaL9fAE8jXeWfh8d5f
d+G+fAzILtqd/L+G7a0vRGKuhNhdbi+WSBRiJIyh9VwvBGGsEl0jmse8swez
KKPqarQKFyrRNRjsAy+5nt/gktNZXXLjmyy8gwqDY3Dtd5awOWfG+nWhQ0Rc
V0myxcjKXAzewcaULTwSLiKKsd9x54rO3ISkNAxSZnMSjcT50MQi6l35kKL6
p0+C2aA9mrtxa/xOzpyXjtYnoa+hteuI0otaRPy1+usMIDt9ejGe95RTy2th
v5kknXrIg3AnhOGY1ovc0H3lKjZ7dVo4eb4dgLz0JIFMULolDWQriWDEuhpC
2S14udKT8BayP4VBSGcOk1Y8qRaN34PvFqv59nODnsbofe2ErWsq4cnWVnpT
Wsv+4guRERQB6klAiLnT4iPCuTWE62EDcF9AHvdUSPpB2fTtsO5CpTox5u/P
xA0zgeOzqXrpZP1vzrpkpgRan9ySWzWVRX3s0DUrp4eVcwRSzZYYsdWiVtO9
hfVpEIPD5vgJscVkUbRT+ut95edtvemzmWU2Pioe0R0KUtLRFwR+bVo4ORnd
rOo17fXqAAc67rQdqFjIZGOMH7U6s8D3spDOaw3NIQQdJXwsPjcuuIWiWhiE
os0MU1RaLesVReVya5Yf2GuIW8WNkhBBIeFfGAqWKPBr2DifGVvgPob1+BeQ
rVSAjV5efXq+fRQ4Ea5mP/AD0+84FgMAuVG6RmwckuV3X0wH1reqTnyb9wx1
8ZZKH6vwzcfsp3KSIeIwiuS6WhXvV4EUMt4ggwgM2dOjw6h/8Lt8LGZQ/Ema
J0Xjdsiiq21bLJVWqZTR97plhVgSjUSGeQXwsml6fd9u+dSjjLBBbZrku2t1
0MGWfBUvqhJSREy5/mNSDE0GA5ov/8VtIwRdVSaImduWEQ3eU0vG26rmI5DP
yTTo2nF2sMNLB/tmkXU+vdr2q0TIt0IDaHSNdjf2/Ltgu8eUaNDCdL2DNEj8
UX3nvlkque9XCpgy1KpBXfbYmI0imHttcEpAwfCR4K3Xyy+A6XWKGU7kUGqO
n9IXMq0KIxuKyM4B0HUq1SMSmSzyNY2ihZgZ+H7lwHhR4917tqdEGOb381AO
dBE1CpD7lHGycTesqCWD+KN1NkqAFd3vHmZ6gizGvJuxNIcoEktmXt4b4wqD
YxxnR0yMiguY1VFY0f7k2NwYhoalc/EkAQKpEcZuizyT1HcKIFFlTaRlhedF
7+iqC7VfMPesB8tXwyBCbtFJRokbnlKOIswH/oTqrwlFtSZKZeHIgIu+ho2u
spOXoPKxzsisl9VARXuKYMh0n4GHvAqW55tmMsVOAmqHkIiPC5a1VA/+R0Bv
xa40UEohhXSjstB3KMeBSfJQ/omoklq2xmJHoQqE8wZpTSFesGp6mQKCE6CV
F3zEmc/fx3HyQAjazWiTLyBCzliD44Hu42AaPykhzv58Vb/0/XTuXk51d8+Z
afE6fs+8FY4OS9Zjkq54zapZeQTkDK1rtCXSmknJP82Q7+7+TriUls+EAW97
Olwa7Y9TwR9iTIb87Ltd+iAxkNr5LM6mmaS6NZ6j/5NXaW55GblNAFX5c5XA
2Rivn0XOo2KVh+w6HzlFx4ryxn7+Fe0ZcBBZ5mmdIuAvrwJ5GC9MYwbUyUlu
Bz1qfcOJDOq6HDvuSItAEJX6gHsXWtdmFmRUiYIKJJnOZnHj0NzLTyn5O9Ez
lfBl0DN5UKLyCp8riMNsFe+HmiTdiQzOBlrJLrpzSonvPju5TbEfRabEw8A9
fMZ8zh/Wy6vo64KDlKlWPTvA19NJ6mmkVWk+ZqSybZ976RbKpT8B2DA1ZhYm
UPd4UjOx2k/GPp2Q5laJFIWkaw8MhIvy+7o2hUyyjw9lgQmQT4cCZfoDw8LT
OeJV2LykZeDOP5cU2aXeVpf6aM1GP/+IhU88HTC6T7yWxJoAWniGZQk6Z3aR
kwXUv5n9rqJZFYtrDnwAmT6iFLCZObm8WFf7VV33DEcyolYyVk2JcfEOjfat
DNWzQY/KEJU4jJMdGvvsVfEIlUBCaPuQ8pqWFSYF62g3tX/tmYKl6Jy68j9F
+nX12IUwckYTqp9WU4IEe3ZpYMw58ITpnNwshveClJPo+mYAX6Kgz/ZvHjZh
8vbzIBHXne1WWbSdfGeVWMWhiRMvEogGktkDEh4TmNvytxBYA679mMbqL6m6
LSgFQhY5Uvc0GuYlm+3UR99S+PgizQ02GfO9pyGcXse5pMs0VK1yJfvM1yiv
7ZYQ1OQ94bbBW1tbMOo8lv8rwdL5r8R7RvcNm9BCqeV+Ya/+f1sIYVhuuTEO
j7sjef08GI1CaXitz3E5qT69tCIdibK8CL4VzTlefioSJTKCnB3VXi+kzlS8
4znAvhPkhwQJBKsv4uLBR3Kjy/7FUPOUOGD7otTk2IqC00Y2FqYSkOoVZjy2
T2jfeVicykUI9fZ8BePFFDyogW1ENee0ZFQZ47fgS6jTqUnBYM4y1wtcyF0B
PjwpFCWjrxxh5NLAQDMcKT+6gKRjtzDGTzigiGg6NJvNdRfQD3+DqEQq83hy
UA3GJ5vxBZulgG/a5ndvm9FM1YIn4RP2m64PUaNqW6Dp8Fm9gRT5XK5cwDiK
QgMmYEBR1dkX6kpZI1zzSzYPSEFfPTW3Fr/Pak2wS8JQIER4mGyEBNpppZjd
gHOEvYTt7GM2Yy+P2aHSfi5Bo4bZCqmic8bOBMGNipocU15OlMLpwdsQ2dod
CLnax+WHELHItqcMcGDykuUNCw8KKVqYM2bBafB0fPeLB479GmVc3j656pKb
mksE0UqFLSOaeQVkEy4m3AVCAEwQ1Tai3WSOvpa0t6kmiylsXg/sV9MskscA
7NmmKfThTcu4/bDn8tvCJeyKni0Fu3KRmRaeZwgD7b1Toj28Qs6Xo49fux5j
cLUwzoF1eCh0o0j2lMi95EbLWWHPTOXLvpa/wy7RfT1PVeS3YG8ksh8uBaPl
h9TNVnArtUAqBxu8dXoswVIs/q75MPXME51dVPD5Xwm5DHkOttnDo+CLnmKm
JajcCSqECznh+Ivxla1J68kAfa6vD85HnMlw6k0fTrHMdlhslWfIWkCsRp/6
hVXHph+f0E2zy8Sg4In+dDnUWlZchKQbaZSLIOFfyDRRmp7GH7KbY4V9/Bwd
7DNmtpwTfQanIoyhltkWjC2OkzTALlkYg5nXaK1u6vGHcL5ozBVXCLVxM531
fHSoMJljFWk19TBQudy4Kxxt7/OXlROpLwTIP7hcRpnoRrb1qg/fvIoMy4QS
sMCEoe5Axm1Pvocc7Tg1dMf3VrJM6F1vIAsAg8Dku76nBCTmtbjVmAlrGftf
rapyWvkkwYVrGmxK7CAf8v7vRZyblhDMH/Ak2Fyw7ZC7WT1i2u9FBnZIbyEM
W5vnYrnzX77gugd0VoWjIAfWjiUb4+vMBjAdblIkMgt0eANh+q+PTGF/NJte
V9SqF9qy6qn3KSa9vyNeK/CbhN/x/cOXOIPENh9aPTKB3c8QCO2Ye9wkRmE/
ilymVI3nbOdm8sROmMzM3fFFMeyHBkJxY46Gcmi2AGkmQ3uic8C9LksDTrQC
s9670uJ4Hqm9P8noCAq+9ZuZ1g5VLIzsMHdgH2KQAZnFEeQrdTng/D6j0eZF
fIVHwZjP5FOwJ/dOWYPbpNPL7pjT8F35MMMuCI5q4dGlI6DdfSBOYBkfRCwW
0muMgtiI10Vn65JLKu31UqlE9arQH7FlwLoFVIX2CebCf3efNG7QuDI81eAZ
GHT5B6u/xUlQO+aTlYZfDwO99vxx5z5d+jNq+KEP0ZlDXjo/7ERBN1DzdWGF
5KmM6YR4hkazsaaT+CuWOLovxKetiqld8nrLwvnfB0PtWbJw/r59rhGwyOXS
WRvAq6NZUCaO9R7rCF06SDKErLHUI1RUhT/WvvN53YKLtjmZvf/s/11HVmfg
Sa8HZAljFQudGmlNOHwq+VsT+fEq91CQ7NLf7it7GM7lx1FyXlWUGLq03s9N
lBgkTPRCvd7e7lU2K3vzDOy5zFA3pVp+/hFUrbDDgUVGTdan/cDhZd2XiUqo
B/zg4MndHlKQ/C29zGpcmZQsfF62gx6v54/GPV2GSkpmufSj4jyRZIpMlkDT
S+/TdzFkglLqG9Mmd5DwRQdqZJpHCCg2ZlbggQ4d60r7pXeUZf81EY80d0ni
dqX9XvSEvbAm/bKlmt7FipTZhGOPWDjqd3ms9nA5e93/OPqP0+3RDOhgqCHa
aNArdPJmgvVi7sMlm+ioJS9tqIRLdjLwdflL4oqLbl5KUOhWQmeiwka4d3V1
49ykM4klLTTyLjA1SBQ9NiGQg8dAvggSNEplv5i34M79bBcgCtbjQCxYiyAP
WgceuOBfvhgZwbPwpxRgu+ld0MPIXPSPKBhsNicavL/iBennqMklF3b6qy4T
ma53NIMTiRk81hJw3L+1MbK4DvfrnURQUPVsgu2Dy5rYu7F2a2PlP1YdEF6l
G/ZT+et3DxRKsPm4+5ICERzOs5bPJitt7wi2TL554c/4/QYhqzy48WxU9bJT
1UzrQOw31/+LYjmq1A8zDNlLYN994N+sUPjS5NU9rVgYhidrkPAjZz0gDZES
fqKF2RsEFJ9BRS9Umew3OYb5sjVULtTq0DOzR6IszRol7nqNKoC8SGv8BqE0
U3mrCJ0y/qKByXj8Wp9C3NwKyZDiIRNV+O4nQQqj22pRG/q5y0l4RzBGaSuL
xR6Ky3APVrK+Eddjy98VwfOFnuk56LiF2ij8h1WInV8w2iKMC8cTPXInWPrq
PyxLCpt7FY8f5tT5JJuGSGJzcodS4gUuB+llqVzflIWhGS349YAOxgWeJhAE
AqaqHAn4njmyYSpC11NWtgpTp2PhmrMnor6GDffFsIW2VZs+h5bjV8LbV2Yn
C0UFg6Eha8ZmD3paT8OUzGEN19vflT856l82Y4a0eDxlYDaj5eL75+C14s0t
wVIJpeVrfkOlv840V7hZru0PTY8EfZbOSPq5BAWRmAhWn3v6AAnWAlosg8Et
RYObAds32jPLRK/JQUPd3G6jNbjHz/v9tBvGqqmDrK3MoMdnoKSvUbhlMzbG
gUMNzmctFiBQ0pR1yCZ+ehJ9DDNdMwEiPgMCBLNQYhqIFI0VSZVThw5iDTN3
s/RZInTnydTAmGUGcjAe9qWxbdJQXOAqjDU1uuo/U0iuJvlFVpypEQVyHOg2
fJXjciWA8Z+MWtlFnlxWqj91QWKrybDYvJBlk3cj1cyLB9MZ2zhB52wYMmBb
j9LL+ut+44PQWp1ctLhqtNDMEqB9i58epSrCIJH0sbOX6gluFOnuNx21gTll
9SLBoaXHP4Sa51VQVtm38jjbYH1O3LTg8UTTn0pW17MkCc+3ZU+bC5WoKeSW
QG58fNyF8Fi44gxYHtr+ESUUclXes84lfogS4vuLi15TYGvNw+hx8beiVUDY
sH1f22mgIiE4yr72OQnMQC3QXiE6jub+7emkyLDIl6ACbX8lhY4OTs9Tn5jw
lXZ2xq4BPyUudHLc+C9jFw1GLS75r4psPrMPFCKIDzTVyAWE01cvSIrgQZ4n
uJShFzwf9IVSG39U7erOYbeZhVEGDDeGdofJVQpuBhLTkiIHl+z53jgsFeCp
IbhKgk/bMB0cZp096nB0VBepLzXZaqddjSgwzPJyrHxuKrXwP59jsOnfMPbP
shCTtlfO1AdmI9tjIHECZOcLajAjl9hixoV4I/KelFHutbkt64HAK1RU7xu5
jxBfrPhmelkOQMB/bNOfrylMbG+R7kVz+acxm6iHcLd6KPqimGxQHIun1LS4
QKrMc9TR+FKygRYpIcFDdsZ38okNVxEhkFIFAGT52f8GZK0WxW5kMXupFtSB
PiGVDj25vkkg5Ie79nJwmxcElPKLTkCG//ZDeeqyzozA3knzEdFL+ZQ6FMvz
oV+i8hk5IVyEPyx7eRtC/j61BKcSvg3uNHmZk9vsPjE19cGtMICDAjL+VaBe
HR2XniIg0k0qcB2WpEbZGaa1vR7UGSKO3QS3tGuUWzUS8bvGFrs/sy7kRz3y
d7n4G9+I1GiImumooxcUj6Yp9w6meLFThVYAsxhGs4ym322E04ntIHGFi4QE
5saQa4L70iqohhGn6rYdpPNy/n8FLXtWQSGaPR4t5ug6LOdo8rwcaBvN4JMT
XCpJxZAQU6FMhKGFfP+dp9jRNjB1fWPhZZbvmituGH/WaR+WMBLN0khVLjN8
FFE6QxDGBH7Z/PHCWt35/NN4/OlYXpEqRGALZedpdoN8ryf/SQhxkfP82qn0
Fzs5me3xYIzy3SlTHRXORSoWn7sc5TrkoWU9O0l0vYyaQOa1cUq/IR/Inr/Z
W0JWFw1L916vGBUBSEd/hXH3T/cm3sx7+dHp+FY/0u7C57ESVmBKeYWIV4d+
CcYqXKRdaiIRQk/lOjT5uQgVy1C8NII9hNC/1QE2lFFNtBknB5iDIXdWrR2o
Ex33/LLdzV2exYFU3VZaO0MQzqsM8qGiBVuCsSzX+RiTkrzGx9XhS7V88fBA
2H3SL23iHf/QxUI4wognfOVDZx5TbdGfBw2Kgbb2t+Ns0Svp/QO1b56/12wL
TZ5x0onBP9wXRMoYN5/syZ4lU42TE8M8W2wY1ImfKqMVpmFVHADPcTjZvT6y
28phZinCApPM/9A1Xl9o3n4r4GgzwWv0oiFIFvI9YleMEgB+5JJ1AKM491Dg
H1p0QI6Blabde5YQ/8PT7QAX/mZQHI17j7t+8vpfJntpo/Z/sOqlB+VQrxz0
CkeQI9Riv4A9wWdnhQALN00xVhQ2ZDouuDU5m1lpDNFEEIs/LTXvoKxIfo5f
Bj/kXuGQ3fXnDFsNAOveT9aWyUfxCrfEzWEXBokiPfl69mkMf31R4i7Yor/b
xaOq8Ji+JISphOLl3ypjcLJNpxJTM4uuHl7YjIzvFqT7IWqUWqzOP4ukDRlv
HLUYwOC811OBmTu2IBT5CPc6vw345Y4y53VUDaBku4nfm1OovzC4KQARKIE4
ODUP7P3njj5vU9VZsj80cwvqXOKC9wqIVrypSgN3wYAWlICscZWBnFu7jgoY
P4oY+8Dcji1fkfTmnheSX0X3xl1yA5rAuSM2dmkI30gsz4u0eoJyXQYTJf09
KJVdkqTE7HMSIgB/rZyyibj2acC0D+BalU2RwUXeen47M54GaFNu4nuSFkVY
llYl664moDjvAEe9SotLBDeZA64A+aamnDT3xRAd20N9IK0ldMlweLr2/grs
f/xoBlkRcw34OsZhDf4E1PIanpXRBhLEyDIYvApN1yeiRMERjhVdTzNriiu+
+GC2YeuKo9FlFUAkFZimG60vU6SxemVfiA8f38v70ZA01dT7kz3zWkGcY0qx
2NwDpPYkQ2FyrV4yyqM2Cnm6TN8H05Ut8dtcLi9UB4gS1SgQejhNtSBuY58L
co0KpDa8m6YHt8PbiEQ/8Rorp8zwRxJKUgC0hmWY6KPykPFAFFhqQ1BuBMmS
wpa+F77A/vcfiKkw7x+dO4zInE8GlubcluxqJlughrfyu/tt5w9GTTvYFMcQ
I+QCvRBLybX6aJkiSGqdwuhnLqWfBZWIg0SUJdZARTd/bu5aAGNEtzdegHJR
ldEdSe0RLP87j3YLlJDk+NdUzTN55pJ84f3XjuWM68G2v315I9GCr89oflRe
VhZN2e5F5qFXElS9V5xM6+n+z9pFQ7BtntqF27xM5ukvjrGfrJVk4IuBywSM
eqaeO/fkxHTzf9LNd/PPtrPdk+uoeSWpg1ZUwap5+ffHCKQEJ4I3HhpxmW9I
GxtrEdqcq1AJbQVMFwIFpgkX+j4BUqXHQidFIPgkVMs0coZWtBJFAWjPMM60
aFuUr8lMOax3RK48+cOGZQBnJtDC8fdkKzggMJTUB7+lTundlm8qD6byBYYN
+r/G/mCHFZ+dRNKz6ssSzhaW0G1p+U7IoLIx8OSLDLwh6mNfACnMpkeSe2vA
kwo4eGmrNfT+79O/qsIgJwG8B1Ev5HiOrsFG7RZQGGcem2qi362Az2VeElLA
a3MPgSDyilcm46MaOh6boLlZvECO1sYJ4T3MwxyVRzJV2Xh4I/T//eKnxf/z
eV8zJsCombsERFBdyULgpGfQ/vW/M1hqoczuuVfSPubGVN6GzCcASnPN/cVd
aatH8yRrAZLjy+lmtW8fI/+3opw2CCIHkNCaOApIJwzJ4w2LLMNETom17cAq
rBnzFUkgeU7qf0o3w39oM+VfQ0huvuCDbvG82I+cbbEWV5MP6Id2T5Dn7W9/
hKKKjui7w0PXLj6rmssFdHhLIeiihJL+VSji1LtpZYTZ74NpeNHAQHbV4TBH
42Koxi5JmIrPRbro3LLswBq+jTsShpCq8eDegNRF9S3MVtU3VDJLa6M9AVUq
F4/qdw8L9vqSK6ei5aHeud0RrD1U7z8Y+9q2YDjVJcIJTGf9FOszrsyQ4vqR
UhHV/LrNdgQo62Eh2ER/wPpsuGiijmanBZfRkQ3LWAk2yrgVByrEgh+zX8VD
MuHd9J8MCYklPeLzIYkByYCd325z6lOUA6zxtjdFhH+Az4rCRlmljqhBgu9a
UsJbNkpHxixC+qBgsVhQ4AIN4Fn0XJi+Irxw7k1G7SR0ZkLTsvsqvcOyyGyh
oTcnUC2z6umo0RtSgon9Ydza1QBUILzf4lDPBYXSm3fhF5E9P85AjhJ+jqhk
yDep4r45R6B8Y/pW/4lnmQO4m6FzDRHf1oqvUFZpUoJ7+auvhOgVQPVEGW6O
+gRjtFjEGQDSkXXUdVBli4PBL6WCzKf32xZNBWZDXx21v+Ormh6xtNxlFUVG
NDr7qo/6i9lnpMV/vfOpBj25nLTbUSIV6AG5hjvcFjzwAhFXIXh8BTZzxfNM
HAnrJCHaENUMw7etSZA3b+ZyQhFzPjVDooUlVfHEubnHFKPChYKIcSvAh/Mc
VqDbLYQSwsOziWNMsccjI7+u0rFq+qlaKKDCDiny0vGGH28hvv5VbLAEGVkm
XylEUVDM0fetUM//frzwpjnsDpwetFai5QHf2nf0c1DlJ843OtUsSrsyY2Ul
bzcthrAYumH8/F1eP7yYstjdt1c7VYyXQDfj347GsX5X9cvYjS9ffJpv3YsK
F8nTgz9wrUfywWlteTC2XojIVym8/W8lxOTTKkMLFqkrrG7tpOunOWcgAcfr
AHaZR5o71myPBJlP8VMf5Y3NssIdpLQy2WWWpewr7OvTciy6dk8WsO5xWGdP
1ZtbsMBCueS5LN802NhYEhaV3Qsue+Wo7hlU2jkNYkORqsVuLCB1Ce1umoX3
0ngz2q7HtuyM9LhA766WVimfVp0o1AbaGbVEsooA1GRQgxqAlsgnp6uycywM
A2iSH1ceSiDzg73TKHtix3R4QgwYbH9kfDUKVQxn5lif9+l47BKV4e8e9JLM
bt3+tRw1kGRLv1h7DrQoAqMT1ss56+uz6kSURAGNHzEizlZ5ZzL1wWYTiuhS
zVP/MN2aZ/ECyAuWS/IlV/rCX5rw/VHI4NdOZYkSJAtg1x1ox5Oyy17s1tgv
XFIjCcQ9ThCkEJJGLSy8HBkBI5ayBNadO6Cv+TI2xVwgtashcDU3ON2tnemk
kwRTABA8m+czipCbLN+ML/MxJfhH/sC4H0Y8cZHtP7rUhhIarMy1TLBymTjk
kbwWuOhAC2poea5dFB1EU/O5ZAhrR2OCjobCUBBuw7Cr5+sR9zevLGL/Tl6/
N2gsRSz+VBIAQohjTkNbHLbHtsBPUcT35DJ9jjx3D4mIaekZTB9wAj22ZK9z
OuPsCvYoZd5dg2Y3Xpez8wPLFOyvT9i7EJoJlqm+gj28QCOgnNLyFqXcL7T0
pwqJztTmPy946cgf2Kk16btYSEojci1KiI+IfN4zx8pHWkqaVWzhOYA58IQQ
bPlPtgEKo3+RfM77a+gwL4pNoGBjl3WNOtE4RBPsVLMpk8sNJnUpj8EKNMCY
ukTB7YbeatA2G4knFy3R4WhVZUba+kAZFB8OnVs3ECV5bMXRDm15zdZ7EWGz
emqU/XZ43x1pjOGczDdg1gEwVtVZXDdhuwx4yx3gN0yWy3TTuPiigSFfed+I
7ucfgEtK+naSjh3bVPGJGENd5gdlyPLCFOWeOPdMMmPKG0zwl/fDSCNDAXrp
wf0enOhK+qHG1LY9kuemnRmnBtQQ+ZUxcT0TVjeAld5uwapFBRnsuALjuNww
fQXFJtxmbq007wglA9L7TDKX48Jl+C9PLt1zkyOB9bkPEc3608FbBs4IZyNI
Ou3FOwchedbbboPhnjhOObhCIQecqZlZq4PpntskFJ4y5m0C48kDbEBwvq8y
s6TQa2vd8SoWpIYj9vocRAMClOWWePfMaIKr73VAS+7g9jeZSmk32wGdJCzF
Qxfohh3UIqI+GSmZJuc1BLE6KSDKM+e8oRlu8xLMWnro6v6ov2uEc95VfBhv
t5LifrPOe1E3Rgo/8MmE8e0inUKHGB3XOsDu4WiFNBWWP5ihUYQIFis3ppDw
o0XoRTOD0MYrK+R/1hlDZZVU8VEtCsiQ2RUkoQejbub8Ta5TTjB2yPf4yNjf
WkUHkDF5rmmBEx0iKckxwJlyyKdt8Zaoh7Iq26sOYEyDO9MGtz/IKeGv+U5W
ULL0r6D36ge3akyOap4Z4OeH5KnmKdei7BaIdMqokLnwdF3w3Qnxz8dWupFD
dJrGZP5kuDnOko/5phnufdrmguwJ15YqrB5dzw8RUs5xcnu9gD8HMZKQ9+0P
1PZmUAkXB1uMKyJLjQgKfAiinCXXdjdjQeAF/8VT1TWHfHMXz4UCjTjY7YAF
9hmTL3CjVcmy6MCvt0yyIII8d16GtZ1q3ef/4mbtvoo3qn+FZLOUW8z6HE8x
38G1sAcquQLCaB8IA1pyQ1PUUro5pK2rTPXe6p7KLYqxZVxFJIyl6P0pgmub
jH8S4Vby1ObumFr3D6R5DrKUBag6c1eSB9MTq2CMkDdGBtvfci5m+lugNsUm
NrZiTwtcbeMY2qQBsnB1wnK9TSqvuIjYuXTVX94LxAtt0aEPzqacfKraY2ex
iF03+NddLfKCvOg9iybquyONoyjAtflztL7E2dmZca7yWoh+S18Hcg9cIlIr
NNq55XK90k4TRjSlYE/p5X0BBB6Xju4mS2lV4v8Skm0SGl4p7Z34wrWZRlP4
ycKdtULnlZs/mFf8wRCUWSbi7D4LhzdmOiu6Ysi5FuRoaXHnTrAZNmMlU3G4
wPxS/tKDQtrTq1IwbhAy7HKbcipZSY3fUST9HHfLxvEA+Hk1HGEKSiUDChAG
O/17a00gZFnPaRCTQshyV9d19NRgzhZVDCXTYodRtmuV1p7t7u/EOEg9OKQg
S2/gvoMQB1YOXg3zW0cR9gHY7weQ8wcIVw0gOpf9QwHDDk7lUmczCIlouzZ5
yS6Q65HmJihBaUksJXzDI1B2tf/abBxL5bloOvhjgfH16d6x4CjzOyLi9Hhz
25qBfFsfaoI6zAN82rrrzKqAFgw1Z08s4iXVAAK4cL2lb9GKztriajuIfIwJ
1FOppDSIwEqGTryOzCmjY5RapB9rAD580rWxhiZ5rJnRudljNBG6b+EiDZB3
4td8/osKxHWeNWLktQaiuNAOsBEu393V9zfIJUvXU6tytEOohi1VfDZL/lNk
lSkESvF3UkXsLq/tIytrkjXj0/O99vDbICPCMnK5RI7v0h21hTSpYc7vZKvQ
jO/gtDti/Wr9Zq9M4wYVF+uhS0s0AF0L/kTuJl+doryWjy8mEKr7qOQy42k3
3wP2hJj08D1O61UFFBWH1s+0fSLq8cFnKK4PbAngCHWPg6z3HT1j9t5OHqND
/x0d5lJRHVjNDSunXjNWZZ7Y1PeGmBeffn8K6gLEUOywNKGc0VEuDSs2Q9s0
scmUy0mNlsI/AkHrboU33lhVXeDf5ncw64JszbLR1i1D4TW7rLBiIiEUjYZf
sjVXNwRRvRbD1ZcbwDDo/tLd9dkFmV4tClZ+ayhvXuWU4UbtR51LcjXLX2iG
D/3HKOnsnTSxjsJ62JNIWMjDUCil77Hp//Kkoq862BoWXzKtSJlHT84TF60i
LU1BKjhLyoMDUk5D4AHTnzKGWt6oZh1uykNcLy72r0QdbBuPNh9jOeAiK+cQ
z7r563mfFGnyiCGupLaWprUStwxG516Ir+zVMF8G/qz3xGKElc5nJ7NRjCEY
8nCI1+jlSv0zao/DhqbaUasnA4sx91yuORYpUqKuHpO0Xa6X/fADiBXKtK/K
Emi+sdW9L8B0K55AvviIdLshjAFGXMm6wUwy6eTEITZZ2vy0vtLnRr5dul6C
QURumJM8RfaoFUQClOmmK/1rqJCvKmbQT+YlvvV/6Hli9K19p/1e5xrgdL3Q
HnGqxOURQIGHvvqwyZX1Tie6ZPkXUI3OcfTvYx9Cgi8PuEGyc4h28X3lmymP
K6Zwy7vJ+gDfZOuK1f98Y4vPNxpN4VYfMGS0p+AmbKLNkWEB6E3uN/GWBON8
CbxHpWOZWZLkhkxMdufuVZFqT/25UWjO/0DZy/KfWgOmPVsJyKczAH1WnlZb
JuD1wUQ4Af29mBebLUmUBrGcc4r2Auo3VTav2hRQrR9PsdQc79GkdJlQ8t6o
QkSr67a5hTiXjVBFOyZyazP4xLaSqsDaZIHRzsTE+73TOcUv4PCvQKGqUhv/
qyh1xmNFuIyhKcJAHZ+Tgg+xInRj2zqS4vvkoa2GCz1Yj+9yLedlBHkcJW/9
vlztT/lhAIRty+eKR94tkRfaRx1V7wLh8GN9BuhnAS854bquSXWY34figErl
mMMS7dfIcd2UN9AyWM5q1WCaIv4eDz6Iz98QfPOs0ZChyGviApXTvEoZGde0
kwisVpxMwbBxGaj3U1uZf+a7Rmi7EAPH6YBGD7iuqFgF5Kaf2sQCoNCU3H49
413xAxEkDqLiKRvk3/2F6Hfn815m9mJIR0acXgCRP10dCE6KqTlelQU8E5sY
Elhpw1oXqg7nK96Howt37UsOGBwi+Tmc3blblkAllTsfwZVUD3dUTY8Xc7UV
P5NWr02kXYKaAL/jfHbdykt/iVhidnbUyRF7hkLsl8mUDKbNugUW5TJH/9Sd
iYnx81Tlo/YyQUnwZdbNwCPjZZYx3BzoLRl/YJGtLAo2+bj8cGvjDJR52hU3
RghQn+4T1ZRSK6h8ZuugI4/Hu3yrziecDUcm5u0hVqlnAh4e9UTvuKyKEKe4
nsuX0EsbwRpouE0gaNKs1e6oGOsXRZzY1VTMGckip3AfXzkPvlo591qOpn3l
ryku7LsvNw07oJ5xK+w6Bu8EDv4M4M7ccCS07vcp+jajC8QUtEzCxaPvZmsd
4Unb6p9xXcGSfR5hWnrFVFPg8joWF9ykB+ma0PK3JnZEkJKkVd6GArBx7wVi
io2Ja/6tSJpd9js1rBlXZPZLdmfCh4bmETrqDuN4XXbGkp+GVtn3m4my1oVQ
ZwDtpXvF9HZPkr9nVGa5C8jls5HolFDVBWqKEcF46uYSh8yzFOeu1u2+eX02
HbwbTyfIptg2j55oj2S8adcOKXEmGbf1iPEJatYeSQpXW+cEKpWcJU2WIaew
GPUNLEt1iz5NrJdbSU4u3G5XVndjbFg4d4Q0DU4/Ah2Kd8y838EIP3fKQDqU
ffbKfrPlTklAs4GR5hJV213R+sPtu/8iC1zL0wr3guUpQ3FjW+LDg+ObDdnz
iAkHRlTwhoKFwwE8RmxpSzd8i3ZFRyPtm4FBdAW/EBAPJjjc692Sm53BmA9r
EqXhAZD24nNeBs+zXM4qFu8YjtthKy3/T5ph5CKjZo+ojYC6hg6qS3xS27pW
9YhpSV3hszHVAyyKhEz3RIih2cHFFhqXtwn1Srd37M3RVkE9M2Zg6XFkqu3t
f3lMJJhLTsbTWdoxuRAil4DUcvmIInK31WY9RLa4rNV36P7IaujVv5Jo0ipl
4vXdA27TsivCi5INe29sRuUxyx418VusTvxcv7WNsrRKGRsu8qeGu4Rs99QF
VHZwZFL3pxpWPD3YVwssD4MOXJnYHSArNzNjPgNVG1deltlDhDmgq2z2CnHW
mpDZ276ufs05Wf41U48j5NSz6l1kdleHt5SDhmCYu/+dGrAtMkitIurgYtJI
L8bHUT2Fy0PPaK11nyStpDDmGIIV4UOM6XWd38Vr4YpFp8mejxXbISdOd8Um
SFZWbeOnP5dNwoW9ZKcwf2/EOiFKeZD0igw4pH523jtzkDX50zUdtWMImDx1
wxdPBEouLgnO0tLXCqLCEEbQtExVB4+Q1F9/ULQjVUlbLUWoAxhIwuC7dppD
9ngmNynxbuni1JakArjA/zIHxWZt8XD151wtzxsrQiD9BiuFq8zyT5xZ1Fqb
XSGgW60VzvjxcKtEZx8RoeZzgFvgS7dydqx2IIbvZwi4PXhVrsi+mE4CzAJF
wqaeJMItl2ln/43XbcKnISdRcSX0OnkNLElzb4nnTExP25+krTaAXN1gox/3
ciyKYj0TuXPavfmwNfYuzjalIPUDjhO+cDBWWnqgDCLyxG+Q3ijt6skIAtmD
Ausx7Sv2UBcEG0iwyyhPXqqa+HH3Eloo9UasdRqsDtiPXeGEXRzVWtjQN94t
AKvMOK92AZeUTgSq//cZMIHQiMmhRCKFrK/1tAN2rmo79ujZdvoKjAFhynk6
kd7mC9CS1PKzCBcCiGO7chE5sz28nfOR4S8b08SUyL6LYMcyav1lWUbI61W0
/JwAYOrjPsTHrCrKKHvrPQDsAA+1O5oAL9Ch6TnUcsOf11Kf5OScJjFNy6xc
vcgf/bhqUV5uxicOf4ZcowPGK2V9pRIERg89eJzX12etl/xTBli7jmDj1Ut6
E1VtAjwgq0i1XmdgWoCZIzbY2fvCy1MdWnNk7kg/Erd/8Elt5OqrNVtKDN2F
4vUkh24o2yMrGcUQefCmx2Z+tYVmNUq7zGV8ddxFz3p3spgAwra3EHkzLVvZ
gMS/kVvmiX4ENNCBFfIWKF1O0w2rXyKAp4EdPuoUmhOC5v9+Lt2y/3jNxpxx
tLJ36MX78MEMur+EPCSlqdiO+Vh6RJkgwggK1xz+mr94QqfxVLxzE8nH/ktn
AbbCH2C/f4ONvYgSx5fYYZOnCWscRMScXGRkxs7VcQRTBR+be9gag2Oe2Afg
G7MdbnYF3X9iT/0EfKh9FrKnTWx+EcLtXfI7VOMseT3rjGVVNHRY1fKDuRbv
sBIzXq2jpspylsNYMV+yo2chOzjH3B9x3WxVugEfMHvORJ4MytsBLuSROao1
bAXtnKOMo5mqSJFja2zLFH1/qw4cs+uNeqsP1Obtsbyd159bxDGt5EyjKZQe
XWm2RKpi8jX0Qpc5cIhNIJxg3ktXe6aaSxw/8FV9glfiCm6wNtlkiSZR5PxP
JlIRR314wofljWBVG4+ZydWWpYeki42snvbCvcPTIVALx7miBRVE92/Ns6PE
PIbN94LE5lDstge1xYGqchDhIhaexaNPUV3gIrZ0YDoqQrgku5OE5HXbXn/9
4IzXvCSHtAcIygbkyCGiY4kcN1HeqmPltBmbz8KPZ3ASG5/RAeocDWjfOMiJ
Rc7Zsm8r25yOEme7U2IgDm8XNePP3Xp14DEzck67hppzVY21/jAFvN1K4L0Q
85SdGJLIa3cu6ik4/rMN/7Pe5FteL7rjK9WojLZyDiBqKEsGnXBOJa+k0Hwt
0oKXERXvQVaT8dgWcm3iimtsrPYdlS9/Oi0f9SvAfUyUzThAcrMn7Td+lmEw
9eyyiG/GfbNo4wTy9UNhItV6iP6XiLZ2NiN9Nrp242aZicZuYbSHeg5v3jIz
5Efu3uoaIPn2SFdn7Jyiq1/K1f8fHR1+jWGf1ntkCXbZ505MUeI0GFYALZe4
anLUYa7e2Ngja7c69nzTOBxGHTJMPnwnC65fWhDCdKrB4IO/d5QgbLDhApKI
vYP5eIn6EFH0HtLKT8z/43wolMFrDooLvmFWnCA0f8m8cSRPKWVTDJt9kHB5
VpxrCK1eIiKOUDMWm3iPyv5ZxfSabz1RGQdgGcweavw1XJkeSDNrEM0lNzRW
dxxJEWrOcRB8JRbPeKuFP7dwel441TUW+ick8lz10pVd0bY5Kl74bkOoZcyn
YSjWIKvIbknA9T9ntMQ6mSDug0ShL0vQWmIDsRXuth5gxyMOBfI1sB5B7AJr
ae/9BlWcQT+CzLr9IZsfmANl1/AWcr/m5ESrFmqMiRvpVVTYkv6T6uDNPYaG
hsOlI+URbuVcyBonAeRF4lXNk64JPVaHDM0A8lPMgxTJtvo6ko0HHHpGjHbS
7LGcF0GKYTIbH4OFuAnHQGXyl7NgUQH+2Jb6B4KUx63RScdUF8FOczprdFnm
2mQU20Js+x197s69JNXjooHkjrcIpOxiziCPik47T0v5BdbQwHyAbhHe9+9Q
Bj/l+oBQp6XDtMD+fMp7ZE+IhI3tgwH2vuE+0s/4eASRD2vYkuEHf+WrIknj
sj0GbJGSfuO2udnYLyiyWaSrpHMUGKb7aFhPM+58uyGHQ/T85QvNoYHllDcb
E6FJTvPzuNRCBAhAjkcBfY67FWrsrQTBMhO5RcDudBT99f5kHbZOd2zbxpiV
Pxt6Di6KsVnewRRIFPrsdMp6fYrscI+JGKyjIDXTOeyIboQGPUYhAxn8dp5B
Aw3rweF3HytRMbYM8CBtstAObfcUiWvwdBi7bWgZaYNoQip0eGcqh7OIN/MM
s5ylegXJdxlHkUEk27IEZaYFnze+Sl8ZJIqQEglhnGOV94UA+Z3Y5kEADz8N
iYM5a9Bg/tWD6m1152OOSdP+4KnY9tuco+RZIF6L/vO8hvFjv+EBq4zQzIK5
V6tFmjmgt3YJQy0QhdsPxFlww3kaO2tal8LkijnfUhgeP0KdokrualvboiS2
9QtvtDzSEHDUpU4+Jf9WTE7Pt/i9gQKCsagqMzyC1Ii3ia/4U59dwSM/RniI
Ut7uWJyWVCNl+mTJdkl2Kb0D3SGrzWask3KoprZilxKjZEp0UUOur798aVZS
6nI1i0IsQNSXe39v5tEEnxkBgJ+g3XiiDYjUluUdp5z+AbJK9ZSVZhcBlz8w
u+UIurAEEVq5o+g+UNaA1r4vR++tnHfluyOt23GJoC/J8gYTCLTQmUO9KtvQ
OETKWhO25Zhe3Q1J/hjka1nHbkdg8fJk2N/DhVKKal1qk6EusoWZpbUjXLEe
Ce+gcd7PfS8Y97xrU8yct8qndbrhNKnqOiTpgsy1TlYcC0P4alXOTiUyMDwq
ixmjbxuXkoJoU3z4sZ9sXBIdxd4I2h4sBGNk90kwEDDnP6NQKrKf2+TLmCW3
Vxyzu4NChJwFWbSXUUzA+y9REctEnCzOYgIJQ4xPdwUk9UpF/Ai8rovKsX3h
98zZu5tRlpuiHpIHPFDevK9M1w7BNeUaY8PDXa3JyNJXPwHMLf+4/m6P0HoD
pziHxa3k0YRWOPpBNgbHzMiCAV54BQtr+I0OhucEvUm8e7vwXxLlpBQ6PAh8
sfLn/Loarsiyb8eXyaev0jOZJa9XSCHzzlOMCYwShZ3uJMFIKbqmo+tjHe7z
nRP/1gmxYVZXGIQjXP+KTs4ZY/usfMNqNxIhWJArbGcZZ94+uNNqLRiN3S5O
6i4ccoq5VT4Vac67LEeDlLrNvwrCOazlOdEaCKdwneT5CwsU+YFoRIH6QtyF
My2E62Y6HMpPTFM9XeXH0J2B+yPY7rXqIlQ5DnHFBDrqg+dWJS/a3KJ2xA1r
/2Fi3KWMOM484YsNZmXmeuij5CVdMDluXtTDU+6YPZ8sEUhdUg/tMtRKWKHA
BnL58zT3itxthm3SCwl78uKRhEPmf2OmMErJQmztAE0RLaD6gVsr49PnaCE0
WVOj21lAc/cTalpfLIeA5Jn9BdJ94gPzuos+Ab0PLaYh+9AwjDzmkjZ6a7vL
6aWdIa6S6+xTu6hBCeQ8ARGTYdIoRYeP+HHpmYEOcwuyZ1tmFDwTM9UG06xP
/tOukxcHWyU6byA8hQEwgSDtewSj57Tl96tZlGHSDJVPL7ZfgQuLyYMgr/Zv
rDzJwXgkoj5Bg0DbS0G5NOOkwQDaOu/WFIxo0t/DS+QtelGLIscyKWLh54cq
Hx8UEt1zrfFM5+lpK5S1AsXE0RtafwA8ezdCq1XYNPUZN8JkXtSxAytZM07I
jUqXF/sBS/uUpe1ZP1FvZ9onEmtK6Qt9zfVMf3GxDrzxMm/0Wb+EdrKSNLkb
VuxddNRJ7ZdkoN804+gM+hEaOVJ2x5ECx8soB/gi8XKk03dMEege0KNclNNH
U10GKbTa7oaG+t55Z/z17+dV2XHEtaTcS8jTH84ObFXmHcxFIb5B3BSnvM9n
71E+RThhP/Vsw+F7gMnWGu6o2MSJg6OAoy0CmmzaO/oKbLjNbE4NdNkO++y9
CFmnJUtuRlzbJlTPUS5wcZiDL4UVtfAzDX8/0GqBiH1YsxYGftn4amabSrqz
cJrJxndi+e7n470o5sDfJUdP+EVspubgeI1y6ZuItlDSp40lwGjy4ZmNhKvK
cE9cpMyVySCBSszmmZSZS4oF5nvjdckeilk9q7SDXO08kiO8EGoFaWkmGEF7
GlkPOGcsSB7bpqZTRKgd6wJUXZCxN/veq/vOgKjTPPMy8w87dPeTG3jeJWIL
BO3wdkecGwZYUzPWjO1IaJNUE77jDgtIu85FLTYZuRjfGbHEw41ctNZGafp1
pQqhpa65JbUZPzSn89HJ867dDop4nVtRPV6T2+1esMx0c5huGZOOfhoYeXaZ
eDF4l0Ok7fmUhVWUH76c4dNOYUUpXj/hAfgbPPkAjY6IIsuY+/sThXcpenU2
+LIQfGx6MXS27+oDt78q5WwuI8xI70dPPbu+Xr5Wj8XbJFFQoT+xJxL9gh+m
Xxng2VEd+MPUs0wpOuxYDZBanto7W7DBHxBZqE6Q7D0VI5eZ+/moWUv+ROdU
4NKYAlm/wuOuC+2y0+JvbMm+FJbLR5C9orIR3j7kjYVdaybmbRvRlTpIYiqG
T7ByOtBdfUDCZ1REe4RB5eQutJzjkDQDIoQ1l5sNRylJbdujNUgYfvugG6JM
8LkAvImhgOrdiKCH+rFG7k4YhuWsCVfpOMh8h0UrwOBHRpNJIDipEBv7owSd
Eq9tsjuOwW/x5UQoRBJpN7re2W3Mugx1joiiZs4JsScrER0W12JvFQ1lNEvu
oiTpUWihaxY27HA0CPPOlHr3dch2ogv7V8jgUqvvHMuu3VPvZTTsz3FfJ8Ei
Clno2vMkEjwypm3omALmNTo6XInsrS51zBd+3Ewmk+loIujOqrqetIprsNTr
PIi6CIbKVesfY15hZk++WeF5gLU1R2cm3kUI4uyyUDQIUut9NvSOK6irF0i+
jgxX0ibmrs0L42wO/6Qsx0OHCN8b7jBDSDOyx+2nfWKsPSeHdEzUIdClvYiD
+kWNE0Hm1pQuSva53LpK0HOcgr9xbTnHIFFyu3zcGApJFP9lkGkFMRtTM03p
qzDZuLc0PXbCoBL+rJmL9U4hpoyLyzXVG6K29fzN1DETT0UKtgO2U+AWxBbZ
MqrDHDIUKprw/oiGx6/vhv3pppHsMcFxIFRts6r2FO3bv/EkCByOLVhmwsSE
oxtfBSFFxiS2tsRdr/VWUbSLkllR22dregkLMPo/TxV8BS0AbAhIXkBqgJnN
TJPYx51z/zBJVdLkQZhNE8vD7lP0e2oKrotRMMpRhFyVR/KqI1Y88TVftibt
3LHklqEb9elYvbWP62Kx4Plb4G+Sbh4KZ2v+rY3G7ufjR9igOFE26f0apBQg
d5DuOniqyUQwY5keKjv4xGqri6YbqIhEQ9SqRjeIT9AcOuWV0oGY9NC2jl6e
qBoGm+8FoY1NHF0+OTT7SWNjiyxwfT1SVd4WPBCcdf7hKzY5Oyai/WfDOjI5
fw/SzEsU++/ChtBIwW3KrB54bjmFtTl+jKhYBbT+7S0MeRea+xIUCvKnXNbb
tY/+ZD1/3LgtmxmagzAwAbQz4c+XocJdPvEEMRKpfnzXPkXaNZ+xXEXdUKvJ
5YUiwUhQi2s4aTJDZ2oP61l+0kYYeF6QDiHYodTp6JwAPwXi31AkMdVn42dY
q7xxnCp0MsbBUMzDVyTJBweIOR9H4qjhVM9cMaX9lag5kD/vUkhbToAl08tb
/LYkt+AkpaD2WRoSNkJM2GPJxpfXpDwfthit+U4SilEvebnRragPr6NI8pTg
VvduUo1F28enhnEiADIm7kWneX/C82mCQfCeMpQvmyV9OWAFY8F2iycpS5Rz
aWRZChgw5qyl5Gt5P/cqEvlsdzlFS2I8ywsIVKc/lT7Qi/bgybE9YjB8fPGp
k391mkg9XbkPCK7G9xUuJZCXbDEZEntJpYTizzQCRru7xUkAMcW1IzVx2Bec
tWFL+zumaWDnXjBBkgFkJ1Msb16+bu7DcgwCjFgukqBV/Nf3Hu5SF2tlWQz4
UXRGbzAR5fHHJAPOOMul3QcIpvhYuf/UceQDdHqTHYrjAvKrPsqd5f1yQTtw
HZ/MJM4sfcnCCIiyi5rMGmwmYsL8eT/miVAVcBe0zwAD1xKsNGDa6SXr7lS1
2AHhGPF/8nVGSHqnK9vGylGhZDbyd/S8oFcxk4/g5IlWPiUqtIfL6ZWU5Wmo
++VQAuTBVQUn8BfmenHsPHZMcH8X2v9bxHVT8A0XdswXPQwLKTUvx7VWBPEA
RtzZ0tAtCuskzYAU19ZdmWACuTXt/gizn6OwAwn3Sv7MEgat/W929VWfAfQb
2pMrVX4WCy4EEWi+KhSEsFFoZhLjVpjQUMkF5+ZUrlY1Xzt0FpGhM+yg6baM
x+ltW9Actqe7plwC//3IyPwib/8GIPqjyWtJCJc5AvzGddrF16lFAJ6fFsFC
j4cO/iPM3c5YjY5f+CyB1va+KVJ7q1rmfLKpWPus7V0KZKnOFjhvBFditkCg
EYgg9UJGNB3X+zQx5vVhpxMZ4jCp+5S0nd4gJ72ECaxaX3hLNv2DwHjNDwtw
Q8ZRIX3rS8dztOGQF9841eOh+PXnflUZf7rSXAbrX+AkYVgPeMRYfpDBqKPK
vS4dURZBfyvoJl1A6rRfYy2YsxZSNSF12p/OQL1w4JtAA+T8h+77Azs9bzfW
tSrfsOBPHFF9mgFZKllnjSlCNCK+FXMflw/9qKayATVbrYq5d2Xv6xSTBeNN
N7TmaK+cp5GBdh54jI51DTX2VobW0Ksa8DFWq/ncfEr8IogTaDtRv3KPPfod
8DWQMrAFEbPIK3WCcCNkDI6nxCv86SGph9Pf1dXwCpbZAZRIdX9+DOg+UxG3
pPWonn+AnyAxAKkWxVPCQeErl2xK7JMoYNuI4C+eiqBmhbWe04E72smUatfA
PaAzTItJsG/M3AkIBtyZKpjntgSsIqBJFfTE2D/QNRv62INWTewEan3GfVf5
KWDa6576yWyLeZNA1hmyEMVaokplQ7ag7VA7lP5D/M0bs6zQmVTRu/fp5snq
nPwB1jA/i+tEJasFeTg+Fcfzom/iLKpDwlAbJuSLrShG5yzEjaXjtXTpB+/h
g1Zbm6lJIyb6PrRVQnO6boCqZbCCR0Ky81DNTyxu/hB0uBnMPonLz7qq3TQ0
cMeFqqaxxCd/NeP/o9IIe45MdKXgXfjPGlvuSPPI7QQtOn5ZG+G2pgHnTdio
tE575hrZ8lQUpA7GNN4NC6T8CGhGfKDl63Im2G8lHW8XAqEMi35u6wT2FG+N
An8sJR4z1j9oIk7jKNJ/aew+ecfikA37MUGR9AxOxGxcFSfnizYkAqGGXZSX
/he2gG6ZuTMkNfKmYiYU8TfEaKqul2JSMpBAbDv85Ca+pDoRFnKij9be+y2E
0w1kbHWGR88/XYuXDjOF6Lwd9OENUjEsm2rQBkBVN3wsJQd5aWmC3VSM409W
pREBeNAQQtzACI9BHeP0NUFiOtwvZuqeCFz3Apm7QuorrxBuaQD4WXMjLA7D
yb1U021azuzFZG3/xnuK2UPVnQdvy67JZpfX4bgItncaKX3ZYOwr1v81ntB+
OvaPXRKDkCUu6J6FMIEsfIpRG9hpq717GxK+bzr42w20xN/sPlWSMO82v/c3
Fd/RTbozh2hqx9oF49Dnn3MpuTeI3k7iJqk63XJ2qmMm4KMTGugOn0SkBAlQ
r0gnq4rZg+SQLo2WGrdabvac6yNQTUWD/Xs6wiFiWTyA3oD592RYZUy2pf29
RYVylLimpRiU/VQYST4ouywkV5Css2nd6ruFW1opgqt+hkmSCfW9/RezJZ90
oyMgfHh1un01keK0wprFrSf5Mg5FF08s9qja0/a4gszM4BQv3kcn9BOExGj7
hAO5HLn1r5cMt4rGE+vszKpFb8F2Ko3e9MhV2NI+5MBopW37a6xEmvpPYeHI
+3lu6ZMJn0a4NwcUG6unqXv/SMIIk0rW3LNxC4FvBPoLj0z9SRJLECw0zUJ2
mT/EIxIjS7HcmhihU2qtRLt1GuuhF4oEgeJQXqwj4jXniyBLkrR2QI1NKbqG
hjPn7n5FeY6cTStYfYuM4dg5mw3cNByUJGR3xniXd+Si4oQqw4XVV3WSmSA/
mhaKhptg8w1huYDeuL2E7BUrn9T3FuIipd65j/j9YTUVrqn1KBDqUiC2Zb4e
6HcWfDmjG3oPlAwzNHPrjjIuwi0XYo5IOtIq7lj1FWY/Gv58s8p2SOhBAcpT
jE2mvOFybWP4TI0kcq3IncbtDdrV/pDHJtPtNkOSRBSXxjh8BDxEEw3DvnoO
ikGYlsBRAmIrB5KTAKKbiHIh7VXupdFh5eBlryxYmur54Z1efzWq9Anw2xpj
UT4WiKyDo+lsH8FBFBIZyB/L6dMVfbbIzMC+WDmMcd5oFXYljA3nutqjzVXZ
NrhUTq5zzAIRRZvOsPIxu5zBFvAhk/9piB+itXqTOAdG4TyxEizuaAZrf11A
bgnEu1nL7DbpuwPhSWZAQ1swv0vWuZ/ZpZrUvGiPK2DsNDugicARoNX9Yr9l
EvwRNI/6nwZB8OtBWRN3eFrOiX+YqrwUpCqhQ9SPkiEZFl58WkxDY7/PEZ79
N/qvxUDkPg5gHhaqjlYJJGgQzz/1MDtYeoq8QHZto1tu0wdxU3jGGDzKX2F5
V8SAZ8lkYmShJ6x5CuN8/+QEA0u9lm8+Pye6JRCx/pCUHlvwTu0Vm/RfxSSx
eXN9GF+8a0h2IXgxGj/7AwXQzeHyTXCV8Klde/VAqd8ZYTtMLtBc8ozy6Ayp
GlttuyWuVvTvNg+xcFh/DvPRIdL2J2uR8kMvPRydzcGX34extiVO5kh9JQg6
j/B4aw+c+vyhivmBeBKkp+LAE+45XUDghZbT7RUfCEFQxOX4hIAYYTmD9VqT
QGcc/4bfV2hiJ1q3ijwCPofNSf4WyJA6MAQqhRdz4FO6MhpiAfFNAkSazMQU
HLJrq3kC1qvVEq2VcAMgg7A0381K8tRT3j+gBjQ73+UopezJrviNcN0MzbBW
SAdRi8LYp1Wbi80uoCyIw4uoX/w98y24RXYgSCjkT4qY4nXf2lKcSKWezW3V
vds27KRBJaUaYv/xa2M5HN+1dA+84dEoKfeBQ4JsrbvLYDL8zNx1kZZdWpee
pZnNTtlAX2P/7zkNDHLX7g1czaANcS1ZMgFgypcPLqdWan9qXm0vJ62OOc8k
cwTFHMcTZuHvlcisFAfq1DmqJnRQHa44seMrjo27Hgg8EE28vxO75dm/JHA/
t2QQRWc6/+tinz4M0Rcyn9FYkqYRjtlm8b/YVRu7ITI9Yc/oMmHEof1+yUOt
SgUJfYCmMA0OAjCndLR+yUGoC9PPu/b0a+VbRlKDMHnNHDAgJn90XYxGmilK
BZQWxo2Ozo+dtCtii3F2xumpGKvcyfA5nhhRDZ6keehxlpBRodEbz8f4iI+T
mK4X0rOm93BWyNKFSxf3JWomdwPsEMGFUSGNqCTk58wp8mtF2k9XtJR1p0ml
dliAP0rtiP4ZZhE02IQJGep+qbPUa+jB0HSHtr/sH0whoH9ZGG5Wl/UgAVMz
eLybz0pgTOYzTMk5mkQ7uD5M/3n00pwMNMesJumz5RIc4vAGT74bRcs/Corq
QiTW3DbqsvfDYp8Kte4taikZLRBb1KqDB/bcNrZaTFMvCURDvecmt1qyEaOa
4dUFgW1Ujk0UhknPA6PvFY/AseeDKbngkN2NjnO+LKADMytVU3tUqqwhWvDy
uX4r5NG4IZy2eQWTkonHdiqgVKiKT7mkD26fK/YoAFkZXSmkzhWN18ZjSwXt
yMvWAIuzdQbQbvMUp+2EOgGZ04ge0R1UUUi8PE+g+rT7n4g3WDDG3DWC9qoW
cW7chwmYU1tQErvSqZknWQxJVcq8CIRm1S2jfuWyIl4z9Fu2vBXk1EVwZTg5
cSg1oEddlRjnkvtRN5tetAk4oWZoSA5m44ENweSopokZkgVDTureBCxLqJjF
dpPuqLx2xgZgsO7GcXL6aC3G3+J+s5fy6uYLHLc0SUt6wlPXH7jNEGGjuYuU
8S4t5GIBwfoyWz3UaXcxmz6VEHdBBSis2b4GWIATqrKlWNiCm0bSogVuJE04
EPtBnjSw8k3bcE9lwOLH3mS3OY5S7MzPbT+lvce7OWwunj0fJgCz6+Na9HT8
Wl9FZfb4MSEENiWaIQyxFWA1zDyIZqjWeHmWHwTPi9wD+rZlqpCd9pnIFh4U
eAbojt9nkoijP++GqqSSHboTrc/XTkAulEyswdsw1DyANgl8BVIS7dOwmW2k
NqEnPROfSkLH7uFKaJ9SiAt59QCcsxtxN7hQC8a+1bMPeajiLpEL1Q/ZeYzS
YDoNDr8zjqF4ZNC4GKu3rXDBzLXyqL1cvCVxAyY1uubxttUDNhlGJrqPqPXE
39r4QquyWNuDCbGq/45LO45WF0pegNIweoEnYzbhERCsMpKgYVqgDOHpAaSf
oiDy3JV4ngGNmxz+jzu8MU0F9usHIm5Nqc6eFNGg0+ouxQWkGXJ/WPX+P/2m
6KExMsYTDel0P2He4tSNSiRzjE3Ax1AFNMaaX/+owpPxgRJzhIpmOsiWf2RE
oCBgEUbZ/kIm90aJOVb5x/h4jK1RkjZHY1PSkksyhkjYDTmQJ2YPw1ou4Y6G
Lu9stCFzUu/YJdlSTi2LRkpuHV/8zHkh4QwahTmuVUzlib9bBc6EIpIWIX+y
tw58rw5N0c3l702twguugjQ97MWv0SbveRb8kX+XnXM0mS0KPlIRxo5ndDjC
SfhhZsS3ynK259YFG0y1XUHkK7vx0FDpRGoAMX7a/XbkNaVGagVOf+zpBBiO
nTOpKKacQfmqC+LhIHg7+JAQC1VZpvzH8Ymp62YrGCVd5XeTRWQODdz8zMEc
LvIdV9JQKoNJ7IhfJCDyWmznKoMmEvyNCMgyvEtNb9dwIH2N2wUqoEOBGn30
MIrGaZJ4+jOj5Emi668K5dBs7NUPSdzaaoXMyM0WT22gkAkIMSqHx3EjLYbT
RJ2qdBUWjbo/M2edG8sGiIXw96yP5c3tqtgtDlyENjjhfDAsQeL+rwgtCdel
C4OjfgFrpnvAH/DiUCN1vPnwJqggsuWbUxjvG/WZfWSvelgSnU9x15evvm3M
xQOULL/1cLk7J03L8ZiDr3J/5SYKh+PggjS+OuS2RnzqXxSNwM/tpeGBxAKy
kI5B8UGuPW2crDWsMJwklFpSOriwXnLItM/HhxQwVRya4U2o/7qRLKtmVvPw
dsQ52vWIQ9VIrb8inJUudNlEYrqajwmmi0GwxP6XmaM+N6txVTXsNtCYANM9
5UoAGT+e89jREiLcLYZ0nkS0v9/lOY/MpvkkWd5T7tnpYIocrgVEPnUjC17V
AdTqgq7BQsy4WaBNdFAR4bCN+21NJy/Twp9rNURSgzhuf00IH2NyylgbZbOr
SecqxIouuHGUBpekPzbnazpzmKrUD50k6obRW05CuArCMSKoKH3CgxuMISjd
/bC5Vo1Z/5uZt6hkFvfWCCb+UGKFFamWGkVVaBAAoWI6t28WVKo2ThfXTFo1
HIdZdmEGekCgPMwfJmPrvVoNpCS5LTJ1uLQV5lXlhICsBcbE0BRhOZYi14Su
m2c1CpSBRpP7GjeHr6qu7kNw99WzKNhMwqRG+5H5wkdtPOcxmoFOyVl2qtIo
rSy46MVZb6euL3fUvsd1L345ZGUA8wro0f7sOjQLPAKRsFYN4Lk47Id/Zen2
fRPoZjP3WgUDiuyMAZ5q89hsXICfbMkkjwrcdeoaz2nV/cGW05U6QmmxZexr
LdMJUadNWiLji8eFm4Ev9hmgSrEY47Di9E7vuFYSZpriOnFxthD7vubWidEG
Od/VpBhUDZhuI7wRIucVctohDlu1d/7eaH4+FbgnixiA0IaRTKpKzrbJbwUz
50Ymjev7+xtdx1GLaJWd0cgm9X4OZrp3ZbSC8AGEix/EnFfDbkj/e/HluwhI
xmB5fWQuwr/UWf+sCPLdu2vKU1dWSSc2U37cmNCp8HYjlc8J32nCP0jfDHQm
cq/kzD5GP1EbTLISMsLYCR4YDi/U65FekA+IWOF0PIplFskL2zECdFxM0ZmR
ZgiCLNkdijEYIsx0+/yJur4qScmn5i742ce52yZQCaAUIlhdxlQSVjJPUjh7
FXxA3ghkNsBTgWs312Ar2DyXMiaRyd8WhWWMhfzVjGRxi3xXR9gh3wFTOg6P
jktOOGJjfGgvXsBgbbzRXvPMlK0V7F6kClgvRAAysbndKazs2iFyksvXTr1+
8coN0dI8MV/Zq5DTll5v/+oyfyqqMSIAoJ/4NjT+6dkhfwLhG/HxjCzoleMJ
sGgVkTD3aSNc/Vf97emdjDlzGTlbtXR9stDzgfROszlzxFzUGVko1gIeIseT
L9tEF3VoXsDTPCGhxNy60uODuhy2XSn1LAV826SJjkOfY3DKQ3ivrgw/vxnY
I4ZuR1wS4MHfLvl5DwUqwik0PZkNXuQhdMIsI5LYGJXcC22LN75YlccKc5GJ
KQF8QeK4a61222s/oU0WLjnXOD/Cc37MkJiJrvtAunop5qIKkhazXwR9EaCt
6tCzwB7jqhZQx1Vew2jYrl4TGrNbH/rgHlMH+15OTD1ZjB/Ss+OIZhGmK868
EOBIZrsyoBk11qySgN1D8rDEyWnMSd6+ZIphUxvRLnYsxoulBpRHzx9a35Xa
sJFZ7dEQZVMvxWgo8kcTPanQUEw3/ZdO1V9JHR0KJw/09s+2i2lqXg/tDPOB
Lp07yU6ozbK+mgyOBm0f5S0dFnzh5iVUNiQ71WIFO2RPlGIlOjc9KKbGQqu5
qVncyc5cQaseQRbnmkh6Gxq9pcYuTTggAnCQQGYKeP3V7uzNvi0Ofnz0Muil
QTYCRHAT6YlOpYBT0/Ezx7zFNruv+0fMpN4C40DmSs4eFd9l2CUvgq76V0+U
sCFBz1cm5JqfpvjKYjlIj47OrE1Ci49XDm3xq1ENmfq7dUd7XJWhBoP5GWLM
yFb6TM9WY/165sHYDp8KNCEu4ybh0fDxFOdOAbJYpbIC2JYW0SYTFSnK1i4o
QXTnLAXXr9JvLZH0HzlljGJgReE4R1sGRMK/Ix/orPYxtHH+OkOTcMx1GTXB
P09+G2rFac89ppcZ+jey+RiAOEesOBCcu1rANZUDN4pfHr1E0dYEfqwZHPpm
TPbxLHktsLFTe5GNgX8PoQsZr21SEhuhguyr+tx1b8U+6f9IMgalJGBZSzUI
IhpE6FPJUWjKrYwXsHDOgY3IyJiEOegP9X3qeHtJCZlviUvlVru7STJEgD0S
M06a2y9k+Gcv2TCOjTAGYeVkDhnBfw90BPdAjUNY4c2zy7gUTxn98sDAJPsf
7eeIkgPC8ydRqSavxQZkAUZX9cLjJwCzEt0z5Lv3kvfgSSR3sNkxDtq+Frsa
GwQHNELpvcF6h/42s2B6cCnQUjGPKv2SkNZHi7WAdyxuBFfxNPLjyX1W1Iw0
mGaDYEXwtNVT7yNP7Nzvwm1mq1bGC02cY6KQQUZtRgJciaIY/Jup6jIih/ZJ
MskJ0viU9JerH5lpuGdLq8T6Z5GGacgtauAOy2Mrv2eCkcBEka8BLCKMchwN
k0BN676NESZKYG8vEyf3XZmvxhHf9JIJWj8B+Q4m/nECW0gGB0skQ1Zj760m
MnYw+lvYrfPPEryCaMrREFCGcQEDpQgzBYAyeySopjggBIx1mhRWrrpvIwRA
EyPwQ1jysUDHh1989LTH/oy1xhFFOgUGKo+LMnJxVx1HIoZHtNqNapeyOxiZ
oA0saph+cwdOnXz7Qz8mGTbdehBQo1vodZvN/8AT5OKAbFLDIuJzxNX8NEMH
p+Xc2zyG/OIEeD/HOlXAUd4SgypL1H6netIvyMc2+2dors19AeSV4qCuqRHY
tSbGJwmSueegUNyb0WGpVCsTt1mBuobI9tLbw4Um6tdodzT1n87pfFdLFfwi
IB+JYxMW3ao3ClEnPRbSutt9KgtH6kkdxT0MSwYCHKn/fYUPZw/EBXoCdHXo
HqLUP+vePRhTwMG39DXh3QODOMemaAZ28b0kVRfaPhgFUWkzDkhjsHuQvmh/
A3+AUiIf6d7/I0MTxu4WsiLn0h4rD5z3fXG61aZh9EUTfpd4zh/8ihZJPRxP
1+yUuk6xqctfIYkz5qZrrNQHj5Oz8HyHNv8L8petmBKaV8MqwJRCq1WacNhd
R1iHFPstF+wP5JbUUIlXxKrImq3kzBeHy7fFUuxTukVpCXa8nxFlf4HBKhpD
77qhWsg2sBibM1Or9Xc5aRyRHBiLxH5WLdj66NvBbYioCZFo88FCO79qYKGL
KQM0MeaGoyqD1sDv+p9v2mcusPg+llwA19Cm5LMk1ioZT5luERrqPVox7xbg
O9LTGAajhkpgKXXrCAyD1YnxKYmUbfSDkXrFkPfK4swjQpiFKKEQdqeybjSN
Hd1rc6+XyqId57b+3JPdBquIepNBa2n1I2ZNBhltYo/fsdNTR2uHiZuPugXz
leGocTzmuGabo+QnUIeGf1JhwaeHT7OXNJKW3EGR7RXYs+2kCxu/BTnFpUD1
o0HZlNGfRMafQOSrq0907rUg+bVhQykejpcTvldDpvdC/2usckX9iClaKsNX
Z2hBIdtvL+Sl2p+Dx9vostrDRBaHPs+oOnAHIe5HtGqy2hO2/i/ltx2jCvOP
cuTMsM5pwyHz+QMBGXhBaKIw79Jm+Ssbd6NIDxf4Tb8f3QyUoGxdmBGnhV21
7rhiPMz2wjJwEvw2Y/iOhgnvG58pu53jnMQbm8nGrpETsq9AR1CSgYpsbmcB
PNSdvarYEuO5xnC9FEYWiUghv/F8N8M1pDZTrkix/l7VZuNxnUsUhG/Xkjwn
SlcOv9pWR4324yjYK30OsxjpUtNo5jf3eQ7Wn19AKxE4jPuc6ahlyTzo5/lx
sDmxR+prIBRA979hI9e0aqtqFXl8D68pw9FsS4jkH+7gJU+t0gbfkju/9wLi
1x0wZXVHaLqGGJUdfBc1JxNujeLXGFZIvn8kFJzq4b6GZWtUaCnCy5aPdQmy
qAIR6uMcLTURsvNeATO5TsU7soYqBbZRzZwva5ohURH945LxnK9Kui0JPhgc
u3c0ddk6UQ9xtW/GEpW1AOOizAZcO5ZGjwKqpPpIU0oanurnL28M9199MNVc
QcUJt2UfMksJdgXiITuTwcjLE0KebbIZigVku3zH9S+mRsnmP19euiIcwh/L
v6nxaZdOHKDwCx/97j8OsoSeiFhQBc7N83Yho6/Sv0cu3uKs1yE6JucpYQFf
5Ef3BHlqx0ayOB4y+3MddFjTouo1aSw+jGBqsQE6KdkVCf3LXPLgKy6PhL3Z
ODTcd4TS6b/1lNEtqv3fRgABjF2Xh3/2RIKv73HwvDmtVI1GgxkOHsE6DwfH
+KAsN1pL9EE2iZhvo6xZrzHXebX5fC05aCHFQ5fCxua9Mt32JX5n+VDSXzDH
+Ofv1Sm10FaV6pacR/PplrGKFgvzt7XMEYcB7g1wUM0XYCvPm5QfMddWLoQ9
PibcoF66+fKNiS4xLi1ODSeuTorRsoRElNQbFdrLbUG5hhyFT1iQCQK3hk7H
umQTNGm5fFDCsmui6tNntkz1n3eValXjMWcEys8BtLTRwBv41Bx9OkFEdhC9
P3yVSVVJPonv3lH6nEtItvIPciR2PMywTDvM5HDtp+zXYrOGyaHv/qlHl2gp
38VeOAzViteuOvI757bfFJ3ie9UjT7Zo5U4MtorieDuz3BVyx6h6BhR80hYh
zhw8WhJMHu9DZjVudeA3uCXYaYV9nQEi7Nvt1mFdUva710E6x5CLUTS3FR2Z
pGikDydfPHX7Sww7++i9d924ggt8yqFxngdthOLMNAIHFu81BnF6w9J2KPLJ
ces2S6ABtjviD9MmNRXU28dpcr/gX++wCtCCMgbOkC3SJcuVVpN4CI+gBLuJ
5QUmT2K4NUAYTjYpNwURzoysC7CRnDdKmfsPahbxIYQxe32ja+tihWrcIXrm
e1P1UPysS7bXBmy1eXUQkcWs05m/q11HmiaBElojbv99/t3LlzqMjsulzQKk
BWTG2F7OV15tznznrQ1uyJhqRWRxkx1FKBTe9iSA+eLohB8pWfR7Q4kPFNvy
KlBNQCdzUYM5WI8te9Zf124FvxpJoWcq2zE3sWfKAoJOaS25gd87Ke6jegB1
HjfsHhlKL8xm0Ru/afq725iY4YqZDxFUpyudMHCERH3jn89hzSG0DtP8ubpo
efGxaS1wgWPfoJ1bm7GfiakMXWKWhvnID0YZQrlB2NjE5u2rV64Ma4vKOhgM
zscQvA5gabVxX2YOA2nJkbxPi0D42n9COS7Plb49+LD4AskSc6DJkHCaW1Y6
RGaCg74Dkbb+iZbf9q6HlUT7OAuhj6pGrwVoYoFIz+0+jeM4BNDeYyNwqaYp
QtHBzBxwJKZ/ccJ9E2IHQjLrcEXhRsaT6p7mxGwGR60Q6+oZ9w3/Nj6qGXV7
pf2ehIbq6Tvtt/apVZFR36TJa5UAxhnMt9ssqlzo4RJUNL1mZqVP+DhHNcaW
/hNCoc3fiN/fVdNTIktniyhdSoIY7drpHfQLycZyOEgvbNJTh7C1aNGR7f2Z
RgDPQzGry99THC1fzHiMvt3KyxxCCPkVG+DwY4G2NwcE7tLbClWrVGmteGwJ
m8VZ4GU8+Q0mPR/jjVAys5/QaXXeEeXuLFTSIn6ETw/9+bptNmJAj4x+foYY
JZ3h1BP1h3b+yGy4B2CDbzGvAym5GW7tm3gKMof+uKMRKlhKyI2XhrYk8fAs
NVbgOwIFbWoJqd4/dC3Dew1bjYNIpYVaIkjm4je3T+Q7luoKYfIck8vaEt7/
VIMEw4BaTGfKfQxq8kBFEkr5GGSMKhwKFCO8CK2QGpavz8N8872K6gtemYZr
kGoDWP6l8F7c4OvQfFxXt+8pkYSBqOBArtdx+jemJSmBxnWw/gGbYri1SW/g
SP5XGRNNuJF4snbERBfFET7wNNdoxTdpFtiOfC5T7nNEMeB4rmKbkwLhu88R
K7cOH/s4j5GRXCyHG8MtNxps67DYmjgBi5xbjCBocAnGdLejetPVVKLXaN8m
VH+tkZjAgnBPDO73upYyT+KzcQeGlPBmRCQaoGLiV94G8uKxwIr7gb7EQGR9
7Dcr0s0e7oxJhKjGiOp5XfdzUdKVeqGww+Bq4JV5BZdFOJhE4c0YjR7+KpsG
C8/1ZW05TwKiR307DMy1+YRXhVm49g9II3KxLmsJU/e7mySi3mbAjh+Rh0B0
Adib9ogWc8QTRZZPFr4UAXRurL2yhpWstsebur7LcUKAoWrTNyGNqhFRjFGL
ih1RA2Z29o2dKwPO+lunEgovjhal+M7B28tDhPPCLdq1ynl3mbKx7aOhlhXm
D0LnSHa5zRoJ2wmyK3gp3pIkAWiSmlo499LNXIMts8mHaZilq8z/OydxInRh
LmU/06vk9aPqcVF6NT+q8JI241nl38jYyLawjzm31NFDFwR2CAGqlKbwfgcT
0y0S/+YTfy4Iee0taNNghRyANekSDVX2oYtVOoAz2+1BIl/kK4+2kHVxVPJh
Qv5Xzn/43XICxekL1t6cqmfx1J3xMaZ3KsUYqazFlsqTW0BbGLuRrcDvGu5e
sZjgNFF4KE5WXO8/WBBi9nh+GIZEEKqpj+SMNTW7BNeYpkb9YLHqAHCJjdm7
e6/nI5BsH2K4qfk4igFHtz7HXIMDDA+1JOIBkfcKdED3UVVpQErdw5VJIvSy
cyqebhiJARFzskdX6GXZX/6qfzAL5kW25lCe8qlMb+nFeT+M4+LXYeKx9GX7
j6yASVQbh6J2wYcQnZdOZ+IjgqoFC8lCwrAzzrZSEPx9t12DxQTTYSGZwtfF
xPhesXR30p4rbQL+xjRtHaRqjvjT0E2fKjpX+J+uqzcVDXVF9+nwZW3F/C09
XaKyNQhNo0TLjfbeo0EdzBVxgY83oKNO+KEJqlvsBrNf7hcmZnVHkzJTk4xv
2N1QOfPO4CNsdMQ0p+twKGFx3dNsetIifW78zlrnw27UTRKwejvfcY8tzRxg
/o/GfkBTUOQ8hgZQ1lF/I7mYea5uueJQsYSgwBCNEDAclEZf1hqLaapTdSvs
SRM8CMy+bUJRlM20KFLX4uUzQzqEx6uu6Z69RoTt8M++fr35AjeaSYa0qRl1
gMhiXS0M3N/3Me7oUKve5Ck6rrjiWn0vDCpUgUX4vMC/NtdZxdE0lFsQorWp
7gKgnuelbvhE2cL7Gtrm+HL1qcmbVwJuN+PbR4cBqcE0QQLxLUCr/41bVssz
690yXnck/zqqMw8DSKBxybxUuodHO+4KTNa3XpGy13Fo+DYXclWceFeQfKdp
AgcD37sUykkmhRyWDdnMReBuZArVxHKWrvJypyBlxl/2yW4eR865AwlvlE1t
L+VwIclLB/JpfF//4pfuUPhMnQ2+TaWUO4AgV0XL6ppf4FshU55yGiXma2Mp
TKgFVWgS/JsWfCzK13Hlw74b5T5ij0Iq4l0boweMK7NmY59xwAZ5bT8vdUzg
2MTaHS7tjb2rfUbJNlKT9LdjmKZiTwLCtfXV6TlK2WG5zDie4iMOCM0mn/9i
+AjDVeStDwnKw8Ny5sEHcNDZaNYzm5xXYl6+RqodAEib3WGKo4gUKPUV2Jmy
9BNgZbu+sjn6gmUiw2NfXZgZjYXbsJnGJfpNEleWVJ846ZyRgLns9RN8eePe
f183uTVJAwVK5YDoq1cROpZhodQzST2xjzIwxQwJyyaaV6DFpgtC1wArHNFc
oH0MdU7hsPMGh7vctp5QItIZ5lzWS0NETkVahntFJDQipAcW0qAHIn7A3Xv/
WYGmeBHrktkXDGmBeE4qfSzRQpwdVLhzYJSPmECIjeZ2cGiIQuvdGbTVuBAa
mZPI1h+agM3Gtm+Ua5WdilIrClwe2nA2cnpKtP2+OGr/VxFpnTM3JSAwpoJu
DIWhX2iPL6Cuy9LBY4So0BXlSfHzzCBSoNhpWx1+VA3FHZso6EGSQM6mojk2
fqrLwXe74EJx5cnYoOe5ccZeUebfEHUjPt1cHR1dul0NFoJC59OcCqUDLivG
wW8C5G1AaDmU4rQkQKWEuRIOAEUfbXUquVJQSGsCWlG9YW8jt502YRt7gjnS
9G/E8JRkWQXJJz/g2phj6W7ua92z0zYcvdE0NsED4I1CApVoI8p5/SlCETZK
clhjWpuxkTCuePeEgANAN1Rr3JlaD/pJjTG4yme6OCY4oQyj0HX7odd2ni7E
i8rNl8XBf7H1qEad0/W1Nm6l8sM7lvEwiVKztcsqUQPEQbT07FP7GKCVsr4w
7mupmpaWjSjmiZjv6tfx6LCGghlWFHUNR6rBdFN0XxaGOuZqEum1TQ2E4daZ
+wxRHL3eKGUZ4VpZlehsnxZH9H6wAgTCCBbi8Vu0AiQuHy4oj4Cl1H2rOJCK
QiZImE3V8ZP0ZJKoA7yAj1yu1TAzeRVOUyz8AFa57Jv1CciW3qh00CZb5zWA
1RQYB5pNoc+S1IoPg3X2iwVwnMbR65I3nHaOHekp17wItyTdbHR3j7JIIK4N
GegRfSEngrdM4A3/YU6UXiQEXncguZIyu8zZjzBKKfYH1x3cLW3Q5k/VO76U
6B19cjUHE4KxZ+6MCh+rlnJyifVyJoZraLNadBaG+koHtx+7fE3BlxPEgZFt
H7gP5zXQwudWAZhKrWZDzaxSFd7lFcs+7hfkmJnKxRQntVdRDQoMqHy2Jwl6
AFI2ghkgs0fKahBkBWZCoLLDoTPAPJARNzb7Yc2S24gqJRFLjrxXPTP6Ikut
yy7Rgj4HWs5xXeh3R3Uv4xAgbM/wr5iUZfbD54NtszDaojvtC7e8ecCqi2sY
7RwIC6CiI+TJ4lZxvnutJDF5732drc+uZUg7CrKyNVZvPq1Eu1JmvvLHE+7l
6XtlPmmWf7U0mj8ejJc3hfh/3RbXKslTtohUh11ClGXmBttwCpYpNT5qxWQp
r0EfDxQau7f6CH9dUO8ZQQHXQUYqzDmESal5X8INhJfq2kvVjvm1aJb/gRoX
HPziUR0zUdrWAoSVwc6FUA/0bR3UB4EP1IaiabT412ufNnvFsTvYgcA3JBI3
jXmCv/p3ScBg9Bxrpx3gwl+qiIFs0GVIY65IO9ZXwevI9vvH/+/aUJlNUQTr
pY2zzJnpqKkoDtALcBdlj9gg0VBSxAnsOWQZpfIKf9g3JLsUoBJSllsW3/lM
KDIm026wzpLU+G6A8JX2Xu8YrySPQQAitEBg1e3lCjiji9fsOVo3l7yI50Ia
mjnozo4kNSoisglJHqoDiVgHxtgtxnBHQgFoscPaQBLJE+h6i+ga5ctCSh1I
bOzmcsncNPc39mQ51hoWv3KdSoIxJNJidpBp0BwOO41QQTDro+DQQsz16+MK
txyeKg3ZWLB5TLmcXYLV5k3qYQ8JBq4RGsIMi/dxoJlC3uUfFy4P1BGYGTgc
xOYy1Wpb4LXhPT97+FiSmpEbku7mLfgDPVtaBYsKA8JfJaGyWks44pl7EYc9
P0qmbf8DzjTppWzn5vcRHrxYrSfopMp9dYMudtHxYx7tX2VSMyfPVAoqS0fc
cGcay+s809HOmpu/nBWPwra6uLOJXwtzIhDbN3Al3UOzV59JxdiNkv5i95vZ
LJOqmbS2AQU+6UpY1Bik7vyJ0U/HfTIdUt/copW1oxyyBc6ke2mQONhadweu
zAClWU+FzTUYAhUdVODHY/g+AdRsXa6w9T04hOK1Mh0CeLMM8y5V0JWDQk8N
zZ/+JMbs8sasHhFZxQy7qAlgJQQcX1M8703zluA3YflpR5dKepzrRgDu5DkY
e/zgqAQLt/IF22w/3YrWTuSTIaM7OZL+9+2YHxDPLfV9NWeskSIBNv3S//Rb
2dWzHNCozV1+Le7ITyTNqthCJx8H2E9crq+A+0XQz7MkfSwi3HUbK4XEjTDm
0+CsqoXceR69IW1UdcMlovgVx1G06QAalPBdsF+RRuUMjRXIgyZ/RZO/pX6g
ahqVTPP19CFPvNDJZgW7tZoE/3VY+ZH3orx05e4xdnSDHhy/s3sU9luABj9f
eSbBwyW4KuGOmEADYLSJbJ5wKl3vka6bUMsvab7UzCmvQepfaOzpOhY6uZsk
cn6pw2XGSRGwsbGijmxial//wjNncXcn4r3Zzffd4HGqTiqA7OlcXC2TWLpt
A15jVt2Y6TrLRk5RnSr55+vSDvjrVXI/9c5AkMJ1Ih/iXBLA26QusZfRocte
i9haec0P0+a21VtO1vmJX3lyuH/MVMdugjm3V0s+8rlzze2ma1UpaET1qp4v
rYo1wHe4MCD2ZqyBmJQH0duu2kqDF47IPG492Hl3/DvJQw4+XgIKGBvR18E5
SoUbjeTP3clsawc6f+V3sCYV5rTmhlXJxJg3AhwPNa7xcJ5wGnFoAuAIssbP
6CEO4YRdE7tIvmjXXMSz170P/cSassk6d8YB/+v3lOBj+7QG5aLGVMww1hyj
amhWvUxef84Trx0295Fkj/NsOaxsPQpWm3L3qMAw2Xqj9TG6ga3QuQC8jktu
b4U1mdIesmXhC37nCchj/4fUF9nJcg1EolHo8KdGVf83OOLIkg8giEHADaoF
AXpqJlJltcR8TNKcuuGN1CGz53CK27ip7OsPseIeoRElNZvUV9SVFkqRtDFM
GyCngEQhtwK/dz8PQ26bikwJQDbILPov8QLfnIeYq+WTFFUYwsQIrLFmZNGL
JXQsIRsHEIA6XiONgiq91ZLrncoPzlLqPKSfTDHjX1261dcPY11l9Grrrrse
c2dSOAVuWKdLtJHOMdw1n98p45gBTE4C1gqXJS7L1iBYIJ5mJil6VvDVbHnK
ja0pWncbN+XcuHe66uTntVUkPX3/yPESWrn7rijoTCmUWNifUYNK4zoR/fiE
hFfs+uKPesJHC+G/CxCRmjinqUAOqwACqqHLy4e+p/C7W0On7qp2SBdRtUaq
vYILg5Hq0pauULmntmWg9VcS8FUKb8RThGBaK6/pdgqveE2Gw5c4KOGGZm3d
h0IswqEPNI3v+47VD/cJCDXiqnX42jDzsfov0S5NhQ9xDw8DdbiT9NFGJ02v
pXyPDTbbwz8Rwc2HQW/OnoO1CJ+fu5poqNyPNzCRHQqLscPjAjjffQPQAtwL
Pe03JtydIUNDSHrrQQBGfOWI8AkE0E2v/6R3EFYTc+MRyLDblier/A2+U+ac
OMhEymx3C1Kay+bFV0V6zjG5Zz9RFP0z/HA3HzXqEHz77jdYOc1VKGsqAoeP
x3SGNedtVrSNxC/iuk23pPM1xliKH9cFIdfbhTX/0v6V0hrddLMB4nJsbkaF
1qL0vxvSd+rj25tSzVmaUxuFOKU9ChOQ3R9PVeFJtAlxNMgsQN7O4qoMICzo
wyzHGedJmgtaknS8taO2lo2RePh4GPnEfhKqONRGIUgXOZjKH/aZ8WOz9X8K
RicN3l1JPIrIP3Jdb3lpE8TfEvzDDCRc5S8Kh5Y4L/U0YBugCl92viFQikhw
pYoPY4feLhbLzJXbmhVuQPrYeGXISN48K/o/o0SuXRpZ9plgcC0TfbYqk2QA
F0FtawlGmCXrDq0sm0vAMbMlwvOwhqs3Rc/oMFFeuc5eUx8TbReVMpszvD4K
UUyibYI9rHv7ZmN8UcyWy3NUvX5XzAwnsMXi9mTMx7OUnRy9QtcsJ7iWZwUm
gHx7e+oi2f6ZRdAEoLVHwBf3IvNUqC+eKr+He0G5x7Fz+HqqZG1sK4v7IZ14
65OfRtKCcbmyyTTfoOilCf4Tb8NwyX08lF/nzEXr1W8AjmS1ZDr5dh5kx7/B
M5uC0jLR8P3QtDWLdKwxU/EYPwhBDEJVCcKcuDIQZd4ZpazomcVyUUJHJ5gj
AhSmsnRJ1cah76PNGZDldUatiOUOctwXJ+R3lJ7JP8nGiP88efkAXoS2n5uB
McQEFYM5KTthhFhQ0FGVbehrlDzyS25uFG+DOIOYuK9N2Zz7/B9Bybn5q1Ic
4KjKahqESgV+z1HL8GJJFJ7G7SaMNiyNsZBdN4P5yvGFo7M+xyeaNLvCY3Z/
VcKky1MO+oCFXGxSRv9I7d98hFP58hTQT6uAFTkImVjYq8MWabHrdW5L8uwq
Yd/CsyUJxBYNiWr/m3dutntM+SWp9endcYlIPGhynOrIZFLezS0T/+YUL1Y+
yJdGUnzDZjpKWaSXdZ87vDgT8S65ehHGhKwMdDcl3HLBy5WxMeLlvjrTSw+p
4s36YoiPus+3teWfMQGqROJkqgL5PFIKZGUxYImP4iakowl0ax/lRrmgS+Ci
42YVwKo+mjArscqdBML70EgJ5Pmw8KoijOySTzM6aAbhuSZBPdwR1JSCS0Er
d5UOo2hy0ZM5ahXtGIvDYGnIx9EtSvjVR6pzwO0sLJpJugIYiiMBADbJUbJJ
MDioizF8C57mI3ckpH+Mp9NEPlCXcL2Wvkm8SMQLMIrA3e4YYjL1oUTdUZme
Rx+MToxkjakytXNbVNEakBwFSt4GOQjUwrO/rw1FlZs8Fi0xqcGrF0jqPJwI
r69cZ8hkGbJb8jI+iTn2KhCnBkE05/f+N9ZkoXixWzT/1STKCjL2XA21trSl
I2U09pLukB3JOrgkB8cVGX/7qWMxyj05HZfLL4wg6x0ooJWDakpMRY/Ltcad
dyk/C21tFTFaF9uAL7vUgsj8AlH87WmJpd4/aTcMIcXqKCpAkRz5BJOSxImE
c/3YtQXaUyPawO//F0vf3ahUaB9BRxdweCblDFd52sifNZoMd+PY37Gfn44w
5HSc4TUVyjDWZ4dGc3Ypt1+SQ7DHMos8+IirE/f4uZlvZ3OL9QQsyR4bK7i6
gHUXKZqkXAm+taYJAr34XDJRpmx33GF30g0AS6l9cdFxCXOXCtEFIXlxXDaX
SWP36gt4FRGOGNfUhtUKCmnaMKg70dCt2B3osjtKyPlEeecxSTQG9gDKEt8H
MG8/XgJLDiucWQt7Q0hq/uhDMVlCRnOV0QlRk58wACQoFlaCWvDPcMr4j/J8
ciHxvhIk6nNCxNcgQ4gVSjH5/h7eiF81lhTOXkzOOFeMfl5h6MKiv2t7AbtJ
OMPhvj4UAmO4NG1ALCSjbYmTZlib1TVoFKPxrp0WedVlDjpmAbY+Yt8HYUlk
y93x3wHNXSTSzb76ct9hpkWf3GtQ32bji7H8+owOvr0IeoLgtYfQxtNoo7XJ
niuCJCvagCR+FL1JHYV+0W2kmOEUK1rZDpe1zyAr7fuCz5PlVEIyh698nV6V
fZjvqY2eenm6sQLvQUZ15FbIJ7XDuVNLUwKWl3bGYN8GMgFAn0cqwFYg2MPZ
3sxXUHOLXm+hNzjSHofekxud7CSd5DKoF+Iq0pwJMZxN2NG4i5P/j1JOge9U
TDCmBiJj/wCxJ6iHmvCI8BtI1dWNwrSBmiSt/jMLQnMttp/U5+HNq77cOxkI
GcVIjz39/po0LoOvO8AMNKiaMx34DVYTnj0DoIT15XlbFdRVgelJDnnn6dbx
VJWeKZFTPRhFDdQ5i55sxLYI+xfrOxX+9nXiF+MHQNhseuA30xZxsGDz98V4
SkLBVf+7SzbVenN3MhbyS+Q10lmyCt7GrIMv4NiLwK9R4nuHGFIi/HDPnvP6
G5boVQ+BbvJJYHHndJJKWUS+P2IaIp07AIysuu/MrmHHgzQMXit6gOuqHFDC
qcp4JMhq24ligxd1trvcrKphpchF2JoJ50W8Hl31kDw4bVqJrsXy+mZK391m
jtadFdEkpQ4aZS+1BtCB3vtMi/yEG/honRDpLa6sqREk4pGYty3nTYWL+Ygc
f1LXaVSTEfEXzoIet93Cd5gOE9jAO6wLGxgyIVE9/yyDopALhp90Xm7QIObO
ik+T/l0Nj8z3pV15z7DOvV9QMaMyAYMXaZ1d4WZB/XYCmmVPEo8rZUK3t1hv
uCXJd1xJdE8/jiyKkI5TxtSJfocmUHjMHtl9AxPl35PBo7vWFIY/nFZYMX/Y
tO7ehugV0KdNpY3s4GQd/tT247KdvEPS1ymqFfrAHUH6NW2dL80jedTh6ojK
ZT769MKNSMFrLQ3392RNqN2BJ72nxl6BQqyOrGHxasQz+KdBqd8/SqTEomDl
0x9NBPoOmjPWMilZHg08VX5R6OujP/P1/f1jUxH8Uoj1Eft2z9J13Hywb2dn
7QAK+rTsOJMXFUfJijUAu7nE7qU5Yt6fvSrlePmkZw3eBhVbQl04anODsWT5
TEeyBGk8O5gD2zBJeaDUmUHpEYqSsGKb6RCCnKBKCikK6GMF+NaDLwXaCTuq
4PJtAzVtEALk6enO/tKg7a6DfEyIXaOgFnPcZnLlkQzfHJrxRch8C2VXPM+5
pJTxa30xBtw+d73ZZFfpPCwN33xbiQllOZZUG8/bCJtYaDGG9/L13cNr9Vgy
kTf3yvV8fFOfoQNvGQZgKj2fcj7vpeCuAXokGmBUvWI+f9TbYW2gD2zaWKpH
sWwDNHIW68xu8hfshh0SbOlikLvhXhxXJbKTSUNP5ifnKywM6w0eu8v5+b58
6LF2Z8DlRRt1upmRSvmSdY5NJmB1emDXS2QYqkmgfu9pQD63NDX+UjdtfUee
6ESOUojBtD7CkkLx1ldd8R7ueprpvVmjBBLCMZlgo6WGST2O9IO5T38Tk9IM
5tM7uA91zKxlpPQewj79o4THhzW60plqz/+wD5+9Da65qvq2qesS1o6XOtDA
qbMO7KHzm4/5ddJPgjRGNfjRJFT10682RJfgsz7woLhst+ZBIXW3IFLzIBrW
8O70RSzoKKdAkcBBXlR9o+0Kru2a3DPJUOFa/blKmmPIgA7lPvLcGZ1Lk8Q0
LdFgR57Pl7ZUwdH4ONqc8aTqr4LEXGww1O6d2HcTBXn+lwkq81cO/+qJJYbZ
psiefuALcZWj1L++HP5OhoE0VebtOtTov9ddA/gGKYp2X/dUvKrRRjHaf0UL
P6f08K8tJLWEN7sbiwkBG6x1qMUUv3QpeV7KuvHgAT2qVNKF8TA6jTTMIHwy
nHJSIRv3EngyunxJgqJbh6vbYRDZmMqFKOnaIm3rrr1GZHKSdjznsBXkGzhw
DImxJib7bAN4ZwJIO8J9/Cbk0qvKKahzN/rLOJOVo2qeM2VlwNE6C+GUBKoo
luk9XvHXLwI2TmG6sCL6gdHgN4uueKw3ny3mtBi4Yxo4Tjiy+Gm/3ICu4UkJ
41xYydWgMW9/clc3nGClRfi9vTG5ARya6a2BNXihQN21D72mEjfC1RDAYyZ/
/RymNJqSl9bcjLcVO7fdvOdJs4qzcJNFmIvRWrWpsYe4hvIrWA9mzHo74a5W
q08CEdwrtl2a91NoZSs0fM6nJ9Pxr977Tz6lnq/bWcWEOYfCoMUMXB7cNWRi
oc0SkMwYpfsW7NkKzsLqyfhWNbHfUI6WiTi9w+pq8xV8nQWDOa0WDEM5HSrZ
L19YmMwIqGatA4AQbm/FvLTz11LY484BA+4oDjxVakCVmPqPX6T1MBMUljaG
3PnLyT/ilAwww/kSjHvlyKCdsr4mdsv3Ihl8jXPOHNZxx7p7zQNnyVCgcFjh
szjujc7TFcQbLVSN2rDbIest/KzlFd7WmDdEHa581TPf/zhf+BFmnV1xMiNi
lj/STjmlUQN+/DSkfU2vy4zOO700sXsZvtXWDicP6xONHKeCG50uaRaNP8dH
zNs8og+vSiteLvETwHilHRNK9lMwBhuOpu3HmmmmqKbUzP4gLYvi78cQE2rP
PXvtKOu2bzFp21QrQwJjN9iGUxffTjJOctrdJrJq9A1Ifl5zGn6E21sD81Ou
Wu7axPfMZ5x96IYAyUFJfiXhgnJPOmMPU8I4NWVNJHST9WTu33H5NsjIyyx2
K+y1puxbN06lsuoEvT61rzRuiaCxg8XpgsyDS9sj78NBolcYhAKuYWa20msX
0l8jTpbJDy9Q10l+yN7MTCvWJSJ+gqO3Q6PKG2zxu+rKpk3KMRrgtEXkyUNB
Py109GcOUbnniYkt5OL9P/JmM5st9Esm3spxdTcnH3j6X1njxBNDG/KduqeS
z/exayaSEyMBAluzUT2IDMBljayUMzlqg9YorcW1YqUbI6nDFQWiK8/kmQqB
uETElmvaj7F+O+0ErXtM0xvaY72PyPRGvbJTBLzj3WFa7ApQuSFQaYy3zyjG
2qwnNqVRJVo8Pg5QfsgwVDoK/8ZzjfJQ8MwT6gBXqqzQqlXQlBGffd34FwRi
Qw/0y6aysFPqESXLJiC85IAIF25lLF8GYLh8bYhZxWnx7vm9cH4NIiGsREs5
/AITD+LVnHlv45+PBxcyYVS4WkzhB/Rr8pg2mlqQEPo+QndF4hQoIounHisN
rPQb1wTQc5ffVMYKhiFzxRLZ/PdMKSXTCZQjwOmvNQEwELxL0Io//WotpO34
kSsFQ6i+CmmxRB2lbJo82k7qb1LXV4Mfp1n6tEs8wxjtyoZq7RQNyqgN3GST
3rWm3ZHbdOFVckIffRF5zyjRRLbJxLmyErQIdp/oBB1iaTewcSXvqaMJqV+N
N/wbNJqc91N8c4LrnF456J0RtuSvheJJqYLPJBEy3OaovmXneQ4rubqLWbqA
KdAh9UNxQgiqllRRNmaO4USL9vPQJJWrfyDf1ocRYGsJLFw/QRoPellFav4E
e0JMgWEQsdVCEtbhXYKchH0MP1Yg6w6OnptnsWFjhMfNe96MWzvM7gvOCdop
+zKRvmLhHRpZnN61dlmGCVk3cQ0QHgM25hA/a6xAmxu7+m03xBKW6tGKcCFT
GkJlVukvVGu+ngrHrbN4mUykwF8gDXsr/Amz46I7wkT34UOzXXwKozanFw8b
wsvKcBzcPeAmuI7vUuTYF4yK9ve0N9n4C+L3nC1pPetFqvS/GeS3stpyW/cT
8hrmUEVMKt886NeQd2ofqYIpQpe/6EB+0cxkSgZUI1nIVS3nAUDnbZbRhFJd
OsMkuiUYeY86EHK0PNA0N8dUYmeGdIgYVc6MUfTFqgwHnFVFb2+1yx6zELDc
oKuUIBe3VAi3nSTQdOTdTfU5oslxOIhmPJjSr/PYfft0Jl1zOYaol85TVCeM
N6e7J7nX/ai+mRmKppcdrm8SKbD7prTvmQHGP+B56bC9fLjkkS4i1Z56kclJ
0tlrvzbbs1Or4C2lsCWCLwvGS/HktU1VSH3GJQQuWuSq2VpV+8wJ/F+5DpN0
FElomsI/kG3K9I3fUcft67dIZTYfyohF9W3DyTQm2Rtt3JlqX2oOu1pRUSoZ
sXtIn3gy9hroYxfveD5Qh96onOlun250tM+Df8avEqhcTHlEF1e+jiLUKaBA
OHOlYIuOxEN/uYQPBVa41f84wzZp3ucaNPiDLCc1Sjgfu1mrwzoAFoFetLJE
glBcDsH7llLfnhh5+arvrgwgz0EGdMbspYyCSJcR30zoXwioXUCixSXFaTQ/
5qwuQVd9WzPtwt6AzyzdJAz6HOXzysXj0r+fBdOpcI6U38AHp3o78Gtk5jh4
tO6xmJxfQ46FzSBL/nJZo72F1f0w8MIQQ3/Iv+7W9sllTvHNR6yv85nfNkIC
XclsoMWR5pTzmNxEeqjZnV+XPZ/IoO5BpwcLEhnRQMysWx8+GSzX5ucKrth9
mHAwOdT8d59BnrmxuhymDtNWo6KH08u8tC5qNRqXhRemEB3jGnpr3ZlgN7wx
LIkrZ67zR2nlcWlpAZ78Hq/+/YXK9Y8usD8VxutUgtsmZ8xjXLyLLRN/vbKC
ahEza3QHE3k1aJGkX7PVWfQoNEevuNGicF3SYTlUve9B31yYr3s/3v4j0L9V
OyP94+2L0ZDXgTIf4gX9h/Cm+sx/QBENvRvpQex/sE8CjtBvQs6I8+QVgSoX
hQcsN10PbY1La3WWvKS50DGwJiAvo1pb24IXl2+f6SwAM/y6JEWs+qs+G+OS
d2TiE0RddJK6LWq9EEZE4wBrajxlq8nXKeLxbtXAHX/aD2U6APC+OfTF+4m8
eJkmmryXMhRtwYYaD+Xu2C4vrA9tNCK//s1NqiseJVuKN+rYDap+inVtcEdV
sAY8M36gkeBdYJ+66k5mn58C6jW+FTH1nJgcDLHpdRiSmscE7i9UMgzAGxhb
bskM0AdAjBQl6Jdorbt89ARxlVJAarA9431FfGMF25uFr3H4pnIjHVCBVPB/
2psQ6RMKRcjxnSexao4ZMSlczIgz6L2XAgtTtf1cwOKbgBFBGF3hLYku2D6F
3HcdGslY5O7/FV0SAlrhH/YQ+6jto0fhw4t8/aX55kmvGdwjcilnLlXyQWz7
MeA9aV6LEjBoPGtvtJSuhCo8zElSMgQ5ZjyRXUNYWOueGs9mwtvKzTBt0nL9
ZoFC8sfCL4KYL7D1oOpi9fZrI9qiBNl0+xGEb/jUMH3CuMze9IgQnOmnbMPt
tAd0PWSjrCYHo0KfX6vtivF8OYmdXpcZbjT2gkZfD31Jt8Bw2ZcyobFl5D6+
eElKEJ3oj0lKHX7MuLIiksD4rgTC9/EUT3PjoYUFobO/vNaV/nHI0zwKpESv
7PTUdWdG2Bqb6xc8RsK9LJzldUQ7VwBJRW2S+u3Dc7aLcheJ+JQB8l9EVch0
wQ4PRhWw/hKDGuZ/lUZb5TrfHINmZ07GdIJHEMiD3PxTruiSV9VZlpuRUnba
lUJpMcxa/iYIL4OlHb5gx/WQ2vDgTM4OjUBWLjZrXY64I6UX4euD6fb+U//u
an/I62nSJIIR/2oim/vA1PWzmHWqvyAo0c269j30Zdah2r1Fvqk5moTGcuXB
VYuoNrHs7xa4PIqYblPW0vW8fKqs7eLZADcm72cQpu7RWh6w3bph53Yyo6cA
IACV3q/mHSq21wiWpCNXLdu6xEMJQkI+UUoHupQ9fsB9A0Fh6NysS8vq3q1E
TIwyfml83rbyg89AIEskPXH7Qul4r4h7AfUlI2BQUsOA54jVUte0QBPJ5hn8
E4z9dWtPQo7IB7XT6eoc9MMPCChip1MyGrsPKnQs64R94UC84H3ANavnAhu8
BAGNPpXsdo0ixEkb9P6WO41wdDLZkbIH4qfxvCjv0aKB4rSQjLQW3Pf6dar2
+x9xcGaAbwnIKewFOBTRrVltYXaU0+0EBGCUcA5k2QS7/Gs9S9NagzkWt84X
w69pJb3Dc6DMl8wXBUdVeaoLUZeex9i9TgvX8aQsr/CU30zwmNeGdd+WAl2y
Rhc43m9n4F0d9zNskL2hSyHCPlQcF7pqjOO3CykTCxMdqwerX/c4S2c31Jh5
iJosbvaVNBBejD7cNh3YGkV1n6NV1i+cXmvxL2O73p8Nb8kS+JFLXcyvm/o/
RlKZ8Rx8i/nKhlOwigXkoBVn30ld59/2oQ6Lu3njYHG/tNfcv4lDoJuZmZIO
MRC+CDa2H6vbT5VMXTryAAGh1L6M7k1+W5my6CrF7g465L+/9g+EpWTDfru3
ko6thYCjJWxUHEXEpTXRicPn04hZ63T9bwe7rQ/NP4F1EXnfOFEnIfTGL+Gg
901q/l3QIAIYTsDAXOW+22QuCcj/hmucnaWO+T9EMGjpNh5HopdXV5D3NcyX
fMz4uh0jfvbsjqFO8L4r+3drjcCGP3A2m2rLuR3X53ATfpAyiBIeH3Kzt2Am
MBIiAsWKaNYnQhQIP8dhvGR/4wtNIm6FDlGathVdIxOJUAok10/ZinOz3IJm
jBdQPIQ4oId5P6mJCGhTnALV9Jfk8Ehg31T5sxpCq7ePCp9omBhBH9zDsNgM
M1DCprrRa9sM/IEcMqL7cH0lHNa3E58qe3V7V8mZctf5PBbkbC1Ziiod6YNp
0Wxb4KIsROJONcj8FI7InwqyhjE8h0fdpJyNI6y3tZG5a+6xiXTFSu/iAqcv
RWrXQJwTsaTplae6Fj0sZlyRL98fuj33sgwhbJiM3naAJS3ncs46RpOwSw4V
YjR3hKX1BopcQJpsYu0wvN8FAcrGkW20RbOXQEg+AhBotGfIgpPtFCnykshs
sayCAxiYLZh4xF4dHt6FLhx6Ml+t/bVDcI9IPkVu7+tHIqsNdBqYjO8Yhh+C
BDUBf56U0gGNXAykfyCqT3Ap4dz//uPB9ctPItFQ6+1kTKYpPSJuZXstOL3b
cqaMCiArgzR/9n/bvs/lVIjv/sa2xVAsSrJVh6RHwmvVyNty9G5ypDq8hRf4
dgt2ShKbzfxbpkKHopP+zZtoCtF5IXVgs5hu2bfNZzL2LSi8Sn7pCQ0tXnuS
9BqaQwJcffHNE1frZ/6eVi6RxLAAtrdG4eM7x1Z0DhGjh8GzjERfMo1xBDjv
laekMnPZ4z/W80V7b+75KBt/ANfm+Gaw8HJpxVWeBGsY021jij5aL806hPK4
hnuK55MZywo0D6D+A+gY4jdiYnwIKmAIO1W4O7L/fq3QbNefMy6cVDjjSV9+
4IWATIsHa5B3DymonqykY3bVU5CGb0sdRHCq/aEPbDaBbIfJJ54aIjP0uv0k
5Hnt11lfAP6ijKdl2gaM4Ap6STm/kAb0C9zh9PlJ1TV6ifiM41Z2fA91/hqT
3la7BB/I2wsKHwGL0ks2sxAGEw+r0xajmH2Q+553KoDZjlqQA0KH5VURYOkY
VntQWU+yG89vB8/CdvrS0jiP8JYKfIV6smJct6b6WHIFxfkoILigV5+J4/jw
MsHg0XJmegIkSCCc4XTRFcYYPz5PSsZwq+mGjK1ouodzZMylWQlo1JeNU8H2
YXqq5Jk2HYTLxyhqJZin52XhKfI1q05UjFNvZT/3EGecczpZHrKtuuOLO4xf
6UpNFJZ8efI8Sx5j9HRrWAv8ZCfVYPxL0//80T1H5Qe6sEgOot4GLrztoa1Z
XbuwzbCD2ocl9tjo1wSIJi/tBPQiwiI7Mg5HK7MFvnEZiKvjNI4nX1C6WEeZ
gx5hMLQ4vRpVGpTvGiwMUyN1OwXXF47X0h+dt66aAF+TgvjzryEz1MBVJzvy
0pyP1JUBllWa4YVX8nRUpvu1g0S43gEikULE5ToQM1wNIeW7bb7WSrKjD/Ay
DDZ7IhRWAxGalqtwLdMvGyGj8cnLrpYcw5gGIHAlj5tFqgh569r5Rz2kFTxg
v55Q8v3KewC+OCiQ1kqvoCJMqirRABj3HUBzNSAGrq0Zi1BEm+1d+8LmeDdC
J7MbcnOiKhVk2RYe99ADwOkAlVUP65+rHurEtS9sHzEgvLLXZgnZeUvt9Uqf
naciQJOqshjqP0wFCl7XWBQKrdQ4xr2fkmTs/tykZG0Q74ZsbZotG05PCkgs
8Bu7UI1VjXpTXDw2WG0EEiTeVR4sA3u4ejGmvJq/xipke9q9j89//ISFLEwS
JHg3PLwLn/eoOtl04es6FWcLwROHfNHPrEWZRDvypSBl5Tc13SO++ikg3WwQ
C2mgyCXEP0UBWGmRKt9tx9LJeFK4AgQnjzcjmz/145mPFvMiN3Cms5zwKrs3
MpTCKo9GV02oQwr7V+JVZX6BLUs3n/HZulZUCig9fkYB9CKv0JZMrDt1zs7W
L4XmKZ6VOVvB1RhVt+Jsv/0GVxMrNMfDFmq9DFd/H4vDe/99gkQ4i1YnadDd
Q3ZmaS5agGdkWminR3s4LGVVWfnsMMypfraW+YIMdbCmbcYQXqaepWEUGSI/
miZVVthntNxGQHSgPzrC+VAtQjYV7NGYF/37iasFFVhpIe17M/WEgnTpgJB0
1a85ABPU1kODotySjB9gQfJlpqJRWF2CeLmmu3TP+5aJkBMUe2WLXbkJGRBQ
tk3hqwxDgTduks4uI65+cRl4v68QNimOLN7mKjs3R46eJ4NIU7VCrZgc6fpm
6roVwWO2WYrH5oo9siDEpD4kwrL4sOPlAeaXB/N/2PQ50o+JRfdDWoHsSkod
Q4lv5ip+pjlEVTzOdgSf7qE63lK1fxv5vXsl8APVOQ8wBgzbiNHsUDeHUfAW
IxN0FRRzfQz72mYdM7kqo4z6ve4YfOW9mk2RQoperaiCAgNSeFWZLIzwLit7
yL6RMb4FUYcytDSOmLQPHVZ8X8fhySkYW0oWm2DPir6kP9+mGpf++aqijVz4
/XRZ1WWj5ESi3qnF1s4C8qbCNc8ElWv0A2/WKMXje2oeVDzeH4OEMblX05uR
cJHkskKs6wV3accqmR0JGeDo5f4dxOd9zWLbhK1+ZGmruzq9tUutZig+oatx
v/n0o5Bo/PxymAe5ksMLdpTxEn3zFjY4kTb7CiSuV0Oy4CkonXha3H4y6NiO
l1qD8FNeMC3rcDDlt1SUqPkzKJ6ySAF6vW+WoLMfEcYqSuKaifd3c9Lu55nH
yFvq7LyPaIEC3Vp6+u1/PkscVeuGToYRrrE/sqxLLUcZL7AVqMXI1yZH+feT
PXQwPbDupOceGjksPn9GT8oXmX0b3mDV5KrjZkmV7Gvtd7UIk5yw0PVz3qvU
Elyz/UoxrUyTnV1PoEIWTwq8e+fnuWwOz4DNbWOKcYCckSSQcXwzYMKEu0bv
E7WRy2v4Jt6SrpHPIOA85YtmO8GzIta3SdyfGin966XQpyQ4faNRVi39jC1X
gT32Zv/zCd3KL6zkfzNqhvvAQMM7qQmmZtX1GmDaZm0zathDN/xJNhMZAw4c
5uqpmZ59Vr/Ac6fbFEuB0XcB9zrQ7ouZUHNNp93zHxaj0qfBCZedMrOLt4K2
khDibstubo3qTTk4+BqUwcInbVWy7GAvnCy2sBSyFRfg9rvkALMFC2s8oBnV
sHjfJShv8dLDa+Z4Fi8et4mYbkjq1gbjdvBKDhb45EQXocQF6Z3vb1sVF7Ef
FDmFfzVgF6y0Guv0h34u+ldBwjdohuF2D7INMIbKLVMm6xp7lUaZQ3g3Zc0/
ebyfjDYTBKvoKNMT95qDZ4UoPHAz1USyTcVQmgFMJFEyQgr+bPz+4lF56yKN
Onz9wA/FsenOPAsiadwdnw27Q+IiV4wMVu3sZRhdWboayAmN7v76MIStUokS
T/UmYTb4P+cF09Y3U4VQ8MOQ2ibxX7oXj4VFlRamK2B8iwHjMl364T+I0FtS
fDO2wjHj7GvGQzvG903otEP2ctZv8Fa4X7lkkqxy7qGibONUssMgsmLFdHQe
5P4zoEDN3KIBfUFCRmRbkpVG7BOmGkda/a3Q6sPvDwO6xCAoCYyTyeyZm01v
nmsTc6DAhRIxTrXURSZyPPT+AM/R8IWha8hoErj42KSwMeTEoE4kNkmQxLG7
9v2+2dyHnf3MIqvvwPaZ564XtwBCxKcGKuT8eIUvdzG03giDGlYu27CTGOa+
fc5yeCmNDdZbrUVRJCxsmk8vu7qL+D6kprKpiIZqxzpA+de9VFxcAe69Y84a
Nq/Oorcpe84e+dgrf/LqdZDgFg0wBGqTW9k/JYWaYRRPwIN8LEXweYscvcXO
z0xno6LJtMDXRnEwvjjosCYO1IAh6rzPHtPabBI4RDEIlnaGdvRvgcRdaSdo
r07uzpGA2a2tnLAEwEZcVp2amDX3qSYqJfCRRNb9VEbg+ObcmvfdOW931oiK
8AHDRRG7LEWiHqYrQPi0x6J2T+KFH0cCxmi1mfarviSnn7q5wVlBMe7liUoT
ryU72KcP0GKNFNCb5T8AMxmUGDGQJQEVguceU91tk4IKIbUgqeNvtGIOvk5y
HqM2Qu8gR1fMAZ0xW3sgf1Z1a2Cseml765NjTrlHGwXDXKNLa1clcZB+/P21
yT5dpo57k+OWUpCEPrSWoPBBJuQJob7wQdKWU49/EVLxGeQC8XMjTYF2XGbf
wL1R4WTJtTPmMaL2NJXQLzftc1W0XCg8NUOkMeSiz1u/6ioQOjGRNycBe757
QEzaUwXJnngSPFHMFyk6N6oXpdHmqJVnn4V19tXZBtMabrRNThEOY9aCjIos
fZVxLt74JaNypr0ixRrrJXO9NEJXAe8RWNvIvcLwDXudC3GPLgBljVv2y3vC
4KT/srlvMbZOhSwXvTjuN20KiggxdwR+U40mzK5Si2Bej1/e+LqSQHUr/aiq
iBLGrLXGv1egiC2BbHK7jEF48SSrSSvgEcRHWD6YkW13E6hMwRKzuesAv7zA
l7JojF3DpOrhaw0xs8JAwoca/aj41xTIwS0a2CShpFnZf8ulsAWWQjvgFWu1
x1s3Z8gvideSaGnnuBP0D/CiUPAH0QADjjlRh2ZeDMe2kKofC6rYYUVQ9QNw
KZ8w0UORnyaxaa/o9Lq45VrPQtVqjlHbyeApv6NHR5Rrs6wFEsTTZRWWEST6
Iz/pu7m2C1fuJ57GcwPOKGwUa5hG006/se0RxTOtetOYkEaOzVcDWOHcDWtc
ZxH+ep2sRQNJ9SU/AIoyLr69uQEkmQ4cE3eloxOxyz3SL+LpqQQJKyvUk0s9
38hNufbu+z3i+6Lpw92A0i2gsiK+TK0Fw2Y8bIM/vwOOBxESEjrHH1ibhqM1
jSlooFashaGX2WoP6BFLih3xU04W76/7w5V8VlNGSAtJFznzUyU9k7rNvaUa
6XxyB6/z38l+pkbDR1A167ggR7AoS7nbBuLWIGvs4iM2Pir2UqFGu/Ax4WnN
fZDLQJ2Vt/zW3kGnplErgkyg6YmKIQxsYOHaf1Fcbp9gnWRpOSAD6WAqQFDz
uEHWDBGAMEKtpa4kQPNHZH+CHM8VulibuW9ifODGRJe1ZTdC8Fskn2/Ts/Gd
eDtPQ4hXrSW0B76w0B7czDssykO6NNLRkDvyCuCjdDt2oApMttq1+PCyZsIX
xvj5ylqssDjNjj6ANkeLfKyVyW1+ZshEiu2YMQwalJzbKc6cyX4zg7+h4ep8
i0qXvKc+xiaAMvenRkmE5rEvo3xZqmdDNudfAkb3ywubHG1MHf6iIc0HSzxU
RjvNio7DJ/vKiuQ2N8u9ld2LBZVMMh7eQwDdXDa7A2F66vCdv5SYYRa6vz9a
5fInfPE5/IHXrGDe9dMzWNoqyLUOjYEgqE3x/GREj6cl3cK/lA2zfvpum8BY
0Fps+wGLXxZfBOb+yLjGsZiQs8pTq48oDLsegF8GU8Y4McGhrgST9L/8hZEq
NtSbD2z6E2KknpI0YG5kI0ZQiMmT4HXxa1XBSvh7kYRag09ia0B5fef2qLw/
N7nkOKk22ZfDxUJX7Aj1ImLzsV9DT3PCRDT+njskK1hiBlbGsTepQqN6Zyo8
3Zwd8oQW1LuqGpTEwr0fje13cNsXuCViK0CHWMNLGVe+1jMT+6oLdFxh76QE
FU0TRP7RJNC9JM4uu0vgNuOLB0fdhSETn0cSfnqpO3clKJZYvrGXkH7XdUli
u4UWTerqdKP0bqwtFXGdBOzHxYUQ1f/rVJocc4aPt9AlfCIRYPzoiNv8oLD4
XVnmohB8s+cgwuNcw9K6LJycQ45OM484K7TaleiIKu0Y/S48VUez6/WFQ9Ft
IUxodz6uavx+eCVEO5R3pYN8SHyBcZtuyuwBM12ud7IWXCC7Yaul/99BObLz
trsnT9qLAGvSRzddwRDpa8eMaiBzxi7dBFqZPrtfw2fH6MIYenmiu2Q30f8h
2ryF73G9U/DGmUhZafdeULsXYb3fCRZzEVUDS0PNzyHEsGCKs8//3fHBX8EV
pB3L3C8DqXO3+b8RU7l3lx/JJY+MtzlF0Ae+fD84LEoDJ3bnuuJdqG+8zgE/
tQACp88IiCIA/hY+oruscKt4ltRKZCPERNSxbFImIMnyaW+mxsya+FMLz7ik
sOoZ2QtfccArtIuDysgvTYhrBzxoYLlMWlSqXF3W+4N6WeeDA4XZV0i3sZZR
A70+ctPsqcIF+EdAIAlD8pu9ivXeoop28vwkcUb1jjGZ6dzloImbKMrqbw3S
FyF5MTdl4+BBixozX/wlj6fl6+x8KOPQtZPGyYexdi+1EJ2PiOmucfLICCLZ
pu1GlZIYHPxYSH5JhP5CInNm9LrjSzUieZj5G+kea1PnUUVHqR2e7Cn0hGNq
chOq/9SDWcPm1PhtZuE8852jrC7xzezKDh1Px1HJYbTNa1+b0pH+hZGjalAY
6K8qxpamPRuixIJ3YrdlWR06azGEtcJ7Ru5HFvpmuBpuGb99wojG+E001aA4
UxtgJWFeEgOtmhJZVeN2PyL4Fd+sduarOV2xQrJBMNf1d6whveaj4dw0bkuf
AD9+ObJymi5cMrui+HV/QbDvLFKaThYvV6jTXx6ycOWIs6NEN1XLuBrzf2q5
exfNFQy7lXRcb3kK/gAG1AHB53uColtRUFgQ9PFLLLZodQa5bvyC72i3Ec00
N7HuVzNQ0esqKDzVQM9wCRxA46y5b3NNGFc3ATGWse2XhNoHMYT3AnFRMyAr
zm7oKuP3cHtAUfmUV0kyuV/jmwHJ5lLxsNJdd3onmAG69MHMVN53li8jsa8i
xrnkheSrY2cPi9MQJPNausH4I2traa/cbT2wa48Tob1oaP/fPD0hzlhNkNz3
4ZFZT7zMGBI6lLShzoGk1pI2NnilOj9z32l2jvsnQ39B8En3HhVTX3Vk6kbX
MKj3bDacxXWC4ONNhgd2FUiHsnC3pNmfPG48FFrR0naewvPTPGERhgNySN9C
8Z6cBWem582hgv33s19lF3NmgubIhPESuzr9TNlgVEQvs4BeJmSdgAmTw8ry
pQvUzOpZQEbjG3BAnapR5K9pqfflNAfN/LYSBr9VVScc7/aSLsnW8BH8Vuay
kL2g/NP4dlZeVH9ydORZzw/lmj/AH76bGmLPoBTbuCk1ln0AuhSIw9SqagPX
Cudm+eCyfjHJCjHr+eBQUZd7Iw8iNE3R0vobk2wuSwPoAex1QMBP/CFeQ2TI
maARH6zsqoNxvzBsD2JQkBhOtL2IzSrt/aCc/xz2aylAtFggc1CykqHU3An4
tMI3llWFgx/5qiwPZDuLFIlNwSg/VYOOqTCUfQ/h+1hxWAfjKcdk8tf4HY2b
HeXT00bKvY3y6ItSj8wKoKhdP1xLVhCBXfnM3QN4p7FApgTnymXugkKpWVno
pZ5RzZq9th+pwtEvAVwcUJMBxazXl1x0tWuMyyiDCSxq+G8BvMIHY9Zl4km2
PazUyCvf8CEiILcBUqGKmSspUy2bjPV9m6VWjLutnGbgZ0Y9kNp2XtAUG92r
S5DkHg/azGKJjbYP8hpM5aWhz1oWGeEUiChJdTyIxCg3NryjJL48C2cZwvBz
64Jb6dwN0PH56VXFWfy99dp6UtiU2cHqNJysVF6zLVwnS7o5LLBRGwAi2U1W
kkFWGKhIR0HCqBk0dbmXLvXrCWhg4TiVMx+4i7MbH1k2S+8XQvgWJ7GZsw/4
+GRaVY0T1fOXru6vbV6YIsFdYNqw0hJofGE4Ji+/1nWDQTjGzxfuZ4UV/+ys
f5DGN6Jl/SR1DbLKvXo2xgIv4tobu9W823PP2pgZSBNcY11jc/33HuUxe873
QJP1F80KLufKFszJEtNMpyqn5cRbHcdM5VP22fHDl7uNaOYPGHpWM/4DV9p+
13WbCjF9yzx8cfT7mNQvetRaJNdRbCf/cf49hVkTP32WtTxDz/T4m8UEmLrF
8yM/xYNbq/KjSbbmo4CEOpVvjQeAbcVmfHIu4GJe+vQmt58luZqW2LO796zQ
ieMVqg/g7Ih4iJDl+rysR04w6rrKj60LsrqSM/CWSuOq7GrDvpoCYW2CJP6Z
9N0naRNwelO6oXAbleIHuiUHG6UI4eevZc+HmaxqdoWlkXz8S23dxkEKCdoQ
qhUuyDDDW1ED6geeBDthn1xURxI2EKm5kw9CEAlK9cXE6KrD5P5xNDVRkww1
m6gP6Io1FXwlQ2P+AFP4ZUFddIlGCmaxSr+PLI/e9GjOv/tNlUtPlVkOG/Sa
PEMbQ3T4muSVPfXaPSlpWaWNfZhu/HN58HYKxY9SfaIQcgfnO4++yJf16KVt
J/zS1wcjk5if4OhF08YVmp1104AcPWXAKlXhRSLizTYIJuYDaE5EUEljiXgg
YRDstVhZzA4Ghi319/c2ESujqxvbpb+kno3F+TD05/V+57CrHfjHxPy//TQ1
ngo68t9P9UHRoGnDCzy0ucNUHAZFOl6ur9/gR4gA5e0kNSns7EM/XI19E+10
5HPL7iORZdHhRpDKYtjW0RjKyNsN3f7ruR6QxybwDPX6SzhYxb5vPOGeQoC3
y0rJYEsydAOTA9i37kPv9VU0B2MM6GYqFx4X+3iQzFUu5ZNi/Hg4wuZU/HQZ
0ARzm72SmBlfnFUUT+w9TbsiDRlPcCMFFIs8aiMi+zYfHYZD5ZoteSP7H0kp
WIzIIqhaMlqD6K7CHoqnm0/PP2haogysnzxc0pSuXi1xAYBtu0Dm+y4uy9U3
4Gz6bnY8ADxf5D8F05xdf3uadrUfGNVOU/hbXAdpAEmrEULFDEdoXTizttbB
1RXPHh6E1iNBNYbUMdsTSEvqGzBnQdSo7OP95gKoEIEOdgMEZ72aNG6DdsJ3
FFQa9LFjrlizLNGtZ30Lromox9EiVHS0067KlARaIkNdMd1O7HPkwjtbBnRC
WpIhaA+1muj5/vZVR+tQoD4HLNaf1keN9eNv0i1OtdU5BjHrfliutNp4NXiB
vNfzupp5mAGGyodaAMkFNOqJQ10bBwYdaYOkdl2Yyup+9+JsH3YLqEOC8zjn
rtoPz21aYZPXRQjkcaulIE8gvYQMrJQcidDUAALem7z2V9KaSa2NbrJOlN73
53lx3cy4pbv6G6vf0Q9KwFj00Vjboe9audJ6MhgyDE6rtqOJhoQBEB8JOavd
TkFa7mVN7Knm4QFG+zDhYcL6+XYWupgf3C+qxRBBnqHP/3DtcLORVu3xbigt
BohykY5huUTZEL16kKdFf9GbzxYAUNj1LpjHLOHiFA2qPUSfgYUxAemxjk/h
HBPhWf2U0aT/lFCBgkjgYajaFe2Qi3e+gPVB8FcybPMAVt7P0gWEV+uo+nx+
hC4Y902s3FqgT0GjQwyosXiE2487uvm/xk4xk1LKWW1mKJkGhOdQymOvtQya
tuHQuvGkfOYL/wUnhrrnBnwyEwoVdNIdKQGFn9Unpdoqb7B25jrSCbw3C0PV
RCF4nGLEwdD1yr6zEGROLhAs7usdrFjcggLiZygcOICmG//kHYFxfo/woJHp
PesL9IU6WihsSSg64rrzgtDWW15uYc4EemY9VwRP4+e0T/G1c8Q4owp9HouK
MgrobJqJgi5/h6A7PFDmKcOKAwHu6RtKhPEHqQw9uoMOWlRNgzDklHty52ph
w/xtdZPCtI5m9KtDtYogM6z6QgXDPcDPXmQHuZWY/m5iP44WsuU/K4zhqed6
DRBv+yNJliRtk0CV2TdDJfgMGv0CfxATsqePRbNS6+6OaTg5fdVwJXy2lmhY
7/shX0OQgGyVDCw3XJOHQ+cCWfezLJWjmytcel4BGn18fkJcJ7KJA8LLX5jB
ngIhZKthLZuAdZQDL1ti23G0KUsZatyuOaP9UGM7HcUsdc+/Yj987zPZV5zN
W9Idt99l8ANoEJ082HuRp9b1voDkJef28NRxDvHKe8A2pYkhMK4AHO2KA3Ts
oD9/jbncR76022ZM1A6+k7z6jq6909rjqEEyBTfXhSwH9nW+r+F/KUv42hFs
MmEtxDM0nSR0Vyy4sXqcB12vmaLSokp/2T9G7wATU5Ek49oUJ4lh2QyARlx+
lfpdWASfM5rkCPPvpe8LlPcumue8T6oJFZi6h7lDGthdVvg1TqdlEHYkt9kr
ZhdSO5xT6uWznn54Hvm4k0YPj6ekTKM+Qj8toHTIpuD4p1dLXuweRIV/uQJj
T+Yl90sO7vvYr/o+eDlP6vVr6nTqrKkhNAbBuEvZnompg24Oi2hjovGFbDAg
P6Aip10ss+ytntMLSiBdkHsmXJuiy91jJc08iS+V6irhzLxxG3ukE0Drro7J
t+hfx3gzuldtccCy2l+zSSIZ3fG7g35crvo+xTxm4PFbw+yIw6IbVe0ZZ+cs
AtBI8AcYsU1TtNuFO9y+jMFW63U2JEaM6FxlrqZAehcCS5/NxsNLE4+FklaT
EhKOhyKpwcEdUvwUwv/EJD4ifDsFFJnJUiXyp/NjjeYVYc6Qb8XA3z2ahrNM
jkNwRWVdgLVvsJlwZ8e4GvYywK4NZcY93eO5WtF7WK14Zt841/aihdSf4mGv
DXAwP/sAghzeLwvhusOa9gXbFuNcx4vHwfHJeD7YRX8OY8vfty73DA1vnKyd
QYrSgOXXQXLahZTjbYS0Y7Za6gy+uyMSpVZU7Bcd82EOAnhtBTzzInFCKn0m
4ZK8x5WI3KLU1n2cbpqC8EyfctFFJOsKWQj2JpcJ9rqx1GPWSXJbpYluCGYW
vjnbHcUZ5R/G2n8/aqOcpUwGDW69DCh/s2vvDhX1iXxEMoN2oENEdtv/h2gv
m1trVp4ebFBD7yKQxrk46GoagqcCdR3cUtB9aG8/Ce4Kh2yZs3w1iTPRZmz5
3lm88hreYvmMN+VnXXyknkgSFjfMRnk8HsPdRwQ0OaviWO7Ib7eP7DNkQ1Sq
WEiWPBt0377caXzyybeMs7Z170oPq7m5Qgz5PLS8dWYjWPHJYdBpbp3PTiFP
waQEHEsQPKY0dvg16WOojVvGVmM3c3hsal4hBLF3IMwfFi5trfhD1+Ixjq/L
Q/r5m4h/ccNdcPbx7/lL7WMhwjevQmjoYLaYnKsvdCRiikphiEn4k4hIUBSM
5WJWKk1C74RWLdsbkebFF8NZzJqhCsZ8S92K7jMhJ92RkgRA0YQUbKJFiNoR
v3+CDUg5hwzQWqppLgyHqZH0mU5hgXy1l5nKFjo2SJodfpybBerr5pvuQmB9
9F2dABuMWZeW1SWP0CJJuSbuGQhDBaeTpJNDFQd1AyjyCE+fKpK6jySoW0OW
Z04lqtS8Zb5NnVHy4H6EvIk7kP8nwb0IaS6EwP7z2bRKCB9fzhI1KeMue+Ao
jR7D4I5tW4Q0T8U50QjjEI208u9Vs2n8TqMqNScnizTj+R1HcIBlLCZcy0mZ
wh2JlnWoofgFufgL0l3wQtaeJ0gYxxJxhvHUIkIDrdYL2WrpKRXA67++XLxD
8ug9+NdxAIj+2YjoKXqfVT7HxJQVX8t+FBbazHHgwm1pZURPqnyiRIzXd5kk
uU3nnC8rWYkkGj8w1DZY8aLMLl0+m8tpwjZ6oNDLaqjuRas88USpnhx9893N
0rk7GqYWZsGKOR0pPJT+1ms0X6YRDC+esLxe+if/o90VtbYYZKBVXCI6p+kK
HopNJ44PMvp9Hfp3YJHaAIqIK+MeQEuXRI+NKACkWl+4rAuqzTwUgNp5xSIn
XhI29C7439UFOohJxCTScSKaDOcmrcDE2buDm0PlhC5aIZ1VdKRQWQB68A4L
VxRJ2HwGgIEYuKMDq4NdpyQisyKFa7h+CRnDQrOnRGmf05B3dol67Qo1h9F7
Vs7TFCTdDa1juuudxHBqdmCBEaunpR0LNqxe+qc0AtfgVfpZ8nGilAnClpzZ
vUpn6kJXRiLPLuCA2w/+dSOmA31F7U+j6wnQApdKYzHiSSDCMZaX5Yw9gUgr
yVSXCOlh8oZNHzgFbramjQBbucwu1Vi/27DTFll6OmPFAlmdl42ZzsBXquAV
apAcjZOwGf8k2EjjLlk7maUi8D34iiOuHf6KXCZYmZNYA1622geCGIyFN9py
ZoHTGFXzBAyTcfoKbucbEX7w6Dl0faFUXqnProhK0oTu8QXng5q7MJ30J/97
Gzu1xP4YTPNUqN2tmREmJcVj+wduoohB/uZSHCF3fSQigEjRtXBYmfIVE3EW
zjeOjDuaSaWc0Gii/24gDnwLgcbNp020EhJFyngwOboJ/gbmPOoVPibsFWW3
RdaLHRjLJqC70bTOcry4NKZt8If7RNp5D1YgmZVDFrsHwSO8/KvAhfkL2efh
2HDNrp0UF1Qu7Rsvtb5UBVCi1q/V/noM5JypHS5yH6owKglKSA2l7jR9xZ+E
eox82JhUSap7wNlCBGcswfvm1FOO3gGc8+ZYdnyZJMBL+HEbc0/l4K2CIIcS
oYzkM32g80/Rg12KwFnUSgiQ0WlJHAuOpXCsJKNIrpb2ISPJI6hScwMWnuz0
BpUcLGZSuatMIkpv+onTUyzRLHgMhFtFpZB/uo+5R+P7ZX7e7gILtk0k+Sxe
FqvoyfUZccwRd2QoI8EjafQRtUGxGlV5seiPtZQgIsacrR4oYp75WT6T63LI
YNV6gtghY2gnbsYxf90t+hsUYl1/zK0WnlLVdo1i+rLlcpU4VTGNqycCodgP
4ZG/KE5dAFeZJlGuGkvIF48uN92dpE8PLONZNYEZMaIR9kzcKIUSG8KLdQFX
+o9RIyE/3MMDJ6qeIPh86WK5Pe4hlpyFKvsTIY46MVls6hQsvkxnd3QXGcQp
z/EhuYTZNj5N+XaAQ5THLxPX3q06KqnA8DwSsvuNjmqQCov4i+r5IoMxfcAg
TGkIKa5OBnVHrxHM1IcXBOI2laIXGdBmAUu8nK6ZqAsHdbl7Vrrv+Kg8XZ1f
HXjOiTaPQ6sb3ovc/HLYsEaB7v/mhSFBMiCl0BExSzbRXM+JXwB9Y8x5tM1M
MzSOYb7lYc5+0/Ya2FP0DSHoPEt88+kZ+OZisSON4FwgTTS0GhRdrejDuMHv
lj/200bfZug8/st2XG908+4Ab8mcPRmFxMg79bGfUrSzrumZhxXQ8OAkNLfJ
fAygsYFP7eGvQgfQD/DUOvglBqUlK+kNbYl+wNc8ychpOqWZ7lsHneM01y0e
MzFvFxZlWiGk54l/RP96wu8W/WzGXgBWpWNBJojUZ+F2xy3izo/oyWrQk60W
UbZ42DmNwyQ/DIRnnV2tgFbIISJ3VUGAj6iufyWy13Y5Dv0koTCqfHtyblZZ
4YK4qSiPi8Zll6WgfNZQ6xozZ7mQmtIp1hHocEjJaYHS4HwpZ62da8kQUkXo
2TfN2M15PHUo7/l9k3UuV+7l5nBMEiegO9fW8MZSIrMS6/emDIlveqXliaZw
nwQeCKdyFfumWgcd7FJTYMkcoW4+ARAly79JBWMQjvQneuXYNzgGwFDaG7Wx
6j5gYn2XRPo/8Xa6kuo8tuHkJDbpL+kPMDsnKul0GIFZVx2V/GVSDSdwehEN
P4UB1gIP3AWJY4pR5unoG+LhkQcV8hgkAY/AVJOCOElz0L2V2wmh5ve603Ww
AubpbA2G7Kr0jABoA1BOeVbwHKiXNUqTUS9WH3XmmzUZv8xGkCdpNG7QHm6B
XYfn6M8L+lBvV/vE8Y3c1aYBu1lGg6cd6GiggryK2hygcB8vgZ4eVRMa0JHx
O1YZP1zc07B/R4daChMxrbxqW7Hm9Ic/1/qx46nzVMbgrhTOv7kCO0QMrIOi
61XEcPOqw4KH+SIL28P5AZRKtnpdwlxCWg7kYelfo7jt7inv0GywncWYFUWE
KyYw5NHIUVZXEOLkYjZqGu/96qaPYRaFGDRMqslR5itJpyHK6WuYuEO8AvkM
JStU0cchNZfmDVeTg0fErTQio/19b76dp4XHyTLddi39GPupA1yQX2asn8+N
1vdz2QA2gzUBhPkwJRncU9OrrjaGCgWRyNB3prn9DA/u3Nz8wWDF4OWktMoP
f7Ink/Izqw++v9GNO5IN97A1QlfwaCitNncPziBZ2wt4TzuJj4siGvbW8UYV
ZKCK8jK1AoHS+cfCrQzIrBh+ovP2UBFqN9YdCG12nu7Z9Lb1ESjuIb0mtiES
ZU9sWS/jRH62jSpL8PSRz2/N3AhFujXY0ENOSjck57RbL2V9hnuk78L8w496
QI5zSoV9BTT/Gfp+sy+kBW9aHZ3ea4OyeADmAvU7ncxhSdnJTEIy7RrLORs+
bDnrTPQ37xoJrW3o9oLGxdsvr1Jf4QK0mRLRqPpqOONg2AfTD1gZHd8RUt0j
LIofB0WZjW+zUU64CdVG+UJJjedxrUA1SVf3HN5MnnoQqB3SN+TV30W+0+9H
35wGXqbmmmxI+62DkzgYKvQB6ubqs3qihD/NG97K4yZl8yhVDGskxxeNXjJ3
V3CrUnStAhY2PH1Z69u84NosKKiXDQKA5ZaDNyyLgLSqbRb2LLOEwsjnpqHj
OxKPmgTrqUlNDjVUy8oln135WT3Pq8ksQHT5xiXYFuG3fp9IwDbr4uROmjmF
pF34M8iPaPd/uTaBFtJ/x2jjcTF76KWyEWLWIJmkvcdBJ8Fnxm9xj+MO86MN
Mxrc54ZvctRaJF592J1J0hmEmqSDorEOuUb1L27GcL/Z6EXU9v9y5++W8x/L
DHEw4QTXha2P2xQZtMFEp/JG5huvHYxno/T6H8mL+CGzrU2ItEiNPUXAg8Vo
D8FN8Di+MiiQ5dyPSm5NrN7l2QfwathumfKxG9rGMvPKOiMWb9DPieekKrau
X7SW5+AlDwvMPEHvGsNMooG8FzErCxbDTA4fZOAY2Xz/4H6UFOAPPpOgzQZd
Ai2xBBEqJJL1pVKFToHEhgS/UrZZ6+loS8nqupJ9gJudH124aATlIa/iE86B
+VLHbIaen1kFRVfsFg5VRmmcTkFu4XU128D+1honhGr9WO2EsBj41v6OyRQS
VVh8l+FG5KhTbjYgEy6vFiMtgU+UJLtx2vNW6luH8yngb83lLiWYsscChf0C
mT+Cq3U+8GktFG5kFqeVWI/seUp/sppFtHLW32+bIPrepP0WUzM8XeOPJVCP
wo4Smjys07pkB+QruaXwQ6PzE/PlHttp73YjT9Q0S/bwmVw05VAf60DGjmj5
b5wjwp+MTZAxdL58unhl0UR6osUDKyd4jun4HJw0yv/ILToTaboMepxf60rV
jPBA1G+jozUHg0AvzHAVNVX6Ncw5rcLKJ9Z8cjpxJSs4FqyqvFMbiPUJquWe
PzG6bqjZ6rV4NsvgxVggOf+tkolE5WNawgLEOO/xavlti/2TzorHTnFLNftj
J4cIeF9gjSk4v3UkV27jTIS4KMzJXRmYldtWhbAbn1qccZdgIsHN/WHIgGtu
yUbwNM5NydGDe38aMpZIVbFHHqlry9gEtVZce9v677OtyCz3OxTEXazKTU99
A/Av/2I+ilpXHlP8oRh49zJsp4M6jofLZgO2Ty9hlv03AhOA5WapntTOE2Ud
Er++cU5Qm21EC5R8kskDjPEJUtSGUWDMS4aa5bq1wH/gV3KvcROUvXm6NopQ
u6b1zY1mph+X9J738UrbGEuBnLaBxiZyosY7v2+u6WJnUvrNjDqhxcoUqe/C
aDrIWE8+NHabAaatLSnjo4+GBB4opHEvn3ZPhTs4z4vyks6XFVsG2IQsIo/W
T68ikICam8wKAtjC1iSED5o+vqs5GLzcfLj6xPPnJvlyxAtDVpGL3884WxaL
YCENGcBJTKfZSRfSZeynUeu6X/s3IbUAEieOS7BgfqCLz/lraMKP4C8rvHb+
l6HOReL+of89RsQtoAZ2XUjrHeuoH8hyb9nJ8SCkbeMsY9MLHEtZ1TJJOCO8
YjLvNJrsjzIcjEKn/ZWOZ/k/cvjmS/kYNPyD0XgCjei6UctqdU8EF4TWvUQ4
1+xM2jUBhZeF6EnjNbsolxMBwcJNK2Tne1lpyoGuh1goTO96NMIN9W01Hoqe
yaJ1xOT8mnc/glrNy7bXtTN/5Gx+OttN3HoRYiQNo3IDe5jvoL5sQTLfaAWQ
G5J4D5LD38a8vL2bDjTQKif3OargIpO8DutXIP+49sc50cXSXk7iYMcPfpo4
CYrVlzylfhi+Pse9Is2muNs9pqUdlavI18WGa0RkfwRLhyPCF0I2XH5AxKOj
8ZGBnOo9ko3EEz1igzywL8ymdZfwUUaFYN/r6NJZxMx6IgvEF6eUEeWQjMBX
UFLL7eTeeG0WxgCINpflmQHxQjnciFpS4ItJymsaRTthTmJAM7OCR3mxgRsE
FH3Lz2xD9gKhEPnzHZcT4X3MKoLqGD7mh8hCw/IYzBG2lf1V4D6NPT05TBKn
cJ4lRxew0cG2KI2mt2jY37DGQNTCuNR8wSVljp42qoHQ9/wH8WBwUDi5f7cR
KSvUTgWnNOR7a3+Wg0eaSWDu6LPrB1iZ9IF1Qo0EaddF+Ow+510CDXs8eC79
zp9us+7Voqk7DiZiR+kqMsu+WBJM8R9Yl8F/FUnN9vtW5SKS+H7WTZqbUwTa
9In5ROiihJlLy4HwE8Vz8+Qqaf5JZ1OqkCDDxAvl571BjnC5SH9/rboyl5re
qu6+nGhSeLEq27Y9JbrKWacl2FKUthkcBabksCEnqVItUPYTlR1E8JDFf/7C
mdQFWwFv+/Y/5WtPzohm1timf4xOraeZZVp5UJZ1+5RBT+5fLHBRcm1WjI0F
acVMv1JxAt5L6f+kpu9HQCrI5SLHCp79NZWau5KWVTgGtWULlLnFWVbV+Lay
vuaeGrA3yIYl4V1+p4k86MPxgwl7Ciiwsa3Aun4FJC/kApMp06HkDD581713
8ogXx/0KjYqBsEN03rra1rTcv3C7+7JNL93ZQRi45Zawc9epTw+nrQZW0Cdm
Txe5MN7+0bmJqOV8wkALkXvjD7GO6TPOcsmGO1IMvVz6VUz0270XlO1j/u3Z
zyvQp4tMALFXuY3KjVpK0bja54fW3hInbAfKiT4Wld677AgyIdp79tqsupLo
wg5EWGj+NEGVMRH3HARgJgKbOPrTs/w69T2c3nIOxZQtMr5mK3bNrCmAUNx0
4rR87PDoOaDtlYT8DEV62EWNwrVocFTN1HqA6+7sCauUaz8NYtkjRxi3z6h5
UFYSAl33Y7rPveXbieLBDQ4pJtfvnEgV3UENHLsv4c37Gd5vUGHrJyk+GM9V
gzTYVtapRWEewo6iTMe7x5b9DsUTgk6lo8OJ8jAiH+RFdDL9ObG9agtTYrR7
Z7BjYG0hhXOaG0PCDvZO119XofMa2lfPBDxaGTO53gs6TfuLsuD90qHnKXdE
7bP0+m5TooKWQV9l1bvupZVrmgmKIu26siQInVosl/ubjSkYT9Sa0ByYQ6GA
7DDjCzZWIQMPZ9tG4G6gRRBU95Rb+nMka3UkMU0Ta3UX9GkeXgrkNY++rSe1
84JU2NJpsYRKHOD18DahtTRFrTGKFH1Tqwh19d4E6Iuqx10P5ysrPrJ+l7Qb
wHGmWZASUan3aSeDDT0CTEZ83qEIDT5B43rBMw0/thAW/iq1jOgBSqOy5bRB
j4ydzuJzCfG659RiHnNh4R4O/ueBOfQnn79hxtADzWwXS84f6mIZeIu6CROm
6y4AwKtBJdcSNTbJJZG5L9GiPeIGhDMP/OrKtCNs5QA0LtwGu5MnLjljCYQx
wEcX8A01UfyPDOSOABHIGsOIzsCRm+VSrnS+jH36zqQ9A6rNEFyBup5ZZ0XQ
TSQoqRThrRQ0QzJXRHXCOI461lrEDuMbUPMLpI+VbZrummTbKEvNZOLxSUlh
imjlbyfQQMfLLiBuXSx38R5x5skXNFJAbvvwos8eecAYYPtTGhj2/VBsxG6w
XKoUaPgo+CdLiRAvbVqX+0A5w4vuTY5tJp6OBtxFPjVfBifJHslcseWPbJp9
6ixOTVCzMH6ysbczEPOzf7dNU7sSDepsfwqc4lvnrjN3JwjLYAOGZpmDgFzm
TJhApH5Oje7H0G5ZnDf7WUTqfCeUAUsjsB9Jrz7mEC5qJ7P9OKhIqX+1QIPV
c+iK8xEOGx1Wc7k1x1jW8x2ertIh8lSsvS4J/UeK3hRd5u3ekd/Ryxsw+EoU
Bzy9m+VqZhF72Zmfsj+xDJutICl2k9T9yqW4hHtAkoI9fSWtM4cDFb4JILcL
aONLNIW1+F7vvx7ha1hbhzIe8S3DCjE2Pz2LaqAwzaPuLD6IDg9GGsh0eRgK
D7aOz7Jro1ZHjwwF3UjQufoVi58bLd81HhMBEBToQEI3nxDYBVt6OorRshwV
Z0uoHjfLd21Ksfr5aN3OWFZvtR2fQ8POzIWCN69b5kAb1Umd3GqHpW3/vbUO
bRCyQwJzNlePBzBAhY91MODi/ndTfUuRyvJMbhfyDBC+p3jUgIdSkj2YXyut
/lU+pSgT+Dj/lojUrx437e32vGkQ2RxnDkL1pO6vvizivazWlvbT/vR0Mgir
Bxtvmj1wtIdCXjDofejEQO9U0zgHP0zJz0lTXHdhJHcJWRHnfqtCcJ2jPZ7h
eHN6ksOQFlFfkZ7DlcdEBrDnrvIaSbt19YTX9uw9SwjG9w5yO3U+FZ6geXDQ
mzzjiCCYS7+sW0/SBDBRWakXjT5QFtWxw270a1qSSbUEFJlKKtd9cn5/i+sH
I51pDLZe7i0vx+QciRltqaWwooXZCcTP8E6BQGUvZG78i+fJH9tn/VaykMOG
ik1Tp3Iom5Vf5Wzgv0NO8FZQLBk7ayn05W2opQ6ZOWwDjRCodHYPronFOTXd
rQudF4PzimNH37i9JHXOYTW9ZqC30DUINtK8RHOlvdGiwLzE3CVgu62ZJ/ha
t0Th16+8sQ/FIoj4oWfgpvttoMUx2dG3VFc8NH1yLXJfDfD2N1qRT2fHuPb3
FrbGzWkRc/+zu2NX/eGSQlweJGRSAoSc9EE7I/kOSvxBdHoRnVeqtB6ITmiT
XiYRzW8TiiZ04UfeMiggxdlrpEieUYb2sb48+zjwPUwFtrGV/195XFaDqcvR
bMfyvbHisq2VoNw0ymEeKHt83wM9hbm/j7XVHgSU8zHGnmqfiaDp03G16dcj
GT0FeTkFw6TSj31n3+v7BEMSPVbkuqPb8vsCSaEC9t1fkyx5XQQ2LCVNkPiW
RmUNcVKsSv/Ac9YeYjogweRVPoTohu+oQmr3j5N/Nzhc1Gi5+FgaKLkaAKeb
7nWHdKmGN37KoYIZwO7mqbKqhQvugSPdnB6j0gZcUHkRqcjl19eCCFiZbPE1
IAdsDEmZufSr4NtLpMi0dgBBb6/6cgjPI1Ycm8S/YRzGadmD5foM10FfV8ZO
waiEHKDWvp2gJ1MzFSRYQYrwW6jMNIcgJme6FE8bSeSE/D3v3xmK4DMKfpyZ
akreAThQmHpl0aITilSlrIyW26kagiyOz1y/5E1pVSvd2E7V+bk9me7QL2Mw
QuIO0Q2vPo1zFvoyMIPTFEHi+L3bliRfYZcBjpvzBWyaeqIns/D4egrH9c5g
CggDPjuqUaB0vSkICgIOW2Wd0D9K2iFFtAsHWKhYJ8c7i4hJb8RaZWpFJFpq
WWR1mCxkZHHFmc61WKdDtQv8r5NQQT6mpfbQc6Bh/l+bF/V6c5/7Jf9UDH8x
hIksdm1Qz436Ity/PdAv/Ecpq32I1CDYUaM7SOW5ed3E+QeksFqFTsjafPhz
gQgBMhWbA/iypOjoE5eEk/Mr72lBeGa5H/jGgWzjlgRPWFy+H17a7xxy66uk
OyLWHu3EK/ynNSvDuuao+yCsbn2wKNCM5v4yx9PhR2ProxMWzQDYUtWkWp1I
DZRLj8UX0bgjSIX873qMUWhOgiBV8MrXvGoCbHGHm6y8+FqWoE+5N2ErW7v+
wjQ5rq9j1WE+J7ZHeDqZePCucRcrBcl+GNFxhY5zqZUCm/RJGh/LdhM17GGl
GXCYz1ceV/Y82SikMrCbwiHf2Q+DEcvaxHICrsVFjOwR0UDFASLlRHdHL4+u
IZpfF6fM94jgEZFXOX0867jYf8enKKMIgwjhzwvy6XzFsTxuPZo/PiF7Y8Qo
TTWD80vXe0ocUmn6FMWJ7HaG64NMJ6D/OYe3ZwWqYww05ymo4IFHg+Kekmjp
EIzpBplT4bun/X9Akc6o7n7ySEkjEMCDjI369eN+CpFhu9m1TEnrgSK6PSQY
ulBi4Y85QsEVS969VNoV4AtjzD5FNH67X0XhMXWARfyIj7j6HXS3dXUjzH8X
m7MBhn+f09ieigGtPJtQ+oiwG4Q6r7Wk+MyIW4x+Ydyhy87e1ELHgiemYqQb
RulRcdXaJxH3GlnBiB7BZbnRfD0TXgvh1hIVSfPgN8HpKC+Zh8AY7rqAY7UY
FDe81NGFNCxrQ2fTGT837qwYrlc9ApDmcrFBBZVR8Pjb/BG/H33I6FoHXvZ/
rN576z/3rg3uK40Wzc76Rm3e8TseikWyNWID2v4bvZHaiQ0aNtwdwa/bnRFT
ZokdUBKW8nf0OcewsB39OXjf0VNtWlwb0YVmnxFyAanmm/Zt7xtudbxqPwGi
WuEd5mfALtRtu85ZvivN7dOYpwDOUFrHrL26OpHfPSN3P3PQFe0F2LWmgXfX
zvj6OeYQfmI7IM7wl7JHQ5wbyEWTDblmAMLF926OXw0QpqWkv9GCSu0cfNdS
5syOX457rNJRT3c+2AeU+147c8lGzL5NCZYXZ+v7Wjzjl6+YsnsIKrpRbep2
1CkmXNPf736Qq/gOZZ4FJHCsvfkGipPuxfXMph2rJGiRGRycMhW9ug7ALBIW
LtAjz3CrcEwEYTsivk8kqVh82JE8Kn7BsOkTS340ebR1it2jk4/xN52jT86q
hgleiI8pB+lM5WYvGjKQtoZirAtirNavdLbrhj39n6mMQ8yAXJmrokhQDZlX
MRqiXesN4JXmYR+uAU1O0qRjIg0ihaH5nQ6T4TykIJIV7wezONsGKCR22iBJ
3zsFqUfGsBo1uvw4JYI3f2t5F7HfQN8OmBLfYOdDj40FoVe2eYSwYphWTml7
WwmP9N9Lf5bzD3ow+E0Qr+ly+Z+MNnJqdBhUai5BZxa85vyOr8Vi7SYtfrf0
40wszGnGzM0se7s3EB62eoNlyG7JAPiV5s2195wu0+GgI5WxW40O6e3ylf0/
i2vZTOA1RxdeOlMjsXULyxbDhMntiaUXOYiFLSSm15/uMPOMWcDFIvhQfe1e
XEGJJXDJ3VbG8pO4YOOsF++nXV+rvYCszgHlmJ3N8yMjVKz3pc0bSJwvH9Qg
9iUBi7j47w2k8IpcXqmpuaTktu4PPvdjH/11OERG+KHioo1ADpEtxgR1gl8i
Nuz29AUWhN2HGziPOpmbAyDHyvB7e3kwro+3RarXP//1cs+22hgUBo1m1uDA
4iS1INkN8fIoCPtcYe86Az/acJhHSAV9YwL8LpXpyQSaYoqIfdzOTGplYwfc
tf74Kuf169S7vMwHWLinuAUYhierSUKTe/vwW528yNWbeEu86TPMoYDefXmt
Yp/EeGsH/l3Zt2L8Au8JgsPXk4GPrIEzA9g6u/+fZWLwXB0uDYXUIZMtgB9b
F8NX2vSGaMo09JQjOLD3mmtaPoc0nmpv3QBHz3KnhvzCLNeb1ZDFX+e2ZjqL
8MlmV1AhqfiQbiaKltmp5ZiHpau8kPy1mgGLuwdI9uLBcdI404nf1yjaWxh+
9LF8BNqFw43SmqkGCcQQaQM5QaAWwBzuUiiCFqfVSOYa2ioRgOAsQ9qPvlVf
XeoQ/CymmftIaM0btoMOtP1sC+6cjTev9LG4cFf0rsrbsBVgGF5jDvcLux4H
gX8XpxM9is6djeUQjg1a5JqJnABt5mfFHzihhNtMH3XchpTo2R+QQoV7sFnE
LHZ8cTEF145m1ByQV2LmKx7JjWVjpqntSv+hq4OmsB954QVyDfdIhZ2F86/y
xaBM1tzO4x3yXJtSQRUxd/Y6BWvrI4sMSA8xe5JCSHK3mWo0b8CVjekyR/J1
eMnahxNheSSwPTCjb4ROTjQc6fk1k/3F1TrUE/k2fvpo5C5Q7Bzvo833i8a7
7zLGj3RpGhBRN5NkZVznNWwgSEa1BqVnRwJ8IveSW57UMrnrmLxRVprXkz0S
uDd26OfmeLc8eLc+2DASYfyN+nbxMLQQ44z17fFGuOBDqmMJ7UXV2O8mn9s8
Ik4tdXT9z7Bc0fBsKuAL8iTisHuOpttrgBoGmN85k/81QZHmaB8o8TC1NGUk
SVwwZam7iRTnTkyzONFXdFGlfAdqIrBuS28DQJbTQFJdyXWYAqKhq29RZ3/q
9gZiXHh0JklMD6N3sVhVi4FXLlnqf5/8hXK4jMuzkuazWOm9MPIuoEGOcb/i
4xQ0vs0Vv2qmWvNMCBsGuqqTWMUpL5Phi5UAwaOArKyt99gIjUJCNELH8ce6
x4MXCg22o3/nHP1a+B0NEi3F59Kzlgt35yfsmxd6G0498xeR21HRiEFoCUUo
+31tVMIeMMhEmqw+H28Tm5B/tbg6eCyxsKOrGqdFW5CWLtDdiwmvXaUicPNk
9Sw6Ho30PsaKdOJQqqBL5C+8GzMe8xshW1Zt1NMKp3XaMDYbA+u9JbP+1wIh
p7CsP97y9X6WlQjZRbdNHXQkkt8VxYkpCPIISOmt3s/XuiqyB5t6j74TyDOu
AMrnMn4NlLO3ncS2eB/dO9ogIfftzRbTQ5l4O9RfIbte3q6IowU8Oztm5Orf
4RUrA3KGACErQ+0pqATyDCcrjsoBN/hl2dYOXf7R30br9qaROLkDpYX0wJdF
BTM8k7skiiflHlP1qCB25CfKo6mjoPpuoQSbR3LziteJ/M/QVykJCQ+KwnQl
+kv+mE+jm2M3qfxJV8x0zWs6A98AkGMOEc0XPLA+rD5dQ5nkzdN25NxD4NMD
UGH8L3b8l+GfArkA9Hs53KsvBSq8A6CpnjpWOvZ0SJP2uNRPGJaA4nVUKmsZ
TIwxWjcQF54gUksSIZdaem/OOFckPLLXZp4Fo44HwVol/IDpylMj7HVactR7
sjE1yU/2PyffqXKFOnvJ12esFNLGFi7QK9+DZcbBu3CP62GnimITrZNHq0kE
Kr9l/YAfccMeIYZQJDTHLz9aN/LIQL4lxQw0jkFFmLvgQQOJhuFpIUXpZQ4L
2OOygnUBzaXVzS45HG0E40jybUcciP+KbOp1Y/jzp8eRcR+QPiTHYvEsOI9t
/AS+pp4EMswkSLy9vJ/+UMeEIIyji80s9MaZPa+JmfafuVvaODUmcGTgqEOK
Y1Q0GKM2fnWJvtOJdx1prWIvm+6PwSX5jVM2UgUIRmJvD2E9klddx5xbNgY9
cFBH98WNDy///H7tjl3Td3QUn8lfbW15oBSWYy3k/NfYEYesMq82L9yUXJnU
yAPmQYbCtQMuAE0uADJsFvUaSQAuFd7MP5ZfhVvcC18o4Xi6PMJXClMkF3vz
lov//7LR16vDjE08nXZsol2kwOZWDlUtEodUxKLBISNvWZbn9KCUfcBzhQA5
xten3T2SSeOjeBucJLA5zJNE6H4EfdR7s9/2kX8tB2JUmeAAW6xzM9D1bpjd
bvorGrykSmET2YB/Fjnk4HfIr0Haxb6fxumxhO1emTXYrYPyxr27MsRbrzh3
j8mwNUZw28XjyLIsMW0KeMV/tISlRUM2GBVS/qWu4QN1RqAUsqH1Djw9zzjz
N56/uWOtj3LwZh+VSVWicnh3FHq+z8VfCFfqhs/8hbZG0ekF/IaS65++6tIA
EHuKBevWIQ7dLFa6pXjjYxWb1u7Gn8SDljC6aKUj9p123eUJqKSJvvLB9wtR
GcHa6SOBAkFD16xdaOxEzuc+ZQf/llU/MlU9atyyiG1Osblp2uxtk3TnR3Gp
Jw41YtAn9iap1ybDWKBO6ht+MV1rkxnPm4qXr84UHIeBL+wErdpHvtgwyv6X
B+ONGutthf8U8pJPNGAtISnnYzUNcu0z+Z0amGD3EeFfyoXggp8jM2Vgs6qR
GpolLn/YwiLJ7vBeED4pMWhqcOUTGLZYKHzeONVTNrG2CIWf6Wswa22ar66g
96Egz7WbSjXfNlPpILKo8Ni4m8wmREqbSAcrPRQgBaJf6FUpAWCO2l9TPy0p
5tiTqq/vMDtkmSAiwq7Fbx+oGZuDd0AXcHApB9WYvpk9viUHqcaxtmLC2pg5
W88npYL02uWw9b1CzehN/2qQ59hY4qbbzmlH4Q0c659X11Mxhc+DI70k9Zk/
i6oAjfHg/82tmeWiia+bwK1EENj8UEB3D6RguTx/mmttn8oQfa1+YFK8zdUF
RTlgNORkX9XHn0dHeRsxzT3VJTK77ubGKkzmUsyUYmW6fAlIWVe07AKI+Rb2
6spoKQpL+CFu/olIEo8HTjLVppyJ5YAydffYxdjXaUznA7rsxj3uHDMl7r59
XFqz0ia9ijcFYc1f4sVk+qGlJYogIbHo/eiLx9Sm5QROuF508qF0Kzx5LDqw
kEREuz6h3OShGXoA00t/y1L8ILnE6qE/P9srz9fXzNFHvCqb8MB6KxIXULK+
yeOR3Fj7UlnuNwESG5VYR1AeVXn077ziVjZSFp1WT7MzATLdY+S/mteShtQA
NzwGTLVmIhNO5de5Jdedrp4yEnEOKLBcDXJJ3dDX7s2L+y9Y+CGRfM88lf4m
z5KoOLsieDkuEnxk7KCXtvohUKl3zlPdUnngCRmu1i3uqJrLtOPEBv4KH93v
oKMImq/KbGGuRwUbbASGnB/xwFM3fZfdCDjOZVT/YBrxZlHuzTjMxkcWkSoK
q9VYFypDPU9bdS4QI2iwHIUVLq2kkjw5fluDZq1+BPBBFeKzSSKZ7GzcE41E
UzFt4VBhLA0sYTmAiq8gg+k459BGjDaNB2h7RMitvNI0UHCG/bThXqLrtXht
E7GpLTOmOWAvSCu8oWufVnclv/q5Q1QnATYm2Eoo2xovpgM1lLJKfEstM29R
m+V5WWGAuJpdENqHb0cPlffg3xgpbINFO8c2A9bbI4XqOdJf62NxJbI1TFH4
OYX/rVJFzlEEihL6w2dV4H1nwSEYP6hCzIJBoh1xZ8GuivNOFtSeIo1u/Z0g
9+HgoyJRKz+OhS6G4gW4Yo5rBPUIA8XYx2kg40TLJtgji7VPv7CmBVfNupFi
9jRp7Q7ygW54gtpSvmV6/JiHPOpA7GjTaFlkKFPIPgmipkpVCJl674bqJD48
PvdQ85Aiuxwtj/ABIX2HkYtMZUR7QbYLitFzNfzqIaWuurPcO4GwNGafT9hk
3rNTjJjKWOtSOYVSm7Y+rqznc1FdxsIMKoKikkYt0oI15l2gsy46PkZvD2DA
9/pRKg2BMN3HqriZ6/DJFvGk4L8Rwcffwj+sPus0g8mrnKXK3cplZ9987WD8
HFZt4WefqID/kq9O/SccZPRfXLu+ZgSm23+oqX0L8DGWZQfSV8wRDW3B1Ty6
i+r4TlB6yRmcHMU0pTEsZT4KkxrUksHb4As8CfZ0b4mpz+y3LFta22GQ2k8e
cQbYf6yvTAVb+8DH/F4aodkHrBPweHwrwNUKceS76jV5N2SZiBAbJr/1wz6p
6cJsgsvYWY/2SlSie9ItwvQXZLshHWj1yuCqaLzeEvBzeE9K0U5i4klGX5oA
aYn+XQ2XfBZ2FtvFqtUdx44FG8jeDD8gE8ObT7E8TN42ieYlKUM8GoSKlo3L
8RKo2v9ixjLrFkBnSK/35jBuQZZp0JSgCZ5EaIqic3D0688SmAZN8jSaAXj5
6k95/9LaW1fsFV8xOV7cv5nNiRap0RROR1FKq6XTdymKI5LgXD17KuzVFSrc
uhE6Uz5Cq53gdJXP/9296v+wSwpJkiz4PMgo/8wxeuZCTkPbkqtjuEYZSv6c
0ToAgh17cI6HMPauVZpNzkAPwkLz2bf1qDq3u/X9KDzSIzdl3kGHY25gnMi2
zjUeMam0qvZ5h8IwtPP3eOH215fUfXSQBNA9a4TvJp/QJMPpLc1TLwo5m+tB
lDPayfilAiikB3eb63K5/aXkJ6D8rzWhlfSdnQVFqM2ET5imV1huuPGnKo89
oU+0iKXwLwATGxUmv7/q+LsyGzmv3CNUlJNvsmgmdvS66JZqzYH/F7KSf3tn
rxmlKxajvOWPbqKly+zg+a9SrsFl37iiwXJAnodTLnMPPchnM/voPZy81zrT
OsS6CxuDHPwpVysJtKiLZHpDBszAHonI9bzfktCzSKGLVeqamKcbuGieEQyh
Um/pBRK4QCOqZB1cC2hfcm1ON/LGwZiVvN0ReoXIFHU6Ad1X/5ao2EBQxwge
GXyakL6cYJmt1x7Rlj9+86t60K8XpiEztGJ1jCikfwSVGYnb/O2i/+4VCfZ2
uxA5mc/EzBuUN7yPKfdMvRPFnMpkhrPEWGFwrHsMtkzD8yLlK9YxFMNZsOa9
J7sqoa2crWeViEca3Jtem+WFUTLzkyM/L7xfeYtANqNOvW3KkG22+Zn4+CYO
FFe0lFcOLWNGDrzEtrLF/pK2V2HPjXNf4GwtaEleDTUAzMSX/7Q0b8e87a0B
j5J4uoHCgoLndEvcPtrFlm9UOUevUrO4bfAL+JVzL2jRzHQYHAELui+dvJA5
YrEOSiiDQC1VoTk1QgLcVIxMZ4kBrjUzRa1c2Z4HMGYDEUS8G6HqYJ/aS+0o
ICAIpXVKeAu7GQJRqxrrxgahs243ET6EJkf+5Wye7OIe3fSf5o1IFPvzMu9J
OZWl0r1YCFNFog7GglNNaWlkx5lCyBZqmedoZ4LO3CuVQohCwk2qh/RESkEz
wWHM05qVGCjcftgVSoMDdskTEh46u9Fham/VH1GlXHnKlgC6/c/sCIc6QnwN
mxpuV+GgsE/CxU1TEYpR5kYi9nonQ9FkDEyyVUCR9ciW68dVIW8XKEuxqCaF
rMpI7nCPQ/P7UpTDAorxojTHxo2kjNpTiKbD/MDWIw4dR4havbHS/zfYcTjI
Ytwi2uCbL01axUD0kG2GLCRK0SccEbbP3F+f9K4Rp/RPrsoyhckB1Ef9r4C1
a/rG+HJvTiPiobSk2ZahQUf0U9FcjJlERT1bYhGYAwjEpWOXHM1Sy2mSjZVl
x3DHHUCgrVqCY+sG7dLPGuWPGlAWMq207XSaAmn6D7BQuQ42V/jW5E+T96f6
QSpRB0ccdbJeU1RERNpG91U5wwcPf3MetEacG8EGGwZMjfv97xcQB7c0HQbd
kGdTuvU0QVSOaQCQnQ26oVSCep3xurNYK4FVwvH7M4UCU6r8LgyetvQYls8/
v2XTI3KrX3YPo/TPZQcottbG6No7A81gZh8sHOnx/wetHx9tb6NBG4PfE4Sk
zdb/g76fjbag8FZoPY0KBvNxR78Khu5loA3TDjLpR53Xdbie2gPfxrmJHmog
eySVR1zPPfUDuExEAaOtynpPr8mXnowekqDeh6BkbebyLqdmiuXxK9xgE36U
VzP+mLvE2aU1GNI3HkDPLNHgYeqXEC7Yrm8nFY8MsmBsoLs3OZi9d+re1mOq
R0U5epB9WHXF1I3pnvRb05UHNC4XIeCWUc5DUXP+gGt37Y3yDsHHF97vb+yt
D8Qb/bGK6nKxZMyCEkkGQ01xAS4n54ciivFP6jkj+u+gw3uO3P7HUZebzh2J
Iwez5AeIneJNq44i2uj06XrQ9rssjHL4LE7mZvTzgOYD5DoUxkUS5NNPrzET
pLfaSqn+mcA3Eb2yzQXRD/bpv/EOqH++HSMcLgFZ0aabMW2GkH6N+jJUlMoc
qAg50zaqE1EWuNf/RWhrTCUe3Gd5tB69IlE8xAuBM4mWVRjejI8tv4CSrAlY
Hf5zz+YvKw/r/6RLLbDF2I7YGWd30kXqS1KegWegW+hZ5//odRFjt7xo/VIF
hw+8YOKtZegN36CTybioHSQoxwiMBbIiXTOWjTeKaPZofmPZB7J3qNwfwlgO
dwr1oQu8IAQ0/fYqwC59hk73ZW6hi/7MRtjZvrtd6Bi9yObLlW+F61yjpFsC
0qlsHZbLZwKtK2WbS75+G3HbR0e0uCgU7PQK+el6ZcsmZOIpWwzV+VLVXLl4
kESVAkafa7Hv/Gc8w47J/xNID0Tg5BiQLEqJM/A5hKEQDDBJC4RUHIxESf0W
490u91M3JnA3gaYvEizCx7FIuA8gHO8jxAqBh29AmECQxvxiCgwc4YqvqxSl
m6dW7rijANUixHv1GFLwNKrA4On/sseO/j5ZT+CoxCBgUWc+hFFgBlrij2lf
oxh3N6+wf4HhmbYbY5Uk/rnuiZxOkIjngFND8U4mdNYzfmKGz6PaJd8duaX8
0cKnJwP/7Wx1bzm6IlzbEOK60AHye3a0WD69QlYjZ2crn4Eq0AfR1U0AUtDn
i26BSG09F9eqNJx4JAXr6d+djHgFvjMFTr5tp1w6zgY/MbtEIk+SdjB1MlUH
Ky2HzJLYy6wAOMaisaO6jIH4ojrDTap4aimedY/OCTVTqsQ7BQ5n20Z7qz3B
mEJ6RN5wBVPbDxti2I9eeXmYz8RJw4eG0kI5a7XFGKPFXdJ66EKDLReFOLDY
uI3Nbf0b1iPryv5VebFdrNi59yT5OmDvo/bGoX2atX0Hxi4E7wYvJ3kcbM9C
L69B0qSOAOi2TY/f4vEdGFB/orrB9qyoTxCIwsq2R1Y6J20oKWR/Y8k3ZFdS
edSKA4zh6d5FhxsH74wZd/9WxiPpykEgXaMlB8M+WAGfNkB+uKgp3BRWAVWg
nAVzVa/QI/CEp1UYz3eazyhBFE54BXHnDGHaPoPMUqHbryjD6rhnkr57VNmf
EbbA98x9qX0ReJsmixKg8kZWpwL9HDBoGlKcr0pAtoU/drMq+dWqzHWghffX
MuxhnOYliaShVrGMdD6DGnddzwvZ5Ya5Gsb0uy9DTjfOD1F995hA95gxkpv1
F5oDnPl5qhL8XyjgEMLSELUdJwO1ERDulRx8CYJA0KQCxrwulbCfMUmt3uc8
5EOJyjEoKhGPB+qFrbcjNaHe2ZKA1YPz+Dj9yruPGWfnasHuYQxbeH9nJNLs
ZwzCyi5GEc5HS0ONUR267hIHiJbRF0UBEhZgRtnrCwNYdnS0/9DsFWjuDorw
WFj/O/qcr3luGyzDUn0pa++yzi8nOUmVyFk4J/m9qRDvJ52PLEwlSGKK/ezD
e2rqPKzLXBWN/gNeiW8umbP4FD0nOs2Mwbsf5EUYkg4mIsXXl+oWj1joIDIK
WNez+IM2+5acFY8P28Sq4v1z9udFU1M8i0TUJBhZTUzvbq6tkTpBQXvbTQI8
cXP7BMMMLmzHLyLfAztIqAkSq8DuBTDLiZk+VEkpnTUHhC1ZDBuGlTqraSAh
Rc3OqwvG2QDptxJcP+JnBbepZGl94Q4dnyUXsTUgEvbDOSuK+lRBrq4zmHu4
8uPNMBOwtaQNEdyEO425ccjpjxwfaC5EMQgtxG3oPJU52pAbN/uK5rF/LjK6
NeJJ4FYLC/fAkD4lu3cYdKRE5bGNBFzEBqcIKGPGNZZfzmcsPYY+KoMAaHZS
xeeF0AS/ixfvgAH7pUCIG1n6wpJLVGG6zmCICa4NQO2V/LMZJpoWT01nHLvU
c9xFGVWNsI+8ZyHdoHcsnBdLt4/gSrPU5ZvJYfhKffPOqlADqNT2t628sBmn
x5w0x/6peCKVs1y2z65o8DLTJeknzHY1MWIvyQ5Kz5t7q87mEQa9GNIvmK1m
6hnynreLI6VYNGWWUeBSoRMHH6Sl2MLKr50AErQNjnxHXY8+QWfEb5EZ+v6K
bxau12WoSLbCgu1eMRdpYayim61n2piec52Aza8QhbyUvgrj0nXBNPTHHD7X
louiu8BlX0/yCfkiBuL5rVX7O6QW81z1Y3ouDlB2akvpc+19TBTyU/G7ocYv
QqvQXn9cERmebPqomXfrIqK+TLcH3PC+ft3taisOiQI53IGGkkCMX9S1oAS6
wQRU51GNsbhDic8jq9C457ob6E1vzbQ49Cgn8YUWdD9bRnnwRpiir1qtwy4d
sDcSBDuGF5+p7mQUxQigMWAVx5mWxaPKGHDx/Jpd2zHvBw6YrVoM1s9SH26u
XatWl3vgBB2NiFv1tvWvPJt8FWx/4PUM5lY9Psw1KQcu7jcJA5S1qaV+LUMV
wVT4ExlQIHE6wvrTItTRfqCPRm6lY5QgXJOT7cpKw1whLfi6KpVtqkYCuPwN
ba/0xWHDO4+M5hZeBdbFgB2C1Px89VBP8zFp9o4W1S/YKTVniIgC5w3kFTU9
BMhJYQnpHfbvvkFzlsNGyZYpDqF4q+CnnVCMJQU6B5NDlgYo2Fx3ypVbBIoK
C8NzFHso2tuQFfv0LTpi49x2RpSCMztJRBC78jzA3HJfjMKLIYdC3QW82zhZ
QfNvKfKw7+df6Rs56ttoetb7rm46VErWYGghKjgNDxFbgAoYTXYUxpZ5aRBB
5a7Q/K5ZhOwC6FeGQPf0ruVzNfnDIvoMEzkh35b9AYHoYXRn7sz4X2Cn/q/m
sh23qhAylpXH0yX1q1nJfMCi+UUQSnCYGe8Qwb800zk6yR59z8S5DjKLpmRS
gmX5RvaqL6JHZYgf4lDOHGeysAok9V1CnPxGyJlKJcbhySogQLG2/cn+53OW
gn/gRjKaHellCfdrTcFIxmilE/BX3J2A9w/S5Sv236Fv7pAypVTTXaPk6CUO
2PqNLtqdcGcbpFoGwYojTlSe4j0vf7BsX8oQj5YzqqG2g8Cb4b2QLYYJNqM9
8wu2/x/cab41zHFXHeyQaYkIrI3HdokkVdroc8Pp6tAg/KYk0oPXO91E4Ndi
FQdgC/8qtJpEmlTDfMbXpGIQ1uRRfio8eqSyruuYX3An4DMpOAb/+ysp0ugJ
KE92d7korAJzJeYkzL4CZCPqzzYoXVsBETixJbavM9fyJ7pYa2o5h8KEIovW
B1KfZupqOjSNGISEgHR2obpihRXajL47P636Zr5PU+EFyp9H2kTXTRWYGEHR
ny5MT7ztUSnW6pnabR1Iq4OIKFqSSCHYiBkAZUxeIpz2Wb4M5GfmfxR1R4NW
OBAgrm2OLRBW5TshZ4py3re87Bz0SUv2Fr0oj3HEi6+VZr5ghBnwxMi0B0VG
kRvOMXDXi3Oe8+/Q4ZKoDflVbN3sr94kFozktSZKGAEgIHnf9oKLKoNjRXpG
eTwyxYEzKDEdzWG7SpHXY0aOSL7G1c6ZUXpxdBIKOg/cyvSzlSMIHs0J2R+b
h+rh0Q2/2gOUtvP4rplCJ5CS45PjhK82XJV8RRJvfAfCjzgAXW148fQRfOAF
aTI5bQ7UBCEKq/D06gyBCYByewrsMoMApzZnjS7NTBplN6ZPIy38F+BRVOFi
YgFc7qJ4ltVm8B6BTKpYTV+nCtcQZBy8cTEWnPRNVh3skTYnFVPuI7W3Mk4I
zDU4hWYXL5XD/wUU9rz4GjROKos9RJyrlMI0aMMadHzfNlpysZHvSP8wEZJ4
s00vMCG4FDypR1SuXCwt0wCGSX0gHdwmPZ7gHYUPFRWVmG86HQP7ja1Q/Jyv
je5ugbP9QoULVCPCqhYIPX5nRCyqpmeh/kXR47TT5pctdIDjLzFKn3DvwdV/
iYUYGYnIP0DfBdKoPI7hllD+B7UxomIZ0JZDiOElQdq5fmsiacQgB1X5Vk4A
9U7Oybx1GNI9HQPJWAvmkJ5ZYbVvwY/Ge9xbq+REZZ6h58AmJcUt1d0kwMOd
5yEhYB1jhsQufwhNX47id0Ujhp1x8FVDPvISrMnZXbFrMyHqAAHkxIsUJxhC
FKQPFyL0l3Vm6+SumlwaacLgsv1mA3hA//6yrcxeh+D06Uf4khFXttdihgZg
OuITrM9IclblywKiNJHsqCwLeUmDHbIes9k8DBQJuOtTQDMuWVlMIWsgLSAn
/5z7qd46fxOfNJRrS7LC9dOZTSGNY1/LKU8rVYmS3DYln6wUBtqliGLiWq0q
MrDgV/BdFHzu4UWTRWArUTJ7LIjP59qIFQIL+rbdKz5mvFazBp16D6CO5I4S
b9WzBaCnhMVGhowlv3CB/ps54bkE3m+B19hvwXLNU3zssKzipl0voEcDMAQ/
DrN1lm1bE7pMno3nUWupYUr65quNECmAUtW6v240I/DUko5Nbkwib9lMOCKf
Cb6ZPSLpWRlP8J66I16GToYJPwhLTun1YyA2dck0Zc6jV0HvZfjFPPw6kHOn
vAtgb5hlGD9neSyn46ajB2984tJDDz4aMT5lxDbKnGHr3PrFfU3IBx2j8X0N
niUfQNrzEg63IO7bQiSjAQHt5/FqYUW20D0zRlVbfyCMQFeChm2wBRVBjbYO
a/kMsXtokWAVWtp1CjchzIZRJtLx1ISF38X7QR8P8UafMwoLMPovPo1WWGCl
xAd4FuFqJgtb2aL3gQp0e5XQLPJK605rnc1DusYQHtNfy5NsOK3UMMHjRIc8
weLncQV6mwCHZzORJVhjmoUM3Ktxu7gEVgovOdknbIOtw54w5qV0tWz7wZV2
qFpVsIezsDmB7MFpdgM/DQxXBSVqQ8MeFVO22EkySPbUfAuTcAa8BETLbFQ8
QIMPEmeO/XURPcjqakhwp4zEA12BJZX+w27Vy7WpKFOvM/TZXegMABW29Bb9
TAWO8P/IXUwGgSXzQ9Q7eYf/w0HJHOClfrWkJbqSFdUK25btCObh4Gvxjvp9
kofdwLXjOcRKCtpu4Dli4Z+zexk+//OP4piITGaMr5hW/4xpN8mS+aaw7Znc
OKbnsEBU1WVDq7iVZTGwfLJnYwFCnrkcRjUcF0YCmOKxa5K03YGtq7GALGKT
2LkE6s3QIk8qU4DLyU2v96F1ZZH8NLQWJmGQcJx2IXskry2n7o+aTPu8qzUL
CsGG3Gh7hbO4HRlVo7tTeQDFnXte64MvgFVXQDoO8omYkqItvlWzF0KJvZxU
TKCFy2PwYpe1Ximnmce25DEHDh3Uyp+pf9MDB/vLiP3IjpcQjvKKd/riDMNU
w56L/dpKkzazs6VNjn+32Uj37S8/AgIQ2wHaohDAvjmMMus0j9Wlwjqh86G/
b9cZEKNX4JvjAfl7CNcpVCIrI34AyoYnf334aiAFO2SPX8DyrHEpW3uzMv9o
Yh+urwgv8JSKkQemcVeFoB8CiEPURWx6OP5G4ZsMHMtcUZ3YYF9coJiB3WwV
/SwQeKEfFaMiMhiWjQ66IJdeF6wWQXXdBfnb9KwO4XjwsAiW2ACJXLmzdt8X
MspRlzDMh6VZMoX7FccAhOh4Cqup1tPORiyjWhvTowzyNRBURoLqLEBuxsij
s+/2oXOkAIoTsbXSo3T7v9WeIfnL+G5yM5RGE4HEX+zle5KfTomFLdUddQlG
15Y3C3Ux5GgfxxA6F46MLeNYkB0iFcDIjblLJnt8uKT3NC38Msp2icku3EIE
1ZeRSU2YNiUgdScjpf4nM6BTseu6ViBpz/SmN+CPXcU7B7BHXmEDKQ7yizTq
yKpR05K14Db8tACWryrjXthoBMRONGB6mkuW0y2+ij70/ppijyTl92SWIx7Y
NzSS4ORF5O2WryGDBN+KntkIZTviifQigBIHrfO5g4PxwzIX+Zy0EiUFwJTW
uvAipdFpZyo4BcsuZlKE0idjyTgSIOFWllfZ5G4d0kKWcPwRapdpJU3xehH4
EuRW2olBats635vd/7+Maj+3fg/Frw629xDMt0R2ApysNS02iDBkPhpbeLcw
hJIB7cZCok5Q70QiuwNJUBoYXDpOnVe33exKKkzEzNdOF2QsZe1rNDxxoZCu
uXElycoxdRxDqfvTi3gwQHytLWvWqpLSS+h0BeiaXVzhicfJcjw0ZOnknC3U
PljKcXAlzpqVc/EbPhZDeUT81H6UJ3zJAMvGRygVVKIIN5sjI6VbV2PKPrF7
cO4ZQAACKDUsjcIDg+rTFgtI9HGftzk3LOppNSlIMnr2XMRq+PmnHWUF/V1v
2dywZhgoDJt4bYZ2fntoInUekBHrz8pJIXSFWF0rUOfcLqHE8UrncZucXZdw
tIf7VYryX0hvPKt+Dq3UElPJh/DpFC40A9tPgy+OFbGujxdi+0UJTGiRmeh5
mBPyiRiESOmLBoIKhGq++xASFHqCXHb0AOqa56FVs/sOs/677neus8ekNF2d
L/um4vBY0D794c2A/CSUNNa112vT4i+UjFqM95pJGVyKSVaaJrE52l8p+XYV
ExEeJLH0bSGeUGCiB8kEBQx6BMofCkytXzp3eZKn6rxTUxngC47EQuz/yXb7
ua5+WYlTwcPLZnexR1rB9FYbpCXZM4KaMWwtXZ4pz7gtqVYPlV/fqojvvEE8
9x7qrsTS6KZcLqdRPZp4q5PJ8ItgYMm5D6MyN5/bUTkUW4iE4qBKaSEkh+Lu
+1Pdp5giaog92CTp9rBwdmmaZ3VbaJLXXtRMQocx+j3VTxGiqbMTFIxWeAxG
r0WajZSRd+Z1TTBKquO2gIlLjO3R0WfCkl7zk8QsDIOOWitz9BKkVnbgCX4M
jzb2EAu6l8CJ3ns2h2vCl4+NnTVUtXMUm788ZPozygTp5z6I07FmWtt/jsdc
hGaAPqcXyg7g4krCCgBEgbrMFlVzG0pnm1R6FfCM79pwW/Vfnoi3HScotTmk
5a6yxP+maOFuu+HKd9Ta8Kqo2PNctq3du+odXVcPYUkR6w9P8NNo26kehdfs
P8Nhowxi2SvHAi4tEENCUd0D6yMd6u3LKExveH5adLaN4AMyCxGlUaVQTJqV
p6TJP+XRChfrPoMgsP92YO0cjCDubnJMLSU5UVLXXi3FZs6B/CSzlbt6bqWi
Qz9HMN6yCjfNirrXDGSz/3GotcX2SJz94+mOpNQU47/quR8c0Zj/bVaqloTg
G1ky+HN0GK4M6gmITb/SFZus/mjdq+H4kBl5txcnx1hI62SUxMEmCUW/ovPk
SL47bWpwvPqqBLbPN6iaET3oX1eMsN4VNOmCdN1CX4jbRT6pQtnLcH4m+h8K
O5zK1/JN74xNQtCecSs6hlBqjg5DmKCyenfFUtG88UV+eFBw44OtdiYH9wFD
oPwZ7bw2fyagaftc4f6wYkehL6jh/eJVJVPfeTZsNnnBh5ZBbB/so6oeqcEw
TBzmZdBnKbxhyDpQfYX0BGstgZN+sfJZnWzQK8+HS0Wu+TFM6wpuZCPmeM1R
QS8DnvgvsJkZQyA53osCsr1FUJf1Fs6QHZ8YDSTjPuXq+HG6a7eb4lmqZCnL
YHrJXvHno+4Ddl6JYNtMuErZwLfohrgPaWizlHQWNJg3PvRq7YB3e1NZvyXz
jiZWU4iNgKPa+SZTfYGZ0cKfxfQ8h1Okt2OxGEu61cPUlbyBURt/OogQ+a8Y
eBIKShiPuUh6IE19Fw21FOKU4Ua/E75KVzdjGcSUeCu6fIQxdA1zrhyVB6NH
SCdM/JaN6ww26+Vw8c6iamI9IrHoZbBrbElOsyv9Jr873J0sZGYJ5ueBXC0C
T0InMs839l+cDChpPHDxXl8LNpD8YTdEe+f0N5dz0uTW4b5irlamcNVNTqwO
69W0K2IPqM00gPXCX3J+qNWZmDwlEXkzk98S4lTTTiOctgMNClQNC0Zdq/Nd
GiyhJwDUcCYp3Ywc7aEtmdot61SPV14UCwp7o4lU4eb4QDUOYByVD20rvVQb
bI+euqBXMkVnfp+8FYMUJxVxIFOAi+V5BkXMgA2EBeifA+5D4jUDuaCHBEx/
q3ikweo4xy57gdlWaxWJ30pLhfnjeThTuliQxN0lGOhI4xXXnko/QvCb9dgF
uhM3kTim8LJM5d/46eDUVdRIGarvF5EXZLQJwJBlMACQH6ySVX5WvjE62Hwe
r5QYy72TptOWgY5/tsmoNfsGExkpcXBu4lHymBVErBetXRACuuNzydemSA47
W75X6yBFcU4I4j31jdznP9F0fnH6LsKfowDwJcbLExxhHzvMNY1q3tRzKLEy
fNyBD8Mt5cWGX7LQ/gOdxSt7tV0zQcZamfF0C7aGrVKSUVfzwApl74+Om2uc
SMKbgmceEkcu2RGzJwVH6X0WPR88PQasYdagGFitZkvvOcP9GB0Dg0cFNRGB
WljVdpH3jyhRITzJPWhZbHpX94zv+TyxpRTRQYeFQ7Q/bTuOIrqpDL14Sji9
Cm/w2I97+WxR7PdlkxL+l8cQUC+fDf8EgccwZvT5IWOPE/xWVBJNf1ZiLAD/
a798n0eMWeErJrFHiroDHQ4jyTeA9dxo7FakIPb1Vu1y+39JWkcxA6bJKhF8
/Z6OTaovN9KunIOxtVrB3DBCM4XZP2FcfZsOHq1hFW0pmYaH8RrgdyP+bfgC
vjtgdM10ClUhiLkHkw5UddTVkaahjjDqcjibEc3uTO47+2NHgSPpy57VBvsJ
jhx3x7oNgGIvCZsxHimpddz4rVBV0IuBm6Qh9gYR1mwvHkkqs+OAdjYIS22T
NEly25jyzacZkynB5iGe3eRn9h+63BfAXKGVLCIwdyeKeMrne8qQxBoVtvdZ
eui084JSY/58rZI86qHkIApdWoeKUrwAo77CqWevoFkGa+L8wAIAq70icBfK
JFe8OXAscf5hW7mJ8wGNIsRSvSkEAIGXt8C7XMhssnhbk5tfBTfF6ZuLBll+
cGs08WbOq9tnQqbt3FOAzXKHm7Wo9EPV+whZSoiMStcQOXMyHpOGHSSEyRgO
Np9isV0c/wzewElt6fM6ZnIf6Tkli3PFLr36bZ1ZqzgMXzDeIqcDBcow8bRa
hvkG9N9qPjHYxNhYs/A8gf1jdJxbJnvCv4k5fYoUJAyAsA4GO3sRhc3N8or0
bcBbF43ba9e4OpUexQ3thgqGYJ060k9S2USABHwfm4RXzEXkbTKaofCJ5nwQ
rjxhRCd2tbxfDjUwEEHTRDHgOicNHO3HegMQnRI2p8HhAiFKUxSMvtc09ou7
AKHo7U0s+e2EERBd9WfeVk1MVXSvuTnRh1q8AR8/uVBqHw1vB59Yx21l5qry
Q2C9Hk5wupB6KQzfJeG4Q8vftX0CnkCWXXeEs/Om8ssKG59I9oRkM1MHs/1P
jOTY6JupGHaxVb/48kDqDcdTbouAwKD9jFu61ZGb6I7fHaQJTTFECnJ9s3ex
DaDJPz495xkMIoMttJWd/c27ap2ZCZBcACDWPcK8FUtyQF7+rv286OT8/Bm/
Yc6SsSCXatucBdVCWhKomeQ6pdKoIvw/806AYZLi+ekrQGpD6CCX5d8x7Bk0
xcVTXtp8tGzg+LUrXYnSGKh4TQfbqt9VOX7jQUa4toTsZzZjdyg4OaGDfE7W
AE41ujqXZNhu58Dqz42LnxusCB3lNY4v9noXk4Csxq54kLA40RLZ+Sc9O3sF
ksj/NdHjy9v1gaM0e0TSGdVX3KG6B138hTVcdnbIJw3quboQLmGPa8rFmcNp
rrj/1GaHpQxXV0DzwvYYzU08m6uvcivb+f8R9Pk1pxFaFporG2PLXOMFkU2G
YJ/2bNsAvK+tD8NwDvKEHPRHNbFOEm/bfJsjoujZydXQju5gQjby7yinLKrX
qUT6Ea6lo0PflD4NjtU/A44gGjLN9uNAbjX6ntWvLGvEFtUXglAmKuiKnDPm
mUvNoNSdO3oeYQmenNQjP23voxv2PzqVLv+i3YB5Okz7Juud+M4BwoaWecNd
UXC2E1hx8uNsy0lW1RnIl757dRf8bwauWwiEHmn35GE4ahMa6+/1XpHYtnbq
8lyzfd9MK61EiPRfsamWyEhp2TDyzsx7YiSYW0uaY7D7OMDWuV7W1q4J3IUJ
MXwfLzUAGklvyzIBwgQZseapWIbGKEKseAY1572Hd6rSG2nuolaMJuTXwKTM
Dsd4HcW3r+4GxMEkPxh2GxcvrO3YTJgJAq26gje4NO3cfDtbfsVa+ok0QUZC
8GScpDNMFqZSyNGISqILq9JrhjO0ghMnprA7hwiqA1AihsUtf3YlhRN6pDA1
rxp3V14EkuHbGntuY4rWZWCW10sU0slNCYWslgXu9NjQYja0IP+xXlTxYCG4
Dv8Zjs/NJz4iv9XYJ723FDn2eC6+ob1RL/iErrxof5IJjmp6SCFuXosCI9u2
qWqdd5lN22XGq+jeNZVw4U86BRI1USs9VAIgtyggXMdYSc6p7bAXEtjwzeiZ
8ePu8nkypHF31u2QQO5FfRyV97Mbne0PlGCE8oVZ/bBnqxpXSUC8lyZO96Ox
Hq6mYP5zeruEd0Aolej5HlbnTa2eRZ8stIpHUqQ4qvjf3uFNRD9vGcSQVA6C
ytY+cz7AYwttl6AwXqOm4b1TRxJzScUKQpuPop4r7sOkKFeSgLwT5AgxaXgw
9dCfmAK8Rg58SNTz4ZeOJpn82D0TYaFfJQJJj68Mm+0eURnWPZpjMNWsqY65
bySL4aShovaLMymbXO30X5kTlTuaUTS709fv/PODvN/9vuH10rw9AbVveEC7
ZcZp9tSk/UpQL0vW24sytmlyALRGGQl/J6Jjam+fpSaJo6DxWvpk8MWIacsC
A4gstm0i6rYQLGk40CN47PUVqtuyLQa7vZiQjjQSy1LIcLNHJqYSlmoy4GLm
nwtN/oifTJ81zXRCz9lDILKp3mYPPCeU/hyYTEmrgmOC/Mxl5U2RT0o1eDyv
l3KDVa5IoFsf2dFOJZ245pziCRkBukTCDMMjaLJJdJAFvTVvM3XyouZLKzXI
bGJq4Hki8EQyS96YtCHcceyZBr0MXefQJaa9IPHiZ973tmPjkuy3sC3uP0/g
CwudETJOwjHFG//ba3sBvLKja++AeOHdKzGOdB4cXrEDE+6rH1pI19bKj03T
o9AiSJYYG125xO1BMJhN3JiesahMREexgINGZ/lX4m4w72x9sz+ZrxBfP9m4
pxFjCO1ze2OPtVRYk72OynBVj31Uh0cbJh8DwHuQ5q3P5oSBdm7Tb30Db1fU
OoCkPvgpopTF+HvHL4tmi2q08MO5xBSp0Flya2nkq2C8uabGy9fm+8yZLvcj
UJMOQ9ubK7PfbBtNByRKWoKxgSukOe2hOMkrx+pDP5+0pYLAbvWce9JK6Fj+
SLwptSRKETyh3xW+WEBcbfa93NYxSRwm7obRsHKZHpc7J0GFuKVfR5sOZEFL
CvgNDSd+clqQHq1uF83N1DFiD3E+k6gF+fxeny5yJwqwHosYc/w1Yg3it/xN
iac2kHie+fyhGzQWJ5uzk0Ai4TIDYAsYnAwd5rBdOPJdTMDXAAWM82NVngYs
FhqQ5EMjxR1ECYKGnVOHPXZ1yaZ7U92HhWFfj3PsBKMtII1P0xHqv0TdO1Yh
EKXmvo2sfuyKIOtjRM99DKVPLkFKe9XErEg140PLCDy/Z5kWXGhWUPZrEwdw
1SGyy8EwUj9j/mOIyNiAze2wzv4pNg4koksp1Lgetkcx3N5222yIEJa7D+bF
cQPIvGzyHsvS6tIeYbQiPjBKGwsqOQnKl7ODDH9b12LeUQ15xZd0qBZzfXyn
fDOdXmcEcNS4m/ftcH8Em4863Y07+pHOAl9cy6XcN+sNFdkiZftjghaN2KyS
YpWvmDb/5zcI1+40HtYrDvcg15NjqeoLZNKEnXPS2pKnvDLhEP//KZU/H9+S
6MDwOcflb0hdOzFzX35xwH/+THBjANllgcXm/NXgorvC+NRVjL4nstG079xg
iALqentHq5IJDshyFD0an8MRPSqzPpYyWjmqNkCrCCGMTg0awiDAsx0q+f+y
HJywqybRbAk5Zd85BAatYzGFkoE4YbIkRnPVHxu0IzuDDzYWTOcoFAEIXgQ9
Z5QqEwp9ZsHlQfWbRd7rmAqzve5fAl4+20mj7HwNAE9C8UNr85tVwcdR/KEI
J0TRO8UmK2K0FxV7kyvPjFGsIjxzRZ/vEjo4dPDUzRKp7f0E8GsKb2I3nwxp
/6i9YYILZbCLKyM3AJZBwyjKw9c4VaKJIgi7OM5fmdb/r+4ooxKry5MFUyy5
WBwhjqt52VDisKQkgjoAIIo7efonGhAz3Gy0oIPoGmQC4sFYcsvw1/s0RcKe
St12dnTz1M7uKS9UXgxzE/hiUSwx3geFQFP1i45a7Yzg9PfpSQoCaWWftNof
Zno/q1svfC2A6KTglFZbpKEQIqTnMinaXBg987FKzFRXPmL3Sby90WLo7kSJ
2QAJC8oi285kKxO1lZVOe5pPpoJHhlDaGqBlz/qcbyKeUgcYBEpxJ0Gajoe/
uQ6JH9QoxBRHZVbo7JTxDbacU44CGxPzXgyLlyU9nPMmax5BNBx2izjnr+5y
f8BCXlpi8yNDkgGX8e3SmAQg2chxBp/fwkkQLjSb11hmyuNg2O9kdeoc+Zo0
Vv0f11CL6pUDd4/1Ej3FMO64njJEUsdJeDL3SL025V6mknKN4zs/nXQNFD2V
Db5V7ovx2VKyvJvFkGUxwk24ei4RjqLRDzT54jDQa6vi0JhHyGNQAUWBOVOp
Oi7YK3ofNTZfC4nX1XT/3/UclciTyRQWW64bIHqh4AJiaX79GNqOB/laA6UL
/+x9EOAH8OkKLuYQmLCpFv7M6GEBDwzPVQRJTJaIE0fGipGd2XKSBH78EDMU
zpmiIz/qNhsgVYk1CT++Px+5weBamA2IjJ78tEbxG/7n6ChHqDdUvKCDug5S
+mam6+HTQL23p8j/1My4FH4BErJZ0hfXYhi/PShaOnpsnAW7N0a1+et7hD2V
Ww/6yha3ZLzFnYq+Z4BsB/ejxjsHZ0/JXZgzDxZQs9uJdpWI0QSVJ8ftNqye
0Hr/GGvJnm/+AjQFSv1+8phjYfebK/kicXgjC6EROseNFXOkbwfT5aFXRhH3
uScJFFm5Djvy/eo+CEUQJvKQ/abQP3BdBk1jP6joCe526XE0rKos/uUSR4Zy
PnpylRbj/7rE4vCVfgPwgKDPC8iXcSOkvUHKV015efP2AzwzMuQzTVRL5bp5
bXdGcnDiGiLqCA3Hmi1ykKpBHOmyrCJXS5wb6W+qpEZFVlHTgwn83b3hsPnF
mGuDcjVoJUg7mpp3eeG+zQ6+GB6TnbdFSh80h8d2NTyt9215YUGxUT0gABAr
DauKR5rUH3uqgvAEDWjUxwaQ98hMduTC4rFedPizXEsYvRIeF/EaoawA7Qgi
h+RBWDDDlHeYzRJvuf4LMSAiUwOekEiRJp3n+7RxXviPUkOkuizeNlI9YQyg
RKzQ8IQooaKqKpNWZwJ2JeRR4wBaq0W8rMqBAoGtJHut/6kqOGIuTzzcVmLK
oXz+fZkejbh7GTrhWvKE9Cngwm1YEOSKsD+4luLywVOKMlU6R3QpmowpaU6W
GRRAIBY8FBRBaE1qew2K9JSQ0IJu6rXFs16hmsTIusN0igIlc9McZFyZep1p
rXuhDOOMWYdW501IflBl/os6BYwQ29YSdWKLvuc/j4KEfIjeFbNyD8w4Gnd2
J0cZ2K+P7B4zLjRqGbd1akFu/E5wt4INJdBjS/7JojGmIZbLtwnoi1VdJFzO
Ut6TKAE4bWiod+U0azeD4s80qmiCb8AfUm32M3K0QdPTPDrgpKi6tZDqLiGt
jxeVsBX1uWNFe+Yo4Od4Hbs/NoP1CI93B2iZlsYAUAIudtOTIVXKJ2fhlnud
gQYC9JJvHppksdTSaZLWiAOxAMr+NKygrHBD6QAlmu8x0cGYwPXRyzYQQ/iW
B3IPL+J0q5FxJZMqNefY9nY5536EkJ56ZjK4YTbPzNZJE5AR/yIhGWmGaS06
bgMSRcG1ETNkEE1LVhOFHltal6Xh+cPNP+ujr+yIfigB+RAcEWOfTi53cDUM
NQYXzokrtxvUw+v0rcuMbhVKcsNzSMtHB27FsFDVLH6o+C/5xZQiC4CH4S0z
83q97zqsKeGWnLeJfZoqfhIXzKfD/s5hyhvGJNqAg7MGsc0pgW5qaYux1Z0M
IQsNypPPD/SoV66330Lvo8vnlzi7M3tM4XyHb3OSPCKNqZdAqQlqcamWGKod
QD4rYbbW+TttPtw6C5ZpMWtopSZf5+u9x7QBFi0VuNtakCiAudsba/aMGVZ0
fLGMEp+sqbv143O4vGdWyR0fOgKZU8j5YdUAquZ2tfoV+plkg/UR/5GYO8cv
0SdsDcIjhz5uWfmF0bKAMDO0DkGPnC7AqKa+UFP+JiKI3MLq1cNxXkNc+dtE
gW9ljdlZV0pe1x/M3q6PdhgGNvKmtmJB9Mu2B8wrWX1w6nRRlhP+/DTk4p7e
0V3E2UAqj8e1Jua7fmEK0usYhsYvWv0+AF49rXU9gMrGsZQplwKm24bjhe7C
h6CzZhqWvLU/SZckugDLgM7upVAtavv4BT4QJicnFDIZc1SXFnB58Py2enQU
NLJNNOfyTuoR5YuCUP/VYGo3kV7kqrUYkuPyYeFqfUbom4AN17dnKj0z2TFl
IRBYYVkSkhrMP4imR8PWhEBdkrWrs45IwupcH0oiR+5UAonU3DrIqr/kNhFy
rPJIEUpkB6ISQjknHrwLq6PZS6RgrtgjMisYINhB9AXjJwjAFtjd+SYR5wfF
PrPBjquV5AyEsrcc9uzpjCgl++pDV3azkQWpO/wjoOLhC6cTNEJ6kXqPncWl
giptVSQx0VunLRnCdktbk4pEJTCaBr0LY5qZzXE4aq+fIEo7Hk0tlI7H2YBi
yaCh7IfJvZMO6wfWBlgWi2q3acgSuex9qMJgRPTpyfGjhscvC6/7ZOdUtdfD
ktFg3PVTxPaC3p8D6Cd9uXmVHSVfP6KB306aGyHgoBiQBze8GzvcWhZ2d3rz
jJIoK39cgXz+x8RerCCJe9z8HNwkzN3t5iBRil2DU+DT6aLjk8NdDmqA5too
k3iOUWHneQ/cHA7jiOScPlZfDOfTq+3O5faUVknzGVy4+izASdu8ROWQAxPs
kcfJ8dEdALEB6DFjatTYrgoO7akBDJ1NCobNdUFcorfwiKeuLwqEqxOboFOb
10Ae3z8HHl9NG2GxJWpLgK+4XBj5jMblyyfrkUe9ObbBWkPD7eS4vd4Tz56V
QVw35pWfwTSN8fw21To5p73dWVu4dGYf3XyHMNNk52uD58LsTxEP2q0nOj4p
XTGwVh5taRGeMBg7nXJ7C8jJdKhYe0gcN0+EYEWfqEp7SmisN2zCJhAr4oc8
yrpEciNz0BDSNq4PbSDQ5UXkAxUq8eVZGXWIi4MfNKjyf69FdYnq6pvkzEhB
vrf9FYvon8dt5VDKpS2B32aHTF5HABLTkpl+urx2lebMfAahAl1SYE0xjvfS
D3pPpZZSRwvByyxlGYX0jHIyOX71wvzyg3Xqr9dhOuE92ZMfHtaogn8lfTRn
puhdD2oMS/ipY7Z6Byw/CqsQ2Ghi2haxqXc2uH0PuTC5f2TSB//xE4tEKzmW
459pqQSoDF/v44kmYCjT8ibQmwF04Gf1dDEG4Km9ySYFLHD1sWOusn4JovQ5
kPCJEFJ1ZS+QpQ/VOlN/KVpVVhfZeYjRpdhKZD6BmhB9yqUxW98XmDcOwK8Y
70qPBTKLU+JHJy9qIyv1ET+cz3pflCAA3ly3ZEN6Aylsa6OIupFtm7UfqKG1
c7YGX6G5MFcQLF5lXIm960aE9vhFUhN1Za7BaOFK+zYajsWd8mgH6OgEgt7s
ItEWL7pngHRYYKblZrpNd2ISAodywVnrnCBmlalK/IbhTAVUU8GK9SGR1r+2
wqiKwS7c4TlPIweAUoMt717aSb/nQe+8MzqluIvgeZ2QT4aho3Ch6JKY7gf7
BDHa43KE/pEB9aqCcRI15Tgf36PfsjtFvt0SUA+X9yj/WSCfGFnInZtI1S2x
ygHvyvQV2VIFMhBqjnEKba9hl6ZbT7WSygG7b3UWQy+50HXM+AEFcnpv1Sfg
dKrSIPppVY1KpecRtEkKjAhRBZRih1njDJN22DEJxORg2Bgzo/UqO6kdGP+h
znW5x7+nM4IrnqjM2ooRJK5ddRjPskINfIGaEyJDEEs22EmJblHT0dlM52y1
9tW7brVRT5h8nUDAkEdXlq0hlVZm9dMkkTOHaqKsXWSl4FOa+9Zi8zq8M46S
v99qWIIU6U4aKXpcsgf2E1SrnRC2m9eGHW6lUNtu/N+vGl0Nd2b3QfbHqHRS
0qm7OHtms3TqinAadxAYwOkVh823nJVkOHU3KK1tSN7YGjLp/bcmW5MBLGWW
AFG8wNrk14m74HCm3noel876vlBeSw8ViXLSMsKZQEIRv8r5sXbXvOjF6VS7
fIJWBMeGsRA3Zrgk0SzDkoLXRwJwmJmJcwH+i6zmNrBOuAg4++NmqpB41P/i
I+3cknhoxaygeKwzRRZEhlcIUEr0gG+GD1eHThYDmSRohTTodrJzZvQFTtyt
mkOrm8S6DBn4YZnkLzQ1nl2UTiVUmkaRlBk1O3wlc1qcA6rka2lokXEBEq4r
YikZytvYd+ZBMzWOViMZEeFFnp3W4QMf2SFkk995lD1xgHiv7Ntbko/n0qK2
WMYRVnIqDbEqVKZZN3lVytUWPXW9W+RN/eG7P+two0+3MNKCmj3mpwXm1VZ+
MVpn4GdYVgNFQi0UfqSJqmzqvGmtx6oQYCtA2ZsDXkHrilD7Usnm9T2nb65C
MaTimUUAi13sAdJffamwASMI/ky/fDe1oykoFK/UhFhAzTTxQA1h6waEgiy/
eK8f7rfv5VYODNqj8hK2HXhsMJwJz7UFljMsoXJJ5bAQj2tzgDgQj3xTQIS0
Rt2nup7WEVSNwhLj2aKQJU0ddXIbOD5EeOxtjeMar66zPxBgMti+8tR4Kb6Y
9qUIDsptjjSjtjSOpxAsIsFBSP4uCVrY2wtq9L5vwh7dHgrMtlIgxXkRvqyO
cz7A3uZIhXxCZJtXjlijEUE0mhqiNGWfywdem8yVoW7S3RTVqMuE1FO3Mpsh
eimIvzfJW5sqWdQezwnAAmXW/gz3LDe4AXuqgeTL6TuHrI4HUk4nFrWrbdrd
CHcy1PJmuEVQ6xA+gATXh4NzHJfOnSPhb/HXkvBAoXKcRuTjQM9wneSPWeyK
MdNJSLwpj5arvlN2DIUplu1zWZfKILKYn0Qrh/Ih3fdoPCKLOpeMcMHlJRU/
I+RsFjZH+eTY7kvHMMy5MdFwLzTWGPTraKLN/3dTP/XC1H5C04ECpEDBleLF
7TZ/7vP9h+UNEBGM5gWQGOWisDpeXFBhpky9+W0/Yv3AZO42twYcUNHZjrqU
ie4lfVQHbGcMGQdAgNjgVtNmitdavznMl9HMJJy07HiQFXHgey/EfsptJZYY
/kVy7/t17iscu+ReAKysoFXT89mamq5KwP0oXANHOFHcPfmLbFONiA6TIRcm
B09T1IVovevm/OduI9zO/Tnu0dEmsLXPjl5tfyc0ChdlSAgj9RpdWVilhtmn
f8zSeiolPexiHrzfuXWtWil5XiakMp/3dVbKqu7+WffrUWZcmqeUx3/R3etW
gWhKzuj2mvx78MB9CqX6auPT4PTcgeqoKwh8UpBEwTqXpbd4JPrPQwSv7STp
NotUn17YxbxJ7/Oxuh6YiqP/glahGCnBZWFJqaGOXTwAWvD7FHXUf+s2RvkQ
eaxBaPVvYDrzpvAyRrWEm8LLx/t/LbxIwOKlLVpQSvqLF4XI79tpZ43ZJjTa
z5FR/yur/DWufkeuKZjMFDIJTxAPojpVytMV9kt2YGD7+XoUS39zv5UZcv2B
SBmyFTFPu+jIP+rZs/6A+CtXQk1j5tyRWzjbMezj5sQuYPZpakrDWxblYyxz
9EziRhgXTFT8adxkpWK6RADvPiqfF2fozLL5AcI72QGWrH+j/PBMqbKQ90aO
/UXBPruaAFMmd99pXTP9J0rPnV8U7QQeafvzFeXDKyQ+ydFp0qd2OWV/ZMER
MSdfQ0xayToyDn7Ygpma4eL1HFUZTiE5VtVy+Iv1o+dhdAuVwqyLVF5r+Scn
lC5tYuihnoD/Z3tPQqMKAgFn90mKbJt2p2owPu66PHrnWCyJeP12AwPLj4jY
s6V6jJ7nyx/fA0nI0quyxn8/eQeJ0dDCpT6R6OHXtG6hx47ssTVaYvNx3Npf
hXZGNvPe2HdnnrETjv8g7oWFmlTmxbYQqpQFanNs5fLry32L5sQyOienO5z8
Ty4+iOgiFKPdrkB/4LERU8Ro5ld5VTYfPlhIoPiyiQwYwRi4+uXsdVaQTOqd
ImJLpUrBzX012J2BiKnpJBYdDG7ooypuT5zmQpYjSvxdh8tUe5MIU4KwrEop
Z1+5NsFSVpJ4AUk8nSTbGWMg4ZKq/upwxmQ6Op89k47Va6SHK5vPbYCTMu+g
bkxMXAk7NPkNAkCSSbcFcrxUPzyRWn+gR4c1hKznSCpi7I6/0t1nuzG2gDCG
J06RsTgSjWs56I2gar/9V1FuKSNDHFs40rx4lq7Q36dDHzMN6hF9fL1hoeza
59vzLfV6t0oR9GATF1j7KswUH/rEQcJOZ7V0C5oWe8TjWoSG3h/uIT8W6mUf
j1w+rz+5xWAh8nwU/MX00jTFUtqQV9R7aWHjzS8jngC4kKbnBWqO3ziQ4GGE
Wxzw+YWF/T6XbclGgrl1d5NEtlpklYHg1e38aAbWsOINDysBDosGqn2BtP9w
EOOa9snURlOytrN8y351kHt+y5US5YS8aZkN2dLzYOM5mEINm+RpB4lKDOsV
2BdOGsBmr7w1I+ugwS0HG6KO7yG9RfxCvcNIQEziCecu8+tgRzidIoAincVI
7OhadKZPyJD99uylaVh7PLLZbOPvup8qubTCaYRkYBgUGeYt/Op4IzX5Nirj
ztfPalUO2DegXIbbjGlV3SIaEJeitssIgsMHAMqYQ3CjEQ2mNuyDSaIwXtLL
qaxPOz4ODRUi/+ehmAEofPrLYt/WZlmCFRChIR7hVZzSX7+qipjY+M6fA2ch
5XkJH5vRYZ7wNSfcH9J7N0LdwnGwLn4QY+NBfPqnm3TV8akk9URPkE+ZNBdE
LgAGWlK7e2jxed2Vee4rlug9T9GbhXM58QiY4Zp6ECv2Gt9kWzqCal4IyK44
AwPL3T/oVBS+qDPLid2UPF4z8D4/PuCjo7SQe/mSXfTrNskzF5Nio1E/g4kp
q+2ejleSADBAsQ0oPR+jMP9de4bOf3uaWciMd1qfJwWz5I6GQeZjjv2veLpN
drr62UiAaGRvzCmXA0ehz7ir2lq97dABT8ib9rPXs27fcqEHQiF4Zj0LoCkN
SLjxpqRkSSg6d90gWFyGW1K165BESTdMIMJjeVyopix0AhTm/ZD6TVP9TSPN
Qt1Q4vPkkDWZKUMh1+AEzQVqpDPA9p586EtCUWe7bYGnDZ0Felu8vltpcGFj
/cJcFxSZoh/Cz6Z6GNP0KtzpjVM2lxVf7ieAl4428gHRonllgt/zjGZ7vHpg
r4IasZkm0QwqyY+bjFR0xm4Qp9DWEMnZocbHLiuV709ZbYGBbPTEmXkVcZGM
afolzk2EgRpwkDFxrhKbCiswp7Cm9fmggUh5KFs/NKKc8w0+UyIHQ81nwYBH
2MVAWMU2uKokRwjJi1F2RYRsTBhUhcgY7i6TH0yWrR+kZvCEUIxy2YHXMtCR
j2FWGC6ZPr8vIzfhFSDuweM/DoC0TFdFjsDK1+J8bG2oD+Jo7mWe1bSrWyjR
M4CF8RS28lqI1NfIPOVdPj9amfyHvz2+2XPTDTiUnOX64wnjHgJfjFtYcMZT
XR5U4XcZHkT8/QKOCOupzgp/NYncnpyPTZ7UjFjNXAQPxmCR/EVMe6MGlCzs
kY+Bf4Su8Xv5eFPKSCwRQ2GBOME6cG0CBOjzLsZliuMaC8pVddG68Gqo6Z7V
JlpHYdIZX63Wu6zONIp0m1ViRi+tSAFrxw91TBVg3oPmDVeyAucKlMZ8YLGM
SyoBGjsiy/QzS2LtTx1bu41P7giKzCfKHW63h/KAEy52QueV38xauQj9sc7T
QxZAqCSbe1kDlOKjDbXc5pUUXpopVBOdgeuccMn1BFWevfpWAKclK1XFUCys
/ClwAFBVCTNs2FB0OQRI9cmVNDhW/zsYWzZSFQp/AQLtlJF96upDh+wFWMCV
GPDnjG+lrB+tEzXgd2E0/iTl2zUoVVsLAZTX/viDLpPsOR83TR4764vkz9Zt
70Itiuv4CJVeXZDNruuBKaTH6i+KMU/0IXDY2Lw6y2vSpirwV5yHFE0j3iJ4
M/R6I9X1MzIYK6tbE2jCMAJwlKYWRqMBnVbkoI1A4kz57mpql5Si0vrnMn3z
LXSw60+Tz7dAzXrnFqNZexOqCpECfANZZ1ePCoOn1WysyCU4KB9JVRiiDhUz
y97cIQAJXz04cdlH09czUyEmzo8IU5ut6dwQeqPMcIy/kBtilCRwpPuLbWHG
st+gfKv/RNRfWZ1ZxQI5NvJAIeHZCHSVkPbC0jmNuv9YyjQ1hadtEl+3qqoE
KIVZLZCbR522bisItN5WV9OpfWTj4KieWOkuKeMb25V1hcLzAiRdKQgkqCP1
czlnJExUNBj6WX2e2w14HH41iUXBQPq2BFiDmMVi1vtEMba8ZmtdcAtorqHt
OU55vAIYFl+9wqXWzlOCfPrQpwcCFknnVNN1DEoxaK4H36FJNjCEqnNdkx4+
D+acPrqRFghEc2Zn4Kt8T2VA7FDMB5sy2IA+S+RGSFlmdZkiYHrfjxYSw515
jceyGnwVgDUFN4EVInUTrIxTMVbBZxU44lkrtCfU5e7ULXp3x2V3dLcf9tQb
xsEvp0cffWh4kKUhahH3mdlbrBAvPmY30s4mdzAzTKCFyqm/oeDmFKvAco4J
tPmnDdbLXilJFqPNfVKTHLtsbYhe2ws9s1P1/p3crChcgqQRUhzaT1uAvu5G
mPWMGVAyD0NoorxsSnvVvXhH47hhDPI8UdxUTYroqR3ZLoQRA1XriQgoDTC3
BBoNHM+NaJ5iETNzeL+oV3Y/REmMAE7/6BJOGaCd1JPM3UQd9SzKk8gtXFjW
nydFRPFdm8szvhxJCZcEiKoFRz4k6Czkr80juTm1B+86R6q4reVXNX3o7glm
sKpNTAX1uXR8R6gzuCinDDZG+lfZ25BqnvsiZ7lMNh2mnXf/nhUmcvUMzGMX
c61dIoDN3bqEIndsmh6DKkVBEAhigfagFw+HVd1/rW+icm8Ls5UPCTz5KlT0
KnmyPlJvmyJEUyJyW1GwW3RzlMcOHwn/WDA4PpsdEnA/3SGZTVwsERTU0f0Z
oxvZq1Oxk3C7NHvKJ2gNgEVbSGFw/nSLVkGW6qmpCr6XVOfpuinfEVnGsAKV
79iP6yVvg6kGTA1ktsVJKGIoPYer7oXOQJtAyTasee0AxLzvvm6UC9CD6p/n
a7eJ3Z+OBRhbZQcePJRaiKpkxUR8ENm5UUnWbTJO9wIMGXTGpfYR5ljv+RyC
Y9iCRu3rW2EX0lpmgBK9tXuXAI37ywKcQd/An44T73imFfH2PoU8O4Yxk25O
4XlFL9I/hiTfSzSpbYQlhhWjqjRNxQ0chBMw3umkLyyog0JIg6S5cmkOeOD9
GWw0MjXXaqbLRjIHnWlqRLpZS35hX8DhjRBnSYXfXo9Bfwe9PkfkDl5AfQt4
1Dwg3XBaRryl2Ajks4vteezKDQ1xclABTT7wLLVaS+iWqABt/0Ikw64xu+Qe
J76vHV0CczeKKsi2OONJsCkbHPxBhCGnRPoc5DYHD8YXUdLBw2rrJgQaZrg6
mxYC67uGV8/ykbHFS9dUFZ4qoGbmeSKavPwlUtv9o9rTBV/g24jfFRAZTj95
quvhEnHXEMzbzevt+56UJZ95AQC7CnfK51cwrJIxyGiODmq8zU1OXG7fyx1b
9uNjuSB16wClUxx2i+56ugqBTUFnGtVFpKQlzB/YEQt4+a4wMYy+8yRSOr+B
mWU4vtp5cT0gckfvrz79I0G7bUdC+1tw29Lsysl9wE+bESaMnAr7Nw2pYCzR
YDUQS3ym+rNB34Hlh0JUAxmqo+z/wbJp2MAGYbgOW/t/nlRbE9xn07cV3W/o
RxufezxjqtGLxYsN8MuvjPLqnaJtMzwwq/uI5eE8KqQS9uJloQnIUeZzy+Ky
kpNFMAayoWVnlTQo//XiQP2lHUPLdp4rlVRNx5vyvbvKwfR5JV36Ck5wSrE+
DWWIzRwp3GkeZ8dOd+j7qWBzlX0x2lzcENj+zrOwdXOnu6L8rc8zS3ndbcMR
M04VQEVZk/A5//tqOd2hEbe8+A0ek3FGSZlhDkf+kw63XrBagSqpXnnNBG4D
bjFqpVvjW7lGCsdquzUXuPPTkgeCygFsw9GLZm8IXxBcRfYGduNfE+ZyEui4
nZaKQjRjx6/amBJf7rNvimxIqHwsEpv0ncXTPwOTetnSeJa70uHJ2HyEzyAX
SJ2U2IMn8zNsSfIVEx0q+neOlbNPU5TTnIDQc5dlv9HDvHwfDQGqjluwqc12
e1xHrbJH/RxkeER9swtdPeKZN5ww4Hcn+ZDClxJFYvaS2aMqzdK7eeFNrojS
tWUiIlPcoaj9hoIdF9qsMRa4v2q8Fv8F78G3nmCOMUQdbWbQIhWIKvWy2l+x
RN9PgfJR/Hb4DgFPFwCq6nFzNhaJ49friJ6HDaDMuGOnDqICIBn+AKPW98I0
CJO6wJRgwn91Uulgtl5oWHSFD9KqH+fHcOCaLQ/fl+fV8hph5eGWoi4RopWA
/APt0nTknexq31loLN2jzE2nMaEJcINNYXWK+BukD6ZN79RPrtcV+4IYE6Wl
tAyg7VOAMIjMi5OHDalXDkGcr6U494PQzymWZiMMxydCKCcQP3jMN8fbCWTp
qiCeOiA12cZj3x1JdJxZ3L9qtSeeXPsvNls924BgdT8Hctq77heWrWMMa0gF
peUZHHcZ0o1xf6j7YgYHEJ+hevH4XRm/PM7xMI3OpiC8im038XyPOho2qXXU
EJSROwMqqtkc+g9vg0ridevYP2h+v8NRlK5F24u6s/Ie/nU7L2Y78zLbumW7
U/sgp3mUxMylD0AJEqmYz9BHdj6X5YknSgTjuFfUyx7ydbZjEtNT3y+iMjxb
X4YZv1mF3WRfvX9gcCrSwPW7DqSu1zhFxK1nxn0rfYjrUh1m+oPgzsxGssKA
aLQj75zG6L2vrySeskQzzctmMHA6uAZThhSzInXHH88DeT3jcsKvloBeZDpN
+Rv3ZUvXlCZLDlTncwQnJohG2dkaEcZgbxbeLFJA/c9QlOG3hZBelQ13ilLx
A4QLrN+U52JxsnnzPMmMmaKjHRa+YBMacidaimEME6YTJxUU08P7YzG89TEJ
uOkJFDesDULZ/DVc3nLrLBk77qsAaD47fUDNEO6Aaxc1B4/DE98mORgQpuEY
p6heTmteWRkPJFNUVot/tJ8rFi2lbzDxJZX+2ViUID3v26kKscc9Ye0qWQg0
Jnzn9FYbJ0OXMlMjMKejifq6LvQaeRYyH5TLIZQgmRni4//Zn86UpEI6Tb1/
PnfPOw/quyeSKfxj/gEr9o8LtXBMiHGaFRKZ6IhOZlMrYEuzV4nsyVFSeYtV
x5WDn3OQ8dafaupwSTMzlXJg3+jW0YrX9Rki2YmNF1kf2p96FKnZB+CxO3sk
sG0eNZxBvrOFs91INNCUkXn5Vpl+8zNQpJ8yv2RkibLwNJGMiZOSua7yQ0tq
5altl5FaZ4VVXEfxjeC2d78kjbcSpncCiXMeeAmrjMnn0m4UFwYAUUeSwxmn
rzGy5Nr733FIloZV/69Ut/oeucBAA/2pLF7wtFLkANWwY2ZJDnVAp3miABGk
0lxyieQs/PPBLeo06C+uKR3ULk5nYxnhrNmB3zLdDSU29f8ptCAnnuh43nU3
EBn/4ltEbl0QDY3H/hyjvaouglFODIWkWnoKLuGqAQFc6upUKQf213jcOgRp
a5WEYBpVjL5SfDT2IJCOd7JuQMzlH1wl0H33F2DtE9lhx8CDKU1JV9bBDAL0
TELIeWrwKjFGtU2/BV7iftGsgObZ2rFpaMTsgO39+eTd/SeUpJarCTdy+tB9
NfYYnZNVCYW/WINiBOkqOoBboogiUK7rziIIkESaXQT8drI89aDxFyDpOI8T
DO4GBmPtzEZotDiuZ68hVCaSoJ1q9JaMuyYarC2fUjfwmTDRW0DJLkP2+ohP
1tigcYQS1TlY2Vv9DJrgqq9q29bVaunIFiHXS37eKoSKW6mrs2UUA3AlyhPh
JAdqH2y1da1C1ji0t6x84jcCZyfBzywUfbopp1MJX9iT24YKogZbGyKa5hm9
DirFGNTgPwnvSFos2kb0OKCP5bVRqVR3vQ0jQ6Ub/c3jsqRmJ7oxIw9sDrqF
4oMER/f5BpwkeXymVfjkDcMp+wr/aRRnXzGMc3v4daflR4LnoLTcYNr87Rtp
MxN1VaPeHpTgNp0d/X34lI8aX8PKGV6ki6lLnedUAyfzrvyQy4wILACRqaUc
b2WnqqKLbBHjXdp4pn7n4oLU95KfZ/HBtsr18TvoE/OX4IehAxD9eaH5TVWF
JjAZNB097FqhyeQzJ+jDukpGgVvgmgBsfcJNSorba7fp2rlsOKkmtf+Fkc0O
n8XHUsQFj99gwqGmaN3dOeKJ/QHdBia5tr9vBG5dkP5pgjbKgR0yHqmuhaIq
HrsTVFIOFhXAmZ1JDeh5N0PXRAY9uDcUaY9RsfpxH68J0I0/3LkOqvSvCMKe
gsErciEfSJdbcdI7RlQT2wH+OuNOkwx2zySPs9fahiOFVUoFHZDOXgzr5i22
OELehNJu/KZlWjvvwicpp4ifeQn1tygQSzHk7qlsYXNtUGr2KZoBhoJ9c/Qy
QGSv02gsLlzGT53V4u6OS3prkp5YVnAMp+TsOGN64MOoWtPlF0rwTD3JnEe1
cZcqVUc9tW3AjmWbJ+e82wfTNP568UNJs6cYDsYekqu/NHRrWjfHeavVVroZ
1kGBDi+soqO/+CY1C/h9mFOaqHMnAdUXM/J7j/7FeVroG4VpfYTe9FMBR42G
1MNlA/El8bA/EyK7k8CTmkucSereaAYEU/BGxuMxA74kjinaNlSTKAtOLqPz
psGp/oHQ4STaj6BimrErv9ib6Mtc67RwrwiEzooWxwGI2Z1696p5r8Nwe5zB
0v6Z7APFmxTd4YMuQrGr5WE5rw0c1UDX5XGzsdE3k3GMRgLoHhpGZvbcSn0i
qqfIFYu3evHRNSK/v0eK8WJvyl3vZ1OWX8DUDd+3vcYgm/6NGs21No3s2Dba
/hfBQzqenioeorLhinyam/CufIDIa3882WvM/cVDogTmD2KBuFoxb/qmioQR
IQoWN7XNbP850enstud6jB8hK5NJ8hnUZSE5YYSHHElA7//nIU2FC1Wh3s7c
T8rSiQ3erWIp0ouBLMxxvTUiEKmwaei3jNGjJgM+JKlasaeKTIedWJWY4bJn
L4oRqXTslrYBKutl6b6Y3XLxlT4kvx1nvb/r8yqTSxpAQLdTXliQDZlFcJFK
rvEhbBsO3JKGOVDTR0Jv/v38oJ/xxXQvS2yYMHYBAw4HUmBt6P9wiDtpZXW7
nV489XkkHW/3iO80+Lea7X8SjLyxlczJ7Tpru5tHrGsbu7z/ikF4H/3QxCMZ
5lF2bwpR2Xt1aTIGqqVfE45esutE3H3VBypM++EU3DEf6kBz334av2SosItK
0wYKNyd37JouCNcenywFUUYeLyR0BWDt2DYnScvsHspD37tT7is89kbfxJsj
CdKpG53cBr/pT7/mZw/HVZEsyAMBJ127iVYwMQ7+lUajrRGKXlKv4FqgrT/W
ZTaOAiIKieUa0fbgdAUAH/zygH7rh/W+nO/tQ3AKI7fYIeGivjVZrCRWzTS6
989jYIQsVtPJ1t8Witig5JAOV5UD74lRyp0hQK9kxK7lcCQtqrNZox2W9Wuu
q8+WijfeX8q+PuYHIAojiD2Qwd90MkDQQSC/m+zvn96ZfnwWTz4Vp+uZcMgz
AFvdXL4pWCHiov7Wm9UsjTUc9lnPVg/wYFyhOWv5zzmneG4gJ5Cpi2CmIGVL
aAuWSnBBOYe1e9Guut8XnGIkoTj/0ToeMuaYBMfy+SL2s2WEJ43+j06FLXtA
ZnS02GrTQKxkTxnqCR/otJnRKsGaE54phXE9eg1Uvp7Xgeg1pA2OrO2KTKfh
LwlXTXZuMYVl3je9sE1tgWSq1S5Eit84JR0Ny0h2inh81MsLZeKm2AUqKlRt
xYyYXEW05shPOwBYmaRvgQBzk7TNdE3meJEDshn8/gE8NefdGAUjKdp1p9Zq
K4u74MBCKfyjqPkM0ezzMqzHqs3krVWcfaepLRNoKtDN0t1A5KSwxL0PymLv
BlAx/+Ld8U0+XLFURLk9ocbS0KfxRCokMWSyicxrItFcRP7kdKm0G9uWN1f2
Pz3F5eHAz9P4eHv2Uy4fCRwIJ4aSHEafJHQDjw4s4A/f29a/JVUQNasbaDwQ
hbW+pJGq6cVeftZRbC7WpCj9i7Ylj4xN9KCR4xbb5PVpks8U33wIRvVbEFky
ev8yXU6NNDVndH3CEhoONQHphmNOxiosSztThJ0ps3oDbmelv867dd8Ai016
Ey02NHl20scV25jGc/6twJyoTpFOC6A82p/7udPKloMyAcGvflYAC6rd18fJ
OhY3rP+MudKovW8Ofp8KoHYQzKeG/V2vjQpHkj/wPsy69KaLfHsCfDiAL6ik
JCLtVB1aH+tsPhWmbxg4AS9A76jZDGbC1fup7Je2c8wCNxHeP0YkZKHsYDLy
2eUZvsSTivwiyfoJF4ELEs/rWQ3wHQtPv4/qRawarxCKCWEIcbXp7llu/7yb
eB2UjZ3FMzj5anipOH6IljMx4FSr7Co0o+K8sxE6H/Xuc9j1+VfcCfFqyMpX
SecLKT3BlgexHjJJFAPpw38jFCR4jFjbvcAY06lsxQvRw3Py/cxchhU++SUx
4ql70j3xfDVsa+3UYK9ifQlCmk+yK1EaGcRNsfbOcLMZJ8ATYzXcyxQitd7k
BSOceGfkLUQe2rZ8a3RIPl87P/kKc3G5/hCDdwhnNEeWqHCgZOKTAtu0rK2h
vpg5MT6CFU7ScU/QMc11AMtI4FA08VXk0Uklwtr3wwp5lYzZRQMBOR9Eg0Py
epI/OR0NP+rQkDxryV/a8AaY8b6HKicYzFPu+eis0di45ITUBLbcaDUQabAh
c7aLsRi/Of5IGaGy13SRaufjYco4ZB3u/FTcv4JZbQV8uPUrdFCUlSXgpp9Q
Yd0qeNgMzDWyYTadsKaYtEHcvgMJLmEIRTBbY/Wy+MwDMomJ7SNWacwn9pgz
/TB4c4z9M49gR4BicSXxHCVRuq7kxgPEXrbnjODgj8jZ46cpG0pWADJQLPtn
VF0hV4LFsb9nYtQBVm8jLwMdLXOU8M/klYNOkd7lL1cqU80BSdPDtomhPq1k
52WYOy04UPYQtKnfZZQJgjg2OAM2R0c3LkASfBh6L9OGBeJ7h0MeJGUXUY+y
HHzJbRHk8tkS6k8kSKeKfkGkwDwq4k7m9akPExt+yz7BMEGyYdEwxtQwwMVV
417Mfk9OdUXir+dACbk9v640WDkQs5/5r7DntldPj2uOm6YpCYA6s9A4oOfZ
0Seo2L8ZtALX5bN/1jKwf/9TLd8luTx4UkkhtjULEQwRVbKYlxtkscCwQH35
H2qsme0sJFeaxtDL4N4uHkrCzRcD71RKmpeQTji3loA0b1EIrU/gCKT6sT8x
UKFunOkunCEeLvzZlEpXN6MF2VvbsqbuzBcdTEzVHJAZVy2sqIWXhRV66O7S
Xe6CWJT2X3x5XEm+enV5rx0Ie01xngBwHfEEImxckW/nZ6WiX1k/pLK9vaCW
M/ULWhNXC7DE2ppTngTHlr8jkuJdF45cER4RWCCGdQgxqS856QA97NE5kz/m
hhJFKWKHBShatELZHZUDnjzJ3Y+4VWaaUQZ0KlSGslpG2Dk8acGzYAIJYUvx
aqoiWpL0mFfMbMcr2xviqfD5Vc1GIz3eAmn3b/6LOMvuwUd2cuWmh5HwkZp9
t9wMhem9TTbx80R4pjB8eafjSgK9KV4O3V6gpY87xB8NAdHbnOOyk8z7qqNG
5tooCgpImzenBidfz9yovjdP6Pv43n4Ftuhs7O+pZy3y27hBKM1u22MnsaES
bkCV5Ht7V+Nr7QqaD+AHCjWnxWagM6G7Q5C2H3NWfPO4rGBf5MUjfxObyXiF
QFpTOhm9kGqB5/bhSF3SVkNlf0xepJNikJuoapfgmccPiIDJviJH2PE9fP78
A7wR545fMgIIbBkeIyxwWhFQz2o8lNd5JayFYGc76NtRpnk3sta0zvXyNL1P
1QMBdXHwLQzP+1I35nw22pjaK2s9iEMpZMVK99dSsTeTSCDbJIJq6E3XoXtv
GuHTUMNiNyp3je0/XC6zojqLUg8rwLc7I060bjBG3n2sPkcMav8s2nukD8zd
O3+r4UvbUAyHP1f8DvIqbIpSa5R6UmcG+bDTvveneG4ile1urO4nH608+jcH
ys8U7NWz8te4nYshBvAs0uSXJ5sIsNSzv00U/7PEiGz44jXux+FRMW+u96I0
PDKickI/w+RGS+vH7/n2QWePHDRo+vuTYMGrmE1QKkhb4bySCiNN4N/jwbOY
wDUvA1jaHniglPr0/hGhF2yiXZLAker2En5KoJU5ed+javXDz6cEL2PoD2H6
5LpYGDnLn8tbyKPek2c9F5MA0Nf2YItlSL5XYIGRk1lsIYfzGpp37Qci9C9V
NQGcVMXoXwS6zmHCkqRF0zKzGTlbug30xD5oMC2fUuuVt/vFQwZJ2Y542cT0
DxsHLpYSxU93J0kw0YS0uUSRRJOsSg7/UmZlj9fglpivvNujVu+d0estVKsh
qcVpLuCQEtYR3dk9kfUja6gbqftrl9lruGrhADnqTu4ZO8eAAKNVkslUAgwt
ajomp43gBtBeudVaOR2IvL9os9CTdKy7euLymroybEcFpeSMqmZP+HEAUUTF
1PP2Pwybv5apCWYQinvEwK+UZ/uWGWUB/17XJxmP1U8RK6+WWOdCEtC/oa7g
UHkRrE8YHnIftnMepoDVu7BMV8mFlhnU9SwAzaAEuQbLhFriojPQmqcsc7cg
ir2hAVJ0V5QVhIiWvz36fKhIstEUp37JbOz3TVucMuldlc1vIs00UNNz0JKX
NggwUDeyQl4MZDwC6C0hZOvULfViGtuQFA+2xLRA06pCOOXlGeGU9I0+B3Tk
OBu7xFlSSn3VDEn/w0iSRWFMQl+wp29/gOWv1TqS87tOFydImt0W8jOVXBru
BlK6nVccVVsKMZjf3c6by5exmv92dXVCE8gNrBiMNRGgUh+r6Ndh4naorgu0
GqInb+fZRqxQka5YdAXjz/AgNLOdyNqn1i30UcOj5L6kTRPGPyYC0PiinBmM
vehaLIwyFU0ph9zw81OsXNhUDqHJZqXyUDJ1HEAcrBuJhV/rCmW/WKS5BduX
yx2PTLCozueCPI1dpbmOUv0sh9VKjjSHBp46HDMuPq8eWqEiNQiI+mM1PZbt
PNEMhJ3J/GOip3nm/hM+IrDUwaf1Ci8zs384rkAgYtp43NEKF5t+vFk+V9xH
O7c5Be6u0tBH00xJhq5jptIQcxTAeZe8QvrAaiJtOfEwRyMTu3hUfnjOXzhN
0gyG5TJMu+Oz7n9u8vWnDIigUhobtbfsaHGvkmYxYa3RJVVRNz2GEeUlaUTQ
LyhfBTFPuZVPEwEjLspeq48TUZoP5lqAtTEE63JFXCa7vjR/fIF3Fnjtjwla
773LW0nQPy88JJUuPveTpUOhgHMWt+/UbiEG6jPHoT7YeKz/7WKiNCSVrxm2
I4BBgwy6M1SNZ97A+qu0xNFezP5e2BC61xM9/WNSI59HyERafM5o0BZpK2UT
7H7xI9eNfQFnCing+onirfF1V2Z3APitXL5asR8soTCYxsYD5DieEVhv8fwO
KlTs0Op9CkhI6SJk5/ZggjFVVnDSPeij53KJA2jaEIF/O8uvOKnS3Cgjzs2N
pBJQbBf3XB3VF6RA2qDoZzKgoFY6PlbRqapZI19pQry/DM/r7CV/gw/C7j5H
5QkkJtQjHhYyhu6QOmcMaQU7Gmt7zvjxXapxsLNCrXJUVLYCtyGZXDqwjKuT
mRiukkqS+j9tFMqe34GEgWE3ecNsEEosf5UNznGCY+LbJMXWytr1oEUopP8C
wUhaYO1QfrBL2XATQU2kHUragLbzaB3v0EBLmtykP6Or6tPff+V56MJizkml
8/ALojJiL83gHxTTluCgEhtyrBlbuRO86pZ20IfsaMH7KiV12IB2g97r76rl
cUxEeMubrX19zZUMvvhwB7YKrS2cjpTg9GOsL3ndsdQNbmBaIzLjedVGfHtO
xhhE5dDCDe+QSxYntuPgBgGSIMiQ5uY1B1INv+v/ucnX1fZKyPnRkwHVMUrV
2M0xGGH88EAgKCrilM7mue4PzCSp3L0Ps2noxTPt28RAg3SEkXPxq4SyHoT2
Q4Eoj4CTET8OVgKPdBmscIEClDVE/LH/is3wFyYdDbCsb6Ffiucd5yjIq/bV
7baIsZnN9SSbSFnuf9RIBbiwpNy3wTt1Vbq180PzhGB14eziahJKnGyzv2c/
Bvhbs+6KFMCNGOdOAkOsduTSj+URQHD8hGw+knTKVHvA05jJLHOtOUWobK+e
s9PZ7xbIdNUGDVRYx9O84o4BLlGJZNI/MNWGjQiaiPV5pc9rVanQZfmE2ltF
/R4IhcVAq66dAlmHd8MKTQyC2/PJwpgxp0N5EIu3XULGGpqnHfxq/IKcJnUu
m1P/zOvIpy2di18vxkuWJ0ohLJkc0shm0EyU+sdTSP8PPH8b75hlAARGTvx0
O7B3Sfs8y5a8INRlElnHSvJc0SAuNWn3GjI56fBOWM/riqSugzEKqdpSTMwX
b7m8w8Y+YycWEyGzljSAavdfQc8+qhmY7o7SQwrsJiUlkjqitFrpmI8CfINu
sp3ePkQ7VL8POlbNgLTGE5aSX6UIgawaB08J7vEQLebDVccRdtAAfJew6EIJ
vG69I8vYmsNhbqKYqJPFDquolTlhuoHMkJT+7oZuEKbDL+d/msNcD/p2opAQ
kXeZVdC5xyj6k4Nnd8HzoY7xNmDB87ZPRY9uI3zGobMrE03ssZthxlX2UflH
iFvpiaxBRJlqpjF6pYaF4EYevhR4OpbfI5S2o6h6GTG+nunzkIM3mi+YGQFF
WpZb2xM+I9Pde6KRn9DeB41nUD8sOhoVt34dwSsmZXEQ/PLE6HuHItx+HPIt
OqUxzMMzWSZVOkS/o/PhIPmmEGjZ88f7V4RHDffcS/01OpONqUN+Pl9z2z4c
o82ek7c3ek+ShNMFKFkcGYV5KqAi5wGxCaSiVUmRWT8Wm0feQmbEzW17fa4Y
JVhIcudlrvscI1FRHo5zNmXQgTuhEeuJv9QWguidOZrwX+AwuFtPEAw9zvF1
q5g1yi+EtKul51UJqJOZ3wgYad4tFSEICLD2Yp1H8c/sms3xAnyVI5bbxQ+b
XtHOgRTvq00ERU9rwG3yAK0O3cHDz0TSLPnFhT3IjVCoGP/okkTaoTPiQpQJ
E4w64TZ4Ma2SRDT2XDmPQLV8cZb7fYonQ7AzOZR7DEbr2RtkIE1yQbLTjWUp
8/6tnSfKISmpwii2oQbVvUmSmsUZR6o8iIT8Kbef5PdW7oCR9Gni87vKcZzN
389/zmu8r19dxJjF4ueOxIyjXgSdchCwGFAD+3W6KVWd6E2tAISq9GSd0PEu
1PVSccxfbvY2BqIFbNlW3kPpKV2KP3nnFu/dSLpvZPQiSPHQOcdOCwE9Oz9L
cIPdjDS7BZ/vcOWD/tvo93AS8Yp8zUrj1EgwNWiE3Oc3ljeHM+5mAgiSQSKG
6zy9rH8vrEb2MberzzUirClIARznSj6fXNVvCms+ZQRaH6nbUuEPcIjEG3cL
T57leLf0kiM8PnItlVvA3hKlRFxWB5aRa5wbO+GRNXiJCEV3XGwbCkkErnLc
vIdoTo1oP4K1fejJbf6zU2NHjni8Cb4envRZeUgxZFPSP1k+FHXGRUX4qszr
su3t8FSxc+ieQdwC4U5tULQKCDzqgN643uy+pzt6UNR/gGDMZfXm+j23zqLY
6FzB0Jc42c+Z7NEGK12vC0k6yBZPH/m3vL+G1+vUk82oo39iEBcIUMSdqPjF
Tlb+pJt91P021Rh+3u9aI6tWdMVOKJXaJl3w6obkgrQvbT2cgMkqSHgBhLOm
IsK77l0x6va6KqlKh9rePWAF/vNa76yQQ+PCoHjxmxqDvmurqjfcL3WUaDiJ
dwsdd9RqwOebn7gk6QF9S9FZLL6pAgBZscr65KNCZO72YJeQo0/1Gc6pplqt
cPuNHAAPCaBNddi3dNsqLiFYFS60osn62aTeahn5PgabQiKSlafyumrv1OI/
NxME8R5ULANsvYsZ1z7GpwZHnrB6ogVKJL3wOxrMCYA81WzcWjcYAzZmIVyL
ScEHdUeIipn8OH2Fw4IZbYfOgmews2Owo0OqzqoSa4ql1+cSiAF/IZI2wPvK
GbBrfNokBqRB5JDlfnK8flNRb/SoTykqI8XlsHFA7meMy65fdZabbzRFUdNf
mMit9XpVSBql4ngyMG+9Vrh13dfbof0UlCjYnwmstLC6F9FMDLIpsGWf4Whj
MNGOmlfA/20UJFbutgmIvoK59OrP/kTBYfuih4HQ4vga4PzwsWPF7kmMSEn6
RWjLAN2ZP8FRa+eiP2czWP+rHwnqPl0jMO6t0BuN8nYK3xY9AKjyU9yZUGFW
rZ/Y6X3OhjdSxjHkHgX42nHzXIKWqMgq/0QBy3aoKond72O8fTc+NATIxWzW
SSgipb6YgfletCQqIdZDsBWjZuzK6nkMsHa0S3WkrMN9QnpWdKtI/CugO3o7
PmHKtoKushP5nfGCvdY/Zlnk3I2hnKyes3DWErlHL/OVPQ5atI6Jjps6Cnjy
VggtT96ffmeHgyHQ1/ikvzCtU6tVZBTvhiDb6gEJo6MvsDkPS9JIJKTY764i
cWfRKRc+ySl5WECFaxKhsTkXgmigVIVatbHkVUOwTkHpohZxHnt/0ajxn6kw
gTAQTbGNbaOvdf1oOJQI96NJzsXxdG7Lo7/mvO5QSw01zwZHtS96MOqYr20l
i08ACZ887giAKI2QzOy5DxcU+WN8vg7GP8+kbsiawfZb6WOh4ULRDEn7+dNj
XmOoGFOy6O9QvoACkifVINT+AJXCCRvKVzB0LVAAIXhuEoTNBB3G+ba/jlr0
LctuUd4kLpPx+LwECvkzqZ7d52hXkwX4zM0EQA0vtG8EpHYPE9hyQ3hElug9
zPQ30gs2UGLNF6BANSwAdfO4eJVS77xQvsI/QqqJ7lfG/P8YZ7L/HPivb7OR
rGpPsyA00q3+5k79VD97/fpYQCSguAtnWfbkkomswx2mdc/mpbclerO7+Xo0
gHmzqPl1ZPFE+tkZ+1FgQ4/4AvMN312mzKvEq1/qFFcls8lryxUnYyOOxDzY
usYkmz779qY1XpYIWaxG0NF79dyOGNJu6+5IQvTBqNo8KxjmulqObdfCyn3V
xaonOIxBRduLxPVvs5AiFl/8bMg2IYlAXfH8dZIvsMyOZF2dMfqIR2bA58hV
YPcfnM8xJAqDC6yyJFnU/by4voRU0KD/Ccvs3YkNy8E/XuvCbJfftKQpXqSa
ChU1xjPEa5o18QGuPmnKmDQRaIrbXG/PVBV3YjB5r60yYXjz3oheuvqT8R1V
WCycdUN16ZVMR6DBCckh1s1m36IJiCtUlGC8soOtvHTom68JqlkJP2Ze2+Se
8kApipvFtuGcgPoXqfaOVGIV/T9fXjMwLgjWZQBffXoE6tZ88zCeMau4Zlmv
1MeRX6meHtL3VJWj+y2Ds9AmJAoqORzmBsns4wAawjLJ5Wp9oC9/Q0jCGlFG
0m/hkAwFQ53YjkdBpgEaAQX1zbYMx/R+7HXJKMVJjlm8peuqT5NmnBRjXtek
xByPmvH0YAs9I31AycZkan42vMvphveCeADR2hw6NDGBuUWoDsISSgZw4iET
aEYRXmV9f2czj/efO4/aLrXMPWzxkctlv4c+UIqHe18r0Lv7mTQJVLWPB0ki
p5TIXx519qAdYNOmx0cEO3Txgh2V5kQiBYKwQhunIfpZKeQ3tUjrUZkxeykH
E+OKqGn08Ox4pbWMmbdzi8NRcN/djezM8vK61jNVeN7+ajXybR9PAMBjkuxO
Qf3yPKWbe4HgZeiNJH6fUC9+nzPRapf8kDX3de+SApY3vRiqOm7kg1oraj3v
Nm8QKH436jAoAZ1QRY7GuomDs5nTT7+u6XI4fPgpp+Z+Mv/CkY0P+UQ4MSl7
CLmsjZgAzCyKpBzKWtligEMIB6WpWBHjOX40dG5URDO5BSmPCqBriZPloSoR
70ZiOZXy8cpUZtS/dI/UW+9qcuigFV9yxgSAGkgecJxVpKEopu1+AcT6DWKx
LJxmiSPBU7zwiyuy2YDVuSIc4jbt94vLbhLwwBMM1ALLxuJ1csPSXYbmeK1p
Gp2c2PuGkx1ARIsFP4aakYa4AQUlFiYCQSUHJgcLICy1UBMMKknM2DBI2m47
+ZJ5Qcem1V5pl4s/2mY74kYUu8MdKaFz+HKGKoY9UrtVjbeCSkDDTl035VpS
VI2jNzeQZlInGG4mne3Z+Dp1pY6qXB7U2w3jhM/YiNNldas7SkhP9ukzFjjw
VkD2Geq3PBKGVQryCcJhVEfS1WF1lZdSTJS+nIw2CiwopVr74FEnAbj8bsvH
sfhxz89ZGqc1MCCPQomEF52tWrKJGelE7PK1ei7NAAsTZNS8qxM9Ikwze4Dl
mfdu53KdHP0IS7VE20sx0ZoufFvH+F92l4U+0XXdIRBN48LZMLsrh6csfO4m
kAhyCfCRUuUDkc5z4M/8e+ddKkeAiE3JGPGAj1TudtnXC6UUff5X3QO7XdDV
i7zxFssZeBvoj6iI5jto/E+16KqgF7MnWdUhhBR1GbEP+klCDVh2LAjf7R+J
cEWTJpqBSawEKRfOuVWHdPATqLqcTTH3iDsxZoIzcWvJ3rB1jlir7pXfks8w
rs3MUi7x8NcXviSBM5LkbZ3aKS8OKibRnXvOkfBrwqRnDmCkzQcBhhzFMWuy
/V6Vz5W5mFZMq69ELtjAwB2bXflkDAZkpOsAEfr8dkV59qcDBpheRUU+AaWz
eSZQp9m8t8mya4BiDAeke1R/mosn4I1SU+p5hLD/lcSskUBDw4kNhNYh7KXe
OtGaeDLj6Y7I1YPGtkgXVMoAdWy0KpdzdFW7X6M6xEHXHa5jstpXA9oN2KWL
L+KCRfcdaVwNR+dnhf0a21CPoQLlb4vBaQsb9h4HQhZfYoU5KQnROzPzcvuJ
Pm79ykGDR+nvqdnFQ/BOrpq1jwp4/3bBkfeWPso8ZfxaDVzBLpB8hy4mfjTE
TSpSpadeQ5seHnw1AMZmsdZby/ZRTBq+CFpHw5yEMKYB79o9gIHU9KMeJspe
zZK9PHGBuWzSZv4HiSBC++pU//239gT+DS4yelS4N3NMlDYA79eLeFx4Miyy
/Qx/X1yhZDqWD9URl6XtxaMhPpE28X+O4XS7lhO21aWD9qXeDHXdCq2gz3vA
Xa3R5xI2fHm7HZGlu/bgyMcznH5vIAVUKnpccuiiNu+bbz26hDcNq63/TK0g
2zDNWmp8tKVnCa4Lk8Oj78FEO/mNA7Sg4Ftffah+umI7SHRPb8sQtC/enf/X
oBxQLy0TbpRji1ZDhXqPSCCwLMDTg5hEwfXSYxuXOOgwyyf8RdScfZgoIGLL
+c+dyg6IZ5Wfz5hHyzMJ85POnGifB78180d987FtSOWyRr4oDAG3QlXVQQ/I
hIi6I6fSNk6VsE731xSr1iJPd1FirnNALqeSiaMTddPtL+6tlqvGvH6Kp88+
T6Wsumpclmp/p8Eq437J4hucieG0xyjTD14ej1Ex9OQLnlHu/t6FswlYsf9K
4AwIlX1D8nstWxss29f5RkIF6symXDDUolBMMnAcogACRyxUzMSkaMBjGG7W
B/PLGlvqulQlJMfyqJrKyBFrG/dHRRcqqdKy67f3ppPn8vT1ZRTGGhfKZCFl
DyZ4RisL775aawqcJIOnLC9eyyLpp2tlIQJtKcbhIko2nQYeeExMBRmEUbMn
zFDdwPnbmFRzI7pOOFeKBowR3O6Z28e5Ut79DmeuswBrUUV4nYX2w18KUeh/
iV9jmGcxD+D5WkStaUE9UtEJ647zjn+ICTCS4oJraquzX2Dy2tkavfdr9qO5
5WAGbNSG0Lz7nOb/Hqs7BbirYwzChCRCCmu4KHb9/hJBskEyKSz8NcA7SLIW
qNa2fpvqeNnompWOig04sySSb4X1wvBc1aPZIgIGL6a6HxtE72VP6368FE2Z
AGwGq+BsyRz6lj02QxueYRlq+mu6dSkGY0VB4TxfA4pJQYipECA4AtA4XnfO
svkWbkpxYdXFgrga0XcfSfPHhUP6PUhtB6vBgPp01ZN5Yqf8PTGed13XDPC/
tXbwkdY1WkFL9S8W3/KiEmZItNx1ZazVSHT7kGZ3XXgpaPKmuKd5eaxvWeBs
PHi0fJDzLgSVgzuSeUUrZ7URAjE06SBOJgIY2RFcOitalshVV3kjmjwQxYYL
E0sbXuEmybSlotkDO654dnfpkuP603pmUypRVeaRZc7501IoO9PC1tpLIVRT
vvFEKrMm15oixABWwAPMyT2upjDrZPebVaCcOI3zsyGlQnABOUBbSDZAqujk
In2oT4b4vENYJfXiPjvAxxwVzCprCY7AGNC5rjIDT+r0J+XLiEtWF2DfbGcK
cdbg5zhnCGGOq5VRayg0Ud8zwNhrxfYZ51cDoGs+ZM4RbXZUARK3kHdObtCZ
nXNPwPBqMdhtq3pEQgy7qUj9qnL9LmHAGRke7Oo0RExBmZLBfyhsY1QBfG8/
Z5CVC3mqc57Q7tcMHRmDepI6W9uaE8uIf4pHgUQ0ks80P6BhKbo+5JsDQS6T
qXn6eDCSGQl4+u7QttE8TQ1AlWNgcytyaVAFriaiHV6Yg4Bt7KxWsv4iG8fa
HOWlhfKMIwV3LU3BMLGH0py/dMzymFiT/ONvxqjEGWgFwl0j19KICRrhgXWg
OIonbn8WoK+SCUprweLsBJlESimrX4w0AdT8c9rfEdZeDkiLt1nlqewwbo7n
72yLCX5LTE/HIZufLqm5lG3tH+NkcWtb1NhriWjRApsrPj5eXJZdWDYsdBOQ
8R+2MSx8xkPPcuCVyNqTowe1WSVAmZWuYgGl2US/jBg+FbjAWGM8LiRI8Vsy
VHVp6tZPDD1BuwJA0CADyiPTqbn6AdhLtkggxzMVEmN7IUOGHlD1oZ3vlG9b
tfkBeber+YXtrWQRlOMNPmzarTDC2D5zZosGDzO9fXBOGbvbbqfYKiZpbqLO
nZZuOXpCn9JhnAM+FpoGglS93ZuJ7M6KmqfVF0khoUv7jH7hFfY4XvFRte7u
XSLch/Z9P/qmMlrUzNTeGjFk62GqQLRpiLeu+50grgUVODFKFo4h7x5NfRP+
0tYIrrKDZ2YQM5SBxEiFhjocudTUbxAjUwRS7RsxHgyjZnr1QZp+nIeexdf1
5ti6eKGj7pnXJijK3rzh3LpI/cVsrJz7g5uStpEl6mjxFZH0wnP6F+uZDJup
Yfzm2d1MVG9GS+HK4aUSJqikuYkRhs5cSddf2ekN2qbuBImRNFWdgD9gNmJI
5qnvVMa4n+54Dn+dW0Q1NkYS1kEXJzTIFEWrzBA9QC8RKKxEXMw8/J1SGBxr
8wlQ3sAAmlsqf6r51/L3xJXsn8J5pXVasXzNzAAoUY05MNsLUNttOfr3c5CW
C7Xb/PJ7/8hVbwWoYwBIAu6t7+Z8Ot/lobAH+x/CmxKmxixyLHozuVYieXpZ
t9ITpgMSDZdNTqo5R+tXYqwQ2Gjrw3MkM180/UjTUAH9anqkE0JoPp55qW4h
ZtcWmgz5sYp6XukXFREU1hZ8SBaETgYfZ6P0jGtQj+H4tefE5LQ2oJ4x5Vah
P0GMX7CVQgswDwP3pOCm8ItRUhj4PmlbJzjCVBLbWeH6W6xAy+caS4lwPOWJ
4Bl3EXwBk3v7okft1GwqlrPXGWC5kfPAFLHfAnvOQkGZxQT3SxyETHeCORHZ
aHe1jZn9A4D7jpI1DcsugtxLAWksAA759QUSsbCzuzfiqKI0lbuTq4SFF8YL
ptwCypY2IW6aVYpqZvRbCY1xQi1Lp6l+B5LZLZOZzD2tCBg8eLTS25USNLEe
0bc8tJVwsnFK1JqEjIjwp9ohF5lz1kAQkZGCT5/pfchx0+gKTykcWmw1ooIM
GwCIpaSHGajsx/Q0ztzbs/mTrNP7xvqtaBdjbtcZLgZnpL25XQNSWFF2Nad2
27dvHJsN6ZDubjCSuUOm8gwYLPsLXg5uj5dEU322K68xDjdOd4vqj16NZewm
NptEWOoEijEVtG6geB0DGf8aP7bQ4nbRQI1ocUH0wsxMF6tsvZFQyy0SAuu7
pqtg/2CwHyzZYcJ3h2TvQRsLpTMGLEOelWQyHSXp5qcfzwb/2MfgPWzpjRsY
1yACHHkesYLFhWt+DXq/iaaUG1K2XvYWcSZ0z3OEWPWCCr3kFlnHTKqindM7
xSyaogKhdNL+o1o/yjGUuPYFVYHmjjH8giE6XkV0VHkQF1zlxoCcqNQ6DCAG
w0s+OXM+kC6mikzK2NQxvwjPT0ei7JohHW0epHmO2lEtaAgMvWLhH9R1eZ24
H1QayIPEYGwxyyOrhgdw/hopJHuBDo8dZI0HlLvJDsH4PabGi/V7WL1IF2ca
ydpl+iHLlzmyjzjG4Vxn5ny2Lc84QKlAKAaZ8wD8A5vYVFn1rudKbTcYw/Rq
5X6J6EYqCwZXdTABDPRvYbQ6MDMiiPsUQaHNptBg70RwMyKjcS1cU0VzWInM
pMII9Xbc6eubniBSH/SesgO/LW6EAoIAZS+WTY3LhmkuAAOVWJHVRnRbK73r
WDEjAakYUwmfxe8ccEPMoVMU/t+eHn/BFjswjgr2lgmktqaiFBrWLM3tXuiq
6V7xps0GC47qXiG3zFkqxUfSVDFjt278C5bUkFoFXrjgLPOu7B5SOFCQPNTE
rKjCUfSKBl/XI/EAErTb0oiU3ysuyWTtRjhQ6+ONzUwT2Mh7FRI0kAXTjcs6
O5BrGvPHjmichmICHmB+E/OdlB0KoUuNx+yxLCwYzhyj1fN6oToRP/4NPyrl
MAxI0Q9ro5BR7QqSHtzhCYAJfIU9RnR04xbYnT97xc6BuGQFGMQfxVCrINru
Ct7SFIvFg6MqZvbR3Brhh6NTrnvRdsUuql4ruXcm6mHrongXzQrJ672YuKSz
jXFcAJbHGPWw2RPEm3MT1fTRqBtFFDxNsWKDVOLFOp1L1pt5aodzXgjYkZLX
hpqgSuR4cYsolDwikM2rV4HFHhe6zvW6eKJKrA0SnhRzC9Djws+CL/nIhqKp
zP5+lPgeGPhkBlNiQnY2AMD8WZPms/XigBFA6YcBNYVqnIIbnFQnbf3z9Ybq
zoj4Go+3a0TTBSiWLzymE5sbPoqNt+2vVrdAsyai0FgSFZ1yKqZf8Kysx9EA
5AChcOvdFl0Jalo2VQc70NRlgv3HSn2TanbtrRuuaQnJax3yaRUA9jLvxPCv
zTsGzZF6D0mZk4fmrUlHAzR4qIEcJe2pzJiBo3xkelaa8NTUVyQMKwxQu69J
iH14C9IIw1rVkCg01sYjdZDUORaNYnIYMKlA+WopMoALw541lnPshQqQQ8TH
TYk0Ot73aad/hlOOUaqoMjdz0Lr2FG0Dck+yJZrpFwVMlhh5gaq4dJyCAgDs
d/8yFkoTUzCJ7dNHrGBTkggkxm0blIxhFSprnHkyBk5tN9KWpccvFdANxSZd
Hb376fDSQ21ZuLlHqUXv6V34MJTjVNVRFCl0co8pfus/bVbsaOWW7YJfsEMG
SkjtJ27FEF1DcqYgj0L1ZLOveIkshsaNIQYEZZB755CrGq8fnJ8bU75fXpO/
GogVehnuu2VdXfVb06WIjA3eoZj+fs+1C0H5isirGGEuc5kzED2AuAiroXZV
aIBFPvX7tgVAGEviWuSziNYbckoajEREPl355oVe0n5EL+rf3ysdzcbH1Miy
MvJb9jMepkjALI/0KaBcymv+J+o+SvmLh7567JQ0a87eWaTicBuUIu384OQ9
5ddW3PDjIzkKtcx1x2SqCzCIzmQIsHAuvpp172+Rr5E45wneJgmzxdSgHEo9
rWp89aShXf8Dpykp5T8EcHBlDpFf+ApQRPqq9TIbtpJJpFf7TSkM8QmWkPqO
gG2fs42f1VDI2XDd1x8NH1I0uzc7Q6mdd1kUgQXItrCQSjL5V6M8kU3wg30Q
SkiNMlTIl3lg+7t6k3zWFSu2SaVD776ZUspEH1Y/Vb5elTvIn4VXyjtbxIIN
QpaRz6CphrNLD4fkAQ9HViAHh9p473K0MpPo+bxs1oqnujBJ1rAhPqvTLsRn
+Ifg08Wrr7HJqNWwF1F28BiTDNPOzlgMnVJqJhPe/uFb5xWlwpbaZAWD9878
HZ6IromQO54hdXkr+ccS7ixp6SjGk28JI7qJqt2DDsEX0K8JBdlUg7D0FqY8
5dj6Q4Vtop5AcZxBO+7MRw36ndptWgdR+OZtkvr/cBE9H7kO3VBgty6a0NT/
9JVNX8v9hAG23rCpLkQI7uJkj0CwddsBpx5UqWrAE28KKutHn7QUcN9WfPDq
Ds0i+ckvQBrLZTfuMY+OdbE1MLqoj7WD1QdBhf3O+KW4lQd6G4SflsoGfTux
aH1dskt+R8bdc67c1hxKhso9G8Q64GQE0r2O+grVil1iyq6zOl/nZA248UEx
IUmKf1tSpyI8cp3+afuu/WyZZMQbiliTMlVMyx8fLROlgRIqEyDX7imwtM3X
odea1Q6JfTKJMlvUGRdX+GV9p/1WiMOaar+nKN1waoHJ3hwP15u3pVukSJNq
ceK1lNGDdnseQZInrHUjosl3cBTopmmz8NIGp295VLgQ7wd2pDWUVyz/Koth
UdtJNV8mCb4epUR2XqcQi8BdmrjbSuzAsMg8FFtG7oj3pDYm8n8j6o6GXMlf
q6dkBHDBhnRWq0mehtLscjMgMcqoDOXucEAp7UnU9N1iL0Y4bI8350QQg0xf
wTDozYfCsrmgSu9cp2HUPt7vYNa90FRBYdQaLkQcpwTwCT4BYzh7cygxk4iv
+bG86cgWDI6jMVqHV2AJNwnfOxODHet5yH2RpeOcDaub7lC4u8L6bqPzx7Jj
aBQBR+Hj9ErlZ/CLrgeWAr5hEbx2t8NECW411wmVnFzLqOpzCJpmSXFVdTAP
GaVpSR23OkZpWtIiKmgCi3JHEy/cTkrHrF2yFwSpVF7nI5IIxaSQQUrCGewY
ESRSWGTvn74XnrwuFNE0Q76KY5IR2PpjfjfLTJR3SWUeoyr5ZLVb6SsjfxjC
gmrbbkiH68kHAobFFvAZZ/uBGDBJO0YTxFwoQKWMTs5fk5gFOhk3wTVxcX3l
BWP7Lrfgd6u81/gVgNl8y1qD8z2RLuIq1P0cGlNc6ztaQMCCmcg8sqmVj3BC
OvEqwb8QACXzKifqS2rV2xBCLoUP4K4ibpWBRvBadcV7+olBx1tTNHpV9E5f
8wqOByJpK5HmIrKfSM8Eb/kkNjiVP8g2TWLIXTexXtDqDq/aMSdlthopH5N8
EQApY+MJWfUi54CL73BMuwhuo4fB0FvHQlIorARzf0I7Eg3QyAC05/V2i7aW
Yv9GljwhG0jBk/F27s3Ice4E6QC6TtKcAi0hvLUxX8oiNWJraoe8mjwdRkct
Pm69v9z941xn9lxXq9tCutI3OcLmZamRtNnqVYP1Sx4kcHc7LmO6hFKEuRZX
zG8RbJbEk9IwHeIv/L/sqDfRadmiQ94V8/K20LIEtDVbhtcn5hvxRuZvMcxF
ers0h6S/beDLbIEzKd+FHN4w8RxWZfHp6BUzrMs2Tg4mP9iKtTJBKwiz3Dso
qD9gajj3RPEnNzyzu1AEmrMSFvCKJhGGYJ2VoN3iscpYZpjHGn0rtEdHpLpp
joxh5opHPGKdeUqq6YX1jQJ2xsNoj8Cyn5H8kwpXoSa1HTb+GOx6W4SsQ1n/
lVEFzOgRMRFVIwKyv0/lxKbp25vIwFKqfxdBY/GNva8TEUgdjPwyTRhjOdvD
1GdYaCFvgKW7EsEmp5/kLaR36l8QODYXOoW3W/dDdg2aNhkOnXfLTSwEpTHn
x9NGGN6SNxkzrXyqL32FQ82jOhSkg2FAH/Wto7paEpSfvZJSI0rRnhrJxOdW
rgNIH7A2T+bzy+y582va1DpXcS2Prr7BsGo9xMRnWC0+5dB2vi6jTIDBz97u
wSAfv5ohsG4u4AqTwYL44DUGlVMOR60Cq2aNxogaTRaRgu2tQyyrAXcm+ZtZ
lrv5ZXXE6jUxlqdF+cG5MVBCrgXgxiv9FRfzVRRcLInw1A822fQc8EgRF3sZ
JmiXoM4xYBlg/AK3ktbc4NziwnHGB/7FaPXYLbhpdakksBlAC4WgHcebN28U
ovF7iHGjgc4yT6uhCPwss4i2Z5I7/TlCT8D2W8htXoAWeuRFiRK86/hRqlaL
R6vIgHRevLSX5hBXzJ0sKuWWdvx2BMxTuZnr5oRapJkdTPdUfC5YOaWRhp7s
6YtpyA/+MFLqbKLdNB7ts1b5iDQrINykiFIyR17iHe0Y9R8B6DCLhqg4qxH4
rBX9bnbhPEmZLrOc1gkMdyomsRq1Z9jmbzqbmAY2DAEq7Kns/tisbKcVsFsf
JtSXbQUuSFO7tGbcvFHLZK817sXtyK91Mlh6gwL2s44DdVrwcxBFGWmyrPp7
piUyqIVrPOvxlNkvQJe8RWdh0+E8hdEIHISs1NCVS7n46FlfgCzFMg2RGQKf
JCjndIunTcVlaGrbafIjuK9vkhmgvsYwSYLBLa3EFeTdENN0rwrtMxRRt04U
8zWpmtBeena3HAg7RF7zUoMvDoD2OXlXLLkOVStOGIqAIy8+pgAHOsIg8iar
tu5A/+flBfIWZ/DPqlBhcoASsTj8hb7IiR7sPwqq3id3RwwvKAfB/mapoAx+
36qupecU5i6MM9vzK/TCMJ6le9y/X1MSZcVc+MebQDRDf7beQmenn0fkWl/5
XA6YSuCBZXkckiXGQTUN+pfwFDbsCWslFWEMwL356gtEysYWbfL5B9ivZXGy
7qOvDuO4iAOEdsbp/dGxPNGL4mzeiqNMdb5+GmpIX3dKYiBxdLwsNU6EOUWY
tsGORXMtZdmCPsGaljaUemRsff3l7zHADzhNS/lgzWQnCqR7iYtPfn0uVxW0
pcPggluO0xG39BXnS/m4ht3JtQTUg5zSL4HI/p9vnYBNmGXVvH+n4NexrZmp
TiWm3gmfx6WBNpRTiTilM67O/0jb7TuG4WCilfvb2wQ/pMdGslntDeD4ayrG
dYNuixeJr3Cf1wOECxXrkY/e01638N0s/GCaHgE0WXLW2Kcu8IlsiYSivrsu
orrUCx9Jylibll9dkAFNfgA8KrP3dqdZUs9DfhaTv3lcTTvPABWhC+AeNhS0
6lsCY6lGRRyFpCIIbK9lOfiMqEzrWtpfYB28q1TVqQqErXgZeUEKAcGhG2C0
lwOy6CmfakWcZC5YHXi81sFSyh10jvdw3Jf0b5tpFxbnhjdoQsibuEFSb/PQ
GqMOWGUrF1R9nFS3AnsFze2hQhx2uz4zIchnVwWLi1O3OtbgRPbb4vnNEx5K
r7FI8CoKT/Z8IQU5/9RAu1wVT4IAHlhy7Dpyc110RQBZm9yTaKIZObzl3Vmj
9v4zT3flu05BK/t8o1fnq4RK3eib/U1DZdhjbWPO0FYqF+eMiMEBqMKFbbI9
uaUbDsw9FOGQK+Xyw5xtg6ATvCjJkFlu9l1rkdBKcme+PoY1zQB4gr27ulIc
uktMg2g9EMEIGL118BMoKyZ/Q13w+DA3mUQ9srFHTIUfF0ACOWAoSWOqh4xH
tIIlQxd9oqlkg3D1C9vwdD4SdG+fNnsC8ajrET0hEHJog2dw+t4Rs3V2x/K1
4j2ARF74ESZ2Ems6HMIv4u0DJ2GwHZkuTeu3yDNAjMQ8xsGK+2IfUpEtXIgf
yxrBoed8MamqP/lXbDQlISyGFr+qyBfP13+ggFQBXgnrWK6eBJ3u+pMiBbxU
dsCOGFq1fh3Ukx9Yeg0WLEhwejTqt4n6Ll/nfvdrVaos2bobI7uOpK2zohID
qYYH1+mDa1rjI4YtOdlrG8c/9TE9wo/u6WfY/s/pnq3AFW5aMAHjKdPhjKHG
NSjo7r0f4SVvHJC1S2pXqnvGMuieZUYcwqIJdLpLYCWgYA/6/40jsnbM6eE2
mM+elMvQEWvyWM7vFxtccdIaG9ZhMju4TMXDLv8MEP0K+NZLowEWIlcXFX5s
EYmPCOjL4bXc2vpM/pDXxjW9p5UEiZjvhMvz+kH19YDXn+H3bni6AOIRHHfj
7AMsd8uHulhwPorqkCjarve4C7ilF4Pz5A4T0963zjE6jkf5WJ0tBoyzWbl5
QbhOlur6NoKPnfSRGrVlr7dbaQNEGHMPw8HyMyy/2sY992KF7TsoCkZp238P
kSmPAIS+VgrnTphHFMcVX+WRxQYrkWIJwzuQhFs+YxY1sz1F/Gr3czdIygEo
fM6iR6FsysYUgkqqkkAKcWqOTjfVqpjlR0BsiJaOih1MbR1tOM8aaYuYTUSp
gsWZ0OOz/visdnDvYljfebhhepo5FqAbDqQtG3EeEy+EzdTKVmEv+zfLbFyK
1CiNSZDF1euuziNu5N4e9TlldiW/YipViMwEgUU719nTt0ub4Sxm74VfH5kf
WLPV5W97JN2LoSrbPPklGdp7SkyeogKRvLIU57r/LL3S0egNgji3rl/+1WB8
8v90SM5hhhc9v2jTcU5rk+I3sc/ASIAApz5938CFx9q7zZb6b6xyFrO+gIeA
hztRmOB5NuDnRG/QVP7Zfttcpd0jCx4ShrbUzcpC7iacF9Zf6XSqT9EeBYDi
1G+Hs6q5O4mtd7m4gnMdP0dJuZIdprvw84OSwJmpyreWW90uOWuv8aHa3cnA
wxZFBIstc1Z6j0EXXN5riLlM1wtQrfou6s3PMQXqDu7s9u5qFQG02+4omHdl
m1RIpez5THXV0hnA9fLQjeM6RPagGwcT1yTFudvbgJvDMMYlzPPxYFjPB2PR
UUX6APQdR5PGbgM2Kuyy9y5qe5+5g0ym9uV4UN0YUbu2UW29/vvUAVGP/9qt
Ae8ezLEsUcaDjXAdFPKsfPN7NBZvsAKYmYsMc7YK5eSeqYH4RCfiqok+WqfI
j9uzcDqV6+SsVg9unhV3NuO6m/12NgaZkcJWIgQFsUMfVZWh+4MezGzNBcRd
z4a9sfgz2NLf+mF/4Y4/RWx1YuXHQ6ikQcuguLZkAnptSwbjjZ4iWJzLU4R4
EYXB0rbXf0ME+ANX/tx0xNEishFfP1pGmt2ASjBYfmzkGgNWiulRAf6ygrqB
zCRr0TcwrvxLYc3gof0qfxEL03xup+FTVZzDsoGNqtSjx8fYSui5wbcrbHpp
lwcPBxVolODWOHg4knve8ShuUJSogbPSzGWZlHX+4YuFIEm/wbSk6vjQqnml
39rmHc1z8SgUMJ4zZ/1N6j4sb+OVm/VB6CmMBgcRuf+ak1/IIqfV1ZSbkb5s
e5Wo1MKzSomyig2gbgfyv7S1urgkwk1uMvTZdPS0kwYldWFwC0pheL1XHPza
uEaQ++UNh2A4OAYYdgOHZgWvu2Tw79N+0XJjBgqqQ2XiKEcRoCN2oGPbr4n+
TOcau4WPTKuSOPZXKUcIeLmmvcrWjse5yTWzBKF2al3ZoVXadT8p0jyBzv8C
K3br5UDyNrSl4XxmGf/7hXkcUUMjpRTI03w9cQzupgY7cxMIRebd8M+Vivzi
9lDwXrPMS9V2vsqCsFPMDoq+ks7iBKhptSLC1QtwENY5S6ut8/p16h8a33qg
erCR9oH+Zis7D05Tqjtc6fbIw/6uw7OPmKnwSMH9vFaLJ3QLTrVJipeM+lx7
waVa2W/yRJMat8Dtw9JZJ5XZ0E6a/CR/FvQ/dShw8UNE8Di0O08Cu86TWVNT
Lw2FlUGiiBiglZojyOrxYmn36Dd09pLO0QNv5pEFLv85JfozPx50TEmDc6l8
FpVed2GJ+F5jym5TRIDCDkTlVWb1K2oVqZsw80Rq9QyDngJCjQg/w8Ir3KXK
Kd0fSxfOqO6oRM5EWcPZcGubjA9gMSPK6KMV4d8/6ARF/QUlDukTwNZSOPpo
aKaPb6q5kZwnRVL+0Zimas0rAmwLR03HZP7fah4RWPOKxhrjtV2j8+Zp9TW2
/SAxfSwaKcH79DzD4WRoIKHKTpHpF1qVE0Ea/Ojn92zhYw3/Z6G2rrJGOqPF
layu4Gsf0aDBMzVi9wjsZ8q1lfR/ZXafHXN/A/5BdaH/7BnY5ij30B0RcCd+
rPxJByFIAR4llYuo/qQv2QfYbCa2i3YRVVlf/XxXtmfQ+Wv09Qwwv0drSsz5
jKYnuLLUZlsDnzgKRIyh0gi9wPF2yxkVjXBf5LUUQmoUOL0QAHRemzruRvAu
9bEtsL5KtPINH2gy1zF+5D7QG7NYENc/iu7KLPlMgxftRielVYhEQ5HiFQGk
NxA94yvXA6QA24IFg/cTFbpWlyPMcbs/uXsNuBle0I83LpjIF2tSJNjexpHq
IQX3rGk2z1MFr8n1mMcTOARHJ1BofGUXuGNEmmZYLD2jFVth/BfZTIlgsIlx
O0mhLS1wjlM2/xe5KDKpMURb22OcnOU/5N0DAVsBIBfcMla1CVr40TdyjTeC
lV6QwP0xaX/3FpP+x7DGwsNBGPjZQ978/q7gcFehZXmBaMYS2QtS9P0c13+d
uUTaWohQ5aik3yuDhVLzgq5Q1w7vEsUZsE9CfP8p+IjWPHq6BOJ3Az4JgQzZ
iVzZaIaINbBZnXaOIJ3ZwYzFNKvRDanmMFj6DwBX5mjXRoZebBLdHcsk8WcW
CmeQmhKElkP3s9bbTEl7/WxcRDAgkHX0hOA7RU4PWci7x9+mFgZfn8w4fSDb
l7ey3l/2CI7w2yQAVQoFf0Tlytw486ydldFwV6Jp/IPxFcF7JVQfwD/+JbxM
y1CfmkU/zEyTdSMTTMCOiv5p3nXeamxMTqzfcKi1NhVHnv0WAWARn6Cb1vV6
EcskEY2OiFPuMI4heTW/NKTkH/gqZGt+WiWg5xjPTBo29bLNWJNXOTsQpvaW
ZQHtYKrdbyTUDbjaWlqvkFmKR9LBd0ZC71OK+rpZ7y5uoJzbskXbDrEO33ka
DaGnPc6c1PAaaKxAQynlHWeMX0t4hP/lZtN9x5Dl/+GJI0H8zTUWGwkyXY9b
lA5YUHpxf9dJF6iPfZqrBNC56Xb4LahMKKPMvlJD2G+JwE1YqpqLGTuIr5Nb
fYWkMFMFT0qahwDqisKRtFGh2rkLZCu1fP03hWJO4dhfIn+ey1YQEsDEDN0p
UwoKssCWkpTQx3/LGvUZV7ou5zqun4OllUWEX9i0A6zPKyb+JbGJwGsC6jIH
r6JCB1sZbDNU5iHYrOmId5ny1H4WpGHwZkhsceslmxEnFUt8Ct5GTvpHpWNw
Na9dZSt+R5XT0OEgi0XK/I2bswtsIZEBPHV5VwuZdJIcQsWyj39rrITp0RqR
XmwCQ7a+WlFdP5gwFJ7ceVUkM5cpeNv0qKn7HEF3YqFxxtHPeS2LNe4e+YGR
ceOmd1wBdekRyEhKVHh+aos/2A2+JBHD70zJxjh3IN+I8kiZLsNS4Ig/4UYi
hJcMcv7l/V+ogDmTAH+a0tNH1KUuLcacv8BBTOKD2pLjOGpqqki6XAzE6ams
864496H/pEM+fQrqWr7mxdkKKJeaQXgt783to1xVLbWfBGpayddhdVHA06Iv
vMJczDRj85Z1oK4WZpxaS2/iCyzvXRQ+cogfn3AoMlrRIFYsURyA0T9KcfLY
rQxvgzEToIaJssnMeXkiQNb6hb/guvCE3QDEhWTjE2VU3Rw5Fm47A8f2paRm
GqByuZuUJIWrVItcBAP2Wvsd++14SCgXdH8HqJSNEW8kWCmDzfE8eyYmQ0+K
eD9Bt30Q44FyDV4kTtT33+lq3j49XWroovUTsP/NzWTidAL8g/PF4GTvzv6a
mEX1t262xWU7u8gKFmJ8vaGRS11tGPa+lAaQxR9Xr2wgEgunuvfqrF4JM+Z7
9sSaKWSNSzHqvxx0YmCEVEwtJthHpARKXHvl8bIBGh4bKxrivKb+W3LOJHqM
hY3cbnducmfQYb5G/BAuPmjUWoKBuLbhlK55ctDoPQYOaY6Bm4uhErgm4TrP
Zp16KPFuaZwPIhnS9b6IkGzMAfKdcx3zhJZf8/K/3QF22Uy2cK8HIrusLMZ7
bRx9nS54IRPA/mp2qU+Wk6n4Kqe+QlK2z6XqqEUui46O3RaBd7KUm2F5aP4l
qtci3jdTzl8X/MUb2b+Q3ZkivbRnYIUv7EjJpBg61gtGbepVOlqYTRhhDKre
PeUMm6JQZ9LLEuSvCH5nGmusnAcg2j6Zg0vxKcsWL/H+n7MMUK7E/RW1bQgv
Voi0luJNxW7oRsS/0gCbfLyZAHUJ/6bdEDvouxJ7OV2sagIRfJNfEB8lKUgC
Zgeo2NDaaO0dgd5OYlL3cKGjwE2j+N/hHc2iVY7BK4ZrAAr3zZypoBRN6x4M
ejoM9Kq44o/ablMU4SCT66JTG7dFNlGJ6KXD0QQmulu8rzQJiw29HCEO1anv
dF+i+Npov3pVDq821AvNWi0pH/avLyBtsoYQ9DzmgPrX3mrxCwF7dDJcz1sF
CWbdoqaAtYeyLiLoI1+9XM2onWg53pGLRyP+zqBv99gMgrxLbqzhzrddKv7m
CKoFold6BCT9zdsXGOxoDkp6WwofC33mEnTrmm7bykLBPNk4KpyEL2Jm0ja5
JswTo0HfNPMRlMmmfWVFdK6BSfW7IBySMYOpUw5adElfeyvssCbhu8IfOnTf
2r6WMURqoixeDY9DQk7ov1nXzG/iFCTor980fFBcVzKB8La/XWuhgJVp0IB1
/7Vf79Pk7hiJ7zDQ9OJ2+deLE4fHrea66ZbC88ACoYpUQf46jO1nfrIEO9K0
uxVgyYpDGWSoicUxVGzq6ditFrObyOInZTfKHzOs+RFqxXgIWb+yvQO8G2GG
j56sT5HXpGkyulH/ubrIrq/usMSlNLshBe4RBbJILzUCeRlhMg1ywAUnjqkG
dTSdSyERCrbrS3cwKw8UEsIvAHrpJ5WRR10UFjxYgoK9Edxpe+MsU7ykMPW2
If2GDOG1kfXd33Z6sqgdDDwh8bL+rQ12C7TwOjptgwUsIIeCdiQfYDOsqx91
tOiF0aJuixxBHCG8jxJwoHXAAVDb1HfRkmcN3cFF3OaL12JCvF2yypHDequU
MDmInD1cwo1Zzp4eWfmFSz/qjfGduvftkec+Y3pEsqe8qY2T8SSqPazPPQXY
TGa4J/Tu8+rGDQH2o+LdpEdPUN4HmgsIacuHZwsZZPFkGe3th8JFA2F6bF1y
ErjjagAUBEyn3fWlWCrhBHvF9FyXRNWIaVQdv/gw+IFdx2dQ73sUP8KqymT2
+oXjhuNkVFMOAwlESegZCU3vP3S43LjodGbgHUl9hictwfENRZotwQQnvt/h
HJiZBv7uQQlpPYxKIOW305wYZ0/akEmfhuwDn6ScThX77umO/5igpTl3VFWi
e8hiRmy7ki8H34iC+cUjjmJjIQfJnxMNemTtNNOHzgxwNw/hVjsl0BMzr0Wj
V7VjvF1oQsnII6D4QVagnpzdt4q1kb52rX44+do8NIZS15WE+r/gWzq6BvOy
AwcNVrmd0byACaJGAIDpVQjFbc94KIe6jdg5o/C15iRMtHYaE9dPoC4PwZAr
ADXxz6ER4cuUXOFJ5Gmwg5GEuU518HAXL855nvBk/hbBLvNCU99a7QihQV94
D4yMYSRxYh8rsIu+5nAtrSEitifZDFwIaZCbB596nG1SozXn5Aw3xCMm+AgI
SKmr+ALMIvfGo43Mw8dFO18DK1ScLCFpUWUyt5NEI2pqleS6JbUQftXAXbw7
0TT+8QpL8a8TwyPOH/VS5liqCXDtf/B3+uUcwG9MAujvHNRhmNnQ/wYPHI86
UOhqVcdD5q723WWN4H9gMaEPIPN00BL1rOAugRw4guPNkBCiBZuzFe+QcFk+
LeqmZ1YicU9sKsM4LaCnJRLZfYERPMtBRU34NkucFN5LQlPRs9C1ZtBtpu8T
fJ5JR4uQ/umkqglkgrcq7bKVZBlmWkJ5ibjzjnW32Wtt6B+B8oZIaxrcftdT
wlkfFG3fT0b/WYsnfQBoSyXXITKQuRJEhlkdNMVbl/PaoAiFlY5L3krECud5
CLATjLTvZS2SVUcptF5/AtrZhqs7KYsvvsdsZAAZh/MhYtlp4a5hPAsK5TLh
g1Zvv6qXDMnMzV9yt3K7t7OIwbg9As0ZRdfEhVU/+lgMhE5icUjm6Uwyzing
7GfXS0zrTfwP7EB2ED9pqKMxgqb8Rjh5GXK1XnkWn+3ljfh+t7OYsvFbgWhv
x1+kYxT659RhRcTmmPb+uo+Se69ivxOieZxH/XkA46fB5f8R5UTj0QmB0M1O
S8nEn7V9IEgYQiSP3CZxvervKvRFLDcTfpXJZrjCpzJoBV47Fd+uzKoLuj4t
etreG0BamDvXZQabNO1Z2gIq/OW2RfiePF7priz4dPKQq+iZGqqcLOjCfKmt
Pp75GAD++2aFrwTB4YkKuhrs+1kLBYi8Bq23aSruiP1G5Jyw9ZXY3GbemgiO
f9pd5epGjeuR1GhwsKYUtTdlD9s7QJztxEX3CILKkp8LlGO+IGrYwc7y8RX/
aF8BYcZ2K7f2A+CP6WLGi1HnKpdJCj/ErR3q+FRqYirJqpMHfQKb4NXqCGrP
UuvT/o3CU/K25Lh+YlnluOmD1+QX+C83/ybDR0xua2vuiWPkyAgqz5AhOzj/
ZWVsYpHlr0UEsfb4OSDfzTejEYq27Rn51BA0NzPWDNpaao64ZYvuWYSwCGLq
F06UJfPJDFTi2RDLxAGGIYGvkZyBKJYCaMQjPIBLgPAUdGzsDIsnpJH2pU7y
vQH6EXl7UZojRMovRHhozVNkQaCCx4DZ5fkaKHRq344SJsT8+Ef3d5coUAUW
+RWqYfJ0RcfPxHf+ZhNW/P6O5+rK3RPrpoFsnDghODpVd7nk0SwzG7nc80BN
/QD2v7WXX1RsqVVnyW91bEfRddGAVPW33hZefnJo8xpwnQYsuvlBnxQ0Pqu4
+zmCYjUzejz+VKyV9A5y+ycp9iAYUGq6aN0f0wgt+vqysMkoVDaEgBsaslyS
ynSQuN42CGVo48U5eu+QGVBdlt/Wmdp3V8/ck62gibp+6FkDdYbjB8xe9o6R
x1/TTLLKDfi8YcM7QnLETnYNgJWVzVbaY/erL7pKL2JxWCLU6gkl6g3opGFS
hWnCsGX5yW/iCm9wA7ynEbqVATGVebKFDlF1gZEPt5lvydZwOn53aBvVWnJ6
nHRkiM05Qvu1IJJi+hN1Dia9XO0qsMm4OknLfwsq3yRrMkEg5ErYV37w+Za1
oHzdgLh6A8VWyqVl54McZXBmV3uF9SJGPe3+D0Snm0CvPDDeB/gvdbcW2L6T
8dk/yaKwLHzqtTDX+YRyAvQn7WLt7BvQkWQKvxxf31e385YP/hwFPoCAQMqy
qMDlnttcywr00fp4/K26LW/znZZRTCf4HlWpaKD8Qk1FsUfVn+WMjPO9j/FT
VUj3kJHT5y017KlWPtumh6FYeO1rbJYRXvNVrWzd45PPIGg8X1+SXQZGb+Og
a7riGfWoMxZaRgQUq0/7ckBGB8z8RFLw9h1xLcgfQTyCtjTPk92rcoJZCmUd
19WKG+j97rssAhZCAtvWa7XQZvMMT//WP9fJfhCp2FHSQv4WFMJqKugDHyBp
YpSuKSFb9+++f4EMv7KcZCM2BVpcVkMH+tbk16TI5YpWaKtZyMzPhC+Z1vZd
sH4SRHIjsxX2iQAQYoESA7QYBGREDh8ZcnxIgyHm6cMvdLIxE4kwwjM+7mJI
KbtAUJLozyjdU31VBAykupn/vmLQqbDmnB2cURLotCPPv2BYkLiWD6114NlB
+oPNJ93gvcrq8hs9z3uSB0Cs2w7J165URxNWCCYK/fF+qunf7oNJO+qdKJ/V
juMh1taw8i9pJO63wHHcHXvy0h1Ouf+/+hHUj1wCbX+8jXzOYIZVag6cMaQX
uXm95R8JkNa4wl+q5PLtrUuM/28OB0SXf9E4ADWHGZaF3F6auir+zCxsEcPZ
2JicoxNDeu9WEiF66nd+BNc/8teAGnItMQYcvIrOTz5ZVn3mVLaWTDB5VaaS
l8bBWJfg2WHawXNvaTNsW+sTUPKc2LOyKwPJrrkoYFqKoq0AQ83MgoCEOrWW
dZjvsgNzRamUXaPGS1mqVw1wsvc9Sc2CYBTBUW5NHTzeiSgTzpeN+SybTjOr
R3dnbiTbQO89O/eoX2BvONglE7hlSpsawPkXZF0hTY/W5ctLO+BqR9HUdxvc
2qEUBZ4H23Lk8CeaeMEMtcoXs4wdNgSZpEZB0FqOnaIoLdd5TLFy4W0imvvu
8RiL0xv9Vi3PtaC2qxMwFxVfRVjXtIKVvupEh4Jo8GKGaxmxfQFHtMLqY4zH
KsynJ+X6DWHztWExrJBq2TMPvgoY5o4SQ/6FpoPu0h5X7m4eT3RLI4tQCvc1
oqbJwGKkkT6GlXCc5SgV+gkjLJ7+U0B7DUXKYS9WVea1hPmz0InJT9l+y+d1
Dc9XsWRJ4Bu+X/5V72ZtrZg1ncUJBYyZfevRbOZ0IJiVwfO/JnXq38Ntto6k
uHWV2GX9azwPtq5+gdm9Qv5oIOmXIgZhI54K7TjDu2EY11KAbQnEtlHOYZXv
aGIam46Ux7VKAT3yVUTycjWQ3wYStyEaAVHjmHVMyZpcA2xxt6yxrDDY5v8Z
J1mbYdhe5HSFp1e6syALraJWNPiMUqp1F5GtyoJSE/i0BDtEHuJDETDAlQik
q/lyrcou0gV2KOvENPiTIlMU1SrSTrGqQQZtXWH+lzIwsxEyPdZZwcasMh6v
lrB6fepP9Quok3cmjowZIKfXh3tMPbwy/nl2CmVJMRtWD5l320qaEhOJabVG
8h6E9FozkPYlHse43smO3jJswA03N0CYiUJVqJDXweu1ah9m97ZB8GUTTRHc
KlMqRk+1XTNfKX6od2koctELDYTYXbop0dhC6air7CXze2oR6t3nqeqQku5J
RlHy5elqvmYaNnR6hkG2lHwb31CNb0jBDh/e/QmP1l8hpKSdYzg2FlXP2PN7
Zm8k6OeEaUxgdJd0Wop6d2Ih1Qky+AkGTthistx12C3weVRwnq2xQqIeJkr0
yCbskMB/+N1eCEfaaFwrU2swo2KwQtVsz+gj4hMleHyNEPy83yTCnq1MO/Nz
nfGJ2PQQZ3ZnYjCwQIUD6wIPe1fDS0EpeTZIDCylX3aHDTK50TXLkMNo2F1/
0rAd345ccg9kIZyJ/LtfArdxg1NHTelFENNJ+n8klNR9ryATTEL+PCRT/KVT
0M3bZz/Cy0yI+dNmHboXqDOKwq87I8+x3iyyo2GAQksTpsG1r9PSa+/iJEZ6
+A6SsdhvjG3BGKMhUoMasEDQ9k+NJAQ47MAl+PdateBj+wdw+/a8HZ1YPQj3
3JUR6atRqYHvUxH4FbuwNipLg0qp9RRpIFXN8T4c39zuqu+3lZlx1vM81sJ3
fDiVLg3+jWfNZFM4ASMuuHjqRgG1cfTIU/DTkA+KVL8ByFo4DtJbWBt1v79l
NGTSWqkQWjOCaUMtAvw+Fkhs3JFPxs8WQ4p2znUvqL4qevUrI1Mva/gCtRxw
wblLXoXm4doRf+Gckpx9EVa92ZhQV9LPl0mUvwar23m9GVrk+Sr6T1p4aDwE
GJ0yjr4NEcLUl8Fx+nI6UNzPU0XlLpuc9S1gFmkGSpC5dHLyMr39XqVJDu0f
7qXpB0MNUnhHikHckd2V/b+tvxnZ464iwCkrbOxrkHbrW6MRmWaCNJrwSo37
Br3LGO40dlW00EfzHVlQuNN8pM6T7rlT5CinX3SUSornajcTngLQlnRAulbH
jdbZavJlIDbw9+E8vvTHHwwmCbu93e7+maUy6pQHdGjNH/VlMCifiVuQRXv8
rIrSQid+2j8qlTmWMtsfOxlWqLUfJsP33/HiByztYW56xLHQpS5u8Od3uoe9
q0HAOsPd/xm7IB0+OvcTVZAkyZBI1OFdYRFkq7lmnpz4X9QsvCPviEnhM8Wq
vaikO2Ayc44a0lXXPT0FuMpe4oyVNYJH6zmnakjWl6NiJHWmlO93L8yCsTIs
WFkiqFKVXhCwu+neIm7L0s+Ufeh+a2XRwJFOWQNeA5R/RKJgVgD+3JrtAo8/
9a+I7bO4wESGBsH+FlaqKLS1GUkrV0RyXt0/Ylv+owdXCMPuWt1cm5jnyz6H
Wd97hA7bBZroEdRFUM3pb/FVDc5peHbzlM8sVmYFKHE/1V3noU48nBfCWo2N
3DsvTp6x0m3WBZpm6pSU0mq1c+/73iJuzMkYTyPxE/jni2dYSdAYePFSaihf
vaf7Es9UOp1szc23wldRK63cPudAFAo7aPfQ0x0W4OvD/fZ4KElY93o2cEPj
Dd5brh+of+YYcXge8FhNYGKjreyMTpFP/jNdocRo8SN6Tywr6uZg1fJdfORU
EKXk6gV8kchMNfcMPxD62FDnutZbFPhMvbbMQMNOA1njM44kni/yb8usaNAs
OICmZZN3v4cJKvK77BZI5y0aHh74qWxvUvY57nhLwC3xUje+y/WDmDdOOvgz
sbHdrAoD3Mt6Gevd635kWmaVQhk+ZoOELF0Uc2+/Oo5fghApsT1LpNac7Ypb
rNZw5rBOY8P1Ypv1cyexZ3+mROhClukFfNiSiR5HjYrZWSohF2kaW7O7ltVQ
NFAa+5JItSyfIMXLfGT2xzZoKf6LzwdWtX/W3gjlu4wTJwbLS6EWHgTwWGlZ
gbmM8Elfv1EErXfxDVqayqnqdf9l/Z7c+n3j3vw6E6wYz7PQPrt4aKCaSbBR
eFm4Z6xygwM6jNZcfwp2/VLX7gOaRBXxWxQOgr9Dzw5qVCpn7oFVUBsFOLJd
P79jVwwp4ZIRdPHc+7tgdouUGjfsj/j4NS8nZeRzJK46KXB0ARuA7QYs06TF
Rc4HcM6d8YbWqjn2yPnT5FK1FxBsWyDEcb+m1kKeVU5UKC6p1UJ5rLHOMmkT
VIn4jZKMd8/HffV1yNSWyRswF12N8iHk52sWiLtcNz8W7Rtlbzbw6WvPXrQa
Y//DCY8pOqlkt5hvUsQSAat/mndj+IupehI9/w2OzoGm0Zqw/890zy46u4zd
OAIKJmPgGpp8TaowTAJ2UrGMHKkknSGmh2yI4QJuCRMPXlMqTdpxMW4NQBdV
t+11n2/QuqDbH68EyEl0yaix8He+a/wDMvLohel8v/WHxdriAnOMv/dTmqQz
T6Pe+xR3OuDaqTs81GOY3H1ofJZCF4blbFfQDMQ3BKwPHqxMEJtm443RNM9Y
vylwPlgLTk5/qbv/AkNwE0mTI2oTurM63NBo1epNHO4lfVX3J2HHI3C+2w7A
SJUA/iYBkEMYfa/Qerdnsujvv0UGMPuacCJPZygWMaxACYjXMDQOWOJnw/YH
+Dqd3itbjq1NFH/Y+DM02qSifXEVqJZENGxQ/5pJo/7fI60dI4hFalIvoR9d
FfCMv2rYIYNxgFWEmH+OPgHtbnLntWYWHldvNVd1KJiAWPGxLaqnCvegJDU9
dXczxBr0jatOJ5OkylZx/xdAvwtpGAIvFrpFD4HUoOA5dCDZcUBvmH1+UzmH
Z1Gt/M+YJWUHAxLg4bF6QfqdjlHJEzOiDs0Evaf7s8Tw3vf7Pfj3PW9zNRfT
vZpEKADqfCG+vCceNx6QgWJFQq8N8dnMlcGlfZSwtpEQf39nF2FLHfK8DIVm
3KLKeJvNuHCfU8Be2REh45V/0dm/xzTABrZclv3QauAd4m8EbjJMPg5saE23
GeiefOMiPXk87vaXIKVxkLcOylYdyMTBuX1mVrLsu/tDgnP+WDP42x5SsAFi
JDMCcGxIM9KaKRnjsFeCbSxWYQAQGsFELFflvX9zODTQK0cawHJCya54RTzx
DgCMgFdYfGEd05PTXZo0ivwn1JIBF2k4zfiio+NPNdqnBH7JCCornYltxB6c
qJaEMQIR5rLECxx3jsikDFcSo8pWiQvEvMbjNvqOEWoaRhWgTS3pt7+nZ3VM
qRHTGan5zZphL/ekQPDTMTkn6MHxRbzSTqwX6exp6gxQGRIE2M9SczUAKqbr
3nQWuU5IIujItABThDLVyi5MZHwveSGW0ukT5pQaXB+IjwZ4yDF6F0wQvHdc
71y6TYFU9Ar919w7n5IEkLrXv1pv4hsEDQ+7qHl1rfMJ4aTCIN3SP+af2AS6
s6C4CXleLIjRucPJzFZ55dkDJqkkik5E0altrYtmP44wfEnvxAol2gAnw4Mo
ccP592o5uRV7I4/5S/qqJ4zBrieCRfS0orgFcZcdQrs6dHpjb4JDTMaf7V8G
sEVFcBJ9SksDtYz48GeI++cipchr8h/j2hhNOyImzZ8Q+JQtQwCTppzS7xEg
Q/tq+ZKH2tiAuQNr8hu1a9d4+UApbv0LNNxl6Hi5nzlKJAbbs1BWzS4CWsJm
lZoA+DWZaGR839mI7PXtA59hcxHMY83xCh3K73QKBT09iit9Nzv4iV/X4wxX
NEugP18zv7ZjOPsIGjKC/ZZfXqEpFfaAA9uxYm4V+EGYkclSpvZGeVRgiiWC
DfS3tT/FLONaTgYU2ZoXykpKb3Y12PSYSIwXYonCcU/Qg/yQeUrxa4Vc+DgD
5q9nhzlUtRrBQRxWrv56z1ghs4Z2sJgP6ino/BRpFdHmRDcCqy8yoikfqFoA
R5EGC3H2KjZZ++/OVLGqrpwnk0ED8dqXQXIKd5a6VoFuDpsVXypoLbPUO8oV
r9o5qsFI+4nAZI6DG3CNFt475e9g2bi2qlxVCPH1uW51HuommdI6p3WO2zpp
KbDSf6B+aADyHi4Wl679SvkS+m9/NXpW+SP9u6OjT8nxTdU8v/huipt/tOkl
oeFwKBu2fwrollQ5v++5ufa7T/G7VpMys38PzS7htKn9JOccpGHjII5NFsvh
RiaGqYnlne/rSFQD+EVajAm9w6NG+fTIS6WPKnE9LJaminSJzz1F69N/uz+o
XWg2ump0iTv+i4SK1eau6uoQbI4LKK6K9UN+ayrcOs4xwqqK2YuFFO0Eb9wx
FAcDl4tw22yi8OvQXqw7jS4aGfneftqWR+ZLNSSl7yYmk8zAfxRMclZ2U1v0
cTkwQeLU+I2P5s+gN0QuemZrQuhP3RnGAw9grO6CZG7Kxg8N1O6kpl+yGbD/
HcBo+Wh8EK8rxv3hs9PUopnkqEm9Zcyv3SBYRK62hnA5RpmOxx23xghIdx0z
9i8gNeWqRrywbekEMgKXFPC+t76rJRXxq9sW1MMh5MAY7S+dbhpHSqjjCKn/
tDG4o4iNG9FQ4PLd4krlhd1qQvDHAPn1vtWhX1zxxW7L3X4LXrCsESspbzNb
F2ahGx1bL6dINqxlQKzGU8UiDjqqUhaX1y4gtbcLAcKaJ0yPe66KM/3OiBiD
3yKdueczE1OaF24q8+3/ukTZ7I0mPz6Yl/GXkW1umiadPaFDQ2AP8jqRTJtU
3OC1Vn4vFvMuFcLUa2Ns+iS8xHvRnmThjKniFFf0nvmEp3RfnXnosXmdoZ1s
LiUl9NLgdaTOrBdbyCE47S6SicCoys9UVRS8QWiLX8Q6I1AIVKtsNH78zcEj
/XfzJG14/2cruWcKFge6HKpQmdA1xm8J7nAEwWpUFTKA8RfXrtU44ld6bpPP
lGt4ky3uEVvjuSczb9LbutYITp39FD+tpn/HT20/UQeg4dAq34f9RH90g4hj
kE+81LtSwjDjqU7Am1jCQaGK1XIzxMK5ssbN8tDG+j5exLK7V71fg8YU8sDX
sB0FrIWnuKwD5jo7qMt7Ry2TE3TwVPk6TWYptABD8EQ5kexmdSZPDxhnLOig
Bas7SQq+J35zR1Z8in/N8OqjYK1LMuGIQdkE8xeGcEoOTpwA8lepKWWN1pti
XzTbFg/25x8RBzOeY9gTuFTQ5ENQyo7PHdOnngBly0SruW68ymVE3Wqwic5i
tE2NTUBhI+/pyXEJHAtO1HckZu1IhXV399224na72SZ06nx02mYC9kZYXIUa
Cxf9R2PD4KxO+lMtO1em3sn6MBGvvTrZP+9FzNRgGTHvbtMhjISDZ2eYcLQ5
mL7fO8GtTyjXAHd8nmUgbbGOlmUM++8rBHH1GbGMIm1iKRq+MAtt27zIG50s
gqcvqOVvp6u5HPOWlEFbn7YIqJL02tSpYLAW8unOP9ktqIEBq+6JjF71h4Uf
k6mkZlQ8eSDeaVDH7hpgdkh2H4q1L6i7R01sTqgGmPPqTiIJOsPK5Zz8DVuE
Pag6+vf53tC9kaDtMejBsoPgGLxOkXchhCFQtUt8ZwR1ffo+J0kVFGTwM5Oc
1vehwcjQ6dyBxNmzMSil1164Du6jApwkGy9ym/xiBfjK0L1+L9L8pud3Hl3y
4th48UO0nCN/vU6d14zOAORPIhTqZZ6+PY0Id2Js+qqVvCSsCh/+jwQXWHe9
2BA9YutOBf+v6sbiU1/39jZ4DHFTriSgp97CYlBhqm2irK4UBM5EM/yiHQeh
Vepih0KB3fG0A1kV6rC0G1kqyQ/c2y+wYJ9m2aFIqDguPkDr4VA3FX33EUGM
pftVjRZC+7y7F9vNf5qX8hk6Ppvg0KNjWmvw2StUVby3mYYzsa7b1n+PTD0e
aB8fPD/xBD4bkPq3eQPZvaQ3cg/TjzsrokHAtULcXdGc4Bv7rdLVsfEs7yeB
bxX6BU5zgazUA71eNo1P9L8hBbRa+qSWfEBiai0VCekDtte4l0+iwkTdzmhY
eEOHVFp86Z5CUWQbA0dTQp7Ik9/4Fqcp59mPRwhoMx9y5WI8PBtOox0iAeNh
GWqtwNt9MWhrbGBrO0subf6sJs3tBBdDM96W5Cl04BsuccIJAsfoLfTZlwAo
IBEBUR8rBjNLstZogxlSxOD1vHGoRzLRi5GtSsLWvKca0QIGj5Oi6EYfCFGu
VUowde/coJNH6LnVJfXgKH6PXYTwN9vUPa6Ll7l3A6ByluVbOieSttFjcxir
Y1qOpKy+k5wfFHRuk2uorAeUp6569RDLPZJSn1gNfVmOZ+hTnvCnBdQ5sLu6
WlMaDROb5rYV2XcuejAw8pNQB+YTXqJhMqXSvHzgwLoZvM9WyydvYQADcC1b
h6NyapgmHBTAmRqT/h/iIohlcph2AqY+H0cZxvU6Ru23ebLmvhRxqnLpn7My
LO7xWyoAJDtLUKXQRUmEQ12SPx3tZavrLo+DOwDJPWPXa012kYITDJ0KH6FI
beym6CnqtJDYfNX9rADcnlreiDMwTdUkIbhTVWV/fc28eCxaiyUuqTfnRnfb
lE87v/52IOLkowqmsNuj+5mIpl8OIhCYB3xDS5MMD5eEhy1O4lEEdoIQWX82
DOswwE3QQo2hr2wLCqw1Yl9KVcrjUfPCDUIuMbIaKxsLIG5fvijCIdBbgdez
lLhkRcBKLt34uhC3onvjFr4ESCkKnxuULiZXT569A5vhvu0bm9xNc7X1h6Us
i4yL21rDB2A0fnQtXR6Z+0lLTTYWPX+8SKwewhgfxaHm9u1T28m/8jgvwqWE
/LJYa84w88JQXZAr0gNL2LIGl+q5XkpYw3VIsyBZ7sQAFBHU+eGf3QQ7x8+i
VV+6ARm0G8IO5zdSXiIZUG2fHg5hGMu2kBhWBqva5vP7S05BFn54KHYFajVk
cQhVtEMOT1gn50kyJS8e1waat3uKHlbBsoUhfyc/HnGL0w5wowzJtSlS7OPq
l26J9j/uQQrqQdXGIrriscfFf9o7mJFqwICWU9by4Y1hriG1TbixcltN4cX9
sEOai+7vcs88Sf3ToupssGt/kP0cwZhcFZJo7mfipX/3DZOSAY2d+17J/TSs
MBD0ZuIpYDbpIqNiXzt0w5RidgACiE4WOJh/j+1P4P9sqTyftaWT8XLym+lb
Xl41rmnfoJVMt6eGngj7oIUS2xSUfVJMBjAdmksA0QN/2y+uS6bfEBAOC9z4
G0gbV7fYNrRvQYY9m0A7EAmgY42JmUaJiig/Riic6w2jut8BQ8hATA86h++Z
fwTw5P3bnRiRCNkE1Pw+gqqgrcbToKoOl5UaZPfwp9AelwJQaw5PDZK+41u9
V9BsbjWW2Wi5xAulVFTqEqE6kN7e6lBccaeDXBIj+7Z/E2BElWo4f5cZ9TK1
XFmNE5VY5x1F+wocUeVtseR1vRZ/PMMadfPjlBqiGEjKEN0udn+KcemVb196
QtKkADwXQtfPVdVNfooy56Azo2BfodGau7PtHS12BgXjYCMXQEmRlRC74fVV
LVWPawqzlr5KwyA6QT8oLJ/NRKmVb1O3MlrqQL00s4jTYP5chyLQY/0kbJxY
/m+32XLNXaxEqRXqROYkAfq1eXKw5aXWQoYVysRMIxsbuV+e9uwK9KMmvDAk
+ykCVk5+hXjCqkUDizrWNgZi8ID+YFiFMQ2M/HKNAyb2d+avfFJx9FGClNQp
dyd0fgA08o9OcxpAFiTLbC42CgqAJo9DEVh9m5Gs3KwrbEKJ4WTytnxyHlLS
otQ5Ej0rWazjUX7mDUtGWA5IhJJIhwYReNMbRocnBfQcsQQR4jV8IsA6lS/a
1wWVbAPWS2EF1lJbOIsspnQPoGjxvJ1au313RvF+7zx0t/RqwtRWHEhoYUk0
Z572RR8MG237tGnL7VcFrUNxqKLi75/5wvy8+6VYzeVTersb42CqXnGu9gep
d6crOI2G4033FIuE0lSjTHkvZ+LzBpFJZgEWfeCjeKWzHcTNIYX6nEuQtwCv
vAJNZ+D52/S6oJW3A43hJ9s1Xl708Dbwweip1fjKLB6pmWGBaXGZ11hCOEGX
Ch//AEj0gszNl7wxyONXuR2JbrB00B3ZEO258NSWTNGHt2MCHJZ2nAA1SXp3
1rKWS/zZJA6lYHKcyIt2/Bynb8wTbl9DOZu5Rm7sL8LUk1Sz+7kfq2uJgbEk
qTEBeFKnWsQYdYxiPz5ksC+3lh7ZKf+3qBYgM3ewKeXT6BHfOWQkSSEs0+Sa
lhtj4XriCHFr94VBEgTKc0X3SPOwGAMotWW4IaSZY0io7gSZlZUkxmv/aGxN
kkBbvDtJGeOyG/cAir/CjTZrfGFWtinPkmqKxMe1/q4wQIz4pMYRfEZbZDDr
ouMgz8qepBDNFLNjl0a90xLqL3xo9nqifxtQof45S4b1bcCjxicV81p7UtHS
w5Ovd04h8VYr4R7iOaNh+zn6MaGa+P14ugrfJhUbCbJeYleY6bmdHfxKNGfg
HoXOj3VFd8lrY+l+0BfyCN7wR9nkVV7JkQGMmDGAYU/h8Dz67UWAw7u0gaV3
oDJuYVsvqx8tHeJ0jPXyfC+eiW8f2DAbVR1q+zU+unlngQYq9Pq76dbEWEA9
ocBH+WAK6rx39wEy/R4JlItM/FNo3XywZtr1QzMmK51EDw3VgiwmJ44/DAV6
GzGkfnRq/Smd5r4xuFLrlZR6LDeQd3ZLZRPCxGDBLCoiSLVZxy46AcEIFYSH
KN1eUlcLqE2xhQ9d7wFqvN7xV+LmzCA96w2qeNNan8sVyRmhxU4CPivKSmHe
Qcb0lirfJn3W2l7wRAvOgUskIKZ6ZVrWShFIA9qREjcCo2nFRXvVhx7vekqO
ocdjkGhMzyGfyK7rx7YMTEswWKYulRZgwwhsxvXLP5JVJyIfaGWSEYq0UvQd
LB40/cbYgpeQRCZmSQGtgzw9GjUfGOMgEW70U+gftkKJDFltwoRnXz68enp5
/9eX6ThinjqXVNX4P9q8v74u3lE+DA4RsGKyLYNYXSVBIynyFQAIw/Alfg3Q
IiYmY148ysmYv0vWfz4TIvekiCqnJkeyiby2pdbwSbHNqbKjitdkCG3NEFBC
6tLESp5VB0JDiEqz4BIFT/O8d0AvcnpniXl6RYicEaXnqU/jLDQyTHkriW2Q
98LoJ73noHkA6ufGOakYwJy5l8NxbXm6zfJ1ju04Shjq/p5NEuK///stnBRb
Jwgm07C4vXkHKAnzAX8dpqzFWks5MzzZYeWnT7J4jrEtnKd2XEKhehNqSQLR
IZfKo3JarlxkkeOv4dXJDnozZmUIK1PvW3igAvAeqeOU75riaYmb3p7JNWQ3
m5cioCmJM41HWLqt1vRqgXfkSVgxMLTDILp2QHS3KtvW1dp7XdwYaCL3tx4I
1+DIMWgyAA+W+GjO2ISGtFGXK08FmUt3ii4KMsICk8fJPb0tEh/J8DPK19cE
XgG5wq2cyw3F9HggZCMita1SljE43r2wVyCAJZlUaU+5orJx/ipi6qydTUk7
UAp45J9D0c3Qx7PEEXj+2BtGI9BUJGUmNihwRAMQNA1sUhrLUy325GbdKLux
csNPhCQw5OfgqUngFZQsX8QiRxFhGYhKktjPU+pwFkzgtd4tt/tyGn3Xpt6O
eGZl+dVSRy9dvMgsGc2EOsUay95RTJq94cRF6pdJ+82qBQu6HfxM9/j2F/Fc
rmAX+28CXpHWMKv9hELg9lSp0lomCoHgVbs8pwLF+Tqond+s+vCaunaqNO34
vHaCBANidAKJEtkT8lVMnQpZ2kQdoqLy58+CKlS2dQwYFW89RPz9YFV0Cwxh
YWwntu+8BLagzbcOA+GYNqgt4ni+t7/UUD8s2vjZypHTxCXId4mEoIgDDe+4
QQ+9ZwfrCOLUtaK5OS47kdye8CayxLZY426xuODzc6ahooraliiH9UTJpzet
R3pFD+Cd+A3rdhFesNVgbdLpW2sNHyVtyKJ3m8PlVyd41+fDgzpx/65laZWA
yFw6bm0cphUh0GqVP7Qb6yWlP8zbvs3L9uVoll7+4Q6b+ToIKQ8LHSWe9TTE
RDi0IbIZIBGKMrYyTm2QWncztXGsvLCtsj6xOyNfSvMEPNQYnuVVmQ/bqrW/
nnH5Yk2zWnKatP7KQmCmRdjBKQ1df8npSczCls8t8LTnLwZYIH/kZtp6+9NG
EexObM34LG+k8hNmDUEvhiKVI9/HdLYeHSMkV8JlM8b8d3l790SyrD0zUw3A
38y0K3DgaOq+Z0X9/Y8DZAoPqx9o7vF1XcrOqu15y6XJT1EkrGmb80ruBRnl
3ItHBFVL7Qm7Lr+O2Vv/RP/euyEG1ALlY/4Mc1qmGYX6uK1e+u0ULvrMqalF
z44jdng5snqzPsYSMdO8x+oWh2O8DG7qX7Vu5xCX/XZ7t03LY04HjIqYzKxf
cQ2/zQy5KMN7SJ1dEF0C2ry4K/PguiQZiU1hFaIqOoLUtcUtZMLZGYYQa4LU
108BvuLgJYd7J0hXVbrrGXVCkcQGeU6gM1zrPjHYbNZN4fLUQkVEidY7nVxg
70CLsvPVjkiJhxIl5HqZYQ2deEOHPOTWLP1YZcK5UEKhjQX4eR6hAnZjEg58
77vGY9CmJ2+irDWooXMWAsURLakYNnWDneO6E6nSdPZozMN4BF4v+5ZEEpMo
ovIZaUIBeyFiB8OLQQtOg6PkbWljx7WyFASA8ERMg8D7j9m8bvEsWua3nUDT
4T28EvdEoEnTvFOsLaMJBW4cVhE3BqVd9/DaujJsTO0D7BczbMC3AARD/GBb
VPcnHLltCd3CCSzJKBPwPwZ9HoGNcFlwvigVRN2ZZ4hZN/Adro2m2EkYAymc
hRqEQ4kVb7BLqpb8XMn+4BqNAtAcC1k5/9HRNsullBqeOrEzkVgJSmyW1Drc
wyRg0iIfSenV+5cDJxS0DgVWc8j8j4gDMUrbFCQZBiiszAGMrVgQv6bM0AsX
m/l6e5+KbpFHGoZ0Rq3M+U9tN5KBnCGkN5taE90m52ataovPh68/m4psiL24
JTFEKSQVEKz3jSIBFrmkxF4m6VXiJp1DrQmUvAulOfDJIzjoh5RJizMtvNxL
QH+gKzkM7oU9YzlV9h9MUZJ7YAOI56G39k7pVlVCUQku/PS9fk+B93x8lRVO
xDWYXZsB6UDVquWNtUj8NGv7RPj8BjQ7pdtKMgUhxbYXksMaIajytHOhS2Pq
3QCzSGZLFTrWAJNghowoQh+Ucru9aKctK9145lTqLJZ656+GEljyg0kPVoG0
s+H0xpsI4tHzFfeh82AHgEUkHhp5fXYTpoa058SlWF5w5WKYlyOnNxbwCXN+
3AcZSRZK5j84k/iQvaKRvvvTghkopA69aS8ydLyvJDFBan2JLiR9Q/RO+gqJ
mOC73mD8HtiFAiRHFP6S6JpVI2sFN2/6T2n4ApjdgJtdMKqoi+5ZZ2DLYSYb
btHIZObQFhgBcJjNzt0clBrRtnwvLIWAEuTPhvWF2VkLb66be4W8IhfLaFlM
Enmim9AEBC1vwVB7z7OiDLzgvvdD6Vz47k+qUmGa20ksv0YmUE4KnrK5c5I2
LiCvEzswLJ2KaEsc4TC4dihpNle0zhUeBHDLbG72Z96Txd1cnHdwyh19C/wk
V2+5jcC29rjFH7XNtUwVbWDQDz/P9m1o8osn+2+tehGBdmkiDZrb6loFX9Nc
KLsBzGUKMtoERtq3DbW3+gftrtEePSpA30CXL9yNwM5NZczReJJY1kv3M4s7
fFPr8pD78eZXsjZ45hZel0gUmXhEhfY9lTfbSqGMIijNARN+G4GHpyXuHx3L
M9tkLMxazr6YWr2uatOsk1M01fNQkUlI9DJd6eUY5iReF6AV0uBlEA6JT6M0
aF616cT5lEPWPy2Bzx1ErkXlV0qFGTh1sgVRZsrS7mvDEFzKZgAP6CkFhhA+
ACbVj2RTa6PEPmf6DCVYlap446F4Vc+/tiQpzo+KVxn1jYMTWDNIvB3LCrnU
wj8U+dTww+GdiSFdUxjo9yF+xhALVQt7BUGOBBUT9NS3zlX5yhaPI2Tg1Tlr
BYNS7j+/ULDWaLkCT2N5bTJ9SYc5VP8fN1ieGx7bgI18QF870O6J8iSfeFwe
QgfcsdFKb6tLDldY1sSrTFX7ByYSj2EFy7W5uspaKXmX1p2whgAxRwfhD8KZ
Ds+9TqxFw9+vvaoaKjT4TNZDcSOT59VSTmKaHloBRROf83X8O2dYb7XnI7xS
z4EobAupu4DfXuPKMuYqq2H1p2aa4KDbLULTzjmK2rpiDS02ky0a+QZt4f+U
j3/lA9msEuAggEoi+4IeCoklSIDHeeS0C9hxMfYfHQrb3QmUXuxWbfxNkw++
2knOcSnQrJ8P9s6MehDeReMtfTwDWmGa8nn8TRmtI52gs0AOm1gGx/X3Kbuy
gMFRoCU3lGJ6FadEiDrtF2+yQgP4EDwq/KtZ6eiTSPbK8ZgkurFN9n7quJLD
zVwTPnLsvR7sct8bOJ1q3INqNN6sLI5mipZ2OC37mlYbmQnSh+bomY3Udr7Y
NofYz5wT9Aco3lcM4YUUzt/GyIz6PHWCBjZ5/eDvNDKdgsfsLzRN7Qrfpt5c
H7EGdId3cuQgW5N4NWj6YQUSQsqtm4P9wRcq6QDiET9S5lxJ9ee0yL+9qKmU
AvTgr23rc+5S21DHYbYsLGDanBLo4uZeKfSSIcIFgJcv/hpZfcVeP0+/iiYq
Gnt/SqxUQiSYMb3furdXsOs9FIgZ4sK0CdYq8pTiqydIuP9EZmIfarEB0yl2
jdcZfYj6TiXWgCVEl4UuI6z+Nf6bO2f/UH1GyyyZW0pX8noqyl4lpvmmoYAx
noPm/lSvQBnEvdyj3j76+rjsvFR3ahBxdUGLkiBz7I6SUOR3T4xdZAP9zC6H
dwpCiYlwX5hsrIxVhrpoqK3TzZapR+0J3uyvDJ/rhTaRtyOIy+4CF+o7fZ3b
2aQcJiiUaA2tfALbEz3r1ydxE83vvN4HdkE5gSbzkQPxV/Qj/YVTnHX9dP4N
OGngMYgG99SOnfwr/DZIdbR4Q9jYxG4uctsKlfoBHitWS4zlvW1FekobeFpu
guQZco9F69yxsFVNkQ26vRBFjmcGeaK0y8nB3QRw6dwcOw5AnmelKMg6jbxS
k7UZNsacoIRiKjGt8oPOieNRJKudNXHxdJ3/zri1k5lRRIBeNhVtFyFdsXkm
Yhei6PF+RL2jUwx3LLa2eA+DTGukdcKwxzTcDVTyKIlZdSQtZzLN4LI0yLMB
DQ06OT3Vg2mJFex3aprzRE96JCG0jbAySpLgwIX5wSsSsJBbW1CBupjyDBrk
Jm0my5l5a7EtiRZHmzj0W1kj9cbUlQPcu6Q5L/qTmZU4sRhgYCsnYJVRlk1I
7doeUvfNl7A492zamrHlmnHCrI0IMX01QMNHEi54phJ9HL5hfQhrievozr9g
r7b6zpP3SxwqSGL84TPuWmVhBtg7h40jY6zfz+oIjuK8UFGUUiIZRN3nCKho
kvRrE3xwrQkrcIT0dNPGTjsMBQyEAUaUwmzRYskDsTB0ocberEPAMhGM73L1
CWdegiruGZshjkqUDaSZJBZNNuimbDCPLKwiMgQIf5SJr/ql+keyd3imiz3e
bzjHa2VkfqaIxzKXcq26NlqjC3M5sJLTl4OB5xRFQUGOmI4/0MZC8bnSM+eL
7rUr72GGHlzejzYBCcCA3ZNmJnzBCbMYxjvf75nDwaxSRTA/96151Uv04a2R
8W30cc9J3C48IfKKpQy4AoIbeDeK27+W/Cb3WiEyPMFWX+h9D+t5KlCKxGJQ
F/ZVD4F/ogxzqou0UAo+utML9j2K1sym1GNpohF4uk6OTyH8j74omtO1Ap/X
A+GP5raDkTHim/BAImV39iqZaMwZJ4XiYrarKl+YRh0hptx+JIRBOnYdHGKu
YgPb6nmP/dO5pBO/S65FW4eSpAdOWS1BmMn7GeUNfqQxzDB2Rg56UhgkC1Tt
A05zEV37KwLQuad7g89UN4C1Qk4J5vnVOkdyAfsTdiuPlcdogewbig4H7zmM
9qXCvFz6spaKKHg88IdCsFjveLx38vX+PK3JLoYXl8muumnvr1ZYyWVdPYq5
PgrdSa/q3qzPPLSnk7WspDWjjSkJjzEHEQ13QbCWs1nzvWI8CvNloqCRUpDi
FP0LW9muR8DUwWFMyYBFFWUQ2zkgDvWpegykBiyB3rPKyDj4Xv/k+rzS6kCj
O8ph91yuvQ8ELXz+hFUeyxm72pJ06AHwNO5LKALpGr2M+oj0EaWUsqbR1/uK
/9AS7nLfOL2B+eDP418bHqPk0acmHhFWFzXlEPst+WiBXNGKx14qfPpgh0M+
PZO/arWfj801LmqRoBrIHGgrsBv5h20QB/BNwgs3rhQXtAjgkufR30L97mbm
vHOGdV7nuAUG6Kk8g025dUKEndlKB4SVgQV54gOdi+/Yy5j2CmJkqyQ5EpoN
mQVRSPJ97Oli49NofofAND0X61n00ArsL5e80MRd9rqgV/4OldWb5/XriTq2
9W2I+g2x3aDUV5F8+LlzXIKylTKqkrpZyqJg+CMSrvhuI3paWJL7rQt4ty1Z
ao2cnEuhd2KiGvDbTaU2H44HVacykzCZttmstLPea0nJFqP5tFD+6cKTGkQP
5PRxTbBEyLwwd9x18iQot2DsX8f3G0NDnJOLdFqNx0Fl5SKzOfbTGIz6xVVA
VBgCNnmk/qMOamOvnFcckiCI3tqPTXIISnmB23FZ2TXekE5diQqRUKvIaAeq
xrSaQrdAv7v2Uh0HPVTv1zvqbr/5elEYUW1e4p7cWfLpFnpQOC8w5J7S9fFC
pHwMbDUaqkjGcHkU1/DAadnww7UMFUYg9cCDc6VxxX+KeQRCsctht0yvfoeu
/o8EIjwgkevweETp0auyy+JpiG8F6FFm9cTr/VH9ttwzF2ceYYBoNnKe9FDC
GB3ncV/wXrZYJ/FGEN5vFyAC0cUpzgxoJqumYvxoNBKoHnFuscpkSF549DaU
q/pEwYLNuhP1i4vPpQM4s2dvpGLdf8nitF2rHq94fekDK86n6M8AMp1eQgJx
puid7YuKyhsZZhfxAzGVvkwow/GtkpvOd1gjKjd+nC6TVAOf7fjAuVkHwZtZ
o+pdn0Toh2OXSP321ekM4BIwf3kKrVrARkzW+nD/THKMdCOqzBcpodWBtJj9
zIqeguZ9Ct4cwmm0j0yldRGb0XVSsghHUNHd2VLcDXFtziLe4E5rOR3FiKEA
B2zdsjQXlNU3wVrhfD9vZBKleTcUWs4iuNIyhH+G+0MKaWjJ690KWMye+fzF
j9KtPdeEn9WFW9CqRmT2jdlfz8SI0U8AWt7MnuERhmsSB50Jy+keEaHm6BUt
11TjnJoAVeDYozcEKX/uW3ad78ihYlEcEI18r6lBUKT9JrNHSLiF3Q119Clf
OJT8+Jd8gPniRtqbSITjXBd5dPJHyImqQKbPiaKoL53I8XdJ5ExbQM6U8y5F
CyIb6IONDESIr2/vPso5Oym/rPxE1qChBekIxJZ0+pvNPNqxaJGNxgVpKXZr
k1KOwcfM8kArpeTzFOfxjNPLLiSB+YXhYtBBZQU5qk2rHU9oqngwtZAXbRmW
JHzXKeL4drPSQcAUaf320ix46tlWUmfPuoLaa4pErCK+mdbOBC14o57X8CNI
itt93X7OOlJdffd0CK938rY6m4gxkxxYTrX0yT69Fas2l21MrRnJCrZF/SQs
BpkCtraEt9ZHPfYqc18I4JM3m4EeLqWVtrFQKcqbIac18MqhT/Lpsd/KoTmY
hsDJom+n2IVWRezox98RzLIoBjFfprddhUq0LleJo/d52gvGQMZkm+r4vsRd
p0ctP9amQBKCCvTw9Ayw9DBtOuPy4cNOhDBMBp0YiJX7nlOCIcALJ5YyRDPo
oMy77DSPbDk+ohsBYVnO2Ytz1onNM8ZsKC5uT5Tm/P3FQXsP70nrqW1T0b0S
sl95eChILg3fKaK7hQ3+uXNTEWE5jktKeTn+kx8FIUSFttjrsHLEdQgL8A9r
elBIMXKGwcDW/WmqZwijKZqh9igQQcyDtjA3jkaF79I3Afh3OYO+9/VRVaG6
WrYTPi94FC/olqIaHDCHhvK+0+rk3qIcyL1R0VMHVfx522OTIpZNVM58WmRD
LTPlfjvVLhBfAjpyvi6hEMh1uIeViGaUoi/gCzBPS+5MK8+dVEV8cdImKynr
AkfSZ21w3AHOjbMJqm9rsEgGmpcKUfzDn5ZTg8Fq3/DQ4OxC9FGokhjRAdnT
56lbogCO76VDdB4t7MTtWQM+ZI+33WBTeXMmA1hMUQgz2HUyOjWRC6r7YCIf
pzfg39mrar8F9fE6ghgyqHGMI4M+UoDosgh3u2S3+pdaEc0DC/nPjr2Au/px
VzNm0MV0thpduaGLRBs4bWb0REQlzWhUv853Oyu47tpgojMmz4HRw8ebxjeW
hITQBsAiRbjYP/sLZC36Bi9pypD0Ka/d2gB/7MPw1aBisTTflqDcYI64btSu
Ivfh9Jec5Vq96Vl/rhIsyAN0l7rEBqxDbx2rCjjmjGuGrTnj1ffFp4Q9uRNT
4W771/eDxr7q3RyBwK6vXH3f4xFrIY2wwoGc5YTk0CQR3zauaelWyJL+hMkG
0dYB6IS1Pmoh/JAsZq0go9cMjC94drO+xlaV9Radjo+oIfrNOmL046gn5qAY
GU/2MQpAUBnVXk4XNTr8JqfDSIsg3eOCWsPlOHuv6+XKRX4FwR6z0vW2lMmA
liK/OVCuc8uuXm2fDvkaB9HvTOc6im/uM2hhUL4IWfelqllW1rJkihHbrKGu
Ve8itKWMVHukyDOGF+cuv60HBSwkvlO8762ewt1yCX0I5gxT5kDQnO3ev2he
zfK9DXn/phXhDzhMaVMm/7q8gYqmAlRMZEBkp+MFRI/W1NWA97tfleFt54k1
xpjFuTKWWjSr1xoNp09gEFDTx+MB2M3pHm4WxTXscLGrMr54ZBCtfVYNeAVk
YJuO5nKuU0o2Ut7SOz2bgEyAd2L+uxlaiFWPh8DDk7E6ChDiuBP9Ue1qMslp
2mLHgJRMYAsUSu8nHNRGW9QsqHdYCSvSQIg7Hxj4CBakHSYXmMp8sb/tnYP/
k+N35+IJ2YGcacndlJlVUZqUnyDLoiQ2IGXNg116fsNmLyfsN+JO8yeQgenS
4ZAoTXDw6lc1/qwnpdJfa+sYONV7qpmcBvdrV8Z3D5V19U8z6vW+MD5Ksl0D
E5GvwfjJNgJzBaXup7tK2NHm7u3Ncb4tw1ZtGDeoEarELzaxiX2b0m1PWUFd
tnoSjM9Vy97nufJ0VImvUOTb4mcOzaxkJhnzGfuU4gDY8gVCo6CjQipzN0Gb
/Ixm+N48YHKjh0NnHgykMq1c4/hPIQdtuCZp9q8r829/OEjd19X7HW59yBMW
MTMMJhZdtstLWHre0jfaK7R5WdVEgq4FBw8GcDBKJb7bKbnril6pdBLiqsyt
llExen5XuKDj8j0E+RWXfObhFI2eTjYgDsp5B+F9R/VB42nNnAG86YCzNdzy
ScxFXanAi4RYtYsqe0tAo+a6vyGmBDi6KOmwYU1ZuysyWjXR/l7dtiDowJAE
2Jw+M2v72LpedWyeONKEFBcbxJ7kuFhoLs6N+o9kvpWJYCgl9PBQ2oNkc3n2
Rghq6Dpab5e/nMD4UzlaunuxCb+ijjKC/PtvL7clxAB5+gxdn8HgciNMPZ1L
yPbcZ0loj5VOePMqBbUfAThyFh98qBlMu3lf4F4LfxasqMRlZ/ekgVZcx9hm
5cqaX6Ptyo5sayCGssrKAUZWBMU/sea1y/WpuByDoVTXmF2xNSSR/xYITFSw
psQSXyli80acWHX2rupVNEmEcSBLSF6SZOFW45yUB549MKrR5cXNHqAX22vF
4ubS9DbhdnS9US2BXjhqhZOxKjflT1YfdTy7AtXopSeH8GOtPvhItIgCf5pE
sXgutPhVzWHWTUaOsq5oLtizbVs9I1uBa1tsAg/g3PNkmZqm6wR7rpARJaTC
4TvKegyDYseppa1Sw7uAm//1VjpTob2UUuWybvpAIb4JsjzXXWA8EaTAvpDL
s6ZpDno9e0O6QQoZ9C6qOQEeY1IK0d22+KIx9MGOHBNPe9OgOxh2HdM3vxvK
vMn4ZDeuL1KiX70Pem9mFeP/ppKRiwv/SXmiRkZNiItj7Re0qpVwxK4uLPAv
YaD62PCKJsFiYVXnj4ixEB8A1qdLz41VcI/u++xlK44jYHhKfbgAQXrdeRPV
gFBeZLNNbql4fIiZ6X6uwoYkjcNm5eceJzVH0jTvAv8KfXBr/7mv9Y8NZrps
qDeeko0O10OgtQNS/CaLqoAqlYKSlJAU7lPRH0yiPwz2tAA+T6FRBNOCormv
jiJhsa1zJfvJ/72xnmwaAQ0cIIXIkJBrq3X8B3puy7Tr5ALrh5wkOu1zf7GT
DzjxZE5hN53Fb7K7H2Uv9/QKyu5NW7kD4uxi9h1hQlKaMU5d7NFWujz9VwlA
E1ETqGXgYblbs9KBhUa4lCnd1swiQZtHlEHvAB6kBKJoe7P5AYItsydxvFtN
X/2Uc96xRYeisOg+oUFtyv1gnNRKXS7YArkOJZWv6OFfFjZeCeask84eH1cn
Sxy4lyjX/Ca4GQA30x5LseBoME6P7MbLGJfhO874asGnjQ3lnlcV9YzDdhyh
oYpCXwBzhHCYriFX8JSLocGBNIcFTl2hi4OQT5lEEEP40Yy3CyNa4uBrafB0
KbK0ioT2D1Gaf7ng1paudULBupo0h7De3fbeQeQtIytPBiP//24t48xgZife
0BxLYtaDUS+SSLLj2/euqmgEm10zcdA1Tv0nAHYlCvNj/5doE7iuwsNawP9k
waNiMOtxISNDX3tLtDX3tC7habIZV2CWRK7FdKfGTM11PN1wC9e63pcleLUz
0jrlc6teT2GYq48bmTgQvf88qSm6cHl2TRiEsyu+a2XGjRbvTc3le0o0XTGU
ahzYxMVo6URBUsaTCM22Szy/aFpb0t9zh6+uLaZ+fpaiCAV4CwzrhgRoulM/
qiZ1quKvfcF/bLEQlyLSl11ZBbjAC0WQYkZ1+IL8hXutgQH8cCyf7ZVgHgpa
SJdKR5Dzibmo5HpZduuVIA+fNOZAdURnQbjd95Agl9ocdySQIEX8fT08W89c
vj95o5VX3EAf71WE3X/qxTeZhQi+2fcgI2mj1QCyv6KNpq7wP1F6V7bMR4uv
2ZTYvje7fPPI5UPNfpHE5eYAzqYSZBkQgCGCcwIX3YJFSEqzIXGIP1fWytMq
ZwXlR0brcoIPn9PBStqMTvM7IO/wlLWmY8kFP4EnheXifX174DhhgPhhVhEg
0kABONWa+2Amo6GclUja3o26jC1i1uLpyIbs/8DjQ50UKWW4Nrbqbye8JuAY
FEpe8ZkBXqXgKOoNWI4L9HwyTcvGSybZIs7GboMp6X+AXXoeaQXbk/Hi3gJC
ARF/GHNWmknmS2Ke87ym/5ka4v5hUKAktiuEwf5lpdV7y8Rg2cuRs1ilvrxk
rCsSkXg+e9me8epT1gh/L4KRndgbvrU+6itTH9LOjcE2ZmMGUgNR1NGCWhZH
YBLx8qHrqWPZ2pPVv8gOMNguPtFpfHwDeP7DW0Z9/JSLc3IU5GdF/A9dcUN9
eO4rI9qyF41ZBEn3hHOehxXF91dQ2DnswFCKRcB6PgRYLscctLNzX8hwXC0A
exSLbWFs7Cv2cmCurBojmSo5EsvchFsEFeTxMT47KPWJYUV0JuPF7nviU+tQ
YrLDduR68Gp+9Kog3YUIoTXEAU2v7vEXNIV1S/G6avF18UvDZtdXueMvM9bT
2UCLSba1dsWXb8Ceskn77B7YBG824XoxtoA3PdHwHIc7RhN46fIp9c2xk4p/
PR8NWjp0t2XNf1+1jWtv64nzw0HOI8dwbZ0QgzPhlAS8lgrnA3LWzF9prs/p
mkC3Pfne7x85eWOoz8/vxtQiHaNaskSHIi2/wN4ABqDQpltq6+1cUDdyx9kG
GWkmI9bc6mR0ecuZJxAQMK3COBph7g09D18FKH0jXhh+VUJO9TjW1QgAOfDa
SurpUcBfh+ege5yho3fhzXgvECTcvk+ScfBrjrUVLb6CYFF7+DvtNf726Mln
gHHpZhhdHT9B1g3+5HC97b2o/rrQb2bBuED/H7wnq7enbTGclO6a5Z59PIiW
n75gJsVJvrslxGcqd2+nCROyQs4YM2PaeT+bW6gjaQbQyxowtvR1Pmv4Smr0
ncU5hJmTXNhxSaN88qEP2eSv5BgVqwBEZzpVEVHHNYgetC3LVTpq7WK0F7kw
5N5eLWqq3fsxW+EMb1p1YnejgJEwiARo3jxnnB4FMlVZTGcOKOnNjG1zTYZQ
xHpkqUc43xsXSgBrru/JJdcSp/X4xDCQnYTiwNF/ShvIp9o3oFiLapva5Kyu
X9CZ0jAv4cFV8WXJAHwWlP/il7+OOo6+lh54wWcA+yq9cZhlqPksQVbyIPgN
6J4IpJsPgjaIOa7vBfFrlsl+6lqpQk2wLbz6V0qJbNN1M843xpfLMGarVa23
HMc261TjAY6td4/voWd/hMTLZ1OkAXiB4wyLQyTIHbAANsohiUGm7J9hrh5i
HsKnXqGAc7RDjuE7sBXmQjf4Xo4/Q4/2bkZHDlACzErFplFJZIJc9oyODtKJ
fOn0LjwduMYQ8RmYzXXDKU8RY3HoqflENjNmxJPjBXDyJO2oLWG2m7z+cGuG
0l77haWgjgm1LnX3onuPybbVY2TCuPllePs+bXRLC9mXA8fy060Ed8q3cWkN
s321H8RDkA9o01WyxyOL4Od5rfBr8aHuURsg1kHnq7wqM2nOihWZMYZkp1xa
qFfsZpww/qXK+hR42+2XlaS9rjxaePVs0oTWi5QuwhIJ5Ny2SMYI9MQmRbLV
OSLxD1CkaY8Vj5EMtJkd40mWrRYY8mWklRg4Qc668xVmWypSWmsc5c27784N
E8J0pDLnQUa4JytdzajlGD0Cm/YVqFeSy3EOb9hQz8oD5xgFgyX02QvCBe6B
Aoc18b+OnaG/tMy9gj3fwUlIKZPR1tTFYh+eGbdwxVWTB2AkLOAhCFFd1U8f
ZvNgbBcnr4f+yI5NH9ORY52ULWNNr+TwpzCTSQz4k7uqvVjNx1uUsssRZaAH
8h8c3oEz3rBPPHx7XBCbYioDypG27U+kqb+oPnhkB3QPlPzWWIOiw1ubxuME
cjDJSpq/xheO4WgmonOBxKVStLJMpX9nqh8++Dnnud4RDqqhqssbL7ALqoHU
19n6LgG5UtwzYeuzFaRSR/f1KnylMuIvOwvTzEpYwScD8Yxj3R7bKlJGpchT
G8LFaJe20x2WUWEBxN1blacdOlfjJK92Tt3IXBGuvo1MJRplwjg/tr1TIVBS
HHxTG1xpmL9XgcTzeTD3XeTpL/sXBHQE1+PpWJauWPKeE9Wk8OxwrQFvMi7r
hkpFpQZONjP8D6Udm2tJGt5EimQzxV8YP0bZA3+xPgTBTSr4ZAYhXphfi8pV
Uy4c36eSZarfzjadL03+1ZGwToMWD+nbuyImhhptq1F4ExdgR4pUCQ/l1TKp
O6mcklxRHhOBAk9CNqwKcnT63NOtqqxdfaUqyIXqfv83Os8TqUHQHMpvO8Xb
rntJlX/uAjCnWKJ6QmXPUhm9AaBnTuXYVNpNIt2TyZ7qzcvsH+/pEH/4KYHO
3ZwNCM6+UkFTUfJtm+lZcv+w8gDKzw5XrQJkvQGxiFrOhAFlUK/zIvt6GSqS
Hpf/qu6c0Pmj62QVRGfPVA/3fITS8e/1fEEqniYDIIelmEHiLZv7twdxrAne
5mLKPfPOk+zBX7LqBDmXJ5oe2Rh2LilkTPfmqxEYPUru1HzQcUH9ZuEhWwf+
YmdEkO8VBVUt725vTu3Du04yDh1yp0R59ltkeC/Uy/+HEmSnZP6jYyaUQm2K
DUnjGt0WEA2pp5racHv+IChxyDSZm7lfcVnR0zxnIYL1cMGmK2n2N95wPWqB
LV+SPqfS9Y3qWRhFDp3IS9RRhDhet+Dqjr/H3q3lxZBD0w9H/fRUejwRwZB5
+eGuA8jHPMeZQv4ni9adaAuJUldt2wBiOJ31ysqmyndM4rlqO+cD0+J0rXL6
/2vIOVqUo8jMx1tOHbj8ZISZTm+uQfnrU8fw2OZ9BcyGHqpYVjFZDNpZGyp1
CLTX2kqNfHnDXS49o5zi7gtese5BP2wSBsodiL0Nv/+7680RztjMVo4cgWTN
0jmApUcGy210dW+d0QMIf8z5mR+t133z3Essq48r+k/I6C2Qsj6E7hIgv15+
hv9otP8i2NtuHYJEWtRJ/67DrDSdi4muVeLkejb4lD1zTTzSnU3MWS610hTo
bmLCfV+lW+WiUPwk2jo3yBA89PHT4FigUtf9JU5f9TdvZ5q9PKFeB48xdYLD
49+L+lcl/y/eXS2F8ygrdEcen2ppnpl717200Vo3aF12VEl/DeTR1bee9Ckb
pJqZq2yp2O6errI9ei+7L+PSoiOiUnWAMvqMeHxx6blNmCAkR/Pg/S4WVwfv
KjTtnp5BiCrRihJfWwtWP2/qfqQO0XTcsAyn6QIlFUpkKi3rvrJRxFilzo2B
4KBM77bf0Um7uEIdBCRtgbVWZCdSJ0nh6QX0rJ2gz0sBG3SchuSjvXyLi5ZN
WGzty2uu/ySSd8o5w1Sj1WjV4P28FSbFJ8sgQBZac66Vv1vMTYdcgwZpSoSW
aJdcbCzmRMtoMPghnPhY+6BRBtIMU+gxYSyyE6A7UP/7ngbyKRlCz5P8KhAA
S+5DKPCtKpCOsMpyaV940z24gX98bEzusQprJUoMj3qUsQjm2DjvWXgPsI9Q
Au4cyS90QZSYMJK2Gr8iFq923atMVcI4PfWeVqUTUuuNnYuFmdv6JB1mnVcH
IFGLE4U+YqLHQG3Me8qiXS+OwDDnDd4wZqTBa5JMNSukAch4v1+degiUjvBm
XBOE9zZGiTytLQcf94Fi5J4sEMyWl5IeLC+493IupvToV4HzymYnM0kVFMk7
5TX5H7zpJpUSvDBosmfP7C/Rsdj3C4kibJ/nchZ6Viv8hB9qfSiRfO0r3UqU
xk70OWfgZ7U4KTFHHvyEIgbKEByJxdnbuvtFs8weAtpXNYrKf9BSEyiSGlUR
n0cwB93f0RQf+r52Ur8nVq3GVv27gAAnr0CL54QZuU7K9Vx96EkaVo8HJ3OF
nGCD70hEtJSHugsJj4W56pRkRJvEYvNFR6eZXP9du4sCGqf5G1R2qaYPDlf2
dLCbvvRvLfcyhjclZiTDiv0GfojkfA8gNfewWHbc9aHygTihzmZasYNz5k7k
dJI93F0zhxxPApMTc/LilRtX3RYDoX645+S48fknt9SvaCBqzKeM8VqxuFS3
3tTlkiWAHYUhn/lys3+GV8EQzJLQUfRKMXT7o+8HqsVuyeJ7m5PuaHa3dyLs
652WJGd8ub8ANuxK8b+LFYeLpwn5N/YXGK+FQOnAp5fErpRthkG+kcppX5nG
PrAWQtPKpp25cgGFkCVjXIrJvvQkjl5gK7Gj2mPzc+OiSQx/ulNXV8d0x45b
GUP6YWgmTXZwzkDglosUPxY8euvykimu/VAd/LymCihyQQJVE4VFCswUvwUd
U+3B9PFb0lbOHHw6ZTOyBDzpFE6O5N21zQ/HkKYy3BPedj0V8c4M2ESxGYG7
YYpxwq/PqM9pCKvddPn/eKtSuc1J1CnfFulEnTb9qHPb91ynHa2B+6U2aGrh
iEySHBCbeLT/Eymubc/H6LIHPMrMyZ72J+KoMQ8APKwQOj+IMLxUiJuqzYAc
SqB7utqiLPHJBhpNgSkVINAw+OTu48nC1Vov2u6a4drb1UUnlG4B16r0H/9C
tJRkhQsukfYHBb0VTZRqSsRB52tDVZZu+/DJghJ+VE0caslzpvMqLJq3D038
vYRq14RP7JYqUFVyvWjeYwOBK/NUGM1IDGLON0mGIePZpZmWyTtowJ0HXr0E
wN5SxnSHiLzIKLSmpkzQgIv0qf8bBgtAP3+cXU+bli8Wn/5I6xuH3RfFJSzk
InJLc52BLpA/lzMqw1iBaxPvR9rkP3a1FxLu4+cg1Icg3O+5W+AcxVCFq8dm
e9S9y3Oy4/j08pSpU11vnQqSVMPvGM8NQy4PM9KyxrbDNDeSO+HiWz0iigIp
7TkwlvLMIKHB+ClKEJGx9AOEsLXygUC54OrrWpHDukH4sPDN5O9Hl8iEMYiw
kkx5L0IWn+zev6AC6GCLFKrP/TlmNQB5x93YN+gOVXMmKHr6tDeMeC2Rhkut
QHodjAPLubehYFb7wkZn81h25AMazV0qh7KkYPxosH1gHjaX4RiwS08uYM89
9182jU5TJJuTlOfQpSiFn4wubCP5lQQCxuA2wYF3S7EAXT3PtV/C+uEYI1yT
ysYiwYy04Cqc+tDFVHxRPoRqa5oyQRjrKjVRoU7rADCWJGfAPLCLzAtJ2DHL
toHdWmwiJ1SAa6kcRxF2K8SqD7RW5h1bq5mJZ8QNeJUQQBSraEUG28Vz3xEh
OuwTDk46bXkONhtzQxeamFI6lG/Z1KY/r0NexkV5DKRBbWDFOqNXc0GcWnG+
uyjLou4MJXHfjbvL0FrV41D8GsmHJhnYr96KQ35BDosFb1I//Wjp9+HDdhlB
L3fEKLr46HcB6SmngAbSVtkNcWi1Nkn/2EHqPy2ywvCSQ4V9/IvQ3FdH8Qcy
pt79bweQFDetIbGD+dC/X2lVuIuXd3C+zRXU6TXjgCfUHQccneY3oWL/cvl8
xIsfJoEOzs8wlQo5O8FR2ORmXehAveRM9lYIhiZ9wtqFitefl8Glhmrk1bY+
VP5ggJE5m7bqu+Ua0b3fHjc1rKRP8NwJlIAvdHNAaYC+jWmRCHpP8M52AyUJ
/3b659GVOkotFBysYqt6P1t5DtGaSUhoAQfSzlVXWLkqugU9NkT7cQgZJONg
GLWNF3MLD4v+WotFz7SCGYueaqtBbsAWtz09mWfZsF690vm1ixIbuVO57YZW
5FTA6DGxlukztQ4LiDbj1xrhzhnhJjqmZnOD0pvb5cHSRB90GCMT4izQeVdv
RUIqwfPZQZ/sAyVxzrAag+rKxVqxd/c+WkayvXqnar3jQAbeKnlSTLTmBt3B
V5gsvziEld5IjxHv+R0xOfGds8AzFx/H3HNbLrSbkGduqhQmdVFtmYqQoLoN
pj1GXBWpkPGYxO11s7nVLyd8m8Svv8VF+Pi80vheDZhBx2vN5/TR4RXgATqG
WQKo6U4RfIQ/hojDpvkr4eh7LvkUqxTTRzMlPnvPof2Yasj9h9utw5zitO0W
YzVBypowc+TGFbOXHlX+tSEZHLQXcP9i0FzQVdG8RJ0M0Dl6XIX8QdBM9h50
4HLI0aSq56/3AKuiLf5MspCQvL9n9k7bllZ55GquKye5AHt0H2THtyVElFVD
NC4hLzQQbzaeV03dPRtzI2IWwqfOHmVfGyjK5DNNs33nMK2Em/zGmGC3ngT1
7kHTKzLakMCSAxGzaTQSb+SMAmMYZCHGKAza6Y1bsA3Vx46RTErV5oNHYK/L
6dQdAoYfk+UhB/NMZ83o5oJKMoZbUzjfG3E++su4L1o0Mwn7W8YKz0cUdB3M
AvEkxSIvkqNsHdyKDRRudJwiZLZsjy0hMsmnT3+YTnalLDGsbAGNwY+V/47j
8i4tcVCXRbWHYfDb1whVGMcQLNA3f8XRpcQIyySPXBssaZ5Se7tOC2Bc9QFn
XUthrPfynBYhJLfOF4bVOyJdorskzt3c7ZbFzduY+Xh5XeEivnITRmXNx/Jn
LAp10F5ZkzoLdYnlVhtYjnn9Sl7RHVQHSXMJiGnSf1N4A7aKWKIT4LJSQQTM
E0p0xJA6NU2aUb0fytGgFGTj/v10UKWTk2MeeAKrqqYQk9GE+kV6BcQC4EjR
c6W5h1VoPsMmMfZ7JHiIVnhel4FFcQdpcueddk2Kic4W75/q72aYHG8+M3fg
GNfTKnR5FaKtLLGj69xo9teEgqXcTHxKMo6JF+LvJfau3amt9znuJd5AViCv
xLorNoOb0Q4nbKVBZ/k0k9ZIQj+utisQQh9nskmH5yXC7LJrW8gYCaEjSoC4
iEkMyx6c5K5TWDyCXQMQvSS6FxG7fXtjJIqlVoUKlq5I5zsIRAwjlQbRqkLH
M4z6r2tJSZHSlktH7rAzannM4ySDPIjuV9XyP4XIIWb/OP5bldM0guJJBkTC
3u0CbwELCWGBxS2ZkbvGR53YtYoAZFTBw8+EH8Y8BitoJ6I4qYRLHSmbceTA
1T0XAu+l78EJiuS/sZHfvHYE0T7fh9SB6qMHGNGrgMSvCYDOuP6hKTdNs83K
3fETIa5cyVSjGl3YK6dqD9ToHUdSIBtXrwm3sXqQyI/7mL8uett/xxzQz3ZT
jixEzHNQrmgYLeRAJt5PPhQtzH3+CUhAjEhSqdApqN3EIEE5+MUv7eLHRvNY
3U0m7RIysd2XQNqQwDVw0Wz4nmm3TdKcwwIdHTw4+KTkVyrUVZbOWgzBZpgs
jx1/CWKcZ1+cC2ghRJ+AWnRUNzpd0aDF3D4AyB+g5LbQjyyXamgz4ltnvIze
ZYDHrI1YQCtQevrQx7JnrdTKyqIQB/8vRsUYCm7E8amGRNpbmZ9I04JvHU1C
r6ecGluVSQyQeyG62sADzY1kFkCYQPlOlf+FOeY5JdpbBdaoEW36AM9shPbM
XmqTpDSQsKe+XTBvKhEeBXwA5ShxGqsZbkFJwuf5BbKQrtmFGNyNwIBGx61v
9vw/SqfGRAVOzShjiss4Pd+hVFPxyUuw+/CC9w1RkFRgbGL4BVRLGCr2Prsk
p8TFoDg+TvC2x/iUsxCrTPWeghLyNILLtwsYKXG9xZ3dflw2NQP3uVd3eg8L
AgXabFUFc/yr6fzTrNJ+zCVLBB5RbCG4W4LUrfgbw2mXDn1is0wiCCpQX9qO
Jq8xj2+kCbgLyJDbwvCtnuwqwSPWDKs+1psihIRaL8xDLg20Y6665mJrH5Wf
S4EFVHsD+xEFXA2lHKndb4NX1RO+d6h6l82pHvsip4PCTppjtCBWycKfB9bC
mJEuOXmcU0inCvj8iEe8UAT5uJOHCJb8olJgZg0ekwV7jaz/FnzaLKwS6v2U
ZCPqjNCsnajakqjJeirmmBPmMRwMNcbsOzk4AoM5lyzDlRHOD894bV6p7gXl
7iqn9niO4a4MBFehaqZv36ORquWWwmtqv+LA2i8rML5bgBWjE8/c6cBCPBaS
ZNyNN8jMFA9N2gtNKaOwxR1/bX5360jCWV3StjwWNOGX9ZmUGz8On1jLLIpd
Jn3SlN23TXPWrfSds1XifGSTOkaqLQFhw75scGXBB5wo5/+VbI7taqREZU8Q
jL0iHisu7BqddX2nWwewxcpVq1cIl5jJS88AP7ugZvmQwvu7HeGaeKHjS/D2
1EGEEmiME+E9uYA/1vDWe1D+8UP+fgTMPB+PBlo8hA1IsMyFPNMbNiMm545r
9DpMLK6znAyFXtNouhHdpdGJEzVkYbZW63zkSjkmv4CfzDGMGKTourLINebQ
0qFeE3jjyvceXWGD/zbHd0wafn8AJXv+cZ6jmoA6xpeyQGAWf/mbwOJmiK7r
hLCwX+auouupZqph3vPujTVUA3RUfxB0E0ELcJ6APfs8151m7U8ZkPDJIrf+
9aIrF1ZjpAgcernmjNzeFGTHZjtInOqfILAKfX1R1zBRnhv1lE9PrvumO7yH
7Mp+NlPLDUOHMx0m6LrpYPNLOqgy+nLptNafyUQNz8BmhrGSCGkOux8RcvOu
hBiGzFPEBKixiO2pxJwI1CnLYP2agcY+6/VTKs61QhBKeS46rQiTxI9+wA4q
gO4HzsyBm32PWnY9oN2qL4j3M0GDN/xmE6QATGwBmNw0sKPTf4BO+KMa9ntq
4wvfAMUAa+Q6LIhD9GCmmj2Olpjczg+CLxho3OZGdvQvVEDkKaXzzltTopwv
cY8GwNowi6ARbTtb9tJCSnz4LjJukqCg1A1tN/AcGqb7xqhR1ziXr7Bq71rq
fvDIBF0h3KFEPU0Jxct2/8FsvaHCSAKFINzvT/e3H8/jYueF5zDmSyeilLDg
j8wFDb6Ew1JxQGRsa8/kRx5+ZLzkZ2EAcWTYbWd9wHfVCP1XXsps/lCuDrZD
/NHRPPOuSuYIY9+VtONTFN8ynpkAvY4ZkCQAKZWstg1w+rdpjS4EtEHv70TI
PE/9FyCrhAabKJ3AcxUXfECgp5svoBo9j06KzZLbFzluHCvnYnriaLEw0XPP
aCj0VAU6N3G1YYjrrAwFpf6fxbtBLPwqqkPIpxu15Rr6gnNDZzjUP02vzcAN
WTK/AoypeAnM+ZIy1HP31Imak6YilL+vFTylcp67a2Iqr3Lq5x9VzX9GW3hE
6v0+ohc25VQvnEJQkonTDufcd3LNBSiqyJf1773pP6SeISEdgWs9jpl3lbOG
QRmIHUEokSv91S8I1VQvDHqAg+S4LtyCiRgm+8qZIb6rLymsTHOuJLytIkYz
bA9HCGENWffTydQqGyEcB5hJklfjQ4kWQaWq01GCHvV6pufUH+Z5aemH54IU
iJRrE3rWM4e0NB2ZFjgClmc5tFhVcVibSNK3yIeov1MjeSi6LMhLjt387Pb1
rEZFQY7e/6ybiGbQzMBbO7yob5BAyNin4XxUnt/IiEdvnPd0MRo5ed9hQw+X
MXWG9okJq2RhS4J2iOLnEnvk6E2oswg+odPUu4nUbg0i/qlrehvSYv0p90+K
m+pe9JGIKOBtGMfkXuEf69MnfFbC9wsdx/BBXgf+5F42bVO7IlcFPHv3DNbr
XUgnJ3ARfIHG+A93YWZG+EWoVdbvXaMb0/M5o1a0NJ4E06lvOwYPRZDLlrRb
xYhLY3NyuXvYieFrcwcTO2zqiJZir0u0CFjw9KLJQZ+GREdO/4igmN3ZK9pL
7+AyE7gxsK9px5nf7uMIBGwYclUH5kOAGNT/CoDeAD0U0i2NQXbx7gZWkUHk
4z8bQtvntZ3ZgyuvVCk9LIzxiYR+WB284V4BjVnQKQmgdq3ZbLhpaq/XzK4J
sPTX0LtCG/d7/9XLcP9vvtQIE2jiN9CMbNZ9F3BvzgpQ2lMMu0OvMEy1JyHO
Cx58EmQee1/EqJAlndT0GMV05rtxwwfZ10c0pRRoKeUPOecWGgGSnsj0osIE
vqKBzIdPPkpnZRHrg2yvFdzXRxrwZw8iwTXKlNkIy1DY9Hk6GMDL+L8tFuZC
Bjeel9blw6dVoJCDKxWbNBdqrLZPhSEDuM0nAlPSEiSJdN8XrN8v8sklXbPC
jD+6Fy0XC/CNACg81YW8DbJZjw31wrRp6YrkoxhM3aCM2glqHWsOyDCEEVwB
xol60rnb2EbtqaQYDUIlwdpV3wLn0awkniJr4Hg9h07WT7n/KNQZ7+7JcNz3
Rq7haK5biMjWodp9PWBLnEp21zTP7+NgIxjeI9SjxyEZFFUGCu27ekAsnAvr
A0WYJI9zu+LjvaXMUp7dXNPGv6kqXB9aHWqZDlkMSYcheBEm5oVZWU8yJ1uW
abwNRqLIcju2MG12b+T/pZBA2uiS/emPlRvDd3Q2uPGdT3nKshxjnjt4qwVx
QY9ylBUWkKsTNNsTdv/GxOvkti9nmLGmJ6CDkGSrQUvnctaoDkhX3Jzi9TYO
9DLPLJr4dYIhYnAxdU9G7O7mk0JPNMh4z/4Rccb2edtnLI3DWoXG1Ab7w6wX
ZcSFsVbFi08zBPC3XjPolYl3s+7zN8yCUF0SoBLA3JS8STmtDfdwxY6gqCGI
mISzhgJYdWdHiRagbWlfVj6SGVVXzpQ48tBLINcSNtsAGKiLWedtzHpiTClZ
lJoGHMEIOXH0ZhP0Nmh4QI4d5dmLAaFSCJTWzOvHtWaoZS4JAMUuFE0tVHlK
oALl632DogOZqSQ7io3rbap9m2LS6Yj28NWQJqe8P9SwZfxjbBKZ/Os7fB3b
J+09Qoi4DhLpqaV7M/W6VW1iXoTj9jLZtaKOSOh2VPgfOcg5Z68EIPc2dDaQ
35uLPNR+2hRLIGVGla0LnNkaQjfpbrLDKnDNJgHHyNVaC8inFo5V3qaxLOiE
Iyg3gwChQtcc2GbU26zNOjm5H7W5gE/yY2FPHEnOdGQRpRItnDyNc9YdzqMl
ZppOFunbEM44BbAydejUa+2Ktgs5RZg0/BfyT2nZJcorKdVDoj9EDGlbxDpE
N6fAygLMnCofr0hdmQHk2u1+Zpj52IXOqiHGmg32Z7Aj39mbvSO9soplsn4t
m1j5oyUZZzhzeWO26TGGIDVSYMbWRGo0xBZTnxelfbeBrTnAIljcIz/N0pLy
o0xN6nNsKPAUbwfSLc41tBDbYwyULzBQNbh/3ZJedRuJDrlqlkc5se8t0/XE
Z3zOuVAegfKpdEkgiX0D4Dkmj6wohKaXqu6MRKCvzZWVL11AjQFN7qELU8A5
VsmiMsq7TBL+IBNYm1zQY2h1CpE6f1uosElcbQ6TYu/Z21oUZLEpZmLaNs9P
eazkm6s0f3n29XTzKYBZM7oQBQkqmjWYenw8zPnfBiqrM1bkzDX2QToUNCWo
ZiO+oDRqH/LqUrCkFnITUauzmsoXoF+Qrv14mObPnECUys5PBErRektyOgSa
1SMEvi/5L82tPSuAZiKeGRXEU3qhfm42qX8h+UCpwb7bL9juedout5qLFotX
/4+bs41zrCUe82VsoOC83nkhFRDrJkk8DfUu9sNeTlgdKgj2FLLRS/oTFnD4
pz0sJVD8IZMHcfJL67DosyMFfH6Vc1dqNHvXxRFwcAlCCfIt9pFgsuvfUUf5
O/xZ/HubKawEB6dVBrSKm8Vua1+dtEn91e1B7Opx2S3C3LbBdk0qePzaIHUP
qbC1rrvd7AfMd2UGaxCgBqFoJJUVwzy5jsli2tcUkaxkujAB8c6q9yUTXjfc
906edb7oe7a0wxb0zRs8+a4z7yLo1rWSEcI3D11aCvNlpGNp53OIsXKvyiYl
9xBxmU+Mal4jzY515se1UshutMv6Nr7o4ZlZS7341xQ1GLBCDQWdY1Yo/6eJ
22y3MUVaDz/fQwns+6WtPa5cl1zGS8xvj0RVnDjCTa5nBoVoCs6b4zmchzS4
7y0zHxqzncGKI6h/FMVDLmuv/+835NQ1uw9RujUdMKkHfl/OocN2A8WjBQEX
7RsOHpzuhhfgRbY/qPaj4YHLDjdNigYNSkDNXWFo1AnPjC02oRzqKSgB+oAp
QKz7ZFhOCzO0hoGon9N3AHnyY0X/n91iE55k9eu1EQnF7T3yxrHqwvqu7/Re
9q80P4Q6yW3EUJY5kQpybpJzFo2zl/aAo8SPfMcNaqrllD50epG/cKEucDG7
atAjLtsI8mYo5Rn1QRBVxMC8ZQC4knUGxUAR1wQoxv1FCznzYyzw2bta/nRg
NY1h6lCW4zmnN5kD9tlorePzAq/JbGdfGaqDKmXaaSykAURvwyu3ZYREXrdn
10Wo1qf7jpPlAfJsIefnfqZW/eZ+pM2o8AMVwlPcu8XZD8uG6sBkBnggGuMR
tWRLfVWvDrAu1TpD0r8hL59x3iE3R9yRJW4wHWw3xzAjxfARaGhnXl3XoYH/
mjqQMVz4UBCuOKvRUbuQwSwNKJCIEKpKrH6vfpxwtgHT4wsTNKMkP0H5qc/z
7aqAui60Sey3D7C3u9U0yXx/codz9Fs6B5sN7ayxhR86GixXMBw3X5XJmZsF
948DQ8wrEhPH9xr8MoUZ26x+HHlmRFGQ5Ma+xpu9FAr10gMOKYcGs+zWdssC
seZhCE3b/OVN9wMHNMbmtpKoEMizM/H6zn5hCF2CS0k7ozEU1UsBCfIppZyn
bLvkaifilpPcithtaO6AbmPucvhokKZkfY5Eh3/Uj1/Fn5knf4+RHK/1eog5
4czbIXj2hi2fNt44ooNV3Q/zZvMOVnDbnI1y915Q5nU8/DdrQKa0/TewN6Id
PpZ5fOgXGzqmje9j4ZlLBshW0nQsIlR0xogUSTspFP3XU0728EIqIZzn+ma+
9s5nVTLQZx4ORoaAQvWVLVNsN+9OIUKSqNgm0LQEGcJVYzmtgE2CS8P5ycne
zRjFFJhHKY0lrNAR2WyCtrVseCPwwYVZIMjntE42LYM/09M0lbVzFZiF2s47
NEz2QVNEva/m6lla0GYG7fOTjQPhe4hh8DnaXblJ4Vd7tOzRaZ7dxkbm3P85
P+rJBMwIQXb9imtWBCPvf5D8ds3+0tBv4OdMfo6wRKIrjP6LB8AG8ns1RnPh
22G1gfTCGxqwATdJaWgW/kOpfoszj/rNTVKka1Fh4n2V17+jz51Zyb5plK9Z
FZsAoWXo5jfzTdsUTGN96H+sZqAxNVBcV26n0ZWEEVHGI3YPvnbEyUGXKAzq
Erto9GGkgvaKOu09a52zb4nUXu9QdT4dwT/cw3e+IIpLacqszp/4YWJYR4aB
QtMPgnCK4AsMGavdEolUZ+QxUAxaumsQrOr7eB1df4zrqkZMPU8t+RDgEHFx
KxrVTjV+qg1DwbkTLdOie3kada4i1A0CFSZ5XaiJCGnYWSnLg4tnz9FHUb/O
bKq3MO1Q8eN0bib20fPhxrYdd7XFO+Tz39wdJb0NmDMLmotBe9BUDOH7335n
dfR6eo0YZeD3q7ALOVikwAWvx77L5czxNDZgdOlB4BLasZ4c2mc0uhSmXR+i
Affnb2AJArT0hhibaRh13/jY6iZkpm4Soni3V2jjtEetX4iEz+ia8Sd+kF87
1uDwMSrbxbi+6YpLgkIXbuFBw9SbCP3RmaMcgQEQdehrUHfkU/e4glognDRD
jsICXH3JNrh7Yrb2AdHG95PR3b3a64yvNRsff6le/e2UbM0/07cCCYUs7Dbf
3W5CCFAo9Z15GhxR1tOhd1ftZ8mwOiCdnl3LGWj3SxftAONDOoXn6er8drGR
GGY/BCNQ7LrJ96SlF/nXlSetdgK17U5ah2Dadb5YeyPX0CYpCtjf+dMi0KV3
ricKFOZAE1PpLjCm454D9/YmB4I4Xn+oq7GXjk0g1aw7QiQ6tkDmkZwPwNCu
Y7riH5N9x+qgEOUuz6e6rVXaWt9U98zyvze7diBUeDdO2VMgWdHjDpxmtopl
uXHn7ayl3vu0zNAoC/pcysVe0x+/DN55H1C11LAzf1wxGVhGu7P2LrYmsxCY
UrlO9MWhu3UN39hDKUKAm1qFxm1czeSqDSv2dxcJTn/tAseCL5ZUSTu+BhmR
mPrR1kfO2oxF/s8MHXakDUaU5FDc2CA4LGwOiBh5km6hiXIMLUpLyF/jnHw5
JM+xZRb097Gzs/TmRg+4b4rktd+IEdI6F9JyjoXc1GJDxuXMbS8R0oc048Fy
nP4+lZ5hIwohdGrIl8vts3v6lAUP+g49UT7z6aMe4yFNoAZBoPlzKxokkcjn
KSQMxsnQSOx5bdkhDUFA67OBX+/gUIJCd+pri3L/+sboYByGH3WkxeLEaJu6
xnTl7nDlE58bx/iHGxEQwOa/KhudnTm7LHpAM5itlV8v8XyE+ydi5uSSmbes
mNxggiRY3eO9nvgj66eb1Dm7wbbwHpi77UbT0IPgaF7PDUAYk0OTtcoxlkB7
7U3yxCsnEFMS05Tqb9lM1Bz4bMRk717D27iFOOCiQ6Cci431DMUk0U1QvbDn
ALOuSn8OLY/Yg0YmB8pE5tJf2LluPh08Fg2RwoAiJiv35tG9eA580huR7SeI
r8lVnGnRcbarqlvNAWnUTHABAWmDdhHvDrbFWTeKorrcc2UN0Iltv+rpBicM
OSWcww8Y7dsESN6kNMHVyxxPcibt97n4CxR2CseBx1pBPZC0qhtxiSlQHzGk
5pTvhEsSAJ0mokbI8dFBr6DZaeQHoIv0xWTvHkynD3AMJG/y8c+TAqsTctuW
bSVnTJ1ISIM6dntQrs+P4q1+tBrEr5JnZZ/lHwHAZhYu3K3Ad8myFy80nXIm
YGOjzR3Jd/oni/jv6zX8M5J2Hl+6X3OOjEC0ZnSdTyh0SwiHAeHC7C3sJFc6
Ig95HISRoX9INd65oBu9WelFgWmypT24yYvW7muKY3XsHeRPcxxI2st6yFpP
CXGDqIEVHpYUPt7r2gLiy8kv5lFR3Ig654lzIAv0pLngId+3/QV8mvj34QPj
oRcszUYYQ65+J9zYX5cqFFLgfrEwLU022wliQLAk91XYI0CdCsi5k8zBaVXE
iA+pCsatUvb7DoC16hl4HrgqlI4pVBmoHsqhwjkAJ9FHQkPnQ/Uzo8x6dxZL
e30rT0YmAG4XZLT3fLLEpAcnw8VR5uynRMxzvIoSfyrB2Q3IS42dm/vv/cZt
jIBqZeXFJQlT8fodWiCgT7B9aY/rK448gXXPm/aYQ+6dqAVou1a0t8JyzSot
7Skt50OwJ9J7l8aGTfa8mnnKhuwczJlOc1F9ZWem7/wUJJ6eZCh5uQiEfDvw
mD5HjKd/St58p48aAdbn7iRJtDOWX9kq4ji/u+//B+8iXtBNwl3HZmMnxKsC
RZNAFdt/nU8N8cdc32/hmjrgad8+uFgXE7cHKpj4Uh7Mfn0/KxKC4FDMDLep
R2WAkIfN7kD0PbY5HDUMSoNUPwzEZpUqearVpnILet4S6udz+csXsBqJn4un
+jw3IbYlUZO3jO8Fjd1dOSz3By7BTS9U4ldNCuvn9KyaQAjJTR8zJzc4rikF
XqZAIo/vs47xGilqgxLeWGppcz71XT+wJfsHTDFikwksNG+kOvYSg3VldYAZ
9Ip+T6Uo8IzcuRLkcTtuAgGGJ3efovUFFM+//OhtA9FxIWhFfVVdmvDQL3H7
lcKIbRGxJUdn7az+QY0Cx8xSJBmLg15/AppaabhmRvSgGdRysaXrRzs4ux7y
6fY2imf4OuM5+vPGtJ8ApqxFviGi+GnBYr/UDW07SDO6Ob8n1165NmxdF0pv
wWkrj+SBGz6c0dM1HUp7X7YdZLrpvNt4z8Pk9Io2iviVvxVncpx58dftN/z+
+a3LQ+k0whljNEVaGXsjLcAEwDGKRXuDB+OA8V3lYXO0eNq1gxkzEKK0Fi59
YAg6xeAA4aQxl8CXNgM0uq8NQgmdg5FNEa7ibbsrbZD95SVY4azdwOz4E2PG
K7xSrTVUoDcXN3r5q2AygowQoCd5XJROFiVKx0WQS8dYbgzYYcJYypkLh8h4
uslY8wCO/kR9Lhut0yWAYC4tgEeCvXTbVrgdACJTEoNcgRUf4aFzdhLfa8PM
itBdf94YBK0cCCmlbGmgQRDgnWbgekZUf0JuvGdB1MjgMGlDxg0lmK775MAK
oPkKsMFDSds35sbjgM2wWBcJSI3SPPl3JHYtQWfcyY+eLNNfMyK6LlUszYWd
OwKJoGXlDOJuN7Z8176y9M9O+A2AxsofEH6zu4WF67iMjzBrjnFkz6/N1QFC
Hen8+ticGvY+J7x5asoo7jBvTF+7GD+kuWBs1wKZOsp/IAec1fe14g/qKXvy
HKrxSsqKCY34P8rsJ17cv0jRTtgFnOm0qdKImc7sWrSRAfiNX6QuHAEedwIo
pSafSp/rxSVotdX01SZmjXPHy/HNbXUUHoBPR2DS8ScnvoOKp3Uf36GXclrr
9UnxgbXwNXz576QdPj2ckvcF/3Lxapd5KSG/qrnl6gN4eZ1XngwQ9Grfz4jk
6QvfHQGfU6Uk/djFQzypwN8pwSHjSrkcWbsFQrfoGmWB5eKAa1Ox1Y7PVZv6
GP1bcXHDwwkvGajVP27P1uCqqV/hwyrH4myXD4MLcuJ7ewqUzMPQp/NEburl
l/2JfTHBeQ/jUSPnrOsQ+FFs9dhZcaOM2YGiydk8qPCnXr45X2BT5fbuTO9e
YzhmwC6PAHVUPDQ1GjlRlFPRJcTYZbBHLAe01TAefhqSPmXclumqa+p1VqEJ
eBWPwTHMc//p+qnTt6udYDn249KljZ8nANC4w9z4097mqUjbE9Ggja4AjEeZ
0J/4Jq3z9yiPFOaN3/SljE+NUH9hQKR/OrtVl5NnG7L3uYdene06CNCnBtX4
96qLLh3iXWFClwaW7UFrMACTrk5BX8qQRRuRf+ngPNOl6pNgwu/tjy/mFkYK
eop+gfG8XgNxoe9w1di2qIPpgRxlHQsED6r8KcCVZS0ysWTshi4ag7hzP5Et
Y41Dji2bQsnj0XXUA7OES3hSmr/4EPZdTB9y3wYlW2lu4N0Hsb/BdMxugluT
CMnXbarGZpeIxGCLYEcz246RQsx103lU0jHn8eXnAJLqPgKhtSQei8qYVlEH
jyjOxvkfuZNuEhMQsp4ziPP8p79saYp250BEmNlqvWY4nw+Z9SOuJFRMApnj
oTWNg4AEWpXsLZ+NNVaycrca50tAiJ6tXAV73dX9sDW1C+ble8o47YXmQEr6
/N70MWKKgVvEYeOIyqknAkKGdI4UcpyVn9F4OAp6ChmdA4n1losVhiEDtXDi
PuY1+at0vIm1EAz5cSJWPQ8Z+CVzpXQ/nxR6AiFTnNmGPg4cH3IZtfou/aEv
Dp8SxnbVP7N3edtC67C90sRb9TKyTc5wefJ86quTJibxO8SFnHhDLaDMb52x
B3aCaYjAtIJDg0OaIeNTuer0w85VBbCiKm1yiUifaxCfAb6ELu06U9IZ6OUD
ww6zaLhkEJR5xLlY9sDFMzAR5wHAHSF+WKCZRbk5Kapvx/Ts3BuxF6032Geo
1kAkABgs3AU3jKmPwF5flSi0+56iNTH0Iv6FffooCBlvQoHkUPaDWJJ2Lr+H
1Q46XIL5HzhRXvOOfAS0xbkTVmoN8yiaUi2tRUBcE41aJTVsLb2TFfUxC48I
gHNEHKuU8XTVFPcseIymCiA5mkUXlAyGVK54nm3h34FGgolyzWHndFuP/Qxg
kZc3yOIyTeJeoqox4Jx12VhXG/UVkdXgRKr55YAz8TA47Da5Qp/nsn6QI7gP
dgdhA+v89hGG7a0zrqQqpogoWnTAPRv7jcjo3lfSUtamypWqTD8D8BI035j5
+uaXUE9eoH+7tfk0XeNWIF8splOLLV1bBFRYn0JnH9qZws4ijqtERAupoaoY
EMh8VG1JLzfbbbaoUqS3NCJeSwVedRPGp2lZQ4282G1zY5FU3HT9G/9o77C0
wVAzrqPmAgxzhIn9oJ679hKtGeZlwi/w8ICyJpwbNrd47vcoM8fNH4wtxvSg
fiUbwvzmBwfiiKvKT0fSOwC3dyLNZod0UIvVT13oyGQN0OWJchsjGrBlh7r3
7gF8J/Sv3j8mkJTSUuKVcWLqS9o0wb0WuIvziWp4yrwGvGQQq3Um/HJ5jrN9
9pOxlRHpit5BPuvWAEwKJJ0xI8D6BhZXjG1u/3j4w3EO5tdfDSevkJaVhund
nRj8443EMRCCfWOtP8NZoqpT4Al8l6FOzvnZkMWVTesXHivWTlgvPNpuaM8V
i7vnrWOfrX3tGV6HMAi0qpHfguPtoIJDt0D/iWG+vsVP9C8r7NWOUu/lrDKk
SqyAcmdPIwqjmdFyyiTIGTS2HDH84+mVfn+zZJ5524FFRgKYcSU6iLJwKx56
xCWYFQULu5Fzo0IQFu31LPmtxXwkbGxomQndMxL4Mi95tLD2P0Jwra9PSIQu
4FX6h94h4GpqytToDngYiFz+JFK7Zf2I9G+Zc4avvEWaXAEl2jVc6JFbNBGE
SD9658OfyiDvloaNY60NnlQH7Y/CqMPVAKPhbaoUL9L983bNfD4RDb/CzP77
0/YdMX9+/IT8gLS+Lztd2l2cCkLaZpYA0Q5fAgNdIXQuOHQ4GiY6pYTFAd6Q
2lUpejuZvREagqVJHAUKcHpZzV6N9wanCmUMZNMtUaPo+Nt8UhwqzBGabNgs
EtXrYkIoq9zBIcgWCQfxyn8qmb3uTRI4YwvEFX+m+pSpnjkm9w/NyLdGLshW
dswNngI/cLUB7MkbP+6BTS1M/wzRabB+TXD5nH2sbC/k0xULomN1ilTr8vBp
O8OLl8tB3BDzuT0kdTFJjlXw7dX7wCnBSKuCgPNNSDi4eNblZo2PK/CS2bw0
/WifU6YSrgxXOyF/8P2kWQTLCIeu9/JMpfJSc/kIuXbJZ2r3OvYATpujOssy
hB6IDK5lI+GrHmEswjXnWP7hPeKHXeDA+zfTivolPYDgDprb2ME1I6eYT8pI
jw7lRVHWq/xQwjfE3+anPgKPZ/j1+9atUsuVbHegh30jddoTKakLx5lOlWoj
U5WjdSGtL3YnF3NrxEyNHTP+fHfOXNG6y7BIfemniJ3CQM2x57QbUp60+jmu
7uTUJid8zCcbvxXDTMu8ID4bleMEPFKfArZHRBRSe9d9poXj8I9WEd8u0XC5
c8KVLb9mnjlVtNOzgwHaM43i0BxvfBPLqaM7ei3atBREZHch5BERB++QiPpH
5s4x3QQRVWsc7bRhSsr41zEs/+uQeLTyUYN/hnf8XxwoW7gYkbms7ygs9u2r
eQLyHU7fiV7wF3vNNxtAH2xWKKcz0E8hWkiVKeXFBtjLggndhM/Xh9XlZM5z
oWhz28R1vmzLiYVs8tYLHXYC1HGRcdLw67KBadIk8xciTPMA03cshyhlAApG
0DTAA32lJOSePBk+/CkV8IWPC9qVoiZ2FfFUkO4LjcSHr0gA8snQX/X01Ht6
0C8w1YeqajdnwUBeGuiLi7mkwOSf6Vzl2lzAitC4AJ2qr9k6vIH3LoWn1apk
9qg4H8rz01cUVfTrwt6J0T428Y75tbIlCutT2N9+hRxoheOVzLSbeKRp9Ckh
PgXDJ4DsZcuEho/O/+h/oj6zKyxqIdJsMvotWS5+C6SprcRVgr2dhtFCIyh7
+hieOqgtBUEiwA51u0wW8IJN72n4hZwUzHnqX7zoEJJuRjBTCH/mII1H0TOT
frq/RD7BKbzWrbAgzbEd8NakqJwsmzpIUvHwsZ28HXZkiKPzOhjkEKVNub2H
mMj8dNECYrvBHcLyfJZA1sr0OX1ZMR2ywe/0eOwGp0cwaoStvFtlBOjWqCEW
QdsQF5q38GRVqkAtEqDZvyOf4fzc5628gZMt6L03Eb4QogBv3PFtQkDElIZ7
nA2o0SLfWJHlnfZt2g6CmsGBEoqpAH6ejN7szJXLvuEhzIF3mBDG971FcOFS
00KHyaW7dSjSADttXmrdYMX4o6pKUzYU6pQp0YDVqv5sGSF8jKOCAEm0jTPa
0IDrPGkXcIrUWe3zMvQ1YfvOBINKH2sQKX3FKb63V8buqrxvORDbIjxlZk46
nsKuvx6Lj68N8CIoXioQVDuE6eAydTtPcOAlYUCGn6cmwf0T8sHsJRTTLSTG
Q0xt1K5pAo222fSDki/MFIeuMrm33XPODhQHERIYLDowXAjHUqGvj+CBrqw0
rxm2fFSrCzo5xowGx1jMrT49Dnp0ipP2+RIpnlkjsgi3OyqAXM6m1+VFMx0W
sw5wnHxPIJA8GpOoT4qQNwj6V7XRUXIQir1MHd6Cvsb8Ie9THa5SoSXcmyPH
KKHeB/WG1d7GdsFoyjlMpEjEd4hh/sd8nrxgYOlhXZqO1LbsylIGiZIWBE3l
otkTN6EkPoFhkVZVBt13i3XRObpjrXceIY3A2fNAS/7YVhKEKsA2wia2HOSR
0rDyKtNyzLsC6WHnZfSdCXftwjjbQwHdeg99cm6df59oxoNxYdk+SkMHSG1+
hoSpESMnC+4SZMgCrtpfKmrRc4NKvEi9pyBw8zUrKECRkRiwWwXIAVtou1WG
YBXDxgILhNlwdGGyBZgALGS10G/lgJAQ3yplJuoWnJR9TNUgQExOLfOPUs8g
iBPKHJGUTDIMYv+ax6sZuJBnsWyjS0ZbDI12CZGqFrk+R9ifjQ4cHaiOfObU
ARi7AWRP5QVfT3JMuSZwX8WQ7S0T1V3ivzjn2JajG/ZhcysNZxFvBVUJ9Uiw
8amRXpKRjcoZjFFv7Qg52U4gmUVWWKtqWCle8u4GUyplRj1ri+tvNU7e2esW
waC3+eKSkIHbCEiLKJJNPJ+WwwlpJ1B9KLSVENlZFzaixGe9+UvXp2QB78W5
PSvt9Knww8eEqKabNWBIvzNSmJgdmMsQ3vE0lKGRKw0FhoF5MyoXpIAf7xgs
Xok1xQ0Ns+hgCt2dGoudsj7q1v1pVJAJL0KhRGXrwjhLUPZm0TClUJVDwDvn
zXEV/YShlEJkcEr78XXVHqIMKrLgWgFV8202t9JPOlmGSVdt0Ltfvbm+4hJ6
0Kd6WqnvAScTRnvLoLzefgrdfqkV6WXtwFMQR2H6PJMcKsh5vEVZVuRAejED
per3MLxMZ7BsRt1hENCSRKJ6eI1Q/9gxQwfvzAbA6T1wS0VLG58zVHKlas05
0iM/s/9L6QDNagS0cXM4FUJpZs9/Bmp8y7AA9zMiPbNTbmjReP3qFTbYcaw8
FS8bfy5kg9SaVZqLpudEQr5rTcjWoV/hvpbqUjHnBjGU+ZAJAYiO6LNLmgTx
nFdfhmWZtmpt6HOoI7N4RyRsS5wo44A+aoKh0KFmETPYX8Hc+YlZv8sGy//G
B8VTsP1P7oF6n7Rmfy9EVYq/cpPOOPyadvL4m8uIkb2B8qynsO7gYx3DpXPJ
bMQ5de5U+U1s21wa7SDcWee5UAhfrnclh4yFsuM3iueD7I74G0+aJyeli2kZ
ML8/cGLByj4nMcxdzAoUEnzJh0jz0bfXfTmH8u0m3GkBAVytJhE4Jojju4z0
kuPBu2D8/0qq4vqENS66aU1MwleIS/mkmi4TZbOpCE/yFp3GwDrmk2YCgwP6
MQwMj0LpkoKoU4pay1jC4vnbrR8QJQbOl5Vq8GxiThG5TC/23l+gu3PlEW28
+tcPJvkeNBbSpn2Kco9apdK5TgA3enpti6+brI1gfehpGCd/1SGa6SUrE1eT
JQqYloS17TkKmOHk/KDY0v5w8ae/bMCKKUYIzD0k9qn7zJ6BHRCuiVBsvSda
5a5iIfYRTPbDFM4hJJUDeib214yyr0tnazxP23jqcuGDQzjSwjO+ERQeRcMz
7o17fMrDzmMTnDloMZKViJxST993Ba5P+FcQ99eo7+kQ90kRg/M5KUiXAeS7
W8h3Vc36CR2mm6Ch3pXC1XC4gFaBxMK8/3v+L58qp3adRZJDXBrsjI1P01MI
99AnhE0K3wtP4h6cNyePlJOzm37NqOaQodoMeCJ0LTzOCW/pTpqY/gi4NaJ9
TLgoIeqBjgERT6d6dS7eWhsv2OMJ2W22SzTi4E2Pv8tyKwyG27H8tsPKwvZJ
El8+GpJ1eZdYwLO8Gdj/MPBYu+XeEcV/jb1nMJuY3HNvlScoSTcByvuJFgCA
1BTA3RgZepHpTOCxtaqLqGT/h1KUxyF+FbMDUpUh4hrE3lA9Cps1ve0K8R0L
icFTlh+VSGPmH/frCqh3zDJbMXdV4kjsKPhB2a8iqJOetsGtiy4Jks1XmYUS
+1qIxLoF5Sfpi6mYUmNJjXE/ohuHcTrM+fpTzQf/oFt1vsHw9p7IXSMDBaIG
naiRcqO3gVcg7iCwKcAUh5acox5zYs4vetR9hWWdAQ8Sv3u1qVewPBjXfhWd
fBB6cVPKmgQPlS0e2LMxYJ15iLC4UpL4IlfOXJKpDGv/dZaqAZg2zdoJZWhe
Xgi6MiapqiOZM0v1/NKgaIx8kI09HQRikZOfdKH17EOaQ9tM6fZyiL9jo36L
b1Mj1Wf9OA/54dIa9CLO7NIU2YhjB5+CI1xET/7ofOyjPBVhxFUOIR18dQiI
KSvjr2M4mSD4nNgMowISBQsnvpMywNR0HxRKsIcFfZQUeOuMWwXzmkqFWSD6
8AQ0Tp560s2xhlfZ8jKDXAJ6Hh9+rmbTuNdf6bgId0/YAs1e2/Yh/EB2KqwE
mSb6oRlIrH0HQjeymQpQkzsAPYpmLsQ0xcY/FBDjoY9ZwdiIF2A1M2x1o5SN
in63FvzLERFXy6bP1KhS4mUBVLz6YpopjgOh4PoMP7lIpDJZ5uIGVB3rT+vf
AJ0LL2m497wdqZ8gtpwoePrkkcNlsW8Ya0KNcuUSNsmx4FR895isTbvBVSJV
fRynxZk726GCoCEWtIhpoTG2k4Xewqx4bM1QjQA/lsFspjGe36Owk/ojrr1O
WtXu5nn7TicLfDIBhJZENF6rBbhVNxZd6umSam/USKTW4/qOxzzpCcyKc8OV
ZAOr1EVwbq0i2rGe8EaeSskf49L3BfABtpgjdIXcLvcmDlXahVlIOvFK7hZW
ZCPqlcl9P5VN+ZjABlKuvIfjQMM2E1vrPz96kdN1EihbFhfzZGihk1mHzHCa
qs95B7m3ih4k13rRjz20rxbcBnd9KByuWcdr73uFudpkrykz9hkoNlkbxEz/
fYeb+M6Uw4cmUPRBPLPd7/Y+otCExHusoJ3dpAXURCWL+nEdtbxRoR01clR7
8ewk6Tp/Jzt0ta81M1NmuZqaxIW8pDBTdzjUGS5ODxyEe9NIgw3DLSDaIBfb
te0Ex0uTovG4J4IJMFClCy0XBLNiXtsr+RUWa+s5/b3OD07Z3IgM78brABZe
8JXhkD29QuIIyYmM9pZrw4HnrMjP6kxJbOxg6ed8JJpPK2MJ5lQE1S+Yv+Xe
5/ugaa0QJA3/lsk0ETLjIq5PfittxYAd4xSOXtj8LG/k484EzZKulzTc2drC
FzQ6hrZ/f0CWE1ghhnP2bfolrJtaUs/CIE2umyCJRnj/m1kPq0nlcCk8kqsB
EX8cD5hlOQIm59zyrEpCh+KULcXk5RKXvqRj5YzFIk96rDcfDUMkG3LnoMPm
VOCXjxiiJUQi8b/Qfpg8jHq/JzcQEOFy4mLbtae9UGmA7VPX3tF0S+WfI5r9
NZ+3qd7lGG8f4+I2Vp1KCPVoIle/m5bnSW2HRSnVZ78xIDFf24b6CpEefG9q
XFJMtsSb1xB5AfOSA6mmORCiGQX0AeyoRlFDitrj7v1o8CS6fywKX/Km7Y6R
//KcEfBiwv+EZq/iKEUkU+ssdKol+9b8MNnIJ7WsKeVUFzCgiHjGnymvPsvX
uM/BgT82DiU2kyRdw3UK+TFLn/ybpY5OWV/OFFtfCCOnPp5EzCSz14d/vWsu
vAhB7bRM5fwEXUkfo36D4PBW8wi5u8T7EUGWLsZz7Z+yZmuGFfcyxUIQucrh
9rjjwu8xabv79dZw2T1boyJNuOxTgRaKR1DXNRj4ov/+KPCDVJwMhxjMurW7
s/Dsv1yfRtz/ush7PVrzMcYS3RDiXby99ELeJjT9OoXGtV110i4VOUCAQBzy
zzaalsflZRt4yzmm9DYikR4Scj4l/ex4n8I84rf8hVTDYPrlTlJwnqX0m+i+
0vwEG8t/Q1TteJGi6wCwu9g/+8sQgDYPZooi74E77aiZNK4d2fqAtzi2GPU+
HW/CpQDgILT5fxmRfstZHoS8PTgZijxuD7CuLz3gTnfWd+NnxzTIuHXmi7FG
ZnpFGqa4P1TgGbIa3fb0Y5a4qNigkZO2sgpb1XFN3VGvL9auTIHyq0EVZBEn
ztBm86MduweQl+3MBHZEVn6Pz9gPs+HDHaMlFD4Y1E5/4kTAmYbxM8YIiZW5
CKaxdLcTpDcm3YQ8HEVIouBO4CNJTYionvPeGzCYgm2V2ihS8Bah6AZT3fS7
25NW2G3Xj8PACT/bZLXkfikV9DlEZ2D+XEhH+rgIq+u3v/5+rB+XJ4zrTxCg
1xzILSA9axTK211y1tNyIhaWuIYdz601+D8BLqK9QTwe92btbSy+vgPROUqo
KsJqifs8rnMJcQEDA4nHeaS6pwUL8axjmkgMVDq8SaaK/bPcjl8brpPBECvN
5DvrYuawml0bM9KwdH3Q1PdlFM0UbocqpH9FOOvmIVLKKGWJIoi3Onptj9ur
rBozjVFgYVHFjOAdya2/nm3ZcsZEOb1tixCSvMhN04vFoQH90L9MkcTHJCy5
oPkqAXpfhP7UnqTsLl7fixKw+YSdAup6cvhT54kiBUxTTNDxgo0NR1C6mckk
EiULmYgcE4nW3CNi9X5GjDJfAZkVBIsU/mlMZsbGwZWE5ukRFA60hs0grhha
5YRGzYNcF/+Isg2Z2qi6FKmvXBVKfMVn2Aqh0BooqDEgKApaOqronsoxiNXy
pm1CxKHuAJAEsjQlMbHLsIMT1+5jTKODCaNH7dqS/TlhxIbLGHqbLu+7dHA8
KsHh63du+tI0TbKtLGOYMwwCWbg1M1rUSbcwkNLcHu/VgsnRVEjsMWWRr3jp
F9NyQVbTnNLEfq1v9Q9lpvuhPW15QjlLUSJ27MM60r0gcs5ax27Kx+PTuNf+
KEeUtc2OEYnVAqUL9vLmMPNj4dWWt6VyOfQKqA9Fv34FxD0tA3v/qybgfp6v
KOn5AZDqvFVu8PzvXDsOOevLoCzjoSoJDOFb7uSkbmZjqL+bqrq7j1QrdMaN
kx5ziEyTQpT75NrPSZAN0JJkfvnWEwH/NZsqcMd8lpSM569Y46eFIZmOamPd
YO9TuJX3/Jpsca1Pp/aEqiV0qVUD8AKksWm4ixsMDEkudeLZUPO5lGsv9su3
pCgfzxjCYjp1bpIJfbHZHHX5aSyh2Xzt7+B6AFVuQZi58nxJbxJIOVj4lUvm
kuuCMCgQ/+BnNqHpWb1TIs5dWoKWs5DbV77prHIqPm3rtqhTGYnlvJuGa6oo
x9fvGyd4ivjqkpRw0PsXBMeDG2SP693OufGx/7UaUGO/zXzD9zjQ+0+NSt1b
bz6U80X/kcyoRWZfJ1lIhg0AqqFrxvM3xU5QoW/C8ki6d4FVxD5KTGQAtBp9
WXlU0VvTPjTufKkT0GNPyUGJoVLZ2w8mY8ypKWlvgnvAwG8FZxPpUbJjq2yZ
n5L6RqIqGnAEPUqBu6/3r40SRNXiobhCNTy4lUbPhtPh/aJnodxaXfKhw8X6
6l/bqiCgXe+mCWCH5O/AJ7UWeGPoMDKaR+lOaEIbSGkjMgc5UJdGsCCEtEja
4kalqFH6k/YOZUMpfBjeqkXj4X/Fk6KIy9FTsqHOXLcuDVjtLr/5mdDvKXjW
I9kM1pENeBfvD7fFbsMI52ZBeGP/CC/jvZl3CLhnhlxX6bEBQbTmvAcOSRit
xynLBi8bbsvWXY4BFDI+X5wAMdTNoGaDDtbJeWrvIsnnvLLT/RbrdYno3qy0
iye4ni8bsGSb3RcAFcdC6mR1JRx+HLlt79kfVIRLT95bi6JqEG+4asNQlQcc
dDreagSBipqAu+IDcdIyVTI2cLrZfISs23RUdLuRBp3gQRYvx6NWHx8IYOjn
2qCoNkD6iYRiC0eHizleYxRs984/+eDOZR0FapFVQJr4Lat2qwK2gBrqzIAM
vs78qaeV/Vh5gbQntZ+Y/rqcVB9TBdqbpWT+zgJV0hTw6rS3q2jEoj6MQ/mI
PRXENWI21l5qlWCAImC4cxtnI0JbWEG9DXrvdOCv2AyX0XiFAQ7o1UiV6Iud
+ifoM4vggJuUfJkh0XnKlZjvapjKCA3fC4+cl4cmjfwswJ8sUw981bloWphh
VCm4Z8RYyohtg7PfAnKE+wirvFzediiujwlbkGYWNFf+N0MR1f4IykTH105J
IWAF4a4jHgW2sU4a9fvTrF3vmEc7GtHL+QrLPCSEFLNk9RIWAB/RaN773iI1
CAEJ08oAyG2Vp3HZyFZ/SXWo2NuUpXwOw+ZUyAvgr3H9jHLR6D99+vTGEXDz
NeKRhWSgbjA2Dho93IzQ4NY7jxv+JdiNHh25lP1aGIk7D91XrviWJub5mJ1K
xQS/XvJkjSdjmd/mdst0gEJHyy4nHQcQNdFXWwI8w+YDmnn5SEqXatS+GlTi
vZUWbe4INnXIKq+bTzPA8jP162CdxzdtQGTZyx0teSh1nhnVe41hsQ+hGpm9
qRtu+vgo51G65ZWL6iRTPHUgzgC/I5WC4tc3ODXu9B8k3H49CHBoXO0XIzSe
mDPM40M2y/nKsAnnir10s/mDXexInlZ5PnMGQr02jYX/9Q2P5czAmyP+rpLU
Do1RYixVr1wXCrt3LLQh8xqqcoAarX8KA0hYIlea+RPKSafWMSzrJ33fGBNk
5xItvY9ElulCT6G9Lx/PBcUf9JxJoVpFEay8iQePE7sNF0PKXvbMy7PlBjrt
y3wWX/SlfH90S/5y1y3zt9aNqCBfFzWEkHL3W//4dwkJtEhvhktR3QtY1GGU
drrpNCZufyVHY0WLZYVg1uUrm+jvSPlXodwDsH5+S4/hfC7n2tODdvLBbQOi
KCTdiniNTtqAELDvmId1cdNmuRbCImmDEPoOAipYEjUBSHK/eYQ/JHjtI71E
k76p61FNvcxuLCyRjp8ZRxU/KgpyBfcwZvyPY7ba19hARfQs3KjS4V6hwo29
0162JnGlrhKd0wDfnXoyQkJEqK9qT22oknTBCEz30+bTdJWUNa8Onfh6wqWO
nojWcYBhah7vr4BKlVm0OgTqDSokskf1OlBvlX7aHwhw5RCb7UlGiFfmV15u
yZzQl7ATHEeH9YoNlXEy5IcAgqYveJBXXE55tAfkW1JJiX6+g8iktBMMJDwQ
Ijwp35NnJjHDRnL0MLOIcW5TEXl7xBUx56JpUej9Fwgbe17PtOFTgVkSiej1
5DLdveotCGETSi2D6+7JI06Juc/jjD5/9s68nDzRMTmzHF9Tx1GmgVz27xeQ
h1PPIQvI3sY9Gi2m39x50DqF3XA80zekNtOvM04k6DBfL/XEucWY2A1BYQkk
QqkXCT12LTEPV4NM99sNZrBG7Hpza4AzMf+UqaP6M1G+y+Uw1q0L6NIeD6so
nvj7H39xF7aUjZM07nsWoGFOUExUIW4uQBQTXtzqnFEIciEaNz/hj49HAOyZ
TnJR+9Itn9g1IL1fnx2gXeOpmjwN9v4x9N26S9D34ZvUVcJImGycxh1p4YuE
/Z+q10OzLE85Zt+me9ZWsXZ1OmkQj3LDsdhnbr8EcMn6d5fTbnCAB6A60pvl
jGJXvmp0v7IYwYjq6s5KgYwW3MiBbp5FaoeJs8cIw4g6cDR0352pBX1EOfoi
M6JIjb5LxMzrPH8oFjYmrXEFCxXU8dojNL6HpKWCgAf3mpGaj3Oulw0aGohQ
3OItl4WtMRfe6FKl5eXml/VzNlVCt1DLTep+GF8bM6Kw2pYeIhJ9wY9x0zw4
uSCI3YeGMcymA+75siCQMiDztOOXWKzlmlVDhseUXL6grMhTrhYYuHSOBwDF
4vz3+CwFarijS6LzxFU4Y84tiZU9gnCWp8KmAu/hqD/1OVPO6iSqoD0cbbgx
upll2zi0UCcSPtnBkazq3T0WMzI/h94Ge3nwossOnkp3a36ek6okxmQ6rTwQ
qKZS+qDRhAf2jcV1qUt57xngPZYoPSqwjj6+Ps7C3CK5GS0HShBk8kMayHtk
vtXyWEgi7oOtemwkvivuxWYPTAgewM7hlYlqHWRywEBydvseyNkmKfe5Tnh9
I01bp3pzzkhnVpYzDywMxaLypSoQwlCfkTZpL/p86OibbB8ZqO3s+xPiki3X
lbb3BGOZFs20+hXYU2a3hcb2Bc7Rn2gmLFuoKbfXVDQk4twAVe9F0y6MvbIw
pW5qrkMo1LIrKkBALUb8u62WvmKcFXpq9Kd8xvGND6ZUn9c6+pq4yFVWzZsY
FFcVydLFCUGrp0zXCTwfjhWZvpv4D+iadt+3BPingEj1DPV0w03EQ00CkmSO
R/CU/eTRXP4K1928PASYHFupkCmBRO8NDKYVtLMMVfZssIkOgTA8eviBGDrj
+wqRZI8hA3svPC0k2dUtpmzjffYTV/IouCUS+EXFWaNb6fwuAzZMcWJlXcSO
i7oviR3Bazmxc1E9WQkWoN+0G4Do9pFC8uK93nWQ3cztFOR7i2/jf7+vayaj
s1q8www/ZPMQ7dgCzQjoRGLhjdF2wlOTOmTXrf6D/IUTgrvsUHmtLtyK+Vhu
p58j1soeUpJl8eMgTYupIDSfsO3tjiZslolGaeeO0P+WA5s79vmpXUBEK/7t
JtNwb8o5DUurH0D8QAxiQL3LKPO5wyxWQbGRx/aCAGqDGPXoLKNZrSgSLFZ3
I55e6XZ3hXPMNE/mbBtp0zCETYd/t0hEuyae5aYGex6BLKRAHTJDMBicPrz7
YqpVkLl0bgoOikDF0aWasRzSgpn9igFtrhSOB1s0/rYDZwndDkcWn3+J/3Jb
fdKCrZ6A+yoP4gPWcBsenH4Yd8XwHnKsR3ToFdnM4ihtIHvGt8Nlp++kJed7
kUtn39mlZPism6sdIqB8HO/xYSdEsrzG98TfhMysJ+SuofWDVpKB9zJNWQAy
JDgrW1NBpVUhA7z7OawXh9KEnL0sN5IgS1Ff6OwX6yHkNLraGb5UcgQgYn1K
PzFTwsCNwtrKFp3MSP/py9DLZ++8E9aLKotx2gCEUSA6rw6D7rcl7/j0WeZr
oT7CUgNDwdHMUbX1ByCYNUKh7SdSOd09WSJpRN73rltfXJf3IHvEBbWLMIkg
Go2TWpnuZkmLbawEkLsFiTJZ82WS5GOzKXw3OBMDaN1ajgAdzgcS524ZH8MD
6+SOlEPbbWyURLY61uIS9660NCl5/fp5+rewoVGkBW8tPzjWf6AiI+j2kjxf
7I5VWaqivXU3xNM2jxhYPUWhLAtK6u9+6DWDrkekY0oWXm1XxbUe3GrxwwQR
SV8FYuE7ozwYc16/Bul8Pkigqkfp1s8Um8EQwLrMUGxw8FVPlF/I+lRaivOs
qEPBSgXQmRhme8wnw/67TijTCBDLo+MhljM5NrnuQJ7EuZLGHUc68lhhpRHd
KDzuTLuH62mhkMDbOUrk9OZDLICB/gdO/wysWDsy4AaPbm+bO7a+6TF9W5L5
IjTUV/hOC5WDLDHyZLgy/PBVMymZVIckeaS1gqQIasimGU0amEWrKL6+pQ0X
PtjqgvIEIlgzk64Pf2cfUBYX2DvDRK8CkOPv618CwjtcP6zOFIcuA7GCSCL0
CybkJkezXXzL5ilPkJZ1kI+wvoJgpcCaln2vJZkJZW/8p5guJB4mXb8Rpu1m
wEduQ4031rei5v6lSpuIlR2BGB5ui4xOeTztm0AW3TPUfEm9sabxUXw1LxqH
491DJsM1gvpbBgZnuZQdKwNiuz8WqW82DZ0dMdOeDx7XjA70b2DEZE5tizjf
fhM/4egMqHIhJvyxwZendA1ahS0o/vvFPTfvxLan6hOW0XaR0hxCHLi25uGe
ZkC81zDlJls4+YPONW6OuwzowuJ9JwoolJqiEuin8oPSeZbALBqjkPfcDJ3+
JK3k51MBWKLCzhP4djEdb9YyUKstfVMsViztlAZeXSaVZNszhVwFzj5lKpHZ
W4E4Cw/tvWSYn01RcXTLKPCAxKIqhqHMHcb+mr07fyEIpCkBOwVzuNnOIs+L
hOyp6KlhNCgKPesjC84ZFGwHUPdp1fi4q72SjGR1+z6HU1JvFG3CyY2uRAQZ
WzKALuRiqNB76/AKLHr3YgzJ9JmeO9lnbNnxZi9VzG/Mq7wVU9XuDP8vtPxr
o9fKH2R7h/PhArVpBIJAg0GSgdSa/EUEnEkT+/2darJqX61Mm2328/3McPKv
h1Rl5crCWNxq/cZ0/+Cy7cQ+/IGS106NQ1biDSdK0G7rwpayHnM6RiTfJ65d
2F+9yj1V32mqRgIc5YSPUt/DcynPikAZ2kNgKmGvN4eH15ZfPHSsr+RnSxUo
VLMnu8m58e22ViGey33wXO5Mj0tIYrINYT94ZVmw+U8qwl/HvUzRoddoyBQk
KRE2QFUKn61AzTTRaB1/b7ry+mzdQR7vIrWKm6ooA1IqXt6BnAWbSwRN6MXL
YkRG6ilA6i2Vze8OoE4FWY/wUWLJqrQLW+fF42JA0FPeD8MzMEghklmJw9L/
Km/mqxcTIS55z4GexsDZ1qGrImiT1SHHiq3Ldba1JeduzlCb0CHVjlbL8Btr
Shesta/wXXe3JdOcUWFqTK2stMb+5RjVm+tE6fv2pcxD2aKEmto6NNiKJDrE
0CpYr6JYrlSShM1rlQNxNUAx4Z/ELbIIRV/sUCYGAY0ws1veCBhPOcQceOL7
VlyViblM+vcnid3BYCQeOMujD+6fQ+MWjHJSFtq/6sPmCIDt/TEOdFqve2uO
D24/E4/c1umjP8BOKA0kBPqAG4+2QUTbNk2eKQVOcRlI2SybNt5La0GS1Zpd
4/feYSh0CFZAUkcZA69Xk/zV9dFvfF/rQg/tFt3GmBVKY5v1iHkcDmeT6wA+
vLghd06TwSNeBrOwOw3RDYeO8m15nqkeNz7kSv8hEqo/XVWUuuFQ69TGpivK
GGZaE/j8DawRrXsmenOok8kyer28z0WiKfnYDM+2QzSjK/8L7IltZVqw5JrO
twqWbWibnSdAP4ASixj5zEz+ZWDPUN4oycshWPz0tHxll5A3Ss0F3bUEhZtv
EvWu5wJ/9zXqPmO0oIg6PPbwLUka5WHGEEKEDRXwb8OCWNBe50opfeRPpUao
Dv4Ki3FUq1x1uoaiY7puxRhVognTI2fHq3XXI9RGJltoEznnVlejoOGAq2cJ
kZV7j0+0gaobuO0FMgd2IXhY3xRQjNsm6uNm634Bvv/lu+LM+R7xW7mARHc0
5Xx4QTazauM1jucEOBbAe5Y1UdPLE6uIU1pf11fVKJDdnzZX9korXUc8aA9R
/sgO664OzU5JgL5pHhKjZV/pTBTHpkGBnQSzp+2EUguBOnEXsA7tJTtG6wzS
Gd+5U3LBSGPRxyHlyHO50L0TZu2m3NzGmJ3jI5RwgC8WqCJzvZ4JlotlSDwz
LKm3FJyRPtFk6Z63RPpQUCVQGG6oentzxjDJqqglbVEYkTLPeyWLlwNirxe6
YRn+9grVfAuONGElf5VRfobwoAPFfWnXZ/qlsATHygCp4GuAiwEJJWcvinvA
VI4E+sAHBriUwXxvC8IZE4KYIuaybWjvbnJQBAbZ6wNLw/gJFGKuxdkCC7xd
cRgzls2dKW3tNbNybvwTRxMa51Berwb1AqnD1CiVaw/toVKupgxLZEof/JTh
sbn8VI45avoH+xhnmDSckxdom7CrWlmQ/OAiUsmVyV5mNBqHz9JJahHUJNks
t8fsZQktKUPcpJklqzJhLGl1xuHB8axmADwATALtZ2t+9rsEA2RBJq1BYJIm
RolXqhXXry7JfkG/O9jDkKM7dxgAHYXyyb5KTnwQvqtuWbSCQheEPNPln+ja
fmHay8DOpWgybGNim+v5v507qvHD/6GP4WIxg1oRbMMeSn1Ly160EhOCKDqO
CSB4ctMPD8EIQur6N5Au17qGLNAKmKtq8ftVFYAocvBs6DK/rftu8jQKFe+d
tbL02hu0xg0v+cW5z/o1z96f0bHANFahFAdXwLpJmqbyzHBqFaKshgo1E3Hp
PB8ZkP/OZPi2YhTW6ztQugFw1DzIPzTLkszSJnLNJkFRazqKRFJdn0bisKye
rcneWc56zPlBpPXffzX0kXm9UwDDo/gqsxB/okEs9CSg/Eg09vp9hD4iOm/p
2wT2Don57FOgycCptvpxkG3PKcKzLR86in2IwiWWwm1q3dKQmKfxlQg+A7NZ
Gm+tmILQ2p15A5qPrvQBHeWAwCYTZHVjhn6R0J9axjxCiBbyPoFhycuSmXvx
4B66AbFIpN7ZmgUk4X9x09Kr1g8WmN9fahY2gvPbTcI6rX9bs1CPrO6A43SS
5PGz7yHeFMS1tRImmZpfGQcj0tdEr7pUFc7WhvKPqC5HEDH79MNgj8h8VPJ5
RXJB4VP9HL6k0Y1UEtbXXXyLeaEXXQ59BO8C0vJch3Ed2vTY9D4IciRDhQEX
oKZfe0Fo2aFoPEMC/3M8qrGCXKxwoKPh04heHupAOuuL/yluIzpp1Js1ooC5
lCdsRV45K2mgda+BzOVXe4n0nHxHyCopxrStXR9mVWyxCq4X59jbWXAJcE1w
ppWpmzx5VQ6XYYAWhE9lY1cd+UKTMDOaZyj451HW253WN+E2zDIe7zUia50g
Cp8YSiL3h8GNlCODgdXa54tiKTe/xrkZhGdEiHGuJBuqueL6J50g0KgxLhHA
VWdi6tDPGb41QGHcRiYEjPZwhG3H3LoegI41nnDyBgZqT2TkZyf/qdcjENiv
QkDiTKYD0P/OMYMlnNnLS/UqAf1USAHoZMKiIfFOBToqUjjVw0SEADUIOP1M
jUnA84NI90R4aRy5G68C7vUkw6WqIIMqFXoPsFls3LMXuOo5L1//Ihsq91S7
U21Zgu0YKMzX1QYEXBOSZHdbO+qqZQs8XfE7SvJI5d4PSPJ95Kp1BUxE/srE
3/1Y07+rDTbvJ8g/wCI/cFSnw3aCugwmDxLT1/yNwZkwqoTDg4jmYPQ4bZE4
UQiE/vqwIFO5dMcAQMnqKujS9E/CE7D26BXFNLNsLgC02TW7raKmZFbW4eua
paSnh/BMVhuS2pH+/HrlaQ6MDQTIuNViXrxjiEWEmv5Tr6HYahj/3QaTkooB
/n4ncO5RWLlTP6e8DZyg7oneaSIhtXWEV2iqdq1/edkeUufz3WgqjiRTllZo
BCjHBxbsWWW1I88U7V3wRJXrAwEPBsVjVvg5HxaT++tcGbzazsCNoNOzyixp
KvNc2U4O7HclYp0q6iOIeMtGmQAWpmTCoMvR/ec/M6AW2zk3Sj8EZXCKglj8
qcAzshkjgvu2L+OsI4n9Dsiq6qSqwrPu7P82w4n5j96jQ7pxhgdXz/Jnm3yd
o1+Y6cr5bbbC7Ks6WGCgiOasBJMXqzezGjWom3xCsMCk2LRAapy8BK7+wFS1
uQ9efPV619Z3MwPMiE/tlrL8dyMTOTUKrG4Ul4vPx0fu7myh4aJpwXykVPUM
pZNdTsw6QiOAuKqrdrVkLYSCwA58Kg0GChpRxO1CGacXkTgHg0Ig2ZOr6jcC
mTz9DIIoIWjKcf18RBkxbZxFGBOeRdPBTzlybfrM+L2S5Bvs9IVFhajJJ/H1
WahaXKVzG1I5Fk6FZqV0E3VFiOAjSz4Xel0C02b1dLtESrJNSrVvQF5wwv8d
t9s2TDnpLGrG6AH/oKWd2CG8XpliBovZ6vvMqW1dXp/6m/iJAf/Dn5jU1y2Z
uXHBVPTCvDNSG94g+K+KqbvLDbaH0IOaOJF3eM6k/Bv6rH9vHKRzE7G3Alfb
8SQeM0vSdKQCCKIrPcQx3wg0FYwHteaFm7ygsvwXH4bmu/5lerb/cmh4GTM8
lKbsr+uPzGUnzKpa/OLhHbJQCsdPIClrNo00c0QtBPIrbR1jwW1CZKiB+aGW
LfeCmpWR/iAqB7/vyGc4qJpTxORJHLPHig/dxxd8BsLsTyp/oJ1iwoVYXPjU
tIZXD0EKPyHgFGFH4aQooltfc6Qx0EVmUM+GSyepJgS5G+toyVDj3uL3o9oe
9GoTu8CuPi5pbEwWIcQBPKflWecYFv9j0laK7DT9DiLZ5BQGJKxYRTuwD+dJ
q9Fj0t3WmWo/Xu6+ttssu538BLhpvlQcvtRqnOYiruZIPV/+/l/2/zCiBlA1
C2MQHK7X5kfxQt6bhsYfYpqPiZM1UuLJpxlueZKRFVn94sxnCchqrJ0Aq7Qb
uSKQn43TN3IzxeidTGmyW3Qo5cQe4ia0xU8apEcEYvOPPTQIz1Jdtgge8bG9
IS353haJBY/eyNlaggNmuUJScW7TKIvvTCSOtcU66e21B8/T2ug70YnypyHs
LsHeArekjmSIJnCqMN3mnydcMSx1NQQS0uJD2es/NLAxLTe45Gk3y8hJILRA
An5fycPsYqJtew9h2vV175UPJW5WGzvYwuKHgWOAqbB0kP0gJ7gu0rXl2Y4o
4CazUzyJAY7V4CctH7FQjNIgkl2x79zL8GnSPbF05perVDX4kwHfvoGDtGXU
aPb28phw/L1JLomJudkDgiqAPMwcw7/B+BehD6FSs0oLwjTgKS/g7X8Ry90j
YPUPoIAqg4b3Q+r9i9MWLFN1Pt3A5OvJBKOQYMd/AJPwqWuEYck6047xNGu3
7rtUn8JToCSYY55V5uDHI7gxHfq4q7XnWm8bNp2N9uKynDuMWa4s3b8OwQBB
VL/c2qAUDf38DK2Wuj0HNB2vgLV4mRBTF2v92DMsGEcQ9d2S8//ZZjqic8pc
8/oGgGulcU22uqGVmliYZtaniyta5pPexcSZ8PN1OnuPirHZ9CEQx2T2WlS2
XZ6wllOuBU9cjaD/N+Fu2YR3x04Q5006PUCU8e7fzqr9/NmNzUuwPR2wRngt
58gXwsCzU4gD+ZnqhoaLLDzO/OX4w/eGSCSThO0ZuxctNKVQeK+xkKCGUWXE
M02giP79Di/BuCPjC198JWuwdd576O8gW99vc2pn0FpdG+ol18ZFXXNpsbqM
tOyKCK3nLp5Exuie/jnJEF65YroY0kHJGeUEqGnLNNHSGfwELXj9KuSbV4os
cYtW+pAxwNPhFbLvqDFSLXQrzHyxMugU5ciYO4EjMgK+a8D3jUvakXk3jtLy
24sGMazGX2+WEsFMcjP1b/fCtE2lLNOQiimnCOZ6TtVXALir1IgRn9NbRuvo
jqZI5zCxByho5FZcWl0OrRqReX8JP6IsE38/pIOC5nu6G/zWVCqvZSFjWnMA
aXkBt6JnKm776MPJrX22u286l3FduIKfvlRKQUPts14pL78ePU/KUKcMtwsj
rRTy6792w3RwD8wq/MO6hFHcKUbxgLoEzIdVTuR1NMi6mOWI13MfFwgmKYAf
wnbLRNeJVb/nuXPf3kBgESkBfcbmWieJgbK5THcqj/rCPc28/S1Jq7dlnW+O
IO/kEphcueSwL4y/UvMaa+PzsiF2ZWsJPVXRHEYYG72DHo2Q5VINzWKmNAXv
VT7ieyFDngsdgSoDOnuyReGaKkBZt94sbj82YzQnrsgy+cD5WdJz6/EAXZfI
pi4eBy36Orcf22clKXavnDgks/HNUNYDyPCUqWo4vYyb0ExDsGc/sCNNd4W0
UbJaL+Sf9Vig4Y5lTeYeTF+mU13cV6rf64I1yIFUR2nVxa4WQviwIj/pYrm5
j8LqjWPvdNIQFJzvZYZvSd7dSCo61zk9bOIVADMPdh06s9bGeugPPFPH9sHW
Flu4IXdxHn17sp14oGD1RK3f76e+JOFkNPzEFfeDcnE0mhiH38Sa1OWyuqWN
TLCamZtiQgOBTq1E1yRfdEQSRLUWkQ7YategDRwe1N2D2knN6QqMPOWI29+i
gVjEJ/HHsIOLzuTtBtLy0ZImJobIGXK4iy3yG3PgJ/euAGjxgUQMV3zv9/IU
dya9HCi2n4/eMlsn1TAgr8O5ZIrbVScfTORN59x+bfMbY23tVr3IWMnycsmN
2fbIRYTEtbtMwg55jr4+8FudWqWG55dNSKX7FdTPus09pYP8OGZZQKqvqWPD
0t+JxY1NQC4wa/hIFtKunqnNWitc26OEgVvwR/8gXSx7uhfNE1m2TikaEO7W
XdS3Wnb9EmFVfnpc84fPB3WtpNGvC1Ovwz8NTMAuAS+DY6tlmsqIgozRSY/l
+AF7M+AnT7nChDCtJTefbkJIHtqbMHgbNwUGm9hN8aVwkb9hNxSghCzjhXvM
59ov4AUWAtJuFoyXB/xmFYdR0OcRr7TM022ZT2DODOi2zz3VeHUZ8hU5Hdyu
TjXpps6MUIDWhI4P/GbnzivkkkS3zq+245Wuz5/XjwaafvUAvIErAxYkxvCv
ppr+O/ol4AhXGNA5QCdEQYj0bm1kmghZH3hfJdGfxKiK6TZ+5U4FR3+CxT5F
Tqh0UswJREYulcTND6kuoov3So+G2DFNpBxvVtnPQ8VPWmkxyKCZIQgr1XK8
sH8og0g3CQOM+nJqUEggVg+J/aAdDaAGuRkIGZje0pefTxT7lk8w66nPnyZP
oWcaCWnJLs6fJtrCGiOlcrcQAMGruEHHOC0YbWybVGKH1sDciS7tSyx7zsU8
iIGI5ubAj/uv6EqinrV08LEaPYIv7LvParpXiEUIspChjGFqa1RPsOaBbM2h
EY++rzmW4FqLZWjuR9msuPV3DV7YJdcsFz0hTHAQA8oy4KU7z4i9CMEXzagQ
Tuh4K+x8p56ugtn/O4bxEsvoL/zZc3mJuO7Z6YlgEYHjYiLgrb1xjZK000LD
BR4K8u+hu6SKx5SPCo/3C/liA03Zyob+gmeVSuaDLCnnB2fZVk5WM1cx7/RI
xNSQAYAlbU77fXMIVxAHpUYCKnopx7DbS35UPmAuCPYY9hHCQ9+D/O8LCKFQ
ZRZFq3TN099KSLtwpGa3qMntG0543xpWKafKLdC/Y5LWwZOdUkepS7VH6ZO8
gupE0OaDl922hEYecevFR53zq9UXeY26k9UGJ/hKdf8vvcFE4twgm+q8cqDj
OZexeDp093Q+igSq6qFe6e5USIF9ojiNTZI8rLWTdOOMYbHx8wTSF+YwPWf1
yaXp7XAGfaYF4nikORRxcQqX/6PD3wuJakZSeDpTFqTPwLZ6R8AggwvmDsBL
2H2fyc9ha5XmROfKMp0JTrBA161wc2whH6ndIEXBeytD/Gx+M4BYPFE8gg+j
RuLsZhZwpKfJSNR0r1urFhXBhQKP6uxr46qpkBqVH1hShHhETmZa8bOmy7pV
+AL5O5IWEA8y6Vf4X89E5DELNrG2Bn4GbsRYzcelig2f0VtN69vjjV7prTgZ
vso1Xe1/FBB6EJhcZmVTHdUsBgQNDeOiHRdaiuf6Dq8uvdL/OB3IEeaxsSZ3
fB8TXptZFBKQiIAKtJ1rPPuoD1ZY/mgEBRUEkpr53TiPnxAWysge8eFUkU9/
Z9Q4VDMSdQifkCNrI2P7Zfx3uiMJePBez6Bp1ULK/0cVpYxmxF+46wcM+E86
6zCsWfaQhPPTcsp9GDUaqz1JB0z3x403Hv3Z6pZcgtNkUgS+HvjFW1+Iqp6h
CaoDgRDsMEId6jympXB+EdhoX80xH1oxxqVR7QtKZMLSR6TeZiKd4CNZ5CwU
8PIWUZga6E7CLqpKqSRV58kzUQMteVxsfGRj4EMGyg6rYtbbEKa/0pMM1ZuM
MvLVh8MLNNdoGkWx9Y5jvfRfXBlHAlXo9lOAWlGK3BtQ4rzgyh5yULh5Ay+4
fT2VtSAN+EUkjMX6BOjYv77tlQSYPxC7gT5/vEV9T/SNaccerQE/DRAP/O7+
15zIcGafkUC7azqzQzJ5SatjB7YhXGugy/jXtuYv7x2gH+Trsz8O3s5fyPxK
M8pWdLwxjh+UnFEXAjFYVGyoT5ztcTnOpusfwrbdj9CjbaEPq7yz3FQeNryE
gpFRGSRsJx4/n9Fpe5N2w2o1cHLeapdMmNEliKkixs/rqbhFbg88zJ1ImWrF
uVmemoOtNBfaZvOIm8Aw1l0KOTgzCEcLL5i/uNC7z25Azi9VZYW+QmZe/KNR
qga6vmhA89LLREi4DTrZb73UWagp4aXa9wCPRJK2j/m3Y6xatMK+UzHQn32I
swkqm+Jmy0rygPR2l4pkjRPpUMI2sducb/Q3JVjt7aBi6Xw/11DWiBKFg/lN
6DhfAuJmLPZCEuyQVyfZRAVDPs289rozCpwLGBB0YohP0MgOKags127CAckx
0QAiY724fVDbXtFAEXOa3+ktpDaNh2HShEwddKv8TsfpaKqidWv5CM36XYnH
LwZLrll6Sn81dbFpaX261snXGNlvpVbHFMkU3T9+YVpGGMdnDUUp25+cfnsm
yYouUa8/o88gFjbDLbAt7WMR4xyZrMVBtzPhWo5gbwVW0VGaAHXgliLvyaeE
K9/IgDXyJsW1E+fR3QkKACUjKR9qSQRMaQUT6Kk0nBopCDhIfzrDVyEKGfeQ
hYmo8BmZcnfSZnZDfMT9Ecy54LSfdTgPjDrNySzqw0AmqivCPyUSpJquA9sb
Lgh1YFXN2NxuMG95roJnnxIrFOJxJ6chei9N/3yTvk3zQgnOU31oppmjZDet
hmkru78smU6EVWLpi1BqiAy5ntewXTwwdII+n2n73T7roVPwczuIdWCxSCLa
YlMDTjHZuech4WiGyqxqVKHMGyVufF/6S9ZExaW3g2ilvujpSO4gVcjje5El
XY4rUGTlqOPjbW5y/fvyD0A4V0JbsFFu4NDf0G3SUMXQ05wunqfhFwCoe+os
q9+j5DzOxHnrFjOnW0CgPNJEnD0Q37TDPDOh7wJMuKdOZmxgKrYmQRKFTHpd
43Jb/WIUDAXG9QydcHHUy4ED8xRE/h06LjaeA8IjLnAwGS4nkpMj3EjR7wbS
zGWLaOpKy8dJ5d3InjIIhCooEv4HqKNOKqEFxFXd3Eo3l0k27HaLq8YxngYs
1pVBT6gw7oFPZX0Jcv9oZpmNm9sAiq5CIKgZiskbtFzniwcRZieDQIUu7fAd
Rn09vgrgKSkLrmynId5/1jvuKjlPTS5QKMY/vQOloWLDzypsXSX4obzGJGs9
zNIw5mMPtzf1EdfUl29+NGCw1x34oJIG1Ksfb2MBBRL5BsJMH1fHDF9S2bgl
EpAg2IcVbd+qazarYWF/jusgBkMZCQ9Ov5HCde0ZywxFI15YRUIVeaAWGM/w
9A3WIDJPaMPgNwQHfMT4gUuUkM6W7xYjX2GYH3lC9YCyJIOvp+oau2cjYxOd
+2QhUeb4ESy4QsU/BsxbcBV3MQzVAvIOSV3fuMuJZ66U3Q6iFWmHXjnY1xix
yKd80gSLy1IJ92bF2PAEmNDEXL0Aos38zdiSb5xkNneelDUGDZ0I5LS30H5k
ZcZPoY9zJsvguBXFqdYetouO2YHEJsK9kyG7jSn6FCgK6bm/T2x6fLMzeXuN
6Qv7UdDn2R8b1tHHuqZunmvCstS+fF5V9xlzS6LajkfeeE2z3eQvQVz/Tt4m
qw/NoUVokupgJNbxrCJy7fe/5LgAsRVEd/3WE3OE4Vt2taFZ3HHkVrC/xM3q
n3Yu/fkPOSzN1Yh6g6PtKqNwF+48wppSwHgr93qjnB7vgX+GFXcEeia9t0s3
c2ztEXe6z9/ojjPcR02FISGJrYaeuRRuAdWDMUZVdVgZDomdfPRd7seythHW
DbsP4/WjlBigfkSyy0LFnzrTYJn/2mWzlV2Kk2uE9W4RIu91P2EareP4vfmQ
5oRJ5I4NbBaJr+/juMBde+50qM6AZKt6j+TOXq5YtB3HaLAyQlvjhCPPGFws
1VaLPXkx+PzxjjRO0fopEJ0DDDH0kbV3Qr7iQXMmDQFxPBcQ5HeLq8BKqYuN
BxJZMvjVgNk7MYH7gFMTZZZzpAyGH8AvtgejsKKI0JfC/It4WH/oMTsS8L0i
JN4oR6SXffDQlSLxCgGGkjK04E3qv+VQTyq6qd/DNp5thdODopcgPi/KEPB/
2lKgsTCNdrqHHMsmM13TzRcDfcKebxiyLfiEyhC7/0QcrZuHz+DmCSqmzk2w
hjrTJmcVOcSBxkWZtAyV1TVLVZWKqj+2bVGqGguFsGl3xg4B4MvBoMPLWhih
c4wl21Ego0mf4r6XWoJ/gubwxRgzPx6P7pbJb+LFM97fz6cTocS/Qjmnh49c
zL4gOu7axmLggRQ7H7LwUcCnFE4dw1uv1tnmP9jZhV+j23xDdmHDoMtj8yX3
wpPfM6WWXo4TTOH6jkg4DLKi4voYGvjuIHbQ/Zbff2iDsjknUHYcWpkSiBFA
TpnMMNjrXndA1gB2sN3zXaAdLlqWnV475DNDRc1GbWnFAUc5Qfr65MyhaUiE
8Zki7z/AeqnKnHTd+OWD0LGFKFzh+vcUxSbWB4AvHlBApY2lebP7FS1x0o7G
ImkbN+5j4sPAIho0ACzMU8EwmXDiz4eJP8hpQ33YKYaMSun8NH/oPxPg0G87
r6Ki6HX4OY13oV2OAyabyvCbrqVS0Se9Qm9aKoANHzNoNm9raJbzTzkhctFs
tFcTqZIWvJkOXHccZ5HGk0zgk2+ozS1MsCbFXx1hcKfJAgywB3xuPiv70Vgd
f2kjdJ/3IZTD/SCBEkId1bNKE5toScPzRJe74cBR1Qq17pqymgtjG2+COalW
9hWf8TeSEJAax4X3P14snVcifjnJlvR0pbBXZzVxUlenwQkX68jTWf/lf+en
QIryekzw5oZkNt9FPjpBhaF3C7Hyw0+RhPrfeA4cWVJhfxRjMoN09GAT0wWA
a16WLyM6aSXpBKRbcT/nC5otNJIcB9NtHdYUlddpx5FijIickDeyCZuH+jPM
Z6GLFyEcnZZLeFdkmDnPwSJ+LtCDinI1XaocYlpMgkEqwExV1HpAuwpS9HSU
gwZiFTTQ+qYQSMv7SeKkiWt2jR4fGkJBXku9CUrFx6n94+PqqnTF9ouvrcRv
fbUDuBCakkJHsy0+WeMtZod5ru4e4v63ACiFvVYc92isa0C96tZ+41H12Be4
wtXXLNTY9cT6RZpjLU5pyKtQVb2wYuohK3H5wJlcSPYuUujRwGR350ufR7ER
x4+2X83xEF5WrNA/bogtlK/ZhAphXGr0bgg3DkuoZtFDERr8bQ9JgvMzhL+6
jfv5lC1ahcXRq/9zMIgGtie6t9czy2kedSTA6jizcFVUIKH9DTMNp73SGrbT
Q2r3V4j99u5wgk20GVr1eZI95Zek0V+9BbtNip8725YPH2w9bcecP2RrKlQf
Gq0Dc1bme2X14F05527k13flJZzJ9nyGE58jVSy5LxM9ToTsHRZ5FK39lLv6
JtsWsg9hYP/EoWyR3xj2dqE9sFcOa3A3tmaImdnvyganmqxbwFPe5bBELMTC
AuQTG6mI6P+OrAw3U8iQ5eqPnSMo7BEGpOy0IGPr9D1vEUrO0zXe5GqguhEh
M9XHU0fsQiyLannWJNJJq9w4f1DxkcUkLs30l/VUmB85oqaRZWeodIoWqRVI
ai45NoJES5kypRzilGVgQJ2UoU09q6PvhVMgGwB3oqfVKhZUIgNwgAj8LRTB
U0sfs4kmlcSDJ4Px60fN/eD0Qo9zlFiff9rqc3kmJG+6YvXn+qGqLP7CUskl
8/WH9NUEX8tnz72KlDuwiEMnZ4BxGMrPzEIecgat2sZXcymhjTyWr+gr4bSP
PsKMb/TNAMl/aun02kywY3I682CU4JKiM549Ys+YO7HxgAYySFUoDR9vH7Mf
TXyNgo3AYUuP3E06w7XaGC0LH1xswWteIxpJT+OK3Fl2X2DG6MWDiJrKoM3V
XrMKmeN3qUxj8ztTQtchnsjWcT6lVW26qVbASehzQEWxbaV3Z7x7JD84q6P0
Lb30HjvuYtHpd477XjwUVjeuligDeqqGuNxQPLvuZBCYYaaAmHCqQsh+I5Y5
Ww9XyXp/IYIfg3aesffhG8xu1NGBdA4T8YK3wgTY36tO3KJKm4L1QWb8wpmw
EIpuuht56SkNDtxhKtYAVcvPa/hd5KPwtS6Zx3SyiS3jm+ovUgY++3c4qF+u
dbHtiV3Ey61VcLahMByEUzpaop6q41Ox0l7U13HNuLweZqBnRLuYGzKSgla1
HOgzdSC8hhMfOpOwXzF6BOBWhDnsik0ZAIcZpv88LEuE3p2eAVMUoDoSVk7i
8ll6VkZ6hcK009JJcapkNHr0S4b4t9mzRXcLbhZShu+fQvP65e3ZJ5j9lkIr
FP4r6FQ24k874++NpwX/NTX09Y34QKNmwUNke4yHMIQmXQfH/wrsRXF/HQrF
rp/wksJAJIPyolwD3lv4+fQbUhGxVVxnZ+Vw9TGd7Q0hW2LNTgy4LqY9VtGz
amhjcd1zgnbZRsOE5tD/se/VX+Duf+J3F2BsuK/uM584+gJDP+MSzAoZ8eVG
fU1l/S3UNonVg1y8CYGQXVCNIODKMm/SVpQsmdZ4d94fukZF5Ok+l5s8g4ha
zwVqgyopIdrF1/gVl0+1Ju3JlnT8xUC1Uop+g3lmGhmpkQz+vHeC4+rTIfLu
qufzmfkUbdma46y+qY68UiLAhp06yzNulxWi1tNwjk4lUQ4TIzcWipogjeQ7
IWfF0a4Um9uMsbFUaT8W8BRO7bGg06fpSbyh2bwR9pSiDZ46vXXZb3wvQxDv
EilqeRk6NQUWv3UefAKSiWglUUuKpKfCNDuy5TWEsv/uBhoGHuVThArsf9Zi
OjqjT4qH5+upj996k+Y1A3zudC8pg8ttOBT1enTOwscP7zJVoLEWxHHqZgGK
ftupviq11iEFLzI+LDZ0PvsT5cGpevAW3CvLnRK79pXdQ2F2oew+quFfTuHl
nzcQg62QGBtWtXCDWmdF6+oxcc7+10pbv9C8C7lw1fSA15ySXu+nDxE/fVAi
owvZdrhkF/3+memMK3V66KCpXu0hDQY7MCQAwvJXYSfKdXvpiaIIjPEoa/Ta
mUTGjOhzKUforbsaS0SvLLm62083qm3px/UmbLrX8uqr8tr6wsC/vD91GIZF
8/5A9rPXlfkGd4dF9T+J/SJ7p8p0445UPyDFy4NRFWt0vrAljkJ51Eueb7PX
22m38S9THucDizKJoHjcITPF1IZTl+pJN0pPYrox/hUukYTDARkI2cE/PxAy
6PG/gMb2IH5riiHMqSZp7CTURBOoqnr9zrK+W3HMvt9Ti4RiTXefYwpfeWkq
B0D7vYil7xcxx9d4m3LfGZvh/IHZbs9C1vWUfkZgBGK+1ZIlhr9VzU7Ovni/
anZuHvcR+qb+kewIgpAnkkccwQv/6OUpM2LMjSEk5DBxmRK/ogU0iWHqC2IX
WQcy29vJt2FMuFIyzE0OLL1ewKha5yGls4Vu2MfivI2FVJ1vs8UnD4/aGyPs
KIqmSO6XOCD6Orf/d3XLjqGGEwKEBlJF7o+EgJZrmEku5k957fgb9HkR2pWJ
n/mTbrP5anx0gK2+LyWBrsBpJLghpCu5CUvXOUGhLpAc6j1Svgta3YJfAPJh
poo/r/oOFSi7ftjKAY1v2fda9yvdg16r0hmKwVC9eTqysDj4QB3UqJsKnrcY
MzNs4SEXSq9Y62DuCBphRpN9POrZjZ6Kk78mybK+sO4yCgSuwfn9GSjbUqzs
zXqU6g/WWba+scUN5BLV5biOL7OxefP/nsz2uMUckqNWqfG6FhAxRZJ2fQKZ
BofM0BYS8A+eF00JdvpclvQ5FtRNc79PFqzEp8Mx1M/IBFn4VDVB+j17xeyN
y8v4UlKcVyOZcfcZ3Me0DR94xDRt5Y3nCgkxfpsnGHWQXeRw0x/IPs6aXAAV
Bu8NCaNbhvJbHIdE1fO1xGuGbgAy07ed7ZNdWyFLBT52HZi0MUMIgdlshGm3
uUkl+eFYA6iLT8dz7V35fmeg0z6qLawkItFOz/PXuMKn8l2cow0U0HZevDeP
TgjZmTNyIyq/T3ZGaUZ9D3hkRK44BhtFe99WHnNWrsEF2RX2BsxuMKMWDa4s
YgpCX+E8taEVOYrfAFlO9f1sf3QSvRJ5NSIsA8Jn1eWH3J8KqrzcGO7Y9HWO
VVZpKmW8cM3swrUt/KBeF+jTsJHm9IjRmVPuwNCBL8lTpg0uVPxsdIWThSWd
fYPj9kt0V5cNkNJYqJGwOdRCLI+aBqJrY0Glb658HVov5rMWz5A8Bs5207OS
mtD2f03TQQd2qLLSBIuqDCJRPWzMg/yg71CLPqSo7t7q9H1DDg6IngOVgQ98
1SOCfuq8REgK/qBBiLjqiHGNsfTlbmlNSplAiuLYq/brOPWqWvKuLX01v8zu
sz0gS2JJt9rCLQW+U4UWpaND4JoLbPRixxas0Ar3xHdEDcgXlHGIDaszPolP
5cFZK5cGOuI/NO8flPWUONlqdRLyydC47f4/i5rNNHOwHOQi+yqnijPtd0tW
H3xAl9SDf8tZlIZd8NlwW2dIGzcvCHnU0QMZQuu/CtSBUbN4Xsqm31kJ0yiq
s2XNL/wLzKn8Uu1ozfL4/46i6f9VwZnqQg2uHuzEJdaAEYUT9YYueWZSN4jl
iBlh7mQ4sKDotwOkKIihfXEk70HODlep0Tf1Ha3nL1wtO10UzCPnNAAcclpg
8P+vX0Uv6OqJkqkSddqjIlEGCl1p4exsL726mVGr+NcIV5m5mwgKR8tEzy8v
g0zJ4SIePQZQAGJD1mwus5scGfz/g02ROuV3Kh3i65XbAzFRXrowLJQVZ8pG
U6QLwJItQ/jJynK720yuTz7I/+Z4Lg00K7EX1f8lDhwrwnercBxB7oQYfBEU
QhrxYY4M81XLaqFEdabvgdpDecrp52jas8SLOgVBo3rO6YphbYF2Qcl1gsLp
6e0foPXt/ETWPrChPuerUrmpEcW0FCVPhhIXzTbzsjaxyPCTepEjv6CLiSKb
THqkLeip3m+L/aaB+ZA67XWuxN0Vjjg2i5L2zObkXEC8FOPhLlWm9XC6xNwB
0UEOMsVglEpOT/JzC5QhlXKztsza9iUXOBKEGA8iqHB/xcTthqsvXoiN6HIB
Mxg0BEsrcUJkOXb5iEFh23AfMIE+c0xAOsCjNHVwQKYbvYexns5no+Z47cYT
eg107bbE+CVg29/2GvCxBD7qI9adygYlO+q00xMWHQ7kccxZ1o+oYNhz7rhy
W/Uf0QSr4mg+3Vr7Vf0XVjAPIJZU9ofKS8dki2H02l2+avYXG7smeek34Cp+
Tamo/dv5d3370vnvQ0Q/FLJArPC/nd82kstaEQxqzao0rKsFQ6dEyxXHHbCo
myEWIxKiflcEKuNd5L/HeN0obFk3ZeNXRQhWNVoH5bUb1mI2TaM4wOKYG+hI
1hn+DMIEbqj45lkIEd46pGlfgHijUBdLke1MB7Ezli54InOvquiJ9DdmSPWs
L1HCuX1mjQ4ujTZYRKjwkMdWxVcsbm9EuhurSkJDhgRAGQmS6Eb/07y52SI7
+jXs1ztYB9jSSVml/Aitto8RMhyTODXDDfzgKIGSyYTjSZjqCzHVVuTUIGQr
Ur13xGvgOIZYWhqK1YLnHdnCSsLGJ+BQyVoMH9s9Mx+36AhmhYJ9CulHvKJ9
GqpTiSVbR5GberKbzmYoqyf/aKYYUI2/dCDC+B3KhFBKGI+V11BB+vfCIfb7
JwllLRKI3Yo7g1xqk0qQpM0kmg73rVU89vz5HA1DPi8vB3mExGAhCIYhn4jv
iySXuCYMdYM1YH04n7fOYLY+HMjEFcWKz1/8lqmb09QOCOfWEUonH83HpId3
v9j6VRImyGGSd+q/uncz9Wgetb3JRk4GLixmYmV5y8MuK2PLT95jxWbMIYOq
WZvaWpvr58rHIeT9JF/8E95QscooibEpPuN2x+uBptYHtBO+5OpyD63KBczB
bWfjC0vDSDGcoYVDvFxIR6dEQkFf8ESwiEpIlHFSn6g4YEfDWkPrxv4Rw6p2
IZmnPJz6CIxDKlFfSphQqP9RKIDGbzmGTKMTA/nf5ENwNrQw9UPeGEYh/EaI
41SrD0b7brqVi498Ga+w62HzVmSIiBWoUIUHY9SYaen544iKmcBD7PtArpG7
6d1PfcF9ZUhbu+kTUAskvp0dXtK7rW6R2+uhUvcDtVNYEfvr2rfaVhBCNtZz
vZvQ9kol9lKXsdJSX9O+es1qzvTVMi7D48/ByPKb54b/WCPwymRIAQeYUjwT
I0iNg3aTUPN0CD5s/eH3xXOv4rUxuBZlPV18WpsNniewvqUq172nC2++RJOD
JVWnlahAu0t5Uvng5+bYzWnVih5vJ7jvuBPq0Zo8r8CKRh3qIKmJI4FnFmrc
uLQ9sfelqhwWhVfgKgzbR5nlGrDjg14FJT1le2OIa3S+okqNsb4f/7LpnqTu
72urJcJUvHekG7E9fPkawpS88939PmE2OSrbO8RkXx0GrvTQwgIiK3LsEs85
UeSvM/PSNCB3ZGjDadpMOZYpGdVnV7lgeMO4JYFG6JULsSMDzBfN7D8VmVGT
EDf08r+2U5HZPNTD9PvJVmjHgHqrBlLn2yGL79IW++IidSw15ZqYe2xD9N44
U9uAV/F6SkqTj/MVC35dEox+KrQXDc9oRyeTrJ03UlQBIh62vGn2qBjVGrrL
qNOrWGe0z2C3b9l7nDC3hzMkHeAD5ht3Sl/p17AYOtzHosqLEQyIdxRAw/B8
8U42AUOUqwde6XLnDBIU6ilLjWL5CFd+aKooQrOy8I5lDieVnbeaNn6b7r/r
HilyiICDSFhSws0NKYGsw64vLBfA3xZV4TQE+ul1EmR1umKWvVxwtCIydhKn
+HqvPJ8DJu7TyCs7E1+vhNI4QBI35og3M+OCdLjI3IgZsO4rv00IYPH0H6rJ
l9MXBr3lRV1Nn/YLreOD/QZ4cXDX0z0U8kEJ3kSalXkNK6842RY2wLOGUNqH
3r/Pw3YutIs4ZypG6gFar1cRbwePUUoev9iNvf+xdmVUjuz3CcHZr4QgYrCZ
mpo1TyInnZb1UEknsaizPJrLhoNpuNC+1q1IiC4O2a+ApyEU4CH9dh4Vdf1O
IIFMAdz2Nw2ZEriHY+VssFCdExMwA7gk1RdL7Ff3H9R1FWBL9fAJtrgAxD0X
swBmgC6RDxCx8BL50ebQtLCw7b2xkhRGM8SYwDGbmhSj7zEVVdvwg8znz1uz
xlgj6b2TEHRkks8hc5WgR73BnavaP/owIQMeHe6IeDEu8hlyyOlmAeR6wPPc
MnWzFzdltv8hBa83MlDwO0+A5TW9oeSR0ZD1XfVrqLHy8GpoP2FegX0Rvgr9
6+MG0/sx/OxV2Fe0E6Bm+xA/KUbQE3SwzZvjpoGEq6GW+F/hOqO1FxSQJgRq
b01lYscNU/zjlzHE036oliD76xDWIajVHRdpK66aweig5q8DPHA/lOQ7aBg4
vkwQ5sreh0W93sI9ET0qerhH20+uBtfhxXIgqRS3eyfAZiFz3+AT9naAwTrW
Mjh5kQ0Wco3zOfOxdiMvCLbIziVBPhHVkIDlY92wPPqAJqEEL5/e74lnfmKb
xqBBMAsYB4lxi3xB5z2DwNNeU0c8pr6UUFf7CpqqvwUkTB/uYAvJCQ5LxDKK
eJ2k+t/QpARUms06clEtpcc3ZIcUOpCUXfKBLJEpf28HPVhWM20P04Q2UtX7
uJUeJ9Bu7SdxZ4o6DyD+gOJtrw90k8lKvBx/MB3PJIUVB8HbXYPFKBaPFN/V
qrRVdj7KLInLKuW1mCnlvh79KhSHbmnqEmRA3zDu11e5B+PZaMVk8ldIhQQs
kKGidziApP3CrAM7GXdVzv0P1YTcyr4zkVsolLyyHtmDuGdNkOv10Ny501wz
umU4I1emQMFUPZRpN3sqE0q9NDeBczQQCVwUmwClAA2CrQgJwetQVDhS4TVi
dkEN5iZErXftY1JBOClJsm/wVaJY2J84duOJiG0yu3bQgQe8h7l56y5QCEiH
nvY7WGvVxmoOWwEy1lWlX72odkN+NoJeph+ClcPM0Mc6moCJu9T5S6zk1Ww3
9uncpOBygYwrKv+Q7oR9KY21IL4P+hObLeB9BT97YJ0z5SqJE/FarReUHjHx
0Y3Zj0Xe7ap3Bu7FjkPPC2VZxu4P/DvQpXWm4sGT8AC0az/ITmLKXITbZvMV
ga9QMzGvTwBtwBuET3SJxuxhsN7N+J0ayThkGqKbJNGyiY2Z13FVdK7XU+u1
CDwaiC8d/0rKKlHMRKjt77I8SvI+dpP/VIQbzaDlb3bGAMRTz2JtesmVPa+t
99PpgjD4NI2apOAKIW9NCZS7BWNWQPouasnGlU5IaYtkWIwDRpZj9j7gVyw4
BeX+YG9r3Rv/j5aDIkrU3yLqO14sitTleKpUUJOP5xmTV3HXULF/saXAG71Q
UUOaBIe45DP9DIXN6kAg7h4b/Vu4CQHWGETGm5BzmBlOybUtV8ALxMZTuEgV
sINMYfeXcS44wdaIkPwyX+W/zdSY/ihV7ZH1B/AtcwhMBLyO7+N53u8tBd55
HY6tMRSJVI622kBkEkk054mvYBKmHHj5fteUlaK+yJQ3DaFDiPCn5P+KuVSE
Lc8XzBAloYB0InUVSMpX/bd9olvYJO44j2EWy5UArSMBMLYY8Jf6nA5L5qGY
mNce2lPYA2Z3J8e6ft+4038uaW5SjxoHJMOtGzOMErnMDSF+SwPE/IhnM8he
evBC3dSMO9HDa//PgBp7Ox3VoxDZldf4ISURO7vo8OfmUY7dJz16BL3x70Jz
AyJmJH0moNik5z52ptGyo9IKJfJnobnh7QavdUu6ldLGpkFO8mqM9kr6VzAo
59X1aZDsAL4WqqFlMrIbnKdDr96aJ5ZT55xwMvc4A9nTHsvintck8mHfW4Uk
3vGfxuukWGBVDNo7BNBpz4ggxbNC6X+AkYc0vYCgViFAf/JpG5/Dat4Mn7bz
vq/Xjcrr4oYMJicIZ5FWigd5qhRjzvQJK/kzHWf84iNLE7Pd1ZPBCKOZn4ve
Jb4vjZt1Pz+5/jjJyMNrGTqOru1XoKcCCkN9N2MeToQZX5KjuOtUwrYXLk77
INx+/ETS1mJNJ3VkrdmSEZR90zDUWWemIPlIwatXrjZF+zOw7zlClPkGAQBi
TwgbIppRLqxYVuYnwTxmFMuo8g8pRrSQF1f/4BqtlNJZqG0grGXCgegH7uP+
vvjtFL5cqHu6Dmw9q27JowJb2/pqaCoVTU8Wg2PYpAPTaFEUMp5+/upfpa1N
1IpGRSNqwI6IeENJD5wvksmVb0kv+Gd6tO7Z5LA1lLZS0pXmFBipDgB03HV/
zEXmkNxw256ojmliA+K83RGKA8knVcNdYvi9eqZFtF0le386gWHNTloaI0A8
H3Gjwu+Kx5iLB/1j/R4dC8vVEjW4opMyf6QB6CzEHFv0Xi8DhZM8q665eXmo
1VyF7sWa0GLzM945cKCoKLTVJ7F79Tp29+Z+fRBWOb5KF/mrJgT2seLzHG5U
BkPj9c3vvYI1f3g8WtPmB57lX/YbPhwXARdKLHmPKdATy78Eewub+nyheP/G
XmDZSIZQLVsyhgHpGUQXm8HV5Yg1FNWt9XznzTjg3OEw/wa4zVYxbmwAc/g9
fFeb22dCTggXSa3j0B9nk9mW/bZqUmWLsry9tmL0BFgBfqqVAP6NBBSsp0FL
RoFxkb/iqkIwOfbx3Mbz6PV6QrKX6ZD3swE8Z/rbqbdvLcsHkQOXlTThJY+5
SYnmDxsA1yCINHGYQq6DRiLXJxlo6Sigu0fHzQN69gbQbDXFrznEfTwRi/R4
YAWsS3tu8Uh+PDNmF6p/YfcOiIjO6AlF83cTmRr82PY30cyrFIp6XjQv7R7B
0YRj2X/Zy0cKy4oplwzrQcMx5p0VjilrvLcFe56tSvYdzpDurYJUO0+7xOOf
cdGoCs6vtguMu9T0QPOfW9tuloH5J4prUMgtv3OiTKoKYqKStCyoTWsMAeqp
wViE7J7RTYqAhW0VWUcpWVHZEtovLARoFqlnMkS9Hjsi8/LKMlcDp9D0qL8X
uikEIkzDTuT2d0/44B2+m4fTfRhVvwvs1QykYpf8/fdTde51KUym5MJfxUaO
NyLfYEfRKverbm2xwzs3AZ96Vm8dI2JzvByL5iUvZ9cicz/wvD9dL1HMHOJs
rbu20FEovtxy4vx06bV5zNZwyDsweKYvub6DgnanxY/SccoskMZ12WQVs4Fo
qo5MsEoeNjUt5i3jpmAiDfx02G3Bcwz1IJdSl/Gup/eohZseqAT8izbjEDvs
T1R2ZQz4MJV2yy/TXDt2dTNopPSGY4dyyJyLqkgio/9UQRQ+1B1bgmIN+VRt
qXzQsG5wefQ5u3aQgmj8w10ZSKmxsHGzMWYPcwT/jV4xKYfzdHEbvmMnFeIO
ydpgQNRlqk6pBkIIzhcpaEt2AYWh8/ytSmKVTbmjYvJrSRT1IGFx6ZARWXUk
vcHcCdB4fCU64VZ/lARK8G3PyYICJ76oA5zIdzkUkI052j7C9RIvmiS8WPGh
8Z5gVyUBq9BHGn4pkCbkb1jckXmwKuhepnzzyC0CbZrMDWFeloLikZAbov2s
CsO4adTu254nxBTsbiU8J1BqBhJgZYBf9ygnv/oVOzCwwqqkO+zodnP18B0D
mRUOfQ2Ltyy3FjD+idUb5I1QuxZMA7TtCRjB5yezRgeBfx2LNLACADDN361o
RrMP8KBrgf6FD8dSO2xV94QnDyp+STF5drG3q9N9sc/jZzakeARFf9mKsBmv
PpIexM7d8AZ05olMz575SM40CLF5vYtK3GfRJqB6mPY2d/WHs59JGfsVgW2m
K14qZBt+QyaYH0HsVeQKQwW37UBbgzFHlPsKPER3Rgomwd9hcG0WVxavT/pU
bodvDdM+URVKGZk6u3Drjr/32MAk3JnshAsv1d4zhMeS6lPC7vdqEB3K4A+x
4ofM8EkCT7W5eSyJia6k+jZP1NtJmxk1QJ7EFnnTBhESHhe1Z+hJS9K/gPOs
ShglXYu0QotvTJZ4gsXmnVY0x3EYbz/NR1eEsdK+gK9U8ndWGCJrDEEhQSMx
DxL09vkxkZQoL2hXIZ9yPB2AqErdZNEPRZLIlYjfkhbFVQXBuZfUsbVCEs/0
1V8iYji4y5dEvLhndQWD7ZKOEt+IxTwjZ7/ULO5/1Vx5txjH4Wd+jd9Li5b+
m2BQJonKvrAD0aicY4BfivlkwJFom70CnBE8wcof2CQd0V2XoO8LlOOHUEm4
kEQ0WM3RB3BhYNdUybrbofinm1BTCRzVpI75GG/GUqhG8ogpAS+2fQt9pZvx
3xK3SuvTzA5J2OAcQLLBZylW02ANqfckNZqAjI15xrT71mOx1/tFiSA+dyu4
uLh614dJHe1XcVoXvEXnRL29zXZNK3sn1Gh2ZiPITP5sllzUpTzb2C/mkNro
AUK9fWKgiCFgS0O45Q/M+n3/4GB8slAnPOrBmje8zq2Qn02gGChjymJuYO46
KyPhDjhgp+G4PGzTmZk82zn0l4i7wBk7u7L31N/fucFdP0MlfHrDLDOqsY9e
+BEGLe52B60oym5qD6j1UJz7AzBQViwmHN5MjGBFsBH00JN/S54p9cHfMlpj
zskhYqFqWIVMbMCSJzRuOZ8Qyc1R5dLyPvmJRSiJ27SMGA4ezwER8AmQZrat
Gzr5LxAZQxd0bJfMO58PZmeiQoIzY1c8WpazTxBqWs0hQY/NHzK9Fmp7Ju5R
ocUQO+q230bmSuqBcRUmotcqv65r0zDvQuFRRqCnVenf7w1r4cjHr0vN301f
tw6wBRs99p1iEvflZ+vJus+xwADBZ+DSX+8o4BfxPiZT5u6SKQjQ2TzPWLVO
TOeEksIm/FUrrZcj16NxkcsfltEi1erFPQIxidl/UZ3nSeXcweKvYE12uJCp
mc2nLZbm1C8J8JH+zFzlH5Q3TaQJdhxSB3oMDznJ/BXfamaTprrI2OsEH0hI
xD8IYdW+c7SNsKaI/01IwE4LawOMuL2EhUEtOo7JSNc+U9FqcD0jMqOi4Mt+
0wzzDxsTrKd3PSfBepRWr5BGC1DAkmoL2k19Np14MoaVg/r50LG+TnHeKLeW
ASPXfu0hf+COqIz+CLtENqegpZTFvk+S67gYxdzGu9Azj5gN/loFX/WUKaqL
BDVnE2pJ/rK1UjTjYVNUDIz8skKbzPgQH/MxNB87ZYBkyis1c/dOv4BX/Zci
ACks/LedpFyhUpY16AW6/MuWIdbWWRHndgUvun44U9Tz6gTDwHQL88a0Lin3
9jxJXT1q6auPTfFhasRpxVGlWCqm+09FLNlmtuidJCoU8Pow6Q0S0TaIWlqa
cyxmy/e7iVfXEAdiP4EmWNlOLU/zKj4liaFW5SojKx7ADjjJudscPm40WMB1
UvBiuoWzHNUVukJyLfA42zooVC9qFjYYrxAGHkncn1yjzJtlFZrdtmHRtDTa
QoemepfD6lcvVddqS+976ppIZNeqRXWLzuEFZ8PtMkRx4igw6EWxkXTgaGWe
qgqaoawDe3JydvKAy5e/GAE6f17tD9t+RubC05FrDMEV/ACFjOlXcp8zrc17
zoJEVc2LdqRT21mYW/MmECwGYdcUzOzTI13QN3r+2ceS9w3sdREvdFr2+D32
fr4R96Btfp40VNKllPbQnngPaCZdT074lN9zcDiZWVw8xfJJIMRWSVL4CHo7
rT3ktsROKQdcljZuunyUwK2FgEmVB76PYitEl0KQDiMzv+8/xWVp28b/6pjd
tRl6SbZI2xrVyZBmEKhJZ/84NlsgjMQgYc56MM7rNE89r5MWe7NUMXAMCUto
h11L82Y7p0Nj03m16/IOwkKG8ixLjynDsy6WwTv6SOaiu5La1XNBILojatkd
b/n+CuW3fIepOHNAEjwkeJwM3trsZSukECYqUs8TaUZ4/6nGLOBnwEzttNdF
172MgzLBmvhVC2GRW5FMwSrxNHgxcDaBrCizHtwNMMWnlAV16iKD+kQXSTZs
dpSJt0kW2mXm4fJY2DfqJYPFzP3Qtc6/Axeb9xytPbV81ocJ69tgR/Wqmwra
tDR8sueceVjthszG8aXlji96RaDnnv2ASJgEtzU9LXr5w5Zib8GcDPJ9OYL1
7BUfylx+jLq5IEfM9NhWnXQQk/zv2KWFhQVyGLLh3tTI+/U0VcQRaQsBSiwm
//vge5lFIjO3KNEQSvlOeZKK7EdOLILAomvH7oyJmWa5G1x2ZBmv8LEuoFIN
eeX5Ll/CZGghWWX2kTyF+5ZjCtFDNOFegcXj38Dyj+PLHdWzK9OrnnqSlEFp
c+3Or5F9XI5EUHWqPXSusbXoHoYkPvO95LX3mctyW/vX+Z87bktSXzk9Krjd
K23rRbI+4A5XKv1DWzmVLh51rHrKVFGkNBeeLznV8VtWoCA83ysefNCz8nAE
BL6/hrKWYjiKy7egIlLxsAPRbppDNj8DQcd7shivZKSxW+7eNmVgFVdw2KmQ
69rZKhsM1Q+JVJGKsc1anzYiYZQwfLiPAwILuGrnBeupF8frw9lInPDYvVMR
7sQ0zJ6Se9pyO7zOcSsgomLe7Ri8uxzR8VB3wpuXeYD2oIXwpcps4/akLuGz
1SE2JpPNjUZsRGtr64Xwalynj260O8lJxD3puL29a+plTHnqnK99lVwtPWMQ
owOJxyqz/0YqJr08ni4I2UHLnkRBsfRjf/zTDiJmJFsa7SdJ36OPE3X7driY
3Z7WoJmaDzODpl7THegEBiltxZD4hFlgYTn6LG6deF3Q8IhtcQEBw58Whyvg
jraDC9IWVj8X8hGES+MbNBePKBu5wyGgjIxr+mNll4V5gGe6aYld/tjc7d4D
k9v/OECNFQt+27e8OkBFzKjmo/VFpugZYTv5zcGjE8+kVqUPdD7/FyJVcGKL
ZZ3MN1463wQW3HvTP2iQCc+kHxilKoriEWoqcsixBiY+15x5rNOTPXMOJdK7
o/ZulsowqdBoouUTxeSRqzTBfOPJObKR99sxQ30YvNpECTH6jrA/XU2/ix7K
E2ObR+VmUoz5OnqCtjR3mwW1YeArxbCjDz5RMOR6meZLBC5C+R4gLX4Dkfs1
LCBBYntupgPAK7BHXGfoe5Eo9C8rso2c8w8UEdtUmPYZIa2OpGRzTX9x8ERH
oey69G4foAyRjk1s3g/A80Na/ynJacZ8ws1PlNW8eYiCXZQo6iIm+VqLoltN
50ArmHCuLj6+E7OUYyLvrPx5jfYb5XnQAFzFzw1ongBmAX0xuH1ItAwRktpQ
IDhBV4lwc+5oQzaBTiq0h9y0e5aB2Rd87+9I3secGFnzo8PZn1bH3Na4QIdE
aRUU5oJJtqjbHMTzLidZRWrMC/krQs7+ckpM/TR9SdGBI53UYYe77lDBps4n
ktJMGxgRHh/8MOJ5MA4IuRbJ+Byurn0yIYXNjK5w441BByy+btok/2fSpdlL
zOgYmyxE1A9wmvC1D2/Xnxs2dgi4oXnPsuWj9Xz3MhWu5kMmD2VOxcqcZ3wC
7ghNSzGiOZmpi2vcHovmIjVjoH8xgaaW2RsSz1F9NyIc/5YsiAmO2aM1mADm
rsRWWZctRTdTygRvsRC/CXE6HCI2iAZD8GZFN/BlpjRHFqC2HM806Iv7nVgi
Ubc16JwiHVTDAcf5NES7zYe5ICdoID+VMg9eZPM6KilwsdCidaC0DFfZ4khH
0PVb6oc/nU3zDtRx1dZCjWRywU73ePYkIZUaL9Q20KFP7ikSuYF90wY7IbiA
a951UT1nMxuhiD745oEmKL2x2rTqUcoRJX2UHLtwQA3MJhK9mxYI42FM52kH
YsVa1OLder4TJj1uXyIp8wYZd65UlqoEWp9qP9KVXJ2Ks2XhiMaLvxuFFfta
2hXJAHsqgp2sP81N8jQ9IceuzHrnD/3pMIewQeHMJbsI5yLDih0qdvT9M1rk
IdA+Ae80aFtVbO+qs4B+0Pp4Zs6mTkZLPCe1ephYBKbavhtXsS4KbVW+xF5f
sQaen6FJ64BhQrgwHKotqQzVd7FzLr4JRfz7pH5wya5sZnSA07nwGGc6GBCT
5jJmzW9UCO2pUb/SNIWo9yca322gZzB9pz+/sfOlbMwYxHIgI5vud0QCYN8i
ZtxQiOPIIxdxSLM2pJnRmMtt/klXNI64NKYmaJM6GVaicylsr4HDFBDktPs1
V0Esa/dhxDdFMzdHxz/0Iap2zOMW3p0zjjS2uUD290maQDMVa56Omi5efs7i
iNNFNPyiBiIdBtGmFvJP84Ahuv99tVo9011sVXJHcL9YMuz1zQfFp9Xm5hVU
oc63saH3GUW1v4HF+mnd1Nb4kRROKfpgaGtHKKrX19QNTJPiI2EcTFF2mY9/
erjGPReIqY2vHzG2Lf9TWpzc2c73elixfMiB+YVU+TmBu7I6AdUt+JSQmn9o
EixMFuUFCdmQXGug832POYzQmm+LbXdaVVMOUuGjSGXokibO1HpfMZKYraTT
RdH5+rmVSQdoE3dNgVi/9TwNFofrobYW1PpgNiQr8TVVvoNuFHDc6BfBL0wv
gpHlFAJQP3L4tdpz8pXkYU7WudSTewhJ5X+pA4VNpWxHIEk7TQn2N8dVf3nT
NlScEPMqjJrlj3gmNR6Atg1g7JJzeHrJ0dwweeKhl98igV3N6+gEg0+NDl1P
/GxHaWe413bAcEy7hWrsZ7lfKQaGKUECsb6UzjharxPKliMdEjYI761cii04
cS6JFcmU5HymqqfYQFv2WMLc2MdrijpF87qxwuYfC8K3pqNRGAa1SqtqrFbm
FDNvnvFlIibdGR1FsHdtbQNyGb/N93RJOZ4ZfAPYGMAP5AfHpG5ZEovs2/KA
TFCql+HsSUiecbkgfiYAzfXKcchpg89SnknPwRJkb4o4KJbYPpVg0+1z9c7a
hTPYjvO4O9n9rFcpOek+u9oh2WrPnJJlMuyO1NT7o/7YqS35FnyVC2w/HF5x
Y9XRRwmR8oZB1K2zu70GCy+YrRjV6dAGKsWdVNU2sBRQoIEOuIHs6Vd8NpqR
uQY2Fi5RugZ9CntcoukNIv+WNMD4Dexo4XSh1poewKfMKZOKSjdRjufVy/uh
0rrnG3JalaoWJFlZnKn7YBhh/eTvNPZcW+Vqd6BDgsBRCMducwwNXo/lWWm3
JxfvmPVOsavcONnwvCyLGLy4SYPdB7+bCR4pGOlb2BMWoAYBIOtFI7dwWo7d
M/5s4AZmKcp8LGIdzkP2tbXyLIOK2/Y2xpanpjdd/JkJEvE8Zs5HPKel4VwQ
zQCfwjBRcUvxVbam29x8lKG6G/0Gh91Nqnlwwxlzn0+O4tcetdT/CeeLUjHO
7Kq232pnChpz3w5ij1zOXFncTn+vByFDCc+xShTrfLgtsDaFIYI+FeO6YGVD
KunR8YJTo0HENsAhwLmzqTdZA5SzCZZPtBZYr/VGHxOPF/aN7I/wYUSTJP3J
LHTvIll9eCT0KXbTcm72GUTsn0nJizpZ8SBb0q9Vveqsfn/CGwUc6u/QdV7E
JypjVTVTxTTDBSvK5jxSAH2DS2zTybxovy+yjyPGKxxn/SJsx2Tn0MhL+wBY
k8Xp9oTML7gqYv+IsLHsIeEfIfKpt/yQI6qqMgu9bpVG/4v7cNbwQgIv1uVc
S7osx/UPyhcdf/OlAIMh4Ms9gHPzS6K0pOlRB9VLLaooz4t0F2VKoLCiVauH
D0UkAZx5N5CXrtuiPZ6Iush73Xfg8rF5JSXAAXWva8NZG2GdDn7aDq4x9WGx
jU2VgXU93l5Xdu/RYMagXXekxHldT+EVaQv9tZXLi6G1uFWgM6o4GMnS7/eq
KOgYsFUeLnf0opLeK6DaelxKC77n4xe9kXPGWcD0LS3T3G+G9ZNx/EmTzr2p
n9uPgiwSRijzf0CaaQryNCX9f93go3/2Z/zR9qPle1/ow/qeIWOsE54mHMVn
//VPkyoyDbU6Z4WCgQ0UoBECZv5KAoecJvtTBIbU0wJDrlm8xVkF5K0Grce1
1xsZztg7DE5PZL+Hr5rttB6nmMcL8Oo8Y53F1cqLt2Qfx684DjGY3HFLCdgy
uBQDbRuRELs2a4uKOAtYlJ3tjtd58uy1/ke9ctFiflmogu/8bTVSnIg0/PNe
PghQzA1OWrAU2qiV0p52iRBQ2XjSAnaFMlRLzomrhnACcaVxijOKtDIz6RnO
/aQjET0mBhMshMpYv3ggoxZS+SoNQO4JTzDzuOaTijqZstjsaQ9kTev+E9Uj
0JsHxuPvgalHgblfO4rBjAXRxrhOphT8B5MlFduM/YN6SVMrJvNUQuq++nLg
We9mMQXanmQHWYIWMS7vXYWNP2S3XhPg6f/QyXWvFs1icA9xI8fN+ulp6Lfl
Q1JGxFs362NBAPf1uneGfr2pswzuQOeLMOI9i23+wGjmf7oZ7hdpIN2AgUzg
1wEfsT2xf8fSNn9vmHyI9jBD02Td6luwOqPo3Z/NDgaSWYmd1aZAcQx8FKRA
5q4XgDjQ21UqsDnj6Q1wTwat7Em/gi+U/3hsa7DVmjsalbenBcXmGeefWNR0
fQcD53zlJbfRn7AAMziJ8JxntLlqGuS0bzyYMUvdnbK7IOtUaeO1b6s+MLSB
DhNWIV4fNQzKKLZZmwgebtKckIXcpbmVbUjrs1l0Dnahtp1S9XyZnXibGCll
qgPyJQ4EuVpBo8TIzzWCC5ChWfJEzxW402+lpU6gMti1oO3vN5mHgcJA3e90
XAeo/YZS5i4UihyUC1U2gpfSoNtoEWRJIf9AmMq5iSOml1AfLk1bZ7hSM3Or
P+hG0DrLXgByy+UFmn/7eDgu039utr83zNsi0/57irhUHHVYPiudE4VWC3bG
E1kZ97068LYsq878+EAKqCkf7k8qJasKoQENcFKewWbdLlZop4n6B7ZIlTz1
G0zyObJdU9gn/xKV3l6Pi7e8oyLcXAHHSSetJh6qOa8OKxGygAVeZjISgAxD
/IaxQAp1OCY3NCuNXNo2mLcdf1LJhF4wAqPecJC7P0yjTUDdyXxIDx+4mIqR
ZBCOUDcueUM0nag090SXYnylgISZ7rw8FZMuyszdBb70vS1u7hxolMXeSUFg
cAwdxbBrTKz3QBgAi/4SawbU3nAtu1f4RapOV1o32OFGa02sKQuk+I3cv3QB
8cAUR334mgSvI72/b9p1gECgxm99ddO99VJVFnt7HppMEq9AlOtCA8DBmFB/
hyjTdLoHKzCnp8YgNSg+jDMyVnIR3corZb0BMlxplOGkvEZlgcbyiATXVlGV
9/1YhPU1nYn3ci3vUKEB75CbEbPQTFTNnPe2HKF+Mz76eaFzyhXRjzL4rS8V
M+L53qkqIlvlci9PAWSuiTpdnTFIwcHtsRii3wFN95leyoJv7yEP3Zr3p82B
sx183h29wLuKUnIcL05U0nTc69xwjQ6gvU48xjdADtkt7WkgeYcIqtLsay7p
WTDCYF+ZgU/GBZvFTA3LXYdq6L4zou6ZRMn3Ox7ZpJmmAaujLmFC2ULRlZNy
SB0clwZ/yCQH45HLL6ieDClsfhb3kGlopmnu+OkqUR0wpIgB36hNDV2auFxQ
Op1Gnq4IPSU0b8Rr5umUhI5D4sVr6S2aNydsNZeGBF8ge773ehNAM2OhxiU+
RTVtCKly3xL7+05MtsA8rYcSV8mNfikVbnB1wbhIXJmq5ZyIDISfFnARsDW9
r9OGxo+6pdqmcLz3MeDeHwLwMCjmVw4a6eRz29wS2ZashnQ6VV6dd14k7sCA
UVFScR61ubLHjtkUHeGXThq1agsHp5v5qwNUQ1tKFvNui5j5YiHWjDB6YoYd
Y2r1+CTDDHfHFTX7oxBV6iplY1WjvVKZrsVQifNGNxYQVfTUWIYr7uRcCP2Z
PLx1aYEq+1cXxuzD8iv7AcqSL4LunoTFZpNRUem5IRhmganbMqP8GFu1l94U
zcYC4IlzMmBMpfDtB2IhTzlBTeSr7chFIj69xr2aO8hMnKfqzlV2hwndet+r
g0VRBWnIfuW3jVq9awv1VPunnb1qgCQKb3dPrTWTywhGpiuH/EVrGD2TCF0G
ql870Ut8mmef2tyU5DUhqEvffOGAPoUR+X/BRs8fxqA5mrBx8RYpBzp+Q/Pt
H4IQsxArlM2z3gBHBcjl0oDKdOCu1ZDOIvJeRPJbBfokGzGrvBMuULcK39vM
owgtRUn0MNwlXtySaGeVx7BlRNpYZoOh6mE5QdLtI29G/gc62igGyuq50PJM
HdmpEU6SxJmF1hez8QDBeOUKzEQVqW6g5yU4t4nuMOpiIZjPtoGjMwlG+piW
zbAJm0wDvS70BETKKNSGxjKZETXdL5yluRrHztWkFFf43AXL3TkQsTtlcAmC
tZs32ZOMOKy3HfYaaHcvxnOJQUOX/MHkgIAhfSD6BYrm3FJQ3u1aob1Tsv6p
Vd2VxRawfzYo4em8uohwVidzNPiKu1hTg9i8CGZgbwP+5laYnwqMC7brHGGG
dIooRyShOSUAdMjk4vhcyYPp8+C2bl1WPvxvAB6IPq1SwcVfqyVgudFpB+rC
qlyPqLdti1hxJ7pa2othBvzSIoewpFceE/V9cgQzZhECrgXLD6SOigBN3kid
C1Wg+Tu1H5grDzR1a7VQA6hRG/ItuO7hxQtQLgH7sRLQHWxZFT14uBaw23Ld
f0A+UrwXhuNMur7xzJ1Bzc34j+OwiRJqFdUhIdseMse6f35TFz/XW0NPaG4X
8zPB46ibvkKHWF1DYgQsPA+MUl+19iaskqRPGRY5Whsqm81ibHxv8jW9aeOG
yK5GhEsmu5u20bE3o4mthAnQPkVT2njjDDHhSOl36f3k21H3BAEIL8pSgNFe
vR8f/Ks078TNpTDXWcvmgUU0brChymPAIRpsgV+FmGwxjObgBgAg50uiRPGz
nR/JOuzJzIBj0iwGnUpZWsYpawKn2oMC+XLJSAZW29wrzLaKNxyXWp2QhcWW
j+s++T+8XWjRioe3/xiQkwnnRaI7+nhUzcLUXhkFrPvWIYAaJem9Yf6YAysZ
nWxbXn9mQGBUhtimAEjcZa10Sv6/aI6UgMqd3sHSAex08BKLRevT9jCVS3GQ
l/pGxw6AGiVuBkiVOkUJ/Ok1d3jqZClP1IeIW//42FQhaazjqbU/AnKTHN9n
UmY1zSTB083YO6VIN92aml5XVu4nq5IMGvm7Y1ee+EzqoE88VNEeIsSkGB6D
eZDhRicdYXVXx4tJiHCHCauP3zo0wZ7/QSU54mIk4uI3N8ugJAqXn67w0Sn6
uMidsgVNC07UqnZL9v0ivFiWoAubmw1nIvsJsU8TnfKAU0uIJHN19njtE/n8
5iV6jSF+upsojA+C8opSE1lszQmIUfPMtrjo4/4j4XenTbW8ayApFj8q6HJt
c/uQgcINO7Q5kG2dWWfoVz8SwuzNJBuU5T3tgJYciiNYuQxRzYdiOZtjN7Q9
OBw0BO8q2OBXfYQhv0JhoLOMAy0SYoDukh0pR1ngwMnUsd9rgel9+5Gtqk44
pLlzjxgmY929Ovg+2TP2gkkXA321P4azYEtH1cOBtzCGRI2Kw6gc0uuZT0Y3
l2dV102aS3CNfP2FvQY/pZfN6MdOL7qAV3iraYBs3zM5W7N1/nGM71jUSUXB
WOVolRdzDA6fsC2hMLkNAfSXsuzSjRh2XY3S8KUBO/JHBc6C3TTTJCur0AuI
lusOX82rHsgcbreZRxq2CkbjKbHHNnhUD4AnCFvSylh1u2e6vJSDIT3a1dVi
pVpKV0nQ3jpHPGKErs0PvplSXDe5Y0NdExDqe6Mldnm1HNYNkjM7kCmJOU92
PHK2uxaFick8LK+peqm/FdUYM8J1N1zhi/gI64D/8eHhSImkGqwdhKu4/NcF
z3rUnEIRXSCukMOTM4g245i8Gxna/wERyBIsgGU2a+I/aZp47Sr8vwCkXZWy
LpUhqaYU8TO5JXfr+ptcB4/p+Gj3ximlVqwe+8VGgBZmSHSdwvCcVhJ6Yb90
LrpeUJe5t9Z7Os/qjkqsxl4niy2f6XMMKzwaHA9Q9uwSHJraPHP2UHgdD+MC
BLh2MU2D0R6j4BrnJK6nhq9nCZmx9ORFbWl6ZGPJequygQOwAhMfy6BGwy5v
rz9+K4MXDJ2KHQa7EFfc6zQDHqO/uF9D8B+g7MrMGfGxF8QxfDa7Tyv7AibZ
QtRA8nnpPlDaMhLA1dloeykAFZtfxLmuOXDKkQZPInChagXxPGjazUoDL4I9
FtLMLOYBTwa6rsRx28CeEP/dTx/r5ENulx8j0hzC1qfAWucVcQ+SATVnaKK9
D8EptJioIfc6Jc9n1/QfgluH+L7N3HplbgBpJfRmWpq+btJX6wcjUNSY/GcM
sKMquVzJ+qA6ccItMcKJEn3I/Af3hv79yFTqIi3qEjXEpkmIhMqsRi1hi2Wm
8MKQaTcr3G+VHAgTD0FIUvfoQiYTP6blcyE6ugM7Rf8p/T8UG0kETe/lIVvp
gai/pjMbf0dEN68ISAUpIw20gzUwRm7ga1uexEjPU0Q7P5ePKgPRySjm6/9T
UI26tt5hKv8PR0PtTpZPjbQ+JwctijCZvJeBF5Mw14LW1ad3plWardCnCI7V
uqNhC7Z9I+sOm505VZ628deTRTe6beziE8IwU6eFOrQA5HIYG16WlVMwsdMN
W5RWJsGPoXaAE4pTX2g2sG53nwZEyWqPTcsaAbsd00qpkEDD00Ucf4YENJrC
TtsbhezYrIIv/1VmC/VTLoq0/GWkKXa1yVtrsL7wFjsnUziKQAYRsNenuPKz
hqR7MzqRHcmxKw1Hk/n8roWTNBIZX1QGA4+jXUTcnw11MhPrZJqeWa8r5kQL
xvhOkl7SyhDaupPrXB+rXdPdd9Lj0sL7MrhVikTfpxKKgrKsZWnIfMFZun8g
Vq1QESCseElceBJDPFhblSfR1KBd88xrPJQyW4prq/Md91osrzFe8V1UQ91e
oXFwS19OiWI8jDhgN7C3JRTRuod0Q6FhEbeNbW0+QqU3+72l82u2VPg7hnfu
4gagolN9gSYJhKKu8EWPlKxiGqt7O7ZYC5IzpHL9pDpWkqDXAQLwTtBsZUK/
Kpcb51uC7bef/nMhgmVzzZiZOU9SDOS4ivQGuH1UNfcxz1L+7Sv0OyhP5Yki
BcJAkwYV+IwaH8I/KzP+lS8++l9KS/u5h438/JcpB/UvQ8b4Nu7ZdLtRZ7Fn
yMdkLp3hG0RY98XBPErtErhrfE+wcQJkClzUeaK54Bgthb2wyYB5i+SuPuwz
1iwpGmv8p4gUR6+9KCGSMPwHooAKYwGr4rIm41N7aYnDAaRM829b4+GHsZa7
vmyQGfK27xeIP4wi0NEMgi+b393W7FLpB1XxhGyQ5WIoIjzuq9tArbaXuHTz
BZ7ez/Caw1W6Jvw8nCDbwudi8alxNKleVXp8E8/23qzODU3dZZS29fRafAbj
jN0gQfJyU/bB1YLu2HRTz/3hQOUGOW+5HONshFyiIz3g2DY5wzYQAth9GcL1
D5kZG7O96B6yH0EpwaZRBxygWrqAjoL/UXQH5y/k/fiaI21pXhYPY6GOiVdr
aG1JB7BxLu/B4/TprHpCwk7ynN9nFm+AWTgpmWHF/3pEd59LOVBLFBNeB6RW
MxeJUNwG4Gpw5JeKqo+CVQIVuZIyD8ZMt33PzQF+gobKAcNUZo5+u6DEcXdJ
mpelG05uAvKzI568tdpSZKNciPkv9ulYs7PoOXxnffR+GS2sw/UwEsIhIxD9
WFUX9heYQ14qn+1UaxbEvw9Zybkoows2REnE3mAGYnkqdiFpYadSUz3vFILT
RE1/hVgvV6OLpGu0MCuAGu5VAqGQUdO3+8RJYoG1EUq+/9Z6M2EKIBgAZKqw
QFgz1pMLElvx6SIPBK/TOLADTd8sIKSmrn3AZ3KGLhVN10qYhs1N1PdrgMTC
fcGe89gGE7VzoBUce7IIDnR4iiU6Dy8JiTeoqw+UOORe7PxuKibA8L5aJ44A
O6nkN6hWPMmVYlYTjQyNjbGMcDiO1PgtIWwdCDrhDpNGtiSqQ7rp8y2WRESv
dWwZAnG1dmhpfEJTS775Z1fKpn7u7XDYA+h58ldSsYCU9yfqEBKdlT2ZN/Ud
NPqGwKA/8E7gjXcgyuFFwG/3R8e4tuT4Tcm7u900YvJt5WE69S0YtIM9TVm1
7J7g+OQnC865d/6i1RSfbD9SbYUb+WhI9S6PgRxByGtRBJ+zqR+HmTxeyfix
osPZs24f9cIzsoQcqEL3LJmOrWFE263hS3KEEvOUcFOQLlOUoMFGQ+Rer11H
zSjuOYUbCyuz9WejmpjosL0wLJbELgYAYsDaupC/agpYNL/bqdemU1qM6mQ+
5uKNiMbNltGqZenXvmJE8y078zniK1nGzgIWou28XvB3p7d9hAOUqYhQQfg0
iuGOGRPhQH+JhdcCtE/G03cJlq+PClfS1tsjUtiWAegyGBjf36GJ6XPkrr4O
vFs6JP95SXrWPlwCauVlbJa05RWFYRUM1lI4V5XkjmzuqJOWOV7yqweOLZNc
G0zqfeOL4KwEC6YxMXpbykUeZgvuxmrYwPBBWM2UFmDMDVEp7847Uvt3pvCl
TNVDgLgrmfOxlV9G5oDmS/Tw4H4g/0l7sMXAz0Hos5kVqsSVBp9bSZaefy15
SOjXdeF7RcfKvJdxEoRCd1/4sDdjZIaKNsvRMXeu12uAQBbMufpea3PZFE78
dNd+yQWSRhX3QkpbmlorKlkZCiWpQSO7fGZXrHFia+yc/a6zOFurhrVaCYSd
vCevt/W9wZB2JkKsscQRa6y36xloBbUWNXpqpU4jEzwtzS4fkFdFNiKvo1B1
JcWI2siezndXs2LMKhWc2UqCpjemdPuf+NskA91d1Rayt3NWKvgisQY8vfv1
Z2EW8nsqRCWcQS36cNEe8M7sGeUgWbXQ4rhqaaippIKqHkLCahFgp9A/jfIY
2PviT85cFEphYmCCvm2MQ671byLRV3RI7mgvca8pdx1jhCnrSSDQbvqU/nds
uZn7UU7MK0AoEUzGXvkQ+2OBhRnDAJXC/L2qfeFeG6sswcTYWiFtM8vroh0b
AEcssi+rKbZCkLQHv96Os9n6JAU1OU3hF+3W9McA1fw//el927Bz4BoMko35
fcranlIhn5Rz802nF0K0WgkU66fWt3IfskV9DrW4ArjxZjWOiboT0RSB6C08
A0VDJzdwSWIypZTJm1Dg7NVmOif6KPJNotDOBoazh1lxAXkPO1/nS30Or1mQ
XVGSUEoI2uTgsTyDspKkrX9fiXS0/3tsWEDY44w30w40RDEO/sX59NyYdhZA
XrIIakLB6lZgidtWZk08iQu5uETHeffAM2kwLhTPPAywQJil7F5bhQXLQ2fn
D6qGkYLNSPTsIdUiO7cSeadaPplq6Pw6xoMT+7IbJ4DywlaL+KjMy1Kij104
n1bHT6cQoE5x5Q1//GwgIJKtjd1HyIzv3lzsq8Cg9M3MVAvRLxTUStPzamZL
JKFMYzX07l7y8ym3PTH64zishsEkxV++6VmWIPl3qW5yjVUZ7fOU6Yz1lSzN
QRZKBy9Ke/KzbnbeY9x4PCjqGOD3bc1KEsPp9BOePyVnoIsF0lMFCXmY9RH2
Z0gkUAN6T90SQyuJwykytLh18g1ocMvocrKJwgF+L+Z4KrdLTIQw8Q0uyaHg
OSycAlTUnIkr/dbCvff3UuJOitdAzxrABx8uE0ddoOkchSK4PwUAz5WYngVm
yhgcq1vIB23G4OYbQGC0jMqAm/ZLnm448iuUhaXGBbr3YL8U7TJ4Tt1rzQQB
+bWYOvfcNEs0C99DnIFZ+yZyiVZOy37K7Ot8w5FhNTnWnsYSacvZx473XpnO
cmBAvbcznkOsAdpzLYouLq8e5v17Oz0kfK9/Xo1G6AAl0THJsU5rVZx6TUtx
TYSYJeJZ3Ym0rBCgR8ylAZ0+vqO7UXwFNIaan9SYkNIBcxhGHw3fB2Orco3p
meXIMRkM2+vK8WuL6kHgZPdbalM/3qdC/Lc+m+sMCORRILpcjs1RyVnyToj2
nOEFprWTGr4/Qye0uU56eBS4Be63/kn+UmzcIkd6vSPJqrT5WFYB+x4Al8mm
69SPh24/48WNERsOGfUY7IvR1WiY0L0n+kkk8QQnNdBLdaU1jWpYVxyj0l/z
kWYnOJ6swweZaEYzVquaNlfuqRx+kb3A3lk59rZ21x3WjK+cK9IFvupRjIUm
6aZw5HhmIWivTk/tBnV09qYo/UQYS1beqVYaiFi0G/CnglPL3mRBO9Qfkn0c
UPkddQpmo4AUXRVUSaD3IB9hXDNoNaBFPm0SK2SOhuDP2CzBG5t6yz43aHPn
IeVe914/AmF1wT7XFo+Sj+AUFcVrKpCxeg1AXxkKkbFZXMqbC8A5YUa52R/B
VblL5TIdLs4fvdLGNHxXpdLAEMrkKXC0m0Q7jSKvACL3NHEPEUlV039P/xK1
7Avg6fIpjwzhKoIwBq/vjyOmUyIcA9NuxffZBnU2xESobj3CsApm9KG9pAkH
s1U2lgq6uKE+ry1RUryiG413P9V43tvhsAfB5DGiUFk7/3DrRNINtBNELuHp
B3ZCwvuSW1EAWBKoldCZfELhJqmWP5a9ISfpTSUF/0zZdAEcHv2wgDJ4nDkU
uCZeEsr8KzzaFT09tKWUwjLFJbP2sPU1y3Hz7aClFycxl77SfCj+MoSnIkWy
BLiSPexwNcu7elKtvJ/At7Ixwvhcg6Qh2rc/T7EPMNqx51NN3bOIXV3/yrPW
5ARLrr6dIuamTnuejSbGv7MNh0Je6q7VGEq9LSRCfJ3gi3RluR5Cn3k7zlBn
1dBlo8uYLOEV+FK1GFA0hksqXj6vHD4FXOCCRaYjivSknM+XpoLzc6F/x6fk
RwpepC8MdysJUF/vT2v2CnLRTl4tcWATddjx2HJuUf5eDaWzPooqo+Wj0YCQ
rlAz8QlrB2hhv7MoLyPyHQHUdl/VIRwoHqMeplFqJ85ujxj3Hd0oZ9yk3Bvx
+Fizrs5PqwvhK+MDptoDShG+y/ZC9eme+gIoqyTTAaYjPY7/j8Q09M8lHRiV
mKQqndIU3dLLVO+03MZPym9RHBHWzmgbeYNbwJh3i92INdNU/esx3nDLqrBf
BF+plPED0EK1EFiDTvp0QPc7N7UC8TJogIfHDGA0Sfn99gJeNhAh4p/MFsNw
J/Z/lhEncVGqdWf5EoBIgsvlnyeM+4w/5OM/HIBTXSa5HdomgXGzMH+fOj31
DlZ4Rrbd4njP2BjCJH/bbL1G6fcgV7CzO14zVLhgTAzgQ8v/AwiC6N3VwalS
GK3DzfZ0l00cz+0VRCiLryessDSwKTcO2vHfY1qObojIPFIF9lwpXvn5MNhJ
4zIEB2xAMSdcRpjQV2XQLqTXByo84fGd5zl3p4AOx0sWsrzSt8yZHMvLvPWI
cb2KLbqzgqJJ+PXF9QzuiIluyzznOvIrkLMQeOscyqnXVyLCJDH3YLwZoSFc
FvgsYy92ObOZkL/sSerJbaugRWCOtminr0jiMk0Mfb3SDVihdPMzZ1Clkhnk
RsoyQizGZtQywEIumi00WQYhIEg9INc+cDfXkXA2CydBWWv9wLhA5w7ZH+0J
SpcUDMqsO6+bC6L/WUWDsaWloI+BTxroUs5dyz4ih+SmRePowCBBrVFo3ifO
Rf3tHQAL3tVF+Ox+Y9eFaT0Ow2Qb9vC5BIyjOfMRP3opHBvV60/0mzQQOR06
NOXjwzifHzDIIha36ggllIOl7NCKdrxFvlo/wXGNsAGXW8HriAxRhm5hZdZo
mSr6I3luK5YdOX2Z8/Nz6JnEVonzKRENNTE80ifxjM63vprO8DwtKwAkAu+g
Mr4bC+KSEcD69NyfpjEXDH+kg3suRVJes611kQnvYbedxyEFn/LddLnZn6Cu
8pd+DA6YvsZ99l2RWK2os2dysOTKxE0ZgcSdsqKJM1myOLSnUsWpHMFid1T2
aajKucYH7bfvLheDVq3q4+JmJQcx6dIJPWn9u2VMkqQmEhcMHGdMay4MpW6t
AFJsAWpNCZAmlHedO17HSQNHE6ZenOhAoyTuzSNVBGhHFgOP3kbeydrzr9m/
seRMN9zn/MRyHw/cdbkmgwMA516GIfGcYR9cKLdIxt6GCs9wLLgzjEpNLx5h
fz2WVIzOhUQHT5Z6Dm9xYXyhbwWf+/Pjid8YvxS9ozwka6lMa5f6ZOo8LarR
xO1b04Qg4Cs/b1eb43UvHqNV68CGhTIiaOH5aW9X+WvOQSuAcBnX63tvEu6A
nfHXXTsQQxLup4RiSfhBLgYZO+3/ctUWCWtwwT5V3eBgQjamoP+op4kheOqa
KkLM3uWI8MXnv28lYuAtQPIlYjyYxGma79vlMILtWJR8I0+OoU9AlYDEud8x
vTaBy67tNveSiYMVFQzC/esDnYn1vdrTYtwzMNyzp1ImAMzDCTc68snHAGCe
bwRdbm8ASQ+Tg+kTR01BTXYmsriwbRSbpZaFa9NeQMuoHBss7MBbprJUC63b
UNiO0DtnJqgAvX0ZxnfIO1vHJSGhwc+4LBxj87NAt2w8hRKtoV/oZ6P6mXIM
KaGFFQEVCs6PhlJxvpLMdpR9rYXJjFPhR0lachnldGWbq+qkz/e51kLY//xd
u4aIhIoX1fxQSmSFbpcN1iZB7NRDOpjTMr5/17WgLnecC8ROgESVDNaSFBr9
X3xx2+u4YbNHaz50bq2pbVVYiWttEBBkZkSjbScPDs9rnun3jpYg61k3JjwQ
IJwmC6AthyUgGTKWQTONCk/Dx6RsvLyYiIXp/rfONuWS8/yqnfi7mtzI5rV/
lZ03/4xZba0B8c5nazCOm8ZsD0t9MXVMfKhxj+k7Hm5DpxZ8oyfE9bF9kMnh
sCJy2Tp/W4VMgZwWAXRRmFvd9P3+geN52Q7A5f75piSOSP+6WvPBxu/+icxy
4ZJgiewbD9U7dW+Bv1GQmQme3ouwSLe/CqPHqEXHOSpcqsA1zJ7MFBsbGAz0
/5WDG0S/c2Goun3R+UoEVNgdtXFkNlFfcstbDPyjJ90/fKkYXzGXYZpIdLsW
OYCy45lg2r7Tub/8ZROaIrL1UdDqIih94uxPCbsb0IhpNToKiEpLEfW2zhjG
zP9YQnXnHLTn56WqDDTVIuHcwIXqua7mRniKkR1CbSOcbmukh60BXTyN4kJt
yPkPfIftmFQ3sGlamzv5fiqjQrgUXDsTwdoMq1t95Wb5IcdXXxBMNgohB5jE
nercOfWIYchPy1vzJVD6pXj23U+j7LA8vhC9fRP+fRl/9iiWR5F5PtumYHh1
fUDKA2BQ+Ns5ArgQowypY7fFEuWvtMD4FeeVICeSDjAGp1FmbOGKrh6iDuXa
GI5aeB2R8L7I7zVT+oVoG5tfww91fbP56tpPtrpaKBeyxI95hlUI54fH71bz
CsVE/YvrchQ8BJ3M4EXnEqjXSc3wJYm1ydSXOeZi87KUQnMnNZvJdajQbeK0
67Hlo8Wym737IigVTQ3VbBegvhmKbMAhr2zSBE+2Il89gVGPqipxPuI6ECBD
t+b0twv7+B4KGkNBbS/4dr+Rn1mnZATp+aZQWNp7p51rFF0CaaPZPiF0RfAn
r0pWRa9g2BxHLlvZw+UYRJGv33dyvasVA4Q5F3HZ0rxyEBsGScSxsHku3noj
ip1kSV+Af25sWms6xsr5cGlTzxJxZf5Crm29HPnhXiHDsoaOug/Yfb15ct49
H19xGyUM3VbDGrGBBDIAOOYNUN1OPE8+QsRq5LzqEVJCu1F90BF4PIWBur5G
7+qeePkS4pEmJnXIgqzX9AOAYBqLVwfGIYSgE8f103TZrbQFrXjcbHg9lW+7
B/j8X2RvvqQIdaPhCygtUZeN3ZfeF1H2QyXNFJpxUtGux/3+uQUPPF3eS0Qk
Zs8Y9VW2ClJImFg3Xx+G0IXIq1o9Z+C0By6SraEzQYBrMbicpurlxGQ1Hlsd
xz9FEjzAmGsWQ7IRxkEt363+GZ5NyJ1Lv4161t5bhkhkFP+OHls0l3q6QNBV
dPAbuYG4xbVAdGR0I7VvwIe0u3hChvfz10xA0b8Xm33lHe3XwZrx4+lzqwCb
fdb+qmhB5i8mkXPtL9QLUaMsjDQWtOwjTgYMd6LiPvN5Ja8Z0dEc3EC1x28s
jUB6SHcCyFP3b22cqG0o63/DVfufWypy+9qxHVAnGQsAjsmVP7ytebXYzHqN
j9J8rg7pNK15ZVV9mmPy8SBJaQQBPx0OXGbnXyhEbNfG14218xar4Zoj1Bvo
qnYasA714Jhalu7yaEEdQJSayXgWBIhk3mixqPc9St43gmBRZdRNDiP7/QLo
UvclYvM1o+cppGl1gQYLe4HOCucM8zY+SY2c9XNb7CRmixpl/FvDoe8fdboC
bK8V+zZYR1oa00sM9ilKqvzGnNkTsyUwUn66RhLGZu9gY9zKbKFlKKFCa5b9
nW4d/2Vj4q5QXRPiPsyI7H/toZBuqqaXX0VAPFKZ2AXe5FlFkCk1/sL74Apt
CwXPGJt9ZNm0hsDlz1rp7czowEaqjxFv3m3DOeAA0BOzbLahI0Wtc85DUUNT
L7BNVZgngeR9OP6OfJ9it4wHa4A13+mY/KofonivtFi49PC9lCxriT8fWknV
cn6GVj4+pJodMrnEt+vdrt4EBjwW49Pze0KS6aMiayB2w6Th/LE0CHdS3Zn1
/6cbeVjCzTEbnso05+Ten5dCGW6koLIHk5Yztot6GWMFJAyWUIgV2BHUR+CD
FL+PsDZpgEy6maj6+EguqQWygbjmWTBF+WOmZwo1PZzWioUz5bE7TGxEPMgO
GJCRyWKr4v0hGmPx5cZ/8PtCLcnpc2eCbVd/p65RM/POMZduAPxv4vbVMBdi
0hEvBVxLxwIpTT/i+mGERh00mouHWyo5IH6v743um819O6zjxd0lusbI/sqE
qdGSVWRdAzDB3DgT1KTKa6eZzdb/ZfixIdLiJZc7CJ+f8z/YIuSaJTdMZGAb
JAeZwaPqDCnwIzcqgdbsKYmd0B24+U+40/WKyLeT+T6xvnhkDF9V56I7XpAA
0+z8ucCSWCcswb01WkIiJbZ5VES/SXW6Mt+SNsj5WmXRPrLfzjmqyIhm7ugm
y9yldzD3lf6YufSKe/glMm5ZHrcQAFVSKWylxEwWUZSE0rigxAWJYh3W9eQ+
Wa/JWHMW1XYa1nWksOgWyWYpix5tOc2hLOaclKwbmyN3W2I6/muMQiggoIiD
4fatcT7yaHWLpERzStmA2feM6skAHatdtQdSEm1ZmHTLjKvcHpOS7vtdaNAP
n9dPuqzv3HdNvh7x+XTJ7p3/3ZCSUoHLLJ3LUQVAJ2vdW44j+mBQ9BY2hsmy
0gCsfXnu2AcqyJoJ/D2V6ucSNxa78WxmMYJhC7/TrBg9TIoAvuVzuIBidoJ+
zQtr4BsSE6jn9fouDAD9fLBPndtutjimHcEhwbyL1B7q3NwTAaVqwcyKFxco
For6LZDWn6PoI310fX10ezTGP+L+D8nYwpAH2jE3SdD9wNvy6eIouIAKiaCr
HH31dOvjXjgZNR/Fy2FD27w5rIL4sfwlh8eIcgcM45EPJmzpYTSIr8zZ9j1Q
Gc3HanusQIJsmSHFogooIkA6Oikss8QVyfPOAs1zHJlT6Ax0ffo+6GJG/2lF
qlR5MlvUOkqelKtIPB1teU+slkxNTDjhkByeYcs5P4vR3vXXXcVcroO35clb
9pvCo10sg+2v1Ah42esvweuaAUh9qUZ5iaYsmxySQjqDV7gyYQZ7OVL1tY8a
YyM3aOyV569CfeS8cN59Ext5X78RlXWqRA1SJzWWhAnhZqYgUYy97umDjlvr
O7bnJ8xFz5UAmSc6CSo3nUbf6SrCYv3DcgRMi5QabcqNQ66D83J/w+ocXkDk
o3sWjgCLFKrd3tbooF/ONgcbdaJTj+f9Z2lTb/ftiRsYtYZHCVHyES158EyN
1b8AkDwtw8SF8FsDfWome9gsTl/dAv+biQcbbFGyqgm2sJV2YR6bcBn9wXjy
Gliow8nWc2OnsBVoD+6ogrCpsFX33AalJKMP0STs96dsy0fbIlfoiUhqY+Lo
GYHXKF4xMbYhAgjrHVJoQ8jL8af1RlAs0N2rdp1TTfQidecXeHRjXDr9aVee
WcFQXiH6poGlYDmGnttJ8RO+1+GD2CoJD99xdvbfjkEc2B9SRHd+kqyDhNda
xxYEHTsD83WWb9+xXHFYKzwk+aAETDc0/1jIc6l7und7EBk7rtHc8Moz5xGN
lb5+Y5pKXF2dDzoeYVvYOFAY5zzT8/jWTPE09sep2PuqCbHUw5vil1MvQnOR
PjHkiztxQJQ+DuQeUn2RujvHG4zkrN+nRZFgt/DBwDZg8jyy1+WpSeFBeQj4
cQKZJekRaCSOcKnrve1AV3zVg/80shFHS/wWV6nzlcRTiizYWNxANHqeR5j4
Syi4JnAjMWrB+XqcCwT+YHeGBKkdnGCqJ69zzft6eieGkFY5zFa0k0KQA093
20fSHX8cSGDT20JEnoiv092ofWTvXjAXg7VMh12Ylsq/yV+V0NbTV8Cz/q4Q
3e848VeYvpFNu8o1/XEaWRNpxP5p7dD4b3Rq/36uQHrloocTNUhXiE1rpoPn
2S+rezIv7L0urPq+C05JAIAR/YbOPPzKIwmeUINKSBepR8fnsgpIOSBjpXGa
BxfRJjdDcIpIfq4sRO2I3FjTNltzJQuC/B1iQr1mXRVo03RopLthK0cm1MQ/
OrZqUBlLSYdVCm5tvGCR/Eu8RElMp5/jkfIC85kIeI2aw4iZ6mQNC2z2svEI
NJmxD+46MvUt8w2vJYKQHkTS/stH1yo66AvDFTCsSCzGWw5Az4OlJZEDgJBU
IL+dI5gdRgCfcXmtgdt7k1NsCT211EHU8q4djSC4aSGmNkyiZlrXI3uN2cc5
3Hd7mEq8LG6upxiuMuqdtdGc8FAhnKEv1fp5EqBQZ4DpH7jzBwrpojmS3/UK
XNNZI3myQl4TzKwR8xqaq1+8ZwhDHLCKs6wfpKqcVSUSMQfYvsbwdUf8LN7j
HygoutELsTd6FsEeXjF91LbvUdVfgt9QBeODAxbRV9SnC0GIulD6odg6nDeP
gy3aEof8ed+IgiqpkImiWQFQXSLXp1cGOhChEQioClheCuL4ftyE6bMsDTrn
WgAVKA1sWh52yEjyCBhgDNTf7hEnBj6HZP8XjVdmO6jyjkHqLxYpZw7CGT1t
OZXxAEPpJXaCt05dKULAVfr9CKh0MghAhwZVWT8nhnBifVVok0bO/XjcyLnv
Zs7lTUpuWdkXvMjBXDY/tE/9QWid0WmO6zcmXAxwe2q/fVqjG9ZJQV8xJ/dr
R7RPq42aPDm4RfXblLtvab97oNU64Us0HHrj6Z938U9ucLMr07VfBmzyG+5k
BYBLBhrEQsbiMnJSeJjCCbueOOGZj2VxKPhqyNsfaDQEVVCOt46jwSuyOj6R
rvs1HgEVo/xgZqp2Lio5F//gb4JAas4w1d1C4LC9SuXuWil0668E44Rf8eLf
Ke4YuO4rcm0xuTB3HY7vVw08hPnI+t24RjvpEV56Z46TRzPHhiWa4quy+YLU
UVXO2UnL6fz37c9e0VJlgipGv1+CYhhO25pf1ztwNbrMKYnE1XqXMtyFuDCJ
nnzzQk6qMHGjI0VE1Rz+xckR9jdqVOSin/1QjKrnzKya1FEabbrea4TUVaRz
g3Gf0ziNkZHXmVyPI0CcHnuOqkiztEtGiCRcmgEMjH/8FakZZBDCfRM9zEo5
YIDpMd2qsXxU2Nzc5Ow/H5AOuRxEpJYFs1XKT8RKeNabb93tKY7HEfahLHTG
ir0a+jlJobNp4i7xovmeJ6xAiDtUp+OgjCmuKwfS54vofLErg8FdlRlkP+Vg
nno20OqSM/mSEKYcohRB55QdevZ+G0acAx8oJq/32fNWRaZ054sAMUWUeS+F
3uajwwLMSIAT6oQlA8sJVI36l0LdtWXmfh9ukAWMeTQMiuUQ3BGQO++tr9ZE
VxO6wddg7mh7uY0rhrB3mWR0TRow2gl5ER3J2JOr1qlVOSE6GSVwtnBTfgsy
6xet+1JiCJ8T/b4K5NXqLJw3eLLhq21kc635zy9hysEAhUtMrZEviixrdpJR
H2KT4qW52GQ5NKBgGPQicoosmNpWQRZfFcmE8yIgguIJU4tEoiOmVlDOv7Qq
mHUGz0S4wPt7/yrhMcuMQel2TsO5vQYa/lclX5z0O88W3FdNDRKeDjw43/br
nuETWht93rI+1xibRRnzM11IBCGtF4iSJ71SbO2TqK1VpFnolYptM/JASOwT
GmO09nuMovWinFBTLFXbhfxENO6Mvek7G1VU2p8evh+WCxE3BxoCYDuc/Pav
sNVT2g0kTZip2UkviBxfljW5JqaI5jo3FDG5EGCidPS6BJh9NJF9AW5Y7HTp
FP627Ai9yWs5X2CfQt3noxt9meWrl+E6vW9sRNZU3SmiafpNT/fWXUMp1L6Z
rYZuegGsj3uAi/o87QXdQ2FjjE2NRTMNX3ArAqlTsG4mp+6bu/Qa49a/y/1l
4RFBD7jhZMyXpCYi1WE3X6Vu6p22bD0SRSdfAEdn9heDcTD9njmrkNc3e+iM
34fcI94xPcMKzYcR8dgvGhbgu9cHn7fncf7pBA+7CYxjuqs7V5NDIQMyFAUB
AASoruRPqrX+oM2wZoNgTqTNF7ZEwv4Up6lS8Y1ejEHNRmvpTsKTCemxmPQR
73DPi9lFQ+lmEYXI4RBS9790yWH7tqpS+W6rnoLz6l/Ueeup8zqB0kCUF/zb
wgpff91ElHBo9E0q3nWuIWPwp/Qqf/09zB/SFA3iMNlw3n0EneiWprnBnLHg
RXTlEysW4HUAR4xhyazhfgFLpyaNy8iS8j6zSyWMhKkjZtAWL09WegSC+KGQ
JalqyOLSbldp7eaZd5TZj3+NwO4J79hFZWAJA6A79gMcN0r2eZZvt5qehe66
ZR9FSmov144qqZfmiMGE488+UsWw8QgjxceczG6KVAEVqVUj+AGO++071o7g
9t/76mqk1WvjS5LUGMOFpCxvOVWRKMsLIP5qqGj+VpOqWkdrEeeBaccI8SxT
rTX0F6rv6NkmID+Yqx7n1sih9yq/P3YP+DWCqD4MRBFV1VZh2LpDwaIGkEzZ
8pZdCulVnQsutByYty2XtUziWyohnqPIQuCdSTJFSLtxmd+4/k7FTHEdgBN/
kgj5dDFvCLvmUL5q85xPpV0uue4D4lE+lLHt0TxGat8A2nxpoRI4/eK/JbI7
greqF563yzskEgB/118kKrvDZ/4t/kfHSFSQ2qIss1NonKRJNBBzYZVJ7JWx
U34TsZw+9zVcYgiAKiiXGETy2ex0zFgLxsFDn3rrkzy5rbKzKpqnxnFjhtIs
khv7SBPMW6zfU7YBl8zTue9hUF2t0qr1njLBDd9DTMa4U0k7FHaIw4U5189C
5g6oO43VRAtkbQI1Qqwht8tbZZjZx4QzR4S63FA9fKIuEcG50CP8kbDwQ47J
nEkxcwcfXEd74TPW3tEhqK8ayIiGL6KOW+e1v/7VrRpjmNKjQLcGnC3oXDIx
gV2MOgJOMVu9NH5dgT49OxXVYs5HpHK36oHQgeTjXyO6X4ACDIXyNQiNFF0D
MaoGSZLs8LN5Pu8jsqcBPrrOnwN/QG3jqXjguTCoWb0G4NR1NlRvGNrq7Ccu
NNJTgbLbf8CAZTLYIEHIBhctG5FYAGRyldhQ3fqGqYki/NJb+KcsybKpkA2r
2yTGghPVVCRCaZKKQpjXVz6xuWupRnC+Ju+Yg9IvpktBdMOLiuGrF1+OZC7W
pDyL+ggSC+m3fNwYANsc3459mTKEEu0wKSHwfnglz6zaE+TZk1KgSr5ygUVf
xQeTYQ3+Xj+Q14UKfgF08eWVdMkeel9MlCCRmB3CMjpX+C6h0ojCgjGWCGIA
Ssm55eCjbv4FhIaOATVwaJAl/A6mRoWTfUdBpqxHDNfYLifxi43byGV2T/LY
x9iiUbvKlzxeqsvOCoo96oTERM12BI4iuxeNhIg2R0CcBIspLlGNKGS+42e6
0FrdyHidzF7adL5aP6WDFwzC+hDEQhAfMO8n6rZsmWlOIRRMbrC5WU1P1Y2c
34wnDCLXrBzu9gGm0LCbWmIIhy6oV2pt6XYOElAJbHQ4VYd7DkPPm/Tgo7R4
tY4zpqU0awIgb9UWf2WRQ7uaQ57Gs8OjFCPLbET02sdHmSrv712eaFNJKLPu
Sr8g7HoxFQrqICDUWc3ZaGymJmYJzFykrXRJQBd3IVkTz445Owo/+lqUX4w+
SuQe6lpzEJc/ViPQC+iTelclAO8XlHhG/P2AIazboeQiP2V9CVdpIhxEQuHC
epZtceSKQlFcMJV5WKHwPlEwxVOqZk/E1lab9KEDYNhEo27iPd2UeSBrefme
mHOx9YBsWh7UGB20K5oPHIxuc4jN9c5dmuHUm8Z0pO/Y36zBa7TXs/wrghNu
3HOAIWzqA+z4AWNeGvsJt/A1q37zS2q7e+RUTpMftGmtKzhE/yfXwRizvmYJ
9ZaAxIVtKDckJsKvOkAbuiTbEWY/9SHuBsPbbzV/xTbF/SetQUSex0tKNbkZ
NmLrXnt96HlhKVOmCehBCm8xnwcP9V1FDMZfrCnmJE/b8bd/olJI6K99rCps
eMBdbR+bMDLKo2+dj8lqGW2MTZs36JqxqrggGFvHjeucZzNiOvRzrs8rcAza
WVevwfYrAUIcw1qjOm/yalA++MFTPYgQv3VEFtLg6RDhWmbGo1ZhtPQB8P1u
jj+0um7gHxMnziVxh1FpC93WGrjzb8miyHrsTu7xPzTJVyJ43xcvpP1JhLfl
ZxEdk4o5AhTI/ecVBDo4u67qDLfOAwXKqyve0QSSSaH2qjX4Lg88prxnrMts
g47+1ynXCl6YV+otC9pXSdlZ2VuzboExCPTprHO0p7V5z+IVJ0nWyZ7Qam+8
3Yz080+yFg1saiQ36wKR8y7RZE04C3CoNWBccShJN3NPnjlfIXXfW72C3VMw
lno78TbHwrxNjr52VQN8EP38eVDL6KHsC4T3tUhMHs91uIe/WWi7IpH13uiw
oROZzrAxE/mB57XaLHwM4ZGP1t7mYzpoHDpp4CnZpcw4QzeJZbZMVvgQRZrI
A+QjlFnDtj5v8mgnCJx+OAmQz3VA28Ld0Rv+YkOeXeQQ9TzFsFESKui4TAhc
+oix4OGSDSO+4KOTF4H0T6bAWGJUvnRU/VqM9ZJKCzSCh22aKZZcDMktR5FM
+vccu+PBkUgfpLb5bYzCE3dvJLf0O5PHvfOgFZV2H0pKjlKN3GFEdnT5Apub
TZFwgPWMb1GO/ZNNZAKFLDMNgeOQP+Iq3G7SHYjdto65ubQizArwlMHoaVja
NDDJ+VoWU7eChUjsFHokbCRvN20cq0oyQLETMmI+cFBeVCQH4b0N8yUIEstu
m1jxhs1pQJ8WnqBaFzinqkt/7ICJpsKrcEjh7NzMd4RATV0lkJBz7OmffIwM
T2icti3bf+wCn7Ylgw3109MCvABTJRLpO1M/DbJL1/lnZLKBH9KcuLz96Sxl
veYZHd2qJOzm749eaOZQPV5+YaCj/38yJBVq0SyX9k0VGojHjP01cewKebOI
AEuI6mwo3wOtcKl0+2Jkk/oxa3XVWUJpcvuQy00H8MKsKH2y93lft2jn1MQs
yrmItMQeOOdBCvg3C6Wyi1swiKN5DnQm2Qvh7ikqtOjdGkNUXpccC7JbkUr6
p/6RFn0Nc41MV6AQgDucPX48uou/tnGKH9Ao6tDrAR/IJs6IqgkgaXEdMS/y
WnT2I0w8fkPfvwDmTwAlQ8eRUJQOnS2xeK3b8FD0tXmBMDlrh7EI09KvutWi
TwsAf9Hl4Gt9t4/5l5FOSEHt+GYshjI0vaZbDNwqBsL6jjQxq2s4ws85j3w/
DH39oBdKAsmMHkBjvoDi+kKHMf9iwB6BT65gJgtxRbjCIpjIRn2JFWSQWwYX
hVmiQtqsu6Crn63p+XfHs7xDg37NTLur8JrcFjGm4Vm+VbYXrhirAv6DLaX/
nKpcohGqpmGURtNkyRdN8x6On8s2mQLp/URus/kgMFLwQ/Q8HUVKmX4Lbdt8
vUQ9JkO9quSMCLwMqugDK+K4Fn0x8Wuxbw7tUPIdTV0R3y27bYGf/097YoGn
gOd0Of1Dmf2NhOkK6FG06GbsFoaudHd1/3FrhfBdvHOXODfkSsKniKDnh6XM
FGP5XnIaP/D+9bQDQkY0bnD+6rpc3nr7+g9PH9p/zthNOU0YWHilSQUuJgxN
9GQEwcQWXKti38dhHjuWT0TKCN99Mk3OkDQtKVV6ODkNkXdS1mpwvr66BXl8
20b3f3IGEUQ6GiX8NHXqRs8Ju4XG0cl2JYETSRyl1kTEOZKwNuJp+sxvmsNM
xgcXFUpBK8W0NchaAEnJlWFtOBF0CFuAw9QDFiLFxoHFnUnPTXJLnP0L0+vA
wFVWfVryXcUb31/6auv93v76D1Bn687xtsNJCMqix3P9C2Qakacwm9as2QVx
GGRiCY/g5LWt7tlkK513oPElC51haSnkCeZxoiHiEPmb8x48+bj5uI6ecpaE
DQZIAvSwke1u26Zb/UpZWTEWJhXlosC/D03DTx4xyRcOfSXj3LKE/+gg5vsN
XSLx4TyXc48hI0S4F28YQ8RAVBvlbyesAyslskggb8zrKR1xcT6NradEBn74
Dp77l1pTWiTGO/ELgQNvilVRwGCn/1yarHsZKz1mr7OAG3fe9ctjVCg33Q/n
Wxh4eLK968U0rNaUSBGbil9k1lORnkCNDBNljPERhmapRBJ5KqDlGfGMUEmu
wO+DJfsYzB+jH1/bJwQa4hXsRyP8DRvIGKmleM+MAJoUvCld6vjz8TDsCjge
fi6NfQ3jmeZ26JmxxqoRUHoyNuzK7f7fqdfuiMa28EJSXzyfYIXH9IMO8gY3
Mtn3W7JmAEf7jxlD7B6yaWeJa0/mnn0HPvnet11lo/e/ugvshXHDf6yEQ6ui
/gRER7wQr10nHugep9jm3rHLtEX6bQmEwb76QskOr9T5l04ZXlerWrazszww
wOvlmg9tzJeVcL9vwQfIof2SEqI+gQUPTwGZMH+jKSvLxmhi8esqdwXPbY+X
lSsnTwtGsxhxObFLXtl9qk7AfQJdgga0HViz6QsqIdAyMsVh5a+jcrGe2o3F
OElLXQfGuk8hCDOpWuhrr5LEj7Z8sv/kSO128SnfK6pwkEWUYU9zx44Gb4IS
NN1uoepTmhjHnmEPU8MU5zbeTtUvVJJ084Wy01nMqmyHWjxudqrhzx/+0Apo
AHEpbxw1XPo6dMRqCOuHlqPO4OoLF4l1TF8gpacRqwPy1ZeptaABG5f6ZEvu
5VTHf6vCNVPtUWuGx7vgLN6fZVxqtkRKceUhwB4tdmixO1i7o799OHnaX6Es
FgHS4FLMvQPIHdAnuFZKcPBM46HbHKWigMwpmsaQmKhKQY82rNfz2xedlwsp
cfgTkweyVq/IOgqH03ZUWcJMKqqPnTL6w/RYScveP7W2Jv0UCoRbAkAh54AD
+MrteAYXldryR8hgERclWqxekhKrXj8fjaWpcoKfz0ozw//9s2xRoInzOvRT
czfyS9eRxd8PlMxNZyaC9o90CpaNapW80ri7dHEGkGobADLz8gv5OUxA00Bb
C3YO4/2SecrOAs5X7fXEp2CLFtQwcCUqpoGCKka0fbx9CP+f958cU8Yyjd7G
KiFFIh2zhsnTfvCeOPy9PYORhNnD6jVRNV5CkEeddMIC1/EvISam1cQ0OK0L
jdgpW5ZJIVWblhQVkLuKbgTDtqM5XofzYiEPAGmt5ZNgqnGj1gVkJen5a+rI
helYZVexXZK3P0rOj0+pMMDVF67DlibSgm/kUV/shelQKeAk45XwoVFt2xhK
pnOPxTBJY5B/0q+Rlj/0H8o/dwg/OC3LCXsFldhY46JbAc1bGbKjQ7cu8WnJ
nirZ1t5Kq99Fgc7YU7VNQxKhJ4mgZEvElKCiE/IcNfhHBpqjQ7YDL08dYHsa
mVo7aEh2INN8R/Qojco8P2jvF2HX4yLv3RZ1fIlxrc+Jh9BJxYZ76I/8b+Qz
uHQRmtsDL42NUEE7kJHSUZNkshE2lV85qosAhhbAAAmgAemM3FdwmXHTyypB
N4ZxoruOh9Kx8iqw+SYO1dvYG6ZbVgrY7N/HF3x1GThCBkB8xfrIOGGbEE2U
BuwglsK30/C1S6NE4NRG5NBq5ClGDBdvjzh4WwLIMbZFTRcldKF5mlcE9Wra
1yX87rqRcC+6KuXy/bl9tnhFvdF7um5bYaoejfA8DRFaXaXHHD/8+2Mq+nTo
HG42K6hsqwTcT6C21Rlid1uLBS3jVlq2Ni5wzn4CQybC71MefocChokLYrPI
dy6DI7T9T5wqG4c0Z8NqInyd4f8HIsj9y77KRXyDpUSBdUO9+skZYBqEFH6/
YJbyJqzoVuL2kIp/XSzIf8EvdxGPZWpZwzwZxUoa7xeCIGGZ7vYw8lygfcfm
mJns64/R6Vc5k5eY3HvvDwO/h8TZAih89DTZbJNepgiN/Kgo6oJLu3/28Fva
NTrsWG9Kmm+SBVRa6yLGJhx+4Zgv2zg5OfoDiAd+mH1tA+OFv5QR4bf+k23C
Rn1ZuyWbiz0Jqtll/VP0RHVQgL48E+i4dnBwmIQmFCIUFe7NvbZx6pGPrESX
CAw4kfdkwjBqzxkdDLs8zZTQB//TD+l70fDVI0NtSmwEgIeRmSIL0/19WKGg
03EAuohIh6ByfMwnkUYZhubT2rzB9XQhds9GBZyi1gz187+yTiT+B//+MORy
2Ls5ITUkzhC8Z1WgyYaK16H/8DqFV9GmrNfJgpvg6g7FEy/cn1Em+/Vn6abJ
IfY+DcXLZpO72ZUOUubZvhzzhGYbhBvU5ljlq2tvE0Zmh04hGCjsxvfTieXY
Vw5RXEq9Nda8bzzHa3dUDYG1UJEMLR2yYQefO0N2sg3hDLdHcqBqUNixpD2K
5dUyPgkOEt53LmobOEK0bIRakc6lhqUvEsHFKTV1UIfv8Dx2fBQyhBbU0rCe
bcYVnR31XYLFz9Eqx9ZHO3a+b+0IkltLEoDIH1SWy6HSAoyIat0h/7m6zw83
KDm/9fBRSk0yDv7mPUtOMivdvlihz7vE0ckdpXN7XRFBsiRt2/JxIIsq3uhQ
H5ehOEQWSMNF0bJ/M/ScDkEwqyQGiP5Nupw5INXr0YWI9fM98MQc3A7QF9CL
C5oD1yUxCAhr2EHBFJcJTc6jWp8cU6smdn5BAzHocxUs+vAkJBEtZHI01y6j
m1iNKHnJLG6h5EJXAlArEXB6sQpGtwrU1l9LYVBA5qem6SWdtYejJpEi5UOA
sOj+IEAOqcZlpisd+KzoplfpJ377gK5yQzGCAJXmY162NciOpsvGLaw5M+U8
3OKblmGlM8Eoz47iYmlXDbJbU1+mGv7xDgjVUzjX6KUvaxRf4VvtQYlpEUEP
+3LtVof4GeK/kkuIm6ync57hsu+Xge+BYjxsbRogiPlEkdZ/KFfcOFnYVgpV
khjzR+BIkXpVDFaY3uCVSjjsAvC2nm0KYxb8Za5qxHsTyIT5L/pZ6vITtgho
QgZQTW1Ufcxqu6GpLgQ/C9seW1jg2B7llFKoMhA7tRPqL9u9GpJTeSB4c+qd
M/kVppfo9Mt5mnkGQYjxbiPq/gfXApOmMwZrIBx+ET/a33MWYGnsyoOPxHSx
v6wrjxBuzCzeRJFDvECSEb0KrwY/pQxQU88zbN24YTsAy3RjZdhb4OOqOzZl
pzhKoW+HrHntLNGrcM4m74IMPNokfKAbAra8CtSqzEL0nkuC3DplrPvtvoti
LWKWYdXrE9RGF8fJk2ekvuTZWO/zmq9HOl7j7byaEfQQktDi1cK7UdKK/lDO
TwV85iSSAbz7R9qwhpEdpgNdqyLpWyRbdfMwDjPTMCtuuY4riRyhpTj7P7XJ
lfh+x7GHLZ1LMb++t1WI0IPlHRcUx9WJYQrvttYfx9/1Y8I4nm0OQ6LyOOSD
8lFcm1KU4+grajWbGH5YiUWtWaiu4mVs+QgxddzrjveAJ/ZcFsfPn/Eln5xy
43/NEEHsxHFjLy43M1saLkrfxz+Uu0Ad00r6AZaKi18KnrahKcYgGpcQV8Zt
QV7tJBeH3Bjdi2HlzJrwMalLsZQ5b/R4xFwH78SDyo898RPcPNWmY1ucKW9a
3lMx4hBIpFPFYsIarBclZLod414hOtK2d0/3ay5aIrCGm+YnjQTm4egPx120
fHkABM4eq9pzgFcCXTCExuWUq7WX18T2t/ScqpDtsyJ/EWDNgCoqDRUNxMF3
ZQg0GKjhDmkCa+N4XJmt5CGpgPrnQpqcmaBxTHA+Q7J9+zBVJ3Ac/lmD+yPI
PGXzicSylEtHa/uoKf5W0hrjvU0xs75cKOFpsmw4c9gyjHfPkpHUMCnYTU7X
KHiZeSoktAT6RAGWC905BpvwI0PYqu3g0VMb5obUWwTq9xHvw7yrK6F9z3a5
RC962saqurxefFgcwLCUikQ9Ev8LSgMTdIQTDZAcknqE6ssCuBGOjGeQafCJ
2UAV6LaNrc3XCOTdQXyr3x2c0rRCxnHXoemFBr1MWbdc+XqE/r7jkCczQmwI
Cyc3BHY+YhS/a51PAllEA4qbDnWfWudvhvf1aOFTvLY5jb1SROZFlBD6XSax
Mfamhx0qjHvffR+vAGqjFz5MRsZTbRnOIwEVVRVqnWARLz6iNzn16vUp0BSJ
5amD7sZFtvSC5rWOiugXaLkSCh4/Q2dgrnE+3y+tlNGRN1dKKN0+nNr16jAd
CKy6tr85WGBMga90Ba7T0UuhDBbapHpRbcMGE5LaKPHWOPi+ta05ZnOrZ0tP
hg3oVjQXqbahC6CqSAEkxtN+xRy8dKKijCpuZv0gKIXkSUdUD3NyNztE3bNM
WdJo7HO+hq+1ABn0u8AmlrHncpK4rX/WbfICus5VW8zCJZDdq6eXRYuNogd5
/GuCDiIxRa7ChQxOFQpCOay1gaPlczjZRujGPDmAMWfKcEgG2kEQqX/4jM6e
o0y+HJsOoNuOEiCBPEi8cBZCfkPY0IP18DA5kvXQJ4eZc8fsDQIO8jOcAhH+
mpOXS94BtyX8X1kVGKWeuhGC7NLQs17qq02sCdOQTo5WhMtRT0zvrpoAMu+M
5zTKgZmFupfWl68v+1YBYd7Sp3j1GxJhLHRtIAjAhhdEUoZgw/d/os5eITBk
Y5/t/4XasSAlFmyiorryKvvZtW4bAfB9im9nYu03sNR+Be2jaajpM09Cpa91
gBhwY/JOnE2XkQ3HkeVdAmA+kYnguhkyhmngUvE7xXtZ1LmNclmA44MSFuOW
WYSIIe7wLMeRqqQTfyZMVIySzSIcgVanvLMg4iSghlk2MlkfIvMJN/oKYYqJ
SNgUr91E96Q1kJ+Pn3KVH1M3AZnpX6kuIhCAQut/MQZ/sa9TB/OvwpuggxpU
hWdg57LKDHRKv230rmILvreZhIb1/a1wY9lTYUXv83atQsa2/ZAv2LVNLtq4
+fdoGsumQTsa4r6Z9i6/wrwT0iHwAQs00vxIqjvo4Kcn5vmNvzSDXRUIpWU7
SzyqXFnC2BBgz5M3gyrL5CI3YEP4rtIPQhuKHwwry0ZI+tb9Yml8Yr8SOna5
mnJVJeLbdFbIxbr8FQxCLQJAK39wJ52srOsTJ8kQO+kxjdO58OADc5S9j4zL
4H+HZXUpaGy5SWPd56oiCKlHdetYxQrk6z6u/KLBTDHtv2Pc6GkxLKZRDHha
9JfGnGNoiifRK6SJXb0uMcwu4GQRBaA0QOZ8cohjzHfU22cJSHqnT7xMT+k1
Xrl/nCfwMtJyL1wYm/oyfZOU8zP2j39B6JNKmgC4Zuo9xHnhfAJetQe3l2Do
j7rXsdARqpcBXmQIvpYBgipTpn0mjSOJNkLuZfZfpPdq54jwqhtBnfTdlzTx
pAGchriIxDyUGfDpnqhD/d3MnsmCPQRah0ZveEEPUV6qx3LASqBYPVvDPv86
rHqgdd+VjIqp6kuE1clmIbUhrFI3OdHn3jBCSafCfE9dwKoD+TrH2tCfOdnb
jMuPXuuH446cEC7+GLT1mwLGsRRy49P+krabcjkIc68bq0ditOB93vS1Lb7L
iGWZHEsW+dTUcx+x5f65LOKG7vi4MYHPPZzKqWhpzHeghVdEf2g8bfI9Jo/y
2AsOVSrWdDBjEJxI/N65PTdhkGN5mf0ffOnSLukeJTtHnd0evVg1SFugslsr
IzuaqRmSI+iV9U1bPKHGyz6ydNvbMd/6CMP6znArhGapXSQU/Jfx1lKIb8v1
FbbbUWVAcSwKbZTr1IPH1ROhD2VW9ACG79zWWtjIX6iphQRLMKEqY9JbrL6G
4bgd6oYx5PFzVNB2HSwQ2KP4BxGFNAbfpHl0F0IsxQjdMIM644dcN6UtQ9tc
qCDQbDNAI8LEXU6uCFVLeV8TgNcw3ulA2wXGHeyYXxMDfPTBmR38MX8W1hQJ
5M6U4RfQTsEJyyzjrsfBmQc5z6743ovRJby8QBk4+smdCLXYPTjSOJ+VTRd/
2WBTx2BZvGgeVoSPNhuOAyGQTabj/YpJRi/TO8z46BIr2Ou7IZTK3gz/FCTL
DwDclPulmVvKw3a+5Zs2qr4c4XekwyT1wSyogwD5UlM9pVJW+ptGouQIlne0
7IAKazfxjD2NbrTKfzt7fv6fZm4fc06giLKx7HwxR+/sty3Eq14x9ZbuYBJ0
/SjvqbQpZqVgSZ34aFQiRD8oOt8rNJWjNHUXSEsC4noyu6e67d2A/cd2VQyY
Te0R2AZwbnZIcmf6HbyMuXeSXh91PHzMfqfq1ZazuR73bWJH4w7rXt4m1uls
sb0TCIzXNLsDGk2PY4rdm8I+7y2Xr7FLoq6zn3NfQiYWREgRQrHruZYSYLG+
L1iuDIKzTlrhvWSf1BUQEjMd5vj4pR3QlVSrFfZ/o3vRImPQG+JDuZ0vGsoc
nrLN0v31sXDsXeQpudP7jkAvNzrrbVrfMPD7a17wjqaCyrWBASPNLXCztpYG
rAajjwPPB1vXb+mRGHp8Npxz3f5OwB9z50Da2lAdCBF8QpeSV3YmrH7fDm3L
kfLsbOHC/8r/OVHFOSdt/PlxPMAfYDKwNsj2GvDl52d/dP/3L5dKga2aqpUR
8cve3UZkQ0MVNQSh9BTY+2RpJM6N7KCxVVQOu7Y4RHNV3MTgZeqnYTPEn9Go
CjAie9rINkExBa+imT2gRsDv0L5O/QwQGiTI30oDj8BF2dKPxdaIvoVllRPS
3cd0FPe6GzYgWjR951eFtPgVHLyWkJyyalrhgQ+1BSv5JdcT1jroQw52aXEP
KQHMMJPzTu+OBHQ4F4mxTOkQdylU+yBGOGK34gJzw/kNGNVI9tlqjYTfAUaJ
1V759DCD7UzEG8tBvOZnVFNXED4jvemYwMw990db4HpkbbjfLD56mWBCTukB
tbUTaTNFAgN+JFFoiwVQieiiNsugZMtIU5CkMgD2SUhESgZkvWDTYh+AK8Fc
TRvxJaloFvTvY8RkP0I4HGpnH6kVviCyOIc85OGCkMxQsoezboATGyDIOTS1
mQb/94siqOTe4tXUwxs8/ylfE41nfUjWfzovSFg10qJggebaDQ+/xo8k8l3K
FDS4w4lBGHIq1Wb4egY04+Jcoluo3dVnzvp470DKJdhCp7uZl8/9Oha7jBZE
vRmDCGh9NCLaomYpgnJT4FRgkgjlRyCjBuIPsm5wTPNmZoJmaRvpsxM+nuR8
ijLFHn5HgdLTS5sn6XLu/AexQID61WwoV+rdlcVAoU9RzVeRalS+cLi6zNvV
oEcOWl/zkc391RaH3kgkDjtnu1cw+HfO470GV8kx1Eg+CPxGtXifPg0C52Md
Bg0bWVStB5m0yM3/ijRMyuoUuaaSqdKTg1slc44gLzEloG5Sa1c+OjxFL+1H
HN5J5cUdM3NTjeSWjGqby6yubaeevzxcHScTu1qOuVOePKmaRdQ33OXPfL3R
EyS2Qq6asEbRfvF+CvWLW3jmZJeG3XQWWWD62c7Eo32FLuIZoM24fV2sZC0t
kI+z0EpICdD2RPnVS5A6r4IKkxkaEHFPHXqnYAeHeanQId121WtI+cJUqx7K
k4COEQt8cHzUv1LvqJy5hqiP9ej5GODkp63GmD3LS8yponmzPuyZ3ajNLtjZ
wCD8wIDgSVgkryGSusrJli3xV/VrxovXOBylz5JiBotbKp+bVve7/sADwXgJ
hjunxhRYQQFCsh4IFGORf8aA99q5/wPRE5/A4DNO4QyCT+vniYNMDEoFdbrN
2/p24Cny5PZlYyELlPbZtIsjI0O9Fc6tvFkAijnebSQ9gTAWXeTJyEqO87M/
WeeK/2Mq0m5FjwkoY6FqQIvFNoMGZJE0A1aoGoanOxlOo29uRZboz4tCUbv+
PzWg5EZOpU8L83KjVAbv5ac2HUcVJmgal64XG5/ZxQ8IkKcedM37AhFrdxf3
Ad/lA0XLR+bgLLEOmRYTgNEO0lK2Z2ujOVE+mpagXSKjb2HRgO9Ew4yK2uR/
a//5EgFI5gC/35A/hT/oTt9HXJh+LaBwyytYl96GOUOZh9g6wErazI4miDLx
fgeY60/MJR7vQorePWG4tpn6W75K0Y5qLemcluEP/JIyqDXv8ZNUM22OFUC1
FiE3PRhvpQyAq8Awe0NARhNBnrQSApp1vNE1ZfugwpHEFHLtjg8jExAQw7lb
QD3oRYLf6+/Up/Lzlunk2UVmXaZlr3vLKObsFkcv8MeNgN1MpMtyxL1xAs5I
TGwpPkHmExllLBUbfsN3oM94xjF3xGw9whI89h2sgP9GGwXhe8mZDEJLr8yg
sXJjyRCxQzWyxlS7tEzGlT7Qit/q1upljf3ZfV26OLfjEesU/zIiTvj8hvkx
HmAsdbkMWsUcRale4bVpdNHLdD8UsdC9Qx+1MzK7alh75N8T/KRkDHFvJu8y
7HG63FdLzxBMih6Inv55r+D107lD1K0sT9rIUdD6lyCp7B4aAe6oLArRvk4D
9n/g0km9ajKuwY4rC3LV0JpURAYGh8lZ5zxDdkM+C80FrVcKa1bdl6EEC8YT
3WIsYLMN9qFha6brO/7uVIX+Z6pfC18xlPnPFTIysy4BMBj1a0tZywTtHQ1e
s/xuEjlJWWOIv9U9ODH/BIgvb/c9XHYv0MkwbYIXWY+ftPkKsB7qXpk9D/jF
6dks0Sx8Hfw+VCo1Id8yg5LtfQuwfpj6VF9CvqZbbiIgu6Q9NrFCY2EbyS/Y
T0F/5Y8K9wrOIZcwcDlXB9CMzmqa3i2mwsHFuCKpODiEg8MUoWKzb4tgVaU9
2jl8EW5byE5be06/hRrAVW2NPD7MCwdSY3aq8K5wsK+7G2ylYIn3opHR/N3g
qoGfHpqgftAYalbwJsLvmhswysj/Zr9WVYuXvNJRKlyqHDZrmuoR9+suSUlK
b6WTkFX3MgVBtx6VEpB2ahEGhlAgpQYZhvlCylWZLcdBKj6V88dCxgKWVqyo
tU2tNHb0F1Hc2jCzdf+I6PqgyKra66trIKSGaFJPRj5dgd97T+EbVKy3njLy
jaAjCwDlX1xTuijzGeIfHDSKwn5FykS5cR94y9k2RoB7TdNej8W1iUjgrb7X
IJp86cQxL7RDd71q9sdx4jR10swwchI6tT1NyzG1bAmIxdYjlVrvnWSSZPOS
dfBA0xHnJfO6pqNlVeGd8A5kK8E7jmbGwmF5kkdFLJ/+AC7n1MV7/7+YST7X
Akbr3TCm8dMD/rz5yvDg5gW3gejIgJ+R5AmQ+pC5+4Ihw1WqTvsCkIpMoIWV
M2LLdh7HSbkU8H8ScWh3tPL36Q3mVCDQzEhLmBIeRr8Wf4NjemmHJTrdUEYp
FnU3r1Y8Rn/nsFeB8GXnW2Uhhjgg/Z1bwZr27MPvZ/cGn0NGHcmoFlAp3anI
gjWo/qVNrkZGF6bI+ZBIi/YLLEVWdUzPCAcpFQQYWJtedENamjBt6itcnE4B
yEM99bUpDCMMXJfLs1BCBIzOOS5FN6rvmXElbX4R29xXTVjtwl7qSuv6gW7D
VRQ+CFpL+jHpFvkDm2WtaIjLAoiOYMFzB/Vf/+J33XDoF6U10wtMwjwuwPtp
FdIv5uv+EclwtKJEZquUdQlZG1EBEe5VJ7mn4SeAdyXKqKcFo5vf42n3xL5d
VYXoUOwv3/ZNe8ZF2L1L/41fmigp+fSPBzeYAczJhnv49uzPYAi8U4kucaB/
byWvx225H7R6PZvFQp9uAaddMKPpAIW6cVol+ecGmwfypfyUi4XJ4d1xF5af
oVdcvt259z/CduhsnPmdFORom592z+NzkrCRR3tXUaDuqbJla7uhA1zY3dxk
6Qfpj+ow3NHAQZGjmP+QtLIoI103YKF8IqITHAVvPoZ+84q0A7uP+HE80aYg
3gzyOOMIu2BkkWbgsXNuJUvh6bv8QF25jTQNETNfqLHfWO+Tt1d/7m/7aDtO
0nKP0wwdFDK0pYLCYK3cCUShr+snpmlqONkiGkWAThn8a17LOeo6SQ1l8TVs
k6TzmXZCKSeKagnrW8fXLNolpqo2QMjsYYJwb7oBfQqUmerobtwOOw6oAJE4
SBShFBCds6MfeFdi/iX6l0UkT07MnvJ4GxsrOk4L98VX7LhFxiC7+baylOO8
o0K6z8o4QucWmjOfUWzZZF6FrsrNhbxmmVuYP2x/1R+IIsp6yziZ61d78gGk
/iv5ENVsO7gX5vdObI7mHHuyWnGPpgkgME7WxS2gmO27LXZZZYO8gPpaNp5x
zOr+MJvccT+WkBQwhyof+Xe9lSTwKEuLmV5aI7utnd+Qcn5AdHXCQqIe/pJo
s3xR6dGDcu77aEvkfjCUZfL3IpGf0amrGaXPoS7qyLSJGgUEmQPAkPWnTBej
KrrHVZSFThjMSrRR7UqKAD8WGK+G03IXcsAKSyTiZ8Q7YadjKZUL63+UMWFH
Kj4YlpGu0Mf+p8oEOrrLyWFFU5rsPsjYD5rYTJJsLsChBVTsX20wpXgFMXBC
9IEsjuxa4MhgO0K4nad+etLNFLZIWd7rbKi6QqUkslxi3/paWcc6IUQr1RcA
I4QWESnmV6Upycau3OPjI6NtKgGpRHI/b7fCoRkFnB4RUCBF6PZ/ypFRX1OI
zJauCIX4sYKD5iEXwASvCnU6/jqGshbiTYM5wd85T5PmQgRHPQ/UhnK0Qlsr
pZ5KswuLEIFNF5mAbO6ydz3WW6B7Bc4Yi3I8gNwIiHp8PrwCjVEOlbLJLzjP
f04/RxeGVv5cRoMvkj4BVVHWzonDBnlS6nJ4TRC49vNxDMnBpStfcY+o3aXZ
7IGiJsXhV2RB5PFtvFl0qz6dKK02RMcT1RS/x3FlrgreRqm+XZ2ts+Lp9p/O
6XAWXemRN/Z7lQYuIfHnZ0tuHpgqSgwHZ7IRmU7LW0mWswc8x3bPt9hWqKJf
hZFQkjXGipkqaBVt5pVjSz0KnYFGaq6hx6YaCOMJOMuFkoIwdeFpdYRe2pcu
g+r90mOaok4cqDNbR6CuJ8UZWiS24aA/3ljSULCwfU6qijz1bz6XAmH4xr44
0EIvRQPGWN31+A2QhWVg26DasC1rckfbz353CkgC5d1FF0NIZcYJ0gPPrVC7
wBLFbFKPakkm3wXPDjW82+Ug+Ds+dV8KUxwjT1dEuTDugEgG2h+4OvgUSN/M
MJ1glPBHetAYjZt/YkzFAwqPTQ1JRr5PE53hMXcaLFmxXjl22eGs+OC3pEg0
/NKBnrUztcrN9K4WFasSu4kqCc9YwB/SKCmBhXpFnzmLF0dsNbgWAz+fpxUk
S8j+iKP89LNfIqAAVu2iOXEjWMmwslLZ0Eyj5DcTmLzRFhXxCx8SpVxxoTeZ
DOY87zIizxqkHlFsdnObagJdEsdXYzbAeFl3FEcLAyLV9C5gN+ov+iSIv4UW
sWr2zMqgXlL6dXbdFJXuQp7TvZK3YJy2trP0ip/DJrU63Dd9RSkl8e1Un2eN
3Umsg+8L5wjJ7Oj5st+zZPio+oBKKsiRMN01fn4rbaXlMKUNYXH9eBnJPpzZ
MWUETnJKM0aDtTsaOurgaz6CNox70uFuKE62voSuKkoFnV75ey5KEze2qZEU
pRiAmEWM01srlseFSAiKvPlxovi7va6fP1Wh/5tr/9PFIan3rVWah/DztWlQ
Ttyv7Lo9TXznGXNX+cE7A/QmgnEB9py+pjBiqVClqzBVMwaQn3eNnnrxVk5K
GZ6lyLP0LZCb+ffvwbudEAZX9pMAZOKzW164FowXenj3eCFlBGUHjlj8tzv8
eLiiCCYE6lep6j4dfviUhMrseDFp6FSoH1+fXeoYxjUXWHy9AEjG1Ba0qfW+
ytScPeSej90mK89Ux74gNXpBdtaov3V3YUfmTXSjnZyFGZUffvOfAKSwZ/Dt
8k1K82zQG/BJ9ArlqfbyEWLPqnZatS8GZqHa95ZwPah4wQALIgErNP7+FbBD
fD7cl5suiKnXXjKDGpR1QjX/7rEyQbGvRv0GUbIzOmDEYzNmat+rnRL0Xs/h
F3gQ6DgGRa1U0O5/J7Jznx3CAIrELKcmLCgweu8eHmFpEqeYLG2ec7ZgNFKj
TAzUhSUcLU6VlXJmlvoIprLlpbaf1qWUPKhFOhJ+jH9+IE3/Rz8l0irTzOBS
yX0v6DcTqOHjqxQ4GYI+hEjigiM8F+6WgrJTAgqVsA8bGEaA0FItp4QUKEHZ
z5IHkfTW+9tM+kl7mjShn1ulL/MvqDqTP2SLbn+NZW+AhbJ1jlyjf2XU5ca/
mkjqWuffjhhq7U2SGQmPGwqDNEphlAjFAHX4W+euYkLTXdYC+QQF0qzI5VwP
si1eYAp8pnOg+m2zV6e/q/cyETbrxyyzLeha5hMP13r9nnfUFHbmn638i8mO
vf9L2nCfl5AhDxIQRHZtr733LVcYzXpHoyT7cjwv0hrk9XHAol4VyUO0RfWe
SgYMt+1B7ZB3fb93NnzxmBB28w9zvME18fZ+0tRkHAQKwICus0r2AXcsifUS
7Akdx99at7MiLyD1PkCxmLrJlk7nS4ZCCsH5YuNemoNFr3Mjnb4msqUJDeS5
l/cYwVDvlIVLcBYMcQ/pG3jQZ5KXG0fc6jgwwchDrT4gUqF5Agc2GJfgAUm2
9djCP3WCgyN10pu3SKltIgubf97VK7vlfJS4K7J+0SJDo022YSX+9hRofm21
S0LJWFpYEp02fBeQCIaQeD7Vxf5oawDtSgEEqLrnzQI1rNMdZr5rIx7UNKNZ
TVWGdprlKkDDGb4f9fXLtzfiUTVeSfvB1cZ7DmoLZG5jD/QXHi0P3cv4jAPj
DWuGIQaj4mbdcQH5CnmCeExAsE4AvYz5V4X80Kuq8rv3CLCACjWXlSqDly2B
3SoVnrN5xoiROIN5HreljdQG30R2s1GOCrjlNwShmdjmx+ooOhqvvTMndyIu
eAMJR74p/iaclNuUINSUsdkqgHkYWu1ynUMtaUrxpbznKdgpJoa991Ye1H4C
RCOShzrkOgpVP0DNLc/HeroCjgauffkpgeIonu8sBfLnQqC8kofYYvH6MU4t
rgTsepnSRIhVQ6B8cDcg9Jnf7OJ03rkWmU5kxtMN0EJInlVZZ7SfbRfwbDeJ
gPL0JepGLKxryRtxqzvAW41tRhGyio2diB0gf3bevxBxSScX/6pT80Ym5gkW
BPZ8ura66qUvDZcth7TSU0jZ7HzFQCixJPxgIB++qZE+uxGlUYzx0yfRttQB
IgHkAZMgnIU3rWYNyNJSRkJhu8u0MTVW1a6mnWuMp0u4kzaVtUxKkPR/Iyp1
dsxEteB9tTsq3g5RXYFtkm1iLIvLibey8K33X+0eU9Hi45fxlvo4QhumEg5t
FlfpcIrxnSAnWjIl3smNyPxnU6q6i9M86L96EzDOmONf5SeLsF4+EqwcivGM
2zeczt3oVw4kufXC8UnolR2fhw1J3Gr9eKFWLzO9HC9hL02I476E6N25iEDD
wZgii8N3yBdIYTUf3DBow7FeVWy6VXo/CcGwKXEbBxXcxrJeEmpcgEoRfenC
tita04YjLXE20IKCXsOE+PWK+DVcKGdxjnFJ1ThfFfMOwIl7earEc6eEz1os
M9o0CMB9OvlT34GdmBQYRtqAuVf56DQXgErZhiQlF8P9LEyTDkxlVAWEmS0m
TOlkqQcYvdy0uioL1Z6BBhoPQkHlI4TuD8fSTNK9eq+XHDaeqx8lvD4FDCLM
Y/aZZV1cUe0MQEWq8m4qhFGKQbQOcqJwsBhyX7qNUTc2zVxCdNn0U7JQHa4V
I7d95JibjRFRAEMGG8h8/LGgL2MOiw6HUq6lCPUSFwjIyP4SSj39Sgg5qPXM
2Y+X6WWzPXSh5oqsWpn79Jy7xkJrQDE9aB/Hwavk0P1nl0yzWyBWSErBpWUY
8dovPkFKKyAAul2frnysNdFijzuximu9iTe9M53ml7GknSFtdUuv21KeXFbV
ylPlMy4WiGhS3pBlwDNfrkVJ3X1oF2IPKZM/2Ao/GLsVZXMmmB6sWbWpIkbk
tZJ0ksx7EtmIhBiQA5Id4HzFF8wpsk/VffBy1oI+F4imv3eooQAUNRl5meA7
olQjVJ39u2HnFoA5qwAx47D4wn4Q4GroNRlKabPa2g6mLnZcgCVK7P9qemHl
4dS9Yod346O4zJh+e8VrCeIBqcrXAWacfTiLm2Ao0MiEm0ovZ9H06sNqBHBN
KbgZuVyjRNwd6jjIEF7vI4SlsiMdBfKq0qd38PvwP8EaOjAOJFFx1sVlyTwT
jM7xACx6LAsL6s8igK9mcBIo37Siz0hji3b+bxtQWYGYzz49wOMs4bTSu5og
sU5b+T8a+FrBr5XpqVviYHfPuVME7cYqi7kqKwRIxxurlZuFDpj77OF3V37C
5qNYtrBKuaEc/4eV68e/FEg0nOE8sRB9A/QkNY5iTOKLNJlPj5FAjPpLYamd
kC5N0+PzNowsruwcW5SqQ5AmKUHZTxPRlYtq/IWtk0OIiJ2ObUkLhdlAKXAb
4Zf3+l0UFySAt3WmgNIsFCTqi7ZQhgE7ajmgycR2Tq6iEJI7e5CHX2yKpa72
FrOuVZSw00k0CQTjPyK+d+5Sszi7mOJfdZprCQM9jAYJrgj2M+h4UQy5bJ0i
7a0vaREYioLMhozg/K9XILVIGPZ3i7Mcc3Yw+2QXVGjfN0eu6LJ6jLRdB5Rg
bOAG3WOEF0sm2KNkunl5HdHInuWFubP8oEHDZ2MZYIFNisULf9yzuC67VV4P
VMj0ygh8vf5wFcyV5hReEyelfjxAy8ZlVnbM9088nooupbTyZ/wXsgK5f8JK
SWhfAx5ztNslbI9luNRCOlHbCJhRdNLgGG/2RAUgJ5tXgT6jia+lw+tcIXfL
rVyWII6OJ2VczOkeE27BZ0l4MloqMNxJYXeEoMbQ3rQfeoo2jBS2xiohxDmm
GM6X5NJzvGXgreou2jYNzVRCNrGuQnBhS4in7mexuE3+mDh/ApRGrTCKp4Ag
09Ig+RSfcLQAlHZBssSTKj8GqN2MDBU4afkNxFjEHoBXqYjiI5tIuqZ9cLKJ
WQUoK+U2dRQJyZNF+JwV/kRbtbDzFF/gNUz4sA0xLb/RcG2sOAPwMET3TGtP
mE0VT/UXVFu31nTz4s1LlgcQAojva+456rQK7uR1khaIe5AlxMRFhX3+Lca7
BTsFXLJWXLMhaGo85wi0a9s8xSIEM/7CzKHRLTF23zwXxnknvTrSNm4ip7XJ
f6ieN6BMOmuHJu8awMtxRibxSxC540nhOjsbLtQ90mXVayZsPORVG7NGIW6W
8bbD5V0a5X2IbRdhFBLH/blc4o5GXH81qHMPvDJvMy9i9BGtmzmPHrR1H6Oa
dU35Dmbex9Now3PGdpyGp+6uHb0hFtVzG8aPcPfO4scr8oFUB0nn4AnVCz9R
XoBn5qAc9vVKtmF0CEag0l7PXi75E1PdFeEtn9ngM3tabOYGS/RHmUK7K15W
YZwl4erYyu91qHTL9JjQ3ZHB4V0GXPav8dlSQEHi51e3nA0Dgk2oTaCBd/Qv
nf154bCiY5NcQ2chRl7TF6g/WldwiJYqdekIbpdvABP3LgQDJiitocGhe0jx
bpLJbrC9WukQbXT0khEIBoFe2l4/YFff0Jcy1oNbgMeo/3pr+QU6TscwJeDm
1994jrSLwsBOb6sRruNXGMn7woVqhINIPQspE7rKHVyar5XLI7GkRRzlWrCN
s7sdGJSStD3xz4vXVEoLLFqcPKdOvFfLNDrQZkgEjicXkBzk8H1/JHR+pNuG
UAtyya590nWEOiMQL29M0gHRxqHp81u3mHZvH9ZkZUiZpjfatnzMolVMaL2g
WQWdebkqu8LFFH9KVQnCSq8U1VL0FOyHEBTfZoDyxADOHpxhYMZnSXwjlHDc
GRA5M6nvS58+qw1FOeNH0nTeVoSux50yL+INJeZBA6HdqlHKYpG6At0cRi/1
HfkeYPtUYQwOATF8AZLnTAMIJ4mOjp6C69Q9eoxNjcim/NnOidDwFT7dyKFZ
r09xd+DIBtsfjrlYdvOEKgjW5rLuAGPjepHCMqlQqZUdEoH8hpPowkJwith5
9QDJWXcNZWrXUNE/S8nBxkE/W6JJbV2ddTdmYcprbCaJquW41pt2Kf7K5t39
sKzKfSyOQaGlTXPyWv8g7ZUx+jwvG4Ic0q892a8V/LbYJjUsVnISZV+0P6Y5
+JylvTsgd59cqzrp51lyxFo2SX1qX5TQiRroGncjqpX0k61QVzR2ul0cIvTz
RxS4vXwHCt1/n3c1Uk/huAM1JnUEV34BzCCnjpcayR5KBcMX6uNMqEh+HI8r
jOC2yO8KS8bUzUT5UAgSK8kP4Fv4o7Jvu3eKErX/LEErO+GHGBKVGxPhdCKh
J9ZFm6eD3Al+PWn+qpLr4Cv8jQmF6w04nvwX3LAHs73L17H56zGybsuU+594
ACsWjmBpwlrRjoWnT3YuwBS6yajPsVFUoUMsCnKwn70paoacMJa9X2YLRFj4
YHphB83NTMjYdKH7mJXgJJe3VYYNqVscn3hXWzd5ULjmYijizk9Si+N5ggts
9Ff3E8hXoXEFwBafqzHIeWJKJRgFxigg7+OPm168SQSRfSPDhzuKH5NGR+8z
4sJX5/UkALvE6AWNYthSWCwVz22+QIwkwaa6pzVdU2dLo8GU2JCiXdZFlrKA
4P5Rw8w4uYZtPTuY4J3JffeuPq0Vlga0AqCMiCdbDG7f65Luy8fTtDVY7czL
nMR3zW2wnOYwMuGYAYA4qo8doCuSIo/HsoU56q6uYNK77Ku+Lpb+tMc3LZBT
645beF9kXxVqYI9E+fLYxw8vxlXTEIDTJLNBMreq3dp4lHc7BydS4wnCXYwP
tdVXoHSjmFOvNsFLCBcpJvAU2MuqdE6gt/U6KEv14V05Kudz6YhNCdyAh3fS
kW41iN41bTxNzg9yIZGs9gbMlcVfE1q0U2CxlwQxGzMBPO7ISRToQM6zJG+N
uejhgxYYqtS0v/GKkizy34g/QzZEiP8yXIQxrtC61/xTrVT/5glB6RO0JCS6
jzElo2iD9uZ8Jm2Ukg1q32wJfVv9EMURiAvQQqC3y7yDjZdQiN5dhcoWT35t
WNQDIG6y+TSQhFprpR5DAahZn4hKfUKcDm0BE+A1whyAHUWNfTNOKZt/gcbS
9rzzvOmKjQs2CbNrSj6gPBn4SWQzjozlJeqgp9crHCXKjk4sg9MekWLul1X3
6tA2NlaOCPm9CKq6OChMftltAQEAAJbz36FC7oeIBeMiZX8Q9RAFD0nVIn6x
57jr9gFw9/Gg3u1PMGx2Gd4SuU2QqPHQ/MCd2iLsr6Y3kKPxpgmxMUx/Nnr2
XqBNWCso71S5gPKxx9kzTfFDXQykW4BDyF/66vFat3HVM3xNztXpAGExTnK6
0NzngHnHuSTiFY5nKhoyOf9GyqIj8KCXKuUuuS/qejEWKqdBIi/BxSjDxrNA
JdCPLnFzOO23OyXPQdYWnul/r7kBY6zXEmI5x4at1pGOj4ZUvE365W8Bhnf8
0/EczyfR9EHGiQj7aZCEc6qDOYDJYSfTly5R+yIZJr5J7ULTAhRVmtjZQ+cy
QVlxF6NcPGvwXp1cQYNorzC2V30xVBpIGvACr+v8dMe9ted+zPqXPpBJ4Wgq
hNM/7TSGeP1rVX//875vmoDJAsngqGnA0uwkfhZPAQCHpX00z+4M9LGHmGkF
YzXC+iKQ+Qv3yKatqb3YfqlCGBTA319T/JM0jcyj/kv/NhpNmQcrlzPcLnTu
hdAYknb+kdzNCf1vG9E8ikKnteUIpQCjnGb9L7ICdFvFFCirztH9jWh0JK2D
fTbpCciQLc6OZgW3KElP4qBiHaj5xSCPqhV6ItkD0CDnKEhEFTX8iDRgyHay
XiLiNacq3QfBlnrXdEbScD6hG4Nl4yhTxQ7NDt+ax6+i4dmYOeJht/oZHmMw
gpR3Grx2PBm21+bZOxi6/qAkC59QUrXhsRFR/ntStOYItHXMvr1otD00nXiv
o1ciejwD8Hv9zvUhhD5R5OCjKtFHmnq9apvcSoB0LgEMWv3JOApJOiKTdlph
zYz939ewT2YTQufGA88XTsOuxV3wK1loTnnkFONywz+oaOrB77Aps4uLFz6y
LwNk45+vHQAmudVIPL5L2Jm35MHHE7trbKHL665SafCtvJnGmmkGMOFpRgMS
IVA6pVk7KvVN2Y/FnewWFmIXxGqA6YgNXqY6bP5M4Uiu30LjlknzldcCQRgO
EbkcrrE4O9iZZvCWhBRe6RVNvDPBnQ/Hv/3w7j0j0KpKYvrAJeeY9ucy27ZX
ImVtOsE5JVCgx5uXMrTk+8uub26nPpicV+WNdNv2r3OusNs23kh3c/+MQCD0
88m0QrJHiXtsI2MNxsB2epaC+PkjCY5/sB/JN23zdFtaGhc7jOMEwgF60ZqJ
C87jzHxFAzycNkQT7R8IA16oOSbEDPzgULOCO8AU9b6dGP25kpjHBovf7pRZ
vU8zGYxncy2JTIKJFC3RfMcIHBQkmZohHowsecxhh3uBj+4ENYBOFF3npOB1
4YusaPc7R2T2XOYJCHMoa3GAoq7NogZ6HwxQasKDuPm0OgWWu18NVXul6Qk6
kPaphC5msTCr4u8YtnVS+pseMnzJQ2/K6eu14VaTOtUPd7oCHqMIUB9z3wOX
51CFjiFdA18wrck37vImt0tma+ILMNdHVJOuw2EfWu26dl9Y94QPQr5Zs3wB
yqtiWf9bBTJX1a8l1wckqyxyTaiWdirXT1neBtNFf6ei1CxHPz4kZ8zeiP+f
QaAG6zGs8si//9OwCrJpmFTnUS/ycktXfCMU6HkHufy+1eUZwSENyq7dkgN9
HvOUQYWhLDzUhxNFzzJ4GlB3w27L7EJNjyPn0Odzo/mdBz6YWSRza3evWjpK
AF7XljxKFq/3ShPT4Vd/GY71HDdhVEfxtWi4+EJFCGXEoCtie4Md55TKlj/2
CcdRt/WJElqXA7kSq/H7g2Fq5Het+iaOHxOpJyqZNAVPkpf2pOHFd0mhOamC
zzgfT8L/zezFTJtt/7kz9nHIQZh3lUiBNU0u1S5fGTG5fwVQhcrL/Z8/sOkV
SaTLBQetu7lTlxWiARDCy/Bjo25nQXNVyq0Mv6OiVDwIm7OQMkT7QBsnqUjY
/yyeTLZnnrbmSpogr0JTsmnj+Un2Gmxic58xqDh/jVnBIsRgXdf85eC4uaGO
56nwWkLGeB1tdH1gck23oKzLf3BY5+26a3XPcP/p3aTpakGSx10ToN/eT3G1
P3dnhOZULhLdcRjJOJnIn4P1394jubDZ0aDCGQaUpELo1ZwBbFVxmQoSw8K1
NTbK30HBXasEtqblpD64z2P2pP6CbHSwy8hrKtdtPbAHB3tIMpPs3OphTiry
+4c9bcwCzpzBc539Gykthrrex4MgylE69pL26Pb/Dvie8gFW4ilOpSo3Qs0G
3Ntm8Z5r7cxyqB3RMwvwip4iex6qlFVpsx8OP+LE0J9WWqO95xcJcswOx3ZN
8hAS53QExARlgt/DVOnAuxwpQgMlJMgJAsSGP5rcIDm0yV+qLH0FllRa3d30
BhWVLeTKI2zdTIoORAMKYvYheyjVuRfy9vBGWI4hXbdowUtq9XkM7NOTS3ba
aP0dVFs3baz0SCYC/1Rpkw+ZgCzZBd2YgnOc11gyrhRsFrH/HOPKQNM4Fh7P
5QyLBZXV8eeXaFkszj7DM510TWaYyjBIsCF/BTlo9IDz0NqxhL6Bdx6H/P/o
B08jzXWRqkUPBbp2GEN90EsEG2lQO9FLHTLtuDnMFYifSxzIpwxjC0JP8p+R
wcT7Jgns8R6uwCUWgZ98UMCxrbhT8NuKNFxV4JP0JAWLgxLf/+4uGI4WDRuL
ZXQ4QIXNRngsKbIHHkOzE76pwQGhy6KRUKJlGLjaoGz+mW1ej1UPZS9xDvIb
s3XEy4yu8IW295qPS5RkGGBRprIsJbBiNIismWMjJXnJ8LRjd0/Ovd/Ydu3V
DRwr6lFjhpoip//ZZ9QQvHo4+QuM0cyPz3ynx6SjQV6sw+f4t9hf+cH8qty+
kQD9gjtGDSgJ8+ZdW/iSvmTlBCBHD5F6WHbkDLnaab+l16LlYVOjTH4S7eOA
vjBZ4LIxMedwlXr1A84+DrvKp/3upy2FOZBhlbdHGTuE64mmA5bm7mGhdG6W
pv9FwGXVHcwGhjVyIsKPQTnwoajqPOZx6D4dXCBcc4+j0BdTB0QTLtqviPCE
EdMq2wwAcZAdanViSJja0bENpLtqdaAjqlWKZyYcUC/qzxogrYTb0kzW8HxZ
mSScRsAutfZq/UGwRgNC4XcV3F5K3nPcWFGKrtSHSZSzBdRwJpxEqOUctenO
n+7G4U2hA6mga0Z9/O8Grij6FBhqcjmxpSMALFQOC2pehJ2n94qo5FjUmuih
Qo/dW/Wk0TzRoeeuH18wUb+B71hvFr8C98CfEkUNYVZqVNgtZ/cFOwm4OT9W
V9p3AnVG+knqpNwiI0kLuxQJJVlVl62ud0BAUM8NabHreLxCeCaOF+4fZVnv
53Y6sXX3QUa0TD48ZAZbpJioSbbfbOBUAufpcYChxPDBOYeM0J9BABQh1O3Q
VQZ7vp+yOnj8JnpTjM9OC0JwQvxY52TlmMckInjSR1JToRmjoAo9Zgk6XdO8
lIRHYGu95yAT42NsSIx4756pLlIGMUKeZMO1s3Up0gJzVACJdt2ManJQsNBy
zAsQc2a6XZAc0zrT1X/1GAsz34jER2HwR0bOuD/sRDMV3/9KgW8RmOLed6We
sd7wuEJNkmlh0grA3eFjSMzVzRnsL8P0KdlEiof2VT6V6B1ML2KR40fCR/P/
/tPvfyWAWk2pUSWOsFSWLxh4mHEOux5ITErygjY2cPnsbP2EIu9zWxXEcDB8
y5S5tH2noKdnA3P+PAiojPWiGjndOXanWcbNBBuQPTfcnrrf+Dw3X+8MpzXG
6ojHXpF6n8DSstGRr17CXyc0sG3jRu6beG0ccrFApD/b3RflEb85dkCyfKmf
62HfKEEtoNy/hRuLNGkjiAecS27C8T2aRfUEgXagFJ8iyiU9xdn4FUmdkDVC
gxcct26fxyDjOWVPdFMJCG4/v/eIy1KPA76D4RO4NHUySHzsiAsUBellIs6g
9u7KfrqgbQj1JTZc3w/tRaGjFaw0dX/bBGNPWF9bvIHvwK/UjurEyTRNh6MZ
R/pl6K26w/S98czg+pb6hgio2du0bRjMDxTCv1CN4VaLXjISGTvQMYXBNKvK
gqYjfimdKAi5bybWXS51kYPeyoFLEweZP+aJ45Q1jKkUJnVjeuFhmwPyWhK6
PAT8oGzTA+KOnx0rLt9jXUDoB4CgRjE//g+vHLDmInQbtnBEA7bkf0RF19/K
hMhtZZpTbos234NYemv36DNHm8cQzaqEh2iD8TnfL2wnPqwc2seF/6vN+oes
yR/iRXkF2k+nezaVCTHw8QUapgwuCIjhc0cuZnziI8o3ZrhzoaEVz62mJ5g3
3YkcD04QA9XkT0CySuXnoxMONzGwxZbINOn4/29y3EJVrNUHn48qLkGeTJya
mH7g9f/kge7xrP1P0pjUq/rjfMws8T+56ECWvQj26smctscMs8PpzElVuLyE
B4DJoeNj2tEpI1Zkw0iaWKM5xQGaMxDoNn+2s4MzZBmdn7+EVIUrdVS01wuX
eMKwa7OBVEO1HAD2nKOdXFQ+IrAUzpnWsr4KbRvmX2w3JGrwfkpk80FHSt0w
uNeuuna40+1IzmtfLv2Djf/5nrMlemVQft++XX1oP9dy0rws5LEiWMx+gWb3
CTJSxtKJ4OKM/s92ai2/M+0Bwlxf//Lct09pgwqUj3H0lLTSh3W43N6QSMZM
FzjUz7K3MpBtdCWasmMg5eWHcWa/oofnyb/3iecDRNxeTvDVcSEjIXkwSLwr
ntKpDeeOiyDeMobL1Q1RkganspdAhZnsWBU1jBCkQXdLsehMqNPf/eCRLBbu
rV5vuKz5zJ4HMjeRdilhZ6U6TAEXmKDhA3X0nx02F6N01VyfWKXPHEkrMjUM
txBv4Suvuq0IWK+cr069M/LBwLIkDh5pbImtU8LAyU4Rd06K5rHFvsI76coa
u7OTWvVXoPHa62Hkcl7GO3qnJWK1PYfhEsmIRDitQpT/PO9xLq2CI4wLyYRQ
LRznP6E9ZrnUCzLTYJd3uc8vRTLvvLs2tNC4mX+HPZu+08IdB87lWhexux7T
1+qaTES+f17s+KuAT7YzNgIWWDhjJMyF1qHwfWi55WE6YPHReeNnPGKzE1ko
wwenWx9tV50dKMZUa13+aHk2f+OcTymTKAy06Lr0cfYT7zVmMvpldBtAgLQe
7SPzoG1hlOgSH6uB0o7nKZyJRieqccyvXcHSzbkCiBvjg/xX8dk7I2rwOxGy
q0bECAj2RGwMGjnNiZwagkIAzjyYeVWUm1FviywEZAUY5w2ZPxjoo/KfpwMS
2Jm28lYY/3/DsVkgWtucfQEUlGcVb57oO4fgXdzGUUkPNkMzPbSngKcjI4Ev
1U8QJE4cp51lIHGch+kUpsY148Sn4vYBcs/HVfgjO5WCqT3caG5j+r/RfNfQ
J6Jtq7x7lXOaDm7PdYuzKwuhuEtuLfsKAaVGmoqSTu006VUIbOFRM2Xbgf0t
lnm8Xi5m2mK3Nu0MTuB1K06K++HZ0wH/UhRVy0Gw+B540wQULFi+ECLjsUm1
weRWojFHk8C1CXyxOxwf3Po5mwMFlbmwQ1/jZrx3uw+nP2SPSvBx1cJ5iQ8k
7i8JmgATTwu12/jLCsFGJtfI/MJR/h01Qj51sLHhnTTf/B7KbFe0FcuEvymp
asA3gcIELp4LMuuQfFigxyIWuluk5Lvrb/YoZi+joj73NExNCPhzsqQnfYAd
cMmJjkknECnbKhLMjXuZzejZ0FQupJag7ezxZ92ypnfvmIoGwN2wKR09i4eU
EgZ0BB4e1D8w4uduk8sH1Vdr7OBUkQLjGAQ4K1C2fS0ZobmYP6tILKCdZiHd
by6kRdZmL+xeK2JYIJ/Ghb9g3lrYBytYG1cg2Q0MAXv6jHSZv0g7f4ps70/D
hiUkKbi74Pq0kl6za4YwE0ZseaPMKGp4AU85F8wArXn9pfQbrZr4VDm6U/HD
dx8GD23cuhee8sUNCuoNOhml0B6v+WIvYX2s4MBspWgVG1hyQRuhTrGIbS5Q
NMAm4lhM3lxIyPFU51+Mz6VYPuMTjf5EIFkvl8kb6ocFHtOntKhmvWVI3PXe
/T0IoWHVYTQq5H9qH7S4R5m/t6O7TFCbDBrVoxikA3K3H7GCTNTuNBSOVHrk
ipOZOIHJDD0fqLML05Fy40DdSxKU9TpgM7fBj8NA1jtDKt9LK9jUTlF5eHJn
N2cCaHyVvbGjtdZzRrva28fa4dISzkrFyw+hebkEVhbEac8ZRg0zR2GedtwD
EA8K/3WZQxfDiSn2YgL3wUKPzy6OuHucpv0/H3nX04ZmvY2DtIZqLq2XOcLj
RyApoxtCKTyZG9jn2tbeaP5BvFI3sGTp/xOBkTnBQXsFva2f5cAJt/oPEV68
iODRJpi3rKl9R8YTG/Ue5F7p9CBxh+5pJHt85L3y6V9IahNADw2sk39BFNjG
w4JqKiNi/W67pz00+tMLPPQvQCrnQJV18YxrdHXf1wMEDBOzE3RBEHGYYbK0
E6n083f9/0WLIFkj5lUx71/ebuwL4eCqIlULH2WFH4UAq+GBIj8JeRHJwNOh
tX8sN9nYcL58lKedDMMcuEFIx9AyFSE2Jy1C0INkVr1NmDzKT8iIc2ZRb/ms
6Jrbno3WyOY9y14PseNodtvZXaElIgrvKOWMOHtcefsSudINdkByrutVIM8+
TIjgF+o/3v5ENAtGigNxOCcJGfz7JWfsxvKGSdOiUbfYTwbcKPMlWoVTrBia
6/UXFHjzbQjHDT4mJGZBym+HMl4VH22Awt8NNbL/mqlo3VTFoOysL/9gpgkC
0/gcCwuODppu9XonfGufRzmY3A+qabH69n5k27bRnmtAQUotYgVHfW48sJhW
4wqYOsj8kG7OQZTReEGFK4q954L7nDw6d6x7uvh1KnkqZ3cq1/nHMigql6AX
jM+qYd6O+z0/W944kBK9k4eCbW8AGmKJ7Mbs9lCAep7IkxGjw7riXFjRAUFE
7DM0HCYqXeJ69y4reIDCg2QMYGtjAUxbjTOM3DgumBDsf1IDNbmcj2HQlHl4
S+Av4FAfcbhKr/3B5gXau6OuV9jx9Spx5iHulKEuXGEGYVmd4m/ffkXxGaBf
WE41m+935qaYfurkj70yPuoHQocs6uaQW2jfn09QRHKAeyUBB+c76sV45Chq
uGIz+lC7wMT7rSDNe3GoSI8QNlWPRgVOGX87Nt2xUS9FwndPmUghdREKNFCb
At/5RjWdRk4QyF+QsQnI+pTXgqJ35pepEtja+LQG1v51Bxggm/fTBRlhx0Gt
AAI78KPafVsjZdPHtZEEmTyrtBJFvSoDnhDpiwxC6P7TO+STce1sbdVTT0By
H8np9dq3OP1DIPbANMoork/UyOLkXRR44q+8dOnCvMfbUZ4k967SoLOInD8u
AbHj+z3nUbXt1Xshnv2Tsihftp0BcYaeDjSZy0WoDVZhWGnJTTi5VC/MYZNN
578cTWJ3Fdtsdvn/PpteeT2+7g+7ONhGuK1AZEFItsyxR/lGSKBuFwusH+XM
oXI57INbd4YffQd8+EgP//AZeI0C9SmUpWAeCH6Dnya7oiSJfkzE7P0HduHJ
Bd32ZyDZ0u3f5aNnJecMeGPs1Vro3tOUqSQEr3gApBPVPkMCuTo1uisPU9vz
CvlOPUxNYy1ZUI+cGdRenzrg5qqzAgw5gS1OdBUO0oNsgnjOQyr+TdvWzThs
l1o5iOB1hzjDqWMnoJHo++cMaSCBw8gTo0cGw2hygODYXxavgqCLctyNoEe1
kKYbhI+5Z5YJwNU4JmQ3V7F5uyEsf72xfGoNgtwzhvxNnx8yR5hwXscjMpSU
/zf+WzUziVzliwAtNGPPPdX33P0foytgcqPb6QCDw6LrFxGRBYZhQpAkHAOG
gUZ99YgyzDJ8DRJVH9pvgtLNxpmde5AG4++iPkHgu2If7oHSgU2yMaXvYElP
iCHMExr6eER2IU+Z9iwtP8nQVvIOoAI17favh69sjTyPeAZaY0nIklUNZALA
eE1GkQ6Jmp8AGKgW3xx7NhgOnjI2abz9efZTzMRrC2HJZa++rz+uzS3sjEWR
YcmzgJ1NBWUBqmaxdhXfWK3ym4ySiNoy4aS2VHgNkFbUnSptMNk7gjxI9wTH
Ia+ajZXHoaF9UVgMoNStU2F1/fLkx/jvCxbsAGNIV1DFUgG/YKM9AiM6ERRc
U+5zRwLlBcwXFzSy8uBKpXze9WojYwac0TsHh0VbemJ87OEBn75QNiMl+kky
mK4zgu149u1uptdQtTVO1ckf8AtjDyncCL7gdF/+dLkOkgTT0hl5b7Drn3e4
tVEJhHVgjOGy3ydHqY0l9ylQS1tGnM1uNilxEYEYYDPEmaYsflm6TiTTgKfb
EK6jleKcf/zrMs2ez6ZWopXtXldTydxX97TPc4aeMUnPOlLTx3Agi8jM3iiE
OFLR3kmIS7gPwqCCsVXmbnE/q56KkMoq5U2C3p0MASzk+poyll8cwmrzsrQ/
WEeO1lDzpQFZw4lu9sfYsdPvrPCs5IV8TLStavIli2hjCtIS4nljpQ3oXijO
rRbS3xCa82dq7is/AyH45nSOv8JKswqBEL/XhGffS0PhfZ5N0r7jEDFlF4jZ
ps1TbmgnCtuCltQMlqmaHXO22u2Yr0Vhh2eTELesJXb1w1D4Rcc7Y1mDUYOj
53PVanY6AxiK0Na9BQjr03IYb+W9FY9YLuPo52HNudATP1AEaiFrccPRWmtS
7ZDGxAI/PkUkuYvSTKSYhzV0KEsmViWLxveA2NJDj3BAEQbLWkoekXlscWsc
nyq/FeLJ+i/tZFu3FoF3AHKq2JlfRL73tj2f4jcNf7F/xMC5wuCoGwspD1Ho
pC9/UCDzpHv4mcEKqYM343Cm1uC7JWVKTYzs0dwpdHaRuRRNi5g91MX4CTuS
GRGuGYdV11YD0S8CotTol2ghqBmNoP+wczN606vSzE1WWpk15aJtal0qWgqM
/X8j7UJqlCp+3BJzOPPlEJ/0JQmElDquHPXL1p7CDUHII5qUXwM1zPojdiJx
uDfyL+yML0olP1KJtL+oqco2THRlEQbWPM2EzJk4P0ryVeGAW3Jv8swhOmut
DYhVS6tqNFregIGo5JCAqWaj/0JtBO4kOPpWKOiMvJuyp+at3afFUZKWkLZ+
qwKcIQtFba+geCP3AIi4SK3iT415DfAaRZr8NXV6SACBk4NDd5a4hFcIntH5
vGb4ZLoiMD1RoLhEsHhMfHrxqE4DxvZNa4ptK7c1zUmUe7XbXbcR/trgHB9B
DTWN+xq6voCVly8uFj9Hm5BmHoGDGajbpglMv94cROf2OSF3gCuAFfRlN3Pd
lYAOp7/vlUlWn/pzag4trSa/pnnn0AcUwombNJcekAEXNX5WkW99jsLbuhef
GLfzW2upufMfhGzEJFdspDiKBjMzxfSCnogZJA4eKfq5ngUfWI3xh4YehyiN
83LcSrGbPTpER08HNgjAVa7wAmPS7JhgYycVhn+0CP1OiamD5E+ExsLLSZSP
c7fqLv16iVeCwH2+6k1G2j3jyBPeDzzkKFwALaGq2jdPIbNbCzXW1kZ3pDUh
IlGsCfpMLEBBaCJDvNGQJRwW9Pjl9dkHaewq775BDOsztvlBHEs1VYlcjBXt
Pxl2dkKjMnu0X6YhCV4BWGF13NEWfGBnF+BWCWC/nUm5s3/fXIptX6sl0FAk
4+TUEhHYXZjL4YXCNH5yWtDgYd7b+n3tE+7DeN4KNJLC7C+xVqnMEdRXIUKb
NgRiz/o66/HO6ygGVeF4a3uJmbD6aH7ZhN5dCnSYFJRbnBWWW6BXTc9adhMW
csVljXIXo/nB9ytj/eB72eapf4C1R65mnP0KQufSWrn7Q8GifzKvR/prAO/B
7jheJuzajNIWlyg/RvRBen/GlDNW3W0c5jQz4F7UeMQztZYgYyU/X2Z/ZI5S
vlvL9/0cO2+E4TKOj8D2RbRCY9qo/sSzcZZlyduDR3pEk6q7CGYtFxbJbJaJ
GDWOkaXZTZQpqVJ/65mrv5n4XGGNrfkqhlVG9581w/JodF17ofnf4HoWXh88
KNYBIC+oWP+46Bdz1i35Np4jz3RCDHr0TAKl0UKeShnJccHH0mPWmp4JsMBr
lp6BPVQB1URT35Ta3P9bALPbml7Ou9mhRPZPSUYcVtUd4Zqo98N7N4Kpd03Y
VuFeg5ieant+e7in46FsJdlB+v1JC1I4nQ67IgrKSC5aGMXiqBehR7qPeMhG
HnQk4gkl0POhOLFbtGYClcu1Uk875qmqGFwbYmrUhFoqSUv22H25ErsqM4Yn
ehkgerArNORyujlzKtyC+YhTmV/rU60JtwaKG1Z6A0NL09lmISuf3ZdlEKAU
Ocwh3OPtp6cq+LXL6Ve50yA1Y9F2YyIChN4sSUsbVK2Hk0OFrHbzdcV8Nrb+
fe1+xss79PfREqZIjEBjFQxnlwA7/GEQXGSqBeA3E75YpwNYOEc4y5zI4Uyi
PbztCsr+GjXVZqa9jh0L5ExYlmBxrlAP45J6AlBDxTVjz04xsCAVDuqCOXNt
90w43wYLIjai8N+qB/KxbocDYziS1pdmbnuDeY9knLL8F6lHaXIsV60ud1hs
K9Xh2MrhUNzqGLNaBbB9hTMWpVF97zJmm6NDzP+ACN94ruivce8rIvl0FH5A
kpMnuNvuVHSQfCZJjNldb3lGTnvHt5lOsTmHzaQuXG5Qyg/OBOPozVuYyvk+
NyljRI8v1sC5aaPTkdZVsYlI1YX4HCJNdIP6BloL9rSCo+KfY+hGFcjjU+5l
CkOmx+Hay6rQVp/vPQaOp9bAe+k6RM1Da+O2Ffj32YVZShpQTtxnLOnExQzk
asJRBrf8/A8YeVn+Q8wQ+EzjG8kPCyOT1J0uBwUCKl4eyCYQGePIY0onzZe/
aomLRSh5xby7l6Zd/ORjo6Idp5MNVWIyDgmTXtexLokie6XNmz5Y2eO4PI4N
u7jFMRcsxF5GxfluOGDM620zVPANhvR7RPXqemsbXY7LCeFOWhha0lKgN6qM
NdF+tnsvbNO2tKca3li0lxDTfZKE7SgG1xKORLSVsv3jfblh5Ss918eAZdCp
nefuxyviSep0B8XzdAzpnmSJ20oEU2NUDfa3UL0d/t/e/+xCgmP23mmJVl45
TykZ1zwTSrtJRbX1469G3O2zIgYJd/FdT/rVNslWKLYse41tHrNI0Dw5J2wj
dHJObZaITihg/D0mAQEpr5p5+Faroifg0RsAm+IrNbHTCfTvwfZ6BjQrnmWR
9c7KjrWpeVhmumim0oochMUSSE+NJtWdpg/tsPzvWWi1ahB9Nlebxxgty+qJ
6nNNgI2Hf/c96nQUjw/CaKC7u+xQoIx9pquPuVU8ImBBgjdQn0PQORrYdsZs
5SCoyLZpEagHu3cbteuB9pArAW0nxA0NotwwIWWI9Pe5JLe5ukb1MsIHQceZ
SyVaTtCg2uZj9k2kwoTEy/gPzkexo6wFhgQPNDuTDYgsRUDuK6bSnp1ry1yb
0T+Dr0Pj0Km5W7yd+wyEH3L+THHqNshyKzI9ktCdo8Q+o82PtPPl3FBbHYDq
/eD6r7mc7du30Ek02X3fxWQHM5tfKTikdD7ZCvYdpX1PEwHOs9d6e3DgQIQl
8Re9AEcqOzVr5pg6jT8NTT+5dXZWgemdqwauBNFzgMEz9FW0sgCxlpKohv8u
wSWrWyM8Cg9HcUwkkpAKouBZeYtoa51SioNgaPm8s5550G6nkbdRKaVM6GrV
tiR0w9eZGQQsIjnB2paaMaSIFYlXLudhLhRf/55cw813DI4lwJ5MqYLy3uzA
MJZIiOHHkhPmg73S+bLbyra3RXmU8HpLRhsIe+KdGk7AKBV0ip3EL1fTtKBv
jBE7np2du2PwRSGPsBdm8C9Tc3wTZzII1ijMcyziLGON5lG2JNdzaG+A8GmF
uPEBbI5jMuFNkhe+jSpxRbAc1vLINgGwnSNHce80kscFXa3YK7KSzp4dmkRj
gEPm4MpC4K8nFwWOfSjhUG0BhpbMOswFT5nq+7OvJr6pH8hOM//nD2Xqgsry
X+X3tvaCWRNqlDGNn/gNuwMwhPV4Mvgknp9KPCfg1KtBABcwirz1ouW/w7I9
FUVr9o6WEyH1p/gznqWUTvdc50hBZSyoejDHB5QSr41NncFL9Va2biqBDVeg
xrEjXMIk1kSY/N1qm3A9cf+mWIYUSm7oQWdzVvFPqwH+zvU6Bpd7jvAhBH+0
jjuqgg3NB+6Fa/IcP3Mr6m4JDTARNzr2wqovuz8jUUEhb5IdzP/9qnw3F9ZT
XSv2NtA27cHGy3e5FvC6EAWE6iM65UrEZ7vLvJFKPM0Ktqy5DkM8lLkpIle3
UbzrFtdH4qOSO55DnOj9b4bgUfgL0hzsWRRPAtFmifYZ+AMtp/117/vlSkst
K9Tc1MFu6qqi274ad+XCTnqTk/2+r/9/nXzu/2s2l8S3YSKfEjtwdKPpACAd
ZkspLeqK5nZJSotKp/6gjyqKP3w3+6Fem6bxCV5gMQ8Jk0/zHee1jB8uAnvc
F6yzDqNzOYYIkrBesvI+LGqV+KBSibej0frgPNo0pYpNL7TRPGJOEx7wN14i
e+iuOcqeAh5hWEqxI0Dp2heJO/sgFOGYxbmDPNcI9+cj8wfxeAP2RG4ySQGq
YsZAhLimoIw6B3bLxWNlz2WvFYx+jqidbwc+/1xWgFgJojWRfuzVNhUsF7bX
sT0bj51OPeuK32QT2RkdD6ZwaToEbJVVRJJfQbeIZyvRjtnbXJ8BvwRezm80
OR+cK1wRBfB0v0fhBL7C4lwFJ4QClW3Lkmay8fTpO4TyAuer3D+g9Eqxxwe2
oY6E+Ef99idYSsS++z+ATT7NUYxkZ3ebvfXZB9j3O+7urIYruAGWn9gV8W0S
BHDn577Kg52hzeQCnB4jg4n3rmihNA7CJV5Jaim5b0WnPj+4XbnFJz0iS2xq
LHaUTsyj49UJOBQfjT31FxbAikFpum3T6vHmXUhIIebXr7XzfqPjOA4tF/Sq
qaiUn0UvJWVXd3GAuZFkY+qrs6NfNx3TxUresELytHSsUj5GC2wNNZrj3lRB
jR0P+eQWjP5TmIWvZ+FaYznGIgsWi4EimSNeHZwdCgkw1SoiuXAgn0IMd2R8
+NA4hu7wmNwwJBATr+7DLKb42x3qd0wznr8Ibvy2DpbmAOXFKkPyHFv5+ANw
cRISWoJ+jJ2B03O63nBHyi7am4R6ZYD8icwX0Y6JxfCDmsZP0gZuxf/v9iNc
l3kjtc0VtM3+6AeuWMeTQL4dkqiWIeGI+6Kwkf4giBI8e4jc0dS4S4ghOG7F
Z1dR7kb4knUnmo8Ifay+6HXWT4YH30hMGzx84R9n9UOTZYwrFrYX4HHnuOIp
SKxOt03vTv+yIWGT6cDRlC1LsmOe/ZtCWSxy/biGtjxhSfhkWeeu0m3E7tHc
dmU+gPJLFQEpjsna2bhZt0RtbI/K5MeorVVHLKXWVazAlGB1ghI8VV+a5Uwk
MKdfXI6DxO43jBRlfcdPibXiy7e1WIT6RwOEr41xnH/7YNsjnaZm/ps1N93H
+Fi6jo4nISgPklQh9kYnH06hvaNWNt6gcjb/Pgzr7NzYcwhN9F7E+Y5Vuf2t
JapZX0QnHpolvAhBDE5AWSdab6Tsw+1nLKYa+xSrwxX7tLUuSEhP6771gk/n
ueYibfo62EM2Q5lUy0D5ZCfdDQA9dnMlmwSgpGMULzBLWi7ADHl/SPOarfIf
wWVeuAxOQt26hM8vHqf4cbUgT4UYbpn6mNfq2C87nI4bEDZA655NDiESxREn
57k3NvTdnAYqqkFYaaAz1s0yh0bWkzcqHGABjosm2iMCABt/TtvKnBF8+RQn
mviP6WNpygmnhibxtauQ+H/eHvFKLuoFQ64ooKRcMCK0JIpfXTwrmnTes7kB
qKB+0ujyF9agc0718hXV1DdlquTmDrEy6xeKNvZqgRewLUPMDdnMyGRI3yEf
xUfxQN+sxm/wEuRriPgMsYn7Axgcxy0nNifwcgmBcOgL3X6XsRAl9d8TzsbW
iTChM8klVX7y7XFXoHjiU7Kk+qRTdiIR184TgGvkqRXK82jKjhffTMoM8fpw
AXNzlT+dP0igfCaMgBCK2kt/QtPL894bKtFNUEuK1lSMoBeBvm7AbFP3TMf/
rE+ZXJMaVZGCvymE3eqETySCu2com75y0nU12G3HfgcSYNhvynEUjjRgJgk1
gk5eLev7pJUG0Ss8bMXEyjrB2Q48WyN0YWinMMMninHGsblPhePRPiI6LIfl
5u5oE8k9v+Mcl1nTq8npzPeSnMZgP6FkWu11A2bXTPy1ddO5LB9NamF5Zwpx
CyWX8TYdsjO/yyAtu3riS/cqQCCq2cS0NoBlcEFOll9l6MKuGTNLYJmz7eOi
tRQIcjyoZUL3wbPhEFAXW+XmvN4f532HC3xHUBXlijm8iWxwIUczip+8OeEQ
zyPgjGfSIMj+iMeNmZi2UmNoX6BhF0RrDl/HajGTBNKbGviTMCSKWxzhcRq/
6C0d56CvHBIdWAAvzFNMfrXGbVRAGjXGxcLVcyaDRsWAMmw7nPpfCUrSN4F1
MPlVZcDv9y0Sbo7oWTf9mirSsRhzWHTqr2NElfLgxSteIprRlgz6wgUbnMpy
+mOrAB7ogY4h8D586xWDuvYjSX033vY10zaXpHWC2IMzx7UTqUPixRl6iS9X
ImQIEmP/lWmpM68C8BXJTYSS5jpm4PxwWXRG5EklJAXc85LImTdkRFg3jYE3
MA+S26/ubyQxE/OWNaakOoijqapzmMwB8aOz1dI6273EEqp1TPu05hs1XWEL
/zwX3M5/sAIwzZGbiKuc+xq703x444uC1uD+win9JlrcYcMTrOkoWQ9z73pc
UcuzVkm1EtFp/pmWUIJQqOKj+FzA4Bz0B0Pm3BR3E6SQCj1zch4OfYRG+MLO
NTOAuNxkt4k0e+MfPv4CurTSTmnzNnuV5LdtrHQPUeI4SfrXK+LIACFmuk6+
j9Vc+EQKYQ1HIwA4y+s3wAqdPrZwDVly2sXhA0nRmJd1NHcV7K2yKJ6Xl7Gf
Q8aI+MOE0bKwKtjQa3CZLoLUwT42K5hfZvitKmmEQjOhQEnlqp67YDJB8CBh
RU5nZq366D8XsQiJyNLhkWEK+oLwUI0UBaKYVJ7LvNElIairuDORGmb8CFuQ
R8bfZqEmaHFnRlzb3NwhdbQ1xLEWCIaf1xYq0EoJE4tF4IMEs1trkrgvce3G
aCKREUyhUvDHaZVI3fwk/MlXWR1HEIRIWVCfm77FcPawjMDSr8aBAmbcKsDO
OVZuvpXO+gCWckfMYyEN7rWdWtcIHdoMH+TDmVHxgndPxNYzLCP+jHoRSPZE
kdGf3u0oOx6K8ju57EtvvUXaIo8mc/OyIDVfPZxgrZ6odWa7q2f6UXiynyAX
fXqnqv0/53iMXsvRL5V888eHPU0ypoPLGq7hrJARx/+UX0NmElb7J7euNMG3
AALjK0Q3B35fMfOZ2V+8LNVtk+zYD44vj8/TVSti5uOJpeB9aof+xhgKuCE7
vHhFarmYlbsjQthlbTHweNDTYB/ndZ7aYXzjTO7kJT6o3xG2gpR8o2pZMC5S
azJO8quMoRrrYirAo3Ex8tKGos0/tDkBH4xi6W0WbU5W9gT9CyW3izAgyW5G
WHJg2v/KzvSHv8OxxVr8s1IcmbbCZQHB7zyK9lS3MWHdcgFJ+gAbGRTO2VPM
tvylrOmX1gwqCMdKl65vcKOtM5Zzpp5VALwLKy0wAqzdENgmhOsVq5Tylsf7
Xjc74pb1bnIKlBGEI2fi3Z1tcmVPCOqAtPTGHEJh5Fint0JBkr0MS5weQsDA
VQvCR0kKS8wiTqO6QaSFEhMykzjeSmZVdaOCLa3M1vRUpiRMJLwYi2oBIaZX
qwPN0JMOAekdl0nAo/L4OahfK4WqfEyDkB2qk8CYlq8aFiO9BVscGAWrA2r6
n4UuCVzkvOnNYPfumXuNJArOaOriZwFcNJzlYVe5hrs+8N/EhqtM78Mc+r5u
hFxcm3quOAgGmW/QOsvTn92oFtoHHl+VBAotaXGXJfuykf4EBGoROysEPoQf
pUlNZiJmJcBNTO9rRYIretsA9AowRkW10bWIkfRn2uAkE/p+9/uP5ymRGRR5
Q9q+G2dW2L97KfZVM9zmvzSMH79jB+kPoASWQgEU+pUvSWWz4kZ4/TO1JoQE
gQ+RUi1tbh3HaHOCEVjUBTbnB/woA4cQFOTZqe0QfEBBu7tAHvu+DOcBE0K/
CUw8aTSwcOme7b+YihnPEWPs7sjCz5GB3dWigjHyEP8tTY4rInMMqZmcwhkl
MhdBTzdxmG4ifKKVok5Jl7W2ktvCw2oSNfGzX0OCjhHzcrOy7UOpcPFIhR9y
K9/ccDIS/5BMH/Rbk7s78YH8JdjAXSluA/x1xE9enfqNbX5VHV5AiSMPtMBI
Zx3ypd8Oj3Y6PzuNyi2yq46thH7yRLLpsAPe7LyYUhhUXWBxiKEbxetgg89a
BI8kmwvvgndraGTkCBlDkV6wbmrViWHEI9G1ENVzb6bPGB2OpCoVlF1q6MWf
QFC6rjP029b3hX3u7YtyrJtI/emwpp3EIT397te6XEDKPZKn4hjbHntU3LF5
my/SY+w9r16NRpwS2Wce+eEtN2E6SlMDHD96RhJttw3yLNJzcCm10FggadVN
/AEavEZRY+4/GCdX8fH4byc4vJd4sj443YkiuOf1z4S/MhksyAhx4p8r2rs0
n3bdNPcYr5JCHfFmqBNZkJlG65DB6uDGYmjUhm+sDhHLrarxmf4ZqP5mb79A
Du3jZCcoi+4dP5on6ObskfcdpBaJarfstj0IPUkcGIX6Fn27r3a5xJGsMP3X
qYaB2AJeeQ0UO5VQ73Z69Ekb7PMU/EM8lt6VouUd0ilBNPYzCrBJH8xalOaY
j0ZtTVhzqtui2HBZVYsrIaVfKIciUG5h7GPqxcaaW0BbG36H/rneQM4VJ3HH
bs91Hv4NZfOlz+gyMt+nMPsdxvGEoCuRw9jPOORaR9qlhjGj9h9eu2fCoMkw
qMfS6M/hG92Atmv8iJU9xErHY9Jmwao1uJYEyNEcW6IQlzdecRQBzCsByZ68
V9upPN2leuNO5/PeMEzopYo4vD4kN4Hr+/IzaKBPJ7O7LeD9RXSjhCECADC7
gSeAQHn8bPa9JKEBDoFhjTxQMCy35FSDOne5FhFkLoURf2vOjd830UmpfMeI
JIO3eRPJcbrttk5jJtM5+PNaXQ89uUqGcCqciOxIAsGVsa58NmnvB8djB4oN
Pia7hbH9OZAziklt9d7Cvz5Lm5gb9N+fJBibKNuRCTQxor08w6Hx2P6x5q4B
0G8DIVgOOtOPae2YQz+iOu601UrrRdq3goZvkBWndCb1LtNoBqekpFCmsxPW
tlnL2tAAMpKihpMVT2iQ93RNULwzDzBCKgabPk7vgbgCZ8VXh6Fn2uW79zGo
SLtIj8cY6pwDOJhu8+I2WrU780Di7RX31P+N+2P8J7BxaYeYs6rTuXGcErm5
g6jtN8WQDZ+qlARBP2OcUmg5o9uZ8xPjOaDhRrODDWVKpRGb6OZPp+Q4e2YT
Z+pG+Gd74xO/VciFcDRgfAkWAp1L1c4i6EgFI5b9ljnm5j+OoCa8qEMizn/G
JKyiEWfi7k6/Xk81pwrRNYev3senUlSJE1OWdr4KaEg1fttcJBvD0E3Noy9Q
+Cnbod20+qTkQD3eBMMJuS/omPfMvoxRuS8sc0/qB8IefckbJTxwjR1CpZAB
O/n3OJz4v+Z7GqETXD6plAfN7yUsaSZ4dqDuEKwslGBedBUl4b91ck6xbhlr
9KNQl2ix1WrT5IhpCY2g/5SJXGIoqKCaryD2kAfRvUoZt0cEXtZcbCe4+kVW
rhyi5Et6pnBMnPjThECReh9mhCou3UmL36xdoTkuf4Ci6Mdjn1QJ8PjFLGW1
EX2O86czub5f548isnlVN37FSm26m4ze4JR1e+MJRwCfjZ9fW3WwMzNnmXtX
mcO9ozFbs7SpG5+k+tNhCURzdTZ3r9TXkMEeEsI/L/AWACialK/3kN7Opckd
r2fcA59qp49Y5ch2bPgsdo7PPSB2rkHrFHj8rhk1mXdSE3MPgGYWgTHsrk8s
IaUohmDEyLOdb08C9BR2KT2+jI6jzWgoURQr6mHuRlbjvBtIfQ8/Wir9dSVB
5Xa8h8kHfdhrrYqTRev60En+nEb4gdZCe4g24cgKwe2+CbbEhpKpaK1iTwCZ
VB3Jv/Y0OlJmBntuelllQm/ak1HxZWFnrKfsMXqgOA3GVgRPxDgxfAuoolVw
64JYYgbaNn2uZ/cYbgA2SqeylAEPeCQZ2eoy9LThKwbH4GU4sQMr2gMU6cSd
8KQh5sIb2uk5/F9ejvYTcJZJrm0RAm9h7a/YGYb8F1DSw8C59k6jHNE3Fujh
9BiUjJWECIL74Kd7DgIVNrqiqypRk565aj65cOd1rT/XW/+A7W1x5gd7wB/m
DY3sD9DKNHQn7MBcMjMe64nM2l4ciOXrwSVnqO2rwm8RGNrUrzJq2Bn2zbsf
a12A3tPJBpQ/z80JjrXwpCqkgsetcv/G5WZ9Qx2aEmjqOfZ13Ep6N+xLOhtB
5529b4I6g/HpVC8TH2sGcjnJhnDkHtvZdwQLsu/vT8tx6NzEUFDWSwQeWDou
qWS6hs/Pw2YneTPAS0z6ae8sVMKtCwjGP289Xg1xCOaDKZ9AB5QKi0fE0WHl
nMLrGYphZymjTheesBYvPtn7N8UYcmJDMXGP8h5NW7f2epMx01vkqeaUwTsq
jk56jYm2xzA7y2jR1wLoufuJt+E2tZTj2eDY1MWTggqtc3kKuLn7fTVoKAGF
zjoCEXh36kG9AzK3ZykTpZWChauszlhwfNDUaCuqC85f9T5L0pW+CDNmc3HL
YgaxPVId3Btc3MXm+1ktx9eGpiHJLj0JImyRzOaZRAy/IhJp+z7Z6O3UR5wl
6PwLx5tM7Bf2ccr0a2XNAZtEJDkmOgNjMp8vnMikwW5hgQHhML8cpCgcsa7S
gf1kPsoJFBrVGUdGIGTfPQzngYm9VQk7sWezRVeyGDxTpKXz2l/0QzO6KKii
UF4ruYPOM4UsGO66Pa3JqVnRAgZU+b1MKtxKMntzbS7CSAr8g9vQKdtr9SGz
HgWuH8EIsiD2ZXGZ54pwxAoOlFZrzl2gaziFRgx32s6QH5yOOsAnZGmirxRR
lGat6MNoCU4hnEQnkXTfyAdJ0QwLlcjyXQ5rBnLYGVDU5SuLXDDKt0IlT9LR
6s55a86u5ozaHDoyrxpxFcTT/NBc2B2bp2vRPKMXZFH2VOj9S9oAdFRh1JUa
HKRrZVXRNKqY8Mlh29hgZb9CkjeY23Iwh6WJ6QKYiTRDL6C5jEobEXfc9Iw2
oh4tcD6d99DBsqfVE94nConAXQ76gRPhOAv4DgDLsnIVnWH3Jr1Eaz0DirqB
9TAzlNUyGNCNnTirUKFKbfvup2e+kf+dQjTqy4X0Ov4rE6JdRAlfCWYEX4RZ
DuDNk1U49CHFHsLKU2afblbN1aK1Tdg5kA0BFC82sB9HtreqvNbYy4dcgNsx
8g76PPXegZw6FwkeKmqr2amieMikw80vq6aLTVdlCGO+xWH1bJnXUZsu7jWr
k8S25ZOzf3gqf2JjT50zVpPsmfAysX6zUTsHIN2r0rjDB7vNVUNhEfJLgNNB
P8E0AIn0WoR1rSDR4U/yW5YVNPMRm3mkWBkBbboQgWVekoJBblibD8fIBaSu
tRy57y2jAeCklXHCP5+FRU/7DHohc6xkKfJJwMQcHT+/9gZd/6PP24OmqdPl
o+nEPh2jQpNC0/3v2W5Q4S1kziAUQQy3PpwfIzUG8hVeWobzz3n3OrliieOv
brwUf13HTJZ8uiENXAx8PEYmhlwFfp6PlaLwTx4wzyyEoqo3f16GnYZQZV5T
Rmbjs+UNt9bTqfqX/xg1sLS01rR6ZA4e5nULOPIocT395e/MkhRO/ARD/MEy
HpELsZEguHNQUHfw4cQX60nINah8oagWWKct17kSt7M4JwJZMX5WVwByjP3A
aZy+gJm/WByBXWN47yfCTwpE68wFjKnPhp//mmHZdnwpG4QdwNa7eFYqvqEW
snFOvqBscOK22FrdkhEsxPWFz3shXYH3DSjfGMGTWryeWSgXEBblrvGDBI7o
Pvsu07y3U3//o9DCFrCgWNrX/EuE7UYvsvp7hVh4IiWf1f1eXjf6Hxth9RZu
nxDFHhBSQ4HZyciPBqc4V/BS87OwarZ81X7Z4J0fgT6hhGs5/b/m8YJdADqb
wA/CQMOzXXSVy+z97UlyGoaaLp4M8RDl6C3p+pTQ6F7veBwFJHRixafsLXM8
ltWn3bq/M0BOxjAYqnkG3vV6CFIC5z22O1kcWgU9CspM3dnxAxqFVFnHBj3P
LtYdB4f5ZVByw+TwPK7u17H16Pxipn51eX6VDEOqmwK2GOkDLsiXFoCnajOy
v5LWoOGdeHATD9+XQIzDGpU0u9ksNoPZFr9VDZuUzKjh38v9X6G1yLcl3TFn
5L2I/XiyT8oWpwIwM9ArG65TdI5XdSl1uyO+PxWp/LW9YNkRib5EApnHNMCo
7Rb6+QnYfqIpx4367KFbcRPbc1jnT0Yt/3BBOKJBgxdQjysj+10ebcVDL8y8
pyucbd6fLO+Ub9mxdIRqAjZAzWSR1glLhX1KXtiFCTTK4fImZkHfLsFVecyb
JU5i4K/n/RW7d4X1ZnvfrMLwCyM1G02/LIcC/FxnVzmSm8DtmUhdUL9oeY0u
FnEHa7giBUTkAC7A60ZBeHjKmV8EIoqtFqVl69yhtv/kRCle5G/NuI+ea7YX
VOzkpxrXaKlLgKn7rn/cMcHJvo6aw+Kvh6z1I6wWMcUdwX08CmVvXJGhsCp0
NBnlPX5jVjzFZRQ1XZq+T80EtqImfqFsKmFtNhLMW83MqUsOEz8kMqRAFK8S
Q4lbvUW584mEkuwsNa69rf/yixi/4wLkOtuO2VOCa+MqyyC6HxNt+XPB7iuL
RxvjZoa/HpuAn3Lo/vqO+Qn8/f33g04T33Y7Qri2N170uG3bi8OmXyrvTgtW
GS8ChFTV501zKUKgr18XYP6MMe8Bp+pJxZDpy35qnlstuifs97nHf6oh2bSH
mDH0q491WV7pmZ3DD1mNFO/Fem5oPBTXjTsbHHlxQu2opE3vIghOXZJ/0dMl
PyYBkFv2NKkg2kba2my4BNWC0dAGUxe71TPUf2HgG1iCDje4QvbKel1Jat43
jiiWMIM+P0JvXBYStesgtQhXXMb6/vCHaIB5c75s2Y2zQKAmSwI67GcrVssq
8gDPaP8PTeWUwKGzhYfAKHe2wHwCTlC8rqLGqSj8Q0sNDxBNkQJOGb74dRhF
TGzXkta0aYQwbpnYF8yf1ANkMl0w9SDDBP+eXHDCxkJasYmb9SX/d2p27/dz
HpLIxwgiM+BzmR3tYL+mqOglS9Cdfzd4+VNrFFV0Qyrv2eiFCVbd/iaUlQkN
TgBzhmQ+ewnOCjtds8/u+GQFvpvdPZK52l1RFvprRfXZjVcZtpc3c4dvz7Vk
8IMyYccSo14s3q8LpGdq3o2M1tfLIAwjXcYyWenZ60Ja7lflpskOw6JJ9nBf
QMWtLqTjpMEO+gVD2RRIRN4X3Son70uzDl4CCLb8+cbyYqLEJaG5LXAatPYP
vajAQzj120Hpl4JFsvPrVCFmJ/Ux9VQJaoFDfvUY0O9uZ4oR30i2M00xO+e6
T/vUkeTIOaUeXnIdANtMzt2gcNVk26C4rYRLhXHrPx2cm+dxzTQA8J1YsTkb
xRFH3dht22fl6FcSCYgDnceP0mdx8aaRhDl9goKjjn0Pslz6YuI6dtyXVppq
yeGa9Gq64XeHO7hwDleeoRCNdvkiZjnodzrTy3iGnwfd8LvCCvaG6Ab5UZJK
BRqzU/HUIwZMgbf4r5I2IqSqvrP43SNoFPSy3YRXu/5JaJXc3UdEhbJLqonx
d7MhLKwrYuoGD18tmaZdRdM+XunvSkwdPMxNDyUk1z8Jd7Tj60xMrDymfT+g
dy9ytL5FbQRJv7Bguu7FW1GoSrMpsypuP+phxPxSFL8Wy9O2NMR5eILytsRf
lujhNkIpy2VFsDToWXACnrV7uSKHD6tEjexz4GJZanlntoHAySKC0v144Pp2
AFV63BY9V+1yUXnLf+Lm5DC+ALVaS3ETgsCYTdL0BUm/Rzf0TJvLxqMW8BMb
DCRS2M3ui75YD8LJdnhT0esfmgGe2XYDklR9kJdjGLEUdIsFmVQA5tggzlHF
HpCSce+7pc7ws3L9zv9psd8RG48DIJv9BxcCBL+LVL2JKbI7TJStfYWqjmOI
wJwdWswMrb1lL3UxGMgTC85scMuU6bQVGTeNZuwHAKXJdclYBYuNUhZNSv/k
NBsecl2yjX270OoFGBSEGSlGfW5kPC2v9Oc/IQAVDY3SAOOT/dOxqRZPlwub
Rh8736nPdOXH/WZxSD4IXy3aNbQgie99nVCOM7MJIpQx+ercEd/Bh63Dk/ed
QeQrNRJ8r2wO6PwqbHIDb1m38w9E2LyFznX5kUD5fvysExoZgOrYKTQZ+8j1
dhz8t5GFmtC8tETKDSnerqujMIWqjuHwXigceavOkAQ7Q98I5dVyWzwxcpfz
IUnDzgg9CizFPZdK4nDOLmFXQJw3MtxBatF9q4ilha9iX08bapYaMTYhUuIX
viQpAYG/zD4LpQI9eE4fo1gwdhWYfozUsMad1v7GnDis5oFjeEoXWu7f6Ja9
udTF1hvpms7mQSvG8JtGFjNHfi3JIMzfQyHpwmtLPsxgH5ktwnvwR89qKsai
lv06oI2uNksyVY+53ybD0G3krqh6WIyKRaBotcx47JV3D3re8CW6/QAUc7rE
h/RxXNj6FVCLsHLWkgc6cxE8aaiwsfgXPxb8/uazkwHpQiUikswc3eGQG6dD
3b50r1tlrJR4yvtMRvs/ebKeg/pVvoRJVUhFCHT8wQ5nfvV44ipH0AgezLTd
cxV17ZakFabVZX4XG0aLu8I1ZDkNiEyhInwX/qXKcWZ5S3bwocUCaotqEZ1M
KG88aRv05zkmINEgK2CYlAm9zDsWaBD7sicefk64vdEniR8yx3sNueMr1dCo
7/KIGEMT0TUmFUkFylkn5yKnGftjWi4GYD6P2YdlPAOSBf5S9yRFNLIH+Ff7
PmjwF3jNcNHPq29FxXXOvO2u0itE4sAUE+zDqncb2pyj63bXYN5asqYSLBV4
7s/cJJFT+KrB7eqRlhYWLtd7XBka2J/Ah59Z4SNoLihlUHJUPlbHuEdLrUGj
gSD5WU9GICJogJaxNnaDRlKbTN2FxFranVtbi2mYi1GKBhco9b1gaZ77jDNS
1Hd3ZE7yXy9pyjerRAoVnGJ5Mkjng6cqAIomh6ehdc2NkknoTET8S/Lf8iDk
AcdgcD5JQzHQhHY94KEzPvHlkQQQpaCTc+lFh//CQoDfQGcAtb3W3xG1PwWx
rLYZWWA+CtLyX/0r2xQh/iHdfZ+T4n9ts/5M37bxn0ug8Rg69AVkgVhQplxp
QF1hWsdcmcVE/XKP0sMbNcIjCZi4CutBF2FdTQ7VHe1z8y//b7Rw4/ip+OJb
xG+i8L/1dhIpD15ukVeDjWeuR/QoYlO1tg0wqpdzR+7WeayeV79enSEgR9CZ
3klwJwBqwcPMJ9GYmqABKaFqnAGiaJEwcwXqIkBVF05JbwvUfnjiaT6I7uqC
9nX/ZecnSTEJ0yenM9d8d2PuuU/kxk5UQ85FAjZv5VGhP3t/cyAzWBpZsq6q
BphFoF0jG+mrTynEgVqsNctRWaI883PBzmvrv+Zrk6vkNT++O13A3xAX6yez
U8H6Q//XMu/3rYsrVlBxt4sppduNpSfmzHipCGAQVBMh8B74RUzqmfTShfvn
76ng+5G0otFx3XYxD5PPK3LvdJG8cR/QEEQGytT8zlHzx97DvtDTVa9y1CRG
v31USWzJ0QHiYgYrYmjbJ/6NyheeOv3fGVHHmNIdQKl0UbT+TQxE6RZ+ZBEE
YG/g4N2m7xFzu9tkPmUvb/n4Zx7fsAmiDtu0OjKqA9bm0b+mpJoJTRMfRZvN
8JdSzREG6fKa29PFziTtBz76nutmydCK+4VubQLlM0iH3Ki7K5T9URAsE4X+
z243djmHcOdOQL6r8Sa1rDYlSrRuMu3zvYN7RdzsXj+snXFNtuHHpwQqvdxm
2xeaZjjfd1q2wAvNkuT/RmodnRDki+MrW6JVVqr0v+rUm+PGFVPr3C7mhGUq
U1c01WDNdhEIGrjRfsMo3d4Pi/x7aoqQ6xdOVG2ejYQePOZ9ic5DBwadYIAt
DYFlLugFp0rVtvhCKS9+ltydm8YjsYJIrLrTqSovaGiLAprnogjV53+EUPQe
+qUvJNa9YqV76mSps2CoJO3WvR8xoz4yMmnS+VmKLNWrZlLE76yJ7tg/gqxj
yEgzmLFj0qflotcGjxRRhMdmPg+zN0T9QXuchzPZZjQtsW7lMaUk5u9JJtlO
vySy1exmB7wXvnjjwAtpwX/Q1IcHYkgjjagWW/2hqBWmKxOj3FLmrsdFn2LB
920Wbf4H1aGVSzNKafAf+cQMaH/mLOwrxfKsv2OJBt+AoiNPp8KkWk53+Ycc
cGyJxQHN3NEkh/ZSFvmhdZtjVO7uhNv2NvWLKRytMkp534FxaKel2Vwdxibt
RNuXOaTjMHEoX8eoK56yXg/1jPfJ7ahWkv0ccR1h0EYjE3vAoQVCU/7PMSQ4
qjT4jsW2kTnctuaeWtw8lE8WeFrZKhfNGlxTKJVtKUV+D1/3rVdoxMto/bRi
j4DUcv9gTEkGcIDQK4N34+hGvKJR2zCsvPdicdgcsobYHEYcy1vsn3fNooVT
mw4aDvZkxAl7sHVumdrYrHvjHxbGAUoGwLwoPnK/1P7rD7e3tUF/MLx036bK
lGpfBvHX7R9XlrX0i/chcN7u0P26cGpc1p9WK3tNZnkU04voudXxP9Zn5SmV
pu+8bKc9RusbMscXogdIbn8w1lD9K9mIqS7+7jwfG2D+Bpssp1IxBRdDrvv3
yVcPIVXnxsOB0cg9czCwa5cSQNjRYEHwxrD6mDVyllRJ6Zmp1BSFIRwWbFhp
V8T16IMW4tAwTUoW17ZAVEJJD0LHXgUS4zuRmHu/nK7Bn9XrgrNaa83/wh7t
ARNKAGbtK9czNeBWMUdXcAHXrb1d8UUd18ixPLuOw/vTI4nDgC1Mdf0cN51d
ByroyM4vbNJutORVrbuxjgvTB/agfC6arFu39Y9uBrCA2QSCkUtsTYrlrszv
rPVG8Ib5uSx2F3PBoORdJVja3zRbAuA4CgAep1w5ApsIU+59UNiJb8EcIe8o
wBsNjK7x8dnzeBkFRez7Yo9bGh4UZjnRONH/Ma5LZnI1ZkM6P/e1TQqpGLZB
EMDZf7YCaIeyNQd8DxfTNJINP7jyQg9Wby/ZWVMN6vn9b6FEFz9QPVSP86O/
SH9F7ajDzs24LIsQXkMOdszqj83t2OCmmFS+F7QYMBxwsFBG8MAgIbbGU+LN
UsJepCNKjfrPeHjtZvMOft4zZdWvKt7ERTjXxhF7xFp2jmx50CTSm11Muqn/
/F0iCxM2Y8+Z89PddS6pl2Ax9eCIpgXwId/sliz76Dnaxiy+DUCVO+Xaoyi6
y0cOuisfk22MQaoRBtJDcqloT2lEAUDSZkewnZtc1SlSH8obDIZeFtjjoN3z
CNoVFb5iHUCsg/OWz/RMUwHmJUIz1mmJjmNoC41g4S/29RiUZwxChXqmCPIc
inJBhQYgh7xQ/33LAKc5baFHf5rgjVrLBRhM48OY3OCFjik10Az/pHlX/4+q
cJ8y7s+fZEpG1AWgOpIeamctfK7IZs9pw9eJDuCo8pZUrpMHOsMDJAP3LfwY
WMqc2etiU+02bLNLY/tJIV3cg+ZhjgcD3EBCG3V7gFMQBWjWnNuMnHjQThyx
sMuO+s5lIvYpCgCxVA+YLyIM3V8V+xpKAwcrjc5wXm5fme/pPhXpxoJdYxLv
U1JiAL3LcOA9fz7x5QQzGphnPxKu2ZPYE+nsUrmftBb6VQ7di/0AHLWCNF0r
RtfjZReU9LrQNfa3HhRrsg0ruVZP8E2Fe11e9RfxSO3G8lXmyAXx2v93XE0b
XSckWP5paHgg13b4/YFHJUMC2MSKsl3zv58iHUDvWxPUO8VenQdUvvPRzNVn
ubNXeg6uNmrJl8VjwpbpxecyjYziRUOpppjK70Nv5vvrnT9CHjkfKd/XlPuo
6LjGYFAAZBiQlBVTGmBVTKWei50jCCr0N7kmCxBcH20CBG39wY0LFfILcvzG
gR6JWbgwbXMqHHDUIqBWtT3G6BvR7KS+yyDTsHGf51l9wZGHhU5r1lWlZouA
jIuOnE+ZXJH3A/MLDHnqbmrBU3cfjD0zvqQsErHQa8cVmtyJ2RFO02Xc5G7h
nkaEvm6CCQ2joYenvR5gPbhm14G+qNnEryekIwgYaGmUitRzEXjz4v1VPWxR
/HHuEKi23S7VcO12ozUXQAqJZQTg8wmEtKws9+5OpiitGeEmkvu/DBA8ds1o
kUWu2BPhgA1iRPQ78GkTlBB010Honk09wflnKHrgdwkSlJvwc8SW/+WWbnCh
rKoeJO2GdbSUQ49LkfB1aiksTJIEXJbFBS2StYeJz7pAwl4SDatOczwLwTcN
seJmt6J5QW/G15he0GPplgVUBRb7N8vlHe5E5Q2CuDGrAiN6rG7oMPnYxeiX
/oHa+rFh9ksYkxaSs84z7Rn2udsZDYYP/CVk4LoLOU17FoOrOnCq7I/a/Z3e
KbQ2mimVX1UZru9O+jYn6vaSPvv5IPCIRbQOfPqLP/zKt70LF3xO6NtWPcvp
GuI4NuH3/QbRDbknr1UDfTe6oL8VKGWEiXoRB9vbYEcXa/WdJg4r3KGYrVR6
KNgUGUfNL+DLlsqP3MA9IpOKhKfDIoF/Fd7hfekCD6p9oazBxSTUNJLi2tHI
KiiqmZ5tMSJnX6uCKuuGc/cpbm48vtZtikiyDp4y/B6+05efcEDa8dV/1BaG
DG5cImN4sBxHmgGrwIhlx0c/8l8Q0z8v5ex4FAD3N45US2qblP9Rg9fOS/AO
OeBIMnWjuhQrvp8YvU30N8s1CSlcRVcmFWJ70njKC//1hhKxnRHZarSgqhht
84a8kA29wFqnlK7hz/eiHoQtosJ27cjXjNMypAtkpYC1ffXsGic0z7R4kPZc
L4ZlbMHnNo62651Ay8KZoUG9/suPo21NX42QSC4T00SVRmDELdXoMj6ndbGr
8p4CvLzQyuQu7mOUMnEhQ3rCXMzkUQVZf3biR2meoAHa/wKj/QXSN94vu7IJ
e3ZK4/639xnHU2WPMOu22o/yKvlpqnmDsJRGiZ9BqdTM4dwe5+v3qlRLFdjZ
DLdhusVi7C+aQZ9CgahRvr0/uZOho6mvnZKrcDcErlkJfuVQ6MGw1ggnqnBK
tJZJOI/fXV3F0J6rkpgaxUIcBP347pkS9Fk7lT/g/wNkW4pY6d/Uy0UMZBw7
c6WIaalvgTVm63YwMZX463tgUWN5pGPgExXinBFruw2Hl8OmZPHamH5EL/Q9
+j5UKt7doEs+/fEqm8K3Zw8T+JNNdKsEyUEIm9GBGkUC7O9L3YvQDuoehFCj
DUBF5nOllzVW1afrVgC3Yapd1jplxOzxpVDz1IpfES0y2gSsZb4N02vC6uFj
bSuLRNZngA4ILjB6WcDXUzBhqrEjBDHqt0hLzXhX/bVm/fp1afbJTxI62mOr
bwveOZ2ROOv49BXIyNEWxPnFbM+qg73GE2O4xPfd73CJ5T9qYqTQ17zKt4EJ
cYF9z4us7YkOTMW/+tuSIiQx6MFpQ1jTUmREjdF5u4H16kuoXay3HghQur62
O7aMsd8uttHyfs9esthAYBHWQhnz2Ybx1j2+5HB4y1xdYoJtRLTtXlY7Sw0W
qlu22aA9rsO5UlXaYpuKxveAGL09Q5c/WcvwTZHcfymkgPA231Pevdq/gkSo
mZN6rhvpQyeB/CxoiW8j2oTTnaTHd3RF2puEBljkMu8gomSd4HmMAXNqHa2u
5uj7b7owEsS2rS+yJjoOXGx2+88+/o4sdjTEXvNKB7S+8oLiiSjo3McyRprb
JWftRbgQL8r/ziR4mzWUKv4ooX7SnrGC1YO/gKiA/4qtD6u4jiID++5Fmvuu
QoeLjOqNy8obhKDaQImWZ4OFl7mti/TWAwO9HdEGS/GqOMmA0Ok/EGnkCiTV
duNouM/xNpTHiBYDES3iu5Vbyys3iHihXqv02+tszBX0aQDZzqEkm7BumT1P
k8grvH4k2b6Urz/O2uF1ClfZElWbz2vPp7e26X3DDu+ShWL8DhbXHVzfwdVm
Viw9f00T2berC27lkyk2ataT74F+G8oIGNif3yKpkCw2TFvClNNOl76p4ghh
aY8IxtCErgJdCErCz/EMEzSFyDsvzmqEu0grbVPtqnB6IjxunVASsNXhKVav
pGDpaHNxxrLeHKFINuYPwgeWDtwjO3zVZ6GLgr1qEw2YWBaqTTMT1tsIDRWD
DlihcXDF4ArzxF4C5eKaBWioJl1TGj9QN8B1mVxvzWgw2thZXbHyR3yHfz6q
0PkClIbzkgUfwbMLo1Ibynu7JVdITSVhj2IeqLwPN05d8ytLxD/GZdnj366o
IVl3tdIjObTFxQKJ55EEPe6mYSQpYlUEoDoEysjBnvQfHxTwqqkLxrnXxqqn
tooEa/lz1/SXo6C4pUQKpzCk+PCroICbnsTY8oP3EkGRG6Qa8hAz3I/Yh7zR
B12bvgRQPXjPZyull8WgJ5HqIgHO6ecPwYnh/2h3m7oMwH3ZPmtADfefedaK
l7+kH9CY+ouKYGNvHJ8qbLDDftTKidrkUhsfvpfcMuaFFEYX16HfMpYQ4H0V
man01mzrHOnhEHg+4S6pHRT8OS4t0QXqRIIP565rBWVV2yklMDe23RwHkQnq
8fyUzmgJPMVwNh42Bm+BskDmZSFGGX0mMfl78rHq6DcO4acxiJcyzR97f7/f
49/iGCWOPlwHogTQFUSK9HSF+cS1Xn3D8MSRWfAiG7l9xMb1Zq4pB+RWUbY3
Wz4tI8NsKQTAXKB+W/JgS/SaCEyd1OfHLSh7DwGvlxuFgMkfgnOeczZNc4Ky
I5P9RczoT+ZGt78nIfXgb39B98uPNkE+fO+3blKGdEpvOpTXv3jAOWszfCAg
bOx8YgXRhF7verYJIZmThiV5kOS8oGd6j3E+XPjieAY0VwEaN6jGZ38S5P8o
JcFN4B6mZwk9oANZAffyYs3K+fXPkWBZKeUO4B9UVK0dr4qioWRrBFB61Bzl
4xNP/pd5Q9LxT06kTAjbMQUL4C89Hp/XXc+hrjbvPoQfsL780IL9x03Nl9kS
egFgwNKX9uvc2tKpWJpqFDLWXGvzVeGMNTX/Guh2y5+3FAb+2EONJW/oVLEH
c1aSDBLiVvu9ZzGcJK1HOjUWPFvN+mi+43lOYqe5xTZzJlww5c6m3LPsUHVC
CuAvCMKL+PBfzinxDUImVo6sTcwg5dggFpI5buuWxmjEBFdco9/Xl/S3W9FQ
xEY/qHTTLxOloibPwjCKPIY0ciyYJ2yzhSG+97IrLjZM+Y50jWdGgw/YLCaE
u9RhZFCNtwu/TQIXVJruq+HY96aVwl2ZWlrlivx63L1+0GQdmv1NFZhTMQm+
7Ed7tnbhhEabh+iNhObexlrfdNmDgn54u1ecmTUFgJ0scxpdhJtzdlyv7+sK
hsOdJT0C+ffqU1/57mb3ySTBw3c6IP4sEfVU1fjT/o1zC+oHffaMxWDgO/Dw
4A57OChI3yQVv/tMfjRFtaGhtUIWa7PFlHQdbkTjWvO818eCfRTvhzSajXf4
gqKn6R73us9LzNp+KsQpHu3TfDi8lUoo08sy+WYxOIlsgwTtCDKyqrx+HyNK
+R6av/PYalVykOMnalR9LZpRu13Y7EbS8+2XHaMtyi6pWflx/yMHbyiizBfQ
vBFXSY6ZgnKNJpSXyqYCipmLd6mrL/8bMPHe2rKllX4YOiG/8yGwsftzQFtd
DUTggdLR0rXTVc5ni1IKM7j4p0yqXzsTb4Cd41+GXTxSdeChp8TxClF6EoCq
6Y6+ajbvb+Lz3oo+V7OUoQc52g0Vdej/T7D4zn3dxQUmknMgK1lV0qCn65XA
ojg9TczhDh4wCEdk/vAfUkS1NpCXVRmoqoOLsGbi0LbSCASIq/jFw6aML1qb
8yjydU3SV1xrIWt5HtwzXqrrPA9tAc8B7h6KMA9emNKAtU3E4dylWe1x8dDQ
VY7aU3yrPBNntVYs9q0kbPSWZcHYD2ASritfNoSjx3gwJj0V0XxSNUAYdW/5
UIfyOs7Pe1BwCKNlfQE7EVvlZtPhvpgMwibdhgQbZAXAv7Ck3zXByfVJ4GSf
gMfnSiO3DphL/PXuvfzZGDmj7SpXT/exes951si368O7ZN3BL4lugm29VQ0f
jmQjOz7dIwVqcjsIpvt0dJWPW2OuONARSbIsgwfZyZ+Uv9oGjx7BOgyOSlrh
xbHWj8RMHolZpIv0jYrR2bzuuXKmDs3qUZpqFYd379ckBg6ec3zfJF+ZJIRE
Pprq81DMy6X2VSqPgMvytxro2aFcNo4ZXVZPaGKnZe926QQiiCQ9Ep45qG+H
QNS2UItH6s7SM/0mpNTkbQW62L69vEjcYvvLDTOK0POI0ZjW073jkqeVgORc
88ANKLQm8VxuLrWJNnqkO0K7b0GfIHQHr6X/vVZJh5lwJEXacq8MDYJyXkSz
7DhBOWXi9AVHgLFOq/5cZusZW2WwwjXFFSf+kDH3t4qjP28gmVBeMr/P9v+4
if+2FLklh4P4KRTIWBYtDXtjXqcK5BEeA7ZCK3mS7ooDni/79Vz5DgS/Jvr2
ibPedCulqd1WbEOGMA5ZqB47Sw6Y4W32kg56N86JDAgX5PJKiiKVCvOd35i7
g/oyeK0iA6GrnAPDRRP6BYZw1uqCnT5ivJG3c01L+lNlsVeHjGOaDm4rU2A8
tfEgZEA3JAc98foYG2msgpO4+EHWZJnawXarVk3rfuK0g+sQ/UEzSQ3SR0NG
zvZlhDUUJzBAcR+Os6KvTNRObuEzAeF3TfAnayuIb/BKAQJr10zek6+NczWh
60PEdP42Bo+JeM45s0SAtM2R24PyO23xH4YFL71yUac2SVczLMGYo3kWcbjn
mPwB2HVvpQ3nWWs90JwbVzVNG0nwNYcnCLASHyVKbYkVVDjcFzxL45hqPE9j
s4KD3Sv1g3A059FFRVyty0/IuWcnkGJXJji8GhhOj9I3Fs22ajYrk/it+KQG
PfmKbofUXCPZX1Uv/eIbcOrxWQW2Q6j1eCrV372+op9sfKBPz84qBKsH0wpa
yM/VgA+mLRRQ6QeuoBuu8e7Q8u0h7HC558Tue2jVrzncqAYCvrj/dn2bOzuF
x3gDDtKQlGtYwESBZuSm9FvjaIKY9xrvsXvERjQylepHPvnvOAfS9MK9zCYI
mxjubb8gq8tlyaIr5OFaTHl3yj84EPbsMMOl4NRD7T7P/Hoy4EJpGZ7xPA+S
zqPSNZDtFeIWdj3cvlNB6nN0iQl0/yKqyamyLEMbZ0QVG+Vv0zs7kIIvhTrA
9Hd1maxdRQ7owyL1du7dgYP4vXcvfQaOIzri3+2KypIHdwuvvq8AJJJDg8UL
W09M27yJ5908Yb1S6QHt65K5tLql2ah8kvxTPOctpTYQRffyV9xeJNZQu6Ub
HX7DxBobdBSFgSIaQxZp7TdjgOoqrU/IlY8OOiwO2NSIczhjUFips4EJvM43
TiMb7ydXXfF8+t4btR+VuVuVMfgu2/xd6VpX3qn+2gTnKaCUmj9YvKfV6zjQ
WhDbbXVskdOi8wdVS2SyRp1k7c6ULD6x9HNT9py1JZdxRKmNoGx7suAbEA5n
fTlFltPRr89bwweXFLTHB9Q3Khs6+0dtg3mW9I/el2NLg2offvG5iRGqcSd3
DhcU+duIf4MCI9d9RsuftWC6YffdymCoDCwKGe0HUoyH+uZgDkXhm2SWj/vF
lpCEdnIBfMdmWEGyL8HMaN10ES4TER7yO7H55c14rA4xQADDvGteVBOdnCVj
ji21BniidkLv14CA3Ivv8t354hZqH7PDamlS4p0Ntpn326NiQmucgyGHVcS9
N2x4f9FLLmzPfIVrViQWaVu4ozsQoO1oLOD1UuyVn+0C5LPwz0dN7hoZwGCh
w3nwfJP5fSmFitk0WcQUR/0lf85TpM1M46Qt7Y6A196Coc/xRPyDeNPSN5Kl
OYAOcNntbuWxGvwVuHSZVhRhQ2YhT3uj4zPU14V+pXwT39JlshEaVV0t/q3j
fmRYROQxXrgBVfG1quA2pRKZMiWffzy90Ilj7Sf9xA23Jq3M0bzE+isxzc7Z
Rk1povPDtfWs3rmSn5DJgPYwrKh8ySLfd3Mn9TiL9a+UAMhdwCi7m/Q+7Tu5
kNNgC1Z5qZRKw1XfTmyY9rBqaxerHIGQBkuu/Q9ckaN/uQlwP7dL/rbF5hkO
Rw/rXFeSvG8rhNfbB4os3Q00hYMKfIQsTp1/lsh9A8n62gZlIOQ0QiOAEM0v
/1gkJCDYgHKj72F78jk1EncFVEpskwEMOXxnL2EY7bBMidYkiWAmOUTR913s
maSHN9OcXDyc/9EFI8ky1VbP7vhVhw/p2cdy2oMA0jhtC/4o3QkWorfNw0cS
7cm0HBmnKONNMs8/odsMFdyaXKP3nS7t8WC/Z/KevyMrNnvX6GDq8ygVybKZ
Jl/siFT9un+HRz2sU7XoI34Sp5bb7W2BycLy735/csH/0H0zwzM8P5XETNpO
2HQwOdR9KAvKPvb56evQlgMLKVKTwLnOCm+SSr3iLWEp+9n2TkhM4/20DAu9
WPMFkxu/P+aBeyNroPgjvMIBW1+s6lgoJaE+t8TcGYlGt1eMkA/JJstz1uvo
eoDpfL78D3V813sImGMoVrUI73k6W6YBXFrScM7s3avLvtpJeX6bLc2I6Dws
PWsuUwlULyHLPY7c2ermAx8g9oSWnduzFMzL0iAWSHta2IcR2zIJznW7xnb+
8hzSQq6n2keWlzq7kQEEEyGjsxjLrvraUrNzGOz2c4f9y+oNeTBbf//TKu4q
g/JF0NpM9xWUpSYL6d3KXIjLKwOJynI0pPAOki3txiMvAEHLZoZGpgCexfoS
KOzLoRwI3lYUz1lNjS/DmZaCUg1LiYkF5+aArBqi2rFjIRMzrlztjgcTn1hS
bnlganYSMjmy1gjbOdGeFIm70RoFItLq7RQ/88R+6pThyy3qRkqEqWiy6Q5m
Z9ALQi23JTn5v5BAt2ML68aTJdS+EJUGqhGQyZvmmadeQOv/Aee9F4sLGhQR
Jzy/iikJoUbRK8Fv2CcEkyRo6V6FC4szTwdLkW2h67qPYsw71YJCJrG9wqU+
BEBO+MuOEjUUjgNKs8GL7oVzcg9e2TvPp4SbHLOBMlfNgx/CIg5zy+3ChX3Q
AL7bviyosWtruU3BR9JwjTTmWrDtqbWMgWhv/zagZvLriWmtvfWxOeqJ6KsG
y0v6I7qZldgFnAgEgvWvUt4KgogRB3mGejWKmIQpuSNwxSJ0EujfbtgG8COV
vjgeG7Ox0ck5dQ0ZFIr6YZNxWUwQDQiLftdrGSTsGLBrekPtCy4sJ+d4bU/i
P1e++WVu2BgogGczhmVOyqcqojRzQZO79joZI3vQ8emTe4jLCd3bvzc7Xc0M
orlWRJvIOyPOLwnia8Wbpewo43JswhXtZjMZdoZIdwvv19VZXs1adU7gbOGJ
QvF9OFQEAioCrPpW63EBbN1Oj+mwJXRecPR8RM4qy8mN60aAg/26WG21nBcK
Z+BsFftHKR5yRr5xxu4MGBbdjHAdTV4izNHqKMp95qH1wZ8eMkz81+wohKw2
hec3depTQXXt7glVngTWZtIYKOQbu0LIGH/TK5W+xWe8Ckns4qOWOegDs6gb
T4ktsrV97lQGc8A6SpkxqYJZgjyCk/H8IOqFMsZWI0ul0I+ExSN+E/v4QQHJ
TkngO7zYbTpLDi3aQ2OqbYZnJqhv1JasQaxANXI/t6UmNDDOVUZs2xj+n0dN
0IBtIkfH7UxtIj9plc9KCghZNthgwgd0rpK+hrlIc2EKKnGMJZyrTist2Mqv
H1hBYX1uXiJoqPUjdzUVCU9h3mkiRgR9Lp/npU3xZlH6F30cLmKotv+dvBpr
vx1pbLdbpcpzQ3E+EFxoWo8lJ6+/2zE3IOmaiLVj1erBd5ZWogKfv5evtwTD
Ivs2QSyC53fp41s/Q9XXJ9Qr0ViqFV4WR+CS19RIMz93DNelkAw/fXIXot3D
naDD4xh26Ei2Tg5EZfzhRoxkVf/DoB3SHhD2CbwTZ36EJO0ZCfpUTpUqdiRg
Kchmwg7JjWNFMdSkp7rbvDmsjjcjnl0ymH9oyKtud1ybrpRmwn2mG6k8LlAG
rnc4goXFWIwuOTh9iCacyi6EXcuMWNSI9iDrD4/CnvGHVRQ6zf4xCXzEChC4
vYipFBxCvRBKWOHCGY/8MOh+uSZhtonpZLgiuXNb6em5Lrc9bxbh3uFOWyev
S/6RI7VBAQf0Ue0sC9VobntWi8r3iVk0iJqM1fKxWFXktmHfI2xLxkIkDY4q
6ZUDBT0zOoL97DjjMDZdDxeTNXWvv6hVnHvlnFubOzzwRcgO5OuvV6dqLJxw
rMzs+EmCTYBgZiglB3b7cM6BjNJW+KfuDUo5/U3+sV8rwXP+hhDbc2vsXT5k
TzqaSqU8CYNHnmy6CrlszzqOPcEYzIXNK7KhvMxAr+QrsGJAiKPyiir/YOcC
GX9hOikOunM6xaILLpkahHLtQPPbM+aU30QaYKvAcLNUitucM+vyCWupfSxW
maUwpfgILHKXbhTGFO1+dBHYrf4biMjMpL5yYD32WTDE+umHKBIaewoxYM2L
9HQ1cX6LiOCj0dipTj1LmBN8SsloqSsylPSf7xF63K2Q7BIUpuTRuUnkwaUk
/3h2PRYkUHO4eKwjBHhVZ9lmJ3bbqLqRHGc5n2AIQKcoavaa1ULKkuicf+I9
URBLTFntSXmojqeNf/HZElz4EMSK75qTd0o7lxEp8OWSl2MBkutx0edOIjDG
RnJJO37k6puPEUB5d7hYJq7f2RgmdB4NeHnuTdYwMt6ADxAsWy7IwzLk1bO7
wdsWgiA3S2RR3vm5FzVdHgrPNZzXVZxwT54GjzkmhT1e/TIp8ahV/hVQNoCq
V/rLL80B/zlZu1GoFu0SvHCiRQRP2JJ1W0DA2FUGuAfLvDUSFZSaer4EuGxz
7iZZzRCnkCGgfPnMhEu+hbwI5bSVqi4rYzgihhLybHRGuMCxRizHcnre/BCL
TTaJv05u42Os6Ra+9XV1p1h9y5wvz7TkxKJRKcl/krTbz5HLO5yrByvF6Ckb
JkOl3tmxrqKQaPvLtQnrKdJphRSdgJoU7ZO1bymQJ+VaEluuBvzshXe3ICfF
4UeJI7sYEbUUJaIBdCyyV65wtR0qC8LUjSGhnAsFxrJknN031Fn+WkN2ZAf4
bLAXbvaK2X3aeJxFts2VZZlQRxD8qjKDccVyyexis3fsnlAZkSg5bC6jJyjA
gA6H9JB0Hmridd6xy64UNmJenyNVmsaMZr+AgTCxjvJ+EZD9amCHlfjSUVum
a+9x7ZxjmTGjEmlw7gNJMfaTxThSNlTla1MSCaYvKb904sIxQ1nkvlURfRmB
sn60jc48KX/jg5BcBAI/DZY5peGMF8WQ7rINlwDx7emBjWujIWtcY/MA9iIE
ncJ00DbLaiwhuqH13g995nH+PPn6mldXbn45E3VzRFHZmFoPPgJusoaT1XI0
vXuPjKLyWBPvn3r2CQcDgM7D6WHBOpmyyiHael3bRORfPcMTaX30R3FE0eh0
tGpbrWIbMcxVIZvBcbbteOEmFRr8HNDHlmcz8Mvq3HhxuujMy8EO1h9zf9AK
K3+1UVWYXtuW44bK2xdIUa4K37XdZy8LyU+g0R9/3LbgDvFFJctsiXVslSpO
Jtsnt4tYMgIEtGZti+RkspfAlobha6MbZJvoOAzGTvpYdAo8uzb2fhSD1YWX
smhGUbmafdP6lnCz4WyYaTtSGIC+JTqa601+0U8LE8LYP/oLIfIidmBAOcbv
gwRqhxWvf6rsRRCuAlaVo8XxfxdNQMSm3HtA8B2IM+SZKB3wgdi9Zp3aYKGM
U1q1IAhfQ0EZKgILu6/DZInPHFQfHb5fLkHwmD6W2aBZ/PTUFlkXDj+I6JX2
c9sCuGwG+iFaV2m0fY8H4o3TCQMytogPdcyUzg7q+eEDX0icoQamHHBQTQCZ
mYMPSoNiTz5+KIbQrzqKrGqrC8u4hv7ii9VLsM0by+XpMrmWe7EmcT4W7xtB
V1u0N0SAwc8x87Hmb7R4a/iwJwda7RT1JMhzPwvp1yZZQN4EV0BsRxv8jfek
N7C7fbz9UAn/Q6Oie+rWVPSKrEVPcEuU9tHLsVCjfYgnJAg0H2BR3/D1uE8y
F+fuhGNqGmL+TaXlrDLy/KKI1LfGVYWzoBxFAV9OBsM0JhWHocnB3N8sjsRK
PG9SsVXqGmCkIXmxO8nMYup3/f/LiM/ZDzYflR0AjwXAPjvOIiCPdIuMCJ54
q+xXHNOQ51NRQod58qrXQWGYrBD4Dci91E4hk/PxcLeakAdhUxalaFG+reMa
apu65u/j5QcyYzcqkPJ+EjulBL5YnIK0rblqcbtznwRQZentFA2/Mjvf0O6D
tu87g/kJTiTQd85EfOZ6GjH2lK+UtuiihbifZwHk+/Tk4YDSIwrjn9QvdetW
pXajjkr1ai/PsyPts23hC/DV0y9RIXpkWCrRk4g+1XmvyBgghqHmS4xCFexE
jB5FZGaEiJUAHyD+mPYxLTHOic0pI7wJRK8N4RR/fFDEpid4g2saMCW0B3zQ
TtCD8Eq24lMg7euJK0jSUAZcdmI7Pi7SvwkS6mK4Z8Gf/KiB9PwdFiep708u
Ec3ieU9qa9xGlAmdBjeICdIqogLdk0H1z3zn9JG1GR+Y8PlrMqk1hJyCPFbq
hT+LB3bRf3v+3+wID0FwegYErVuxoztrWoL5z+idrgplzzEnjdYDbDGfOrGd
Ogcp8fJP24SZBUv4hBfzR9oOE8k/aQ25WyKiX5mlcNB/D9sQBhvmVx2RjLFc
S4YBOHVj3WwThYXA0LELEQkaZJhrsQDaoaS/ulS/BW8jPuEZnYTDkiYDfzxA
7kLFOxldQQfaaWXzlnBQjO+gCcKfhXCiSyP+vrof42s4UmDoG+SmPJNFNAOW
KwcB8UusFzwe2JaqKAWJkdSoUIFGsy9ZMdFUDiv6DTGvYOuUdlq7vqoM9OXH
jhWbMxTSoj1Y1rFcyEp3ydJzaGCrf9acF9iJVAkw1kQMjl+32YkvSSyYPW+r
BCPc7kTYVFLOYjrOIpWapqH9Ga+nAdtVKXuXYu+b2/8zlO6VlO8bz6FoJ6iJ
1hkg0UlkAnrm1ATmrIpWtKbEYNDWsviCaHU2GFL34lPfCo4Pjofyd0ra0IlH
EyL5BeRf77z3wy33dPhcSUB8c5ZGJwu/jcHl1d0zsHK6UJz/pQqgSiOeb92h
s2WNwd42LSMD2Do3EQ1XpHLk9k+xLM6GyjO70qcQsr+cSUf4CmRhJIoMM75b
nbcfjyYbVD42ffEI2Dpz46tHYWirk0SvzqlB7BiK8LQ6ZQGWmQuUqYLcdbs5
Ph68igoQjAzIJkLhPECluTsZDYdiLeswljgh31Mu3h4mC0XruVckmQprIYm5
7XjsrNmWvtegYmBLGRiEYd+wVj30TRWNaRD53ZzzxJH36QMGxjNR2mxQ1qXm
gX3ZpBPGOscDNJpyFJ0X/53zb+MSnmbKWgrpAllhNUStDC8MgyFS1xMoDjBL
mJGxva7U+v4/P0RSDsoC4lqJ4jbsdr7KKV6kGOuzZT8w+J0sxoFUE1diNBrc
XzFpYApujr5Ppf0irymOk4qYGRjI5bYCy/NQjULEVuYoO4qI53lWrfI4FR5I
4r17symKl++MWv1PJH1mGkKCZAGtaojyvswXbO/w4cEIwQln6a/ZRqSrjZXu
UgwdfK1LsEMhNpf+zM2oZT2EUq9RTmsXrebMQAA/RUJiTXlOTyMp2xjB/YUt
ZBOYtFzF3mh3YHUFe3yMZCjimsRpojr7F+rEhPd5SLwXAUQMJUZyHFy8K6Iv
Cuuzfn/GWQ8uCKsTj5Nq51jEUN+DMNjGWintvLZNCgDb9S6BB5HQ0PtRtzL+
8lyheopO0O7oNkzfYo2m47wfMatQs4KgaHu4+J7kzbh49DUKdXYSkMy0F8lX
EYx4cI43GPl+ZtiPaVJvm2XUCRFGcSWT3Oy2wZN1+mx1FRSmoyLNEWuvYuUc
kGKoDL18PXQOu2u010EWNB1RYnysByFN2hU14LP2XjCACZt0d6NckrBMFDvH
QpGF9KYITDt/I+PodP+pGbTTIzqd1EgJwd/q30WD8K7gvfjkhRfdMxmy1obH
HyMtdhYV8+pVVWVcIDsAz2GEtxfAupuSQ++bZ5ZNjun6karrSGI6fF0vPVBz
/Kifty0p53Uc6MBb1KBbRUDoaXtYbcHG5GIpSd+j/zOM9MzJhR4EVcRkTgw0
5oX6FFlb441ZSUvoDz4TL+JEBe1eAcLvw9tZW5wIZol9UkRdtx1wWW2G5FhS
OZkb4MvEhYZOTLkaOiB+l37HX5h/VEPFxGcU5MFfKMYKyhyG5ly8JJdFYMIW
GFIQ4kiOl+zrxoxsRASwa+Ta0B/autFLMOc2rvf9NeDwoFjzhpEzcIAERzkj
8QWViyHU9kJWEmoqyGP1BqjQtFqdAuLZnUTEL9LHqxkvU7HNuMmi2htwAJTM
oVfSQWP+Ehthe+30G7lu4V7y818OCmkbNQD16i9fu2wEzFn6UycP09G6FEQP
+F5gTlfpn5boPpESVig7Qcdr+1M3+sTuLPBc809cfcRYKDYeRYb9Id6G1HPw
OXoomcvymGHsEAcSyHx1Z2SF7QQW2UPGyMj4fVniJcwzqI+z0tGkGpOfsdBr
y+9iNThUNy5tnLgoxH2e4NnC1+Cn4QM0g6eN7NrbYKeZTprEckNo94pVVE+g
Uy5Bz/UXmOtIRlTjDbAKJ5rUgJ5AraTFYtxZIawXpQSaXv/wUppGxAB5SsKE
0Cs9E+KzAwkuaM20nXM7S6XCN7TmCxGDzoYyeXNvvQ6OBeDOIk74BUxQMMVh
vqah4hjWrIo1ouhBh/67atEa4zqcVZ/bW8ZDDCQjQVZZWD3EGfY1hhoslh+h
/sWzP8an9g70o8utyUpIfWwvFAYAetLThUHwzaglnEiZEyAvnRbpjQWeUby1
LCvHuavoqm02P/pYZD5Yvxefo1rUTrZAdDu3teS2pnJi4WMcLO2KOADBRqLA
ZM+iM2P3YaJ/LGlf0sZ/9JM7oLoZ75MJ7bu7ehp/ccDOfONYYxELfXJDvUNE
J6rKLj1M87OTaGFJFOeF93kFCIbL8J0sWt1mlgN/WpoMD+tuPyeEUPAjxg3I
aTscRnKPlPaC75y2w9qofD5HJNbibdvQ8SVvDzLK300ITq/tNF3Tj3x24D6p
bvREfs+YzikpUePKgtxCIFQ1hOGYidpNnF8uZ3jsOGu1ORS7dRRreVkYbRJS
YB5X55/42d3MZWLf994hbluCvKDyvUqJomkIvSNni20pR5yRk3N1P9LYxAUp
uyy7OIPOQ7btzTmgowtVShykcmQAOdFHJ/Ue1NzJPslNZohVpWxbCFgmIJBb
im0kviASa5YbD/6fxGIOdZ2UctAmqCmhFj2dagew8jf2zMD3RCUoykLv2jqL
ELSOnFJuVTipwSaL5HvUCvhdAjB/cnYVLvZBG3ieUfarQjKvwYQXhSMw0qAw
kWh7sOJWZ5/nUCxBLd6fn5sf/n7AUM5p304iL8970V07z0s9SukntiUavMua
OCS8PRkVlPgX6dGZRwXENJ5JY7csBxn/4CeatvRohqykR4IphPSd6T9iU0OE
BGmof6EXKdjAzmlSPi4x8RLhGK0GGUVHRTgV3FVbYyLTExv7SGXZXtdCij+h
aWqhcOjXXVUO7yDHtQcHj3t5hAOGxp6BpG6sWvkn3b5AlPC8oq1wN04kRx8B
98CK5/NLmQXfV4DOjxm5bTxS/FuVnut9ergfLsflLlQ3x1IANoXpgXZvZ5qd
HeJcw00dtDxb6Dri4eoO5/SSRHoTrOSGgIHw6LLtdcH+xeTGAqh73P2Bm1RM
byMODtM0y/TTrBU5aexoaDd5XPX5epRV04TW2nZDzmOyapgDgZwEnIw5cJTE
1oCCYpFU2r3xSgz6aafnDNHYtJAX3wumrxifPHY4yTAsvToGlm13abzW3jnc
JoHeYDiWqVT4K3uOKYZxc5c6190A0DNA8Z/oVnENi90h+8Y96nRmHmpHYfCJ
qowPoKtdvbOVdEtYadki1jYLTJwEFbugsid8QSdsdqDw59uX2xQnZJMSRyhh
FfwNRtKPoyMEE+XBZSvwdf9mCbAAV1uwS2bp8/TyDaiEOGcfB4vCWAXgzjfR
WWggVIhjp9vhomVJM9p9pYHwwHmXYCc1CtotgpnrE+EjVAvC+8sKilgBUGsD
dxKh3TXcIIe4JPTef0KNB8fDAXTaqoWvARVSpnpyCqNbiQSRiUCsrPWpv0hL
pdPleQFwIjPxsfpLSw4wJomUJP5wBq3nBFkd/jMW36zh5q/JWrrXMjrVDxof
XvSZRsiIaTxsZgLHXaucVsYlZ7LahJ9051CM703Azmmw4gZm/yqVOpxjSczd
G0T9rANEaE4XgSaBlUIq7OXE8yAOhiWD5XD6mBrWrHGU48AAoDJm7U6lRNyd
RmIQXdt6/ktUSDM2rksDmmLeGReDXxfOsSvTb/fI1sFBcPSPk7EFGCe14gpa
w4ykm8PNkNK/DndC/RTynAFNqws0jaHdUXHLku0BPsFF34mcYoePuKf47FqX
cLfrk7fLFJYNgx5mpzkQw17COZFuIb8PO5wtNT1S7TOzMee2cUzEM+aqFk0G
OGuZDlX1cecmTs0G1Y4Gylp7aR7laof4hNZi3NzB6mG/qn4Pfa/SpCw75XxV
DUvTxrMnIk//Fnr5aOlmvraPwaIcC2DBWMcmNSjyCEoNKKwSNxQ8Sy9f/idB
I39T2lpGmcZkACPh5jYj2NwRegu9JV1k33UUlOjMUYN7R8kg17GJesCIMWWj
2uPAZiuRzZPhXW76J3qITUf3qBylFhdVbQqJujrIPyc1aJLejfpMri2k9WRM
cCBHZ7Z//7BsZAqTKfWRDbk6SqMozDqBuk58707vEI68rP+1iVyCtmLJGgZ/
R67CzGeJ1TK+xV56bvOqWxNWGM+Z7Onp5zuYPR0BefgnvhZWemJMsIzhrxcq
ugBu6kxder9MVeYSzRvA7rI2hYVb8q5f1PvDGzkfpgKTM8gd0k2Qm1x0j2kr
Xvvy71t8irvQEu/kNJNP7GScj8t5B+BrArKHy49VUQp/RpM4fEAHbz/hn1gD
WHt7CqwIiobHYQOYqbvhDah40KDli8O7RLSBiy9jHxsxq4af8qCahrBmBKDJ
FbsEIoTjST68K/nxMLAuRNbX0jupvHGK9WtWZF6RkVQ4qRLm4nTNAg81Z474
2v3y36RpQxOjjsZNfbqjbo24zkuSkfPZxIZmrdjOQMRoQbdVcxCpeaedCIhu
4xHNA75D1sAQZd3yFkzrFQ+7VfBZeQAugKi1DMS/amy08r/MDut7gDfUO35U
GqfZweWRvQ0dQ3EkIeQwNEj3hZSnUSXd5YSn3mzP/ksjW6+sU6BHMtr/aMvF
1k+svLCOmHF1pqHJkLSP+6mYyEoDPRjuO645mPyamZrKFr3hX4YZdy3hSLhx
89igKbbw4CzXk4LI9zOVKMxFOi4F3w4RYJRUrozKn6n2nTU7Ae19yMpVurT8
5bSpZkFRduCLnpf295SWZc3lbnrRMbHyU2I3cn/NNIQUdNYQWTZdsda0zwld
g9GI9q/QgIEsB+NcXkO6to1FRt97zDv4Q1sGSp6fFq41ao1bA1ic7/eiwXAa
NtGpSz/LqZeDemHO129k4nEZXAT6Sm97DKrtyGqJaJmuq8EMxEMQ90XvzSl6
Q6hK8SY0jcuIrfP8Zycio+dNDreuXvALguaR70UYEh+Mmn9NLA/q44PCojtO
qVFXdjKDLtff/HxLOiMK2JQWEi/E6NoQOrVRiGGQK/rwSJCQ8VFe6Sx5Zf5o
Z+mCDANLuabEaUDi/ycRYS3YfxAlngfEbNTGQg/4a35XBIUypXhB+cU8Zx+e
+opF5953oGDrbTCX8qCynhGcArnSRuaNTG5s+yvHK2Uvjuj+gfj/Lz/DcOsN
I208bisX88hgO0X/rOGRfrIIf+aJJk8DsIQ34ZQKYTNQnpw9ys2x+K/ZXKC7
Nk1sVMvR2RL/vQaWDQ5dGWDIYdbhEOrCpPGVWmO5Csxevmv4kxfuStA0BsWN
V09fPGj9A4qlcE9Ao5mzCVTaskS+EaVB5QzSyn9ZqPGTxhBdpYvHDlvN3sab
25Ozgy3mGb2nalfmC5sjSR9X0/Dm+XWW7WQYqbgIowkJ/q7X3LXc/d5yh+re
lVE1VWgesqqnwAyuSpSq4qfBlmGDUIzbvOIwJA8wFbcBHLZf9PNty+lTSlAf
AZQg49o5mnALcVPy8f8p9EBHaKJHNTpifYeiMzmKMVMRBJCthmPNOYM7OPzP
pL3kCzNGGxupZoOku7SZ/YCKddNenalWyP3OE83Ni17ntoQ6fOKpt4vabPCU
keLtrAP0fzpzwVM62XBOkfkD6CWH7DCgmGp6Ex/BlT4kYQJrAFn/LV7xH+Iz
QlqWNVMNpHdR5SLZXLm8w0XAumayidvpfnvGDp1XBOQoWNgS+tlag+NdCUcz
dLJmW1VbzR5tNs0tyQTx+WZ/sqxCRIJQbMH+kZ63C87q2SmQ70XDYW8e3A/W
SgwgriDCYsbsc1irMK2cHuzO7Fq0gr06DWGE2K0mVwb9eVWsE5LM8ZYJV8vC
cqOhwmKvPQpJlAwQIzraVXOPlCJCHRbSaooyWiTgx3JPd+qBIPYXVAXAG/0F
nkbmXt4JIm6N4Y0zbO5KCdWtnbcyuVLk4DVXIHNuPSm5QSkfOPyKeMbx2tFz
nmXcuhWevXbpjyP+XNI/tsbSW/1lZaYqhnnlzxnr/N2EWKcmFi7p4XjeiLQy
jhB8GtaDJezWlNe5qbjO/Isb4kgzKxrVah2Z8971wstNG7Gtag0kE/SQ0Rvl
FtIL1QSH1Ia/sl88G/rD+lymNNCxvbpGF+oJafCnpuh5fbF7Zo0lwKpZCfOe
e4gYB0R6o+4SCmqGYx/MiIJmbRJofrOurHkwcberuR7/37HxZkppKp9b5iDY
KLKdpNO8ZOyjneh6MuE0og+cA/AkzPJUsbqJYPa8fpYd0t4iOMaM9FiufAwg
Efm0W3Wp5U9VC1rBQdNn8oD8ZJNpsTcASSVZeZedvupZRhKpYkc+FDiuMoJh
m7hBi5HW9YT/UOGvFLrNX0ItfhPZgpJliw2u7XBQqBwm1wbYusjCkmcFDLL+
yQ6+YNGdX51rxiBRU1436h0mWHXLQ5h7fYKSs8vyTPaBIrmy/cEr96tye3ti
ySm8XncJNy62fogXvelG1V4iD9FOQmMXtbHuWHsMec8NCGsIaEqqg3Qc7NGG
OWQiqZhvfdX3lqPr1w6CZ3YmhjLT4U7FRERw+ktnoBrLpRSm/WL8k8nv3Umh
Qm10L1o45ixevDFW79hj+4MI3E6B8BXSBqLrRknEl62z4jluSTBl48i8mmQb
cEqWZY3IFKCaZ9wrtK51GZ8543p0fXpJ4W1ONxJ32dQVsO0Fygo+Pt2JR6UA
oxWfZpYBF0bsUhnYt5soEFUWyBenwnUtygyJyDrfIdX2BLo7yEZ9IuVJX4bI
Cx1B0SrdjuME1uasajD08O97UAh2bB/dwMgdT3BEdYqQ/3J5gDN3ziG5uK6M
d5LxKzT8slazLG9/jF6K/Rd9Q39bA6a/8aYAhShSHDKX8FB7FZYoVTJF6TtS
4Zn6jGGlFi1veYMPUf9oPX+DiOIOQee3bCaBmQeMht7AEC/HVhJvHuZhAtG6
cG6pbxG6MoT9G6Ly3iOOX/Av1J5fF6uJBXnBYr3yO9HeY7Cy0eNmn9HjQkDQ
VyWFouk0uXeqj1e5bUfYK4iIr5aMXGq8LTuXw8Dh6I/KaevYsQ81P4nO9lJ3
SzTOuL5nP8+gqEXEcUAnVdnI79DmwD1AiZ76VkmrQc84Nxda24IT2Ko5fL7D
LVl+VkIYMJVr0w2gBEpLT3C7BMavh3s8xJdipDocwWItfbceKXcgc8kaUU+Y
Lhla8PuuqS7sbgLLLS2NXJCCnFk+Jc1QuhuMSKpjiEnS7GHuI0zgbfyGSFtV
BMH/6zPEu+IA7jUIPoztjwLkJdZcflGOebdQW+xO8SGnk57OHBez8ZaD3Nel
Bnh9uEsFsmXjPEXrDin6eB9f0+KhMU8fHi8gKQkr6l4s5jXjWpW6U8qV0l/a
wNiZnc+RAfUsB+h/yYYl4GtxIv6CU9+Z7VcTtXIoMAdYoFBDvop44R7/UgIQ
7ygawNohv/aNeH6EmAjjAVVHjEwb0q8Zop6cGaRPWpbQ862rqHsoxhrpkaBK
plNMSdn+d4i/r4CpdjvbynTzyjk12ZG/5LMljN8sJcKXA//OpLXa6efQ4Cm/
ykQs5GS8vh97QamzkU1+n5bEPYT2IVFSb8dvKO8e+3NP45bqXcrkV+R4J4h0
qFC0rBSdf22MkiHdAQ5AcqXDH01PdeL/csdxVObe/B35TGteLlDHmrXzhw6p
Oy6s5sJ77JnZsjM5hDjKCioYKcCOAvaFshVRkQGfCOkMPhNBA4/WXvBsD5PT
L9cFBB9K0QtIV03XxOriYdst02PFfgBvUlVww5W79hFNWrCN4Pf1Goyl3fBK
nsBFNwyHmieTfJq2rQNOK8pi4EoSG/xs5UKeXsa5rbvN6iZPRL8DNiHL38Yl
gsG2aDvBtjsTYISzKh8uF4Kc8R/bQjvDJDFFxA42qPsGkmCTZTumbeMMVm8e
+GhRmAwx6fVLQ2zDycRL7CLgGm7d4iRwnWLXrLG+zjoBEpthlBNbJEbZwk2f
QgqqmQi9idTBQkQe4GZNmKHeUrNIcZsDiZVPGy+C6LKh+JgQMNqiymbUU5UN
EbBB2dOtxcOwtbQplG7uv5krN9WXfZRZCV/JuD8FeHlvEmLsNX9lUczjFXpk
9/Y25Z7cmKTPuSTvUxWeQPesmtch3DJnfGb2+7gHWQ5I3bDWlg0rfbEqneLo
33k5kP4sfQ4uWBnUGnSn3hqjDZFzsv5jI8sVXSyTz6ZSR0O0WBQ+GF/qTDwB
csRcqrCkivzzaNTAGFhayew1Rfv9IRNuWy54+4Bxo6/EL9gRtAlslrCA6vWV
xKA++4wF5uYe4OcIwnDg3m1ZPuzGQ1VU2kI3TKsZZqmKFRePBo8OW0aMdllB
mzd18FQfhxu4oOraChD8aHZRGXMCjjOFUtBAMDYkoupqYW1cDchvPv2LCr7H
7BS1kcfFmmVaFopEUwFODWWfjy3WW/c2DYfOPLM79BZJSiDdpfL3+OttaKbH
4mJARsBXuOgEGxR08bxEfiNdZFrr04RmMY4bD/iQw5kO/hdsHkQrU4jRl+kC
+G6+NZRESU5GyDVxPxdP7eVViU5cEzzGV3m6Mkpdb3JQtCogjgUtJdgopO/t
kBBcADHVuJL6LT7tIu6nn4CqWBs4rMRVKT75nE/vzP7Om4/nG9eoCca/C3mm
UHnbAuAUuu3Oz4C7eU4vRI4Ltk+mzG4iaA09Istz4FtY5vWV0HROKEbx0zwY
0f9VOJ/m5ku00/V/TFAcGwKamunsCC/DhaiG2zTsQFYQrMd0FmBqzQZ0dHOK
vNA2JXGLLq/UsstBdZ162pTAe+vfyoVDXguXshmvbFEU+Rm/G0xWOFPASER8
ZImztu90Z/RNMQ6U0WMgM9Xvxrww8m3emZNl3EFkUZvpaWekW1CzGx+xC3uY
2/z3NNexxUBv9en25Ov/4wxY6AGJhCLl0v95lRLj21DO5VbyVzbcoUJivXhj
WPTZI9F0w0exNHPzfj4YML21s4cy6VCQjXebIqtv6SWImnacnbrK/yzZ+diU
F9JtX2WZqf/zGvW+/JSldEf+9+YIrW/LTqdjKWxFLJNKdA3U65Rg4KoYWSD8
80xbhAKdQs8otZspjpONV2OlBafIefz9iMXO999FM4zItzxusmruopjNZYOX
ZAkIenhAZDd4TavW4+vbw7g2weVpuW3Vdx7bv7CmQLFYthER+BQUNxzDeEgF
j+KTP4fBnimKvFQ4y3JRUqda/6C8qhA1BpXllYO4XgjeJWqPdXZdDBiWVmFk
bynSHORkbJ9szToseJmWP9IZNUYXhisi7btKafKdWYFUVLEMU0CkXgWPX5vu
oZz+X7hpvSLzUYpzZs5lw/v6aD/n5Ns05mLXXLAlA0p086gjrNMljIQHwexH
4UB9p1FHK3GCCZqMofjDiNhOqhe7oHF1J5NuhCANH8M0NHIuN19WEzxZMAaX
0+RSX+PJ1hNE3hCYYnfpyU2hUam2Xc1amPuuBt1Vi299Ao8AYwfNAnTQmo6o
gdMW0do/oerx1/W25IblACt66zi65jyUxjBY8cC+Im+vC9xPJ+IdG8W+/OuH
fDgFr5A6SbNRCUThAsV0IK37YfwMcfuyiUoM3TvyXQJBgRQXT/ETerKr5YJz
7AKC+ciMPIkzzmIXijfsz/fVWiuZTRuijo17TZSfNpfdNkOGYtHx8kPhLx0p
FY2KHSlWYkF8w1ybzSV2kToOSMyXUQaJR3ZdFgL8g9QXFoQcq1ddFGB47fyX
EOYCQlj8ett3NAjtEZgljQilyWW0FScBv/UmrXa7453Vh15U09DL5oAFetvV
Vv2VB4IBrcCvZHCTXhiYzbyHiqKiNUW2qij/joQm1Ro+uoGeqCsSxKF0Esaq
pHfWJo0wBo+ZtLVXORKBpPYMcEoRSuwNvG0LyNxUn8yEsRFjEqh8gyA933XT
ZbYLt0AyqRPyQHc9LfFYevdKmbwDag+wxk67Eqs345ewlDnf8aBGPgxkgPBU
itTKJRdQ80sdgygX1W/J40yt0lckS0Pjl/9XAf108GziuwS0jNcLy9k+bIfm
TbTQFdbT2DkKscGnvTO9Arv+vN+eA/Js/QIrdlBLH1zV2oacU7JY7LgG2evB
OaNnbcgRUYnLdP9kxi3A+V9DCfE9gYgFUG8s7S5BfeMeLB3pOllbDwdDk2H9
scEHpqeMxIVYH/vcrwyCt7IZxqoofC9pR/ZKC/FWG+RGQ5u/DEUjjHdsfo+6
CrDjwIToRkx88SJwEHyM0bqQs8BVroKWuNERzPhehFQ6h7K/0FUITa2wdKis
7pGWsF5o5lsct9P8aEeis/jsmfZoFwatR0ORdqQ71Y5En4p4UmXDXlYSBcWM
mj0eBhA3mxGdWCpPM8Ib+dwn7CTrvs54IoT5LH2PAyseUQpc1Cr+J91UtxnY
wOnx//XGb4w2Ky7qVq5m6O0qRR3ZG4dQn0w4bt+L+b0midMavQh9BpqOsbk7
xeSt6dLHUv/J9/palgXhGNVUylnCM2EEVE6FFk865oB9f+ROgNGJ+FoBWfMG
GUU4nMxv/ZbWQXrjCHHznmY/UAEwpeF2jw9V9u27Q+fS0QIdjpf/B4E8Ljgz
oMpQd+Jlv06Oq5vjY/blgkqpjeU0qdckgiia5D4w5tOAmwSkLBlzR9tvWmN/
04zaHgyGyFJxnXWzO91Y9SJjUXfTjAWPYYSU0Wc+iSc2YouqffBs/w0FoEWg
QiOJnHrN8L7jqbWVVhLCm09Fc8cHH69UU1OTBBWf7ZuFnxrBk2Qpsz3LsLq+
l52j3HTvx8seUELTKRQC1O7kWxPYWrGOuacXiocnMczwafbscxSMGC41RKOG
UYcXeXBJZ7nrGzO7DeSNaflbzWkDcm6KoZzzFloEJ3bVzblPl8nuD21odDUH
xPQQJFKjqlAZnTrlYizce8EY/RDTBRBQySO8FjcbpssWIVYbpB/URnNXQfNV
ivhW+XiAQ/lsPZRituhOUuPzZezd8Bo8D38qkH5ic6Rro+ldF+ASXEgIPjBD
wNqOxgjpd9nHE4O2nvYQ54h/qiMryrereyRGQcT/L1b89Vwxdpkm9Eb2nJWI
rOR9oJJ99Elptx3Jdqyhn3SyUnhFxPjD9PHMxPSVYRVq3Jlk7vmaAYPBlYZO
ZopRi+yG4Xuqtq+cN6e2pqJDAur0e+H3ds25PtwpvyAdHGBxviGeJtuwIZGA
7VEpb0mRyrpKG+wldNVGuADWpRcPDH6aqTbHgjTYam/GJgkCxEEJpM6LD27V
iOBW0t7wCtX4IsqPMnfhEdQyTzqTHUuXH0E8ne6onwXbV9+SXOdh7foNz1CK
/q/pk3ti/qzyOgMwuCU+8FPAwyXiMx/XZET79xV2BJNH2dp2dRS7cz8/l56l
lX0j+PRwO1QripVTOt4DoHwB4VTFTvhxDRNGLtJ2v4tkASmuhbXt8HB9KAY5
bXaZE2lWBMapr0Fye0P/t9xoDNcRNp97anehBEEowXkn1KWbLr8SvaqaRp0v
hdVXKvjjk87XmnZCWYeFShzpP4WME6QIkInjES7eALCFs0QSSzuU8l4OEffZ
b9uYDdNuo1uIQU/YTlrp1dt3BUpYlgYpb5xtSGMgFspr3fyMNNhTaW4hJIZJ
q185NPISvQjaYZcBRrG4PGYkvJZcloRMrZ2Vd50PordllrwD0NliyR09beuu
IslzytXBcB1CV91ZHy3Z23w7h7ckRUJB5o6GN7qn0BuNBZlm5OYpXIDEOyY/
AdD3ZDB3W0rHeDB/P5g52cmMBLOerUymgTnypOj+H3xrGBcd+JlinndSXfKH
e4khnJsm/5d3+ifjoO6uxAqO3AtKuZ8WwWWTwak9+uvy/DCs0KI6Ok4PeuHG
gFEWWq8remBSXLDlel+2hhxaai1W2npWBMaeguxl/NP8RCLmSamjV1tDory6
ZMdgjvtuCnvuo7so+KPZGfeHhrnMldAdbdov06z+dVL+LoLxR90RLJHAInJ7
F/KHlcNrxZaifc/GGZk74LEkOiEqZUZj7gXpQDoSTQ/usaih/oqGtcX7N3uV
F+tGAx3wuAmYgEsM+O3a6rec8bakSoZeZoXucx/IMB0FGw/6NZMzbmorqYDi
3asIXZc7G+IuRmVB/Nd/Y0IORb6K9atT1OFmm70UagsTD0UqQ4woi5UgyFkC
wb55039mIJn4gQlPA+k1ZHAi7sR80ekj7JQ6IVyY9qls277N9iIsjzQprPX2
c1gkWJbK1iya12YXxlkMnVdwQ7FyMK4I7zbYB/7hr3mHGtyhXwS4u38OsM1d
7ZPKMxQKApri6k6Kj/9020jxmYHU7SnAHTMWRG4OE+DYnrSsZpbq8QdXuj5I
F4dK/H7s/hzDaqfevUBSb9rrG0HiawbbSBX0mqouFdW0SRm/sTnvTXJg+rah
49sRH5nZQqCCIZy/fIqLFtKkbekwFQkTl6lfsj24v+uw9UTG5cTHpYcwmxh/
dWnVVDY1duCPuOFS1Ht4Reua6Rq7pSqr3cfb0MqCCCbQFQQp71zSAKGfv0Jp
b3PCcX/DAqxL5Zf47JVN8dkZ8OlQpPhZwpG/3X5nwg/9QbKHwvk4sqwu84JS
ZeXS6sFTqPWt6coXvKwqhhjxxic/nkKWQe+s6+61aImFc9poA34731stw38f
odscQ4o1DVXqrVaBXtwAveITeOeFXvCICTZL39PLrqVkPp5mezbOIHvvWp+V
gAc3thPYBjqAdp8xkGHiyu9P+Qg6gTs0Ibb2yzuo5GfP0H+eFK9km4PFGT4u
d9+sqsIR54kbWC6hey3kXDuV1B2wRvZNjwn3xIP0Jrm01L4QsfeYbuF9/vcG
0xW7t0g5a5j2z96y5m9Yd2fZxtLc+/ZfD4sTuKVQ5jQy1JPM4BznF0+BZ774
jU/HrjiONQSQVn1MhsG9K147nbuNy/rIIPti6LuoXYf1OfjT/mmDiXf1Goih
fjeZ4m5S21T/4+Bt27HO2E9WeWpLrqMG1kpxxhGqtxMTgL7stbh1Egm/LBZH
U1RanqbLcYnPrd+fCYCbrmvTU49N8W0CdMdgKrf8snBYtdZK9gBo52hlV/yg
UoLkX1nAHKdeSYOHDmFv35mNawUn94jChjWE9C2hF+qmFN9qgl1BqNLexxKj
ASJC7UzNFOo4d1T5GJZVgHKIrpIgseXndR6XNEN1itiKIhTckdD7mbr+X2VN
z//bnZnS3xAUzH42MCqgvW/bDGdQhLs+AH+XoqjDuQrwWV4v8d1Ly8Ek0QPp
x0OKNmNC390o73EQuBpVQl5LGlBcXuZv9rYYGTPDWs75PexRUZdi2AyT+FnM
wAzzr3EDHjtUR7yQ4GYkl11ZzwlFmY0hfEFheaxzE85N0QmSLQOG87V1yoXc
cDoNUgrDsCa2odNZqT1OkdxdiNIUcN/oRM73LJn6fYbxzMZflrjRvVdvPbRs
eElKxiIhgWOS7xFfgPmRwoIvijMUXucaybDq0d1ASdZwzmzZhZZUiSZ8FZ5O
HHzO5WpGA0Fxn0GyvMtPbb5bBgotbHs6a75wZYXZaNMteP0v5in1viOvKjlQ
Iem8wICqvPWw7yMnEpVPe7Jzl3MQkka26b08s5Xcw6qsBet1T0U6BeyFrdxR
yY7minOn1qR+DDZ//sKb4NetPkuiqGv/svgBfXJZO9DpxVOEHa7GaOO5IU3B
CzQi/TGXyxg9fBkoLzNfcWSBi5Qk8I6vUDbFLdks3MzadT50tzU+Sge5xyIj
jw0vXLT+a4BvI5rxyvbohPhsWsFcdV1DJX5TlHMKRyLCybYK376DKoQZRE6b
g9hw3RuPefFApuu9oDI9r+XYiTUoVWm0AvlRU/S2mh7RvbLBRwtmHuxAQJw4
NMoRJeR1LPFRNuKVwiuXk5//2U5QwVptLP5UYtkWAvTVNOZiNvADF8B6yk50
H6Z5A3YBpXVMuJG0VRIHp3p/ObGxO0oU1hzrEetn7u14+50603HX7N/WPl8i
Sv468O/ihvukLx9eTziuPJV46kNou3qujCGIrN8AIQMsYsPr9YD1nSTrK2Lo
ZlXCbeL4qktBzBtb++7ALUf9fWguMe5LOy1mzHgkL5pml/VHC/1tzDuJ3B0u
AmqktLZfGN1m8I0anxv4iK3CMGGglF2h0yE02MpVQwt0zDKNnX0+XXXAwaQq
OtUoXGViRBGynmL1+TXbgajmle/nxHvQtyI7UsLtg4hl4Q2pZyQVucVN4zLI
Qfdba6w3V5Mg5JRcZaiWTSz9W30VUm9sjsVnUuXYsecYySf11JGs3x/iMnZv
AcJjWcR3EAFyZaZyQnlxQ/lrfNOTbj8QhOOdUfcPA/KPtelq0YiPz8bxOpzD
F78z/RxISFkL+4vXS7fSH3/xYE8AmUsFFN2Z/Dn2cZjmg76AIRs9kYo6/s+7
k+aZJJODI8hMM4V7eYlZtiGWete4PkxqVVfP4VNtj1L/lwOJNyrP9/DwaVAk
4hpYbeg8oUmhd0Kg24JFktZ+S3qnPZXprFhuUNo9juEzRGRCo+6fvi1p8HGY
NKJ1/wBfJkIOueKVX1WJ49g6KRRwZwoIL8NDJ+Lm5lvoL51R0DKcEBPuszul
jfJ19n2kp5RId01lknpcyvOw0QD2MPuqKpcOp8TB8/V1ibLsrzP0LNy7dn0J
6CeXjYvXTwO9uqfkPfuKEbtwNLB50YE4m2BKOkfPfY9QU5lwvC0S/p/wP6gd
Kr64fgEggNfptpoHtIPL9N67Dh/7CZJKAl1V7k9PMYzqTuknsPYdm0qUqk3X
gnjvI5A5g6wRvBZOUnkwYD9iTFoILOVgfYS/nZflCWJpdWSg+fJBllDVY/lb
V5zq7BJ2YJep5VE2JUmmRTHL6beQi/KRL8TBtcxKrwcQlMYxIJ4DFN8zquYx
fkbkVZ3VHr/pFhh1yISAgs+vrmTjeyUlox80g0KWGBBDNpz2fdz91UmqbUMx
aUoSO6x3JeXwwRvgYwZUIao4+ryCP8BiFfUoVCRwdwqxHbDTyILBCMhc+Sqe
ve81HoojQJ1I/bT2Qw6h3rs69BdBuV+ymQJbLv1potoDP2RsQorWQzktrHat
yDadH9bDQ+z0qI/N1s8gBGrTt1QO128aWLsqBSMpJCjOUVvUdYsXh0N+LopW
29NvBgl5YnyI/lQzWpE8ugR9U0omGpnXwKGnlYJcPVwlkJ4Cr8gWZ+Dvk5ua
VAPH/5GtZ2iQmpRh0RIvftyJ47wnfewW13XrRjshW28njl6hF939nl8OrFy3
uIIq6JMoU1BtOwQ5xLKhMrqzWHBSZ3/kMsREjYytLDg85jE6KN7wFTmsoIfy
vC42qrN+zgXwupt+ZP7gY3CdGc0vCRW/P/8YTsAGR2PYEgo+85L5AnLnYln+
wJCJARtfVcmarzPd4MdcwV5/9Sa8VGZROMnN1zfzpVsY9z56WLJf4g3BwWY1
WofDCZq+AtzjtYFJR+ed6xlh4BQOz6A2E7OoMYU7iSeOvrthl3Wz3dHFhi2b
tpQBD/d6J2n+Z7GjUCLzGyPmDjyvAp2wukK7JPmtUgHDr69HC73x90qy/RfN
8FmakKnXOp6w3tNuroIeTDAmU/M4b9hvclA+0WpCu95I47nUYZMqU+ZpORIh
3YfvlLMPWvPDP18GRR5ypDAZKZbvV5EVqcOrxYtnB9gDE0mDhwOpB/a/QnCk
5N/JGitShsU5oYlsFzjH1Z/3CxKWeYmNhifrukY0gaVQdF8DXfE0C6h4s2wC
ZkwSwvb8wHqcaZGYLx/tyGXb08ksyOgtcRTOQba2b8obk0TgI86o9fCrMOQ1
a6LMgsXo7nVvmKYOlqV3bvjmmnGhxzjW5fxg029lsUhuIg96cnx+IefrhWCi
bCQe9eSujAluMQDG6t0jPZzSXy5c+tQ0X+OK6wWOtnHqGKlqNrvBP4DeCCVL
bvHiwjqSSJ13v3b4jhGPCmDPFhksc03FeqVO4kvpAet3ELK+u+bBI1zvDJAR
bRiJ7DPfvgSlEEDBWNKgOU0dMmKUh3uoUOTnqU3HHkdl0SOCYnC/eG3ZJhMR
HNaoMxViFUbGabiAZMvSO9X3sR3dT37V8PMWY4IOBQaGla02e9b5zZxlMCNU
4tDG9Ulslh4j/77MPnAjuft5rB+IVenp4tBgNqaMryg/2/C89qGrGjj/JC4x
E6bfrCBGoox6j4lluLYVxx+ZzSxHW6in+tD/1NQKo9rIc8yGuiBoek5TqKQf
vGFfD3/W18C4xKL8csYm1Y/X5h0dBkV0MkO/m1UDiJIKSqGfYGOP8Mfc/+Yc
wYiPvLQZSqa0Ol8cFgTRMjVBTbX8X4m48R7YDIGWuPRNHJ1PbxK3fahugNRg
g85TmP3sQZP+6ul9Y9AYL8KW/hJWR40lAv8LTt89zexgSO0eVTWufOEWOFPM
frbZ/aqkeq4LVHUBG6nKhGVroIJqKlaGbrFEopdJKLVupCNW+iO7eiiLjQbF
mj98LhQL1YLWiuh2wE8AnxF89ShZBHwbywvbz8uEe3UNGZ/qcUh/yVVRPE+W
DpC5x7i9jN+Tp3tPJMGbjxHK8BmhdO9HyFLnhi7q8dfVg0ymnnPToaHSe8MQ
XZWnteMXfmcTUsrumon3g2lan2p/57s9xnk8wV92dX1sxeMk8OnuTITDT7l0
lJ0AFrcm+nBAd2r65I5FIYs+btbL6zXFOf+/zdRMuhexFP6X6CGVwPI0TCxR
W04t3MsIQ6KFpGKD13a2OtoxX1YgJY74Cqbz3cFtOITqhdTA4DBFZMG2wX5p
Ij8R0Z/AIOj+bfstJ6IewMcG4g6n0ANah3IikJCpXnUCARCrdoE/m0b8wYfL
Czwm7EDmeEf0HnmyaGY4ubcteNEoU/znJK+7cl9cSLS36baB9FeNUK80cGSr
2SpnQI/4Iks5EuN7nHmfbMuKxdIeulUIGCEPNZWj4y6ouVLU82UJ1+otx/Y8
4rh2z0cIpFTGzYkCu0W879GbNx0+AcbF7qDuoXqKLDbtoVCkyMR509PkXepb
L46MWxQ/j1LK8kA2b1Hu2T1oksWZPWKrobdlsUCGvbDEuebifysTz2quR5/H
v+RRCBfeyr9VU03QnEiTUSc+P1Za1r7vFrDuWCvRRrjDwZG/BIQwzdZ9sZ+4
0qpRplQZbzhzjU3knguTNta8Q+y6qHcaFrOrYZytzSQ91/M1Ia2H7XrbeYB4
B3xJNRkVHn0g28Ca/hFW5j41Wz8a6u1MOtreYiW7jdiYTiSqtsqoE2Y/4sgH
LadiRoZOBeMfUVWPzW1TRf+MV7ppJWeRj1yH1ZBP5F64MzJvvDxuHOyj+r0d
qWKIS+XWLvNvgf3kEgq/KXgJ9cZqaiUkCvmwIgyXt9D71yEOv9he1fj5ZpNT
HTy1kMA/aM3/Q4jdFZyTv5g/CvQjW+UezlQevereSm3b4VqClAR8S04/R89O
C3kGFwTkQVzwsoEM3e6fPRMxLdnJXgJS2cd5Lf8XWDFWhhympNAVziUSSY1J
gruMF5JlU3dQmFaSJJkBc9U1HaSWNcCrvwKwMA8dnd2BU3rgzk4RokcrqYL+
X8ImgQRO3isy9EGaEke5Bz8Cq4B5PnEyIlLFmplOdDQGkrodxO5hcDU9IP3L
EmcbI/es+YGbVrr168NgO2ky7H4AbO+eNtIlapNG7Fvdxu8wGGmwmItyWt0e
IWBC+KxyFA9/45VGHwdX2NA38gJRu1srbZKTcXHmN/aFGebdOyXmT3OZrKyn
ciJhYVEdWDwK+PQHOzhKVwpve6nYpO2lDAfue6/URJFg3olatSBlC8OSg83b
lvRPRaa2Kg49QpnZYoMZBRqZtEEiQ2+rrqxtNndkDdDQnc3RwB0FLx/+M7L4
bUNzJImP9Y+qgWyFiUAxNqisSuFQ+CQBe9g5w7JEPoc0/Z9DjAxSiyiuqYzd
MnwO/6/NvRduYRWJdL/+MVxjj8rWz5fTDXI3tiMxE3A0VRR+HUxe2UVnoyVO
2iNRCpISfekp6moqNdl3g6RR2yCzRgKtr9NpN0ZPr1euosT+TngkN5a0i5Z7
8SZ+Laaebudu2C67NH8TKhzxG0tcJbOaBpMa8o4y9AscDpQkuv//FaoCEsr8
dIlKNwcbWYQuPU+gcq0DC73ezy3JEy0Kxv9m4PODqwbOvJbrBk33gAriDc9Z
pJ8eVBR0RzCRcsGObHa3fZnf9ai++PRqh6Qc2ot6g/7SzNHTm54zhzCTv//e
uTGwNPH5HALP2207BMos471zjRcDn7cWP3yDVfIKnO54In5isR09P6uaQG2i
IstFvkCR9cOWqnh4SXxJ4BOHpEMy9kjaCzAfeIx/UpTnV8FatXrBV71OjkKL
qeyG9xyIKKG8mLIUpfWD0RDwY0fdZMOJNhd6MUm/ZX16phK6i7dUPUHacXw1
sjq4MKe6BvMKVnL1GFrwS2oXGnJoaVZdT+N2VRTI+UTqUMEptAe863+Pm1qI
Jcm+OTbh9o5tNkduJIaSpGrCyDSP1leSxu8sUWzq3fSfmyQSM9KouXtl1QgT
uhPrms8b0B2RVfoJbiWh21fFUbpCEr8j3lksAS4JJBI4vOyY6tAAkTXzzLTq
3J9AUc9lpI2nSwpnd0t224naa/Wmafx7qB/xmqsorvSzg9aSjItcBu5nGKxD
6JqoUDr3VHn9FPhLLmym7HXQcfFvWqu8Y3iysQ00LizBnhcjIByJEQHZQw0r
/J+7oqN6BRqSb84tkonshHiLokV4Eh8NhTS6CpkZ4IwM7NhEgPxQcwAl6W/t
Clzb63YvZWD2zhgpEfGL0WkoJvMFIABzY0e6QW7JBkuGvjg9Ku/SoVVQXt+f
wtgAlg5BhVjgxDYTAUYdYLXTy9xQFrLDWf4XbyPWq4War4gYwK9MxJ2xxKeU
32F8Mrd+VKzfTeYxudsdlQp+P3vMeo57eu52WnTQCB5vwNj1p27JP2rD7dYr
+7U4w3kff3BMlaivzoBisKdtk7k624XQhArs/Rznpu8QYpb+7g/pqk7zJuZk
3e1km75UpTYGgSjLjCUGjoSLMqnQC23OIx+ZjAA/kVQn8nvWGz2a5Cl+E5Mk
d3GLZ9vFVhJNj6P8te9fuU4JDYI88ior2VMlEuJTgJPy7IELJSFRs7Pr+h+u
TNVDzw99nwGMX8S08y/HMREbH0kwg2aL1MZGYmpFYxF3kzMX0gS2QSNmdzRN
iYqZa7/749+cJDprPlCiLl8Uwroj3TqZVUkcVaowqwj17RuYyA1e5hgj0XWF
Z7gGzh2ikb/f5Vmot46Kg62/1pFHiLRSmeFuRB40qLky4iUsbMD3ANxDRe89
5oXRQR8pN8DLLFl4rUOn/9a2X/vPLjgO3lDPO2Z2lTcFsSaGIlEjOO0BNfRE
X8LVzhiQD206s90kqmNMcWUgkTDVM3+euEq7F+RRqqMmXkjMgEwkXgptmT5y
PycezlqS+oAvDw8PqH2Nsq7PJpp+TwUlN9cardIUY9s/3oEZF5XC6Hgn5ln8
3OalAAcYV+YxMtwi4gUPsxtxV2PThaPbTRKIIko9kfvQITrCb0og98Khv+GW
obc+6yhVyfUbDpRVbB3TU47UW1vslbob3/k8EM5EeNvl8lZYpZNVd99EidsA
gI+qA1sAWCTXGcphD5jPJVYQ5WuGgt6vzNf2qrnWQmbfF2qaOFcfDE2Tg2Ts
CMp8xlbIBuoFp96UIl0uZttmhkDAdpV5mbZ060+mijfCAWCm+fUg5Ae5OWED
LU++MslONUf8APDRO7cjU+ZHjfc9OtDClQhz5g36si/DjXQ0Bg7kuPF71H5f
M7i+tzu61gWsQMfJgPNX3t+wJHMhnHmNTj+/iiTIprPMZelVHvYKVe4SdYn8
pBEj5IQJsgOsEfEXQX8SQEJ6cw98f2f/ytdw+F6l34CeJ60xT6NAI37dZCl6
bd0BwmqqlS8g5/wjPP+khI9K26rHr/7zG1DBphye6qGSfaKKtzM4udpf1WsP
UtzSeyuSaLTrwtxurU7v/PE7HIZX4ZVN5sBh+AfPKC+xUAZkZWjdHVHQVa+I
/N2PtZppM2JZVWwhO/o/FdclarQPKDp8buu3inaFIMYxB2gAU/bx3YQ6dosX
YJG34UUxvrngOk2AkNiY/iifaDbiRPYltaVLg3k+khG6FtAqVbEl0gj7STVj
jECOGWAMlxiWcB+a1l8CcjdHwW4EPPZ9m+ApW4yfBZd16/9ejoelbUG8UCVC
138Xeetk2PB1fz+rU00WTXHP6bjyn8NVS2sF7BDIh2S/xKAeJ44mv2jPqQD8
94Yj30t6J5ZJY8ar2PfNTDnoldQ37fBX4DMtvuaKUjVS7Ou/KkyKqiEpwiBq
9PnztNJrPcCCqIz20nmKNwrR1N/bQ0pfquNlM7Fh1LQwMliZTwqxRJGekGKv
7HxdjQ7WGXcXAjQ59shosj9U5lqQ672AFYVD0nIN5qSPiF/TQMnCnBcrUYGw
dqqOvpljCOW5cHgnLLPBe1eWPTEqxAAkWBAhHvCpjALOCJb8umeKKO37xSD8
D0RQwAPCMj/UpNcwKSNYTObKLzzE8mHu5vVkMIWaOg7i/MkzcBwTmFNeUuUc
ODmAi4BPo0bGa1cKtTl6bhT4T75o3ZlMIaLqKeYmbLz+dWWKbDsQNgOlaKtm
gQ24RaAdGpwZbY8pyYjDpOovaRFaDZ+b/qtI9g97LEv09a+TAJYaqHVb5VVh
0egoA+mFmqZdB2aApHW7/Jab1yo2bgkrCdHZqL7buOzZp5VHuTSj+bT7OZTb
Z/ZFhb15hpkbI4jzTuqVxhMrN0AaROVZNHpei9nKhxDTVg/Q9n0+I+DqVI4/
4egtNAJ+aTSX6wMME7KvK0DIf1vpLb8vRqJtZKgDECBsKJ9+Kj/KP1cUpAIO
MfHcSTXejCUr6IM2Dn/CL88iYl5/+64wgiqzUGBAvFKkVJmSnnieMgqLDcpB
17nxabH3u6lCiiSx5UqXrpRWqL2vq/avuRC5ZXe/8BQaK7pPmr4w/VD5+oVa
wxHTN/LM13sRi4JcPIZhoxnHRIue913NBo8eVU5qJMGWHECfgJjPj085uxPo
VYx5KDwk9XB8AYIt5AejsHGptTiX44v1HTQtzKi62GZ2gSHsIjmIAG7XUIp+
uS3LFdtDNvoG5XqsmctgnSu0V7WSHqQvDEKlY9vboyPPj+pW8m0tjtsiloU4
avtb/q1o8hGakNzTBimtrN92Ou6FXVDcP0zFVoz0J+uhMcLKW4eTumj3bzIw
Yw0zbUVl3HS0n4nH+RfNJzNJI4wmDSQoWXOxd0hxYifsf4FEa3DbNZoGJq5s
1V5wuBhAKSahXo7tRePyYvEkNs/ClPbybqJAhCDTd3Y9kWMX67H/K7rq1Yyu
roAA5LVr6Wh5rE3NOQIEqCbCP2YOgZ45/1TpGVDR69s7qLHtgb+EYHzoUt4M
o5LII4gCXyQv+PZld2opyAs+sOpWsNfj+u4lfH02WgjRuZCGR5seHHBMZky3
yeAPy3EicujrAxGF4DqEGcYPZd+y3U0uVfLqDwdWicAjTvXZxrWaFuE41i00
6gPWp3TVH2FDbYEIlPT4u49ICoc5iv8P/HwbBZKnGTSEgvANqkWNIRacF4/K
xToCk47TcE2tpCTmxiyIB59KtqDVXK11risFVnBy2/OlKGq0pVdW9PH0mh+6
MS2O80aF1eiW6H6L2GGewslHOBgLqIhmN+ScAD4Zh/CF21QaX4sY3pUhiKKS
yyvKgdKwYItCwa9MuweGg+KAzafgnpz1J6Gi37qJlwxEdLwjEfgJ2VelUcui
FJGHiIdiT1uobo7hBtKyIP5XSU0hVYYWvP0Rjty84ZDrIKvGdmipurGdl8q6
ax4OspWaQlYFB9zjPVb4A1yL6d1jUZWKPP+DMej8CY6qzj337WD99eVxkzMV
6xixmB5RXWiN887fxxDI+cgZ7IevxPBLjVN3cheLYaoiaPJ4wOFo+4isWgbh
gBDMv6+CwbKBqWfaP4U4FIE1RRxVAzdBfEJ8kaskhsFvWHlxJftpw49o84Mj
LKhJS/5AGvw5Di9Sqev7QVIKi/Mw6csu2ApHDgEF/8Jbxjo3qDUrU3P1kjEF
ujcDNchFiZH+k0hr6+0YJkKUH+5cbQJBjcnlbM8JowRXg30UmjkKHdzp2Mxo
am1z3ThjaoT2zmaoT7jwSSpbBN+VuMYjZgj9xhiOSOV4igt8rc4XmGuDe31R
AY+Rq8yCm0tZL6KYaCOo3jxClQE3wpiPh9WRh29exb0yK3dlhfmvtIXUWMkI
xBHTgU4Zzr0F7GpVdrG7rBggSukZlbNgHRSEyxYqY+1NYL0boZ8R8BHO1nL4
925r6AlTOJqN568V/18jpk1uRMMxckkAhsyr8g4h/MnxAd5ImD5MLRO9babU
xsiVznoEl/VzDiq4HcLOlJ4/PLgnr/dfBoEVkCmKl1v4nqDaq71d0FZGWAAe
Mf/3/NHLi/nLa8MD6wCon9Agj+CnnhRvSdrMwCjg01815MBSBeku8C067U/U
XnjOVjAd6S0WdQP4VTcNs+SfywGuYyyScf5SD5bB5mROZXbwPlypETEpJPFn
itcOn3uRbi+wrbfJHXTRSV3Et9DzJXL2ge+l8oFq1wJ+cSlygq53SuStbjUC
6Xeplr/s7veMi0ommnkydTHP8/6b8U6Y8089NJozCPPK1lcjOiLY0r4iHckc
5f8YEqOVCgd5CBji7Ge+FpoA6aQJ9zkHW7mDSzf8s4NEbiJYMfDxYTru1Unc
HqzkciMtulyvlrb24CJPOiqA9eztvGyBtxychxKUMwBAgI6wTYmfFy8ra6H3
VKoI0IkxTpKxUUNsunsqm36wzdbRVZcGeaXfIuFLTCBxxHkyZWH0F5DALGH+
kyf33goESvHFBSZ2/lC3Cp9g1xNWxboLfj41JIXG4H56Q0ypuf8I0eW3+32A
fDnV2MHliV+9P7QMmOvPSjSOTJZZT/z+wKOpzpClhohF+Z/k+x78W71393eE
ntymBD4ZTwXig6ahwEbPQ+rii3fWJ7dHt6nEfGRHzGQSWXKHHM0T8gSiUsav
EBsZpz4mjsgQcHsp/3SZdpGPMHpWCNtIKOJwgeLx4dCZxpYd2OpgIDY5JZov
YXF5k/v5KsxDYJ/KuDbgcMKcVnm4XZaGU/LiigQGMPO6JnmU552UzBFan15i
Efc0leNDjH2KvHYbQ8/2NRvQU5vc1Yve6vn9hYIe6QNnhCdeYJ+O7Rbw2kcv
szFDwudwHlINqlpcG0XWy7tUJuPpWAeGSL3nEyYMySHNBmK1GiJMZdWAy0h4
QEacZeq07MrpgsS6vhs8BDz0+BCWekqhqtwnOGTHrrlRD4ZGc8+JmP5zxtmQ
uwNOPWQtZv6EfMXh0m+PqERaCU3Q+ekS+RwMpEN9zqjNro4cCsVhrv+ZE6gj
nl66JoxvZA4s1zGHx8jUjVCqtIZlmnkUAGe9fGMAnbLVt66jkIfI9nsr2aYr
N7BiFuyla4wH9jcYzmbDdCK7f/LjOS8VQ7DFG2sBeWdYKHcZVP4Jkqn4K143
YI6ftPW55RRORCfTDTQkX3Qy88MP0kdBUsQZ1Y6zxgrYDRFSuT0MHJ47Ia+G
wIs5qBUrcslRtEcSyLUoOgR6aOWHHfDP2F9cVuEkjp798SJFwH+vBBg3Heby
Co1Gwehd/M5mn8JdvSmN/mC3HAU/KPTPIFVuAtmdsuzDdpx+VFYnBpwOLItn
8m8uDaEdG45keDn8QEu92cSO4JaLtfCDTPTnos74scWbZOXjh09d1UG4h1Qy
uQqbrcWjwDVzb6z9rdVojvR+UFLA4bEQyI5K5C2MkrnzGEqTzBJ4jm5GjnSk
UgC1rzJi2rYymO6PM2LbHC3GqnFr2vhHdQUIMaa4MCVTVfPWyjOqrSZ3k6sL
TQOdfLwAzAqSSutm4+tMz7fSv/WzdQDy59P5t/s+LFUvvbcJ4Nh2n8ZZ8PL6
51YzU1qul6CHgjkRBFyBsipjyjt6/l5QceyccX4gl/WY1/qG7jomw0mHoOKa
zRgBdy1gw3aeAvcur29axP642upCHqtecXp7HsfDiuDhPn6tQTUNP8ucIBrf
LlX/uYraKYfOjx8132E/i6WPq4cSnFcPBHlgXtLCBBiWE/Z53eHo8LPTLLAp
m0JxYukIjPyw4JoNupYPauaUG6VHXrPQo9sx6TllreuksTN0IZalVp6f5+Ag
W8/urqax7dkxSlJ1dxSLUAVPKhnwJG06kD2N3ApRYSYUAqlLZKItwlfvtaG2
/bSKVXkADyjfzAkRRNQZta32oozvOoGNUOTqdQSu7qOmb5lAOQea/NnWgDuf
3tzL8r5YCVdrThgMm+xopFaPDJIhDri+7uAdjFdgblqwykNuCK7t7TX6w0wT
7DiiC+/A7OgU5+DFXKC2PAgnD2yVPkCY8E16NOM1SrGgDgTblynilqTi211G
gNXM/DhKbBPYFCF8BSlm+c64Z+jIw1IjcItMHweMEtOlIMzjl5+1F1KPtbqD
YPl+Wtb6zlwRwb6OgkIvY7uVBVqiDJEAOMVEKIJ/vwmgllMhrxM9gqaKAEyN
ORDfCTxla/1VXIAwHZR9SDUPoOj0lUAdGfEuPyJE7l07QjntGaOyvSpPOGhI
ZMD/wmYycuzef0/nIIKLBCVUCAVg438bTYut1IItDdY78FIFg7DLno00R8iu
y1rIUohD/IfmzpeuyMNv6LH0LxvTUJdMrcL0g4B4flOBDcKWzA9t+vtgLa2c
7rSPXFFW5gj1QssFFzwIvN2QA/dUgvtFQQHzTL3RE8YoQylrbfypdug/CA9S
6XMDvNfforpEGpF5Ei0jjyz9OixVlTq2QRqN/Mqr9vgEcX1ueQPENkL3yQDV
Hcdi1/aeJXP+R7iCq2bhvt0NCYTQapJYIcS25M7r45DkpfdQl2yh0jZ0qFLD
vmA2VB7y6C2Dti8eejoIZoT2OuIv2zHZVX3qh9JrcHoXTwiuybABisdYGwZF
99vGESeSc098uVETEzOYzXvcfbX0mxCkeCAfuu5AdX9KqPj3UI91Mbp2BBDX
P0m8RgUPZZ4PUcdTQECihsySnL3J/3gqrb84og1V73ob/9rDaBwvO2BJfng5
1x7Lj/kxuyHLj3qyInkcGBZnTw7Ht0UG4lfMq1JED3jjnXDRAbM6H5OEWdv2
GCt68vjlVg0tXa+uRCb0KKOCtckY6wN4Ff3YGnKD36LxiknOtTT8loqPFhmt
JrO44JqvvVFMBFotACcCWKLYf8lylV2Smy0nRp3SHtmLV6mtYd0oQPIrh9kK
RB04KXZm6y7Q3fU/43sRuHDT1QinQm1YQ18ht3w2Z5w8OST1CyBZjL3RJlya
NOEeEGLDtnzSHMgRnx9VREjCtUgOlKQ3wpMdjsPdF6WaW/Lp4ACJokpxUM6N
YnmFSzwa2FORlwZnBANXeYi704IzjZ06iIdKoOXOuXSpKTNEeYHrt6hEr2a2
T9K8/PbkQ8JPe9D8HlW7X2x3YO25t7p1df1NNCHwBr0ZCwVkLXzZYC4lkFkp
azLbvtGAnBayQtRjtrSoyVDwzykK4V/R5KIubbtWm3Y145RFG7ynzpuX+4me
SykRlSbwtbKt8SJvctXib/sr5BtKMFRtvn/K5AwM3Cfka2HrxWDDbv/nCVJv
BYXyb41ckdUslbmFaMBXFtQ3Sz4vzr79ZyI+VuxSWjcAGu1I8OwHUUzYn/gn
h+DhhxdBbuF4WNn9Of/1SaQ/0dnLsrWWdaLpT6u2uf7j40UWWarpL0VLtz03
cLuO3kGtX63ZdcjvVjsGOEf8FfTArxG4wHwAADlIU/ZDjwFBmjIgDjnkf6Ok
NSNVnoE8HHHVDuYynTJdtFHjzVxqPcIqNzBy8GNXUNTTW4E6sC6U4s8qzetN
OAhUcCI6ryrIkxj+MLXDEsFuXUl6MjMvWGGbXQ3062j/ezN8aNGHBLT6YlD9
5t9qijpUKNlRUS3/rLDWxy8n+cTk6p86ZsmxX7OE6ZC1w7LGba8qYROdETPk
48ely/AWbF3jk209hiz+tVc6bXw9jFTiuFYgpzaJAG2PrU2CjeJTZ3oumQ6J
hWJf3PCyaxOLRnLJaNDxu55/jH7xIhCCFq7cRp/mUS/btdZHnh7GwqnR74uz
3m4Ys2HZrrx93wf6pnfF3dyPKHl6NDmcGU4havhmWGba++pEUBmLyY0RxIBE
YYF6JXg9o9SdeIfcrqih7E5ElKP69YYz4Z6qd1vi5dxAx3+cGqioCsBBvZXc
LoMqtyM6954FY1UpvNq44phw5wGPUV1yhofUwUnBjO3rSES501rrXPy0psS7
j/M/Etv7TfaEUa0CNZF/kLapNNuQ7wFnAHrlTYwtgT+86OaOIbASZWedAV5F
stHpTmC4FXza/xOHu+dEIAHF9shjY//+cRXTxXiex/fxR6e4k9ItSvDqfRa8
Uv1euuLzri8uJo4GOIOQAJHLLUTtrzGGE+lWK+E7rU2L7nW4+jN88sMIffpM
qOa5oR1uEiLwV8Syv92wgtViC1trmhmltNBKwb8RGLngah1NrOOuu+GfjYqP
isnmks/uhzF9//hk01wFSVxkCsxpNr6b5VNBXDO7wUXRoill516PPo5W7T+J
wzX/UOnU7QB+I2WLOTvkhteRTi8SnPDf5mBuR2Vk+RAPU9Q8x7uKxFOt/uPX
3/Hv5PzFb9gmM3uGf9Kdi6W2RL7iPSeb98LGWzq+BObGoZ17HHvYt5kx7+vT
mCt639R7TYhnStlRr/H5svtGep5Ds1ZqFBbPkG2Vf4GPQpP1BDbmtSZVwRFl
qhPLqcDtou7ua7Hv0UDVqIDqiQfHnTjp/j2phr7HOAb8/fIXL5fy8xK33FnT
t48tTyA//679d9SoDDk6gYdzvx4uKsEbjAucZYzW5EQhNGxAIx91zu1sxnZU
9ZtduxLmIFjN77c4lax5dhZZt0t1jDyjCupwnArZbkrr8qoZeZYy2jkEYcaF
M9DSKQmu1/sMPZMy3SEqdTn8aueG8xwO0FfnGBpGtT9LlQ/tIZtySZDNZ4+L
PMbdfVG/Pt4wUNayJW7Rypa76CIEEJJ2k9++pJAEkfx1QPixHb9CsvKXtzKx
z2zzttlpO1+F87o9tjCc+3AGV+RpbX210edOISZqlcOvvwD9chQNSILtOyHR
UAsPK5hpZ07n1HGRX/KAHKNwLHehC/0Mb/2mRUrTOwbwyOS3Y16xJ9c1RDJD
R2Jn6rm62AFcsJCQmrGVLCCqQQWM30yje9oHex4iniVCwKJVqA6XDNgkUDva
imGrT7Gc7U/bUvKyXK6G1lDhn2Rg6A++SvysK0H2RFX6dzh/EDL6XfKJdEY/
BIgpWINcp1/Zgnr3zjN4yGLV+7xT0IeUg9pMJ6SfwLpceLFeip3hxSeZy8ri
Z+hOlrmWvtajRmyKGgA0eAIfeWroquYuCoYjvkjxTUE2hQQe7JC5xA7k+LOf
U7TDZybvizH4xwESCwLPULNpDOgqmTcoD5eqdGR4KV7aD12w3J1yvnZWnf53
cfbmW8qDw8e/Ga8mVkUkWXjzR7b146AUSm8BkDvB8IsnOwzYsqXWcyzvTq9+
4xhU0ciORh4h4zEDkLavl3Hi0xn00AuCSoN1mdhWGhhDMJGbejdlxoZUmhNI
8u7J6YskzUAylfwKZ9tDi3gy//mbDfpxhyjtR35R8T/d5Xkvvwlk9JcOaMZa
i0iAhA9iJq4XbcaZxeRUqNRuOA0kcgxifCih9oM2MDHSVgypWWxM5vATHgA8
ySJ6R/z7k+BY/mR6BIKMXw4KExFB4ArrU4tIcobbzO31Tgg3SLI5FaI4ATdi
vKChO7Qp3c+3JeNPgbvjDhmh8M3zKp0y4QT4krs66l7ydraVSp8ia3uZnM5H
x1+C5zVm+rTyZpP199cvuieNwd47l0QDfBmRMfdj+qKEJ52ST7fXyRlPDvOA
fJB0NvS8iEnDYRswxMPhoEuUaFSq/uDclaldvensIrGARKxSIblSkRgP8Pad
FYWGlPToGEMNfotpqpvSW4vfUkwxZyAmgDVD6xgNJFJtkoBc/4n6uj9kNkVJ
Z1Cvh3Eea0g5bpz2O4qlydIuFGacO5Ms+WNENy6Jwa+NZaPDTJqXkVBVaBrW
4t9IjgYjAUuXwW51TbrzAONhJJyocqwWl+dPgxukJ7aWUXGvHoLeK+laB4GF
vqQ3W+UKoYEzWUeoXNTIB8eJvC03qhaQgMsORzDsVMvH9i5Jz0eAXklw4hpI
2GKkMFF91fwIwCrq/e3GEFr+54IdlFFTluwVI1P1Q5zC2hKQnKZmpDmRZ08i
qw79kH37bD3L6ObMdiPYbH3HPlfEP4R6C5ZHUDcT6uw1IbClvhNLv2VPOtsr
5xLKBLP7w9ikv6ezcauVe/FTfLnEcRKKhDkVueCnVur/9s53EJs61tBxXljq
7WE9E6fHtdhk87zfnnQ7q5CGOlc3oDob/efN1JC/1s12LMjcNondUHmUyZea
5j/bdlF9BP/nyRyEanXrOhisCaerg3otS4F366ZwtiwKK88XJ/il68FssB08
GfniTsNol4WPdH+0/eWGzEaw/PeYqjZ1Al6yr0N9sTGZhVFXGS7qcI268/TP
4kPojhhOTCbHbwiZo0HaNn4qQG2yai532Z9+tZrxb+g2eoT1jJHltuUyEYp8
vRf6iG0ywymd9tgzTktVTBJZ0yZw1DQwIfdUzlgP1JUHr7j9uHZ0506XWqxz
KDLZotw9NRZkxbPBcfl2SE8k+uqbWrCKBTpSQ5H6vxmPopTp+ZHjn5BlFFhe
Sns1SPuleMAbYKkxcxTO7hh5SJMGm77Xg1kVwIe9oyV8ZleRb4Cc0c6PGF91
1JMt9iG48JPMcpJ8CE0IyjecbVPzIAAGd3xTBKNzduEMYjg3+go4xDRmNEpA
RrNlB24MERbClLeAkPe6UN2BSLtO2kik/t2XzlO1eb5nNm5yQdOCqCR9Q9NE
0uftc+nS6AWfcvk6GyW4Du2MABZg7jq2Dv/1cEshERT0F70iZtYol2t72Gda
ZXPBSZo36irVxfarXF904+rt36gQXOi5EraYyaVBvhV7Xg9yYX2G2rJKYB/d
R+BsUM0K+0bUaWXOfGtKxoMkmwiaVtB+QxAxtKmJsqMgo5VxieLaBzDIBoKT
fOLWnivZ/Fkub0H7IJF4zhmjI6Bq5hWEypXT3t86lsl1JZqp0gCXbMvysK2x
HcfnjOCwiqLZDm/4H9x2awMk+oX1cLUVyJq9wQctKYFG2n41z4NIbACcHi6c
fbyjO0xh/C79cWjX4/Blf2DUCLMNhLbPLavgNAnjcDUNqBNnDgWK2X/y5Ag5
Fb8nBsvCokEb0OuliMY3I8/bzg1jyEZQQGdiECGYAdpfRpMPnwZSzbB8Cgol
+tDv/tKb1tRj4WrFYH3GSdLf3lo+s5z7j8esIZmq0K6hcTQWDMgoHpgtSwpr
c2ngKxDFdRTu3z+M8d1Vwt9TF3F4rj5dvMQrHW5Q6NRNduaaUHwvxIs41Rqn
SzrV1+rXtsWU7d5qdxNLvQmJYmlUfKyyayD9KpiJvWz7MsifJKrFPEm6kg5r
upUJwnVOAoxIlGoQpP1GtF9srOR/iqZ70FQBndPosx9pYeYe4a2Da11MNTdk
v/kwbQuNideCeMd6QXhfPoMOU7jLAuT+MeL9oXJtjfcUbNLWUt7/E/WjqlKk
q3tyNEkChGa7Co3Ba2HTWQy3jeDeG1HEvU/Ev5rlKJggrV5GPFUor3hf9uDt
zgS+XWPGw/KpelBuQigRfvgtn065XJenwhd19vWoEp0g1AhkASIs7X6pseJW
p2LqMX5SKfF8hu/DxvYQLDcdzYBPGewCjhh331op3wYsSLC6taPN9QU4fQEg
GvBSnazfVk5HnUYGA01NuhUOjBhplEv3qowKaD6dJVRBLqN2vPNNx3w71oc/
jDDbXPgYVtrGo1Omy2G6vaE/P/3A6ADHRNRBz6YUN1kUXOSWIPJ9tHZd1FNk
s501KvskdQ3I4TvltrJErrF6ggX+vy4kkWxxNajV+qZmb8ZFd9FMMum2idTI
VEXesoGz++OyYT1ArEugoc9/1+dJdj9eMZUdDpsnuFTDeiL5QwTWBQKiT/Q0
LwSFYG9SDx+a56HtwN6t/+BfHgV+oRFJeHc6qmHuSQmA84Qj6RGj5jvuGb+3
qjOOdqUQonABUj6Ovv/JZ64GQgOGG/6cMEeRoeg5V9hsN2p2ggktnXhsaUkf
wFbYz+5f22V5mgsGIyLg2HOrrfMu7YgGS1dWD2P814bEAnzDpNsJthFzFzzq
XTgL6Igq2tfUFX5LUMUnBJg6/4YMBXjvL3u3+WVu0rHBLRfrSfdkhrVuTURQ
xA3syM3XxzI/ceVYbxtx5JMEZmaIjtZAtomKNwe7vFZplgZiss1f8qEXi/aX
jGyQcUVu8EPdEwx4hYzicRjehvbacJp9J2ElG9ow/rtW5BbfdfPz/PIUmIIO
oKH+bOwlMC8v0FJtRQr/DlVbb+KfkXYvbq5H3C63zq4X3W6wWl7f5qhIqowv
ds3XBGsrDBCyX9d7yhhbNCfg0rt3SLUmXI3LgenZAd0lhVH1jHMsxcFmL/0U
jmj8/whUMAf0cOmmA0DDHlqyU9bxMiRU2ZTMu0sWKUfdrP2SMXJt2QhcwrqD
JhBbcf6OJc1GEK5gUTTeZ9S53EFpJpvRe7OS0rq+LfcaT4MYzkmH6bfgFXpw
h+oDbAOu8VlbBF/aAbavvkQH+WzUa6MemO4MlK4+StvvGlFLGU6qXw+sRKI8
Zv0/Q+zOmA3nhZwcy7ZUqjPAmPXYaYN0jUWiiinJeXaWMawWXVauyXWfA2pi
mGJv96WgPwlO7vFqtH9b+YFTUpvnfLmKT6NVGGqyQR/eJWNDnm5UU/DRovsm
usjw/cNm5xqHyJzxwUVMfDogcZq7rVqPZpmDN2ULDvLF1kuakjAbtoRlPoE1
hApaHZRcmIESQbt8hdYYXoUpKzIEg3RsgGxwQNvGKO/WkQSXtwYLLQPNKpRn
jkzhFz6shUALWtcJCwEpefq3iv5BkLNjhj4btHLGAjE4W+M1UwpZB7eDkwq6
o3V2rlR06DKFf8iwN5sSURgyolHQok88opJejclj4u3r/XXVaSNMnnXNmx9c
8l5LFYU69Voz7oLnUcW+XsM3PiEKvsJw+2fpgRp1p6csIvOQAkHT3DwccnMI
ovhnJu2otr3r8+vzGj4vzgPu0NXWAaPOOn3p6CEq3y15Rro8fz8YzZ0tr2Qr
ARJtM5I9c7sfaLveGGqHwArOQt8nQVV+JdNikRwV5/s05z/GdXiK2XwCXA+3
aZcbeoXK1FkBeCcULu0PNJNgOw1+rnZFiSWWJkYha1iW7sm9pr1bPC8ncDgw
Hka8pd1c92h/VO6k7wyjLx7DuKyehnZXqGx4AR08NngYMQE0BcqVYVR6l0r0
RYIYXrPZWBQrfolsYFYRNPUQckmG979rIeKStdk+LtqSYz/lMrvTrYAjYUwb
RQp9TAHsMj3r80+LVMk33CNGoc2cXH9NJTi86dMR3j8cSVEY8DKZQVaXAgTX
0aju+bZbGWHORbANmW85zKWhc9/zOnBQg5g8k+i57FN3DCFHfGVjJfTym1b6
RLt5ig2qu+2yzzV66FLu3ox+H/e4BOivdUKVu3jLwmhGBocTAlES76lm7ohc
QL/pBThycq6yQzaHzz2cgKtFzS2sXdI/lT+9y5Dfh1igYA87JCOtBziO/B7n
vIv1xKmTyS6DOoIgfHmTDrsY4yxYugEzzK24OMmr5wKjDqkhVrChv7H8sksF
KdtfILeWlptg7+HmDD2bbEw0wq56DfeMwcg+B7hzEP7NVpHcGstmsK5EcB43
ZNEf7aN/T/P05wATf+4Nk+Ph7a0sOx0BO9XRsTZZ4mG5Uurb7hyAYHaGjXkI
EDduAmWDgpX4lX/6OrIm+ylPYmhpCtxtJTNuJLiaj2JIQgo4osaH/ecRr2bO
TENn/eE+otUse+/D1MwyC5UItVsgBV0KmQr4A562CAI8VcJj9GWtkExHRmK4
uqoYCi/qeUssKDoti926H5Fzq5CKPpO0sL2PenLdUlkOlQ4g9YtcB8Dp00jd
5QHW/5milU08r7vB+V+jhM21krW5YpaykVkn5EzZaGdmKqrztfVhHzRdts11
htCuRdFT3O8gJyRIZSmcA8cyooTIg2mt4fPy0JFEhUjg7pQOfLWUODz250ZR
ZqGVXfItCal2aAJWxCOSKb57DNyG+T6LSGsOmmKIOTh8s7sPqpE7F1ARhxHJ
WYEZOgPDEM1+qj9GcKXGszURUIfs5vQQqDdWidQ9sZevqjmB5sr4Xv6GmWwc
UWHRPZWgnRv9qWT7eFcQ9Q8fzK/vXmiwzB4BvZUquiDeUF/fVNFo9YmCGBY1
2iT9YKCVbjbDRuYydgRBC8xp9RlckRPdVc6mr9XLsqnJheB2ZXDYpd4HbwK/
q4hWc+2i0zeyvhs7BaJdyteGUlCQGAQiOkef46VyWpWkM7CJOkj5l5BwB51s
Wqxo1o3UQu5VKA/9qt6GbbIWUwaqeddEJm6J5kDnnsuFqPm2mQJsDQ3WAI1i
6T98+H9TX7M8/6mj0CJ6a/KyTtjket6riIjsm6DP855Jng184NEW22IHCyXI
z2gmDus9WptWWzRmQYzGGFuC+2CQHXpDxOGQnoOhTRo/fnbM2ENRTF7ZiT2n
EfxQVZWcWp1+5306NHk5BFU8mJh44dfl6ZNj3ePEKF4aKd0E0n5mtaeKWhJT
uz/7pnhnAwLRSS4S21GCxHH9krHSZYq02y4P3A3M97tuafXls1dUy0r/Pqwa
j8+je6AbgXfGmZt8J55/HtfOQPu6RbtATe1z80zDU5ubTZpW5KkQtb+mtQ9n
n/3w/gg1Knhd85p41Iw2wlM3U0cPKBCxAVZQGj5R1kdx3ehpPEUQSpewPwpe
ipqF8xv0h0er8dfkGMwSw3ux+0MpAFCruaNg/y1YICuGBIgKK7U5ebGcwhbW
8RNT+m7amwcKuyz/donp2NGuD+yTetcRStFetbOUA3wygq3T1iYnbGwNeyK4
4nF6n0YAtZnu/e/IXBg/Tqv+D6+TxU75Ma2Ih3Vv8Sp6YY3Royk8UdEq39Nm
i744Y84XWVAmvyC+kSjRlBo4AY/k0R5GZQSCoHQOrdPDfj2PBw0h62W3slmy
G2lxVdMR4aYVDz9HxqRKeLOZAMqDlIz5wMsTzrUWx5LOQc/4nKU4TRNs4uDA
teLRLuaBNPSF5Do6dPZGi4vqPCh9Fj+CiGiymgLy2Jl+B9WVwbtlzdHWKNPU
TJaUkuvJ2d9GNbrSqb7BReP4Tm24uGrwida7oW+GN3xw2QDOtCiytlZRX94K
pU4pLd4czarUFy9on495+MEgsRctAuNi64n0sWOjT1MppyH3NobEYXGCtYbM
aUPe5ggn8odtnO/DZ/RnsSYhUTSkRv5SKGsvrEbsHHvzPKeppqaEK1JtaqYt
+tTlqiPssmgEIMYS6NbVvWdF9qDQeIXK+ukvc10MbWW+oy4GUFWHzyu1gxWr
vFM/2O5vhAHMyf6mVnyCQaI0Kk9POCc5lfrlKZV5/7Glx/r6gE0UQuPeyGZA
jpmJEubLy0l1SWEDxlHejWOOIhjjkwlCcF6oHFAxciKRL/Mg2YqM+Y3omFtu
+ySczt0n5G5/MJCn6MXdG9X1XwfbYlFVqzyYGm9JtolJqPYKQhehnR+9izIu
rRqUGMa8CcbwSH7dl7mro4ZVbSRdJdySC8J/OQWk4OZGq42su8I4mL1hqS5f
1qqttDyVdd0cY6n5lCOwWHCZ/ewK4uigjQuAK3aQhCkIxNdaqVxLKWXs0v6T
DFmd6NjkFZ1L8MfX9AaSsuEaJt+Rqm/Cu1c0j3udIibLF471E614QgdFI+EY
Ia84fyZn9fA0rWDUqUglU4K1nY+O0kzzQeOU2D0PdQa6MN3pwg6CYs/63YE2
QJMLfj3UOaVE48FexBE19E0oPKEcjZXDV7vgBhEwHl9M1szXrbnIFpASAcK3
I6t52VXp6/lJTN7+UCSoGr4TKzd97N3yT1rB2S1bSKmTb75GRdY77yr16ZQh
aeN+1VGP9VTiEY9ih2QZNnmtSFS+mJ9QK9/6y21VH/6Orvmi8fi0EKXK2dma
CusBysFmI4F7+BJp9pi/pHuJc09JiLEBHTS64OQUhYoNI6lvRfCyA26SAl1E
BPX7eaVj8qHX4MjtPeM4pse/AEk1dWZ+8x0c1PLnR9XoGFqFTdvJ+lv1gDZE
K7FCeeDQu9KKHujqXHFYf1pCuWYrl+XVUeiYZnp1Itkcsa6UGEJcgsztCIWt
9mjdDi91acmRRkm0fU6xcDxB1UZ7RyonRu5dpU4qPKREXcORtJRn0lnBH8SI
qRJVt3VnzhP3ppsaWGjtWlZzOvIOOk4R/BUYVfSP5rixBv0hbZNf7bCwOmu6
69n00sAbnOCnWhvda+MFOUNVwxqDZ4MEC0RgY+07udC7FXuSnb/9eoMFYIS+
nwjufFInxOKqk20bS+AHvhLVQ6Jsh7VzAIagmmxZ6n4VrYiXMkJ9UPPXkOPq
tzR4a94ytzuAX5QnBEM4Rd4Ei7wFtzHno2YDYKr1A3vrL3lLyuCyaiBR+b9Q
xlhDvRb1GHbCGjBmhXSWtQ/U8CEnr8pBW6XrU5QJPka+bM9ug4WYurS6EfUG
mhPfzepynYCjhRyJ4BCggrKkH4Ksyfln8Lk2A4gefKJDu+BXhUkvhPVmiLtR
NRvAEAYPe80luPibmWNYbaNYhx+PzGtcvEruDNVe+sGGAQR0xwP5YY0aYeIq
BW8nKqDBg6pk5nhf+C2S8RML/QcE4shlvpQWwHpl2rnP6yvw8lNjA4MNEDPl
AmuiTU7JlVpIsxSm6MYrbW/RFLIlcx+MafIJs4yP9UbIe3UBf4goOcg8GMIm
+/APdN/KeL798zA5D51gqjUF8vrIcyYUn5RK59DorYiSZzZULpaJ8ZdsfNHf
gkCEua+29SlJUA1iDzIUa43nlILpjV62Wq2UAlK0+HyKDBnUgSXy2Hj59wIT
EGurpoS3Iv6V5FVKfeQgyGJjJRS7OBs29YSfqBgtcNFmftEUXojfCSQTrAla
AtTGdYjZmw/eAQ/L7HmKQtZT9k5U5L/9SSVznaVsPDnhciu8FxNZFhjdp6WR
T6xO9pFaZ0a0NCpMWKL9k09tJw5P7y6ZZbT26/Gy5wSHziO6pgjwA/lsiUA6
0ZHdEgWd7VM+y7uVag8aCdQite4RHRxSDCLBu9qFRxmUaC6etGZ1A8Pt9oSA
CTUJqAkK+esUxlCWi5MxtocD0O2ojbCpOr2EV9pDc2KooMe8YN+LyB1Slcer
AJpHwveMpeGE84EuJ2t0hk3sdLPkvOX1fAt3FeJDp0/QInxp7jD3J8vtQqg6
wJCBa8WwU+8aWq6BNbKS+lZwCg6Cd4PiRoxipxd34q3kVyA8xA3kGk4j+2O2
UJSJO0qmN+NvrHnK20zTZb54xZoNUyotXYORzOypzj7cxh70P31m0OyxfQ4K
FOlIEvUDBj/BoW43XhK+mcXe9VgUpq65yCRG+P4XuDfj1HY1up2czAIlMGu2
CQ5H2ky1x31pzvMzyUfpH9AaFrkyfgpbTCyvZ3TupMpH05pO7T/1sSE4CQxe
E/xQj0fNmqrVDFPF9twc6gumVLK8GSbwkr4DlfypDxNYz/42tcLNgdl1s9Ub
zbdoUjJ2M/H/SN2XGXBwyYk4TuiT3NDolCH8anaejuEIrfdgY5WFxRDr/vqY
/kc5VNIpS6Dr+OrHq4Vms3tiMxswXKPyjE0qbtZ55xmv2gJBeTWuMHiQpZjg
X9Lcy2rAZARjFEIEEHiorm/HxGkNM2lOVc2mXl6PUE++8smeqpx160OSaBae
noyCkMzvQNYJdr5kQBtSN8ykbx1CsDTtDzUBJEQV3QDUYs9P847+7mfsbX+x
djtSTqqCvFUoHqp4l2K0IaTw73Jdl6Bn/MY+LXhj3n+ZEaoGbbD75DnBhsrX
kH7l/HDIo892Ej0+XFe4+3eRSWNWAcPdIXCfJUx2laWbhPCGx8bNJAkv+wVZ
3zpHQmjITyuw2VRQ2zQ+rFdjqjtrcId9A30M5fIzPY6r5r+OcZplAdRiSadL
oERv6YUIJeafS+MSHDNK/D5VZhvz5cZG/7dFZQteyod64o+R1H/1LNxYvLYq
MncTshNubeLqmsm0qIBqqyN+RVpjmAiMKNBofK9x70kQ3nUWyRaXxqPyLNwT
4tpPHlCR9O+IXZW2GziF0f9Ow+ogFTGjxYDwbnViueDJ6O8XxurMH1hwXP3Y
H+L7ipoenGvXmMBMUiM7KXztKX2Xvqle6Do02H2WNBHN9hM35J0O7czqLqgb
laM0nVdh9SnO7JxN+VbchczxOQNMxXE7hUJ56Z7I2C39IAp2V53eFkgMfqgK
QG0ay6S2GyCSOC0oRIOqyBWUtAoPAoJFSYgONpRZl7urNmUffUp3KFTs/VPl
0kaBif7P8snr/qklXd6GSiqG+/anB9/eFvE6gmBpoGXuY/c8VY/3bi/yTLyT
RxN9D/mdyN/5bY+6JU+VChLEfSJ7Te5GbO7QOtgrDaZhChH7SlKNFJcJCJOW
0dyMSEIxUafcmc2ruhMxuUUrPj9gTJvB8svPHse9hGiEfIA6HeJIl1u/GfpL
LxSSkPhPJmyks+P9X+vmDBF6fQVpjsWctSj0nHCqnLrpfJCobhqbH+Hwl8BU
XL4nCQXpRgp/B3/PVUwPfIY37uqn5iAr2bFmsA4ZgHaUYUHcZ07o4v4RwjJX
MEo/PPRq1F9OjgFw2sp0TjQpxh+40KMTL0LqnidE3REaosAy5fRrhymYFlR7
WnXSqeyzmRyRdBF+CFyqaM8UpqHCa1HLYck0thMVSIkybRYjA2yMa9sKO/fT
8rFpYhAxL74DE0ZwpANtdaT7D2ndjykq344UX/qS6rHwM1+xfXIoVdlSemRY
XvqXs83nIYOvIDGcNZAoeNo7+gQHWdzSYKIpAFk58Ts/GWJVbAcnc/Wv1gtL
B2UfE3dqYLAqrbQRhC+IEnRJFFReV3/GvgouowPtKCwahGpyZgPYFqpBRPH1
iGqhEs4IDMd2r7MpYWxUBbxrXecB7vmRRQHibP2Ye1q2XBKu9TeThCtOPwsa
05ZhGje7ULnZrfZmDAULVU3A8mGvVT5FOwjpEL/HWzWZ9TCF8eGEDOxac+c+
AwrkwSkp5AiCrxGRCRahJS9DMuHv57CC6IwlXEqoBhSMNguCrl+ezC9ozZzC
+R8fyPJntF5gRvy+QUccetHloKoPSresbpapKLGR9lowQLC5cE2T8JQhkedw
ZqjH3fKvPUs5uhGlKSiewKKCSr7kFFYmVn6dvyfbcTu5z6uohEdzTooSmpmN
UPm5SeAyQ7u2oR6akntlaZJDWjkn7Ke/zBHMSuYc1PCCnUdgimNGsllaN1T0
bSs1fDIQ88+XJEvmfWJd9FgDUkgYIaNDf7AKM5hgR566zza5QtzIcODOmfSc
OqkX5ORrzv65rSIru6Uq5G+je48a6wDtKIUO2fy5jRdN7qV6Qyb9Cbh1s743
NY7dOsgRXnC7PNtFMV9z+vSAZLLZzD9NWADmUCKyFgIUGZ7voS2Ptny0lJ8I
bsuxPtIlG/aA3i0kkTuMyInwD780Yg5glYjoHFXqO8GNP0raqW/6R+y4NQrE
QcX0lzdat+LpIGh1WlLtR75z/x1uP0LgfA4oYXVGFcppLjimj/JLScyd4V3H
ZLmLxtswQYyKtO1c1Pl3gr+7nobjAmc2Fd5QTNNVk24ZzGgh6eFW/sjCfURI
P0Cz7z+5ZrJdrUU/I/ImlLv0Lra2g0zr0rA771ByKNgHxijA9mZ2uHufpiJ9
Uz/73uhAWOSePH0yIQ8/jDroAu1RJK3nuQSrPl9MJgfSdH08U6eMDI4OFKXU
gdPFujGou9KQuPCQDtrFkDfdWOBj3AtX345v3rdUIXkQ8AbEj4rlpCjThtHf
1xjTln6OKleL0ybJaQpXl7Xm+bHS6PzYPbiN7Wa3WArgwVuBQnTH/OijAgGr
bh3MQuRvOI91IlPJ8S3bkExoHk797Ze1fr1JE+O8kGzIHd/wOuFfX4h5HgWk
85R9R53hl41cZL2r16salntiGA4y53CMrKNqAq4hO8Szb2ZLUg9fRFVTl1wC
0AW0FELQ2COSXHhEQOAaA5SNI02OXiCbTfNGbx/1c4bFb/LUUD75KGp/8Zk7
Ws27P/wOtJwo0YuqYrOnjx59nkF3VarRyNiczyeoKh9uXa0oURgSMhlUB05A
+N52ywpW1iONNcJN5H/LUOL/eFVBumH0E8l3Wxz+/4pGHltxrsWgal+NWmHc
jg/S5rixyGWiY4x/9c6eQAwkyJtY4QHyFGeD+oK1kPS87BObI05CDLKLiv//
zRFdFvndkdtWfkgSwhXbrPawE2xEi3zwonTtwTuuNQLsVPls9Gi38xeSjd4D
s6NnCrhvXtkbvrSdzhmD2GfzevxX20LR9HP2c2/I51LOzbfo7c6dD/fRaEhC
MWUpBTamEfXMm+wOfFZ3NqfLFYsTPEZNdWHRPlcwqqBCk28Xs8dqxsKiYGN8
NdBbBpGrheJBlVYEqWwY1gqPa4tuBBY3zGGBjEcf3nrmPOQZ2hbjZJQ5fzwJ
lZfBjEThJOrn3W5U9uZERplZyG4FWxk7h8U6O5SyJHSD7bXOsG/CMr2BYYwa
Lt+i+ez/7AFWdw35p61lt4r1ZQnIFfU8K8OnxnrUfAEFAuvwbSeeWwQt9cQ6
MZsE9mVyby9X0tPHn9KZNCAwkbsXzS0kAJHEteBcTqht2ldCvQT2AxdBD+Ia
bXtNMyAqBdRLsKlJvisQE2sDwQfHQYC8mCn/Z1TfsNPrFv05u5CiUTOBtnki
OYlx2xDXc2JakupQ6oHIaUFiPcYISvIVON8oWrJiEyupZkG0hShnWjqfUuqD
X0RLdimYCHHGpkg0+Z7UyY+hZ9ajJbRDXvfM8JW4U7IdO2BJp2ie8JwS9rP8
qcJypxfA5ptXaeAmtMUu0pVbiUJ37gE53x57xO5bZGrBIlQH2woSML7KcDx/
yYo6PkAhBv4kNeieeM9t0wKkTyROiyIFs5wMGsm4DpjalXqQPnlUoMBQgRbU
ky76fOw0vMrPbyGcn9eSjisA2vfb6+kImiGh2P5ZWApoolmxE/hrnT55hVMc
xsfRKQ0P08yMkVpr3a6vsyaKLfVVCl+dzEGr2WS1YnsCHMLE9p78heR+fwyg
12sWK5Hx4/brHU7sK4Wsf+jGC0ITz2ImHHw1dD6rVetg+CLGV/wVLCTVHMsj
ByATh32nvy/9qT+Sg3pglTH7p6V99TjpeD7j/SIVHemzLYwQIy3/ETbkRpOw
Y26JkBsCyVOCNgb8rALkKXvL3fYBjc1aQRQo1viU+NebdsFurh7nq1JYsNy0
nfmjfR+mE9eLCLdcfxCaf0ctFMSrlcvEVbz8xph9Sh3l9DQMoJskOGuJ2FuX
qsln/IvkR0TuJhmjrFT8i1Y8T4wNaP76J4wYPxUDAG0fQpF5dMes8U9LEHka
jTYLXy3FYhRxEJ5hRPYYkRQGcj81oalJMsW4s/QsztI+tqKhM2EeTxTnwkL+
pq9MouX3DI8BtefXzv02eEul643ycjfFi5z5xaDA96JlxLAEHm7haKJA0cep
Mk00tG3eyyqRqQs+BziMYDItC50BBht1GMNz9rXy1iWYr9NXSi+FIRCuq2AT
byhVqm6MBeK9IzUudzd3azdnYtGLFEd5WY6vDaBpvx27dZEiMx63vc8lny6V
QjCKBnOtmqodXZbcj7j/Xi65c8Fq2smp+OKIRLbj1BFi72RXyslQCmr3hn5a
Xi9i4+o0CW20S5Czs8HMCKnmhlnssWxTWB8EiQ/Bq83jAVj/C7NiJ/hi03fw
sAh7a0tapG/a5rQGEOFFxVHWMc/XWNSzQra5ScK3Utuz2Odt7bmFTuKd9ehj
qtbvFOHBvIeRvB3bNGJX7TBpgnIwYpr3ccL9P2mO/RijU3GT2X9zXeNIg4qw
LPSpCHf3DGN0lGeJhjmsbdQ06OLtd4Hi1MzdVU+DkaHcQasP2BwNyXSvEvKE
zfG7nC3t2uFTDy78aMMFXw2CSQh5oVD94+eaFIAym8kKkllhMd/BdKjNj4Cm
WnLSG18lT7NACyelBKg4h4xS/fO+hOgE/eoOI0WdhGfGNcRa5GIcQKRMHMYY
hDu7xo37Bkld/Ypi9YxYfvHPoq68+3/57mu/bhfwWNvJHgfKCzbdSoxnz0ys
ShyR9fbEgKekr4m6liCRfmdlGdA6OeEEyYsZoVX1Win35E5e0wqYc0kxAPHk
02Z+n6uFBfRK+dThUAHw0kTw5C3X3dKZS2FpeUDp71F//6wcqzWtCZdijgmQ
zm1eYP91//QTyeKr40Ged/+TtdLHloufJWvMLGgq5F89fvOo0lS/taF34YXk
zLtkPjflAwt3dfKfEhpxJpH3dzHvfRVPqnmij2qZG/wZc7oF9P8VAjUSJ3QE
Xbgaax4caGA90bMT0Nla9em/7g/DO+PrcfD6UbA5/WsMnMm241SuvTD5mq9X
FjGgqhSa5Exh0xFgIPRgtpsWKV7l6ssAPpgBpozrOJMpx3SquRob7Y7NErOg
WwKZdQwsaTIoXtPtnG3Amc12EJGLWEZq46EHGaQQ8BVri522JymSwIflc2Bo
mzeUhBby3JAYtYlpy0hwxRcH2qfpWYlevaJgCELg6VoaFzCpeZ589zWWB3sD
zomP4niYFXERFxuhXQgZrP77RONb9x2UAq3Koy30C/L4qZbaOLkA+2BDMPnx
zo7qT3TdkG6PcaY4aJkPzGcvmMN4jsqI6Xdb9vd5W1vOxdSJPHZaetNs8oj5
yZzNB1slWldOwQT8Ut9CBB6neSA4TX8tx8nyyrgXdSpgJBygqFKEcIF5RRiT
DC2268mXhmpZzGQCG3zfvbwh0vfhvpabWUzcDqIGU8Zy2p06cJJS4dOxnrPg
nbU68yshFQl+GbUSw2gnEmL4/4uFil72Z21IpNkte8WM3uIyf8gbzDoGB7XY
VIL+imdztpRIzN5ufRmI9L06/R0O6yrZJK44MisTjOVGKQlwFQLiBVk2Cdac
UjXscq4T/f2bB3/tyOl/lUEaPte6gx4WkOQH935IDfy8i52FDAYgWVksw4Uo
D1+KcaHwA+H14YusMvj54HBdgg53ce6aa4vjIVoQX3y2UUV6r+b19PZMUS/e
XJSlqWQP4aDFADxGbDNFILCEJKA1YVvzsRebTz6I7CjMzLS4JCh0UFhDiYyG
EDvdhlFLrc76JKFLDVPeWBEsZ0r0EjBGSg/8CkrcfU0izTwoEpOb8lvKQ+Pp
fmbb2w5qEODqu3598Y0I3usH/kg9QrAI4uptmzQVFirjRd7wEpNIVQdlhgzp
4/xZFSYHkpkyXFRLXF5/IR8oHSM2vXlxkiNCjHuGakFuGzk/nOXKS8O4ZGHj
L/Rah6qPAphuwlz5493scCnZo2AYXuvVfMJJkHj9ut7nknlGJAafMnPiTOuc
M9QK5CGKNQ18eRWDk0HysxPR2StMsOUVqL08ke9iwQsIClc61za1/FqImDR5
c0IBa6LDhvKgiCd6935YDczLwrVmhStpYA02wIh4m3ny8WwM4TMJE7g/A3QH
eb2q+n9jtG+Gu21I7tn0RTgTd8zpPrF5SVjBCAeat4/ORbb4tVgJVLukjh5k
I/GWWyC2dreEg5D5TwrchMA6xGP2U8tx8Qncw4U+sGSq6hLB8k40IkJDRFMB
3fGEAg9Q8qH1mh7oENfbgZ/UEh+9jDxzt+uUjQXdeN/LfzBzsR30kcF4vHwV
1+4e5uDKRoga+Q96Zn4InL6FJY5EEhk64uDfExq1pOWxOBQwoIS4eDB+Wusx
nGrNoFhV8BfinQRRY6wburFQO8zFTSPm0vVJxWbkN9+fl/fsFn/X7ZQW7+1Y
VuPNwi+rd26FzZ96+0QJ+qgW1Ej4DVuJbS1xjV1CsEQk/ttInjP2GzeF/Js0
yUvvkeWm/d3Zs7Lq/wzW+5dyjHhr2D6JsPd02s7mN3YItLHlDqJxLgbSs1F0
cMAytm/5MIT2t99JB9uMz5CTnVCUm99qYrjQwRVnLkaQzQO8eiqqwFwD6J4P
KvRboz0cl5PTvL1Qi4XDvOO5eqidtl3qs+NhkcJmeSUDJhb3S8K892TtEDb7
za7YPzzw5a517edKvbgFwfGmXcZIoFpzbTz9z8IDaV2ND7gSzMn3IcHmfrtc
uQdsF3BZO07Ex+n9IilU8vueaU12m+9nkdAZW5TD5NPgAUSRO07EfOrpfY/j
GhT5I4h5U72YZtmmQMlNpRULmtzC6GfjNHhMACIoYpVfG6M9repSBjWr+4wm
u73eJ2Go5rHQSJr4gOQfx4MedDlRHFNMkK+VyUhsp0QRDJJVXPLMzii88POh
E0/pS/9aKS3+hPYTzKTZ3yEFZneLd4M1O3VIRbvq4id8CkDgOWGiv4fGn0W8
RzwTaYOg9IXpkiddKH5Jh6Qj8QqAEPb+bNBz1TDXLpfWUoDFARF4cNEPVEKI
1YXZRA5LFLTYbzeyJIhq9iI6lqT4LR0cwGmeQyx9/FtUyu0eskjcNo9nOchW
R9qeytKytj6SL3fgC52G4IHZJ+lag4yZy8j5NYWr2wjICfg51jwKoWC5ELdN
dVc0eDmJL8h6aSq7Um+VKAhuRfIgiqpcSfO8qsDrvaICDROsYIVeS7r3amD0
oATEHWdex/8KZ4PItdKV+tuDWUF+Kf0kX8Xg/RxCCJFd+7CZiU3g28UQPT7G
3BWNB40rJ1X/XuSDqwI2Ajc12pBvd0va56FM8CqUNblLy0sERqqEwjY0h8AA
Dnl9S5/Z298KfaYWfu/j9heHdfasZSWhmV0Zvab8NFvW/Lu0CJwgsE/bFXNw
hxu94nBBtbirc6DhsVLKun120/AxuqvUiWwN2S7zXwPOcWLp677UQ7uCF3TA
uhuCOu2TtfaqpTsIzept+w4xWcnJg4GsS34wn8n5y8MeYa38mM/ZjF0nFbNB
i10QVHcBJSaSj7g3TVJN982z5PQ67pXOAfog64FyzGp8EINLJRqv7xxc/bv2
caAOPV0X/FnY7bKePQVZN8CbqRKSSJcpPOQsDY4HdoYCT6ZCJnyyOVUG12+6
N7z5WYAD9xKddt7vujlz2Z9++duRajBW8/nQTIfrdn9OgmzRGtsYkCohsClq
uEaY5EfYedT43a1chpPOZq6P3jQYb0NW3NBwwuZHpyGx+Z0SWuDadAkcUHIx
TyOtEJYpE5hbGZFaptfrtD01Mz0XEoCoi6RVLkXksa3IPPzPeNx8hL1+jSxk
f9vf+jI7tH+uqnnrw0y1Uvywq22FkdYJ7tAGqsIYKXKIXmI3d7oASsAI9U7e
MReIurFYNMfHIxQlHBgG3L95lY313cHHKuUp/t/fz0nP5kf+Ekf5VtRQ0au1
G+nNcruKftrjTJ8/FoK5lEhWE1+A7941dDLXdmTae5Z7SRCzRCjluujku7GQ
Bdh5IUQbTXmVr0POqxCQPQUfjOQmdSCDQpX0k8aA2i/Ks0PebbEgBmZNFyIV
dC2jQjDIXOaKawVT9YVpeMNCng+0KLmMtZDHmvOl/DSyNoz1Ai1V/v6Odn8r
VYfCLVWPVQmuS5NnU7gwwnON4LS9l5rksxq0lmsQqNjp3MU5ZXhox27w9heP
g2IUeJrO547PXn5Mj7YlaNUxe74zZcoixgDaFqtcP/XV6zdoW009nUzoe3LX
V48ht3AonjBeWv9nMnw85HzyqeqqqKBmq7tXQt0M6jmgY0LyYaVgBEfjpca4
K3/wTlCAR0i39iYkNc9HHpkmQZSB9BrAgeiLxWNTfWGCU5v6fpeKae7JBEDJ
/iBq7DWgi1VHmZ4IOhH54/JPlya8xFnw2165UwDQR6YMAwe391nhFFUXZ04U
/6GavMvDyTCy3YxrB1VGea59fOJSSqqt/f2FP4gGc+kCX4s8JMME9zzxkkrp
CQYzto17fKJTKSiqOOXIm83xHzKcbYtqvrzo4/yGCs6uGJ2LB8PE/E/3VGot
O7zSVhaUvaGPf5bCtji5KB31nEozqdKdNHsuIf5bfVgls+lXfSWc9hvyCNes
u/joyX0ciQCQ/AZkBc5P5hamNkpMGxsWqRWXoEnlh79BcHuPFkhmYKnfsBop
QeTqoPEPOq2T1eqVhvnUDDTZBurnKKsDPUXuJERURZdugoUEKcpxBc3zYxYg
XZjfefX+A8LgqG5p+hpXJEvpc1eSBQwmgAj9fGKVzKLJ5HoIicOSw8viIyZi
ahHYqOowwTFTyxyyoLhJvdctEDkhbASh3vgEJ2uPPsnuVugavoxZVKxbdevb
xt1bVgMHRhB7mnIICxqDjQaFK20qzqV4qNemqxlbcgEUwqb6IQuXAzexngdG
FRlzugE9fOI1dHSy/Inhdpvj9hM4XaQp3T1MJZRFhjPw6BngUVm+MT3JwqFd
0hFkVWDc9HpErr9n1q2/ml1xwD3x1yjl9wpXHLTFTQGV907J4hrH+rIByYzP
yLVJbn3u6QTGWgY6PE28iMPawznd1E1aKvdekBM2FUU7c5AnNorTckk8LCLk
eFlBrX1f4vYlxm0GL0Ee3b/1PRsNBZr5lMFZoBgL2u89Peg/Ql9xOJazOapM
y3Xsqj+RVb64kWVvMTqkaK/5f1jpLOaazzmb8yoGAqdC9Bkj8xKSq2r5DTJd
Q8OX5welMcUw9TuY89KlecqgKYXjjR/Bq98MEWu5QI3nKQDgwGoUFbF43si6
xny18WtLNE36LHHGZYypMoRdMxbRx9LvytNhi9HPRzk5D+4vwJ6+bqemSH9E
9+4zAYw7EfWyvuQxpwuU8AyUvpfFEFVd2zo641s59KqOs0dJS4eBfThckCCa
iLw9JljcE8bCFp5Ui26O4ZGhkD9nLKtKq+fnH0i7O0WBhbQPMZaJwljDQO3b
Og8cELbUKILbPZ6Sz5y/SYZndzG1Cwld8TLDLoHGWx7jnjBjlw/Vb/PZsSo+
XOWkMvIO4TA+m/qqy2Wgp76jBddLkp9riwC2nkHByv+VE2qbpdCOslzHDyyF
/c8cGwOo2/Z2IMTV75YnvnhZX19PXmuVG7q5fVbkE+9zkIzHiF79kHG8TUaS
p0g9tp3UROuFaCUFPtWGK6MNE7xwLL7pineYRa2LctOGHoylry+w5fpIC00X
ZpqCE9RMqUhQGO4lEx7cODXRFGeK9KkkkLBhYMgw1TkYE+mX3vFXM9dEugUZ
1Nkroix/5Jb3PVT8BtisW3SnRq9aJk3+nvs4k7tIbq8ygfsximWRbe7Kbg5W
gJcfKzBPdwpSCTZeXWoW12ctT1kkcr2gEPLWkf1ZYs/5n5SKQfA29cArrz2S
4VexOBVTBEKQv31JdbiYXgYvBA//NEBvjtUgtw5bWBPQiU/q8VUJRO4Uz31T
XGkQD+QybZCwQm1NMh9T7zL398YvQuKtkXDuViBIlmla2n5zxxX++pDh9BKV
3CyhPUNx1moTERetgAS8cwuFONpA/oM3AEFUJKuApCt9fr6Jyw8FBKh28V2m
tsH3Jq/E2leKhHLGkqwJLRFrhXJ1DXIu00+vUUVG9P5qom5HaEjYUiiS2OXW
7DzEuLwvUZq+dSyApSW839JOWhGBs4N9JQkKDFgU3Zx1eahTnhQMPJVxQr4o
M/MhWTiWkTKhO2BgVyktIFqSNWPBo0FtYAcsAM1IsnRdS53Yxv4h8Li6GalY
YqR65oSCVF5xFax74gk5xiwEBBkEt56cxVTnSqlR4wk9WW4kMdcuH1rcLNfd
v8ABSpQcSH45JS/qR/Jg9i3O8FXOp/sx2nsbzsRYysQmjyfjJYOrSOD8seSw
t+Dw6/S9Wb4J+IQwWoGpTcFfSwHBxcS6Nx1h4oJz1lQ6e4gNIXqH3irEe+B2
pZXiJ5+e/zS2QKOUn06qmNk28JbJGa6HZcib2TKHXoXebs+qvZ3ZKuvBt+Bk
v0PIvJ6xNGfgqspBlYMBzgHkCxW0Q3mkwpvPs1PIhnSP/g/Rbw3N4k224ORX
vyln2zyY6O2EzlQpfilSN6ryh5CeST2YxKoAraW2rv29lXLdmvXQ2UMOPvYd
bsBDHMwLjLQQO8fGPOXELdaBky6LmAsyDG1abzaxEkuYlTxXQtcnAtIPy/AN
WQkSDJ4GYsDH8rJCRXCZ7JGQizW9BP/T3r1SM/oBnXmssglj2mgJRRmjnnJy
PRhwHTL2QcD6mWgYsFaU2vOXW/8c1/49VFGHi7/x4RrKhBcrA7JRmuluETv4
tsI9Jj2NL3MR0AiO78twSsYDoAX4hE2bbTBNslBYu6tnCMlk/rGSNUIT8Dzk
ThHpgm0MtsU8mjk/c9ZLSTpFJQQMesjPX8xIcKuttPIrQB1n9cQ9TCkCSl+J
3UFbWNnJ6kMk+/NK36iIEAfxizAR6yOAQp5GXOmnMvBcNzB7S986CB6awro/
Q8Rxwe3XCTYlVLg9ayepDWtjWuvIe19Y9FUkr3SG+UZ94+H/EmoozfAILlrO
fc1dLKP0wfeHjfwSxfU82hLqY9nvSeC+Hf89WFTsqhUQod/6tp6362Dknmod
ujBx6c63QvAcULlu5UhKAWoPamEbG+Q9zuLN6AOSYBKt8VlcNVBNzsbySQIb
RYPA1uVeIdvaLVPJDZ0+t11ZLjp1gPsP9ZeUXOwcW1rTDizYBFE4N1zGFgNj
6fJiJRKz65bO0NwVhQwrM7ZyklGcOHcaenneUid8CMdIWP3AM3XbjTRCsMsL
tgtq79IZXuf9V2ITiYIe0xLF2EBF2y/C8Qz5HOfTzDa3warWc3rK8OT9QfYe
k4liF5Cd0d1MUNQnpJuA6vVTinDygmVi1F4RrAroWqPVn9URS7gQGitgLnZx
t0ZFrIP/PosC5MMxMvgg24J9oqJBv+0WIxoaRDQOQFc9GS21V0Tcg3hbufsv
Zd8UPpaj3ljmw1upNLTyP7vRwqOsPZZtT8g9nPdiq+jUPkbHCAbtZpLZf3lw
UbioQMR5LUaC3ViBJGh/R7vvWPdNdC7t2WiQdT4PA5dG58HGTjCAYhm5dTZh
S1cUpaSY+rqhE/1uVbYvcbOAI0yd5cMqilpf6M4qx6nskX9o0XYYadmsIPde
EBZSHmFiw/+BRAUGRZBOdu6EfLd1iR+VUHoFCRZ1qU1+8btmlqfVM3MXup5I
k1MsHph+4tr7ExakIGTPCDiHwLFUSfBC2b9hDhGS10wwvsPwigg8MaKgSout
5L/HPA/W16Z7Vov+E55IWKri3+HV85ttnHlAtAteEnL13iYFd4/qgojaSN5M
Lc3inyLr5ISt8JRq5rPFJOlH0bWxxW3ZkMHZIHwVm7xoE+GQBsN3d97ymoFV
3s5StzYW1ha0gYg/q6gwQFx/SjIXTl1V0zxtEPX9YaEi+ZuRp/O22vrySiZQ
IlLnQrJDZ0f69ou/d7qir3YZpxAE2lGGL59z+1LlJizAik54T0mTIxp6ZPxZ
3Emqxct5dHnjYnGaDpVcQSDZUQKjCgPRLBOtaDTRaz4JXb8v8a1myTlOHXul
322f+hMAIN8BVIa0UXRIJH3REhfhmmAeEkTWuKgA7sb5aTEhaON/V5ZYJyS2
deHD/Z7vdQE/dq1CuINxTjcwrcsxjxC7G0X31pPfLjeMv9o61M2VQA7yR5TO
NuNlOlThtrYx3S4GY7NrEGFQiQE62jn9A1kEXY5Qd/2Z2f9QnxrdAhZWVX4j
khQ25QwriBWqdMGAO0+jzGZ7LOfA3E0FptpwfQytGCosjI0/pScNDP6eDInJ
7/SiADmqEN9YUrOC/v2sbmTRPF4Hfehee3iqFDnyOHI9X/05L5aUmn8WiTDC
B1zApdTHUHakoDFjrmFVHJTvJQYdzDAdY2xK0vfmVKd5pcIT7v+tlcJ39vfn
iwdRTi03bkfttrFLkvyk/BAN/9E3yCyjduy+WSgBEQk4QSlwZJ/vsgaWIbg6
bUynQ6JuBMM0HOXghDxRzxarj7txflH4SA4Y7PwoDETUn4G/LzQTgcZaMMaK
1V4IDGyZK8/SquPJunMeWOVI6Hl3KagFAHKgQJ9atk0966Ttzic3xxDdtzK0
xOxKJekK02wlB2AAeI6arFWLp3evPlEGxugce9NCbt+hewHPECHwE/JGLQKq
AlYCNAok/8HFpNJDuEEWv63OacerUgreXBA1nkmt3jfomL4kdoxjc3XCJwOY
JNGv7CTljHIr7AYm+ubjvnKhb+8DQdAW+IVIJqDOK6X2bS0dTymZOG724lW0
qZJTyE9vhMYt9Or9HIIKzZFkFLqG+MqnGkk3mabJKZVhbIkm4WwnWKw8Y3Hq
Lf7ovvfbf6EaN8W9LSQBkHTk9VkFSjSvMj/RtuGElg1dp9dac0yzno0/D8lj
gzZGKLbWPQ/RDrGqDxI9YeePhbbnouvydz4PhJLCdqRG+6HDRgxc0hwTzh1S
D9IGsJBefZIuEs0uNWTptROclNHKk+2Au7RfpohEhm95b6Y8Z4HuDTS91c01
/h7N0FDTBk5idgIuryqbbEAOrc/Rtfv/1mFrAMzxQj8CYpSpoI9ZXSCyUFp2
fL3qv7F9/djdnJocjr0vbQzHi9IsposlAjLclBU0jquPMzj0ikRgZp64DapO
C4B/mOqCE/ktDP8yxvLllDBF/QZv7v7BFMZ7oCY4K4b4zqlR5JPWTBEyJjp8
VuZZLtsHUxnPst62cJ1X8qGa4JsxRxV35rbV3Zc6QeetPRp4HTDCbi2VoaJf
DvIv8C+pzg7arnG1/iDbFVFcqWAJS1Us6qaZM+fpLnMosYilul7OlakCCsS8
co7TZ3bf+36iKYyBswKLwVwPswGNcH/KrFq4w57hlJypLy1OFV9/fZfKX7gu
4PG5Fbq5yTFjKhB9ekC21gMgjR7gr8GeO+bf7MH0MauTaoPqsvNJNiOAE7Ny
gIi2qUgQaX2VFgFgY8tCxXhwrPEVlOSCPkX3hu8kDlS9ARyWEuge51plugnK
VEb30BG9mMtnEilUQ7PbkMDg4uI98ItBgXTitaFkoeCBCV8F2nDsQFX8X7BZ
It/knCDD2tJnC7iDVK6/PL0GyWbi4k9crmZdudx+wDwntTunJxwF7P2qW425
JDmZeIYlXWevyVy4vH4owbzDu+aeb8Btu61EY9BFlxh65cPy3Ga3BpZbwNgr
CoKit49KOTFDffsolH5kND4M09cq8Ew5sGeactcRx/i6lb+aEQwBCqCgPWO7
tf0Hp2tg6aDZNjwQAwyMD9cvNddNX5vBc1YA1X+9YgS++FWpU+56bbMQkX4m
BKQ+LndFnCtN+R6UIrAUu9cwH2LRh8m3dL1oOJsOFNIBWPXbOaKsotOMhoEx
pzRdmiVtYPRI4yuI9GiGMnpXsEUyfurMJffJ456TjIbX8qMHJk9QoR8hB4HD
7EcnRbRBD1cE3gveJFqtZan7X55qWFuN5zIB/OeS/6c0LAM5VflRlg2iJfbU
nmCRliAAZ/zuBtdL7pOf13pC5b6phf/3WGZmIYotLGzqB+JOp9xJ3aoxzZjD
SWesT0CnskS74c5+siuDRqIWeX5I7rK3tWv5zlIpCPHNzLnPXqnogQ8+Tp86
xL5Z2zXahBSPycRRgmYsihc19pOa+CWTRWt+CC2OyMKuZHT/ucSXnZvpxOiP
oARnEEW1XEloVPZnskyu7tMqagzbODupnmE8HnFXOt6hwAM7cL/7QmGR/Oy6
bKqaovEtUyk4Yp24NRvuQ0JfeuD/dUXW2e+LIEHZML8uH+a1DRPefa77wqZ4
X3OD9E7O21DssTBY7iX3GVABr5GyLODphxZKi2AfLgWA/ZBMdggTZ0yoKKoQ
2LGfvklGLLoV+tpg+i+DnQjKSFxx0AI6ul5X1DF+1o4X2Dk85rFqonZ2PPCU
kP+XHxIefUqCoZdGj044FXRDAZWewAP00jlcPFKht3MzBqHka3b4GZDjuy1H
1MXUKqGckFKrngS95g3qxXFImGczgBsHqdcNKAMJ8Pjk5UOyrzTP2uX77XmL
9GoJ3Wl80BwsMmMi8oR6/mld1cw9BlcIKC8syUIlfr7P7n7oS0g0JB4fZZzV
0/LxpeILYO+3NmOU/laE4pCWbGFk33RydoqrxCfZ4PyKI0yElRKp8bEzjjWe
XfoaqpXc3YDawFEqDlxYhAW69t/eBkMF0uA34jt69Dq2iG8EboZRM25kXX10
6a7gG73OEvOtcT+ViMYzHtOVvo68ihC1hghD4wPmGQUhFaEcdUbc7ABjg7ua
Q/I9huA7e0ap2GzjHuC/3HtUIkvT8YOOZ/w0iBkRA9EYyDbaNd1MTZnKuGzQ
rtmv/b2Vj8oi/Iq/uE2cgIz7aboRawKwQs4Lhfpu/N3gPgHq5YfAyyjuzigQ
tvHRusD8D8lSufPm8V2S4UsbYc8M5h9trcC86vahE2c9MhuydBv5xjEv2+zx
TiUPCTkw8KLYt0LcqyWB4Mg/m/TQkJ5eKmiChkzRZ8pypJq6QUsQb0Yag/w8
LM88A7yMUdJ0sH7HHH4TnyUziFnKTLSIrjIDki9vN+U1NgrYLrCVpDEOOYMO
bmcuagCLs4sx5h3taKY5Th2EZc8yvt6I6WxBK1PxE4wm6yW4oguPtUPfieOC
rTYgWcP0stclQLuQSZqvrNCBIzDF0maKJYcrE/YwoectYQn6IkKOuB0HKO86
PvchWUrojvjjKXEx81YshDgRV+8OfczCW4bLRqfwszzWKy9R6JGbbmJpD4zI
V2Y+a0b7PvGqJu7Li18+/QSePEjZbBXwVvNXZRhQfopvsYoUzc6vry+EgiYn
JfQ9KT1pEPMAwxGIO5D1zU8aq+y9BT6Xza2ZaqB2ag1QRn23jWuge7mVFMYm
sWbkcDRglwesh2vhSn0TSBcq/k3rO7nRBNZKcBuBlWllJ5UBOh5Xq94c1voI
3fjXzr42S+ihNQiycwuk7a3QeXWTM25QnFFO/DgCaskMChfC5lZLjbdVDiLl
Q8fOFYwMIUys3u4vSdaZqmzZtewlC0vcsJUikGrl6l+v+82y8AyNZbE9eGvz
ov3azGH3Zq39vatvUOcB6x8h2s4KTofYB7V72XMzT3s7RVFqGv/hksyFJCcy
kLC6RAL3hRV6z8w0eX6e93U03c4TZ/l9RtC+4BAQQJnONbT3F2pIbZ73kqCJ
uwpfZE9aeCbDce1YOhY3LOyXT7MBRwMrEKBqora2zlKMHCUrrFtv6uMiH/SS
h2ZgM2PSuka1aIL062VmeK1oK8rhP1aE+PiBQyJ7mWt5N1y/vILaU92eqJa+
RLLrvLCeeZiPZDlnvXFMX7In1wdonIVu42BP3qqJEikrCksFxaKpBH1w7sz2
EBMDxuUNnpM2QfEQc11G1okgMnWeGMZJ+DlkZMpStDkK1isklTo/KH0tAKv9
nzxe5xrMKjTjo/HX6unCmVTZqiepxUw4ErP7rzGGsEAFkhI/OktGYaPekQas
UmrYmED3T4XkrW3M1/edlANK1s1nhfJhVJ9teyq/6gWhjH8RPtUsWvJ0ifRG
WC918vL0mD7UcpKGOEmv168ZerplAmGJdbDMzT0TAzvOPL31YsDef2YkEh1G
V53JTXU8TBODrHqSA3+27mwtJvAhEUj5IvWYaIJqIDgV91zu4Av4G66RpJ51
AKDi1hWYX+Nu7hQIlu04L9ki7uI/U54S6Uk3lxa1I9QD29SnxCTJbjPu9PPa
EGcW7yOJlFByyKC63Fdfx8ePQ/KvoPbDVR1VWvcwzrQoc7cBd4uSSmj/KGvD
59wkRfsB9Rjkanc4SJYboB8w3jwuj702CDjt9Dq2YrXHwKZOcAxzcwVTjdZO
5t4bFMhgd9p21s5JkQN0NzkTxQApmzzCxlJD6VVmGSUuoXLhCB1Z0kzsotn0
L65BHVvOf2VDQRt2tXG2vuy9Fs47N/SoWyzPHeXWqD2JnxaY/WLSRjJGvWhC
QK1ruwhfiIrqSb4eAlJJveDljjw4QUqleLbtsbUhhV0QMqvlMSi7kW+IacgN
ngus0EoYWj+iKgS8w3yRuGBf6iBbnjlXMm/I/Tzh1T5gIcOV45dCgVQyDzDs
JkJm3W1PMAFdRl+WggXdEkbdsJi/mZAoNBDVUVqw97iw+dl5a8CwEviD7Dvp
/oGDeGhyts0yk6yxhsirRJGbhNIxdmRZMpWyTYXaHGWr548ExU8ni/H0ZtxB
HMV4i0OHRhxTE+uQVqMQwjQUb07BMNDCWHkJ8QfJ495HQnnx6rGmhBS8L0uZ
yjjB5nbiJ2hGWUFDBkHZNVKzyZgciLnhyx6+WBjT5oX8rLjFBbvOAqjS1tVV
GXNWNqj/6wFC9IIfKzGDIjhy6iRfAk0CDbSs8o4NDZmGUhGIZY3M8cztEZfG
0VIWhmgO9ESHgKok6bKGvlaPfMgKB+96D8E9VROVA1z2CVh6fhvWyHtNxFcZ
Puo/LaOAMTn7uwG9ABYqGkUX9zlXAQrDYfyb1+GTwfqVA9UMnKn1eG1L4D9X
wLMjKpnlJnDT3WpS7K+aJuFEPLZMcQF0fnw6HWD8/AigGvMJMyPXaHtWtgRm
hQd08VI2lLA4cmQQW9C9KmLnvODyGASedyJfJRfrSL8Uz86hUHHeGEIdOqlp
9wfJXrWfh2WIBpD5zgO9jE3sl3Q13TX5lx/RoeenhzZWItB9jos3It2L4U4O
+CVSZJlYV3slM54uNEcN2dKpjSxw5gp74yOT46iA0npZBCpl5QxQ7t9uHfTt
OOPrX30ltIGqZqoNhgruIAgc142MVree9ihO197mw4FbyLYLUgV0EjwOD8vP
NJ9YIIttX3EvdzzEJKBuKVoYQBGK/9NHPNUd/Pqlft1EuBybykYaXRsf2S0N
7vsTFLEafue4qRjZxePbxE8gnhuZHlGLBx70mG0JS5diqV+QAV6D3B4VuFap
yzXDct26cwcgXNPD74SkG7nXpTCEO+pqJZ5LPI9pPIxVzla9roDgLR/IPrtT
Lw/+4XPe9IomZDVwj0su+CUfmpPKBOSYQsEzV41hCs2vBa5SZPbHydQ65GcE
O9cVfTdtBQqzj1Jd0bX3b2+UZDtzwrCgzqwpHv6DwCbuJ4xl39G9fhNPIUr4
nhV/I/G9oHX9b15WqJwCJpk5leneDfXv17gL/W8T9Y4Vn/RwtR5otGKVM12D
to7uHWAFutLIrGl6mMyVurFoy4aGGLKtZQBnu6y0zAL3esX/TXl9LFYd4i5Q
KFEy2L1tBJxvk3rXc+rHe0fDV64ICz1VF5di33wIsJya+wbthdzWleJYkH6Q
RV6piWIK4yQmqKnoGSULSvSopZnvFypsRFWNgqnAwjEOmURfoyKHMuYRZVIB
9MznMw02VOpple2yCr/38/d4QZI7nsRcV/kfcGgMk6p5GhXob+fZJCm/zxnH
3STerw8rOgxa4IubmJ/DwHFeKGRTb8HpISNH3ORIhIFPG/em9wTjdvWyLZH5
TnmDgdVSxGfkCdpetRLIUPdMkpltK347zywa1cmXK6FawsymSZW1zVU34Zv7
gvlgjYsOXAVwTCe5vVv7J8fYMF/x9gYwBPm+/i6eDN1xLZDSkImq/mCwYWHO
N4D8fhRyJlcAIvqPJATNXTgthTMkdGN8667BF5s4lSJAvVzZ17FO+Cqnjzrb
Tx0GZM8Mm4KmXDLEUahnQUrk4pX2IJTp26t1ZOC+Qu4bhBr4Rn6b4mz78USy
0IWrsUHVSdiK5WwAC7hZtTPxR+tfFYQAVHoOU50rY+KNua7Xzd8IovMRIUf+
rVuP4jb/tEti1ljqdnYrAjS7cRu4aKMCZfIOudN+/zrIDGlAS7xegpQKwA+5
m4DrE/LUuisekhXxYxrKzbfTipJ1l3G0vf3ViAnAqevf6rVlKswYbs2vCirM
LykAMU/7KDDtxb/IMhZ/kyb99rg2w/JyQCjqYHvn+YVU2amqm7BCWFFI6dN2
2Ly0POg2zM2IJc/KpbDVQrrm8Xuq74BgDSNIhrM8rGKx/zsuMSn+5jf1irxG
HzkD1A7ND3pS93cuXtg/XhTDd6mGh2rtm26LajofCf55U9bWA9l8rwa1bUBr
1NbqyKA0DWEemMbvPHAdQPBJQg06N8ehmuqni3ir8uk0kf5bRBZMkADvnMkw
Ll6XaEYBMebjVk4HWG82cetSoPhr1SKKHTi+2ikHzrTowRLUUGIq0tb3ku1f
XVEZjIHRvBFkf8gO11kGvQvqHttxp8niP6zWVdy3m2w9PVyoa3UZEn3iVvs7
a3v8sZP1vBWEUBUS912vlfor8mVIzzvtzR5CyIfuNKs0lCywQEj5VujGWdVq
q9ZDKLSYZld3CJQ49lX//cNMUI1O2nZbKEC57mxFKRWxUGZyj6THXMH+H53B
+vu50gaZU1J5Zjol3QwvRibqDjwAwM43OHwZE02UTDMsQEdzx3XiLmU8SqEe
2CnB/Mb6nkh/RdpT+/LWfoLmhePmoNt0kGpmM/YyaAsdlrF3zHHbASSFLtpp
DbL1m8S14jJv4JtEE3vf1RlWyEFYTwmaVLHeSvdBW5wX3RHYD4EzWIBJootg
I1QQF5EeNLKCx0fgNNjU6ctJ7VkmcW+jCnVy2JbJJ8JKl2ccSvgLzGmwSUuk
xi/4DgB0zvQd5VnhlfCztNIY+see8mXEr0ay2RKfwaTUteWqOGdmeQSbgCnN
jnXUkha6vTzapU84dPs/zbE768vpcoDY7AS/SVotcoYlkXyvqmFTOYE8ovf5
D0nh9jZrbk4H8L1iqMJDWstW4srlFd9M1XLm6FvQgsbuodSYqxvYkEw72zYL
skYhAXSmFtEk31atdYT/9SoAIoXCyhiF0ESuxdKk8faWyAo3tHUL45Ep5MId
QDBFDU3yWLjwRIa/shWtm9BC7EvTE59Sdrqr4imcy1/9Ir5rbzV7Tyjm0lUy
jwv1RRNKfo/NwvDN/XsA290O7TTzBkyoBWWllnhp89BOgIeNlJJVQ4UvHb0x
iDgFw0ZGUg+xHSfHKwY5k9q1rElRIXdA+lpgWgQwAsr929F7KYTfoWx4DQ2S
qVL+mWZjRKsek7GskLUVAg85999jPJnXRwy9Jky8iefSo0SiaR/ZmfaS9Etj
23fmRsKprlRoMvhxWr7u3w/UXSZIExaFze5fW8Cc03tFsJAaudRDiuMjOkAP
QrYpX6oeDgYQ0dWzSO9KVVnhpTMqAFET7XdahXCOZgTBafYReNIun5TfCpZ2
3WmpiBGTC79QvdsJ/hJhwEMZaZjmlLVyXcCZ0eevQmLUgAxle+UoI5nl32qS
n1VmFn14+eK2eqcWUeRqgP5fDGGPBxbV21TgsAyDdLxBwX7e7WnpqyJzzf5b
1Nm+C4aaMeQzcxr9WODjt31iHUGDY7qaEmWWtlriU710NZPZyv4nr/xL1Y76
u1McxXiowrRMDqOSiZQz41vMncLs/QkdYnPu+Ra1RUiYQgjiYJPyeHlEjZ8o
h0MZVHGsHqqG77Ib6IzW6vIUvw+kXfVaEnGar6YjwwKVE6h/bRkzttvxDcIg
9Fot7X6JPG/S1rAyWGTiQFGaF1gCumewOw8P+z2O87EFnavcfqRA4jpFZ6Fw
++UbyZFpzyrWjE/z2igwo7fMRJeI41lXMofAnbuSPG4X4UKU0mUla4I0s4Q7
rDGsqNYpskMcN2j3FlUlPHj9dsDmIfuHd9c1gQcmBcGWgjK/2Hr/ONKn15qE
pjC9PVliEHYn1sC8hmoXgwJWhV0wMLfLG0ZA1nU/OawuW+rlC0GwEIi3P99T
sTthUbzZjSPrrSEvZWgi28ZAGDkgjGga+pAsA8YzR8EoLpu2KOqQln6zvMEy
ytMlDOastGVClEMmLaZMba/fkvzWbM+aAnbP/cr9+GvkmprDEOcX3Sr5Agml
uxPPQLGCUkcZKikF9ZAsp2qxUMxfZRcr6+xLQOofwdMsiXPKKtKvJbv/qyQ+
ERD7aglOKW4s2ZE5dces0KWaLc7CRCyaX/2Xo7N3ZW6VhbtsC9r4beAPjx7t
5vZ1sJ7u+hJWJ5L0EY4jNbQOcysELkOGBYmIDna1023VHnb5dDub6sqz5K43
T+eaZcSUoDNSt5unVPmFuWSloUIXuvfdLJH4wMoLRnncj2UFjsqni+3z40mL
t6fPeujbKi1TFB+5nnuhrGVNf2SABI2sXCXtHR410BW9rHyoCHW7SXSojzGq
wgp2n5h3hY1fcdxwGTAr9kl917W98Fb/CnlKC2aBvatlFzSVad0Z/JDuFO8A
uoOkhyQOJ3a5o6OJ/BWcxQ+/J3UEpujZ7T5T25ALDQSJ3FRydY/5W8Eby96c
VsSr7gvaLeCWRd6/EJvubRBST4qo6oLQxJQD3tJgkYl4z0Rlg8ghCZx/U2TT
+DNYRsm9yyFx6zn+CTY/Ktqd9BqlrRgGeNL/8ZtC+733UYS/2i10nAnooq26
Roh/UrpPCQ4/FaWVRzpwxgb+sTQwLdZ7kMkbqt/HMTFRBaJ6BVYvoOrpoZD9
v339MBH5lvVuZ+MYdQx7ZIeNBfrHPwgsMiCJzBmrCnxnKJyXBpXNLJN/xnsy
Cs31PAs6P/tPg+fIXeFxMFQY1hFxErSW3Y8fNcSS5l+qKwN7xf5NKNEFt6Ti
lymBeJWWRTvoWPFcyCF4/9ZYaU98TNGjkhLQtCOajTmlfLx5jN1NhjvEQTWR
r3rmw5SWyvE+PHu6aC7F3nF7YPZzjol96c3KPGJEDs+jKDTHhB6Cy262U52a
uXXQ2YECYSByHta060miIfCbI8HqYfTBuOxQcFRn3w6jSAVLXWGNm+vhFRSM
jvSfCfabypwwPT1nV5i2KDGRG1lBO829xlxYpgSZzU0xapGWWa779EKzyEPd
c0bMrJar0qtSjlT9q0mwC6wCQ3t6YUoM6uwp+OTbLP8dpDJaJbSmySOBg3No
438C3CSmCGX8RC1yGJ/iojeAobJyCa6Z8K0lQ4GUVUHeQyImXX9AAT4reDv/
92r18lbM84vyV/N0NVOxxCBvlB0T+RsipzSHNj21mWq4VyQcUTvQHrGvrdY6
nCAadZuixdyl1bthWhGmDvLMx1YEkWDZd8g2tF1nrcEnZwJCKLZ6JM81HWUc
VNQqPh5kPh8zisXjDNlk+IsIvuApy4AzFQsuZRcsnN4OvNJS8A2wIKbmSiR3
I7S4t4f7T1aLvoK58RHlnRc+lHyq5qA2bDQKwUREZt0htYvp9LW+1AT3HgAf
/07Kbae5p2yvscZqJo3gRauOBnnrqZjP6j6mS3P8+eagfsMlaewyMLhUeCAy
t4p1e4ztUkKLKKWg3Qpg7WWLifkKi+uLX2xM7kFuaM4clPdH9UILIF5jfJEB
jKfM3yDpDzIO16wNUtKe9J0fwHBnp/LVO5rZceEusZesPPTv5N0ZFCUt4B5b
Kkf/z+aNlnXzFzmHijbdwYDpj64cW0RNFm2CKyTRjnF6zAo32eNMqy3nlOy/
qshuEDCKfDEcfCqHlg2wym76ug90jWXk0l5mCltYzADLhMGmt5DYVw5faCDr
HdqnURt3lzp8H/TQ9PPHYA6HR4xcxr0uc/rUelyTfXINXNLK9ACVSBE4rvM1
8XvIuuc0DKjvoZPVAH60giwuFb0RpFlXHo8rIA13AQrh7Cnj61VFY4nVWiLN
B7a3KWhlLyP9+I9tEizy5D87ac6IuunG3saWOTve9voctYIkg1cE8qwRViFO
Hp3hKcBnrWvCRsPs7ccu5PaFUVhjHf5D2pWMAhkaAtEWzMYmeIWCvNkzPEC5
mcRfvMslJZYJDocOBCj6WjOmDJcItzm5/SaM0w7F/pE862dSu63lVtfBG7Xx
NzvS1VKEbHcQ4KTed6Mjori7z05tj/jrwJBrcxDbMVMypw5HOxCPvblqN5Nh
qq8rXedQWcaN1CadV5w8lGlTvPQbF0PiR0be3MxqANRWElrtqxkTexOPtUKB
A1NKP7vJBjgBv0VHqx7hS4xG6DrpPlJvPkEoJ4VbFGcr3ZdK/tnG+Qs3QnAQ
Ma7OSYqNdsr3ZxsO950HVOKuBQmYHO7v4NDFJOd3jesixZrnWcmRaoE3x/73
iF2/Ou60keoPfukUJJujrtCFta1nN/v2scOJveXIvHIgnPxeHvzDp4Tt1ftv
XNLiqyUc3+cFpeqA8E4yIGroH1bi09FZL/yabG3M0B90zMnYq+B+nM3owORx
S6CCDrdlzZYXRMOmLA0ijxMrQ1fbjVuA+H7J9VQ2Lm46K5bovNBlXMi8vwIa
315D9w3oMmNMlcxNYShlUvY3flJl6aqayjOE96M/xz+Qnzx8NkesXkg6W+YM
ItNXHC5yhUOe3MknCieNkwrgX2lMAIYVqJwK095u52ok29iLHYWIkZIzYdDp
KUxbkq2G+1Qpt+ohg8hXV08N9NdQKK+7at5uTd1pUjIOWuGps7/6lsIOTPl2
nOU6H5bJJzZxYbv9dzEuCQiqBdBq8a29fP605txtTaNpEZ1JW7tqe8RrBssf
RqRTD6CV61o2cLvCzprMbeJyjm+tSe0WA8Vjd2jPskoSoboLz6N7LgWb1PY2
/ItgEYHlekkN+Qnigb2n7M1D+LTgAU7V4/4A6fNO3/VIPLSpmR/iQXvoUXG7
OBIohHIo7K3nqrk1Yp+y3ZNw5M3QxMnQOxrpreQLYffSps8q2D5JfjDO8STN
nssix6LjXALc64ZQMm8Iw3V4RBEdfI6w/uR5UniSAsqZ8HseWlf1dfOjwndd
PG1FAD3bxZ9RqlJFBiKmYwmg+UMTKieThSb/1wFOd09A0xxroW00gOzsfUet
2dUS9FwbB9EnSbUsTo2Tl7ZdzbCVteqe1kUkfeW3I6WFVYecyZlFV1mgofSY
GFJRy0mjO/8a82NwgoyAKwqPSCo/xg7wf3/0g+vpdqa/xq+suAZBWDRZLI6b
ZZZilkpSiY+QGxGqmmbNAavkJc7dEgXDTyuT+ZIfL0Xx2Dwzf4RjZOmIeqKO
om/uhB7N9djgFWQ/ee3vk0/XdBsNfIKPOTZ6Yf8ZYpLEpgGSHoOu7fCK65Zw
Td7GiNN1pkLe+xYZNpxRXUTAdPjChVmv7YRL6u6Au+b6ewGpcOZVyz/FMMJv
fR3kuxhqzrRSvPGvIb17qEH0l3JkD6BzytPxR1rwy7/ngP8DIP6i0SaU5dx4
+rXnHiD6mQMrDP7LsyKaH76O9IgdtmJ24tZNYk+nu/ytFS+9ST9ybOxeGjYr
outC5JF4wo1gVMDshH3rNZeWg3qaxSBt0GcFM3egfDs1TsYpa5ZwUAq3gfA4
25sngwFJ2k9IaMAIE3hivcoVfmNLjicw6iBulvOi80HyTx3totHhXchFIIDJ
LVj60rNcsBAmEo61G+IHz6piZnWwl2Dty1PhYtVYlePrS8WyrvLJTtZ7JFdh
AvX07AiSwsH45UfxUSWXuggq4hn5SPKu2tCrXScCTUcbUJqD2dOvfeAS3rF1
+IDZOuIsilWZab1TMum5x/KsZicY1uFcq5SvupqpuVVX5mc6dEW/IE5kq2tN
K0RPcAp7gAwqDz5L4ctW87p77lpid6uYVNovumQJFCA1hv4iNVGCX5LcVg+k
N5qX+VJgno1OFJvoAbY7vVnq53cIZK3CcC3fKdBDQOjy4cIJYtex4K3T3yEz
Vyeq4HAWQ1IfV3qJspAAOunFpEDIp7hS+8boOSxn5jPraNALHGkKzENURJdw
A5iZixDDi1PcaQsLkqSpOzpZzcB3PoRJ6LkOdSW2rnZPKT7lI8eSe9fBZjem
PtUiiBFdTuBR14q/ez4YREndRhQ0ckkLTkSzCCQEo9UoEdGjrqnRh9W+0ywA
mNKfaCC01+slX1+8qaKh95bDpiN2FRAMOpTWRfGZyOnmDoBxVOgv1ORsOtRO
bESvcp1hy3NEIiNFUoYTz31qb124OdzgC5rZlL1qqljBVpfIju0xEHqB7kuu
O3t6vEGjUD0fCWjZ330FXH0ha+DW0vL8LugHil+1BFpQwrn+eHrvJh0gqZ9a
eOdJaQm9sjBruF1dZzjaGOiZ5F04uGtcZLaKkiAGzeDWoGAwnnQusy6oQCgY
pjhwQn2GwrpgHcQPV4WZy34p3cXEaFRGxP0T6cPJcalNWAkV2uAtwMRjMzOP
8YHIueESPAB0Rg5rOpGyFhZNzF9f3ehSLg0hlrQqoumeNrPDWOYRBJU0G6tf
Wg83kHwe3lJ8ZryFaQVlbiKN9opXK+1cwZhAQOVac0dRWpbhEdBLPbBE1C92
BSzyFt15mVrUkTZkpSyqLJRNkvh7RhcutMqdhee7H1NAfakqg698TRNy3cAJ
ftfcub4JwVIYujESeSykpk7i+SSXyLtYSrA/o54SINLS5a59UPOgZWhQpxai
Ld48ff6WxjAd1an3gMozCFB7ZYodfkTVcYBwVgoRvA+psgXScNxBGrAdj8bk
yOPJcAeb7Mi4YT3FQhIcJ1XwsIHf5KsGFFPDKq9o58ZMesXNn2o7NFk3G78v
BFhs4S60NwyCkJ9ShLfYbSfZeVK05h6vaf3mfgmgUYXQo4K8yMwl5c7j9hS7
sAhsPM+yCrzjKj36AFxlrPbPxx++t6j5pp9x1GLBVv1e96Rr2DntfNfi/tph
gmOPcAsADWBm3V7DHevhuVwA4FJ8e2ST837izU330OAoOVBJFPnRXRFs7koF
kAkHWj89g49Ukp2F7AEv9pqdZOvNJt+rGKQNtJvGz+NO2zDWfrDn1ygZOLHn
jyFo89oTAzcCzMxvW5IHuaqHCi7qBvGBxtxbimg5xodbac+h9cgK19QwXrNZ
gsXMcFPzdsMZGss4hlE+fvg6gQvdXc1tplQ7k/PWvoW7XGtwFraHVToBpDBn
uDFoy6X+y6CmrxHQD1nOh7Lj3JPRxHh1Q3GrB0PEmdhQwccG0xSgMOQszCXj
eMSO8Jv04LoXPAjCk/KHdwx2tN6ykMBN5N58wqYuuHjLKmGMSCuntt+1IZY3
3STY8lK+ctMGKttpNt9Azxaee5mSw7AHR6a8xKuRNuFhJ4vcCtQkzgzzjiLQ
0XQvHqaEtBM7iyogIvijDbTm9yKYQXpu76CVnrv7iHwUc2uVemsO7Iov6jji
PGx/UfrvMYPWfsLyaVTZWy+jI9dMwSUGqK0fovMxA93XrA/w0Y0DAqOFNiu+
EojaQ1BysJuI8jwxPOW0IGc+SofbQTcDkKyx87XedgrQZF7QBuPF1XwbvNbi
WM1WZsWwIqUfpIUVhQ/9q79bDLeI+T/3JPwdFW2Gw7hN6dJ00i40L1n8Qavj
EN2a7qcnvzWX2Cm5vyjPnlLDwP6pJCwl9C8NAxXdEFiRq7e5UECltuqnUrQD
9iDx9w9Qyvy0HxXDzMgig1jWkuRA0O3L8Qln1HicfiMTlV6ywguVRCBZG2rl
/6d6xrCo7ooPn/ws3KG3xWciPkWZp0r70FoPc8fMUX7k4it3dVNeDcD7Olpm
hVmLEzxGKTWtqJWMoAcs0ZC307RnzmrpfqRuh7WLR7zb8Ds0TIPDEmdWcgX5
wqLiT9DukdaIsTWOBeThgJzDAHSGFNKmyGNW/eJnO+oTPOl+oqGthZJpJeMK
0cV/rufQvY9FaD7I+KkuV7mwAPM1egsYTJYKfiFvkFXXlIBMGMQkHmAhPs+q
Ak/WdbivG6K8M0bX7SHFekQCVBelknZi4XJfSqQ64c7inOkeMhyeIB3G1RR3
91FMR5fNfzA1K0/dlkwEyAgOj3iPixy5IAw+HIxk0QzrluymFvIYChd00YEZ
YIR4Lvkcfw03xHOscBI/4fbf52s8gC/GdSlDz28BRxFZwHWM+EkpnKmjRiL6
BZe+2jaI/8r1iv2Z28qpchegL+DkN6yal/6wesFyUVCeOUdz1ximgE3vxTaf
3Ln1XGAXkCR6H4bG0R9f8rC0rIWe8a+sBkKQnp+jqA7B3Ua1kelyj3wwQfJP
fUJfmKFi8gkXyyTWDLp/d2oLurzu1/SAZHlvuDm7KJoPcX+fowMDZ2Ui9sdX
CrtXAvw6/TDtYEb29Qo89r/XGl2inIhgv6BvSzpJW73y1E6dEwzVjcmKZ7YS
Cu1P5NaQG6Ej3f4PYnicQ3JFFhZEagGbib1zm5mNjQR6WKeNen1m8wy9gVxQ
UgBo0MjeZ/bVqWNW+nCIt9eq5PcvPcuuW/fSNatWQsl2kB6u2bAx/LcRJCoa
WfLS2cDzbDAcRcjYYujP6Zag97ConJ58C659cYFMDkWv9czQnSOla1qZIDqR
KDH/yOV0r1Eu07MOdhHDC6yEF67RQq/KtJzgHN3DMyjk+SmgJXZlF4PNooQc
6WMnpC3SNoxDDsdEi5/2ORbJNHVk28sINjWitSCm/c1x3nTSvUPviEIfQJQ3
h47wKxU2BSGKRdXzR6pRvQ2M+olj4N2iZqMpOIizH+v8RAzcPT9hC8Y4Ih8J
hN5GxEl6S2uwPXhy+GF9PJlxUCMTc+fkFhzjXMUY1W90ZqrzNGsMFx61oqdP
DmoNfcou4ilHg6ciDoQ4BU2/Kxih0uJEvsM//Pst0lS1w+vrCscjIdxA7Ur2
fC1/pRfT/LERLJqyLXlSQfEQpetb9DatpvLhx2lCPaLXYeEnS9H/RaL1E0Bw
2ywXEqDi5MImLqj6HAhs6ygnLAh5KkBo91A46fwNrS5gI/odPkbwDjm1BGQl
ObsxgtHVnN2pnpfu5id3BBNLc+mhEX0uO/5QeuzCqY6qgQV3ihJq5MfBBsCd
USlEnHTsQWLfJhhb9AbecYNw4fh1+t1IbkrbX5+HKB86avZqYyC19iF7Cuzh
AF7mPs+/WJwMdZ7vL1pWc/80RYxs64cFN0mZxrdKW1wtvDuH1Soa2QBL8/y8
76SREd2iA/1UwWfNLR/3db07xdQTrsmOCYwYA5ME/qnAGlHoIOpQtxpwmRz8
5o8ftigadMv2wQu4ATUL/QutdFlZY/MW1kKsGT8wyFAipFi0s2KbHo/vaeG5
VolbglpcDnt4qEV5xnqdVeSopHsbRZHFMQUu2WGC/buXkG+KnRs1MPLYqfab
PDyuvXApoXzgWGZaPE265OkG5WhfQ1oMWFwDopw9BtzAlspwm0rsS68gAEz5
mZkI4BJEwy223dUJyPfX4HvqWyhze5CGOJjxkGPulOelcIjvgyIEpHY3QHXe
mSjrg+HevNpKLetBM0w7QXP4FHzKgFSskEHXphDeuxZDF7fctmFuzeAM0LU5
zn7+dEdeZ13U56psCIqXRi0DLf79FGJjqjO6cJ5wFeZfXZEpAJgcYhwYFPd3
so4WLUoU5FLXjy9l4iFwwtDlA0haRCv10wWr3Exw7gMZjhshV0z/xtcX4or4
Nd8cgRbH5kNVb6Af2BvIvar8OcnKADxJvf+i7I+rjMZqdj/41oxOpSNyh0+1
FdY/4uQbRvUetWGnTPJadMyVr1658qpNFYcuORaI5qIvFKbmf88+90q8Ox27
AOTxLeKpFDwrG1r3xH1nJ33m9Lj0JZfh+/7+sKmq8SPqhO6AxQWRjhM/k+b0
qk6yaDAHJVAc1cyusVH2pGhdi8GJCytVCFgCrwEhaBujgkxOrbdNLHr+6Ju5
mvnxORRd3+XcCcf3xCsdnp3wRyTWxHaC3xC4QSXcR2C7T2J8y0ucrfP6tBdL
dFPyFgXJp2sTJdEa5vM1TZ9eQyAXb6zr66FXFHS1iH0ENi0qy0CtsF2FCSs6
On5cdeVbT4Yfksb9wVWyTfEzBjURmB5DUxhLVdnvFSdXag6NvTMD7mXneugq
Djf5mtkidomrk+3UMeN7YIyt/okiB0558ICgjOBKKWDRr/RCFNGv86CATfrw
JMgjQ9DA1PFEcgmwa1Ldpxf8+M+CIunFofiQNJb6TExGwADYFc+FoyYg7N3m
7jXwpSbjivt6W2GL/fRV+egysixTSkux0hQgbOJuod8fv0ypLdxilSH2yFY5
7BmAzl2bdk3tAWZx8jdRWY5cJ/J4AJ64jtgGKrckds1bHIG5mBjZHj2BbIJs
fWL5KYlAW/KQjuY4kUEFHC5qgGzeqxLZpJ19kT7z6FuEFcBTi9oSfkGRyo1j
gFlFwaKE4nVKc/3SaOCBWonhf1THR/1C/2zwUKie31/SRXV3WYzAKoZ7Dy2M
dfdKHSwLyzf4gIm2Z3H6dvYwspUIXTw8wMB49CcyurOVR6FSILlw3+CNSK6r
x1wxah5YnSqiJpzUb4nGlNuRAQPZaPHlVutcp8Ojy1lRDJ2A74W3EhXCS8x2
HIApaft45K5wtNQBUOpJvi+XUaixJ4dgxZ5qv3rxjOOT/ZXLphH+lGBjIAxL
0j3CudNG7TOIWMlfYxC9HW7As9el8F2IgZE51MQlzvtu0NGWgRTeaIzq5Ah9
EUdpA4w0imFG7RQ9XxlHX1dyoZkOqCBOdX/hIHtJzDVs2FbzSPeDF991asEM
NWzNcM7F2HWqOV7Ln9HaiTM1UZP+zuWhXqFUzcRl97aVr8Q9gRYvmiEth6bc
V4PyGNfCTV7a7AY09LxdEyXKlF53b046+64bHFjTEg8cUX94fCffPG3+z2G0
W1G2KHMoOg1hSazJKfydzA0p8ic+LMRMGSMWT0e/taWYr3JRSmLVpnqKI0jC
sa6R8A4LRjI4dUPLk+4leBXEZ9PYd19ypryN0JdHxpiQP1YyaeT2AtT4Xcyy
6HFwA3HFtSBfZTKbzx/JKUR+AzItEvB+0J08v1ifC7WknNACL8O6/G4mp9Cf
YvLkA1vrHx8m0BmRYRjOuQhKXZDF4VS0HTUi3qtveW0UW2q2y2kXxOK9t1gI
xrBkIred9PT2uwLaglZT1ryU0VJyG0wg16A3CUk0wnCVVq1JYqyRI+BjV0Kd
9+OdsSAwnO41uutHJQu3uRHndddRjrGU/pUDgbbz4bKPDid91F1LdUx+H0Nn
HnZRrEo0oM9QK4Gi33SbiCYPVkNaTmY+yXrGRzh3DBr6v/IShOKrcHfoIYeA
L+BTco8H6dOZdIi8R/kF80BM0K+3BrVMKwequMR5arGHrbPUD3TXRPf16yo6
TKwAvvG8nrJ7ZQYXD73As6vlXmgowvqhrJtfC73HUYSAyglHaw+vJMUdo9V9
I5u13paHLyRq5z76o7NF+bO5NgPbm83WfyPIi9OMf3LJ6AGrSMAtITlboYo8
D4VdQN2wCIfqr4886Oveer7eDAbUpOZLLA7jTHKqdNq8lSBA9CI4kyca/dxH
5s2l0y/Y9/nCcxmqJFNDV0XQVflnKbYrWpDEqhZwp/7VMeUTeOPhD/HZk9Md
d767FVu1pSICkua1KsuzotT/65NtzjLP4LC6jFanZavJQ8MfICvBDzhgTW1D
FgErl5SyjevR+GfIAr5TMIczdGf3aGl4vbRSoMNfJDH4XPZBEDS4/guQ/15p
R2A1i2FVQMye0Bx/5+K3bju+F+0NrmXFRT0em09/xYDML0TImdCARaXFHWp3
xXBeDQcDnPs+r1U5odf26bHHvhMjNmtTV+X0+IUj1iCrIWiwY0NtI532DI5C
wkVD8KvJmK/+oFin4CX1nN3lbZ4kyeyVmc4Lw6zBkYnpXLZsyU+pvHR5PLDk
uAcHP6Y39gLFK0VQCJLxQguSh+LnwRMto/ucKMqKtujC9ByzyhQbq6f/n2AU
gnjRhySVBeV9t29uqhQ9VZ/kDd+htdgnmPEtA9ioxUHA0LiW2BcHFu14xy/J
TdL1WbnjsXqGz9WFKLmmw/IqLL/caXOuJI5fy+zVLLWW8gMF3keQFJiWOgoA
Xe9FGnh1t12GRmtOcfBOdIEti+6PJ23QbEY3M9KGGr0j5WHAMjsMDtpKvRj5
W2/j7Sq7A1HkJ33PzmjAsHom+3c2SYH0zOJaMKcmLOT3QKk5EBs5WjQb9cu+
zOGJdBupRmmbF6DO/ByZZuHf0SgbJ/oT/0yde8Naquj6DziK2UiYSDVFa14k
k1YJstC0XYuBsUVNu4vbCXvu2ewXR0S95L2JXS5XfJWUh6z+D09SU6aZIE0n
S9+BqR99emQL5JCxttvDRnXofm6tToxZ/3VNs4mjkV2obnpjak2QVuHHhhjv
GbU2li0IMmablDy5jusZmsPvbIcToq6yHzeNf6G5yRc8Ei8mWDqz7G0Risej
WPMOL4zfL/LRbuiopEh30kCq0L2/uhlCWmTRHW+/0fOmTvU3uewe2gJlDkt8
C7JPZn3Ij+InRNLx24pRP0QN2HA5KBKf7fqwV1urJkTJzPNCUAhbLXvja68I
3I4uKDFC9M1OXI38RqOWVkJleNKsc1ytYAmtHPib0XVoPRPZwlIB+lRpBQUE
kGlg4mMrWHiXknXxKJSK+g2yI2AW4+2cliNF9L11IJBabq85Kwz4d2LqtKZk
tI3S/xqog5R12gKt1RMbW+qs09Bmjs/pHOWwMUKk18zw7j/B6/VFksTcjvMm
/TFuB6sWgwdVo6bz8HdOoU2krDgJw87NaOEtJxhVl+rcIRkhXsaj+lrvVhrj
QVNtgwFVTDdlcETd6eL7MT7F+NwFKgKBTgGeQ7A3InPbe5o2ysNT3KeVMrIx
1erqM5nqK1wwJUeSKWyLMYcCZy+ru/nRR7rOAXiHPaFlucsopf+IuihHX9sb
+VP9zZuzhz2IpKUb/EYWeZ9JzBA4avDU+NnBjtb4vBGbHfVpsjl6/NfQJQbC
aPrEuGsT4HoSxY6psT+LcDufhnozMb5vzmUC59wsB9UzzmcKbJuzBLQKIYWk
zGwgaDmX5QVjIrN+p/sCkugEBXB4LQhE+ubv/IM/OfS4aG0dvH11ahphVy7A
BglJXw3WTr7olewx7QKKpsuj5pxv5pg6+zKJMwMmx78i/bUH+M2WErIFc3QR
hvdZuaEX+Zmj48ddj9oyQuwRJlnJSyG991v8ff129ACyygYtPlXSwW5KfjhS
eltjgKfy2buHycDH2kb9tHRwQLBw5NJRV1vBRnPzC1Gij7c1cGStud1fNssf
ANxitl6dieTIiZ+QSpz5nhkiI7qtil7Oaug4z9hVr+kVEWFm+Z8FIlkwEtO/
VKF5Mgt8PxO/8gFGjI6jEU2ScUQXtC0jGEMNMoEIm7AhugrjunHXtsV+JcKW
DRONQv/FlAKgRCF4Uw6UqrJvU7m00so3qm/bmcesFIQoeA3YtOaTbY0QtWX3
D/K5kUsLWFETKXtTAjcn1/EVmGgAQaEGw6mrsMx4SdjGLXc3oVKQss3sbapb
ygjaYUnzQTD1WWQjYTWsotaeuwTKCPxlQy+7NMI/iFv12QZfkGAGBH6nmQ3e
vRxCHxjSPAvDyLgQa+oyrS4f7Y/uNBgLWfh+QzymuWeoncW+TbScqSZBcujS
g29seeOAjKQypioXJepTYGzCoM8FcUV/7g4mBbEJUjB4DQfVy9VZaBQS+ZfO
A6W08S5vCLtGXCJnMv8QOQbTh40TfrMPQDBQRLAYe5uDcJyLFNqmJrRvx6Gw
/xgcjUGh5HMcvbwX8AzB4iVM+7xMjO8h6ubM3hCP0S5T2r/yvKElZk/td1jR
5VAJRNhk/Q7kSiIvLWFoNuZ9Vdy2/xyhz0/Fod7QcK6T5Razu1DmBydFTEhs
KZjrTT7mBA2QBEWlPyUAQayfN6jjPi/Bnb5cffGSLh+9L+5CE6Bi0oQHrZxN
5UIpQ6/kqy0FczE/9Wj9sMwJqmjjws9Aprfhls86zHw/FB7kAAG9AnM1OePh
C1NDjTZkPAqjrBhOTSDJ62zGm8Zp55SadzTlmKvvQCoWEa02QOmRBgpzHBeY
vwf3luNx75q6hc8D5vUxbgMPbdF4B/SE3Nwe82kCcxhAVqYwQVKvGtebeXAE
a2CtUhatqn/FFYsa+UDK/XANp0LiWEaKXnkKUxvLEUtavNax6C9HffCiNbZ3
eAKV4yhDf3tM2gW9lRtijDBHgaIOBuEoQoRue0WZ2MWA2smscyf4uWsMYhZN
/mjAvrUmkYZA2nSAvow4DbRvs8obDGECf0aF5xLZY50Q37Wjo4jkURlIh38R
cC5ZFcrIfiAlKZYFZDbEF1Tw9tOKAZTj7j7+qciJTVs4KKJQDXJ11Y+iVhhR
LtLr85vuueuaW2qVh/0KX5xP/j3lKEhMWRHvj9/m1VuCOXeIesZwDlbj7NUA
gqKyOfEyX7IXrS/BzTzr8zqMJdhwPCSqDeKQdyBfLf50mbpVcNewt6flyt6p
sJLZyvHL0x9SPB03mRP3RcZSK6BbQ2XeVLeLO19gHuLGGyA95Upo1+olR5K9
35XAwkctMN9+YahxzKIpK1gq20ops0oK3ENqR0f0Ikny1sAYkKZwD5wDYWmm
M9w0Uo1TdQ+PRSu3/afSrItuU6tzCSKAP2aiFk6AiNdHwQ4kdF8r9fM8S3T1
LWLsCZw9P9ziTPHlz/xHbWDEkOlqxFkfuudNIdQa8Z8gZ6G5c6/nAQVE1MhK
IUh+U9UKTsO3f5PQmgC/51DY8lD27W+aOYgXOAdMgnQbyJ8WNkp19js9z9yj
BJgexZjRfIAJccvyPeUKf6gBe3bJinIhTIOx6wPBgBIG2MZWwBngciZylRE+
/wf2NHayM0eJMQ7fk9Ew+bNwe40pXSNuLP7b0F+/HKCqJQTSvsMrN/wdfNwo
A7xLvzVG4MWFmcN88XvAVS/YfhUQ8HYPVOKxQNeK+E4TLv/KNy6j5j1kIVdq
yVGgI+7wvi3rlbff6yb2CWWDb4Vbt/OzPYjNY7GFe0rsOGGxQZWieKvb/rxP
nWAfkuR/6ilOUN63SAdvoauYjUax8vafiLJ1wRP87bxi1V9v3vi/edgiri97
xwx+Fp+g1p/zQKYAoFhgEQ0xfsbaA2wGCZWdxMNSXOV2azKyh1EPnebH28vP
VPYbhgOqR+HJbOCGQN7X8HlnmO7pEcKziyn9xVfoQ296QuVtz/x2l8C1jim5
ET6+mvUhGosDrRaVSi3GgHknSJAf+ulOz7GS6y48Km6HquTX1geEl5zXjGXv
X9bdxHn8n25Ke8Cuc9sSna2C83xntLxs6kPsFXHyqQwZ2Za8MGNRFWYyUHMG
V2gYry8R0qP+T8UsFV5Qw1WEfF4V7FHCSLOmsjOP/lWy4RJBgmAp+1oH5Mf3
tW8x2gcprCxNVd6jtSSDq/q1phvMxKNV+nXvKRCQqq6bdPwOGuK1BKq9ddSe
Soq7LBJVUIH7TPLg5FgK65luytiaT3LP6jN8iztvIGQamGM9L8KR+ev10eh7
pmtiHMR3lQ1YWY865PxgaRMNPGJ7cwoVyaxIi24u0LirLH6roOSvCwWy22mW
WOfqBGpBgNZFwN2cue37oXrU/Wg/2L+7DSLE4BEynTogXQ6R3CEqjZ7Kdkc7
oBmo0iFi0srNZPP5aLhgTb9wy5UvL1oOD36pRPMaUx58+QBMgInqx2qYWRgO
0tArzmFajRfJl5lviCMBMxwPxu8g6NW9SbctbbrxW4CX9jS+z41VVGJroRZ0
iz+x8MJdBH8X98m8Qja+GuoLFL0I6/1IxT+L8ezsmxBx9VefF02mm0DvSG4r
WWnMfKi2rOtxrW9EuzPmFPgojWPde54MrsVd7+zGGr8Kc9jrrK3+2FqpfUvO
WeDyVQ7sAtV4+3wEq7e17Ww09fra+Pblk0gwriIdQgeAfJX0M+liM81Jxfyc
iMpLiHAD2NI8B+bQwU9Dnor/EpyKhQC0LknWLkBnTKz6ITSwIPjud+O8Vl+M
FBU+VYrBkVp60Ghb/Fz38qE2RL8R2Wxq3pZRigSXMAw+kh/p2qiAi/cRywJA
s/2puZafMRBbAkctUdGkZ9PNKHJkSb0MXwp4RK+1Ur83paE9Mbuq8xPDWY4b
ZqslfeSRWPL0mLVOZA3J25CYzZOs3v4QAamS5WVvHZQYpF5rdPp0fzoAU81E
sFa1FETBBojCrYcWP7wiwmY1Dy+keII/GZ6ucyqa/ERV9y++yWpGSJP2OZEQ
cXFvYtuVusew7rtZ1sx6LR4BUR3w7+sNRRKpV+V5eKIhCZTELb4DwDz3Ayl0
5oA+x4QO9wUCUq8L1Up43dDYjmNqlxQL5b9eZ0RY876MHtwXM0aUbjZOFplj
tWJm+HRPBsTx2p+g11H6YnngrRNPTMGu1LUE+e70/Mm8p9bg8fsrYP9zBCLm
RZ1xmACfRUTAxEpwvZfwjz/9+MDFubRY3JWiY3aPO35LPYPocNd/7wGMD0Cu
+8sZ8TpeqgugglhIU455Bg+EG/Ys+nFzHRkG3Iba/EpJ1pHiFlFH+iTnPfZW
5nPgt5YtN3+oRLFb6C8lTxnCecYEKg7Mg7IWr93mipyjg7LS+K/HCt1eFZQB
TJBTFvz8sHp/MGQNuJmaRuft0Y5g4VVkASP/uiZOoZr7XMFf34ksWhVSoG6i
0CKWirjLGmOiKPr8AKPfcb5HqWZU878KLcQEZCrEola7kne1CEzXlpxDthvP
j0fd26UWXqxsweSqUQHWAWBi4DzlX65zLYDUMJ4mY5H6hkoOuhmQF+J6NObO
Bb8lOCYZftaISPArQvNXOpYKABLptPlCJtkq+NVesrmbKr+6W+goW98uEPTI
XvdcIJhZhLGaTMAACBWch6zA/5dVwQY0M+/hU92nzYUDtBSLjbB3jfenSRQV
1B7h3reTHarU4vKULAF1VKR0relHDfn1sSSdN1YUZFPxXvXIxLE7EDHsg/dc
efv9R5n/dMZbMqBeW7d9Vd+ws0Ul8luJvaymBcnFyAXQfFXkJPnskeJDve+E
K3KCTL+T+1lpmlehXE4EZNek4LZkDI/yrMi0zMGzP7i0gOvgeNrqkUD7LgcY
BS1sQfuo+/kXtvacl4Bb2fJ0JHY4CTN6uEMt5R8Fla1nnYn0Ja/86a6zDR31
3XFKJHCJiCepMEMXZAcSTyW6vNZd231ghrH1gRrqlNy37guuMEAT1WHKGnaG
e+8XwP1iUPjJrldqTFvDK3qgavQMLxrAEu2KFPZztmNYu4SmU0j//dUeRTyP
CcUKPxdxQqui3Q0Q2gV27xdjGsp14SNelVP9LPdhqvUTVmJFPMWfm55tjfAu
DaYouQdBigjBbcJnKX4jNgkJ0k/pbjS+JaE1juu72QthwvKq3tUAnIHQoez2
s6xxLdUYTzj0IYws7g0NJcIXATc2Nrp1QBpdtHrvCYPbepnYB0+54VEVgD84
ZnJFW3QHKIejOJFWQs5BA5/06bnkmdMf8V35vSkTA78WlbU7sjx/vjPvHgz+
EY9Xg+DCGsMXebGrHMRb2hblW7vpjorqriBE/K0HDWX0hSX1YDowE0l+uARO
J2c1gnpipEnM8fdw728c7ciboe6PH4XVoRgME/VL224W76vWFctEmnj+w25y
OYog8lxPOIxq0AU5gW9IG44PNJh6X6yrrXoAqCD0kkYLY2iWIk7c4O4509yH
dj/wy4looh4x9lR+TtcmwBPIUt+g6lXSYAD+axEBoXTczIY25+iVPK6yo5ww
C32tQJnskcGZZj2OPEkGPkigCq3oux5jjKuzxJKdfoTnurtPw8U/soyIBdlH
54gfxWBBGEeZ8JA+ELuTKB62XvbPansnRMbbBKDgk920CF18PBPBLXj80j2g
l674e8XeUy7wMX0CFAIvbc7nByFao8k3dQ1IYk5TerpoPDDf7zZMz2iW2/3d
GVaFT2ODqkzEk9ET1m2AYRS4WLyoiDhcA0ZURJakxE3yJuGFCR/sSqC/pI9v
R4aW7KwPeb/Ci4HqrQseBLvp7rF2Sevo7sDfgDT00S6AkLSj7nhEIYV+z+Yq
+2iAuKuU+FYWYwYEiQ0g7r7oUyZY6APPU+HuZ1QwjULscPjUAzVyC7/+tLEY
K41q/gx2uTvZqlymEnuLL/cPKHmgRvBgiteNb5oBAOCUDuBh3JJYPtYspGJL
KD2AFF6ZB/jeLWlneim19uG31NKO+B+rB5VOLym9PN+rQ2CfgSB+umiY1B3B
9Waa018eLBE1Kfakr5m5riMQLdxbXYULKD+x2oYUgtlt1+43SxBzuGRd47LV
EqlRSIiJdoQ2WOkdUQBVcmJKwvsdYhHsse12zpZ2wnA9S3bl+bkad3/qkmMz
033LsN9ipuOCT0HYC3dY2bZYXIkvvWL5gpL8ZCtWhJFNXqAw3uaDUVkKq6TA
MfSuJhJM6TNSFASQWIrDaR6NgErc2XU0pFsRY0p/6u1GT6Ae83EvhN3cVtv9
0TSM2NmUSDoTa/ETCakomK5DOO5bfNWUtoLBZsKL0HR9cStpesx+JF6yPtaP
uxxex/4R9qaZs+vo16BvvxV9AU6AfCowC75r/Z5HUaRE6wYCr5+fAwxB6RXx
dDoRNu2ZW9ggeF9LrSpqZcyw7Ds+um9d3flBahOqsRUsaQmy11zOvMOcwg1o
LexeVMZxeGw6EuAiP55QBpv3PIt+hvO3lLUZBJYtP3B1/NRtuNWLfMAWfQ73
B7vYC0dpparNKI4rpWOTh2Xbs2eA4sQ7rmHNr1oW3x83ckPpLJjLreQWJ4Al
wg5RbSH/1CYUw8lW70iOaANvbZ/+axOXP2N4V8Cf4aE2w5u0mjvBH98yvob/
fJiJQLEOwOORAUu1GnN0XyxjjMyW8AhYK+CT68UlomPNeiUc+V/2jByjqetK
PinhF54aYIariLZ3Uohd3TE4yv8L/zCkxF/xOzfePat9o+aMiY5HQJxNmZlV
qhWgQ+7UN7mCjePMMLhp3h2rOJB/jUCQOlq3385NW2EgQjtWkask0QTtPuIw
Yc7KpQBm64f69x9tEx7udxGISxjZf0PJfnWHE2ylAsArUe/pWfB8EqfXWhRh
Z5Uag0uB41zJtHPz4XpQisSCorV3ndTR6OMil0L9X90KBHR6Rx/as3+Kp1Pz
yFzQSpik9huxyBNGHiRVuShCyMOD9FpmqOjUjR1/TWwviDxXADE6YoudPc65
SxUi7YoBLeXy/IVo++Mz1CRHKRjNsUGMxHlFlYFiSbDPHR9rR4ugMYVzfcmv
HeBwcbAuUhaQS2MToM+vCW0lwXE8bk9GrIrjTjNc0gD/+cpMlpnXhmHARglD
umY/eaSvp5gVO5Wg/DseqCxZUCBq2mBv21GhgmM1wJib+oKBy6OZKxNXIcTJ
nqe26uyoPUIvEeGKHQrxfKcJCihPoZjXbRIPenrzoM3bRq4K76FA0x4KU8YU
VQcstAyCqk7jtgbDo0vJJ57PhzoqZ/5ctwQDfLPHO8ttKuWysymwaMJfN3gN
MplGH1ZgFFaQmw9pcNDcPbMFcNZBqhEHIm+WV6fDMifL7GCvaBjj5W+bG4FK
160TE7UWorcx/fuJpuJaa/L2QbVNSCMXUAj6tYrIZ2GwjU5vpHy1D4mard32
u6qa5h/DzPSquGnVGFcOrzGsoqJRd+wfuH3F2Lbc5hBwa7hpYLuEQVvBe8t5
4TB51a/YyPetWjRDOq72aHi7G5+wVZ7DTos+H++GnDDNsf5t6/3J79tFUtll
hxYCIlwyaz29+ovvraXcs0rc2bWsFoWUVZ8L1V1Ym+X+xCoe0UBg6hvYTTzF
PMBIwbPGObFX4fbgIx45A1zJSbVhBPmNmbDhFgEyns3+vWiSq+8Z+r3CAM51
+OwXhHDyseEeB7xTCy5hy4mosiN+ttiPYTXh1lsJLxLc9/Mv2i6JgTP5ChL3
nwTiIKkAJs8LIaS1LC62h1+kTjM1x8mluUAXm4Qwn3KKH2QWgbKWPA5t4OD8
+VUZtln96WK7gxtiLNozYkKHrtZPP3qvPZsaqFYWKbPoOLWaR2BLdTgCpHy+
g4C9LUlPFatH1Dl4AaxRnhiIl6HR+oz9Xj9YAPUxRzrJ7VPXpiMCoDCuOScu
w4dms+TEXZn8xLnbw2jiP+HPJXiNZ6nhv1VHfEEn466oPuPRbi6czam0ETYx
cdj9FR/g8Sk8iar2N5MRPgIcD7kYo6bRBZ5mCcZOMuiVtMiY8zbloOzvUry8
sTb8Ghka/yyL+XmmFqHE9+2OgMrgRSVlDpgeIrsz+T06gIyfvPz1JpGAvMyG
FBAOPvh4ab4yuEWkoyvk2zlVvsKhELmsD5oGuxo+ElX87+IKIEHzDrJjmHxO
QpQUPVnRv5VJuQG5ESCgy88Wnbx2dKkZgOXXnIwkeMOPehMTYfJZlMxeOmTO
8y75+tFBmXlAfsZ858qLPs+dazOSIekUUkVIEv4AknLy2LR5L5SrO1gCqI85
mBsBrmvRLlVAHsWLDmYJ0gteHb0/sWsW3X02QRByay9sk0LNLHtyURU2boXe
OgKWJPLdgnKpqCRKCZ46xDv08gRdKYf1lPC9rgn6inAkiHmoR919PDusEAC/
iPY7irnqOA7TlKS0KDGxRcUnVy9lPXW3r25QQCEDF6HTYEJq4pHAjcU/y0yF
ZGlxk/AvwnuSTtJJ20iXExow9Dg+MzRaXfAPAgSjOMg8+d2LMWZiaXb0Er+f
VlxQYeIGX7mjAIDRiFIPJJBW6Ny5N8s1EhTbL/dwtwFqt9HKnwuMBuZGz7Lh
FFwmJzLcrLBPqMF8PypYdWfhD2u5p4s1a0pBGGcPMuR7Va42G8fHotoTQMzQ
e+jaRn0dEy0SkPJQVNEy9Z1YbFIgkwhs+KDW2YN4CGfyeIxNhMFng17uhUi5
z1ivBw79rIHOxdcpMwFa9hP4N3z+SYqT7xrByetWUR5sxxrBMtfQd6/or6zW
jrOmDpKqBLHwlNYoGHVY/Asl5L9u/JkgoZwmQkL0a2Xe9tEWitc2ApkqE8VE
Rp4X0Q+qBHP/FIE2qnYgrleA/Hv/CGp1DCGjLMAxYpVA/cc+S3lmY7wOHXwN
AIgc1L8Zo+HUPGy79J+alxXj1ctgQWvTDAZqVttwcTHpp5IORECJaZO88N+j
nrE/zPcGnxDIjdh2iJSjwlRpJ16A9qnm61qm472HuzPpvrEISUJqEgy7sL3k
1QCHjZFqdW5l1nEwZTrTVaZ0xUXYBy8URcmbrwzyyMIdTv/5NN1UcnzHsQpu
8Qzfy1lDJEbx101GxpYkUX9sIRwMDZbDodeUb9/pag0jV7AYhWGNTvumV+q0
2xd/GeW7vUePnyvzh2eAhirqLaAQ7Ost8GRW/x9lQcUZVqzyk4BSofqlQzLt
VOQe+wlyV3qB/GX0QG+Cf3mmM2AwZHqRZ609Fi75zzoBfQRzJzHiRmmMouSo
sqIfmafPwcm++3EpQ3pMumnrg+QrvTIyYkqua+AH4jZkYJo2AcFLg26BKvP4
QslZyVaz+CJ7izL3PEpTda9TBf93vutTBC2Lm1dPxRtdDwwsw7Rn3WVyS7C3
aRmls2h4SAXTGUb+QQdHx+oDKHnXGbpgdrcQTR+7LKedkqzRlzt/bQj4uWKq
+57mp5eEw3SAPx47rIdtNFd4qtD8rVooqACrwmlyzuezGdTjXER4Fpnl9sDN
dH8MnFeKbXybS7YsACSdftM4dS9vuO4nb4pvrnfbiuk1hXZFUx4Iq2MlE5y+
rAq8jj7pWI5+Y6Rk3bKJPOA1KsrDu9P7V9MWC6gTrl+K8c9Wv3CG22cL5CHZ
5Robgl5oyvm3ZhPgj3KV6I+pWjmrcBOf7kyJFg5treLhnj7Au2IRAzwbKIjp
pBGvS/eP6g/GTvX6Mt03zdw4tG0E4O8GCz++LzfbtnjBHLIZmODaTae15M6b
ToV8cly3Z36ucDWrfmX1kHz/cF6XDjlbVNPOYwf8nWDe+6QY8owoUJM0esTV
QgutjhltDbjdMZvECmPbJgGJjNmskT12nyeK7Kd2RW8LotSEq12pQ1DFUvCF
pKl6vhvxRVZvO+/U5FWNPrEw9TCX+YBiniynxwdPs2Hjfl5mkJTp1/6NeKRV
asAk9utOF556A/GAEm7hWvCjwJHnAAoyjmgNjrh4R1ED0dPMy+vOy6HgNg2z
t7WCf2BJxzsmSbFetxy2U+UIY1W8AArZ5dq4wFYs8zxAbcfPMoXaIg+UMAwh
6alxOkvDwwMpF0m1OEjGUSII630s/dfUz6v7dr15V5FHAB8snxSEVZIZayN/
rpAs3nRK8jOZc2jS+8oORWRgU7LB3OglJ4n+FvEm7Zzoc2rwfmpN9n/CAUQc
zFeJDXwhXyO7mV11bsYp9u6dv4Wy8V5pTQDT7AvDO/wGbiNS3aShSE7g/LE2
r1uH2OVNiLHKu/TQCvTZSp49bWiHeYJ3G0P0JCK//UYm99KCvQYJ9DDvyVO7
7j6CwqGNaWRXJ/u+KIABD1HSjWIzBaVI0x5ccKQbw7z6wap8TB3c4FYCq9Ws
RepcbuP566kq0D8hyfuz8Rm2Rd11Afi4lGO/u8Jh+lfSH+cLi/C6b+raaK2h
5IGYVkn6fuySVpLBzZi35JK7TKZFHuVZ2SKWTJ4nCDKeXODNv15p53rXk5d3
YH1kwt8BsusR3yMghiL2WinpnG3I1wrnm+SSknO2KIZ7/UWXTHDwrGKUYVU5
s+lMc+HTKTvNHnJwml+vt/5t16H0UIYRHFMubyat65m1Uu0S3V+guUHgsZeq
awu6rNgcU0YuYJ6m9L+1J5C47/AdWt4fAoLFFow8hb5XuNy/EglDOA7EMPfd
/ROZyIvMlYexmuxa0zSOF7CgNjgipj5+sb9bTRM5KyUKKOioZvqpIZ7E/9Gb
jLetNaHuGDYE0KGOdTW9s1TqpLBPs/qjlHsVhrNJACgVU2zw5PVo1PmOhjJv
hJI5j99/ofmS/zLLUQCNjfISNM4wu4gr5iBHT15vgOjcGx/jR3fz9dF/IqlL
WHMzyKr32Bx9DG2tZWCwIkrXQJtfHR5a2wqjn0YUVjxRyvBMruKOpyXLGt8+
dcHrPNYqvbGOYSxRM12/qfMUO3BIL83s6akvm+zsuoY30x9eI5GRaByNllMg
iy+CSNUgQiRL426u17k0jjz6l1CLy50/OLoESswZo9gu5+jerOImP/l1Locp
gGkAoMazgUrQr70UEeDn0kMNnXBKDfPbNxgLfPQR6/QT2n0Rx/0F6P3TQYaH
TG7ZcXJS+ca81kMOOYseEw3MJYkZNnhMkQM6m7mhNVr+Sg7kYfA/pGucKYxb
zo1zKOBVQxIk+8I6bj/moDyAyFM4WJMWmDJlQ2Her6DlnXBuHxIvm0r0EwNo
SoWA13O8vxH1F3RCMFUYjrP+FMh+fkKZJkBxmlzpb5DmVu2tLcMCpC18GCTp
bl4InPSPXOABSJEM5+Wa8rOVz3zDgciuoq9wLmbW2JyQemSJpGikprgaiRe7
o4rqz7SUOtgZ0wt9zvMvGIzvyky2b6bDP/h4u4pVykVPv9uOSgNfyGxxiQS/
ELcBMC18YtKtw/FkBlE49evXhrGKVyev8R7H8CcAnWLrfpwqEhgiqDal97DN
R7z3StpoQvwaQn/1gMNeMPfTzjzxmUD6Wit4ns4PJjofceE2ohpvsjel3pu4
M94qPwfiw8rAaTw8aYjvQK3MCFR+NArZkbVjUgNUQU5pWM7AdIYdDPQdCvY5
QwT/yCWSq9KuwuWpahv49N6KcvD9Q19ttuPlZco7zjls0Sgbpeo9kpj2G39H
XfIL00hxCCw04mjz9Du1CH7gpmbGYBKU12kqi44M8UWC0pZRe6gJp7W9ckQy
GbaPft/tWkiBm229H/BwMQdGnkKxytM48UuhUnMwRVR9dMrNdrS+Ngurg7X+
/LWVWnZlPRb8JPjZPLCoEX0TwIi5trU80rI4neGS0ZM6vC8MN0Vkj/z3APCf
5a5lxTc8CvxvfyqyumbDq1ef5d5U56WgnB3QAZ2Wu8eKbOVi3Pb99mon38c9
w+Z14MN3KSRR+TERS0OUu7kAanKDVxZFdE2/wJRUWrxWN1y04b1dAb5pzmab
St9FMCAdzBJG2cRXJXtCK6mDm3uLThFJFsO37C4AeoRFDv3H626OYE/PpkwJ
MUVwU9ke8WttXLyhT7r2xXtxnG0QAIWG7/URvTAPT0/maAE4gpZ6xRup0XPc
V8AtlZ9BEw4F+J/4rKLTsfGA+Taqnz0IscJWTwzv+9tBTMhFxLQBIyD8b6XQ
fAH8Lgxt9hr7PFVlfFDndvo2b2tSRYbelH+yIxhepwxmS54V7YwIPVjkyRBS
zyytn7cm7y/YN4xX88zETt6T2m9+mN0RcuiSAbmMAOhlWQ79a1BcZrLKAKRP
caPVIFGBqENFeqNn4cjU3uCpR0VHzjt2fbDaFm0xYz5oWjUtQIWhcSmaltfe
aNCx46izy0P7HwT3MIf8sq+zgDA0WpCKTGu6BKtKmZHI5OI37vHmfEKtuPN2
CvX6uoUmjzknlqyN0Wv6i24WlFcddIAhP6CCgV/QR49TPiFRZ+AGr42O/aK8
yDPojG/FHFGVooa6NdGSUbL+fr7WfK1jrbm3Mv4RjjdqYQuFLu7Yu+gN1HHH
Cj0OBIWjdF4vfWIqy+o+EpjIeCzX9/n0yTPyNdCRH7lpBp4g7gvsHMN/yGBB
DiiCUMvgaQDqRYqr29B+S+vsy3nmkBHaS3LY5sgnejeV4ij/OlAVl0/lw7ZX
rd6pOltyo1yfCazDBVXbYpqJZECSrR/vT+j2l5VGeCK6HZ/c5vFI7zN4b3qB
chhWKfJLc6aL5l2hQ5vI60oJQJ73rDKw/RfaQlg8Ah9YTXVDKDNYPIEGgVh2
Aq33PpUK9PphidSzpP9nTn8gkaL3r6pC7VKMAbMppSAaM1tJQMKuI/x4emxZ
TO8BXHpZm9kANqH7TLQWbk6c5FUjVKG2ga/y5HXBkU9u5ZJzIBrE3Nukzm9L
DlHAPHbZ60mxHepsMDNJZdPgtzNbBooRzy0pwFV5R5FQ/FhvyguyHKTTgEP2
0SrF4xw9D/IhKKx85BtjMF+jRgqDygApxoL9+p/O8fJ0tDjSZGeKoFFBtINg
o4smjDajcqAk1ByWFQwf0G/awz3vH2wWankR+QDGv9PjchnJGl0ms5HxdAlM
rvaIzVmwzd401pwK3cfTIGKk9f0eHfNBbQ10X6BZu3gSdS76zDkeGycLQHMy
6DvTDw/alvKrh09/3cM0Iol9UKYe0lJKTvlb5MRA2FAbHAQLz0mea0dpUYUC
PFvpcGAZVDhNVqLIPI0Hr0dCqFpesy6ZUjy5DRBMnO3dP10/zb9cVn9ot0w3
Ah2faD57sZrNTo3nqb+TgcrtJvdOmqj/k8X6lrJo02hxKJt/rzMGV5RtbSSF
okB+MK/CIyxHYw0Zcs0tLZ4H5u0AZsv2lHSZfr4971vDItzlYrpLv8y9MO0n
8JEFTYJMvojtzOuFDfNzQwl95bghCeehSmdfBSLkbwDuFGTa3NtWskgIry7z
347igMsmcHqBWOnKoaIkgUgW2xT5/VP78aZjG+tWJDN72QC8YpAR7It3vDDd
fVxLhif7UoxeuAtrlGPN0XsxoPeX89AjFkLontDjAdIVRzVYnzscpr6W3Xqh
R3LheADKuTWNXfInLHnggWxL7h4x5ZBCAj9fWa+0YaWJOJyW1RmlWz7aRMiW
OLfFqjreFNjX8029qIzyJ1xQPsi6qBoCuF1wpZWscJ61ir6jXmz5XYLhHo6s
f4pnUZBrzr/CV5TmAsYiLBr9/daZ0AlFcdRUXNyNbL1sPhaSZxkYRHQgY7bj
dgLSsjEEQtZ3EIORCqsiIQepTzFc+CpEiTQ5nD6rarrGoLREukTozSduzHLG
WG/CvaoXOXvPrCbju0Xb8awr1jJw0dDkjMq1mtMDvcBCGTLMR7JJUfa0PfC1
ikCKJKZC49kt0pTd+JkAd+tAEFuJP6GdJsAkj3sesXnmHinM0VqJ5DLRF+uZ
SdUouT+U8MbJOLlj+tAV2JVo9qayEBIxQ1MRDskzApwjyFzxue/RWblHpFeK
nDSG1Z6COD9NVyyM6X4k7ul0QEdL6rib8A8VKT4fm0CUlSa2ft8cV9dxAzB8
SWYNjNj0uNrdNUGoJ/i7C+pKlGf44MEm2/Oi5kwxgV3N/yWbTsQLhGhN4BL/
k1f6HcJ8o/46pMK1icu4t0ySOuNIC2htt47AawnLiI9RPgDjOalkFJLqFiZc
QzOAks7dlYMacIRh3tpLoqEBEs/8vYqUKRM3Yf0R7sepQ6E4MIJZnuGDu4qa
DB9OZKydDQJG6B+Wb0R9SNbjPtwrZCZx+yOLeQ6ImJfVKFJKAo7gcDJC426n
pXw5P8oYidTy6sYiNj/ZCezLhL5z/xD3iJlXMwyHsZ8XOX0beuPZYz020j0/
0YwXDc2r3Z6bpqMUILN76JboaWC11Z8e7qKo/vkAW0IhyWLZ6XxL6Z2lTYm4
lmibHIuFBqi5NNL7HRD7nZZIJGG8jgjwIgDtDkZM61JSz5BMffOd3k+VzEqa
kbCG1h/u8uhd0hqLacVJXS9O2k5Uc6aR2prOw7TMevPMUqeE1jWx4n3TbrEp
f/2rAULLoSrp/1GvXAMMHzSV1j79KWhyQONDGzHX0jgtDezrxFAvXlUG7XIw
oQ3+0Rt4Hi/D031j1CDpYj7G4K0FLtPfxboPOy2dxivc2Gr7iutvqZp7fRNn
bbrE4nl6dCG+QTHLtpIvVN5ByuEX/9u0O2AlZ3vmTOrjxBZsScQGsB2fy5Cq
GqJAo7Qj+7MKdc4dOCAMLHANepAQBoBQnKvr/xPqVYfJWLBj/+lN1jc2/pwJ
lNptyzmOiT4fl55ijPdqVtxeQ74QlslWuCJ6mNNDpelkLYgvceUikeQNnzSI
d6wrdEbm68IbFsQArZb4zBNC5Jv5Zbo9V/aQjtDqTXIPljySmX1PpdDYqhN2
5/E+JrLQ9qXPkt97KEcue/7Oid9d+cG+dpsvgGOAcM8fpTTj+YCYKaNO+ObN
rlshOR+q+QdOOI+D8j/zUjlEXiQip+HI+fi5B5Ycf629wH+8YWNRRJROHXYF
Qr2nsO6ZbnyWWP7Vx5T+P8ha6v7SPrbeDmkP00+FSo7a5L/oYv4sQ5JTxRFP
Bszoeqrk4e6LaJ1iJcxEaDbgH9BLdj0q/iXfe0pIGcjmHwOiqEK1isnI08gX
muo26TyXgf1ruEff+KpqOZRLGb2R1+ZEk/lJP29SFpJuwSOWQNgtipWLmmVR
fgPhaJAAJtQNfCPrVPNjFmuZdWfUFtyIACUYDnNvq7wbWhNvgcl/CoB5Z9+e
PQXZr98mNAm92pub0L1oJ8qMETiqZAFdTrOb1PPjSDj5zwnLhq4aF+Gu9e8n
tAl7x5VdHmby9g4ecHM8b+1S2nDuhqA9p2vnaR/45EuuenQUDftXvfgJlTOY
OWMfXT0oXnKEhAWdg+QQ660oru8rrUmLsxtoXz9okpBk6hbb8QjPiPNTonXF
mV/s2Z4Pa3+Q6mFZlpasM/OW0b9apaqgVhA6YwyrZL8Kk903Z01G7v1Hniwo
zWYJMaFxvQ40b3UwLqSb/N5cOyI++EWZGYEUAHzwIRzd/2n95NIW1x3GxIYQ
tss2IGWQHHpLwKBro2EymaHXV2/mOYsJyrUuHqYM/gwHZEZqGJnpWTs1QOfg
x7H7b9b8vrsxONdmsWlzyYZWzpNpyNKpLRmp25UsNECTPyFeueNodDOHyznN
ww4Ypls9f/eFK9qn0pdkgO1O73L0tczTRjifwpbf6fVqviBoYrUvBs/qFZ/U
IXVvhUuT/0S+R0CSyh24xVrtoqnjAxJ31kQxhPQsp0yaIBhSZgy4rNWi/ZlQ
X/xSL9EKBhOya8bQv8VqvS5xXL+bp0Obj4h8MjRLdDEAwXW2RA4yktpRSTya
4HBbXnvgctJNSJ1RuuwMIaCW1NP2chLTiM7UGt6YncLKyKYGeFZASc9V2KkQ
YXklDX9LLnFZbzaQmyW/jqjj90XDFXPyLq6YzIEACU+52d5VszVw+jvaIfzQ
sFbC2ed7XlCdfQZdzNgD3kDgF0SegHi+/tS9hlhuL/ljDZZL2xCaF7ukvhr2
x1y7u/1nn1+Sl+pTwXru/xYGPgW8MBZXAbNY3BPayuLSI7+V/9zlGSz45hg3
u1yr5ApNXvCNT9vAE3hFK/f7S1tgp6GRNGpcQXGhaINMb1IgMtJUlW/wiK9C
pU35J2E+LuQqZy21kPwxAY/pj4xzbaeyU9aX59+4QJNne2ZKPFPnEkOt/3vQ
ZFPAq2EItM4mKgC9ToKbNkjgDcL8yuBN2xfiJ5WYIg1PWoFK7lo7bAdyGHiV
0OUeJUBw+4xjbGZtCejCu72tqsA2qyY4+ILWf+MSGgoEIFw0KhYDBPrTr1Nj
V6UQbsBucXwwaoey9RzgIZHT8/R59FaZsOFyx+ktqqS1gJnnLdTfY3QNy2iM
y9FeHbggzfI4Eo0pOvaV+j9rqsgqChFNQrBjQfVa9Fpt8YCQ04Haul7CAejr
dv4J3tRU4QFBuZP/g6SJhETUDFTHdbSSJYxqJ2L3hdgbOxMF4A7LlvwyHxrn
VUmh/QrEPA4JrvAZTTXRWegn3OERIeb1lUZKwMcySdcxQnl854CZvpi5SRAu
6iNIYre+PPDPst/GO7vy6xHlmZdQHMY9dZ+smnKakjJseZbrQm6Bwz5sXiEq
CR7fal5R5FhafbQRL3pqL1w7OwjjTrIKUKPCzDbi9AGPcqruOjoWMZxtJ2vz
5DpVj2zOVRTvjNAJ9hF8audncHvRMHPGdBXTYe0tCXykxysPS+2WZqRc8C98
wGc7lmqEFCloSKeN8+bsirvfANciSeX9lYIsA68BlvFbQQeY5xm7UXctleTu
tfOmV6/v0aRUaaa17DNy5scyHLpKQcbyFAicCJJPr+0a2D5xBJ0QQIiQ1btl
8u3AQ+AFbpmH6Rqnz1ht2M+wl0Q4juSkSUTCTDRqqQl4yXioDb3lfZb70h4j
PWBk3H6blM+HtimPDpuRPzoUb4nQlg0cmG19ecFfFjINSC5dHLxmaA3bhKNW
piF0M/MwVjpre+PgpvMBZ2ktuSxXDo1Zx0Di8DDAcuJvztlJBM2t7G/oQ60Z
fCxIltgwCc/o+mQ4jJRyeVAmM0wjQUyYWCeWwUUpyNTra740DBOBKGJnJaHq
OXdXOXGb5dI+VZaCVx2J2ioZ5z9K2nS9PRcDgH/J3RRprEb7qlCWq+K/opp5
aI0qoRQbGoVmi/X/SiEqhY1BOaXclWX2MR/TSiCB60AqI7UZuoUZUzbAUyOa
A8avfnyb05fDiuboYRwyAr3meWpSCTH3aeRU5s3gIGmODA5LHlXmIxL1qIUa
S3TaMXBDgmegfY3eZL3K1zbdO6fTdSv2w9mvf3qWtgvPT5BC4wm4c8f059B1
ir+7JWzkkYeQEHm8lMcykpOFdcPVKY8nfloW5oQo8ybOLRWApOKp7Zz8pxcu
Fqrev4PfrCbFdAjNtpfiuQUrhq9lEE7fA2kXk/kI0kUAwF3AJtdLxDXktiro
pRF2q6soSdgeeoKgXNL6tnDgPGySaJxuMDWzQwkOlW5PqFfxE9G9lYvY1BSM
tOrbda5BNi32cIDbpxC3Pxfe005pnKTAXDILTHEwqoT1rvoMEb0ejy/MEKr4
kVwyXap3LDuz+zXyWDVjyey/1doeayXLL17dsTT/AiQraypy/El11KrL86Fe
OJXwOwIIRcC6P+mYV7ncQ/E6B9EzQKM4346dRbZ1JSQp2zgZsk7kN/UrD/AI
oT7+Xtx45HtKSyu28JpZDohMuXeRAm1LQ3bEmTV6iyZ7pC0fsRw5Qq1FDvZA
KtIHuFjCcu+nqPASgnWaKq5C3IGcWug44cJgyX499JQy5LYnMNQ6V7k6UrD5
wKD6aeDC90jXhqnDUx9b9bZugX0WU7Um4vdbNu15isfWmZ1qiaMccchRJ/e3
GOEnyIeCtWCSplaQn0cf1SuljfDSTOV44kwXUVnVtEci6RW92Im1uxGwmB03
Bvn6WcJgjRbhqCYoiSB233SBdBJHQFLP+Xkgh09p9uQCpzT8+pkYvvG9hMaA
UblMLPF7awgHQEh0BvMuTDbMY9YxDI3sPTK7jxp+nNkT4ao6RLyGwLdvqBZz
3Wyd+yEjiTYP9z4OshO/y7VptLzQOCdivRvhMu6dR+Tgz1+94TvJ4k6Ho6Q8
p5LHfRv9LOSLQLXfVNuvIUQviU3qxL8u380eAMxsq+WC+Z6Jk856565YFHkn
LOT7W1soE6FkP3yareg4CugFul6C0WhtCO11qbceRQ662iR1duTAQQa5qC/E
o6DgPicymODuviokYaGC/R6CB6D6ofvDMm8+SE/KH388BBeXfdtXDisOiqhE
Wx/jGtNaODgl5L26G+MG0oIPQUVj6+4jQP/G0sYeoMM3hZ7uITDH9SvPMzM2
UH7bNm1chGfCGUBUOyLH0E20HlyfiTV3fphD1kgqX+OQNyqyKAhATqYOl1ZF
UOSoOYal8c7PBG9BI1oiXsQcGrb26VN1hlgDMf/9kDsOctSL66Z3+nGI1lpk
IKPNCxtD5Bqdu1TsJOGs+RK/MDeAvoN4QPAZdHuM3cNeiUO0SZLoJ6y07z0B
V66l+amorgrEisbEf0h0zVeLBIG+AzoIdU+UBrHOkHbstCrlnv8MSnsHUEzn
JIwzpInLIm3Cj6jb5PJWLAIU7gV0cHkZ8S28RYahljf1jbvbMfhkVu6fvZOG
vy18BANss6l8JUnBXy2uEm970TIx0PCjF6IP+QhDrQuKMRkrXHByZf/yzWzp
bHUuhVO13v4yXe56Ah4Bvn7B+ihyZAPR7GlNG/S4GWyKTgHAImqQ0lTrHW1l
3f/UZBajT28QTpUyMYnlwBGgiqxagla4F9j/Ymro4WniGkI/hs9OSye/5kbH
QaFr24qzxxFhI+X93dgULI0yYf4DRTH5W1oGXUHN78nDC32y//tSfUJd9V+c
YYIN0AGHpQ294KqpPEemAnzOBj2PJlNUNbPyGnYK5/0s74dmTcXaeMZt/Yfl
ciPMaz/3YXd+65tqErFkN9+o41gx1wahEQDdJX8fWWPpIHAgRJKGnD4d2RXp
lgvnrsORazQenJ79gu8fZ978uoe1cOZ2e9lxLoLDxquEGXCTEScgmztfRfmH
dwngz1IDHxLw3ZvNDrdHvniTsCaharxYgwovdzZGOLLn/KNqaWYKw1OiTv5g
NzYfdVxggAZVSNmg0y/d+pDhMu5SD2nzwOpN488y5go/KGoshYBo00zX661k
6RtuwLqhE63oqVul56I5km/QyiIKaibIM2cjweTefcBad1JJl26ZM+QeMLrL
Glq7tZmtUNfhgnaUQGE75qEolF6tHu4VqLqhk+kG/YPnokh9iWXqAepBvu52
ThNgrlVCDj84sqYc93Jt5i6Wlbja9+gVTSuzVYwsAbv9DU3PKEeLRjxG+WlE
u9liAxhCm9Rdl1psFpYp4zzBfVkcgYcTXeTvVqIeUDgWoP4us3M4lc6Cf5Hk
CzE9+/uiwMuiVZ0BsAa+adW1WlbQwHfOTj/aN38VoVsesohXzxm7JHjpEFBG
Uagn5cVOF6+3eZEpD15M7isKRyJWUHwOYmA66JY9QMhjyoGkA9jmYvpBQ5tt
WGcCQZVRTezDeLiazTrN597y714sZxrs06kGbru1VDbRpYW/VrjFWQcpcwGG
IPzuomVlZ4ugrSsDc8Ag1rCpKFLv07RVEeV1Ayygh1Vuu9YCIfuIVKeV3oUE
mV9Dd/oZwYfFgi9Z2SvF6rG2h97f4GHUmCHae4HDnmhsFcyQjE+KuYgp+weR
r+p3OZY5y5MjLrpCeDt3Ua8aFhDKwj1bJpPUDjWB83uwMXdY56fXaLpBH5av
QrJ+Mfb8ppPUc8aXTYxmyVa9ADGFNTHAcJNNKZQ+YPfvW7xFfA95w5cs4PXK
g8uMzKdwjJDxfuhrwNO5zTdBDE23OJXocFSzgGzfycMZIqjjhe/tjGblKCTR
fB0uE2jouCFeCYC+OgkXzaAEPN5suvlkxzXlZbjsP0lSR/WPbVkriIopkRul
UMrnQEf/3bT5Di/VEwrcEMTGn3fBPb5kEJ6fpePM3h6SJKgQAcriLSJdQozd
OH09VRGZTRdfvVMxgqXOU6IfcBx6LqQ1APqGB4PClAB8FhiHRmyFX52m8yrk
ukt9tjhzP0oJWmHNI4SgSawBXxGGemd1zGv3JvEJEtCPNcTOVTNhRXyEakI5
dBhXrn7C4SDz5m85MNXu/3x7ha0OpZM8qfctv/ETVQWx89jA2uJwQ7m3ZMiB
2fCSGX3IpUTHfyhaOQpOtz2vt9d08WxGNkT40URpRtaD12++FNjyYR0EBmh5
7nrTDUzC4iva76GFCiLxF+r6Xx3dCP/4UlulRxJXBzbUOO2cZwAfA+ityzVn
v3KPsC0NNPzO6VFVK8mXdxKO4VVpSOnc+8WxV1FnqbHIa+UCIK2Pd3UXmYYx
N8byFP9rGT5xafz6X2FLEyfUvaT8iWbHYC8fU+Bv++WpOeJFpzS4K5gKxsgh
hNqjyeDdQpJwdHwJXReIkPlV9B2qmkA9gMaFPdXCFI2m4oUQwzuqZFZN+LYg
yKUWLdK3xkq6brUm6wDsjoa3lI60HFODCdsBzatmI/GiceL7ngWxhe2O/HoG
ABKz+GFxCOiG+es2wjtNb5wF40SlB2nyMH3tslFxhJlp6jjFUKFCLN1oCKeR
HBgYWyH4pOeiuCaBtUcYCl/luhNhZeyhoRTP4Ili+LoKhWugZnBzBkM06pAe
8h7xPHLPMgKX1Ca3fV4u8mSTowKhXpJtAvXfyyGbrETK04X1wrQhj8mVTNrj
7RH6ZFrixHWkKKpyCSG97CZAZXCkp0iefih+Nd6rXDgkHh2eOF2gj3MIQZch
Y7OAxtVm+oR2VnbNpbF9WvrWMZaeUdYbmWpcE9S6ud01UKRgiwZTHSGiBL8Q
9fk3TOQee1E8JDaYg0XnAW/PszKsGXWUNwStF52UiAawcSp9zbFQWfeidcHA
sEKQWgp6NA1QfE4YSa1QRzHf5GuJGf6SBqVHUbFjVQ88ndGne+zi8uuLCjQ3
dL0N+hClbxZ3JNpzWfpxEOAeHk567LkKLMXHKgy6rX7SpsYiKAwAvHpuWWLS
OgBTZ+1/kPtGV5M+dcMquVvyszKKKpTy0FPcD5jAZQLzjkWZUNyg2AP03Lmh
57vYVJ5JRyy/CuVWDdDUFoEL9tWuVcPjWdrwFmguQTJyU8DrBnhuksojdRET
PBQKJ6T2ftTQTRTwW33YTpQ630tTBQAQ8bgVzA0IOXpvKkQauS10AhZfkmP5
kZVY2OMweXSmWo0qsBnldYjMcQ2Lg2lx40pStH+GptqB49WSJBHGSbKqUhk0
2A29uKIkgSzr42YrcQl52amXFnkVUcVwQ/wdeiTA8veEO2kJCleUuoiLddpg
U5K5LTGscNKxDP4yfSld9LHzn9gX2RXjBkbd/7hebTqrsWsfqVKbDlz/5Jg1
vHuq9qP2UX8LtRvOPpvN+wkKIN5z5wRLiyEqFE306JuqZXHwpZUqmRE/ebh9
kgkQyYQji2FVBCCp6mpifsLwLuS66CyyndxYhzAvumkeRjI1r3+Wm1VEE593
EYv6wk4+XPcrJBnqwS7cSAerAtd16ljwZk8t3i6bc4vztVL2mmZhBxdxstNq
teiQbLM5K9GY2JwtAzYkea02UtQ7V0SAx6H7yo3+OogbGShnzf65DNRcMGrE
A5SeVpYV5nJCWTWouZRbuc6/Vkizy5BIdPoLT6Yh+/DP+MxpWwwPVhJf/dIg
qJZP1YiImgaKVlaKU3Ad2FMtnwWJbIRYhw8wf+PfGrpoh+Pg6EDrF4x/hynX
irPM9objlZ52N5wIi7AD5FkVvwINz28Uznpnn01A2Uce0I7ZZWmQbeZZNZcQ
53F73yguY0WtlqiqG/uZDBckVoJYc3y1EazTBSi/gEywxX81CrJB59eLfTQY
MacZESQcIZ/ZSfuwELScFiQhD9aKd9Cpso2A6Lcffcn1i/VB5QWKIa/cL7XJ
vI5MndnzyiWy+OtTzKPkmSYzoOfRYM25Mb0NqrZpcSFotmGprEJKGcOUr9JR
VY4p77OI8Bo03jXIAT5cWOSa1E7Wd364DzLWNwrS0Rzz5FrdpuRM45IbFhKx
Vab9nriXiVtawBJJS+SQrDno+Qg4Zx2VX7VKjEQCyhNTGVkzM+ILJfYJfEQP
24F8isW50LrBOa4DCr+jZE8x57J50J8WP+CYobPJCqDbgEQ6EFS1dbG6QXWm
Dp8FR2qpH7SbAdi3CcJVSiz6MUYaVr0tbrAWHFv7N9LYd4hvih9qqg7HuCmZ
8NBHczAbuZrwQq5rqtVp2ex1RiOPXQRr+mRxdJhuiNgkMRlpe7b6ipix1rZk
FSDG9G5JltuWHAj9KCu9qN9WdE5Dcf8mjYS/3unmuwSSHKX4BS9oWp+xcJtl
ZMa6V49Uclv1n9DKbbhcWXVBJfYMudtsYlfIJpeZ8SHOJ0joKlw9YWHFJRlC
8owHEQhSaf29RHeDERtpjvtF2is2xYaQ5PhGWLQ3Qo2/B+tq2Rjy/mMvq3DB
JYu60JSpmNHiBHg6VSlNiW3nKnVncHGF3bFDDKE2v+ME2aHJfs0XJ1kUFSR0
pwFYRQoB9hGRmBIG9dh0E/qOO0O4EmsbhxUHpiGwIwrww4Ks3+a2aVQRlqfZ
hkQimVeMmYwORc92FvXFHWWbwBDSkdWU4uUU3QMfJ0Pov4JEaXrv6sHzgQ5h
IkoFOcyYljpJQBnZfswrymPrzZeb7vReFWpsydpyUlV+6OnaX1Aa93JeRTkb
3rgKbxdsXO+vAUOdype3WKeAr7/k08ZRJzwYjFe/+aT4GX3Cl2xxgkWZt3bj
L3nQbCNEVS/RyPrWgYtWCllO5A5uhJsRiwiUWcC9w8EwovZSwSSanYtKn2b1
uDzXNu7t71leKo3fWSkFieZKpsF4Xg91sqEk8S6t5g7Xj4qMMAWKb5vuvNsE
nJN5lyWYz8k0QBwgZDgV5d7Wk9/ZhGiRKS9647/RoCW976G7nTftis+jasQq
J6vJNyIDT2EL9yjt0e6R9/+Uxout3dKHPxR/dynXhJeQzeK9MulcPJVfQHOA
fLT8ShFMzpdnfN0Zsv3lJcCPNrYz+IC9IqmmOU3Gj1jLbSMoN5Qjyy7nz3zM
OUgEEYI6wlLHwUXeJpZZrfWrK0so0gjiKwfItUYXCBuhCRpSKqXyLKTtsilw
VDYS03Jg4+1anWKfKqgoU1oD02ALI6jC19y5vEILZDC0qbXE/GsSym7vvtSq
yiWMmU2gDl2bA8L4nuOCy9oycE+EH7G3SE5nby8UqD6gK8z0B2Qpp1iEQMrY
6yCOzd1NVC+X3f5XN+UhhcTMae/3qFy3CfeGkxGmY3o9DII3UF7u4BJYgYEa
SSM7tEoH881baDN/dO9OP+efcPS+OKBhKqSPY7RjYqLAiOIiXE78Za+tGG3R
TX4erhTdUNp5DAY6KuueEBgfqmpWBgU9+2n+IljigGN/fJNmwFD4mlCwv4YW
NerMyfaqQNUvR5HYn42yXE2Mi0LIQIIQz6lr3Xf5mwslsQ3jod1cP9E1zQv4
ylCqQdKkWsHXFt2P0DMYz3C0GgB26fwCTr8NSnUjCk6SFd+TVenJm/+xmr8O
VX/RWFfRnF7bgrkw+nKcc6J5fpo0/CsFhX4q/ap5g7pkOxWT0U4KPIki3d/f
n1vtPh5vhBhvE8WOZEr+FIbBsxZM8QmhJ+W4hFGH0RoTy2TGb/2pSyPL8ng7
1S788gWIcK53HmTtC3v/Zw2jff1KUQzlzDxwzuGEBVBGPBiZ5bUqteNqrsIn
lpVc1+PT5/Ry6x3L/G5loqc43h16CgZiAz0RznqwmAVCGSMSPcbq/WOX2RmW
aL7FRoJ0iZyzoTz08rJyl9554GA4LX/8HXsXbL8SrHzd3wcIhKaIlgfUjH7Q
ZaqIToSofHS1s5Uu8/fMhbrRVeNNswTXvDsd7SJBaU00tazv21DxykPqFMHn
p7Se9q0iXTMolXOb/ROPCXg0ddwIDQlKWVXplc0IasYNVkJIX9b4ivNOVzSU
VwUugoic8C9S/5GPIpyagthqiH5MLLHEoGQNhkty/3UsixPRnvzFKroXB+Lf
IX9+evnkAz9tuugtkIZE7QQ/viFGyZlZliexVxUZBTZpy4PnrkxCATVErxFI
rJjxDVxRNlvSpbRAqw2QirWSEyRbl4my70pqq7XGQqMBbRPmO7NgOUuxqohC
uC/kaynmQ28dcTB3tqODeyPB0xsB0tdovyTA+rxkvsQao0Nt+kVvCZbnbWx4
8k5GFVdE8SC+9ZhqVuF3C64xOfUv+x2HPh8u8yRpMmF842sAnI4qdou+5Nrr
5rbTmcFE5BNo1F93OrT93FJok7JebAV7Bp2b6WP6sPLJUZ29bveGdoteyFJz
+z16s7hco4pgeH/AC97RMQ+gENSRNTaokbLxH7KVD5NmS4ScPJjHWe5/0j/7
ciETz1ddIyNQ1gtGXrgJAINte/mFRvlr4At42YmNwK69wwpCdGQ3rmY6ebs3
SjhtHaJfQxuOK450gP7EGAnwHipGNXyc1NK6pSXCKZZkjJikB/aw21YuyFR8
yDqCAZh3NoOW5GzNCR8y/7cl2T1QpWhjSTb5419M7dm1zFFkBjsDx0NqeYTb
0TcmpbzZp8WpmAzhpDvehv8eRGJ1+9YlacJMVc+Thpzxrxwnwsx3kGxPf9F/
I6uJTYxCFba7DYxZPcUTf6BKKFBH7rPZsCVGUEnNCiU24/xTXXq852G0tMfz
oLV7tlVXD/IDxT7qGselFp8DvDV3UZBqBW/SuKD3hmnn6HFjjJdUeixIevH8
8mPM1zxDxOFbNECsiqpJCbQHaqgf8+HDRQD/5dMv9NiwooVnDehahnNKZxJz
zq8fje3+5Sm7q2EPzCVEgQxVY4myQ6RxoH0YTvNClRJKuuiPIKv6hEsDvTwD
Pq2W4HHddfTaHeQMbUJKJkIbOo7Opg8etL7aAz8VdRgHe9Lfo4xVp0O3keDx
/HlKU0sSL+jutt6ImTtojYuJxCwu7cg1aK6qXqhXS5qdxNHoSnyaX0GBbpXj
965aG/1bgpLBMDojR+eM7y+NnDaUelH33tvqmtA+bHzvGf7r9Br9DrhTh6HH
QllxFAgILMUNzn3lYFkFaEi/un3z97/h1F8ymY2fVuuliFvM7r2x4drMovRK
lTWRbuQIlHax19R0HSA92pCtH4Q8USBgZ5Clai4Val7lz3TqNuc3+lNFMbLe
iyAgGjvjjcgrto41yWloSJGt26Kth2z2E4bIAvq2XfaXH1BgUY7YW4WwebBQ
BCGygperk456BzsSNglzCH8oMwGJszuk00ouGb3XINZRnwAVNFOMyHpcm7RQ
M1mvse/59zOEvHVz0jP4xE0q8qxVDobrz8PBIipFnV2UlvHHC2Ere1K9+pVi
vJkT3xhMZPky3eJApXd0GdMvhV2K49cuWvMeLP+VWwqJmC/seAFU+u1VTog3
yiG3rSwWd304Qi8cxJvH+1oNcNBXJ4bchm5cSgH0zHUnbZulC2YzqVnmlkYe
5/3msrrNKie+QrjJpXoeZu7eoaNndlFNVGjJ1VqahevheC/In64V+dzc0OT1
vu76nyTQlYfEQezD79U6JvT+WDrXVvNj6lOEXy+HtUicRmql6l7nSfupeJ2P
v6zdh6k0RY2WocJzNRCxcP+rW0srw+HpcfHUBUHe7TJz3QI8RIxk6kuDT7e2
CNA1VZdqfGEc7FQKWFaR4B6LUBInXca7P5HSk1wo/UBpPTl/5sSXYW5R3Sr2
4YEJgw4xRHjs2bgFlxbp/nqa0Cs3fGAxLfqWULojoz9J8cJOdeswNjfuYJCb
3oj1o0JRNj3A6M9gtlw9FJ19Y9QivpslY2vJRQ8+BZxstJVtzI5mWsU5IYLe
6HIYXvW7yGNQPd9Loic0MhMnlPHu0Vcvac+bF3mVmcHRWnlryo1PQyxXM8Tt
lwGNIfsXt03CeX4VMQ83n9XxNGsPoaVutLkryvSU2w8ijol/OuTfkAZIYFrz
s66POt/wj8aH3z7C+tQA2EvRtXMKDf3k0GxuIoZmK/gqpdgPzKi1O0+hw52d
cAmNQRWQkP63P6nAsx09i8EPOgoadmFVaMobX87M/5gSZcVlVPqq3wMu7IOS
6nEk9iXgedsxCyrDN4cXt4rNdxtbZc3K69fAvQBy0foVBLQx+x6+m7EVM+GN
86rRN7Ohsqn8KJkzR0lkKXjb2IBxZ+qSc93uhW66EIqH08dB1eqd2vH8ghyM
CNmRncKaDZ1H1LI78hWPcxquPGxXfvAM1YrCBJEFrakpzOzt8hpQGQYQub15
jFkgeZPwx+TmWwf8L8GInrPuFMwJn95ILZi+cw/prIH7Ii4CAAKCKQ6iJHJo
/qTR75EvooTNI0vxdhbKtROUYL5wfSOCo+zectcq7T8+TBwCM9YVpKGmn57p
1lU+4p0JVAh824aWesQuBo4af4wW6JEAs2uHVRU2O8L8Huy9otXyZAanuO1V
0hrayUqr8YtkpdCJkApgT6E4dDosn5A0R4nnzY6NoGALaI8Cbb4Va/pudrIK
LlKJUk+FeUXd5XnyUmU+lNyIjNb5oorJ1WOd9D4dhlbYD4YQ8pM9bp68+NN9
m1MY3Yl+LtWNpTw6eHn4NrrEu/s+nEOpMQq0oUapvvSs1RQ76rM7b8NDf9Lz
ohOEKIbvDoaBqpXvgldPlcEoEoZIwdKnX8hp8s2rH+tiJLbWjXfso9uEMMer
Oqb8x7YTwmcwmHKSczn3SEJTK1XBsPDQyGvUqTjIbqXpI6S5cfydsvc2fDry
Sf7vtkn75iib4gDwFGibEOrKc/mNWqPMC7bkpW0AwCrBgsH4h1yzYeSUxDxZ
74/ZBPVJQxBtiO40mtNByH8WlKwLIn6cDtoYMqGiOtrLrFHu1HZYVAz0BIiy
HT3dfN8CCfLcCPEHAmYCGv0cb+ZFG3RrusU5glS/5eVx0e1e0ruApNJXd9FD
Ia9cOT5bJ5pTc6r2sOJHACzUBIvZpfiLjRCasCdMzo/940xgN+dfyRLAS5BJ
4Pd3Q0601jeKUHidalVF42pEIbR9YqMzMFETCcItvHOwU2Dx21RxQ7815q+a
ab290a3WMd7UY1EKfWdCLiSUTfGwRHR8mKiEhS7V1vna+xr7i5SeLrH8QRwY
Dv3dlgWw9nnOsALwnnJt72cUVcBtncyLeuzHCu1oW1273IBtqtam+Zw9DPVa
HdE3P5cSpXbW27Q/kFdrReea02PM6YBltN9cAIk+e7po9aJ4qeGmLVyYmV+2
IP0uaFqQbkXULZFnfNyvof8T+umpyR5iYWJzY+KJRsHQbpow8fyjTiWYJiBw
T5pLVNy0I2UcdXNGUK6WGZVGEPGGinOd4n6OygjjYrH3rOz43cJOinhZaNSk
LMvlMe4EXFsD/jnGcBcSiXiNUhr7f7uhurAAepKHAqf2k/1S3b0GfiDevtFC
CyIcjMd6w8sd98dOgqd4RHTZjnR8mZbtkoOTGR1SuaykL4d6+sdBjgFTCeSz
m9icLCavtWnVo0mEAsVWZn+OIBooL9lr7ZUczPwG5JYAc6wHggGKEoB+AUnm
jibfM3FX9K1xTWcL38UWZ4BNKhPOZhgsbJI2HMNUuk2vVPWNW7XXpGeJhEEq
OTfYv3q5ZQgUVBqmfRr4qPUH1jqbBcEAqtmtMbAV//lETGTK5IaXn0JNVGQ1
lf3GKbMORbqoQUUU18T1GOGJkL/9P4D9gnmHIyJpohimYUwjffublJs1TSCH
Mw+pRToJqf4Rj9LGQLPnGjyq0gbw/juOGbQxYBKW+ZTL1WMKOgt4zZL+xT33
vp+pYQFGyjYah5zIbrj/XsU3ioLAONGV/J+9rV7L15JmBrvLmeknisheQODP
I8sCKc/KPV0gd3UGPFV0mM1XiJqj9ey81/46VhtQJhSfGoYn++OQBXXRvLK9
zdbKSAP9r3Azf1J58Beh6nk6PCi+2OboDght8MpbOZYA7c6Stz7KSpzUg5Lx
+sajZmVaagyuJJyNxm+S7Ryr63fN41aAIFVhvzrEDJSQm0AK1pH7g9IlRKB7
mudsZP2LSN3g0b48064tzA8OEPt4ez0GJ7zjzI2Hec1N0/Pgj/tYqhC+5imL
zMA/MiIs3Jpddl6t6JXduLph3xHVsHEEt/+hLNLng/iHNlRC0Lgjtd6+ved3
IQfFKazOmiTU3TzsvEWYU90LfJ+ztBNfJqnRoKOgLR6kiJt8DUD/1h3peEDa
E5b58qy/S2P4XX9cl/OvsvCCEe8eT4dBosDtATyLnRk2gbKio5QiE+Zx6BqB
ev5ScAHujFBgOiwXRLwaBBZ6Zu+XQW0hzOc45S1fn7CCCf5ygHka66klxHsU
pbvEUCFQwVKzvmTbS0gh6u2/B0FZRdHF3GjUDP2ZQfMGUGYts7ex1xPsICUO
rjRjYm+Qge2ukxxq+xYFznzSDAiLaHUx3yMhCBVeYy+diSCh9cIDMN1AIiDG
Xv4GsYkeQCMUL9HfOr46uBvdFxjyLDsqsa7qFk3J/CbF8Bz95uWazg0ifUAP
DwDH5B9ByqfTPAHnr7IdUT5LFUZjIeSMnDIAdzvi2/3kEW/r6ar3eOYB2XmR
VK0MYdA0wMtbG+Paf2KbHXEnI9dh0fKBFvB4kc2pa5gLx/YEkSk1wh79iqUn
00vFckpT2FSVUZt+gX5bItJE1BiY4aiXM7EiWWVva2VWaXXAGp+AoxWjezku
dXXp5fhs1QfQKpfGxGNjHkv25fK3n+v0QPQqKlA/m5vfnpBJG+RTXT8Mglv1
tNVEorSGYRe/PfRlFjmc9c9IfAhhI/rLkkgRq+2RZFC0r3y9w5BqoStIcbaZ
+LoDL0pRmKjcvQ4uDGASOMI0Yvi4x116wrIfthcbw3lCpZiED8Sztnr6Kk3R
k0ANyUHmGO3oGSOktPCQHOY7siTzPk9rdNVIXsljc6zDtPkerollsVCVxsej
whxgAqMBauln4h8IZbVY3fC8cB514SNiJ6jL+cO7tGunMqA2cHIUi4Kbyh/5
TLP8HhhEr4qwW+HjBHhtk+WeAbHBQN5mXnSW8bHl2YEBMvhW5a/65XyMF4Lm
2Qk3EVFg5v6Q/6SDWdbSF6FtsGDvz4emcwXAFZKivKjGgrsoxFgWJtIc630l
xqC3N7JASCuLsDvkPvy7bDxG4ec4REjRnO/WSSo0VXtCMuRSYV0eYG86nNU/
BJt2B+gEZdeH+72CjDqh6LgsfaTTFw5y6dJlM9OJ2GghkiCzHIrPvGPjgvwH
zghyOSwtsD3pDauk/5KRaxjQVkSzm2jfVi1X4bqV4r43jMZ7eBXfTN8EoXCv
gN84EV7JFmaNYNPh7YCIH1e20L+tQIrahjDIVq7QysYWoPovxTQ+TQ2gGhkY
OZn36YLIiRjdR0D+nptiVOtKOMl72OQwEf2Z6+kSSGppnrzF62Rk/4Byyo4V
CT53xjbFa/9fRpNoHJOFB4yCo07nBhHNXOxg+UODtEmnvGPLaOxH6GK9Xp9s
qbkXAV/tvvKfixzWlOsmXrkm6Q+jW4Nw4YDMP0AfO9oZvb8QgVTqajnMZKz8
gHS/EbAi7VkUAou0nmvnbv5qEYCm+JpimOP1IiNdXhiAjTnF3Cv2Op9YhtSJ
A1zB90tzFYnGMYs7DqkSb2ZuIq2DKRr/VpUZoR6/9QUwtw6HVAiNa14XWae9
qHWilkOKBhdDLuPlCFGZEziGs+xpUdxysXKoTj9ixoEm81WPxVjWQWx9r8MR
pdHkSgxUN9SVC3RzyC+EJ8urWXOZsmRcrMnLY6+IBM3r+N0tnNDTNviOaRVb
AnHBzxDTZSZ7CZMA57k1NgR9GzveyQw1cJ2Wwnh/VPQMKVc9SKaNQvytJOnu
xSBRUwIib11PLG2fGEbfGEvQjPgWZELImtMSVwSVv4VHWqQIt/6EItPepVTt
bvrY20wNlzMwltCluc3CTGPQQ1YF+BpYFGM3/2kq7gK7qRMXpQVYvLZ5zF8h
RpjKdOQYH0WrMnc4NsZ+eXvg5XmgBwI1cLe38o3Kf0hWUG4nkuQwQaG13f2s
Xt+c4KZlJSjtlYc2v+hxQdaJ0SF1oeTBJP40RUIexwPq7+cWrQOADIUDLlL4
0WTwKhQCkq+1c17yMnqHd70JIK1TvYmiOlU1mSBOUD1YJ7WEj3p5P02YXOvm
JzaFcklyuY4uLNHnzZw40DATpq1dcsfvK9WBlTCqk4N/srUGcJgQQ+8tR3YV
RihEAHkJ/jRUCjFCz2TaK0XOBAnWpQO29Sz3xy5riiFnNt2V7fVtAjP5ZbKw
OCngbkOoMso97SilXAxWvV7A/+7lMM8efyl7InoflXgPyzbPJw8o3GBgBFC9
6+vceh0I+vut/WOeraYl0xTEo0iENbm+2W3gaVNU7IqHKJBbJQqK6JQeW45M
IjbxY6rI0Ww01/O9tyZF97PXcUWuMGfzgZoeNuaLPa2mY7OA7iWVb+zbO3f4
EPTAGkuMrmJ93jA/7iNySgKcEMJOH3xiOVA2VsFueCnW07klZ38RzADgXRgx
HBLksa3RvfL1SQfy6YUrqdWHDm3LEari9TAYJIq5IBdfkoNqgogw7XgZzaCn
2qYwhYpTwpjOHmAlDG28RjiAyTTg5pQUa8duopUdoMUe17L8Ke97QVQTd3ff
vnqxrxo+wp1q3yr0LpalKICUBuOAcJjH4UxPW0WpM03DBeMmIHvGeUP1+iTt
+dhgY6SEndT52ek2ZGR/xfPfOnCTSuzPpsjbiIN1NkqJtz25yBex5czoWIef
dgCTnCnfrjAkVXN27SArsDBQ7bWG9KycThBLPEoIY66WlIG8Vc0GfSGdqPOz
5mRz3sGampksW3R42t6MTbmBq7l9elwjp242dolBlwTIGoeHwqZHbuxJJxic
8RZ9cWCenV4KE+inWM+pW49+4L3EJKRd2IpLJkvsJ43Msjt9ZFmRQsQmgZ/m
mOzAff5cg2oaqOs2U3MKNm5IgxDPHod6aeqX6Bfjf3E9WefoTbDsIjinB7qg
jHILv3P0omRfkng8fOKi9/LykZetqod6juemPPtGeDBy4jIKAXd23QjyT6GN
1uqRh19IxoV1g5PSZBaSxDLJ4fExDf7t0WudK5m31aWacDNmFkWo/AiXxPiX
zk1cKz7nD1mDnky8J8TpaYf+LfU+5mCc2DXXj/G3Fd1HW0gqO9Q+XjbPPHxk
jz58jxBAYVH+QbeA7TgzeMiNnzEeUHus2MwtexijDPdcmQzFKL7EYsRciWZq
9olBR6/y9HWU7x4DEB6dDfg36v/PVXsciOPo8xY16PjPF31KKk//gc63GqvD
lfIq0hFa67C+6uhqZPnO69h96MGTnUYfzzkzOOk92KUsb8L70ZAN5ppEKhck
v8oJZgPToiStHPme8t7p2z+HJhqpeRt5JrMMTFWExLOhfXNonfeg1//2paQS
8RqDHlezjy9YPlWrPFviRyHuL49UexNhw+ZYLw6nxxUqLq+a28FSTGnxiyYb
kv2AkzmM5U2lRtK6pRtrjC+YGNyJ4//gTMOOFCqyBtnzIBqyA2PoDEC1vc0F
ZlNsTXasCLKdIWjXatXI2/EgYvANQCHGd4BtXGpzL69xffyU2gStDiXTWhcO
lcPhc3sBtck59F7zSiccbzAymy+ZrZtG7RH5A0Jbpo2sESsnI1R0QkTWP5ff
o4zq2VNuPjMW9D6XXlntvT9gXWssmdeR1fSn5Kk6LWpR3Yns4A2xKzHAUhoi
DX86nBoAshvUVJ0NyuUnDaiYFoel8gXFRmnNHQt7ni6flL9Oh/frx7DsUTjU
coifLrj1rLrmf/dS11FNmtgHQ3XRN/NBH4qLodr8sWwp1T5mZNRLwKZerVaB
C8CL8m/Fd+VU6fsA4lzzIB81V805jr1nQV+wl4qZUSs9nxwS+uXRSeaMxBM7
jHCfeuo2s2qE1S6tBHcY+sEox37JbMYgeAFV4R4jBCwek/i0y5q2HcIHBQ8j
4TFCi5/EUiSfmswcSZMtSLGc2qjf5g+v8hiasi12+GxZysQ3vtQcTMU+ZKAX
P76A4PHkpjjrV1WjA0ag8OY3DwyUVKgsU+QCPwfT1SrCZUPI9ZgiXlAEg+93
4Swg+sm/M/siV1r9DSGxdU07iRwRlPr06joZ1xaUffo+txzbLNrDTzOI/0oV
Lb6EGON7XyUtA1lGGmd6RqwtC1MKTKxLBFRpQhIPYJYgUNfOedwcwNzO6jqc
GhRfbE6akG4jU3J3bq9N2N9reQB/84EMzq+ZG5efYwP2WAU3Sa4nl3ck5PsD
48QarzQdI55y1kTH6NGRvEHUkhqyWf8j40sZhhvPTVlSFYYafWNy7PuDU2ZB
oLdQ0M8kd3PB75dA9Bj/5sYp4neTAO9TECAVgej8tXwppplEHXO3SMI7rj3U
BNoe6Pu7/PxxUx+9LBV53ep+6/Rzu3lFPdS9Uvf+oKulOPCmwfu9TbPXbOD9
uju1kMez5Y4XEGH46X+8/EYUX87De84jZ+ULNtb1lApyOqr8JJRB4J91UzDZ
apw5Kxoxz58sipzqssWjbrLDMgFSzxwx5GEcLNWWm1Wf1UD0RYReDs2prC59
Gcs9P3/mebCKbh3Q0N4axGwg0Hx4XHR/BFOUmIYB34RWdpc+oRLUpLDQt8oi
3nFOZxH9aSQRKpXGCkf79jMEmxRnmcoXcDj0MuxSoZefwkXUpVz64vYNBEKY
cSmqwPAGRehAYwTTVLqhl/BlzDpN7zqx26Z0EkxykhShYM+9H4bVARAEC5ww
KAEvAFENzVaYBd47Ej2arn14nr6Jydc6s4vvqABhxVHDWAUxZepkKZIZaNo7
Kd9wBLvUqsU+yHjWGX8ddP1REDBoFfsBJv8gtaIC5ugRjNChunt47zUNE+lK
UrLPkpH6ovWSljb6bcZpA3n7+Y0/wBwN2TmE/Uq/+fjUB2Knus7CqiK7DnlC
srH5C/Yq4e+k5Awo+sxCaifyVg193NMsow6WZKOfuseTAE0M2sCSS3f/kQPM
VB+zWBmR5UYWSV1NEAKXrS3yZtjta3LpJjlrdbs/53MVr3aWvEqCPDz0sYAg
k6KfbPpZyNPhxHFo8g4XwcTGFh6tlOGorVoVhHKmg6vL4aodUhFcQzL91Iph
aiaqH8QjlP0SVSlqdEKBB9RcI1TZ7UDbSjLxfJ/bArMqHfrve63V9MtRV+z3
Gez2DqmMOUjHADaFBsz6I2do2XCVFTNuStD7fZNBVTV7TbM73Gbbv9iyiZUY
W64QKfpJIfoDYswU1jVoCbq2fc1kmql3B1XREGeiX/PgbI/v4bJqjusn+NO3
EpIIVfheC/QGp4vIQoKpPvF04q+bDGcIUMySDsLt8ALAocgLMHq5YBZZAjgy
4aS+DxN8tjCaN1sGMj9qpbzS7KED2swjPYyg2bf0ZjtNsZEnJgrW7UnjEjpk
HO57HQCkQX32xllLEvWVShbEv9ZNMCg3XTLzkFKAv8+Lugc6z47peFZjeAht
eIy2iVphMnBXUvj3zyBkwqOhiaqV7EQIdP2SCpSZMxKwOy0VvSyAoISQERIL
/KLiAIcjVyp+wmbioDeB9Y3WJoDeV3zcK0bf2wEzkQskBxN3J5yZHNqyYKfT
MnnSPa6Wchc2Z4h4erlc+TqgeIG9PHJAhLvkQBybRwwl1YhQexBUnwpnmD68
1ONgLJrrTmoxL9AcoZ6m7V9HOxRoSaBDKLESlJMuihIHKKU26cD3dFQ6eb+z
Ft4mdfyaVEj51aDhMfTDle9vS5LJ3rkv8L1VtoERmWGex2DTBZoKtMyhirXy
9m2ciJ+30Bl5/QZCvOI0Lb4wKhw32OxC5nMnxIRuLvPSZqnWZFiyJqzC7WCP
YU0/AfsqWia+a7KFbYIYbQ90Wx4e7wUloVfzMWveP9Iy0zDcs8DCyXCwWwm5
YdFh004VgIXXasexBQ5CAOso9G7FcLC+qoWyEY+/QxCLKz73ZbDfbQUZDBG+
2oW+v8Du6qpFIQ4PkCb18hWX/F5Xhf4xbRFZFdViltmuFv6cGHZVLvTHrFaM
4NDnBJqcG146hHHoUmCbq9cR0sP24KbvFq0ST5DOIYXwlNDQ2iyNNavCduxc
CJ+9CtSv7Fm9zkKgYwbdjkEuz0FMjFzo3U/GLzseXiWu5wfOS5DD0qwHMzCf
EBVdqwHnvYWlq5zbTxjYnOtd9VwroTxIAFc4U67DGimrgHIEjYcPpl2F/ZNN
HnAaJyrNYtVOjzilGRohGxJKWgA2zCycejlrER50lH8ZGJ+A5aNXEeMvx6rL
ynQJZ2lDWKe5MUejtOJGNOyDzRZp3UEzi9llKmRdPg8m3qT0uOwt+wVF8zT/
4gKACffHM0hIpCmneto/VzVhwNcI9Efi4iUeWHVTyl5Z2G4kQqo0wNVSHtr7
nvOUx2JJqS7HqbPp6DS9EqCGui7sHt2p6VTRUOcsjZCzd6hbjNHFbjLLTwlv
o1e7+fOF8Dk3QWc0LT2ibqboFSmCuM5V+nVfiNNCRxzqv5NRzDTwe6JKk9Qq
/y8SwkJ4/OnCMpNa+h2pJjurONpEoKIp1ICPb7MjHng88a1h6Qsd2cBJDK58
Io5QEnN7QkYSB9KtQ3jdB8VRb9Z5wqaa+WXujfY1SqPdCGhr4x0JVlL4g9d9
yv4TMaz95loy3uIFJNOPJgEez7oAIsifAl7ptwxN9AU3nkYhzsFB2qp74XDi
GW/Al/TCrGM59SBDZ4JuV2qmmMMuZL5qmJEYfmfVjexVjr+4YBcS/5U7p5Z6
RPTuR0aANZ8w/ZaWucSpY3d1KWwNXhMX3q++SiKsimqc7rwEnQnD9oPxZcI1
rTZAaUr/FMgUasMYgsqNpLoG3oahhSCMKwxmc92YMq4Mss0Qqgv8RvE9qbaz
xi0+zHTukbaIIlW++kmzq0GpR6QqehWmLSa/yzcM8zAHE2LkxY23YKrEWQh5
OZoAzmn+smoqJCLaum8/qme02l/JgtlbI2RgvB+2ZjNMAGYAuVy98TiRSpU5
k9KdPayOlVlAkaRRfWPzSXBC8fB8ZHzAGYdnIusfel6J5VeSFvrcZTbUYvue
q1XEk8DeqdW1e5sMbmixRJm7uIWCZZ973ZmHvcJ9C0UqqEH1YpipkzgpMySd
9q21DmuxHbNRFXmidkqepD0Nc8DmlFuYSVemxlOBH874j2iWvUTepQV7a4Wk
/BW1hJCHkKFlstSEyZF+YuRMF3OTu3gzaodX7JKuT1pSS5A81Bu1wC3pcgpq
1lN9R10YIvk81uKIV9WoFbx+ZZPoTJ3FZwTTPz2ZSN/zr8kDy1UYO9t6LIf4
WNUDtXVZLGKl7tjkyCGHBsAmIlZISiP7U9ovEpPL6AmXl81oEDKYmLT9SeAS
irpKGDA903Z5fyYamTMs47m+oaCyr/mQVhCGpxsy41LY56fmYsbj2/H0Ldms
Gwr4/SRjfvwoc+lWwpYF4TDF3iEzkw715UtXrIuyxqLBJ54G+/vDS2aa/FkS
nUIi+UFiJke14RZOPTJAPtk834TAC4R2DETdWT8AmxrvRkYYIkyBTIdAEDWC
SZzR63A1apzlYXhP8fU3xBdS0iy0sqRkYWx20dcSj4f0S398PFH50+g/8zo6
7yxw5n+ePsS5r1L4TAkDLAamJhkeYSbApVb1syIljV00pQQKHKmWZ1yT5tMu
9n831FpTa2qPP2wviWvOs2PkulJEa2UWvdi9PkzCTppehhvg04FlbOHiM+z0
gy4vsoJjPYjwAjP76rZfnJCIPJW4eWaDuoGPe9qugcZLoZoMGDSDv5llVATG
YKqyKel2SJQo1LtACRNqKa89ch9RuBfX45MPGiiet5YanCFZ8jl9I7AZ5577
xKQ5Nq7kJZnmStjHzfq149izfkEAemB+APSjHsj2TO36vM5VdnyFY90xX70w
c5NpiGTj5WS52E6F0pTiShgX6x5znuAb281Jq8Glki3eruNLTs9EYAtDJ0oC
p6S45YKkrJBq+/ZGZkLhNMA3vrL5IGlXCz2obMBsvGlZgKihsHtuuuMuSMXR
korfLYXYUhjd2z5QExfaHqaEfGZ1NI6Qub5hHiXe1OStec2JxnD4f6KLckKQ
YOQ/mdT7S9KxtQxdnXWwU9nonVMkSByYaWHjn5z8ffPARE/RKX81zsgxP8wn
Maew765yEjdiU40gqAALmZHdzZ11IVn0iphwfcjb6Fer9aPTRoBJsplUbtGL
wLyV4nze2btDE8hamCKcap5ieqdnPRWzE6ixv3okPkr8QQ6apD44IE4NoYO1
cu0R0GuT7A7fknPOgmHt5THNLm7YomDg8FIOFbqlKa6Wo5yx9j1LHJmAuHLo
nPD6hvhuAz9MTRU4SlamCaYYkRoybev2TCUWL98X4lnibn9SeBFETqikU0B+
U7F1nVV4RMg/DvIWA4EwtWJDJ1GYliKJVkVQtQjW+88v8QTZ/eq54zlz3zNW
BvzpKONElPuwR0dtXksz4R37UCtpElLRZi7+kp+YwHLburUPub0mu44jqaRY
RmEOMPSt7qDm5L2S3nQTVio13M0MeDVafyOGwW39AaNJPiHB5YWPHyJX6LmC
JO88eVMhs95PiW7YtIAZhzOV2Tbj1WTrbU743Wurx1uZwOPIiW7xO9SolhR8
8ZSXbqDGw6leoLOtp+eVNfdd7Y6qyDfKbOC2kZzCewrbbRkSwy9+TQ+s+h+p
KXtiN/WmZyHfVDxpuFIyKFN1uJikuLYb0rnRN1qVMhhS1hwUSJntIisrbL7Z
Xxr5MjO8qEYQd8K8dNIpNMrx2uJxLy3vgqEdGx1MBS71cGpBATSsGzJffjdZ
7yb+Jd4yZgNqWtQ+xE9+yIImr/hhfG8QXXk9OwLAHT6Ksyqzk7rk3HD+xbog
Lkql7TNcEzSsvPEA5NxKh1Vq2OBs280/GAdoDDlPHQ633ndCpLzp/xjeYA9Q
+zHv1lUV07aZgY9mSh2t9UvaAvf5C/sXuSPmFKLShWWZJMtPtjtvC5CGDA3p
CnZ5KKzqwmBcksXmhLPyAU3LbNN4tYEz6iCW70+009OzQOQAs54FO5Ux//mW
6YzMD++fyMRWEoMdvYCSjiR7utDxr79CEPil3Xn/qzEJbAMkePKouZkn/q+y
SNOXSRfDNCqj3t4EdQDhgsvZvfpDh8YIV0NDO+Il0nQcRpv3k3yZh1xhmgU0
uEmvNUKezHoww3bRKhbRUKeu3OFk4cyGMPOpSszl2gyqEHrE6L7CUj31iisn
kTT39IIx9M+2ZcKS+aO8dLeM5WI/I8zsDUUjvS3pzNUGXhBTW4PZuwYmyuI9
bj2xSo8rrLJ+2uJg/dAhUJb4B3BWwYi38KQiId/jK+wQ8deaC+APW7Z8aCIi
oZtwCDArmpIPLigM2LACoYsS79imABtW6rM7C6mMsbz/NSVi84Ey38tk9/UK
Bbe/eKZ+Kcyd5iFTfybQMB70Nv4iW6v7LZlSXxojJca4C9G0jQuYZ8NIfgXP
e0FnzYuAez5iYe45yyv/j4BxFzQN2swW+gEPx8Hg9NR+GPeX6lqeXXqdwcV0
QwB4KCy65kBGg4nd8F49/NLj7XT0KOGwBeeANNTeDkn6kbGOXdxGfayPeXDL
uXHxaG/AsWHVaRcz8+uIzToi6Y3ZAXbINJrBwBV307eh3opcEPaJNxEQqOm6
AUj9zM7/qLfDLFUxkQCT7zAtmIgU/PKSAKpG6jKcKFiZUZ6zWaBh7J+6vlQS
f2lNMxTJjoKEcxedGhbS1IffAUetAEcx0SwMMmBEy2pdhmweOwuZQVHXmvT3
CH1jW3VBi/DAOcb4uoMGmDarOM8kfCrrENJCk6SqhNMOzzwFq393xZTgzx9t
pj1QK3Jic6aBh72NASBodu9e2ric8cr7EvPoWgXiNfGU9qV7ES0MEhaoRJYn
nW6V7hvxYeFZm+fDKp+VR92MUlV08kpJpXGDqTGCAPyYIPH+nhfh379ahFvw
0wzBT0WqrVvI4NwHz7X/VKt5rBxlSSmpflCGsTrG8ecxEWK24FoKfWzLHDUz
VfhltmMQOMyRs/H6JiXIepNDMQGxgffo0AbmM9O5HmFsViq0WP1a79NDLvzS
Kh4DzG+gdO0dHWzkUHpqQD2F7yVMV2+RwJQQg+BiefJIJMDSLjDeHqZiUWbV
lEvZGrRp+alqND6OHjoohkGagfFJi1Z3MqE5gyQSDNTwID58po7oPhGoDu3j
KUmkaHCAwy4+l+ChL77xIKpiIR2poQgQSfv6vAErqkl4+wIU5aKuLXDG3/9x
wx0rnnuX5jTjCo3Cvtv3HW52W/YJA8kJ8ATVQQlEF+9K/oRUWDLAg2P0VD4j
k5mCY+KUGzO4Z7Q+WqAI1yqA/KSlbfF6HiZTYs6pMlX9kj2IFr3yEEdLcbET
/G+tvhbd85HLFD01QP9tG5CLJsYrq+LRna0j2B3DrRv9oZKLIlp0iyM0TpSr
gkG/BfCwcArWMjFwbyYbL3tA895duI2SowNDuTHUJnNWpotLJRuZ+/I6NwhR
/bVtD7gBazH8nOqIqGnozPFNG5wSl2dqZ632cKJhxuyIQXIAIIKE82rFFXnk
KWwg1nTFG3cLxocsyxUJnrjk0KIDAN3kvDwLpgtMnDhmCASboQhJlA6TvSB5
mjETeQyw+D3u0Ja/9CK46wSDWU5Tm1jEghWqxEYO3umLt53Ke6PwO7TMK8oT
hlLrZVhS7RZbD62I3tDkeziJzgn37xAjz0QRjQURDOf6C9XNJ8D7MaU55okH
uvYu73bj5CyKEJvi434EAypZ/Zjz/JYy2KN9SRthKZ3tZDQ/ig7tZFCOx+Gn
v57UsDa4OzdD7R61E8Wz7nZOeGTJTcKl5c6FtFgouUd5HpnR/X1x0m5ELXZ4
AUci2Tsb7XvWVQlgrId2PF246HuKQo0NDbJXeHM/bgM8Uu4omrrMXeSuay6n
WMseOm8KgHSPCcgk8+oi9fj/JTup5lHdKGVViPdCeBuNDqa3BkeGfWATU5Lh
7LB6okPc2invXg/H/x/QQwokEjskykOifwNWnulVkwI+6IZ9QHuuEHG56Lcy
ZivCRqM6FCYD9NkLfMj5VeQX+wq97pG04YGPpaPZgbkwfP1L/E5ik/3WAJwu
R0oMqvPhHtMhCoz3lSv0GMHQ0NcNyJFBS8ixe16cRXFmLp5E0dHRGHBdJfrQ
OZhTno54NJC31n4pWD8KDb7Mgt7OX799pI4c4FfE+P4mOHGs0kLWabAo9h6f
Xez/l4+ypCCxdgrFqH3mQ0g6uqgVuDsmf4N+PO14kIX6aQGofgkdNOTYo60Q
xHNRbGrCTWi4LoPyOzMSeXCgyK9WHbn3lwYYrzCTnoWLdkeZKLbBpINhrdgr
6U1QIkrjMxmAFcKYz4uvSAyUI1erFMiEqnI22+Q3vx6u2hMacUlE+ndl6Zhq
Yfh7Oxd65SW+OSQK9dbv3jZqp4/CZ+MGQklfjakgKt5ibbmGJi/wpL0TaERT
ZjIpFCh1FsbZCxcutZLObBHZ9RLYZJudsmbS0a98AmMTEdVT0XTkk83DJbmI
WW+zOUDKpJswglzHWmmaIu4rtduakUdL2TcW//PJwZTPSEH+R7f3NzOWXfJE
EiAO2F78onrYkpiGtGYEoDpUJGXxsIYyuEGpUsTJD75N3eI8V8oFu8o8SH3i
y+XjHXLj1sCQAYkZOHHBd7qBHIprzVuoQejERQu+Q1n0EXc5OMgTi+Tmjhj/
lNpnI6M7akTMnwJPgycVCrkyhp1Yn8NuB5W418i9YCBYQZhEXhFiIJiqkC5r
tsBtymsYf7sFsGdkrM07HYS1yG+2GahglSOFmiB5ih6mjCg2rBaMaosfWVTA
Qs4PMwReyPm7DlB9mkIIFhTboYei0xGSkHnCBT8/09+xkOfL03jJw76Nz0vL
VS5P+btuTxg6fGZ+7tF54gj+uO+qz5CAWVEhmNWvGn4DxJmNCNyPDKuxH48p
cTm71j6c2sHcparoAltPYsvifKkM5nYu6jem4Ofw+qCA7QWsdMYDh4FSfKXk
pNQ3r1Ey31Rk9RzBwRl33GjXJC45qVCz1qUEgKQ0rP8/mQSABfTXPcOV5XUu
ut0UH9K/Ujg+pTZiFETdRbVMKaUy5zSomzm8fU7zFdrWkYIQ1gf3qcEOtdeK
heeyM+WGviViZZMMk1Xc3pyBZLuME96uz0fT/zFQ+r3PpeH5gKKNOYS/Dg6l
brzq9fh2DZ6wGMAz8B16QjVR6aRdspA9ywothaL7bMERFoPtIl6EaIq6zuTc
pT9YgDdqAjvMjSfewPbbblLUI0GR+kFFvPDa2J/5/gWIU38oTN7aI7yWMEzb
0WD9PzdHeBG2KuNKcIgMSV5CSl4fgsisTA+Vq2j/5NyUrujhOzE8tOLipIJx
YR59OWA+1u1OG+r7mRct99yGDdExiHoGDBHVW3hWe5tp4QDklITVlbW4wrhH
PG4bv16/jguNbR0U1S6TvVZaG8eBWp0K+okWJqLWc4AFu4KsrOFdPx/Vw5WR
SCKozTiqPgKyJB2XMcThyc5QxDIuqSvaUrwHVw9DDlnwW/eqZU6KJhFRAnm7
t71+FQkvDxEbU+KBhxGena6hVibH1OOo504UgzEXvKpQpEtJ1gMrEjzIbkux
wL/sV4qCjc0KioZCE4suHSlvya0w7ObIBX3Kl4rQOwRvm6cj2jbbisJvLgta
MYf2ozUo9ploUpOY6PHDaVcaDXoWGz+suZCS6NgC5U7MU82UnHKMo+oARmBO
d6oZ5pobX3hpoKBPsRZ5Q83hTLj1MEmaYERwixdwv0oqmjR+kIVnAhDhjD+j
tpjcd96neuNheR4X8TzzcJGo0zst0PGW5eCR9p8htwsqdWiJCQko/RNG5pV9
+sxuggCrV9a3Sgusy2S/2rwhxAFSX6Dzg72qJVJ3sPcVmBsCDPPlMLLT/kJ7
BKi65CIHoqwtCpC6ZpjSI0Fqsf351PILBfYBj/fydlil8EyD1jtJu473jrae
M3nS0SRCiDquICSRkSz3mtYr/9tv0OOvH8zGMS/qFf6t/g4jQzDsU4B5vawz
YmuZyHup9zE27PSpXqslIXtv2QI6XgzHYwcw1858AgS0M8u63HTEsBmA7EBC
vq0kR2/KDNcjZrmsYr5UbGrg4U75LSR/+xSrxAG1eojp0/NCP99/dyi9RMCg
ZzyPTVvxpMSvBMEHG6AMH8aqDYxUlh8aaldkbDipUQKgrML9e+94qsH+FIpd
C+Aw88wyuTA1NQFBhemVTR87ky9oMaVZIq7xIjcujcctR5q3oFylTog+VzuQ
r25Bpv9lQF5+5PloPas8Wc45SaUGx2Q3dhQfPRKIVgTZOotgd9eulBb1tUlT
ztByxyaCy95gRuoSkL+iY6fano+ovRGlDXstCybmBhmsEu8R9/6U/J+brr9/
JMqZfSRt7M2bQ6eUYKwJwML1Z6j54v1kx8QXRKiN2gIveLAH24O2CwcevcEM
Pb0w7L5GwAtUKL5iLIwTNwZIFXdUQjuceketCyJkEI3fPvmuDhR9I7vtYccS
h8SaCKPTz5N/7+UxXbaa2Ly46uzDBbGb22KA5p1O9x+l81Y7awNj/PedhusX
7EwDMQ+c2HAS1v2DiWqx6j7I50nGIod7K/pjJP4/WpdStXfMW7D0HWjr++iM
hhQ71sOZ7wHrBL4EXjrdnGgTiBbWru4P/SpMEwvQOhs51L2oqTczJlrG4QYL
if8LOs3TPHiLNTB5hkGpZjKRDXwEJPTuW3UC4gEMAZFkr2I+30Ou7HFr0Oqz
ghVuEL13MYBx9/0Ut/NRUfo+/XQReNXtPtck7R5jMEYbwCcfqtm3QSGVivP8
jGKtKa6k2JoZr+85V4L+5ObUZpEMLdRMfLdaLTqtTuVEYDr+NlXVRE7W4Zzs
msVRmD6iHwjxEeWi5JxFtSb28rFd5lw8jGmwHsG3lS6kSsryz5BJ/e18NTQ0
iP0l7YmCANLICGFrHyk4sJKFUKwPgXdPDlSeHDT9KRpnKFk0fDgs6opmzowM
X9wvatEfUN4jgcASbaxYAYQSZxY9l/5Q0TiaUxTAHaz3wIPGxDeSHTAPLhBM
mDmfQ8ZibKT99XjhbiqQ1nqpKvlWySEFabGrbIqHZpwn4YhpBn5oeald+lCv
RsUMdC9Ao+zRj6vyNOdeGruiXq8dYN0gYZVwWICkoCgSHVV8IkObTy/2HxO5
4fI1+dh8YBDxpJKu711UMoSA0KfIfrplmXLbTDQioEVSSxMbwIvP3CJaxRUO
Zy6/trBvkhYXAeT2XxEQWex/LCMehyZ9qkgn3qJdHEehfNSQxvl3amSAUFqk
kMQkJCwUdYHfPGXLi/7XxIYnOyjelGioDK73M1IWiDLnTgVh0JpBEycCb5aF
yTVaUpKiNUdHHEyBBCYHHTnAg6wLd4wRgk5d1a80L7xhG8rOrSBzZRUaCjbz
aFJhY4iPZYGl3AzkFHdn5T8OBp6uAnSnWQVr9PzVKtnniVny0xgcS8nm2EqF
cG9S6uaPgCSPj7//pQLr+H7+Lj746ZMyPwaHq6DvWImv4VBAFOrAsZ1fqaGt
fr4/mZJPp3UOs+zYxQ9oMsZqbbeTJ6lYgmA5Bkhjw6OwxUJxLzs1V+Tw7T0k
dt1xX4hNF2fUhJRo6Btn1jzH0st8fevyyQfFXW9YqOk9gMIqnbpS+4ijT07A
uTZvVNVo31OYLtvr4mggM6luTxSbJn0q2lxAsXM+nr4bFSkI63vC1hXiyNrN
ZgpeeWA2dyNcmQW1qVKzTcqcly359wBEDPngyn/AZqnuLn2Xe5B6zpgTi7V+
we5bsnkf1effvsepuN8lOYJz7yQQ9fvwwdsCwy4FK9Sw595hB2l6vqCQsDeq
I+P1PHqT5o5fe1naKYBlXaSB0sgORWZ0eoP63zqCIFy2899M/XBd+tbNyli4
8zeIM6ZzXDgi0RA71p4ZImuOMsnFA/Nbrm4PNXzYr2MJ6L6oApU2gXIYd5XO
fajbrk0KrVrZCpSPSgQTtaq+HvXVu4qCXIbnnHPq1B6i2T54coTlmHHDi3/N
oDrAFpf9hathENEsSSFPPEXU/UwWG+OfG+a3uqRjFZkOBFvXB6HCTDfuT1k5
d7MMvw8Owgp+zhe+tDGBiGx5E3viCjZsCOB9boW3UFNYsiWM1zLyrvfH1OWw
CLjfze+ruw1QgBub2FARXkgYEWIWnbRYO2ilDI3r9JD0KCavo5kXVNU+4ugl
YcW3EFrf79dS7OiA+WRYHitwbt4JAd8ayTfSCUmI/u7nPMj/J9ArnPfbd0m+
gumI2GlcBgqq9G7xbfnSD+5zxhMy44tRtbp0gQI5NOV7PZSDxbb0yZmyNo9w
wZVoj4uk432valZ8v9IsZBqpi7WYA3AQIPQd8qamWBHecrwhQNoEShswDwLO
uVZR2iUfuU11X2s1CGTO/AVmLmOz8137vlyYc2ZGDObHp1H+3Si1llySp/69
rSEaYkcs0NWrcmcyA//MY+ZN9y21KdEtI2UaUaIQgpmae5tiyveRkO1N0Utu
coIVMrIIlIpel4KzhtS9d9wBMZb9oI/qw5S2/iiKtBduEqwrCdxaQbIqUW2f
u7VMt9HSlE2+b6y3dulpX91De22U4TtVVCQA5NOg85VvGhMzsW5XZEcQEQcy
OUiBaGZbPFp3a1HHZkxhtYntBaqYKR9iE9NMLnmcxr7EvxGkQYrriYS5pY2n
BsynCkB1mudu0PhZDEUHM0GyrltwYCV49d9lri4NtGPoRc2TsR8NB+lTIUin
CHnYZelkA+ER34FHER+ZG4R3+Y1QW5gPCRU3DRzFXDWKV3VzzLbFbzjb3cBR
McUonjgOFMqUepFSPJzW+2PmFw2CTmZCo2YrpQ4ElzuAr+DjYXoBQPGeuvTb
8/ZltvBtYOIZ7UNXJiFPd3K23vVhRXu6Z2kp9mCItt+qj1FcwwRw9w1c5F60
rKBdO4XeneAxOtw5bucw5HlWrOSAYifEB928hpvQyBmNCGcbtsJZF+NTYDuI
JTwHidxmYp3feqYoiXLzYRWsX37aZosww2DaQKeAeqjinpUzLuJP3mdLL5SB
sVbsoFi/znqunnm24SSYo2RMmbihJYa7boi28HE8IBkqmkq4JRmmVxPPeZo4
G4OnvTtbJvEtSxBgcIavgGeDSv+T3k85lqD/qbwnBbic/LxnIjCjw1t6E22R
fGYCyP5mb5DnoLF/BRsykyY+9Bf1M/qe4R12u0M4WTiDuQKedqqZuzVxM64e
G5URm9oj22W3ti1TtR25I5y3vRtAehppBRl/ifKEGZ6Mr/6WohVD62H7NqtG
tUxq/WJ07r57nS7IFFYeMr34ZjMro5HOqqCDgJuV+YlVwYZ+EgKorJbgTDsM
/bhkv09fN3UiHlIrbvtTK7sm4n7Kn3Cb8yOIvxGanttLvUIMZ20pa4WCiUcz
dQUPsvNVbp6MM9JhzNf2A3UUYNQwCVzXX1XlTJO4EsVw+WoqUWe3thsgLvN8
xCoAf02xJmBk9oNQu/Mo9S5pHUc/hEWnGr4px3DuBA8O6fcrvdyQa2GJBV30
ppJLjsVh9sgDOHyJ6gPH2C/36u2AVOJMaj5a/Qat2wLG2ppjJ0dDa5BkyX7W
21663gYyd+EyqKtDFrcmTRMjaqUDi+jdKzGV3/Fn/FDOnO24eqzbUWXgJMaJ
Y39LqspZ5lxcauwV8E6gp6ZPw2vj2Xg/Fjc+u1SKhxeenInTXfkvVJhBn79+
wRpQU3TqZ68J+tjXHn5JpX33q4Gi3hP6EVy6pOgYkBc0O4at/7TyTbC3/YXU
ETsZ+DszXtgoCsNLKYgEsEmDnJL9pERF9exBK6fDtxKEVFnzNGy/KTC2nSR2
HPqlE0s9YstsByAA9vyQFGfZJ6/CyzG+gXWr1/gBQhIxCteAIDSqo4TzxHhk
JUm3qkJz7RXQbJ466MwkByVDE/dRcZWQls9QzSZu48RWTuVcvlVJu5FOELWw
R+anPfFIRfovOLkGcZy1XzWQOj07hjntgUt7JqwD+TviHqX1+m66NJnOORO/
jihL9BBOq2CT4oK+Afc03bXokSddS6nFzHItkgCuIWBAGpnZHC1x9EO/WIm4
luJNzofUetRhbgIynqNcViq/dYigc2hESW1TdvKcCiCUL68UahLzw0RTXCPI
3W620omJ4lTASsYcGp5oEOFVQeKb7AFPHG0+nPDZtXqMd9PBn5fENgXykM/h
asvHPDHIBN9FQNcsyEq0hptzQViJIl+CmwxBUtVgPn2ZIU70eKwb4QmTJBce
2b0hEoK8So+lriSxQw6Yf9h50DWDmul9mx6cNIUwVcwrGjr6RVq6w0iVA+Hv
3yx6M876DNKqAoxDfN4yAN7ki6MZHBygeEk9uVuzhveSN0KUbiNvhi0PiOsd
WcwoEgWvWio5V7OpTte3Xt94B2N6SFOBtabwAUK/Pzlq9zTMPUoTx7Lun0/c
en5+mHAGf2+s+YZXAMY2WirHvejaRbZVNN2mMn0StkeRKjY56ZdqOcoj/67u
dgIUf/tKQRPUBGCEPcn3ox3FbctrYBCakW3Nk09HSf+VTqMOsJlQRQNafQYH
DTB1a5ODu00XAzVjE0QOPgjDxqPuQBK2KGrxGVfrt/PyzfqOY4CX90QwvJRv
tPi+lg6cjILYigVSdXcNvVkKXcd7fBJ92sZ7V5o7LXf7RW7A/+JNHm4kVKUi
JTeTmSsr1+0sVh4QA+RURMZ4TxBERKcYcd+b2raeZV3VdncxMOEKX6lWIHZi
dTeDTYAgQgy1g6ZpnOybTTCiDJJgdY/MWLwMeDfPNLUJYiWsOSf5ue7jk8ef
7QedfflSXoGplxS85Ko2ix473k8H5MibkrQKfSeXwWjgYau83F51gqViUbAJ
W30opyhmD/BwRVl43bmzRy2bYShcge83Q8OYS2WNF5AiQG7LwT1gLODeV/dO
KQyaRZTF+NRLA/9mW7dw1gycPesG3umBQccomyx3YQYeu3vhHn2/nTTMTMDo
YX+oDSWvJkDB+1ryzsS5A3heNWZTrdiEH+clVNiBpsWbqzIS8HpSNPrAmmlI
8CrxV+1/T4C/3LaTwKGI3U1kuQlia35roo4JiMhcflptd6sgig3I0VsNHPg4
f5BbfvKCR6Gz8dJTMHUNmhDObK2feIr8ZygL+U2qrhzcCi/feEiUNxFxv9UV
6DOuev9OY+3VqXvTTDyF/+zheIxAmoZJ24JDYqon+nkqC5qNtJj6yU01M/n/
DtlzdaM5LkbtiUkZkeAe3wjb2tHT7sgiXrfvxKpsSlzuyocvstFNuQe9wyLk
2uszUnkKrSj5bzU2yEfL2dB7q9eY6xFpPCQocnQ0rPgnEJLqIEcHi2F6peIB
Lj0YcQ3exZw8KGKzMNB4OeZG/EVQyt81AqpT6R9Ymo19H3fYryXOgVjh/Smc
nQKt5GouVq1nrJIsupqltzje3Q23z3kI5M/nKloIatGexfQ3W8dUHiXOfCFD
Fc3AS1QcpMg4SWkBfixKYYqJsnyN7rseAqUr9h+VtdBKim0TDTZ/GHZpkqaI
NT3krJ4TxZfUHQ3lFnZfVxcbWHwGzMoYq1Y+UVawlLS9PUmOb5qKZx/YgmIm
NypgnU2Vvn0TMQmZBfcrvM+qI630WfZwC0vB5pF1sMx2FuG8KAtPmZNID/Ku
qqaTYTvfGj5/oTKKfpTW/GokVDKT7PcVf+PRdvzMOKgfOoWSoT+n3sXdIwsb
Fzzt88B+5gZM9YJ1RlviU/Eg40BU0pIRuU1I0ByBHpJBIpb/mWr+VdVdWX2r
aRc5jdckY0GfV1aCNtD5cA3f5lRdcP2dNEhY+7KVFd/BeuGQAgg843V/GDxa
1sxeTwXUXBdTryDydTdZ5LWO6Yrhfh3NdnwTLtn+4tO9u+5/jwOqQOs0bM3I
Hy2dgxh6RNq3pApgrsjeBqz3njIUtgkUdiIpkFVUuqrlEYMnWDdItoM4WBo6
W6qyc2h4GTULP6utsFLvYzHMW+PTRXzsYF6mmbyRcQrjPoAp5/+J1UR/vMAB
JZydSg34ZVk0WRQg3usur5ewOgecA30Ian6iNo+JGPt0UIqsyBr8Bs8bnHTk
y7Ak+KxmYo702RVqYimJYoj0D1DMTbeDANnErcSWkMAzIkQN9QGiO7efRMSS
pcMGqb+djqPMAd+keQ0/4E4V9ZiT9XfuDTvk67/ecivWO3dZ3JbvWhmrn01l
m2H+bWo8qyV7AD7zEinfofWqIrwzqk59nKpXfPAMiN3qhvYqI27bqJ18NX29
cGswb4s0xklyncEKuGwFeaVEXHiAjjPMttcwtByYKRZFW/7DjRoqr7WI400Y
tMIZt75Ysr71w9J3wzjWE5lMygzorsRLDaPDEGvlb1dUHMCp2PKDOTBODL8H
aIcSb8hQgC3Yh9Qo7gD7gBb2qM3YgQVOFb0tMZ+F8Ztz6af1YIx2DBm+cxup
nrnrZo+6zBYmc8QCcviIHRfXVAY4VfyIbTY1eWhBMxe20DECpqktXfJAsJe5
zrgSv8RR5dpRdPl7zKv4hVo8XC/k4F9E01uHyunds7Jo5V5REHj9v0D+u3Lc
6PJ3+CuclSzvJvoCVYYKogmINZFh4CpgjpePDNJeQ3ybQOTyBwVIzfjfSvi8
CI1G/dbzQFq08hFBddFpzOJ6cQwjCoMqQEFIR2KScHgS8b8R8lcaKwzius5E
xEhvAi7aSHKs6A+FpPjwAe/qiV3C3/hlQBMYI064+gKcQmJfjEv5vdCP3pnn
7LQLvmvoXlVidV+3fHbH+8C+RMzDdBs8GBjpSbic1BkS3O6gefRqb26Jh3fg
zB8h4uI5mLHLbB0LsItZ3vo+3JZ+7xnZeF8G8llgeXS645FW0pCi+TA9QwfN
6rOPK7cv0+JELVIm2f2rlTRaSoBtWGjTQol78mKqRb6Zxil4q8dF88nDKu7P
zswJ4qHCfRu3LvufjZ6bis2GNoea5wL1VQK8gO76ge77ZS07qUSeeZzYWIYF
ljVyju+OxCi8FkzrszihXbg4cObkIBMAjxKC9dt0G4HlB+TBds2KG/vjzwQl
/RxEpQe12yuOSfHza8nPIPJC3+Tdwcc+O/09A5sAYj5zZyqrmYmk1rp+rMPt
LA+Lj5cNYJMSgPqoV1Vi6NW7YhHeJDn3ggh9p54t+OYDHim6IdJD3d1PO59B
lpzZtJfbrf1DTPheJmVM+S9wMyEW2sRX3O+78Q6+JDR6jwA2/WHT/ioOCopS
eG70jp4HvKCmz/RSdBSO1E87w6bpF04EU9J8PozixjXPtDAvcbInl4RuUFxl
8/79ZHO8/zXKOcjABNgC42JsQAEPLqxNWAu1x1Qix/CO0mzfHfbdqbfs3Z1S
8H5zKU6eps/O0sg8+Ed1rRleA3tK/boJJo8FzOlcudz4v8PBj5B6I/3yNShZ
mr6kaFbNyvIilK+hMwrwPZyA5iK+aQ/btjlvPXZuHqrhjvxyHJ46FfC1HZTb
lmx8+pXFkHsmwiiOUmHgjYWasqDR8KXAbJBu/6koc60tDSr2mypVSfzfBxbS
kI6APSS2vH3fL+h0iYnhb6X0fwFvlW/ZFJG/pkkxSo/SJnwSzIOEtVY2n42t
5cKAykKgTO8WdVBKm6k4euv+BtUluxzpH6jGRydJ82hCxotxl6EJY2RIz+fv
HMFoRKrehJSaSP6/7g3T1tstvHLEmY3Z1SliJKNrYhZzRO0nMQVqrkdQdyBD
rYXPuJeusiVZQcoQAl56UIta8ZsEEYTdQewDPiyuQVEN3Atm98HEVnPfKnfX
hAw2sQ4uIJptJbDyU8X+jgPaynuopwrrakkn4B/lK1rBcf0PnY/cnScpvW8U
F4SiRNsibj5WXRfM0itqehafv4KndfcFFNhjZvnrVbX9N85QF+j0nnFTpIU5
fF3fSm8inCtJHlo46AX/oFDkpPfoIpZ/PKkhVARnfIcNZeLfvIwCsn2W8F+9
7Z89yFDH4pt/M0DFuOvKmKW/lPfSjJAI262reGAzWwTK2IODvNXqfx87S4n5
GlzIgsuujhgHO8XX5cTyShHNmY8XYZdS08WEM4KsGgQAlvabXRCpF9fZuprI
0iAahYdz90x+nDoMbkJwn9BTsLLLZh5tWyMa8O/HCTqV0lY0hUYyd9tt9WiR
iGhaPNC1vUwlu2+sv5hCFWYJlPRHtrRaD6sC4vmK3OPNH1REBAR9Xhe7TrG9
qu4qil+tUZJ+hLwOR/+WKtG9YdZOBapjJt817+PizK4xdJMj8JXqQUPatlI3
2FBPVJho7Y2tf1LKWEvePwvEQx7g9pCeHlHRVM8NPBXJ99jgDrA6qirmPCjO
dD7ghWqUsr/kjCCpHOT6vFXddzWS6Y46/msbihacwAdR6EK0qEzqI9SmK+H2
NIJt0ygtH9p0P4Kojc4NstAkd/fl4wLQkFe8lkuTUcWT/RqCLsQHV21d4zzK
MeBVF18zmuLZ8R8D0o8jgSh6Lqe5m0SbNS1s5YbDSQSwyQfIJVd5BntSBHiY
nuaPCv+pbPHjDF/7GOtYUXVaNMi/UqPqxm3FVNSu48Eb6vRrItB+xdhu7A90
fFkonyG8qzTo51FQkPzra1lePGAKG5L+55k0S3E+KJjlHI+bFK9vKwPBNI7T
r2IGuGT8nWMwWNPMLSyR5ERNFoWvXkP58aEkpXrmMFGVpJGJ8fkvL9lA4IrQ
GpQ9noSUwvJeriPD3yycFJ4yYmE5Ptm7omQP0AuyEVcwWEPVlPGW7y95EVRs
WL0X08pq9MrL75AGJx2wO26y/TooNym6X/J1Tb+C7etDac4KdcQ2ktmIscpF
OEmkuzRPXxe1uslo42cYZmmzywhRY6kBTjGMH/xZ/A0EUx16Fw06pppc+IKI
xRs9JnkbsxaQRd3/dTxIw20F68Wpa7phUW87xRpSxvKz99HOjnPwxtrfkJw4
K/5WR0uwumtUvLfnZQJXKS/98biImlwBrncVKI7uDQcTEkus6IR3PLYTbPV/
evfEiGXp4F1awcGwb+cg6BZgQLImGiO9S2FX0MCimvGC/J7wei2h0XdYUe+A
XpenLRBRh05amDhqYlY+o3p2YsyDkT3ot2gOnSLR8pIXF5QgAoh7Vq39FCJO
VqysnywlRkyaB2ayFbkodfH2UVYq5JEr8o73L2yLnjsManTkx+xtwYA9xZbp
13GO8mWcmzBeJIPwgBeN9C0jBJPBHe8sL/LHJ4M/k4NoErL6oIKFO6vXko3t
rXOE5JBAPG1vfrK/bsUkBqqqr0X3Tu6Q50S1QP53qJq+OuNZoPK4REdVJ2yH
NzPmeKKS0cya6YpAmbdpiOaScwpLReX2DLzLSc0Tm/ZpL+rjlmm2WPqWqzfZ
a8aFbHcsaYntDokOYdXeXFzhGsMYmNTlwVZ7ryAA0gomH1wRMf5Z9XAr3Ox/
aNSJHjd12LPw+MA14RrAenCl/xhX6siMG2tDnPi1L++DFV8JpZCfcx6brTj2
Mdn5wIHSSxXB1hYtFxZRnOgtuFrFXaqpJJ6fwRvaWZD0vDRjQ6Vq/aNEeEo8
HMmZzWy007Z/WN1If3+i8qzm8UKTVPrBDg3610Iy+ywIkCsX3ffoN57+lEGZ
UfgytDF/m45/aCTgvjp3kMDmttHNAs7NNozHwwU56WSi3+s2pSd12BOb9a3o
fFM2e373iG0/ON7SCc/yObXokRPQZ9P6dFzqKfS2WOANwuWiL2ynKNNWuEOw
rl5Tu+AOSC6e28syVWMklkNwo/NG20kpBAU1SxwYt90cWWs0b/xRkT2APU0s
PfR15ajDPfwLuPfk/+4EJB/pwoGipPuW4u3/cTMjhIEB2a8hdTVvXwW/VEhT
U7m7MljmB+OsJ9JeAhcj0o91E+3g2BMJj7lAk65hqgOPjRDuOWDuSLLrf40G
ji1NbWGxiYdUW+yQwijBdSwHrLJDD3CJsoz8EcJw39UnQM5lU42DTW3Yp3JA
EiT5nNRpZPbUYYou5liGIvcn7sySlgpGJjruHVpIPptVDiBCJ+k7+3/OCmb9
ZwsppZlIHMefjyRvTo63vk+KkS5j5Zp9HHm0OhWS1xgx+aCCqVRv+/tAFWQt
KTgSJVZ2RabcIny6gfYSN8DsfPnzmpOu2xIqoITdEuIUS8+fgRihShsQf2kC
MDWpc/5Vwp4chBvA0inned1ERuCy+GJmqQIo7ok/FWBhO1JqBWLr/LSXjSlX
BpnbpitCsMRcrZI5ZcUWfeVCy/mStPnoZmNbvtDnAvbWx9Y718PWypEFRUew
VtBKFELO6/pu9GqyUm0uqg25rDq7wSYODy1mg8xndP1AnVv8ZOha+4PqP5Uv
djYE364sNvuvVcTQHsH03JrgIC+6hgRW9q/TUwO8iXsup6WX+Iv3u8uyMYGQ
KMFXue+lZ3AqqKnXdeyIRi1Yl6CuAbPmkucuOTTdrRTNKrEnoeKSI9XkdA3r
SDMK0pPeqUWC3RO0Uovbp8h7Y5scoA4v93CqWU+HhXJHRXBf9CY93CKcFXIt
NRacgL7D5n26b4CYeYJBQJsoUiKkSDWAx56Yp3Dy6XruZyM80CIREJ5jQE6Y
3x0qru59NtB0ntuTi+MeN5lWWjQP5L2pfoKxMW5XUv3mSlKpwe/K56AFP7tb
vmaoxHQWEBESQEeHD0DTJIdvzB7fBA/IZpv/MRW9GdoDtqDNjejBnEENj+rl
Mstgo6sYvpayJ9C9sFDLFUcl0Uqr+aREo7yoqCAZKBOI2BZUKheK1DLn3bkN
SgjfteOmbd7LnO0a81Wvm3qWKj69/mh6HLFDGGr4n8vLhTULa60/4R4xiK2r
+DyPrcEFct8wcAQKRu7UgdwzR+lQMxBKYWDNW1L3fjl0+2w0i8h0dtiTjnEH
nplJSFbaITfGhG0hOkodDUE5X57OHCTHJaqDkDmNJJ/QAmQ9ELT7VjLczQ1w
NqD8op3BYY9ppD4NZ+AXocfRO+OtMAee6buvIOZdIhO+mAkYYKUe20o4W2Xd
+GaP4ylZG8cYWkO20y8u9bQouP1B0TI0Sh2MI4KNiLHhbFfajoUEBLH9nYi9
xUTBO0ztUytSIlAC4/1r9rXWuQC0LNOIloa+eFuuU6fvbpPna30zqVoI2KO+
9Gyqhxzt5sCF+WWHsJm6pld3w83gAVMy8si1VUjTg2VAvlwc/EGLEDXNiYtN
7ZP5qf+syYekU1/zgQ6eKO2SbjmrsFCcESoaVbbepbqERpVRsBJLBbim1wAa
o8vVI6DGffNYjQPV1ujlTqeWYPeemyoZhmimriRTf6S/Nf4Uj3b4zX117sNn
ndQDaMHk0x14qgn+UFtto8pRiK5P7EoeKR0MipYR7R/h48l8DuWor4vFp5Rq
57Znb0jQS+mXXS2A0B4mmWlLWSdddzvRwzj7G3NKCjyep4MKgnHZNe9zcCJ0
x1CpEf6LaHhx+bc+OAx/8pDom7Ribghc5mMaBjUw/vAm+6aZ/RXyiuf3LkSU
R9+b8LF0hmvnynpIgUYelfn6+q5vvi+4Qk7Xh32ppd8K21VU/K5qnhSwPeE1
xTBjJ6PXnFtyndHFpLrXD8FQR0n02NbhwhKMoQjxblwyh5gROeuyYgvT+RaD
64aVjdB5EXLi/KrmDV9AoNEKJXxnwAfHlyEMlZVfl6JeXFpuMiZVDq3kgcn9
X0WianGzKcl+SjjvT6GR+4kE2j0gQCwxL+RoBjBqA5GU/pSou7y9OtiNL9Z5
Mn2QMT6iP7GZsOGkxX0aFbcpddkIGdjbbji3UcyItSFcW2S4/eoohdbIKEIa
jy3BV9P1uxnDStXQBeH5la3lH52MPV9XPklTZ5xMRJSNckvxTA/3n9XSLUnW
s1Fi+k8mIBMtDKYCNGFFHG38oP9tDeFyWtZiOipTDkC0W1f9phgT++jonj1Q
/r3gDI9UkL55VkPU3jZg7is1jJWcpKfsWpG3+LHPJeG6Z8K4X/2kS2oOOzXy
sA60Wa3TojlmDeEUTcUrfBgVlYWg43lSF+d5DWfPOKvMlFCxinrxJbjHtLEF
0a0TzsXbwjdQWwtztM7blaPt+pWPFkijPEQjlj5iCy/KjITDhjg6plfE9YJe
jUbhKOoEnMpRasS8/apQz4sahYi76fJgm8R5OHL0FsUI4I+iueMJkyDJEfwX
Ckx8X5yEJvL3yJDx+FrOk4sbBFID8s5WAPS9QQrrFkmJdUSs8Uk5FRZilR3x
iQ/m3iMCspbWzo2Vtjk7lNY3aQ+21BNJjKZFPKZJ3k0HabTbxgXjjF4RD+wL
p4HX/zO64M75tZKkKShrolcNXWi2Y2bafjaKKehiVad8ZyXPJsXup/pSknNW
pRDRi+iu3t2pyuEN875/X6o0A5lp04dS8bulAcMqZs4+wnVC5A4/FijH8VYO
MKTPOo1eXQX03UEqb/dXZrsh/7CdqI5WmeRx+vtPzf/N3fkuzLwwubWlXqJV
mx1y822fYendhXX92QOK7ogit1YIw6MUJPl7to1CXEC82ckVrDTQVjfRECnz
hqzszBh7zGJKcV1NVXCjeUnrQnwoHKLXNKSh1qHzdUPdogKbMTEqggeyRrah
7XSyFn2osgvr1QKQn8PAoU5PHMrftPYn3ZAPxl8mnJAMWSQDq10rnWiyI8ln
a0QwZn1VKFscjUsJZHALp8HMozax/MwcSWabyW5XHhMVkfYqURG0XAB111KD
utVKH+0IU5fK2MNxNrPQNwQF7IHVNQi4BK+Rnml2FmSllU5H2p++g3eTZU9V
cgXS+fYvDBgpeh/xwdj7gVEAJBLCxNLVnSfcJVV3T51wjNqwvOeNitVRcGcz
J1M/qT2uWuCA3dELSGJBkXpLq5Cal01YPeKZ/ktoLIiTZzq2/vUB5aAC4sb0
TelRNjY+QNGJWE/F/bnXS49xkAjQ3LEQDLj9ovGq2CM1BmssLyCO1WQNaMmR
oHj1jaiJRzrsA3RXJlHnAWfBgMITjm2nuIVXhAjtSgk9+k30QvXhpKQ6GWiB
ILTjJHe71B1fEsO6Y7mKZqDRLeBXsAkQNyENNJQR11AhH83BQxn6MqK5RBGg
iTG8UBEcBf2TWaTP7Z1JdSLds8AZPV+/irJ36lndYcdnNiymlB0+5o4J1nDB
P7C7ElwyduwBFgZM+0YcUb3yKWEPXc+bxrbqAPiJdmlfqFX8qrgSL9kmBUHr
gQF2IDc4xAdIdLOy4sGRYYv0bB7ZUaNnp5WJIVQx9JO2V0iLhUMRNxXwo71h
j6O9c7/V5Vb4KfHOb2ZHDwD7Pk4wP+TenRYGDCVKKurxftIs6xVtmp9YNdH4
Z1oF64D4owXFUDDcz9QdEAezGGji9F1krbDYfwJD/DSnwPKoIjZTZhRLaPyN
PBzySYwM4quVyNJIE28wOJvH3d1BWQQG+5R6Nx/QsNUPAFOpiQvk3HPen2Up
f0F2plSJEUS5fJo5K/x6L4z9kBR3ayXxHnr7Yyx0/fnAh6vYnVRGo5gWoVRu
TmpOr0McZKaCH1EBX8f7Og+tUwVTunUMiIrHTWo/tu+MdJe0bJ8TES/PU5uS
yM087MdUM6YhUiX5zVMODthKUIVtF9KU5dxt04FMsK3yFDHQ+Eg0Pfsz/3R6
TNZl+pZMatIVqSbQC9TaZKM1c3Bo9GcDMYISJljcDdDN5x346KgBNLrdWeY0
yeLJlXKAwUgVuAbvA8Tup23H4d5S+CoB1lh+dcDF769eBOxfr3b/V+qb8T4y
kJFvJ/HKWixeRpdFmAx93NAkZvmV7i7ZX/zlsv2QowWxqTbPA9/1IldBAWR/
8+qBKZyHXRGCFVeulSWuQZMxqQUd39DfBmxQKwLQXBEcfQUXAyUQ89P7ZMMR
mDosPOjqqnWUs8/KfQjq/bFEnArppBm3DtSvt8G2qdFQdDyupY2HIPA6up2S
r5WoazAAbj6UhEIm9V11kqsFomh/Q+/WG2hyrto1fjnJ0L1P/4BpES+Tifjy
HwolEEXlL1QetJS9so1m5OKzoXGbB+cL2a9sSuNWwDhTK08mTwDPOQum/z+u
lxbslv4VA7LS9qBQWITFAa7ZJ8cqO5Cmbaw2VweFAcO6x5Br/0DAgdcQV4sW
Kd5sSUFB45Bgua6ZR8WCt4UcC44kC1H4iT6gH8RUosn3Xur7+Q965x7QKaT5
Bwf1GO0KklHFST21iwTOeT3rQ2RLfu1JDUETvq8Mtww3EtlS74QFNgJv/g8D
GgxktLGw1X5vWbt8Ce7hzW9Ell+OZD8/fTobr9f6CCLblql+9MWweSmKtuQ1
3wrDsDd5+uMeNd67vXC3KGAbbSd43FG9mCMSesXnhEwAkiK5+7RlBA+TwIRO
LvMPoK7QP0H/rTbogCmlKaQEREvgH5voyi/MyOJ9LlPWDIuiwCV+J+oWG1Vf
8tBy2Mih21DsDgt85HqFQmWYIOAbn+4WT+fooHKIChLW3+33z5pJHKcSY/YM
AkoHxV8xF7k5jg4jy2kkM8UA8dgVnsm+15zvB8ALdPlYJOAd9+Yl9tqVUy1W
10tDb4oin+ADpCxteJcVxOUZ1qpGEnzhqBC7caQilvUCYpJtaYwklBNQegil
HxBdGksEPKBjghF6FDJPjJfZt1tG2SLUhoPoJHLXYF/Dr1Wt7GUR+cCBaT0/
DF6bcZFmd1Z8E9dbMmk2/8rds1Ku2A09FQpGd+bKNTQIRWx8wyuD8HziTkCu
pB/Gy7IXMfvXcYsWV+bb6AyXLkueJ/1Df/CV7TWt8AlrxOBI/YaMAB9KUpFw
/lBTFTOUk1FJcU9QxSoAnoZ/i0NHmJ4tIVCx2fshZIjKgpsBzwLQ3uC3/kmI
nHMtwHlts0zuscmMZ/s7mTEGH2cUu0gHeKuiLCNsZLCqWVDA4OOZJdciGpWC
A8Poe4rSioNBzQ7MOE9G7NgwIKTXOsTu4YVs/HKOGdSEqqS/eUl1Mex14zf+
8HI34JF26id99PsP3VbpxwQ7m6jdS07ts+Q6yVS9RuJriDWY63LJFQso7Tlo
LVwG8hBCQHyGqS4ZuNBUWND+IpXmbBu22qs4LsK5uZx9MsR1BPfiR6Ey8Wa6
kiqiW3dWpWg5FkcgeA/gj7OSA3tUtDcu/0fTmRT6zn8Ql1wW5CCPmQGrP5wg
n650iK1qiBeo3A47ctVt3LCzhTtv0BbstQlrdH/ZGaBG7/1vCXcec/Gpa7HM
Z2Y/LC8aXSMPjZ4uJb1FVkAyaJ5sznG76aJSaoxK2w4sC718UeYBleIQnoD1
UDTGV/oQO1WknolcoLg1FGfWyCIqHgoMFOq5hcpyNGbtJWAFirgc3oeClw/t
fImqOFa/LqWcGNkNX90Yc0s2IlKym4A8QCxMl8RQwB5k5aB1WkFehAM4cDv0
RRAI9KTGX3TX6N044IEvPt6vSs3q0c3yCPk4DoriUt5vwOqq9A0GSMhkM+Dy
SXfUYlLHSYCMilOFk1yN2bjsTcaFlwd8z17ZD0xd8+rwUguEPvqxr8PAABKa
LNzRwcNw+lyLFkgqAKeXT22sBZQJHoy2pzJ2IyZb2MWp4m4IEU7d8wRkwxrm
5RL9Fpy/3P52hiRVPmMJEivk0OZF+aijXzMVeUg2ikylZkwRlXWIufy5Cafu
Kxg4y5YsL6bpsfPNUqEGqO81JxrZw2Wd8EzcGP4kBfbZ/7UhKTnD6Szhog3L
xo3xIB68btFzeeQt/I1OzfYh4TLyeqAOO5++fBBJ7z+mEoYtpVqJRvAaa9lz
+Mj2EqapqGo14O0yuHIJKUwy5RehYxKQfYgEqO5TpKQqC1GFI+iv1lu4jwby
O3TWm+kIwKNatovifNuemSygOYDJ+Cx3RKe9NoecJRbSFS6RGWfo5MO21aU4
pbJLijpmAXFcSyWdwwzeUllRr8tD0VrqX5iQGeTv61VgrKg+ZjVhNMMYoQiC
31JDB7RcRA2WM8ZUIocY6j1caGlY7RqtTrlJ6dc+J3ReAWhxyPJsyMiELI6n
+iiVYcbeYrg31t+KOsn/4VjoF7rNIONLg3Bb0JZJW1iQi8xTeF9sM0Nnm+j9
IO26Ly5BsNxNbN0gxdl56gwKxQUVD+hRpl90iTu5jbji7oWN+FK3QWlnTcjg
RU1in1BDfHjFaDmZajtuic2JOzU09c3dBtrdPfK6k0/n+bJVTXQx5gOlUZ/X
YqEhPsBDv1v44jHlyNM5jYdLFrOhcv/gVrhCZ/DQNS88stxeDyBcq82QzdUj
S67HP/CfrBFUkxeH2yc2TymAlAGzBnyc4RL13iroqJfRpd87l6KyIlJnk+1Q
8s61qFODxE8hRimV8MEfjyXh8i4qZpifiuFk/dcTM3EgIjDRmmfsDRhqo8Oz
EdQRy97Ud5FozO6E8ju4UwTYH5k96KryDr9kwDanOxM1EypFs9dW2Z+AUJMU
Yat4YjV5/lzaYN/Ou4V3EencehjpUtng58pKowBhtipRo59v6jufXL4Rehhj
cY0+bQsa6Mlewk4NbkdNGEVROMStx1+QW7pJD500QxOfitkEAS1WJaTJvkG8
r++hvv6qrL5CWstjP4HzN/I5KXu/FhQ8SiMJW2rNPqWFPqW4zmyNyrsaCA0W
jEKd4McRd+r4sGGaTtOrY9puHOPHCaBNWWR8VdrmBRkNCRll0zUkLqAHKMGY
+auFuNTzDd6XVk2aSr4FOvIk3sBjzaDsYMHZMV/d4QT1iy8ZJJ98ofYkPfT8
8oQqcErw4+SfAYusfj74ewNVxHc/LIu2A+nC6OwxJPoHWXAGvlWfuzKz0b+B
JYA/h3WY74bfeD/g3F8B4wZDScWk8fN+WOjp5xFIzRuW7Tb/f1EYgbxu17+d
j2LLZZD/Hiu7KbVkXodadW9G5orbSOWTiczMje4Ad8jIqfPUeIlx/+LC7RpX
3On8I3CWYw4xql+sbbLhVvsE/SkAwzx56EtBRRsebHo4RCqdq57f87UrDcvc
Nf3Iw7ofLNC6+xQo6HbQYBG7aWLpJqSwiBzTkDY8R0ZiasHrfecz9zCom4y+
TldIinAXFol2bowtW8gDk3LJKEkUJ4J47OIJg3vB0rU6DkqRXB8gmkJy0bwo
WsKgF9rwSbg+09neddamf3pyenfIDkMXfq/h3OadCB4QkrVumsIgaxSvYQl7
NxbvUry+UW+4fxlBsrcl/JYbO2xrDCLpx1ppKorgoXsTVgn5RIWK1x5nweP/
b4Y77rV1NpD/VpOBww95XGJZTv1bm38NIabtx9DvwBwUMSC0mN5nYQDcWZgf
LXyE3NlQClw6XbUSFqZR4QFxMUxI4+0XBYYoluNBeue8r5DjbgBAARQKZbxk
C2xf02naZ25l0ZRWAGiqTr2H8QeHPIG4tE53zybsEP8VAdnFOQbZBWsDuyNr
22/NmagP7ZcnOGlzoDMkoQPRVpzJHEtJMup3yymco5N08UGKEahc7reH58hx
Hsl4z5EnX2IPqP/oHkgaHtWf2aYW8DlW50Fh+4T8xIU3g6s21ZcwH+W09xiU
CO9mjUn9xPOF8jmeMiJhBWJIPVAXS2D/a8DRgcjtJvNLviyWeNqVWYwUW/HA
6qD5l1SQSZDiBuRaP8QMi41h2ZuUq9PlZqI8KBje1YyJCn2Ag2SI8rO/cqzI
uumqdTXhOWdtoSreDDmCYcOQTLphyK9sPm3htfQKeFw7fWxrrBo4sAbU+yIh
Gtz/uOPS6J23EtA1V73VcPRKK6xmiKNKCy4Y8V/NSDYOttl+87vwzYwWLJTH
KwgmKlgnpjNmhuwH61Ozx77Ct9XeQxXAquAd1R+fW5t19zkSYA9NDFQfYEtO
1JPBAshZKylCvmYjPccrXkithgpEJd9hBhUlqJmmwBmvOnCfQ7I/2jfraBk4
9VQjorwxjFPXw8bzXPdB+BLrb5mU8Djp1mGn2r34t3YN1L0fh/aANDib+ZCK
vdeN+17W7ECGnW3uoyLvSpR9DfmeSJConi+REgxOl1IcFmpGSL/Z+RNA7ViU
vdxQuXrzZjmQQLAmTCTRvtj4BM3d35p3Keu33g5VwDuKQ+e2Gx48K3HlfuCu
tHl0oClgN4OQVb1uV3Dg7IB8UU1g1g2B3BIpDOf3ZuccWwcg1tXktB3HS820
rSPGF/qN0ZcH5dK6jYz12p96Vvpsj/4lu42OsdrGZ5DxQcF/X7lV9W0/QPbX
2XnutlixEBwVZbMlHndPRqStilyWUuJxNRum4VlH4FyB4yI27+/ljmx5ppV6
8yD+jQ0oswLLmB7RRgWD5GV/FyH0l2T/TNc0VfvLpa2GhGb3jJLE5XZnHtw5
x3a3mMysLKj6j1N5J/Vvgd6Gi8SmspbSmHI9fhA0vAm9hHoZJr94oi+d35wh
BBKUPQQPNdDNDLlBnqgvYJqUJiMS/Ejm30YMSuUlaextqdwgh3XILEr+cS5u
+1noaOVU8LFp97hURbexLntx3uG8WzgehinH0expFLcUTwOT+0KWYmyeXlrF
y+g2XfLNe5lTU6cfy8drNYytHQ3iZj6tnb9ntpI8eETL6pAYypXCFtXRHSHE
ar4Nkv7NPAgOUxMSPxKOXqlnn3vqltyMDUmJufl9eVBvP66Iw0TgS2Dr2S1B
UTpUAybwbosbqJmLp1Nw/iZ0lSco3lDcc5kJZ7kn4x6LYE2UEJ7CeEGsMdKY
IA8cQ8hWW+sM6gYpqFAYKfBeWpmRdeJvceNPo1KrU/YEY6HVVR9UUSCdr1hV
qPuVmnjfZac8fN9M5zl/SgO8a4RcxdQk9UD9QYNgxv58mwLXC0O9DdrXZZEG
eStDg7TOYmDeb1AcSh7D4Gl9D3GfXOuB8vF7H3UWBjqODKuiOO8VxyCgvwqc
zARz2P8Gx19iau5oiB0RSqpllQv3jsCZwbq6dHPew8BUp/54VmIccexB9PLX
0zf8qJJ5tIsS3388a7fU8EN5gmN+RlIJWvrEgtKY3kc3DVF0NcKLZMJTJAzY
szp+dzTY63rgrGjuczaXfe/fhEQHlk7MgksHLFucoKkRWa5wdOHbuR+9OYV/
CYvbnX7O6l2EbgFXubMk+yqwX9/jJD8RvL0g5coHihC+Eb0SXE5tLr4MJpdk
Ycsn7nSSne9AAQHEG70MEiEAFsyB0hlqjB221KOR28MD8VI+DHKc2hwBhk4R
NyKkQbeJAjLrG9rLNWHvMRR+VhyK7PG4Hdi8X3AR/fyTWSm3JLsTpC+xpT8Q
DcFsETmyOrK7BdauiLVDjv4oAFZxERMqIeLaL26rmFHxjVSRQMWOsCoD6qaz
l/5p+sSqGRjbaZ7PPnrt5OOqlq9AbIPC2l3HPDjgV7mP5dKbyc46tM7OKuFy
u4mtp1lSKku86smNjuF9aX2mjK0w41LuIfpvmH5f2V6L7y+fY6QH75sLaZvL
XfZ+PKtEwZx4zQiNZ/qtSIsFuH3cDGO8l6oyWdX/YtG/cwA5SwRmFTbQEUxf
rq7AdnO4mrgHMZBgoZCFyrjd0kM7Y/bg0Iz4y5y99K5Sd/i+UjucZmkxCOE+
h+xrvsA+f3nRYmkl8/fjFtoINjvy5HxKjZu8GDCPBBNCKR91AOZLzMsEa25m
R9I4U4ATqFfb88lnnHVLn7fdPgNfq/8d/+h+HCJl8hlEUnrG7gXJZWh1ctC0
HAIW3gQiIwMwM+6asMxw4RCQICA/+HWGmnF3RhsSLQTRLrTJVdqtQ9FOxvhm
F96VoshvyBZvv0gcN16I8ESWC3JLozyel62q8fAWBqCMbpVv8qyFIwLCl0z5
KNgOBHRu9+z78ra69lofHyKGahU7RY+Jf/1qJgt9NXbsCkZ0ziHuVKkKYMMS
eyKjg7+49MQsSIuA/D3D/6Fdsruja1Gzqc8XkGTohfBXqB8yluaQ4dCQCBwR
F+Kpd14Uq9UiKNdr4t5kkLStVYr8jUxEIR9+kLEatGJ+1BjXdD0F1She+gzl
VUFAw2gPrYmn2GU227sLw98RyD0NEN0TC9tgELZ3gOyTGsOLAvXXVjs9cWpe
tyzknOrUh4WNYl6bhdtNv55n2pViFqdy+JmBoKtCSbU44A8k8G+p/F26gE2/
udgc+BnM1PwaSKxV0SWnV7iiGpNN9ODw5zKove1vhetpEnWToIWLV50hSFZK
nfDz5SNPgi3M6LVND8NXrDh0t9sb65Q2GZjCE+HB52QJft4gWBGf5Yf3sJN2
k3HSeFQidI+KCvLAs6J+Yoh4f0h6R2fqpNIjRpEOcIU+bt4ZtUMwO2TBIq+u
9ZyHqozoyL+CzwMeoZePLmOuW0NyAOEWMdJDoF/X63/yDj4d/21GZ4m2dNFX
3mvy9AGByujVS4xD0n3z8MT1k/0IMDoFoE0I7KdwAbKpMpHvOjEM4U2sgUTl
TAIpD45xhsCAtKI7oW+szOI2vfxim9QSm3xyez8SyemJ+jTA2ohjI7KuUDLO
vn9l8zjoI/3flFyGIMQQSDLkaiLDDhdEdtqcXd7TiVD9lW7l0WpYXAQCnOnK
DqIYFACi8WLqcr6s3z+ABlCZLIbZP2PIChnz+GLfelqgZaSqQeCO6VgHyslU
HCK8g7wt1JXWrDryaJTtI9uCVpHmL8EjKw3qsB8krqUBWoqmydXdzihtKzZ2
6Zv4iYw3AjD2wJnKlGnZtwAV3CGXMxcHYM1Y75AVj4fkHxpsbE1D75+bY5E3
7wdC9e37wJkkK2pjhL0Ra5VrTwjE/6JA0sgt1vdGhkgPcpy9PwS54YVr6THZ
5CzRRMnHvd7R0UDBRRdVrXot+NPM3ce68fehI9ZOVGnWZf3rTEb2kURX31kz
oCivIbQfdv5JaE66uZsZVV4unChEPHo2tBY1aCcG1ZsXDBCY3cYre8cD/lD9
d8tRCmDuFwBcSAcew+h7K7JlMy26o7Ft7UqiIvzp7RBm+UxUS5rVf8JkjKqS
aCDOgyeTcthpaffnsYrCW58oRpkFngjSXDBFGUFwNTzWX4a6uQGFECk7PzJF
eSuhUzkU1b994fn1PDVY32pGETqcHQZ42FcstER/7UZMm+orcp9szPpzuUpU
4+m6GEB8JvG8rcs4WQIHBm1voHBEeAmNsN4WHI4+6/Vv7ZHIDixIux1CFkc9
nHxjCv0z2Kn7gDoHCR2iHrmcg/amHYghArlg08jY14WIthPVTV75KVt/aMn/
OuJ7WwkBgx/G63F/+8MN7RBMkFS2sWpiVSP4Skg4+D2u2mc3bTo5YRakIpIV
ziFpvBKs4QnXPozoCVo8ZrI2ik6S1sGHfDCvSSQj5iw1N3uqBjvpqG8YG/Lw
EcRKLzbtE7bfgWAwGdGigFlqYfgYAG4B4ADFy8serqMw4g6au4VWj6gKWVtF
ySKMKRITFt+jJrZkNAAGj2VIe4+025Q68+19YxttnpQJFUYqgFOJjFex+BH9
zzPQvKX37hy+y4T2XSVpxqBpyivwpM0MQydrk82E/w91e8YywVtYL+EY79OX
SaieLpamlN6mz0UWYErJ3B4PF/UINRqpOpO3BPwCW5lZ1ykdCphlwzAghSbb
Rb85KBqGcCDeTk6l+VUIEEVt/dkLF/9fXIpe97b2iuOeGk3/y4YC9mYPdvvG
xwHjE/ZbCt3iSc7M+2xalpybaoCUNcPsH9L0KSP2mtRsNadkXsT4qxOD+9gW
tV9xydnE2MWlxCjjGIGagUwAJs18ZVaCN1RcYv1G12aQTCo4R/K6w39ca/oE
nATGjmXh/Hb2a0KoaVL/ZKTBRWv2cjnoiI97NbofhmfWkuYw7XgmxpFjRsh6
Yp5lXPWdTqPqDKJCvbV36xe2UtPqNMQjr1xkdPgsNQqT1UYdSMeZZlX5Vh+n
NcuUE03GqR3gNOhXMFx93gr+EH7iUFAuNw/OsJDNAgw8hGauPssZTybVQkDe
6VA+QQv/Mlryu4u+pDR9kn5bM6kQWVjbpwoTnlCgrX07t+lJye4yWXY9hXZS
e7uh6WHIaEtcAa4Mb2zBEuRGiYaZ/WT041wXlvUZZacef9egKGIXytLxnQf3
XJJQroTI5p9KDu3mqXIAKKqNUefOuUeSrBplFvo7eXRAnH0a1AB48gPsMvPY
dOJrvI/RwI0LyyROlhVG6FkwQOHZOgeKdGUp9W8nllbFl9AKLy/1VkV0trkp
ayCFOcMcpCqk38Eg/54sDQR2rP+wZhQ4Q14oNrg6fhumhCEX5oaBOqCCCgkA
K+ZRNDBa5YM/UtoWgVn7P9u8Zko7t1002xc3lv9C5O3VTx8Vr/dxuBez36cu
TuqXsmFM7IN4Jhz6M6LrOrVkV9yVGdaN9wZYgWf8ILdm+/o99JdN2btQGeXU
JHIrgghKjo3ilW3RJ2qa0kVjpqtWv4g1KautFv5AmYNN0n6RJOu5XfNE9xlh
nYbTlNo4NAxavsq93WwCKe2+yLmR6gqKXnHcWBJNGjjZP6A6iah/g+OpOeG2
RwruzzCvuE5YTnjVSTEHyHF0vrr7vub3n0HJ7ym8FZ5LEeGx0dsPWdTzExA7
zhOnoToyXHmAtOc2ZyGgcVIVE9FudS8v3sX9rRlWN0srGgv0Jd0bIIYtS8mD
JFNJ9Z4oSFBMww4/LMkOT3VBWc914eRdstYeQhInsOU/JHhiOLH/h9J5C6BR
llVBaQamPu1PRWyy9b6xrOv3w+P8ILCDlER/iyKkNoyPhk8DyMplcEq7D2Dz
cNav8st636mjhOxnJAseYRym0GQhdF22YDp6jd7o0SUp5hYyYQSJa4HL6jTO
I9RtVug67AXgy/lSuWW+RZO64vylM+yhXDgrnE3br1sKpRRalUEotIzeXK4T
TGEP/74LUW4ckZ1KbdTJfkieNfKlXq7v0ZXAB35axaMVKBwGIXAoM8h8/0a2
GQpuKliG6D9OOofkfSl95SfUndgdxmLdT0oqwMls7SfjbVF5/mbjl6Uzx15J
gPqNlnxZXnVRoJO+ZMwIvMqn2VAda8rwe9SStDQVCUOR1yO5t3HROPDK8GvU
PNvFNFL+0x5bp46vSlhC+gXfFkO1aW6/4SGM+ZEzOkXUSkEd+KSs9ouvotVY
3Xt/GFZ3OgB67NyYB0YjVVPYkQnNC8/QtZAiBt5BWOckV1TyA5k0gG5Z01xl
eKS+mDOfX2ZDUOxSMdnrBHWIjVeU/fVfQUaQGn2+vjpdOh0oqlm7Tdlsvik+
+jGAdakhZJQv76qT/QkoyOavkyzxwNcbVW6qM2Yka8RTxeVPwJX2tRsS+0es
0a+H4MkFLmGTmoCE6En0awoVbhC5RGO27DSybSH99MtWD4wgyobSwrKghKgJ
YGokF6PK+EKWnyK392/NtkOMLpdJEhVkfYFD3cQ6eVolcTPjO9ABXxDjzg7S
dFnKIdZiapMu51SmjcS757oymXNFBBaXNDNRddeqto31kuLXMO5XKG+ML6nR
ledLc2xLQjiNYAmxOeAHCudSmx13luDdJhxiP+En72ArnI+HRIMAsh6tfk+0
xoRTiAM5whMx/X5quEy7BrUH32NckjBrJjjgQy5rzgZdG7XiiAte2LILGNRz
oAjDeXJs5RVCzS/U3c/jbfvqO0ytu1NVfm2o5cbvWMoFeNgzz7TdkMw1iYdD
HJZ+CMikZl776RtHHdzDqIaUfcU30bBbGzoTMbLdQtkQjbApmluVaGbfTQFm
DIT2LWTL0uMM6myj0J9q6RPtMQmoXQ942QAKjnXDxtXt+MLLgk6bq7jvUdyS
vCDHt2DEt0o5fWidJE+M2/LRaW7XHmZa1MczeBJ5zUc7yaFDLgS74pu3rqCc
Fd9gwPl1XdG0r5IAtM2blPhMFvD3P76FstOFL8e3KFexif3mXZBurtx4mw6R
zbbohG0ZNd7EcAdVifwyo6Cm08XmnLJfWrRAW1Aor2VyGJpaQjK0s6f6tx29
3iTJoXPYHDGAswndH5WyhCk3/qZhgeToNkEpK5phoDg3sckDzI8UhlwfYu0f
XnK3g2qsb5Ubx5GvUp/7fi7GUzISB0LWygLNkWrvpwpGoZr3XXlWCrIKXSr2
Tlg7NzFOJt+dMCTCGk3DuSPPjkKeTa6+bYgLue9EG/DKHI0qXYilOOhlrNDJ
k60qUMARioSwa8R2MgDFkhV7d8fGMdXfAfkqqHaDd8RaMbKg+8P+8S18lePW
cccTvXtkGwXrSZ0QBT4aZOhauddEgA9P8iRbiz6BoZR10Vicap2BS0wqsxpb
Xu2Avi4zgNFrL+xwEXlaoVVO/J/Su2s8s0/nwMMT8UqTOvwwmyxXTfCjJ4qP
5J5f5nedyv5alx886oR14FgLj01ySefL546tI2xRL2s7BHVz5jXlRspeoSvy
RVt7mRhv2uqQkpGF/2GReXjmyosEqclhD8LwyyfqquZT/vDLiEgXzQsUlTFZ
6Ti5MXJ0BORV/KE2CA7t7BbpDsY1PgkhMUJcLeN0rTaoCMq6Eb985Rc9AKwM
rt2mBhCtBiRjUq0yXRfBHS1JWuvP7tQppsqPGx/FmEDvpLU95nqWxfEvK+I5
F9yYpBNbrVDShlB5EpTZFD2loDM9ZdBiq8aRw3/8OnXIaihxi/nww0TtT+gU
6p4nVn6TRoD5g7ENcn7pcUkhTS/MYs6l15Clm1ncT6W+exyoRNq3GdngSZ5m
NRX2M/SyDsmEHiE5BYbU1arRUAhtIhCKe1VHyJlWMEhXdquBTLbSvbk7vReN
Aqn01gVCIXXD05NL8ro+OKKwVQfICx+5DKcgtqrSgPSjFjMSCxjSxQX5fudO
y/x7/M9XVClRSKclxrNezhWBxnhIAV5piLtE91HoO7BP541Hif8AC+Z9WVl+
Z2XYEl4xj/ihARJG5/UHbOftfobscdZ80yCv8H53KXV3FSF+AEA5nYRRqI5a
x5qSZJEI3rhlLfT1Pttg0uI4qTxXiaVQX4QuYmzB2TRgL3WD9JvtBnwnzppR
7RwOXkUtVfJ9MMD5NCVGTdSQJR9pOdvEbp63ORRjlv0rsPdZqnNltHxXL0AE
n8m+8GBe8BiXKUKViWp8fxOzi0aN3gJpUs6HUeA1I/Itv/bC0ffHSwIR23pO
pdZU/7zNpNngwMup233B8gTdc9Ybqj29+9Ysfi0r7e5GZT5LClGfQfuxikjL
p+qpMIrSWhRS82byk5oRVb8sTKk6xB6WPIu5FQeJ8tT3dpG7rQSJ2r7M/tui
scZ7MaZQJ0o5pJK9eqm6R1AG078UplCtCHIfh9ms4Zmqfb4KqkcC5R6cADwo
Ei1VyD7yIbco+Ft4vQqg8Qvu4tH4lBmtdgJzkHDDXcVvsG4KmTm8D0oBN9EX
Jc12gJfCyn5l9Zh69ChB2fxoLzUFhLRAKIBFNpUTgnvZCNxYTu4HxP7j3FCW
5c+HAUwzqt8IOX72B290cLvbEDj0gAr2dfW/iAVPjDnigPB/e0nLKmDXMOL0
owIlMrRAq4Tzft84iEROSbfsrCY4OPRw47QvUa2KaPAhd3eKN2HjAfTMJAZq
BZd6bzd9dJwsilnutKbw0N0Q+FT6Z61VK/70gPwkEHoOXx+YfhvWlLiuT/MC
ompSbUR5Gvt4XaFODJS8/rp7b8uF2rCeFBUES/3+MBRqfQY/gD2/UHEAfU8d
Y5Wi79mlH4k9nKHQp4l/JmUeiR79KyiWe2Yhk4LcDnqjSZTNtvobsiDkASTB
eWwg9qoGZGYkCsUXES+x32uSWHwr/7aDQXkZ7CUFqhO8eT2HuSeOUgANzW0Y
fms4bBql70YOa7kqN6wp8Hm3pUVG2ByLL76S3iVz7WPCVhGPlYfgi/fKaqXk
yMize/hm0AaRXT234YSQU9yYATv6rSJ1/Hd7cvK7D4Ai9uaNO18ufddKyJNM
u4qzC9WlWJcCXsJYAPFarwjIxDDLNmtgr8Aq7IWCqnGFo0W6SJozgFDtcj7C
M7aYYtNAt/3WlECQSKIPmwqjHePvHHOf2vWCPsqZ++CZiHyRATgQHfXpZR6T
06iKyDAWUPimpQQcF6jRCAcMrx9XQUo/lrtxYmYIa4JS5xy+N5pjJD4J63jL
6mZ/v3Fs/RQAM+q2vQVQlIWT6hb5HgZHPdi9W90oPrzd0eYcG+5T/CPYhtom
dsj2w4uMcPajl2NDiQ4BYMwo8ewZFj/PvH8NC8Y84gJAgD5D6jsm+iXsZ0U2
ZGqDuvkpcXRJr4RXD/LTWDv/yCvFO6e2v8S9I6Ri+sLFc1Il5ooCKCjGPFmZ
1REI/MhnjC1gnAo4YBRGZmcDBeqnaUdD9uKvIyAb6SLo9ZLsGEqy0AjVxKbr
hkXRf+MlMi8xklldvQnvf+8YfhtnQyHozn02b/LVCvn04JLgSCmEl7duYr+z
CgjjuRHN4ORyG7RQAWc0ALEI6AUcRRFa4w/AUc8J2sRn6/8qY8GfcRAwBVkf
K+WyJlPYuLV1xPfVxwWtAjrPYFwIa+fIcYDrWBVvZAS7EwKG79W+etL5Dc7T
VG0ZuPKlX7q3vWwRfDrR/uVUOIHBuOq1WL7utUtLSy+EoVnL7nLLysAXAMMz
TYO1c6wdtwIqBeXzumA9ReGyuaHkvRFRnz1VK8Qz895F4O1M2Bh5pQBCn952
pRHtieHWmktSuBRwMYXVuCMJI8pjIErua0Ysqm07YBiAPfvarTgXXtNCa+Gw
zu8+B4gEIBX+Bf4muPt3ivcs1pbTSWiDC79kk9fEtGdvVMaFm38KCmobsfuT
bNZExxFPo1NHaCi6jstdjpbxDV+ZF4PK4VWNNGjMXvSjjcxMjDOobFDeekjl
GUwDUk573rj6nIQbpDwzqraUAOu6gLA/kp5sWUo2nUBCmBVqNnEMg+Bftdwl
eiQS9F2Q3y1MmROQCpCBahu0sAUGvTTJGiuOelKqiV80KUitvZ4c+jD+n/y6
yjJdnpI8iDBp+AXoQMBbcJJpVwvIN5TE559mLL/L4OoASuTLVFQcxtjcSts5
zTRxiVf+UzGrEb9i4q2/hMQ/iokaPgpfapAlA+QGqfSIdHtHvEWKTKEWYuiF
YwGASA8vus8vQdCmCyqH+zkbX8qMDSLw9UnYvdE9yoYM9MSzjuBmGRyt+lXV
Cn8WrCpOjt7QIGoY78iHFEl/gp5A7upt//7KgJvsg1U9GFxxOC5lVXGYihTf
UeK4Pu1H6PXOGrKk2i/WjiQAJI3PJKyrg7vF79x1zNynIQ4/kiuJoKpAFTmx
Ms9hJMuG1WG00h2cionwuc72Lg3+PsTFQOQGV7zlRkkhqNMxejs99fSJhNzz
2Ds+cUkVcHShuf9ddK4BI4SmxCHIkTqwpeWzkNhA+lLRhYY6pRfPB2rIHPEr
nniw7NdK78SwWJkmkuPaGjyJPIxtohN3gtlsGsg4EcV9Ok7VD/G2h2XR+FWw
ilTZBUIrQDfGin6oKMvKCnBpX8aATmL+0XpqCyzW4U6GQ4BEX0HcL2kKM1RB
sSY7VSmQL0YJtmNUV4QcdNCYQ9hUARWE3uYWpyU1hIiR3igmWJr4u2mVDbVh
2a/oWe/gBfIlw4sDmBITEPmaLtVdkK9t0eN9OnFeRIyAcV11vWQvOp0Pyt87
9ux7dAufDFnCHmHs2caOYsgZuGVEnIJhK9pCc0J01ZZeAa22Wee/fNP6tU6v
C6bVAUdffkqdfYFlWlJ7rswEy/PK2udym0oA1Czfh+oQmFByb63cHLLvnlWv
//fxJnzWOv2s3Hb564IvdzRfLzBQlKrxYtEIdvx21PZH0SOtyKuwLSotdtcY
AhY7PVyjZog8++1Lx9FSX5Vd+rZNzI3qoXEJwCtsiw0uK0cLOsIQ9IxC51uY
R1SSjY413LmdDyxFIWy+Yb1+AWrHTbGCAEnuXc1cTXzF7eJ+6rzziKLUsnP3
82R3GXeT0L9OJuPknVMEPiZ3vu1Nq4mstTUdXbdiT8Yk+wxozHYFFNOkH/FS
VAcNL34wMdW5RqwVpDtgUzofXcmxzh8HbuKCrOZN5LlxSrie35k/7XhfIY06
X+9bKH0e1a+pZscM4wqOqa1BAxqCHfBSAYjhiyvgMgEZvXOaqvCEeJ2f801B
mrePr49imdpZL5oXI6bmqlrstnbmeqkWqBabQm8U65AFpbyRqvYp5HYDvaHD
XfyCsBGQuN1lbjjJsqIzcnDgbz3v4IS2XTWECAJV20I+OcjRxQ8GBd5OUJXR
oqrwUcTREdkwWZ2ATH08n4fcP2DYyS/CDgAIQ4rJapHcHGE+MxcVdBUj0G9X
U5ZaqLXsSVh4AiyeLAkLUKzOI2T/KOlQXJo67SWocfwQjXo+bV827k76FE7w
wDtjeNwJ5eHSjk1g1X8yBW9aDAe8mQkqpmOi8HQW7cpNbXO+KmWxC/HqkZVi
DoFRLqty7zIahssl3gSaDOYx92zpOGLD9AKmvVQsB2nSkkkMfVd8xqBNotu7
HX3snrmz6/HwgIftpFZ2LfhWqxx+8n3DBNcDPoRanjxz/8RBfbQXGZ+5CcXl
0IKiMxctMqnVOQOexOiDKwSKi6bFNOgHpxkRtMtR7U8dP9BdHEcNziP1Qwqj
nAzJPznBIbkyH/lS6dJXSEiH823wfDmJlJBVLzBf5WGcEm/eYDvAf6uqcPIn
G5amnnroB1JQTQXNDqz0p08HVDS75R5XMCtYh4u8zshxWV5Q4JlJBx5TC2ni
jJwxdhWouBXhqdPZHovtHutAJHSZOxU6RUx24gxliAKGGehntBUo4jUeLEfn
tXQHXyXkFASoYep3qWz76ihE+2KkAaKvGJ5qfp8ANc0c/s3ZlifvvNaZNWPf
EiKpklpSvSaeKKS7KvcWtXOkLjuOuL3ZV6UEJy3yX3V7hTpjvGLn1anu1oHN
T/faR8rCdtapYtMvjReaVQynURur0X5rCjRaogt5ma/zrHyceb2eidoY7T7V
dX41A5pTkqeQSTVBQ4PvYvX1s/Tx00UArOtizI6tI05ALCxREihbWP0aRFFO
LYD6T23BWqmB+NtKNaXnmaR0cAQUKkEroKMWobqq6q+kB7PFzYDWQ8RjpgCw
oMCW2ZyFX+bxk1k5zn0kJk2IYxBUJd358CjblKbpO2/r3+EK4jka+1d/fij5
qkp80Qo2DclqHQTcPTYB4560tsnOI1EhuS3kXS0HEuZBYMYf3l4Pkz74gQv+
w/CfdVxv/vywd35X/kN72d8O7BJaFlkazBO9d8CjOd9FLOczBeNVxuqkAcQe
aNFG18X5u/izqc71dEhbVF57x9ZHKS2ngQmo+Dt7KgKWiZ+m+/mDyIzenEdI
DTJtozsNyrqu+hE4CyTPxLrlulG1Nw9QmcXtdhiodqc05R+ytfYgLhNkAZ4k
KafbCQkqAqMhjluKz7pkIINv12eu1PCtH3HDXt2oiZvY4Nj6d3PK5AYpC/Hf
5l/Ze7diFgXpYp+uxXVlw40iz+kLoC8w7DYN/VcSOsweznWaywacdKe5OKpa
l/baycAwyaEeKd0a3KL508NmmvuWm8VWV8FEBUQfaIqWRPgCmKKurWH+X02j
dBkseiUtHsna5rdMM+qDmdzWoIDNf6DkyxwzXJwhg8/2NdDOixd+IGtxBPB8
68ekl1lItnOaSTvchtk6D0YOa2dsaqydc3Pz2abup0VardNlYgKVCNw2Ft3Y
lJW5pytJQyTTL/gdCz2+Ojksv00y4qc59Qw+v1AVePGIwbeylrTo14BD1+sl
QOspxTDRienq68tPqe3TYdMifA4TiMjCqvRLbyThsx3fFXe6S2O4Vgcz/Vz4
fzml3sKEbtWWySJVovA9xdMGpXlruGc9w3r3dVFkYt7CtjctE0LfvxPb0biY
RwLEWNyvTGqyCzEu9pZ4Z0gE7zMLK683II6OYkJsbz8q9UWggpLp/Ik67FH4
qEGFqRvxTPXS0ukEoYwSLjnVLMOOwCQchIvSM7GjxLSJ7SWw7keG6ukN1KEs
dNYz3gRT8UJk+XGuP08Kb4rLlwNaj+jhOO+oxdM/EJVH+GIjsb3SsR1fva7Z
1mPXPNZEZmd+XlG1mX8AfdzlrpVxGUXN0AHuiytOzUIk3tB+2iFixGHiwwgh
R3ixKvnfNCGjM2uqAATzLaNjAKEU8Pi983Nw86QWVEYYVtj48OLcDhF4qU9h
AQakx0NinThmB0k8CSanBU8X4JoE/aQed51C5SHAlsHQ4Q0OxD0oUGmMx4m4
fu+ozhcTLYrcV4shRYSy4oUpZNCtc38oU/I70ho/+i99UOVwaglVxLJmXg/d
mDeDNHjwGGQwoS7zOZZNEYtDj82DPRerjqHs/FlBtP1nNgP/4YiQXcwQ1uMU
oy4kDbkfViAysLfZ1y5qFCPSkt8bmpHPH6MuCkZDWcyRo+LnOZUGpeNSJ6Gs
otibLLIEcCKMRuoy54t05I9uL6jh/OAksfZfiRx0hoUpaLzKUXcmJgg9IPWy
far/+ukW7qyxEfOEiWT4jnz/jqghYcc8j1zGR/+rJLmMG55r/uv09/PejWHp
PfESpxr3Lcno8VnUi0Tp6pHMvQjH5DFDamoBk/kjQtwprJABKObVKTpHucnx
Or4uwGDGjbDQ9iQnvKPJLYnK6YNYsa7WBl/ar1J7cxHcnHPeUlfNJHLenW4B
NDsfPALMQR/VaV5otlyAUynDYwlRr7h6tXYVi9OmI+fhWNp0IGnF5uDVq4Br
GKM44CStqXkQHbUoyL/WkbngtOz/ZllpedsCIyxRhA7cjuu0QQfH5Z3zcVJf
rikihhD6NFTyyjVv+sYyrKe7L9z9OEtSYMHA2hLbLEVqDlkJuccEDNB75Sgh
Dg8Hkq7OMBSttjX4bEa8M67DYkRIXm5lYRawORbW8+LGsMoxCyiLgRv0NANa
bZzrjBa6B2KJNNsb4Kcz779NCg245+mLgtGnWxqOu/9yWdWqeFFQLywV+rT2
EKNV8tfQVNfz5iGi5Inf4QVmofIZVikUks7MsupwP/lAAr6e2IBzeKsu/UYy
NFj++HTgLu6hv/7NFKP0cpDLZMX9fP/i7HWTjiKurdPYscVbr6GNWLxPN0ly
okJoYJSEwr7/M2oyWXZQ2A17xTxZC0tUdnBIkJGC81Hp7fJFTpuZzlmBWOxL
GhEwVpY2nYsXs/t50f+c76l85+kITC8yausKfYgSBpW6pKMqsrya1XyAt8PZ
dyDPPKV4qLSv8IKOoH0XjiDiDtt7fQIZIkQwwNWGiOOyhBQTfwj2ZrXPg8jg
mIbOOXTa8RI0fPaBHmtAw2EZ9uBVlpQo/u0RWS/VLsw1Lt6AI7c0itX0f22t
8t5ROKDxVZqP/eK3kHbb0eW0eldf1XxC50yZ4x2w23Cm/BaR2jkUCz2d9t2c
U3N6m27YhOqro5HR4A9JcpKDE0fBLJ/wRSx7l/dxcVDcJdsiDxwZRevTnD17
5dlG7RudEhFxqaHtYl7OiVQJ9pLl9grAsXZb7myuYE795DSL75VRBrm0vX4L
K05l3kcTBBBri+ypStAUG9bK+XHIY8WRZN/S+3JahwfWwv0jS5IP/jNcadY1
zEzzMsuSJl0j7O9N7G6v+WU1PjFqR/Y78VBsdh75f71BKJKqO5T9O5Biy+37
VlweslLhqgzABuh+BMFiFSQnwBVQFdEp6lPjTzxnDmr/KxJxCA0e6L2YdMWp
OZ1c+FQwKS+z4pJ8Kl3BS+h8CZB+NUgbbxcDhZZP27+lBLwSvyoOGyyXWtL3
WwItFDWlvl9Lwe2Tq8YL6ccOcO7VN7yhuWrllA2Ox6BWOf3uVxR20fr2ZR3I
piG5QmCk24MrhYsoJRXPhYfzm+M65PQHfwdhdFISXafCcKCDWncO5pr/2j1H
IIm/xYgeeMqzJ85oKizsqnMf2VuGnqHcNK8qUlrbEBrSEVvnB5cyuts3KD6b
b95SMqK1cSpO9KnQ4608j3VzsZJYufS7bvVok93vyL9w9MNpKKgyb0Jf1pWa
JVMATVRwbjDDoKspNXlydhiL7rAg+3e9+gaUxwHv/8oHXTuH+hBN+8f2GmxO
pCMoMgfEkGingxyv0MACo1qLplrktI8Pl1E0Whr0AQ34lsZqmGqce3bTz4k9
SKuKk1A0psv4Pisv26StBKaMPu7NbBaTzdJIfsK93zkQXmBBcUiHfxpiz+hd
G9wzPru6t8P0IPnx0pf+Y/GOMw0czK75MvZNPVrsazqHtFsYVzX4FTfNyMof
+85BlZa9Nz7jNdLxYAA2YhN6Ydv+V2G0E84QdIAtxQm/SW+TQD9FawBsT4R8
ddyTW05MwhPZac5GWONfCZV2SCQk8NK7eivOAaXR5ocwpRoC+u7FBTCA51/E
OT2L9fii7clY6TSek/fyX3sQyRDVRtGKTjSiMP67aG7QM2qgIppbAOmQ9G3D
BaNFdszTSG5H8b2zKjBG+/UKfoQvGRoBgJBHkCaoX4Ka6pQIvuiAYt9w3+0o
q+i0+RywEJ5agazZsYcLNdmF843bGOOlfZOtcv67KJr7zmg7AdrHlIcPdv52
lbeZQIyeNGp57BZcv9xnC8vNPuh0+ZC1145gRAybLyxbDU9Fv/qJZHtOnu8F
PcHVfvWpA3bN4uJcrfr3IN1E+uns2y+Vv1HKbPUYJZZ3mpA7N+xwLxq9wDpR
T3uK1D1WA9D261Y1WOBrxxbOqT6bjaQ0K23HBfsQWjUYmP+i6nQ9XXfzAO+Z
4WnFgkCabDaVx5NJMkuQYTbEnRL6LV8D35+WDtbeWGTUqKJjhFS273ls2ZIq
F2Z2cctEy1VSgZoy1gXWv2w9N9Wk3ECABILSfMw7wsk0qGaEUvkYzb78S6tx
XKOkCqNHjZuyIe8sAHvERK4p4gykj6hYFNYhJynux28Itzt1e0uPa3DjTyVA
Axd31FbVH8R/TdKvXTrRbD1Vu7tpG5P8rPDSuCC5080xs4nKTxo+EcBEIzSL
1jB3XGxP6A7C3zMgXB0x0WrNpzhe0kOtPoZNLuitRj+aNZHS2B01oqCI4T5k
VxTh0E8nlhjcXx/Nm5+iLp5+DcxfdO0xGWyY+C9KMJR/q8a+82NDN7zwEgtf
8eTfXPFpPeIGN8LnSID+t0Zd0gaACIGiTrMBtZMXXbdPAjIuhe2L7sUkWm5f
pRP22K8RJsblM2gaeFO364soRSwh3wbksGIaObszRHbyzBiZJehYMMJX0mz/
pr3zySVmgmM0ujndzKKN3LCRkgNLBYwmn39+rC8/yGLWQ6m6cQ4HLLnwB9cW
HUfmVxtiCGyvplRR8igw811yqp8Ha5XNGgVZZ5Ea5xXRFIM6PEW5LqsZ6LGQ
5VmjvYzCuOxU3GoqRt5XKG3HD1xmPLhhxYJdSV7K2F+hbavMwEP6Jtreb5Z2
XGDR2+T54gLk+T4B7o4g/ZLkn54uSDiH91tV+a230YDFJ8Ldbxq+907YcQnA
89E2esvUMEp2V8/kxPZ5oa9Y/yRwlPWk/93xM6V6ZCPqW7K1pc7Ds1oKSiQl
zvPOsMPHoV4BiCmbyv2gmfkxtf6VAk2oBhaRi3v8hW+CyQ6CCZCITtMMEq5y
MWr4q3dZIP0nZporQvrzgSRd2jDz9Q14cfBxxz8sAZICZyNkKhiUBZo3rdLB
lcBJh2ZhbmVIlah6BTz2J7yFaYvqcWLRVn7HdJdyZksBvD7XDdfG1oSdlgZ2
bd1QBstBPHDsZYpx6Wf2is/j4xlpofZtffgOx7gOKqSL+6y4oyXrBwLUu0d5
6zjjl0mpR7vbhSQ7wKpFnFjuzhTxIYIyPfPNQmhgR/cmWl+MMYV915C7NMLp
yRqRQ6IlScCFxWFKcM8gPy8Dhzjy4S0F+ssXvTVJdSBad5Mtel7TCpG+fJoZ
gYjbNouUK56E39WWBKKAwTeLoo1TFGCOOsPKCcrh35ADBWH3phacwmTFtPEg
DGaLCuFVqwxC3g7NnJR+H4xvsLmK0F3Uj5vXz026uD//2RIkqkemc1cRhuY7
nMwbKK1HpWgCETkh1q6pHso90ylsYXhzHVqQB+QM2Y3Iy8BTHecYiMn13Utt
lRlcmjn/216Sl84grZzLZzy5RfGvLZGYdnDxed/caBSWvyEyFZP0O5bMK3j6
iXNSeFq5sd2csXVToUAKzPhRuRrctCJgq1SpFzjicDTuSPHF8ihj1xbsMV/l
8AHP4njD0nJcGZzNQDnnUBNEfp3jlG0kKY4Wbqr+8LFQMQ9I0R1tp7hCGYT0
sre0FNDG5iE5O5Tm2Xn1dCVg3HzIAVOuvHHmTZY4fEExQJh/1Js8kDe7sEoi
Zd8F+JyUi3at3KhLNpfIRZSlbJo8m5WF5B7IeidiS8pp1kXXmp+wnx/3yfBu
82aSly4VUgqgLWJFPueQ5lCKqmiG07hOZjG+a6AkX0Ag5vERdfcCcltJ7xCH
qOTwj0PdbsElXOBhw4TXwUtoYSA//fji7yKsvV+9a76bQD6qCt+MjL1RGyIf
094fVDeRZT9UnKVETC7DU70//ZBSV2qXw/dHS6yXWl51VHoX2sJD4h67XOdN
ha+aDcNxYvPM09O8oDpYj0Tjc6SwlHVR3wahXyZq0cbvjuAjqIgvQOm0Qq85
c0q8H19vJruWcZI1H/8B430wQxCfRIPyj7BiVWQ+DPHz67vbHK2w7M/cSyDT
eoE/H51XZ7ncD0SUfjnxto3JiSb6B6WXSw5gBh0t9+ZVXpqG9gGKf9HMmVlx
wabfGmzVv5eYjY56/gj/UATu8SbSpK6JWDDl4Vn5xWEUxQAcjscKcB085N/D
t+wqyMuZN4qBNu4citcCRptu/uGwIzbdtFuZwub28FL6AEHMMzmjGmKdPjMy
I7DWcoydZ53S/ZThP29BNflmSOZO7m3STiJr3NxLuvl9//4Dsdxr0RgafWQ4
cbRC06Tzemg3xrdRGyRSLjzM/4+18xlfMhSM0woyQ+k4qDtsk9qZ5QtQy9jL
Be/4F0HJkicRfGdeacSh5Y2bY41NfhpFUxJ9Zy0WSq7axPFj9qds7lOKcai6
+eNraW4TDNRjYuMWHvgjCRxSkpu9t1YY+pxyJ0etqz5UrZqfT8mSOeYYWz/J
+klGM/szv/2aqX/a53iF04IcP7xqA3IWK1YjMLdYWxQCMImdiZJuQelLUqkw
23Ryd1ChFi32kPj1MBYGiAAyKN3N6lPEcZQtaXsm9uNp9yO67wHDFVzSKaDn
YshgANlF7Fb1aRD5A21r2HWUyXW347C/l0pWbCqMGG+0ADL6aCdCT7jdothe
N17Zkn8By5p3UlHkIzFj6ZEF6xYnEf6UsvP72X4TC3/Pam0fZIrm4+mwEW7h
uqkRSD3TcLs5YuG90YAXraw5/jXlWFy7UKmvqTqWkwcpX2pRkixcjH+m7vxU
1IE+FpJNP6DnYUlITtvtC0NaInrVO5PhjodqFPcVI2LtLBsA18DpvLkL5GP0
1PdFdqswiGZPesGFBlSUWQL/AXARAuV8qwU9MuQN43VL/16/9m8vU1qBo7g0
GTbTNyIK0af3i/tgx19dKLuwGxweDneBqKITmTJavZrP5b/oVUDVD0QOiSVo
lNh63Oi+hWIFw3jRg7G5bPn0xRW352lVkBcMvSHfraKpvGytBBGEoPjIVmWc
LMhlnwG4pLEiJQvLEhuhJOtIf9U6sA74Y/VNK/e75BY036y4aw+ruQEKyyhb
k/pJ1UlngvXzSEA8WcaJgbX261Q4JPV3NSwsq83MfZYjUHCudw6MQMEPJ5Lw
EJKoJUoC0iDNWVoQ8pr1UicpPH5XTcVRi76GplWNXC9vV0dDChrM2PzVcDWZ
dtpU3RFvwwHXq3mOZLKG1ui31FG6DEPkcEv6m0lURHKW1/MshjBOag+pcJFt
VX8o3B0+l699kPkImd2mx/A27TvKdlowef2PeB6+nCmUIMRNRlxbcrDIRZZ/
qxLco+nyJMjXQZA2Ww/WkylZUhgPI7VVzP4duYVifQWhMFMFAkg9DNUIsdg8
5VKSII3DdoyOuOPA4hsRAVp9FaZsbhqCdoQlugHlZecDm+l3SPLzwRed20Ao
svCZB4AkWOYaCrsPhVKb4LgrphXU9X5FW29UQVMfj8/V7eoJUN2v4Rubt4Yw
N8GPlsRe6qflvvwQzGucTnU4wnZt24l2H7o/uk6/l+GFFXZIb300dBIQEvDA
BpkFHc47uu8I7XWhYOZ7YMQX0MA/8uNALWsjTrU0xPJ6Bta7tTzEX2BVKO6j
VXGO+qT4QQRncRsciv20qV/TsrmMlcNN5N8IqNZoitJsIkMVorXbrB/5oL5X
dEEhqmbbhJcao5y1/E5lw99RAXSDZOHoRcfZaZWQwzTewmpx3hK4/HExOLyq
GydP0e7yfLYqL/ffLzB7BCoS2mq6o+qvvFIoBLlIwPgGwsIPH9Oz7Ig68zzU
+jdthP4zxVwh+ymJIT/UK3bKQSMum7lCPMwNXDe/qjVP0zLNT8yu9svR3goI
zzGVUu+7kNNQjDG2qds3Jsyg9XOqcyob/z7no2/EmDq5OscJCF/J6vGZqXBU
wR3zMkM+q48EnvaRma/CKM3K4OF7UgkbujI/ANU08EUfjj61OYWIV1y1f4kz
gIAY9WTe0vtiamewMfmqvWoCNwRdEsyTrd6pDMPQpe0xojCYOYM85mZWYEHG
sD6Ht08Rz8VY9mEuSjtmc61UkmaGYoxYjOLcwFu326HsxWX0VOa4sHn4efcZ
x3WiaICvSoRCT9z4K2HiZ56BYRH29sAwC/gxZf3uKe4iwx15Ur/qR8EchPNe
Lr0faed+TNzoZUyiFjZIplWOingrNpgRKtXP/pUM3zcyxXydFyix3RyLcOlM
RPp+Y+ICVcus0s1A/YpPK5B6266Il9w6/bzRhiELVC7ql5zVLhc3iXmmdcNL
jVGn5CHlQd9mH8HTwB012OKDR+plx+7ROEF8HvJkMdUaX9KWE1gCzxxcgJ78
LKNPypO7Uj/EaOjNQzjQtqwmS8jkjZwNtTjXxSd4SuL40pBMT1cYoj3M6Rgj
hPOd3MWfCrX0/Z0lNp4gk5zY5vgmgMmTRJGBiYaaPeN1Xq3floKEvFTl05Xp
aUKsdjtSBfLkbB2jRKSmFzRHWuhInY1gPgOFMDYE0/bRAEnkRIAkVZlLSDfq
1bh1qPJmKfrJCSP4cF/36YdgmxKqH9RLb4aJw6uNSGGeXyjftQyYm0f0BAkg
hI+SkxQCWdeO3ANLWFP43td1z7BkBmDvqteP7vflmwvM8OW3wC8I06Wxbi8b
5fEiC/1H3WPqPFaIus7E2W4hvhDA8IROqrtFyWB0l721taBVWXR2GZLqi8f2
GsDNnv7fG8NOUt7ro11MBNxgtveIGjX2G8eZHQOG8+fXdcwdeo+U/eUyHjeV
nRa2qexG3tjzJpgKkRH7o9lDZX2FDLfELtzAdezUxzbyaZJiPO2KzDmHaizz
hI0nTk1N+4okRwz/uuTIZMado3Ev+9bnEZX3lrwT1cQP7mqfPi4gAmsmb/iU
EtC4M92KogA6sZRo0+6NHAnO5dJ2+hdCzcMNacnjd7mk2OExq6jqJqgTofIl
ejZNsOF3LL62xUkQqSy7Odt/tZaw1KCNLz6XNxIIyzXPfbitl259KA6qKHWz
VqihjhDU3bjZallUOa9Jv38mz3A/0+4TgkxHNiA/ewqGkGYdS2UrXWPNuiay
fQAv2tNsYAHfoS563W1IoCpfGs1FsxW1ng8cWHqtJRlSMvkmamd3TTJUAHUq
V61372J682yp576ar5eJXx3c+guNlUZ+6eyySAXHlaKTqkpD0gw2LCNIMZIf
27sT22UTaqReWb7QfIHy4eGMCiryrPMmH0Bpue8VeIqoHAgmwR1r0iN5QIg3
vVBE7O2dq3uzl0tF8FAzwHnb4JJaMetpH9kN9XAXJDYGfy+jhYoa3F6Ey78K
t6chc04XbxoosWHjbc7xx53qw9TIIcYNAaKpcda2lD5IWzzwupRxkgmuLIrY
9cgXChT+Tmo27zYqTeWtjUi6JoGcO3gTfmmAy8ktJ5oL5zaP1Zj1xhNVMjLz
y4Zn8MwQGofEZhoYSj0wqkqFjGx+QgiFcBjkhfMeNqzgURQc4oSezQ9zkxlz
paEXsV0C6Ly8ECJMVwk+L/NqDqDtVrjmpMA4Sm47xZ+lW/RnT3yqEK5TqFL/
/82ewJh2DGTd8nfXHrX0iHqhuC+NJr2RwsP3YMtYaKvgRnGiC2/jDOH1DG2t
gR8Bw/p/EvbLyUA2/MHBuqXC/EekRR7wAzVAgKt7IVBRWRmA3EgvkLvERiQ0
KpCA7AOcT/u7B1HgSoOvM7GOJIgqTbU5PO4uFldx3rkb+yxwWMZTTKED3WK/
dv7n6X3m7TsxVyqqnLw2e1KzfGEqQF+BTO5woNVZBgdDKdweY7Xn1eYLMY47
0l2qr6tRyE/R3fSPuNThZmYkq+KYZFS6UzLijb22ldww9Tv3UG2xP1BpAP0k
2k7sO6CHdMG2YQeR/U24e5hj/OlxmhVBeM3mkYMD4m7oacGxol0liojQ27ON
zY2Y1pOEAm2ZGM6BN32IVXhcAc+2KG3s6bGnO5GlGg2nexsfCff4VBp3S0B4
pp+yIXxo6BIXkCdE3MCcihwbOofjCoznqTUVZvh5LDrqYfIj3OsMmqbJWc4Y
gISxNc/oikbrCPalB3Tkecxj3X+GVYeBlXX7xY7aKrrP5f3QD0+un32NazpX
Z5ovvKIuqxlzvE8GdVFfXt+P2hslU2XF7wXhu5isjglRb19tyViKdHB7RSvq
+yViGDaly+gOjETdJwDThiGkX64hqSWM8CEGxIoqC3otXMJiKvh5ixZ1Mkvy
RfNUMVIY6rVIKo8ci9XX11D6FBztrMOXkZrdz7mMvLAmAioeWj4yKeZmS4NH
M//f01/AyIXeWE8PsIf7lpCdbj3Wpd/dU6ZEyRfHWz+rxRXt+F5JwAazo3eP
UEihWxe+V0U3ohm6pkiUSpEX2u81DRGQxdEmV4KUT8gjPGGSQVEzV/bmT0q2
Oz2soIsbyCbFYV+ohJ+dN2emutcmH+yq9mzte4CkKDBJ/KtaEkWqG6o4Idx/
+UUa5HbvPXVwjvXnbFhwxPQWW7kuelY6JVDHfWz2FtIoBchdBZ910MqIlyZR
72zY6spyJqILRFDxYUBxVoBG/ZZ93j1idUFWT0ahLI1c+ircXYma/iNzOFD/
g+NCW6EbCbsV+9TfsBaLJXfWA/r0vsrkEucUDQR78qWu747ZiJIMW0mR5tuA
D/C36XMHukngyucSdKz+KCC6hBfiemjX/BGrejw2WB/KqjntK47or83J7QMc
iKx27xaSUX/vFgOspiyrftTQGba2ziq4xps1gLmJx1IHX84P+q8r+AeujoUA
N40GUFcWAXifWqsrJKnED2esvc23WE2nyDGp5NX34BZMSXX3lRR++xOesvGK
qdvdn63ExoB36TOnMH6EFc14U53vW6LbxAcgR87zhjK7PBSwJ8F9LpyCq+b1
kzwHERujFZqfF8P08s/gdf7g2uRND/PiyuXqJ2lvB57z1vir9NfDQel6pjRA
H/dipRbmBOQO95ldTrwiNW8wZ0GpJ4DEzZy2Fs33T9bT/ismsyJLiP0pA3YM
6s4pnotJ1CatiFJ4aqA7Yv4qt66XvAHR+uQGT48/Ik+22aW79habfw2v9I38
mrsAwsIO0AUzxTqHZuqdbqJb0QrezEDo2Zg0VAn7YVDHo4nTWYkmW1ZzNeId
B0u62wItSVVcweYa/qr1CRblBLXr1etbrG5zVbylBKQ3a4W57+LYw0i/rM3A
QTA2bj0cO/g+rs78DAyPcidebBf/UCJQGLBhU3oO1cr5e4QkSsl1ZwKU+hOA
KND9miA+gqPQ1WnClmweg/UUcYzXWq21EqO7QzQaHQYTggZOOENaaOrVH6gx
Ez/pSKLtGqRw0i2V0BPF6SfZcqVLsdYpSlYk9t/6eh8nF5BKuOjlhqwkd3cf
LUZaFFGYCRWyf+l1YVpRXseIG8zwF03azY1oudIpfFLJ8yprrgcDy4lBSw8+
ztBbZfjdQsfjJ5DNzGvYlOCS1/MCjIoKJGtpYQBwg89Vv5/iIrJOUsebQL9y
e7VcDtYSe99EvRhAQE0PLzaRUzMzkUUuLrxRLiSmonwmEU8ysBmdh2MBrjFi
SGwaqdNQC2mUOUKjkEAz/itUVqDO6ixGDNDZgE5072ogxdwTnMR2BjlzBvEW
892rxwtSpwnx/NyUVQPS7TrNNS2qRPPVNV6viy+p7eREK2aTWmdjRqu/0edM
mPpcYyZ6L8HaW/t6iqV7NaQ+ab0vA7V9ebEzwevcAFsU4/IdY9KWh1zuwQSF
1Bg8mZPn5VsH1alwV5aYYQuL7/Vop0jCN1AlpnFcxWIDYSS7ApkMxyA52/p4
Wmn0aqtjbs4o4/PglfPVM4LEgrqILCaFknSnnQbxalpEZwh/Rq3TXqLUTBVp
sZfO0mtCoN+XKU+V5zwG/+KAvnoB2DZG7yXyAPh0drT/WuJJjUaZPX1X4fCA
uS0hQwaH3RSFLD4+y4PxCTY7oEm3QAoH3pxBqbc91trXoveH3vIXsSfLlovz
nRQD3FPZUHxf0n75mrQqodIRrYKvF8QzF/gPQG5uCAKfz6zGsTUsExR1dfJ0
18xuOl0O2gN/Ee3FPfnJ/iSbdKfmiQLfJV8V5cR3a0Yf4YRwR9hsf4sLHU+b
kCfbv6tICdrBPN1w+jbnMzw/q48xfbIMnEVLeUVSF0Q2Xw44l/nFRPhvywmn
70rpgevr5eoGLO/vGPY0yCz3dEICkOT5p+TXF2qX+1FnJq08P3xTTzK0Q8mk
+OjY8xr8f72Ev5mdueeZtpjMuruv6j5Tg9Z+iKuEFknxUT+2+qGOMcTYx4UF
Rfpt6y3878r7HjHZRlPXKaDRopKYtxqLjaCyVv79DBBDkOZWDkmVDNxrdoDI
/LXtVGcC8wFxmtWj/7B0npo2lUIohjh+6oaLCc4VTYUys08kK+0snGYWTomS
CtSKzpH8zXjYBRVJJNbPJYIwrbpBx25Z/mbdDk1L7ZTaCuPdht0i2CHqT4LM
aQR6+DaDAF9T5Um3QOqXA7bhyNMXajN3aWLfQ/5t921YT2feW9cy8lMTeBl8
WmsjWY9N5BtIX+fwIHtp3m5Cifn6zDMRDSSuZDLaUHlNwHIGh5Xk/14d5du8
53y3XRJ4Cu2E/qrMMxIlWnqktDjorQxhQFtmOV+GaJm+seSLsrJKkMzajCPP
cgw9CZ0WaxgH3gROz+XHYJL1dbgaD9v0gllR93hTY4IRE9IxxT/vNYgU97xV
zJNB1wAfsjFveHErnS/OV2uWueLGs3QKMj9kfh1HkcTh1P+pU4+HuR4glLsi
SDGiaDwLAdGcalBqrthe77vtOY0i2kVD2HLnsfsNdstvxHZolrnyrbR3efyI
4pD55VS6644gRUs+o+cYWvNDRfPPQ9XtG19uBeV1KW9i7inI8J2RSNr7z/lP
7HQAf4BHquIeIKannL2K8LJ2AUt6gpyCjfHzsCEePS55WDF73I0w76T7/SX1
pDoPUx+GNs0zyfs9akp+8AslOMPrpoYao4LWIozgFISY861lApRW1BtLqIgy
hp7gawR9i1ybYwcKj+R/vxFUl/dpW0M/m5Gf56ZiJByAmyHGLbY61ycFj+Rl
E+a1n+9Lw99NAuLOciIqGLRaCgdM/KpigDa4lmjeb7OhKz395H1oUemeMO/z
e7e4e4hBCEHbQaFq8iEG53oq74TzJPoYKhJyfMrU59RqEh1pmEJIWru3c4RE
lOaRVX0qdAlxdzUTlt8vN9g/h5X9EtYUPskFtpdPYuNNV9KKnGEb2bjqS7DH
nfnjTWIZeO73zaPSXPs2Jqr6NaumCGXgx73ct61DW9EMt/DmtJkx4KvShoTd
ZNGsETdFZpSku+DJnbYs2pQd+CvHJAKO5LcnJ/0fREmysSe/kVlvSthr2lx8
yI7z4FffB2fwQJ/o8VpTzOI6vTS0aoiLEM+EhGL/dPRGjJvKPDzvHB2uWEK+
eF9TeNFBM4PHFLhKDYD++cOddenXfxpZ/cot+Sm3mouvEA07gTi+fEn1BbIH
xBws8v82pCy3yK3rz8SvzytEgskJyLf7dspggNyRNQssyrAzHZnTfzp4OYXU
IVFfCk4WmlQ1YDY64g0IYylaFJu7GyVlGWE322DyVSwYxXfh6TsAdmWw4Z3L
vuyPXrFyMy/cHN9aYH1iJHZKegZk4IYO2lcdgq1rm/F2lS2lK7BLm6CUf6hK
X6mw5dIzE1RJVlKkT/YTsMtY8zlKjE7mw0dX/wNxmFHOtG4OfAkoEsVoJdPE
VWgM6ZFDkCpG7dVJVGrhWyUtElW17keUe5jYjQS3W6QBriYD7juaKLZYgtt2
TmYcE+FLmdVwGkHssmRBqgUkUMxucZY46tc1gN3yCLkg6g4Kl5hxq9yE0Fr0
HTczRDiGsafa4IFVgvpYH2UnImQSgwvOlE6VXxTIwCoP4mUv0ncta/qLs7E9
qFAaECieBdnr3j582mwHf/UWnRV8E42A5j6jQ7pBefgGvh8ef2ohS3FJf3mT
o7JKpIXaSeQ+ZXBaJXtZlVOIfzOuce+lv4H0wGX7sunkDhFMlerjG9r/8dqh
7AX7Wh3IV46AdPguCxRLcRIQ0sWJyuRNU5cjswJSOuSgHHwR4sLpLB3lFDpR
OxgTIswTiTwQ3O7S1LGyUD5CltGX1WZD5TKrcBqoJ0zBYF6fiH9w0ET0srp1
MmgMMsBxlCQSqZzMMCDCUPc6zlpwE4sY3crDt5bHdZCB23+5dSuafBnB77Gu
LLs/lPMgB8fHR6AT8+mosGw/LwdoPj5xOsTw1mEhNEUHGUbla77uoR+mbzj+
rcbWxBgd16yYLrzJxWZXkvEUNvs10E50DGqYtswUAPVhLGRaWvR+P+6Bp99B
4FSKxzNb+ubTuugcHKV0yeLmhPyaY1sSFzblIJoUe7FNmQM70iACQmRQGQ7x
2tZuAN34h6tElGEVxGYHG2I8nRLfVqwuxVR+awJgx29J9vGOvaLVJXrph/wC
+8wXfIw5cH7Ca6VTogMnyTYsyalAySaaTwDg8vKTzyvtUaGjUtmd8tGRHKYW
OHOjvMnQMQsavfAe4+n0vFxXfUjVVpcv4nk4Bg13CUslCalepUCfEwOiQICQ
NHeL5GRujyKMEs4ks1qRdUKfvf50R88w1CoJE9EWfcz7myCll+/zhnW8oClN
uZJlGuT+Rrsb4xOcQmT+6e86dBY+uXkoWWN6tsXLOa/IP/NpWBv6hMVR7061
MPZzgaN28CnGb32f4jHCxEAy9h+Z2p8c9vF9A8bqbikiNHI+o6J2jNaSctjT
1gEe8nNOfvG1BUZpkrlC3F3q5SR7q83MD6jHV5mbaaWnc/XlYZ04XeA6sN4i
fJBgC4zAkyVvi1DgajdVH4Q+U09JGQR733u9TsVKNGqlI8c9MSxIWsqNSrGs
O9rvFYSS4ieF5TG6pkAQ1weejMlVw5Cd2Iw1VNs4gjBIgX6p5yABSCPRvGyg
4gzUgE+c0pEeEyd7fBOgkjikDYjnwY+ZKAsTo3AgTQenKpyJCNCV6RP+9VyH
1WFh2uRDqt7Vv6lbTffuJ2YBnWWzN6PDX9itAQRrppYTVpypI79wX7wEuURq
XR+r3rpQfFN8M+FluQE1I36JAd0fubRJ8FhYv6qhVhfNhnI2e22ZbaaIDGU+
cPh4daw6LjMMWdxNfnTrIRFnaXe603+CTO/Q0+RqqYVPb7pXsYiBM2ThkMmX
bXKKtyC4PYtg9watVVNuVlygLA/bGuA9/hNY5TBZnZohQCXBM/JX3qrDZYy8
u76pnddje2x+APV6ig9Sl1jvF6RoN+aiFfgtocDDv8Tj5E9UUAoifH9QgnjD
PMXh0MLFERZAr4YLQg4IJ7urDcT9+gA7Kj+1lKKm3im7/0xnocnjCZzAg6nv
Ch4QZu1rU5kyS23tYKnhfTZnt0dd8Ce+2/nadbVPbJe9ECI7gUgN+bMecHgo
1+kO8fS8NdeHFa6hESbee0dq7j5LuOBXG7mW9xwqXWb9Xr1SJvSjLEEoqBsz
EBiw3KMBiFPOgs1+NQgiK5CMCyom/jedeS/M30Tw+pHeLdmKMjK1YCuaB7Pe
qlo6IP/ro1WfPqrw5c1lFxFRyBrdqAjCrUfdPlZvLROTUfr25Z3n3hIIcw7O
PyaNQP9NoRnqRCf38XO6sWXjC0XZbQAwT/nybqTBoJITH9DpY6A2kvsmFiWH
W48/QpnIFc2aeFOjdqaTVEyWyYeSjOSCuSWvvxbubNnOh1kTd9kr9qcZi1Nc
lT6t81+83K1ZaFXK9ef8CkAGmk/ak0Jca3viPxMEMUdbiLbj0meEqXBh4nJ2
qp8DkgmEgt1JteQsoG3p+wHKseoROqip5+uhGaEh1lhW5tNVKfne5xNDghNm
C49N5KxOcwXbjMmcUVX2J87hgysu1dqZbPvjB/YC3vL3ub8yJPZa1W1iguZv
sFQ2YWr2yvHPKuWNOjj/hkd41WeBjvz0ofHnanSr7jLGXDSXIRq83Iv6pnws
A0YrmmQkBKXvC953YOnEgB2uJUOfeKwUu8F2Vzd59XEgcXMrah/KOSry4ljG
timEKNl2iBX0xPVKVmOtAoGDfFc+UY9KNPCSKtV5PFr6zbrr4p7aN23fI4vV
UziUYOFBwDluPNeqA0GPMPPZjWiPYFK0Q7dT6ftwZW0h1bWXkXTXq1Rmz3Db
b9IaCl4NYKQuEV1fWbG03ksk3nijGQXSWL0sLBeyLLwgNNBeokDW+ot9G4vr
VwcMXDxAnHOAHqExJyHOQqC+W3ucu8SAUv5GZMbGJy/Fk16606c14deZQTa2
4mWoTNxqqMhwu1drWWpAQKo7rCvIB+Iktne6oZyRuTK11+SGJXVy5/KL03rp
TB7xXKzotyV+DtomBueif5TcWfFzHataRJujhvfqQeTzWiU0zQtJvEu+XZqM
2ep92XAFGmCGPBba+TmoeqMxlgTManlomwOJj/UMWK7uiYWucpLdW/SZnxju
/+lB+UxA70paPUii0MlZKKXaEmvMLAdNlx2QgfM195UerLlsi81IXNR9Qpcy
WVx4NOxw1zE/zzzWatxiv4UBS/3Vwa2BVaUwR1IckeYJZOJqBtMaMMBSNlY+
OX96/JEY2XLfvJsi1eTsojKK5ZOJLxLjZzAQUXwWuaAMnhCL65rPcROKkIzS
hvNnNLZZRLsK6TmRDOpfgqwQ4UA7FX2yQ3X2mcirSqpBHWnMKXA8vuCp7lic
ZXqqQxnRK1px8aws7eRoXVY43V+xLWeZnZMPWCH2RF3nfoBfNxo+SzFZQZdE
acchktfPxJye0WBFpGhLt0RjI887qMvQEB1FJoKxM6MI/Ot/WH378QeKf1pg
IDbcbGe/vLFOPuhel1oyOupVOJTTTYL98oSqDFAPvb2y88J54YAtIMTO4VJz
XyVO458743zJEKswvBCaIHfeb864fSK2vQXnD2/nmZckNXBfJ3DBXZDyiz4s
GCOiu7JNUa0NKJwVCCpb1YwtxMLn5HUujbeABcGNmVXE7kC/Yg4etVSPjbwE
bT4dxJP8GWWaye8dANQcvZ6v9Vo6XEiCRtYkt4NsNBTH+4palihtQxAXvcm5
6wzxmbodmv8SRy9dnErtDjtp2mDkn6SaZ170PuqZew/dQiFAO1MvWfu8qgGs
qDQyCtZyyUDnkMz18Dh+ARHI0mquIKn6Sr/fhPg+3IHSU65S0SK4j0zDFk87
/23btivb8DHP+liqHswzM9qDS+GYKHAaaL2y2wynskTrStSosTTykvjZimPo
GdHg/H5ZD/P5icqysRcCejR/H778reMEkIHG90zjXnWBwuyqawsYXu6VO39Y
q/KH653idmUSbTYRlGRraZLPHwttnKfdMX5OV8vwH8qFDuvrU4eKrvcdd/Mp
/b7NBr5Ux8T+fiy+JYHbkPIYYdVJrswN9xG4FcjGlos5TCFUbIsjKLTFB8S/
4Bc/T6MfFS/gq1fcD8Th44tMEK+PQUxu9XP+ht3razDuNjLOaM01O6YIafiT
p+a2k+Dc+T7tmuX7HvG0XWj9sGQ73YIz0NtXsRuwrO1Dm/Ah/9pgjYpDENbv
GCEdijp9xq9Z3mrmN+dQmdC2/x0Plz6lKEKnUwpUujr3e+Xbrvq1H+ivD+0b
Lh2W6gLXSNPPjbqcXxOrWPi5NA3Y/PIVmwOA+ZCVm/ypfAXRZGXNjHV8ZNoo
G+fPjU9rzGoHUxIjkqH8GgH+Yv7BVgf7kfgAFy76kEhXBYs7CLdPskBJcCeB
A+mk/ftuCBLHY0Ez2HCSwRR+9Bmp78Eme8WcmzWuNpiyJ9jYXCtmZGmpsTYk
mo8G3sN60RGC1TPELIw+OBEiMtPFOCtVHHihH5pXigWFq8YxPyEAo9O1hDKx
iA4JgZrQ3GSQwTPMs3L//PARggHB/d6P/cFtsZaaGuqjOM2DtfTLfNygnw1z
AmMd4RWzEt0Y0vJmzn0UlFmDU6bBMEs/4W76GFrqL3xMEJaxlhReIXzECcv8
7jasUVxRANWCMhrRNei5Lnw1sK0oHhOXsBixor2OxnnxE+jQxMcE/LQ0S3RW
MeMwiooJAjt+9QuNVXBP99RrRrPnpAVNdw9Eb9eAaI1/hJHFxsD2737B1Ajn
oVUow8YrNfPpz0xrrdxZdudlZ+i5bjnwZZUo/FjCvJWqX2xActAucyCCNKry
VtH01Rr4V91OVaF8EMJyky0RorYF2KEJdUdTZVD5FGSMdyXZau7K/jA3fraX
gQGL8wjeKrj9SSLLmCrg8mXbjg1glyiRotRzylPdDg+YO3c5EtNRfka5W9+D
jSgW59UHEfgiUYqoiyf9XQQX2WUaQA+k6OR79p+jSUbdZTxMjH3WmXaQPzS4
CoMHoyS55dMpps7fiKwWrYvmd8Gti8n4I2b60ixnTRem57nwN2PsWlP3WaQC
0PIKXnsGOQJObhiNCSh7m0NOKJkrXJru54YTqt/6OKNBTlRpgOD/r3efFAoI
sjbQUO1TdIBrUvKIxO1zBmSZgPu3KPVzPUvoChcG+DEiIRJFvAANSdCRadbx
oTt0uaiQ6/l10KAlMhEg/VmZ/4VcvF3jepTbkVGQ9Ca1dDtAPF93LghUbpgU
QQw+s1l70qTZkMa+uvn8BANI0NWsvSuvZq2ImklXejTx5rLf7KWRZuT1bTKS
+gw+KCroC3kS6/ZexpxsSj84LKBySimHc1Dvo3Qksi6laYbkeR68UreLWqZb
VX35H3Dy1+/u3wONJYx63qJv2m0+FtK8zsZNsnzeH/LHoYcmj+RdGHZSUMeG
HE6zTLJaq/KX6hlVW/xX8CZQ74fKJ55i3tfG2/naiVLC2KtMgjGrKxYK2ydp
Dcdd3xP5oZTJw6WSheaIG33BSDKL4og2jemi7K7DseDJgumJTa8mUFc2GTap
B5KonDyRTEK4MYIMZfyLTiwMJ5ztjkog+Bm08Ja87AHFSK1M+vSBPNui/0rn
hxyueb+3oUBdWnZRaUi9jTpprUxJNflcElj/ABbgcukA5+cqoJJBKh4HFCzY
Sw14JGoemnd9ylhlCnotfQFneCV709ltZc/qRXiMEWXgfQqSrd9jibBaCUl1
qmrijqEZAN/ckIIEwgbYbgae/QFwqo21WePn2i7mBj5m5ZTts6dLt4k1x6lO
0jTZHnYVUUaNQo5aPEKcwsXFaBXraowxgJA4hwpih3/nxQ7ERz7ZjGHWZpRR
bY56Jl5mv5zANseqYLT6L4zWUgNlWOamFk47xK/awIrFhUnoSTm0ZCZz7lA4
tGIsd/tyeQ5Tvg8cFHWjciFoOVNbyKW1l566dwv2cwKgDvWatL4no5H8l9/Z
7JVvEFNS1ZIFgQgsan6R5rnVrZScYC7y4W9kNsE9tOoDIHkAx+fEzQQPtlxr
68932ZprorOKpXBWustjX9xe1aHSJKtOBkdEXAp+J0rr5vk+5s933SHkwrTK
5WYEnXjOWZ5e24rc8egUAzoSUH2AtjngFKHTTYl9zI9iULgKUSwouhOxprfN
/wf0GtryAnipzVmmUzX1XfBwJpToXf5+UXzdHVX+sKYMnrJ1ZW58IiyezJZs
yyIR8MfMNdWmdmMcV8nVIZ4yVdVxWI0hM5SN2CqDspxvdn+RpyjNWseJYJlt
1jqRXGhelAPFjyIXLlTFEAnqtCUeet2A31YfyrrtVoILmpN0DgIKHGv6Rqem
hustHIuG0x8aF3zoVlWJf0r2c1dCzNZ9QKGEP30B2k36NYcdI0IpQ8mb9Ldf
1OOeyTgs52ywtyfUP/gurUYv8aKPlR2JIfSfb5xSFNkBqMsghE2TFcyfL7iY
xNC6mjxC+J6F/sTmFo1gHl3gOkt89ANMvJwE+u4SeOAK7ukFuxnufydUbBAF
GZalBMfwQ8RqI/2GJ03lZn2WosXxgzXi5FNIqBPDld8EU5EJJnjLCn9YLzan
VMgBsjPJl4jPPrCv4KD510PGTtWXldN3zJ6nedIN8cjKDerHSrBbscWYNPA1
gLKzF/R89q0QzHbox9aPh4Pgc+5/uuQWd2YNPh/2aA9/iZeJg4W9NFLqzDoc
hFpSm0sP/yZdFRSOFxNExh74umlB6xyIOIqp/fijmaN+zUjunikMD2kNkyK9
m2cYjZ0DF4QfDiX5eyKNby23hrQfCXcydFA4GrjKr/jGtRxXsqoUjMhJYqca
psINb7CLZNtn8/nv805W5H6rrkfm/qiTZGOIYAYSC9/pcGLlGl52jy3tGAs3
tllPnGqDPGzaiPxWNuumZ4W+UoGW2OLCGXoeLc1t2pNeZvOOFcOzB4R4Xjyn
itNIA37OZrtzQkR+dIfuuyKGsSnQt27ydG4uALRcM0640Di9HAat1lpAYuaF
xEWZ+6pQ2WJAKYeVLLlgpJV/vSnm9YJaQZ4b+Tw4Cdj35aFk3sijAcrMU9is
4c9tGYS3Y7DcRAQwuP1MxaqSNsQ8Z/ouuRVCHmDpHVL1uQ/c2AvSvtlLqg8e
lxJlEXj77uHzNquXjdvnz2g+SXIOhjOUsnZTye3j7TrP4aYE0RvmIlyqGWc+
oAhuIqo1NHjHQqFZ4OG+otYWTVaebW/NezLxZtdxAUAh0GQjDiKSZjlJiTnL
fIwoB/S/BO6mS49tEvAOjOfxPecuPCDlys0yFDJXOSWLNBuj92cu71oK/WI/
3YTVtPUfUz1gdMGidTLJyPyQSDQjmWeckTliCMz34KAmWJQHDyVIPMmVoGBd
eMlt6gpHETFk3d5Q+UYYZS8eIYYRroFkLL6Prn8bPRIhKbFvOiHcP3+PhF7i
1HErCef4oCZGKYyOJFHfQHWdZ1BLJb7+tZvPeRPnSvIUuc1+QmkFq1EWNewc
yJbWTT5WrqW9rf+NBfLb8+Xtyb4haMeWLsI2f/1YTenQF0+6uO+Rxa3DiC/r
NsK+t1ieVCvWXqo8NQbbfA78qkH3oMZVgyZGAnbej27l6t3z2oz4NPHpkRoz
QJsDF1lcYjtSj4pAat7i0KfhzqNZkvm5l0lI7r+YqXMMNpTTRiihrV9zfYoe
6tCzTavvQAh4KF71A2mXxsW5ucsZ9ONtH6dIUvxNC5YbejQBIWWGxDjGFRyt
pJPM1ItaMmqJnoBfCK5BsrbYI5J4YY3BtCo8WBhz9mkfLGhm5vSWNX86ITgY
/DEAh3vf8x4+A0S5iP6r8U2kzGbnB14GtAZwIV9bThOHZYL0m4PW0NDqWQK+
novrUMKTeyhpqLGZFsOWunTV9qOMIgnwlge3XuyEmLnFNqKI+nHfI2b+E+yo
AyY6uzryGGlAVAcq4BmcjkDf3AZCU0SeQ5KjNpgSW/M/QvruD99Q83KCZQi7
u06var3SmZidx3jj3Flq/Td07Y+MCtnTMOdwoxCDMi2P/4RkMxjyA0zVbqQc
zzSub5Cl08E9H/iPT1+aXzittE9ftofKsxvPFtUvtB3hIjX2W394z9IZNLAN
wf69//t6tQLyXV8L63jI/qaLJBC4BkVvX69SAu0wTcaPSTx4jGR/BwwERgmZ
xra31OrV/psKTgEJfNSkmUgCVaHH513ZsLWSnSQzzHuy558bbrW7eAcxBSVQ
Yjal8QrXkKcwxRpvD9UCr2osERsuywa6ti4M5TzeJJe+Pmv6iDAxVR0cQ8L9
PpOe3mA4KDaIr7auJDsuALJxCXZj5iQniUvXSUN/YLmegvsn603v3ukg1KHa
XHGBNb0+/klz6XwigcW29rQ3dRY+NBKBTxn4hmWe197+XnPS7oMBLm0YKnk3
boF4+t/SmBbfQ1utMNO5GOgrPuxiEY6TeZV3Z0VxDipUaSnF0MYcHVzAPc2G
7ro79BIV+qZEOZAbyX5/Px2utbN25w976X7EpeEwFUkwpAZFmOvGT7xgaOUa
4GmaCbnQrJSJmrGkUq4OpKszz/EaacuyXCGRcsg8UmmGmzxS2eGIK7OniBti
E5wUrT6cwqVP7vpu9lJSsDkjy5tMdMFGVVoNe4m7KffSQ9qZdvutsqVw0n7S
RJNNwszESUmdz8zBdEmVahDF20Fx6jy9E+YsEU7ZlLCREnlvfSnvaKAneCnW
YeVUn+MvtPpikB8C0OQeHOWTlR+C1Yf1ClDbS3V6k8LzsfIsERml88a5o/4n
7v1Oc8qO/kKR9uC+TGzqnZSdVD/0kx0TmIzZBEdFtD9XrU+f7dyA0HCzZ5m/
BWnbqdlvhCNrucF0x4SwUu0y4pxEJYsP/KlhAwmLpY9owDPEr+4G3e8QLO9/
UQHsvm4bsoCb1hep0M+NIrkWdizBPt7fRexo5YhZZSt6kApBBhKJG2iotBau
oZ3Rcj0D9naL3tdye8tlUG+xIpf9mePjs5Oc4B7Od1Adn0mCiHPHXDjU7itw
dtN9qYdjeU9WbLtH6gF8yImwn04wjMVY+aIicmBOeDREQaRFladz2VsTwhCH
fE2i1dys5m/UtRCIuZqilPxPEDS6jm2e7kGzFg0px+21qUTXaJLCQS1RyyfP
OEgSi4qNNWEZLZT9pin1Crhc2F/z2a5jjdNnL8QO69v4SQ90/0mzOw+Q53Zv
IPtdWLH1sXnnOu+x7TMOaGCCz10fWYpt4F/A7QN3oobtUvDkKrZkW74+prgy
IlAOMPPlQmI3GblQxiDf5E8I94pHLjjNNvlLMc6hFYxMWtmq5BeG9RHi5Mds
zqKzzfb1qmHE8t0zw1mg1BxB2Bnfbg4EMLsf94UYz2gxtkXLxV6xll0IdRyP
6vY++HHTUtLj1nyblnp5UseGFeQ2jcnoLEuevkxGY/Le7aOFEhLaDuv6P5zG
UKh5VFY3ACvHAHNs0BiOqmH/nuSukrWAKLik1bVQUwdcIpfywwJ+mm4I8g8d
/+a2Y2FfaRfSEmn0yvwA8pQU85b4qtjxObRvB0nV8GOc9fTHkBNnje0SLzHH
f28fkeEf+wxnj10AxGcMAhgVCuAEdu7eQNYluQmkBYdlHaIcbjYr8y9Vjjhu
lz/ZMZCh5eRDibzZCI47NdcEMjr8zOlKyU18kFleFvjrMJ6oiNi7/LBI4EZ4
zh1VH48GQPXY00fnWSEuA7Hfjgm7+tI9257YoDVp+J4xxOaIAvRWIwuw+2Yo
3czP8K+sld7xA/JUuRrWMqV9RrVDB2dDo0Id91SQzQS+358S8dM1JXWNbg1p
cBmBQgK8SHPPOnWUW+z6wwUh0jagHns5CivPZkbaNhcqtu+yryypaaiRUuYV
YFE35B0K/9Za/rdkVZv18PHaaPAh5JLZAiIXsH+IjLtOJJHxgo2B3L65V/KC
yY4aHhG9TLIG2fZx98GPk52Zcdd2Xjc8n8tkE1gUjC0mlT8f7Rtbj33e5KAy
kNhN9TjdJeAMNDk2Q6jwZASNrAkJTHByEb2f5bEyCiJJPC78gzfQEvo5IbM7
Xc2CNIL7AukYWAtV+v3sBlrT+IAVXIrmSJvHZSu9U8v6Uj25p4+kkmJuBGTK
DkK6ynhhZGJXL/pM80yCOAvkXRqlNnEFtyVlYYpysx0LDhEXh3oQPeKvezlV
hXzZvtuK9pmYuTTGlsrl23pVvuev2ps1uZK+ro5jb2w/oPj6EEaJoal595at
V2bGMlBJO+eR1bI20aiOxjHtMpTODZLjuxFfeBZGCRWgyWu8BWvNvj2fRz1F
mp4uTxGkt8a/bMxwhu0ZJxtRVQeMR99nZNxYt1xkojyw2h0GX68j0RH8nn18
b/GQjsp4kIYcu2GtP3LluIPDEX/XJwFS5/JhrIIljW/8qOkEHKB2FIOdab3l
3tcI8fvnY0D5U/+TxpXOJIx7Y9FFxCqt9tBIqV64eLDmyatwoe/PqUNhbhOx
HHEdM7WuiMAZyl6XOPFAFx7TrIlM4Vju5GDZei1U9QL3TQ393i1TyWUWpUfW
1JX7TA3oBQTc+dP6pVok157MvvJoXUMtgETiHHNzh0JjSUQgf2+1SJeco8q3
KeOF5/dGd87V5mEzu7m1B3syexM/YUtiG4nhxuN1loL1X+ArPQfDG/srm6Ad
Xk9rjvheT29QqpUQBtQLnSUU8avI1RsJ6U1KwR0h6ob13vLP2ZxNhNQ6KXAK
ORdb5S4vVBw8DTctXLDVhsOWURHZtVkUn7uzcAJBbyO87caKQPGjYJdl5062
G3f8J/Zdq+lFGTJ1737+liidVUOjZ4d4N62NDaR+mqG6r+clV2b/3sODE9zJ
RHxn+rxr2YFBECqWjAVrH7ViJh09x2cYU1i6pgoHgBew6dsMYpv3zargXwwO
SbkD+kJLx6JkZQFB+fGLPm/gD1OD6wthUuObuFO7JW2DAEptxt3h8aAcCvQQ
wvcd+zkjKNnQ4y/cgWVO7tND/X2rqXs/ZC1n4O1xdZmzlGn2qq/Eal+X7FAZ
XLizt8tFSTjbqfirz8l51LF6sC23AwgiKUAfG/DfLPFCdlr0QWOsccobZ5ki
C132PWBlz4MF1D1XSjznT0KqrjOV9kbuGjS0d3i8gKaUolcEsUvghvYPqk10
KTPy6VXymCUchGok0eqYs2wF65Cg3bzDwzNzyMbujR0l14m0YPJ74mBZGqqH
skamsLe807n08MujYHqsaxSDbdomyGr/p1tBmnqfnW2rrwmO0cqZ0oOqyYOn
PF0GAg/THXuMN7RbUnOfZuHOJocoGV5K6kLg+icIJGWf2laTlgefknf8ZBVv
K6YMoHor3InV+/ZeDcgXz/RhcKfirtfci7xyKH1UMdyJy9EkJ/ALgnGpdUcP
dgmOArIIbJM9mmUUnlO24QsyfUQE6G8EHLBq3aQYwJmBtQCBWhg1JMzof3uq
VmisM5tHsV6cdi41oneF4RUNUilYNpMxJv/uyNqMxOQ9WfmV6UFMQF/VV1F+
5N1ZnIgZTimBv6aIiNIHF6/s0hyCZJNdFqDaYb6cyxKJ/e6oydjrLqNwZ+0c
4kdjNFh8VYcXr5WAGNOYCqSOvuWJi/RFCiL9aXVO+Fdlnv04HTsjlfn0pev7
eW+qd3AhZhCw2MV6b3XJ7n34IJTzBc4E5ho82/D/Ceu0xE59pexc7bbThnXV
fLuy+loiKs37iK9LipIZIvs3gFKdSQRmw0L9GmQYCAr6Z72JTXBi25V5CwHb
Y73dWFkP1QareiDdl7P1wkdIP6o63hq8H5d7pcmPGzIExkC3HA2Or16impj1
Znkmh8vbh8o/cxErc2Ye7InbHcQqhCxcsDJcn+P8aiQl+Q6w3rJRFwKQ16xh
9zGh1es04l1srwW7RtjXTSXuGXUmabnVXThq/N0TwzMMaU0jZx+9NSJOOaFa
srNQRvvX/U+4wKAUsTaWJP8/5hWYussjRqbYjGSu+W5nAhIU3MOPa1mTARHC
+ynCcRE0Ui5wpnmwdsy+BwhenyBcjSokEp7KfibKp0c8/WAaamog7k3fAHJC
zEtHIbhywZ4Cl5wgPVAebhMAkLtF1nllBeLAe69yUGnwCcxlckLNbVsrO3uJ
UFhTUsW7Bl+Uf3yz2moOuRf1XJ5ADbunDOp4VGCEoqoa/I0H46mVd2600uuA
4PEOsPY+ANpyGm6zE2GJ5YlQ1DJCBmMjuZ0CZUly8mYAfpCH8GgFpqMrOIES
sOXM7HmCiNVaCtN97OqAD8tOKqJQ1JORE/Crc0BHFweRBHWw81KZAb0mZFkw
cg9uGpY+AVyt1dv5slQKAlyAY26acWkPn54AtC/fjuCofTLVZFoIXqHqhlo5
8p9GS8fRzoP6a24bVbyiOOHfEyqn+XAGBXVZjNc2+LM/DwNANnwFqAY5O9Sh
O/ZnCluGx8xdX9nTj1JWGcpR+mXfIQJ14UCPqu11J++aURfFzcDCpyvTwEdH
gQZPhxDJSGQOlhcDYJgMSz9Qr8xyWw+xBA61FyaZauBn38rUPHZpydlrnG3O
CQMhNfG6Z1669EyIfvASulSHttVljp9bzTruOVBvp2Gj0pm3HljuhAYAQBMu
CRsX1c1MxJ1ABj2aWNnaVuVA+DA2yHlwsCa6kjMQRkWyphg/A8W6RxBqG6Lb
a9xKlsd5GJrStywIPme5D8PJDu8eFh2pZhwIhguqKpdvkbA4SjA8JZ2YP4cJ
VzgNCrR45ou/i7cKV+hAQCRxwqHUe7Gy1vt2RdCQQUCOSX5K3lR37PeHe2eB
FXw6ZbPTuBqFEJMSdoGPV9gvxEcfhfYcYZPEUgBQzI5Oq1vWb7MOmYtN8ne0
Wg8BwznHiR3I+LRV8cjPk6aa2ruhMUBveUArsd4nhwnbhpWY8cMOEGNn6suJ
Vo2Funm+BZqEY2o1XormUICfMnF2koaDp9n2RUhDcjzWJ2acpb3pyrs/1DEq
5/jAX2sVdjZpMSAFseD+EF6Hi0mS6vbAYmmZP9j7oJ/QBylzksrPoTyDziLg
hUm3OhFau04rb4SvyHsUZkb+6YewvbCHeOdzW7X6gT79bfy6I0q1OJFUxXR9
tVR94TV+++Hur0Gl4FLC67vAODiRgkiLP1TcviFjEwl+2ZM1oHkbT6xJA7WO
rogv9yuur9TKNaXYKJzHyIDuNmeU7Z1Ovuj08TgoLcnrJcs6aWf+OnPFCoTl
7vSg99/ig+kPTTILoeBgtkrmZigAkTPpI1HEAi/oILmhbbeMGUjVP2+YGVVU
P7ytcj0zSxux+csGbHgHCxAk4LQXHF874AD5alLtxfX0/1fdvxvMKtqs15SM
dKAP+R/cSdaxML5cn/jq7rErV9IRjd/52HB7S4/sCwKBluN9px8pbvk7/NT7
WOW+1F7c0UmoD+Lzo3LX8r1+Wpq7A7hg+7si9c2ZgHpjcotGl0dl6ZpRneM8
fQEsOPoji3qN4MvWdVX3kC+l5SFN1Hexs3Kn4hcgGtBYvLx1K6ePF0BnqT3w
Z60tfufEk25Ch2YLhtRMx8KaHTlClbyZ2OnqV8f9pjbDzfJa5ahQHRgyqdJQ
qo7oxU2X83YCG96b48Dc+Ui8Czor6mcHpS+OENy1Y9ouYRjGoxD+WwsLx98x
ViWfTtiDWI3p6/kD4+Lq5Sb35FOFJbDmBYuzoSp87G9uv7bG6N9jdGmJFYZq
RgsGU+tQntOllJuFfJLSD55hc5VDEO3KKVrQ2n+nCit5O4lmhid62ZUCYN5w
9GZxskGncF/+r7LPWuuu34TR8YWgBU6vCCtXTh9XmW4TGcVNU6dWWuxtkIMx
ArCSAaEh29Uj1OAnMb7wmOJEA3E/ipVdlAZnNuJHkdPLfBwSpRqG0tqdF6Zx
lLQTF6qICRM5FWFalpOiGfXNT0kiybF5UT1kQAITSS1J7W8px0NnLoGoEDHW
zZFcafKWsKQZQXxgh2k4rlK5+z7hlEK2gvYLtogDSi3mWwirQyen6uH+DtGS
2iRZrtXALBSVjWyDw5Kmm0nyqD1h8g+RUK3NbS81WCHzpO3dTNQTqMihanlx
1xzgxERB85rvvCrPji/ntNXWv38iTGBN+5puXakMxp6STqY1n5Xwok82NuXS
RQ7w3Lynyu4OMxCv1I5yp/tkDuqu/Mkaqz7TJqaCsfShzJRMywuf8O3fdOb1
5nwxn3Z9K5irWJWwogaELGApwjFiDOOE3o4KZvsrMTb0gsGcyzenSk/I9CbA
d+F2I59gkQrY3qS+EAGdYuKs6S98/dUU4fzAQGDHSvU+7a2h/Bb9W2m0T9xC
QMELCV63VcTZhaobvas454+Z3lXctEWZFss8Eg3YRL6mYRWN/kUFmH/eamdm
kz8kwecq/tbLLjj2SXIIaV61OX4CwQuAtj+lP5sNwO7WKQqsxZuQm982/hxS
sRN7D70AgtIU/aCAZ49oRiAFepbLc6FGyic/Y9EMqtzbuiRa2KO2VNG2Dxu7
fGfbgR8VkDAleySUxydiNUBFHkMBuo1IX2AevxS8Gy6D2BNH3dXyrBeLPp1n
pYwdOPHTXMomoMlC9Z3uIzsccJ5B9aMatDkhyf0gFDZeepPZZrvAJFLrjh8N
4vuLpx9sFTSE9Tsa/c8KHOU3ZbgEDbju9UFmwyC8hCzru8ixGJbC/JAjftqo
qi5tEIzw0qRTQGT6iHBOZoYTBIKZt9+PZcUuzWVFNrZqTjQbaRseKlPBIMBG
+o/52zq3csR27bNLMLpkKRQzCup5/t1YzXnBIpNqzpQq6ST9s4J05guRMLgv
2leY8twAIzSxX+pwNGUBtmQ9d1er9zmztI0WjC0wWVQdVXR+un5NN6nqb/gf
aHXVnurz8dH0HDnx7GMl9jqVr5swA3DF9AiRuYzMfOgA/1uExzj2hh8KS1OB
5aFrwN4fmlf/aPlN8zX/yan5UiEuPKXCfaYKmchF8N6lAMAiCqkowXrEhD+M
1iCkh5aBJeimvssPo8jsHyu3B5Zux2+2mOqfsBr484eQACYu4aTEm2Fgjc6k
Ha8tuzbjyXkK38AYep+wz/IIsACqB2SIXXbx4UxqxkdJ+JHA5gAwEkoowzUI
gmld+GAJAONbEX6VV+uinhsS+kFN/Ox9S9eupQTNOLqQEcTtel8RLGUCbKGk
NgI29DXkOm+dbJkdPhI5tU9ZIagWK8vlmAu8mftY98NUJhMMdiHo0HJ9CnaX
IWb0ehs6jymS5QoVH/BzjYG96JkR1BgloAg82QFrsRVZD4AAJ3iPkrBgLZBI
8CJ00tg2GrehOcSNAhqqcQSnjGtp5XqPmmkeETmWlMsHycWmETrLSeSpMfBT
aGLfRi5d/2pKcvssFl50S/DbGVDCE5p8epOsKRuW6xRPxY3k3xnJWZFOylY8
/8LDaQ8bhnDc3qNqj5Gu1SW2HYklfkKxdcshaerMQQ8pz63oYprQfy5bQC1P
yizQBrgW6c88un+XLYd65wIkEvXMPvnts5ds4aQQo/XglIz1zwtT5n13GZPA
PRynWGMOkoraXYUSYdjAZNAwk89/RzxY7xVx3YA4H+bgPbCMyHcsQma5gAd1
haFBbuC5AqJDZ+5m3QlDlD5n7C8nCosIB1sD+2aCk6GExGbdYG3xiDFyqI34
aQCMXHSanAwzfpP9EXCgqcsoRaPoA2LU5PcR/PsOP/L+xkv9sZ/78va4uyhL
eKhkQMP8CXDyO+cdBYNBK7m+wOUzKZNmGK8pDrKE+sbHfuhqAQvyzt1l3zST
KzmDO4PIisNyU0Y0rMe5/npREelRFzpUj6D2vkH6Q7izsWNSpGZ/pmYUWXUB
ZQ2HhJ8XU9UQT8VM1V6mLGuqnXVuvzkDiCCjqhdUbYImR0m36xE5lnedWu63
n2VSuSddFzbwwddu0raXqCLEHNp/1nF0GBlt/sQbyr+n7zLMEzmetQs6MYFj
J18cRwWJhYcdGLlY7HhTFlIUKtYXezJJ6GwnThULHgdEok3XWXb1G9pV++zr
gMqG+uvLtS9Xn+ddcsrliSFCw/z2WKjGi7SvK9TBQlSeePFr3lemxZuji9KJ
bPPnXELEwyaq30F0Sr9Ahh4coR80SOaWzseKsX5ta+ytGCkypIBLPRMjw6TM
NTTPPdSEzNFjcIHxLiJLgJSpMHvzFMmW08F3bt/3QVRI+L7bLTmHfwhAXNhb
MX+5A7CMjHeYBpY59mQEl6KqOxZ0o/JSc8nRRI5DobWGbK7w7S55raTmU3Rb
pSgpgOjq7P9MHCC95NP5BiE+J8+enSLZL5fgbPhpiduBdkLjxY8jbCDg3rbR
wEutxvtBNsbEuanEX0lN6IBjy1S8buFcHyPt8HeoJtNid2xVjnle9vYdwwzt
xHJBMeW2ia/AcNo5gdihXHIEcJkepKD3KjXZ4VrAmXL3e7fhn06fxbYHuZwf
3Ade37Z1OhjiQFW3m+YNRS1c6ZurNHnjZ2etZYp+FOHa0gX31dy42EjKVES0
5PC6S2Ec2e/qjIN2jo7StcWyBFsTWUBGZ5cPaszyK92yoOxCwwGD6u1Eqa4w
G7aqlSidd0/vUm3pkCZg74Imrjksg244k+0nW2OmtZWMB/z7sQCLkeSdCmAK
T3QZU2XnHsARH33Y8SOUJ9S8OOoIonQjtLwooBqY/S2It2Q0nDQiGJ7ToA7R
7dxQCmLyjwid6ru7gaaHVYnqekxG3NKmmiDqrT4QpsInifRmJk13BhV5P0B4
uQ+JlUyGcJGovENIW1w6xTUOkyPMT5DKikfBJ9Y/H6YMpDIr0LNUI7UWld5T
p3y43SegZALNWtPVTIF3TCxQT1JF7hGFmPlrjT2i2gtNtK0PL0slrZXLb7h7
eV4o3LQZhdNEU1kG/NZwgW7xmCuOxHJevcT98UDgMkgLt6weohuaFLR/bmYP
FG7V50CS7xKMwweBV+N8KvT+tcbY7Z6LzyJrKfL5y0sf2jPNbHtEN7U5yl2y
7A3E+sEeXNgyLU4AuBO1Y5veeJGsDrPsYAa0BdFADWZJM2USVkdNyaiyOOLP
p+j/tBWLWqwCs9pOL8VwgGueCDtgx1MKbGbaDkxsVY9P6jSTWH+X7AJ9boLO
+UzN78N/F8Mo8KixNYiMQ2/zJqv4gyLQShbRfD13J2JBlXnOq2kEXbMKnTHF
9DWw100jV9zyIahBtyOIOF/UUDXYmAPswpNbQeGJaQSHsRtKAp9ngSUa1mkn
VBaYq6yv+w9+Q6euPn7EDV/Far5YFAPH9wunJK2J3B95GpNLlh/pL+4JZR2S
ob+XISZ7U57S+qFgQEuZZM9G/XqTJ2ZCb2tU4usz/eFe8t++b4NpG1euFHsQ
p3ElbslN0/mPwI7/RLi3S6n5HFam9Ny65NN1yTi8YGT5f8khIA0CQeCiLujP
9PHbkhGtpe874Sw9YUNCv54wssq/6ipVi760uVUwRhQ+aLOnKqag+8WPPueV
+Jm33Asa89QPAhfGYXFLDeMXpe29E1kPF0y95VLLxTidXG54ulDuZ7G0O80+
uObAzMcQlxcOw/xaX0GHd1co378EYAXLIylsdsJvmx+4L+x8F44xO2gf6fOA
aUp8AUCKLot/NUSVmov9YVMkHo+Lnhd8yG7NA6ilBYjdHRyRdKBa2qTxNVhH
obNMggZPFmChx97CNHEvY8wvaJl2omE4r/NKsMFnz9K1pTl62bPgZXMAS7FQ
bH87UEJEWNfhVe8Djl+D1pwg3UCK4NKCCD+yZp7gK1CoZzSm5SkFkl1jeZ0I
n8fpabHBFrcNIz+sgugo6MLTehTXRHX1jTP0QHV+pS2JrwXTbiQr24Lwekd8
WTs3dupGXnkhai7d+qfUaH8INWviMochMqUYlptCHVOf9OcaY5gaTT3ysJPX
m+YmI6bb553YUBoVuk5zDPbBzFhnAqEfOZ9ZvZjkyI/hnPKQcBIpeTamvsjo
TQ3naYo8jnfEUt/lVQsP2S7dhWjQ9F13gJUNhgrDXdczuWnYat7nX/NEYygk
cu+y9VF0wF06E4dGWbyy6HRznvQkot0VAiQletPslXm9d8rzeWZqxMzCXuGF
xwY52TGvNjezeGieuxUWVLXg8esmg1/GVqNIqzHsvPf219Wj6GGzFt/h8w2u
Nn6CMRIvOc72mNkKJwOT5P0frt4zGCl86hDyVWOctmUCMFITsYVLe1Wik7iP
Kos10fYYBlMkgHWu+13TNBsp2zPGl8v1lBRXoihH+VxosiKDfzqqTg8nqMKa
/cpqzDpoOnWQdMqN6uPUXOcXUcTWs8/W5VAZebq5u/9WZvpNVcVPcYRc10X3
G+zQlGQSIBNMeWVZffFdZrqMwurfJLplm/Q7PhIRU3HHMlV/msFKuVf5hG4U
HJ0z6u8Kr/iZsTvhcBHWjtJemBEppJKL5dfXn0jQh4QNam9gc1b7j4K+yKSJ
L+LoGufogZOTRs5OVcW4TJ0TiL/r7Ot4YgUhJy7txOVatMJDE/7CNY723Psb
o/XFcROwuGdRh4HWhD4SVOE9Tqj0dxgXTDv3oqWEzt/hAXymKy70Nem70Pl0
5B/Tbwj92wf5cRT7l61SbNqJgIvJ6j/H+fMHTSwm4jNkkXAyKF24HV8h2otj
r2GVduuLxyFDv77kecKFPhP5wDVPmsM1GHAODA+VNm2pIZ2TCFJGv8yqbB9N
2OfC8LVnGPOAEQVQYPt2Pxk9xZBBw3EdHvO0QF80O85q4bscXMwae16bQ9Mc
idqbPxDOSxehYNmuT0fVIKWUNC9ViJ52DrXL1vq5M5x1AJFh4+9AAsCFmohy
WFPuwurF4GxXInR9Ez1+dhiFBcpiZi5mZ2dlfpgRupFKdkKT6QdXM02wFM80
TuSwXTpAeKSpYYZfItODLHMME1I8h2/keEkiK63cJ8sDIoI6oz8CCcrACyBo
uG/EBSAfPw8JJqz7ao09oAqkKCznZ+5CJ2d6xw9zpI/Ypf3xKRFUyHHZW/Q1
CxoE8V/F34DhIzvF8mUB5Pxv/fyxTsyM/BrfElLoZJhTBp68jKcZpdofG+7V
EhLFECyKLNRYTAS6/LY6ePfXWrz6ysnui4V1oT62MFVyVRxLJZgcR+aHzWmP
yc+Gm56G446Lj3/8odTVmWm+Yk+AGNyJ1E7TMJu8DirbJltBX652pLeVUTCX
zqCatGAwBYbUDVFMEF7BKro77WSk6jskmv/+5mb4GnXj44gobC2hyG66nAcc
pY2FrsyvYAeENsPdf8yslMbcMsRSKUmQkZ96C4WMLLCGhTxgX56Fu3Tlwvsa
uOXRn+06q1b4drWF9SfJ07cKqHSZHiTTOl1YUmfmI9mH26wWNLmIhV6+k9Re
4aBMVFpXs6QubzQTrBI8XT/BYiZSeXakisbgol6/7eano1P9uuJ3OhCIoatM
skJsJOoVey2IttFNUcR8HRChvdtwGSO985FZtEeXVE9iJQvfcOhQF7MFsFYA
9mY3E2U16DXH6XjrGHRE/tfXEJMx1tU2izOK6JNBZIix82ceH428hspKyz2s
tzJu2Jwn1DnN/edcMjkWZDSpk2obx6HZvUapoUdpHkhPpFKaFa79qe7t/x1O
ctDMwP9xn1wakKG16666nOGFnBnh8PDms3VHpzvPUXtY1uB261Q6secmIbdH
9lO0TWTgcEZVFkT0OmP25YXUVzV/UZ2Eyp7umXx2gAr1Pt7p5Y2r5zhYAaPb
XkhFcihPqDRYNzIpi6O4iNZ7t3Tamnuz57/CVqOyJzwO4P911cdiAMl2iJAa
44aA9VQ/rH4aLzYVRBtdtemt9onG8HMdqkvjjz+f5VTkNKJu2+5ujlvCiekU
ZEA1N5GDuqZ+fTWAxldulUBVipY4SZehDMQkpqe8tBFzvHUQxMSjs24QQVM7
DTuoX6ontYpzp/oRsjgsmSIMLThWvsDJiY03+KCHOQaJaXytOmtgOVzh/Fg8
zYcgqvfsJHRSjGR8vLP53V0ZiWZ+kzti5wPNPOEuiwTXpHJd1KzscDyN7BGr
MhITqWEaw/lJLuIsfEWDiImhAOwfemeXWjswayLALkjOBJLffEMUR2bNnaPe
yVgWHQOuOXddDw9gBrM3kFIMQ86pUmwheD5z8i9nZUMW+l6bIBwHpSwMBz2O
tAvur5MRGDT0Ovnsmu88fYz0FWzhRpNlM728c28kKA6FIhLuKCiNVx9QSroy
hP05l8erDNNs34bn/vntB0DpC8BY4GnBCRAOKUkSlyBGm3YugtEJIrAMTPSu
UG0zwQoJMWq/NxEQmfMHK1CnTDp8LaMj2g/IPuu7s55JlMW/us3cwnspkH0P
M51HjyoilSYCRKmxLZOe54rDCoCx+8l1Zp3i9hblvjToYFziRnWskqC7QGr/
0rkQC0IucUA2ziOoXjvr9N0qHjY4brhDYjDOBDurJ73QxS+UZ67SOH+ybXKk
IM254lJNocuo2AkaKM3IIwnGDZWSA744KOp5SGdzT+ASk05NygBtR3H8FtyH
MrXkEMvsnboE23km9dT6knh4rOma3y99WPG/LcKrwWVND066OaFcOrxXmiL5
a0se9aSgjSLoZu9/fO8pju5bIBbOCgyiGCRmqBsXfrzuoW2ihIlr4uHpWqu8
FROs1t1NHybcIhUvU+1FVyw4eskuoQvdpzOWBWAHb+FMvTB36e8a94DozmMI
GPnjUoRBXuH6PCF6hk1icSDjAnzStICJakqORpoOijYq/AJdNXScllYtqGKo
GxFOIxa8DY3DbFzPCAB20qgTVOZ9xk7SDR+6+iW99rVxep5mgUjiPXHuaM4G
Iz+6W+ALeLg9XCpPo7e3AUqGhmidzcUWtSJDW8bTUYIpvNVyhyvE3ua8nRsg
h6i3t3KOVijfmvUb1FjKHkMioBaSGkTFkVFUg+Z2n+NAsVshQBq5DpWiJUkH
3R6YvtI5l/sv86iSdUIVo5YCGb8afs2KeH2SE9cYt7Y5ewC0j7bB9L3EFeG0
BA92DKJt9tJuoLGUDcL4ul5Oqaqm8Dn7GUU80os3zpmeGXvMJnYV81vY+jhg
BQ4CQfQF/HtBeK5WQksqy28pNR/wNBeZnsY8EMnN33djtGNwsQ+udPXlwLTb
M3Ewv9Y64KBMMlzPhpB+yd6zDgWPLWdaMqZLnUE4iwAFqN98os6i/9nNODtD
w84gc2O3uSuvQZlsv7R+D+hwZFt2koJKqg9BzNBj4XTUe4UUzgPyGLUA86cl
++APITMr6pqV3Y+4is0/OZQnNqW6K7xqemMQPIOHDJIVbQ6ZhXKgZqT7afnC
hyaeyKjHT9+8sJrDjUCfzZSZ6tAMNomPwu1iIG9WCu0ASXjyGDG8KvDLazeR
9CuMzV0d58lTsmEqBnraJWyCHGT6gWLoefg/u101mdivAbwmq8+yRXu3EA4r
JuKmtbJdQaHaCNttCsG1mMgTz71x8CP/O/bMFlY0RhKTNwV/vkHW/x4k4UoG
A027Mx+oD0vNRtQIdC9WykZ26yOYR4Og77b34KFfLdlFvroC8qSjMlTYcWbA
f4+kXiUy06YELvHhv0iJ4FyPSEKhLrHdqfb9Ma5VMsNHmFcaiXk3GbGYhwAa
8nM+v/sNeGDeDhys9DhCHUD1bLuoEXCd1kpWB4r/kjkiR8wg2cWXnhcdFczf
LHwNKbehb8xAMbHpyFI6miwLDDZm+H0nsoftPpJtqTa52VmJXhWh3tBl/ECw
b4c+FOCHiJK/DXQloUNpKWm+UQ3o4Gsmyu/4W7w7IFvuckETR8SXuA4bBOoG
u3+G8FB2AFDfpFW+2dW/iU7qxGQ3460iia22ckF2dy+/t3lbZcomNbur/FvP
gqGDdlHwZdnjVR1FkEs3MT+vdXe3m39KODPadNg0UmNd0y5zW8aGf4cvmur8
/c75KO+3O30jIIYMooQWccAGXC4m9zHwEIa00nb8i/vHKXSXQWbtkOWlghwF
gui9VO+ow5XBOw+6U+AcZufX75clmaNQXAUJFQsUSPJZUGlPra2Gq5F0JeQV
VUzcDuLjoybd5Daxyn2KlLPN2beP3trxCI4qA1jQpPTwBr5ONttn0U+zDl+6
Dm1FKFWwZz+oSswoI5AE4ooBZZB7zed1QGpu34IXgGY2O/W835TvgrlHpGvL
vAgQUelauYuJAg+EL3zHirjtr5N2suixhLRtDDLPSrL4XU0KJJbYy0E3RoLH
+qtn/oZeiX+1ERgovjYN4Lc1UVXHNbJQmDJVYMfnogIvTtW/prHkRJ33Zz1s
jUaVutq+7C/9GRjufKp8szU1Swj0nPsnErYFXAfsNYVN5ZEv3z/3xKPexJd2
9sO05OrwM3Y9FZiODx7aTirj+QIHfXb0UayoQH9Ve+S2/rra7ZrVP8e5QSBn
+1jpaKvmlkhb3QXwpFDtHoIrzPvSyfFnJZUmlcEXJYBMhele+LOsiczdAGxK
Imup5defeGQCBzAXPgUjDPNDTmM2dMHPPyFDDrpwjvafavI85eisJZBeoZjI
3+VAJ9nAKv79CCDtvGUAa0XxvuqSKargbE0uZnCNSu6ryMdnxPR5W4h0tVDS
cXMq0LIdbnwTbMwC0U3S+ai7BkFDDdRDF2pmqNtHwsmMarT/mQs9vVeEgnpC
/dS2iWVzcZNM3tVm8mNL3VbN5S8sRLkqtiwksTzSRNp94+35adx6oT0YN9Dq
c29gXDd3ji8qFYKjGZl2aM0oHGwzxct/YV44dnXp/17CXuStVfP8MJt+iyrA
oM9U5JNKFu4nbTfB35eEdwZP6PNTb8N9lHBV7zPyKx4lzeDyK2/PjJRnEFB7
ozH41oQJGEuHAtbneNObje82PtKOgByu8RC4t2v3/Yt32SzMCptTvqkLKTAt
B+EVZAv/2Ttx3+gnaJ4Jj3goGppkvh8QQZXn5yF/9E+sjNd0zMcI5N3WDJIR
T9NAwJLIBTsz+RfbPToORZNosU6bnfaTiCzd9Thr/Sy/y/5jIQxVGmisYVZv
OZl9ak3or5wDznDKuTh5g5j7ysi6q7/EoSf+6Mcr8YuFOjIyYgkcermdAymP
FuORT1x4lPT14alRm6e4QL+jAiPId0gxUUgS+XpA4ygeZ/RarX9UOSQ99qe1
74aSF9FX+FfwGdp3pzp7Z3eoBgAGhly4anynFnHggCfNZ+ax8K+5jnSlh4XB
4EULDQO3JYGyB+UE+OS5VI2dfMoUUUlwAw0OlV5E2A+ft1vj0iCmJpeg33Sf
EL3jski25gEXEm4pvAdEj3cURQpa0Er/dMJ2S+UAyw7ICaQpFb6i7J0X2EmE
3d9rvt9iUqmo/sF9Tyk+dIN9D26eJQmMauFAu+K5TBAZs2aithnShhko2G4N
7E/bayksbHGDvFqe7FQi+uvmEdudZo2uZzue5aYHZ63UDIZcNxRw92ZWkRlV
xA4FewjsRKOH4HUpNRJj8Uoc8Y8YIBiOvHTnTgkUQGoWZDlp/BTBjL999gBg
y4tipkxGV42cGhW2yOODrvsggWlreS7SsFj6OtmggH09ZsEr5RCrOIugMyNU
BMDtzEHgQJOiYJmaX4EB9uSGeueCXRyDZDCMjly3+vLuYBd6/4uLGpBw6A7b
kQYw1wt9NqfD5gXxRcny1x6Evb/R3zpmkFtQD/FjCoaVo/3DtYT90NcyYYNB
e3Hf5DG9dnitU4qgP1h3qkcLfTYvFfi7jzobYWvJnGIxvTIPnB2+EuR9YNy1
cm82vsLkffT5PG8g1gzD47ktER6woBwfaSbAaBNrkMparo/CH1WSqKNoMmUU
y7zE69OXYaKUOHAzN9mbmEvdQWbagpV3x9rWFW/A0Ev45Bvpp8kxGAmLaZY/
32E+EQuBPb4Rs5k+hq3krk4MW+9LvsLBV8H5FH57CiTNyH/7axzUn3nJT3fi
l8UlJ1bLhvxP4+wjhPRFw3Ugi5INPK0CAPTLFK3PJa6N5pM+nqg2jLtc4HGl
WS1PCZ/mcRYhOxJI4aC+emgd6Fpj5YBF8f3OprJkI9mCqYbxvuvmsFSNg4Gf
low0ZM/Y5lzTF3GW52JDb3nQ7wgr5WHk//u65vlG+aC6XpUJu6z6/SZh8TtZ
a4aBoS6ooD8TIkWBAsLVVAgcyoxnx1f6P8UsPS2+6yOvMtXd6LCU0+26tZHG
bI/gDUWewQ1jCsjPmB4o93cxsxiImd0AnXYhG5841FTCvIwZYJDbdCPV7yOz
I8AdXPWrmbM3VYYY+6FXCd5H4SlxEPJFIY4RA3r8tTm3v3iqVb2yQrEJ4iSm
+r6DWQ2gOa8XmODJ+6rDZr0DER+yH9lvIUwLl5/8/OCx2G4YqlLPRMGLW2Vr
AxpDTINANt9uDCTo011rfcNVDvJ8LNgEt/0rzhRbBrpW6eDhfGWpkxUPjUzC
Ug6/pyjc8dikBeq9Pkdk9zFosgM8w+q/nJj1OP84fqv0lrpV5SjDBSnv9c58
7XsX0yJ4Qzzx0kL9FWj8rVBQNbmODQCIRUp6cueXHQySM9V9us6pm9ZucWQc
pJkK9WxsgqBePAJnw3e5NR3mlGidEVByqW7fySbCnamU7iXLBnFAbqlsHRyG
i4P2fNeq+XaebAG6v0W+P79CBzLYHKxHYAnVr10tu+LeCzxwuCKtuClAtmL1
QdMxw1kVcNJqUoCjpcwkaVomv9iwAgMBdw57XcAuTklKNqElcL9intLj37Or
KkgPuHOk2KYLvX6Z4PYI398oeV4t28HgDWKpMgpqtX71PhQ9apasOLB7DHcM
ITscozRMxaH2PyykB8M3C7t5CX3Ra9YjsXzvMShYLZ7/CtbDNiJwNZmFYHaE
Uwld+jSb6S7GG+neS3RHOZjiyweUlcVpXLVgKeMTrWAiuEYmyzjnv2m0i+MZ
0mNRCC03uinjIrecm5I5WDfO8tVUEfjLY7JJQvHYYsOh3Kq1H8U3DjiTHBwf
3NwGwmQtcDpuW1xfFgYWLceo5uwsBUHMMVT8gW85oPiuT9pU0n2qYsYJ1O1n
EOl4ZBJdvbVza2dHNURQ/kXbDqQQBF9QIlWx4U7cgGAY9stmNQaphwpCyVtU
UmSy2OKMqAX68FI/PMcIU6m7j6SL5HKA6z4AV7PZsowXwO0Iy2YFJcuPEOgC
S+tRLA5stKOpQ+Z4Tws9k0H6FKK9MNOMkmJJ/kYQZR0sViSyGQkLZBycNsd4
XvHzFx4ZK2Ro/poHkFKtnqNE8cnJ5lVqcGKe+blXBORBDhIPrO/tH5XITx0B
7j109VteoWCeh7u2hNoXoW1LlHgsSmSW5B76yClHogD8Ksl9ESVwExkX3v87
YBniiWz6VJ5MMGHMTbGm9rXw65AkvYk0SmcFqKh1STULlj3pHyF9FL4Q/T/g
f8cWV5Xki8K3MxGFiOP4SgNRyOj3yAgxBQdpA0MVemV0wvk5RqowhFBbZ2HL
1oSu/8fzFeHFpPJxyrHfIxaWyiOuLBGQ9ZS/ArKEURbhKqzTPMMTc42TaVdf
PdN4WSFJutejM+pzTQ4fFHa1V7lr2aCDrmkqzbM/xOVvzBnFGTBy1eLbzIIL
AkYYjLthsUVVsEIsaNi47z7htrF3cTSA4GMsLqiAtD0hz0hGMV2kj61Spgy6
tj7MBD1M7Gug2xxZp9qEjihKPGSdOD72ZIxRMWfyRgMPBPosFXqXhZOQdg8U
6fQKKEp/t4yXK2fKu7nw3SK+5oO4+vNibENuHt6MedTwnma9DCPK0tXCWRtv
h39oTaPcYrWLqcIaL2ddEUAiJdeMv3Rc5XYKUz2jfoXc+oF94j4nH16lruu9
zR3L9Wj4dnOI72ITo0CDRlAMki7V2WQUQ5B88KAU1wuZRe1YP1OlNYgs/z+X
YHqxthbETAyurruZJxNIw5OlLMFeg0rekWB03D28Rc1YaYIhw1bjwli6EMDf
+GnMv6a/36SXWeYtbHp7HGMDgxEt345eihRWOoqbvyRfLJIfMuYDIlbqj6ej
EfcAuw+6Dt7zZ548nK/6KbwBy5BcLd17bFO+1lU5DJJha2w6OpuLaLUHPTuS
6GDNXUwlFNrJiXH4EcaSpBMVMTO71P0fZc5y4v2Y8DLOJ1Zg/2BUzDA8Jjra
X3QjLFb8vmy8tZxKOsiwwnJNmke8+mAUvd9aYiDur9Axeje+Itxp553t7HAv
IKbHx2FEXchVOsvrXJpfWPYdGpwnTXU2Gdaq7EpZix79/QUfMimwadp0SbcK
nWldRra5TO/b+zUKydfdw+KxXTljN2g2i12PWxaaLLjerHLjDX4GFVP/X7z8
tN89uhOdywXY1XU7bryD0klN0rczXyFhoTpmm4y0C+0ue/2oC+zM0PE2NMsc
MYC4LXHPYSp9+OOkyifckXg51bA2BS2Uhy1EMit4LVAWhmh9NvYdnkokBISC
3eWOgQuIIpDkte20x/+JV8+GPELGZ2ckEfm2esU9CV7MCGBk5sMeo6yZrZ+g
+I6x3INp926h5F0KkgcCa8XKOBJVoDLbqi2iJR8b1T3ruY1Ce1ucZljgepO0
rOr68UEPCaF1CzTusmK8iRMm0BVfQ7SmNQPSY8P3Luhup/OQUldX2SLiFfTK
NhHb9bKM3xgRuPPQGRLXeVxgrd7CBxqMEXZssY9yWjBlRtbcimboRMNNLWdS
xXKyrClxYJKpAgyr6LlbqCC4DDhzra0nxyD1R40CXBaHKYKdtI54NuEUJwhN
GedDl2ugX9M67BZVxYsoMcD0cL8Ksw6mdch/bUxsz3Y5i2PnFZSbfJW7nCe/
d120eBQVwe2AQY70bEE0xg5RQLItfkLFt/NqtobpTQGIQqGcbteSlK5ywi/z
vORDxHvBMqMQyFc/JEVXCOT6oFn3uA8paz3UE4bvm1ZR/vABzZgw2p6YQmgX
I2vC8uxvKPmt2WXQcw/JyaRrFOf1jO2AbBD3XpFXiq0XOmRpBpGQum3jyA+J
Y6AMW0c6+B02AIR9ifBrZj4kzK98oTuO59LCiNZyi64TYO6ydo1zowVqwveG
aR9uJNe+eVCC9RY586i8/mqYWBliWerWwF0FOm4VSFvTwfVhWMiUq1wRoftC
m4+z+CjlemKt8Arg88JnbFK05816O4xvgCRvF3zA7HAEUxJEzPFRuV3kivQm
YnjZQBYYCeOmKfNmYmp4lcfEqV8pG/BiRz490bqFsMG1u2MVDVqHG8yn70yh
Z2C6H7BjBF5l0CGmsTMLxJas1FOGagQkk1Gij2h8f33PLTl5vXxKZ9vVdzeV
AdfuevWV8FVtBSh1W08f63zz0mQLXgm8im9x0+QAkByZjrahfFaliIiRFNJg
+nJ3MIpkBZBiTSpYyCt/KcDclmNwBsIicZo7YZbumc17OQilRnY14LXVjYu8
wm53O9JFTQiRFxx1chu3R/Z/HXoy9T9Ss7r4xy5jKrghB2WNO0qp7sbp+hqL
hbWNH6Itsy1iwsPPRDPkyhCO37VWMIWxwzZTFKJGQ/norpAqkLgDdYJ2KTL3
LJaAwcJdNlNRSKxj07nXXMlMNPT34zUyrGHoWiLA/NQrNUk0tBGyS+G/cM6O
bgN6FeQ1yiZL9tYSZilJPALZzXElioBkpQQ4xbI1cH6zF+TXjxDVskiowAMu
rulAuuX4b1qYvR/iixb/V5U00J+6nKEb6CwTNfKvBdvSNsF1oFtNGgrgdPcg
TQoe4FS4sW1fNJO2joj819FX6vOA2sXjW4xj8bPq+Oq0/jOmBbbzpWAYd0r8
NItxy/zCZnHbt/lgdPX2e6wEFz2I8JKpvLeVZVbGzG++9ysRm4CdsLNtWbnG
N+8BaExAMk035OVfG/owg7gcyGvq8WY6Yj1274R594/EAUbLXSWsVjxJ7MVx
iYii6i3fpCjmt/4SLkWxRg5tQTXEMEhXvcjQBdJf/MuBRpEnUjKd1cl/Yl6y
r0RgdpUyVbr1BceyvKnDD6mcj4wxIqDHu2ddkP77IFgppAdBfdIeYX1bFED2
e/llDy+Ge4hWuH0dWqkJElrtmAyY0yukIqNH7wcEgn2zLhY4Xy6iKob3eL0j
iky0SBAYDZ1004HLdFGEcP05LcLctFIOgwxOzTqjB6wP7DQ7i4WaWNbDZcIe
/5Sz5SYmlBmxgX5/x7EfjnH9QoTX4Yzs0cBoG5bXbRTiDoAjokf1i5YFbCJj
N/cDVa3ED3IYqldE4CDqbe5vi8z1hrOr+jygM1XW69BQZRUvL8VyPsAraOv2
8ivFKnGMp9LjEkn2FAERCK+cZcU3XE46TL5y5hLad4RIjdeLelLivPH8u3kD
V3Qya3GXvUZ2mDCSDGRmj6U4/pYmLXtAMRnNEA+zDfeZ5BMpUFyUj3Ko0W61
VKmBzI3rZFMNl4JVZ9DmNTTNjM2vYbEU1kMHSnbB3VPu/x9WbfXuo0CwBSZz
xa77PDjMh8q1jXCS0JUvjUaItr6V2Ca0/FCefGN9aExOUMfR/pamQx1JeEM2
zx47P9kBKzfDOst+uKUj8mSit4K8C8HCG0ghCqz1Nf+w4f2Jn0XQe6ernUS1
lfz64vH+NimButIpvkWaS7wRTFcQQz/jPSqUeZwwpJs/GprqCyB4KCtn8FIy
lTOJhKLTpahBw3Pj8ZW3tIKqbiZkCWMB9a42dGUp9kLAfE0tryHDqeObf016
NT+Z16/j8q2MUydl6nOfhRnFO7Ph2ZctWX3TzPvAOv4CJQcJ8xhnKH3T7QJZ
4xls7LCQTaZd4AMDrop04d3zDvH4iSVxcI93uHCUKNsnDvof9rGwTu3Iw+Il
+69m2fJ5ZBp1TL6Tc/EiAQLNwPMtT+Y0elZiJNZYliWJZT3Yhi72vY4jZ8Qf
ZYEgW6/E2YHYC5zHps6a+KTLhVbXWmFkUMvX6InvYLCkerlaj9hmBDgHs9kR
YoxKRspFv1CeNSv9EamnyeAYRFvpoV2bpmi7vZTxQwCrMSrGCAnN4HDjoaJj
AdXUi6C5z88Br7dNrQh3TzCJqTHUfpAs0pDIN5RpY+z4jJU4VHGLYQwk30P+
+mwxN07iM/TrmGQT1GgqK0Cxg/o4LGKxSVHTOieD9V7gLLaVhzqK3AivTQ2n
vSfyb0V2BKt0U1ojKYBHE85NxF95MA3kjV/vh/JpNY9WsfaUwlmsVYh6hrSm
XhXASi3zfvQy0NwW8vwtmLc8QWcutxNSq+mA6zqMM2SkxuS3r5HGVWkyU9RG
mn8/pCre+xGyFtq9QzIDgJq63FtpICyDekZW22j1kMiIlC+MV2L/4IOd4kHB
GPLtP0ZSVydD0QCJkL+Ul4w95bRub4nWzaP+BArGfi7bywwowJ38uQCKNeE6
JKAyqEZ/AgOTlm/se1DsX68GLN4pNIfqrKwc8/hSx6LeJakfomA9Qdph+rhh
igOBJBO+7X9y3KC3/YNVLlUs32iCS3nbiEVWNGJcyMfvZoGHwhqkoL/S7S4U
TIVIuA/NhJ5mtmWGrkpCcgORMuLru6S0ZGmoPuqBOR0zjf/Ks6CBUILGI5Ro
g8IY/fji9WyyRgpr4W8X9XGe7y2Z8zKH2Hc2NroMcTUP6R9NIvJRlH3b5Ue5
h5l8E7xqoNtMnQ3YWkxYP6K2F64BSX6RZojDZHfFVOtw/92+1PQNMAk5QrmM
ktTTT7FnEh9ftrBG9GgcYOPEG2epYRfFn+h0m9Uw4s+TeKnv41c9wBt2YaFY
9TQQQ+NJINRHIaVP1+nBCVDDLMuJN027pSl9u8JSY7fNxsdOf3qwNVw1YJ/9
yneHM+ulzLBWGTC4xsoEnCbMWIZJ7NGlwO1jKGU77lMr0kjAK0KFFW3nvcWo
rO87pqoY/0Dkt4xj8q69oA0DQaFgch3O//0Kmlv0rjBcDMiitAoAG+y3lPhW
bw/mbOcNZG+MBMW66/R7rCHBFkOvnQV630FT/uAFg/vzPPRQrVXdQeJhdzuQ
Eq/4jSrv/BGQt2uRKBvKjBWJwXgbrSakiWbidHcp3HY5446JWcVWYyN94B6o
7RPRUL+LojOFDtuGZ1R7RZVyeKdZjCSoZQhgHA+DVmihF5IFeMPCTIfob0Q9
09SNhJRNNKz6OyfRwen4KaKze5yDBgn/a5uiERVrGA1VXPHLjCnQNYUTaC4f
5Gq4pxU9YElhKgMOwJU/BILT0PMrPC/J7TCuAr0k/xiYo/t7m7dnJkdykzPZ
2a/Q/L2WxfyI5RlcDt8IXQ+KZzeGLPKbpE0/PfKFmyIogVwYMgDjFdY1JT5t
enFY7UCJAppeDnra9Kw5RUrD0HYPn48brdmxB8LejdszRKZnoBg01qZ165e9
Lja0Eec/LtXgABQV9X/qJrKy3FxLehfuMivYzonO5iKZRApE/yG+r22Ph8aD
GrcJlefM+7aybIuGzzgAX/k7lOP/rARRqLVgQF2pAoCgHa5mvOHyv/6LgEMR
o87yn/lfiel2QExIM08uNH5Uu0/iZ4VtXkhsuHkhWwnPQLVSAVUQ4hzxdvby
xfl70X8DRpIdxOQK2x3Kh6A1QXx3cRsdd7HjaB7rwcrQ0oZETAy5Kx4BpAqz
+fSTtAZCMekyz2MwI2qifkB+5IFWa6jSm3Ck4JU3qoQP+mRgtb6+be5v3/p8
xB+W5A5wJf1oxqHInsgFyiqgs36von1uuzq9DYGtIaltKSSyV4SN3h0SqIMq
SU3zhnSHL9Sy9mbU0ivQRCbtnCL918NQ7cHFUOz4H9xJ2timK318YHBz+nyz
XAZApcyQdtFjYcdv5kTJtsMOuv2E9/Qflo7Hod+VwgovpmADK0UrfB8RM8LF
5vYGgnJoDIPjl2BSLLuRNmmrBYJzVA3L1zNhsRd0vYr7+Wh7oMOpH3Ca1iFH
Afujyr5KmWKAOZAItmJF56DY9m3oFAvmBncARKKIlbo2I6hrKPRdVIvsH9hk
rLyqS1HDCcLtCJelZFH5P3VJaMQQjvsyPJ8oIWudJzlHdZlzL/lPxn/Kk1RO
P+yajrBDoMpLG/2SIClWihErP7f1eKfpDrzrWdNQbxyZk570c9tsiAM+5Yo0
E7L6RwM5ENdEFH5N2KzC1VbJDmwsf2yl7r0mcX2n1llJ4pTzWn0I9QvVjBgr
hmLsndYDylZLGhwM+f0e579ppjIH1trwhlvNlZ1hQZ4Ml8Wn2vtZzEkUpgh8
Q60HLGcbbAi0qPxMYyAOAJm6ttEC5GgxHw2l5FdrpiHtWWnJRYYCy7rtFoGU
qv7flD2AjhM69evrUBlMTW83NL66sAibeQjFSCnUCdo8swgHn6dvMWpNlsnQ
N8s9y3ioArQRWJpipqHZ5DipNMjUlv3/Dx+UeWrgVu794q70u6C5d/g69bZT
hHMgan39WKSvxyzbtViF8eXG2OsINCoEbPi6vi561c6nUhz+8ZlzotrJRtGq
TLuyHeYmEQM6FRwB0gMZNZ9x2fczM6OAXVK0o6fxItFBOATQAv4kPYzLsEI2
uGEq9Y15k8PssuDkVsdzrN+ASNmUUZ4SOLSjX0lwvaxmC6YXTLilwBsjYyUF
S9ADFukqtcutYJyTKWGSOkcoFYO8es2G9AqY6xQ4fdrSqzxzJeONd2HQlHmQ
1DAXhFw5ilFh3IAdiW1j10R4pTuur8bMEoxcziSjXBaGOZuFKAUxYAhwG13I
CBizJ5YpoQc1zmGxwxqJ2ccJ2N2ii0VyMNQJi6XHa36eGEW6A9lm2FObFPUR
B2AZShYq+/jqC7EU3cmrpQL3K52/l6KLj8hpYultWvBcyE17IaJcBf0q+yWM
hsdIkWtUgyrVximP31r/R82mWI6JZSBZjJ1q9Riw0GTzbmDLNUq1UI4IQTey
NMXx6F5TXGrn8wOoYPGumRyhoGJ+Gye+4rbDIT8AjeX3EQwLLD2Yj+cMvQaf
3ZdZa9P3LMWvZP4qvvyq9sicjOWkVbhfZMpq4eLo91q10gKx8XzDuBJz/O7m
1/Y3Alvq7EyKx4l8FYEE15T0LV6+jFGY6BX8RHqFQ4PVgCAZvS0KVt6ju5fM
UrYWGM/fxNjUAXkFrANloqaQ/3iIkzAtuMs4E8/SnkfeVZVkR5ayphx6vE/6
ioRf3tGFwlb0ROA3lgiuX+vzN5/PHuQUXRjfOX0fIkQotc2GnGC5INDHfAex
euAMPhurhwuzeq8FcVFTOYJcCC5pKM9kdauXUyzDH5RwDvMjvymikBGRqCeF
YAzL1jw8u1v2Cx25bK7UkTJAAhWdIb3984z5eSQuaz7y4FXNxLVM8Hccb2ph
cAi1DPRucrOWQsyUiDqGsA2K1/b5A22KHpCjQd7PwoqiLF6gvU/DAXxUIY1N
n0BsXpctiA81XkZL9zl6jTTMa2/USpBWmoEXXqHkQLG72hCDgG833RfGuzaO
/+olVQl2uG0SkvbPdgrLCAUniJCKcmG7Z4v9xfYXC0mFpbonhDbMuKs2fr3/
IlO+GYxjzUrITlS+5MrE998L9Wi9Nh0Y2+3CAuxFy/Ak9tHUnya5TVuMSq+a
oZgTX5lVIpkZ9DqmLM0WYIWZ/HXkO8N7TMPMDZxyfKOkpi48nan82LTz9dvR
n+QDO3PqDAmntzESy4nHrHETY6WuQKoQpDWATBy/Wf/HfegRvZ22EMRF2IuB
ahFn1M1jF3E9438ilZPF6+oauoymqjJ7zHXRiJ8AE4h1rOtDCp1KB7Gfjmsy
DlmaaAO//GGNXHtvWW871aDmTsiQm9uKTAiFOxmgmamI4Eo0S+9OIbyx6DMZ
wCL2kd8wMM07ylF7fQHal4jUDv2DXwrq42QL3Vz0sL/m6OHxhTl8ME5uXeoo
GBR+AEas2ZvqB+M3/3uO2hTqmJCrD8Q0jmtLL8rRCOVDxHehvXmx9Y92UaPE
UmbAij+mWfFTtlxU1xzO1ywVvf7LXibmsG8wNvPtdyix9IuGRAVTbROMH39E
9iHD3fUUDE4Lge1R74SAil6mXdoGeAubmReGJUgjyjw7G1XpDkdzNekaBJPU
9Ods01pgcKhN2u+eOQozHaTQw6Osi1HwfTKgKjH6Y37VSywKd7/SHzEGcW52
IOUWU5jgOxS+L9lTr0yb3dMj34qAXuu94LDrE3vYhnze5T9CZPi6eZNHtkNW
3ycqjudgHaYskPMesl84PIurKj1cmzYpBH2Ky2O2HytqbuwFFq7kyXg777oC
jRrQl4zLbnD4kHLtU8oRfGRlqnt1zcnQKvLL7PMofroS3QdXw9WIXB27rkpE
3xJkIc2TdRnhivbDz9izwcK8q6xp5+r8SZfgysWBTfzE2UiG5xd0SqkBep9j
yjrqilIlcVTCvL4Vn2OEF88x/rd2Oa0f7JAE62W2S81AUhmIpplBAl2LuDrv
CO6cg2gpaw00Cbic//ib/k5gElO4+3v3UZio2Ulpdu96jas4OZ32OZM7RH1U
xxv+fZ+uSgZTdxLgd5KbnrN2uCwm0y3AobkUH0UY7pQjEtMw9uC/md1EYd4w
fcS/S8oRMlrU+lHc9KV/3dBl4STiR+PPGGyFMp15L3UezEmj/vU86bjkvxTZ
u8W1WJHf0OKePsIISU4aCbYkdevsKkWJqrtSFRD4VoCmaBCP3yQ9J8Ih0Mse
IoWWlbbD12MOMhHX7jXkPp5eAotjI7ra7CmofwjgRosxKAOPrXlEAQExYSD3
EtqEAL0u+Xy48pTvgxFNju5u00ooa8hXZ41KvU0fegWVABlj5YOH+wDIA9St
lXUasq50GO8anDnmoPZjJJj2YedSCmbPYrz71C/guaoZj40wP1uiZd0xPfY5
I3gN1/Mr10ztsdp0rTAfozzIQthRMHhFBvgf0Db4vXHb1nSIike0bQmdGJIQ
nUO6roNQLiSateYcDJcVJQuZFhKxD3Jmbw5QoMe6C5EXGa3R3cqhYDQnh6Rq
iVp3xGPon0IGv74C0gfROPX9tkxB6uTYNwTggLOg1oWVzORZVGoDWD8BLBQ4
bkC8ck+xpOGeVudqnACsn3LGhiZZYF9UwztddwRsqgMTUpYhJh/hdUlNRyqY
ccHEoe0g7CWeol+y0/W0yHnQYaNppLGjXP6mOtaO+BMnpFQAp5z+IiOtiVU0
FiozG+Sn3YwYWAl04wmeq9qRNSiUUG0g04iWLLBip5K+gc+by8m5V2s12vLj
mkejX2oa05hCf9UskgOV7PV4tNVGahZNlz6UDLcoF1SdkGSA849xOrIgUIdD
zKXjhoAtJJYOOwO51xrbzsrf4YEPT5OU2z6/m+7nLwsPHOaqIAbaNiTGtp4K
sBk2/IzcCSZdjCljwVKZxx9oBXJTnerkp/lhxjVZRaTXiWUOW7c/fuxnLk2H
v/WDZuUyITiXmbmHlyGaJ7dzvuA6sSYC1f0bu/H4yIPk/gWVJJdQsQiGucRC
mSv7ixkR39YDHIo7gtg/MoqWqXUNLC7/Ka+FEWCTIGwiwsQqCGbaLFHMuZ2h
5zeR4vWR2ZSIePiHDnI0jDdZDMLud382ELuf7lT4/b9Xn+NVx/UHoeUjke3S
iTjJNgzNc751VhzOTVzrzTZ2VCjQClMOOQgd+mk4HXwYuv/rxqnWPxvF5xt/
q4+wefrz/XTM3iZAshYmzfym/AWhtPUIlfGC25xJOCvNq1BURlnoVFKkK2cJ
eCqbgedU8lvm8DpqdJdBVU1+Tqp0sn5QID3OT6hNLyG8P/QJX+5FG4B7gNje
GwtaC/fqlb5h/bZdQazxPZVhAVBFTQKMWVV3Qgj3WdzgU561rcMVwD88Ss/J
n0+7B8v05a9xkakIMqx5JgeC5S4kebeYh6J8d/3Q0Z+EpjtPilJOWpGuYW23
H6yOkg+p8dde0vBeGjYSI1DMW6CErPNr1DHfG/8FziR19lKf0DAN8PzkkWzx
274rcxgukdsUmjFWLpNoyD3ahAZLnjtyDxut8RyqwQ5aZZlSNrZVyFB3YtLe
xpPuPW+AGQmi/mddF5gQ9VCwK2MOcw3lSkk6w6VnsrD9wz8PXtubgXqUt+3A
KdpWhZpXjGXIch2BCaDewG/uMDKhoK1kkzWROTiG56DCdVj0XAC4tJMFWPqI
uCiS7yYBzDfP0OziW3OaT2lFFlejyULLZZj7xlOKz/3fQTZAK0id/Qy30H7w
WpZmjlolNDRBkiGeIslqGSMNMAY6pIDrexJwF4SPMM11LPd9U+LlhB6rKQhh
pGT3xXlYgsWI6+xoLr8m/LTxkqZjoYaWw7VDQQ1Y0F+UnD6avS3JpKcXkunW
wSm1vKb3VBaDrmd7MtWIa6V2tzRqubhLCG984aCxCS0856mUEft32BLjAFoT
rBhqkmggKwJGXzBfbQsm7ftGTvAPzkLp2CMiHxSkC3FZbKO6/Ogflz2eoDYy
JnK3GwUpJDJ8F4/TaMFmhqRCA/1HrmP6qYh2jIOX454arJ4QzNXT+45wcrIe
M5S4CAmav/CSR9Lkucjap6LMs2NrjwmWnGV+vqfXzK9g909qaZhJS5PndO3k
KJZlyx6jD/l6/5Bv36M+VfJzMatotg4gg55slD0i7TbBmMasBCLajNRgquP3
nxzJRTW9zlY6oDZBMoQfF/5Q3wrITUlqLi1w8RFqnRKiJGkLXTOja9vIucXb
FiExlJ1pT8ILGva8L6DC3cjqJg2ubaCB15TVG6kl3/tuMye+PxAHJ5pt4BVg
J+ZXY/UkZnIMiVU0bdrUDXx5FaUXcODaox5XIT1NVisFhNT+05prC/nj9rFv
G1IEtT+3rH/k46eKNc22X3t4W6jd5ktPQnjbaUJMG4k5e0woIDqBQEWwDamo
jJFM/Cq5XxpbqqpNOUQRf2NAuD237KJmgaR1uDC+/rGPvpKmu/HkLWOWXJk0
kqHZP5V9aJw6htmKHHHFG2cbIu7CkFA4XEMot23K+poQj2p+t8JpG63gjZF0
086rz83NmMinss93eJXQpYHn3puw4BGk/mxH88EqrVrj06Dv26rojY7jJ71z
9DbjBAi3uriuL9cyX7bR0bixUbv71nW1RRdK/eognsM3XMOpG0q5I2ukabdB
HjJN7EL31s8wjnsa+HuN/2rVvuFY454lcBi6BLantEmfqRuO2ZCjlNv5F7gF
a9kWR9raWWyCe1hQNcaA2HqqlgPp8wHKkOIHT8a08eLTUfGQk8nC7977iIH8
PifzOxAEwcOY1s/hmfDkpJ4N3KUl6cLfr+hb5PlVTz5LAjYVFanPrjPeyWaN
QlGHit5KYmMNfBTyWhJxvhnQ4A+Ufiz+UrnL1C2/U6xXcMqNLyJeQuVQFftU
yETxolXG2sIpL6x0EjfVdzTHXOolz8kr/raKfCdWn1tZ0t4Dl9jv8Yyau0Vx
4NmdochB1A1MDd1OQ8ao1u3eOPanCpRCSyte/p1LixqngK1wk87I+tBAizZ6
+jY9pa8rczf+ygb54Xk7ealSR/BqdHOELTO5nesJ4JGBcpb+J3RaSAuZx1WC
PacrRXgHBYduttM81RnndS6V2clp4XpASSKhvqJ5X+a2iBtinHTXY4WfSf8q
nwPYmitiDyqS0Q/zUdKIr45zaO9ENGGOBwDNE61DGhaClpEL/NT6dHbe1ccY
z9hK01iJzdLHSRwwHelYP2+BsqOcbKM3CKaSi2eJpMrMAsI4HcgSlmg4HuXa
ali3YUwe90ub0igQjIZ3i0QoFGQhReWV6sQqRcHdit9wR8H2lIFi86HTXgKI
FZbGZdA464GIrCS/8Mdww0vY/uLN8wg92R54sHB8WWMgn28kQMaIqOEWlce5
9UovonUL/huR5d8d98mlkYPVrmCYm9Ee6GzKm91Yeucy/gSqfwlke8E5Ypz5
lTABCKZGAcWLd3XqSQ/Gpa92mfco8hY4zOKD6nEYkyfa2kGb8UYT8jxZxFnq
/iGYS5rep3iIMKKFxVjOHjqiSrsB0tQRGvJrIRsU4aL0cqGZGC7up2Gj8I6x
BY0dgBeieAAVAqUJsfBT9j+WOhze8BfWJAtMtxsnxLrx0RRfqbUVjuSX36n4
fNCQz8xlK3Zr/A41g5lvvhMNaGmh/nSqNJza8MDCElcVP3zJQacipIHRCYjG
gLymlaUZdIeMORjPCNVlrDwH5prqnheSWjHy0Je/LQUgyPZjTR+8CKbI8WAf
zsR/i6SWD/BTz1yZDkGoVc7cgHp3e3Dy27QYjBK1hEg/YVaPUpf9k+IeLqA/
43JEjTSeFkBtqim8MsNotdZi+qeZJx86IUZ83QLpvElrFkcjgeZvnTVacCEd
6gqsVBbdtVufhsJqCPzX0izNknzq+CwDlV0rt6Zusf7NMFdp7KI+vuu6R3hJ
kYGPAdXXRPee9m2H/L50fM6jzQtMuELx4R9RhjcHQ6QWt4izlx4SOaZDPnyd
dZgAZ1swgmudqVzcbEpOuSQucW8a+yloaHejbRnhxgDEkeg+P5xBkPlGTYLj
s0X/N8e09NNMLARnO0uf7uAFQLUDl64v9ecsNkbjn5cENbkL+kUIC3Lk4XZm
eud9SJFiIh3CYCGc4Kbcr4AIZRAy3jjA9qA5TqGoAbbNC7x8CUV3lvBv3yWM
pbx41Xd7etf20aj0lSVxfdMjs4qS8PjadIQPR0PcbYmpbbVMxsvapkntG5xD
h397YagMUKwvlgjh7FbPWHPobJOiz+Hw3IrCf4+EWC8PALrWLXdjLLtts72X
JUQC8SiGoWc91VMSEk3E5CMfceufBnv9kXRTbLMjlcYgE5HX/P89540khqlK
jZFXNFz8P37yMcLtBJ2zoKbmy1Np3ALDifXRHXpy17+JyV1QrRexnp9jXSqc
r9Ugm+Yk9OOkoYa/iqocn8Fn3MgspNLS9bjliEbtLl/1k6A744r8HYwcGkDJ
NwUlGfngtw1IdeMQo/fP/ZyT7CkC7FINymJQoMwxFyEtm7vesQUCi2LDkmm0
EU90QYHBcAmYvX2AqXXFLlhAd2sgcxcBrdGCQG0TfnoAx+/KHpc3wl0fZChC
7qbjO5t05L2lbhFoqnr2KyD/CEKemLycrO/1SUPOoYW+nCf0QfRASIfq5d71
bAX36AzMf26i5koFM/IoGVdIn4Z51JCEttMAKUaRXA5oT94pHY8S2LWVLGVt
K7+HfxflRw7FD0ZRChhmbZVEdtEIgjCpd5gLzAkRjUbdhFD9Ai5G7NA5E4uz
/2PmtCW4vzojaI9kF5Ys4dyWjCoFeikykWJS+VL9sylwf10IPeHcEkO/sP5m
sMZS/DU4sZbKOYbwh2lcnPgByk3LkXOPMMb7udy5YFCdl9vSWwmeEx6Ss3om
So0ZVkSNkrz7ntmBe7qDdGDgIrw9FKELDCF+f2yZklSiTPGk6gaCF5a8AW4I
euaL7o7XWgQyFP8wguyzswxW2cr8bD9pl18ySvS01QW4pu1r2e12uwk3d8eY
scL1rIHKW1iObfAG1hDVrM3Nqwx3K++reO5tIWuXYeiAjt80sWuudiGnMGAa
8cL9B+zFZfNd7vpYXt17vnIDJdScMfy5MexgMdaWYSZYM1avSHj0sx6K1kDb
X5VMP+6iFrrYQnD50F1BcqUIY/qdQdf0v0ky8MwpcqCq9qoOFZcRxNgE/Fgh
Vbb4CGxfeBxbqjKWUJtjgmqUeIDMAnkgQIGJ3Jt08LbG94NUJ9nmaISpEdoi
RIJFwxA18T+UupLzLtN0yJfAYrr8RNg+klJ/u+4e0HbIB9NHYNRXiaveJt55
5OD1het43XBEAqwVF4lBrw4Caz6UEhk73kwridVXLaDEKSk1KOv9IQvIIFd5
N5MnTRIU3Pz56lT/QL1/fcisLe/FpLSnUnHE+k72tkfkShm6/gcTzuPxwlqF
3zT6cKN3mLxHfbseJTQESyH462vg/blPEyumez4Usf0Y5Vj+TdMuu3NlNKVt
Fv+bm6mc2Ugya5RUglS5HuCQpRwxFcxBJK5HO0jjmJyxQ25iWS671RouOH3u
cGPtdYVobP32HZMC91wpQyC1mEConwZZKGAkpOmqp4erVRqbQRtGfMpEggNi
fylNQPuJyofcyZ0VUr7XzmgWdeIX2HriDVr8TH2zupQo/Ojpq/toPyYDrqkQ
Y95ClFBFy3IcV/vqi4DXtLYnzpokFRxO45YRefc2DkzblCm4b0wauQh519Me
0DZSoinJfSBrGNgU7++Be85pbjHpsBSAghIYTuc821hcgPraCC+EtMb/AFHx
KHUR72CzYwuSlk3trErOhllwQpC+bJ0vbnVwh4kf+voOX1tNaYJ9r19iHQmy
LH2ZHZQy2382dUulPhl9HQ7uSbwXRS6TzHDOWEzzo1M7FqOJ013gd0KqNmp4
ZH4OjxeSR3s1WY8uRRKJGszusFMx5PXkV6UTxbY2MsGpyq4d/R3g1Y6jpZaV
Vv36ry8naP56zdmUBkqYQvqdbHfp+K9b9nIOfO4tu/7+r2su8QnYL4V+OY1g
anibuOoOoVuAdSqslA40q7Vnja6OCv/iglS9uaj4110dOGkylUCv6KKI/Z4L
BJJdA7g4X1p3I0sHSf3Ghn1fw03dy+s4wjgMwDbkuYac64DRWPM8TsXmAm0V
GHKGPAZ2+4yfU5clPtfdbcXD8gfQqvE4C4aHTyiySszUKarpke2Dhs88m0SH
dVoCfETNrjpfPBIitkjF+2jwpLGS10/lmgrlOGI/xVMV8lREEFmp7Bu7B7Fi
W1nI4x+WnaXQCzAe66hA8ulxYlnXKHBb8Wrq64nye7NGKeVNC3mKjm3xLCRH
aRted9I4xK+XbGT6eAyzRgsJ7JS6PQGcX5LHILckPGbcGuvlmWjZjeifU+kK
gw9I6z8agkW8rrneGpjV/BT1TWp6MCrSyxDRy9WHl9YtpXRF9iT3sJNCxtXt
KOolxKrf0Yr4VwpTiZuaOWTYUgZ3vvHBluu2creYmharRziQQrEQsV4wjrnq
OUJ9OAtrTuQ9it2OXd2uBkNY7OdgKrK0/Qn5QLAjAfQ7MvfsH/y3LUaJRVgw
e8wLN/f8wx5LvVjWNlEdj/7xUPnccF4ZgsbmEmHrHJyaY3em1+iGZkMIYXHi
t+71sQaXBdBtmNa3AO9dBm/MxBuPaZq80RUOaBx5InNiGdKwDAN6hnEQbHpj
nx1oF0hW17zqSarTe7xlslgjjSKzSjORGsQs3TZH5jBDJ6VHNONBjMEY4BGU
LZl7PqbCSjjbyymkyHfc+3lBggi7CfRgQyk4njRc82gE+T6GxkJvmQD+cjqP
OtNV3mUksLod/+44xtxrpveZ/CFf1mrYTJATxTT94LKZqKGMSFYG4OeWnRw9
nhI6+tPSYBL/GKzdqe2zEMG3mDIwExbVqYhGNuH6sHRo/jGkoEBQ0J6l/QFY
KgDCAQisRoUGHSQKeVN7W7yKE6NrVCLsH3IgeMgdc/B6gr9NfXrC2JojMms8
IUb3nLpU+w9MiGl2CW5hBfaTJgd4tUcMOjDH9EN19KyR1RfzmwVlRHi+jWIw
UXXHoO0cLpcLiDiMx2e/yhgqqpBsjrOh+ui6PQIiKfiQfTZkrEPBEb+sNdag
+p8oU6qoUotxOl22IkQlId+1yygK6V+TDKTHSfvj7ubnjM6mUTjYOIdpd22a
JdyFutJQM+JacotCwKWniS4n1p9tRoSvHhM2t+0VmTfSoyLJAOiipxglBdiG
z+gSLq5/S6/tAj4jKYEc3I5BvtCDA0jwLbHQU0cfF49Oh0UKie1anU9obKd9
E3ZsUxkfabbnaczgcgxLF2J6dHiLiSricXvddWwAHIW4MbZyo385PzlXJ0R0
rn7RgCGx6aMuHz+FlrWrbPhY2dqkx0Ps2WQHkfIH6Pk6fSWojER2wACNECma
I1aWRdvNKI2ratri+1nVKkt+L8TaCGA4cpEV2xdHy8h7PkUnP0yK+se0soAA
LneemZZ87btASxBJV7Qr/Zp8HO00xCdymir2kyPf91DhPzUB2hrt+GTCIfuB
xYFSp6LQwMmHBCpp3hFmQvTC4rMjVqT0KsCqRBgrmBHOuLxlDC9RDc8LB1bd
7KEFgpDU0ofcHaCsg/lKIyGNkjximcnxEVztErlutmzSbd7QEJpmJleq/VTQ
1NB3DHRuJ3MFgF0BR7Wze3GwI5ebI+RzMfiz/8D0zNAY8QR1JwlOQ62I614A
giNkY7UZEn1EL2CoaRAK4QIqG7ZOcTE/jll79eyN3bLCfG2dlLhwTdvhfOfC
YudSSSxCeRFtltOcWVQ5aonTW/3voNTETG09F/48et0v2y5iWOoCJROb9E/Q
97br7Ugn6rvK2JE49trwg6uKODV+790pp6Tyfy8te0vDJ2Zu+idEcNWmWQML
gC47yAz/QSNv4LbyiShu50tuaEmthFCNAyPOfrwZwuU74bAW2cwMACRtR3Fr
pCkzV6erv39PAtDAiaQ9L32h3jUp/1nttatXgVWbwRArIrPUlkoGw9h12FSl
f1vGwm1yPaWnrHCrv1j1dYB+tX1eWjsf0VAnTynwsszyL8z3Whb8riNR7NMd
QnOtp5Q2uNOEuTA9T8FUGZkrMhZ/aReaQ1ErlUICqxEV3rMrcS2SxTWjFlx9
th3CeY4+ZXkIX7zjfTHna039deJKmKbVUMyioljmvg69GvVYrPcIPuceQtMy
sniOfYj+PVgGPQppOqLrcSBlLtogpy/hCJaBDKKTjaPEaS68Wz18g8vZSTn7
0GKC8g4Xpc8IvXhGtSsC2HKU6HVG71Wm9qsJIQ5NG+rH/QfVvWdcBV9pBH+i
PvzDLnqXezoqgr1yTzG/iFSUbT9MEvJ2bRgASDMj9zkkmOBivhTHAhmjh3QI
b97J1wUNpLADqwNXtvplJA8k3wDqOyKCxExrUg9Rcy/RqBBpjAACvN7Cr1fV
drvh8Uv6L25L9mkHHdL77QgRIcSN7CD370vvwAo6d4xm+bprFTPYabl/PJJY
RFlSSQ4DJMaMS3GpvO7A0CkZA8wdWX/bTMgYZuMA1sPzPIAJrldYBpHiJSpI
2C2HRFzi9NKS/emcuEyz2Als5OTBb2YttiY9gXg7XeuPBSrdiFd/cvv2R/Uy
iDHIer0rmV0s3G7Q54AhnIIUFlrCTKBn7XAtPfh4kKXzls0REAFAQhUMKGbS
0vvC/6YFW0xgF7b7Y7+Hr13QhOIB3lv1e1SN3JzaPbAIJ7B/cfi1FM/EkZti
wDBQ1y2MyUcsGzpjjsckd/fwBXrpfIGrP8AeAY6IjVnBWvqv658vJFwSunsl
HfrQw8ozn4WQxl2fqvIePiU4P5/IZ5l4adeeJ7Szdh4jM4KioNwjqkXcC0ym
hsTqe49yMxsZYLvpuzYPtV4lLCKBNEkg34G1wuVCQ9vmCcJ1yMDdqVh5bqrB
g8is2RGgCNxIjtoqgWadkidK7BmevD4mSRF9rZSYvj/FIz8ro2ypEH+YpPEQ
p0HhmonaHNJzT+OHP3Wzsq7BqEZDuQlba4l/1hS2wpeRh+H1lVfGYErRQ/aC
mSHt8PGNLtcEHZL6ljMRpsDddTk3mQVTPD6si6EXpN0CBGz0eoqrFq2iccV8
xDiYm/ZpHSi0RFZMrdhemLrH8nDVwTkH5/Yj2I6f29cYyS2ZtHOIoz7hE5tU
nkjXavISuHIBrEyF7sF0d1JSka5gisiK/ykrTVf7IVIxQ3jcHpoy4PqzRCxw
EsLm3FdorWlkuS/knG0A0ASbBtBPrU5fgu22FmtyYVAZs27rlnly/ikPseBE
Jll+OTs+EFaSO8ioCk6kYYlVwYSYp8j/MdhxVwkPZTrMPzSIpFVn10TxtG4B
ShOdTVA+mPpo/JuxJSxYhCoTT0z8ouVbxGfuhq7WEKq8W4HG5fce0MHXoqUM
DmmQN0ClOe7OZ1kVjBetLYjip9X4U46pOZJX8332pCMG4ZIZpVH2uCAujkyL
yAywXz1BkzQG+TLxTHzg/MaDKKRkIzKV1DfUBhZ2o0jm/HN3olYbCiPXT2Gu
nXMmYXEzUiyf0ips0b0BoOjzmHX0EZmew3VU265FU6uFTWK5mIN5SX0lzekh
kQel6bjxiMJZyry10HW2O0pMGi8jfLD5E+3cTw3C5Q7Q1pDjSfvBQa7uKsHd
Ywneqo+K3dvIIv+JNpRpiW9AJ9APzvtrlBh4lxib6kM1Ex7l+fs2L2NbtwjZ
G8QfYy0dPKYn68vXfiq29VOlJtXoI9g7LStJPNqlYrxGgCflGxWtPSDZknBZ
x5bxMi1ZJKGaHNTZ2QHmaibeJLQ9oKDuRlHBuHx3yBUhy5mca34Kw7/BqX/+
jMEApOMSQHnksh0H+oM5ZT8cENhDuXHLVyTOwHjeS4XmkaXwTJAZSXFlVBat
f9923KV0uh4RA/M1PB/EvfDYrwnHr7o1ti05AQERnGFLmVKrlI4AwvkkSM64
jaRxhzKmylxnWdhUrzHCEHAmMpgc5wdK6ur8RiXoMN3fJ1hKOwE1DLOBGmUF
T+8y2UDiaEyYUq+ejqAKA9cRWICOHJzNE8xHpJYsWBXn4PFtjgBBmVyZzPrb
SPhLE70evR84r+gcZhzT5zB9MWmW6OHsoRjVFhn34aWCPbUbtts0+ehtxPFH
9ZXzwXxRMRER00hHpbsXdX1dS7a4f2rkVFQy/R016o+X+W82MFsteq48+Dyc
fOLx64tFKLFtn53tbn87i+7a4vTHWWRyYM6TbjGKn/lIkZZ4QPkBQgbHEu3G
fI5tynrSrdl85yGjluu3xWH8FrENBMKz6RGlJOitJucBlMgh2GIfXN8lYlzc
4AYVnD2ti6baxIQ4wiYO8EVQ8i88lB0Tvn8eI1NWorHQc4kTsV2CE3Uzxkew
wTrKM5utsJ/0g3KSXLx4Izsg7NSx0YjlR+3O8LVz2odc0ogakQChlx3NZpt3
cwFadi0NM617f5Qj2cDMSnIGKW0SOvy9zSiBONNOEYHIEBslCH94jCU9QRW+
MyuJUKRC0Vp1pe9Pu2TBNzna50E+PP0KRqjJ+WAE/3yyLeZ59/ls32H680lE
zbDulz7UtdmQKVhsv692MSZBwmYj98s/tKyw/WsTRD0mHmF9/mqpq8myW9PF
zIj8lzJnr9VzfyDl18ppndNveGMxwl0TfPBIKDrRZGPFrzhXYRHg0K24Iw+/
KYOTgeA7oK4rRe0NxM+kCsRpokix3DiM80uJl4y8m2ghqLMIzz/EeyJDX5JD
4Uz0Gbzi0tVKOlrTK1Dzuv4XRbD6ic5ggCyctm9GsTbkI0TTvEF5NKb3ExTU
QOrtouwEPvP0DF+1S8EBxWgCd65VMy6zkKt1TVhuEy1fHZnohrN0rrrf47N0
RxIvmzLfzDW6MVFeXMJs93bOEdQXPeC1oUvTKgOnJjojmfG4HdwylIRfIjx4
9s9LztM8kc1sw00c25HFfLb35NIzYnE7jRc4t6I7SoWjYHPxHrG8lV9cHTcJ
eYZY7+qVP0A2v3kgTZVJB+Fh8CdX45PMr4iA2DyW8DViT3UfDFjxWXS7x3Gd
M57PrDdiKY5O27xqbsNBwN+MT2tKCSFdjN1faNoyfica7sQVBi19qddmj6kq
9WJQOL1dbT+0Dl13kG6faOql7AmcT62xIEjmns8IOsaCmv8Uv7634PrlqUlo
Wr6Zn/6oXNF60H4UjgfzdPVWHf5TVRaNcFmLkcsZXOTERMwbfB5OkMOYSCWD
el2EItAjP7HV6uul2Vs8mt8fOgH3T3WFnRZ5i1pkVg+ET3uyauEvZr9gBwza
J/GxfvI31mbwrcc9jZ/WlyY3fjBqdki+LsfghCpkeD5fQpJjWxKahFJcLXIW
mH1V+qCNd0V5DKfe3n3ojo/fY69YDzlXUwwmBvuPbe+OxeDvJbCwwtmpXYOA
v/fYylxSlLPWP4fh/jg81e191oG2KBAraMFiIRCqV0WUuLX3HAYRuZqQRi0q
RBtWfBLsdTq1WDGV3B/c95M028fUOvSkKowlM7jhzncGCLMS8BHXXWQjWLzc
T6twe6WslZLJa9hdpmQ37mtV0q14ogow1NLmL+VWZeL/msBwuJ0uqu5Rprgi
adogcksXKXNsAVIji2Ea38OBPs5uxLTZIBLFy73E39vyCLZYgFHRRUomTLGC
orMcC7r2Am3OxEHN4+tNTTAW3h2tYmvvz9vcLpVlKh4IIC9CjC3DZ9DidZ5x
y1tD2YfWAnXa4on7GqOAhRhA+TeLkQGFBrLmGXofaXqQzjrWO2y19MnyCspP
xMwQiFOwn2XreKtHJAI6mBYJfFYEpSzeO/Sp4+0Fedz3eVs09Ke6/BjZDkQf
gcig9mh7epP8XTeEO/xK5B3S/WF+6w8YqKVbPc2NshLCDlISUdExWXWqpf71
huI86Z35J2fltQPnI2xQsnE6OoVzS0mDgZbL4rT0yow5JpuGuvjbD3J+POVO
v68AkVO7I7mPfLomYe5ynn1EY9wqtba8fAX+JI1W4foYPTmgyw9p86FF6unR
ccD1hIAX0itUlapbIzC+B0BkXp/3vPIkcUznOsOoiPEFvLRVmbxeJynvh95F
v+2SK4zCq63/VPmKygGCr6mu2JgPy3gkvRsGfG2vfv71LijEWYrIaYRQSeZy
jozicrm7xy3mqHelmEB71HVch8Vqv2w6Uer3HOtkHylCgMYq3qKmN6plLZLD
gvfUVZQWSblHFswEAHFQ00UPQpmi7XmLU0kcR05grSWRuIhIx3QN+PuMB1SQ
M676dK7EcoucSdQ1M+av6hGhPNKBcYEZ4DO99wze4FPovG6LNZcFG6TzkYQk
IUPt+VI41X4HpggYlFgN88vdFkxAMoEjAr0MuDBbzLsErH0pAcF4wy3dBNvm
GQEeCeWmXBnaapJOcc99bY8cqkTE/NjLVvjnPZTkX6V+bOOoyiIU1ZEM6EVl
2hjAAN5xqzaMsGSjsNmpT/LI2HyMFcqjaJt5besaobwTCBv9yhaAfrkHxhQy
wZJCbuSiUpZfqKoO0PuxLsWEOd96ofbxWNrOMcR4zQOEc7pWUJkx2OpIjkI7
1bRW4uRcdFHA5tHpg9FYib7o6plzb/ekUVojW8AZhtW1OX9xXcpt9BjFc7Vb
xlsldeNHcwbE8qMvb89ScVDGLhDvwDJujjyHCO4rJqLWWOYj2ezZbc+xjl3f
BLVK0IKkljBssgfkbPXWOiTeBzGB9q2u7Pp2EYam0wKzK9Fs98i6DR3AEZtQ
ZV10g8H2r+73x0tUXRByAvDj/qJ+UG6V0S0TA1H9mDH+EtEW2PSCW37JSixB
RGSjRWtVI0elnw2+SHR6Bnezm6n2Z0v4xtUEnhzfD3d5rZLcPPXcHzHUp2Z8
kfPbEKBObV8jLnN1uEZN7DfQcjUX34IBAQBTLWGSJcLE1UIkGBInxFQFb3vX
BjFiwAZwePh3GxXrHw2mbhDESLGNXmQfq5s+jeyoI37MsgNH6ZO/bsy1AxGo
6PkIZHL6b/z02aMENKbMg74Cy1ew+0S8T+vgVLx3yJivRI0IJK9IvJp/3Crb
S8NS71eQdSkwhwBcqYm9IhfYthjowtJ1WyEQ3KuZzoIrgjsSMufQCejK3NSp
LJi7wNgGAaGY5vPD6YdtDUnPkz9gJf6fMxfBQ1B966MVZadx8Hb3EqjM43+a
oMtMLs/8sq1MW9SHdm27bv4whn8XvIlQZjICKykIvH0Puntbyz9C3XElxZ/U
tU99uVA+cA0z4Ptr05ogxbGEOOZjsuzSF/b5mF9quc/+Vjz1QrH4eRcu2hyT
Bd5YittMYlOB10vfAtyxxhLuHHnrJnEVyFEFWeYiTL90QhXCAELIEzEf7Bav
OJlfbRp9Wj9MU0ng6GoKjOKm24rGg9RLDlB8EV3uE5f/Dfmf21KgIQabnrsK
BO48rHKJFsx56apYzJb+xj60NsI28UouYEv3A0kMDphTMvNSqI/QgGDiJPXy
cX/lu8GC8TJp02Kb65xFKsjoeXm+sWGMHCQWSTTBfFxaoK+gOw8NiIw1r7fL
kyF1RL88eAqbLJXQ4uJAr/yImoFEGwV0awRBPrUdAS+VfCQKYnnrZ5xAg1bz
cwItS0ggi9fTsBrimA/bmInEprEOUIhVGF345wKhD9ToelY6EqWQh4ZPu+kb
99hWytuzGORpf7PA7rZFstt4LHM7gTv8rSbMYZ3zBOIqlcJ7ncIwbJ7Kg1KR
HxkAjowdBdHs4/OFw5t7TuZPCKL4aI5OFN2DoSv48lP2F25e5jO9CFk3nrXR
GOz8gsGRCjhKJCVBEYs65REJsSy5FB8EocokR6ObM5P1/CjfVgjFG9JCoN0s
pFv886kPXmsVfTW0GU1BwFqaPnCmb8HvEkfqMP0bsyLGMS2htp6+jaefHN42
DdHRic87cF5k3JH5qad1zWN+Afu5am56JnyTLoS8TwMqzTco395Tw90RljUA
8JHTT/FwtRnuiY3Un3TXW+M3G+UPcIvXinEjey8BE3P2h8nshDJThhNaSQdY
16n2sigvGcWBDhq6rHf31n1w41Gbfe2jTrCnq0qXZ5MIFap4apmAXEP3ZeMS
vleFnx4SNou4lZtIGE3uJj+YLFCwmrXin1+SX+tILTHh+6LOt5rb0bATOXGO
vFvj5IwRySEv4rkgg1VpRzCgBZY3Z4iIoxATvRvh2sc9cuZmmLCDiLn27aAC
/RwIF13c9Hhc1a8gtXfUpkV0tUnF8y3zMMFIOXOlQHOjJQbZootCzm6uSynr
m4NKynyXohOP14qlWTArUSWerVK3h7hdurJcyc38gZcP/1TGPLXfUjJJ/xlE
oIduZBBYEk5+nED+R0MBgR9Nchbaee7FPv1wifuN03t0TTtDs0o/iYGCLy3E
XC6C0F8pH4r6FdwXhfEoi5S0wo9QO8ZCBhnCdXMJLNHytL+NEUtpIxVXrX3k
Jiyl0qci6tgfpZYQ3UU3/VmpFP0GGs6SRLg376PJW/qvg1CuOZO6Yo57s0U+
Fg2nIHqGSTIxnLl+ZZAeUV20COq9iwHNrz8TXUoKBN1tAy/gGqfTOnvp17Hf
RHgqNG1MQIYHWPLKpBVwsEmzrXGjXkxiaZu5ZxIGYNoixRlQCl/QYOFSIO5N
tpCY2TU1uJSUQzHDALezVxse3AHKIhPbSR3gjjB6xg6Rk8fpRGRtK1iae+Ec
LviGU13LH6dhyywJgWeVvoXGUuJASrS353JPoX+lVvOvLZ5FVZJQW5aYZ7p4
mAClYP0DNvnIiWJ5NezXAqF6axiEiUrywGmfwFQula9UUEsk69SzY/EQycdW
AHOiTtvzwGjzIxwwg4wnyaNdb1n3gVSUXi3KgUbm4hBjms1VUt2HrtRIsEve
v9Eqv6gNNi8tGkaLaprUTCEgEHfmB4g71iobWdLnnGUCCAIbxDLAYpr+FPvv
nQdeiHBxoR9Fkaet53eagzhMwBN6ODP77jOTiubZ7lHNHfnCDcPQbj8aEEyD
QD/YYYDvL43rhWV5oEEnX5oRzUGmLNM4BU6ZxAsY5IScegTm7z9evop9KIBT
8P/MWNkF6xUaFv+JB0j4M8PGtgXveX2dmN07g13SNe/kqDambEb6+E9CEtQ7
wyekIwEP+UeRlhY0719OHrGjd6mw6w464QuiSn1SlEilueyhBIvwKb1NXfyo
CiNdEiiHzcq3NQJlJsQ42vpT4FcqL7R2I5LqMKqqcI+UgFdtvngp3iYSg51W
aFX3HtpBzG8B+Uews+r/foldP9+sq41rsyTiifE+IMdmpH8CfKzqR6ZxqNCn
4R8zPV67VrISADJZoK5ILJBK8KjhHvNxs8iop+/QmOzGAhvL/xzEmS/qwEAp
Cjpy2pSLs0nK7xq4VDTzLQaR51ozOQcHceD1aShS7zR3hg6S6/PY1gVXzO4K
9JdE63a1PuDvmkBSkCPCk+TkPuhZQ9mij7okBPZ0zw2fz+7XikwakVKD4rnr
9jXwcLG4aZAX32K0mDVgb16I4+XMItJknC8hS0kYEKqz5bU2iMty9DGvy6f7
j1FYomEM6xPZiReNOl0QjGtM6pVmlxdufSHkjjOtGhCW2k9y2aJfUJMSotlz
L5O27t/8lAj1pnhjxeMXZRIzmtidNgZeNVaLIBDj+1kX+A6K/UF/xix7T9/h
QUpzWqSB2y2gza/8VoCsRkVfV5dFV87WIL5vF6XOnCHi+kS6UkEMgHJDmovr
HRrrK5v9fMsL6DEYOz9LhoiRovgJ64bVS/wFbcjF6dcnWaqNOwrZG98lRrrd
ZeZdbUVbZGcAmk0gfTmO59OjOQET13r2+76bhXsGx9fqJKiK1IfaQpN8g/Ta
IK1E1PMrJfTrqdJ17TFeLf4uSLugtUg044EwMxoJfxYEV7NXiTuSW7YSazE2
n4X28vdt5eA1OERnsbmHfNKt0o71t8aXA5OUQtJrKs4iknnQHX7vfLrFGfZa
c2DhrkSU/4NLY9r524Doufihtyz2pO1S4PHcy1x4wKGiIx0ow3RvQL7TSzYK
BoikWTUrmzSwZ88I0RAD9OoVTTCQ6hm3nozDihr6v0NVlO1BNJuUiCFHcHs+
VjMp3rnC51mO64wCUA5Ynj80WQLWU9RPU/klrtJy22JI9frwYlzmSk46D3mv
R0vFf70EM16X+fAHRy6Of8RdmaZu7xGi+uPl7eZm/ilx4J7skl67UYyxjB3M
XeGhwiWU/P5bsYeKTVGWRO+RGCuzRNm2TaY1suHCqWWVvUds7mlkuYODiQTE
cf79j+xkqnX/+fFsNNEkRFCZkTnsYo0su/2OfdqQIUB3m/2ndrNoodrz2P9s
oAcvA551c0hu9bbFm1szDBYNQsua8HlstcuSS3oE/D8Wl58arBQHwXPFiyES
Eg2uvlY7WoRjjafUR898/vVABVySYtLb1wz9fRYpvTa3gczAPhgwYtD9bwj1
SEUDmZx8604v/ZA9PF3UMSBTz37yHZElz3no3KeHOQw53b5wbgsuzt6eOsvb
qt3x+f67Q1kyv6P4u2I4KGLCvYGwuie8azZV2derH9o1SF8zPnR2ud+JJBtK
QZUJd8fo5r9IVxy7VKzHuuglGpXU5IFaR8Qpz6Sb9jNZ3YjY2CxXcQL07zNQ
BBCb1S66m0FdQYGgc3PQdaPYOjkOKl6ZuN+ORIIu0LJ21OgR6XgSLvIlr81Q
efPK6Ijalgdbjw5Pr24RbBWTjH8l3W3SD3Yt5t+nFFAzfdbBOzPGNtv5R0eW
hwSgJsH6ORl9PyRzxIWasB/SZ1PYUVJIaoYd+waiMVDVy/mdHQk4Xer0L0Jq
UNhvOp5anMM1IpzRvjHBDYgJ6Lm/zi7SUFX2S7g17O6tk33d+bq18vmPryr2
AHJ3a0/NM60/DiHfIu4XpEj2O2HOuj6jIh9iyYgHULgMr+w03EHoCUn5rRAA
H5RAt/nQfCuiY/3Z5AbblRN1zwy/PCvFQKy0/E7FgDIwRjM4L8xvuHXoc6hS
VzfRLS9h3dLhMearDoZSADqV/mVEUo6y+zRg8y0v498EgsN2qz5gekG+MmU2
xxRR7LObtadA5iCDJWhOYPM90i1x94rivbqx1rkKJfGAes3g514W6LOtohbW
RuUo0KIkJWoiRE3HVstMlaQL4lpTsicogY63OoB89PpgNWDyXpPAlMPTdtMa
BfI9WVj9HV1m9cB1Oo4mSSaj35I5Wc0lUC4BQkowY2ugLQk/EvOACqHt5c5v
0QubaVNw6jFzwYuS3CqtpMH7Plx2jgqIj/LI0prS8sUM+0I2/oTZevDyIfAF
bGCtcYGZOV9+LlSIrpdu/oLUZrS2gqtrNRW4ikLDSQ4y4eYv0fHsvNXnV74R
dFOilmBfsARogC2/zD4JRHfhG12dAZf/MKyw5zEMYLXl1ArD/BMHiHRq5/qt
u36+2NiFmNCe7EO0DZUCQWm5wuZ2bO5Vjoxjw3FJPpFwMWquEj3LzaTMux26
Fm+37Stl8ivBKkdtpK6fVMLrcB/MV5mOFXfaJj73CBbNPKh/2pVxUdCOTHFR
Pzb/p2Sp2wElVOAxZEQwFqW6rsSHwUUltLmWU/ecXEWB2Qc5r9x22fSlTiyP
ElmZfmQIFjrrMppB+ebmg+vrQnoV7MfyX/EYMYQPqsY2Jk4/LlQe7Yc3NfIi
tw9IzYr6liShNq2XF0MvfwKLN0z/vS3VcIpXbzFwuo9y1eCnuif9Ru2hwEY5
AgNCK44vmUKCy8N+QtaTAJLatl8uEzv/iv3sBA3je7uSqGPg9evkfz+TK477
5Eg1KS/bNBQ1C+hnlHKiaK/u8PVxCsQG0D6fKgCTEBAuvzJKCcZhHCf+b8kh
eXbr3bwcSy1axvC2EijPvse7iL6aYPevNDDGsICyAaymjNRiZmHPtqERouT5
bJxCS7hwV89FRL3RD8bZa7la4MdlG8qtvN2AGiduzY525gsc4K8gT3KFGHZj
klA45yeu4JVSjZiMtKki+GepBEFpcmtM7fJklKu5O+hyj6Cs/hhOiIdl14eG
JMc+/4l3Oe4XsAXTYxGeVbmSPeUpnnAJr1r2NXcgUVJS3OBRzC+wPDN7pGxj
dJJp0bk/IdifrTLWTg4SMgEkm+KFyWIKOIQu+CcJZxBsAbHY+wqFYgtPTiuG
9NjJngFn1VVQbHCrj2zLjqMi2EwpfXv/8oRwN8e8+d49aI9kyw3KavMno34N
ofqg9ofx6NB6DFIFhgi0jMk+yXrMCg8uACsPDBU10Uwqa+EtxOc0FjQI/7BZ
4GMNLWgM71PoMRtX6bOSAbWDFjx8PoPvxaM0prb2h9uDGh4mQJYQJauiRRWr
TpYSssnvdSWC4dbTYmptPxmA3W0lGmCudTvscYLQWOzjLxbtKMRISzKfWSbg
oXM5B81AUA1OX1pwznHDp5JIzfnsztPWqoa4OI2NSdW63DcerOsGH9LYY5Mj
114SpBnvuzd+8JcdaJUX2KFzmbKVvklBITOTik6eFupzf7FtxhTLxjLZt5Jr
u2HXrZKRxnKgVokNvW3pa4+Ao7iE84Clt5TVncY4LIuRITIYJazS7lQLo3Ck
BtpzIasIWA0BLhJtfa+GsiMvf9BcgMr7RU1yUq+Th5dDFGHtN1d2TDg83XPb
o1gYV4hvcKlfURUWWv4pfz1mERiwd7eaYY2M+4ypFrRc9oZdWIt43Ac4WaXO
ePSf+fMggRMS/YKOCxbYdYmjL8ItCCCAvWHh1haLptKFaAyieFTUW1bUpq3/
c+k4jGqb7FbddZcDJ+lDULoj8OuBFSvp3HUNX5qDlv/xeAyNGRAgzU60oatU
eILZvF3yg2F2NgVMvpFbDtzbEMUXfrfwHp1EKsMGiEIsjYAVTcQUaqb++A6j
wdmLK0XJFURsLXdjcNHLobZmnY2064bKKaSNCwbcjcOGHsma7pRX0wjhjWVT
vf8+Ekm1xY03gBV1siGcqydQakmW4q4xtxFpMCEucZFKmkjevfMi0IA6BDLY
WnJaq/q9ZnAnNiW1X3FUlMxGx1U4rnKvkp1iZ8BVDN7a46n5/Mh5RRGfHFWl
pSJLuqUgzpz2bBbXk1lEHCdBqC9vl4EkUSRpn2s/FNZPXbDnRtJfaehVsezj
HxnzXgWVevcV2RxjG/a/2OvzG6MMSpvEntL7eXmsJWGp+V1Xq3sP13KVk1hj
5EhV4EbWYALrxbgWXmG1k8A3ATJFwtxLd6QPgOeVp5DNjw/MSVeIeN1R+RdL
zeNIx3WC8OCzEUfOAOZ3aDAhir5q4e6/Ub7VQOjBrnzZxYS2ygJ0vboMTc+1
7CydzmJ/Yggde3TgAYC6hhd+hwKILkEwxVF+ebn8LLVFjfOY8Dbj0uwufO4E
+xWIfTSjDBLT1jS/an8l4SX7b4wIYVhgpm+pzxNzm4KTwzEg/vzxSVutXeBk
tRY0r4111DnT3qvJbI8zpKkCPdNGrgiqV9zqwvis/fYR914Cj5V66r5iFr4T
lVnzC75FciRNquoBhU6hScIox5PQ9Bk0pEkOWKXQ8V7MzvjMRoQrn0/YF6x/
MNIwRtAmBoHPZK3r8pqlm5nziKzz1BfvZsq0R59+SI0+kBauPtcZ14t3YY+H
d2PkO51IqmAXKVYravA5rTnvuSCOA7XEPNLgxze4uh9KadgwxilDxZBBcwGD
tvlKfDuKS5OA9gF4c9YFf5sa30Xyf9YBQi1MmkJY+TC4vlOQAlR3L4Rvpc80
WjYDvA2n12v00zBj3MPlO5QHHlXxsRl/nDSZAL3lgPvzpJxb2lDD7EAY0W6k
6dSBp57Qf5msB9/NAtoQnjsyZC0FkvjvKfpj5Q7ut+eMqSpWCVrGmq5lrY4J
C8UrNvd90ktk1DTJWFimWo6Tywfd9mSo8g6rG4dK04Ph+O+dgb5Oi/VhtZf6
b1Buo4YT/6fhMcQZqxhlX/V51z0Sb9mdgO6Q8qByOlRST1EKZ+RP3ECARuRa
CKBOQSvF3sbDDfsbPnqxY1OqdG+zrI8gBGTYSlCtk1tRKWIWyl5OOEveeNe+
QHbEXj8+GbViOifD27hCk1utGdFGBULUoTLrssxA3IBKpG/Myfw/IuwSxqMB
yQ4S/1i2YlcByHLCI0tMpf20HBbKMmt2C4wHFTTp12rHlqCByt2G9HjY9SDe
cRusT7Ve7Pn8u98F8IgNX4xJVm+9Z9sjTzW9lSWMK9iw+vGosNc7wSGwJc3L
ebvpJZuNVvDKctQbZb5oOhpHotXgKyPQD8OpaMg/b7W5cYiDGm/rLuYmot4g
SHQ8oBbUl4L2rEo9mKkA4JDdjJt1MqweDRnnxePJfQ9o/mgoIOtB+nipPcmW
/Y7HgHTbfyfEQQu7kqc8ODd8Na8E2jMEz1O1RSIe1/ZPbaT00+gsWKEzoJaF
75jFlOfINhSPWEWqR6PPgCanMNJh8ZPQIENfulobourCmpp+nGaHHSTC+cN+
3hSy6IPYGL099S/pn/WiZB5dBnIbjwVmdC9IQKWmUWy9G13kYUjQMAeKdCu6
A7de9j5Rr5tFVELB7yyjL0Vame8CMrWW5UkPf0dQg6fJmTFB8mdb8AkNeCBn
3eG2mFTO4wOnd6Iid/QvxfA6RFzJ6mi2oZjJxKRFnp80zZiwpxhtR86eizFP
CNzzCxLNXawzEKNDD7hJnKahnnJBOh+4AXXNyEWNSjRd+n6zo/l56z5zWmRl
6aTyYN3NABj1SWh18gvOaKH/CdJaEtYpEfzSpJtQZJIKFF+Zt9aXu4DJrOHi
giR0vebgREqtkFUC5ajnNcVTtJ4Wx541fZQH1Rg8diWPxx9Eza0j/e5JotSj
GyLXAl3OMAZTj8zCSrLN+LpThL64OvGr6ppw2ObfjXbaHCDWwcY3Q/lf2qZA
pUwnWo5QEa5PtW2lBWwVGswk3iLeb/TQLzs6Owg5604B2C5AXz8K0v7xQOxt
tWCw9gsK3Q1JD4bz87YIjgyq3+IGmFqofHzpm9hawf2AxkSC2JhJgFBoeXXb
jqKl2Xd2CEj92qM72BnXt5gIwI5S4Ee6SF5aIYIzRhG0sAdGy/WzCECgQYfA
gGlkRg3Oa1MxUGQcbfI/VTfKCr5BG68/VZNOy31pSgQHTgkLtNiO84GdJBpJ
4Sr6WRr0UwqndIMgtUoiR7DlCXJ4Sgd4IhQQPti9q4dtmZz4/D9Wps+fXH+Z
GmTKBPmMOAedXq5i8CagCUsLVbb3S+/sXgIW4bC8I7I1r6OWRToCC/UPgOn2
JQVOQuKZgXa98Equbsc+auMhVAEjOxqTCgZHs3qAE09cdlF+M1lPF7whKW11
e7MAUXouUxejYBexps5S/UziAuqHWQt4z9R7cBO0BknN346t2zYEjU22yeXh
6dGtzVLUtaZDyEl9avZqhP2X0PwNgMNsYgrw1uoOEvtY20+fpTjKpwsSPJj4
Z+9hzqx5Bx5i0lfWawgmyWAT37K6f1xWdkihr057zKdlUzQvbmyyeAazsWkg
iDhMAbxt/wY7xpT/uPOMj2eG/OzMZqL2RfiD+ZUrneiQAm9ket1ZztzGkjmT
mlvVEmXRWBE0MXVFAO9E5+AfbemNkJKB47SVHFhJnOouW3p+npFHUtI/7nwY
9reQpOZnZciHUyebIspKLuVsFYu2DTGcTFplF+9BJqUcrWW7kIAyWv5LzRdd
2h0xHek1P5pz2Tgr68rCzzuaP3G1X8tdU+NL2PLboY+sbh6p0QX2IR2Q+dCt
g/ka5hiDzoSgs8v094xADAb0Rmzbw5AbEDzWbw6jJBO5VIrf+5Pcgk0DyC5S
gK6OLDPUP7FzFmRHi+yHOb35AN1FTY/SWZW9p3icpJY3bXpC3lSrJqRdTUSl
qII3f4fDqKRfvoZqPTZDPQO4Xor55DAaRbHEvXzCbcmQz2JlPQl9pEwKe82e
X3SXh5QkHjOLDtepQbV0CdOaGur+SBU6tD+77AxmP/bIqaimw2YeTcoEnAff
ZNUy42OvMzEpKlY9pHBiwweg2uCD+HHNh4jd5+5bpNqDxXCpQMaPhSx7hGh5
bT8dqdJqFoPRFFgUsu39rluEmImmT2/4ZbwLdt87YpVrFnxzrRAVJWUNTbbw
bw3Lyh2d4IFcvdhYUFyLGy5kNa3JmBi3FyLRPwNBpseiddbzynAm/4KucSAo
ApV1hARu/wdwvi+dvMhBYiyIIGmSGfZYcVDNiHlQUxhtQFayhNYmzz+o3Sx9
2XBBUv5hyakrP2f+IZnfWjtR8a+VfhMM8Fj91Rg5ndkua0ZCUvuks4tCVGUw
PwRojfno0rD9B9f5xp/6s1H8PgQJgrrTZT0sQZMM1lbC1VnW8F1V/dkXNTW9
ZUlTFe4fEGjOJ3tbO0YHdGwYGdBjeCGmJ7UIsU14VQy5PqyGInLTJUhMev0C
+BwVTUMDYtZJDGactPpX2hcV3Uqblvk4QjhmAxNhrCbDqDo/XGSvT/mWPrc+
rc00U5z0hv/u8BxTOKOMteIQp7zfyrPSRjn2FmQdLnRlDcTTd0FRZZ/e9jcj
jzr4HeQg/4lBodF20QTqL+a598He+M1hOMwCpg+8WkMku9qiVLRxqVmAmIfi
01luS1hiH1PBY5D+7T8Yzet24ANWspuWjJ9FyB8RVFODQX+cjEOBDIHN18Mw
CaDCq85kKsX7BdMoZMcutXBU/MKW2vOeq9vu8K94EbzewQl/8kL/eAt9F3SM
/MQXiPbi4i3vhGKwjJQVIqg8KBjcBkrgg1h/WiTdGGhSHtMXMZzlcAu+Jc+S
Dkt5t28uIFEKKIJ3KIghtuXi6qcIjXe+P91iw0FJMe8cuqU4DfOk2SKb7qPy
N2aGXdZ7s+eL09oUwVb0/Y2vFSWLR1Luj0oKSBvpUMAvj0bqXZPrE8f650q9
WSDPZsI70Aw4TPK66Tu++Jg0K8/0l8oXLD06kaxcBcHdidSSI7uD1LhLoeI/
V2DDld0t3RakIjl4r4R8CB7WOE/JYbrS78uuDLbC1BF7D/UMP/QT4UaeWgHw
Oed7F1X/xTa+/DST0/l/AivektYqbsE0qqTjY6heaFb8TSpQ2KTGydXyYXBd
kJhLk/PRN+CcRqDjifUkUQA7N2/wf1NZOHy5tPz8lnVERc4twtT4D7N13JqQ
mbyGEwi9wgUi3UFcfx5D+3ygQlDpYsKjTsyUWVTuWKgnJQqCkQvxbPdBgBLY
0AhfIMXixrRNknuFR6vRYZj60SlRMRsto9QP0/0Kf8MXjrBBuPdpsiXm9bKD
JOvgWAz4SsX9wK3Mr2+jyYa+J1/g22BHZ6Ku+p3XUNLa3xAJXG+Qs5/mQYvm
BScOOhzqEbfIW+1qagimQzXKob8E4RZb7ml2xIjgzciM8dM4Mh66K+7GaKfh
zKvOP1YbPsdA2X7tJjZ2QvHH0KgpbcoQEJu1mVDo5lkCXAaPlt7joYYJdYj+
ZJbgsuNk8Mg1WPTfZtOQ/YxHayN2wpwEwEbd9c3z7utsRnoO1nVHD/ah+Huh
3eEZydtTlClxPi3iVnIjZuzS/SR9WrLgoswSpjR3T/3B0LfKcClQgl0i0PpR
Sg6Dfnd4A5NuF5DOyvd0GYyqYn18oLpSavEuJwXbVa9Ee+CL9yA2Lr7xfAml
IRHgxjrPvT/+TLfr2P38eZTDgwUryGaRd0kj/RZFbcDgo0UbkortJbuHZvKK
pmEUiU0T3UxC7XoI49Hragndw3tNZP3n7WyYdwtBNMKRhCgn2uZKUt+SWBpG
WhrHuG4sWWXeuvia1hVXYsB1oJl5Hp+FN3SGSScGPM/0KAvAY+VL6xNsO0wR
rtGFd5t6TEjOVCpca0mFP5T/nZ3/dfldQj5ASbq988zLuGl2bBBjGqCXxQTe
zCdhwcX/prjT6kUuc/pU7orwnL8S9dxNp+b/j6Gbm4Qz8DEIrHJhuvoHNCNA
wqFJIGzewsSfhy/tWtMx5bMYICtjbVlis7lmFqjX31DFsa1jNqZxs+7cPuzl
4Z5e66HjxCqeyou1z8EVFLP/JGc3pVC5UnJI7CjCu3UV4ML1bl27hOL4FSvD
shzK5AXVGTutDAtFEYxZ2zWcCOFMZDCv5FCZF73Usiy3DK2uqfqT+QHvTRWZ
C3LmXFvfsOgoL9pG/cHbbIZ5UulqeWdiI/3/3sYh8Q+7RPCfKhR5DxBBGpET
9T8gZERe14DdxAqLIrdxrMK+BHIuG0qkKWWv71i72NYO7eowfwFRy2HMZvv5
mj0XuRyM9m2u5Izr+LNwV6M0AYS/9woliOgkLPnnWt9wLSQrn/uxNoqctAVd
gO+EreT6OUivJg1KyQyjSg9OQ6BwY8CUihjAChPM1S0Fjr0cYz0oOOCvMgIq
oKFei1et6c/QOH1vk11UGpqfFkR9JOAwL6sS/GUvJlQ1H/7SxnsfJcz1LBqP
8lRMbuIMXXQEo6zVOvhMwHvqZPjrpuzCyGzwtjSw5oixdqnXU0Jdlwcj66sP
3vZNHnazCxnPLYdsqq+cJlOsIVtjVQ/TDw1Wp4D3qPvMZDuydl/OOqiCCBMH
Ntln9GpjbDAk7Pg4uhFs89EHFqstGfm9gL2WOSdaM7pslqHWICYC0iTfkyRu
kImG3mgeKU2S83j+FeDA5YDQsgDar8HzdCisSl++1BTrvlvAzVU8N6xJ7PKb
QuPwDDiGjsc36eyaB972anTVAzXbs1NPGGFqNwQgzquDNEbVvTTZUdwFFZ9A
w8HQRIdjuJPP/drAyip+OJniq17L0FDFynZVhCzOX/V3aHMVhjPdBKCr3oBx
hCNQ3S+LrVOKF7dRMvXO+M6VoflqqjJCREVa/abcJl01xUkEd5fzifFaMzH5
dN9GjYOfurXLNVrTbsyzVYaVOQM+TybLMCFvQ5y4Laf0A9VhWVg3m5+BU7JP
xZDNk/HZ1hLP5744402gakdeBZSi7Nu5Mbu+8zv6Ro5dOl2SIveNCo0Yv4nG
SoZTSuEltdx0k35JOw8kb1M3u/f568p/mVeWMj6RVUYqNJm6hHhwbjls9RV5
S9PP7xbSLdgGgsZdeQooQ9ETrh8y3bWQpcF9KIYoN0lFHx/UWB+BtB7sImPE
5xuDGknMs0Vmt8uTNK231yw0NU8F+DfFS8/Lz0W6PwTDyIDdoUF82/Z2aRlY
NGWgXTeRAKAk9FXSx4J4KTs/tYVY9vW0ICQpTlwe9LaN3Vy3bH99sB9PnASe
xJWEqWz49Bi4nVDZJokuXw+c5O2OENeAFXydnZil+C2ATSzTnn3B2cHkXmzs
mFufMGGk/PJgG6aJMM6An6k3pLKoIBzJRjT0ejjL11ldM3t/Mvl/k/FV3MO9
Uuwco807+D04nwARjx7OuD7nn91f6iwMn6Owx38BaBEDRIXhDntXkDbsdn/x
VYAtqsBPuTy9CdpyUDrXWYvgP+HUYs2mRBkfml+PId0Xr/3bMEwUT5IyEJsN
ppghSN5RpFXALEaL7GJ+ji5wn2zjWeQg78J1oIveSTEk/z3uj03i/W4ubclU
1O2ENMBRla+HyIj/w2mZ9TQSqybR439vBQKfOWbiq2g3CKWv4ussvMdsBPWJ
W0Ef+dbdbwztYu1WMVOmIKMI6C29OWIWbsyziIc6TbVkT1bUohFlkXhCrtV+
THXQMTzc6gEJDlKvCTX8TmWdlovH3BQaQNTdorVqtSI4uDw7G+vgP9WULBEx
qqZoHDxbyTwNWf+6CMosBV8TKkr9r3OmV5GO+X196asAzrpYQACrdx1bhqLW
3tgZL69AYFs4yZ98gsCvqWNAaf+GPbjJqA9kg1InTWnsb7azHReGMGXQIoBV
/vdVF7k0KONuu/xipL/kF13ohZLTea5gMZ9B+HpqlpKCw505UDujBft4fX4/
seNL9tUgBLtc1Gu8Og4CVLCydYe2k66EdobFyvB6csNSPwjz3BHJ1pZ7we22
KQH2tPWgcE2XpMEXTgV5V6kbjd1fwLsn23HjwdtNFsJ6OTfDKpaf/MHGm458
jS3izbJZPqbhG9XCs8OKef+0BNjcG43ZsuS8bKWmSlEC4NuZkkKgmC/++b5K
jiB84vpD+CeS5Iy1igmgNb0aLEHlr9tki4oC5mtQMQxMuyyt+uEm5EKiqS/h
oDRB58jVx3i8b9PdEWiAorFTWNdXC7acUrTIaTYlwskSVEssl5RZIKfutgmN
nyxLyYQolcFORZ6ZPPaLsjB2vpz32Q/a5bBEpM1k332TTqLuZ+D459N/fvmN
9Q3ba/wFYJH4lso3aqUSuZJgeFmlSuRUaNBEe0fIRT6c9uUFHADovSp0T9qD
3229HXNAprWxZAdrtG5fggUJ3GmZvVlsTn0olO0C74Z2jUnJByxUk5LvzrHB
pgP+D7wdnNyRAOjNomS96Z8p2RosUp0RKgn1bRfRmvIt/OgmiSrWGxecFqHt
ayi5yAOC0jcPMYgwb9HytcfQWAintuE/8rhc7xcPeCz0pWXltrmgjPzhFEO/
r+C5uMK1k0t/uilGBH2aGT5kLhYPZZHFtGb6VQ0AtEaj1XcnkzaboUTNe0nQ
C5ESnq5NugHHRERXVvndTYLNQJT5NgA0JN2OSGDgHZ8jz4zgIt1bJCI1Iok1
+bo8AhRxkWkwhw2pZBIbwjKuUgc3GgM4ic2LEIWVSpIfsqKQCWY8boe3TCwh
LNuZ2Xzc2a/W6gizOiJpWWKgzdXF0YRgZVSFh+UA6Ft7nWaxknGa6Yr2esdo
1Nqrt0cv3qzdI4+gAiq6ATCeAUmKYexghcPL+KkJBkIc7KkH+bL+nCGEw1Ev
QiTGOaXDErOXW9K8lO9MjGnnu5pYQ9LXGyBwkBBQtJpfUhdw5Csw4i+fLwL0
Ce3/i4yUiNwLZepjebMhh5FKw5Th+MgJp05Idr3XsWAvI2fFj0Fc7nURqnlg
BkcCZnJkWUcWOx4I7r7eTLjXHsIEGzCBnm4w1/EMYD50iW8PssTjheds/JSd
zFOyTb4O1QBAUw9nOmRi146Syn1kBX717QbjbCRX0PislgnNBOb0Q3qTkfpm
beUy/WeQOz7ceZWZ319tFlS9DzoOVmJuwYwoRDAK5uuIO3HTCae98WyorpP4
vIzPX3DEBdXMqjseAx/C+dsOGy/Jt5kxQYfBq6UmObE+1/Jt1TUA2kMCq+uR
GGfjgrKny+UNSet8okAgKUMB2bzvYENahF6Z+zNFg1I7ZlwolcM0gQUf5SVX
6DserwyY9dgItu2XvoF/E58tqII8/z5EbyhewTS1K21vfpJBzSZQbkGYfsJL
2bv3CYqipe6rJ5fiRdgTyyMdYNFIoBONlbz1EWm7iGWQfsDQ9ofJksQyWhJH
BEp4PnyAJof2mlusQGEh0EHWpuS14Kc/hVIYa9uY8+/8evvdFKXKH6+kHYg6
IjEZmRc06RpyvrZSFTqsF9QK8f8G6bxbssWawV4DQFGfi5XnDbUf5MvUC4eC
7J4UzPIE9AjTRRp3b+IFtB6iNF/c52U6+RmmHeTk3DrK/+ltUmciHShrZQ0h
NIctKG6W6lA0PivCR+zR1/ryj+6Nm+nTHHD/dN8hq/mUbAIm3hJDgpsrHJJ7
f4IfkEm5dyhNhJduSKqAEcLRX7iRaqqi24J8r++FojyNLrjQCxUrSEK86i9t
RLh+lM89soe1c6Y99crO2H1dtByI6tyglNm7iSDV1WN+W/0nJANgccFsxFZC
/oKOTqtM4W+rD4qPllRYiKbMxRfvZizLezIYdP50bfoU9Z0e4eqdjH3KLUR2
VXO1vIqJuRfJoaCqUA7AZuklDX/GgxTg/y713ZM8IeXMO1Mo91+K083dH1mm
dpNCFWiZ2QrJ3pPaE6tew93152mOJkCHUCuwtNcgMmt5z95lNREpK1Uj2h5X
EL31grVjeGE09R2E1yLL4zMZ/y0d8LQHoFZ9B4sthAOZXwjOch6ZoiJWHWod
p9jzZCMEsADn2ZrYNerHIpAwhVVlK/fwdKDgYClI8iORNk+tdiahFGTAN5P6
bDKRO50dnkjOCoEQ5DqLhEHTxmfMbafXSzUcRRNAjncktB0Csktkgb/wJPE/
gmSGjevbQotiMYCSnybAl0lKzK3QtOmsUX05yic/AYZvBETLMLvTGXPnj0/w
x+VYx9ONhtb7fheCPYPvtxHy8vrncla/ijkTn4yyBcFAxghvWaWoZUK0m9/B
Z3G1OEnX4roROaNpJV4sT1sDNqIp4NFvqFG4UoSgEotVi669/DkWkZ4dKfNK
KN3FNRNI79G3swfBQrAgLqV4zENbb6fhxnjrRRLtQEwT0LRalaHmetrr3KL2
Q352068uzzFpyRvcSRyjMtZ46dqOgvZSCVfWtVtvsKiUkUaSjkUVAhgEnFIW
RZT+qzCreS/LlmMHGMQYDIZAy4iSquzkS7wAPL2hIT3M8XfHnYv6jRvtnDiD
TvKtJtXtv1J2LB7ToPFUaFcaqLQl/K+rZVMtCWj5L0/FZpvmidJIhNC1yKoF
5zRqoOkiBLhP8GMj7AqSRgsDTUfOYGphHPIchz4ehnEvhTEUIrj0EmEgDVvR
gmmO523b2oQ7hmdcTq8MaqTbK1i11cjeRVjax4CqvbMz5Us52ixnXg0qDz8E
ABQQe8czcBwvmrk4JktFejsAI+wqr2VCqviZFT3I9TLIcg8s2pHTzq4a9JLd
imV4QbB7Pl3EtcCCMNUvp2FK1KLdxtIaOXU//tPffxrH9J4bo0yJ+DsQKN6i
31DPl9TryY3Eo0kX/TSTAugVBwOh6lcLMB6f33+KBVE7ar6gR0X9n0P0KLg7
m5axozKppRU/VbGfoXje7F98don91Ob1csiB4vR2j1MoRLoZLhBRAmsIKdbp
gnIs2cx8V/VzE2tNcDTqHUddHIMm51RuH7Tbn2+332vbK1bozMxdR3QR578Q
DYl3ozeSu0umZ8HNI+8vDn7g3Do+lS3LSdOcDSg0p6ELtWy9T1NbwMxYkRL9
gA4tCjmLc/LF1Utv3vUSBQFFnnMaFzmBRKvgVqRhD5Jry2ZxoL5eCoEb66VT
mq5h4guVacVUxnUySeGKhSx+GNG+HPSLHvk+lU42bHks70uyg+2i26mVi3Se
Tojk1sW+h51p3UcEXeN6bnM0a9YenxnCQ9t6OYE+jE+EGjTpQKiSU7QzxHc4
Sk4+Fp2oJLpKJ0roVY5jg9EoRsMptiPqiSBD2NfeiTmUsGIaWS3PJQtytxs2
2m4qgmxA5d1ypRGmlRWjnV2mK8dRUXqY5aH1MIvCGq5kWMpESIxmr54ZSfX4
at8mJE6LI9oYClEwejwRFNe1xhA2LHhVLc3Z0cUtDYMZm0p4g35U/Pc+rTwU
04YwPErMJ0CUfdIQMpkSH5qGhRQAmwcKA2qxHB/DqazT0FH3PYP7ly3oaUJe
eZfqgQVCw3QOZ8MhuA7HnbZcfRh+ESAmGT9nJHid+yPYqofS7yjj9iCo4knZ
CatXwZra4EB6BOSBkGOLtodxH44T+jzOWVgpOL6bu1r9OjLIJAf6KPf6kb22
nSCTv8t97/apugU23P5LlDVIfTkUdib8nY1SmL4eneLa6GvP4uz8MsXi42US
Yy73GB3ksQo7mZLwn7Vy84inv5MtDlunOI2VSrEsPtqEkO/M8toqF7Ge43VX
21KPo7Nm+eol7n2usPPWUr0CWT3ktlyXfUn7VPuj38wo/caa4dh2pjBlqTsX
uFvW+Ux3TJJr7ndnZefO12pzJVQL4GxpAcxRmHVKRQIiF722ix1EvVgWuSG9
yYQSSbh8GCTuDzR9RwpC99UhbTZs49QON72H4GCdARnc7ZG5rtDIJDSGPyRL
2KUf6/kalNXqWZehmVwHyK4w6WigrsOXxrwna3MERnC3QeOhw6+6T7s2J+Kk
mnGQvm9LvVOhmR9OnUuMj3mI9/yn3iF5GbvbBLOZUtivOl76ibDlX+8IpGwH
uB7dg5xYirXAECGchVQ47/nbOUyfa4T6e44gFQTnIfQb6iRn8i7CHPRV0rWB
8jcjobbUpLxq9vXkiUJUcURGR17Ls28+/HjWJbivGU/48mieGiogrsJTy8g8
lAokimVnGAM7IAdrwiagzRrFkqrvG7rC07A32OwODKwQmUnZtiBEomMOnAqm
IfO7ZR7vE5Yt88bEVKut2rDKOHVBcfFmRqt2i7TpKH007Hu1AHGb12lScJDq
0tbZ8J1wZcEm7DIQcaeS1bE1JjhKKDt0knW+rdIiSzo7O40kx5E8wfstGZsp
/yu5jWhGM181oSj7yfY+tHNTe9XRodH6L4gvA7JbOGhVSfqxIxxyI/yab6Ae
AAq33dFj6PlxjES+LqNda2nYMwzGldsiM4IKlSvDsijrUJEEKGp3VF9jU9em
ge+P/GXBZ7l5pC3v+t0Ww3M4tF7MH42Tgu7g0TI7gARiqV/D5us7YLNQ+Dkn
OZ9oRZOA1AYHheissMzq7u5YVTEpHX/hPdc0GlRQtL8JkDcjSyWU0BYt3q0I
3QPCZCv5XB5orvVQjwMK0NKBVS8dnKW6v8sq1oVl9CYIMa8xfTNMbkmujWOz
2SQ68Rdg9SfSnk6wz6Gon1pF3Z+fJ7RLuUdAHFiAmYsvsgjX9Z/9p4/HJLkI
/7AF3wi9kHz+tqKG9CeuxVnrs78lRMaCHq3RrrH4ieX9oJncfkq2pcWK39ib
tBoYrui/8ozGMubp2XPlotf8HG7xwA3Yfk2ygjqmGaqHvwySvxCPPwwlrifk
KqBW3Geetp8tBxQK2m6Rbqz2CsiiESTIsapb/PFM4cYlprwY3AwQzMf+BSnm
yTkB9Y4k5k7nvsw8/Bwh6kZcG/Shmk/t2mUdONf/TSnHrLJZvRC1ebQi7mg+
GIQVWt+MYZVHIl6aultOZGO4EY1gHlHX4ma2GlBAYSz/jeXrixs9R0ltvFKJ
HXb3Fk67lvfy7VRJUZKaMfcEm3aWAUn+7xmlDsXg/bw132pDLm+a9Of3xn4f
vYhIqPAsPsoEL7IEERlR/+4U6bIabXFuREqUyovabPLoj/zUavRN3mIer6Pj
zK6fLqP9DwKBMjmJyVNkJ08NtetNkFoOhOfIALER8+ca4uvAS0WlIGTqe0om
cJMj9blHknbllFXf5f2k/mg4rkM2vYmA7GcaE0+W9nIFRa9J3/WopdCkQBBA
jwI25ulbXomKrzOAnRS2UCBnCCGILK2C8ESXX3hZg9u1/o4hj9Szr55f77N+
5MMjqJrvNPoKvJOXplKp/RfoFt6TfvrXWmfOq40huVdM/JpyT2Mt0lFStI3B
ThkjKAjUHPTzl5BA0iT4JjUDiw1P83uNBuYncKzKkd93lkcohs6m4I2sHNVM
Hxg+/hj5jiH8aQ7SnVdtsk7MIUnkMObPPSFYFVztY3iFyQ4NNjDAoBulTsqg
seVMc5XXkzRmFQ2U+LiPb6V2Ap5N5nQFs7gxiwOhig6fw+Rq6GRm5UVQmivy
7wrqI0MJ9yHbks1jdhF96mQghUEOJEDqJEdcxyV6fNdfNsMNQTtXuqS0HCdp
PdH24FJVy7n14FcmUrv2fmrTdD91QcZva7/7nJA+s7fYeJ9zgaQwpvx+buMB
ZTm2++ctoz/irrWhhJvgMNHiAmHpQEZhaKT1bMMw5IibrM1rMXdUSBj2s2/+
kZI28hHnToGehcFH89G/bh4FUCZAbhnGFh1k4QxdJE4sKINrfgoYuBfJLOHj
gU7BvBQ2ERcE7rDbX48/rPjylLbMenD9E3ynxpWqvggMJ81V8dmQNgGHtwf7
Xm+8Okqd9pD/5Bo5bIKsFhDmlTj/je2DzDV0yszqQHkgpHxKOhSY/qPvCxF5
9/VJhZPoW3JVaR6l6zVR0P2PiGj9f+bUASs9mPVLN9JTgwym1r2Ixhgx751W
y9svhvjXtZeAHtlgEo2ck8Rv4w24MQ+Z4d5t48gN7LIV9Yxy1lkDGWnMMp6f
jJT7BiHqI8wJDM0g7oJGF7prOauyGvNgVXkj+vrDpi7/w+bXnQeCk0XDYA+y
mbACE3aBLHpP73ttCPxgaQZXxGPuGQPzrIrWhC21fJT8FbiMaFsjqitkBWMc
LVlzVTD55Ar1w+FVrafGKt4uzK4BGHYkWJN7vqhtsBgBTBleoEob3jU7E7mq
U7xV2X/Qtto6fuvGaEXsUoKSjhZ6mfoznI0vI021Wsq1g9Fb9AZe0O4QNksZ
lTQV8uK1vY+tBW2AQSS8ff3CVn2uz9Zw9WUn+EISJzW8I183sZzZky4+rYro
OH9bYYB7X/HLoRvaR0z1GzsSB+BD93OIqlYu+1o/dy1skYdBgXIAxIcHNm8M
Yy/vX7C8k0SR04bJTEV7g3sMvVj0y/kCY308k6NxtRjzBGYPSUZWjyKM5aMV
rg20zwXAuecwt8mXRVl54nGwEh+dypsv4UKHXqLrzBF0Yzh0ScFi/ZzP3/Df
STugvs417WV2N8L7avbayFTsng8L6/SB4QLjWHokq3wyYUNEI6gO0UC+ShqK
w200wPfOPrPyiotyFvWl6pmbpce9Rh3sGArUuTDGTMdq/uFtazhPSJAH65RJ
abI5/+DZTELcqydRunwT5s6Djhie6YghuqMvtKhkDvuQS9XQ/NeUgAOsiu5s
6wSJ+e7DCbZP0J8pSuwpgDhS2vdOKedAI3RMTiSZwgKFZ51QOmOmK7MbG1qk
/v3VyWa3miJPLVidgIC9rvPe0DC1RE2RdQUWFSKuDcv4dQ0OOOmT8QJEATrG
7uJcmF8aXVFIF8S2T1WOHYXUVA4CgEJec7cjbDyhcDCdQcdXlIt1PFAxTKO1
i5OfiuZXICjNq69WPgyBpIsJu25KJmIx2bIOuSEXqCUvopKkxd4MAdwrPGBp
E1TbZVjHV9sveD36+t0zr1sOtD8yfMSdnFNZnotJQxufR3bor6TukeqRWw2l
WjDlvhRWj1ShDsAiTKeyfaLZz0xfXnLuTbgRAJMChOy/PhLiLRwa+iCCorBC
PR+OFZcpf20kO0/FHIwD58/O7p11Ow6vYkCnX0K7IKC7KmwTtWVi6YK4xZgX
nVCU7nVZQy+hAlyoHuIBHxbGbUak2thX9/Ab8zXa7Gmk40dRIsSeQPxP79LF
ve/EtlN2atA+DcB9W6REtJz/SawxxrjPMpu+RDsfXefKTWcpXC0UQQ7H9Alf
kQBWDLDzHoSMxU8uswIxNspxS0ja/18QaE2dRUzdIi7M4ViJaxHLb2ydMFVF
MwEkR0JoGV9v/ksm3Vl1eQix+koSXIHMzHuEO6wxMMVuR2ETkJ21J4rXlFpN
uWiPJAo9S8RMb0ecr73/v5ob02YTgFE+SszOBPrylBDASi9F+/1lYl1aIl4A
NaCmvQ8i8wxJOqaFeirxxgqE+coJgaOHFPZ1L9DqTwAfjfZfhVnF1HWfBjPa
dd+C0F8ZlA2O5l3CmI8ND6zi+RyCGvIQVXSxlfZppQCH+sdvedcUyfXnsfAf
vpB34+aJw5kZBq7tCT8eK267wRYs3i4XTuKeBiJT0Oo0lra1p4RdHZvBNoTk
xzjNcfijp2tVUKuc9YulSKBgluDbwgbbZR2WoliVdpnPImvna6AftfFeHMqD
7wU7qS90K2z/Amg791WK13Zdt3dmca+xQJG6qkVGQIu+C7vYfQxXUcds1Wpj
XTupoGbNQgaOgnsUGmAngF/YZCM7pK6lEQrTwUBQHSPZiL9zKVyTDaKewt4l
X0ck2ODLSlv54jBzP65KNuDnjJb14X/dhtX1HAiEwFjki3JMMFsBvgAKTw9D
wpFA9lYyd7kEDue5nl2kqyhoIg5JZGAbbrB96T/3WgB/CdT/xr+XMtTcmw3I
9RgXInGeUJ8uzfPTDF/v9mkc6UZQUmdkrr8Th1Qmojl3amAS5YgU0ODwfGqx
P5sHTrlE4BJTcf7RWauAbswBmrbaxekI6DlLvgHbRMorbuofDYK9Gcb9/ZTv
WuKnoxQVyHkjppOkLzRAvddIJuMB9YOsmAGaubVaddetbm+I8MokGK0VeDEZ
sP5aEWt32UN+D+o7+MmGjxTdBwlyzcvTunSX4iQiChWdMBxrujX19p/Zvw01
CCJWi5WOF0iO/Ge7wnDER5vKQzgcl4+AAaxZkaQWrCWzhdaAhQmyjYXSuSKa
L2Gd1wtqyd/AqiO6R+RoemyKnGBm2p5I/kMo5fK/L3XBzwOeJZudu3HJWJpP
WX1yTmi61dCOfDn+xSVy1c35UKftUIKFXtmo3xJjhKz+1stTAX8eS2dR5fyU
V+DBiey+NmUaa/nUlZC6jnJQDI3+dS1bCyysbPe0S8r3Q2ac0VBqVOgAtPqc
dRdqBjL6TqVokCTYPhk1IoJ5jMo3Mtnh6AfCQL20nEO2yCYMlAqhI1sB+5Yn
gRT5xh8gPjmHjDIwMWjY9qQmAiwKsiWMeu3NTOuNu7S343ggwKCnGnPhIwfT
pXMgBy6Do3knHwZFJgr13fkk/6M0XpOKY0ytlLsFH26mzRnbnN/1KjSwN2X9
S4sHC4hh5fqlShu89/TbcmEd6dnmp4eh/G9GAbmdJntD4hExUiuzGlV/SmcF
AZreJC+mgZE3c36rkB8+16OMl/AN8SHUvj2mxEvSB37NtMWh/aTnPT0Nz/KY
XVFn62EDRVlt3CBwU16z40ks+D1ubbCKwKU1VOCkPjzRVGa1OIfR1qAqIcx5
dMCytsq0OncuTYCNGMYPdIhJ4NM9I46tDZC0gXg0zIJTPYSQKr27H7n9Pw/u
t3BgEIhmK5ZNVr3sc8KID3q3fLtX6VlqrGXR9myYqhspHasA7n2R7aYaAqDi
6YHdLUAJUC63umX6H8uJncCMKlF90UctfNSB5fjUHwUGHjrwAkptENxDD5xc
gclhlUli801xW1KxIGWnANBtnDxab6agdt4GkwaBLrnvSmUTbEp8VaIw0YeN
dVPj4D2PLxz1uZ5v5arCR5r+6QwGMp8uBDYSlWZeDp5I/uQma1tVu9l5kmO7
J7zF2WmR6q/j+tqiqE9FJOe1f3HZ7dMWnkxWsM6E4tbA5bW3NyI5K3Qiv3m6
Awvt2BY3tbgYBSk2rRfAa9OEq1WSXa3Amn2ukVabCBDbXh2Zy0jitI67x0Ml
RdUKcEJyfPB1YO1C0EFmwZfcIJohPbNMfwMTbzac6nPZR/muCXfdXwp4ExR+
nvdKfDLe53JcO16rYD+o78vX0qVcpz7xVw4hgGl+hKkiTthTS8SAyW+euGfU
pGwuevLoraw2QmFermbsmbxJ1mhCldJS6sRN+9vSiq3NragBgqJ9A/rHWwnb
X+cPxj846YK1sL7pyIbCh46a2K5VvbL4wniE1nA6EMekJ/8+/Y09pn/WAfUL
e6TG3QEWD+6NLIo5w2nHeNJQLJDLDNLQR8GI82SdwFD1qEwWYoOTFuDwqIz2
sjvrCofAgjimjTFfzjVXfgg/z3CpaCh7i5Eo24s2HZGP7J94jovAmYoNEopn
vtmrRghhakPzVOejKNSysBoHYj270Ih091JXgv/uyxyTP3gQniZKrAptF8Nk
ZWBn7oLkWwIG/VYeMKXzRb3bodKAAXA3VCzdzMbv1YMEOIJIe4Dkq58jktEb
gaOC7iw1vbIKlzIM+Vas2JGOIcagiH9yR5TBLzTgJh+310fgriV4BAblmpzD
u+EUIZKJNKRykXzekiLj3QdL3n1PzYq/BtyvDTWebeCTZ5SfoY9WJdZ5i54T
t7lf+kbrVyBKusDRTcBYE96l3zSe/rUx4LIS4OfF83n839KpxUi2DK0gN+mo
7h/ZVS/vpCzRjJSrHB4YEZW7DZn5o09txLUipK8+MAWq961n8XubRJb2UDsK
RYSk/f7WCfpaQJ83QFyo1lZtuYMdiS0qNbfrBeg9K+Vz2bHhbXlEfFF8UMzh
+Wdcb3Vn9kuf/4zadRfGqn7y1Kp4o8ni2M2rZq8QVX16hDewaHpQGDJEFET9
yixculwuj1gjqgGyZH+eeZ4xTqUB96Ts/RyJVBIXuD4XCSyDlx/+1gbFv3JU
HOM2uXY8XjD2VI3KlNZa902LToT94SWJnvNgWhLwT3fQ15twPZLWEhc/d3JR
NSJ9nUNZmzDJSPfaFu9C8tC0inzFBFS8vp/st7KAK3p9sskFFX6pRiasbJKG
kdwH3liR9PNFBqhvEqIc144KZwSQIzElI96MAjq8IshkJCMOf02OxmZfBY5E
m4jipMjhznkEt8tJz6PGmj4+B5kgGBR6m2dW2Kv/TI2KwxtezYAkChYX2YSz
GrCkR7lWEpkg3Kkne4NHA6MwME0bqAGRXauhKb6f9QoT4OsdhasGTwR7KVJd
XC1uLHc+BHbdlKRdmwT3V12QMOWmMp5jkwguPO/Jx4GDZCU4Z+E5Kvw4cNgk
1erHD3hHyLlZvlniS3dNy2jr2f9zOVM31vC/c0DcYgyPPLmKls7+8oKNylgg
fIQHiDkvXPUALmxaJFbSj1z+XvhBx3m3Edg3eWow/w1n3NgTkaaY84ShkC9r
kQFQlcj/9VE+ELsrEu1sHY2mycy1pWZVXu4HVMh0jkLruoPPZeDsTp5LkNoC
do5x3USbuuupYkY2VmlcWHdeY7qGY/CsKTQif/TwQ7x6NDkGlBNPgWVVSsn/
OEth2BweJPxdS3onoQpnFCeGJuRWCGkvWC2sExRu/gHgzxBPK5aZOm7nQhJV
wywE+CFt1URl9TuBMzDtPxhpVw2kP7KgzhZ3gt7D1nQTwfBGvSS6OlIrw1MM
p6A5g4Om5afvg/sXyaz9sl8Ej5XMbFrVogeOUfZXYaXizqXrxXwyY/fOx2n4
EUjSnZvOPT1WP+VjWcBtioosIzUs4LN8XON6CG/hlB2nDqQr522Ia+CZdjlT
W858wksEpvhhVDd78OYPvva4/1pgP/MtqY0H8tfBFUgsB/IFV+VDVQ8Xp1Kj
fl099VpZyq6PRRb9kF3zVlTMYrzjvavmzNiGzSluaKAzzu3P9jKE9cLrftiX
EJ+pIC6MDQNMUYi9h5PARlXkcXVTUMbo/9rPXFnYXAK7luJBKSHDLyj+mxms
7gj6Dh2zTCjeS1jfDJUkL3WouzzgDqv6omDQrihYfO0HBPKxtsv3wb97VTN8
WH/zPCh7bDo1fUVkhQrSgVdpKMmXB+1NPtF+5GHl43L4/p7DM6XzUNvBGnlW
8tFQuIF0Ic+ZpP+/6VV63dMICxsu+t+bVwPLdT3juLXGFkglvLi/g49cOsOX
qQ12rfAN66Z8yAybvmPPqoW7BnaRYyKGK/6WXg8NLg/Q5c9ZoCMl2smcL2av
e+4LhmA0pV57D1TxzXf8SbTBPcqPExnKDOA1GUKIy33yjNT0AmqghDUEgFIO
it0xbdHeLCaHqZWHaWIGPEDrmnUKIVe0X5leKjG3AUF/LhhapGN1EVVj3ym4
AGZDRuY1jziVHyHP9l4XUHAhz6UqMbKD6k3d93aVJlg2OzjfFzEx9UXFHwSx
gjQ8e0A6mqrsZdFY4dfUU2Jm/OBNCaIKlrquCmzcMkQ7cgWglxoCZREU/rEH
rQS7jLhCP4+nIMbP0MV8rfgVHaRs63ln6j4Wl2NU1RyBPqdteEp24gKpMi2l
0J/XIP1VpjzNSxY9gEvh6W8zbwXLGbDu8PdzMqMQ31ppxpWcceMJManswcbR
Bk/qIdbFk4FY+gCLsJgi9ynT8Mcjsi1zzSNiMcoTqJHRCaw2fqiTENVe+vNt
idmRMVB9iXQotEpx9Rhcv/Zbjg1OwH0TKuKJoaTKqGIS/xT3aqe0rp1+b+Ke
gnnGyROZrIBDwixlhFS9kfzXYYFim+dLpmf+2Lcth1IpqHBkYgUvqYJp5E2m
88VvZacN7/dK1n3JGBEJ9YH0L6M+VtLZjrVifpEuxhOCUAc+BY0ytVPzMwdW
F1JbnUr2SKoUONn4L/uv8IgkK+MfnOL88kotN8iZcI2J4SV2PUw547o6jNXl
iC0aXRHrEPhJifKMfbmWiOHn9LDjia5EE7KFoDS90ED3g/jmD0ViNf3bV4bb
B8sTh6NS7RnAoPSGsl+1jyBPAfImULB7l6fJPwpWQH0OcuywOAJI9OPWtw+6
n6ZBYw13B1yNzpzi752QZ3Is3um9tiTuM67lSKMD+DujzS7eAKwot0W47zos
L5H3eIUY0ZH3oz3hgFelJuiJAF9/brbcN/dZSRCTowvYF5UhTPpUtJ3VO/Rj
c20Knf0MpJ9k5xKbsAqKy+YRSiv/ylNe1gjDw/j+9AS1TY8RgxL2oECOu2oj
588CGmxmFSB2OLsJpEGcTEQRMiMIwZ5aq/ydKwXlxM97cW5apIKfzlWfXWPa
FUFjdShGtBDghlIAA/OmWUUTnkA4b0M1bwpgBVSy92HMn53itu/58Q/sg/75
I3ztOIFGk2AL7NaFMWKEltfqGuwYKXxW+HKTkWaevzhKlrDkRKxnwK9BLhaL
ZepA4J24Upnzyt+2+cJEOF+7wpcVfMzpIjCJTks4ysGJVRWfhBShz4cRaKhj
2OXOFRKIsb2fjBl/BZIR1ev30qswA+Xb0q0/4J0MTli8NA5880mk87UuwEm0
8PFZtwxA4mqNshr9rLIy8pEG8PzweIQtQef0d1qa8QvOYTkVTLXySRywTHI2
zrr7liKGLbxenub38dgJj14Us6p03RgLP5Wk4UiRo/u61m6j+t6xudOaxVLv
BE1vsct+w6aY/q7n0e1xpTerPLixQhfRA23Gou5AQ5IpSkHUL6ld8fIzecOg
DrY2Hz4Tn+bh/imZY7b1IF+76XZ43USAQjh5SMLvGyBe4Q7oEjUlEuhUM+5Y
QyXd7Gch8rcxbDeaxxPIv/vbw2EO3FPvQN6INxH9t04BJIuJIDgUM3vJcstt
8spfoZyxkXAX28qmlZfoYBW2QERr22gLs7EPYLWcOIlWXw+KAIIx954s9OcQ
3aFjH8XdDSHRmXYcZnOSfwcDOtmX8ZBu+O06RT2gPsQZnCRWuHwP2CfoylsF
FOG6kZeAtdHGjwaIhmkvRxZ6KsaxP6NzXYCHGI+sXeTNIO9hM3tSazuB4yX+
MWuTwO4DKOGJ4z1MqcQO7nabiLQE4ODV+7myNOgWy5ObQrkPCqy6fLjZm1YR
dll/QQkAta8+cQM3Tgy2+lQL2xjySJGKl1/nbA3HvHf5ol8peauwOazqduCP
EFr2jkVnDqJF0D+gOdoudg0nFXUqopum31dzRSgSzgHgS2JEVA3SLkPl0oxa
ZvXeF+vl/5D0E2GV/vQ8kL+DDwdbIcu3J++EO2BmJrouAGWSuo5GMRWO3MCc
etA4FSNDljh7872tuw54LrZutdr2I6YEHmGzsJRarQxI7PN4kCL1gMvxd5MQ
IckFyA3gNJx9Zi0tb/BDph6I0H61AV8J940GIb7HlbmzVSjDAokY5cYe02rt
hcunfWdW3FurZTcWKwsVWGUDcqYYGTT3dOCFVeJmyBWxNupBuoEeOX1Vevwp
KXJgi0QAT8mcFqYM9u+qi08+Iii1UCb46WmuZWV9L5vqaUo43VFd3echAQhn
hd1ynKB0UM1s+U7NZwr+Jd2mcjDyYznl3VbxuBirM7km146HJe9X2GheCKZu
C90FzLG+O6bT+O+kctcfmBvirOzuxdVkDbrPaPtTjWVlRG1N35Fc0hy0aIMj
8NxHfumYf2pAyxE+wzZs5tP6xREoczYBW48p6tRt8uiyFvrHZZPKrn8T/1uo
8oe3F1gJecWNH2k15h5an3kG/9YFe2U7qKJFl5l5aVUemlWFWHr/sj0CssI9
4x+1sn9Yr09kF86rkMLbnM2T6TNDcXQl+ACHEcha9RBurPe2VbHzxZQVP3nE
jDdWG3VZI3Cq81UG+XmZKFk3LbXPelwCTEC8PgLmtg/yEKk1DC5uS7PyjTGY
Xj2mESKjUwBfk1u7Wd4rEt8/+XxQBxX9h94f2vre6P6KPevNdC3U/vjwnZpn
UvMxr9rQiPToVBoBZYrP9XpUbqWBmDXcH5Gr8zRWY0ikaKUI0pbNW2WwHNAj
CyPS/XB8A4fs196arPy1MoG9gfP9DhCPJE/AO3i1y/swvK4iQDf4Brt3s4/l
CtBFGoXOrmlzrfUtKDFLxlGXo4NfffLkYOCpzb/Q533LBksvtGnFcDAc2aHA
pBRFcFXM9JzmlzVa7WUgyZVw4WJgERtqsNXNUoDSrRpkrXuPe+IDWAP6kz6X
2Rhtol7KwPrQabiBTu7fnoIud1RfgJSmStL+gh9uqa0pmGELWk+I+KdoXOwm
SECBQEbtDbxnMwWTmMoik2PKMyEE85LLXNfTs+YNy0idtihQJgpgQP7Bdlgo
9lrMaKPYErqFsW123hKKbksNH4ol8MNAmBCrWFoTzvKtzl0984eK0SjOpZxP
2G8y468p+386cqYqiZLmbXqMrBZoo3UymLMNtPHFG2Frv/W4asE3uJKWpERr
nLDxwAgsTuEolROZid6SHDAin+Iag+ncfR+mBC8gv1M+VZ8hL819lm8oJsRE
q/pO+oaDargn16BtESXTMr4G2jP41cZadFAqFUWPlkUw1yLZIc2DUfC70+MV
BN+myWsPwVOyChllj6XQM5o4ADwUKpdjbiioD+KBx17LxMtP7JEaiCQA9bU0
8SkFiSIXpWJOK3wPy8R8w7m5mlpeMGF83bvGOGaK0R0NshaUFETMUb2u2dYD
M/jVLho5s4Fr+IGh3e7HZ5IXiureXk+d7AkweJNFRpJ3VcoLD4T55F+G90TA
/b45+1AL0yeMQ35BIGSZgyuESc6T2lW2qo2bAqSXLipaVh4z28EsEBBn43wm
JRd9VFgJZYpVRsxDwWK0y5kV+O6FG6wuO9gb3FecWXWjnTWk3IF/nsP+AvCY
8hRlMoygPvZGqLl2R43G2BG9M43/K5tsCsZVXcnHZ7E1Zw4+3qorBM7iFt3m
q5vTyzHIpTWc3MelS3SUq0isu54dKuSMRisGtM0l1YLiSHa3L8k6PiYmF7Fn
WxGUt1YWZ2tN2dsYuRPvpKJsluDBMrSjlFYyjz6qc2x24y8juiirIeKG/eP5
abOFGXYxN8Y8RfdgreBxCAf4LcFkdIbS/+UFUvoXZ/PVh/8zbJJqWE+4eo9v
Btty3bd3/i123r+EKImA+52p85yI5tnGiyjTnTHC2wjhVk6XQi51uEOGqYQL
yEgAVcMkAC//0YmNjjQomoM8IyJB0yxqUQWe/8NHIfr3P1fXSeDA799mb4Bx
2gbnDcIUiPFZ+hu7V7b+cbiYPPtQrR6Ge/52HNCgehdBq4gPiULNvBTREdXj
nfck32r7LfyQp9Y2rvn9i/CLHxpk90e6JAFume7P/94fnv+9JsGAhwdFuUzw
RCGXKYHHwCA/ZIqM/hcMqyyQQlJyNJ6g9V8haTuVqgfgtoj94eoadM+ollVW
HCC1fucul/Kea/RHCsVRB09r7g3eZIVohGu1cjFnkV5zk13mUq49465IYDmS
jy66uDNZrXT52GcN0g9gSAF3O7Algs6pP1W+dY58KZ8BjlAHJho3JeZu5Tu9
uqyeb0elelDFb3wQmHUOEh+Js+ib4zBZD6ofPDesCOBS2yfp+ofbnLBJxYIN
8IwZVGesDtRxwAdSu6mb1boJ1qSALtP5giypBxhnqIEa9v7na/MXW5NtykPv
RvRRgcdQauQKjNEdF4gnhsyUrtLyXOYfXsMN+QauK/Ilv7yS57vwjABhHcL8
t2qqzn637CpgB82Y00McWsHqvVYrRIs2PjrvvWpgfTsophwdwCVomRyx/IT5
nuteUvJd+ixEnuicE7yozF0KaW6+Y7OcIUpAGPe9umNmQXQ1/9uUqANZVDDr
cSssqVPTX+Gczan6DkN8NdXgkkQAPIb6Rmua9HEh+ZvVBLogCTLtOXuRDyH2
axytGbdaeZGOicfzK9/ADmQkJ/9vSCgQc2TWaTqwNRsou+GHkvQkg9cNH1vJ
1oIQBiyT2U5I+ozERxrYq1WHU0cpPqkOXVaDxVrVoXlYbBELNoj7rKv/2vU8
mMnUnOEmQ384DtwSqiqBSaz6+75hZzqkhnt44W2S8c+b/1vCl9fHk6fxLZWT
CT4Lnuklv4YNeEY/AfvQ4zV72xmuVh6AKjck2ukiw6qHdybJ7fMeU/U/KAOM
00UWB27FLx6Tc+yLBx9lKah+3LG4NZxxcoj7jgBn/n+TZilPQfROLQmbUrVA
qcJgRWfwHMDU8hS4w1F4eb57jiqdxurCSg6AuV5SvGDp0P25VTKPA2mT2uX/
l5YnY9uW5nWT9owrLdvgSvMgNsR3rE3/p6yGNL6OcT92uk8H4Sa/lnvx/eUZ
DxDKG3VhV2sF4mxYODiyhro+UOzUTroq1F/SKJmL20ZWeV9NEig+uH3tqqdl
Jl1WPDsTv7skw31D1fApM59IU28JbprVK5XFBMjLr8/ed5MaO1yc/LlIZtAU
VwZS7XPkQwqMxYGz6NsO5oCf5hWB/cGGEAZYcUKtN9BR4K33MOKBonH3PQd/
0k66nCj0crGMZk8fDQ8rYklbswmREZc9kSqfnv/CG3VMdQkb0yO39p1YXn65
L66wd+9jJV19GRLU1AX400Bf1qUO1q49mBawNl79KH3vhb/irR+ZUb3mO81X
DIY2/GC+In8zDdoBnLSUjETAsOnw4e7haw9ntKWWZ28gdmNuMmfjkulk9Xta
ykzTt0JarCYawTfMNFJAEqqBTJZZycwgB5k8XrStPhBtPGj6Y6zXi5Jlps7R
6hbUw6yR+fIHmCtjKLAGfFRDLOmW7UYvvnLH4NeeOn5eAN0ch1II0elSlvT6
H5qkzafuUeJl8Ejdlcp2WMbbBJo4qkmbIQH7kaIDVrvYnuKfB2ss4o+x6m/d
Drp4d9RGpbgPPl6SGA351dPF0hegKAFsjXAH/g9EgT+jCZYZCJ9zNSKp9yhW
jnXI5De0gUN1YMn1ASyLCr/MsJQ8QYbIBYpYIES4NgxHRscvOqW0R7HmKZxv
jG1zVMrdB50iIY9Q7gd//EckCc9Fr7Wcmx9u2/Onaghy118RST1wh8oMKfm3
BB+yTXRVjQZQG7L/3ibTjZyKZQuG1wK8WKp7/HCpIlPvuFJCXriF+cJ2SD8P
liMzoQXpu24btIHlbOLx3klwNALNAHziPkbHh3uktcOFXsu+eFxvFxTgvmZ2
2pLbVbvWKG/TUEhYpxc2ULzdlYc/iH/1fbaf9wWzZZgnHJ7X0rC5ICDibTuz
Ptbo1/6Cm9uRl+jZ5cPfT2Ria2LhElJcbP87YNUYBX0DldRRZnhbamdVNIv4
xIjKtYvA+kluSE9iLrs0KqoPQQt793RNBeAPv00go0SY+qZz7VJU0fdwRDqC
jNGmDF5aXwrsJJL5g1LKhaFf6CvK1atMZkh66qXI/w3Ej8AUrTXx8F3mMteg
gwHElL12OJV4LQOGtsPTU90NLKQd6OFHT0tTFlp3XkmjBix0H2cEyY6y19B1
HqHnJqyEmL/I6Wfqg2LamyeY94B8qo8hrXy1tYmj/CxUW23tZZfUVP5kr8He
p2kS3IcJSQZkB535vlBVAK2xaHLMs7GhauucmAcMH40NlvJqVRRlx/a/k76P
YA/iKF2Ql//PTSrYptQIrY8MDAowosdbSMUeAE1cn4g7tnrg+5AFoRjoaYzv
OkuVnptxVGNjnvBTw1uNmtZgDgGWPXVTej+oAvZ0lh4UxpepcMPMr/M9QZiI
y9hjtRiNAXnZuj85r1bLofg1NcU8w3HH9hdbf39s4vE3CbdtaX8/vXbAYR1Z
bPYH8L05mp0PT7F6rcotOrFzPDVrLVfYiJyLIN5mTo7WVLHXZ81tH6jVe66V
U6PPaWWaojvV74QjRiZ+uppDzYaLypu212lRh1wSfu6HoWiycjhphhyLrwSk
WMGbtXHnatSKcE2MrLI7VPBmsOaeM+FZlzOtRRh0yMuUxIvnEF4eodU5gOMS
nbKC+arkLiticJqHW0rqsldXzmaSt9r+VR4Siyfjxkwxxb9XFiFV8G+Q/owP
J5OaYOA5nIWDrdvCD3S/2/WgXDA/Xhw6G48lyrGGjg1JCIb77smeh011xN01
NSuYNLtEPYFH+/do9Y23JrS2qddW1A5W+2/2eU141+hYt+7sE+Q0XWUQsfD/
rwkm2EIxuYEpjuSSu+UzABIe1gy27VLvXy7d0MnmddkjBBCHhc0qUy10ACJO
h9OMygO/TELLeMl8lj9JYz2Mmg0AgYYnvZ0MpRlIhZFRb+nIRSOVSacrfoDb
5nmyY4vkRciolJa4UAUlJ1VirRBYFJ8u7qIQUy0iK1m5DoUcpT7qRntOq793
nVX8hE/KD1L6wVx7UpoAnktc/OGzk7HUD47VRpyvX/Ux1jMlWTw1MyHSv/ww
4j5nZ8Xw+4xR94rLWsPiV6l9Vj2v4wvZsz4s4lt3VpRFHDj58Wuu0LIOl2gt
8ltAOysHJZwPbp3RwnELkCy+YDb1hFU9RvW233miJK2WXOhHMoAwd7j7aHpB
XNjgrqoci1glQjXIYxm+W3phP6DIRRi4jmpm88qFTeVdt67YfAJQjLiFhv07
oMc+uNS9TjKItps48jKeF+2K2OZwi6Y/ZlTWgcwnvwaXVIAjLXCUa9KINdi2
u8Za4Yplcki1cg0Ka4w20QYAUknn5pxHBnHoAANXWm0TOEyBHshoIKN8OV6L
bTrZapKaSe/Zn5cRGAqjDYCCx6bqYsjT1Jlw9B9ID7kC3YvCQD1f4NqwNVM6
SHZnLIjkHlktJorv3uPmb35jSSebaAHlSk4yu6XJY2x2bQQh0iBjU4X6iQl9
PYZv71DFHb8khP31Uj2ZQqYif88HjKqIBosZhPdUUyinXZi0ajtLk2Y2QHGM
X9lOHRtV43oVrlI9umabW2+jd6LKX3OMCbzeLBVNGyAUCPLU8rCuKDgdZmGW
NF8YjaTuI18dus3XfhThwGeo3qtaM8bvDrBf1aXga4OA1u3k7vGc8SY7pC85
jXIyZxBSYlQsYyHUDC5HhxVb0R9JfwzyimRY34CR6jIClqzRol/iml+CdlRo
Iw07NMFgGkbzHClThN8brQNxyZSJIntJ7uxUGiUKw47MJN9S5q4hq5PoDusU
vnm/Qhfq8pFNN74iQV2jhV4qs0DqIdLVgv6ybqoNtZ1/a6xSrT00KWNAJSCi
97ifklIis54iDK0BFdSsJ3ooPVgk69IrxjyQ+8FhXIOsiuyQUIsZVUVIwYcx
y8wMf8kG3CS5Ec7WbRaMUE0VQt6QEuE2W13h5ouGARqQmekfFVQGTuH+gsCs
WIdCK6vee85ZiudZoY2mb/e+tzzb3m9MhnQW3JfxDEct4XB055pEkWFFgwEs
9aTGtqqyiB0Qzm7vAdtcbyIy6UI5P7X+B6imxFfGEVSWXFpmJHPVvh0mKkEP
/IPU7bRbrcOmXih2ffqikL0Y10GIV5sZdZ16RIIr8lO78pfgNEj4qyWwZsqk
fwWPDzaA1SKqLi1JTv7oP+Rpn6FAWPnjVQLSBvayis6v5BuxQTo5Hmv63gz0
4mxYwE2y8dYq4Jey59L2nPGf/5fXzyIpVXrkz1jNsL3Sbr1iv2BJhvxCyrMM
uJkz00aTEsgWOcFdtN6zPCJ6hwDIIOObfWkPEbPEgJ6X0D9fCKSS6Ae9Tgyc
6kyIhxRV7h7DaHPcZH6C6qG6vao9J1Maiow9sRQxZ4fwllKJBmPQ8KQMfnft
e8mMIdt6RJ5OrX9f4e470ZSvnmG9xAkyVKkL5Gi11Tck46Oa/FWqmolkOvq3
6WA1LQHsuUpVbOqi/KrN+H6GeO3xLcareiAXeAALsedo0BFjAYJcoRgQKPXD
yu8tWEqFSz87J2FvhRKdaGRWD55thdXRFUta9g1ItHaaob47bQXV57alGCcL
Bbe9d7KG/Woz+S4KQQhz5cDkmTokfm1RNwUvDKbpZCvgkkoFdEWBknBbkXSX
nKrG+1f4u7Z0dmVXdIFoyqva3EYidwhOLOpcWamWQni+tkxOfK5CjoeAIh1h
cr3Bnaz3o67TYaINoCpRl1P4re61e8+MJYHWceZks7DtaASGcRjBXtXYyHkx
hS5DVpSXd/ImF/y/yBx+hru/u7EzAqhuPBjOz6Jb96H4dxFJyOsTZTcopGlH
aLE1IgFc/yVQT3gVmXdWrY4aGT0yF1CADny/zw9jXLN+qmnbHKKO/0PExtTP
rCDKOdC2k7jJhOkD3VxhY07q4RN4lVJTgCNxntM0sTGW5MguGTl82y9sV3kw
fP2zPyVtNha1/xyzVqkBY/zNwX6z4tcLPvpzUn2kwhdlbzmzSrTppcyr0i/l
5KCZJu/u7buDAcQTH76ZZ+ZLISLCBZq6hoqz9NfENy9pmgLEOSnvnhIZ/1JL
IPRtIhdqsUVE1cgv9JG/VYKKKBIhEI1bC8xQyor32aKFYLidrfX+jPDNNrdr
rgIX9SolkFF7lYz/UfCc+xinz07peRmt8GYKlfB0m6UomyhNJN1IrzUFvfNW
aphDSXPlc4PB/RDs9/361OCR+j4gFrxXxAl21Sh1Kv37NUSd448YDdnHMc/L
EwnGKWtHtq4PYh3/UyuX3LK67P/k2MdeJgD3AsyY0QDTFR65hPthcxC51wZb
KnxFoilIQoko9ImSuRWzp2TFCON4hiDUcy4P5UZe7rsVMmTNJMfRAZgm5wgI
dNBrv+A82oTd2YuTzk5f6s0plpObmmZ+vm3qUJfvJ/Ijn/Df761rbSm1d5VJ
rWd2yezRO9iL4qK8BHXIWlqYqfRe/n4IOkrgDrPsAVCqRllxKYQUR2+ru4Mf
Rg40byHFdzZWj1hiZdkngTPPiA47mKEhEQPdCvVO+D/alhOgPO/oplJ7q62y
sCvhu3KiMAurc5bCIjegSB/oNnqTu1FJFyWIuhfVd18JfywPjgyxjCAf6rDU
aPiMSCCK4HGDvCCiEK8RVldkrA/sS7lYLwc3Kn7muqOFtfW7yhYDGNyvJ1ld
+No5W5vj5CnEGPAfkpX0EpByjzkJ5yLp3uxXsDdRRWZ0zOxuEyRsY+DUJ0Vp
1kM6xoMObUDLD+WstbpUogeXj3IrIBvLUMCIjDDuA3EnrUDU3ScpN7+k8lKx
4q/NFJ+L4k2Jlt0exBrxcFG6QpGBxLyCnTMdXJZGxBGBZrhdruWoDeT0YDc9
d1yKnXDAiKOpjeJ/l/sxsCCbLvP5lrJV/zYiM0G1oHlDwYOa7qS7EdHOILMg
3i8+ztZawS+qz/O0c+7n/aihPygE+6I3bza70YY6qCDxgYJZW3reWxH//ZvR
d4p1JT+tJBrZzq/+OYRFakEygQoooaipTa7HJHw6Mz9IpZQWFLVN0w6dPg23
Icx+TIJXL5RUU4Us+O7Ss0EQFcJsovpmjU8FCVhfXcmNuoWPkRUEuVPzZQPB
QGvEasiJetRs4PvFh7HtxFXcvO11DD/51SrUWTi9a7JKOfa1jnUjZiD1OWzG
8e3UZ2fwjl82hJDfJUkAl+GRSyAszymglomfbyF4xXO31DAnpYVQwbWeRGMR
vsCvEPjr9eEh05WJfEQ4qgnZksg37RgH8s0VrDaouB0iXpvE3dqYVhelqL33
zeBC4svLtoF4KD4Qh5V0ch4FNVfYN37/tKuu+YhKmOoRXWEQONKhwDsctrlq
GsGrF3xZAPMYzrWDCMtYFRySnjMAkj7JYnN0LrXCvpplmAQBgpk2+GAjgICz
aBB8AcZYPT23uu0D7ualDvQxidYPqGy5fTtVhmgaFMiupZPqKPRO2XUpvl6U
NYdot1paG+JG////BSsZUyBvZb7VRGNjAggXgwPr1pKsq7O1C13Q4VIjhvHo
0qnQLTBR6fQGKh3y7uTrt8+Q6jphxtKk5R0MYzNiI6LLPvRvWhNhWQFestQY
cb8SBF9UaITtU2e2bH+X5+dQkYzTbBiJZ9mSVNEUIWbrLSKgIa9/vS/6Zoyk
jxNknoZM1Kd10jqQ86zPPm6LXYMrTIqUCl+5pqbYosypm3vMv0M7t27aJyl0
rSFBKCFzwpojqqvxWj/ic491zDIxT7fpEGDmcPFVUFEi708kP7q13vSSu2RG
1I1ZdUUkyBzPMiwmDoKReDzdlJPdACC1JzljQG6UABMzul9wnFN/vBhUzptE
VKlGCO3vzVDo1937gd600+pHYTBr5AQGdirMHlspaPY7wX3pNxkchSXRcoR5
2A5u/LEKzdfqMDmOVZz425XN6D2ZL9Ha/VQ/N73KV16T+t2E4e+fZHmE+rNe
rxiOMLUHUUOsmc4jXg+vkNiS6xfCtXRp0Xw5eNtslSOtGXJvn8OwHNVe6gXx
/BVWPYal6ckgfHc0Mp5aER3SeWy1vTnobNd+2sZfrlzfn6IRszXQ1Hxi22Mw
GF+LfsxpSyZPY2qtrxNYxyv/oH4TOKEBcwyEfBTpJezOgc7NP0s8jxhu+owr
j8aVi96MJ7Vw4JGIVCh7xeCqkxHnEXcmamIfvqWjrrcg5UvaHOmARmIY2Vr2
XuNXF41Gc7P5IEx5iQ//mC8HTja+XvD58NlMIjI2LWctkYJkkue4wz/5ibcq
efpNi8n0ckxXLtLdd3k+E0sYuvc1DU6bFHWj688CJ8r8pyY1rdaRxOsKt5gi
3UC1Ku/p0LcQxQ8Gwd1N1qEU+W9qL74KthaBZXtH8CxqIQuxBJzMXiLloDx+
TV1kdPiqLdcmkN3OGF8I0bf95hpJFThe2H/+vkOpeebChFvTMSEuv447cBgG
yts5oWEY2vUfEyQzsBU+hRQnvFd1ojLoHoHQuy5YY8T7cDIsa15pnnIv/x9j
AyKeNSQdTm8Qha9g6qGVjGHwAd3fRcAZRDNWJv8+zkMRTQW0zHlGapXthrAq
VyJ2txnMP5F7FRv8kaNXwDQLZfzBaSc4Y/+Z5r57if9hv303LtfTfapSInbd
XTKynVE5jXMxd5PPYYUZRXz4GhCkJlCxHaTgDlgfdag/NnXp9HBw+08V1XWX
Q7mXbaaX3m5ybnMa+FVrJ7rC/jpCgsKu4tv8udXU57ZGmOlo+TF1mb48jWb1
IdczFJuLK4cfT5Epp3sAXGs461EYkPIERm2n5zR3eYqOpS4J4o3DrcYnCz+k
OqP3n/R8XeiW1/jzKkvpilcWF5S8V71i36PiCiACNsys9ZWSs2O0f6OSgqhE
IrqXC5KAXSJpNFReXLdD2B1gl7uNB23mPH/jud6gT5tJ3ChihNuFxggsTqsh
boYvntJrwd8QM6/n7mknK2LPeWiq3l5Q0JrxBPHEBDgUji/CihC26jV6SotZ
d1eX6chCEUUlmIykAW7PFswrvRWQjARcY7GaMgiTtdC97nLUICs3T8l1Xi+p
7GxQK1iJbZP/xig+ttSqB+S/ZrUc7CDd0UBNFUX4bIGH6Cv6QYMnQfsRSKku
FKZat1bZ8oBFNk7PfTtbb7MHv1BtkilmXokfClY3AXgesI+uAczIXw6TXMqv
EkrkZPMWg7BHqCno50zm56Yr7AwPq8hLereuMA0ptBHUD9oBS0s2BwXihN6F
Yac764wHTdq/g4WDFmdcfshsMKlrrBlQJg9CxA71Rey0Oww+LihksYsdx/+m
tPq52msnUVJIE4f0BtYHBu8MzRr9uuvL7eW/yvj9e7OKYdHTa2qdvMEg+yG+
4E4h9WtZChKeNztadCCA0sYpvk/QSBIlY4AqoIousMzWRmvmF4NFBgouUhN7
xhGDn8PrqmGcqCCmDgrpDU7wkAwfz6Pc7xFD8K8Jqt+3ABUe0PwSGlgdBTZ+
o13pyDaeY2RWiBn4K3MBA9Amhnb/x7+WU69Vzmok4kK49af9M5jqgzmNgBXx
rYvoc9S9+GwNtWFvb+AfGF/0zLi360KkYQwgFflAxQfqkCf9XPwYFI/Cl8Sx
blV1FtQW5wPZo8k1kN1XgbZ/j0YxK1q7IPS3/r7D8hftOakGriz/Zhd/tEcT
meZS1KaIJfIB8heIOMN7uds+YljFN+jr6UO9pC8F6aPThyZu5+VK9wb8ajQF
yMjcArDR54mvXz6nTmVEXiwajkGp8VS3CGus4t1KiLeMdDYuRhBPNUJ/Qcor
C42pXK36ncnHGxi20gruVPgPU2L3V5LnGjQJ7G4rtglieOsn/rGl5hUz6Vpm
2FlHZARTZt5WGyjYmg6SO8YLQ86B/WJYEjiBjAFCGJGl2HxTvUh3p9XsNPBa
uXmCynhPvvTVlrdzRGXaZcuetdvCZQzAb080xkCRg0ShxMGJQFb4C+WtdG5K
p0qT1vZURti6F4Q0qNT4EGw3n8rHcE83us/hVfKotntxO6+t/m/o/N0krgFU
nhfvZyBq7V0Jf4SdHIFH2zcY4B50HRVBhmiiYb58RRoP/uG34nd6x7j5fOuP
HpVB28gF0ojvYwdcdw53MZZ79PGX2f1ENJVKAACcD5QOq3TlRCLi9goAoJSs
vn55y/7h/SII880IprBnxzuf4wJ5XuNmGLtUsnkOhuo/7fbzkeurTz1aXCeG
4ZEMshaUcdpBI9HQL8tbGa19SU4Up0BTkx6BV7xkMBdWxijh+HdGHW67JFaK
hY9wSkKQXV6RCWW6K8deH/35fcw1qMMTpXHxDhLgU+3T7ORhkK/4BNG3mP1N
0GqZxFgJYaX6xefu3kyMTHyDwp05KbGSwsrYtpmFWSG3pWDXPhWMUIPDVo1g
oyv0gxxIHV/SZNdoT0UKzJ+TWMZTXU5iVp2P/dqj6byXsoX20r2akIgnl8Ym
FT78yjxLJqtIyORvOYlTXUEyf5aLQOtIWL7ro50AlfymYmKJp3j9WAJZB8cC
xn4q7TTdDEXLCnkqM14TPlU21qZqsi9KE2FhY6tPU0jxgoZNlgH9HMkHHFRn
f6bSSxW2de0YRgjGz0QjBP2TXbEQQucBz+MyN/h9nwkXyyXzozfoVznxvpc9
hb91XS4kuMyNFNedf8IqbNnMz9bQjHym3yb19MVKcHK95klxUh57SaiEOPrh
qBgIWF3JiU3gx8kT2w5/M3fp6ZXccxBqdkAKzeneS2SVRVf4Zx6jIuYu2iHG
LGlDwUt/nYTFqS9Swqi+9abr4EkvWVsgnYVgxEBoPZhXtvZjEkDI38TpYf4g
fC0yHdn2OBCTGg8QzDKOLzztLclZhmldZHlG1X7qYfTawtTE55a1r7EHwNvk
cw8M03nOp8929KpVGtYAxOOOELc9Wu1zdjAzxcie734GKwE1PijYCxUHL8Hy
/l8I6ZpVQoBPMAgkt60lCB1HtVDz4BBtcoJNsPg6fQvuyrMuw7XkhdPe40Qs
CfI8lXwWNxaecx1clj9VLeFoL6NFO/8F+1juW1J0orBSiohuvWxv1aJ87goN
9gSk/jEXbVzGpaIDKOnazzi7E/Zcs2Kw4U0v2y83JoFbl3JbDowTP/yDj7qq
RIgONyQ/9CvKZuAS6Vu2LFFSTKGk6IY43yxR4W20ndBmIGoYrU+0wFlQkQTz
igVRwcezY+4wM5Q1YOAs3QKwVOXa3Feb9AnzDwH/fi6sbNySTS5wFtAr5UUV
YbXkFahXJK8t9xnMqIq/EE6VKZ68C6saN9dvhGCfdTIiO/q3o4o0HgZn3pGs
Caeht2P88xRwdKuaa6vPR0RhcMIpEewA6Of2s1i3f0rBmSjzT76VS2OA7mTm
4POVmGNc3WAbNh+Whhc8L9lrZhpp03k7ys6TDcnZfV0/Ja+4dd+g3bNRcTXF
yT122K+k7Jttmiyi/knLcl8o49SCVIfhB40Rg6u1flI8JKtj9SNuybAg/T6s
HtbzZkavOjZo9hCVaVuIiT0WSJ+ZSEfkhaioGNyuivH/CX6AaKY1Q76Tl3cj
niVDmsXivFoMXEH4ft2VUECDmX7lln5HyDpkdASHKndWzmU79V9kC4AJ75DT
Rz/OWq4zXtYduEWmB9QFE2lmE43OHZ0CQpfyvMtCNwwUCeqR+Gly+OSNVI/x
8I6D69lrjN7tYTSqzBHZCn/xMo/7f8dZJZUh8niYVXBvqy/bcWwMW+93vZQ9
nhPIoZTmuyH+b4VYBTIk/FopLgyPz/arqxRawaX0SBm8yijc0qQic+F5yo67
kBaWtF8ftPuA5qVN8IkIaNYERIQkKnCmzRRbT5PomQNZeQvWmTG2gDtmb/3v
Yi7kc6pndT49hYGVQJAJ2RLV2p7fNuAKZGNTlTkwjHGMMz1bGv7KCQgwtxxg
o6oFEIeXgOcXm3YrHeOiPcD/ZYq+siRasQxex91oiJjdIPYZHW5iU+RKYLGt
IyrwEGeovvRMeQGhch8aOpaQs23YjlNUOv8lro1TeAEg2119r+ohnlG99pMO
SeJFaU6U6fHO+INZgylc4ODaAPcmGMGlXGx+9ZGz6SgS+6dcKfJ0HEV+wjHE
To4oYI1ZbCpK6c951kAWG4qheJ4PQtJh3NoUJygVHRktkPGlDR3sTzt0ZhlM
8TdjOJ8rHAgA6HR5cipQWF2CDuLFVmjI7oQVct5b4pGsAcnn21FPfB9msjxr
FC7MvN3JAPj++YDdOw1UpqaR0haz1OxDErPkZ8n3Aq71/ampzOGeXqxtx50C
BFGhHmatTfg74UgYiuNi1UiGiq0TmSQbqQufeIn/w1EqFq6BOKZlM7id0ICH
IU0ADOJ9afxth8YVm3EURXGiaiNl4xWdWLeWUEj8vWfJg6ypP6CFxThBWLtE
N2Eb9qrFXonOP8LUYKPkvDhOHjOo+qaoexwG1PA2seICQzf1CiKw0Zy6L4GY
0XUkkk2riAuxnjxDIeraV6voCF0bqFGdz864Fk4FlvDlN5+i9MMu7XPLnvX2
u+vBQ0G3bg/oSvs4C9AkDm48nBpH2zwM0CWjLfmoDxJDT0WbT1KkUu8iaZgF
ncKIuH9lvMf3Ap9v7HsR8g7PZHyRGu3b0ja48KwiCuPd3JS5yOzl5cC95Pbj
VBEQChOtMvPCINR+AUPA6WPdC885JUnfhwcaHQQft+yu9XsYSeGKtBdum478
el8xAM003orgDS4eKHnyHD0cUw8ISxW8CwGBkWHFZHbgpMngk+zp0wwhq5oG
xun975//vm6/bFtqgXheh+RDe+7m5qmVsfQE0k89fEkHcxzP3bndbH24D0Io
Xo7zX6kc0ZFVlxTzd/cdNlRBsmkNl1IAW41FzgsCpCDTKOMZOzOQiGyzUm6M
vLx1Sh2oKJTNRXDoiUT3ymi+mqsBasV8OpqwKzzwVQUAwn73ZGXTxCO1YeRh
rlLO6G0KcCOHUzvfcxQF292SaRRz+nhDiSYryNtfZf1z0M9TB5f/8a5Wsv1Y
YkMk5G63ORMzd0BOCoFRlRjv0nEbs9rfRkJqE7+3+ObkG0NVYq2mMLKbpiA9
fawTwn61WOjPTq6pjilLa4hQivriR3ZlaO7nwXJ5WjT5bWGZVwGMLL6eIS4M
Op30TrxDiq+9ezfuwCbkJqTScp3Kqq2ZMJQ157fqKa8mKXsAzrYu4lonXvnd
ifo4ANpQt6GJ4KqzICDXyTjcbXR1APusa5AkGSedw9WT5GJnqz7TboJHZytg
V/KgrPAOWfihjqQn1NsXa55vb+tbuHP3T+dLccZ23UxgTXMsPI19HW8fDiXw
9i0qYdDWqBe180elerdJebYg0wjXyrqYhETrOexvyp3Gd4EmhIK8NUB9pVZg
JrNPrkS/2SVq/juu30Q494vItA2R4bwZZZ/0JmMJkwO2S4EmbmOzzCTLF6G+
gY6ibVdIWjlu6OejIn+G4dgJzl+eKy7TlEQ4U24F7BkmPs7bKUWG/RpdFR+o
+dbzUIcRmjfo/jWFD3eYGi2Tb5FZGkORmI7p+BGh2S0W8fnHXgG1nHCIalG/
00Ll7Jnw+aZ3t2IKelfILYEx6Ezjj3jZyII6XhZQDTdLyi9MvhiYwUOvTyJu
6i+5j3ISCEH2Vi0DACQt92+miz4GvTetlstXAJdB5ceKZUBgiJcbJFot1RJD
B4uPXutj7/h+bSEc9ED8DYS27I2iDVuZQKfQuUaL4eDCzFwdPEFMmEMRCpQT
AJctzYMlau/n0VH90fhTnwYdlX/FeJynwjZknZ9DviGl+9UicySSNfqKCl0o
zu0NMeo4PRb8UB1wA4t4Ii0PVUizhs9KugTlth44OiUuHA+ul2TpKq5PNsHT
+o3OdJfTU6YjuXlyd9i6fKRXBfOdViEaJepxt8bWztrj9Iv2N0zzv9mb2kaO
DLS8GDObFgosQHAw/d5crXritLU5FHDr0IKSCpzYLULiI8Y1zNlHyG2954Co
mPOT5g3tciEKGvQ/4ffDk6SHqrO+jsyitAGywl+zpx+gSvaj9SPJdH/CLmIp
/IrfnzzILjmfzvO25ee9c9moDnWWum7qw7ZVYzzT11W0Vr9Ok96KS0TwJR/9
fBawgG30VbSKSbMEqAWlMGzmHc4BCsRgGMtVg2Os8k/9CDrwjLyJWmnZHzdh
8V5BIPf+2oa9OWODcG81AinMQE1FR2wl/rtOHqGnBK+Z/bIRBadUPoNRDZxO
ZKvJH0+yJ0wBd+/+n985KwTjVOniIh5LucawLXbYiy6pf6hqPAy3ycf75Dn7
MGV4+oSOVGk8pR1QGUzeGJEsMDIq1pmc6TeLbbyvRyk82tVByhsZegq6706r
wnR/ZVKgAZbHPf8CEN/+5oEVW1FVMo4MKa00qS5EWMbL7myBagTO31aA6KIk
e05A56K0ofYiWyd4HxX2qHlgEXfW5Angdt4R1kJbkiBJrrqChBfyaObzYCrO
vP2L095FouglnSa3sL7CzETBN3HL+DxHSRlwK1DDxi52MfFz5+E4nrD657sE
OaQa1Eke6+Yhtp6Xfdasn77d9PVdEqyT64BWt1UUSoeZ6uGChjsjUAReH6AA
h6uty5Cf9UhUUsMElO9pC+pIzx6M8+LO/cYF3XMhO6uFHl4bjHsW++aeZema
IFDrSF1hiAU3ZOnSchmyckHVD8eyqZpujgfMeIDDiOz/GDos59xQCk2ndaY9
7hZsmvlZUbzORbjVAau5wsV3uQ2lF4Qx+UHapVKlkVYzbRaBbJfmF64XF4Ln
fm8pUgwZMEM1GJ4O7U4oNdz9+4tf2gZcgQ1nqVBjWSIKpWF8HKvlyxAUKq5i
1eq5p7BPQgKQyx17A4crKY5cvG+w7dPXA5pGD28fTINxRO1NJGI75r581g4K
cx1fYz8wf5ZSfAjYa39R9XVQt8hZl2vC+vloTUVG4Gfo7yOz/ySi5L7Tnyb4
NoixvuXmw7/t6iXbQl3z/F5BLr+56jSBz9sNqiflTpdq6CRCQK1SdTPqP+pL
RitI1fZbHH7Hikg7dG9A3euieSAKHsMT25gt04zEqHeBfTOJb1c2ryKljTu8
An+aH0LJbneMaofbRfvJSW5qJsd8e3tHOW++ZdaeBmj62NpY3rktr5a8kO+M
yNQL+wNSDbpJQw+m4Gf49oOR5R+L8N3guqRGALg+5qWWiyKZ4cWxO+wrxWFz
rELVlSjqkg4D4J6j/BSQvWI0jxggETjlHJTt0E8+nd7cf3yrgp/pSWJXo9NT
4eH3K4/K0u6p0JHDpcvvBrB6IAcSoB45spSUkV4OvZaDkXzj98slqW3o1dGY
GAm2Z0JwsPrwzcS41eSv+RdYqOF/K5C4Tke2t/1Jo/+r50MDCkhNfLV2QL0j
a5954IhitwywdS8wnw+LKV3bPB6r+vhQH5N8HNmeCb4hvU7GHuvBHZtDvjmZ
z9Zv9pYqFeDpGDL2QY9/7WVXGah4YvOhgNmgi3AAK6bqp5zZ+zLsFfrJO/DW
1nDs1/snr0DvG7ZsKVIBK2Z16Wc2slEJS92pXWD90gOfRrQpkNa2fELNptUc
1CJB0G7636B/FHgZrRqOKrHavVl6ksVeMcojaEdJdCQKXG8v2KQv8I+WG/mo
U+Bb9/sbw96tf81SoYMJyfRggUCT4YrqUkzy01ujR7BozSnso1zAzLSvbS3k
LUZZkP5dv6TiOiOs/ZG/Y6ti4Pm6SQMxbZKi7sKYpFJBjLpaoEpuFeSEmvhz
j+v0dy0Dzk2UMsh9l5OUN6E1L44A1XEkfmifOkwBpbJCVlKFDXBXmZHzypy4
tSvpwDTvk/AkgVJ2f5HZCHv5pXVAFYB/2nPCj5eSAVcKxazjYsZRdVdVdiRD
39bW0HS5RDQ0gS4vj1E70fGYYX3u5net4lazynToQZPpunDhT01z/nzF3g50
ri4eFu3lFao5SCamr8viAIqj6+OUS8wwzWB2os9Ht3eoqoIueHVkBsHjccu2
3NU8OsZwtfACzxJuVN0UxJVCo9ElEFxAN8wwry5shWl/pOueA36tVhEOrgvU
SLOxKlJGYA3sJ0olql8Ux0pqjnn++kZmS9Od2+2k5BRQoIe+naLvLTSYijax
QB0WuKW+AMe6YJzvge+W6eaCttyBNwNLtV6tCfoGeVygu6C1/5kiBaVM+waw
YlkRG4C3r3QJ0cy5dbHtTIW69qHED6wYWgOYGo/vVeTMuDPkg1KpTu2yLlCT
mO7Z5n7L+TSMapdTPLu+/kUe5unVhYItgELdglxRepA2rkYE8+yQlXpRnhWa
FLzVP+7M84otVcFb6hElSA+ZJbZ5JuWkN7vOhecEY58Z6sTjr9ZCxLHY6N7D
oUiLpd9obxKrz2jBLdT05IVKs/ZJY/ixkPtgFdIo/X4oONQNasoANWC8tY7m
2gutZiB6YUIKo2a9/lD2G5gi1wort+D1e17CkA407LQFMQNRZjZWUDdEGPiY
Nk98IBpa4kBz40aKuoHem2vz/wXqMftPnOv98Nzg4Mvh2qlyPYWLjHEv12bj
nhkqsBCuu3ozlzJZvneyVWMu03cXTcz1qRl3TnFfBpSB3M/su2fEWHJKsrNW
+4kmTK+72Bd9DbGOa+VnIRXlrTEAv/+m4KQMXDSZeINQQdEmeRoM1URXpLIE
HpYpztcrZPkxVuIJjQ7iG6Y6QGMbFL3tlSTc8pj9iytrk4wdG44kU9TfpOoj
1pP7XW0G48ZWxSv9DVVoee0oUFj7NtYoTeNTmXGspEdod/qczgkufawLCNzU
GeefxNdZkGaJTS7P7KFF1EaCK7Wpd7xFkSZaNYurxttv5j/WREq6mUOcjVMp
RCD7ct8jrf7jp1pm2FPSrtlK5GAdVUIwXmd9uKIms5xXioVce4m9Bia50DeM
bjhbno/bzWWAhnmcbeIPRLwTITiHjcETCKG0ovb0TAX82DBSdNYLFfa3q4Kr
hgLW5LB2mw09PRiuZ2dm4n92AAG4rcXBHeVH827zZm1vWfhNHPL/gzVPWXe5
CCo9VviS/BJ/gudrjbeVnZ7u5BxSQqjJWoPwdX+20HL4SqKnlD1DhXeyPIET
q+/pYQvh0TxhnnOxLMm1yD+2sifWH2I1RVDXdf9uKompiIBqVukvh7vVryND
DPJ7N/pNs26LfIK6Qro8qXGBYEQ/mjq/hpZSz51KAr58vJr1DVjXQf9lTfBF
SZONk+GrhqDqSx018cnnZVaD9+7WsQWQWuxXLUTo7+BKUYyTGp4G9NtQB9KE
fF7NJz/TarRKVequfNhtEA3CNuItIx3e16Tlw3a5J4HvLq+KY97RfiK30Bd9
MMdNYYRt6uFstMA2vW8AagFRwp4NxPIb+D9sPw6e7dmPLrbBp61JL7WHrEmI
5Fi/FUsDN8zFidGj6mTeo0+lfN/vB5u4BgVu1vD1B4R7EUUwLLh56s3VhXxi
7FVdPhmgHHbN3Li9mSyzsMW0d3QCq65lcxZa3RR3o1tfT2Jhm0zkmNU2lnPg
WDbRlYakI2Z89x6SW/CP+I+3FF46S/Vwi6/AAaqVIiHicf6JvW6NVnlhrWjs
3SnoFV0iCV5Mj/5XpGhJqv60MPVyavxqSzx09o/oCmvP2iFBB219qhAGEk3g
KyxKdXnuC+9lB6M78isneec2z3sp91JDS/YdFZ2CynJRJzSZ+ewjAbedUw0v
WOPQnbpUe9YScGHiEMqSoUu3co2P4NqvWfClbcc/RX3ncBwIA6TGaALtJJUf
3k0i9gr03IHYJIVsKcHtK8LrRwo9zrnvo4MOv8PbJkWTGQ9GSR0jUbPn1bJw
0OZC57436/Tf2Z2iuLRLNMAbKeK8mkxhnjniLxjdmwaFZbZBgSiAMaTVl0cg
Jlap9zHr0VXalMJzWtfu38snISANKP1x14cTAF9I+n7RCj1wvLz7uxO0WOx2
OA2XkXFC26dc4egOgS3vmd7pVGUGHOgIXNFMTR9FccsK03hjGb8a7GBnxCCt
T97a7oT3W6LjudGRVmrqfmjo9/25ULIfryB3bIccDEvpRlRCaZXXDToSpa67
FbzGO7ibPRQZ4OyY5oJGHp4xklRsEC9B0SqksZAKVYfpHF+wUPz5xf7UsBkd
jt0R1hnoarH9haJ4YwY/Q2/7/kza7Z10dO89eMTfMd5dfI/EKNBxJ1/9C00D
NRPYyuyNqn11Its/FCWFSJim7JZ2Zy9cvimgKAYPUk7+CjhTdbOyzQ0PsbZi
bea3fc0ulHQfVyTMN+G48UhVcq2OBWpqZwH6hTRT7HUjuIV0wgvzX+BpbFRX
KoVbgtkRYpAlpm9PhA8cqx7zteO0dAVUH1mGDa2VXQN5usKlomquVRZSUSLq
Q55fWReQ1o5U+nQnPLIylqP2wVd6pdKlz3qSpB2UTWd+yZLMqey2zkL3ME8V
TItyBlE30Su3hOD3uqs+yzZYaho9M2DoADCjn2aZopXFoR442PrNGBPL095h
G5RtwsBvsyPVL5N8ZIQtE3aBsyCrwjQGjQnC1W2Vn1GTf1RMWOy4Nut8+4I3
uAlZyELkd3n4yo1FvFFwH2cSBbCMaw3z+Q5NuNdfqweCjHusn11226lr9NJW
33H1JA/r0iIocP5ZEUEJBKGiuJTSfqRVFn/83odwGggvx3pzAhFsLwcGe4g1
0bnkvHA9bQ/bZhKlh92NyOszmRtaX25sZLycNU2Luhkdu1yuEB42z3thO9i3
+1NiCkUK0Y7YSAfajqQy3md7RG6svZmIO7qZ2JTINxE/EE4WONwohWivcnvg
3Zk+N6+icr/lukTqvtgmutS6wGGKn8Ij4gHviJDXcrTNmnLVIFlfko5+H9R5
tHS2pRvx8aaxPK/R6Nmh4p0u5A8CprbdNZnSQYwG607uhEb76DeVZVtVqNux
iZA12ijTlFhymk0V1JDmnZw5XCuG09DRH3YMJsjP2AT3OhrUhwAe0l1M1+8Z
hGopRgSfPYXOGRvP/P6YBjzOn8Waya3uYDqnnWn1avgiInBZij+X9S8ldyUQ
puO8lRbUuQcIAYtvc7EWA+ZBVnEBrrIeoQPtQ4zG2LljKlaLvDjRMgu2h+2v
jWQRsk2WeUtCaROmbYAct0ZdpqU9Cn6aiwqa2bIihD2CS7ZZRPq5ziJ2h6Ys
4jQ74FL6NEJqaYbheDkE++QFN5YoSinWuSJVG+IHtvkSRb1mupdjdGlYMbUk
9cPp/uwJWM8cmNyl2fqaLbu5N1U1kD3EIuykdL5Hzt78EmWGiF87UQZehJBH
kP0g0ADPbs/K59tFxrVJkZ8ujdBHTqbjDyOzVY4Kp9X754og/6XSViw+d2j0
FGqqXzc8FImqehqqxF4fXAP6NS11/tLRHzmeqq+8uy8Ob9AXRLUyfyDKO8It
C8iJbFo4PSSq2MZw+Rses7WeJWlbykpMd2VY0BIKxLulQbPMzhjdgmjt5gJO
UzbVmrFzo2z7CpNBGritmmVjWgTapsZPd14rt4bUFonezS1Ot3J5vlDDZ7Jo
a2LY8Nbcb1c84NpxDRcnWzuHdnA8BkQYNuSpjDNHKGQrhs2fAYw/N0H9KDwS
EF70aVqtFag9PJwkcdKz8F2mSvC1djO1R1HjmDxbCkcy2ik6NgCPRjYc1dPx
Nbk9iAQ/snEs27xmVhTGA6b7n674M8X1ACvPtJpESdh50dkaTh2p+HSlSoeo
P5cqtec+aTnV5UbHIGlOcTgqeQWSZSC5qG3ij13ijZsjiL0BazrtzveseryO
qB1KP2t0ZI/ckDuO5+0F9gMZB6nrcv906yfL4ZCpxXld+/5aJG86n5Gnu+pK
e0XzV7hrOt6vXIYRtt87KZ/BI8my8eULJ0eXVstHt5cD/sAp7HygnlMutRbm
/x+evtGx5TlrBGjmcJJtD8lBcVmI5ujQUiI8CpEOtZSouZEXO2hYK99eNjmU
6HT3GtAhhy10XPFRyyYhQ0HKyuFTli86QUauwhUrFYUsE5s3Q5LB5wc32gZ9
/S4NYDHO0LFHopVbkHCIatNaC9gDhd+/RBOZMptIRbqzVajGMnSRWg0BTDAk
YKLPEqLbitdoD27ljBzgUqWil/fTIcX3aYVOPRerdCbefWi7Bh9CTFMYS7kl
cWQzUPpq7lDX0FeJqINeNMJjzm5ZmFpd3FvOLhc/V0CgokxjhbcO73fIN8tB
Tmxx0yewumQ8kUfPZgDoZgKgeYGHOt6LLxpUtuNBj4g+YkZE+Rna9gs3lmeE
oPa0GYjiGtLgVs7CVF1fFpA6CeXE0s1/5WKrMYDwLqY66vnk9C3Y+hrFRO58
WeHWBzgd3yeESE36UBdhRhsliuALtoE3l0+fMb7MeiVNF7RUnD1VnN+aPcL9
4SfV4UAFmVwBPygddAhTUwsfGqP8/pXzofQf8hc/2p8IFzeMugeoY90DdwxJ
mbcayAKWAsYd5easjGVNvsPoB33XCcL7U5N4/0laOoTL8JyBKVFc7aUVKHfc
OS4pURGdi83iGxDDz+nPcnJyKuzQHhvgdK+vGQ6HI55PiSVdbnP22XHleRBn
l5QPeEJFxTcaqwK3UIWq9lRwyLrmpomABaduwzdpJiqkMIfPu43daqdP/QhJ
dzSTgMWhtp46YB3rC+j0OhgXF/njJn8sjsQMvTLUY04mhXJoq3LmU/K93lxd
RnQD9lgpchJIQPX5TYb+pIJE0tO5vnLc2N00v3jBbXZP1vxcw1HXQRVCRj7e
biRcDWtPKlVNgfq5is2QhSxfeEmikINbOHzxjwhSz22WW0g2fmxupTAyTtiL
1Fp2Cike21vg0ZUDvGOri/hXutDjEHJVYq1JOXxePXDZQvuh6goPD0aDRWnQ
uwtQRB721/RHUxMVJyvlBO1yaZ/zxMumu5TdAqcgpU27xuespLJfIB0uoJ0m
FVbYhNPJXEK0G/70xIFVrj+ojreZsJ/uQfboOTIGYiaOquo2co49TBeGTe8o
c8+HAAAJRYwCt4L6T1pxMMRiorrUHVLybfaAXM1VOV48tZRKR3DOIlwG6riA
KxdpsMfgpP50ckqP9S+rwq+heUqYlH9xhznuWgDbQkYYuoqKFLSdt2JOF019
C5JvQrytXVdLUsf2NsZHD6XMBGaIDgeTnI7DAHNfodmPNC12t8Oun+yGD6zN
g9R9HRyUqI3IJI5Vqp0pSdp50tqfB7Fmk2/Goz68yaOfTxOSbQjA/glLWF3E
MwnS27DBzeqK9aQp6+S1rKF5Kw7iG00vJnWX0zqSlcA1dz6XyHa6YxMwGg4g
3Il5D3wJL027sO0PsEgsjqoIXHAkF7NURptTLP2UlEnjYZcuhh4aeI+Fv1S+
GeicZP+fIDuY3c7ny58GE5RCcyr4wFT8YwYTDxxeroTE+1N+8GEBq/d8SQMG
HjdiMdClgyDN4Ntcf7iCjXV6zLijZuo444PLZUnzE1WLZFFSce9CtnTw5fx/
qpPjYr9/rXCrGKBqBcfKtt3F8xI318/yMiQm8WdZ03vHGwFah82wNfpYZhrQ
vbwDezcuJCxInyNeIjbwkzz1QDtSMVhBWoImWN95t8sje9S9Rzugrl+8bP/y
C4S9vtd16QWD4PGKmfdqcFljjF1V4qBKwoIA9tzqAzZbJ5PYL094IpRXqP5Q
/ZTWOPmqbpVAz5Y+5BAKfnHlpHNyLtsyXgUPlGk6ltVx1iJyqFFMVPwB3cUn
OHhfRakT76QysMbgacXPlujF0kpWicmXikhyc3bXpiIFLyRXN3bmUaK1aWcU
f0s9QV1bMi8JrGM1iTL+Um3b3nlkGsnr7ntD2OgXn7KY44MFkrgiLVVC69vj
KOQRxAgb3o/19rQ0LfLw+eLWvgpnTCC6wetH5ibIF9v5bnUaY7jcHITaPviU
u1BguR70MhqcjazMl2qRDYExUkrNSsTIP8IkvCWjSuJXwcBAyLwAVil3AkIb
zjGIPjXntdrG6TiUmr+ZciSDHIHV+f8B+7c3nCouZksxCaDeHWP6hVqdukNP
jb1nD1Z5va+/1/OXTyrwp1h0oW95sE7tjVquqUFMvS7mQftSG3wj1pQ0umA8
1Q0KYaWa4fs6Bz4KndKLNafdw8sazmmdbg6n+gKg6qkw63MQ0I9Q7Kg8m6+M
ltArIoloEM/94kzjPqKZqr2Q6Y+ZGU3HNGrsBf5KtlOq8e4olnGpxTEZGQZv
snnsp71L7vTFrI+DEUNIoW6UEUI/BwQ9Pf+Nro+SsO/ip3gx6dc+wRf/EqtQ
OW1sWu+I8T5MNJxweojgIGxajNmT3rQfDV3PsuPEN0yxB1F1OQdWcbEDpiBL
ecWCvlmUNHvCvvZ35wOxzJxY7Ukjzoq8UB78gKzSy6myY8npHdsxIfbt17zX
wP8lsKWSFK+yYG5aS1VQuL9Cggzm9h0ikLNmT8nKhPTFXfHwnDCSg3Q0QGE/
9VaNzzmFIlcxNg991HkJj7p858OQ5lxQKyqoPVm3lkfv+kfN2p3kQeIC2OU+
KyV5zeHXXwhAhJaCZfkqg3Gww9B6LKU7ePyH+vhR6KP9JuFcA1ETNlUb/OBi
U6hjDP3V4xt/yLtTpJuLaFZ+Mcv8hBpcJcAaGklDCMYLAaM+8e7uGzmLh7KS
6Ek6hUgABxVVqQgJqnc8kW/dEPJmQkQjaNamzZc+qDNPWObD/uJwd2dCuD4d
K0L9gnpRWpaKVdY9BFkb07k4UOkFDWJHDWEPmKKyrU8BMtIHpJ3nQJ2lLCSq
yDtUFq/rZNjg/EX2mbZpwlvLgoCw6BKRCd1ZVL49261TT0/ya0ceZghLi6JJ
hRl3mdWhKJy8Lh3pDs1Xp9wfSM7qXgpSa/RxCgFF+1TMNgV77p0zhkyyWMtW
ZsCof+jgZGlYSSFvlOeBrbpGDRS/5gEdj4x+DzMPN9hrREsjQ2XxRTuzKwPl
wzj4Mazw4H53wEu0DzfAZdnVpqySTtaX4fbGLTBZKcqv1cwZDRuMTOONxlZW
N6YdkFVPFnPu91jjCFqEHlbcvgfjtZ/wjGRIRkU6QwIq+GZ/x4L3SeSc35YJ
3DXzs5B0CRAuvMtWhBUha7+uoV3mLa4EwDHrd+cpULMVyx174/hyxbPK1KWu
rMxtBzl5sicT3x6S/6F2bBaKj7Q8ColC5VuOPnEa3gwgz9rGJgT2mvx0ua4p
pGXPtviYuYs0+ivduywKqxW7qf/mTNzLHKQ17lcGTL86Fp//4Wtj7CKs7t58
vh1q0ih/ikWuP7TmSPth1Vgy4L12fbW/+eVg+25iGf38zuJsWJmShGxhlO9a
8ASfH76MnNUUXSsyxkpNP9FYNF7XgwUjeVOtPEbOkNQuaw0j2Rsfxg3lSFvR
2qhIovz/l7piowZ30BoUQsS1DoEqqZmUZaVZuCzrNiWTq4EnS9+lq+hz7Am/
tGYNjycRlOrGGt5aMTQP6w0/85xzJDnGiVbpd+IDk1lcwtZIF5CTAIKiJJaB
VukDZFjMSKD5M4+m2HqADdgm+jtN9289Rxuxr/a+VZPSFmK6LtXnJLIb07A4
w6eEvl7aCi9vfz9wM6JIZu736crh/jO50sCVGpUfeqZzzSirK6aqzSDfo6Ru
9GIFNBgWTxwP/ZFQWrzOVLBlKqNN/GKE2TIitHiTdGhr27X6qeLfPPBdpaKx
ekgYEsm2jWpN/xoV12FiEm3zUkW1DnKnBSPP9StsuVocHoSpNvnDZBUYC7vr
tA3Ukh2BMztUvM9d2xQV/Wg5jx/RiGPAorah7gZCZWYJGDRr7Yhd9vQlXFv3
FksdcT+eYCnQY6m5ARB8sLnEATNOTllBtr/qwBaHwMV+gpDkwdBao5IzxzoZ
Ue4xFx23j02KITFyTaAJM3+6hsT5X35pzw7wE+v636QSUz6850MCXJ4YCpcm
CBypyMkaPULmJ+t1QFDFVPN4R96h46UEdbX3fSYMIRtMy6ma+SNFvJFZ80p3
e3bredBjj+BFCeTMKwjtMCy43Kfu0UvGsY/jP6QzXHUJfezCAx0jc6hX+8/S
3Bawj67ZdxXPt3saXw+REII9RE8Md2Yrn2owXkyS7qFyxtahJPp0YokFcMfe
tBBbxf+a4jDD1xwIKe0APmn4ju8ngiBUpoITIM3HBpPKPjw4lpxy7+/Adcsr
zc22P7+1yVyA9WyxalSIoHHU2kRozZKuGla4cE/Ri8+YukbOBxbyILKN2htm
744qVwInzzocjf26aY9lSpL3E/xz6zX9reQ5ej9kHGtd3+c8cJZGbEal7kx2
AvqrZ8sixJckPasJggjbnXUrHiD4if/gjz4dM0SWO1iL1w5zIHTyk3B5tnW0
yoU9bDqAoc8EoOYckft5LwAVHf5X3ojGfhylkuHORWZ3Ls9zHFychy2YQRxL
oiF4p24l96+c2tOz+N4osygr1z+xiRcKDUGBuJlmaeltUZLWOTfjUtpXFpm8
yomVCtWi+n4mA4Xo8/CWCv8Mv+zdNBKrWHXuw+52op+ZpthkVnrH/b4iEJO/
ICGHEQi0zUH54UEBfwC0tQ1TwBT7a8EPOHwbA7Ho6Aolh2j6qnmgnYz2NuqS
Sm001n6OzhneFoXwCtPif/vS0WgF6YfidM8VjR3yy7c1Mu9B5Ud0NNr8+neY
Mfr/N0pE3e5nrfBuNkYxVu66oduCwhNIxMB6VEiyoxGTXFvvoPKBRwsALP3G
+kZk9Dt5goGJEDuseLYxEYD6Bw2jCkmg8oPHv2SMGgBasRzDoqrvYtvdKZac
1g96FiSOlUiKTtysZezEdNLLd6pWBWqyajk1T2KXu6Z/g7lD8K9+l5PQiUcE
vmapWA4uuwrpRBNiCvwj9PgIBSqPf1B4Rz+JgCl04oyBf2cgaKivIzgnCmDV
VuqmjaADiQTdRyzhR4AT+u79s2fLizSAiNxWApsnbYtUN1X9l784c1vcjyf5
N/BdQKAE70ThAulqiXDQZPRcxzg6KRRvTBd0o64BPKWzigmB4PIgZNhZfc6b
M+ff7YSCFZW6EVGTSI4RETrOQjX/QnMDdzPRDGSmF1RvBYW4xHk1SAlHLD19
eAZXzzxp6qd0N3ym3Ae4QG45rY0x6QWyVqVRgmyMRz/89MpXJH8O4qjvsnc6
ASADbZ5iww8KSJRZnr7V5gdWZgtOns8PeajPYM5VyJUC+m9MLlo9A/SOXLb8
Wgr+h0bx7ZUBdMwds50ICioM1X2aHGYwCUEFoVCt0y8UB9M9q4OdT/pI1yE2
izEq1XYmeKLzxwGOx6Vnc1vftUybEVbNDurbFBKiPkygNXj/P8xwoO0DPVRF
0QUE1Ujm7G5ao+ZuGYzyJyNDdmkbhJfUkO8jboYfNVbymope64vE052AOYlM
e1m/MwaDKkYCZ8qlA1OtiQYKo/8Zi130TdUrrNerXiFMoL592k/+UPaOuA20
juttZX+BZfhN0JiEHlUb7hmN2m2oen2kI/QCbiqndTgzBijuia8y5ykg0L2N
ODJyCG4xbY3Zxq2NIUQYhDog+rIuuuii02gZDHQotp2+P3p9kUedv4bMoEsN
NwMBMc2BJmkoMx8nYVimCnXLDNDxGTOoGEHZaMW3qagt7mh34PBaLJ80DbA5
+a+s8fE0HwSdbsaXucTxKVImpHgxOIRJ3tHcdaMr/wVvi0iQINfuLW7lEub2
RoXdzemGDsnxbL0etpKliUoyOekNH2l0u6G2OG53a6YnDEufwwMe1lh1uY7M
q4K2MDKcTAJoBV4RYfHjbWT7HytxirXbutqerlX0qk0zHUr7SJnIC/hESKud
/6lleOFsG9JcWGcPFxZjt7ZlAFNjw+eLs5o4+KMbFsy8akQoj/nnL5lxDUzO
oAr1KBpmr5BfW28qCDhaE85KFYKP8MP9DzraNXOR4MO5c8ZZeH0HOchv3GfI
FpcP0tbCtRvhfY/PR9UzKcc8tsLhkBx9B9jG3Wn1g3PgfWUB9gKtNcoIkngT
MUbKIC7SOnCvjG/oDTvQraJg0wyJ/DmERM9KUZGducLTIj5C1LyyeuUC3t8/
ntrVEhHXjbSLqYEPfKxZ7T90eScFf7oOgAYPAzboL+Xs/cObWkuYx9708cdo
c28UV10bVnXy9Crf1cSrXD8+yj5pYrHrkZhA3lJuvX297B1sUzN7dkvqv1mt
ql8X+p8j19S1zN27JUMc2kZmeD5grxySVlnTafGz2M6np3Quk8SX2pvo8n7g
jtHRcfciWGKJWf1rapBSROejtJl7/yDOT/O9qg8+zxH7U0z/O+r7yhNzLdxE
q/S3EKFwk37T4ODx5wHAlolxxgzoUQgrHHo1y9cxl0N2UxSX0vySGPYK6voK
kt5RGLMUaW8+7ifloX2otJVmgoe8La5OYMtvwO2YAv47VMA/sd3mSVFEzKLJ
pCSaZcCh8iXg24sincMOv6wNF3Aicb7tkLjmnBl6y3Yu2jaAKdQ/gIYfmUO+
MEtb4lXvenfjjq+7SyYVaItHeIkDH7Exs0pLTmaT6Er6gCgrrStU7vUrUwn0
WSjbH9sq6Zt4zMG0LGZ8t9P/ZFc+ASCzzUOVXYpcvu4U+ga4jifkHDOE8MGk
WD5jJFZ58/x6BeuoV+Pb+zAtq2dUBWQBFLDs/dudcBmUV+NhKTZ+vzmmWEKp
omCpKx0d5vw2cGTlTRP3sXicrBtZfYUHXqouh3H1HiPENkheL//8MDvo5Kfz
ApiPK8tzuvURMzXS4dgk9NyjkXq83VXDr88VI8BLsKDNDuFSmbrwfXcekaoJ
rgS+PR0soGaNdvOvHI6Y5sX43kHduk9zUAdITsuleI1rJ9uTeqUlAx6G0hKn
PO4A+EZp0EwU5efw8wCLXbbGAbvfVn0ppK+7p0nGFR7RkHq89lUbXHmuJHqf
3ss1CNrFJAzVvOJ6/bvOGjuatxy6EqEjKdwlLrbSut+Qb/w+3ML3m2036D9C
BE99BwEPeQus4Gb+I0Sj0B0k55AXeJRFGg0T3WYIqB5MtgiZk4q7TXSvkfHr
jsgOibSqImyQKKVCpTuy8W6nHxFhNtX5k5o6yzmDYmLIKBaJePJTgeCXh5T3
GSShLheWgoN/2NSHYkxW5MO/Qj7vsym4e5NO3e2gJ5KnLQ5YJ9MOuHlR6p0b
kb9NbJ2EDyMxkiHuPjyV02Th17o+1Yv3vyT9bHkqdC3zmFsWkpgedMBH2YOk
6BDozG454uHGyt57z7kGqb/UtoE8i6Z9lfthG2UnWtdiPr7raCqO2afIEYNc
+n8um19816zImyOxNLshC3DbXYMpFEkHvUMfWpadCYutjKb7Laafrtwq1Idx
VvW6WYVXTCARqn6oxlcjCa/uk/1tdSjmYxGa981T+62qv6zsyIVBeCzIbHWg
ez8/jXLx38qU19PIe2l0fNwt1HmMOgtL3lOsAiPClkZHr/Y/quNlQsuLjECu
xUnyDE3BSFXq+Snf6g9+PYI6i4Uus/Qlu277XNvBrSi+rXZ5uaVthg2qishW
wJOvEpTqz3ibQ56R7WtgigRad0vEnJMXOs2uDDjHlT9UWsHSzHi7Hr9GoNMM
TRS3bXJSGow/Yps0KaJHLYe9SdfwUQist8sL49X+ETgEk5oHGbYTOYQTr3ur
t7AwvfZiVedzNKmMjG2e6stnDeG5S582VBYfmBEvU96rUe+guR+DBpI8sNF6
B317EYoyfmnj9Y3dp1DmHWcRQZoIIQgBl5tlJuIeX+rV5arW4l4W/1QpUIpr
IGj+UoRX1S94cDb+88A4C+f41sYgW9KjtSOzL5hiI0DJIsXt2r74YvTjUUjC
FBnVCqJ+5QfR3zpfELWk1RcRgjh42RFxw930o8TGpdTfPtNe2AEWI/Gj8o+i
c4m/U8jxPdEvNe4lLb2+Xi01+WlolewQFZDKszomkIxDTYdgr7+zNZDSD8BP
b1DBX09E++fgqbR863FYZ2o8IcnHjy2Q3Q4sg3lrpA3UFO+s9YbgBVvkMXfT
xgFupMn7iwO0uvaFETBvWeCJkQwP5D5rvJDXwVUVFefNSAYeFkF8GEymy74l
igpJfcqXhYYoEySO45giI6t+Fsso2n4VcsUtMyF5WQEkWIQgGwFZ7WvnSj3A
ddx0BR6ms/st1ICX7+8py2zkaaqTJ5dPiRZArQZqAC8iyF7MiQb/8JTb78/n
M4nbzkkPHndgND0ywYiTgzHWCkGAA5W4fX9uDFEL/LkCj1YERZrgNi2sWlX0
ADRJ3vn+h+kYvgONBZFqpoPTgQTKvFXyF2t6zw+QepW5QCCifVyZHdO3mej2
4O0uaktUSTtkAwliqqJnBfYS1Ys+Q70dbwfhdqQKtfFM/17BnNd78/KgEwVi
S1kMo1uHA50xDeTxUMa5voxcL2ODFRwhzxWubPdBmu95lZkh5VCQhRSwl4nq
u2l5qsYtrQJBiUFGryHY59wlCvizAMqPuNeuY5Oic4I0fQfT93m78IiqzBC6
6KeVsr+ekhu2pXTmT9hjxdMLjk1T1j45NJ+qIHTojvHcvSP2H1My3v8u2tXU
AbgDWIGBVogK1eLOc57gQzQaysPJGMqnxlVl2KLWjjLkKkMG0xWrWr/xlY4m
xwKNIX3zgUa6s8xjuZEyFuWZXVfE1FQXhTGDxqFjNFUU0+GRtSi1tYFchLnc
S2ml4a4c82ETLu/xcvG6OPSByEsPyl/zTyaEXsKT3pIervKc18mT3vhLzAL3
+X6FIDBzTvToso+rQ3yhR/vCQLIpnu/XDfBOFzj/JxMxY//Q4dgArQUQz+wW
fjZ7FHgB2E7yIdlhFGDISEVKuxIh3S7N9v1HzKWNluQHwbyniVRiDChzrGck
+9hTpfe29wjuLdp1QJj19SFA8BnzYrLf5MXiypkmiM6tffyoveReZ+1fAgNv
QdKVa4XdtZTHr0J6cOJnSFy155cac36joACV0hGRHWUdEUnnYDNUg2Vd+bqW
OaUVPd0roHtjKmGq8W0kNLAE7Q8rlgWDH8mcET1EUGuBx7MGAYktq9QBW88F
nPrNFqRXVeM9KcnEWDsVz0QbtF8kcMyPMCHOQFmm4H03NTmpWM6AnS6fYCol
w534B93UpPENU/FhsoGK/xhKxPE+WHEmB0eb2WGQkC7gdloQ+3JyT3Y1fzsY
MCR9FSWELPHSub+xw6oS1+85HRR9MNu4B0TU8dXgadEBHUqCQ+b0xOefuPEs
e8Mu7z6OVffKpclSIPXks9Lm59LePW+5sj7iFYb89kWcEUIYTX4wUMrDpCR/
IoXxJH1ZKLNCmukX90w/NgWHkCmZU+0xP1ZInQoDBkD9icuZvZiZrP6zT2vt
JOHxGWUlgBnVXKiT0zL1Sq59AwXbD2joeYFZ3l40OCISegFXBVtZBobrVGci
aQfWATK7IVA0OZAUuHY5S4lwHWNU9cCY2FAeMHhcVNPWn6TZsUCujxA99zf9
3IKcZCmpt45Itdskig9/f21HMTKi8abpwHOF7zAiXG7DZ8cUhhchRvxFwF3a
WgrhUY98PbYUEmqSv+e0jg/4CVpXHbSA6Jc/h1UHS51iNI9PiqoAdr10g0vx
+KhieyskRb5k455Qdp6H54pmGiDnFEOKMCct5i894ga5SwXUkhfhr7ntUsIC
64Uc0mddw0x2FnsNImbYQLOpPNGPNhmBBL54pjjbJsCV9KTkNwWP0lckzDgy
1pOu7gGUQPrdIiRm7DVUKOAIzF3Zjwnx+YHRlVrAUaLEtYfSMQdwFTBdYDUo
oVQgE8KO+2Tm1clc5sbpQz9EZ9RdJOAPhHUBro5GFaN1cTb5MTkLRbiIVFue
bsbn8mV5ZP9BSw9LHmlfa4IJBTGfsvwO3iemoDKJ8jICX3ieZUnB4MnOnZae
msnxf3Sc4SYduazuhXrbUXADs5YBe5mfBpl3DY1RoqxHS+9UuWfrQXHAvhMV
qUNyP6S4apvkAp1RxODyOd8dXDR99k1mz2+LQKAx0YC9Y9EmxsAzMFsuQr8S
+60ioCC0PKQzuKrln4N4WhMDqX4a3luHN29DrvSobYlXoJOXdYBPDU8qe9G0
wtGZ6H7VjwOHbUJ8h4y7eVNYWrfjirO4+Xxa1Y0UNgywJNuXqvjZqxDB9LUQ
nun8P3J/IEVb1ODcRzoetZI+mxlYu7z9xY0fR9fD6xm0r6vSFaAoM0TjYqcw
iKFas/vMOiX7uROJPVB+Nik1OOteIYHiyOzsp/cProdNo12ZK+msp7/f8+cz
CBUM6ecj5bfqoCq/7HA9Hvo+lIWtWf7BvdSeLPjjn872X/zT9huD3Yc3vvb5
d8ODehiUvNaesvonQg7ENN8JODMiDZw9hJro0S8zegqQqv0UfSz2EZLE/Hjb
p1DIJy/MbQo0QuDVYsA8Ea7VeHe+VPSNGdBtWtYzjM358ez+sw29Zp3nSc+T
b8qE6OJUUhKktlNh0cvcrBKl9ftOSfZt9oN+eP73ynKLQAtJvDhpm8HKg1Ob
lj061L+0YMVTu9S/okQLAWQu5qq8Z4X84Rq7icfE02LCdlUZoezrP6H14R/Q
HJWHD+xqxUZ9dWOZbw1BSIHryUGuTG0ZQETdePCM+N41VnS1SMYHMQ7BknYS
FkEh4YWhCMatqCvTPpZAX0ZHoyVoIZGlv50Qd5W0PT+AjnNk963NDkq7p3NM
GwvVfzjTA4izmTqAJg7gj2254Xkteyw4SX/ZXJ2kcRTnp9Nci8EeIZzVDD1Q
C9Rq1wIc0KY2FWOyfcJt7rjJtaxFLKjt8xVwHnWARA3Pfdz9swiflkppAgwe
i3YTrw++T8yX4IwWGiHWhQPmeI51O72W3TnDJY2KXbGNL/cPrVF9cZpHv3yN
qbH0EOJ2uSb5rw45uEJ/lKMKARGpRS9caZyYWk+vLqTNsz+ABzwLDJY2L4jJ
MJiwUOxug0BUUQpM9ZOMkCwft6c3NXChouUcsET4yrCGdOCgmsTactKaQRvA
50iWTXd+6ezqJgp1trA1h2Y/3CD29WtQ5SJeyeSpeLUS4Gqbmuc+RkRf+oxF
MNDtOb0D/m1Yq128T3iojBMbkjhDNYb2VU7byOb7SKOOCZypHGwkFZJV/g6w
JEBfrxBKrWGjcvNgZ+30TztsgNJnbilcks2gEfjU8s86O8WRYAubphasp3VG
aEZq56qWSA9joHNCBqT6oqkAFHlkJAG+FjeGaySWY5bRH1fHiSIeot/cSdtY
lbSbROG6E2aF8CBvL8C3d3FA5bIQ4vVoNO9PD/ielV31PWabGibRbj0O8PUl
0E8Bd4IP25ZRLTy1iqIcTdZ8YBvL6FjBRitlpHtnfPiGiIn+KB6ofeqYvjyJ
eE9DIXhCiwecL4hvpGin8q3dd96cgRfngroqKgeRR5/E9rK2M42JJrhE6dTZ
4fRp70YXHQvUlYipbddMvEml28kkqsOvRHMR+RwBqIYUGwogm24UX4s0FYR+
RxdS5cvzkAVKqomkXp2ykY9gJGu+k0CR6TD5TS/+rFltTIiQpnvXwByyF5TU
nKJONDWTPY6cbW7cOZToQcCAXeTAf9qNqWTLWa4ke3yEQsZ/3Jg2iw4gAo2F
/5ZN+dakYSGZQtFTf8Ej7+UwwMXVUiS33I006oCjBCq7Miyns0iAB8UgfRyB
tKl+g9llzCP8kdTTXlcBtwFloe1g6dPwyTa/62tTmOg1nge0xla4Kcce5G96
/CevVMtPPhgqhJZtUQ1nPhfFgwPcTSQbj7vZp3V3YJkc1+kA6pOr7nCoBzcR
3hhZ9naRBugCaBw53n5VtTJ2Q8SikOVqNULAKSDUKD6V2RCrKqKqADDw3StQ
MCJuolmR26oURMbr9Cx9csJlpckllOjHqu4KkLtQtahSpxE3uPAzOpRoUCeu
ZJJMhAw9/nb0clAuki7HYYNAm4MvI9/RGVxiulxvO9qRrLUR4A5h6Jt5+t//
JxuACQhXdWRYZZUqN2Jp9oSrIAaKBOD3AKzmzpG/BL4VECgvayU1w8kflmhc
3/BNmQIZpPmTS188exRPmA1a8OWZWYzE/DQC/K1ZrXpV6TeQipm030UN3Bvj
VWkuwU3EQUgq38vh9Z+0OybIlWBpkl3XBG4r6/fGn9vKh4d861Hiw9lPjFDc
TYK2gJTYhJmxVdwjfyMNaRhY3m+JiVPyA+Bj9w0v+jdKtsAs8tr3Wgd0j+tw
oFTTyWCQIiyomAZ0sEn8vNRr+1MqLVu6jlygKGS6Za/2ZczcDS4zYD0b3jZZ
qxA7Vahn7n+3dE+ipO3f2+ktYSG0WvsMvnVy5legrzcQ5PZgQKIzcQRMLcFS
mb1aJeRF/huUvz2tFS1apcfSoXv5MLVUuAjYC3Mg+NTUBsW1CjcWDkhuS7jA
3KfRhoeholX4AZ9azEoThw7+VSZCi0epkmFWZdnkseYxEwRyidqpSqBP/OQE
t+3WattodmoVESQAx1/VADn2EisG5EHdXESelPJS41WMJtnNmhRllPtjyJf/
A3ZIZ8LojAMju0gkOPM//IwKyUC9MHYMjcnIfraQE/inzA0cZjjLSnoijXtD
l/Er4z8xG4gVS+1qr2kpTDfy4JxuNEPO9mYwwSoge7FRoD7E92W0rr/DzuQN
6Q0vHdQgDukl9ekErWzIcJo6mxGbHL0QLU/KLz2y/t0JqHHM+fXgsDnEMB10
KHpcj0CF1pD3hccZJcTYI4DC7TTRB6hCuglSAkpcTSTfyMuegq1uDWAUnHmY
lMN7wqmRnJq4AiiCZczUzrajsH5kYSeA3bbtQzGGoo3NzjaZOjPOvtodQPEG
HuOVXRCDqRzcl0r+LHXHm+uT87sgjjCSeEEOsPoAmqW6BQ8F093Vefkn5UsQ
W06sGwq4n3/bVh9dVlqnlwwNRxO3r/y4yXHIok3sSg1vIroTk3K2Ehl460AS
IylipVQ3VeVjL8ycTCKV3qfeocf40qh5uVNkOrRlMw70M20Nv1QxV7UEBTo3
CuHwbjc4G8kXxDublOr44srQB9DTuJmYsdbSdqZ2mzWOcLhVYXMb3HVZ+Of/
jIEzje5PBjJhnrQbcJ2zprvlou0V+9b5uDggyklRiuIO2WTkwtKaJVBsUf2a
wGtgN/PTIrzmc/w6AYIdVn3+zyna7ttU39hOLLaKVGUYPeABbQ4rdtij8GtL
fLcCoyf4TS/GXpcsE7Id7T9dxj6ZTlNgvanoyaBPjjbir8a6vVht/Hhrt+sm
BgX1619IfUpYxKuR+2KxIYyni/4PI5es8dGL84LLbJl6YKP628mN9V3ca34M
eeXio6aw8J/8styBd04QwclJK34wLiv7cNx+t9DgspMwBUFJQk2ZUDbqXWku
w4nN1nj3x+NO/TmzevIL6yv8yeA7AciNMt3uHFiOi2cZc7+g6SSufwwI15se
q1RkhoCaMeEm7/uM5euS7wEv905N/RuR0O/w0GFGba3LuD+JimVBRlvZOy4/
fxr8gAodONERkYpuAAKNWdFvtf8IxNa1/zlQWsdainZ7AtYFfbi6TJSxF36o
XmDtTk7wvMeLPr4erpQTmbYLbzIW2y6iOrE1z97UA7vOFeOSZhyN9YjAuAax
kKlB/s+wIFyI8DrkywRD6CD/52i1x4qHEtI42imqh/VvGI1NOoOxLNZ9jS/+
O0Tstg3OLcSVkkveW9WWm+0okhYv7SZuk2cD/jPPDV7CsclxsZ0fDATRN+np
NNfZVm8B93suA/94hq5StaeOoJi+TCFY9EODx2b243+J7dJyqvRC0VThplo4
XvJhr+TwPFETk+x5pvdRYt00io6bLwYZd1GU5HwFH3+Bp68PO4z5sHSX92W5
XxtVyaG45yBSDEYB35hQrHPQgWEpQ2jQuz0V58HIGhzG0G3SjKVd/N4rcm4B
OL4wkPJQvG3eKvt1BAK6+6J14uy5HeB2KVRppMT9Kxaf+FTKIRm3eHEbEC3q
mROLNIttCzQsum4tnchoYnA3xpYpcB7f67uKD9UiIHChFKfsE2ysMIvmmQFd
5E1zXesrxLGxkRLXDTva87/BWsAks19Wpke4XbT55gpeNNNgSpmq7gtllxCw
uNK8/XIcm4GxjmVCH8Ss6xgpW9SQdlbI5j5U8+/wdrkZJNSIjbPiSnea6nyC
W5uca6D5BwEhREmiN8/NDGE/tYRjH9sl3zapRnLO74nw6wahz9HPnFO20XC1
uwj8r5Cm3kkybiBP7yEmbN/d72bwx1VfJ1Ui8NJdryJWMoW+3kbWFW8zEUA+
0zyrNjkchXQVWKmu9F18NNGTcs0OwA23P2568RBO9LuHv/o+YzMy7LPTgPtB
9q20JKSjDOL/k0kTD5pXqYtGLhoJ9fbvNgW5ZzLVDFN1sX7RfYAxfyoC0sM1
IBpliv9TLal0V2mrZ00YVHCHH7TLDSQcn8x5GLG7TduSumBbW9+XrCv7hJby
l3SNlu1hNw5I5Y0qzcCFOwC+fNyJpve/tYRp72ElIzAg1661Lx2rzTwh5dn3
gSZmjr6cpFfWBekiAqylz9Bp0Doos2Zo8EO38FKjmZjUbOa8rXAthbPFe5w6
D4RNZG5gU4jnshrrBRoCEG9ryX4sp0aUgCGQaTPeXE220lf1QO4CPIjLtrsV
Ywk3jjarfnHgSjM+COCYNS5QGHTzqw37QK+2Z4GO6jBmrllFEulRJocHVOhR
rGcoG9Yg3FUb1ldwzujWJss+QXQazAQYSmJ3PnEu2VNHI4FsjaKphZJZyby3
YRig6hDCTnThkuFWtMv5bzV++kknKq6R867E0+XBy7QmVwsXUkoaB+nrY0dE
FSAfXuvKqmMk9jUUrLRVdbv63sv6ni5yWdNeMmTsuLucFjFYeoum84NBCw4U
E7VsUClRbT43i8XWBvniGDD84kep0/ccP1kPktGBOVp4tR9Wnd9Cx5RSOHLS
OcTPSH6JBN2xNeDPtnT3SGbGcAhS4E/T6YnOSrMvK19ddiq8AmGPiN9DCFrc
/281pqR4OmtSIsJ2tYPOPDzNwt+rFuONBuFQnQjQyWqtdoc64aYRs//walHr
A/gUKmeamDHXkPhR6I+/nBnCxWMZk148f5NuAQu49Xboe0zI9gYKTXwcf0QD
WOENbCv3rfb+GzdnGNt6Tda2Jiu/iVqBmuhjD5JARgYTGIHFL2lXnri0M62M
1pLx7q9qq7v76vnHBODNos3kSYC2nPgQXHPDDcPExX2xr0OKhJ9XWciih26m
FwGwXUzU52EyglzW49pZTfRDiuK0TflBgDmGoa2PDpiwmSHeQzkM/c36F18r
DzDzktsPl1i3rY100UptUi+ckk+3iLu/7zdVB19w0L+69YSa8yg+g7wNCoML
/L9SyPKL2hMRHcRlfW7h5fnP5+xI6a1dGyyszza43vxbigDqwOAXxgqK5kWy
qbnLTAwxedxy+K1NtmoFVVzhRch9aAqyskY5qroM9BHEyVbpZEpW5GMmkMfk
prWE5QbOixX+Bdxv6og8heg+H94ul/QVDH/aCFCWtb4NGxUFj2h0E1Hjq7TI
BnWh4GF56GRZxPd6A6WPeXNf22Y+jBEs65HJ2c+K/TDUiuEcho0btOuT7Xet
NOt+ZFzkAYS9SmPiJ7hTGKeCnyLaUAR1IUXyMtIcfg6AI6x1DCJXPv5Z4cWd
CGWXg0saad3vzRJq73bb1TXPCiW3v3P03DG33jWLZ0/sqZz7KRvnHe//gbqA
iQiLSJkcR4qX+GkjZP6zl+Y1dXiKgk8uzAU5Ght7nKAps8h9p5qj24GvPfGx
eZX9ZH+WZGPRy0dywOexk2aIll3M3it4Q7SAIeYcC20Yn4hd/V04UaTxrPZJ
ENT4JvkrokkkyIzpoNj/nBXUGdi7UbgI/i6FCeShTbEyhaATMTH59Xx+ocBk
lzjWpnIp2ZH5kVOotZCVIapFkzu3yJAnZAM4hAcB82ybs5FSeERRAaS4Ewp6
NwowwxFgV/208MAkCYw+uRk6vgRmJrRycXz8DQBRvyeM/x68TcoS20cSaX7O
pxK6BdarZmclXyKSslsEsdLFRsrFSen76M/qYl6UzFN1oWZFz4yZsbOAklJF
Fy97kfyMNehtId9chgxH9LgnAryfqr/V1OFQwiu4NowmbSNEJkvNrv8y0VwQ
Q0ESQsljSdzqxtWjgZ+lER4c+iqz5bue2qkkyfGqP8cjbpDztSxKpZjD7bbg
anmbkSo8WS7mXVdRv8ybB1v/7KO/U4fRiVh+pDhG+gOce0LrxfoVa9wxulm2
Okr9t1q8TO5jAOpGf27HmaHINXGXPAs0geHaNWfKU5a/tTNoyLOsKx0ptM06
jMlpvfPFYEIU1J3oDDpb36QSO7Ks3SO0ZexoCqY4B4GtfWKOFAP7TggxQaQj
/m/B3PoIToTpWHx3HyVyfSQe1PdDHK7GwxD+4wKWyqNZ97rcS1bZEq4bX7dQ
vOzpUeim8Lk/iyQpmjFkNU5JNu+/VDviV8qOeO69smwJbrv4ynG4KjJIXI3K
wr2yqERaDVOMazIvRsxcq4Agy8A8bWf5plonFor7DOugtY3uUtKmzo7bzPts
iPa5CRmYan5aE40qWZ88t430LMTEQVfK0PGk4EsLgs53ErjT7gTbLx4uJF4t
OfadgCn/sLP5MbLT8iSkby5lZ4pA8LZaXu934tTYuGfZuzHGjNwZrnxxOOOm
3/bL9Akhi52Nzosf7OiMbLX/aS6lf2Py2zwZ2I8XmWtQDbX2SWTQqVW/jZRd
TfIbCZAkPemdxYxRVHdKcgJmJgSGipJOCgxNRBsx8E7uon7CdKhM6t9zlTB6
VMYBCMsnL7OQbjvxDz+/1uDAJr5oWmLTjPqWUeTik6uARfuM0piNir5mI1kc
517Xqotx3YENFc9+cB1qwoS727MqD093xLLkuQf08pTDdm1yAQefsFgJ/WES
9twnOan4lFE+c0srz5u07TlHdQGJqL1PMyQa8V7MAmDGNVpUxNuTxCL3+GLG
eUbLa4nHr1haX3vQfWUZJCL1u8KrkwMz9qNYSyucFJweGKEvi7U6gbr2A9M4
XsWG0kY2xa4CC5X2Of4ofLyXlgCU4lVXTddN7y6DE9KBa14Bb6Jyub5NfVt+
nf9tOWbUSZcKSf745O34ASRvhAoDaZwacWu1EeEHpeFd5YqNPgC+6+cML+EF
b4l0+6H73z2VZi6zg/BQmXXsXGt6E1skRQ9Oy0fJxVi2AfkXUlPoT5/RIL8D
z3/XhZCRUtqhm53gR6plNSes5/3jkLujKbzLjprYFUCbze5KM7GVP9YcqSUZ
FDjpi7soarNmI7JNJhf8vrZs/4K61jVJC8rvkix6nkyJqn35hbGPmxeTxgIx
vd3xIGBHa9DgpbhDEqTUBdWbrArDbV6E0qE1cDsEYibK3/45gvtE0zpMjdcd
T2ExYVAYpFH+ULFQjYA0Lpf7OeLfrhwYAA+EJymX3wlsRz9s6ZmOqvcXyprc
dJw0+2fFKmgbLFj7E1QIM34/wz7900C6XQfLz6xlBe4sLuZl2D9SYPye5FWt
2qV09WM+f46hJeBLx/rR3F3l/h+tpUP4reV2luENXkDblsVZq3xR7Lfrt1DW
SAp4iYJW7ZNVBPhO59YHH/LUWiLXMsoFAEj3Ni6v6z5L4xbsw+plATrlKjQC
Glc/7GxKBrDHycYYhSgHtbrjbrCCSgi6tXUtar0qQc97GmRGRf/dJz9h1E9N
AwqqOaisLn6aAHcvG5jEnA8c6rLjJ81zZjL9W4kgRJxVTKrVtHCKuHasj/HO
juolbtl+D1lQdFV0FEandEvWS7loYPRX2e/+em+swhBU2xF20GFhdZp2U9ZK
sLyvKtqZ2rhirsuTshqjAuNKOQS9wS4UmXXF8eVuuWgtV+nv4Ww9yWxAMBFn
V21xmcQcOQr6aP7Za5po2bbR+lCEhEoH3Iizavkw0mz74C1VzWSX45h4r9GK
lCl3c+mq7Kf3CiD1xHKRO5MaY+RbEF17DqgEeUj8pdAAO2pBBx/bRT30XQOX
o9+80brRli21JoOr447izfWQycSPQgq6kfnORS9H7yaQCZRqWU8yIZLyAgQh
uQ0N+5mmRY7GXoLs+HLCnTHigGE9OFzfGruHSUXb4Yv0yV/P9Ly01PBeNKE7
5xBIgXFotfHMGNWic0Xta5CYRlWoolBuRgKbIro+GU2rIvwwlieaN5013atl
WsOdS9/jpIGsH8B8ygUjdetTQelZTUQcGrkZuZ+k+h0eK3tM7e7nLjVzyM+B
cleuissVVTLhSP6lpKoK+KWpOCGlBQtnyIyD8ThtF7eX3nx7vQOXRtQnJQlw
3ZR5vYM3WGN+3mc4C5Ol3oqybTKLZYz/GBE+/ss29b4EhpwHBp1Xjriq1zjG
g/JIsl0dks73szgwwbVDKcv8vXCPVF0X0dUhhqY9zL8W9Qqvqnz/BXzqcNIR
7TKH3P0u6ZCdukEtlm7OTELR0r0ZWo9GzRcc3cFLx/TMmkrgG9vKNTmLYoz2
c0oEpEXnpryMtBJ9JzCdfLKOmoCwMCPa/xkxgFjp6ajr4G8bK1fNHzRXQc5D
pDYWM7/WkqOO0QFGGoP3YuUUhMU3gRvmzPGM/CowTW02hz4RHkWIJ4dxpxLV
W9kT9vi+ecaQngW/K+BgibVPQlx/7HkzIgx3C64YFDvOdoko+Dfy8Efm38A6
dKfTXT52Wt29viJj7QbDcTBWRx5A7IWKUN1gqELkSEj++ric9lQd7hH+0DAn
uMtuGeUHhvw4r9UcXA0/Fat9x+CJi1pIPtqx/1IAWzT3B4015SoVwj7SUc6y
sKt17wK4CJETEH0tQ4QJHAQ6oB2HbtPLTXlf6O9XqghBSLNmoFhN/J1T1poL
xG7fhHxc8+BypwQJgA0SLn9tvCLXbGDb6S8ZcFRS/NUsgNhXmmSf9bh2ATTF
xwouvfMs0kbfhbxlj2/fuRIuSDicJH0XYrWmy+cmgfIpNP//BIliqn23jwR7
wkUOkLJXKGabRAnRZkW4VGpFQEvoihViIhC0f4y3rPIhsKOT7/+Hl7jkaDs4
kvH5WRVzXnEhFnyF8IhT09QQD36iBy2DeldxsOXLzI1UYNAubViMemie+xDe
tB9v2G0S8uOEkJ72Ol1/5V00wOnFi1hUPlDRFA7cC7J4Dr7YVb9pDnwWEUhW
pQAJSouOIQaXyOmLfhrrD8TApvyMX5U9d/oz14VYCQv6lFwij8t0WIYnQlUo
2N0FtiUL91T6tyMzidgCOp/YdjKkL9IG8L2N+8eNmDk5D1e943wmzWZT49ob
4L8T2FHMnIVWH8zDnl6xcG1+6D3TEakNX0EH7q3eh+Caj68RxuULpkyBCUHw
c1soxXZbLFttZUD+KmdFIU8fzlLNu0fLP+jAf5Rt6H5TdR+kxDjmxrZlUo3o
LPV6Xx6sOCQWQPy5zLehwNPGm6L1U8TB9ATYey3iR6rJfUqSKgG7hzYUz3b7
LkF4yjVEfBa3aMtqCt/12/UYDiYQmMXcOpHj5Irj4d/gTbm9Ecex5/E4u+YU
T8JUKuYiG6Ix78aRlidNq2WwEQ52XirhilEVXUK6RNTS1YnSKCoffsP6gjtQ
BSJPD+CaLt50oJFyo741uDiVt+Jl8cYma45O1BbjDOALshPLTpB58RXPhQyC
TX45hncHBlFPSPhmLQ7SQxgxLGpgHmvQG+thmHgUX2cXy1TzXQ8hQyCUrPY+
zpsh1abtpg09qeb4D9WZA3eoS/Dy9ZALmpKnZI5hybXrBmJAVHCZI5f7UPOH
+rdUznOe7j9Zw0qLVvXOcDdqXEi/m4qoU25zmPqP4eZM5bI7be32ynNjpBWS
FUcGxVRNWT8r2e8g7Yrma2FJ7sYSWVTh7WSt3knoIOGC0bFheiJqsUrZQtSA
xcysDpUXZtYasVy/8UpLoB3FUaKO8Vr8E7vVU08xYUzEUo2NgSZtaja4fkLg
rzT3wvMircq+CV/+JD+wAd5frwXLZNd/ZG/ulsTfT91aO2Zl9lZNh0qZ/l/t
5jUhEZgOP7Zsm/XS7/dLndNiYOmMct+lllmG+dot9W5b7WmzuGBAk9Ju5Dmu
CeOJ7Cb1yz9Kx2BRnYsY5ay7fXRvUDP9ovtm/Y0F1iqd7LoJceNt5yIyX+0n
ZG03mC7aimPUkpS5BGPzOybhHILsVWitxS/3lm5a39agPOaJAo1idMaqIXER
lDW4psmNwZ0r5H6SgjR1S1Y1AZmyk6JAFBPM+4U4vhWjo8C4bkMeoGtfZsr3
s+SGEUCMGKYC7ywHhlr7RgMFJwhZrTjoxwoTutF0byVAaYAuY6BYI+QyZSNW
NS9o8Bu3hAFfTquFJGFerl4FskvCxf9LB/rTnCeBJNeKFTY+0D9jclI0Hhtp
NEHmNQw1gqZn+xq/269eglxO/yYaBQsrjYO6vP8g9Dy6O93T/3EDU6BhwqQB
FkuZ7NV2GoHPcLn9iFk7MKvHEagJfyMIFueCX2Fg+4eTczu1kWDaOzuqDSAK
8Q8cCborB8BNCMU4np3xnmIYRrsuvO44wM/pHaT4wVQ4V4YBSFMPV1dgdFjr
Ly0o2+jrmZxyjwcjztxQTfgUvebdHQKur9uA9H+5zK36YQf5TQPTpUBSgTac
PCN1Lp0dnKanuEx6faPPR/7IKtSRAKkJrPp6FrYPMrw7Yi4DV6vPX5UFTE7j
yvITlQMhOnZ6yji9lh6UxAD8Kr+TxxYALdHQxh8mfWgCzc25AkwNRPb77vRD
jWkpvhkX5SViu12JUlhIxa082BX7PqR3M7i2iXdmWSWBqdRzUJbw60YDM3gH
jn18idzVyHOwspK7RliBKfkIk9WqLmM/OYm2u74oWqV88bYFWCX7xshv1xxN
AoPp6NTnxN4/tH8wu1hjZZ2VM3mn0ezWitjloeljhBISoEmnZOhwni2sJVMT
GR4wh+9cwTW0Vlg943tW6nyjLhNAwfLSfYw5XCJ73Oe5Ctib0rAifqWEmQfR
IEDkUZRiFz0oPc1T1rj02sZzf6e0nH1PKrTJoJ2AFixZy4quWrsCSP5hQizw
gks4gzSfE8VjvV+VqN98a3FIQem3ThUoJdr8Wy0Ymr+bthpdjZjowg4o5qmd
BUR2IAxogUTORnToWFY904XGgKQkFteH23tp3QxVDgybzKudaS/5lxSmzv9k
y0kdZjGCiYq2+u1uwyEy/GaV6IQsJr7DtKXA+GvRrKNY+B6IOU1z3fKPk/Ai
eOIbyr86KlP7pBSLkfuEsu87Bn3NEIQddOnWVNw3RLVGTBFSQYajSPa34Qsw
0XYcaYyoN0UhNsSww2EM/h7daysdJIdVBbJTMeAssbzbdQxn0pwI8eTmePbW
GAP0C55fjDDN/dRkXNz0/MOfOMokdiW8S7ga7WEpvBMKjnVatDhDAKqG0/7r
sBTItiGofIGiGFXcf3GksUQhHm4dNwol6k81/z6jAHS2vyva4Hj/UShNsH+q
cmLI6t+2bz7C9peoKyFgEYC9i4iv03BZTsZ2Az+gla95Kt7ZkqKP8O8z3j+B
nuevEs5XWhSKlVnFPnQlKmTkheuYfftKqFi/r6tJDlLZk2i+RQcnsoIobFSF
FvTtbXjpmU6j6JB+Vnqbf3GuLT4XnD6NubOdRC461rdQC9Q1uxP/kSAublTE
rLYdZ4Y7FmyvtMFis08LAhnZMsmecg2OHep4SR6uD26XxGEQSNmCKgRNW85H
TZFoa9VUAiCVGGdB8Cx6/45zBP7K+qOloxnXb94uqnRRG4qO3IlIx7AWxT9I
5GbISD2/X/PyC62XzxnPz3I9BpAgTdP0oH8+cKy7dUNiTYxgZtChdfOS+6ZT
gUWhiFLii9E37dK3Go9xqMjCgMDvfU7PkToNzDyBdVSMxAXJSM+SeF37dhHn
9ZT1Bt9JzmOv+zitZ82tCWupfipaOLDpAVXYIk6O2x4vIybel7HVeHf5NsbY
1LvmWxXnCWIKQ5VUDv+8ykHxoX8WMcIGJ9bDQ359Wfei7Jehw7bHa0Yk9ch3
Srcmyv3lwEanHZ8NrjNRypP/Aw7K/Qk0iJZ+S3RvngSJOaTcEulxwRxxZmiQ
7wG3EWJjMVdgt6vBF/VFUFlndC+4tpRXOyrUoy1T9qcsPv4HVY8j37xZ56pq
xDZ9R+IJ8sxOS/gWoHW3lviRT3o6ycIvB2H9oNs+S8q8KK8gDbivQf/PNNkf
5dv2xxiqR/FlQITJLOlHYtflBgawe6wicaVut39GvecCNBEggeXkOUBzQh0w
xeZdKXjbKknag/kk/TAhuEO9SXuWrcK59YcpYrmP2SwD+wtaCROQgWm7MKkC
P5ucRspIXrX+93YrzCXgRgn9ozBDzt5YGyo0JeUYepsmxdOPQzqc19TpwQR6
kF4dn1soP99fMCZ8kKsodopxl4RAgGCfIJUrGmrqX1fP2mcl1sUGuVh0tCbF
Q6AO6NQktHAr7l7C1dLK4VcvklJHfkjnGzsC4C8ZfQHyHlRqO8YudE9aqPJc
dS3bDuc/PYKrthbZzl57j0gAnwHN8ojZKyHmwSzERTLtUKX5yvVQIbtBWS6x
5nYEWs95hwptpPgC5pbrUwuLJbPV4wfOhrpMCsXEMCHl42LAVCyZ0gdwS0bj
gEqSTcxZUK2x6flKME9M+75QTLigUgPBLFoGNSZfBsy60iT2phq20LH+s/4x
LJ8aEAEnqp14xOe3DENhfhnkV2Yx0KogIRyQvgFpyCfkce1hoh1zcBizL0yL
/wx2zuVttWK72IZoViCveNDNYyP85ubNO0ZShRZroAd6or7J2NugrNS1Q3Ru
m6Bdwf6YA5HOXlIxeqx4H1mZj+PpFOC0R0bzej5QHtuUsqB5E3NFTanlvb7B
czYFw16QbGaIvjYD2fF7GjuX8BCF7c8RdvCg1MyOkXoMZmUyyDgEbK0eGW6W
jPtWTzF7hXDLpI6nSaJCuyl6URPKmbErxWSUhsOMxWleO2xDOTWhI2I1qxJe
7rUDDFlMTmXgrse3htzDceDUpl/Xy3VJzgnV2ujepMbQTHnvvxi1Q/j8X/af
ahzZNSPgYofVcVJ5LgEswPgYiW1HTzCTPvvsJg67KxfgMHwqxuab23b/g17B
7Q7DK/dFlLM7D2C2STt9z9mj3MRaxNtj/frBU5D43alwcIRDjfjqmmvUbpyp
1PSSzRINu1M62gpsa/l0zgphfLwXmrHrJAoGUInwutSSAFdy4/+0i9/3gBGG
MQ3JcdP7+Sg4MiqxkqIkyLchlXAgRrPYnum4mBEHmHA1oGu4GLOXQVeqyQtW
yG5ONPzb6Cgct9LPAUIq94I/KODbJYmS4puFyZhILUDvpxqlxMdxdyjtZl3o
REFJTAaPbtLOWlNPp7m3SgMavfDL+dk1wIVbBsjWUGsPYl2sWcuTavmG5wJr
9QK0wD1ms2MgxEyfgJrlvBJwqd/ghRhiioShGWUwyd+X2ccRdzIbM8ZGisTP
nxYh1SsNg20flGp2HF46lpcSTa9Zg/09GSTuGxZpuK62dovTR/qptX2RrfwZ
aH2Sl8TtG3tFGA0nde0TtzBPSBIWhyDqoZDwKZNjRHl1uZ/TMkJq6lMamc4Z
4Inkc/HMw9JCWXGHZ8G66o1+7W67eL4AmSFny2OiBXx5J/jk/FgI/Ch7PRX/
68I6eE2KckZY4/i8xuGHuBolZEQIWx+0Ye5O6M3MlHuuA6O7Xyxiut/TpCdg
cVx18lHmmK5lQ9Tb4bO5SlFB33ofFh6LzgaYx5sUV4t2o1ODqA8sHuh1dVDj
hOfFcFk1VaSbsoiBrs9CZi+cB020XhZCFOF4X6ZoBmxQy6uKAeqaflrt+af7
sR1yqYOzWLxLnEaqWHLUEIlArnEQL6n7LufFYTcXL1eqVZOUZbPh0ZyzRvGU
hf1jJ/5t8Q5ykDt1sN14mC3N3/oWKwGB8LOdcWttf/jYuFDpWlP+Rodfw1xb
1qvX5Ok0Ge3qmMwpDSosgTH129DGAGwOJBfom719RHWL18nsSRPy+oqHtEfj
423cYy3OV3zp9uurwyzoM7NO21pKgXblSbVTgyX8Hr1qmCHXogR86xanKdwQ
22RFyW5hwgbvzYXmSzSTvtu/LkgqLXT87w+AdrWseZi2dytN5MrRd6ZECIq+
FL4PoAlLoRNfAtFSdEeVmvN8Bkf57g8BgRHNtXJKesBLxYqx4eOZK9lFI+rs
fyjCPwnLfnMdrmQKaFSG2a4cdcRI8yjhSSm128qs65Q4cxIHlJ6UpgU3bGfU
NCykIeuPDYbPqdPWvzSz9ZqhpmvJ0Izd2uKJhTUt4Y+wCp2C0MZ3xlRV4YPu
noIsApBjkBHrKscoJUO/y5HECRxDwjUpo+HHXQYaS8m1sSzbRS6NA22Fioct
3FjgL2rv9LSvvprsf0nTe3WBY8F/g/NAOoX8i/J5+614xmziLhauOLUh5dNx
4/6NwBgbxmT0CPYqLqnS6qhtpODPLIbbJGxDB5ucDJDey/KoGPA/msoAZGOu
BgFgONBQ61m6Ce70C2l+cmICuO88nwF1KoRRLtfcRtoU0U9/QnGPPcpWp5NB
Noefc6Q98H6eqTgRtjBr5ARQpaHbTf305+QQ6fpW6iRm0gX/GVJJUIe3l6+N
TJCWfZ9IXxPrd/KGDNOXbDRB7aWsEMBjb7azGZUn58jb3c85LqSMeLgulnju
DPrVB710Sp5uwiJaOnNjnBqzoN6uMRRBdTOAGMVxK29hYA9xHZbHUPHXOcf+
OiTWQYB2eXPKHgaSSLokBFVO+z7WTR97rXMaQXF590fcbwiRI6YLjhjDbEuy
sL3yeyN+xkAgrVTQXavmpfz8eiqwCB7hjEtQjW3nhv2by2hUN7hB4MdJxD+h
FaANiFsHPU8NztIbaPyPfhrAnbB77q329KlchPEidDcbs/kbW+htgKEYycLq
wIQUeqfZSm94XuualC1dnB/KWvNtQXEjRMeCUJ908x40IjybG5AHmPtsB9tf
VVOBdHFGBOXfbFFesVg3ydQ6NHOP+e66lHNTWRW/aFPNLbjO9SYyZ1Vau8zd
pPyyaBapaw5nkqH0qu8oroK6rtNOlWYr0fq7iGudALog+CyiZ36BeIyvZJbO
0uNPgWM5JlAbYcZhX/sy8lahzXXwR/EJAf85It8GPmMu/vfUarWaerscU0AU
aVqKjQWjUc3E3NlPOIj6aRJ1kBIoS6N7CWjJFOlwvigTHHxc3re0UboVe9hV
IIck6KRCanP+6zrnTRn535kiefwL5omK96gQgRK7djpTB+TomcrdXJ03RB1M
c4f3iucu2PqLZievLmCxp5GKd6e2oPdlJf+pAkAsCd6Uc85lPeDZPKcoXyYC
vxPqcP0FIyZbQCKXAEz4vTFsvvcgT4aS0IXop7UNx2yuFKDhQNY5/QF5wbhO
2fZH3lo6B0AKeXNsFOjElwlcRVmNoBMOl78ohrjHQuJVMlLoiFJlHWDXi6es
dqG+07UcNJKGldTnJxE7pao5Tg/uDA5IzQ8xh2wUO4VB2zYTS+ELtC/fwLvd
IJMx3ungGc2UVR/LAY/8yQpdcYn6YI7gXMc/rgkKsjX2oOIQK9pUSEW4SI4Q
Umr35ygKM6//NatbdhARYHucaiUmfr9BaGDpByakOFuUPWsPM5fw+XKmo3MT
i72zhaxGOxB+eIBFULr967ZIWom+MIzP05V2OcdNLAFjAV3EFbC6mr7MZhgo
xkya8FqHQ8bbk/cHINAZxJOnkYFZf7oRe8le7Sw82f2c+XAdfcx44N36lCPi
0OKSNDvbnqt//XoQz+qoVA5rjoio7b5ECkFpXv5WsVyL4MG9JboV4/Fn/Jkr
LnvJs3dfPX+y3VpYy16SwTEBCJQZoHdnGo5BNz62Oq+KN+Qx60WIPx9L4qRy
NiGSYL4L5XJjKtnIxSBd0QjhigyS57k0BEwKKtBMyigZ9DBZ1AF+4J92Svh8
eYLinYVjQiwvILu6nyANzN3Sv8ntv3xmz824LZtaGF5EvMyUymc6VmB/GFPd
NJIVfRKX0VuxPiLUxHsgV3mJRclqwCwsMPImSANuYZwL3nxiAcTAo3EOqgB+
BWWiOMgfSVV5+zfyV/gQVODy00lp6JmKNBQj8mIh2qfi3RR5CD+NjETNVfjD
e55mXcb9rxrbLbfuRcFF/4sZplVfdLR1PG/Idd7ZdxBtNlqvMHhkZ7jr1WjO
U/gTBuKN19JJGzdDDUz5OmitLZSRIjFl4HzKfeQipbjV4XG0JIllS9KV9vJh
BsDjTERjQKiMGTtKA7EnBNPlTGnyAyfi/ksVZ+QzN7ganojUmhN3fb0bLx1X
lxz+ee97AdhOuzqcU2e5XolMycDTLJJqnmrEdDeGjeuO+9Uh96r5U9n+KVS2
Li6SsAq0+7iucmfhWu02hTO8aQri2bpL09JS0QR03VeY8cfPBicYZO+gZkWB
PV8yAjZA8k4JUyoLSlSfd3XpXwvw1RIpIlBzmgJbBwwyX54OOvbKyeBZuyWG
+Gk1azZCqN+7CsITuH5qapdUT7U7oWhXm94+pVew3fnQspl3EMu81vk7P+w0
KNewLlL2d6mE8R3gfv57hxUnDkWeMbUk/OZvIma1A2JwwSqv3CprvgxdVxmH
swmVakVjc72wdjE17dzwOJgegdXABgXXLezAOCGySOevTRUx/EDxvV3NBwli
nQvk0RK3LTTd8Lfs6XtxMmUbLOkjJ4tta7DuQzBe3fLSsUE7EWeicxZhL0Az
t+0t0N50NsLXe9Q8uH8eg+yw02AEyEV4ksy5+X7Lstx8RiK+gV4/JAjYR6U1
YsoHdTirOjJapbnf3VmxhDtESn9CNxoRNLUlqBbK4XQEErlYDKZtFFPrRoJW
z0HTSdDP9QcMyI2akDNgjeIfjoJzELEDIltNF96NeVMpka+eSubnF4qXQNT0
xPZ07QiRUeduu2AB2LqRmc1DIfeDmpI/jJLowhjgKz/W5S+59gWTDss8jDFo
h+9VhvTzlPHf4PoA9ajy/7+zqex7PnXgz46SOafbkhb09oLGuctpVChoXRFj
DDUu3pUyiU0Pv0uaM72m5fEH33GTfwIbJB8U7nCuNzKcRq0Cxfxx7kAHDqdN
6NEk8Ru4uBtn8cgT1UJiQiAyn9PMrNsSc7Z/6qrbk9wd6gi5wUwLpALRxAps
7Xed1lKTbn11cRn5wz42Tg9UQOcJIDjmViwxrTuwwiuska9iLoMFY4cLCSu5
GVPZpkEKYEthSI2tyqBw3LO6ARDDV/SldgU2oB6FlT2xcvSAUkVPWRjzDZJu
c/It87aRw/+n3m/YS3szQAfj2QRJ6tV8uXpemCZYMWp/Y0ot9wnBllyPPQAa
F7Xv+bc6bMHw0Ed4VCX36wkZ2gRDjlbG3b1YkV1MQJz4elRldllLIEaUlNVO
lYKh2kU1H8O1uOKg461v8LN6keRcFwVnqItaoRnmsO+OPpNvoMKLgu0FhPmB
Ch1D64kvBMEYYQokbAclo106XO2LF5rTq13kFqjVlrDPOlswzvgPq5PWlNlY
Qru81+XXP3QPFXKrEA6LCL8Qvwk14htEgElKeb9YiPX4ZU3tfzGBfAO3Vz7+
3Q1AzvBRtTbpWIH6jAIJ3+ZqOmZ+kPPVwguz24ienTnQjFRXp8R7yIC6iMJU
WgGsx/YY34YRFjVOfCh59qdXlFpJcMg/aQ7RJ4GckVcyAVkCDnXNn/OVpCVr
ZjihYIVPFlIPR5oE04FVVb1J4eGNpRAO6ORpEH+oKaOg3kXQ+epJHyhdj6aK
SK+UfPWU5D5IH1ZqnmB37A6lC3tXxSDYe64TS7Wc1Dd6K49bHdGAkA05aDhT
i34/9MvEyUPj7/mALStZgJgtaHxIbH8k0atd93uWqrUh834lze4Qg81NQmKr
aslFCHc0WiCC1T3Q203M+HP5Qj8Xm8zp8g5yxVNlFBr68XlaK8A6ovqFy3Fj
i0WptI2sRoi3MXb7QISiisdwrExvsG0eRfEH8EXzpS8WPenjjnQdlBuEIsDq
IQnb6GM3JuUxNPaOBQgRlw7ODDaqI0SKp2bifRq833ejNSOV+aEGZIS80USh
D2s2jQBukqSbDI2UMMzaOwuZGJfLn/GeeSH5CkhHX/Ma4ZwA7/VuoH62yic0
M5zDkM6kwIWXAA50O4FLb5ufgyCBn5itIJjbq1ntbZLg2JPZmAaNkLYdM5t6
4O8Fv1GnybXViy8x60Qi5+jExxlZDAu3o/rrgAjcsV316rO6YfKG1YM13Xh3
Rs7+AM+e1mUHICjfuuKeDTjKRKdptKybhAAZ/tkaZtYX+uH61hXK9heVdDUe
d6NB/NOWhG++3Jsxp/8YZSqcb5cGcqRVLuu6xCn8PpXE3MnLxm/Q8US9xw0O
88v9PObKa2kAItYNfQtoEN4p9bzvvWMiR3dq+G+ltJ4ZWoSxS1egXD2ucfpG
HyHYTxkaMoMAfz/g9OOVMIrizWtJVMU2lHlr4yTK6V/oCu+Af2GWpCY6VzUx
R8e4JSLzxZzPW9/30GPphb+RTrl5f1BhJOuBoTAgRFn5uvL5lgoS8UFAEkEy
ChV3P+wqUyUOfV8yBLpn3LYxDoMLC/i1AvRXujxb1V2ONYZkkvVt/g5rp0OE
vRk3suNsh+R16W0torigYPlwfDwHTx8+b2/KKFqnJ5qBALHtqJYUTHHSJEYo
uiyXyaD8+/1Vkxgv10UzWvtomv45Yvf7peSrbm9j+NALeSvNqw6AoZLaThAf
N96IeH37pNuyHRDXO+tafE2Vf1lh1l0iaDIO3OGDREB0o98dNlT1E6D29nPR
/g/Zt1RwrHdb8/21FpfXSf9QgT3oonbb2l1IzoD0pmfXIlIb+5dF3vJZI06F
fxa886TTsvD8hT3p4v4HAO3r64o3rx2PSH7z+NBwDX03aNeB3NhqYTCbCaFI
BTsv7wasiTg7XsqaWktgnLKggAhnyIN17ijRh13F8q/VHahHGHhDVh4+pYxV
5AT0wRtCNTmtihKCYQ3ZCLtYXEp/9TAdCJTtTJTiiTtY4b4tGUJgF60wqGnD
VXa+6/kcv1asFcU1HgeRXRsf3ZU7Ru++wQjApdBZtwiXcMzNoZd4b+75LEYx
hd84p27VJynW3n5mcs/9SbVAYkfs9a7GlMbsBKMs7vSztkfiTmJLr6XtpnWK
xpT1Dy0c5glC7MsTLjDpSadyA2vXPHu5/oQ91aL13CG4fGGPG28MFnvOnP5E
0RHDXA+gQVAebtcb8kHkTaDdKRfzd+f1xQNPA7cdrpJcQMiGkTAH3JKACpGM
CBtBvQ9yqpmUpGUlczK5RDyZuNGs1/q8kugETGea9xE/QpHaONFc84lxjIm8
To8iCyDjOIp/lOPTsp8ldClPPDFQJk/jW5E7nHntwYaOWNqB+CABd0xM/nu6
4uuqoJTQ5I5FCvBWoAUBpMoRI7SeyWwDK6zN+8kkHKr5fPlHd8/zURGPnaOS
jHvfG6IoJ846+8fOoMc9wW3wmdoeNQ6b3k3fJd2s/g1pM7RlyEqJLfe6dgQt
I8wP2asLGTTLY01lAXtACzj/xL6O7kW5MZwS2wl6F8TQgygTog9nbVgPR+0M
cd95F7mK9koBhJ9TKuh3x0fxPM/EHefEDAhQn2LZv5Uhz8CmTP+IjYC0DlUe
4JbiZpqNR1hXQstVyjt7rHg6mchFJh25ZAtSXn1Z34KnPYqXL1Eey1v3rSoj
JYQMei+BaVWaHNKmvRgWWIPiI0zf8JMhKlXzEyfoJi4p0pIWyKHhNXqUulP/
kHbT84obCUok7EjR9PE7jpcT7ihj6xd9AtI+Lu7sqI2+h6y2O27confog/5I
UP03nYNGNCRmVK47/2kSn5grKZXU5ztwhNwrdEoHihVFXJXit2I1P4tIybDQ
e9HL78Cj1aVKSYUV9gylR8OTmv3tntCFxVPg8HBuPJjx4AUSbioGPZDZ92tS
L/fL9V0DG72GucfVMG9+7nC6tfSb+ONDfCFmNPzoppkdfbQl2lAWvijkW99c
ijml0qiWKzdhzMZwOiNyJIYvGmcWfxzfvSmIeoTWJ1enMnHduLJu3kbi1Vn3
SBJlju3NkgTRLNz+aTdUVwwmOavIcUnyDQ6qvbx7Jbc+mxMP6e+nwBpQpQfB
8QfopB3GMIIGw8gtsvZHSxmlhfipA21LDuwxr9+NsQZlckMkG9xv5AX8/BsB
zhhBVOA4GS4GU5g/+ZUvggZFoLYFYuwh2MYOU/gWG8CzRfScM9yLeIP6xM6B
nG4MWvxmOpDofVBjKH5kZnrDFzwsiM/qJOAYcP6HsZ8sc0rWSYLteQPo+1EG
/CtJGSAtM3BBdqcqisOmEgt8Q8kjVwHdN1W31fQm0pF43BJHX/Ac3gcn9GWU
R/AqG62gvF0owQPKcA05O9Ggq/wofeb0ihH5rameFVmLHESTahC0af81D0+i
InTPw7Bd5SGKRGWjVAFbzlrzYLzqZJbYhY0m5dtwY/RwJwFpegUG2muOiwSa
mdbc4bTY3mcg5eq0cfGmdHpJOqqdYiztYQdyD0XSD9OQyVNuKhY+6161ZiyZ
El2N9V6iDR57uPpWbENcvnm/l/61xDhjDJa6ri7/wGY0u3w/A5dLYuINVXHW
jrkX30RSk4E/MZCD3ZKCUJCNbqQUj0BPat8RMGXtcGKRZEegjt1shJzvwJQm
NtvV+EGPI5GWiBeIwTu+90wx7pcsbx2i+gRZ/ybiVDj3xzdN/++Jx9ujHKqz
OwCQgBMnHMUAmqb7xeV3VuAq74RrXT99+FkgH4Mc/MF524bFchNIFanpYG40
CuZutOj0mUL3LbTGTbF/s3HMzZ0RbsHoBpmESiiWT9Xr7wiE5PRZUflae5SM
XFh9NkN0Z2OIIPi9CFqe9tflp5TeYfdDUXztPEn37FgvkXI+pkgHpQBE+jAg
l5Wyxj/KFcsx1QmGOOZrIdBSTJX8J2sH3qHgLbBlXloXV0MKDdq30qjCbbx9
aDIXbIEOzAMqHwswg/lxrZKG4OYJ1pA9guSQmirUkofL9yvTl6PeoDKQDQ1M
W1bup/LMM3q8zahjXLq4K4JWEXxtOKbOi7U761JlCmoWV1pqWLj8kbmx+F8Q
h4R7bg19IiTGCtU6YmgfRhtHMV7qZC+REM2bAeclPMQtQl7tQo5dFH35WMR5
njSUYz1h8eFMmoHaK6yLQSTxWl4kCgryVFxjEOmfkwXgkXmMeF8622RSSOpx
ir58o/P9pYEU5VQd6IqtnY1EmVRGHyKqm28HCSZW8y/VCRAHe2/HdM6PJQSS
P60FyXIkbtwQcHE1uy3r4KI4h3OlLqQRsSWHRi/eF381f/sFKi/I1QxvZZYG
RsSS0WKTOXNXz4/ZURMjetu3CtMb8zZsJXgJZNPjdCwfcOqTDxT1qOKQ3ExA
u8sXyuHvWFsYz9g5IBnFJOaUolZUoFuM3JthBpM5yM4KJ5Uut4dzQA5vW4/s
It6PGabB45YOqUwus3iUcP6LAm+v16d/mdYUtunjw0yfOXYgtC7DyBPtWOY7
sYrRiV0yndpbH4eVJlzSldCOTE9heGZLWswdx7b5U1UvNSFwHi9Ooul+6bJc
5zL3kndjlpEHegPWh1u2KJla65Ob8hbKmGQ7XkkHVhJxZK57U08F6y6k2aMZ
nuo8Pti/QUOqLzzSwQdaEXvoTeK0j1GIIWDzn3dFVV4EXZBV7vAlgwh7SD71
DSPw/XCi/DFWPQkNGEcRN80CPNp1cksmH/5SpN1iBIZmopvSrP7fQRuOwc+D
QVdts3TgT+ioWvq14qv1XzOfrT23wD6JRVEhy/ghaumqehnRLEPLm0P1a8hU
FnIhkU8Ojo9boixA9eyFyT8+yj8yiI5ztXLsJdc3Gh9K+jSfU9bbRuIvcRfo
gGtKep1JwwV+QYK4nu0STo6JIC2XPtxhnTFWbVXKDMPVMe6zEl4LaonVCoud
qxnyAWs8EU2D/798laufsgtCw65yWJ/F8vPo8mM6hWRRoorGXaOCoE4MH3hz
QWZSOOKD8yO6NoubP/cUfyluBBL/2LMgZALO6VrRIJY78GFJNTZzql8co5WN
9yeNWVOLepY08qcg7Ydgd+MKZz655IOBXJlLx0hqqfVFnqhkQl91vTtVOljf
WFriZ0l2LlS8r21ArPKVth27FY/otnob2vU4uPl+zNqacACxRxIsO3OQAw/B
KVa8HH1WK2D7zJl45Tg5N3WftOCTHHWvEdAscaNUD7YPzkD3jIblZYw/iek4
hzR8HLvYmbmkK17Aw3f0Ef5tPd8Jbz8IzJReqfdGp3H3UtPsPvRRYrf9rG3u
L1F4IoP5ZNrSCTWP2s++eMuz9SGtH63VFq4YQSD9iQGPD7vSYu1jpxlJ86X7
ml2WIZkuViq7iO4O4BrhnqBXfRgdKTRzsfqRok0LsYjX5qS7L9/AvFxtmtek
rwauTRAECkgWxiND2XzRQc+mq5GJakErtQBVTt9F5Xf4NFJaPlb+4qJsM0d2
tDOpYqjxHZt6CQP7h8SUJNi7Hbd2c74nrZPImnjNiE4vgXofKQlU58vrUfQc
sPGai5wuVupBuCb/iMB/+pvfz2Rs9SZ3h2VbXDG3P9GyZNCQh7uHesxYOQoC
Vxh1xiPhevwmeeBylHOSLPJA76MC/BpdcFvNPs8EYylAI/+QOqehKLOLPEsN
JZTs1Sv+n/Zkxrgy+9D0ZsEmXiG/inFmybQQYh78NNatAseGvsB0cFmLgxnr
B+5JU3zsVUhppmjvtEjKqDP8VEw3YGrDvLH08WMXBodA7q1YiWkFYuNQX7pD
9SavYUIskvix2lOwCxvj9UJJx4f7ZiXHCymVbnqlAqiobvKMYG4Ac0OsRr5R
LpP2g1O9wtnH2QUU7tmcCfnO9qyvJSxBR9jsjQ3MDUlKdp/8bJLkd/x314aH
o/T+1evwBWYzdc0tAiCBbL6rAMu/Vx58WkxwneVRVYTUmSL+RJVQb6HOMgYE
gS5Ohrt74Iq7WgkNqKfjQNV64jiAttXen3/OrGe5d0zFhfnmj3SZsSV1J1Y/
ugNeL3BJDwBKbu2+IEhNXAp+iXOQ2PJWX5xbIYjE4mE5xGzUHBQQY+ZTgHbh
v4RG0WAF0LShGYcISdNmzR4h2ljr87BZTgKrS/n4gW/+d+i+Gm/hOFITlbuC
zowVfnmCsoydsG2F0wEsVM6HiBYzEKnGtTDD/lFXp0OWZpb40dMKzkkh6rvw
AlrVLE2HQmEfa7D6PgIYA/Rz1kWLf8MLYDQ+7tLJlxJxVoX+JKjqeWLROPPq
P1F/Bf7MlqPcaUnnwlO1otHEe8kwoyO1tjgVMPP4s60yg9tpgTj/z8hv3sAG
Q0P6x7kxxtydq/y85yk7zEPvg62CfB9o1IxCBDcrJDbYg59upcwwfZMdHlwx
RUtP2vb07QKQVWUi3rXnl5i/8jEV8RE7uqGZlouyRpjn+hjdDVwgMDBWqwz/
43YODN7bl62Mj4ukk7w29XgwX+XeysplS/vyZQSq4w05io9oIaYvTHxMIfEk
iICmxqp4mrW4gIHk8B4wJfk8L523o2WnQIEqWxBMTrjXiF6Jw98m/1LJ65l1
R/qJjYd1JdatZQLzk1eWsBP0te9rRA5XRS1DynY2kfaRoV3bP9Vo4nOQC3BM
JsvkY9Z6nHIVSn9vElYoCMqa4Ekg7UEygMkA63PQ9en8OfxMHnkyr1UXlO3T
YRVWtNDnP8knZIsAFHRalAqN4M/CRSnK63zA20v69cOkOrQZJ9H81aeeOHda
a+/19SY6lupvybF0AX8Cb4GSIF6NeUPkcS+slb+GUmDxTb5NAyDeqpX45YJ1
FXp6twAy/wNByN9dy1dVtKxIJUGLlKqMes/3S3PRN0ppJ2hfyct5Nid1jOhJ
3o7eH+doKO1tKrvCAVm8pQMzHPoMXfqQKExao6Ld8s+zf9zFhPz4Pj6qaemF
a8AywhFcAQrVzzis3+1dttqqE6ENv7lQdrPuiXyVfgpIHMcL+imZMqVyMN7L
y6hAUmFVEJZz1beKiF3hiu5cVlFj7rzWTHG5tkIDha6LvaCC8NIq1z7N5W2G
xprc5C/7GvNmis+TpP00kbGDlSvk+rgs7Ylq8dbAT8j52NcQDUU703EF6wZU
f912FGpbgs1nyqkIrhqkHXssQ0V0BuBWU9njc3k3eCLzSgUYb1LL7nR6DgE5
m8nN0rxjxwBW0v3nvOrkFn9GFUeKfztVYwObhqxmxj0l5L06Mce//y1kCnwx
oyh/ojLkFhHbxvgHm3Y5yF/MgL/lcN2b+HE/1k/IC1m/TzKPJjuPBr01pplE
AqOBkJlkYtCdWkwCUe2v0jbqJ5EbSoDe+clJkeAUCku4UOdX5aTq1Uy5SJJf
cpl6L41SZmcLqtPPmN6fQD9M/LUIlUhqRhjaFHvXGmLQdV429C2EiMfFa2XF
bYP8Olz+ZX8/FqM3Qoi0zMwfZitwe2K0oSgsYQY1rvyXkyzLf3a8ZTUIkhlt
EqlqePTg7ybBBjYo3VRH7vcjrpeM0BAR4EoatkOlQoFbdnkakLXQdGAvt/3K
3+pAqPczW9FgODOMDA/QDnFcTYznQCFyRdcShEp94XQDLn7qp1v4Klta7kPR
0z8fc5+tUxMa20pZggq43eUkTMo8VyfcQEcPBv1wG7Rlm7EuGtEwcjNklxCG
qJifK1ehwVrEl38LP5V705Y/u2uXl6rvBGGhmB5KJqW/UIudHgmXsFrvraZ5
bBAViN856E3xc/4kO3UGGc+rAX5X1k2IS+WTOdHCP1byque9Q+mVApfTP3Kw
VVC8m3prJUD5wfQMthVaHS1Nxk39thI2NiarRdczdUb9CpRCPEz7TnuU46Od
n/vN3ZKPjclICaNvyqd17yR4na1rtWIEKh2tdwdkpmUsrjtQmlvtyb9IcLT4
8mqPnlsrPB+uA5fQHACB30Wgx8hO+U+mfkjZ6aS+1/VBL8F5jIZuz+cynAQ9
hp4GP+NCQCjKx9yDO/4dUibSC4FAgaWfTma9UQs1R3MNSC/5x14Sv+i+9V9n
lmDktvWBYo4biYDCTAGPdX68ozyqpm366r1iqUAcMaVtjmiZ52ECNV095BjU
+nNXhxPocDqO8FExKkim0w9lylND/hc8rneMdCNWTwF4ij/N098VPoMAi108
imuBPku7PrbKG8Ey8fDxK7xCSuYN/qhAJ+F88Yaw8E1vpQKmTBMSPL7mVbsK
UiC6UKP3978adY2SMXL+wQYTewHYLreSHxsgWjeEf32g2828YY5EKca1jUsB
XS3vMTAjYgF7TYRHAQQ6xE0fW2TVZBrB44aT9g0WlwHxZ5W04fYpG5O/bYw+
C0UPSBWCLm212xqVqS8KoAm8iB+Ii5FBHHlSWCP+X+7uI7x66XTvQ/1IACEY
LfTDD55BKBxKe3B3zhCXQJkx7/C3l998FCgA2D5U1bm3IihMzdeD5RNFc2CJ
TZnxpLRhq+1fa7MedRzB3UUuTk2Ltls+gnXSTVnUKATx5pa7vBTQNat9gFN7
8fizQwqTA8Zw+dpwyx025yLgLM3R9nQ+6mkdpP9dt3gqGSMHwnd8p9Q8BAym
1N+Wg1IyxU7gqt3yHlsDbOfWa0nqO3UQBIIhBoxcNIVPhK6446sSDVQdh5OK
8Q9x2fSmhFsIbl6E+KsZ3iL9KDU+w7IGsfzNYKfCAz2rxnfVpNKqEdr8Ctym
QMJHwuoUladzR/LBmYYLS1Aa24VoOkWWKt2AdDB8bCQKYsvq/QBk30u3oRD8
dHipmuCHJ94IXUWnRlNV6DP0J1ymuEggZgWkd7jMYcDmiZugLBoDtGaMXqTB
K7/fJn7M4zvWbCjsMVBY15CfA7GTALNaKGkrel0K7k+Vp1RIqB5ZQJ44C/bA
/2gZxkdtbatqSO4X0cbhsDiFN/bm0bRonYWfoTfznJV1J8i4FSm8eUX9w+M7
kBNQIAgOYqIcLoZbFPwjqNq37V/ygoIXgOelD06f7RXi7gWHAAIL76EzTBEs
rdw4zbZ38uIGcka/bnEizI2wFqQ0mGfxPFt5I8R//p3rLsEkEgw77nf9gYQU
XspoWsioE/1wrO0sShscwTfO6PM4a6XNfZqFXH0GyjgbO8SxrV2z56ZjkphI
aIW9cSL19CT+9kEqdEsZTGAiKpPLevYhi2lb+R54beMLwvOHjfuKZrM6bmWt
Ol3rrrgtFdOwBbsfxB9mMujKSgDcnZM8m2JqMR8LkIXPwM4IRAJa4xamk5n+
lzkYiZzn46KFp6AQCbdx/9yJStEcCgy0Gvus0524kOddAUDxqpT/Sp0rGJbS
7vDn9ybhkDG/n0gBypxfRbidWc5g3ixp53VogWSINniY69BO9MZKmZAw7enQ
DbzJOozmCkMd9IbseBdxiww5czlO0R55ajbGqxNUIrwJnR9fvGjakt7EYyo3
2V36nINZY/VvkZ/XgX6+g3BecZstRpnQRF1LHhBWBjEaNdU13xWpAZsDNhus
peVfu0YWsq0IMlCmsujo87uNUKHpUxETyDp9HZ/yxfs8RSOEZ0pq0Q0IMszr
nagej9Z0Y5GzkxyGKXIjKmrHu9zIxnEjI7YVgJT5hWCwwWgfD1+Dxr0v89ip
z+1WilB//zUo/JAKGRMTDEkaBxFlHym8ovGMRrBHweNhLEqZHGiG7yv7KDyp
FbIc7346eravTl4UBig/uTNLkvVcv8LIlGukAyHiNValowlbmgC0sWqifng3
UKOHnkNas368qxsjQZOgwwfC+1zlfK4jEGFvziOIhsy+EAYUCcH1MqQKYQzS
X4AlHmUjyw1xQ8LRORET50PQbwVuC+LCDIkxMdGQzkP66Dml8dWouRoWI97Y
q/UYc6NrIbbBSISl4ECmNeKjJsBuWDaigsVaAolUB9p0DIkmq592WXMa/att
84FMtB7iH7t/8ejLCCGs0np4XhMwirKvRFfqS8XxfIogJlhX9rLj8o7muKQK
e1frE5ovHoMHUWN8IeG8lCYqvh0pzQE3jiUc4+vf3vKqZcikRAYvcD3TkObX
BmJPCPMRSWhUtdmQbPfzedFuKrd7wwP3csRrmws4Cb7MOL38RJilg10u7Ng7
zbfRrFHTH9otaz8YkqSiQB2wsF9ncFoX2RZAx7HJV+2bxei8JDyCFFI6AVeM
tB4MVz1HZa71QM/dl1nXUj9GaARyoC6pZS+eXKNbjK7xCXNRLXQnnt4JG9q3
5qw8Pzi3EuO16nAFIel0zzxR5Lz6VRXuY5MQD/pW8sKYEItqqSYfLC3jFLRk
bbRXwzMX0yvoWpGdh6UaW6qiB4Bfvdp/FcH1Yf7K+8oe8sm7thJRlFKM7yjy
W22dUUD0d5qRnwWZCWpCBXt2fY7foZtFd0nxrnzGngxGZWCEH3lqvFCJFG3x
9tWA02PL0ATGiF1oU+5yD4uktUWQMICSaa0aA0Ge4XLyCmrkeb/oHuLVD8LX
oWoaqG+mhjzOuDL/BnnKZjdO6WJCe1T+2SYUSwJ33JhuuMixNKDssKQXsJRH
1ByhecLanyIZZRtXeyRfFwIRWsP5aMMRk6eHLfQKR0zvOioBYQFFCFuTdRGh
X/YXAxroFWFUvKDdDt+w9kPkJskIi1addYzbQM8LcYpr+hJCS98Ik4O5ClNw
k/eumFTHfRSCqv9gG4t7dRRmZlS8QDOyd00h439CRtuwVcnAl2rhJpxXd+6k
8cYumV3WkWniatvb4nhIIEk7w9rA0gX8/LCMqCaNrNIhTn8nteqVWe0njtko
gBNcUMx/zABNRMEyW/Kzi41RKep3d6N3lJypt83QJLcytR6eSsM/vRf3LZf9
oxYHc1w1TgasdEFSLGOeiXXBZTODTfCAG9+Q2Q6YGieiVGs6EaGd33Fg8sDj
bQfXS9PGGJQA4SSuRkRGRYOtmK1O9+P23w50xSF4ums0rv06FQy63420FnYV
VV20FW/ole2XW1jHmxZ+zaZXxZnvdTaHFPvTj0Xr6Bo5L3iSijSdq/xIeWMF
BOpmQ/PStardpCnn09zaS5moKRSTgdsyRts1KSspRNUyYbjLLbE3T33KGJSz
acj8S9/gY/nTAUIbW6aLuM3jLdEeijwIrJFQytyf8DvdzKuJqo7gn/iDLYwL
M6DsQKdTmsbOxoazkwCCBmhkIyhcAPMBcGDGuKwT1PaIP9oReg9hin4HJUb8
/VzxIjJjTSvk3yUCzIHMmVt0Ya3Q7ay5D13RAbHHSRhErAQ7Um+niJUB+3F3
6A0q+NuFw3QX8yRwbVp8SSGAScDb4CuzCbmdA/zZ1HQ6v+2dbVGz2G4UpVVe
j9XGiZLJ+V1EQqTLLv8dP8juWB4XH+1zNzju1Ce4hj0NGo2iugrh+erHKO0D
95EXUlrymsYT0MCXhpp2/nef1uKvpxdHDrkFcJ4f5t4VcCWucWhW8VIMgPPs
xDpYu/M7SzjqWf9j83FK/Q3bYRxtMBL01OADK0v1BeyBwOoto/NNzoORCUeu
pElQfKZYGwOdzOaK5RZZ+PwPGNoeIFX/fDTX2rE122djzBEubNVWPd9bWVVM
aJ/spWt6NlwH8Yy8OFHFNweW00RALG33SZPy9+qP+lUWj88RHex6cWLV86M5
2ta9eAO/+cXpaWskhZGh7qdpx7jofsJgJRUFfMulSB26w0YYLf9YzGq2mKEa
PNh21IvlEDjf2+PHFC7QbRaxi77iK/7QWSDWoMoUJXw3JEnCKpHhODSZYmt6
pRGEV6Y2Q/Xzmn/VjR/WaWLSIFKjJDwtVCZeo06AsPvBPhvFyA9H6nBI82fV
32NyG/WRQHe922NybOab2vcTsPfPNoDmqRcWK6+lcttAkvJErDeX8FgYN5X5
4cmZEVh/1cCyWvbr9rcYak283LZ2+CcqJSf8oEQf71/mmH3G21meNzaaMlmv
Rw1+5pt/P9MlsH0l5PvGwdNoFQvZXcFWIXw71ttiKzyJVKdglON2jNZflEyI
C3OXTNBoo5YG8Btf1SsaavH6zVyYvSL4daL+BuoGGRZLKnrV71kSlGFWHJW+
loSKPQ9BcoS+lu88tk7WMcqFQs7gnC4Hq6K5HWCvJgSjqLvhVy5Xe7DMjQvu
aRTiQR0XasUPIsBT0cgWiBezApKuVQbaLOJVFo3Dqz/3f6xoQqNbm98WKCo0
NAhkMdV6AbE1sT74acjCzo4wYhYqieFO98OJDwlUrRvPazEDAfd6XVrXFMGb
UogmOPhPKBtPK5bwp5ZSi69HDtrPRXa3LGyOoPXuq9OgVjpTDtFTlojZe2lK
RCec8sSFCVYS9+frS388snoqR3swugWSMxFgJ5fJKIz5r0BomSLZ+j1u2rK0
PG2XQ/+D+YVcQ1BRz3GuAAjNA/WGWJcNICADC0nfpVpaBLy967QmrZs48sk1
/mIf4LTusIC1tO9+ZYOFyVTQ8LKjhytOZHtI0WxBJYOumnYyR5KB+iyeWAWY
rELHe6Hr/sB6kAGkgIRuGONlnr2+lVCn9WxBl2f5eNqFH8wLonDChlG/oHym
jnrxKPW1idwznnKC/zSww4A7IGnN4lmylFzYrxxxAzSZS9f2nSpe6GtkImoV
IUzPNdWTzAMr3xt6mN1IesXOT89uaP4htegh8WX+Qh2XksBvM7CHlTn+d+rb
iI3dWBu51BRvRSHJlpFjZPwOaZMbLkEN2+XjPZAf4JyqF3Gh4wp7MkhIsiZQ
2JJrFrv+HEXYqsgI8bEtStWkJFJNbjnz7QVH76/n8nBs3EROB32+/YwJ4qMp
adV6RnprK/kWcmho8DjpxpFs4aSzEKsUomM4DDejUBk2J6y7OdTyX6+oanl1
6L28tjhZLFZK6OGlCF9oW3LYZHMeV4+8/btKelF/gK4DBbp524Bpbd+vJ03h
Zc+l3AbeJWWZvDPPuwCUeaoaDB56zm6srExsoEdEMI9QtsHI+xij5v5xciot
9saezIiqH4wS/kx4aoWR1vzsXiDdDu9wxNvj7JpvWP67HYgbgNx3x1Tv/pRQ
MSWhITeaOh5b0FDjoVzsGQnaeSlgnNVXWJVP2kOJ69Qn1lo/5eIaUdILeRfZ
ck6Hx4zJcXr6D8w0qPd5hEGn/vakNurfcuasnGNzBvJNndcq8BwgDnjPS8oK
Zn148c4Pl29WJPGeVwgsQBBafNFJtryT7xlbeezfak88Qv7RpRKDb6k17S52
jxXAH3oDA5lcmAHQVOyqupsDq33xhdaXRfNErJRPcjYQtX0QxU1YFu3eblve
u+aSSv/zig5iLQ0nrrTeYvnAhlZKQNlTgm3jWH3KwIpiHJ9jWEVw8nLyMVPi
JdxQkzFnahZNYxXGcWMCV6jC46QEzEHxmgOC9OKv3mPATu5Mj/xt5nPjzyLl
K39O3R4KEhs2HBNBFC/p27skioYSjtY3HO9Jyiex+9dvJGR9O1PwG/3b+Wk0
ftJuforinC9qQ2KerR3aTrw48lYMRDKsYXSU4s0+IXEOO0IY9S3qZXss68Zt
v1L4wXn85EusqxmTp9bpqD5ItdyQ8t4pXps+p95I0UcerRLAUdUikwhQEQ3p
GjF34UgFBnqBYcYHm7NUyqZhek5YdlOzgSKGEnfYyy97DEy8IInhL7bjpd69
dFtk/yLoS58GCRkujiQrVGmTMvwWrvBcJjLf5hMbrnKLz5C1n/ow09Wapnb7
uVEXkt1KwngR4JiO9gb6Pa/Ryh9cf9heVGXE6z11m9R6w/6wBszdM+9HLxu1
IjGXlptXZn5nQgcNHlRhzO836FOY1s9Kz9DDNMpruwE/zShmIRcLZ94aRQro
77d2QdhH/mIttTKvcTlaJYadoUfgN+VwSfjM2bdoZr45aWJs2CzFONNLF+4g
fpUGYxHPRq/f1Hr90L7LmRhZT3ebuDRUOn+RRJUyVfLS5JPHxRm0F8LwaKs3
p10F+y92Cu+1kAKgKwyug9T8bsQyJKO3EflK/99+5ZMoOT3f7mh5x6/BU9Hj
lmNihXGT1RsiIJmsoAdO9uhYVc7E+POZjo2k9IzXsxa9fz7EkF851W9ZCBaR
8XKglTR5Lqom4r/btWOR5JstEI3q1O7iVVXOGRfeA/PUP/92gjnWj7/+bJWq
9DJyoDjIoc8N9ZAE1wS1lztRgNmBWVvX6Y8zZ0+DxFhKxHPwACDg9dh8Hi75
wTmTSIP8QpKjcP3mJb7HQfa2d7vCrpZckKVK/DHp3Wr+5XU8mq7SI2vuvdmr
6VWtbdMsX6oRggUrsqt9L72dBR/8j/xvizlF1GIcEbngZQd8DfisNnb7a5F7
PYnWSkSH9ByemK9uNaW2kaW81Ig3/bYECZEyMI9TZpPJ0+fpesHskS47fmjJ
aWVT2P6/XIJvPp6nbsjqL3P0tncDeLSGJMWB2OMFqMSHyeqoARAORacnaF0J
Kb6bEA+Na7TuWgESUTV2uP2H/zG+x8O4CKiMxwoBM7fgeAwMTMEOD7qaalus
eSU40dKnUd29y0HnTaayJnI0EQ0JzHobEbhl4fN0jcXCj7rfBjQKlUcIciBv
c5/aNXSL4X98SjO5D8KymJZMHVCP8mcCS5/DD0OBUlvXMyyXFuU0w2b74tXT
h5Ry8CawX8n98vOiHnGBnucLnJZIbTPQ5UBcDxrcLe0Brbm5uKl4IDBHTM4y
UUI2ODnc4GaILYGk3jX87zCzkmbh3rRKyitC5ZxJ8Ht3IKfmNsawtnTNMlo4
L7PV7nLu78jOs0SiOj6010jgqkifVid9JZHBm609dJlA+1JdMRSRiOZeQd57
l54IBt8G789Qz2fwc4vzEZIjWL/GtvpP454TM49Y69A0iDpbVMZZ5hi56n8M
cWTD90mvvGEYp+/uYkqkEDIiDf7OfhE9hj3hHy1/Mv7plupRmApYzB0dnudH
xutLX+nK9g8Gc8+swUSnVaex0zTYlWoV5NIpxUhzA/z/3eycaOTvaa+dP/S4
y4pg52JFRcHUwmU7NTIGvFchc5DvbSwDAeRapFEEAsXnXwSP8hc22n1S8KMe
7DOw+WkqBpGPcbIPLphOaCIe5nV2NyHXFQ4MR3KcTAujC1kBiwzHkr0R8xw7
/S1EisfRLdvdjql6ECbSjvbR4kK/ROzMNvI1lS4lbz8JX/YCpsaAvy41N6Gx
ASWxS/Tuq9j8kstv79KeBg3jqTkUGFtWYOsNoQNAx2Bbh2koMiqY71K9yaTf
CZEuRiVphxoQa7JlBlu99DRlLhRMbW3Y3WsBOMDFwlJa8Ss7FIg7ppGrWYMU
TQom/TtRZbiEaYXlhMGZXD3jxgagVyZ2NOY9qm5xd0jXuHI3DZi+4BdfSlXp
kiSUDhsIPBV4P7V0efL4ccN1llkOf+8RL9HpMuGb4xxzlYFhSN1NNgwQ2xjv
xXcgfaKiI7HGoMcLrILD9uo7Ekpj/K/YJCN80hlhCrRrIXzbyr1L1BaMIBd1
lACGcLnuHyUjMXE8PUOK93P7nQ+vv1vrcMYKxFgfV/kJ6K42SNDNLE/Lyt0u
F/MitYoA61SbiFHT2kvxZHbIzBJuYws1++kiua9l77jC5q+UDFocZEUFXtJl
wPxW3bKq5QoafpDCu06ER0PBlCYqCxAcbwWkdAZBnBhLe1HlRe8qPaWRHJfh
vL33LFiCEdn7Z/hjf6UCPIG3T1PrdwpDOBXEkdfTu5uf0fd4+YxS0YFd3lGu
ZBG8ckKenm43Vp5mjSYQxLBYD4Q2G9dB5j25gWT9maBlnbPoX5qrNFLwcTOA
2CVem5kaDKCScfZHGEXqXjB9ZcJEGcz158E3qwoMB1LeEH7WXNI+AaulRip2
lXPcGzyA/RiOB9kw7XdFdTBwPF1ZpYsFEdmbBWQOo8AasQEN7V2y+8j9ZB3I
VanT0AlXNSardun/prx5EHW1fWUZu0HR9aD5kQcpGSg8898n9JY9ds7V/vxL
+SzLzNNh+7uF3WGKlBZxc0HcHC77cPG/I2QEYDgcle//bBgLvKPrz9JlKTEs
PaT9AnRZK1wwy7ElWqSMrIsjALmjQgpnPs+nAlsrfFxeyoM76yQhHzLjHRrz
IIfr7lShXCYFn/mlvLOrv1lVErYWcflVgiVTC93BIANA8EPHjM3hX7/cE4lG
xwJ97zNsKVASIMc0Hr4yFNY20OqUP6qv9qkb1w6N1e8vj9wp/8PzqpcwOi05
ZsP5+BUalUKfMlKA6Qtwvg4wv4m5CdppmsqeyA+Oyr+Sk65nl5KnWAJUIGey
nnrvdlPIZkJw63unVXhPm6e7yTFhDrhZFOcyCpDbmLtF3isd4qb2/k49s30K
SJ2nyfEdtJqtdoUIxadlCndZmiP5uVlAYe0JPH64yOExZpWELTCo3GcCSgMU
sLdeqkq85wR2TmiGCTinCun6bUK9LLM3L5XwBkl495pSnpNdwkOeZAtRdAeY
uESDBXAlBlwBAb1OMRf1ex4m6BDguQPBJqmLUEPkWYI2/k/J4M0TF0wzKo6U
h4cP5k9bWkF1XLZy8EfXS+4OlzDRGzCmHsQU+Og4b51WgbNvj4QjmpnTveUA
BcOHBsrcyN6+S9u2pF5YIF4x+acWrUbENFT+Ig0HjbayElRyjFllR+yFh6gi
uhkKJI9LZOLmmcoqC3LoyK+RjT2OoKNpE4XHN0CvBPGeSnnCrk/0/DJq/7gQ
D8/kqqA/UWiWSq0x9fcBdT6JtnwOb8XxQ8bf7fYp8gtjDjOe34c87wxuF3hh
BnWSQuwfKeuYcVLBHDHFlmiLvmp99CLe0f4RdRd5dZxNbdHoIQhmav+s1yi3
UjcSWKFSSChxb7djTt2IAHKx8mOA25kaKWP2BDOmcJk5VYP53V4LreNNNdho
2rCvEekXWUlgrwmtkAzQfb/lfxZjUvZqZTv3IQZjW34HjPy8cq85bgK/+HA0
1hUMvGYxYdKnCVKEDLv/i/HJLYbHf0BQE2FMR7Rzrc0xqb0wnIv0tZhFr0kQ
Xag/hNnaFBFKRia5i+d1VL36sejPEYJxBcXrLtMs6QAnx4EyobLVKvif0ntP
CigiwId2catGevFj7Ivue83VSR2/ei/P28/05xmwvTs46gIVilYpoyzO4qRG
1u2aWUBbbf4qxtEzARPgg3pypk3MCTE6i18X6cbmy7Hq1FEw14hMUy2k1R8I
JkJLNsIamBpTbS+ja4Kf14Pc4VRq3BLJzCrTTRa50bWORW/WHrrE55383FV5
AMepSjyXgGKNhx6s1j3f73nnWAmgvZDUh2WNfE46uXIdSICguodGdFi+cmRq
5ynNouMP80FQRN4952jqBL3EH7nwj+Ny3KpxzW+OdDkqtHmTQSWUXMN42+pl
NwZbO2Y4HkIuKPagc+2AikIce0ILIm41BhMiKC5W9dM0Hp/VkfMvFif90/5C
8my2ZBXJsK8ziGmOtFZ3dxLSW8e8eJHuRuFS0u9f+rYDESLT7A3VAdAGV+Jq
Kb2WE2mPW87dKOiBSEQKBE6Nxoop2I+StIE2FoLVkEiOjRs++pZr/2EmB5Q8
YiTL9RfWAaPcMWoac+NyB9KwX2D6/HOmPRzTJzMR2SKfRvZ/LkQO2Xw6qgEb
n5SDvnuYt2Wdwb1qZNZv0ZKMCnTM7eqZCkazDVtzsa0oeTgy13TXUl6hZu8k
91urUP31iCEmK4Nsxx4+6GzJw+CsmdeyMbxBVweN2bpJXtZhrGG785NtEffx
jMtkArcnDpBbhqJu1zpEwf+3/aCMKFNApTq5/x9gT1Ik497QVgXLL3VjFqT7
AIPKugLMousTbeM73JMg/NAcGa7HMJgOBYvjoCl7bh8HW/PXjN/BkHWCuVLJ
u6Z/dAKl4RL90BMGrfDLcm0wc/JIONAUX0IEM4Nd6Dba39Fwd500NmsfVQh9
LikJ6IgPOyIjBj6J3njfO+QvTJ8kwy3Els/llGLL0gFqEegSUPhFNvcfkP8E
q370lJRBUXINYqqdA7w5xlQwuMUsptVZKJKXGgqnXBfR8fW2ZwwFlQWrrLiX
sg0LCZqwn8WMUlAHm5L84G0YfkWwg8HndK/OJuOtaXRvQ4dlqAh2tc1hDIwL
pMAxd0mCq2Casjda24nedPGX6gj1VFsDjJK762r3VT8ALX8C7mqpgSuWHJih
1XWCSGTnkCUApK++HEqNkiIoQKs2MSTHGOlcJc5RueofH152rAXA5ZJ4/E9e
0yROXxFnhQMRZ1JUdNuTWQc1UavDXN5UO29M8Ecarcem6wwehRNCrHX4a1Wz
X3ZcEfAiawyNYiisiKxym+mNYlnCorEOVloS7WrN1RruE2jCM215dNw/2zet
Gq0teI0Cvykido7GGjey6SNz4a3PQVUpkTiQNcKT3mitMpaxS/Jd2/avqRI3
+LiNOFIygE/xOXR8o1tr4rZaTBk3eENaFrE5SC9KTrTOYKejqM6TqRRl5oL1
nVQve5pvw5KFiBjAGldT6KLEoLYO9tLmvJFO89pPYGjThzVRX20Ucu07UnNg
/yjSj9qJneQV+76g+kd5Qu+RP+jns8udjfhkFaQauV5JPg3VoOxC7te5KPha
QkFhLpfevGWRmKrDQiWvOPsVonQQaqWSp/nyCLOaJHoWKHwQvX6ULPRTClCz
CnV/yeve2VRSEPZ2gFOKMtgcw7n8tDxI1V3Ir7FbiCIl/6H0HULrBwNNafa4
S37E1cRSXYvbCDgvNmj4ua94uvzZvAo0zJhtEjgtp35T2v8PtvlJrM7zIZ2+
rSjz/a5nFR61u3ENGc63TK/L4rDnlK3oiunahP8utnK9XRGg8O3et6TkTuX9
X5s/+41Uv2db1CpCCuYMYrudX8Gh0ELu1cTFlxyjMadj4VeDpbKTkNshDnvJ
5Gg50/6wTRq3HqYWgl2aMNQQ7LMRNPqAWVE1kQSQakMgkEHz+WdsawIM7+6i
c7EQauA/xcSsTto+skwdr2mFaJPyrCK6GTQOjsp9Pu8RSYe31NyWQcTi6/u0
XuMUR44qCzTTOfqKa4QwW5TcTqJvv9iejmCEX0FQZJlIs7Txt49GTgbJr+4H
eMnIyeEASccIolZEXvxCWwHXUEpv8dkqDhPSa6BxgZ3CKFCo4i7de3DioRSP
4FWF2h60QNVU34giIbAOpIuY2K2+fFarc7q/8KBiI0/ToAmNp3hYIOzUswGE
1RBNul0/S72NqqjWvIOpKDWyLnQxR55z1wGFf6OkMWq97DKFU/9jO318xkcs
YApWUUA1T86JIP0gmsCh+Sgv4ZVJ+hkiw114eJIZaXCCsIn2AYchhc+68KX/
oU2SzGyYN33R5V6JJgAY5pBqetNSTOYHs3O0sKBIQB+NzEFEy2kQDv42+hzJ
oBaLFfplRzW1HhTiR4U1KpVEzKGlVw5Hz3hLqkMnN+hrrm105H2vBEZ9//zn
mYYSXwK3MlY5h+M+Jn3JZf3qLGtvfAhcH91ZaTceCrxGYQaw/RQRCVfcAsWv
81H9N2ff6I1MnMCA0gcUF7uV6anRLdi7DKq4oCoJ/KtR9YGQhEeJMpFk0H0K
eDPWkyIlB0jHIS/hnT8LlyB3MIM3EFp/l9BDoDAY9UjYRusnBHxlQr/pZTiJ
iFwVOOwIzErLrCA8IEjDsRhsHZ9YfCjyO0hdJAjqLEkWXZN6pj+RTphqqq4f
4k3/JwbOuk8cLcR9hX4puuDAmwFJOxDhM9pLsXOuRKXiM2TNBur5/TIgCzDg
8Luwh43YVsU7dCUOE6uHM08vAeV2iDkvHJND0op3kypz5W86FtokPzPkafll
/FDRNvmw9ySsan9Wcci2o0KZu4n0M8dzOWScOKbAcVsPuqW6VasdE7i4GZxr
7k9bq8vVG6u7GFWOTuLCOH7Con+6bz4NmaIhBUdgL9fElmdcVseDPaIonZvj
wlp6WsSzby9p1qL7hX+2187Wy00/q5N/6SbWEixDUBBh81ki9qnJ8XEyEm/V
fLjXwewKOLQ6oS8Z68pqv95y03PzQgFZbxTvbQ3Isfn6l9TRwX3VcDjd4idp
EJYDgkg8ZWrYCNEg1RXd5c9lSkKNwS/v+PjDAIeTMkjAuRKqiBlwmCBD7HkV
JPh7pqh14dJp9mNS7+zckqWFA3v8aTf5V0ep+wqaBmVTVoguFV3qrAk4ViAE
9w97kinmMQJ8Ek53zs+NvRYJr2sOWq1QvkhzwOcV0JGy9e/QvWhUXkMRTMC7
/kBGO5hNo6qLotZSGcCmx+2/6iI/pFNql0BC51UthtLMMIq14cEn/8RA1Nl3
eFxAcgKwhqqlf/Ym7YARZrL5gmm/VHrNT7t1RC1LsGmujHVFZIOnE+6KOM0z
4XZ9IWAAS157ACLBNDB4AHOpf3c+Yy96BHL7GoKYzj7NLwKOKL+GWZuwMcjy
/5i1s3eeVwZfx4HE2TkxzGTZEoypWdrsDX82xELeVsDsE1cuXNnWrp1X5nuU
HGgdIMMK+xuCBaOqY0PlFCAZW4XU6ioPb9+BLj99RRdg+Fta/ZrtIHiDJhzp
inNu5YSocQ+js9NSKtgnDymg6xt+wb31vzOSq/4V+eo8/06XBNvrTWKcGlwj
Re27z9KgmVbGGvxSojZjhyytgArldwPtqm23sc+0wdychgehZ+tTw0Nn0CA7
KtJmLtTl2WAkff56k8YkNab1kvkYNOMkcZ+M7FcrH86qpiT4Go9duQNvTLUC
PqTeRnnyO58c9QQMkq3hQw3LDyUoAxCEBNK5TP0RWJCfY+NVavqdPHdlrlbq
1h2rZJ8bynvBAnEh/0OJRO6l/crC2VKpLoj/EX1+HwQvfykW4OtPXOXv1TBr
8K7kRqZJqtpmvKdY1aP4CbaljVzhr7ApQta3mLpQqM4LqCTo8/hwyVZ86qLT
8XSoXD9weJr05S12YyrPseWRY1mstNn1AZp328DBb4nGwSwGgJoxoMxBr503
9YCkccCZ7dv2e/6c2k68gEb9k9FHMZUYaB1mo9En9aZ4bsUU5hZAgSaVU7KO
rLLicI9hfJJNcSkWdJiKQgNIlNNwlrYSL4G+XY75BZzQf/hcj7VQo8kxpwRT
LSDn0hmjhuJnq1CqYZIYzEXPJxyHA9SpAkoiWYa5jpT0d9YIRjFM1/sv349m
0PCovL4mxeNEArDvHR2CDPSEPVs8QETJnxezMsVah+htbl0pMbU/m3TzX2nK
lLmt4Ad8u/nn+fEXgCNCt7tgTCnxolkrwhiuHVe6ZDK0BlcpTyc72cjWrSs3
N4hrjmvapwPZx23PLBLGSafDTb1gIjI2dz2Opd0xHYhOPB2fAtBDPLwyZoPC
gDdIVC1mRlx9jisAnUE03CstQd4NBkwBS5yyyd3D5D9y1RF+k31uXfiw+X9G
CDFro4RIrDed3a/WLtEgop2Q1BIwhps/iQgb0peGZ4WDdBhZ/UaLqgzzNJnv
d3pfrGvb8ax65hHQZLxFlb8GQyJMnmVFHccJ/nfwKU+4KlO7SahR3ddEJu+H
DVMCAxwkbi7lov09yt0yOUphQMt4mYJQZZw0mFSinbK6bT8eEJoeA0QgQv3L
xNu1WDOgGDPywnAKdDcAOu7WcBFu6bGVnMeGorr/Yz46C9nQ1KxevfS25MXZ
kLF5kICZTp4L+3RIy3M/6xfwyqCSRBk9+wtibn+7ySPqju5XSob5UJ2d5OdC
BkvoH5QyUftRvTqMnGJvtk5DPmEBvXtwPcKOsTAOyAnfLVmjXwYRdyNDbw7K
P1C70jQUwIgaivrSieIN39ye7OgE/Tc2VBuWOvloBPME7Rn4DtiCSQbqVDA0
o7440Wd1dmrpUnCpp29Zy1n/9pmTi/JqnANxqaR4aJANBbtb8q/SRvCn4DS0
I7m5AdGpylQeLBzKkVKLdJTdY2+2mV8mzpU7AhS+8zCxlMwbEkY+VJ1GOOnw
z9m+8mUtv0EYxb9uZ2N7I3HtqvPQg37P+Mm4zy7mWsZIeWotijAGb+5CRqeG
6BKZqB4W/Y++DLKNwphjVg9IT1PHTwHJbAB/Z4SkJ5BS+7kxF9sYFlOoB3MS
sFFTGK3Ubnq1cWPRDQ3p4aoa/095dmur9HK7ImN9GUG6gzoXyXa5KWK/gr5O
Zm7wL+H3Rxqk33knuGdsd/2OKHuVf+nGQDNmgdWK6WSvNSxdTF+pm8GBd6C+
89AS7zwMa6bIWKq9TTp5KjCEYWRT47O25lgwn81ujARnl2CBnayErlEPTelz
1d+YpqH0B0GvqHlGcIMuGYslo3xYZo/348d0uyB/r58NZ0ugGgTx4X8IQX/J
6bdgECeB7mWCJT07zdaSjlD1fY91+lITqtQclSlZgvkEZSOZ/XJsST2GcmNE
bkGpHOf31RIp7yQkcxwaLISSQfMw35i+wMqjUM1o+wD1HuvoZbAZJNWaW6hh
Es14owC/fBsGMqb6f9HpqMPhIbP4KSuUVrhS0OuDB9H7kuHkbSpyUoT01ewE
Ks0p9TiizC80SR9N6nOwCUVJTOMuvs+/dYmhKIUaI+n6gWu88WafOHoGLqsA
wDaK4mTbdzZ8+zTW5fm/Z1fOPEf2Vjab47yGgYDO3ji6pB1a6yDNqgUdncc0
2ToXiLFa1NSMQ9WxwBveS5YuDhzb72zi/4samUuUIer/EBlWzEOTr/Hhma5+
Ti933P15Q3mfwI01ezJCXBrl9gXrxZIUBfxCZB1P9JmVDPtUTTiy2RPeoH/r
gDQvD0M4MzH7j7Ac+OjeS7AHtyQCH8koHvJ6+U9AGrGyBQEQELoCSfavGODP
t8HQEPSTFeLhJnTCXtvB/uJFhQRebJ9FsOH1tVwA3JlMGNpY5oj1Mn/JuKT9
xLGOKA/fpkozHRiwq2BpaZUew8IHWdiilU5BKb4+fvuCDUSbOwzTI3cRsVUE
G8zNNlj86IRRrRHpKUS6+wqqXVaAesHPR2UH57h7tF43Y9TAkTL5R/14X0hM
N9oxwhaUeWLnX3XcsDEn7kbVSyKCfxfB3ekdso+/L0+gogz8EaPX6bv+le8R
trbi5SurTJNcObkVrv3049fjZ4oeiorn2Gr7Jue7lEu99ze9lD8QuMnCj009
UEBor4sl64dT96yxhV8YCg8UvbRCHVmayQw8khdwo7n4Kv/dtID+1OrnngkU
rdsSsu4eLze9LPxyZso3M7MHE/5bpLTy6jU0nQApWPmrmucjexYRlYmWHcOx
suyQHpiDVTW8NDC54qowW8mmKw5S3CaPDTngOiEVDGDS9qHtnUzmbDycqqlW
u+C9dtWtzGj3JTmNsuj1HIUoKw1obzS7oQjhnzCWqEFep38TknRhLXbHsZ2Z
MWJKC+2AmvOYVe6d2L8yHcDNSc4XUp3QFrLSjx1MhkSKMqdmzBSZavsDNrJc
aroPVkq9/pSao2w3NIzt2cylknR6v9JdYwUYhsGYimayt0nDZ2XPRsSEnwoL
xdpfTq/9mEvhs5yYPcvVyIbnCtJEsSr4ITZBpuCmS7KvZQodkv8UIG7A/nX0
mP2Wi5BSJJW8r2w+nFqXBRXVduVwCv3C5cLLoGGs/RCY/gZgOZPupQFuLudF
u9SnLeoKdympE7kP8WxqBTENRLRL5iBj3t7Ro7+q8tGmNUPaCAU8t0wA0Qal
sfLZnly7vojBRewoWuIKj1a42CuWNhLnyZWgrgGIE53PtjeKHY89o6IGRKNV
pC3Z5jcn2254qs3C40fEuinXLr2lI3kKsMxYVOptdaCHDLuQAY26Ikh7lcY+
vbNUpkRbg+ASn7iOTolNmbVlNAJTp/+mkeBhYbeu0IbnbBC4s4j/Q2Es20Hg
xi3BwfghtxPGaG7VUk+JBhPd+P2fbWYKhRh4qQxQW21AJIXAIW6sicIibkmf
bawTub0OWmS6FYFUjuE1Y6VnPdGkrX7woLZNpqwFRC081wMDVMg1taNAMeHH
CWNTUApvNhxtJpswqJh8iyTUXf2oMpUOF0qkAuXEyeiDDCZz89YJhgpXulqq
SK65xBd8YG7g2zAC++J1PR7i+3W7aZIPQyPEpumDX0a70Xpe9CmCB6gv2siv
byO/GmO3n1ooGFGojyRITQ0FbJYzdq/8GV1agiC0OmBqbm6eIMgCfcfsCXRg
i8zZ0UBExHJJp9umi5uHcCWSXMLYUvGx8Z3oICOUX+cH5+DoS2cBQV8ugJcX
1yL0VMPRjSEuERYjJbRwV/5CvqgUeeOOICEs/mi9ILMXpzGQzjGAug1DdRn+
bFmW79mOAAps2BqvsSZmOut9+cSCFR+wrUShqtKa0rO9VpwAq7V6J/miWsKw
janMhh6yidf5Us3nOu3xXidPQC07EHesaz2RnTY6rmluFMDdTm6+ZihSFTO5
8O+P9qJa6DCR3No43PkG8pwe5tt9vI9Wxxd5QIaSQ3iBpS7EMxxZCZRskCQ2
c+S0mBxlBdzJ6hqPPO8Ci+esqaAqx+In8zG6zq2sxVQYy2IGNBRbbBXI82KV
OgPRXoT5QSj5iZn4u3kWNPtZAH5rSFpyS4n/1l+/AAOSsDCBDxW8lIRKnvuc
dodEPGyU+FTlmSxa2wLFnmZAVbEmJGKSNFmlxDPeIJvnmp2vQOCQYqhwnJYo
Ld5f2CL0p9vxU1qcysFV17e3qmHSfmI4y+Z9MNyMprBdzjy33znrZaq3Um1W
G+9GZ0w5uiedf7NPowm7JmKHk4ZEL3vVtOK3v/UfeRmffBOihSUxh5ESW9VH
TRfFGrT/7wwVsnYfhpDByRlxSVh5sp4rCtQd26zyeJPjM99z386xpmB7ni/A
7cWvMdROmVQXTb0bdpFLYsxAqGnyzeWBH7PaLK8acEtGFiUZ3eqiGFd6OJuE
yKHK8CiNDO5EhNzJE5JzEUC8e5mNl5qKFN7LE74OTVzChal7g2tZpbk8or8t
R60f2CDa9V7cVQUMaz/LWdDHkVHLW11o5wyimwCjX9ms9w5R9IgfuUV9Auf7
at9yLOr4E8PJV5zyFwAhUhGHDUibybGGlYy0FLBIGj1P3MMMZpU+Kb7ztF/d
vfL5lcNOAtRt8Qkjs8Np5En0DuOvHidd/4sd16Cforwrk/DdJ8hW7bF6SfUi
SohWfFFO8Bn9NpwSkrbimC+MvWQmZMtC4hILEPbUBdbcSZLkB5oKCy9bQ+vs
JBjJnR2K4Xmi0bG05S6nWHYbVj3ifuJWsXTHdGZFvtr8O806coEy7p29manO
S2zwBOV100uAlMCfZ8mexasjmU0kDe1gXX9bOrPqrn4uZRxFGPlUWEZuCDQO
FNc59e2rspksd3HyLrg4eufBOuc8k2CG8Wp5IlwORswgx6RuSqqHn/suSJP1
S1/onS9juhJYl/pSOajjLOCf4rBFkIrLzJw3WK0rPEGqAJKjflALH6PaSVjP
heg5yNs/AY4gnCYPC193mZRn9DrGIXVP7Dr1BxQEsCvSTmV02ORzml7cI1B+
M+SFwXK0xmU1vBashBrAgMd0wshkHneBC+rJCk6io14KsRg1CKvE/ah3ybhZ
QB66i4BSwmX8kOZXS9iCjJZSVfdQ4DxFXy9BQlVcSRXeDQLHNYcTTSyyRkuz
gHaxz0ZL0qi26lfDBZHZe/bHhijg0jIGoEMaYpP7ZuC31H5Db8kbqnVdJysc
7X12NuHkZjAIV0KEAp+nkwcnmPIWahjhFqGBkUt6PB9gKT3iCO+pU6gZoKJ/
68BMiKrarg1HYmmSCE/7v6egIPy7+jAwY4EHyCdRVTEKFe/0rtNJXxpw4SKT
kVURzldjt3yw/Wja/LlEdsZxRsOcral5sDAX51cREV+O51tmWaxS1fi/c+or
Lo8PGar6hTDsczYFcl1N0HBpv7KaoEZSKJJokXM+loWEryARrzZDU4JjyyHm
HmC8eHikIWiS+h9rch4S4kiVPtFYy3O0XiX/3Nh3ASFwURjTzz8VIuuzc57r
qUM51te9GK3bm16I5xXIeI0DwIi+uyhNtcXHpsYB/zlXCf+Rf7i0RSw5Vppi
r39c4ppap3uz1lLRm7JKc7KPkVWcN7QLbXgf8J0FEPNfEZboD/H4QVC6sahQ
C6+xgocTn4cqiefc3dAv3PrxxrszP1Ahx7MdUzDUF29gpA4Dl1vYK2rJ2WE8
cLDRT6dze7VOZdSO4WdsIr6xxf0SeNJOMcsam4+ooYTOtVC8RUEf47DE0j19
EV7hVxgk8zKZDfGwrgoxFnnIVL7d9HfErFQ1Cv5Xk4O/T7UdSvWpFzRV5v3W
GnuAliioUt5U4bda1mkExxmGpjXNmcHWLz9stkj1KRfVZawL7II/v9BdzLFV
OeWOLgGKJYKFkwEraJqpb7E9ISSM5duZ6TGgpJCQmlJCpOJUpAB6jScRpi9z
FFSUNNoUDbs2HPGHSs0T1FRMEGQ/0+9tWuwqGsa9r7nO5SZo4cNA/4Cu/m4H
UZN1klwHOu6IAmX9q5PRo+tCPRd+spEgWd5nhxmkrJz7Ogj7LGgoe7XYpeOn
DAdZ1xpqG1XOx3vDABOsR7KNNllsPMpFTluG2i3KtzvL6u3JmoujIbxutkfs
peyeOyOTlb2kt2YbXmFd1QET9hoRc+6Cw3nDZAK1bD+Fnyx3ir7sS/hflW5P
48zBgpMqNCXl4NC1zx3u1mq8bwhENo/MFumRhGGkecNAFL5POEaWdlEHoumt
tBIW7n6OMSw+ky8OebQyCYW9fKwvnAUokkOkAV9ipRu/PNuUFqhBt2xYAomv
uDLeN63pB7hSyDkIUsUNXWenQ322JrGWINY68Wwq53Q1+7rbC3zR/xbOR7ZN
WD0bW3pw+uDsNLeuLWTdEuztgaitXYW2mXEScwdzpoTCCTFw8Fxcfr3BrY/G
Ayold33CBZWUXwtdTpTLR36w5D+CysR6YGr/AUvsGzAyR0F84fFxnMgxWgdZ
H7qxyLvLwVzvxKR8Ag92mc7wmUwv7huC351OqL+lW7+Tg/kA2rtVolm4wyGi
pbJBME9btg6cQte0jd/VnuVuaYVECFSLLjt8pdUgwelS8FtyyYBi45XK+Eeo
iRXKgfLIVKbWFgUI573HbCm3nkBpp8oyu/BwCROPN75BPjj+8jehIU9HftHo
M/cvFGjvkYVqCIHBCsCLIuuxFpT4jVTp2hk6V1Wcbib3qQEA0o06mQxUsoqh
ux+EkE5VyuI8Mxu2qVqqDGwuUiGw0jdp/AqZ9bVPkZS3EdYQxoxVaJMHIRxI
xJ40rJx9xl6TZSdjq30dLnfgJ/m2a/g9Z/rxu2NKpHoFXBVC+wHI6lNekR3R
n6HdLpImZL/PxxSIG0tTgVJv628kSC5MStxYGYwx0vxbNODaPIk/Ihg6q24l
BIBX/y/hr9v6sy1GvternLKVW81fqyzXb2dCT1xWhGXdof9gZTM/LyV3hUNQ
E0H/GRezYvfRBphBsBZtQdYURI7R4dL0lSIOQ1AFLNYvUX0S6b/f5wM5zPyo
t7nob9Sc+/4K9etUMjwQ0qSd8sZ9u9qnK8bHQPxZHMbFYNRgiTI/am7YSjA9
Fsd9zvA7A3lkzj1LMTsuyitY9Fgp2n8I+pnPpVXrJGD/2JlCMabup3Y6FaIA
QTdLYZissNZSNyRxpwHqAbFJRus7x4lRQdHS5tDpN8kKU+6dTwrxgdEdoW1h
ju8KpRwwZMDrSjJUaJk/i0TGTGD6UOGRfwXS69eVKTa0Xt0nagg1FXZprD0e
jF9PZbanTp9GyQsEZv2bctikHBUIWVw6Nf/V9jy/H/j81NOecfGYRupTkGvU
Pxjvkw92w4gqp72JQ+d51SCrW8Syvirlgj0AgcSIzoLAbQ0MaFoE3AZXLUhz
/MCvMnuJ4bNw+UJy8CqnNib/fDAZovywaqibx+pujOHKFirM8W5MsPthBZt8
0bXsjplg2ZPpxWZ26e2lR55vQCowt0n0qBQBt4Zz/HDsp0X5PlMTwPQs5+OR
KVB4MBIpsdiUUnQ8yZlODgnqCI+XZqcxjzLWb6QMbKN6VoIaVMIDkdj0uEZ4
aPMxEjENTHR9YGR3mFhbIQiPMN5G1xt9Wai8qRucXzMumMxZDM5NeOOCgOTx
abY8trNiU611Zq1u0rKbTChGE6HRflrpwFFj6GpVjLAOlT2R1RDvNs3Ebhr7
UppSDLcieFvlM5BI6ntwep+OfoBeUZ9+wRvhSOcRtaA1XHp2fprQFTKr3kJ5
atdei9Jf+ziC3SVN+Zj+07CH3jMUtgZ0UyDSbngfMOwtxoSTMywEZQBVNL1l
y7/ka/Cte1LbzLerUO4rz3cEdn5QeTheEE1dV/iLLSJXeu6kHD9a4xGcnNAo
TdQ292VDO+BhuyZEGtPtfrzKQUbL9HzRZZR+Z5Re61cJqmx5NMAl0KHx2WV3
MFo7NYSoyxfEOez5ANfm80XoE5L8e0eS9YRbEQnHKZmdHmvZShgOOsp8JG2f
HUcQSGR6WwfE0ME/0Yx3c8SvqIwpvt0jP66JZDKO2Q57d4LxbZHdJxWBqd2A
LZEm+l88nPj1+p7SkUE5xT9yXv5FN8nWipc4ZMWD1GolysV/jHiss5mLqatn
ZBigojSUCBW817OMkeaQa/vjlQ1DN2AxcpTKLV+0DcqgXcnWNUY6TFZE9HRj
ZawmoYdek6gasYFWC9PgEiq+xAb3jvahqjAnyPQ8qPH1uCe1AkZg+7LePjL+
CoCzJCagLrrpkxOlCb6v5aaIWZ3A5/t+HvhGtyQ6ksBxgz/e4qYG4B0Gj+iI
b4oTD5VhDA7D7DsnbCdsRyj8bq5/pz7uH93XjroiTnXX+FilPtcZO52TKwdL
K672AoXqT+5O3zExmTnWrY1PSTbEC+zY1K7OghEdR0PASu4GpO3pK4XKOdew
/wyg5skDI51mWDY9SMjhMtKjanaJYi1EIoX2TIWOcDYg9d8Zz20p/dUn9d4o
XO9Wz+kkjLGk9n5QYxBSPrf24JsEoTDmZP3WqaKEKDVSVQdBUx9GjzIoMWvA
JbKDGYdYtSqnGB5HYGVUZ0siFXMN93ZUW9PWy+tVjNgcLdkxlPSImLbtqS+n
0tj0+8JKWKDyZRcyX/mGOcu2IiL2pB1WTawb7/Tfks1J88tF6bQQvQMNZtmU
QvHuYaU7YM6uZmUQnviBZZ/4gDZQvZ/tpF79M+Xs97qtXKV0qqLghZGAGEK2
jyVjNVz5XXm4a2/Vex4MfE4gM3Vkl3bj7yTXLO6i7VeLPA6v3lhBRpbGEwfC
zvsp4Wf8dUlaewQyK32V0IpMS7w00FMzjNcf4svOT3FVqCtpZdbqq5pZ2Bo9
uKTHHL+lYlWU9924ifOLRzdRxT4k5yOROIk1HewlFHlEXgEKq9utDaF/kH80
JaAOlCNJwnGokpkZaSg8oEu8b3vR6CQXMsEhHC+AAMg6mM/9YUR4lDGo9d9W
si16QPjxMat9KZKubrPCkzhA2mQ615yvH1SDi92NUHLnBnz83qi/80pbB13W
S7k+upwnWsLwV/fuelc2ix5WUBNol+gtiZlHz39J5CoDP3r4hGme1+Batylf
UlrZGCKSMM4r1mVkWkc0lfmhAxjkaiy3R6Sty9I2AQWI0JSyJF9XQ2CZvq5p
MxnaDE4L4b9uLIss6itPKFZ1z440uTfRgJf+g2IXOpmRyC2Z5cSXCOlxmpn/
G0DNYSn9tEiu24jsBDJ0KldKUO3o1/tSbCyqEQcY2G6hrBhn5aVwU28WZhyW
AW2f84D4yS9NLfKCWsD4+ivyv+v5zRzMZ7k9Vee97QVqANwEjWQlLGVwBJHH
CUPe0buy8X2/zVrBEzJtaUgl+ajgHjA8luOCAbw0QeEtlaPA0TbVNI4yOmN2
hyM8U4Zep+QOEHdn57DbsVJeWqyAwFdyeRHzIrN8IS7+FOLF+XOKg5QGNSQk
FT3lyRX9Yr4TQu70vcppcLmlAkKEi1owxGgZ4Hew6tcSOj3nHYJ8HSPkCT6t
t/psac0QjPnz503P5fwDhOhtFxANWf+06u832f7RRcfIi4xC+WEcDNvPudAi
HXvgWB1ZXVQ5n2w1TIt66Z8dBAJoUrDripA1w906qTbNIwvRApMPmlmoGXAJ
ePpNH9CxtV3GAVhOdcfcO0CwRfNfGXP7YCdBbIiRlzG3M7bBfXFM64b+T6I+
Srd2v5LXVeX9ro89+wEB/hO7koSZmQfYelZK3GbXJp+0L1woRG93VOuozQiF
ue+AfAvqz44r0QWRE3GHfQ5gN+/MA0k1PQ92mDcU6ay1O2BhLJKlqwk+/y5C
N+6f3i5mpEm7q/n1xixy02Fx/DjcVRYZo0ImFRT2sFZgdikSb2aaDKf1k4eT
8Xvq2Uv/ZAhAZjiBtxWzbfK0YnWO9kDodR/7U85FRvxy/DdfXv4u4WtUmF/U
QJ9xb2uVMLzBM1BWE8ROVAxzwVcjqsf7fSPdnTgFjD+l5tH4D5q8MlRPhO5m
C68QgOdyS62mPiOkQkI5l0V8+ztWhu1P1EQRdHWK+YQj9idLhstU+WouxmDn
/EAhKhg3Whx3q9GWBRbzyKcTsSium3Ka5qHtF438/eR48t+FkY4uHuc9FA0C
51zlbF3EQ3ivo104OUE8jdGrT3YUMu1oO73IlDEVTUp4LB4vUYfnrRvS4mv5
6KNrnlcXOX0a9flAMziIeGupy6RWoW5LNYC3Qb7ybhbrWbVRgEzodgUqZXxJ
BCCd1HfLb2ef0vemPcTnhEOFFz2Uuz2pCuovnz7oARG6NGvSl/G1nb2/GhJq
5v3BaE3JPuEicbbXy3S3+NBLiFZxh3bDEbpbq1qPPw1EUnqteFdx0XMhrDvn
0ZSWReesoKwWKaAniUkCjIidRzjFg/cbo6IaiDYVQFDz85I241h+whGh3XF6
2R1C5wlM7hNTflz1O6sfQIl7XiHVCPAZhJ3u9ycL/LZ8qfhvcicpQwZ9xV7P
3IoFlPM7T/VcZzgpEhVrwgtrY27n0rqCtx27s5CuIfHLZK4o4cBhOdgTLB80
tnqENpHiokFDVIkNOMKctAmD7s29a8+35Z2CDU4Z/SZ3h04aidghiNicIm9d
OSFC8AdtRibgtnFlq7714o7SXN0FzpY+YThU0PY+ttSpgpACy+1q9990wvtE
V/iM6D7zBNjjncGokFWbfYGGkv4sV5G30yvQ1QzV1KQZ6bsZeJCijiPQN89e
5Mtxj/YsbghHpKEX+b+NxUNsP3iFVKQ+XcAY3osW3horNGUNdVxdPyLslVUj
+p3EcZqCRaPWbnVBLPmraCq2MgDKsWLnPNaIB73Sx3xzaosFHt/EBuT9vb0L
xZA8PBgirI59h0827TbnXuw5EW1+YiKIep4WaaHNkL4QPzIqknxehjoQNc7e
w/KHtCNApSXq5akyEo3xuFRh4oRQEUXHHhiz8EF5Ru1cdtVpe7bi27Blsmv8
NbMAtyj2S4vIz8qvCqDtK7U0GvjQgX9K0/lm1EB6plsPi+XXBpuPSZOvxWYC
6YtNUD9zrJ7wfuHcy6tWxjQnwrtAIN163wzLAhEOTOuyPp3DM2T1nh8mIKOk
2W2OwNHgrjzkTWOnyx+RG/pcxG31+/V9XS1Jek2/ztbNk6RtSr/w6DHKv20N
2ld74SfD4WTEMrpAXlKdAcvc2hp6nwUtOBX7xLQ9HT8RSInFgEzGKMiB72xS
Z9jTGUmdOlcgyCxptRJdKb8emJibot76fmPP32dInVNJCSN4smUPk860A6o4
lT25DDxCZrT7xqKx6LVaMiuKB4MRU9Hy1B5ibfZm80uFlH2oXkAMGPXPyyA9
zUiqt/xqJ8EB0hwO3drQQFHIDHrQRUKuaRXuIZ4PQOKchMIH9t/jSDT0TFsI
RWUroxsygTaxkVxDgG5r2kASjnQvr7PcXgVHRHOfUGuhQjNZX+H2P1yanG4t
ZXHh+r1VDMAV4CHeyMO7imeUy3ka75TXm5uppl2OrQqclTy5GHniv+95JxX0
AogFkTEpEEShvCafjzKIU47VA5qzY+cxEHDiRKXDacE9W3CCyjvfyRgutPO7
3P8ZLzPCe0gCCQ/tiLSXHyToJ0eSv0KsbAj/ing3N+wbUKSrIUB4S2TeqKEj
tzkaOiaIBhGf/VS1StfzTPPSiT3jl8QRoU450YHjrMo7sa/XAIQ+bMM1l+0B
P+kSz0dFQJ67G+3GW8B1dPkByR3xxx+5YSOdUcCDbHeF0rDaObV0axRBvHYg
Ptn7n6eX7KSk41dHnDX9RT0peIAftf78T356tv4NjQAb2FcRds+n9vMHwulU
C19mz81I6S/w7rPSS+ls5MXHGKzs9oz/iPjZs7vrAftv/VAVPFyy31yDnYo6
R26LKsvWFKh2mJRrQrmB87GL12tmEAgWN2GjqX8n0zBUEXnSP2KKruzCsK4Z
Oi9v7Qd5zY+DXkQu/6kJWv8CtmsDGvnZDoHWdPXaDf2Ri6Msn79+hjShQ/5p
HlG9ePIe6x9JEa8DLhIUERbi4C4bdaQmuQ2g670E9OBY4SR+k6zaeEh1Go7q
EPUCkWACkRomIeWNEb8KdUBX3a2XpfymtlVQHzQZEc5DKWJYdR/GiwocqLAx
ueGuWAL7Lt1mMJz9Qp2yu8FVm4L0nnEJWUq7Li9ADRE0JSg7wy7IhykevouU
ARsx88Ku3XeTPASwuUsGEowTO9NZw2uorUxYtW30W9lpPZFX1Ij9dIrqY1zb
pKZB2njOlU/iwoedU9BgNOxMAnD5W4iF5KxGQmN2ix3OZgV9iccE400U5QwH
Rb1i3Kv6NlhodqwIYBnPRHXWUr1xomCbhefWfcU2o63uXVna0WB7w8SlMxvh
5AHxe+pw3/6xNL+1NS4V+Lus4rJ8j4mMIiHM3Q482Bxo10VGQoEVpz/hX9lc
FZokcSYiSWG5aFA05TfUJwHzsSdzgPrqFDqqWGmvzqN9+T0GMlTdiA3/sqUo
TsLZTS2/VXN5uCg7bX5LvuJqTgA/8nnXQ5PzUP0ggkRfAXKFjnlUB3B4pHKO
CNOYovtFP1UP0lRCizxBPcpsqsgeevcHC0EKzeNVH9fkKVH52wN6QPu3QS86
6DS18rH39K8VCkTv8XhAGxb3Ds49DAshYcAuvr0r2ksqoFU9NOafHxobP4+H
PASx5IOfkWS7ioBgTZ14LHgIIjDUmNYrlmMuWY1ie75LzKrXaIx9HhQ/xCYy
mHO160fm3i9sgKIaYZrytsweKyBJVtQ04jC7EJGeUwho6QRwu6/dA3/15oP9
k8CoAtBiUNEMpfp6NfW32iyhNryJQNO9EsZcZQEE2XBKLsFHUsGzwXzu8+NH
zaLTVHIe1UsGQixOWj9WhEnI4tslUAtyazqXVT/j/jIi5ln5IzNgG/Uk0PoO
fWf7eDNPZ053ZQ2n6trdCVJ9GK8I7i+k+glOPQ8KSoNubcG/CfoG6DzwjPqV
7+e7nOcTZx6rou/LS3K5oxE9NAKrC08Y1SGMF7jf4fAUTCb9pZc2AoQWC550
VAgX/83t+iyJT0W88oGVaD40wGyUDDJ1VuDusgG4RCTSoztzeA0ICRsyn4BZ
OX2IXVshrNcNAgNWpByN05yaxA2s0vIDfEaRY2oEU7zLzL+QCyRLzNzYgPvV
lQyibdr6G/iRd5Fty1xibKSRbs4iz57kc0e1ZSb5ecxwVlPU9ddkJFsMHN8S
HVi08QuFsqC46wIZZZ/ckcV5rrrqlxD2HOHrnUWTPUzzjt4Z7YESObg57jfT
BKdNTtfeCwP5ghHAKE7RZZ59HiuPzCDjFkRFWDDWOzdRqGVsKxuUext6U2Zk
4SGlfhh4OftibGcOoJhwel6yOhtEBKDr9KcRGPpwH18Q4cyWsZk6z3i9JNoY
vehYcuPZiOx7eVa8GQM1qSaUEb8ExdoCWC2cFuys2frBxqTfauPd0V4WCnHP
aFdEI9hMNyrC2urI61FiTjpePkRYkLysAQDQNiKPQ9B+V+GL1xCry8aeDWZ2
8QACABdifvUt1m32O6S2ccVvMLXqsoxD5xO5M7KwoTsljC/CUxsKDbVe8pK2
dJAngvj7+86fL4AIM1KPBlVcuua4S3DMHdhDV3aTknIKgkp5rQWGnTc3/VA3
nDEO32cwGQ0DO6z1w8NVkeT31eH2Mu1bMmOyey/e+xhY6dAO+eVxRmWIGuR7
rWB/gpvfdiVVgoe3ZUzHYkIDhZ7ca6B3nzRmIoA8wzAg6C9DevAOXtsY4yzQ
nPmw1Mdy9UYX5lNNQQx4SMWhudbVnE1UxV0eHn6BZ9sZRekrYFL5jR3G8ddp
1+RZAIWD5aqoJ8O0pqKrgLLn0O6L4y1SxFo7DLFFVkfNu1nVSXtitpXIwnR3
npxR+CXLGPfahW2OsXhRYc+gShVH+Gaoaspo4RXk4snuUszTjMFQd/MfwfB3
pPq3DmXPDNM/ciVkSQfmtItGldGIf5y3AYCbYyeuQMTsPVoUQIuJx5RXQsDj
JazhpROz5SvDM6F8p2tna+3tv1C34PHpha0jmy0cWaDlZh9eAx8zciJDkDqR
ppo4jeAqhFO5/4FUX37+foWDSKEjqguOTM5dsoGTKYYTSvRT/neUysHXJpW6
sFHr48/eWdSao9TnzJGca6QbZh10Kcc9jcwtM6McoKI8giuOP0sk72wG6i3U
0KS5VhymLBrObc1lIUVhqu32tmH5oUtIVvsYiMdU83M61yEqJvatTqFHhvQn
vzuyiVyVgvHO9vKXESYS4JAZ1U3crb2SeOm90GNMmgtN3Hivef82NyCQ43oU
JtxILVc8YTtP8Hu6JUsQR2qgdMqbZg01oGYJa8HHhivc032sTxVovG2S+VV6
rpKNa4rBPE0p7TBqGfvOaWOdGuZiUz294w1vJxsJK3wXBwuukPFNcsolOguz
514k1jvvmNc4xO7JcxI3OYFBJptBgdl1pAa+NIqKZizlbCcn3GGJnrIvqjPo
wmtsivcIblqgBswIjJkRG7ncE+SlP7sN1vEG97GwBvPcG161suJMcFFkh8FK
d+fCI/OxKAvYfl4+xpPyh9DH5IEiiSuVwkgw1J4wpXPsFrjwuMpbvLfbnrpK
Hq+n1RxCPxrUfBqtlFqV8QJmfTyHqMN4TwRMibhmQC81Dii4B/89MuCYGK1F
k8bN/gsiGlU9oU1R/XAYV0rIxlVdBa6qazEKymlP5PVMqZADu4TupTg6ARv2
3oDTtphPsLwVBWHq9OqoA8VWFTpZiIVy5pImpCJzsw/x27Bb0ltu+0vYtEnq
nOsufFAXSCqDmRvTwYh00rRS0LSMLYE72uX4Emz+3Z0DN3N0DPs5gcb8vejw
/Oa8zipkjEECi5q/9tbrOqDRTVy0imi2ho4FJ/oM//hjQjZTqsN2XSQqeynN
1lvhltbyqdXo7towU5xo4ETi6WSbh3q+zPbFr8WkEPXIYlLdKfWEWo4w3ikt
1q3jLQ826362tYhFXYE6ri8gDz2sQ1/ObVAHzeVSC3gKc829HeHh6+pwV6wd
G1Bbj2poUh0GHBygb3cq8QYK9yJOrpM/9I+9071wNd9VhmSuRY9UmLJxIcGP
id3NJvIvWQqtGjqs/ioQbB3N+MJlOiZKRtjz2mCL5V3C1/TYL7d0xrGurPyd
CSjlFof5uOs+lekfv1Y7bxq9l22XqZI/UZU0eByL9tgFFglwCmI/bRj3ktD3
qvXl1ApgQeU+4ywkskEOR9fNldh2Onx6B/q9R0PEUDl9Cq0UmPvyL+BbfKDE
1lAvN/cnc9ZCaXqQqLd4ir3irWrbvYH+nQglxdMhg1XCPBmJEHmGdu1LTR/6
2WmzipWYcSGa2TU73FbJuRs5Ey6RqGIP0p7GArGlBVNbR3YvaLD2A2xD9wXD
2B0ANq44kPGncRjgyfshk0Vt0pDhQysEhWb3rTEoNB0ctk+agjL7kkyB/lXb
y69Ox7T6/DouhgIiLk/WAuPVVCaS1iTcqk5ujnsqTGBmVyt1Sc6jdJYlZhb2
WyL89fyW4u5YpfMp6ifCRs8eGcdQNxHWQnoGcXnCQzHtkIUu1XJ151GwdmPm
l5008iwgi8JEStqiOZtQ1FnRr8WOs0v+dUlG+gStD/BnXl+LfLEGJDH8VbNL
qin6puOLejkIuD4GxlNwPJwX0Z+a0F7snOJpoT+xpB88GiJM9+dUURm+IvH1
Y2hHmgYgTICGf95L2DQIQ4c8MY23Q2dj37LPrLcwTyFptmzFccLj67cs5ysW
WsIvv6ZidszBTZEW+5lUo86QMPLjBWeFZqY21TR9T9IOO3puutNOcSxPlysC
kHRfYUxDGAT6UOuQE1478PUZ4Rnc9Ulz3rntAreEUnKq9sQ6vnErNkGlcIwX
71zJu+TqUhl5NkTVPrffxOF7IaEmOk2YlYriihC3Rpzs49wMFh4RRyNlchWM
OLHJY6U6Tqkw3toK47RWduAxdnZvwh/aEF5jshR+v3oIl9YEY8T/1h+rM261
vpYNnorPr/QVgwp5fWO0ujXniSdDR/513on3g8D+JGdl2UPyBlykjghuwPD/
mVBYmavNuETS9fwTNqrrO2otF/leiQbQw6ieDd04dtZb44vukbk55CpZUk8x
M0n/Gpv6RcdB7Onr7xr5t9s87HqRQ2MoM6s/EtUZADquJr+syxJI4z3J28zU
aZDA/wmfDn3Xn39y3rXgeuT6AGZa0p767UuDpeXoy43AmOQg/8sGvGq0CS6X
uJXsqoezwDHN4g2G4hqlMJnsW7B32gPV8utQ2wCjgu7eguyIMjwrQtvJB07H
X85nLVuejmiIwk+OM/323pC6NBB//VImNJFGuhHqPUiUg0jXtLNuOREA7REB
VSZMO7hk3OiuQBz0c4RruX780oLBw7EbMrVAp5aXwMTGdijDIQTCemiEKj0H
T1Cp8N4ISjVZTvOewZ3zAM91SGv1T5y2IIbxsRtfH0igHYRgv0U6XwucB9jF
0sVHYlV6VbaqdimuW80kTFSJGwGPNhBB/LCb4p7/zUG1uSXn7t0CSjO8GiGU
f61bpYiy1wL4qOGXsNFXEzTHgzKnUnAua9cDKoM/FgKLEKbSAVbHpU2wr3w5
lpeoOo/O0d26i2xwPp8jFL8EOCFRircb7LJxEAy472YyGIRU/j7vUONyhVhJ
X3ZD5zHiiLGynaCFMjQin/GurWCyMzmJwrKCQltARiD9JkzVkJ3o/sC+dTfl
iY28dPhk7sXn0vmvjYIeSD3EttU6VduR4pEs5i+GBicvc0JJsLQwCntQMv1s
hHVb0zEnRffAp1QWDDRJz3uHnBojoSEwAMHq7aUY4OFiwq3W9GKiBkkY9pa3
XyUdw6MIJZtbmRpoeAzLdYctJihCWJFpnrE2IDDO3yF+vWLGD6dCZOmtJF77
LGGmHJcdlQKXbxHGR09XwJBxCEgp0bcHWOhtICo3TihwN6ldrGswCShS6VU+
QeQKORdrKhgQIeQhsW8C8DxMZJmVPOEf2p1XBwuOhMa31T5EDiw3QrHVz0ER
8YvhmR1DyRntK2A7MAg6+L1mxz0rgFCNRo9ACf2qVKkK7bNpyJhMUHxrbogy
Pp1N0UWG4wTzoMR5ceV69nSfbtcggVvhIefhRwlscm8+/xYWB7XtKB9dmX4s
BniSpszeyoq4ZUJMz4YgehNEZb3IyEwo6kgsKwUEtys0pfM/GMLeAhn4w3hl
U7rgpfMqc86GECAn6mbAIUZl1Jy4jSQzKNeaxYIlaxKhe/RIp21aVGThWmiY
GNOU7P9OCh5qGmRHZB3HRVg91tDzCjhJjZV5jpIm+pmOrzlbKtI+1WNYNpzj
9NGqP3IncmCSWQEAQetAuj2q+JRMFlzVDuE+PfECi6jBXy0oyNW5dJIDaLKo
hQuc8xswRMdhHbm1+7Ai2e/Ixbd/xP3V8BvkFP5io5lukHqo0EUyBrFaTmJd
ayRwJl89PLbHFSnMkOL+sNa/YrVyUROQ+NR+A0YFwysFw+RVuL+hZrSjcfi1
fkN70c5HeOpOZxv+2l35mELI7F/WkWJFsQqC4gY/zLbNw8i3eCugzGzDIxvd
+PvC58+uHEePDofcMJAUjemKkZDnCRlePMm4QmLw9/sCwrvdRl9RcZLbC3uq
DIG6A+JvW08xWKDevEeafNQIKriixFQOzY0Img75QYj6KXbxIejdgShhmda4
uCCvG6Zd3SfOwThMzCRjPVgXzHGhXodFKku7P2IIFTqUNG45kF5TXvcIJl4E
T+qH/lsrV9OZF4F1Imm0ZdOh+VzlK8cAqplRqgdZL68E6CSabnk4oXCLBgiP
NXdmHlQA8Qo3nXRx9M03+qcgTgir6V5lt1glf49/l5s2yeUtDwDTJCY1LpSj
UQiebaKGBZtg7ObM73WIeUoay3/ezDa/ghOc+mlTQi0u58DLf/RXRQ9FCM7H
1f/zXOez9CJI/npE3fgDczXfjKJRZOrjZY6yMGt/5rhXc4S9TUSjG1GRsYTB
6mDJX1pmVkMBPjFjB7k2/JlNsZ+JJLVR4NHVJE6YxSx8ugLZyxz0Vd4EO8uu
CBrGC9ySI0qsQ1TRw0Tt+hjIqui4CYUnA6VhDuB6fWPOVK/O7MTe7YwBKi38
sDzwQVqP3uhNCOEfhXGngPE11kD1H56lRA3loMDeeOSmP4AqnYe4KH17LDMM
72/wmBQk2v5R8DHlVnYbmt7LOr2CEc6vJ25J0+jdlYqzVxxTAsa3amxBPY7n
GU2o01mjswXwXTDlQsQEKCPyfiq7q3232nys+KnKsdEOSgKUBMWch1tTznCi
a6mhct0LRIRznBeiFySrSU5WUJBCY5ziB/hiDa7sAKdBl/ZFUFlzZxsupnIB
sWc8GjPb3KkwNYy4yB29Hvx9EZJDjZNc1O3Jpy2omAexVScPabGzSdPZyaw0
XFqHqmIRqAliDwDpWF+QG1Grmt9gdY5IRJ2eJxaA/G8KPd5mUMLfoDhaimBX
AZ+Hcs7ByI/UHYD6v7f3yH78UELrHS6K5YhDNJBGH5cFZ34gjBcW2LcL28wK
Si/dV3453qwTQCrYCk98N6LdF1+GRciY95hMtz5KCaSxFnANq4A4ayGM3/Aq
G9NEwj/TWGwveOeKyU21t5sPPQPXApkdI+MgaNK5T/XD+OW/vsnhpFA6aNMe
GQd8zSAbMg1CF2uxNqU1DCnH0Q8kpGlKvVr/IWHFQirP3awCS9NLpaJHjlEJ
eyzRfM581xWF2WuUvNJffh1ajWggtAqYyqND3dQX6GVF8iW41xgC8j89xpNP
qkTdCiVtRFSXI6tu7Ak1RSuVTiFixXvt4nFmqTHQ0NdYVkHOZnRgP5L1qU62
k/CqnNXIE3hdRYAHkRxBGvPAI5jT3smy9Ps52vh6XPi8qfrmdS3HEd+q6dOq
2Y/HRWR6fjCKP+jsb1HR8UtfQhDMYpDjUHNlS4VCLGPMJhiHGUhtWIjrjpw3
wDKO6z38uD8Zm5hd5pdhBpGrTycGGunUma/CiPtWKAR89866AOvAyklf1Nzw
CXVks6SNB8FEBT1QsXzgSvdLxli5vwL1WA3P0UOqagPhXDwRUzLpaO0t+Tvi
YWwGSRAgSKGu9xHBlAUV6F/jxRjp5/qvNtPovGvqIp30MhtgUQ9xNX5w5cZk
Eex/TqwQMUorvVqpECNCGsWVCmNYzl7CYWaxEO8ZhQ2HxPNGwhop1XWXXMt/
UpviDuW4cX+ozmT48Z/s4xvZmdaP9fxcuLIsMARj+uU4di381Jzn3Ka8lyh2
C2oHXj0fmi9L/ybxmnbXwcKKVUglS/gB+GQVOj8VEkm4gmDriwO0LJlmtp2T
H5iVofKfFMVfMvyYXjaaSmTEQVVVKwQs6SuBucgVxeVOqMZZ5oZIm9UPlume
SpGlIjefoo0e5iyzntWzieTvbqJntxdBw683TBQ6O/zgyufhQeKUw0rVjQQX
Mg9VDekXG4+5bcPj7wZFsRRGghKD9dEP2wjCuRNViWi0aZQXr7rclqbD6eWy
OqjIx8fowvuFbNRQF9w766gqgW6+8dMgCmRnHJ2bVDttKzsOCKbbz+HUDI84
LZdwW6M/La6+dLQuszSPMMCV0uG5tzq6MZ5ekwwcRQYFNhkeVZ/xDna1TuP6
NDK7O3NxuLF/l0IPGmQUeSDM1FMmlVCjeN2oCphSA1BZ9y2wcJEbiOGL1aEk
7eaJB+ISXgab0kjfWu4UlB6MotzD7SWEHfFGFkMFmjXwVWbqyq7Ts7dUKQ4V
lhYRKLnYLjlTHLY2qj0OcmbDhPeodd3x9HN9KumFA6YWM/1g9CsYUUYb95Gx
3FjnxOy85oOlKsd0a4VVADlviriL+3omrmonLx+AwBaZI6PqrBhbRyCoFF/Z
N07SG3MzWz7wQWnd4+QQystQOKa0ut8oy5iBWC4zQQfSeCbgIAox84QHAbra
XED/Cll6CLok5lzxJuNFHO5M1ERZZ7xeTcW5QZgRhTsoaB2Ex6snqhILU7QF
R3j8q6C7hm7GeW6S6dYM37wlA2IHRSVcPQwjh5b2FBmcfibwZ2bmTVAFrGSy
bXWA5cWzKonnMbDsumAPpWJmuzANPYVRVUhykSFSBA10FyPF+Bjg+0Dp62yI
8FVMRE7uBxiMlhifE2Fk4vg1liPUc7JgScrsfW2G3I73JADcuWCNSt3/GWdW
Q+7IWVjN5S62GClwfpweZugIT+b9dmxniMA7PkSWTDNUpQ5uCykZuGWwAMD+
9Ts3io38vl4Oz0J87bbjb/5nKZqtSgaCbnRLOjAglS/IKQt69hd4QEpRFzlk
0Cg+qLm3cVYWBTenHXMPShEg0ePPh675+aeIfT1uyvRqvtyvkgpq6cULBJKY
Y8sBDZD/aRLZPCTx8+9YHDBV39+aATMPut1MLPXBno5ARkIyIEDrz1YM9o4m
rUbJlWMEhCtwji9MgXYBWUmD1JQlO10T6dWr/fiWw1LmQiiBbzjkvrPNT4bd
2lQQp8SF8rwGzvRlxrZ2fb7Jaus5nQPOvyiNiK6BpbkX/j6gg1eJVl7uYvc0
lXM7BXtI8ND6IpPTIqnXSCqAJ0ztCtRwEIcvCTz7yjDlUUFuczeq8G/y5uws
h5EBcKoKZF1RZ07o7FRpEPClcK7YD1YaMsihtonp9WUA//iVjYkE3224N/AK
e3vN31G3LgKv1u5K+J/qIYnx43Pkn6uhX+c/CWs9cO9WqgYd8S45iedXAORR
VVaglxPY3BROtEAxKMk4i4yDVFsG/mjRP+ApXFQeR0XSu+vYWzUszJqI2c+i
ch9uQqlW1HrcUZf2d2XEzriy6P1BTX/7Sa+YlCtmw83gsQGhOSssgR7Qg0vN
QGeEt2xD1GP+rcRKIdcbgRFLGKPLOpgD3ga3TwEpOgjuKwuvI8F8pnDuCFwo
3YSF/3PbgV2wWkfMgNguvBCQQ3dzRB615QphSEsSA7QsaD8yIwHzQYAb8LsT
3dRk3UH8xHE6IRmstjifo8yZ1JL/wZb++qIDu8QjnnwHqawsfpKK5YtQMgbS
J3rCI5FOP783WvlR4QIFy569kOR8i/BP+5WQxxFhbkFuS4on7xKYGRWX6HlZ
iQnisxwvWrgPRiyLxIX8eWfkm25hjEl6zccm3eKSIfT01NPvdAWHabvqYHLV
JT97xJlVgx5RQoVFNhRV+xdZxe6ZuKo9O3lLCu9GzcZSr58ailwNRaaqrp8W
bBbm7zE8plikeyYegousYoaMDJOA4nu3aZaXzXopXk0lphxSHyIttO9V1ady
ZSggXy51mX1husDJ92IzNA8hsvcYO8t4bi5I2ITNiY+ecV57GGzJhlHVLPwW
1/qQTsCwhOVWH3jSTZK+SomZcGjatd8H0QO1N0K202sexrNCTafGiWuq9jUT
wR7AU7hT+GyTOq3A44uZfLe59tAfJmNb3ybzBeIUEJV78kgYPL8mhnFlDHfw
MEhJQu0hpVbAR6MytEZBgwDYhDXXRLIEhYD7CSrtDLiZXb9UuMB08W8kfv9a
EVrnlZx1NOWCtSorJxq1qeG94dpuG1T2b39uefJguz8Qfa/Tb7MatmD/apKR
RsZ21lYryV5cYQQE3Gf7HHjRU3OsHH+n/hyp2U7DIS4tQCFVOGDR7HYhTBHn
rZiFNb6HHz/kPfdG80US1miCra2xScsftZze4uJp2qLY3YRdYOcT9r43x58b
NQQagkEPPmJgdgsrrbCLdqFQfgwSsLLM00yu4mneRxI9WDsSgL9PWyGoTDMr
9bIaqA8jnIFT+9K8/ICpfjg5Hw0dZmcBdqMYlKD9umP5Ag4sWCOCkEyJQ4Js
ZaQnez12osiL1icEclr4fVgvpSkJbR2V13fb2T2RKupbZVRpf19OKv1nyMlZ
BNKnOFnJsH8izrfJW9ZTmYqy1bAeJl4av3+/QYrCaj1u8V6nxThbgWzGsjAt
6LBxXOnFgXmQqvqTdtXuMAMcldnOEteEwhl21EexMJ2XerY8XoZEsv/ERvu+
GtKeLWT3ab6JVxz5eeh0H/JTr7+/9T0ZhbD4ifW1ew5SsKBaSBAbdfSA6ZlN
b3ILTXAHldw+J8RUEWUcPMDVm4/iSHjM5cZhcj9J9ivmAGIu0185YzYnVONV
vkDutN04qSKi4Yw+JyvdAxeVINRDJ2j8bubzX3C++xKn/8I7ObWuWa/WCRKI
DYdzQlVSVbxppJ0PGriJk8bWNIvqJBYu1PR1Hqfzz5a0ziCLck61aaZfzg+s
6NZUOSetCMD/uTtT4H5NTGIWrpRyL1wbcfpDh9NCQXSXyTpwiV7r+dUzB3fl
pei/Nr/F2e0+Nuke6s91LODtUcxNGDz/wfeLBVvMRD4icj0NCT6W2+5ChvzR
+41PSz+bIibQoPirIk1nPPuKmbBfGaBPW5wRC0GLlpqLDpGoNLSvV/jUvImd
fOGlMWzTswp4g4N36fTGPMxWYlWxalHtyN6fafJ64mkhAR1WAAoQ+QIj5stQ
6E93qQ++RQp0RcvhNFif1sXk/QeERDBFiY3+gml5g5g+xFH6KfHcWAXZYB3e
wX9ISoeTaKX4E3UcFBQ5C+drdE0tDyi+Qy8KvEWyCb30bfjnl8zsxVVFqbfz
0PkF0IW4HMEkrJgpIwYQW954aYQYytGB7uOWsz8uV4ZAVnA5d+KBT8dfwtv/
kkATJFRylhGjxLwbA6PALyYcgf+ncvwHws6nRaLSjn5jQai7W1b+O4s2gfO2
uCTUl62DM08O13/m2UK9AEGWhW9VjqICQre/nmfwHs/DEYPY4NmzwZulodgs
TqXXH/ghilhByO1rnT7sbIyHr0HmwI3+u1cWvMisht1jw8s/EzSKEJoKjJvh
r9Au0GIHmlc40DRLUcuIfBdoMMD8RBS7NaMESIFRm6cm8xFk6HTWqO6tNd+M
Ah/3aknJL26ALRp/+LcJ5h2u4tkNVDuUDl5lqiLeRn8GVGOaTiGU4oB4/YsE
OrZ2TTe8kW4EOM7BC+8TG4L4OBRqY+tNVF8JG7SFJKsxTuSsukw6+h/Ntlh7
JLB3nLLTrDtRdxBAuP7sTWZWtoNQgRvp3t3gASavhIt44VTYCbsIozguzzP/
LqWuoL8lYeEzUsG0LYSBsoxHsE8hdpZ2nDh6lC/Kt6/CALM1NQkNs8vIv8/m
4aVlZ8PCpNG44nUL8SOiK71WhOE4RAp0YxW612PoRqgTDuOj4LHDlvlRFBVr
Ue0jLQrF08tzpfQ+1C24PilJiksgM2h6Z2BX3KL9TYe8Kg/l1ZjcP/WB2tyc
gZAo+16qwsZHkzqL26jdwna0pa7Bq1OqgfLF0MY0aiioZXbIRmjRVRLNy/CF
8SLz0WBY36ZllbbwRLwWcqtQcJYFCPXXgQPgBTjEEgaw9VbwJRJulOi5TSAe
ck218xR+v9ZOk7HM9pAncVnq753bW4yECRISYH4wyQt5i/wpG0/b8PKrJF9R
j56qk5g9Pa9Q9G+rD+GVLXH/1mdZFLYw1ceyDT93jr1wM6bluuhlI+TahPOk
BIjy7D8ChAPHZLY6FJb8QiPBljFvFVuobCZKYaUHV2upo1ZOji2D7u0mfu4G
sKGyBVuVazqKYQbkA/Dff37vFEg/PFROLvHuhHACyZT7jFSbe8eM1H3jrBFH
W+SGrNrZYcTnhM8GM1zQKhAyDGQvbLp9o0B24Sph2fSzP3gIhgDt4+uSqGHM
Mz/QuCmwVN18Au9SHc4rUhJGXOXZ/yK/iGlQL4NxuoLnO+3YWQwXFVQZvmNw
zFeWeGPyemwAsHrhXeIBiB/25JSgaPW4CO4+FAEUCziewSiDBZWDQ5JJ389x
9HVB5DXF2jvG6qaAk2sg3rIK4MXBjAKes8iCW5MloZT4LWu/VgnZWv9ylaxL
2AXp7m0yBNtTZYEWKpLkuYyJZgKx+BPonBS+HCLyrxD/9dzdPa7f4I7//s+w
8Rsf1ll4M8dF7DlrWee2ra2sO/yVePFNCDiN+yXI9FniBVvSYHOzMFOJerp4
ujcW+1hIZk9i3N1GINsIvBZHjwAdy7HBpySDau2CKTywnH7NJqfM/nxT+Epo
oPgUMFaHPfWTILOcF/Lf6YH7pZJSdOiP6bcSpzY0S79rkQqNkU5RVr30cSK7
FdeSIkTNcqEtOQSZnthxdQ28qB5H2CU3DtvOvEmkHuBxDq4KBVf3cl0qri7D
AB1xy6rvBe95P5Z8W+b63YcRqzoWYZgWt+WEtnHRVopt8o4NiOQPg9iIaRR0
syNrcqvEPkq1lJonawaZb9kPU6Hq2l4KNcC+WCAEYV16IzUXkzrMrkFsE6Rk
rGBBzPVJKqqIX4SWZdeXQFpjwuSIO5AxLdDdO6jZDOPxlKNOOSFyVLyLk3Ss
Y2esl4ymadqkVLy03Bda686yU0lkCOHpxnuWcUEwcCsOBlLNEsHK1o7wJtRa
gRAGV2ZZZ+yqELjGDuHiyjXbrVWdQkPUBj3iSidgGIQ+wn/3oF/4Ne3vrFQ9
OvUwggje456WSk4zG9KmZ6muPb3jweRrZXtzco2UMh7YfElbljK0vanm9c33
LXJc8AIp4BN3lydscFNFx9qC7Ahy7DBShMlTDr+FNnINDxOtW9sSIFTylf97
ODpBZ4snRcRVLWpW5bSXH275XKJkpundaWu31M7IzM0YG59Vx2f67KoGgOQZ
qFLjmLhDWIzTTmCXrb59ABR4jlUtbwubMkYIRWS85tI0xxc6IJGJqAu8a0VT
DiUEg5IeUsWN0cUaTAe14C3DzDUwRYe7ZyYdfKWHq3ENXQoueWTvsm6OQAyy
FXpZmYnm2Qn7rY0qz3UViurAOXnwLiT9YZHs/cam/lgs9ftj3IdJ3/ToVn0u
xRYVaQXfTK3GNEt9zam5T+cHIkPYjsAHun4NwOq9xJjw8fP1YW7ujUm1aS1x
iTxKsUwigNVqPhtMsJfRx6fFQUvVXRPQKAcCEgD7mYgP7Jz2y7+ha9oC30E8
+ArDDbFXXjISe5tj19jikN6clk9jF5oPFJZWSka/bI3zwvGbWhnmbPFZCsXJ
HGH0qJ/jVOW2n4w/BDHwLqeoRNSeU5p43tLWQs+lcSbFlNmE1mgzVPjg3Vr3
aKtwFYQiFncK2pNGXKeMPlaiC1HdK3OEwZPhdJYIMqT3b+b7BhOYWBw79O/B
jzDBRJvC+1S5uKzjbkekIKCoprMG5KRbf51omjGiOmA1AeehPiyA+C+jtZw5
1hsoohnfjQQ8blWg61U3Bvkhm0E++adzen/m62VvfL5QDr3IlXRmTQE1JuAW
ZSJ9HLh71f6KSGfgtEuOvix8NuLQu2FUU/1xb1xcR/gE/Wkk931E14xgwoqy
NgDbVjvQZ0hd+WTHkHtdd+Y/1P7BHKzUpAX/MnTOVDSa3iktFKE1XAhtxjAK
YoX4tSVnTb7W2Ivw0h4Lb7ITGdHtQo1wnEi3JEe4N2mJ0W0bUKWBZ70xFLA3
k4lPZC9XWGcK8PSaP3RZgkV0+YWdoldP7zo1vQNM5vLpFBR0Vv1qTMHiigwL
ei4cMyC+OYVgiMa6VM4qIaiBnW1rB9t/NRWafCUT88MpgkmAVrORVSqY8IxV
J1tPpCLCNrGOIlhgPjhBx98Q0oBsI8Y1LBA2jzTW3AM9qXL/fVKdH1o925JE
Z+DCoEbKkGtqC7ojn5llllobXOZyt4p8A/IbBWxjIxL4pjXMrD3FlJnrGEF5
3aLDX1MtJfOzSH3rkZwHT935x6HBdCPk+mIZzWzlqagmtazqh2aeLMYn1zx0
VXoUHXCRuCHnJCa9tHGndyK9TeOA3kHwT/mSxA7mWD8Ho1T+V0Tc7VXG41Fb
BTCF6B9kfUTGvqQCp6OCjglPjYJKVctI+0/e3OPrJIy19PEXl7YDtbTBoIBn
5UuBcK6OvvQhSvHeryBHeSsNns4TY3dgjMdKLfh8626Dq+eE2N7dGjM/ksQT
KlMUqZqfrO7GCaP/GNszYB6RBPD6VYf2g2uHp/wvejOfcZRMl9us9dg6z6U7
EdrrW0uwhgQcz+mnm+so36v70RHIHk01T9NBVozRrRmQdhL1eeRnvXZ4712R
KTWYYkMQIAj3+g95I7sMJcAWojIxEfVMtP0uG3HHbar/fEACK7MzfC1JaAFm
OZ+O97asx4FKmRMerlb3OlebeD05v85p8BNrPorsWVSITlM1JUn/I8EXStJ7
TlenPZuonQmZaIZLjELGd3+fCXV8EUleeAqlwatKVAb8hR6cDshAVvfq+BBQ
O7Ox+3RgqBQU2nItadFozrU0izxIwn+wO0BVsIRtEem1qlpuXjO5iiWvQI1q
DHrKYCquMF4+H/3gt3IjOkGzzow48qSPn4rw20fqLNPTzlFbyEofHe8gXsKV
r5ssun/XkI5Tr8RTQh/YqzbiJOdelgzrFCi8vBxh6BBZ29GiSrd9ERJy9sQ+
SMaO8L291T/0k0eZy6aKrbNhxxCq+YuLTROMESsGy7Wh3fkgwPLYK2aq1vAa
wraGEAzORV1HWLSMkwVVKYtdj4ixOtg8N47iJR8hLhGXVrtE9UQTdCaBLwVv
Yek2U6gqWUqiTzBKZJ7t3MhZ3k01bHyURfyPEH6qKlqB5+8sS6Fylp4BpLvb
cetBwYxz592jDJiHtK53yFs70/0aqusUHQjVq2jTKL9nHDKUBkFhvz7F/Wyk
jdoQEl2TrjlrKNDC9AQrVxelonBgLtA8DAair0pyw8s/SiiZzE24UYjKbi1X
WJyCsYDM84rqh9H2Mw7/6DNVpcRaVOptDDqgCpeVTrChKR4UO5QvfuccKIRB
dWOfmIalk+X55oVcfCphLXm+k8zZAdoFFoYhUmGcM6kDxEf2B2BZMCggyqpI
Oxmi9jEiyVKzSH6BbXG+hUAGcC+1BhzQVrKuQ31DXBdRGXX9t7FrNAg0Vq4Q
950RDmKuQoUhklWSquY4LaEDBvOdWuXaVk6IG2o+fbtkQ6q78lVsuGdeCZM1
BLX6ZoRsmsM71gV3CEBwnmmmQVKHQEzYnc7N9gS1DmYZW4c853eeMcuI9yjD
fj7RdaVqILAIXx74ABVxRLepQEarwwr3G/bk17askYMKl3ZDHzYG7HWMDXk3
gdKopMTJmWklf86kjJN1AqvdZsvuJXVZYpCBmWRGdR6bSRFdCVMU0NtREA71
ZZ1lNdDNdKyGHGGetazSWybjk63CFZaNXcbAWyS2lqy3ajqwGraKqYZIns0A
B8N7OPMt5kIPDuVyXW4KXNS7AmWar+Ov0mtw3mBGOX4KVFuYzpyFioTxETj1
8M2iZOTcCzbG/dITU1dDtjvgF9zG4iam/L4Mu3nwSZSbf9o7SfSV+nkgzf1F
DTF6MC6H6yR9Essm4qohpz52VP3xA91TgdWpMKcFIZ6dbuAmcNUt/zdnyqca
6p226QlAsc2TuZHWIS8svSw6+3ykzWHoNZM9MjHoeBbxFGlC0PuawnQ6Qv5a
+cTh8WJjpc7lcA5niRiRJeSqPJxZvbRr6YOj+h7klMnTVTl6BnLq4cNyqkz4
GQosGOVoCv6wCzvwzmLKhqIi/kevmAxM+Ecx40Ur2o2ps1YsJlUL5uVhIB/k
D+JKCQb+Luo68JOx1Br7gA0HPzn7leDuOlJMF8FyyO+jf/lkZZ36PZq0nWrL
dCTuDDOPBYjGJ+dvPGjvl18dFsnUDtRtTPShznQNHb3O9y/P65T6GJmREl7a
Tvstf3O9ql3VUxnrqqo4nPjsly8VV67wtA0LKaM8CVIL6dFvxIWrkhzEEkzG
GG5w1vD0NHsoSJX7NLuXJtdHfmMq6VJXAODM5upTPpdrZIx3OmoPQLshwt53
3l3RiKRFw01p4JSU/LZ612PcLhwsHELjqBW6jT9RM39MY8zlpvhE7BS3sJTP
HnAm2gyJme7lrl7l6Ni6PVRnskq571Xt20g3hLrlAqJL1iU9mgg1CfUzEHoZ
hE0/GFzbHyycJ4ryoe4wspHvUFyDwDVvZLzlMx/r/Z35tsvNuJHp8qSWFmGs
oL900eUQb7lO/8GV650klri0xMb92IU24zga45l78v6Cb9tvUvYbb4y9PdHj
4pzJbFr8/Zpl+aR2H/zzW1pU738FEnOnJV4P3hquTMvI4Xx5500AJinT7Nsi
Q/UYEgQUrDuE55jdy928aj8ud7av5tQx5R/4o4KtLIS9NA9nf3QTMZ4QctaP
THkBd3bGMBJ7bYGYPEFUTPzxGTjOQ2atCCfQPUNAEO4bOcecxrSem/I6E3KW
rg+MGutDS1ZWf+2xJ9tB5e2gzrgbT8QLMAoTdCl4sNBAg9Jn/5P3dPKO0dr1
aSzKZrBcudBz6uMKgVdG5uSI16jC0iPGg9h4uaW/n+/14H2s6SipR4024Bj7
ZJTGEKKXUkygfvTQ+ZSHM1Zo8VhALiifMn4atb071AjtCNcaq0sfgNl+4uQS
zCv9VqsOdrpoWjIJUXGxY1G1iNG+46vX3hBpJF3skeYnf7HyHdHXcQg8C/G/
YDuxxwwCSHsAE11VVwDIHXzlL8eG9yKCWCimpthYxrBajnmSxpOGnpledBlU
9pPst9tBV5aNB24EG56YaLfBAeU4QsXDGUoDlpksnN9znqnEsFnJ+f4OiQlV
aiHD62Nj8qa2eA+6z9QWSNJIuUH9naJljLUItl2Vs4Epa9qQgVCUwDQ13fHb
UifyMzDDEUDZrksBnixJpzIWl3NkS26jhGRaANzwSH3ik4ZG4Db0O0NP3bf9
XdglMxiOpLA/Gg7DdrIjmCbbjEn3uSs60r3FgNMMyXlMNvH42Jb/WF14AwY5
9maHQfXvaFj3o97erqPydU3Svs5VoisAduO/gDbU8TtaQsobgMXE8yiO+R/F
hqpgkDNzgcfuPfhIXwppwqccXadlJW+kL7vEdIc925tYSEpSXd6x+rzcNrN2
6YbMHLZM2saUEpGSoomwv60yYPF5QSSwqCMwxbM4vxOXgrO1amdbOZtaFKpE
tKM/jK+/TrHbnhASNV7VPFmPjUzdsqboB5dU//rTpNayREIN+lFc7fZg0TM0
wPFaSXTLhSTNdAlxuM2iO6B6QbRt2+tQ8G2G5p/HMH4AusSt3sLm19t59f0K
LYZEmIqVxf1CAjWxu1TKQdpjIEMYfzuKW0jSTUBFBZUg5bWxMAAE2pHE/n3s
YmPYH+fVUgTZDdsM2V9/hk7TVawNTnw2Qm6mrrHsXC3T19QEQmoFB37FdG7P
XhC9jmjpRxbpBKU5PyVmvGSXshxzp4VUabd8yc74mjG/9asSrIfUzbAJ5BoW
vJ2V7LaBct8ZrUhfj8UtF5FwZLcev+C9qWlRn2VU/nmSWM47TTw+b1uP6BXz
+OGJQFmBHGVOajnXGDFT3en4uKobI2/Y6/dMi9K8cxX21he71Uo12nGMDksR
PMWKcQ9MaXRGs/zwVP9hdIV2HerYDb+psQBX0AUh4EisQPj0ajgzRIEM3/I3
NIRpdqzV97529oeCGzIVLml/kzTYciKrgROgqOdqcTXmMxYIs97HsXwFjpoe
P773qK7nTvm8kGUCgN/IBWr4VWSH/SDRu11dyx0dnr67kBzXwx+0nyixsant
pqmri/KEX5jsOKGu/JYBJGSn2S5uvO4dJxiUntzhOLFs/oYcVIUa+YB342yW
sXogA4/RfdTpR6QNOKFgirTgEferHAOnEItDjca4hZENxuyctcYoMWsR3qgO
j8cVscc8OTBTbjNURCgZ61EKqF9TDsqft1k85rBKRiUb+gtKfniZSdZmilnj
6/qaXTpt5TTUyC2zaCzQTZzkTCmbWBlqqjz56wc2wAukZMoxOjkVMVZ4zpqv
KmAz/Xyakzlqk4zoB9v1o6l9sCMZX/VXNQWhM8W7VB0EXG+Ji6f9wL0LScn5
WNGL9i6rKMQbrVbjyPR4i7D3kE0mMIxMydwyAcTiU0zy4tw3756BIzl78ZUx
OPHCrAHYMPa8xH0nwa1Wts8vfWUkZ5FS3VXMPcSW5UMrdn95Ucg5WGstuK6P
Sd+7331eonCGH9oGaImJXhmL9rtMF4+tFxZcNQAZgtjfbeUksjoyEVoYD6du
e1jxSWTTe8PiBauoPFD/uxd3BDzjxvNoqgfng2fMEvB2itF7adOvGXRT5k9J
jPBjedMgeCqz6k/WFAfDH+DklFva003Ytj8fkW5NfFstgEpUjBV2vVRjCVBt
SYMeRF2iMjY5FjhCWoX948ppAIoITO68VgPzCq54RFSMgNKN7aILM6ljI8Yp
1uTAjdcQ9Miu66b0FjEZjuWYaxESVkQ82jZbtHiiSkIkuBkx5umAVR6JmCfn
j4Jv67h0Re3gm4s0qX+tYFkSzfeKFPQn+DuEsw0brbn4RttQ5OJlZa8kHt9P
8INWMr2aUcUlgsZkJC23eL395nzWd1yUNhnt3cd2UrjiMLFCnpGsE4R79HJi
3KY09+gEm+wNvCKQAtfRIuY26BQIXhFSjZasyp+PpTc8Ebb0cCa1tio4vGkr
Uh4Qzavvy/UpCBBUey1Xm2OI1gkHJk3ruFE/oC+hiCNV3tcqYk5bE66ZArr3
bvgv2numD7F1clVRE/g3EgRXfywLE7dhaF7f5xDN0nltjEvAQNS4xBzvAgGq
9ImWQAy+axbkawT9wIkM3JlyYqGdKv2eeqbvGRjOaqBC+NVrBcgQYmn/Jkhf
wnVtf1J/iHSG9LSKYBLSDZ64G98/Hlpfy7LUcf0tL4QpOajNkK3TTfIUghN2
oHPJERWdlLD3BaEIL1wO63BDr+D9i8bv1huOVU487iWzFiJnV8xuqGQzhHKG
NNC0Avn3/UwBm6kZclah28HESvwhk6A/lVt5FsQ3p9zCRUtV2NOARUAxAr/W
H2Ch/u8oxHLv/P3WTJJ4upEi84V8uxAUhMoH80OY/URu/g3k1F2HyLsLeLYq
UxqtoU9aGzm0T1nzjgYwqfk4BMZhfxs5iE2ANtFOR7RL1vxKCSm4KScVUSdX
0RJ2+W9vvQAmMsQhoNDezcrxGjeaOqGzM92Cml9pZjQ1ztM/l25S3EFEx66B
IeGVaLT6w6ETOx8MOUHp4Owq5OzZHx6k+h2dO6ZjEQpp0YRR705CGdVC/wT4
jgDkBGbUHkHQnL60MdLEoznmlw9wtG1WRaphj7S1FTyQvqMLEmL3ybqnrQdI
nfObLQWvf1hLoDf9Cars3fZYRvAVfSAG5Hz0CNcVVGJS+0MfaElXqnfLfyeg
UABhvXwF+lonp8zUjoIsi/SDnKXYOYnYnvfUoZ4xz6OVpC8kmqiBnrCW65TE
28QJH4BUewPf1hXCLDe1yM9IO/dR7IsvlOpvUEN1WQZqA3jYe7+mxvHqkKmz
QwChTvGqPuRcmDuWxBaSDsVt9p9KR9MKqWnRqgY3eGkfL8W3a/UURLcR3fSU
NCocaUnqHMTtJaVestqkVtIn4kZS1iQcajvoJh1XZX8KlFHw49NyVYCkEgct
UDdJAaek3ohCQzrtHLJYuo6gRx0gK7+Sq9HhiXwgMvLFEFtD9TB26yz09Tyt
kZTGRfb56cenSYYLXGG8+rgTOUHP6lYih+f/AFVl8caqDasNy5PQKY3jzAZ0
MG9qDAioClb6gej2LkrkbPutbELQyLcIdcNUC/0hyJUHYlLpmWlFnqWyZKd9
oFTFNeUFkQ/B8+30RWxeQw/1eIo8iHn0qN1DEhVpkX8zOQtdpbtbRiu3ZiZ2
8CA6aKwjBIuRMfLU0UxSIsEVn3wQ5swLWBOv/NRnWpSH++9FBrujyu1ya/8/
Wozv+7Yq9j9c6ZIxrIhpyDomSq2wbASvkm+GxPgqRAG8F9pK6Dbs1PEI/Rmf
jxMVapqiqyuSheCOSFBxWCnw7ZHoBlxZlLXJ86HCNBjIkilRkwd7CzwibHmx
QzdsKHgchaP9r1N4TbRmiSF5fZHqWfypgIDoo3Nps1Cb5cZ0FOppKMLmitVw
+o1eFHh8xlmbKRXwzaBD/tln1ghkDmn38ispk0fadwv9H2tGoLAOHJCyQ8tf
/hgJ4ltMHlsdIgT6nWbYE2g9kNcotclgbUyEfqHkVkW1gKvTWz2Hkk4D1dWn
v0KKiMJJyGtbvBDFlCtw3X89EKDo+AoICdnK5BQScXM7uVOEI7ktdonX/F6o
YWcQ9rc8rSnzy2zQc/HGiNer8YJmP7HaT3Y45QTIITCX+SkubQDTPtWs2sDr
iGzvTbQ8jdTUZJpCXfYIcHU/V03tIxqIzOEQH9BuXFdmEvKYNhX79uefZUsG
fgFi1Xwd/KC5F7FCQmykpu/cPdKuUWOmoaN5iSEWvariBwYKqajJZVDmHYCL
jaGHDszmXizI+V81Q6RCRGVrbSkXs36eZbjTas6w796e7Ov6VjtxtIInJE8Q
WPt/JnbXPUWo8ZRdfDKvUcOIGW2zZlSKQwM/pN0mN8DIVqhAj8ArrGdRXvn4
I0iV6ShJyX8FSyvp9ooKg9Ap20+02WN1/h0gWYrF/6nvgMtJXAUzzYY3NqNt
6dN7CwzzYNgGVtFVKykuAAFbSen+EbIBzxIpi/kjLUSPxnSo1G6EVTpPEjH8
ut/8umnwn+90D0Q/NwA4q7L9JkgxEkrRheqQAMth8/6/OljRS6G5zSq/SKWT
A92LyOUxw8AyJjIZu64GgZhBDMv882cnOXDnv6+BwSDeToxCe471F5nc751D
o9th9BShSO86iCeDVjYHkDna5gaeATES0WKjjtMf6Qx2qCNSs5gQZ6yXhbB9
iNVRG3d6wf+MSXsEwGUNxgR7tMGHbWcO1opbB7U37tj1aGysFxz+31Yo6T4q
pTBgnOYjCToVxm41yVedbsZ1UU1lWw1KcpJ/pD2txyXGMNnsVec9rmLW/4+H
Xzyw0YEsXQOTI2jwZMCrTctSHMhBLfUBVzjBcfGxbiAR5F482PalB8SxToOC
Miav0mXxa3yBcIXc8n3aZktVPUw1w1uyWfOe0uN42JtgLsOauBe3GJdjOHP0
ePPgaPBjcqlLvAeIfAomQrtGbYpO+/MMXgECTs5br5yhw+fQU8LCcfnVdjdD
/6UfmmAOf/If0IFrMoYKWOJ3LjyFQ6bqpNtpUeXWVAsNA2wk1SHDWL/SpcEf
ER48x8mGTOHfLFa714gUV3xQWIm7wgR39pITUKXHagN1+wSht4yj+z0HioZR
X9wiXPGhVNuzOrW9gQ+GNHxGX+hJVL2y0ST1iymyTASWefnkWysE+NU9QMKF
uV9imVgPiT8BE6skFtV/Vp9eS8yUeF34OwPxNYDVCN2sX5/ud2MUa56mc/MP
hmmv7xlApvNh2a9M+Tu+lTe0zZsze1fgvpeuB5XouFL01g8Tz3AtKxP7Co5m
Azs/MgOh6qSwEBehqG9QEsezX71x5ITqz546rxIKql/6AmXE61InvD2zQ6vQ
hAiKxDdICtBLkmdCs+uwM8k58lgZEuiL87jQisWQfe0lVsddoLOWqFnn1TiN
7k+tRwuIQzVR+p28iThtDhHXaPUcv8za1uixLIecObwppdcpyRJZ8oxvenNo
LlgCnRwk2B7BHZFvhiq9aJZGc54OVNlJxHCSosodVx732OO9/7SGbdOxS9ru
4uGG+//vAoEo7qCiEl4ChG+qeHy2/7/2e8n51UF/jsfmKLCQbS343Ww8bj12
x/A6H+0Fuxv9FFef5yXbe4kfCT/dN7zOUJS0DrvDZhYeTg0PD7IeG1g7E4nf
XYUHE/v2uxA7JnR2mizomE7ShmWf21FOQ672caMCOHPSPapghV7nWNahboeZ
Z0txxHETqwyMeCmXDRnebynKBsfigOCSRyrTv/e+4hujiZ6Y6xpaFxOKLE/6
xtiRM++CufJSHF2qESf/Z6acAjhxinzOd23hi3ty13G9+WoJfDsuW65cafgL
FWwg1nrQQ8E2R6xqOSKElmBChzdVrmgqh8G02HVpZ8JCDwOX2FYOW9gLxfkf
j4vzciNGkDL3iy95apxCJErWIkAtZadLVOf8gL9j6lqqwBo5OvDkQ/SXqr6O
6M1JdXo/8Wwa1Kj3VYPPd0g4dbrziNuQ4010HYtHoPJscLupeZAaB6YFPldU
bjxDoAlqgpMXSxL3LEGQV/e8CkL7vR2I/uXkDE2NPgBRaygGS0v7OGyN29OX
ZneXl/khOk0TRvVRzBc6EOvS1zrLoZW52qqefcViEGHgANHxe1bnJw+6KsCn
KjyWfzwSzwymu0cFlsK0RVDo9AP2mHbjj9Vx59Cd2zBbA2RPUOHCBOJDXSxf
kENOgkq5dEEfAE39Ct9Hzq8jEXO5p8VNaqzYZkvHBE0KepSGZvJNuQZTRwBo
XG9m1SI1wAWSzxgBTOQivEKZ/wzFg4YsWaLbvmHzT5dQV0na2xwVoI7azZqT
6EtMCNkVfEvU3fFqqBOu2fnYLv7vE2UuhxUNIIFr8NHqaffx48CfRusThy6f
8kMS+tyWpYmmmhjvpxDpfEEX9VSiohJqDemdaevDjK9FaYnCLKSPdt1MFxJR
gXL6D3kvnmDhPoxQhefjyNSY45xdVwV7y/P2BWs12eTfTacUYR5QPQ+cDEBZ
VAhxACTWIrVSQFECiIylBrN0aJzGH479S1pVd9LlzbC1JpwpUtYWjEAmIMKx
m8IcUxaUQUWZfra//nUmPjpII06rnQe8Gy56IyIQ18mI/5cy4XieFHpEuVWX
KAosw02vuSx3zm+7Am3o7kWXSDscYwer+NQsDpCvBJG9Hy1LyVR5l4umTQLo
CRYCmrmx94Ii6nyFFq8zKjMqcq1YShG9CjYZe2JHLO6DjGHwaGJpvABMGgAu
wfSHlX01sDstIj41CBuaL5LQBQ1up/a2zJ5IGmwuVijhO7obpFMVXnYv+I1K
rOWLvEG6ga+eenCtKrWxoGtaasIMmg7Bq/tXYrMVqflCxXTr3rL+KO6ScPXX
nGGIsIYYasruT/L5oHIF/azU9JrX9Y6s/JgkYoWbJsrItl66IxzzwvMctL4l
wFO/CCr+jEMxs/e0pSteDFnhAYXsu1HGy2JtQA2wffya04Qw+O1YrjRUJlnD
kFTP0hz4jLArvIBzCx6HTtertJBkapBTQk8ZvlgsdE6OOLfv+c1gvheVKaAr
zb5FnMeo25W0sJkxWJqvVyicpPq2DbOEgBB5eO03xPO2T2gplUWQAfW1CPI7
9IZmxxsh/HyJTo60jbJ5I8MxZA9rYhzNWczwo7h2w7TLXCGnVID/AwJW68+k
SjN8FTVDlknfMUz4pUUdPkb+kqL5RpVeILFQQP6NNWBXzaCJ9YhmMUY9EnE9
ddagiSe6ER9TIsWm3uLBNYf12BmM/iuPcnTZ6Buk4zgf8R+D3XI8xVIbeIav
eFPJWV5bKk02lEFesrNQhfMUu8etpkZMamXlWg8pg5aU02PiowidRmBdbrMQ
stS32r3KMe3NONG/v7uILt0DYQ9rhxE1ERfucKLwyuHJNvs57n/9oryNjCjT
vivgabh4YIx8lWZ5fvH3rSE7BgailJleg3mD0W8MF85FH16FkiLb40Lzkpzj
3KnX1RrptZCFfNpN399Vvk5MvWHwcNgEeBLUIkj5NTdeR6XdzFDLn3o08+DM
mwVh8d9fw1Jb1h3J/Ihgkn27aWVfYKBjZmR6UcyLOLpJvQdJ+EN/8Bh6YiuH
OrWFdSJpMe8W+7alqOORhg10zoKG6hF8dwKYaCY/rNV2Qfp0C7zdiM0pFsl6
aToo1Z3gxi09IDv79jKl+MNquf0CZNSBf61sWj+A5jqclIsEW833/Eyz0U38
idc+NagnGyTD+mzIBInJaO9VBDhnVFl9n/rWN+G2XKF7d46Acp6xfndGQPtn
Y5HeQjycJqtqBUawdOjyCYa1okbEoz2bT6LRD+WhgN373Nz6UQ8d8hsCP6Fl
4+Q/DyJEWktL145xm9zec5X39sy+PuiGuk4mxpARx5QglJcRNFdm4y+SezWs
Gj9qlOFBxaz4Ywu3+LdW+FSljb2K3DLl2CL4HRewHHOCsuuDFWfFR206q5z7
m13Dsk6H62yVkue4fEjxbMUAbtZXHDyglhS8yFYwhY3MtrCoMRrDzojjcXTP
D4j/CPqOSNU53cyAHhRTzZ4W9LSg5UuWNtpFzAawDCQghtKYAkq0OwV1bO70
jioSHegd9gVMBR4C1ouIiLWZmV4Mpj5kG6fc9z7b64Gy64QRi0bHC58xoKbC
KCsM79Q+aVOIVx+wVUjCCmj9I6lQLbG4DVnyU5cmypoPhRrc5QfyzA0dCxRu
5aU47WYAvhQHIFszLAYzYSew6GgaKPqSvl1Ae2ePGWybSY6ScELMUJdZUGPU
mr2xqG9ivL+D3D8uotpSD531/U+SMIYw2Ct6XxZQQVuId0F0pEQ1TdkNj+YY
G8PNREK+2xKwaGVAZgk7fGVVrcXnl3/Y5aUbMXw8zhFAdPpFSq1nucygnBJC
8WWr0BbgiyWm3UMwyswC0tZK/GU/Ix+RL6W1qxXoa6ks/irazhyPxKBLz9BB
OXuMcnpRgkx338GsIHF8w+k5GuOXnbr/l3XdNdjVrrbZjpVH7Td015E6NVV6
c/Nqy/ZXfKsha3RetuQ0/luQ6HAvaQCuImsS2CeKyMnfYLm2XHu+Nmcc4S1b
XD9fdtNw7u5ZWz8H1XoKoXZRIoAu8lucPpZuJYG8HD/OyRFVgg1zyOdBDEku
f29bMJg6WYiV/EfG41pzh09ShyxYb5YgXfh1TY6eEipx/qmg1AYZSWuQDqbO
RmAmTCW9iSMB1Wj2aatAZCgI/bEHzts67Uqo9tF8Evc9TPWWPjLT/R/BDPWx
LlWQkLXcZwdCn+WvBdws0eqthEAZ/YEEFOf7ypuj2O3OxF67ksYAKNwTuvz2
nMgTN5cdhAYsTXRhc95BSyD3k60LWzW5GPzEKqaV8VrkArrsUCrx8fgBYu9W
ZgMFULrH44pc/uQibWFcuQfnk62XaZjZ/w8Uz7QTYOtxQxnLX/fRUwUWpvUZ
0kZlRKsPnu+PUVvmxmqkIeoiYTCKhhkcqOo5QUEGGSsMhjlAtoslzBTWyWUU
CUslJA39kKfu/XOpzCKSSf80XSYopNVhBY66QPKFSFXM1JQRx1/58DWbSLoo
L77aRn3MGomO+Wuzfgo0XNQNJMgAz0aTrCF6klooIdykEdfihPjjTfiiVwxp
Pi2CLmS4v+U1HJ2H05rF01smCMCG/yJepHkbELteWrLTRuSuP9E4WL1Zsi+3
XgxU8/XG0B5PfkNPQi9SwxHwFQYkuBrtyybsb3PRAX30WiCrUU7uoFR9z74/
rtt0pHI96ZBLh8hybKKLiJkEqTlETJindpn/ilWh46gjNxVPDY00dvTlmSpS
R1V3jk/HclY78Np2fXZp9z3aGJIhRM9o7SarDSWyPgTMQqD1V/9p2o3I4JkF
BCDWrvXR1YqDTh6dyFzzdHiBzGafRM7bvV8DmWobp7RpkQWVRUtGWw5TQut5
/3tbMUonwFs+ARcZCPTVJm7v+kohAJUZqusV8EdKdCkyxosVNSToMSno7RJW
rlZN79gv1R97MAv4x5ZUcbZY8zZrkhqk1MU+1ODzN73CwYlEcyT5+3/o7G8m
a4kmuOsBi6jOq+zOw9W2W/xUY7TD14H3P5sYyFVoviYnQz52BYC1VNTOUVWi
g14va1YM2aCe1u/li+wAsh9922OILGZBhgeA4c/5GBCWQaw6n5bNzVWwwplc
h2V50SC5kt40BU82Od6EAaWY/Wt5yo05aTdEW0F6xJiqCxG2d4QjThLvAklq
xrLIacCjT7FfLVGwMszmipVCH6C7T0lDtY/sHfHYGygypmafA7m0yCKpqFe9
rV5gETz+v1JVbVubupL0gm8OXTgrNjnwTbX4L04OcRqNIMk33YzMXYKBNabE
j/Yz14LQiZ4/9MGNCWdL6u4PKnJlYfzRM4EAOpghvoCk/o0QAY0ABpsk3YHL
aBnh6n4uNNpHaDGZMhqtLxgTZKQYLC1hJAFxAilkUbGWphyysnooejDuNorc
oUeM7pcjaTUYrIW4aNkXoiZPL8FLmkegHpMH6AfmDE8z6mPmlho7teJNpwZd
WUK/nd9ZRtjutnMuxiDuxhvVbvDN+5plLObVN1kf3LSQt7pDHYrgbmnm6Bvr
J6A5NdA9SBIQSCzggw3wai/huMlpSBF+yySbzlCOmxgi+8Wtq6zw8diro/LF
QUNJcpf3AY20LJsqiY/wHw7mbSWg2SaiivuVnPCRDZTIkEL4y8wqXdaudb7W
soR+u5+oAwOI67ZjoVr0d8tWRWJanlKxWLxyeWxpcnvFWe5b2LMtcTEoDWhT
K5wEEN4itwJzMH26cXsivlxCe3JGnDvZc8pcbF9I0SGEuCfGFvR3b3ETdRv7
aqU86E3/MGcEL0EJdV7f2AxeCzRw1JlmeiCE4vnf599JCbfAWfmQ8Aqlf7P4
IFZiYwnmqtNGWkcbJfQH7GZtUNrEjlJaJbhYrTjsKy/GCjZ+HA517cAydpZM
ygQuV0HxU+zlLw8nvccbUF40l/P9geKQBYjwNrt2scFlkAPLtRvzfsi1dMCN
6m/wRQnZtxtaJfO9eXCZOhhhWcJZE+ltTa3xk+GA2e96gtM+A52sShX/G0zw
YoFUb2MKZXoyjxgF57GoqIgmiRhjJVnv/nkEz7jU/ykw0ZOtqTzSx9zYg2JR
WD9G0yz+NTvi4pR0PDqPd1g/PYj3LJQ6zivtQejM3Y03IEb+1fFC8KSk7LHR
63YrCOaBSqRl2EXSp4NRN5GmI/j8nUQgxi17jSY9qQkKvDXmOQ5k9YvYu4LQ
djRIPfzz1WlfhZoUjc5T7yq+ZvXd/y78N+7AZNFoh4Ks0JWnLPz7ev+Vh9Y2
wrwWgAYmFNDPnOytWW/TH6CiB9LRJecAlH5Ahy+Abo5NmfJHYgqJ8K/xqeeg
u68kCNEbsTk1x33JJ+IKFiun5mKlw7cy1HBgDraCku3U4xKBx5BJUzslDr3V
hgm7zdNNOAZCXQromxTXKJkpccWkSDvXUAnMLlLKcgy911cOgRAasAQRb/vE
bjk2J3rJngRZc5BpaNp3RZM43ktgryBXJPD0qZtRMzTy/LGDPuN928TVUcU7
ZLExzXRgDlR3ZkyZ8pknzyYT6cXxfOwFcuyRA0DeYaN8UfPLvRkz//XkD7ft
2ivAb6ymXJbylHRcZ71dX9F9fH1mzEYg32RwHhY5wZ+JNhTJEnJ3sjYvMK86
Z2EHwMSZn1gIjzO8YSqKSzWE0WQy5/eUe333reLE7MNdpi8zAFAZIXz8qjL0
pQgU6aTjIOiKIn1B0gSmX+oCOvB1tX8JNxk3/pJrHznxpKAsXShi8MVrbVon
7O6U80NlX6BeU2FVnYYE0RC4y7XsBoSJvchbUmsxj5/1dJeiJ2QVSw3AxKVP
6Ed4HTPURMv8dgZ7swAKpK9o5CFNzltnSXZK3rtMDuViBW/F8R7aiuqaSPz4
7hZ7G8R6NvZeXZUKRc07TtJww0iUtJ6Jeor1jOlNk1Yfvg7ECsODvdMZgziy
vC8iCRk1fbQkWhXHlsxGnaKoykZYE01lSemrEejtBvErpLYrRaVNGNgPWLFv
sUn9ScQGm3Lo6n1TYjuV+k040tBVz7tzSUwNBtU8yKhDz+JpQqGfB7jG65M/
khh6SVwrIeXmiNIuHRmZHZjWD0cU7g5e3R54TLrzv3DyQB7DKijVqChI9Tq/
GHE9pizA3BlykWZBH9ipg5gjYm20+eXfJRKSDRhchXpXB9YvHR7ISD48/do2
svkpCZZrkgwdZ5thwj0SKgz53kL06MXCjyX434RR1Wr7KwKUpAAPJFGBxSZn
vMPp1IyOCnbmd9q/SM3ITVVBcrTp7jtY9Zim2QY5FAq/mWbFmlVAEYHLz0wU
MvRX9w9x3SOu3bcs8JikzfcJWv3MGE18Vj9fFwLDwxsvXWPjTpGdrpXaEEYI
hMSjxt9Rp/FapeF5ccMc+tZwYgNNGl1b+rUZuWjPT3Fc7CeGUmbv1W0/JJqD
cKdaU8KNi9tDZuUgb9O9kSd4dLTCOYJf4sEj/9tkC0jo/Qs/HLwpqJzioDG/
i3BbSD+PV/Cx9dZJZCCHjyzjyUAEb7EAvXabsz8f/kYogHgwek5CtCcVNQT5
GwxK5XjKuGs/EO28EcRfxmVYJ8rUwj1b9Bk847JZ9vj+jfUGOKnXAtNslgHC
b9P9hYE4FN0psIAe8KgB7n2AUrRLeMN1ktgNZJWPADvQdzNcFtDbBLWCnyHf
WH5F5gLNhcLFu40F0ljC4K6Qlw6cWt76/xh4TPMQhuBP3gEnV3a7PSdykK8a
oJ/2kmBSrUbEvCLENnr5c+J5FXFpDXy0CoOQppLY0dnDpmBLqdi8AVoll/in
s2v9VORQzsrD0Oa/9C8UKiNM30Ra20DvuLW75+vRN/jwh/K9V0uQ/vcV1HAV
WtGY6HfOd/S/6aVQeUWmVUH4D+JEwO3TUv1QMbLpsaRVBBKNVl15+PdEZkPq
vrFtkbc44QNhthQHTraZFqMlgrtduWrSvb2ytNb1vckr3zGMiVKVFWlfprPU
tsi5BtEWX+In5DyGunr16KLmmm3Jgq8kFfsbRPZI5fSk0dzGmfvoiG5OcOjd
73h6sUhecXcmZNtACEJyGJt2NKgZsVy1x6PaWM6sSIZcmXtyc7a3pJVGhlDD
Wlwqzcy+3wWFdZ1ugF8qo2w6+tzzVbkNEP07O3aG38sIW+8gMtXAhsl0myd3
FVi+8oGhTK3QVAy9U3Lf8SgNjQV5dWn9MomiVT8MACMoWcZm9nwJWOGEO3fX
2lDKiR+1oqcBhDA6RmuhPq+b2xrAwym8SJschHw/slmxNPFVzcGSHfrEh6Rk
Hzu4FxzQwOtD4TSVI1me6twWQUKlCC1HqJfkvWLYHiEPBD29wNg0xWDIfDvA
tpCgCdlDEXNVvx1RlauyS2f5t6D4bxYBrzHt1tcm93KC8dRbAGztVeMsSn4B
FIt9nNLeNcyhxFHHA9B+n7UdoL818iKi1sgNFKmu9cHU6tvr5H+6KMGKxgh1
iIJR78FeOhb1sr84XCiPF2r6De/3n1r+l9yHNZxndYedVEar2d3qK9gmhQXi
yalMdpb/4mKPBOzdZ8pEs/cJAC7YouR0JHcYBoJ8yQH6PrxSXdxE8DXc+EKY
EbBTun4ZU/QIPOvZRL8EnDvCDlcAxPjciu+CTitlMMqrXNKyj/mJdFOdFLl3
IWm5lws6ee/fXL0BGyOZfj5Jyq/TcmLOjtHp9FZwQgxS+wZm74YSgBbZDU/f
ijfJPaxpLgVXevvMHhKAKzy9CHlLBEo5hjz38YT0ZM47EpImydDduhINIFgZ
zzy5eCXX3fizp4PH+/3TrY/6Dna/EyLKnZhM+XMIFCyFDFx8D+fiAyC0d6yc
13kFH2HF1rHNouAhXl9/Wm8hQJNdfFkWZASw5zqLAuZYMp1gq3RBWZqVV+ZG
wGNh6+LLC9BxZMXqIo3ZtmYLujpNt7R1Lv6kPRD8QwDj9SKW/TELUjG8xuXS
w2/jgoKFXuNhmNcxQS0swpA9P7kj0poyCJeaQQetV2XgToe2tl2GV41WgXDH
SyW/r3+A5HBSTFmkzjbEjS5/wlKxLdpbp45cARY0y/lrhT19+zxRqrNkhod6
+SOge97XTq5Rgr1q57KSJ/d7XNDdC57EOFvgf30Yx5rECZpt4NebaXSsvYTt
kNgTyR2hM3HgBtNme/yhI7TZS43o79iHKALlXVfdksCx1QeNUhe0Bavv3hOW
5gHbmYlTVOFRNAP0PQItWg4X3xHngERQ2VvgdgreNXrHrhGV/KlbajHUjgKR
+/bO30OQdwOHcsaIu4GxTC6FWzsYVObW6mRAaqxoEpjkDi6ZVQYIXDQLhhf0
YwxF1tjD7IDQhY60L5Fzpb5eq/YBV3lFmN+btlYSxDa7FSq2SISQytqWC+fe
P1bqY3pfXcvEKDg51RYPm7HiPeXzV/7B6ESfKLSMksBl7htT41MH3bqjU+4O
ajmDAJCuOgzxnEy/JXJeKyp8JO/FQjJ9BXx0wNAiD6kNo0rQd5ZlNPST4Wjz
UbOoz5dX48zA02wTXR2Mw54NI3vNXLaDBsCZbBV7fQgVT0PerCTfXjjlTrQF
2X8osxNTkG4VtnboaQdvJhm6yqP4TWs+U02XAH/kSAuWNFXG7PlvXypTZ+QN
X0TJ/PsUlGCVbVk1TCp0VsSsvrPPjkw8d6oTeejc5KtuTNZhX2ZlBqGFZxYt
kD6jCnUfpeGjY378u+dxzBQmvplU9pmzWNsRTxtgncC9rP+6Yszb+jBtKAYd
PUH3B2gKKfaVKc6ZG5JgoR/8vuqE/i5wd7OehlYEibCd4b5gOSivWt2UvYxB
1FpKwJIhgJ546jdKsACUR5jV+Xqry5IRSAUFWOoiK6pYewIqx1WAWsCuOBIl
3RKtfU5itZiW5vDYDb6oSBSD1yE3vkMA2zA7ZuDtcE7bJ2nJ6ptAsGWTfQfi
swQRa4E0zFU97Ye9XQeQKoc3JlMSD/jypghlwElEKX2CfxKMsXbZ9NXlLdNI
CJgcbv4kqnpOlAT8Ufs+HhsQi1dVEazy7F9DFV2r8fEXKcwD/14LONoAesT1
swizdSYpTqtTckaBRCwVh6C0PzfilQXgZgWagg/c1fqpkujLV4IHe20la+Od
c29k8N4yPjY4UNnkr60GV9bCGTyMWPC0G3u6QYJ25SxCOf7oLdk/Sdh9gxlg
yOYWauZ0IyVMbrwhhnKE4mYwZYjuHBkUC5NHmToFPddjZ0YfFql5NjtyeVft
Af0kQ4CcPygJpc7ZJYb7nokII2DT1whI0mr/DKOCAXK7rK5O192my/tpdwWN
ma1RDHmrAet3rArnT6rpxAUY7BhV2YS2Tz5ndSoDnslMwIXH7Nz5d7m+QP7G
j5R2u31ibCEwkYG7qrRZU5YgUJb6e+4o6P3cD83r0ugMJoGwHM5mqN7U7oSB
78oWFmv1SSlALGZ0NVO91wwiyCmgtTTLTPJRz1zW1OLoTbM3bxfZ0mtHo7Fn
vL5STScWeMOoHc80beI0clJLORyLoGAhbS7JqB8Dk1xmbIrsKMPZnK056ygd
zu6ddxksYHTQAXIPg9dLuREyIEUmsl6jPdWcbufZGRDXsdG5V9yu9o6rQPBo
AwtDVM5QuFnM0YfXL7t7PQJfr013eOCf7bWk1f0Ynj3LGlMV4zYQR1tpkt3c
Sx1vJeu59KdgH6R4FFZikZyy/joanl76H1K3/ANLJd+iduMeZIx87MPnBPmk
pBPfNQbI3m8Oulqoj/NfCaUOdFr3LhgF31aEQcH7Mp4zJRlubxwDN/iNaNuu
VEwVdCcQcpnw2DdVtGabgQgfa0J1l2md7xHYg2afsl/ygQLeFyppZIXKWH9E
cyp6ustHY7LBsi0TvYgm8dc5+YD0AQcfYUq0077IAYxIpOY/n0IVTrKi9pWr
uXEmzYYxpi1/12Vmhncjcg3j0CI2RhhW1f4DuDBjMYTtT4/fs+nEusSkYuml
KWVp5Iq8d8DwzMmSKuDK8kkPJNWqI1Hu8E9StCO9bAEYMG1PNiszNskOBPI4
ijX5HErPoGui67wlr44c3pn0XsyjoQAVAiLIbbIZnuVDQ4RJEGVBJ3MqZzMg
PSHD7wOFJHGidpVLyWF8gcuQCnauXVWWRMaZIF3ntjH9JjdN2xNWWSA0wJ0b
91rwL9T1T1Td83CkG8wcRd72a5Qfi8yqrCHkbOEwT/Dwh5ihJ4llLJmWvFnw
L82TIFSS8O4zLQyvvdt8l7yW0V/txwWQbWo2/Gl6s12jnr710oLUe9Yrsd0V
lRKTaGGyUP372WC3uPGAfnkF8NMUt5lZBNPECcj0np+/qCHATr+u330agyqW
LaBhD0gl+DgzgGxccFMOtd6rZC1C4uaY4nuM5QlEBMOM28M9qMxV2SRbTbRe
FXqqv6A8WnMJM9V1jFkpZ3Md9MyN+yB12GN4I51Y5iYydClmyRd4pZOF7K4W
cvVQO9ZXe7nHS2Eg8hygZz0QVmS+wErNJw6SaaXkJv3RrkU6tvZggH2dvB4U
hCZSW4mMFZ/fBwcw8gi4Rk/niKJ8ZuV4yU/GCTuIYCqxBR6KfVXxjNiLUME8
XYK/hjPGN/Z9uEjI1NRR56mns8JC6fgBX1XsuuYvQptLXFO6jMr5TWlAZWkF
nu993HIUc7//KpxTrm0JDsxZRV9qbR6DrbF9xU5sk1v7BFEU4bmb66FC/bBc
XdY7MrXrTcanjaUivO6in+5Q6hk4QkAuggv8+pnShP5bZTpI1T3axAojsvsm
skgk11ydRXN9ZnRjZk1fcXGqYIvw0wZR+490P0xncv0evog4jO8+wcbA+m3W
lu4GHocXRVMpYpPafdjYWM2ZT1tBEhKLMPB9BVQpsX1GmkXjr7buk+2l4Z2M
mJJaJp02jDXEZBsBP7ikiDhpBtNDTXHV1TwJ0gHZwMeMyWA+XR9AwZVVFDpx
rM71E3FHuCzr70X4wB489BQUy/LHqy8ln3MJKobPhb4Rxcl+HM/j7wG1x1OI
HATaxp04bKa133OBxvxT1OHV2iyDabHO1MtKNmMtd3TDGuKq3NV1RYsWNeUA
FL84s1Vr/hRf7VYIGwjMW47MfwBdfE2V86eLRWm9aVh7geIpEwfSpOfHbmPG
OkitZk2xAHU0jU5Z4upi8OlEL81hW5ABJhZbBV3kSOEe6kJY5h5RjJ8pPNkl
7krr2IDXAqQlcNoKnuWxOI5TOB3IWCDgLk5b/2jONA3B5iKyd77vKiTcmr10
nWs6vJMY0JhqmLCqFz4Zk6DeBgeiGrx9xaWECZ2iNdyRo7ew3HuCjxGdTI/l
FE60q2JQ+kKC9G/zxAgqDZ5Le3CKs1vjHG9jeM0EcDmMUiJqDrYI0rYf0zSp
k2O7nW736JPr/d0+56k3SqswTIbFZl6OcB1L9+voRM3b3tvmOZh/GY5pkfYZ
7h9fU7pUPyhkEJVp++ACN4jHisaRuTSoMOah4Wo1xco6K/zxW6PTCI6EjuYO
+8p55NW+uWMAsggwYZoE4vjSCbnZtjTA5BHYIUEtSFvxGsR4LPowr90DLfPF
LDoQuVZl8/FM1ogZ6xRQgJxNDUHb1pq8O50qBgd0gqGFsl80kLZuMKJ3TR9u
jDScYOC51Q7+L2P9EnfVg49OUC+4aNPl7i/EgROVvg737E/DfSNRC4bMg+6l
q0RkbJftH/EADgiavHLTG8Ksnspz32VchzIWfnE4ZT75iTd52ld8DJ31wS9p
fQkClNhgK00PgM4GghgzR7KFaH7Ao8wjy4+UebyoRL14kjiy2GWritUF6Fn3
y78JVrIX7f6HEJJbRWMR8r/0xGTBHdQC29+tubPIdSnc8SqIE+/ieUun6pcI
CZ4ujVO43X/bBRCJrZ8WZQOPr7h4EUoYCz+/1QX+PYcPH9pAboI1f6tc8oh4
pZ+q0hFkAtfhevHhv8/j+pSRXhQk6iSkIhWHmic0mxgYmOH/EskezugTEO6M
K1Tv8fmarJyg5HSQBcUVCeUngZqqw4y9/9fJEz+PaTpyh7TsKQ+UJZT8NYFD
aEfjIoRFAHK52gbfUUkJFKFZSz6eBGc9MVPI2f08+AcQ3M3bIyaeFvO9LpUC
iEODI1TyopX0IsZ/+r22X5vZPIvYSooa+lq1uYvmZnNi7n7OUr4FQ6b/oh+o
aWLK0nHdW5711cuoK5KfGd4tiSHInwzxOktKujeIjdKQaDmVPcoqIJSYjVXp
WAfemmIwx8r8vkmZ6evU3XC/yrzxGudDGsMP1AnuvAVomVZZhKtAQUtkGI2Y
QeE9pRROsSlTKTSzffG4FpP2Sr3xnLN1RHpitztQqrXVZYRC0QqOl2nq6bzh
K2LsalMsh7BEc9aQ6zlrrJ2Soqcha5u+czzWq5vRhVyxk4p536Oi3QhEztDC
uuLTn5Riqo3eBwPOINdnEqa+7S4KsEcP+N9hNjDUdtqEX5zLO/mM+9kIbnvr
cPDrrV5Rca1jgl0mb88H2xY66DYnu9AbPxhC5BGbdfd23B/cYW5ntxja3luZ
zX1Xy+FUYXbBG1LpCSIP/ULiL1CHSP4FbbnKd/5QKf6GCLHHOQFQlRv0Fv3/
KYMlypC0sWEhGY5lP0zJhB50fjnQk3htYkaH1nVefbwD0CUzSFyCug7wVCi9
udGPQWr2zKVW3dMM8VJWx1TKAqsIBxU2uxDDwDTiOKJPd9E1L5SJB1jAXlIz
bqlJ9vFXVO76iw2IOhlo+plRHxmM24KvCd75otrzgG8iANgfmi5hOEndcQyZ
CETxUwyFHbduLNGeDEziHUSPe4Y55sqWlgfpDyU2GD53/I0q1x7KQINNHgKW
o99uOICyRTpCSRiSo6AmCOXQjASGxpKMvfehANXlg3NNV+wOmQl/X1x4mFsk
Hf7ry8c4FWXOhE9Ngmyu7vktrDmb6oaO2uIVL0iiU6fvIUJ/YCMoq4diwAx/
NCeKCHxAi0iBTeGDsBEZhQk9CYqQtFXByZ1RCl4LOxRbiTZ8/5waoPiaWntG
pzbRIzb61BX22W/G/gEejUDRYeIJeGQsRKf3v/Ek3wpUWZ+fF2nCrmKYOx4M
ewaPy7UQqiZ/Ykymk0nj3Tui/sHxyhhw9/k2IpJdEk9pZmFW2EmoIJAxnaEd
ccTGFu/Ep+y4lfu03K0gG0ehDXJU4En6KUCO1le3A8ZKPjQSVFRyOCoMd2bX
40YrVfyMg2VLlYYu4LyEgkC8/gXMOq5oa13aVJ5WDHHswJb2mfdziF+yeq9+
FJQ+HfrsdBQsZf1SZQtDtGSh3E4GkwENYF296E1PU2cseKfy5AHKe2EApKYt
0ikTq+HwnewOVAno79QFEezwqNyZeBu/8XK/TouZi9xrJgFjUe4fxTiewZ3y
tbNshJZBWgTHIisdJLmOUZi49T1dwlRzY9VttQA5Hamc9/lg7HpwlFD9Ac1d
PBlon6pemgNF9eJd0q7u+12tBPxKTQTltdVHltJlbLPCa9rQ6kphdXjBrTkL
3l/mpQcKkcZEKvCfp5/42ma5dDEkdaN/XK8Ja3S0xp36fXJAh5FJaHGNYkS7
8wq8JZPp6xjecxd0Q3m8XxL8RZJidKFuh/lcO2vrhDAXaMLbyC1y6i8y0hbg
TFEb0FAUNPOlGEulSbQcBsn0bNMDwW44e94xXQ6H8jQR+8YXqSH6xErbIQRv
Fml4BJZG1cIxATxdlKX1lJxY43n/rXslM/F/sdeipc9A27LNMpDN57WPmalh
FlrAzA6/Pm24m1fJq2F4gKKmTfYPd/EUTZdb8YjrIDsj4/MBq4ZL4jXe4t/R
jLk5zcENuv+yREU2qI6Sohn1TjsLQ3EFh4HVc6XroGymS0qKK3xSZD1dL/a0
VVQ1/uLks91NEualo+DAzC+iTkcRTHjiZuyiomER5FdFXriF1GUkQgViSWxI
JijoWVvgXagolVst+cg5/K9VrC70NOeS9HojI37apk+YhkqVKWGvREcEMgZB
S1tdOYZlczkJaSqX2G0lIc9YgG/DfV+ttI2GbVTCaj4xudpitVROfBd2oPDZ
NUkmyGM6+460N6K7ZwLFndyN6GOZ8TeKbH3I7y1TdgANbV9yXx/KMdYBKXC+
U7WwIY/BnO9bKFkLh5pmoeY2k0KKhwx/LWSHfIV4Mm/Tj1PHyWaNUFeeukJa
dvD5m7nEDYpkvlopQp4UMrFeQmKUe314ZyDnk4blwOo6NEUme8y05teC7Op+
NQKVbFbBsjWZN1ktuzoIPYrKjK30qdQ/ePfNppXiD194hJ9ctbiHAjPbT0EJ
Xe8os+AkausaBzi+gQhIFg3bw25am8bwpN5MrIiY6iKQaH1zFAvGmzaRhLwk
0FuT0lDUWhaDebrf7qtjaX5k8+q6MD+v9qO+3gxEEjcy/rBIfoNPPDW1qIKx
z4jMcFZhip8qa8NNnVbdQjozt5pBUpja1j8+569aMOn9nJKvo1pfY8cVvn0f
JniUtq+pj9JfxlvV0p8PzpKdE3ELFRBbq9jhh+7i7KgXdlN8h8IpJrFYtE1T
GSxWu9uogCnARuD7HeoF9V+uCCpFBZk6nFVRUFvQrLnmV79TlkqpvrT9yFfz
2FlWYgg2nNsppnJaNvSRQV1bhFbXJH83m+IjnsD6ByyBimrUb8kgrGgs8UVu
5T4yNEhuC3rQsH1Q35Bz3P7QXhn8ZK0rV/pweRVK3dJBsZBi9fPayjVYLsQU
WTQizMzVF6+R+BZC2MA95OVRqFhw55GoPNZaIolDJ2N8sOx3moKaH62dOXEd
Dg55KK/Jh9RDVOURdILeVYCmiJb2G5EwkuZ+TlYmgxkPmFLSCzoMD44/CODS
ANS4WuAnfSoFmyXsMJa2aFzXcGfuLd+RI3Vt/xSkkQaCstX+tJrys4Yu7MH1
3iSwN3ZWkRWGBrw5AtAMkW3BFw29advhsr891O1xvojB/hbN1DLJQwi64n7X
x3i4ZKrZUFkPeCDCimOdTOD2PaGcvz9SeQ4gofVhueJg0qgzwlKlFDmxY2Y0
jaLce/pikIMZ22PC91IrdmaRoLusDTyaJ9KkgfO5ZSPDnnHLMwSMjl8rv2Dt
Kgg5ir0vpHm8881nL3Bp1tEzB9VSvCtGIW6t2ww1TTJrgckE3ZZO7Z7zePGQ
ZM55UCVTmBQHZM7QlEpDb04kOTQMkfMjwu25x6q1nLaeB+10cKgOuC4ZtPAR
AnBiV7PBliR5sHEbjyy4s5MQpvtUJTd9FkgAiHvb9Xt9uJFLbgFwJatdjod9
9Iv+PhFy+g3kt4Kn7NDKiNcW13N7kjXVC2ztU0a4ajniFnSr1wfnzjkhh3f+
EfrEeFk6GrXL9Rt6YqIUAdSe295SMdZWNu//CZz+IlMT/LWOe1fzKIAXqvVg
2qYbnznBFWOG2Ebp1z6rIaVCRp4OHmyByd0gGGRD6p6liSdNh8o+P6nt81JM
AKcLUcbuPgHaP9zBFl0nZ+d2bBZutLQ24caOFc/byqnwxEYDR7ANDIfI2qEK
8Z0tmmYgQ/wQw17Kb2sCNMKNSDV1/5OTAy6U5cgkLbWjrdZ4nLMQQsBo2aQ/
+SEBfDUbWc+EeEpShMzYiljcwvAk56ptGwNtEtBLwfdD8hQYEyC+HfjKIxbh
l3xerjqDtTtpqStmtK/pFWu9w+bxQqQJSc3fLBz6Ia1RX2t3Grw4EkSq76BB
IuhoT8YbYoGxOuzW0PJQU9NYfoHK0NIjm9obokvueQNXHpBWRC5TFVbwWlfg
4Kwu632Oi3j4U3onirqfo/LLVriE7vSRUUvO0EIUMq8rZdnTeD9Ar5XMtBSd
gLUh/tmCFnodd0EZcxX5FlgyllalnaYaGFhVG6ItlaiKzfBNPBKBjSayhvF+
cz/a61FlgePlru0QfGofmxkvQqoLcq1wOLsbhnsmdyqTQtM0fdxk2hiEHvYD
r2VXfTHlF60WKq/a+Ve6TDK4ZlRYWV0chV4/mu6OCUv1OIWLcekSf+hxmVEt
EfhX0WEv+oXvj+UECH/JoTJmQXNPvMJ3CZm9c2470z+J2TobAupzH2ANyYKK
dTz7C0n8MyuGopQxkEhtX6uNc/OjNm4nd71uXOWp86AXJ154lAM2F+BRdaQC
ap1xN8E7ITV6/XjlTf0nk2mhl1ouoMnMjsgCcLlR97KMGVvshCerzlCpZ69q
yCVPMz50AOYDugCMtOrHm+oEbLT3Me2oqdL9Q6lxhmPMWYBEhCY3g8u88NnG
XPMzlj8w7TO8DBv734BxeLk/hFRuM9+BtUi0RAedYuOTcT59P/vIYluYrvRQ
+HgS9jeNny0aUA4QYNqEQCc6i7alreY5O0BThLpobevAAa+4GWm9L6z62cDP
Sgtf/P05MLg6jbERhRnoNkO4AgffJqQr/T7wdRIA7SsH2NXD+8JKDhluqy7g
kdXAN3sOAQiELxRn1qjEttLvLviAUGjY33hMo5qX+7wjgyeVVeI5qQNYOaUg
g/6enmdmVfJZsFlr44FRbGwyDGOHv54Zo0SQ8glcTelh+K8Oj/yjvcJx0ciC
HYeJd7xSSYfXbAXEEaTHHEKzvabQ58DA2yBsMAfGPsyupYLqF5X7Ri248Oxb
h0M4b37apVXGZltRsIwDZ8dSnNmTcK2kaA8XU93MLfiXmSKIodQo4rxNiFY1
eSucgoI9pEehsEjEfqRra9X+xhHAkHFnB52vWLRGIZwgaML/+pLvBs6dvj/F
hegdjID2WFGnY/H1kXJZi0/SsohTjZ/8FE0QAkDfPQYXLsv+8hOYaTKgBQww
Svl/kEN5HHHvRSkUZA99Bv7hdFHsGSGcmsMWsxdinFeh8XhzPsNhD3YLQ9Cx
ZAeH2c4y4McUjaoUyVdGktKvY+LydPMuEKA7T/2HZwlSlVGcfZI2Kv+hoYAW
luHpMEOp4QIliHLD+X0RJDeEDQvXZe5M+jernVpKfCzgAalvzxc6D1EIr7j4
xQoiGFfQ9S3Ryum8qyy70UBuGox1c1EdS2OwyM8tNkv7MXmymBvvp05UZMl8
eYoLRGV0vZFQdN46d/r+Ur1egwhoFhPb4oGyCbPHcOC/SeNfY48C6yz5/mp4
6cGoKl4TZ3dIVFVaoPcEjLxWteDPvwJeNxbbwJIByBBS7B4juaUBM4bY7df1
/D4hjf2yyVWDlkBcVPJZPI70jV0c/M1lcUnPU1Tg4jCnccXRz05TR6R4NusP
1OBvAz6u6nzsuy3ZtN++zh0BC4SEoDcEDdWvgGnSbNbmNECA7K+2TuL4xInj
peZzr1+eBVQ4oOt8LBWcxd8gkBOoesq3IWch5NuU89qfXZYwjASymlZOASgJ
UYsvQ7/zKrYTqJ5e4jICI0Eq/2kPf3rxwwnAQwGQq293msWBPp+TbRUxwF3U
k8TQt+TxOo1bqDyr6SgUbiLU7XWJ9bEZCMKhpOzAr69QmMiCNgUzy56ktUam
ChtSWHJBtcmWLlwSYrV+Bcz7AxYfz5uB0HR/KdclLTmDw4kWJZ9Yrn/WLuvz
iAJeJvkheCS9BxGZhheCoVTdaBDpQpqWiBNOzVJBI85nPSt0HtX5YtUCXovY
k0vtwHSIq8x0/fVDqJasC4S0OE0j3f1i1fyoDoFEqIbl+oTqk3i0YNolgqTU
SMqNlD0uXajS4sCnMqlXew5NObI9Z1IqPa0npLftVJUnmZCwBZzEIsWkrzzm
r4dgvgd59hEspMVuCa8eWevxQE4v+XNflLAcgYBTlDRwAHSNcKog0SobtetJ
4Pf1DV8MIS62FMRCo1SJvh07DYcGIqOX3xSrCiZA2HEvBS1TP75+2RhYFaE4
oLHdya/5pizOEy1kQ+EzWtEpkRXY+wiI2p3bRGaXC78EUfhva5u9yv5npOCf
0sCKbuTnwJ4W4hu9r4DyJ0a5ga9Oycv7BbaU55Vp6YTWAHuROCM8EYRE/UNK
NT9miIGinF8qCpNe79Zz4T06rWu2fhx7zDn2xaJCgGUnX8c49JGCBLgV2+Ad
6InXEDM/+Pcnd6nxymhhS32L0mUngg/23gNNUaauFvnaY1+kYlEgbRx0RfYx
N8ESOw12XbTfYEIE0xc2VWVEUj3mGgundraexJ5fpVSKipGGgOYbtMDdAcnI
jcIE6hUD8og9a6bx0gX1n9dFn1mF+KMlMnL8MB+65Dy0s7k59nN8MorsVzgo
hLkDOFRArbg1SlGM5v1O8YRs/Js45Fo3vgSfF/1x0HgJXRueYL0JEkxlctZ/
B8Ov2RO6aTMp+Uqc26lu5qSLpxHBcGkrE56aAToCoZAjc6/NMVMnJ3kWGqP1
h0ofIUL0BLiW/r+EGoCeDfZ+L0eTH5Zz0zvp5r9AXJ4x1pW9IuIA9CsXciL9
FcDUVAIFeC4k5XzhNUb0U8f8l0i9O6xQbHbgL8o49kd3mjLLfM5pYd2vEbr6
aWsKMFFPciEwhOd43aMotvf+1fmMogHbF6sHjXB7Nw/XIiCviYOfOKbx7Fxh
XMyq7HK17WQNfneh6MM/zKG+wZFv/6mpII1INmV/E5d7oTfg8639mIKt6pL1
g74Nhf/+o7Dtqe+FBvKkZB9IrkSruZEnPS2pu7qUGRAbcgdUofTPgNaFdz1X
rSEgW3Bii8Bf20+p62lKaMLGr7fMimLr0n/K9cK0kd4hu8y0jvzfRRJq6LNr
8itDh3YCDbIGSnQ6lWLbWOmMwnE2V9CHiPoegit2Uo1Hbb7eM5B43aeA45Rc
nIb1QwNX8LnZ9CAfcqqxlBfJEDzgD3akqky/qvWbCoxxdbB9wVnRVZGu0qgy
etIOC1pioZbtDzdxyk/l/RfQU7NhceU+eDt/1ZakkXkSIiNStxeIFJvP2wqk
B3cekudBb20VIkHb7k/lsOR3kUaCfdwzElJFFS7FHkrzkWhW5mBSJaoUZc/P
8ugl3BRlUHxaHmiBPLarDd9CEkDyierB6xxzgW3U1AdqTmXHRFqkJFSQA4QR
YAZU/cT6j1nB3hO/FIXOXXjSdV/4V1TeLl4KUotBtZHkgVRqreobS7DhSqwc
svLg/Ngnl5kj4tsN28IuT7DR5jnKUMkbEiSdyP8S1f/7IrlJgHo2V6CHK7xn
2e1nJXyJ1ABxs63N89EXnaT24s023QWt1WfWHn1e/a+7WrW/X6kDtyu9gHFt
rfy4A+pb7QL7CZIFs/owCW4qegnqKJ3NizS+Zr3L7JhhFOl64MgDEhBzkhXj
NPrvloC+7penozJGDHbz1alQni+YpnLp8uOTECiQCmEPvJ9dT1K2vcMUq7Oy
Qv3ARHBgGhi9ey0XnazHhvISblxqfV3Ea/0qEPh6rGVfD3YcC8mARHnSnFQP
vYs90EVQH4UAr6hbVLoIYnWd+Rg8uxd5SAalxvJMqt3zWSUdAZlK3B9tN1Cf
J/kUOIjAONFjCaKxHR2izGqOztzl629sxTgyX54Nk3Rg5Mmj43rfhBhyQXN2
9eGu+J+ql9/hQwJFQnpnyrDRKIV6zJAXZZ5S3mGFBO2MVltNcB8ZQh9sPhZS
bYTpD1zCbZ0C1a74W5snKx6WU2q9qFjQOsFjpPqpoTcxeyIut3GoXVygmpA7
/oF/S1tIOcFXyx2Aza76CqTBjHOoqarP/xUSPMBGcQlPP3sEdTsB9oeeeA9s
gITe8uNAVsaffbFa61mky5qPUNInvm8bUFqAmTlfyL9lxJXrOCaqPxf2HK4y
z19E54KRm2dd44lc7RgwzFi/bjnC3belJ+bSUVSl4FMX6Z7LdMwwyiBzwAF1
brlyFAxCIn76AZWgIkJCWW7I5U7+lNEl4al9FidEhCTuEFHBaWdRzbBUzdGq
Wi2nKlwnpsCAk05/wGB/Ulw9YgrTFb1IT9Q6pTEIjmSwzEzB5YnJNDiZCVO+
7VI+6PQgwuuRCj6pgZhHoRfHvzi/G2W+Od/Bkd+k8skELmIjzx9A1oCCESEq
Jn1IrDHXj60fqlQ9dSQKUs4ylFMasI6zFFI2dXIS9wrkHonIujJ2N7rSMugu
jMQGJCbfiNnB0fIFmXcRIDpJG88wjAx3t6d/6+bv6TIPUQKriVUBmHURzM99
C3fDc0cOP5pVID/V8+oaxnOrQArqldjWDsvOv7VbWr1xUC8UA/FTkXrfrv4N
HPcPjlbnySwwRo6uxV00fIjPGCUSJ7bKJKq1Mh2vEwnm3wztD2KTJxh0GBFx
/anfKJaMLjGhUMNBu10Zm+BQwbC2NvVj6uvDB0OcIBIk4zNfEMErHHRVVrto
yROZxY7I/2o9EMfshwW0JxHbJmF3+8/UBCm+cdTQcAcpSwaHdOoZBHcbvkba
kBOHFXr5CutmuxXRI4oTi7XhJFsrOW87pPlB9pgOD/F2f1tN3p2uZ0YgfWwE
yX20LH//50PaPlJe6wyZbW918eFK6SZRbahdDq819+qxTfQjzo7xK5NEKbSw
f9sqW3RA42E0mWa6/I23IbLCYKBF0/IYQ9oLZIH3YbICtFgk7MIRKTWQM2fv
NOWnGyUI2Jh1geekMYv9iMQRzjuEW0/B0a9km4QBe5Gn3CaYMsGotWzWHnkm
qJ+1jf7xRIhG3Qz1dXYWl7oyYY3Qqez1Z+3T4dmy5t4nDdg4K3o9QFZ3SxMN
1UwLUOK2Ra8VksqpKY9B4KByqCiKf+lwGT2pj3FkjZtNCESFb6S/uvukojHs
eVtjmhW6Nv6lD5flXceHvTqY4keqsZfg1FHvw2I5WXVC1Jw2oMzcny5H3JvV
TZbU234AikcVvDLwe1LQa/AX05OSD0mqnSrqyWF2MsHXKR6PzpxW2Fblt0Ok
//Pq4thKx+XR9E72c+Zbu4dmP9D63ooztj/fra5SCp9c+ONgVBCRbhjLQNrb
LhDMQ7+VgxbuoAzelPdZdW13tSIbwHBf3KZl/pXyTqSr9a1NIEneEVbqWFq/
Dc04JHlGdO8EGxCJDOPXeO9KXQNSfc9QkZSxawT5QRR8NpyFdIFlP3BYYSBn
rgVLXODYSuMY9mngohHrbDbH0uYbNGrRPesgFU2KUCNtYYvys4obFncXHwTB
ORQRvOxR2yjdYVA/UAS7bTPHkX4HJh8Zk3aXGr7GjElvtinY2G/rd1NSRzc2
gAZIKL+TebOfPWzA8d1Z+BKe17f9je8QRRWFmNXMsJtFChJcfJMj3rq9YM4+
5OV2wrEhNpHa1u7ydrSp2gs8XEfwK5s7wjTPYYNL2tfwLPHU8ylFLuK6Rlxr
3QbaMidyCOp22ja7RlFbYJh3m3gmNo810u8LZVnNStvvt+gGwBQ4gP7agrE+
UGuKSdiw6X9j7g4V7mvPo8nrAZWX8huTfRKfOX6IxlRWIfYbEL72b1evJg85
mx9TRlNlsq/rSWdwWg1gtXLRaYfEl3cWA7WWvBBQnsBn5eYl/BJcMB8xlX9G
wKI7su10T2PgfYmViDQjCVPXUJOPa2w3K5Y74SWuPJvQOresSQr/w4466Ka7
JFklLA8w5ZapPysnIxLgLjXWKHOR+9zs6IEcAtyCFQIIEw277u5h6rl3Ghwc
7JhBMFMy/g+deUtZR7WK0nmFROTa9KioJjKIawKpPqDCZ/fnvYq5mYxK6OBN
zxO14Nv+F0AWV0Dlm77QUcx9UODFsqLiFOe/1nLcChfFnm3Ere9x4kKRjTRR
ax6Erzm1BY/rjEjay7/U+xhDezo+8/fOgjy0W8ZDdjmjh5BAitXmb4NlxIEv
5zyZ66HZLfG3iYVbEvoexcLFRyBxfDBiDEfEgYG3cqrbC9dr07LsQIlqZfjC
pPSmFLGCnw3xB/y4IpfdgL2IFVyAHFeZtqYKEgNXb1lwsldF3W/njXuzk/7/
5LHMSrY6e7iv1SUpVOCoW887l8t5ifExcI9WVU6/gFd2SmkApJX4RiDvcXnd
oQnMUwr8S12/gJEDz+B6PNIEZVeCi2hG+0ac+pVi2CsOVPZQMjKnrl+co7AQ
pDH58s3J1+CY6PukJVlXfYuOGK3buE7fxJqFpEL2YKmhDZ5IDmmJkB1P2nRI
7v9MTvpuzDUEKx/mBMbc4u/HlG2BfnI3rPkPL+ewWHA+QF35WS3E+W7mxTyg
xdsneAu97+4V9Dhj5dHI7bVxXxFJP60RTI5kAiZbGihiidrBn7LQO7YSztGR
IqwsiBOTIG2epzvWwNFJDN12b7WUzQMJOB0bhkToy7iGHBzTc4FSkVD6hoCj
Uqg3AYzqYOm2KU8C5N9BtB9Hz0K3thy/uopPhTbBtheGX+8EyRKbhk+Ks/oA
7pTgP3qCu37N37MilIeTJx2HxS6sJBsISXgFjd1OHgEAEfw57SBtqo9G1Vet
hAX+Ceek39wXybaU9Dsb6hWXQJVmc1wLq0IxtPMEaUomZV0xizquFjaBuvUR
QVXeBetJC/102S1cJHbhS6YTo5BdACXqLPFSk8UuJ+/InpZR6GQOmFI+5D6M
/ZnxzJA5d8qnhPQF27RJhHv+UM6XRI7hIALyzsmq/VsIAkPMZoyUcNvwBqZ7
fVXSXvstGds8mvEvNQz1UqYj6BWf3Kw2ZxgIHJdDNkNxZf1GK9a0FgZRicCE
BoVhMRd6h+iSG18AFGtgl52NkocyVO7X0mYWd+L3o9TgW8NQELSBMZai6Opu
PEimPfkLOKfQslQGXyPjNsNgHjhLE+99UqsviNwFZXW/QVf3ce4L0edB/8Qu
zO0XiqEZAz3j5dC0WnNtMhGssBk/FWJxCZ5EBSjVSwxdP19r+m/0KijzO94L
gT3XaIMPzt809zZM1zIdgBm+HU8paXi2YSAdZhcB56zi/2OGHvbLT3i3cK/p
jHzSYubboeVyCnzaDIsMb293WHQ7mApaQO7xNWINt2x6ptArtlOrG8rDkoIe
A3gc+yk2PQ8SPQeHEf25c5iqZLjoIBnOSIkBUfmsBH+KoWpMDbnrf91FABzd
9Uch8xbOlc2u4PblmomrcshKQuyn0jkM3sHAtWhpmtKsVtbvPXmLoMaJd6lU
WRpl6eP4Gbpw15OE/H71cfiVcB2YiqORkiTvdzIfcFzHkR/MwaU4g/B8EgAl
Pgv1u3DY6KWyKO5W9sVcExXwIL5kAOUwC5UVSqTUGyt9AB5EPs37yiwqTlwJ
iKS6pCGQiz/Xr/JUqIAylbNKBhOMlsZLaetZ54cW7E6G8J3XbaNitDd5eQXd
xYR90XCPxCAa6mluSe4SDqiyuxRjplA2WuC9bQ2eLWyN/AY4VQwU1cQMogGQ
Nx6j3DlqWYfUQgioWwmZ2aKTCfEYlK6wwH0NpTlsSOIKog1YPKSEMPvI3HlS
nrJA26ClirQlpitEreICpAw70djsvZ96keZ+/pR+wkv325JjuZ93xVIOXFeF
v4mhpENP3qC7zJwXq5KZA7Udt8JmYj8hB53PnWK05MHZAz3tFTdKCAZVHjB0
kyGBH0xzHZ0uihDvbrPX9cTSIZyt6xXc0C34WlWTuusKLzLhibTVWvGlwYNB
lK5js67prIAGE6R48E5ymOH8e+Jb8aFsg2puBb7H1DJE8kADJ9d37NRksDLq
nyF3cgOATp0+GnyQSkstT8SgLlv16EVHV5GUoMDIywgUv3t445yz+Hrl1iur
IrxcGm2sCWKoX+TvKO5TK88TOIAo+E9IxJeIRxCKwFnAerOVkvfxZ4mo4PTK
cWHgHFqXBWXqeLMpeAyi7Qdb8K+Pm7Ly8XX2r3cnRIgq9futaSI+g6E6OuI3
p/oTAVrsgHbNAYLjVoux4TxNmktIvT0Y9jfYbjTLOs/khDw5aI94JzAoyJ/s
fKdzcHmXrCiX3saNIrvtPiRNPbTP8BbN2VW7wtdgWsNORfFvsQ/XbKJuOpj6
mx2S7UsR+Zys5udfbEt7v67WQguQJgCywJRiRPzMhQRry5sAt2DocMbx1+ts
WpY3YZNbrHDMWA2FVoe/Q2GiMJNUw3O2t70kpUHcG6WlKG1RTya3aqJCyMLg
cEjDgq3UwDytMQruLJMt6Vr7aSvcUNyXER0/2O9svTBxqp/kA93rtfmnONMq
fAocDPehR1MIFyFsrZjaBhL+8TrGOwgh7MklmPxX8xazGYqdZdkDN/PdRnus
mDCRfmE230CSzzwAyxYBQYXtiw0j9XzmfaZ+AQOfjGJC939k1fWk84xNEOOE
iGWIfZLH5vrAEAX1zBjM3srgxL9FfekNyiCZhnLNNs/44KhVWX4XvEwHocur
eBaQsbp31cQYhDHXXLFx6HyQCopsFqDZ8deJHxOxAVUt1nml31wKw7bF6pfx
ZVgulOh7Enx96p+/KMP7v8Rzn+R3mFltzt4LrOmaBzpU/ZDx4sFtlVTckl00
yaVXj946RoIs6k7VBB/07Q5hL30Zz9eTAASTyMhoQojvgSsS156GnSN0VLKn
JpcF4HEbnMyxy1dA71UDubuj2UkdGGie3RyD8xMk3mgPiKIaHtE0Rf2Q495z
Pjq4rq+NyF29My1WWUsywwjTqRC4OHC4t20TGT1AtNPZM8KiLzq1h7nYVhuk
JInQH+v1TLa3G2VsUObaz1cvtpwkcyF3vw5RZClBvkEzbSeXuIOxL0CpFJ5C
v08qzQsNRG8lqRI+ElzQNj8sTN6ToPkhGvNqTEXP5Pt1PqjOvaerNP54qf0f
kG/W9Q5PMdxHUZe3q/oUazluja5GFoRe3mr4WFh7OJH+r8tL7vg0xQGnl/nZ
QziQZqoY61b+TMFGKF57LNnn5AdBMzdmJtnFguIZjfE8HFF+fbvkYxBZz324
14xWEdfwGMdBzYWKKCn491BrAj9Jd/a/ERN0vlQuAkxxQIPpSPpXEK+i/r/E
0fK4czZGZowmUSqk+KykPOuVrsxgTd/EwaAjzvwBkAzDNPQDlP7k94eYiwNh
r5F34St89jsGvcRAX4wO4Eschr7bJFI0QdLhvVQBrU1lsSkoo1HLBGxWjaoe
KSaDow0aOJq6gsIB4YV0WyIZWFdw4zhVxzpCX5RdmtI0jLVh8qTKjzGiX/UK
USrRoDcFAh/nEpzJ39qthhGdF0UM+zpwfpG+Jz08RGCYjqh8Yo9KKW4Ixz0W
pyxkq2DVYwjtOCfoF0wkJxoy1fs/rqvPjkAS+PhX0RmEdZlKbkZh0uUU9irr
Em10dB/LASBopteB1Bktky5rmSCgkgdg7u4/AR4WqjxB9lS6qR2D8SDknHCk
xuZWMXhFT108mq+gLk7+CJ6rhoxdeYcUkKS3waXa38YpcGpCLELD3jHQq1EM
MAxTuP3ot7bjUM/4OnIFV4jnelJX3hUv5592eIfW5ZzazVmxDSMQEZNcyX2B
9AX8jQPka98+kWJhrvnyf+UZvnz4MfCoOKmzleNUtkp5KeZtgvXqJYA03yGN
23U6yC/tR/PnR1+g6xU4dfgxKV79MoSL60n1Hb6WIVu7K1aq5/jFXVh3prw+
uK4pUkKEq3fQcuaC54pUO3HGgPRLEcpn3seRr5Vx/ONwgSW2OT3UVp3EPqAI
NnXTEJOdnZCF5scgWgqgIITYl0IAOY82M9BTiNOQKids2WDfz1QmQJIB5lnm
IYR+Ndc+wjURk4grx9z62BeaVWYugM9cF31TylDnIb0GGqndfAtP5bhe1Chm
xG0JFmFSP69Wdcbb/2Hk9ryUuHuSXcxGiepBs10EAB+aaUUAmzVuKEEX0icn
G1gMw+a6Yh32BtBMg1UqBmbAa9st1w2NihxDJSbPZ8pvaNte5mbRsjEyiCPJ
iZpm49Ggm9ULiNqWpFpYWVTzs3ngLgoZleKDFHUaBXGENJa4gXRqF+NH9h+H
asEXecnGOe5+T6PkB7tmlpceLtYFHYB+2/Wpm8S8Q57yR2vNzMa0HFR+sxIK
lmndBddLeisB/irjgSIpOW/V5f3MrPPNIaOu2cYi1ueng5ucNz5SlpL1Bd8Z
HRmjc2N52x5/OnWzRfOzJDI4ylrbx1UijwIRNcgO6wum5svb50UBNF1CWc94
Po6u86wLIXApRzFcLUlrl/C98rSiLQcw43gWxJbExPDdaxj88/WhEfmppXCO
MNiPZe6IE/FiQK/FrrvHfRwcMV+TZ0xP8guEnorg58chjY8Y2qGhpStk53tK
6bOHr0RHNfQj58aKvUz8gmQWo2vY3lOGqTQAwQI8ImlcPvLtRBPDZSJG2Zq6
SV2fOtI9E/1PtgBZ6ONtF3NuZMMX+CWfvQ4G9EaAA+UilLHpS6JShlh/rIjK
kWi8z9kFFt1H/2aXCdCl3AnabV3lKEA9bmoGcJ7/GQj96viD++/r0JKxOXID
cXs2JzumF3QSlRO0uEGSO7H1bEx73NNQKgvl8xG7cP9MUHyOuBnmWwUWm0sy
eLV4jr3mB121fVR1GTidT5RFSrbAIT5SUoEppHFePUsTbPyoKmmWMGr0HISp
cb104hg8ShTWSFMBH4cymG+skq6r8DU34dgwQiB0i33WhRG/drAihDjn3iXe
KFjG5xJQm6hJnMp8UD7cnA80aGLUOzfGVQOnsppwd8Pw+JxOkbdhnaTQgbH3
itxtDSGRQkDJClEaU/r+3e2UyCYnEhT++RMAoiDxvmRwH1YntIYWz1zKwevQ
YKvqNXxzPuTEcTTDjYIGL+YgHR/IQRVsS5Gt05b+uE/wIPCD0veBbxgY+tXg
XSGkfA1r09SfQOZXEo6HX0D0cakCDv9On6ikzVHIoPwR3+oyX2fC9cEk9k2V
5wn51FYCMhhN8PBdUD/o6FOCckjEPiDUs3grdKfT0AMFP3D4s4YDvrC8OpeT
lhk1vbGizKjRR4GHpCFAaswzQDNzLTggI1KIDQBRokcYjukC/Riy5IN1nlQF
fhxyTPH/FFl0VAL+2O9hVAGdVzuHtD+KKH4Vb1erAOsE3eE6qJ38L1Fjz+Df
QUk/4dGZ8v62KaMvvV2hRL/ZCMJJljRd5y5OvjLiLID+U3uwSHxJ2Gq6rpFZ
HIGZDTLheRwC1kK76htdfUAgiH8VnGz7HqawzrJAnmiheEVMsloe4IIiCqOK
lofAHhdakvka1sdh8Tz60W9CWSyL+s/pBcc8SvW2H654qxDlV2SyJb8vA9ez
cV1pVsZ6T71jQ/lf1BmQWXi7YthZvoRVW41AIrQHZZjVf308o7gqPeMiRl/s
CZL2zfMcGP27NAPdU0OsmZK6lz2MQkVlPYdmLGVa+5UFO6dFKnFCZGIVut60
dNDB3YCleh+E7B1LygJQVFWQtZEVwLZKcOSjmQG5M02x85vDl5h7PsUsx7sq
N79dn9uWnXdw3/TmO3v8zG62ui6hAiyL4XHGThXejN4ykhqWe2KQ4D9l2yxW
K0+8XYNhUSZpPs/wJv3jMzNQjv9hcqj6X++XT7DKP9+x/UBx88EEdadqzwLX
7q93LjppofKK+bq3W74EVAIvyQzVJEpJb6+YMVedm9ODbDr9xd4Xrqe6Xc/X
TvjRJZ4uzDFAIYj1hmnEivfI0Dr4LFv2lDBOh9yAYNdgu0cjadgYmkvZWL8p
STkPqsF9Dvkv1VKTrnB4nhFwywGnFcBlDvQM3nYx0mPOzhR1i217h7ls4Qb8
YuQIUINjeSRFVWWFmDpA4HftweVvVFQEId94/ZZnRN4Gv5cyr9z6I6V6uENy
VxetM2Xtv7Ae/3hlleixX7tsYhaf4AW8OUjG6Tvj6hem/hoveI+dLVIg4Eza
YL3EFrPnuM5uTL+omvHPxdT880IowImFu64u5YDGXFJbK/K4+pF7udjITaM4
gm0rPjNv4mZMd7TApzxNX6kW9hrxS1dyGUV34ud58rLSo8vPKJSKGHgcZwpL
acfZ6qO1hFy9Bn54abN59GrE9/s7MDL2RH7HEmxgsPXevIWeQNv/spW87aIL
R4j97c2VD3xFVL1p/uveWZewt3Yzwl4qxrWO2C7rkQdYhyX92zPJ9uFiJuDX
D74Hx7a4O1RbXzXW1RvAC/7dRgn7knVffY9S+F2Gl9h1q2WQrG+OdfHtV1FD
aRWupHxOzVTyTfnowIDYvstQKEaSbiWGXVsQQRU16Dz9LJvJ9t1C6dq1mpYH
sd1OLKftl5OTVUamjVftOlq3YpXhW6ZnnsTdS3BI/f40gckZsmovzjXKfLqD
5nAfN054xJhH2cZNOqlfSCZzZftFbWeU6qRxALJWZeXK6gVtxOCXI1+/Q4fr
FF8xAIbQYx12F71l0BRSvdbEQvA2SnYmEe9WK68O5gAL5cZohZlNhEkERjW9
83boqCiDI27VwBxvs3C91ycLQMzhfG0birvBgScp0bAkFOWXG7iSftk346vs
7LRq38JgynEGcswl1xkdwYsh/EgDWhRz0vMZ6Qqlyz2bYBjbUGj6XE2AmwkS
RgqoCqJwrmLDevolUk4VGd89akfsGEczgrmwVtj/1AbUv7cm84gd0/wiIJkG
BlMdzrbVeQ4UXiSJrl1OsrUDlXe6aFLqAZFdY6T6VqzP/ACN6Id1D109JGjr
U/HW3KL5GHAZTP+6AjyfvQA3RoWRfb0tWequ9tUvbAV52/06YQwFLRqzxzC4
122JAdGchDz5SPbbBP3jXIRgrHokh7JYnOoahOZEPcAgbhdtfhsr94/bLumE
6daZj8enqNXHDm62yqXN5pfOzgHBninSHBh8o8NTnhwxpn/qsmXdiDK1yWvG
zWd2v0HUvHfZNgTZTTZL44MMQnuR4oMMQAdde6LIE6qqf6hDqFQ5SRanyeJJ
MDormqJq2D1lB6gSYBxs+MP7vyAs4wOcIaW7QbkqXmxsUMxOZQ+Z8yMNaCOk
6zxaJtrslzGGRTevlPBVUVNVQvBwKCxC/KFBtK5pq8N7DRFywWREg2I4+YRW
pAptZzPX0sl3JKdZUV6dan2JjRumAjCXBIBIUa86k/wOecqcLo2CHBxrswzr
Ian0qjmobKPvUABD7kpr0Kx9ner3uP9SouFEyh1FhaWwC4gOlQ2OHfOjMmRA
bL5y4FAMGCRB2zFaE3WHY/t4m7pxEMhYuHyTDAWDBMVeFQzfeQjrP7lhKIH9
C9QmopaXsWy9xpOJwZf0HLLCO/zr5HX5tnx8BWeGSOD59zJBX2ckRWo/KdAD
D/OmRqz6Kwv0d6hUuliNEQzfAa4zRN/8qCzTLjJvI69mSBnkUcPB550jPASq
DrAhvZabUhEwcefkrXs9gk5E/vGbBe0ykqb/KMQ7SdwA0CpmuxrmlRyo/mOG
DgVH17f6tcrO4+WmWRqfOUKmll34oYoCApQCt/S+Rhv0VUhUtGh0wapxT92w
SFkjRqmzy7zZwVmFs17cZT5avboXPdUHDvZqNug1X5VbKGhrQl+16oUPJGJ+
1tFeuhMK5871fcR5y3NNUVNlJ0VNcy9xUO1pMOV0ojyTybWl9F2RwiUjnwkz
FVzNXY1iIFjyM7gSltZ5kF8Qg5zWZUTTtvNW2wB7buSv002Uu2Fq2NQBNSCY
XGO1dmsfPPVjQcCpuEpEP2F6VSmHAgkZzlnzsNA7xyUViiGRyAzQd1QgOgcL
gSazrI/9Qeh+7ApBcxwukjuwx4M5kk+B5SbBe23daX4HVHvCQlMYUXgm09Ms
lFFlhH5R/P+lAyqAQ55I6fmaUOQV9iw11lXlBEogaFKuQ1O9D157zr1vYeAB
a3M8SpfC0mpmkSS1Wi+dEtu9dexDoo4DVHNIX2+OpbIcodCBxsHJI6ML0H/d
F4+Zb7D+o0mw1ontVpcdTTEt0LBoo/0ViKzaH9Veej1sdjvDLR4pZWAwx/Mx
q6x1EQRWdFIwl7OFWNKyWctSOBTnCPqBXdzfgGFHikDdeYuM0mluI8HcQskN
Zf/JQIj+DsEyb5OG9shw4avdut5rZSct7hxCmOyOWI13O7fuPBoWJNiEvmqg
V8Xml/R4Kw9/3iAIvJfdqg1KjxmAvOCwYuEPvIRos1Pwp5xLo3199V2RbeTU
pGFgaTPRCDJ/kBXLRyhTglcRYNCZwdcmCyiwhZr+JrL6TosqNYDNHvoHqdxD
m14MbXkfmOmR2uZplFRDOIaHn++AnleEXZtU9cb1j41fZv9tpNAVf3ksLO9X
kwHRj8J5rxoCcDimqRFLfZ4esXPyQQ4+hxU31RUNQdIWGnmciv7sxmJcO9nt
LQ25NevLPHeXnPCGP8ktsD5FFG73xaQsaXOxd5lvZZJYGlURCP9QRWcwhHPs
X8AIkpMhFMwWXYNQ0AKCWrj6ikH94rIV1Hf7Vgw9vex87ma1qrmUPRl5DYt0
ewYRpLFcFl0lxN43F7lA2kI7tI74w8VomLklrhrPlhkVIM8KuSkbKiFCQTOI
f37fnfr83eEiGJYYP/8P/9p7uQuibOVnUOT4hBX6zwvQdhkZfZZvTecoSr1z
Gxs2PoMfU4jjprLCER6kCRWiFMeTV3DovmaCH6xYug1dgP8llNqwb6YlxN4t
MiY6cLeZkc9XYNsS8t4gn4eWnLQjAv+n1Rz4Fw12Pq6M64pmDLMAi+tE/x1f
dUuNtuoy5y+EkURGK0PHt/RzqmP6esU6z3Vee2oKupw8D4C+gmpCcfZZ2dVg
FfotLMEZigzBzGRQXZIihg2PXJfPondI2X98nWnWWtcIH95KK1JeP78lUpjF
IxfWAmqFF80eJdyge3YTvmVCapPfZrxb0amZXrwjrsK7Ztocdofv0Dyr0XEv
uN9Do+Mkp3pLE96LS+yWUZ0HyPQ2ukQHWtbPVUPJm1ba1RDzt+PIUwvNs8lY
nOUyVlC8Z7XDJUtFe7NiEKHD+uNLIvbXAv89lVGSA/K2olq9oBiZmNgTdPqy
HZGKLd14ZdIS9msW/WbW060Twm1R3i8dEX2Zu8eqcsuWeGBWAE5vmyYNq0vM
XrajT7exFaEctEAs5suDLNsn5nCemV42LxLgB6bM82J8sBDyLka7zsYnOT/f
irifVOHy4jC265GVSftVsRXZoBTU91HiGqQQTxenP2ZgWHvT9zDNMFU7jXeY
yr29WiSMFvk/kWqS2wAU+7aSZ+Li9LLsq7muA1U6y+rtySiSt3OlmnYJqKd3
cGWPcLbU79OJumA3qlbo4BEBe4fcD713q8eKmP2glHI5WFFLqCzPl92vLMQc
YN8famdC/FL7yG30+hAu86VWhl/cjpGKwJwQ+/SVzR6+8NnagXD2y4V0WLE/
tzOd8dfgq4nmtjvuDmIw3APdvEmiO+SFrl2wMoG2r/OIn2jUL50NWLpeFFsz
zsPxBVUldP2KhZ62yhAD8MCP6z6PcC6tO4LROzYCMBr2o1FdBdLxh2728txw
L46mcB54CyGe5VucrvkXBt2JT53gycfCx2DitrTEGmyhfz7wMRLFaI/WfzPQ
koPMYrPMnwtxXKaU17eNQ2QbHde6dr1aeARiINCe20uQ9hEP+SLR1WyRUJUV
pIQkf06b9WF6d/K6tjZlGxx1gz5AR0uLdFN8hW+IgWiHeEF8qGC1WNJ5doCF
pQrRobbz/eIQu+AgtSTJK96lQcfTQTDykfGV4cG4PUCbbY4GbT0sSD5zD8F0
XBhpxPX/rIUCjxjKvR/++tWTVHvzOqtLT+tXcvEsjPu1PrR82/MaJXovlWZl
cVnb0d6dSXTBlDSviuGTgIfQuHCiVOMmk5YCW3AV8oSoN+Yqm/coZovinSlf
TOu6d6qs0pJ3jzwxpHY/uwrQJnprDCCCzVaNV3sems/NiFjdoJzwG8yt1Hlq
LN9KzP+zxeAO72ORASUaKXtPODHZ18NI354MGEv9xkmQp1yeBmrYacwlt9P1
TAvxSDtmZgQTfuz2oUic2OS52EldWhCFFmOpRQC516/HPlbL1KTrdY1wCU86
omsXV+PdFIFJADu4LJPkUbNpkfq+0O0MvafoqmZ1Dz7mf/y35uXIrE0sB8lT
1eBP8DRr8XbXF/egP4NODv/J21eGx33sMWLROTwjSgs975hzASq4/pNCutV5
jz6U4zjiXl74bX+CIwtmdMzBed1BnEKPkWNolfesfIBLuhsINBsCJqUbFVOZ
SVvWXOpvJaVsMS4V1TG4FrQi47hycGHK3F65vWRfrhIvsFxBLcMglOMkB9b8
qeth1JYpBUxSPJHWD5NfaypzHgn5jVLLkVXP+ZsMIbZLs31PHQ4yyHYANYBp
loWwWPVVwvBKqovNCV8yfaX1VN8DCjvC+0vch3Jwj+KV8v5eHZAepMeGQeB2
bCHTmdxApWp/7xVfraEzQGe9DKBqUBDxiNu0Fx/cc5v9EJTpVVDtJX5nws/C
18/7LIFWel1lBRi83oAVtuXWo5IGiDgXa38YDub8K2AoZYbZ7Z0x8H4z8XGT
q7jaN4CgtnJ2Tl9MSop+e0D12hVZWiwaIJ8ZM1tzkpvj/UOp1Mi3vjdyvS8b
OXr9BODsjiL/fkpFJj9ztn0oLCQ5u6HgyD+8Ihu4+5Vr/INpTT1TM04GGFbh
FECh9osV2DRbnT6vLFgOKSHQ7Y5JqZO/zwbCh8+1EcDilP16qfOBWQjKhOIx
M6sbYGEeuggg6+xU+gl0O9ba7V8BDvs2JYhip7JnWfd6pDXnQDRSGSY1tH/b
HTjddv/iIw1g+9NO1WNU/X6PpfXDtpz+2wLdcVkgKrPt7Al3NNEu9FVi+Llz
9xv6LLyR5s/55KPymltgaGgT5QpHKC5v9h/AUlQBWN4Vz5e5+d2WmmrALEJQ
l14gghUCpswLKxKN/S6p5fozeZqfl6+1cCFjcmxsTtwg0kzKZ0m/LGAK3flV
8KkMNAW8dCLhomSoQCxcU+zlsyEIxToHT3s6Yk4neTffPW+Vs73X3A0NOhqN
NWkymsdn1t54lfv3qGERv7T7NDsiCaYFF+GMaEXZjzsBthq0AwFOWFYHRrll
8JN2jwvw/uwwQattC4pRx/rBguE4rLY6i8Z0Wu5D/sBP2wZGHcY//L1eqVWp
HRK/LM3kotGhu6bZ0KiVd4F13/8pjVf/teqh1WvmcMLUa9i2JIgjXozGGv3U
+tWjiT8JHoI6vVnfXSz5Gy9jd6RNgGeytsH153IAC3AGgrKMhVc2ALzW7dyb
cKKSDSv9MBY5GWpfqFM36MrEEctG1wE+GKGJX5aCoL+ryTn8FuP9wYz/Xf+d
xWmvskHJgDo1f/pvWpFETl3sjAitMphdj2wTynwvggVkBfSuRFevDJcht1UM
CCJmncwQq85sco/Z1vD/339jxPyIOoTkklf9kjE42Jv88+zO758xnyG5ZuKO
ZgLYa8VOv+Y4RTZa8cgJLe3A2cfd901B3tGuII7/7GUK2VAeVACcVM4TLS/0
K6nFMWzFoGKZnRfZZORPXHZXuwH6lAy06lcCaMV3gDUEt7BJLGTBnHi3++N7
GwJ/zCWfgIjVl3QITANq2ORT7pCozWx05z+ehnfLgEXOg/9YeNJXIQ6cSb0T
2vZEpo6qO1gusAuYc+FXuQkyud68YzczOzH1kAH8jGditf3VPp2JRO/Cw+jM
o/1I4t/sF3vzLkAxPe0QpcDOky8Vvpu6wjPPx58fMSwCTHdqClNkQ/NgoH4G
KBrV6z6V9tK8u0tifli5B0bTEaQqP6ISA7T4/m0Ip+H86G5GwFph0vGF4011
CGA/Zp8aDnZLx68mXsU5NdO2vE5nm2xkLUuA5iB7mlvV0W07itE4IqWNYla1
/Uw3ia4cT42mVAa9Ymq/Nav3Y7wOJAu7o+SNWa8bT1ZF1Wz4hmw8STfNvIJq
bDWBScJPG/7m5mH1FEllcS9KV5eEQyuYyY3DvB2yKHzDUZVGqb5NhiHEXYN1
8Nn3IVmwjpKWSST+rxyIky679E19Wlfzbi8vmNw9zwPruQkiLnXmnIO9DJOu
XxDc1Nl8M7bW72Q6KgFnnOe4U/AyGftSv36O1q3cPXAwvRnEnkW+mnVosaQT
whQ7/FWXeA+WN7nyd17lJXAEP/CnvUfedDQ+cZq3877MVzcjNvmyEbadmWWo
zFo9cTcZiBLRgYcOdicD0pJpX/akXEW7/8RZHLfJkVQX96OcvoPRk8sUGvRy
2hMajggGM8gNiICIZX6i/Sdek781kVhb3RkrsEZ6gLpkV03NRGedrB7rJRV8
rIa7flDiSZ0Xv9EOsuZa9642pLSWXxXtEgUBKWQ6BFpD1cxd3p4muzw3TRqd
nyRftzNqc9Wb2eY0SVUDJ7LlNI9+GO9EXUDnZDON1eRgopeazIm+x128CuP/
tVRlXOYEWerJ1lJnfMltHTcOgrlIB/VkoYL+/NOeqnFVDT4cBsVWuLTLpNut
1b955YFtzL9iiH2IUpHyIExkbJ186IeU4uXVTFsC5AehW2Q8PTSbug5oWVh0
kunvqwgMHlOwdIxq3+e/EfudA29bYudeZ0bfVpSJw54Fa+0jYwf76SW1cXe4
GdlhwlSo4sYua6gxfMuC0u/1ts6vOKjQYdMdj/Je9CvZjgHBaExSNrXsJO+Y
kdMX9bIUin8Ho/7Duo0lwOuFb0ddZvPdGte0Udz2kWilj/5shucS47HKYWWH
3JtXryBzbc4witVqxwhDEnuAyiSHDcZnhMdKSDyn5cR2VFqKlqVsPBWDQgUj
n7Xqh1NtPKAt28uwEPJnWwP8ubSLJRqW9pe/ZhH3SoiMZwM0WDCfaPkrme1d
7ZhaFVpFyZqy42PILheREcw+V+lyh5PDU79P5hEvI3GLPfyelswOZL4IMVq9
AwuozVLHOExC9izluBu74o2RQV9w4C36lCaD/pASDKed7dSd0ciqRo63l0Jj
sNxInqZL7YaHSobD00Met4DIcePVs0dDJImmNLlTa6qS6MRewHHOgc1itlJW
dTHwvBVhdfnWoBwrsjcEkU228xLOqaGOTPVLYY9+bK4r5yj6OdY21kHRjuFq
Kq8e2UZ7aildoRFAhRFrBkRYy1GKf/B2xx/PAXbgCCzPD6sWHd2ZFob0LniV
8iSE2W392ZOMhqVyHKhGCDCBugX4jrR0iX4xv2uEAyQCoEhFd9t0Ak5Y3jjv
7S27wehYUmt1FB7WkgfdC01eyusqyqCyLEptgb/DUsFQ48exi1I969Sqtdld
vGdsvhZY0ZgxL1cchg4/bH058s3odBk4RtbRfYmqGieGofkL1tFO7Cixy70K
Q6QrNzPZrDWuc98J9ZefTAYH8sTNAa5sr+iPq6XxDSTME7NfANB6iDwwSx0v
orvqo6eiU3w1H5tNrUoetY/2e5v09U5vgMYvbjqXplZqNFlTEHPDiyl3QlZD
J+KrwAt7TFQzAkpIJB3jP4IMWjNDkYApsqGzkswZIDMHo26i8xxuHZyjGkkO
wVol3cOFFQnz5VqCEUYV6nzgyppI/sruapKn9DHsoCBLEs8rWeo+O91xWdCo
9FujCUL91Eh8HJUGGYdJNKVMF/834vSEay5OjiD6IPZUzOFK5OVdkCwriX1b
6GBhppy9rP+Cm9ZUmWCoGywoPoaLKy6HXt262YARPCGKoH1EeR6mCUpYQSFj
YKPuHpV6JVGC9wTTYc4Pyuqx2oJHs8i7v55f4NbyHpPaxy6Crg2vY8y7IJKM
6BZNWzk76api8Pt5jIKSmumNfMBD7fJhecr49EhyFUs0/XBIYmFId+HOIHGY
SMKNjyWcqYqeGbhd6Uit8a5faMP9bGK8yK+nPhXBBNAPYpCBRSzPKNF5caU+
FfjB7GyVMrwZ0qdqiOclmKGf2ehDHPzRU8n3TU9XgzAml4naD4VpsfP6ma/T
Mi0BM2UbJxUVqk+mrlU+dH10Vx3xn9g0ZuinozFHX/ZlwcdUSFhyV7jXF3cr
y69bx7DEf2KIUHI3ICZox9K8cwNEWT3xqJsRX8pZxtfAb2HfQN7/KSkIieDY
O2VcsEK/bt3BMoFpohE0orDs1kPAQVP+Gmcwb2Yp/Chjftg8c/5F48aEQbGn
9uvfrgj87ctXX7sgDs1pZgNN3LZRBXe8BcPAO8SIqyufMOBtjfaleslA4vLd
/EahyB781DowXr8ZH3rNXtzq9TVIVY1sqXL6vSvKY1QujrWhjXF5KbZiCdjZ
0kn+E6M5ACPCLLjKsxl6nnC/6W+ibqEX9Is+OS9liouPorTNYvgH9PnRyKlE
mIaTnc/s4JxewGWDaRKqkYDMs1D9hxWNB6D97i4lX1x+o/H0Lsc+/pX4BwPW
Riv0f6z45zsmLs+fre/+poIcIjGvXgqSVKbgfeFbk3Y7U0ee2lkqmjxliZhd
J4LfpLq5Xx914hMRqf5gAIXqmM2NLRPOF+m5Mi/kFVV8CMTqY2e/V35NzO3l
1Jt3NL5ONKBKg80/bOgX36el4jaOZVGuk38N30tJniY42NN4DsyrIHm4z6jk
hQGyurLudEPqwPD3N2M1ZFvVmaTVYWyuWWZDEwuH9jRq46zT1oz//d4ChJy/
3cXDwu42rfMOgrw7yxIARuxhhMp20iUobCuXIVwaXH0hmLTADxWOvjUQuk5d
16qbcb6e90m1CnSgKgsrmnc89g1hhvS9AaA1lwUdb/zRFbRc5xQBKkFg55IC
M/tqbJ+7RjKvr8TmQTsV8u9pMkqDP11/3ICXujbtP76YW+Fxd3c9jyESxTXn
yQeZaQ7Qg6W4bB7QQwCjyRW8+9bnjW/FGLjLLhGsEeQom9TkvUnMWCNtkom2
KN3hRyK8MieSKE34U2dLJvKXXxL4D5iynRMf3faeZobxey1EeyaWNdDIN55M
hPXzh1Wv/hlIiGPlZKTLDOsvbeSZSWyjjpyQqM+bQP6knobPdGga87myRyDU
mN1xOTSR63NZlRb5MJfBHGn4VQ7KoCMnZC3orHCCa+ITcSoyGV5+ZZgYhEcS
B4uTX1mHZ6aiBjxkncnhGmOAqY7DEU+fFAxB/XyEU+qdnf/OO3UKwDQ5Wvh6
yXwxBS+kFks9wINMYV69QdwoHxKXi6phb01iZ9PLO3JKw+CPyz++StJDYaaW
t7vSqJjig/S+s9QVfAOd63qNnMRR/KmLzBRqgkVJkIKggNYb10MSzScDje+g
yVs2+Cp66WVJMVdwO9u8IVETMrXFatbJ6fSm0Lj+lpiqAIOkUQRDK+Mny95x
HRpnnRUmTBZ9AFUszjCsKJTpeRj5Ue+bnLjjJpWcgktfSqlMurlPW4Rnf0na
sA/rnbA9guypHcESjG6+wxY0j2rzNhmxiPTJxhS9PLouL2xY0x76dthZwUZh
1hs1QErn98GLZIxsPEFUgdU6HdviPp2GkxDsvjt4cUmtGChw7ulxUcry66bH
CiEJJy10GyGBG1L3nQdZ1qQ3NUH33MAalc2uyKL5TgkkIJR6rqZ32h8PxdsK
islD7QYk25dub4x3Is6VJCQ4LYyj/24sVnZ61YT3DDaHohzS8bsHLs0DRn2H
Gm3w6xn69udcRLEsEi+hxcitnUsQnK8gAV0LIkAEJCbkEWi6iKglrjKY3U7K
OfFNzt0CkeUTNBZEHyMbNdqLqdoNgk4orLa9xp/UaEl43M1IXRrQ2RMpc6ov
0v63slBXyATH3kUWQGHkPW8gqoHpda/N5D3P8ni1F3wttL8j8BnG05KUs/cB
KJRhYlIckZztDdxiGztbHaCseK40ONvAkK0fZAf2mc8ArB+yeuinP7rDhQz6
86GTPmxfr06jappvTe83avhVXkF+FQlr6hZsemGt+8DQ6YFIXo4KItJcJfvv
OI1HAJO1/hJHWvhG4kaSs0t69M6nmN6Y7hu38LayPpUIlYZ6GgjnyI3VA0+m
ZS3iescT+97kU1Z5AmVuiOTgSJN2q0Q8L/lU9pS/0I/LtjrdO24oiFfu5PBJ
Q8QpPAIyD/hsYjBFg5MgLBLB7D/2I73WBVNBuffQwR+oCHku57HtskR2DAND
zIFViJ/L8iMiZVja8NVqxJPBrZTm4An8IymRW+dF2RxHf4rL7GeI8Z0T3Ceu
YFvvSyob1RM4ziMzPMB3drPMS73CquEkIuGMVbFXQxC+BswS75GBNlG62kux
lIJfxHWl2mJm+9gVY0yVnaUDBrCimwU+DkoXmJCapvRVkwiz11DpmuyUTiZK
c0bdIL+oBAA/Q34jhNYNkXpFCZP8Xh2Qg6kZsssHV6Im8vQMR2eEkhQABXlO
jPkHQnJN0RR0wf5z4bdXi2Clijb0prXU71n/qUO1MgDVHFrlz0nqqfIVkvv4
cmtsuTtGVJge1g6/+qwVeg1MlJObGC9E6VsoqTZMwsrCDrVTsszBk/ZB0vYI
uV1yIXPIK7QHlEQLaEpZvNZ4TIEWMZn97Audjx8PpunjnpiSfDQCEm9nVG4x
eBzTyFt6MudUZmyyjY3h5+rQeN7XaCGJdbHqAvjHzaqaHqG0G/Cn0IYMGZRQ
Cmqm3SHQ+IYBoubp9b45gHjcSdw+F4tcWL4pcolKTXhBtTnI9L/l/FMuPRPl
2ysr6uoeEb1+lMV8s8hTTMVhvAWW+M+5qBLzPW1IV62m1EpJ/HfCwdbz+Yex
QqXkOmQw7h+G6WwrZ8//ZNVA1ECb6D0WQz0mizdXuG0QfSqvFqfRWdyMVJmE
cgAZxZRWJpqZq2KdRMX11b18zLtL+Rawjrq6pv8crw68v3uMLVu7qddpKUFc
HN3jLsj/l6KO66GojVo3s+1t35HFNBojVa9b7RVwj184tK3FcOMe1PGxTR7/
UJFVdPsUPJuKGE559bE19IcNSecBqU+vGCqEAdQhx9Oj3gZE+jQP0O4HJFKz
anDpnrktC6ZSnke8M8XQ1KVwPTrj5nfkeKe2Au9bVD0SjRRJ0LN413tohfld
FJUuDsmzszmpDcOqvZTij0xp98AUiRI1heoSMQIu8VoD5dahp2R5ab57jADx
9KaZwCZJDcYaGWFYOuJUTaH0duEviD+4J9gZVLXTnpzc28bw2wZQvu+t/Cie
UCuqmsuKNBNLIXerALFiVqaY9rAuwz8MXdKYIPf492ulumj38RuJFxk2vXpg
9pxBsJxqVPgaWeAiCrFM3SA5xuxxGuJtJCXabG+TbnATTwokX2fQpxRyCeqU
05Htb8iOSKaw1jSIWPunIxEA6tkMVm1n3NT9v4CHFzb1ElOogXZrWOLEH5ZT
8nqTuhBIxwqDToMJ2uxSOvpV4AD4RcJDnO2G8VPD24g5uVuaSQ2mFkNWV73K
eOEotaEgjmJacw+RJoajozBt82f4A0WUTWfEe/11Qu6q0pqZA52uJTCeKy/5
VEG/G2WAe8aO5/A4JvvM5vYGMOJe60WIMPmSSy68VglLcU4Fw6lbek85SiDV
Nl/FLrEMu9eQn7YB3ZHrRO/oPdEHCDy/JfT7gwS55qqUDdtKiRf+0IUFBvao
ElK2GgBFdOX9wlZM+sFfi0hsY7AJv/EClXDTKBjHx4p2ehMegxokRYGYfgW/
8jTLnLAOEuZnWeGp4JxxG24XW1AqpnhOmxRgxqcvijBH654b1uKRkhafV3A5
tw2I15aYUktiLMweVtBZCedMi0Ja/25C7W+dvdmhEFp+VXVy990/LZ5hJWKE
d60P/444tJC15Wq7FJReIqUi0Lbo+TSab2nTjSCgyR39m4rDjIYHRe4omuGf
TckmwhmXZq8/0F3v/FhUI2UgTME/EiNITkF/pC8KpyjWzV5WevaIhNzWBxpv
2D3KDANDtdV+sW7D/QtENjrmI8ncAhk8fhZGFPmIVl4FhZppjSncIdroCkzb
pXwEfPtF4oCId7YaybE/D4VDOGsNToTBE9QDWk8khd1B0MA2RaQ4OnNFZyVN
jiV8cwDPiVP2QCuXv2PFjOsd7CRbxrYSLdbKt86xQYjQNX3uwvC7Yz/M4Uyh
I7e4kIT37p0vBtAPKCzcnwXuEMDb+1LT02eZYQoj07CjCj47Fd+G1FZ4arah
/rCj5nucOKlE0pTIiDKMPP53acaukpsbWQv0HRX21RVK3R1wMgTzVgagkRxh
fFjOo/E80yCc50tENSz2GP4FSyzyCSR0oiVclGyvFnLDkIsvYgIr60eN1kz+
Rrz+/gQj2LkN5yosSbfUOO3KGv24XyMJGkiHOXblNSByr9H6OML1fqOHNp8A
/HWSnaxH4ro1w1vB/mPCkAwwBa66nMom8qEhm8RasZlwp2o35hEOolxXOnbR
k25sTi7/K6WqOeCwP+RVMMeGyPb5k97zztuF+9hJAaPOTTBsvNUPMLOk2jF8
pcWkVlfFKFWGKhkBeSsmGFKcaR2dgyaEUulmdd6PeSWscWRskRVzJ66lXyMT
ulhGSzBreNaX61hknizWi85X7b4tbNYoFHAazJbg+0Ok3r11nYeE8X4EVTWO
2TJp+zydUpU0sY/kapGvbwnFMvcqq9D5BN5bY4vUoSqzdTy2zFdjNUlfq438
URM0dZHSS6b0WgpaF6vARQHGoTyO7W8po6xgbmSN7CLD5h0xvaQ2eFtZAfV0
FPQ8liuxBaQtzDV0HtaqOZHm81MH8B3kHoGg5KYNpUlXQDJi6l1E6vz5QJUq
vY8wrre1+dcp83fZSx1vf7G9Om3ch1ad/DOdsbu9pm9SXsD0i0sMQZgloTYP
l7pQXoB9v22SRiKGiTtocJKiO2C/LK+55X5OSewswdbrUrBqz+az8Q5B+glf
/BfE9uhzLx9bN34ZcQ0cQvD9E6lW036Ob5SrH4a2ThmPhBmBzQAz04CzQsle
FifTPWe7fG4lx4twtH1bQPZitSJoJlRYMCz2pWedngRDQqAUJbzlG6kdpkyW
fVbRWjECGv9xrROkh/Pc+0CZ4bmPglCsXUqotD9VKncUgL8hM7hA8xGmZqut
D9/RHckYl458Y84A2FWR6FQeaw2rQgb7+jZ0eMFKJxMokh/+AuvfQ1fuUt3S
KhKTjnCxH7zo/9HdKnD1gNHGVZs1ukIrp1jYBEPMMyeJEOJIpgTHvaF5j39A
XBzAZnhgAA7+mgI3IDUrGegLM7HSv+Q6wa/GjB9EppRosYdtOC3ciMjQelsQ
Nc9+T7T5xLeROYUPDxcw0lzFZXdNtz66tIivxHxtEhd0oIY4+nurGo81y4pl
cfyOtFo+qidmXwxgIKHUBY+l5mM9ZAsMXGcQA1mkBE8DczuHZDxSPByo7ltg
0YS+kXStSJEvj6ye+XZIYElJP+P7W/JVw5NqQjeyiCuFFgfvOnUHeNy2KbAq
jwyB+4gqGW+Dy+yfpxhTDmU8Ol1GmyeJFyifs6PFgFz3nnBlAvm41zl88NVZ
kZqqRaEDW2VTBzZGbs3pij5r0w1TVlc3MfHeofjY1cBQTOHciM8jyuSxUHVZ
SZA95VBg2HTmApU47hojJQ4cJbt1G/vQ2f9fCQcsIDEpeC0vgiwtlyvFedji
4hy0QW2G81zDPl2xuwiXh5TUFJ7+d1/rl6+FeKtI/+pnKrj0nIoWxdRsxMN6
pwPpzIjZu4NzFyD1/wT51NtHhP3avK9oy6pC6p/kJ/00LriGDhw6zpaOy4Mr
j5318So7iknrVJDs8dIt614jsh2gJUwpB+g9BR8TBWDE/cvew3XTHiBPodlb
cyq2QZ1UT7RxtRvU+isI1SmpvUmpDTU4UoMEYTzoVp9yVjDzNu28qi3Vxorb
xwPXmh28LN4Dc3QRQYANzeRQ0FLCU1dEE+G+FKw8Zxz8+qXJ15PQ4udg4Qaq
hViJDzUIjElr75c4wGDKUZgkCmsMEcJOOcOIRLHUJ3xRC9K1FTJl61ypqmLT
T23cV3FHmD+86ZgMQbrAVdMZfZVXFNDooRaoSeAlqg1FSqT2iEWt5CBel9PE
nEYAfGpSOxiHGtZLECzfKvvaxP9sV5Ac6f2EwhVaQFr73BGEBrLYE3Lv2NUk
fuZVyMaOaJyzzdHfpR3UKUWwfe7K+lkOTyCkTSCkR49YupBPJ5PRbfM1zqcZ
GbJtxgJRhiV0Cp/dXkaxcvB2fu5tk1kfYtAYcrB5BwL2Bo7tJLUep2K+QIrK
tpJljnD0csboi+M+ToB6kHvDF2wmBfpEJfrT1R49jrxGtAK0gFbLABAdVUs/
f+BkwdpQd83cdwlBuQFo+pYtY/qX9I92KNaRfPkS19PDwZdZJnlpkj9eEu9e
G3JYwKbSxt4CRtNTOnZgeCeG0F9jFiVecsxV03RcdSnEUzTDeNgrtFQbIU7r
N0eqexnRsV3ZfMR0/QESLksT+4duveTjV7fQL9lvSykyPY5mzSGbwE6SybMe
p8VebLxKCEDVTYakv++6DGMwl29PU3nhA7Ax1La+K3JoBl4eIKYnZNiGHHSk
WaDdD6d0m9167T0XwDtm/qSBshWBQlZouw7fdEo/sJHM72dXNReKCXtEYm73
o1nTDxKBXrk875Gge7gndWqgiEO8+wPlSHo5zAHX6ycCMzGGw3SGqkMR36k5
p6rQyRwOFyCywEvIEpdsyzkUk1JS/rtDiUgVHmCyYTknXJI58RVghRCnT0Mz
QvUjtp6Ggd84djrSVLYElEnmVIkRtn1hRK0iAJwlUzu2N0UG5W0KQY+10NZf
EXM+tQugbS4G1TEBbEtKYHacEzAn4znLIyji/MLLgU0tLHdwwUgrw9aRzBDv
Ffl5vT3d30U1kz+0PzF3O6BEvGWMKzlVBoybeYSKFjlbW31YR4BDOUbvnYLj
4H6OdUXwZgBqVsXQ0jutG5R81lqeIV/QHls+gM+rS35P5aDgaoSRA1gI2vcq
6XL8E8MWvwjzoDIoVa9VAu9P4AS6cF1hZp2KlFxZuN7xQOYd12k7HCHdJgs/
gtaf6NYuGlsYsa5MK/HLxY9LYMqKIdZrdQW3eS0cZ7DpnD14LUIxSqGeN3qc
7jpLxD59iCDCb7WFO9wx4Otx8PM6qcqZ9zAN1bdAP30cX7O8+nabbIIsSPpT
1MRANSBXT1jbJF+N9BNB9etS1++ql/r5HAbvojpZ7eNyia0JJp/QbJ0QerCt
t3EFDZBsPFhMgolB794ssmVpMPXASOrMubvvo/MY4ptRtFPqiO59jgYHVA2z
a7U4zPoxTnF1Yoe+IAmcF40OoSVRcA5/vQP0SYKsGi4+ycXj3pSHIEciz4G4
5oJ0vbLqBWz1Ms2eeOtVhyX38xSqj5sx16j18PAeV0zb013PJowCmxVIwmne
QcFe0lAkqra7x7Lug92ltQRwzKvIwe6E8dJNQKoAcHdMNtsH3uD4zXksHi1/
CBKncd3HoJ2vmPXGkSomn0PLkCN7PN7EBhoXO+tfcBndA5qdOSOOSPt64SSm
T+z3JWJa97CLo5SmmWNltp03QTUdMQ3NjbaEtqhDIRahiFz6Cy7zeVh18LFD
RLGl4hVlsFHjj/6q0faA/n3D+tQU2HQSm2CQRFVF042cNc70aLZ7gf5Hb0RD
lqQBVtj/Tu2qM4oEZPc24V0yJh7ENsFlzy7NfDWzO5t30Lrndk4HfnsD10rC
xPLTtQ8qGUxYgHmFVirpjCNyZ1etuo+ZTg7nHMCdJKah4XcUBau87+/vfsnV
3Fn0UyRd1FcoN6ZW8hRuTgEYrcHS5ZS4sfGhzZT8wBqhEz6TntOxgfLx5eHQ
gRT7TpQI9xirnmrHZEq8hZup3nL/qhMnR6IuNFOIzhgBZulF3PXKcRQN6tsW
QisrgDsgX0RAo8wrzlYg452dnu0vPZSvuxLSaCg3QdTgsVrx+SOnd79t3oXj
MVt4SI23vHq0wow7yUYOIw9YNfoGtQRKJJJPe27InC6OWViIAjWB6rXNDMti
Z3rwrBLlgvEa2ppq2GKRKJAljCjJVWVdHr8Ey9Pf3pY31QAsjKJBbxX6x/Vb
0dicyXHq9HwQggIqD92l/+QmHNKmJ46yyJT8olEOIs2R0mAPH5JH+xFzn6Qz
uOrtlWb9UpfVu4HVXDkkr/ULm7zVcEe50C7YeOunJ/7Mc+8LdkDiiNNFaZ/W
IBTo0Guv3ehlh3OhbPS9XeE1ETcY5eqfVuqdgyNBaMad2dRV05P7cAYKisrQ
kb4HpYsZPAQ1BEnAqskGDH6tgIInGGmOp7QMSgP1lHzwXILX3VcOUEzOkPv/
CbpPfOQLpq8pjgl2TNcujhMZdwXlKdk1Oszss749wPIX6UV1Z19mmpnR8BVG
XIfYdsxLOOG2ShZZFJAQ5UOpHtgKdmf7lVvgTGGFcn7LqpqRVULSq5I/iHox
l8781acf1s7aDejXe/+SQcShNpXcb33iVSiCT6jIhT/dcWP6pLJQQ6kU38nU
DvcneWVzaU0Oxf151F802Bz+FDGPDt7eCMmFg4LRWxHK8JsuglYQKKJEqsHN
OBRykNd2EB+uwyAu1/ObdG4pN3ihWikgN+74JLuCztY0ZpZ5Qsd/k5lKH64l
4NNLiRXWr2nPxRlSdpHhWJUiemASZ3U5WF7j0KBt538bavavM2uhDdVjpPn+
8e4DkinsWSGoXpEhKBUI4MScsRCsRPVYkUUH4yn79VUNfi9HGKF0v/Vpkal7
g36d0vUV/41FR6nLIE7mNdggYFb2lMdNwNIXL2Ws56neHZqWmrmfVSJAPPVx
Ngw0MNZ3o+Y4m+aIHVzwOlx7YLqpfSXKRpHgJW8bT1R7ghFfN9beOURU7EO7
UdX3bzjMQTyoBr6bQLvkznd0QEZfFhc9HKjsadfK9K73XHZQFVXuy39rwGzs
OrSj2t3bm6PJ1vm1PlnQhSy72inNe+EPJa9CB7SrphROvcTydGIySBID63R7
2kw8iwXUx7cYTXg0ZQOLmJG70hchDGFQk8w3CCUZUrSzBod8A9ji1Kb6JqL5
8/MzMCI/N2PVMtesualbWf2y9iot/1LkadoifEDkgnYtOxOhXo+++BHtIbmG
vE2u11x9GgIzgM1aw4uoAesSZwWAb35DH4NjIqBzLvpvIODhQrGonOA691fN
3q4+B/G08wMa1cuwCc/rLps/YumXn/LH4pWfu+jNal3xTXpG09ysrUTLuT6g
bPyZcw/IKYmNvT+/aefIwIv4uUJ9S65psZxvxypcuxl3vecD6h3OlsVGyXBp
ZwhibyVvM2gb4Gv0OpJtU0e4BwEDiARcY0dONFpiYJeiKJWqS60jIwgiIBpi
mj0eWHk6BH5GdhRYmvr6Dx09eTdGbEF9c9vNnUWh6kqlRREgrvTSPfYTy3Lk
qQRs8TsKca8GwnJEWuBnWPLQHtVaNicEcJo/XqHKpNCd88IObE3PtcdNVC3s
nZsd1BAyMIQggCm7k8UdMqzpq+qiD9T0fwmp03b3bObu5BGAvrTRub7AjdhT
PTZHUHPeg7/meLPzVaVFmx35BcTos6NbjJyS5WqYErI4ZBF+N4Rkl3AyAW20
lorWmfCyL11BIAi9DxHgZUc+hEUS36sCbrY3BSJkHk/7ASfA3H8D+ZFyuqk/
dR1peX3zzxA9N0rw8V+AwRjg/0HOFpmK+ZN6Z4lB7azqDo+Z8qWcuKPcfW4E
zxHs07iZeZNbQoatwe4HmDgmPSqz+IDqywfka0s0jSLARrX7+YXTQSqRC82q
TyapPtEiv3/MIS1exoBNN81imGCcrPk+/80Uf3tf5hgQtECoyk284EhdJMw9
4A+pejlTUdlV9aoVMtek83XfYvI/7n4H28qGC47o0sSMO6J9xak5F7/wEazm
2fxJFGjkQheMca+1k4Qf8VFBE6KzKCjvVDJ4uVoODCbqBGvhJsGGFZeLauVl
J6wjaUnmwPrgIXW8axmrTGCaVdYpJlBX0QVC+iH2yCYH8U9gCtWWzZgtjQ1k
t063a5DPjbgvq7Mbxmpqhd+tlV+318RdF+qxNzQsdF+W2aE8kHYGKjIU/IHg
YnC7l64G8zKR6ueMpxr0YI/nL+gRX/608JGjqpe4N+vvODToXUM8f3YzaNeE
Ozrx8yT/8vUcoYop5u2EWmA/YgudBHrsJmTVWKCs90k/z0a7oy0Wr0AqDQ5U
LPjwANoiyEdoB1vVftKHn2CzCua/H/7NnkpPQY/oVBC7n2v7zZgRRXPwD9Xe
11YLs/aqW6jKxaljBAUscnX1s3TD6Hkuly0vCDXOQJL+k4epcV37C871AWoX
VVWowvd4uhaqEjct75NChVaCuvM6lVGqXvAQwBWdde6xb8bCdfYfXgxR34iJ
QKtKsLl0t1+Ll0wdGHJRW83W328/GiE8Nkjsnf2FYbaQjYTfEkLPwdx+/nTo
m/UWvEwjR/PKD3vCQ2DPNQu+z5o9DRSzKDXqKowOFFs91IAJ5qCVKQDKbGq+
VFd/iqxtZMiYgzactHXBPn/b+unBXlntZBpYFMrPEDGU4n4XF1Ke19ENybdf
rg2vurf/nmgZCwESpVaV1Vvxnda2YOXtEAcqOv8Ge9LT+KtoWV8NJEi1lqKP
PE8danunDmIEzcbLZicZd51kD7OzyDiVlvb2tnbkhOLZcEvu4b/ilAfMwMOW
M4Z9ggLOkWcsmVj/p/aasHhzRkHCc4WqEW3Nsl3J0Xf/XjX8Tx8tQhfp6186
fTIDXRtMasM6jQcEH4rsAh48T7yD8B4NdySRyfUhrn4pwyu7lOp6FAJCyNnl
98MRQOYylMP1wf2wViRj5tIHJ0DKxHVnVPT+RW5qk4gb+hYh2rD3H9hH5CbW
cuqpwuh4kmz32xNJanC87x/zjCseViFKHQdBb86N5FxzuifbWyiIPSuSp8I2
LA2AqjNGti6x8SZIxAysJTG5QqTzGyxmD3537uiiGHalAzcd4SH257DJYHSH
SrGu0d1eB0jCvZOvOn5JmF2+FgDABHwuZfZ9UYK0FImoyc/hsFWd/5nt+9Y1
Bi72Lg02E5qsqGg8cXfncs6B+gsSQJV0a9SGBkUkhubb86v73TWyoZnS3wlJ
1gam7gOC+G9iy3qWzW1EkeXHOMYVXLskECoOSUcmFeOxwChEMRCLWycPbVeu
kRTv+g+9AOMcwXb5pWwPg9aYDp1vdh6cV5360sq4Z4yjvMyGOrsift8D/f5x
WN69vUNthtXzITgJrb8vjJewdg48GKqrNrErae/oBr/C6i+npTqBxx64Ks/Z
TjcjUimnCl3ESoAiYNPVJgYLxXt7888s5HslJBejv78nFxNZE4d64mlle0vP
IvWDQvh0T3q+083AXkBAKUP/7ysph81tFmSAx8tRApZ46Mv3LYqdM5DOx6BK
u+MCeMJf5hXm30f9OgCak2OOPLkCXRN/lY/ZrEjW47whFtuzBktf8pgTLQpV
OLk3RguYMXliI/Uvrg7QYXgvB4wUTFutejUqO05zyu7XNbzBWNhlcBSygOCh
PZt0qxV6tVCswO0cyRy9hf4uDOIJDzINnMZow1oMQZfp8WO8TNbeq4GxK/n+
HzJLZVEmhSdkiTQv6dp5asNfMHEWLLoq/lwivThgIJbsgCmdv1YbVWbwVRFV
Der+XSf577cp3vwBLaIdIu62fGuZPrq3GSfDuREgtYeujhFsRCLbsiuuf2Bq
o797vUFrdgFM+0aK1BhHiLMgRYD3I3ipmDsIUlTO3wGMgkot64VUUYwKrH5O
HrRwERdBQO7zj4L1bFegYizyZwD190weLVecI50BSuRSFrwUIbhO+V6gRzoW
3v8XnvaLVdSse9Yp7J7dtp1pjUMhqMvUC7xpBMKxxggGLMYRYtZwqGHYLs1V
drnPA+ZdttcI2p1HnDGMMQed4IuqTcW+POKTH8xpJ+6TUerKouV+B/Fpw3tI
OlYKXTNtJQDqSkf6yd4g34Ay8U9ynJpMsJDJu/OgDo2pEOMViHN2iNX/bpbc
5KUW7yQQZXyFyPWyjkVqe0B6VSD5HLcZYAIEVj78nxWTp8gcvmDY8Bp9wWt3
tpfnbtskGdLtqqN8eZDgbU0Kw5WRHS1p769rF0gFn+CgVY+il1XvIKvAW3Ua
cd1CdpFgAqWqyBPUX+r3QzN446qJpooGXxKiz23VY0Qwto0JyEX0oiufjBMc
WpxRIWLHNA0mZCTIgW3KuvBm+1OtrBdWrUOwWhA8Ehy/hBDeaVAu9H1yK7rn
UuZJ9Wdgq7GitHEkXS1PQwaMUH547dZdyjIWNnylh9EwhwrKJyOh25KfmN1q
f3C75qNQLx6GMhlTiDENB/lhjTu5VvMqktxTaCZ1bSmi6ULZzY06CClTWgbF
VbyQupmHXSKEg3Yd/YQqYlRjXI5Wgnhhc1/NzG7AkDy9UWpYvDAxBzMLYIa0
uoR1RE5DaaCIN9zI5Gg0lpLUTH1H0rb/6X0l5hyMtNcwt0EUX2AN2raRMyo4
2HThWA8x7Zqta0pAVyU/0y3Q9D1y9LQv+L9bJtJPIPfGOQol9df0tWCL17Ee
QG6GFYpu95EF71SM0VoY/3oUB5geGCxOgW1w6o/DIpcWGvz3pnEVDv4F4Lfi
7iv9LaOOvCApyL/dFpXKQlepZleRtPTx2ZbJmzT9L6s02PI7aTQ8iNySmfl4
JmV5g1t8xj/3yaMJ3sX9X4GI68U28CD6vwwvMeODvIh0DBCYNCfJ+sylbG36
CDFJ8+zmheDfdRxhckNYFJng9UxpTghhUb5V4iepBkXPnHIzHtjqWd7N4WPX
/a4qqMIbNvyc/Ii7uRZlOoaDUIVsc5fv8TTeIBSFf8DASeMB+sJ4NtdfFMss
hDAjXBud5ve33Td6WWUARNynQuL8iHUjCrCsmYu6HZ2LUIVXVPYZ4qYqMKAU
DV2JQsK0sXhBqGLa+kWE1SaJHQUmBevrvfEaYEgJnLepvSU9BofjMf58W//L
/MVujqqL138e9S3AVaK7kHxvtWjmtSLY7TrZtj/vlztY7josNnwqYMglzOn4
O9KsiCC6rj20PNGg8tebQZyVX0PRuEqe5RT0kXRi3SnUCzvz1UQOm25qgSed
SBmh/YSdUEMymoe81S+vzKht0DkqOKL/eebIiU69Ajopn0t7eBDCUEzZ6Epo
nDit3brPBqB6eegEzDmmOMjzOitJilMr4z8fOUVrdrLSydMUOoEF1dZmkXBI
GlODK7hOcCWj4GRbcudn+VPrsN/VWdQuI0mwiQssZH9E3hX7iosdTXQEUssn
qEccUOflG8IRWAgV6zTfYYpJss1RYjIgQ45Ij7mxz06i0ggSOhvgSBtgMtku
yQnmQ9+Ks0vcX0rpYZqTtaj7p0aYsQQIQNrAg+NerNXeE5qV1uOhLmzDGDUF
BMIir4916ARzkMKdOUFz/H75Hhor+d6gZQ9lMfYj0mU9vIw+IF6hEJuMv4af
Uf23Fz74c3fuU6G+EY9G/qEDymq4vp0cVB7T7GC0ak+fkKMzDWdBORRdnxBt
wKsshGogpr2uW3E0GdFFndycYjJiwW3oM2npL7w1j9HCvIWpBZ1FFIfosFR5
rtaFuV7m0r7V1l4wSaQax5alMxBjh8l4CdK1NMkesjdN2nxqReuXPelFH0PE
ehXG4j10t+LTce99xIVrfaVvo7jzzqhRTTWlnx+CRjS+aJtFL13gjiHH0Y87
biAlZ6/vHqVHg35xh5w7B59o+8vrH79k9DL68MwT9b1Jpk1rZG2UaIl1MTYf
2aI6sAEmU7GLP/dPRTqZ7cMRJgQPqtyxAI3O+yatdhI12yFQPOUOm0E0kF4j
phB4ghIauLlaRHlRs63MwJ7j/oINcyYJjKlHEjY3DHAb81HuW024Gqcm89sD
p/n66A2sH6n2BAfd6IuqLoanJjkIJNDty6YNZEFwPcXj1ZjqY+B7xuk4xM0Q
ooe+qGxcXlAxpHCdkxQ6PhwhTYC+tXt9Zo1oXJXmAIj2a4djyxDGWUyjuaOX
wAm9s9I/RU9UN0EeraPskJSqPNJD0bgIlqMNXdy2Yi59qXsvVxUpYq2osLxe
xBwZIuFmQhaIAcGk+uiqqP4nB2BDOqmXocWm3dZ1DLs70QoOX9fazjkB3Mmp
8rTVYp8HIv//0Y8fcKMp1k1AwVZn+5Iss1IeVfOhn7hNg7GHFEOaKC3pZO3c
yYZfP1aMgU3B+rJ7NxeO3cPZC17Hg2SFyLnCeMe2rUWgHaQdhJWbv6+9/Qil
a0Nfqkr91ay68tbQL+OuFyEMaBqp/E2PN8ypzRLQI47HFsu7s6hD4Sr9E2q9
V8kIRnUBGRYXXQhQ+Ah/U56A0NyTCbqMhjDnh3CXtaIgaXXR/nB4LqD1xMtu
UFWnhoyBvmueUsSHAYeslYmOLLnAcDN6wCmh38V4po4mJ8Xb8BFxhH9J7F+k
tUk4O7NcvsK0Ebp//cV+hMpZMBONRjpS8f+cuIr6w/A+yebiN56xSR5+xIul
GXu5cnjMwfDS6wQWZI/H7JmrUIK4zhickqBiayta66m6ettUos0u6oTbrkU0
fz+P7lKVgrel/ccFq5Z5M0bgSPfK1rFRjZRli5bPQYc3gvDyzT2TtukfSguM
41UbcEYGax2kiqGSvD+SZububYQxFjCYGR5nH2hn86lUHZdzFhgzWBo5EZRn
3CNYk1dKbMP6IEHfd1K/opJDP8Kj2aRJ0c0pVmHjmpBqv/Wq/PGWzDxo/5nk
gtyhhkOckqdJJcuEzIc4r9AwRfjRcTKiGgB9rnNNX0ExxzdIG9eDgA+vKvH0
a9MBEFGCkjPIOLBap2iRQHvaJQA2A9hFQNRD2ntRpwOYcthGR03PT+EgJQek
CzzLX5L3PX2viXRakohZt9ehKzQuznkXzFacZYUS17YlHQxk6sVpcFURYNpP
ha7WldmGkwg+ABlCQIDvLVwKhCR58T2BCBOuc+tcV5ZuTUMRucmnxJ3CGnbn
rb8IpKWF34ZHw54W0NqElkzI+erm78O8vaZzThxbxkZTu75qKgS5/WTy5tvA
tsfiM9/UBGEgcHt4ajqThN4Rp+f0pIVowouzPV3Z3PguVJdJsLh8s9D5eHM+
YXtwVTdA0xUZYxuu0fhpieSIshj7oJ/I/gx7V58z+7K9Z3fYtcgW9CUvGmtZ
i0XTLmxuHM/bGBOH73Ov1BPMCQ5FXkX2wAmph9O8M7SD3H4Mmvjx/r3xYmNS
hT6ONjeeVWkcJwyXzSbdLZ1Tqv9MvGNW0Gcmojt6Xy868UWkZhzvIkUkoDby
D0H8SrtRfnZLp1KkFhg9I1wxKER8cwqZ3MIRLXpd9qc8htxAZoJDNXnhLQG6
pn63oPdiun8C172wtYctM9Y6jvTNETr97zzulxw47PTdXqskU91CJLF5CsGC
ngLiFfKVMuHVS44to6V4gMkhpxHWQ6f9hhkGMRApozvkrR/NuainpMJ2+LQL
a+/Y6DQqhHS32lyLMVxFdyVh9IVRXu1+5EUPziOxDSwm4wXeXi3W9QOXTaXj
Doh0IDL+OMvZ3DmouOKm1xT31wadkgu2V87yP9DRIvWzZ/OJTM6wL+iFO+4J
XzABQeshPYWKgBCh4HpT2FCY/lebBjWA8pXEiBq5cxj4A7Ye/E7MTNmvDpFg
4mmFzxDXyi7bUCNgnP4yjKMXDlSdR9ntGzMM+GR4FyPiYQq5w2tr1kngaPV9
S6IJpi4j+udkHEDen5lPHwze2mA4MopjXXIRYNLvvLMsEOT7y+6vxCZ8sjcg
t/HJH4L6N2T2vi01zx0BcIZVz37U4jOglNT4yUwXAR3g63aV5VUSAnJ5kzx2
IzEl+Cx6+OvyH/IuVtx1/LPC1x6oNFn3c9cJyDO8xE6NZkTVZMLNXjXkbK0R
yAsItnNJPLOYvhIdN7gqqnmI+jCFIakA9tJvloJDBkcgBmz282oBM0JvhVg7
CJrMnNsFvOp9sm+KPY20kksKqvObkhcntDNhfu8in9Dn/TYDx63usH2u+6lu
OFZZ9QQBECS6rqWqwvfx0UIepwZ/GL7WYu0szAmal7LLO9kw0Eo5f+7Hu+yG
adjuwaaNH8p1ArWq2ykZpbA1cG7SE107VF+kQH1JbYhk7tORv3fh2NFwmzPf
gk4hMvpYVyxr02bWvkeGl56kcfCZvLWBbFHn7uH8UyGLbT/3VwGk/FyjXCug
dxAGIcBokiMxTIzdQI3OiuZaMh53fu4IsDgX4Njn9GA1Ia47CHYIOUH/l+dn
Sy2cZtuXyPTjD/k8F/7dfmGxDds/P4OzP8mBZzpqXf62wKHWQCxD9qpmsjRd
QG1RyocVWFti5c3o2kDzoZ5l3zF+Oq0xcXyZvJyCcLntzOWk3jydkMXp3Qji
/Jb5rkBnkJs+6icBvI+wX9uDTeHLRBcke52RPNeSlPeBVdrgRBpbXoUlK8FZ
HP3XhIqS9ax2ZbVUmptfTX9GBWkDmZdhta9gClh4T6/jYsPlqg7irz6+k5BK
uD7ZYEvY4FCVSNEF2ftQSyttKSRZWhROIEaLY1M85r+mYRiAqxnuydnYOj9+
W/2F5rdJ9rsWW3uOv8RrdZR/G9xpP0gKStMe2y72S+9NU+l3EPSufUM30Dlb
ciZEjNZ9cSs1KjD0PQ9gw/7HdG1aO7/3ZgvTkurw4qD6CGTtTxP6m7+tgab3
oBHhWnM6nzy9WCagbEvYNuOC1Mvnqe1qaznBVKK6QiLNiad2j67KsZT/2O5H
A6SDIylFK/Cm69Pzw9tCopRsT+0PkIHur6MCTanARY+xtELwkScgrLd7Gv0g
bAbBLS6pfajh02JHUbrK6tNCmUVJ6RDwTZ0ZrUHjefoQP5jJehuvwziN+/mu
RiVMel+QpbX0Du9+sS8sLuDe2cyhTKsT/szOhZSD13CKR0ttA4/M8JXzwpwO
gd1gttnNx2P4Fs2uRIi0LN99XXwbPlTD1SMbr7RFmH2AL6FO9VcrwAzMsHrW
+rwYEeU9S7CmjB9TLfpQkNLfJc18esjvB+KXCGHrdaaynSY6mgc5enXiRwaP
PGoyy1wg2rm6PEdZQrQCfkjw0cbEsiyO1+Dmk10YgHgsOQbwg2R4G2v2TAvr
uQLEk6/mI5QdP2TedN+Khk9fb5kNxEVwOgnVXC1KCa0jJEA0JWmx9vungVnz
As1u10ZMDO3bgOa36B1waWNTaLY//C0sfxY1t0/UCwKzXQtytqPzGkt4Sqxa
EKCmnIDi1LlpgzlsBVELszQd/UE+q4ufdaLtrxuUf51bV4ei8WP1a2IdybbP
yHoWbaOb+oaEqW74JAW/yDdKeYi90k+2gcqmWlxOHRWko2rRQWlKF8AOJSHf
4+hMHyTTGUda6qenLvagOFzutFvVKgJImcTZdMzrJ+sVTuFC360hI8TKUkQz
olm1EQOK8fODhVwPGbIB7Ut4o71mQw6QSl5Plm5j3Tqr66xT2R0oKjF/3Vvj
ttPlTl1VXZFOEP9Ax4gVbqA1FsR5k+2chXz9VUBbzwWx43KW81OUA09xrH3m
+rO5dp4ZZuPo+5lf7QkpopHV5COnwkbHXgQDCuP/uCRmswZxVBTZpnQGSClP
Ol+2rWBbQGSm09LkejLNrlJQfRcEUlXSM1BOog8HgVmDPpZ74wM7jPbSjFAg
rCVoajV6gHLzSEcFflVv6JRIIMyvVHf0tP+jSz7smtmOHU5CGX8+UFxX7Cgz
GBhHzEBKm41+CbrsODe55Hgd7dqiNQNuFDdgJ7/ebkadfJvuOslHU6lkK5JT
N8AZd4lq+9qIvtVS/rQVbF9ppY7dtZDOC8FRfJrCkCEMbzmlfD8n2FfTbFev
QbWWw2zpRDtwr6yOQN5VkjxgH5eruql5mSzuzG7sYaax4IeyUqzOrOjykHMK
hzmF41GONg85z6YhEgEhHlV62CoNrkmwfuMvo47BnxWPBcf4cQePZS8qFDrt
3yVcs+USAZy7tB/HTALrOPJwFM/69lzcivSOZMbnn4zqks09F1RTs8nMHm/5
3LiJg6w2lfEyJYMleib8ioGZDtyjCN3nZfp5pSo4cjrWwUcDtwPL/Xoct3uA
cFUR5bZWz5SyZdXuys5UHjTB9J59E69NdKqBfeqiuDTPvTHi0lZAQLta19k6
u6I0YeQ8g6HaC1r6lnTKIYm5iy6A7E9qkQOZps78KeKRzCGl91CuynZ3OV1p
gBF6BT/QavgNFp6q0RhUB4uyAKZ12UoxjL5DJFVXVJGLdKtLy5xThvBg3xdG
C4o1l/PXV45RFkLQhZl3UKhbIos+9MZokLHTx0LOMEtVyIwlKtuEMAlslbpf
o+ZEHtXpGwVqiHZbkKayhZaPa/362wkSsx/A25kt/hR6QA3vbyJDXpVBgsB0
X0ULFqpHY3/AdiPRdqbc5u1K4rX0E+xwPsD7a5ro0u5ERjAqJLpSTWH7Xsfx
zg7LbAlWNIw7JE+XcYFhISYOMhiMzOhkSxnHAacteUVtEg4V1JG134/f/vMg
v1+Y0Gj0hrqn4zowTWQoyMzl5oTeSiP+jKFb7ARZUhWZA6hZU31nhwc7bWFj
61956fzu7bFp88YQaZlAgS6cOxztf5/zFA0XiN4JdRhLuEyd9p5S0KIpcpZx
O7whR/rY6L4F9l9Sy6JaDYzkwCVdV4WpquiXlL2lyPND3w4fU+rTr5DCimPB
lx4ZWRdAcYNGrdYQL3LjCXcw81dy7dFjnplSbHLOShUiXnVcUt/4zJeybz13
t23Genclra/gowOSlTWbTPzWipd3m0jm9OKvLEPX+Ab8MDaEFVdYsRKxy7Xu
sY9vCLR+A49Adl2hG5wdU7Zen3AXgepNYd5iB3K5jwfMJLeR66MGuWr4qdxK
9oHtKMzLgSK/A9jLflaJVuHqcdY1zIjntqCdDB1Bxz46p8QUdJgfMcobOPTq
BH5PLweato72VvRYk/AY3USXCKc359BvciXpdMTm1e8XVV+IcsFWpHh3DjPp
TXSFKJCVIlmRrTJXqCvwkqkiCuwQa3R9LaaUAto0v6hJNoIJM9VdtXzYWKIA
F95rB0plUtGMo6q1KYOf7wo0Kl1tvc9LbB6qCygiBJFZ3CK/7XVC96K/50Ax
eQeaGkb9qSmpcKpCyk3l8fqSHiUvhNrIPlTT6iTd79+AXr1DaD1/2xPF7SAP
KkToaKzU6U2xqDVCESAahcSHUVW+sKmKvTyHQsR325wVkaBuJAVMZ2ln53o4
E3QHFnHMiRCs/l3yujeuh+QtAAnTQ04c99Z1khYMJ0731ExM1i3cp1jPwFgw
iag6iF825TnI+/EHRonG22VzEKTownHPvxnQkCBphe22wr0hPpjT8zML4CJh
l/7z+tbAGABOuR89i862RFMYYJN8tjOXbQDmiG5HSygOm6z5l25/SgODadlb
alojR9j8rsO2NGKaVa5OY8ZaJ9wMga+Fd3jf5+PoRq9Cqoh/XzXXE/PQbsWy
WehxX9Scyv15VpOidefw4S9alQMO8r6RCnmycuVMYDbeNnAzxi3LSay0xZFZ
EpAjkEd08qo2A8pb3Xi61jsWrmFWlkg71Qwhj/w6U9jHDvbyi7CmIvHP3ctD
T58svo7dILVLfD17YrrDO/PV0X6SucuWT6DJKWcIOCEKs7WMUr4MhBUa2Vv3
QT1+OdIRkpVrupQ8dHj6QPBBoLG9FFfgDMImyeR3J+j7ES8qquHWevLhHqCy
fvRH6mQc1BKpNmxS2P4U2pPq8fjygf9cg+KBix7S407igTYw3FK/bUMP8KB0
vhSs97Mt1KGFyC6UIf0MoUPAf/Yz/ZkbRjZuWHQ7Iast+YVtHl4NkwIZ7Rya
iPsP/OVCuQa6j892Tny3Ff8Z3COGYUgHVlZQrfxj+c564pGcsV53TUGpILTU
OWJPXHdeOk4yryvSx2s1ZmDxeXRDdgvheunlZo7uN0GHqDEUhwvkD9rj68f8
TpAvi4OzMRTaZmd7kwGaR+nauVoQLLE+MOfYKsJe4SUPVugq1swzd/qumR5y
KOievQv36OiBUDR3SMGRk4sVW+SRcFSX+3wi/XTT36E1W2TW8RzbCl0r2LPq
OYB6oOuOi/rGRvP56CTSVVutTKe3QUbKgEdbd9oQZOoJV0K8Ibps2AuiSydh
Jhe7M1wkStV1WS4IE9zZGR2KoCI8NKQmIMoNfBFz2CuvfTI7y3D84WQ7f9Yq
jjD1V1CCAZ7UwgZm4IWoSKSeXbe9KmnqGVu3IaPCc+hcnk1aqtpmMB+DV5zX
PgLrFYTIJ09ZfyOH1vxAqE2jFwswUKoABlDQT8Hk3+BnWpqx/owvrb2M22ur
6uNc+1PJAW9jq5Qx4whr1oP1r9movl4fx5m74JGhOjw6OOmuqpqN3Npsf27G
BCWm+5Z1+R+omHnHatyG+OWP0DiuMxhg1IwQ47sDTpZXphoTAS/IqYZFIavO
CAXh9FOOfBW2bj9guLwj1MWpwBwvoWfOlXHZTVLQEz32LBwnKjd4UL0WOEYB
bYlckXUD3VwoDo92wuYyxOWbMz0tmMs4UZ/jH3YHnSTlD2UQqKlOIPIlxYP1
l01t6+Sv+pGdAH8WaXwmZpcKoGYxr7JMqFVoDUWVzH/yPVf3jXOvOp8cBiQb
HmERpkVXf0QzwcUefLz/bMqNJTLZCJZ2yQKQ0Lgsdy8u3RcIiqnrUQ7sbnCI
ZpU9iLoJ6nYdhNAJ3wjHIsybZDZf9wif1hST5zpD+pKfJ7XHOblkfyIevxS9
y5NGrWg8uhACQ4Z+tJO21J/OqMxZ6v5VpKLfw+s53z+djAHJcP1ccQh5wSFQ
abMvHjMS9wRCLYGvpgcRzXKjW6bzaFosmEI9Nqfe1+h/pnDBuyqMUDB35fLh
QM0bcr7QU4rD4urUWoCIRmyd3GVuz1TQ+3zgS08mDto4UcMLRSJq01tjQTVk
0Wwg0V6iwQvHgu8St148v0V/442PsrHnzXqQS0JcTloZmvTd0tt/mbrS9TGD
jqJJBf1IC7IcFBeiyKpMHWf24MGeBmAwlBuuv5kVYqcOvNUF2iX2OEG9jFOk
namqXPD3dpDEeKXPZ5TbL3q/GFK9rqGG+aJX9I1uDgOw375y7R0IQ6VkgUXQ
ufzlfA6CGP0yVWZY1KK2k73yNLB3hA0yKXoyEH65NjP63M1UiUEh1+tUt15P
EDnLKxx8y2XIjnGFx57e6P0ai8GYMb3xjSY/HyxZdekKdbvDABNRCIdJV1pf
SEqAwjkJ31pKZYQ4HKwruZ+67IYvm+t2CHM42w7gjfR7BCJb2hsL4wkRcXL0
mMwisIVfBHD1PGj5FuzlAOgEfPjCy5xxdxy3BqRVDz99/rCry5UqUVFDtgsx
dp6wERYLft+FoEus6R2Um607dsq+XUsALZgnxJRzr1vqy1ZNY45C4YAW5lLU
i5/LHECK3vYslKrpyAQKB2WQOgrM9hxiMH1vs2nCMTfkQZwaipt/dEO36j9F
/YCk3TuYbzbxHW07KMst+OuV9n3kCw/LPy2aPP3AjK5ZVIjVWh9wZfdpmdQp
JSb0hGxmWd7sRrzDqHuBI5J2FJtH9H+o9HDz0wpQGrJFfW6k02+CD806+7nK
g9W+bqpE3Fy45L8G8yVC/evY1JyDthB9x9yc4ZV7GtZX9sRcs4nsM4bsWnn4
c8ZEBVlOT7t+6jp/fY5HQICH27zBk/lJmJN4ruFiiblW6oVR+Kz9Xkv2DChy
a6xhhbC3mPU15XUFpmDzUoGpEYAcxHfhgxrllyGZFc5RojQQisR1ec5kETKv
dreUUBQ9XHAtti8VVWEVRhCN2uUkXb7Mp9pZrn7mdYSOiFQagvp/sbVx4lO2
G8Rz87/x752wDCcLRi3l083ChFgU6n8lgpQENKykDM1NSizPJLspDf7abX3n
yQroQMabMyXybA8IhalsJskcmzLfZKw1aU173CZb82ZTXowheaDgZKRQz4uO
xwGYeP8RoNf48k5g28c2rBLqbtJTGQJarpHxANAtGaEc72oZG61UkpjrxeEZ
i2Sfz4Nj7DW+vLwPH0p/cFrjGF+1oViVQqIjvlgkIz0N8vSxz8phGUxG8ROe
TytZHxh8WCi/XUx4dBxY3P7mW9JsNUE8PmzlyGbU0XoNrtudFBLrH85FQ+qD
dx7Z4fTEBj7aq3Pff82qZCAVyIk2rsaS5onzfVAWB11cmnX756AO1otniS4G
2A0/WkXPWrwG81COBRbmZ8zYN0QRb8mXxAF7lFKHRQbZ9AwNq9s0f90iV37d
9AhnOt7vttGrQhlwESzMwujZFtHziky7TIugiP6OpdacY5KlynbIPJIjBenE
oExQJdQh0CjhKKuT2i8Bp0m7cFc+uCpEXTJbUANSTFHSP6MrFT0YlBHt7aIS
7o/E3hUt9aQWDvSouDex2YtxPYHTqC80nwDil2QyoErnpo9VIo2RRVvzJ1JV
dEFLCejgnfzOyxDH589/hVnH8KddBnpOYa3DjKAj7rFmRuWbZQr/jo4F0Spn
vLmtCcXad4EzeYn9PfAKGGvE3oyFwyQY4OIKDXYXpYTkRuP2p4LznEXDTByo
xHAEL4Mg5mrMQLmFoRImny4Lup9e6aBCq3EcnFYWufWYWLQPLfaS+YdtrlYh
u4eM52oeB9Yan+AiM679Zvpb+N5LEwGS+ryUFmDgFAP+n2ayk1vxbh0YLMJ6
ULvx6j9YiJj4GNPNSJyZOSqHIjz9nd2nAhu6Dhxn/wRvNx8gXEDsWl2+0x5p
jOkNoWqaeteBZXPl1VN2bew3CsvKxxKfkhC0O6gCdC2h0RZ1yJIzyC8uI5xT
8RolmAxruPmWhwp0otXvONBk0pVd94HiXKZ5jnIU4q22lTbEZeV+6dYEoLb5
zfT0sMbPdT98vLZrcyN/n33fhQh+kXUpSl9jLxGm0yP02a51KPMbsW2MkjhV
gb/AAvCnCmiWUKXMVU/2elcxY4d2SG3uPO96+OiXKy4kJcjeZ6uclRZVgPW7
RqcnTnp+g6447VdUxb8k9Op5PDT/PO0iV943/ErFH0/FOb2Hg8sb4FuEf2aY
wHfATKbH/nexbilg6jNbQtDYNe8cPotiZjUD/pYMnDdtootwZeNOVuLXqB6g
BkcKwEVXrTVVvIYgCN11OkJDsRJZ4CDoYp2dinN4NcxWK8urz+DqH510KYyQ
Tv5fCqbgSry0w9XI77/fji8cTj5D2DpdMzbZEOJccG/pF17W/jKHcQxTjkXW
kFO05fVvqzmiUNYYiSAHZ4YnwOIebvZnoymBymMsa1m1INzv9yDZCY3sq+Y4
ekTGMAeE8RRBISUKNIiWAYegohbIhtRsvWptcLMQuGU74Bi4MFYOXtjMurbu
Gt8rr8XkpiOSoSHbIQMUeAYY8uItbZdCSEFTpiZdAbYpTRt96vPcaHFSBsQh
DsiUirV1I4d07/wZcOBAHrspyp7y68umZ2zT2ODLjsrMvB0KnkYwlgNUQQof
kfo5pWaclf2nELIXkZLp4xNNFGyI2vMYw1Ms8ZMIKccElFWh97trzvL6DRbk
l94G3MxWc7eADl5y8GQwhS7OyRnJiT+qqC0ui0Uzck9KH9k4NDkHd06XZYHC
OtXyAunCxLdgBSSx5Qf++hP0ainOXbuPF036KGPVbDuup1vHFY0o2nGpNSOB
ab1Q64Ozv/FujdINwZU7LAhJuqy6bXjWMHyEKF66EG8GShFi1DHdWM77Ovq0
FK7588NtF8gctcysib9PqEP+7F/02boL59vo0FO+FJpt4WTLilvsLr7P21xh
7rgd2xqp3/t6y3GuSZqTw/fhbO8YzOxVsf0MrYYnoKSRoc3ed52BxX2pVMm6
CPAstbMi0pVkeu4FPIkbhYOpng+JHXikLAtAsGPoQhxp4VDKEwuF7c72j+lS
K5upbKjzHJPTuW7ZznJuQdaN0UE/cDGZd1IRk90/io8KOSHwdCRfDn5rYxvQ
0JZG5csfbVPNrX1eU2y78CCce6X+eBY2z2lJPwb90hOwuqFRe7JyCW9y2umr
7zlp2GJSHQ1wb0Oz+N3H+tRtq33S5HMwVuqWkDapkZL59CenmawlbhPnos4b
3+jrBSYpD62MwRozfgY9vWtG9FYwpqGNAsdhTeis+Su0JfG4WnLySaKmjbiW
2iQmpV8nNmAweXwBLA96Hn3DLkhEDLD44wji2T2d3Dkb4D0qMfhUmTJ7qYAj
D3RmMNuMe/ExwieWW3iSAbsV9djNm4FsjvOSHY1SKy8BDNE9SNASDg1BmP+s
+dOiesbLPjwE/THgAF1g7aMwdzvMf0jCdgMh4DPr7kvoT6y329+ar6l3ugEn
wQarwr3J5ltpcju39YDJFW1WQV9b/ajYUXnUIFV2bKkMYuWdH75n0KDvWUh6
pSJAf12WgBXVegnjaD+0rvhlFSUIFF6Tcqq8DHvcauztkMzJjEdNnbjtGmuD
cVOpluI/jWHoFpnFtD/WFf4z7fxJq7GZR9RlcwcF0w/yDGu1C18d5cXEDoL9
AMZzzFc8i+YtFbn2K2Dh/8aSaDZLnP2GuQ/ISsOX0G2fR1hPsmA4YfU9JBCJ
cLY81CtgixpGXCrV5bou4bvMLHDr00dTvXWXhA+8W8zWq+uI7F3m6KF0IEu+
oHv2OgWjR19Tyb+DSrKT4+xvL20TJ7wfsBInW6SHEmkfCxyaGaoQ1FcOiVzx
KZZGJ1KJOZB3dYVLLvnaNQVYkIOmcPi5o2pIDllni6avRwuggTn8Woq0AmV1
j5KvlpIKSVCl3plNV6RUB0NWbCzycK8ZYclcGe05Jt+V+gM8Ir3Nmgm+/7CN
pNt3f2UqjQOKVaNUQe0bNei2D6V8VfbHQyQfcaFEVC3Y3/AQx73fO4DUMV80
PIHKSe54xVudHDcTVKyqoy3QU9lF8MnWLERfYP44E8uhb04R5cijMESQrZG5
3Z9irWtJDXd4fe8wahnKmVlRN7SO4yqgAnx25+SrujJk+jdrvi1A8e1FBju9
Bvj9HzrMx56poTW3Nsjd969FWHrXGcUDxPBTan9C/2Tu42J4wuHzTWvSFVrY
ZmHYrnMP9vRQNZ27WKcsciTv2GO0jbM5XC9VNRZFAbIrM6hGn4vfrK2sPYbY
+W473lgGaX3+JkU6+XxBHHFAr6y+YWVNyHTYx/KVCkQNRm4MWKuzIwuuJNJX
SwqGM1vbAyeWWF0vmq3jUgXxCpPN6GNWtWHJ/zyfscQxXL/xu2nSxQ7lSMFo
CcBpZQHI01B0DNNVaeLNowHEg1FDA/PDQj7As1vwwOJxyBQM71U+9xIm/05n
VEp+OzWVmMiIJjr019MFrApocxDLXb5keGs68LNjaORVasOnn3rnrRTuCwlk
/OsCABcEIErhcBvRUeEG7QE8KkCOkebWirRvBFHLO/nxpXNyOStSxZtwTZNw
Y7mtlYyRywsxi09sHvLjnkkomz0sqRe207Igr19pcScGTeb0KnR4ezPuK2qv
gnHdsAGp6vYBR6WDCqpSuplEnQae4RZYhE5q8t00BD84uO4J40+7RhetBj9/
zQKJnb8+3H+aYozI0FRMTcPnzNiIclW6XsOlcsoGxJHWKggnnxGA+HGKxVux
tAXpVamEtg/eH1ORC+W04XdZZpxIIvXhfQRNlUz4PtoCSfIOFKPsQZObDxoN
JUtFhD6WiDTxw+qQvSQf/QtcAzu64HeEX7K2QCIzLY94WT2k2dX31b/vVatD
oRG0DYSry136Lb4pzPPrflxDpNJev2XX2piCk+0fmoQ7P9KPP/uOVvFL3LFr
AZIXFPB+oycxK74mZq0rceUK9gZ34GTygXWvqYIyJXCS+afzGVJuuiXuCxYA
ms+p6/iBK6UxJMYkppB3NbqpEhpqZpT2vrZaDMpvWM+gRZ8vHR6YbuWqXeO/
6ZSwrXbAkuYZHCWlSt0h46BTbMZCR+R+dhUyC4SA/2BBmjTo6RAy46O39Q6c
Lh0vyqm5W/rFaKOeFgMuVwq2vC/Dr4dCX6C2uFJeWsElrFNB+pjo1GvlFxBE
QA45LglKgxoBoQPUR9sCpd3ffmNthm8YWdmzPmV+V+xamEwh02FR23te/2CP
JLGLXwYYDIJXCu6FZ/6AUVKMDCtVQDU9R6/6g0d8UJJizXSfeYREbdl8moDF
S3BgSxnHYf8MgpyhGzG8vg7m7iy+nQN4pmKdbUvbNDXKh24ZzvllrHrlVhVs
w9t5Yu7q1Qr9VrgJ68jTPQbbBgeS7pz4SdkIvdK2Ef912ZpAe8x0vHXBbJLH
IQGYC9Ho0hSQjcVXJz4pGujD86hPxEongLmVdc5hgszfomqWg7KlbeCEHsxN
a5JiTLg4jZpfdDAUpdHiyVKoqi9+breC0K2CGWKnHKDO0yc0/OHFBcDKiPx/
G0TaMD3FRTSouLLQfPLLKwU9zZ3erA4G7N3OvwvRTqJook5yVqxKaAUu2ULJ
L/+6dBHq3YnZpqEYwE6g4qCGX//GA+9xMJQ+5ElStGXbXGH06FdtTq6km2jx
/DQUFdsAeOFSqNLQtBDXU4btBPAGfg9Tw602ka1VUVC/nlbRNHmZYyLAPhxJ
Q5i9zuZCS6+IKsBMTGpgpCLdZ9Ecb5BmyxEtpgNrtBj7Az+iQ9PpytL5U45W
xOrR2MVD9InP2oKbLcfXAgyoV1WK9PcN3icAiax47gKPYmxb7RdzFKV2bqi/
nbOelNtPkql9qArxPATX4Wp60odrQF6Y+8/jqJO4tMn0qSnYKH8pWGBCbR2a
aSYqg0H7MDiPrvI5IQpEjY1WH3Ie6isVKous1rofp4Lg8MmxwZEufE4jZaA+
bZ2PAw5B7UawfA22uuuIWL1RE/Vzm5ce2uxwdaPvZAPUG+iCj8Js6V33Z+6e
OiweOpjZC9HPI7CT5S213xXm8VFMaxOQGhIBGwNn+vc6wax1p0hKODP2VK21
dHyk4EeOMCoLf64kKMKhbusUagOvyNCGGEEQSCouVdUu9iubKcX3871Trh1Z
AWrCo59apDLsB/TkkvhmnI7lf8CA35RYJPu9JQvdQcUe8vq3mwhN+59cqXNM
D88jQY3a7qW1eAGYpAFE8V9S+T9em9dFHw2eOSRVb0JaTHKklnipn6Af3z+x
camB8aCs4QuK55KOgjgBvvUgE8KiE6vgSWCpsbrFtYTjQhqwtB/VqJqw4H0M
Q+Px1/szn0Q4J3VPdUYDXY7AtN2uQ3eJIkKLvO0GI0Gt9lsvCJvp0DaDf/E7
WLdN42SZexYKKvlVxScFpkoPP7nG5lfTwyawzT2B1RgQcHi3B3+e1LjryX7B
6czC6hJQBNnRu9XEYFmJ3txLsSI430bwv0Ss6AJzJXzwdRI0Ck1UC23LtPit
/XwlYPC+x68Oxz9zDy1+1bJen2kyFl89btDld8j56pojXDGuN3G5R1oQTmPo
LcuXJtO0920Um43JOyGXiXtTM1yuqyWxeZmaZOdsJ51+NVrHmUyW0f0xF27W
h17Gk5d1dSILlHpSWFT+L01rbvqqYzmbliV1hB1iNuefB619vLiUjOoaXGdH
QAubGexV8EwDoSLH/uAku1EcHnMUnbsCV6/UMMvrdw/yrvcEp1lEL8Q2Ib5O
2HbCvTqi/dmZtQb87qo/vNi/kWNyUPndy1x2ZC+Hi2mT8nV8Zv93C2M0pIhR
5dxE50XWaaKOXqq909moRCeYk8NzjhvtK/0vKLKJgiOPq6oy289SSmfQnd10
FALn571WLTQcrHnDTSTtTXSqNU40ditbJcjDu0mM1SlnDtk6iQv58DbXWd8O
BwVct0lEaFMHrk606emUV478qLmkMKUFPDMg8iHkVarhhQQxDEOmGxvFv5/f
VbF77yKJTd9DeUNNNIGp87HG8E0IOMwn7W+3dAxkwERCIlpRyEJ7uQ4E1g+U
WJHCvHidFVI1bX9grm8MyNKw94JwhEBV31oz6b0E7aJvIgq10hkukDAAGBYu
ngf2aMimOV3kS2+I0OuCNzudqVNvTOLx2+9JVjaCvHF9EsaL3p+0ZGZaqe/4
G0tnDIGgkOlFWfJf6ohxCFnOr9gcedSokM0BveZ0sJZgOPdKt6487T/Q1fcz
luNm/WLZWE30krIxed9kPB3seDYcz0IUduaQ8739JA8/1L49T9sWo6aWFePl
IMvarCEBEwNEvpwanTqAfO0Vp6m0xa/CpGr9Cp537D02aCKnBgufd58DitKr
NO1gAOP8Cnis4+ThgdZFVncvY61mWiHbNIGkbdvuaTZIaLSi13U1S9Ry5/Lb
rWAhkU0wDsyxuPjqKTsJBXWMdUy7UR2iW/ZzFGZX5kha4C+/scTtIbwpslPN
YyVoVPoqi4fkjc8Y3Lk9gt8NVDNO2wEIL5GbKBl5vifeUkq4D0wf3IIt38u6
x6B0noQWPjxN4q1E4cw+bj5poWcrk4KiFC/23acnl5A0nQL1uYZfh37eHbWn
6w3CjJmNH/VA3YIKmtsad9eoJaqRi9u1rx8wudTccLeZGelvp4SMQOZHPniS
Ex/+dLGCQSzyOBP2qfeKFz6Ek28r19Ps/8baNo5hsB9Jxjx+IaDOZZ9lPei8
NaoMnV/Rj5camyHTqu5IMOjnJ+cXyZMOxrrHFym5exj0hTeQVrr8wBHXUr3X
FRYBxX0httqMJFB0kT+kmq7QM+GYYzNDuv6fyFzjGUTxdc8lNFjeh77l2K3x
JWKv6sO/pDFV8/BKdFhxSd6zT2rdtgziKZkXJiB/EfUtReoINZtR9EKFT1Ts
S5bwdvEmqMSKVqO4uX4FhQymKbh9Ac0ake6+Yrgq6iqL6CzSHw6p8mYiUfRo
kv70VzeDaDuP9D2lDnSg7Rb2i0ecFZuYTMf2tAAwpO5oQp5z3WXT73NssZuL
34PX2aBVCJHi/UXgbA4H5Yn0mTHTBzJDT5aT7uFbWZH/kEC0fm56VRp7+EtE
QUUn2OADfjcQkpWcLCJ5R3XEpmZKy6Ki5U8C6FXyG16oc3wnV7rrnmIIBJDl
wHlxUsNYVZD9Bdg4Dm6+GsCpJBh8KyzbxDJyHtCYc14DVJGr30QQDJT+x+OZ
JbmTbckSAerCUyePI3ujSBhzqVaQGJBqC8Thm/TZi2rtzd+4DDibD9xoLERk
DV3FvlEQ5j+HLBcICwfp1/NeXr49xtznMmcCUzn/jTXoSl2NZufnBKcgcqv4
mLoscrgMaVsVnc2lclzcKKRZz3sGtIsLZlsobwNpBpxxVNG77r8HR39k0UyW
SsWb5brIprCBXRpo0eJYQVk+Kz4bqBb7So4swIAaiNle2N8x5B5cZYtvvxXo
psP9PBU/7CXfD2m7aQOfqELHbtPnDmdxECS8tc4AF4keMaRFyK1HeN4Nn5mK
LYRJ8dKMEhSozaRegbwwNtQMVgGcnKZp2+uhF3ZD1v+hxVwb+riHzPKBqXN8
4GEvfl5hbAj5j7FCfow0BIW8c+MjC3gQEZDz1Qwh2jyxM+NPxTKi+KwugaeO
xkzrEZcUMGtYztZrnOD8Rhv07pFieyI4WcgpSJM7BzyHyFYK1yo59BE9fy8G
mN9pIOj+1JtIjj16e7HKj5CVWpFKkEZDJkeNrliG7rweEh+vGNxTKxo7HIS0
9ddri8QBYfKq9pE9GMATeXuvlPTwxwJB+1LIxOwJLUkFmFpI9bgEg55qnpK6
V/++k06IgVo3TTJR19iv9vBUuWjftuxgR7sKRKqyQBahETlgP7S41jdz431s
QsqV5uAsx0Ywj2G+Oyx+Hrg/6kDsdqzai9pEglzjL9cFIjNgjF916jBtQ4+O
qsRk1Q8tNYHOOKmnekDdHcNQa/CdjlkoOQUC3DLWugrPVCUpTO4xW2+TqtRV
8wLbbxpUR+AI77owDiitsyyj+OhYKd7Zq1AAM+qFkqNEjTHOiUweXNEVmhps
TSJtFJMu07E80m3vMFspPCCAcrJL3aL7v3eO7YkC+uj04/MHfgufQkYr5EHA
tJbzwuiJUSfjLXbc0Uc4d9NwwEfA8mEO6TaonImU+0e348JrCrSsfPCKSCfP
+kexZw7p/jE18MTgAPbYmpIhEo+lPxCfKa8RwGBbjFP9DSxjX89+ZnwsBw6I
w0B5cPFWVaH3AHraXbqpTmbu7qCjcmvIc3FotJtKPVzIOm2cxRB2fR8TPm0Z
dtkno80VMKpxCMKCCZ4XTHxCZZQF9k0YD+K1208LX8pmp8XXKFm97+HPB+gR
+QKvQ/mzwXVZKNZznRJjJzrV3PVzwF2IL2AITcSR2y6fL5mcP6Zc7zKyO9Ru
25wCWtCTG5d2D0txYAEkeE12QTWWDYvFNjBJZ48c6L/DszxKW+hymkynZ+pO
4bbuwGsEiys7HdaY9dSNb3/VWOG4Swe56wQxecw4K/BXB0nKECbAY1g+e+8r
rSpItnsiRp1dbxu1JqXsQXsBV/WGlGhJbuWuuuwyqaV5+rOKUti5IoGeSmV1
Q9uW1sdTdII0dtBbv539ervDeFU+NlUY83PDmxQBjYq9kaNYlwqXcn0esmlJ
V6cM/XzzGwZHVRU0hLI25uEW5ttZxJCzZP2N5bBwqcEqc8vUPNJrEOsP6CxJ
GJs2p6XqOQHSaWDB4V4ju+ebGj187Lm5HUSK9Pxtnp/m+46aJTnZ8cmwngaS
buua8hEcVBZdbtHqj6GY9/6HURXNOoz5Eg6bN8GvGBMvx8sIlTpnVn3Nk+0S
3MmP8c7mOzTDQr376iblncCceRzRN7nQMPy1kTYI4Qdx4zrsWcrrJ4oWGzaZ
dUFeKdU9/SOh2/PgbmmqqqpRr7Q1V/tcteor0fTW1sJs0oT4gbh55gk6B/fT
u1wmrwZ9yG/i+Cw62G/dTzMm6GgK0k4AZusnIBvrwWu1oiVvrYruIXC4u5JF
ObdLovWWcZaWKcqedThQBq+V/nSTmT30agBOO79hiGjids8Fikiru3SQRLTN
V7zpT52Geel+gqrHv+fgFl409PWcE5nPNv/fK6KzriCITJwWXVDiiuYvJH/E
POSiGRBcnS/+MRhZXNTeNvpzjhZMRx2QN5S/0bmfosjZM9vFoe+NPPbz5qzI
4ma9uFYfxu/ow04Mb4SSrboqXhRwKGktrUIo5g5fz4ww1HOLxEx7CNfb27Ek
rBfIW/mr/ERXO6+rREI4/uOUMiU0gKhzyy1+7/xUKrpIqnu/4IXvDYsz2e14
eStaq1CJvQVB1k+MhzfsDxvNf6uLZqB46WfXJOoK9+yS956PNHyXDPhBjJV+
ZKjLIhFxPqNd+3lKOB9z9XKXjpuwPUTSSXKe9AxM/TH1nu6/rpNhqPxtB2gR
rO94D2oDufwCXhLPMRIFRCugxet3UnAc0wsLsajkE5VZ/riODzBvBMggK2VB
9iSrIGotKAilh0vZVKz6ebArwujtDWtVeeLwAv+JWhrCRi9UmnSmsu8y+hNS
70jAOP5jAdktXx+g490/83Z5dRrsrLNpjZLqmeUSTXG6ltc3XpBOm2Lu8hdQ
3BvkEnKs0jgKX/WvU2h3ahZ2ofPEcOMFvekThGSpxDI956XUvMln/PDgNR5S
+0FCPZTOfaguhBlLIX6fOFbfPsmX6GckaEkosUDILGp1mBqvfoJsRMTPO5V9
ApDL2QjXNa7wwQzI2GEF97TUi0CqrllWoWIZDNW5JJXBIYtG9BgZN6yefpmF
jQlAtPGCsRUSDbNiouO3YLriH/Bbw57yTEFPwZaRDrESGv2zraAxbmuS04h9
iYekP0g9x2sOmw1h+Qv2eXQ26hAr3H15Xs9rE44x7uVxKzg60kAplYvzmhdS
zyp0OptqZz4c2bhwxUUh9DOzBYhNIV3UUPenuy7hgB4kQDGdAubA0wVxGXkm
sVawZ+FgouO29P/qSjYio1edlCxHihhAkM1v1SR3c/SRyfcBbJZPxuI5BWQl
kR/t77dHbvqXbAbOb/mG7c+ovCDzUKSOrPYIz0lMZZhDezWcs2iq+HWg0NF8
RplLmHndBXTmJpJOrr5fWBIqPZyH3vnyCnE5xdnpXbBQ6txYSfBsrHm4QLXz
E4YEsv/ndnFJYWAYhG/R7cfrwmqqgG6+ps33eNKkpTHJ+SZQVpGfHm8gZalJ
OYFWeOY3aQPBVZe4zTPYMZcOyylv0Tvtc8E8Aw41F+obdATwrkPOBUlvIpZD
kDOiiQYlln/xiSH8+a2ZhH+EdpNe5/ElNtpFK9la1Me9TKySbKpkrWhbSpQl
CtepBQaHPp5CtpghRnkG80IjaB/dLrrdCObz2cRXIyawEkwCS5rFTbregdqT
k67x0mHV86OxUbW2aa+iGOQpz7HoGubwx9c6XRBxYKLGBJOaqKIPjoy7L6Mr
TEAH2yQOacgacmUDZcs71sEFWemax1EuIu7HFV3XnVqiX9a+JduEGGT8Olu8
mgz5RV2s/AJShE97av8WdpSVU9EICxRTBhJ6DXTD3Fiq2XmNDyAU0d9+LDsG
g/UB+r9AEXdAGGjzUP256E1NcN4Wh4Jv0hTK3vNbOQzR86uvuKejIb7Lnf59
ouLQ47x0yUYCfyLm3y+w7ntmFGx0bdQivNs3RBuLmHD97/Zop9PwCY8PTeTG
t7l51Us1lLm/abRzPqfQhT+TTtV6gUdt/SX/PJlP/dUH7tCcrnE0qDkWf2EQ
oW8Ry2ajn8vnB+DFij7aHly4EQoz/owYgpxSh6AzRoKNxxt3QIrWTzHiXuDB
sM+c/AadYp9Gx/P99wNKtAWw4mFIe2ASO06du9yRVO5MLwFDqyhMtrX6uAJD
Q5WRHA6cTTgcmX/9XDckpsqtvWQkR/lH6pbowfL3c9C8OWb2uWEZUcI2Gog6
PW6mhcMBVc+Cm8/B51CpbJzAYlTDdHG8jX8evYLoAZq0YhkoXm4GyJsr1qlM
cMKrYZ/ZIXRZ8jjlQKvoHq59NnVR88OcrO3BoU6s8FOmdZbWDys4OTL3+TfG
RwtdAw6GtwsdB75vpkNN7pWUh4UQ6PQtKsTUkO422qINHFHpIqCU+RemEpxv
4ToPLIryqBTorNOoPqnf+iSDJHzHW8tB/JFGYyivwFOSuNGkfwP2i8/h4bZo
Gg7RaYqKytHzlomSKMXfvu8oRi1fVb4+Tp5E4cvm0C0oCB6As/C90hGGzFus
eNgmYs+Io/q/B6V3qdzluso9wzr50HP35chC4Ph97gq+jYX+N2zV+R/GBFea
tsS8+cRDfLjJUOQtGkBmo/Wkcgz8uOWSG/P4/Z3RjHmSmJu0oHQrSGCX32Y+
qwg828W4OEUI9Peh35G0PN2r8fpsb/UfZCUBcIGa5ITwQr264Kkbvl34wlZI
bbM/Q0YTimjQ4LxfAD1wNCYeqP/vUp1iq4JS4LGEmcPEqbYoY1jHh6sDZktd
Fhc8I8Av18B627zsChLsS5a8z4nFC4L1v0zVfBagWsa6oRf9FJKPNLJWMbpn
kx1UPSM+Op6a+WvjK1mixTGhAcsGSaodN8ygoQFaL82qwOjun0ONGCKiBiYJ
jNPA4q7xY6O+ZFWzilU4yF3A+AYR9rfFQIqiTBa7uuffJZ+xmJv7NIzWuwlg
NbkiEIhbveB3gJwT/lzJ0b347Q1G36TagKqtRDQZYfYChlibJtO/Wvbhn5Yg
4yuwIjKEVJZOXV+xkw8F0ivNQWgj6JKxuQKqIYXHFT8rk9eO8L+rrT/3DGic
WLL2UfGFd1K6IYsl4VdPJHr4zbfHhdAIyhnVcKh9yg2nce3sel9gl46QfDpK
xxjakmq1CdGx9ozXVs/BcFVaVQSLec9vRcC5ygDkMpowk6HG/J7ZBcLwtBc4
xCXMd2g8ZJ3Yagm2drr9xk0H9w7ghAwj2792dkl++FT+yYIRawunCcGsjpax
9crLHxMEm45QGMWW9Iql1AX0/KsD9xsPVZv6wlp4NOKJCKWonPkDr1ABo7id
Sv3K9zKqmhu9PqAjuqqI/lwFJmEsfa/za1qyJmgStpla8zV5IaNVcT4sxeuT
sS+l/oI/7CYgTwJEdvqInSMN+Je3CZJAXAeez3H6IUN0vin5z9DNSFygZVt0
7oGXUMCst2Je487u6TqTHIH5PAQN/8U3RdVHylCScXW9FQZEP/bSppLfZAU+
zdWvL2KzS2rOFrL66JSR6wYU6ry2E87fkLtHGfCK35jOkaFdIDTCd+zxId4y
1MCLxSr/meiv5fVxh669DunlPia34cCLyK6xKxJbrjPKu8qkPA1lir2tSxaj
rF9UnCFQtcqQu5uHZbVkND17dQtu/0wPilYfDznmAfEkdhuve9HwBJjiCEIg
5w2Q+Duw17qw3NtzkciMufR5tXJLwJRrVTUyXWa5PNJMQ0d4dB3w675BDRin
zpNjPmIyM4BDSE0zZ6RamU7t8qPYpMvOqg4BQrPdxgrTaDyN0B00WVr/aJ03
MLbkZ5W1xRYjz767zjLDrVJEmYVyF6J483gfxzfiJ2Gxg/5/Xj0Pwd+T7MWD
X/NwMIrL5tR/PGHpj84WpUE1oTCQvlqWHoaKprxhAWG4i+TpBbk6Jvstza0P
Q7v4GDODhAWbblXzdZbxC1lvWqQQnbDZNgJhHJ5HKrCgzFcNL6Gsw1PYHLpv
IWN/UABY+P58HXLHpzoS79LoCWegCNboDmyGfL24vdBu70gBLtOfWYqxKZpk
CyEhvjzWZt7vxt2jFFDi16a7nWJXQ1AAL+n8OAImn2nAnvHZNzISVJ3Xo0LC
7JFP/eECq0cRw6PG/d9R10lETlRw9yKCw7l9/YZKSrf+2dXwjC5G8aZ0MiVM
b2C60iGj3nJYF8UQpgSrUgeKXV8Z5yVS7mCbkSeFKBQnK0JBgEsxlzdgL3Qn
5pp8Gja7VmfTW1YflSUQjckZ4hqipU+ttwUr0+wTLmRQQnsklO7SZVhpkWig
YmKtUh/PjWAASkTxAcFVRS7x8/bTspv/K6F5JPM3O0ANUy88CZ4opvbTDRwP
wJRn4CVpUPWVuviMIDgatk5LOg7j0razx6cpy0S71VHa90KC1039mrLUcymC
MQ4jLLWefuMhvNAfS2UU9UPHZ406WPhViha1qxqcQNw+u1Voohd2qzZf65P0
9eyZNYg+CpcGSTrkKwn9ucTwDKq8jSCiF4i0LqQIyyfk4apS7hW1YboUek4d
HNos3WSrfSAjljjGqFSNT6CfzTQKklJNXcTboi/S3+sTmRsjXjLbO+6vAyWc
d3DjeCIyZBc9kR65d9EN9WqEjQDYB3ZZza1tHGHJ0IUhUyKt/74/2N0VqaRS
FvfQCVu5SpJiXyHIvMtziPFfWc28Cq9UAoGK2yBfqcODXhCTT5M4O/1MJMf5
p/6KIWbzgkxqmTOTEZwDHsza4AVMZX8DwWVrJrO/QoxKe3kpNisZ9prvm1sT
Zdvfvz+dK1m00oTbuoudWEbNxt/8tyRLdlQw4o8Dq01bsEdyMxHkZomtetCD
eXhj0l3riiRM4Nu+XjTrVuXyFvsWTU+7VEe6ziBwNZBn7dsc2b6dfLYuCH4t
Ve7U4Qz9XohXtB6LK015IQy2UXeOtRjsusbzMtc4Xy2OKgHELFRX0qcgGA6v
pAZUEdRuA6vw+e/tOu/5qua7KndaMmYAPy2ciKerwCfk2zZN9633YBOexISP
2RxxUh4xezooNGkqRzNyfgKXxOPlcYhnQVifXD6BW26ZmcheKuNC4d+9fg51
X+HB26XlkE1Qcy0uD+lMKrsxlQWZLESxhg7nUJZDlqiQFDXO5w0pbtMp0i7+
EwijhdkhuMpfoBP+jMfWEqfOoDSy2PVU/tQzZv/5eOCR27Cx0WqnioGeS4ph
0F+yIiZ6M16Atq+1//Nuf6c/czX7AB/eQXIgfQMPmpdWSJEDFd+QAwt1RuDI
AT2jVav12IDdrnX/gdOzQfQKeVgV9molj7rQILzdpoJJ2FrLEeTSXzUe5Qet
8w7cDmtw+nHcDLu0byrTMJXwJAHWIDTlX+Xx4VLfOOx+wzx2pEhrntAPGegn
armmjHrARetJzTrwa4p4ShT6qhegTtbXrn0/22reUs5PUCnHcyK0b2pjjRa6
A19URDemaZrXkS5/IMzcgQBtIcZfxo0zzat7wb69VOiVQzOOCxTylb/AZgiB
5ydObOjYVN+PmUoHxbvhboudzqGqyttGmvczy4sqkLzd/SmwrRjkX/6jJcb6
uAb2B1Ylu4+en4naP0Eb0R8ljl54Wk3aBizsYXtG1V3sEmjw8H/3ncES4wpV
+KXiplbRR9d//JzrcmexCTGOPjqtJs41F3QwpZQpDlWkHpfq9X9+3FOBRGAL
pTFTTAQOWj3EP/jEU5oFE2fovCsyffxF8/vd4gV5Zk42M89a3GMa6Gkfq5AT
no28oQleOAbPLvuhyM1QTnMuoGhOO9XtVXJpK1pYL3zEVBi6tk0HwFs1PsWB
+fFicp32QHhAi9j3l1AU7wk2W0e0DNkn0/BY8FSj0jA354bYqOXCKafHZknw
npvqh+6GC38d/cGKQYj+RiSqsf//4EQZXk21d+Y/WBmQt+a09OostcDDLNgM
nD9N4y+quRqYFQnTV9ZDqzwTKxUEFQZYqagF35jXU0pRTPLTjsj2XqxrdABc
qm+q/QNL7bYSYiA0pDN7tCyiPGDuUJ7Ur8ratvly0y+AWnR+ez7GpYhbA9Q2
T9JUgdrwaXozQXM1t/4vt/B5sAJTglmY6CAUkEWRqGseE5lRux2BNTcMEit/
8aqanW98VuDV+JyAksZ4XC7rqUdcv1iqpEAmLuHujm3d3S26QJk4Ckjibysj
ZhGC6RR3xEFm+sAeb2bs9kXUIkAJUBnCfPTq6E4WvIWrN3pSLog4Zx1rv37j
BNEMVDN80jv3gKsd8EGZhXotrSk0zD6JgGJ1R+Q33Q7C4D3hVfx+HasToyes
yUl7JUOZc0vmW/ePpZfDRdE81vytcwjHKVlrgxZAQ2vW/yPQFERQEbyrTdk4
uAIIRDC9a4CbEAkNxg6hXMG3J9om9VNFJFLEezkp+/8HootrOVjt3XH1NRoj
ezuvNbEDa3/vGyce+uq9UjNMfKIBY4rjMC4JeDkFlwZmp4hFyogzsEYppt8i
TeJUJOagJY77AovMSr8HWYzNLK0EgZUPaP6+Mztd1MhXBedtE+lMBsLtiGKK
cjylq7b5S2rqbav6kBcQViQjnEDXlpG6CzIWmdAGHIOeu1x+c3f+VvNJoUFE
aNZb2eYniosZwmAxMo9HXUQdvjYp0NPP1SIVHFsAlP1h6bVfi4TP1EupExqd
Z2jM/U9pIqUkwx+7+huf/Axyft1snChQpNJE2Qc6ajFXJTwOHDFC2eMpNicD
KFc8eJUQrKjDt2oQfKweHCTDLp5MmDkODdd0QapKMy28yVEmyBwuyNYyorZD
qF3Kh/pHSrKlG2VaEpSlxydYQfK0plc8UM1OEVQuOt2+UuHYumSunaSSLU4D
7Ac1PB5GhHUEtHM6gWAVFhnSvcXX5tiQD/lkaeAVH7S+XeIfZgfAZ9opU7Fr
WElpv75yXOJgMPHsi4eP5LBpJFsxRYYUCwSnouSnm9pG3aD12OtW7QKo6zuq
VUB200Sayvlepl/8nJq/rjodI6mFXOVaU619brIFojUMedt6OOJtdyQiiwDW
DkJ4XjESM0CO3x4J346CG3jsfeZ2FntPIRDAC3hv7kTHF7Ds/J7bDr/GXPvS
awitdUQ9Yb5T0B9NKq/h3+T2Ov6WPpAdLq5wcm0u1GVnj8QSMs+O6/sriIje
0+PsyWqDK9H57/2Z1t+WYCdKLIpQ6WkrdAHqzkn0WliRV/lMZKXzbw1TCdTx
hG9HqH8aZbDdsv1U6ZiIcBH6Gj2eRXxUAEI60alu5rXCRgX+KvUwx9iDjcVQ
cmBMWE+ZtWU25ACELQItbg/5iuVv6Ziy4sYqYcmYYHpyNLLm/7aVoyqvumR3
9op5AUw6K547lyk+EkE5MlJQPrN0sf3TG67gnqW8zEvfTAcuz3jhN0SfZlh8
ncg0OqaeN2bbfK0oNPetWGJ/DNTZeTl2DWUx8w6TAqZbN2MBFEMI54Mb98SI
m+WeQ7lERnEL1VI8CFQC0Y5dlVILR5blkAMGuueFKtq08605hDgzuWitm8qX
a3b2gRXsT6Ofq2jN+jq/e3SOnHu8EM3ZfQ+hIyl9j/vPCBQMzLCsfJKER0Dg
UhDjJjg07UOCUaPs7Gavsv2geSCJmR3ho75ax+5i0KXTCshnmeR6fSraGrsR
hE06lqHh9ZUzIuYEAM5BgO+IAUR3cig6ey00Xk2PwJXxGZf52f4n977WPUU8
itiQAi85V/HJ4EMK8nLI1jOkwlFbD0R5yDg/0sw/cxf0Y5D68TUQgFDe8u1O
Emu2WqO0AKabUWUHIGyp5TZpV2nCKgRO4HxiTADsrAPPWksTIKdS66IyFeY4
z2IQ5vFxBqgctpeM5EoTql0ba9xVUAC4+dpLdtFZ8WsOhnN93Zt9xzUxy83w
HWk23jgkGaNu+a2Fa3hdBT5/bGvI+rnvv2yECtVeJHEZI86UZOsggXCDIcAc
pcjv2X85V5d/GvXJM5IAhoueYPm669OpusJqDiBhLSDnUzP75vnG5AkqKB8o
pnv7/kXFtpuS7X6GyJ6hDB9OwdMPCVG01cgo6rOqVSsNWCbtBdoXRuj64Vdu
VLaoKmnnhISR+lqdllDFFSUUMjZPhGHXjx41dzdfS4H+jo1D8Oxxa+ugd3Na
q4kKrYa3wlw4iPvDaBP0PQbR6+qqZQyIPJ1dB6/U5XxG7HxR08wGcP0et8ym
DHvOMM5oY+eqIKb/JrcqZOsG2FxjYuXWdJRpUkuLYUyJJqc+B90MX1zUBjNF
WVwD6dqYKnrZEocdrYk84MKy7NF5XtxZYYTvod160P7ozsWHyiOVd7gR+XNr
CkhDnyUu136pwVdk4Fz0jOfpeMYDStifxZrHnJalg7aGsn7aw21MEFERXq51
K2i+Gz0+CBT1vsmW82514fNcFPNMQG22AMST+Y4E/i1ny+06oFP5PhP6DybD
I1uVlFOBM7Zz8DHIZclXekd9A5ZSjU4oTwVT+JNHqw/uZgJALsfNdeWPW/KS
oOvvWusl/P4mkl8TeehR+7P8N+GP/7UTrBHxLz5W8F8lbKsLo4tAPV9eC2Ze
7HpFtsZMZHUOB/No2GiPE85PB0XvNpz1cqDdz08whHdhfFhfAanLFKQAkl5Z
jM10nInyHGzICfG8piWVO7aMPjQxlsgOzMOZ0OPw6VWe657H2C4OWzUoGtIV
7oPjDx/N3wDi21+/cY+NHSC7RnYFUUScA4VgNs3qp26oqvaC23fwMz319bm6
Dc32yJatLIlrn/QZaLTwEQwjPYBZRbXt071rh4F/BGGUm3cBFz2TySdclReU
AtZ3jC8Q9I74AJe8ADvZwbIgFDSFCvHfr24zueRMWsvbEyyVqrXtrwwF4Uhi
iSt0z9XwAs4Vw6n4W1aAEQvDRGziFXyOMzv3PrPxxEnxx/BwW9avhX+xBi0P
hSZkrT2AOeUzUBU5af0jowRFw3qobYS4bZYMOo5/qZ8RiUQurFOAybGQgbqt
GCfCNuvk7zI58e+szii9P3X0an06UfHjCgOWOJpGEqaZsp2I5dOaR6SKtAYu
rBop1WtG+9tdoCjMRkBL7dPYk+fmTsSxoiYM05t7oNVGJF7u6dKuYHKJ/J7/
lGkbIDa4G40wO0ArM4ytFqSCrIhssF86nvmXwdXa2ByoJkEYAmBPO+O/TZFB
N+rEY6oSxnIM23Dqxpz5P4c0g3FMEEHab1J+5wyA/8qbwtsuWOJUkXEAOKEe
n8r7dlXeGlsHYS0FDBdip89c+TngHZ05pqwHKlflopyMeZ7OBICIqvi/5DVl
s9HdA9O/ttR8ql90qpVMDB9BFm805CywL1YDxE4i0XugxO++JY0t/NLjTXBs
5d9Kd3dCyT9sLbI+Vb5B1pGWisziQkE8xFQUEupBeqHIOjT3asiSS5XLoZCX
LoQq4BGuXKY5W7Qp/EvIIR+XhUFU/WWcKznfHcNfXKsxvf+h/UpXwCM7/vzA
kSuGvQvL0WvEC7fxbICoMRHmbxackykAXXmAhTJjjDPwyrTeefxjirmS35g5
8VQ/wSSDPmp5dT1keub2ctYrb26SSaT37RrYbKL/t06jTibj2F3lRX2Oz5/S
pLR7an54bcCALKTYmrtFctS5ocnqqhL2XdQZE1OE1kcvl7nb6JGKfQr+bIwc
7thfZTw7NKBqBRM4qZK82FLf5NqQXwPd6XndP5EZtDBju0M0uv9sKAsAHFJg
2XEP/IlPmulPUIMWBULGlh5I7L0hhcnj5n6GAxneuShD9+k15JmOyu5G914s
1d6M1rRwkuONJDfbWg3WwdlxsiDNN7IqDHGqPEMAvp0x7UjBvfsRfYRCacVZ
PqrdWfo8CP8rpWtmRjHICfWTISd0b04CJlq7UErxydRDp9rk5/g+JVnI4hji
EQc4njwQMQuNE/m8BKviVLMG5odknP8ro6G7uNyKWxJ44tum6Hia3n4tPfKW
bFh81/0NhItAwOdBj9fDFhfWR6qiVWAnFf+rxGcieuKfer6z65Rtn1/bkPuA
blIoHwvcIMzQhQ3lmD6mGPSf6HdVfwimuVdnuqJB/UYz/RZK9vYaAw69FDPk
IcTxm11z3jGaFpO7mpYTWO333tqV6OTNx6ovh4/LWAWdQkwZyoGIt/qqeYP1
RzY0MiTeOYhktkkF39tXLFoaOn2B7WKkq8mmRg4OpZe2J8kg0pBLI1luZivA
xJ8hgga+jdQpQZPTGoKXrCuntNqt42pghZrQHqcbcUKzXG93VSayAVIqSolU
WZJjIhdYTocGVM8gvO+Iwvggj6joewbmDhM4pjibViirLepI0XmOo8QwxLJ3
zVg61AYn1ugqwqhGcD9TNn6ll//v5LeNvnKgAw/f/XL5mOeg+nZS2NonoalX
kqWidi6++A3G9HzIsvuoCxPSuxW19TXY8eUlqJFxIDJiqmyj9JO0QT0mqgep
9tKM089JfBF79ciCGF1evduNDRiZOpqlpPi3DwefaKCzHzNyArf+wRLvbB3a
85QfsHDKeL6F/cxz60FGhbHMoilDvTuAFSET9CV3o4u3JYlzhJj5uKCjiB7z
/qTvhR8MFMJyuw4puD3Rw6z53IHZPo1XaEUSjOlGFZO+3OM0bRqvRMpi/U4n
q3UEMSqnFp9XMKXnCW+O3/KHzAGVKobKKdMOAtr7zGuMyzMeWt2Ku6j2f5Ml
Qj1VQ/htiGv3ayGHL5FqiDLxpAJPLWSmR+CpA52YOPPF1l7M3cJ/gY8pbyCa
FeByIdy+5GTgROFGM3Sr8pQqR8Owf+2fm9WuhYlCzCh8Gg/uwqJscyqW+1Hj
QKcnXTBUpgTJD1pwMKUUjmc/fokIiPlXOn5Ox/XCHr17+YKCBPK3HVMg1PmL
LJ+qLERFyLS0fxhT75aVuedQdFW8IV7uuLKZThwqcNHStvaX3ggnyO5/m4fa
nfH1++OtJXeQC+lrUBXDyrLdqzyKpm6t55d82rrt/MyJ5ZQTT+TbGMnIbqTA
X6kWOWp3SiY8yGTFR0vbwwdtwirefxMFw6uUjiIyrG6udgq8ZSxXu1o5a+0A
0iOhbLn4OUkocruEwJV5u5keYoldJLYTAfBB8WhGnS18Z0oYIf79zC1gqfU6
thZP6QAleDE9BnLfBbIrTVL39N75EwEOoBlkiwzbQsg40zqsmSlCKGTpNwiL
hhJ8lyWLKVMznNwpIwyWDzN3Hw/oC9aHohN3H7xB05pSc30oXFB3LvvdUKP/
nKgVkKFPKE3TW7A3akQnDhxFiJxgzT+MJrbsppw7J7Y2oDi6albqTmHao+m8
B1liWqIUYH0cJSNJiuJ6vjvYfntVVCT80GB5APK21Cbx8drba4RLxPA88PUv
WB0DJJqiR/ImdogpWHMXQZztns5SOWYkAEAODQea3vPJPqjCd6Uwpu2kD+Cr
KGHYUGgtNeXTIKCtcntgelspnhZFQT/4ASEYZ5nn+O9j7zk2tDP4iNSF6MMb
h+/RLpgMxpvumKUVbLrmdQCxUu3pgB0Kknqxj8YyKeHWnSgWXkH6AbPbGrML
rE9OmhEZLEx17d0d/zzRa8B65tAoA0H8Nm/8A3ViH0D8MoihDt7YnJsbsz3O
Coa+g+ev5Y1zb/B26qhjEOFpPIqw0Rd7wBX/ZpIAQ8iuB+rLkpm6EP2GHl+7
AS5XVJ4Q4KxdyWtEm4MNm78INkj5Cq0K/nOuohk4MYt2Q/1Ax7wVuxkx6lzq
WUdaMqdpyvgJ9WP8hqTXBqA4kaHtWGcak2TBOOW451rdpRiPcLIOQO4ghMEy
fWuzDWtJ4mZhrH8xFedeHbpBU60Bj7apV4vAs+kRUmGJ+5lhVSKSk2kCxap+
d2o/mV7PTouacba1leb05t9z2xIcukZdZ4H3tNr/ixOfEQkh+97zSUF7+P5+
zFjECFd3CZV+cod1ZPzThqxj3qtRzj3FZEb7TtukhAT3WPlRfe37XG7xg3NC
xnYmlNJ6yFI8ndBYAopMCjXeKoiUhW117tN7ucDFnRpQ+g5Ht/cz7r39adOK
UhHB6X3XY0mfIHu6pggN8uIQF9l7tOgyJ7vpjq6kAeOSnvzhgSnRPeaQv8hy
p6IZpdnEFzp9Lh70kWF/u9nt7Mmtng2MnD/27Gce/XhAlGAZeutHdHYk6AnX
PBs8efIx6e/FZ38pd2PNytLHYJ1B1JIQ4UpB89cNn7Oy0gr+kptgCsOylZQQ
SG71j+alhjzgz+V9Vuw40COUNwnTs7FvYyBcpqW/Tb2D2Po0GscUYcFwcFVy
Yw/HtAYvn9DdfRhFGGuuU1qMnE9Y109kee810skjFVjh/nx6VWIx3Hhd2jPZ
L4EN5hwi5N5GGW9RvdJxsECfGMhK1a4EfI2dDu+Ue87D1AK8ZexYLzfSwm5o
2f2LmFMT4Gnua2vSLTAJizTtYDzfk77vtALCEdSWDjO5pdyqDXgGYs4xMmWj
8nxwPb6jRk7Xo8R1ZpAw7kqZ/EzJXfzbMIFSqj7BX6dmmolTsLyDke4rvQ/4
q7vLqNkYU3mbdVijBIykIz7+0hsaIbdFC2hnz5DfrDY1vjtcrd0gTPk+WtZ5
bEX2TN2YDLwQ1rHpm9LcJbLTkWBIT5XABIhpcH5sD6lL84bFcEn49BFBRsnM
k/pGFR3MzsRXrYSm30JwSzLri/U/X5gSyYi3tWp9c04mKJrJ/L6Ty2auqLXN
q8quoLkRUHgik95tOnoKZ10t09Bctgk8Swvn/oUZjz3TQBo1gE+YNSTnahhX
ebqM/Cmumjx5I/WC4osLaWHpiojXYLVCorP0QDeTsJsk2gxx9HFYYIqw2wUl
Hy3chp4A0eevb8yeSs9NM1xIAlurrtygOIEo5RUOoILbxjn2v2DtBL0BpUbv
Bfr4pv2wNING58bQfPYc2ZtVTCoL2vI0zURbpH4POdl98bQabcagmcmNA83i
T8ze39NKWiyjpgt8Re7Ljg7cZlIiURTSFoV7vpGE+Vs9wNCPIdez1yOYGsmO
ur+OATxk5idbNB0LqcB8J+64aDk3eYpLG1WTViSl8Fg4ZRUK5zHu3FlirLYT
AoHwVW8aBE/fQVD8DVxFXlaQXVfFkAF346grtfPs1f27fW+L7DFcVe6O5k0X
4vza3jWKl2jeWcoihRAzWznKqaYF2USgE7DxVHvUcGRT8d0q0diOE15wzRdP
fpUwGuyg8pcEslU2AjCjD/6NV4BIXS9IE6vgZduXKdYuacY7X+8a5quXAtM0
gpe3z2gkFKq4hDq4YidUmLl0xgNhRTeDGhbKIBcYaC6BZlgXwN+u36ECdVMe
9IgEHqVJ6YfpJroJHdoBqCtX5xST4L5uBflKPkWK2oZZRXbkDhIroetH5Q35
G0ABeZ8HJ8jJ2hVNIelZ0BCoCfLijPFzl3yVNu+cEWhm4ePh11E9Tr9GNZod
NEDvOZ+XvZFahAcY865JfzYoJyohQJQrikCrXXv1PvBflkvRzPaYP5HX1/ZH
gOMwaj3kAQqnFEyFkrNA2G942WSQTZ101SOsAIESIEOMp57zhwpzfBtzsV0g
iIu7YY6SO4OuAFuIJNBZgjHzdWflcqwuk4shGIjls3gQL6P7qlXfWmwVTZFY
VX0YMDuNK1Y7faLi2Hw3RgH8EAd4VoH5kKFnsmAU6zNfgV0QsrvZ7dQdiZNx
GDzx6kwSa6yC8QWtNO+LvB78stBI6gNPLwx1FN5KNZvqKJr3veN5lHMPAt7x
GQ8cIEvnrxVgNU668O3IR9MJ/5jnHuV6k6cUVCpYUyH2fKcvX1VNJIe2QKMB
hJvp17/uyWcVk48Ffbji08vs/sZyeVqfndpu1/1ZAALQmnx5rNwpfi6WXsHp
hQJMEuj1DHnGqMMm1Ac+gDwDEW/0nb9yVpoIkbRZTiEhnUY1WbV9AtFe9iXK
gVQFY94wr6Rjabfs1fZJ7i6uhom45x9DQ1TLVZkYV+qtF/xdt8P3XH+nm2T1
kAJwTFu9qJfaluNMnLB07nLncbvyptIdRwsYc+5d+WMXrZJ7XIPnqXR+q+Vr
ZeFhamsn+YaZ4ezmU+3By6jL+4iCfdIj+SxfGiFxuTNkiNXJsfzgSOEyDbcD
nddVZSENZ8R3OZu9CgGGCyp39KahJSv8HHZWcw4JVjwzpJMiUH8cNfRzw/nd
l8otMpiC/BJVJyTatLZGKU8Bz4GH9YLP5s32+anJhvL+oQyyC9/m8OmyEoq+
dCBt3zuigqU4jd26DQ6XW7jlFReKFq4ZDhg72qGxC4URKPl/U4GGmS5D7XwM
FFOlbQImG16ifibrC10qe1Ym22AslhJwBw2F2V4cAaMjZ9ZWr84jDew5AyVi
Rz0Xt6wf0QFft4erRIm+3K3fJXXlvpc7qbRslY/kqN9nyFWjBuS4dI5c+63c
JUQ+MzHnxrlLtaPfAZV0d9DdAF2WVwCE17KicM94pPlgg60ffzXGr8JdS+o4
rU878B1uzglAntUTm2RfK1sVejbxG0QnWtA4U6bw7XHCDyHNwbcA6gVacw4P
AkVA/yCUV4mhs+W2F8DUFswJ8iJuZEc3p+w3x0yF3eGRm4U/xbYps9TrkV9Q
eHMZdzIXD+2/FLDDh6AL3XHLDMqjQvHikM0pa6ehb8BP8BWmbouqjYekIs/0
Y2ltWZfSAMUlUqhzkwoeO5F3OTHBZCc8f3djP7K1kFypPkoDGlyzaR4ixHES
3rPpCJiKx6KB5clI6xNneXd8PnrSvJeuWmslg1uma20oUJEt8WeAHp4ZVtP3
NX1WXwngRqLeounSyyoOK8JUs8BdQoseB7i7R358YgDezCD/Apsz8w4pWe2s
FOyZ1GrMV/uAOrneuWJawHJ+8wAL/oSO/h8zEeF0D85vzqwTJy3vl4iq5Aqk
/KWE56hSJTwdyJrqLqjmX2gT2kcynSkttXnUn0QN9iTsSMgTFeCwfKOZxpUp
bcbgc6bk+LgEe6n38TeldCqxIgJcpV2kda7emdeTIRqBv+Qw8fIUN6EnJ+E5
2wtFEjaicp21w0fyNgLDET4DiBFa9W4OxO4UVCADj2JnsHD26wlZXOqyZ4KG
4zM7x0ELRTPrD82aRCzALN4RfThKWh2jlLfQNOskdym+6Qb3oQkqBLTiI3ez
kwYAlrlSUPsu2S6ryTg4CHwug4RjhUFb8f9gO95VxTL9EvkQFhDn7j4rRWRt
Ctop3pzdj9vXtn+uBlyMczFwOIp8YB3jn2VbAvcO4K2vlTwQqTxYG8nZyvWW
qDk1ESX7T9MfVH+Rk/HhyrdifmKQ8TXsPY3kABnNIBqwihV9BALwy81d9PAN
DIq1qW27UDaIg3iDZzR5QNOu0KNpJpuCwsGrlNmWJkWofD/rRviFFz3PLfWY
e5IAaO9FIOYwuP2qEqEs3AYDj+4GN/Qh9JpCSgz1M8c0F6iTLEBs4aKGjZdV
3vsrdGxWBMAWutMf0eWC9gEpnTyFMF7MyC86h6YvME5R7uZCVFM+wlTfmohh
tHKr1CCo/IWoZdXnIhKehopDIg0pTYLY7qHR+GlY+Y+/e+F9ZDGF6d3xJoYP
O5cNMzscn2H16k0h2ZKcPLp/eLw7Th2f0cJ9dk+KlFhCS6LNbwrcZZBrmTui
SZxXSCOy+J8+QiWYPE+GCKNFZo3+n0647GJ/Ja2QxO/0Dpp7yI7v1T3N5FSq
voIa3UzGOTQn2XmBgrudBTpOAmaNaWoANw0G4V7n78lQiahH0GiEv6MpAwGZ
3gnXgGW9lvZGMOZSIzDF7YkaT5uSck+gfDuUnRb0jAOK0zT5AN4DB4ncTy92
v/OFcW711xfEx7B4k6qt7Lo+V2uErSFveAPAc81pvuMs6jYio7iuO/NHx7sM
B/ZI+yWhIExwWlFUPHekV5+zO73o0jYt5S2ALWBqQL5zWd9xx9mWP6m7jwRb
wNgTERjHzgvBt+8YfyDJCOdO5GpUdKCsN1ICpcuh7cFZzXGaqG31KSL65DpR
qTaxYm8lLphJEifapZ6GP9jc9a/LOy55CpaPNRoPKLg4XYKlTAyGzN7RRn0c
cyek6oNP6+X2qLzVrRUo++rBP98B3kbHuTe+OJBx9xo66+cZdbLjhNZ8b60G
iEqZvpBkyA8zrdHLgbAF6F8QTXfGwByA7vwWdX5Oi37JSTetpt5sHX8UulQE
GCAaDZLNnWTZG88H9QFJZYClfK/ackGB2qXYbrHcolyHJ9cksTb4odqQXIwj
5W6SqQFWN+En+TjNYtQj1Ca0bS951zCJXf6u6k9HMLp6kvTfKHfnWkr43692
j1DfLnU+hGbw9OFZOGo7r7oNavETwgGuiw7/LIdmIN6cP72MkUC9MfR162fr
/Dz8DEZODQBqza7r2R9kjXfViirzrM4vtJ7Gx5Equj+7z9m+hmtgTdkyzj60
55zxIWW+S3l/UUEOleeLK1y0Lly5wtqczNo7zALCkbg9yxpFctyZc/jA4+BX
GEngKa+YDcCqFtB+cutbVUux0MJx2FT1q8ZzKrgd8DWjI0kv95xE2Ls2Vks2
aC16Lpa+XW7r92BroGpPZgqE0OKFPPJ5pe8QjEq1IuUqxJkiVEe/TkDb8+3j
tgTDmPmxVAwcvWuB42wy6JDLW9sz7PG0r1K7UkGsJ9Y1m+tgkPBGm+hbnJiY
NaRjF+ZR38NI0zxmrrWamqGxQD2Yn1z8XQc/DvzybTAA9t/nSg14eKi8r9O7
Zfz8aNC8CNgwna7KdvVP9956s33ydg1tcjj/CXL87V1Mr2xYNMbhz4Cwbu/N
P6v6QEsoBfB0SnKPRFNVyJcCMaBql9THoyqX8488v5C6Zwd7fThXoZy3PmlM
blGSxgBG4qp/oLoUFoGYfBRA2SzzIrh3kJDVrtFlKcwBvyO7t0sIGOO9JBg8
ubVXa16roVoYn0WHT0omymfZ5BUlTj0ob5mF5nLhNhg73Z/XTRWt8MjJPRAA
A/sbRF2BEemTPN4eNC6Q3l65xok3l/CiNbfScrkIbvip4WhWbOlO9Qq/50i+
A6WuroHHBbg/5qXRSN8j1XCEUZLTxBCeB0/c4hcULIGYL1uamEY2RtR6Q63P
wN2S0e71E9F/mN5T8dDha5hMwCix78L1rSGOyLuN1ElCebl2enha4s4t9/5A
WPmGPo8yMXajnXK6N9w0DiYUiaIVSWodAIfhcU6lBjTJ/dR37sZVDPamUGEG
QOab8k41RhhpPWaO5lZuP7rjo4gtY0D6PeCzagEZWlxVkwf60MsWDj0+MhNc
mLEwKBg9fjjTdCWQBrfTYOcTLLKyn0T2tyh3o0Upj3uI7x1FR6DdzJNR00u9
2TYW8ziUOH3LCC+ZZXOUNtLt4seQY3EPOtPHmbBskgu+P8DywI6/nsm29tXY
8LVGPERbKxmxdN3WlPj0qBTGRWFnJB1R+9XlioGa/AAF65pjtytBCO5shk46
vG8v4i8aJjEqGHM5QVlFf3ImShjNrs2hnnQg3GL1tyhCfVcCMg42zIHA63RJ
2Dkaaxz3KDWId5RpR09HkN566DScFkOJ/sdBZU84eWrzkwAjXMnoLhKx7ZOa
8wtQ/VDuos6jlB5uO9a6qzQkw+WB5c3olODdigm4uJQi1+2a+K7FpadTz9J7
ilMmpsJPAEViRdAq2M/d23ThB7duY9bXWVRDzGqLBqfXdz4hRNi+3wIR1e4F
7yB+ZHmWLVgVUdW2VhVXGTjF3bBlH2TdXu3tGzCaBiXxEXeFQSv3uIAFOXxB
dxsWB4/8oiAgHBWaLGRDnyTm9DZJzmzCuZZuatHY/uYKm6Xofk/m5ZLmv2Po
d0CjTLg97ny4eulL0FjPdAT+na5nFzHg/laMPm/hR6c0KFhvWXpZZP1ythDJ
bMr38jezhxHHxAcv5J8FM8g8Nni6/okLf8pXiGKMR+QMACo1D0XTOL4z6kAt
ftzaIlAS+OxD8GO89cd8mekNgiQ46efHsgrq8m0BESo7HkomFoPEzKIN7P/1
fvKsSeaTYu8uWjiR64thDqFt/hwAOuU1zCGPXXI7otM5eovJlP+1VAaULcvj
LV12MScMxYYGCVQZ5H1TfSIQj2TedLqNne6Hw88+RHr4hCW5xzQO+SWSjlDt
Dn80A3euEanxLSK3cSiFuBqNHsnLxqXY84ZdvSbKE4r2id8GvNZAJ3O2bI5m
KyZ0xE28zgOJ8bviHQgBVQ3Z9Ajx1ZmuyP38n/JSop1G5JEMJy13dyDGOOGf
WNvMp46dGKA9/BVWhi7s5YlAwKwS+ySl428VzjSe2CtKI8kPyKeOdsYsNHvg
ki7Xh08m/LF14Sd/aUFCfKxne6aawsYFsiynABTpeasEBTDmfF7H5grQ0qcE
ayuR3q2j62gb/rFnAzHA2PUtj0Q/pTJZKb7Qm1QQI/SEsYwl8ockFqOUx3c8
RAEJg66EkixZbVfpznMwDH3mwaZalMkgeUixmV+VyZ0LoWpI8lu85VuKp5xV
BnXvWZAP4VRCwq7URJoqUZT/zgXB2xAkIJ/D5Njj3z5i1gqi0oPKiMSeKNBb
qXHhU0x7Ny6R6uvvNCmVUHcGmJgVoaiApvg9lXqp641Kg4nJVeADKpcA2xby
lxskR6e5r7uNCMqm4ZL4HKOflKKou1f+Wl7Cy6rNMySlwoC0oALmml0L08Jn
b7yuKz9QF6cjs1MTkGScNmyXnth5Y+Fv1ifPubpocYyIgTs8N3b8SPMMmUv6
WLkYdU8/ugSMScCPn+EVAWWSei9dmWY0cBd7h7l95+xNrMgav8LhcxkG5PQ8
Je6eZPErTr9TETAVPZIJaQFYr3F4UCGdVlH7ba30b9Mq9iO4SzApU/2DpiCT
kMx2CNpAljCvt/EqaxxJJJHhYOhfgxrO1vGj5h25Y1PxU68bRCt4RtiyW2sp
xqLBEUYDvTeoNYovMgYA+AKrQiuoUUGVnRQLdpxvqGnnzJ4vK43ORZrtPTlc
eOedUSCVEkcUganlNDBJA44AQTlHc+aXmDxkVRsnr73CIZXjCvaQOMzzBbSg
LgLY3BJR9PQRoVrZLMXQxRU+RsNMglsCXfd40ZXRBUqc77iee38uDLYXiJK2
KZ31u0HXIff6qbIlKU9U+dZAqXcfIkCmBhG7FSNGCAH+Ie8PoWvYgdX/QEVL
01OmmnVUCORZqhbL9x91OLj7KsrXQh8RWMbGuQGMXLbtS0T5RqEEJnw6C4GC
OiVyO7/TDnfxs9abfDGOJcj2dmx3PXTILZ+ikRcXp6G1I3vJepS4gRHCoCT1
5L93IqEmojDlt6uNwe2prDX/bkK/otq6n1FpYW4h4r9ogUPkl3ohJNAnvtEB
36Dp6NGqrJUbU451nn3b0O/BVut4aSe8TwxZQ87O4dleFTufbsqdrUgZN8b4
K72tDvd53Qbhy19T6Ge0eNqFlcS5t4U/fxW6lznCtqavRNEGVRSVpYZizEAt
+XffykgS01nYN73Vp2bd7MuCk6ffdbH9X1rtBx1lPMaN6UdiYnWMO+TIbsgN
E1poCQj1TsKlRoVqlDTMQkuVRNPa28NhyAZyQp5KkbGy9gR//fC6SjUEKKbo
k3erIKaiyJ1QVxNFHqKLVZzy3pEgeZxjWYjh+ZLErOOgQSYMms/oN2uUt8km
JdRX8rCwMHXL49M1h6lbRO6OPH5rBj/H1JOxTWVg3a3J88UvTYrKrf+T8bah
D+tMjZgoVt7Wa3qz4UjG58anpVwO3Zmq9xX12vygwcmhToprUq65uKn3LlXz
/6D0RUpREgv/BH1zAOzdUagiCOuQ1r+VA0UGeVq5HGzAWdbIgpEThkGDyWgA
ejOsR45pjF3emh/0uHE/eyxEnN/06zPYYqf6nUMLrSJmFCpqupt4hNXXPTU8
vRKxntbOOfZs8N9gTQo+lYEp+whfnSVWyQEt4Dot1WpCSeZTVrmUse+ow6ez
SbN1C20KSes4FfKFKTmPoAA1qTiUU3qfzygzZNMz2UE39puhDBOi6eAGGgEu
NjMHE69HeaW2j2AkwH4Oa8C222Kjk3zrqaXr2174WVvByc4am1+A+GygpAmB
TGVdXAcKIXhjgHz7DrijDLViFxcr5+VFavP15f1Vy/MgJG/3fwst1smcohrG
KP8jdA5t4vLi7/LxLh5UewjebrCstJbKmCErf185VyvM7sNx68R+CbvlRjDA
9V9q

`pragma protect end_protected
