// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sp7cbldmjpuTNWi/7MNPFnCbov7PB6y82S3lCpRYgRdH12c7uKkagkSEvVKt
WMppu7M/MrDg3xWefzMfGpKCFWHjp3G43gU5EMD6cw5p8cseaE2O95tJ5J0W
rfTWJ9p4EhKBOuO9UyIQk9UWPAgzQUZxukewl6+E5y34XGT3BW6UC4wQ1pcP
3LVgQjCWFmm1FcE7iaTneypoF+CI/ua/S1/m6yGoudzA/M5cVnj4y2w0nWPI
+uvb7WSL3N9w7+VyZu/7Wpf6SfqAaCNWdCPnwxvMDVprOTxwpJxrD/AElMsg
6y8ZNx1mpJpv1ZJznBPS+Ov5MDtDaEwkNcyiGJFWXg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H/b70ufYrJ16ifU71L1z+e3DLmhIRDxO4Wim8lymAdvTILzODI66rHuFyypJ
Eg3Tor1yLv43RDzWEX85mmM99NuiIotyLPtQeM9/aOG7aZVbifAf2q/EwRvD
z6jeWVbOT8AcBUtRUhLREGklmsRAwa+E/AbK5ufVW73xEFgo539grkbsPBjS
q0oV2oShZ5NSW7Zinx38swIMMX6I1Uy/nH2m7TxjIoLIj0+aoenOrlxRZBy6
D6AY5uaFHP80aU6WwwsJjQFG4Uo/gurYkaaHSxDoKTILuLCs1CTnwZLTqK0N
am9IuLbLOciDoHWWywbUfvbiAM0a/BuEqonLEq3mRg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RDCtz3vxk+Arabtf5xCX4zVRpIVfjEkxelvzOxLOPwh6lL0mP1mb1hRj4nB9
t6ylwI8pHdTa8M4s75CkBY4LyEq4KVugcDPKB5Ys/VN1i7fWskP/ZIfn/JuJ
KEef46oW4gOD+VHIT7bXtWv9NBrdvdbDicJe7WGqRzbcGhXRW7hK4hfibvBQ
r/qoQ65HM5qwoxXMglv6l3Ej8f6tBeQFH5imARahiJKpf4/NZ1lvKY0rE8nD
FV5NVI+jzEpJKHWcXu4po0qM5rmc+5FT6zBGXIRjQWX1HYVTsOGP1cxB50R4
zIbr5okgwy2E+QW4PxfRF09h+6XXqauKF+DKZ+inzQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W55gL4kRqos0k+BCtE5aAw3npM1pcrTwMMfupsahsUNh5pCDu6BaymXZZM86
3ufwQHnNAsJ1S/ajF9qwOu7Y0CK0FflMcchzpPMzvMAslcz/TemYF8aP6Ane
6PGgeRoHh7oAOEWNOU4RNFSGATRF7q81i8QQ0OxCjHAlZ36PInU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
QAfQ3Up9LWrOzyEf7IsiubLgLAD3xiNo5hp59EWEprSB1+Xg5xahL0Oand+u
cNdYKhJVxbRRkF3hbA5yZBbsUOeBh+WK4JIwmQJgW5mb48pSyZifRfU9YINU
+BwtvX/IRTE0ffdwd27D+jmX6TSttO9A3+LfAUJQdvemFINmE+iLCbwEDY6G
VfhZ6oH8dGx59JDfG51Smy9ouqEBvmgyQINNG53fOOa+OTpB50m5GW56KGcu
k4hAn2Mz1nR6Cb6BFyCjH8hyH1QRKG96yKPsWH5JarsCm+pzN+s9n3e0vlmT
XtIfTgahZ8MxXby4HHLlgDbvvXl3H/+OWXO6KtKAaIqHzOHswcdneSmvK202
wXH6Ff0a73bFPGSBUvA2Mwt7MtQMLj3dyxIdbwbf+mN1f6x2DUMSW20UinRw
IVuTkkXqyih35nFBwMPYz80k289qccWd2xqhN1pzl06TU0OnoZjMqCCbBS/l
SGWudQL8GXrM0XkkKZDtG2BZbUwfa8/c


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
t2p+qLD31Mac+iXySHE8jOYnky/5N0iQxYWvcOvK/PyBtOI7JFF9imj/2/No
B2PX36D8MLK6oxUFFhAPEaFLqzWW6xrz4GwvS8NxV9j2nS5uYBRlfW0NraMK
R46gQ9BynioO1kGDrRoIcLkLXnIrIsonk/YpxQUh1vgdobSUGW4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SEfAs3XIqTAsDRQWGn+6fxQEBF8f+BvDLiF8EgJNwyBdIwhVPEKZ3Xj+AhZn
ojnO8RUdlvNH9Bf7XjSXAErxBFaNgqhMdRxZL/V2WhcpfhmFj5mKiE/lytzO
8mHUL6oOIH/g8PJEkUbFszYxUo40Npw+dzVvo8jJyZDnPBp/kkI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 24112)
`pragma protect data_block
TDzTaccyd0nPDO5gPcUFpJBKRKt5OhA8w3HmdbXrPaFvvMsLOkK2+gJ4m88M
DJB4arZv4BUFC+hUwDk7Aa8axp+H9+J+LuWQ6LoBGEzj5h7uqeVlo9fVYqIY
+CZwbq7sWdyr/7ntt1/XpBbJfBevJJtSb6aWHtF4JmagRjZBoRzxTxRvjl4p
DG21ktXosw7wIoPpMTdCl4RbpZuhcnAOUsQ22qE1hk5uqwG8Q53AvX/WQXcO
JRGtt9gnmbr5oOuAl/HkhAkPyL66QpJYrs0oidmfgKPHvIaRarkt1KWDsnOJ
QVmon4hxM2QoCivH9JWTq8lydUnxR/L6d5xfSbGeADAJVy5obA8jetKZf84Z
wr+5tDSIcDXkl/fcXJSprebXhJb3wmoe1hZz0RoeJ0Ltm7UIiXkLZDbBUb2F
ri8V+Os/FLOtLUZlE2iHtnCF1BCG8N7e8XGZQF88ByEyYOqWAoWyhLYVt2BM
Opa6z7JVg3wKI5VKo3pO+xZ1ZoDjpiIMxTbEk8TxWxKyKKDRbwpyroNe5hcI
RsW+UXiWpm6OrGGYbR0nh+xooLWGAjun+z+RJ2uu89y2FnypkfadbvgX2vv9
j6KmxmEc35VvQGQSx38ndwUcS9B53K6z4E0Q22HnWp/zq+YVYWtv71clO9n5
p9jFTHpFR6XLNbBCyqCpf5dyGlgpMjhQYf/x9qX0XXr6jJ5XgAij9/voCE3j
vUvJ9Wz5TXdBTL3a3Hq0mKmz9/7QuyIPI5MiL4WSW0vdRCTcYhzB9Lgs8pKS
uobVk4zO9tgc5XaJw9cII7iy8tCfW8KAo0OK62BIt6VpfUYoeoB6ptfZrlGa
+aKruDUi0dxXoL3EPGFj3CeF1cfcFVjqx46MK5k7TEv9BnDCup0W51YZn8SG
c5TARO+53FGyvfu235Cl8J+MIwKvlFsG15sEIKxjwO/kD+S4siubCjDG/sJL
PQf4nZeOc4Lu9OUeriJTZjxxHHpq9YqgLYmg2Gdg4D1v2t/yM3mGAJQ9VywS
zDcixpkcQQV+O9gWj7eQX0/3MDEQQt6Y9oPYHp+ioD7Nbsoudh8yhodn2Qli
sJREQaxvOfsI69JQkOdhCSXmUtVpmwLeVP/KnmCX4fVQM0FoyISaNU5rnDA7
+Jn9+lO7jvRsAyhAVbdSM80RbEWhixgdR1oC0HDTq6RBkcVXhLFdUeobDIM0
1ZRiJ6MLqwj14XMY4XdUuoAflJHffXl7X0uX3wm/tNsCwYiUV98fUkAW2d2s
B3cW/6QbW67pAjXdS536Gs81ebrGjS3iHKpr6OFZ2Cf1+RqesVoC0qmn5U2O
0iUNrk5w/98UgPJH675RLdGYf/QkgoRReMA2+Jee2/0HdZare7Z2ieEUMc5j
qHiFZznCraeCzJD0pblSiJsVTW0kKhHUVCINAVOTh09OsJClaC7aakgFfNQi
NIZ0p2hOfexcAXeMZ1eXBnLwYAss5sgpUkfX+NWb5DFZH586RUpVXvlfPwzh
ODJxngurQAosc8yjE5Tkep82uMO7qhvcMkZwAdh/HAW1k5Ky+fEADdRz1QxU
thAeAU+m2TcRZtQgqr4ygDPM+k4H/V+gGm1TuC2fnLtxXt7e7uBfGjOyUQeb
OEv2Df1a69FvutDkP5EVGZkU7hhaHkUoYO18yTJJKnCMqK81zOvJqZDbezfY
2UqLFj1AHNwPmaGKX40nbBniKSDOGmmi19KYZAbX/nW7vIHw3vezNWoII8lU
utouloMLGCE7cKeEGlgKY9noAqMa2dg7YBTAxnSa0OlvpvxhJGQnqPqwtpVt
7ZRcBRVTPVXofAtK3EC7UBoY501Kpb0y+lGj1OFLWBJ1RbULattC2t3VQZF8
95AtCT9RMKbg2KP9cy3n/0GcEKmrxs6ine6N1r2no+n02xxXOlr7kqd1UyYn
S5SfDnaJbiX5bCgSwvA7Dt1R1ccMzFo2fuQiUWoXbT+kE3rIqfvZEW80leh0
Nyuhupx5xAJVxVgiWnq2BQ1beT3RBEgJFGBVUKqkPK+dskmcJD3iSRR30Kyh
UpX1xFNqJOSLYmxaeIptlHIXAR2SCmJdsxy3GFJWsNx72d1fseZbDowvc9il
dagDWVSI5GvPGgu++mPi6d0oQ1ZvOJL/qXPCQ5E76BCDLK7f1Q+tTEPOhcnG
pl+UR2SibmhCJbGJmk5hyCJPUMXE6IpXqAQxlXL9mQcBYcXjkI51Hgu9IWZQ
297KsHBuDDwgNY1BoQWFJLmRlGV57zSnq7mbh1lD+fZgrcJ3RaO3YB9bhJaK
CcQWRAh1rm9whbVOWXILs2FxPCEj13nu2LqUSO9vByJhDYl9f8GzPQ0Z/FH8
jpGYzMO1WGsryPAoMkkY/8jugNp1/nkBHHdV+JyxTc2+Wd4L/3s5yrIMIEyO
FuH5CljOoy8NS+D0F+N9LNT/nc0zmwGK5M0yUL7Pmewz6Q3wwrjxcs+k8cQK
tikLi6g4zqHW04KxXQWKZyuRknFMg7D4YN4hpKTJu21hA/6OPIzfnc+1RkY4
UBLgTlzvzklVpR+0mdXNDcdJygpe/bnKZXwTFEHDmqpzbHEjabUAmpRSdH9U
ZCXFmI2LjHeT3QXA2LqqK5Vrtd6cctazh3w7BUvKwzSg031QrMUhZt5r2LVU
CFtuuiQuuo8vzXKUcqLZI2ZweeGBOzbZxIJfq/Zb+PkR26/ldmWtYXeLh5Fb
tdHa1mQJHgewbplRoaRfDuSdT6QX0ZGNIjcYDesNKi6LXm+xoUlYtW7/UDoy
WI8jDsgpXaB7X2ORz05dPrFCshWS8tD6R9MIXSIOkSqcISH4tD383d+kUStg
Yg7mqTEre5FeD+/c287Ffx1gW5Dr2aYNcMyuqyh6gwSCucA2r20BZd5RDPh1
6Fb4FkESd85Xy22/OCbSM1Thnmfk9GBbhg2bSOanrY9SzLmTLOkmrotiLFgs
kfeXvNdyBinrLeixiFwTdb2tyxXX/N53FoFh2TMTG1MVe5rZ5BsLPLspknLo
oVF9BksvA6rc0LxUTt7POme9/+22/b5kUZ/FJL8R2klCdbSBFtRSqLn616+s
ElOjlmdkCfMKUA9oc+uJ3C+HzlRZ2Z+k9LH5rTPkbTc+rCEOHUp77kBmUSRX
J9bpENZxlvq33rKG7wbFYV+u3iOGGvPJ8cZmvdDzKgLeZTwRZXbaGVW0N/HC
RGmPiLq0K0YEclmJt139qDGUS5Ug+Ic8SptbTu3FTDIL5qjP29O8k0Db/3fk
4w2Ohg8QJ3oqNfGxTjpTUFPmCoQo5FyxhMGdrnDudzhpSxg3zEW7vbS7OzCc
RJTNvzQvNQZFyAAYOC9wSjod/N8GG5euEwAVdk1cwJczQKjiWNs913AxB53w
vcbWaucU1VhRJGtfqpwngtxqaa3uo3zbvndcSMDHXpg0qV96QGQ4Moj4oEym
zjpbLPhsh67OssA11csJES6vojLJbfVJpqx304MCyWHkWCt/wOTTgnRFPPUN
f0M9uqpTvRN4S3TuePkAtSlRu90zkiNZ8IfikoEiOf+hFdcL8mXro7WZUM2b
TAz9jcGTWpqOuzOMhuYlVH2t2vdbTljDbAQ68erETrl5zRXCBx1WvDMEavfm
EXG5IWSU3C68kg87GhSUub+ymx9DjdWuHZ50ei1C7e3DgZAydTft2la2E/Ng
CzvlsK2Jx39VDMaEHWw++lMp0YyoGghqH2BPlMOlaomHU8dWh7OwG3/bu1xH
UnuLRl9mwFsfmd4V5nN97G5isqtN+2lmgiCX5pHjq1LIyP1KvrcHT6o/+K/1
nwxqG5JMt2FwVAoNswQPw2geVzXMJ6nOdBaR6AkGDH5aruVOXpvf3YIBBDI9
eR6c9qzyaxf8YxpFZHRqTBgus6ecW3v5ATKbii5cYiNccDYhAvBcxrX+HgO+
6TslqVEhSZrqz3UPEZoiHwokpIhlU/QdmkCWnsBcwGxvgRTodpbfhFxL6Iae
+2jxzqWKarA2irPr/53VMgo5Hvbsv8t/YmYpM/PDhi1ea2Ewi0yFrXO0RTBO
vGYbdsnACn7QA9yHdrtChBTHc4HNlGaIcs5+LarvLAHf+0RnFv2kH+zKURx7
KvilpIfwqercpbjtYEvq/trI0iwU2qPM9hJO/sNlvXI+JUvfPKTOeOtzaNAf
OTz5terbHQ28nnU1SOzxFduUZHWBHTWXwQ7Eaj1b9tQbLoUZwykAWML1s/wa
L0/Hzr7hIMKSg3jY94an4IjisBF8+6kvZG40pS0oG1jBkztBg40ipF5e7oOK
cQfopNUAmP60iZE58kui7EKLLSWWzxC0BYQOkXAC/KYan2JhmucKSD54NcP2
wCUBHa3HUXgqUJq8aU7FgDxj6Dg0kgJgEwTfdSnBykwtI+WleOXCoKnRC16M
YlIvSsfbF+PeyVOgPDoVzKWGGoVapKCIC6qBb1UdCFoh29TIJdA5gxDEXdFn
+G3ulI3hJlXy5p1z2Rau8t830ZMwoqwHvRAnlcKnmZQhL/e+DFh1rVoL/SMr
C6g2wcWPEqAzTeMEGdRvRdycyn+B0ko54F618iVLGGG7Oof3s19QeHBByKCo
ayM9w1htD6QF1QX9ZzkG6nfiNaQDc5NP7iWHetMNrNxkvZutOfYuvECz0nsL
MfFVYt9wwoh+zxWyiHYqV0/hR6oR4vj7xecz86U8lULU/kw5n0yxwrOiOXvM
ZJgi45uPYJnRFwEUV62n5fMoxiTuESQa/Wefm4VobJ1EFs4kwe72uEEeFQAT
qzn9oxsZ0Xpr6uWIGR4UoBYW8nF/ZRWKOBBAeJNGf9t0jCuPX4crbIrnrPCs
wlFAaTlNHDo7XWc2A8ihqMr4SXUx5KmibPeXxNxbv/EUWCbu0sJSKS0ETrGF
aY6Chldq/jfl29w7kUf2ZUnsB65x/P0c/iS2W5rseRLZanU+SPOTZZnBOzah
qeU8RhmkyslXyoq/fS1T6IHoq5rpKwOnCF3y69+mDoJMiD8K+TkWQOtI/ieJ
Rrk91f+tZ768Kh3gH55+F/0rQ8i4xeHkmP+jiBJ8hpoeMaIBxnhMv+Q8swaS
9STbDnqGAfP+1hvrjg1VTfYWX10M+PTsqsblxAdcpw2OkPyCGnwBlrEHKfPO
j5avUyB73ImFBXp/zlqLTV6PMRHePFq184u/o/oTRG/F1gTRLml+uZa0Tpdd
+/RkVYmZh1CZATce9mR2C7gJmOhPVIw0Ma+1fuRlFi6HVo9TZ9OW05/AGP21
/aeftkuqp1qnacPy0lNj4yTcVPKOTznD14VJ0A7OejGrMk+WPpZG39BjKoUL
tJmIbrLRh64iLcdIYu/bF8aKnNdFyoYUQYaKgoBYkMjMzjW2UNGAfu367htx
aXR9CWbotHUD4btePbTNs9+Kd0N1n7fjB0+U2eNMFQupNPO6ACtYRD1v1rFw
l2Y4U1bcVkteae+5nVikrA+/2b89HKOp57IjCroSgja0r1nQxtTouNwpbF1Y
rCibgbdQ8dUjjsbt3PJc3ZJjKjX0/vIsl/GWmc5PsNs6JlaGWXuDGbrzDyNT
fh3vTGL8hYH/VJWTWFQfHf6OjIlNvY5IhBoWA96Y+phegId4SrGDovMHWBXw
f8PqVRPUNktZUq2S3KZcp+MJezSy3rn/uiclzGh019NcNrIQeR+1tmZM4gfK
mgTdLIPDU/4LgM8ZDuBzknUg87CNPcm1ut70Y00L3AYaDihrMy8bXzWRcKJG
1xmYGdAiLSYygAu8BXzPE1BupsHmEoQh8slKZP19VfEMX7XeMrfukFHvwZF7
Hly7QEeYlWcr6HEb2Zb71Y+rmdAQo3UELpBXvZ+IMZBV3dcN5hcrFM4aQAX+
6N+bC36go2SUe705l8tfgBUP04mGnVQiCXnenz+rkn9v09iBz6ZDceeCgMtH
VZAt9OAGRfp62C9bnr31EvWdGjDAogOBbawbR7wExIspURRUfzkkxreMYDOu
ThGVo5eaQqPJyQuOHmjRfcQHTvsCZ+UyryyUfbovHAS0AfTAaDIYLFJMbedq
nfhDFJWT0De7HMFSq+6yp8Jg9WFtHwFy8jqlzkTBvGeuIFSDe3QLbYrNKYa6
Ke2vqRsJY5GXjZ/8UQkkj6U/xzQbbEwtCgYbHmbhtIt8CjEYAjCCWjqE9wZY
L29HfaSdChBJHZgX+Sr0kxR84J/lt2CWHVHqZ6dUjWdsmWUjioaBM6EJcNLh
ab2Lr/5NaflPuhllZ6y6SHWkRZU8G5051R86fxpBWdD5rNBihYvmRYhLdxOR
Xe5//lH9MfsQ2/sDnnH1kT7zL4FhVAAmBtV3CS2h3u10N7jmJZUu0XSAo92D
KVmn4jSo/EiikwiBIi2j7neT3xtU3ps1/Em5j70cJXvzY4jDDV/uWhNfP+v5
BWzOI7PvUb8YdfGUg8f2vknTuLuU29hY5OvyrYgVIGKR3qChKyCbtNlIwwbo
igs7/MWj/LrqVb2LX0rRtK6T4oXc9B9LTrW09kH4Hm1cTags6AnARjL62B/I
wD43DCe2F+QU7jzVo3GtMyjcAumOQYrd5dejFkS09gbmO5X+AwKZjsuUVCzN
ffao28WmPFNhoO1l6L8el+O7fHhXa/GC9Or8l5ESin1nE24BhXQpfB62O5F8
ueFBcvOBY2OPgMQvCTh2Q/4RXTDYTGqagUfCfwX8dJZ0+Uhnr6inhRfyTmrs
S1USBs++FzYxdyzMWtEu+4qubtDWXLzJzTBXttztSaCBKz8LPRX4cX5hAnnu
f+w2AtpTweZYNyjYIG47xtJurGuHLKkBmKlknJNfupCsskOG7TbllWIZ1+Cz
rkqHgNRRRqbKOztTMo4Qg2+xE8fuhrtu+g+xsFIgMvFK4QPTxwQ5q0yYNHmq
7uIhIifmm6Xtz92DaHMB5ZyFHR5HsOfoK1bEKrKWyXf1XbZup9QeGUL/NOEC
/8BvZlBTzjPtNhzHX60rGDXfoFtc5oHEOElNCo+1JBwYu1Aqnbb25NeDFEck
gxh6onXDk7HnCxA2T7OK4+hVJ/oP2+jafjyNkkO+bDZXCU2Rdw/dD19QIM03
cLnuCq+Kdbwo4pRDquhkn9f0YG1u9UM7tUPWKR4kI2N4D7G7mSxLiSt9XJPo
SSoMAg11s5QPJmiFVH0NQHI6lVa8/j6INf8Wg3EqKFZdyoPLw1muWmq05JYc
NAlky3Hx3T6cTPCdq4XxS2oyXQJqalxi/AJuwc3m3bhXm3I7TdiduYxstx4F
Gp17G7ORLwdG5PFMPrPVdHYoXNGnpal32t+xHed/sSdf+BbosIgl1qQ8Ylt6
K+ztOCsR3UE7WJ7n5hHAmeB+L+E9gSsruYVUFmMeSYv3P20gZS0Sx4MoXrSQ
axuk2bKWxj4k1mjMCULtnZPfY5pzkg5HhK4eOKEeelNybWVEMjwTEsj6NE0e
kNa6Vf9VMasJNVpzoNfs1m1oEDVk9UyNujuXLIefiQwvpRMdOenhB3Fl0XRC
DuZaRizPG4gOXPxCwQvQ3ySh+/oQ9WMXuzozJl7LayT5WK3POIhAMcAIllzS
SGlPbw+1ay+Bftv0B/TJtk5h29XhqUlhpx9+hp9H7Li6deogp0lRSAz7VKU5
3JSJOiwACsbjrUIj6o8a19D+MqICGDzGtDFPo1aG1CpBh1hUxe8losqiOa4y
WzL9Vy3FVsUBSjTPoIBzn1Qvu9H8i7cY7LJGuQtmmXKkPFC0kKznfqHUiAHU
m4mDhGUXd9Ta4BNfXpyGXS6BFWUs3qtUi7ACvqjglxgzyNQ7K5zdYl8atghq
JE9WFBIWNleCtvfvv+MoXzHC1dI97semVTOMOvCbdWvkeyPDl1zxDMwAFxg3
8S6GDWvxRnFg5EGqFfxM69ikaQOTcscZyzLgi/D10G+d1JZrHVo7Zjbz4CyN
h4vEemMk38LI+7b3AVc0FB2ZUcXAl+UWnd4oijNUmzGH6J92t+dsoARMhcQj
QNKyCO2lS8PLuVmRBPNbZbf0XMRqCS4cLLV5yVHuos1EfxfmqXHYrseFbjJJ
jMlV3DWgT4BSiCCODEAMNIohfaidnzOwSCXj4hmwEAy4NYFxvJ8NQyNCrwJc
H6w63A30j802bTAV7COwOAOMsYXP64jLOgDM+OpmEWARdfZf+9HUnWjan4Gq
knLlpOCaN6HF0JUQqtFZ/t/YRp5rhe/jeiDUQ0I1kFvtqgRhfZVdXDYxawm8
ClGNV313dILc5e5DjRoMKA74VDX22/dES6GsS5xMdl59hH4RgMCtq3RkI1lq
NsNFcfEiU6zWe9FoQgm4+TlfRvPGNBYzc+WY2g9UbWGc/lrGKY6xqyqNt7yh
EjKy1qG+jA3EKavghJ3rbAM7496PfCRWgnZuoUHfmVT9qRAU8zV4hBZdtMEW
ZcbUlk2esUI3shgnkz5kdutl3HRa112UMs5m36D1vgDXB4Sx2jEwK3/K78kQ
4lAt8Pvv8ZDmKaf4PbONYOCh4XL5ZfPgyd3k671cY50KZHTyIFG7Raq0B1Ca
2BpQBowzHBoPqg6Y/1vf0vmY41JSkR/1loiuQr/YWSXj1Ay21NcgALKQwoy5
veSfZqrxztXpmTBmOjK51jxne3SLSNz9AWBtv9Uosak720ez+Opod7mRUDK5
9RmKZ0U3iIYt2RjqUtgWnSaESDnXEVaC6eoJFQCphU2qPXssAJihISlE+jcK
faTKbdVt+1tpEhKdJuasGPWnHiRLcssKUtjMpVFbgPcxWAdw3C9fsPlxhcPJ
LRciubWMyalbK7p+TJ+n6ilTu3FyQkFllPT0JhPMG/h5kzSpYvPR/CAQS6iA
JN+S6rDXf807KPEeAYLZ08F7fwsUpHQklbCGBc/mD8nAqcAIaVPkWzk++Ikg
b3CckR5Ett4PU0mnELVCADzTs1XsRtG5s2vU5AiyJ5XpSXorxR6Mc8RAsKcg
sQuh7BIYDHGAdWK355iwY/STmvQxuxZUKrijTRPEmyw2SyYz8F6PhfHVIGyJ
hq5RPOjL3isAXybb/97DXXAJDqH5kA48Bwv2nO5oRJ0AeU8VPM6BRMedmshE
R2Yi/Ro7LMrrn+2ewXShcFDO4gIj8i6Fyg3tGnTb2PdBFYpFc0UhTVSS8wu1
ZJiH7zMPt8P5sJGYE5Ai1wk0EuyTr2oevfsbbz3GpzI/k3B8CBGByEO8tkP9
yQN1hiRaHT11/5mlaC2mqMCTY4iMmTUPja+4h6YnSrAaqYt0RlJArlT0WQCH
FKQZxPdlry5XZfY5Zna4w3IIMXU7yWiPTM7i0eq7TlGZuACfLPhUZA+KNsio
x7V267+5JHuzvbewk1hszY7ZMWJE9j+9z5AeLiLMFQD6Im0MAc9mqw/JqLiB
BmLNLzm4jzON083vkpiNGt6sLr9+Y0Fg+8Xe3nJ4Bwp3wq9HPIRktT+7KlQ0
2zJ7j8/iFJ0f/QhCm1VepxXQh0bqwYuc8U25StZjDC0U2Y0JzD6LpM4HBnCG
oNmccgnaoIQng5DR0etY0SQu1e+p/enxxpFfp1qzj/gVUs1QV1vmHF3hEQMM
bCm7aJI2f8B7Tc46izQToZCljkn7r8ShADJDrhjhy4esSf6ZO0s+B7bmta4a
cKWgoocTLB3mgkzq7u1pJXFJHLRksf097MUpGjxnMxLYz25uKOkYZFFLwjLp
mVDWd8ZVJ4CLUeaVZCJpN+AYkOpQsrWAmOUw8ATsskNhO07HcEUwQLYYNZxw
aLYNinSN9jDPz618yrWKd7wDpVHA/2hWPrnfCo/3khSKASkYQ+2aFLwcAXJL
YfbV/KJ0SSAv265c9yzoSAtHE9ZGrbwfaecaWH86A4hKCB7PiqaTSt+gYN2c
tocCweITO2yKWAMbPUINtHFAQYgfj7pjJWBP2hKZr9rHga/pPHOhrnQ6MiAU
TKkppmoabtWStonxGmdlOahbF9dgYk32CNNpzxqUexwM7FDo4gpOzNENTv+3
TCIYH7ORCDseu1udj6FNocj88y5gqrwfSBqpg4vPYt09vPneaS0rcJ2cU4oh
Se6AKi2kaolGo6dzWtf0R5saTZTpJpKCW1i2oycKmBdimRIjhx5Wk4CNNAtR
PyY/Po6hqhh3kfrnxRQD7wK1GRUZ+dPIKy1kzCD9SU8uj3n21Zqh1evw+WPP
craLiPczEO326EPU38onS7Qkto3uQlYRQPSoSzJXHhKVbueuRt4DEbi2rotm
4XGQ8C09z1qE2gnTfsepmF1wELh3o63qOKdXvh2iFS0BYX+cw10rMhJpTa5k
5uJX5EyU4QB8zNZGB+BXg2DQcQ20B2E+BfMYyc6xcy0qet3JWhP0WcZ5w9Cy
mA6o+ZX+DT7kPTxw7EjX+fJP7zSLeSRs5WEi05uQo/nacf+xUUMRFdlFhQZJ
BYkR7PcWwjSJihMp8yvXYzfEhYSD00RSfNyDBDH3tRly7y21NXEYAqYMp47Y
LhxeV2tWAOooDNjwztVJM3/I95q6yC+c3tDOdpmp7Z9xnHIwZB/C9zWkXqkZ
jAuq3/8c5nCCC7darN0oHSvCvjG/g2Y8oEaP0OGyxTUz7iD2aNcAML3/VoQn
e6CktSA2qg93EYEpyXpgKdNdqxvVHOZONJaeNBuCYJnZFyMGaC9G3FlFeOMM
rSI97hvM1jpWh4tmNNmw5In0GOOZhVBWfJRf/OOz4ca8ES2f23DtRa/ZxcQk
PBORXkqRN/axfzEJAPxoJLm26ur90B5T0tLP4Auyh42HRcKJ9O+/4TtVJr9f
6o4d40EjmrWxiC8xMAC+0vOiIsvXvxsyhwIsuXNHzAlTXHdbJ2PxEfYBSzm7
Whf+zQ7L1pnFSGcAMrboJAff3zHelOOHbLpTQGacfkT8WMOp1tq+x27/tc5O
jyfj5LSk9MvU6qBpa83pRDNd1vA+KafuIXOz1hf/kEYFiCAIK59+Nim6kZxn
KlNM2CYJFvPDy7f2KxYIPTvT59a3vMUPiecrwk987DjmnO0B0CtdWC8bQu1j
vlC/5P6N4BGcHh3N1cMyMaYijcgW5UxMl0bShEaALmXbHjp3dp1+VOtWNPmu
2RS1UuuNXDCZWfokOGyGicIwI06M5eD1vwfwG9opWCooKhFFxRTfFWyIosna
Jvtq/S9yCNFTtU3wRO+3TW8AIqwG1/5ryPsFIhZxXD/XGj2spCNalYdCYAI7
B+Tdoipx6bm/+wv3es75gO8KaSNjzq4X+38W34kktbzgr2+0KpLSMy6Q3VOT
bNVx9/PgkcAtpNluRmk9aWbj6bumBGP4saOFG8nnCK4+Km8w5AIFNMfi+uEU
hCI7ovca9Dh40dVLEzoWiCvTMusQxKqKkmaBIx8Xpaov38V5O4W5EbqrRfqJ
rSLus7jF1Qjt0fZ/EjyGV6FMAprk3oQZ8tBugFkUroxxHEVlXdK30JU2cbZO
PLxzNEuglb1O6OI2aOS6MmR0UPcmvd5AwJWlN8kym9XEXRXV0cqGWJStoC82
5LOyYiSU4pgPNE0UHPd1qvTJm8hs0wojRqSyP+6brsNEWPLDeIywV6tFGBpN
CBBX00SDdu6YnYBsdGPm9V2xm/z6Pqj6vvjS81ryKLmHbuK+DPBbcW0aiY38
rH2FXx24iN2JcsTysbcA8LBjYsR5Q7wZ7GCrcq+DOMksi+81OAtUcnX7nuaH
ujQTyf8GOigb/bsU9WCQB3AwDVAtMDqE/hZxTycYHsJzzrNHGr6VKmDm6UUL
FGZBy3xJlisancKg3XG2SrQvX5MSlir7NrH31oo49Rv8fU1nHSRD0NUruUuW
LWPZ4PHArWcpCP1bO2FTUfGkDbPSIKM/i0stkfytpMLlsusF9+MQmDwaGQc3
KO5YddZUAH1jfH+eyNvy+CPzLvp/HE0gy1dpitjatjINi/4WHgzAgZ3xQanm
tU+UVCSBJrHmARjNJWkOEcmaDRlPk8A0ce9L1E/KRHKi6GJ3wZUNQTXH/T21
H1u56JcZPjMh1mW6tmwBPZv+0UlTMmm771PJtfA4QPYTaLXH1TUwhFf6zoui
hxvwdKO01yRDnR+2hNyc4OAMtUIax+sk4BokI4iV+RU8AjFT6BgUsSzmFAgg
FohXBLjvJjmaX3jlwWEksbuVXTXkRC2kRzF1SenIs4Tvj8qbr+fLedq700wP
0QhutIXME3zrhUkgqMMei6MB1l5DWa2pc95uRVXJ4fyqc4hmwp3SNNfsvn+1
pxzLLnlbrFjsqnkebxHgCVpORugKRBZC/wKCIHigq0iew8fBTgNBo4BFXubd
Ew0qUrufD9CwFnSqfxYoS6TJhZU3x21gMmtCFgO3N6mAz6vWzau9nQ7jTony
0xayU4s0ChCtQfY/3wLcuWfgGkWaGoQnimPdtQ5HkrUuEE+wqeClyio9hIpE
3QK5HtxbHfNQcB6juqzmlDNbJufSk1RfdJN3nAeeVsD6gxRKwDnHSLBlGAvB
Jn0YQy8ura8y9cnEByf+B5BcJRxEvR2SM6YfuEO0nQBv+cqKgdmQ/kdMisqd
3F8M9MR5bXZiu/ysL99raLvffzakdRDj4TD9GUvCcT8wkve4TOeQ5BpbI8GK
Whwy/Tu0XSR2ofQ7URfQjcZ+B0LadmXHnDqAXbfTv1Zte5VFu1FirHkPgO4n
ihT31uObGuuZ26sC78/XvwBNaS9u6Ni5glul4IlNBzNcf6QwtN0xW5kQT7H7
pPIzgjL7+pehJ3vwmUejLHiHYfnyn7aUHzghY0VzBr98zjmFmzzJ6AbSDMDP
MEbx4mkveY5UPNRSfhw/7rP/Fsga5pSaqMse3TBAnysEVzRzYZUMO2lUx545
a1DMC/iXU95iotVUm865Cx+PaYTj9G+zdkXXL6uNzGND45f9ctbjWFr1BZ25
hPjJyBxKjhpT19f+5aqu2ap28hdt/B+1BaapkF2zxaLeIFpbf2Ta0JmDKuk3
6RKwtQkUFO9zWyWQsTFsnKz8umxV3Psh0OuN8kmJylDMo/ICN+mbAocRElVu
FWXXbKsba4KZVYOC4ynLa+D8u62CGTIltNrnWp4kKZoMU8tlyZRPhL6HF+w2
H5vtcpad5oQ/1D2iZaV4NRqSrQ31Y6HqT8tZj2xNKeNoKj247SQbItmO9H4P
nrtYbwnpxkcFhSIXM4R/cK5ZGZBdeoiso1yCJy93/fiuk/Fw+DIhhF81wNWS
dnGqnCcaCNUOqkUIfLypRwu0v/fos8NlEIWraflvM9c55+fBiSzwamlnGVXr
Tp5b7+Zh1KIO4EFfN/n18KEmcJ1mO/5sUHQ5bl2C1wf8sJO5Kj4aiVGd7Cp/
jiWciZSeM1QpEhBIAogPpzVTRJbCg1devjtmDf5MM13vKpbXAkKB1En7NlsC
LPhZaINWSWJ2fR+jjDQIK4U9xQ4x2+iuXxhTgLN9Fe6tVdXgryIGTf3nKiuU
cf4SUtlI7136oGgf1cjq0hlgLSnNVgDUwxDN9h3JERgKFMAmKjmXfcEICBVF
lvX1cP5nvk+z6Al86P+MLX85n6S6p3djYaeDQBD24opARLCnksM1Z0XNVd4l
sY3ew9LPak4P77cRaOMRLfIwY+U0+qY0f4MyHbKKGMurPwh/cap6EXAcAdHk
/wxv0hKSG5jYDPeNWrwY4MoYHTZC+BeMN4EjWPGMBnwFTf2RpGr8rZ7BaNJL
eYFn+mpeYPu0l3xBzDaeEcVZGbwEopIAt3A45j/5NZvJwzqNE12O5YLA8sac
TBZRmPYo0OPolLTjkJlPtQtcBY9iSnlLwPNEQxQ5pEP0IJH6ot2EBMU8S+gh
yMOtjh+HNbD3CnYxdM10ukkIKIF20bQPwYzx0m6WQ72mC2i7ew1ltsyGu/dK
Zrt+n6BcuCqDLnxg4CCd8FiSGfHrgOfGDjgm797lYpdO/ANPNKf8ZhaDFwgi
WeNdQ4hCSLgEHqjh6Xl6zwU3U1mtDKvyAj/QfBbfv44tCZkhWIQr7/KRgeQv
/1PS4QZsVQjBQwNsuzl2SXwJbGX+bF5rh/m6ItAL54iGchoix7owW/qdDWf7
faeDdc7vxKHVZ6AUMwdHiJgNOApIJoTzq40s1Jjo/40AcMAon8soueTrt7Qx
5jFakQxWIp94ZokyowqxBrmmt+1/cWKGDp5g4qEfWf7VfaBymNaQ8WxrmrfZ
Uydhu7VP0QhrFyu/HuCbeOr17ZYsNOqH/mj7a0C1Lwmm5jzWIvWnDwajWPCx
emmjacL1TdzdEQpOhhLhW49VrCjKW/ZTnQiE0C2dhhjntzCenfsMr1JmHsXA
iJQv/EkSKIzF8mexwhdyp/sdV5dh51Hb7n9zYz6G13oOIQwk/aiBY3sN5d3P
2gm9wpTr1OUX6j6URP2Bv+yJ/orAKvTtisI7Ndco/tSqJ1nYA5Deb6s/NQyT
9nRBa3B0xCFdzYf/dEXD814LeTN/Du5kE8uoxZ7VMVEj1cD5jw8HCL0066c/
EWFkVjDz3OSqrb+J1a1inGYBYlBW/eILzxyGtsKNhI2Ido78ydp+2W0pm3hm
ECUO7JUGiIPUPuF32BuW8ZFk1Fd9YyeBtJyZQVCrYf10xksOOVEu/76tpAv9
1vUhe6sXKsE+kEat92VsSQvK09sA2OYyf0AecH4D6EbWHShWY1VYs2yTlsNW
0lwRpO8HSzyuAVyQ+S8fN991T5MfLC278WXMMJLuYiTJylHrR7Vd1MquKN3v
HFeIF8uQbivKPYyrnKWLR4oVUKAU+XUUNEc7meQqHTwXMYXMsxeOERubE8cu
9/1EhWPtbQdJNp8hvWpyXSu3lIu5x/4M73spNsQw6AIr7ifFNmQkrpbR87jl
aDTQrCB2mHM+ItmdeoP1rUGNi/k/9lfJIqfhtdXqg3n9ICW3b+sYvusNthvj
620/RRbwY4qGjxRvh6Xnl0c0d/3LqTTKeYJWDf70tsPW7O1eNeaOeymE5N3i
mT5BQt/bW2Jc+LNNk5mKs6iaehPW09XcxeS74aWal398g+9K9ArHe+UyStcH
ZM07BCnxH6fShRXFL0Nx4CFIjfl7qm4HkTKPu6QcwwJXUvXTx87iyAEa4LdS
Y28KwDzT2F4DXyPdaw/xZFBwP5WmsXe40X16WyITXxDm3rBKzwfTt14fUmYi
OotBS/ivkPCeF5qmn5nrgr/E3FbhJhy+0gbW27AMg1ZwEBKDQ1vOUGMtRyUr
NVr48tlgJllLkY31e+Yru7GnahOMNSl8nh7hBx4jwss8B2iY1RSgdhRdBgJj
XCs4V1ivpk60QgVN7CtdvcUnWLqpKvu4jdVPeXNd/fhK8g47vLJKpat/a/6S
Hln7UnU9Fk3qLOcDMqMF13Ov2udSW/dw/xE1zkKBpaPwzxum/4FHfgysLKTh
LyE79zCT9lXvSgv5at3Pujjiezhe2336QiyawvK4P4sAcn49F5u0jfgBYJdh
Oqc40vT88XytwtYXT5vJwbWex+gQtsmkqHI8R/3at1f0LJoWl3ynKmVEYq9T
otMzlvv3AagXkpACzP1HZEZYk22tzuryZd9a5MW480AbztLfYlCxa/dVdbEp
Q97H+AJKdCRp5TQyUSNdNJQ7PuEGpk5WDV8T5OIn7llYwDIlh6Z+Sjs2+cVO
8mpvRmLJc4vPYyQdtjdKkznwh6RGrLEV0ygCmYrUSKVduTpWBT+/J6JZ+sq1
G9vv/XDG7ZxkGtA2m2IPQ/t15DHSKq0XiBVGu1VRZkHwPnF8JVE53gY5m0jy
QJ3Wwj5keE8anCGNjbCwWJSoRR2gdC4nAJl//KLI9r6sfzpgAhiyw1UgGNfC
BpW0fI2OTFni0rYoAx5TLtp6Ag3meSTupVNlaupVwevjnbTACRuuuIIicImU
mGyc5qQB+Ox7EEm+nXJmBWWFfosKsZIOFhGlESm5BGVd0lTt8TVk92uAwZX2
22tbT5i2lVw/yM7s6JHesv0Soi90eO2apUeqfo5sGt8Cd6vAC4hTSJ8whu9I
a8X1JJ6HZimhFMb5QL6Nnpn/ZzBsG/pvU3Q56MnhRZ8higc7rCnxkJOiQGfu
1NvAxM4Wjm1bpF5eZ/qOc/nzrpIyfrQthDb1H5otcbkb2/ANRZzC6ma5jLnj
Z1uQHdbnfnhG8CqEW+hKyENOwuF7W4ESn1KoeIAHwRlLOO8GMK/n67+X2MoR
g6EkPzBJhit5Z45g+zxdSDM08iHoM7/Sc28Fb6PS4ylxUc8OcGBzg45QsoIV
g6oD2R7dvUnd/vte/dW0u/zEcyGcj7/l7ONl3VI0X87XSj4qJvZV3YqS+l1f
uGZHU3Q8IzsK17gsgEA8/KSHanssbk6MxHZicpjEi7uLk1XzgApGTTqBGgBY
3tu/FpgTioOE060zMXDWRhijJMxJZWpMoC7QPva9MOEsQvyqpDX4n2s0/198
4bT4xNRh6gpEe8I/MU0T/ISws1LvBuenutUEU7igVLaoHQ35Jf+hs87TKYa8
y0PMnFLXlWTuaIb+SlqIz3xkuzv+FBr5lFJkeHbuUzjtAGmEPY6ByrNwJTQF
ZMUGHSP7GwLAaCNiEh0TL4QiA98w1JqAyouDiObpvRBqTQKaFfz/OgI7LtYa
LFGVxQsqeeXQwkKoKUNH7FGFNfaZAdQUWuRHzG3qSh3vMmPaDA01U9+fNmcR
7Y61LhILEYm1fX1A6KctURqYmrIN+I3mKsa6lpQdA35GgY4VSZdKICaR6QO1
6rKEyJ6oO10imU4n8d/ZxGbwfWTurqiga8U8W1eLwNG9iZYUMeUO+LO/xenf
v1AMLOWWCLtTgB5EfnU9LpY6b7tKQxLaStBTsHWvQrAOv+xaM24evoKwAPqq
vQz/Pr0tRs7XPzLwic+H83j2BBlqsmhwJi8xCvPmfXhQ2YNKUn9qQoFUL1wU
6fvS2bEmh8Su0NY/swGNGJ9h+lr6LJFcO5tbmbeD8khI9iGMTjpd/5sVjkE2
GeI3fYV0t53lctwyGCKUXRkDPHig5F5+l86P7xuV7Ns+fao9aTrQOajlY2ZJ
DQUZlaJoqW2YTtesDtwUdN3wwbH6W7V7W87wWmeDO+tqLcvRb0k9e5e1b3z3
OWV0HHp9Vh7rdCMBa3N3KLOc9qdFkMJ9d6VbjilU0YiAnVdiF97SJMfkie1U
w4fuevnHw5oonMXKshts5RU/++LMsDmzWpVJ7LaK01uIwuoT71Lh4Fh6qtqg
2bDcqu6oIY3jq0YG+RmtyVgOf8LJMmICX3JGCHAQ8VnQvtTW0RQJs36/IPra
DadQWGtgxKccg6zzXgEhDlz168JmjiPlMFvUMAF3mPxod9psyV1IWZr9ZIXq
TbP449J/VwMIdJsT3oPNY/S2MAerI+LQ9UB4LjfjPTZf2wQA1OnbBz/1NFad
JIL1JJnvpuTbGTXlsKyheawj7Ed78U7GkQ1Hd8VpKTGwzos4wndrC2R+0uEU
rs0ELQ1xxwt+lvIWWMlOqqogSA5l5e7FiHhNiwabqHqpnEb29PLAkeXD7DHo
XZorCCGri9ZWEEZ110s9Vl4nlKmCFfEdJpXgMtn2nsX/BGVsuFOcnKlQaYLi
F9Z82EKKxO3xunQh+zI5bss77MDb9I1B9lCt/gsji3RnqaWFNn/LTTKHDYAD
XRxBSehjaDbCseXt8BeHo5knaSIFfmFCuhGa8qUDEHfbFC/JPBiN5XJx17Tb
LPB1n+XOrgRqC21YHpUp4Eu/WW3sB8mmCWjblwed+1CJOdjM1IKz56XTrwa4
d35VLVf1EAlVwlPSEtoTNjwaoBFbH9WFfXAGyracQpEQ1mOeTlodL3z2n50w
VmtwmVDT/Bq8Zacu3/zm49d+4zEukz5DN8ecMBo16PDEy0Hv0uI6LQ1f2gEI
MrLY5WIX1urgmUodUOswmp+1zAt11OmPseL1/KSfe52iHsV0+IgLhOg2dsAb
9WPvGXSPapHV1zMCYJRAvflPlRrGG7WEUkbdlst+9EB1OGpv3imtPCvg1JG6
kBAqvIXwHt/Ehr6GGFslL7YQ2CLQZdsroNNbltCmRZXEPew3depzXCi+ezLM
jdtcDsCo5YcmeuVW3x4KV/5Gy6Jef/BRZp4pqDvzFtEc/H20+pTAAWPldHY2
9jTFHwHN/m1RkQ2qiLb3NMR1MZUZQoqHK/jBbkyToPhC/j2x8a9UhtAChLyF
N90/pbiNArDbErBaG9hi0oOE7V/bs2ZHoVdkLwGOo7ARyVX6lKr6E3M6WF1h
9omZ/3aGcI8Oas6XTYZrwl6K5LNByILZqRN+O0W3AqRXCcrFiT+z4YEA6F4w
wtyFcRScMSUu//4BsAsYosxfDpUn3suihuZARTLgTH1v29UkbPWW63q99aE3
481FmQhhuQhupHHpKie3vp0rlQGKtmTniY6dfzaj2ZmVYLqfrTyRh96spH/Z
BhHzcjomp0t+Omx36b9VQUxjlYziKTS08DZiQ4DFEppzHPcxDBmumPfse96W
zlZa+i+dUPF5yF9XPqAiDFeViluBSRnyfPgUb6P63HcP1i0qxbbn7ozfDvdH
9Ir4cuzetuE38Qry1kGMM/AeXt7ncu3GIO8I7wWy7cZOxW19XPhuG7xMTh6O
K4wRaAK5dGBQ9vIT1pNAnKRfBxUpZXqEjtcfNoooMr3M6vO7H1B6wDFDtCxY
I8snA6ntJrnveMBvkX3dMreMZCit9nsknP4CWU4ELzfWpPmHPqmO00GYUZKE
euJI5pZeq8hPKy87i14XK4oML+pfGEGYREvnUbzgyRlNhQUzQHNIOUpNvon+
5HlUWDr0CMiRKbNy2e3f9OqsGxCYfntOgR7R03YmkKUncjLFdxcJsob47/ew
mSAC7hss9GUtQdM3JVQnrXYkg8K3EwMkCWOC5IP3Id1pQ9dbeIDyJtHjl7Wp
xgAQtz9FiCjtAxAWuGEm7NJElnBudI/5Ui73raGULHNb0NGOp13boRc0CsXY
nGHv+Ha5WjtyswLlP/asGZ+BO48YoE43H4in1MrDuHIB2dB1S8Ok5qPKiEBt
ncIs1CzjazL1g6lw5KBbc/8KMbsGTalPIITl2SX94XUU5RZmy9DicSY2aeKp
arHm8EcRkYsOyKHm7i4NWohpvR1bFNYgzroafMNzyGM0+8MWfHZvWcWKgk3M
h7wLCQLBX50UGIoTrUS0wPPhobMBnFh0X5ahitrLbLb6bK+fUGCgPLT0YizZ
HiwBAxehxa8dom7L+Emtf6oOjJiklvIflTjPszlA2buTh4qpsoAnNdi6ToB5
D2DigF+ZrnMRoxStfbyO5ztwxR9jsoR/g+q0P3m47rZo+5c7hZytf5+ce1Bm
+gx5XhJ1xkiLcVQxGOxARwCUw6Y6MMkZm07xtLCi8usmzJ46NZ9yt+h4rGln
xEBvHW9KQhXS+7PWSU4Gz7nuzCWE9D63Q7MYwMlccsobrdYqexaaGa3hl9cm
rOB+bW+AYZz8v3Oua/wJozqWK9zjZF1DcJJymBSSzfTyFUROBPZGJuc23+hs
GgghzvxT43O8Bm6N1WqafnA8b7KaSWKBHbqOpLPAWTvTvpn28rlxWz3DU8iJ
vK1NLpDz71cuD8yD99ThoJf6gI5Jfrf7/oXgt47YJtTvaXdJWW4vnyFgIKGR
4/KaLVqGHCo0Gh6aN3TRhXhGSItyz4OnTbiE3puMWkCxKEqNJde2XxNG1KiK
8fmvEyJSuedVZs3QWKquGY59ezIaV6oke6T14gENa+bAY9M9uKbD3MBMe2gN
09ZX8XGyPskLWaykg5aVtMxmErPC8Q1HdWVGizK9Sf6wB6FTkQ8aVCEyOzLz
Y3bPDii9WVhJ6dt3fV35iTurx4BPYmW5jROneqphx56TQwQKCjEMY0MfmzAj
Kmhcycj9viGHLc0tqasSZd8QmqQjDPSxVQmfrfVOVlN8yzdWwvQ3SFRfpsiS
QPo5N1NlazYYO1h8jsbo9E3RfNIMOXzbZ68vpeUK3iCEbJXVS7fm3QFhiPfJ
Gso1G2VvKU21aGNgZCZQHp1gCDWWhYmVFNOFZYhINv0XeyNUUNcsQTyMgtCw
HIwmB6UV3dhxZZjYLdU4hSCT2csVccotXfSGQSxreO9AlHkUtyT1niS0nj79
w5fYcpFWVcK2D5+/jpO/iqzodGFNSoK2Nkwzy8BfKWeDHes9jK1gDn4T5uFw
hlh3fAuZfOi1j2tRWpnGmVQJPZM/ImOBI22wXWXal86FAQ4pcjO++ayRM3Q5
po0sPu8LN5PIi6xJNQjSZ8Fm52LE4dRdQHCA0lEWwTb+54LX/BW0fn8z+JKt
OQfzU4cSLTyoEaUqSdAiCW4Bomn6Gc511WEoYwa2Y+Yq183PpV0nVcaO1YYf
iiZR1ejAfaKWzY5uO6xu8ixSZkC89bec04vVZftm+tWw1PC/bodhyb6+fZyv
nJHvQKcYk3W3LhmTvazsfZCOd5GroDMscf1mby1mMd6h9/t+oK2YdL5vxETE
Qm+G53pkkeaU/kN5+8tNnwF1/t0Sb+uNQ9aBJoiNo5W3hcOajz6Vlv+b6Ve+
ihQwJxKXITTVSjqaAiQYW8iQYm4j93n4pLP3vs4yO8RqG8VL2bhKQv5+JQ3w
Zf0Nvzat6ZGSe+xujh3i/4ZOmzJe1z5bCa1Cu4aI5NDlpu3oTycuBOT6luZs
5J00WzPEa1P+yeKPqqROQCXXH6H94sHPsTJBH19XC5Ap7wAUQjCW1NuUbk3q
Ys5xJDF+OPEAxYCL5pXLei6g/NL+AU640ygWOqrwx596P8dhOEuA/eIztwVL
K2qgiX/X5R47ehmAAa8oPLqd2tTcLt71xwk/vr5duFCJfvgKekECu71Q87oO
EjQPeY1UzBH+6nRXAsGpGVzv9qtmXnt3ccqNycTMhRLuUdc310KCletbojYU
vfItl6ujgZUd3ElhexruCvhA76kYcPcY4CW2/34YV44VweHlZ+znWySXrLHo
nVHY96RAyJqpOllxEQyi4W3IqWEATAXBwyWUqPLwwBKlcwLoj60zeXcyzF5i
kUMuJ5E4uwQqzNb/MQy+wujPJ3qNslVqGbDvG41L1Bgifgjq2VH6IJUdURrC
x5aUMWHlFSKbqb1n7NI/D5Yf7zYiEtuXPvRKVEHwVzrgKZgskSPUjpKza3fV
soq9EIqNKmHt4FU/gPz6/+L3i/X01sTBQY1BXFT6oL0tgWJ7IgQ/jCL7ZX8u
WFgGmv+sXHG1C8X9PqDWispi3tC8QP0znd62Vu8dctg7TifkUUfVbyiUm4og
lxO8Ufgc24Eghphd2z+2AMkDt/2lWspjIYvUkI5NCnHlk1Hm/QxLauTvqFwf
SIRIjz0/4MG0i3BgexFGvjiw3bh4A9hYGArE/J8TpjzAAbd/A9m82tBQl5tQ
fQApDgXJRCVvdoQ8R2vlLY8qDJdW1+SKGtBNbBb/K+LCJXOjTATqKAmRGE4Y
EHueP+wAs58SrV1do7Tj/PHVI+75GWMTj6UCg50xosPo993WljrhTwq+kLb/
A9hlhqrfHxWaklOLmeNOXb2C/jKBCl9ozaYxNc/ZDI4Ts6MSFiDKLbrU+y25
xHw8ifnS7S0RU53+++xqHGjqH30KJ0ODnRknyfrNXqzAHWpZ10An7asiMo7b
lceylifHAxW26jnhNZGqqRZa/EjYpZGOZIiMZFnxIMZeXE/SIeFqIyh/vcmB
cFpqFM5NDqXaI/LC6HZGRgxFJJwppCMq+qmBAjSiFwfJlbDIXPt9yK3a2zv2
Zvd/8WGpHzcU5RI0lOZ8W3vYpzPszwQKDfLoLZJOMgSLhjaBTQZSp67QsXNG
yEZ8skzC1EHTLTTtn5kY1Gmcb1bZr7IULq6J3fdwKnFKtFhJg555xozRoUIA
ZBYtCsCe4OP74EVf2/xknDgu9+t0k9W5tlevaZa0QoKa48Vjex5vzTOLGcEc
N6efLEJM2ANWL0UWys/q6N0nb8ORub02jdjoYkCcWFWGpZGFssKLNoYBhHOp
y4FSJWTD6xRs4fWESNqfxXhHXuBSa7nf+bdc0TwOJD9GlwVeVu3RPlgwdL+5
CbEFi/BUAgg0c3nRgq+gQkZwRnstD5CRdIgdWUzJvh6i/4Lt2haPdJEA57W1
o/oPMsbLiWFoY331+poVta3WdJcwJ22W1fAWv4L6lnwh2BnNAydGPQGTIq6a
Zc7hEmp9GnEAPMn9Dq9r5X59aXQr1N/s4wWo1FRKOcjAcgHd1//HLTeouwgp
VhR+li1wSvUN7ofqgpNZRFS9MWKyADMIQXpWwD16dQj+WSQBlN6SZvVWS8ZN
lfxvoRQgcHFCKxwgDTEa5RMezmgyVWyqFb+xtIlTn8YviEk6Io4ocMkA4nmH
4qO09f6ZUmySfCu1iv41g7C3aTstFTW8HhzTpb/DERhPonHDDIDD+Gcuwgss
Px349GiErbE+yZJ5mdhck5p1cyqZPhfnnFdbz+lbLpzbBkU838R83FsLsXFy
4jItp/tgQikNHBvlXQyZRyF37motN73uaL2Z/4cIUw71gHH/Crh5fUqtYySh
U24RFPrCMIH/UtGQPNP+CLlhuWfmGj7wAONWlr5+zVU8OGkvK81tQdHq+FkO
Fex5+qsIp64Qo3grvUrTKPk3qudtrm4mXjPqCfUWbwKvpYnXxeOrGiV9cB+K
lFtXhWKMWJTfvi2bV9Dbp0rB6+eWObynzmY55jXuvGB+QJQzN/qBuPdJK86e
g6BrKgO9/uMNXm06Wef2hiwZa4L0hwSnaROyyNvI0xVO1wg3qMYj4vOTMiHe
jOVoQuZPNWEkR5tSX6w/VkGDA6zx2ANXYFaPAzYk4s3+btohS73PCE4rYoqD
iKijLLKtqafZKvyyhcYmJr7VYpp6u36r0rT2ZMcf3qzGVEXqMP2WLaQoKZ0B
MKXMJfC7M6BPnlnYveeRDYciesuNSOCqvQyDvFQ30ITQpnuFllxEWvWGQ03b
Jdba2f4C2GMdwYhUSIp5O1lfGUH4OJkz1hOYCtM6KUx6TXizSQqfaGiRnGp7
L01b9ygwHaw/RD+hNXhOfIswfuFXA1nbaoza4gbnoeh8oyVw36voM3+6nj9H
fBb+4E/ejlitWCnIJJnUAExwS+xOnNqx0vHrqnAMEQlLxW1vJbzVCE3NVn+i
lFB47Mfkjln2udF6LWf57Nni1t+46dBvGFi3zA9eH+TyJr88w+jkDFax5pS/
XtetY4OXe98ctRcE8IGclGCyyTf8rQ/g+4B+LJLKW02+hGEVWgL+wj5sbo7L
GP8nkBITp9VjKl9aRxxGj4mArUhvVwxPmzEPYMYfN4+/mujA/Ih/xea6SgkY
FSTgapsQNdAwhf7EUjOq1jCR8VDuWP8ODMYmuq0qDUUj+0b4OrXKRRH3HKmT
eJw1NKaKh55E0ORpHNSzsPzc8ScD4S3KMXbFH92dvO81x2AIMSr7tcSG1KJ0
PfKceR8RpZi0mqlGM0KmOvSpY/5nie0ZlvXCY/a18+iLtAzz8nzO4zzMrw+B
me5+YciFAiWZQvfm8+SOy0dRIvY19FsY5mtFrOjEwLocxDIePD8DNJLOhoNX
54eBKyMQsPCi82Xped817ZR2xDsUqXOOWkzbNJuVTCtCs1wAXwqFCOChwSc4
COJL/2TuTzmDATiZl/p3RjfgGnUoNo64xGMWtyWZk9Kufsvsl9rkizcixTJW
NGtueQyqjXZt46NM56I5hkxwwxuPkXRmBi51vuLTaoXe9fSF+mMhW0zVk2Ed
DQArDKT7OSBZBj0OsQRg9dAsmXEnBuY5mAKWgDM11I0CjEgYqhujFMIEt4QO
DY09BTRXbwUYw08w+jofp2N0bGam7chkuiHAy5wQ/fvk7qdJfCjM2DQ8mpbJ
AW7xjriiHcPvWWXqUfBjm2E1K8ZKJcpL6v+y7BO7Ec/jJ302ZkMGIWpLUR2R
p8cPrx5o7X/TPJpf9rwrPaUk5sQID1uiHaDpzLzQCS7c2HY0L+0Y77ykBiRb
2X7RpMCpckE07Io/LSXVS8qxMbqxwqR5PlSa+akelVX9TVeVq5KqO4fg6tQF
vgjwyX/Ac4/rgdewxBK5+getKFeCddjiHZRrVzRYdnJy3cFyepb5BnUD7lJ1
pPWAAzg6QWtzkdD18peP8RBnt2aP+mPJuS2963u9jlSRDcEj6HUse4uFx+y/
TZ+N2d8UfwDr20ai79+Bjfag0AAGg03Ia/0q2pfCWFW5ef86MQOv+K8EJ5O3
g+wGDXZYSbDSauhKbKzCP7Y4Wn3oarZAEGtrOoU/Hx7UkPdkBsXNM3XI331W
f4Np440nCFrJhHQjkemMReyGAu4tVaJ0zUtVZDy0f0OEkHbH22ZCI7kTsLTG
bMkZX88AUgTqR+Ond0A/Yb1oFItoCcI7o+pyPuzuA/b9T8MY/ioyQ+10rEHV
1FL8PIV5wo0oyvQn3WNkhJzpStderobH/W4fwnyrEV/sBFv85d1yR2B1RD+f
zG/8+cJaSCs9MvihcHWq/oj1mUHIPTNcP7FMh33jX0SGzV/x+1r3yGDpD/Md
wMb99WAzPw+0fQ4bvD9mIhaBDWdbdeS2GO1RYZTXqoGzcNc1Q982BU9ViJv0
xDK4hzhb5Hue77YeiiIIOPDlijcd5jNyYPCKvi2RLZYxMUHCTehcc/WhtWYJ
6bk6CUbsmbiEHTXqO2l539P9I0EYrjxRRyPzCMF9OlOKlnF9HgKE1oGIHeNR
0l6Ywng5VAw4FTUA2+tql+nzdzWZM2DgscQXJjBSXrL4HlaXEo76mcIiD/Mm
leiLw/LbB7R2DGfPwKti1a1g1XtFB3ZD3tT4VRR807cpTfpU0Lzhp0toqvYL
fhI0LtOXVHgjfA7BuhPLWMpovop143jaDkrzfiK71RHJPDsYt4Fk5DhxWdoj
cfEwSdejN9kuMUUVrKKZFrbnNEJo2hTEEeRYB2LGSidvpLDz87klBYC6CtPx
J6bYqvv6XxOQ0BB4EKbKIuOq3tbBiDuXTt0oFNk9emSmEJDtSZ/kDE7JQe8E
bDsbMgTkzwt+ya24gk8/1n3YYcSraia8PDteYwJ7mJvU/lszJ2sNomvD3LPv
o63E/zKRfhpC+I5UhTXBtlOxwJpvJS0t8eic6gIqln+/BTOGRdDW3mSzaifp
/ZW2WrOXlvv0O/Qt5NDE/og5mJWxoX4ldnpj5TDc78ERrPsWoJy8zMk3Y/QN
l6vuwHckcyXA1we8NPsAqyb/oEQqGArEu1HnmoO/pC36KGofzeR0gI5kDcmq
KaqLKtvD05C6POSaRXJY9JL7AnAzDXtG2RmTufsiPK4tyCb4enIqQl/koasy
aIeIZ/rmbuzGO9cHWvbINjcUoT3vd4KPxRfX8BWoA70oEPW2ffzwD52UK2ig
iqvj34ZtmT0CxOPtC8G9BDgb2XdUDX7USSIYcbERqCz1NZti/qJKZ9boK9Fh
xHcx7ILYdfzPurcDksp8nW8zUBS44Ptpjc0e3ymLjTl6zIzoCj/yv6Dyi4Z/
cyF9Z8Y+YJQkNt/Vl+FL2b1a3q2e0LvB+Hpdh6/O+3X7n+lIi0z+6HUEfBVd
AB58qxWT9J3/luia+gcM5w1b1P7Q1DoYOZQypFT9JjT31P9aQRMOl2GhVRle
zbpWE5QgmzJ9pNe6ycIjgaXNRNS70wV4Q25AyJB16S7gK86v4TsTBbs/QkIt
J3PCy5q0ZOl7JQXKpitIvSC5aLqF3kz6tQEo1RuIpu689k3eBxW8OZq7Ac9r
slOlbdNrmMYUcBWF9ohnWpcHjFO8XV63zlF0sP0MDHk46KY6IwGVY5YIhDpM
n5iOLc50dudEN7sZv2lvfMbPS85OrRnnz/uTvp+s6L4+CBvMWT2FLsSnUsmZ
epKHf6Vi8149HbQzbDSk4r4gCYbLqZ/EYI4Y2wsR3a7gBVd0/WO4xAiG3UTG
wcV0+iXfo8UOYqmLXdk52EgnYLpfIUmVjyh8BH9eXHg7p9/dUJXMwYK5xx9Z
uJ9gTncW39OUfeO48NzEw2A8VQsIE04+VktZjBXAL8k8+0+HnvJvzDPomdQ4
U1Q4dDKSs2Z+4YIz8T3RX/bN8HgaFztDBjGZsxueWxWowruNz1OmRjUeLL36
yUb5DsSJ0ZBjLhARc+cJ9y3mLRyg5Y9Eys56prJJCzVpfX/P1IRIU0qSgr+R
Dg1q/ClH3WNJOkDvbiRnJoC5h1qdcdv9wqzMlTSOjMV5Vqo77pDzIfK7BTqt
32MTX32i6eto5nu3ZdodLhHekpypL9+5vS4SDs7iIzYvEGZKByUUjy12fr6h
Tb9Af8whn/5rADn+1ukNpBvFtKut20yfr7D6xOg4aoKS1M1Jd5JUc0q9IFju
H7CRezYtgGNrZ3Pe87pmSZtsfmJ3XURx98CIhUOn8iRvsN7FEiHzUh4LRsr0
8Z//hfXtwZrehLkSROkDchJZR/IDUCfCs4TsAPOQNjEtBJsGcLMMf6oCYJwh
E5x472kR6LUI+sPILWpbq6wRs95MOHRRHbWq2hT+GM3LhzSFwTN4p8qMnrF6
m3jfqTctyqr+i6ugbgqHaGdiVOyn10/NMJzRo/3+AwMUkt+d1ULW5zBU1wER
7e22baHtG/hFVHBbiUopY8cbC91DcAVciE9VgwhsD6Q3BvoGEv5pZP2qN14z
GndCXBAnyi1tIBXFFjulGf7tiwXm+r21TZ3BY5y86FuFUVg8pScZpLFmlrg6
V+OMCFvLoN34ytFCic1Iew7wkp+SH85u396Dnsjedj7B+o2SHrSw05arlybO
vVAph1TcTAoWs2mRXzqCbRQJT5cdJLpn/6Znfc1VVO0t0b39/1Hol/zRsu1b
D+LIjiSJBTVRG809bSoYsVZmBFz9BSIiLFcE8kL6sUEO8V1Zu9EsNUedUQXe
dni1PhUP6fPIaRdoOMMXjvM8d5a+Q4YVOjj4NnlKxhcLR4oFSc0+iD3hJdmK
wUbKx34F3bbmjoERio6oS5CiKqnQdhkOUf2u53SV/Zt44ogG3P+gIbEWMG4x
s3S4tZPn+heq7VUMw5nRpervLRgD2ufMw9TZkeRVnoF+ZRnFcbQNM7dYOw8J
f0BQY35BgfhHcAZRmqYvEsJzZYk8Fx5cnqVbje34BAwHViv52XMC4o+Py0+j
ipRdiPmZhrdnoCQEf1TlaoetWxmx7A8ULnY7//0pIR/fVr96wCHoEjK40DgY
/wxfWjTSWT0GltXo9HL+0mVRdDzf2YKeHmWnjDoMSIJH9kU6nalXBDztGs1g
l7hnBp9Yf+dibrFVcKohd69f7p90lRZUkVBCgED2naHmelz6L8ajFzM65Qdf
KW3AyDlJ4ZUTX5jlwq2dGzuPcMu+igVFXxvJMsFbYbfGXbk1JShP+S6P/eeN
Frp6XNBqRtOG3hzwk+baIkmneEOeEHdFPtO4QXQlbPAs4PgD8Q9w2y+sUb0+
/EaPwqFc1GsgmngFtWQLu0XIKnbgwFXzhL4DXV/fRDKYYDWOhwAUy5eIYwVh
+Tmhz/RqHRPrADpMu2nhXFxXSAHT/pv+T4bnJip3Wa+rmJO0SAU38DkVQ24q
aafACtqXTN1MdTmljbUkkcBSFktkBrx5me5kNkmtIxPPPKB8vv/wEQlmWPgG
UXgNZMRukU1vJWJHYfs044dsYJjSyvJQ1v48tlNecR/ScjnOcqd5eRum2tas
Av4/+Xm8OPlapEWkTceUvGSZGzcwl38CL5iEA3Vhh0/z/t+BdWMOLN9j1dau
B2FsoCSUsicl77FzydbMUAWVMOLwRPE4inkkefEQLzmjYUZMps6W88dFTWTL
/O2ysxa/jKlEiaZICAUrK3ObuK6fFp5g5WIMJyB4/dgwkWysiFcGkFtcRDfA
3p3VWmgGAevxEDAJH4931GdnPF2U75+ZhCPArIpnQttYH2jsBN2HP2Fzs/QI
5CciZQjmiHvH3RQpqte3DflJGGMmLwdjowM671yUbr8sXHs23GkjqhsJyr7m
c6/hw6Mr3Tjp5H2d4cbhmKwLLhsJTnJK9JmJ8hMGgAnUvIzGMxtlT9dNQo4L
WawHsbFQImrh4ns868uUavME61twxUsy4MIvexk1KOc5TeixHd7kJruY/ueK
exz5jsX0ntG4reHJF/biTivGW1uPyDrayvJZHpg5RM+fc8KTJt5duBB3sJkp
P/VpyC7dbQGD2RNSBa3AqF1cA7uz6Drupbk4oPxBDbT0UJGZph/hEpNdv7C2
r20u2yu/5W15vsRSXG7CBcwOkx/YHCC7Jf6F4h23FGHs0B9XA/NbyDZGmuVi
bu/pNI1JpjTvB81kVsjhXftSPo0WlH086VEuU0f6s2QctqmGZbbEHR32h1Ns
/uJTFgVyGDWp4q7nT+L923tNnGinNQsDyWJqluhtdyFHGhU80ULMbhGxHk+3
a09ycDBzcoHfm4v4g2W5pHLjYkYjHoLb8FrkPGLFxq+bH12e+m1Fc5vsVmqe
vFQNrwqxHV067S4sTjAh7TtZY0t7yYclhqgR4P/xy74/mbw+SoNE60dmoWzQ
F0LgrWTLwilJupgw4Q6yzFA4JSL71qwvrhlJ0xlynRmmy+aW5Rkn3WV+5cA3
8xXX0CyRVl6gX71cRDp7nwh2HR//MColKxYXuX5DUUb9DCWDYuLCZMnhUqjN
FGtq7IhMm2zDhqZhBjntHDJ4jdg2zVPT3xUKIHTKaVcxUpJ9yXXFLwkkw/4a
RwWc+Ul+Cqbu+npTrBYBRV37h1uzCCUSiMFbU8hUkiCR9CZpnVLIdCODoXO8
mEIf+k6JMUt74oOarsX9ZrIDaPLoCJKSs6s1ZRiSuM3aNmb5mwUdOZsfhoei
S7TDgvgJXPnxC9MQMZpEBzVz4CxfDVybf6/Vdz0nJaaqdEYUHvbY4w7mKW+q
kczrtkLG1krZOxMecYtUIjB/q02yUbL19jUBTHne7xEt3BQFHw51IHxXvJ/1
+jENE2MQ6oOYvw5l311Tk9Oe4BiczNcTB4G0G/qVlGphKrlxfAEaaOlZqY8A
WFwf0vb/ul+r7yfFgz5wSQNxY1eZM1GTtlaCXJ2T09eoUhvBMqe3m1Lr+uYJ
h2mPjwWoAI8wNLCMzDvnEdR0xUPkYpRqQIK/wZlDrSGYF3DLAhdKHSGCHcd0
WAXCOi4TuEOqbo3ZiLTSNkB5ZRtdxhlvAeVZuzi3EZJ7IiVLCNZPP27ONj55
+/IgqvPvx2U4DIxoFsmjl8LFDffFZ+T+/wJrtDGOPo2bPGwLw6VBQp8N4PTl
FKDe7Wl3i6NC+zVjAWjRZ3uXsAnc3p6FwoqG2KDvvl3tbQXrWEU7Ujm7CAJJ
rPyOs5DSxAN9FF8f+SnN8biPZ/TzUwYfRYtU5m1p/Qps4LtebU3jTMVC7NEV
wTR4qElE34xRS6tkU7YIjtMFo5BcwCNR0rTLCb4Xe6Yo4BjM0SbxK423JvHV
P4bxXyiEu5wFT00Ge/cIoXekX/k5sjR3Ff8Ta8rhKb+E1PPh3yd/ndssZJUM
StNKPclA+hwHG/KowxdsibgZIq5pP438BolSSxEyytAOWgUKY1iV8n2IAK3R
g78btDRyOaSwxE9dofquuW8rCgKdh8Zj8uX2+XWwlCtKPmWw2P00vdrXGYe4
GMcFmwVVRl9bVeQPMqWYXBRe1I5C7GM7YttcKKpxJBNAdiqqQ8++eQ3cvv8S
YAB3OWmexlSQjyJ+nG74lnmtgMgO2TArX/yNzhFFUG47JJlrg2Fe3waUzpB/
ZvCfdzZhCFcv9L8AoaBlQxYwokrNBC6cTvFp7/8iOz92dbN9n3TOOERVRJAx
nafcVE1gZpbcexFDuMLJIWy4SncfncCrF9Nq2s5qK6otW1gPIThWw+NJt0BO
Rvef306JP6eU7bUFnFmwClYKdPAjPwaIihoPpuvbLXH4A2t3W5uu7xPNiNd6
xHQRvgyxzZ7Gd0UXKxaryxPBbjBhbvjvv3HDmeOyke9EeFNt1qu5JCzqxKjn
oBZu6ygEslb/ABOnBRGpDOtszCfTYFdAta63zi+us6GEtMWTfF3CfNivvQO6
cvT5hKpA+KUHLtxnrVh/mqsd9hGcyQ/nZtU7nPSxHB2nEWbv//M9ImBqxE/8
jpr+4RIZJfJnFFvyrbj/bDG2ZM2WfvrPo10CgIMpOLotNdOjsMMVIEkJC29D
pargpti/QUCPNtUBV5ya7xoY4h7GMAgBrKx1oD70r+qYiN8apsfUMK7xp8k/
w/ko9zlXPn3SglwKujj45oNFehPjW1//HRfPb1fUziY5a5czQ7GhrSaRp/27
WlEmAtVtfPHZGiGUWWtvwCjySmH8sah9LXV6pvloxuGjaC5RWKfoRDMW8ryY
3EwwNt4B8jdrLLVWWrjLGnhjmhjx52WzSN6kGB8g8bsbS728usuF30j7balM
Dy34jQ9RzAMPHcFYLvzvM1aRljvA3+hai5Qk5kqbCWxmwC9keHo0Zb6F3ulk
R0ypfFBn5dUntLsnjD6WesOC0BFXlu37K+niZxvHm+SG/kXAbldLIHuMeFz2
b/q/moPBB7gsYd4RAwVpXsXMm1/4SJZ68NCx6rr30JQdBmbV15gla0VI+a1A
s5baFE+Hkq2QBuw+zYjDnflJ3GbCu13PjMUYzQZ9E3QWg85fYWtftrqTOE5k
Se/oCAEkiF20C0313FJ2FURiWAoRLwwKJ0+Hl/ppBjv01iAUrtcNLechHdeL
DIHv1aSvio0MT96E8TSYnR/fmpCYF01VsrjR0SWK3q3VBkN6hhA/63T0KHbA
4AyBFRrlHeJH2HYbrbQM4kUBLMISk9BfaqN4tyrTm7KT4MWaj3+7F1dUKL09
YugTrLy6kUs3b909En3Y5IugznFxgVRQdQ2Qu6Q/kLoHrSdsO26dJGO6kpJj
BXtvcDP1NxtLmOL9fZK+2y4mIIpWMNFGd7NF/XknKPRDForB9yldR/DUwRku
QjmAY9aJg9PSHG/O+YHPmfIEF7t3kSKlBUxRAkcciGWFWdJymzqpNRogEodo
Hw1l8mBFNwx1yxs7u5Uc4my4LhoZk+QinWJEDyJydnTmHk6nNlz8DStpKUdK
aS9I6olJKWdgepzCRbzWYdm0IonI4DY7jPjPgNJ3fNQSqafdK6LtZvYq7fxK
bSqHbPeAu+UDBgLMuYJtM0Iq+klZDSMknp9towEaoKMpR+XIlcdKJgfZi3kE
hHEo8njQuXydgGyQX+G7sjq6ekKqWyNcKrZD4Zv/1R0hIP0ldXJBMUECB9+1
cDzgnLRjtme8IVbtG1rTYfpbHMhBSZV94PoPkRG5iLSCcY1XmtSPpkGj3hiI
XwLruJhgTstMbhIMvdV18TTBoO2Cb6Wffd+a9xUJUhXsw1524XLHusg3CPIF
COIM3lfvjAOzmZKq+ikc497aQjlLavF5n4yFUkFT0h03zuYromnALUxggPDw
/5AOVPuJdfPzNHzH5dVEFPLX0BAb6bfc4qsAf24jSoEWGK7LCq6Php57rb1H
ONKuV4BTU9+7USTAtfQfs6ybMHIbRLIshVzapm2dznzXc4k7pNybfD/8VRtn
Ty7aM6NU97iZCxRlA31bWLgHCAK8//CVhc11fAln+qwt8brO6SVwFTs9J6dh
QM4EEOWmzUZtnP6WM0qHpurzfua+xXN+R+SwNSuI7yjCXa7hS6RKcqwV65Oh
W7JXiGLqFvvRiTZ8blCoDRLM3l/x4ANXZwiBnSdJTU+ZjK8eRFpDi7oUJ8dP
CVtDTxP8rQkPs74D2WnKnk72CzAnbV0JcsWNUO2NJckgGudLQUkwk7Zxcz0s
taaRp/JbWG5I4s1JBPCAsXdisEvbo/EGnJ2yl3LgUAwwajVGLIBHU25mZwgs
Cwe/y7LpEKVejDPGIGE++yjfpjILWIJjIG8i22heGPQaBj21EOEI1IGgCuQv
CsmwDPwYAirCesCzzYDGm0kKoCp3fNu55E0cTlX4pU0blOhO3k80iF+FlkY/
lggCEgripeZhZhWzo52h8x1XGxv2vbvjKtaqVNjudCJTVsZSkZqlZLE68uSS
t871NcP8F8XxMizGZuojBfWaWpl3uvBN7cuqaavFV+QzUFLzcDUHo+zO5Px7
10qtf0cRUKMqNDXpdX/v6YvHzmMx4gtgWe4mhnzGvFRm2oot5m4oQPW5nG30
V6OMczLl0YLpdfWz6CC7F9Z+ielDRYD30ylQl2bzJ1ipuqcBH3TPCcd2/XYR
ZHoS6VNrZwqdiGrGSMLxbX2rCxkIJqJIeKC4c6aq5pwn5TNg0EFS9MxcQJgV
YNUVUBlIHkJR697gGMmuoVM6PCd0GkXz9Ry2lty35u4r3FjZBacAnm41QoyM
HlZtxsH46VkDT/iZeJPuRiRMSfKwrs6C4e4ph+VhRqWeI/WweujtOgbrVdh9
0YzaVWR+ii0ttzhArpD9cwI4pIwdNsggDmJxqIEmS0KBNP83Kg==

`pragma protect end_protected
