// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
U4ktkxcTF5GtEZf9EP4Oy50+BgZN2e/rkoeLg4UQW0rC/AmqOMGmcjysDJF2RfUMShWF0pi1M6gN
wmIqb18m2w6qYkhlxgYBW1ZVXyXmDdVnGhAmubDlMoyrJcnhevMlw2ZdsLlbIzzG/X4YWdp4HK4T
+dgxBRjGP8q9vrlvQ3qSMiQ0Vsu2GjwO/pZPbqIdfTvRM6Urg6iqQ4ecVxGV1cCep2eaSFglYB+D
1r8Id88OeM783InBuJeVOlqeH3JYAUbXV+MjVDOHgZPxEDR0rUnquQE1qGiFtlL7+rAxxKnDMCJR
u6acpDvIOXOxgZKKapSy65C496EGgDR+3U/O9A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7040)
PWxIP4yLixoX3mYt8VJcrywn/uNu/ZEfILHN4bRFAXW2sjFjhiBV1tPGrUmmgUZquiMhDI+WaWH9
IaAQ4Uj0/10ALK4r87jfFUpsdPNFV91CmssZajrj4KFHrGN3YAv3Ne+V0/z1JHk7LIwtPkP2o1wM
cXZWT5QRDZlmpR8uEMllQcLlfY1cBjzhRz0ApHwHWlcpA+P3LNcjnh0Z5+K81od8VaaIFUL5bzVa
4O4Z/sQ4JVTSmG94km6x2YMgB7WXfgwIXnJX4Z95fhhZXhQasxzgHy67JKgjHY5b/OqzGsblDUXu
y9ZyV3XfYO4j7Fdf10vlHz9lI0NMfj70o7+ID7yR/e3tw8//r8zqPRrDCuFDekaoxHl/boU6VXV2
1xWoNO2uab4evmydYxumQ1Hx2x/A/v3fOmlWpQe6QpPt3nSGyLqAp6i4vbeWDnCtVpvjNJPOGaaM
FkIs8Ij3V+krMtE98tJRtmuT2srwVNRCuf0wAmOMHuCJBDdr4y4JCXz4a/drfA1fv4+rO7AqVabI
jqMp0yDT8TxHi5IErbadZ2zncGdJ9H1UaLKZqgzicedpoarlqpFpeQvT/7Z7hfBRLxaGJ++qPEDV
mWPK3BkmfUX5EG6+ytFXDLLrwLuKBfYptVk9C5s4IvHrpocW906MHlynYH9Qqae20DAKnWDGF2Z7
2Dpq53hNuj+yaC73XjPf00uKM2c34Msxw/RWZVA5zA1X7qG5IfWxwzoWX3sGmTTNkpX/dPNzm/Dv
WSrjD5FHGc+yq0uNwBuCLNCuaetJ9sY5PtwxT9m6tLQ4s4OUtxhD8aQzH6SK+o1GeFQmKngmsYBD
IrYEimUnRYh3SMtThSl6x+2HZarnpcO4zZY0R4dEP2Zhn8j8M+LUU4vY58qVrzY9vRHOkq6pIeNX
2A/h5jgBRf3ngNBIxVf0a3as6gO4JOTYEc7ms1bRpjJ4H1E1o54ZQUnGcxyavodBItco07iXxL8D
binWYzD83PRBH4bQJhZNKUDPYGeBxSGnyOjbqjZth2sQwgoc6K+Qkh8KUT7HKVVqAM+2DC0bW14l
MA3deBhXghMxreOC/V5GGDnFLBXU5P75YKtbdNVW5q1cwZQckEJhRSam0L9MRfuk3rVenp9+S61V
Gwl20vD295hRyy5y02flz+1BRjrC1MEl4eMGYnbDlNEjYIhUUTSoJeadLmgLs91Gm//3trVis4em
1dBtq3JMJSevn3Aptedp4N/va72m0kxSL3fWed0ZmiYH8MrfyoM+7i73Qv7rbMstj7AFgGnue9qI
g8QW2LHsAIy40v15PsVKdQyIAUrrjBbMwPC9XvtY4WRAXr+2KU4IeFHstC1Ms3WzLifeuUTP+SBu
jx9iD49K8t6svGE0htc2sTACnGsjxK6qtg1N9Kx9wXg1fPxnRMIZ6J+C8VPNvLGlVwfQjRqDhBTm
72/chIoxGAS4bCD7vpwBeRWiwsccbLXNEUtuCtHlreR913eOAGSB+sQzGstyoVwUzi3fhJI5/BBz
YXDxCDaoNpmQZ4ad2B+kcAbFSO7vxF5NwE1lBmqxNLEnm8dGNCEEyj32pFgG7gsZfxjDzw0dxQhk
2X8OJ1ifucelvQrSCKxOYiWT2GGBLKcS9PPJ/vUVv2P3ngwBXMeG7lBlNoD7/8q+QY/SCyVtpE1a
5dx1Jo5jbILQemEtEWd5E1OvotPwqhcKAxkKX9MicRfjBG8Cb9RmfFCofetL34M2LEUpb9HFqGPu
BiRmfvYxESvKeOjuR9spVQK80OU+Y0ksWgmxTjg9mZuWqmCNqO1JzJvWu4H6OhZFvsyKAbxB2wXr
Al+jnESZV3yIRj1kXcmT13tOHfHHs4IL8YxHnakmyDnPeox96SOUeT1h4ByIX7X2ci3+n1pVnbBI
G9XuCWf7boXxny+NwQ1KnS4YbnTOl3rIDR1L8/tQgquVaM4vSq2gpJ0SSogIJNHMYjwT10Rt+MPR
HNkHKzO3GwOuDijJu4BnnQ5zlcb6DuwdxHWngG+pmukLH8H8YgFNf7WVIU0zGtEpPD6OiRY7CZaS
xXEJ7t7TxaVnYPU/O+s7LnNV0Ik3Lk4A/f+9GAdXhsb9IMiqsP3QHVnMN5EOEx6Tw0bBjGf0lHSL
ROPPLQlMn7OhT4JafSn8ESnnBFemPx4htj7XT4XVdUYWfo18vKTLUfUvgMPGtIBNx7uA4CN3mWei
DOk5qjn8NMMBhwmQeLHsCarAVo+ANUTAELt7O8sWnwXpm1vwy9B9J6luqvKPWjWb6lZyOXj0qOk3
RnUEmEjX12w/7kbmtgO3Zyrx7B+85SB40g37M9R1yOuuxeLXVy5J6dXofn8D+1SUby0SIRSCdYsE
0CDhX3fiZXhcRpqui94nizvaOToZEmeMvSFtRWOw1KKmBhk8AnCSlyIU9xMke4S/9gtzLvMXUOio
VXnuXbvNl3nNRR0qLkvATvV2ICKDznk3fJHGnIFw13Y2T5wNsynY676cjkyQwq6RdiwJc6b4Ffgg
jM87TTX99l7ZOwT4S8dG/ZcZhA3rsSe7gIl3RWnhnNRTL2xzehl0YrH0MKDb33KyjVoUaiN+03vH
vzZHX1Nof7oBO+UiKydM2A0BseuLNoAN/C2Ys9Pmd2SLXolrObn1O6WwCGy2cba7v39V2N67Jv9h
UXvgb54YUn9sXniREele+d8E3ymV8sikidwwao52icqXvnQrvKGG1dUBBRTTUA9hjEmL5FCAvMSm
hQsm9HZ5jQZphqRO+zFujsc76UfjeuhiF4wE/DJc8rPhpf4+XKKr+nUiVmOC4uTGA1r1jBAzJrQt
a5B2cP9nQiQ5uRzsarZlEYLm2tlrKViRzbjyRF3EnrvxKGL4+egRshzg6+qb9If3bxIaBRrEVSuK
QDyQFM3jIR3dj/Cuwx6zx4DLl6P5+6MVo7vsfWQQptZmXufgsH83M9yU4S2jDH8tNhAGqyTcfCmp
XGIfTY73+NOv+/YnUasxElY0xIXv6/qgrnmvZ50vN2N8ByVBP5ef2AkZO80pW93BMj21guFupumA
gU+YNIBDsrDk23/vq/HiRYmWXfsNL6T8z3Xiak6WZKeg13t9djekxyuuieS4b4jGQwjetyJVx1gA
MmfRfxz7WZ3+L1+lRK5Oe6wDKnkNEDxLqNLz2CWqkFSrz/B4pcVtCT8y/GbdFFk15dfwvVp4uF4a
mFGHUiid1wrLjXS3y3ZEw74DchD+8mNi5dPBrKnzUo7evxNWUh+9q+9pHXwY97jjybalirlwu7Bt
OtzRlfp2wpr+/FrptgUk/gw1zQ5UCgHku50etFa4+9xI1PXA9NwfCs5ZmIWuDWyJ/JThsz8UX6rw
5Ryl/LIlHd4f9G8PzCzQes4oOaYfPBRd7IwYwr10OBVMEM/BO3nccw/g5dAo+nVXEHsE7wK+MM4d
5wmZHtfo9ORqGR5kEncUKrt4azPNqaQ5HC4c2kB2xcTMLCwU4nZ/C0/GgfYnAdxILSdMtlp5ZTqR
nww+/rvtPctSEs+XnvMZUH2tpRYiuVIv/XEdVBoCMmHbJC3Aaq8azdRTG+/yhchJo9yOGv6eBgsn
cyjlBNvLxloJwuiRM55NXaRCdZdnFc5/EpGeHYTxCx3cFoMlZYfcEVZWpwfDSiKcm2K4UaqU5OFy
szChsHgmlMiaXvOoblHIlum8Hm0EEqWzK499LLcO9qDjVCdqXbG1yqXKmZvXcUsu0d+ijXlTxOh+
PGmDR0qlixyfXnHHOMEURqnniEhbaXyeIZyt0e4O1hGpJ44rPWc16CWwQHQqCg03ROzRKykCWI5q
0OofvodSL2HXWxDgaywSHshIJ0XHqLz2Wpg+CTTt/WAZaYHjip3RXtoTmAGy+p+gOGIWabCssfsX
2EVnhm7vomomY1m+pl2AKwzrpIa2Yq4kyjWWJU7lofHuQjsL8tSFY0CjTAgJNkxtplUuLMGY/VKv
Ikdzgk8daM2cuzznAYdFc0B/J8pwKfoNO0y1TmMSMF/LoiCYKK+CTB2pyTal85Jwf3USytWqCq3S
qjGUmfn7iAi2ILdE4Zrc+wk/wjls5HWNomXimmf8saaeMIMTV7Zs8cjs1TywhxP5KhmZFlobEaFz
Q1mEDXcZEn509wNRdjbAkbesE05pUqk8AKWaXvy+v2pgvcsx8RRmlTeJoUROgaYRwEZ7kgIDE2ub
4lKq9O1s1qdKmf6ooVYizhNniGI0WQ5od64Z9eOd5ZNGya86Cclidef1xfPUkOESs6qXoQdnzkEQ
hgvKXcW8HiiSv3JwhhvtiEjzM26ueSCIzx4Yd3J3FUYcQUqux7ZY1wZPKRJQaQ/SwwOPRSoykQwW
5C17DiOIBu1XXq0uAEC4WsPN4JYCqm2Y73+eRpLzIWHMKRhPgfwJflzA9PUO6MUinbTaBLuy7xfB
h8ItL1+DcQq7JulYhc8wCkzcRZazouz3rC2Pu0WUG/R7RBzJ6ssHKC5BnCuY+FBGa8sYDh7EriPP
3tot0a7cDSg6ZsmS2sFk5X/8V6ZSImKtN9bE0mcKfVgYqkgq3hoO9VDSXFSRGYfWfT1M5bTn5Tdb
C3lc04sdrcl7qwa/zW6Mu3AWpZvJswbSDoiV1G7mhWm4ZWOm2/M5QFUxpqOX/0niA3hF37jC7mnX
coVZW1L/u5TaCdjf8XJyV0zhWf7jaGMAJtFE9YQKZiD3w4GbUuRrJcQwoD7k654QiZ6/6QMNwXse
91GWYtynv1cgTc6zfTLIVqA3rPBRFR3bblceGTDGQGTVdQG9J7xc5w3trSxicQ01rTpxwXTjJBxF
e3skgHRSy94IshCMk1QCz3l94aCEz/oAP29wGVihA1g5Vbu2BYykWbCNcQvH6pUmvnJ1VAruxMQJ
zZGfrUhiZAlGHOu4mcqg7UbtNV+Z2jE59uy760bvm/U/saqJNTOhcYGd2Qy7YZ1PgSso0Yen8k3B
TWAXB01RJEwOiq5u1ywU3eJEqzDPpnvivtxZEl8USK+xK6LTsgUbDaL76cIrbyxz97McNcSGycSW
sNsNDzqKOw5c+aG5lRrFWMhyW/vg8Bb+YVFsq7padpM0eawht1pHgZyKmmHWC20Sck/FSqA7xZA7
iZseXtYGD+vbMrwdfm8zkrq3eWnbfqn/h2x0Aflu2fztf0t8EjtMp+L9UtmPTpLeZCX0FT9vjSwK
ljxxAdZ0HkGSROvz0ibqiPqXeZpC0pmRFyn51JEIpuu+g49dxwG1/V92VsGTunhQBU3miHlvcF77
g/OcGdkeKWAr3wIJfXUIrHw82tQAiq2VNrTZiYvTt6tPpI016KPwADsL6u0UEBK3T0Prtda1UscM
A6EZTZB2fWvpK7jMajHydDnnzKB67+3AvfvuHPkDyQYVH60IYWYjzXfZeSd401B1Xjl3/nbqymFd
dbRKMViJPxPCruWMaxfwr0URXt53wStoXyWsy1cqZ7Z6S2vehkpGyQg7no+AulooFxhZvJDNcexd
ym5CPk43dv3DtO0NKDlbJ6pJSvV299zqNeuDJ8n93eQ+LiZ4nDI5I8fXjBUEEWGgVp/1vcUorDyB
J643qKwP6xS3s66zzRJIHSme8CfYG4eX/ZNkkqGei/oy3GRrYHfnOauHG+kKQpZuM8tMJhE9q0ur
6Zydlp5YG8r/JDltY0O3q8dPYEyyVnxXdtmMz2sMvIym6cuGS7cG26wBATNW6fCSziPy3F0wqqbz
AVHLMJoax/PZnIPQK3TeVwjfrd5MIMP+NY7iZGxG6Qz243vgrV9p6aN+1FthIb7SIboyKy9k3c+1
cpVfQLItsTUDn/3HotSHgwGBCns5TBIAGhLNJqqXBAbqCelL3lzoBDQLM+Zbh8Gn/RyjKNpa5tun
5bEdfyJY04PvtdYoMJ8796ZbQ8IXAMhYeeiu4c8msjn0y8Io3fOnDXakHc9oda+lbKTVN0I/gV5s
tDMozHSsG6/y+gErKi3X0yOpuIQsqlL1oPpUx/4MY61tIWDyxmIPj973DD8RHeu5zIsmxWtihMnp
lg5GD3xp69CCkdmdaAmwNffcLdYr10hclbAOvjr/Q00suWABDcwU/U9JZBRGQVVLaLNh8vqcXUB/
ohU6tN8LR9hTEPc/AmDTbPwDb4210Nvi2UV34Rt3NWidOspQmpjepRuMGFD1iaBDVOxWvbAfW09n
P3U38W9p2te7nnDrPLUDtGSAIuxnKcpvYsH0J8Z+yd6CfjEry8cT1KO0an9b8r728eqZg9WzIpmX
y8U6l9nVyFm2nfHj0norsU+z/kpRcoHsi/u740jZTiIlG8fhx0sNfvG5a0n0mKSYfZwcUC+8SK2f
sV3maKZEFRWfkQ6rz0YOO4nouP8uUrv5IqkBSNVEJILEMFRD2ZY+dRnCOITXM0YSWsOHlb39QkCg
JwJWnnmEmY/CAbCDRJ5bu2kRDZQEe/3hfRE4bwK8u/ZBi988xRcFJURPlDNMlT5TkhkLMyip2zLH
g2qTPlxlLVMOTbPWlMvY9jT73nGtxPBOD55ZQnWh8awC1AlYUzqJPaMllRdY68WQAM/jE//PTcIe
S/ysE5tN8csiwdNKvS5iDiiMRl9ZnF7eWdHz02sWcct4l//kgzCrAxgayLNgDFp94Loh/nDwfTKF
qH6F7x6BHOKxn6ce67RtkW5wsJfo4nyfK9RDP3uYJKVynHuDJq16GNUn0SLg2IL2kgfRRtp7k3vt
nFJqh6W+djuCpkWa8BI3MTyctV7nVf087tVM8A1Lc09TvssJP0s9v4KR/IratLZ/kPpCX68cvXP5
vON5p2ulr6yiMvVL1rxpmuKeuiseR5Azl5g9kHeHdywt8zO4Bd9iF6V0zJ2UhXM5NZEOQGYiGb7y
SqeRJ1MYcoQeodEDXe+RAEq8tUzBFTweoss7q0pMd7mQqLwW32OvBPpIh6PkQsEL0aKWHQR97BUA
GrRlb5pNb24xjM6/BkcW2oS/DB56wLQ6T8aZum5nitdBFUsRtPYPcS8O/mqgiw5NCLzs5+br9x8i
iW2p20TZDh4i+p0lnXFJJyqg7uyryxdw+L63WMPoYmsarOcEg1pA/JUicAAAO9AOD9hIGMDyhmTe
ClOfL6McCns8cyrBGPFC3gwY1xQGy8vtKk7nwjFqtoN74Khnzo0WNf2v+sQz8eXeDA+4ZZ5EWLPJ
JuTiqRZKSHhpjSNMXI5N7rWOFQsZta4RAyv+KYeGeEfz6whS2QpwMLOeH0b0LMpdurWPGCspFwYu
VHuMfid/ggoZc5tOWgMETsYP1y8wqbNWBNisK+QlgEnHqzkdbiclNwe5P0B4UJthgrwLahBRyh4o
yrTgo5N84xwH/d1Q72ZPpSxjQVT/YYHnlxdX628xwfsP3Lc85MT6wweFBpInxsgrtZCJkLP6q+08
O5pL5LbVzOS5XfsTSVuTaXPL3c/beugZIcLhbD+XsT8OeIOAmVrSOFzK14WZ8zUgmkJmyyrfcevz
PCCCoXfn4bBjn7oJd6HWyiovarmwSprGCwa3g35hZc9KUOryaKBDDAmuIxt+yanc/XU5zHfu4nIB
bNh3uWwP8b/aA2AM5VPODM+C+sQzKpMyV9wyNcRnqTceU8MkeQzFFGhipvlJeDn8f3nGMxhe7Q4R
n0QPqhOaSPDM9EMMDp+FU9LwMnnI2aZEQJzl9PrwgU+CjXF6GPOl2/KCFo+nFwfX8QVFidJOOmB1
WuYJqs02ghTWK9YkPL600J4ElHyrABk09tQP5YjSnv/mY+/KK43V3ULkDHBbQv5FbpX7jGIqEJQ5
l17ZJELvPxubqjfg/dar0nxGpC7oqTGz0ZKmuOXEX0igHEnlKDY+M4z260fTbK3ptXUPJUrQ7Hb1
/q5nC04LKBKWNrO5P19nr6Yy/nOswO48tDPG3x9iRQ8RkulDsdQ4xvAT0dyR9XKvBApfoiIhY4dY
knrq5pjFq3WAGdocSeurMMKdAJvhKOwDY70ro9mLdjiJ7CJYGeUJUCNVZacFTeR4BJCj0KmP8ZO6
BaquTnZXKhFz+XHk38f3o3kqAiitPyemd4exWUYiaZBV9Jz/DjlNePsqxJRcd9bQzug8lUusDdAh
PjpAmCvT9eiZvIiQt5Ald1swGn1WOAtRT+MwU8Tpq6BijFqVBpPuY+dJR0/Pgf4ENfBpNidj2wNR
NgDr3AW/lUEPOMesVv9l6GUhAa5m1tGtkmA3jOvm8kAkK2/hX3eyo5hGSj9/43K7pT8vq/a21Fn0
6sFqxz2ikT5WALlHB3YZXeKw//RJpyncX8hCBUfH82F9jXowHrwcRAmGXn33RmX/vTZW5PLJikC8
/x7O6e4lHakL1HA1Py2CSP9N8OQEI+hAKR5ecP54QAOAIVoD1QBY1oPdiNeSLtqfSawKvI6J1uxH
Plj23Y5uFlbiZSNxBA7q9z2ocmdMyPMF6zJX+kLjqCvs9dpJRUGG5WVpbEhK+9DQruLCuBTXiLOW
GebifL8wMRN6urt6Ds8KPnBBf2jCyKa+MwcldxKI2GJdioPyEUEB6MJkKpXgRqkJqn6FOqujhE7X
ez1TAAbI/kqUmwX1o/jOpmweZ1ajzJBptRYSSqjL1BrSAKbvShF2UWK/4WtCbmiQZpIcRUYb04eZ
FfqktZV+7kv97dqNGzXJMZIykqiFSeQrctRVWV82OZ9W5iNMRL/93neKMDL0FWwCOtxWP516CbQ0
T9wxcwI4Dda9j/wzMg2ri8ZZDS6LD47+NgMytW9rAk8FyNWsd+71SMYNW8xAvNj+xShhud90q7cj
w/8zBOv3XxH0SOM5frCjig3Gj+DMjCF53wNbyPoBFjIwJgc/mtiAZiVqysQ/srrTV9SzCjeROGsh
hprloZwmmpUKrQ8kglTyjjqXNrCvCLgfnO/oRdasQe+Nv40HufplFyoapQnEf+o/ND1/uYEVz1mA
rc+PPF6s82nAt7QKl3TZONHr70AgwWXp32gTCtCFc/OKy8XfmehlwwwlwIps7q3UgUsHy8p5LQh2
VwYK0TbWfOFZs8WjENF2zCj0TcdbURoQLrUNdF62qwv0NWP4eNzSE1KMbSqx/RUGyGd8lf7tM3sg
uyWxj+L+omPG8s5tQ2Sgy/Nmpmh7P95i9xZvtV9q4bRTzpt3R1ZdII8cM91IHwzeY6n3+FTR3S2y
g4P+yhpihmZqwV4k4JcfwiYZEzyGo5uVrjHbnGkaz1wBrqTUEvZWKXFZHxgfNsJyr1Vm00XkM/+z
ZC3LmAS1MXWogCbjggLh6QMAlLAbZ7CPp9Sj+Gd4jLLN5Hpb8zGwi4eGS/k/ly2Q5QDrXjdYqyeW
yuwQF6+Qi09Cga34ofjkq8E/63zN2xYjByDxMhc6rZDCxPct1mV3m6VjR0wQmszZCLHG23KdNE2d
UP8hXnV5gLcnhAQ55nVJpxHo/XmxmYSDB2eJ850=
`pragma protect end_protected
