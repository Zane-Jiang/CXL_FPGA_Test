`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
F7fu+/LXTQmGy3nrJaZFgTj8dRcckBPVPCoeMd03TPqzzh+i7M/zOSNRjU3lYhHi
iXIkmSW06Un8vfj1ItqBMQYwJsbDgsi7qu9VZKcrzEc6Nw6LnBX18puKtpW1OUFi
azWcp4remXUype32vL4gt+bk5tOh84uKNta7FFGsVtk=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10416), data_block
Fia5jEIgq9XGo2rD9ruOBHkcsHHS8XR8wescTsftlb9rzqIgCAE5ji8/TT0c6kfm
EucirR0GLxqqg9lbo0hgwFePeqdaixmcIEluByKOgNhjzm2gm9UH6FETTJxkf9rW
GeaUZtjWYtuoWJEkufRxUOF5jq84h6FSNLoS1V2kyxl6K69uHWNA2T2IL9ekvkkx
gYWm1gDdqOZYh345fWEmsHHkQWeBtAxSoXERtTV5hSlPmrNCqYpCx62h0Ula6YRA
3pkdEfAOTL8oXLnG3DFlCy7lXdGABeVKWUpsmhzPzS0ZiU++pgpsmYCEN/OWbl0P
u8+pouZSHJLkznZ811XOpUD/s3HU4ny4XA5kKswOx8tcdZL7/hoUltmPUsFo6wQ3
dbYjTmAIiwvfTq+Z/W0c7bYrb/5WypAVhzNCqVLVH1bRakn/lq8/tDbhPi5LpUm1
hg1zDPEz5qRXvJ/xY8CLu4UiXuB7p1WrPeHfIpOwlhALLnnrUEjOPw69sTR9bBth
ZgKc4AxI3TzTk7gnkE0Cm6p/ZqYw8Tto/s2eL8NQVGXYN9HIP1Tg3CNk8aDNkyIF
moH3zUb/hJfmnpgF1F2ogTFNuyfdKn7kQXpop8YASaBLPW3jLH6I64WuyqqlRgfE
L8ljfTy2II46nmHM7tElcDHVhVJtNrvsLu7i16L5gztvk/nazvo9qPtWilol8Dz5
X1fT3DzWO5sBCit4azRceF+TqfDrgiQ2pdcoFojdQdhvofbdJLJVXwUegpicHjM5
i0jiAzuQpfxjfsehuPRxNLsAkpio8F9sx6iU5abHSUuCYRtog+5y9HN0+Zo4f+gQ
DX1mSABOA6EmAJtOIdFKSHZ+ierQ5Oqxn20c+TCEXmvGM8z3OVjlfHGIgaZ3t3TF
CtDU/GUoRgSwdbDHY0o/0tsV6buoJBErmeqSPJbVB57HgQQN5DSeUeYE9E3P18+7
u2YUBCOY7XCNZnby3c5NEA1EqbxlGikzAfG+TKno7gL45ghOeM0XQof8X45nBmlD
uyoRLxFmqHXy5+iuPgycT32D7nBA9zuh9twBv0GMDJ7tnzkq43i/3OS7c1G3DPTS
UZhWp03fbN37qQVzxRG5eOMpivxw/eIfyIdruqKBZkI17JKOk/id5E7JMqbS8oDT
3VMFDTobCoa56+YoCnjDALzKBbZLVGUNP1QBVvCp2yOqiIkDIXAvnQ2rpYRvUxg2
hVSzF3WRkybzpz8466hGF3lUbZjluu5DPN0Xo6Ir2bSFByUoEp8UkCagnFghjzKH
+DHZ2Z8jHUurG3n+HdoWjVSaD42lz9GAwsTmCKBstk5Wt4izzt9e578PUQtSIafV
uXcLKoeSoyg7t0bdA2zOPQTHcGVt896a4pPbLc/MRPxnvz6VeeFi7J9JpTv+OFm+
1Rl1/DybCPgfhPWhaH1oY9a6XWRXWmMl4kibufnv4cxM4odlqjbEMpKoKUuUZY0q
6Yj7BfEj3WCzFAzsxy0+YjMq8C+yyr3TCFpyGOpaugIrXEZ0llv05oyGCYtS+C56
N/CkRSVbLpLkPnfenapfirjw8FCDOp8DN2fxEjNKmPvoUtv1kiLOIelKCNyR6g19
1/WrTKpmDwDdRmY1OmcApr2AV+x0I5/HVGY0LS+5RURZUZBG8mGJ95tvNt/ZJcKR
kfdk6v75RsiCaosZ3pKBxDaDrJScpO7YRLy1PzTFF/yijqVjv39x/XIfWRtzwyJS
upZrUlj/WSJXmmWjpm1Ox9vfKHIIkUZwvooB2KuamGoMCKzcuEuSSoPeZg3uLeUD
5zZQWwU2bFKW9DB2eW3x61N1rBOM+jkRpCNaIPHu6KdbNrO3Muy6Tcfv4fqchfLm
ewCbrIUD0AptAiC8kzTFnXwHkemAqYYjSedZLVWaqBu/EdHU021+zqzwcU+sakWX
ZrALzKdr/+glbOXwfYSPszsKC2nejhp6Eatf7bcdPUjayZyPrfNWhZgLe+WOaUjg
jyhXXmdkvRjxZ4o8cYVKwW57czx4cQvYbVtPaUIiWHaxO9CilhI0PaPJK3cVUvu9
nK0h7pguYZIvzlga5oFefOzN1Zah1lrSuRmTKgBzMlPzaIog9tPKftndVIbcd9Qb
ystusjE71GmUsBPQh5e9s3Rnrn+RVcjmt5/l8ke1KxhuV/MJQM/XDq/qKzVNzu1e
kIdPIEK7lTs3vL/7H5NdfutKVONIsup6ba4WX6ZwuSdsTlFxW2mMBZBAiFu+n5yS
g885OqyXTEAtnMqG2gbyQXfWWJ8qDZ8ihaOrVsd/HJwYZKSOemYkoMWiZ+hGkd5e
wo93fKG/x7L+237Azpo8ZjM33AjbW3J9u8NLs5fSx6JatbYRoAAc9nCWMgifyKIO
LvlrVM6sfBVgewvEYmlaKf1OLXhIYai/fU1s3JSpMT2fIWHO1+1lWX8YdRGg01pt
ZLrR0Ov6NbMkPwKtnAtN6H+BYyVDw6qbDyrfTNWider8EC5RiRtYU69zNXTAJv2H
lPmFlJEUjxRTsOMVMtXX7c0CdX/0WL+a9FVfAoDQsIEUi6WhTIdSgIEVHLaCLOXe
SnEj025hKRXtFBW7SH8GQPo2hblIJ06IvU0njrt5mrLhbRzf9Gwp4xxO3K6wA0qW
DMRL5qp3Wn/Y6ijnlTu9W84yK+0IYLqPe3tNIaBohEbXnrmkptjLcF/KTCNVvg6c
WirD/P1iZmN/RNu6En776xwrAbZCVa8SpPUGdaQJkZ8nDZp4TE5FZ9mEZlO2rPX/
41W8OF2Fy5tptt1lFvbLpDP+gJx2muiyIuZBrTW6Fz7U+FlrgIaclE5Ku7Y8VCJ/
V/IlOT86cr9WJUUDHWtkSbnqUcR6EnLJt3rBAQQ4dqkx1Y/+I+NeZDLCcNuRF2TD
y3OWhyz1vumOmCILTyfPW7f4SvsUIIwnqmFZj46reZWICDLFoTs67DYUIzfwqcd5
z50sta5AoCyAU3mZOF1Gvwq/Ix8zEbpf6vSxEwcm841a5RSgdUXrilVHGRSJgklD
mrfN6yW6ZyJNZGM4tprdzEmB8ohmgCJq2oR1+uKUO55+TlOuD9jLXzIcty49T3cj
tRbqPq/9GJO3tuNt7AiuoSwY7w40sFsfzxC+ojYrxmqVXaXgr1QdXQCHC3zTvXP5
0iISa+Ra/fiav2r3AeDG586LUhGOcSxC34f0UoMYr/TU5sIBg8+5tit9/CYw6hL2
sTRkO1c6WhIjjjVjeKnFDE47Dtlj9NYKQk0Z1GiXuqGmuKVZWff0vp947wMNaY/a
8R8fTvnlfi3BuKTYErXggv+rJ17DeQnevmdqnCQNQNLsxHdKJbtcq1TENC32FmGK
liitIICSr5o/99+Be6+7ksLCKQRP5x9H5pkEgh6iImtsMd3s/6yqpkfNDqsT045r
/jM6aVjPe6JfgXeIO8FxFwuhoZHDfylYMyOgg8PL8CyRcFlCi5dIqCWF2m70At2+
OskTiqHTNbD+lUI33iLypKTyqPKARezap5YJ5GvisJnRMUX7S2Ea7/BRMGWsz8qw
f6IRZV2vVfH6d/39chtOhFDafZVPuxRNbq4+07QUeuwPdcifSw4nfI7dYNHKW4R2
MP/l+ts6GKxuhMTS7sj9tTWEHtvdohGkaBZIGYwdjQR+U2P6+Tds0UKb+xwyZ4YQ
NxZdpiDL3OKa+dQNJef2INeUDd6aNLreyRUtUkiaTPgPxkbrMJEH1wJV8pnBihx8
C/LauNXwjkutk58HgVJQum6P2HDOQUiuCz7mj4GZvRNYZ+WnZA4LR/3dZhHYVYPm
N42ltN+YjngEIBRUHQgUCHpNJ0Y3ccqK/OUR3hM0Twbk0xJGkMsz6BRIJt3ZLv08
G6vcWGZ9qAFfQG8Jn8YkDZrlm1YkDjZq/G1M4mQpNVsYPYe2HU06zvW91HEgXmQ5
yj8ASKZsinUkvz7coeA1wyFtJ5VKwMId8bQMU56XbfoznVoEX0IzyJ736E5d36ui
cx+DpurVPUN4rOOMiklkZnxlTYobEL6IJV0WXbHEL006Y/ZYkHdqQoehMo2RUA8E
jLP3CS1Pif8BkLUkeF5cR1xpkOW3FNHCUabtW/tsu4GXO2PnXfnO9W60nN6pJwDX
Hjdnzo7qto0UzFexFO6VUKtF0koNBbK4xWWhr1B2exM7KBHpw8X59M2wqjadeuCL
o+FVVPlePemDZxiiAFhuwtp5MUriM6CpZixhvHAEU1ph0v7Eo5Iyh67O+K+QYONo
iEQLRA2pS3W4t1QxqYFpP9mwILEAzpbXWHvTxbBCbV2y93FC1AkucIXb/2eYmVkW
aJSlyHcQObX+LAOUbC17BXTG6FXG/3174+aJ4wNoxemmBFsxT3Snsu4EeNWC1RHI
Qurc6s/NihxfAk3ezrTKJnv6iu0IVKBqGFcw61/IAfE7kg1fW80qMkxo0fhwUvv7
knV6t3z0m5xa6yWRVph6Pu0YrJ8VR2W1p3OCJ3vHKpmZI+nECd4Dg99Owhx0ZweW
XyXT+g7ajSxf81ieMAnEvRY33gHV493pyV++UDCu0kK3znsmSGtN1xmoCF0GWxqK
h28H/r82XjWmmRe9gSMgbJaqr9uO5/p+QdPdZPfyceEPGleBeXBySRM9+hkyLpSC
FCodTRNu2YRzbtowyFX0g2c/GEU+A1B9Lz6cqaPimZYPpuIGrIU2v9kjdvaddkr1
UQUrO4b4S7OrAF+C6gaqUfIbB5+mM1U2Ubh8E5K3I7/c86yFbqayyfV4oVrPWlqk
3zU0gskYkgFCDtEUT1/mOo0TaI3/AI1hO2uumXrYxVG8ZLgE/4lA044heuHZwA2d
8OjWkaLocIBE9XJuo0Na+fVrGKV+nj5Ttv4ppieRE1S6hk0NkB2Akldlm5OJWPRn
OLFhfr/Qp7/JWJm42USMJ2x7d/J7lKyPql/fJ5AQtfURPqU5oL4LasLm2mvGRIHD
iz3O5+lk8tEnOTlfy+TUWpRaKvy+aUQjOJEzTqoBWXdD+z8bjQ+UMCinNyiOIsPy
tyxLE3lckVlwV34GlGxioFYnJdfO0aBnZVU5lJNgiUoAfCsgRGS+ScWkNx1UWGz+
yOQ8fH2vgYmgH0J2D5DWlJHuSYgXMZhOW9XMX8a3+F++P6aO3mXbOif7wqrWScIk
SJKhl96vX+9BV8X9VPTL/dJ08jBz21oO88ui3zEXap7uK7ekcIZkJ4luMWOUhJB5
qn5m2XpNFx+A/Kck/BrWGRrYEB03T0bcTAHBBK7KM0e4Dj6B4hHhhvp5B6GfB5ES
9VnCNwhLmQRkTyiiJwIJTFDhPPLrB3xYKMujHbm4GJKYxaX3upjqmiPuBtwW3gve
2ZK03qEMVKj2ABIn3ohLBKU//EWVY16wPbXTAoSKE7vB7C6DpFgqgL7w+PJbzRC0
P22n8CNiPQz3Z9i8a2q/IwBO14zCLlPvuLUWQyA2N/PhfmYJoEeg2j8HHmCkxZiJ
Dm2kLDmvvg20kZraEauSJrbRizDeBW+sTbNSpWfye7OxQ/AYVzulsR2SN4GFs2o2
1gfB0aEjXm0xojiENFcNEOgbEQbfPSvKaX68YBDHRLuXGbzTJmvjVVtXzYzrmhEm
Mk5Om/NQQSEvUPZyp/g5ved4X9nSbRM+pNkCQYJCc/FQe7mHj3bGGUjOwBo0Wguk
Y8g6Ti1gIQTbCbmc5f4RASCv4bXwk8jDBlw2iok73rKdAU0rmCaLFeMCexkFQ5qk
5v7D9HTXZbAwq3YBfigM0wCrQrz4+6VsSo5Kn7CL+rqHIVj8nbATJZ6mvA5Z8yWw
oTwT3UYS6IVJIJ266XNKDAIRMg0ZEdSljgErxkw3Ed/S0T2Avl9wuFYGx6k4Z0Lf
5V5N//cSfAAryvEiolnHak5x9bPfBANTdJSHEZiP0nYOWmFz9F39mnFu5DvjUSFx
fLDHVx3XDhrmXsmpW+HdPy5iRc5Zom/vWvDXZ3ql6cT6G8HMdaDR7AayOljl74Z7
EYJhi1Cp368DGQrDL90EMJ+S/B4bt1mogWiWCZu4GAh/Y/TCoPeGnWt0MkSCs86c
tXNZ77hKI3SJLYBvjXWkt4fB9TuupGPNXgNAhqP95pKeg0zDIwspY/yz/XUmffam
GkQCQ1CCdNmeFrXL35BErlH/FBLlHS4Alq5q+W1d6a1d9OC5FKcwy7gOy3/CLnut
SfqAJns5QZeqdo9sobQi9Cl0QtcFy8Sab3S+VglyuSo97ukKH2u1KU0P83+3gcjR
XQaeHkz8YVi3P+CteV3WI9mQh5BeIxz0XuunhVbdRXAa9t1YMbuXKetIRsR5yueB
aX/33yIe1KUf6+lpR0rlmmU6Q+O4TxVbYvgM/QPEUn1+PufoYnlrLIKUJHVFASn+
HCOYYhDQ1azFuvoUzOWib1p3zf6L560g+r4GaFcw2m1npPzM13S11E6pfeG1wZM3
trk+EU8a1+2T3yxWv3jIFowcEcNsBeA92SgGS6anYyvjhlfhZ3tEPXIFIvk0waaa
udhLqITmDawom+Wndhfx43Pas6oK3l8P3K29DnrRWwomS3qIoJ8fahWRGmjBoVY5
6W6pfSzXXv1if4GsWrGsQdEaKRT8Vos4c0zvWFw3F5VzjlZiw21QBNuIiUoUFrMO
75HCRRc/wN+ZoAJysZe+tz2mlnL4yQ8DUZs/Hhd2QyNpdZUiBXnYC/7rveOmgeIX
o5JaiP+KxAuw77A8d8aql022BN/XYsg0YJWwr6ubqKRElKCdihPXhoFLpY/K8w2K
A3i0+96kInrFQJFeRXsRa6viu8lSmdS4uWqshnfA/kxe4P+UGIjWxki7BnDnk0HM
9P1a0iVMxVXJMfPzaqn/iKOjuShrImLb5i1NZVivD3LC8CEUkpii+lSve1hapYc8
z0ucVaarR22jnmGH7GVZlWfrr0Ux5swf64iDGX7sk/pQvNlKaTME6jSkILvqLcFr
dYp9kD1xupHFUFy0OraSx/ZQUmIDWTurIZPyvuMHvtmx7PCRZ5TZYQRanSYlJ8ll
GXGYdPl+AnbjnuffRI/T2wCDUHPPrsw/bJFIOykz2hWSEwTpa8AybUcfAVodzglT
vYyrwHA4ip3kycqH1J2q6VXiA//Ygn8O3K2+Wt0Pa+xq5mlSv6K4LfCR7/pczPRQ
LfNLGIoLvhYSxBmojCGYTxNu+mi4odesZ8BSFWKxTOJ/mwKOjg/yjx178C6z1aAX
vUYkKT7D71jgLn+Nyyev9e1DzYUUE1kMRdh4ijxFXjpuZdt9GmElKD/EdhHQUkKK
H/NVJWJAiiUFblVrlBfuqRoIRODYwUAMJEifl/T50nBka46Hqx9UbI/FixjRVLNT
yiukgb9es9pD0fSt3Bb5nR9HquQveuAY9oSloEfmEBaHDtpXYij+lr6PqpQRzEG6
1PU9rJ0MrrpUQqOBkQHkm483ERCBHcHottfGJUqPA832Q9sMBcSG0Ee70bQS6qso
2YKcMKI+I36I9I//eUuK+V+JCq7UF2/8F5WkH6GnseIVK8e5xsnlE8glDyP0dp8u
AFWMAsj5xUODyz8mZ6oxVK3IpMlsEyCS79dYTBbMnTXnyIzIOlExSlzFCcAv5H8b
4iNfg+7iRNU83secIqeXzmEMeENu/+btvHk2dsn87eAgtHejZr2NPIKfl0X2HfTA
Jw3lfpp0jPrn58cPfPRrxTHGEclEmHV26UH7vQF5JnSUJWXuSm1/WlTvlHD0ywqv
RoZ5nBW4AWG5XGDDOI0mTjrmDHkIWMZ9I41XbH6kTwi7Bm2gEXzXY52j4k3nlQrH
wvglFM3/ai4274AdoQIBtkJzctCF66zKeiPzuPHwZHUNk9irxS7AaPBGb52kPnKL
ttm3QY/PdqbmmZQLC6tNiwbTMyHkfYW7CVjUW8ZEcBgDRePKGNvjFGL3isuXbaJA
NTxb49zyQWCsIDgSh3KgDcAD1RXOnxrok1vSqvKNzeO5nsZ+k6KoWPw4CdT7xV5y
RGmTethu/dwtA7VhH3uORw0dGDUjPouCpCSTBxV8BoQc7GRSwsDP0+z7GT9IEb2R
py/BAeIdbGgTEIDnJj0npC7iW+u1xOz4/anS0n1BZ0zNP4tYYn4QRzcpuA1sJEff
WNCwE5ebqFU4bXGzIn0OdD5NuWAmQ1X4PHXkrXMXuRc1v5HCR1Wts/B7VQnI1bc+
AUG5zTvPIVdHK6tKw+YUWOIcLZ70aEENAilhYmBk0dK6XIlZum/ElnAO9DD0r44s
YK653uUkvOfOzn7ZsesLEIvVHQW0GxYF6NnwRmWTdDPyUxy/InavXzDRI24u6EwA
7NihJY95yrxu0WVsnR22xzfaz+trTpoI4VW8z/WAJpiF/B2eajUteSrAmM35Ysos
AkteM/Y0k7Gxnor8UTz6u8zsp4nI/sSVIFHHl+dTruaDko0EZWeuC7M+iF4nHSH8
VjIuHb31LukrxQw9m2DXNNUqCqxwHIjWkJCuBrDIchm8iviseqDlSRONOpfCSwY+
EpkqqCDTd+evH3gCCgfrz+JBhrLA/G6g9UmAzkfep37hoc9ZUfKnk6a7kS/OfiZF
GAyJgGcNsjyLUjEpn0mts/mO6bh9St/J2xC2ni7Qt/DwzCKDJFvDnv66wTHx4koz
GhGjuFlkxrM2TUZhKjTVUhiesf8i3ivfzmZOz4J7ySovDfcng63/L52cS7O3fcHB
DcoNP7wbFUFxg6zdFrx8U3OuMxxm+pZ1pZuj1fFJqajjxE3f0ZmggZiz0SGnCFJ0
6a5eLySO/Tq0MfnYyBSr2MtEKE36esSEo9gcYDVYz12AmMipuYSqmNas5NLxGAll
djeOELqM3nhWDMXsDwYCneGpt9SCtYP+aYdcoizI9eEzOKAqmpMuKssXKVdIMbI3
XfsnZP8tbvvbgrXQtzI4anm/clEyAk3G2LhGqvH/gjL/21FMDfhB4lo7V57EWpFi
W4DzqwHsRmxwx1IHMJgmIp6PWK9E74NHByxKPRil4CuGkSe64OR1GLxHOWj7rbtp
7AiaNVIqm8Bq1uJQd0ONUJYgcQOMhGyDKs6XvmBg/k7kUd3j8b4tkcRYSH57C95h
VntPO0jMUv8hH9UYU1O4/dlR9LChr2SNYFcu6CYaXCyY2g58RsqXamXGt2AGjQrk
Xh74uGzVFU8+XUqy+4L4kNQz3sWaukAi/+weQqHbihWiPallgNEB4LGExn+L0f2K
x7pvsCYEallbdTdr5O5GIYY2OgkWTEPxBBTWi2DV2WQEUQK59psiUZlVXF1oT+z4
3YKeAgq5lJqTYmtuAPnJgpTRxphhQdgaQ3pLQ/6irlgXuJFrMMtWv5uwREaWPSDK
fh0VkkZoJDTW0aMawdAgPnLa+6lhT+Zou2mPjf775jLCDQvoKFQMCqRAYtvzdf1r
73QkXrAqI0qd+UqpNX+IbE5y4HwMlaHoTQh1D46S/J9z+aPLPRqjnmOlSSWLGM4b
txaIFYtJvrtZPVpq1mwmMkOglltv2892lxPA68HgF37B14uXSm10giwm7drK6xOz
ISOFFqAWBAVJDOXD3Vzmr8esVcLqHMjJHGCI7mqIz//y5QWLpkwdTT3nNGVjKHRK
vGYWyrLHxHEFtZS7J3/wEhli6DDoUM3v9izGJJnWhZSSP3rqc1e2TZL4k/OPsc8U
kuwzGvph8S1M+PVTvrFOZoU3ygFmm2+JVLuzy7yyyAUv9KxpHF8c2queXA3BhyZc
BPoeon39J+IYGluko2c8a+/KhJXKe3JQ/snBoX27SRubvtxTwMe7h/fr+B0eCVdS
0fiBV4oMQvbx+pGM+voFUoDAnHVRX6P2E0Ig0dsjfq78CB5AwMYhkOqc6KqZmi0n
2BUeaK2uTz1MkKLwQotbpdz+6fMQ3V161hSQD01EVGmGbRmtBzu/OCfBFlsOil/u
StabNzgog/IinhRvPK5LxoC/+5gZpP9Z+hKtMDXKEB4+OOyAt65kEOzmMQ667v65
nHpBOq5auePHZxGL25cEkvtYxW6IBqrbpdgSJiE8aIEdPqELP4PXlBR+DIZLQjK3
gipAeyHPtHZz0LZ/4xiq6VV+MMzdBHilqhjaE9IFmLmEHy/TPPitpoo5coy9PFuW
RrzA14zpcvPMLxI3dDvn7qCAyQ5qgRao+DoQJKLgl7lnIUUPOwAO+nDD/SakJrno
/GoRf1PWe6ULff07USnsRRoz7WEL3G4EDyXmHd03DeP6umplhjEJ4r4HRdKkuYsr
UZIdP3kQdfLOqMQWquSgRdPqkYDrF/gHRji6tCgnAjckrdL57dvQD+eG2WyrOJWc
WTJyJYhL1sYSuTFSiMpuzRkj3rm63kTaTBCTK4LAXwDMqiX+T0faIAJDP3o3+URV
EA1pK/MKz8Sd0g7NNLuERTZSzAXgq3jSpHu4sXXq+e5b5wdfovINQ4D7uvfj5bUU
JWzkzYvS+XU+Kf3r5L7iXu2RQUu0GmIjl2VSvkPgzKRQUN1wp/dFNrgFOyLsLbOt
nVMYFULmOA6K9gRc327jmHSmOKBDtPhexN5Sh+xdNls2FRn/2GcFwkiirnTLaj4j
Utb7f37mPZbWT5DISwmvdziPvx9nb1/iApy30QD//UKjPDwsGi94GcgjsCCQ20M3
Hf+docX5UPHdpd9rA6ktFpkUZtLRp5ycNUX5ww+OtAVFxbM/ijBh/EWy820OomMw
Ni8zyioNzJJysZUkbFCrQJ2OsBFjbqv6cHm3iPVHDq+iG6qwOcq66SD9ImFnedev
1JoIHTQQiMFgW4EFx7OIkLbGL1lEs+VGeYRSt9n3ijdNLXQkhj/GS8Eonr3opqK8
t0Xcns7ghKyzSpjXHdseOs2Yopm8gUeuJ5dWCy27aEAdRkgg5mkCRkiWnk4O0zcT
FPWOB1V7ERRVKvuI8/Wlecfhm4uMLgYUelOnVS1W330e9yRoGNRcTwnKXAoVt8za
M121wu179hDevmHH+ZiWuoXSSXefZvFzfaXr5hFdAAyP/cuE81J99rx+xAA/uESJ
9+e5+xfZ0tURWUQTc57pPX3NUApeT6x1jwn0wlYG+a1eUJTCWkx1qlx+AJWAu4pd
6PQZsY+Zh9sSs9G90Scv5gfawIlCk7AF+8N9x+6NlM28hU0dqISMv2j73GP/IEbO
VrsvDRcTeRUWCChsPNNtHBP+OiMAOshOarhmfOWwQrywjZZ9efIoI1EjtsE2PdqO
xqmJkqyvzogdLch/zd14NK7OI+RM3ijwtxigYGylt9n7EinW5X8QoL/bXVqA287F
ThgbHu5AK8i+PuDemwFnshy5UukXYH1sWUIHFkm9UaUhs65xplOlSziv/zntwpDV
ziknASULRI0a6AJ47E9CFmpX0byJYEwtbKjOIVwY728HMY+5HHvTFZoGq4euTXGr
hFHDytjH2EHVofcSKyKW3dC+WF/CV8DILEIEQ1pDkwTJYsditd1Axx2Qq/2LqDvE
J9rv9CWH9b/wUgf/4RY4A8Kg7iqldmCio67gP1eHT0u79+5/Kj8Avbyft7Z/uWDg
ONPmKehOfPEeH5uMqlbpiatstIhFPRZcSrLK4XKWgT7IjiNV1BQCCjooFM83bvmW
0mj43O1AvEovrRSOhLFq4ehoV3IO9ZlFr3aq18TzI0TJI0DPK5E1vA0msFs8A3a0
/VKo2SA1U2DM7Ipv761Nx/wde8kco0Uy/YodMoj5XNIMLPrsIACLZvDA78DL1JF2
O1GeE+kAvOdvo4hxzwvQqkZT/aotoMyRvbl20A24bmf/dcCfugg0+4+G/8TePWzS
rXRvA+MxfWvL/wJIMN8j0ji/jWs/njiTHEXteMahxxG4XFsfAy1MWpREXTK3Yeof
zv6+jVlw8td6uZni9r7tDWGxaM6zuiGFH3ZRNgJpR36S7dEIIoi8RS9oqei0wYOH
ejXmAzRTr6gGe/j7Xt0eeAULnKt1FHbjOe1B5YngvEsCGt67FqFgK+tqbI437sT2
ocj2qHHSYxeCpV/3QQ5v3aMGpTLbj4bnUnQk4lbu13iAgYUj9d7gAo1bj1om94RA
3h+qXVWjUI1TiFJCRtac3rhG/2/olPA/2uMXOQPFXTuRHHt2tx7+ZCa22At5eUCb
cMvfXnDNA8GiR+FC1PIMyif5y1UJyRWsHwCpMErTaxTIRYZxa0Gjlj6ET8c7dOHu
ekt7PAtmf4o8xCSLQC4O+NccS1pvgJKCFQZ/BrfpZ/9PJaQT8awqIV1RlyaWGcfI
QX7tCDqusFQuTnlNnVREpCywFeLnMsESzQj+bG22mUXfOdQLBpy48w+KFtrlVuEq
r6yKrMDHrxesWshEAKcNk2h3ucLUY5k5usvCUoTF6lJBDyPvuPH5N7VocX7IQreo
2mpheMI7PFeV52jbDckmqiKU+yTF6FSR1jy4NcY0VtZNcq5DniPScGm5PRpo1IjS
jXlnsS1akMsKJoiqneYilTQ2g9ZRJtqVHXJjvS+r+Xp7Ol2HiNT+5T92E6eQEDn4
Q9vU0L9uUnPz3h8HktblEXEdNORS3/FceMAv/dqMElv16HWxjF67o0nZNjaKCGwz
DeWPgeRhvTWVIU3soGXgs3GP2r5x0IyK697s95344i/n6rYdTPRcsxVPP+ox0LEK
BScUKdlfIF4zqYm7Nxj1/4B7BwW4OTpDZ+hi/syGHtAJKrC+rliPAWaR4/je/2nx
76chgDBO1egTmZ9OlWmOOCh61dLlcDZPyfyvkmT8hEQk8sumQgPo79/+PGIFPPH9
/ClCnZW7Zw7zoIZk8sMfW1WXBocYC5sYHB+xOz6T0AgY6YvtJ9hLlOTsglSTptbr
KS5pLLsQcMwFZbj3HlXyePGUvowZ/v7Nc3wfZUuiYq49237MpHRKBt9lMd8vfFR6
PypoAm03WDU+HeEIsSEozkW1fZIsA87MOu/al+I96WvyoCdl9GvK3WpbTonX7G1L
RkfFScsRiMUuaMEMnbcFpOf8QK1wPGwmYqYt3e7FRz3qqPpOU0imp3zVEtxSwID6
hYuHwSCHqpDUzI76bIomEHxkCbh3RgHuOZ+nid84eEHAYPlg3GYjevis2ycM8up0
9JN67mIg3KK9z/YEQ3zJQLDPZWKj0T7HkMsnY7SIAKli53sLkGtYiyWSSBjBL76M
djlv1HmYykmUxEmEr5uZZgV6d72lRhDMIQi2aPXT/sGto6upQEMU7ka/GJluzoP8
FNpLG2bWMRdQHS9+orvxKKY2fDdW4UXY3PTjMeNZltJ137uJZhIdDtqRvTtqiLxe
oMYxWvP8VxZGzU+QCm2QrvsM3P3oBboj3L8YPEwajAQ1akvVtcKTVISVlLwSRYQK
qc/ws6gHQC5Pw6Mg0ZUAGzSOCyau1hV8Iqc7sUdCZLKho9ru3YrNa1Ku5rvFQP6/
B3DYoQ985b5WlZEQqahaBDNnha9RtlyMygl+GMHeptnxfHbg5O5pbPSctn91Asge
bk6BP8f6Ni52E3msDSUNmnWqh5mxU1Nt0l0WtSgoS1MRNEBfJqDwivzeBQ9dOAJL
9HO0X45//K8WDXdUvOt2drKL1a/j3hgm54fIJxnocm4DWL6TrqnsHzVSnLDxZfDy
rP8/KQHnjvL5Abb0EBOzp/CJmAnw2bMzQiL5r+icl56pesTv8+M43VMmktNsipI1
DuKWEjNAkRNvR4M3D/aYZzf4S5wSB9wIPFJCqM0yaDrTbnRmkBYIhmaO2CTvAxFV
os7SIN40+yyY+Om70ASKEV3hWm4+NM3UrhQzR6PONMOa5WYjkZLVOIVc1gM547tE
gkXL45MiYfaM/5DzrXoVjVllhl0YUWbZjKkk6glGKAdpzmk+21tmv+B7BfNQI5Dm
cq8Qt0a2ADKBDFCtc+1OzQuadKg0BpwZy2qthOI8s/QFyV8wSX9k86I5zqyn2tTz
2hCIMotvM/eigTLR/i1QHbzLk/vI8dkBvkV8sEtZO7AMX7LCYieRa9XUApdLq1bl
`pragma protect end_protected
