// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XwthqjMQkzIfqDB5+UT23H9WOrLFHz3F9wqW9Odth7KxtYf+1MONFAi0hjT5
PxFGOz53T78XxFEDN5Gnb56rf9qk8akOmCaDX1RRnK6xSWnhuTSUNNBYabwt
+/Vb9MAsU3P9IxX3kkZCrfhMwv0f4IlS19KO7d+daOeorPVMpKXrtFs72Gcj
HD9N4bdqq1EAYyffb5yCBjdNwPMhY8Gur6/qZOwT64lUEC+j5WPGm0p3ZxLe
MdmKwEIzWcTohfnpOki64m/vBkh7H1umVz8uYccyN6TByg3uELTqQ6m2kfEa
xOrOUH7GlJwvrHkgJ2waM17vTi6JZIVujvAwHbYOwA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IrUyNwrzz/rlABGLhgJZzSpxDPV4oJEnhPBsbfs8X1DDXvY9k4KXBUajAm9M
eXeXKXmUf4a4Wnic3RHdsrFj9CkNKSGOKMs0wiy5YlxewCQIifSRXOQaTWjv
AEuwksi7kPsb82uJJGuFAdYJQH4mZYdY/sRX71N8GDwn0d3BrddCC264Jwi+
9gyoCrckOtwwxJoVveviOOBs2x1u21Gb7gt9ud5sFRw5bctqlMB8iRkN21js
w5RYqjG1hC0T8wdoKff3qbNCboCddU4PTSjs7Bh3SiUHMPjO4aqx1+Ua+b89
YepLyT6vTFDxGoGIx0Jdgy3AOz3zHl5ls9Vc3BFQJQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FN4in4BenjReV+xA8QGWecUq+/p4gfwo1iAnrN9VNLvu+M9E6XYCKFBq4T9M
s10M35QvDIq/JTGpjaoiIjTJOmXuTEx/GyGu4TzG08b8KaW+61asnmREj5n1
d4W0NpdQa4iMbCPTI0AYowHLkKF96TqNJ7eWvKZD3DbYLPKVnNiUEaVdPdPg
oUFxDT9BKhS8zl0nk5Z4fqk5ACqoyuYzQAIb+2niEXZCalDMipYSpFjq5Bs7
urs6UF+pKFlODrIwvGnaEbfF/WsRaOm+kapiSWt6pVEdgXHMJ4jWBK+O6OTk
NEhlU2Nna5tuVMcgj4HcqLLsVKq/QdVxuOrdKsZMdg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y0/LN2mcEm9Xc/XnM2Wp/ecaBUZ4Z6Q4nfA/CadH3GkzJzeZTFzHzNIEBYWu
lKlWm3NJyZnPMrFAOOzkrwUuzdWexDNSuDd4tpLeIAtb1WsgrPm0s+ZygGyX
ammCFDL4rX+4kPcNCVUZwN4tNzKIRgVpoX4uj5WYI/1zbgTSdRg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sH/Uh20b5HJglx9q2CeU7JYRD2X+PFb5VCOiVws7XqFEYZ9hzU/KaFvtBpBE
YsMhV/ijUol3SNGTgAdqHPA3YzbJsgYZLTyCmmPO78DL+SeBix9Lt+NXfohE
aOSNzphj12B9kdtNnxq3dt/gQ6nbcCVgwfY1AX6hAxkbrnfnoGVe4Ttxw+mc
bd0pcAnHwLPmGhncRqLmuElrH3gi5d2lEop4YczOKn4letLRErlaLZoXUpLn
g8xnO1UEIjS4T9yZqtrW6XXHGn9XbIZ6eioGQWv8Yew+33QN1hBHp+Syqc+H
q8SHR+m/rJB7bnKS+lY7WWsnt72uOMoylMqsSjPyeIT1iwySuDIScF+Z7WoD
L8ZLoUS7xYzx9GTh9E3M1MKNNUroBCPlue7WNUdVshjT8hznbwZYMixwvg9p
sUVCwXJ6YHDYOqj/VRTXye3hczj+0NOgSSss3BjEb2NyIVtsypdu7YpLNSOt
1kBi121nCvTy+AsyI9u6cGjb10sE5FTN


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ckDTQ0ICS1EfKYYxqq/DT7lrML0chBsDeNiFklD1QX6kC7DpswJGPXiqHqPi
mz3yUQS6suazxw5YunOZr8QXgjVxTTqtdFFI/IhFvzoxTQoTmZLjZwZmhTZj
7LsX/jTcyFPh6Ts11Qnz69Qt7ezwYJ7iDCgBFu6E2HkEK9fYe9o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sStqn96XyGTdFyTnB+rh8IkYPPK6h8Dr5mqQrBm4pfVW3p1DuyFFlwxrW8mM
/yjMIB/vmUd1y6UJRh7xlpJ5Tr6raxEjtC3Puii0SwQjIrErDXlpfr1tDSGX
rC2aIY6XEFMzWZJ02kXUfX6rXeH3bzPW//+3NyBbC4WP5riRtvQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28352)
`pragma protect data_block
Zumwacp4+PJ7bSQPI0rFQvwwJN7xZW29jXa8VFmCdIsS8TigZm/d5dD6s7yb
oYNNncvXkcd6pXRkocFFUAlPueQmQIi8KHDsmz+7TQLBbX0z2VT7kZ4DEb5o
S3UL28VRnoRyKdpNXNfDPSVeS+X7HaO+AeUhEE1oH3Yi/xN/BeIXXNthCRuY
/LQ7fdBhYGixCMWPTSI0H7ZEB+5o08vu1efxWjc/NdeEuycx8xwik3pg9+13
s2JUrXJULzq53dIeA/bKY6bK9ofE2yNJy7KOw9tWIQL1KJomOWS5tuFnk+YY
vaq3zJu7w/clHaeNk1zq3nEskLAos1Q5Wtb7oQbHuIlSNvT+XxHXhrZNk7vm
U8urMAGq5B1Uc4d6IImev3YqXMmzA7Y/3naFTtrg4or5Cj7uhFeskiT86X1d
s25e/bnZ16uXskFoaBcmb4TFkpBUqEvhRLO4hAZGd+pgelHEWdOXhMHm6tWl
YPMnZR6DJ2YDbyd4U0lCbibz3DWedL5vdnnZzafH8+xE9W7+OUe1pADKGG7B
zAcwwhGi0DfHCe7bMuj/BzWk3r+ZNrzq9AWwx8Og5JPW+s7aAQZAYH/iaOm1
twYUU9i+qbEAnVYBglTGSq8ggFt69Zp2mXX447cRR15bh0ubTWKKjkvuvXY/
9FCBxWxpnCtOr4gxhj7mx313pwoVmhWAjMwpPulEnNQl8PttVjSI+TkshUk+
d0X5rAJ2VtgTjoSHjsvB4XX0gr/w2RhDJz4XSWFpmJFKgeIjcuJTkPsvGyPo
LQ7sX/1asYBHifAk7qBeRv0C+2jkmGE51i+rUFuvfV6iqs1e4AzhfmSbYtKo
V/gN7adZf8KJrwL5N/8fzkUzHoeo4pf7keZZRDCbDSsKpOE0H36VwdLXz5ct
+Pj+NtHxBdP6bN/3m+KBJxJ2ZyCdyCL5XZy/JMPNlHWJtrCWxk+u8PGOMEm6
Ppse++3FaZVxPGyZ2C+NJCJ9TYmpOEoWFkssONfXnChEHciUfPn886q2xhTF
Cmv+u7nvmcikqn0XBHeYQTw4uJoUCMG3bPu5PR1unhJ8QBsb4aefjy1XyKHf
7sE7NDAlYrkKIgDECy1KB1wQc+gfJztXfSTv1aM/O7Eoyn/aJFMeBiuLv45U
tU7ax/Q56pG/dFVuYsf2GhrdW75QIl543g/3eOdT2R15lcOUGdZQr4dsSV8w
WZFZvw2qbhlqzsVk7T1oDJpRIKTVwCEqw4jTNC4WBUhAr/yAisBZKKyeugYH
c4vi+WCUSz/T1D64c6FpGhvXBeNC37Hvsrl5ru3X2keSSnxaWvAjldvMBmXN
bc4mLQP/k5PsYdU7LGSk8ZTt0uBScJ7mycjrbc2e+UJCnMdgf4BrkItD67Mf
I56NjmHKi60PBcg1fqyybO8klW3fYWxF3bWQ+KQKvUDmqQn4se12Nc97hhZu
/LPELIviqg9q/CBdtt0x8JVpP92tFmMMwSgUX778eDUuLmrxXgetVNVo5+XA
cnghlWKEoxObNWQNafZMGTUwnDcm01qU/NX09/vRtr6CgAbcLzRPK3bdLw+z
IkZn9boYcynuOlsL81G06XMonLH16rH0t8twqZ+phMvKU4xFrh94+v6Tydp8
0ZITIRqHqfiW5Ay0WRMLxuVPMMwoeFtzsJUtGFqsfG1dzQ1gtI+im4IPikVB
pWddFxrBu16h6MBvyWj/LXJlPkOIGJJoETz10/96dIuKDEzWMsD409NOD7Mg
MAT5fhi3/SWUedM5kNYFXRASzmMMNa5+yS/JLhNLixRS7C0x/caDUH4ZPTQw
YCEdj1dmp5v16bU351g5gTLbsJsHokP6oDnYgKDz80fb4e5WxOqJdNyxI8p3
X/FJqHLnvVRivzVJWROUwuLKN9KYjDuZEm5jzWCcR0A0n//NVbdfsAxEyBCA
WKvbLrYO22nZssPMLPxOfdIue510dwq0WLbLNuDw02fbnvHbaoUeY407bFfM
m4q/+z5rmlXfADqae68HWVwNhwrwS49RC0aaRO+bjsYv71kNNzsn243dpV+Y
cFI8VRcbKVY0SHrFHDD80vd6WSgnSllKLBo6dNy6hChb9sfTv1ErzGO4bGkj
NSJB4ByqdCIKCy2mVpgC3YhajkRKRCmNcAO5MpzlAqDIVzhBMrUbqyHvuwxX
vJ2Tb3Xhm416q0JLZZ4TB1I+3OWESSOuMY6fpIkztkfdQZK0NaZkX81FlWLV
eN1IW9Okl1vgrmcF6CeJTVV7nidU4mEjVYxqzEaxCxBk0JqrEnOJZ61fZCH/
lGqGoI59gGpfOZkqCGVuF2Vc0qk2MU3UU7iVZPs9gIEchckb1lXiGU8ebC3D
Em9TVsTStt+LOffiDKbMRxmlaHp+1Y1khefGfRZg2n74gHEBEHhMBhL0mt2O
u6v5JL1PT2r+065l3BYu+3Wn5neOuhmdhWLGOmF7vTeYfpJXPXztZ93yDgf6
sK1ntLdTb45h9mgjnU9P1XpzdgvVYtgInBLzPa7gT7DD6ytsA6YEav6BljSm
K1YaEsbb+5PRMm7yYYOsz2BO1qYWcd4JyndlGhsmR4kwezOGHd6cYAX7zO3P
oUxJ21WD04Fpbr0Rs3xUvA2dNmNsV9/foLmChcIhre35x6y90QyKVYab+KnY
RDhPBtf+h9+GQuVeXGnWOWFF3yXgEAn8f94j7VuVMw33BOtAtLnr9TgrRXln
bckZpzZOzl0qD3v+B1gVaWZTQx0LVjEgAI2k5kXHMKIc5GHTqdmwXw+u9Dh+
LsVNPd+SWe2mkN9WQssDxeer2fqSVvD5Fn5GqHDN/16yS6G+lcPbRyYQVfCU
u0SeVs3WyLZn2UKfIqcnIMebda7men3bdolKWcjyzRogzgvaQj3vrkRZmNGL
44Cj2RDq7WIv6poCxSzNJyJn+iM+dgnW2pebXifa6kc2WdjK8kqyaT8/8nck
he6tafabnQ9qUfbqCpkiNeE0Wy96ydAhp8BAhQLJ+dhIaYsUNCXbqDPpM2iL
UYfeC+bkbhBGQ1kK/eX8De0LhVzRDgh8qenhe2tKRRk1OWNF295j2nnl4Soi
OCuKZcVg6rZEGmH9O5wOBfl10r1edJJJpThFKF4VdD3ytc484imFnp7xOujR
MgNRgitdzEpPqyaruABQiIgJQWY7Clnn0CgB4yniuFR8xqWBOrFdi8gp+tXM
uU4GObDTAvxmZqxlQkUhbeAprTVbGhhysE8MZ4Ihx8WjLidiD/u1QM/wlu6i
PmVe9mrp9fG54TlBwQzh+He/nf+II/iX2jFboAP3tZK7qGLKkIn5g/GE60qo
TtqCd9WY7ThzjccD/Q0j6gj5MwI/PC/EzTBpx0eQWnRaiuEzYEAiVl/UdCN5
yfVt+TZaq7mil/W1hUdIcZ8I+HK/pFnh+lF4oWpn2YuKs2AQRJqqmmfs3qkH
rfIILyibRqqxHavc2gCB6MAt1kcpNZG4pAhoIQ3ViceS2itLX3kcPcyYpEkf
H42UAwaea+l98gpkD6bvQ2IErU0nVxPym3ATn3GohDPJYXx7gnKIsQfbtg59
eU7qWT4e4djSVuxT5nan9jGUtVJMh24eoqOREAwKntD+or/vOTOh4j9MB1NG
QqQ2hCrvrH49z0zoUvBtQTaUT8rvgc0DPfzn9V3LYMtK3FwyiZ1u58jmiE6C
KV50BfjsnCsi6tEh6m8KLo+cuA5rKuLyabjOwVN9lMgpOnlwPmViPTtk/o0x
MRKFTbL3AgH4eRbErBf/Gv4z7y+qCtNuztTIBqtn0elXc7Ni3EXvJpzuBGds
zykmDkuV9T3bQvHbuEJzwQZ3m+CJgjzALvifNacO2uW28GQ0CxaWlvLXO+1S
JzB7jc4ce6nM82e9u8jdlawYlgOj6AAhO1Gni2PK6t9OVrMU4MVUBA8D9yZP
ptliIDkSeFqBqEPOUAGB54uDN/zT1c5a9K4Ku2w5cxes7y2AotHgE4cz06VQ
lsgiA73tmJfE+LoY6K7hnlPYL84voL4z4dLOVE4PWlj+kTHBy/00au9EAynu
wlUOr65KZXEnlHcVzKeObkVwWPA/4o5RJ9VuxF94MlgiZ2lxUzPfJqtR0lf1
WdcwP1Y22BM31B3fKGKURVgdjuOOmB/E/yJVGkDAfxRLL5GPePc5986zbgvK
WeTyxM/IqlswpM7Qg5Yxmf01pJc4SJBJ9aT4glRy1ZOo77MDgdfSsMAzNEJU
655whXO729eOz+99yWyXvU6hc8w1YYsqWo6mt3uGpb7+60XAdTr9x93QQBar
h9Hx6xyRfoqj6a4mOEMypwjq005fm7cwec5pPjtHy3zUmGwE8heNfX/ij+nG
1bHwe+NHIkiLFAwtxEJqW9BKJu3TXkhOvJKcJw2+sRquUO3E1bZwjYC4YYGK
hqcKbB4KwTTtKOXtsuak4dYp2pBUgMx4H8tdRi32mMSjUtgD45WL+8yo1iAn
xn9Q87leATsTSL4KdMw8m7+tzJsh/7s1jMNwv7Fe/dq4VOvaYBBspVsO8ipZ
O/rCh+KIE3pzcBLck2q3ZTQFwJ7s2HltrPE1M6bT1owWzjMRsSELGxv3Ekt4
zmXC0tgnbErLWP9IOALXki04XREWf/SKFEuvsqk4lWoT1ILb0BoLTDbBLMid
hT6ruv6SjrC49L4amhZ5eod6Og3sdhrn5wJzxNhjqGV+kujh8fdt2gnu+zUH
fz8hhJf23qzCNkIcLfeGiJwWEBJYMa8FO7832xdOFW8faxBJfa0mSVvM+Kb5
ivTujMMuq9ngPjprX9GF29nULtmWFJUiawUWiRRlVwabtTX4iRb3/xrhdr57
ZtPeePt2XsymBkKkcgykseAFS23kmzpS1z2mgCWSjJrXiu0xBTYwwwNnx4An
hgtsyUFWmEpySdW40B8m0HI9Oo4pB/5PFts6TK4Pm2kKWlpEhsONXnKUfA9T
0KZ5yNnsbxf4X0jzuezmyqV2HHv0WPl4mX/MO8tdWzuRuqAgBVcIvNdHoUsB
kav0etgE1D2+D7UlqC3+f/uwFreuyUjXWRdx8izjrvPxokePrP9y5mBOBExC
Z4dPYUP+LJb8FkKzACYAK7CnmaRYpiBW8CxkeL5Cl+R9wR/WtGvgZGQrtiy/
ORdT0Cq7eIflYYOJJow44lJ9De7UvzGmrIc+V+nyzL9/ew+Ngr/Mfm3PdBuv
rhcpcFAK6RFSZgAbfndWB3Mpg+wfQil6aLUSGfXsgFKYhAA6quoKbt80/vJj
Cvix9QTI2RLidDZ/jvBfbCvrhbtjmkq1GQPAku1pkLAxLau4evPACn+Yz5Pk
PeXH79pRAVdeIP61INHCC6z3rWHIwXq23I61jQO2y1tXL/8L9bftxOjhkP2G
1qckjrOJtRKSGrl/GazAZJ7ltVPOtdcZ9QoAZlEi037BhP8UwlgXVfDj9xI9
dyAVtlTU9QYeqzOtgeUL10UOFXIpIIURitvUhIed1/15iBxEk/iSSUFMLeQL
nA07vRvAYqqCEuJAOLh+l+YU5f0Zp4egb1TkXr0UbMNeA3N8shlZOeaQmkrX
4GGqvyn2VL8cTIVAZC3UvPlq5Vj4HnR582ayIfBv8dieUVjoMnlb8X6xzeRG
aC0uyeyxBkdPad8CBcF15qWMEfBUbEsXdPk8VhMXVWi/8CyW32bOxAk0jXIw
IMZYT3FnGuHJYT3+l4TzlcoFC3bIjqhf0Vih2wA6QvGglNUURj/552BVEw5e
pOxHGaMno6Sbwi+SOua0tEzHyEHgzETnQvi7M4yniuNFV2YGMwWmEWbokTG/
/O+s4lv1c4AR/VJKSSvgrYnotkMQNy9WhIwqSReN2tlie5DCN5Qy41LB0ENo
HLLJ74UOZnnZofvPJISwth3QfzVWiJwx066DjFkyNEDXk2bgzT3SAgujE1WK
yxG3aR6RwWdSTO/dLkn22FyAlyYLpwsCmXa1mj6IsnSWazAcktqb2Krtt2s3
7IfoGSazkq5Q3u6ZdSnCFEn10CG0adKeSBwwi7D84udNOhEoRz1c1GhERh/G
F0s3pPVLC41QW2JKazLt2YRLULDf3b75XJPfo3E7H4jCP5ekVfiXihf20HDV
2yDDMp5uI3u3NkyfOYrDUmrD8JiXDgbDPfyLAbUGdvuFuDxBav/mcbLNsJU6
d1KutfUaAUCvcPkqnKsJdYzLVmz1/5y5FAQSE2qD+ib68MLpZwkqajydtBuD
tA21ES0/gDNB1KQSl9najG5eXDnwtXoYw5p94QzoCS6v8ZkFzIv8Mwb819Kf
D/ZNZRahi4DLYIuvSaXzdrRgE8dCOpWHsRuY8vtLsS+/gM6jt6iyvILKF5CP
rqQa3kMfB9xyQwElSRgiB5P8UABwn8TCvStxYrbCLU0lERTjyspPcGKbVrkw
ArKsoRG8IVfgn7OnLq9vcWx/XOz1fPD5Gl0jjp6GkyD3m+q4Uth4zgQrZPeZ
oYizJ7LRR8ipH6oTZVkc3sy/oW9qdHBhb4OkprlhHU3REYLuMgWiWaB3kplG
LgCisPvgBu2ONoh2hlfGvVY/upSLga+5svtcqbFfG7xiSsmcYN2T6qPWJs8i
pcN4ZD7Cp10+oqs7drCLyFVzEsK4WxYgEaSgn5yQz1m7uWtASqpYKif+BvlF
4ZfUIFm2xbmVRMDw1Yr8T6QJ7qUEkpnZL30G421azK2ULROjvxrV6kHlDun2
4tJMixqA31V6lIdX2FnBqAPyhY0wefap0l6c0SGELj28WEEAN4l18PgcLrDZ
PdFZqqj+wSZ8BUiGiabB2L59kRDBsYZHvaRCDw3IhELWjsia4g5TkmKnbIsG
/HtUF8+uD2hNw4sVd4+FJiTPS1D8PuZRIcKKvq2h+XJxtiNfaSqBt8Hy+LSL
TvajygZlJ7cPAFezMrZllpBz3rtCDtWYaz8IqpO7oOyYuvbk97M/FpkvYRoF
m81jU7gnPmxfOqBZOoTUtWddiglqjT+4hkzU+iRVV2Bi+MuiyXFKqbAyB25r
QyzB4GDn+9T/RRXjb0zxO+ZVJRLhm4l6yFXXD7NAE0p/sSiesEYc78dHzmk+
rD9TYBpCnzOUghiYVUiQzR9eM3pUH/D7jMqHhGZEDC4d6tgjNRAmUZb676Ol
Gk2eiJvNLoysOEjHCtru+3oGKw3o5o0BH4Ko2Swmbyoh9wd9NmrK8TdUAXKm
KX9r3GZ+AneWXJ36NSg0LiOoOZLSJ9ndbsydvNb0nbSbURg6Qw53tRMmZvN3
Nqh7Btj5DBT4srR4l1Bj7G82FEclkl9kPRJF8DbUv07TdYG3yOm6nsudo6FY
7Cv4N/F8mFvN+20fHypzEEVAy4M22mTW/zdU/F9JC0h+7LJkLUmF12BM9ql6
sQShHFgXqDi8eaou28EAvheeb/AdHwBiTWlm9we8h+HEP/eLzGpMrO799St4
cqu0tYbrMDCX0SMdW3PqeQ0j3FVDUhuRZGEf5JPkffa+N0Y92+4jdhW47NLI
m7AG43NcpNvty36feyyLXu/eH6c6u7q+dVjniCsPhdY3MUPJcrHP7w4GwHUS
ov0mx9p+nAzQlbN9FYcn5VvsPmEnyETehNPHY5ZmxgFV2hHk8oFx15zj0Y1B
8oEVnywH2m2YAq7M/wO6LNyrToww0raJwg1JmLqsUmU6HP4mXODO94zfWQeq
QYhP0Dgpjg15PQVveh9gZhi+ZWFQqXSqi/oRKmwgwxbB5CIrZSj1RsQLJBvQ
etPXivLGTXc4W8AaIGVFDTAuzGbUnRRSHN6P9Va/IZtxU2uGtszzu/8VdmAJ
jK0psOJFmr5ss6UNOw1hn8+iqWlOhu3F6HPy5SxDRC2tGNjdXQGrLa7WJ6cE
lx+VJYI8wsqHmyToW7fomsO9UDdA9MHBob4BCI/HlaPFpXhtB0MT9PwVjcWC
w8eWH7g5njB6qredEtWIajaTm5UWv25O1PDe+E6vn+7iVaI4mAaT6rlOUzxH
DrJbMP5QK4lKbIcqWfYsKhKJWTq52s3Zea71YU2PBWGhAWXBd5rmPXNuC957
YNunjHutYht/bJ/FcEaUKHJnqcGLF7yTjtxGhJc+kgi0W4VIgWVwRd3LCxPz
Yj04qZFBk2WFakWN4ZgVIS+KYu5/nqxhHzHv+q7AJKEWGERyGk9yslKuY+TC
L3LSXNiKMrabb2TB6DiCmHv/+pi9Br5j2GQ0PsYtr++ozDDlY79YliAU12FU
IcooMgk+7s7AsnU1NcScTESzaw7H3GoaSQY2Pa+ew1K4oZqfWQy7VhRoGuw8
6h2lb5jhAToe0N/ez6x5Ze6RiqeZEZ9dG9gZOnJ8/5fD0xAvUUpWOpJud5ss
rOPqTs2xNrK4t3vr5w485gNr8hhjukCuaF5tQ1Aj1xJuNylELWaQgeQ20Tl1
1o6j95K33sDJu7RtxeczyYFs7tdociDMBUeG0RZYCWU3gYgoZLuEZR16MKIs
g5b5PzZlws5/54Zm2IVzYM47i/25BYCY69DWtbwZ1i4k6Yy5hNVAteAP/bWO
DR8HH0THU5FYN9Oz82cHuMUIRTfIw1e9rRiXf7IKJUNaSfzqzHX6KCYPA3cU
F08hA7DR5/QQXSXQ2GYHogEoghZp1FOI0F+QbUGecUz+EvFb7296WUlsNZIL
p1M/ziXZLXV94KPfvjX4uG1KgJ7V2vp/7BbbPETWJGonGv5usO3SqN2TuQei
gyQ3uWSOM0PczHFuPMprkgxQb1cMcpBu7oZFS/i0HuuH+mJ86b+3oeZGnUmx
ghluGBtUi+YMQYN/chAF1/FnjlmmoA091Ga67KPvGhW2ScbaSQjaPeRVKiLZ
96SX4V3TQ3Qa6u7RNp7WpnuwoPlh62/FJFts1gjHaUbcAWtZTx0COjBe/BcM
hvBhKsy6kVgmzSFv15y3zr8WC45TNLlRthDRGxPIJAAeRxOAeqhIlU9Sqme3
gXuzUGh5suf6p79irbyDHb++tckaIIQwIZjNnj2JQCPpEJbk770s5XdlfSIn
N/CwSO1Nbrdq+8st1GHpuV71EdhP5mARZWcaODYRCCwxDhZOfGiGGKS15694
IniPL62P3l985VjdKi4wGv2A1ErwcLUfu3NUmBPpPDfiZG+ICmrDGlsc6r2H
lt2lFsJhsaOc4QmzDX18YMXLgHCF4t+77YOa74cL5mcy7yqUwR3MPULZ8tFa
C/bbO32PcvJMHG8Hkm8cbRwWO8nk6bgPp1t+/RaydBirWXwDdlr/f41rclSt
TvHvxd/0z7uEkZIb0IfTY4vBEzbDI3tUVy6GWMy2rYXlSIFdFxq1Rd9tq4I/
Osb1UNnI1eRFl2UTx9knrHcvKQDtDii0me16TAyIF/lcdn4SVs1OwgxANr31
fEnLX7hR04ICKmK1YmcIQL4PPlAPoR5XO+dz8cG4afZJC9Ozw2uBlZF7/M8q
qWKcW85n50k0GvLSt6CBRjZeEBe8MkoF822NTF6OMaYKy9dgkB67m8EWH4fV
OaCySOQXtyJmKdpgQYVCdqdHp6w7pgb0D5oEQZQH2SfnaTbBp0qBohs7JPSZ
7z+psUJtCQGo1qqOjHunloAp/ZDCFN3znF0XewGNAIDEVqymJNXVUrVlIEZN
PAbKHD4CJ8zdpAHX9PJyWqdupJKfkGgz0KpAvDzxcPjZlAX3U26F+n6bSRnF
Nin0GZViNaCyA7btKyZEbSYe3KyQx3gppvgPBkX9l/QtAm5KVDWZeGnZM1vy
eRYLflcktKeq+dJSyNFolI7bCig3Z1hHnQT9tGTAw9/pGmX1bfuAvRT3cMnv
hZ8zMBlGlDf41OhIkkJ6+Igt3zwiAc4FamNOzZxuy6j8sqdLjil0uZjmauu2
T0eyIotK1ZtZN0ehGV9z+q1lLWgfgF0S9M7hLgo77VWTDXhV6lwxURcRJxrp
kp51IkMNb77KUlY8E8WDETgY2S0dh9n9txiRovT5cilz4XKP2tCUvYe14+Wj
QKSvskBTayeCCDGftJk79l8pzk9STxP4+q4cVQzN7Drk/4k35W/+g4oEOD3p
i92RpfPeOecp9OtzZDE/9cWsPxHM8GYuUa4LJkAiZm8Styvm1bruC/WnBeoV
TVJxW6kBHFm6Aev1NxJSIYztPdpTrq0rwlEkeMa05noVDJ+f+bz8sqhnPTPj
nLmmNfTELnMqJXbX75dAQ4Juk9AqRYPzGbx8GRHT/knyXiPeMRbxbAtzWLF9
1h+bwSMUDW/n8oElHVtyfbE0Lp49nXG/biIUeO2HLojoPB2XjqfGq3Fzyi+s
Xl20/DP1wGi/GxVpXJxNnQ10hcsCV/gHXxdSr/KBs5mWfPZk6AMCs3K1MmbN
uV2TwBa+TLw1duR6lB5/t8BmRVIrUd3PODaKTKrwICQv46BJOCglLANdalgA
xdh9FqVcXvCL6uXi6FN6aea2Hpbs4FjW1AH1SNiMR2dwy0wnFcj6GVAffnnI
ZcV0EQhHRATgbdzJ5HEgWboO4EI81kEryBEL5B2R29Mwj3QLOrYG0gRcbonc
+5IkUNeyhqsdn4FjBSpe4PCPVLLq+8ISW2BMhXCaMdY3QwiyAbaWgfC5kV8v
9+McsdyHg/AL5HyLh5A6yZlkyZAmMM/C2hVZRTY09Fda+xCLChgRfbxTuo0P
ABy8KW2l5XmNomnR/Kp+adBCwrVlXo/iWo6vpBvrZxBKZg4ZMlPMoEvXGKw7
QTD87Z2fXE0s+aPiS1/jUCAI2kBxRxGhYqb9PC0w6QMckP45Dc3suLM68y5W
WOfF7F3WqXPsrxmy5COAmoyeTa1ZIM4iRIfvnPEM4nWvJ9pT+HtK56UyPhAf
e8PgnO3+wllDi6ITB9SrQ7XT2bZlyGD/ZHB3NAkpD/MtAzTPNnQh+NK7QHnJ
mwqH8ggwfgYIVHed/JBA8W8ubQIQOfaGaZoVMpxpnY5YZVDkRSyuivFIviu8
mVLZ3RXOxniONqIy9ilEOALBHnXgo/IhxmqPBK8b1vO/CCXUzPsYogMiedOf
4hpJSnkeb9jHgm0lg2lhY+UA+r4AedIewF5kPbzyL61mPx8hD26hV4FcJbE4
abCehxybjoA/F5mRy9a/h51UGFspuxsKQm6tzul5WF1HQxvSe0y/BQwMWXzb
7yCrszuFxSXWBY/B/pFeeXaNMeTbMupSjejW3ctZFJbvAekClLkprHXRkKSd
7+zCYuZJjxaZim+IbLBnHb+6xbbrsJvjEz5qNDtU0ItdrDQ/+b8oouHc25Sf
+ZBdc713tDXezb+M2WbRZzBXGeoBX/kgq79O5ERUTR+ytr6hCGrkmkx7wrNk
TUUDhx8jM0n6uvYVXEnMjPJDEmTbI2rrph8/Ko6D1bijuxIgYpLH3UcA5lt7
HuiPoiszLFqWZANU936vXdYISutIrYVFAgEwfzy4NZcpZdFLuOUNYzf9Qr6K
WDcqTiDR+L8r2v/WyoMU0/cVXFSaThV9GgYBIJWs/i2BU3gjA+iOye7RnrdJ
OUdEBgm7qhO6LSnQ6/msNJdTAW1D4fGJZ2pi/LXNT6Bhqh3fH4xFtmswcI80
5GBKS+LXpDb+1K19uMu2oPFxVDCMLBJwSAEmfcF0eQhXDINMoo+EXKjXjmff
XcH1rxHEe7Lh7+vfCqSwC593rrsFi1+MRcv3B7w4UnsRGWvxR37rXpstktH5
2PMcrrAt49Yne0vxILxU+gLQ88fTZiKc0XziyaNxCwiOqE6Ge2+VJutfBXgr
8NSXIeakHdvwzJN44h2szzIrtRVOYhV/TrsJLNH+rd0c+Ue3fizbe707niPo
axi3BezQlJ/WhE1BsgDI7cSTo/2n75XSEa+5b9rdYa0Ech3QOnwK6UZP4ZM6
0EudxpkpSMEoPGiVHxkPRVzI7uxA0j6PNy0LiAOPcgAVvGuyViVzwk37K1UJ
kbzb1lSgpWUSHGYELcoWPXF3aU7ViOwi+HlspfIKnwyvzOYOUKVyJupmK0VH
sAfOfqV+Ky89euZ+LV156dQX3W/2WSBG7hKwJJ5W1DVwUGT2CWvEgYrIx9f9
GubnTcP9ts7hX5L0GjYve71MCd1S+YGs9YcjHQJq/XutNjozLthTQnI8gRnw
yC9f29gEYkKNYgukok6RHPl6ThRrd/x4MYWcope9P1ySjAyR/Uc4tNJutEya
pK0wqqhnLtZ9GfRG/MeUSFjzbciH2EcC3OwdF30KQlfdbbIMRvfzumgzqJIl
LiM77QGsyr1R/fzuY2XATekMqOWJ5wkiyzVuFxSORfcJBy3G2EjiUzbgtg9u
sf0wbkvc6niqzzpUE1D8v4+EmTmQyZ/Ude7tanITpSOao5pBOUdgn4curni2
EpmBsOH5oo5bD3r3ytCqdzruAG6B88MDFbHfKXiBG4k352LEaAqz1m3alInj
DZZWl5AnDU93uVseDA0skhByF8TCIIsRYPBNQ3a0VRkkaeh+7DlbjV0uyJAW
RSIXpSalgQWdHhs1cwG6x+fOuZ/MxuT+oYvzqUYM5hc1rZgAhab9trbCFjK6
Fao2e6o1oUwnQwhBPV+Dg3m0pXQP+R0riZeXZPAQUiFLGGbFEV/KRnQgpX/Y
ZkkrxUqqixpEKqChBLIMzDTkRfYcyRvghMNUbXNNUyD86Jp4Uw5R8SGGjXTO
+nAmwbMARTr7JZB97Bod8e5d8jEEquMZzeWz86icioAbaTJH4bCMBQ6uQnX+
OzZsoU6iUp8E2aG9UTbdyTCLZ1gMqv2YhkI2nUkNBlKM6pR8gxotCP8b+9S4
7XbXA3mdF940Hvj631lkl3uz/zBj7lUFxcDoMTflYQiu0NggrpVn2U6p0HmS
ePSkqd9xxfmCDdiIvxsOFlMxuZSjg4lBcHiAea11c3htp5Tj1AGjBQNHpTO2
TFN44XSrXJoqF/w6bTKuaP0yRNSuAfisWZtegiNy0yC3RkvGUNRDyhjzs89o
Il+AQ+90lxSw6X+yf+gEUwKUB1kw2D7PcN94MmjdtcD3wG5swK3/yES+FiKy
R47QVUW1pU/J5zeWwWeXyiVjRUDlIguq/fSoC2uE14WUn2MaMaTIZSSJ0N0j
autyYsjZ8B39GypKh2h4iE9Gr0Kk4HR9W+Xy8cQK0dM7CT+Wu6XQUP35gB6u
rktSTflRh/Eg6zlWybeQU009U6k7yFfx+h15TRlHpcdNvLYyea8I8emhNh7X
HANVofMNeJ/CwK8oyMZmycnDAEPfaOaGNKSmO+YOKFA7YQKnhbZks/GfCGV2
LgD3Vc/7kfZe/Yuir6AcK398/kGsilDSUWU9D3lGu6cFb3j4uIu3nxBXj1FE
24p6dk5i3Yl7DTKgoj9zMbCma0IeMAqrycNBUtgOoQPbNq0wl3sIk8H+VrgO
fHLw7VMAeWiJm1VUnJksGbym6XNfcf0z055VJZ/BMr+CIATWrnrpqtkrE31t
dsJPKiMcDzCOd1e1fiu5ksXgGuCOhQlxVbddlK+DcbaL24JJEnkum61cMXeO
lxOIWtZgSXIpHDIUEzBrTym1I4JsvTd6Tzxo6TiOc12/CoBLJd27Qi0urEli
NqlJRwWZD1DTAkXhF78OVn8+Bdm6k9xd5voIL+X8Thc6rCV8xYwiEi5xC5sm
PKnJZKORtUmB1kjnZybdneISKdiok2M4BUo86S4S0KhFwURjAy3cZ8rRkoRb
32MFXKNFe875HEzZ2seUF2CPqu/mmJqSPaZYm9qRKUF93zb5eIaToBw+O1ss
AsPax0dNTxNGuccPJESFKJEULGEEHQLNt1o7dOQdyED+migc9/WAhXyx/ODh
H0q9DUu03khEdIOLJlVeDjtUhPlHqiyjFj/qNKIli39V2H9G+cUyPAbi1I91
zgL9P3ule65f6uz2LXSdpdKcp75MVHLG6cD5DQvAP0t0+RRyVXL9bfApYq7/
25LvlIL+BteKZp8jSVaADhbe3nERJ5GJy7zhSfS27eIKQNIwOpFAb0M7m7S+
kTHRlvGw7H3ipI05YAEtbI871rXGZXHKztdhDvmN9/6yVjMtUmqoAfiCoF8Z
HsxS9856P/0fh7AGdb808LQRTiZ7NZqin9ClXnhmLms6oLHI00+jMjGkZtsH
tertChsAgFqKJnIDjXsTJIoyLQ6omgL3hONM2MlNpyifuBQrxLVD1cVHtV4f
SioOewajhsTgCUAgO+HQqbHiZwL+2HzO0PLESsHcHvMl+AYUW0WYHEfjptnQ
0yJCXzjUXn+isqd3L9nOyezPcLHndxWpWNHxSUQA2fXhBOXkfUSftl5NJMXo
bHiXgWxc8l+m55w2DQkLBGSE/F8ucJOf3vFf4pl0v1sjchQ+9lslWjFnhLzK
dvB86WvNsYa1/dulSMcrpiauuhFLrfCVd9msL7AXelPRrU6tvTNdYr1obCDa
uxmjAB6DGlV7jfT54q5raVPQZrELTSgOOsxUD4eIKfHWZnumEcIqiD+DvNK0
+iNJKacO8+1tKjMWI3nr8/GusiXDDNLyzIW8mntzT5stJ/I6bJ6IA7RWH9m2
EFYiiqFayLrBqDYkgpOmDz+p3tMaVrYsPHKfGaiN0QkXrP3bynjy8JGCt0Gb
F0yfU5WGykCD/tqvam3HkF46UPfA20g3WTLVZu3o6en/XGJ44ZU+X5PeJj4r
PofbsR8H2bODjp3G6INemBzFSeiM7XvPa1uyNPYYdBk8hDcfDOzfXhuxfHPD
Ko9iB4gM4hpemjOuKd3dtr5EMnOI581R+Go70Ds8TkTXebpLJ2S7fEA7PhWb
g8JNocLWfUkWqUvVC3S2zVCqj9ZAVmwMGIFxNcH2IWwSGWL4VpoJP9GiEmhf
i7f8cDYYWDkcW5dswsGSixUWfSbLlD79s+bw05S+bBBjgNZIA5pfHa5l1nzZ
57KBHgRD6uZK0jeBtURloUvSbVTaNx8yen2r2wqfeCBNrpuJgkHUsi8U4deo
thAR79/kIB8XKkfFOvt8V0RZWCzaNFu8CVRP16NMviPDI/8MxunArmsX3BiK
E7R336PTyk5uyeflgzkIFOOEpOrRDSEFdUplRMOlpRxC/9840mS1tFJuLpgo
0IS4kdoXtwA93LBQ+IJTlP2c68okYMOBoWDHmtQn60bv1644zTzysKOZl9tn
vvPWX4LqEm91shHSzGl/oCd42G/melwTrLBkwBgmM8w0yCiVeUTYnkB7z7FK
20hDwJqxAwLCQ93NK/leZkVDIhnJN01kXimxKw2/rTbYzY9LFLEhgy5bYz39
ZSzLZJDuqot/qSIOQRy+eno0mjxCqEt6hWKZxYzb3A9F3GeKK37hQZ/v7oYB
mf1waMqSoaYH/m7FUhQxB79WoNs5uj2TR53OQfdX/a/duiUVdCYDdwHgw5nu
8/BwKKI3Y9Hs1voG+uYc8BJdvWVyLeNaOFzi+rwqBA7Ubtu+exjdUyxbRcCE
KYe9jMB/sOYkzcK+lSFARWAmGWCk4hwTgkvs5hDWUxwwy3qOoQaUJXSmtW7/
mvDNP7SjdaFExbboU7+R0XHEwnkYrkFD7lL8S0bRkxmjdVS2ovt3N4wn0gIi
foZeFCTDrVSjcxBtnhLYQYechgBNweN8S+GWSCVy7jNch4WuNBFSQ2+kSMwc
y3i2uadEMeCCksK3w+6UoDgQzoyXqXqB7uM7C5OUTaAmwcUkrh/jRhcWpKZC
bkZZQsz9znyrGAXvUci77fx0LowwwPoQi9qThuIx6OxyQUBNXKUcz1JFc+1E
1vpzEWNDLfkcJ4zqho+tnRbKTNBK8Glu7ejZ1eGpPb8luIGH96MSwKL7hBKI
JtLFKBCACg1q3jRTi+saglcsk1Nwen1rvw2dMJjFvC5tMqe5wfMxHgHAtvjF
5HnlpC4rvJLDqrV6iXs8L9ZKSFRBne6Ddp1SgFXAZ3Tar8+g2RudmZ69WbkZ
AbiTctkWrr55OODty1Uvupdcp3WwC6iGz1ch+/rywFKz/LRaEEyvbLaP5c+m
VdAYRO02cloO6RSbSsLG0QqNqUrhtQnE+Qp4Rjq0i0ud6kJ7ZVl/oKLWdLvs
Ci6zCW2oJj612oklVsS8SwEgFkqzYIyJ/OcXLO9EixUW9I1gtsQHutQ36tKt
rjgoL2xrbepPJABPaCTWv5TEhueH6tr7E/OZJOKe9yYa1V9ONDH/1dgcd9HK
aEHjVv1gXglptlVVdQSCCh/AAMypVD/dtLp9cksD+Dx8fj4W8NndtpZlNM6b
8qC1fwsSNaU3GyodPrXLWZftBOqCLWvjAYpacdvaR9QrIqPESxqtQ5HeMY5K
VRSwq6Cb+OvkmF81qjg/v9jfi3mRIDJdjPWkC980zzCvNXlFJlof7vpSCRf7
M5PYpBO3fF6JyKI0wdReVJHnbgGXNe3htN/jihQF9WrIBRGzboBgl9oVCDgK
EA9h2JPLPyjVcsXFg0TvUKqGUL1Qd2XYFUGNVH6811Gv/9YaxQbJJZQXM5qo
V2msVLNah6ke4uLHe6wRc/Zx6jFnK2Q/btTjF2TASy59M782RK7iFZGK9TEh
y5AuTldTKUvoHJ2TVwZSsujVMRPtSmpDtnp8ZwRU3queDHZ/fAEez/1wisbN
j/6opA9jb3foCroaYgBzeMHpFAKVY6TyVsY2dNUgBZAvsA4ZupOI+K9GLtr4
heF1uJ7RND1g3Ep4f/khOwJYm0Yu4DrmKf1uuBy0uxq/No/Kkdb5s3Kh+TAD
ODVwPPF8QEO9tbTKAezAzGHuzD2bgRifaDZWXZy8DBVlnT8I+KQXM1hU72bq
XA7tV6u4Oar/FTOFkbdha6YoYN9Mypwg7jRHb2BcSY38x65es2zHXIFofkTl
Mi1ixuMUDmvOJp7YcS81IR3g81EBO/hrh6LDuimXAre473uLsu0Vy1LTHxTC
BQanI6LX6K148WBl94K1t7zqVneEjl5hDybrXQGzFgKO/pxlx6xqWs7NeRK8
N1kbBs9ue731Abu4iT+Q6qIJ50ICtS6dfKRyxpwErkerer5gBhbP+ysJC4k1
lyHBnjxIZ6q8ZRa8JJlEAAteqtlilqj3I28x8sFnlU/2KTBLCJlfphZG4UMo
oLfjxOv4wW3VveqylNsLqPMw4f4cPC6VGQ2Cej6S5jlMTuW0vBj7MI9+wx89
kBjWOzg6VF8L/0rbQkShZGDpruxWJRXzNP2lc6cGrJpxU4aeY9b8C4oqtIoL
vCuxZwWpwvp+Rj0Sy2uJPGkPbSeEvV9+DYmi7BQxWAaBd0lZBxIATPcAQr3j
EVy+71aeKyWzIIepQF2xgze4gIjKQWOQr2xDOCB7MiK/Nqdc4O0od3UbwXc4
hAfE9qMkwW9+zBJvj/2sxDisfl3C6ToyM8lhMyKYuos/B47hixmMpRKssynI
icQaGu2zUogKcc2wIf1iVV8O61MTkY00H3EuVE5jRyVAjz/TSIXGwn/AXUYI
ySqWfrTvpgS7V3E3PHbg4ASJ34ttyJYn0Ge2+Kfl7b4sAgjFNW0I5Bhl7N8q
9wqir4TZy0KlPPDb04F1oQ+Q5cup37RLf3mTqhRuUxokSJnuMWPo1wqDRfs1
8CQpTYklAIvZ51NqjQXnYk+Mmm+vV0b377kC4Nd0piB0lw2xC+3xh3ZcikiI
a0+8b8NMW9Ch7bXDltGuwtK8iyXXlTk2+x/ptQfbFwJy1dg7uY0zB3PusYAa
18GVN6oCjVDvkJrqK08zEXarKy8npmCnEN7D9O71L80q9Iqhzw8f5vlKAKDl
O2m9LHQ7CaEdo7l3qWACwEJvI5zSCK9JxlBUdKsVplZK9gP3T3sipmwupvSi
mCQmHzE+tI1j6jGG7J52SE360JaC0wmW5PvCkai2WLdzy8i4dbG4rceSX6J0
nd+nPCdTCV45EsMF8RBoXV0aUntn1Iq0SgOJJBQZpR40JeK1bFRmhabvyxfR
9MoOJiYJe2OT/sA9ZJqGD7igx+6evOK35MdSdS4OViS15KIHunR0uDet+x+0
cmCDP7k0OHEK77iI5jifkae/Aku9elPxRab5VF64BU3t8gqN4pMaPQvJIhWD
YfredGlVx5M7AHuOPpfIJ8ValOO00bI0DnfxrhtlvBblxrB2EtqAdJT27KNG
smBHSh8Xig+Wf/PaT2EqAbUpOgPukurRAX8K+tJOgn4lXocbhAAodfhqI95y
gH1IRkOtDJqvAVMQk8NCY0xC6Fuv78nnCzDUHNogTCdIPQ24CHGedCl6kuTs
gMAwoU0hWGr+7qvdusbe1vQHTlAiWZLULYxKvZkEL2hPfoi1RmIuBl0wHqNz
R4zf01cPmc15PW5HBvgQAZCn4G+ExtrxI0I2ONj2XlSMq/aa50NlYosDAR9h
pJPOQlUy1jRE/Jiq2wmKRFPoHF17RlSaXinGmmgqkCx8L5cTBAIPWQtnXLbz
BvzYXR9jLuw0cAnfBlB+3yGtoU2da/POti8uZ+dX66Q6iV21W+bUf8WfCIxn
jie8DqkxNQuoRtYAiPTYJIpZxY1dNfAx4iYuQb4Smz5QqgDsGoNiYqWrBrNe
2E4OQB/zZ817pfrQfPOmreQ7H2Bep64yl58sdyyCbPhOfkS0gPrIdfK1tP0q
SWCsHCv2hMuL6lrJFl467gfoF+jIfI+D24agJDqFzbvPICv0vUK51mHDA8EJ
CH8qWdYLeyEuo9FSWx5rSRRd38c/EblqcTM+O+DBjk4LM05RAfaP/qj0fAK0
T1rlBhAlWUpnkme0Zyi12zp/WfE7T6zBxF8zAownU22Gaqc3nShN1fiK5b8H
gBDaqnpoVrNjLUKGCLdaSu3rVU+TZQbL+D5NPmwYJzM+SVs5Kpm4sy0PqgxL
dUmsUqWPuy1BzYsPcicUkfwON9npkz8JR2REoSGotgYbqLvKaRyWz+W2B51V
yjEn1ig5kwO2A3NYTd+JUXjTS+YH1+ajiM4+TVm6Ho1f5ag+wx1E1kvcjBGS
KuCpROh3Nm4xSxeIQlBhqiZMZ4ApE4aBf7m7Mto0yNbBZpUdYOQev+C6MTBZ
6DebUgSyuIyVolWfqzsIchB0EQwwMnMv/ISUlnfNaKw4s5Q/TVNznSI4lvj/
yeHcaa3NhjAdCFryRc17JDU379fC+kbHEpIeMDLJrZ0dQNBVVyVTsOa0EPZt
uNjBOJCurei+px9hTd25pfERhNcfzUlrQaOtuFpaqxcMkj6BxH+WrVWdNIdr
KyU/yv67+lJikCINSTYd5AppWqXXLPuKSifQ0fyG8nS3GZlv+qiQFyM1PwwQ
eAnK/jN/C3tbNtbXcEFFcJu/LbST8VXIf9gUabNe7cvPSg8WUPCXas6XP1xs
Aph2JMDc4zLPna6SLMJtFdDHkIghV0x+8PhBzgo07kn0CDf7fOUc2ZH8Aavj
JJZoklRGDOgn8ef0bzjCwUVVPv6EwB1+rSws5M9pqrk5QHbKdU+z+3vcwvxp
BrCn4W3n2aQIlAjP3HE6ntoDEhC829vN/HvbDettKY0sgCW1FbMOaY3rLh30
rWi9l3GZycqL7AGJqbul5WoU4ATe+TwK9PKXnCLcxTakF9KaoVL60scZnugL
Eu9ZdII+HEffId7icGuEj18jTAxB0BjAIUIncTcH1BY4iup6j6qaXhQzJYOy
S8vHZOGkD0lOiGeeCwsRFBxW9SJejtfrIm6qQcdxhV4xOfuvY9F8keeRzOA0
5HNb8C4CLosKOY3SDA+kI8BTFunneCBqBkvqcpTP9hdvA5LVNEVev5ja1ceP
Iacht0OG2wT/mpn+vlddlSUSFmnVFo9ApVoJu5O82f8Je2zp+mO1inzXUTrT
UuBDQXXwtN5DvtcxtCApjgh3DWuOdikOes6ud2YkHhBeI2mZaiYeSuDvi+M+
5OD6dkld26Bt88NQ6yqMoxyMbVQk6eCN9C5WFlo8umU0Sfamgpw7qmr3lbBZ
XqW4ChETKXCkhhQ09sEGmFOLrR4++Uug4qW/IzuGsRlowjN/twc7ngoXD14t
Fak1DvDetCyRSs2An3Epr6ZBpZ3USVbRDNljdMjlX35YzDV9bBOmHeyUxe5+
vsB5/hG2YA/FgarxD07YZDnyeld0xfP0YAs+ub3X2ifOuiM+cDsl++lpmiKq
YztH8/LGVnWr8mlg+Cn8sTiS/+s3Ic4icbXAsgZ//3rxirof3gWpXWswR6pL
iVH9Rlss7+t59BRtCPLHm0YSO0Aiy9WZuMt3ar4+ZYFSbtRDDP0P8F/lMWlF
ebZihcIH1POf4ISrFeI/Jcud+EY332sNqEuJ5b9TbEeHG3rZLVBZgv2HHxz3
UvJFPVrT9rQUuChlEzckfUqUxcVOioe5bZEdVtV00GlgZZHp0pvQyO1YmDWI
Z5Ra76WsyGpfDQlSGfiLxMlEyBCdYUZk9pqzQ0e73r6FCA1tiJZqslp8KPr2
X7dhK6ezU8wMDBiP5SxWXFoBP0DM89Oq57eUh2wKIw8R45wXxf07ZgwAXhxH
+zoWwwWEaFrPkbdL4I7nSO5UfBwn58sXnx4WVBEMO5RUlbTfl0dfQ395An2I
A+c0wlAu+m7Hfqxoiy6L6R1OrnPkBMLGC+9hBpOSJ2ay+SzZ6bfcPDkU6MFY
gAYmfqSF6ry5fP3ra/WuRU9FpQYG1lBvffqFlhZ3NIgEWPuE56A9sYUxMxbh
MfDWuC3Ji5+NJW2Ex2/qwHV2BXBy+zHX4Q+HYqo73aC9XCUODg//frSo7QxE
f3zTI54yDQpvCkkXq/cQxFbjRvefb/ouvK2LUx3Hsr7En9+2rbkgjNsuJLtd
6AKaqU9+CRfvk18WD0PASfDgGsiejbLTPOWuwjicoU6k0U5/gF81uSgXamf8
b6rdTsymTDmU/p5kfjaYJ9AT0UkUfmL0IkyMioqm/a4S11nQXYPFLMLRQCGI
G1Lm4XgIE/kcEDUgoWorDR9Aw/kyfZxpWyBSHQSdaPsrwiG4HxncFFkTzsSj
/QpUn2aEa4i7AcXcJga3lH9hZPLk3hHUNLdTW3/7NvUmn47Plro+ccKNrIuJ
JGWOlMo0zSXcANneRmQmRhDoNGZIDR9997M0f08PF+qdXCIhHuBkkjlx9LoY
6QHbP1m/D93gRb3kjcitkkyJWHAYW+5xaiiq2NRPs3KV7vC2oVZbIAsgjo3P
KLPd0k3JBo6c38fjvTIMCK3TAXR7gGY9WTM0gA9UvmQywR1hfp85S3MwIDlo
Obtb5NzjJB2sC4mM1ZxZgCIEPAq+U+xZapybAtiItQ33/L0POobmpTLwFq8B
WEH/IvRgefkf0Kc5b+sOO+6jcftw2um3hcMCEI2jRuirzwLJctKmea/HNngS
MRjVxQYEF1e5BZbiVKSkpNieJzgEGMoyJTL+uP1Z0zrwU8iIUvbdjWDT4WGQ
QuxOGoUc2/kiZZsfoX7AibxyIoOGYlYtF6poTO+GbnkGg9QaGcKcaT0Q1PQC
fVbW5EDR6robdr4gkGCfBIfkhoqANb7t/APYX8hJwl8ZA2bT6NmfJWwhdOTj
HiT+8sa+pD/Wim6e9pikjMXSm8lGRaIhywZmIMk4fKfI5qFB0DjUfyMPAD1S
OejgUw8HUeaplAg9eDXq8mqv1ujAQ4dvf/NvEh8BZZrXMVvUEpr5jVw7PqFK
ELgl0b89uUlQbjbWcXs9T70BOt/isjCx0YuLgNH0W/tXRACNPWYB9X0P35Uv
WEZHFuHNqzNR1YP2YtupA6ZLw3ovJTAUSh6WcXCz/QmBcks8tradCFjFgnYq
ydTOSb8TZjCMPBFD3oe/HpLHPN4F+CS7wYV2LgoH0YFy8syg7bdRSBdEqIP+
J+F0BqsLGNavDU2hoS9fyrJhe2E6PZXPgtB0WDdDk0Y/Ips22a9PohsD5xJH
eH4sg5TN3bEALESwsvwjz6jXJAK2zBzxY4ZUzuRiunQIEr/5vRGkohqBuBkc
ZJWeosJ2n987nKTqshz2pkDHVJDOCQ9wnUEoYd3iEHPw18f1mOsjqd/tEkVv
Ll2flH+Y4umJD9jkiveWOOt58vdCksue4nuiBHsa29U6Dh6zU+rRdA9dRui3
uA0WUqQ/oICbDfUhqZiPHr6U2IHXPJ/xeQI0XgQFivBmZtx1pQ++kL4uadqi
50nCJhgROsmeMqeH46hkbiQWz/F74wxcFzMg6pR4OOq8nLzLmxCnAwTwv73i
AqvbxLVtqVNb4INmTv+dMihXasw+5u+qVTffZU0Qduo2Xbd53PLaUNwdLnwL
hepNGMjkSLyJenOuBcXiEhn04JNRFyMHFD2PiFWxwQeHyfZn4qIFPGGTi6w8
9owAtW4n9473nqCfL05iSLafT/3sj7mS6xNmhFN4PU1HxZRN+E75f15FxdRS
vmZUchiQtRCJxpQyMFvCjhNQHdJ95EAHW2UmNqvB4un6G63c6JDUVN87UmWw
8YazPENgEL9mNM8Enmp2UaoJdgW68fbZ6TkyifhmuytTRjw03sfoQvE/yiPZ
q+a13gRuuG4cibrEVyO4jUHpxRgDLbFy8hdnWW96LbTUhFDwxErEW4z6sYQk
dya3TL6hYYtByEZ0Ppcro6kkEFVIbImq5lhpWx1MEPD+vHO0VqQ6/OFklEw6
RX7mcv2acyK+18KolEulyPz9Oxoxxu9Xl6rD0uKU6GPRRouQ4n1P2Z8VhwJ3
1sHyF1gw6o7XTU+cuFN02etyDQUvBXAbToQEDVgblqdR0Rz6QJIZUc1t5Ex6
VDBLEqcfo8bWGlm6NKnxemR5c9khMq8/b9Qr8kM4tt71dfwSIZQ1IIYMVq3r
fqFhGSHhPTlpFI62JzrFWpHXSvTgAPE/TGioJnTYTo70HtoWfKpB75xmyl1U
MS6Xd8yBGLbsujmNDiFtuFDa9hn94weQ2HESscr+DJA2oDr+zF9gYYuQgvaN
SckB0k0zHWqIwEbuijQBQ2LeUBSCW66cZTtSDGO0QbS0DTOYsDXh+t60CvGg
wIkmh20Wd5wE/5aGMcsfZj4PtNmHHvCZeFe78pP0kaW6afc5hYvs02/x3DUQ
gfBdSbv63srhwEZK1U8d93PehfljrbG9fxxbNhstwS9AhSHGPb8AyRMRBdDC
500lOungLX1JV3yxdiUsq32zuzEkBKUsRbxQtS9BpWMDotLZGljzyTKcQuNr
1yZggqm00kgGlZVJ73rmhfjQisVmURFgMCc1V20uDtjbImOKjLCUZRKYKPkL
tjXEE9DMew4NlIo+T1NZPzCxGSSZTX4nBNFVyu4rGkeZQ1a4XKB2ZPIFWSF1
kct0VnGoQwgLdKbupc1WpV/baE91JBYGcySnuVtLqJ/nWKZS+NNcHhCXfE1A
LRf/tHFVnXP5ZON77nv4HtqeH1KTaHBPAs1ASZJSCKUevTfFk5dpgza8JtlN
3tCPU+YSAck5dq7s7u4kGY/Pvuk8wAd/RtbuJLPbQwFf4+Oir3iY+l7V2aTN
fH/VkxTtMmXZhFdUrQvOW/+oRbXvY5/E/35PLbdLFnjUpYYD4wYSrc5qRLKJ
SWccTscWqIivuYYPg1KJoAyd8++dS0ug699Tkz2SP0OSTwtk701Q0YUbrUM3
mHyDzQEukrLmxemqZ+JzMFISxs+FMvzUzlGRT0u1lD6OdLUMpTHbN5oFzt58
XyQpbhMIllY99fwVqurYknjoxHE5gmORAaNYOaBgVONiX2Cl9QiggS9IE5Ls
qG2pxw4Gj73nfqFBL8AyTJGmkOPo/51YAR0+B4xtP1K+smCZ1KHnKIVjbIUh
6fbUJpgmObTBHEt9K2MmRGX9IezZLQDTcnPmLvYZ+7JBoweH06aRXrA5Sizp
f1szN8ylvP28zzE10TwbYlw9FdWdgCOjnwNWjeg0IxCDYVcYIKk33gy0TIFs
UCxXDklUbKQrDs32CTwXOsYylTkRwGOOKwq5poah89LLD0K5EHbPj7Fp6xLr
iJp5eaY3MGls2w4PZ8DZciG5vz5PrpZKffbh8dv0GFPY3J/Jo5M0UBnFjWsg
48BkYx3tkY3b2HVv50JgyfkQxT3jKf99AbHYXXSS9zWI2VBrSrqTMAaZFcPK
4BPZTekhWCXGMpPZTb3DDt8qeAMlMd/XtDVIKAoCndcsqfZdDgOpRMfqEVj6
vAT7vKnRwnMvtwkLvwTKRdkGFwem+UyM6PszrJdQTFvsDOxmQGrXf02O+k4Z
zK8TxdYLbdYTz3QOACeglclhC8sxePfXkyFnohYouJYf2fIbf0AAo19uNtSW
MAwqYro2wqmsqmFYhptn7Tut87qEl24AmUMViXIooeeLgC46NWYYe1uSL823
yXQEMWJFQVJEH9+NWKjXPxjRpauG/VLIaQnSmEEFAmyUX+6s/xTPGz5VuNTj
JFpwsYwmxZE05K73+1nWdIq9W3vDqZDzebUrZbWVZUQr3RMvXSREbRcKg+HG
wekWVBL2vyhoWkkh+tGfFrtWD5WipmlqGX65VRWwJ0zA9b0xBgYLe0E57da7
n3VL9GYw/b+kUpaiKR1e0w2TsYiIX3ic47ELZiH5lhLuI19uzvLWy8jm1a1C
CNOmfXUN0hR/Z8xV29r2mdX42w1Dd/e56Cl2suOTjKLilRvjKhmblK6pamzU
IP6mn3Hrar8hGdd/DEO0MvB7wGS9l8SboWw/R48/2jq8zG8FNLBWmsGZc5mr
S81NQ7JzjnF0MK9QJkrxRbvJHvv6/gDgH9Qd5ZHiPjt8ZcAwF2jPv+p6oM8e
MU3vdu9Hz/mi80PcODrzNNFnEXGLud0G8+EADia/hDpGF/yTTZDsaoOzJs/e
2phngjedA92J422HHOyCxM90F0IXs6yeqS/yb6DZiTp5y2iu4E4cMgH/P0of
Dx2TbSkk612b5O6esxmQ+jcRMC2XfvDlgO6Hd4Vdyty+d68WsO6Jqf+/btj8
HuqrC1TaoNK/U0iwOQR6Uhx6MYdJDL2UC6K3pFDQF4aHxyesH4oWu2Sw9Lrn
FQq1OmFTrJEy3m/vE9YGVLaD9CUE8PIKkxIMvqtfgPpyDWG/KuMNkOPjkuqB
ok8XEN68kB3pj6ZOGKfPJHhhBPCU+7449C07pmIJtkIOBbAI1yv2QQ2YbATy
WsE/0C6MsIrZCbLFCcuBlekLiFper6huNr+xyFvqwPRmAOe73wrb4mhRPFyN
yZqR0jHOdc4X21EnoXU6mwdxTJyke2fBnYsfQtZGPlSmM6UmzKl2OjO0jMNm
3zhV9Uz/pITFxTWmbQpPhBgDe9b5I5rvPWsAi9JkCioUux6garpE1+JuhMuR
NuBgxi5AGtVvdUTbWH5wW4St/dIUMtqd/stSHb3crHQUb15CXjoIcQStH+wx
gzjdPdP5Zg50mjzrLSQop0U+pO92Mr3DPE+4ybqfIHSxzUwxwiRB62jnTFgO
vsPyJBt05xVyYUyFTWizBGswz3eoLzlvg3Wc7i73IM2awv9FHxujLloMF0zR
mWneNmCS2TgQbaax5az+AF6Pm1vSjcrSnVgSYM8XyDxVuQNjb4nGBFKORzkV
wM6JuA7bFzddBB636BEHaESkkS/nXH29ftF//H0hEmziotGFKA5GHMBs4PsK
Le+8W/rPjI2lReQCX70lfDNoEGUoRtnBTr+lg5FDp8QdgBoMLDKuRhBO1zgz
q7HdPP1G2r2UC7MxzznOqgkBMqnuWFycskQumB5i8jMaxTwWo3l7blRoUSE0
uGXDag7DFeuTy3+zN6EhHBfbaR5d2aBjrgOy/SKU6N8bgS6v4+ZJX3pEiaPL
A7oxFl11UXQkMvugo699SypHvcQx0AvUGjr5GEKweX/de7ixKDnLdvVYFIwW
6PV+wk2TT9+DVkz+ISslzUKPdwyHxZ8rjKNtPD5yAnQrXiiJJaEhZ5WLMsuG
UPaGrLLFTA61bVp2sBCszrsFlbU3Re18wJlxIjdOjpwfEAT1hV0USSk9okNl
DY6AlIiKxqZF1hLYXIUtSkb+7cdF5jguTeFkXgJyr7a0OFOAPlN0GhMvzWNc
aRgEsvsEe9SazW8bca6ueAG/cy+lDWKQr2pHfvAatuVnGgXA5oFAAlf+77Up
J0d36gCHp3Rl1brYm8LIxbPZHojn6l0ZO0Madc0ZbGbcsxFdL+0HSKiJTiPu
ktTnuTOgAGzul1+uzt6NQ/ykW0PkMuPBPJhDdMykMqr+3o8Lri8GMqJ1Dm1T
AKHHmu8ZMlbMkS3yN1TTs6g+1bMan++PD85bc9IZgGCInnKDnTt/ALUzL8Xq
lyFzh+pSt+KK//Kdi94fgyTjw5DAfDH5MTvfJxEAjuPjj2LaXN/dZCigBXLy
0DX1M2lDlLLveict0RXo2UKTwGBhi9C+f3CclGw4T6bDokUeyBzZnCgHdWnU
KA2CB8iuNDGzea1I/WhGO+hnis0kPuxtBZEOOY8Z2rekpGKHbsg+VNwt+uIU
xcluncDpdOBR79iTTyUOgh8Wr2KR4EMd1y18kMkglLzvN9oq+d/7kc+yFVAa
Fby/BJyTSzTNPUZIYk1CvGNL9Rg9fdB9ILXbt3rwZpjQhRzUDgkmZQJLTeQ7
H3eaenAlK0hSlzxbGEYePyj4evxYEss7BFj4ynjy41YZSt9ZHYu3bsORdm4w
uqfV5XHysNlTC1PmNSqXreuAjTPYNlLeQ8/TOa7eOhqquD1Q3ptYkfpCqAim
SLQrBIHMOKyirhmODwD2pGzF7jZL+PExrt7SWu4r2ZRno8t7sOqsJbau0yvS
bVEnYWwXbpWoXJyV305qGVA7SA3ZMcCyTYmNGas405I/YLJlhhkEFuDKCmAH
CsTqBuLOoNe8mEz7/7Pgh+1JPPIw6iCg/5708W3xY4+I4X/7ve9AudbdmNEA
PVbFxuw2uUXDlS6gcjblrXr2GojKGv0+P8799OKRvghLEERyEPRgjFomY+/s
NTcWm/Apa47TVY9JgQGXvF4dNa3B6SRc5HGVD7mcYJMEu2EZxXPZRJnRfct+
i8bTAnnADe4OHlxKBEQKEP9VVsBZyd9VQtiGPgKqV7rpcSy90wxS8W6p0Ki4
CRLJtewrzVrypwTVQsxoTGcI5GdiXia9iPq6tgISB0IP4WUHOGnvCf8N4gS9
IDyGQVyUHVUYF7Y1j6KubsAc87ZZoa8Z8lzXYfY6LHm3H/TMrnnx+cqnOOUh
VsMxUeMm9h2di/M/UknLJaTEye6Fk//Sq9yguGAd5jdKekcHOANtmBQ1IshS
LX5eQ1gpx+qB9uW2eHIJ50+X4DUEMKzAMYKZyU4f8s4xwj+OKXs5iDB5bpIj
nDvKYQiAz1IgGhCKTalVa3/o5sCYnnoyFIcNtEZNOuEgqUssKmYZAiZj1iAB
/mU9mWi+KwA/ZsoJthdvJY05p8zWYVHdmhWIiAXiEKNarkXF8FarCB/6Dos2
zdmGEjDe+cHk1X6Uc+0zXMqzc/xUHVZ+HgR8NK52M1wTVwjkP1xIoKU2K1/N
0BBcxUJ8LDyrdjNGOJcOkzoCK3cpSdv1d5urfgy82ht9WWz+MMQjBUArrznZ
ZSye2icsUJorDLWLUOPMGscvDPSUdJUWNEZ/6j8byZAeP7kNqGfTSrFEhjeS
DrwrZor0QWv7UFXIp/he5DQFBZ2z6NfVie3RW46mNHX4lmVsfF73GDLiFvL5
BYqiV5x1ugqTOHCIgKNEyJcACdh7otjXf0Izet0JaQ7/iJFUzBK80h6DYT2X
OHKbTCkZFuxi5cTwaIguakAtMKy2gnz6yeJJrHNKxCeKVpVvGVH9O8xph5zT
rDBV1cXkL+iZFX3K55GUWdc0x/MwkCs5W0EP55RVYeQQHaQ4a1EIlTuEnnHl
MPIzoh0jbB1eL+FAPn+z5XKq/HRZtoFOWJxkALE9kx8zV8xSR89bzDVw55j8
AAm5tVErV+KFlhPdKy81/v6pL9jbqGuF86nmywfFUB8z+0zHKl/we0eEPQn/
HnKaMpyGzhI/4kprxq6I5TZGOmb9NYmPBxes2Jr04mKiN4JjcIrmE9Nmuz5g
4uGIaL4R9fy2uRiKUloEuETKjv7oCo0GvEg/V58g/y4yNhMyzqBr9taDjFmX
mJkgJJSyZDjn+3FjvfqAtnkz2mSIVSHq1CdJeRVnKd/+RX201c1va+GsNEGU
IAGVjDYUbPKFK0/frkZVefHhzjWon0V0dYrYoSSujr9ge4UUikd/+fmMYI/n
UZ47UywV2Lyp2QwibkvOMZ6Nz5PoGHYdgazblGh0f0ntAbT5hlpGRROjSkJ7
qYdhi8oqiQo2WfJuDD8NxOMfd9nWb/0mBqTX7IcxPt6vX6MKMTyEjwvHftPi
nIyCHRgh2mjFnOc9ZOK/uOThUZfbUTVd+26GrvyUx0oxM96U/wp0+BHlUNcA
KdKz+ccbXOQoXCoIhQ63bRK8SXTazvRJoC+QSiRa7vHS7obFFbS+VUAdzuC4
WAgYOfA35ZMFAeVxTwrPsIhnvBrXXJYKPvzQ0fVk5FEfH0OapdkLrFDyxfyF
HDY027tTh4zSsq443DHfSy6R3mOMTnC3GO5bieEnIgRzKFnom7xtnOhSnK7I
S6fRMQuwx9WlVm/NmnwvkZ4D1aRzIvdhXGY6S4basE8YftEFG8bz0g5H5MLR
+49uYw1JPY8VVWQFJQ7FQNZ0iTMWgViI+7cC8G1e3/ckkkxhR1eux8nQsQKi
YMAWqaw1rECgm+MgpBNfwEZjIbJO5BbijAlqBu0DY7u7WssOYUK/M5JzGomZ
YGdHhCyc4/u8gL8kFgPgDEU5C9HKH09Wq1kfvryXX/12qr5xEYkNR7Q+eAxN
aAlxlnPfCqla91mwBTtoqmzDrvgft3LK+UIZBhMIU/NamUrRstaqYmEpfojS
ikX932syhntcv9T7Vj6FyzwTVKdvgkJJfXeeyVNDKmyfhOTcOmXq9asJcd+8
fpHXuIKNH89HMVzlGbxHPRw6VD1aIOcvejKu1AK3/DJhrldumYHR1WZpEt3J
4gHytlSGmf4tvuF/KsIMcT+FpSPG1zlUyDGlu89QXNBAQAuMsTszneY0JLWM
IPhdYSGHsSIMVCwffx4giCqCKlp8N/aAlzyyCwGS69X3WgfpWFDWhUPHPfpq
YWDnYCCz21NF0JnIduxendDEMHlppjPZHTD+9XU/DHd9wWMZuSA+ygGPgWJ3
gLOPb2Tqt25RBmAtj6TVHy7b9/HG2wTaX5THp3bRt+UYuWCI2VgCcSqzBKaQ
AIaxiTeodqY8+eFdFXDmauuGJkLSO2d2mIQhHwWq0dj9IFW/17yXfs0n4W16
l+IBWBl1MypCK6mLFLHV18uPC1PRU3J1KobvmeF+F+qVNzIK3cQhYJb4D11A
9rc3L72v0QJs0lmoybosYWrzsRrbhMTb7slNTNe5yJtgXUZjvkamu23fm2JA
2XjPUiAwK0nVsSpPWNNxfaVe22G+tluHg8Bk8XtP8oc49jG76RKiEAoqhhf3
p07WY0uXinMbhyaqgmdF/KeT/rvCPyybokcX6B8JseI3jn/jowHbkv8OxWFq
pkbBNRU+AS5RZ2JwNbKenNYcTZfb+RBpRz2sRW2MkKEBJQJnqv6CwlvA8D+L
PF+feLGzkbLCOpqDvg2k/Gp2bzAZwwpQsSCdhen1avKZAs4aRzCxoVFEnZ5f
OyuqylxnP/LOP9cVyBws/+ABX9qk3l1Tr4Q9/xFTArz+8s5DoA30tiwV3N3D
dEgWSiYyqldza6WsNXaQmq9F5avpk7DVAhwVhvtJxeIQPNSmmqXfJBNgTPlS
P+dmnZGQvOD7brb81Fm2QZW6990xbflzAXGEdU+PNhY8B/YJZn3vgJ0bXCCv
6xKFpu8xN6jDB7h+tAqBAQQxIMJVNT2jgZQb0BP3JY96TUEOSlgDG6ElvJPo
ak8emBcEBzG1H4C3LDGdhr0kiEGbltzIN5WuR+zvGPAbPIG3/3pV82yFKWRZ
Po+5rjzQ0O2XYu8ExCID0DkbA7f/29V5E/5XB6veQWxwUSMb50obAfvQUUGM
JOqktoZH5/c6HacLXPiOsTdogxs1Ghe421j1YA75HXv5wO7pmt+AEWS/ACuL
isjEalUkldueB7SpF0MakZlUWSIWflQAGglVPOrEzWX68N5pn86xdzM2dnas
j2vz+Ij8mjUCA52vgqcCT+AK6G/qjK/p7hO2L4Or/eMJHWH1H/ttl8I+59YC
jpXFRvQLi8VeGdeWqzAP0K4aSb3W0q+I7WvYvAvgFPu0KbR0uo0VoAAcioZY
lhaN5aDGi639trZ6E6oJE6ltzHFW0p63UhNM7XuuEfTbYslEsQHyRDeo2fb3
1a4VahJiMcSHfErHzy96mfkOjzTjSIedKgMGhzOHehRU0pWdmjaASI60p+15
9tverpH4HeC3KteN6TnykM7gl/OnM1tAvT8dxg7/ojB0VTx19YJMZ4vGNq4N
5H7NDYjK4qzrWIIRVdArCfRR67xWyHtTYth1SoXLNTWm+drbMapo/rJyDrch
xtP8AKSV/1xVB0pYfqFgZ/1IDHOn9xFqHcP0XbLCKpfaHSO+NH0shR3CE1qq
JI7Ig+Zu521YwMfNnLLPTPWPo+Z42qMWG4/1+4YBUHaZXpF58prqQdpMo4l+
QWOJ2icowqpdslbjh2ku1ENPTpOEovV5j3hlXVE/e5SuqvA0fKTzQZuVoN5N
v2sJFW09D8UerFZbGpqAFp7YqShghDqpuuqp9GHuma9GcKxYPgurbKLIH+zc
sO1g4sNSrSa/JXpk+S0PPmvqiJocz+wUwl0XP82dzhp2Av2vUESi97/3nIk/
nPzd9W+YMrS25hA/TTc1bVI2NkV/wOc0jz69ekvOdE7mcCw4kbXh2rrQZOAi
hNyD4/5T+1NOwpSNCixbdkWdrw6AbmtS4W/c+XKx5/92eRz3CLd3gF/4rDLj
ffI1Gk4A7y8cXJt67bdsCxTetR2EZ1mzLLymC3hFLd/MBJw6SNyPLwIf6HFZ
n8bvrA8v9xg1obASoZF7MJf7l4vgtjjj1B/kHg/CO9PpfmP538kjJ2Jw1/0N
fN698TkNdUyIcIg1gh0ig2rO6uQrSl9Mp+K2d8e1nSnH6A1xYLAR/C3Fc4zT
LQgbfjgeUsdrkXT5LwEPo4qL2h+/XuBVDc9F5unS5QE9yb+6Jtt11F6Jtgpl
Nx8rKDp2EjdVtC/mxvCk4R05PA/PoY8hvh1B+MNb9LXDsXfMZrFawQTPNiX1
eaj8EDC2PTc3FLVm3TCB6Z4euSvla4XLzitws1XdY4OssVwTNaGAQ+yYzefu
crgtKKrp4YVXy7cqOsAQ+Z+ENFwpbrLTHPZhzm9/r81ov6tGgpyqe4TScBrM
Q548Q5te7AX3QuD71mqSgd4h1WQG2zHC/u6qG9yXU3Q/pRV0kP5RSNeed6cb
j3UU3+NWK14bI2sAzoGWnYD6q3E/cIrDhRChQfcnPvFQoHhKid3bd+VkjvzB
ae4/huMNqAgj1WFpdRwLUpX9AkiedrOQsY2MegDoc0DaZYGA1kFrZJKOA5Ws
08pkwqF03vSFHq/XjF4f23hGyYZ8bugzt1shCv094vVXHdHkuDdaG1eQHbxy
EtzvTHsT04+R33NnAdD6C7WAxY2TcwDGQZ3+82ETkAXYGr2AdNllwFIZR3Cz
kyS+fdpK4CfLFJNKqE6h+2h0ycERoF/LNTX2uvfrd++HPJN5jv96o28D1mFK
JljdEwNa7y1qG5b3YHwVethdnXD4WvehpbzjGTvxgQKFR2ks9YhMH1Rhaa6d
GENe6/imvSEFAC5VAKO6UdaSN8WAz3OzO5Lhido6vVuCtA/M16FtPA7IpeAP
VZGzIQfNWNpwst3Er6oyf+K17HE7nb/Ok5BJf4nLDZyFQWZ1uu3xstPI0wjH
PMCIEV5sjLZlprgBBTQcoPxIv7fOOkEnIzRp3mtaiHeRWWsgN7BYahXQkHgv
btSF01hQiA8r04ptgW61Rq282rdJKbeGYQISCiGUGXR+9YC2UzmBNtrYPQQr
bzumCKz9m9R7WDu/fsI40oC3HDve/kJFvDMlpnadt4fnaQvbxXMuJ2idsQfm
bh/AwtasDApNaisift5GcJxmW+xeIjXwisIC3cnsqIRAAfQxoDU/t2CHJEoC
jyDyaSj/si5rITurxsiV1HjvQaK/B2mL196YIruddrgqZUD7ih49zG1Qtlg8
7qeREuRUrC9l7bUO9kI4NpxrsrcVjXOVmznRSZtD0TaFnMC+U3iVFigzdo0z
cMvzNfaJcSX4M28ZdIzhxr2mne/WmPu8Ltw9iyLPyk0+Gk5gE/0/AAg+yvE/
J5x/BCwMu6EfvQItr4wbS/4L1vzgps0FvUAsbAiy7a9NCMyG6Sy7afcjEhJp
+DybgWyhao7SFlwMnkIO5NlqzVJYBGUMH+j8EF9TAaTutq3SP/LDc+Aqhrvi
/vc8fEItntaxIb2V2VbOQl1soydeTP2b3o5qDqmSHC+zl1VwDu04L1/eWG3a
8NldDbcCeV+yJxfZb2A8+LPLTi6LZYCxswSd5cqIM/rz1OEin8dsYPW5iH7O
/zNotB6jG75CTpKCQcaXMswkunSlZSmBpU86XyqXm0vTgEl+qilfJ1lkq9ii
u4f1XRUzyUG7MJ2EMf0yOhi9/Zt+/uAWTO/3q4tSPLFhqXvjKoKg03gT2jQO
EDWA0cYUQWaG//Ef+l6zfJuki0ZOJxiijOC+TIGiOlFLtfk1whwvkAJAZdEH
XBZ2jk7Z37qMitL1c3VhggaDdy9xXweL66hud3Dz4jdXjZETec6oh5ylnQ1b
amkUZO+UNUG+o4QmmsZcNX5CY94jTD1kCxzbZfGFALO0Dgw8PNgfcXJmNwMF
7W4muk9Jk3/4d8mZq+szPCAVunmoTZcI74Jyrnw9F3nzc1T/q1HQWvHAF1ye
FVWs1D5x8yKXHoK+1nPZSR46N6nukcCmur2RDFO2J5M8BVlTwVal1UJKq5RO
Z0VkeHfKZ16sqGnfuMSh/nVD1D2IpiU688wsGaAv+sxZK1CiAS9A7+5V6+Ls
ucAH0R4mLrNlh7qR6uWsxNl5Q81pDobm/yqqJhAeaQh9ka1S4Lofc7CZydLK
Oa/Uhho0xfbFC6Palk9DlE0hmnSsArqvDRB2V3fBNL8hf8/gsItx6ByELpf1
lkmSNC9aBkEmg3kaU2qvFoazBxJHzUf0qkplTugHOslyx/CX1U8qOj2Lh8L9
ydhgCgROYWY7PSPIIqPHdHyxdpIgpEWGoB7GxRaBw6O9CrJd0WKk8kP45/7V
BJ22yJuKqYLume6K19lKejlenGPVUo/2FF1gX8T0biJHBDkrX1euUn0BbqTF
5OP72CP6dI5V2GCkbaU89WtnueqRt7MtixBHQ3wppI074lmSwFgx9OcDf5Pf
gD7jtfA0jhDnFhuN+1kQNT6R/KFK31f1ns3Jq5IS9XQ0dgHQ1eJ75Rxgkwjh
DM4DHVkkznYfq+XQpm7wC6ojlaGyYBF9z5qLFFzHrpYuLB3RR9Fj/yzEBOLV
CsuuJ629qowpMVOIsw/yWtLaRKiW6UC77xFTnOftObO1WEpLn3YnF8Uuz/79
HBZYJ5PVMfg8xKJl0EN9bd1oNRp7StkGH4w54dATw+bMFNGfdiNGmVCzP4hz
o2ZqkO7nT+VbREIphTaUeE9JHTHmknmyZT4HboSy74qWauemgJKyNiT8WhVy
jiJSASVpHxsb2BI2sacV6JdfiT5mAHI3xDRALvt9yCzWp1p8X5kKogELjQ+K
0K9NNz33OnCbJwZJTwxBF6zsS89LS9jWJlHqyjIDR7Qb8Y+iYvkIKddFD0Rh
TuMkn+vUjEBMYj79bEV9u7JFeSSsoU1TAbKjrb0vtoerEsKJzQrsS+4tTwvv
bycTuBi+vvbTTiqaLSXzLpaMsLGqViBnDFpywUXau7Umgyic64bg+Wi3psvQ
1P9TqVpjHpXYaftLj+MgeuGUAGHgLCFU99CwhE/GIfsjUWqYImpHiHrNwUO+
cFjQ3ss1zhc1aerBN2yQ+K2wJ9uz4/szbh+1q3UChguzZE+bqDMBP1viwPu0
z/QyaMM0GBnCwDWTho8NXYht6s+EEEuR0cV9vWoNKgc/1qA/a5t/HHMsOiJn
sbEm80VZ6GwO8JA/Wp6gAsSKDfRAOSCCyGVoaQlAYQ4jqhupd9GXvws9ezdC
YQvaDIfXBqrx6S1TSujrsbOiOLnveK77efQYlaXmHoYtVEKUPrzYPhlgiE/d
6Q9GGaFUuWa5PdUil/Z4oAuw62vMy7VrnakfQ+gzzUzvY84kLmT/Sh1jyigM
hDnduTf8Q7nqWAnc9ddK2zhhxR8IPrQFw+FwXFWtbNmd8QJL1dLdAo7Rujtd
Ynl5UrPiXCHmCcZCk0838x1WHcC0/TmYiooe8IKyMPYRUtTwwFayWWOoexCs
1HzWbO20bv3ZNk3ZnyuyISyuief0juG66WFHQZmjw5hTvo3OkQSpZvY4lBeX
y7i+h+/7AOcXFtnxfNMY1vKuF+D/21EueggWdfEQgK8ef+8B3LWehR7P++VF
vi6N7bLLIh767zRm7JDOHMH/P/6gYDGFopRQZ97Ezw2ylVm7Dx/JxrfcPAof
a4ixMIctePRgQvOXpKs9un7eISvJcnBNOCQM22ME1hPOjsOGFA7jjL1BZBBx
Hc9T20SmU7cO472o7hN7nnqTROuVp4Rf38olOfO14Y01qCKbHoxuqyFUZLYC
YRuwRbxIz/VHlDGdUjfdMfC05xuq1xavpPkApDbJ8wGRZG38X5NVBOpnnbvk
ZmB92hblFCa/rveS1bcZPtkJd6h4LdentritsoGY560oX2FAlb505glKQX1E
k84+4jWOy0ZXZVg+uV4BLga3UqYTvjn0A4430qNF5WXKqrmM0ISVZA2cJGDl
auY2B1ly7SZuyO9zO1NNhTdrI14myrb9tsP7sS5uhcP9NY7rYjIXBFxeCXkh
VteeMsz6SZI3zn02R4g3OXvLWkR6Q6bs1Ep4Uac5fP1s6K/mPs8ShErG8vJZ
0AQB6IVZmo3f1OGv3VsNBbN2fNIAwMIiH6pCMFAuW8RPwrsc5lWZcrWzHA4q
kidwBQ5I7F7T5Yy5ril18Jed/sKLGfw2TWcTk13zbybc18mnOVVZA4n/BYOI
8pYFgR88973yFbLm8OwO68hA7vSWW1tEhrxCrGeT9pDRvxU7GrDdok8J1xWD
X4KWRmJzlGqJd+cYiooK2/RkHy8GZQuM5nAAVGIAuI7PAPGP619rpagqIxhC
wkUVTxFX/ynz+viwruvOfkCetoB0TqXQ7+dHEuierT2NX/7K7aNwBEhQdfuS
LxMrObc8aD/7H58jS1Q2iMFPtsB/X8vnF+iV7YCzgsGjcJE2SkL/sp6gfB9P
Nbh4Xj4qO5qq83mxarUYihqZpqYX26OTwfJZh8cljh8TAjnkVTiRjGggZmXs
+RwTd7wguYP8bsPMVMMjpmVC+5OFu+mpD/UF75I/6sSj0Nez1tSCHTnwhpNK
jPYYEkP8rEtFNUF+2AXtE44ViyCwlqG21InirX9pVilYWtJ5kXLQgBGWl5G+
1V0ecpuaqecELz7xXsR6oauhM7IaGFRJPS9A5MV/eiP+jWBuoXyY0uItYnk6
9BgABGGc6ZtNGS9k33MnHtHTlWdKxL/c3N9SqFL16OMxPIt8VjPdTYHOnGRQ
maM529tNJtV/daINFyq2KZt3SAq8VQdDBX4NWwdr6g3z0EikJGuU6C94szfc
AoDiwRd0yooqlSStt8aMWI0Qu+DOuDNqMkV/ejc5GPIpEZp86G3a/3R0OYmQ
LH7MiL+LxYN1AqdLfkCNqXTmnmC0nUp049VEAsJzVA9cGTO8caAQu1Kw1U4h
Ic3mhcxd1y0Rv3y7g/JIUdo0FdFobDeF5dIeH61GS2WnRn7cMlNy5e8Qd6xo
a525DX+agFgeFSgrCAME2/d74P5KNKN9axeGKiiVpt/NqzFMTbzVMl6YZuzp
v2k08Ex7dB6WOz6IGakOJcTPxphq8eVcrh8SvUUTZoLScAwJaPkPirolWIKT
xQduZyMkMlQrerWMqWRWKOhZag6CimMZ0GkRGE9OLQXedLBBxEZlaxWZ7Yhd
e3PhpHJmseznuJlVPqrfrn/mMwZp7vE84As3rI8a+5tpQ4ZeKfUWF+iYhpWw
6EXxkrWew0yrq1rg3+FGuQAsNR9xnBcQIRmopUpHYv3t+y8RaeFiAYZYX0qW
s3bPbaoeflWetmV0e3YTi/uUv+AixsxY/3N1AgWCRsuuS57s/xHRX3odfnQU
cXNBbOMka73J8Delpl+++dA4KdFXPmUwotcYDazS8IvW1J4nxM8WYz71oSbZ
R4f6Arx/76Et+EDiz/T7IUl4eQ/eAlVCEU9Wl0poZpBSMGdhEIY/Oib4J5W4
pmXzpszKCa/ksXHjAgshjdTuUw8Bc3FutMZlkZiiW8Iw+F56NPpN0uO1Lb4U
ps8pr1q6Nbgq5H43eGmzO27SUsyoDYpIWaywJARmW3bbN4kl8Af4AxtwTuTb
V05+QbrrU/NnYu8qeEUeiATY6ovECIJXBfvGsaMxWR2oDlP1DfNQcZYaIc8j
3pjUqkIpW8KkvgTWztsYv4SLlMh/eN3HGtgXi4tgExOy3dNRDKsFONigoj5o
dWaxUl0FNmCcZWj338tL2/CkBTyVgHtgbhHF0Ak553n+rMGNMKZqW7cMxrKR
hgIbOq0Kw0r7TEL+hL8w8DQxC+pF/ZcjT2Gvd2z9Zso3qfSZAy/Xvp1kk8qK
IxvCMUcfuVCRN6IXTDPqpSB3pqkSTFLdrg1uRoc5uYSsARubKwLhf9q7QDYh
qUEwyRP0G38WlKd5JEV8yCjHrL8NcUVKM6ItCJK1P8AsEALayjdSoB5ybeli
b7Ht0wfIeKNlVYJHKqhUIkOcv5cgFYlGjQaBgT6YWtUPMuBvCKfwoOQDW+Gy
fXCuzmOYJfD3kOjvdJEeiMQzVmHAu9TMOvtIPZeOQE9DShgx0M1pXOKVo7Sr
GdHOUakwgvJw54BpPkLL9BC+0sQ4mJMNGopKUZcPv4AXV0JTmoTzXeUbgFBT
sqXrfYcXYGwO4wNL6cHri/coL6aYStnphCGfoGXpO2t0Jgb/MkEOodp8N8pV
INgGo3ysPZzqkJVnVHkdigeTnfloBGZLNQ6zoOK4GGTUak00ljIitM9uPSuo
OJLkVcowXv6RTzeiSsx6bt5eDWPh/jiUNIOqoIwJGozaa8sxXvZmaBFpXoY4
GNMIuEBihoxu2RVOA4dk6vHXkhDiT5G8P/X4Kual7Eu81tYB/WO9jGtoIRCs
MJV2nOb2lKzN7hj89SxvJZUdsoU+TZalzp62T6M1I4aEKtwaO4CUowQmucPZ
bPR/PSZ2PvxaBEH6to/RvEAEwf4n0ICJXmdg6nPdaD02XGZm0LChfMMWn1Jt
EDy0nUyYdqEv+jFAZczLTQVPfQ7B5b+qsZtb/CG3Qaz274WH06a2v0KVc5Bs
VP/p4NnHRKXBgZZ0e5bzt+SKW8hlFE1eiNvAHABYImygSor+rvKea8WSTlio
8jmm8xNDTgtsOS/AnkkKPUmXloKqhN3nRix8MlH7y7eHqDbmlo6bX4yjg7y/
rA4YiKheOJFZXem62HAaGELL89WndQK4DXl6gr4RZlwSNSK38yC68cgQ/RS8
v54DoJT+ulsISmwXNwexOiin9XsVVWXK8MQ8+Psor8qLdkXtYrcwz70ptXMb
5vE5kWL1rFNKU9YnmWt/nfPO4wbNSA5omJ0n+N3sDfMyH2dKzczEaHFGOva4
90n3lXo+WSbYlTY0H1TvaX47+if5PjPezJE9c0GCcfVlCXErzW6Qu2WJRX1P
asssOdiZpnJovXUytMDq/ZzlfjrPiYn94JMWbbv3ls74ZzZ22BmHkDbOEBON
ZLDNX1E41dLT6RtpOmL8IbpQgi3MtAeOcnNgWve1CBR5sPuAZQgw+2huYmAu
LG3mzbI3KZqJLB/xUbulUH89XxpIJrcqa1qwj1Q/413nZk1gjEShJM+65v3J
/bZUBuOubi48boradsfJRZ4So1lATAG6otJcfQnyTL9Eb5cx2GTZBG/iVk1g
Qo0Uw1n6VOQnNK8e3/tcleJniC8vi/T1nDUMbXT3bq34Uotbtg9eMGBOkFzA
H0c=

`pragma protect end_protected
