// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pYbZ9WCGN0fYCHp5YuyU/sQn32cmpcCa3YpTVpPVt+TqSzya6r1LM4i1U1bbyDg6EV0VFi4qrm9I
W+yrXuZjZH8WI0ybJwD/Sjw01PxoS9V5E8ojy9VxNCX0LtcLk4uw63SUp87olA9MWy06eLHgKfhl
FWIZnvg5r+dBK0MjagbplcafVyjvKqBEobBlsY0Fxzgh3487qeVPjsSpYI1kHULLpKPmuhn/2sT+
Jxc4p6FdFqE5RvqQIpWa5VVZydEIPmAJMkUfAwrtRAmOPZAnqQF1RfBOQNav/bXehKPLiJiabnbd
sF8hLlaD1BVY7a13OL6cWyz92X6dR7w7VY/mnQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9536)
SxEBk86K2C2+dm3YompLXTJJQrrYYs1r9a8hW92fd+7xDsxrpn4MpBphQx2iZ7A8atvyivH2RL70
FD9uId/mNB6ZCCpyjxNq2xvI7Y45yij/y4RQ8npuj9xHzN9mLJQ40acPNePtmpj0Pl3fj3wWEaD2
Vr7mZaTgXkyh6J/N15STXBuXKlmsrP3CH+EKYNzQiXYZvooYVES6tb5I5l8YjIzK/eyFmaHNjIOT
obwKcrbT/1ZQ/kAZYbgS17uWYNMChCHzJoEQkVWmeYdRHnjsclPXks9nzGgD8/4lpgE8qG7NuOXO
xzgp69rxif3rZIEuDr5tJktY1kjRyK6GChXkndGhskbX7CiFBMlknI6ZFZCsmi55rAmPmioYp9PH
LUtOXB5LbuEEyBBw0H3vpfYRU4QPec7huDadZKzylQrONUuHNG6iOjz/FdpuDHm2wSUUKhgupimk
u7PGvRDz/iM3F75SBRvYcUine7BAlKH0RdpYiHVc2SxcTK7j1isfyuKqgpbXr1WuVS07Ba8FHQLr
Qm5HbVfEC4OD850HVVQ4F9Gy7mvKBnNZe+quq5qgmfNc8S8Eotn4bxhXKLypnPQOeHBQGvZXXl6f
ypf6euAJgYvL5gzGt9jaZbOqThMmlcMr6poGuG0jA7HMYaGmzwsbtcsjdlh3erQpN61lOnoorVyX
2y9T6LDOSNMqvhEgRxjuZN2ejTCXEs1NXV/5KqTN5VZyCe9VrXDnxFmo8tL+HrXJZz3mibFmJp1B
wMLibtXEaPGAnVXsVAUxxGXKMWQx9eLRHyt/fKJT9wT8B0649oYDy08NttsBx5+Q6DOrlOm/iAUy
dtM57EqYLmDYooF/o+AKgn5Pg4KSDTITeUEEgnHhtUKNEz1o8XSI0iTAKSyvPqlxzxkPDLe4JGIW
G4r2pFIn7WJWJZNVXIF3/YlYofblDzDySVIPvxFywIg7XHv2yGbI859wK1chD8y12qw9Js9xQKXR
+K1hvTAXaD4rpkJiKsrxTfU2VXozNcQO1ZUr7a20IseEsUFCI+T5VRi6BlJII5M8FkWDslB07FRw
o6LpjUmEnLfb6i3bgWkmXV+1xDLGDuE0Mh/BA/XMlODy2u/OBgsHFtveiChDH3VQXe4MzIFXkpbj
tfWxOUjOjIkFb4FUBz6dEa9AFWE41P6fzNb1o4Nd/UXgXU4K29is/mLVyHo9AMnk5nzSUYMpMc+2
CNLnMLOz8EYy6T6Mok4LhUwPnW2BHOVDbnV4DHrPkLy8RQmwxmLlJCmLqDz+xxPT0vWkuDMYCpf2
DA/3l2lqi/KaeMbBGmckkvEpaqH3BpMFj73Uvy7JlwRXYsOSTM3gCj14CLvzn97RN2wa2KRLQAA2
k9/m9HYb6ZgXJbpkqcDERA1qRXt4euXha2G7q/IuZyuFYsKyYGMfTda3g5VZDKaSAdLbkhZouo8o
/ZQPQJl9GfVDk2+0OUEuWOiyyfR03E2TV6HpdIWaU26uH8+mcpBwwHgWhWMWLrRLcpxzvXjCzMDI
bWYoDtzH97jdEdxWod85knh8AZbdwINzS70AOv/y0jh1WD8hoveqRRD+66+GdUztcnJH8uHO7MWw
0S/fphN4An+WRZ24kJkqlNlWLlObBqwnJKuPned7LFhUPv2GK0OTGdZ8tJ4EP+J9X5zSpSvwmisU
YIxuQNBZ0nH67GvquF3ZLTdk+bTW33uoJ2DEeOEzNrUPeQp8tQIMmHUatel39aqAQwKfvPTdl/Uu
GJ6PKKiicFLUO+RNuQhrp8oyxMH+zW8V3ZY2tnkNw6eKgsQxhvAbnGrnCfBvRJW+PvlkSw6NxIKA
l6H4wj2ShlUt0mQXV1PazoBZvnZ61gp1R57il7gPGQhJdc/UrlTwHH6bj0o59CrowY2b0eM/EKZW
IvIXoA2tUKQzRFoUrWJ2fsHSsz4OryXcgmXQpHApw3xiOQubcLzk9oQK+7HuNH+hruqRAbh1oMJw
EySqVmbm0eJVaMQ6ccsFd3UnYHtqPIOiVEwb4Uc26ggf2YkLo3MlqfJZYKvlWlpRxPc0ZuGzS7HF
kNZhEtMI/3gNmBURXDCnOuGJSaQLhjG7VdIec06Ml+iaWBZ3jSk+tVTEICkJCZ/wO+ve7xm+K4Zg
/4BlmklwCGFc7ZpSE6Ag80scTC3Xe9X9fDCCXkm6kOezhR3BpUYSs8NGtYglOrJeoC4fQ83G/MfK
tZhfhLb9J+GgBDgDJOvuTd8driVFjmcd7G7Ga9x7OwZ9TvRMFmHhWvW2EAKndXMrBGrLP0GP3RcF
zYc+sRNq4oCROiSFRzfGp2E2hsvVVyERY925MENtHgokwaj4pGGsPFhpfKPe2zZT4Xr4KH7VkB3W
NjswyQW57tON0cJv90GpYhVLlleISUmBrPMlyH9c0bYWSTFGUQjKBRNQwx4hHHjL/qbLxRLILtSi
fpyxp0avPDJSmqjn4mU9zJ57LucQlYWMGY5zMZO/lWfjlNgpQj2KMCsbVXNtBOAszKZyYymKKvIi
Pkz4TMSom+h6Cz/gKJ8DDcFx9xC1WpnbzA1wvRQvxJxjrK94xZes6I//ufFp9ee6VJ7kpPh9pNW/
f43hj8QcbkxkyEZi4qRW3Ij5gGxpXj0vTuSrFn/F9pBp+YDJHeFfpuKuqkFiqKSOIOyDbRsNld4t
kqYwAv6p3xnzyebqaRy6i88+WaG+DWMzyPc1bqAofIVM7Gd54k4dwiTPTNHzfkewqzVLgf7rIqmI
2rbmo7ZzoJDna5J7rU4w4y06NRi1EuTm6k7v74V89sacrJoJUtVNio8Zvo/gXxycEKSpnKwgb2bV
5SwZh6sU+d6jLOnMI79KgG7mJj90jREmmVD1hLd7HVQkzM2hx4lX5EDiLx4vrq7Imb6/Oi3JYBVj
nznYnKXyTzy78m4LV3urzJa//mplumXvesYQIxWnG6wKnt3oh++J+w4PXQrTFqBvsZwA946g/Gi6
Da/sSy+fODzIPAMG2AyZR7OxTgpJH+tFQnUuAwMdRs+3DFlc+6um17UZdqPDClUniZMdYOPeqjZ3
lrAjj4pJgxc0ry6w1zhp30UWO/Wu5LDoIvzYTMqPiI4SfxxMu3eVxkk+FEGe14bMARP2AuNyrWPA
iHm4m/W15JIkLtJpjSVR1b4iKEz4zeptLaC9pkuhYyqJaORfW2pLlv8YE9Zt/d1F32lQ7V8aCdzZ
EnC71Y9AJznS6st0Jk9u+VCT/UAw7HAMP+V169K2gC680jSifKip5eRCOzD0ccmZfBdtVUUPg8yU
/9JUda+zmAzZHMYn+Sn7mGg+tF8NXcJgtAb3dHOE33lqmYi1XqwBK7xMjIz+NCNW/PX5d2nZWVGe
Duh0uuhIydUxYwZN8bb/t3JoaNnlwp28BM68jIOQOUCDx/e0+EqKf7IWXKT3JKHC0iw7juAqEcKa
SqB9K0PD6ZNkRXTCWd8DPAQOswbRHK/jvoj2r9CxuVvnHUj1dn7ebwVrhOet7dx7L1V5OEvw/YgX
bpjvyY/Hp0iRtqTYtIM5pYaPEb0xIIclg955fwQq2LgQ13KAGsQyWyj7ahZa7OY2mHR2pO7x7vE3
ewqEJCtZiankBavmqtFaKoJ9PmBxsqyi9xQsfEci2ZuxPe3CvlCDqZdTeMjc5rITOzE8iPk4tui1
/dgbh6wWBT4wSZkLa5Cu+gcBzGzs7c97R5+ZMBIkTVZpfwJ99CEFtrZkRrvV6CnO/nZILWxrY832
FOerOdU2bZ1hC/R5SeeL488EOj/BczJ03GUSqO+ONKBuj5jPlODTYAX8Xag7iSxEBmVerIpXMZJb
kN+8OQjV23dqNJVOYocM8wmMmG8ZHNfyTaczeq3X2V2uvcIjnobiloBB4qZ5DgbibQPqTDUJJ06e
HX3cvcowuimIZkxTADJiUmbP5WmlL9sNe1LmdSkiDM39Rp1R+pl4BnVD7ANkMtqLsXCjYhDuREdq
2kMrMumt8oc/mmq4EODidl71aL7daXHGlkOx+2+rAEmSToXF46khRDNlq+NVKzzgeckCP5ulGsuL
MG7w9w4i0cammo8GAh+2hzvRUiqzsrdGqU6W0+mBCrrNPhajZv+qGtrxA2Z8xXM4CqtIY1ZaJ4bU
HNWc8CYeRT9f+J56S+dcVQNbuvU3I/DyIwcSKLsLxJAxmc0UPm/G+MXV4x2VaYU2xyQ0Lg4eaPYl
+s9bq/lrtIZRlcDtfMA5dzTiRo9yiekgDR1ej0OIT0am8H07P85XXRmc64p3Mu10hlKlw4V9qrWe
cQRpweCm8lf98rncI3wf0K+K0TXe4lsJe+O5RN7RcndN8L7gWx8l1DCw4+Yesc+4ziL2P5/lnLEI
/5OtUoidONa8axH6QrIjqNNEugQGWgqhtlqB4L309thWlgsxJUB+FVhvxvlLnoXV3Z2f0VnaIWe+
OzGRVLK/qC+evnVQhW7z2N/8a6Eq8HKmPcSmu3ygIhv3QOo4gZn7tWOjUm+0RwIwpHrKzLazAZaq
dUKJSLshdAGCZbGJwvV1Z1HEIEK3CSgZEAXxuMmZjQPD6qtFeZLxeOOWjplc3+SzXtJb4UK7lYHt
1v7ZquSTC0pV964BOnhWZMrL9xOZIOL5dJjnyPqZMalmKgcXboRuWqKWAa0Xp/9B6wz5tku+zkZl
lupr9eIZYWO6WYWgsu4jITzy7WBN0MVnKFtKxfBuoAeeMkS6LESJ5DMEpduTSUvpq3+lj7V6lP7a
PkZaf8d3f+rrr1M3w9k8KigEWQ1SdhN8jBjGNywQthizXPMK+uBLVVjY6F14AguvkD/psUjYFFBs
U3COf7ux/uDX25YoyIGDH9jxd093/ONXvwCG5baFRQC2faU4J1GklBRhgp2GLg9BsIBzAt5isCMa
Zhl5VigLNUYzRgrhaqIZMq3nF0VfuT2VDOq5V6fQGkzux56miAuNpv4fM9PT7TOTRLNG/89cAcWh
aZg6+BFMIt8kxVPzj14pnwXOCaBFwhrj95qn/0M0Pdmr+7I5ZEJsfY7BoLtIE/lm9IFn6flsS/hi
3GYG3TuB/W+HJC+N1kGFjB9zZbc64o0pD1c8vzJhFmJ4Vkil12buCtXp31cCaRo210x1F5iHPyc8
siM3pkfTsjJe796dwGpbBZAXEe+tehIsUkVuDZolf5uZtTtN9k7rL1d3h6J+t0vbkM2jORtp04p5
ePGJoztAZwOfI/F/ywikcveW+voyfOoFHKO6N+Ly7uwWUIbtCjmX0WZ8WCW78UrBmh4T2KXldUuk
j1eVDIMwxAVpbO7jd9BbSmErv+0lTtVGAIQbkGskeovECbqI5t94Fz8g5qEfW0CAlDfbZg8FgLAf
DDdYzqEKcaEscLvBQpSkyC7hIZ6V6MQcJnZPKQiyLQG9+alxEK19UzR2kXKPbDsphpOLBwdcft0m
qZG2ndHJx/nciWc/zXCRplWu96BdqCWx+WSPfZM+7mOtlPNdGZHrNpqe3RFLdCvXsT34KzHP94b6
xJVz+fWEieJ9LXBh0OWcc0Ab+IELMNLSSXZM0NAJLGSBBXDXu8cEwKpBYB8lGtdIzhY2xmpzP13R
QBdAwHidDRgldw37Sc5HPAHhZDtOPv7XHcmBxtBtRaWeMJhe+z43BklbR5nTeSzgoIhhJh1B0iz8
nxJNlKlganifxSJnbZ4Y7qMQzgnEWMSI7BYRcxuagXSZzlWnha/7NplgopYrp0uVqUZU9woHmMhr
exbAZv6lGyMW+GNIJvKV5WBTTh8t/5iQ2avmpXgRxhYOWWm53J3DCukKO/G5gMH70umeMtRPg50p
ghCJToWgYpEq1eyMIDmTwYizvqqcrd2wZRx5jNEOI8znoTCJiBVqEZ13Xs5yS/1b5brCkC9MoLzq
QCJO3f0I4zr/3EtfnzXFxo0AuhxXrXZsv7jqKGpa6ui9A6dlXFQLVJSNR19Pn+c50R3QTuFsks8K
169pOHoiXRFti3MrKgrC+AtGGTtB/ADw6fodhXfJQmfOx5j4GW0Hbgj730NRcrEUdq6qCTKMQdGH
1eRTsJ4JjiK9uI0vjVnlvutgS4RaR3ikKrKPOODk9XbsGMbAb5NLpDJudbMQU+fYJhkLyXswRLy6
TaVAAtbdDiRfNh/EW+kqmm5ZcsDxIkkULAgvrlNP0CRSi1uAvlUfidKTTqIBtH4ekq5NTJidI+sg
mW/vbMWTiGWsCpb3+yqE/5IaXNZJ6EGHsXj8QwiGJ6RoMH1xUNO/06oer4D3wX7SlhGsy/UsFzVL
ilUJ7Hku4f9GiTPDkNsuyBpFJ9vlNP+7ru4gIyP2ooiYgJKyV0e7pmBvMsgQukJbXavojRUhmi4L
2hWDf1Fs/Aylxuq5KWDhf5CiJ+QdgAS3VoQcP/LsSKU68g+d4JUNvW1YAMHfJ4QNwSLhsnzzKp5s
FHJljyRUq8qchPbix6Ww9yUbg2jufoj5xC2fNrb2plO2Ic58Q1P94VUCtEj2w1PbjtjPFgiFJp9n
8bXsn/g84NdO64w3xYq2LIuTlsf8GiaUdcMW31lxurebiMGx0R64tGmBu9VrGhqXYBLv/SoXQEih
W7biW3NrH4WafOyn7KUr9B7FG6DybNWFj3SqkM8WdmHmoWTaQxFSO89rApkaSns8ioHw1MSGrHkK
WVS7Czw4Ne3xx7MvkIY4O+WZUXbEkbm2EbH5Ub9ymIK2jJA3SebnQspNIv96qovd+9d5FHCW+rdU
MrP+I69rx3cgLprLPnSLrH9L7ZX+Fm7X8J6TOgOorwrSSDUbOREM2pu744jhXFjEwrIM0Y0PtN1+
lIWYB0ckQl4uJ5ikA/f8/yqYZAqaYt5/Xov0hL/uR9PDASnFnIl5e9P6oIHHKGj7GcWQasbWINIO
p5kbrxY8gJvlo+PkCKUyWWR6YjsfVTmr4U2tDc+Zh6LXGC5e8031/9EyC1byGT43gFFnQixc4efp
lrXoHltOAtrmacNrozA3cRcazQZ7enf/YUUzN5RKHuuaviMwdB1sofp2e6RFePCh3Ea8imcY74Xe
xhdaZpReXFH15tz1WcyMl8MiBVmNeMYAIGVtTtz1z1sLchV+Izv7SiG3xD3FP3Cg2QFoCJ8cFNUl
7AJnHnDmHdDJq+zVzpo/sgmW8pvnEeHPRf+8Aona8KoaMNkJaZyqi+I6i1GOXTkPVk2jd0RCRML4
e6i4XHJqPRUjDWfnuguyJXiptUtkn9i1ZGEwN85NIAmygf06koVWD14EITJWseMmBTOZHg0Lb4ZQ
yrdPQfA/qlbBvpQErGaizYnyk6HzV2ByrMXooe/BNKYjZ8KX4WH7wYKPY/tpW7itK6tR9xMfwv4d
YnqAfEFa3+/uh/u444LL506yGKhCRsT7dWioXXLkjWqcxmyBqqcIFnOaCqutl+Az0BAvVAAMES1B
/Ol49zLzfZKI3bbd06yZKkI5PXMIY0Secx+FYEtkcCNsfUr0O5JWJsFrtU2CeIO+Jtu3FQ3qVR89
ZqytrRJPg8PGr5c/BYgOGhveI5LvLjGF5x5tnslwjcBdbGatVYJg8Em1sW6y/ByGW4neZnxoh4aU
Bai0lZmhQRiDJBS8rgZT1Ht7FBQHg6tgWQr7WdAVjOCM6wjvMcgP4C3qO/cpRtRfOJCMh3U9ebtf
lzBAjLIJduvnsJvAy3ZJaW68B3JMPKDeDCi7z0sl9udyc3hpbkyHHTcPUds+EkdEEWpuP2UXk/lj
wjbgyV6T2HvM0jHJWl4077jyCb1agmrWPLTP54SJsjqRyzwfnH5VM3L0PN1RPjDtaH0gNgyJjs+Z
W9/Azg5sTTK6VKi+XSOP2F989oMMs+g4/RcOBY4ng9DkqvgP/VpL05sfbcPMira5o4cGKkwP6E59
9MZ84AMIsau+gLOr+a/BEC3uznQzfk/T/x2lGiAn5GR4zGBvI0HmY4qO+J+sdLXGKkwl45cCPn0i
HEL87I4Fpfar+GScuvCa3WdaBYBB0IyLrLDccIyq27vE1J3Isg+pLsdKwV4IBSlWhQRUU4EcbG9V
hBuNqqHEHJnKmYYCbj03X+8jE7q5qV+98IXqTvgRzz9/yViQ35WNc75xAgMrQRG/JHlpOjLSuOJp
MNUyNRz478Q8AmLhkBEPD46At7cHdkPZNZfrPXFAH3wMSJwxmeaoAN4Zc8uO/DIFiVHYWHcaT3Zu
UQL8yS2UPSvjcesVDyP2z+MDBBpia3f1Sx9ny7X5DSe9prgjRRbjpjKcpWEOURdvEbYI8nBrBbce
IcSfVHL3DuSt1/+/r1t/x6Hf1/nH/oHSuGPzhCalUfY1rYG8Xj0kTEZpib1xRX1Iw+/miCDlNxas
fPelL3MFUqrBYS6Z+k4SZ7pukX7UpA46535rQIDnXpPbiVGUMtWFnbnGIK6Ky7oOCSQzLLmAhc+U
q9p6n0oPcaifsr+jvuZEmnAps+WTyTN+p8ZNc07w4PL/rK0v9Q+48M5hEum0MOTHL6qimrK3xl6A
kClIM9xCoqA4/KmuIVyDRifusmmNOt3hTCvni9PYfcHWRQHTH6TawWSDGlC/udMH/rSLsT8WNS/D
mDfNuX03Xzrpkj4CliAlMFD7ld3c8Skfe3GCytHwU6nohhU7Q6ygttm05w5QtyqtJGlIIREOEQOT
cDKwqUbpHX92e5u2X9yKMvX9AHQG9w7T5lUE18VHyAtwyw5PbST+wffOTBkHBhRY5GE0BTrl40Jz
12gKFgwUL1K/bqwc6iCYHRsvJZHMK8Yxgqhsh8jB4TYdvD4EYFnMHPgVGWOZJyL9S87Zin4CNxZs
pXZXU8o8C0XzhA54/yDbdqH927W0gZ1odsI1Qtlwdx5+Kh8c/sFPBArk+TBvAi4TOw5rovzo2fsO
TZ/sOZWOGg4TJEwfeB/j6wbaMutUL8jtmrQFbk4WMbd15QISXRAJjztvnUkEZQ7qBsmhOLURGhIc
bo3GSZ6VM/gytpGV9CEoPvItMNgPLMaU50nN6KZYXAWF0wZNP85EXGl1tQDzwu3pNkPbq83k8S/w
pcqVsrHa4v0zD+qkFkN4CFanIY+GnI0JA6LPnH4E9hXP/jMkWSP/ph9g/g2rhwIkNu8/7afeB4Gg
J1ra+TZ/UPoBOJ2eIgEu5n1+YaDeKb5Q3qjnBxg6P1dnPBpPI9me6qdB2k/w118abj/TR2kpVKaO
VH3kF2HmeH71U7aGjCONoNUTctbZDE37cr0IYb+1LHQxGx/bbg6ov9N2bVp/D9BPv7vl3HrzEDXB
PJ9wG1fNjd6OgAcxRwuUzzmSTRK30wUqYZTMeOv60CYLjEkIRNuIt9zqboApvsMREq+S/Sd7BWK3
G7Ns8rpzP+ro/S1fBsvSeNerbAmZpjVs93hwjJgEyhRF7e937rtw/94UQv4dSbEBcZLQaNX1NDjm
lCW27IX8q2895wTB1QNU7wcWmraz/FTUrhKxdtBxoGEKu04FZMfRkWzgy+harqThLgcnkqA0pebo
wLLEiHDZWOoBH1iPVSKwEfP33HaCwy/aoCQaxy/lL8CHXKIIOCfrQPpK8l8KjHq5fzj+Wm9E9zja
rFXmlEnj8T/cDMGsTRo5hZQJ8E2tfPJ2qA6LBWrhZs9LT+F2id+8HOVIvdJO0G57mPmEC7MjaEc0
zKav4lR4iqiB2q5Oy6GjVQKL7QLL6TVl528HSkQOmW0RfOknxd63mKdwAbuQij1aIQSJNp/hd+Kf
mkF8R8vtkHewVIstdvumsYt1XL/X966Lw2l/kMNfxia4sonjAbvcx+H88Hukxin45MWVaSTzvWTf
OSP0RJKye7zVKVaR0bcq3G7EnZDY1U4RFXQVVdERae91rPQ7ZJPVf0faAbdMBXeRB+0nHAGHjVnP
UFOz0azDNVkLusSD5kKFbUXTSu0fXZR9o6e9R6Xa+xCcicIfoKAxc9V/LsIsUO0gCdD+1XjsztjN
hpMoSrmrcEQ434oXH8JCLHUUu/ws/CyZ0goLP9aqtm5Bf75KMGVv55K0aGsi0ci2kfNAitWQVsHU
eNZHaOGxh33niv6ohvfSeBiAM7AJDBluxE3ZVaiD2gxD8aMIEttzwpo4MjjhSr6D4mofPk9ryBu2
RzIvPFjcaT212EQ7tWV2rnhDHZ/lYqSRT8dvCE67Adgklgdb3udE8TpspnIeXEH+t9qlUMbK3297
IabvHVghER8sEHZrkxFJfq81NvCz/8/Bv4LIykYaOCzliVnLb5gSiM5PuT62Xfffj4ZePKDf1ro8
SmdJ44n7SbNRss7i/No8DlbvqiRZcmLplRUdW7tUcKqSRGuL5S2HU//ZzzTIJDpniewB3X3HufM2
nsR16wQ8UkyuAKqjnjIGZA+86DM7Nl+no+HHExvRIXqe9FVhmVXTXaq2jDGztQ+U9FhDGWwcTzCP
iDSf9gEqzdi0o68AlgnvTvn9ToOd6xEuUTiM7VXsk76HUI3b/jMEYcWiF0jaewTU8l2Y88D+JAAH
o41ZtFIjdoD5E5DgBMBZUOPvo1YDjCGNZlLE74CLY6FGtGXC0I33gk5Dr/MaMnOOj00WZTdqtQC6
g8OKTj2Yy/dtyRD1WRCrRThHUG3Nxz0ZojdKimvPdFMCjifHaLAP/4a0B4MsGan3PMST9XLOYNeZ
a0d5CviKWgl6kw3n07Ghzxp53Zk+bsdLkloJRxYoaaFoRjzeUJecMzqWsm+KAx2m1bGnQd4hvykR
HdnRxRvnLaa+ynOhiW44caw+NsCsgnMK9wHi24nICNd69dnu91qEXYWiXNHC+gqUqcDEd5IPr3+F
3cxJoIg+f6qGjmaOmrHoqJvko+UjZzXHxnIqq8pm85r/Dr/ThlgLpcKBcsyenDqAO+n0mWOwB/my
vHsvSHCBMfmFbaldjqthaCHpz0DfQWHaSfKNckzXIE4XjfT9XDJ+5/TeBjor0dsG6LVuAxeoo2h8
lyrDuvaOiLb0MHN+l+tsMGAh63REDna+8aSvwa64mGvkGbRQ/enGnH+atmgajWBTPoNH0ynQ8o0g
fnI9PUF+p0nTVDDbugmP3Ki0xTPZS1eB4DA9SBITlJykVLrCxrWNSyDvJ5mu2oUoIoPbY2u+EpFu
ZEE616X7dUJy+4+YVkFw7QHvlC8FsGTK1yUfrbZ0198nWw+6d9/5rDdVNbJr1s6w8hgW1XHO1XQA
fI2JcDf0AUUgJlzAQBwfp/1xQdGSDp1XsJXPbnKDRR0X/zei05hjsTTX4Ah8URKxcOCNj7nmT9yj
uxV/d2mqDfAt+xCAmc2SSv2c501BLxD6h1jleaLDqtWoMSOTswIlIK+il74OYmAtaugYQs7WZxX1
1bPI5RhwvzS7Oni1s8DMvIt8mTGu+RAEYCJiI88ItrVzr6t70gwzrADJTBG4AeVUyRf/fF41L11J
+oblU0NF/xwZd7ySDOdJkeVcy7UCub0atuWaWhRXr69RhaVNKrILHHe860r4utwmdhUkKvHPTxs0
nzV+3RtF5nnmBmovpsrhbBtKpY27P1mjNxi0v8tb6FzMzefyIUoaxYkF1HkpVTpmIA0FY3ABwKBx
aTv0M30SuPmougl8WvSADa7T85Fjvv+rlqvR/gacBp4pbR+Ds6OM/6libjzj+Cojotzp8VoBB6Mp
w8dtiB0+0cL7NX5lcLFz/WlibPx7qwmZ8UmSm4f8T9NKBep2z8YxeboA3t93sBSETdMEq/05GpE3
vnIXpe+fLZuuWA3AzhoK0/U9HdrVToVkBkPI0Aj+gpU/+juVPKYlHNLCyL4oeYac2MD4T0NTKKmS
jH+Wp/h+Dx+/H0YCV527eJ5n+tridt/qKwinY9o3x69uuY2S28EdXiwZy+c3+srS2lBnI5Cfe0xt
2tkCBugMAuN7RdNt4TR7T8UmasFGlYbfVG1l0hof1kvAHyDkZrtUjiEPIs2YeJcBzeBaQWl2zM8p
623wpinrUvL3fE3pcGqu6YzofAikCbcddfsEdHmDsWDuiaVEhixG6PY89KcDmuAknYG5HC/d/tOr
Kvhy0wueiEHwxOGPsonakzktwZsoA7fkGX0ONczYexyQd1Fqz2v9/+EtW/cjpwJxBSIlIyVg724F
LL61eFQ3A0iIRv6sZfcVIdtiF7Mzx9LK2cUnd/sfrHn5THuH5ACwSY/6qjfwro1xZGX0DRrzfhhS
wmn3pkIcj9iQk+zual2zsYllWCFSe/cs8oTYpEjjX/pUrUWhaVpmkIdnwb0rJLPTD/dfqd4wSmed
9apBZxc8yLPMh/TkPCTYO9ZdmTIEb9ywbq26UvCJ/T5NSHVi0dKk0NtWxO2Vop18uCNS27xxBkkY
midl4izlOJMe+w9jj0QgkhhcyZd6U5Iz8rDA6CdAOISJcOa9BOd0JsSHJh5iE/PGZ8Q4Y/y+t8an
u+HUZqu63GXjpJD52OSptsthHki+HSyk26tPc9fLoonVkl82Chxfa1aLva0J5bO4MN6YnmBmU2B2
TUhGI0lWro4GgSfs3D8WEAmifgZ5yRPvMukE2dIZ4eHdGgor+8+M4H5olsD88bnEKs5aGQDe0RFi
HN+bRWlcgB10x567laMygz6DxCxKWxPYvkShx9vZb+1P3sUWzUp+bzAbN84JmA+mSYs8b4vTocU7
s05CADRkWaYiqeiIFJ8BhHlAbgjRpo9z34w7+G5Zpz/6prO7vCZYx56PXHZGUiYRk3+UdQo8aJDf
j4pYgMd0ui3bG7jk5rh6fGhihS9Qkbm60RfatZW2pm0c2snPmTgWEblMCPY4TuOQUMmtK3RRrP/i
q8mjWDxlEpTUs+DK0kGk+FE=
`pragma protect end_protected
