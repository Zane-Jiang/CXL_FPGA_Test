// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UCT8O9LuT00xKZv5ti5LdNb7Nkx3+i7z7zlsCC8Ee9f298nykrcIsWmFhcyl
HeRq77yhvv+hH9p7J7vOGtOcLd8rzPjm8mHFUVA0XfVJ+m95JBzsStBMSSzO
goXYlK7RxY2Mw16ggySCezvfgKVgg83DlCNbuaREiRLKSNR7IjPd5xJpEhqJ
Ax6exFEg29O6mtKNv9VH6mJhbX8EyDQn4EZy41ZFMB2iL1qxJmbTkHwOBuN7
HvBraaxpsGe9m0HH8acXN3YKYRwMbs7CLkzhKtiWkOkG2uE1Y5yOH6cGq/AY
P/1kuah1sTCH3pjZHhVBCHaMwAMY9Ts235OPxP4bDw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VjSyCF0b6dwvI0ZrysTiR6UAZiM87jNcbgBDBZHiuaBjotsYZRO8fR8AWBY7
3s0Gr0j6NJoIRUK+R+KXSF0FwrQkqyO4nYzNnS/CIzHi8QiF0v0WhEEgdaZt
CV+MtHV6SoU0/c8TGt6jgh5PzGE+qpVlBNsd8bbUNBdg95Jn1+BFwR1DkP0C
8a/Y1+OcS9UheFazTe3oDofevT+IQ4eTSiOXuo/j3PL4hZxh8gWuLsl2H03V
eqGbmgdEVfSV0jbntT96zrccHIypSEcYcvfcu+Cqr3N5Y09Zk4STIRUZA++y
hM3SJbKN5wkoYFbJRYEIXH5lhbUrIDsnukd5nrpxtg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oqOoJdZPVQMWeqI7DMAyLl1hXd9kpiMlbDfvb+uKKttJnz9u2MpGP5rr/AoU
VpmaGzEJxL/qTklHpXN28CirockDu1tGIP5M4TFtL9VqOz5n/oRO9xsdhSHh
ByHOHe9oaqq8ZXaxqT3nvQRiH3pccW3fPUrpygwY1iAzxuYa0KxQVGz/evLw
khvdZkwKmyNnALVBjyjRRXXyAfOAcdy8d9J5J9BpTkYmAdjSnVdDwuwhK97r
nme0u2aQL3ra+pGK7uFKR3BajKmp0I8HZQqV/kfHIwDlT3qTpcD5DAoKgtBY
vh/BtN19u0l/An99Rp80Hjze0M+fN/bEoBtiYsKUPQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iSoN7PMeMe8H9pJq1oHHl2sxeOw4IOAuqGQjz9n/hlHPCaA26uCmDxuGz9DP
H18q/EkdDlLzvVtuP/FboHvVcSUY5aJq6jy9gko4+0QC/kifunGH++RQuLpn
PSf5XYMlyREoXodhQ6rHZTPGdgnnlXkCMq4LjRT+LRm9osQOOK0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kGtguYQGJT08JwkiDUS5/z+QL65QS+h+eXH2EBByt85m8KLZdRt0Ce7lOl7z
bHm/d7s5OWQvlKaVcmmxTYtCOMKjnadk1MJbytmmv6hWDU/5wHfMZ9un5HRv
itopVuhcsbjUR7HlMYDXYosAxuRI+8aBcbisq5qOGIM6TayrksnDPbEYMZSr
3T8VdT4eAbNmbVTsmFIphRx9FRrGbLmg7CCRHaSv7IxPfpYD0qu2/Bw32zE/
Y/7IryKQtWDITOfxZEGW8flfBpeQXOL/EQFIbHejzqgexmIbErRkURgf95te
bN5xoC7s3rpPbPcmYSDxsLL/pGXTbC6BilFohZe6XIrgkxXOlUvT/58RvOcD
6vINgxYV4E5EH51cEes43gxDjPkiHNJPnX5NJZJkBiPYo/PWICQU2CM+8/ff
D3Rr7Zyu8SSGpy+tGFf8DYv6Z6hvX1sAsOhSzspU7XSXYq1tWpbAq6E/s59n
XCRcKVs9b4dI+aahAFRq3nOHnU0XDr2h


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Hualyf/78/yYnRNZBnBnAf/bmbCuPpxm91y09v7m5np06uZ3dg+gJTgx8lPP
TtP9BqMvTnf7X8qDJmjgNHhZN4ehtL5IRc/GXz1Ra59lnrVCpjTOcsLx3IhS
1N/DYExOI7wM+VVTaWoDJSnqoXu8GXMTvQeCKl2Wfi1LKdQnMhA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Gdc3hGTqNRoqiICYnIlPjRE/Q0bPGPrA7/4qTbB3AznHfDVhO5Cxoc1L+35P
QFjjr5dSPMTpa7g8DyuDi/Rz3CVKP340kM6TrmaEg8FRxZiVz6Tg0TYkBvYD
MFcWw9zVNJviA2KxROJNIH2qY9Qq942MqGI3/rMEWdkE+oyqYGo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3952)
`pragma protect data_block
MaqOXxqbxLQmh65Qn6KELbpDHgFCrfF94IGef15Dh1zCHgLdd4AvdvzF1EBA
VbzIvTv5dw01biPulJEMN1PhLAaruP39IY8ueJxQixFQbTh4hloIw7FiLLKI
KnFHjIJRjk4GXiWZVjJlUkz6iS2iUr6ia3LCxmtnboPhT6vsOHoLhLRU1+ca
Gnwp5i2ljw56d19fzMiTMBBGyBitYk0fA/N/UHHlmmNkhPmAOpfdepigbm3p
vNvBfMELVbNIM5cM9B9carK7MhBZIkOd+gLBUaHq0lZCNL0ZJNymsi9+CZVU
oEJbx2+/PfvfoVt1uZKa30TxPyJnrD/RGQIKNjknBWK3++otZR6Y1ibIjDYV
guoPTT3RGXDmF/7Ebsq34vFNCvcfJaB+PGcp1QAGe6E/2Yev2tuG1Q4GsMlI
bqsRWoK8cSUNSkHB6dk/yQ9Mn677xgGR2pA0m+v0eMk7v2x6XN49iISEE4ae
vjR7B3p1K/DfqYvC/JOqFRh1uRQssfKyWMzYr1gbFQXebPDaT0GC/AIP/XIX
pCBBw4qmf46VsW4/6uLivBMLLk4zKfyL17tx0gA7a0zq1wQlFOgEdQIwlw02
ppxHuTPG3WmP7Z2zbgixtDy/iJXRtobQX9x3jdEQ3LUFcvdDhIlMJG9QNPrm
BaBzyQ1C19n0n/P9/S/v7HVydIVpj7aDxUMmRUqXPtuKifveuvGEkoJY2zE7
eZAweVQi3FiKDFbAbC5bDcn/pHEOJ/LBhrIbCpsw0TINouM9emesumZT0t3P
m5KMFcIXRJdo4VGztOxw+ViZbEMNXTWg9KOS2AEne1wtMpXQCCBUAB3QXZLO
JA/ngHojj5SAcKXWHXde3pSXxd2gWagvqHwOspMAluCdOScZw5uw6EX+/b04
hrPmweOQ+9QNBQic1J8yZz0w+wEkptFmx4Ow1HjwfrRie5KTbx4sc068qs4J
v60bUtPwwAbRmN6avDLf4mGWcRvRyvGl1cXDMqWfw6aONrVYEd50wyErAyiP
xvCl7gTrNCb/lBvQDp8H7M36c6ToULR5TLYe47s96uTVWMa6DCXkyq1a9g1J
UMxSjNJzTN7szL480ZB3uTiB6U7QTN6O8/XBStK8FCSJms7Z7dohZzLYXD4v
07631EIRHYLt3PUPG3bA2kfaV2GtcHoWwg9igvX01djaFCKxP0RRy3FxBLV+
ZjSX42yuClK3U8HGTWuw0RgdtkwXxxMlP6Ykp3pKHBxDXroOx+4XdytgFXyb
WUq6rdsv4xtdQzEtAmmDwoM4hyDar87Tn9N0D1rqKsQPk93ZdKACo05Z1ijO
yzInb+HknaNhVm+n8E5xWqIGQnc6HsMfQWQsoRIWdr4CgfqoO3a8f2niVca9
xb8+0wcgHPokRoid/tGdGa14YoAh9Ku1YXM6apXfBVREVv+5AI/D+CnoOq+m
NqzmCGH7I1X8ercCPUfc2fd5AZCTujvQtIxhYvzahkh5TFoCjvpFzTAjNdLm
1zB2775+UImRnzhhn6ErjW3ulYsYBRMuDXlwhMKBGIM6KnazwlmDHJSEi7b1
002d7bGkgqd4KmbACb39FTfNnWrY+ViBu8+VVYBiYfdlL8FTrqfy6gN0dzeP
x9FdfYnv46XIYkbCuHMR1QfKTsI684ke8iJkioPR9zo2kq348w6WIv0dUUZS
jGXdDWGKNjBN5ZwP30j48EcHBuB+1JEWCl4Y4EpfXa3NHr/mi01be5gx4oCn
ecsYe0WuiDZcQsbMM7ZMKcmCVVO7GWgQEF2GzV/P7k/IgdikMag5RI69Btnh
UXjxPX44fr7vjRqaSDhmlALSZA6GtkmzFy3IKphqxE+2p+3ntl/J3K8Ynj90
JaWBG+VjHTIozWW65ioeWw2PHmoibslziwHcY0MJatggDA5UFXaLmxYrU+62
aO9vSPge+XFb2P8On3x5HWKD2THWUzBg014wIYK/E0bssHIVWO5CXLHEqv8h
sWyR6IngfLeqNtLjdcJYEslbz483xurVaE5UksrWWcdBVC/eL9ltwqZSOjjy
Y6s42IUP86nXzl3TiOCAyxlZFVH5z/bC+4GWwaFfQduP+ImLMO/f39Rfotdu
ioDwpB4kqstarOdfS046B0xk5pB8nZQB82/HTdD1Z4/05VlSxsOxHL7qJGkt
nB9j4OqVTXvPQr6Wz157xuyhl+e7EbNX9kE/U+kxKv3IHcaHleN7wqEcy2+D
rbYvmf3npYoGWg7l//InVvkDi0ccoXFiyvYRllcyHcJQUsfIvkLHuRAce5o/
IvtkAioIPC0+oglKx0WmiScCSCSFJm1rltWRa+O5o66IU19nLyeLgqa2yD0p
9OIJ2a+xVTFxomH/kRQHQFK0e7mMl3d+TtTHj/HexMAqim/hS45eScfuxiIt
tZXDh+0mqEEkZaBgTDnF1QQUghDV/4DxDR+4kTCM0bLVoYfOmqVTENsUazzL
GTZOuFkT09/xG8T/X5lsEzpvXLxdheljRjUW2f1INVxAiyREQ09Qw+9yt98y
r9aYfrjS5FVsUQN7FtEGZD4MmN6ES2SB/NTkVqPkZ3/cASBYGFiWJkUThky7
4Pn5IAiG0c4si0rPr92sQXUEL0YlLJsAPRAMezMReAf/qzXheu69WOpBe9EK
/ZKggCV1cpDJwrg/2ya6Ah+fEpFJFY2ZQBV5p4FoUeIxuYNYyiGsPyEgFOET
xaBsAELoIBubfGYY19efF+GN6p0WwsnkzvC8ietooXVhZOEGRROzhbA2sI0W
peG+crA3KrBaGfWX1z2nbcefu7Wqt7SpqVQii1PQ3HiAV5l7GeT+M5Devs1m
52NPUvbGaTxeIg8fjARm/pMGvgywRz0JoqpUL0Gv9H6CNb6q7oSOSSV82hU0
7TY6fyBTntw5kk/OwLUFQfUj3yyC97ItUhwDWFeEMTnoaWa9XZgv9qZ/ZgKK
WB13XTT1vf87iK1oStJZzBFqfzl+0SnwDKuCpu0vnXObLSMK+j8fa8YXFXew
CRI3I9dOrrJ2Lyn9+osTOmI8jE1oi31+y1occXeo+dMvwDhU1+d4y8QB8Cr6
X2zFhgdSBMTEUJSa+kaRcV1UEjQD4c2sidhRXPgsb6XPiCtcz1oPv9LV7rOo
d/jAx97bgMSwFc8u7U0pw3ZmwfsJ+Fd+sdsOSzcdI7u5AUJTPl1xtm/rbZtl
j0BhSYy5+D9db/mjVqjZj66QYtvcBuutB0ccRVslQBFPcoNE2/Jan1ul8OgZ
YaXdu2g1jFF+DHoOxE53/X+XjDrtKeTgUjH1F5zmbz6DPTCaon/y32OY2cl7
vA8Xs2prqsfkPfnjHlsGIuE9rdQt0jwJBP9GETKKXHnPp+EAEx6FbTl1Ghna
4F54aE5ytLA6oYS0NLCQa0Jgd+I2Y0rZ7mraC3OCHfmfTq6ULiIfsvmXmyH3
TjBf6AetaRNyRFlHofUyNjtwa+INFesmmWyLe3MYL7Xg/z7I14EoG/N+col+
/K/FgoIZqSAuo/JCBos2hD9AcIKeQ6HR7gauNCrJZnA2gPYdNgyHgGsaBts5
JmAiAyP/Dy/R3LO7b5vpGvhc+hGxXiB4RbbV19fykAtvyMEH6WXmBn4rUc+2
Xq+TUZhuGn38KHxeQOzfweXZ6d6Be7/gmvQ/NpCGNvEPECVbe28lTUeeJsVe
5e3PY42WCXizwOZ00A7Wb2e64XJ2L5aV0T1WXHWeghs3nmAEyKdMaTVKfH+Z
U8+eAbFKjoR9139UZQN7D9vh1/IzyB+Hc7g+vBxSC+ePCNPxNlWnp7hgTdOd
gO41vs+nJ9SFGVqjIHoNweetpVnonNLspJqUGYhlScxmYdOlhHASkxC6nY6m
PRYjf2VzTLZwFxKRp8o6HQpbRPDLdIBcJd5fF8l5UQLNdiaGTiGuCFKUctwp
pbuCDFqmNxBIytwW57YwazHw0pHMsSVxCaF6pA2/4meIrX6mfKR8RNyPc6X2
fVMheNHH4D/7JujtmBnj3zf73O4JxuVZtrIRDURZOSrWZuGjVMG5ruja7l6N
lcXDvozyXD8XkP+hdnajqCzhDwqVzDDtUngg3nDmp5SOu0lWz0e/xedTFoAh
PMfE7byCgZQVMR18u42reZfJSeBwVE9J9UnJiAXrxV9eDKVJM4ykf3fjw8/p
/rWRwldV+uZohCONKzDa82U9fCLo1h6ziTZYav1vCFXCZDHuI8e1s2ji3Sao
znVxEmYnz2GRYhS78eY8Fkl3BWG0MXYpzDPKJFODPveZcMHQLywCN12ypDy3
suy5EUeEH+TOQuBB3TsJU7nsFSNzAfZPi/mhQi10uq2nGeyLVoyL/Zh1SeWi
gU163PKQxrIkM54D8qhmqO1mLHZMB/teyzp4fCVIMsi08uft55Fb3FmKRfRr
zHit5udjeRYX1DABAe7Z/q9+UTcLlwJ1t0fxmjQqGY+hydK9aImhx/4gFYLj
iKV6ocvMCvYDW3Uzre7yb+VdVIuTVyNCpYd/mgUlfLqu/4UZgztwJC/rGTAf
v+1f4VGOUyrTLtwWdjDGj8RQ44ZZT8vxCK+u6rO9/hy+DQcV0w4gTNXLpGbl
JNvSrXo+vObABaG0JlUh7uTl6ccEu0VFKWzy77c5s0D9vdoA5uI9gHcbSEQk
7Lp6oKu65ew5WCGkHPxBuEmOocrSE+8BC92nch/H6VnbRjnssK184s3IUzbA
SC/5WXd+xRIZiN/OTPhS7lmirh5PSx+SPk1/tKJBsYwOgJGxEtdZLS/n3hJt
bWa+fcZsT4gShYatUKQ+9h1C4yaZnAXqWwENpR88MNUAbOwqOV3FAW8vKXjv
9YYyctLzzl2970OadUTRxv/VHD3TLr4wUEIA+L1VQJcMBXNHzDjaWqsOJh2Z
v9LKy81/0Ze+t7KTpqJGTxs+58z/RAtgq7Ht2cihSmhABCx6yExj2snSxi7g
QcjpY4+YRwl6RNeP13Ynx9gt2VHbkI4iXDjMGLWf1FKa1FZgFlqWoKaqNIFT
W4TCvkRNtp6WKLXOFWoYvrYqsE9Xw6BMeF48I/09tP3yNzlA0JsKBcJh+Kvn
LQaLQfBn4P9xmj4mqjmJl2iDqou/ETVSjjqHsSAF+UeFgMiGpMXhHrL1MdV9
hIOgMaiQQqfCi7xgP061UzIUjQXBQH4yoQ+AWOg5fFPq8xrxDK4TneTdKcIB
hNn3aO6WhEOuLSP0qEMp9oKbbaTBusVdPfpd2UFmzGoaIIV7DdATCd+cQhmj
G4qLSZsoqjRIApqS8P6LrdWreZcQIEu9PlXZn7w4OsyuNFwFww==

`pragma protect end_protected
