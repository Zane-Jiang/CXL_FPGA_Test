// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
l8nE6m6Y0uXJKF5ay+8OH7u9ucc90YmbS49nAwUD99aLlJ1o3z4OGa1vpDeTgmUQ05LUwmG6uxKq
u5Qu2rcqo9HdoDcjWlTKhELpSkvu1kKI0Zm/ck+WHXQuaKlZe9upZxj6RQpCdNQQF0UYYtnOLWr/
26PtYsC/AaeG2XuyGx04/wjjxtLUmTKbguQHyXNR+UGQcQl70vJcJUtZUPPqU95yQFLUCoZOyF0o
JOO67QdmWItHDKP1inqewYfZ5qkoIGlvZQVHinqTnkx6LjauC0/GXra+t4OWq6wRfdJwcEceULL4
mc3VBf7Xzo2omHlyoA2eHw//5wt9GfMgXGPCYw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6896)
o2yIVmV9NNl3c3RSXXCr7CM9uxGcYgKG0HkMzg2G44A2Fly2Dsk6e5r3qQoAeWRYVgMlzwWxCCUi
AWKkSwqtWxNnQoHJJWbvvp5DpfohVk0Swm5NeuhFJ2AlDcgwXufxqoPqv5vGIEdSqNjNtSuZJVEb
IzCnOZeS9fS4IpnxDk/jIH/0WnEtyK3jXqZOemfyoeT8zx4oK618GvTQaiGoG5SimQKQYxJ3VeAe
B6JSpMZVCYptA8JVKpvcQy2I8XtZU4YymImylpm/d5RHMVOHU+/QsT8GGWlw+to5JliwpW3Hd7z7
TvUiM+joBzmNZhNuT+pm1YqaP+XSMUoZhFO1KmYHT1Kz+lYffT0zFkCkdEotudVoO6pfFrDVuH/p
Pi/yhCS/rmbOYyjADN5N0l9ZYHlk3Z6aneclnMKYfzTA/MnOQHRApSESbp8TT0/hUabOGRyGa24Y
jayg66mjKH66cOP/Qf8mIkGADBa74WRnCa9c8rySuuoniVr/5LHvqoc13ZkZ81b5RU4qTlMx9UNW
QRrOqUsMBOIJ9VyZhSYk0qJgKzH7qJZFiZ3AG+kxzS6YKPcAPwcYKaWkgjPSYxkoju7+efhjfJbc
tuPw/HIEl/WZYupVfGgr6gdgq4pWavSS0EqArPePTm73kj69hge2HSp41nn4fQ7TjPTRmuZaRo5j
vnOazFNmR3yat+/A35n8VTqG5kc4ek7icVX6cX/XayMkDOpckFo5kn8Ac01X9kb/KsUdZuF/vKD2
qDM6r3I+IScVzYsw17iyiSS+Zo8tkjXhES/lc2XxzbsQD904GJ2nZBdShvaHQQZd88ggw+lCFW0l
tgvZKWV4C1RSMdN87QdEqfR7CEiVLk7d1jbp2bkfCjjDtmwTXcD3MbU3fIj4S/pucDSk9/6rtAzu
f6+KQapO1o3ykPgpv7OART7TVvSbgzPLKkoAlGor0QhSVt5zv307ZADvloJZ9Ezm+0Puqy67sBGY
dzzoREd3CXx6+akKbeU7bkxC1Mm5Dq0wnrIDLU+55eqOyU/dgVBawOHfSmBGDk4Akw4oeFUJQmmK
MZNbimS1DfgCyQOTDdadVTfCTiI0Pa7HfjDnMl6MuyfzPoZMIfIfAMMXK4t9yQZInPXk/HrR5mQv
GYu6ioqu9ZJEM8oYnTI2U095DquWTKWo9+0s0gwBKQstHbPWmQq2dcgnMemxapZ4UuvpdHuUeIA1
UTfVI4h9OTg65/6huUsip1E4OZAxWm2mj1nsW7IMaresYr8kvWF5xyeVHu5/B0E+7y3oF1ClKNwN
CYruWBCbOMgMmHoQyZjxSZPJ7TG7jFFslaqRpzZg+3Ja1RSlQgUdvtMtLZY/3SFXMYh006pgXOHr
unE687S8gvKbZ28tDpqNovh761xtrsLCgweVyzWtqa+PiAM5lBgyO19gA6Os117C7aTMjuyHTQtz
UjYqEA6cUyqtwIyzkrpdecTrG6+oCZEJ/Ekg1QSDT8B0Q6VxstTJY4E2jbrNUSr3eFkHEmhBuZmN
bkWl0prUS9A+pJIVZBLeUQazl9PI8ekNNL4BDHSwgwnH+JPvfnEv6jUtEybR+Do8cjuzWo7Jc5mw
vy+kLkp1hB+VccqLpesFlQCCW++UniFXDwS/n+HiEIOqnA3nL9L1NMagZvJrNhH1wUiyZ7Lh+/Kl
mIeCC3leicRVWkMr9a1Qd825dD+F63bvImcuOMjRLkhHiQmWnhB4HChb1l3xwZuWvfoUoHVgZ7S7
RVklaBhnM80MnWhi/kVIxciojeHFvlN4a6Soc9lefDB9OAmd+GnbNgdQ7SUdcUTqLLtwTGvey5On
z7dfR5NAz7zRQi2to85wjHighYExlumLVH1qVAN4BEXI7DkFeQI7wtqEG7iGKndtR0VJNrl8fSBy
shkObOm8l+MM38v4/7/ZccJ5rGxf5MnFkU0mL/adtB6Em/HqAYeNi9QRfZsUeSiE761svjv0ZkF/
x6VUUyO6JO8O7IWRtFZqxTLrCN1TTMsRCYYmSSoBh33NJmNEQgVm5VTYXEXxOHGqtm1MpxbkeWXK
PHnB4O21EgGgSOofILzt06wRdABBtjavCxCXYFciyJ4FFUTuQBbfpfHANPziH69SUCyNvSuMb3PB
XSbofDhO1wNfqVVk4HN7wMIbha2aqzbdFq/VEK7Toe1uZ7zHvopmaX+HNHidFswF32usvO160FeO
UuYXdD8lbm7AkMPb620eJiBG7LxGbCmD7/y2RFHLFqwjP8a0vB6/R4E74DyX+g+IS7Uf1qDu0GIc
DB3jgbDHrO0h1kSXXzUo9XW10ENndbByYEqsbViydrjpE2Do5WdqhcyJ/JZX8t+PKzU610qQ1wu6
Ygm2AiCC7LKAbp0LlE34qOxKSmWdwp7x7PumekOgOMyMCLUs1h6U8mCLHA5JXupX65RJo75noghs
IJH9gGgHlyp0ivw6ygT35WC80t655T/8bqll8lnlB+7cLx5O2oE39ti1NpPT5/q4hhNXfj4h/Dfb
KInzc/8yf7m1/+NF5NZwt4HB0Vk6HmU4JBHUU4NEZcRDtecrZxbfpha3chcaec5hbZHLharXsQJN
C8+M1ZdCFmbWckGrukXH0Rz9oYMAH6d4HQI+i48uGir8yxVAvuUGJ7qyZBPscQcUREM1GGJ3Guhr
aaeqHR3MA6oQXu+MVZdWuaf253dDWu2lQrNOArDaUuexhJxX7yL2kPiUCMMe3RP9SW/M32J3crT/
MbW27BI7FajDVooES3uBBDEVSCQ2NHy9KMTrhIvN2A/ZgY2nQ++GjAjR8jkru4O8BKoMpIUGto4R
oCT7Wb12DBc2KgyBNqqKk/3spuzaTjQBl46isbM2FmDzxVKYzVcaseloy1tyLxzTdwHn0CLMb5N5
sZslfw4hIplO6i0Brpc+MMZ8/YNH+TNOcW9y6xBd0TJe1zEEyNF6bRvZSwP6jCPhZPrHIs+l0het
EOHDuypSTN6J7xpM50P+KNMn7/krVpFbV1LgmgfQMw7zq7pZUzCZrcBASJpJeAiKz6Z5tQ4iCqA0
3hd2KdljRbA9KRgnE5ncEPsmFjf0gd3vbXT6oLTrPBXlY5kHcVDjcttmY6SBDydzXfbkqDDWJ8oJ
aeQ0QhOV82Zxsm6rvu5a5rAoRwr4lFwIII2mI8Yd82PONx7wb/d7errjGqDEpXd1fOq5lo1we1r4
AboL8fueUIk2PBkQjL0+5W+rhUwi6efdWKJtp8AE0kCSUaZeDrcVTpPOg60vL7QmoGR8ZQgw0oxx
/gZYihYUI8yix2209XV2SOkFj9f0IT5+TZOHZRjDvMUau4sy7wpt2VmvN3sF0hm60sWttAkry0U2
ngb7UZN7NXhKCKi/1/DeQ130UShgrzrGR4EL9JdyxkG1RKLIENZWF+jBPwNCA1zS8T+pbkP+TxSf
2v9Esgjq2ZSRs83M2NNWmAfHbu9jZZ/Qbl/2uMloQB3ILDqDVqwjhIlUPdIcQGskSjvb6K2/ylnP
hOKCBMQRUl8FnKWC0lm+dRtZBV4MlZKlIzfu62OXpnGd6EAAAlyIbF/FOqKwmgXPGFVJk6YMhNnI
wk0OH6h45F1EN+Qvwh3/8hXf5PInT92BHLhLXePATKpXWtfNqJKYN3dXIZ3TcPndY0sPVKPeAl+3
C2t+1gxjrHxBVArvteEoPm+8J5hoND0evuKVwb3BWLNafJUkEiSh4R781o9E1lVonnmofpHs4yak
QfArCNzV8QY8EQatmKfZINMbZ7iKL6JrJhJ17a9BvBAGj/DbFOj2gX39Hs6QxKlk/Ef80JkILVAG
A2JMuqoA5FHhjhHztSWrbsaKPwLm582I8x2F5FYSSWw+bMm3d7hlc7qGw6U0hiU8ISirTAFumNMn
CfpfWM/oNIgmhwcM5GvPjudxRhCiioLDqj7X9eZDKJJM+gCXympjtkobiP7dXrjWm5poxJc6E60W
tD5aXrg+suf3PF9Q4D9o9HzgSblPEhcO2u/b9V3vp9eS2vqvJ3ICzn3AW2BEAjx6PD+XUGIHq5n0
i62byY9bgIvchKWM1GFlpOd9Rj/lqEMXhYYza/+dL33qqep5/Kyly8KAaWToF9Z8j0ET2jCOXSq1
MWZNItT1hOIKDYnbOMHbqxA1Jonct7LQPMsr73vJga6d1/TfDFgo9cLFgbn/F2DYTLoj1a8SAvpt
Zenuj6gB4Lg5ZUefTJA8v7I28DTGFi8OX37lvauizbR2s2EbDO04EhXxflNGXnJfrvsi2eo019IQ
WWBAr8hzqR+94CgDIwjXxesASvjZvILxdB2yww0KFy0x0EtkEM5A9ubZVDYD/WAsSWjBodUYyVNI
7cE2Ftf0uyJRZ1UcD2Av+D6XaBEyukPl72r0bH0uBNlAhJybtRS8ilyIgrkg86fdSBMRSy+mjZZK
lJXSUDygb5OzgljYjuXt2fFmod7l93CcdlC2PjfrbNGAO9tLERaMD5Zvkpu5tukO1gr38LiY61Wo
eYpU+rjQGNOHTCrQ8WTG2DZG0KNitqwe5F0uMl7IqwHGWSI7lsH0pNxoWA8MtpWPOIhSRowzQGVj
L/iphwPd/7iqt+j7aGm3R43Yo68tIYz3ot3+qrlyZYvnB1tO1G/3E9lbmN14P1PUhXkoLDTbGuWP
hkbZr+yHYOosZZM8s7fwb5qxIKUBw2ce3J2CBlKpPS4r1hZFPWosEZmXs5xxCZrica2l5tVH8HHN
hXQe90VJoaFkPbbSTaZngblI1K6QwdA8WMKwSWT6PS9sbsqolwVA3GMVsjoH31YcInSrvG3cansc
oZYf5+cvVrYEDbfD9dvppAfaPF587BWxXy+WV/0YB92pya0OZr5ov5vJjS19rrM5ApXFXTP7vhW8
/1yEGwsMrcrmeNkVgbEDnq3hzMLcTLYTOZQ7rbtE6kwavj2+92lVXWtqWaguzPA+8Jv4mBBTzPLX
BDO3GTpIVPVMRYbAI1RcMXldRX2sXkoufhEcaC3So/GMZQDe4kULeAK5fDDvyCi1cinGa4xW4RA+
A+C9C61nrAFjW3snlFBslNnYzAccz1lwPGfX9cRdS7Gs1GkBV3JL7YjcAUJnU/LNlkiEmgISVSWk
02XTu+MkPZXuOx8BUrYQs8Dut0aTOfCWkzGZowDNFQ2x+BcB7btCO831sWO2i6TT7GvRLQtIlVyb
a5mhSKmuQluRVjXPPS3qXBlzMlKe9uSQbrS/HOFcdepuPN4vonRd/EBE8Wh1Dz7l9UaCqGvAmPrb
30ZqXkIzqKkmEC2xeEJBedoOlehHX3TrPc8ynqKzXBf84iz2+Sz9Q04QsPpPKelj8LZkjRLWedNK
hHpx+xW1bcQaB9I9X9mw7gFRJWK3mw5kUpwuKz9NIYY6aiKnHaPEgZG6sSouC2WMh/9yoLaTSKvs
eWyoxQwe0AsxHagkbrw7sKLWbuNbjmTnN50tphkSplLU5d9OBxog7m3KJsYKZbdebNv/gGcA8WWE
kj63LzV+sBHCk7MQTgZQB4SpMeCMMDyKxG0heKqeIP1EXKEYBbiwlwfIlwuUkO7e1t6STA1cBdUI
NPgFfe9CZZy2WAzAzmxyfsw9byY7fwARR/x0lotq9uH0j/fj3rSAkEy4SPoMjtoBt8pnLniKWZG8
S6+NfQOOrB8GnMPVM1Za+jUXNT4xMeNTiXQXCEEsOSc1kQXgVl9OLicuxtyTMP7fPChkQqvWQLAQ
YncgJj1PhBxcbsRxUKom70k06RSstDBZVcj9j5uAPxnelRXKrsw73L5InrEHDcBxIOlDaU6kK9/s
zlgMbZDPiqrq4rJF3R8oLB0G5jSxtLMk8mJZ/1sBG6nKQkE3+25OyA47viIdEnkU7kgyMO1OaQpg
OqPw+RdcBlIpxn/hH/PQGyocJVseuU2BmGmPWe/2jmxTCiVhpMAYKhLcusxOQPigfz9eYAzQFblV
mcpBlcqPxGtkK4uWFVzhTfZYvqyOLyQiqwwpoEf31AnJxqxYz+yaJmBuXghINjXX4t26BjUYh/Uh
XcDrCu2m7Z5w8bl2VZ6sxWKsAbTcsi3n+pO3b+aLXnnbeJtbFmh48/nrp4OeznucWBznGvOydIfM
vPTWwD2za3EJD/E9WrtdqQubtK8efJC+hx4caLchtk+Ev0i2CvhGXIP89/OCBYGTthC+x28v6CTx
tTer4rfnsTgKqSJPrjKcXjTywFlDnQqOD/0rPb3tHyatH0Dk7ygXZW9fmL114YiuaKz+xuyRx3iZ
LqMu7k2Y0JZ04nu4TarWQ24Lvyj561HwCCRgqHdKDp4xfttVHsxsSkAywZbeji9VXgp8jPJG2Dr/
ImePSyC/sMkh2umi3Shm8b8LVkOd8nMgaM70NEhKryeMUWFb/0SsqxuqP0sIsdq2eF96/C4oyPFG
2w+l0NqYzfRHoPyDjIHJsi+9bjg8XdSKPbwAI42tkeDOZQmEaJCJHCJgxbS6O5/8OAs+1+nl6An/
BFuxzPSNAbbmK3sPJHZOgE1/mzDsnbHOgJTiGq+1YUKwMGfFE1H5ysXbGTVY4eEEz+SyO3sQiVv2
YXwdsA0bK4KSQspkid8e6myrDTTR6BlaS7CQDijPq9SzeYstQnsVRmbM7pAiXzoCv8E16KnAq8vS
LYHGe0HaKl0GcBMFqCgDT/ApUKRbpaMebr4L57BHwdm8fRFj3xcT/+z1YqwWaj7w9A/RQ/yBO/uL
4oLzjykZ6vFErvnyPrE+gNQbUopAXGpdM5ljJ94AERf/8ijbdiu1z2ua4K84jCYFMzgHI71PyRGk
FN40FK8o92faSyjiAsA6Em/BiZFDHqTd2c5Q2BrFTxwHjB2KZYrHwg01xbOuALagyt1aNYylnx4B
WVzjOlTJ8dpLaey9mi8hDQaEsqEB3HutYeJ4tequZQpJcvI+uYXwnvU856T8YX50VsDZIOEIK1kX
UuzPmL4W6C1EpOfjVnQnmcaXU1hz3SYA16nQEfrzZds8Vc7LY6QIhy/jsaFIRcr5h4YiexlMxcj9
BBHYJUG31yHAMO7t7YRDfZYgEQniH/NerTvRdfrrWpg0UthAg00IZi8efW5qKFI/AU86PvJDGFPX
xnZpCfSjI6qCNlzf0bVh3pJyRflQtgQOB9ZMrgb6VFWK6m0IDeT+ulhNyDx2kcddz1T4JoOMlZ6A
8AdWLC1fnfu3HjxXZM6fiAfFzacddxiiltrMoGJWrGznppCLYpowuOLmkm5lNyDIt7t8gbUPYI8G
pOfJw7zlEyV8rFkaHHo3FymAJr1tBGjSC9V2IK75SKXGCUOetmDCMBMU4NV8qMLVjp2ZTBtzeC3W
2Nd/ZivjiSD/QlNS4Pw4rruIe5NY9jli40hoFkAxaVvfUzpRbI1GRlrpOy7T2WdKMZyIwLg3Fw7F
fwI0rILhHtTXI4YgBHOBxCmq33hekh8ExUavkDicCsQUSh5cTqcf5EVA9f7WF0QfdfL3B3bAfaHY
5hMlkKW8TgqPJBbYjdvFEqFJq/3mmOtxgW9ln3wwgJbsJNP6pQv6f4DzaRjb9UKfGECV5n0RFisi
t+U4+O8ZKF8jGtGBwVr8JP4D0iFrJClHkdFP4m8rFX5ByUJB/m2aRxiLVqhNO3KmN36xTMNtgoEd
i9wRPHTAtQkCb4ovTDoAFKZkZw+k69vvaBJsPA4pkl5X5mxALX4/56HAA11vRTVrgrCMpqGP3b/W
l0Gdl1Y1Diqlv63ypieM0acIUBQtp3BbSbgfSSU+i+c4y8dAmWDcq1qJEe2GN0ktEHQs4lLxpq++
2HwkIwFhgUoWf0wXM3EIC7tgZdqipu86ZwrEtIDXuGfnxfKcT2MQGblFu+7zcdUTpgK+u51CNeyf
TlFWQSfDjlFcJrZHulqMMgwfeJCnROvjga206O7IU/oPB5ucOPfJTlU2T0tfTKDHTYhlY9kXP/Eb
WZkRuRca421Z9amm8AS1Xtknid1HKqHOkD8gm9k/wlpPiTU+1JFD5d91IQbLMEvR8xOQNMibBVeV
JqH9beahAk6JbOnxput3E7U+lilddteg2pa1tGmoZN7yaU5SjimXK9uVgRnSy9Py31ciLnL55AWX
ASUQezJH6WK/zE11b0+snqK5nr5WoixRDWK/EZr78m492m94zL4p+sR4sKOu7v2suujMxQZULEm5
q3Cz17XJqyjFkVLyOVs4BaY44be+aOpyH6qXDQ1CxKDUnWD6sSZ3EFh4qbv2c+vgTVXlrx5TpkR2
oLhcU73ckOEKF6fwwhZuIYNqCItxxlVkUHVSog55i5i9c0Kmpnhiuwkd9ZqW9pohBXep6PP0v1ug
d3gQiJ9y+DA7pGRuoD1eKHmLtEog2Bvu52PD9MsvFMemO2KUchwPmyb6qzbGJimk2CqnU3QjEZmv
1QoRY7yL29pLSwQbxOCyB/Hw8pO58G4LFmOsaN12/Dy18FvaNqLEcJPsCpb2mnubJQlig1tGDYDX
58ZpBg8EoM2DQhQkjulUFBcy+36iRX/poJSjX6BmkBmGx4GCorame3WgirDA5aW7FrlsNcCLFYGv
gSaA/a85AGcA06LZaCrT7jKZD/1bVnYKy0WmXuQzFTuQKqf/gW6k78vt+9gRfpbkaFtr5bAEDJYg
lC3OY2O2W8NAVZpu1ZPoJshCitVWNxdqXtkkccN8eoVCsIdNMIN35rJNs/2k2SsOOcBNs/Ceh83/
/ClTz9LNeTDFB/w1dIw3xUK8blfQ9UzaH7vKmkD5jUrUVoZz4mDPY4MjjuOYAw7snq+LAYLFNZlO
HX84AIzBEJypm/RHnfZzs2ePKJLFabOYBWAqjyxf1jo2jQa7mEvAq5eT+SOQvCjqF7d+bIVLOXOq
ksk9RDcldnaSgfL3QAReFdaRyjAqgW2QE2YK5j9Hi4cOz9zmPBT1yzuIjwhzOp1NSnizG4Q81OdS
MMLwPA69kR4Of1WdiQxOCfcrl8J45XiLosihv3l7CKC8GVgFbqa52zsSLazIsl8JWjX9f8k3RE4i
PJli0TskPwYD1XO9MhwytCSTXuzjSpPM4lCwBdGNlw8Rk54hAdRdQA3EFRpqZIQPHLdIyiYNqLZk
ICaL1DX7kNgBorLserHb+CFVcSMP1Bkk2iXMnRvrTwm5ZD5N1q0V5MslRuO+CnVadRozmbcz2gdH
edDvfuwTMbE/GG9Ux81nFKl1Fu/ba6kXlwyMwhawEs+Qw53RXbm4q4bytOppiHgnlrVwgoKiOoM=
`pragma protect end_protected
