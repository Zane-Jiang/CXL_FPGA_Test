// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
McMR4wmcXoCdo8nqE/86K+7NQkE/xBfv2nR+DMcKY1bWMWog0m0YiXceIXnyqQr9YIsVT0KxvPNC
9tTBfFnqjQloV7nLuDbPWsMfqs01HfFrl+E5gvln095A1NJrMX85beVac7UxvENxz943WC30JZd2
yDZeqeKPGPK2oqRO4C4UI2WgnBe/9h7HwvKmprXCO3FagF4tDR+KYgsa0/YmZo82Dir55V2CUWt6
OSdqB5KF+0HtBfZ0mxn+SOZvF493pk53t8Dh57Nut4pC4864a4yUSiStb2xx9tESE25To3plUQhY
o+HG+6nTtu8+sW9dZ4/jJ/wLbPGADI/HXTZiqw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 25728)
nNPCmixBUkWzH4EuiSgyK32EZU8sc8/DZ6A8ud5WMmq9UqPK0TKpvouMDb2mBLUMegBgRvqc+1dp
BIxzIFvQxJP8/caj7STzX3la4HddAZZQwbVLxe7d8l8uWwHB1pAaQAUbAY0UeUVSGMd78V1a5wyI
TSPkOeZ3QljC8DxqfmaDaBc8sOYgWV0yTo0o7MtuCEn7Y3TdFpmHE2m/0vQaq8Vuxl51VkMgVOcz
rMTeJVk+3XvcxHzRSZ0EsUI6ANZAdpg4dROyVuHPeCGrn965M0lO7kAsbmqxmjsoY704PsGMav1Q
iyd79082D6/c0qqnMpK4WE4+u/oTc2hLdEql91CbOGN7zUyA45+ipBLDuwczjtUS8nV6iSgTYQhw
W7CiS6h0pxA2B0dGpUlTrd8PP6MrIiBjw5PndrBuUb4Zh8TaANUrfUS/0Cu2pii0DTXdY8lTQ6Uy
Q9zB6a1kfRQ5PqrllfkpoELZO6BACuHx6twpwWzUQJOKsRwPWkRtCRm5Cx0qPJhoMKC8O8jloz8o
npEA7UxQmRNmOdNTI3NP9Xw+lgI6/dGep5EM5tgeoyABIkjen6Zv3Q+iJjuPjB1kPI83wmC152Oq
Nm19Qg96isR/ivEA2yUPwU0JC7XGwtVSj95cwj7wtUWvHAkh8Yh7MtQML7YX5gleUJ50sKqf36ZH
HX6N4j10y7YUE+apne8dmXNdSZ5IUIsiiZhBZnbqn4t/dVlV9T2ssLFL8gRyhqI5qmRzwq+Ok5KA
NFkA/EMTa4icM3RXIXuXloJGh8+251u7hw3+655krOx6L4tSXP4ZrMrujy+GijsoTh3iuxqKz2R6
XOxjlBYypo+mv5l82z5nLu1enp2Ie4NDxuBrPu+RUnOtpZYc42mcuArFpv1978bHca/8uqVAEO44
jfpRsvvl1ph4VGFqeHHAbrxs9kjlRzxjXeEd8gQVCLkr3LVtrv2APQT2uZ5MrI6o1hpYmD6LjprW
lvBuFQ5QWlr/YmoGSSfxWg2i96CVX7P4F/TPI7l6SY6xL1raOFG809ABSS1f7/K+2AcH+wIsl741
+rCuN6bzMJhBXSPGF3xNVXir3oXpxWPzWKgei5+1nCygx1nual5xj1CCigdJqJVwE/YCQV1KUG7f
3wh9D3kN+0QvIKlUueb2fbZYZZWgBfaACA4nex4u1dOInQ0Eum4W+F01eejdBpl/DynMBhkKcHpZ
7PgQ1kSkT8wv7L0nk3KVpHs0OZSUj9APym8hIZ+rmSMFREAYe4YuzGKXvYI3QraUccproG3COgyQ
bcISLEcIoythsxm1PPG2Rws0/ypxZQoH/JphDlUmeqSgVMQmsJtXdkc6iOuc1Ts9XBXYv3pAqfoD
mCrXYwXBG8zzt9A5fexZbA9357to5NDl5m/clhddyyNi2h0b3iC6ZNCeU5c16+YMTRpChGmAx2CP
9b05087mbWIp2UpmZ+UP+tyJnjokkUvRj8ictPv+4on9FA29IspF5LJG+J1aBI3WRF8SZ6HmZHW7
vc8dsdPrRwLpibLHLDtSAXcaMUPiGVClte5spOFw2xUBt7dg/hco1vTxmL5b7+kTSGf1DkDRq7be
7fbAdVRoh0yTfSqOyQXmgRjjzUbhM2jqSzQ1TVvFfcLRFxo38ldGsT3m4mxcPDet2tMuzenoNuez
k0FAhi98DcWNmoeNKdvT32EtnXIMVy7D6SVJZH55LHkhz0kuVeA1oKpM6jNBP4w2pobaE2KQQLCR
vSXpztlc7Jz1JS1Ukrtl66WnutBcnGZ0eKfwWg9Uzg0kcywtAPGwGQDHoRMdpBGHtnjwIfdVr36T
M57oxQ7v1uCVu/nu8pn34aAEIZfIWR6xcy5VMLbhckzaS7UU+0yeSJxV3aJY2TobIoGVTdUXVGDi
GHFerLcQAQARCRMHsrO8wV5xKMLvSjTaAz0MzsgCjwqtxFgq963UIRHESMlQJO2NFCcGfPeggskR
39s/0jDUv472KmWXEU/UqRb1kUP/B/nIc/6LTVVzFFfPEZEmCquJHIHEmmRJZH7xz2ZISRhLpp7Q
LjEPNYTVvBK98cSP9iuBg4zOXyNbp/ZvaKgPjsRtbMRHrpsopCcMFpmE813aQuGvR/S0fGUiqpTT
DQ0uYusVgqpseLHSjzm6K3cmsz8h1h/eF1dOfyZB2xCDifXqRNRFHbIs3f+BuQDv4yeAI0Bn4hxT
wGQIY5mqF4ig7PxmHIinkI/Sa5wG1uBrsV5NKhsAdpY7cjBXcpJD5UjIMJxYN9HWhw6pq7RFOyu8
3+J1F2DnTGnpKWQo9fxI230My7KUhBbE0xVQD4T4uqoMscpuznoFDJ6fk6XpsvIBZmbMAOC8sAFy
no37M+gKoIcPf3jbaayeFgP0OcwGra2Tv5GHb/GMhIGCW9Kfdi3LFw30n9vt0LoEv6ycoCyw70Ab
YaqS9Y6OHtzGxTf68+7ome/SzW8SV2rUl1ZGlx5sMn5gaPewsJ25QYf7LCzhQ7E+LClk43V78A/q
XLtQIwvsIjjvfH5VG/NJo8+1CGmiibjsnaZv/Fo6yX9vmCIyRXc6TMHkiQiairNYKoyQPdWXFrvf
5H8FnPAX1x7R05xWq7Wup35EN5tDOsOosV5b7TP3lVAdvCtM1SWMPtz/ObDT7qiiZmp5ORD9LYm7
Dzw9ogyxRPEflHe6nX0PtkETuPD3snw9uc4fFXIcJXzYvSXIfbmR5Q0DUIYwc03CJQrGQbxxLKGK
/sg2Cl06cqqMHyryg5TpEmcHBMOSLRQoeUvUH5uDoRIOSR5ZZbJpClR0vPtvxkNjMhyTBi7vI2II
+m94Kne30mflS4bhFZwzAeMWTJT+kNqWApX4CE5ULsE8wv3t3gbOQ5dL1RTVVmcMqqff5yUumWIt
CBkqFLs7NNsyp/5tRwlA2oEbHTh23yqPnBGhs6tZMHzrKTE4s1dB5tOaz6Sl6Rxlo/XLKpYbtiQv
nX/E+i5lFeqzKl2Y9XHN8yvx0IbBjP+AT7n6wgx/aNz9KyweT6NlkRLGnJ4QjcIHkFnuhMeBhrXm
EVK8nIqueBr9kK3HYSs/wIlAZPKI0Tsp9jIoeE1V++DxUpXreKINJJ2utCXWXLYnXxx5lK2x/xXJ
XqSSbiE2oajWS5lEAfqbUBDUS9uWU/1OGCwR3MgJ6zMHhM4CPmTSFHDleSzuWl7N5KS7ySTYklwH
H9+lAlH3X9WnncWaJua7JME4O+qZhf7f8u2Rdv0CYyGpH2ZYELP2JkI6diVXK2gUoAKo8GdVUX6S
HfbQSpMNJ6qdg/xsjR1AQhrXFaha/wRE8qQuQ6bizHC44IyTpUdN1nZUzJG4VfJrs9UXdCMokqqj
ySEZc4aIh+a3KEXeDtN57E27YaN77L76LoQL2gMAvYR0X6PxD/q13V39nzIMFcqoFVQ7TgbiQ/sq
sxw4BI/tcl0nbvNS+LXvcyZDJ5B8yyFvXhRUflf21Xt5QTUvjsoBimg/2UBrpL7BwyxbXrCS3vgz
hxMpntMHzpJH57LpX1RxY9Qr/1T6lvIUgipQz4/MdafOHMjSC+ftmUlLm008S/F2RfwgE29s/uJl
sqhA4VXYhFYgB0fhef4v96PaXeXCBCp7jB9P9G9WJ8la2Y7VaV+2pekO8Sa7njaKHeBY7oNT8MCY
iy3bsLaOwmPPPfblAPmLxLD683TJQpN/4VHgh3k06tptMbINw7TFZdWw9VF5kUYn/F/pBBcepw2j
FgvPoQ2eBG6w9Wy6Pp96xwbJ5snbmAte/sjV1QxV9mILmijVKp/y1fdm9etY7NbjEltk7v9iSYuX
ynOe+m3WnzWH4y08OBmOShgb2jI+GqeBRX+3BLjSN6lW5Y1ZaD3mQcpg0gTUoRbvIXZBoW2vOBFR
PCTScQymUQ8Q99gSg78uwD/3tiXbFphNAlk3YQArYnR8mC0tjMAJPTRiYoiT4YdKIOemkfXpjB8y
WQpjMxgIPOqQJjX9d4Ng1/NfgH7TYkSXra9PnCwepE2SqpZD8tPlfelGW3NUVcRlsULlvDbALeys
q0v0HtBfe7aVJgWlqYHQTXgJF51IhTNrR9d0wJ833PRGMwz0R7Gonml+35DnCHwHOY92tHmt1XwR
JxDa8cGf+QVCB2v726qwrBrWXa0j2XauG+FW6w23+8uEXBPSUo1ZDaCQExxuyS5dp1co3W3c79UL
foAnV4E9eFaotCOeqJBfBlukDqv2c8lysncO0ZgzHqwqHlHcpu5rI1AVoZDoa55z55nTDC0RbnlF
56GnUngUecRs4kjd/pkdHkhcuD+sMI6b9hwINud6VgGq2z7PTkDePpy74VQZFu4XWvlOBUe0dKff
lyMt4oYXuZL66W27jELo/Hrxxi6189hyNZeRjiNS66txlcHJbbotmIlSv3q8U7AuDad+DZOu1dyf
T5+GeR7up/d3KWEK7qhpN+wNwpktzeCh/q2IciGr6WTRufzUFGOgOPdbYvA+PC7KKgAIxoMTDw+C
KfVrRF0ejph5csyV0e2rgRUHt9EXJcQXnUYiwPQfN+5/LWJH87SMkqM5XdXRGHgxuBGxtyU4pMmA
AeZX0s3D2ugYp2VxuK+vejN32WYNO7sbxuFbLO+F+HcjRvfBm/P9PlmRfh+0WPJDN40H9FIfqnFY
ZxEDMLOX+VnmmLfJ6EKwdgaA0T5f/bmxhxakzlnocx0eYDqEeO5AqilRqHIDKNCsOGiIPL7T6B3n
YDXEv+nUcJNLC2Mln/oC9kHpCQ1LyL4UCnagI8GlHSnNQPxvZ5MTPw31Q/hu3CwTfqjMaTOET5yS
Bo7UmDzWbw/HJxPF4DoGnD0m3NG7hHGOz+mtUPQjcKjlUZ3TDjtUtRXs63bmq4qI4YYD5/7bmfAL
YZj3uUjvuy2r0hM03BLyRZ822+op+IXyll4gYQhLgCZnZ7ViSQWT8ctAQpIWxWwmviefyt5ajz5P
FlRhwshTOJs7q4Ah525/nPDuOUbWVF1GUSRIK3kn9PeIu6dvwQKh0qinbhDRd0c/+YSrGWcS2Dt7
Fq6QpeYSNLfJ9DlQn8IvpVJvMnqWk6YtXhVoWV4Sil9EQZzVLlGnhnXp8KCI3ouT6kHf0z1zjY/B
yRVeydzDGkC62Jw4Rt33teHwD0GHUMyibrHhBp7outnQBNOKpy+6PFxml72I6MjFCH1cgY3BHdBR
gl7qDt+j2GEhvrOOr4G/r9+NYAR5pqz9BI9ZZ572Hc0MO/XO/6VKkTdXueh7cEFEmUqZ/HKFAknq
4Qdw10UEgCbPtqi3sJnd1I3DUIyWKpPy3x/isAPfJSgrnNy2NCX8I6Pp112TK+HPKdh0T7POZ7I6
IVXIQPQ9ACHeFnUeQXKzY4s/9PP6DCa1U3VwmXVJ1iKRZb/VbsvC8T1Y770JuANtSeE96UobkmJA
613YC6XOVjsNqwou4ruOwilwcSv2fPNWKZYcVNBFctoAD4N/urBeMNmY4wu+dJ8Z5ag2lut5Uord
j0qV50uMTbtOO+cxhe+PImF622bF8WiJCeUPv/ekZ/1M4ihx3aIuftYdQRb2b0fqvjhtpCOPC4SB
X7okJK8pTD3WyCDtW1EcxlRt8+WHkzf0tu0AqeFKCVtSmK9HK2waHEXW3mkJSzfG/lYIrGHfPcFC
bQKu9uqHWZTVEYUlsXaOSPE3H1BdFLxsYsiGn+VDXO/CHdIh1narRpukM2u063qPHy/JdcftedZt
Lb+qU7mgnMX5Kq/n4XSibEH6G52RzxiFqed2pCTsWI3CJwaBvMkmAbuJTI4Y5z4RxftGOLrIKhlA
1SatBmKyP10uB8P5YcRTdXCH/kQNCcXq7EKy0u3PiimYDlA1SA0o+8wRGB/Ieb0krYq1Pnl/tY0F
qtgATHwUJvkT65pHd/WJ74len23LhJn3xWn4DOgSMxNhLnCfPpjVdVj/z1wpm8S+vH4NYXZwb2iI
vQesrZvF/oMkEhLS20mz8AMqxouueq2Z+8ESInSsq/QpfY9fhYfk8RzIJ/sLKLVG/bBhGF6mlq8T
dG4vMw4Nhu5acI9LgjLLqBnjuVN63G4cElAI8njXZoIQ9BBDPoNGRq7j21l4Yw/k2buDX3zTp85z
FxX0l0QET81SM6MNtaoEejWbk+qRu5g0i8K+eCJ+jnqST7tUJkGfu/A271aYogzYe32BXmJdahrm
yLVwrkhWVvpceZMJ25R+LudIoC2Z1sH+pHrIrFTwW0lrR6hRhMR59lhFUpBNRAXhYpzO0hUHGiOJ
yqXG4LDOPqMgvZj7j0AxHhb6pkk9fjHtBUaUFQk6BO4QjO2mFeHnZiz9zGYI9ClJTd2bEQ/S1DaU
76BriHNedBHu7qNvquPwFxdw6F9LfaWTgR8mwy25SgNTUl4KwTcERjTWoIAnMBNNOLLp0gfQ+AlR
p++Mfsl0oNhD7bdz9ucZ6EwUMJBKuCC6pO/2M/KAA54JfoB0OBo2cFO2u/zgNg25jXhZ4w/d+uLf
syaEHvzjuEJo414H2vU/K6m4+VtkcsCz47sDZs80sjQB7CCosuBqBPHRUw2hJpFv96ZRpZU005/b
G9yNwNPUXmjWZ1i3SIS0I7dh2ndIVBalbI0VHYe9XS28/O6cWrApmzJRNepWq35c6RZQa3/PkZuN
J+B+Q5eD6CtLyuil8rxPQsPRz/A88ywYiW/27fcnTjIFYRfFxrN4uMwUz7nF15sfsMy8ma70DpfV
qazuiajXBiLaroac7s4IM4tVx8bnzvwfUEf0OiLikzL9FNc0K/Jtetusww+sjTx+G3dwoXhNvMDi
w6g2BgAx79jxHzneLlAsTinRT4oLKPnEnlufvyu0I+ZOu3MJjvq5gLSg4wKL2pQcJuFMzXa2h+03
2yhf4pQWAjNP1H6O0eHL7JC5qILVUbkaAxpthpVWzEo+C9V5Du3h03DYju4po+CRSwfmspoM9piE
+mvt+cfoCvPqG0T7bYd+Uhjd1YX4hxvg23bLi8VW6QpyTe+SCoowdgDI4TQp6kb8KvELG9SkNR9j
emEvqrW1/FHl0ZVw5PW3UaS/gCJaPkQMJKepw5aYdaLxdRhE6SIyeXMF0k2fARMiSHFdTD83+9i8
f+bwd2Kp9gbJ7K5EoUPicutiQt2ifBQv6S7d2KTMiG3R3WPN0E4hsUpMeryfB3iGUrk9D+isZr8U
Kp7yHmAkwEtvsuXMf+VShZXU93bDs+s865HOZT4ulMZ2XvIh65k6qjV8RxA9MTa8uTptkx53EQ7P
cdprUfvBZP0gcchNy6lLtyEQnXITP/F57MAfK+78NGW8IgATt6xQ7nZf4zRTaay5Aatca63vY7sm
crynPKG7jAC00sdnTX+cRvZ8nikqtv3zkeQ+0bUCNn20OYiVI14H0713bDGn9HwW+MxVou/x3UKR
LDLxXNwX8lXUHEN29lfLkYs7FRrXQ7a2xZz2MjQkXQxZoesDYUwVQd4qIGN6gW4ZZsUZrqxSmtJk
wAnaP2uhTbwHQmX5UyLs6HnsCs6qF6fWgRmWRIHUCT/6rn/NwIgAwxcVo4ychyGXlwbGoaTq4JVf
91ryWPrJ9wIdmmTzMDWh+8ECUO+etCDUJEithjzpKFD0pYbYERFpixdrw8eCK5kQ4wdMo+heldna
59IkjPxce33Bb5CffyRxLFAKT+pm41Anhyx9c99e/mEnV7NoTU2AiMjp0QBWS7Lw6w30TD8Q3umO
FHYqNX+HSHuvwtHo6wD0JMypJssFgaapNbgyTHtOZKqqTG7cdkfmCt7Sju4PDt7ZlYajZ1GI9wIS
GesO8dNRwK7rzaj+m9e4NIPJXcYFiszYRhNZKHNJ2nlvmm8BXxvCxKDmmKUBxjRgyjD24n4CjAVd
Iom5UTNhBWu52ySWZUKOajdKooSQcPVR8avXAgmJvYraG6DTsScfyHAF3xmVC8S0cixzDDKX3djG
RmX3gvYaqBTr2o/244hZZsY/da26rGdzfSZuVmNXd5QRPoo6UT11P7DEFH2bWIVVzC4ZFpD+wo8s
kMErxpnBRwHliNd4WYcNkk3tklB7s/dQ88ZPBeXW5ApemrhKz4WlKah1DToso3wsdZs+M+xaWWQk
Ujpo03xOifbgEuLb7CcO2/NLfXqFkNI8OUuRXr6K1Ms+QHEm8B4mHnuxNwzhMdTOKA52P9bi0amy
9qCB8pJnVBRkXQmdE3yK2yyy4e/ZN7v71JHaTFvtaBAVqogLZ1bAFK5FcgL0+yqwaOCVB4ozIDhF
BuzNxsYcICmlQfSgtMzFeCGohNWiVk4krcmOpGGHJv+ikI3VoxpSLfswYkuUzMHj9k5IfEEAtjHN
PVbREZyU6hjZzzT3ilT9aTf5IIQxpTvL0YiBVf8C+zkRtt9rpvK0yIUZM5kitBEf17iertEs51t1
shqwYT66k5mRVd+t/QoRlak/9v6ovJ/aAaZoyfyaWHEv/dNRJUcxQZDnOHB0MGlc91Gz53O4NpuT
c1LefdOKIZ6yfqjOA6Rkp0cUzwYGkhDOPGk6r//f9RLqvEBXRix0maPRzPBlRZUGpofkq2+wJCPT
HgcnTe+qigL9+Qr1MXukVD7gnRYMsUUP+MARBHa+9gpDwJVXzQGs+NX9CxFwbyobAg2cNlXbS2Az
G5er6vVmeX/33PGvMfqlN8b6AJZbRow5Nrt1wrJJkbRlRaiKYQUxz0byU4fGoucqn2fY/9zaxnBK
xgFv3VkX2A6gZb0pEyvNovV2gTrDRtKFIrFlF0j0+WFfgdnvB/ll2wRXzKxczFpNuhLFnBH1peul
mRb2VpmPPLSuvGh8ZrkMzaPGJipgNv9bc8zlGyaKFfEseG8LAcFPQ7xK1LsrrZNIAdWp25iop+8X
QqF76Qrc/GoO7d9GxbrT0SKKl/KKtVHUtQh2QZbwoaMWWFKJAc8wAA9yTdleFzT+zUus/3gMlU0B
yBwKaRAG3UkW9/BcYNgEt/M5qD8T+uL2vvW33aRUu2OxrxWGoDu4LvXrFXc8EoJ5yD5gmd1nhXCL
vrij4euiFgGogIgjs/GnxY/t2p2dVcvRtG3cRqooBKGchXlQHIcBGIn+8R7NSWLEmvqbVYqxSLcW
dSLOiaIL7pFgegZxD/LS0NK+hKHWDRIMhMJg7gqxhGkIJfok1vE81fhMW1hy5Xl0sNyAI5KAHSO+
bJyV/y+KMonezJYCRh3bEPnktKff2a3KlbJPd7N/6IiG67Uf1eWL1RmAhPyUrIaqDj82Yg5Xwb3F
BaAJB4dLD4Bg0jQi6MY3w+4JDqb0APpIcvKUfUSLqOfr4L4+1BhO/icMMmTpKF0sXO9v8Sx/qk2y
WqDt4desXd/oSecAHoF14thXkL+tqndbWiN2I/A0sLxe6ubTn4CknYPnPFlrbro66wEnNWkd4ht2
L/UWwOitsPuMT6lM9lWLqkSDTiHHjORLlhPpE6kCXiWBkNsEuVrlpH+MusUK7ZC203lnmI0K+6CY
BVKXhmplcWYK3cuni1amnqnwDke95zhJZR97pjNrvTBMPa2A/uHsunzO/lSCsUEiuwK6W1YU7LoK
7gHaiptVRC42cdOgei+YkIIPCOS4Z03LughIU1Wi19VCCmYsQKlROC7WxMBac1JXyA2vjIFgWLdE
bRsMinNZZl5O5EnQxzk0MYoqB3S8AsHRH9xY6d9kizDX3Qg0H1u5Jw5lF6fjK0D4DCyLLr5OtGZe
zA7c6owZVk84GbYc5Min7N7VDnlKSRvSa4vMAl6J7BH9lOZFw3/vF1NnBZO1NB6S/N8IjrlhZ6Gj
gpbAmBSw9rbREfhHUZwscmQb3l2YpuE2FEt+bPAgWQdyt7NdZaS/THAd9JARFqFFnVutYBVKfvou
LaUkW7gvvxArdQcqAL3RKcKtS3ZlQMOiWXrXc/fBQBgcHpOF74yPn/eXML2rqIgx6/4hAfJDk/s1
iBbm/vcMBZ30gLPInSaAwesx6R0/781juYMKzjD4Qr27W7/yecghCX4uSK/LlD0EKaE+NSYONQ2a
Y+m7RjhDYC+KVv8MWMnOvfoqiHaHizYAioTo8+fwTJ5k5BpBZ/gyvjjTnh26YqIqxBMQPk9gjN7X
rMZwxzTaVupuFV81yZsFsOVBcPYySSXlrzAjPKL4EjIAIU/p08Xr9uZLSbNLn2IMc2HkuznCl4fY
q9nK+5m4svzZUmHAsnQRbyiQprvWJQlqHdtQiGLEz4Tpt4bmL8k6O/ztm9lTa6HmX7+LqQ8zPZuA
J2G8gCCsSQJ3GZGAE+yUrGtQt0SBYaE8EI6Uu9IqSR+VEPgSOpL/qv3g0tmhoc/dM0gfIRTd9oGf
GRperoPnoicGtuLzx4Qvi4+8mbgNI3Onyqvq14UYCNoawSLhMldlmRZQMs7DyAqaBP0gpJElvkVv
Nfb+T4M1Lw2TzzuRHBkBHD9eCmiExTI+yZN3CV5VcRo2o4QTlMS0TyrvrF0LPPIxwTWd5lp9E8xu
KPSA+hnmQ+xie0+qTHa17n/YuWAftVlFS7tkVrfCbAJ9PF5bof6eRTP2YQzIE51cb/hYtuSFpwkJ
F4xOeW9SJcVUjnAZbndv3HmtWPSoHI6gNBtrLt4o6fBEsSelby3c32rl/p+qNno4LkV9rAP5UQv+
vhemPMfKhEUHqB0VmceE+2ASdZDb9wI6/Zs3j8of5bbD7TjNYj05pbkUB1TrcJRtwLFNOPgwmPjg
ne0kcWWDKfaKaE/G9FkIGRaseCDhqzeeMvAHBIXK+lcfLVVCK0orkTEf4UTzGmfrAZFPuShzcLZ8
/T4ADpcNBnKMPhP5DauZR+ddXteQ6+eM+upg8XG1K3AkY14Cx+R41EqO45DoVrdsOQKbYcDktB4g
AkKu0Fm3VDW9+p8s30oJ+zBWWa6dZb8Es2cvgLLQ0BY7i0IewW0EbjyuC/Mj7cyd0kFGf1ItMPsj
2N0X9OVEvhMmMldYkEV7RBsNr+hXiPcBrscwh1apdekz9apoXlow6MgcfMpC7/wUpz+oP7x29nyo
l0nfyA5FRfgQE/yqGPCwGtt+vXDWI0NsBEAX+6/EW1fOYrPEDSMiyKUSQ+/4PEvvsta4BnZWQ8r1
Ji7Y9bWBgRzSmG6IDME/K4kpVadRMkZp/OnXrKTL3roAGW6zRuEI9xwQ7uGtLQ51SztXpdbe9rRs
GOIU9LFIMIKDNC5PoQ/CsToZY1wWUHF21mf3A/NxUUf0xLZ8ln0AfiJa2tuzhazM3Ztfd9WAekoP
wuenqa3rr86IZOvfl7dBt5vnjVuD22ena9hstdfSQX4xqaUhp09XbBMDgGIMb0y7l/lx+FZZIcSy
a14JojoQmUOi9AXzdGtSGilDLZYYCOxSFQFsLpHBDPMzdjE8HC6qxnq7XeO5V8txEbYvP0r4Zqkz
djU9nlOEiyUh+Rc0medy+6c3u6n2at4z8KmUDSV5nbXDTh7sh5kVizKjU/Jdt9j5lIlA3+mBzsTi
Btw/R6Ycu8Jssxpy9j20uz4ZzbxM1Ml0YIl3kgXZZZwVNWF+cpgGEp3mhfUdnu6gAkLgZwLjHnUP
BnTCFrQNjOmCxokt9x7zSmghpLgKA2tQzibx8yXQvNDKOmF8+VSIcU4TTCnWp/LR1XwVw9LhVT8i
8Guvbjz1zP2meYrdz/mrwoq6j3hYfj1nERp2lAl6ns3g6rSGFIKyh+s/HZBnGkwl/BV1bk9G7zn5
hOeX/eZODYLqFi0k4UpVXlYvvNUIzLCwWU2DqHFXqQ7PkMT5D+tyoZCp0syOcYWylTr1i+IWfj3f
Xv0cxvaMaRmlY1LXb0xYNWzVum2C8B4JK/dHa3KCIITz2HyVwXtaGsTNQsCCx5YcGmTg61Xt1ZNE
QtxGvv0CYgftMLjeOGeOloBqB+fpXrt3EqMRascu8hQihN+sKfAy+VIPDySUnLPRO3J5hlaZty2V
y0ffmUtVtywp3ovvbY7HrlFvE/J44HnmHQLCwwc2WwgFdYErJms7dF/deE8SoCeYQ97TpEk6A4O+
qZH7eFD6DAfTwyuzWBEIbxjp2/1Albxa1haeiCXfmUP0WnxVWFlzx6DCjOnmwmyhbW7E+YFI6kXV
9vbjRf3+nu4/ys0o5Gpsdj59YEG2dvwbDdNcwmuMJHOGKYvHwfX85Qo911gyVT8Nq5BwpzbJ3bL8
XJw+qJXfy9eV35yekkRhgtnhWOGN2JSnRWYtKb7acdPjeOmAzb3rkzDF0ERbgrU6YuoeYNmgA32s
lIBrN0kKfLvSknJDAdeRgqADq8Ok1w4xgCJS15+KfcRsGQs4F4Vl8iklV03wBMcH9F3lbMxKL0mH
pkwccD7yAylnGfM/AlGAb25lHo/DGTQcrcaDtzed80ScH94O3Mb27TMrPw9MuFiL7iBrH8Xqiw2H
6HaC0QoA3Zpeei6e6ivuqCuKFuxcqmCTXOWnQaqgdAMeovaNnWAHjR/tgM04fMUBfvtFTt7ZRv8A
Vsx64jxgc3Ph+ddt4f+dRh5MRCODWvyXHTN7c4uw7HA4BeFGjim8gUE/jm1jvdGu4bAfaSrDYqre
1073Wo5udTILIvduFyhg23yuZXG9lK6evQqJztjA+OuVqzn/4zz9wmPbaSX1gphmnHjux8IVl0ZN
yapcwpV6s6sonOpEa/wap5bQap0zt4ydp269qVGFv1k6iqxKld1OOYNDxyv0ZRIBoGGfQowMdpHA
XQWUy23RszQzUurhrg9mq1LFSlMqQC6GfUCAlqZBRRHXJX6zLSyIKjB3nU2gX7sYIdJ4L4ONykzJ
oyKEhOdV1PcavvgTpbAcskhRaj01N2OzVtzqt5vnRzFXof071Re5RORBknu4ebPETmEdrtMy+qCf
ir8OzVifq9YZa6kgnllkRlWw5wJw8g+3swYpvSImwMBQe3I6jlfXYOxLUTW1WHxCoPNn5PJHuoXx
8YtAWKW1fkJs0X3XiHNYw6f4pUSb2B25tOUk9fCdYoDgZlRKqD/NNnMx91ACZ2mhS0FhIiJwZURi
7LajWIOuNbxcR6PeM1fiSzl1KGTrtfAfOQmXPbseAIRSvbJsqpZfrGBv3+oPZiAp1aJht8bh28hO
u+a6E3IEgSnosfHjP5cxw6rouyW+zYfyxUETtp3aT0gu1bLZfume1zFZK/CnzNdKPUTp71Ei1S/o
eZRNf5BOmlvZ9PMtqKNmRHoBw+bm5zNbxwmelV/rd1IR2XrPodqTOkHZEz2IX4PBtmEe9X+B1Epd
LaLvobpgiOxZDHjZ1QCGIynh6vj+bbkg8iC7dFold/L7olo79TrlgkxQLR6z/aPZ3CZuudg23gLg
FV7SVvMJVsBSp+LH00Y2VC9mVjlL+vyojCe0K1pVe24LCAzFTBd2xYNlsJBXrA9WEoU4owTY81KZ
TK1ORiHIQk83+GkMCl1w7O6ms+R2Ve9AZM9zcyHyb57FV2o0Sy9u8HXDvUDexwpokX5AZPVETI/T
KN5gcfkYREx+QbVs8+jkHcH30JUlbDAaedTW/WrSjZ09ixZg5Dpashy5n9LCANqZQN9UrDFh8SMt
mV8aGAeA6eW8JNy28qtSELfCI1fz/XzhX9I7RANsCuKqqv3vuXiYc2zLGW/ObaBpsjm244VoYZCz
9kgCZY/mrxfIspHrjk8kNBFZ395762uF6NlitvIHn0lA8pcTj4YVW2LL/8jFcVBN7vp0fsF/+OOb
qfAUdH5B2DtVbpvlQDHrEZM3jKRxHBrAzNIK6IxxHoGoCsk8R9rSCrPh5yHNf2XkGFbW/6jPv/E7
ckibWqzaDSqAGlaUUfVtqg9V416jwYB6PqEDgNkyrsKZEwDMMZi35BIqe9qwb4fENywDjvzq+tNJ
cIFR7md/thrOF8DRXSahPoEAE/VT5u1Lc+DIqvLh/gNxcGmPFytaLDcS4gvU6+lgHGobrv/uFtwl
8uC6TCjuNQV7yTkoO6o2N+KPmBnhMxBugH+3yH+xCRCMM5pvva4Px7HDDB5zrvcDwy4OdC2+eFBw
m/BPanJ47kyoIYH3VPG4oM6bivSaAax+vnkwbGaqUo+0TvB/C4gGiTBCGIsNu3BqdhQYhvwKMhu3
XHzbRs6s9/w5y8k9EEitGxXRdxp8VJIIHnqrI1QXB6fW3QvXUWSg3Xq83iJqW4f2ZXDEMUAqtFBx
pwLNgV2zJyZ/rbkdnBrNL2CbY3TiAcMUQQ2q9p7UH6hBRp8D8u0AGOwalCOrBEnKv8xPfkPLvl0u
mIaiWg+Hb3bHQexuz40NLbxY+G1zXcrDHNFyDqwzHrR5K0PSB1J/O+MgVizycBuzSstUD1g5gFVi
TClnw4WfhY0JqJ5onTC034D0fPNtMwA/TpzLWZyZmmNoVSrmOhPHpe910WaQNitpMvx+oIXezK6L
q54Hiv7/beLm2xppaiWK0XqPjVLM6sgvO77ftTnbmxaIP1PUEcmeEDHAt03nRYb9kZ9pOeDnvgga
IG62iohhUrYuJbrRZ2anGzidZ1OS39dtpvvchRdoX5TGOGuLml4SSaewAkubDC8YOPOdbrRVGpvK
9rnljCSJJF7Y1orPHNc2gpVTeEjSTYTqeYykUvXZzuUXWVyrucT1dFPTdKZa8tqj6OIuozw303Dk
WB2ZwHQoWuoN0XT7xh/AoIkv0iGB7b+wPWPrDvX7Ckafd6xSXYmTEAdBvSqSoZxMigCAMV7gES+t
dCeZlbZWwK6D8yzhFU1C4t55s2OL5dj30Kv2Z77uUqkOKyVPaZriCcWdDNOiKtE1mdMhWwANfvdV
PTfrENsFNfe++l7cLutcJ3I/Hih/a6WvHirN1orQ0xGCsXLhbKnn7o4Bo3CnmluY/mH2hs7+/XdT
sHnNPNcXRUv3Nu6z47e8HYjFIaM6YZaTw55EpdMpkb8WxWOz5LHkkyJug3MDCy24HJMnrW2fYqK6
DQXFJCA+CUiBKBslua/5jrPng/QmD6RXZ0EclYVlf+kvTrRaSuZb6PwsCdgvFOJXVRDnTePnUDTV
XT17bjldpQUMn6j9FlJYJXXIkhG4DLBZyRhFzEBQ7SJQSvRU+hIF2O626k8+sxob8HiyvWWZxgh+
Rl3cMa+aXaa38FC7dWd5SvA7pX/ngCI5oYI+zX8OtHWeOcq70AoBjZ51XLmykdlpMTw5RwC8lEMi
RnN8Ts6bDjgHGNAcSlBEMvDF4tlQgVal/8+eRVVJDCK1jjKIU2vK4iupji18FiCMIn3o1yCR8APl
WB3fl+2xOUzAm31tg21xtXkjWoysIOtDazSu4k24zezNjyXY9F+Ruw7Ovnk6mii0Jq6nYFb8kQG9
0u6bOC8V+P6POWVaP2khYKL8EmGfzwHgyr8TV/4vzjDaAXUiA66Dqb9mZlHST/6a6JiBJb+h0DLi
xxal5VdDZR6vek96PGb5BXCZgt3tEbhjEvMF5xBnSHAPwlCOTBor2RBuo2/uLCniHd+JxehkjEu7
OtIEuVPkniSDNQFsRKG4L9mddz1UuqDHhvFaDBSJzdUihfptgNekz5PRiWGdqLcWbeGe/ecwNmos
n5MwaQDpx8FZdg31p1mFFDpnqgvIdAjnYacAtR170wAoHxJVirHp0QLipUy5gKKytH7P4skGocUm
Pyi2Sri6/kQs4A7yvajaleW9gbCeisalOgxMoWKUW34DJvx4nDQ8iA5SSRYX4lU0GgeXIgNtDTEr
Sk8mii+na21eoWLzjd4YALS7Nzw60mhrLTSN/h6HQXsqLydVw83qLU4haBk0YzFXt2w63K8nO/Yj
Bcs8OGDby+f+lv1k8U6d0DcqTTuzcmBIiTTVMetIDbhd7M61o3x593Dg3qX3jC6b7vuWXgaNEI++
DlZfr6U+uV6OVu5GIsVJKuVstz9bM+1kwC9qoetvc7iHwm1fIo6M32iqt7gWCWHehhTdteXrmhqq
BV5UmIZfPl43klSMmVeUlcUHK09G1TWPmqBOV7kmCKShzdgQVe0LSgKtg53EpPYmdLeRqeS1o9BE
1oRZXVD9ItOg+VMapr32aHFcZ4CW8FEPhq6bOnyAbXnLT5amo6RWDrEfVFdunxte5vB82iC0Z39c
Zzm2U9GvZB0mPcwBP07lmWSXhVjvuc5f7CfFIN0xymIy8/MjRMJrz/hdEPRV8cFSlDX07VZVhfdb
rGpALoID1C20KLsx/vW80PcP3Ki2YsZf14lJY5xyAf5vialQifPIsPiLJ3HHhKKLbG6ITonjWZ7I
81RPUr2K7UUhxSD41bpRVIX9z/NlKenfPraRXdWP9ekAOBw7pnheeDG4UQqQmwQWBXVzxIvxSLqn
KBmLXN6913NyFf6o71LkRJ6hYXRFN+Fuy6bzFEbYREkfet0WeLsbH2xe1oNxquegAJMsTsUOcxRH
OMIndg/5c9TnkxxpTro3g9GN3hBn831Id1f1LC2VyQmLJA3c2F+CtksVKymPBB8vFsNk9rmGPBpP
WMOGhkqtr5A8zrBUd1oBSl98p9qeo92/c83+EwFgUlP8pue15n3ljxocDuJiAavxcR9qnSRFuObl
HITAQ9wOgq/J5c/EFS/ymaTP1BMUcdE4No+9kgiLSLCpXYPZfOTh7N7wUPQdpJboGE2NOpl88MgE
xedOXgKMUCHWzNItlLXzdx73oj4ltRW3pcyp0UhQ0hqvikpwQsHWWqqL8nYpGUd7LjeUI0GaZtAf
mzLrrEoMohEAqm/Rf0Xi+H9jK3yax1XlRenQQRuNwW3gScCii/5obowgegdzGqYK+e+dvvb74yaB
2O+Do5Eq8SRzC6G4PsK9xcIsHMRf5CoVpT0D2ya7qvvHtP+V6QeWN1gVZvzharjbQz51aXd/v5sp
aIiv/7T8pcyYMgIxsClTvKyAfjg2th0HoIk5g4E1tPqUICS2BY/bRCbPK2FzCfifszBBpIZ084S8
FHDitrjWMDmV4ZvK642J+iVgJvOsQ0qLGZSQ2P09cs1S4eaa9lh7meLSAMzjPuFSMqjoXNYoRgSz
6iWzYxXI8Skc5rK1fgdUtVo+8gKFoWbpMFbo5hVKzZS29bxgdSijdEvtApTtVtI4Ftaye/cQe7sz
piKK5uteDT1JGgChr/4kUccKIt+jUiJKFExwLqSRgZ+o1jlzWmTLCwYtgAEAE0+a6hB2JrexT2vQ
3GXobkfyfKHu8xk+MtSwNYQL/tavXAuXCIArrOfl+Up4p3A7OmjJ+EOEttBAq3ivbw9CgwpswYBF
7Eoqa14hvESHfSDCGm5qOY2nDogINJeEUR4w3kk62ldQyPNo1BWgeeei8A4Lw+Vav2oKj7MdMoEY
6lc8wi/SaNYWZxb/GhUFNOH/xbihkXXqoUzYvyrsR8PJuxtJMBV/F1N9CgITWXd4XlljDNiC53Z5
n+UagA1KEjs8zO2nt7u1dI16YWZu4+giWbSYKwLlw4idmRgONjgK9lsyOUINUrmcWg6M6qD5/Rsr
KppjIjihcKsPmtuK4aG2G3QUNxcEowh04WhDVajZ6Ms9moGxA4Qx2xAnY5kBglDlhjomISr1I+WP
DuvRJ7T6vPsE9x+6fQntS2cs3k8GCxI2NnUGo4nKC9UkCwSVVcLua/OLXlSLjgfB67dc1j/i6QaK
KWd6awjBdLf76wsWA7ZYE8tPB/tmCigOSYzOhE4td1xifUzraoD3m37XSfxnUlLv/ApAHPSuysLp
Fd7ICBHyJ6qFaU0rloHegeIksdiTIYdGl2g6XzgOKxOcBZfP88O0au6+24wi7R6y8J4CEUhXTer4
CzITIFdGpTBnuCbxuAr0XjvtDxRCSDcehC/QKJab40G95YknQKFxkzmJfg1mFLMAmMa7jGtof2hG
7/9m/Z2tgwx/KF8HomKEZXs2yZhcFQuqAxOxGU0beSxNATqTJQw+ktsvIVLestZu0xKtnFc5bnT+
8Pp5YCGaJ5dwRDnJ8yr0/H+PWiiFil4V58LeMD3LUzdh5kReKrN8A6XcwjDpXEYe7Pcx6gOJJNyx
GoTKWyBc0IeV41jF8h83ArGplBcW5EVGqeVavhElhW/ujH/uErapUFQ1y58e22zfrROW7w5BjCeY
M4Y5Pi9Bd2gmvM5yc4/yfA1H6DRjml4PHMaLiHKBR3BLgk4prW/y84IpXc0O0Cecbn7OdpHKnB/u
S98wLSZGVi+BofzIffhim0b3MG3a1iUhfjcKEqhjasMCahfQeuOAReNDZ5d9UYHbeXM/YvJ3TjXU
k3pEkRCFH2QG9+hwBSozb4AYrQba6TYZhstePrwZVyG+GraOyY06I+x0fVtQY5yWGaRsF2hFI/cY
DC/zcOcMFLzFhAJoOtTt1LMtlQKyCE3GB9Cuq7cgqtwh+l1krQ/4VwytMgNWEcz8aE3AkSWqcHdf
Jc2m8NJrmrQnfcg2mOmerxHWfdAHxTo1vu8uZBznaSFBDqvpzCPAeTTdWs4q2BDt0xfHLVFKYXS5
mkJwfEq6J3j2Gr6O/mgj1q6R6is7AeFV3lpgdKu+fPk7woBZ2iU/tcXlAQcruHCI0DiAXlo883OB
z6rQtPfffUZwZwVO+NqcEX/87PSyho4u0q/xDJOcG2HQxOuCbf+vh8FIgW69pPnl2oR+/3bMfvRt
GcbQE4qy0yyA7iBHTfjDfahvAGpCL2kyA2JxeLTowVafBvY2jbqFESAVaP78Ik1dh1U2ba2nPyki
l/lTn3GvaDFKR/nDT3Jy14KYHUxqrXj/4L31FHQw1Wc2K4LBEmzo6zDuOX5q0/SYz2qk5piqFzJs
4+sR/LLTXJyyORq6wpVnuhzZuSO4hTVUmFKs/uaa1ByoYMGGBS7853QjZ8u2QBwOV8an353S6ADy
swXZZlt2DYoGYgE1Wz9inc8fHhb3mgLfLDY5C8u3hVjXYfwD2a9hVtliqQ8CKPsevvpqcLgl83bV
cVPY3JdvpLncmT+mKvQeg8b8OgfcMkjHxXbKCgbV6brm6xhTe9sTuvLtaXqe8+C+R4Dbwe4nAlzb
xHvGwVLgt7sUdxcJznIR114XN5ddD/lz+a9uPVefymF6Qb3HizqXjaOcbS9O9DxemLvhsEyimoHl
kLW3XkeFteIPSt4hwU54t4kedcbl/CaBfOh8RBRwu/GLDBRwd61o/wgpYQkzw36l9/bAx2RAjfRh
cHvv+fdgehAQbko06wvGU4Gla+eywHxEd7BwSiWvX77BVLKC5wYT2BBk7mbMw9T+AkW82zr7BpGD
wcXkLFiFRtGBgx8IpUW658SBZx2dE3qyGCBzOpyvcW8gdVFpXCKsYYHbt3IrY3PnJspXXOQeP6Nz
rxXydkFelwq+qn/vf2srxNa2idtxqDH+3B6zaQ36p2TOgzFZvKsBQeFaikoo5gsfuY/ptYvPzRr4
/ckgCiQma29cfYMbHiTacrAO1U8dMNQWRsGucQI1aXQb8WC4+ilN/ZV0LDWQrqJzAmhZDk1eErRr
Yw9CgK3N7xQpaPKoSvU9kMbl+DjCb4wNwWRpV+2Uq4yVkD5MAOvRn70O3Kawh2U4o7HgmL8VnlP7
DcbclD0m2bWimrd9Npg6Pb2Z5vc2F6PLAQZ1nJ/YDa5M0vL5O+DMhlux+n2UELIoIDTK2MSsY9Go
i+oxi4Ol9dZP1U0a7COYpkT0XImdT2XNwMCfalAL8TRd5v0ae5vhL22wvNDCVq8L1v2LSYOfKJWY
raijWto5keHeQ5Me9YpSTt/qscUzKg7y135c5YlZjSx85bkNHGUuhb43oqzbebzSHK6zy0CJn1W9
8+Krs24nEQuiATQVRuWpOx9+PPbZ8VimLKvECN5apY7+NVIBU6vKhS8SZyUpsilCPIryCe39JYDY
qJzN3/iJ2z+L9cHjfuMOqIPWS0z6+ZRBOVItiy6wGrUJtNkU7W/93GeCqSCXr/e8R+bhyo1iUVIn
XrJDd6F+i51YwHJGVGvQzOKUXVT9jDFW9x7wnsR6gOxGPwYMzBSdn7forGu2FrQEf1psxbIxnSF1
TdtGa3libKVcZUbGtbur5fIXPs81xxN3yLTYleAIcmiYAQNEGp7s2BOfluvtWQT9NOVs38kFg+SN
vlCZRZbmVk5g7BBPUiCWgF0+7Ytrg1IbTKDFB/uw6vEftQyKcrXsmAGYr9fA6FxWYUnc11s5d1SJ
VRKlqvJGc4AmccHln179cd76LhmOG2tnAdAvzL72HBvXPjioIo91d5zWe2+4FFmbmFBS8F9gbaYA
IFMLsLgtDMlROERWh3D3i3H6BKnobbXbWziU3bQs1THX6PQJ6kbAym4QPsNwn4cEerxsV70sxk20
UBbVxfHXT+2Gfa6cbeMhlnu04UIGG7MwMIPF1Yv3tYkixJS2U/B9Q6kKLvusZDO6MQT2hyPx6KdN
Y6Xoecxt5NvmBo96/Im2E+2QLkaDIhi8wBraZMVV0UZWMIouaIeZpd3xctUeXkkAQ0oNIgX+bNF4
V9TWmG0wnhVkOI4NTuQECooatTo66Fk+Jsw/seUEGoDsvkA3VTnnCsfY3uRSPad48SdR0D12K2tz
QJWDz9S63w6A51w5mViNGn7XxeATtB3jvYtGc8hX/qrFBxkkBFfe7aEKFNK960lkuhQjsyk6W6rU
iMWvVowsdICCXtqofmbG/81mcbbALYCc1lv3/ooqWe5mgGE8kj+WuYyqLX+lpYazSb7EaoeRoW/I
abTXsE/P8NFrnOTmu6Udy1vpkYeP8y0cSx8uHlGcQi5+oKddPMgYxAcPTFE9HfnOGjIibhx6HctJ
/yiWFydoVXWGUXMnMw/sIVreu5GYmteaOFfd3zvoM7wT7T5juLEop61jp2IyJj1EFHn76kdghY1F
bF7Wd5E8094iHTi7SQBKAj6ygH3lsZXlgqTqyAjzdgGHaWt+DXHNpz9TD1szB5maTc91Tu69++v+
7W8gKau8Tucs+06+46+fgsoft+tKYjgGKg4wX8rr6/f7gz2vS16fgrdq2jc9O/2qPN7bEkNGRMFX
XiVtgac33hr+6vhio6JmQNXjnz79ucmvJzSyhVhsPIvfpLGRfDtlxcfKRCa6amm87hm8v8Q31S7Z
TwEbuLEB3eihtC0IPeDPrn2GIWKw0UQ7WD8qJosX0cJfJRwPXDmGz0M1Ofq96ae4McQEEjwBnTtk
9Su0MYRigwUirzufCtf5hJXP9gP8hmZrc1wiWLdNtS0VESbhaH4h6CENATyultJHlSAKAYTlp0ZF
GscNdhMs9QzTG8aZbyFgkhnUfR797l9zcwyR3jIVESaKY6gGePCpqy2p/56Ng2MR1NnbpP4mgkA/
5lXtuqqZORbX+KzI4kxavbheRGZ48ZvuNPjhKV2CKdRWsLX7hgARWSfi8Vgcw2KJ0t00WyhTBkcQ
XpoPCKdrIUv9GcQVwbqM1liWGqsIpN9w8zMgiZoqjPybKYJkuLpgXStvjCeev64fjGDA2dm2faI7
yw6NNCwl8FUD20tvoH4mxA8imWWH3w8MyEb9VknpGGpSkePSwdhoZ6oSkpLsCU7QQcHstnV7rb7D
gMx5L/obXUSJksJTMWztV82Q45TxU3Tqt7KTsMagNePSA7hVVgxLufgdFLt7poTdrr4CC51uodnA
bxRQufVIppmcIy4LKwA60UTePPDGt5DCZLd0EXq2UOmRJ+IXBYgLYOumIlxNOSldSS3F9nBmPiQI
h4FwcfKIfCUbN2c9VwJ6jC3u+HmFMc0uYiDJW91xYEJWqtnPA0zuTyXyV+c6HA1yI/y+n6pYhTmm
WMrvCWWO8Bu3yMWnKyBt/L8SIzD87G8Fd+525GhBNKNtHsf9V45yEUgXQZnaECormPVJ+sxbrk2r
typFhBEQIus3JU5w1lSq0Vm/40XiKljfII7epwezHeaPmvl+nEp8tsHyBRhZRf01Wq3SLNfDzgrQ
/YfHvWIOI+8viPyKtpjrEmG5HI6yY/LY+MiBYEbp2DsQ0FZMev98m61JU6H0DDusSn58V+zEVoWM
4J1VU25ee7+mc1uDEhxBxdUw0jg1XMyHXPDLRGsYSHTBZZa9KL0dONq/91D5cR9+RF8g56zOqB0p
gl7ZELhTGYl3x3x1e7gABrERZEHrUqMuay0fi8uN6R0Cf5Q6q4ooK6xcIfN9ibH/gA5JDAfM9LxC
2rmHKIqZ+oLAxmO1507i/Foe9OEVKF4BmmVBI0S8hyE3p3qa3nGAR9JfWWXl7SEyNgQSFn7dG+Gu
G2PS7xGbQ2iHbGI7qVP/UAtzglcDxDDYWgPF4BtMcgLLdZb4Mrz0IIKqoMwMhJbUAFX1nZ2Rdi9t
btHePoMO9gDj5u4TcRUYIE9clqfLCbkAq83ehblKTxHTPEg35xIlU7h7UYxXBPiO0OhF9oLYekq3
QTseRujcljfBX5rWVM9rdpgJFe0edmhXavCLKuvRTMkzUgrKn377fiqWAFmggQwwozQd1ef5c4qn
JUfgc/4iSdy3OCR5m6V4sYdB6P45IOHw6oboc2AoawMhLid4zV1UWp6p6BkCJ37S7eDPNAeabkl7
4y9FDCJfMsTt8+0qqJ1p+SoSWC9JtaiWBZMU5VIneKH5A0V+PUYA8dH+A0vv/9pVeLMAjRVIuXq6
Wd2jie1XjnI2VQl5lqBF+eUbq+pEMw2CvdPEGg+a33I4Ofrtq4PJxOa+aqX8AZW41363B0tU8DJ5
yLmPn7VrR0GH8d4Np0pQoqBJYuo7IsxtCjM6NO2KgkYDwo2wXA+Oe6Q/wx5/4EHn5eXMdTI5rE45
nwdJAHSD3gMZyBB/SjyLRnW7FVJD5rfI9zixpYcHc8feGbxm/iiSXXc0d4u8dQhgEmANXfhOWyC9
MyAJAfsmBdKiturvXZLoeS8h6fcBEqq6I2j07mW9+AolbL83fGP7Dt4//VeglvfhvILEPbw8pywv
/peQxXLnxAz7oEcMHiOUOtJXaLZ59uzzc+P6x4o1yjEZOoVw7kWnUeddqCGIUwvVjb+cq1RLt5eB
c+AVHVBZ0b1QWcB82lNLh56Boc25lU0jj0+86aJNltFJzNHdSNVVUY7QBSv/Bd/8RKvIwqB37u/U
SIpuCkFXLVpcOfjf2HYXz6vg+ZgKkvgOxlZV+yeQSw49NVMxpHvxUcSkb/MFNFZXTB6chkjt3VMP
W+TQuYAQ2Yi6RG++c+GzD1Fe+uRY7L1xWeJ8674skqm9Km118pPHGtAfyu7nWQZKmdH/TKxQVtJ9
iJBY84xcuYtbVOfrrofiPAcPVcqEsdCpZjrlsw8C3WIz4l+CSrMkpsc94C4RUt5nzO+YVBpE6q8h
Zo0LWqb2aN1dj4dMa/KvOz2ePY5V6bfcaELRU7mjHvWKyC8D2jjALdNbkqdqrM9lZEtOxlke6040
w6sL99v1tmVL8w9+7Vu5iNan56HsOOBRjcaY8NLscnv14L4SQ4lNfwY6Z6s4soRxNjoy087A6L2C
O82C8SuQh4aRDDTg7GwzMyjOsx3YL2lWhwfL5F6fMecdRC4bMtxYS0qdDB9Yli3QcSEPdBxLBrOu
oOsDPvCrnDuR7KiFQehNmGjrLhihPSOxNOwN9Gr2DycDiodo+cMMTOQOB9pQokogLSj2NVukwH3P
TkigZM8n/ZUmgVBS4wQ1IBaCP9tf9nGQVkaZHnXAHpn5lXo1+VwPKEHKMOUvpLE449MPnHE39oAO
MiOxNFHpcVM2glah/IGFFdjof1AHfCBa9rYRZdEdSfQqOdyiBh8P2//hHnLWur2bhd5BH1pcLKkr
/gciqB0DesajBx6irpg3czd05NmMDkPFct97HBnczdcMxlssAK+nE2EiVjmplFxs8tnvI/ZKAOfZ
KHMA7RiUr8g/56OG11YYRbCDgQJvxyPaD2+Lg0aUk0xH4QBXM0mMKe3fsS04r3IY//HqQuBZNiuE
bzxuelzOH83BCiunKI5h8oH+DpHa+RZjnUY0geg4rp/57tJ9ksu4rDqLqSDLTGFdopgftBbFvgoc
cMdoe69IVZo4CCJ9MQhWYqG552Osh+eJQGB+hblpgRlkjPQRI3Fth3NmcOisqfRQzdQx14aX9hjk
lj8Gn66KLlDWEHAmgcV2lMyuDKtlZvaPS5i5oC003ElIR6YA+CibngW6skNoqdyFSrZsYxgiRJyg
IOVTF1PPeiGo/2CjSDgt/JK7j1aDGlCkJXLEruVakaHCpHqqTZ5nwIxDAxOsNpHxYF8S64G6XnpU
U1+ytAWtDP3M/fAxJ+Vl15Ke36Qd6m3EYFBJxy40k2MqO7EpyhVPZzbPdFploES7RlRo/4NbahmP
+Tgsti2pfow0XV2ErHxpZI33CNP2Pv4O2MCmRFOQqjYkgdR2mAKKzKGFsysfTCKDMGxsC3zU773B
DzIfpmwIwdOROUuf4CHrNtS+GP9gOTEbkTwRsBwv3npus/qDrKL9TqaPw9eUnTw1TAgqF/BhKo/X
IT0Lf8LVN5YCPBVJBRRUshkt/Zyc0DW4CzpbPFdU+imx4j5GXYt108GqMVsq3QkRJlEAB8c2pKso
FjBiaDsJUmwZI+ja++DnKHrEssMpTTjaxPW9eNRu8cF5wp7c7DsaN47q2hfEpUrMdZeYfZlAuV7+
tlKIFy53zU/pwh94UnjuwJ5xzZt1zn0zYugHlwfpDyGA3H9GhbWHd6mp5MxoQ34XWy/wRZ3Zt/ly
37KzemSvD4cNOmJc3L3MAoUHoUSyqRp4aWxokXLEpwHT+BUFpmOOCR5OGKjDURzl5IpATK/ZITie
1+nOccgGlw5JR0SiOjeCoo+Gh8aVlxb/YXS4LmsXYjEgQBDzfGCLQDy8fensx4Cwu23qBcY2oGww
DAV1C5sVQ6EETqeKmt7Js+hboHrq/q7DL6rHYaNtm4xJdGgiXf+Qa79zOiRUecKt04UVdIi9lLgK
s8KEyBMBvi1VIkhRdh8AlRuWK1P62vgSk1XpHDDPQ3oqgyh5gvvonPuwVXVusewuWE2lGTmuz6w2
Mer05DQUE6x0S+sb99qWBetMb9k5feMeSSopNzl6lfn/qdEhZRhY+rWgtOL17cgcr6FiemZE/zVO
1R5jFS598Hc1OlwL7KOXV+gBvJ4dLybhQixBxN+1rxMVqhkJ7ut1P8kFxDXB7sCuantWBXVrPAWx
TT5CBnntOK5FQbxDBE07c7cb9nqefOxhR3bdkUmPMwIb5cr3n3nloapGQkS62ag6ywYJTVKvMbYF
6aA13HPbNpFCRr9S09xkOTUDdZFUZkObv52D3fTEMnFhKFg1meLeBfNYnn34plE16baYqdMcPc3O
63JZ7Y4VieS3RfdjnzyfQgBtTX6xvgqEF4XsNq82Ge5hDnTgx+2apPbOSTsvr4n3qljdiagzz/oI
VdDQZcXIXDcaLOLV2giZztXYusFNrJ+J0Fl6mSE4f2DpZE7hhTrm+wmaKxkc/pm45Fov6lBzUgjP
OB55tdHxFoUAW/DiREVeq5RbfwZ3RlGIQWQ8WOSMLhlIXkZg6XAQITEPuyxu6PfCfmWqwqeB5ym1
vhsiG1TC8pisNkvljGZhAu6b7Rx1yYZQ8TJuxKjGcK6o63jmWle5cMx49zYtLuAcpcvbIZoFdqHb
6N17LFyId7iBmr30bC2378kwyobecd2zCCRilembb6SFaOF5Yf1LunhU1h9QnBWBPNf7jCy3Rsft
oB0beq8gBz3ae/vRfCePtRSkJ5nvo/gedtw0JJSnPygqLyn6QfA+zHWienpJa7tUfsiSWjZMOmnG
XIV5dVkiKroFrqlIS/H47yiEgoSpWbgJm5MbihqRi6VikJCViYV0ievbv0Dzq7sumuNx+gNUCdL8
7FFfdBN0iFTlFIjMEwV6cAHRiT6kM9lYx8moSYqFXKskzPHmLX+esLrrapdGH2Yccm+jwSUSaM8m
vPuS2JcASmA0+k4ZNyQXSAx8QZxhQaPbWIPskWWQpOpGrQnX9jgSh7pXzxboE1/hfTosfDuKWmIO
GCIjFAidln32Z0vDkYvC2MGkoqwqrpF0KbdsPCEMg8DeXsiZJnvyOlkcUG4HYWaPqGrgYXl9nsIv
NrX3PYFWQ+BtQGY4hlsdhJd45v3oyUyW7KXNuFrtq8xs0UKF2LGYKqCb5snkR0EKt49Cf15CSLc/
hz94MSLfrLpkTQKiA/yk0HOW5gpDc5oYGMxxLhUYjf7fY06btWmdtb//z0zf7dltUu9uUBW0rxbk
CnxEbV/lXnN9K13L6+DejS1qjyGo0NRF/PTz5ZBrh0O4IVSReRXWM6Nx0z6HLKN8wzYihP04afrE
QIdUTTdbut5d9kqKy/aKH3uZtcuG0ASiiUdDt3UCrkgMNn+8oDJZ7HKUOrWnuElngfJ/J035Kumw
EyogOWWimQLVyJ5WHias+0P1OSPCsjsvBSRCWAUyLxR90YfucwCM5Wf+ppTfmNcJvcAna5HeCxHs
Og9T0XD2qZfBlmiRJImOP1Xbi2cA82ypvRDaL/eOwyyWcpml/TeksHyXEzlgihD2piPkg8BaU8Y1
88F9F6SLNJ9BKCsfZtfgMVaaKso35sN7lTrTbJoJzS7FltIcWg9z7698Ogni6JfJTYatlD0DgSHf
RstMItjZ5w9xqUYHens26xbu0oKw+lQWx+ptM9GDrF6p0H1IQq3SER505jTBuIoF7IZrU0srg9jB
bXUhQPNN/O5G4PejBOUOYBRAHWh/gKyEYe3L/V/drA2kQOHhe6ZctGVrHktAidJ/AK1kTTZ9PYGQ
UZA1og+uGUed+rlClVelX1KRbtygUUSM1v/6Nmed8MWsN6+l9f5RAnGjReRBvoboqjCjWaeFo75L
QMMUQY5oVVgi8ImDRR71r/YGnYwGKFRNzUyPtwUs9t25nf2awvO0Y4fKQyEISEAT6DGxTVOoGSKj
qFx4GQ5LpKN0n3KFwJVIRcpiChEAPXX/hkpgMHdO26h+wk+2ZqVkZuORDcYa6GCYIK2sEkCo2S7v
0tLRHzyMAoUligzWq81ujoy74McI2CvjxgrKkQ2iDTpE+C6UE9EWkAVENYZI184oeZAiLid7VqtZ
h01GXhZE0jx7ESbYA22hsB3ydWp5cc4aukn+rAZG07ulLbuxwe9p+17B3Aj2Z3ssQK7T+rwyGy4c
inpUrmW9yPvu9CAxLPf87bWAti08rx6C4xzzcFcK2itKMckTe0h25R73gEMau+wSTeID6IRiAQqx
Q+vt7NGFGi6WgdUqJS/TW0J+BiEN31CDz/u82cwCc0p6SBnhR5lpP0IkV9f8N37T7pkqBwzzDJJj
60uw5ijAcL1O8vRahncc9bA5Cr1SLHnkNua6aDnkta+/onENX0gCiFdIH9aoyK68U39x3OHjVXsV
Oamk+dSxhN9HEYykMcK40yxgz8qHp9v69Dh/W+E537/q+n9/lKq3S5m1pWgFdCWa4E7sPT04zlOW
qXSqSlekDqhvfnW6Uj3+/cEihX3Jf30fZv7p5VpNq5vti3TL+vI7ZJJMPL6Li6hCDokgyPJL0BAT
6ReUQ53XpCc7NuRKBJM2TqiQ/WJeaZvOSzigHpvguSMloy1xvO2NoDNHL8JvfYjirEFQ0XVrTZgK
akBx9qoxbytwjTGnb3CKqsCW15hZPFVqLh3cYa3BlBIbJ86iei8eGzr91NNbirUgN3hc3R+Y5Mee
SOVgU8nKl/1S7QkCxiy8HgIz8RtWGhdfdPPO4A4IPHEhO1KoppsoLS5a237Tc/gCjVovyC9u5C/u
NP2WDn69CnQUiJWRdpx3e7xW4y7R4IrBplaNS3SBNQZ3IBKVaELjSEcHIoljNz2pzWypXnOb0gCZ
S1r9/xF+nHTA4ZcRLjpOgwaoHgD5fhqQDD4dgbNPn0rJFWBfolrzAs1XGpDSSWUEncTLs9Yi7eAy
yj5D9B+c7Oj23JdavQ2/Zx3uIPxJjHeAXzTdZN8zHyHU9Hk5qUU3tevPzSo8HrbG3Ks8owGvd3Rg
LizM5hOSCr12/1YigNvWHXRKs451Bg1biz2cGwnbxOieDwuwVAQQ3ZSnBfRsc7rBrq189TvK44R1
/48r3HWHlh8wzA2xX5/qtfk4lp7KmYfDib/+FYB2IFFEINBcMlvrtYDufqpEayz8DYa8ku5djzG7
H156a8DM6OnSlseMH3LSo48NAXkpwpBzQUm6pVFWkrdhtl8Um5kAeXHf8VqI/nYl4SZOBqGUH4HA
E3LCddS7AZwMEpy6hoz5hW43RDF4e6xqET6OifpnI6GqnMor8+bbAK74oqAXFWFZC8J4CZvWwbab
GdO+8R20p0EsRYevAYttS2JyylMUGLBaM2zNRZz0awLjdPDKl3XLGH4/50DULKJcaGw5RwCXFuyl
uKqOjTi4I9nWAr1OFz1z+UAloU3tITWRalLMRahwLxYlmAUTJ9IV0YwlNBBq5XRUaRkIvYqal9E5
Tq3Gp3LP+Y4E6EHaY+WxaTZW4qZOSNgDG3UrmTA49S5DGZJLA6bm+1/PgU6D8L60y9mI33pZ3Zv6
dl8XoTbBP6rbd3R+LD/moF2Uy2KV8W/bn9uZqs0ODk8kp5oxAn9Pi2qhzY0KLhyAJTyZJyahhGZz
qDNhGY89q6CQuPQ4Iu0MW0RVhh18oR6VLd5/tK0i9DO16PbLq93iwDjeRsDtYiasu0pv0yvxZ3c+
2wGAC4Hnn7jSGRQVmGtrwdMa+C/BE/u/5wmiXVNVzBfV0tsK9VDW3w25JH4hV39ugJY2Q6N/28zR
tSIyGjcFFNy/Gwf/i4hawMvG7nnXZWlPINCcDX/khjA6PkGfBjDcMJTsakiUq85ARoX8wKctqBsk
1soIZn3SolD/BslptdWdtAGOLRtGT9DoytQbf1R18imtOEtaCkikxpJ1gFQifG5w43FR4sVwc9wd
aUOkIpaBA2h1bsZh5CR0rd2A2k7SjeAl7Ix9Vib6HppvoJbW2FumZ4I5wF37vt8zpdUzYlnx4BcK
XS1FJoNI36SzYcL0mincioba5/SA1o77U5bVy6+MS+E8GnnVjC1xL6BgGkSXsV3ZoQYl8jDNWxKA
u0imjw0NEculhpJlDy40jxBAW8u/4FPWBGUmLKIJ5lU61Kayk5KvYMLY7HmiTKzwqVV4HzmBUWxw
SOmS0AgI38lnBWzX3p+E6q8xDcQkNEOkSkzmzbRiw0NzHPt0gRSqWSdx1kqV00uz2NJ5u1wP7fQB
0QQA/3wksmPtOfLQb46w4k5Rw4b9xAP/OqTapeVP7fQvEfbdxJxBVWvNYTVd9y8WrgD86UDK3Bas
dS567n5xFvbFvRW01tpaTkyAdxG4BhQ/aCeLud8ntFKZgB/xs/AQM50mHBN8pbE1odmNZqYCfPC7
JnP1RFEX90bm2C7i/LJHdaFg4Z/ASlicQxlAWNl6FAH4KKrqxVDd34UC+R4QoJ8pFDeBucrG2KlL
Ux1uOk6qAHLKUJih03v7kaDJzmtfS6oNExF0wOToLt8K/b9tufkpvPVo3PotbC/s8pqJBGafSgSN
Ji0jBWS2DR6D3qOY7WQCeq150JvA35hkRMgON3BksE0TXnCZWwCxpK3hOTkY+p4VIcVNK1SO+5ZF
x/5QPPpij2A1eluhDCGUj2NHElFGy2+dYHP12dlkh1aXUQZyuQF27sN2MpC5Y4qBWvyn8sJ9xUb/
uJuLHqLcPJFpKX7y3besImXf658KotVRhjN7LYiOlJ2bq+bwyJafajSIbDnHe0PHNOkWM//lc+iX
wlpH+EVnhfWVVDVvECXPOp+drJ5kg5XehW12oRjnh4A7/XQuGI558z48f1VaNDt5tzEjA0FrvQBa
3bP5RN0TNTPw7BJTLMZX3vPlE5SsAneCA6FCPawHymEwHYpX9G6URvN7mLRE1BHSam88+8Q7itbG
bBbwKDekjn7Lr7l1ZhpW4IF5XE32pXa7OHw6yPXsPBj18g7+Z491ySA9QICFcinmU5o+9s/KkTif
H1OIkWGTOmTxQv4i676kWrVCUg+vtHxp3X12uvsE4dLx80EQjgOvyn46M2R6aJyQvjI2nF+R22F2
9L/2NXOwY8C0aNwolFqKSX90V9lNvsOl+4g1GTrXUJdjTqdz9iEkbSMZ60h9jd3T37VkfPWxca4A
FrOspKw1QV8PXjxskMEfprVyk8eSckXdajy6TJV1epD2v5/Yc1gLal9UoSUNg6yoE1FyfBBCffCa
SOgaUjWldlXhDWJTUfUway7SxbG8PI0THTPn0mead3crs7mq/EBD8VqYPRkwCYAc5kddBgHRdY7q
tqx8nZOSHY+Pj/XMZsdws49yhGD/j07YEOXXL1lgowxdC/0SHMowpG3vTm8lw18p6YMqW8HITtx5
+3f0gtBBIQVW5N49K9LkDyrFVPYMx7CGBpDt/yYSVqZEyAqJMR7FrwEvnBaZpzkqz/I8sDkpLhnU
hu8RMLLsYsp0OYn2h94i+iyRoQxCYLUkmivrUeSapFmoLkfrRj7+9L91xlH9l9/6Hm30NDGlBGZ+
TPIxMbyI5bOR7gjco2mS3utc/PRhczDOMkbkmxsMMk4lZylvZpSvAATGljmR7y+Kf8a9s6/DSsXd
1KGMrxeC6nugF50kmx+Qwww564L2ea48I2BRNUnZCdlAm7pHFEx/UaCECJT88YT6B2UdQ/vJc2Cz
7/LVn/O1hLdKktfxQmhGYpJIP6Fz/q3pRPDF+BA8sqLuhFX7RU2BO01MlivnGuNdaKTXmBrfb7AQ
DOHK/p+cUkZPXRg+tzPp9z7KmsSMzrM84POXVaXURsdITyQKvUStz3ecNlvaGCfuZG9BVLQgYdqK
X8yOpFJZCj0SfBATULsY9uTTO8/QLSTu4ITiUKc1vwBVExQyq2xLXx0/TmLxExS0fh4ykEiX7rBW
GxAcvDRFlqFAP3wIkxyKD5l9gMA6G4wPwC1z+95TjjlQfp2VZPN0XvdyAlEpthtPW9kP8QUws55Z
xik4R0jCrzsxcn8EolCcRs6R280z4ahW03wvv3uoNC3puCgLzNqM9TMDq2mpTM9DQ5jKk6BOh60l
XB/HT19aUnDcamsXsCFDNHmExVYEIWMipj40jia1s1J6gbeDqLjpnCIbOSXNeiiIwDiQMF7RRq9S
krR1GhaMZDx6LRranQiFxHPt4uU7owjFRk6+vvOs+gXYxXiXNyo88vFUkiFZUadu5Fca1qYpeXrh
EYq36S+exbDej/uLa9nF+egyzD8QV7cJ2rouU9LiU24ox/VKGtr3Wt7uv11re4ftJ1FyPE4iCT9K
hBGX3RHZGtJo0eaGThh538aiVo69userjkX8GFJlNHTah+WaKLYobIIoerGEr4/UIz43C0bZcGI5
oNVWTNNqzH9GpcgxNr6RbKFY8NPy/KFcrhxyi4UIMzSPOd0BgXRDLoJsBm7MrMS4AFnFssY0EWQ+
R27GbCuzWXRpK2EwBLPFI5jZsVtHvkFXqY2zW1DUXJHSItAx7N75oivYocM+RPBHYk4z25U5bX6/
UkMyGYcNOo6qXfuz6RjS2BHl9kWgsz3UEPoc0n8t3I8o7H85rzkCK0oO9hxGLVNvo+5l/uyySCVp
oDx49lLaqL/QO/Gl5Gy3GGq+EB5AjhME6bty5YTNJol3Il85rqmirkPrCoiQ6vuIat52xUW2N93G
v0vwgC4PxMV98ux53heTr+DiJdR9nTONsO4r6uHg+sHeGeb+kCbE1yiqmLcLNDGsJqVCU9TDhbmH
XjZ8xiW1y0JSsN5I2/Ngr8GUUuwsdMiT8lJzLdt+gM2Y5fuQn9jMDBJpRWYq8VAWQm+kQCNwKyOy
Vmr/D+RwgBzoK1SbY4a8Swvbsj+B+fPjVK82X1hkwtWEUiY+MR5yPtFLxSQLYVAHGb9L+uHpmg/j
GQHuLYgwiisj2bmK9xY01GFTteO58OhsrFYXRMpzLIhULuGHEiscIYxQ+GPJA2j8GJfmsjswx5bP
CwMxIBCCK4uOlFPpfo+WN/vF1IdZ+zdsf0RqMBvA0PVctX1qGU0uywZKypGd04yX6gB6gmnzbU3G
oU65cPBKBBtbIMhR7hizY4rO2s5gnenLcbJTaVJOEPsOJeSY7/nc0G8GO75p9Wa2bTW/6XrmveSx
ZTkMQ2DHckDQXcMemLXJ01EGrWKiH/3WBoibacBmD70JMoRepdR+wbFgWHAN+uI7l9T+uf03oC3H
dZlSoW208ug6HH3B2NrBJV0QMwS0fAAepBm9htRl/zb3IDcLv7K1tGXN4u7IDyKkaO87yyXHvYkI
0GBzoNBJDssakNQj4a/N75/YAfQP+xy3FyANUofVsyrxC9fgSPX5pqMGJA4T/c2yFBMe9tl60vqg
WsWSUC015yVWc7h5Oc4QDTeWzRNhToNuBIrGdYmIFunbjn+V+5ho6y2N6rCFH/ZfeySAJ9+eabU7
Pog2v2R2a0syydAEIAiVFKmagaHMxrrUUhwXgEhZ/4F//U194ucleuc3DaAHBRvkKbNleDfhj88j
6lm8kTPTm3peuyB7WoDpHF4WqlCp7SPSZMuGkWxjmp2JyPlaNUaVt2LkihRN1LYLut6+rcIBzHhx
v4QCE10wISiW178BCNywM7LdhVusEM0aclUjiUUcgDUNDNGspoqw9IaFPZukJZq7DiX778zO/bdW
413bL1CvWf47JFjhSx5Es7dqJHqgjEVE+PhH4gnQSXziEQmpJwsX22r9JTTDB3CB7H516SvVhVW7
BCxXJAAv4dMfmbdoHrgL+zqvtlwToEoFS2sk3pwfNyUKh3A5sH7RGn8JCjDt+6EnhaRtBKiSueQt
ThwE79Qf3JMrT+wTvkli7jOnJUiK7CxzzhHIAt1W4Zy1dfp+wkZdx4Xcsdh4BIIiBHGAP4aQSn0L
KOEb/GdHD6t4wCHITzuUIH7sfyFUdZVE/aiZrC/TRjnZbpwiV5pwtrhkFCU6RlUjpOuYYUy+qb/R
gyleRAaIjKlX/tHYKiqqIdPhO1zRmzYvFTchDywaCXY8iKyuKnDme4zExqKxAGmMEjeFMIr66K6d
pieYXwPJF6TCIrwhm103l0L736MR8CzdyydvG9eEMFimD72LFExkpKWGSjKe3phY9Xy/K3KrBgsi
6bjEf08Ysb21MgVXPZrEyOPTcHKJn+Ci+AXMqH55FqOcYkNKAhIrTgVUH6xkb6yLgh5Twr2xGHlW
saNSXrbDul5qN1GkhlpFpbAfnnkXTZS7lxHz0t/Ga4rWtpoHiaXyftKqQ4CTPoN98TDw1O9IIdsr
xgLgKm0oh/nwmnJxRaAEWJL7gJDwSCccNxY7cG8qWgvrAgC/8b+HDli2PH1oq8MJ89ROoayfTo0j
7KLSC9XAeEbRfOqLGvTy+QqLz9XXi054HwSL84X4kraP7D59kcw7XJ2AZ6znT6qD8EpRfJRF3YIR
hOg48oPTDs2G8B9Sl7YaasCeAA/t/tGO6BBP2mKmfiHal7bJWM2EAzVkO8Z11r2BaJHbTKS88mqd
rINw+LeIC304l2DyKIJACACh8joGnadiK+rzdzSZey/hok1XezGFiDjsnq4NV7G84RbCeNLX6D1l
wFjCAWNcR/sKohFiK5xm0AtL1qCTLpAJL2B3sJroS8UGAdjJGK/9hNQ7C6wFyRn30SfefYmw6m3G
zl/632bi0cj1TZvkFvfZyDhjO7nCO6cDPWcf88NhbcS/VJEwD2LppQY05A4UDpYoKuXgLcBp2W7i
AEZBrJJIixYcJB5iO0A8VCXuLJkNl/PQKVu9pbsQvCOh9RK8laWrEasJt8UML81bSJkUqUv/qPhZ
KC0IMywgvy8WvFJwX4uSJqmNCWqON3USAOLhOUUHGhH0E2yIsgcd4SEBmvqd3u2JV6AJah923XZR
5k3ZqJrNh+vWnTxGMjul6a0m8gBPU4NVyoBwBfowhZtPnNM90NfHYEtlujpzrhe+t+r0q0Hnj80p
mAEqrkZz3ux6ElEDTyyEEJdSr/G2B4C3rrD3mJgDfdmSs+GD1+jVRl3yScCJOj6X3DhfIPphzbPG
wdRpZKJc8DOTihEO9Sn38X2TR0tgEF8PE8KqkG0AgqqLRE625POAru5B0BZXqki9OT3/2zy5YqRZ
+OnlipAJujo5se21KfsoE82gFJw0t/Hd0H97MlQatEeof+cNeHrNiFwRTYAkyieyp+X209vDYoK9
XC5AIpAEXCnJJU+ERTkSxipfxwhM4bpoICwJFNFQdi1lElevtny6+pBjofxcx/wwNS7Aq1Fr4Ilv
AZPSPCOJi8FCx6fHu2VKk18Pw5BZRd16nZiE5+YDfFpJE8YvJqWbW2lQigbpf2qhZtfrzs2iPNZs
J7ZYw704O+8Odln9gsjavO6KOyd8MiFDcdn4ljQHEbOnyeNXatnAtrFN5NvrFS/4BpTadpU9hY7i
+uMZjGwQT2AE0hHA1Kcf6jIAeQGG/jwq3M1x9CztNPgtxWIKLBUdCk+xAQ36QdVJAgjYQhGdvDfp
di3GZ8MAy+43yaQH+uBTwzZlnxHIlGb0qoRVrepYqKuwbgtQxpYGKSYtBRBbkgeMpU9TP0OA52gl
0MdrG9Bo7tSmyPp1YQOu0J0EdzSx
`pragma protect end_protected
