// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
leMfNUBsRwCJJFrQtWk7LWMwsOyVDLhzdm85Am6d2EJB1hpW2xcHZhZVkQzsJHct
lJiMpdwpF/XKJqNw3WUqX2b/rl3OtzoSHTHOa/QaWl2OJ1vzO/qpvygtJBv7ZCLY
IKAEG0Sw0XmL7qmo2Tb2uTbZWCsuu9wO2km7slB2NEE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1080496 )
`pragma protect data_block
OfzqEvSzLmHp7V6mj2DBjmdc5rGOJobA03K/ngp52YKSvw7B7oofouuI78jx5iYB
E7yHOB8L0+1MrrocqDshtT891gzNsXSj4v7tqfiKUn9VKk3FjS6oO9A7ujjeoKuC
w3o14Xk5IgyW27c2/PAyL89vXkBkUqQjvJdaRkCNCAUzm19tU5CVlOdU12hnXaoM
Ll6todtMKPg61wWCf0qXtOJ5k12Va1MdARpdkT/9oZ39VbGvWm/sTrpgAofYwy9A
ll1Igrt6TYEkiAEAD7Qa3KItLarBLzCdnitouZBBcTUy8JT2FHbUMK0AsblkJJkL
piiFe5Id74SpDV6oIz/PdVcKaS/Fkle09njzvIwf+3A5sMy9KzetVxxqPTVOgQCp
b4Q7kSJMOJ+oOBddOOTqk/XfjmGjHan6TXxTdDs1AjpEyeHEO45wIPjRIE5XVQGK
EMS+ZItuNSRjBSqkDIzjO45vI1Zyr8VasXADUuvcinVqmaCBmRiObR4YvZvAFoXa
qO/UROACY7SdR26zE8UcbHIJHIdeunHbfoUeUo/tMqzeYMm7MB3/3P0TOfF8KXWB
lur90dVq1jsKUBHkoEGnkA/gPeitlHpcMqFp/vLvY+ATG8VE5yAqQpZRAFtr/FJp
6yEpqd5nvHoa+dT6ufbdiL1Q3AZIFe0DysAzZw7Pd4EUqeyvtbxQggS5fwLw3Qyc
OAMCV+HoO+rkx0mPVmv4CdjGjqpvPdSaKj817t0CrMxjVedaTSIMgQzwsTEHKQL5
fiDrCmsm5KU1hV/U0BpLbV1J8daMkKjlwfVViTI4qbAUB9/YH7f677Xas82FjHT3
kWCst5KkvGdjzudak/mRbiRib44Ix/GRVUBAA8pup2JEaTVToHtjpESYQ3UMWnWa
QHUMaiqXH+l+0nPfGADeRSFx0mrqgklTza6qBboyX2zWE30oMKNR+4PV+Gl53Dxr
XQ8KUMMu3GxRxki7ftGcy9H38M4vLXzeiKSXv+QHV/d2CyMRYy3DszCKNwabUDmE
4CNIIdEDbm0Xu5OGcJxrhC7CEzycnWFA+0K+sBwG878nKJhzXs7W8GctFfC86NZs
r7e9JtayUVCP8oRyBCqmSHjsGGrnOcthb3d56uiMQVPGisCNpv7Qt4flDs+E6MFu
7+fqGFnmls2943FaEv8iKLHAbLfa8iD49CnwNVi27NZLmvh6pXEh7ImX2YmCycCc
fm6GEO8YTjESdKGuhXLv7att4ntEJB3xSSOUT5LUxAZjLCwOIXKk8755Nks4Yb6e
drqsj7XxtIRm3w1OjMxu5CsUAynamM7QiA1kr55vhe7MMw3F5+BsM/W8bpwHdQSb
YAE1FxIz61VOU0Kx4tWt7INuP/FveQE5I38giNKq/SX6FkeI3ZpueEhRE4jBjIVn
6CFMx7O83RszIok+1Lxk09no3TDNCAUxU7fRksQ188s4BoiMk/9DwEhq4obkmsTn
CQrgj/PgXukt5yzyL8FcWpz9D6nS9+eIrK7mOlBHC7xyuDr2Stg9buANwEl94PPF
T4zDrjfbakCBOJLCyJPwW/hxfHqRKmrlvwAXa/URTF6YwS0I89a5hpU8t9SGxWZT
91QmZ/hEgszUejIMFbZ9Kjf+i8dXQ5c9SsBAB5oUIHfqYwdQjhXhd/Elmp576oJu
E969w0EAMQ6S8RM11ph7qZVhVx/RPhSPjDOSHoHWAaM0AeQUdOp+frvdoNupemGM
pUVAA24jY5u9IJP5rFpgKKYlWaoQiSoAUwtTZH4hGbnfPMQNNLSZKgEriMDgVprI
QKO1Y/a8J2eLyFPiuTR1/80GbQx2744XzSMo7Xdgk0+PpMTcQvSKomZjYzx/OH/P
55B8FCQhXdzTUTVNyhsYN8XKnoKVPvbtOTBzl7OKyiawHwlRz75UHNB4JfvvbEi1
fEvsR8IF0HqM21YekHKjtPdEBY3uBGGMnWKhwDRX4jri9lNQT//aVV2WZsfdw85b
CbakfRyzxNr5DWJe9JBz5QIO4ZeoAtEJ41iB/3GbGBD3p95jHA/333ATYTfpORBa
QgRo6v/HA5rZtrUOz9ch9xDMT4/RREOtiib6dOg7yd5gJfZFcImhQTSDWk6S2VEL
YisacOh8LgxapqzAEIQXj/O7B+Zb1+5YK4qjNZpmvOKwk1vFjh1g0HAmwuqmEhRW
/sPsE8KjObLwPeW2dQExmPILNfPRzZlttoVilJqUQuSvOZrNOAbftRKISeKBZcDV
XPGZvIoL+rNH4sFKmpjiY9rUf0oBBYFSYqsogfqZ+lYKDT6ueVEpsi2qU9JzhjBp
hipcIednQhVcIk7uqxK1dAn0d0L2BlJTudJHSgs57PLuRysC4ssIrOOEpU0w2gK2
oUw6nTIEqhzjv8WOwyUqXKkpQd7o0HZzKj14aeD/Gk27UgQNilJQ25ECeiXdJrbv
atK2x2XNmFzWn2aT70gBI5l9avniDI8Xe84qfqAsvP8JfoyTs5Up6drmjqiRWesE
GBQ38Pf7/V+sTb0DgknzyFncX+HnsD7QTr+gqh8o6NYjIkVuZX9d6brmbOcdtXjP
XuBoP1MVllumSFbkbu0pGMfmUm4y6g4xoiCcN3Ky3sTZjwQ+NgP+97whtFly6MKn
TBvQNDPhWxOZGfZ3BDMoN6l1/cOn/On3XKfcT5XtSNRpKg1joVpP3jYmgr7jPQQ/
XMNPlVt/EZoSNks3fcr5/Uvpof38Uy5N6mapns32vMX6uwiBTJUeHR5lHz7b4YAI
b6GgVnVgYttFKFyME0YO5plv1gs/XvqMe3rZYMe21k3vQ/bfrUZDRcsw6CIy0sUg
2N0GRru9SC8/QXNFGXzBOX4KSmD+cquZY24uKB2KvfdcjCwgwkx0zRie/Q610RO7
6beQv9/IzqyB75zEpcUif2YXeE5NqM1iRob2fTm26ImIJHH98lkIj5PBUn7SVLkY
/wQYhSpYojIKSN+w4rm/hrCkx0n5nufzQ8Q+ncdpQJ68JV6a02y2Nk0/3n+7Lyti
FWBRLzkPdBImx9Us39AXnlqzxikEPv4/PQW5E6zT3S80KhjA7n9JijogrKJJuNWU
+lqd3aahqVv6p+E32sUjMwzw3eN3uFpIZ0NbVCVheTjW+5ZXBT2L3TvkFMXlLbZq
2ri0OhZi5g9XJXZK7gHvNtApr4KP4BRb4C9rVzFV8DVJspMyR+0ZUsvPmN7/ndLm
9JnBNzuGZGefoJwh7zr8RnRExXYVkkPnv7iQ1WovmpgwM2uwm/eo4oVyAFCNC/i9
uLCt35JYbXmNARlQHscoU29WejLAY+t5uExo5ISRzYu0QZRFjz8Et8MLCDe+xhzz
qpPGzKTw+TcdZIp3ptcMjoFmeFbeXaAnlZv5zZzwxwYaev0fR1kEvFB7/tZjb4hR
MF9kHuSUL30akKqPyAJ9DylhthEsHilYvew3ze5MwIhjc8wUAVAmEQLq/lKjcEKW
DuJgkMsYVPiGCRZLmjLgsIhXSdh0AbCgDwpI5VOS+vvxRJfyzan8dVzEW/+SmqkV
oa7qc2DHPnzbE1ZHYYOOAwFqiEJqbpTsjoparo3ZCeu0tcbE6K5ccOpKZ6X1X5QM
plik30MxuwLBCo7At4SzQxrkS0Q3RT4FaD+wwyRnzF4ZR0NfBToJ60ubboPTUvEK
HflVWBFtPOyT1vUyLqSb5nU79fcwlnPfuqPZxqDX4k7zQ9/CbKyGV7LBuH6guIZS
FG2NutWoc3nz6S+kjW67VlG0BHyZ2ON/n/mk+u+bpaL9nvpWQbDthc8OdDy7/LWD
E7+vM2OeoOznZM82PUN2kH2r465eaPfO2eljkw+yU43tBWEhaYq7cj7vSGKeQErO
JBFma873ymdHQWBvr9lyhBkngg8y7pvB+HgyhbFvGqKvQIB5leL6qRSJbYMaYdBM
FPSMQx8CSoYjNobl4i0Vg9gqZJZjx8+HL68GtC63o1UIITEartoAk9lqIsAuaLYi
ctiognnbPP+unCcIfSvgKIRPDI524JHohQ5sLKxFd3sgN8Yd3zsfCT/W/5bisRfo
ijomvPIIUVdpgQFX0FNwV2+a7EX4PO0knfHMoHa/NQWfVPsKFTPR2xYQBXB+AICv
oGNhWp2gPXgm0gpBDAL8PGNZFRoGSageStqi81wNmnPWaGl9Ajcq5KCxjicH/4It
wgCqrEUq0O79dh0Ui3iN+UaTkiK3ESuW8qp1y/XGw6w+BzeprpeJiDl/r/9v2DNn
NhuQ+Zup1EcT3erItWxuHKvRBWqTUrm5ZgMJ6JDXP8Max+lRChXxCajr3U93vN7k
QtBiqU0FUCER0wPmYi1z8bWfTYop8Pu9g5inz+GEe7NGgLABH/70bh6Jol3n0d7X
pnwIF5l4harsBpZ+dFA+kZ+I0Vy55RxR7nm/3uwYGgOjxZLWqQNRO6h4nAymXQlz
k2wXFdX26Kkj3xjsHvpQYBSr0xFPDiBcHedoS3K4elSugY5lyJWtoEUvflGfd6Ms
40EAjNJtdNrqjPuOqw5godeLbMg3qYmBhMRqZE2lVRldcWiyDf+wmRff+tHKxx4g
n8bXbWTbpwZkjZHrIHg1MpKxlZHiGJGOTccZOZsUdeKOxtsy8+xxVXndgrZA+5Ey
4So4MkIox/iKsqhA8RgZIlIpqbNe7MPPa9yDIf4nXUXpfmw9OGzeGI24Z4k6aGa5
0qecoY28et8MwpdfjimhM9H43/+jv4B+jQoEsB5Go6ImeENUJO7RsqWI3LWhKRGC
k0iAshPddinZesODib13bOXyirM0iv1sCfAwf5QqdYS04xRSV1DD3+Mib1N1Mans
bJnd4uUK9n5Q7JfPYSR5iunN+gK74exu2ovDfD6L/dKQ3hDU5AMyOp0FXQ8l4nOv
IhjV6CMmk1dCKnoYVdYd4Lzg9Zwd2u2ER3cviSUNAJhuBsyst3f1zfWYUoh9sIm+
yzLy2ZcSw7pTUGnQf1cBZ6OMvE4rXgKAW5VnagOS3w2qeTU5MyYPqrkdmfHMFbSJ
Pcna9jlZJC9SqG21xPl2x0JcEiNQc3JOBw5K/6B1dlpGymyFqftbGqAWuuZmaz1l
ZzQAOK7WH5tr1BmPTDA3gKc4BhD2IUPgl/N9kp2XhUD1xG2PaRc6M+63xHxX+0mM
whLOp9G5w055o9jvn5TSm8/jjt/DbFD7Cp/B/DfdOzsdiykbpwfdlWKDlMZcPqLR
Ezd5FHQY2lrgYyq0CdvA4NqaC+LLm4cvt8/NTtnWFfF1LF6gC8EiV+SOo9MdpJyX
9lVPnjP8yML6gOeEYVdlEzQxYmoTLd12bTExwdXzgxI0dilSQByLgOqGLshDWVap
a9gMp8zkJaD6LsZQsFL1WfFD32GQqhTJtvXDTiqcXdYW4Uyr8JZ6rfyy1GEBWO4T
UkbDodgMiY76gpp/ZFLEiADQQnHsejOmqCw1PQA0QN3Z5qul/hdYNFWaaTBmIkng
XHcbb3uWFqnwhNvMdnMmGOGAb22ZrqhzNqQJE+jbfqy+K1MQzXi9D7twLVHOuhll
7r/Whf46vSkQy+5jGBBlImtCfmUPQ1zssNiOKT7WdILuJGgmsbC1df+fF/IlqKo+
QK9j/t0wUE2JFbdnR/icFXgxqNEDWhFomats8HHWXKB5R+imKjRsnb97QIgBHsfK
sdjzLx+x1KY8GvU5UkVrJ1hB12umKWMN7Lr1o6sC/A/9HmECPLlrqrZtcI4Jz0ZS
E3YILqfxRAS52W0uL/inEL1C5Uhq784qOBiv01BSj4zmELg+XD6ohiTk6UA8sESz
PAsvAhRaBPA+988G7/frOPyfyKNhyGUk6zzzHjRZD4QV5YcJYxPFimKTl5x6/dh+
HePsl89I+I8bct74lsINE++hMKifky9HYPUv4TAyHv/v3KH/tn8at8dWlSGLjMOU
cXb5XEaqEFgMOuqQ1xhQQyzAXCR2KqziGMQwRzSwGrL0cFtb+UtMzIn6uJ40kqDH
CBkqAjsMzMeM5aYPVoc4AfZSSoMTkdzkWWcRH6gJgNLSA0X/eMDOKOnkrZmk9zTm
jjC4M0w5POKfq6HLNg75dD5SJCwQhOb11rP8h+Uixc45Z1Yryf8AOoPqHgX+QUAn
iN41ejKrpvIAnarxwEcDfGbYepBSZS9e1RUOgV0gyyQBSnju1+9xYwE0nT4t+YQN
EY7PwdQkgsBpKO54NdL88J4oGNwpheH2mDRUGdvZnocqZnTfk9REs6RYMlj1aamE
qNz1AZAuqfgS6WTZ4toY37QCDTvnFeb6WJhVxmi9TVBaKBGq+paT6hAxG/VrUXHR
coMeOCC9Rb8xZhpf1BVHNg92Xk7mF7aXaX3npXx0H7a0C0fA/fw6TS0an3rTpNC2
A9IAMGuJtPOYRNSMY2xIUVn/q68Bt0WHQxdIV0PAyLTRs22JgD9F+e/ee+fPsWED
Z598Ka4/7El5cYH17m73AozVtU68KTwKRP9jI6x74rPpSMVoWFY5HQkoI2wmJFlT
oXACrF3VRA/Gvx/4aWrtcMN7RnxfHsM5gShGwTc/2wBIaNMUJQyYvM11JEczMwcN
oGg01e0dG/ISRPoe0X6sCU60e7cwT5XEhJG88mGd2hbW9JqT6O7Czxd9Laf9ea7M
Ogj4OyW9lk1KerfTi6lxoedBRN532xB71bLVxnOsIYETeuabylMEaFDkkiPkKp+i
KgIlmB15lU/z6xX2uOU6qatpld8zuB3tiGw0QxvNePQLh0mxspp2eaSSJ7XarqcK
foTM4cZ4yvR+BSC2YM012l26RDCpjPtzQl8zG7NOFi9DhxZIEUy9NfHo8xFS2D/B
KB6xP3iYo6YIKl8i19FuYfWro1LiwzopFQanl2PUPf7eNKvaKqdIB1byfoKYfi7+
R2iiOqS6ljw6g8qTCLncRKehzhrUIA4L1qUhwG+mCYfLuAL6frcK8t0NNgCeRmTh
JoIkAhO/TZInUCKrSP8Rhp8KNB8R1hYUSaIVW+os2MuqKXm01PjMRsjcM/v4ngXg
5q6fFgv/TsrXU334/FC/hinjOBKl2oBbOmUnYNyX3jpBedNE6pl7xT4sJ6Kr4ntD
4xmoHiF+yeLQtgTGD3f+TqcRBk+Yh5UGYPg419GVwdLYxQ9InoNJn3lxXB+nqlsy
+VJdt4OBK7x0JFyzMWLuhRAQlAlXxlhdbUnnaichcbDSRbLyQRWJnXPDDzbzKx/Z
zGCuAQrxw8YJjU8P076X0JDDvM1N/zU4xet7SwN3tWW2mWxwjpXHuL4mxOb2XehO
rQAAwfatcksyXG21UoMTsvm9Oz+TJ7kq95yyIariDpowMFDwOk+Q64YIuWpQas+r
e6VA4UN+Y6ZDDslbxlsIuV9oJH/KdSrLT1Qd74ZS/nWQSNbazwdcELaMgBUPK/H9
cqnZ6cxUGGpLpOmpH41Cp/R1zBCIfnTmkCgZM8nQTJrQuf2hLJy8j/Y0288y44Hj
qop3XnJMsQjcj0VTULcpV5hId6K8a3fw1qyV6mtEaENB3qyBNeA/ARL5O0ItmgLC
dFEsFZrSV+rcrwwgddV37IQQ+nbYXK8475+fw6pvu1TILof115MAKeWb8J106OaB
7e/VCLgFmy8MegOJwyrHv0Fl7i+GQtyQenQNZ+iSm20hWMgXnl+iiK7YJwKdNhX0
j8wzrNjEd9a2UVTtO2SkeJc7NqAb6UbreGllGQCc5ZUaNIenxxS87eXMiZf6wXg5
Mdjc4dRq723po1X2u9JVva8kF0EQXCM/xkQTQ5h+QaZyHCctzQNoNgCghBj78xsZ
6u71J9DcwWLsnJvi0hPHzkP4z1K04wPvPPWEeFTrqXc4a6YG0JQVUWG0oHxveH/H
bTGs7CPHfNEqQwKv1hbtrnap05ETCnt9uPXdImc9kMj4cxFGj2GVxAtOzmZ7y0M8
T9BzspC2+gTRYqJOC71cPMCOIa0z7F55FP2zWxlOAEgQW5Yxj2PMOu9u4UBg1/x3
zjJLBlLOKrMi0eCLF04YMXG7dKghGumQWzSsBiOuLhIJmN7SsZLOwWyNPJnY8cM/
Yppcm5fu6cUQsrihV9+YncuzV9F0bCeUl3t6ups80H85PvCJrBUEe2IxD7yhBcIW
34VlDa32HrTod1305X8j8t6Ir+ugdf0f4H0rPH2rfihOUqCi4VO0Nhlgh3xJTVgu
589dNrbP2PZsHh5JXX7aYahaq5cr7CnBrmgrFNpjjd+AMEI8r+dtpPhKKYRpKCnN
yhRaKPmyZNiTeCfalPnbca2hdTg8R1AOSYNmPJiGcl6d7yS05q2X8SCNZx0mcigj
fwMYfpoVaCYpOA4K6wm3F7xbLHxLGp2pvewWJbUJ6Lg8p3OGmKA2iGV+I4anovof
psjIfpsyAK9YFQI/eM0/clw4FTYpD1zoHhbUeGPYWcXfttZ4ylKe+6hq7DKOtjXp
Tocft0cNzKhvOtxyhsOUBNd7OMGQDka5PCVxwmJP6YXkNgFN4Q+cIyUuMpWTsqL5
cPwoFppU1nprJYu8wBoHiyczCDa0qPWb/4+29hoNr780gdybGMVNT0no/OJ5Q7e0
GOfudGHAYOFrwbmDVxCQcOUa4Vvx57ScfK2Z+lAsDjM/HCH+EIF2Tm7xiGPwfeqV
wVn3tgnZ73BHDOw/RbfBw1EfpXhCKAJet0jmoMd00HGz5OnRZQnkgvEIizolYe6y
wqOfmwN2AcKzvowhiR4uPMuXq+YOeHaml45l3I51ctrRsaUMSyTgBvHLYK/ldE/b
0Fz3+5ARTtrL7y6ORNKK/t6bAuoTU//eY/hI2I+dQoa7v2R0o+w5d1zxXG8w62Yh
RkjBbufwzraT2t3jIQCLBdst+mcr+YFYk5qBYhBtAJY5fUMkcJ0DVxz4RE4Ml5Sq
WTc/RhMWbJ94U5hZ+FMYvSXpOCgWdf84srlqIgcARHmXgLsMhcIIgBTMZKouHFnd
8yithPfS69Sg48Kb7ILwbcgEj7EHG+eTvqpaEwy9sBIbErDQicdMq0/zzLRF+33Z
x5HYUsRMbF6ueeTW9DF27jE6hQjovOFWmVAN9GRmcTPiLa3ooKbqWdJ7V3TYgFuX
SD3Isd1Jw7HnVVkUythPJ1etP328T9sBPONgKooOfjk+O5wKaaC5s5z1dSJlEzx9
We+VGcgx2afLacQOloVWtZ2RRqfV/DvFX5v7OM2t19tMf+nJGm3TFTkWpUPlyWkA
0X7WVc973u2bFe/VTs8p+/juR+Bz6Ern/EsY2LuLCJ8i1te/VmZLziQsOun4dOFy
I5uILbTCfbRtuwTWGhKFd4rvy0gWVTyIxsno1x1xOJ9bJmUcSyy1dDBylq+n2NPh
7g6qQdkaWGThpZOLnibmgR22GIYB9n/0AuX7fclDDtm1I/P6cixciP89zQKPqnbr
24sbcge4evVRWG1xXrjH+T2a8vRCVqqN1m725RZ7aVftTi6eu9kpAyHKMCHNWu+3
Js42onaXHTof/jyohvyjhsB4141s7ZS+Lpr+N9dwsccVbs6hE1SNaiOOfGDrjIXY
0mM3FzHIDxb6UC/4Dj9qmbW60SksRbO/Hn6ZOTJQ6wT3BngDKlywolzcP+rgc59l
QlpdO4HAZaLPSk8IK/R4I0nxiz5u8Upoh9+KLQ1cU6WlyoeBdqyV27ou+Q5vwifu
/YnJJpmHpBbg69W2NIcOWo1gqZWQncxLv0WQ5QvCiPNFPupGtRqRMILeWompRI9l
05idXsNkU6ZX/Wh+FVgY2QtpoS6vRNWspZ1cmJXNXAuNDXhxudfx0z0afK2AGK+u
mYo910nW6s+OxyihQ8fgZpv3HEV2FtthXWCgXm4uHgdsJRZhl/0b59b/Tt2jtRcE
qg3iaZpYM8QVXSFv1NxljwHMdkcbUz+PXUbTo3+jX09VI9oaqTXqhP5/c/EBK8rA
y+wkJ4V/9kRWomntgFbgrJPxLX1mSRl0uIB1HRak/hqBlrLwkV0gihAuQtr9riKf
CyV2F5JooVJV/xXPdhl0VuwoktNdNyibBp/2xIZLSo1bXexTBFFmrX8VR2pfLlS8
LtNkCdzKCrwdr4Vr5+Xky3yWX85SVjAryRKsRLZ3hBjPqk8gv5/Ey9FotZ6kWg63
YkNTJ6GLGdmyamEaP0YaZGIrrF4VMZXB5n3qlocfssDWvXLiq5HkCCLkYp3RKcSI
CeLzoxM/qIlmoVfE/1IH/Q6C1Ovvxq9wQJnkCl0CTKixynHBdf0sEWvTU4kvnctY
iycadice31Ih3yGbqTwGf4tvmmbVvbjXIHne+dPaeI3EPCJ7psFRBr9RNWtwU3oy
lsRJFNp4u//YLkv0/Ms3yd6t4k+puGOKpNFfyGV/KRRilNlZ+Rjc0IA23Ma44zQt
3tfYagl3t20+9hYEyakcVVJqbWZN15C0Z0qlgCxXnttcQkZckn6QCOdeh/mvwHxG
PgxdUu3WD5RSY5vMQ8xJhsq2G9Ctg5GhRZ6tzqJtOX1OvNhTd047d441meTUpkGY
1Q5wpE1l1aihQ87CBYUyTDImJ/sbIhEdwPVrTFu4jr1YoxASreSI636ZR2VoIRW6
tpOdk03sLxXZrfxdjQ1tonOSNI4+GtoQpshm+L7zrpWib6bPSpYmj5XK4FiuHJ3Q
pKeOSX50k9we8YvL5RX+jSkih4qEOgVZZu4LB+S508m3kUxwNb5LJgyjy/HeyC0h
NW0DGNbbRAO58wkBQ8K1KaLQg7YouHpem8XFhTLz9RfRtwOjXkRRM2+QucrkFPau
gvkVEPL78xVtFpzpPYQnPVxOxCB0o6Pc/ZZRElVHatnl6GKADCQVzH75pedZurfX
PjxP+eDQIX56USXblqahJeCpWTlbiqfxhlFPlmdQVecRXsfZJtL69A+hgmc6qHD0
kdTZVIO6bqaqyo4HfXQLUT+/gZQD1X2or8GvCUFaWaPrdpUlSBEDqPaudQZfqFpY
meUx4GROln6TKoVvJuB2v9+ugjUoAnoNgfULBxfZbOCd4CjCL7cvMULt7RHzejx1
HR6RoXCiqDFU8Xi9FPJxlfGPdtlwLEsadeWm9D+ZhmHR5jHWG54RYIN3woUiN0Zd
/+szDANOzwUiVkXJKOLs6T2ghDDuhi8nFFYjKPmkTb3kduWxZKNbfav0cst8JrjU
d5uVUS8RDhj3HzXh1XWzk5Ql1y24inYj5r9sF20Jq9uhfVv7JMuscQQ5x0Gpq61c
Nfd5VEsP7I021iU1rXjwGE03NUaNFj+ATAaSQJwS1ndhThcAlGYbD0mrTYScNhPs
xdykFadkM0Zx2BxIu8YEomlYGH8KI1gTMpeUUV8PHaPQaicULJkLfr6U9DKHksMF
J8gdIvSSWwLe8vUmJSvNZqw6NbhzUUHJ2+pzJqpdGjZW9Vn5NVseWsG3Frr9oaFV
hZTjdRoPjQrtQrw6H+gO0Wz+P2bsBGJLFS/anE+2RQwdTwhfT4H6AKkj7fUzQuYN
erHRbYAdf8BfvyRvfXxx+MRf/KC7f9355IXQojMX/ggz82qlL0A74eZxL0lCyRtC
xA7SnZSZSSGHG1bBtA2OnpNqKKLvsOTtO+JUbTQBP2a8RAgQfCBApVEOPGcpUAjG
/2sfEy4MJCKipVhvGeyiIu7ZO6MCfXtWb6RfqX7hmbkNvWBAQjuecIahQOdCheIg
8msetKwCpnQ0aag1Q7l+JW0ZzVAjfUuVtLKhLzPY0GQk2htvZSML946ygamECCBi
xYhY+FMNHTUcy8ExkcUvFmXpjtO/haN+zD+RxJrTbnimyWuB2DV+vtwfrdq5CTfd
ZFF0CEQw10Tp1LhX9wtCCGDx3kpNsHUrceRJBsWFQwgVPrtBlXO+oPbVJgDPtpu2
9E7VLbolimJiwuEges91piH8LoC0pIp5gZcD+/ELTFuYpHaY4xrJ5cDTgcsHoYbK
P34GLz12p2yV8+r0hG/Vf7HS31u6PI2C64zuIKwgePApo18Grh1pFS+queGtIzaZ
UEGyIzDRIOj8Izkfe/8uZ5n5Y+fYN+khENzJYCMhRzRkH23ikABlB1LThrwsGBa6
rP9fiXfFfkVZ8OYtTCRp3dJI/lR/eahcIwWamVY3wR28xqlYw9hHfzMTxMy6ZC46
kE3O2w7n/WQ+Pl2gn04+7dMb/wNOY9UutsUR8BrXWS/nD6u5d2m1bqW+i3I0KchB
rSLMxF8a5hIm8KUQoyHUFnQcX+rKa6r4ryzP2zevtQ9LeHXgMzBiHu2t1sNQuFsa
uxvZtvMIDvAhVatrd/4KzOoU6ZPHZfIJR4May/on3xrRpVCcIHIfvIghmbevEG0N
eE0sWHRcO6T6GxumroTrcoYZuAhKHtQCCA1jRMLhVvwL/mDB5ZyNJkW1trolAkkS
FnD7Nth4IfdcEd0Ph666qxp2+LqDb1Stlbak3wVeM0BeJ/Gqvg+CyDsyt5CojgEt
/94L4cfcBUXIdrRKfi5Uq9Xi1exJrvChr+wJn5iJRi9D05y7MK8gq4SkT8bbe+hi
gV0jRodUoTb3nGESB7fxqqREZPwztkXMshWUQhpzmM/AtaEluX6vqXrdrSuG830s
weRoNLoAtuHacuSmaplBhmsG/hM8pQvOR7HvgXuCzRO6BjjW/sP+MCAgM7Axr9Rc
wmzK7IzWsiizXGXa107jIjxe+dOF2goqxq0Vu1b202IFKbZt8IVFQ7Re7RQbiX61
KHXjvEPXv3dpncOjxkMC4+DPj1Pq5XCXio+mOY/QbXz+4mcdeAIRTh112hoYJSvF
OQ2Y7B/r8r4jQW14c9zLI++zSPB/F+EyPxMaNIqNiqPoWB/PNFX/KiUeu+oynC+g
LPVholXsWD9o6SenG9zp9Anot7u2mTCcKDLr/vI09MxyxcKC15vYZBeA4tOCuhac
8AsB3YjFGh8PqHpssA9qw1A3x+fVCIgWYQoD6jSa/SpLqIJ+AVDiIMxhMEE2++Fm
DsnQoVT/jc/spkaJvbf0O60OiKNQsdNEOMep2w5/ZK/wYX/BNSvTngboSqpGrcZo
8m2zDaeepNeOKZRYa7ZIUof/Dpuy5UavPW//Cv77iJoNqub9+DElQonU15P8WMwb
RW0pr9rfp0pswQNnW4X7We2EQ826aFOJKXUJvDBost2IARMlMQlmBE1+Q+CGriaD
/X994FL11D0n6ElsFoxkPgVjz/0yU5VDP3vkGrgeHqaFubvEHGfj4SSNMETkHL2G
Dg61tN9k8jJilnOqlpsZDuSGyQNrb7XqWW2CZi9nCNWNKB/Yd4YNAFWUR2gQ98k4
Ah/gXjPcCj5q75OPnPm9qj9IQZfPZGFMqS4k+g94/ES3MnSbvrzBqyJeQsRjhnfg
XMwBxgEwcmSqqmvbRKuLX112jnd6i50lqODKv8WrX285tKFPh3eAOjdlkgvSB50t
YrIKBKqap2NyNghxAjRC9HP05MpQ2HwHKHfACRMzKR8Sun9scJ5pHXyNDTP9trxC
1/b/+et0v2iqgw8wSi7ELZEG4CsclCBq6F+T2lzb+CsfJO2Dtoy+P2MxJg1OeUQH
jb6lUoImPyEkeCmdbb0F7Rb6DU19JqDfONflyfuKrDVmHl1VxgDUGp8crGuyBzNL
IIADhlj13qCSs7MvblMs8Dj2xEuw+lmRDq47wFz7P4MjItX670TPlyuT/FixRwc8
pDHYlkDmm1MjqonymaLmvMSwp2vq4arW0pUA8bhiRD3KOBqEnnAWzqNeNm/9r4pq
aSigfXN5G1IOBJRMOCE1qEqC69tVYl6mxRsgssAOWGbwjoEVTWS41HvtWs2WTTGr
NzXA6mDGTre1dfdH0eOWipJmDxylbGy6fqucNVK3jfbw5D0eYj2F0Urw2BAf7kxz
8rdxQ6eyI5UICS1dOxqX5iNDQpPqlf7rK46LPfiLgJjiskh2QERNNkUUn6CbAn3y
sqeQJXOAdEslhj9MBO3eZ4bUThJGg8QY5FNRGtQrAF0Z8zp1PUi5Pl9Zfpnf7MoX
EAuCXLHg3uKmozN3zkqVzqhUVHD3NeqPjodHp5qgFpGPzZukRnmo/p7u3Zxp0PJ0
9/X4akoLQa/Lkxr4Mju0h/+ymAvbMIwcujwwV99Ed6Ye1FHfOVlmhPsbDUFaZUVh
OeYa4rsoRdoEIf4B1rQi9s88PN+aRe5BlaW09zSN4w/AVHtZErjl5OJrLP6himwW
LfB/HeTMIGYRAeKld9e7gkKgp/WDazfRA/3fs+Qbh1BRyPj/85skNN8zzBmLMhsn
eqjjHYegbrqg+y7n9hlZ7XprnWiCyJt7dCRsBakhk+H/smc33uqyvLp7vtjlQtnz
VxdSMM/PfsqsVTHYSQy39O6YzHj4F3mZEe1e3nmppUpPaUliOggTPj31bxNN07Qa
UO065V4I2BjU9Y9lpPDrMHa2aQ+y/xdXWZkYblvMEO6WtUM4SztCw5fd/kNGBnmy
7au1FtLyt8o6aXrjKvv+LTTw3v0cnIk+VeF0cnpMc+XtVOvZkq26cx95ym+C10fu
yIp43xGH2D9Awpu2K72mv87hSa6F+hmCYFkXeUlxlAAa2EUDsRBdHSZrgLhDJfkq
BqYjC7Sr58/JuniUmLrDr3a440btczkR0+ws3+1lqZmgldMq6lktzpq16kzO12lE
4IwkgXeyfXIsqvoRlT+Vaqc6XYSK+m7uKGf7FGj1+dnJ3/HoSt4SJrxf9DqJDHyV
SY9SiEqIBwm+nZZmtCILE/esoQl2jl+keqoX+dh7RZg4AClIqwzT89+2qoSwAcgL
MB894sui2+359MGiES8hgwhu6AJ/avAD7vv6AKNJR551pGABFrzx0u20Xrk7IJXP
D8Qb+hmcQM7hbB/bsZl5p9rrRvABnDvs/U8x09/cr9zX1kfkiMj2maHujPcIGYqD
YlCKgXgDiG40BlIfmkV4/5AWeT+pbyWsqLcnKOSfWvYF2dAxqw0ZoFr5WUD0GLM1
kBORMtcvTIMaZQaKFYIndqKkMxskSpIKiBvSpwfMutonbKP9X3MKEZimn6mO5e/L
xatbZMnW7C3CXggwa8ZAPwBJRtFM1KaHhF4veJz7E9YrFe4NhHhJrZuKnee4CJG3
R38rMFfvLKgMd8/d1RWnTI2xx0oB9adjgCYYhyCBdDYbXGvYDT1r+0dk7LbuR47P
PFXSQ+jAi6jZdP3wFv3mS6F1ZxVDJEJbXgrJA3kyiGtUDzbbmsHLmbZGK20C0E36
XNoSfFaIgRmCEt8KV1jImRMk4hdrJcDUAjdyC+x6F7GN8D3dQXnn4fo1TG1EqFKe
gAT/xlpEIU9PYs8ViNy8J5RvcHMZ+LHyVYDyqgws9OsS933O0UVJuBF0GILDxdPv
hMeiVi+r3XZ27fK3MUtrOYb/MuAgS3Xereo0WS9U/u1dnZUY4smMs/PdMNhLWIAC
ZJPPgP9yu2/fXHbJLw3tpNNZiGwQ/3lG/dvuPavb5urLOeaMq/C2lEa896v0OenJ
yefYEcDwhxKjzb/LcikHbbsl1LqirRxcYp8num+QN9bnYqJ0eDPDCALOltWy07dv
g4+j5RGbvQ6sNfnrXAD1CGA9QC9NKuPUjbPy4tSZCoeAGmKg2NHcD33jKEjGXF6D
egPn90GyWtb9as0nrfobB1Qy9XVC3SiXUktJaXnKJs7Ui8tt+F/xnCvIjRki2qms
VN5NfFEpK0hxcsoWqYWEpnu8fZbv9+ZgZUWm+S/sM8/j6BEvSYVvtgOepv+gvXSX
6b6z8pmTU4yMP8aMp61q1EZ6D5VMUg9wbpTtifeTTCxrIjEVh5Xd3E+oT7So3KHW
oeyjhnYjdlisEO2A3dRcTWxqz86MfVc3qRH00RLVpj++vNPhkHFNeyDlRXOUuvqN
ar5h99mv6egRSX+dbOnbTdu7MxFyy8O/xVK+bg3ofUU3hGmwBs4m8/UGbTR+lJmw
Mql4sNdqulbvm6BlpNsUN5RPs1uvUAzfO62Y0/VWNuBo7jHR3dR5k53B4HleFYzF
b5M24mbp6zROLqPgMxTUQF0ADldqlaZGMUNT8nidf3pZNKoNXTHl1j2iTodfErEe
6OGOLeng5RPnmXuHl8iuhbkQeziPm1ZWWVAjPc2YbfqlqB4VUQm5iq2M1coTOxNr
KJgnBDJK1eKlExt38CR8TX6vmcXN7oWKFlc2L68pDb3S8hU0sNwb0zx9nQ9q1/Gv
jmAtctpa8k3PgPNiZYgi3Fq/nVXSabkQSuYN29fr1mD7wdN//Z7hdC8Jhj3mozWf
zud2ueOL/wCDZA84c4vQ2CVlaD4H34QmeQatkGRibdNzO1TNob+h/GncpRO7QPG3
8IdZFZrfICRbelP2tjtXgFhQzH5JrufDTWEMejt/2WYjhIUxMa6o1ahf/N1p5/Hj
3cJW8SttMpRj4lE3ERxnVqpfDvXCpqDDS+vPhwim6JKLbBFmGl3P9w3c3WpIMSGM
IiVmIcgYM+6LN0X796g83xvVY1WXsELdE/oC/B/ncp1lTCCQ0JCnqlPX+F/VsrIO
HzO2lcssNsUKfjA4Rotljy7VBl/p+bO9rIdESVhriiDe71/nu9eBrPv9WznOJ0P0
bD98GpNaDcBO6dEkdqw2ENx8giCmEyYszVLlkoveWIm2Ffvh53rKXsbYIKhYq3M1
K51fQP8i6aXCwtPca10hQ9VqWnXkeerqDqsLkKqFvdbBEr68oFxwEGFA8dsunKLD
edtDwPQfeGj6vduosWptCmOZ9VvPTS98PBBxF4/vAg9LzKydD+ZqcU1EpJBUix5x
6rOZjWWIUIQqI/OnAUbQH5vFrl52/5FSoGL+4VjGKiUJVAvAseHWaai4bO+opYZ7
y7rhmi41aJBnVVTOFbo8eAjd7sdLLZH1pAQa5H2kwIJIJ7s42x6idD36fptVTqC9
P3WnNX+TzEmluce/3waJ/WNi13gi3xjzyzNA5dKrNxehle1Io38FK13abnmWZ90W
yv/1JUwY0DRUFmPC4GlGGCn4QC7w6oXc0c8V1vi3YYR9MWCXH2JOGK+gJ1rJUVDd
r1B8XI+38Gih0LK4jpmHs3dSBsXIZrtvNC+wJ3R9eqZrDQS2ikhBPnaRAA+WL42s
vWtye2w0whooht7XuczhjhMg2H+gAoICmksE/cmOj0i4Scgsldkx5RnhuVQ4SSsR
UUTtKqPdqUjuug8aHc6yaoSlZrnBriJB1SbY/E1HlFGH1Q01/FLJfhRkx3u2Arn9
QHcwCATPufOLFKfFBuljjoBrYWVBLFnH1tRYvUrslgMm5n8vtEWXlLGF2Jb0wvaI
Nl1N3eqPYgd9qDh3VROByNr9qilmYSZkbKCCa4fPiQ85u0VNkg6TEJ2OcKhcGjsg
i/IsqRrxR3VBhaTV37EQOqr/dhCS/r/fBK5+kbOYgde8oEPuu+jdI9vpqIJU9tQP
LQ92BJ0tQcVoH/3Fb64qeREPnGhQhXgZQ+f0d/Z6ibmjqu2wFoodN9bNj+1GYIV2
8bc1tPl0205E0K2VoONJD4rCw9ACgtNZuPl9bb+F7qT5b3bjQ+4d7S/vJ3ya2H97
f1RYRS7BUESYh1tUI8iGsBieOOEkzR2ToeGhwgXbB+r9Q87sVzhiIVOJXvrWDJGG
8053d2HK3YLzEOKvi0r1YX6oyBlsvpayRcojTO4WZ0hrTkD1wUlWwrSXwBoHsCCN
F7nGurVWFkt3okJ9OA32iQyGcRabCA7fhXsFi1CfkSZGSS1UF9ZAMkoAxQauwtcI
5/IvGSeOtAgFHAfl705qcKp6iKZUSzbeyWMSUPk9phmqoyKLMN00OtJssVaUp7DF
H7aTAadFR71OI307UcXXeumODAZByprMeT5AZnBcZ8Jfdb/N9vbTfl9HcJfXfn5p
pFlpdwE5iB+jvQS5sZZ74iaci66V4Ko8EOXr+Cyv9wzmha8X3yv28MxWboTTpzAC
w4GMESVILagsJ+hOeORbaKxrRmUNlccgUXNQpcYjfJend1JBbMGx1sMPTRE3U8Z5
StDA7pATvE7x2ckxlXmgb+bJ0XfpISREq/yxTATTHhJuTNPeSSHY49tHh4lhrKFy
OX6lCKlW22vcbEy6/qaCLoC+uUShCRfHo7e4zasjdbz0rxJaKOz/qi2841hURyN9
n7od8d7N9ak8Syc8qLtCTdDIJUXXecfopQ73R+f5NbOOpkmC1MxxGIWjekAAo2VJ
W7QT8uIEBDDR4dQkLy3C5NEsfl9hW4nnMveRoNnZttxqO5mtoNxtJCerI+NDWe7U
4x8NsNd7r1z+lNdiM0GW0Q0I19wYbncxjqGjldfUsGjj2syA1KnKoMvDIGDbsBxL
IF70jkq9s1AHSVgW/JS7fhun59P0kD9Z5dhCx1PykNHj1RNTZUCp3oLk8wEUPZO+
CO+Sy8189EWeNMPZ/UHKNuAWxRzU/ErBCn9fXWgOJmdlzdTB4jehzTYpbdGQCECG
pwvhJaHXYr+vzf5Wt06qBYxm9k71rj1q0LiKE483OTdqKsOsM1KHQEeUBwM7jxi9
ccdGERS8lw/Ai0ntTGOmrF1Jz3KMNb0OK9Zh9ebyljM+IQBOwIukXq/7n1g2VIGs
K9WQQJtDKUwdGZT6OLV7ffr5aQ51oqaJZpbJtASfKkDRSWIywXE4XQIGVDeK4tjd
7C5FW/qbxufNLIVqTPm4qtijP/pzx2Xz2ivFIyEdb3jDXc+aJ5UHCXLP1mpLOzAI
nf0JfiGFldg4UmdP8B3jjQqgfq0L/AjzV9+QWfoy41d8XzbkazWWU9gVDpzwR8Wo
YYefJsUBBVjQ8d+WAXke01ek53V6vWbn1EfZuejRo9ZJ8frRrJxSlwSIw6kRQf04
yi/hrV3T1z5m0n0OiqVoXNut+MGuhufiOaixzFq7Sgqf/bBBybzJTA6TI649hO2D
X8dZmUMC0IS0K9dmMnrY7iuTo3bFruXwAqLUVt6vICFosJoA6mqw4k0hHNk9P7R6
Okx0V+zsXgABh+CL3BT0WU34Yrin82w2EPO7uGDey5XNgjC7B/LZNH/j6AbtB6rg
VGEBIbZliwil84MUVkWruPDtEMkdFT2qfdAHbo4xh8pGZZQxbtDfyabXdZIxIRYp
WPzTaSZ4uCrgzcbGAF/9unAWHzsF+WNszFlPUoPzkjdy9PXTnIkdy5BsAlt9qdrM
PC/zNRTnd4zlK02+QOUKLzyVJG0SK34VfyAH2fQZ2XR2MKGbyI2kjV2flNGS/LLx
zBaNs9TSlCf5vIi1eCwReOqGpklxjgDQmzKsRAXO91hyuXiPhBg1rbJe80N0hBZH
JB0Y1aclhpw/lYgq3CSUFMt67wviX4xoP4dyx5W2cbjkC2wgFAoqj09qAfS/yzXP
k7drvY/CerERPnOOmLfDmamP1mfOnvTKmJZpf4AmMa0LoW7VoZcAP4jV3H4SaHAI
Npunsl2PK8YudHUTcplIJGXBv5XxLFr/tvnE9iK4SlIDsSOLD6qzhQHrraZTMFNI
bsaMIX1YyAJz0AbCxnrzesl1oMVyFaZVTtZIyan1S16U09ALMbDxmm5oaZW4kNzN
5EPWxj7nVFUOx6JXxQ81pGzOUYrn/gioHI3fYe/GIxEINXWQMQRNNjYJj9WZe71J
xgjny3BqXLsz/iw+bQut21g9rmaXkAjWERssdYd3UDUNxMG4dGu7eL0O7SwPtetJ
LXpma5QJ3LxfWxeYljziLDlrgyTrH4Za/6qnixm8ByGa8bb4ZSyEor93LfF2CK0+
TtSYe1L1pzNK0YHjE4F9Gl5Q7Kj8G++QPO3nxYwgrrFTyWOmhABJGZIHGVmbyiAQ
xpjxOOBLKDzRb/javr3EAEkgiNqy+Z5p31v6ukZFhMbxLw34lRo6jrxz7Y83V/67
/7vuNPsuW/3JAWsmcqJmSISap3vdo6c/KadYZebz22UuKn2OeVM4uKDuQeSSS2LQ
WeWgLKkl5V+dnnX+dcjNbDoZr2osV8AyCmKK+cyOM3X9rq0Z6VC6tKvPof6mn8I2
JWg509iFW52Th+ChYw09dXB6i0BojGFM7LChAAACcRlbrwycBT6RVdNVDBh6fj7q
ygFWNxwlVa7Rw4ng42o4k0+wxkWgOwrkzKMcfAgZ0M2T6KNfl5UIynjR8szZwo6n
ByzSZsZmIVTX30gHF3xIBXXoUwctFGIdOAfZzww6C8AYFSpFHxDEQJXw0+R9d9Ka
Q/kLoxRrgvWguDlyygXJczNbd+KTi29iLICx5b3uy/umTGIqF/s/RPMzAi5/YgJa
1KfyRSu0Bc5ITrwlrKB9nstN3+2AtK7RjmHjIS1kSfgFfMAORnC4EWqCeq6OoR7j
gXBIhhzPx+PDiWazNUvzQ+bYnvPbJj8lDU3mN3yhg4rSxb0xK66VZywu/ltcby2E
9/P4vtMwsZ3aFmR/+3u9KFY6GGccBpd7fWW8xR+tQeKWXAz3IXseOo0ulF9ByCgP
c/uRoa+1h8G7Wo2ndh3Ih3yUNBPZQXYctYOBBcsxg3ep0JwhEIog7lklvSFmk72u
q9qf/BJ1FfU4mYuXkqx/gxNblU8Se3XYYwjBmi+BaBLDsX5wnbN2V4acJ13q57Xn
VwfSOUcqJppUsQTr+DHUcZS0C/bGdIcL3AvuBdkJHX/dunmoIbXbvtxDhJ2SIrYN
GjnvAFt6ctNmxfywXpjTZvHgGwtX7eNUUErqnX3Yp/XwBZ3YjBDVhAUIIsWYXf/m
4JLgiqCpALoxpz/nKEs8Uzfs5kbCQJPUm6ZvtTECGYCI7rgoCDPP2uuMUlkRFR1D
Yae+Z/IbhboB+ntVyKMOGcDMqgjUNCBefGOYQfc/GgRjgydpAZ/DDbHQ7szTsTJX
ix6I20rnEuIfpOjiPUvB4/gmWw+of8V4Nc0Z927WxO3XVZj4eI9HQ1s1UEck2RRx
H+8BId/p+tV9ZhHX4rcTBwNHjslZXKiGN01SNz32Yx+ujKaxLiLOjBKe3wZZM1Gg
YuhaZDfWgC+MvemPX+lwMABnVg3LBotoViLFFgmezXErIyRAkLMwpmbubVUTKiBK
ABfROyOZZdb4IhM6z7hS27mxwfeN4iArlY8bbIXpF1S2sWP+oCKzjEGMD/b2oMd/
6/fNoaGejANXgAf+VJS4IKhN/MkSCZfBG5ug9EfyWQkWwpXHHuoRxDC2e7a+RRC/
3+Ro9jvOMqet9J3wp94FhsyFIV6lPJDZNzMXEGFzk5oATo5RJJWnrpNu984paSsJ
BNEMEW60IQPojvwetBUFa5jFZMBY7J/645evlZJe5ILC98GwlvQkl/BP5aE9Xgbc
cbxXOxdbO6aP8/tLg7+4GXp+h/T/++HrbawzAsKZDAVVrYdfR8zH9fcxLqTXKZET
ZEG3Se18i1gYoiKN1xarGLemJ0dUDrzyKDkhgisHcikhJ/ggraQFgaODaXJNZGxW
2CVjjnmJRuC0ZdMrVWnwyLozTS2GVMv9GuDyOq0IDLM1HoNKxerPm/Bgmeo5icuE
X7UJN0ocAvnX5qM6aFPq3r3X0WNGxenqawC0toAovwWkELykiMRQ/qNI6Lcvo+jx
ZyNC8Axz+I442Mpjgbq9atN6H0cX9cqaSQYp1+MxJc3veT82xnkN3L4XVccC6G8b
FIa6rnrgXGtaXf0XzmWCkknhp/MK7TVuqNKMOLNmSZ1aP6CbA1BegjcxgXn3OWIw
IaemHmWXtgOvNe9E2nueIigY1ojRqdaHfuXceLx1esFzeI/fnvDdJgqaA314uxHE
zVpOHDueKXEApWF7HnODDtyhgih/cKzfzsGlPuO0VbxapITNOeJMleCGyHC9tFem
4Xk/Eo5s6+GweviYHLlfNkhq0lu3weI2TVb1B1QUHJs9vaf569Xa7r4TvXHJJo3q
JiP8HR8YZv7osTF3ROt54iqOO246OAExrMRrVQk+yBNvJBTCZHiToXqKJJKstNy/
+zRyZajc12wQSwBe5jItTW1kaF9JgfRM4fj6JnDu8DHZNoeKfk4lDxtHf3a8RH9B
qBiw0Y4ajv0rxSj5rvXRwJ3+NvpU6Hen+Mz+LZkLmVuhlRZQFXIsX1k5YFaUaUNm
rEl2rlJBLGaNCiafhcdr+t3huO8aiCFYnfflynYlwjPZfXJPfOWnt6523Eg9hIR2
mndtwzFL/F4F9c4ej1IabIqEhdMrDrTxUtQQlL6dLP7IzGNbkDrYx315wXLnPXzt
Hk02MDEHzkn+e2TKED61xNR3UfvWwC0FjYw5x1k5FCgnihx6X6yDNGWsK66Bvd+D
IoRJYzJAmLXRn+k3y178w6szLOUu7qcqXdOuBxQNxRmdSGpakaWWaZAymZ092Dki
rOrIiLN5RrFi3trH6Ap/mCtESkoVX43deVR6z9FcMwFBmiUc05EcSTQ0VbF2jd+r
FkEVkiXh8WNCswXIlFMY35EV817m9h0I0l3mtB89W/kG51Q0QDXE4jsF9PrBgdWX
n/7KSO+YCnNTL7IEB/pEzsQBKcTGAN3o8UV1xMZoiuFTJUUK8bo1pehozGW7yFq4
4j5s4Tsyu6C5z5Uqs/EkhFJrz++GIOCPQY0+J8tqwyW+k1HTP/Q28VQUFVgz3G3h
5bgpPYmNvUwZrqNf7Ubfjvu0p0y8rlS+RESshJZrIgmEhm7NJJqHQ0w5vfHydnUK
MqCsPjD2lNydxhwzop28lE3D6nn8QKvwdDhelE0wnqIwV2UOg6PRXA0J7R49jrC6
BHbsec8qCQ3rGd5FkIHnHx+X3/UsIUKdacF0ucz7TLIDVKt2MqB2AzaXXnjKz/vb
7BfmCFLKP9oPNpOHMDEs+PAmTEqY9rokVkgn2H8+E9pkt0rPCajAOznvU8SLHKiU
J+/k1rZt/fKQO0Q7LiFL7dTSCyL9DokquO/M+OUWyKvaya11knPQAPBtOHknEV7C
x0dDjvvy2Wm9OiKZ8VT6wPXNvUyW2Fv0Hb7AZbZwz2PxBk3YWeypFIUFSAlD84bS
p0l6NCBscuUm2gcLdxccLr8STtYBsTRpdWQtHvloDSNbpiKofpvDnHEDBdbp07zY
t6aOC2N7uBkjdpPJtD5p1DcyNX9SmML14A2NmpbN/tjFu4DWVCNWqO6Ew9359Bca
uw1r8l2QKqJzeq0QVDyOP9j9VC2NTD/tcgtp7v8n+fYZfYlYIr8xzoXfhS/CMxGl
nCSPcfLKRD/+8dF0jgsRt/VYpqftTz/y++PLnBAdia4vY79nJtfO4XvGllNNP7FQ
SHOhcU4xO02ZWYIxhIyQ6nBlCOk6a2xKeY01F+YMBOxk1nI/rzQBPaCvJYyMfTS0
R6h+12/6u4Z9tko58pu0aTv562yiMxKsj7vJnY/bUh9zRnOAt5GpLB4DOsR4Sbta
nB3E9b56yOTAM4qx7OJRhhpxcEkoOUhnTEurF9sTgzcGylECK01r4YuMnWcKJNKS
Az27RqgW3EU9+R5xYAIcJzNonizdt5o6mY+3uFK1OuSgZqRhdKb3RCRLY3yac9+9
I/YyTizDt/2X8VljVTvtI7UZXUOhsYbC5PTUJEHaHCVkVATDrrTkC2aqweeMwwE2
Sh676gwIqMHWAR2aJpHFZeHbfYHDAN/zlcUjOXaOZjonTX/ZdafSKjh5hXhuVmd9
XsQBLwJnNBW6WM0B8GYzhV67vv6SqWgRF0l0lRY16h7nZiqPjm77VXU+cmjW8UTb
OqQQ/E3A8w4dASPC03NwrIoz7C0VIChCe7muKgpYZR9qV+5CUOMjjfhyRpIgUS8b
yoO3bMVcBJLkvx5H4rebD6UzvKYzDNCqzK36AYVR7EFdyIzWKX6oz47whSUJymEC
q9dYMn1ax+EWYDOKgpp+YftKHk2IGwYVLM+3Pc02nDsvdMXhMB6IUWjNSN6ehmnq
EpHPRAKl/HNf/o/2JAzK6MgV0necWbAvRbPHDnYD2VQ2Q8DUWyO4MuhmH/W9Pz5s
ZDTgYOWSorUIG4hHPDexvlbOG2dufvEFARmFGJHX5JRHnbPngAd88sllIOH5Qp9t
5f6XgMKFLo51f8LVsWhr+xevPB6QUYxU8P5aMLzjeqh0MayhUFp4HIiGKSSnawGn
4j5oX/e6iBMFVTQqd44N3AskcYpQug7E/hzqp2GGppMGOrjFdx6ypQeFBab+XCyV
6mGRfAskEk56YfyMx40p+xeSf6B6f7s8zj39/nNZcF+yv9xs6fZQBrx+HKsbfNiT
G4lvNB67d/AFninfUQtLXnvT75ap6ICpnVvShRY5apxao9jbtVpLesSNeCYxeCdM
zTph1LDAmMRj+66Upce+8OqKFd5gc5lGoCOr90b70K2tKoTGSPwfMqzsJrsSjzSE
Z1ZdqjNmSOjQP3oxf1VselbW6fnfgOJf1hpPeUsjTXvQZaVenNDYEx4WEiVg1+rW
VMSFImOeV5Yhgh0hqAGG0DFInu9bk3+qX3qCo9p/PS+p5WOxl3VEz5UcwqUNtUhq
bi5oZdEkHOzAaJwpoVVq9UirnkDUUQOZKu4N3ijVxynHCZXa7flAhCZT3deQIw+7
qXDb7TK83fMws6r6+OcW8vQtZkHo2qWkUIdcNDRP9jQS9L6Vq0eRIVE1GlQDcrLy
J4BTg/DkDpcY0HcW023ZiO02F00ZCqtXCZkUgRlHpgaoXGAwOj1iNu1SzOMPVF3a
8riS8bpBlAHZsZtOgbvoJqeP4YFSzGvNwKh8Akj01laVD/HwN0VRM1m4Jc5vaLwW
Aka9Jh0TRdcqvcYtmFOTaFzBaSqOcbifWcPMU6uk5wS7dyMDUWl0mOtsBPgWJktU
kciBpjMcPhRtiC665PlHvAHLX1rJc2Zjsa/uSRixrU3xX+CcD6fA1oPR1BmWE46n
SUWG4RUYFBrE2C/LIyobFlNLtBLhbCkehYuN4oV0erW4fSiyXfyYxRXmJnGvu7r4
ECyI2HNWfT8GcGYhOGCPbuEo9IAlarHCWJeyrzHWfTKNzxspkhxII1VJrfh/a0w4
xM5aKHCkiIieI3FuqDfmrrZDmZXu4wD8n+Qr2Om4Q5sUlpogA6uWXzwNkT7Mdiwy
DF8qJ+A4h/ae4kf9dqH8/1hTVjztO4XIRV8CXiYW+xfjucLIbeuClmGqbhS2+5yw
zkFJuRheHFWVCxYbtqAKqxPaPIp8/MW3pjBO98C/dR8qCLd4GrIC3pmJAxeAlK4P
dpObCdrVh+LGzFJPuzEDQ1fRPbHzyfIasR0mGLykmNWjrVe4gNrWf5zslkUvAgVA
dHu01GuKrvptKZOOHSqPPfYTZl7piK7edBkG9A59ER9LzYbrsmwtyolgOrbfnBXP
vhhj3a3hgN0xa94n7J4knQKlR1nQSW4cap4ADrant17WyZ619E7CS8jMWW3Rcd87
zpc/3Hj6kDtaXkUurUq+2O5eQMF/Jxim6B8rKjMKbIsIo/w/ON+9ihMDEwEk4ul/
bT/xIEWDRMCsk2p+YEEAGkSgvCNd2BZA/NUGmoZuMJnZQ/wdy6qN1C8CR5V9yFr0
PIGQ7iDRhkg+VYwRHrEjF15S3V2HXtwsy4jGPaxLm5snNiFoZYLsgsPuOd0IXBIp
sClbnIWy/5xaDhzCHWvb0MfX6M9uhYYcTRpWaSQyU6GB/NY9zs4BzWnhMy/PfAPM
PP7l5LDxzqG80A4woCa1l/WvUuAh7VK+ctOVE8EhPKjgD9Eq0/0/+Cx+MbWMN2e3
os1TwCnyXnkKXj3lIK+korDS2hHGIFnsL/8wP9nb4goNmkcpjy5HIHRXLHJ6uUNP
Ta3iI23KVP9/JnLeSlpuQ/nJlnzOCkNoOJP4wiA+ulPXG8B/45YRUG8CK2gClH+5
Wlq7PZFarE5cbjtWyKrAr1uq5ZHklZuT3jra/5HqR52IJ7JO46DpHBaZxKIYFPIL
1p5b0way+8HICJAXiEP5ILjBqKBQDum7sk/4/uXiKn/SjMP9cf13q85mudEeEM10
bMMGefYi8jpXC8hhLeKSbVC35ttI2uixlFFSae5sxlOf8Uto/cTcUTbjGgEgQ76j
514AA5NN1Yf1XM6e/rO0O/ADczN1DbgdR79mv4JiLrhR3UZO/pK9yeG6C6rpGwr/
cQ6A4/1c5ddqKwkLfcg85l1UD1gQSicV0h2KH2M+Mo0Kf0ONRIZnZUsDPDXQL6Ox
1+GgV9YZ8QOYWGEWuNuosP82henAn1VjSlSFj+1sum6L42GImqyg11ESkiTyQU0B
z8JtvTf1tsx0pJuyUz7rAvByZGoMkSCQjOJ5YEC9NjNLS7QHiFR8PoCysAll7Dmv
dh3Gmdq4Gyd7LrM+4cxYhIlucaO2YIZ16p3niao/n1E2V2Qp/0mc4RC2J3lzwSEY
Qb5ZGlXDq4p/baeNIlisQRWn7FNwfUjQ91gxw9VfOeMriL4GYeROt9UXzKlqUgP8
o13iIB3Nm8TdL47CpCE5q1c9TDlz+ZhG62aSfjkZ3Fl/YzYppgF5GxYk9uldimms
uP9YmmNYoR/DC0KKAir/LmwEyIAlGirCrdsKp0f3lmaGay4YphDmt3Rc1EQmWBIw
tF44EJ7pZENifr9cwNiAj0PbjPJz1jQPr8EzchniF8wwIl+ny9XYyAHNqJHb66Eu
ho45aBIDi2VDBBD0ji353+GVfMmT7kwY9XiPmR9h9hF+c+7jnFCLcxq/UuS/SzT9
XRxy4mklfvcwzoRsq2qGIPHTdiMn2pWyxwPtX610ayqfq3/UEF23XKuja62HMMHW
S47PhRgR0N1WL5+S/N7Y9j+y6uFtwCR80/TiaNsNaaJNBn1Udbx6jIdpzaXwxWs3
J8Vnnb5WYe7J68fvhPBxtA9cb4DAG9VQCMlENBREw8ZWWSuSFfhgQoXJ5uksrABu
G9HRxJF/ArTHMU1kZJZUgHcAvgByTSiMAlYFmGVI5YV+5bOZMmX+0JCztflFo/iX
i8MF/2+l+uAB2hSRwzFqv5hmFQRngPnOHORBXGRuQHRiXFuhteGA0ouNkxtvrNwe
jM3V3IE93YEPmMb13hMQMvOmXEvP/AK7GOhbGi5/n2XjWsjgaWYCnBR4yNkCRjTt
DZ8fZK5LUQv/9cbXA6wD3xQ6oDOCxAo2rfI0sLPeImW8GVzFeEYAXre5tYk8rsa+
iRuvsf90lajHq0q8bDvSrsfuxp4slGKeJ61a8br1dX5ZThOERgf/l2fNVJ7svsTn
rqgRdecU/OEReCuyaHmLGAFX8D0emuZV1vgddfWvm1H2IG3rIoP8SQbl4XIF7NOX
FV7VRB7FqEl/1F1CMcVn508JJ6UjYQE1PdaLs9TZCZMD1V7OiIGUx0BsEWTEYgDW
vH7UMcvs8Vwn7ThccT+Z11a/6ZsuUUFFEZNjtgvqSV7KHCB344Qljf5lN8mgoOJs
axFq7QuT7hnLN62nTGjlz9WDg+QLqcbdZnS0Apa+Nv+VHQ+voq9cJXc594B1ZPYs
HeVMwKvdldyrLomoiPehHdBd7uNCYb817uAB9QW61rRrMZZLotbvrpxWC+4ZxVoM
JC/Ekdss+etjoBhB/9oMv3glGgcN9y4BaDXCK3VskecoOfM/aPF143UTUtzu/g8l
v677fgFfCrnU9Cs9oS8wLlHtumlnAeFEkrKb36e2l7JhlGNm8HCR/ncYB10imZsD
tfwDrtjZf3P/ldCnyJutTtyuR/VWJibit3RzaH41o7c8LykHVa2HX/d00Fn+to/d
kNee7AMksppwHeB7uYngWh5XGCUwUnAoOx9o4pblaEgqOA3UI32LS6t3tf3PmSBP
W5F/3jNz79J9L9fqkwFXidFiX+fycG4u2uU9OEYdmkiEzzf5CdCAMKCgW7mGetXB
atGJhrd0frWQjeC1Pogx6uXjTQeCJTo+CAc8AET6FDcJ+r2p19KHKdnRc+Uomu9D
Sux3C0XNWINhYPmg4yLucw96Uuqivwfmt67Nv+C6S4Nt9b0HBV57X7j7NJ/8LFoW
vNRxdsqkj9JBFjufiEKYM36kVbiYuiMnVw4vhwcVM2QFdvhqTnQeno6NiDBTnmki
q1IwG12zYbtO2jju4WXr6keFLkN/kgE16I71Eb57NkAxpgyEfuPAfsNU4bZ0Y37G
o0UOpDVSwz+SWSrs3IKiBz9yGs3JaX5dWwZUEPcPA2kVD/qB3mkKQdV88Cs4QWPX
J1Mb7M1GhdgK3gtv33RVO8ohYQpiM0BonxQ0Op0nluteT0jddImK9DstuayvQtJ5
/EQG/2rDtbpldl8rbhIZUUVi9Fs4OYDJKAZOvxjhx3zDzeJwDb3JEwakjO8W+0VF
8YEQizqyUOL9+PTtgJyHIfCTScDP2eCgw6NEw2luZxSWcY2SY4zGtjxMIWFJ40lt
vBWVyDqxdus0nwsVDVYEsxDEIiAFU+/3v72uVjzRxCpXY29paSBwVSqDDplKGbM6
P/ZdkN/j3dRJD/zTn+sZgnsmI5yup7yAHLGXP43KENAa42yUIBmnx6q8jC9u+Nhw
z7zXJuUJ/SurA27Fbv5Oq1tHk+TbvusExvr5D1Bpmn4TccZTtwKlJyLvph+BJNe4
b94/HJAiy8VCaiXH9WTdUZj1Q6mKZdTMTLdLukzvxHfBSmbkzmbVIhk1llHRY5/k
BsR+GYapzB0sV336gxEtgRcnZYT9zxSBsesk5SvAER15pvIXVB18WaUhd1vpbBwJ
rgq5NFciEPa28+XNoVaCTxRS4XduDSoZ6n5HD+6/eiA7K0eIdXz0220//R+6IoRj
hQ+Q1sVBs6mNJT7uRcnNt0FvlajMAS2TBlCQNH4t6sgZmIBiSBilPXXyQBuhkh1Q
qfSitiZm0sdFvQ6TTs4A849UBhL4EZZxLb6wWyDa3zotMUB1T/hyz0J9HYY2DuLT
+NBlD0tUhag5CC+yq6kC/TixvWSkrdutnpGVCWVnGZHyJ+egJhKz3z/JA4exseUD
CwFTIRAAVPPtvZDsqe9eRUkdPJmILRjdwQerMpSN3nZiJRZeu1DsLC3IYKq+jbRe
VZOPPthCOPUCa14tFzIsEhwV7uNIA4PYd+3wxK3LTVdDSDx64FXOiriWSGdf1pWl
PlG4E0wZo/L8dDSj6zFvhORWtQTpsyDj6D2ydIdXWZxkRHxgrS43gKJD8ysp3ft/
MvFrlPIo9BL9RwAyUebxf2t9VoWXjgiRBnZ5lOPPze8XWGFX9XSsKPQmW7KMyrIE
8rG26C+3iLQmtQA6vyoXIvGVtL2pRs+oL2rh15LLlQuCPtcJFsEMbfwiotiL3XyD
gGQKI8rV2fJH3BBxUbmzahkWtZhbM7ISBcZ9Ccv2ibn1n6psaOxPg6KPOaJWlPV1
pJp7df4TGdR3aaPszVAvFELJPnSfehl5WlmnRIHva6q63BCygQQto7VXPU9myYqD
6R++bE7U/M3xdma5GxPGq8JnhpO5C/nOkicQp6ZJEmtmbxduxGOqOTGpUlg3gMqq
l+P2IiKOvw1VQZD+xnOFQ27qHIG5AM/Qp5m5xi4P/UCxcznDJpyD0/KcyUTj7boK
BAsrc+OFlz+CAOlIX46NY+dYEM36nDCW1pM1FrVpHGOFbX1euUrh+QrnlP+c7ddA
72SImCa27eWBEv09RFT8AwXX+8oTMTKICya8smRZDRrfgEv0WLysmkjlLhrEvFmo
ZKt5YazLqtPJrfNBaweX5E4NmnPciBPciHGVn31GUkDz5qMA96xkwFoUA/vMVpYD
2LsqPoMMiaCn/wmZ6L2pLafbfeVf+X6GzqUSqq4xQGHXQ0EIv+8QOPi/M2ipiWPR
sqxU6Ep0UL0gjnoAMneumxwyC4N2fEKUTISFJcbqZWpAxJzcdewP6IYA01IFAY8M
qBx3jG97YSNS3kjLRnWZN5Wm1Zke7fQdasoXydl+Oy29G1vMTSKAdvdzFIoygM0o
ER2Y0zCeOdOPm33rlFHvZbbMwcdZlCoOGxC1NEc3m7mempFoH29zP51vgMofWXiL
KIn2e3uoPRUewLasGvCLESmftKODF6oJ5qWDyKaLegLwj7gxr1c23eZa1Os4EeR2
Oej/lZuxTpqY2/eFJGiamErp2NnHYtOHmqUdV/P+cIYivj9k+VJl8VPrqgoUOlu2
Jj3othTTvu7ZKS0SDDQ5MmvEzsVsPvGqle4BrsPzZkGguVa1Grwms7oTjOE3LOE3
fdhVrQZN711HSteriQCbG8I7eGhXTw20sVLydQ06mqCl0tPifxlSzikGf6KWDN56
Am/FyeicEOom31HctCrGGGFzioNPdlB3Rcr1MqJ6klRCmv8btM3jbzmTZ1Qv4RPc
2OlFaV4wY4V5rS3eVIWAT7rA8AFvUjCjBC1X4ffYc4Gbeu2z9I88kaOC9TOZdmWf
jT1dKifuq9q1lcW20rSnL391SiYuDrXMuCHkS0HTouv+66t65IzzXgTeGVWISyYJ
qUcfkW3Am+yLNEsdbGVFtTfKAD9K7wXgWcu8gQq+vKbcJVG0BWaJgpvfbD67t+o+
1rmfD5+MqXR0Zcph4rKtfY0uzeeHVpYq+5q7B07baZAbGzvBR0Jm+6CZRvikQWS6
osmslHjhtb9fcV90EdX+RvBxPHtih0kr5MwRPdKazGAab26EyEMAs1nVLu2saX82
J+PYf/Vwk0a2IhvPNqHJs3zxrIfougYxTfHE5NytXEmhA9SFe1w/bKIsLsxJ8Mhu
/m8b/ElKQ8V0sjz7qs47xgnXz6w67bUxR0PJ7YIn9ttGeOVMdbJ6FB9/HZbauOb/
4gP1hYoWNyrMtGBA2oCb2OQ3J1EJS/M/nNOCEIJrCxZ4Luo2r/vLYxh1oUay2qK9
zldd5GHAD8rUEdj155m+PDckiQ1rNtgapo3119vc/DG0jxtIBtpTvo8B3DgG4EGl
cPDQHRWWExJKmKse2pEUoyFiW95rNpsM+n58oiwRrAf+s8M63U/wibtiGFGsgz0L
5cOvqwlImx8ahGx2MnMjhnuhczDG/LmIfF2UN+9Mk21DvaaDj+O73VQWC4WrjROV
1b3TunPwG0URPYBqZB2/qgBAKh61ETBzQkJ8sRyQrmyfWN0rydx+UIl0IHGe+KYm
illGuri3LzKD9OxX4mNDoAlpHoIQhqDtWclK8Abmc79lIrexhJOvigAqOEe3+5bt
uEuvjq0SrloSitFpxlA0rI27WldrmBGrvUjyXTpQffEaPdVc9SkUmawini38Y8US
H1j5LCPljQldfeCkr2id1mjjPsY1DHSk1bgK6aQiF+VAF2PKZIxuY2KyfoiULOGV
2ztUZoPh80n7Ajlj1BPodCZuA1Elkxg6fqro86/g2JmWti+wuEbuF7zFOcjPs17g
m8t+6ub+Lj9K+MJOFiQNVixsPuGbKs0Dh+hSaDQPRdL9kGZccgrixiH2SUwCtD2C
BYb02s3AxbDIu4xFPLKGNmqk1vKQnLwhL85xI8m6aT6Y52eJx5tOw7dRg2ZnSps3
iRN2S03WcIKqwM9UjUh7DjGAhMUmAKPHApw7/hEldxNF/A53KJ/Piz9hNwJe635U
b4PAFAGJm0XlRc38V3k9V3uQACGih1fa8coNUe7wloKzY5nQbPoYU2UvqcakUgXG
bEX7khqKKNmgYfmnOnWpJ3pFM//8zd/Oak+37idRDOYCVen8jjsF6rHx8ALOUQjy
1JKe8KFz64TbOnAQd3Vk1SFIZGB8ofr/wx4YuEB/pUlFOSArsr3f8AtjRDthv2M8
4YZXbD/hRRS5eQ/iNTmb92XIEhmonNk39cp9N1QlKQAiCFKIVDlncuQ8TD2dmIVE
KJ1NxUK38+eZkZeseXX4A8yOrcJCi/xovQqkUa/Ej05Le7gwAMaQQ5F12ki3j2mf
N/idv1sMoB04qkcRbxbT54eMDzZGkmuq9wsJN3wfdXiScgMAedg6O/DOuYlCYZgF
cNRvHYAcyW2dU2h1Adg0/IN09shM9Ag0a3yCmI7gJx26BR4dFmfBb8vP1L9GSdOK
QDaSTibCgUmnxZBqi6j38xvbJJn6kW5ohWIe9TQuR0sbe1ttnQXtN17lRzdLXIqH
p83qq7Giz0z23jeYuqUmZJPuNgiXXgD1l7dDUwBF2puS5RL6EnasL/ltAwP8yZRY
EHi3XCIwNfeKsZkMbwYmcG21+DHaxc61xye5x/EbyAjPiBIy9Dql45kiXvw4z3PL
e8GTjnN3gNbn6/Qo7Gb8Qi3kx8ZLDLOTF0xec9PsPNvrL305BVLhIlh/6WTweGZW
FD+zYlgGmv3Eql67PxY6cJrZhdpvhkdcO43DsV0autA4hegJfcFi3j4nUMOwofIR
tetWn3o88GkYouBk6twqsSI2gqblD2xeoejV98myQU+NdroJHygxsne1K5/L4DhI
vdnKZXp0l4c35Xq37PwfZ2eb++Sv15PmHk9n0qCWkkYmyAeDWZ/jro3BlHKv3WiL
CCHGfmH4y9R/tjnSZXAMIUxSkybeDS44KuPWELgBlWGPlEOqfgEL647VvdsOdkqQ
Qp+++rcPN54wRVpJCo99wliS7+dWnkZ9c/AaIF5IszgpMJtMtqJBMh1SbCdm4T3H
EGHzFv85DAMpHGYt23bWL0skhrxwA3dWfKgl6K0dLMDSPCLmuVwMsZmcL5UbbPEG
yDtrOxVc0oCGtYsIQNvYdWUtLG8LSa4C0UfeFEOyQ9Le/xWk2FIDhZTFPWLLhsRQ
VMS/SYiJ0mPkP1eh2XRO86PfzvgxXgjqTylAchNCpLBAa4VRn8LIDUN5I7GR9Qem
ZMFN6TEXZi3fu8HEWgRUjTcxENMYX1f8xA12PkzwvC9hCLJrZ2Z7d4iUxPd8ieLu
5u+M5ZKEzKFa8W96MMXs8duh+/0tT3dMMIQiov0eRvJIl4cMzL22G4pczDfasE+v
vBfUcITSlQjRkm9qpvK7H/tB/vfW3SO+CVAIzrXmsiZ+Mhid0V+itoXDDBC+yzZI
waXPvK7NmKnYobGOmw0sl/YeuxJ0SFF6pafxGGzrnImoVIpznk4ASUu5Lf30oOlA
GU10kX4WwZ5qO8+z4J+FN0HGyUQtiv0CaU3cF39BAhI3BElRyyzXgwKBqgWVYBtR
F9vjk7FjH9IYt6dhVocaDrPkrbooR9fXFbMNhAHH03g0PJuEvC150P3WBrODs4lA
g4QQvtHhHg2h3hkyVx1Ft7jO3b41hhiDsWnLtR4EYl5i6dB6Fbv9WpEVmeTYxmgf
ajc+EwTKlR7aZ0WLbv3Rpxhwhi1zy6CCwIK/AzmqqlkqB1v9bywhcxFn9UstQWLv
hgLZ7J1k7wXssNFMyUu1vQnLo48L6fSyzBGWI1kIIZtoDIf1GOTQnM3iEgTZPkdF
rniyQ1f72R3updFo2v6EH0zSkBdUMZBLFCIp2qScGtGzVh0PxU0IiwFyJjFvc7Zq
E38JFf2x1qoXaH0T70iuM+Fbn71aqWkTV+BWXuZRD5NwBpyhbwMijveC6BNSJ0M6
LSxCmwO2TTvS12gTZZzWlEw7MTogx+TPapm1p3TAUV/xXP5n32bGClQFzNS6qNOd
CISKAAAPizClvu8mms2WrZreGI0gnMVdtzVGfpb4YWt6WaDisRfmOgiUojvGxZKa
dnYeECtcv3eKjlgo8bns2Uqtke7sumDfpLV141olfS+7o4CsdC/xXvGcpBazySKd
SsLDv3E8UBT4e8XCko/CB/BIns3QFK3GxC8QfzJyCwhMHWqLFow5AdDpqncSp3RP
8++PkM1CcHQ4R8oPrl2z66uLbFdofRiwoQWq0JTfEU5szR6dx/cUVrnxBerSSMg0
60rgRpAaCrurboVhLhnskAI4xhQ93jNbygW0Ot7BHE0PwxjUo+iJsq/olzRiatNJ
fHCZ9FOVehIjBFgVaTd9bMsUYtMa/xbh9GFMAzV2K7HMDgbrNlceQDTp9VOGGUgf
TTZ/1O2WbyiZD1xa5DaW9PgY37qJCo4U6kicTS/PMok5Uayfq86CkeSm6O1/V2bk
64Wuso3YVJmKpNQ7lu3zi1BaOTeH9xkBdjkZgRwWMb5ek1R/mb8XxPu3zBY1tuHB
2MlD/uQv51nZTHm3mc9JxW+EVgqn6u5KAQhjdafWmBUQyf5BK2dxVLt3l6VtRyEN
Y5lFLlKe+TmpG1MKMOT5fJvO1pn5V+QDMREGnS0vYaZIIKpaSv7EPtryPfIhi+sy
llGQidKupYvITLMCCg6FVrcfZX+NGayo1bZ9HyAwq9m60przxPHh4me7tVJQGlyo
mmnhOtkmGc+yseMt49W8P1VmGEVYgHzhJlMgIeVZfQDJ4SrAFBHw+8R2UADwCitt
qq+AkcEnKzdGy8fwDpQgULSvLXeLUEyhkETPkHjjwuSinHDWd0xItDbfmWQScAsf
OtFsT2L/Xbp1Xvg5AtTkp1SB8hdKfeOQILaek1YZJwLbHfXV8/qRk8/oi6gNUKuJ
SvQ20sD3+TPI7TzXoGGBIIaGciq9HeuahwULABd8dsc+1PyMTXwGbkZ24wpQy5/l
pNOWv69YijS8rmX4zLQQb3FhZNQQW38HmmFuRzp+HzFYdBS0DtYa1MbHzzFoYA+q
jUpLmCe4L+Aw8UU9GMQXlFUSOWqESUi5JYj6Md+iJrLjOdmz5Lz0oGA86+hpbcm/
0SVYm9LqGsbIo7wFsMOfS1Evu3qNger16KbPiScyoQC5qW4+gxjgms3guYqVj4z8
xNAmrEECNis+2KwA3tqf2P8nlQ220OWfxfsZMk9UA4PCOnQJW+V83uQmvtb3yIJm
WCRi9zpUhk9+JV8croX04Ab6ZcIhq4+gYiKO1qHxauLyGhy3rVjAB0Zs1qIasktO
MEPWmaAWumIe4Iw1B340P/bK2F0inQXEC4ASb1ZvPT5jqwzLMybJLKhEMvsmb/9Q
sN9M/ThHwYL+evBtmTPyVAl9xRV73SyG/aHVgP8yOt9Em46AZYo/3VQrJfPIYUOb
k/E2rbrxEn4sex74tgCP13FU8H154kwj1Sgcf0tuwtvJnSLqElaPIRmIWfqbTmN/
0QFr2jAzMlYQmwBk72IPjS8dMAVk/oOguE/xhGTDl8UPu+ng0n+YH8z8meSMJ8x/
2oVdsfC4jDPHvwqLXQOvnQ2XPzJUgvIltv73gZ4q78W2pZrvELOs8mtKhIG06/ju
8XkESZfLRPTnlUH3pGPcOL5LfSWhQj5pNFxL6/k2zigu1VyHj7UJe1pzFHgk17AN
2aFXgSfcnttuE2TmnjC1wnSOegAVVCcXdAYW46P/EPlPcc632mMVrAnZm0tUAQLU
CCtpV1SQr+meHGxA92YY0pIc8HgPhne+6VpJCf8YzyLSEz4SPkd9xFVhcOflaIc0
MTf6pGYY3utFbKUTED4UdrWd51l+etWj5yc72xdClEUMCpmOZWKNqnqmSOfYhZ3n
bnmwtVgLD6H1PqkfYo9lxjxZ9Af28BrD99TLYD+fVK8RW5sWu+Ad2fw9IkkYTbxj
5PriY5Pj5hxcqilOBzy4fcdMpEwqh0dsl+B3faulqTkHwlSrtFuwMV3oQWkhheMT
E1AsM4y+C8v9jVEUm27WANw4yZ8w7spCspCwUmFraYc9J2PIyklhHL5arjfyphZo
tx5zhQ7oawWmGbJxf6qJSw0/bxHyJX5WlM9pEd7SGfm5ik1wVW6rwFE6+2atZXJl
1voUXoVVRLyqa61ToS4rLWra/4Q0hSqvsK8RjL1En3BqW0AJpeNmOQf0crqrwvMA
/z+NSjBGX7lsyI2HaXZTJZ1Aae+dDj3tNs8p6DQRBxFtWPZ9121Qe+Bn1jxdjKfX
0l0G0fkgAdsdcyYVKNrDh2CADQOYuwA3y972cC+zKe0N1Bi9tgUoNPD+RfE0ps4k
z+ylNX0I2W4H8AqY4lQHVr9Szt0Zyj3hCE2rp8aBtHyEjJKgwzygU08a3C/aYig9
xSchPqv1dzpSF8wdARDIcOTR6AzmXhuN+S1/IgbxsYl9+OFdZh75Mqu9MERmc5V7
8glMnLI5br9ZOLKP3roEllZwU8jr4KR0G3MomyBKgR6MpzEZZgSQlbm8dg7XiNG7
3WDdtHxpwsFUWLIehSgnc2mYZlBgDue4kjN32DBo0TgnJ6Y4a+N6DrDrlJK1RoKK
tZtshWzAhiGqMA2icvdttyQ+mv69U0zbKP+8jiaDhgcNYGFBirQfCNNGJ2b9t+fc
2wphNVR7Y0WkwoSqjjO+0SCEeyTCHZLA9S8GmH9prn5X8+LBRYBxLPXz+f82XEH/
kVF0DwpbdH1usxlSXR2hbRk89vQEYKzlj5UUpACfyL6kn7hw1jFcP+zFDIChNw1x
Ud5EdMeeIgC+QnK50vNZwg91AFXZ4Mg2/A8Qz2l6PylR0ZnVhdaBlBAjTJ491qq3
NouzVh4TsdmwVU01GhrobRUAYQ0WMYCcj+48iic0/7RgSm3pMfyaUIpNpcVZvVyA
/3fvqBK0rlcNREr4meTchLQ/I3BieHTVmNR9CE9xqzuG0Kxf7b54s/Fo8cCVQ4pH
xDJPGjZnJ10cosLki9aYLOEGnJ00Shc7WTILSXjOWo3abtuBJhzsWYEsbXAhlR16
lYGAg3FkuPIl6j1m2CaPv6tDu62xJ68YNYqAoryByQuezwj88guWYwp44zwS9DU6
4LlwcH2+LcFzd4eHY71xbgyvgIRP/4pRnTeJBMeM06RKUea9XC9JxSm2mwRqwhmt
Qwd4DCAss+6wG/IRlG0dCMWh9DFmZoMVXNhHR+8wBhORAFLQtf13tgevuW4yn/yv
tV5Dh/uOGEAGg55WSlhbwBrxo+Qh8bhRSMiXozxQ6St7CxPAXlT/O1EgHhYYVWFC
zZDO4X+WLLfC4NZd918IUJ5wTGcSDM+P3/wrKfgDLO7t4nvArBiH3vNHZW49Y3n6
FRF2ffbj8lilZLHT53ymuaXLhXMsm6Vbz99jmnlZ07gxa5XLw5aLFAAKW6B+xc1v
pn7Ct/CYJUDb0BvWNGgQoYunVRzkeXrnaywqRAfPf5PFxVwNJjeUEcaB+b/anE1q
gghVUo73nfUgnaA5eRYTYrbiC0bKIfBwuVF2L+7O866mv8Mz8OtAE6YoT1/D5Ael
rl3tZedJudEEAL+YN21TTazA81DyhXpu8LEEV5uv433E0/Cd4K2wzyVV60+jdCk6
AVS5G1QEnLdmxA00gOrRnoMYX5ESn2Jp66QHkHSMrB40ZWt1T0i62q/lCgL5IV9N
m7EFyvfmgYwAo6CwnHANPoL92Zvr3ZOQ0z/M1sMwR4pB0t4sghAl/FUDBq1f8Kf5
rFMYNw3nG6G5XTHQ97SpnBzhaxvavY1ZS9Tzt2XMLpVDhKQul343M2PI7wJjeVeL
Cw0GqU9CNp9g4QMJEny7cSNP5op+wOQlxOnKqro5WPUUUr0TYE3LjmOOEnpiaG78
i6zkP+fyCDL3CB127w/eb8JsLBfTsmujiPvakzipkO9iHYJvzhvIUQezGbS+lklr
gU65MdPKOklfipsfZQxcCRnahgxyQF6f9IkZHF3lHuqs68AlUMn4fL5ckVA22Liz
KsueKzSpRxWmeZ9Rw2UD2dUhDzB7BTsRTcujbqJSS1WWjvTshNokoLSzQv1USYYh
4gMPFol4P/z6MVsAkE3toE+jrxL8BQGoc7KwiP/wxIN8oXf6MkKQVgvFpD7jqgxt
UJMQoOmEvDOfWxkjFxMJoiOvtMh5KhEw006WvYYf1M1gOTk+MDMFJCLIEoNdd6cB
0+YeWONCioTvMZJ9Zv9RTQOChdKVf5i5mSoE+Dw2RE4jykRnI9r2RqlGkTOU1a5s
85yKLrPTmbcuhbIMuAdZ+Ei1XuRZzZliuM6LEX3+SH48I3TGXmifwxtDEx8KOGDH
o/nwphTaNuoPOQnlERu99d7k2Zl7BEkMJl9/6mwwXaOTvRwpW4t40Dnn47ibpkUn
eDul7GLp70eL079B6zv1rsdH1eEM2S8zYlpbeLMsoLK6o0YoUCOIFXT/ZcyF8Nu3
SKR0KJZBtkeg+BhPakJL97m3DGYnuqIju0DyBGR70la9iZZFy+fVZu9ZLflJB9zj
A6PRxAeE7LVlVVyALV2GyS4cL/1xz9LHiMTTkbuwKF6Xl9W4DXBAk5CS6o0mKRis
hhWnIVEN3y59x21i/Pe1oOWtR4Bd94NvobjDxH3TJd3LbB+pebI1nP07Egvz0nqq
36uZrEi0uKuV4zMS1u3504bwwjNSSUxD/fiDRSrdTyLWzyweErynStY/76nPaGp8
Ec6DjXyWw6HWoQJx22HeqL7ai0Mek/iEWoG4m0agcZza4+jGl3BQOLZPGrlTHlJd
5cerWkH+stflI2bqwTggz2GrsP1hd/a1e+3QBgf5Nso2Q17KzhZn7i14kuT6lwtP
dAto1cy/AfY3dzhP7NbWlpnE497n2xOC+EoshPRhZXzoHapwdJydzb+JRJnn8AzE
NqRMx04hg5jK/hOmXpBIqLYxy0+WJoOb3G8R2fqHJR1EnuFMOw9aWgyD69gVyUEq
VVX/yy+axsFrMASwcdlwqE2mUFI+2NdpX/yb9xwVJ6jp5wjmTzFtlxCC6pMWBXFe
QNAy/4DXnt6wilN98JVxAq6rajtGyinqLz51URbVoB67tMuxyph4YxdA/hWRGWCk
t/FPIje4wCXLJ0X3FrCe1NXD3WJW+0cw4zbkjG7MajGmpbSn/+Ltmf8NewYg1OuW
1KSft+X5wtk1e7lxEI+InTT69JUixB8FSlGTHv+KlYW8hWBQP/omcZgGsTVD9iGd
U87GwD6ERTphz2iwptR4OmYnoedICUv4T6BdaG2zwUr4AMJ+5iwC97+YK8AU/9ym
CxMpaUdhiCU/J0RSGxkgSUPveIIF8FdbwctvuB/ZUs/2ODjd4VY3reQ96Jtvit4+
drBolvTCKffifxMLvtH7CkrZ89QI69EbU2/yxVEAk+gOj0WFTuy8GlBlJNpYz5KC
HTyHJ3tNcKDv18XoKOdl1GBHMvV1/4beJVC5Yu+khultSZukFNcJFIrDkSFjrQ9Q
9JzLYHEz0We+L10vj1EuSOAYtIH2pZfsTfXsCJJPfFAWKGVi5wG0MByczGbu1xXs
tAxBvTRcitUuVAWlkhbycmDrnAhzyccimQ3aDbALz/PNkPRyb7CO1HMzFxsynv18
6SaVof3SbVXzKrcdM2sRlijshxpYBE4egLYrocgCDwg1MI2OtCwA9iXgNrncFF96
KPtXQhrSpTbM/SxTW/nKxmAadXJiH6Gsb5A2kjhgEG+FbWCRTiMWWq9ZIGDsH1fN
z6KUp896YRS4AVa2qPOcbBcWMDiXG/w84ym5iSU7/HPER9n5oOnbBmV9BUrvR8rV
3EFqyKI0NJUEXRRZ0JLUNGQkiB7PhilYxxVWmiw1DqGqV+hxox/MJoAl5b6nKLmw
qbT/b4SbNhK9WV1tlj2uHZsF57AmvxL6AdOJqzDT4lQc1GqnnlyrwDuLSyAi4D0V
a6vaVBsadLtiHkLAEBC4pyANAN1YKrlSenmCKDnGMgqnYi6TnHePAlxH+rlMNAX9
33hL4wrEyL6ndmKgnH5mlD3Yc74A5DEWaI9mtvb4UqDobaaqZPpuR36FphFTgouV
Zst7cGVTI5i4fSZlRAn+DG0v1Z/jiyjlWFH6FBF12FKGBLjboOlqGXPCh+dLlLc0
i7PHv/3mC14axVMtpHiS7vaBkFphzOEh+9Bz6qRA+GOj4pW3B4ksBXMpZWamqRMS
kO5tMiTq+cCWfckbK33RlcoNtMuxRlcQk2RpmzxMBNAh2eSHS0bqHtqKorirVTK1
EtFsqHhDGuyKPadi2Id54znFdWlqNcqQimesNDSEedvJXvW/5wXMil8FcE8TC3hg
+FD1H+d/Htqlk33xzZEWMxsZuUdjtor63uzeASLyBtUyCeTAAdj3cP1eZJ8HfxuF
/YECyOEo/MoH/scbj82E9+aVZPApvRAjzg0ZiCzq0atH0RLB9cAejQxd+nd9WxN8
NKEs28EAj1xRqodLwtkT72BNNGUHdP074i0Bjr2SCoD8d4LzcivQED2RcOcY7U8o
Pg9YaoHs9DytTIlo1PK2na5+UIYoKlWTU8mjQ/NHxL2krNwA9k+WkD4RYpXzm9AC
2EAqBPfObdOtupZrMu3z43JLzZjJ6oSvD1Aq4wDWMOA38i/bbx0VabeDfzom7iW4
8MDIuKrL/WbQY+R1qj++P2ct8JmT28zoBSlY92jj4oIP4WW8bh1yBUaFUhzOfiaR
/xqfZboGSo6bKe+SbjJ+e+LW6zx5//akak/mmZOGOCnA+tTK40xo8bLmuqM16Ri3
ZG7/YD8GepCecQwRE4aPprNXK/kzfksz3YqroyWu/UVHRpBqA0uftQDrJhhMt3VB
JPrx3c+IoJT/PO9FX/YWD65MQYdLdsGkwrmA2lj7x/DOI2ZkRa6JQfFRgdxG0g1m
gzyLT+jFUVatdMlu4UWrkeTi5uzo6xlXRG2TtBPlINToEnnLFWJ7QJCdCYXSx5do
AJvQuCpKuCC8n+xR1cGa4pB0vBvZ0wlhJH76/Mcivdh66RUnfxD8XD8kghYCb5Ms
pB9NPSIXUpg4CnA45ikGc1Lry3WhuKVTPEAWrRLBTCqdVgsPlDnOBxWirXY12yxE
o/I6QRWz7O0QpR1XVWqQb+CJcCtOMWPqAp1IBaTliYfpg2fEIu2Isau34W9dnVlF
1ajgcVa2D7WdPpyl4Wjf/TvVovcY75eNEoim8RHOork5GgcycxyEfTuvWQ28T+U9
X6Z4r0F+Fo5d/BEO2chFSQZWDsmRjox4/warOUXaXAvtXeFoFcU+/27GZ1D2h94P
lWXAdoMI1SW/8GUIbfcuqCOFkm5ex+4eKt33h9Rdd2q0hzGMHNnsECXGdFHIGaD5
wV/9NcPsxQjrWD929jHaYbQgFujZado8O1g00emQNp+/OmOa9ntUO5iOoQhrrv2z
mBtH3Q+bNiCwuj57aC/cW9YwMXOjd7o4bOxAHxWdHUl4tZccBEBUQQXnP8jHUcDB
SaNRcwPMEVUdGA20MmRd7ou18z7SUes8hR7+dTzXa+59dPH5Cd02GPnroTrYuawK
aE1DeN/kBj1HFf9aqyDYdvzAfUSKN6hDRBIP1VI6MysRuXK4+EeUkd08qievvIHL
LIXNOyZCJAVOPTcQBGmJIwXAsIXBbEtf+BCWomxvWK9b8OJ5QOG1r3PEZi60zsr5
QJyD1i3DXWpxyx2rh+heGsVYonr7iIgHGWtknVvZC6EUzRRD6EgW3pq9GnZdhuoR
CwEv8icRy71pICTrIqQAC7iA3mUl2OnPZlnToowS8WEc12UyACdECeNg8mPXneNg
wl/TSWHs4n2j2SnwlQkAGlvOu+P+H9H/01dX1FS00fSQF0O2WxwxAkllZM1nPcpA
XFTXFcQq2gvhABFRMkZGDsGtQLgOBHBB0cP4s4GXD45rWuvmduV4vSjUz20tKyfD
COdb2OBGv+7gqxRVv2Uohz6MbbTyzkYHM2SO0HxWKdvrQutQc6PeBfv2t+RtJZ45
clUxs1Hl7VXDlDTsrKbSNbXUCqYq8ZhqKM5+/A32Ucq21ClH8MtIaUGwac3+oPvv
ZtJCuUuJ64+LJeEdt+6j4XrwaPjUVQ5i28C6WsmntENdM3c1WdilMul64gzENvc6
pktKsvj2B8ne36rTcOTIT3gOb8HaMTcWI6HNIBcxnzLEPRdW41dKun3nVSzDdnZZ
vgHr7RE/aYPeDzPo7KoWHIUcUkX6D/41wMRtWOAjhEAcci6fOk64sl7UqaXgclE8
9r0myo7zYLVFXBuqRwSTm0kFSx2TYHIkAbu+CyViCJvkqynPUk2DklUnKl3+yiNX
786fC5H/B/HaA2uIdIo0fNq0TuNXumZm1LNC6dkXO3x/Epc80QZcEZ8xSThuPHDG
UASOTsyYfamh1yDzknmjjvHia3hZMtIE84s64MNCxsHSsGn4btAFa6543TdHdSEJ
atp06FNBZyIL2eNRz8U4uSVRKSmH4L1BrNmHphDqpnUzuND9aj9DwpBRhM58MIr6
WcMNoASlzib1J5U6vFNHVhIyrluvq0Stu2M0H9emt1jJIH1Cbe7zWj1IoxRm7CZS
+4JKpISmbs/Dd03u5Vqc+Oan9iRQ/AU/ZmKTvG4F9tq/L/NUL4Blh9h1joMppMM9
kyEDu9SwMaxj9m9T+aa1MmGTS0Y1IPV5U7N8NXk0TgCNNzFsTH29T3enlvciht60
SK6NiSJf57B9K6iXC9eqpNz01uIEVHQ1KLdVxZPWeVrRgytXvUqvOd9I4HLL6qcr
6qoTha1nJU5W77UpXsR3mqfTBMRFZtXBt3Okx8pJvHCdwMr0oWgzoEGBFKk21+XI
9HUUAyTsTwR7o2l/E9NcH5hZpxwFE6UbuVPcHZg6W50ACN9Oj2N5cwD8B/MESnry
8KaL5Z44oYy3JTBUorXlvvaVAwG3YN/U6QgtsL6GPj7aqCGCgHHWEfkjnK1xNQri
OyMygrvD4PkK/LUsH/AqCoDcEwYOkJorC7XiehCW/MqDsCZEgaEoqmX99/47vXwA
i4ocq6ZspO0lQ6W34juSoIYc4j5Gss+iOzc8QTgkfaPrStnOJeedgsNeLGchKV+i
XqaZiHY9KzebGsT/xHkGMVNKWAKrpOwXteDnrvDgYCC9aRl0McZ3/judr2xTwdwH
seswCUc73wcWhUQlLemdNQxN7d7pxj87oqnzZoTET/uuvxKjuo/nJP8WXcPJUiu6
KpSTx5jRtLMPqm6Dkj0b5DD4dWFlK89DoC/iN2B57eHPGCZqWU8d7+3FzY8528JC
QMCuO6N2RYIdTBdOkfLD6cBiPoq2QGfCdKzI/pARoaSz2Q0x7Lc8wdtGE5kPgeVT
Ep4OddbzBAfuFspapsvK8yGFuQ/3gkw6IaHzVhn0tUz7U/KtFX3YtBmsPcQXBfFE
5ljQDi20kKaJ3eAjKZR9KtAVL9gA3Ba0VQYL/7Ihq3dG3CAyho4xhyvkRD+wtKzE
XycInVLa7Td0i3708u9XIjwP3DgyXmwfxYHy5HpEg+ESBF4WJE2nCbsXjTwyo/30
29tf8tjcz1I/GyI+xmG/u+He0dhJ8dg9u/8oqOu07JGpNeQ0hbQVMuGdGYc3/TjF
vaD0tK5FT5Cxwri932+USpu41miz1zQIp0n+DCbJv1NmPtw1psk/dM4VGfV0WPF/
56TNFjR6xf6XOue/YTiaWuaiqXRVzqBGYoSx01y1smXxWlYLMoRMEhY9Xj5mB4x8
vmH/kGSOYS6dmgVvOBH9J7qLYF10mvDKL7UQW70laKYOGjSqM+w0wyYP6CwgyPKI
Z7SkuTgPcxND6plPCZ5t9frluIx8lp9JiXxOQjaz0W9XFFoHWBVplkW/XjKgMvXK
yGYwUsEaHqyV2W3LbKcZkakjwnICP2wCwyiuYZtR4mz1JdancSrL6Oo4ivnvB3u2
Ph0AFsWlh97IUtfPuZr0B950aImI8yrR9awdWej0OEjvq4dPDTSs00szOrKB2j2N
2EJcGF425O/LfwK8W4SS8G4I/YoCgFr6yDH6aZIwBRNpdy0M0nQ9/GdNgBC4c7kc
Dg5QfBApci+IgVx+UGOcw85h23TBzgWxx6G0hITO9GS+KRylT+LwsDenbbxym20U
8W02Qqnvu3evGp8UcsynKnynk/7wtathXZWRkL4YU6rgQ/8GfdgXiE/PjMGv7FPh
hZFoakFXLcCxXkXidXxbxDKtcgcTzLO8ThDmIQT5kQhVfeGR8nPXTrGOJqD54arp
GKtwQwbORtkZ5O3tVGTNksWFrxKh2Gyf7qcxzuHJvv2EJM1bGjvdR5NrRklMDshL
xOF/hXHgU/2JfcBU1MkBIg+l1Zr5WcB8sqHRpQWKrQDnsC6a5ymcJosFvNRJTj4X
of0sIWx1SK6zOeexzKNmyDW4mA9a5mLZ1i98x7y5oTsTmpYuE7Y0Ftr/7yvxarod
ebFTKV9TGkMEg8hqfVGRmo832eRZZqx0PSsQ7JE8q64neIQP1qGXL2wqM8lfTkJK
2NcwljaYO2OXKGAn/E6Obiv8oBC4rPWwdYoa8fFWRj2+GmXGa4NnBUk5EWRPMB82
yv0vzi/sAnwv3B0AuLmFe2cnxpkS5dTbgir536Dlt2JAduLOxYSAzGz227PVqxUQ
x/llWwr5px+oGwp5bpsoDPR33km2YvaAiAvaKV+Vp8m7nSziV5Uf6ebinKAtNPRd
iJ3zKYeeZtQHD2zp759BXyCEfTWJ0lU0I21f6Li1ZY6jYzugiV35rSJZtd3dPkqy
jkrlrMe62N584uNjHf91bpxHCaW/ZcfIV8YaZSZrgzjeWIL/TfI1e3twCtpEyOJz
fhql6h9q27vfzatfjCpJ2KmI/H/mhxZ1fFkhTfeSIETTZm0x6YJk7kG/6KXQNpV2
o+LUCiD5LBReDnpnGlxECssh8Z/Kc54JLrhK+3hc3tpUYQMJXydsKnGGMmtViDBk
2Tn9iXoj5lutdwedUM0LG3Z+J9WxpTUs7C/dgV+miYG0L8PDJxLpyE/9PPliWMgU
iUZBOrCQmKMGxis+HSr31jIamz4hYmEyGKiEfI62g4kpx77CPhpKa+WFRP1gtdFK
zbMkfNxf/TmeBYYpJ1U+Tvh7hLs2w1GPrOq2gtppnShDpPRfM1YX6scKFxP0pXEe
CYKu8dRXWRdl7RHbkuYPZ0z6EBsNr+zSpz1oOyZVnnGQ1mlgXU32TFqUqcaD7ClE
ptJLitm5Q4eRB6EKHscJuQMuav2RHFVP+SFwTbQSbPgO8FAdFdnY0G/fDqfutJfm
BmOSwBrtyL2nnlQXeaxfowjVwCJUjAfgTnlNwIEPqztYkJ7dQj84YBHweaMZMKl3
mvYLBLU/2oU8fJNya7r4pXjtuXaiUL3iM8JYFxtdSNNDHdRb0kKMzuKnH5D5U2NY
BAgClcsuAGI/eK0tbnMuFxXYMQCRBUIVnzHGJZg4RRLZ47fvcd8bx/QWujQ/sXyL
rojcTv2gpyS3fWayGyybuI2Q5rzY4RCSBOXu/bj3//WJ6V0jyDmlqZr/ylcglwjZ
WTzGrmIfuNpcF65UqdJC5MuRFMqDHnEBHUVbYtuuOOWkdRL6iPKMBDbHiuwY7Hrh
oB9SNrbuy4AZSG8XpvQZqVP6qFp5IQGOg1HKaQu2R9R2CFNUS22TnQXpM8/IsUxr
XaC+xMdd5Ce/daJ6wLxKDmih0ri2mYo/GxZLDxv6ObC7Ov27IC2DrsQBy6JXeOQa
12n8WOmW6DVvF19wo7o9k8Oa0kfeyKT1ZmdfJEAPmR41lKorJkh2JJYtYRaT7XPR
Hi04Fi5On8h/tZjlBbMRFVHX3Q+Tg/uUdCpi608ut+z/SuDxDcFQF9SwZopzUxad
XilmejhCNHeSR50J9KeeYPfMjaQHXmR96Unw9Yi9uRA9EPGHhutRs3+cbRNgtI2U
0cG5bJsNYXa5yO4YsstFOXaCeMVlI4k7vR+1DVCXYDhKvlZjh/MF2ab7/w0LjAXO
61reDLo58SoAWlnI6lfG71B4fMu6ZcJrsehwtCL9m8HiQEW/77Whr+pYjX7HnqMA
1lvY+9RpEhxBhpn39THGTfooISjILI1eKEUNEtoh/N696fU1PKvvIv5yRs2G3B9K
yfK5zAA69RuV7fSaaBZD1128QK+lYiYXWAPQ54HZjgWUU6yJXhp/++K8RIxC1d9A
t+oMQS73I1BbBhuGabrKgQuCkiiD0Mbs1BUAVn+li+PtaisEIz3iRzl4qBLWUJYh
H14wquLK3s2mB3AWaN8XN/coqwK4KcfmeyOF+bLTYQb/AYOgSTAkvPMzZ7o+G8r3
rheNyd3uHaJxYO/hFAuo9onUQLf6AQxafa/aBNALE9ttRgAKYmKECm2dNUEPI9C8
2LYaddjPRM60mKMd+OiyiiwdkbPW6Oi3b0hhar5JV/7yR5QlLuTD/mnQC7U4C0sD
NJUlWb8uiuN9XugjnJq+6bMHpf0wtevXRuNtFn0dhmPQOBjM/BPDDLvG8nfob+OK
1KEvSnC82ZDEtM6H3JomZHeH0kgGWEPBel9kMwupmQAf2/1vgTn9jAUKD5+d7ZX9
jfjpLBc3odM6/OPIjNsY6ku2HI7cUMsQh7SAosd0+R9ls9HGX6r3QK0rlQJJsF+I
hjMrk4htIfqbkg6yGJw7RnqxHF1/UaWFUNeJcZHGGnd2DdgJSzGZoVCEccU2TFUB
P5+y1FyuiaPvhcnNKWJC2SPoV7A82m1FB7Aq6DqHSeyVRSCOPMEGtM51R3Cl4uOB
49u6zxVSgiZk59J7cOCP+QU9J3YpshcmHC5ejHLJpVBOBQEaNRuwU5dmwTcQpX8X
J3/siuGmmkX3DqEKFBmt9b7F29Nud9oFckLMwiATCOTHaAM52ma/vqrSnD4IhdYn
Vwh85UABGs8Kb1npwKh1UNPyLTcsDHnJyKFxxoHfHvfqi1L/L46oa4eP3/d0/Hz1
1ZHfKfvn+Kdbtlw2Mt8/gUrWF2KsMRllf6ytq2WbAe0VuCZtab+HWVizmvQ/kYli
j3TqaKcQrnFUI5g9KKIOl5ATBo0xpi8yYZRnlai+/njr8MLhOuL/RB4B/7umfiOY
hKblgkvxbRMuZCWhhQLg8LToJPZZo8fUwArZuyZ764MFWVNh0Cw1OExL0GIbjlP8
avqkNkb3t7shk1YMEegkVf1xCn414uojDLkhdFKX0KvVBaoj3VOF3Csbtr35fi88
OiQE68bK6o6eB16+KBNgot8lU+F+9Gie7RtyDURRQIRoAUBGh/nzXG23zObWcqeT
7fbGNmLFdnD15JUh7FC3TcH5Nyv12xkaIHO3rzRaxZhITM4VoxbXWFNXsM2Hg7O5
NAMG2qBmPo7A9PdFMrki92OlzYDqvN80mk5ZYTi40UnDA4wUtrgCz+1xSPX7j1Zg
yaHTRlMcv2iW5VnKerpXBCJkZCGOPWZhkSzEbTDUnzoafKZK0k7L0UVBlaBgezo+
9vhzJ/pdkZGj1uaD5Ezp/bGFgBJi0kopOVWonJyFpZvQEDmfQMdh5CH2vUUXcJgB
ZQ1UE+8BWBtPkEO8VbHpJeESCTPw90dz1mP6fDCprJcW6HPepMCN71oBJmKcYuqZ
OODPjAB8Yb3vMJluVSvulkXhLd0MaZGXfPorpFIHs5xLYJEciFnndBuotCKCgsHD
8DAY+YFSpSS12j2VhY41WuhcRxHsvUQT/K85nDpmUnHxqDm1ISxYlLeSXwh1EIMy
Q/+KpPjQ7SFdVLN/u9fmBTU0JzTMvRro0wok7iLNyNzcoNt/rGn+labx8KC+VLuI
LXN4FFB7KcqRmIirvE5F3pJ7DWcMpi4QDq3JJvylOiteTfhy9Cx4N/mkDfB3IiFV
RsKi9BMbmAxjBqtvBJbXslERgJ0tmtGxFk5h6Lyh7U1/zF93tEVQ0KAlCKK2PdVG
/Ef1MQmPJnNw76FvHiMp8NHuuxcRRkWEDOlCl1HgjBWv0ApkODitu082TgfkM2Ey
7ugxEiwv5HtTbhCsQWh9wcR8gfdnsDuMb/FDKQ22fszEKqxNAEOjEhwoTWGLzTz6
xuLql6ebmINJOjKsS1OUX/pT+UQrrzINlWjnJQmNrfC4qic3u3WC0jAY2uM47KP0
4oxX/uFN9q/+N6rowedl76jvQ0RIPImdrI8hHGd90dKFHOUe07dC4yxxC/dR4A27
layOcvVBIeF2QNGnJeOr2+PqOETVRPOYVjUvNH6cy6Oor676nbhQ2wbdcLiBR6qL
h6/0mt0iF/LGamaIkrPr4eDy6BuC4Jjo9BqnaXfwmtQn2h54HHo/Ir2Mf7HgC6Pe
s1VgW8BkCsgwVY9RstAh2ToSB5HJo5XVcss86hT6VUdhHL5HAXYYZq91x2SJ3ejI
+1flYfoL9P6RIMbs63K0+5qbtc7NgWnAbFtM31BJiuKYCmFgWlPO1+4+UYTPAdsD
YNi9VyCONMerQqRariTzzRfyMkIk1nzRJDZTXhOUsen+OMcho1kt42seOb7+ZdLf
hRpVZTGyXjf+8xjYugAlC3kpwiZAonsjmQ2Mqr0yFCu1/bHwwlwOV3S9sEVYvFIT
uUvu+dApC02IC8VJGr72N8wrmmk65/RcTJ74CshqtbCmTl4gw9Si74X98WU4VZNt
5zEw9Pay7TkO1jrC7nE+r3y/q79icyDayRsqJXv1HfS2X2snoXp1pBr9gRjxVfoQ
KuFl4po4cBbuaNl6oFDBd2TXQ2YKNyWv98W3i4f2pR+AmsOTZu8MLhdJNwq/u62h
lRQn4IVAV34QtToJkDcZte9yxBdSvM5YxchEAz8+e6WIGBZPiLxulMcqqCqyy6GX
+P2PrhdMsFXFU7gV8gJ8BW4jpA7qTTv/lLPzeyfIMTpa3hBXGWRDVYFl/78gxhwS
GlqZC+FTopS7jj15beJzSrPVKQqNzmq/o15hL3vEtPjTBo21ODxe/PYoGaiXhYkz
G8LP4KUh2poXLIk69j91cfV+KmRrQTJBLzhzQIwygIiHjyNG0Sh4IfyPvWfLKefn
kshWIspLIPyZCZgunUFXxTIprbxfLS4I3Pv9s3OMgJq2LPA8GvF4vF1R93XWdfKO
35aiixAEu3Fh8yMPVc6HlWVsiTYYqN+XsdxYiVS1AaaJVAFeh6iefAqng3CXW2vG
lXox4YCCnmkkImndNhssMo1+KMut9VOmB/RfCcZ7lU4+TnDrZOC/qq+nkSqVekJm
49xKa44FjOirqHcVdT+PGHr/YVI2Yo6F8WLntr/RG/RHEE7lPmyiqtfNw/tmb59Y
YBWc/tKZOYLcwtcipRDoiSuFP0L8Lgp6HPSZCJd8EIXKnebo5adRNaOfC+QCNHZV
OgFHyflfn6hVj1tTZe4Rd3VOcBr8sUc8EuJ2Gp/tQrr3D1319uI5wBXcVKP8jIRh
0+Spa6thnYfCsJpSzfjre0mXmYzPtLe2053tfdrL4deAcjqBx4B+izeijEkyHjgT
AcVhnkVR+PYDWuv5wtFkkJqtjvEySp8vGohZZJrPdZvtXxuu/JakiTDrjg5YW9DS
oFrXjBiI6qS7tPiZ5JaQvDe1lXpeFnCehKnw/P/TnEsvUReMkvvpRwkV9pJofE5Q
TZsWtAtYdA1/F8ZNlhc1mscuFrzf8wNL0a2QG2aerFcm7LErvmL7mY5/7otT4Dc9
atl1KxJQ99SeyTxVPajoA8mz0gdlqcXxCplAAQ/djJiGsb5OVIz6M5nUxKOeXbFY
/myO/dpsPcxRThr8EMSq6TbleZu//vBfIhGf8WbGo5WdMzJwCHmTHnGQ8m/sUgWs
P3+x3Jdy+K+yP8vXHgfijfG6xSbh5VP0qKgMpY1YAYdW5NLPP8BvKPvp8gWRuKrT
HofrgwL1F5fhdveonkDeWV2Wcskxi+1D3aa8cfNtb4A373/fs5vXrgbN7RPlzHIz
l1trpsEhuPSKMzg1JiQalruhGg8Q8UIx7pK4t1Nb6EfFP6RIJfn/tgtOCScZuaMl
m41DapRyN3B3PZX/sQ/vt8Y6jiwk7f62zPsYmy2NYzgQsNrT+g5dmIsuOqgVe2vm
AU4WjNDf/o/jYYTiE6yDQNMWM1Xwklc933o4LMXmQ5DLZfLHzVSOdUJ+MOo3FrCJ
GDspmWlG2klHwhDCqW4Hs9mrVvi0VaYbsdAm+ndK3b1V6psjEPbQS32vu9tJM4EA
WH5tuata7GyCP+cYX4mhxezApEBEdnO3OsGJ2c1fmtR3vEPNmS9HLlDQ5iVyLObf
1D0/7pQhOIiscbHZtbw0AEPik9I6obQ/hV5gPKI27eltXhUxNJfTkAs1TRJNwL/q
m9dPGGXTRHfqVIuUBwOu161IhzBQW7nCxLTZZgHRE3Wi5b2QiwgB9aP5o5cakEiS
CHIRZB3rAJFH8tEHB10M5B3wMSt0L11SR9Ca6Nr7J7aMEtuTZBUnQKRsDkbmHorp
4gE3iRXXRulejFdssjTRPrXZ1grrx6hhCmYBUnsv+nhmUOMr32k8L8dv+qO1fOmX
7ksYPU4rp/6rhp+4HZOeJBd/Pr71t83E8K3zStplupsWcQV9RT5TNrxPQn5Gnfb8
2Q/m7Fbkj3h7MZVcskECSZlf22+ofmE676VsTtuljg5jZiKugrcjz93OA6Ny9NDv
+b+3QzfTYGoa+6bHmtz4PCiC2Pi6fQM7wFgC3RWmRqyvXvxOoEjqmeKMxCLbdex0
xzHIBHZoDARk5BK6SfjNrJUqgbZMEgndl0J/srpaSfwyjLGaOvvqUj1fHKkvC76B
ldyzAG/O3JOK2FIK7CQzPLl/sWZwwKVvlqKL+ftxxBNVrAy5Uq9OjkWDC9ubIf2A
I2UKHPbkZQP5cs+DBL8Pom8Q6zHd8QYigLLY+oLbzXzFKind8v1aZnyS0Qk15qXt
hJy1bhjkbdg0YmggaXAlLevovzerkSRfwsFN/IaFHrysxGI9VfY1mJynnMXPX4R5
u7GPVYRpRHXN0ipAxaYTp6xPXAW3JmP4rLVHDBzw40DDd5mRS9bHpvUYemws+pqt
k/1zovKwOJHtV6GkCaRNJcmtonL0oZmcBs2D9YCoUEnAKBMgEH/RiZQJtWQfjCaM
0JsrlcKJgTfY8asSe3CnY4Ml1OrVh5FLQ4cDEi1MLBvzU4RCq2Bz7FOZneWuaKkf
2jDfJwkSvcOaftwJkGbFuvKsUGA08WEOOvznUiZ+gnkHqC1kz0zNvAYuIBjOLTE+
wDHcqOQUVMi2HH8pH6IVGG73fWGrcfpBGv4Rjb5WGKuz38gGA8rnNzILWiBNcXRL
DVd5vc0KgNsX9WWKPPvrPmE2x4dxmltN9hkaoNlzyJ8YhoqdqLqz7fpwyaBIv/gr
x7p2tkOuL5F+vULuB40boz4hHpvMjuzjyaAX6ptVNuQ0LyEBu/8ic9utCUHd0zK4
Kta1Po9tsV8QpHb5O68B99udcIpo2urjAulb63yOCVYyMMNRzGMdTJTOtFkoFxU0
4xBG/i0KmEnNISLzGwI1QM9py4rr3Fm/ylGJRGuSpVlfrzy1cw4HnqF+K8QcwhSa
KN10/M9PM25EZ7KsWvlmDzXGpPPrXajsw0uNXwUGRrz/+Mt+CjYcK/EEYodokfFc
2pKTJ1p2ewkPg12Y0BJuglQ26JxX4KjM4nxXhani0BE0q/xzfjNnOwSUvmDagkKX
rZUauDgj4xTmD06iQeIFjM370JLMGXRUJrqthHsCzVG0yJfBFePaQ/NdDEQUeZNA
+ItCyeWBBJyjXr0V9HhaJqFeclnv4zYajN6tJ0RzD41+Z4FBIT3obqRG94ViGe8z
RttMmaSiymYwdgdC3xDKubuHYhq6SoUUwUjkOMDyZMApVJxM8i+vMpKHbR6jP5YR
seZJp9jfUpihh+UzMY7LOMMkJNX1pmLPFd51n+QgdWrRTqyXvWOX9LSfeZIsnByA
cPi1y5QhF4gldGmzUMjQDcYn757sZmAfUUZ9h4BCJcx5GdxtvvUNxeB2El1Ie9Rf
jMfGJ3PlCu4Ck+7niVsTuH2r2geJE3gs+5dnpr0J5OJpoIRKsanSLRnt1UpDY+N7
hTE1AhiUvKAtyj7A+d1DE4DzoRT9sqXpa0bKrZDHHfvxABRGE6cyUw9QHD3sZJrZ
Wt0SJncGX+dxnU9Ks7rDOgP6+DFvVOHSEMHsO1IVtZAkcPoHtEDNnLc+cd4cz/2r
frAdv3W+56KHQlJ+zBIzaE400nUXFj5+4jlxXihIEJC6IEvXkEZYivrXuyh0AYTx
dO/unmlzTw+JUP5TAYP5LStsEwNNZARUpWozY8E8W+BjmvOWGqutPnc2r68tMdol
kzIKTnNV7BhQN/QGrZNgEdxn0FhywC2tRby9l/2V2tqqMkKOvw0D8kXwH3X5q91C
JZ5UqqUZ2zZOB5bm3SYweHDJ8OjYE8D2km4X3YMfW5+evSttUJ2l48rVKtw4EeVe
QVvLJRUOa+OCB2k8eLpURF3q6IBPc+shbDmsYcB186nNtnLbBSy4TXOAMF7vU8HD
GdMKjk0vGJT/+87wOKchutCRv0eKHlFmLCM2TB24gvb1DdXBoR4KDCuiozdDgamm
D8vxxiV2LhS9OF7kdB5gzxXMVIzYcMuTyO6Secgay5LWZOwOiMHCYmWOQrPko/MV
s2WixUQew/wCD1XuVqqB5HHxclnL/mpcO+9vmll45OHx5mMC5t6P8IGSiKoFODJ4
9NAnyy7zGIXhM4hAEHQnoBk+JXP0GlOQxzabDdYPOFLQIF892OiV4cZTtn8smMhC
jzVy3wtQugsKxDsQ3T9/8LqlTAbXuV1s4oUY4QexM8SK9rBpoh8WI0F063MBb5YE
52mA0BX1YF09CjCAJrqpKayb9zQm/NTQ64+rmK4KfaGaKPu3r3xdM/pwPNWzPD7U
BCPn47Zaw6rY0zs9ZljTNtmLVDpFWRYdWr+UZPet7pfVx0t/82pLR4okNb6eiCBV
NzVKacnNDPvAQ5SeJr2y3Q9ZfJRCGer4IcVe+Rz1W1yNDPezweO8m0v7WroV+jQU
/N8P9QEYFCgVhQMKiB2rSkrhzuVO5Idqvlzu08szHr20Vno5y2Tie2uw8+1aUsHC
7hFgasfAKewFttilGRJpFR00nJLXALV4zGs9+9vwbL0nLX4tJVLIwbYU1jWA9sls
Qpaw5YiSxz6eA5Pw7kpqe8UNwQAbbaGb/pNWEhqHEWoNJKZvSejzblayZP7Ag823
B91y3pCKYbAbjYNCxgkDWojweRZ3QdCiZvBbTHPvqzoxE7RKOnEkQoZPL9E3wnmv
v5SkS6iISOjCKzqevIHXJohTUq3hyB9s+InAJyyLN4Ev4eTNpg5vgieGE2f9k9Gm
Onsz/re2mCUa6jtmhuIGk3B67UmtCBcMs5bL/aIUH01BzAwNg+BYZv63qo0s35tU
VfOg0HzIBWNyoLt04ItQ/wHcBRyzEBmH81vZUFT8zCtgG5BXlh5mhXAC6JYgEwIa
6AE4iFqE5cuWV/5K5vL53RzguSloIxIpDytmc7WsNt8zj21GCr/4asMfz8CrXSQs
4ZTHP4d2lOc9OVPbsDdHPDx3OL5QIg2kogD5PkKfIEUUMT3S6YwJkjFGn9s5dnBC
LBR5LuqZfe++OWlDB64D/rJKIP1TUQcxUgu/1d54OvRG3ZcYjH+ulpZSDHMcYnkn
cOXuQtVFfTnqhgtJIkbEY6TS48vd/ob12CX9d6BmI7hmdjbin3GP1DwCVBCzYp4W
AkupmAvRX8gJStNlyqPKXfeLGt6KVx85BJSUBlwHGlVvqYUZQyFQmAR9DqG5Yfhj
Da79VPk8uSqJZ3O1msDozmkl2/U7ztj1xhsVJZYz0pVFS1eKa8zLK7JKyf6FZ1aV
XvfsgwMMBRmYw04pg+CRVqRvqffHZ73nTP+lhXFCTGbuRRRpbY8hgpUlzj8dy7a+
GoGQ4sXmtUWk79OnDYMpNUrWa76ehEvHWCM5IeSfIHMw3ELTDPzq7t4ytbAQpolH
6SHFKRl8QFuJWF7VLc4vBC5tqIx6zvxoAO/qglgtdLFdTA0c95y9Xv/rHDnW5UCs
zqToJHSQeJIr31k1OvGd+zLhlQmdVVayKai4TzojyhfbPF67XL8je4k01b2nJ4gd
mR6MwqW+VJOfHmp9pQQUdQFwrQO1DhEyRcym/UTfeMnxJXszqAiLs4R8iG5YXsXl
zjVS3rot0ydz9fUafrMP7BxA/aC0JNYeRvFk/fvQdvCA/ivylc5kA3SFwDhnIzJX
M35EuXMtD5H/286PAWT7UWZXoKGileeTnAnln3wf639N0x2PI2qzaYKlryjby0GT
EnR7Jv6WO6LalOrGJkg7NnL1WGMa/Zba6/7ROpU9SrWkx0lwvkfzRZ9nW23rbdJ2
rT/767gVHT5m1qn8Klhz/FioyS1OoK07F0cctqwOqWjc8bmyn8DaEYUBa50Ed5Jc
tGNZR3DR+CqY56DpJcUD4WIqFV3QiydjXOIXAhlOT1cjcnymYpow2rDkKBzcz7zq
bAzjQkgUZ4GfVYn74ZiEcweY77KfQUuN9am+aBg2BxBFwjvg2LHRpu/otQWfpvzF
mymzKSo8Bvp6nTi97BhBZ2gcSXrx/TX2VAf5nL8o1ezyXKnm5027hWF6wACYkIT6
SlxjIAUtfDQ0Rfira4I0RCmt5GvvScS+iUppbs9JGN9HlvgH2NlLKwLI/Rl13qUg
YgilC/h5TX8txt/B96XvORyBok6z5cVVnc5IcBdo16wfS5iUq6xHHX+bWcBjKYLu
oKsTOmjhTvY1Nzw/a2ijpVh6CK92OAXPGOr7vgfwtt1MHJhno//S1MYPbWBbo2GG
tChixujPNLAGc7zu9CX6Mnkm5kjU6EV/6bDv9rX8ZPkKXztkkQ20ye4g9TK0nBdq
sQ06gfxhf9qO9i7cKYf/zYPYrmLZZADm1FRIjxhXnQXViCC6M1ikjAMvMGTPe/sA
q41e1qagKMdzkgMwMf/lG65yT17KwfsRGNNdeM4vALISfo7MGmuCuAdr9ZzP5aJj
jh7Uln4RIAyiFCJ/ifQxaSyR0j7pU3Oo8Ye9b+hCOkeBM0ypZKjvgUdHJ8Z46uXq
+viAk1VV8CC9MMMczt+N0O9XO548ULa+BsaCh82gn3XTCv2V5EZoBWafKSHbdPcO
NViYZJxwsSmfGSzmqVIIxqY+XTI/HcbqlVc/HLPFbsYcSu15TflAmGXCjkF1GSY5
ivzLUrspxc9z+j255aVzYlWCDZqu+pKW9/bA6/pQEeq8ur82wFOsp9i2NBt+b31P
Ntu9KimZgo5PvvnDjmMHlbQ5TjfPLoHspK1o+yAswGNMmBHRXKTh31EnXqc1r9hA
KAR0/0nWI/oqcF0Ostx6loTMrdb2ULAmII5Y7k527HhgGJV+2H0Y38BborawdRf0
8GOxQ2neddA9js2YEw4Lo0e2SNrwKxOO2MmI31+aR9siGS1xSDyf6ZUkVWU8sCmG
smoNw+/24BiBcxVF05XXVHwd37WmCBJ6LXIFldz81sBapFYQyzpaY2en6a3vO4hJ
PgziGFia5CQzPxBQOgW/e1OVdxnPGSmybxKEor/AYZnV0N4k+ParZMDdKQ0jIbHv
T7+BDPYfkneCfdMImg1lQOFDMFTq+hKy4ruQLDg3+aBKpHogFG7uAnTznfMbVpSH
nTtaAHDHgPWgVizCIS7QaprlE2LFkur01uFsaU4pJ5HELgW5pXE6bbyQQ6T+gY3N
TVRK6wVg0COaKNQML/Qr5379HAE4ueB4kymoSgHmY7g3jwiI4J7senmafW1wRFL0
b86lHd5Q6XHFwHBQ92LHOr83DBYNsm3DO/ET7FOG72dQKXsK8iz+2AlVIlAytUf4
secGsFTcvJn4SVHylYA2FUuPFXdi2vHychOKEGQZqEhkhmtBYCrgF/YpMDB1eINO
BPJ8eMmCtBkKGE7lrvMyafcBuRw1Ox1hIE9GZvXJ4Z6Edvd5rfHm+yy0RO6O5/VJ
zmbQ9nDrhuKGT4su4+0G1CucIoCl8gA+ujxFO0YpLDa0jM33GDIdcvTSkJbWqcNu
tjWrUhXLZq3Dj3L6y1AmOtQPnbzSi1UexRsJ3jqMf/x2cweKLeBAR51LEbc+mMU2
VH3dDe49nA1RTve+uMU2vB4ukzuAFehhe9LJc2YQBitYG6GRht63HMCEZ/A4KGkj
BQqXHce8OnY3q06ImvulOp3AWM5ym2ErwLinFuFUoY/Gvzd+dYlxpsge3IPSuOIu
wU21ayf3hSKy2z5PCLUCmSL2ZZa0cYrM3TeaGRcQvZjY99P//1GYRpJWpGFWsbNk
D+OWYZHW56yJWib2iB5HXqMGm+vju7sBY/nfFQYl+rRqf1vwBQJ531JgR+EKgYWf
2la5JjVr7g8Fl11qJP/l5PHtILKERslE1R1ncntVbWof4WtHh1zVUgSyCF+WMYXW
ZaAUE0B91UYtkN3FrIObsKrdtIwz1sRlO25rZoux7taoPNwyqQ35Jum5vXhqOBUF
d+n//J71rvOsyP0TulZ8gsIhYZ4Jdh2z6fG9zxLdTbnNdUXQGixeEOwXEjn5H7bk
Eg7VnAj3Ntwq4R5+/bis4RAHz+YRbL5U+6tFSkn0E6cZtCxbBhvWtJ4ZFpQd48Kf
EDRCj4FKrLgZmx1WCE6CjA1W/2EFOGbit7bkJdmb64hmZe1uI6/fljRNEiq9MJzT
Y59X2lqGVsar3W49VQw5ynokIfIKo/1MFM32hYeKmUgBAL+T8LH8NXODTKeGKBEU
oeCgwo6/HvFBMo4cir0tgX7/VRJ7X+f12zE/hkk1rHBMQsBj6MoUxYupuzTbEuSF
LXZPYTqY/4tc+aTyjcy0o82Srwueb0mEwa/w3c5kXL7lIu3YtVIaIp+mdPFobPKX
vMhihX5gLtyub5Kk0O6qVHAy1KZ1zSZwemSU8FKOQlUywUFER7txfVa1BdzRn3nl
gbq9XZJ4hNLBv8IBhnn9vcjpzLxoczPi82E5JXeDj8pa15M1uhLhP0J4dzhl5JJc
H2BiR2uUnYw3kkjEHCp6Eq1CLMgdB3anejEcLygF4X8DSjJCY9igOQh+SECxBKgF
P/YqkOPBIv1OkehlJkskHrniOb+AovLOUAmpRs9rq6Mxd4emOqVytooqjyKgI2xk
ZXyzXPZEyl7sS1pA3ja1Wv7ekqT887omry04sFpWjSb9k+0FGiuMIx82N0ngH+xD
/LoGgwRjLNlRsUIjW8A5SajSv57kVb44i7l1VAbfTEkheHYRhj2GclyWI+umDBUj
PJMGRwnQvyHU+Ibco4hsJoJu1l5vLD+tVuO2iy5HbKbmniZKVODfiAJ7MenmPIF3
NRjw/yRyFQZNC/VTpk1C/8+n9nuHFpkKEbOrXV2zxCBWNy/dD/CsAWTHGO6sZ4xX
DDUmKTX8FP0W0N3wWkjq8PJdKmrLtd91DwOr0WKHfQSB4lZmoeOg4kYRJw4H1wCH
vRP+Rd2RUuHliCn0Oqtg1D2TF3mresstxZZtyzw7Jot4dZ1hro525yPgFEFo1qoM
V1xg3MsYlEHH6Gp2Z+97nQRWvcaJ6CkkxQR9zRKGJCbzA5zd10q7a87cIAr7zw3m
Qto8WWp+Aq6dpm8OriTvMB80fq2U07JPSWVTD8FWSZpe982L9T7BGtogCgw8+uB4
s/eSxI/goHJR1UcqaRxY9HGlm5m+J9dwO14xrGXxY9roJzzomXyGCxoC4q0Ky11H
iU5PW7YVqP0zIpQFASxl/W49X40mI9cdjrEs8tZbgEUQUIHFfkUGBADXp3MUh+Ms
RgyrRlrfVPF7ZHtgjTZm5v1s76Dx8oKPHlNKVChjbg1D6qpy2c9ZFXMJllFPc2pC
leqTi9C4j+PJ0uTP3cWrLlAA9iO1dBTfLzxMg9793NE89dOWhLLlLWXzIHb7LDVM
Xd82yRCfatimDUIUK9F33xZQ9oUEmTzhgaXncy3SfaW+wlExdci1sDUJ5mZhsGY/
mW+aKnI0uS+qQsaRDB6lITcpYBVKwV/zvjSo6pdQu8/ZvR+aulYN72Qao6Xx+zJq
IzBYPiA/xIetam+2jgXuEzXQaL9hREHckFFTPJ9Gj/ydpGPEoeOU+heoM02Vr81z
LNlvD/Qn3b5O85QIpjoVRTc+tBNofET3slr3wGN9qdS0j4xwCJHb75+HAoGxWWix
i5cjWuOs/VhUPQgvJ2TZN1HKEBs+z8jqFEamXteoUTGRZaY4reppKX1H5sBAFgON
zJSoRzcKt1fxqbvBTL+1jNEEInk53WTzwmconFTVq4X2EHQdbzbb67yy7d2+I3C/
AlRXND8evXfvPZja3XhR8bPf2ZryjfJlSyqRfxWhUMrxYcIzw7FPhemVt8z1pey1
1BPLratQatKQspqtymb9H3zkBussY0MzqD4dw/xfhVvxGOlxoOQwbdqYkhEdqAca
BhaonHNUcvCqk+ml4c4stGI8ohhJ/JB+2Q5S1YWrK8vc/um3HBLIUVzTOachODw1
Usb1z7IQAE+3kNaHRXGe7dlCWMfJG4cPFxbUGDvgYSFkNyhZCkvP/qzaAZcwGJRR
hrtdxgrig1M2nS98+iPZxV8iJunyi2IBdsKiJ0VpMdJMw7MfvuupxkmSpOENeFm1
9QCt0OPbGBflnb+DE0Y06Bg7oMos2YNNe3zWB9gcKl6tPJCnGNZGjUA5Q8mt4+Fm
UCYgsCv37Y1e0WI2F/8LX+4LsqfgR/KFjUnF5cXi8IGGk24bS88+ksnes9OuATud
Kx+gdF5FnuxvDE0ITCGGwPQZlC9TDXT8faZ/OvpCEwlDN/N9MNeT5jagCHiXOFp/
XT1Os5OqIEWejLL7tnOaop4Nzs4F0Ke1kkV7FCdKH1txGM7+Dfat3FEzIcjgkfVS
YywjTg2Hjm878AhPVOy7g8qopgK1LndqSqGxtlmT2JKc7tNbVN3m7ihOi0+EqBgQ
7XoozOPud8gCspaaFzoIWzR8BITqrSqavQN+GQukPy3RYAikHU9eu3hprqyyW2OG
+zkCGNA6uNpowDqAiTkBaz3+Hd0rM1/X68NKx6f1oPWN/b0pVuLDOqzMoL0blqn+
oaAKsq7Rt5V2YQQWkDhW8B1tRPazmQ4ZrhAg4ZKfa3w9pWyt5mFuJ5CcvJE+oCmu
vID5anz6zFJr07WnqPwt7v8kDzEILr9EzjDUbSzlWsk472bQv91AglAXXR2ZQwU3
6LlsDZLrGNCkbvlEN8Te7oCybBjPy3NRvApGXUmgkFM+scoCBVZc96AY5WyZfisl
/5ymRvTmwoqCJuG+S8K9yyyyv2LFTThPtSE9ap6mOItvtHAh/icKDtSLzKPTtvj6
7eXJ0qoTmX1Asmx/7ICW7ayvT/vLbQ66vdbq6I9gNdZ4890hu7d5b+GuQVHDNbpS
gt4ONm1A6xpnk5IqS5pQQ16XhB2HxB17yJGy4uAu4ub6nWDR5rHVmhMwzrBoh8MC
1iViotDOE8E7Bq/1s0stju8iT40UgA4RAXuTAnrSbkGui2KSVgpnen3gypvN8pcH
gUH8ohkfVSzbO5SGF35YK+i7Os4jWc0c8JfFZ8ng8EAezJ5pFZOBNjoHDBxoHCRH
89U2+ut5+FJiITzDa3C6EKEXdz8AwsFU+0upqNpks8RMxBV/l9hsL0K5uBseThR0
+zvuO1YOwdwAyKyESiIyjw0OnkNsFo7kc4OyfZTfRBM6S14QVPcm5KARwHRAJJQf
4gP+CCV+VBMR4STPmJ6gzgTGYCwkDKpYpNMjObuK3OoUszKmuAPRXTVLRh0QOPVv
YAHHR968609Qk8uLVEHTW6lDDYqo8MMN8LN4l4bYGCH4qnypdWIkUAb4A5Ip25Rz
6xbbt37Kx1vJF9ia4WhzCxjAyNxHYkJxa8WF1qC3ZMjuGYBfPrgFiOp2SK8qi0/L
UCXdsAK40KeY0nuKl318ZX0iVJC1fk53s0IEEzto+RpVxME4eql+P3lQtBiHAUpD
h6SbLICeuCiDXhQTCoEqZyxiq/A2+2kz9dhzu5C2RBOudF4P/qbkP2t5PwF68pS2
Gul3jgjj7h++cETDd6WVVSM0oJQ0iLPfQfyC6Z8QZq89eiIbnZb6sSui4NOBOWw2
qA1SQZLkz1z0wIVWxErHSJ4ubcyScKc+fecvojWp4Z2J6sHI/TxBf9E7FQoiA6FN
ImCR9D0r2OImriIwG4kWWCDsTz/mWReSI2xWuxC3Udc3dNfrpH7wJ3NJ2P5AzaBT
dKzrkFXLyxhOyV+/6WgWBvhOLAe/MZG684wwTxwnRgCh3wWU9yb6L3Z1/yWVQhpR
EtXDgwnRqDtIXl8pwe+OvhE/wVqtE0Sq11pqMMEJxwT9/upYAG4/AkArKAcJbfkL
e3xi97ioJwTzbXsI/95q7sb3/N8Cr46v2Uj1Hn86ZBFJJZXHtIAsxQq/FovQZb4r
ax5iaF6BLWLwLT956SWh3+mu+cDYQ1+nFhvBmINVA+6TafHOkM5bIGn1oHplA8WQ
Zh3aAo69JYPrWEFAYxrdNlMWP3I3Meqk1QFTitAUwrQzou1bUcW5+VoaED3mc1nJ
lL0sy9lZnRIDSDQyyKdH/jSILMu7i7VLfVuyMcvyxlWT+PT3zF+bVagy0lv3qGse
9qeK4kzNJdLBVCG0pkS3ECkAC1SyUv0YbjtK1uoJkqYG84Oz904BgYye29g0DBRc
L58PolIw5sH7y7ychGhTbp1BeVnM9z1e55/3bwTVTrI1RYLwjZ81SHfdRreXLvYj
UVn5IZEjYjlDSwWus/2c5qbp/dva5IBOPQaOri/Z9f1Jsmx9CmynI+YPaqtacVnZ
aKP0gUb8PxCkgNuJDOH7dUre3Ly+q+czOUgHexSNU+4eSA1lWuEHc2ASEGuqFPfE
sVSoVj29l4UynyVIgRGfDdhyt5VlykdF25X2YDjIGolNOyOYe7gOgVDCcr/ITG+C
Y3qeE7LexEGdr2tJkIZlLWk9L6WOrbtwGMNir3yV7hncBOqRuS8zyViNlhOtQ88g
c3t0Qg8+3w8+3zB88UC2F57li/ycEZI6/GcLyA5c+in1SdwrBsnfqO+Lb+3YzcnM
B9nlDXlcZ78kMgm7sFz99CY5C+jswQJqS33NyoAvILRmligFfFitjLb5RXq8j6H7
6pVoUTx3UIjG0BGOCOFGi/CInydIID6GUnwXHFuPFmdjrb1jmC6Rp3k6XySmqE3v
KT9eZOezsI4jDNwIQbl/B1+KsRhhk7NEXWhVlu8oRMMxuYM+yp8fYdp0QWnGBRui
srFm2goVC7Yj/620Mtq5pJUte4drdVT5QAMzFgi8V8JM9bAsaWFmShQeCWVNbdB0
dT7HgGiG1irhB/WmPAFoKFNaFNz+MMcKJMD4h1LC/Zy8+2mwXfUsgEziwnwSU21q
iIEJQ2y8AOKbILTPERRtOzqnaa4Y2Jg7RNdbT+MufS1i89WBRcvjptoNr6t6w6Ob
rYnRokGNLz7xkGfFYy5hZmEGAA8bSBkOowoZb6bEAmKn3UpAwwnBstSOjtPO+vPB
O5wP1EEhSXZeO7mR6UPhofTjpdvR86tqwhW6uynQl5722mINHAfcb9HYboYuapvm
93lYgKcmNask01VUwY3RngDPO0R8Hw4cLhZ9tAduDvjNPfBFoZUhCtsMVqxndmiC
m5RkKIactBqgb+TAYBvWp+UI0Xy9jJb15IVsT4wM6puWIxWmRAoduqnDIHGZYRCw
3RQAJu7oqAy11l5CiZUms4KHBYvtpg3c+qU0JqX5tBiFagX6kGdOK/ZsP+r3j1zV
Q7DvtFRdWDvJNnmCT0btydEYejbX6QPdFh8j3cSkm5I9+NMtiDreiNhpjQUVrn9d
ax938VLExviX2gO+sQ7RyoGsLucmFc8ERe60OA59KZH4OC9ZcGZ/BHVxE/9SGEnn
0ecTaxfzevbo7c4XYmJwMPwGLpVyK2XpSWWfg59E94jJQ865qPE8jj0yki3qbSlH
Uk5nYNSFFtcdhFP67OtEsoiDUShJAsFK+2gwpxgZEZC6aPxpgyVEuVeQ6kKe62FA
BcY8L3r2X9Qa49m58YsNxIiz8uoIAxoEOedQgvTjnA194tVcKsb5YPMSyk4enAta
QH4Ad9YAOs6fOdidxIv3BDRowFR+AcfeAArIjH0/cJkV8Se5k6tXF1iJQOp76GY/
s9GhdQEme8E1wRRx52hj3k5zL1CTEFZYiFKcYCTEFhgEMf02Hn1rMilh3F4xzcBE
EqirVZpL0ckEQO+oFYPdykJ2IaA4KVjP/Yfx8BPJVsYr27ILKKz1I+dpRT43hsc2
eV8J6JbI+hI1pWhdOeuumKYlurWjYP+JOQpna12EQCHlac4iBu2XRBcBlPpkWyYm
N05M8etvvkLlnpKF3GyLtRfazy/t2Eq1Pd/JQzhq7RNJLEVF5eGH7qlCN9tDgwuY
IvyshXEgkzMLwpl8VrKudAILv4wRnx2rEeW3INp88Ct0ptDLOBHBSNF+C+FiohFv
Z2uITQD4kerWUxVj2hZEWFvXpgf8oYSuJTN2QQLELDywtBglG79NTajq09xGEaAB
2GJR/0xXdp1r4//JqC839JiToED5qL9vYUb8c4pySWdI5Xo0KldpfQ3jvnjv1bQP
yMI1ihS6zIU6yGQd9Y+7m+L2Y9Qefe47brC7ItKi+NqSdEy0vJbREPyr4Kp53HqV
Atd81p3wBhkEYv4f+EASnBzVj952fUUG8As3+ogxnvbvuNhS04Y44dpKF9hQiTfs
reA4HqqOqwfIRg48JXq0tE7LLURTZyibeDl3TwN9OHvPzmG73McmJ1F6Llb1ANYe
c6RG02KEBmPT7jz+F12ozlBzIcAn83Jna54/8hhkWdZWR95Yb9ncBN1zk3a9g/c4
z99gU7mkZAxGhJseVQRGIRcxHFOrQZYXLR1sDHmDK9AWqqnYdO0fytCHSUywN1VT
qYdd7GOPsRt3JTRBVYi7rrAshe9ieSqU34bZegXvl3qkMC1FBBKR2ke+xhE9jTFp
XXCs2zmmombg5lKf4qSkljDzY1WnCAjnjazHZGZvsj+/cNmubY6u9X74RTs7SNJ8
4HvSvu7hvh2uiydO6/jX74cVMzxiJw5+6TzR56fr+/fKLyR+MiU4rvbrdnIkAgFO
ZEVooE1TcUN56Js3kHRIptjYhq7Sbf4TP1rXgsm56KuWbc+PSKMOaWQTVesjjARd
tm54HqmQ5VPuGUP9FWkRZxQI+VxNBrb13z9DaZ7sHhgtL0j+GJ02H+g2f4GlNs71
qE9Gl1BiKxUsi86aAWzBomgqgIvpx0kb2VNt4Sk/vwvBAmGmNAf+OkSIUXz8LY/5
pgsCkEVHzQbpewaQy7yvC8+rn2PmYexrptF+n6hFycA0zBau8CmaBLm2lqLUOyIZ
ZXSY0d5UFPGEimee1XRiybApo2RM1pXnE/wMj9BXxHbEmhKGQJux0lu4Nao9VgBz
RslkiSndXvn9Xn/sTjYKN4buVRtzDlSddiROmFDgAbmgVJ5GgFZ0HCi+ySw1CYqE
3hE8WQ+GobfvM+vyLbHNNYfZSHeOyDE1BjepJZwe0cXk57i7jKem+xwOJ3JHvrAp
w7VS8kuXUbRmWsovnd3CY2K/xso7ZWbxf6dlzZBVM9C+lStdugVwKQQOheSdV9cu
zeTU3MccbL5StcB/v56352bLgRo4hOgfz3oRKvpLIXan7qfeFoLONuzk8pc90F8Y
sXk+sLWXiQisf1bXRu57RJDssoYLZw2T3bVm0OSPuRtp4BfrLOzMrYIshsyT0Lw+
sT2qIvAeVdg5Ew+xI4ReSliz05vxM6ngwxG34v6LhvhPtgKW7wpK0t8VhNV2vmHe
lCDKR7JSXNXLWikkKQEVcPNgBEioWzNCgqPBRPnHSPGqwbjhsXaKfU4dm/ToIFCw
sK5+97xmxbrYUGXVuEC7fxxumSqE2iI80Qj3RS81bHnQfoR7KUOWAMBqwslymAX8
UOd68KvkCMG/eFD2n+QsT/xJnkwi/nEsvholAxb0I+lp1ZiBV92ZyATLMpGRgJcf
psNP2kr6TifyDTRHokRg8TAHkk/H8wS7UfE29lbycvOnZhdzetUn8EuU3i7TrfAP
yurKp+dCDsjg5CebdD+CV2Vf5ITaHtAILaSsEMF2DZYksMoLRPT7XeApNisXOSz8
pVDsFIw3zsR0MsHiOodzoDZXc1TZ/8mcOtH+XR8p1HYGCKM/favqWGwDSL+NuIBP
9HDPb8lwbP2qNtzMu+gARL0KQXTs8Ic6t01XAaiwaFhbZFw89MmxNPXe1rzANnfo
U7tpsNYlDQwzeASPnOPmHy3hFzqQV+IyJ94xBcMgY7sM+3f3Sq5ZeP5x1/mHYj5M
iNmbd4okx/PKTFd5VQWw/RV0IhGp0p0otcte5KjyrOWHvI67vOiBeJe0ZYHq5E0H
jBa977cDNC4dwRYrlNKFSEsmJ0OJC58qNFk3r9ksB00fmT/rfVdEhFjaWjvFykI8
MMxZAVkKjv53dGWSaWU8iSnTy+Mh1hv7IkXzvC1A7hYmKaa1TCwWoIqk/ut9t8vx
PvPdw3ULxveBQoGMJrxsMOmAgpb8881QTJ+GwPeNLm50njZcTp+Die0TomBlD8f8
m7cKGN2cWqcIlMZmX32cO2NzSP4B7pzwyOVNqV90WHtjriV7mcwDgSe+JCDjK7iC
WP1niZF6Qn1WS7adS9c5gKsZFPFZrmIIDV8SaJXQLQdeAnVX7TnKegWwPp14hRGa
QtfylBmCmLI3e6IfcrLrr6VRinAWlHyb0UjVGKTSjmriP8RXGw02CvO/PpnLqRTq
lDjjI8ab+abCXyB5BLSiL9x8wUu+t9sBSx6HpQloasHH38fK1UpoCtLhWsKt1PdC
hI/DuwOxKhIo6yXhlxNMrq/g2FbBt6aRqyJj5JHdEldyCcMxi+FrqmDI5CrKtjZq
wjBguKyGtwcwWqoOw7MtOnomlibVaicZAilys6iJgCzXqZqzP+OGqJcnYDy8lUZv
yIAa1O0vd0ffu02wpuw9BON0DtlASdDrfcqJHnZHqYLVoYap/m7KSjaZqDuUy5fr
wLGugOn44xVD5KoxA6zztKOymLr/gyTOHk+cWSdUZFILybDxZByKyPEKQ5MljwO4
ymzniI10CiD3gIXEVcAgyZ7abnSWSmbzC7ksFxWiwqZFUl2oYiATNgDYD/mg2heD
IUzR4rAxsDHHBTZdpmYWk1xXZ/OMa7qlb4uQ6vf3jMyM1PfYgJdBTJDLBrovo1dm
ee47KxwImjozT7q19wL5CNIbQoPNHGi13YlM3TakSJrGzao6+ittLsE80klGBCVv
mayEwbGaqDrT9iBHXoOtLAQU9wYwumfBH3zeBqh2qgA8ES1znmwxCd+BbN/ncWx2
ZJLqmuC0Hcgu9Zje5bt015o7VVmFMxe5HuhC7lIzgD7yFfBfe2F66Auv4Wd0Ngs8
Za5uK/JOJo+NeP7O4DxjK6GKQUTPvl4eD2dJlbsDZaSPKzhjc8FmenEPymVVuA38
+cxLVbalPEU2sgNNYVAs7C2ZDjCi6kF/vGyI55seWtguTli/5tDlvM7K86nBtJP4
KpYOQgKQmwTEWqUfKPoLJ8Zy+NNOBs+V95eC8SI9bT1h466zO9WapDb7bNVvD0cQ
iXYTnfhy70ZdJXonHYt3oURCMCCfAsu2y37Mg7dYyWnNuWj36cukRX5rRwfvjj/l
721tCJV80lMCuhe4DefYfKPOs0bOaE0h9r8ej/gs3Grw0zpcDC8rvojuNlSrXZ7T
mTfskyhwjLZiUZoKyktSl/wWMEHV54GEUnrWqZlmJ2aZpJcUarj/YbQOp5UUX5E1
rtxSmXV5xt+ZRl+zHtLfiXGxgpyuWhA8U5PfNKL9ZObJE3ckrdH137rqkC00UTp2
tOy5Wvgs0S6XkIDzH2iL3OkdWb21Wz3TOgum2FjWIytQ6CMqqrc4EQNXihj2r90H
spE+Ifd9yfFvEiTm80qiy7wOaUWR7y8CBWtofOHfqFYj6lemU0CggWdxVg4rUU6m
kOuLwjZn1LZ0zDenoVK3HNIRxxMBl42C1CnmjILFhTJWO5WtUFlepYzIEWl5Ya46
2grV0zwNdc/wiRGxj4d6ppGjPakVbxhGBL3nbATWyRoELCsTRTZw108Sd9+OQAkw
1KMZ9vxPryT2hasc1NbSFXIL5sRCkfsYB/tINcPFJmAP6u8jTsADBvg0VXyVAbaK
yvgTi0knFpvm8yoUKyZpS7PG/kxg2hTZo2CDkJTIcRPfz/wW8YqdIY9EQgl9bFrU
238PA0mCf3MXIBWB9+Fwub0VTvcASOMl4yFv0uLftK7BahSxeSXrDeJvyPEaYkwA
J5vr/FV8VKtjWF3U2nPNSwc7A00Hdc/zlTFyzzZsqKv+5gMYvIyX0xK96K93fwIN
c6IQ/IpQmClqxWjcsET1+tKp3+QNcT542rM3VIUoBYjSQnT+SxY67qpM+hEXiuzv
IdMXQ204+SO6mB6SaJ8voZM7FP1JUhVE0rfBNyEEBEMd4X1UHb+AAQ37/PCt4bQ9
5v3rous2iJCb2N0BEWmKOeqBEuPix7bfGz5L8FlTrB9mmZbVOgP2JFGq8Yy1SiGS
PPJ16qhX54Q9LstvgKMVVeVM1PHEfhY6Gx3o0nD9Cefw6jXA0a1bJcnRJUJeA8Gg
SlO7kVWN4WXcFa4dCkym1T7lmgS8XtERAHEfDhtX9IetWD4Crb/cvKB8Ij4XSDde
01KD0LkIb/fROT72Ecn5UerE9A4TEVERczGsLE+i5VCoeT46xPQLmM0qMUGvUNl6
Q/P5hzfAesEYK3oBtfj8CRw+3iZNLnsUCXgYyJSnO68G8rw/iXODqae5l4F4khCN
1Mjs24ZnsFBzN3XDYP1DE0dZGTmo1JjRTOjwZioTixsYiM+1cC+27B+Vwjs943uM
keEQ7VVk5TvF+gf7RBcLhoBOTQ00/9fD9xQrvCjMhmoUhT/N23jYcX2LmiP6Q8rf
AGjuRvo0cifB0HFp85J+nLAlBIKioQ/5xKCVV6toDZwDQDIaJx57VvfY1xQIr7cE
fiz34hZ/q4u0CsrI4EHRFbdzg2fnEumR8CKbXgbrSAkhEJOvaLqL6m9SVh/yOzCk
ZTKoD4wc4UB86BKgj8tTm/yuqqRTDi5V4r0uo9mbH4LC/9KYuzZEPZ1b1/VjJ6ns
O5bwsuk8sxQbFSINLl4CAaq6TrGnscoU+owNCD9YUKLkG04V8ZZB5G+MVlMyO8dW
69MgGHhLki+nr/Xr8n8j+rCGVo2Zdh58+ss4xd/K2Tl1BMlgwM8lkNbMXraI/b/I
R5l3Do6l6tLfyGo5/1H+G/0lL9GVWb3VSQqt5xunOS5d2C3bKZwXXyB0mCkyWakJ
IpWWzMdvJl+4or1zWCHWAQ4ISoNXr0pkmgW/iPSfrc3aTbVeSoDxtRs4XPL5Bh/2
Ie/KndunbLfVizz6nnCARWcfgtiZEyQCevtx+CAEHauLAKTHwzrnbYcwN8P/x0NF
Aq55UKZUPd5I4U8cpShgo82PPm9UYSgNsEwCUTWGp3kRLiBjwqn/4H43JP/6Pp0o
2jRONQbBDY+4SICbTDCmq8Hoz4H/86ZiRW59CecZHBKk2DGiPlhiiFyEj5oyI7WC
Z7OBjMhf1ehryWc+9XZE6rmDJfNsIumWQWJXDqlJmSNh/xBieCJIvxQIqOVDd2us
8AKVb1m3CJ3/XVvBgezNI8OGDIFOHA5mwJDYRHjr1rVnIAqeRZGCT0O/jOfe1i3u
c3XRZ0geffmFQJf1OM58/7heGx8cUAAdGc9gu5HE2qSfPcJggrAt7KN7yxPM2920
ipmo645nvfJJFfAgjTiVstA+F2RqL8FWX3T6u8JwFd/Vv49fCK0n3wCPmVc+OWbH
H2q9CoucnnbWDLOx/KC0O8U8VZ/M5hYcPki+4OXI9sKYkdtT0ov3OhioK7JDsxax
8lOmYfk+eBk7JnOdWIqCO5KF83SZelYgVwn7x1nSx9Kj9Ei2w5ts9JBocbOw0AZK
z3Ad934QXGFPUsEbWqDAWZQBGZZX8a6keHJSCTDi63/eU9KadmrGJuuQPLnqYxWz
vnvLHYE4kM3PQt3Dl27QiQfaC2m1Ez8YhFqKDdftmbccGqnzQzmLzBdaBMG9StSk
cfPLI5DN70SpkQewPntdcptnB5f2Zkr6bTn5TdmPIRzRwZxID/8t05IxaMaUceWO
RswG5Wg3tvIAmYvc3yt2lO816BwKzOW60Hx8v2cdYRMMYhi88uuL/YpSCa+WD247
HDMJucGe0NpN5QxczaXMYNh9a083G8v9rUjUomtPKf6cV/rHKK+TTLAFH6tyynuW
apJPibv7aBiqhbSwI2tfOm39obkFBTwse80uJuZSaU5FG7o5nSjT9ki+HGoHGj1y
Akg/TVsVFJg/j0exqHHdcfef9cnwcWPNefIgHjwtEG3e7pAQUDrbK7mLfL/ifxc/
UItWNfT6vSShMZqakim7RxN1LKlvCjP6pZxF5Q90kEYob+Btc9WnQ47hl+5zHIld
/Q4pvA1EWL2UYnZOSILa9pRd8KK7qki0OsSg4erO18UQVN4DZmI1gJW/mHNlvntV
xVoHOfRBH4tMYOTFc58119KBICEvcK912QrKOtHJqXDOzJmcGwLaPLR2vhYdwx6P
29bIulTtMJZDZ7L1rKm2blK2nnyWxk/CKs+5r/b5YjEdBirldDffwfBXaTXAri4R
7yV4Hrm2pYRH7V4Z0M8p6QsU83cyyPkh6Bew84RS4mKvv/V+pGMp1S2qD+6g8+r+
plTLkXZq/4sn1U/N+yNvgHCPrV+eRu2M/jS5JvGV07yeAjbm5fHN0/BG49a9Yj1p
nCo7lwP/AwwUy+9VNlEFE+yY6+WVwONDi95958/TjZ4/wkqQF5Eu95fxiDH11+2y
k84LHskkymw9CQBAjpIgggwAijD5ZvrKw/GEmKY74q2i+a6bJiJw7wCo8TwMOoxj
IgQ4X2Hv0Z3KbAs8npxM/BmzvKAc4tSiRcNweapzJVHK481V+z2xH0k5q1Pvt8A3
7M6nhkyXm97YTiq3h2aUXHKNgOoH7h06Z3u0/DuiRSIhl2rHKMbZWOvDGa2eTTDG
t40BoOCm0XBD9Y6YNZ/kjteydYFKao4xYnp2QSI9pM5qleHgVS/FLQZ2Zutdv+GU
BT90exBzWx3rH9XmhVpjeuhPHe9iof5Enp7CQvE0piBjQ0jAhKcl5cZIlIdBILwZ
WvtGXL/3dmkfzpKQ6Ma4enIR+T5yZa6z4f3sg+4M7rfMdQ8z6+CAEFUhChOum1FV
pY2HYOUW1fXQiaZZMxPIE/yeGKQtd3aW8T2JQZBDgocxCMK9pnGHH5RIe6vUjLKO
+UToEXt+b8neOCUr8zeVVXsu+Z+U7jU96XfXT3Or/D8GoRmyReb7CHSNFg5Ifpns
zakikyoJBqpbD87fHrTAQMv+xVEaRL5mSyrsdasSC1+tOSgeXVfdo1EvtPdQGaFD
eNU+g24AjNiJddj7PFdD9/tl8G4quBctPATn3hI5Skt3FSOGt8uf0BrprxR7CjfQ
V2G50kcXNwJoCSBwK0VIbZqPZHnmjj2woxL8SVnqVQvi3CHYjHr+H78Tb+j9HUdW
x0UVEObnM1ctFr274rGsOPO9W7BHnPi5GdoA56nuxqMS0zjWKeOrcyFzJOmq3f+p
45yNphn18o64n9yAq3pUKV9xj9U/CNdlF+MndcdYqFUY6vU/Z3pbfWZvt+mu2hKG
hCpGw+1HtJjIaQ6s0IJaZenZhay7CG3hO6Bz560C08VFtmngN9dbECk08rutwVGF
eLIGefhKpAyb8P/SIosHz1lau+02lKYQ5PnVywhZSH4jH77ghJbfLwIMx16f0BNs
e43BHEz9Jx+WfteIvHbaasF5rmMSq29D7qEktmMZWlj/FMagwWATN01edFONcdIF
uyJJ4Wo5mksHKq4YfyPoe788YCaQJG73hq/f7RBo36ReaJ1bSLzLday33w47zZDX
GGOsNy3n99pJlvJrRfWTvVvOFHFRUpZ9xbkh7STZsvqtsRGwK+CtV5KmyPAEtC50
AGG2q3Eh21v3qHgwLoeb7LkmA6ezGZYeXF1WmC/SGrkG6l8PuXpJV5D8+aKU9jG7
Gd6Go+wEqJvecfPQLiL+oTJuYLrxvfUlcNmuoIoxw5SVc0H33hFIqJGw7YIJ0Za5
B/zeI7v7vF0f1FCLbv2X+JJMmeja2owRT0IvycffcUT3hY13ZU0/RMoyiXfNURV7
nHCSl8XMvq6bFLpsjLDzH+94fUeAz7o/Semeo6ufpyP/T1jkbUXZJKZ37WYSI7Xt
6kShpIxg/Z1KXlK1zMnwv3h0cqWdm7vTo8Cg36E8+RNyc6LuoMu0lcDAsJXBr4vH
D2hcmihlW/KTF/OZVdEmF4w7Y1KmiSiod/O0oV+nF1AmWFm6xOoIYrzJoYOd+crj
jcMmQb/RuAN6K9TqtHdJrBVH2Z+F6aLYlNa8lxdi/d1qT4oDVQFaOXsStFoFdX0B
Guz259rsMuBb7YJtWSRXHYKZCnUb5o/elwh2JjdljxHWhwaF9orAzk6+RKuclWNn
JfEF+iBMvFmfDzR2knbQ6iX/fUxUBqBO4t8bUgKuG3pwcJMj4HiY/qLYIiJHuUAT
o6lXIUFNQ8kQdgrPaFuuXix+LDMiyTR0zl+VDe7PCeI0agirVrp+0lZvLwHHuU58
lYIeFjOtu6IURipVOVhH824xTJN0JoxCQgzpSm1XX73I8lkV8tnnDXLSaEc74hra
icvgduMyG1uWpZFNfNoRWaVolF+ZNFnuBSBadSWQctoVgqxml2CfoZZWOMvjVDQY
Es3i7E39UTirhxmmgxYeNTITrWT119zn4FA15mYIPPm4KSWK3Pdk+I/ggv87gBco
v/9nSE0WoMCfO3ZpMpNJQUr8fOziqQQR13sp2jrXCI72BYCpfj4dikqyJ4Ii+2yy
X/vRnsSQ06YJzd1m9pLpdQXgm5YBKzKqjBJMnZYtqFIqWL4IMDiSuqCH5ezk17sr
AmZrB/8JM4x0FHWdT9IB8vuMwkCsibIbMXMvyvo1YT3L2xMfnL+mgfREbAk1lSnM
7sbf8XYfHbPcHvva4K265j64LbYuE9+iPznFhpgbLhA45mHVxysYIXKtdHQbScXz
xEab8zkj+tuEA/jkNAm2AbAfmhkbra9tKWb9l8GWBRSAU6MjbuyyxXY80ZtFaI16
OgN/alte+s2hqCKvk1cwKFxoWCrAOL/hwOcPpOdALaoIkCqBsZUoIUywJ/YmKRXI
uiJ3gAMWTYLrfRzsLV5WjVIdfo+6yPqmOBHwYuIvWAZI9T50SeQF1bzPoO8XMPEE
ipq4DRQIqd9VrOkpFd5X8zrzvyV6g9ttrJsit2HI6544BOrhCYXpHhsrALv56Fj1
Tf5pOjW7thLKpuyAJZa+4mELhEVtOsOyp/b4bg+/ahBFBSMUBVC1+1wtLLPqixYd
eXMeHbewei8Qdiw52osETjP9UVYRdFtp0cqcW2MscwLTgXy1l6q2MMQvuGJBHbvt
X8YnwCkBV0xnOT8bAmFHQGcpnh9eVnK3C4xq7sTRR4yY+I/WYA/2z3opo4qHUQcP
RASZ3btk6CgQi5dJm1JPHKR8JFwiqavGo7HvaeZryc+4DJ2MnI4d9AkAynRgrlAv
1C7nP6grtQZzF5hxlb/2IfGvenU3qpbTuH4b2sCdSAXhmF9JhwhjrPYZsX6TLJpL
dBaHmw+RWLLgWThewl6STuy0IhuaLffMujlFdgaSEMYl3RVqRxx4Yw/iWP0x8thm
jo+SaTxTJWK54ewsAhwL0ikZyVcdDbTG3yWELjRr8eFKFjR6M3FSmRUVcDklTQgG
d33zxu8oVBpsUTQPugWQiW6hA68Aw/QV8sxLbrgIdqdoRdcyN36USSKb1yVettWH
+MVEOz2KHrGl/Ql6ShbDx6/KsXVK5bMG6rNa15BL0tKJF2Al4VVQ3D6t7K7l8kJI
xyefArsS+SIhpltVQrJqYAQQOsrx/1rOPWTsZy3iDc79ffLGspo9A/Eor9ZOb9xv
ZJ9XWo/7b6h6lUtYK6NdAUj/VqVdiPqYtfrKPFrzuvTrBrGOMlmwNJ5E/1IhcnVI
C3l6sCOo+ab7UR4tsObc6+g9iFxPACYK3JP0ZPVSOxqzCWxfPM8eVhaXA8UsD8rk
lDhpggkrwN91tIwsB5PnGGnnwnQinIGuE8jbFTzMBt48cHCeux05GkHpEcY4VHcR
Du6AJYi0XDngqUaX4p0JUZLk3HESttelZZ0HcJ25zF0W97x0GFYDcV7OyNTgaHR4
53RSDQPJeABqWAOLTCqPEP5boXVaQHSq0/orOgcOhe+ZNh4270emNizZElT8djc7
oc9S42jzPVz86nSrJ2/UWVZc6k2GFtU2P6JSG/BrXt5IDvaZGcpmlD9bWn6Hg7EA
hfyzJKazJbsITSmGdHi9UnckzasDcparpGy3F1bECzgZV8Qqg8ozOV86Kj/BY73I
NZuaLMIgKP2jXWyPovGOiwfgVkDU1y0ZN4neKiR3v4sY66wq2+lVTKNR1JBB7Qev
aiapE2lQQ6M0mOrboOz+hXYD+6WOhV0ZihThmLpxUb0xYaMgbE9SX1Z4kj9Tq1OS
OEQ7oZwwb4m64tsx0jHiMrfPj6gSqO1wisF+ZeaQk9YgKIKlQ5DjB6aHZ6SR+NQy
hm4j0whXL/0e0jG1JYeUC5YfgNFCMvjeh13zeSDkIKQVNsC2MUIq+EGd5s5yutqC
AM1jtiYuZNyfTgLOgssE/JRyVT9gzfsp9fD0/JuyXkJk4OSRNVHszAzumKGwBjjQ
rv9/eLH7Icq2F0bC7vxqgJxU1LsN7Qgbs3I39d0N5FYGhXz8l/oj+e8Wd9fG7xLy
O4qM9fIbmi2wM3Nq/i7jFUhHBAatHCXHd6RUZVDHwEzCqtilr9xWYhQEzioMyDqT
RGWvKg48cKT+vcormOrvANTDx2I3HF+T56joI5aUB77fzB24RYJ7EzLR7QokTCjO
6GY41d5zjiKudpXAUJDTO9m0PCs8nG8uOqalc7Hgdz6NxN/dqGCIZjI8gSWcM8TJ
Vanoyku5S7FhpIEyt8yH4WhW+LvKS3ZcT4gwnhlna8EybFC95j16siBxAakPvBB4
ib7sqVeixJ1T2nxr6JYLOYzzHs1Gd/3FmkCIp/u7wogvMv+ObQik2Ofb+Pw0LNJD
ihsJJMLS8Mp9O9HQp4NqfQTgU0RKfM2wRxNdbZKVHPIDvQvqyXfWCsShBoAxiiHr
Gv2kPn4BGG5mbvObVGyCydtmNbZu1X2ln1+yWODRmVflkD7NQBLehYHmZFDR1uxc
H/1vhj7/Upbg4WaAjUZjVa7lDXVu6/v/58qYRPF2B2zhtUPp5HEGnQRrEtcCvxOE
rtsI4/Y1yY+pG8yx9VNOSRh5BfctgwJsKPajrm0ZI2jQhigGg+oVFeFeaqPToepE
GW5T73OVqJuPQkyBWLI/yVnClYNPFE6kaVoLYfAJY+pr4A5KAXvo8rTo8bi0wufY
wuNjY7FdXzrPbcN7U8iuG+q8qHlTU3l+lTCQ3cHREiq1h6Np0u2UCRQW5QpNt5m7
soJR49gFCB+xmQ6GuhGA2fQeqp8JmIw6P4QDuI0W85Nqt6bchfbVgTHqB7JoSkmn
G/qxAa/LNInW893ltkB4idKcQyRzhZmPBucR6IfOu4cl/DWQiaYONisrDab7Jnoi
pZTh7pIysclR4HjmI2OcIEiCaZ+neAZ9/koyCKt3vmdeQqVKB2hEP16i4RPUT3y3
RtpUttuKHxyygwwgy5+ww9/XhFIb+09aRrCjxbtbrmKTthsTsflPY0GK4k9AbTLT
RsW1cC78vlhNVRc5XVnDLyrb/QKBwAEre0rYj1e6mIkjWg/Aszth3pBBCYH0rl27
GEkzZda56Ed2BAIK8KePZQDQBLNLRI5UK4+c9YdcUrpnQV4LORUHsro4b58B21ue
B+vOVRC/kCAi+FPDqkskUmZdrndriRdFcuYUZ28kJz6TNOVJBPFZRGpdgjWsE982
15zEzgJvk2OzKgkMKxAjZoFbW6w1LlFhC7GSQxogx39y+JZ2Kox6s4iU/EFqU2dj
daI4vsbjRauOAKc7zIBtJlIwqgHCMJtyhvapFX8mhe9i1pfb1Ld3l+sO02bsfgYT
Cnjy4QHCn+L2+BBm2VCO+AJ76AUW2Fof10VtpAviiCv+AC1vpD0rKxD47/df0vVR
rodgX7I95aVbwQRqOpqnQ/uPHH46clI3/3T5fcWYl3Xg024OniJ4JcSvR8DPbNbz
MfZLa8LKuqpIpi9U2TFqrqejtle9KLEea/jJGCqL0UTc+okjlTShIvtTDJw2Q9J8
eCdI7MUpphww2BtHirAuKh2zlMYUDeb/o/keagD24np9dS42jKv8oERbAW+aV5WG
ahu2Be4xHGjmR0fM0RF+fO84GYKIYtrH12I/UKZTR0u+mY5lXmGqLkbL2/1dxv4G
Y8BDspS4AR0WmkxMm/8beH0+0Rgr92paLj06sc0y3Z37Tvbkw9X7kMWJb2LWfRyX
eHkvuwGdaEFYZJt6IB/0mPky//ZH/vM8xpLL2ku8v7Ya4Qf097mWMZY+6vkWiG+k
AeXo6I0mu7FvWI63v64+dNDEMcVSZ8n1E0rdL7waMAyByJNHRj/oPE5IrCaFM2bK
+mBp+vEexhCZw3c1r6YYhdHdXVZaVh8gIANVnSAJOGlkVOH8welm1GKUXodkoqYF
Ji5QgiMw26sJxjuzx0fk3HPNDLYO9mAKOlyfYt6Hfg+84gHLmifBWR+wUql0Nsnx
kicq3tLBlL9NOp7CIKSXiOnYt/T17fZT4xR6wnIvkQBXiF7wwKHbYE/Tzy/vNC12
IyQb2tVS3xjuPoCIOjL8W0QUowyR+/8ehhqRnhL4z1/HxTUckwB4oOUXdFIA+3vZ
Tcgrp0VoZZt7yi3ah9qjZ9pG55tpgPkN7BjxYz6xC6ZwP8nJds1Xji5tGZIcDhNy
WKCp6zSzUpxSYSvhvLe/ykIA/RqKdiJwU8v1r3Uz97HvlDpW/be8WcQXZGnR1I9I
/1oR48kvaOIDcAs7rfaUfzs6wbol4cqI9/68zxUYDGwR/qdwevp8b7/6kEs/TzFf
b/cYzoLn2ZIEvsrIDUW+6mcy81o5vqP6ZXpXsP8sLJMAY//JE1zIod44eJ2JhL7k
l8KtKoDFmMwDMPH9MgLk7sK7R/BfVAElPke3rIt9ONLOl5eIt8r0pdQCbu8Ow/xq
ADJSpEo9I/Wp5CZIAV0CprJUdB8nhSMZ4NN9Yxouu3pi1C6UNRPj1H4C5VbJhfsh
rSVaW6XccV0QiJUKxu10YEiAP8HkfkkltEHkvRpM4YGsFK4Aphx9J95Ge6Hw3G63
xx27Dme/kFdYbwIp6IGemPQGHy7edJEKyFoIKYNKvDeVFG4P3ZShW5GriY+gw7yX
j0KVduNE069mICLvoTyG98rAQEArwqIw93JrPj5yD6PFHRk9phjPWJ6IsF3HfVKx
i2LmZfUYU20pJYOLZPkOwJjyBpcNbYom77BBW1WvadD9IW4xh27fhQU2YB0CdzRO
DJa9FUmvJAum66OSisqgozHTAkxt15W6fzK9kwAsIgyVKQxu20n8bTrmiy0QHhiG
rJ+i2mIJmt5siNxxMkgf1RfbUDKZjcDMQmy2FXRHGgPOKbTTg3/60QI3Etrtj7zb
TTUvrWLi6zJSlT7xviBOGf0h5I1Kk40ZZRCaamNnIcUlP4Q3L6bJPMA3GDFr3t1X
yBhK9sU/4hz5T1MzENUjufCDDgtgdUaJomF3mjdQPOyBKyT4sjH/ApzKzImTNR+V
hFUewRdQRDVKodrwbwG3eCoQZI5OYtIQKupVtQNHuGPmR4n28YZaYgQIqf/r9r1y
ls2Vp+0XsMnxSfPDRZA16qeQTeHy1Seetw/tE2wgqBs6Ka+ArKFCEHGhelEfm1ql
4WHPLoffMBQtQiJEQV+YW7ElWE5Q1yL645nEHichsAl0y4n4ZfqG+Jfz50Ke+YmW
l3NjtutbBz3k5wm8vk5wbIKL9/t/yuoaV0lm44x8KF/9/MomIxkJ+qDeCOWsHhnp
eAWqHYDouWumF1ZX6xuY53vM6c3gKpqChe5viM/03TFZCX0Z07BK5xb0oYx8yZFH
/6C3a5YnI9HsvWkdF6ysVI393kxbhfewZ0L6/J9iQwQMqseNAv1FOpkCsnMENaxP
bPbnuwlKYFz0fiSosHmM68/Td1WYRN0pWx7cZqSGgzEdw+zXRfoXK6cLY4hrQ1LI
VcI6SKtRb5Q2babVphsYxB3AQZlusDGvWvU4Njq6jHASSKspmOjkYFrYW8dPInBD
AbKia0DO3HSasupMRciqufjidUY30Koc6DteMoqlQCXBaihSKbzFBiOuylK62nJn
5HD6BJZT5vT1G4CCtwdjGG9gWrbqGuuH9U7Qz47rQJN7PUzZhJPtTVyG7xSXOEMw
L0kDjxmqSylRtJ/AZsDVqHWXPmxDaEJ/SCVVzi5Gw1fpx3X9A9TJ1qWR6aW/w5Tj
CR0nnJgv9oE3yXcucebJQZ1FqqU/Vou6EvMT7LfKaMNZPfZoI2gEmaKWF0mJdEVz
D6bH6Ixt9eH58YA3LEssNkFJZwyMjlRp7WSpNVfsdmR+6vKdHK4lmZOIInFPWiOK
X98O3qUrWcEcRbPKF9/w2gtJ10cX/sJaPO30/bKSmfyMojlf4GiJGhP/bNRh/U0e
q67AjZE3EVGIUuTeG+WcavjTVG3kFEIo/ECEaW9MGatxfXDBfihiaze8aeXg5keJ
q1UKdPs5yZVTDEPpopkzxl1phvKcJNjnz8aeudrtIi0t4+TMr74TZiLR6ABCdQyU
wcn7qYOoQcm6MTmpftXsxC1QwsAyc5DYcQr3WqJSdWkgvCojiM4RKmTk5b8sDUng
76TlHV3/ZR1KLLKgLF1k02WTfV+EB08VKUAOUcxaFdgCwDQWJa1F8D2SP9kPDTVo
JOE0XBgGxaVGCs3z6jzj2lAcKz8LuNH/KuwBN3DXHOwZSVSMzk+qfjG2wSqWylkl
LOrRN+kgetZHaJA0PPt0tztRKwoLYJoTtRJ8yOLaEU5GUCTB5qog23oI9vb6L2H0
K1ameLZPUBxMV4am/lyWHx4KxAGVSx+WeqfZbwy5VfoNXZlSFeiGlMlVwQpjAAXL
jNCULLg40HDa3dRIwSTATdN7rGOG5ExqwQV+EMQUbDG93YLYfwRTOAww4xY3UzAj
Kam1ESFiEYZTDurmb6ECjv+rLLePuRVaAQrklW3NgQEllhlIFaR85DHXdZlxpRrC
aIJqRmTd+onZpAw7O2cK13hmxNGBT9nvq1+5xxuWeX2vHa21Z8bKbgVVCFwfVXE5
8oyQ5r3xHWs4n7pb+3vfl1oQonYPb4t81wqfPZwCkbLevQSluWP5FR52eevbKdos
2HwFwuPx6+kaqE6OIXLInemg2zTxmO+5eO8msRzu4qOzYa6bQA5hnz9Hq72znPTw
djERKk/6UKqupIInaiPhGdu8BoKLGaF0hX1wfksZTJJv42tDBfF/kdZtBngZfvha
LgnMsVDmVKDg4ACeCSF1bb66VmTkp4b2j8Dz9YokPjxunIim4/IU9RzmKJpQ4xKG
WexTUmQZwjEsApi1oxcaN9WIvqNgJt3MwrmZTw2cuhN6v4yR9tUpZjeyWphitSd5
5irOkVR3j+gDYjNsRLFalZuMQg8KZt+LoiqB82mQXNBd+9yXJYqb1r0IjgmvSv0K
zV/B3R5YFCJnyVIYVqiwU1RKjBTavgbVwmu6tuuvwMO+xCF5fXFpwOZDK9V1JBPN
IXtoidjl7iwmeEFPzCFrUvF6jEi4tLve9Ga4xtVNzLRaY3F2q6GjIgrNLNf+jSsj
bNzCKr5UnUPNPkyT2sqT7jQ5JHus8dMjq9tvCNCz6Ev/5p04961Inc1FdWw91UST
k5LPP1KCwQrptjTKUrNw9wTJ9Lv7g4e7zjqPfHPxPhE1bJ/BtXumk3l+I1P6cuFK
ze/0sDqMJhk4blG81Ol7g0V6j8HeY8Lwkmk0yeIcZx7Sq2wXzgQBxrZLvbwKGryh
+HbuqxbZQTGPrMMcMpvFtxKnhQ1VrZRtipxjKSCI9kI/31Itz4Gr7VDVb5hvaKZJ
rRtm8WKO/Fj+mAtvWoOxyUFJl7QugXA7Jg8yjsL+ZXJYVVGPyJtuxmwRDLmTJ6rE
5ZPLIxmNF/Wf9iMvP1YdeFd8xL23TK65qxGRece9MwpsF8g2kAJRGaoYHmAamWog
P8G17/1k5gcRcB88bvTop04oPsMgPbGxcRtVgOX16D8+7IRcLWPJYgXkgsdtMojY
w6cdrTjleORZ2dIQUNmgyHgqCemFv4rQw+3rOpTgOkF9VE0f1D+9D6ummy9+hFgw
3HCZ0je4TlxrN4jZkQNCctwgnB/JbGTEjDmLjjPiWjV6l1nZ4GVnJp9W4tNIjVWs
YdP0CXWIUJY4dpsIGA0UPmz46ZKTJixrd+PFjVyJ+TmckciOnhNZjKzbXfWegObt
wN7XbZjqp2OyCGAGf0byZOnijV4HSkbQw/piupw8GhpNYFlq7E1vUbA36Wq2MCOe
zzIPVg6cyMwES22QOw3q4oPLXvi20BXpfCWYpUxmqEYnZVZpNMA59LLhWmFU4fTn
7OElT3fhCUsfuJYk4EyAgKOxvVkj7YSgXgHobVi+c8OXt76/heUqQn8JczmcyATw
gnVhP4jyxbHpEAb4Yy8dURpo1xQn6MUaOkUBNZHFxYcHfG1HFhVTKnzlKLDKYLTU
JJHq8R0nv51r5udO87JsEU8FS3IOOBYiNF8FDK8aT7jB83IESsjQbN4fKtp6b5Ce
YgEoOJBU3U266XQEXxAfFxj37D3N7EOIjRsaycbHXCnvAAv1orpzkwaHs3GyTMpN
vxXyOYxXVHocBIUyTlXpiNvEVWzeZ4ue+kIk1xctv1GWXsEPWgn6uRuGhVWx8qt3
PAX+wenpuIxnUrzACfDPTtslw8XSO97h13lCk9yxr32SLhY3CBgCkn1AYWMUCMQC
gi1mGwOitImNNUFa4Eu1HrRoUf7RVPaVABQbt+ITN+OaYSwM8zlkR62adr+3ECSi
6s98iYuLMEZUJoDhqvTKBtBqIhn95Kzzhkd1iLWUxlMLWVs6UIBZ3Z01huhqgasj
LFXUfgYRvATR23823g3dIhUqalj0qyRAUZ4yx7QmseIRs9LJwyE4dvvreSIg20Ss
W44867aW6oPBkMpO5PywaaNKJsJY8y94x2/dEaNU4Fzb48Aanq9DQlQ18dphz8Sz
J1mFSHoMNqcJsjXqruWsn6eLwIR1ZvqQaokkT97NCPFt8Qb/KLsXp7kXaORE/3Yl
D+wQ+QdqrYOMLK/XxyeqBZ2RYEx/P48vSZubOD4R+uO0q+3/4Mg2gbyut+Lixnt2
hiHegz8/E6br8yzhglzgkMNyQGvFuYcfu9ssJCX42D4La7BSEIZMUEsxd1+s7jDW
eXUhJd443Ayt8ttgaKi2rLFub2nKPLb/my5/XSSMf+GJNDbHDtK/iD8yoRPIJ60r
dD1K1GkklwXwnxK/eEcnv9zmcwZjXOxGzXrNo/NNZ+ngHwmfXAbJrdc04J5hhnSi
F9WWjX3V4myklFvNEnxCK+8x3148YkIZSlUrQ0OJcwPlChpE4sVKGwZLoVJWFknz
u2L/bEyR6YBcM/2/aCZ6VZgzY9O8cdd6eJJskvRdJ/9P0Vgo871K7juilRvtBOnW
kx91LjXoklcVB7RUo1LXVwpYok0rYCnH1vC5v9BYWy+3QiwvE+UuGR3WC6o4yyX2
Aa8D8oKnb//pD55hI9phpciuPK3yQnX5mknOrRtm1fXlQgEb8xsepvdRbyXqpEQV
laIVV9IEbZJhkuGgb2gkLEw7mWpB1ugwmS1SUJxxzJGeCwIzYbRNy05dsVQua45Z
PnkuJJV26EdarSoEEl5ZxzzojaKIhALGvVy+jpnOTheQYDw4mW0+TjzOuDLiHGOg
tOyg2/ehSIP2aCr0ObfB0X1GgKS9A7o4kW2H+8QKVR31jknXlmBwnkegd4ggeyRr
9MC5qWEWKz44AzuXwncsiQXtAdP4nAccxfrXQDBlNtHXxkbOJ93xBsS7YPX9tp4a
s1dge/Uz8vO+nss/sGkFVzJjVKslXMwNXTzpdVvubn8pVCQaSpo7BbbI1eqdEYcz
4lcNFaA+X/63L+fqt/W0ZTy9LZphozL6DqY47UOwDbMq0EeX2C/7dRym+lfHl83H
gfHARf0bgamMknH42/2rocVGx/V3Fs8GZPQnLURs/tAZ7WUyiSpqF3dRrjmsNBc4
o/+xOm5R+ZNZNPRqQ93eBcJM12nh7z2XG83kI6DzOdf7oCpCTNQiLajnYJLfFLz4
HMVDmAeaEfaVbfCsYaEGriPCh69KFows7TCd3NHrbPsHQbx58ub9zvaRCKhYEdBI
nA+gb5nlFuhx5dS9ZSJCn+iYxLLDcLvTWc+ByykxLyiS+TirP/hYKxCWtlkmfhUf
zCTykFcOB/+SaVhDB7igj1A3EJ5TUTlw1jUn/sbcs73u2n+5wGEVPEDtdCTM6QU8
CD1bTEn0A1N7makjul3HyU6xCwl/5g9zaeEw3pIeARFn8FsgicRr3/e3kIzhuzU1
rE+tmwOP25UAbXjhTuWw185S4gBAdPzNFq9J7uBcre0ABc9bwQynTnsGxEItZZjK
WQ4qSuIO7HLPaXGVxRhdWsAQNzmT56RRD1q29QyF8Q6259TAfTSPTwDDu1Ux6mPz
QErJLYQFI9M2y26jyzSNWlaVNGGYALuXtMVbzvJIocFr/aXJdHWOuyoqQXnbs7Gf
MG151OJBayFjG9vwatB14ArVzsFc/ZjTxfXV8v5kd1G1cL5FRZQRzVxiEXz8D1KR
xe8YcsK2O5FoUznKXJEpCDmLqzO/Vj/N4EjWc+XyHZSqITgteh2e2xFac1OvaHgS
uKuRemdSsx7YhBg/tr+4N321Q8GYm7aZ3aa5sY7qUKxrc28M5ckcKIJDMkMys9z7
P6PvuNXAAF8n/eHjqWEP6T0KX8lSk8YWLbaoAxmaqDIkoEGD5AUvB7ue/AO9ZbqB
fkrdoJl3agvp7UXz83pxOoXHOfxLHNDi2FQRgFYO77+NR+0UlLlez1NFXWH5qMev
jjiRQ6yCv4FZ8TP3W16wYtSUtkmttfpIMsBd2aSFM7/6sdwrxMKWkJEKn1Gk2Cei
jgd/KBSkOpbX2wYaTnzE91yG6sY6YTLVP7JAW+Dq/G/GuV8e/3obYhKnWrbuu+NO
MD69DHLobWXwMgcQGFsOKL03hjMIMOA9764SnPZDzMgT0tIoSBvHm/nKi+8voWD0
/NAls8grLpD5F1Vb07qFE/ZTj1zu/8DRBpCivCxXZugoaRne2GfhLLIikM1uump7
9N/tU07FxMJfr1ZpkRTp2TDxsXty7OX2/iAxQpLz07BVsWVqKIa08rJZvmP0m9d4
er7KQIh3YZI6cma6xH80j9AaQDM0k4J3CnqjIU8Fyyy1eVtDai17jtuVi+ZQ8pMe
+SPNJEbu8vfK8SeGW5Tlu2zm7CiCEH7FX8/ZV/+MokVDvdYIVbing0xfCFkPvkLp
Sw3LPy/TFiRTkHRsf56059hg0gIJdAqyPxSVSvRuwL2jp9uNiaJPgMM5TXGU8pmr
ZtRq33GjIeW5O4qooiaaLGH6YCVi2aimaWba2vDQogUyNp9XlDGbAB874SQKb1Mr
DNTbNCXzwMPqkFnC4uwDdmb5oYHR46w6T5OdMichT05AA0F5SNJJfWni4YbKOPIr
JtCHuyllV9IgIeBRcZdaM+wT58xErdH9t+5zyqPpeAfIuPT60ExWSp1Vzl7FhLuw
27fmH3+ZVkyc31CZByuOh4ErU3vPhLeSVqrdEisDzgr3vOQVlIFq6zPAY7Zls0Eb
3lmsm2vnyVf7GkSVlYJBFq+99Q2u4GxbgWnu2NjY/MArs2+G4YKU/RLKR6opemA7
j7zdWXYyK0VaKo8IBbnANBBOT79XY56xkncd+FTUXSnDXDEakmcfgbjKqaoXQ4Fd
UkLbH7RUn2TuAlF/VJt6/VRJdaMgrEIeBRRcIJ1uowah61DP/UAFxH5db85AI/G7
ljLms7fP1+SKD87cioA9TilTt2tS0JFJ/S+OD+eI9k7iKU6Ip9O8cZ4nACPzPoqI
CdtkyKym2CoZZFnU7cBRa4IwffMuHHU4yBu4NrrOieYaur71EQpspJnacKslghN8
qEztrqVffh25PDp/6EC48kdPGP+bwSxahVXG2jfWHnlMpVG8R6tg6QrcZLCTORUu
9Cy6tJQnj3V3z24ZbVo6RL/Z5iHRedeoeuWE3WqJinmJszTBcGLEc3RkF/YEyq8j
uxofF40VvpqiFyAByN80AR/yYgrh7UK/579D3kqiijUIVLwpYuXO/JSrs0gGgPWH
k3Zp9x6Fdl7p3rZ8yss+k5idKTQlyuCfWizT5X2f3J5MgsNXufND83JlFHYQBFfF
x94VS/wRIwOMtNKGOHj4Y6PT2JQZprKpEY8iWAEhboTW4GyRhmQQECNGfrM9P3e1
cx+kJxJJAlo02/6qeqPmE9JFQJmO6cnhhGAq8EEGxRCvE/JgDLh1rZFSQRy2yn2p
sLVHzOgO9vmnrcAlkbOOmEMUdzHGlpdrk3sC3vrXAHtpxUZNXQQ1zOR9p/AV/5WM
plvHUzxC/R8YwjLh5gWPq5tVNqCVh9OiPSNTX7XJJwEFPkwFmYgm0zmQHtXDnbrk
+yXI0U+f9l7n7CJ0fIkqGayDAdigxPsPGRAtu+V1QeOv1hDfqq546kQhxGn00/qi
Bl2J+UL/6oDIfQ5+KwDcClwoTJjKc3CwxDDy7tHEjtqaonugxOSifjQOKM9mCWbc
vY9YL+PGd8rJTbzSPQNo+yzEPtPKC4eTNKAcGUX0wM7AOg8TouKIgx1lCHikOQX2
hGwOmFjAfX+m5E2TKszdC27TnvePpWGaqEBQtRzHzMOh+5jTf5zup2P6qg00pt1r
pah3XSnADgNgXcJMnyOPmWrhJpZ789E5OOjaEwPkg7dBLMTkoBZ2sVQ4KqGdDk2m
xmy7HUVwyfNFN2wORC2ikJ0s+28ig2AO7vsAa+ZYCthm363aV8A6lMzOHXfWjjDT
VR2ifj/OaeUUdLa7jNFgsDMbFGdOEa+HMPlAke6hKnJUziXDscDn9jqAvevDu9la
J5hCF22ce3s2/l0LDJeU3eVJ9TgqtKxJFqcupXTMKnQ89/+bNgsc4f39J45ar3Ou
iO2mXdVdlbCkxoLZmqaQk8k0oNR6v62r7Q2/enAGNMkkAjrr0NP/2Je3pICl3XBR
0IRMBFnIqtwvlL51vr48yHHIXiGybNZsNc0TmgFwcuLSvByQmWoyt1ux2YdVVvne
X0Vp0boJL4vg6v8Alf0AuW8Nhnge1V0JZGkNOUTC83Aj3POj/BWMSZEpPCV7tdJK
+0vKfY8nTkHJHJVvcCKsz3j2MaTc9KSQPF3tUw+mxRw76CFV0wymPOa4s75jW5di
7fvqXuOf/Jt04Ri0Ais3205YpmBIGOeSNT5bzKs4tyPtaQ/ZXnDFgMAE2cxKVYIQ
AK/awBN3LChu/M3bEFF9/EFXOnNMSyy7D9x8xHKcHJwq0GZmqGrQo5K4hZTtu0bP
3fgHP4L1lHSJJVXBY+3k/KO/SjYEsXrAY5RBIGDfuhQZxPM6YM0meNwjMjYrLUXM
ZkeYH0P5JTNPnqh7RINTGZO+LMmHrjVpiAjRs7woiw4JPTEOXAFoFeQGTwBevmpl
R7hN5WJebGVLJTPIsg7gSK5NulrmsD8dfkJZild+XfDWLh1TKVCKONmw0QzZzIs9
tvrHJH3zOCR2XhldfHbGkd1/Ehdcmgn/ezvRp8vL8ViyI+GbgX9g8orHBCSYbtWx
r0Jz0I7Tay9FXdGWZULJpwymTRgVSh9IMaOhDLszYQ5HQdXvg6X28bF4/Rc+UfCe
anDr1DNz8g+xGuNPw8ZkKOszARvbmfU9V+E2HONasfgXAh2E1xUBEnlmDzMfG9+A
nCyYJ1F0Ny2eridsovg0ZPyrqGnwI3J3JSFWtY/93D0OT9hpzlVSb+ixdD+WXidi
I8FOJZETkpTnNvTSlsI0skFGVIi+w6NCwMKuEZdXSHJOC46qCA/f6yTf+BOd11/n
Yy3cpwvPYZwJly9/2EesEHrrGVg4Aw6gu+4ROgDWWN1wCN//C9Wij1LgEvJIA2j2
ERqrXNwMfeAVS+aa+zSrO65svLgWa4r2MnTxpxTk303+j1mmpzQqM5ghMubQW2vR
obuD1UMnVzu367DR9X/n7dnQ3n2ud7gJoFyYj9SbAKbgtiXPQQoFvyPI/vjYVMOI
ArOG/yPa1wEp4zu1cNyfRwz9VJbZnFJCCVL3u/s7vHzbqHYmydMh55Wyi38rZNVY
JvRc9rg9pqQ7ylXiErsu8+UDkWXua/9F94uFA/hXjsCAbpmeiPEMHqjAGfHRO+4J
f4+D3ag9WmNlXYSvrD4dInZwHZ95xyd0MU/NvSlNBe1ROm1iRoAqcFanKEVCMd3x
FUk3U93NtCOQMA/N5/V2/n6WAWgtUoD96gIep9+XRr61rcc3DSNBjg0GAZIl967X
gczrxX2pNn0sKWY83DK6I+lpcqfbnnvs1vx+Ho6NHY+goGxh7E9tVM9THQ/xzGJh
jTlJGunHMGLHDSdI5hcATMnYZqxKHac/igReZjreua/+zsvuFsglvQWgrKH8N6bO
3Izdwxf9bkD7B4AZM+Sc8z1uPPs3y41SoPA4AX/0/Z2clvlqjftPKCNLD745UYFA
2IWdA1EKayw1sdEumJFJsXpw9JGAJ/m21ta1Jk/pN8Nun2zepmvZvu2cK6O3i8UN
yR4MT5OdfkD43XwZIyTtaP6f/Gl69CpMgchgWLEt74i1uWNskLvz/bjzbG2Awye2
vBy7Be34kR4Tu/YJlqbUO43VBu0ICFcXY92NIdNqL3GGb4UyWhN2pHRyLGy66FOg
2QOCODu06zqTGaX/r4HMHIcMHNwg3cZXcYDgved0Gt/OcsyMM4gKcJ6B3DI7lf3w
hFfuRwWHaiAmh2y+Ft1PuIFxRxqoxUIhwiSqvRGGi2Uj8oKYZsGuIKjDOqUJl2Ix
Rb9T+xoPGTDDOcM2BSQW07VwZIXwy+YIvDn/qNyE90irTb2E0IkGuJplzKMfvqbH
bxbs5nRNZMp++QV58W3MUhvcsoFOWcn/CQBqb7FJomq8LPoCFlwtOkYc5uCyACQ4
POxfKHuZN+iu54dcId+ZhUJ+fKbSR/fmkPWJvr/bxX+EapYtQ5nb1wpypANDaPEQ
MPPOtNfXQnsKbbqpfG/q8kJwT0laWjqj1KIqYId45vJ7nbJ8o1p98kf71I5jtUWd
jcyZqAlvJ8zmNbSvzit6Y2KEUX/RxY1iEz32BIGq0M+jBPfYmpqriWvjAvohfPXj
UkMLSyKtfzo0uecUaYqmsI1BjLnmoedTEczN/Kc1wJ6KCqZFpRKf8axcoEaAGPcl
ic/CUttYzlndJewUDtDFHKNkDfhACr4euXMfcq9rU4ynFDFe6aSxLCpvU/fV23Yq
qxMZzEUommHrZe3RbvHwwrj9GMSNc0kArz1SF4gvam+4JDGqQoD5sSs6oJjscxPd
DhlsZynWq/MRvZXdUYlbPzgXaHeOzqF5qRMHudOYu5gOiHTyp7L9+ra/m9XFAcdl
K0M0khYND4Zd9mqyjGVSZYESZH3q8J7Tke5+G0e2oWKCFfv5KoorljWaPGvgt5sh
8B3djDvJwIkwb33V7lTsC5R6cUfIP7xhDHpZgKceoSyYD8VGgpge67hCaENV/lf0
3wWnGpp61lQOqnb4EqizfkhxkCPx/2YUgYdAtzLKaLM1/qI6Z5OfC93n7lUkk3O1
z3kCXVC3s1niUT/38z9XOkhs3UjMMzk2rf0ojXfBa0CX3uqdiobBxMN2Vn6uIsw8
WCOKTONRHJKCsHmVTJd1bqRFpyYJCrHMJTsKC5V4rBFiVIogGcFw8+AwpWrXwhkK
Wsa6LXft/hTO9/QYelNhWi0v/N8Dnapx885v77Q0NcggJ+AbtzLHx3mBVVtyMAk5
a4qnYJa5nge7mtT5a9W4Dsn1DZ3f8H459NtE5OmvaddBYlAJXFR+UHZrk9uAhEW5
WNXhymVVop47jeENcj0XD3CHSgFQEQSSAdc/+vLdRyinthOZDbAUs4XDHsYNvgrl
O5vJzSRzBnKekvBuM1uqJMegwqpynNeban21+P8CL6uKFYkyKg9pgr112hBf9O8I
30oeHrDvweHq5RpEpHZgWI9OYaBDnMlrClFi9Adl3Htb1xQLdBwmVjITyVepMSct
ua5nwH7mLQ3iTp1q0DkacM9zZ4zk1QwyUV56Mlv13Vs5LtKyQKXUQiwpXkgFHvIw
9yEKu3VRzSIzP6oiRH6ebuhhA2pQsd/gdoXtpF/paD2lHQYJO4BXVeBc47p//aPr
oY5dckjlx4Uw6uTn4RCkUKvCQk2siAaLsv0BgkvV5V13fTUN03yBcR3opL1xYQLF
CyeMnkwNHg78PJLMs9J1dqjkMc1mLgu6/cYmkNKTHYeeMnRvEXv8dDtIX56zjxev
5iY+g6d9nm+pymvvYEdcmJqo4/7ZB47jPRhLC+xPKaqunz5FgzU7HceWiG1HV4Hw
tSxY9e79aP84rRfaeGtkZeK88d67KFOhi3AM0zJVadG43Fn/WXBNI5kNb/sdQLY8
sWQIfl2WSn4jvhxGPs7XTpBovEtXpZ8nz5bsGMNc27VBFQ0Y0nNmAxjP8OUM56Sy
ov/sf7d0KHnk3esSqS9bpQUxzdIBxATIRcaeRELLa5WPdYJyfn3sH7g6BI4DF6yI
d3uZ2ZwuV7oHU9XhD53Vj/MBAPpbsAatvnFFw/XUEpRBU6kJqybZEHRc0yApXxRk
GQr/QSa1K7Y+G4qtokdZnyTBqe/rEtbZ6X0f6yVPtMZq4WR+m4huuXOb+UhzgyaX
vWcmip7v9qV+3JOsyFcDFFnM5xZ10v6zIk8K1zHSclOZrpxW4jfpHl2lx0GpOAED
a2bxauYwgxmHkCO52Oy8ioNB+AtLfVNdmBeHh7DgbBB+oCnA8DBcn8zdfEuvkwsj
npcFBNy6J0trqi5AitkiB3YO4/A4ex0yAdxIFLonhcBbYw7gax1Mmc3vnw3zKGl3
1Bb86pHWaai9VfBDRBG5+xLYTqK6KC2YhctdJrH7bunKwxncxOz9cGycpG+hf4bx
NZhJWzvtYYGvS0022R9lD6PMC8N3lxfvUFdoO7EOOci9pGgBDbSwUc4YuUEjVjVw
YOY8dTtsAiVPQa43vN28H3z4y+XdcEXA0w1y27Km8fNDhSqIkWgMegxsa/wTR/ZE
STFSGI6qysxhbHLrhmfaGXlfy3eL+94cEBBJ1zPV2UbzrrBwkxv9eUj1RGJkSgI+
I/BRMcMB5hnb3QQ/ef3HIfqPEVjvcNWZrwnlyhfSe/9OZPrXBUSDsWbkiZ1pBx8c
LrjADWR7MEgIpaPa7CdGWE14Aigr2roMx4wNhsMWzdVd4XWtpUio501UOMqT8GWp
wxHl+8yOsV/pEMhUi67+atOvpG1bY8P9nwMtKeGeIq68Hd97B1SH3cDqmlXXBrn1
dLPLyrHEyISBkyMq+XTLAck4YynKZsQz9GEySbGBVD/qgd8UXj4oRd2B8IU5J39f
knILAFPqNnPfuq/qv7R54cdUJuvhVAIjjcUnyYkq6mQsuc6NIl50ldewz7Y9y4va
2HdEWLAizACUDc0tHC80hsfMi9soKphDPksxyV7qiJkX8y3SECyfCK0gXTH8BE0E
0hLtzlY2iAvQQqdu7T193iWezFla5he9V+niiCN1eCcvI8c6F27XPnu9ZbmMM/gD
rLNM9M4OLsPqMEjdigcM+oOLAXfmLV5o5Wlhqqqg9Rd+cs4OAi/DhS1bWMjCF1rK
K+7oF5qEhtqErIEg0xdpVFzaz3JGMGKjaBNvkzEfMtL7EEqx5GV5wUJW6HFV6uVL
+Lu37s0kWcE5VXTLPfwxpitG8dpcEI8krYDWGS0pNf3kWqEkk3diUzAXB8XYIsbu
0iVYsLG9nDWvnT8DOYgGI4Wq33ElGdt3EOQ3EAQmQtwPbXFWbjefZA56C11nBFe5
lxfzQywbZEVImXPe63oBNTQosEQYruXqSEA8UIEjQN5kq56pMFDlM43meRzPCE2D
NNHNouUcwUgniwI1pxxdlqctniImiAmWvvzTtUuznbNPHgnzNJrbJnzQkSgMuHFD
BN8vMyCL5l8FLl13IJ0KRejtUvWdsqR8RH7eSe9CUYU7qjRe1El/czSqbTGiLVPh
IAZEGobcyY8bdg6HQRdf2NbQQMRi6JyHjx+xgipiPNFwmV3TWiP8O5ndv9RfnEmF
BFzep7iXyw54tAHDMJaY2RWvrWhatIk4p0XS2F2lXX3/vufgU7aAUPkm36Bn8LU2
sazFagovVyo/uRfinhtpFigbS80id0gdwQKawEob2RflCYaka1N02Lhm+j2BZRLI
DLC5TvECbh5OmTNJUwL/vleCQJJfDg5YH4YZJ1zNk+1VSO2946cwAOF1xazpjhUI
sgmhNDzcKx5kAkRwGrYwDdwzQYnO9ZFQiF05bsxkH9V8mp/KtYdkdG2NzOAiYhJu
t1Y7qcI3d3q+LXkq0Ia256tKvgy/B22f5Ajgc13bTL8E5ZtHVaRf/19k8pu7otHy
XzGsjEQQ8Gh2B0dnLQjlUa5atyXDVPPszmIfrHNdZjiPWNZRdTgpBbG3BRRG865L
MWVzpq3hT0UckAJVau9SZEWOPcZ+gtMQ88uTsDeCAL3HvY78AvV/oouU9QDrVtCh
9PQ/6HeD+64lowxHLv/gp5FfUvSbobqrYivjGmVVnR2RUtFVpImoBg7nIbF+/M8D
hnmSknrpiuqJzfg53OOcK8GuEiM+wNlB2BWjnWN7VQ9DG7zMa7eI1ujxAAk/U2Mm
SYMNvJzanifnRur8R9sL2RNeOHEZsdoRPxy8QCrIKlo3lZ7d+DJuaiI8D5xVBFHa
mF2gxzh5IFJOrC+zqnPaOlL3aSgB0NL1p2JIJAKHlm7a/WI6Dty8zBZ98mPQGPfv
eKIoy4C3k7WXNx44oSFQVPAynkBIYT6t3AdDV+jdPm7295WXwyWmbiGMC8HZQttt
SHLYEhT7bdm26+sc+dd3LcacbiDjwxdEPK7yNNg6e2PlI1cLy4gQn67AVElQQiXm
Jl/qED+czxyZ82I7iVnTfSGKXxD+9wRUv1ThOk9jlIE2qkTbNSqRRL+8Kji7rumD
ihFn4Tf3OU2ZGjjRUQonsqisk9QVTs3o3Ez+V/UvkL94iylymNsCMgQH6gCvfKlV
30IAZl7ULVilABSXNp/qNvRUavJyMV5mFI3bLm1mEoOzwcH/LWdT0Q2BQFmVmfAG
7l4lGwEqaxuGFudgyUJif3h4+ZLUoiT4uyrqs/agPa9dnMvkNho7lGnYDAqbKEP5
E9lT6D0FvUYK4b540Fo+GIXmga6G2yuKx/X/ItIU3abcybxkdsOdxfSvhRBka0f4
atIH4gkCwZNOT1N9N577aOy+WDrTb65/yepWITDIJWepydxjYeUEgN3Ob5n/W7Ei
t6Qn7x5Ux067WlwYZzEwRd4a2ZaoGN7kj2o2oSQdbAjozPI8dPhHkkccYog+Mcgh
3F7Do6hDOwZo+nYi6vNUXJAC9HMxtIcV7XM8rLI4FkERJELBWaxqmG2+1Cj0V4ym
f9mLFhEX3Fta8D9e1tuy3NxSiHGVkEqJV3GSLRvS8BkJ2VW79uPIP/AJQwRPpO0y
d+6pFQZqcKiL4lCbZzt3iLr9oTYUgWTWgTda1YcwWUL3ra6OZHh5Cf2VzbktFeZp
kzdUvlGlc1NFR7ohIX2jIYqk8Hjbkjjx9Jx/tQLzrYoy5t34TOSrEae3WLstdUBX
fhf8widHw7NzxqkS82FsGIXWh6pIeCmuMIGSCZgLh6DtPIjyDq8SXAEgnwo6YknP
cfND6kWMYmQg5ywHLjDCmqDFiii1tiOaD88FcfqfmL6W84+c/ih1GDbpP4xGc+rS
jKm9aZgY9/lyOLIbXjxpWYpBUs3QM0rJhjRwMSNGyZPBu5EYcfi0DjRGgMz4va5m
OmVBIGHhqlsUU37QqXksSFd8DqWZGPTbrQoIaiGsslJdHNyFcN9dfs7S7RgsGyzc
oZxKeyRPIP6xOskQaUehS1rvSQ2nSeH48EDl1fSopAu/25mMkt0y6VlHwfD8k2TE
NHBzTf8ULTG1ujIN+I/cU6oXTVK91CXdfnWEXC6FOzkXXeFX+tW0jgytMHbcZI1u
eiSgqqMgUf4vze34Py7atEgHhGP77Qg80k25DpYm/U8spVB1fo1pwgvbyoqOoLfN
BK2OD0opYvGbrKTH1Bg7DsQUe/po4tyo+HfssmKvsWycqLmK2gxC36mhHcJKyTcM
w1/4uDOBk+bbNAtoMh/jI/C0Zjl4NFnGyGfW/WPeUVlvKP6phyDVKpC2KddTWbCi
1tGh853cWPZrXMZV7gkCLHRbUfZmveqx8vVfaty4N81QpIiN2qvogzMDRGdkKxLA
hd+vkyhQPMnaJiC7NACZrPLoS6Zq/ykszh88rxeu2iBRgYJMm1+6gBBqPCaOC1hM
oxVj7MVrsjMtWdk7En+0YzjHzw2rKb+WjHgULJIHxR5TAbH9RDAIvCWfVQK/4hrJ
Hzx4MntLJacZVIGeheoVRwb+j//vNMEXIdw612gCk6zic9iXbaeqTXFEQMiZd0rB
p4KbrIQgO5tmXkR53Ro6vEpdrOEyr2j7WgSlubt+CMbZODsq3FXeyp6fcitDkGYL
llBKSBrhVAsI0n9TZX4wZc8ox4YSfUWOrSMaxpllwtt4SHkmwEiH17MimttKsaFP
mmE3zTv+mtFJ69vAy4lY9OzhTYR1fZTvRc7FzQ1bl6gSh1TRD0jfGUx4OBti0YBR
d+AH7KZTss0OeBbe/y8WDO0VotNmXAUZz8BB4ItcGJb6iyZ1+4nueupeInUyzmq2
RHdX/1agSkt1xAhLjoVXqlVNgnelc0FL3aW5j53XX8MzoSIoqW8iS2tNQh4DRdVI
n4wuk+tkcMi4+odx051dVNgAFgIaAr5YP+DcYs9/JE0TY4JJs/D7jcM/D8a0BqMQ
MqgJoAHYkHMmbsYMN1SZRC5z/R8Bss6VTKPCLhrmWesN0JlOMW237QejD5L72EuR
kuSQXrH2ze+N9ZzlZQwxgaIRLD31Yyheeq9l/IRxx0zdZ8EojJWAf9/BbvpRaGhQ
VN8eVdgg45qpryJwACivGE2sIfjUsrJFXMjZSLDnNjcBtCIz25GCiZ5X3++22vJR
EZGTjvzTw2WaHP1xMmB1V2TzHAVCBgD3YMPyRZlZF93AuWvDzlZHd+rHo9Dkx9Or
MqwdX+tfe4nrp+HxTbMdR/+qW+nTofXNeSeogASiWA6GCYLSDTyzmmI28c0HKomU
D9mM9Dx2GqfCKGmTgd2Kz0bfcjG9lFYsQ9yGhgNnv2NP15v/BaJ8ebIA7+5gRBc6
ub/9JMNMNIYzmDijufBTghllT31w1/BGwYE5AjLc2OqwkP/6p22ZQnpo536WsC8n
MDuS42vFF0MFna+SFak/AjPvUMc8PD5j+F4vqGDzH49RlNKOw6oM+IariUFmmG+c
oy9H3ZlWWi4zZTakhyCMcdHL58d7n8dERM2oUWl4nJJwf+Z7iBmjuVWOrX47Ab1b
1slHVmwvcsXNrYM+ufIbzJxRrEEL7O+AVx8m6NvIdyI3OodBg60v2Ld2dqiUcuML
BhcJu0SEF4QbadGXhJkcCD/f5AQ9PlkW1IrcwWhp9PrwPPv+N3FoIQyfqWphSHl/
abdt8cljUUTw6GBj4oz8Ij/tO/H+wqk6fSllX5oX5eI/6i96xe3fDCLLbvTexIfq
NDlYYGsk+pFJ70oP1NjGHYat57XCR2xpwAWtdW28oyKvQHplWNHn07PJS7cwNFEO
ZSZIOM843I21ki0MpV9EL/TpxMNuhyfC3zZmdRfty4zEE+KFBRxGnODvq2EXC22T
/KXPPYzodEyTPTv6aTEG14tfrcjPdIKedyHDGCakVFbSmFg9PJLJIOYNcO1AsJ6w
nCoFOYTlENA8m4+IqOWTPahsuxHQaJHZlb/8Z9bEi26ynzd3C8Sv4q7M0SppJ6OP
iYrwghzFxLEmGvMCTOVGW6yCy0dICWrLAZhXGYb80VdZo0HT0Q+d0/2/lpsuwB2t
jN7q2wQMC0dBY4/CnC3EW/7Sej8RASe1T8BTtHcKQYoW0MVHWfCzVxP42yPRqDfY
LsI94jYQ54LBXogfik0ozJz586Tw0zVmq51y4G+vUVbjBFuvKCnhskT/jyvc8kyJ
TouP1XIrhgCSxD4FIGsYO9DJJ7vxcimLrpSWTqbjOb/ttdi8LxP9L5AVYOexqA3I
TFnXe9+IAd0/HxdROvPe7IGjBn4JR6dijHyWdF5Lbc9HQcOORXsIv1onYsoX2cMN
xGwrGAj9X0T3Hr3gCQLYfts/LVQl664pJKHgU4gEIorBN8iojnJ6fYlD6Kmek81c
UH61KQW5ppVG5mH3OgdwC9/qDAUnQoxInBBdQ8CSTjTkNAvVwshh+M+/xwVCVs3U
RgcyhcuiEJOD4asMk/aRt41RgJ5jWBY0ht6WTPTLgjLKkn4tVwxfgKgrKLV44jCE
bOVfPaZObNTXiNgYtzo9uklXwIcOZ870CklIR5v5OfiDR8VM1rdXSUgP9PH67dh1
hySvsufM+z244UhQQNSPQEik3OKiKDCammbEuFafiJEa287nBzb3HwLS9YiHC39p
BiADgFtvOCCLiaYETfpLZ3rBb6Yqeyx9eYY/EXb3t5WIp+x+cx94dMJShK01RJ4y
7siLbwcwm6Gbhfj3kTezLQ0zOne9vCCarmVpW+musdrbHsJl807+jrWcL59FlRg7
TPlpZj5NP7/l0mjai9FS2puNDrSc4pGI6NeHsBaG9Z7ZDq0qdZel5kr4lEXD1bPj
tPZRne9aUyYEeL0iq8Jor/aoK5l1J+p9TVczy7OvcE35QVtUFLR01uYdPDk5CVVJ
UKwLk3Av+wULgO6C4XOjKL29C4mRvSTD/6GzFm4HXyKStJclpmCVUpiCdNFYHR2D
iJ+Ka0YLnYL8FyeE5IpvRqKgTHVSA2M8s4dCzt/uCno0Zj4I22tgeF+X5GZavHRQ
eDzKN/pcIMFP4dgUrHhSWvM00wWf33mBxzM70osG4aHyzFXkBB6BC548CVcXkZkf
AMyHCGMNad2n4zBOJLLKWfgRDYdVU5y8tMOcdJbbL4RSwwsRx8cbyrAZ80Mc8BwT
Qp7LLa2ABC0hss6GnRDLCtAxxPchWMzhprLDO2FNfXMqt7DPmP4rZ8sc0/Yp1bVk
oJ8CJ4ELvAWxm/vt8aSc/amolF7brljPE2/bje1tQcCHizQyfgT5BysE0DZzEwez
isF79z1GIhYL3+AuTwn01VRnIdITKv4PyBqIpF4EtoYWLmDWK79HQyqm2EwAajdR
4htoy25iohAv/zb69m4JLUMzBpYSReSc1hq0dokB0h9F25nVT+LdtPbv1XneLY9Q
kZlZ61JDPNPFYvsYJi18vGKcvnwqmo8VZNiXjWCDAelouEcyjRjoJ3D0SUGVJy9X
Hy9dOULCKQFqR0o4BMSl7YCJgk6KVtxLpBvGG9YHiIT+mK9AeFntztb43+iGNVRS
gubmGUXkwQpi24kO4xC+0MLd8IcRbOIeqjIXhVgLFNE5VI49cheHtVYVUK4gACYF
QYnizjlrxk8fcP3MsKbHIDZ/wPJLZWZZuQDXGRulQvYy/EU84TfljK5daU8+FmVM
ZMqDB91IXt7YVsjTHqz5l2+OPTfqf7AGI+9a5ct21a/Q6bUo1t1D6Yfh21dq2s3c
7gQ6yPwAEaYxEl+BJnLgMVzgaGRI0XsKTTaDVITRdO7cMZD/fSTmilhCjh0igrUN
cNwqBrrPhr2ku3yq5tzS4uMW1woCbNRSWDYC4oLorC3yonwVbuEJ4WCaccGPe6/f
7mha9qBipyTBwmLlOpbZawu6Vb00LqX6Uq0Z/+31OJs9gqhP3X6ft41TQrM2haTJ
+ZiBlhA5JF8IlJvjKh1xqdVWl9T8yUak5tDWkm7XhhT0djecCGAJZWGy4KvzY/Qf
tAEXOK20KMxPmqbNJFzX5rLF+JVEmcOztESWqVxJOPw74E6b7KTCDX3ydBZ+w9qz
yXJ7S0riDCUoWEBI8niTRRnH6Q4FDm/522Qc9whbxokBH+CW5ioXg8qynELfNOls
4437DERT6DMaBRkUQHq3xvywQWXkXTvy2/Jg1hng3RquBRPBgteGaWu1vbvEPHES
+kIqbgTRk7VjxQfMSet5u8g9H3WgN7C/4EWfHjRrHpfZluNCneAvH8BIIT6EdckA
dMSXjX1kOcGFGAZSVvLc+ldUa70FeivE3Z8PQuXMvTEQVHuCJubAqcQ4QcN7OGIn
UvgIZu7Pd0rEeR5oU6RUCkNqtGWXCQVwTrtOXh/cHSJmjEb8I4MYBbyRh4GpwuU7
2QJa79ZF3C6uxrMPBuGyIYUJl22XAtjdJKEHr6V7RDUINvIk8/RH+c0YyH0Odofh
LyACWSdvu3Sae4lh8H4Ye4qEVdE0MYczj9VofjV5U61NIr2SaK4aw+r0QmvT9frN
QpkJhJ6nJBv47t3EEHfQLQaCTJvVBXya+C5+X00PdOEcPwaw0RyU+ECK4fiY2hKc
EkvaqrIZptT0tNZW63Mkf5DdFEElxENnxFJSpuXaf1I9FicRMijCG78Gg1mewCIg
JYOgl1ea2FjUmX04x45BNi4mkQG6+vKfBp4f2/+BmETWSgXX0yN3yWw4DFfls9CR
FCOScfqwmDBDG1YptKo/HPmAZELm+nNrAGJt87fXdKVLO6ynecG4hu8D9iApXBmH
4z3bz2aR2EknjlWGnK/jNC+0rc3kJ+B6LjEbsanQffFalM9g8D7LnKpTCthCi9tp
yaAoYj2uett6L8kT7e7U7T9QMwlZC+Y+hGNjYxtRV+kRwQJVm67rDpYty1RVrols
XJj633BsPEsOUtKP3Uue2PGrhuIcHzG0fc9Mq9ztHx9i8ULx0Gz/lpBZFNPn83Ub
KY9lcxpyvQFNr2MSvsI7+CP+tEXLV/vZYmYlFKz7YQFC6W3IBgPnCCz+XL6fBU4x
nJeB1DjmOOvR7xcJOXPDk71ihpGQJfIJZtYpKPvNVNKhD906sHF06YPVA7aqaI7F
NKSJEIF4AQLzO/oQDmccaFnv3fQhHSu9zJbGOtksWCPPt03AUsIGnioMmmFuUe+Z
S2CwjC7oMnztjE0NRG85w0mEYZGtLggBt2zpRdUfxN8usyCoydztwg5tv3hmeS1t
uCO1E69kbffFcdTnHYMyon3Hw/kCx76H3BBlQnOLuFUPku0+Pw3Cpr+KCbMUK/sp
1FJzpnIegrLLW8qVhU4JnjkS6B1JFE/8MknQNuuuPox24HospuSQnhvlfShTyvY8
fXNb59om5AmF4a5HBdzrFfMyW6DHFE5fNXqw0AucjQcAyWmabRGbWOJ0UL/f/Npm
iv8xh7ZIV6ob8fd6KSEvfQFnTTdX+st+Cbb551SQCamluFVy543wVlQ17cMAvX2U
rMGigwv9+nDpNlvT9siSKBoiDakR6AQhQiw4/gBShQw++NVS4cZUf6f8K10r1d5W
Z63dXB9xJR8nosie/iMP7Pe6jpEoAEtjCNdV+gIg2gVe9CzNhWHD39OpYix8Kl2f
kJ7jWaI0kR0MmQTLFZR82JVA7vaE2Qf8+wxN/nz8tcFYPFPDupSrbaNY7FrCKDj7
2iSBoq8JMFF1y8j/Xa89+qykKWRKpniOFshs9V5UI0fy6i7P6zoD0a6qp3MjSpBY
WF/6BQwe3f1Of6xxPfcKTdHWsmWJiaV1wvh4gCNAShy6s03UE6NzDZ0GLKnDCzZR
ZzoIrKSDu6dWdYjBQsj6hKPOjBtnjYvixtcAeYrICZRKgColQlonFn4BOT+RzIdq
HWuZl03q1mDaxIPbE8KNBjr/0DKy61X4O8EFXJg6RL33GfZwdP/TWJKSbFT4eg6M
maHQ3gcd90Um9cQTdm1TJHOxxtBNbgVE2phpCbJTGkGBuZkrEh44yqVDGKxK3YOg
hk+U05cXTqgQd5f04fdHp45CKa2BAv6BbDKJYxvRHLwvqk6Ev9A7m3kuaTQz82rv
5rNajeaD3bPm81ygjfRVmovA8Bxps5gzn3+/JxqYhqBKfybwBpAkzw6+ffPeM0/h
s3zzy2HB6cuR7/bBhHgXer0cZ11yAXJJpY/a1khORm/q5NxQAGbY5Fvq+NkDS5Kv
kdODa8sxWpOXHWds6qi6EtQ01xWOlpvjrDjA2m4LYW1XMU05vHbq/za0xKRVVwUy
D2j/WIXybHylpUbgVF/2mAX5Oov0YwD018WfiS/VNTPLEwjeG9QtnVgIZir76h1J
xhZjKqmbD7GXcT1dvh/PS8UYlIgbzQZBaSHijqjmELrAWVjRL3oAxTC8+7cnvdSh
XCLWtpKnRWbz1q8EPXE4IO1MZWuJQp1cPJtVyls//AkYIPjxcUHjU89Q+Smx+Iy6
gUlUY0wh83ZeRHEUgQAZp/mi+Tid0eXIrDkcg8gyEUSb8u+5QEv9jO5uBhrW/zeE
9kvjwnbEA8BtchwTRbE34Xf6mICxKuAz5NLxGuJFJaGTG2sYwm1YFR5dAPtmgBUx
qOMCElg59eZqjd5yVntj/UyurNZuOvBNZLWP3/W6cwCC8ECpaUCxBE1TMp/1p6Y7
gBnZcSePDsBZS8Mm94JhSWuRC8TqgEN2ywaOEdORwAMM3EDZKcBhMn+7/jTpspNB
Jz9TJc2SSUbP6cpmhFdPcYjh7+fRah21vAqhWZZNCdcOYFuw8K2xcV9Uz4iX4uSR
7qZHvUniB5Veo1TH2TXHScfuYGb5JsSie57Qc2OJkkaYbzqZjBhRQV8ZcsT2V/cC
W0Ui+NAbpGBFneOecH8Gmm/OBCR8fAhMce8cAWn44zUmivAyIF+9LyCq0Ku41zqp
knTJ3AqTiOvq07YBAJSyuxKDEOsAVB5Qyb/sClgjtlUvgaOZ/ye2NhJ2p1Fowyze
MWG1y3erhKougBhjtnGEKiRem6smJ7ZXChU4YKU4a5xzSSk/tTq0JwNQG7ySzYlb
+Kw0vhgFisNGGYBWwqfiV+DSlyBdFpfARgvtVtrZx8clUFLML0OMizefaDSdMQGO
tNuT4OgjmfRvXKAKV1rZFFgA39bu4GpjrS7D8ZnOJRUB9Mh9ufrWu94GjVSGEQ95
e+UwfaX5mU44palsQ0BqPuvr1xCsP5yp1iAhtZ4lxLfx2Q8+mw8IZtk33bvTvA7r
qdg1AH77MDRYpZwn5HSe07XpMuuZoq7VOMKm1y23ZhXMDPPQ4LnsOqM3x27bFE1W
QxgtaET+NXF8dFdoFk+FjP5kMGc/H3DJAjNSMn5kHKHcYXjBw7lecfszDitUlLyX
pXEUW5KPTjNCPxirr50wmbcZBvmYWkmHa5Azj5UPDY5khzwsx5WkgPGV8qoxwBmD
zrl0fur1qh4fKopFBGAcBKC3lFsVo8Sx6A3ZmIr5uIlu36UFN5IuNMuFXs+RMIzV
DXjNN8ZCwTF4jSzhAxq4/GY0t67uUsXkIo/yaZTOJN2RjxskRWsO8IqzgZlqSlPo
PT5GIo0VRrUN/glr6YYIxe+4k9kZWANZz1Tbio3ESo0Wi5VfqwPMBS2WTiJH81FS
82elbS5lj7bii4PSuuTsFHzvgd23121cXJ7yPy7SBJJufXQhyfOOzX6fah9HTWIE
81ynOT9bIu5LoetMUnvpHClTgxrVXF1spuW0qajzlxakaPQlQqC6g0ntWzf14RP6
lJxSbFLZv+PaNl5iZiGN2WsiMXf/PsRVEcFAs27Jft/0YiSMcJ7A3ZvijnOc1Ky3
TORJ89jL/zbcYO6yprnDIF/l1A4cWqZpumcNMpC+vDEWEVn8PXQJf2ILHRN/17zO
4QLzHudHSuCEx3Cq74rNTmQhbnv6EXlPWMr5256rN8q6pZKISa756yh+2lQEcYK8
S/TakNdwZI6Ul+gxgxe5NE54qBCtSwfurVjZkiFuHcoR1EPz0CR4LS6/oWpIuGEN
iGVaRgPc0QomFlpuKK9p2CELZ7v/Zg0celGSQGGzv6QZjYgI8Ue/VK/MDM01yJAS
XLbunfqA8ORPZjJJNDB2S7emB1Lhz9M9huHbRtEjqOer9Xgy0Bw0v+jq3sN6qDc7
FA+qJqWTGiqmUHPBgo02LEwB6BM6ZoZe9vMOwulBiewVJXJYRlOawFxFGYPUnwrh
ZoTNepKnqLDaXlxvYVEfGsRJbzFWf2rGpYYN1Mc/V0PV/9krWClnzjezlknCbLcQ
cZ8HLL+xWNG+SJzsGZOPcsn624IjemEzaw5h2TRvQ06DEz1r8KO2UBg3pwxS5zg2
8NXQAhv66iY+YNZdu5Wo+y98KkieaAEyoN11Lqb/ax9/73PE6b0D85dHIY0KznRq
0siggNfhLOT1i4nWRCq4KVtO9fI6jiqohm3gxvqtz6aNhbbqxwcnQY1x2IebUR3l
vSC8mRa2d+HouUuydy3bCR7AP1kh+sFUQOnWOxRwbRSU6jk9zvG6NY3yvBcqbIr9
uWilTWIzOWdbdgnVT7Harircaf9GARJEkWEGubtpAE24sxYwNGPbl7RENbIF/Ov1
zJ26D4FD0HHEpdGdaipiWQZqn6asO+GacMBhqQMyR1VAWTaioFq9SoP6k0MtQV97
jGcydi0vXEuH17LkPSdtctImquHnf6nG0xwz3gjWdcZbP9Ek1a9em/jDYoN3OH+F
jOVSSE8BsCkySlCjypdKhg5uvzUP/14TbdN1FEausRmVSG2+wvyxGfRcPwO+OagU
jJEjcEw6ykmy0iG0B2Sh4jmN+mr+ylbdcho9i8+TTaTHsGHNowSIBMwYF8fwztO0
rL3SjQGhps+wrO2JurGlxdgbLyKcblOeBl94IrN21ysj8V1xYNLf5O5yYkLzq3Qk
j3ry0ZyFJPm8KxvL2htRbOlxDTBvPi3XjnQNXDdnmoAcLvM3t9huFpz993IHdlMc
WuCr7MfzUPVx/1llb/1yBNwlz+l0sJuGCSmPjBEATFxv0hfyF+oJiPTm/SA6Hb+V
afDPxN1bfqEpSIep9O/Tnr8q4gKScGwrU8Fei7Jsbx6O3jFf0inpYyey8uy49M7H
Zd+2fYRYAnH7QSDhzYXM/NYfxyeGBBcg/bHjwBzQeLTiwxI7P3xcPkgajkATumZL
0w65ZzUGyTkKOOaUBG9MRwcfWsggeKfKGSOs6BPcm+JxLH7xCg0MoBHyUzT+yUkk
STIaVob7HtbqI7ydZ2GZNckpZMJMsVphIHCuRfck4po7cTUcmPBPtcorJ9/2RJqq
5zlxlHoTas4askUYtCAsuvpeD3Gg4553sEl89Cv11PB2aNOlY7lFFjsyGUlIpUsN
09hF92IA7UaUgzze/jGwIJzQbaF58iqXssWZE8UOxK9GYO1WM1c5RNPadkUKDtuB
W8+5kiOLOST+YZPFoC8BhlkXwho7ISOFWQIdKAhD9XbdRFGJ1RDJ3IXNJfmpBwZB
hzV5hFMJOWlyb1MwHCsyuwYjhDE8odmuCQEVQ9toXvgtfaeDwiPnu7k24QkYyuRd
lPpiHdXU6BFMuQLP94dIMnIHMKJ0OCY69La4mR0mzEVokn1VcOF+nr5cFW2rRfWg
OQlRLmZw14daQxTF4M0hg1etk3ORYyuTMz/m1AUlnA3OvD1fDNyfAGvC6CuvCPRY
cFs5nvygdd7kem/QxCrJ1QcJj9yD/H6Khhmnz1CTLH11JiJnej/uhdQ3aNqgfcWR
Hp6FD3f40rhhZG1loMliyCCcoLBcq/VNpObucVjyDDfwD1isdnwEQu2CDTxkqbc7
VsD5Mcnedwzu1pkM8BQoXEuDPlbESMA2Mi+4X7ZqBqOHLEkjtmIPFF2krDhic3Ws
fC2070i25dHyRtHOMuJ4cWfvawkTKZScqSR4QMZre3x+FqBzDpKQWHEGrWDDBmE+
sQnpJYIgaoCcenBgQEMaLQfdpMMTjv4UXBq8u+JoVUfGT6R9uNoEIeQzi7eoGUtX
hjxbgWWdg7Lmrln+kBoCn0nRoW8ssk7ispbjv56Btm/2kwHOVvzRFUmbtnD1aZ7U
j+wq3r7W7CNSPgMFd2680XyU0RccCtpVM+cQ3RP/KveEnUBjlO+tuxRWusu7ao2B
M43sio/DTwUXpZP1ThlhdBnrBDVPpGfn0jHH5wGG9jhrDC/W6h9eoRDBtX87raNR
uM7Cdts++6DgojFdH2t3vP2gH3lnkBg0BGNlwOUORBFzUXEhilwnscb/HyyPooz8
m1sxCqL9za3THkl+Hf5df4XZidIYecYZX7cLHF/J/6O0uShghxBgaF+03MPRTjjY
fRpJifg8JyAabt6ZE9xEsZoBZIMo/u8BF4PDNqAjrzc7TFHXIrY3WzCeU/KXjdoX
X63f069rQn/WfSewtm+T1KuFslJYmnn1z8R8KsZI0jqvVMqg9FUMv08sUsrudVfy
340+dQfLg9vulOpLudHym3NnOFwOhrC3PhMDr4sxxE5cDstqUe0Y8jo0NpCgUbtv
e9wHk2aRM7W/Fz7t6frIEWctO6/w7E8n54/NTWFW/eVBsTP25fYdWwAwUzkvnSmR
wb4vTV7nZJLSYlAiiFxQIq0cH0wt1VvgPPbjoZzBnd55ELvldsOAdIHRioiscwSw
bLL0EJmUf5V/tgz8iXKPscNOetzwIFfNiKceymzWjs0LEaIZcmfv9q+v2ahSHtwa
IIeqnOYz2z0/a+sDBPaoLwRySZzcPNpluGVN8iCVzbmUAwZYF/srjeXeNmMiOMrs
bojCP8k8n6Fi1joTdtZ8paEpOnEIaIuIzqRhV2TMs/12vTuiePX42afkLarvi2a4
AC95kfckNtUC9Pl+nywU12n6FJ7KPN912piQIJoaX8JKu427Y0naoyn0RfoN6aqf
VLOLc+Gu7pJx3HXPs07WMIsiiDn0T5AhAvO9pCmVDa8fTcT3tQxVFb8tL7fUHz7h
EwUiDC20qIo19uKQBxYzNbk1utXGKivCv38Jk+dfNP6wYjICRS4PAtBgZNB6H75a
qkN6dW5EAYmMtEpCo7z4b40n3jBgipwa89G1Tw+nw6WtDSDN33WX8Wuw7n7RwiMi
e6uiSkqzwoYRTpmieQ9ZZybS7aYSGMq+frqWsHtjnDvSxdbmPSZOFFwDVmCNnsnM
PJLjRAnME10W1i6iT3Wx7wyNVVhwB/jwe+ZemAi1RRC1Sj5ACRSJGFxnDH6sIKGg
6HjmEZYzv9IgvqFTmguadmorrfiHUCmQQCJQ2q860g02J4Bigyj7ojeKqXQ7qJ3K
439x8L08GqYDEoDX1//ybKYfleCGj4ZZZfY6EmxaGEpiKI7AHFNfj9qgg+RqRc5A
jgQ18jsN41Jq8LRryfu3our7DtEgXIn8c2K1ZokwE1JOSloKsywe0FTizAfMo+zw
9nQ3T6Y83SOY3l7sHAkmg86drIeyXKaE47fyZ3JypBJG+y72pPpzg378uVpaEfHu
zXstsuMmdA0uK3y2iH29OaOiAZ6YIv5jtcBkfJ+X8o9IbJDujDBW7HkW3xTFcz0t
753BarAR/cFJsiCgw5rNUZYtd+J+Hx37KPcfK56EvsHfBPR+pyZ3g3HCMSakqf25
FY7hYIyvw+H5g8pxdqS+uQFyAFt1/XCZgDCWtbPyuu3omOOi+R1qfA7k1enPYuBW
53G49UP8G8DNbIySCJBP8Vpwr86gPNH4TKPKSBBiciloJ6RwP6OP2oqkebdFU6U8
nKYElzMSWWbm+kMNdL+xSf62CE2+emYsVD7479IpQ7BotOzrTp+tpCCCR1oMwHKd
+vq1PBFlbV74TrQ4kWBnUOGS58fnwDKzbNW14ICHWMF13yDZTKCQWoCXmnmr17XL
Lnl2HJE0qBPiLSqjvdM3TRFMUp8u/MwVGXx+zvdGUFyZNRvgygUAtOVI9QB73vrm
nAvb+OZaoxS034MgqvCKlrHlHJ6NenJzaNV3L6kgOu+0u6ZdxUA0tENlMy8PsXyn
OI1sJii+dlwlMJpYE0ZJxeNMCsb/nK1YtYbkY5t2tdP0OsQ0hznfYM6vpJ8/HVt2
wITIlFT+sh9UaX+4B9NYarMcJXG+AlSxfEYcxLM7XKFRM4+Gj3l57OG8bmrDGa5M
ZUpNTpG+WONOb1o1HvfPsiDLi7yMCoVzHcnzJN0pvdg9qeAUvexa9aExNblIlFdL
aMRiG1vNEUkPMMdSb+5cFMR5A8KUMB0iCx4ExXjiXcntss5cMe4zFUy5XpyPNlaj
/XZnz2D0LFQj5LESEstQJJtB6rKyO3OOA5AvnAGDfRv/3WvpSUQVXh2R7TLesq5n
dRcvPRMNgfvW3svkf1vmG2SjCvV1f5WAZOrwBvUkIlJAjUtXj7gsOT6DDip+RkTs
4kk4G1OGGmWW/KVXYR/zV8jLFNTA4alLLZOHtEoJYPkgxE9q7gwCXKt7Jr87IlfB
+wEQs4t8liFsRh9uLKbAQhft6PekmCvxTpJ8O8Ndb+L/8dbqvdvZSPshSP7/9cgG
TSIURTJk+qhsyPK95AwHYGs4Lgb/9Fjui7vbFqNWAt9v1y4R8q7hP2FhUbCFPixW
5XJSN+f58lzwNgZHr3XBCfUS7ruxxR855wmG4k+aioYZ+P9SqOwsR3RFP2nqFElg
pJBgoWZ2Mmtt3AwOWrAJt6iae7pw2nYn47PAU7VBjuNv79CFfAkggd+V/aNa4hWU
2XAtIBA7R1H3havY93lmqq3eyulWBy18jLPVdBgAWdoCQ7BBP52KDlW//dXtjfpH
G0E8J8mFFgNJXDR3TMfAg9ED0Lkybz9Bpeulgva9oKAMrjrkjeZV4A9Az7SIzBC/
SktYjtfOTYZgKnK/ksNIU6GV/BlyhUoBz4e89TkPlC/X4xHzCcGSUauOTAJWFkeT
ae3N8AKEHFXfwUt+KrdayUbVjYZ+TK4KBtylOBSTVd5d6dTEdNXA5wGr+e+yYJeh
8f/lpKgKSSOcZuCLPCf+uNmOW3skA8PHxBX4SUgsxi9ArOgO5c5VYDV4FfbEu1Ua
0Ywas6PJr18FgvF/5USnRNaW4SM9etFXB+6eZ6/tRKCqwcvfBlBAPViRx0oUIjY0
Bv236hvYOl5qjCeCv5+rm7gqpN3IGTfUKY0tJAFklXWDOSG8BC41wrG1L5/fuXq3
avgi8Fvv1CRwF1u+HP8t49R9O+oN2JAc8f5IOCx/IBOKsxFcCjYmVIXdvwP1s58V
ojNI/2E9/S4PSD/YfNLq4MowMcP1N1UaZc8XFd8n4/zoil6Qf0e7ZgjPJS9pSf+Z
NPVyJlQs7gNFXV8IxJWTsxoaqGmRMzn9y9/LPfM2D64PUyjk+Cgv+qWIO3AbcCWl
tgPPTwpgPrS43/hL2g1fByeOD32PikUMxgcqCS8XqNL1Ge2PrQYsP60WUM1c5xLb
Bx2498LkuHjJfmaYwDDc4HQY4+yiAh+anaBnBtf33N2O6BLaHcOInt8WljLdxChN
CFSyd5aA2WyBzqxlOygShwE9yfFhs9VXlG9472cZVHZ8vx55Tq+nyIoYjlwNUdS6
LPhCc034NR4hJVC+Q1x4dSXUR/d77h4+Mlyamvz9VDRSRG9uS6gIhuV0wk/tQzfE
mPLL+0oEoO+qTe9k0cEOboacZq2sjrHQQvxe7/TuNkOoI6qVnqZG8oAeEnjQaP35
tpAgegnaq9hyUSZ1+wTXbJqWL4jIkzGxHaZYnO+T8aTFDeT+f5xLOUsZUTC6LSzN
C9DO4kzZW2ttTTINIhA5h9ZuuaetXty+j9U3ZmjXAow3yQ239Vc4UPps24BbUojM
4U9o8rBLYfWzD9catsW0Rbrahq4rOUqkIysp5RcgPyAAyiwfBcUhB2Z1ZCyJaeXS
CGfdu7BJwQhugfFIcfuMLPIV02mf4b8UNdvY6CvOpitVnq1ZvPJK6qbWRDB3SDVa
BYKw/nqLbm2r/sXgxJp9sEDDD1EtzQfI5YFu7OVJ8F6SQuxG/6SV8jekIvENcJHU
+xXGeDobpv1bG1KnufSMyt2bXz2H66O+dppHWLFhYUmzSbBbZKO5J0TRtSRIH6cs
ErOcq843sUuXQ9SjFQQA+uyVtmjjgxN9lO5RtSoek85p5Qc9ndoKFKFk7km6fZmh
C5zAsBGqb7qWQuLfvrKvFyWpBl5k7+0eTPLOS2iYXO0/s9nkn/uep7EfRcgZ5ke6
oKS9imkVe8kYW/8o9EU8iOsrJEY+9FWZCcadXhXJ8lndjS/Blp07bj18ND1ZKyEY
W2fIAtjh9LqwULKPIcCFxXdJypRC9OHlIxPOE9pRrnh/OYEHpaG2DmwX4HziwDyo
8AhB8Mlgb1vcR+ZrdP6B4FEOu+uvHS96gDny8OJEqPdn2baFOR3jgzUIW37r3XBB
7wPSKVlX11VgF2nEqWvsAuaU/jabi/lRqE970kGF6KPw4+nlGPXs9vP/Da2Na09G
HnqhGSxKk3PJd857W7LKJMOg3A/ZMntx6DMj93TZheSg5QzVxD1nzHtfMTA+cdhf
pdej7tdToOxzGffoDBo4klDV39izsgcbyIzRLQRoz8Q+yuiVGdGd1SiAspj5Djgi
2SQApmm3hUfqczizTSQbBk1eWxXOx0K97hOOtqDIOEGnoTJfDEkEDx82RTSUTXfQ
+kWlgYXl7+5Ee7EtStbeQAbQ5vxNd4loJkYbusl7zfqoyRZjhNoXkZBeUK9aRZ6y
jYtmmgMkNQOLLOf8hVK1eAtsKsGHlwhv8Th6zCVYY+nvq3avPOT9aP1cquWJjobR
JmbkEIfTeaIuUMibvgwhjYjQApUfau2DQ6yX7Glyv/T4f3ELQQIqXaLrJ82HzuUY
1AMgUi8/w4BL1FxQywHo/H7Kz/0mwwecHZPV8g1xZjUnFEAeSipn12sSoiRhaZmy
GaHi4EZOKtmFfXtEVXXidLGLgNJXa14pMdxgnyf9DCbYqngLXcMD4K84Wy3r/LJ6
ssWzkswz9kpLEkXFBW7jVtwaduusFEcFtlO0I6wdvAHq70KOBqovUsorB5tktA9o
nsLFKYGCqMkvZ7XIOcHl7fcqy1xmTZKIbL1bG+MC+uvBVkMZmpQuyx7KAGEWOk93
2Qn1R+CHIv7iK/TGOXDVjEt6FJZ3mDUzaxrRhCrdAsDsQXVfTt1j12C44ELco38z
dCDlxx8+im3LA/81kOI40fkBFPNzpmCI0NH4pN8AxrJN68myNgkEBu9bTG30AUTL
AmNdCGr+chIzlxxMJ37BjHrBbq9N+XVQ+CCtCywLer4zw0MLSmNyhX9dy3DToyvv
aWdViIKMWxasFt1ohdGIsT7N9XwmaZMtN5ND/Koksd2LTSNaTYjXEkYikKzX6rWp
gLuZskFHjfGhsldHV10UAka8M5s0pOJFejeN3yCkEnBKCA9m4il/XpE+MylCqKHn
F6O+Is/IvmOBrFr5XAPQG64YUKgSn0a8k96X0fWJy4mq/Zxe1d7ZOdIDtOAUAUjM
+qmF7wNFmyLKBw650AUe2b0bDhdVmLAXZb5ytLn0r/PQfWWHkU9jVBRA2JnkvwJJ
gnaRVz1Dm4jnrGfs71uvrM87av/mMQy08pdzV3dn+zOPpEuNs5MjGeCheVrX1Gwo
hpI9c3cg4Ew4UIX1SLFHOqKIDSlRX3+Ex91lOiyrXheTx29uSwSHbqMcyNVb/n3W
CTpGaINkhHOlFzpUc0zK597YhcPiao+LFhI7YT5w02W3mQUVYAUimXKK6YTw3NeR
DTp+rgfNde964n9fRb4aBkJHM4Ar6udIeQlb8rwexr+g9weNS61q1LDi8L2a2Ia1
5BZ6MafjFI133IwjBLnL6SYSr4bhpIrmirHHdLL4TiNHJ5gW6M796Np2RX4bjd/5
BHeSwMSDDlmkGgFGhK4uHCYwpRkQXvTbwUJxfoGzmSnVOlPaZpR0Wv3wcG7SvePP
i9sK92UX3snVuFwgofWxHEIPzXzJgUaCnVQORjJLVzvbJcdiLU4jFt31+7IOsD13
hUEv6hMgLVJZPnOlH5suUQv5gnG21uVU5BQeLgg0wY1MM7P+EcxhP9WI3GhNpYsy
aHdCLMdBGKoo8VxE46+U9SLboyQvLOT5hqBdMrh01nJf/e0DpO7dotUMMtfA9hYv
HgQFrZ2qJ3Qvq4r1fugCSWEZiYDcKTZQ1rGzEhvjKEcoxaN7kusAg0TZROIwgk5j
7cqNSJIfq2nyFIY95NJnWO26wZ4qRRGquFx5ZxxNOHy5E5R9qWRMZDkKvKeLLGKk
Bd2vXaAwVWNAuIqoeSPkCIXrYQcWoNJucBbLqOie0VCY0DxSK8tlJMn/4nTUteU6
QDE1gQVs/EU4rbW9JTADSshvAeeHFRAncjH9WXQKi/AySgNkQ09Sm0xJXaWDTcDA
JJ7ALDNKzjayNAiq6+jKJuJIcxm/uu4ExhYB2/vBJz98Xy4pD45iTfh6DAhdKLuj
TX/mh3XHBSj3R1Mzfe2d201Wyb+Lw3Rs6PdvGQ5PrMgMR+BEuFu5oEpeCIlpq55o
QaRjjmxCPLlLOZ/PXFnjqgP1tyH+iCWUtt4iH1XQJCoctRoiJGoHFTy+D55OpujF
dx9QVJSSx00gDVIIUR2gnE50WrhsYnOWU20ceEl9oXfr9vVKpNW/SkCv4jL27Rr4
MR8OBXVEacKNCDxg/PpjJP7oMcfLZjlaSiS9SYdzfy4yy/uyiv+ezKdd+bAdvsVg
uaxEtz+H27W41pxL+8FocL0BkNCRKjPjmnXun2Rco+zgPpeFbgDH6JCSG7RoFC/Z
KbpM66+p01ZojMYida/qi8vL9f1uGbBXuYvHsCyk2D9u94BorlCICs0At0h0dBz/
iYpcXn8trEsYrKLAJi9nDMHSDf/L+6kk5Z+9U1HM05ZBPDgnU+9v8BK/G4HQZdaB
WPMsU+KRcWEQRitzPhijnOMof1iJ7wYurWm2aWIVnp04NIPZb86zwlm3APOEwZ8v
AnLioZtAcGLCEqpPenIEoR+BIFePQvRfYnY2IOJbLr6PgmFK5k3OQxCWGlj/F4Bs
iLJ+JGtESgPYTizHuk9h7V/XwtNy3tcAjkehKHpyeyBGeNc5JrBBKVzYKz/QVfxO
2mA7p17LMWPTDX4Ti3d00H7rmAYSeIwX/KErjEG9ab+b9XQNFO7KESWKjFiO4r7j
syok0xvo3YgNCBWl0CHnodpApSjxffh8wzdfMhk4IUEggTz7Len1KBESFg4chv8s
X7yaDhdklxl/qjan98aFBi15bpIjtiZIgZ9VmnedBC/N8djnVqTHs7P3OqoN1Wc6
2VPqW3sAa5y2QfaZsJHgsLUH9dvWqF4L9Hz6oKEoEiGLsP4H4e8JpRi1CkT94kMV
nwPqtD1HnXrufHgC2WMA9XmSAqzv14o0APOldMGhHeeNYy/KlioklHGxAjczAGwj
FdNbYOVvnodS5bSEPI5JraSt8k7ip5niN1PD4tdNuYIyU6tjaACZPrGYlyQECQqs
Px92iZeG7pGyllQpc2NfGb5rxbnM/hKdMNI/t7eVEVTt7z1g1rZFDI1zynU1KunT
wNiKCBfGcmN+1ww/MIbSjs8jFMzY3IvnyIi5CtLJgnLbFJt+gC45oUfvgJvIcjzw
KyUcTc1ZFdqzSIOrMcjFLg80hHLsjOJZKgcLWcMRgXFV0EKKUEBTMtCLCh+ElyyN
i/3VF//doi8HIvt5rltl6c6UVMYgTjDuN53OL8Cp3l5vMpMDuvvXVKxaelIiHLmM
1SYFcBcDzRhbJJgLpLO6YvW/m7OwcNnLTzCdlNmylkS7lLWeAxhSUmlMr9BTqmu+
iPc27rB1RPzVlape6F15hPD0Q9gVvQz8FAXntUQcPtElsbXqtF2nkSz02zkpugij
1pv9nDspv70cFY0RaUQqKOAZqgLeaOW21ZQa0FmndTYCxm6Ve6kulXVR9i77Mh9g
rTzC7tbD0BZ6eIbffd5XDrPV/j36mRDkETavGrHStHbcfipMC6TsAVtb9pMl4Wbv
IDmpJ3ZoR9Is8/hFbq3nhRCYR+OvlsonyPDit+nS+gdWLH1AYADrC7jgdJKgyqm0
447+6dcqA58GGq277hw7vwpHOBsTXFOpIWhkk5Qx82I22ye8hutQ+CSuKr9+PjoX
P/FwdcReqx9eq0AqE3+TEtmNOaEc14CPr+RWLwLLFQ+xRc8om6KYzJ58V0ajqJLH
vv9rQne081hNjcXTtIU6wtkT6eCokh0o1bQ91ysEbRsm/8shXVHU9qe5M70JKq5r
3ZPE24CHl60bKdozhifNDPcUeMRu3lJqubeF86Q5Nmivbff48ST4/eQsuLLE/f2J
Vo3lanM2+wIvjlI1jk4LUtvqrhVyohOqiwJiAo1kwKHxtkO2y/dQflzrZIp6aOEV
5IIuhNt8Zi6ylphdv0ycZfMvy1aE+DGu0MPBFTv3NNcOoM3XMFhk9FEX6yvJeX33
Uf4hGy8ZXxVyHLreF47yNtRFJKwOmi7wirfPozLupdGuvd07wcEMhYqz4Vb9YgU9
pEBE5NMg4GcKi00EB3mcFv/oaDmvD1YEcKjXP/fGmcc6hpuwboQJEuWw8hcb4+d6
PV25x3ovuukCrwWNa9YxeYOsepkZNW/Ll1C+BwmnC8INqtyrPqsPM3gyrAgMCiR0
tGP02DJFO7zAfLVLZB7W13/Q9sn5S9ziSl3iXqog12vlouW/gdSpfN8Ijt87tSjQ
KTnfQg/E3wY17TQw0qk9kC0S5BqU1hS1HKFmEk9f8VvFB6kbbOuToNYFU3y9Iie5
sl9Raf8GdLPFGb/E3varP5mijJFzAt0agufkx+PahSQyafFT1vNwQtzlbhyvlx6P
WfGLMSRVA8ncnJIDmY5mgXcgSAv6Td8qT4dT/iwmK2fxMItaqy1zLMd/FFGo/nWD
JeDiGz/ioFCnjDLBLiN4nE8X9vWx/6b2P5svH5Qs/pSCO94kxsONBBkM3ncSZ5TI
+u++YbT+ycX3l7ibhEUJqhukeFIPZ0XvC+ljEr+Md6o6RuN8cTdq4rQhDZcG361F
wSn1wD8MX5uViXie1r93US6n3V52mTqZAivhoUxGrtMO8KqdL52VQSOCprX/6EHE
lY8A9Q7Etf/NlgAbpvVYubeuYjaC3KvGhuk5sLW1dfQCf73phgQL+XVd0ZeqbNGr
pjgSXcnWJznE+PGojoHQg5ELJMtHyyLtcqtdm+kSbHiN4cpWJgzj+8ALLJjP8mod
TVbq7L4R7J338ourQtORxES+J352wUE8n4TPE03wDY4UW5BoCr5Zmh11YKiISA2V
paMvMN1xhwbUr7spHrEjhbvMaV2j9V7NdDwc+decqAcLxMsMAhejiW4jzlwG4TV2
oB+Bpb+78e6r2lcNSGJ8n+Sh/K07cW3xnJyA/d7mwYEfetqqIUGylmXGvwzoRxX1
BNDR5Wukxr6I2zI8+JvvvyLgVMW9UATEsqAiobu5fe2GNr1x7ip10hSBR8kxQkpG
SFMs+oXSQhNGSkzOnz5kRdLE+bX80/sPdr11OadjgygJxJF+ODOvGxr43rnv2nT8
0a+pxpM45MFcpA2q7czB0usF/jc59+UW1tMOjE2NoBUTxe8gYke6dZHiRrAM0K81
xDI0KPm6o/LqBDiYhsBbYGXZP0EIQF9gOXTOhgZByANUG1XvH5smqSCC8Ct3lKhe
Wvgnlu22k3iDdXkzQBeJMpKJJwbmU4V3AQ2j8CqihcXr4VS4CO4MW9jJau9C7EXL
c3Kacci7OV/NXfeb1ZJQMEXCd0W35Ezr+TDl9hXgYZ+G0iFW7a/TW9dXI6RUjRkU
0sYusds4YGl+FnMgBxdbIQZooGyHPlg9bmMz4u/gaB2f8EGhejOntyybrqThd7Jh
Cxo9nfvjXpnS4EBWvmbud8PNcyrtjwdxyTpH0tBWWtThWBYUXi05ULrbEjANPKU4
bm8glrELUTj9xspunp016kpL7l/U1HN07d+CMCj2Zf8uw+r0CkbhMrIGx/Q86Nb1
k/zYjH+Y5Bt+iVNg1y12uGS9Zv8btUkQakp0YuT7rn3iZKmqC3sEXiIlBgMpT0IR
BcJVs4V3PkshxbO+v4r60/vpyDPAMKF0v1ZSN4vnVIp1k6u/rU/6RJbCqcPKl1uc
N1KcIVL9A7ez9x7XOOqW0/kVaKnxzvS0Eaa5ic/b02vhOsdFHX8QmpLlSsMwx7SC
ggfQT5LOGdC1LYj01l37eQtt+akELT6X9nUqVy0WGNHsAfCnO9MkaJnWtvgxWvpv
rq7N5Uz3lbK75BRa5kHmGgZqvJzAm4AW22r+ryP1NkhQernICKC4r47/hurYRtkH
fYBAKycqJzZw2BW01IgiP4Mmj3jGs0Ja0MZIZAhSpkfavoHU1oA5UJyDU4aLDP9u
OqcOko52TnTdzaz2SXPI/mdcEv9Jte19YhqCGrsojDyfe9VE0Nlxuwjp7klCSX7n
WtLhOlVc+ExiW1OCycQ8fYy56kkuEHtJPHu9LoqA7Mkp/925+xmMyW53VX+yQOi7
BQQFs6wAfwvTizI2pzZSOZLCFu15CMwaiaHv6xxbdzFTTc9Cti28odCre0Qtmp8s
oc0kRSEECDtYvNZaAiBA/KTxxRJFZSwHuX8lOCCgCq2Fb1Q1avgR7FsGr05Q1ILv
rd7uZc6kHaLyphkGDyM0ZCPXOvlKuncvH18Mw3EWJLR0Q5TsANXvbxF1PoUfaT7m
RBqPPy1C3ueT2EkV1AwMPylfR/HoOxmMdlNlmXOixy6Zv8MqoVLiCiXQEWm7fjPG
nuqR8BMsJTbDlHEOsORRF+FCrwvoFGpmvFyg7SI5za1QhsghXVtuafy6LZD6QZYB
x8cGrtn/Q6YLdipCU0Yeqiy4J6EPyfjtRZEBYbTwEExWzLBbD1HXkOKzum370nxb
iSq8Jl+afXddcECR7RvuZ9TuazJGOettEeBtqRXB4iv3KRwqLDQHDROxFsALWT0L
Y2e1FRdDGvpgWy12AG+TFsrHh5QIYMDHqXM+CoBZCkRH6oivM/z/wB6GkID0e2tm
prqB91JqTAC3GZy8KxQp2h5Z03fi6JTB2dFvDweIC16ASpWt/619GxM5UVqoEaoq
XACPIsN/NkO1+e5qXH4LJL3wJf2K8jC65bjqP91lAiZ1SlY5UjCIC/aORN/ERAW2
We4iPTND3H5h0jk14YDzn7WS29+AELrWCG41E8y0om4X52kIfiU1L1isn5ZNQakY
5i4hCLEV8YWQG9Axw+2icoUV/BwuPUXOjYH0/zMbOjffSYIfwroaBURmT7f7Z1ry
EtLJ62Kpofk6L6dwIzk5x+172F33kuTICFTzd5VzxxhqtaN7bJtSlQjuFqVih3I2
oNPhLFCcvTDX+0g9o/uhZa10yrwUCEES4av61Tq9WBAnncKIGBznn0JaZWKdk/z3
4VSvgD1ontNKnV4j8bHxtDdbxyrG6/2Jy1N+8C170+ZY4WdlClseEzrqlmPXjS3y
mu23UF9i18ZRN3g9tOL0vXY75c33BvLP1QcoW/UyZQXIgQI9vd9Rlc2hcRPiFHCi
OdAgiSz6ZFea7J0Dtb7qYrfFgRQRNLt6gGaZAwywwEjNQAEojq6fE77mc9J/q0Gp
H466EZoiiR4+QVKYX3xw4QOvv3CHKpj7NVcEeCnt4VJ+vLi614I8WESPk9uD23s8
vwB4VzeWvFU03KeYyxjagJxW/GYTvSCmqq/UMf6fVreglEMkW3wOUKSOWxqjSDrz
SQtyDiiezJYU3oveknYppgJ34oHu3ymI+9B/3VhZOs0LG5V0E1mdiExdcL52xrWh
9wXCVqyLB3ZgdDLcDAalAASg+rcfhGeBOWFrPpLs8BVYne0d0QwHh3mk0zffg797
dC4yAC9UgNZJRBl7Tj/3PndHjGWTBLWOw95Vvvgx5WpAzByF+TlHxiLJdJtB6vlp
OoRiNeRhk500nKWka8LNRV6ir21U5ScyCXoenQwpkwdjlS0X7AHltz3EMSFfL43w
SazIkG6RWNBseayf0hmY/XFTZT2OnPg9GNQH7ghfLeydZ5LXFb7OZHxXxhOZwFC/
dg3mt2aRuhWzVc0mF1gexRwlXArRYFYszFUlfVbDCymbJ6n7gFP8GRAUmlUYeXyd
I+I606EmmBtBHDkkNSAW4mba9eCRa8eqRHsfHiV5QoAS6bupqyqTtR6oS70250ml
ztWQz3PKr7xWt/VoV8ZdC5P25Ukmse2f1ZoVkcn1aBVCcF4YLYAgNG6ONM6j7IsK
ygLyx/MxICHLyN7XdyfKy443RApxI8/yb5vWuLk+obHbI6WjY2DfcfjrIaDfGj0I
+DN3enqtTob4/QFFbOrNVIKMS2vbECY3QIqpXyZ/RxMFbDoW8q3+w7yWzjcS2kBI
jMg63WXyUDnHLytok5N3P96vErcCUHnQUniKHg3xSiG2RbTukYDNcXtoxpJKenxc
OCAeyt+XQax4A6nJRORGtKx/pMAuAZ/iTpStD/o1J3WlkuFhmsDoLPgJI27NIDux
I7H7LcUTcT3RKQ+1xU37bWpvkCEfsNifBWSJEF50Z2s89DllG7OgxzznMGBQIppr
ZsCAktIT7pDR+qCr1eJ2t5CxZsjdeeqKkdTOggHRG7J/hSmEsz80/gfZE498B60H
3qeamhqJS86Rcy/0Er/sRXpGNO8afIv7eer9gisaWA7IYvqomaWhcmaiz7XLOBLQ
5eJ8UGZ57dgPgMOdROHngA01RBu4QfmhUJBk+Ch0LoJHP5a20vV6qRR1wY/wWuIq
wU9Y43YCw7NL633EEzgKKaqtGPzwaWuKh1azWDrZE9Ya1XYslFOn2k1X640K7sIk
Q61EU0MU4NPMmGg8jAq5fO1NsoTWDHplJZYr+5shX3/esNZ9vn5awC+Efu31F++f
nD2WxxbTVOxHvdmhRdUdDnPix7KwhiyoxDNt19tTDtC5hPjcZ44rD8ogPgRmH3aC
5BYkRyyJSOBqyB+F27KE0XeN/RaUzwwdIx6avSkOde2kV2dMivo7aSIJj+NmaZeL
baOBnSqOx5xtVza8yHkiVl/Pndum23EBsM4K7du+JnQ3zjITv9qiTCqD8KYIqwXH
4ifaSGpdLhcl8O7Ni0Z/9kbG0H05ZojeyET+kd92YQae21kG0wrT7nDQp531HpNL
FFC02O4d15l3/4B1ZR3q+CvobOzrya53Q86WKHQKgrHCaipmyTDELsAElVcpjlID
1rEaG4mkmbsSf0HTUI2sV1igxC+e4GsFeTeBIFhCQxtM5qZYz2kv6Mm3fTtnht+q
mC7QBBqN3BmM60hCaqIdO8G+By9yzXXxLoERpNCoEYJcgyfiMuKFzqACea2Zg/LK
m8O8qRxgIDyyLfPqB+FZy02tz0JhJSL7Cun1bJw21NpqTE2t4Kq5VisshjnWtJ/w
+/0zQKkGhj7Q6ZSnZV+U4ZTu9sJ4GXFWTM8ypvI8E2p7orF+gdv4fa+TZa4clPZF
O/cWSUM6oPYOwCGqExXo2Y+//LCqeWJD3FWkTp8zlrI6QkC4gWb7jyT6iuysKk4f
fTMxKHzTHMO1WxFRMlBqclJNWz4DewER94IYiP7eM11xyN3Xxu2aRAdOjnwDKuEp
Ig096vgHMlpdFCJeAuGBjF4bKik56OHj4uv73Ok5wJpD7fRLHQcMbkdX/kerGPpv
KRYzDQb566L8F23A4SDfexgRgzbCu26tcrDqiJQqro5+V/IlyzDe1wckrL5dVdWD
FML7EjGvht3B8cVYiYECc1Ki4YmXpCCUR6GJiehQaJr3OGxr80rh6vpXxnSCczsY
1QFEz/dZ87N0/CF3dl1Jibt7GBmj5ykZN+tYxqU/7k0tDlp/BoT7ep/ZHHLg84v6
7DzE0uGIw89bQAR0uYTehil276jhxnx1K/7WKB6iOw+oW7oJ+OrB4xUKkNVp4+mI
EmTw9gaf5t7SwqQ94FB9Lg+h0yoJBR66OEGMPlwCgSFwdosR6wRhQyxAIQR6PhhN
wOzZk2+fqJt0QobEdGxBLhs1I8EHLz17hWUYqoARPqX8RM+gn3jLLkkZo59XEy0V
kIzWf9J18ZfzKdZpDFFDJYigQcu34FskonnUOpPJkS7pytQBzMzZeV+MRFJmzjDG
EQM+D4/uww6CWkerfHjGxg7Y3jF3nscXP7YywEhkdn+4YT1QDzXv9vuItycKIDYS
z+DMpF1XkyKrSwpuYX6kd9WH2QCMo7wWwFUE7vrCBAMYNv5oDyCw82x64SR0wWcV
6G4Cmqn+MwI5g4rYl1hzRCkY+7clxRjxl0Zh+7s6Ms6JtbT60+pcudARxu/0r6w0
Z2R0d2U5ZPsx1U0HxZVFXUAAVQOxqhMf6nVeWhYMa6pL5GXG6UYYk8o2DCrtb5g2
Z98WTXWTPRLMMt/HKt3VhGM16c/RUrO8GNcenWINT7kex7r11RsIiqlT+qNs619M
2wrg5qX7PqivKagCgkG+m6bKgd4u+ZwY9PJamCXrqnrWez+NSvRRXyIDlRd4E1c1
madHZYU38lvl8BCiDcgoBHyMrWTG1ip/yYX/xoS3HS56Ks5ahucDRNCG/lHQlPzK
hKuEbWpgWUOQw2kUrvPTjpgXABgonjMh5+h7LYHt0MB6K8zAxRqOMri3gGDZ6Iyr
nyldMblITNMnbEM1F+QDyocvA9H4suExRQ3sMHIJk4pjHARBPWHI/MJUyG6qNDhf
VGuMF4zlWg2WStJveXYU41rwM79d88qTOn+W/JxxBz/5G5LFMFt3qkQW6KFXEuEl
RjWV5wmZee19XoQhbGG5VUkiFMP5gktEFoAf+Wvqqyf3/4jDPnJlbH2AeqABCNv0
gZA/zHilo94NNJj4owMutNK1hVlBVkuEb4IjHFcg1fPUBdf9Z7XMuEqCLw+1wFl3
9JGwYEit6PHUBkkxQwwIVnWJ/W1zZIFwYHnBtISzEhRj9d3PPO+2aWdalyzqPP0T
S2LI/ISt5dE4mjtR+/RY2XCHxFEazDKl4PsdKLWL2hJ6pnCyzzK2E6MOjgc2ggr9
B/rbW4THcTth+bckXOMTJiB1ZO2wyWZ9CpMk9bWMcwUjLX67Rd3L1xaPy9/h1IcN
hQchFut5IPSPCrpAoSR/0d/Za5clJr1qIoGkPhbHBNAapzB45ouFsCWiUZZDPoEV
lZnzM4pL1liCdJsq/WeEf2mGi5h/IYUvknVE06USFJ8fKxGhk5OCohdh4+y1RImS
mGRlexLC9BrqDEytAOYiha/jtPO3bMYtiK0mMdUEt34gpLJGAlAlPsTc6WJIF4UZ
8DbPtUYigEOYjRfI9mgOno9C1TUVdtLruTJ2ZgfFfS8O+s+bIZa6qrXyBOK9e+u9
7ePuJarKL0rUpr51Hp6Le6y5ZMlOBLXL+GcR9F1QeG6YIEGK/8nHQ/mg5ngwP2Qz
TyT55JC+VIIYy0RPzOtw0xqLn7SAh5EsZX5mNIDDKnP+DT923g09/+hVr9Hc9YrU
ID3iN15Nmxi/Nspy+mgJUCb1kpo3K9wta/3EIrtoAA4hp/F0kF/q/PXrFDhg+Ak5
eG+yFj6eog3Mp7BstnI2j2QW87rzguViJqJLAdEdWgk9+lkIQZmGBxKPdix99kh1
PsesaCABXgoAx6qXqHjNzXNuqTcA1Kr4C68UJjRNGK/FtAkd/dwxkqt86f82K29T
68g+RiBxD/srtDq5nqVu+TKzIfsMbzqKWuvwsANoc1cXma5wxx8DjDmF8shdGUnv
88GZjtx+7TH7GIoRBALGNZYAAUuSrNVLg7duWwON6H1wf9QWimo8kekIlZBAAdy7
4px8ZvD4C5J5VEeUEQRk9W2eJ9u2cmRNMBqOrTq+UMEb5jbDeppAlpYvxWylhv4i
VkvB1o4GOy4hfGkvdo8n+zmMWtB50I/bCvXbcSZapNT3xqemW0/oLCuLvUniamqR
oTJFhvMVRqmYwzek0PWxahG1FuQPOz+H4jk82R16EZEyxNtNrEvyfQCSL1gKlpjG
1uWuj4711a4wA/uPIj141okZGd/XAHASHQKFcntYzTXluryg8N8chD3mj9pabeez
3FgLbESBUEsSmkUmYKzCvJ/0ncdTW+cacB3sKiSYFwg+u7NUKLJuS/GkoWJElI5p
RmSkyOqMdcZ05kCTDpMTjf80yxOcxSJ5l44xa1s0QcnKwtT3Mtz7eBIaOF6Iv6an
enUNBD1Rk/Kyb4VqX4JpulOh7IV2TAFP79wimq9a8kqnUhqvABjXZ7W/X/AHLmQl
/6DwLg3IeRgOZLVzT/AhEtA80x8ahTK4+c/+PHfnx8rv+tJUo4GAxeCelHrZ9B4w
3ka2ZcrymUhJqNIpnYmM6u8/pHeWy4bpWHHquEMxfzrXZpPhpR/wAVESMcosp2yi
LZxruLQk/LdIQvvVmht05vndr2NNp3cjUy+EnJAfQPs88BhSeY2QxD253SBhwSK6
3YGYA3Yw6lzG/Ql8C6Phfz3+37YCce23rBiChxEGjhrLhlrK96N3pXDJph2ZzJVd
LDNAYNkdf6cc8mk1kL+CKSR7UA4rj+VWNdzo9hWOQ2UbwYMaHl3oSmulVVXpjtJ+
5xn+JHP+ARne4K3oLAeMjfoSAEtqwOoCcxUbU0DbY+d4UgHfNj2tjk8rr5CCTDJJ
IA5ugXUffuX2g5it/ID1q45n48eF6XqyFWe9VIJSqvpoP1grvdh+PZYGssY049Lv
fanF5rp+cmjRPPyzVFxIlxfXzwj1NTdTt7pzt73O+o35GIxjPNBwq4v/t8khgc69
jmyOWvQvcnzWyPYLAWTnneIAmNq2snEOZyiB0V4TbJp1KkP+nLU9PN4QkD5rP97w
oaciwrg4YjTCHxqDQK9ZRiIvbGRESdm81SQFIuo5rAlyjYEZEKLmsrbknsIK5Pd7
6BpDWzuv4ZG9VC2jjyLAr/2El52s8R6hf1t0RshTAFBgOLaDB7FRsWcO1hOcOSNz
h5W+Sx8Tt5NByilVjBPIPXIhUgaaxuUraGvi3UQp4MxTRgav8kfNao4FJE1Hs4cW
J7C4GS273my1kqVJQB4viTPkQK1VH2YeJagHv2vnBgytI5sQ1+VV4dAkH6I4cnFy
aFXwl/O/Je9qa+eXWm3Vc/yN18L4zaMzDg7B0tS+AnOUuPTFq1fYG8iCKxubKn02
J1QMUGWubAtHVuLGfSFQo2+T/I9Z9kqBygQHM4fw3dG2YRX16iNX+ImcObvUFWLF
FksrvQsFZHyjCmVLBxRHDBmKdjL6tSPUoSHAOq/AVDx0jlnZwDYvhJIHkBCATtzR
8zy+aKogQud3GzhcVRYjpzQwseRV02tOC7tRXqXBpTxnAzPYQexC35H50NZUcGrG
nVV+4mwk8+1QV01iknBusLGc2uFnguJh6eyOk6hlYssJ0UdZbba6DX2ImCJ11bq+
BMSFJkMQbMxECpaS98LQaOvos1sU2ppt9hw24s9TRnWY5Rp9r3QqBTTHtRzqmzOW
oHOX7gIRs5WMPUHJ8gtTTV+QXKY60xqC1RFJ33YfLtBj2FgSZ8uiz627nE437v23
r/ho2v4OrSGJrizrlII8ciRXC2sykwMi8QRE5ynpQA0fCyu6A/i0G0J9CcmdvpW/
wu5yrdeUgcrurmusrhImiDGsaitZd27UmepeNtebvTrE4NB6Pwh69H0ZA4tg1NMk
YWzisShPthNoY/Zckzg2aKiNi30bibNlZRbY1HKo8MQfwASzr5iDbCBCZxHkX9W+
gONZVzH6bVek2nRN0yRL8pRIapKREMmR+2esDgn/QLHpVyrWuwZwQtAU9+EogOKG
KyAaPtVg9qwagFNhnVzhMQgaviXappkhnVzKlmeR6jHvx4SrTRzeyKax0efN6+uw
0OSMutPyeaJUCDStRf49P3egtn7NmwBu4dhXKXD+CIE0EkLNJsJEernI7jp06lBr
KAfBuX8iDLQMXlPHMRxJV6PZAO89bkr+9dFVFlPzf2AhxTr7vp/heM+FNWUyDOhg
CVkIxxdGC7PThbV2BFAinGlXFaA2rSY9lp1TNRX0/idCnP3TV9ZQhS9UURlXTHGb
BLgr83MFM8LEOvlakR/zpYGEHADJLi0hi9vbFxappyC/rZ9VyI/YTpWVDguK+/1S
crvrq/uPEeuk5qxhi/3pyckkOgH153B54QpFyc0pExYM0D64nLk+KlYIjcijctIF
M0OfQBqnBooyvNEUuaYI2GTYvKvTXXCaIOV8iP6AoXN97uNUAyNUyEY/jRrypEMC
6CgvjdhlcOKZuiBOaAeYFCH22yrmsehu3glczlObdPoxDFMHEZw/lxI49XVdJY4b
Yr3zqgyESWPWzvnRlo9L2X7ee+4lxQIwnAoOIUss3/ZAtcmR+04eGDf3zpGUKn+J
wvqbNyLe7LpkMsFolShvj5LbRiCthbSLutlfj/ocYwNncnvNo6AIBnhg7yiTrA8H
ziSqB+ZeqgebO4kDywqZdzcMyLHAsbsRIUPwZRnYPdt5DQn2VbxrOKitMojip4p6
353oPkf0arYe/WVFz/v/chlYWYo7t7JqxqOLPoape942QDiDxKyQeLepzviMkf76
2ufy1Y4S1avfdy2NCuSeWRqKA8Ur8yDtZigi4LkwN9oZnbWshjMmhUiBcSUo9WUG
pd1bR5p+nWyzZrHvZDbrE7KV/GSNezQp+gv/EKZx6wBZBn9dNtJAmJ/rtndjI9dZ
bspdcLz77jpEm6AzNHZsCtHDtnQz/78AVeIJUZua75pZnVrNWWC/6/n0Uak2OQmD
HXMlx/lXmzJZyr7fCWTnT+JvXilmR8bbpOuZNugAOTvkDZ+K39ERMRDN+wGyvbqD
b3J/rreuLwldMvV9tvNAAAjCBaLxKBscXAMABDYWX+NNrZtnDM4H4VwUuEyfPHcG
/hUunEGZpVsk7BUpef6HWtjGUV5VmbAYiRF3eQnARRPwPHKpFZdSCmMSqKswriAT
pCDhxvwx/izp02GgkEb4lkSxLmKxYQOmVf6yUx0cuwjQWx62LyWE2o2mB/J6+txt
UgeNRXnhq6R5lCAV/x/WC3m+CqYqL7NhLyqz7Q6RCy7l/wMVfZZr2ktDs88wmWWM
T9fgAHh4lE8xV17oq+SJhI7HRMrwHIV3SSzSS9k3K8xB9p5mK1aV6foGFgVJY3gq
feoJWAM/2RsanZ/xDaqheRIx0g8SOXcYe+SCRag+2jI1VUKV2yIrGY85IpHPfVa7
xJ0IrFNgbPvhvOd2crxNPdoDI0NIlsgYdiLvBKYpuXykawW9NwUllX97G2nIz+Wi
wevWBk7nBkjbZCdUouKFEPD+2Afw6oriXGxYImpi2uRXsXJD05vHp8DtBDBQGyaA
cEEpCkBonkp5uWEq6oa4htsA+JpCqe2UIG372vTZXyG5nv2jfr43Uglswed9Sus/
jxfSIDT23wJpw0ml2q7ntFlm8UE6LCXd8D7P5glW61XBs1PmZcbqiDnCc0GEQqU8
nZaNGBNK/mswjYUDZ6QzIzbLq5X5IAMheCFSPLrbyy9pOLJAQ82livpKz9n5d15c
lHfMWZE8ZULwQJMz+IZmRb5uoj5/pnArZIukK8vrXC6isy+z8nNu9cob8eqTdZWf
2NDlG0NzfPNb9C+6cqq0XtwKnm7n82ngdyVlYYSyd5tLxMdHkL9iCTbAqFWDmXLd
fTYwmaSgQoC0bZTdIrRvTcIJAZIHsaBfpbgHDBGGRdyDuwillQTMCQbHo1+A+2jG
tcCkJYDdAX8xaz1EUjvxf569784NDqI276NpHQ00aT8t95kQrJollnzBiuRr9HD/
qF+B76XYqGGIwEGE9Ce9XyD3JClFbkStJE76GfSuB9LjCTMO3dKQG+/fXFN5JamF
x0Dl7wm/ToQ+euvWy3jl7Cnd2JPFv+WlsTp5wk1fWj99eVYuXNJs2hcwX4E4JpFw
nwQijWYQVfU5Wx5ly8Vk2EOLXrzh2G/cb6Jx8MCbwi85Mma+7kx/ilSMZdXkfrHk
i32GqKH0OQKDTCB8pyXfE/TokqFtsUJM9EpvlXxEeHGqk1R9RG9cRpHGKudhis97
yoV7uVCGvvBoa/ZZkxeZ6x+mnY/f/F1tvbxat67BTavBiGcwZlh5m5vfIFjCl96D
s6Nw2eKWObNt2WDrHACBToWGqH8eKeoNgCcKQO+i0L8YG4SgIfircEjypxrjZiD7
5WfJk3MfXYw9+bsnYc7S4SWWnetdyMlZCEgnlsrKaBBBRWQ4Z2TtMMJ6dzFMOydg
y1fNQNM1/4TRVftl+ssypOGjHKDw27mnoB+rQRFH8sIt7D1cCH1/lzjnh+ULyWlG
IFcHtHrtCzqhjXO7AU3vixq5jQb5X11mXOWPEDjPqXDY/P5o/f0xvlImN7YPkrPj
chyZ69yN1qMjnVQwGMD8gi8Wd/mtIgJ6K+g6ubYc+n7fPRLGZShGfgiLKMizZMWp
76uJHHJ2jBKPGdryAPP05qPbQv3eW94CUDL9UhRHK7LUwCzNTzyK4ln6YjMB3LqG
yOi4joPOtO3zsb7tEv5Fatx4sD4MgjX+RpbPW1uTVzIbwj98I+ds0MkuLnziqjFR
fPlueLlz5RnzL4zr3WNyOEe3HknPuVOJKQgrjUdbzDVDJcRnVqbiuhCuFGWvTNYM
SHS//4isoedc3pv8oevrUNZAWsSjDVvEkPEm6B1d5gfhzexRFh/RIv2vgm1EhLpv
5o9VEnxRlgcK6B/wLiS6f1nLglMAoojZ5mglPbpXXwNpZU/eSRE7Tgrd9tzaZGjN
pfnv/KKO7kPJmlJ5ab22oirlMXwh4vbvathuKJWDAdAjFIvdCbFFQ0x7gCo3UGlW
gCWJMerWDisGucxQOZWCdPFWIDGw6e2xbqS1V+TqOgmFzZqgZpIsTw2Df/RrSc5q
+S+wJI0lLjD9THw2ItZXzOKz1SgS7ZAqRBHbw4lQ/0jnsHRDTbJmhUvgbMtcOrBQ
n86yp1MyIN28XzqXjGEfAQ2K0glxNddLg2DBldrx7j4G0iy6Ys6EDoC4l2c2mzZk
HWD4425+iaUZ9o2IwO7xEKIy0+++CnPEiHrDtoU3Ij841eilr1xooJMDzc8JYInR
xF45ee+EJeajXgUyc6JRkBiwmKPzXmA1V4VJ5ZxlOieNd1Ch5SGucx9o5lf8xdeT
hq22l/EZcF9EjQIqIayFDTexd/e1974C3+2bOI9fKmmmEUcYZvENPRGTkKqdD5JA
FzAXu7HvoR2UyYEtakelK+cZ3312ETGj9gTLBZXVzyOfpPWSXp5pAXptHyGyGHbk
LaFMI0eMOrPQwSokUE6dUMFloBExpgvIxnOKi/8zZXx/6GpNltONOyxNfslVJnKk
rmu3m6tdpUrFdAT9t7wX+7JTcEKdPbN0pEdDkXcY4dWdEK9XOSFTx8EwxsuKvOxx
aOWIXkSIrjSUgENCF845E+rXo9eO4X4W4JXhhR+U4PkJIxNYwJDs3aetIVCkRJg9
TETZzb+WZuxXzBKQo8KEtDC4EBGJrOYYerRVfpdLRjMVVxGy7pR5PqdSCHghNA6x
5vYDTa1J5VKfZ+wiGqcf7aLtg2UwbWxSvNgHXD6ml03QX6XE5fTlN5qanbDeSKhS
vebFujGqeCInkhKGymvafdDGXHDOKQYmFwixUgVwgMChmZtvoQQKVA+bQoof/LW0
t6KtbYy08Sh28biAJIZ5XLV6PdnbE4mGb0lssV1RvhO1ht8hwDp4WwXIGJKVJSG6
i7JtLO3n0hmgfQIxN7cM1Zi6HKqpaqFIu90uZXs/rztE0+r3Nr66DSop8ybl3Lle
F+iweRpBnZ3EXm8MmvU90diX1T3hePmVvS2Qx5BWoOo/aZVyd8Ob/UxG1FbkKTzP
v6VaJMUDiJH8ytCVGzbacaWDAJ0+VuQCnmiDwwGZb6O3l1FR9seDGU8D3wlCbQok
ROD/uFTivoyQL+VZNk8zo1E1XbfUAvJRCTPhbzZFm78/1im8KlJnGD9NLbJo93Fo
troCusfD8cRsb11pdBnKblIY2ngMEjKTYWpNGCrQlYzYFE4UFt7P7xggxbg/f8+t
ypJtnEe5HhWicTEwXCwc3HH+VeypZsqekQ8KUEVyY8Jt4rm0Fv+50qomvo2pb5GH
wfYmvw4gKLOoEGIUivG6hjnz1zhcS4ZPQfKmMM+JP8YYZCKkfS3dwbN1nwTTXdcf
2L5WxIOZfHc/uEuzLabnGcbj8CJkTE+GToOSDaSQTbEA2e44/3NPzHHKdXzvD9UP
OFJDJP0MRwb0hyu7Tq2jJQI1HIjD39ZP4ECLDoQhECA6lA1JpYfGbipQlC40I4tx
JZxfYNiiUdF+LlCV9hlTpvkhThZtI5BIJ3Y2Pq9m8nxzxyeGXQZSDSIZYzNAHtx1
o1hQIZ1t5mewnvqUyA6g8ktUDi1WU1ekO5hajugCiuZg2xPB8rEnCw7GYWCRv9zY
Vi8YN5W2z1ikT30jodn/TvIZ6Ngoum6i/EJhW+6YNmlQETpfs84Ov9TQ/MDuGkPG
MR/p1UmJwo8Q7YHMPVBpYSzvpSf2Jf/0KRFJ3Pry52PpI3JSTXwYrnYuDF8UVmIn
IZMiJGVeiwcLIyb/+zTGAFXmEayBh1RNZr3jwu5qnsHuYOFxnPlECl1/9asr1m3M
w0BguhjYZQ5N8NugaTHUqBpqDdg/5DHppAC7+2rr2+5XmTIv+TNHxRsrxywQ51yx
h+OLjcjk3X++FyRZqor1bzxWckuhPkUcQ/q9gzPJws904srqmEUCls0yCkGFVWjH
LR8wrGA6sY9HvD9iIDZL/ujxVKnEdyGgCaXNiZybNN14gb7kOr3R86yjZCac2+lG
Vjoomp1cMJ22Z7uEatHxCeCY3zPVg16ClUeoIDa6JyM115zRfKPrRJsuwW/mddAf
M5bBL42JQrsFQTxZ8NuvBTiKD7QDvStAZjZSWWTqdsnr/C2H7Cz8kBZpJB1CjhPx
6nrKnn+XG+nFY0wRndgLDHg/xkG8oUEMNLX1S23qE4s/MqE67GYk4g/px5KclRBQ
wxbC0cVqKSqp0unHDqhMd4WaVLmXpZBd6ovBmZq9ZmR+kF/Y3eugEpUA30uwN/hx
GyqtKlTaJ2qGrq6lYy8Ncb5ERtVAZI7qvccaSo/ytBJG0VXg70bz7/CHkZNMwwMs
RpccGyqnwNdpP2zzTfM68uETLFHtFpxOyGt7iGfdBm01Afe2hld2zcvThCRDBMHW
nqJ07zCZsFqC8RwjirZ4w46YG1QsvVoW1n84LCYu79q9TOneT4gK7A5u5qy5tJ9w
V5LPb4jvplTQ6Vbo6m8CQKlkiTcXvhomDPT/iauu3E4YQHIoIv7/vUUiARHiNdzR
GEzI4XQOfR0xzwN74L8jW7og3BRr62HivF80v71knJc+lrOkPu6d2ZTrJyzuIZ3t
pqzpTazNIp/buFvq86QpT9TvA645DEsxSiAvl9np0dGjXhHBOHY0fPvbH+/h3jf0
PM76N8w0n7AYcZ0a3DVmkB34WXY6nl0UeCY8Dfgjp6HCCUX8RRl/TtLDEiQMElSK
9FsQq5kSXqKq1lT7RZM+9aOWkYRymuFWAmTX3NMsgpUJDV5MXL6lPsdThq14iROr
eToO+480Wy7bUGokGYmgQesbWGhRgn2+QCbl2pswPxv+9On5GAfdEbbc0yQZUzd6
KD6x/4Mzl7JtlyV/ZpzZIWU64GSTa+zq7CsQnuC6zIt+AlpnXuJyDMqhubD+BNDw
0byRioh7T+gD1qpqY6CFH5L9NaynC4VVpEh4JNmUiTxxBNPxW1SuGn5jNYZxLc7T
1mCgxV42eYTnbVvHooliuFThblM+WaVBs4ZAV3+Fta9Rau03Di7Zyhm8QIZNnFlz
FcpOUtWuTqJwXSGpe0j+GnPs6daaFXxwJDmEb5cWF7q4FwypWAdvLR9bLyAm2QTX
k3m7BQhnMsMaO+zlKpJv9s5BJwz+hy7N1CVKucB3W22RZnkJsjN9g6SlHggFxyin
8s27WQ0u3BOCfnX2inFC4OMyu4QPERSL9jpzY5wVvp0P8d8yVk3FtW0tDPMqrLvf
FtedlCO4SKvYQljyajp9xfRKm+mQYgTY8Qn9sEr+4Zf+CQk1tyTZWVs514sVbU7D
w/fLWr+GYEpOzfePDbfnXLuT/9ocZuSRjHOE7/qPMRFzD+8/Rd3hfQDxhstqMUda
1TLz4XFwuEc2+j5OjWGFq5uET/HzJVoj1kBl9Y7FxmRIsETvU3RsqN3mqGD1LTJ7
Q4ML3by5Sn8vSGtUEmGynah/TpahRmz8uQAWILcFAicrB6ZonptOjCtzxIAl6B3Y
uxlRkASppavwGHnsyzvZVh1twUSssLEmx+OpEa2nUUz6MdvVrGmdwc36XPSBZzVa
JF1bJYEGh/eJegPB54m6vWkVSjLgkB2mUgvWEp60UtWVkV+fy4H0f69+nNBsO/jZ
/mGwyb6Bfs3t4ymrZ2nUFr4LgKbRBBtadFWg9DXsUUFwA5p/SR8e5wUzER+eFY8f
VhfS847l9Pj9ln5JkeXANRVl+Bob3bVDF4PMM58NMjCoVsTgkI6nXSBJzEl9JhCA
Fi+RqonSQzpOcH9dXIljWznM+j76KyhEGvuerf3+i/dTDSDSDP4WNO3HFJtljHQl
mw/R3TUVJilK6lg/dfbQm5rtSytBqi/s+qQY0qxNiVvXJrTyJx5wTviC4IIoUSZ0
N57jsikTHgGgOFNdvmFC0CYqjrh/gf8s6308rd9EKAq66dGvDUBZ6usj0u9fXbNW
BsgnBWxqpVAhst4CVNe0/lhJNLWJ0sWshejPmL6i4Mcstw0xgQqPBmWQpLwL12g7
iLNATfSxGosizlCmrfxSlmMDytUiBmnA1XCLwB3Ap+MTtlFaw2Rrc/bv8N+KwQ5T
Bk6aEvD/RfROrYn2aQqKMZw39vXzdY+CWfr6md1WyauTlLR9iJnvkjkHjPiFmz67
kieK7pkQGFjZljixA0h/CUpdwSxI/6wvudHzcr96XGKV2uVYlbfTXJwxlltheha8
vmuytAtBgaGFss+uXntdN5iWtl2KQyAEiQ9N46DqbnwE75xUNFtqOI5nnnQ1vVZ3
smhlI77LBnxpuTLJEQXUgV6KIEfUkW04zSOw1+hd8/JSfDXyZ0aOBTlcOzwJ4eMK
lEFJxLzQNr+YGFMn7x9yZTYCeBZ2xrF8fHLNLhJ32/Tlh3d659jMa40OcKvHlPlI
M/p85+zICvg9nKSkJuIad4Qsm6HMBHqk7Bv5onaPC6zBzTdx88oAtejWeXI9SWZv
Y8pGsvbNGdMG/8ZQD2fx8bkDgId7iPQR/XPfSK7plC+dE9Uu95GekRrtSCHJ4Ft9
0+qnmk/U+SlMi/8klJuNRKBeYVSI9wAdlz2tnId1Ji8b9leJ7siiI6mu8nT1dIVR
YKPDxbjG4Pp5cs+av3LBNc7ywaJD8BqksYditRxA9ik2+WFjfSX2yWbtq0Bd6Ug0
1r8EVcST1BgQegpROw7pXjHjX5w9qQpI4FO8dUtm9OPbQ2vQIJmK+028g4JiY9Ff
20cP9JMr2Di5z08AHS9GpJWq2ySCVfqDHGDEg/JZLfQdiypbtKXP7GAAEz38OYeB
PdI0rDOFbNLNu8XImEutNtkTkp4DPxcIDgeJNz4U7uvDqTWrHcYgfRBJYL4WCKd5
jS6CE862+uqTThHtBS3mVaLmBYnz8l9ECCQf5UpZqqEIJsQ/u/jKEjVfmqbgnmDa
2NHwteju5AaeJ1fTq/oUn6eVk40eoDEuVv3NjIwLfIF7Qtll1y//lN0neOt401rt
OxuP387LpFQ8f+wTDCGGCKpNEb7mUUYXWOlQmyZ6D4jw8P66eOrAPnuJtztaNuJF
kBCLlCI6YF2M0aNrEIyi/xm6Ux+PG/n1B2/WfwCPOUTwclkduMWpwF8zFPiqP/Ql
cjSa4krMco/pg1PbDV5Vj0o+VwmfYzs18vTpK4DlQrxg2FbUYesO7b4rKhzQPBcR
wrwJxIraSl6Cj7tgez0nXhPd61wwv8/VqQqT6b7D42XCn/TcYzkVw+RwkXekpQtF
vFBy4MMm2FEdcA0zpe4F0cWJ4Te/bD2S/uKObcdz6hUXtmrRbIf1SAMi2+60s5I6
/mYliIuwVs51/XsmzH89Ql8/o/DJaj08Rn3qhTczn2lGXy2T1G5hxS7Vll5XVP+x
6Mcfz3hudwYJzRnMQ8zHK1dtzz/Z5f1yTpXriPP/mE/cttg20Kswt2ordr8l9fcH
E/33cGrIHhskD0dc+E2F27wiLqPqClNdPkXDLi0zbNlbT9u7A7skR9TeBDeXAiaL
jQxeQ6TAugQcKYVSsmauz4VVv2G17x5tnTymfjDVyBLXU0EXnqJVR7d5Ntg15YZC
LwiThB2tgM74g+s1OCA+MpUV4m6FPI7dv23QZl8CGvLIDDaBfUBfYy1qQNiV0Cmz
Y3d+85/t3o8eVh9bL+Ot4ygTQE8g8Si9KewwH/r3ydexZMrrfYOMufvbZV2yBJs/
wxqfVOxmFwzFrFhvJeLCvT1SiTXUwzD6NjWE4f0kOwNevGIIoCGs51IFvuafEzF5
FYuYaYJwYAOjGYO0VeJtL/WLZ2gO/a6lSd33sHiM9XuRM2OZXlDSimOGD+eKqQX4
fzY/fiaunLf89G/rvl65XMuM94V1RxQKViziH+mx47cN7zYNtuvSy7+jzCmE09Yr
hI1pkjqBSusVujX/DuQxz32WxMBxA3YmA71z70W/6o1r11jLYMzYBROWGI7D1zge
Q5zN8gcArgpHlvX8yfZi1P20hkCMK10Yb8n8/NYiFrC4ZElXThOjXIxlYX2CJuZG
aP+Fy5dVCxqhaFEcLKSDmllREHMSwb5bmExd55n46/sZNLyIhfJOxVU7o3/qbyHZ
ZMM+DuUHJRT/xByUCPyH+EgzddaYXJrjfSwZZ3BxtdTck6NLZv8bMCz05e3JZALZ
alSnO1J2rnZWjBUu9ObBEGTdRSRIvADnNrtu9x6k1e02d2b8kVzsZzQ6Z0Uu892o
j1hWbHkgOgnv1LuT1kcIMDO7ls84Gs0XK6oW+tSS4aB+oPmzihQ8VYz8GVhb/L3y
k8m92NJtfHKOGKzG8xMIVnw1E7QcjWHAqoIYvv99cd3REydODAhFrfeieXL6UkGY
ldtlqcHw6feyYh6T1YywldC8ujujhSUTL3f0xwez9w5LvQAkYRbE2zQ0uFW89mOH
kAoaRxvpSijW37uiE1+TOjnb1aPsXxijsCnS5jSvXlrzIwbMgTFaofazopYKpKS1
zkhgNyQ1po87uPZgVi8H+KIdA9D56viNTISRlkzMJgilznp7XJeWvao6+Q0IKgQr
dmTmcUYTM+EP2RFgrHuAnd35IbhEESo3+TN+NoBpgjXg21PkTdUQH0F7xredshNr
ixlfpLzrKtr4m94pGSKWo3mkHBQanfwFn6dATgdKkIb+sB1wTfJylNcJbZmuUOh0
x7gx140CnL3MuSpO+ODnDbIX2SMfrrGK4JUlVSfv54+9JDgWc/1BXiGj1TZV8Nw3
ya8kUnXe/yDP8qmUPAo6IRDdbDu94hPcmWg+vg3M4PIkoVjrZpzUjbxIvJ54P/It
GsAXNWzllb3ebmDfVQ+gUK0qWxBKe1lHeFhxoT7UErmo9F5kBvSt85QzstaWg5uw
NiW4O/6HN937euMHA3owL3hjRQYaDe0286SNu8CKcp3WLTKH1e3Pbn/Arp1zzg6u
jsdUbTZW43RnTbYvUFDSsMXB+1og0tCnEuToe9Dct7XZolCegJh4xUldVv6ZSi01
DWFhJZoLggqpLxTCZKEFjZRqkYu1p6kT+y+f7Wc689Byvx7VPM3qT/lUD6CzHNDV
l20h2u8UFRj47cdNU+1HUB3IE+MhCchLEdZF/LM24F2qrugQA8qRV4MCyKiULDuN
83xwmLHQR1uReIYbdUToNjaDKcjLe+BTTQESR3fLrObhqemJZKXcC2iZFIoEM+cb
/wT86nwZSVWkNnHRdX/S0Dl0YuwWfZheXBLs/OuVGaCKa0ehe+rQ0kDEsZkeWVSw
aBwcsGAw6AqmKQB7y6KFMAsoOzk0RrpZS51yETSy4v0ara894ErYEU9fYt/Xy5ra
M0tzuFFDt0UlB7CZOPs3a0MeiVjpq3MflLvMfzT1C+Cr1scNMoVD2TaSp/UxfipE
Fvi1HdmPHrxcm7ns9luos3MOxx1hijf51SBcbpgI22bVy0YUA1faiPn4JtDLGN5B
9i2AXhL5r5oq4Qb3F2jLOBd9ihDUumte9BA+pApbvfH9AjMpVv9hNqQP2M4m4mbE
kJL/CS3qFzahTnfrTCL2txBgVVdEEWkKAKMVNSonCdJWHnSTGxkJkg4wzNr02+rj
EnYJSpS7VlL2YfoA8QjxPHoAddk7IDa5HtVtw9vbmzun6Mr+V3FRLSM1ZsPTKVLF
1IkQlxBfJoosaCxYet7U5IYXaNBDw95IOshvx95osbgRIVAK/IX1OO8cUKM2A3Sr
pP5ZSEKQI+/Tee11Nloh/Sf5mAEfc+km/mAs+6K5RKBeWi7fwEcja/9/i0pvI1t8
fCNGInbLQXHnbwCzskFteDXUpli86fxDT6YjsptJIiN4l3vmIxAONZV7gyTfjTtN
wdyFDpgIn3QZrblrU2NTrP8AD5375ihLeyQPVQ+lWb2miETzJL8aze7WlMqwWXnl
TCX9ge4YOx3IhG8jY+VDv1xwFdwu+8eZHVJ0FF9OfMuQUdin5CnQmeFeDk7N01oa
Uxk8B++D/FbmhYemyjgcNqmqrF/upH7HeW4MtsLX3F5CPXLaNI2BL0NBYPhSgUzy
Pk9rI4IuhjSXH7/NK/paauOM/i7wmkx5rOL45xAm47lD9V31+0pt5L+1OyP9f903
ADPCD1Olf4fgo9BbY8SBlFoHFFAK8KZDOi3LvI2mChFkj6rAYScVae73TK7Kcr2E
qBdSZIU2OUjJwI7wRmzVfchFqVRhrJ3knLo8zFyltY6oZxytvNh7n+ydGjK/lYzW
ALahPNWEWbOYWeLmCUanixjNIjf7T9TOhXRVNktVOHltFPTpOY4kWnIoLxvDot8U
WEZOxsbQO5slkqrqKIvbuXrLr4DCaq4ivyS0PSuMiXzm7BltCBw8IjQ/LuT4QDzL
jbtcEzWgFS2gT8CVSm3PqZkFLV5CnyFKgzQ+6iSUnFzcgan/PLn5dkbnlwa09nED
wYaUDhRaQ4upTFqnulGUNIflelMdeU/sYxutNqdNF8p9Ut5xFYQ71M2VT60Ej/Nm
9E8TE6nvSa7kiVVC1Qz2r3ILOFej97k+saVGth7bwb9cDIF7LEALGMqsGAjCBSru
7dM1UJhv1IYt7loqsKIUNnaPR8H2BWrYkUKEACi9E9mMA5Lh7va/UZHtBO79m7za
mw3u7mvVlIEcN0B+elndNEFXBhhvLWyNF/9Bb1oGyeVC0pwIOCqzMSfcDYnk6+eU
uUZm/j5SNhZsGtrVnkXovE2itxv2WewC+1Agc/IsHhx0lhS/YyhFPIoaTcY3LFtq
uUJsqPhyD2GcsED14NX41jJoQtGFp/LGvy6fY50JeqQ78P3wHKiMRXQP9sp2Xp5t
GxrLvl7kCA9NbyqfGFV0XNZ1dS8KxjNGQr7/O9s9eYcDPv+jfKPlBJb+Xm7lvjxB
KD0GcAM+uyEltM0gP7VIekVq9a1Z/e6g2LGw8Oiq6tdxJDgdOGACBPDKO3CI11lJ
GmuSVEAMYidRcD183fCLtgtrJPnBcTdEwlBDWRk9CBjNJvTP9TmSpjky3cHztMuK
bW7AZCL+lRvsP+c0sUGR491iqjHjkLWFdBC+9xQhTmWxItOWgJbV5vriPglUGNZo
b6Umspf98alZJF3QWQTqoYY42NHJTS4CLcYbtD05AYt4qF2P2Iui7vsbaAFQ/XCF
bNqOjbUi0g7wUAx71xKDoF8oFx/vTSYAk2rnKIp4eAQ0/4g/eDnEpYix8RIv6p5h
7P16LVStE/EsbLJgB3OUR4t3Gb5qrNYnb9G/UZpIlcNGC9/zHkoEz4+mYiksnQjl
qVVdbf1PC9RGncDMsdn/Y7f5GTs2th26qtjNbsRKMS4hWMop7gjFPMDo27SpuM6z
KunuodsBh0DMgCZ6rikbnkN7pU2UHGw7xWw1x8CbtN6+pQMnr/SVo/FT8m3Wy6Wk
eFqYVKl30f/acDgRlno5xSZAM1Rp1H80pvqcDzVHCWoMUVmL1K7NXZOsnTRNiejq
vnOGr48uZfBq3f940bMkbaIR7gi4G27+E8VWUrFqOqV1lQwtgbs/F5XCQX/BRaxX
SHGb5sOHNb0Dhsb1EFpt/C5jWL5rXdMf8f9bxf+7kGRGbRmeHkV+9nKELj0qceVG
tmp31xxS0MaAMJ7GHiE4gnwXIYTVQ6p+hYMk0pKzecXvJ5PnicAdp9q9Q8SUbmsJ
FH0BpWFh5lAiid0qNuKpZ6XZenD82fAbR8XntE3Vksn/80o7BN7T0Og3b5TSGzJw
VBnTIwVwU8qSCGMD0rB60baAqCOgPe8D1YWyD/VGHd1jfbjKxArXkYzEHsYGEfjt
zN0CQBl5SHXlWZljvyjBnTlhA5rdQ+qedcHoYgwRdke9gTsABnpSv4x8v6+haiQq
gf9mUAouxF3pm6w8QEA4y9D+NNKqqegJvmsYirz5ykyPwpVqSMXIwivPM4gSMpWK
AhKATpeq0KBZJyG5SNypEzGwfeZ+rTzD/Mm3ev/FFgbW5Fyz1UZs1UQALLNdwTzS
ksTICQNnW1wnqM51SLAbNjizkJXDphbw0rUeEEVXzuibG5090FtvQbdRdWjV7C1o
MO/n5EiaLKfkMqeYj6tewUlEYJ79OAf6aYBj2J7vTsnKVrsJeXto7oJrDFdLK+V2
SBH6TyJUJzzrb3fXXgXkcKo8UXU4Vuue1CGGmpnmQmL7SqizUCqn+xDgmugHyWHj
pG8HXq1CoseLQK/gh40uphT8dZExeSDUUQfhKCeHaJv/VOn5nTpuuNlE8FoLzkp2
CrNgxoKsrdRxs7L5oL8qqKG71yEZUfKbOERJdf4UfaGho/LiHyFft/G4ykcftMie
7k2fjdm96NiCec/PzMZEJddnPxg/l1lqZiiAW+ycIlvxhr19tIEsAD9Aoa6VAFfX
H5FIM5w8DlC1M42625kHtjE32+PA1P98GgV9fG4K1cBYxuSUZDbl2fOpzw3wJthW
WHYpxxsK6/ql0e6Rh8EJm9funYzQyS7hyPJrnUVHzfaYJHdCFmOzykNd3uJ2crDF
lU++tsxQlcLnjpcoiSeYXmoYdnRZGjrYnVLX9R7MYXj6Hy8WacAy3QbWB5yqs4su
HPaKBfcvi7pvXkcUGBUOt1BfkJs5oEdGnRrs8/h8p6pSo56h3iJW3gyreyPtI6fW
OfkN1hIHXUN3/r6htaSCF7NXjR1TTBDjVEtmmYek8pgxsU8lwf+Px5Xulo9kJ0T/
IaVB79kMNTp+yfChcapF1QWhXMzzbFjyVu22QxpFBaLjON7ifCbY1cwmMpOxngoD
IOv5s0toKDFsHWNxI/4Td9v8GikbF5kd3OL0rM4ZG+CdX4X9EQbPI3e5vIVqNXvk
JZIdaXV9ROhhfPDBuCsmI+xalYTWvVqBFjTiloiCcQ+u/MJjH1OMON7welJl2MJl
mImv7cd3yJRD1r8vj2SFaIk6Ak//RNMug/Yg5isbM6KAbImsl1CRf1Ro/zJXXPtG
PkAocJITEanc/+vDt5n44RTc2xqH374+m05gFDyGe0u78X3eZzqAXwhKCljJZgWl
DyscH1f4MAr+1cv5Lz6jy3Knqey8scvencMMVqmWNQbttiQuD5snRyd910483LVl
5b3RWJ6B6tJGZ9YSZ0BpjeKKYROaZB4ERpjV4AQzPGC7u9v3EaKwgIMZpKv721V1
0RDC0qwvlo632FumWCDV8z8XvL/QjwY9WHONGp2UtozrpjPL6OiXZGcS9uhpI+Bv
wacOvu6Xq71AK4HH7Qs/I427hgTPXL1dd970hrMTf1Y4gcekE/Ey0uCDE2MiQt/K
a17FE8WUfdlKON8FIIocEGq13/St8JunvSWUWjSVkU5H3aED3ynQNNmelfbG+IC7
/WM0z03bdbbMbXCu7lgGVvKRLCCohKIrHO+IaPtcLkYWgezv8z2H+a1EEONDfZfm
px2HtoXn4QnD8djot9YaDQCfFsd7TvOsiyIXYfbK1RQAY3B5UqI8u1aUfvF4q9vn
IwH0ZZPNsV33RoPcZP6ytGhXjwPOWfqnapWio5aHYnpsUTBmNziNudlsUmZvRogq
myRnr7p7cBJUVntj703+p5w7MCcs2/QPma0iEy7Zxqrklv1k2Kkjn7btUpJCqzVk
5jQ8HbtaooEqPEj36beOLhkQqnmrX9OQJaEIhizZ4JAzsIl4fCmeYVe2YfMM2rZ9
SICzVxjdeYlKH9mrJPykS5+h1EX6KDz0y+ykH2xiyn1VWtGcd9Q7h5tgJ86uN7++
tSLANGa0JeBjYHzuWuwpB7YyGXOEcHjUtDxaxPyC9Feyw+dHgQ+89SIKfELikmyz
6d1HHxQDaj7yCWm/w8OOrliSaoMjAdmzPTNJwjCaLMh4UNLiF8PxjvjCJuUETSY5
kMNnnb+QcSZVos65FERzidGLfaQka/0+mtM7PUGA8xWYQYqtOry4rV3kaS/Rta0D
N8nk0PUv16vFYv4PKjo2TfvlvOOIDF4+tgURUzxqyGjUsSphXY+fi+CHiJu6Mxvv
n+XwxipkM9s2FK5OrIkH5eA6GQvIPvAbo2q2hqaLcOjYc8S6yJY9qaHfcXkB9OtC
7q1CaghPYWEBnG6KImetfNyCGrcTJnmvdoYBTv9Trjl2ZXEAnQsXBAsPoa2GoezU
UweM8bm4tOKMMjXyLvAbIQcbL8p9ly85Mn8fy2/eZzXqK9V6V6QR0VOyD0rvRCEe
xf3BxjKzUzmcJE0GRkYmWa8rWjcRXWAtAyxvUDf62a6yYm90fHiLptqKehBmHDoG
Zjn1oXdFnz0iApsMTIU33wyNxb2XYzX8oeh0YZPS8u8HwpRJktGTf5UNSwzh/p0t
s4TYQIANPNbF7O1Mbud+qKht4JhIrNVAJPW69rO6VJz5kRO1SuqRQ9fZWUDnUhpX
+8ZmX0NA1dAJHOjQaXKAHlRFeivYihCE0DkdJq/GNzyp8Nj7Z+OHddEiFscxwY74
+HPysMl+9zVj2AbSy90lLOKEQSEdo13Si4uEkSPnEvUfz7qWG+DIv4jfC5rGoqDG
G4bfE2rcQRVjr8AMRl2XLpzX/ZjGPWoI3Juc7RR1m6t9ntgwCQsBKug4spNqu8vU
hrNJNLf1o8V5gjxyS/ssI2wEoGf22AfC1rtqPXwsehhf8876BaMYpiV7CDjPOhWY
H8YoHRrk5wOf5x2gkxJv56EBHTOzGm6SRiS5P1GSgo/st22IRuWWt/ZsNCkSqVHm
G+6oNYGLY8h7EbtCkCsXtmZYZWTb6F2Q1DMOZJdwmV+1Abw2OohvHxWD5r33bNX2
BPkcrUsgseovJFM+2h6I9/n+8JsIuaud09YI0//hdUg8elpMWkozC1k7Ki7mYXES
L3fXr60MsxF7q4xKM+QBdKXnOHP6skC45G5xMWIGpXmh8JV9ktTdc36m8IHOGzEG
0xIFKNtBKAqKC0NrWnLLEhHQBt7xqTtTGvr6x9cvQLZyirOE7r69GzBGRRcZ9ke8
ZavFwnDbtr20w/VanQfL0cgRnIbuDQStvMtGPZ7sUKJeJpzsKeRTlSu343r68eym
Xz5uCErMkrrIK5rBIbFqLX4CevXcVvtdrM+Aq5Gd8yK6MOHc5YIuKFn/w/r2wqRs
PXSLKVNnBvyIx1FUli+K9G5+Cd1HXyVB+kBxdQpG+/gelgqlmymuamHC4KiUUXv6
UVk/pBVKaUuog955QlGan4SKx1lUM4QZqya6k6tarxZG6YSgEvDxLjD6chY5HVTG
r9aKFTB95Zd6JkhFIm5rH/u6sDbTXhGU3xTp/qEBA1SDC8SOWuJ0bohL6/E0EQNU
RhxbMVh3aqDPQeBaitfPRBKEUQjCHpv/4Eza1adNE7XFXr3wxm3LpBePUoJiA6UZ
bOg5fxhtsZxdPzYLc9XGgomCBH8V0ym4T5VA5/hWgwQonUGoWpehjCEMzJhDmeS3
IHHHeGJC39pGy77ApztN9ms3sjxKtdCKlLlWxPSnThrPb0lgBaesSfSjl2lVRAgk
sk7X/jUWBAJzNiaAkzcPoQxRf+2hnLXV5QkbAmfbYf/YdkXFF3gZxWtmAIq1WZRI
U1BtwaKfX8nSMCRV9zBxqfUzykLVdkthFVlxjKadiUFud/I7Tahg17DQBbX46YAi
p/VVcflfJPaYVeZJjxKpnpT31B8O0MUvZ72l+efJHJ5nZ5+vnDZb/x4P5Pc+VDFn
kr9yZOnjQhhVbP+YRY8Z1mTRVGygf9/dREyWcmS7wfCmL1br+qlhOeHvyLtMdt4O
Z6LrE9GY2QC570lMIwvTHABjo4Y2upTz22gMS0MGO0TEM1RfoChB0+JAMUBgz5NN
3M9Drr4+3tFqVGmpBaIsrb+abgDR4koXPoVQUTzELsnkh9oyGnICBLCvm4U5ceFz
JxkB5ZLOUTfO0PSOXv6Gc6kJSRSpCZ7ktPwZJ+L0RJaevwyvNaYhdrWtKrcjVVbZ
5FMHsPMO2cdTNjNR4goebfdlm4R6pZWJXSo3Ct7clQjHlerU5UE8fzoR72mXiEKw
rjUTB1CPgGdDkpvZ7mTz4f3L2GSHvkXe0lmmRDLvamW8Ns/E2q7UqAaKJ1zCdSEK
ZmWKwmEODiTYKuOqdp9ZzsAZNgyE5oplAyZKV+nSHUgi5zbtSsiRi6vkncJyZN2H
lvGbWjbNX5hkEusf8ERJbrHYbD4fooCcZ75urH/ybLPT2De32GlCB0d/auqxiFtv
PmSrdkkwDXZp9a2uMtEd6BcUGqWHmze3vLyIBiWQT08x43FiCaZGpTBKJxoAD7Vo
x3MtY0NNwT0IcU7RhGZsnPCn/1agX14bse0FPNPpB99jiM4dmdkDQK0cexeg9etl
SZieZu6x7A/ZYwOf2e+7/Vz+YdzSJU8398DNdg0Jl70j0EPpC9Jh8eB/IDL+BcY/
AtJ7zfrjLYJpDSV/7yooymvgwKgcENdDQ9Raejw+yu2LWipqU4PTNSyPD9NylXSV
Yx6HRVQgQOiLEZpe8XHzCyW19LwosnLsWrEuqghoHQpIN04OI22B9g99DMK7I3s7
M8SdzW5gvwLUbVnr+uWnEnfYwKA0FsUIT0BD/pV38eRUIt0UoMkv6sNecZuhoM0U
vpipX1OL73+/CNWFpzSzysCYG1ffvdezZal1SD39aNZfZIfVYtsZKA0e94E5m774
ZUCcgWFDnBU2lBkSihMnUIFefoZYJwbtOmQ/rceOVTB5WhPQZKFYV6P7vggdWIZE
4O8EAze8XAY9REVJYl+pq0rx0B92mXd4RJFPkQwlWch7mBkh5+OrG+iaqmzZe8YI
B493E2NLdLgR3Dve4hHLtsOLD0JtRQ/pZ+ezaWteTQx8IwCNRJlYuUbhCpF2JN+Z
71G9VKzAgJ9jgJw+72FNnFMr8o/A4vPtJKWUUzp+o/RMKrm54YZfPQT6VRFVW4HP
uzXgEDKKHqBwOkf2a4PSilIXMNKMhdhLtUWxrcX7E0gCD+xVz2JzYh1pRQhanM9x
Bd8ur1YtUWu8eX0QpNvBoR2D6j71zkotTax8lKoAiYBL4Tu8OHMQeb5wBVA6eW96
+LTO1ag+rA7YQ9q7nW28m82VKHmK/p3+6T7yHzI5smXi2kZv3Che74adP1PzGB/G
FasW/AnoNaTRwoOnLZhrDt6PwC+iqJA8pfPGG3fJJNT8qyOeFx4Shpsh5S4lFH5k
eFwTQGUeqf5oW6laZB576hx/Xe7Kog5BRTb3PlFApJFR8b7xTq11gUthUnoEyW1K
90hLNtClxNyxjzhMwTXpAA/1u0gFIY0q+SZl72TeXcCKXAGZzCtR1fUJtt8Z+PZI
AGiknfnWD7KPbLF2Wm3Q9wdxEYJosIVD8E9bv5EtgaAvHr5QShT3GxJo4x0aWjAP
/wbGIwW9nMPdMeuNwS6qKRGpdw+NU7WwYd13ehBSLO5fswD2LEqOaRgIQC7p6MOQ
N89QqttepBQqQht3caU01uFsxX1hXUkAJbBw9mCAAVzga8YhFwkD28WmDHqkf4SQ
DXByMBmEsXrh31i420B8b+SIJt3lo4Z8nt7dCvVs9T/gMlVh/qiE53hWtN6OMGDc
wq0tVnNXThp29OBCAgpQnDImqGfxW8S/izNtGqSdAX6Vn0hxHcyf2QKBfMaftNHx
A0/R8stsc4WmyNCLIWUHDb7S38QfhNZzElDFKJJXayzRYSvEYno5B6YCXi/WPZZb
Q7Adx61a3DyVroCHggy8xi6pEKSDzS/Gi94x1lbamROCwpYgu4Ar0hjzbjczdKLf
5smJ7DS27cj/rTFj5NRdPUtBfJnB42adQB4/oP6625dRUp1/vwD1GdAU8NHtZU/p
Xdm6/Bpji0rp1sGJ3rSPEH/XiJdh0qhupXAQ0w4pGT7sjA533l7AFeyini2NgDeC
akKxXs9Zeotzzq2poRr17BCzjTRyVY4BlE0dX9HCyOUo3yG5bHFoxMiXHF5GYYKA
PR7c8FlS4ldYjIyOdAkdYTzzEsbTzR8H0DsfFaDnxn4KtdUtBZOxxz7ULlsdIHqs
712Yt1G/kmlYqFZnTY6YK44Wx/KpcJpHMN/rKkKIBKM/szbgJ8a3ArTx/kFhtAHu
tH2vePx1ENJ/5OLWxcOu4ZVx/ENVLNFi2l1NCpGGOpHHuFApAdSeq7m4h4fJ9RsV
BcnKzI4O8PYy2wl6QuWCTnL+yWPwvkV4WqvwXYU5bTSTOWXZV+5TDp4qvkXsRP6b
a32HlVZX4NU+hzxrXfC6usEDMjg+5u5Ys0ZHDwRZ8bZxmuOUK0Qebf2DFSdAp7vN
XZOeDlAsGPmBNRQlZSMfnvYFRKqDC6JQF40BdOpY+XEbV7BgKIh4jDvxqh3L2qm4
IdFkUOGX0ymiVw08ha96Gh2bX3S+1A7fz3qqLNJ/NfcwGZAwgq+8Ooyba3hP9vI2
lhOAdQy1A5zo+urIGgNmm3aZqd2B5suzr7brFW9NCjc2auhcNuP3wKWKQ9TmmV8S
6rYYux1hbf28atGWm+y5LWmDZpmi97uZwuODbmRwlY4sPX8lrbR8f5U6lL4NmhgD
DjsUURUP5ykpLoSHag6W2R415uDKm+VsUfZef6esPe5DVDIM7lf3+Or+bpyEHG4a
SJnpVvK+30MJ/wIyPwTIGnuRwz8n3mtGtrT8UUaSIMGdGFLMtwlAf98RK4nh7vMC
s6mH0OaxFdsOfIaeXyreO9lv6rIG5XfXm6uhPcFC5erwQn8pvNtd7dxXNx61tCN7
7mawq7EPrWunIx07e4pQPqrQK6kBOra00B7C5g6aJGamTeDPB25dxkslRwVaEvgi
WCeZyxASz/tOfSMRAmSuLgXzsv9RLt1J6fwj/8PdtOBmHfDz++qtSA0Shc5ZwZ02
I7pihSNXQKNg61s2QnMHKM8dABI9qvTGHPQoP6WbBlLRyRYGZg4NpjqK/FMwdEwl
8Bvzsr8XpZvIQzAvfkN/j993J9VCRrcpvDFNe3Cp/zleK5TP7uRgKchfJa1vVVoY
JEdatJquU/+6vBcM6pZwadOrZZZyiDrqRd8MF5NcRzPNfvytpvJa/tYUb3O60yGl
Zn4W5TV/Go80ob11Uq2yDC+r0rCYyA+3lcw43IdtasHIYFOc1XGqQiSWs6JAitOL
/cEvZsgH6NgIseoqI6wanqbY30MvyaXAV7GIBFwWp1VfWAXEeLViTg1MB8qkxTYP
Bao6N3i76yj3wYSivYcZyv+dMiKP9ontKiUzGzVmu+CCWtymJlhj4db6UnkeTDWr
h6WXlYD3TkAj9zcSuGhWQFgQViRthniajPOuYURr7yXwEvzND7sbEj1OhRk0HnhQ
Q6Z8xMYctSWQcmlEB15CDS2iFaNULU+lzlKChmvI5FmnDaPlsLgkQWrJZWYqkqA/
hfKRv6rAiuZPYb5YWzAS4exZ32VH25aCzYM7hBZkCiE0LNpdmW+h+WWtL/g/tuQ6
keFKK3DonF5iOdZH6/Y1JsJupDyz+hAKIk9s7OuYbXMwduUqXYoQljIVeNFoh5hz
X4ASWLc+s+bYaloSP32brSUPbcSgo0moinVxNkGLv1T3hUbdaH38dIuXF5o18INH
EVx2UxL4dMt/NRSmdON4m7x4TVWL2YPb91gqFXOmF8anXEPcrZC9G0LknaHRlZf6
0/yaAsOZ0y9X3dlvXBcaSxZBlF18U9KH5q6EkiF2fBprrJT13fmTYHo2uRI3FkvF
Cz9EA99BYV1uyNq7drgO9LrEuCbQiC/XdXJijp4zunmb/pAvcTcZ4gYCoztLaarc
nB8IzKFRPeCJnC7I05/AhwudsLfSLtknE1j7nKZmT4PO2YPhIUSc8dQi1OUKjNmI
X31zah9rN21EUVINvIml2yIPFOzR2uen13aloCAJ06c34ap0eucFCNMIXwKTyBv6
GM9McIWWIXxjZKTzYVa4n2CyI5UNGeNtdflMN4Cm7c7eCE47gr6qJx4vtgWYCPQs
X7Uuwfh+rnTKlFdtpl7/Zoiwq08CMcpsMWLGwmfMn1p5WRtXfi30AJuDejXZ1ZIZ
p1u4xQHAKzKsbrqL40tAvhgo9LFOnG9djY6MsVirf1ctbP/n/vSo91sreEtf2hkw
5FoU9ArqUUdc1QyLx234LfbCFchWNkouE/NJATDj1FdRm5iCBZcn5CO0Sl9XYYce
0UmyQrEk4sEvQlUEJMuNEGn/W4ptj2KyB+z0rl/TA+20cU/0byiQ7UC3empzrrZL
Ar2o4BevEDCqaI5wJE5eMaTyvWTLNVW7YvoHKpCNVxtKulDt/EMHZ2x9tdRPvq9d
LwADpDlbrTuzO+mIwQ5oJyAcuPT5ArofK8k2B1fHfOAHCU27YOQLLuFfpQQtX12M
14AbNh5+jE86UnMkJHTW0G83PHQk6zj+nUZ53k8HIm2ssvvZayOW17bXycxVbUMq
q5IypWaVwNWjdp3DZLncy4TgwrN+oO7Lcd1RXYA8Xywz3j+MEJDGLktqHMEDMafZ
JPAvWYMjqY0LQyYN26WwBAdEXAaLuCMry/OrBfm/Z5xWQgrB9+wCj7xWwt8NeBHD
uqyujnfy9AiMRnfDIUl2a5PkEx84Glk0rq9LpXH626ZZ5YY4zwR6owe94i49pZrG
ChewZw6AKvu9KAkuYEV9TzHoQ1kwB0SHJrLg6bARSOT03Vn1wyDGZI2HUBND9C6a
C0piYEaXDBWjRjPqbv+wGQYe8x+3Kul0PBalqK4O7SXFBeTACVN4tlEOGmMk5+/i
0xroboXozA3MCDnz6XeatxtdP0ri6jusnCTah/tgZuv3a2oFXdwJiHd0BUEQzuAl
/+ooZgEwT4OkLzoK/+r/hoYNzsWT+YKUri1QEs1aasOXQebCOqBtnH1mWEmdcI0/
TAxgEfcQLp66CoubS+6zwG7RZvuJR3Z2qjQF9OP86XytQZZeMK8ejDFri/3aO2UD
mBW0G9Bxj0LC4z9ZE0CZo6bnV7+qZ3UMLYgh0/EgkREBi+V92SmTG0bdvP+l6h0S
fxAt7vQPAfNH2FoO57QXJ4lmrws1weO9u4CR0t2JuYPWvXoil6p5aqKoz+KsohEI
mz1YbtaWi8f+ZC4eNY3ywyDUmL1OCo/Z7QBRnM83aJBNfYXXdEifz6fR8gXNkgL7
bds0UOZ40WATX386AB8S7NAns0E8v76a58Na9YVbhfqt5QfyQeZ4YkEPM6iOQ1Ql
GBLfummjK8H3qogQwP8+EJo8GClik0rLfcYXB2362uInkwo6LnN5Z4By8qHlQedw
DMgt+Is/zc3beyBxIw/eGa/l/VSyqVZuM4m09s8wvbTvBMXJQoAviKZb2nLfgMej
CNqijU4nNLgVYMiFgxd+9C0OaYXZSQTOM9LydNxf3XAy49V2fpKZGAExVCSiAt/l
YGO5TYeCyB36Nr91T211KuxPV7zGlUalOVMY/Ug3nqbCiAk1zon+VhqJ7dDik1QQ
hq6upg3V2dG7V3tPNRaE/iY3o+gIDTzYdmd/mghAAT32acOq3UQ3OPeq6yIH2gKb
W0uhtov6BvH6bBAHpHSaf+53oYgm5CikC+cPi8fnAYOMwdmxp727BoFm/mYKWfeC
pfP/a7S1fmo28wMafkvRFnsCjZgNvKNCr45UIqpPwCXa8tk3RjpXP5OquLBfsTJC
sbhx0Dbx7rg6WQn1APQrFeVxXvl61jUbX4kTf1JzZLBIN/b02b3VpWF0Mf5x7DOq
MisCnQst8Ts0UXOBZRj9pqCL2yVJhM7G99W/xisguamCgtxx3O3IIqn2Lqp7qLx3
ghN+VUaqo5OwuePQl1YswH27Fbw5fTfJVZf4RjrOlnuy3A0Bt8Y+SKwVceV4NPHg
4FvJ+0A4LVHEAHFD7GjLvUwsD2EMDMVDXgnlx9LXUgvELZmvlQAej+6PgxnM5EzF
2ZV8mCgdKiuLhCGNPNLFGBFseHkkDLhTZ1IEJycDkAea1Clr8VJR2cD9Fits+rNL
/6ysYX3xxankLcRtMKX1OABiAP6ETRxWAKM+VyG5u4EEj3oHzE0ZFYHNCpI7k1Md
7dhBs7LU4mL3I6rFFZDVuy4SRYgq9YcPeuJ2KiijJmHKpHGulKFmZ0rm0yGces9N
QFYoAHJZr9lp4WS00ydk+OizXgn3+fEP0HDyKNjpqbMcygin+TD6tM4ZQKb4LH3n
HeBy5b+vyYnzkyPmb0+/6gEH/gwVCKGqc8fu6fi3yG9tUAugEqkp1w+AviDBw04p
RHpN8cYEPAw0HFitzeYBha0CowoVqfNvwm+epbC+Eb7qW0nMXJXjCTSuqqpv5M05
pKfWW1ipP+JYEZ/xtXeWPDmmTlGstmnVhUDIfR57SQSmo1+hPw3Hu4SvJ/x7YBQn
cNy/KHIOSyQuAWsTpakcBYA+W5F7MqFsYp5VkyqFWpZoBp+7d8p2NMhfrY7zse4T
Mw3bBRGRaoYVCz5bP2hNYhRLGO6o+Wqpocvw1JEwwZLxbOinNxfeIzgIIN9BQvDX
tB/W8lGhXsSSutJyM6d7hGPKHA3LFNpBjDz+Qx3+U54Li5gNv97Kgj7EtlU6BZCn
orpxWeyV5rAa1aOpUA8vI2Ao3XkXSSVyj9MPeioLCK7WHHF00limVoCdoihVZDQt
1QufEIHFrE8kqK0yBvqL913ThlLrAxHeNSVCy7lf7tpBX1AnAv1lB+NTmPt8PbvD
Sz31cauVDx4UL/30kcm/HyV763qc3yn4IeWY/gU6ADmNh/xqu5Z8TOUMO43hV+Rx
xSEBexTCzryB2MHec7L4xy+EcD5ufiILGkKJZ7eGmK9WyMxF4Ux1b0vPN+8pS/b6
jHNFCgHv6yZ+OES1wv9SPxOJrJTvjFEJFRddYOEKRH20fCsZJZaIxMrKQj6hXFmK
iggdi4/1LTHuCtbhLdH51IDaw+Wvb9oXnDBLzRD4KSiSFajh45gP00z9NZz2QgzF
QGbydqdI3TnJSAh+ORX+URcCIwW33GLMVRsFFHiPZSY25V3Ryi6rH+kK3B4KbcJK
3AwANRyDKEjAKBhg6TEo6TfFD28oZTejFlZuky+roRK1OkYUZY7KYBtvMQFD+qyd
OTulPFn20hMy2IB4uj6OAgwkTfLD/liJI6fOsAHDNX1OBsQF0YtOysFmZh0b+tmF
ysSC3scOJeEgcBkWWQOqBv3Y5RG+is/KoWbJMkzVYJfmuwncikQaoZ1LZgmkDDvj
+bnNf+kQk3KjrTHD71CLu4BdvljEQyuSttVSG4nsa8M7/L3U1AzwWLSWXewtuKpz
kP1xFWwdOOBAcCQZ07utYEQLllNCzsP0lBT0p44rHiVzHlB+3p3rDO3ITnF13eyC
/YNWxAdGeE7uBEmNecFB2yEfexkBgmzSLk5sQrfMq+snNHIl48/B35HMUcjptRIl
KoD0tvVPhKVUSyfuaHPip7/H3QKNiwSXVBpwNqkitzUBl9iG5nOjraD3dRkBnVbD
m8iA6/TQeYUl+NT4pa0Fvxc6uZUXhCuyHVndm3NTgNk0IVYgy1TCguU+2Hih+gu2
kXuneRku6XaQr9LaRVqwj9eZbpkTIUTnsiYve3qDdxYiPL0e5VdRsxm9a1gS2G+n
5JZrRFhwz1YWcIFz/ASgv092I/qtVJa/QvhPihh2g7i2nmc96gtf9FrkTa5153cC
Vl49/lCg6163G4Li+2thBSk/+avvCoP/8VP078k7libSvEgjr/NwzVvE1oQwe1Kl
jroCY7Kdkmzf2lt5c8uAMfDOgpTcbhvs0yNVE04CuUDF9GWKpvBuddfeO8DKZmmF
XAEDm0XWui5i47VYuPm+QrvlDuThXhnge1JOwO5gsChVF37NYS86qhZFQSxpJ8g9
LHrUCFCyMuHiP1RIEMAW+QjtCEonrnHzNWrmjeoOAR2vbegZmMAXF4dW8kqKAkXp
8+n9k1oTnkO/d2CtaWpNm6gd3LXCkfyekCach/8eMFR2DB9q5n3Zm5FD6I94p83a
4ioqE5BZkQoNKCn4OQfM0c9aG1/JES9jIwEogBtzFMpVztMgIY5yTuSBWNoHXKTS
kQ2eM184GG7bhNFbtYTVmszV0uw/MCdFBGoeT8rbt9jLvNGpPUL1LBLUUrUjIXWa
DseodCqObtQj5LT3nXdHTrf3JiJQNsqqdrwNnfDL52srqkeAzrx/ArqeY/LpO00R
LmnY0juuFWZvbhHXGpYa6hcObAYGOc4sC7SWqCcARQMrcVML+6nXvGFP4S9/GkAW
x9H2D+z7taQ9UVaAEm9VGcTS19NqE7/OD/D+clLxCz8FqHeuOYDAGxOim9JGVb6Y
2P5JlCyzxjHGDhtWEO9YEbC/rUGyxyCtil7+0FNjbBCDoJn0UioK5QPaX8dKPZbQ
zAugz++f2nk2K+xRSAmaLtJwDsJw1KiuoZmCDpfu/IMUXE/lgEJ/AESgIa/mUqi4
tMgFnfB4RjLtsLnUfx+Uilk87udcSqKP7xhA6JqT/+dNEIcgUKpRbACOLB90Im0j
ZaxVGm0+7OYnkaXHdWzUAvLNEATA7LCpt6Tg1lMIHEg7m6YZiB2+g1UaiPs7z82Q
wnZquOvqJ20OKmVrqsZLashsuzF4HAvH6ym6Mjg7SKzEbEJ0nGq+P6AXmOyIIuHd
SVhS9t3zU+cqhUf6o4Rz5+p+ylS5bnj3l1vhiB35RDjAVNyfkmG/FXu3gO9bpCyC
sHpmGBkjY5cYDmxJ8yjLPjTR74jk/tMo7OHTJXYQi+Alh23owNhkADbUmN1JqQ6P
86gKiUqvUkPyTMdO59g2HURXgwD2QHkn0W6xjbcRHnSUWkG2uhk/k6mOx2da0gEZ
bhwuB8+JQ0XJNTHhtgBqW1z8u0WOA/JtlxBPKW9RbBALaPm3Vqx7ToSReS31nOSU
nzfxrjXlp4PcDVOpdXa/mTtw7qyX+MEiOHucyk2f5TmSlx8vQjta8nUBfXhVeRIx
I3tnS6GPcHUnBs54sdqGy/ILFMoNF32eBYpEo/bFPFXFJ3wy+dgnxIFdcFBuityw
+Q/N6UrxIe6kCqtP9TRai+F+CdY1YJ8zA911JQENxH0X/2vSRD6Jxr+TiWA6E5Po
qVPe7MA06IRulD+9oh+tPlNuE1eDbNki50h+Ndr6D0fTHT+gbZzKOdIIRLqGpJew
RNKUuKkTAAHMuZeRchxQ+67JMAE0/oQHqRQsz4WVLoSHy7h5VXeoVJGLUifgt7Xk
fGAsUFiGQ9yvlGq57Rot3HfPu6hXnVuR2QzQ+SDbXtpx8NdHNZUSZ8qPhUKKe7l+
rbgBlwwVk39BVPrWiH6edR9RQ/pb+Hl4JdUf1DvaMey/mmqvszd+paqKldGn2RMD
nR2qwrbty6Q37hR91E8RamMP4LmBDYeekLB71grfP2eK1GRyu8557bxhrJ3meUIV
rAeA+2pprwwzzT5AdAjZu3vjE8BXo3LR9rajrL2RbHjC6hYgjf+RdmG/UPTUlx22
05aeqtfPv5EovWxrHqKYWMPvz2FS/BrPbtRQFsv6BiMXrOj7YWVszFl/4vinEsfb
f1AjlHlemP365wHXMLu6Ep0XUf06YaN17W3eKuckDceLe+negawCKMsN8o3fwRtv
c0Ms3zQwnG/HK65o1Z+TsPBHf2jjKxR5HC1TD9RbEV9yDY6HmJSKRyNZo0oshznn
EUIIYii0dWUA2tu1DU6uYuFzfT0f1O4Vec43abYVUg+CCKCfAJ5OfqYVsLuaJTfo
i5bttPP+mVTzHluCAgNi31JSlxHiPR3xt1E0k2iKn/OvC0X16/U2SFCKcHvolPwz
LNrD1/+u6TAXOOju8WFw83lswjGJklZgB+bcr5X6V7KGIQlIN7bS3HS91+A0RQ5i
snaVKGhlOQy6+GRLQbeUW5BEg7WSc9NLWVq+B7DVSWS/3dLkjqtnY2pMri8Dfc7x
nAAlp1pwIw1D+QTNP7EWxXlOpVtT0jjzVR8DUQ+3r+ugZoXjjh2L9acIi3g9uGM7
M/mlAadkstTu5BfLpMFaQzhE1B1AbY4ZZ5LyHXGRlJAwr7euvUposFIly2WQg/SY
XIlFVuyDxeG758agUQedopHaWI8pO5klZOCv2SzIG8JYRH1ufDBvLdaARsVEi+tb
lUVSS/VRgWeO2fNcm8jjP9wdvsttaulrzfG8nWFjVeiTPrmTopO/7/xBqB3nrE1X
ofeoEIoz4MQScoAeKWZS8x6lwOvOZzvaqozF6b3+xY0NpO+1yzS36YUnryhZl0Ym
gY2tItJkUctYc3O/0qS5XjIPlG5bz8nDX5anZ1Y8oubF21s2Cn1WzWDxr/nk5AJn
mihP2lQ/qoKB5KINw9m2h158hxhSeMHqAzPlt9Ymo5te6Y/3np0iEeNVxyqREaMX
bLbpxbhKeU7Wu6WVdeMeF5pG6y85I4lXQBV/09zGUYh25jh+10Xr7advbGdFZLs6
ICWt6rHisJn59oapkBtTOwfPgn58VNnxCKLsILFsx8+ttkg1DuvhGAfPDdV6D21W
Gk4AkT195WmnRiWJ7Zy4/Q6QARcSWt7tsiMeQxnzWjqB8jnsVJvs7t5iRZQeGOLR
qMjoNf2oU5F+3pfNrK3ayP1C20FfvRyPPSqlSJoR6A01OhNSgz2QXqeOIajWYA40
Su/JtZSo/2tjjtcbqlwgYIDZw6AT2wzVc31zHcTVccY1/4xjChR2AWV9B4Y6AaXC
+OuhkmZQRMXvbllE0JVPB9rDj03z+W3GXx4E4xzibuiKXy6IoW2sXsqhGRzIFwf5
sDsUnfrjYxCpQRtRGoBMogLdBvxgzgBpV3YV1/Nly/UgAWuN7QToojl9mwuzbfSA
UAsEku8nLALHFRHmirIY52toU7PTZWoz28uphT13TSJD3Mu5cGVQ7Ky9jSY3VKMK
8zrlyxxXXiduTyHBSInWvC3EgLq4Tl0yYp7bJi7r46eqv8s/0XiQbPwLjt9/bRFm
GyHbbZH0iTUcEkGe4Kh08eWrlblCyqkMj5+UsGyxdLWVLDVCrY6W6hMf1Fx1u8nu
ulx0bSpb8FskjOeWQFMBuM9l8xuTVZNgCNQ5R8jOXgoDeGVuZf5EAUVDjiBAYBWh
YOR7q+wiJblu8frn0QFyxNpLgdNrGhJQU68SZKl5ELwidZsQb9pXZba0vu38MB7m
atryBKruVKxspX1gSwebxb8NfLIR2k897nBwRROA9byFsjhrRWcmVICgk4J6NvDE
cqYDPYR3C6/bNHTTJrt7+SZeV2O9QVK6nDjYEUvVE+zoO5LUu2UfZfo/xj+9dT4N
K6DABetAhkWQZVjKpEzHmBYV0bzBvUxi7bYA6XgAiZDqC/heiMY32tJ+Av1II1ZR
qaDr2J0baOEcfk8bBNN7MqFLcTv8tkVmF456N8rIRK8jqARXRqoq9nvq0ZuirNSp
UO8B08fuAJgn7zCaaHvKAVzuaT8C2gwfqhDhR2liZcTp/tFM3rvpPQqXpnJPAwZE
BRDNJQVms/VdgQKjQpEWnp687urJRNrZvh4jcGQsfIq7TZmfAzRUTCZ76kn1lfdi
EWhEgCz+ZwW9L3ONMZNlqmNm9FCt3OkqGGGCgT4KtKo4n+AC2aObVlkp3U85PloX
j1UF7/v1o7JXuzecISMcnRG2iyyWiEmf0T7ACqnsadpW/RmEBFP8kVDn0e11Y9ax
CxpB4phUFbrArDJP040eNg6j+aAJQrx0L+BrTgigxM+NNPOR014oDdem6Bmq0Op8
0GFGMcjI/F/YrpTJVuGA/UrE/nBkWyEzajI/iMNW5yreeJVLeE7FmIWa8b7UJqX6
WqpNM6Q4Lyl6PwZgzRPOhLfCnVJ8HrWwn6gU3/0VDdvBYOjJ8UHRhh3xPDBmM0jq
bbjkaYYG8J7opIaiga2dsOLE4VrQ7YEM2uktR5di36WKylcNWRkWEX8Bsts/LM6Z
5rhRhVXkQduT1mdjiMGBf9kldPp8bP9mP0m6EHyn2HRIFD5nNKFhEPuiWgOwp5t4
CfcQl6LbF8WoyOQWf1jWhsXsQZOrxlkekHzyWbRnrllZJ42fRXfHy2FbPiRbUAVu
QdvDs1r7upVQvgHoM0/U0gSJQ6jFyggnPskkFQifrsP1Uhjrxe3awrFD82krBvHo
jxdvgtPsEQfyEnNzrrYANMrJiwqaLTHGnEKwXZKJMJnxU6VzVsaht6/2Jiig2i+o
NG4Jy6qb+ZGcWFEWJ2eK/SH558aXceBltCTRZ+70uR8E84eD+M1mgqLDafr81A7L
z4fRu/YD1AnI3QQ9vvEX0fZWS254DysfFm1LkFJSQ5IA9tRfBX6bzx3rGtjg9iB5
NheAuUIiosnlj9ZAiK72WbR6pzJAaDmT8jVpvh1UNVpeMDFtbmpeFBYZyihuULqw
xH7SwFzP2EzNPoukCeKr9wkeG0a+2GOaYyH65wICKyrkXIKgQsGKJgrhhOEvuI2A
fzenXBJOI78wLT+uWyIJ00BqGN1Wzwu57VVxORllsikRk9NnUGwTm0S9K1bj9DH3
AuCxVhDa9tMnmjjPI2HUlWSAtikLfpm1bVV4fx+I6Ms4UdksizArJc7MRG+K5zJi
55YEz+irR/7QinA5ogrSoJ2jVKfbbTWDL7U1RPjfURD0GtcMKBk1dtHndxnCNyTn
j9BTGujnq76GugMC3jGHqFo3v1vS5bwTyEjwgtxf/nA6qHFACy3WNAqYjfr5wMWj
haNDZy7w9XCDzIhzI1zropg9CeU5SqGrN2ARc1z8qCSKxirLgiWyqXFSgTZCAgE9
uxrKtjDtXyhsaZ4rtzPe2OYOSWuvSiWZ7kGOQhaZaq89gVQLY29G/WvE6iqJ9F5q
aEe9Q5pkecbOMmjzOzoIi6Yw7PhxgqUwfMWpkTI1xHDLvtJdQ9i9yYhg8s5h71Yd
kQeB5ux01tgwUXCcoRbmyfChqhAY7qivJuF8LZkWAPTaSOZ8Gd0uEW2rMpWgnxow
lT/eazDrjPctadOvNxlAQ7dxSJVBfYDGgb81+ilIDrOpxg4f2zsSPXsGxh44izNs
SNjfykNZ6STNP0qMtX0+zfRfBe76Cjeft3/FrF7ZJQRFtuSmcmvcfMfX9hlC47SJ
Gt5Jk3Wx+bGjDuWfROl5PHrn2+DwDv88dEJDy39E/B32OEHFkMmn/Nue5Sag7v76
QhDfcGduhLkDPt7ExnTQhKfyWmKhbhtooIDdh7uGJOsTIgfWBPNbxJq/IocjZw3U
/d+LZstnemA+r++7xWgdEuNSdj8wW12FlRd2uhupXl081whHM8BLeFDZgVtfFjBc
MnMtJ3e9+CnOTjfCBj5T9Pan0YuFxkVOf8B/7PBVNvgu1IaMGsAqcBtd7nQ4aFvk
gwbtPxzLR3/6biYXRsKJEvunHD/tAOo9Wkp32RcKTe+dG4pq4uBBIqlXr9S6uWPW
PlKvnAZnDDeeE7eyZb62MKJM1W9AJbEnk6CnyKecDtFUkBRyZvdCVhCNaO9V9bAB
+j0PNN4m/JVU0ADEno4+b+zMrSibGBQup7ttNY48+//wxsSqzgrcuZx6s7RGjSE1
SPtgMqBKRimUKggZtdvUnoGBy508pr4KoAAL1roXngrEpyPJ/T184P4jnO7Ivx81
mHgMSiE/ZS9U5yzmk2HtJ8NiM/jYKiDBd0wJgmaVDeVilHxAv9HTBayCUWTTSbWC
188LVFEzQdGNEkM/RlI34UczRUDc8twXagQncysouJrpoLK2i3vxqcs/iXUDN9GH
JqnyEeNHXY1qi15D1+K1Cn5lYrVBZsSRgZBDhiiH+JCouYiLICrkH8w36gYXD5Kz
W1dlyT4CFIFVIfSWs6slg+310dq4lKZyvIst5qBqwB/70oD8vFAe5cjCaT6IXd/C
9YBWTCCfqCCqLYwVpDjctPU5BLkUtauFkGlp64Lw5jL+9FRYs3lWl/v0L4ANhD5g
s2Qw6db2rvKGTpB0cvTMPeFP7V4gUg+4L2B33dHLao5xLZ46su9vGeZD0yFqv2eu
/Tz3oWRKIKNKMmFdVb5VG+26BdXv2kWiCpWOk7zCmns54lnUEvNgzX2czPb8DdOq
IAGydvpVdofuXpHAj6fbXbz0pX2PY6Jqw4o2AdlNOqd16jU5E8p/3/6ImpGyrx5r
hDlgSkWw6KYSqgzt3l+EOHfQ0TUN/TQ8G5ptYC4ZKE6B2wVWi9Kr1kA4kew480T0
ChuXZUD4zEgOkzv+Td4qTalcG/ngB1GbxpnfBAzv8EQJezets8QTBTrO5l5M9NG0
Svd4hw3QeK2+iXngNIRiYO7972AFIafzhWKr1DnUM2EgOR4wo//JHKArYsa8/KAn
Qj9GkLiFf7QfkXoH37EI/HhqCJOcO3S1KncYSx7wt3n/M1ScMqtweEn5xd2GORKI
nqP512GEDtWLUclp2+oUJw2n4qulC8NC4s0QZxr5+Ecn8sbl3qZsv7P5eoMyEXSb
+Mm4Al/X/Lgj8/WRXU/1Tn9ZnyyutzctyQyDmRDZ2L5YUKLPhCK6GDe8btkhCvUB
moGyx3I4LLGDj5wwaIJTiqPGYvXRXA/JCPXAWWsjfxNvgbk9o/RV+VWv+I1iFm+l
S5oyqZwLoTX1LOtWX4HUVHlG/AtZv4NzBVCOyK3mxRdLjSFCPNKDFzG5RyOJzN9M
FRiUqMzqB2J9LB6ttR84BLWT806+35nlp9pWfpA3NHK68zL09msXKfROpQEgMzFP
UUJSz1m048mr6y8O0tBXooN+xAXGzHyoZF64wn44lFncifP0A6FUZJBLVD7INQkV
lkmtZdoRzRCwjT+fT+i6vprDmXDYWMFx9FEwJyvZP4fEqyOoAkxwivBO/I/13ZI+
L5yykgfklyFA+8qeZ79b5Fj2F74bITaqxpjJHCg8673+WGqX2Acq5UrZx2KZQHLT
rvSREtIvLmtzMNe+4opkMrqJVPMRBrmzjeGHPMYUqGWyIMl9m4uhHxoSFTL/5icf
Iv0JMy6U9jhsJ9BHnDv4E8/sSrr1AnXWKNahywMQzxUSMX5emFn4frRg3Ss92IVC
mSpv1Tehoiw57q66qqgTK90Q5evTpnSieVVetoOr1AcIZI4nVa1Kf1LKyRaNzi5u
8CXJbnMpWNAoBC80oKZEvzQ84O/8c41U1u4msFbvtONb4seU/phmgn65M2DAe9hJ
OtqpLz95BCg6BcUve9vZNf0F9vmVlx7nMfMNyQDTvlc/QTXY4HHeKkJ8dRMG0AN+
nQPXJGjsHLomwB06doFE+hRk6FalpILKCj7pGoTk+VU1+PwRxnPpGNOGiQuGy/Nj
gM4/33tlD0bW6YaLYL3Yac120DqaFYgWVEw38lMxoMnmxJH60U4XvV84yHxw6RQD
hsrBFFh2OwQGvUg9lpW5kvVWEwLn+v8vKaOCBjVbJel22u2T7gctHrmuelc2LOI3
yA/MvjUr1X8eF/O9ABWfaQBz6Aue8MBYByvibI/mv+oXZtTTxybzh1ObWW9r8aIR
PlDScleMIsjGVVWGnDzENdpBmcjoDVBFh9Aw/X3kB2al/A5lP+iQ2IGRaYt/8hUs
LPdAwXCU8gdDSM9ZDCXVt0ljb572PMryVq/M/KnCCwHQyjXsDlJk5uj9fQoj7geN
6pmR+XmpYquapFZaqKWxmLH1F6Sb9dNhXk5GEijGDgtC124fkWSNn1ravbcSErlH
nyHCQ2hzNOkJWxlXNbqorz52ySePWpnyLON61yygoJbYG28tj2UNiqTIabwr/71C
JIkhTmpgVDf30icjINcogKipPZZrt19S/8SW96gq4HfcNUKMZOuYRXisPYqQOIh6
H3mAdGoW/EFBm/cxqLm7ScKGVrMGMwRqUf+1oPrMFKJNyvBTyxHf3HL6VpJASQ4K
oqK1mdbm5+F14W3/0ZZn8rXqQRXrgWtnxIrjKRCHsErJnDMpW0T/fdXb+FVndkCY
k/Ta0ug1VydqXqlqIBAqWTSMQGUw7jdmyszygoGz/NeMnKTpgxd8jYp3tiXc+X6I
mPLU/BCwAJoTqBau+gpjhOauV/O5g3vOFyRRL1NsTGINHKP4ZvtKG9dvRPAVDx+i
zUOCiIQ80kT3FuI+zI9Z3L1fUJ4z6m7jLIVItsxjnwl3Gu8Is8SzaMszdOicTNNW
aVsTKH0AZnAIbY6uXZHuhYnxrmhAMzc0zEPKg3pDi5Y1HuCQ8bis/YwXEMTnZA4r
T2giulgYnQsPZFgenMDPyMy7a1TO8IxGHca/SdjeZTdQiCwvTS+caiV9v3YA5hPj
84aMNET7qzI2BJaoz2QTpdxZjbDy5W6I7Ec5MFO/LHaAsdqlm7Nx2EutsLCshL66
LPDhMvg4fGgYYMpE+tGRj3omOnyjrX+AE5A3StVopdbumfnDb+4i4J3D5co8yRfp
PrwhTWOmSUh6SViQCS+UxQJG6qCnwUpSfnfnfmKtfvGUziQ6UFCHX8lbF1USytHy
S16rflKJrbZ2V/LiJ/ezVpEdEACvt10ik8yU/gi628RxDUIuP1Kq6NHU9wCm/JJh
mtzFbl3uEFoD5d64zvGXnL7L5x6YP//qT8mgg/GFyMlHy0rs+AwS+EFeqWtlFfln
qK0cY5ZkCZtz1P+3rEYcXt+QU3tAQhZqJnjCqQZIP2qy0xembnKsnpVYIbOvI1HF
B15MsbyzzzQL1zBQ/IRa19QrZkFmYzt2IdUsZeI34oT8+m0aQ8CQrGUiy0uQBTiu
8u0qwu4Im4QhlDiNH1C7jPIMQpuEjBVNfg/7nShex1qymPzsTpJMnzTKM5URlD9W
tUV6gg/xnR1IioNZ5J1MpMnYMRJ5wf8zoWtUaV6KL1uX/N5KWmZXQPXfztzvRa7o
Sw279fatuKxGwbNDlHD4e9QHTTedpUdFrvvolxJqRHjm4XjKmnkGcBlNiaoSYVvM
Fk7fV85K8X0nX3Uurk9Yrc1sJM1W6LOhvRNb6hCTnivFy/bKecDdj5zNcAGO2rJV
PAh3mVkWi8Ev0taqgTvBK2f43g4v6eDG1UHl6YgIVAj6weC4ERnvgmPWFU0CSSu/
n6lE27VVfIEsOYR7cux4Ai+mq4rraMyxt0XKYadsbzM9JuMpmIIIkqW2oA4T8iAL
mDOd6U5YrpqZDRmND20Wys2lC30iWgXNolMIUQIvWAlIPAjZsLjp9APQmah9vWS1
IvjDdzE36Jahr1i0KNV5JvMjnsbb/3Pjng4kkofXvHC5HGCFz5dJxjTtLfSKyBsI
12A7D2KsKjARbak3f2huejZIIsGBfHiTdUBTlIF1Pg7gXkLK+xe2ctmoovfD8WVf
iYDQSCkGQEw0qLpgJxK41s/izBCnAE/a6lRG07S2+6ND1koCFEgyEd2iNAcSP8Mg
RoYU+5PEonBgMlzTL1/Xpl97S6D8jNz52e7Bij+0tSLYab4uuiHrfZBEHhvx9Zgb
oUBgn9y8YnUkmz58Dh2pUU1/uLsEZzaQ/8mzUuKzmM8WEXy6i/y8MynEu6TwI723
D9w/qsRzRzrloPvuZA2V1lH5tJxOih4MsNDxA/udfGG2nl7SH+fEjGe7gcSC0IIB
LHIEJ8DsLE6VSCLJrLfxq8x4YaabBeLRddXYkR1ZC4ao7GG6qWN4EVNSs7PsFWEk
rXAQmD4AMD568Chf1A2ojmfRawR+uUqyfsg+M2gPD0oWevCRUOhSw7d6RESbVeqT
L9rciGg/K+ymzJNVdIE/OiWcioDfKtZ19t5Oq4h7T2TDOISgBXwHdXgs8Mp4bspo
dhdwu+hBaG873TUxfizbKhJ2ubKCKfDzYf5A//M1oy0P4qNbkXmEhbuZvR/Mgiop
zmMxr4TUwwHiif+b8VdAGpB61QNmgSoTHcTIlnweXPHk10h5MT5kaQlDwPRF8Z/V
z4++dtbIkdR/jp1qO6B43fWHqw+DoXHsIF0ivD5//TZJSWcKmob5EOYZ98gxZ4xh
fHz5poEd6fSzHhLdDYVUgATZLa3qXWsfmXa+jaxvGNqCBYhcqNBVYRd6n08pnpKZ
k03evaYnQd0OPfPuMaYSrShcDB5gQrSM3MDxs4Y+Duqi48JSFpiirKk+77XW1lEp
ryW+4kg7gdZ/YWYlixdVOIcCGtpvhYJ/nwE/nuNI3ZRde0UDU476IKwSRc9gOPg2
O4gO8gmC6H73/oP0bMGqv7Y3Sc15GkRe+LBmmxg6xNqoyb706EngZvNF89ri2+Kz
rM0KcMOQzIFZPbFdDALyNz+7+FG43Xce4eJ7+HJWjBjeD5fcQU6Sb32OBSWPT/0Y
pVZ5fVKuQG+QfiedjvdCWrL5qKUvrTOjmMxY0PsRw0A+31GnUsr6qGZ2q+K0Gm8R
fiAZqv4zTbplGA2ww05a5ly0B3uekXagQrdLeIYjSpVUKw1R6ozizZYfKiBkStM8
isEV0pa+F69AKgReSDTNJhZccO9V7E0iCOXWlt6wxbh7ANof1QxwpRQlNkPcwMih
FnQ66iJ8GGN+KEo2U9YWxIbGLgNgFibQ+cQWXWkvRL4J2TmLOySpcllYX0eyEEvm
fm2oGbqM9/e62oaF/RI1MkVi8x91KnNsIXkbtILGIt3s2n1Yd5ToobJvu2u1IKLn
RWyMcBKQa6yC9cgBux70vP5YVXkao3ahHZBx6L0+1pXe5vnEHB6puxinOp8h4Mkd
y+81QPB2dAX9+m5Pg78JptLM4mGXz/CVWqmCbTnwhlqd8eVOmgiExYqqk6EBt0D3
PZPc4zoBOCzCt27+JYRdHe9L9VM/McqmRTZYpxXIn7Y81jw3RrYYonxCmSyg//aZ
U3vg8ReT1ZwxGyR3OHjy1Gl+S4qoJ7nXazO5q2Vm8GGxmKHaN9PwUwkOXMLcdxkX
NbvcHjJdz9mJwH44yzT441LLjDEoioGbBvlSo1jV8rMJgvnjxVx2Y8E/+MkBoerv
QfIv013GJBeag+9Y8sW9VuOZasbj6MsEZHQpGdzM9DrM6MXJC+TLAhz9ITFh3vbP
D9veBEXPU4jxyzcbJes/7H7yS+6q6ijYfzTL61/BC+Yih8bHFs1FoZBhlOnX+P2D
gzgiUTLPmgZ2qDE4Ly4f0sJpcmtqJ7JsFOjE1WxeGWgousDe6EQd8S+VREXAOVr6
XfgIq6WPj5xLxpiXiWioz+nAC9Wr2h8GQXxQrq+7486//v7UaFAOGLbWyzGyF5Ef
wBwIqmO+FmgfBYfXkUsQ4CuSmxCDj3mxKHRL0Bgcy+r1L1R29zQ7KmaU53jRvu2a
ZyndUq3BpzJhnQ7DosjChQx2TtQrxOZWDEXfq8O32lLilCCarWs7EgPS+TmcJqUb
hP9LcNzJGRLYtXblVSFEFOjlCvUvYquJ3piMM3s6xtOmcH9B5vd35xazuwV1Ebbd
FFMnO0exEJHMGIjMMzNrH/77AqLjw7aGZzoE4Ve6JnfAnMYM66pdqLGhZVEbOJhb
uorwn87Qd+d+5WTgOzTqL17ythXkaK9SukMRXozulwYpazvvC1CeRr098JFqig5F
9gViWfdBhzUtzSS8ilyxlrk5re7ruX6jmjkKNih5RGTcu3wntSO93WA2ZHKgDE41
lFUWXKRcJI9TzGS1FvBrJOkHQgUWVdeEk2wtytKOR/wef67dRdQwGNQ1Iqsaah/6
iTQRPH1uKWjmRedTRFHst6bmRFivVZmgYfjwwEapBXeLYsHL54CIdb3aHR5wM902
nY4dZJJi3vgOc94Ogvgb1bIAxwpXg3H04SSS4ogKCPKsGdEFl1so+qOOkN1zGwKI
BDqU+3oRYIQOO/CBnxzn1hx8C/VHG0StLzwRfiTAHkp/igDx38c95URUFQjI1c72
TgpL8khFnNAtSBPKSE/dPvJuPbjFKSZ/5ABPHi14ALvelzn6tMNpSTXdewagdicJ
re2eWV9Ki/CbSB4iOf0aoXJcnJMH2g/rXd62TvT/txK1AxBWtnQPcneq2sIXmGaz
Hpt/AmmtSwloYSdptCn5Uan6dnC6WurlhvYafb1MDDTHSLpUYunULIhpK7h8etMQ
ZHEme24n9ylIcMpZaSdRwBSd+RVgiBgcBK7GUHBSqofjzElkn7USB16VZPObl4gf
joxqdtFlRE3kZPb9XMCmXsWWSt440sHmpH2hOr5clnJv23yz6+2IncZHq3++CibW
dwY/uEq1ysxi48eeRMBw23kFXJkYRP/kZ83GQVAvuQQeOFGvftBOUgshcs7XObku
mRlpEbJ9yEElVE7J8q35savsCpMES1BqB5navQwAoFhCEBaLnoh72nrN8q8wHOdR
54SW7XEfK4qE9MAeP7nWKexOXcVOCAuqPNhGXUbSPNspStAPiPkyqpsXRtYblWOI
IJ8znpSUomSMsouUWPtwNgjLkQ6s3e159KlVYYLtDt+wauy6/+X6OSzA81rEyIyJ
jKVuwzhnVFFdrmUh9dGsH45XGo4f+8PQiK1IDog2Tts/Rp4wujvVCZp6djXT3MJr
KlxbZO1ArtfG3FWZGCybspJLNavpv/CM9u6q0s94FoTHW8HekNIDtrPlayPR89bH
wsH45h5BUhlZV92o191EtsAl0BJUZ1I4veU4RbXhlfjuRY9E4eTozHg3Kp4tszDW
cd8lrIbEp6zbn7cTrGvNaiCCkHGIoBAO2+RL1uqt9hUcnIoTia2BApoMZ/bfFHUE
jpH9BSaYtha/VWH3jszfn3xXoI8f3MxPKJE6v7UofnPpfUIAVZ0wQETVTFO8AjdT
gmZY7R2MxdcFvw4EhjJlKA8/3BYuOCNc42Qqqss6doDDrIEBSsNrdO1UzxWp0lb1
dNlceeTUlLW3No9D0LUIOay+zuge9OA62AsXfUu01l8VniuOycnv2VC3z7aJZ+Yq
IjnBM/qckLZztIqlNyu+UWWTfHNJyCH+GFG0sNl846qmgylCKnOkOY9yLy6Ht53F
euxWWNx/mlE0zNq5UKto3nlwcxjYdfThwLrGq/TdH085Ng5qh4CXxQoLVtaAtYHq
It0RfdI99mUmqdkJuGRFVHPbUTbAr4j3/AjuHiR4fMI6w9Oq9N/CDuSfpJN5Q0yK
O5XHijngN9rmw8nTPY7zWQt0rgqdRD4yROZY1VdfTPuPbYLxj4cnDKqE8cUAp25/
ANMaOR3CfqyxNUR7NcbTvNFKVD7mAVqc6NVU0GVxtodDDr5bKwm50TncV7AEkF/J
ELxUKpY9a+z12z5HhV2rb7Wm8PgLoNUfV8DjbFytJA2jGwN6+ojtp7DfkP0kCPwq
V62XA2nYqiWcZXNBjDGZAm8P1hbJaIhJwAtCPzlxROVOQR8kslAuabzvlftA5mbz
jwRspgn17GXqloOjIOqvt/rox+TgL2ihW5hQL4+3WVk3JlnqOdjlEVgmSwGYYj8e
lkn0xtE0kLzw6que6Nfy1ormerjkn5fxeg+xRHqySFrfsIB8BNb5MPYfK/BgnUUY
YgbKy4w7Mw5/1G9WOtIsIaDZikYQ63nuoIzHLsB/Sn6FL4MO4NmToecFPceLOK0J
/hieDfW+nh3hzErf8u3RaW8WpmQjt/jT61y1hl2ZwzEyDmXajNKGIVoYS4bH8mIW
KACBpTnVfX9pu+rD26sRCs+HkXynTJX4OP+DmgGcjpT1M8/uTBtv7LBUIHajYpS8
j0lBfDd7qNXOiSQcQuOq4BdaJfxdEVO1ndq5xdNk8sVhmAzLIpZaUFFzY+WFg6rI
isyOqnrlYkHB9m4ol2w/RmwSJW3CbRI3R2UaVavtlTfmyJB9uInxmYxem/OKinPG
5XSjjsz6zZkjQXdT89jFO6bFrVbq3FonMR5ZY80WCR+x799DQ8potPXVaJ48qCCn
anwL9K3DkbqZNnyT8dvQGvRakBnS2qklQFiaG2UfohnYV5XA1SMfOcJ25derT65C
zgR6AjixLNsf/qjgmcgKwpZ+bsPrqREq8BQEMLULIrzr2FotJmkofTxT1sZyxKsh
4eIUFXyKNHnHyRjJjX6zTSQ++KoqoBS93kY0P/5Y8j7uLdDDdcMoFWjLSXGVTZbT
F7CL5jCnDj00TYsPKEmsH5vV9K001f/FWdx4P3fRMnyw7DFxAsminyO63Q/lxqfO
TU0QiUkq3myLb7UAXhhGxy3q2uVKVEknIgprw386A+w3/JcPMQJBEFaU5XGdDDdC
vNVnzCqIUWfZzidAMTNx2bok/CnXb3x9HT6NmvbNELqDEYTK/uzj2eQ7CljPoyiE
xIazSbUKgKi2Nm4ZAFBm+bOWL1knXIAlonba8kOj/5qQDTQFWUv1kzO6D62/DYhW
o6T2SlVJ+GAqGjzp1JMVJjI4Yna2mZCPt8+1toCMlRAx+mIvJVvCqziz0hcBa4Vo
uyeR+gVKvMo1XhifVScvScBtmV1pVoU/2NTfsGJ/weQ9RahzjdNUdTDw0+bAklDQ
QgVPp6am29GKogbnjRt6i8fhxzvenxCrNrQOVmMOakddQWZn1D4AUP/JDJ/kGJtV
KITeXoBxcYxOn+pkb84V1hvtzLNFjoHT9oUYVgnZEo40LlXaeD4OSSAJ8ZTlxIG9
9xFSOkU8ltLUWBC5QsY1+fwb87+BxkLDQgSPLSaSQk/r6sLR8TOyQx9qyIfs5mT0
KV6i1sUd9uWkOyBo2+ljxLRONDbRnRqkUyhdm0Kzs24Vjz9AGr2DheL6FD7JFHH0
NzoCzTmQ5oRMVp98ev70UHMHogYRRBL+66iC6bnir9aY6j9F7S6sRWHOHEhaC15C
aWqdDyfnRNtVu4cdy7/v1UGyuRDV9egNtCRy7KRQcHl2pXdLV1tlvIsGIhv12Sty
+P6FOdi2FUgvm6DNGVuhdVd9/pIVPLSf6kYl/S2aza29xyvADMOM7SURIdh2/1gA
rWbgT3ZTDuONk/syVbc5Z0nRf6ZypqPNRTRVNwP80CC3iL9aosxP6FFdSyzRHuxn
TUCInrTQvnxUR+7ojkLTFyEhc0IY9dh03rYFEnA5rUtUVrf5rzjei7kt4Bi/lPTl
NxjqptENRTSzTd9TqGUsnAvEqU3C9EBRIErqT1FLhLAtv6VdqGCty9JXQhv9mEgM
ZWUVHrFF9Es0HJyRr3LWGkBakTVxu9IfQpzPkyuDktmSrIaHiTTXOPMCsFP7h8v4
Zb2hshDYYr+uj5LL4mSiCf9FEMbHLVVo4i2nyQbIij73Rp5gZrzZ1HTQ/s8hnxKL
YBhVuSRVif6DNQHUKAPcaBBQwAo3enM3FKh+1If4WBMuBUGc+5DDX3uLP+427M7w
8q6+uZYRmvvNcecHeSMD+cdBzPM9I9h8H62QLaQrXc1EcfE/+RwSMEUzutKmSF13
FpLjDU6lXa5BFeVFW+CbpS8ie3KSfCMscPU7LuWy5HvELnFEW8jjbZYT5mQ95Nmb
fSOJKlWKrx96w+1qGSXfmtfBdrjx6/K4WPzAHIOW8FDs+fE23baSeymem3+TwkzL
PbQFJUJmsIlRYdSaeDeyrd3JOwdyWtVNkW6fYpmN4+FqgwHv2Zab5hqNSQkmmz64
f9KXAeZc2HooSPTs5MCYhc9VafAbtO3e0blTnwdXJO/tej0gqCKfdiCR3YJNXtw1
YILBYNCGY/xN9B90C3u9lOhbeNpnzAswnA2u6nWQxPeIpUKz1TKWd640HqMain+R
SQGvul1kdZp/7atFWO5o/PjMO9lWiQ2uCON4/4NS16yYsgp7GIO2l8CdPpuGfpHh
a06zeEUFl20anKyJWENI5mz1VG5KUKGmVi2+sNgPx1+YPDEA8z47Q6yLV8ajbsF1
mSOet6DPqMij4iFiiHpleRkANzPbcILrknAOXLgzHh5ZZkJTB7wYJI0f86z17DGG
KZL8fZzWtRvthxuYbdOW1DVcx8BAmx1sbq5505RqtHqORmmZTaV1jvwjcLTiJ3bb
P7V9H0HMT1olGyWhZZ8BsKnBbc1Bct9eAD0KCPgH8uM7LletGx3YxE5Tj/6UTafC
XRxR/rgAXv3j3IE/YmAypy34nv6IS62Z6AoUNAt6bf4Rhc3SjnoeYSBa5ajw+5U6
ctQfh526+/rO9RxJ+TVEkxK1358T8X3aNbF+ECDquiHy1HosGFRc/OOfJ6Kz0UVI
AH5DCaei6d0TLsD+Ah2Nceoqlbdel/ClfIJ8us2VlfpcNm3OfxA499qO3vd+vSDV
zq9V8S+TBYiIuz9DB29ij1CWWwiTipon8TFpeh/2PlQHndKL8U/8cwKiHcGsPZR0
S288q+G7i2I8opHj4IjhVTgftVYgRP/N7g6fFtyF6mEQHISvjqQcoeSx2XNJYEMl
9POiYyuoSfScv4lo6e2ika00JCrz9jhmr95zFLI4wJISUObgRamXndC7QheUOKd/
CBzcj06hD7ZXZY/ddxt/m/xUgLoS6/stjkHhkBwlja6EGvLrZo3yiLMvor7fqfmG
L/bTG2FzL7PSbMEAlRgFu9618SK6xv7pf8beYcEyCZNzMq520JjolqBn6FQ8w3l0
MZ1OjGNAbndQC2rmsW1EpTE6BhKB3zs/SGURaMlhsG4t0UypuHvji1NpvnyEDTlD
le6Dqhir6LFCqn6csYS8zxKAzryD4eLfhgPHIt3xwcvPo0fUsXxYY/t5DPRI0OK4
tzmVZsHtPtICn36YjbYBYLtk/U6Hu1GkM6dJyhwEMFYRniGps3Js6Af5XSySMGj1
kX2pzsCiSioXdVRQOFvizTfibCb5fZE+exnB/KF4ADNG0tjEUT87/qFgDQ0gCDbq
YxWSIClJhsFHffqfuquGycmewa1a1HCC8wgbo9LcxQtbpzulSKananU0RuzBVWEj
JgT2Wh1R+1NgLIGZIG0l9dmwBjdT2ytGs/p8aj6JM1iiuxw6SfYoyiH6XmIug8S1
1gwJKgsr73QW7qolWhWnyLzhjbqUXFYqh/QIPUrfvYJnNOb8Bk1tCyZvms1wm59C
PDwNMVxSOh27Kc0rpkoC8cHmbtqvJzhaRHV5ZjYoQAmkZe5UAq+SQCqD4El3sfKF
+mddnM68JGVbJnkW5I7aI/UbqvMrbg1k4zSgqbixZ9DwcEXZEHStfkpxhaXX9JIn
DEN9ohyC7MGlV+feuPN+cndpwnw1J6LWVMh7Thbfs4UiPPi34BS3XJjd9As4ifL0
bszR4r1mAPi/u4ZnoY2NLzWmnI5W6xdt2BX4HZ9si8h4YA17vFnnUgYOUx43WYic
ecQwjshtWt7bkJmsUS2Pai3bn/if+ybe7ACO6bLFZ2LUwSw53hZ55+ddWG573/oX
7jChJxsI90USx3nDKA05k+b1mnX/wmamnREGTtUrl37birlnXV/VztF1UxTSysbs
PKNF7L/fxcf2g2txwzx+ZEhCyAsv4EsllYSbBTaEUHz0Esc2Y/xjSFcmjJEd1MZU
xx08bFqOql8ux6/b+Jsr+Pa03miSh8Ps18qJ77nmn8sSQ+0sJkBNRu5zx58px/qM
wM4YRy5MOds9kA0rzp+dg6kD+2MMq4/CsfQrNRIEzmnq95/sZGNhpOZcWUVkxwyP
9TUAbzJPuSODXt3kUh6nen4MdLNfXdIFJtTSy2bpBZaVZUqFaFe7BnldojHmPp5p
1xD8L/3EMs2wTHt1jHu06jrmib8qHo+Sr/qBT1wp8tH8GAITvgioHmcbK+9ocDf6
UrxA94sdzapUNQDX1faOovaZofWI3nIlklIFQPd3ECMf/ZL2tJ4QxnoV1zQ6+fBL
6xo796lnyGKNecQ6Z2Op0ZRhBM1LKbkkWpWPEBvA6VqJo3FTePlN4XusQtyL328v
guNWTaOpPl3+JM+jARAL4lrRge+U64zMzXFInaHYvrVSMHZUfA9wJwuvfd9v6h8R
St8DarAX6RlN+KAbrCejY73fK7ssXDbsLYkNgWwouDwgs0hTess69Ghc+XwWnJ/U
JUsl76EJSn4qGJSu61COEH0x9kpmNJsGQyrRxkouGg3kPOpKTs1XaSfb/o2PntPa
UE/t6EiSAfABSaZSt5cF4AzqdElTNEgDEch9BHcEa8tdFSnwYF2I5d5tQbZZ6rOa
QvnhqtdThTVWN8z/YS2LTeekE0zJilOEdnXrsNR/KPctVh4lRgZUUesZwu9pqkZn
z6ee5qaTPIH+7LnTw/4y6sydS45tXm/MaxTcrui7zvU+hhldfraxnen33iUiLct6
R7OHc/vKMv11shuVeKCsw08Ho43hmaWlN4jh1whTajnD93//Dv8yyZYerW0VZ6Uc
E4QXNGUmT3IsC+U36o/N4NX1unYXD4O/wTTSLZLqwBSmGYtj+dGpUL1CwznGu4XL
x6is4sOY3MUUOnZCzTIR30BpfgYuiD0JnLr+f+QMckR7ww2SSzh1uRRWLBddkrsZ
SBMTJwgdHz8cIF+dBFnC+XWsKWYiILYsB0IXecf36VGz9fOI8ePpmivJEOnYL80s
FeLw3ekb8cl4z0kxHWtzZT7SiItKwDTCn3ZB6YxcITa9NiIiULVksvjwOoZOh1Zq
IdCNUwJm7TxFk84+JKDKiA407oe6C6FZo0jYU5SsopfWC+q7UnLETbBF00Ov9+mj
jdNQNDswPVun4oiBuW/UZpz7F8zfde/FWonnc6S4pQb2gtDYsYBRoz5pGt0I/8Eu
azHKiObeNGVH12fWbcmGfVMqq2Gq/iBZHXc+1RCAMYwasgaWp8hXDBKg5QEtVnVE
ApaD7rIoh37mn7EkAqxzyMMB06O9wtD8k1t00LDHeuxEjl9fS6IB1pvSSFDy9AOX
dUJQ69WL4qb/ju9BAq9mzmyl7TMpL3At6zMt+nY0avQ3JZ2EV6qK/cqdZgWKf+gp
HQnHjLP7N6YxHp2C0MKMSCnmRCL3KAVIv6rIMKQweqOUv9TrO7kIOVzFjXZxZKiG
n6t3/YIJZJ9b0NttZxci7AWmUVMgxJYHBov/aYvbHXuJY2BAsNb5T5t1GVecWtOf
sSv8B3rTQfxbGIM0eb4DC6lvvT52AnDFRqY/0QwPGjkdk3Plvz6MylMwdQuMbAuQ
18ZEKfvjn2sd/1mGnB52UEQHKEX5yb9nvq/1jU8+L9CnjZl0wUq/J0S65MNSamWD
T6zl/+D3gxcpR6v+kFZ3vUjoOimFMmJnkR8/QvPXYDegrl7ZvQml0u0hFc6iYXZT
JsYbuZstUS5Qb2chFvd3B9d5VA58Is56YFEpdLH3lRhN2dmCYLWPOXXvY6TF+psh
uTUmZeQDvmXgZPJ3F2b02nvrfbxWtoA1GknmoprwjoihehCxIvg8AX4fMYvio29T
uiwDWa7xTqdjrhRhkH856sX46MArKmGRQWr82Ntb7Y8w0hnWEQQF7mbxbR6K4Bp6
UKZP5O9z/Cy204t/Q3QQtWYQulDbmFvMDPm+UdnhvvkE1sGgSG7IRqQUqMT2Srhx
x3vR9rzb5aHDSNHTqGV0RzO195cLcdE81J82xWmrff+TnQlDA7ySZ0i2ZEDuWIj5
Eb9H+/KvgNH3J0qCV3Z+wn9pDHX1YCTq8KHXeXa5IkUIfUgdfS31fSiFC4V9FI3h
j34gwIZEkfWYXGD1qntiAJp4Ah5UdCb5re7ZWW+pnRbTSlRVM7Hp2y6zFdD8cKhM
nMVchuIBTWo0Ug6EMo8siRLhaWAQ0OPxz0XKKi0mpWOmLipq+fHjp2LRFel7Krnk
keJmGCzqzGnovhVF5XVwL1I7nNyp9RGH1KPRtRFj0a2Klqi9vLHK1M1iDWh1inIT
Z/wslS7ILbE6XREChNrfgEWQCJjvlis3v2pCiu47VzDGw33Y/JTzHAqrSpaipCTA
qkJg3i4GnS+FmloS4dHRWAKxJlTeWZIwVduDINRNrp5jJREqgC8ie5Gnhcau63xO
ZlmqfT6sjIYtaMrxfqRbCteRDY8ra3sPtpDHgAD4ViZcIzdD9q+7QLfoOmvJgB+r
Ko8IC/UtcU0OOiwAIU2v0O3akJCkd8Fw7UfOeYqAtEv7n9euX3bEVn7w7U0IY3K2
rdhG+LPjp+XQnKNGKDMLKuwyeqstqVn4k9t6faVLxgWJ/fAExXHyQ77rf8smyWbK
nBJqF6/HAuTloBKzcD2tvRuvsOQT8/r5Rr2iImDy1oEY6/vR6UPSo5BeyHWE9LoK
mcL8/w+e4+tgp5UUDHt/GQiFAO6Oh1VFWLgSa4vnNvXs8Rkd7emjYVEkCfGRLTUj
vBjpjG5igQ8nx6Kq+9k5diBvSSA67RQNwpjc+aM6BjgT1/tXrIdHIXuZpGqShtVW
XwFFXrCppsrEaPQ8arovuK+cQcbzDFt0TW6XnGdAfBxPIM9ZQEh861JQZZ2b+02r
B7+N0x+ZxQmjDyBmA/2JKPhiUMNdDHPVmydq5TZ+3Wb/aPVwTbSn7wU2KCNKnAo2
Am9ROLNW7pAuYFt+/DPzim5syvyvT8vk67hsfWMscLnxhttOmEs87uTZmBcuxbX/
Qk0TfQsopielUg1S7Tl1h9dt8oKcZ061UEceeA1r4Rwth4j+nIcSJReBOO1mFNtX
0PDn5O9OKXYMlZUfb7pqHHH0JuF0Qb11sk86SlbLD+TnIAiBp0+GFGxedZlxNhmH
8dutM5hsR2U//L7HXCh5gLn/PgCxcqQ8TYZpqwBQwN2cZ/RZcupaz8FYax6X4xGo
MfFICINVqBoXigD5Z80lmNh9mzQ88PoCimV/mYwmSdYFagybRNfhPQUhfWBUq0C/
qfCfMMOO8h1SVD+V0DV/YGzvyjrBuPEQcT6Ie7fVGZiTI2hagXS2ER9cbDYqgQra
3tsUhCfXRvE68O6gV5tewtEvW8dT7Z8FmunUvBaEU9Ni/h2PxwV61RQqt+gpXmOW
7ecU4lp5Y9SqqP7Ul2NhscSClbRT/4xFXLYNMRULxKflkFQADUDFl/NHJO8/EZdi
dmQKpEZ20xnUuxg0uKIXZZNOYHlkykWL80qTS+Ceb5WEFaSqmqwWSu0//ylyTE+G
50iND0Ggeqx5hj7szZiig5fUTvxei9EfEiV6LxHbA3Atyz+xHIJ53DLEY42RtVlr
UnRh1pYt6FnK2e2btbh/e2H8xYP3C+7g0dCC7O/YKgMOXUqtObNwPbrh0zCz8ECu
I3l7Apd5hk8iJ2pE1HDt0H9abq7/wBZaYwwyxoixO/ZndGziHzy0XOWb3H0oFlYI
OWktsCuMl9ct9lPD+8KV9WG6TPToPxr51rgBFKXOGbC3w3Z5aMvmThMrQAhTQhlJ
wGFJ206QsZB/TanQ+mn5D1uWrgvecNl1DNBTO7Iuxgc0DSujI6yd26xTdy8+brUX
UAaHggXock+g2DwrBUu1B95senVGwgxl1uJ0P6U7Hvxm5C1TiG1PPLlFXzMLd9t+
BgsNn5o3llQxPnn0rVF0bH4aCKC84LpsG1/aVlWV48c3eVyXmlhZHlnegVkkJRf7
/unFvLfkvnKinkJwv/DW+5HUc5ulp4S6FxxHnmzUGSuTN3oJPwFojEGYCbXRrtTW
6Abnoeb7kYBXZng3FESVxf4cdI1EYy3h/MMQ9WpaIVMGkTF2EBt4pK1neDW9voEI
YvvuOHF2ICravh2kcu6Uvg3tPl2sy1Mu748xcUCkDGK1qmhMO5DWU0uvWehvH/8a
h1vQUkxHt5xa+IWjKVV4aclDmb2FBZie1DTbQuc/OiDg8ol+/yUF8azJIMW341E9
rTXsJL7HFCezxLKUppcyrBsaItQXlZuP8dKqmvXKpSTM0kalWeLyaJjmf9UJpdE2
80KT4Kihk++EsgHs+ay3qIO9hX+4IQasLo/gzrUH48WQLfTQCLmgKoEqVQ2/A+Vu
yHw2oKwybbAK66kj14HqSlXZATI64IANXVtdVY2B/USIrlCgNQiHradzf0aYls/A
ovo1jmClD0lyq/7lqkB/9UHtVbVTt6HklY6pavi5aB2UlYzipt4U5BhGILCwd+k+
RztsjJ0HsawRVB0yPrI30GuwUvLaMLBthLPIDUC3ywBXdDDppxoRPK9/oviNXc//
s1gzQAYU8dSs+93nnrnHNL31c8ovJeS7Ddd4mYnvD4iPTzHDAMMaLQVXeWhPdGaZ
ETErsxlz5LAJVdCoL6JUvYkxRZF3h3mJN3Mx+jktRWspuQetYe04OT9MslP2QbCG
gYQi61cSudfZV+pMvv+klksc7wvcyKRv4EhebQXMyDZ+WLbM1IJatxU+VLhILlSc
J0wpwht3hZceBtxSsR8gYKwAbw9NSXd9/ck9s09YklpcY943K2Ru/ejawx71JZ/i
xu+RLcFB2dMttVw6N4IaogYHv8migsBVYPw+FC5DRotf87fwkMx0hYyJ86NUPmzz
jp1hEAATnTT3V38nGblpK34Ntw55vUv8DX4R198H00TYFgsjcu8B79ZrhDEylkgR
m1RpDxbROQjIekX5qUAdtotqbWt22wRW6/XyhMM/lBuBEHZ4jdnlyakgAnpUgD7D
vB++6O4KXKAQjXYW/KINNbnsV1Rucf8eEgVuQjjdKiksYhgzuT0la6uKqkhD0LHz
txiYcN4FGEYgvB3C4ezO6dJdKAGpReo/PPNQo2wDm6g3yq0dPe2xFP6YyW9CX73n
ZO8K1Gvt5gBiDd11B7Txm00j+ET50sg4LE/AcavCfWVIwIyEGwDTV6q08OZWcSZ2
kAvZrlqjgL2QD2dlkuu9+bt+doqVmx9V0Ti6b9aNS1gZjNgZVjvaTwXyJT0PXwJc
ns6hLh40BKO9N9hY+xuZMdoODzfhHHchpt6WaRtO+xqdHIms3PibbCJDDTVxp0K8
G9p0o8Lu1D7DlKyEeiX19VH9XuIOZ8CxMlW8gS+zLbaUM+Px+DIZUzbPJZoEhPru
AFgC272wBPxg/29Sc8vXsg2470UGYwqZmhNBFrmgTSEK9q/JUnXDFZTXE8OhQfLe
p9bpocl0TSgQQOQfzAE7TlECWXt+NgNzdjYYbwxU/SeCgjL+ezSnAg18mXx+YSzy
ZPaFwH8MNASZ3eXx3LXQFyFPzIQ56MNla58B7wlBE/9QIZ6DV1mBgbSVYHoghxGW
vMqpzHWNPyPHFU1SaTorlAq9MQc5qdi5Po1omZJvTcroW++68JustgExdi+pxWlO
gDGTDbGQ+4y/5omBnND9zJLKDEoWY0pGq8i1bz5+0VYSLretNuCdmCqhlZggwqun
PUntu5XiLZ6bpBFGPZsgUPbUNTD65zjubeGYVmR/SG9zB/lsgL9eniDAfU3dI9bB
KX+IV5EoC/ExtELatD32fu1Gf5oGzw2u+qzxE6u7/QZ4DFcD0HR/OsMo+ClvCBUQ
YDRJVgM0/Yy9WLJ4XnE1OVjX5nusJJHgxNEdIGfoSTKea/IaNbd2FlppfUm9/Xsp
RPcrblmuLdi+oooZ3CmfWd4MITL/F7xqlzVt/5noiZ1e739tZ3221ZEXOh6Th/Em
9FGH56s/mYhVQcajkdKF8DJceMy/fKVXagEp5eaBIQTigbiUVI+A00/pjB9rMfPr
tQRuaTdMGX20jVNDgs6s8ds8kVMS25NS+F4b88NTGhRIFhrbRyXaFbAxl7rPqZUT
xkjiXO3RFe3hGEruo4qHrBRdFHpYJW5n9QwUAHKKNtsuxyFbaqYku/bH/a+wbqn2
/2fQZXhBEo/0IhN6sh/RNcxFG+ySQvQhYTj5++gGpRWZsC9rbBROFDQtrhj5Najj
nuDLUPW4zui+j8cawqycTPXfrhzSeC7OxZOIxb9B5HI228VM4Ul2TvuBqT3/lQBh
ZjmwQF2qZrpGxKupcati9h45Vux9IG+rZiBvJ3GAdNsh3BDYueVrSmsmQYGvf0v3
YFtqSQOXKYbF+naU2QGvpYZzJ5neSMFKLL69V/pAmxVGnpRiVR/wm+Z6yb//93r8
S7sP/8ZElnr2nNImWmG4CCv4KBVRbGM7ZdVKOTf89zXZi64Eb5XEE6tD99vD+Ca5
xWmC0aF0kxmEc3UFoiRCkeKrVJ8LY98hnuiAOw/46zwRqvEaXv2N4kjKQnJagdfQ
ToBOiz0xVxkW6a5uNMec2TWyxPx2pXTRt2Hc9Z14tcyXrglvoTFwhz5x8IBDprJ6
h9wYWNN8JhlUgvTBQrPPW6F1jcJ9jjU61/qg/q4/MuVKk5EvspdNsjiuHdaA8XTp
AnIWlNz3tEJR3QPRHfXRCPVTmKReY9wHHHdH+5ruvdqIkH0RBGa8qk0pkh5vuU/j
Ddk6vBf0bERO2ev2S/XPa8JxJW2aWg/KtM728afpncLhyk8em7q0SVgT8b4qfhwG
i/ZVWiYVKIu9/tO1ONikIDNoCc8gHxp9vpfYcXlJ4PgVsLSzS4wymrmlMCQwT2Ln
TqcbJ5hBah5Z4ScD/JeKPR77fyFM4DcEDfWii4srSlothJ6iMvHgqrn8ljc2m8QH
7Ftluh/MP4rUyr2imOQCtnr3mn5HlLeM5jv0m+WylrdJuPz/IGMWfOsk2Ljmt5Q+
N42WmjURIT2NqF4nCpiHNOnwvhDCUlY+L1n93gEzAJ0kXgD/is/XdkBZR/8gPwzp
9AGED5qIfyiL04OhBIXeilOI2hLNv2Kpw+U9R9tUmkfmqZHDjpW3uWHAoP1I+gK/
VjaN8zxpagVuHLVA6gEGEyqirK3Hs00IS3AmynBsolfmVdcArcNlfFVcnO2Xd/q4
VfeL09moql2TGQYuhJTsxRZxMCdEtWhO17UuKaVmg5YTpKmPbNt2NrJ6BikeJ2TN
Z8ED2YzjMG/CxtWT11WgWz+cVgQWlo6jxx2x1xRM0XZOdMycTk5NxEDoSUHdr7ik
0JGKxyl7juCnVCx1ENXKFdwQ9gm087rHG+Hw9uKqgWFIMr3BJ0pnwXg4WyN+ddf+
hNSlE6l4jbuozrq5t1XiCvhghY+/NyIBdWkZByZDDKBXx2m63NZ4AHIhvFyRwCwB
NxIZbkdkpv7x4hnQvz3EABwD1e+07vVFyqrc0V3K5Gdt5QlaQUrl4qrWw7+C0RD5
3phNR6IPOdNXHrsx3UYcmSBXP0+1xSVQdtL2U0NuR2LGI5Q2mL7EHBeOjuuuzFza
LuwAM+6tjmXyIRN25qRfJQSb/mZAWI1uvQe5+1IE+uaeMzA5e1lUZt79pMnaBXPa
wTA0+OLQSofFib3hVoO61Q3Z23g0UQ9ATCpFvLw3LtwwiVWd4S3Q7RHRnnan4X9z
mhPW96qc6l73MFfMohoGrBJUdHQtQ8fwvWaW6aoBprN5rCxx8YGzmWKrMXPuKoft
XE1sNgY4oUWABRn/rx4AgPxtFI+92lvlMq+NkSG7FwXpVaTVZ1kj49U+6VY/13K5
XAv3xnADWiZCAzT6ctkMyat4eIZXqnRO8Rnvzp3Q5lDN5kMBy2Kmm84pkrZKN/78
kdfwXtsv2rBIodvV+tbqD3r4W58+q2qbazGdxxL7RfpYOOB6vj7qcnHxdU0whlpq
RjpJJvY5nKDQ/XzH0+OTaamZrs79WoaGf3V8veXHhSLUTL9+vuc2Rw9mZl9fsOFP
NrVH1o/zaaIsLBbjYvMov51cbK3CBLjj2C9Rh25LviAIa07NfAwloW7eYujByOf8
NohmYGxkVvcMLfEsw32wlJN1jWgoVlu660bv+cNJjfGJVibO9q77bPwPBPzmDpZR
KdvN9S9zFujqsZ1GXmQ37unaBmwMjToOmub8wgucJU/7nmSWG9EcUdC0VSwyL3zi
gi/HGHawEYeGd6kTfNfrnJiKk8ZMzSboHYauUIZvcmpTHtDtJU1Qo0UOSLf4tzeB
ovkahQ7FKiqIbjRJn0xyp8VDwnFcO9NEVbhv40t0KCOGtvhm6B0lKrgq47IkpBoA
gwlBWDm0fXhhrS2TpS1xqsYiKa+DlrulhEMLcZ0UL1rTbAfRCbBMXqwuUNM2XykR
OvfylqOWTxBnMmtG8iBsqAUxYwh7NSR4+yr0LCCXgLQQ12RX4yhARihqn5TnAa2C
ZnrR4f27pt45c2XOKdKZy0G5H7W9rU7Uux7BjJrxc8MQNR5pa11SNRzchkpZRjUE
RkxoJqwhvrZd2c24QsF+mabQCiZU7CgXdZM/DPTYzMVhrbuFxU2lzJfFUznG6BqB
JaMn0ZEJVq7DehXTbCsY3RTPpsOVsPsXkKZ6I7PIt4fG9vj+wdq45dm2HomjpqeB
swXqoMi/VuZA0f585h4BPFZwxRYGIK76KV427lEND1pr0x3NcmfmNOAfxhTZGa3o
Y4rI3DR2QupkIjopgkB9pehkEdQ1Kqr8luGmkx31jNpYeHYh3SpohdxITQR802Jt
tBnAgBw9dpylNGgocyvLRwKnx3GkHBMEbV21yVXrarHLoSrHvaWC2htAcbYVL9fq
W8yp516uS+CWcVEFGZFoK4UJzwkb4uMdeGBCMLaP5e0qRTRnqGM+1xVJkPqrH4Ae
9EFTJEz5Bld3gmc/l7fa9Og8bAj7lokp9VSBF8QHgxbQE4+ikNeeMrRIsn0fzR9W
suY0BaEnh4ZBeIc7COEDpfkXNpL+xfHH1lXiISJwEGIMyMYH50IDr+pj3e7jpult
jTzuHkYcKbeptLhWZBABRsE8sz1WJEf98B3hQ39qOyt7lBf0H2/e2zFLmKevnsR3
NfvHA3wo6aZNTfWEEWaoeu6zV5K9Ye4JL8dYNRcm8oUO1m9laAk7O9OZ1so7Xi47
LHFQGfeRkjMMnddQkcludRW0gnze88vYXrOLg88pARQ4BhJaO0acAX/ngKxhoNX1
Ijxaatx7hNSKHiw9ptS34ELhefRgMR+xCYwYrUOs77OzVHcJEOBRmBoPPWrJVCK5
IhHwD0mSngcjAV3ZOHh9eFlxvIA0dkmmrxQ/tJaJRQc+GtNMdCMjm+ntNStL2o0h
SOd4m7EfXMMekYR6duK0TpTOCf/+HQRheaQOUWmFhjZZCUf7YKFwUx6KpbrmU6To
pSt3B0EuTlxkOoceMco6W8uQ7O98zmGsHfQZXkfwOO1dspDnO3xd+V6vjFUhS0ff
qaVXCQ8QXJK5RaFoFNgb4DPgCQAQn99D6Esb38pmpp3QErVp6GKsCu2fN76llTL8
ks9kzfuzjWXr+NgWFqNPiIzvwa/4auBZ1la1U69S/XjjYovskNopqOcmeiz3QB1X
uB+DdUDHC/mW2SIsGEZZWN54v9uSfdICr6Jt2/xzFuXQjAYPrywk0cuaqeyrk30T
agfVVBymRz/p3x//XGdNOqC7Lv/VRMv7RZdEv0KjneJzR7iFhCwY0UDQAkgdfbR7
0sSQZnfKcrX/VUeTIo9qI4KbUI+2kfmSL1+3m70BccE6jgOkUz4hwcAR6EubZBff
98DjlFc/++UUeh8KnrCzJYg4KOJmqf8s4iXCVcHKgubCssjCoutc9ptOMgrDRFqt
bcQaSHTSyuukZSQ9LlPHfuWeUG7nG9aIMInV41v+HH9DB7KZeIr361OIo2tyEkoK
BGWGDq84G8RIlrMBb5Wsrp4M1UfjI3LiXOTTCgQKkhNYd1ejEl1P/WL4xRvtEajx
JuQst+NX76F+gZuFEt00cHpp3KnSMl1KuSYSXiltJakIMNFyhHD97GlazsOHqP4a
w4Zbk5++gl4AUqiNesu+84WBs9MCdEN30bVQkdo2crKz9yZX0IXP1hId5R9Plv8r
lBf7hpV3+f1CqAcE4rm9wEVOOtm1vnkbHVGjnTgphdRyQB496225g1hcMCE7oJED
Q3CLdOlUDI7AgClcR2odQxWqtgN5vYCEnm/++Y+VhSxDJ1L5S2shUDfh5ARP93P5
dj9W1otTfkETjXNpv6hC/8pgAShUvN5PTVK/8kVXLl3sXQ9yBQfDRaiq4QvvvxbJ
JGuJUlphoc2JXcIzNKQMGIg4sV2LVVOecq9ltBLkybXcguGbWIZCB45SfyqZ3C7l
NXpg291RJTxtapOoWTk5o1elk72D28gKaNPrbGneeNaDRF773Oszn/1LlaOk9s/t
dEo2ugxovc9E52SfSljiIVCpXYsKZac95IVphmH9y/vN6DzSc92KmYkcjzuO9wuA
OTpqSL9js1GXIYkWKaRn3CqJi9Io4mUOAAoql2AWFXTFzLfI8PHysEZw/0pxExXu
ctHQfcm2bFUBV6E1ERyLy7OsgiPzPhGCxE2ECQ+hiIN9yPLs3yDBOaa//6dLG7QM
/3qbcP5ZlTLhaepqU6/RRhGCnxLoDRUil1UQgGhb+NaPJ5Gxi5w/lWgvTgJObhnx
vHVqkQbKCVR3C1I3wAJBMNrfwC1qXIqmu58KNDZuAe6ycvK1KAOGyQLSDwyM/z22
HIim1nEew6hlq4SYJIwPEdIewxzWvAk4BDdasD2/GZaOX8C366ppI8I39mwMtQiB
Rlc0hvFLcpla79AVAwgC3xjgcuNC9X57uUL+4r0adcx3EZw+aFiSnelmuAlG3sb4
JXUAeQZ822QfQquKZvjAGm8tkg3+MPWu1d/g7jo+pJEDeQnJk/cgkKdu+bEB7xg8
gbiE2x8dmXzDzceVOEBNM6Mr4ighuH6/I7n49HaZNaJ+7VxUDJD39BqW7PrFHVoE
xBwLknHcsbCFC5M8suUw/i2Hy24+8S7aoqSw9mmc/oOgSTu4mRpwkCrm59SAo2lM
xbfO7apMafWv6dgCTmmm/x+3+riWh0Y9OkSahmctA9JgpaUxLmTQlosTnA1k6SW2
O51xnjLrfim3kqXGhe/RCKY8osg4kffKj8rAbskw/Nu2nlIg2nckAQxAiYynYkTX
eZ0h9yMVKas3WVMGkScUqCM8SdcDS/22LtT6QTQxV8ykq9l8Unumaen6js6CO01H
vvTXTzN5bkCVTHpjkvy7CLGMoNOMBxzJZ1wX8qhM2Gt/lskpqZZnu9hE685wHQ1r
5oaqwcfYMzFSM6gx64KM3B+Zt0h2OMPDtt1pYiIHZ7jrsHVaUdjmJMB4pBU/iYQR
TS9Nnc9+LpT4AU3abDIMLuvPgjsDs26EXn296LdJBk0rr5dN0OUbhZlTbkP1l5YQ
HRVYBnkr9RwOuqjdJ+kEEfGH2jCW4hocSd54/BnYtT8Pj2DBeriVFLttKCHeRXdO
eBDnLjoYxLyF+CdTmgLPfuCwCZZQoWfJpAXxmy7n2Qbv0SdXWagcI/yLXhpkQn0Q
b+A08TAXGW7B8HQS8roLH87DT/ekqMqQGGDXOFCdIHky7aT0oLXg/cRWqzIX0d8h
CcIajhyMz9PzrHO5YwAwW7POljvOJpi9W6b3SuIA5WBf2rdJj/YRoUiBL1jt6p7N
HwCJrJ5/QBBUMVkUaBRNtSXa97ShVqWIMoYfFkiZGrbvRUl2F2XsEDHGPIjKiLjQ
UGH4ny6XRSQ394kCMi4jgibUs2EXWlgH3CC9xVMWI1Hq9qXTjiwtmXvk+gZnE3mh
D/1qzq7K6jgIy9fG30BESjL4vOHQzTZWsZ20Qr+4K3TKw/uRq8mvGmxrVb4pqOKM
tbiGna/JpNBYUC/hiZjAqLhHyn1aZFnZj+MxNvA1kee+tClqVKcOBDUSBNz8J3jM
GOphhlILFFtVRa7HuZMXRWfdybL28EqSIE3DYK/YeXp9uAZ+xWsIxkfWFJCG3Z/E
fKFg7kpRDPU165TTSdS9QSKfuPNJB1jG1seInGtQQiFMNe8SX1+1jh3ruHlB3ixA
Aj4kWIOrdcjNlmcmGFmpCe9J5+m+VMEF8NdOy3pwh4tYHxuDCc6tOnXWlVG0TTuB
QwzkEcvWxat6eSPDEvPxnq0Vv+T0s3eGf7qF18yEeQKVXLt9bYdLkfrTiZz19VoC
muGQ/Vi9ZrTtfXfEAa4k2UqLJb/p1BmnH2Yqk0l0VOH9POeqG5MUPEbd4FiZBP0U
jIeLWlhyxpECQQuMGGfujBlJqR0W25hlQ7l7zZqOkDyIFxCXgm/drXFxghH+ENhY
xEErN9IqXSfuLd7gebv7IxemO1RhkaHNeXM04bjKAjm9bXPxuwZi5+br768leH9Q
pKzQFcmIuKFUZv3VUWputltTjZUXNEIP8fZ8O3Rza7sgfkp5UfkkfSFe7pAovWeo
tAyBuSwS4ZIKl/wRJa/hbWXxdBDDE+wiYEzlWFO8V/fjX0Yp9ftjhEk3JeIgG8ZZ
ROReo9wERSl4LfCLqMOJBwqIc1RUP+Lsen0hHHwFDKhgSI9G3VrGn7utgxOGQJwd
qn+RTFHFPhvrP3Rg3IhfcT7gSJvu3oxclVUjPRaaAMbnLkKQdmNmnp+7PZnVqIGZ
nximu8wmF2+CmUzKdr5pXFPVeWk5diBGm3hHb4FO7jpD8wOhEYFCznjnTCkEsubM
hSCYSqL/TnuId5Ld8CXToVVu0XoY6IV1pLTohEGYtgvlBkXWRRBvHM2YjYSyJ4I8
uq0DCyUts7ix1vomono+xPMxaBpvN3B4hy5iH/em9E2eVc30RuGg9alju80y4hz6
pkT5uitkCrbBKpZr4kVIGVscGY+t+RJmh2qDY5kQIQy+/MkVCckV55lsXzngUjFN
nadduR2mB8SdnUNYFcqC6bkj5EcCl7xiOUtyDAB1ZnsMS0e/uJ56Dcn+eAgxB+V6
J/xh6iu7MMYtYO0cfkVkcuOGUmbx6K8hqmrFqmUR1kgApQOWRsVNGr4LNBjH69JZ
o32bO0Tu3YKxL6Vw1GeEp7PP7fUExEFjCjgenFXDHfxfDVJvqLFbvVhFcyJU6F1U
BouSy8eIE4kqZcsXmdFnuBMOKyd05UdOQab3HNLo1mVuuu+TjJBK0gFISZdhuuq5
0cX+2/pueitXbVQH9xC+7ovnmeFc8CtghdCi9MaLz3MlWpSM7lPONLifOjLfwDfL
h+UFdCwEpi8KzMzojeWK9SLwEB5n7AE1n7z0PSCXe/8KUwmtBhaWD28hLMoiEn7c
sxcsNK3TLwv/CjWEWSGyzfVLWY51CpOUleO2conGwZ26+/NSYktY6qUZO13H/qxX
+QWriN/H6ov3rEViBxW+y44HmHUN/Z11QuTNUeac4q39/tJeKS51cfOvYgGz9rHf
uC4aeimi1shMHWzWuEsn8gYCRt13BYP3emKPIZFBvIoVOLxURKmrr61GyoH0oMoj
rWqbeIq3G4/5+7T4XlZFNlL30jDI8DSHBoHp4Kidn6V0UWoJiF5igQX5m8k+HOxb
Kg535ZXOOIWIhlRWluUJK9bBQJn0Hf1bcnqh2wtW+9zXBADXru5651oQpbIusQyv
1r+PnCxcaqBYMZ4Wi+h4ZtzjPVkJtVKu6Yfxw1XGD9EPtRKBBNuC8Umc2tfboIQj
RoM8c5iRB1ZGMDcQ7mxpkg3gu1I/9IcslV118C9s8qDxcgVxq3Yfm22i/IwWjK/d
oKgfK2qm91duFQQiMm3NwWmlY53CT8hKDccWUSLQB4hLwpbUcspkeSbJ785POF0R
34B/iWZimZot5Y5eGs6TWBxt0rH6m7b3Su8os9m43W3Cs1dMdQnUhtFFTLTh+t8z
UWIGmTsY/5561cmPVI5KS7Uivr7s2Itz5rP1BfUn2wj7j4rL1Fx867Fq7lO4WIpu
D+gSNJxhLL2L29XCVZEqP/BvMQDDaXoO+ZdPvxezRIddpjdqRRLR7+Uka2hm0KM4
0Dg3ABR7msh23FTahhDDfZgW7E2cykj1bTzpBF1n2YsoutwogAACndMdRAzht+vP
Kjo05EHt61zDEmR+P2I0ZferERBFfLw3Pgf4EiF4LwleYLqvrXNZlX9UdYim2HMd
s+xkJxC9HA+hUJ+4aZc6sjqsf+thEDCRJ/+842qYlgzvReMOBd35uTjh8ygLWOLI
mjgHODk/ltfnBs8+GA5jSZ5FTuNfiBsnayk1cdHpAUqQtkenojSp6PNiaJjidw3o
4kTlfWIOkqfiyKe7Vqj7itCdzEwGNTRuO4kUGHXdagf/isQuv2i/OrnUqWyRXAgv
Fub7+jDf4c3Ioh9IWbD5T5Br3gBpNov6R2O04O/22nr/obGPRt03lBBNin5zW3Ep
yzC0sJ7fEkJqJCse5XI5Bg2Zo8lSTXTIY2qW9DhustUfgmzWyuoosOFKswXtBGOH
BiuzTJlSg0KIRFOxdrurGcBu+U75iIr47vxev0KIPFlOTn17sC1eqasBme9HKUAm
QUgjkxNHQUdM24Y13fOHWCqp8i+EfhXm3OJ75UKGnibDeETGUaJhZuA5x+sqnVMz
SrodetoRslDHKy6Sdb9zYor28Iuaq0zi7/qbqyxMKzBlxidwWZ/73KAjRZBsQ1xm
j1NjUuSkszkHuQM0hwj2tTRg3tOELLsaEBD4qsC3/LQlrCjfUc0FokFTVFMvHfdV
cHSXEZ6+Hd3XF9amRAtlKSDaiQYh7d2dV4bb5UbQpVdws50bHegS7FI6jIMnFVjn
WmucqCUT6FM3wqo2ApbVB5qSvHXJXc/JTQlHYSXXzKrL8Q57Rd4+AFMYwQCei4aT
TOgusXIGEUaT270DVW08KNv0w9IZLiWUJ8Q75zTd9iBJuXeYFKcfXg94vyb+0nQW
7CpFhasZ4FT9yQI/y9VWBi4Nr9XSlJSwL+/lcZLDTuDOY/0lxt1MtNWbYgPjJ+Zz
Fx7UpQU99USkdJE9kpx16O0hiU8Hxe++IQT2hF/9qz511Eqo5KT2cgYiXgtnlZon
5dl3BpvIqi5JQExTtFmsIxT1u1S5HNrDaLt8s3xzfx1vxYQGdD3A+4dxRRM/xYZy
RqL3bjDMObNcJrfokBizR8lItXErJBu908VUcYt/cfUIQuX5DnldNcSHMCywRdfY
56Se9rJdrGGRfrlc70QxcFFJBd3U8fAc0/8jitXIbrM7/7OVU1qSeBjV9ZSpy38k
MOP9eVLurX4YnTvjOwi8O2IwLUt6De7hUuP0obh+s1xnLce9ZC44K+RIR20nTW06
2TWsFQUAPwn/QhluRBuatEGJ8a9M7vDyW/Ok/MS2B8e9B2D8tJHK3m15b0FdN9ds
BUhNKkCX1x4Qnwug2uonSNrUZOQudz4cCPtoiA+18PYDE/pZWRaVtroFj7BgZdJk
+SxaVueiwOlKUX1agAf5Z9TS7K7owpC9kpeZ6ezvnNnI98+FFPxacwRrlqwsHKIy
uqr1oyc+KBpQJ0A+yBY9h7z7tCqEn15hViyld5hUOYvCFYv8hLXMTyWhVNjTiS8b
mSuoi8t2dLLIJXhGkC8xbZ9Iles9IgJSbspLue6stucxLOHkrcPK8+D9mjZJr6qW
KNeDmDSiDAHljI5EW10WSI9R87YJcLLb+oMQ9rf4HeR7nyEZORXaXGQgXPjy3KNw
5sXhkh2CH7T5pDyiM9fQbYtU0Ag1op1g3vB4wqtx8hxw65nmoHpDnKp48Qu+SRsn
OK2N9iu11hbY2Z4XhxiIyrLajzAfOM6Qijh78Nn5/e8D710lmegbWG3yi6AZFbAY
2gsmYmd02pS9h7I9m17363bi9YhuzFXY9lnMny0djxdZMGCH97rCDmpHrCNUP02W
4T+RYU57w4lTWQSKzgARRqVFBoQsoN858QjejbPd347zqgJkgtOEoQqxySuPdCPC
I9sPMWGBxIwi1e71VzUzqklJpe3bE8tuXuXahSYSd4X7mRpM2/cpf6R3P0XSZzve
xRlUqksThMNSs721R1HYlh1o6PntHltdg0jNGWEXoUn7tXs040AFEpGWhNTQkoz7
9bcmQT08oHnpznZ6Lie6dYtMNOQ5lfWsqglHnUGYsdOKRbidlYp5ar5lSeyxIGyZ
eFBwzqqk8bQroPUXLp7S6WL/p+7FFhlqdyLpsFJm3ptz8bsUpYQsqeNLwmi6ms7L
xkxVrorQmctdq4O415pDt+Egfzdlp5aarYqWGQ5G9y+tA9PaqDl1WAzcjPqGk2Q+
eFm7AZHzrmBVGb6Fxj6MJ3Cgxj1eA7h+sH4GD5Wsu36U+cfec/DEpoDqYGnw6rQf
wB5JD+fYnVRT478Q5XxndVDMvKM+uiL0XDAb1EtBWs7gTbYt5kfWQQUuY7GO7zOG
6Saq9WCYk0XtsRhRGnRUYQARby+8Kp7/9hfPLF483nb4y7JxTQNQBQoIbhvBUo+m
p5cZuw4IAucxaDj0pqK+N5xwiyqI0VY+Ztz/zuJxZTxtUk6EqLoAFS6cVpIkUjUf
EaSK7qzt3i6ziLdflDH1lLXR/uteR+5zMJ5B2OtzMLPFTVfxL+32ePFdogIl/pHn
CkxLG2+zpaVXsVbGzxefWZpTpaSyUDAYhQQ9peF/V6lArTi4O5RbdiMaIM/pAmK7
dL3m+rtI13BG9HtIm5PqQymnMr+55m49lHZHL+sQNphzLxFRN2tbGxPWfKNlC7Qq
AURMGEkURhnVxrY9W+aRIUVSerurco8guVbMIawLDUMA27xqKl7m1KSWPqLQMnaY
j5rJpdh+B3KbU4Swpyw1Zh3Rqj48HP21x1b72yDOocx3cFjnYMijky4V6+JUoRpq
MEWKFpoeSlwXSffGvGdzHv4FNRTfXhfTIfL6NuBsAZundXyUg4le9gdeL/BIdJYa
ef+M10PFfOUykWOHW0JTxrYve9mjRnfYlKdXPpd4CPn7jTeZtdpEiv+jDHbpONTE
SA4xk26QL2zSdv9cZkBG8bleU7/kyH4N+hAWwu4WMsp9lUxs81E+tdt1IKCptxme
jKNf8P/i8Fao3BAFsFU8eQbD9guQheYy338OzNSqp41DOhqe7CQMYTWTyRu+WlRe
QDYxb+uc1FflCD0hWC5tBcKZQodDvpyIZd+J6N6kjsFK1KvDhJC3EiHTQR/rGN3W
6uBxh11PaEWDvy6YpFeThVvSpB1QohgH5tVzkVS7P0grhg1OG9S1w2THikM2fdeH
AP3OXhyks3q9J44cz508X9LHE1uIb6RC7HuWlbt5ZUwtitiYqmfWZgzH9xnG+gDN
tYhEKyd86dx6ezTaUVCVHO3scnQUEJzR3647+F7+uFGCaL4uA/KZAHq52pKqutTH
sHRCyWAl0By9NC2GBIZEbK+D3paLvzz1Yp4doFFz7EgWv/QV+x0ufivieeh7JTRW
RgnRkauKlKu8mOYFFpf4y71GIpkBLbOFu+HUwbMxwuKdtpAcktacRSOI4jAKsIUa
JV1A7dBHN/WZGg2LIpvcNqTocZ473r3wtrdIpd6syWmpnhD6A2AohVpExhCq3oc2
Dmlo/owjti/AhS1FUyi6qn3/XWYkFVCRe2irFASP/YILWnPfpO7fXkO0+2gAWxwc
Z7FvoUvrUkM1ygpYz07uOyNr+gfi5ZnlBrqlKqBF4s61frWszZqZjyFjFWMEmuT6
CB88qc7H1vD/8eowrAqqw2eF0dLLER78AWcHeH8sEZGQT5MquB1eAUCamgHf6BsU
kpFW6F3nLBbxFobts/OiGNGRYwfFxQAA5mwZwQbN+jdLNRnRvyqB/Zb6PLigHSG2
qU3uYW5+aEarQxpw6+nCC6lNgOovA48beKq97fK1iDJhTRMEyJ6qTgGQoEtX3ZWK
4J9StqOi7RNopaZ0bUtS8CFyPbMmkEAf3IWumJ7iG1HP+nBS2AtCWImys0H5K3fh
EifEnACkVcZq1tTfLZMImQd2vqUoEjKEf+4UKyWtkn6Ue1y7W3GyUHjg5+9SPEQG
yRD8RPqCaw0/l5kiBjylB9UJ8Z3G66BfNJ/8i4SSKStQBJF2OhfWuVj+Jn15+lin
M61lloA44hVCw/91Kcj50d7hb7Zp41ynM6q1xah48yAlurS64gnnYK/YfVliWT9Z
F/xT7FUQHRB1RkWJYQdVUmyJVSa2Avc7MJbqz2RYk5Z0Zk79sNjqCAjrM3wDJrte
IatALupnT9EfN6yPY56EX12ekP8tSRP6x77S8R0PkkvXHUxd8H7JjPe7mfhvbOfE
b4NXCSTc2k/+2Zx/8nChssTQ/cQ272ExI5w2P5e0AyyJVNdM9e8H9kmHxF2z39Ch
EHKOz2H+nsW8/JqAWvkNhZVshUeQbIJAkz0/UOTOg9EHhaYYoV8lRSKkXcQKXVgx
eJ46r2nwr18wO+4ydlxvldiE90PSo6chKbZ5z1BywQxp7LqpEihsdq6WF9RqVyJ7
kPRItP7exdERMh9UmtoD//N7j495QDhMgYBxWNcaubYeW66X6jZ29FNh9Te42xJ8
AOin3EJb8siUwWvOclxUp49WRNwMwbq34o/Kaeh6c4SBnOFbKQT3Onn2STHpnjIW
J4pzPW1xWE82VJYiLdwV/KtiB+15IzyjyOGvK3hNASYSdxdu7eZ3D4Hfm/b+ke1A
bdD9wMRNl1QQvRlPB+NJdvHKpcSDRo9Z/Cm3/MLgeWm5NHpv2F39tepkO+FJZlEo
O8NRzML5Gm3kujrQ7qLw1ENWiG9PluSgpg5Am642fE0ydmuVAjcCujoMup/iL0aI
wXM9hhBsizC+xT9e1EErR9hi47xdoOIdsrMUTm2yP5fXGhNmxLsmPO+ov1BpLeLq
fEpjA76fbWXmEJw+HYH7N/fJuMqMwJwMhOJL1HjqSjrT/Xrnt9rL4RcfIxde9W2E
zmKsJv2nH7ANrCH5Rd33eu121UKtbYc1UM9jPfrgCnCNSfvhk7Z9HMsxgq2PMtpu
z9oxJ7TY4lzm+xttn9RDP5BiTjdH8YnHYyRA5GmmXAAaIU8a0KLfXggZnPr8xImS
n/2fP4W7LjUWCgXp5wwmE792hx13xKZTjVbqLKGZr7FDzGMYcpDm4KqTjUVGtCi8
VVSQ10TnPvEtr2GYNsY2i8AcEOyCybZszdd7HxY+nGLDyw/g80akI7dRrPOgfhp4
0eXirV7hTHXwWbvZavRS1CSebQZatfS9u21ZgUAoJCctjxlZfBqySm7Hft3HQ3nd
vDdlJtdrXIXMBQVbscoEal0rodGEL7rIG46x5drlZSr2iunXy/tWX4rq8Q9n9OBP
/lpnaRhvCXJUAgYrggMVqJ4FmBq5guG4gb1qkb03laz0y2VPWe2Rq4JEgPOXSn+W
RN9J59ETQ2JwsTyWXq3gBwUpaXom85RIjU377pecGB8pKmB/LCD2wT8lIZrQDtA1
1jXPGfG5SgII+wZyNqxNpcwMCW2av2ygkloB7Jaz8VgHlr1TgaA8Swv9mtxM4YkA
ah2A9kpWg1L3FtrELE5LTsAGeFFeUdFzd2E9OmYpWpHQASJRkRpo4KdJx4a+2NJT
Mi3Qam2oWTbN74n/b/g4mUzG23ADdEVfpBUMn10+iJqsAIkliFIYosBJuKJ/TEZO
RCP2ts8J2U14e5VRZL3/3vB10Pux9oc5DkrWBYT92j4s/BICqWEtMwf5BuhoV4te
6ICQcSSsi240p4lcdHpUyXAemstMPrxlbT2ov8KkK5sFSwNrangnvCtBKonH90v4
Ah5NgBpcQc4B49Cu9aAv/J3IKWVZSVMNnQcaAk9RePUC3IfP+u5mBUNKJWcR5c5+
UwwtJTga4jqYWgxrV3xkfdfHvwWIdntd8stBUPN+0Dug0/1e9HNlN5AQubYaB5/z
lUIp8lS0TsktVyyq7HdykaMk2rqQ1FNKMM/QF3X7exMJ2TqXnHVr56A3VLj//75X
XvULsdL+xeZIXOXzm62NGQxURzpbUL5ESPu/ErENejGDno5rjCqGZyZUqdJsqYkZ
76RYUjTNJtGNODmA0qv+o60oRX02OTbFzmebdT0473NRQPTjh5IX6JxwkVtgu4PC
jiH5WjqQcacuc4e1ZECgpg2l1HowfII34waDfOzKd3Fy3Ir2x19MDp1PUrgmpP5I
spivfmErH5ouPppA/f2FYZwcLBIONXmtbHsz7BB0BVA1ErZ8AnhAnuLMC2GO2cVo
N2nMmqPE0WmG+luF1uS8L6YHCvuRl5GuDhh3z0/JvhYv1ijxYebXbS8J8uhriNcr
l1zsz6x9hXsYTbt158Eh3rYOmDaojrS7ocLnDVdU95I+mrujA9uDt4iuFvG/ZpGk
PFy/172teT4pYktPUkhujcN/lud5wPln6ItiGBQrlcYOU3TaOKwrnMeG1/Hnv7tN
Feiq5Vf0Zgvoh9oNGokid1TQmrZCDEp0dBBCF+1DeJLPwvpLur0uK3AQoYPSUWiP
/ntahQyZ0juQ09yFUxXrV0eCUXrC5jZ5zIn+LU0Ly2Kgnd5bU/pS048/pBzstQ84
/MAXrT4ND/NEbQhJm+qw8UeDS5SoHBLndj/UxJAFPzhrXVeytvf5aX5LChNOdVm3
wl6MXrmaF8V/KxnJuuT+FrsTCtHxvtyglTsAqbSWvDOTepNXG38kXtriz6w+ofiX
8qKlAbthhKR5+r08T5xCuXC5MqipVQ79bOhHdgI7oJZLyo++f4FaxXxmWpOJ1oUy
sxbzYKJgy2YKR/ioCi3Md1KRRgy09oNWxL+93GOEMt15EwpWK2N44q8UQcBGsHZG
Grq+Sat/WUfBegtA5iMre++b0X33HdpBbGdtoWxel26g/UxXN63A63MvGquo+rBs
m70WOfqhiSVv7lkRxvFKleh6+tgdW9yk+jBnlBARvVIubfNYJV185MtsMLproEcX
DbIGkcDpClYsQx/vw1LBFl9Ym+LAESKn36B4vwLFB43RmaNtpgbfxfYc7Lh7hrPp
JxK1lkrVCVFyz3TESdwLNSAROoRKXhAzKZeT644+p+CImYqPFLWX6DVPVEgQ496Q
4w5IYM9K8YmzKtHr/sHHrOb7Rt0/hMR8lxpg3gvOMgfDQnAJKSUFDU024hCy6ii/
9n6l2jQkNzp8Li9FWDNSBp/gP4zQR9vCAGWtt0uNjK1/iIe7iOmFGcgwFFDE5QxQ
LpbB4AIkJ73Qa1Mjz3xCWpwIB9K5JjOo/v0vVGGLd0jRMOmKY0GmlcqhLeHh6701
qe5XMF09tp9PX+e3RELqA+1yxTBtjm4Vy8lrQQ5NLyv8kCdbA08RQbsUOnTFACFB
/eoFwYyi5pz4dYb+k2nIxT6dhsnqFUyY04DEo9Wop03kkcPGInS4TQtH/x2C+x2R
uHAIZTM1gwkgK4OPCrD7YuQ9IeVbQfzgb4R/f0gP9ybIoXv8qk+AZMacEqrBT/ye
qRZJ8/zt/MmHln+ztdq3uS3TskTief5wElbFj64nWfaXw6WCfDQRivNwmmx14Pin
d+7JjGVqetsnWW7ZYB3nSxjJ1ZOI7gxnzksdEYxx0YhInNASSzO0n1/fk1dYpjQi
NKKvYiJLDzau1NQlMbN+eg7eku/Se0Mu6lOp1t3n7NhR7IuHzV+euanyntZCL8Z3
POGov5/4lC7RPFrXjK/VwoNe+lx3vhIQMBL3FNTzgZVeUB9VpjvZmZl2+i2ztbSD
s68Eu4VD//niCBeGsOKOYTHhSCYxR6BZcktdhCGAjg/EzrKEKcqfEz/pvKMI3Acx
zV0FRUJcLpPadeTuFHrxF8ydVWeA5gCU+kROHB3d7HQfx9dNjdwfpenps1y8IuVB
uHgEHrgCrokgFzYfHp3XdqiRssLz3yJw/n3BlpOaZUDSnhuwRIkBwBLX6vV9LnEk
IoWZv97A4fEZ008l5QdQEQvxzceh5Gn1xNvJPzLEfLCS7Z4VheBJiKC8S2GOpxoq
xmbiScDZ0bV6oG0TOk8KcERKjIKqDbP4s6TOohBV6YibUUVhjtg3FY1XtD/HmOV2
wb4nnPoVh6YEK5CcJGKdvL/lUjC/jxRwhIsqtnrGzVw/Ut9zs5h3KDodwNbv3HVQ
bfgJ7LEnBKqBQxZaT6F4yKazkrUlvDbF31sBsNkJUzmFhM73ks4pllvoAc++KLEr
OQTEZPuTR4mDKeO8+tphok1Dxz/JekB9TmeAZRT4Ul9yX3m55HChNYX49IUxrxP0
g86thPBgWFgLournF1Tuq+QuPMadEcSycUg7AYrsrLKxQxICkfk1Yifzw+H+ajqt
QIsDsNGSb3V+nYPkyOja7ulFoP6OB3L98/3Ta9cGTn22MyZOmCBbGev3dDunLPZw
oyGQW0v8plVCLdtvY8mniT0F5lMjoOqeSCGCQ4e7YuNsxVJl6C+wYIONj4JPAJLW
1eMrOlIfWacitT7Uw2yHHIBaKvudLYIsoAMspAEJEIZX671+fxc1eEJ7paTA+yev
sJHBQPx4VUUlpuEKGXUeEs+ZWkzGfQeeVW664g4fWAi8wc/jylz24LG6yXLUc6TF
/KwxGvbi2ot0WfOiaHBINuJwBH0h3lQJUM0EIEKHQ9anPN8asw/PnEP4nr284uI1
zer2Ynvvpx+AmIQxQEvtU5l8624UkfnrC0NxgoeN21/xjO42KddddEztE1Y/P1O5
jotvb5nrj5WBzgsraTUxAa+Cqf+vNoBk2MtMWFy3dhBi8/alNzUpRAmXHBzhZ3fA
JBpKCY77znz8oK8p2TUartyDVU5ShKzoZdOJghWs7SsQhAAYJCpYmWIK3s5Trffe
2Ot35gBo925XQKoS5krcIX/3085yUOpkgYiuiScDBSx0QTHMMyqnv87drGXYooVP
toVcgg8btXlgwmyi7qabi84+QEuBZxx9ZTuysCaaa+5Nvyh4bwhUeDOQ1K/q4frd
fSD/RIMA6bxniVUUONyoUhxogv/8VwREhkzRWs4jt+ceeouUpZOrrvRlNFmK2zvk
U5xOjLkHXcKKiRjQ10tY8cNTWGFbWFB4pty5kMBuBxgovnTh0Rg2jA0Dn7YZMmhb
IqOqrO5t7VPLxXilNj/OyQuEfysee2F1FjVhtn3hPhCzlLVqhoKtxOIEPddz7Fn2
ejK1j3SizDANh1qEe5j/R+ojOCcM5/zk6K9fRqKdPeSoSzqV7qA+6i6YNmjT78Kr
Ex7/QF9Qpq/eeDMRsBQXqfDZj4p2hqxx938a+PTrwDQDAMnEnToe8x4Q7tzKfljF
I0dvY+2Vkc7yNto7CnbwruIx8ZVlEpDaMWJOTD4Q7mLvjS1BwWO3w5hpSFlU+sJT
B1c8v1YG6ZyfHGVxwE7+dTw9MOg4Mzj0m0AlYf5KProu71enRTYAtqGE8Hpvk+6U
bv0MuB5KZs/L7/lJ6xwbZwF8B49rJSd0+5OWxIpGJSvNMOJGV1sv18l6tA9Eauf7
zGfzHwz4bJjfuYDl3G3PlFDRhpHqrK+6VshquzfV4Z2gaGsUebRsoBCWIURZuOBB
WaXL/RaJM7rrDowSQ6GBzPuqVHsLZqUdb24Ugaxg1Vk28VQdHB++oeZK0xYeKTlx
CVRYhVpgwCz9yWtQX0UYFjb0lEyl9cvHar+mBA+HgyC/9dIAySG0fCqpspR/RQDU
qd1fFYp0XE3006l1QRYcXXfCueF234m9V2w+7SkBnH7Fqbgq44RP5CHfc1BSUm8J
AzelohlI8Z40xkQJh8Tt3rAKRbJsVXK4i9C7oK3QvfS6ptS1rbeVtHPH5EISpgBD
061BxhvsueATLIa/TQXpPka4fz9hfRddU1FVjaEpIAC6mXu5mW4SHc94cAcIyv5m
GsCRLsDDwSo4AbBYVdGudy4xicVW6vx8D+Z+xbIb3iaH7tJsYhBjhHZS0XTFHM9y
u771omuao1JlLJ/VLlKOk7xDnszPDpyMD9bdhzLmk+4ubS858OLnpxeUy0d9cn1l
z3oguSiq3ANpn3szbAj22ilOm9JqLh5pbfQbZ7WhaxyTooURcnnJxvMLW6A5elP5
DhHv9+CbQQ69k64oJokAYyAuo5eZDL7lLFMbuw0xSxdLWfmtr5JEmmJlbCxnH0/D
TnTzG/Ivj4u7iVcz0HcQq+qa8TsZukl08Rk8hWX1//2U3x5hi+jx4SFV4DT4PJQT
kmMGREQoQZZapBeN9sT34f6bQ6drEKANlvs2cf+6KlZTyySPZ2ALGDTAR1KBtJLL
Wn3yW/0Zss7ywM4cqq1g+MQxIsIk/m16g8Ehma1c4UkjUP/g4kHszD8Xk0GGmr3m
hTfHRVjlGMrgwjA90vvnJSYZI2vovjvDgmUKl/XTREO4VMVzW0nnERI3izyTcj1f
tP2SCeVHkt4EkxdCH7GgsY1PpcbNMCGmVj/cFvqnAJV7m982IHf4AZ+FMjfLxbyS
nW3DdWS8zDWctliOaTbPQ3XhL3END0EovEaMdr3Fh750ryf5HwtXZ1s7t9TDBh2q
nKtT0665i5bbonbs8H4ee01zaRMRz0w75cE1UAPTw7Gc4552jrc9mnVKWDQij8yK
A4/JBgxKqbf0S2WDcPitnc5mCCXda851JDhzuDtXM55UgDSUlNT3JpFARDhzGJYx
aQBcNfiQkXH5IiiWnU4c0WRju9730N3KTCK5EkMSFFIrgEsWxc2ixszntkvTZ4fX
sqvLh4qyu2LN1Gse/h3rW3Ctpsk49C6M89rrOd7wMM+eKX3Qiz2C4cFTFjle7XYv
RFu/xENR8EBrhfvAb51x3A0fGWd3oJs/6Aaq4wNfA/fEF3/yOkLUQtAbhxFe+3r0
nKrifqyuTZgEDzUouQXPyfc94ug8UBGyZD++mwTEQW8hbouosGXJhLZN5/5dvRNR
/hiUXNaNcefL1nPm9QMLGzk3PLPb13I3VSdwdzpp1wfrWcSTU9aaWkhxy5Xy6A21
cut/k/HnsZKlk3ZA9iFGUp5llkp4Gw21p/PfgmjJ02ETzlyYGSVZkTEHPX+7BxTf
Fgo3WX8pLmY0sAUx28pprPAU87BUZBxC9hb1h9RHtANsuNRd2w0fHVYlUDSrCdV1
xWAtHlvMaiDG4Pl4ovv6TxUIFxX+uD7lVwlkQAcTAWv4Wxbg1lkHfMdU/JyJhGKH
dZcPf0e56qOUCKQEiAKuIwEHV0E14lLAyRzZWjlyc3G6cF5EbsgrFVZQ1xnB04NI
2JOhvUvbDa4tD5eT17+kvf3/qQusjpylre4aRjgVmXn6UT7BQ1T4WQsKrPv9LT+o
3qE1lriVBRq3E2J20mVej4iaTzXRxi7jOphVRH+ZzL355/bl+dK3uF0lLcYsUScD
7guGGoCfKXcTVy2dxLxyTyxdG+2cB0FGO+klZQ//VMaJ8I62PL91XaEqHgcdUSF1
StDxTszlohQVi0ToSsMEg8h2QjSQ1GBJTr0aj8tJoA6VNSmWa7A4cHig6jCSqsqC
RZgg0xhmsnHyzLb2VrqDMePCv9aMW7pcQ5NSoWQ6UOMLPfk0f7zA8qRcfWrmdRjW
LA+XzS71T+KQMtMGo+3SU4r/DWXl5/hN2pP7pnwNl2iEV5iHmHZ77yFH4uPgs9L5
qjVPL2WFQK7yDLWhVoSs0Euckg/INu2sQR+VTM/fiCSKKE22jiUnVGWvaQCh7Der
A5KuPwVu4MQgTq6SNfzlyXvKl701tD0NZvB0y5/eMDnqSz6eBiG//FoCWxBBEPgu
d6dGWeBJFh4ngHUGNp0nbvH4OO5h+6Kra4AThOkKmSP0B+6pkh7JSP1F6J+69xWu
LFJZz1yFWiqn+po458FdE5BkveF2GfWK+1Ieh8nPgksCkaLrDw6cXD03dplM6MSh
oQzfetMqG/7LcNx9Bpp0ocfffG4x7LE+iNLSlBJX/WDRqNPENzlqcQTVTJ7oNjxG
eVJbY9UT3C1dTLAqR41PkCm39k6YaDMZxSRuz9TujZ3GOkDhJKsIitt+bJI3T1+R
tsgueUciRNlmSCz3hN0palMAVh0dWX/bVtL3yM33A6JcoOkkT0tfD6pbh1ZbiCNk
0CZSU3oJ7IB+1anfTObeFzksoSNXJ4S7Ax0WLu0XyM60ZIpGoioh6RK++P5ptlff
ZcjNJVkrvcCl7f2LHtAiLEn9/rHu5C2BgO3lj6+L0F0viK0cRsZYsXPBjAPLQOcy
wQT56qFd61E/PpSH7AE7gC749ulyIpO8pqOdXSfnQlPcYUXBlZFP6yafaaHZu8/m
aBIAHYVsE/9UCPS/l2aYdeQu75K1dHDLstJyqJ2ZlXQCin6lyVrQc8sahx4AxKzi
hR5T5pZM5WzjsauEMwPdCH3c4LnWbnBEHsEMFQ5VRgcJYEfjw6USuceZ69luyUo9
WA3u/b2lpTLUAuznYlLmBrnWT/EB/VfOQVF93OeLgEGcuFEDnv4Y5eakEuvMsDMq
hsO79JMWo0dFZVk+KV17FhH5Jyh9786LkQb2pwE/qqCppX+MQqRKfauoxtEqIXlW
vJC39nF0G+3vsJZzDYeeOJWJ4KIHkKv/4K3gAJOVAKR3bCu8EApyktjUJY6pUZA8
agPodhi9vabNSHk+ZqtmrGJdVnc6wbf51KHOcDuRVAeWBmi71P7U7Mzdmvj7fRUC
3fH3OsgAGHseu6uBnEpHpXDj+BSAvxrBrYhQNXsTnLqgDxmKd56cjxYoDsJBPYSt
WfRd3UlSD1Cq8cUQU0C4KF9Rq38DEWmpWPxeru6O4CKcepBJi8JrVFPCE/XJ8z5H
a33pyFU+yE9Wv/9LCC2I2aub+VuyWJx1ZGSgoW7OAlrQYBOnC+3e96k2MmeP1Mr5
cK5/oPsG6yr2tKqfP7QJ11Cyd5ZWgxRpjz0Wzaf3XO5odcaxt34eyykBX98iIZeJ
y/0dR0Ollz9C6pEZxgrBo6/iGqtvKs6UxaHmzqq6/kNdrGos9+RfnDNB9zzL2Pax
yz/Rkujv6IdgrxRtbqzLwZFy1aiqrqoC4NTclAIr7KfkAqmCj7IgNMTZ27IKN+xI
og+M70YCqr/PQsemPyH/GsM24H+wab9GBdJJ/mbOKaLLxcBecqYfQ3v14zPMS/Dq
FsbuJywQCKlR3f66JkI7C+CmkVM9evahVou5A6+1Xy39Sg9G+o8/TZleIEjfLKyo
VUdMRtsoPNMrrfcS1edCY/haEwg/FFzbDCdEcSoH1hyShZPzvK94QAnB00TCx3so
FosrtkYEHlfT90VluO5HjjfTacA+/vxx3n28FF4ISilLSrN/SMwoKIG9ivlv13js
+C2LOdiD+3Lf1hWOTwFeH3E2h4JBpEefyRdhIDpC0yIM/P3qNeNb4jUwMcCzbz0p
yeRjUiFmxv5FrMIqtyoAC7B6UKRSQOAWSjMYY5xwYFlc2ljy6x6tfOnOHYWSQ3oC
C0NUMd5XTnieAWeFdUx1ILbjgFJ0DNNp20kHce5VLr4BRFcLBr4sTODbsHBeVYlC
3lVz075JiD0bsG/fwt6booRtIHinJ1IcCyRs+AZxROyljpzwiu/sSnOrj5VYhIok
06kOv49lgQ3JPdpwkpVxyQJ7fngzcqZ8cPrGptQUt29kert14Aunvn3YvRarX+py
yC7shSrj4u7WwM4nyEHSF5cJ3t208Cyndtgl5zH4WovSZBMO1VTvMubMD5Yce1CC
em/alqNKzWD/bpPAGbhw0RFzLb629+fDdIlfefXIfJx7RxSroi/cVG5v9woaQmdl
whM+vZ4DL5m+V+ImknCLIfZvWLsbIsi2ASh1kuUqRR5T9aSNSWTrVeZuCYCMwnN6
oB31SKKQiysPxp8Wys7kk+dmRbKGtkPXcvnvC30CBjspSUE2BBUd3aVcQ9n2D6BQ
jXJiojQ0uqoarUzDvJUUffmcmUnhwaZdcMaxRFDOJtQo9fBnW7Pzv67QrkhchwLM
ZmUZ1J+5LV/zpTr2VGuiW52go/3yIgSjwTWjQ0vbexiX3ptDbOO9+npWZzkyKrqJ
xhNfoUNAznXM24bQFE7GioUKImMKC5HM/tgQKrpyWEf5aJ8K1fJ5WrYRz0LJXf1a
4CsO744Ivtk7havrWCCZQnQUVWngipWy0xYVSZfWMWP57sWKxvNm7PWTPILVrCV1
hc8NC5KMrZOYzIOKwamiYPUiecZelpVNLkdTIJT8HEpROvG0OcEmFccvTCQnJqYI
9+ejB+suRg1kldYl5KJStTRTeSZ2BKSCVimU7sL+jIEMjAm60eBLylxcpZZVNZ4E
p9A13jbEc0LPhakZtnTixidbMEfP32Fazo3rkCpOUV1ZJnJQKUDYJfL3+jDphggP
lHTQBTOil+Pp8IMjemg0Iqejb3O+s9P32tIm9RAQpqhD7XT8ZdVsDIG/gkfeHL8k
dz2ZlFc+uWVOuWJ//WN3MKxecX8TQQdd28AT6EJua2tC2CIIlV0Uyi6VglHAUv14
3lwhLL8a0H/orWGUonAUrVLhLVg+psIZZxK6S9MlmWNNWnq6Zf73I1saf9N5o7NT
dnOL0rGXIOyB+0IVHOj5qfAxFbeGiOPhL0x3WZ2g44RCzzBNJJmmNK51AIA3t9IT
P7SINtHjkE6sMs6hSjIxjclPNAjpNfJk/t7pdK6PUF3SAzWcq0RD09JYnUTkTufF
g0Yui5/agqBegL62uURZf+yqG4NFIfJEqa6Rp9wJ+dILiAO4J323lwS1WOFkV/Q8
XYE6VR00KaiXjz2spI4FxcJNdJ9kbZ8CDp6pLbS6uCjOpz/QBIEiUJpSclJPFvTR
lAomWTVPu06SB/knewBEWI8/T7kaDhtOSVlJ26t8PKKod3q8O6XcaYRk1ihrp8mf
h6xRPKp3A24yrPu5pP7dxhoJ/fP1fTpaMp5f75JSPY5iIsufCZ1P95C7DE+qbnc1
vqGYyab+wjYua17Ef3C5YOXfWleQ0nc7Ba+p6UAe2HLD+1wHBbtwnOnpLj+0FGlP
AzVm9irvf3omRuLpm59sa4I+6qQWnqQyW/yeayTXwWIxzWX7zyDLCw6SxkE9VMLM
HyHXKc6hl1dIF9cL/Y7scRH1q2q+juaFKJppG+IQ+2VDpsOWhmTgdTDj+5HMlkrG
Y7q3F5GmUXs/XxF85RVFYRxLG0kVMwvd0s+Dj1Y8nhkM3XxGZX7azPVhFQr5IWqC
mKLqA38RWjX4jgC4u9Yx1CsTa0uU58NjKK2TjD9PJfHz7ObfaGO7r1uj8Cwry9GW
xkohYu2BhQwsJFI1AxCFvv20ingggeVQPZv3Of7FBIGXRfmlusbQt2zZhDzzcHY/
7OT8SSm6POJx3cbjG07nZRknmvQW9udBcqS2XNYZIjbCeGrZ9jHoNzagNfkp4SfB
S3vke4OiBr6pn0JPVub0/yR4ZNffuClXvUJh87qbnLG2O7SrCffTeJ5NBKEX9XvZ
pr/sq0xxZ6tZhZ3R+D80/YsXtidybRodBCj6GpFpEhAMVqSRPHM3A9ZWy2cn9joo
6p3Z2Qc2p9+3aK4Nk7qAAuB+Qjy6+V3Rg7rH5hvBHs4LTiDlB7q9e3wGpvkljPpE
YZe3iKrF+o1MRZ/fzHuuPWQ2lWUyn0sptvtxCHcxXNh9YES/Ikd8DuTQiJ37qImv
cfiL5KZ1X6gH+RUarelleJGhd0L/zugqA8GFR7lTf4CRwsKH+wL64FMLzXY/tsFg
84IwoCmxXKVoyLSrzg/b8kd4WP1hgSKER4ZIgbH0Dj3u+iyEIUNARkl1bbggn4IC
4uYHTRYnQkGE8rY1hobYwzmJq3OI1pNEzLynY6BPpFyRh6Pk4KFqR1n5tKYb+oeX
A1R7teCuaxj3DB3Qnmtov0IgOsQM/XIyWRPuoAX0NpuyEFCT1jYIXHd3jTysIeDS
Vpz5FHyg1xcLbLYXIJMq9mz4YsfplDWUGsWG5aZFi21IAoNMZdWyxJEuPm41stQ1
501MTpPPitUNGKw5KS3IBwAyUgCJxpxrO9/hmyi3JOdI81OS0xgwCJ+ZS2P1nNru
irAzZsh8aSN/2MXGuXS5RAxkUd4ZPtjiRl7/3JNCp84xAUXTz6ThcUepJoy7flhI
AemUK/GLywy3NkHRGsxMfNnBlCvMuP5KmjzUPLAVc8X8wZFY1b0ErSt5V6rKp6uC
FuMJs200NAAEMOmmxPc6UKheUg+v6KVQGpNMR4gt0PeX79dLBNiBKs02YiFoFHOi
+d3uf3XjqiXff5/qvhKNSsJbtDVTUFigKlGhSeteXm/Kf5UhzAj6OG/Dci1EtrDQ
GzQl7QPoD+1XNHmkkDZ/pgqMjKkZl2TT3G5XzbpZ4ufo4HF/qFcb8PPEELpSuCD6
N4oRxocKNEPPBFPKPv+ocmB8JSNtvIZ2a9mb3CPrjaUI5sOXkOdYrnXCOf/6ghUd
bI6eNMab4g0/OjpCiqwmqIzAwuqA8pnD1wI99pwEFu2f0SQEn9oACoV1YWux42Tu
kJa7nt06EdPrn/LvEeYjYDh8+NMJphn05KIdMJFliYSjgxw7Vw/3QxCg4eH1U+WN
QLwQ3+d9a7ruahAKvDD4yOBo6UFjge4Gxl5HEjTa/rJmvJkfRETUst0SOiGaPQIF
aNNP29PmT+P7nWrPoY9+ZG+4zIPjOZGlTPQnKmvtnyNexI9oEf13sAFaa2Pap9C9
KuiECps1Spn9h28ulUI1IPw6HOG0pfsiwZfM6YaKBmrXnUaAhYcpCHZxkZCjk2q0
jZbT4ncKL8QMGWo8MPfs+bQvgLnRKLVY13yczDh1o87PZfoWE/3KW79zEecaL/wr
iPv2g0aliC40DgHkMeYTd2vPPZREMc4QwBEtvGSpBtwlGe85Ghm/hTxq/k8Ekwa9
GO/+Exl5yRl5oYm8IFqlQJYCYTlJDUFYcpAODmIgvxfD6oTEvzpIy0JJLsYF/chL
B24XAUAezcx4Qvvb33zJ8XFK9OhDthRz/S3oK6pWoRX3n7hhp5I1pLpcaCFj2U8v
PI9ZoBIES5jrMhNHpcuQv33FxtA7N5BLHeb352Bnn2AZk4xCW127xxVdFYovndO5
ZCOR4mJTWnMmgNRWw1XHK1pXFUxia6zbYL4OHZVw6RGZbYQ5p49H1uT3wCiQBVXq
jWnvD6jITyxFrEMsyrPl6UfVOul0E9/N5n/G+xKIoQ4lQosc8QFFSFcplLbW0EVE
xNzMTbqRuc6ZNahCVffozHw5Wc+XqxG+cRKtGmmPZ5c5RgiVvxtDVTm2MF4d+SWe
bLS8tEemW+MqmnF5D3mU6lxrh3hvIJij56DTLFslNAjAU466PkkEL47o568RjzGg
zu7uy36OaX0bnkRZY61dDYMqHpLLxrQeayJlfJA04pc3qy4nJRkRQakGDx0l+NEw
i8EI4D2w46JyGso8sRKHm95xKvnj+T9dlLuavAknaLDyfKAdThet3f06sE73K4Hc
LgOYLcohJ6ZwOur/i/yFUkP8i+0GFsh9EFP4Z4ngzUUoQs9UVUxwJBXaBe2zTStM
A+Wd5TDPv97duTsznW3x9Wm01g8RY2Ak9hi/we4zsw3NUs6/PmWGY6DLnCuRmB2I
CdbAhM5GMJ8Wksk8jcr4c+Lqyu/iv3fUDDUwLaiUhY6lbvbtW2e8ARLn01Krz0Sv
ZUaaed1HLp8ZroFy1uu9E3Q5MjROLKKxbvBqqE0XcvLD+zn+ZxFQ8uAHNCQKLtf4
+tuTPj9UeoyndJqSYsDSgPYIlwcHL5bzkEUcp4zg3d1fGIqya3IPA1xpkMEI7b04
c5Fw4Xff5dZLXaRWjEE/QDivTo+bzxzBoaOJV3c/VC2Mvdo/2UV4cfGzzm+R/BhP
WdjVmWlZkFqYNeVaT+zhN5DKpYtFZVb/0PGatAdBPCRpEcByeoM3QqweKV5J3jZR
Ka3jvK0U0IBYmbdBj3XjaaQX3gUdk3Y/vPts6guT48iGV0mpt1PPAYVWISX5l5gk
RDdToeRuUuKsdP2Dsa5ONBRR/6kTeijHWcx1TmXx3auOTqTtQnraiWO95JwlJgVM
poFSlEfshCljwnoA+OxcDH74y8g84+cbMJPK1mQ5MLQZSaJlvPY77Kl4zR88rmZO
3cLCXX6+ZSqpzOG6o8G1X/dg4DWEHOLRW9m3BF5i54whdUL0J2B2RnqbTLOVn+Kh
uJq2fQl8bHhQqJxYOwZr+OHB3gR451gEpvCoJXCYJCQPxyu9Hifgi0RwcNKW14xP
jWTu1brmnvAd37hnl3udchX5pz+RjbJM9VDwearS1iVs0lPV1spCc5FAXLZfuvaG
+p3TRxVwLrxvH9SR0eX0Et3hLzWUeO6rcSmlgqi3E+B7KEAkvRAt9rncU02QX+mQ
bhPtKpXmFvwGaFTENrQVOjNwL9Nvw87oYre5X8LbpZa2WG/QJMPTplUwNpnCgH55
GxCGP1Tf/lyapekBvBGqka/tEf43NQKXhp8SVIDcQAkEM09VIZkvPe+VzRxvT3q2
CsubV0Cff5y6Ez09xZPOHMU+SCvuB5lviaGmoU+gZQjKvKodWMkXnQZj+KzhAOvt
dcYKd56HkR6Scpy0b2B3dUEE4d+Nie7ou0jDhvf/FjhKhogZShVgizoUpe/rrfme
iqgFzUl8K6gk958jcx+p41uTMriNkHFHmK6GRuQnAn4esUd9OInI51zLc7LiQwJi
t4JeCn2U5yb/TFve1b76gfMSPxKsoXQB+0wbNZRRs/gnML9N58/DG383kjbI1uC6
38Vc4m6MF+kMiG2gY3PDL3NOqhztEqjvLySl65SKDb0svokCElFmwqiUAa5+gto/
VPT4YC/KTh3aADwA9x3HG5YH5609ov70dU1zhu/6nEuQaodRpVSrRfcucAyiUvpg
vXYxnbeMbpOioDxUvXI/hegj3YEpRZtDNCGMu6wzZYC0jdW/KI2tajnUxEyGoMAy
6SobU5qnVPqsZa/fgG/HZBs1RWNeFLRsCMD1xH1rfDrOnY73zH2i3UtCexlw6xYw
Lq8GJPycokKijvWC3toSpqDGe/SW5AYMLgB2hLs6FHFzMqs4gioCzua8FxEmKVUU
MN5O1NHYzZvZzykhwC2V+1tiLFKVjWQZLIkQYjQSojTQiA1LgpI4pxN8+y2jvrcI
J0RhidgW0yqSMrJKqF79m2Eho/snXG8ET4iI94eVBGNMQ+wWYLhZbp349iUjFhYX
cpnDrZ6cGINwBPJprhp25d3tN3sxtgxgtFVWkT5tUgHebjC2aixqgnwJabrULzrV
8CxKtleo8PhjIZW/LdWli1Wn7D8ecvOgmeJOV2PyllbCNRnB+GPY2qxFNihOtanT
3tprCgzV4fk7A3LKlwzOD0zy0zVFhM05b7KesZFtPf7AnmTSCLC1d+sV5WVQGjBI
yVL6M+FmrrxAaTlgjRKVV7ZzSWIn/XzstT4TH/gERS2sLN/GbPMCdsmbypEP1b+4
mWx8frNyC+xLobpjOLOODW7L6k/ukk7BaZMwDOX10ZdZwki02ie47FKuooKCDPSm
9tJpId2Id1Vmg19TEysKU7fdX9jteEQTyqbUrd5QMogFroVtHplh/2TYCx9FpKOe
yy9ZlOnQFL6bpBvwb9RQ9cCO7nxZLHS13ZE3jrfNig9/yjurfUPSdplU4x5uC3bp
pxrAlgc2tkIa+xgdKCDyGTr1q4mTqh6hKrpYA7H29UyMFjXb2CYBHvj05ITmPW3l
flQdTjbeCrmKWNLAFkzvKap3DGAeacnSGPTyvdrGHWzQWwK236jOValFXe/aQ/d7
FKMeTGNO3zG/9XWDpsWzkP5QV+rJNpPMQ6Z0bBMnVuYzKKUiGz1EO9xpim14rlkJ
jtoFPE0S+hsaFqhpdByDrGdru8o+GexUdfOz5PDC5LxTdLtdc8mJtznPr/2vinhL
3llY2ZYBxr+6doCOq5xp3pLdvjZ2xCdpFQ2E7RFAylC6GCYvV/psD3rLxQD4WXMX
rERUjfEjTXRrnKWGklPkXTAum7oDDRz4g08aW8Mzf5DMMxyOV/WL1T0YG7g3LEne
LC0UT3XY5Tn6s1Ube+GFrxyUuEaTXG9S8bQJlUTcBIIc45XsM/tO1Kjots9RDZb1
ccymsTNTDI7hTokokPcm82FhhrGHXHhZxO6rvum5ZNF3wt7SjTE0AN0ayNd0sjex
mLsDqYUjtB6FJ65BW9aDj6JypE4BgBH8L6HxZk1jeoRYtCeQ7o5+JwQQ6awp1QLZ
qNuT6JWVJQyaymqXmGZI7VtZsGdMpRTaAs4XY6GpkKnbNeOge72Z3oMqGzPf0Fdm
1mbJIYf7SqICFsZ11BUo4rKnOi/OafDwTNTFViBxTLV0cOTEcXJ8RSMYGaKLCAwh
dFSg5TW/1/z2NLMOMXTflyPfaoD/yNYyTkUbI7d6eC70zA2Yz8fwjGJxLTxzl+iM
UxcBzkagb8Mx1x9mKlBfbz4VK3BWIqrN0c9mWc21d+POjNrB/kXQBJWt8gA7d4tQ
owpdzO+GmKx61ZKFVeP4FRE+eVDzqiYDfv7yGPLD/Dw6IGn4qWWeXM/3ZLZIjsoz
KE3HaixdPSDh2HzesaYA4hYiBNO0SpX9t+wp0t9OCG5eSGfWN6H9bsmvOCxszf5+
2T8k33r0MUwvM8Yjh8+TQQQGpaFb3gj5HlCnyLfUl1XoXPZtuKj0VFzwboIcdUV5
Y1+wfDUZmrtDloae0bp/TNXHcgHjYg8rh1KV+MH2CSALufzkB9Zziw6kbBs7O1Ju
T103Y22bh2dnKTlYOI9DEGSKfmSblHBNz/XbLtkTi2vxvDOZ//EVgg2Np8hUVzJK
3vWfdJxfHddczowz6yqN4nZwfTcoDOo6Hm9+/GTO3dj29HYjHC2N9rAHJjQ8EY0K
sfgBKKQROy/F/VpMmLQ5VNYBoXYhPWUGUduwDDTJUK3rdsKXMjzANDigmQZkl2lj
BapCIoPR9bSV3En/5IQX52bUXT5BiKsEqOonRB5FDckug0cZ5rUP7UEBSCheprbZ
dlKfyrPEIlMP7ZUeOGPZfgVAaYyTdRboLhN5j1s1Cy8aIOy8z3kWvh0tDoULIO07
0ZPh1t8CZe760IM+zpPQKUrv9cNboKjGQKOEeqR6OClMLlDnZa0W3Tm3xXrwZo8q
ckpo8yAVL6wOylZk4+Gwq8G5ybgKBkQ/opU/SG4L0INWdzPTNfemhcFwn8ew2+3H
EhmHcGH/waX3rLauP3whta8T9yuxo7XVN/FAXEvN0oByL/gT4NvK7fp8ChM23Rjt
DOupsYOXsbgNMLr3+3iUnl6HPRGWjui2ZZdxjhOjRmimAvYNY864xmJWNi8CWpes
AsEMjRmhw8eIy7q8WiqGxcAJYNx29w/JvLG7f1liMzpJDDBYSLgKdIRgLIOc741u
pPPBjyZUdNi0kEhc1moUWWkgIgWulC8A9dq45VMx5Au+RCAyjKruDiMDjw7uZAmj
iWDBVq3Lr/Mvvzf2XqBVGflHyMwu7ScsHhEqDSnVn7vz+LyQIb8UipqMnkaZDwzM
Hwh2NO3vP+Cx5BOxPbm4fE2U0n07DeiPeFkYnVakO07CC2wf8FhfqViOToiNOHd4
6/dWxJonvQ+taAwgUyQiTjs4yOrU8sPDs5fBgsoLNrxnDCOEofP1UfETzDsX/pqd
AK+F5AMHEp4jpC/Y1U1FHvaXnHXHjOjBLH4oC1t44r+v0eW8VsWH2i23EiyiXzt6
3M839qQSLF3X0X7qomwd0y3v8OCdGAbslCH8QQRJMT55kD2ttQOkYbldx8JGAx2p
+/HxWhjJv3zBa9psR2RFaluNsyr5fkohIXj8miJYNacgWzQNui/5zKFivxHHnGFE
GEkQrOqrXPo6+YJxW0ucarVVaHEFbiJGIAqrPVB1+OKjs+2eAWI3M4rcbnQkat2d
i/5ECY0lH/8BDx7737wdb/zrRvriZXfixudbuf3Qei8/prTPyBRs6GsALbhAtncN
YNSqmjqcm+WSDfmK0FuA3dsxdayfFLJlX15hdXEUq2DORKC/A8NFct46/mLwnXBk
I/wgTXnyI5n+dKN4NKkV0Mc36Bu5Yc5IQP+s+DL3ikGiiabh9+OsdlsBzDM4NbSz
0saeMGVikpGoejNTU//R+bCsAnacjmACutN5VBU0isJZyrRDmYhhM3aSXiGt0Luw
1x+bAJFPZWS1w9a/ccWd/UbC0oGMXrU/zbXzE4UMJ2SbeKHj1Ey+3vGoKhhYkWRG
KC7kAoB4fUAjZwxqduy1uLOi3LaO1XKr+YloxGWBjcDdMSjHTB5L/nIc5HC3oWV1
h3cVZCpSBSpl62nCudweUmJa+VYH1d11GbXhwSoZaHJsOZWVunKRYB+Z4I7DYo2D
RSE+5DA24gIfZQWOQ5R8rVIfk7T5iDEtJ+FTFK8/RbnNitApvSmuBIMaGvfMOQYq
IHk4Ab05Zl+OUbuLca7d5moyUaSGeWK99PZMX2NCxerLpV0CpaS9jx5YtCeHXomR
kffSXS6M4Cx4BHjpTdndvojf6yBNI5cdGJJU/MFs7uqqEe7GCtqtF8TPhzEJ07f4
fbNeYyd/lXf3O70RRFLOm1hppDhmuxo78jp4Qr6/wel/I814mXrvsn2N/VCJY7TU
WXlqmRzsqTlxTv3YOQ2HfBOipGjF+mSdr9vEE9jwnafskNXH30PFjvBans8nXQSU
z8EMJ64QGFcA6XVVRggWGh7dTaEGnPi/UqJioPKYkTmBujSd+ckGuubQQ3LplJ1+
xzs9EcFAoKcY7ctKUe3VL7C6PbF8ueUm4X6Oh7Lxzn2NTIkpzjCY6E41220v7bvD
8KYn36xJ8hODc5mvtPB8iUadNEdNgpL2QtPCYAjdn1Go5XtRJVfkELKxXHYHHswP
9HOP55NFdneC/3VrWm/Ur0tAamGdDHa4Lpw1u3Cas1vl2UPIf2XXVsQto9XKeZ0n
anstzBfE40HiuYSOlBbYyAPYmAhdJfT2qi31TTaTyxD4rl5IS5RqbYjJvA0bwVT6
hr2nbnpygXbNAxTrqI06kOvcapoVSyfTv3ovbxrLh1gbohjcxjdqcIxh2fGV483T
Ta0cLE1PJngjhE/fz+PM+74z1a+IwRQHbjKXb3aAiOlgh0RgoRWOAjs5521fxXTp
jGPXyq/7LIflaElbYakTyvVGbkk83o1BEFpzJ1W+Hh+Q4RKCrPKP5nLvjLL2tg8y
fFcv+3BVs6adMllVh82eL4YST4xWVYqQIAMAOxB7m5Z8sVdwqKdIIZRGvTPyUrgi
NguoR98NGFArhVngtjtL8/yrfS8p3IGApl99Kq4rHKBGLCGMiwsDiMGKlF/9BNiE
zydgUs/Zyt5iQ/KWidUFJfe8fP0EuZ/7wisUP7sXy226J/S2p6q/PHufEUjCTx2O
TlKXYUxDiMaKEqNudTBGIIvpEutgWcDS71CYWPlZCoNXqAzyZHQMt/GI2pCfK9Yl
Eah8/eCwt3fIDRlRGoVef0gqOLIqaGrwQ9neTWRMjxV51sRRcxFwFdrroe3MMqhE
C7cnlULjodXEBSMzLJQZGADG1PapPkIim9Hs0HYeAZeooK+Pg6rnAAn/eMh2LDtP
Da0iUwGk1D3YWQjcLR8hTXsBI8ukzI1glWs4x8BOlj3k0BHQhuX0r6Nzn1LwseKg
1qGBEHAMavDEAig5djfVfhbFJCfFcxUsurO+vuOtOnFf5mxVvUdt1SauKguDJxIA
J8k2pbsW180BSQVLOriihCuWOAVJIyaDu8pBNMzV3i8sIlc/wjjunZnDYR7adgSO
oXAlxDHX0QUoIXjnZiCPNMcTTiNszyd/jR/ocMXjUwIfflh797nGo0REABWaCi5L
4m1zrTIEfcn4e2YbmcaHzBpakPoM4CZ/ECIhBn89aE9Kj5+qO0MXdU+r30o+mSxH
wdv/E0QA3mugvkq794eIYBo/FWMLtJMgNfsGsZ2ahtRUYLbzCK5BPbpxRRbRXxA8
1s7NMFeeBrSxB9Vilq6LplwBZeUULn5GhDBRkrBa5SGvMVK4JTpurqtVxU+RGADP
QV7rSBcTmDdRn1x4wE5QP7HEekHmQNyrg+sZzw5Q5V8EFMxv8X4ijOo/SN4b0jwO
rK0J/rSqU8nhexFMj4WR4NDWkFTy0jl/p+QDopR3gc+OmzVec5oTBkJuYhQ+G9uy
JNR5XI77awQ2W5jF05ab9yMwU++oHcfI/F/fLVx0GhgHqWoSTsS8ZzN71TvlfLNs
pA2zTiR2vRS6vUjo2dHAEvAdXiwn2fZLvJVgSv5xYzsjWtOGsEKc2aYD0cS5cbLp
mbEG2qVENPh914D4Wp7gc3Q4j0j9voWGMehF6i2pIgGMUSkTF271SzGuUIKUweib
GHGr4NEy9JUzaVWF1MzXYqkK8BQVxOT57xhSioC2pzlJrr7zfSomX/KHnI4S3QwF
zMOxNAeIE62gYgrBSzVqaMk5WC9mj4FxYjnPQpXFz/3L0qLGNERqplmaH+yeQtT6
cfyUWOP6pIXb2U5N7JovsI2eyG1EH3wSEW/b41JHDByfWviNCPQ98204+xpCIn8v
8K92IVHPkIymmXw+sp31Pvz0sSNTS+o+YVjmEinirwg0Dj1FTFJ69S67EuWnUubY
hXWLiA6/PpcxWaxFCIsEFYFkQ0931+wBCat1Z8NAaYeiTGCW75GCQM6uFUzgLukb
CsKRfkBLyItO7d38N3VnOp2FJlUTpQGr8Xb+bxc6NBGXv1SlFfezl1El4VGaABbU
+P1OsIRcsWOZWyvZCMG1rbDkNu9ZdWgbESp5P9srRHDc1ztv35ltI+SmlLtKhjqK
NwpJU5tuJ/tQQDYFvpR3wvqh75OF81NqMcQRM0EvsPO3xZx8OY6l0D4jJIysRmWQ
aFRo9NOAfKNx3GCUctrV5W/9MZThM4hzWoxPiDa7VQn5WqUG9lKw8NxDbs9nFFnc
noPbLny0KvH/QBHfcdsO0SnGyyD1TM7SHd0TKKheTc2ahBz8LzHP1hCDpZqA/Q5p
H+z7yyU+tqMjC14pir3oLowU2OZh17kl/rEtUNBiztDVYrMDvRhLF7nbGgCr4TjO
sOsI4kiYhvj7o9YHKXEVL+7qky1xTAKMxlw+l0lWzsPdURG7LceUy0JrBiaGcnkt
2K2fGKG5xMnnD8gysRo0apo/kk/6NoUekjyMGNdrMj/eql/TL8XYUiwYAqeZ1W0b
5yfzbYBJ8d3FQKCKSasaTG8yc5tvyxuOCub/kDkF9BajmXFfTtptL7Zm3dEHLE0F
CLBg/ISXZlh9T0AfFbTNoK9T9ojCa1pLjNQBr2uYcGoY3qL+xuz54qXHGgEw/efC
jnosCj2ktCXuvlM9ZFFpDCDA9oaJAkI9DVw0jcNe6KQtHWVmBPrXfxJ76j1+IQFQ
VvnoLjreMNgxIZXJKt6r6LPJz4eYGKgcHGhR+d4B6EdrsZjnILfAk8t9q0NnZzrO
GB3WhsKJC41yvih2zLKrcqkn7MjB2ojhi73ELBfpqOB94NN+uJsqJ2aZwCczw3Kz
7rzpOFU//Pa1ERX6hus8N1yyBrMatQQGOyG695ZA3tgN7A5rhW4MWf9UvECHQOH0
wR7LJuVAEnBo4TSEKKGDSpJDPEnJOWZtoiUIc6olOr8zhi2IfYdnkPOOkqAktagw
koUznxpSpMi/uwPAMH6Qv1mq+qd7uigY/8XdkxDxy2t8dxZrG/TAXhiH3Ff4xepu
N5wPZZ4G/qFJApV26maGLzaW/m4nCkEgvfyL5hjmOhjX8lZDf3UM1o17qgp4Mdlt
2PwMm7HbFgjF3i3vqtN3BibZffAHdMQLee2w9Ccu14cyjAb0XNEXhnfbsY65KqM8
16r5YIuaN0c/OnAj6ZVcatggDdDhX9xN4O1Tvj5/jRSxCxGieiCxoP2vzaj4pzjV
xA2L0llyw0a9RnWkfini0vXDZK4RGwGzUbeNeAoxYZ1ls3UPe9fJC9+mipPHlDzt
tD7ph/rkqUDIaHNthMrsXRliHx1VY0upPQTEF0AvvtAn/OpdDH1XI4rUbyCy820b
tLPk5gM5yFw28P+s2x566iSHep7LSgw7O5eeS+VMBsk3cQvXrayiy6Gtaeb0PaRU
G263jj3vcIs7SV/ckYjWtSp1P0tf5PYDLqlgFwiWwW+HP8DSvlitEqTEhl/hczW9
542m7HxJ2weJYBR1Iup/r6eZHSbb77xVmUdP/3vyYOD2mSOIYef8hT9ODPJneQV8
WuO8e8emsLVpJauoyEA7v9Bf0M3MUhWP9/+VA6M5zm705OqWSsN4jKfOaMiZIhlb
S3vxQ8lvDr/WYtLrYmgOzI8x/rLxYR9TkMhBvK8gJ3v+tS55HnY3mZnXwfb/F+dy
CTlLeK6iAYYvNfH9crggJaOJC7uSh+DEp9z/0BjG83FHo45il08Yq8dReRHYm1ER
fmEEZXAWA8A3ht5TxBVjU1+br4bJrFmITpD5MhRFPYko7vzLKlK342LqA/75wmx0
1AOY2EDhJ+fL3uswjJ3WO2FPzxCDqeUKR9pBp7NDfG7IvGT4QucS0qPGgj4zGrQZ
aOjMwnACoP65s9Vov1jmde6mgqgqPtX5bOp7FmrzFaH9d4cmLyxFOj5+cqiZHrT9
j7S8JbBVZv6+2ShAZsHzqs1EYI+a6FFVnNt5lw8MwKiT1qTIPuAsmbM8rZOD8yq+
W3BU3mu2NG7PNVztZFkeyAcD6LY9jic8XxlMAY9Cs0XdKZd1Ol73KRpJKWNsRdOY
9oZCu3FIS2eQLsyCpNuk3cGFzfA/KLa8xMszFNXx+aXbSdIiAiToGfYPB/XXeF9n
Nk+Bc4HypZdnmlvuA3H1CwkdNZb8vGjkPe+mUAClv7d+BYTvFak+3BE6amB/oNp9
KA0cdkTi2zU5G5b2fRs0vP5Rb6/BeJ4dy7e4SEW+JKK0Wu4XjylKqL0bEoCpmps8
neoJakuYTxkeV+RJs01CGxlF6m9q31z8/JM0bFpsP71GXD9wwBqidZUBEm4OZWXs
MsRIs9XT0thah4GHZqeD34zlaO2KQ50mXRoK9dBFFeBd1fKzU69bCqTU5etSaPsX
FSrTJ4fqxX/+k+DvrdJuCwHUpdn36n6MtX62wA+g5WlkJCIbWX9DMaoEnyGoZorv
g832FYUabU6cTeV/DS8YSechyg0CRLCSwExSzFfzBP4jtlQ04cF8GxHq0pXyvPeX
56xXlhGvd97Og5NR5llRgP777PNVSENrYss0F8UH0bZokyCrR5gi3YrPK6FVqdmb
MqHrFojq2JhRLirXeO6R0nkfqpjvBAUmI7fK1kJjvD0glLnO5RGRl+3G2pg/GGTH
aRo2jCqiyKi0B67ITxCKqmiPeUg5Xf9FTLHCH3MFpF9dByIr06oiDe6HBxdT9ruE
aHRFiAA9LoECm5TA0H/G8lsefzPkGbW2JdAaxhFzua+Ntaw4Ao8Qs1KcRT/18gC6
kiacJoWsSVDYWJiDRZJXEQjkBOOuVzfTjQYrB/1l+ZTR1idxjoZ0S9MkN9wqz3g8
OPxGwOqAAnKe6lwyveSKECEZlQ+i40toKWt1S4wer7txQd4i4Q6RGQUYMc6lTi4K
/pPMFrlmBn/HeGdGgEFmbn89+cE4whxZDbJfMS5EPrVWFjrXrQjmakDbGnjYM2e7
qSR3uWM/B+lgS8cXGoNsh5BFsOR1slEwXmdLwh/YyopIww3gGt+0QLskgjrpdbEp
qCsz6kR4s34xFii37pwW9kIf/1L3r4HtAWsHXQvMxcuRsonaGKKFmvBeDclNZtgo
6rMFcREAbp1I9JOPIeXk363d1DiBvnyXUmQ/AvkZfdYPyDFDUXWC6s+9/AwYkxYs
RKFgaHoXHnYYVdQ+DYNRz/5SalUni1eE/MvRVgI1sisRqgMDTRQUSwswMJGL1eC2
7K2skzvRCjxlzn7Y8v0XANvpRJpcAaDHfttZxgafOBQI9sez9Cnty2wmLt6eShcY
lrTjsycpuHrAABOrlzsy0lBHaI/VoLyrGHFkp7aK8O3dgP3pR19N8l+ew/soPETD
/aJtKsbGeVvQSimhObj9pqqKRIHtXWV5cwXZ/yooICODJEwHnzAp6hdG17kTRUmi
Q7/ey5zpUkN5zCMrMzoLaoIeBvnXzoVxYxw2NMBnixK4IprwvtHLkgpbAHtsbNRi
1qoOkOWWunZ0Qsmj6hYELHOp+9ol0SLBoFZYTeN+JiNQAgJtGqg+fpbe5+ZGbNNr
OLMXGlrISG3SrcUJhqoLnMt6UpKAd/7sAVjFNqTsx3EAkIOCHHP3btjzPhQE960H
IczXLjDYE6VHExstakdpsEOoQjcojhXU2vSf1XIiBLaw/sswOD94KymsEQfejWA+
lA0HC0l9TG3UE5ijSxjF9aZDIIn9bN7rbU483WJDh1yMAzM9XyhDoWD7BEoYem6W
9GgXkrcduGuoXZFYuMn1knWPV+p3ZShhciu+bCJHfxRiIfHMTcPMKd+xVknJ7WIz
QIkdoOVsrn4KgalAOYW2KkpIXAZO9QPJpOoSFbXIlX33TfD1Bv6Wf+QViMb9go6f
Lc01frn6CO1xhtn22g4TdctkMu8JlL5rglCFtnpjcZJMtMhqkwahQk+IsErAToRs
q/52jZoqlE3veg0+Goz/chYTwUbUCcKNQDv2DgAof6qLQyLbKPpttHbnZeuZ2dsm
yuEgR5h+infCLabZwJ7csKkJRPScurBBg5xxFHgE+/HWCeHNxm9Tf7e1L4v1ChCh
qoIS4KV4FIIvZtlP/mzTsFCxrtq1CxrOZRRsKFeZ5ZW4ANcNeA6QaoRXsFC5SXCm
74CjpZDtX6OcdxBUmtToLmLbucfyZKx3y//jQiB6kTc6iY/WiWqcneMHd03u55b0
r8s1skHa5ICG6lEyAJac4+PTQbLJX1QTjYyPOdWWXWT0AaeMLbSCGU7kMwpHcPOg
GpAbPDY8DFSJQ+xwMChJEKu6eOYNF81nh+wS2HwGvUsbExrNccgA0o7pk/S1ygIR
RVOijJJjlt8t2AmEdHaAVsr5ZXYekYBErjrPbsXcgMkzAsWHlqmaLnFBjTvn9AIR
F2WfeDwwV0ZjzORuvaR4r+oHW/OSKHMI18SLyDkj0VEuL5FRsv9nhMHGtQEzQl9k
edu52Ud2JUNCscOU0xPch+XU5uoypAgFcNeomNmVu0J694Ak9hWZhTmkxRQPj7Hb
rPJM3JdMUCefjOHbEPy8oD12gb5xC9hdOTkrpA5FaDzzwgkaq08PhP4nT1LT67So
vNFkSyiFTnyQRIlz3kbFcOvCwFvoLrogpcs4FJLSKS/PpR0mOy2c3d9tSW9BdM1n
CG+04yOv7D6EJWrGsTAxOTXK6x4dQGgihj6pgjwKhDa7NDamJ4x8T+rRsBdl7caw
Csd9/XLZpC2Ig94oeJ4JbyjNoLpISZh3/melzweIJcj4nICtPfPRyL574Z7OutQc
wr4aBD+LgwfWJU1EeMx36oJwbwbFxuwNnBXnUiSxgfmK/t6ZBYhHU1F7r/hwM9ti
BVA0Jib7cGmRGQoGqpW1tKLLdqXgG4ba0DKUmIFvoq7PRN8sPIdSEPzPBjtHrl9v
exCZRymZWra1xWjva8Pirfl0xhA3pQb4/yjeYi30VCW2GDD4OdsOag47QfuvFRTE
bIP0Sej705FpJ//Lwz1+ogpZAqMipGIDaSZZslV+Q77/eubmJ3V8RPm6HGpkj2cJ
CSj8Dl0tufuEsjKiKXlyvkivhqP3+C/r/8WgS0QNiGOVXkpfYrGC9VU4SJ7T8OTj
ZakJg4yyg/bc1OcX/z6VEyJXnOKsv2ZKqEiFMdc5ku+D6fw+JdAxsdOZhCDXEvQj
WWD0BNNbFj9euKeqj6Uc628fdv3DIYaDWHnhAZARxQSYUvO7UKFvQtCwPulAz3+4
xhZOHXegwCF08ZvMLR0u64Cd5xFkB7DnprIngR44VJyfx3a5b4HZ64KCQvDq7+Ou
4tKWc7lb9mMbXjfve8NkjqDbKjXB6NOTVRKyJGv1n93IUk1C9aBH5kyNVsWLJTtb
a9uRbKUc9ZSGmjPhifAv+jWWjD+8Zehhubbft2KFmKcHVkcKVp86zOmaSEQwq/7y
i2ZBpdqWwYMEu3r6QIy5B/ftw1PY5I19TK8cXeXWxF5TECyKjuS1Q2Vxcgx510ML
irObNbUy+6IcC6H7er1u3rkau/+vFxkf5u6wMXzNH2gshtDAP3yyRnRAqWkbC5YE
zXFfuNx0UoKMy/6EEBgLHKGuAePovPCS3RQUVQZ6gTL41alXrxxNun7NWv81KDis
2SiRMBx6NGGxK36K5PzZmCRRQ6aAhTjZdlA+DXuYxwELyFjEEwxNP2woBvUXy6n/
vWANU4tfYLZxAoDin+7clhiQPmmx3eRikkhoyS3juM77H/dEfutREOTrXNbzJF1L
3FV/vVWWsPoNmhD1D/nLkgEGRxc6NXeFCDsIdXBX3QDq9KkZdDVdSVOU1qIIGM5f
vWi/GA0A42Cqi032hefRAp8SoVAmRTEQiXHubc4L+mcMKArB051CNN6LrAxtSIra
9Y3u2kyeN1W5KMCQdWM2BLVYTXQMwEP5Ve+BCbi3xOcMQWWogpCMbZN6dbsMiyCg
bdWIYvdvduTzwzjgQBn4um27h8EKdTIrl87vjdB500i1kzuANdIoeeekfd4Fpq+x
wqiq5Mj/K/YxWoYVPbocbN3Ai+YvAVVjYqZt8BH16ZiZAAmtooCLE4FBz741UqjV
71GanR/cJM22g9YHIgLlxO7gxI5QRNPStB9BGWS+evKiOC+11ErnmzIBPoVAxc2d
7NyXRJgYz2OJOs6Mn9dpex2TCpcasacfDRzJu6CoS43gnKPUAZrv83jyRJUSTgzZ
yU98dT+QDcmoWFs29oZSkKvH22ye25n7a8ljBKUaBeB5E0RHbkVDGkVPPYn9OKAT
zhTCN+f1kpvF5EkZR3c9ZG3pEZknJBAfNsltHtd7xswiOBA5vLkbIwws6C60UeZC
NWFe+BcpqlNw1y7RnXwf57E4MN71SmhzFkr81d83Vk7CBGpo2kolXRi75mV/yo0L
VqTUILwKjPi+4k1hxyBtWaYRRbq72rXbDASsIImjeNHjv+dxiQQDGHm6TZjiARwn
B6+M50fGQ4iEUi+YDVucuDceeTfkG/7Q9U5pzWEIfi57eHjRW8FxBsVfTQ8hEIa8
EY3mqjCGphFeNrKo9UmAafo0CuXcH3pLKTX+UWZzuw5R4Gd1xKx/AnF59TPS53D+
YAdIoDDaM76Wnh5AmWudS0uOLRu8EFbelambi4p2DKySJv5JqhhAA/krFAl1Q/Nb
nCmljcezNyHSeT/znbflZXX6ejBucyylWT0k9H6dmTL+VTphs5mKbqBnn56tyf4x
889puij/uzhZf0kFnYjgUCQv+c6AbI5D1hmAdqBtRsFVYNBN9c3WSEEbrsqJGvFw
TozdEop+m0AmXAGG0J8pOkJ4nYpWIFMh+MYREhMiYPqWTouQS2uXnCMMqLImbXPP
6CJgT36bvWj7hpbYTVQIOwbO58PzC6cYhwNH4ZjIDrNVPC1m1WT01AYMrTRPH4rZ
j2HyN3/G8L9pE0DMf/qFglnpu7/Gy9jYdJcm6RJv8YOUttR49rcW78VAFwwPQimC
0aSvtK2WnorarkOvwHHy5jkf1axaokMGlD1HEsVf/oCnSZozodsNBQXrsE+ExTlF
5kYeMBs1VjTYEUWkt48giYen5EDxLTXuRv5TMtvVLwsshoJ1HJrdbN4AuJJkcoq0
/nBg9bjY8oLzyZl32YRgmtci1XFM6UxBzkwRP/U9mMk5EK0/f494lZdXTyhZBexY
rJF5ZXoDfu3P/QIifu6BDYzh0WKVsyCndlJCARCI361tILh3Y0DGFx/plxTCcj8s
SHd8t/NuSg1s4Vmh0314R4e0xS6Kqim+1f/FJYdHsRlknKRgzyBDSahLyrALAG/B
rlaIz4nz+X18aXmaWh5Fg65ihralPqrTdbPldOZUmhhKZdOn1968Dh6KVQ5ybui9
29mINMxWs1Q4HicnvjQCO4P8X5LS/njEwWw0l3Hw1U0/Uhmh/kFfb9tRlrSSYsgq
zB4NRSrvXmG7QvVgarSgB98jitbFO4lpv8ftceO7dP8ZYbvhpE1+OMp5YUfm6x66
cyoIZ7CuyTtBNEcpOHCQdWZJJ23fvb+YBRTSEMy5oJdXpdqvfcJxOpqG9DdiWMNL
hd1Iz3CmYWJc1SJLHs+ft5gcfDr1u6wHcIvJRiHS9/19IJwaIdum/B0YYzhoPKB7
rbXr44tx4flNeC47SuXUmvBsP6FGLZ157/9X0DaDkAKCstjhTzbt+FB3Tl0jkG0v
D2dwWXmUwARwep12bxX7NJqLoixOcV1mX2oXqh9wFkaNUEZX86x98xjVu1RRev1N
qFoF1hjA0GBBGUjGN94GWelzQuyVJqZTOfr4L6Hc/q8GCdHLHsG+7G6zFKCNoyNp
yQabvmUEoeW86RfJzwUZalEFRC9j1INmcZ8+OTEai4Fafd4UryTdmK0u8ftEu9SH
/KOTC2m9b29S4clis3UF9H88XF/dfVa49jFE7KVQ02v4QB+JPaBYz5WK0pzMqwbp
6AX68+aFCd/FzO18///lmNYQRnZpb/IDhDiF9OvHDVE3EDOZWtzLNAPMMEJqDOv0
GnRF39Ryl40YyJli+7pYeRrmrJBPw/wOnL/rY/OulJOnPELs4F9FoVbR+5nLxpbs
KJ//7oOzVHSVbgD7M6JpLqMSjDQqqiI4IikscSJ2WmwU7rIZD7PjfW5wtYemO69s
p7k0q0Bgof0xbLYQI6Tf/jv5mzzZ+copV5Rik/4vShB6e6HQVd0mJ3DJBvH4YNCN
L3g4ZYK3s3z/TeDAjS4hYrkGK2KGI+otrtxQVvpD9puZQroZwnh2f2vRgjAO7G4k
ui2IKHKbv3bzc99p3rVAFFWp4M0AYmjqye+8EteKJSS97ZGXrxOeBcX4CA7U+unX
1jX0ULk6wOxL+m49puJ/OVJhYSgsZaFyhUVMQAe1fy8jBF+TxKr9PPq1hWuvLry+
il/G6LGP30GJAtsQl238bLKxDI2Xq4cAQvY1cGAHsppmw+5IhH8oW/64FA9uuRQD
DOQGPnefOWWEHyBVecD13bi27+P3NcGZ5oDgu0G7oB/dy/UDQY3mzYnvxYiwyg4d
RxM7SHiS3sG3Qxjwj5hXKTT/nT83tdZ7Ec+pBMXbrOKKmxrqKy28ke+J8ZXD1rCb
bJH+qMrfbramJ3TjfHF9toBFr4vXCdhmk+KlKFL40uaPzIZcrB8FPlyFCDchPbGq
QzsDOs98pwsARreBIAzuxG+Jgv2IVdw1xYdFgH6gv3+8RK2MEH5bUL8UJg267+GM
TJi701Hfgw4hO4mikTCvhyE3FORTQjR4Wcf0TqH+KqT1aOuT4BLodqyj0I7QIe6P
d+zc4w3lXPRyYHHsSRxkDVvYYooB08FKapITpEGtthEdp5qF/zqohOXHTcPdgrL7
Qz2IgR5TJ9kwY9E/6nq3PIm6VXk8ERhZZUAsibvFn6+S//Kbu2kfR6V9IDawt2Na
BUHodXX3iYLgh9Jscgz4Ko7WKzZ6eobXni72Pi3IyAZMYXOH1RK3rN83QDfV2+D8
YqcExQKRQCGjUDkMUKN1APio6sPHJyL9e9ER8FC/TOovOBEF5ehCIHjDgnhlh3KU
OcI+3nH9Yy27jBZF0AxQW3nLh1pJ1NLn/EGKg11VmjdepI/shpwRs004sXbAb18u
EvtP4ck7QFEjf7StnYpAsUznDQqURPw+zYIdAmst/B7gN8iGUrCopXAUWaHS2d49
NsKMd4kDXDubgeFg3cDVbbPjDhNTIXhjbuYcNn1xX7icU2VcDoKq13xagagdW+lw
tHbaN1U6SY4DQTegOptpBju+FoQTYIFd8SJVJjjQ6VX6fqG8ezzvC8rupw/BACPn
/icfTE8GxPAiUkvIMuMcs7rk+SkRW5fsIK9AWilNX3jV/z4dw7dAKM3KSfN7AR3y
lujOs8nOC1gTDGf+e9tDtEfvX3CIVH51InQZctGkrMOJreHq3MSBLlVS1YvWjGWV
Y+GqI6bX+eXj3dQYrrGGv9KRJFocZ/o77oSNc+ecoF+4ByRfH4tM/g4NSmPViRZp
OV8Ilk3O4T4SW4NA6hN/lc2CLDXtUnxPYKpvv+Z/OypI35juM0Qu1orh3ar/b8fx
K8oEcdYxWQxnIOtl8cGj15wnanaQogtC/zxdwc6C0E+BJ3lwXxKUOdE7rfHCn1W0
fVSnz3sy07E/xNfZ/DTS0EBz/K+ixt+s9sGuANeEA8jfgglzlvuvSOGwNuCyD980
JfVebK3leG8wFd6rKUehXamKRiaZ7l+HN/o0E5qZa+fGq4GOOeofL4uwsTY3WurY
39KZsfwsIedqiunqrGSIMWhxkUQXJk2dfnMySPgrGKu7vmTIMX46YtVCqt0waA7D
5gxnOs+VMZ3Qa1X1Rka9ja5Fi9RwROQzYPZ/27r0Hqg+bzle7jgVWqfiRMAdmtbs
SQxqpGhSVfcK5eqmDRGwhnZk7Ilag1tptITG483RnxJkaP8ZccTnYO1kVOTO5fTg
tZVE3e5x8XDYpv3oUkGue/nthmsN+Y6tOKly5kX5a5B2qzLZvPFek6lutam8z13L
9zS4NCHELuTLjL9nUZR5F2qnP42LwiN0R8p+05VLsz2k3jXAyEk37VdooEz+88jl
zRye2UBvaIMFPY9b5g/QJGLq/NwwpZp38/kay1FoF+frf+HGY+EN50cH6PYN92hm
CvHjTHq1JjjBtbXSo/ErKCh+wXRiCM26GJKkiGEFoD3btmm1iJx9yCUJqBiLIXe6
GhCRljppHgWaEo16Cj/9WjMy/WGhSrcn/Y+jNOx10eleyuOz+GSZvNAY322Yui0N
np4pxpMmiZRzUA2+Al2OHGtR3u7khVXVvTHJeCPYWN/JayjGYqAkV1GQeOtkONLW
cG5vxavtheTrezKMudhy80/omizLWHrNnJCPvFzF12xXzL21PbX2tLDzGTTDGL0g
Da63r6eDpdPOAIrcyoYAlPK8nXokp2tVIwj0WmE/5xKHEuSC+0sI5YSclteKqJF4
PsB76anmy2PFgCY0AeOTpvwKMsJMUwmjjNDOUAW6ogQ2Kl/Qef5sKwB0RSWIo75T
fRBcwB+o4GDir6gaVJb8qo5ET7UHa/ca/lz9OAqV98bmjw8TbMpSB9xt7RIez81b
/0xRgMv2s/IjCbwan2Sf/y/gQMySHm6C5hsmM2Ti3fcN/IX+zPbbNx63B6iJcspN
fg1FXzMBQRJ5VkqS3u7ZippMtWqBv+9uaSqfSigC3FMdpMvJF9P1z6HcHA0s/Yv+
DuttF8qQ4bZeSVtEXzvRFYV7YWvduSZlUylGlWvcGRZeaSkVAEnGITH2U5liH++d
RAXdSAIJYKVqLiJXWfQDwlVHEQBnmr0XmGfBrLiZckQzbOwmj5oPWtG++OhqtsLO
uhthM4IgynWkgrxpOZvA5sSm+Qt0z2TWVR20oVsujrgd5/Jx8wORUtytxqnhYU7U
Rm2ckXs1py4ysoZSD8VSicAZTnu8KglhLtv+g+gWtGGc8Z2unMRk5jxSbNolv+3G
jMlygk/eafuLO3jdaDo/JWdmCT4kbxiEMs+LNnPmltr8PrnlnFhAFMuwtWRgjXg0
XRx4IG66+6onHYx0zhZLOIYS8Gd5QnlpP9R8HTcqJwhyrO/sRXtoo2Py24gW6zZR
KctTqwQOfBX+WVX0uRUftHYZA65MMggi9YK7WE6zzzfLdmsAQqd7QJPJrkLQTt4M
NsE5IOP5/vqdoYxpXibpH4KoBu230Yiwi0pmDF1+Ce56ZhAPW6V+pkP41bvaO89f
a2hQL/YOjdHMCwqKqPUqwdnW/nZOAgIEqneaKXmLQ2AKTxdZPL7/Bt6DS/gEwlpb
Phi80uyDrKGfU+vM+Kt3Y4Rlal5jkf00c5VBpmqz7TGs9gFIxSTVB2PlWLFPimbN
S9WEnP5TvJsZyqQT+exYPeuZLnlK4O/9i1p+jqr6H+9jUTnyzuVNkPj6XZW2U3Aw
9srX0MnikVVtP5GlIFYy8Gk3fnVb61ooy+paNt5kq7X9hW21pfoj+STkV+VpdCNW
9EWZJRE7UsVBSSDK3OG6vH/n+KuevRaTSPhHMa+KrNu0Tgc8WFEuBXVDxP4c9UMg
Kulory/MOQl9T1WeTqaHnYutmJjNi5WIHGySo2rN3fvpKnLbKcWR7NnId+aNk3BV
oSEbk+gSYA7VfPGAsaiI8QOT0P9yXUV2WIn5XnpikSSue2/eQnCMzRtzNB+31zbq
EZ36Wd7E0LKr5ENAaZGvuHKfN5ua9UQjby2OKSPfPygJ2zG4cxLcK9IdCSGYWbRC
K2yTUtBLKDyesgFTPM3Vi5RjEYkC1PlnrkS3hP/mmpbGJl7PI3FV5MOkljEmhQpx
gTQB918msbbFRaZWxhh7gWbmeYVYTEFHNRKu8nLeGVYK9xkdOo2aDRenDc15bXEq
zkuWoD3cGq9OIr7sWZdJXD33iU6rkxlwgA0udESTFXW8jWgg+33zh32axZV9Us/l
oLqftqb8xwCZZi8ZUpnSUi4JhOvtDoiOUjJo7RxMYQL3qFp9Fk5T7QTIzpiO3MdS
DGgk8YK++2zMEwNmF/0IzkMSMM6ncg9sVaVB/E6+8YzWqoD/dPcCwwzZqq3cn/5Q
r5fQxgHfT94nsSfzbBCwaBGlIbIy7Sfdw3NJGuQrgzSWOdoZi9ixHKwnOx5fhzD4
X0Z5MnLncFTtBfmuWteIz6Y13sk+VVtr1OpLVK5ENrX13PgcdQ82cIGD7UDr7dd6
le5IIAM8/z2/RfMa4tV/TgTl+yOGVTw9LVSAvo3BGybxSj204KS1+fztrZfwPb1t
lyrmPsQ5fa5d8N0jScuyeDmEx1Pd9NvclDi3HymZZ6ctSU7TfRIvo8zTH4MexJp9
bKbKWAR2yxgF6ADr+LNPIw5fWmNF67XGxDN+0TPb9XP1UXQTKM3wsBtYSrZb8Z+d
1zBUHerBiDfImxjZ3e9sBVS64Xuw24rcHjx9+fh5dFw1/2Chj4DjcO3IRFRVUL7X
BTVNMZu71V6FJx53O8XuLynmBDHjQRCx3+BemK1X0BgxJxjlAfWtxGDRZGboVy0N
7I5Vi2B4y3GoicKcLiI4HEYvUxtJN7wnNJJtnhAybM6U/+q+8SvVRUimn7E/qjUs
NCcznmuhsVEQlYl7wTPElQsfc++ZaGQwFCn0GhD0C7L0kBOOc27tJZmisAqIqek9
L2BsWEzFJcT0U1qE6GDktu0veapSSkBpTdlGnW585ew+IHXFofiRJVL98Rc353ml
beLxqFBUPb7m7XXGwrW9qT5mxCgLEb2eScdqGBpXSJSHgtMtnHv0RLWXZr9NMakm
9kolN9KkRgBScjI4jTOIVKsE2Hlx9nqP3AQiQMq3WtnVKzxVU8vc4dqDg/YWBipb
4UrqqjQmYMUFxZrlmREfBQ+NwOn5yMzsGIkysFKhWaauV7QCPdB8alo+btpYaS8K
wkz6TJ/jizewvUHT7hDDsfObaPXF6Anok/SO8Tukj0H5CZZTx3WGy2w6p2dzzNr6
aViP66GKObvLdHhOTJja8V2BV6HUl7FRkQghMX8lCJ5VFHK84tNR9LhtACZyfbjO
z+YuqCy2xNJMIW/4LfoOzJVr45tJTks9s5D7PjRmvGXPePan3mevNaUgjEAei6IV
DLg/JC12Bct7b8u4VoVGzy0JlorCV2filoTUj2rMOf9OpLUdcFZTkY4/lrAVxgdu
YFMS9p5RjHCuKa4+OERt9bkkAFpAf5qf3sMTjIeqUv53xL/mA0NTRNuIA6Xq0jT2
5ETdC9zuxKPaaX91guioqTSR+PvLqzqj+C0Jsq92J9fQV5oufx9Z+hWFCqIAxjEw
GOgIiHXNBsHipbI7Qg3xVqLRpc+NiKvZa8VqXxiP0jQxoYUzPqzHaU8P5/0yEToS
hSd6blq9cYP92rxjALRHnF7jqshH1Q5GZxMcx+Vagxp9JTabQbWJFPmBbpaoxftP
KWuGJgYpMvTLdbh7kWIkLjrZ0kJDYEDuwKog9ikJOrTDCeu1gDzVS/4bbdK+wXut
gcOyPW0Z0v5KMBW8QZYNsuNgwd4Oly8iq7+uoNzRDvVm8h0LWa8QUdjKWvM4JxJ8
gWkf5ahVUD1fGl0TgMKsTfWTL/Lt6PpBUzBma0mIZaSkV1E3ueZnH090XFY0zxiZ
sKmtpP1kkFQQsnz6o9EAiFXHwvKs4cwy2HQphCtciqMy+sJDlfrKYXdm1gA2I4Ws
tS7j7yoNZUGDeJ0F7HYG1MxaXsa8GA2ht9vv+r08LusHNTxW6h0G+OcQeq2FBwc3
wIgazDsEuuOlMtz+c1MX2toQ/5wpNbCzpOGEY7yHa0lZy6ENltkFw//ahG6cL1Jt
pyXWQLeM5fmMp9QVgYQG1t4jjakRLW/iNVp/jU99dUDxxqAa+3FdDW7hfoPHNVfh
3nehJ2pScRNNJhi6nxGQNyzZ81nNnSWOh2+GYLNfpEfFEwSezJFpwt+n+9PzK/F7
lUjQhz0hXzOQH97pIVbfued+vdOmUTNbwaWLlaB16SOsyUe6S4UBrnqlIamznwBx
Cp3E7Xde2R0DYZL06ocfvWz5udZxWPxCPzlN1yGFz4A94Z83Y/VKCX4SL/ZgEwNm
L3nYcQ4PG3LL1emzk0cYwSS997V5rFzUrxdey0QjR/0ERZGUzn/jhf11uBDtlepG
hmmXpq1yLKXf5Pe2U8TFTQizwOGn6Z8giQZ2R0fMSNw2ZQLn46FSdJVzPbyw411Q
ZhsRo9vYMaIPY5p5JPLAT+KbgmvdsuZSekjStYLYbApe81O4p5OkrbpwfA+ufFNk
b5sm6ZA1Ka9JVshYtxj38ijAmwO0GTGW07Pq5BdvH7sqG4drKLBnxvcv2mJHbOBH
lHUBgrkEM9eo5/cUrOlSy0l9uDmfSLhfpxmKkNI+yltFCa6XAdYo+4Mb/8CSa1AT
WcDSJsCg3mT7Hapm5vyhHNb2C1Wvhm9hfJFjd9McAlUMm3bp54E5iLad8KJsTkMC
YypoDsGfqScNQU64xWeOf+PVgVUc+PYzLhT+bC3P3jIvL2wJPKYj0FfJ3GaNvY7t
T8X7FDPqztyHJ+LcQ0y4BIIFKO5JFYFdogH8pvBZcfVEH1qiqIt3bT8Ci5CibMl0
sbuiheBBz0ge4UaiJ7M2DscU7iBzsiqqopDDFiUg0bL71wKcNyoaywHZmMrafXkT
TSFcqLI6nl1WtxcSEfg5YualcWWUoQN1hQ7b61T9333fDDrND66p9ul7QsVORT54
dtlUIwiwL20HTTxENt4H/7vtRlqCk6qzkDJdTIVn+h2qGwaAPhyo8XdUz9hgpVQW
oGroKEP1fPUapIzt18fvkCqeXG8d2a7XOctUaZkw/jAaCQCW6FhPNStarpM6HY+S
XDzE6aAR2wIcAetoby+rueINY8V18WNAZdCVv3HTNWWVsvK1umow1SY1Pjpbv9kh
3ZfjUmCT/hOU1hzWj0cG0Psux1fZFDa0nd8e4GPRG6Ir+edcJg1kCH4zSKL6uPHW
gEjI8M2wtB0HPDAi56TQ3dIoZZL45iKHghhZAqH/lKRccoswMV6R/yCPxqPEYTj9
5Xk/TVq06R//exKQQI4oE5FQNxXaWDWUVPuAwB7q0ADvkG1pPnAwgfnREk5RJ/ft
CBLnObBoTh59TknjZav+HdJP7kcZ6cyugB9ZgUpiDBuZPZA+ciPgbmt3xoox85e0
CItpdmRQelfBpk51Nr9k2dvpyNRV6WXb8l/ZpZ3JOOxyTngou366FQStMXZtlCO7
6hN65LVOE61bqxGit/Zm/mzCPezP7oITac/aD0LswX5ryW0y0UQOXpwTyC+lXT+m
ifpg0OUVQRFr43dSa90x5KgkbymmZ40376A6WpTcoMSuu6OfSaheA2IAyddnoyG0
HghmSu8bAn8nOaDnDKLtgFkTw41RIPK7iJ+n7w+g8Z1rm7C53Wb0O1BSKDYNOYCb
y0JXbAOPYK7a2XQ8YTIga8/JNli+EJ6npoO/Rultu6JsAlIZxM5nx2lKnUkRQ3GM
w3iW8UZdypvqAKcutdVK53ObJ3chjq8PZxx5TJ+4ArKCSRU2fw9DanhR8ETJHfZB
2cnv16ldncAOGR8CIiDUVVPgp/DDQxrFOZFcGU8K8qTMFQcWS+teAp3vwy5+DMvo
9ilRYxUgkQlSk1zB/HQZZ0MB560u+QOOo9dO8arqzkf9wqQ+fT7qBS02OKtSfINJ
jp2dJ2nGFv8FNwU8qe30jpAjCxEGzF5LibJAnVI7V7QQf4Egb98sN2Z/LxQ+g374
6rAA0lYkNlsAO/pmpz0qN5DdwzVfzRV03JRBGYPVKgCcFqQk7ypBzGDtVitCjzDM
+RMH8TCD9qP69YB9a7QFzPSHYTEGITigqmYgncfhj134bgMqlhPCx9Ksm2a0RlMa
0Ni7uTBLPsJRhB1ynRH3nw6WGUDqQ95+EbdQoZdzl1O1+lBrzzH8Q8yQ2pG8A/aN
XmLGox7FlszuaZjtROGdRGoiRBjzS4lHG7iT4FTjLXxpSxGmWv0j4AoUJZPSKtuY
NEv4TgfREvETyyC/z1FBLtIikTWva7v+TXO3FdMWjyGk8GC0vCQqZvIORAnvN+Gu
4P51pxil73EBBH83wQFWFDAUzrzrEo2jqTPJN9cBL4hMjO7jScxJ1DNy36NWF4Wg
uNllDVmXe8aLDewny5dWbL9pxjPk0p27l5xJiiCuIyTKywReK2fulN5KgGoKBuuL
z40f1hshPpyPJ5jtMTk5c9HbaSiHqtBW4X29vAWaqCULJchxgDYULLUPUdJDZbaH
eBNpYcHRo9FgNpoyadzK/Vg0R648COO3hhARstHF8VGzoFexrmOCxvluJx0+66lY
86S1Q+oaLTBD225en8Y4d/pCAv8zgE1YdMXM6mS4Bh/rwSTpfqVOt6JgvqPr74Ea
I+hTjdlsX6SGpPcp+SdcDhuv9+VP34gArB2qC918Pfu4hl6skQL6xUD6j6IHXkP+
ekP1FqjsjDwOGnNqJiWjmxRtrtVSuecc2G4Xzv2WfO8nggvSAW6jQdYfGFRJFHoP
mcK/QNCU2QizQTNqLOL2EJbw72c28UVLUF9gMbVo+cAfqd9Di+37cdv8PDu8Q4mg
Zqb4CmJSVb7aP6b8wBnzY54El0zu/7hNDaBv0Ng09iVEpb7rSrkV3WVGF59iIOVk
51XSXp3fVo+IMe1BNDMvTbrGyymNUuj6V/VQC10ajLaa2LoazqjWIMd6kLmUQL6K
TU2twochvRdR/07KRygbMlfl/24+dr/uhZpCSkMV2e4WZQrvfNaW58dChQqcaKmS
ZxWO9tv7CYDmU3alkGdInpXFCbTn6b/5t5/bw1Sk42KVfvavLP+GPV28HVr2SkvP
m8ojsW9lFlv2y3DJ8I6NbL2zpW4ayBefVLHiru6Yioi1QfDlVR5XjwyVwW3lI2Gm
6IB5pdMWMREuqF2kfWt7YoNLCN7YM0HvgpDkJYtAsLKW/QKC1DwE9pjXNSQdMS5h
3CHnYymphHvXw1ePl/kftCPYsuB8eDkN+d88/jT0N7Akfv6skT8y67lytFs6l6oT
Tz4jR6ghjdyZgtp7D68zsR/NxXy1B1jMbwVtmAh8FF7hSNGmc0B+vt7M8tvgZ91B
wXah1dxk8xt/Rc4tjUhSx3v9/XhFrjZmStQ3WrbDSzdrE7pwA18IYFH+hcsOaFFi
1H5Phmu9Kys07VefAJmK9dF9ISYlbAm6SXU9bAtfl4XF/2v+Yy0kAmKtOETDPvT9
nMaUX3g4i1z35SFjzhtdeM5KM1wX/qJjO2PrUFxMmoowNGYjLf3dPJDSoltaNgXI
bylFdEP4Xjh/BCP2Ube/LyKf1ZmmE/exaBtPZhvVVs/ZT5A66mSb3Sjdqpe16024
uqgjKAKL7g+j8iKKRVR7cu/iLAq0Gn2MuhkpA6kiCHHJ9BQ03grawsMXlY5rVI5d
AygFnAqHRfrJ4YVGIoIEV+MhYt+54RHO2ZGdmMnD/eJjcIWwwZSTBfr8sLV3mJGR
bnUDqzHINZmK2CqwoH8t9NtNcdXA1ob/z57di56V3dRSKUlT09gOQERZm58hmdVH
tSUKHCJB18XCMmfTDH7uh3JTBO1e/H/Ya7rQc9g9RhfMus/AkLDIK4ZDduGd4P9L
Q2h1MwKdv8vACUrViiXjdslq4EJ9rZTHdd5tKvVvpDuTok5H47tDmE/D8T2uxg4R
2vfTNcFnSjuc8iz58kCVYObGyxNl01cxBZRulMlSAewbL5iBcS5ppXjmS+B0fjQy
yz3p82OUdYq8hCw3oaD0RFAG0DtCp9Y3JQRbZoLHU1v5+kj+EEdccyKccnSl7EQA
bLm4dci+r5KfZqOs9rxENBNNquzXPyU5hkOg/m29L3FBmZN0gZYUy5/AnFStDNJT
exsWvyK2P5tmXtaEsa5rJFxW7j8vmTOShvbuG+IkN5tLR283JY/k4VIabN2Rww6G
H1Z4wQijqqp1fBU0jcsxDCUGjjgSya79bNutE20rMgytpYdx8AWh5TpMQpHbgZAQ
FftrvqGBRJiOd/JkUSkibysCFZ4dtT2gLVf020AMnv3bpIpeaiDi0uBumool5tnx
SFV7u47F8+hQxj5Dv1cFiB8lZY3UA2FVn6FOB5kz1JpAwXWShE7hR0AGpgCxWeEQ
VfR0gVgdTjWFt+jv300c754KJJat8CjXSCrWN0qeUvt081grd08Mqpj86WabfgsW
b6BvAxPnU5rrl4Mk74X5KHjytM310dLuOfIIHpkPkMLc01CTkzyU92RJIjUn+aNJ
ZkbXmHURiP6DtaT94KN1rChdHmHook3LWmGS1jd/ibhPb8p99gaMebhdwSVsDvxH
jW7axohPFaN4eRsf+bvLb0t6enySrX+MpbtTvvv8/eqd2n89uBiXclZPFW1dqUZq
nXfizk4kTrPkznw6Zrcfg3G3DKjodPxkouM/41i8WsH4hHbjGx4tj/NBchHITcJy
SNnl9SDozsbC3+ANi7YndIWNvpk6nygyrbLQpAdkDCcE9lbB/7/sI+Xwb6gf3BkY
yUQAKqVBFwwvH3BicUSlXm7TlBvCTq4zpCilzaO2C/hJ59guGfUUJpGTqfG+9Mgm
HAkc6LbdCQGAfVtoLJW9fD4R35eSlNuvNnrX7V5eYKAURnZx1hXD/Yza0VP26tLW
CsxC9TFGYrZXWn/j4iBxrvgVerPAW2tr7rviUHYgj9zHLaqWoC1/UUYYK0bJOTKs
d7ixuPBWF7Z5pPxcuzJiglRV/Ylq4cvwBHfAjy5kyEBtVslOViY4z4qz1MMw09yM
ffSVdlnUbGwBPKFZMqmxnN4R8xMJ0rBALBTOhkf0f1lxn/GEgBiSNws7sWooTRdU
XHv8LziUdN+ev+y1YRydtjIw/+ZQfhWSK3ZbScoyluIJTUzOiCkQFnMeebPtRF8p
e76yl43LDbYFXWMU+ZzqWoOfXkAHgJ75ETFnkGLgEnEcz+8jsPPToIz0FDYYjL5F
aNl5rCuwzThpOmtalsoSpvFWwtCsX3uGk67wJ1zSXFed1+lKuidNLbns90+exi4I
6bJf7BrNo1dTDKH18daIHe+YZpRxFcT/UhawrIqf44JS5SMuXGHS6+oTTnU/Wnuv
7hnRdKeutuaSLJRzq9K+ZU6lkLk7valB86t23aCt3opYiwoaDOKmVUTx/qKX4v8n
AarKH2BD7BEecy1qw5mgNiLo6vzI1VZTa0fbFgNP2jPXhQbQ4xV7G7a43St/cuKD
xKA/76wwr06sJ2J5XfpPKiokqR+dPB5NRSnEnFClUnh5+rMYzao22zF28olnvOBO
epttbsvLz5ECyCQpIEDtpzaG5s74PGxFG2Qszwh9Oe/Mf+7fVsCEYyfrHkJPvvSv
MNUH05QR27F0wGrhnLdaBPA07+3E5MLXrKDo/nknhbIELrh7jRfC4wlPAh9tczqm
7TtrcDIt4b/cadcpyCNF3ce0gsVUuUpkHALfZX2aNX7t8BHV2CRtXunyPtKDhRFl
WmN0Yr7++0RA0i2NRHvuQYwVDV3ZRz+P5FKx6sxFvjNKX9CEW2DswmmqNyUrloOE
x+ATEZcs80XZJD8MXWOfRv246cSNDJ2pBWWfr8et3WCglpKODZy/hf6S2CWKKyBz
Xyf/ZU76/sHTa8PlYhrhRXZcMBHy4Qzi7OvQlsh2wfXcwpwGVS/bFBxPz0L7HrOv
wiFFY6OEPZ3jDBG2DJVq7XypkQZa300aJQNe8hQmAQBdHdouuRHUYzd1xtm8PFOS
nzW3m/yaxlxYqv5jQR2I+rT7mfRe13qimQrUUahBTJk6LGrQ6WqtVogj5JuKOlrl
I1MUsKT6KSAIEeMcXl+PmW2xheUMeImzlF6ouS2Oq5oECqIwc/FQBuEB1nFr7lIT
foyvAA1Q61rjUFphUeQ8Nr4rAWwOjdZfOouJAp5BN8K246SKgG/FarMk5Whbhfbd
HOYr9+dJdy6RyNR7haY3we3OXt5u499/5xg1yx0EUtYHDrRfP/mbo01m1S4iieTN
rRWaO/+p+xv2JTm2xxg5oofBhxA2QkIBn4A+0/ZCkXAV9mfBfpB3BdZzd5qZuSyC
2pfkScsL2AHpfX7ZO3jMBKCpCs/DraI2tPj33ZCFvQpZPehkSgxBk8G9cGs5k2Jv
yz9WPeSNYuxsF/p+1JYDEZ+gIgcgFNQj94FOhSS8tOBMt7QOEM0CIbpP4oVdQ+ec
KegdrXjE3q/WikK4x+VteAJTi+PjoB4iYNuVHMlofWCK3EYPEOGQFOUKe6hkGf3W
srutlHC3Rm1JfyqIU6jaGo3XEifNUVNl+7+Ui2NHQFAV5Nhv8AEb0V7hd4VLFAYX
f8bC9lHsjGz3vPhp+PKFilPZtOwtmSR1SGKlu5m+vXHv9pWynHs1kCtHa2Gn5miZ
dM/ddso/HlP4rQvr0B8B7rqG/3pBYjn79ah8XuOTmZVj3HXO4KhPtw6MKzyaIeQs
ctA+B5LeRBYd8bxJhlCkltDqg0U33mQPpkcfvPfSfxtwcEs9NSoaoVbRQ0FYlndD
YsrpuUavGAiQSbakxE5DJgwNo00HPDafeRlgzS3YjKukeXKjVwcDxZx0IHqpDO3X
n80V/gkrcj7hGajNX0uK3/IAKJF9yagf/cUt+fYeLF7aYU5Eo9NX9salIS5HYbwH
VkPblviKcLPpaHATPY+krhS8hAqzPQqZTKrihXPwDAk4P49QkSZUG5gh0bT8Xyzk
6kL40hQXlmWEdxvN5YgR3VA3ztqmARoAHjvN0ap5M2IZommBgdEn6MJopVkPOLfy
AH3su/ROXvx/2pTvEf52CDFnquEiN4aUHtJJ7cv1aEOCmmFSSOEIKV48pnJ1SLMb
8U8Ke5OkBFljLxcYHcfXO5BnqOJ3JkFN2UCVq1F0JS/jxDt2mvKDmqj7ssVPffn1
mdjJqftDS/nvmmnqhCDok21mQiLUJXMpyHHJDImPt2gOLe2JIu2wr6hcE7EKAH8G
P0n1P6PL0exdvIxRYTbEYLgz4My13qy/Zy/eKbJeUcCjgKQsUt791BvWvhRBihhw
cRw+JUXbW5/zsWajy7yORHDndzUtBmUBJIXJ1ozMH/MeR7FAP3lQUxbQ1JHKOuNM
HdY6bG4F5b4CD/7WhVWKiAXdWh/N96qi6xT0uOqPVC/Qwfc76uZOKktNKIL+jYDF
gPnDGV19znUTHVtl3MeYEb+nrkcr/y+9wHUkGxPAdRLVZ/gleHmL/ggrEFia5KQX
8J5t3LHGFBWKoADEEjI3ApBU4IaVFjliof5nGIQdrSkzvd21MY86qrUIqaLGLBxg
lm7euDCxEs9XoWIJ9y7oKZHWKpozP8k9w+HQz4WGmI7Wf2TDYCVPTq32/r6OH+dl
VvgeZm2Jfi1W8tWxJfB3FFCPn0CWWVjuKk63etMb9KGvwKxKWcbwstC2wke6TAPl
hPIXH0Hz20AjGrwP8ILpSgLduxmxIFI9mZjpbh7QPAmEJHy2pl8GYMUfI9UdZIik
jzUDvr2HxjtXNooh12klEGxefbDDTmdOVsS8SC/0KK6Fob7x5W30zIHLTIGHtNQZ
ACUNAOswlpKg66ibIOiXkCtzfsxPAvpcIJLiT85v/y84POtbTe86p+SrV52QUq5E
Auq6JSvILTybFt5AGu6dB1YQTuzNC423SfgId2vtCgBP97//ixObfTviF1C70lCU
qh6fxYqJIOxBYUm70pM1mfRDlse3o9Yr0+I6XnA4KW7BRE59XixmeU/DR3BD4YZP
IdsnujfsrIssHeJ5bbcUIQ0K6sXd6ZLgYg4wna3P4xJwSxRFuXpB06sBQq8wsmrG
fDm9p7an0cKjs6KgRslkVXeb1fkjVyNzBcc+ffZcp59U+hgr2BLxnf2OqtGreXBM
WIw7LM+KG9NE06oFlG6j4bErmzJgTrODezQU7lKOILi/kRhZe8nwAO1mOzGCyrAt
9CLXLyHcOeDwDbSNAD7LpHEVSvcnQoZ8rag/BlSxznSN0Ns4augldYHaRbYUD7c5
pMdW4z1jp2uxNeNJJvifY0kvO5J+njksjGN3/5Tiou2o1zwcER9xfmmHv7hH9Ksd
bnryGHH73ZVjMvlsYFsooLSysjS2e54c9zo2IcA6l39gET20xoD/iohfj5R3wTId
IwT5Co8w4tz7TganIzzNuNX5y5TXEmdWz74eH0PMZ6Y4Gfq2RvYmsisLX841Wn+q
PKxYNzWMzxfNjphbA0U3rTCCZtkglgX0ehFeCY90xQvjHMekiLAeEv+Y/B+OI/xk
vrKBxD/5vcpnTFWIfrmk4iDkkmrerHQFX1v6eNATqLPmsuqIlRafSMoLMnSShqwJ
zczyXxdGS9FCQOFOXEkmjVAWYbtinOrH9oZ4vtvE1xPLBzkpabzd7PS/UW/DzEuz
fAlwMt16WHZnPUGcMvDaAA0BEnocH3/8YlSyKNWYU1vyJSoB947BDmt6seeyeQVH
NM+dBkyb2WmbK66fcQ5SMByTdo/uWQBxCmRB4aygqOx92U+R6TxnRziX1LvFQw4p
sCdtVXffKz0m4QSBV99k7lNR1QXqAp49+S2Ud6REA8Gejfxf0mSiXbnrRKSHl/pc
cMdfe2HAtj3HHJl9GoM+HtH6ZjGFq57RJNSINHwNacgrA0RnsJj7xf5xDnpPxRnR
2ONO4YygXr1bouEN+8TjDJ32GNzfb8zT2VKiCHOtR6WDUrwx4AMLDHeFlM28Khw1
DVDVkJ5OxtmzrtnRdQ3AtJz7CfI0Onwms0EqFIdEsJGPHpyLrruLIYJWBNcejWNt
c7KCuXkRAp5xqivcjLPLI8nwbqbsqbhTMo1YjphwfQVbRPWapzWnr7oQn2ctRi2K
Xb+QfEukNQF1ESWD5ActnfD0lId4u47obdRbmjqD6vOT8/ZL/OQKSHrjJI8SbsVb
2R99aOF8nBOfja6o8EpNHjaWsdAqnr+j7udMOxcZa+dpLt8CieRHTz+2RT8qSwZh
vy20DAkO+lk8jPjG27DnmH5QDl1rUrz3YmtiSvbXL3B+F0qBulmXuOApYapL87l9
UogSIU6gWXjdTOtQuxY0bjekL4Vjbz/zX3DNuLOPLZt6250AifKUAbs/tYtomMhI
tdl/YdD27egLFNR6rd8uBcVPnXHg+XulygseF9Pe53l6HVNTrZHVYb80LIEONGyu
OXXBT1CtjosU/tL+LBSW9b3j1kCENcmDpgyc5iEAuM/VPesDPs5HsWj5cZkgavES
sDjde1zfHm9xbyyOdSiXpxhwDg4IvStLyKrFUJz+AQAakU6caM8HGYHyQlXGDi9Q
gUvcpDJ51Th0rYcBQTJdRpXQcnfjoHxoZLfWwhCwnkTj3Y4gkgC1bnxspp6fZ/Ru
2IoaLnjDbl4xqsKDsIz7lq2I5QZLHHzJSLLUgKtzgv2+7NMPO7slYIbffE9dByKY
6PUu0wEX90p+DrRc9hRmahU6S0r5j3XFnF566bT1ersUbMrs0Rri7l9vEE8cZ6oq
HXFpiR66IcBWpsDfQ8lEok7lqHYDbNVxaAzLy+gbWYO0fk8SYcIxyMQCoOZ2nrNx
ZPkKky3AWL5TAYHs4TRwOq0vNeC3hlnTuXLOqdwBMUBDYlqlTcwZB5BbFneOn+sz
HcLFBmusDGDiZnohnS7wZCWvr+Xoy3ETP1r7zMviMDmN9nu4hYpkTIrabtWqJmVC
wQU9yY+jLn31TgZYodiXaqO90yF25DsxgupdDQCEhVR2O9NUp5P7yvFDc3m/bPjm
OE2feTWEyxT5UVLMXoLAjSmBcCjUyvrvmRIGYs1KhP1Aa3FE5jAnY66ODJ7rHvKn
eejNoPmzvjJQC0Ng3mjt7hZHbwmTxEBp8PGmcHN2MJO3q/+EKstP5AwJNAc1uQsL
tNIgcLFK+Wrbu1cPpLLvdS2g0MM30uDhgHv5Qgy2loFsLgdQDNvlAnaw3xyutoaO
D5wvEgAfTy0JiofnvgUyDAXv0/ex4WhWs3rwDFeb2dPlNNs2v+/1XkTFuSMnTYAg
lWGL0odFujdipAnbBvnb78WViQLRNRdgEl7VB+FNfRAUTkWmw0D+dC+/u1Wdpj5g
snjvBbNvvUS1ZnnCAt9M3nhpHB+n0Z793CyzzewAKkTibqQYWOGfwd1IsfqhAMvs
fQ7dIBaVJOsFC9nv8dm2iNpEeJ6W8eXaur4Zi13BOBgspiolxHtaSGNoHkj4Q+iZ
yVwUKHI6WFiAM3CILMkD5evOIYLKW212dBI9DfjnVHZqDKLfQSw/KiJ24c+Lqzbb
U6V4ynqdW66NvLVCExUgpmPerkI/pwVa1sLRwEjF0NIlr23VSrNnY0KmhO5Xwfzc
mmFvzbZ6xyduvCY95V0y7ThIkx1grQTELSgESYC8chL8Hdsbyg7K9G72d3sa01un
S3/lBrjpEAgprjJfGSJH3M16SG8t1SFpkoIOg7guDIOXoXkTVIbXM9gvWGz6DTxe
75SZOGvi5JSpX0SDxXXW+I1rxj5qqUxQ1leL3SRAy4mHrYgSLa8b8T6o+AAkAhjs
7Dqi5w4THUWTkG2fcjyxbX0mP6pTnUBiXb1mEa+LdIGiloECgNSz18MQw10gq7uF
ujGLgd1z7A1Ts2B3GD3czkHaUj9EyMUpTUeLY/fJEbGipYWIfBS7t8lS0HLcnSsF
Z85lqvWQDk1ZdYHn6QHT5DFOSKNoi98KUqxwWZnQky/H0J2nasWLkAIKLysKy0lW
FATgx7ASoklx5GTcc7Jz6sVAb3zwoF4tPf31DsDfLR8VJ9LFv5xGeQ9bnxhm37/s
OOP+XE8uy4SCH2n87Sfo3jg1OmZeHODSRGsS+cC9zzVhYbV80tL0DdYNYx5+cBjI
EHCf6R/d9QbgLkjxMxXXOymsl0+tpLKtxtkrbJNGowUKGXGX+286swE6AuRHoOPu
/g5Zpgr6iN1Ma0tV4k3Nef79HPPmbpu8qZIGpWqssjTAnKAO5+rOfROLRwuKw937
lez9GYfnO9+0vD0tCD+WSN6qKStBDAeU5ffoWSuxswO1l+39k6cnh/i1t0wVv77i
HgS8nrjnrhEnCcmzu2ATG/2s/bGA/lN5Pwyr6zDE0wYKWXlLGWdGTxIbmG3wUZFK
n4+fGzSII0GVszJpO6q8YmW9u4Q4NmstA60jk7J1UV7nnZS3/ys7OopQQRwuNgHj
NEvVHRUN4jb+YUCw5KVAe+6iyfKcfMr9zgyr1q4/5vFo811LWqGxwt/cjicWmkz4
cZEUH/j2zZ88NyqA6QygKHbW4HnkYNwB2BIsYPrOuebwodom1aZyntld7lf3aj2V
PGpRCGMj4cqX/PEj/Kf3YCkjVcpOsl7rjvzbscRXnPyrDuadYvehCA+UoLor2+y1
0qrhwIaIrnng0F7UcJAOeWMMbDJE+xVJMpS2Rb0OYO2ebhelaUJCSCaqXkj2Pyp2
DFsn/O/sYxbA0YF32o4rMzSOcOPXwCT/aoZpl/7YUEawrGG53bql0LaOs/xFhiXj
uuTxW4NA2TgX6UDA9jYGzoQOwbNDfMkpJ8qQmWDFZtGV2LCfv9jf5cwM82rZAc+t
CiR7Iy8cDZBmi0dUFcTFnIyFAni32TCX8G6r95YLCLkQIbKtlFtwEJjiWo3aAeMs
3NfxC+pnhrHUz64mCgDYjph0aEsUIYWrJSe0qaAKUS4ZASOPk/mTc0tGw1WxIG3e
huLPb0pFrB4mwjxmDkghBt5Yn6jA2o8pgewPKI/GUSAYVvNiA0sjxL/A8rjDjtAR
BLuElfWfTfXyFNSudZY3EvEah7z2PQWy8E0oJ+EyWzawyyhaUTjOqiON9jrFHiCO
Vuw1XQN8PXTGbvta/PCtsrkjYXavJ8S9Aodq58GKZSr4K8GHl+1NaEhTjNCP0KS2
k/K8eKG50n2Y2dnhZOfeR4sJo2UfdGQgsxzvZnI599mhu8osX3/BYj4yZbxBo/7M
ACOQ874AjAYzq2azNfMTFoaFvWdv+A2IuAlcHVOK4+5YhbCCwEDZeV2C51Fqax9f
Uh0gIa8W1k10J8t58Ekkwjq5jT5FfSCigRhDFQvtBI1OjA+mfO1uQgsl+5XKhPT+
nDJD9o+BTEoht25Cd+W/ehHHDDdYikXn+C42KloelSch8viZgpJ9AGv0slTgYu0u
GhV9Zau2pCh/8/UDZDH+Qx9wXN/RvnOv1qWncydP0PEBJl0Q1HSt7qeS/DZsAUV0
sGqvJy6kq6/XJRXID9t2fUHjvk3gY3Iu4qHuAhK8Zf89lqAkVoxlo3bGLOyIgP7H
/YvjEysXBpZgYbF97G6Eq2BgnfKHhwETXlntKq3oKDCUw545Pjb3YrC8iqPyKrbX
hV61XjNWRaMOx8co++fLmEeZtbIxMcOYMn6cbjFJMjYtQWfJydWKWT4kh+qSJAKl
Q1bAtqTtplgOdIJ5bsQruZVKTQGSyLemDKkFxVdQLjdHqvqR7K9I/K9ZOJoqhk/f
/Hu4AnSLlYlqE8HBsq4QpgtRLHgax2dIT7mbJeB/fcjdESILu1PERg+EPbHSHkLF
7Wog+ARxYYvThe0kbTKom9mKcLcA1n1rZOksMhOrnRokC8QcmjLziztVmAOVikXm
DHJiLB/Jr5LyYT456x9dI9HFQuThbtOH/7/cwYU3k1Z/wY9Bb7IJXCyQFsg/AHlA
lS6js1x/J4oGyJwCbmGThSK5zV1pSKe77OMT0Q8E0/rHY+dsVGP+0zKYubtDdWXf
3EHezW8jUmvrXnbsAM4O7Qqiyc8nA8ru0aq1kVFd/evEryT54MEGD78DXmyQWzgc
cAFIPFY1qIknW3Iivck064shcWb/HOpxcZACYPwZMiZD+lxTm54ilaIG2PnUtmpx
xOlIyj3XWJt3ecTizs0ZWULKxVWMQcNvIGePulU54Cwoe93GkK0kIdxcPclQGz25
008LF+93NUsMaba6nI+XVCz2BwtcwjTvHZdms2vHi3A4fVxsON8M8+e1N2JaxQcg
H3K4iUECyVFxgNQWD7kK9M7Y5embRl2877N0s7BRe8sbOelHli58B/hMIm66cKtO
wVSuZYsWcJA3ycoMaIPyp076skyE643ZlPFCYfJin+fJKqPC4T8zqXKIqOcYMYkE
5iZQxuVrVj4E1UQ/E/NuqufDdYZeeX8dsCk8DhezW7vPhVemQYX+0ArX0XQlqtEC
B0Ex8krJ91OITIuCNfIlq3oCABccHFNtzXg9sizOeLRHPvN9pbzogzNI0qDOygoS
vumuHluRe84OQ+RUxexrjePhcDn4rYcusDKPAsUWAAmKuKYvyiVSRapSdrdkKiFJ
0uzT98sCB1Bp7ShnL4g+NcNmkUtN5MB0vcvQYeqUf9gX54hscfE81mmPNNi/QTgy
empfLeOwBfyQo9+Uz9d0371EJVSyHFES6RRQzIoWt0AnLK3Zn0T+vWgKBEoeVF63
nYNxWal+RE1Q8nIN3GI2/GoGKm4T+JFfj/8z7T9YFlCysWzOCQDu+ymLF0wax5KB
mo5prMEaXskQ0ObK5fSzwPRRa26eNoUt2/YIYv6kI0IDep3lnLl9Q+N/bN8FKsGD
gJ62WCY8J7P1ombwNu/Lp2qUS29soZvi1fASquxlB9iMsdIWpHYXny8oSNhBe68Y
TyaSd1ym5WGeNHs0YW7cWcJ+epXPbWDz6FYKnAfU7EPfLNM1N5PRn2+8nYdF4fA0
99zGVuPEnkHenRF2Ve3PoXZe9RQfZIgDa3VwySGloYYRPWUFuRwMg+vsKlID9qHY
1uiLnnMDR3P3963lo62j1Z1r6TbX9S0kZF8HJ0nb2PddUCKKYGcoB1rLmahfqP5O
PtSbA8DcSGjGp949iwTaZPi8rYM5QL0M8QBhHvQooVbJd6P+g6wtKNznxU3DLJ/N
9gaK5Q8CqEmIsWa67AFrwEfgrS8/QGvsV7Da5CYIwr+jf9YJa1S6140XGbOveiFe
lwL98xzrwt36sQQdyx1+AN0P+vVIhflDWx72lxkGkvYPKV47ZfbmQUsxXZyjfMz+
QD6OfvXf3OXCsFQH7ZSpgAQjmnMFaCmxX/Ja3R2Y7Pm20DQmiaOhaRNHlnBoJYBU
eagEIeY0fu9pB4454JYjmVaoPUnc3k0b+Bfnnktxt6uXMIvDObdrf+0XdNy2Jk+h
2wQm8JoocoqAabhO6mbIvZYYGCRooavUEggtRq7pjl93zc+kRCGGMufa6xtFt2/Z
JXn4/n738kADhgWUEygFce3ebe9Exv59Im07GOZ1MjgPocq1TJuMpjNZA6zN5P5P
tl8Zt6ekgUcrKGAD9TE3rNAQlPOWsV/GEugZZuAb/PeiBrnYTvpudSgFNl3/o0o4
+aibNkQemBnBreGb8aYaTfaqrOdRvF4/CNefz3G7GOIY6vDPNaarfRdsN1eApnd8
1THyREBMEzYziCcPBv7rcS2GlAGU79LaxWlUL7wLzIw97s8kq2HTAc0No5GMJmQj
cs2vMhfwqOjP+406EhrChrKZ9h63LsW6cPd61oP85vI5q8zOYL+906N3Tyb1TSt7
Pppa/L2T2R+xRrkD3s5+gBKRtVLmyg7XmqcVDpHughC0E75FyFDqgj118ND5tqcL
GOnZhD6atKyGIlzRGvPb7axc0fgZHv/vqRGUApykd64tECSQQSQqOwcqu94Gt0Y0
XXhEFy+pJ2xxYglGpnG6sLr8B5GarnGPFGDO34GSsRLO0elJPPVVI07HTfkmvdC0
YG/Gd7TyKh0qqcPB1tr8CbHuPBV4dIZEx7JDWRKz9ubugCpbYsKw2xIysFSv/O4N
QlVbinx1OjwYW0wGujfIOLSpDxBg8HTT9rKoxeh3VNDAkgKYihJtpX58YtTfP12B
6MbiKZk1bUzFLlP270eOrxA1r5hBJGhXb+JIzLTSVEdXk1k3S1XvK4cyuPhjXAzr
+Q+gsCl8Fe4HOjx60Pby5yZnO4BrnhIrR7vhthK8/+SFwVniabCAUp9mcYuCc5NP
xlmM3wiO4boJbIW2EhV8nS4e3Dzvs04P/ny/CRELlxVSIQswLnWtDbwfWWawjHIF
43jo4sdIdWkz260W5tyN7cgWmCjpBy5j9dAqPcWcpGrK21nbc1X9pfGLganIgecH
K7Hr7IBJ24rtG7ODBWsnhqA1zF4vJl/qWulKpF1wWT+4jSIKIcfO897AeZqQM3Q+
Q9/QSllCat/y+MaTu+gr4vVLSm6Z1v/32BqdorczJzwbQBrXo2d73PnhWbIdNx5d
aFHjxoQ0Y/ZBskbvirc8AgCwSOqIaoGWdFTIaB6936Kj1mu36VJI+QmK6cl1mFBy
s2kAFPCXlRBruTBWKGyxO8SBIFG3pDGp6HA/V8P42LD13aS7C4Z6reas0ersyjYD
Ys92mHyQ3y6PS2jXLGPvTJsgkVfRj+X4+YoJ5/gc8XvzDsFJlGc3TguYxS/ECbnF
NHpel87xxKDFpsIzuOiCvkoyO3MN6o+kw1ZUe29sorFECBt2ZFlop5V1TudmRCT1
OFIN+k7hg1OI7f4zCN8kG1cEAcocAGj3eYGTdtkcXc2jMK/6EX1FnVnA4NGZYKG2
q4V6kFyEjIn1N0jvGTvGamBJmvQS5XY9i7tIDlVDhIZ0P/jqzZTtkCp41TBxB3Qk
zFd4OOxsE1w2fgRIkjAh0LqTNsh9JVPGka/ykFv7StpodkpeVRXY7NZ2LX7fJHcw
tTaq/Dz7gWmdFM+0WCZyQY1o3KAYNubnKWl3fj3oXBJwEhJ1zaG2XUyYvbTs6tvk
0C+V1EkPs80pSCkAbwAeKDPqPkW3qs0saLAbrjdR7sU5rhWsE9j40XOcm82Dcapi
rGPdpk2vNH+6oC1Z8onlEUOltyDSwgXcDCZ41UWYObobOV+gvHiuu4dDkfs06du3
7VNZ7YQQd0bbqVvxnf7SvrjIYbMXXzOQ8Ks4ugYcbhWeU6AiMD43OfIyhjCAgxVL
yGUiskkkF+qshQq9d4OLuS18150atNSeXZ4FbWM6HIL9iMcGgx1XFXEFDfoewS2c
ayq/DxQZAM8TCBqMJ6hrNHaehZbSz6TIjY2y8P0wwWB0PeBpZPaNmxY2Ra47lgwa
pEBo/eYmjjCALELBGEUrI7/BDhC0ukwdN/ujT1Ud+Vhj7Rjbwz7xLSOzGt9W6G4k
GUwjKDychusnJvWaCgEtAdIlSBQ1RL7xiQsroryDMylZXO5gIKx26mkUlSiAH38F
y0YHnJP08uX05XZhPuXVsrcwWB62IbkfF+UjVqEMBg7VEs9M21uKtFRt5K6hjbTw
W5Rp0Aq7vF5bHPyMnyRpUI4/8lWidBA5ByIUkfzMnDEOkDmae9cdr1MeeoDrGmee
M8Zqv578iXamGwmGuO2vlSRzzVLb+kuvzpKpW3ljnBZ3V1V/JbDX/0in7OU+jLGN
SBaoj3vecNU82p/F22bBgNXhRGOpzpQoW0Cvwd1dQC16SLUs2s4dbFUVkdGuE+un
YJCb0fBTnG91AONApDXVYXM5iNgs62lUL4UGtAgcm+Q48ZHuOht/v5IsB1geHS6U
mQ4BR6MROjjKO2IM+qSKP9Pk4bvW3GzPLk2HfHlnogBXsK7xkbQ76QsmyOxxCVav
4WM2NMQmSPmtsuqYpivyWgidOqsCsgDUVXue/+c7woZDahyD5QERO0FLxnLv0f/H
nQFTELYIgS3PCmnoL2ifX989RwtGA5avCsLoZP+ZWiyZXylhd5+V8Lg9XooRwqUZ
leBVz5JmCsNXTDKcal19qL/xxnmxTokIOEYyBeTLbFvsgCUUeG2n1mPNSMt93cX9
iBBW3WsdEG1HSSiWvvkChrNP0ufFRCJRmfxOXKw+YPWWnOvkY7uagMpaZx0X9yO9
NICyHVKEoJWULc2U2yJMLa0phnledSl9Mtwc7PCMPBT4/Pud86odpan6v105CRdl
IyUu+Uglpz1FaPBTZRwDNR4mnTw1TdaJd3qr5DM3UTE2UifLtGaixlb68yHVpGaz
7vTySqQRtr+f3O2jka6YbJr4nkXcT0GWulNVEdyyJJUXCWl2Ov0b80rIqEseBeBZ
SxayBAYSWLL29AJ8ey/j/DpaLpr/WQJ7ogkQJwFHzTSn/+Zc9+RnHd94jyRQyxLW
6NFnLz4nQKW8mGyJx36/Ad/5YOFkKJE4Bi0mqqFktHzXuPYS6B4wfXwsJ5MRTnzI
ptW+9J7ytfs9iP7xWe1wwnhwZaLAI0J3TriBUkYDULibSYQ4iT/q2TeyQzd5QqIB
MHurbAR7KRs0kIXcoi++AcpRKtP047mqsxnakznLyYQrGcLr/HHeDw1prcGC9Yx9
4GQyN4TGhFFX20e452v/2bD4QYyjiya3eyU8kQ217iewRziPMAFoOutKoa1EeLsX
5molAhBq090d79aGzV++dpnEEwLsowgx1xchnNmTCpmxde4oDyWS3UtiKSyCH8h0
LtaihqO6vw+JhgTWC+oZW7G6ltifx029bzzV3WdBsOq76VDMwoKPmUBSZ9YPxYgG
WhPUG6kgo7OQ3eLdkhONTi6G1Z//wcguFpoWTnEs0gSr1K1n65iyTv7vpdm9v3pk
o6hre+r+7ZtIkcm8ESKkaMY9org1p1PjzHJBik2PLf4ZSAmZcc/7/Efd9dUja0q0
SMce4Jd+PGcZspxUWnCzr1bVbHCdSWLTbXuJGYgrnINiYnlDqTrDsvLvbEK8jDce
PNmCrwI4HsbzEufF52qgV3sgCzzSB2wMzBbz+d9H0zFEnVfkfuA8ta6qvrT6Onpw
uTBxRW7glET4zQLi/Ovgy8Tgxg0Qhu3I/goaO0WaKdKsgNLfnPRmi+JTlRJ8WJ2D
mLE7hD20dZO8Du5woRhvVem0S5T0kr0Tstbvg+JZ2Fa2zJlUUjTahyxOMXItPBfU
mZzb5QKupN+oenkym3iJxqOgAdibiu6+U4WO1knfQnrCouAclesquluJxi5/Ox16
cYJHWALHbyQ3oULQ1NKAf/bF/tJVsWsPitgN5uBrcdcUa0qSt3MyN5OUOIMwfkgU
axnrPj1aVqI7qAbuCePSC5JZ+W+mBDov5xikdLg86w2IobPkffqIOcno9vu+vqKI
E7c7JOEfk3IF5FeP9BIr1KS7faXIa+u5MFYEr8Da6tfPYzBu9RWMi17+KOxjdBuz
Z6H8I0DjlKt3LdkWdGBc2KQhp81ak52liY50Rj1i8rcZ+oYaPjwrWC8RtpEjASdL
9yKGOUMVLqLFAI1u6Mmx3CRg3xS5Z+6a0xLGtC4/MOl7AU3q+d6BFxXC2OTnIgvC
tpnjD45/D1WjjurcffS2qSZknjbjAIcLqiOwNVpa74HFNl8lBE7fS/ZDHCnHUUiC
xzkQosFlul0r3uBSZw7JZ9lxeZvfembod2gY4jUYmazzWcRlRmX0ahVjQk/lzccr
0FtkuLlZGXktEcWKz/9vZ8SnTkW++vBseLTUaf7H4r46At9PjT9dAD8iflkITJqV
LFvIpoF1CUGuiCmq9ovIgCmGqm/mf1L4cwJFchTs/GASSFCMs8Pvvylzo7jR4/J7
rhCs7Nym3CNIj3Ax13kpjqOJnBFRAwV8q4aua1E41gzAm6RtsbJDOt6xcRbzqNXZ
ZJvTHmgCuJNsaxRrkkrhpp2vr/lfUnL8D08TzZu7bbTDcNHekilyFiwxlv0E/ttD
H73qaI+gzI4rQ/WDavifbt9hsarUWlxHOLgePy8+sXwHhsdh0Qd0WliKnqMD+ClJ
eAOE/gb+uIUGCvQUIX8J4/PW75tc05ZLTBitsI76IgTsqW3eGmXN0FyFVzBDVk67
DtWcsEUopBSDeOJ7aOBPQEVVZ5XCOZupmrbM8/SEtvaMLpGxvXzFdemLRkKdAVsw
8Fq8/4YPcZD0SFduf2RiS1Jz1E50Y/iSXWQExT7apL2Ziy+eKKTaNbxtfZHb9VhP
dWHkGWAbiuyPTfIYPtXBtWbVqLCLKyEyIgjpvvu5kznk9cRfORq88Mwo8Fq9WZFT
c8XuwtvZljuKiy7l6Nq3+eudMruF8eOSMsF9HT4EVKj1XBgYiXDtgPboVrKE1/Ak
dQyzO3AJm97QXb55CZ9/S4PycNYJ8bUIWpK6D6vdO93gEWeKXGKh2sHqbw+KzZoO
w1gG2CoM371599u9UXHXZOVKyW8WfD9DKB991HmBBLqKNUOmW3kxkXYpciZE15EU
e7LOlirNytaCVlz4rSRyZgExPdXzMuo5uc+YvwTJ9OurxOCmf6AUKy3oDJOgyX60
11Nc7iQJyz+DWKrSLdQcMQUOVOti1sNw6yzqxJFjFVa2WbHkI7uN7brfHMTnfCIO
zbd7Ws6xkCNyPmSsgmMtoPqEKM71MlpbwA8Qju1B/uYirOzyzi9ZL6bcL1I3bTXG
Zdm8Zp7QJ18PWrj5WWHT80I8rHQW+31MqCBEFGtRlQCLGHoLayArSLF6/GFtYf/G
sn5NwnrIMwX+zO48hd0nUtV2KBTkzHo1nrW+OTwYmc4xlyF+z++FFMHW8dyRi1/u
NavhPaQwlwi9sG9IK/q0TG/dqIIx5yP6CmRViVO+DUXW4DDMfLN8SkK5ZJnWPk7D
qG4oijtIq+XcW8sjDwQe/7zvwF6NK3BpWvkdwWmzMfOTpNQoPzBtRJgfXE3Eebkq
rSEuJ1/Hr9dy0C9b0gsJRgkLq+ka4kgHwBY9XGO2dFYrzgrZN7eL58+Sahhjici7
vBmwlzYKDNZoLrsaZehDyuM4Ed/AtpLCQ33exIzJsOP5CAXQBAj/BqOiC4Kdw1U6
EfzPtfPGBMpOliN/gMKMlo8MV3ZfOQWvGJ5++wkhB5dyrc6v4QPqfeiWqJR7x4kD
EcA0wPx/bPohLyc9LisXA79TVol8p/s568scPDXDtLlqmfpgGA0S/7ZzXQGEd1RK
oModHpJ6G0VdrtoxseKUr0rI/OaMsiT/XPsDEiuaLDAS/uhOIboOFaHtftmfDOom
AeLTihSzYoeOupUgNLmkvlXP4qW61Ed4/N1WSxiJmQQuPlfXK7B3sAPKqY8B2wcG
7xAMyKg2NU1tzhsGGvM5Mw3oSi2ekpwgYYU+m0x+O3YmENsiLB1ndfZ6xRlkQHD5
0bRfoVCeM6N24AidJhmn69l6Jxc0Qz8B249anFOgj0WZit1W+vOOZHajTjLpWb+d
I9lh1qEJME0acko0hmsb2p9bmMtZvm2wF/NzRK8XRAvagHyZ9jjDM8kdAvYHwPkr
Q5Bg6ZNnmMEup818j2miIq/C8ye6weUxqCrNeHmwcSRYIjtD4yejb7lodlezSgjm
fWC5/damGklcFJYJ3lgXC+I1FRv24/t+OrjT4gwu2Huz88leJZJawspA3g5fBDSD
EAwOjOcMeyyAwZvS3BKMk96hqzO5OwDBlLhtlNzUo9OaEG2e2zXOfEiM8UbxKS+q
g1xmfKF5CdQaGq2wWix+Ezrm7fof6OAytVzH1NnhRMQ5fUZWCOpuokc6lBpqGjc9
dOl5vtWehGSL3LaYrvB5YPEYcyL361zbK8prEectBTeUUFKUXIUD5dILD2HorTsS
llAofvViyPKFAkf1cEjzsp5kaGQyktymlT6NZmc6zlBQMEEOj7jE8AwgnnCgaZ/H
zlGPC2qQfb5muj5gxJzFNY3BeeUVf2Z7yEQvcCjoT6Wrzzn0XYq1fTb4cwAKBc3t
iGCk15/z6jEn61reachpQQUJmx7FGv8V+07IMLfBInhHzQpojRZDv8gm4ENEMe88
NE/bazgMW+7uu9snukB4cLi2iEQbjz83uAzZnbajiZxOHsSqUu7QEH3/GIwF8wtz
0+u2YOHBurlW8ZMKYLxDv+trgf0VGidnAlOanZT2xU3z/MZXs1X4KdkDJi4THoAI
Q10/Rve2cn/ktDPMF2JQW6d0TlJANlIUGnlskWoUuuetBaQhUr8mAZfopINvPrii
ROH7cCGAgA+5U5DkR7Y9x5OfDQ2z9LQBeAscRe6Y7oMuGF8Gegf0EfAbxFT/6tXQ
Yu8W0Oe8Q79Qjq0BV9MRPNyvJZcK4Y9YiqvzwEddAJHNIueJ4jRkhOokZgx39D7h
be3r8aEzM5nESSmCF+BMA68cXn+WeKHPOAHkT3eigkJleJsTCmTfqlkdjL5pgUzL
5n+0iCE5AgeNEknOLgk8WQEL5TOvinFLyzTLS3BqxuJCF4DGjk3NsOFfApc14mBA
OQOMkxUxth5miVVWDraQuoIZhs106DjuZx/HIwv87UT4ic2LFc/1pWCDi+iSzHlQ
+uRzvBkKV6C/xaXIjKHMgjxI978TCxWZDyObUuOPwrsUT0f72waX4DBFrMBL8V4a
tYhLkLX3iCJVGww4q7wvo4C5leLgWzE7WPz2qkkUt/4ekmV5I0IUFNZ2oiS9UwXY
1WW3mZ1pJyPA9pS/HbVjibj7ufxWZ9BXULMRQxjDiOhgTQmsdVxxxR6Oes59dLWm
IbKmftnwTJjN0+XDQuO2CCX4Zn0rpY7pyHorPhIVeaIc4ibmDISB1FTwcPITuwPZ
yQPubgyoiTpuQf973PvVT1ob6yyvrh2xsyiPDiFhe2WaKsVt0Y/jUjMos/9EdiD3
j0vwe+W0FVrI6/QRsHwUf987W6tjfvNTLRI7ReEUH4E5ofKvEQTEu1c+yAkQlZYi
R9L8TCy/uqXuZayKrPLZDnKEotxUB9n1X8nNdwPl3XGS8UlYEOZqRUxqSTXE6ivg
BGIBA0aBScFAOehT9UosVdxTLlLe3tro4Qphj2XXuwd7uruPpCyvCGw5GcVsonB1
HawvL4/DrtyEZq4K8Do59xhDUIi7cJ4hfNUpRGg5Fql0fLKViv91Lg16UWQqxhQ/
kPvrTfU0rTTz0c4cEUI9d9C+pzjrlNc4r+ChEdagjPzIX978C1KJbumdSMlitmSO
LQOaGkui26eFB+70p6BGBcbljdhV4Mmoed/CQz8JAAXvT3OYr89ljJbngwHV26WL
JiZAUzICFyYxd6Xpe6glCp1PoSxhoaVvwNbz5cYic7Yzm9vSEzTaFvGHqpXJnEmG
leHT5KhQmGDUl+ekZLa5FfQqo05I2vsGo66NPMOuvNJQnsSKqTwGLHAXnen4XI/T
r/9ajEm/dU7kTQQeqo7gZASRc/vV+av3onxsk95d05CkMIMW9NtdTEVhrA3Y2IBZ
WYTq+zeUV0CNxGWzU5JKWp4yQIVbnvNl/2xt2vSv58oBJwD5u/rsOhvYw9ysBCfg
kxrvJ3Pbj5CWrgZZnFCqrKdVD8GNCI2d8Wd531KreMLrBsyBk8hyf2F5ju+Ipgit
aFff8cvswP++30Rm7MCfhYQtvQwwmgjp2MUSKc9gw1GUWJItneqIXl56Lr9vToBn
bd9o5TRJWEUmFLIduswE3scWFvxD8rl2/uHev6h6VnumjUBTR/xt7ULuMb5NZYK9
zGvTLvfAPJ34I4b4z197LXofd6MCunNRKvcOmQbyxeWn0nPxM+CNQmT6J1W0Qu1j
G3wBcsexY2WCkY0iMD9YDtHQMpCQ5S0hYTOK1O+qzUkz+8E+6JE4CCTzkNSPUPoL
7H/947zgrDa1e8nzig+seUL5G5dZjU1PFCvU868oeXe7AmJNFnfKzeFI7i+UL0xY
QB5+i1crjNMpq01FEwelmRCQdeYvyvUxmwUqX8MM+s86G+j4RfJfKT15kFWPB1AW
4YjPZQ1BND2SO3AlUWPfZ92mOhZ3cphEQAfMCSP/z08migQyF/GfjMTCvUvzOO7P
jjYEOGzlRXx+hMyUpevJ0ZxfDlb0nFkF+UP97I82D7HZ+MqeTyL4fhpTNApfIwmr
Doka4e132EDiQA0Xwp0EKEmCAU/RKa2jdQSthTwcX1UAIJe+N7KebsiANSZDlxhs
2/dTW8MVCtfsSBlc5/YkB/Ju1HzoQWqVGAosu2WMCBRzmhRN8e8oQM6ifg6xQ90A
qUpmTngGQgH0Kz7Vx3DSulvLfNPv8qK3Xgml9YfaML6qcCEbzujzPne+3eRdWT2H
nHJFV9MfL4s5GyHxJGJsfJpcxkYI6ZG2Sj8ag0HWY7aaE95/FB178xdAN0tVuPdW
RuqDz0hT1Jkmt93pfkB3s76ezGzi+CkBv/dzjuO3T3tHgGpIG/yUpqS/5ex+friI
24Rz6vaK3X49m3OErNsp63pRrY5q4GY5d59DJSGbX9ReoMmN+xBjFyJftHLJkOR1
9+H7NHn53QhjTiEKjP79akrkcZuo4j2VpVIK4E4nn6vMRppCQhfSScjHpafNwYNq
UO4sh9+NOrkvjtr2ZCJtuLma3khux3KZFhIRl7bn/6H/NkOle63fMxjTIwLDN2nx
fUaxHXSeLvFUoBaisdY1gQgje0vc33g5YHluvpybvfcegJnXd+EKWJDqojU0SQTv
vHcwtBZC56VhSAEts5RHcFsMoFC8SbB2Ctfr2844xqSevhKKG5LwYxcbG1qKQCsJ
O6XPc6Mh2oP5ne788bwQcJ1p89f9S1GH6jnGTDw8n22NDUchaVNU2za8KKYgqrbi
77iVDzfr4eJtZE3+W5aTpB70z++KbH+CB/Ug7aKGinQkBNVFCASZyDpBgqtSXQCm
KQPZEsparyg4jVetUDJAOCjTjyWYRJhNOAEU74FjxJPPJM4+i/jrBwarHl5zMIdG
BimeKngNhlkOyWut1gbffFl8LQ+U7k2e0OZpAbn89dmRL2TwqODCACbQcEC31Al7
z6jn8fc7QmyBllVbHDGqPIicni/E44I2JjnwqDpZcaV0E6j+AC4tFY0v4hwk/zAv
kFE4NeiW3T7byMmf+4SZ0JOpSdwQv8xmcdJHCH/dOXTgzoFkwTEncWa8XCWO16RB
EfHScJKO/0//gKjud/UHErNUmmswF2d5hDhYJnISV2Ryg1L3AWxzUvnUxwBEPLjx
vhAGt9tu+lr4vKbGPJg8QYn64Hiquy69OmqUYA6JSUpvLLG9eBaHY3eRAGz06UUc
Dt8/3rjl5RwYZNggPE2wjjvbJhPmuZrW6o0BL2xHO92p8H2YC3UQzWpai399Wg+9
4YSZDHYvCAbwZDZfPuKnMlo/hvTMS6e4SX3kDT6RpuMNQ7wjBldsHwZPR4j4qdLl
w8YWdoZQGxREbgJ8sCseCYwSdlqtqQFCQGbvy6RTm2OT8TDTG313mOsHAzWePZvs
WRU68gvDapZMsG+kLs+z+be39H7jXNn1nEr/aCvBhl54hnjSgFlDPZDtrLP+qBnc
3er0zLJI00JOGdYQjkWDp76H47TesQNSaNvvl/elzHN9GuUjH/VcSM5K38xJKve7
A/+M7LFmm0VaEKbzh+pFlIZYk4o37cAmDgtm+DXAepepaFzqyu9Ql2RxF41NbESf
8rV8MIw2XyL9fu2aukwHcafNugq5rv9xKCwWbQdnbeVbaG5L+LCavMj9HvWvdkih
uPRgg/wPUiKM9UUxo95dxzYs3MOD7juZHi1hqSgLOBOs68kcbzSaSJNbxzveQJnx
cMEmm4LEGmcIWJwd5+PE1OMj43iu9x8nY6NGzF/J+A8WXyHOTnopAkL93U/3QGDs
yXcM/CjaAr3qWjbr32M+FXLb12J3EazcBK4vZb/MiTMwfufSqmqmLlMw6EdH5yNh
JCYFhdcxkwcg1OqZf87pcPvG2ZFJwqTsdhLLn1q8V1OWARL4JJWU83ojCNIaqsiU
EQftwDmzoJ3j4dZM4iNXSHyJY64kT9/zYFkxJ6Nh32BfKmK6so54mdUKwxfzo6au
Ee6OOC2Pr6nEtIDGTfHD0fWcDSk4LzT6ZaJicDmWUBbzh23UXdi6GsPzb229Xm6Z
0R8iOBHftjqx1U0ARW1Yn63tJfOaCQAK3USR5Hyd5PWx0IbVZFF1QPXt9LYC3C83
pmqMSBHVnghgx1B5niwGK2s4+ZmoejCPTU0swVueY1Gdyh0J7GPA3qDrjT8oPLSv
AbqCKVqRPd5TnC5+kiIJMqkrZ3pQDBBm3hv6wVNdFAQPuz6KpA85lBmvzkenvVh/
lhiB1VcnZ7zvjCw55mOYyxfz4gTOcrXmZgXXaA2QEktTnMeXoyymUxTcYEg4W24b
hrUtCNHJmO4YAacNhr8dyTmVGPux9tDn77A5fIrb2ZdZB4S+F3h9Cg/I8/W/0vCP
7Y1PNT6RG/SLx67i70Ho8tTPqi53pBCSgP1OEDDX6xYuczN7KM1LjIx3O3EiH5cR
aVGL8RkVu0IBqOqbz9OJO3O0aAohWbA5nX4oH7YapElWV5Eh5dl7MAZQJ8y2sgDG
g00KFTiqFdFxqbjNPJ6Y5OKT920Q7zxaZ3Zwt69KB4FUOIasM+MZFzsNDLqmM2ph
8RCdpu/nSR84awY5f7piGUB60fc5+6K+6hEYe3jPvOHUvVdeiXR+i3KLZUUv3UB0
QuVoSIEsat6ybFrVK00xEmNUfIgMy+pQ1b3iQGbQoggHj4WuB4PXfJ+v2gc+87j7
J6sILt9rBydK7kAcCFSGrpFHpbd1+t1e8ffCCZr4anSHGGnQn3jWJrVLJO1wekAS
+f6DaKu7ughp8bqkCarZlg5/g4StfI6HqCmye8j1Sz9Pb4+7PUl/kl2hmIo6HVPw
k9HVCvWet5pYfk0atcXcOorFQnq6FTEQTHMm9oUsRpMv5PZZ3h8vWD12TRywjEL1
ejzB+bxaNpkV4n9l99jqoHDe+SOLWUX8crYAILDO1QHXMSfZro1ThZMxLPdRyeDJ
HRB5Pi5XItBaN4H7+GkRMO0TX4TnrvAI3T8e2TrG6a9AaokmbpbsKDp1/X1VNfzz
0gJ1H92dHq4mkvm47lb16JbPb86U0K8Uo8HIIbr/OjcnOWcd2MJv7j+l0hA9asHF
1j0WziujtuPARCZHx+/TuWsJ764hQJcPgAZ/zrFslRVcn2tguW5oHNocGHVZ+g4d
7lHyhWEfUaarrYPOnXna+2yiE91+xQ0VTXMYXyTRgEURutEQ7HLzWjUa3Z8otBxQ
9V+van815L1cAuRdCQiuM3ZyhWe1ekehgmoKNZREwWpVwXD+n6ugAioL8yVd1P6X
9ijbVIAODT0YiPycgBcxzoN0rcsCJF/ClXYqxWqD387HqhJ0g2hy85qXoYPgJHXq
UgcfIe9pv90gbRkB4HoLfN59V12FNfIxDQg+5+XRmJQyQ6JHhJQlPty1d/FaRQ8g
nfdKDy/TOA+cXIDWxuw3AmG7ybcUdtocc2SgKF+a3eNL9xpCZeBlLyFePsOzIn2b
gz0ahgUXbEyuz6RjC0mqy4m5m1I3dpn0RV0FLdJPdqFsVhNQo0M/fUBeauKZmGc8
L0k/V6EQYb3ZroeU69FEbISbJRWoee2EuyQ2Tol8nyal7DREFB4u5BC26Zb1outT
gzHSqZJmBeqjF4j4Rh6FncujV5OjmGUkTEoIyZLugZn3yV0X/ebuGV9nWY+zp8tS
1zDkEgaC55LVqW7Jngs5ejtk3o0zHZ4zd5msx2K3IT/DiRE43TY/q2Mu39KDryDb
DVfeaHS7aOEMGVrQd1GYvmvpOoSXeD4fnZB5L1QLTMFGIuGpHaQIlRFVzGw3xO1n
WFesqHrWcGtsShRsSzCb/Cg65LnDEvsAFgDG/HU9jUwoIwnhANEcnlHjG4ri2hAR
ORpvxxGNpPY7yZaSPVeNo2gd9CS6tUdCaQLNxwIWg3yNyAjBVbrHGeJy5i0kd6BP
cDxyySuKn9+CsC1SAvw1mdr7SgbT0DFT1zqbox3fh7hAGPm7sbDTrJVqYNC05wSF
A5rwz7CH+IvX7bkjAxhEfzL0xDTeudI+xE03SJ7zyJ1+kkIG8K/oMUVIc9UetYcT
hZnlPeWqcHXdyL2/ozQHLXLyM8OQxIrQaUfZ+YdNE13cwYC+PBfjhY7a4P464gJS
ZiViO8N7lsmIeIrkFKIfT4NA3FVhBzUOEaLnubavgZMo8Xjk3ChePRwJJ6dChxOs
g6EXnyDLa7JYqZZxx2lXh1i/10a4MK+GtdBX+0uaKjO315lj9famwPVzqAFxocBg
Ma4CNUCEJSyVWxiY9LQqBFJ64ssuqxPrbtLYfGV2ICUAeUrZrtQiIH1FJh0aSZw3
8K6dVOD3+ecMjceXyi7+Ubd+rrUZ3eVoxBvdOxA0+ZHoJFlwRAPLJd1C/h6M/mC5
lioopVrg8pXdejZ8i4ewAmS30T5hGcwwoqXwJ6Q3MChbz3ayxxJQljLnPBebloXW
g9UoK/lPaVAViBx2g5euLtq72x6cqLbjk/Tx89TYjv1ivQysXOi9wgNrTOJMVSam
TQRCf7Q1IDzw2Iq2p9WqDyf3wh11gMEtp0G2MzyhOq+Xs2E+EK6VUcjnnY7BjMKU
NwZkCD3GLio0G+38t/w1o9MHiFXQ1GmNKgbi4tPk9y5hpdlWGubrKbeK38CYL5FW
e4nFo9wOxVfm5kG6+qNS6r8jlAEQCA+B90WnFDOjKgcvSgk/7io9WYFFqXTMQB1u
B1ZxcabsMP5904veSyH6Ib0UaN+zwU7LUf8WaoXOwpcu8ddYQfEARfJrzf7C9vjB
CGHtb4SHxiMHDUtwWvNHnP+fhnGh8R5foHaWhJgnkI1HhtGCiwarswKhyEGIdOZr
Sd0jc2TkLa7fp150YqhcljinWB7RbmBUU9jMAbnlN80RPNou7944pYMS0gsBLXV0
NRRNaRLnoJ0khTBU9LgvQx0DeRZKDoXSeV92ZTUwTlxVwJuQ51fBlcT5sE+1YEhs
7pU6duQchNx/tjxMOuwjvM1wG7BVZEu85kgvDBtirQU4tSfnPZqtT25ZVETf6P+7
K8G22USpQDV5U3/aL6suvvlHiHBpHK4FdbP8JSQB+jUeHqe94Ih/IXAoIazwPrvj
tG1a2BvQ5FxfqaNP4oGPUMiTkpavPI20WlPoO9JNr4zpamDmK5tTR3RaDQVHLO6p
+KpibuJxWbJYp39Zupy0kfP1xpua1LAQ906+FRh6kYf2G13IOf4FAWK/k8oiLNYY
imh5QaObkGlxxPK4NFchMrT7xF8tfeJ9DDaZE1BM+p6bagGg122jJ5S3MW9Pqrvk
OO1/0Isi0NHAwbDo7MMRxZ8xNY6NQSWAJByO/1OTkTI6Bv3B0svKUpWIF4jjtXb2
lvYDiMvEhl5RAPhWc34RQC0y2ZifHH91z7W+kUMkPhwj3Q8qn+GufcO+2jIDdtt2
9+srXcPT/t6Rp7pKIiLEbBezhTvW2aEg4sOHGbXe8ptDJxHjqewbr0fW/5wojyx1
cB1uhvM7A2ZebFGj41r1cpHLYg/Yn0aRFCuXS+IGOA2BAnmiIqRSZdIuCdQ20zlz
m4Fb33MWBnfuGhk2QfPzyDji+W7vQkbgMkwinAtNxXQov6r+x/XDAI6x7HpbjtpI
eJKyBrdiS3/8xLWeDJjSEOWHNv4fq4ZFd52CjvA7v3p+Gv+2RoWn450GSiG3kMMR
w4ZXqCHEXbuexybfyq2SFnpz+MHK3c4M5DK36mrLsuf/5mYQixlrtriofxRCnycF
Z+GDIaJ+6LZ4FHiLyOy/pVQCY2U2GIpwj9jzYzs9ZvlrZwLUDjg0bDz+9YeYHZf1
jlSvXKg6B4swBuC4PDGnHYBMaXahsj5FZL0yCnB4kyGuvUUmXodC6Op5KutfZbKI
Uf2/yn064BbKozKOLaQ4kWn5ACxNiHEcN8yH03Jq5b+37/kMFUzI7gcrS/Zv9MYd
uQ15o0avttBuL1t5WbKhPWLNPyKQVAPvcdA386voUr7Wv0fjvJNhbNQa3KpJoo+t
NBppZEt9ap2VxHMl4LxuHl0v8OPbhTyJxUmRdmffYlcMF8tz1LkhS0uePo8N8GmN
rF9KP4dBOw/jcMgziyodoxLzy3mineLUR0xgDn2OPgKzFRuo35nk51/qoF9yFvV1
98RtnkucV9wSBV2C386oc7bVgl/A7QthJ1qVM3FarUufb2/DSmbeFNBPEfFdoxN7
cG8yfCQhtQL+IxN5I6W21Vi/N5jQPvg/X2hBdJ6VlEm+SWbUcZPLyxaXTAPgZBuE
bgsWqP3ZmkThxaDzU4Fz0cR8zdb990HzEHTIPaBvdn9stzaR4tqrumlVpM0nm9Fq
waex3ds176cN/demviGpMTGat2nTCWHdzwvmoiA9TuTb4YqaweHgotGIj3rs21xr
yaGXSHwy2uBeY/m0BXgoul10Dh/W1ZmKT+zfElSlRaVFjME/yXnP/S7ttJuo83nq
eWflCnICCSbrMLKmKnvS9nGvFJHQ1zh93iYedamIs9qFk312ojAtAWCi4ND761sU
jv4TY7ZRPskqzFUnDK29nj8sjIOiGQ4XT+jv0pcaQSZPatoE3vQLXuzeAAFkSV50
OvLEnRxLhwGx59wev4wo80rrDiMi6Sl4nQPgFOVUMvr6jvr2msMFUeSg9AWRV6k+
vRCyBVHA/oCMn7x5GkDXnDrMJwG89/597ooPhSYYKIWVMIAve1t/wilr54ivHolc
9GoO9s9t0sBC8RN/r+JXyUHZWXyb2u8/HnZKRkmEXQiMZFEcMXlwPVPrQTyAtzo4
1853noamp7g1sTWzGhNMqpjnYS88De29a2QefwUWWbo/CUwWnfCC3gyfOTwHDaao
CB51kpiOOHXSMP6RYTK4b4ih0LXLL+LSbkjcZvBqbnX2m1svZVDhq2Cig6nzqv+G
EP6OFtp7MccTr8lI1S9HmIU2+j1AriG6ETOABYeB12D7HFSuusgVq8oi7w3NmKCW
258VdH64rz/iKNSLF8Sdl10jfwh1MbUaIk6o4N/8JJTWKvmIuxmH8C3J3GpJxpOu
8Sy3Y2OFfD7xCJP7dcHdsfUC9IGJ2AqTEIO9pJX4w8ILOiqnHjVJPNIyXhspNdpq
L2n6WESEXaK+dTwwV+X7pSM+bRwJssV7lOEyjNnJ6SJ7TIjT3BtaK9CKa5xh1qYt
4uA/YVNIRV4O06ctF/QfbzU7T5OBnom5DFhiHY4jTRme2xpuUgFOP7WQvCr27xjt
L9DDl8wShvajnN1yT5bU+XKmbADEqprb1DGc7j+kK8SxRn21ovEjWYx6hfzrcKSD
bp2lxy6viHgKsMNeUow2K5frVzxAG7WCBWwU8BJFrFLu2cuhyIOsbb3SbFzpLbSK
/w5hjtJibWdwbekIHpYEoY/+D9dSeyePD5J9iPyUMRjQtS1HjMPBl78515rSvGAu
pWZ+KELrzq5bItuiEegySf5XjDmRPafecJakQqU4mWieEtwlOPlpgv5aRoVk2tIt
XcdptFygHPKF0qCPeLWWHUikTGbsH638sqSESzj7f48PHB0sdhi3QopJBVCjmLh0
sZzOUW814m+O89FHQ1Jv4wgi/OluagNpmFTzFxAFUSTsix6GwIi4DbXrqIqdvKYZ
CZqqG7OtXMHU7kau2j9cHk19TjJfIB1tZdPprMyM1YsV2hi5MDlwwZZEBKfy2GT2
01tV8wBtD6x0gCCR3yd5QzrvM1ygQ9VTKL7iYyNuDA0t3DALYi6CXUMvwcWqugwz
iTwIKSsxkJuduoMRI1Lrvlp0TNYNKWQXuLEEuTTDdD+pPGgquaG63yqueamSMkAr
kSxe8t5OEpR1qcLmieITIYKwU19bL4of7GySNwG/Y6HaJvcWtnD4IjjdaDCrfeI0
NfwASKz6X0HccibGgOogqELewzPtNuClPyFN18qQQG01zYNHsOG0VoZKDqZykd8m
GS1NvzzaQpeNu++zbD/hFCjl3xcFi9AVG1odEzuXNIuKAueWtXFkXvZ0f9Htbxyv
cWmEvznw+M2Dg1egIVwVXkR9Tw1nT034FFaGUunya366+tFoDchwg2nr/4q2Xe0B
vPsz2xi7VDbLrjwtnswk3a+BUjwZXafzxNDEmvFWIVmKz/HFKTEgbuGFPG6c2BxK
PnJMSpXnSUd5EFDi6Ogb7xiuHUHBa8TNo+nCUHIHrU06szwE99B8WMmSpUj+aIPG
q+/GXPWM6XDtixym2aYgEaX3LW6rpKk86A2C7+0miOK0kzZA41PsH4T7dnMr/I7Y
UVASdnxo4t03ipRiePBHdM/QkODiTAIlgefb5WpvQyU5Jwy8LT6l27FBoxOgXAQ4
F4EbL3KBrlIyvgsk14/8WYzOrzI01/X9opi8dISLMgtHiaeyhhgVNCltF0UROfK5
470DP3565LY0ew/ykhenz7IeiB3CyJKaidQP29Kb1n08syaO5TW63JxmZdNKW9Xh
k9qteKsBbCWdImFMT5S36uTQKe7GeSYpBjh7JlGmrgoscCIBDjuT2az/MsRIpen9
ab/r6GFhMTv8AixOan2vgAt/lSLR7JZhrOnM2Dru9Rn3iPB6B6hcR7Zmgb9uiAbN
506+uRmui3VjmSC4RoYnhroHlYlNUG+RsVIMYhCSvr+TUbeDmqGstVxovxV2Bsw1
mnDUsIkzwzSmat+LUH2yhJiWl+OcGAAjzpHIwcV3mEV90Jvg30PAtG0QHc+SZOrk
bwVAN737CvZr1kwsjNUdCmwdsQ0Ly1COocVcyNqO1j1ILWCYYpAP5ghSOD+rV3Os
tGe0V9Tf/nXarnyUtFgR70oesnJ06LScu7jJJ/7jtgztQ/DJAW+duZLG8a/Gu4Kc
wlTtHC7UluKa13wYQUy7/ZAUUlhRIB/tbMTcZFMGt9ClBJg7X1ntzKrmqOf/5fL+
HQRYIcLJUIxKxmt3CuaSfCnaXyLA3SJrYbtnIXlt6C2vucDyW14/W1wACzj6ZR4y
2tGk0LqauNJl5ofTOCw4V3RgxEodTpNPc4Gv/W2jR67H8zXe6DVkIQRdrQGwa53w
4gsinMQJrZeVkmnH6VTXrensSEH+UQJkLfaZBpzDE2MA9LgQ6a6ZmQv6wWbMNd43
v2Dl6Pn7EAbL/ddxBV/r/xBQULoX6PvDiSMzLh5xGsciid4wWZSXk7YPcBULPRsk
rMl+OuGKebn1oP3eLjJsjlRCf8nowlPlS1EvA3OEpxXlUVCdYgzice8RqwTFvZ+y
Bz2t8Lv8pNFQZmd1iGo5atoC45syNHqELt0SsSgiBzCtM3lmLVKp6wleawBkgvTE
ngN6fgqMJBgzWirNLilnAzb4vB4ycp01VYRHNTwNQaRzN0bSly3vFfff4D+JYxd5
QXS3LmInXtdB+qhXsYs9gLmJLRZ/W210ywo6zT6lOaGkjTd5G2NgJz+vWCot+7tB
bcy8QWdcB33Y0MIWzUYPkJBwck4OwUBILU2n20gvoGAcb19tuSkOgENokvhSd7uy
fEKBGNWC76kTjdjP3b+a06tzZ+pGy5kBgiEsbiv2H6JUkV4usPj0EdpmaLFyMtoa
kogJK28ygH+4o0W7GpFNJSJvmAdQNsBsa71mWY4YNUrFptVpyo0uJWnVeY6el9vI
5IG0ObkGfneFMcriulm3sH7pGMFKFQ3AyEHOFN6IZsRM+dP7pN+sQWPsor5WOsLI
7yQ7Bqv1SqgOCuoQDwk4qeqQLmZ3I+vfKnMJQ09l/cshC5kr9Yb1THna7ayRfZib
L+LtGwa+B0MKTmQAmXqZqtJzxo1ybUhM9IO9OLLBH7l9P45a7epUNCKifuXnibw+
ieBihXWpIChvZObi1Ag5x4AL7gKsGTsl8art8k+AgG7VKmxN8/1JjGC0haEPiuVy
LOgkXuCeW4kN/RUm3o70cHwZ81gZQR406bgYUaj1ulYdQ2SLZAeF75VVrPmzIVoN
rgFyuDN6kmF7ehThmgBCZyKvz5nvw8Qflk+rAtMJKJlVC/RxhS9geqDq8x5EgBo7
N5hzYyCKsKiHeTjqqissIzqYTk8lThcpfmn5rQTOnXzDJs/05nUKdPLC3CRTlNJr
iHzzOI0XsZ6Ag8/kCOru611lcZ6GZlYPuhG/gSrgR8dCJdsex8wV9+PwtdFVlMgh
33maB9c1BkYLiVPsb1vMGE+qfGrriark6RpGTjGO/FBXk8OTZdXXMzvXBXQBOsFB
AOh5/6HbErNZpePzdeqNk+OLTYoMum/FPGBCDtomho5SqMxSxLuAbv9W+7jrYjgL
GE2md7g6ZR9njKFGykCmePLdVknKM2EahBqcqM8XX9f2bHEy6YRclHTzABLKGttC
/+CD1ieSfnzqKaz0fZc69AbFfmOMUd7nunPkK+Qjod0UZcLUeMQ88Nnmq3Vys7tS
86Spy7tZA/lnZXcq9XuS6/kpgIBoqXTaPfZ/lRliEDxEP4AbX6KriKCBqZS6AgZs
tY5qzwFAOWd0gMptRzs1bnvQdWFyG2J9uqq4NGSwQDgsI1c8SymZRAOifRB5Xahf
gTRE+l9qGMVleSPA7zPfnuKtsIxED1DiMOqK3mwwlFwYlvdQKd7CCcv3JYauoEMZ
an5A8dTVLUtHiaurTmiZTHHngMWfbbMcHz9j6MJMIy4aB60jDezgnFtGEeI0Zos8
aNHhY40EU8bc+d5Tc3JcTlCgjmj4e+QUXVqOEMU58R+PNt7qg8N1Y+yTFA88Z2iv
apHZL/f2H5nplUisNQ1Ht4Cuz8C740vNbKpnrjJZjw2I+XTRP1l6E+BIjYWaevVR
5VtofAN4LI+HIYipVhCn7P6ZmoimIAVGdb/bEQEKVaELQSowRiBJYoVwu06WTHrR
oipMcqaopdPNSTfECfTNi0SNPBuDfIUs+ppTgV3a3eH4Oh19SXBartROWDFlqseg
z/dw1uiMfqj7hlgHB/joxgzl/dzgCBUf0pwTdGTjhCBwHzdjfjYYYcfrFuwRXaew
HUjD85qiLCUYXwZVS6+6EGb6PJjEPSw8W6wGh14A3p8S0zKwKZdMUBez+acO5mLp
BGHVhoJ3phk+gtyxGoBbxBar8rWsjfG1WS3ve+6kKGze34A/20fSUt7J2yDDz+EL
Iat3udYnlOzVWJHhl6gXHg6OwvomWbv5LKwRVBIxNNEpdi3QlBxNXtc8GmEIvYGG
98B+FL8M361jnq7GjjpEqXxMGhBs4238OyfxgzwbFdE/luV6VHTe4psD0A2qqRVi
jgauwMrMDIxkP4gY+9CUHXKEuTtk259covkdQGP6RUHHtEvnkwFCLHeBFrPI3doe
A+8TPU/M9b59hVDQ1lYqUkPn4MPsG9IQBguHyYdSYqF6xfKLkW/JQTfbUuoqUZ1A
ivuCRhabEhJx1MdJSnOW+Umab2TL7LYRjyN8h2ZiOBar6FOIwSNSxYstBTFgaq21
u/C+gkzhVvGIr7Y3XpDHAJNEHyHOh4SoMMVGQxt+w18Gumwvddkedj8ttlZIqJIu
SWI850qIvR8qlhs5zEcSpB5CfQ1qKt6DUKT7QwCYJRRJcG1HLZt4NVBRfOc1aJY5
bDgb/hlG+Jx4WH/6iyj/gSe0q7EKhH+axu36Mssdv+h3zrDpR/AHiAGmp7DZu/Bx
irpegzgZVdhy3FeOLJ+PNFpbUHQhTjLiZEDYSUsbgd5vM29VIeUatYOMbpFTuuHo
TfknXsx9qclTnWB1PHqy0KNjP4jFXK4ADUcvL9T4gUOxQLdp8RPJp9fzMSAdf6Mn
iQ+XNxv9KFZYjEDUz6ysCcqSM705nBMZ8mnGoGYjQcSMp1d92hyardSpjLUPgBkO
vUDwww6YQ+fVCvUH7Tslgf7XL2ZaiNs9CbJ11Y6hdrnD757ot/axAXKFpg9jRjcA
NoHpR2r4yClVTAHosBoFQxKk3rk/TfDrpHvKbqM17YcNXO1Zw779TQw7uXK8gE2A
xmvaCykPtx/koqox/3HbXE78TqOD0/IdAGyHXQIgeQucy9yyRw+JnJBVKkzIPbmB
sOOjlmcZSlbDBGE9dsgK/XZu06gQlbRvG7jKYNJ4LVxZ2eaOXXAYuEAqHjU5NCCg
Y4n8wqCwvU9RqE1Xva7Cr1rNTL7ouY1nAn69jrJgFKjM9MH6Pf244ykMVZcqYxTC
nEmCmcWfyduoWGgWoGSjlliE7iJkoiNMmHk9bX9uyta4YrptYtfU2vAUfYPHU+V6
iGd5ZV/v7AS3eJf/7VGKuuadUV5VXf4Pl9V0Dsi2UgkmNY3UyjrNTgk0sRsw9RTQ
sUnYMV4js2N2+MJ+231iGkx7yVkbgGM7glaTOi+1rAfkVUKqqRKdwtdtwPNSn2lN
kXib+Lp0ZVlIfDRQU1JMdzYPRCEeYazcpcOhg/UKWdJAFq9y1bedwQUaUqsnrzUm
VF12TBkGjRRGfpl9m31v+Eh7srD/Q/re+uNf/rQ63hAUQdCk49rlYX48a7X5Uxeg
i9mjNnq9rh9zBw2WKW+EyY7N4RD89gJobLjXK6VCETSvgSylnKBgXk2/psmejvBQ
ByYDahzqg6p6GS3V3+QlIyQI7z4mJKR7ILCmijE/0N8hV5pZy9+3Am/WvsejnR1H
RqHX0sA1Kr/tXGGdGi7Hh3a4eXqVsmYgVt4xf2EsBCD+vJ+5qrE2E6WOCk3Ailrl
6QTFnrs4SezzPUnOu36/Wxg2Ief8XFAzzICV+v2shYKajOovZQD1XbBJ9ftIBUmB
+R4fymjx4nkGOJzVbO+vUxGmlPMyuMx1Wk7yv6o+ApBzKyfaP7s7rq0/tWKCnxR+
tsR6c9TlOGfEBbDqFFNyx0MMBZZl/ab9wHxZfIBZQJmCAk9Jdtp82CLaB6qi3/5B
bEIW5q0THi+ZBWjpz5WCmBTnmjEH+tT6kWXGBGPjwxIAKMDQl2rEm4RtIKqk1NFh
NOL3ikrBINH0BVNYihBxwL1m5vZaCEp9cJaYQpckMtFGn+SzcK4wJkD0qEAPOAfq
2B6/FkUX7dtMyRRs22MXosJ354jaPne8uZerEn0fh9UzqSoTENqO8TK3zIE64f+c
yPwku98YHnYAEy8T2sFD9OXUwYlK59dddW82wU+QyKJ1EM97lSnxaKTZJp09nig4
N0ppI7NWbhv3dT0lNPNpSxilOQjDo0ld+EkYoNpP32ug7actLbWbEY5hPWLHQ1aE
6i7PmA8IXyfAp2H38y86gJelAoAsrozwlTYkuPsnym2IraA4N1/SR/MOnHADVjtD
aP7jEiUzk7JflbA4cklplUbBXijFn0xuf+OCMsUwJ8jAJTMWQc3+SU+9Rm0IEP5s
x8yH3xFo7gfo3TbQtmd75gpOZUiVR8VndylTyVAMkClN5b99fKRELR0ZdZUtCm95
hn/vJ71pkT6ubNuaDvhEaVsimP8bHRfzuJyA6hYMkrghAkjv/VEw3GRPOk220NOe
Isuf0cYGDHAPAeypwClO4t4G0n7dcHWGgkUCcGVxtN551OToAx8jEQlgMnV0IfsY
0ro5aLYDhYJ72YS7J2xM+H4r2SJ/tzLvNx1ceag9TCNo4ntKa+P/RaE7LbsQuK52
AjfWHmk3C2P1FMD+1uqvI6x5V0x4YwcMmHrcNI9xfD6uNHCV+KcynEfJS6xBTOSo
VsDtmBJYvM/wIn+zH4G8drXBC+sFLy/lKgYvt9XwMSamMrMS0LaiYVi8qaHLDj2W
0LfsnIvbjnMbwQa+F59hqhwjhc25rqgDUa++h31sTNsN71o6Iz8hzIPne4bPrq+K
/Hnuf6T4dvRBE4U4njpw+vQhEgwtDxOQZueDPkrYLQjLBfnrewhvURa5pnoh6i2p
x2MBftCMoWLFJfq58o9MgGQ/5aJz75A/0j18PU+SfI6A1fYah8zwuqk+7huURn1x
74uBqheCQRcTa7Cqx7JzHSceaVAJbGYWJucHHV6FQ9DCNkMZ3ZHjIoTeVWut+bEY
Xt6QS5FsUsCfcNqP7xUF+fr42MuPEOqpR2tIlX3+sn/K+5BJ3TpzFrMt4dWM0Oks
1rx6Qwu6feHgYnHXDbMKIUjL9Zu7wzf2A+vtcNUTOFY8wEP20pMoyPqxQOXYxPw9
faovpY1oTMxHxRNmvjnIjp7H9Jj+4A2dkoNgJaMtMKWRbQzK8lb3jxQnWv0Nmwiy
u5qAXZApBfSfQFQEKT9UaJF/q8pcsshlwGzN0gbVrGDIEA8qYUnqGeXAqb9wqP3r
rfipoHZV/JXBE24LCIKU8BoJ5Y+C8xln+6n4x+MlamF2HX//pBzb3RxS3ToOIfej
jgBULdJ0Kq3EHoFF7RH9ZrhSNnmQud9j9b9MNG/xSo0E/MFD/TMtUpce+B9JQrjN
c6L4ZyB3Raitd5WSu2twHojDomF2Q9isv9Ra+M7vgHuDvb3VIo55lg3Ncqy6yfgN
3aoAxBqq4BWO7W+rOtjHhxsNofFDDEi34Mr32H9yrHWB5aylG2dJ26NTEgrAaXE0
p+ONKGQ763CFAc6q9vCwQNm0Gw/gOipk34sYH/MDi8i5vPCMHyQ2XeqiuUrrrk+u
qJFlX18mzeXDkcpH2haTqX2mdMvxV6mcKCjMmXP/F9rLbom14hnkiT0k+BKb23vd
rqFYWUVHhG7c5USE/z6bGSztrxDGEbHFKUdo63WMal6ictaN7dQLC1OJW4DnVj97
KfXFJzr6DhdNyzX/vSQahPbj3o7/KwNixbR3BNk8eU7iYMritgy9yevRdo3HxfhX
hR2VvfqgyRxX2hn43rFYRQpw8oawjmw5rr5Fs0dF+4OynoYvDJu/+a2EI2Belv6G
P9eDCtsT4iuY9fwo12HQrdx8A5wOfdxYrTJWOdETcikbP+2Z35kc1uivaidgyiPa
E9VEDqCypQRgg5hADtcpivntC05jkyp8cDnEnvE8a96UIjbeIFAKxNjqSNeIzcmC
U/C3ub0ZmXqfgmVw3EZiykpGZk/48dsavVrlAqmL8LfQEjKYZOHjPcOun0hE9gHd
TRjQq5SWkDU/jcjwi0RFmLwgxEm+EEOkntLkM9s1WMH6NBL/apU+LqwaywG1/rkY
y+PD0sQ7p2fFJv6vyOSNGV968hQf77qRUOgUY+oaucjPjPTbrsrDJUDqYzerAHex
MYyUc7pYEURUybvgXtcr1UYOoLPQ3sDzav/ISM/5RQcd6WLO41tnN//RqVy0AGzq
s9ApPBoh5PSH1lWQDp7kL1Tru/yxjRIVmT8LBwIQskA6c2ZF7UsVOTqBWQTZNmMk
csCt5NZB/eoUsYOAz0ahRk7xDJupk8mYeT6fg3Fig5t4LOCVMNx/z5YT6QACXvFQ
uDegsYVckknvZQn94KndBCXGo2ZRf/K+JAwGfB4o7FaEr8DAGMoVkFy4yhI0G+/5
dUqlJUUBxGWHao+f9523XcelBAlymiC6asTdWWtHd7fX2QNp6N9a55pYr6g4lUQt
Qi9lOLnVLnml29R5lla9HIaf0OSKYW6mfib6em2WCESxc7ztQoPwhWjNYt7D8X7j
730BypdEOYfG9DpPXCy1PURysG8ra+PLLYV7Swmlzk/jyf65hVrRe+HGe3v9MM5z
m2vnGd52sZ6rRpYXeiM4v1lICHYvcUdM+plWtggv0h2MO5nuI7Y4l3v3YpsYjQjo
WLVejP3Or40Rszwx98UNKbuZCQim1MepFPVyZLrgMRgIrkoPx2NP6EpGnrchfuJ+
ipA/pf630NnY48p5gzjZ/98SetxnTLwZN2lqwlh/9ienFVsr4hCqNof1F2by3hk1
5o7/TU85+FBRdia1jaqwm78YnwhiCwrYAqZ+AWc6bGYV2xeDdLha88R49my8AcGv
ko5F2oEEARsomPhqpJUS5hOTSMb2xGGY+UVu/V4VqTCkn29K/p5fM4ZQAwHjJ7Gt
XfzokWIHo9o7R8+ci0tXror34EEsbHQru4IJ9a/YNc1ZcPAc/h8dOmOKUNzvuJK3
guh69twrCRgTEOo/kUH5cK4xfluAH6jg/35F0qPvBGi9+I1A2C6Lv7vUZAD/tr9l
tLmiVmcKzIRgeS5Kw5bm9Yiuxag1MZ0pxtz5dAy4Dw8py63uX3AMyemErvpqizBU
p9E70fMqzyLn/0/1qrG0QlPpd9KNouci3O5dnjp/bTCpM8qldTKYq0msT2CBsL9n
8OXZGWwXvFvemV+Ez4R+SHxTMxBOBVVCs9PkqWJqaKSaNLe57TsWR8jNrq1l41Aa
7rEQ8ZNVvyuR9nTQlWc3v+kY1QG+250SkJeT7eUjVGdewCxxsUP+2K1ZsNghycW5
icjl7REzjt9t3x9O95ksQysIBA+xo0YjD9HpdmzKC4iEFEAE/HlCHpH1QHMdvDcr
szb4VxAJbExdiSXpARP0wWkiu10nmTOc+fkuilLmZGjjHAybKlNmrXJ94jzHBuUZ
MpzGNY3a5krFkbQfzWyYZgCHAzVPOFV0gy0pgL4traQ4iI5SxjggAA4PYCRab9Cv
K0ONhYQ5juUMa0PJ1Kw6nhD0U82xxjaVfm1JECYa5xjWD7Y0VgGoL698EV5cUynP
vJpKMzHJhmp31nIAroUzGQuzCxgyT0xBL3BCaLotuMbcXXp+9QJ+s1vXBf18B5Pc
vIGxWwBR62j+zEFXmPqP+owqgcrMr8xI//RYsQcUOgKtkNSqxGwZeClW9fYvw0eS
o4UNYT3qG+jIgTmEr9HbKwKRmdvUOR0tdOqyB1qVftMc352l3cILMXj8Jowvt7Dx
bZw4nV1L16szKso+5dpAH+M+45H8/STdO/eXBashJUvite4uV4m07qijOyCXhVCA
QeTGEXf4ZwSlQXK2UbBMYGrV2Gt1kupJ0fscn4lqfD00kexI66Wm/v9I+jyG623V
QB8mk0DE6wfvs7sv8dy/DipmWV06rfWgGl1fC4JEUCmQ6AfVdubnv37i7GIo6/yX
YnEp6A0MT/BEmuWm+U0+ou7sE5/Vcw3rDXrgZJ6MPQF0p+CiK5YYRHCENEf0n3Ie
S18vtIL7FwPj2FvaAMFwb49wZ17kcKD1WR0O53Ww0ycBlZ6zgWvjPrupsdbCebTY
pIXaFpjpSz8cQQU9mGb1fPy6NI7Ob+6skZf+znoTOk/tSAgrAdyllvma24cyS/hf
sfUu6ZPhtcnc9YEler9u/7beb/eshtWVntITjkjJTgvhxlDg3IhKTOzno+5RZULf
O1H/fCIBDEX57lDwaUjj2ffs+dq0/hPSsa8gy0rpa8nnovPifm7MEgKyGCvPn61F
NQo/SMDIDCHljBxgtk5ny57+e1h0nsHt1zfZc7qGELHDT81mS6pOYaz9K2cGAZgp
V5laTc4HHxSVC3oceRj4qEhI4yAPNR8zp8xZ42TEwr2PkEz5vybPIm2N+N+oVhFn
nodRNMCydfkTqWsUXYfpaGmz6rqyX0ERiBKBrwZlK37+48vM/ww8l8Q8mtUEy0Wj
YkCnb59qOQrPyXFZM3hiN+hW8ghqg/ozsXywYS0ckqu3B4Z2uhGZ7mi/2hc482L+
VjXSGBGWYDYws9cHRG/gzvpib/X6wjGYeSCmO1nZx9IBGw7ziBdstCeSZS5e5098
q50ToUdJiuaKF57tqWbPv0uYRc0uky8ceYEtzVRIZkOgcA4/+KsLGGE/OsOsolKQ
P7z/KAZaSeV5UkVbKt798vUPLBkG+IJ3NMKQ5h03YTzP5uo4pXfxhqnvqZViI1SZ
K2Gy1TxdBv7UJ5tXS2ch8xtLhcu/sgcae7rjJDQN6OPk6sA2Z3kTHEZ4lupIIoBf
eMWeBXAbcRmmHn+o721VpFogGMksghBkDd89tVFSsB0uRTMsJq5WP8w6W+PeFR9D
YU1uuMuNi5BsqdK9UgjSnbnmzaHsgXWvFxwKkjvzq0NtN1KddXq9BCQPJGJBwu/N
WBF8BKQlHzC+1jwxdfx1dnEtgzJfpGUE6K+ZLg2uHcrQ1BhfADwxANbm47ob483T
WCOfvKaHSI+ETCsYjvyPySsNZcX0QR65DWiYc3mZaq8V1gqNpkil8w4lBRyGJyrL
3wvcjm3JqRhNUBnMPXtIodm2+y+NuxNJs5UR02HzW2qy/ANSuYEEFnphJLYrJzA3
KOde9x1Pb7ReN+oyVtHQlLgua4pGlZqiZIZYeJBV62G5E/Kig5NUto3bRPxUjIT6
OlRz2XJ7h6+z+7hW7M7RNbs5n2fQ6Xn7Dp0X1fmqLXt9s0yjgqn+2tzYMeb0l30/
KnAJOspGKpp4f2eCe1c6H2gEhf+8VWsP2IxNwD0GQfjw3pCxxfupBKKv92R+r1HF
Wr51Jp7wnOv4sexOpxoKj4CkEzm3Ymcyj2xqFOGUU865I4iQbqqDbWMSjmwLMrel
jnqsfCyAyKlud1qk1bnwOgfANcNEYItqjPjvHvJvzogex10sECJZZXRigSaha/w2
RBbOxLb5hAgj9LBoMRP4dEOLcycOZBNibHCPXe6z7pqJW8CIaQkWy/2ZJHo4wrDd
gpqNn30KtEIWCQXcKybaFzPEeyGmSd02d3/IexQyLQdKCw7iicRK9JSvbPPiWu9d
klmJ3nxZZBIWw9xpgBldU9rtD/EI11HekKvNwa0yCnVVLEe1rvYJUbzPVkMYoPe+
JFb/NAxL/ZKU01Ft5ZESXke/LSJIO2e7Q213sVCsNCjfZHbrLPS+r+/imDHYEu8m
Vi6rQS/n6YNJqgaJg7usRNAgpqz9gwMjapBoluBwbHvObu+3awR8YVwXC5uwRmaD
wWznFswais2Evg7/oXtA0l9NhXyf+pxz+EiI+GKnI6VI5++UCp8bYBAnPo9K87PF
dZsgixoEClAQe6VeTlttAKrGYcFB+RqhB9tHdU2HFkE3MS1JUjFCOtXODUBOvnc7
nE7FHx4p+/MCgzAOuq2sFqMrxvNoQ9LFYNYdqJqOQMEPp/zX7p2Dsxm+hLLBnbP7
zEw/K6OsgTAdJ+fc3/XwC+Em5cSibCghmXC84VnJyAn6tvgFiSpqYdYgMYL05fM3
uqR0nYNfmbSEk/5aYYZf3gOT+HrTGhXQ+Yk5sx2NO1UscK5cqWTXtGm+N1Ti5iDC
igDrCkkLLkpWbe8PmLMy+9kwTqZKFW8xraixX4tNDUx0Or3h3HDWInd+f9JrcJo6
jcqYdtGXTgQComFJzZeqh0eGYQKyzTvWpLP5wHSWDNt09ed8ObdHcQfCwo9YeaQU
QiJUHqyvmIxv44Lr2BHBhIXn8VEuwbCFoXclZburrxM04UXTQfL6xqYkHjsgPB+o
0FzmfnjUuiCtCnO92DmkWhUdXkVPWa8pX+/wgSZ32v+kObp+us6LCeQQ4tBV6zZX
03ZgxOIldlru6mbeKn/hJs259GECd0bdOiVNCLBbOfdzjxrZKEdGHp/l2ggMeokx
r3xsE839OjKEbf+ula1jcFFu66MAUYMZCte1GIp0LPfYhdTJPN6Q1fb8Ea5ItvAZ
/gSd8I5brKLnDL+H2wjXw6ybAHYw9XI+pkRHaXvMec/SfpNmJIDFbFOg/TR+Ni88
/eKGA+xRhIFARxf79eLe6ZXdpFTN4mBRlGnTbdIBV/wPJqgxGirYb/GFpBe+29Vh
bkLmak9PNQjRWkiaZuuLh2UFLiLuCoMUgwA6i096VHEU50VqxqsIEef7FuY3ENub
FqBOhc+J8VQhHNybEXCnfHKxRncRXJ34Wd2CQ5w4juGnCqtUElzo4EsSekRIzYcC
ziM5kZ606dny+tMB0T68P97Dt36/U0MWkd9TXm6O8SWTbOFOVUPDQlkmsgLvMhuh
5Kz4FlG1JDhbt6JsDbUKWNjMMdBxaEbAzrHcGOUnxrUAuwT1vJh+wbhUvV6AVxHm
TIU9ltGKfK9GKNq2ZP+xuRd9It/ckdaqzYMOaONtb1+yE9nAa+PocFJKXzWfGQha
fEv6wDzi0nPHYFOofB25GBDHaA6vrc9PwJS1pRFtAXMi49x2Qmc1IXt2WNDooQ6e
ggDv/wmRqWOl3gBGo5rY0sdnPqaiuReP/t8Ty9tU/2ZfvQpoOhI7slWIIuZNbbOc
XzEa2fMVlCxsymiQ2p8jx1zKBClZ2E53EJgxJK7OTZGaL9FHyZ1va1oJUJZkYK5d
Ur4wlx+GEa6mnlDq30IQZ14ktckQqPHENeIslnen5Nag9DbWqbxAxKcduJaeoIl+
X4KeMlVh1d8BaTI8ZQjvBt55/RFw+YW6JdpNhLQlynVlc1jweuylm58Nb/wVAjbk
J7XBdhpzvvkLcvahxadez91zqz0uKQyU3Hv77TI3D5iZo3nk7ZBndiLMQHqCE8bR
pCSD3BEwWz8d7IqPZeJC/5IrTd2IRnfeOHIMHBHWTCASksEevhqO5N0tHDHzcyTR
AEApK4jvSEkCGI+RNCqZT6Aq7C7LDVeQl5E15BqIfKp/lZ9FZoxAT+xWw/xpUsIX
2LpPtjM+ODQUf++hqhiYLa9dlHsGxzgwxpc+cu/5xKfx25K2jj0jN6NbfSjuwXrX
mpg7vsMAZgbdw98DnzaYV45tN/DqQ6HLWBgjckfYqIgp+/iLeSpRkaoweGOe0elh
pCK32Z87VX4mH0ZcSuHiSPIKGqLXC1FUolnarfWz+N5MZvo2KIjxj+1FfB93493Y
2/RknkSSu7GjqNcVhiV8IaRjO7P9ruwCjJ5j91gW0lwfaKUFTxtb9egXJNMWi3yj
tSTqSnh+AM+lkZcPcwsoNDb6okCPi5ETk0YB98t+FLHEIBPS8x2N8cn2m+D5yB27
nfp341Ey7CCTN6PU+ENNUtkWcZ35lbEjkaU2u/aagg5HWZ+aYUIVktha4NaJQOfz
Rp5Yk/uP3Nv8HZJL+lnMs04ARLyd4ZWh0VT5YprDpfy2Mv1T4rJuTPi/D/LPp36r
wWjOQWUuYLr8U34YjKuv2DUR+QO85uL1hvwZOI6Z1jsVxexE9asyG+OEH8VWLvsz
GyAUG7l6ZK0x8cWW+bMqDjBGdiQnfHiHTPM0VLQ4N3G+oQDQqpDQG4HJr5gchi7/
NLIkqebJF9UdAnA1wfq+gXIMwF6L3RdI9xXC5t4F/J7RQ07fAXAddAtDuHjqyv/h
IKzaCT3wcfyll58lXZI//kbWFr/73gsvAJe+phZnIAyDLwwcLb3op9R9STe//+X8
9ikKYL7b9b3SyWpntumKWpKw6MhUN7FN9i7mpKuJsmy/FhGSqLpB7C/4xypr0pm5
OQmvJBOwpD8Nc/01DYQmXgBDAxXyxy0LEIU06j4CFrC5yzO3/NanOaL26J3DzH6m
eQI4VxdZinqFYoslOZZnrtCowliydrhx6LbkKxm2+3HbqHYUqUonzgDQseH+mJ2L
jusq7TNxpdneWUl1fOt5Xsk3v51xFl6AcemGwhWnSlDMRTMnJhyfUD6hQGfmkb/U
2xqZWj2sUs3nyfj/96JqLTEaemq4volIlK+3yUg0ZV90Nuf0K8d1sACnQ444CXpz
0D9QU3Z51uy1xbRSG0YfvyLMXnf2qZ2a9TBANx4jzuFgoaSqf0LSMA6ZAJiHuM8N
NIDgHQYKXNP9qxSpCqoHfrnWcZ28yFyTUKMqvoOiis+8P+oPOmiVadNFn86+1k6P
bC/RpKRceIpKFOa7mCN/Lii4Hj9e8cOf85T5/2uWZ2OcBNJ7g4ktKose9ScP5ndN
yfmGGk4d8gamdC6gDhoLpiEf28RQkCr+uWNBaDMqi0HW3r8F/cgewN+KUXjz4i1y
e3j64B0ujTRCEMnh5Ywky6wBlrp5r/2Y916OC4C+QfnMtfUb4R/aL93keCSk5IAs
2BCWd91ZB/rOrt+bK4uJ/k5BAfwb1+4rO9dgoPT54NP4512pgXlmzDE4RxKMMq4P
H26qr3WvuZ2zWhSJf8oN0Ux0YqgXkAWgO+N+Euv7Wx75G7ppUJjA7IAMpLYSm6Mf
VURVORD0Nj1Tn92pnaSaP98jLXmduk0UBmyWBzQBK2v4EfuZ0apGhRbA8oR++ozq
v8QoUQrdToE9t75CSqv+3HIbG1UrPAG6x9v2E/Bkjp3rB2R6n+34ybWmCWJ13RXl
Bbq/zQGovt1LQzTZS1KYwg0F3jMclX8ROag4oLJgltanOxIRlqiEca5QYK0XzEI/
fJXocWv+n9TVgGO1yqoQQd42RWKindZrE8jRVbBrvoMzzaee+uXp9ORajruWWH9p
U8gkKevzr8s/uqMBdExZDgNENWnS5bghfVo3F2FKT7fU8S5TRrm2rterL7xVW2tY
dGgDCBxWbkdrYQ5NhIpkeg9lHlVmuvGXFo10EOWjuSNMP9rqpARq/+wvRfCWrYNt
FEQQrynAWAtpXOThA9iOorud4TQCguOMc6vKpSgnBhugTa+sIN+bKnosouZ6oOd1
rwmh9NKxGcAUmYenf4ecWToy9o/ea8VRqaiJNQF7v+INYvqlEdyByj25U9kSBKAO
v+o8fUklaGUbMwIPe7XlNaBGkafVlkK46i9qm1RD3fLxPqRrWgvIE/OUMh5jV4bu
JeHm9th3VQFihkcldmimbiaMHuCRgbYlybgORNLDdTLfn+WWj+XOfRPQLvKxqr6p
JDXAbbFaXYz5b6OgbuAOTdvUezGQ6a4Hn/aShcgguY79QcXJjjYhNTjYjgHzr7Kq
iQOlLumAdCz+eCGzXlBz5zk/zE67QJPYXyo19D5YRPMPRUDoaSlp1zcq10VnTVHX
fZL17bFhmtWjHOr6GTOT44rG1mjuwZoeCZPNkvQqJN3/ivYg/6fdKEzM0D30NjsE
c9AemCuOS/TQffPLEUOui/CFQ97L+LBYduKnxeUMjpycPK06HD1R/X+cyP7LdJkW
YnMREDFogKIOtI8GJsoCLZj9kQUtFRqGcRyMF7OM200cAZD2qzGA7H7VwXDABhCe
toVRak2YOVHsbMR1aPs4c4/QQqwAd7NbT417YVcZghVtgA8SGuVYKuXqwJqM5Pi7
h15T8HRzM7rmKIzKZ97Jl0/JbJqzirixaVbYmbK2j/V9hEQumIViTPuFUIIuzWPs
nb23MOMqAkY0J96eC4CjAmu8Lk9pOE0BpCcrVLlTr9p5HmPXSR8ldqhialuJCHa6
XIypORDfmbONNkH5y2yOHegALlK8Zg8icmaqatH93w5sAHs00XYv9OjU4THDAq0y
Y4vYvoQrce0dFlnQaTnbFzIinhYIad5Zi7ryai1UiACk8QMHYgl8DSdWXUuYYL1f
VX3o9Gpd620o5pFHJp6glyoB2+8f18w7bSEZE5rDmnEHyEeEEXNKE02cyEVnjQAj
OLkko4lWyFL+J/z7yMFwfjTO42D1uiPLbcifDmHfuhelxO0Zx1vyz+c86mx2Z7Kr
M7MQoQJlBVciITVa088xiiw6dlPlTC++YIhIhLKi4b4bO3+JSCPOWmN7a602D5ph
0BdGfURfOtizzKAAc8sr9iPyT8Hp4tNckMrQe4T6MvaGymVW4iuHdjjxAQ7aV9lS
B19YegwnJfS1gDdYgtD6K4TP/WBLDFAaWIcEN9THOHZsHClS/4hwbrkezXW3Y4pV
Kj3MGOg1rQ9lC5M5aQ2RufZor5WiCJleSuV1p5D2bbOhr30uKz/M3mVtfr0VZwfi
oSCceytuR0WKoHMWnMieVUGd237QdKYUkPBQINcw3SKYbwmpvskBOmH7GCCxXsP1
esgH1U2Zn2PFcolpcZEd+LKM1TvDmMIUmsXzhy1doA5iNnot/Ya7j5xangqkL8kq
1XaJHA2WZg+j17jDxPLryJ5mlDcoL+Va5Pt4iRM5xZ8RV4Z2XPZJnzrwR2nFyJAd
HVcFAlqR2XYd5iR6nlpi7a+yYlC0jXZsARazSliVFsFPbuyR7jrLdSVwF7UXKkgP
vHUmdUylIqYkcXxWN8QKlRS287ykyg9FVLpRmSV1x5AQxKyDS76Kp4ud1Bup5VxX
gxUwYFBekWA6cSBvLVxHOopa9Y2g0BHq63+PaVn21cdpR+zdqY/4WhHT7X023qG+
/OWcw3ERz1nrMAIuE4clBUWoKFhuEpine6XS8Rs5zPa0WWsJprE9QIiu9ZI2sNMh
Xx1saFNQBkqa+aN1n/zhXme3L2Gpo0uIx7A6uFqtsx7+jUdMQ7VsY88B2tLZ47wv
tX8Asn9Vg6ECgINVJYMjLK5lIzV7xW+PdyYF0p532Iqh+hw/GS2ernQOWtzC8zq5
qLLXdBqyNH8VvbB6qP07Se9FXvFKbdR4dGbtm3jb4BFeu83VjKmWy7iHRkLjsV7F
ThcNy18uD/+HlB62+bMPh5+XT+5bqIkJhxBPhAy8jqohjI4SsFtYm8SuIuLrDguc
1+OrM8yUyu9jxPIJ8h8DNJGS497GDPMap04KFWLkn051kwFzYqB9r8Ve1ICurod7
5DsmfJt244TggLanWIzN9SjdzIsysMu8NyDxMYJGKIGqMzQkkiwMVK1ld4Kf9Y0T
kjKVKLeSfZQmrLipAjwKyiOkMlpE/Rzyztaff960oPI7l7TBRXIL63vcwenpqNms
8U4mPjccA1rEVXeW4wmhQHC8ByiMS4a3dX+1Cdw9WvGzNM1Pw5OFRQI+8htKu2Ze
xV310WxydruZl1WxK1Sd5tyfXh4YWjbYARiepHgRpQk8MxlFGbVJhWHF6UdMPk1M
RGiM0txhwoRoTWF77Pj+BOemvVMQrp2tPKbq+2ZPq6Bu6yYB4fwHE7Zykcbn5E4t
fZ3P3wBZ4Y1EuXrG6/EyqMmcmY2Q31ODdPyEZhL2rwM6MywckzeCKZ78UrJp2vjW
SId+h5L1nwHZdfvRZD0awxOykm+Tt9YgKscGvmhp511ned0R4mqUNq6E6rAQRD2A
a25+DCM7wdvrHly5ZL6GitdOirjLqOOC2vXWC+83Sii9fIxkZh5aDkpeaJpSZlnz
K3EPgz6g8Do2tSVp9EgnerWzo1e9coIH/w/VT0MjQfH56jHrwx3WEXvYungKIJwJ
q340VaWOimp9h+XKVQHNj9EK5lYU3UxzOU1F+SFqQj4BQmQcUFQQj8E127TWYxHT
D/CUCUeXlj4WckQwnoJD4ax/0y5cFwqCob/1tvqlyD6Tc+YpUCQzteM6ZZfgjX0H
5+plidS6BXMKq/FL5XHbKkWqbejGb+dSpIJIjDmg21uEDqPQj2miFyujRpB1sZ/m
WHa2Nyh+an5PQwrMoCea6xpgKE79dubRWKI9WK3G9PpkElH0BKaeQxsiUvVNhB80
W4e+PSoOZiiGKR6GC+WgFS4S3fgMpsAacOMuCk5OIMn8XakPyA/Xar8gjLO48RNg
QR2SHk9wpj1Co6bk0Xsdy4c0L8iK0RS1PePe9HRGS+Zjhq8xQvSKespklnyPa3lb
/GiAobWAHmHYjA0+pFhjTcqdX9qGobZiADU2Ax0WDbfX48buxpRc6bUsRFD8SldK
kJOE9CKL9ctF/p5DpHEVaUSXV9eEOJyGG6v5rxgUbZpGQNDk25RNEVMM6uBFvFwA
2Tz8m2N+rmmJ+sAskKq3ghAud1xglY8wu4+TcAFA8XO3a/f29UbITjxqCtEaosmz
cqHSi0vCQdmJum8Zi6ptydlfZhZCndAWTrqKNgFscxGyNCOw3Y89dM1g0gffmFSk
S5FBOLqQKhTlujzZwUNXE8R6CfUfYtRjJa2DD2Dym4YuHhH7UnI+/+NsUebajPK3
Ozzgn6XX7JkcfoEa90B7E1Q+sev5v4tY2AL6gEzgTjyS9yZyCZhrplFSlWrRSQ8t
VeGwbtF28ZtEG63NFdvgdf4XnsfwAuqyqt24LsNlHZMF4DEZb2ZeY+29QzQ5gqB7
kahf5+9kCj2/Mhe98b35nhWHG4Q8p8JseuGruIkIVdaTHMLxpvWkPBwgTvZwd6wm
1YioVEhSL7V2+JDhDgJOi2LurA2i4ZRrhWNywqIb5Bldiij9VDfSq0HE3Gu9oUhD
RnWAZPiIYBfi6T34Q/TvZl0/PcyF/rJXnYwbTIcJoV1zrr6Jit0n5+kzO8Th7bTz
19pAbb1qVm0LKAYIcIrrGmD1sAJ6jdM1B1YQCTqrJlj5CzN5pftrE/a6gwGbaBbV
MTwdvteVhkTSLLnWr0ja6/yocJyIRhF62RaZn76+DxcHtAA12F/XNnAQuZsg1EDy
2Vi07MYzJMhJ4fdc3nx8l5eWZXnNTfbszrWYV6FwjT59bUA44mo373bu7pNl9TG7
l2jhJt6g0voC4XK6U6TlnQle2DinYF6gxoCQBarIrxDxKFLB6AHZu/8wthFnnsU6
dNUBHysPF68Ikin26gUxK6rrO3yFnLio8Yy+RQxvpk6DikFwTqPmu0jaMnLqRulW
4Rr6NDDiKZwGtD9g0EiwUApP+OOAYvu09dTstyHlSl4uMn9C47nbQkzbrp7J+l2A
qip+OnpPALyAQ0RSQ/54pIaPpw9obItV8EN7nP7JUtCPYWrxNhIffLQw/xrUF4HB
n1KYjbqAkOXIduDLgeKJsSAHiK5KB3OZ31vql50+X73C8aWqki9lsEZEiyfo/WZY
1hRBPgfslk/FYiWe//YC53C8XxE6SN+7uyOtuRXG5yclHJ82Sg2+T5U/POBVABHR
49QPp6m4dGm/m7a7/xH5Y8Lxd5s8gfS8Ajyedb2WXqikBRyLXzZVLShT7gbEoJDh
kU7m7chvZd7A4dD1X72Jt/XAGZCtHoI+m0huBtkX7wEUn6s+qZRBQa+LP1dHJS6O
ohKiqFjuiFvI8LEHAgJF+KUvVYinwXYb9gKcNlRtWi9iQuOzOQKDsatJ/z6clh75
5wkU3wRdsjzHP2CSBkEi3tjH2DQ6hk6JBEP6dZBjwGUrCa2WwePt8HLL/qgs2V6k
gz2I7MOi3uB2LpLb91092K7b2zcYR3P+Em4TL3mcbStEvvZtUQfETvSSBGvNqKnf
ATXqmHsoC1o1/r2xF3YrJ0886vGUUzUJp0LmvygAAQzjTz2JNsHiJIJ97l/zFtQD
+Fh/CmFe8k5EQAGpHPXbnQtb/dIVp+bKdGN4MYhNiv11Ga2xGuHmcwKwhTKBntYq
Ut34J1jv6S8aP2fOZLBOQTWlqGHIfQFhFY1ZGxQyTYEe6U77bGmS9/MYqpjnQvV2
/IeM/NEsM1pzmJM0b0h1wWiu1BdvlSn3pu6tDCBfN//Cvb4Jmx8QzkCZ0ZS3yIQI
kEx3GqewqXdw3Vx4gCKwduw/pOmgi9/qzrlCI6Tng4XMX+/AxipkrN/mZb+qjP4l
9f9PLSNL/L/18IyjmGxuksIfi6+d2QsK8ewEVfz96t4fEwnDp16m/Y9eoYB3iPcj
ArZhXDaD4vmzy/yq6ohjLCA56tB3tU9JqNS6eh0fx4htrwFEv2HeNiZ0Gx4zOO8Y
qjlo2FK8cXnhhwRQ5x4tSPSPVsaUfOD+8oIgF/Ypdh45T8OA2cxyF8zMowmKuAFH
M2zbx5CSoDxMBe3lxqYWR+R+VkgZGewtTp3fE8eJj55BjoS6EdgaKrpftB3XfVY0
/gKfSFVhfdHyinwSWO3CVJw0rtXSRfNSJd0uEw7XKntYrhw+MUEeZXb/1Aq47eyK
W7idwl3J2LAh0vrb4zjaAplLUMx1U/ohPSPVtO3CMzASxN7iC7M6pDY4vmQ6YGoH
r5PWNZNogoarRUlx01Xje9BTBOgG2gnj0Xh9//R/DsTWTTlLicWr6QmOB1WMjE0S
HmnXzyrBALd44/BoYJiuK3jYv5Y9IHmlvvVj7zf0/ipMtGn2MuQDPj0f+cVW6A5G
zuGxIC67cnsYu9vzyHDOK70vCStoHp4YP9BNogivwMexXYxchQgrt2GEU2PhF5mV
gJCVBmRZB6lNY9zzV7SToodmRkhleF7taE9EDhYofsueViS8AsYzW+TRgWDJfQLN
1R13CtP69dMVqMvzc+oBqifC5kQOqCkQBs8lzI9p2uVYVdn0WuJ/sWtz3X+FJ8ko
Hzt4Pe2EXPewVxLcDvm19zNd15S3o5qv/a5SGX4ZbShGvK3McPTZS5mcscEo0SNT
svMsobMrvsqLe/ekL/cLvfIK/qKo8eYiexbr9gYa0osdWvQQiZOqmjWpi5J6lMCd
ccJa+5FWrPZ3JJrcVoRpKheGqhDlibM53XviqG+VtfurQBpv7TdofqmtRsU2xzPu
EFcmJFtdgKB4aP7dJkwyuOAM9QTXOxQNfbDYpYV3XoDd4qQQsFRd2Hm8w9ANlUQJ
LAzgbG7L74ISAA3vYlqV/ZBPht8bQo7eyC4zRpVPn5QQ5sNsUr2rwrPC4GEagwO2
5qM2UhBP2++MJ2FiJBi8LnHSCyVHbhq/lxUFD9rED008M/iQTRuUqt5YodjwiATh
yYSurV7Z0tkNozqiPl970/yPGWihXDmrU8GENL8cnvY2qdKMGWAAKrEMxi/1TMfK
HsIH8ALu/s2vFpBMe/oXK02XMCtzJDKcWbwpONbTOGSJBlyVheeTyjDKi/Bop9W5
6gk3zCO7SAE5N8ZVUH98336viLrDQ6woPEjfUuzrVSexuJY40qCQwZ6PgZa8iGeD
8bggvgtf+D7hADav32epsfiP0cMCEtJRzeiNp62BtTMM0Ha7uS6wTjAYe4b75vlE
0ppe3TpKSe6MoT5HzDqElsFINeULHp4WpAVjfJ0fddtwnOZcGl7vlD9gn5Xg1Ohq
NM5+VpAMdFMeOywfpO8fLAD8Ll/Sc5wTZ9MuAuHj1oOtamZEUUBqVcXu3kglqMRq
M6vvXd0KpJiAdINO13A216zTaImQ9+Bl6y5SX+WhudtyXhlHHBGWsARePuGGCoUx
J1EcZJTMyRVd6vRTM08q4t1ZyKAXFuoydwvwapSHdwgMMUBGc3oVKlzMfvjwnswR
MG0USP98c+Cs2xpeNQkYNyS4dmcVZyTh1ySvFiefESoUCJ03D2Kvy2v4dgiXsw84
u32T5FQVANUbDTdl3/O6afSpC2LvyIzjMsbgIhnOo+CBLcIknEJC1FV+w5QlwkO+
1osyd27K5duscbThtKhHjk/Kcw/zsnEI4pyudHqrRujV1RljkDqy+lHSNi3rA6Xe
P/LIFV78pwGI8DbSa6QIo+PV360g8dMonw52H3HtB4bFmufvRef8McRof1NIDSkm
qHnG8DnMhzSFomJZH4NjVmeE7AsQ/cBKsBinnGdei4VCbqRHgAG17AX3vzYsrwMS
ceYtvc/bzlTHIfZ40Ub6FL2jaAEUL+PiwsmCyTb6APeT6ii+H+UFsByT2/M5VN1Q
VOjGvE1r0X7/cYdoo9N3UrXMstmvqtXnp1/Qg/DnUkOuuoaR77GYC4HQErh+sf0Z
AbCbt9WFAKEHYNzVz4WXxN9QgYdBfcId5obxftDMMtzEhDUstC+94DAh2XNx9QJ0
C2o+0JV6fdaAS2HzCCaLOpgKosXwqDaaR9bs0qwWDNfJUy/H2UdDvMynftixglBj
+1ynW4JwozyL33unuoOlv3zy6/kCEwqO0Fz3rDerur5ja3tprui+AwEoOZQzCuO7
Q+pdLacLWOpw5bUPpv2bJq5QCRBBKJFisiWaA7DxxUGcN30EgMgE87xBNR7ZeMuR
ITSap3sqa8cqXXTb+QVrmI5aUQWUCQfSQBCzDRASyquUN4bWeeKifG2CyUlNiH/m
wtexDIk+6X/8HiXVNoKxiCvTpVaU0MrxqGFLSQ8fWeMmYlmqu6zeGAk9EUGjR3PV
lINJzeht3gVtIAUU7pk7rNxoQucoNpiQaRnWxVjUPsjcLoTtTu/gQfsy0MC3rryc
bFkDS7LLip8bUCpczGzjqbgdS5i2rCq8GgC1ax3blRGCsnMOWx8474AYWXSKbEVp
IGD897L/e6daVcGLNeTbAb7rJef1QnWIpsKUAbTTEHZULvSe1Q6upe12P+08JdIo
IuBZvqCB+Tu+eitAH/BPWC38WOobsCgIa0Ut9NsQ2+9k6MCoXQ7/TcOlym1vxiLQ
nBcF8d0Bahbh2bT6dQT7FtxgLGJcvb/YNW1FUsWtj226s/gZ4hBhs2Z5nqDnBu3R
XJ6co30JhD9Xt5t5XaY45oYP2AYnK2ft+SSn/mfAB+0gvAlYQhwbJTBgBT6AN09R
TAW1lP7vqKMiw5/r86KoD3N5yVMEIRYEbn2hoB+1LRN3bgvmwUijE2d/oiZWbSS5
js0SZE1uzr+1LprBnNunAGffALbUJ5GLLdNECah9hsmaYbpHSuiuFnBHQiWr/mco
t7otBjcfG3AEhgOvF+5aeXUd1Iv6ZopRFvOGOLsdfIYVWtMt3LYRPBTfRs/MX6Cp
8Ul4mLe3I1UZJbYqbgi5O9zA96J1F6uaNwCV3OQaHP2GpRnIJu9wRDmBL2baW05Q
xIuMwvyTzVL4KZ5ffoa93UNqg6DMRimMrtjO676Sq2kEqiJc7H+rvSdNh0Qvp/To
GYIoGmQYZDjbhntmU2rcJLng72iEkAxmnUOiCPYk0NG5QAhzNXCLbwluNIAFWkNm
XdPeUiTplHnUbrZ74kJUF2ECd9jH9CBeoFdsjkgqYDmd2iNmjbc9NGzUvbZyGfTT
2uUGd1oH61dU86HnH0hKf67MRwPv33Fy47aLQ48IVKfvNLBE+TVuSbU1Q9FkzIQw
/K2q2qXYRdBXNdD3ZWAwcVgxbFAH/TAqCy+3tph1mwXVJvzlwrSWWRTpX5ZR/beM
333eOxK1/Cya5+Qys5orlbppQpbh3ghKwhTxxQpnNlB5UAxKyuUHbfaxzF3IvZgG
/T8hHryuBD5iS6IjQLhFmpkLzoVE9a8o39V6MdkYOJkcGv1VlUuzPKbtpXOCXkZg
SSnZ1j/CqFxfsZBy1QqVNNtXLzuUNqHHOcOeRbDIDewMgqcRdkMCZgyElrWLTsL/
RpGcqgm1PCsWyTsneurOQZ7qJMAovMAGNx/dlpKj57LJ1zUCCWQ0izhdvJ0e2yel
jbmaEDfwK/fERU1vAZj9ly94k3/hOxhBR0ZRdvHUqPzEEmQaoC3DyusBCic/7A2q
5D4YDk5uiPG50I3bv65XHJ0CZ3nZvaEP7ctd0XaEc7QKEl2UjuzwZECmIk5viB3q
OyTH/wCJfG0pfMIQYHYEgoBpGn8oObY61h1J8uBAR1MYW5Gp4YIvkuiDiQdegDod
VmG1cBJT7iWewyUftdhgr7xEqhLmI4mhUFSqyrV4T0MJHa0wNpQ7B+eZxvlXMsSQ
NwQXploG4QRFYQVRSt+zSeLjlvCw6f6M++7xKP0S4B0DKB/NeWglgvM6DQIdMg8q
e50cDhGsThJ+u5OCRvr8T9/eQoqNck8+TxZrrQ9WpxtvGdBIgpg9SlboVOJTWgNw
B/tQRTZ7LxKRNYnnYiK7Wl3gEuzPfiGN5g9oZh8kGVE6dvKPIq8G4kiEPoSXiI5G
2fSD3CB4obMQpxwIkaAha9E7r4lZ1l5n3fGTZbjeHxZQGrhY4d9XVPoDXQV017ru
fwBM1kLOgaUipJ5KEjN10iO1NVRN/elmjAEtjXMiX9DIMfyMkqRiQLFCwGKK7rvs
YGoZu9NMWYFIkk5dlOp5dvsQ5EBJ6H7HfG4phhbZrQpEmdgHGJEbxd1SpL9UNMmx
ro/s8OrSPSlZzCfUtCsYgZe+y5dYWYPXY7RQ9feglZv2zktzG5PurlenZK8khYl+
h7KUx8j5FiXQxrRTA+H+HzJKDGSQS6M8szL3N018XuV3ytPz+cNeBHf5Jv7kS4+I
l14z5QwjebOU760mQEzX/yTyUaNOI9ivTe7kbrCK7XguWVzFpNiH/BdFwDMiA7Kb
uIN8n8ymBQxYnig9AEHfuqYAFS8PGHFBPx00CdvOpExFyGYF1sBHuvwe3juVllzd
U+ub94kT41GXTrLJosAhl0svOFPvoAvTHcvM4WKQTYo5P21In5N8cwmQ8O9+rQYW
y0J93IVWIaaP6BkhQJeUc401ef9XANV6l8gWdNVGe1rYE0mKkJz+vq8H0wQAe9X4
GOcxwvHe42E9EDYEfWAIl+oAZvxfEBgooNUKHXwyaAjMrWZ/0gyg0oVnc/2ZZUcP
bF6G4RLY6g4eaaHrpVX65YH9PYY7qAzJCh47uGAKokyshxFMNLiPShm4WJaHSjcl
fnY3dcJ+uMI8jbSkNLBXDyX/Tcn1l5RXfLP6qyFfG8kOAy5h3LNRX9IYPVEeCxbu
JCUkfpDtml4z4m8HkL2Um3awfRX/ftxcmqdFajVGPToHqzTv2NY49xWC8H98jVKv
yl11DwlxK9frLq3Ww/qdiV8ZRtsK/GV9hxVIwGzy8p1sXSRIrtkVFst61DaW8fFK
JzJI297fZs50hPTanJgn4SRAKkDXPn0wOxkwc6V9jwcbZDcleyW1kCXXBeLm0M94
yTnCibWgpqRuqmYHPYjoL/ufcU4wSR2BJhj3FFHezbB3NL+E2PedPoVDVxw1f0WJ
NhFhD4XBWqGOKKc0u3rCOnSKeA/Q9qOekCRkxqUqCBX+dNEffZDnnf+XprrtbS6/
tKnlhg+E/TQsTczVrO1jBWMXDc5AahmLPXLA5Ik4c6UrGQf9kG5tfihWRYCChomg
lo8dTSoHgtyngbTiEXrzqTHSCyXyupUnWcQNEexpzgHOgdfcdQjF5T3iOb7OVIEE
zUUyl95equ+YWNrwSvfuYX5+QSm0ir+KXq1KmPN70ohZH8waYoIWUTFBbWe66yIK
Gvd95M3IC4K0U8OHj5t0Ukfj6BObfyMRvq2QEjQ+CbnlO0rUifa1tO/4vIh8cxt1
G0qP4M/PN/cNi5UeuzkeFEVjpACoHBHtzHIy8OxkaiEwIbgvxqPcKmkFu2gjMD0y
/c80X17pf2hjM48AknkHDI7FaHL8TJKV3j4M37n7U7g3z0yP0aqO2r5ezBnCkne8
VMIJyixXOFQei75+SdCHp59CQnLY1/Xp4tL+37blqXUdr36x28agUTU38XsJk/L7
jEu6HRaOotuwRgiZqp1V51D+K9hByC5AVhHvZGzFnEWRDjej2r8qlDKyCZHeLYs1
SKIlqcq06o8k20s+DWnicvkZfDtQEc79KKnvKDlwO1SdcVtria/RwMyl06ZPuPUB
hRokVgemVkyByJyQr6D0PXNl4YTDAiakLkUrfPtnMapv4bBpmlfKoz4SngLxaLmE
FuGfjeO5eJT3R2ng6wvBNpkimYOopdLUs01ASFr8z2umME4iS6rfiefkh0gx9jU3
e15LcEzBZslZRwXCvaT8o+2H0q63VeEnBiRZjGQ/py0nBNYQgPwHyPRtlcaawCfP
QWH6DKZJ4M9txr2HIyw275BpS3GqduMUlub+1tG3GSt3yPfqJTeXnfymKz4OeG8l
qE8KRqSI6oRNrPIkoG9FwwuKqBGTgyVM8JVlZNL25dHh33aDH7ii7a+5Y0s66ewP
eR6a1ZUAzrN2mbcRJcwiPm4kscJwh/XZhGBxPokWeKO9rOZdVrfhsZL6qQN7RIT3
5VgMZAiaseShbVIlGXi3dfSckCUCn4gDHXjSe76TcBvbCcdVq10Q1jqnCwcjW+QQ
3qP0rwH0U08BrL1IRptF6yReEfENUYVqyEFdjHLuDnLYqWld4iNQSHq0GJQYR5N0
QqrRkeEPhEO+w8X9ZZ4FqBqXFTZLXwEObsQXo1Mn72JW5BgGnnEmaZz4sCSYC/pm
u+65w0QJ9WOAfj68hlBn4jypwZ7NkUKxEh/yGR6q4/PGKNsWgWnQ8IJ7k8bgB2ew
N/5dCMEWfrujt26IxC7E66rsJxUb60wBbHmwJzOqSnynBSCZADqnaQwB/y31etUs
T1MnI+mG5m8WA8FG6G9ODPTMWVPVWIpJNZJg7AozSYqsF/qwpU8vmWZiD0CubKyd
baTkVOcR3JEbttWhczFGAPrlAp6w1d7SNQtb4kZ0vVz26VZ6PlCnLtZw0UOViPFY
fqzCN0xoMB1y6e5P1jdiIH8uADP7xSNk4Y8LFA8cJF8D5S5NfDZL3jeLoT/6KRjU
17tHKBRw7DkMeoLCh+KpeFY+3jhOgv9eCSMpKY1TiGBbfSLpTgkUwV0uQDfY/NHD
6yuQmocL9cSIyRE41P/TDtwWna8Hj+6RuRSU3eF5eZqeIYO6j6jQrapxRWQXZcx5
2c0RIiylibVUN6YYDJeDA82qPKAWObXTV/l99RhVKOsDRZMst1C60gMNCArGGym4
Vuo/qy9lovV6u2hNOvlLQdw5MLsJLPqb+YbFxZBqWImuhFs0F+Rqz2TkQ+JcRXJM
yI2pud8/+Hf3qjNZk0wdswbDH40jFpk1F4SNuY4F3vB+Xgl7Jh2mUyu/6eyJNPb8
B4MzS7+zR5ubv1u/JmpWLVE1FfmQtZl0t5Fs5jNm0Yfo31qWaocQbXrZUutLgfta
p9UVLFauXfpe6Vxoz/zS8Z0F3Zqc+0FL093e1sejtw800AGgr7dPep/p4d5Gs9u2
wh2QgjAeECPNY22VmXkRiqFDOOr6jTe7nqd2P6Wuic7FZUsfIc67CKuEJ9KxxQ5y
9ezPOMnJgMWrqyZ/4XG29o/ytBJ2mZ5Z1UA4OdnsAihkGSC+2N404n3jKgHLu5VK
7DL2LjBTpxo2kZYYTdcRgookmOPLiUrY6zECy9R3mJJ/EwLSAI1NAI2p5da+5bFP
/uCofhjXwYEvd6vKwvp4L+OYLVoAT9hFLXs4fpUbfy5CbvgVAWzyNya7Haf1qH+M
C5EnEaUD4aguGAGNa6g11l8AK7IUcQOsbzM5IcgjPNTU8E9BPYbeJG/aq0k9ll2l
odtbvwMtv/D9QWfoQ18tN4S6D2gKprZjFEQI/J4aXqdgrImO3RNCayszwqz0zOjQ
M5QRapgvsGz4ZUDtXkisxQQA7K/HOIPzh0tx/MR8+011eg3RBfWbTG+2+tixrcCX
J+t0URiCQoUZmAQuVa/Q4Spw070cJXZB1udpdX6QxfEB4ppLoCIeP8q3CgqJbNLt
p5KUw3bA8VVTmsBHM6n0dMrkrLbICqcoth6QY9Y+fZM+1XM62WXekRgIBFijNZb8
o82iAthUmuJqjLx20ELNslcPCt+iY/9/pVIu4FhZgzpzWphgOrrnaU24hjrePkmW
sGMrXczdJriE16rm77u6ScVxZMwj0z/XiU34/m9wAF4odY24s0SsUuH3d3iU0mUb
NMbm/jJxegXQuCTUUChPOX+yNTZjtRYW3lFH1YZC5p1eeKg4hysnJsoUv4m+N3Eg
NBTh8szqn5ntiFaLswWbWCIjIy4NYIgJwwqY6itjCnemBGfsxY6N0L61WkmqMi5/
LFCG4HuNetjUw4TIzFNZ/dvX3PI1N55mVMrW27erNe9hquCq6cKsnbkw/gwhpnKt
oCifxEsWf+dBl8kVfRLrlRkwe/pIXU5pqY9HYi5Z/9ugVdKPppcQMvFgI/xPfMov
l5diuUHNTHz2YLPonC27iXQGqI9dkok3PLyRrztKrQrFxfENnwKGi3QLyW6aKGUL
kPt9hkED/aKX0JFm4kJwTgE/8qt/SosdYGMEsEZqZ+TIQZaOVAjOJ81XF8MO2xST
rEMq/zho5Bf8eJZMdRI10bJ0/xYxI8RwffO4HtmUuKqs/b6fcD+OACPzqHP6niKb
6HpN77WgHpFDi39eiKVBmvDaccl8YaSfz25/08ouxV8q+ebujk4wp8vxCtnuQMQm
Tz3rLYYjaMOaRXsuVWTgxVg2cu/p3+dq6XLxnmFY4BLdUUM2NK8jaxeRxreHXejg
xylM6LdDi3jJTOSjbirpFWe7/x4otZRmiFPNLSLqbYDtaA4Q/3ejza/6O/rSNlOQ
Pz5GRJwZpOsccGMOYmF7RHBVPOVJX/BeqHhi5zs2QR06XYb89uwBdYXljm2OK8Bd
uHHtd4hnXGwCLHAmJnVtBqUjxs+aMwb52iYxstRTe9aTe97ub7V2JU1AMmMv3OE8
mo82uPfcoCb6ltu1LUyDfLhYiptzJ8337/84pr+uZdFN/S5BXDnwkNkTWUEDY4m7
yHAalWbXDqgRSFFhnevXEnQa6riipYKHTf6ZvkdU/O6BVlNdnzonki4mWqPleNXm
VNxd2b+xPOqLgN0gOs+Cub9qs7sB2Ad/ZI15FKVmwESLUITnLFvmHG58PTEP5VHk
AjVfczcPYVKuWW7hVbtKY67P7lpCcSG5IkoIkMezjPp1L2CNLlklxR40BUyjeMoj
wFIj4NxGvbOV23Xz4r5skFPf6N1Jnm8QhwzpcmYczNASBidDbUsP3AZIydAIBqbZ
idSN1LbbkqgWAUm2JPOEOrmZr0sYp6qdJMXdPL9RNWBODPUsxqfPPJ29AeEtNZGv
Ktk6SnTNoSHAEZpsnv5OBgCaHqImiiO4VGqKCn4RXYEDIN8QxiGspGt8J1T9jRt/
viHusd3UCWUKE1DiKUfKLgijBqPY/Ezw6vxEAfVrPIOO4n7As8u26Q07RiPumzFV
DpL9KmPmx/p1XgyOc6pqkP0Km+Fhg1YinSAPmsQbGLhapniJXdg9x8a9kY6+PI5c
/oeB1jFPp6GD/U2SdCCz1Jk6d6B6PAWAsXwDTYvlpy1O51KN9d30trmd0iA23L4D
WOLUPZNoPNz4FREc4azDz2POR2/6VVxe/Eyml0llD+Ua4sqxlE29q4Yv0NZyjC3X
pFiNvZfUyRKWHl+URIRKJKjfddjd52pcXTWuoJyT4dRxa6DIfdRYdJRtj8gWrxkj
/P8G83PSQCsD1jChkT0nLhdEXOO+aGTQmErvhB3cER6jaQdqClvNYZ/g7pGXy2kx
D7gSOVnv3t9GDtLsusPLgnLouJdgN0LSjX+6713vz6iXJlmIFIx2r/Z3pOeLpraD
zirGITuk5EQ4iLtVGF/tc1rdYeorBO9G+Xh4Qf7Ozqn7BACT4afMikJFegS1/hwJ
UnK7k/1J/nh9LH8v6VxXXglkSKK7xyb+lIIMAw4ZWhouMF1dXLI4DoFSX8TeqI2E
kZWSyPyvUTcNM9t8ksSo4WpmMEZRgYIcMBpRNVq4lPa12X3xuiVTBIaovUUS5Pvw
GBnysdk3cV3M10EXj849CRTxtgKgE1YgpnEFrVQxuWkRR2bZiNee7Qilbrixozly
XWNmEInexESifEKu8fLcFtIyTI6gTbegLXwamCXrcrmOdaKRf1a6YGWcHmSgSfxv
sz6SIYtgu9OSn6Z5rogWdASsKDNRFxOF4vfxeRDrSrFMqg3Ebxv3Cb7xHsKEtkr7
1WuiwTWWRG9UDzp/oqZZ7zr6rjuQhgK/xUGb3x8yopQYhhREoTSM/QK8deokBxtN
lB+J+tgzy35SH+uhi0LZwiCIFnuxwBRP6oC8JVhyYS7Jo3l2KhJl5TwmOy53jy5U
hwJTzWz5ucuTZN1+kuNddrNUlZuXpeABXnc+mr9wLy9uivqxGCs/TRerWk1Wnf+V
RbF7qGlmoFwi7Qy8znJYTVa+KrVZ9mS2leE0Ji7HttmdgXcbdA2lPWLDxmOPotei
YQcdiFMS4P2uLKbvJsBx922QbKxD/mBsIiTL86g0JHfYqfkvQ31c4wHbma9GJGVw
n2c65ExLgCYsB+p0YKTHhvwKhCEBVyEjQQD0zFKtS0HL0h1c9aRy/5a1l8v0XX0T
oLfWerN0oxH+WOWaBHBTzcb7Atd+hJNQ9+ra6STnuLv5PY/mBeWhAMvdBEZRufLT
CScTj6Eif16F9GZS0+eoGhN2yyPGMQyKS1rnzLJfhR3eB6iDBVEu0X/ql2ySDRi3
9B8uH63rjt4hUmNXszOgWRzxWy7wK2xr8EdOpYKKtRU6YFM3pyVwy4g3w0hSUs9u
YB9qdktTTkflnb2oqTDDmIMog0au6F1my/WsbPuTfDLpH50+B4bowekEnPG5taYr
zHfx5HlbVJTrO0QpQLLg1Xk9fjvHhXw7KCY2SiElvWvjNRqNyvqki5Vl/KMzGsJo
+fzV10k7oT+Ctf+mToFp1O/LnMliEiyv2/FOGVUDZmmYpgdcuBMuwAwhwB6+Ky6a
p6ammLGyL35r5wciZS9peDxcqiJ43iNDbBe3XVvpyhr0QsIz/hdFzp0kfPpBWBZu
gygUjjhr44jgGnU1hM1bNu0DkBaFPEXoCYY6ewr/0O81DBQIugZZHAubp1TwTj8a
5lW4m4r81MZbjRTdGaq1DG5w4riwc7MWwQVpbK370Li7tLOC2y/dB7zosOeaSaow
f5s5GCVzvbQ/+mZkh0jgOSHljOd8G8tEvosj8q/2XxJdNAaQf8D4yHccMjEiJF9u
tldSX8ja9jr+mpnFmBE6qF+j5E9ssNTi7aQf486fnvMCBq/1vL4NdS99FDJPBd3D
Tast8W+TxyWWnGSRkKMeXJC50mXNAHfAJT3+JOERJN0rZ548ZrtEx4l2rn18TeW3
Ib8JU0JAtiRSFNISTMdyKo/eYtf4jFstWQLyzfs6IuDP6aMwq+f7mwq8r4H31CPl
5Sy+LbD4JbmrmqE04o0XuNMkfLSeKR5+x8+nVcQVtXPiEs3vRPMwFhp6eNPQTSlx
Uw5C0c3ELAakQPY+M5C6bD9KDtLHYPEnAWeAUDYvmB68iQxtE72xAiWHyisLEa8G
sX/WqAbYucDFt+N5Ucj9fo947XIDRMzhRAfJnr1sSkp250Ax2TeTKGPKEvxNjbxt
+frHpAzMJQYOj8mhtuXE5xiGY0Bo3OBmh0XCgnTPKdX55K7hcWCcRIK/kfM4yky+
YxeWf6KsaP9nqmUv+RlBxv+sdJK9gQ4fGtmjusiuP04kpuHH7WLFmzweykbdf2pF
HoSWllYevbHD2a5IN1MyXbuSJuQBuZTuwdMQj0IHP5LestKdX71MNofHCAomekJy
iA4kehfxeJQeT9ky2sb7JGLKdYYFUorsbLGsgmILWkIOIAglQie96iu/h4CJXQIk
H+sk/VijiAO3iro5eLsEBpYold7KrKunv4hoLUSqoNiLpeMfDBLpiLmudVGJX3sl
K/rMfkQ1Hxmxje4g5G+GqAmH+dHzYYo7vBU6PEPhHUirsJwuGARbz9IMivQTwGkL
DmdZg7O7SJTBAwNHDqV441kESImkFRcJMdxWbrk2ni3Bd/fUYftMCPVWKtWqOqZg
65XFNsuTnrZ0FT3VMUj/z1ifWhkuKmsqCFGN3BW9E7vSVUnbCM5wR9VYr9OBdl9B
VaoRteBavQf4PBc8nyDfVamBuim0ee6T/4sw84Pk8iyElY8Om/KGZyeeQOPVG0tZ
YY2897e+dEPQr2CV5AlUz/ECiHXJiBRd2gQIzqvebUWlJ9T28liGJYgJTOzpfMCJ
9K+F70Gj6g1mf3mlS1b9bXvKInrB0ct13c2iew2TfF6eH4Xk6gU3ESIacniDweVf
AYRVls3Ug/u31K2xtC3lgRYIbAHXpDlF3mxVoDK9MOlOxaOj2RF7SQO9UkgyHH0g
zPmMUCJ9uP1YgrpT+hzFWAimVydlkRPd1C83ErCAMOw1ByViA3VI5/sE919fM2H1
+3Lc7CQsCx+BSSzS0Y7QJJRLpQ4Ukk6CXig0q2cY0e+lyo1vz0PEsQEU4kzTHLU3
VxRJCju+j5SksuuSFCQpCGekD45dh5GODFFDxPbHIra5T6Hs6bZIUoDXWoqipCIo
fVlaZ8aiEsmnWYoTJlP8Zx0u+qpAFNyuB96xmAFTQim/+OF/eOFJW6nzg/BDq7Et
wWUCL+K3uRKtgkcC4feX+Coz9PP3pMAHutBkiY8KrStDoyiW0tMIO+6WhwclGGgd
AbW7aLB8e2L9B6Kg81UqrXIVT3Z+VrlPVcG5wwb25jagQ1KfegBGB2c2Y+wIDb3r
ECSBozW3AviRydPOvDms7UOO/slXJIHTzPvsklibMG5qth0maaCBO7yU5dX8PJ9Z
SlaL2mjL6m7YFXMYh6Q5qMjgLHW53teE7Ub+emUcMauXJxlnPimWeSPRQ4RTXSgI
qWcw017R+2oeRC6OXcEMsQh9FyKKjoQFBDu/qxFcO04xWNOY/339e2Kb4zjkLu4W
vX9AkTWLlSspakPRgaMdHr3CAmSioxiRXXZL6QGxPztAEyyfFasydWULbopp4Kq9
2XADkPUt9QhlHbhdU/UNufSxhEYhYDF40G7+7NnRX2Th1xtw1U+w/esx1+eCeI4v
1BJlytLdJFOxAixt9xqLvhD1m3dD7KMRcF+4E1bbrmdJZ1ArLtBCjIv+dabKKALK
2NHcb4AloZyKktZFljDM4NDWP8acomo3LlDmUQTgygDjcC8fzkfSnmrD8vb7KuhU
ixl1hGLIDditvrr2D39ZhqacnL1klfKBM2BWwfhFdZxb2U+jrPBq2W7MjXvGc0+5
XfW648Ul/iK1zNmgRAQ6EPpd37K3Z49V0vl6EM9NLgkOBqd1X6+GhMKj6gIF9T57
PTlXeNFoQc+pBav1mhwPgxfj1Su2lICf+2tywNZWT98vc69Le0NAvmwO/TnL86Wr
8aJHIRCkuisJFEsJbEfHgKvAEC11GEsvDq5D3TxySJ+uVg7hn9ZnULgnBBdiL9gw
wL2CqlCST7+a3V8NEsqcdktYgRZ9VAZXhE5DQQcuc1VxQQNGRdbXbEuEO1+XLxMX
P84rE4uL4cGcV0lcDWdZZT22CJ7h6aimwUXWKC84X9SrfY5ZFhOxRpLn6rFDfN3K
X5OlFn4jWcpGaEe1kEn6QBSfxbdn4T0RoWa6mr/jPhfN2XrkIi6X1gOdB427lbQ8
Ahc++WQeWWACWt4sTqWaJCFjtO6YeYpg+ywzPw52A2mlXYJ7UiLSYJNLNuo9xztt
tnvUFkYiJnUSW5AIL/+APw87/qfUkU8AIWdnq+y3QEg/4llsHa28xpwC5j80vfC8
sTV4JtK8YjQsiHZ5XE3j3JsCXD45iTinTxxHliLhDXgo1afPjS16olVYaKu0hisO
hZvhr+W7oTROjuF13C8ZyiEvJxZ2IFV02l8C8J0iIfR01cugZtp8H3PjGRgdpGRp
srfLAXSYpZWIVDEdYWC5ms764P45KH1eyFsORkO1rEV38xTNEjeVyFTySUJO5UKd
pRCS9imoyZ6K/V89nBvn0p0ujS/0WfOVuczNRJJQLZNCMTvxzVoofVh4qM3kuR6Z
pnSHspwewJzEWhs7igsvJ/P8+qXxua/7yaQ6Yj4B5Akk8QXleFv8Kr74LDEKHs0O
L4pd2yVa85I7v/QUzsc57WXSYnMmivGczFqcGDJvNDnOp6ug8kWnLytJonjZ9Og8
EnH+nancg/PAYuyZKh4x1dIYUd698cLBsMLbw+Q564kEh3Db0KP6TCrjC+1ri/76
telJazqeyAf2ukroK/W4X3Nj0J81lOoMRITNSanXVCeUFw4ifW290QYDgKL7fWxu
zcKAuWtO4b8wdGffLfPI/xdArCFO7kpiOaZf7vqmUQeAhE0DJvvx/IyoqLC7K8C0
y1Accvag/jscFytDnMk5Sumn0KjP+RNBowj/YIwrd/n7uLZwOZJblz1uDSb/Q3me
dqpVrY2M1MfvvAzYicQXwTENR++8U1XZkcTS00AM5B0xanLYEnF5ZIKY/iNVAGE0
cgcfBs0yqe2KZrXfDp7Qey6RWc7jXk4r+dUW6z/0iHCigzqd5AEtUwlZ48NMgprK
14q4RpDwk2+eUNilRTTh7vWfVEMV1tLn8phhQON8HdCwKhZkcwuoXzxknx418rb/
NItQhG27tpet6aevxrivVjqIyVtJlkzqn3Hcjsw//3YYq+WhrObCYg3DP376kTux
NpejpczjcC1CcoFnLp09lInNoFUJJZgaQOxkkzsQQwxKTy/R95RFqvKJhG9ReN1G
2SUImuFgrUwnWAI0a7KW7cf9CN2zzEnhPjxDTbJZx9kC9HA429pm6pT33xHt69R6
mtcHF38ajiRUpBJko3KTQR0aXU+AXIeW/Oi6n5nlkpzVl6cQEEOMF6AWYBOoQJiw
yf2eFN5mLr/Sk3mZ1vWJKyfvq5eiO2tRQQE9INsguEDkIy47jviLSrR6aJSD8TmW
MpKdqoLMR/962wVOJYTxaLVva/NyBHMcX65Zy0EGHmnbfr2sci8SB6bcoyJ2Q9Sb
jSCRjCMiPXVewWB69l5B2A1h21PCbc0yAdauwb5T6qwdFTXcn0nKIHKert3Fv60I
CRFtBE8SCD4yXreGwLwGoaru4elmqAL6gKJbFCtNezQhbtH2AYvQiovp+cAT69dr
EDOLAf6tbW7YIMMFc2Y99VC+d0m46LLa/3ljDF+uuITfq+auLFDDBkSUw3tToOO+
z0d0JsMFzcHa1izl1BKdQD3yc+VICLCbCNfdN7RZDRUY0xV1NkzSJ9YX3k5tejXW
Wz+e246cJUfz8/BZiRfziHj8ome74A9NoRG/pJnA3TCYI385f4+nS7FUpnr0XAeI
5PO+56q7jzZfM0ABAquO5XFXbSy0w/K8bMy4d4XTTIRuM3ODpP/LRuKN3kTreF5D
BGihWyiv9A1kDJrpEiQeI7jgFjVrmdeOnBb5IXiBxSd2VZw7MdfxLW62pEQ9wMhT
TF/9ZPTo/y6cpMkpt9YUp8hbhFJOwHKpfTQ3zRe/QborbtE83lvifIvsMuKqBs8W
gJhNqYTW1fzkHz3//jvm5tckvNRovqnIWdWkSmkowPlV81fZVEnkBq2UiQ14FB3m
1DAI1goQrmH5ZahRwoUN2yitirqk+oXqaYmpeLHfojfzx6NXuGNTsdphLbR7y4w4
HzuzEvuQZjC0j6AJWW6nGm3CmfD+GNjB8emHFV6IhQ7sce/lMmImHsP8mU6UNxg1
njlXBvFompbAnEU40a23851/veWkh4REu0uRpi1Oc+cjW4ZmlekjRVUEIaV+z2z/
1+jS1YZEjdrNE8m6mWmj2YHrssNmXZXSOY4by1NXF9bM7/ETc/iSwOTr6jbwIzoj
InpexVx3VOVPCqvAZBFe+Dlzn+Ujc3yGLi+XRxwuLXW/hbRDBA+QId8F5QUfSMop
Q5REuvFeTy7ebbJmZ9jC5rqnhZOmiKuwBmmSexA57gpHXAAHtCwFvcTCUWVAT9D2
L8p9RCzRQUMekcyQe9hGpjU74kaWO0Z33RShARwaxtgxBCQHh5QH1IMRSQhahJa0
RoXqOIq8Nyrtwwn/89hSaammJYtpTO6KcGMimFx8qgT/zPfrFZggGHBnLQF28slE
eUTkEWi4p8BoY6wW8kXveS9Tp8Io9bQS7RLVzG+NXNlI3iS9iLC8KMjbM/7OWhof
9EHN926lYdHRV+mA1PyJ1N+RRSpM29ub1NpC+hl0ddYpap/b4IxesCZAsYlDWGeG
yDak95DQbfpUucr9t5BSELB0IbgT5Ffd7G+S5TgoeTnEKpPDJIfPA9LLSIyx3IXE
8Sjhu+P+MnaVmui7+irUyoADt/FaNnw2Cyxc0/K8qdG/xQJN91nhe2fSQgPoFHrn
R39Kpf8vVYoMLfSVTvly/Fr4Suxci+PUbRxHKuAd0ixWpUUFGD5LIE1lRHQ4iaqw
B+9TOcXzt2Rc/DqwEF/+qWxIlrkiPlVu9bCC+QTFibNunxJpbbpgx+wr87xJGx7D
/XvG+buc+xgtVMlIkA64EP5eTNd6EV5i+W53SmA3g0x50XdBn/o6RHvcm0vy7gIT
c+ToMDoK0hRxZJwgg2FjCK28iKxQgvSazPfpHIyLX9IGeADFRpSWZf5gdRBQsKWM
qcc4ybhvcYh9lge0nUVzfvgXYdKl5iDdPlb+htFSZSjOpGYrBL+hNRPpAKZWs9GR
Z9EAYzqauQPRCPIkogTOXb6/yyKOXUVlXb8tjtwo1QufwAPQS6rpcv2Muav72bB3
6OIjdxqAg6OhjcCjdbv58tIgzuUchlebxwT+wruHKlaYBjlKxANtkDDoKkEy+vvg
i7xKSPXQswd5EC4vCidtVPdcd5H2sDB2mXIBeGrOcQcLlyX6TBQBq0OokaB/8wrt
onyYeiQVvAKBpST8+Fe2UCofZFIb84r4vc4Tvhm0oDG9PBIZu6yAc8Nn4pmUGYAV
5OoEnC/9q7H+2xVN5d3gKgYwmFNETt1Jt0TG58rvn/CK4eJH38+HqmXC5N1ekn82
wALSJkjfhbLPIBE8rq/CUE5C3tQMsju/6t/OA8SbmOhZHyKZ0KEV6ceKy8fj/I2F
loMKnbRAfXHzdopDTSz6Jvy89oelUUltB/4vx7nq4/9bdlN0okuJG5dpEFPWJ967
C796LpWhAvA45PamEj00TdEM7gVfnOncbAmnMzISN0AEw4KAv2PVzPdRmfu2gz/d
p32DIL20lXWAZgHPnXxYvgObBJvdJybxxnt6mA3WCm5+H2wZlxaQX2ZzSzZCPgT9
X+vY5ugeaQQ9T5MbpeOLBp3eNoADkjmb0tJ8SshRDhhexl124KO0Xs3fXPxekNhA
eSPQtRUKbwlSjajn42cLxNpWhxuSKOSEuFQRIRJAqnAW/gMa45Bre9A+KM3rH/kH
n90AHOJsFXIHjzCq3aoGiArsb4xehQ6Ba0HAtM5WrAM+EfG+Vj0bmJhE8iUddjmZ
viMk9GGa39pmQEHSeirdKPdRCoFVZwO0/yN0F0zspCQhSnlz4GiG7S8Ht98bfQzj
yIBm8fPrZAHstwSvrYpPZbYDKVdJ2QXS3f89/wjTaUxQR8drVxSGxtIEoEKbaWTL
A6lQTObrnJt/mvK/BpRfseBNLQwF+zcv3ruVWsxR+Ap+OGqBZig0sbd7NbX26pSm
i8DEzeiTYeoSlhwvo21ga8dQ4Q5ywgWf1tRyg9sXGVpF3MvR+Mw+WlNtCMbhozXd
I0COfm3QzpxCj8JqsWVbkEb6tkvNyvRFv3o9Qv8F8hCW1abQ6RSzu9HdfE3boUL0
gcgAWEzd1JKKMbv26zspFVXsBdc5T+jrSf1Fnkvlni4eXXtJAbnVrUq8+256Ckib
HxcQFPnLABtrclQy0jZMKS9aQUuNER+igSeyuN/Xp5QccoFhlJZUVn2z+MMdBGI+
iQzprQfHcligOQogMWCnAMlm0+hczg6NBe4XVIy9k68JxXkpbYH7j0SjUWeH1kXq
kq6SBNov9pkCxkuxmPWoouVaS9LxnNG3eNQzFQ2wAO4gEyZSQ9BL2fTCzmbgN0oX
D9jnNvNbMB8PEBCRBZ/ja6hZ1tgIE1RAYE6VBOsONDO3Wc4bT1iQXo6Wb58G0q7x
AptBKo5l8ocrT9uSpCteQJS3k7DCm8uQQFG4mD8dMkzlKDgYUgFAAT+leXZOfYkL
wfDd7FvGT6HBCAR6IlUUIRjdgqinvsuW0rQEDKy/HpyUcmIJ21vc90ceQV9qQFee
GLx51PC5OfcM7E9PcDgr4JNJJUByDkjLzHPbL00cNOvCVgEFqHfWNJfQP5bHV7t2
USAa0UyAocx0fjdP4MYyOc90JzWtySoiXLSPV/kpvLfODub9WRr6DF4YXAQQ+8DC
0KXNyXxThuu3obqipe+6KVktFZuxRndnVghaC+7IpIFcqQAB57QZ6G6RaMyHMiGv
akFt3tbtJk9Mte1UPZbBUie2+vt+LmAUm6/rMPxbRGFsgzFZMsGfzYOWFQZqfhgp
N/fQ3qgHhoiqWyQY2aL67bZopUw9EDtFna/aRuIkxk0sQfkrfI9Tyz+ZIWJiZrdW
qvB2Pv6gzzJU+o0co3zbWDtjqgQdd+VE+8lEr2wroQ5OERKddkAhvLT6d18jLOiS
PALdv7OsARqWydOlBZSZP/TwKDhAaVMcfQynritaxoiPw8CJmlUtHv1FqkJfOEcS
N3Vm6QgV7ob/HRsLLNzBMBA+DD32WPjryC5CiiQaaOh6YXsUtHLsEua9MLd+XeCD
cbgRvBwA1j9zU4TovyLb6zxqyyrsfGIvlvRQUeshHXD3U2/nnoSRbDZND1ZPHXU3
y9uzDQuAKU81A0WeMZTQQ3Da3tryGKzoWmQC7ChrkVir5rc1VvFCkrI0qny2Os6L
2F1/j3CAZChzSuL7opjFWVx3M6lj21oufeo232pFrGHmnv6CifUShxLa4uxdPfSK
xT/gI0ZftIXcXCZmuGdOaO0GVKBlvWqChvcJIz8Zm5P7Q/hekprbLeBf/f+l5J3l
RPDawZlpEpBmjSfahUdWPirt11hUKy1bTwKglpaJB2J+rBgLd3dEAB7Zyi4uGq8p
Mxld3ThSwuuHCmBqt/oBbw0nlMOuClQ0eDSnWwu9HBAbJJNeHSvhjtefh91rbzV7
3sgX61L+UnrDrWeaVQaK0fHor+/lTNYuT7hBgijcCoxfIYD4NCs26T6IHZweZLZX
//jebbFFd4vjz1xT5njPLkvL/9VsDUl+n1Knkvi68I5BYxJfHfOB3HkOlnkjCqol
W1FbIGZNV0rMdo2vOCmdT9On5VyqunXYyg5300ADx1JDMbBgwvbeTCFhae+VaQfe
UMWq/H1Qc8ZXfHjN1I2OJAF005lq7OYu10ii62IohEhu0mEAGjtFce0K6EIl4WUR
tkuQFkODLHnxsaC2xSQCwKF4uUKy5XCit2QtNgWsjS0X/FJPksVru4PUQYK9ypDC
yaLA+pBXxXAMx2yrxF66ZVz9bloBTCddrCIx6QDZoNyNpAZlrB/ti1D0RRntHd5Y
XDK2szvzLWf4D5IqpiJ8fMrq5Fsb2ynCNeifWp1GgHKxHyd0x/YFpRk/hFqNiWtz
ozyOgLPGDABm7PedkG2hN0uq42A4zzrI2i80AQ1KZzTCZjMkWbNnwo9HTDc+u2Y2
dI2wxSXyul/WBR1en97n1ua5/YKHGkgO/0AjKoA63ZOFgfDjpcI9RdcF9qUeqATP
TvwhX6qzKd58Q2BtF+i9kzsd1LFGc8dkgGidmVqCcchHoE9I+M4rCQ/YRIfpuRLt
uVxeljr3zCHzVhOabZ4brr+0tp515SIEszQA+nc8FooJ8hAI/m759TF7XwVMO0oP
ncRDFRgWEBEHpKZYQmOqKmG9AxLJLRNVGLmvI1SmnIRjhZdbnkQMdGf1qVYEmKmB
3i5ZNrGigVQ4NAA+V33AVe/nmATvRVHWrsYs4LXCD6um5tQdz0qbGB0ND7z6BFcV
bBq6SmWaYmn0+VEXw5BHNE8Ino+WjfmFPlzYl7WrNbrMV0ONXZ0TTCS/v2YJC8vu
NpINC6tXW5Z8Ypu1JwOD/tWQCorRLBQT+A2ndiZJEIV6DZnF7atntgnkHBwRwAuN
am5qah6nsg0RFky6yXXM0tdGrJ3BNzPZPe1OFvpNj2Akt3t42mv5BY2fClZm2F7D
eVBHXDIPVayMxQWal8j6jD4VJQLkEEb0j1Y2jBDFfr7yFpRpjtF0/sD9V8Mp0Qae
SY/mM8oKk/vR69UFJu2L92Y2ANiDcCe33J9klL87INMFqpRiwlNTPSOqPDdzhC5Y
61kDBviwpcwUBNr+TU9ieECzt8pLG/GMTJoLikOjLin2qIeSmwuGFM9Oyqy8hbF0
KcMtKdhTCMSyyJrdElfb1a90Ww21Cj6VY17svtuY7aPPyMowAFFat5pnRiRxChhj
8gNC21XsvI3uEE4tW4D/7F+xCrNjWyxlmHfTWivmX/1lCGE1LMSTPO2Ug/9IYZRP
P46fbY78BzeSMz+EVkyUWj4Ft6LDRoIJ6cIRMCOvPMdcYcTj6NjkO5NqXAJVn28j
4w2KTqJ6IGhzK2PT6HXIDBxszalGKsCo+AW+8SA2Ce6KQVBJRMGqWaFAeTAlWWUI
v6AQFZ7Bpjfpup64kVSmikYHM1uGhwmIY44jXB7k8Z+PPjUwFCml0zLJMHnjxC1V
txFxlPpOdfF8oXjQWCCqgzTdjbyC9JAZ6xQUzBt7NngC6K0dxyu/fPpb4CAGDNaV
OqxrZnMdRwD0hFMFwaT6At05eS69o0w5ynVSX/8sRvQe+jK05NdmCM6FX7j3zzDG
i5olJ3by4b7iEz9IPKjyD8Q9eyIBHjjPlUWCZn8CNz8rmI5Sq3qwSvmj50s5VDvq
PpLSiSHMgkRNEvRdN4WhzPmz67T3hoUQZA18zDneM9/K4uZVsUoHP6gri1MPY3Ld
CFX2Sk3m7wYtZ+qAPP8kJPm4adFK4yPswgHmWRjn8r+cET3MvkfNdPz8VxcEEhRc
4QGtEYHr/aZYKpRh5bfr05a6ZxPxNQ77j/omokj5Xn01kmzgbwBzNwVC7wX5IpuO
CRQlMX0Og1jXeZD0k7VNi1xIli8PxXiQNTMeatMcboxtDSxMDyyw619CEYm093jM
M+R6wRchFI3ukJVRKed6C42i/3eI1Tf2ozwbGXuOA09RQ2LaX6MjvSDu9fn/zdWe
X3kdZHPy9T7iXJu4d+6AzZtm+4xDVK0JW1jjZ90aIB8wxyfKUro7qwW0ZcSEwlue
UgmDDZMcYf+H01opduIgjw+sJ+JoYQ8/L7xXbU6DvUEOMcn1hx9hLdafnvtKXCZM
K6IGxmNMrL6BIfU+P9FwJAesFNgANFMdUaP3/80EEKQQPizeIXzyMk/lg2fCblh1
ZDRfaYmqQz9xlEWVsjEOiM/K24mtZRYD2OO1ST5YPYTxeYg/AnRPJlojk7FcEHoj
/jAxtbzItt4vc8Zn/Gzfkl5R35pRcLOZrs0QPv32hEW9fx+mQxWJvKOSoYnXlxK1
+AGkeVJGr5x5Z7x8+KXn6QXDm5SEXOoMbktNmePX59aGIPZbirOf3TxsY3yCiReb
9e9mbT4fiP26bfdRG9jHFeozGUUcj/uQIaq9mDGiks2rqbTDZVL2Ljveq6N+Ge6A
KHvWEbMjY9SDFhdsVlNME/DeCRUP+7u+Xx5tJWtQlF9MG8knH3ijheUU+cGX4HeT
iEHfD9l3GoeeXWNV0i3Co0m7X/j9Bp3uoIP6bfZhP5rpQRUzHVmLx/3toCihRvm/
Chapv9WjMkS05tJ15Oqc4NaKydAp+kpUXq5xAEYKIHzgZrK1q7cZnHdsnI/kiWm4
14RK7osKTkKWh6JiYaVcSDMhnytHJlp7h7fTFzWFkobh2LjGon1u1jUKGK2zpY7v
PaCl7UzFSLOFU7711LDq1QZCfwsKvhZqCVM7Jupfn9tQNBXSINcgwlJ8WpKHHN6y
XRlvccorfqB6BNtriA7wRr/YAzfDAzZ+C2hVnME07S4FD7HNuep2F3jcvIWCRUpa
7XIUllWtQK6EE3TSFPORproGGxlQekR8KRgQy4htA9/3OCNhjZVfIVbST9lgEjga
pkD/D5fQB81ZGjKpqcSEBCcSG2EMg8mEGjMlKMjhNUOGI3978FihyR98liGexvU6
WwE1maFxKys3JGSEBDmiSpqkvcxO5Xg4mWkzkY7bwVgoJOBTxY7t6LdS9GV3s0oG
1KbSbJbvpRTV3NJbzJVDTE8U4XTThlvgyLX72/sYuCU9fRTuZBivtiHvid4pu58s
igo6L131XOoh84kGbk9jdfGrndGI/WVvKWyZSfMVcon7+SnZqe6Uvx3j1rDVh2o+
sHyEwJy8P88N1SdVasKzxzDpokbPbKrCabcyMbHg2qBzOyZlfczk3WjiuYu+Kj63
+A5feLvYjqQL2HwqOY99zm24I0lizcqTH/i2i/DL/hIvqWR7Y5qrzqLIDT3baTVU
vu3205QgduQh0DKfAReEbvD/6SKU2myuMl095QV/hvAVy9BkuqqyDy6HAdWHYsJy
ui2BwvWSkAhSYNhh2755AS0BKeRMj6Du6QSc3LuYJJGPeKwaZTTu6T9eq1wnMWdG
fEfwCmPWzwi8jIy7gcJ2/ZTqUW5BLhpjpAGTV7+Yd3KRiiW4puCU3vatjzzRobjW
M484m3EH7S2emBF0+CEcr7NUk3GUhXXrW+ke+ltJxJRp14B+TGuFsV3Z+U64uAMo
mgYQbVSFlI+0rHQBtVN5p8qRSuV7G+Kim/sLfizFtfdEXjLVry1GydzFP6sn+cQL
0TeLvjjdpta5QtGQV2/r9cYMekSyJMR3ui+yShyUl7SIcszjXCUI5W8QZLAsIIM0
4seJChwmX2rrGPBjZWv7PbErEzb4ndZQxChqBhcAEyZky6biXmasnq5+0a8wzY/J
MshVCe4Ce2kX3UY23BC6cNxz7HuRwGHIMmBvCmiuYjUvFp7DZv5jF0W9zckkoeOS
HWUl/HFTFcQzI0fbnw278iVvaZfBC2+rbc1d3lGQxwuyt0PYkjPzhEoF8S5duTjJ
oBE+zKDL1kKcUaCZKWIQTWbtZ4Lrf07ibwAHPAwb8Rr4Owqu3ZUoXMJsAAeVs1BE
gU6BeW9s+6t1TtTBZSgAwZ9svRgNBRmm+VTEX0TXqlJSdVvfEcnnBCqQ2VsTW8tk
02/OlGzXXfaGY3tUwyY8a3mScC5QLF5yywPAcJH5jvrAjs8U71Iba597qV+NWpIj
SEb2xcppnK7wbBw9v9/Ei6wUdmCEpF9EF3Qcv30ZzNV2NpS7gXXAQVrZOOT6d+Ao
mksGymAMjrRry5pLASmRTQfINhy8WUcNUOYMfguMmqYLfbOcMb6FHEVZpErsTEdE
CjyIvI2nzahacEAUnkx5NuET9JXre5HS5xpLgKbQYEvGzYi1UTBf6BFNXucprech
zLr28WlNJxVg2TtCvXCSyEbXmX8L13SCZYDjEARhbc85ESAZLry+EReGjEAQ//bn
SSX+TNPii9hodtbPj0woM1HcSpY2EFNp/FvAMGco5Z4nKqSUR/+7DfSnGvf5/ts5
e37l2k9SL5RLePPvKgqPAzZSvZ1kBq/ZEEBvNegKrdCeo8W2vlwsQqU1zXZ7r+Gh
v9enLxqQ3AsTUamQk3WadqqmrQ7yclMBLrB/jkSFW4wJrqVaS9pUR5bDkSGtKEcZ
7CexsqPpJzboM73u6U3C0wsg+4ta3yhv9WbzTwfTfR13s4Gfz5EEChMyVAxyj2nm
OqNdOM+4jdfKpU+HIGbpT0GtGDcDFReif26ySvEdey6t2JvrLUQaVB6/zglOQcWT
XmHVzS6HugDU+KRjBJQL8vT08JMOK0Gap80NNQ6NgKgslyYmxLLpJF+L+7wUxREI
M6TBE45NauSrcd8VGZNUahUnDfcuDUue704A9qi+CMLMmpDtT1gbD9ebaOKaZtdX
Yf8bbOOJYkwjuStoE/ktaP+HsNgXuTE8FF7PYaL16SrcuWeb1iLokAwGssIe7/pv
mAOG92xq9dtkAHOtcqjznXY9WmZy34WHfQ8rH6p9DbbZcwCLguF5fwA5tE/QZOZN
dOvTm+QndjrVYY1UglLAVYE5KA/logLwsGDdWKnDC7Nd+8rE463WAheAuho5GmxV
tjOe/klCPpfnWCtoYA8ZLTU4mIEEX3DCOLTisb3XZincsOvzsqN7y4XWp2MCEV0y
wNGHIFdB2/ls3XLsgRVcJvHUMLpAnFqBnHuXYiM+z3Uf49QZLmSKy4PM4rm0+CmO
VXq0PoNC03tzsnqGHaul6CA+eMnwlgQXqSeCNM77euRKCwWEUXXosDfW0vV/V/5F
KwyQmvshjPh/6QZc0R9spYkqZR+63W0f/ebDOey55/weGDFS/k4tMumz8oMR1Jth
/Vwt44ho/SABJbDbbSubjwLn4SDCa3vbmvb1ma4qROyiLcRxLvmHwzHYGTg+4Nbb
umORU02uHgXZVU/rkwi4wl0C1L0XqKqvy944cFNVYau2qYUm1vrkwmFYoBHoqTtD
nCwAGF9T0LjCbfXMcevWqqYXcNqQILspJ4tgL3cTBnPHdZkIXElPYdIfecVGuUF7
PMd+oXRqqxCk3t6f2GIA4YwrOTmok5rEcpSOHUTmJqxY43h/Db0Ie59AlyQ3/Xnn
2PKPgDI8hF+NtVITb1LwsddjOHRQuCJX8U9fVQmXUhf9WlWFWFNX0l4b18KpY9Kw
VBHD/a0+zz4GpTt8W/NoqVqCbabLAth4GPJcCRoAGtyXgAQHn1+HorIvyBTBphds
grlpkwEaHAo5zHfsGbBCzIKD9CLOwJn5NZF6x1b1+Pj6a7Fnzy6qXgFlj+mD0bnd
J+NV27fjqai/BYz32FYkuuZ2HDPeWIVELTneZbgMSn/goqOycunU204mbIzFt4s2
F1BbKUJeWlRkdGlG6ZIRwK8IIYULdv0fSG5vtUoUDE2hanv3as+XfMJhmbuYPS9t
0sAqcA6p+whkwoQ2we98b1aC2cv9Hb24XCPpQJ2m/XdzJNZiJ2R0zPT9LhPVIPqX
BzZefZjAHEsDmHm+wNmzBTE1BFQUjAHaSzW/62fezc89qQIr4D/Ebm9GN2wYzDnC
Xzmt2BFF95h5ZroA0ublVY/ccprzULA+QWmpK7XnhA41jbGs5aBlRRP/c0NYdcZI
PWgVk+kUj6nbxpVTa3p8X68VfGnpCNEH43Vl/vxDWR700/T++IYO+chz2Vh31P9U
W7A/KHAQPMNRFo6MnJo3RqSdPKSCjAONr4RMYJ0ir4r68LzXcMRIzm5OpE/VSqi2
wB7YPH3Xjh9gJVYCWRM8v08jMhSB4PA6OuCd214hJ6BGhExSxXX48owq5XH9csd1
jFZLJjDYUKMyR+7mMEi2IH4+p6kVClb3PnbyCrVVPYwH/gxzD8BrFSWFiWRdFann
5rLj8TzPLNvOY3959EQTbjwkoMHAnELqaA1by53BrnRlqIAD9SNvfQR1JlWgstw9
Xp0iHo8RBdY6s7YvAld5UuC7y4OEbQQZ4XG3KMjrWN2u+0VDwTsrRjLkSkbhAOHV
KogCTukkUkHZmBThsgRibE/0WzrauosD6qeSJ/qdjZYXVZ7B8wQ/a1eEK3/olakr
6IVgGfPjdrtJSowoHykdDXuGu7ErHa/F77kihHmdcM5IsoCdtk5zoxAPM1XM2RvV
iqQz5Qlu20k0qMiy0yM5W9966rhBU4FjL4Bw0m89s1fCi0XLhAHEQluzxBjCjduX
yy1I4N/4dXp1PkxMgc54mhQuNli/j++0vEeLAO12s5MfsqSfTvTNPsBuGt7hA3sK
qXBWfK10uh0Ki+BHMwhxArIF9ez85n+znMlx+rlR6mWp8l23aM+oRONbNe+0OJWi
R+NQO9fpfOKHfINphkYgElPKImdwNzjx6IAQYeLtE/qRws9BoZGahZwsW59sRqDk
aAMc/G1sd8CjZYySdMBeHIHfFquNuR2fsSX1jhNNxz10Vd7aSy848m3VnMVYdCWE
BGyYtXvo4Zc8d/hWbgUnuw9iO24+azOiROuyviWJf0XGi8pb5sJOXkjA1VXsZFyy
uQ6+ePWNk2hEyU2DAECWwFil5+uufSAo5Dqu1DAHygHn3281HnQRGdXsfg3qtYep
/DCSzRsWcEkPYd/nxYBqxZuxpJilqKqO61vFnGVPIdfRkQq4/lYsd37aiiNrbrYm
3peHaDMBbds9z7yXCNd0YHMGfGnfFOGNseqqWzhdYn+jjs3qNlq4i9RaOU32ruX4
vbYWAR1ZMfmjsQfxQPD/cWwVSfp3CVZ+KUzUuJ0qmfrhtMJy0qcPS4EwJm0NeZXJ
TIQglGKBitF43TpJdRVAnSgVkh7wmQG3E0bCKw8jDyR3Y9j6Q46AG9RYYIcA94jm
fT3jiEHzLc06WgrObUdIEOL8G/ihAqZd/ah5d11LiSuEfmcqWl1x6XN+9YdRhQ6Y
Kd66nPabuEtOduFylOUUDv99Hiir90tyju20xKwmu3ycJ5F6kiugDjVmwe3yam8d
3dfOyaANl69pVL08IF2qHWJFJpxPhMu5f5LIuVk+KP6bDBeBNHnFlRbbXySzJ2lA
FYF2qSgdE/FQiDmf37cTPN4G0seT7MXW0YS+AD9SZJYgoX6t/ql0YOwAyakRTrIt
+CBnneJWSgNw4lH0chssX83/CXicxiJoV6m+OvUubFb57mNPVxMYf0SCu3kNXIEn
RN59/ndsu5H6pqpKiG3cvu8MwmP9UM4Ia5IhYkqZBliNAla2OH2i4yCnxJYFEWhx
QeHkNolH5gEeX6fhmHI2zIQSlTmlTtWJpEawH19ZjuSWbcIeFYebOFYpESmOqORm
rQtUA9JHjr+IL09i6qLxTIX3Kh8nKfgdC9YTKCJbU71RCeB4qrHi5iC17wKh8uFm
yllCH7Or6UEyHqDp62lcAKdtPQ5VYyZjkVpc1UQcnSxJJMnzq2b7h6vFd4aQkUK3
lKLrbigcfgV6phyR95/o9LFlD2n+mV75YUfUODsjcefQ/aaWtn8z6u+MtVfezstv
CI5KpumvpxamqhUSyOz0Ovp1lBVUDAKIPLNMPTlnXdzRzNxXkSOGBP+xdQ//g89+
PCmn0XTBnvIuxDZlOOvSirKXM1jMSYiMXtsN7HX4ioazlIy0G7TKdc6TCXXXlFo4
HweQYfnzo0hQTZfNnVxuanwdWpxW2eNucIxL0M/3yOizUfoiVv7pVik3imZBVUuM
80K5DufduLcJGB2YZ1kgCuKqPYTBYrBb/35u8IGnyNN+y/OUQN7XDFmKSjLaDI3C
ChqVlu/4AaDPtqJrbr9K5ZROAADPtCIuRr0o51B9C6+6mHgEJVHDr17KPhTw76/n
Kone0SOs8lO7nmmw13Wk19gDyPWrPOtsoorL/kxK3WnRgN7jrBxjwK6a5ZYw7BXe
9BoD4dWM7W8vLmQaD3kgCRf3LBtw1kVsyU/vOBrRpNW/JgcnwWuNcLL7orffuiTm
FuLTyzF0CoHYfVeAIx8cJjVA6Ho3oRbBi6rgPpjcBo2V/U8gYXybLDx7O4O2lex5
ZxQR0ClBCsejyRQIyB5KVp7VNs8bGDPaOtuL2+/pjPmmDnkgOU6rFFlBNGkTcw6F
OV+EPiZW2e1iMLsfuo8/T3Ir2jybc2JJ/mPwt/WD7F0nuzIyI9BNr6tl6P0jV35+
2rZUfcTCJ8VNcsKvFiDxASactcf08LD7eK8NyeyRWvrKmV0bacK2Z5owoD9ywzw9
+OOwS1rdI3fHTuMB8WT20Zv0JvK+38prIC/vMgNQG9slnDozFnHhTvy+2s0F3N7F
SKpm+7y5Yps9aw3NyPIO4CY/bJXS8iec/G2hpKpvSlVp1Zwfk4ikQGWLvz17X0zS
2O5Unx+1Rl7etulFxIa8IvV+0aaCeor7eE2wXb+rmvDKU/pMIAZBWVFGDOnrRU9c
jILtZ6o/xYs8q+IeLrNDEyM4dOJlSyh70Uke9X27KrmNZnjSYluJvA2fWKnJL1VP
yFtQVgMG2pqSUSttWXHnZ8lbAl7107FIAHw6TREskejOUIj/5eahsh9PIJ09O3n6
mBF6AjwRuEXOIrAG4/mh1Q/jjrIBHfeToNpHtuF2YxlMRumJUg1bgImF7hC3zFLX
d3iazt5HXiWp81N5GejtcvgINr2+6Os7FG+n9G5T108dnKJgYH4+Y0/VurrZyx7K
bsGoNHo1qMDkhRHqHJdmhbLZIo5J+0/0/W+q9VQ76eOZnlbCDR2/+eaYu2oXAjPN
uz+vph86WPk68k7b8cWDt4IpfxpNgYSDDfpE4vO+qtbDFvVX+O3ETC7GQGR3ljij
HIiJdS16bqbciMmuB6w9a7fKhRpQWdd7qStXDGSv1eyu2N1EAAaT0nystACvUoWb
hEIz/iNMTNN+WDg/kdnOg7g2ntCuZccF7pGFda6X+JEh6eS3h0pEc1MrbrbFdxAe
yTI3mLoX5J2UugxTugj7cU8WB1cKaya2RKPM1fYDKVfjHOPiUr+dg0Jec2HOLMGh
+OKDdWD8wxHSj87EYdTROT+4A+Fw4Zvo1ow5noqK24ReEts7guHYFqEWJw1dCut+
8se06Bt4QtERifBF3DTds3udWiHVkJyAtpKosOzkSw/1rFQwyrK/dMeXn7P7ukW1
tPBBjdd3Fn2dl5ohTCJGTAO33UWOWk+lQuEtidVdqUOZ02rvH04tEwp7zCFxpARE
mYD6qH7Xq+XVt7NLMKxH/auu9c3wiR9N6ETw9c4GTlm1WR/iX5HE2mWGJYxe0v1j
f0uYrArY+9O+Z84GL89MJiKozv1uFGDkB8wwPepxtbQbsTEZUlD/nmyxx0/b2S3K
dTzKyyMMAbFCLj351nZlsXytnFOoPfrq8rW7mk43xv8dXprQ2ctELM48wryIxk9j
PXuQSQURBrmOIbq8bvZSMfMY3YEN7p96kVh6PRcpXrD0zwoyE7YdOsDA2fRqkqd4
nNiU4GOEM0R65KZxDdcrNb8/w/uWMstbQsCd03Agxed4MkIx/Z//6oHo6FmRsUBw
suO7YcioUt3JAQz3jGaKdKXUUHRlhyYmB1e4O6AW+xB9ua3UuhWCBD+hioWKrlh2
IPtfzrdDHpwtv9QBaxPHRGMRSiMJphCpe61G+j9VhRwZ0S9WkDlVXUz02/EOXXWW
4xni3wcIJBRkqKuLisQ3ydK5/T0QyD1K6dOVTCj++e4ZlCge37Z05xHDTrNXhmy2
zoEWkmGMtFX1DrutRNxmZm23UwA8glTLCUM2FyfR0QRdwJXCMVnLbtWcIIcGmPJW
c5Tp02sSjqrGw1licb6k8td4g6cm3RiO6Zjte59EOcfacjPfB2wHQtbb4TIuYfCO
pC6ayruWgoLLeoEXjr6vM1O4C3e07uNwKy8cVpvSL7gJW8QwAFqL1fiSEf2l6kLY
/jYovlb8e+2YLTN0ZagLSeV+XOwgac/H7D7X7b03LBud8DLSJrCd9KZJVF5s8S/K
DbLLJ3bNd3iSXLtdrbONx+VIJAZ3dxUWtveVrPEBRNzVxw6oqP4KMzT3sOwhery+
X5oZGtMkLE93FP8pFOQPjOuo0WJR954zZ89LZTeF+8IRr+aA11xCYAlgP89N4/+G
sFMS8w4XVHoi1q4eZxbojmKviVVWs0j+Xw0i0o/3e45ynInoS8RcU85JJYJvYiYO
aS9IgDHqIqLrYG3V+EQzx/ar5ug5a5tg/vZzXAbknecC19PNIGJMlpWfug4sEvG2
/rvZvhmP8X2xb1Npfq+zWwCf7RA5OgORq4Fw44Od3vNB+6WEDulbjzAYJ+zh3Gzv
WoXKig9vVlUxrCVgX2ORqjrrd9YG1xfmx3j6IkKD+dnxVed5r1aEvGvaP7qLpH7Y
LbYxY+Lz+vAKBXBmAB7gEq2B8FYN8GpySX0hM/etDfHvpobtmhwJtmm0LIyCbiFM
b4kHdF1PDp3uFS9KKRh9W1vTLs3i9bGVfKTBnxPuGhclInFK500tj2Ai9HrNghYb
NyNVpZ4EqtvRVMKunnllNtFfZvO8kFqgAKGIQrQ/m2kRXy+6TloNQ1OTUebYfvmn
uCwLHiNNq8vb43MtAbCDLbBVZCfBskYOU5dCgzjYMuHGHjMJNiMvm/2HuKZXNZB8
Do43dc9LkX5ImB3PPXeBGvPbQmBPgAvyo5S2V4VHc8Ybvw9lzPFRB4uQ99SsC5JW
5vnFaAEzlAWb2YazCaILRER3Dx0GdjuN0xErce0Asx6IBsruqFzBy2OPUFXDTwTo
nFKobPwlK8XrUrOiAUPnTAxyAlNpZ763JPU8ouPu2sZm3w4BAkwSHmjCQcaLA+yi
QRe6f5Dd//xuB598K55O9CjYz28q/W21QcUQjYvbg/3Tdqr7Q9tJ7ttBxN9Q6knk
Fcr4q/hQ4T/mbeHBs9UZl92U+PFsnqxsFmgNoSBHzgthvmFoXzEMY8oxptcNV6d+
hfGIswvpGsewd180Vc5lPzxMSF2QrVUS/JgHmp8wBCpThCbgp2Jxh/PTiQKFtORI
8AiWd5zy/DGjfS2GqmX1a8ugQnERO9ZjY8nWGZzIhb6UIDSFGpjIrQtc6708r1Yq
aDMGZ87JPcHnA7Oj1KgRngs7Uq3NfmaT0sp2RxnCZ4qTtWUbNiyR+iKynH1KL/6t
6O/khVcgOrtoGL6UaxQaid/1oMhXpfyDCBmwUKTeu62feer2t6M9YQ6QWFbmeZBM
DJ0sTKAQtNfBmRLe3j760ky12PwJK1URC8FPBjVlxrDPqJikEu7Ki85slGYvSTDr
fpJ2T8WBUK7jZrsZjq7a/5KwsdDHGFoUQ5Lti+1dNv+OgJP2IwoZFUEVRpYYszbP
0FCAyE6qdjvrRrHyUEJMoboF6eI1IHcff7TMEZ5MBLMDAyWI08SN0E6nu0yhB4Fo
CRd86WxZIZQKXRbYy1+yI9E0PrnQ6HYfYoX2b2bAdFPRT0r7rInUWfPRKQ1q4Lgo
wqDCvZYAZC76ymHURfA4rsFhL/8hV7hv2MRGvBCpUndczPeS7lvp28Sj3TgXU/XM
qRPK7u8MM1wE6+q2uxqaFkjoAM4QwWHtQHgqxIKd+d5zMhaNw/JK+MPc1ujuFJnF
7x/Y4hwd2HkbTTM1C61bOICN2E7uM4ICR5BxqkeL+a3LqwZ2PzWyx1kMiJR6cXFA
JvTEWf7CEiyf7k01+dd7jv5MmhNCysBEJM1UnEs/wbkOs3LpzbEAQqb2jilH3kVv
ek5Qd6PtFfKItSV/oQuz7AMuQoIUbFi0PT9rM2BI/lZg4y2C9Yx5HjHagdkUjdww
p5bPYi4Xqd0fQlt7eX1m1G1f6+Sg+3nDl9S24XNofvYZg7XNQOAG8QJAY1z5Ypbx
MrxX0FTDd2jxsFfC+dgSP9IxMN3LqagNvKYwir0lRiiV//I5JAIFHJTEA0dOsrOW
Qbsg29nHmrz6IB+CXaCeIkNOC3SOYCnLgdJPR+lqMK/Y+xAZ0QJilKaYHHGh5PF0
wPLXNtXqvh1IGjn8duqyp4X+W3mOhnz8auUBmS0cr/KlaXjN1myNhDby6ftZ5vIO
Pv6LM+pN9u4v2PWZyMX5OOqST4yV0eCTeNbKMd8HQtB40eKjlrTcmLDJy0cW1IUd
9mn78d+uC1m3nSnaf5MuDfaD+mV14LkaE7uctRoiA3dmD5cNGQ2V9u/IXP1D+heL
iuDUesOdsuIu3LafS7yX6EC21Sr9C0Dt43pMvh3GKZXPDdVZRO4HZGB/ci+XLbdg
m39lbLjHc8TXeQLtxs65MZZofIolEj3qWwTwHH1Z6cDSsrR+sc0diobAoVVUVmXC
Cz+eXnfxylRCIqkyLIWy1fc+kb0jbptlzSZ/4R+OVF+b8fnN4IsTA2egTbwY1w3a
0gqZ4LICAE/gMtg9nPItACjYaJA65BVznws23ZNYuirrtghurwsWkAcbcyk4c9IT
GOqPvwfwKYcpnvNjAEvtZYq/dv18Md+gP46Erv4YhDrWiNvBFb7qQpY8ycrdabWm
Lqc8rtXHSPgO/sfiUr2cKlp27brRYQ5nD+6zie8oXIOThro1FCgNm+ozxBVy3Fhy
kWpYU5AT+TQAuHAYCHrB0VtseyVKIBlUb9wPr7lseCDIWafZIxZg+bRe4AupXjxi
XqatF/H+PgyK1/PAPoVEagYflhjiiX6je2rlM/HiA/7XTz47asIalMU7r3SsfMyw
gUwRBjDxgXS+Vt/k29pTw6EnXtN0iAbLhsxVLPiC/OnDgmde5lrcme4cfNQCo3Kq
CTKsRxfDC3qZSDZ5xKby4j+RbpMH3D2Twmv9hgTQIQzaEATgKY2dXpnxIxQwxoGq
NK5sZhfAZDT1KrUkhbw+cI9N96SlOFfI6HaQovnZKosJrGVSmThCGHyjfjOISahY
PY59g5PLpMa9NYDxky3KSx4FL0TUzq1Bd3/9u7ife/BKTus0HkufwHQCfTDp2pKQ
ChObm7V4T2hVGRag6NMHzWe6ZyFWdNtMCh0SQsNB91MKo4tQ5r7rgNxL7TRVvhLz
P9p8ZI+M5Si6Hec4Sf0MFtHvvcOjS3tIsSKxTszyhWzUHBIu0l6vqTLsI2wXCE7g
KajIya0Tw7UD2ndYCuLpJgzsw+yw+/P/MRbznIFpr47GNFABFPuhfenOb8NRRIcd
gq7RQ2pcsCph8LdwvmngRXZV+jke9B0KpMRdw4EWO09g5/8GpVWjcaI3rnnIJweo
lWy1aGTWWEfTzuHy7Fd3q9FuqkQsu+5AXM2v5c4OH/lT25zG3L3HbfBETU8Tsa4H
yPGq3MmBNCO9f75Xlbb0FV5xh24RUtvPXvISb/5WvSGWFsHpGwsPzcMPqKvYJ4V8
LyJDtdwGozQTDfNOdtSrFsPRTDjf2VWJKRnJuHrl8h5//c7A4UD1fiMR7b9Vu5kN
bqOPEb7/uolEqfcLEvYnNmhDZOkbl+3wBhEZfB9Y3EvCtdpzrrTAKH86hi52U1Gy
yQ+h/XlZR1a9nvcYZp8vN7zBRyQOGhPufGfWR37B9QpfkBTU5Zg6LspVMPfRTFBu
x76Yu077ybHXQoEDtRE0F7adueNtCS/ZVIy4E/KQKteYysE6vjSczL6FGHnoouwa
CY1bAkDGDj/QyOACZSENKu1PlZcb0bG1KvZNuy/fYOZ2A/H4xz/BafeOmaBWUopZ
Dan+LfZ/iHtQiP78ayJCasQsF66mE5PX2RISncqGsjX+WcsxCtjCUhLebaM3pVSZ
hQOQ1Gev1Vd+C5bieuMT4EybmoLQ2tUsXKhDlnRf1z3GTy5sEMEW3BwkR9XBb9ho
NJiB3OA3UHnT+oSoxslMPkmtO5TOw6sQHfUqkMw1hlLc94ikwi2SnFVJoaTYZz7U
93hTssQHX2cIjeYPdslY3ra1pj4L/ArN4XTWqi5Ep2Eb8JtZq390dbSkSkh/85Lx
nYs+j/EDp+jv2qGlu1XEvuRsb15OBSoHWbLikNRaBgEFqDWn4b67fs+l2+g8rX6G
UMus179dm+YJAmWO9z+cZCF2nn3SJnsjhdPzGTpglnbU/Mru3Ka6Yp2KEZpCojht
ydfwFrLCRVb/YZxplxJDvd1dTkUmTN+0FjUA8L4i8CepCxX32VQfZ9N/Z5xLyJud
2H+kfbQVuEy1btWcGy+hJ8XTBAgO+IbPoq7CGZZXpSWs+xkUlLL1YhZOjbIw+UCN
ko6HbxJMHT/ea3U89hYhh8i54DZ7lA/2Y9RsLlspJrDCc+zr22T5j5nPvkys9HL/
TqdaWvP8VyHIY4A5nPuQjNapwlh5Hj4700Mbs/XBW/RK/xsDJtS+YVLYGCYga6A2
9aXB5F2NkR7lKBI+os/RTEP6bS7844xV02tQOh00dbaOutp2Mcc/Ht2Bxqrd/tk7
SscrcR+BMq4BnK9lblYbF4cblreKesS065R77ifxTQRV7AKphSoafVCN42xvZO05
TmvP51nniRIoKBun4RqMx+xu5Dn+exCM8PZJ9JIRt4zavI3poBv5XtKrlE5x4IcH
CriiHXe1s/n+2Sk8OF/9St0Bxjmm+6HSqm/kFAIMm3Lbez00HBabevQvBWP2nxcE
NnMkH7IWnufGu39fCX+0jfKrFJjfMpBHnnamx+ZHGLWxzOoHV1ZKacSB090tZsWo
zX5e1PcJxjm3a/FLcikEpU6vfR4YaKBX9NVGKfNMyf9lpEz1m/nMHVA1lKJAIGMQ
xrjiJPT1LVjVOwEAuXzm0k9vLTFFhYqQRncABACEv4vXztRLQruw4YoAt3gUWKTC
2hWd8VcZEqhBeMfogsVY0zWIEkltUFeRFxZE37PCSLWd0AgFjjQBqv1WIaigI63M
eZWjPGQZhPatO/a25HSJrmScU47l7tNY3agtwmuLvhYLtPv9PQ5h0w7ReTv9a1js
PLZl+FZHSN62H3TFzgaa0f2r38oLhHTXc0Cn9x8WEpgnyDFYYBCaIaELeEEtfuO0
w14UC0uI5tlWEQSCitJZZAFQ9ehu9UkFS3pcJwwALaByPjYJTVBSJrGI9qBAfQtg
/J90g0CX6CDUzDLVxU7nYHDPnzjRmS6B85E1hecGkd3S8+kkrQOsmhPxaBIf2GFe
Cgj8XvNaIkMZQaiOHqHZdYihSnAAqiS7ym2m+Sb8RxDOEKKkbfT8aEM+mM2dlGnd
04e2NuKmGi7LzkqWGgcAD3jl8WCvvzEuTNnSxVT0TNtyw2Kw5NZDP8RxmBi7fVwl
ut+MROJuF4Qhf2v7iMvnLaYVkKyuc27s17egZKrom+GqTpIQNHBWRUjnVSObSGOh
geuDFrmjTcmTmExq/e/7YbVveEmH+XW0QKcJbDsHzZWzvXRkt8lXMNXd+aXayNHT
LYBcfzJlQMHVrn+JNuyB/Tu/Ij48iDNC6WprqEfGi79xgSBf0sk9eEnSX6dljmFt
3FGvwXnZKWDgQkvMD/ZPTqoq2X24y8GKIlQS9NMDC176D7XoVj0jEd1yIZ/1X2dG
t34JUy26MSeAizquy+lETr4YSbWKUl39d9PiLbzZQ7SAXnF4XA/6Fr8PF6lCo0u/
pmA5twFIuv2Dezrl8rh85hJzGWuBh0rFwmWht8NVeYgiClJ8w9ek3A3Viai8bOSd
avU/+XqSfhff1dnf7nliHZh8WVMaJI04fmooiAwH2KkPXF//XNNDWmFDX7K373yw
18YfjUh83jHmYN8wQCLm1tpCL8Ac0OvL8WBJSPtRKWCy+NGl+fbzaJF9KNyEBj+c
hUlTxKsAQbBgZIPY8n0G9puinV232MVfH0jhL8vJKHS7cQXXZK9N2oxXJaZFPwRk
BTCCCWBuX9ndUIWhnUq93Bu0kvXbJMfhU25+CTOZastkJZMzFEkkjY5sz84IW6w2
8yRXGzzd4jcgUmVFrS/D7z1E60pGO/RjP7bv7cvsjET3eBmNj5kdvmPEOwB5ED4n
WhQ+CkIE+FGlLWDN1BuD4zSorvbIJeizXePiJHz0umtzacSyyNFXCtxIzBK/iLRU
OqIDoj+5Gu4kzxjwTVpc/88SxAH1AsLu9SvygOovWPnK0E+OBsgIX325PjUGdw0H
bRvQ14CabCPY6fkIxUNJJFPH9/+lfc1R6iuR04wj/thr6CpLE9aN91+p5MbzFYAs
zmcQGFXXnRWo1lpQ1Kn/2Np05kX47NjGfHvDDhDXFyNnHCLkfp6r6DaAZshxKu/x
YWFTkBbDaTnjykNXT88KXGlJ2pPbB77S1dWb3SB/P+Yp19YwZBy7VnnSelj8TCa9
kmA5TFGGtkqHWnKx62NVSR72abHbnt4HKipuMkH30UNunMAeh6o5zqbSweypyseQ
egSD0wAeeHZOTVONjpZa5iMG94POnJa8Un/JQToCdB77ZMBAlJGzHOHsl+xBYemo
q952rCzk1oCeqSoX6q7eSYy8Eak0nGY7sgHyNYd7taKpj3WFF2LqO2WFxl3Brti7
2WepPiZSggjBUlLuZMgpcg/z5nlvMO+vp1EAzh4j+X5Yi3xYq/NFb0ayVxP0ITCa
A6eJTujG0Nf6deu8QzZ6Ps9SFa0fvk9TmPZv4AN3YtWLZ27lL8jQGUUUvsstwHQ5
JAYw0/j483fN7WiH/zoK5WaoVo/13IspYUY8HSFFeHng0euhLmOEeO9/1zelo7Jq
nge+ttKQ0/R22ce7Rlynmuf6g1c0/VlXNP8j5mYY8znGvORP6sn493EfCTsilsQ+
t9q7Fvgrhqmf5B/z/eDqvpSS4NtI/OKpqRbee7I0a6ubicyK9L4PDvqfRxglSHmB
yqRFvoEfdNaWKfPg4qXCcSLZO5uc/JwryzssWU7bAnpUdFdvA6ZkXIW+n0yG0NB6
xJVPvRdicmoJX8xJ67nAYeWfY/DBu+C9HEM7NYXB5v1Z8aa0Q3bZd0zLLHYEHoob
4fh+ihWxtj3OBdXjvG7xCS6zVxiIC8uc0BC/FnHch+KpJ7e+m8EC+4Y7GJf7rW7N
DkXxUCDf+iykukmN9dR5A2Kaz9oJdZMvf+rg+EsRm+8dxUP64y0XW1E/W7SRDGHy
xOIA54vImq1/Oeo+UVwx9AoxpILBqgkMZtvSSjA7TwaIiNF008KYAR1oPScMOwdx
fMAWZM3T5TWygi0JBpSwYcBBFgbndaSj4nIta1ddOXbHDTpuVe4jmGcyWL+vLiMn
juXDiow6zGXZPPC29huYfQNYhq9sAPpticCj7EPT87UaKu97fPihZwJZz/Kle9k6
nWQ0woPYqx1wzTpkOYDFU07qC/s1y9zmOBSyLs3xg/4oqg5FqHxhAJKGhIThoity
Y46+DIqanDIKBVtMZB8bEFbvJ7rRPw2jaBb/HgfECGy2KjYCkVBTkt/DcrhRI8wG
JpdAIIEKodywLcPEOZ9bCJHG0jQulJ4/eZzgNXlr9SJbXSrGFQVc503NcYZ6AX8V
6h3OpxGyF7+hgTg7tg5nsL6mwgcoGKiT7oCnDLpRyWrX4t6UCpjWKIJwH6/fE/9U
wy/N63S+oChMqTE+qvHQ9DGpTs/S02ZilCbFer0uwZyRBQv2Pj1Vhq/QYHvm5qHs
DlkgGW/Nl75awgzrDV0hviENSkJyKLF1GxaKX/PQ5dX63v1OVrW9dJiKkHIh6D6c
QzAmryLMtUmRb9Q7c9gaXhKlDcMOnA5NQt5/zHI9QpRURFv6QgY8keLW/5iM5gAB
XeQZbaMOrTSv7A2raizPtBB1UyCRE1a/ja/v6dTm5gxjYYco/GBvKzs719UcE+Fj
owTp1X9zTy7SIMy97DogBQdoXZY8YxCQfWyb4b6rfIKAdhVnULoqe5RMa7uFax34
q8eamfuzQm2dhIieRt5e3If7XcSWtt2EQaB+ozB7jGgX3mGNyJpM8otj34EkujtX
ZhPba03jWzWSlJRcwNeDafBlYF84XK2GpY4eIdUhmC+uVL7TdCjQXx0IoLR9rRQG
zloDOv6gse/4jA1wvWWY9PDW4WYv0o4MhEIS/iMobSvbLBGM59mVqv7lIYh/heW7
LOqRfZtvWiAUhc52oYJj/tZDMgiu3NkXxt4h/Bv12scNji7Vz5yM9kd/JxW3sohn
WDkCb6NQ6FY+7lPn9DA8iG6tVPFJsBI47IQlZo76gA++kMKzug4LCRfIc7eknkmk
9olUr0Si0vjiLx+CPQcU6aCGERSKrbWdZmZ2rGxtNyr6IWWupod1IXfBqYJXS6/J
XDworYtnif6cxZ0S6FDItQbukUUz3EDZoX2tAUZokA2QEyy0by5cwMcjir4kw2Yx
qCW3uOdqr7wa87afXYzmt44ZAnXTW7gFY60icM9uXIDy3oeGX117tXGVaGFeXHDH
/KsMqWvX4tSM3NiDARAJVeKlAxMbxLrhW0UbOcgFCVzJehLKYHXQZjXqHbyw28qL
rgeSSUbK8qpXnUVISwUXHyvpr2lYYdv+a+kcitCKzsNA4wK3RuwEpT8SxXS8YjWp
3wUx0vvfdahsP2kRQZi1qy/q5FxqP+90fH5tuEH03fRIgyqPCcBa+joWF5bmJL/5
zBzUwqUDbLbtjZQ74bH/t7WphgwpHfFXyf5Kek+A8BYyIIKe1srbY/1OA0HPYPpp
C9ghCn0SZFgKEe+ZIZMiUeSVZhg2kjp3eQ7kvGTNSQgscU0sZFK4K7+F7lTFxTq3
oRRszXyaurvEPgBou/i2a4eH1WBdxOzaeljs2zCAB/tO6sF0b2nnetfkooWBNIr8
px/ppeEqPAtwl15rMMf1ajjfkpkUGsZIlUFUClQQZ1CYCX2P544wFRLCP77ZVf0J
iX64WzqeQCJxtAsGjYne8WIx6ajFGJeOR55GOpTHT5D1ib2ZfAcso3WrggQv2NMO
9VV6OiN2ocA2giMCvTK61EjgmWR/IyQ1aBxJ5b864TY0UJ0TBc3P9VZWhV9p/Uwz
H/57+0ApHOuMm/L5DTzEBhTgPqeiL4im0bJyb599FgQ/uJwk9YIPQoI+Y1NHDSjs
Mm/ON27Sv7+a9yXnBMytvr6a/4te7eJaPQbiAy4vaj+AaiD0/hVRpzsNUkp82Shv
A2GxscqUZaxDv3JIS3OOlcePbvj6MxBWRa1/md4tLZAxpvI7sNPkQRF2GjqTPZmO
6Nl7q2JuZgMG4bQhuYnVXpvosUf7Hh5Y92Oj544nT32dSGnEejnU2RVZILmd3iZJ
Nok37FAIRAD7FkXEuhV4hxo0fovbyrLw5IZJ/4it/l/5grTG3fjA260xhOpeEQqf
k/ENJa9EA8AgegTphVNy0vBz6AavuzBSLxIljCSUx1+C6ByymSTVaiSFYFHjxc0U
B9AyPE/e+7l1ZaJnK7z3LzkzgM5hpxzq6aX8hlMsGhLT2jQPtd74PxmTEDlWXYeA
okBNziqYW1RmrXH4bWICsGHkihMECoMozIVKu6JJ7Z8ZL6bpJxtSmA5TyHYEqPlG
0gRwDiB6tkCdZ5yvzeI9lAb9GbThAnIVwPjkNoQ1J0FGnpX+F+Nk2Hb5xHkN3XY8
qcQoReW5XFBkJJCrUmjpQStYKtdbovNT5gplmsyDK0qb7MQDGh97hpqUFeB6ljgp
N9W0rAAZ60MikSpXLMk3zrfU2EpXLjkSftkfdfYAd/rnpHsy4RXOekdou70WmJB6
UnLwo6BpomAdDNAof2970V/ftXN/tWgP7NPOYkzAKGo/jiZNcb+aZfWwWfE2XuGH
x+2dmB/dqwvvQ6to42k3p6SpArSxoYHC6t6gwDvBm5vIN6E8PUaWAKrtTxcbciuu
etrGJg9x27DDUZHwbMyit/Tt+Y5Q0S+h39PpDc8zWGRM61/LTz/5Vs2k7fZxH175
++mYMzvwihEzu1+sYamKVUSesN6u8N5/10FBrEv6+QupvXc/YlxOawjkpQJ00gzl
iMrhihMxGYTmerIUyF9vqCX6bmk45HEQKalnLu0h8YKzFVUQYANh1Ho40f6JY0El
UPAtQVD9/PeOIMFCxvTtKWhkCQYoWBJpMqIKo5kMy0mfeYUntE6jgX6S5Yhr+aoE
TbcjalHEsdIxgHSdu4PqSp4fhi24lefqWfjd3wUc5gXh7fnPjORXphqhQMIir9KJ
dWn5a+sgRYs8G7GIMdSP3AOCiUJFqABDK2H0O58ysH/Mycn46GUKgMxyj4LiTDHn
DEZXtwHma9CCMVFiQ9C8NctSpEjJLtNVfuYhOHYvT/aEhGocJgpnwqTbBcFLqbyv
20LQvyH7O6CXf/okOGJW6h0WDyBT/aDbqZKc2LejyigwhFOsL6KCg8hXDx9VZ2a9
OJSRQ7VLWoOMc60EnQFeY1wOVWadyG9rIsU5PjFnVo2XBV4Ay7nTb6GK7v1YQXGp
9C8Mo9PFidxUOEHBhfLDx7nIz4apqc5FHwMdEtv2fVPsj5xE5XqgYoxdOHXIwsUw
fjJxns0UB2G/yGl5wkm3KKGfdcTYcwTRAmdfrWLZbqBpu65wfsVTyELqeu/6IlTS
EVHy3H/y8nTlg4ssZ7ShKk6kIi59ZzWvEitImecNx/FZWAjJS6uMy/3zx6CPgqs4
DSdUpCYlyzpSkExepHqYfy6X0ytDANXFOmEFykqDaynzl8WJ13BHXCAoFK7SjQVL
kBmyYDQnydCQgw9scrts8ZoF7XOwtbKfTTwgBL57dFohIsEvDTMXJoSVIRxNfqR9
Fo6IvZVmazIZVB3qEg45dtP8Qq4ejDG35LoWVdOsEUyay1iHMRRmmQpRO3+lnpPX
KP+Islk+ZEHJq50o1ONpkTun8JFBjnRg0RUhDlHv00py4PPVEVcuHpfz8YvcKsP2
2nl6GkenxeGI6ZIf7ff5/sGzr9qCgmnQgdBQ6bef9h5ivhuJAcYRstbGHGjdy9Bh
Pwx3dDvgL9VWnqYyfrEPHBWgo+0oNEDOenzAa9SAy+RFSx/0zpWmRc7vdIYAvujp
Qlo3eFHrIXxjhwhZKhFVutV83StLHqeMDE6A98KKX4oOupHdPUG4aPDDOH5Ax48D
Clf11U477nSDF4kydcTZavV9LNygycYGRCIeKwYi+cbl2tg7mPKRy76ERD7cU/Rk
d0K60KnMW+vECeGPAn4eVO674fM8+EwAuYfe1ecGT2Tkv6XplwRLb0AhhHgDjjAe
FcUgxX9nzpRXlCztaPPYkWLiIlGwhqfewjAQ5unkY6MtlEWELHcrmwT0eg0vx+Gz
gelgGCwq0y8H5K2biAKNzpqlReNtAFE7kf6di/NHAwuSogR5CXoGrYtm8TYaIrum
baxejCWgWjSybvJS9gt5wenzVLAe27kFl1m9otd1RDHtebeK5C/FnVjDLb+imTWJ
yrP4HbD1HwuTrC7XP1wzVa6WzDM9z1vKr3M41Si3x+/f9fYOWQ8eUXn3X2qSMET8
0TjYwhx2X8isvry/JjMHVrEEBRKFvOQE40ZbNgUR7x9oR6tRZxt/x8e5kyZUhO5q
x1yi72PA8GVl9v2JDw2M7roqi8PRSmzj2eamhg4tzZuYqVPhGFfnJ182Eg4n2njH
2ETgG/wWCQ4/TcXbUdsqPa0hpu6nVaA/owtOcgkMJXFXFe3+1XlGlJiM+q2bNU8d
+mCVtTtBhzmIaTgIHiZWjT1ltNy0qMKPgmWXgmZneFexbxlPbqH/75pwp8D8E/ia
xSol+3dOYuLka3GDc6mOpZ+FVYBbULrlzB9aojnam2eupSNgYDmNIUJfl87mvbN8
a9GV/LhcdMO5ZwCxILKLbSpwqrS95kPZ2EZPJtUkXLkk+rpckyTl+/JLTT9mtsMB
Bjf9FWpKftUDi5N0ovFqC0Y95m8G8K8OCfA2SXGUwMUQp8Urt04Kz3E57dSjpkVV
SsMu5/pOZq7rLtcLn5rNU5RXaC7lewZu/Opxrj3qFWjiTi5vk0++BvAO12Q1I+3v
ufB7LCwzdvIs3ZKO3j3L7xsRM2CIkfaO7uUlwa/3/c9tXimZTU6zw79vU+EQTK4U
qSeyb9KFYzWUdKSIq8usrf2yijcz87cddrUqU1Fvp7Yb8GsnlTl3vAkWV9EYD/mJ
lC6vmLpQAOFQQsmhUuqY6kF9XYd3DVgLRTYZ3y5UCBF9KQe5C3hyVHwelwGz5IJa
SBQrgyob/Ykyl7aH+fvNbHU0LSKp6zlnUp2b9hDNIboKWGcoZPMaW5m1ra/vUhKh
3g2c08/nkT+gSQihgImG2bVHW9pLXkteNh7z9whCS6H7FU0MtPbXZaMozbVKivlq
7bB11cgFLvIsj8mc6RL+lZjBWm/AJlA7HM0xNhleueGOpl43iOvRI6nRhqIrHcSk
wQ46HrnrR55/Rk2ydVKQnVVswgU1/PL54OM9J6qrcAtlvYTBkUx4reaZiMjilfL9
Al2ckBpdM6PVZUfJId2bhzduLsUCDkcmrKAly7FPQolEI0j+Vd952R9MxiDW9E9T
THq47EPo0oNcJ7eK7z19EwFVyE9A47Nrt8SrS9fTi1DaS9ug+dUCvX99/S1jdMTC
cXC6p3OnjZLoLjzEAFzx3ASbVoLfV3gPn8xelovytC9T0cl6tkBUavJ60qEON6s2
VGqDaeowvjQ6yamf9CRUYnChrtW0+Ex+ikZekKoSJP47YDJyhwMrGCZzEXQy1cTA
Q9Oc4D//qnzsec0fnAB1BV172cHwiA849Ib+DiCejSVl/BCKp8Uw8g7WfLbP9O8f
cf23vcUsJnRebo2sDygyg1igcyC2taxe8rqp5fgEDbpwAGdZDDDENVotfOZZVhSV
NcGymyBTTQ0nSQO7kOXcJC0zzH1R9rqGgrTzWR9f/7os9GuojpFMLQi2OIKQp9hx
FW4dXTHm7xzVQcbj8NOdi9nZylfs6bzdAx24fSfER+ptp3cCc48t61T+xh0gjQ7p
LGlk/lc++GRunVhGlHcbf1RDBteDjKV5d0aW0tcA6cdzv6RarRs/SMIB3TVvNR3L
He/J/xp54ErnUEGIniBAPXSdussUX68qnFhorDRBZcjwTjQaToEZEAEXg1kT4fnx
MLrhNoSz4mR7Af+aCy1GIscX+OK9ILwjG5LFzJfpzEUsrXRBN226NvatwPyOMbWJ
BUzwVYRti/IMJSy3i+UIZZACmF+DeHTJIjFa2n4bXF5MRjuFyTQlPp4xax+klvkk
QtnEDix9uny5SI8By/Nf0lBxXPkvqJMvGg/cP7F15rxcPHWFYKvd5JKOiVCwDeHA
QoVjLEza321KlZ7SmXMijvoEWQHyZ6gE7WdcIZnGDmV/IwaPhfBJI0vDBQ7sRRzj
gdH4usp6MuD7TS7q0zZAvmwB4j8PFy0YJNAntDfDfuTsFeW7B52wAeaSEiVO0fR4
VyfalgE+RFxHhKqT9/bwLhv68+9cu5ocG9h1YqPVUr5wSw/BK51a1VaHWEN/ikEs
vWADj4Cw7zl6hlPd37YiHS9NBJLZZKEh9MtTR51OrPKbCVxG6hkdj6Mge8t0sJcY
+ChhOXaoQr9SLHTOByPrgN2x8Lba5BSViiApCAg4Hjo55Xn/6Wi1eYipsDVi30I5
4UeiRBVup7Xl41C4PjGHoRs8rwmjS1LNq47NFF641vPeE1zGtxvbeDRb6KYiYBo0
eWj9mSXN/cJItzWEMg+fAAq2znpVRxl21cBk+HrnamabGr4cgDcEXeKJsUWxiaJ9
bXFftx2ODvQ9Q4jiXdQDl4VE96riUWWrZk71LlHzVk7jWaJD74iZ4dYl/IFLHhRW
8YQRb8Fn4uCik3Sf98jVlajCShR1l+KmRgzGJFDgZ2AXicIAbdxpvUhJmy4NPC3j
dYjhVWwvgm6mvmTSrCDad2NFiW35S4az6E1UV+c09Aagu913iPLjdf35xGVG9GYt
ydbvS0iY93P4I4NCm+UkwMXICogAIuqMqqJZAsLMccNDZPjkusQQh3oIWKUpuTnI
7svBN++/iIManmWNSFOlZe69J4ebVBts6MOwuBVMo3XE+64954s6oG1YbKavSdHR
BddNBpla96LBsKcE9lUCK5xdI0Z+2d2Br3sYoAjcmBEvWRY1AmRi/AtFXjD9zq0u
MsCV4N2sB7sKVJhPuxkxX8DoJSOSCt+b/c4VHWx6TUzSQ5XxxIXljmSI/8hC38+g
u/LAMoNQtWtMw9RKJqJDmmeO/h0VnDK/8Uubbcv+H10I5YThbcuJRzsIU9YvkhDn
9kGrWx/ozm1LjSAda5YwKh+8So5sCZYc/2yE0gp02Ozk5eNxzXi28gk4/IjsUJcb
Zy1gZn5udkKW2aH5/9Yo7ZqkYrAFqE/VLgxYeDuwDt/V1Wn52yMcYX9a8TkFQK0f
/rcDloN32Y2cPT0Io3cSmQEI5KBkfoHqsKYa7PWSTTMIOZ/ixQmLiUDrlh0jX/4x
O18kqrCVB+u4ydSdt8KpyectBceyjWpUx5xywGD89/oQGm5lx5mKVoGIa+/M3uqT
T4AF87ZYJdOImL1y2lgg2BDFzqJBjIEoQAKgmhKgt0A5rSGelkdT9mXJMl/5gstF
O7r0ZNeN5wa8W4giiZffi4WEYfgbMDj2DGMnfda34lx335L6dJNcR93Kh93ebGEZ
6oNmGQRaIOuSef/8SwSuTBt6Ef5ulLX3f/C4+xQ0wN7XnzkZ8g6/FKF7XmMF4/j0
X/hPsYFt7NdR3oWUIxJqGvU7RRFP/vC2HaZjn0vgHYnLlV+CM24G4FgxiOcA6FOm
PwALAzoeweKVCXjTUYgXZ2D1KLl4EG7T3pC5tLsO0MMnSqZ0s2hYczAZ0Ppi8WT+
hE2LAwqIWcw04MbMILcQ6oYnCRR5Mvm51+Rftnn/S+f6An2CbqXhpPjhmF9L/Yqu
KwHN7wZSFiULrzgdLeDiFAxEnzsX5ctwjSGz8uqYnseCR8CJPdn0TWHPaPz8pYm/
f+ByP6yx948F/8W2YG7KWElJDuCWaqk3Gw/gMZJxyS8QoT0h0sXMEhy7QG11mWjk
LrHExeq6I/O01WrAypGmlVnOLH9z+A7kZWfg+EvFVtbCX1Mrvktj+6uzoY6GRBgd
u2G6tTU/ycLeBeHbZtGfHolmECPa1hgm/b4EDUYwVsrUzq98aAXKqbkVQRuYfI5/
vNwALPEleeNRd7sTvpIrpav73QzOlkON1o0GJtFY9gpiVI4P2IgWtYqOww67SDbS
d6qQB5UnGaVrvKi05QtO5vPsgupWWAx2UbOYOJLRP9Dz4rHVh5viIsss9WiIoFLe
sRS6JuEbIOSFbWAb5UUpIlE1VBGIGwR/XAFNQpoJPmu5lAlqXDL90lQSc/2XReTe
mzDC7tdqch8JMvjT8/y1aCgR59qU7kxCgrmZ/SKmoGzydQcoaVRMvm1Om11P0t+q
ohAxl1OPCbatpJUm9UzZNC/4tdr/bDgsu31MWcOEUB4h7bA50Astil/q1ZHS1cMi
TcgehUXPxpSAQJEUlTkW1kIj1Nr/IgpSjXDYV51loNSRSE6ayybo+XPTBShPVlqj
BaywHgjTdpmHB+gE2+NTBnbFzf2MYP00Skr/q0Pl4pYL5+pL5Fx5u6FrdLnEhMf5
uwzZXa2aKXk+sMpwyCnypQ/m7At0/vVBVG/xwsE2qc6hOnsnrir92UDTkCoulYVq
nkI2nVLh8A6oNQ1ONbpxqgpdIU7Ti74Aa8HXHvH5Wc/KhZmK2gzCaSNfGCPIoXlV
RBCYMbD+hZV8J95PgSU0c76jkMb/+MEsxsQzeVwCXljgtHrtjPq+fWJDW2e4O8zs
FR9RxHCI0CxfF7AjiEC12Hx25eCkp6oWOCobFS0sdqBD52tpmLoIjoHc34GdRJjR
0xBo8Z51fx3RLAKX3OYGIL2ZA9I6TtHq6tMYb0iDVkLB1y3PVZUpovfMUfxKA/1A
hj0PrGpr69P8CjEckubi49lG6BFt6sh6XAFTjT95/6kixT9XcAJ5qEkuWav4dFds
A7n3vLypeGIxGkxcYwC4AdbPfOSRduoZYpULQ1amJiWijz0dxP6z3Kp2KFg6UiSa
Vaa/m/jTUHLPT0dYlErSAPl4ptXIMZ/Fu92oM9hShKY967wgHt4glEQ1q0xhWLh5
xW534J3TzUd2KHsYZI6NIesyebmzVNEqKjirb2ymMVWA/lD+rKvQocXgGz/CJtMR
cjTeWeLiH7nHTjACNLBubJh7v/gEhwIKtpyA8Nzr8esm1BX0wWrvaMlqGKvKGYe6
us1pdQoVQIXZwEsqbJux+D4/ixgnABygRiLLbtEmeEuUF+/H4f1+VTFqwNwpA24S
+BiGF7yOcWeVGysB8z549aaiNJw6ni7RtqAiCortl5KdEcI0beC0G5WtF+sLtrDq
L57WIaLEgRZZpW0oj3L6tGSPUiAu4cQUHIKMJ1frGvXdaCY2DVtt2U/CXSGuaLyD
elFc1yCHuDtKRfgL5+zx1/pyffe/vFp1R3gE5ulKLqBWVF89Fg4FShPjDKHoAjKp
gy28pM5rAngWVr/O0CZ1xo88EMF5PH0hMjtEpgn3q9KBPNVmNuKTXjdCN0MNDbis
esTuJmFv2tJHa8CxZn9T1320H92o1iiBu3YaIOK0lSTLnZmDQ0y4OoZPUJ6tG38c
4sbvfM0G/HxlZ5eo6BEOmwHNV61hlt15CPlDBSDws8zuLz+siW2+JUPFomJDBcS4
cLRnJziWT74OmZkNtyik1uDD5JMmoXH/wgQReZqhg1ksrc19KvxJGSlUJ/ssGKG/
R9ZhCE4okxiDmz0gBZrX1glpaTK9mxqILvSsSsR/Yhu22pDDNt9HS67nQMDuhXbw
GaLkfmH63fN5dJoXWzlW4Tb5DtafILsFqKeG34hyg5jLNqbZNfn+BQJFVVklWKD+
QKBttEbYI4bJ8glCvqTEERTU8QRBLope0+Nkuq7pWkSsQAbEpWk7hfdWB7WteB9w
HojiYH/YlkK0Ye6JJkQBlFxJGXMJETwGBlDMLyFvRrFy6BBQMS+RdbjNAg6RI+Uy
V3eY/h9ZHsb3MV2Do5jLl1eDRAu4QAlBDdTXMt7rxmQCIIqBPaggRaDQpLk3gc65
n7t2SxcOZphKAL8dIMfX6fo2fk7zaKwOs+0rDwtQn5xGfgMLp8sRXzIVzxzYGxLt
4yZeH4jYxsaaLUGXrti6GK48PsfJ2NcnXFbP8kMCJSBeZauLFm0pLzsmrKJ+C1za
IkCQT9CCvFXgErbfFO5XuEsF/keHEe3hSvmFV0sFd7w/ve4JZed18+m55C+McA1a
gdPlP45abw5XGvqnxaRZjBYy7VOjK/ObshJXkP9xPfYPOOBsjDQY135LxlLVcMnF
dVnNgKfNKhz+RZC1Ag41O28lgupePk6hVInMqmISDSkdbAuw2G9owuHTr+PrU4nK
5TrLpbEUrVn9T0VQf9gd5G4etxTverLAtuhItyl70d53UjnyLtWI+PxkAeLJ4EXA
hc+n1/sJNPeiDjcnckCa5Nq/93fo5XvA8++UKMgCEOFTOkKwsqs84oQ9S2B8WqJo
rkb62eR1VAmhL+D1fVoqUDlxRrX1wx6aJMVUurI+K9W3y2jDB9fHeaKjTNqEIKxB
RDVu4kaUIWL9XS0ed6QXmTDW89k/rpM2ZC2eimUK1aM/TyL+z2klwZ/cPf90zwfo
oUqAF1b/XqLUTkI0q/OCNC7fSIhOoOCP3yaCn3H9vnhruT68a7g/CV4aVTzrv5Am
qb5Lh2lLCPUrJJNnpO5jyq60UdOLsKxGrmpy/Z5vPJz/shXIUAlz9TunNHKA+Rpu
5rQNVOmnYE5ABmiCCFPtY+Q+cls4g9zx9uXPermDsNxIWlGRQunNh0xQyyHmm9T1
GA+Ttk8OosYq6/RsT5GJWjL/1hNZ5jmQTmT8pwp7WysPs7+jGGy3sbHcm/p+fI5F
iXJGqvcrDG5GJdzYysgQjy4QYej1ea9zyHo3b1hicIT0Vo6eUrhU3oRgqvookPhM
hBHa6saLzGp207NERoW7vavHo0NtvjxJ9vChWVvz/8VBzPCwNBvCwoU/N4foxNyt
pe1SPCA375QHHl1hDYUmDMFfTkoBvFXcjxPoA2TpMkJVvt6yh5pE0Ghnl8/fMg4o
j0umsNaRgU0QuefyFkBAiNX/xTCdPW8A4aV/17vvcTw5OjD9GNUBP3P15aOsSDmX
D3SsuP4KU1sOGZnUCy+HOua5KqhW/BKq2jzg2ls3nNTJwmZBmFXOPVMymXHH855T
Rk6qgrebRSseLp16oUUeUhRxzoax3a1OMZBzNQpXTfaWOJ7wUz9Bi5X1mfhURI6h
/GjOqXfjSc6eM/tOkwi8i93kee4GyqKmE1tUaGA/wmX1Utmn4daRSC1TLL+Y01DX
hEJR5AU4yh4H36TjwJMyDT6dO1tzM4mB2fz4XZ3jJfgpN1wSMgqPMAd7lzEabjtV
PSZIGt+mZ+noptsejfMP0lgdJ3f/8NLJgEVKyn/VRmhD0ycnxNze1fPMIBS9bZfN
e6ADP8XIMB0UeX/613lJ/JQcE5bDZrbWlhV2EtwNXz+adV10iNpyYnaAVnNUJpY7
jtG5YQB9/fCTSxrIZAhzlOnMstNhbz8cYg1c30ByUEqdyNFtG94W6BCP2afEPDu1
dcZ8cnna730OK20oCEOtbTT2UXsLoaqWmJ1hzUsDgRUkfd7jIRyC9DLywbwOUlEU
UPOSJH9vOMXLeeRovdVH5tGC4xa4gBUsqR4/DURJcRKwURFnU7nthAHbyeDEjFLe
WvFUQJSlO2cD9mTUkZFJFxHMmps+CHXpP2YQMNeriJejubs/m4qyq4s4XBAesnQB
MTIAFZbnJ83UItpDPeASt8XJq9Uq5J6z1zQha2LeqIeMnAX0JEeYR5Ed1O20w3ZT
COhuVcS/FE55KWv9QY/knA9rqlindF8EutDZoJ+hmw/C916v+98eHkPcIWHqciKE
lAQB4TNY6EwY/nOU+RvUGTCtxswLtopfZaYLfqoYz6ORGu7dnlNjmrjvliNFu5z4
FLjqHTstjOwQyUfqYJ9aD6ClVnnlky+x4EObyNt9BMqjo5w+VKzx/jQ5EBAexeRS
uOVMeqBIjKMQDmyLHOsG1ePZCWEIuvMqBQ5GgH8DX207LHqhcK/k1aJbHQKOQkR5
nnI3gM3uD0bGH9HVY51Ub//nPoRMEfTPRq4zpEiSj69E9pqA3XT/njknjc02OUrm
nFxcQ5BOSgo2/xQ1i7A2xoFMjj5kBZGozVHYPirYpF4i0woVufDNpwJNT4HDbxHI
WtqYlfkc4H2VynrKDNh5nz//HIcCtKn7MXRK/uteWPTmpGbGXX6z/w9Y6ttT2FLe
qQAPD8LoOCocaYza7MwKDXcSXyNVrHKqNePuNfv9opaFPlHjgD1GZ4grYQL1h8K/
TlxezE3wzs/zCfifGhKXP0kESBt/DFFmcMzDPIqAJ1xeZ+hXUOWY9Z7BVyC3xwIA
RkiretEi3lN5Ouu8PXPXoJ/vW0McfC/9RCVMGfk9wqgGorCS4fZ6pJYVVLar0CRF
HhMUCK78rx4R3eBBxV/wGyIDWtzp9GXp94MpHOzYSb8cUiOeywzR8j/9+UyV3sQQ
CfDoc+ZI4ZLovtzrkjRmdQloIJ4l8VLgcABS+9NwR3jCbhAr9DHPGWLEqTrdP54F
Wn4g536lluB8c1p3jw0HdRz0syb0BuTmruWkyBfOFCZJWy65fSoVWVm6xwtWNkap
Wdf0jNNa2zQK3CMqf5bRxzavcq5CZuEZ/YrsBWA/bwJ4ysRuAWLi/u6FdrOWCuHK
6M+eK+MoL0Rm6JQw44uYTNnGCx+XnMjArXh6H306QLUnAq6f2pQMzRS8Dip5xrWj
S7pQar/obFcIytAkBuMvMoRLhgfYCGYZFNCKbuCj91e58kELNpuHav84NtdOyP3S
3pBlpQApj7ihFekmrRt8QOFYe5SiLBL5VYYIuj6Gu09Mxd4I2aXn3Flr0Z9yp+RY
8hG/vb6F9iKkSA4vkSddNSxak52m6QafRlYky+vE30T5gcFgCKxwIcH7lI3dLIrD
CVFfkYZFYZHgKy3D+T8bJd7nmn8bQJnZHpEsn8ToAwut0tHUCmxMg0X4y0Kn8njV
y4cg3EqrU0ec806uWdNo+Nqo1zg9j8L5SLIGgPh4IXqevjQ07Nej94X+gntt2eZI
iyGWl1HlyjnlKQVAjvIV1DvlXoWjLDpyGzUJxy34ztk5lGX/rvcrdoq2evf2XqqQ
NTYcrhI57M//KTxSwobx2wc0n5xHEerHDJuElQs38pJfWTrs1kcvdW+wgO6z0y5f
YsnUk50YKWKjqePWc5JSWCd98Tqy8QO88ci0YrhS3fF7E85GEWswHoTXmZ12I378
2/mxNj7Ohl+CbdkuPgq6zTmw5I6Rzor5BnKA1sxbh4PcRV+OZ8yGTRy0j3R1vdSt
JDtN1y6Xblai+c+5HWp2LyNTNGiU+WQwnZWSGz0mO/GSY7nG2h2yvqfgW4MVSLGX
Qx/c1n008Qxiiz4PHqFSb8meJUs8d2paRn6LVnA1OW4hi4idyB57cbaRcXxXvMpU
YaSWiRZfESpLMO6R0E8Ab5hVHsnyY6Mn70xulhGAyHlrK1ulLSEYNncoYBfpQRHp
yRx3g1b3SSsXUesNNGAZ4S9noFPd3W0zWVIp3Ke0Z3n9DDn47gnvrLeu3VcfUp7G
Rm40QJ0Uj60I5IeZKBtgdQc7YCN+YnMRGNLYngvR5UB0MlW0BpnD8lUfqM4kYEDu
Sp5LXzYbtImUX85UBeZ/vOO5s5TRKAh6SRXGkIa9SAkAe5d8jWXH0Fr/VHqKIvrb
NBGFwQ1gkbcfeOfhqKjmAUiITLkgGmNF5Iq8U3X3IUcD3Zi1cFVxDJFOQQy6QGUa
fec5c31hWp9IxdSBpUOtbf1UHLvenG2x/Co5+NqlPcOmpbTnwyQB8Pqe9ahVTylu
cPVZZquWBitbrHy5ReSRL5FXJwm4MqAZXHjNhjmNGu2tEb/fa5PxtoovRqXwNFZj
5xX2I1F9dzFy0ENfncTm3Jp1rZPqclscfePPOYR4R+dSWTMvkasg93h89Re+HTS3
J6YoYkOzBCOOgPxWpWKd9khBrn4DzO1YkAqN6GuRJCO+4+r44DnMF92BlABw4SgD
PJHPbeRAkGAiJZ3nGLMimireS0wvzDl24NMBKWTz6nssqnyR2p4JDS5beKRFwJyZ
gd9NpkL4kcZtaRTcxrtFFL/M84NZwrYMbBrRwQLAWhrNsEhWSDDPlEbtMjqM0QwH
N1r6++8mrSt2DRmvRA88FJwbSJKjRDYoawXajg35Dw8Bczk1qhPy73+2e9X5ASj8
k5Oh+iQNmJ8lclJEvb87PAzAbNyeFU2d+sz7XKUloR91DAgH+pKpFqC6oH9blPlo
4RZOWF/iTSTAsVoopnTvXqBhREq9kB3kB8tNpg4PeGKaVcY/1dRbDVXBb7FFo4NR
rHoM5I7APRpKFzD0qbFajAcnRVvCB7i/qZtU91eKWpV/Yq71xPdAboSrQ/iyeD85
B3Y1X7fdfL+Gs1Wc4yQHk5rReTxO9R9BxX8DrCPcDEjPLEqDp/7FlHKQ9C0Ltmx5
5HIF8rlSs41KT0MKr+HL1zf9at7HQqIqApmPUuTr1VbMSuzBlxlczby69kS5hzcl
DxLLjUigP4kAAhrr2AInb7qyBPMSnDzpJSQYmCVEQ9l0QeNjtY2/UjpnQMUHxQrK
OeAIUYTJSCrSgfXRrDMmc4drPjERvFDD8nTeb3ZQujUerJZN1gXtsqLq5tIjpNkJ
h0k9YQfEecgwgECMD4nPInFbvEEczK3sRuRHjgTyHkVDuilgpOADtWwFaorm92k2
HuKfh5st0RrjugOFK9s3V7WXaekLetphv8moSjprz1gt71p0I2ejw6s7eRNr7UPA
a0lnp9/ipzBeEELvSx4L2W1ibNy8WNiZU2eVVnPBHejQLsGTO0jEQVWrEsGjsag8
/+EVDymvwQrwHb8RwJL7fMwPovEoj7XDtpkGZUoT3meH/OD2ji9G1atp+FbgxCi8
01TjETw3YYUtLtpWrKjGFtMfXrsw/QStL9EmURHSL48qsHG7WIAcZ6Wzlz+na2+6
rhbUVbwlVYsb1xEpZPHhIk/kt6XiKfZ4+TN5w4h5x2LtalAae6EzAJp/J9vmNe9p
tlbHVPmfV6VAlCsap5RYQUVgCeNuc1xT++/tAeS8FPb02fLdtYcDqUGXCI0TQbGP
RC7JVhpPXyvbS8m6ETLeLcjuNlK96L/ZkEN/CFz6DHZhzcyO0Aoj3ovS7EpOsyLh
9ajLu2UJR1JgTFtwB8lnGCXz906jOVNFLMS+anEWFgyr645CwQnIH6DxaLBRX1kh
ZykyWIkYpZ3Ay4Sfp74chhWvCqN2cWzmmyqA3HQommZyY2sy4eetPcUPuezUuBAX
51K8GG4J5vg1l+TkPLDatqkYeu/dGBWZZdyQzNr1DPMu0shFl4IwuMHpAWAtqNWW
Le+YUe4hckKqHLAq5+/zmxe+zCcyJqzUYRcZtvUaSBcrVOgNxYagxPnONKKSaQ2u
rVzlb2JaLy2WBTq1X4OTs+CIQ59SPTkddpOOQAN6Trxw9trBw7NtgenCZk0e1j0b
TePZBjNWPG3YOwCU7nuxzyCYvVVEpG/kzuQ21f2LmUhspx65TF4IPmACgZr6fx3/
1DCqxwHT0HR7GHfBP3pHVPKmJyZySEE9aTvcaO9In9OWlhxYb4XDwh16aRIV2idY
00PS1O/ol1BMv/8GdAltzCnD6WwEZjjpp/+7wxfyvpMkftx4tOrRjpWqi/jAyJ6h
wU0zkvKnlzyV1Fm1+Coci8AprFp50BlMMu7hVR2DZX84eJczc4EK91NVJwnfHuJX
r0nvzO2AQeH9IXexg2oDg7DrCbMaC1UuWLf6aZXPzdxk2y8EHZaEkA/bTgHYLO8s
n6QmQFGPEQmxevfhueKYFiGynazNOXGlJWhb+c1p1IKufrGHbSaJ6U09K8rJre/d
T1EL4g+aVRxnXWVapiAzBRglRkML5Zkeb6nhNWAJM6SaG3KNvNEAbwXCnNF0Nuvs
OlncGkDbulyvk3TXWeqcnZcSV6x1jggo1fcAtzE3sjbilVVSlQ2cFigRqJz56adD
g8GqJUFfE3UI13qLFAubsTZ5dosoixrG1d4MwzS7nTMmfDFpMhpgXJ5xohwbHPfU
X2KhMzQfM4QtWMIZJqqRVxM7yZGQIKBnbC7SNILDuKnzUrDckembUCGG4Y/zAI2s
R1tAvG0tNXzqFo4YYlB0pBjVRyhdoekIq6v07qtxqlNIKKAXZDr5BD7+N5T3YP86
7RP004BBjl7AmVSLQVulAGegE+B7rO0E+qA/E3eX04UKp8uGOBm2ZvaWiv0DO0V3
+vVtr7Q6MJHD7i0LO6G4t2aT6is6uQPtseMe7zubw0B2bWnPEFnE8aQ63kw3gQ3K
q4X+5fXzfwr8juIuMtrziT9BWUiVkcY2qkBSJzovGlMKaq8WWwSbkoHTAE7FQJmg
EaF2+mvO/7X7zZdSMZ8RIBBc8a0/9kz/+QHYT4A6SU2E8H2U1V9IByjUupYxLUTk
RB/a9FNpSEruHOOGEvVC8zhkoGROJGnRNs/mMAkk+F/9Nwyhbp72GCgzVckd8Xr1
AZYn1hYnrTzQwabirKMaCBEPwdMmhNjTEfRKLSvWfnIJv3XOEIOdNrg1X21BQzEM
ANvGk6PNJED6jYrrjR6iiUbmTfud3N/XNvcgF+xGoVn94+KrUlKOa6kgKsCQ4/6r
ubBmNnt+P/UynsFwYH1H8gC0HtdpIXQFzmppR6MWqx8HNT9mXOTghuRgollhFW32
AJfwj81rgZtmXVFIW0KmjirTf52BGBdfHqw3JcSp2x3zfTNOufQBctw8C/B3ppnB
vksTphVrKpRaFTwwEwpbVWAC+e87cmyx+ZHq/okt7VgDHBMjLtlsjOhY9Nj3Rkdn
KxF4S9IF57C6Wh++4nkm+F4eq3cp00ZK/TgEgLCc6kbibLfsLmVx30PjJo9Trags
t8s4Lm075weCsUOh2D53Z9SxtFcVMvNdsSi36vgtDT0njxkXEZqN9HiGGt8Yxuc0
0L6/txXirtYl+bpJ8ali28irfKetUAHVdFk8bXYkGmhXTY5jQUe3VYGJXLDc13dW
zMRhl6kqbrOAr5eitnzaOG5ma8gZAM6OceN3g/Fkg7+ZCHOp9B70iaZzyisRCPgx
tq8fYQja9XjP/XK92hdvayw+mLrZK6tr1fv92zApyJ+RVY/bGrsoi6ArwArbKQY3
5yLpwhX6mDvvbEQVRVB6erMteB5Uz4M2cKL//lHKb6i0fphS/v7vOiYp6j2otvzb
EDXiW3JWoE8dXYqxPdtVs9aI+QiYPz6YWKlac43nJhI7+atR4MhD6Cae/bqshKmv
GtLulq8K9N/m8/43vg8SuU5N00bLS3Y2k0gWtkQAHwJpjq4KiT1K1A08UObVHP9d
Qi7Ld1rJcN3I5VprwqUqjPqSni1C3o+9TdjwjxKX/2yxk8FFUISMNDA//IOsfHd1
eP/yCOTkVqXWnUY+PEh9UH7d8pLBlJSrBLS6P51O0WiARrVB0laG7U+uC9Wn9MLM
lWK26lHhvLMufu69rHZC/lOWs3FlnVN3afp0q2yLXv/q+ys+5pzg4z8xjTm1HljO
r43iX9qaPkqSKFtJWX/FasXEaEkXdkgdnQV8oJdxhdP74eaNwF5iZhuEdrlQ2Qlg
6MxylOwb4+CBrIUGeRbRInlp87BEx2CRgyaWVC15z4L+/MbS2sFYQLMhIY34+JcY
7XDpsE26m5v5CmGVuCkYYTPVBjjMeZ/JNLdZD+dIPR/XGEr+pr2BfGVo+ImQPyW/
O5cGaoX1SS5Kj8AH1GYhAWewUnc9oxs+84xQWcXdk32nDv/186Ji0ZBk1e1/Aolz
H5SBPEn3hRvD2xwpbZh3UN5xBkbfh9KBbM8WThnuTi/3Aokk1F5CjIFpXroJE26D
YC7lWwejydl00hQn+o7q2wZDtrXSScPqPKgNJOtvt6CQZJJLcf6iGHwfDKxXlh5H
FVIu2wXfjiicG/56lujY8QtHoiH1knBwDqQiIi0S9Xmz56BcmRElZo0qSyurKD8O
WzTg8CQFBeCK5A9NA35B3l8isrdP8z+NF1YFGv1ZLRbidgkeAlLAB0qEH2+fktHD
IdlfYwdibyeG53mm0hUcSwtPonp47IcwcZBoxQNITRfwyPpuf1RDLPnS3djiJs2X
Xf5FZeZc/3E2Jq+PRrgNcdRzajg21zaVFaJswp5+YbTm77W85xwKWR0jYJLQbhkI
RH/q6QvzZamz/805/5BdYjR8TUN4brYN0DicSKgXYIxqRmEcVHpySpwYCC6I+1OB
oKB8ML17m5t0A6vfbDns1ywd9L0wxgLeBs6OIt9S4La8z7q6d1lynBvjTadj34FZ
lRvw9pGBDMpTes2eKCwiDieESTKDc7xBa9+Ld4czeEfeFvwgkWgFvl30ql2X7+3e
gqIA8Bg4MGCjm2J3YUTKVBAzRODQeH07XdYIu87jbaUJPDNvr2exsi1a2Y9FGr+9
9SzO+qDfFQ1L4ZPrPm/8xFg2Vmny5vb1fj86s2xcORNr+/YOcxhu+V8Y3FMwtsBs
6d2Gtw1msvtdxSR7A1Wwbz4FC1qb1dI2KC7h/4FcWtYmd5RNBmt1InhMHh9NNhYw
0jtB8pPVUpnUL9GA37dVqNY4UO3NvhVHBToFnI8zrcBaQbSwFS69yR8kZ3/+yQ71
90CW66W7UCVPWtlv793QiLmOnGiJ5rlxItn8zSggOQXnmLNdPhX4catS+dWF8Bfp
tUdC3Ro/oazT4K7Wc85i9312tHUY0jK/DYkEj8LIIXT5qCh0IkvfadXv/lVb4tlk
yxeEr/yXlrc5BOcvwZ/c0SGkFMZYODWjhmvbLjRUV8TIHW5Hdlx8y/27qhjLBYtw
YwjxkUgRN/mEY8PCgnBwJlifn9l2PKxWb1BOXKbs3WuqGtlz6LDk9OOaF04Vv28A
3zrCKmquX3AZBxjhTeJJCYhX8X0fHfiyTH6+AOQgoXZZ3krXYEEti5N1G938JxKq
Uo9rH/qup7MLbZ6urqroaG0t7uQhJMCW3UIwN6UrT028DOh1OSn0tS19mSrRwT8f
mNsW2y/UkfmyNIQNwhArz5EM9ehyaVESXqzwWEWM6+5t7kqhOBkfW+glwnzzUyTt
ADBjy/VwJf5hsRhNdh4kdLF6H/yj+VdPVWGsGXjVkbQ18kj3/va8apqLI/cl0hVI
nG6YSGBnVYNLOQ7J9CdjdCpMKqxJ8V1QSL/enzUtZuRtHFVRaqpweV8aRNXqOH1F
Qx6H0eiUVmc0HM26CXHRnh/Att51SalhOU9P3Nagzyl08xC5OYdCINSav1IX7qG/
djuJ0jNHh8RxKo2FzazYB79xZ8iyoooZ/H7dKd5YNhtyGqCEJ/I680JgdpiR3nZN
xQHtbdgH9zRK/z137ytwrNYF1+4CfurIW9KLY/GWed8FAyuocbGU0g6dzzl0As2w
c5f1b8uE0yNV+G8JdriXVny64szYWGDF3GMdx+viPOjehs1CBRRyydvNJm4JwNcr
lrCGmO++k58w/8/FfUh8P9g1Qpjq8FAzVfnc1DR4+JMDgrSkYcmm8gQLfBofTy4d
5x1Nhzed/ccYIj6DodPHzWgNUHsjlX2yiIK3wOqR1CzpL7828MrOaTjGKIPlRLxC
wADrCOYJriyUsKGQPL5YGItvaSaMKmSX5xHepC9XPcYUWVBHVYueh5tcyPmfIvlr
bycx3Rv24Q5Dp5EyvuTMfZK2GBjcCAuUMD1qCEZ0eu1XC/ZbrDpgTYA3tuQq01q5
XomfgXh031NI/zdDQxpE0R3Th7gpcdAfFwQ+yYmv1RCUfhdR9Z20QcD/p1hOlQWf
xDhbrWac9X2oXBPCYwcOnQLGFynA/9Hq6s7In39tl6u9cva5O3X7SdJtU3+GPJ2Z
fwPnDqQlBeocEAxDZd+L4rxXgO7wkA2JBSokp2wQKQenxjOdAR+ClhTwCcNfsxeY
UMDU6AXDRaa43tIVoJhgY6rJP13lcpWTz3jwHKGY3bpN1ALn/10IBuqGaOBcZH+A
2qGDmmtjJAKiZhiKIBqIOawp0A1CZD8bVoC71/1a2gle6jj630vtOE5KgqJxo4Ep
TqGkX0yP8+gDTCIOy++l0NVdSIWIzYaI6Db9uMqjQmFoUfGpZCyJXJWp4eXL0XNV
SjMmPF7UE9UqN7raz2EEkGZM3+dqRQji6JKuwKkCFWf/ouQSodIFmQmIh6ZtpQnl
/i9gbgol/clQnJtfu8O83nymTQo79R6ZHktlF6unMXstzKqPO7kG5IpmsyD+UYMB
wGbXiUyb/sQo8BaChPsHXAJHFLnjnr5v2KPKawdfNK/XyHWDx+WI+Bz0aL088qJn
Z323eR4ccFa0qqLYhJbnUEdFWCkePM6vNLRm40TscVJkL1PNCWxIXji5FhGR5wan
yqgZEPYePe6OZkZ4ctZzyuxHUBsqJm/l4izkKc530iSmnW9rem6h8/tfpAhewmzf
YheY/Ddi6ih3wdLrJG4nE0vAUjXozgBPvSvwK70RtMhh/OCNdMo2LQEtL3TIV7IA
L2o/Ry+Of/2RQ7/IYUHKmE4+XYZpnEQlGqbWWxTIg9m3GtVIhPqXcQVgqZhvG0fO
LPxejYkfgwgR8wNtvsyRriIiUtrwTY5QfQzoIsKcO72vdHC45TBK97x+akjoHc7X
sa08ptoknmEUZ+gncSkVrmDJ256wx26F8u4nKWE+9YVl6eBUyJCL1+patiiS32SF
rgtQJifZS9KyqQPx6+I2cYNaSorOr5UuOaJ14BlCiTB5WBzu7Hy9IUftr1eARznk
eSf7TvBA2pZjsKVMMO0YvAyspf8BLpNwvzNdFW4KmScsYDBTboyaTJsdeHnUNFRC
CU2KKaN7Hu++PED+4DyBlzddhEs+8SFH2ob73mhtNzEo0XspJntb3Z4zzfI1NGu3
PQgbd27HV7mI2753b8YCSD2OPs72eFFlsXJk3ipMl/UwY/HDpbh2tWDYO8ZLcv1G
W9z9Wnb/UZ2ji2atjBKIakTOT2rSmmHJmRRpWFyDn0Ap+6Ac9lBVsiM+USsm1K32
lvdfS6ollQj0Z45G1VmjWULUcQpW7pvDy1jl9+prygjLm4torXkGNwVFxbXbtrt0
KJN097HpIRP2By9mxJbcOAKiqdyeIYvrQfsvLb7deVjKomokRjssbLIxR1i29ed1
NASmkX+aJRS/T/eEuBDMmkV2AC6uiGaxAAPmpdu1Fd27ryzfZq6MnvvDAFHdCcAF
JL0s651SvgvNG5ji2rRD33LHR26eAAsU9fVX6jBJcqVsbive+YcOB/7ieKSfTb09
4T3yppWdypvDo8iTb0gpuXdpFPccToZ25D2RyjP26Dqhrgpf08iTXGLpErSj9+5l
djvJ13Y7FdaDcfBcBsbC3OEzqo7Qgez5gzyvb6BGprr1NVMaPj9dbHybITmWrBwA
iBrI8bHQQv5tDE6A6vWGRxpkkKIhQpZo5sERHqQ+plPOJzvXTBXw9kUT5d3NLLkb
zb6NEXWG41Vp9ASJ6SOEHGYrl2p5+l2KeDRPavpAzlP7LELqymu3x1OGoMxKSdRn
B3/946d4/PIJJ0hbRFzAbGy3ExZ/hmUCVRiASQo5nI83cDEaPQR0dvxDZ7DRfN01
DZq64/LnGdxToRPd/fDa1h1v664lSXj95Ste5uZJ0wkKXsyKFXNnyVrayFlrWw6L
ZFGIHDhINncxqS13YmzNe+Lj2vwPORsJfnPqCsqLa3Q7YCN48ancuWlI9bpuzmDs
2TLpLhszuIPjrrNuBo30DtwSXel8hRJ/xDu53Li3oiZst1A9rzPAmU3PJcMRZbmU
efJ3ILy0BBc7I5fZnwG7dceMf/3v6H1kdzmYNb7aedjQ9MEwGBnPNzKWyxHRFdj0
gtN79fvWgxvqKS+7e1sy1AzQJxoLzKwZdmRM72LwIqZGnecGtWUQsP78Am2MutVd
V10QpmxaxP9xwQ/43R2cKaUhFe7eXOv1GFPZvcNtkfAEQX0ojUJB4xuPxGboSei6
H3L/kiTUfYkyyNh1bsHhkCcM+11iXq4T8IGxZMg3WNAqsTvjodm3TFmO2p1f/Mhs
ibRHJtNF/CQDWBQ0IJYzxZUzzWfXvqBywrMbNTk5BqmpShDOXKzAa8uuu73yTBuV
L1m+A+8CRS7IL5f7gZNFMkHQfCe+cBt1aBikYOGGs96kmAREnGWCq0BCU9G3zYtL
v2yMSIbc0//iPd7kIcFBDb9HM5uKsHOJ4y8/hLs8fFECnUCRZg9mErIsQJkk+zQV
FXzV3KcMwxaaWpfjMiehDPmuBjwzqTgy/KobiazSKGLw1xtBr7OxRRDbUYXRH4Cf
Gxlp2Js6V0Ek+IjUQEdpIk337jPiAHhZwught2nkpNTRmrnXL4RkBD0q0jqxmUs7
xb1tlNJcsub3aoY/LPkCu7V1s6nYM64ZoHSrYtqMs9KooI1ceSX+w7RvwCa4CTx1
QV9VwCSXGXEq0SCjYqmszTSkKbHNGDxgFZu2TIF6JFdrvGpBq0piLP7+pu2HY/vK
VYDtSzRMYp5RT1WoPzRS1k9BFuMwen7al0p1VookNPhYWbRjpEjWxD6kfNR2urL8
1D3WYjUnxB/dW23WILTaHEqe52wWG+u+LDXnRqsjaM0SKQOlIT/nuLhVmYSivJ2x
NgihRxC7xShZjOCfBTSjN/9WBRn6+DozPs3wmtKtmJOGLevI504NKBjYSlwQnzm4
WtwGmHh5aRb1TbshnNzC/rYAhnndca01GS3/zyKh9ehHgvLqoYSzquUEEyKM+BJ2
xm7AD7FRtu0Wt0UApqmBQs3SO62u3N6DDqvcctZwiAgjFM4hpUx0OQoUIziElmBB
SuRCDNa45/Nj77fJkalim4wSm114QgzrvTbnRAkXvPpHtB6wZ6Jb+8VTfeIP0Nbi
Wr20vD1v/mCyziErgYFo1vT8uzlHABNCz5pl8UOKwA9KtB5C6LIjNNMTYVP3QmjO
OBFbkYVPIswnKkjq7QCbyLq5SUDo/uLJ7qpIo47tC0gj31RKGlO7gyg/rOk+KSpi
3GT3WxBZgCvQiSOcWmmHU1hQCu7e20kP7uxzUWBotkyGH/QUZman/ZbS9kjvvNJi
O7tvJWh3MpTznuRN45cNzNumkYdC4YkCWJkUEhMVPZEnRoLvGLpLBudwYACrtjOe
sKZMArBXyZgHMYnmLNnFDbxoKPkkiyXVRtxK+X07skbcCeuXCtKRqXWkYjl3ReMA
Qhq7+dJSqiQxhP8aiAFXnbQZqak//+ZinrIp9WWp+hXUOorSwX/8JypJmheZLtWg
Gzy7M/nW84ETtNg16oEagkQHdDMHiRAQ3j6PlIAiXbiponvaQqH77HraoAjd4T+1
8qVXh5xQWkjeexILOEGF729ckYQ0EWfnX83JQRTKe4DN1H66L4h/I1lk0yttpV3+
6wzU2Z+IC2LxkiEmvijg1Z3jO68ybiieTZZKUqI2KqCpOVy0fC87HWuzOaF67MDa
2plcr8pK9Z0rFyI1YIS/UQKuemot/LE48P1y4H0bvrUmsiUGaInNX1fwVxPxF0zX
qykfep6uI+OzIBe9uj1f5MF9epgLlyaWpB6A2co4nY6Vpk4MRfLCYTKfgMofXH4p
M3WL+iFgxrL61yRjBi+KYF1j0ZrR9kZZj1hITOXPceM/Yp/h6fqWsJ7hejTWouDQ
Pxd9NBt65qQ/ZKjsyZvpQsJBFcT9DYEhlLzPmB2GAQZ+IgxUGTUOnRhPQwBEUYR6
PNSRjEpBYiYKLWlX9IzzSWxPBVoDxoacmg3WItyL+YJjWzou0QbLLJ+WHP/3podi
iPan68DncQSaK1/eEjRPZ/zJ1eEv4uoOQVV8x1iS+ZYzoHTdhjH04//8+FiSiZ21
jVK8J+bgPhmIvao9Mt/M/23J5Kp/hUMrBuOM5UBUlICdBWq/q6CV/Etw1Dpo05rc
MHmnDZSLqwc4IN4lVZk5rTgyctumVFUHVvN+TmvOq+HBdc2uVPyKw0KtJNu8YICZ
PjLumQlLUMh+KS2jLzOFFYzjPnYcBFsjz/ueqr92qpdD47APc++8D659CQbKhqdU
cyvEu/teFdIf785oMK1Y+EAX7+TlNhRvLrgrOjf1SOpAvHAekaYI2UcS2R1WfGfK
J3RniGfNCW7mJ6egymtsUWT9aqsGkCTJMyw8qGlr1mV4tGVZxvjUZ1Mq7p+zYrHl
syWy00IWGbH7WNcgkUvtI6QdGjjRcyw+0Uq2v5D6T/QjqM8ZPoGTi8crTTxxgS17
86OmuEc+hWuoeMt2Kzlkbegpf9RduuK4Le2h39HRAj1L7CRKWpsFI6ZzVObFY+HE
sdqKRiPycrpUzdKF0+o8eT19iK0K5J1Ukp6TNGGvwk/wo5WQVNYx8s9M+176eqi7
abdCOcYzM8HkyNPOFIuDQAubbMOBf++j4LOolBX9sNKcR0rKlv0fq6ELeCnhxEbo
WtQX0jUkCSW3qWLhJlfOqhLlmlE/9x7TIZqtiTcSn3vfueGnvMzsB5A0ItHxWGUd
QgEYyajn+4OTmR/3IxfgvmqUBNpsUfWyxwXIOZUnjYgvdfjHjtO+r4Q8kEtSU/Hp
rbOD/6jKpWz78CSvdEl2BfRRW/h2XQ+NaeJX9KBLztHt5FXWlLUzRvHp8PVpvfUx
rSVyu/LwulOQNKTccxaiz+Z7Md9q1sc79EevaLivcxBeS0Rsfp9wXqgSkSsPqHFu
RJYM+LBzh8PNW2gcrMS8MzBUywuUCJdXi9zsy2bBtWKF97oahHSL00Sy81lx/1MG
mw/hG/rOxWkku2yPsUaTg9xdlwqk5G2ZJJvgwAN0SYDvs+B6c0d7alk5vK93kac0
wmM+8Vy5D8+A9BJw8FS6fdPydl2jBryxYgL2Ipz6ZgemvAvKqEvSro639q88Bw4M
T7k9QcU967RlFPH1y0daU7bqzD7/PaHiWBKknFKOXTW6zIySbwe8EwF487awL/pL
kuIjnZKwH1EAIoLL9a25bnk5W/YVSReRJVfutQ5i+ZKup6AhxPRHL02LncKy/VKM
idD24kkg9VAoR8O/VpSathqjT7GGDSQtNJs5jLSVpAogJkToQzIu4pkyH7PYd4dz
8Enn0ViQsJP4sg8U6QznR6BC+J7gzUgcVO5qcELRHVFvdCurBsXgWvUk4Lk0O67G
RKuNxX6etsoTYIZkENQEoTzxEFa+dG+MplxOCG94Lgio75vDiMww7HSh5ymOZfP1
Q120EJ0gC9CBSgzxgIEVdoz7Mvkven6pdZmb8WpCRvynFcirpkCnikSnSeR9nIHf
H0LfFvQmVCj9ed+IHcvGKjk/uHDf2Po/C/Bii1LqI7LZOeMPZL/GrNlFDQIFGs0d
HLHgDgmMMXSFSEHcgs5FyENub98VLj6m8a7MYSvKPmU3y0B2MqBCK9cb6bzij7Ty
IZTpAP7bgVkRruXYB5jj/h9MPq0g2bbwK3/4hYyFqPV1ZzngtLb6BYLlFX0qViuW
EY0pxkz/oe03pd2wsPhu2ub1WKsYV1F5VyLnRhPxobrW3uIe1V1DNS3Bm/afRMPR
bph0Fb5apva0BRq1jiaS5UBv5ZyDdc0ZfzsQj8TcHEHCjcJqM8e8i8qv+64nYNr/
vV+aBBcDyUV0hKe59VbtQHU1IFWUYLPg+9R5DaVWtxxIX+n8AzWu8JrLsbTf3EsS
W+Y3XMPEG7ZHP2d6rHLVZPKUEuqcxjFW5uJ9MTh1XxjFZ4WwR2EugJP7w5c4mEsd
P+hR/w3VCfoSM4O4hYMzAtzDhn30nEMf+xda/Z9eJ7bls50DvwmVVuhByChrpj2/
QQspBRAlL0hXTXNhQYAURI4gyzVYDEr3W3sQVh97ChQ+k7r1xvuZz0YOJVSGanyr
ahW+yJut+vtyKA5ofy9wyaC4DPocQLBbQ7G+NZRGMtXFLubbH3nKgD8LdMSy256h
JQB9Om0OrNjg5jcFH8VatuAF2cJ8Lgo7aG2Riw6G4t/C5kXrJR+ZJx3UWrUsGAoE
3ggg+yQwiv0ICDDXF3NrKKObIokxhJajRlIeZ8/yvfQNAopA9gpUB3hTydx15/nt
NcW20ZpcFlKOkmvQCST36wj5gojySc/qrdH0FffLiCRsWoevi09JS70yNlr+7tFB
oYC7EucD5T0/1yb1gJq7rcdelLpj25aqHIenOhZgN+kEiD34XcbpctTt07ggNmI6
sRk+Drz7g9ynRg1myFeUGCJTsENkiRJn/hvBDsiF34k7EZewK4TVZk5tYpCO6S0k
T+lod1Z0du1xCBKMGfutNCwI2B+PlXYLM7YKgUOX5HBEk9uNS1+ZDFcOFhvJ+UH7
cbH5hq0d3aK2wVgv9i6pgtqQNGeLTP8NoFkkUJQpcnE4GVJSmtzfRd8lPsLlXyAl
q/T2JxPye4ZLdi7ctxxhKiSjWbRqz5LzyiFqHr4wGe0OQO9bi41XMAzoA0pooLVj
jApfuhf8ECEIaScXQgnwj0+OF6mX4nIL+NGBpnC+AfAGBhlA5ivm8/3Z+oAAb+M7
4tjZbAEyLPw/GHYyoK+wSTox2Yj6gu9/agY8EqWVYldDQK4hFmP6K9pij0rrxoux
MhM02Orf/EJti3mXgtODjHsQ6d73GQLkTIArkvf7RcbMG6NHE0qksN/EIdvJiHgf
Nd5dbUDqBQN+smP6ktjL8nwJl60wv3TtUN9Gqvs8oSi7+kCG/gt1LV+RpKgsCy1I
E+VawN4aCNnlIYpP9xaYFpmeh4CGEQTR43atotQx1NpqNjPJtBEWhnvkWOJNRNeL
c7NRZDVOERR62oXTK8HISRpKFNLo+X2D1H2HReRVhhEgoZy2MTFsVWBvw2M3TS+f
awzDP/E6RArKVMZjip+IsZ+ewO35F7xD8EtXg1bjU1uE66aGr1hann6wyi/EV4Ns
ERWuFxlQA+8+qZeMwzeqoMTuD3PCedQ0EEZB+X/jDnKTHbMSN9EtfCJppXQWfxdq
VlRdZuqD8bEWEr8SKr+aIW5sweTzJ8wudzalDKkCrhQIwY7NhgYxOyBzke+mhfi+
U8zibqhwLpHYcZ32hUfHJv1OQQDASvYiNXkfQhyjhgMNk8J98PRlwMY96SIg3ykS
Bqxt3HQ6BQhgk+F6P9I+FM4viovka3hN1tteGOy7xxB2UF9eCLC3ARMd6OLzqrVu
0Po3MdgtqQ21Zctl3jYGtJgDz/x3qA+JjAX0M2Rj0nM5KL8D+D4sa3/S5iLglFzK
lHm7Kr/BpJeYExpD50ibIZShSlFdhkpOCvhpMHe9RLNXPKqeq15W+leDMbf2vSah
+Oa9url3q2W8vcgw5M0QkD7gCRxlS6WQMvEl989zBPj4mEGJAhV0xcvjjIZkb3I9
h6jB2wvFDrZtpPfdGGWMCVbO/ovTDD1ACQOKPxPhZ9MuxQUgeMxb03Sjnce8c3LY
ouUYFuGC3SxlcF9pbq5jwaTPL6HYphkmcmjGzqIFcCELbpWBqknmdUWdxPeXlK1q
MtGNkM+Z84WxUxzy1vpdLivbjXZHFmmPV40wfMTnntfMmSMapEPBH0KfdhBfsWGI
TJr6qd02MZMc1WzGjjFy7mMsHE79pi+8/AXDGT9haWZQL3y7SMIf0Ms5s+E0uRwO
vKCEx0XKY1BcPm3OXv9+R54e2xqS2qmY4R44umAfEDjRFg+HvYKspbyYcY2Op6u9
mUyZ/RgIRmvreJFaUFu4KeHuv2SgAUr6FFbS75Lud05+FTAh0bxyl9zQBHN4ShFa
DymI8fXsREKPtbw9uI1Bf5fs/odZzFU56IkCIKl5yguXH6DX7zqUeiLULpBBNWdK
RcH8wmxH9aBJDh1oAhJAo2oOvo1W1GSdqnDllq+qosOwOYcepuI+rB1ppAh8Edf+
nzA7CautCTCuqwSFybiVyVogjDOPLyMoNpI3jqIMoUi3OZaKdx0U+qNIZEeRYJiR
g43lSpIhaLu4UmUuuoo8Vggp1vnQIboFnnyvTgkKMgdNi2nzqnXQC3AAzALzslBF
9Bj+2ZjnqN/MoHp1vrOKSmPDiI1zZ9bgfY7Vr/bu2Q+jIxqg4IhmtUicOr0z89qW
sgVJEZsGE6gXWI4wzO4gJGTeNHYw12OmJSvmyWUIW8VgP8J9Lv7Hrys/FHWw2dP7
tQ1YBWMbsF/TX6RoGVW4jWIMTs0chA+Hpdm+edL75JyT3FN9qUT5BzjAWlHh2wE1
HSf89u6JYslbPSQUcwvJg0YjZsjJQIWpFEhU/nZHbxSx1f0vzq081N+nwGLB+JyV
FpxuRU2melHejqonyBNM2Zgz3oq1zyoJz9y3M+sAjqA2fpLRKVbapxkFuws0VDpr
qfsmEtgiDH8ZBmkL1QS/z8EjZnGmFgjoG8fLoF7Gre32vybm/uS2iolyX3sJAc/Z
CjHZyB44NiDuFfnn4k1uUfNgcF4N7jyCmCmk/HK2r+RVAw2Rhk9I9WOpitYm4nhl
1OFqNYdVzxVISZBfe+uFdNugwr28QbwsFyaIXi8ErlqWm0T+y+Kx5WleHbX77nO7
dNmFsnMNaG1i3qFJGC2I2+bcr/n8CYvrbDgweqzUBRHO+ZYoMn5/KglXUH5Ig02W
ggMx9XrtlOFOEKlHTkKBwmm8WRlM0JlLgv+afGO/DVTtmOuQhSzrHwbHN4d9dtlU
qj1A10gkIy6v0WQ+r2m5sThgFh5ohDwC/XNjoK+V20awAeAMaDanh8aRncJ9vSAk
syOXjeUdayYy/GOgUh4J7o4ghPZ7nTdjUQj4lwhC9pZx2auGzbVvsnGFIg97EbPJ
C1VWomRhWzsSZaT38KbzlDRccgF8X9pDUpKgpez4SWwUDP4z1GrmeIhjFtb5VreV
yJ4dP5V1XTJFwXfZDUo9O1/W1fCv/LZRY3mF+9xjV/5+yaDnks7Eqi7NFac26YhH
2GXHk1zhiEwdAHp6YKk+NagoaPBPkeESWPAUooJanGMSQGnFWtNh2GvjKGwsSOYt
OSxnFEIBWMkvaQFQc2NF88KwN8AV7uhgQ+tzhHXX2UhS/6Eokl4QhEJS+Aydt5/e
pqyj2+m7KJlw6oxTRXiwKeZjx8MiyeJ+ar0F21pa/peSTbPDvTdjqghJ1R+1Wd1M
yZbMvaGoPSTWOPihsQUsTG7MDrKVKrhBlMZ5XC+rYOB30Sh9LHuCUcQQzEg11B/p
DsSVCL2lpqALW8+HS1ncKJ70liCsMD3PnqHUq/xCGu1HvRkb1UzS3ZJJZkTKME9S
qpBvfeAcNWHiyPCQIs7cYihFrANLWWHkjCPOVwMcN/ZwIUvfdQJW5Uh0FShnp+Ed
dVFVm0MioXA3YONFKhwaK/gc5pF6d2/q1jJaJC31JF07aujP1yXO6/q8/ri6cfAx
Gzgv3pD3H45k7MNXh8H91KPIXKFRGXcwP0OvhrEuviBCUddOT1/zaVdZTKCIixRZ
DZ1OfS3rr+twF14xVY4mS0VFHvCvTnPb4ufJWJ/mDsrObWRJ/sMB81dt5xERTmt4
l66Kdi4gHUb+nR/qfPnQfejjoGVdNqHjgkzNmIrkdg/XdNjqFxNF3ftQksCvtBBG
jz8S1S594yIXdTUTuQHOBFF22vfpwazeiqkS9z37bNrVPcF4NzcDa2kPxJxrVTc0
Zyz1XwQzq7vrtN7bHXRhuXH2kGOzzQnIkxtBmVW//Mj2rlLs4eQwVfmjMU7tkrYF
tKLEyVRpDXJ1TgCkKTW60OvFXmKBN6xAVjOn/pCSPImoq6CU6PHIUK0/4DFiR6Gn
HUgiCMQDTeR9Z3hFU3kyw4diesW08LNvqOWQf9F9rVrSDdgSoz5aacs8sG3clIHJ
laZs8QYAbaqewtnJDQE1jmELsCF5U6/lNuqd0+IHKCn9pNt53/GNF+gnol+6ewKF
r4+NACDUD7zYfaE5+V2tjHga3SPoORPN2yDdrdmtVKH25gHJgV9otKmw96yy+qnw
Rk8kNBd5VuiCaB8FR3XxXX+UgyKMZfRs+8sESY8lTIM+ACXg1Z1SaPFNzMqDwk17
NUl3Lokst0b+p63IeBLkvakMox8wOOZshemKzNoHXKngJR9vFsZ1yDs0ukD5Zqhj
y6Qwpfh9++2mzxoc4CMBtDaeyikv2zyVRrBEMjbllK1yqjl36QTeEepEaOtpsu1y
HAR6Wuj3iS63pQDx0NB8YrC1qkHy147JN4zvdCKanfAg2yCs7E3PZXntwHmoEmU0
l1EPHoLKshfzlJnk5AmyjdXVbDYf8FAOGAxGhuLUEtWBGf1SuQwPHevEdajHDXsA
egGpCBnYG9+Dr2wu3pqfG/Zuo1zU+oF2dyaXnvwfDj53rz6VxtmUh2b/ch1ZKixa
vJW6xTtr5Rm4scNZl5gRZ52g3jOKhPwHYx/Du/NcTMbblk0BWWp0fG4ktDANAPGu
tX5sdpgloG5DYpqHnjkhKMKHi7MoMElB+CrvWjA4WfLl5P6kqVgJgZdU6yFDgkZN
Z31C3p+Nur+2MOE9SAKECH9shPl4Xns11IiNA8uCNGmgP9NIwbiOBKst7qF16Zx6
gW9nCK7wAVHVo514rdeO0el3a4izhW7alCuT7s6tGL+ox2ohuYpiLhpSJowzj0/2
reh2c3LQFPXMw+ylfthKR8OXGVuVsmuSGq/ZCtrpAlEvqUKlbHZPtMzXhJXhu4iI
h4LDevRu4SC3pAM+71x84AsT0CIZ/CFN57Nq1PQZ4h2fi1J88WoWm8XG9Xeookr3
fQ1SYo8/u+VkiuJTuZxb0mpo9ZuuhfKRxlP17FyF53TXBVvqFE31ylGrgAQ0yO3i
qvt3Yc9p8Jhof+1psokghfdpTtG8sMsMh1plLyXVzvSBhuGBhSfarh0kBvSXeg8R
I3Xq89CnVq/OkNDlBqqHKP0vtJpiJnFTH+kSRV0GOPrMWJbnxZG8i7DIHGiACLMn
94ujwH+5ZYMyT4pKFbPBYbMgI58KcqomODnoHZsC5W3zl2ATcUPY1mfZzxODupYI
6iVebZHObaIVEA78Jvgaf71fe0cemevjsNkERJVV6lWvzUkMduEhoWYywTr6k5Z9
IZk7BmHmrMbrIGCbVKqnk35YEvfJN0YAesuuXqD+nJMgOLdtwtsD0a8vUct82/F3
Yd++uP6wp1oYU98vfBbgq1HAPdJNQ5CoA4Tm3wnON7VWKfSTSOOFAS4S/RnXna3V
ta6o6MtcTSEpjPQ0cNZTv54ReO5DDk3MpA7hCNozBLa9wz0pZFWkfXcJUZWcsMMQ
sdw/NQCgntNpZBskQTtAX7AfiSo6bCd/MOj0+akAHxT8z+/DPS7abGl0wvrHL0FU
u2UsY0x12+ZycFGhu9BTgJd81lPOLJ1f73yCXHg2QzdDJwk5Xl1kWqQ+AWY5Gl9U
9P3xw8vURWOnP8qDrvp/pgqHR5VSXfdSNukGoD7T/WQdWTyoKETq3nrdEtQqkHrZ
CTM+If7oObC9Z52ncynzonESSHNs1Ya7/YDb6vjJAFHlD7RELBZhe2b0dUlI0/j9
EB/L9Pco/9w2NrnNab4ZZ8uEVaRV4XCWY7LJXJo9e3qUqB7INc4jiYGmIF0plaUa
sOBzFZ8+X6YFRxAZ+lQAmYekd4XcZYRw/Dz4VXH+6dwoL3O8N72YXkLVXbqx+IM2
VroIQe5VF/8u87GlWp/uD0t3XT2JwByTFUe8Ig2N6R4MC9MfKbdrkDwOf2ncSEJC
vHeN4wfhke1awQ2pKGo5sKd4l5WcLvy/WVzxZbpQsnKWuC/bBj8AeaZEbgdu/UFG
Nvo1Hr6KB+NF+BgeEIpwRAPGjSgeAMm6izOq6aKlBXkZ2xtXQaeiTW1XNJzKfkPR
IWaM++2KCa1i5TmRi5FXwdNdZbZWnALUUKug7hH7fT+r6blBuL60lHYMwUSGLWp7
nbKqpDv3KhkJa7G9lFZ1v1YVvJs+FIce0DG7AMYFdxHvQyQ/ehyo03kK/cT0St9i
eCZL8yVA5qNZg5JSDI3zcNjTZuGU+Uinko6AZUwvLf/tgcLSkhHOLiYkemAcL6+r
k7IVDazJZxG14Ahr4xW4QVhTUvcbT6fe+XLJPtZo8LRe3M5izG1zeD1Wyy2fG8m9
oqDEY5zqPtedJ8F3d6YEYEmjvVkm7L2TAXCTAXJTFWol4ZBD7bdKZOq81jpk4Phb
2fqrh1Q7pDJNWE3VW+R54VuPcd7msFe8yh+MWkEk1SMoWlDimAFZoustHNpAZ/Av
i/cHwzw1igvyqIdLbOLjoWraRbl3MxbpVaQnc10f4GbOvrQ2OtwrEZC7OYYf17II
Cl5+EoFgcr06oZ4OmUm2S025MWI+NC6u5KQsvRInJYNIir98rLsiTduoTgZnNXVr
JwCD2uTZHnD2UQjDG5WXzeuU/PT3f+D8VO3Qkxm3W75lZojOU2dQNEFgJXVbUbyq
e0bCFhXgH+dV7/9vaTaaNwyc3TajdFCD29JqKPKfs41LJZ4De0cMyoKW5bbUUO4q
etNF6sO6ob0SUihiKNzMUHqkpobS/dZNIQaGH4OBhz23FyzOGgp9DgPZDJncS/jI
akWtmOAGSVGRwZzMcz7+0xve9HcVGt8fWRwTeNTbAIPidPjXJOHuUkXhBhHeJiyT
1RWR+94jsNgTraa08ftS/Nrco1zOnvbCt8Mvq9Bd4YwKGD9RMSFAhOThVcmMr6Vv
30nZt8hQAG8za8src/mz7iwKWmk+5toYHoQJpnjty/u0CzlL5mV7uY4oAabq0YR0
G3CihXYflShuYDHDnhOxlFtj5/zlJWQFyPG6I+K4MCdh//GSvzSwmq5IaghXkGe4
gzd9Mmu94f9coV00VVsCDKsHGQHlK+7Fy1grFAF+bPSkUpQLqNwC7VKDQsYz/6at
k/gx2k/+kYb+gdZMXoJShuB0beO782AZebDS0f8fXSUj62BbJuyotn2W5KTxsy1f
P7KOAxUaSysEWjPXK0dZB40fzTASX4zf3HH4NbVU1XITW3rTjC4M2TWJvwrbj+yM
ZqZAG0SbTOT3PllZfoBzUIKAYnANdn+tRhA9OnOWPcl7sxJHGN7gZPKmlgkL46lG
+ai7LD/PQp99nvZ2jPDT9SEh3PaASW6TD3j1cC8FLzMwWE/0+weAhmnoQvGpDfde
ST7PTZ7I33vApxraVD+OWYS1OyuCrwYpLu9vRP24vvNfYD6kpspM0javcQK+SAyx
MAfXFgi5OquwYVSlZv1Tns/SBflrw9xjak4C5kLd86m4AyXLpkLeB5+DfrLTjFwl
C1r5Du0hvhhComlyx5qwMGRfK6ILu7IuyYlrc/YTijAAVI3J1MTXBV65v5cOl1Ac
6yFCDaKQQBPfjHaFJ+ZY7haZR8PIfpg4Oe6XV5Q1fhiReL6FMyrVMUrcIpQbYIZA
Jzjq7R5rhhd+Av6QCRDIXK3gJQbD7IpKRy1tv4Xgd9HTBGIn9lZAuvvvNSIrEmgW
ld0kDKksfbQe5yBxikUsLI1be3M+AONKXW3M56F9JX8285XIeZcj0+sA0MCN/cfk
cH0Na88b/OlAWV2OxFKL53LnNODPPdsAvMUCVTP8CqqrajoQzGk9WOxmvOv7TKm1
U8UE9ayLJU/tf1Qurfs+74SCh5iljeLkVX/pSiPIuArWybVtWFASqJrJ4Fi8jLSq
YMbkVYsNODecA9qUFLvCyqKyF8otzK8/qz+GJyzkWQUI2PsJdPZyFuc/cn7hS31W
K0Ov1V0gFQmtL2BzZdupIut+oCPnA2KvajGW1Inztc+Xik4S4t7LRskQf+qRyxFL
WW35FXvvl/EFd+HaoUPyw0O80y4Y2D7cXXosReDt/4SxXwnXb6ZwlZ9mW/TPGIIN
8gLqEEnPVczklNgkg2jm93TMpMdlxlr4x/utvjX+IDnA6s8+aSYrEi94cY+Fu+LU
kw4VIBreaTLhMD/HKtLJcq7sNydQWfd6dlJcaaAWhX2liX2XniFKkGUzA5LU0euj
4unfxyNoG+l60i+JH3fd2QOX68kj87lZrE53lhY6qabmpWrFK2teVuiCXalK8kka
K8/LC6JUj0qAMJIVk77TdqzFWwQVXU7fyGECYheUpZkfDZx8vUg+XS6VvFdth7X4
pJ6UlI01TBdcYhZzKFbMVj6VH0fa399vTWKPZgx7K6iZRGfVMVkrURcUyUZ2aS5W
lt2CTFf56nUsvwjscKzv7v8fvsvzh4Jff6jcYNfgi7yNr1dHzuEYXo4kiBrsBcGS
jMA47QlXz2JgL1YGgw/K9gAlis5TdsHLzVHbn+EPi8m2Fhe2Pf1gVd6KpdL+lrv+
VCHWrtxRrp+/pcTmx801LJuypHXadU77UTV/7NybmtSrqsH5yTV1njKiHn0wh0Cr
YT61vbEVxbtF9luavz5BJuE6ej/SgIaXuR5pzn/UEoeEwW1U0vHACaPZIY1bmLqu
tdBXIwkVHvHWrlUPg2wW+51rs2c6o5f2xuSCeCui7WpG0wC7xHr84ppd+Vi5tLky
a00cCf/sYaCuM5wSwXC07pWEkVOIXotrSGa9Mg1ux/rQZ69epbsYHBWiCCg63AJh
ASGn2kok+FsEoK2orG9wrOrnxFwVOIFbJUhWv1ZM+Tdpa80KwFsqGdqb2Kif20Sx
lRYD5cRRc2dlfxEFD7cxdT0liVd9i3neQ8C/JmY+F0B/mxSL7L3FOFLhd3c7EQgn
ooZmzPAcXizlldTiZoMlYHcePazb1cBe+AGOegHUk4T17JXwjKCZ583tkgyykpZL
TDmUtT6emouKms1ENk91MoVzb4L1iULmaa9KcvO7N9ZUqbCy+h22XSW0YkpqPN5F
Yd6+X3dEADlyg+0dzkMfg7Wx2DnYW3eeRnkKOvhvrs0Y5RIpGP81kHutSM58J184
YL9SqdsP/qYEbhxNqYlAYj92ZDPwwW3eS0uT0JtQJGMAflJ9y5tNzAocvfer5FU6
xx5AwBVX6YBjJkhEXl6iarKFKwzs5NurU0RobdP3hBpqXZ6qlukhSKkJZoh6IVkt
iZxmCTITjEF+9Ibn/Ihs0NfbUNqvyYCCt5Ah6wcd5w2Ibo+iNFiUHdU9KctOtGQD
8hB1sL4d4lwCknMi8HaWsRWlM+PP1HDXyyK8lrxcBeHmFRrZe6Y5gIi206BI08+W
L43ci2SNwufwVDib55Xyk8R91ffSCW8m8wMvr3IASV2o9qeGJqAwsCjDMAB57mxY
JIYsoP7ffoCLFUR38Q7CSn8SLykiSg/HBjurDQ1gpwqJlqqx0TwqTXgoWAJqELxH
SeOkI7PHBXQSipt7ozDClvq+Aas5exyd1T6Wci7/4Nfoz5k2+LHR9JH3nGqDYXF2
/A/w9Z3dJoVwMrL9RgjmF3MX2T+vHYpxFNcarW5oJmCkwy4swRNa/H3c3NZh4X7d
ypSkF2ukGNBeVKEuVxJLCXnlhaWx4xLusYZUpyOqwK+62rdwAuSqQcKGoOSv0csC
KBLG+li6VJYUcJKPJ3yQldrMoA5YlbmSRDpf4eBou0MJ3IK+TdE2GG1JqjMyjZNS
JO0qRcjeQzmGZeix3fKodVk/bBIf8BaHegGvkI2FraNdS5jRyG3QbxlmVuqJaIEq
VsHP/a+pknCbvF5iNf6sMVCeNYCWdsRCAMwtkaRqg2tNPmrscddQnb+3nNYFFR6F
0Uax/GwXgOb4wV6BYRArR5eIk81q5CUU5t3t7eshPSVWsRKWB84pLJVUi93svEiY
yI7I1Y0gLhVY787Q8yAxr9S1JyZVFUF6q3Z2IMfHF7Ar+peg3hRjN5y1XS2g77Ip
FG/DNRlJfNxGe07UXbFG8G89xzQI2KgHbWECC3PD/tsob16UVPWZDJRnmMHUaiIo
rmukQfWXKaCCIK6efHqqTO2LlIoYbRpmzttItjLnP5lutLs/YuWZh2ZfXxUOIZzU
3OU66p2o/E0/kZWyYv99eCI6/EPrMytVwhY4jk+gu2Bc6vbcUyMNmoPndEZfYhZO
ls9D50hghz07GptEtOYlIySt815d0B+NFsZln6DoG0lZX/pa2e1FL3jhgWoKFFzV
8mDhO/w85OCow79J0kNnSd4yHwtehuJF95oUfjH2RW//BMsyVkv175nphcQFwtfj
TmxBwha1DBMCEmnaWreTv7XS+stvREwK4vE87Y4/guOvsd+61EAi3A/k03oegg+e
HK6Pgl2H4oquwAa/9xg8F+K6zf1RBS/15bkwyexLSj6mDrl/aGC2elQ17/yUPmbR
yM7ctTZLqdWAEcRwCSkr+1KetpFs1n9Mh1Tois1Dc/qqFhQFyq3tjfOnYQ4R9L+o
HrwqXdAdiBRu/sHg27QNEfaOVJaw9rrogAQ10hVHbCtBS98Tn9rYjb1Nhc+5KK/A
d29TNnX0JBSUNKRVzpEVd7STa16nwpQGzjKrjXboRFF3fnVP1IcIy5f3VZp/Ml46
8hDRE46OinElbZkorPrs139WnsRZ6N5HrA4fg71bu3IABdw/JhysEpqC/rkYGxJ9
o/Y9KJ5qQ6f5or7AFzjD51vClIEgiL1l08xB5oPpZTGwov3U3v23ISf6HhVgvLNE
IjR4WSqQ1ZjOyTxPuQdZtirum1d2Jf8+fpbCmaR9pHImjBlCPqecGJDfVnSq+bhU
F0Z8s4oxEM8axaet/CdqsfbaS2y5zfK0tOclgoikJqLYKTYDFk5gNKe6jMGLjHCB
brknvRIcoJVopZEjR78yzkw+besK9Uf8LSgKFpsZXSXoo3wMTeIr7rHs5BrOH+Ns
jHoryqIJoEGQJee41lBNnrJEARSuNkcDfsZ+48hinUEP36pyV7DJZRsSeS+gSSNH
NfnacIoe00/sCasXouVn2yYF9Bzf+XTMK3rCD8EQAX81VYLMxIDwGCN8XDE+WASI
TR/JSD8koqErTphvrdFuD1tCLPGHQcrbzL4x8KQS/6W1svqQp56OJJX8slWj4a2V
xw+70fme8ia56S4JIslOlvwR3FoKewrC+taWFmkKq+xFOPVqK/3p9mxh7xA4xme2
/2JzPeiUmSlNVti2HUn/qOAjoFE/d+/8e+/kzLIy8+ni4xW+7ayZQFCYqFG/t2Am
EPFbtNBl/ORzulHgM/ai+E7elSvRcl/JWQnDlLLPu89uoD6ScXDbKWXZBfp2PjBN
ELRQdLij+2mgwHTI9Ia4uM6Dpu3nkpPlhDiojJ3icomx3puf9qoaH7/xdb/E4zEi
WKyZXrZFJuTv+yLy/b2qDxcYHYEtBAU2PwsK4I94QKjHs1Omu3vnSXajjKbuQ45q
DUDUo2zKQ+9KCYDlbI1CfI4TK3kKtHtZH55u/jhwblcn3Ba66TBcZHaN+yzcnDOi
3pMGgSdMNo99gZoPtCKckbVzD/TbcJBhf17bioZ2lLkvDgQhqJsMdypAHY0erXmn
v9NDg51zUgfIXs9H8OV/HRRA5LQD+grgVCieLtm401P1WYLuJ3MMQ78JxHIfeqXN
Y5ANVGPJQja32uCEI14IxFlnYlbL2c6vmfRBdcrFUUHzqpibq5fZhWubMdCsOWlF
Ec70Fy2Wy2aKAnsVVui/ipVR/3B3BtzfonJ+HAl+OGi88XNI966gfIb8huriq7L+
//n84x+tCNIGKoQ0nHOirXhrCptKYquFEdSGmNG3axKoX57nSlj0DcIZM7PZqIBX
paG+MpOjKm4ryrDmQBqdp+T6kDrXHvH9gnhxgnUAUIKfi3Nd/CjiPx3DqjnDh/6h
nxv/He4IhBoFP/Nsm7LOhG4vFsJxeAYfX+2XNxcFQoYYy+KeY9Qg86mzjJfg+FDc
ko5EpE859WSW75LhQGJW7+OHwBXnlUAr/rUYl+lPGkHyWUfVpv4L0tNLgDaVPnhU
BameVbshK4qwxBHuNMYYA735PplaNbIAw885BmAycx6Zwimmjvd3Eh6towcGKSgK
ZQdHTRTA5h28NuSjYbmqIm6tPzcmQgpy9SB2ywExEGoT7AL9jhCU1iLbeOrm4Xj0
pALiTNKk0J7ZGPO316y09xD229NY8ouM//T4H/qSfE/1Ocb0Qeid+KloDEhF0S51
5wSy11UB0q32F9bzaqzO/7/Ab10NNCHmBnNKGrCWzTs4EM0md1LoAYkgKW0Gv18s
FmdOHeoa686pcAAlRdC8w9hqwECrkeY/HTEYyeC+735YcqrjkXcyTHIkRayVpu88
JBCpHs6BuYFuhUJI4X+90ofMUmf+oU/ykVSkx2qMo3pZ2dvUKPStIPtU2+TF0g4q
aFTMA+EYBLHASjItA8QOQ+HFgBaMHCMTD4wV0JjsY5iIPsbNGGLJrN74s/zIcc6d
PqkVKd3t6oB3hTjVb4Cq0jiT93m8o3nip0uQf3zIwhfC3NUMDwh5LRw8uWhp0K/C
Izjow49nvmuzLvPpN9rFUIQKw8tF/zAItIg33qmxPh1cEn+w08doKKuEKO3Zy0hL
ZBGHCE0aTGUU2EoXN8EtUz0TvrwKiOjI6sj+WKvxCaSQRLQjuOfEwbSiBwZea1te
BEK2DQ+2j7pwjmo3K02/QXPRtPUu22SCWfxO2VxM/hs97KSZBjLXx1RU53YlozIa
mWfaWXoV8c59hYcL5oyEqdjC7nWN2HM5wmA8Oohe+wtHFJopqA77zzi0ATzm4eso
VpCKRe1rtkcifQ6nQPure/y1T5Rm1Vi75i5EC3jYB1tjneIwVr+JIq+U0i6IQh4H
jp3Mk/AE0GsHUtkXEQxOF2tFhOU8khRcpuxCjIrIZ3JMl4Ym/l5H4+z3P/Wytn4l
pX0PA3D24J5OlzTjQgOesqki9Ty3Nwv78KGPJkocDLQdQwLix5kuaLxDmPyaTvbx
9mjmTaKfMmgZhGum6//EQp3oaZNu/mxW03OCs+F8OJ440pPCIU+AxtXG2JIXZtba
bETt+Zhn5V0imEs8bX/nxGmRzcpNsE+oT9hGtNauzT/ZeNgLQ+TgO2fYoMB0e9LZ
uXmgs6VGhDeEjEeS4FcUpzVal1zaPJEb3ac7fvpO3Ahy0bMNEs2mufYw5fPuzJhv
JMp4UQ9i2HDw6Pqyrke8tICtwkz8ex1S9qjYWgdW2fuQCo+B0A3+3d+siaADb0DK
supOdhJAp7/TcyQhLFFRtMaY6D+Nn0HI1A48vlGwyyYq3MuQ5/07NpQRNlfZwbxg
qEzp9Ws9R89TfVZppk5WfhviclaWzuGVOTjxWH71Llkxq/GkRr16i3uFvoxYP+Tp
+qjrx0SM9DkZnttxR8o7WxIoI23U0fVOHhI6qFKP+EhTLhTZsQ5V7zl2wBTAJkCb
MqPpQq8u41pYZwTLNgZwttsLZ1aIzus/avAWlVXxYcQJka1kvxEDv7Ezub8HqYKJ
Lk/ujeJyCOGNjDOpK6uaqHkvLVGgaD5namMz6l7Jpo+Pz5WLfb7vi+Xn1BYLrxJj
op1ZFKva3c52cjnZiEWTyMmWAaneMfRzMO0sL6Ihy2Mlahcq2Cbn9gRY2/imVj17
ORmPjXHqx2WsztX8wjmanbnYF4Qti/2nkYuAdwsCANa/euHPTvVF0mpTUYLHnHMA
nFl0WpIiXVeK11UbVzE6T07SqWR3u9/0GLcAzNqLVYxc1w1FEuU2W4WOoZ0BoI5X
LdPukhN4yyhlSj18qsg9IxCcB3RlMuECClJBvZ9ZAC4urYARPRnQydDt4prI9WFl
Qh0XXitMu3eu4CRGdR1N61itGFG1SoCpNmJQvxlIKf5cMte3Ux5PZnikJ5sKO6Fy
D7rgbdpRkme21JVXkNnPyS3e0TH4rGK/ifZg1AafFHp0SevFbuaU/S+x58038wWk
UNEAlz++ZzoaWMIcS8UcIi7J/eB7gdU8kLW+PK7ZXKU/d8DUObflLZJmpYrifip/
Fbt6aMGoLd7PWyvqSdRgoHKpYHMWIdPgaMkNRpPloSmQsSV7GrWBMRapRSdQVWcM
cAnHpVDSEpvm2mu9LDxqt/x7Q+NpJ+mSM8uKnShoJeQfNGcPnd8Pg5Wu2W5wTNKP
Jz2VB9wqQDk6VT7tg/numQWWhTr4P7Bm6KVZZJYiOQJpeHiBdWMkdiyyYyLbk/zj
kW68DsQTJ3rcj6JHWe3RLlY5DPbtRzJsK/L3mmcLhR0NhgiTD2QYs4Pwrl8rm4Dq
kNo/qcTP92OGzf6lT36R9Al/R7iO754Ia2c24xLeXvziMsJv2Iq2nddfFCQ8UNCz
19owKozBXEJ884eHSkoMmVZ2k6vdjRQnzE5THPSYB6G99QRlk/03WYv7O9mKxfD1
/kUB5gHUsTGotaZabiYGWuj04uPQnjf/On798NsZ7mropwNqNBK//fk/82EMIizQ
/TdlcPazqcM8eEyN9kFrIX494tA+uKdunjuDxoy54pw6xUToG4x6AefD9gc1KRq1
bBmZtZDp2aAQTdz/zuy10RyxzykccZudaY0Pz+GUd5ZJ2dY+0Mn6Zm7rJ89h5A6S
2HgVEXsAezUvJ1LgLSkpYsKCLPzL5d447chtFlN+WSD76E7P6KshQw1lw1pNLvcd
AirlCrfcMrmwfPusrLipdJD1wkhr8R/3E6iFTSgZ69LOzU1QRCOAaghV8PBBGgdE
AwdGvRoE6TyQg0ZO4SUsnwemqM+xdfpQP832m/l8U/D6nr+t+4NDf3/idd118yi6
OGaCMwGa+vML1Y++spPTC49sNJW6l0yqQtHuH7L8zuJfkkLzxaWxwZIJ4VMKPsto
7OpMkmqhpoEze8EwbIzXykkkW8hkcyd/OgRvl5BOLx6KeyI8o5kRjHpbCC2sUP0w
CPoZ0uIBaPLytfNKeSlzMAJ6dQvLNR/VZld90B6rhPdh+J7ctpZeHkp444oa0nGa
ucti/RhnpXji6cyr0kia0gKLw//7bdHQCVlDWz4YBFLpmACjzASlEet27PhSVz/n
YYSe/0+wMHymz8moQ0bnz8lIHWww0Pta8/dctXW2QfxmwwcjYfO8x9SYLMFFB5Y+
i25lfvgUU5TKvFt26cUx0uI00uljWCGRjthKM+3gD1Vg4Lm0d1ByurK9yVkkiTEe
3ZSwDOpDZD4gQqwavHhM+fM663UVwbSvLYO5Wj+cuxMDHU11UJaszvJL7CUDRTQm
2iuVI4vV/Lhk3fHfUSOeiv08xQB3Byw2LYv/BnZvrWX63J5p6A1gm/2/S/BaYV3G
et4Wsg/FTzTwLD9O8TtuRDyR68xd9kzW3JMNGMbAukX4UXKXWoT2WhCFqEIdBecK
z1hwkpQUaudsKiIBtVEO24ePA87JD1rpfcaRPCGF/3+88ssVpfyaD//hEw1e2qL7
VWfHIN4Gcegt5yC657gcosxcAuWJqgFhZnN/Agkf/z26EzKc4MgY7wVA+9ayEreJ
PSi3uWravaU0WB8Z9cjxoji4IeCAg5pOddfqim2+hSyuE3Eu2AWDuGg/jwVEHz8j
eMt+r4TKeWLCOFMhh6X4rfxTKtihT5MKhWQpQRFzn9aQgIWC4MwbVzUmMvaiac5P
1Huv7snyUJjQ7CaoV83g5mqDz5D5qSm+sO8HPhG58xIZ4EiS+x7L5Re0aExz5H/6
L225jfpp2+QX565B7bsezqdiTaDBYp/uL9wPVueT0qdA3sGGyqBY1xqebWnjWmXh
b5qgrG+btpY4BWxPkE6vZcFfimyJFSewymgvYsCwl5gefeqbMTporEGbT4yoJo2N
L2i30tp3MDa4KurhdT8IJZdUMNZ4IC0Ymuz9NQrh93YBSSnrjSnNM9zl9hO6Qp4g
3+rU74gRZncqUpiIloLFcFytcq2obTfz7yxDfdD0X8fG4D1WepRi0D8E9hb2XPQ+
2QLvSquwNXj8njhelQcR4bTLu6cVmyXyCb2w36vHWdzIIpP/t26oDQrKm3XQopmO
l6JGBxMaECPb7Eh/Rr8MzuDAzwoYosR9lAJRZxNbrPiOWaQTsBF16gGXQUIIqmc3
joIKd7nng+5otTrjNLv0GcjN2mjp4I51/lgmI3+OEPtMHGSIX/zDBWDh5kW0b67O
VFlXeknkKckwXUUgEnt/wWBsysMM/XrY48ipB4TezkOgUe1qiA6+nGuvseVGZxC8
elfNQJvo0ivZO1tH4DpHYHLSf+0DEy0ETK8htDKX/CaxU2fySXK6nk2RHAMdl633
zgeNbpdwqGaf4etoacR+kt+63SIXP8rA4J0lJFyzBL2nH1epYzM4UJVj1rcDeYNr
ts3ne2af9jY6GwJ1yHXguaG+scVwom5aMHZwBE7CLFxTgO4iSqd81fNjWQwT8WdY
eebhQm92/x65l6jjkvA0V0X7bH/QldJ0iDb1JfKtf7kivQb0/X6KAHjiSVmehNK0
Z99PCb1qR+x1XiKrifSPPt2Qx7kdEolt7B64RblcuX8J9Xejo5+pcQya0eWn0NL2
tRynfW1pl/+fMf24TWz1bqDOrc3T12kTKqqrHSAaqM3b2eM8lipnH91uyorHVVzn
WWjUpttCZDCowEqAM6XW114/qJxvJnKcnsAZ8cjgI1WjmFr0HpN3kXh+LgZvL9ZU
dKwG++eNUydJ8oxRWka1yql+7SwVuafyfU6NivB0gk00wyzIyWlOOv6MMfv2lq1O
hLuspUq1ozN0W1edZiWLWMqvJea2A9mfrbxkpb/YlV6BwzJgF1mlVfz88sqjEldQ
sAQ0f4KmiNj+VegJpZUuBfZBp7Kizfw7i96/V5XIVAtvK4tSeGbMZ7P5yUz7ZFlm
hD6MVAMx4hzD/WfTd/qfTXMT4MBm/Bzvie3hXP1aQLaW2dM6iEWf5jhpqEvVQr4h
CiF6aMLsLJNTV+YxgVcCTXcMmpwZBeOraZ/F9YTkrCoFkcjzHsbf7kwj0z7I8V+/
MZ+w3KQuKrSHqmf7zyRVUDRdMaebehPidBcapH8QMX1jwJn8iRbEd13tP+ivg+V6
TrAQ9QUQAv2eAqkTMY3nGVyeKXQbl3P9CiNyPNfG2eYaAGGmOsIWB7UHtOsrwdgg
2LlvypAhZf0QQIS2ome/7NZ2xtlHTL7QyHS4vFOA+VjY4MwEB2lF5ifmOMWxJ75Y
rwlJ6MuEUuB/Hl6ivaCsoUD0Y4qBkmHQbdQ8byruY0wjwQUmP9EVX4BUM4TnguDw
rxWiTA9LNnMDfWkbXWnrvu4yVyLhw9W7EArQEoyJpM7MMwytpuQKOTBCeNDsAPZq
/MuoQyWR1WyIJNVBlzcNZVq+kW27PDb0LdTspjtg3wvRwyf/zwEUVTQsdEntansZ
z6wf8p40sIY9QxvHzaGjgM+Zs2NV9l8tuSjZLRkdXeoxiu/YsAXIGHwCrDRjkdUg
Kyq+HEcpyKESZ2r2+OdksYHecHcbnDyxYRPic/fQQkRjyXrvB2EUmA8nYN1mfOsM
bS78AwrQUjPCdwoiiJVDXQjmg7E86bBe3upU7dc3mmjk8Buc+NUGd2fHanA+Tepp
6ENtmKO1q5c/wl4BrQQKso+cANpmFulDeN0ev6WFIKLseDfQb4XcmTb3LO571v3O
N7o+R2AJ/P8ifn8MUpc3IkCsdNs9BQxNEpTP6FEW5NG5xoVTjrfiUZHIAEGI93fD
fHrarhGUPj/5+Y+yOA+WObVJm0Occ86GXDsnaaoOmK5W05CXuwk+VjTdiIB45yMC
LrUb6Mvpce47j5ad0YCjG8g7tPGoxu+0Vci2qCQfif5/LD/lZZYkwTZF1DnkjorN
H4I1G96p/t9XRw3f89Lk2iTBwJJ/VxBrvrszgO+yVcVsboLGUZbdNnMlcnGFOv1D
ky8F2cpO2+CIDW97Oev+YcD3F7/qjF2Jg4bvRihjuxy7xYuGNGenSahmd3xUShs8
Hp6xgd8LdpoLgce/waLriz+OAUEs1aBm89CqZiolepRbmMWcVpybjSpob2HvRd9l
t38uKf855fCM53Un/n2YLVnpfRhuFJQRWhwDjXqGH/g3URKAmcKSd0uEqGjDUD/V
7/LqhO8DUIDLbSc2Ny0WrJItxyJV2XN8Rc2Uvoy0oyfAZOjkNJsr8J5AeURLnKmJ
1ia80ak7t3YT0B5OP+OGdpjuozNYlEdvw6lOFOJz7alVbnfl2lLiGcDXW5Zq7yVe
DaEby6u+J21LwFPgPsipyMRUX//FvSvAIjcmewNPpxaccBbNBthIykJ7dkCvlFlk
B2kooKM60GtNf9BJqzt8Z77kglHo+20ZeYiT3JxhrlqsTXt+IUMi7+E78nJ1r/nA
mDaTzV7C+TNhpdNiCXy5yIx19NPWD3jY4fD4P8KFvXdpukOF/kjtthcf3jGuAt2X
xIo401txwepk5RnVQXLr0GU6Tj2mRkYiDZykbXgUOqyBHxLeVQHrvypyFhWnxChT
UiD/CAo8pOUvjrlRDFN3vJDP7rje145KTjoilePm7K5e3eqcGMs7PJhA6rGE20FQ
UDGiGT1jR83nzXkRy33H+D0x2Sa5lz8tAXHwss+93IWFddqGmkUHscausPYdzKxZ
PNEV7IjjHGCMunKbeUCsDrdcYO3DLMwZKaDA5gkzHs98rrvItq54P3g/Vfw08SLv
wW69PgaxhEWusDrWtONCUalT8hz6xH2RHulGa9l0afR4Z4TbQxMgb4Y/FMegD5on
ovAu/Z8icndbKKJCGt6VtUssfYV7VmUZofBBb4akPSRHQv7iZ14Im3TP2vtvsh5L
HDAoAY+/5JVGCPQkh03VoBdPkDMKC2XbS3XmqY15ns/5gJsBAx0wUERomBw7rJQd
WUPuTNHxbkOAZykuRIoqRwNA9fqmL/adEwIf47AAJiD2RRMUmBD8+KTC48Ft4V0r
aZ98x103MLTTNKD9Yxm2lKyk2U9fqR3t3YZ2GJvfNjfzidH57fxth0wUAsWR7Nnw
APW6DhtQ53NkmeCmlBIjsK0cNQTS4Wx0RAeZ8Yza28Oa4zEzCIsqDneFvUYlHA1v
ey0WetK9F4QpfHHXYBsIE+HePE6vy9SOC7AunTKjdowfYLeCZYLZH/NHzcv4ZFkC
ykP/wfbNBZCb1vlad7CjmrB8IHsGrYo+XRMjLcmiqKNvTxOWdS3/KrLmTYCJnmxh
lp8BWsufAG6ZYUfP6xdUOy6Rz3kBFI0U/UYS0NoP42Sw9/z2VgrKHJaHoA1PveeV
Rg2Hm++5wtb47zkjr1Mlr1AYWu0UCIN7MJzwzPO5ibLYmjpwVC4UV2H8h2QVE/xm
t7AZ1hPFp2QEKaVtgM0IZCwud5P66jyid8tcfKohHvdUPx1ddYz1atBl2YzpxXTm
yp7DzUhkdwbHqmdh52uUUrOAnjYLkPfvxtOaaVYDMXGodoAG3WnX8Mfn0qRLgoUN
2ukU0QY7vhZzq9XtVfDh11NP4pGlDdxTPTNRz1NOombtH0PdwVKX7VOwwy49QC0Y
GY7NMEdqumZCyroMnPvg8J11YKDzWejdkazkNBableJ0D4AkBa0wWPpBXG9yGQ4s
QwQkhDVCAZA+Su/FvQhl9GXhbV4x80ofZN6Wxn1IcfZ9RKJMboX2RMKEE9T4LpNc
NrOaQOmp+uFXMCszjnzLSRfiYsSeb7AhE5RDe6r+m5IU8wFKJLJmVgndk9rVw13K
uzui7neqvYBJGuNpyQ6ra6c99CLzOtsObjMfx1pwkauEk8pRYyQ4SR88znJNdZv2
3JTfinF9MBTh6Byfj0VwHDDMKHiSlhGsMDxrpdnl1h4kh9dMT9Tm3MLnBKNbDds+
5erK1NHotGvdyOOQLi0HO9+0UZ4AUG+Nysrbq51HyMbYUWhYv3aeUYjPfQXhvcyV
JM2GFm6H8NZyqXoHQ4ELB6xhZz0VXSDHYY4oZY3ptQYG6AAGFVdLX1T40HhbcEmc
kUq++0uLw6B9OsgX3KNuaYFX6kuo+jPQaqpwMAwxboTofXqueqEQvp6cUkyOyoBu
1jbvfUBhwM1yhLWWJ95Q8JVFYlz22GWnrizeeDjL+tCg2A8o4Z2yAHre5791qy5k
Wl17uyL+rPai+j1VfJ5bUQdOXiS8C76OaV+KizFPgGM/M3NNlr8e+OJLbCaFeyDB
zMrYndXswbnL8xsziGuahq85euLEkzVOLBo0ZQcyBtmuVpeyUMQVxq+VIJNwmKei
G4wLhH1rpHmWAUReRfHgQlKAqTvsR6EeoAfceUHuCtaQ63d5R+YeN3BmGHYv/uAr
nB9Wqv7GwOOjIFjvKm1STmjy3sugV5TBQ3iT23FXLeETsLcRrjfOOxNOu4SEiM+2
kn+arRqcvsk+T80r+0YxmHFh/ncbFsu65ucjQ1gXQoQlQvolq3pvkSLc55e6Xeh+
KtD2pAwCZtT3N5n0wMaL33OdrBoDuU6v6bdMkN/qQKG6li9TIpWzm67BfXYEbFtI
M08s2ezNpY3jnUcJgZXWGnHhmUl2XrhCksvHv0DB5QgSihCN3j0QcuNBJ/wQLLfX
bOdpfr9NMzBiCeljJ2lWcR9y3SrTXgppQyTKiPgusKb4IV09SiOHve3190zmylVK
fUFu4dNgKr8PxmTL3KSDknSvNTkeEjWBjxBaVy0IvwGR0OiDSCLdWXrJVksLYnB0
4LLwET1MNzomKxTNk2fW67Er5PRpiubprZcnnuVOKeX2lPjLQgMfzOPQQfo3UcTp
tLap+HC+GZ9+O0UniTcN2rprANv1Y+96YUe1/AX995OK1JcOUBfhR0xbEKiE4SAX
hVebo+JmX7MTasUkupaZQv6mbGfdhkdgalG8XZx7TGCuuKI7qkhPDLhysuZmuusj
R+bE1hkIVTq5vUd0skv59WsghuhWWmzRfGTzvvUwXkLtrP3Ie11mPv2dGPLdlEMj
AKGRChAxZEwcuLgFoy5RrL0nt9chwNOqhuLtW5DINfEwL+LgVoMcjLbtcTTMPkoQ
XgE3NCDdtVK05eq1lGhNsuIY7yWJUgg6b8tCj8Qk4HXatn7UchGi19I0Qt1UnNWK
JGZzdRdDljN7Gq43wYMeOehCLCU2YIYrgB6XmxM+VchDWT6YHAlEoMihW13keg6m
oGlKuHStttGik3RKQKU3r/PLIypRDaKlSC4dRK7sIUemBYZp6V7mfr2OxRPNZMSu
qVlDolXdKQRGTfW5OwoWfeT/7S9EcoC1aQOQozG72Tzv38+9/4ZfOcdjskK+MG3S
+5GmgQqDsSuEOD4qY/ouX03sIYlPEiFNAuoG7mPCAy8b48AVWGqFLWlBgxNEilii
fjTh9YPByJo9kzm6g6VzmctF4aFODodGFsMUm8oEPLRF4hX3kJd4Z8k21IhjxEdZ
XHpkBeDHsu0BiJ8aj0kibZ/c6plfC2O27wMTHXGPJS3HmDu1tQiLvgiRFZBj2WNg
rTWXG4/xWkJVbxQ+DP02/BQm81PbE+f42fpGgxJ/n5hJouqL0An2y1MSjoZWoMGv
PaDTRhw9zwnlFtG/BL6cboivbzXgIhwYxLIsGE1Nt8TZTBwOgh5dRLccLzN5HTQT
I8gCd3yO7JuTExYradX3ZfMn7m31ZSbi+FdWUFQ5Mb9DPDny6pX4v22jv+WDCBfM
U05rejmAz6JFMrrVU42mfmuBEG92hBLz0bR6rXfYqbNXVUyxFXTnHUz10JmUS0Ad
VJpRzBL4P9LIVvnKt443LJFsLRSMnjWPg/SbrEPpqRc6/kA/FfuevZafMlWEisxT
qIH0ab6SW8OtEzKiuQz0ZcMNOXeEe77WmLsa8FeOxAu1uznVxDfIK+sEALxHJyGN
GrtfJQSs7jxqhwGByryLZUE3VIKb4gp3HFaxfEX5QlDGUcf1dh6/oo4CuJxBTB0q
YLdr8Y37juZwqrHODBlbqioF4mFAZ/og4RaJWtU4snu9VzT4/m6vnPTx3omfd5tR
R9GP6RDkP8HEZXueWYFeFNLpKua/UlZA9FRgcXyiPGjcN58V0DT9ZM54lt6g73j9
v4UOibdeDIT5OkyOwkLcCFFC0JJrDb3rr4svRFJwChl4q2qB8hmX9g90N0pGOfdm
+pi6JmtXQ4V7IrvlqtH+ooFgh9+gFe1ROrN4NMRYCw6hGNlPpWZixPDKRLY0UID3
oL7fOOR+nOF8v834HZjfGMokE9VTc0LhnRlzT+FJQmHJXFgLsO7xWaH8q7QuN+Ic
l+EvKjEdcUUipQrjQQRh5KbMyO1D6m+ctqvl+y/zvVbqqo6sUIVpaVvjSLJC21Ln
IEXQ01vHr/K4z19KIMfTOl6/b7bA+2EWmw6J7I7hRtDeT6B8Efg+0d6P3V2Enbot
QY2s5v8c83ceUCA3YTPXhhj2Hd5dw69ZZJDf+ojepbGWw+FdPYlzeQabPDVIUOm1
uY0N3M93mbCiR70DuNLc7AZpc/SN8VMCvbN9PgVjIPgqkdSKko9YmSnkcTycv7Dh
qopJPBwKnOSKAPJDbCL0M3xSTdl3k47ak5Pwp3b9ZLf5HV6lK9Mr88gXWZ3I0dBL
MDeolDeyptP/TVHKmLvmWONPrqydtP14tLvjMlOGt2FrpmwRhXfY/QkQGkWRMuWE
bTOKc6SYr3i2Q5Lyud4jzIX4puj7UGcBXezzf7Lq10NsrSreqmlKkjeD0ahXZ3Sw
60OgtAF/dLQzOvVJqOBpBfHzPhonSI5aMVdGhz98nAMnDLVLGK66JgDA9DoG3B14
sVhl1XCmLfNEcbwDbeud7dbD1nBhCSUB7WMHIzPzIgTvkEesRbWo5k64p4ynBYgI
LqRhOmN8Z2JLJDtnYpVV/REaay1TdGqqgr/H9kq/oZNT0wolc2Bt90II5lMc3TOH
P27s3zpbgKBidGzKsjniuTaOrXnxxEbQQ0KWU9eMn+KvQLhCNzPLxZc3FS4srxOp
nwCyImjt9pJWsvHWiF7rvPyoWjINYvZON+iscdSXYsABj8kCg5+Oa3MsMNyj7v0r
KYJCMcLg0Sn2EqNWjftZtpkXWpj90reWRLbKdEyW631RtZRE4FHAMsRxXreUhbbW
ydUgC5DQWmkWTQ7Hrb6Nwxk8R+0kLl7k6Z/QaEDkWs16OW456ewt5XMmyPt6l+Qc
FrdqACYqfjbdi6UVQeM2RXi/phP/BnxmLLhhBE3NCKsZFfCh1Mel2/J7LRBtNauB
q9Whuuve9SjkeZAoLeQsh1bRqoQVo6U6WPTRXZEBk+e1GQQPf+GNcnK4q1ZDyhhF
ZomnOfOqMIaI4HJIMM26IXMYJIeloP2BGnY/JONG271FaE0yCVJw9fUaplCfFJXw
9DN0P8q2y8jPJvdXJcpyLmHKzVdypBCbda1yWu6ZcCT8r0t4Y3F/0lj8kRF2Rjk8
qLo/PTv/P7YrRCvY4EEIoe2OH4zp6FecVZBzjl5udT1kXKVg1lBsfFEJgUw7brQx
Sxj0g+tV54wOCsGGjBK7+rA8dNYMESc2J2LCh4rkvQEni56XZS8s0U4N7vyx09Br
N0F4Tzcze8XoAnNPfOcE2yYHwifsSxxr0wLtvfIAF7yTIAp7Vw5vmt8jhm27rTE4
sYQnynMM62/focMwK0xvnM6wPPU5l+gKCi+3hbmn8SbQzyK5kzHjzdoTgvI1vaF7
Y0cMNWEpvFAr517d6Fo1ZbAGc713vT87RHv+PvXcs1/pJLx5LRq2XMSPqki4xooE
FQ6TIZn8EgVl2KOctBnT5K9rrdgouyQs10D8kQT0CEwcQTejB3UOxK1JT4AAff3k
ISLrwW0H01ublASLj3e3ocT3GVE5i+r8i71quv4ZabXqF+PmKPbzhgue+i64rMKp
vcCyVPlKRpTnEMJ2yHaS4y3zmMMNYL49LVZqHI3KKPp+jATod7lvkKLFvLesflem
O91puvh0Kng1G3n5DeqjKDQzEygT/j1WSmn1dZdLwFgocagz7Kma/X98yanXeSWq
hhRkLj3NPXHQ6jWFWrE8tYCsdnnu8BvgV8obgzEuO5XMt+2Yr0Jqcj+t2HBvwE72
wf3xyqqq9qx3wcn9IV/pFE2qtwDRp3+OSybaU+Gzk06GUiIrhQIZ+62Quf09ayEz
fsDqCljuIBnizQLHttwPmUAwFzLw8fuk9h3Ht6T7xr2y0l4qIxZkZeYm/Ayn600Q
kVsffRGUf1r4qCzVNzwZHDQ/OJmVZov/HmZ9LVXpRW3B/hwQwX2S0zVddb/M1j4Q
4ER7tJzCEsWUx0H7pjkyYBOtlk9/ZfGSfli8yXwfw6Z9/uTfr20Zcu4NZKzDubGb
BODwi6v5XWtHOERZyWPssJWj1MEUrNfUoiC8Z2I43h4fntNRfq0VAq9hehgHSU3X
6fp6W73uNvCeEcPe5hX+rij43dBh9coo2QL0anmQMDYLYmi8E2XUuEKEZGialhLH
TfaJ1Z48so/z3Htv6AWCQ84T2ANZlSgcd9Qdu6lJGKC7HOojbA0xmSNzHmwrHu7E
C3oH9+TXxHh3GGmENIr+F1BJRgn3lggDe/QrnjsdfRNfIzFQySp2zOEFMALPcfk/
fQbCTwCNFhFAGbkbrJwDloglH2nxwIWHkALplGgTlMAg6dQCgihVctW3008ST943
X77JwSZpy8hzSI4Fwmyjv47JgfuG2UUTqqEZntGVAI2T5UsxBuF5cjNmI0zBrV02
vI2m6PbcR8Q0dH0ZyddQ9Rv05v24zX0ZzJxXJgGqQ4/ST1tR5yxWg+I2tgwwkctJ
qRFVxstgA55yMXyRrEIW+lr4u9EsMYp1FFzrIdLF/NNzbsd36co2dPpvP59QY8Il
KOmj+yomB5V5nzcRB1afqJS4FPbaVVhjyw2kiv3/+2tMt0PhC1zcYqihJhjECaOK
csBx5FFALmBdVP6Gd8oGQ6dWhr33Rw2x2AFqT3ekbq6/1OiD9d72dGKmkQMbImwy
ixQSKwcPwA/WYEmsMynB9G2On931JvvEFnxqFDJLAPzvr1ZN95PDFmjzRK6NNsTd
ODkjckIiCZCBreFVCXUG+6tYX0OZFE2lCYRSNi3DO/4OGnPcQ9rnjOYQ4Z7OSMlv
WIY8PcTjOM1V1g/y9w0UOB7bzoubOII/KCh8IlRmw6TwbkPcd8tA89cSP7Y8iyzK
W7I5QMzpGFTso+2WdZU+XxkNlXhCB8OEk7sd8ho3KyMi7niAHSdDEpudvIB7AxCT
Il03nODNoQ9qJV6oeWhuRbAjHZTs3Vzr2SpPKqWAiGercFZrqFmOE74k1RbQMQmI
Ih5wLgqxSjL9sts6nt9hZG775hXMX1qG/0q9JlefHn6H6yF3fVCorAiNT3inaum+
2J3JsITeXS6R/m2X4pq/gmjCjO9EfP4saGRSoJSfjKXf8n5A41k44Sf/52s8N83O
UBh8P7MabaqByq1gKzfdFbYcpvFeemxS3yqpFevolj3G3NzOupu8ue4LitS9NSaz
sPvm0jeSXJOxBI8ZekYerLFyvuvb5+uSIiKQtgZZvYFdQrgY+CXYBlGjo80gbBIE
uJDrJ/YO8p0ThM9BIuSx2F/mBNSLi2Gw/sDARp83rBzXf3kSxlScgdyej4dYtLOq
2T4x7Gz7dP8AxYdBn8di5b48LYo1IONLIAga0gjvu7X8dEObGfj5pDmNKwkc5Q9S
t+h5wVGQ44aHKpxajVyQHMo4eMWBehZu/Bgay04YF/HgnHicep2TAYmok9VUUg4d
0hF3YlEiOcs508jwJJOq2IK2yg/xPpc6XU0wRoyGtXTq3/hgb7WtsYE6Swcux3qC
u6D9byD6iZPUQJ4oQ7mrnyAsds1Voj5cQwGdHqMJx5jHnpEjLBaqngztn/nXWzto
+hZ1FCHJ9kTXiTaCqklx2ls4MLUuZnl04jfJiR6rxJXqtuUGcJeSC7keexZZt96f
PB2V8CqCxEoU0HCEf8JgqXq0sCHvsMaDRsMQ3M+uGgqeKs9LiIiE20HQZRueQvvs
EowhbnGJ2Qp/NWZ3i7fBEeFwWzLySOGqAc09obTLGJDE6xEAZHvLEZsaWPjvnNZX
zOZ5mZRqqAEKSAw+r9bfBzEyD8pL4cSB1IdwkC0LQcwmIHg4JpbKxu0I3TWCKmuK
3RKsRhc5TQRj2BVk6nE6bLTbF5tLSJ8+RAqY/9dQXSH/CqMQmOTAy6tVvsUObwpb
FFa5f0dQgAJ61h2WEZ6bS23osXjXm01AuPK96WX2YKlbdiLkd54dDgRk8J2PCoGb
ets9xQORFzJZi3gMP55LOPRE9ppLcoEKPZ7McbZuAWiYlNKc1rdTs2kuA8Pa760d
9VHJIabiWCTSBn7abBkLnmL0irtGU/3t9J+mKsDANUcmGsD/x0JnDUHiuj+zTHvD
/nclSPiXeKRp8sOYTCNbWmwkCJmCl1pzsnvG8kgONa10FVY2U8l+y+nIigUa3KNy
3xUFEsDeMBbhikaH62fcUn0HTF/yfGcQcuzJ2S9nu6TLO2wZXvHFcVHbr5yMoGyE
/wqmnoDk8TEvJbKtMExob/5ai+jpEyRkhNtExGT1KC9rbOZW3VRJy0tofvgUOAx+
HaII7UoA7GOD9SuYd2z/Tol0Cj96aygcXWQ2ufx9bTcAQn+wueZkreKBvNx7gYTQ
4QdePbYU8Nn79gBz/RmYgy0QRZk3ZnAZBDBZvimaQ2yYl9y6hPrf8PbP75Ej+SIC
o3XveQ3rBLH06do5Owag1wRErshqdFrUZzpV3rEUo1B94Qi1ZLUd7fbnG/HC2cE+
EyKkWXKeQzc3LbOTbwWf8h9KfeRaDTGd1nGnWG2bcb2LjTMY8O0TOb4S3vlRHvJw
AzXEJpKBQYlVQZUFlxJzSKtxonjhL7mlSShhqQsYct9I8+evXKT4uZTfTkCF5SbF
ndxQzDtxWPHfKIwskmHXDgdECrVv0LVUem1B94eFHIjFZv3j9wVLrOuD4PymLICr
e1r5iZgwkCBzXd/D6vdAN2wf+/BciCS53AsxU1kXzAkWGVLR48G1cLXkQKYrLUQr
bU4o/q63Z2uDaGTFvFyeITWVTN1W5tBLvpFHvekm4nQJhhPdVME20umWwcxMkT+T
B7bQeIaHFwmYX5fnHBFuXpbELRJhYjwOZLt8Pqw7IJc61sPz9OMmR/bRJHE9Dt/W
0GcEQRh+/OK7C97BTjMO43N/c/0gl+pVvJL1RH/Ut7lfTZz1UC509XLvL17FT4mS
UglRqq6bLZhUuD1dk35+PiAcK2iVz4AmGJ8MfyPwoy+VQaN8D0np4an8WgVEFMMy
i4Ozdrq2jUt0btxJ3u1zPOF54fFgSabpTj7DyUEycfygdcpRNW7gTaeeuNq7WyvZ
IZWRPuu9uGrHWb/Lhsq0HYqRRSfQ7Xc7aGrZjxZKD9N7MQ9oE2xp9lHwWutylS9Y
5opUcweRY8Sm3A2ZL6xCBNq5BiP1ldmGUaLf2OC0G57NXmvci0kaMSCnR3y+n6u3
pDZIws5as9bJ6Am9yljCWPBLNFX4V7QxePPoVepGyaiQ+2m3zwO53A7DHOg/nJ2j
IZbRRbxbMbQxZz5ayyCRXDS3oXMpSs/fmfH9NuluWy/d2VkYLiMwG70nA9jPgK2c
4Yyr0+evsdW47rjtzHla3xQhKbKhevJt4fPjS0ILdQvbwIxDsGcudOcjq8kPphTs
Qk0RM4ZtPgQ5flkLaczClmkj5RpirTvfqU8c7UfrhM/HZRhimunRNh5zwxO4eOzY
T/7uCbCLW5rx5phd07bJS0x2zMP6+pq2kLGeYSSe5Ff5oOnPojMl0VPLqasrJvyl
rVZfn715blyinGS5vzTSmsTPN/3EUnBG1JW50QjgbYpOXlXmHgKhUmuvNAbx0gGv
ORu/2O3OiqQPhVIww1I+ET5woPtMOOpbkHT5xqOEs41nkksGF5k1vgH97IQcxjI1
Sq3lDo7glfsnBdlQHjs3ixZT9mtT6c3filmeosh0kWZQv+jXZX6nyiXHVeu4Q+4Q
2Yze22umEJcO52DVSVpBklCEy5kfMom2uZdX81oZNHaitByifJo1VPv+fpUGyOEl
hhuaKDtl9noy6KbziYbYwcz3xA8g87YRW/NZCp2SDQspYwJg4uRejz5Gbl/7O7H5
gpg5qw/f51ykcfJB4MdwKDqnhgukJhXpfHZIX5DUMlLrI1Grk7VZ5feAj1nMJZre
KCpEKu6uLUGuPb6rkeqbjTYG572NQ4w8oasdZqVa1jy+VjGzXw5G09QfxhO1mdtV
DDdFsHLA0i2TRhmuTsls/AMgVpWcww2WYabKaywGwwpuU0uUYZ3j4mQnvztxa/p2
5tQjGC4erFb8K/OBv0+V1thaXR8++efsSRMBDQOUXK6mlyqexqDRnTfA1grCrj4D
Yu4iRjo1WQCO61d0NlbVKh/zfYMM/hJypk00j9grEAFuu00TaMR1vUlaixA2bXU9
qci8N22czgoYQBV8dUgPqcUEN5F9wigiOT8/nDQKdZ1AhMyRyTip+VvZpSIxWEDw
+PNkP0GF95LzOvFzk5a+8yMp8U34J+ocMwZ7HRZ6hwLVsOZQWzjG15n7cBQlKnmr
XNKXqutUncNyS2LsiJRiTQf469n+sI4SNyLxf/oRcLfzfZNAXpmyT9Z+h3e8eoEG
CFkAwB2Anp5J5Xm+hAOZh0JPIYJoQ4FO/jjzp2pTMA/FggINIwjdFdLPuTcQWWW5
uYo28T8LamERJNutl7wjAF3GfA5O67spkuYdaa0HuXPeyQhmYUN78RmEl/SNLw0S
R2CEA2d9My5YAuVePbyJjjR18EBlQvlXXyR/jMo0gxCNXUuu7renwa/QLc8MT/kb
1ykD3TifzVe77LabAHxFHD8aTl07xxZKEE+cc2HAnmOgNxFKRxKJo3lC8p59xVvo
WjtIjE1x4fegJxDTLai9w7Wj+b+QvCw8xCZKukV2ulbU9N+JFeaexULqh8uQuOQy
Ww8q/56exAm8NznDxgC4yYq40VpHHSaFYvPSteQ9WGeN/rZen9/BU9uX2HRc18xL
oEdgt0+yKXHqt+hu/oPS4KFEnM9zGg1SB2K2VWXH/h9j54tuV91fXOC93YsLxxMA
7/h6v6k6xoevy78K+tXLFjCtjYAtVp2haz7U1NM8PNL6MQUgoO6wiHlfv6+OkMTg
UtycIY5T+zJLbCUAidhD15u+QyIrX/pCq//c4pzlvI5uxbKn3pm3qqqiNLgbnqo4
hsCPZKer4uU9ALqBg69r46o82JfuPcAUedR/st1kSoKbnEJ1vyuXH9e1119G3udf
epd7gDrh1ARIQwo8RjmP9whpOzzJC6LXRxy9NbmjyybRN60C7Zm/ZJF5CYkeIShN
UBaEmn2w36oayt81lyLryjlgaJyOhc5gT9RDMoXcV9B/RWMpWQ18t5nFFbdl+MuJ
F4qM2MLcFoX9GsaD2tjNe95e4l5rlMEDRE+glRXE9ZCC7JivAYlk3YHf1P2s5gMv
pb3jtRZ9l2rqH394C7ujl4+SYrdAbMrrUWVIXUKIQsaKqDFI+/Gt14PDqHb8TI0c
NELbvH+8/j7Go01RkWK6odVqWQ59PtvmrWAW7UKQCANdmajcrfYN5aNRWNzmKKkA
zBzB6jmqPEJ+zSdQmX9eRLyYF0uisGElxsXf2uZl4wH42yryTUEFcvDbglmMEpYO
GSp9680/AnaPTZO9tDt5iS6OTMua1mJ3voCyaXpptkuhZoe+XyrdDVaT5UaYJ2hE
zZdJGopm0wVSjG3RuG2/Hs38Xz1d6GPYRNpy8BFAHaljA85nLDny13u7ZJiP3guj
YSNhnVqmINeJRkUbRaO2NDsO9hC6MCm6xrxR30EvMTi9LY5ioymCO9NUILXgXIyq
s8Hb++2nAqXyT2BOiGQMtSZfUFdjQ2FZwbEn7PG4ocqUmvUq7RRvNc6rHUYFAi5t
2ptq/4QlhZsO34ZFu+zpffvsyeRefomXBeK2wt/U9+zW1iZdGmIC+Xcdf/C83pGr
MOZh1ta5XyTMgRZb4zKCJU7ATu/9kHSs5CvAEE4V8oMbQmwsptkLNmwXR702boe1
yvq0Xd0X97rnDe8j0rYQ06WY34l9uVIREG3MK+0zcyFxe8l3ql7Y/dsAgPouRvhF
k1V4VugMOSDyTfp4CAtVVDg0ZSBmSEJpqxtlivnK6W+EDC3KCLgQ2G+TCE5Nc2Mw
6m0RXUgK6OqgYMQUArh1AtSrfpOxh3JKUfhyPdQrYW8uAebnI229glCzgM//+xG6
3VWisEynHmmxiCwLyy0/J40VrHHAkFLJ5ItRmpU4veqTU9Ih1TiMnzZB/8Kn//t3
IyPbq/XKk2TLe+quC6gq3ZU7RRO5G8uy1a/ZST4WLV69HmLA/JsPGs5GiRYYfJup
GSKKs2PgncdzND3LqNgB5ftXP+kneH52VYjeO+8DszpJUKVXDTJotyeg0wWVjmP5
T1qnanzkXSXfS3fh9KdiiKDcK3htId8JXvZizsqwWJZNyTw6MJ7GyZDTnfjSRrs1
wCICDjMUvKlTH12wp0n46ZtX16PVWItjcTHegCiicsT2diBCBfcDRSsCBg0qSx/w
IFFJNRbadW5IcifUISGQkk6TM2UdUzNoeh8IFJqAcdsn7ivETDFAPx8QvtV5AB3Z
wFnMbKMMoO7XhTfvfpqRPYEzmeQazvQ4okTI/r63x8iVCXh3mjVWOgSQrpLQqCNt
NVBf+snt/47gryFfsTV5zxm8YZSzMlsoReeJ9ak8K+1kXpZU06cAI73SzpTOhui7
PSPl2jKMmP24MiTEaoO+j+EzNBxvl125T9fpfIrF5jX7CDeReBNi79cZT+tWCwJR
x85Aibs3/d4PHrd5Uig6YtpRyZFFghKs6xAzkMiULTKfQSB8vFInbAH/32iEUbYB
Q0+d/RkDKFr4BKg61QMZvdG04qkcNsS5bHo0V7N1Rjkuuu+4/hO3U8TzW7pfTM/d
nmm3HKTalYVXq0A41GPLm1Hw9lmmJIl1MCvBN0jhqmJccgbRgTpABEHQ5xi8qYRC
BYxTZkgZPc/0E4Bb+otPCyxcmRIgc1vVirz2/8tt/TziooSvwHHMHtNYIrv6z2MU
ze6goOpeLPY6xSbX4gpMtPpuZ81UJuDFcHgIzZMJEVouHmgC9Ed0+H+77cYCh+Mg
2QaKtb9qQ2oFguEXOX6itURg0wMi3tTRZxBLo9Gp0OmuAKb+MexmZj4Slt2UqgHw
7PtbKRIpGGH/udi9/hgnzz8+F3RwSyorXA+1dJMeSnYC2m3mMjEES+8myHEKbObN
exf67HAOF5r1biAjU2QA4ocPUjdCalzDb0j9jmcXtvE/HtpkxIBLdHrwDqabYlmy
LuO9y2nFHToy2aj8P6RdIJo3aRCkPo0XqzEVfvj78GsWHJXRRi1yEkoZ7ZBNHmuO
ak5f4K9qbEbY/7G4V1m/W4fJqq0fdDhinD8dWzn0lEVsLDFDdldQ4lvgthxB/8K6
x3kT6VO3Ge9n+4La7xqmcvyDG1cZcX8Rvr+gn2KPN/B6VRwSl26BCV1nD8X5zO4R
hc/eWB94Ha4GBKI3PDzVqb4Sc+nsltQBQze7WmQG6ythDTzUZczsYN+d7oZOmyXK
ua9Xjf3kYMr/5sL/intfyPOkoGEm3R8E99TBQOhUDx9JCKkZECl6V31immgaFE1o
dhICkESgy2PchHzok79sHfpyyV2pItpfhqNlJ0p65KYqJVZgSfyg4EK5ulcvEfVP
2rivXqJ2almqpnE2sqcJBkZw4TdGsfe4R7RYxeef9SLU+GKzPI/aeX7+7ygBQWpH
d5Gxp/fJA66ScMvLlIigDlZU3XQPSPfVcLQ34vGOZKhOZJYirrwomhmHLuOisB40
kDiUgSYUdeMcO3OienDCEXVMaYlco3EKxL+DcffoitEfWCeZ8d7xW17N0O336wS+
5JcgzhLC3hksf3U6rxR1sujqtNaFBMPs8q32Pd/q/0SBsIX2tgoq8/tWbrrq80Sa
y5IshA4jvN7yu9G6wByc32NGEWc83bYEPATpb9HEbNzOkFdozn5E8zuUimDdTXIF
YiN5z6o3JcT8wj0JWJTpSoUvyQK/vWOktlEzjVE1pd9sq9czmxLW4a+Y9kV5e05P
/xv4ijIApeo6CUKY/SXxTiYG3caAUGDW6kItK/fR5YUqoZR71kYhlXXPdXIioX5/
uLLauRNPh+JR1p/3+HRFHwb9jTv1GXzCowMs2NsNWMkwh6tQNGT5a+jtGT+UvCbE
ZkaUmFedPzeHWpPTmqE1De1Q5exZDfYv1veGy5qzZSqOi2zlkONR6vLSoffYi1Jf
tA36oEwzYnZuaig6L4Fq4jBRqCyYmL9FfNG7ezX98wGxGn2KtAQJMbfGCK6OVoS7
Eurn5RbjJ0+NJapzqsyi5ebZe5w3LBm0+5q7uxeZaa91Y35Wt31JiIczxjfdhxyt
USxVn1hQ0Vd3nFxVYqoINT0w+eTujCakJz8r4ta56Hjc8lLOeIknBnXFgnzISf+8
NgDstNgAxK1FPgslPYDgbieG8l8allUyvYQH2VtD/hmAihwdlRMSbnuuEjJlIm1x
nIsx9j2TR90mWN2AelG7KjiP58rUEN7Sw2xupyIMyRG7ebGWQhVKSvwETiMLhFBu
lAGS21F1FKXnEU1v9LJjoiM4SMX0oq5jN6kNHEGYI9kg3GOGteRSIeP7nigE1LDq
9uw+jJFwdkJoDH2lh4NJi3R8EYS/juv8Z1EJEQT28o3eUp6eTVISvhZi1zp13w77
CONNvV0XtASTsKqnY5d21h0eNq1QUjc4kPLHDyxpj5/misUwue/XINarZqkvjIRh
LJ3lvTZ3/xq5QxSZAcX4DymSvC0zgnu6kwVKJpYZDVpjSjFC/6nFbBkwCFgL//fJ
jqsMlVZsk6SSbpf+PMD/j1ms2pEdxuAXO27eI6/f7SCRfTM53K8p4S9aQVaH8uey
XwvwcOyqSDXRkaFFbfQx51RILecYPJf/wJX9Hkf0AZ3k5qy9BIR6DshUKsvK98cL
U28z0TuXUYZwxJdguUWvRwR4n6KycsuBS8jVPjsv0/A8DfgbkryZ+iqZrzb4a369
d2BM5QADM3Nt4LqV4OEYwPXNlqbU+jhf6V6wEZKfHzI1eJB+lgChMWVL19F9UZNU
N24sTCYEJQzq3xWqZrnIXH4A4xPfGuoMhNshlHemoBjl/Qlj5nud9O0Lq70Ige0z
C/CF54TxHZDDdQ+C6UWRzRhrf3EIXw0LJ6p54wABS3hZIsa3We2KIIiPRkveZeJ1
zcjbKIXuXL8ep4SrKUEjfzItnnFYX5kp10k2F1wf3xS8vegV/mydpkC8Ss2SCU8d
ZGPtGsbJfvxBxyvogig8wdWvf0um2riR5K2NVgEm0jwaGP8MXtqHcb0gpyLqmXh0
oWraS6+kKFsFfJdMzEUKl45OTC4tnSkhQxw8PiK83UIGCPhGg/axW9vQiYpgo4eK
75jzcKIQb9gGlMiGjJ8Ezu+6fYxY5IJZpQ5YEzwWId/ygPX2qxZ9iNEz+GOyRbQN
ZrL4eelVOKppyy5ShNmpSPB51Mxkel4LnK30MmaN5XB0qDjKGWRAzy78w8MfXXGK
/klGq8pOCqRRkEJDHKuF76FBR9TYFjvj2xz9WjY5jKPPfNmqHhkeptLhkt+X0w3Y
KE/1TMQCAvARcrIy5fWaq2Ff6apb9/rym6Ttk2U4ll/Ahh2Oc6Uams9oyn7ekmOg
N3t0no4UJwVPuJGVl3gzM185aOWsoBLOQsFBvbdsnWoTpZP1RqjZvZL0PQS8Fp8k
vVLwL60oUDliDvalXfA8sJ+Iv+Fq782sTtN8vMEyixvPvuS1kILhmZFiQ3aSLVeg
P/9H6M+5hsx3rW+0jHj7X2xdk7Bk7+lyBvlo06NKVQVpnmMXttfS3XgsgkVNjLuf
bQCFLtt6QP8x44CWpSJPDfod6D3CH3ws4VCoq2DLPe6y44WPtfBkufh+fTyErb6S
f5R9ltheqjm1hV5hrfTP0xawcAZ+M4KLMiPzHBS7TY+St7WCp+X4icwHZeZ8OwjL
lderiIENago3zrpG0qCwC/GYNRMzEcNKYj0Ax1swlGlz/fwQgdznhNyh60d6Xmi2
7dLIy6YXhwMXsczeLI5+syMNRYVfhpDSyZtJfUT30vgxk7/ntX5HP6bKK633VDyI
CmKmYEUO9vqeuwbvvQpeD4lO24VxPdoulWptDa+r+DpHUJiYpL3tYZk6q3lVkIqe
PBLfu8vC3keQr0k+Mu+hGnIwBbvNUVlpJ2HY3HKlLsPUcJKtiZ0mVP8nLfLWbjJC
HvwaYbqe1OdA1UNQdbmUWL7/MBn300Q8gLwm7X66kZCk9rsBLa+t1eDiA7E31k8x
iACGlCR15OrtOUtD2xPdL9kAp8gCF9UycOwyVd9NksdPYGDEb9peGJ2cnjZUHeCB
poa9/QoHWwujGB1O6pkvgaHrsloCyLzC9ogJxmL9JnkvGINaQmV7Ih1X8DY/0VsX
ykDs2r0ZzPi/GVeAgphV4nhyX8++onQg4L9TPACynCdCNnEiL6vxlNfbcdS/6BAT
CiMetMRQisr+kitX6C7GhwuCXntGrQRhh1cbFZzLegh3VnwY/hzD8RfGs60ugrHW
sMcV2dbZEUpEqgfAVXYpsRagwK3ql9Idhp+RPzt8cySrb9G899K4FfGv4NaA4T3a
LKlTX/+slVxk+Exw8m3nyspXlKz0Gm8Xju0/VU0Snr+lmgDz1aPEeTgdrgORaITn
MIvWVUt469eQXHWm4ePemoBDRNz8QDbGLExQTTKmkPoc4iVXMjOS1T5xl/twhNFw
TduZzagPDfrjNEuQ8ql65DVhp6ClkPbFLKTHDZzCEN04kzDMMDI8+nJ5C5A4wypD
lkCSVIl2tN0fIzkNTNjB6fAXYe+pOlDmmy1asOGCtC1tFG2m8hcRu0gc0qhIsdEl
XnJnuj9VXrBmk3oP67s+HfehbYUeEq2diLwmQy9PtidqoxASFKvdi2p7888Gjw6F
gbgvzkIa4x+VhWNra+m0Hj0a4zNibqDRqVJiIILzSyaEYmhqo6iZZgPdXmqXGBr0
jWHbcj+lAgK+9IfcOvW+wqfsrcZpR+/J3ZXaAr3yEcj9MwuQi47p5YtBc0v9P5IP
YmpsvVaKNdH71ZknRS/xYCo0D6lwcNBJlXc0BEOog/Qe/8uZ+DyvgPDPz1gQ0zRS
uiFuOXIquhP6RIAx0hc56T3cNZ50DdCneUvQa3Cq1ocUUExSrZuzPOABlqaFnUmm
+H4QLe4wNM04DJCdbloX/mtOBCzCVgxQqwgWWMjV70DupeT3dmGO1hR5ihUsozUS
jGGr6pJ7J7om8gCF69ubTKyLTyzUiXmttZC5s/Y5tNnDr2aHPE4VHKtyBAZkxSVM
K3b0ckVwszD9LScdZEhGVidfHyNAQUDkMZMr7Q4LJgXXioABYZeK4ICw7rttwcdJ
2E8zYfDEdLv9q4l9wUO9j1Cx5GaVIEQBdMWEJkR+njyS4zUqnpJWdh+Eb41g+Lcp
AyREj6+1VFWTQIeYOGYdXwPMympw69ZvUjgmG4ksjJepqWNsBX8n05ieN2QLus9C
Dz6UQgnujjkzqTJPocSQjOyfKmBEGLfzVTYwLRP/e6t3VTo0Sz/SfXdYOLFirt8/
F/9VlFkIQ3qR9uNs6HFyEsZdi+MCbiTiwlZo1wfIDMPRbCVPWwj6zkxH7q/VZjBT
o8DPPpqM5KzxtMj0WPZshvoAaDnG/VqRiyjl0UcQlNoFqd8mdl/fPqPGMe959OXi
lBi4VetZabFJYBEyZunOFnmknRyl96zVchq7jNGEiTDw2gZT7lN+bKmzyfjWYLvf
SHTEuz0siOnnRkoN6sg8QGVy4fQ0pDOvlDNxs0RrgI6QapIoplsQhCLkTmn/ajZA
X5TVLmJrSWRlvapFf+CVNdGb/9bvA6VpKWL/rlTRixsw/w3VGyxe5v2Jym1CAYZc
V+wiTTCr7yG09HX45hCE29fnFXNNivp+4dRo/F4QxBvD0nSgI1fw7DrEBkb6evq3
VjqdXeNnfLlBFFvuXXHmKTrvvn9IJdwoz9RXQyqkW3KfQGxCfYbhdok+cztFTKpd
tkIJdVEngb+9YZY38QMJtSslaOELonvqb0EDHwriuiX4sXcwZaJFeTnCg1TCNy/U
a/f/aEtw2fI8RSuzlJg9Ejf1W+Lf5I9H0j1pSqjR33omKlWJxwAGrDu5kbghvjif
GjjtPuIwSzvr8hXr3bqOkimOAeXp/mDU6c3J1klwQLojAebayCaeNyBXEyDRdYAB
YwOVZwfKTbB+U7c+LAzpt6gcD6a1uA12JuTJXqRO09AZG97VUmHaiPVKVkdxo3tR
YmkpdEf1M+9hePAp/dLXHZVHDFV+6BFcpTrzpJjaxOn0O5MtVZ3oT/AE2c6rs6Ct
yVPEOYqRKj4KQ37UhQCVrDE9Wp57rTsHeZ5nwYoDusi2tLtIcUq1p1ibKOIERhXd
BAnBzUiAz/YItkkluiwNb39AXP8UgtECj+2el1kFc4V8UlQrk+s2BZq6q9I8gmJX
9QUKP4HD8NZNwABiRDApe84Gix2zbT2wUqe2xxO8bV6p600jTkXLvzH+dhL0D6gQ
eBpyhVBW9s2MyjMmDH6DstIutcDFmav/9gmLyS2YvOTUsW2sYuUa9tHz0X5DahaU
nxvRPOY9bkALkT16SvmFCfxMCoRMAm0x9aW2U722OznXJT+RopJUCvhbsn2ufanY
R+65BF4iBV3kgZwdzH+hVfw5WmYai8WrR05AHJXK0D5RK9iLi63Kjevh4Vj+5Wz9
hWdh5JOrLZnZPtivC4nhBK5oRea8wpScIAD09Wml+GH9Y+PjxdmctYKPPegCIZ7Q
Pgq/eJQQEf/1vWAO//y+MoFFIxqdkc+oR1RtOo7ocBNoDh1uL3ZWl2kH3E3E9JGH
WhVE0dNjNoWwrL27luVBSos3Ts4hAoVhFrI9BQwO6IOXlejfJ+w7WAkdML7f3xgH
8mEg6SXl0qL8dByuMSdAysyNdePqIbc1U4yJc9sgyzVm9iyMCetILOumDVAa42In
tzf+HLfs8SzzKn/HNdtdZo/5dYlJBtLtT8/USgufU1Mpjqw7Eik5us2YUsT7KGfS
jiKoU2NjLv6MDibAvAFsQ6cIhX1G/6SEaAA96fdO61JKOM1XmwK+N7FxdhZ6Hl5x
qTz1zgKeZDUgsv51UOoipzI6jGfdxknLZb0Q55huBYX/6zxwtb6JEYfftDNbcJk6
Vo/DrSmZiTaWssXTmB4Kat26gljc/5awPlAEtktl0h4/OXg0vnJ1lwKyrD54HkdM
vDVoG5zEIAt6RWFXdUVxyrUcKJHr0aePSjbZIJOQ5DKy9OJnxBCZeR8MBOZmGU9O
mtXzsL9IEg+5FVeA4k7FnCEuBpv56sgAYY48nb1maW/BE7yigTLMkZyjXnOTbqty
DG3KrDfPOIORcKXj02v1M5nYoJynSfBBFITZHw5E1/oEHjhWZxmBdDYXoo73qbI8
vMu3s+uy+OzqK6RerlwtROofOnwTV9QNWUrx9uNuBn+GY3fk3eI6j7F9uUvrTeqN
d+BmZ0/wUepbLuFXez5zXU5Uexi9afcAgD62vdrsTTj0Oyy0pfQswjrVsvhrQPro
tVc06h1s1YZru5NdcvmRbJ+iL3rTVaDIrOVAF2f8kSEyhvc2zauJzNSr4TYpGA22
9ltMg5l1QN5wb4Y97JNRIwgzYE0rHRmsESQHeM2w639Nbt1/0t+XwwX1YCz42hzR
F+4NcHGsLVEu8StjyqZlOnKeY9uAJkQM9ccA1WDbTtI/hAFxtYboNfFEA1c2xT1J
HCwjgvkAUxwcmYLQes8eC/GMsnAZ45usAvKgKxO0eNMTJ5vKqo7yk3Qt4xk21xrP
B/T6CkQ48ylZxpDgalXvus1dJ+gI1u5xdPNx71JT9K0Oi3bQ5NItrkJ6tULuy5Hl
XjQcws0QKF4aEEoNpk89OHNVtvF+iIGMJ1er6Vr0rCfOBPgHW4gUKCced62qyB6x
3/pOk0M6SsIn4v0bfa8RAZ32lzCWOKGkMnf/+7YgEU+MQSW0LJFa4DZPXdN8vYCg
qQLwvH8aQKaX1G95hE1/OiBX/LLMSuxCf1X8w0ik1A0QSU7FlrJ7eDpA9QrYSwi8
goMH+ZL5OL2tpwaBr3WFPR0pjCXq4PtPgzlXN7w3gOeX7w7AIObPmXmC+AykAlT8
pKWngaL/k57kmLgKoAouyKzELUz6/6sXsnBMqyFp0U+RPojbaLCJOwRVe3miLRpY
5otCZzzV1/hDkSm6rN0/XlfR2GDZ85juBSy7TLsVoIQBwN7gn50/1gpIuTV7+WAE
e1zGEoo/48lXUFKVnenSZzdwU43Ec6lDmtWzE1FuZ1Aecqb5CIPzbGb3VmnnDm8K
Ex+qqUZjLFEQgJCxoKmWeLlp7oaEcKLqixLF0xr48jMpbr6VuxtaRloetOk+U/Yn
Sl9KY2rwtn1pco5D486MQuGjfTlGHo+Ympl1lYsrrRvxZDWJjoWn1fJ27b1NIZdK
upths1b4yd9sAL57TamJcIUZMCystsdh4wCX8nA2WE3/rzzAxXeVEVNZwwcKmqjk
HjoI0Tn/iUWxX/Agtu/DQ0WmmusLrMtDOXkNFBfm4CYY4j2cKVQjZOc2q+uQ2eFX
YExuUJ5pTzylJb/ihITrnjzWup5H8n6ZON68QthZhE7nbzP/Ssfb4xpoSqYP+5qF
uiaCTGYbL7be7y3dey9c7wfmD7BCYECnvgnk5eY/UqWu2BmFtqJhTjiyF8KX1xR2
kUCj8MgOWAnpIVR3RgBq+G3q2+54GfSu5ZMZd1QNBPjihED5z+FP7cNDe3tjywof
YpYk0Z/1Ep4Z+Kii4zIfPCvF5Zw34AtFHqa17Esvu3OaKYqyAY+84y+7TKoNYdG0
TPBoiVO9f3dNhid4iu2SoRwEJe3phLKun11sde7CGG8huhy1cI7Ha/9JW/UO55SZ
XzS+ay12OIAisatiI8I0BYyPHVbmoHx4Ff6IW8rdmG3uM+RehPa5+B+kWoYOQXMR
z4G2pAeoAncnNpHQgBIj4VzIJf6nk2JMRe3hm/QGGWf7vJbAlIOEvGYl6tWmlyA5
7ieaR4v8bBa60m2zMEJ3XfbrWdquR3dXTJy13tjydoCm1e5qQ+hWeKjf4R2XH/c7
RCf1Bw496ywRFXRasWIfVFfqM+nLP1TEA3Mp8TuQgv1KQGWS9GJrwPBxqrDsBjtQ
QPWjRV+TgP/HA+opKeNko+XeTZPVsjRQuSGiWFwXFnC3HW2G6x3KVUMoGX/1qrkB
+HS0i8EvfftGFjX+dQedR3zs4PdZwxuAv0nV9j0TvScIitmUsokl614RC1OpFJFr
d+ZgT3Uc6sGzLsRm+mlaWhGhyaw95EONYCcetuvhHKSi0GGoKXdW/9ScOnvFRWXj
9j9eVf4Q5fZ4rcx58dutudBohaK26/nK1rNj1PFyI/NgqjiQsLNl1Tpi0n0XYe4n
k0TQ71VNucqrsMFWVPM6nsHxCED3ohBVjjpa1g+uyh1bwa+DgXaTUjSl0WWqJ/WY
7AhB9gIVv+K1JsE08D22uAf4jxDDRIUxdkx8n1GAxoo2emJFb7JORORo7V8up9mB
7Iw4iPQLegkcuOoH0j038rdXNam2bCSMV4O2FqavgrK5PG4QDf6FuE6XzeHqt78H
9C5jG9D5nqHv0WCVpbvcIkgSkgPZ8qtSY251c1XMpO97a2BJzVdnxJ3rTaPbbD+z
fbYjY5nILuTgOD/xksJ4EcNg9NkJjxf3DIwqNAFc5RZBkYBkwz9+5Pvw18zkIpxT
lR8X+w4k/CsjOvO/VilwUtluPmJoLnH099+q1W/MPKF+E5kZr+IFgBzar0ap6la7
dkKuAGPAqFoqTmf0gH6K5hdDmqlSGzfpz7RMYg6TjJyEXnHuKAoHsPIzvDg1J9wU
nTrTsev0e+NZ/vgU/uIoG8MISiSPf9xtFg2142AY7ImpVdu1fsLbNxVPjMHe5dM3
L/qyCvTTX3bHBubHWgC1fb2McXzIZgUlooD/ylpRLICJma/41A7FnNiZk5p7rD8U
wct+ozD2y3EuWJvH9j3KT3LI/Fyc99bOCgKl0X22Z9MO+nyuMcMKzuI1BUEbr1pV
wnvOD9wIhX7kfCI2VAtVS2Yc5wQ1aIuH82L9lZBuWGpqiIJMjjeYgmWefW50P0TK
+eKb+y43KBVUL1/L4d40TTYBIJVvYbVgCPdkTGb8DyWfl5JT7sO8+KM51VMW/sIJ
KZaXcRF1v0fVbMXs8dUK/rrza2HvLj/xXYIi5q+3MbLzHebBh4ODatcI5x4PxV9A
tANGpGhwV07KqOnZcyzv7MbYT4HozOV7Q4mtJG/3j+3si8qTkKBzVugpzg9o+Ks3
z2l/Dfa/FnqJsSQInRTzlEDGWDTX6Q5iPfSpPwvJM8rlr/qCL3SRlB0M6xT5lUQ7
V1B3aFe0un24r5bOkyCyhnpWHsQ2fF+fJBM4jyELNw9SGzC2bhh/OxvXLe4FJ39l
5h6+tOZzuzByX8zzw0i8+hJXxokU7oW6upsWIEvM6KCvOnP9WgmH3q5jXUm9EY4h
xiJHVreO0aZCF1zZiyQA3/Jzdk882TvdezFoVU5BBemnFKd67sx2viUt512HIKlS
4Dy+EmK7CPqDNB5vBZO8OpjRpPG4jVCfXqtVsCH/DMGCBJw3XSlVK0t4peF0DEZp
WWz2Ch27FU9cRj8JpeYvbA4u+KikMsZW/96R1gXA1iZOWinl920K0DKfE+Ub81Wx
5VbZVU0OzwOqxKHYqeHzVTohxtOdFhQYIh+YKDNA9ARYPcWPgQMsUjI6sERflNu7
pL3z/ddeAMY4CgDRv1t+mdIGZHMCoMgErtAa4EW5uhNeBS0P+FB/iY5kmHTRljbc
R49SsZ3Qs+s+LjkvzMGFVyww3AXSTOSyP12bvdMbJRgNbXHcHr5nWLw5D1J/JXd8
x9AGiaXZw38RjOuV5L71bs29sLcPu28gJfarqQeIoCq2MAcinBMPXykrxLbbnFjc
aumIv4Q1td1Vkvt1D0jaZA8QFrW8UIB+qL2Mh5I04jyY2eBFUAXqXmEqrjhUMT/b
lQC0PiNHSj8y8txBL9c2dq4uU44Y5NbfKJGhvnDz8IU3C714iIeqDuAGTJEaEeIn
VfrhvOI5swE7DdfHvLZcIBk/mCV0sRufCznnAZYfStSwwsMNC7NHCBSo94aQFDFm
p18ME38Sbnw6yh1PcZB7d6UZYlJahvxHmtKhQ6tS3ptKzn0MfSVDipOA+HEo7ifQ
16TJZRjvh2TOCmTKOamixgZhPKRydrO21pWwQPqNiuiBMeyTDndxK6Nw5mQ0T+uK
4HnkJEdJKXArXLTjNCMBbRjt1G10WQAlcp2dzeh55Ynxj97SrW3TfYC98jKR+Lkc
9++lGhpojV+sB9Rn2IYMZwstsmMLfAtiV8bSDhs0dQUm01pOAouDxdaSERimt17P
Gi59VAJKhVsXmrHuLBL3Q4f6HdGVuWnvT+6450yfGC0iwoRdxuHQFQj1ufjtY7sI
cQsx5TAXnFTpGHR0pmOmgBurKppA79l2oM4VEPlaatw0GBqgLHR34DZAnx1K2sCV
iVKBIM71+oO8onn+eT1MLtvoeqiG0GT+VCMu5LCWppu9keawwQCTgEuOuhk0fFlT
W7YeJvS5ayjFqogUdwHrkAES3M9H5NcZ+uvPLDHYOvkvHW+9dVfJtD7gP4b2NCon
bPJeD6Fis9YU0UOgeq5FqHvPDSDD7xPga0iktj3fI0/cuAann5XN0B7Xi1unGld2
RvleynGxCChzVc4h2AdBGHtxnF7y7zUdKKr2yoxJXJh2UK09Q0xw8A0+aud2AP8S
t+ymJ9TiLESHuQd2QYY8RuLEUR+5BKIeW1Bcgt9I9cLuRlFlPoO3Isdp4d1wJqtI
rB6jYicU7cask7DbySfMIDWUhWYe/nJlqFBy3c8zPcbwXoM/iE0bHwl7A4RPKDwM
Emg6jzWhu+Cpkz0Fw8MjxD5jkjEDV2zXS1Pm/mOP5FW25LLWvFrYMtL83A4Xj2AD
WvJzAbw4b6WYtHmzs8dZUwb3XMYXEqcyMgFJOX0nJ3Xhy4Da0BrQ9hlW1mfzy/2I
0TNkNARqZGlLyevPWocg2X4cc2BjnA4a0lhLZqZkABAHBwbJVvF8aGB99/pBYB+s
guacAhy6xRELGKt+nphZbGjrmOZXLGTf9J4x4pfB3XvXTOhSO5I81bfMspqLPiSl
ZzvPVP1jWP+VNSxkb82iaA8QZEiQp/PXvAvwATv98WBpDfEDpQIzQWQC7yOBXKQw
wprtUjrv2zBKjL8qsfijUc+RKU0B9PXcXfP2lJV8Pj+2WFHOZMPBYmU2yI0Ea60A
SF+GOZhKcBzdQ9ewAsakrLtE8nXU/eZ4Yd023hldZdeiIMSd++pFZdD7d2+Zp0KE
zHG8hafT9BN8g6sgy/V6X1gWX38klAsZ6pqiz1LakY6dSGh/ERKNeWxa0f70NZw8
S4B2ybKvudRDUWiT9eUiT9u1UQZac0I2QVIdIWpauOYDj7W8o78vRWsoKPqho1f7
aD3S7kXUO1iWoTI+hN1c1BWrowFHukCydbagpG8SlyYuABZxAEqg0ExgZUFax3Vm
+7R8++z5kHHdbtTlvWFRnBk+QbPLB6NSDhml+P1Ly1qV6VnZVBkuVEPZ6xSP7xlt
AYoJ2uKJDjbzDSBPTO1AC++d3OowgkeeV9HQn3yjon5Uy1ouQDDcUDut0jNb9dTI
SN1ZbLQ0gkpybleaO/uebM/r6O7HpsW6N/I7HVZx7VZwUlIeBgcYm9Z06Nklae7m
IirMfH791DxSgddGnZg4rGzlBC2au4QpOpwecEsgnsN7uPCg9weSN3PG5eJ1ss5m
96jW2Bk2xQse+GYwvGTbJl9xw+UXkie3WdJG43NfGh5PM5R4y7wbcWZbk4Vdp/9e
qmMtQpmkBu2dclxflym/7KZomaR1grrX9NTHf9tt1SRzngOB59vYYaP15/wEM53C
znxizICg7NDOeoIRvx3XuRrUbURkRF9UkeS0D0e/MTo+WGigoO3ca/sLwxPIqHND
1cvr4sKhseM2O95CqQFZ8Q09Oj5TDkDVmbhfReskVzjvcQ7jqwnvRJlIxvYHUnS8
vC/aSFwZkjU0DO8DMNr3urS257rlqKoiRNCbWwsMuceDqawtdct1/m1Yb7ZPC5Wj
74HAIHAUYkHOzv/9/YY+HaKp+OsdrQA88YxQnNZO1JuCBHLLHthv5OdsUWig8+OS
/4DZ/z8eThK92z4JXEtGlivBCz8uQKPewrPpEkHjjIXIMPFxcMFVXaOdCjfiWqsz
BhcauZ5+xSUHuEvSpjYr5mzA4nCOzzCAVxsL8vD+fVvvyGu8t1y6AP7xCpNb3J72
IDnFxxFE1nJpHJlRdCjS6/axDW84RP8IX1IwEs7hcyUtASXkcy2AGx5O53nP7kRX
FF5HzMmq7wi/ODr5MJxn9HZCihBwvVJyBC/qM8sn8u9BgfP18b/xzPz+wNIN2pnN
/WeT9Uo6NQO2d5nRyihetAAGRUr0peWGYUeFwVwZMnsCB6auDr9dC0Sa0754C6Ry
bnj2YUSs/KyeFuFLEKfgo9pzgyyhfXxqFxS6bUDg3UUmO8JXTqS2FxfZo8nlpGVU
apNW9mxuA9eazAYX2+KVWv8DEA5/KJ9TOZDgF/QIUPAL324k0yAPPonWB+2Dkizq
yCnelzkWzHO7bVZEPI074ogU5+QKwKOzsIxgZLQymkHdTeDyLGL+mKVwYTPmxNca
zxkY0j76/VW1aXmRV7kRVe1rmiU87HmgPrvHD0N8JTz9tW4x6ON37+LVbSbLVyv5
5oBfHaIZ1PieMgxFx/VnC7u+1vWzesuUa4D7F0/Ch1e8alhCPjeYmADJyZ4WszM2
GwOadGb8ZDgEE3GYq1vbU8/stQbfhb+miabCxV7SqrhhY4vk7LYLO8BOvEncuPyr
oSo9JUoAPsxYfnRCUKqN2rti6ebp0LMS/tOBrEOWCAjHiNp1QHHNjhp6BhOolovs
wASQgTKI0dUDz3lZs+dQ0ooN2s+ztZtAzm5CcQMx/rsmiGtH5xdAZ5u2WQRkK7ND
v541tS1hBIUgc408/DdtDKtt3mVJ9fWGNdKiB4AE3H5XNP+xZeJeW5su+Y/UOn3n
Ti6sPC6tNZidDRO1qUM++vzMS/ifzJDI7BMCZp9g+eFkai75u1VgYDbPlsTRdI1l
PV9Juu/dhFvbATtg6pw/OkQVQXvLvbPbmys7bwFKJEM5anmEcSqb5L8hvpv/nHOT
iixiyqXTxJV+IXfkhfdNT4pRCGSZap9DdDAoig1zHbe1seL9JtdtXMznUPHqRTIl
Jnj/7E47Zi5uBOKm1CaS9zqANbujpyNycp3ipyC7Sc7bbmqKO/dzcc24xslvT3HT
HIfOL6aDIhKOnpdSTNSxIgKstma7Z8O1FFT3GnYGJn5AOVJfgLWlwHcGaKW5jILH
y2+Q3vgR7quPe9ZxJJfoU8QQpajRcFG4IXKOv91u+Nj73tXxQNfKxQTEG5Cx+cDq
hV7wAHQB1J2J6AepPn51XdOwsSvfg6NuRwRAzowxeEUt7gIFuq048SAQLJLpeHWi
4Z4L47q5DmXfY89fcvs6h0n/vIZAqr28gtLGlpYSMUAnohM6qMB6303DxCPEdUM+
WhQ+7szhLl7Dv2qsPoU29+nWt541/EVamFdgeCp/NMtvC8LfzeqY40dDL7mglTE1
QrB32REM5Y4m86UWugH2Hu6CxO8Ql/3CVWdJoDamByvfyypPP1hJDU5cv9QUYYcW
SmESgl584Vn73KzD1mRFSbim2b60RJ5CntBWEqog44fKsVzZIh9hVXmksw2rAzG8
4V18X3/rI1g2pMXDUS0Bv6253es5EHbTZKXJYX3iLyvE5v10XOOTPX05dY67CuQ7
E9XEW83BrUsCBULIiRdNmCJJ5KGtRiwi8n2YoQ8tZJkhxe8w4aqvM1RS7kf7e0Td
RVO531tuHIxXyuohXzJYChaxa0hzX0mXi2Ps8BIiWWmku/c5zfQ40x5bnW3NOJ5d
3VTE6u8KGWvp0GhldBnOTAHT3kjhC8KHtSNy1XC7qDX+ngFJLVH12HNVnBnYCHOq
rUlug0SmtPPd88m8oNUxJ0G/6b1GFaGb4EoTSRhe9NTKNSVmK7hHGYpG3xZd3Ngc
i5pCsOTYodX1YGTwygFM4AXNA/H12+1p0MAeneMEIo9gQ+q2ySAmYl4BTontHoLZ
HApERRJ8v4ee3SkSLnDBy5eCQ2UwO7noSOW3P5zgPZGIS+T/6FhXpTo47flT6duX
h+XjTENDW90xdlrRRa8nGYlUD5vn8RCjJbh83CoXcMcPyCmIfgnFOa2b1yv9sZ2Q
3KZgQZyUeH2nGtA22XTtUaJFHszkiATQpf89tMaT3hrpSO93spiEnfwd6AjEkPD0
iGPEeykIsKc5B77EO0GSAELquJNt8rzevt13Zobl2yicCEpAOozFyxJxybtz0M36
H8kKZuTI/zLE/S6CbSGPEbZrREI2tTPFaBmfLgFelge7/23uXm/JrpvlJ4o86F3f
2aPTK9AuZBWPdqeUsZyTwkNe1Quf6dnYisga96mrDwqWtmnxKqcJ3fygqlX66CJr
FIyl4OpUlJpnfoG82PXTDzYRyOzYJSaiy0XDBpiBdRN1Jo9QGRgon8ehllrRAvgi
aMsTHO0XrAwyUxrSrqilOzC9Rxb6suETvyzM7vE9WPKuJPSEI1lMeItyeZc+9fqm
unCwnEy4Saa7xJKNauXmouMYYEsY92P6mPakAZCKQaVI7vmQIFsLijxkXEgoe7ht
Tk4DcU6O5T0GqUNtCuWygSrckdtnJzG6RH/W3W/QcvTXl88MJMK9Qh0l39elxvCO
ogtVuLhZaBUyUsEUK82T3p+7maFL9Qxkfp8AvTyZLDqKL1XXzKRmYvJiluVL84j1
P5RcJt/lRBlBtvSo8IUalVjm9tKVOcvSONk7YJGQuIbesZ4x7Wgrfs3PJcW+SmZc
g3o9n3QCWMNBcYDSXc1xIWdjZtrpFFVcooAS1shr7jDwvjfacvPY9Ahp+sEmDjq/
0W/twXA8UOzykAx/11j391Qo2E5P/zkp41zmn8OKrUFSydU5hOqGhHrEugjfoMxA
KdEU+ilWi33AKeXC+VMzEU6uHt7NEmwug5610ez7W12ZIzr3XYc8I/jjLkgdwWsB
covRUuW3ZCst8BBlctZhRVKADoyUn54N1VrhrAbx6b8cI/C+kZ/xSPSo+iVULchJ
xeT3K4a0j0C6AwaVDH8Gf6u0UPwOK+wOZ0GjmqM0iSG4+9NIXosBWz9KUyHI/yxV
EqvdP9alPBpCQfUtfzkeBFzFeC7xuReXfm/h/bMdlLUQ9pEaC4W9GEQR/mGwj8Kx
M9hK5okjUoFN1/GY7HvBhwFiOKzLItXhFLJovx+VciQCOebiJIEWm/ewZv/omsKE
38uCrhdmOnBNdeLgxkFKQ1qxCrV3xJr4pJnH7bL/Q/CLna4lHxOIYHQWBdr/Ubvs
2aHtcQEwwu5H60ZqqGIQUAAksmrAR1IRur0R1bub+5s8MgAmNG1fkdOjXnsY82U+
kp/C4GyOps37ijVdMIpH2jyubkAQHnBVpHTPkE4x+Bq8dT8EC5f1ry9e3oEqGnfg
XU1MT0vw1pSIX74BukaSVCTqi4k/5lj3Gnhq5UUtHvvkwN6fz7FiAHkGREOyarUQ
C3KGawj9dDAmWaKSreGhwKcZGHj1Pl2v1jd607q3//6ynXGp80WmwUReumaje2S8
7Sytj7BqAxqhB0hXWKIgBAKl3UQy4bVSip5kK6zMWxAWTsm2Z2vyLec+KlydXQ8h
FO9bSP3AcJE5oTbOKiDnERFSfaUHixij3TExGvZGNBInkREG998QrNOBH3QYxM4e
Cw8EcATXgMDJcZNi17SX5wvUp6smoMoSxklKdu+lc3LC5SBDn6by+R+L/4QASaP6
7uG492c6eQ/DXIHW9rmFcuIZIs3cwCiy4mOMqnjmk/JG1b/ZNZteVhuwyoHJKzYB
9mxAWjKP+PNiWH9BvMzDwvABCb6qNLI8ukUOt0/gIkFVJVWfdl26YQQRcfNMEMkj
tCgDQNFwRs9XdayXranOLfE0+Zb4EhjhbKBo2V9FT5QzS1yc+iUCTTYURygoPomf
WblmBijTYXzbVTO6lyoccf6GTvhWcGy7Ll9lMQ9cuDcgZl6SlETEt0M11V6D+swA
7014I1Z62VGvdYocQ+TspD2GFWyOKoeX567pO4opoSRd/3C9GXYtViArU897HtQz
M8ODOt3YQpetJVMnBMAKR36N4ZWCmXKwKW9JkHCwX6qiJqydFyEX529RApqq3v9n
y0TQJE2wsNQ0WAqQVc9g+/XpEcnn3XlqVVZ1g+CUKMuU4aqj6e9pUsrkIApGq25d
6B8zdDtgmI735bqVaGdbX5+XQNj4BxRBAPQCn2Mcdvg9xkpJyW94E+WlmeOrVErl
QGU+Y1d8MKpTK7EvF8Pw/HAdCsMpQ+KhlubGnBLFrI7GiE5jZW5So6T7M0ybqwgK
hVBCfB1LgxmlvjbxYEpYsnp/9gCkewgX7VG5WXfbrFxF7v/US9SX9OPAZR6gSnTP
iKtzutMm1zgTR2kzmet5NVQMjJkRnTqQ0vf8cZzQ6yveYYGVqH6GWYA7Ws93Yz4a
MkIkDaHNGRy0jixkkYC6/XXd8mo+/sN7uy1aFGujPWg0HEdPs8FFyv2dlcqnKL3D
IiWpp4sIg6bFynE716wyhJHWEEvKqgJNtbeuiqnUpyZZEx86uodLcY+spMGZMj32
nkBvtUJtpu1DXoG5F6faH5fG43w2wNHEW7qpgwofW9pTko0E0yERKhyjm6FQPdCp
IphIO8L+AHWOutPR7jm2l4GoN2lJrgMdiGy2+QWrZZjThkgBCHeZwObXFB7YHID7
CZmWtuCpBF2zrsZ3ykPAlpQ6yCkTdx/ZsTrztxgFr1DV/BGhypvpLeptxoYJTZRT
lyLVc/A9yskZYqDFDMWX/zw66j1HnWwFCmxn/NBkVRxlbEBPL7vJaE70ONPKSrUL
HqrauRqI3frSwNArPkZlf/GfWL51J+ej6G46y9/GwC+yivj26HQv6UtYqCbVYZgF
277q+1MVWXP0d71tnxPdj741QxkSyAz1t8JGkYSyTOEqAlQssXzVJkeHMRPij6jE
AJ/5+4xGlWEzKrDmsx1qxwuswzES9U/iuPy/qaC6r3VhRWaw9uVC4YKNaM6W2Ddv
BSXFYoDOISeeKbB5JAFL3xxcY/noTAdWgrmB1bUL0XivsBo31fBKHZTIQvhVQPRN
k+PkjkMAXEseNr0kDd1HIV98YxbA9TuC0CJppRtoMZ5o7fg4Re8f49PiogUld26d
KNP0j/EEOAj7lslmEjD/P4FpKlnAAhDKUUY400xhbM45w5HWD0G7rfFyYUDyrJYP
wJObrDdUuj4lUxi+b6uMF4wnIacuAX4dFsTUUup9YwtMCWFBOjyh8cmCd8SBPVId
17pIMDmD6H0u8qPJlXQpKi0wagbSbvESsBT9z1TMpVDME4r2qH/O6gtp8i/0modt
MRtEx7/uxUb2CBLIfKCGjySrisvifqluLE+dQlSmfNfXkOYOGGUwyimtHF4aEoPW
ny3bq+bcYP5IBBwICbH6hwpDVOUtCRHCw7Kh7Clz749KJRH748i63Q5w1lnRnQUq
Y0kj0KFLlPA0wsm00QMHcXsc8WebdB46OUh5A4w2HLehANpgEcbp1nwiZRF7Sofe
TtcU4rKYxwrx/f7F1AMYCFScKdulFTGJ09CwDpLAZ0Z3uVr4AvDLsvKpcC9CMpq7
hAdBD09a3SRYc2j03kfKeU2kcuEG9/MfGvUdAQox9sRCcca/Nz2dPMxsBDpbKjJV
0qHEi52rdLQLYEttKM3OixREVbHqj6RzxJ+6J5ATshAVttizbLIycuyYn2dNuNcW
9wVE3U/T13Lp/9XdPbnND42gWI+o+i+TcVmA56PRw8e5Qn9Z22W2Q3SiXKGCEimz
7KBj0KaN87w0AGwe/xFUqaOfWhk0ALXFlx0v1sRL8aY0YWJt8apu/0q/kcvvN0f6
aj56kKrdxaXTdVSD7Qbl9jciUuqRmRg7ZX4hUr2OAIbdF3KQBYYDAaZ965eWclzC
WvaWI+8OmoXmM5oSVCL/GXGH7zYF01t+r34vXcGLjV0RoYkWAGHHqKYw4U7h0/3Q
Anbf6vEV1cg+cv4e051XCE3YqmQ5O0iVSJncLg9Iy1zTFokaw5W7n3QAPPEmkVZK
uQJZSKN2vgZyOddCPSgHOya22YHvHpDAv00cuzSPjU5isawnlkzPOegtF17/FjFO
0HDlPv8QdwJE6A3cObrGZGms9ABLntwUPgayHgI8YAz/ePyVMcRzkIG9uPNN9Bzl
t8vETi92aFz8YxSWQOTVa3AzJ44f8aNkt4FjLCkGyoQX7NTG1AYHKQTU9LT0mAZj
VXHWm1UYYK364sGBjFzeThvXBZrw9T5SnO9toCm2pK+WGW54+XocXSU7h25z0UIj
WbitDxHlDOCrKATAz91XHrtivcKc6KXdOPI9DmY/zDhGSn7K2Ka9t5qtV6fwshI3
7SKURQi2MrWNJET5j7scCVEM5CB0+5OyKUWXdydQ81UzzDhdXCvH11jxQ5WGN5yv
bOwZdoA5cmwquDNDtppUWyqEKhrrTcBIL5sl3JRjgNMNjb/wjQf1O+h9YZptW7T6
BCX0rl6jjmTbKMayqsUMIuF8g4nf3A1qzXOnRjm7/30hnBqMpIBsfDe5olrr1NVC
rvKrp5EU/SyeWVXQhlpbyJzIW6uqzLSnXfHzxw+tGYEaCxDh2nBu3nkbFv9LWFk0
qgDf7lik1IqEWcXfyE4nc0FJD4fTZcWqxcfXHmcfHbFFH7s4QvXsK3+yj2TsZV7+
3dFMAPqOCgRIp6vPht6a/s+TNPndxe+Eo8lFs6966T5EcNYRw5ideTCOpXwciUPh
8WxU4tye31vCBJPd3+vXMwxy9tgtWBJquOMiGvanGnx0WIcJY6Hvn83mg1E8TS9D
R9C4bDS+HI275z/kOUlAGGOWmpcm6vsp40c7qiHHb2ylEp8gCvMPdBmoNxrUXu/5
D1/OumiYpUBGFVur5MsLGR4iusb2km9m4fZbIKgv2t2ak3t9/39Lzls7w2wT0SNI
qNfSq2zs0urjgRLiziQaHvyntJx5KSOqHLgcWHkVSJGnXNT6yaCrdcI9vCQj34jZ
ClU8LHg4CEDaka12r6sK8lyJ4OIBHZeHi/NI9A3wpuhsFZ957usNUD9qBl6MO6go
hBnH60Yo6esjBowj4nPY5WCFwD++ZPnkcFBbvzc1qWFipCSl0HaZn3qd+rfVpuot
kUb3PkefrAT/SKRZ07s3YrSc+/JaroCg3TdgSNAoro0izEiYKajkw00ne3fHdY/I
Ofrc6zJ38MMijmTUm5sCmO4RRRRoA/tjW4NmtrEFLVG8G2Usxt+Dg5wzV+/upJgd
REQpVdaTFQsqq+eKVLxc0OLTcdkU5FXe8SJ/HWr8xDK0is/1Bhhe3ZBpXXdiHpnk
8sMr4pXAm6W8F2eD0SuRF0EiIaAdc0nXJicWnmhH0M0E3B7McyaW/VyZSsivKUYa
7RBoWAs+cy+Tne625C6SgYtflO76M6eVJC86xcbzRzsE7xGbfEaHvC1SicQwynM+
SfNsKPAiaFFYeq881fL8PmgYf8DMw8rrnZx7ICVNOSYsdBxwJTVd9ojntdcS1r7a
j7l3QT9iTD7UIJnREzgZroT8G83za4P8MBsTbsW1G6q/RfzhNT+dbbEkAce16E33
bPNwbwj+GRPQCyFc2Czr7rA2U4b5PmX4JtzYMgJexaKRV8p1m4FqPodREIy9lTvi
WXO/GX633BqPv+9km6sl66xqLAfBbTHBaheSNcXsqKd9atYQbKFDkt9TlXJNfZsw
FAVS9rtA7KDqr9hxL+VV8g1SFYUTGiLTRc3NY8PLaDMdtZljNTeEkEuUyXSTyLdZ
D9SaUYjGqvqvzp6C91eFvI1TOkA1VLz+VxmmmUbPuXbJXFaZEEWau1wpCe65CJwh
lreo5MdfagWrvIOiBhTK3Xh4oBXgnYdyNbvBSCJXhpBNUS0CLMbW5ZAKe6Lr986a
RW74SWm72pIf2Hx1A85EiGBGRy4hsERLql2ouBTJqfiWndxzaKWJfxWnD7Hkqsye
kmHLF0ltDwpd0fSeMKz+514c+t58cc588ubgCQECu7YBfelvzJEHS2UwI61mPivu
pNKxGocQIZT+tL2YjkP2QKFNqp9vt3qysgRUGt4E9IcsTqbM9YVGB5gwdk0pMfaK
nWss4ELmCmjIgAAKrO3y3gDEzzqBu6quYkxZzID3M46I+bxgtW3JMLU5s+mdedHs
TupIF+4RgU+PwqY5F9idF9di412L7u6Zhqijv9jukwTrL17ow2/Gq0Tiz4V269RG
XADUZHMOlEGeXhD2gaAWYhsBwRapNlN9u5b0EFb3SrR6sPztFQDh6X37ICt/X7oF
fDiEaHgu+abkduir8tP0+tgfTHQ4uiEymXfOEG+89Xy/sqrP97NYpYwzk6Rl+euX
4LVF/XLwiv0B2GxswEHaASs4dt3pfwTGZF7FQF6U/k0VJF/DxRGst2C02ne1H7OE
N65Y4GEjyrQL0ZAHnO3MKYQPNT+zzfDcVp4QBQcT36IRvo4oeHHeaGS9zgE0NWn+
ZTSe93V0QaxPl47YIk52XmgqcwNQe6481+iYamqRtu37dzo+lcfK4kckY2Pe1bOh
MWRe2p5dT+jbv4luhX4u/V9Rob+Tiuo4fmk0vvyFQKtK3dYws0EexTIt78ZvCBVB
Y1ndn2L0zw4+iGn10yWIEaMrf2Gx19MSAz5jISkJrF1ABAOwTlCT8r2bhDQZF1fs
L4ywk3slKKn0+UeLVuZTyqJ38aqg9GciGV4v+UKxaEDovDMYZk0M0g8o7f2AYdn+
WuwBwlwv8qHvDCGnP/NWHFnVqjjmeXmZdvOrdBqVKXHrB7C8xW2MW5l+q2HDeyk4
QhzHgMyK7OeP8kFflnY4DLfwcOr20R8Blxfppx9LqC4i2yg8GVL4O+8L+erfLjHz
kzDkZ5C+3Z64kpEx3iV4k0cx3Mf3AGVcOIcpp6+aghnFAvE68DqkiTaObG3GNVL/
AgYL5lSJjaAtBfK3p/YZDHeYvOIuHVR2zx8qw743h9yPwWEBBTf4ZYCC2aSNPF90
HiXITeggAe+d1jCT3g9A7SzgFDR/ysN2IIuJ77ocuuHn5DnzjHe36xp8vkmbrPTQ
4wvrUF4Ru+GQwFbHeXiPxjvq6IIKdxL5+kA6G7KvAFg8/5ibgHkmIu8TyDeudH9t
8Jp/VENKeK53N6woX9f8xYpEiwo1zin1uXOOiL4gYW39/rveDa21YbeKJBC8emEX
xrYiRACCmWzZi0pVFYvpb7jFb1AJciGjMxIeI9im2qmd6D8xDedQZ3Bu883au8CL
GPEt742/c09iMKQSonb1xQfP3CYUD2BkDW0d313L9h1Yph3cHZ3WLZUJRZxqCT2V
37Sn8EfN9tkhtbKuVjNngVd7J6LluqvvJJLxwcjULkt98pmB9KD8XIuisQgnFfBg
rS1CsRyGezppwLPEydw6nNrPrhJ4lyUrS/3z0CTC3buJTFxyuimfEZYo/FvYDlaj
tBrDGsEkvNw/Vx7IZplWBNapW/uHUuCnd6qniW2q6D6VZQ2BBfBeUBy0XnKXvJg2
EpdFN6ejFN/XsEMEoGp7d1M2FxPKpc73uQTtQpaYZ0gfv16XiR+KtCRhDtrQXW5V
XvhA+fBdd4Z4LoGwkE7/rqevDA2akbFPRUOMczzbLjxMv4t8nBZtfpWbVJC5cIGp
GYFBZyrRR2sa2DXPRvHcNQgtFbW7EmIrFABVSmlnZbshCasiZNNF8rrmaygji32O
zkIY7DLu1Qqab3ex7kh6GqtN+GgIvFrRxdqWmWhFtn9RyLxfBYot4on9Ymf9Lk3U
oacUPbRGqI1zufHyM5Xjjws4mRpKyUI+A4iX3E+K6LkU70bOoyphV5D3aWXWkXjs
74Z6KrYczcwA5/j+tD58jwBiOp6+RujuTI23bHuHZVmS5Weo8KUA4WeZjC1nJ08z
PDg9vCQOLBaaniYkOK+4KLRABEB6Prl7c1l6RCL1dziKrYXJRJC2PqL/K/DG2W6z
bkhEX4r2tGQwgeko1Psrb7M4rdAsu0YhjVJGyY21Y3TX3b3X+Pq/kS8wCIXctitd
l2bFE9XW4/9FxVlmmlnpNRzD5Ox72CxB4psPvX7g85vIhXcnRoMHhW1r1Mc/HCEM
NGmOoqd7c0y+PZvRlqgvCgJBvA1xaJM6rJ9pj/4yRXqiehofhxNTJ9myniMYLUeO
naTYdPUe0UXgU03SrirRVzA08+yubn5nAQZn3YUmufqCMZWv+aDjiACx2u5NmWHI
USHe2PGshPDPpz6v6Gc1et29Khdpn8mrh9Ep93BQQcfdXEvNeBXO6DETHco8XW1Y
gpZcvupt2dS2pRjdhgMllEtyldV34F//29GjZxWMQHs5Fg14v0/H57o6DRDln5mh
pnf1lY65I0wd4L1gCnedo0IaQHuzuKNbDN05SfeSS6RnZ2Bfh3vk5mPLBaepl4oB
KYqKEbfrEkIofNyVkpIcjYpXpkftPCVwON/ahNxYiURvryr9PL46q8xGkzxPwS5t
lJ0ELx6wiQjqer5jGX+hkIINvqYTcZHC6sIVmKQMROfTIp/cZgt1TRxGEZVBBsQY
Prm1Ko6yKP7bpuH1ndqM7G7w5PLpk5fNDwTDAJ4SVIP5ukH0yU4mWllV2a3cgnqm
OwIhPs3+rNYLCnJ30KCwriaZKYYXZY5sGwEDB1jB+3OgU4DM1qJJnEugoWFAmlnv
Ns6pGqeVUbSsM5kxST2mtqBKeVjsAGCj8UzTiY2P1WA5qwK3OMMZ/bFKMTRUuZ73
u5uM2GRJmFTvHsO366AW1XA+v796BSMs1hxZRyctGPDk55KNJidBsKHj7QR3ZhA4
ewLU5rZkOXzYIxyrcc45pmQRLDzDOQ4nZcjpMwQe+Qv39MV9pNO/c3xt2WAsIil3
gOuGfiRPWynWZGZQejF2DQ+9p1Rl6mZ9Dz6DZIxQiHsN1ZoRxyRlTCvA+xmyUORx
tkuALrBt48vgWB09sQq6mPfUzdnK+g4O1rO1htHh42qa33K9T9sPAAcynIPIuHRc
kjN/vBLlT4ahSuMG1CB+woNt8rgXj8CoAJeWhcSKzJoCVKyyZOgBourt+a/ZH/1J
fQ620JPoKB+TuQr9InnSf9Sg8ww0F4E00s9d/Tum/a9zxXO9+xl+qgAN1dcqcT2L
ilm3nqueAP39VYiZbCRa7zeiiR/J4lvhQppX0h26k9AELsKfBcVmyNQSPBsCbquy
a3F4x2MwKAQFVreQu5bdRdBnYpDyVsicFCbhlBsA5/8k2ngKjS8UbA8+Zp6ltjgl
zmokeDBv/Ypj3KOv7YPXtK49tkmTHclCiV9/eyXnAH9+4gGVs3KAvWdOgsqHpWMC
rm5L/xpdxUKYLW0BErVwQh1KD0KnepbupM6GcsL+rfDR8r9FHAuwHkHiR4SJeYrt
igKYM5do2n1IStmsIhKyikbpekj6cAqL2Qh3U5g+QpIjzGqXEINAZ+Crw4n7hj5c
6N27KX4r+y7LFqtetrvyAAqtzkhtGNGADEBPoy8nKiYw3S87gi5sg4QHb+HuVVHb
DlyAp++rS+rGjfDz8Va1YRlsEPi3n1HVcvaEdzxy2k58R0way3M+LM0EtwZd7PRU
kFFwzrmr391oFlov7P+2MZc3PNB7GRz4kpA45KKozpzuVN0NZhlOZtbRITXKaCfL
QBcMez43fciA64uPCG/VmOkSyUQuz2j+CogXGiP++7/O7WqrzYS+m/TABo/gDD4m
ND31CZC4RbGQXWEMzKQG0fvOZZqJen9Xp0gawrKg7zCtTNhopdnEqePWBMcP7b7j
n6OItQG9vdWV+YoY5LhPSYw6RZAlGYIyFQRkK4SPbxfiQQR4JSMop5Za3ArbXq+a
BaRf4pLPNxSxp4BhWETZHyjlCe7rWKpzX5xxmcevIuMNW+9fQDRvOhtO861pG36z
XbfgS4ymme8IcFZ/L0v1OriUnbvynNCsewjpIuaLqSMyCKRpRwjVBKvhnTPyGhr0
vaMrMY3cWfAOt7WnRPVgrxeEMGvmDAnumH1NLlCwP8U2Q4Ic68dh86VmytMN6VKf
FCofC1QZVoZMs94AR2vZ/4deZEUI/NvCWgjKLVMABgR8zdOd4bpDQjxvur/NMacE
rYv9iZKTV+PWI37n30qgAyggJxxLH3AGYxfxnVocofvWq0yBAZsoKjxef7Upavwl
ZBsj1MOh5OpG4vY9gaImydg15tKuF4x6JdvLQjI4Irr72PJ8dGuTKPOpSe2bSraZ
5UU5PXmKdCAR3JeG0jpC3fW62xDXHT0fWqlPt3NCGxpRCwuRmXkfg5apb4fWl2ut
61fJxBvjPS/WsH2/vqs3w8/z8lcEiwjHFEruDrSkZT3PiopGaWn84k8NgR1ebrqB
k6h4/kVjXSKhXoSdeZ0crW1Q/3VO/DRcSMVXJOZGHPcoA17wuHmhgt9bKKSxZ3X0
4IYBg2TCERvn2jKBUFVGLTWfmWMVMKFlEQCOVu4E2V7XWYEm/zw+oDNQB/Gm4bn3
5knCqTIvvY9golgb8NtMdh3ifClWMpjXHJBpQrFA005TDmdoFwv0A/+mt7hmgb8f
6FEIZGyCCrAWe1/CKUk/SczGbdfgrxlFY4/jGCS6fAx45M7NHznJZIEcbdHg1Dby
wkiuKKcbTkOH+5JKR0qqx2MeukuyEN0+2lpTqdh73fP5PT7isukEoGx1oqcgFLpc
N2L7z2r0Phx+CO/W0qAPv9jJhhtN4zcos8o8zWPcR43NaZjqY8FVPcf9Uz6W3rb1
qlMq6v9+mwfVduQK3Chaa/AhD2MUPR7mSyFLtWn5wyolKFGDn2JKMiaUVl7kWsQ+
0gV5mpJDh/aAT9y20gwM4UfddzO5C/XvHdcGFFbbcfScYe5tt3DsJd/75tochlIt
jPd+rmKoVX0xScXAUhxLryje4VFOycqSVxem4L1mvy611QfE1xfYbvY9bFI0lY/4
QZ28Dc/M1O9lGwwi6kGzIMotiWpZwyDIhVZg+ualnDWsgZVOdOviGX+aBwFuNcd7
JO+fHJ61HvQXlaKWxt8yLinWjuPdytbQ6iHQ9IpZveh75yRgxYDi79gFxytf46yM
TSpwkg43Hobrpy01ny1wqQbbZaYI8lYr48Er63Pjopd9Rw48jlaZPsNq/N8nFA2G
Kh6EuQIoUPYLQIwCmBuwlpn/xk/zk9FycB8yAEEJwfwY7JQSEBb27MXUxQr4QlHm
5N1qJ51zmlOL+arnzgqEW3IM3LRwJ5ZGB+u0KvYzwY6/OFkIYUB7hEiRdrPmS7wp
4JDXGywQ29o0aGVfmxVjiwmjEydfOsEtTKhhLG7ySJPxnhs0oY2IyMSWHF7LLC/E
UKXHSQ+sDEyFBLAWWJ0AQXfuPSwEbreMXedobwwjykPLR9cTTDMWjQkSkZWQVFVI
dIXBVeNRzny+oNl0sVyt0E5SUVmr/4oNNDHQY+C6j71fy3KUrEO83e/I9nTVEPC2
xALoNPQkGs9MlNygURMONVgc58i5ht/vc3Ot02LFmhTZKsi/kJgKr1nMdlEbYYuu
hszX1m5BK2zq/lRvhTdvruiT44MNoVZEBWKDwvH6F25rFNkhtAkVKq6CGW2miy/K
aCs63Rp8Bs0zrCZAdqGBSDnUmB0lR9uUSnufIbNdJUnkm6/mtNF9Rn8nYqgPMs05
PwmFyL1STfdrZOoWtoSleqeA0wOco1ucdkPJgTrEtY4fyesOBOVs7I888Bh17wuP
9CYbF5MDVJnJGEnUXUt0PAp4sF1b+TqVDKzH6USvI+EPecEPcmpTK2Ryg6Adw++O
P9VmuYxJjA5pXKNGBBw3FYegaaXVd2Z/HBhD/Oi50oHhv89RALTJWIS4AROiK827
b2DEpQ+JeHXsWnYmL4+9B4MuezrUdCdZcty02SXwfjvnsBG/JzrcS88Mwv/v/Sz/
FNO2b+L5Q1Txn0jJkQth5y2eSivRiymPoRdABCDSDNgeAZ8vEaDApFK06RiRTXQN
gNFDwbjqSzKR5pHBC0TeCrE5+CFfDya86DKmljRL5pObwA6kDJPvpeUmBuAeQA8E
5eFE4tmckqeKGRh2vyBQ1aEmlPr0XFpz9DBgvLN7KZz8y/vRSar0Be5Dp/MiiGmh
NGO5Koa8wlDvq3g5XV2HkaRdXAmSGw5QUWDDRJ8/UB0OlqiDaQ1tRyu1EZfMu12t
x3qBqcS0qmSgXZGtjj7tY6Uig1hcd9d322eDRVx4/HrQAvrcrCGRvDIfyHxZYc9z
WtI/CVPyALtOjO/8rTnmYXogeEK/U6I+E8XpL9uamkT0AJYdYlTStCEpAfUN1A5a
aZakBcyUtwaePrNJHvfu+iSPVaaO3nPHR3fLpdKUEam5zE7q1JBKS70BYF2+e+5M
dkfbIGUr+C2JuRtoOLhRoJXzN0C3G8K1dutZla5i50Idq1GN0IYeu0IHRR4Qbs4s
fw1EVDKVmk8VsyIxziY6sRXUeBnm1bGt5Tlgd0i3aXrljQ2O4d02tWWS9B5azOKX
DrIsh3Db0NOT3YK6XzkUlPPPTGMvTDzSa12doqt9nhp7nFtVZax8pSYZ4BY0wS5y
5epLZajWm9p3pp4Gptgi5rr9n4i1uCGLty7buzH8IBlou/UWLIt7OkxlYwWQHtgz
fMtX/Mo4memfJJd3Z3VbrvmCSkraunqk6pzEhrH8UioRsBl7i/So0BiwSNXvy6HL
LaYCX/vGN8LN8SS3eZn+LVVEQJuda/+H8NZbiyacf56hwJLxFVS93tzbMFafh6r1
PS+a7JDfby6eW2meUGXR7cR8nGg8L8/lY5nXFERID/zDRUJahYH3owJvfzK8HpmE
CvqeUp7F1MUkdA/ZIdKB3Dt2bHYJPDxqoPlHvUA9BeFDGgRIUNv7C4HC41DlsqaN
0gArxXbbO2y/f2kQq285FRyxA/l1WXLQgtkiYLNqXdipSNkUB8iDdVMw07PyE3iU
sZptaNrqbviUwmtkXxIW4w4hYsy+3IbbzFL4Tyk8b5Af5gA1XzmTOTs/qce2m0TD
bQeKV8dKNts5pgL1yk01I62dBZy4idKkb51ua3td4rhxRg+zIAmoJLPyBYOsn4Q5
8z7GMX6I6X0oHx4eYmLgkUasSsB0iMZy3IWzJxWl655AYt0ZDRaHseadYApZQP2e
kct5lTu0rJPghR5HEYdN+M4quylFCcghfKrZScar36uRtxUeiUSB4Ao6XHvQEjYR
+OrtCp2Trj/R7T9MdZU5ahMurmXGMX1HsYXKDu9NTX8fvQZTq6HxrZpXEUdoZn8X
pgq7vYLgIoXWFdrKPGdwxCIWRcMbb1rU1NoT8ElX+vu3y/rNAyg1pi5ieogKiX8J
JSdxZmTudIKHzQC1CFUzAZI3n8kvt1JE8dl5hy2Lrteuo0HNlrTVbiwD9nQmaeLH
lS0ht3VBBDaipIrgHPO9gpRGB/oQj5+pu2dO2aKVH2FGLLO8QhOXiw4gr0rn53Ty
bmyIHDQsfKjyOJ2ampzjg8iNWkjs5SUzlAqDNLsVxqkrDGp9RXzKGry74O+RgM6I
jsiSAj7kAD2LFghN0Vg5OKvLCHxOTsVVLNnEf6rIYn/M2s+mu6Hni152BW5uJbmD
Ga66rEIg3v2mtYq4bHd4Rd2V2LWcnKC0YKqDxYG/dorNn22KLCx4YfY+pgh7QfjM
6IJpKj6mPyvq5hSr3O++7FvWcBXXsn+ZvGR0gfxvqWFmUYd/1xeppXCCXBc6UqfX
gM6gMADLRLr7zLuwiF5xo4IXAwojPK7owrDV0Nfwykl3CCgV5DuYamnOOePKw1Ut
2fjbWO8xxvIseHha6TPMWWe7X8de8FneVgHZoWrZjUbDm6Gc7O/YfBwY98Adf2j7
C9OKj19SXghU2JmsVrWLq+sOme+RzlsJsm8hW+JY6UxOYfRYgNnIfiTw1/QVMkcT
yHjEjfCaAvjQC7xKytHP3V1Ul5nqbbvXWMTEjXtPgqdQ5LuYgLY2DilipebgSInR
4LL9GlzIYOgKPszbn8pV7T06L8uI4OxDUkh+rldzEW2+shMgfhJmrl8wXxU+z+iL
vTACLpN74L6gMR7LvwBBJegaK/VJLBAvpNshDDMZbud71JilnPU5IPEClijxVkZw
sz3n2y+pDbp230HjTcHjLModlrmdb/Az0IwCOhL01gDHMQPx7cTay0ksOi0LXBHK
yHWezszk37B+HU18G8mrQQ4B+n6CwFNgBSJ4VQZoSQnXvmiYLwinoT1Sj0LWkRrm
3Mi/iNh9t2V7nGg0BVC/HKN5edv06ypayJfadISv30A+coX8GSpatyWQDsdh1qNy
Q6sHOnNtijSoBltw/3bvqYKSGCruGKaRT0j3rxphiSPVFx/hyWSsxCvtLhWM3ScN
fMniVoEah4FgJEbRpgNPgvO5F2f5v/cu5Ey+u/gvA1LRTtDDs5yajUrMsA9Ql8m7
V5ipHuUypB4/V9QWIAJHVn+gu/POdFIq+0zkqWvrjMRdAP3SEvoHyeeAVynZKkb6
Im6BmTE8WR5u8f7/a7cxtY5KxjaMgtKRjHQzQror/MeBt06eQo46lqJasHR0v4Bk
va01ZR83iHpIK+6FyvQdzWxCPIuZjxAVqAjLGFf06bDWbZg8pqNTIZ7h366kdsBF
6K3ZoYgw8puY7kVJ/QdemGn3AWRMQVloKdU1MG7WuTewM1ZedvMW9PSnVS4vVc60
Z26n1V4DeZwEcp/yVFOrR0z0sZpEInK7UleZJ7j1+VEV5TvdrGdPNGd0o1HYgZ2R
e3vwy+NPABU0Kwko37ZLPiEmKPvuvpMMU8KjINPwMVjh4ynzbdd5C1wB245hpE4/
5iGqxb7sbzI+5CSfPOiqFHvKc8yVLQVRiCsWoJKeDJxIGcqU8rHGg2IMSrAmSMwK
z58YSunrtSVVjuo90ase4MBSGvud0zh/CPVDFwT+Djs9i4//wagrrNRAox0xpgg/
miQqVfwv52xuBNa3/r27DxORkS/UsLfD+danV4KfM53ZORfpA+s9S7Eja1oxYnFy
ZxrTPRWwW3BOE5uS/37onoOSI2Pm1w1CgfB/IDEZNccCCMCDLxaQKrObdIsAnmq9
4bulgrDIMNSntZPlZt8DWO+lHDXxT/BL+voNCLCccKQAuXtqg8yxPvlcUuYn7s89
NzmfMhTzAq9DBEXUR1KWOk/yaSbrvjYGCh4BjlhtMeaoNW/gWFVZTUYC9aNxkkig
MGgaoF9fcKRMUwnzXoYsKu+nsasP9Vp+YWFxNzDWMG90Cq6rgkCqZ/M82+bCfN8D
CbpXQrnJhbWKv/ZQRgbHJqoiBV8RRikvKqxhBHChUbryURblABxRw0t3EsaQrXN6
lPylp2j2QhwGsoJodGfu+U+HLktlPLKWDPDWdnxb+oTC57RpT/2N5RyaQqcio9Hb
eMPCjOjItnch89bs9gX11SDTICWp8tHwgpan5FTX5UrQbo2WMio6xZkhNmQG1vmp
Po8HSON3rHZBDgjYjZ123T7uKKK+DTmWIPp+lVfZC3bXEBFzpt5ZwnVfqVnAoZeK
PTspRrGDxAtv0tntBEkpwLazXvy3KVAivK1RXBLI7XIfPD9pZYN/jvMXSFI6v1cy
Krl6a1wEaSzgUKiAm0mai4rBiDO3aRcoMsn4G9JvTUehPqUGT9K8EgNkf2jLXAx3
KnYxilbn2kBGorXosJUGU1mAxEH67bjAXH/XntkVwbkIRVdfxle7nlrUJCsQbdm8
iXEdOAVsefn6b9yGJOC8SszDrG9dZ0KiphqK2RupUwa0gw++oEDnzb9mfZhcvUiF
Y9RdQwQ5PiVn8lFUDVlGtf88Oh4rmPd+416RX9PvfH/HyfP9ZPljnGcQD8n42mGO
v3jrIanzls0+W7Kw2p8oTX0x95+4VJgY1e8PBsBEq799Kpss6x9tVecjokRwAV6K
4yEpffYQ6ClalgfDcAXe2MLTW1nnxR4bRwbf/foWQYE5mg0rT5QcmKh3dJR42Rwr
9UXNcPMQHeJCK5tC6IrkVQjtcloclR+gbegCRrEq/gDrqyhIcsBXUQJLwdkYYdlS
zihFdO7AaTQy/NTpBUv4wpXhOCqgVzw2lfqnNdVrrxk1kmaXvydcYQ5H8G5zRHiY
4BcC5xhhFA4DdhMYkjvetps6JqJItyYSmDOqX6WrmQR2l3kclHddGew7hkN+P5+c
jLsmxYIm7RsesnTwssn9GFdE5ta9F0awgMgdhAnNR1jR3nhzEPgnkQ3NTrj8Mnnt
avIx0dN5awV+FBAQuLYQa+TV1Vz0gr8LAt7O1G3wUpm13xMfUUVPSPpnHihYiXRi
3864ZBt0VQAL1uolUDwdG2sX/N+itb3O2jOVq25X2L80zjC5d/umGWDT/Z0I4geM
J+gq/Y36/PMvR79ug5cn42peoV1rElbIdOas0R0o/AQk4arS7F7/UQMuEc9u5CKo
bSdMNSQj17xRnDbjs2uNexzUpCqYJm3ZMnCvozpO+78YeFnnW9bGzo5/7BizxHP3
w4MWnrm+0zkDyWNod/WG5oCLTRqZjhGJUw173yKA1XVXahx6ypJuh+RmfZ8f2gTY
hDPkd+VU/AsPMP1cC8adNQvuDjn2MxkZ1+pBnTWVFBGwVtqB0F5T5HrrYjfyS27+
tZSADrq3vDotzfMi0jQLWbtvgSlL8Uy75gAlkm5/lJ40SxgdoDaEK2TSyijkFCph
6BoUJDZlVYuU9BM+iBw3IfYwjtZfq0Wnyqx31fSSdyD0RPLjRzuitHl+RVgQhnO8
4XIcJz71mvLkevl0PsILC55cn8VWnF05KGIBz8FYh0xhCqFXKrtbgYmOBWjIAKdX
mWlHecNuP0au4warH23nI8DrxYqTdH8VHMeWmKWhtg8qi9nlIgHOqkRpy7Z1PW80
ba3bVmWxSFMJzAU3uieDxTWCueOzBCWiAi7O5rVhHSDOU0wPkguUif6Hc4aFJeRi
OLPYC4GMXaaxL9iYEX0uGq/5Vsk7ibT88YLTO38sujAjAWu3hHiRorUI6lMe9cvd
FaIW7k9uQSX7NFNHzl8zp/TBUoOk2DkfQ0by2LHm1tc72bNJfmuhtF3DK47fHTIb
o3pbQkigZ+HwV1YGGVWItt9SR+PfIE8P1q2FzxIEIZDZJbmtwqz9ESFshl+NEG2s
ro3i3jc8KM6+FNpKfE0KX39NAc1+7Z0Xye71MjLGAD9NhLQgP8Nx4Qh8v44WSQb7
HjMtabHkTd4eNbxEj7sYbcjCn+VUSE7eG+EpSmqe1Eh96kJlGGAVVyAbXNQ3vKeH
GgOQHLkJs9ACmDZVibbCdiNoG9Lm+yastvFNSe481y5OZH28Qn4Fynf0cAVvjv4v
oQugc/mLXxMhfNEsN7qJkNWCsh4o3VdmT0BH3gEQOE0CeZ1WxSXjS8N/XZEbpOeL
XJ+G2v7KSP304iq3DTn6J1r/vWvxfWeDdCsAl/RGDhzbNLHPaCfeAmgg6p9EWrID
Uiq2IacP1LUMe6r0jqMkQjyDR5YSs0RuXeyjWkMuZ1P9ysbJ8vML6P62Mv+PVRHh
Fb4ScEsmESw7gVWM3F9l1vutsXZ2DXtLGvy0P+myJFCir6r06nNFsxYIXuJXtY+c
NXSdWhRMsDCHqrk87GVwGZE+d1i7E6/5Jos86bSby42s+DVVFUGNOkbC0eoDni95
TC6Y9b6I0bYcfDHupOV1QrC03XsX/X1LwJsGGNXjs+LJ1AX2XtA+2Wv5InfdtUJX
r7GhN+Ak3io4WK7X2yOs8NZtl6o5oN/Daeu/2afkDMijnyj+W/fOJgIxPdXLBE9U
Qi9eESoKhKz1RbDfJ2WIpG6QGyxJGP7iqw0stCL01LZcj/9AlmCd2ALCaCTdtwUH
9iWAFFTklEyLS+VvOYiMFDK/uas4//mjz4YidO880KGBG+irT+cjN6DkJKwBB75x
y2kowNtjGDLhOSLd5AV/aFIzLrzs/SJ/ksJnhaXrtGrWXTG4v5b5wRBN7aomWck2
j2sb4lmtsFcUMsTpKHbzA4XjkfCw9hAst6ZXZijWVUyHncur+txVofPXOlAahU06
VPjIY0vvVyw3Vp15E27DgfbsD5jEuRMv2M7U+KsdHNeCrBYJqRst14or40k+8OcU
jMHJmvDcOaDMJ2NZrEAbYRdIyVD3DTqwPr3Dnewlj9GbVaTFjNP5cy1ujW06Ahdb
InWLAFhd3IgJ0jLUdHkBukw+AwVv3lFxTXzW8T5Jm/uDNUqNblg96aFpEnNqsSoJ
wluNfUDnRIzjq8ESp/u0sG9pvLs20tPn3MR4GHUcDynoZUiL0GRcQkpX3FrVMSSP
3NQbsmH4Zve6bhLhuelAuHo4xaE1uDfrXVWUFkarvX8iioGNiJqGuZ2ONLU4G/4s
fmlbE0rkd6AVSdR73wf8iSjFcspADgI3A1IbCTsqOyagc967SQoQfAiu+GffsHfZ
cDLAcIR8mkcpHGrVPsFgB+yLqpyfwrT2rNfskmGc4YVVewJpXzwK8LbCk6CWdNzJ
o47aF7V3iEVV7g2rZ3Isex5oKZvi02r68rYr6xFVpucfHC8cnLGFGz5bfkU99rgy
vqfxk0YjQ1oSRavkVXopejIJJN6QIMOi1HXWbnNjZIw1oKzCbMvYHC2LB1NFCpjq
CbsgHBk/D0BclpopZPfL03Bv4yKkfpXzfrnc2fgxRrDU6qSYNB86SxNo+7w8z3fN
q4whfodQSydFYf80P0Mtzmuh/VPwRbQk2GPVdORbkLizOEpFb0ZFoVMEWtb8FPY6
Okry+lnCmgka6am/hRrGwHfE6BjHXzl1Nb1kNwXyMKgZ6lcpiO4dVsAUqhKZqqlZ
apWOaAz0/qFI6N9MB3xPf30nTXaYQBcqyB16FadI8oSVwBnT4CafKrhV8P+z9YKb
4O/VpG1j/uVFHZtOwfLON+qoD9ggwSLpHiprRwLOuOGb+NiJTpEmimj484dWvx5U
+wwoK4ilrZbmu6SxtkB4ZDQV/Qdf8Vz4XxlNf1gyW9kr6ujaDqQurpTHNKT20Lmx
d4wGL4qtbJKJEzihuZABrW/u5iAL8ZXG+RYAkkfs/7CeCF1sGc09Z+2z0OP4yYu2
SWHrkDImFwkM1kG8clM0AlcrGCbmkTZ5fH1dPLa4wHQWirq9p7KqxS+e8n3chW7g
0osqrpZ/18CvLDUhVnQgvEGA+j4uO4UP8uiiVaNI6N9+F1oQ9p6D2XaOg/SDLx2W
MF9zhHXWMe/n+c+mvN7+s/+6anABmo4ygy8rCzhtsts6upBm1toAwLwXLeH6pAOI
iwge9vkWG3Q/Opj8R7I4ftlKIzJAZ60djX3oN7PHto4In4wUZkyCTjoCQ0wdqpPV
1txn43JqK2yNg1dgSe0YdekvRXHKUAke8msXlHvrbr14t2aPh/qlhkgg8nq1XJAR
N2ARVWmevdrokBYodMRU8KuWvjWch8+95UBaTgtr2dvWFBg4j8Os0rCvAoV4giou
jdqKULJD0gbixZrMEuIbEy2iieyFl4+n/6wGPnCdyGZ0hGEL4cOjMe//RdrI1Gof
edfTWJcG5ObLlMJ8zODpkhS8zw08/5NcR8paLs9KJz5XGmdblTvYW05T4qYt7ugj
ww/csBtaG5av1SaldP/TCNSxrt15Ej5C9qgKUvhI/GR1k+NlCzRxVzSPHPLmQX0x
rQgushFY7BvP17Dk5OA336FrPOvQiu2pVmgTCzjtg3HhxLgyS8PCwWhq7l1pLXJr
vp8+iaeSw/UkdJsWqGZGo4vsMiFaStJiCRd5/yZ17ytyAL4oDKX8b8wFkdt7o0QN
EuVzqGUvWM3S3Cg18uaN3/ci6paCnBIUF2UQGidcXIzTG/mibgAdIAArqet4sgfE
zxfPrjuWJqwO1lXtUm9ApF06gRqnTpw+BnFecGNv3LIZfynEKRpfgEEUAzxXrOHc
SAGUjV78iRPtaYv9VVfX4ZG4GzRSg81WBI3buumnuM8PH5t6xs/Zp15uPob1Ih52
l66Jp5rTXCTKPI8hUmYJYmL07BDlY/3PnR9ZnOKZOnTKG1OYDAE5DS3bUTJihD3d
WdLGxBQtOrzdSC6Inoi4bJ1W5Y0WQf34RmNb/5lSH7xogpQDO2D067WWA1kTdTJO
wubzhP1BceRAglbWwrV2Guk+/3ldzrIRkXysJ22iKO8REHlGc1xqDNOcvdNYW4gV
Mmw2Dm2zc0nbED+WnOXZx2H+nzhvUN/vqeKIt8dlEr+AM4aALYIujzI/b+KoGmPY
jImZ+bDj4BC4Mhho0Z6U4zxI29RIjptnWSbTgymKA/O8zmAMhf1AF4MhqWZe/jF5
Rk4IIEn8BuHjOwnJImMz55xM4km7g7sGG3Gw2bKUojJyz/Ry/faudJgJk5YCF45g
d7g5DzjSkX4GMSNmCkrVjbQxoGVSFwSjj/hgsN8B/iI14PNjQ56DCmGkopnQ75+X
XVE39E4r8tj0KQvfhGojpKvzgDjUIy3qxxgz1bUCzhrhWEoGEKoazsg85O4CIeRf
FjlapY9bIeiRL2iIE1LqTSq6G6bv558xdeDUzxSGUpXjcTcOsweENqyVNVVyIHeM
7Gg4jv7Onk8hX2ge+uk1x5ewCSYiU8QDKdjbScfYbAwvgpzcKB1RUbc1nupuL7eP
kdaL76yWa1KdsOWt2zcaGVu7KGTN24HaWuruzPtKKtTXuFPwlm+Aoe6AdcKzdk/m
e6Gne9dkM+PmJ0Ldp4mN/OOag2gEtSR3P9W8MxzwiQ2R/SbWLEMWVaxd5mUp9cul
g/GpTnm5YSxiYhnJdrDeaIZ6QpBWEURHLvpLeoEtOZhc0myf9Btj7mWBmy0GqZpF
tgt+Iacpbv1ysmlQEJ/w+wkiju15IOQsbFhCjpz9x26P1+jx9KUVUWXVJD9d2RA6
f/nTMC6+iRxlGmFjqS3Q7st0gMULCxMKPg7GJ1DCKIxgsQIBDp3bCGM08xzdjHgH
HJ3DN7NexgUjBEffB4lsXjetAE5I8eX2WLNqaBWnYHgoBIla1xe/T2pEoVT5m2rH
bYaz7Fz5FDqX8/jfzqKbYlhBUy7peKGipONVT/WxGlONaBBHiNtPuvt+kusj5TAW
R02/1p4VrpArfztGqktP0+oIKp1hHxlbMRewpibR7bPPn18wNRBAm1Qd7jlqg7HJ
rT6Aja+vrzpOksBHnNL7w3SNJy+2qAOL25u2Kpx4www83z5DElzus1Y3As7F04zE
EdrSltJpasHNlor8XheQ5F0OOA2XSswKd+PoTmsbS0kswE+4cRGmdpXdodS1+t70
a8GDZfFSvELgGv20W2Z0YoAcEjC2/fhBY3qqmoQkUlfXmt60I4jcM3ZIjNAe8PER
Y6OmnPf8KU64Gqgulyiqc8Fqx/lkVDd+53TuBee4tFhVoJ1aA3beOI5Os978D0Dx
ZQnuXv51IVy6y5OwZvQ97rzqc8ZOwZ116EUxdpWT2iuoAz4Xmrsc7w3vNc55VKCB
AiI4r8f2UbOtfmBiA1nazENbOoz3VPoLZ5okBNgNkOftpN9JORbuhm3GlHevD8zI
pZ3gdOTXtlETJ+G8Sjoslk5rB4TNLpUzsdA4c30Dd2zxVEaTgb5XQkQafohEh79z
ThEKaIkSnApB8zlzoYXVuzJqkO4YAFl7Sx0lyTfmzxSnym4iESmYaxeotVG3w7LC
2gPLwTZF6PH/ZrUCRrpfw3n/Hzeoin4hJ3sbq+b0kStosYnbja3iWl9stmn+CXKH
1wV8N0//NkD9C0uQPvA/cmjmgYo6WNidRxfj6rz1RzrXdKHLypCsRwCVbZhDMpR/
aJk9D6c1ufiKDKJ81VT9wfyC7kNo5u5Z/nkzbA3uEhw3EpxfJ4n04OoHECPeaDqp
Uh8q0QaQszBIpLpyRTpbdgeDAZdFmOcPfpXTSHq2Ufe2FxLyA+UPDxhOwSqVkco6
eAfFXQ2XBgV1f3uIt0toWml2B7UzPkwN4WhGwy16//DzCR9ezBl1owU/ytMmQXsS
9NRlag4YINpBjGII1ZhvxpaEwhenaRnrHPVPtd9hH6i0kNotGlu9vGnT7XzUIAZV
u+crALsublmEQ5NNSCfuRpPar2coTLmfbYv68oH23ij1YtmNd3RUYZ61+73+uT0L
6Nm4CxolfOPymJ+/URj6kLuaNI09QG5bjxGHX+N23eNyqTNlF0f30IYjwFzE72tC
aWlXTrriXX4RlGCPR3MXZlMtnU6NrVjt97Zg+JEqpIl5NnHbfoOKcFIRcNPz+f8o
fmwWdM3BB/Ld/sdJBWG5kHD1gW15r/36UL3/8XXHtntvmy1y72obI3Hesf4nDCI9
YHyzIBnTsxOU3XEYpyioHbIvsGqEW3Zhr/mGffPn4tAcbt3MJ0dlwYNIaSeCm6wY
DOytMZ/GtGmFqOTHlVCcRj1JqPTIgz8cntzfIt5yNLraWTDOd9ITtMosbjumQAfV
IU5dVJOI6oxqDm1zmluU9ky4VmYJ+aeTugDo1nl4v91MXbFmfwB+rs66sPaNiMp6
v2D+OHHlareErH3cu1row2nTQxi+UUfKtpmIPH3YYgcTl2BPG0P8wjGhDxdV9B6Q
8MPV89PjrMp56LorZMeL7/5YLv6IFH9XE+KT0woWkdKJPy4K/r8QSZo0x4kLa+3p
bRF1uF7OcAjIljJvh+N7feJd7Hyj9o5yiKStdhPKF0d92BpCRlROIx7cwW+YKk/z
JuF3mHLMjOjaLGCheeooQbOG2hKEHHgyiDGLmuOt32msNvbNrdtNz3DeIU9MdU8G
BPAtgLNPTQyR20/hYGDzXoVfFRpx467Ye0OWRe9/N/rdg8QxGT3YCRpJdskrGCkG
JvvVe8mYba1FcIs1EYEDovcCmdm77eG0yw/EFT9oayLfTk7y7CEt8RDjuz4L8h+t
C3uy392wUJxovydFIEHG60grStMvwqIAFwpbkBsoafjZr68vWdzOY8qQj9wLAAd5
Y6VUGBjhMMFQjkQpZmxcznwDixyQcgb5ep39xt+BJ8qWI+mnYk4ZreESSfSbgxjh
EtNLTy5nTBmvntYXaiiLHLkLOg4l8difNYgENB6m0CDHhlSTqYKja5gRQZ4F7vR+
ufcz8n1EAgk81+vRl4Ymj4w+IF5q7wPFgWC++PcMUG3sPdLqqMIugmcGKynwK8wM
rsRxgpp7PtfGad2YvIGnJ6e6vrUMkye+Wmpba/A3AGUYHHl5Jotf0a9IJZtHDSn0
SzcA+7nuzxImMd8Z+ddXngDexIu00eZehgURw2lV0fKVCijW2aDc9zraLlp2AxyZ
FNrDt2k0U69G5RrJqqCUhhTUWqPGDGi7irObz/QXi2KsPamkRlhM08QGsWEmSs49
nfFlxsvGPCtnz5OzF5WXbmdm41s491c7lk3MLPelFwZkqpSU5olfP3vg8ZdHfdPn
x+tiFdE98DZVc5BmksPg8GDNmAIP4tcVUlePKQeNXsH+fRGCJys/5pRBmW8qJnw3
T8h0HuvOlNUcTYYcQrdLWew5m5xnx0qKlebP/MT+JPNCcfR8tpkX6NtlKGGhWvSM
g1qJvHEmw1yS/PB4Y7kE3j14vmj9PpvcqEQIj+7jqk03hj0DGCYn83D/y8R3Y3CL
ykeQ3zdGvCshZ9h8mfvgI3uNDbGEMyiKZ3dCTbsBWLaJI9bjSk65B5a37pq46D3e
Gtq43R2OaePn8y49tPuEOUoFc6Drg1R++d7BGhz3M3rzjAWG/URpAqhx1yrwWVSj
LcxgatkDyFdynnzpmYstXGjwxNnpC1B1PgSFQ179528d/Zg1NKSkNk5N2RV/Puvp
ym2v0LF4R5pJLGTzbGFo05QgRYzVpj1rbjHZVJa2KGW3wFf6R6WGWlFARzr5DgSw
NlLSokash99yO0MlAi1vvVbf5wu8Vv4+72JW1g0M4V57C5KMr6fXIrndTkAwgtvA
YjrTqeZ4hNNTWG3u/kvgGuv6GsnWHC4sudazZgOA7NYkCb6FHwJv9hLY9zpD2LHI
6TnrnKe/ZnFK9cp8ZZvbX4+n+ArFgCkXkGNlVOUJShmWHxsOgjWjJTYLUo0HZsoe
U1X8VGFBDxISfgV9+8+GVaf/9/mmYBoLaX6HP32OfYoWtN7PQkv42QtKw4WMAEzJ
1EfX9HNPurjBJtaU5E74Yiw6BxeKYEDC23sZLkZAawLKH6wp2LdNt4DiL8LUG2AU
Awn8rzcVYKZ0wFPBRhyg3Q7vgUV/P9xuitqfpqFW4wfI+7Mf5t/kNzFOFLxMVO7b
9qRnYw1gpqb9yMlDnQrXIATNHCl66RzL+LLXuGO5uABfGCXJGXjYia4ro8PilmFl
kUzprRUMNe/mzJORtLCGpjdX38DPNL1F/JpSL3vWUSxh9kU/rEu3fwyxjDRmE9NI
KEJmWbCSZz6gEeoqP1/m2BhGMsqRlqp11IsmAcc5Zgtm8fcS3uplX4ze95SgIk5c
72fhbxR2+0YCriOLhONyRU3U+OpT1SVreQgebmPFi+3maWP/fQW1ldclufzPL0M7
f6Tm7uFpR3a6Cu2oL+G2r7OKLX6FPT7TOFYfGP2Z6BVJKqVDyJT/kXWFAjlShBYg
/NYPuZo/cPY6WlhFsCl86DQCuMKF8Dac/u41Um7JJWol7LwcZPqIvEstQRr/hZNr
wDo09/Q3P6zU9mmAfXw7lYMRuasH8i7PfnbSiapk0u4KxA0HzMghTNp/Rw4cObiP
6WxV3PrYy/9D523Wb4wREIZIC6y8wcL7IveBhYQ0zPtxO87liP+dSJnjkH7qF6be
7qPP8I7ckcJRWbqzj2KNR2WplQs0EqEqikIq3CZMbeT2iv9p6crljrPYvsuLBDg3
eIzwffbckxWZtxl9RQlDSqdQHc7MXI0LQKhf8dJnBsPm850BwogiGd2TL/wSVZmh
IKgCsoAGTArFRBoKEiiH/z15CHytDHxErCrMUsPfXWGFzW3QSkRsSELeWy5bFEKM
t744a4xavpysHzfsjAJ4LYq5X7/WScdCrJL1F62o4I4Hue0YL1miyoC11iPS/tW8
mBtaQQgoTm12BnD4Z/a+qjI8G0zuTU3nkpJuFMQPT7bJTl0f/qms8YjFpofjlZ5F
LJmrEb4Wqakp4tc7PlmMMyjBE80lecMGolH5fJlqhK7FAAi6NnYPjqHFIZI5aLUa
yo4aQ1/VDR98hO73Lx3RoU1YEIuEJnt6aM/x/g8fK7tqT0HBX/Yk9jktmVgw4x/h
j4jOC69Deyz25Aa4GiBOSnqFFsHG6m84lbJRY4X6Nz4SzeDPrRo9TJlMFqHrbmdy
DBKs7oNMEKOrenQ1N6NfKcjxfV8g1/w686uGe3Ttym3Y5L/X+uftoZmV2/PWJ6ab
JMNcgAWXYDRLyvKvQ3MjjIOl3oWkq2BesrQHb3tcVg+GdJUSghWRuxUGXqMrymGn
Qw8e7s/TxDBUoP3uKxN+SuctseBiyV4PqVJaIlpqYoPAO9LjbnI3BIvEKbMYX3kh
FFie+3+sN87Hn/M3OlN1hgVhfk2MyxjSx3aierSfornOu2mNnTjtF9yg7I3zqvyR
40DK1A6iXBlT0VzkKQD6hcx43Jpk3DAFLbPUsVI3IqX+CPNZqDGt9VN1g8wetaWe
TMjTelOKhMhcYKJ7fcrWK4nI8bVo32cJL6hXcdyEU2y/rBzEsWCXAJ6gYnNMfD12
x+yAEB9fncgVIIhKRY7cj3dPw4LEkHwT6NrSp0zT7dY5XpP6qvjze8iPD/HPKH/n
Y/VooZSpjIiwEbcezBd20NBhpRQJtJEzqaXFNK39qkVZd/XSb1XRUGzikidFkxG8
6QI/RuffLhsFIxR9EpJw8u0n+d6NxIl7Nw7r4TeL9G9sq9Im1jG6DjOtGs2KBSDR
6Hc3BmVx85bPmnMj4L4aCZ73Q5AvnWzR/edcWdi+/dSjtkBXjyc4u638xMm+CNJE
K2h0NlHTOcrNEfst/d0zJYuItYLjPNslRVGR8Do7GF9VMlFzzj+wJyCSNQLSKLPG
4d4wUPmvTlXiQb9H+xyv/ab0KtkpSIYsfQSkG75JRHrpVfcL+1C9frEYj0Cd92PP
BmCee1ENVsYTkzt4sfWWTUlzeDBRF6yO2j6oQ+cULrPzXqxqiRo1coRKkci3i11z
0LSRfGNUgsNkAmHaWBX8/DFgKKsGnnl18VDviJZVU13BSu9hBDQ+f5HhHtJwsvwW
u9nOFwjZKhnNG/CETzhIa+jVyumI3fXjqCmN5JUSLF9M8KtyfwA7dfLWgXBf97yr
J6S5LKzSy6rP7JGog8uJ5efgi/3KHShZYULohqYI1NmOKCPJg8LeUMMyB9bxT5Uu
NNFs20um5EPsXx+6nwvjeZV5Wef0uveYjeRTQ7arwGQrDXz0zE+x62LW+fOsW1E8
+jNbg6GAZDPAPcz57m685AfrZe6ihCvrUEbTppprPan84sx3XaxZwLg1LWpj1fJ6
zm1LqXrV7dmwcjgw9Nyha4eUHaK/ch+GzYXRKSRGjrfK0784xWerpK/LvoVFiMD4
cnvPtymP4X+pE/0lCGZN/Z4Xg5EgN3y469R+LI2ek+EShUMlzDIUqVfXSEAenaeE
WdyIpNvET/6BgCw9X2SJc6+FW2l7CraLL+4NqGBD7Iu0Dg0AQIFiH6gCC8QbiwyN
dk0VxCvRRDaIBf9DNpvUQ1ELbxKtQJC001vZ9a2Uzolj3TWoDaCBWsUI8g0MIHvm
L0Yl9hRTAYey3mR1/VycRkN5e1SNx6qmtqBKfAhYdQ/UD8hGqfd3xZwSFAdr2Mv1
Y8d2NH5vrsO7RV7hI1sjHWo+IUSbNESvI5X9dyPoDe8MJ3fiye4PoNfw6Dmb0KdT
PfNnlmN4Ypg0rVLG804j0lOYkIDsBVaryZYl3xHRHyY5MmY37XQmJ31hgwpiksjp
IYV5DVyUDelC006RxSXh91qhl4Sr24QP0rjYhJedqTAFHoi7efkJpiW0yZcoeeHN
LV6U+DWUcHW1n5dj/Nrf4Myy+Wcoght4lFxV9Gi0yStqeMbqXIqyvjq+Kylc/sQ+
ARb2u83LiJagAv1KQikYJEVxMnga3QwnmPa4XlUOh4lk2Cza0NGnPCxQGsYtMo+8
BsVKK49VaQBwVjuPMXJwj5ywqXnyhy34TXBLKS/j/DXtwO3EU0E2INADgsoww+lL
0URINsn7PgN4REa8degAwtXLgB+BLzVGOkX2lLSDX+Zn7LZWOXQMlgL1crjbhMAZ
Gw93n/BtxaHLXqax401GgwQfNYYZ+7zjLGmqteKeSMHHzF2H7yFnrAiJ62R5e0cX
LlChMuoFMAJfIgi7xtWQphRFD3XeNGKLXIM5hy3g3DSTFS7gsM8smBhIQL3Corhl
Hdz4DVRVVIW7v1nik/P5lLKBYdi4E/V6tgiEpw6mZ+fFst4z82f6mSCpSQjFHAeE
zBxCJO376kGABgbnVb8xLbB5YUUgva1B7O0Eke736xiVMKk4LUyxFTuHqw3tb1ih
fdgifJnyXHqGDkfWEx/qdxB0niEuVHhfcrHDaxYnFBxV1cAQh9qZJCxJopOg2URw
xUEaO8/Pk1q8HbSUwGIcEUGLUS+jVb+4S8w61gr1TdZ6RxeJiMFfVYqxNwFOHMSM
GI3Tgxv+XAtRullu4LGjtPTiADldm4I+G6R10QzqmglN5W5jr0LspulOHXphw/Kd
InagLnR0QSddcxaozNTUIZIGWpj9Wk0/JKxMToIm954fNSkRWTQYBfKhj76U4+Ii
rYY67wEGk/ijKG8/4Z3p9iUOF8bGGrzfP1B8r80d69BeGfAhGqfnwjDRqfC9tbdn
1nrO85R89csiOhrwaTSSwHI1naF5bI2kkLxKQWf15Vtp9yIzbzhujBoJRtH7m2Xh
QtE1IJQFreDJeaEm9pQWKY1AgO8iL1E/xANQ1ACW5kZYYHhBBwuxwrXOnJjjDoKi
YTOnSfrsaBrQnH0dt+3fwNSE7c6T8aCAyBUi8rcBZvfz+K6+Ips0fS9GEOelsLSv
0Vix+Bmx6/5svR0MZCWS4RbBwRYasFhpWlpJyBdiWumO6X+wH42bnX22lRoJHhDt
TrIpkWWwHkKKBN4KYJWbJUDzw2TaEa2zbDuKnLpYfveQTO0g+YCmbCxU07GueVax
yMLWvS+IvsZLXSbWvDO/4tcX5T3nk6O/Yi+Su2VWwuShOB+tx1C+Wwsnwb3dyrwD
PTAVs+QfPyl4x7KsxkaKn250n0IjmC7EjEVHgUUaBO+F9pNaCe2x7OhTrpoaGr6/
ME/n2e7L1Q8vsiLlTi98CHciz0GUmFDc5mzE/fX3hmiwwUyWp3WTF9DJSKSh3KAE
iN3Pt72MvGegNCNvabU2kPSJRvp1f0ZxRpaiPIIShuNucfXMN2T0H97y3YaBnwsw
G4FuliYZVBWsrDJyEIschOhW5rZ17W75GFkLOEssUbSPE/bbpCLhfNqKhIt1j0ku
KjEladEKfXyADOTIe7t7UESBWOcRFkMoadj5Dz0ZZAcc14MCoMLB3MVOtCc/rcIj
D8lQ2bhy0gfjv/kSWnTzuIlk22FdWEOn5WqkA4IzX0Um/6VAc+cR5bLXhXGS6JSv
lC1M/yGr/JcTrj0NHnKGjMWreMJ5gPwE26JtGQ1ADDzLBvfkFeoOf6FZglWVfZm9
I6PrJQz3SIjhOx51s0+lOyRjHL3B5cTFJGPW+itMug1OVo+cePtNAG9l4T14Ic8H
83KXO1TnlQvCDhzaGSeKdYQxeR9xgUCzYC/GSZ7DyUGdEwZx2JRel+VP6/hw1jp2
NEyQnebLmQGdGQ8fcepi7eUzVnUfeHDKFAYyMGeaIT3sQcThkwjQ0/9BrLzKPlX/
tqMc+x7YROKXAgAWuAUkjkmbjr7dRxe8CFgegA/NLFC+01FDHMQRcf3sWVyg9hZT
neybLhMNvseuoRabMEPFnCyzGRrqjN8nbrwY/qbGMk8uspezPPChAfktc09Lr2/T
SfUM8N5A09vPhqthhkQwMDrPL2ys/GMFPoGwycNEcYxKF3lhNpN2kZ1SJ4XZ2pw2
gbaTmTg8xdlRkwQ97oZpy8jtiJnzJ7EMml5KJpERKmOlyGdnROS5GeMR773H/Ow0
H0vIjIa3bIMen/VNqkCBQrIHtuuYRLLOaEFakvylEn28BNc6A0dTXT0VEFzkcyFR
Nnzpd+7W/Jl6/kK9Lo5VwVOR0rLN7mznCRQxiOFvywFMVSYM1L3+AQOcfzQ643Qu
SSKZLuBM7sQW6w4n74pwuf6yQnbwBtiqZR+ysmgFamr8W4b8u6nhrxRKeVmtS3S+
gfhqQgRPOs0DyjleY9nVaOjHPayurYM8NDlLtRSOsLnheEr9vsk9wl6gt03+PzDN
hndfr4/vQThyTa2hpjFpNGzuCO25VJmj0hDRkxenAWdfp6ettYR7t5nIf26Zn2Xb
CtxV1q1RGw5t0Gc64xc/ifuJwF82yXlag8aBGfsNXRA+7EwJnzxg0AxfvuFvKW1U
fKIAcTtcoW0H5CYC0YoD9mIQG219wKkUA9+fjsooXFgHCFDDkGtolDE0LT7MZRa+
DihmJHPJQGWiqK5PdPNC1+x+EJHhIZXQvmhz/mzI6UZrsT5LBjJwIWShI2jfTaMD
GhygwebmvVcecIIwz8pmJnSEczUp1bgrM5/d5f1+PzpKIs7+RdDe/kYT7OpFvYHw
K/o/D7VFv//1de4ulx96MTT4H+E1958dMeC8bnXeNSUODqC0LBAE+sxuIvGOzw1O
f6LJ8D9d1YfDiEeDalpt8ROw9K5h1nyyPbm3Uu7gay+GvfK92sBEXnhWGydkB5Rq
Ax8x/rru1x+llvvPDSRshfFMGIXfzMtiHIiTNggvtdeOScuzdjStgJgYiBPTxtLc
LAoh7cXjwF0tv7OdcjZRAMKAtArPfYta5hHFxrSpnN3BqDhApwMlmmfAtylCZLdK
jqNqJ4dRY3klxvrswzUNnpfHbwWTa/yLaIN6oXs/3aoxHdbprGAdhqkaPVhrwhSe
rw4SNEZSAglSPzc3uu0Zl4Y86iKoQ6pEZsou0iKS2HpHF3DXtsEmEIPxxrynukkf
QExtO9j+aGvZ8fOtd19ZF/HkfoBx58KyjJrWwjyaGSeyV3zioHuvzfmpU5zf79AJ
xvqHBAPy3SB3z1ksOAl9AgS2pEYqNPxuYrKSZXjPe8Lf1Bv6Lm7KwhsJt9NaW6iQ
wBTnGlqKQtpAXYEHH11aHxP8Cv4fz3xiVPfdYJUwQmHAHpay7W4McnCWJ0Zt2/Aa
C8PqUKMZryavR1aclhKzasBYr/qFBlZDNFq1odSNJ3+rgqfEjxiEarDhoP6ggnCW
TDcZQV4T42wrQUU26SRGA6x911J3nPAaz4QYtoeShuGb3J0iS3UUd2Teeroc0fXN
KSYUuEYb+hvmyTntwIqvsGYuy50r/SauBI2mYC3QsA4pTuk4EsTNgUmnIZEH9B+F
uI6Pt+EykDlUPFwGdR9Ra5ZFmQ8KY3tfguo3BULAiI6uUgq+ZCB6gfDehn/QliB1
d9ML6tjmhFNwkL2xDRxha3CX62OVRyyylLI16aeX/rezqczFTeVzT+xr+sswFa3N
c0KJGrGxqRO+z0ZcIkoz918sV8HrPEzttUsH7evj5b89pGwp7fP8KZcz/cCz2p+G
5vLBQj5wDX41crCjaTy0bRjmO6qKlJpOSJnaIZ11NcUBb6VSCDQFYVCAIhNEU3bz
EERKr7aFeZrOE0nN7OlR3pBW9DKfipEwEQQpkeo26pdNYFZ4anrd3o16nLzBBgDN
s27W/TYeHDWnl5vkFq87rNnYbQHciIrUG/drL/O4aso6N5Dk6Mw05LJa9oOTVgft
bLvpTIdnxnmHOKtECtCKKqOzRyPYKjD0zSJKVRFjmbcmZnR5mAdw7DZu+YGoVRUn
upcqxuSeLfSSJWahdWiA/FTG3mXRyuf0bXTQS/VAcKw33UzumU+AI+wRq2hYgeg5
vb9W1FeUTVti0oqBwSlR6T1t6PeIjR3Fjjk3MxCd3s+/1LDQrr56udycK49WXvgv
xZAZJ6U0sBmXfUpcAshV2a39/YLqstdUIDHVDyP2R4pwH9AThWHOi8sODV2dGmFb
p3JIctck+Qtf8dA3ocJjYVbkrQsHjC3aKoFvQmpUrmhkU9h04ksWMW+ab5X3ysjX
9lmHMdFQX+Z0g8fusrbXU7VeqUxNn+crnilO/Tgb/GFj+LaOzupBHiBzy0u7JmoP
vLz4hd9+pZVjuK8OrpBAkqccuwR4Z+IeeIR0mqOtnXn+wG1MBMhuGgSp/mrNGhvm
FVm5RpM5Ojv2qCaBKN/hpFhhiCt7VmWnf+J1J/La04dtbeXY9nRjlaHL7967eD+4
gItrHxJAA4P52GoccLmGw4SypzXWDa6wTQZNkTrjHxRFkMM4D0+gKiBIx/JafugY
eO5Cs+zT5K8SewoYIINrP+R1TXrZEVVcgTEf7nNDBchWKxst1PFUxZGOBpXqxl2R
n5v190qlnXImz00ONAaNewPYi7QzIZYu0kMBFDUDwCYXWkrJHDBIkF3YlgfEMXJm
60HgGaD+JIKkRKePXNXmcAWbVf7F3Rx36/5tRWpF+JO1+WVT+lpY8vAIfpWXDLM4
E7yDtQzdvFhPSBy2GsJ2R1KUsAomoxj42jkuqPGx/4TaF943vNkJVcPJSwjqYpAH
5LQwy+EIrGIh0wApLF/lER7X7z3rvEs36ztTt4+RPwS1cMWA/xGflTvZq+RiyR9w
LIIqfAPTGF0U7iRo6gYnDv3IJlnlVReJJ9ANmqjIOLNSPoDB27hKg2rnDguEpPSJ
NGRRSfGx9JOMxzbsBwnmE7E+YQ0jj+vD4jHhlKCr6AcPtGVarPvPZYqLOhcb7kRi
wqMlHUhM/wP2Guy4eB8c1rRZtvabs9ppXu4W9KMBXsbY/RFQOGYMEGv6cstelqKe
UB7693Z5dRiU0dvzwNmzou0SRFwGPZw7Dl8Ynsb40SSmV635Q/k4d/xzLj/bfO5C
w3IPSeL7IgK7JnwaflWGWAZIKgVZ/41MhbzAk6aBUjFr8zfNqitfJ0D1MBsUACzO
XJBsM6gs+BUAhtpLWRsogBfhFe1xcvkR16HDZV/lWWJmAR/pd7tW5jCqjAJv5XAy
uLaOzftE8GZTu3/dlFE56ljCRhgB52lO/qwH7NT1HqKWvWw57ikJLiJDs4/xNeQc
6wAlNRKkOedkH/B6Ifc00FGfMDxvmHdSlAi5McmLXOboCQBk77Vz651HYztcuXv0
WWOMmOHvYrkmpv3M4CVjLlCAn648aCkETHinjZG59mlkk0Hjxjt8yRiQam65C4ui
MBhN4BS+XbPm0103lKFOHxwfXSJW5yAhZX0JLFVNGhTSlgyLU/PBFx8r4B5RmjuY
9pdcxCzTFlfJrTaQTjmg7pOsLYAYFvJHVFJCwJWIza2Ige+LGhi5Wo3kQCCB6ChA
pOZU2RjbpotLebvuTECmcOhRqDHclI+PxVRZx/dv4AM1tyGZFiJ+ETQ9y/D1rTTf
atP4ZURA3NAso5f3lASD8LdZbMmm6N2h/ZxVkmsgFdRHgGlEADwqV7NDzRZaDmGp
rFeY0JubaNF3/k8NBz0+jD23pjAfXc2wvx+xTDjSLaf1Vr0dyixgKrTtKk6uTAav
DJpzESPDM2HubRpZpHGT9KoLA5mjJqRCl9wg8VS1vWOeZisJDjl0M0c9uBEJv7s2
qz6PM6iZekSp2IkPCeC80RGTS6jt4LuKVCmsxa8Y0XvThRevfV+3BNgBG5zocC0R
Ti/LZ2mngnxbdni2K8eA91mbxbGKEFPzuU1+GnmLtRPV2reoIghT88lZk1ATjWMk
zwBhJAEiurLmp+w1TiGFVmyUFR5M1n/HWCPJppieN5FCfYgFZYaMWVLVQPCKIa/+
syfDJ7WD9SclXnG1Aalqzipgq6i8s8Wz00q+I3KqvBrjDCt7AlHEYJwfRJlU4yYd
DHBM4fES4a1Ul0bbKgaayIjf9ZmIZL0UFihIb1VVBs8zzwjNbsJM/GeasbCdmAwE
TrtCkm0zStmrnXxxG6pPv/HKljzWWGLfz3Onf+IrB8aOXDGaFc5dZDXEtPgvl5Bf
lXOt4BkJ9PUItOHyqzhND0QZfCCJw29cMIJVqjJHFT8dUytKm6rMlq7y+KhV4Dvm
4c2GPu7hl6FWTN1DyKZ7/ubAlvmkbZrK0sm/wuR2llthBSCviVHHOsAW7kAZfJve
BX5tLSpGfDcrAdWXlk2uHJw4wsjKc7kLJqSCVzKJ7sNMnr+gthDRaDwPt4jQTyTf
AUpe4RBCtWaTBO/cZYz/s1dLXYGOLldbtmFBcP1Fx135cR3NtYrcGiaqzRg4gsg2
ynelBgjsUs9xrUOdj7Jowy5jwip+8VxZYfR7/Cl6BzTWNV5vUbxnuVFz3/Sqr+Ir
O6iWcor0u4s0sqAKXCGtbRKaqfKqc43MoscxLwDZLsrCZWA6/TjH3LF99GMOkrjG
bnhtmI/vE5yWjHrhqdqDB0k3RXKMrBGq3+DyyJXTx2rVK+z5LA2GD6APG5GlPQu9
77oTzKn1iP5/WsZQBefIgdIvhZOg2lzKelAVlWGzVoeNJ0sW/tkGPeof4VZVqCFv
9ilDRp2hM6KZzrEdun6Gk/LtUm0qYMLxolaFDIIjvJ1umxXCAFGzJd6lJNohjPFz
Cclzh/0FtmT/AStMldVUYW9rfzjwl9RuGzXRGNkUweGcaFQ5B4JVKKAFcQLtdVMJ
JOjPw7OhCDe5xEYeoz03gylfAtaOFwrZrEyMGfHmfkWilXYW+2bFbl+fgNqbukvB
p/7quvWkDWoGSUU57vf1n4tWHC61bm0R59HmwgxYkBw2OdfqPfTGzJG073ovKKSt
AJ3KXDjoPu0KABkbnKKXYQeN4m+ex0ICYfMu7F1VMsecAyqG+vgJFHVwmTJCuhv6
ujWzc2kyFei8LSTzO90lFTKsldbME0L4LmeoaISdJmIicnmsb0QsFiQh7BicQ51x
iziW4cwHemO95Hf7sZs8a4Qfyz3e3vGuRFnSZ7ZFanNzdWFVXzzdzYmYtZ6j/Kk3
DWGhG+v+FzbrOY3ZSQ+UzgGqUb2gsuP8nybLhA0PIbA/pkwDZdI+MRIFf+H/kzm1
/kqEvmlBPF4os7qcLcl0C2xtvBRImSs1n2ZnMSyipsltWdDFBODKRkZ00LU11kyC
sr6mtwooY9Af/Re94fqGejlDS94GAwDG45mEiQ8SUW/STASr4gTCj06YhMpoNJDT
b5+mm0CqD0/VQu/Zo0VKGCLdfwnY1YV1b2eJO00V0Jtab5ZtK0spDXs5BmsYRFcP
kTCAYWgKeUDeF1pf1tPEfEQduuL4MP5QaDH31mUYF/dTL5ugofCoZMmPv5wnTQ77
8KAQlSypqqAvkCNy4o4bmLmnPuGzIyM+w4N+lPUj20dIj8dFUsUtiF4DmfI+sY82
jT0u9DuqbDSRTyZdWA3lcpACBoOHtU8O6l8iZNnkyUEFyMmOxgvFvVJjqbA/m6uk
r/ZTL2aExuHcB7ayj3wEKQl4wIEgZO2oxDjtOO0V2S/bjuZnTuXKgF7G+mywDdhh
+142TofRR8LiCsgVZR5hv5fyjBtGKHQaLIuMYksJTvozbD34GfBo1z6wGsyJgFGh
qtn3m1ybibNARGr5Aqde0DtX72dAiNcIzKFG7+6SAWZ9szoUR8++KHdTeuOdHHbK
GWI2fzARFGBfOWAv5+FHN/MefqTFn519hnKU536mAvsruAr38ltvx0pld/6PZO8S
IDzbv4kh9BesFL0n4cXISaQ7d/5De8wnwUpnf5cNj8bRZeFsoXIB9Zog4HNV3JEg
Tcd5ygvRWqoNdpDxe1zCdU24V3F6Bwj5RRL2vM+5xr74ql4aHne+fIjRPWuk8O/v
GnfARi8LJsVLI615Vb0tEu/j3HsXK5y+NYgy02G85D16bM6n4fURWUQ5/ue1+n90
uu+tc0fgSsZbYFDLaW0NxCn2DDNnhl97i5HT5TessU4k8x7PxPTyusV/BlDYIHiJ
4Cnh4EA/rBUAvcfW+Vd3hBobCUIGy4zGXo4L6kpqxCYuvbtDImz6rHhr6tQf02w8
Vc9iWRSGb/bRiWGWRgelAIe+sKNjeKb28NuXcFb+ShFOrH8Iud/BbcZRekGZCqv5
hRjqNwRXVqE/eyuLcGQcgddgeDQNQDulmm7pFb0OCr+rqaFlcG8+MKAipRvjBPU7
B/fy3HYQ14g7D+Kj7xBqCINLehP/7dAANRdehgoaEK0uWUVqvsQ0HeyEYF6VAGq5
Jhi7z0qfJ1RuLl/x6hPcdCE7+MYrAdnL/Auyu372dT0ltbKabuoT7g3gY0DTBJvm
QvGhPbqcew5dM6eKb3yUlOzQRfrMpzoMR0uBXRtditYe7+c9ZtV/Fe02OwBqaWsS
0N8VYUKKIlrNodDXg2+pTVgYmMrrtSVhfeHq4ssRd001ItNbU/8IO0PWiNMuYRWr
kphbefw5pMVSz0MxBw98ATnEw7AO2j+MGoYiAtfAMGuv9AclmzO8JIhzsXcnvWHi
tfrjYAbdZfXyBloPw+B3a10XpKNsGWm2TaVS77ljmvRVSGeRMRrbF8JIF1V61ZsT
tfIWedSAMPXD7iPIcLuJc/z0X6PwkrJzlKh+Mi6jP1qXxPI4KsOFH43o1+ycDoPa
TJ8sSefewSB1THbrETd6/r7Q1StrKPXNL1b5bVzLmDnf69PdXNcCX6DZqxWrkGhN
M/ooKDHkR6i/zJ5gJ/FqV/iHSpiIRVqBm7gMMbihBYEN8d0o/97Rj9BgVkZxD7R2
CE6uQCxm5+ZMqgoDi+7L826lhjkd/Le0ZNXhSZ5CSbAMCgOYrKquqz7FGpgSx1AR
hDSMIrWICC2xkcITc4z062jc3HBc4Bjs5KvcvoBTUngICLmLIpnXIhaxcYL9kl8N
bqBxgnahVOkMF7tNvnEz+0WboR/ugFKDQYqyUhHa9uPItgVse5BKo5glbsPKdyq4
J3qZFw0m2HpOJWVePpr0cX5sgk2cPVCoUqPbQ6BJLqTHA1MhU2gzu1EBVAEvshM4
HiYechj5NICACKQqvKD9zuUE3NXduHDsnVT/S5vWq8UNSZwFPF76qFTKP6Wyr8r0
hR2h27qblwF0KiUwWu9CkP4VGfjh0anQgDTLZkvrA5RQu3wA/dFEonGEKEDsKWk+
1veDsKdn9HXxE93Owdc3GSLZYwu2qEUVJ0p8n3ZkVQ7M9i5NVQaP91UkBlNzOOBC
pdj13qoaRz4w9yygNoBwjaXuK52jRXwtU4swhzhUcD+SJ6PxXOtoE6uOTYHw7L1q
nUfZKJ2GoZ4zdTMbVedYwUthbr5YPsR45D/cyocAH3qJMPnbcei+/muu1skqn3WP
rPI7ZNzeAPH2fQItNm1+PVkNhjdFmtUMZKa+24fx30D2q8wdz0U1cSFj2DAvJZPH
jOkL/Fw88rcxC23N6iUERogt00WXGoKfN+JI4gTWUnJ4dCn2dRTWQVW9IstcVsRy
G9djeSa1xjRXGxaHHykrwoad4z/Bnf8qANS9PfVH5bDwcrXWkOEhkT9mnuz+k24g
OALDqvPwbxla/BlQeLS7KWRoLdhKDZh4g367JXGpSdkeMV5j8xX+w0/siFJdoi+C
kKsiQom1urlEpfI22E9e0yrNp9O8FsfWPIQl0povtHYnQfk53CRvm8yc36ar3tve
T877G+cS6fa+jxSd8+bkFvWFKZRtEO6dVJJLn7eimXjuPlRj25tyxF3qcdoY4t/D
A7n3pvoDMjBmgbw/MevLJ41fVZ608W5YJFUY0oIZsckLliv86wkpbngT5zgb1+VV
pIKJTO89O0hBZjQDmRFQOuXaLWz/xkX7lMFmmi1eQC5BUPA9Bz/5pkNekX28HLnF
xKIECUpuiKPox4CjdoulRcYSb3jVKc51TVM5CAi7O0FicigAIJT7bO6TdoiBI8Bn
BToPAEje6qpIHrGf6y43C/5wnbqBz48xexhnRVZQZuu/fKpse6Ur+lk9t0sILbsV
exNHCg/On0N/ba0aB0LrIeLGtdCkofry+odN/bsCQ1Ld39WmhPiBPKUkcYO9AjZ1
p7lE4wwjRyDvc06ZbTEhqjKTYbyvtJiTJqcjcbr3mgrCxSpnkvsRKmUTQPObdtEY
6pL5b5iwRKySmDoXdoYv7dtTjhnZa0033DH6XIscLmIJorSY8co0CAKp2b4CTNLh
O3qvwEj5wxDJ+lMPetpjVkHDVnCHfISXausFk7VKBzqaHP81s1ZkxAyf4H3JlmXy
ZUrKbAnVFo9yyJXItCHMmE4nfY4X48stX2IVQ20Qd4wK5L2SY6V12CP93g+cYrkn
hzaVwLAcKEbRZ9rAuEW3AzDLz2RCr35TSqUWp2OvbiCcLXT/I4lHVpXY/7ryHT6p
OSCGUWrVWdSfjl/xX3r1aTbpfNr/CfiLya/4G2de2zJLiWPTLWKx5sxJNuslQg7u
MHwoM7ZA6M/4DDDEKAnXEq2KkZbx1T32++qmf4BgPfjfmGn9mgmqOx3o1YinM7Ri
mqaW9TK48hzq9EUdEh5oK0VHPT7WaJJ2FUZD9dCv35mKdb6LllIlWEb2QH1zyrQV
rMq1oOxNYA4XAJ42qyA8RMj04Q+L5t0iVv4lqhbAbP1nAPnkd8DjFe9gxcFK+ZlY
4idFE1lmSuXidE88jmS6zfmYcrMKM6EVy3LBCz/FOwK14tsCQAQKcbjVcrzO+QRa
tdNE4gYOH8OoqX0MQnfO4UjBBA3D2QdhzrqjR5g0TIJgyMno4s5NbX2sDosvxCjI
2jvmJDKslaiR9BnROBa+7jmKqZn53J8h+muBygnAicYupq5/h5s/scBUFZYOS2JP
Xb2EqAIssZJsb6wSi+0CngJLmsC1oM9iRwlDesqxBvHZaYX5hpho1c47O4zn8rkD
cygRexLvvk51WgMUzUULnxcR1sotufB7g2W0kOmfilzDgH/GODSg/l7zuVnxJ6Fb
TqHmBck0dlRhulR2csbqAsLfRPeVKIp5Kf9DsSSwul/2It9G9E7Eu+q8tH9YHJ6K
LFHYWkLJnYLvab9gNVmqea/ohRI0VhXw9ldHYRPGmCaJDmFlBTXhhZKVO0EOuhM3
j89bF+OID2jQXuHIBjAwbwN6Tz8DwBIZ+V67N5JwZPHlcxY6cAMwbUh+hIgIwjsG
hUgPdOl0xJQPO+AJ50z8S5ySoLLvgxKEPsI+qCYUk1S+57ExsYK9Usg+YwE78ef8
snaNNK6ovaPAqdAdF44iCoPQ/zBUvDTHpBFzUh3CveTgkJWkLNphSaX6svkEW/Rl
EW/GpzrKwY/Gqxz3WL+NDCiLy/44DiIJPn1Q9EJSF5qH335qxFlb6AKxEoC0Wht+
RqZoqBYXHDIdXTKg3HHFRfMXQ4dgftMvDLjpzfcy8+NJYZBU9ILBHYXzZrxJbAZJ
4z+1VNQ350pfrkuw3wDb2L2cUlEkCTyB92CSfqSgKpLIjEFweu0mgaRenOVRK+6y
+owRlAUN+prasm2JmBHNhr56zCxeVsLkBFAEF0hSJFYwj05J8ZnrbhYhDiSETT2j
G/hdKTG0HuucpQcA9qohzlnR2IfNiLv7pLByk+gbDoVZun4zJPho7cGLsqmPeqhh
3zczq4HU0D3P9YLIJxqhYjds4wN+Jgr+LMkLILp9aESj3SSnnMxKkG4VJ9D9gOR3
hvAq9fNz0+YJfkciOjsnnfgN340iyO9WxIUaK8EROguWgMY/vwsh3g9PvjarruXX
hbDVxZhsSqYoXmvXKPmFFNJI73rRiuXLPmKBPP12Leh6YzGrELBWHRE/NEXB0uLG
DRoC02cvifdCiBE2eUKygemHqlEBTGBRREPFQbpqEDP71Eh4KoJawmSf9RKM+JVL
5jTod0s74kWZ2sEZm5w0jKfBk1/NyykHI0B3yAnmt1aGcz0FVB4QvNoOvmFXVaRQ
cgBxLF+wlJluKAwR8DlIOC57LE4hzdcG+eT8H9Q9lg9YmUyOcE6K3kPKyzJ6tOEy
dSh38TluEn9e4A1iFTV6CZwDt6GeYheWwWNm18vDLVTWav7ePOy3oQz+WPcpe7AS
s3gwfwFv9YQM2oIJRE+Ix4lWEo3KLCX/QZ916ByjDGBcvYQlRDqqgGP1Efko6d43
i+o3d1jGQDKss5rMkPoTiR29K4DSHpGW0ew8cbsTn+nPsnzkVN5wPBA+6J9sz4bD
g0sQWPmQpqyUBSrWAYNYq6PqSrJ4BWdDn5UPMA04FRZtD9eRm9Jc1QKcZESSpw8m
EFitJqb1Njih0uGP1srhdzNIgdY2KQRdTQpw+V2oQ30B++KK/28cRHc7wzIKiP1X
EPCmoP1dpwMCUT9o6SWxTqqSjjYitEaiJabK6THDCk3d3E+a25L3MBqh8WsL9ll+
RHDryJVloscTHNtiQz+b8UXY9IZkJufl7h5kkoUssG3lc3c6EGDeEugNWq+hX7Nu
L+07E9BdBa4nbMM493P7QTEzaCvmY8XJ2RE7ixOZ6CJTKwsbjH6JNux/4F1M1YaP
g8tNqx1h095KuDYvk0eF9cf1UMlEUL8RPnjfcgI5KcLNVkh7/pYQbw8oVuR89d9w
BojmvNKremd9DWKHG2mMpGqLGibXA0TXOYkE9Vca4CZhEMTYeHv1lnCYmctnYxTS
JGGt05E2zIF4eVEP7ni6IUPNDDYswuEaaGbueIYIGZl7hc3mx85UA8rUYgQhoXw8
DhgYrJ/cbb2KMvCXnMw3pObQ+yWIwB/HUhlyNrU/wm+O7Ww9LzhOgShmKTEjW+eF
J05edfq9+3wJ8cMQspjn8rVGmtM9d4IIElEuewFJGFw4vbe05yEs4HRMSbHwViPl
Frs/e4Out3T9s51dTDOHsTApsHMx4q2rrcAEeNoBI4xQTJSFOBOKc309XdK6izia
HDahBHh7egrugbzCHBu1aZ6IcnKgJ5yzA1ESaKcDJhI5+XdJqZgsXqx6D+IHIFdD
Fn4PWe6oyuO7efeOHq0IOWgw3qfYUkiMnXaWH9MgORfPrllze4P0YDaB7vN5vYvW
RBPMFdOcS9tbxMM6+iznnQyD0aZOs/pOHngMD92mYqQZ4kfvt85CIfcBw5yjZTGB
kEKIMeCC7sCmT50JqEEVx9m6YSvah9CNBungAmTcxRL0GVvpA2JlOhpMTAVGOvQn
pQimem73Baya88A6vsjXhewvRARVi9CFvFxjqGnoGHn4U/h9kRUVSEYt7JZJgvvv
YAnwbPEj4/MUk/i2wcvd1Q5GkZSYwsLz2wQ/lsBvhT7VOPosob4VeAkFWVcIWy1w
v2UadLOg0xgO5CPyOIJAZMqtXt+sYxTJikA0XRdLi+8veOmRRnr5DofZiXVUHfuH
oKPKY5pE/4n4nEIkRy2K4QY0AIpGsASyItsX+XG5N/JVoMLWpjR/Saba97zVMG5u
BAQ3fMaWw3uu0gfsUQBssAMEr5xwRlJXbJOvzdd6hIl/qMDpuXITnV8gtRvOBq//
p7SMaiqPro2eHG3YlpUVdfkTU+itlLMYN5yy5U3PaSp3n6sJKcGbY8Yl486ggh/g
UB+N/qK2FZym7wT0zflQ4vjXyZ/P/zzY2DORV+RoZM8yrnU2TX6+MpaANsgh1S6K
WadACk5mwKpC8u7vP5CmiVT28XY0w+iX0GRbRyKci7t3ItI22H5+elFrBJrlkGTT
S5TSDF0t40JAnth1Qbn+qa48bVyh1SUao4xJtgxVDAu4SpxAUujqaU4i1WiBxxzh
qN0NgYxbwEniz1GZKB4KKiCoNRT2UTW2uT999LcSfWpWojwN2hmCNGBd3900WbSk
ZK2Clrmu51aJZwS27Yzch9o7jlBk2VpSdl3eU98Y4pazFADFGNG7KatZk6Qz+UEd
PKuoVkLeJHkmd+v5E03mvB78tsqVSmKeRNijzEydKJWA/JKGL4Rqov/zPzHtDa5a
+CY7SNYKmsajcGlhDjOUyuYQi3zCDKaguQ1uUxm1t+mYmyBj6AP9H1za5Q5afVyI
AMcsoqZvcvEfzjOozEMbXGICWmpGT+8u5DOLRE3k1PYsIQuMuACXxPjk2US+iwgP
W1Xwq8V5ETx3yDa5yKAw7xkEMFk8HZGNc7PgsPoX1GbFcAqcUZezeUQucyk48iRK
BZ4Tgn7YvFCO9LN1cB2Q1T4un87A7k0kWcA5WIBhH8DLGG/B3JYCjQZYPUwQSf0A
TO6emw1zeyp5Wg/4VirLnDPuzUqGh5rU0SlaS0TUbodizxEiwSrbCGZV8fu5S9MI
YzzOWjlwlPsChPuDjg9LlZiXiDJBnnuedS4EKuXoLNo/hkIdGJ5P37IO+VpahpcC
yYFnKX/oenwc6GuXoZjAWrQUj2xxTokh2q7hGmHwIaWLJXwUNTI6PC/At6svnOT9
bnUUd5L/yoF5XrZwmYePhah4dqyYG3qAoF4CrZomKwT/CMfsEMFj43FWHDvmPira
ZHk2HM2FOWNhBwhT3zc+2WaZRcu/b0IAJ9cy2GlH1apg8XZh7tedP6ldhCMp+iZU
lha1mNVMqfWCVqTrQQhWAALF4kRDNsrGilyj1hmNRxa2rNXXTkWeRGcTOGae2uGj
qxH53+PxI9Fhpg6i4hGGNLMEqoYm8hefcZXhmHrq7pHb2ElIipUDFKzHkG2FjtaU
vNki7T6GHdER52CsemYKkjz9oCGqvhGK+5slCDXj03vuTYTDe2jg0Dpflc3aTKtI
ZGNwAXCIfgkT2RpQc9LDn1o2CBjjEOxw7vyyB0o43VlBKM2/DiL1TxX/C7pCLnKd
oeaHkw3UHKrtjP0/jD7de6KLICwkBDlCDBmwutxbpWGQnYcjv9QZ8r1oH74gGOo9
n39tt/J5An8eBCKbYdCSwxZ+kWNmjny3X1YC9TJUCpS+hmNoha0az4xPcbMn9IFU
PNeVe6LJrHW1aYHzOV24VX2zNIQWDGAy8bsHC2siIVDrnkqN2coDsIO44kW1eWFq
XufjKk4MJphRTZXXKOU4EuMfOrYxrkoQeVO7YA14XyE37Bjv5ea+8Rpxsy1J0/X0
UTWYJYBVQw8e2OWUngIY+etMUqtZs2zWZTSbNPhesyvy7wageLD7/IL6PtHLqkg1
9TfioVq2tHvHLz4Z1tRf5zOUPh3zQEBx73B84vaC73160cgbfKTGkeaWUD92i+Ec
5dHvzz5GquM2mRLf9k285ttgU10cY4Kjjufsu6As6vajFSS7zd8fzrefqdxMUeCR
2+oQmXOf3uHZB7yaKykWKxaCFx5Ur4bNhPzmXx6INAu9h90ZURpXY0HrwAVep1EG
olfdp/2JveCZlB7QawFGe3/Y9EVIxX/1ZfXlfF/iWgvCiBbTPRib4J3p8PSy/Yuh
KSFmuwKQ0S4gL2ffPNfjapmnRNmvkmXbs8U7SMDDGjbWa4O3fLkTVHePerNeL8xO
GluZBh8WHsuNVw9gAdKATH5+aiiC74rsQtZLItsETr3sdZoFVc6/HEHXB+6sLHoX
lhcj1k9i9yYa52sPHMJScSYnHMZ52MoMsXk1jMpRGY33XRmz98/lNMLHuRo6BYUf
4LtzxhTftMUZLQv4XRfzM6p9FFfE8BhQI2e6j4UYo7/RixPKfpjH7OJ2ERb9vTWi
h3d4RWoZiCn7suhZphCwDxIgggCI8yZRLSFCKemc3f7kWl/uHo3QDp+lE0BfqOQ/
aXCEQ8kl2ixeFvxxXnU0tI3h+k28HpPsijSQe+hy/lnXU0LrC80n1VpwSlQhrtdQ
1nC6Q7b0lxqAz7d0fnVXODafwdMzrWJTrDDEo+E3nWuEj10fuUpdDy5PbKzRvrJG
SOT9Ysz2SHEw5+3LL2U/xKjkarg0CVF1PeHNxBwzxnd2DOjUjhJph6SP5vY9/Quz
bAbnYq0JhoSndP5K1EUF7WKz6J55+p9DvU61qvf77r4mwZsEsQb1f2jFfVGUYkmv
arPGbYZjAchUFYkuRazEnoS5BAeddz7cIr4CiWDKpt5oI/3j6P2h3ak+mK1z1AH3
hYiofe+6nWoafFXlwvhYEPvG2QduztChOHvBkMnHBp9jzXAz1vhJa3kYwGW48cE7
J/LJFqMu4xO2IUdABiuorSwT2YB3rjr4DnlFnlSNvHenSV8COTdJ8eBlhqct7N6c
xffxbhha3DWT7YndvIib1fIOQvSeaTIOAB6krJ8I0xZZBFJGQV0opU0NR3VqdSGu
MocyBorHRRZc1KcZuzXNTWOJw9ta1QJDJBqBMp00OK3FWThCYmVTw8V7136R2W/U
oo4g8Vhd9w687KmKKhuo0jA5JFUGDkmGd0+KkELN5pKQws2zZOOlckUsIMn216ce
iZBgK6PpnuzaSewbkt95DfmPC4OU4+QHVHqH2wDHx2MXkNJIlqLS/RqKe49XyUdQ
hxbs6jPUDaSV7rNNbHy4eAhRn/vRhhc0BXxIXQmgZIjEitfi/c38xVQDpqxKEI4E
AjI5ILdsDNP7gyG4PrM3zjoNZ/3cINOQL7lcxzycX23tAbfYQ/PX5EBmtEwRZO5G
J74iyqeCo0t9Eqld2eN4NKlWv3eivM2wG39xib4AQium6iXjjkEskPIKvNdOKAjz
3AwyvX7Txo45IpD7nKF0Bw6l8/NZ5xKCrTy2tYsmbl+MQ3tV7AdfoWmmgjXesaLX
YE1zFsIM9Bfay1qKWi7keA7FY+rJZxQBRKoZI4eNeuPLmZ4pEPOjeT5oN9wYp5Pl
Lal+F12JRuTmfRETtG207yvXwNRcYJ/yaUexJuaTZc0EnRsSm8iN6Mvk8k3O2i8F
5ckAolk+YZGE0Zl/PHS1EnNNn28ZnJR1R52gLpg6qmvyb6NtUg+8Yii5uKc2LRTL
GWlycDMbI7uqdOwuUZOAt5wvbDuQ90obXi36J0WMd+UA6TBdhbUEVkne/j7StpXv
/PVvs34YEJIkJ/PLtE/30wvbjTbYNuwhW2uZ8k5pJcTAxxQxWZQ0lMZpw2xc2s0z
wOl5tUZgugJhBRYqUjesjWJQ/IuN4mDabdILpyMVekZ3RkBmVNx9HhmHhQCXm9nh
iDyGsyGWRj/a0aOobRofFfdcd7ewzBTrmPgghhiWmvURPsgMAZwN87uqpyjcWPHo
IZZTDDiiMFu4hc+8+BT2Roc0oUsibslyE7HssFP1I1NYzoywrPziJGxT+HMaRbly
51UgOo31wsYNN7U2YnuL15naK0ek7e/hkEem/k9DVZ9uJaGtI08QgFj5sUxz/uIJ
piYlZalvXMi/o/+gpIh3Ze8vuN5eP0Un1T3Je3CVCqN+LcAawt0wjJFD7dbqBnDd
E1xFIh3wZcQr8nG69aE4z2bAJjHhGfMyZsR0BmiFSwVVgMchoIMHRzkOPLW9BGLu
fl6IyyXiWZyxF5xV0KIMmSv/FDaMbGPeh23OIJfJhEdAFivGRFdnNdBP7CxVxNFb
xalTu+lomVicm7OlCCtC7/26NfhnVugK1zGWvO0HWwzuN8nrpIdIQeg47IRQPoxI
HOSr2wVBvtp5HcGz8AidYvxrwQHXznPu9YyM0czeSWrZwVGIc48BS+rigf6NMNFI
rCtCNDO7OI/qE6zFFdXy5HHp1u+DL0tnghDoil8s8HeTKWxqgTxo32arHD62PtHD
Bi/t1qaX7xEmq8UDTWSyJ5qD0XuNwMIo3iesum82C/h27LBFqVGRnQ73FjNxymWq
uDdwioad1ApogyytU9UCLTHoJASQ8lbM5zI2Vm8JrAz347gfIEcdXMVdu3LZtxSy
ikTrNGCOzfZqwp4t6DfT8Sh4Ia7yMNGpjtljTFYLdz+fNzGfVEz5NeWYRVU6TBdQ
8I3yI5f4i0Rf4ZjbjjU/L9b7ENF3O6DLYJTZLlaugBFhrsH31Cl76PXIxDCgMXNl
SmQOVlwGnDKZ7Y6EcuJ4S7l/iSXptvBmcbfSEtwMwxaf5YvKIxTTWG4EEA0sHvYb
Z61S2fKccgGAi4rZ5Fecar5LQs/3EDPEdTKQqkqn4X08PbsUVkjX+NtyWwmK9NaQ
D35bz3BKATyFVROBlj5VoYIirJDGGI7iBgj1VFeXfBrxg8uzcPrFDyQ7WO7dZHdB
YDVmLJkuxaghWTr6gwiuj+EiYuByaXRsxM4v+V2Z+x7g0nUECvpjbxo2/nawB9SV
EyM29SAEmZ3VU6DZAvHni2f4D7gHmSx5La7obONObQBNZs442rBBnBIKQ0rZpBcx
gKxFaBitH/nShyL9fg0P31zYWEJpGgD3ewTJIQAueanFlpJpe2x+0nYfDNX6wCM2
IViQrEjid0GjawVO6wPMNJIoBu+5qbjxTC/w+9R89/3DQTbXna6VFp/HvUs2C+6R
O4NaMCRlarnqqt6b7WfZ1+x5PEAtXuXjlB+axgWRGmHKVgzTskfZ5+RILKoZaVRV
rTZY1wkAB7mdSW5HFozqVLdsX90SsVSQa2HOBeFxWXUQ9eLwi8pxfiuJKhrLIa9O
T5qMrmlGF9IC9h5g8AZyMYb77pPEtPeZZa1Z8ZXEG1EprgTJX9w7GUZYVxlcf9Xk
TCmHS7X7tWmbi4J8SvBOkcv/XzUHm/tklqXhH579LtlkiRDdtvLNT6/V1YJUr85V
doKqhU0Clf0XDcWn43hHxHutUAIUxHp/pXbm5BV7U3jtRG+QcqxChUDm8TNKiyP5
tfQV1ZAFTjW0jkBaAWPpyKZITAD3NKO2RL8HTXqpSijJRZ8hB/zMdYA5umj1PxyO
FIZ/fNlanNVxPcMKKfH2YsJTqEkDK3NyQZq940DISYh2+0RU1eFreaRFl8owaYMg
OWvFo1JrEp6oDfwGSywkiTi/dBEvxx4HPQ0yTisgC20P/p/G3qKwUgN7bP9sxVZn
qySGMa5y1++s6Q5fFONji+k0A7Dwp/UGriKSFJ8o/CCRxxjYVzaX1tk/bv3hKl1b
T1rQ4QtJU1lPiEIPmUWMY/N6G79Tmxu7eO8NH1aSrnH5VuU1Prwmdeq4W9HYryzI
blI+Q+MMEIypHgRcFbokNnsMQrBVVB30l9L/RpEyqkF2n2JU421WXUcuU+bh3xdi
tSmkCrqNIxT4aGQt8M+2hmc/voosaKi4sQaHEmHzm1GA5/nS07nDQTY8BWq2oLgr
AguD3CsBo8fivoV2v0RSo/aHAIQdWJnQqIeic5OYGPnrUiDWydlHwloahJ1DRSRl
xa0EaSerNzkZHhGL6IKbOZeUxHoBeJ++bCih8ll6oYSfu27Lctz35DQE3RIkntkV
skSgALhhDiwbxZkT1YPCY9SLTZrnO0t0FUgxFI++mmbV/KSjzacGi5iZC8bttqkE
tcDGEHz7aYkrVBc17kIdx/RV//7qiK5L551oL1pr5fbhKawH7yMyjBi6C8Sh1duE
gpCX8AZxWgJ1aBtNkCcBocxXqtBHkZMflRmNBsj6t1+NCAmnN9lgSMtAmnMJBzG8
Q2gAAnPwM5EeWPvoUW1N/t6Xw5+lekw5BEvKpiH40JLCitNmExR/GuC3HH7Iba57
ZEy4wQXQ1QaX0V5GH/95uMVr0N5HzTI2hNQpg7DjuZYC9SVjxWT1JwVjBcYaFJKt
PF3TINBpXI95yxbTMzDWZuWgSTXXUWuTlPjpkIbeKHv9UDw4IXeqLo20XYqujs/M
aeOglaghpdHGY1eTC0rPUOd+ntXpWMn+Kecih1h9Q8x88ntOiy2fDJnHUKtj+JBD
OW5739k+6NLqHLHeX8W3t2E6mCXIlfdeo+vLqtsAm8BiLrP12Hr1MKtmZvPMh4QS
OLa1hLNcOsHa090cb4PBSmifq4tYebXZsOjydqWft9ZXxNtNl/CELDgn193UYUm5
j1+eQNnx7qcAV3Q4wtWzP1ZOvfC7dUaNcOusciGqna4BS5wXlx5nGSnnGfRMJZp1
GetOB/CcMV9bnCizeDdTTbIvh+LB96602CkcJlmHFwZu+B0vyW3xDbi3FaKXQGbY
+87QQJIB5NlSQwwcH9foedPQK0Scd2gu0snPp7N2bjiVM9yQO0TMPcCf5iGu7J7m
LfiEUzphPXCe6VX5sltE1pgkbuoMAKnLR9obzIimNOzFU3ouSLgxlV8mcSykeCX6
7gcF9vLtVWomG6apMF8/hh6ACwIuya64yzDjyQobc84TWY0Svr3KJXVo3jS7dn3c
yNA5p99Zms9D9maV2NDtTEhg9rwUIjJSGODr0uJctFOrXbimIsfmlBkleiRU56vs
dys5yMmO1pQIdjKFuqWhbd4TmSa2XxoD/MKAYOm+zsQZIc/oFWluBQz3aP2ECuMg
9+HmUPrpQZh8gD3AbFlRB172vmMKhbIrp4oE5n2ncbzVuwjWKfCiUX+zM6scG/NT
PsJg0wcFh8bYokLnNqCwkL/M07R4xspqDVqjDazr8sKQRv0dVqRyHtl/T6rvgQdp
2Ce22Uaf9fFeUliIxZKOKni8C0ixsiB3WClE+veVfgjw8UHnKppYHOpW13Z5Fund
Qy5Lsk3Kw6KvF1G7LAOhBEZyfSalfsgGbeuU/ctcbsZIeAvBjgDQXNPVB0x7R1lT
df6NuTA5728yd/GJbfWjZhr9aB9re1hOZGLBeaVHvPGU4wT65upB+KO4Y8Gor9L8
FkQcGxtLRRbNiwYfIJbQrR5h4e/lGAue+sviYjvYufKlg5ZzDlxklBq0AwP+oxEr
ao7XjbXHW5M8ML1zG9umOyu6PrVCxEixu+k8aCerlTpWEME200oDb03KaguzfD7a
0ETuohFLffLV6Emvl2Mhcqk1aAMn2tokntTwkndQ0pggb1LMj8QKhKi1LJIGy+cJ
ok4Er5fSoecEQiWd2ihhLFQaWIJP5oz3jYi31VP+4lLOTv3beWHegDANkC4mMBRw
7rI68T06u7SYVWP0J1A3qi+5c8ZeYnFuyEW+3k22dzJV5U5wAfk5yIpUcbjn7J0w
zQPYnYDU1jf5I5P92htv5RyPaOSYeJ6ivx6qlF3z3QenVB/iyeA44PNXR4sf9mSm
59zStLKypUJZRbjfIir5ZjfI0xg9wC8CQ1zS3dgbQRV9dsddSsJq1u7pjjP3v/At
xGwM1hKX0YNzFbR86GCXGmbsD92bJ7+mSy1XN4QaJ+h559TGV8ITp6klmnOcM0d1
nXB14DqtRnpRMcua10tGU2QQh1tnv8vN1pEszfa/HJ6U/RfXNsOOAJEaX/T/0O1L
TAmjkVKKkV8+RuGBKbh5AuLUTT17iZEFKWHBSOwtDgiWOO/brsaAI+VhRHvuQK/y
zpY+sj4Py2RnuOyoWKEC9rGG9pb5WiQs4P7CvmJ3YzuWBN7Oy8zlkibh5kY34ffh
I0Xpr3ZVg7f9/VLR0U1PFIbgUsW3p1IC9HDF8o4btRT/+kz5R/84niUobqqYY/o/
WvIQAORQqKJoi8gnAYviy5jHG7LLyriruc87eMOmH6iznYhzyJhNW2E2HPOu6pPT
517EdZAFhR7IUrc2mIUtWQQ8cURqjnrN5MfQvGCAexn+DhdaLe2sFf9c8q1Vurqi
I8hU+4Z1+F2qUqHyh8h0bkbJ0tMkH+T44RtZMOrwOtNRT+6BCQ9c5i2274UICSuf
sFXyxcm3cSRTtjLiEMGSN+CF4/HJcA2ICQ8CkK2lMkjm72vcklslHExoDYYxfPn2
D8dSJu/4ar2Eq0360gHyKFmuHXhoJ5v+1UYVCnvqKxlGuQYHJXwWiHDKp55p/jsD
VlqBYPc+xGC3vM5OmOb5syziTHlms5KlYTx75qx4IrT58XHKZbZl7VNQIqqg+5bI
upYRi0RgAQhrGpSkf80M38ee3Luy/97IzktkwxtNV0v8LgchVpT3T/J3hcJaBYV2
VXeLm1tgqyBMJDH7elQXqTrJ1TPXNt6ajPjn1PrwN4DwOJKmt7D8blE/jLU3OG6U
VgCj3nwpJq080mg2EVX3pAhfvRcZcwIDrNbNKRG1KTi4fwThBa2vJ81qHz0Twws/
HyjD1aDgAyhpE+TcaAg4o+6rINVHdwAFumltDCVIHKN2xOCr4tDFE3Uuaw47JWMn
M3MxvKh1aYkoqqrbXjSo1/6yIp7uslwQKMOk8stUcMo7RZP/4gUFb9oLAPaj8/Ki
C9xIXtFqLq+XN6fXm7+KtC9Y17vc1/0YzBZ9X2290TIBDTSEdqQzRzE5wALFGtMe
AV8qFn3qNpSWPGCKbKkaLaCH0LO+t3EgOna11tXZcvedKQIR1qVVua/l5ODyjn2R
8KEzxNHWnamMj6GPqxto3yYCfK9msW4Lss33o7WbuMh8TzJpeYy/8OhFBaG8KGE4
DMggWlvYze3Nd7jkF/kYHG3wtUi0JTDuknXOaWrEaROSqKVwCvhDiyzeW0jiOLqu
ZIBnKiwnrmix5pc7Ogx7BAl1s9v6tKtvaKPHAvoKWacir6r3M3zSqqWCWmMagiyC
ijSCDBbrxrbYqUgbNHRqKNw3ee4Y7xBlUp3KXP7Btb6ANf+VKqv4tG9Hyq5w62LL
dB0bsNSQ8E/RKREthvGyf1YE+Yx6OdGeM3MmQbPxZI0C72JoOwOQRxAGRgDUC98E
r43gJjbiyZrmFri3pma13pRHSmNDGr3f9DdXf89PDx6NpNKxCK9jw35/QrGZoBt2
uf4gtarQxHmGeLZMuXImGWOTukc6zHyF5ZNawfl6dP8AbOLdyEtqfFqfqEtnjlCi
IBZ98ghDqgz5v+cmNPExPmz/2ZrgH4zbq8QWlxt9kqUsp08z1Hsk2dbearF48gQc
jAWb0oWcn8Xo0sQjutgPbJ/URg1ZFhYha1mjhu4AVs79PPtJma354aJe7V0Fsmrn
YWjSFfPr+sjiSeqYjIKHrAIj7PJDIBk2eczkp9Ack5NczNVRGuV1AuVybetGm6il
iVD/Rp8u3uyT17aiRmtQ9qf+Qf162cKKwwEw377m9NNwLBQfcnN78kE6u++egXxN
QROfwfLEWKLnFQgB6NbYpq4EPGjilQYYqpsn1kkE2P+2a55rGhjxCyruwa5com7k
BjPsIuGi9a1Mb/fTZPUnQ1lnMvwdQDIrCh+Akp0MmEmAARRc7kz2jntwjmXVgtNd
2q1NSVxP9bgX5ff/QyNYQR5EsEgRhhrRx5vztNPI5Pl3C4ItM96/errsPb0/SrJA
8JvTn0T/CVsc+lEes7Xi2WulGdL/dknVESDnZg7WCwjfFxPSAbdQWr+4gYXPE+od
qTMsx0lUr4BgwF72a5lFdfOQvhng3tnBagdC3JD77CRjLhDRNTYb3xXypmDSzz+u
3CuYyIEHk6pGwcg/dHGjM+swRKAXTlMBspXQxRyuF/M+lyDTYGYhoHtF/+HGUTWf
BnhJTv4rQHmoy1oBShiyT3+AQZNWt5auHTztFN8zAiIc9OHDgsi46HK0LdfuDjiP
gGxM0hBCnR4K2FL9MRBsglnswbThHYyAsa+kb8tmfXdjJmQmJrGmwNtS1xhtRWxk
rFY8Q3MvxOy5GqOnPJGSAxQYybUJBZfi2tuuow04r1Y7tGb/DMw0wAPGVvxCCU/F
znMQWFIkZppmz23gu4w+tJiAFBjqnRJIi4YKvkvlOs0E7fbS+qhORNgDXmzNnMsg
Nhie0wsDntzQQ8K0ECqqpQ55PVQrL7zap9ulrVhePRV/7a7eVzMmwUELaSlGD9lk
A95eQa7Vs0d7j4K0sWjCblbKF84/aTT/Ryi5eppsJvKJVApRdWLq6XwzKBN5BYvG
bjhR6CLYYRr2djLFSUH/d8yOt9Hjj4CfX9+1z4sGUGHdIZ1ymC9eYAIZdd0DIaik
aFhzfYtff8QfEeRKWDxRqV9+VZBoq3hsMuDhJTwpSDXXIKfqll4DWpSjbeorLIi4
cf5p3/0mU+ruh/M+7J4N3v8tcxySuci5Tgdwd7HEm4W0rEfcGTj957DLkp1Fp5fX
6Xnt0lHtO03YHM+PgWSNOlehRumtsvovSET2PXc4oHxxdtlsGQ0LiOvinCCNDnb/
36VAvakZSK5Ke9h4zcA41S+EjU8sftgb048uZ1EM60AIEWmi/iLFdNDQABaKkAyK
r3EY5gEhAKCCgSJd8gZZ3zFdUi4t1mi4/efix0R3qHUvpeqfF0WUawxFu7QRyu9J
1XxOoBaRrXCke614otP29VxaMc4u/a498bXDT4l4qVJRKjNt/507AbeZ0HT4QE1f
S2rtr26ObkFQHJtUmkje9TNwhzxwMeau9tbpMRMg9Y2BLPljtRTTDZ2EyIKu+yCk
m67ZBuFTM3YiLCmv5ljix6JgB5kxrbJ+4c13S2WNf0RJDQmHvifZfJSrtInJgJfB
nsQde5RHewObPSwMZ46o+R12c64ZzqXy8vI+ZLtJg836LVlAxEWkHuDBFtPe/C8u
ix6qWkKsEhBADeWUZfAHR1iGPAX8Ws/JVPVAfUw1+v/3oWeh3LD9UEZjmEDFP51a
aG2E8bU+GVtJK7fuSCT6w0aAIzClXOv/5n/Ysee+nbcLhJVhH3GTY1lSnjlczDX5
JUpGF1fxGvIF6wj+018Mr+A0H++j1/1lNbgpL+jFFfP2ATA9BUZrK4H5YT6HweIG
S+crmgTFRSScnrGGdLVvvy36bqMysF4yUdWhVkx4tiK8gZUDu4bus7cYnbaADWYF
SmNn4MWNAk4KvIlKrjJ82GepkeVIydIPqHd1Ub37Qwe2L4WK4cnVEGvM7Wen2ZkJ
/ctHdMKN2Br+XTY1hg4q5OlUdOTeLpNdN5IIlgWIUWyDiqHm+rpXdKmccUXfff+K
UxvZbIVs5UDsenbVDkfzEisNzBJeZ4pzQ3dmQRsttKAUnSFUtrtDRKTChliQ1aWi
iYq6hRSjkSVxaBCPL4mc0tV3VWwK97XoskIvOtuHgjshlpJSSBm2GwlXUnKvxODQ
aqGjvNdkfOfEa5mnCWcnBbrI0ICtsCnHKIn9Barliuim+DPw0hejSLXYAgS7OO0G
DuuHbkqvy0lmUfX4Yb24zAW9QG2Bg89ZhX6BpxXEnwRniUIg72eHLg/jhashm2+G
hfnLkyvDeyyGU9ekhCxEokxKvEOjZQKave3+Jie/3yAPIBGAP/OiC4gYUHxY9zYn
LvQdeIL2iPfrtf9rJAytFNglYqeQlFKtNMiDJjEBketzDRFerAsyzU9nqjJ7toM2
bn5DqjWlF0tLeZU1fymXy9yYiMAGK75lxz1B8bNsTvadYOQBMYWjauJBqyibDaLZ
iJaKZkoqymiLsRCdUzWpovOiFAA1CGq3j2LRAHpUoic+9pnz3VpVskxoJlS42cZO
D7DtE+P+nGlmG+mfmkKCtqWVywNUahDEQgaL5F/vSqWtPPqirXqNsPzujybb1eRi
z6trpW8PQYirUa0e/zvIRdXyBVARAneLDxuN/W4nrjj35WtqzPRQZRycC1cT3SP4
k2WmhgQHJEhExahleMZotZBRrhFy9DVKn8KG04x0hx44An9pV2Wz86wclEX1G+Bw
iTKzYlc66qaItOp7ucoP0rBF/o1EXhaZVvJbEAMfCbBGLLwOcWewKq49utNyJ6bB
DIn/h3IwiidxA10OzNaAMiN33tu4TUGYOPVH0Qms/z8oJGcdhPKuJta692KHZEPV
Uw220FviPwcsjd0ERC4xgE8nnLMH8j0DXkBIRTmKf/N3NgvdufkzZrDF389ZkCbM
3XgmveyBxeH9dF8iTcXH5s2uD+CoU4VEHLRvTfQC1oUB6oreJYF5WZUV82JbJ/Dp
zDeYCURDuAPCxg0JtBEUq43XRcpqYHcUS873ShBiy/K0GK1F+oXk4UWGY9SG2GCu
SqDZWuFVcZLKQjIhgbt730iE23zEYs0jrSlIA9E582dOFi6VnOoqKWVGYQPQ9g8A
ZiMF7cDrrrgSf3Zs9G0TDI+UNl6zYr8UycdyF0S6LcRsPro1GOhYTUrneIJ1sMuv
qyf+ae92U5a4wqZR9aay9MnBM4TVDo7MGZtG5fO7d5ETRy3Ivbs1RtTV2jMEhQZy
SszaEl7pwfLPlB7gIzsIihoipJF6V+NUIXT2/HJq5MedMlXGFWAlgNvaz4jdLvMw
wL1umRWmJgiOlG4NvxEU5DXbftLN5Gvo26eh57CEj+jRFhDl4r7DU2hfc4wXzouU
xoekTjoUhuxjA2X6RzA4Zl77FQQWLjwILUlcj6Gd56C52APPTAr0TOxwowhg7Aji
igBh2/jxGPY9XyU9P3kPrvlY/Q3mrtZHQlWvGZL70I9MC3ateBLmyD5Bb35HTPL9
Ip6R8a8SP4Fv5+kVutSUwHb0P67Z1NHKL3ZEv6A7/E5fDXrm85WaLm9r+iPs4TOL
2eYEDgSXl/ITYMMdRhkxUHLSrOh6CYjDt4rPO/lJ/8TlfOpl5ztqc40ErqRqejon
T6iVAbQ9Nd3EU+HYKpIE7uP/+UI7E5n0cQNDjUH6rllvhz1BGjMjJ4zaQvpSWXic
XwQJVtr4GTtosKgKagq4xv/SSLj0H8sqzv9YrO+E1xcyChO3KOYgeYdXPj1gB341
dGqI0cmK7ZPrbUhaFKVUnBrpXbF/+L975BBgOWobs+OtHNjYjRtOgQG+WPWZ/TA2
om8DOD5jFqK1e3ajMwcfGQdv9W1/dP0RmDLmwhxtUOzCmncWoctQzssh9GDqBK24
Rhq06TPVNLoPAkW1OU7K8sZd/yhPdMCr4QRzHCn4RkYJYL8YPmNYmFX59ethUNRE
+xeoucMdD4X+qvNHnqyJmUPST+FtVwwPg7mMOF615OZTQVv48mDFLizzi2uWdYZS
tTuWUBwjPZ7WYUvZcE2rAwMuyD0fVhux68ihN4hEYKSpqdQrnjEB0ARff6v4EVUj
s7dSS4irMPTlIWfrzUUUoB+nY5V8c+ODeJbPrXxyus5O36EbX4SZX0UzKMovXzlm
7RuPCgD7tK71IVa+am71GQK1ewFuScDx3HBkdCJKvcY8e1GWfPuj+fW4so6usDpE
Mjwz8qos+brQZBZziAdqNcmrLSfKaG9YjKMPy+gflTAX8+opgDptvRWDt1mpOkeS
exzzsd6f6oW0qwXtEjuRB1tZFLzHc+nvm+yy6PV3ceBsQuwRcaR9jfUaIuLofi+o
E/sXbI9J5ntZhpGC6pnnES5Q+ujFpe1te66TjnQgdtg+dJ0dPjDpjk7H8Ni7TWsw
nOtb4tdBsjBxAPDuAAjGCGT8rAvfOtlnF7aB4zUSFPPTkCgSSwsmfeCiG5GOI+lV
uEXdCtfh8yykYADshSn31dySqMmhjbTbbPL2aHtrAM2ItenDu9Xg8KJuMZx1iFB7
Do/7fMYM4G/Trd1RcWVFam2UZT0j9LGC8eeMuUCeK39CPEMUo5lO8rEixTxgqsBq
o58gvJwyatx5o8BEx/nQQEDWtGvYBgLKDZpHDaXEkWF1mK7BoS0MYKpMwXQmdIst
n1GLpCscGWjVZAFgOYPo75RWA7yNEghuoyFuTDx9Rf+IbXIEqxH2yQVMyVJ0B3iP
avYkTRmZWPJ7izKOwxSkD0DtnS3CPf0SXzytMzASp2e/+TBQY+myCvkqG1fds0tv
N6gyY7Khz22B4HfP4gme1yvj2WTlIYK8+ufXWkQWa/QUn2dz5sTyevrZ+w8FimH4
JsgE6Feq4pry4HiK5PWsRu46zlPG7/qUCNF5mB+CheeRu7gb8Qa7kB82+cD2tkpt
BHn8NGbQ9WqaRGO9hFYnn1WsNFCf0fM6Jz10YFOAyIe9UZWZjPdEHoaGo8AJArO8
pL0BOVTowJUIiuUIdtHxTNi/1Y4kgIZgUx9GPUdh4y7x+pwkz0Z++QKSBI+JeV8e
UG6Zj2cQi2ovkzFXCUnmS5gHN8ASXmnTw1W80kO7RpSWr5sD3g8rwxbPZolBlImN
e8yM+35jX04bvQs0PyaaXyMwWhUbJgzkqGjIdKUgSd+3SRnlnAY3GZXz14LaOrjo
LDeMkM3qSNLpMY1BQsiXVh0pg9EVbQOqWU6uZaszWRk+NBmOtVedHrGa6kTmGboL
8NIQvFFwxhAweck36AydIZkDz1jyw/zY5ng5XcImhLp8t0w3l8L1GvKDbFnxrMYX
bjEs4yfddLGmirBZJWAeczk6mojvkZ4LqgXtr7e4Ofpvxj3bleC+a8QxbWMrwWxn
wYsvSF9QLA7Kuhxn4ZrUqSOX1qfUfc0HlE6Ddgzvxz8hixalhhPBasNvDqKpRacI
j1wADyEYOFpPiJV29p8Ze9TH2c9glOLX0wntpN8tkW+12bixFMHehTt3QiATX1JY
HmgfrXE3fyfGaDOkUIagddfs24hYyya3pgBeQDYzDy8FRjOex7QGPQiXzrtl4uI6
W/iOhN8ABMjEa9Fl0AbBBkZVABf6arNp9sUArTebZS0s17LDifxU7Qe4gfh+mYIm
oAv4FFkr5wqXLofDOrQEnIimpnlv4KwhdTy08b5rmPe5SqnoRg40fIhf/iojK7P2
TXJy+4fnoE9/GKHBFo/T+fdbxbz8/eFFf6VijEykSW7dxCgrru97S0NW/4y7mM7l
cMAmJCQynNAkTLSoYScb0oQ9kvG5fDZhp7a3dtZUyj9KnSXM+QOXEo+wUandkuhY
JAnci4Y/WtMWaYdiE0Gv9SkMtz/P5NTwRMjicsXigUGWQpU+bs8Tq6mr0kB1KXqj
XUFZkfNbdJnkJR15lrVgTGpWSp0g7LTc6towH69rh3dXzgrA5BiFuj5HVr943CUG
LUF/rrFVUGGpEZKDyGk+f9dHIM+RxrFg6OtTWc440aEHd0kDU4XhYu/ExGGVrD9/
s6Ksy1aIBBeSlaZQDWGeKu8xNW+QfCsz5wy6Jq9pYc0S83s5R2ZwTU7AUis0ugc3
Ujf5YqWV7bjuUbOKg0UEC0mfs4XiWSB5rAusnDh6lbdmiYfwjjDMybOhS4WqbAek
/xLSr+itTquM2joP/g2VLFarD4LR9PFf3TvnzIUMJc/ChLIMBBtJPwUVcRlJl+6K
qkHAHuGFvIzNJQtqPjTvBOXHv8WPGUTHU3Juw4XIVi9innS8mbAHMsWTGWYdJv5b
bq6q+yAxAJbIXInJdGvtcak+9hiQgNHEjxwnynST5lM/y43SNBSB1W70cOUJ+eul
I16HqLu8rsDC9fAYr2LljRDO9n3qJiSOpGHpH/BjZHqTiouPpB86bI7oAx5u5p7x
/ABD2OMnp/hD8Q1u7VEdeydqTPosscIyTeny2matd5WCpBh2DVCiwTbE6UT1DVaY
4dXPNZs9xJqR2BwAZbAAJbooDIywPnC2yjsQ22hQQAmSBoocLeGVp33bFHAd5cRt
dlON5MxQMWssTFr4DYaMKG1dgW9wG6IhfpWeCwiQMVxRkr+j8YU77gVRRP+Er4ql
fztTXuwFldDta3W4MKr6bhiJ6nUsV0JSSy6M6cqabq7NoYCl9jznNfFRAWa/BtZa
fDZlBVyzspowWo7LNxQuyLTqIIUEtCiyiSZZ3glyb4rZBXVgrIE1hi6xIeSo25yt
lL8MtOLbwYw/9GSIqYPRwp0593UV3QdC0I/JaUbhh54bhI9FaNs6esx+2IJ2FyTQ
rJdpwMKQoN5YP5W9uHsAU0La8tSL6si2qGBJAUE0yJgIdkbNu1LZAFc6/4EZIRwU
/4YonShvchHSm3sbcqpIt09wu13WYZ7OYWdNXVRwmI03ztKYB4+wWjEI2YUeJDtF
KnOOJ1oVIe7AIQqwIGfXpvXNhnuSSQwvsNBxhDWMIYZr/HEvfhyCc7Ht4iwH1yqG
2tOVtjNopGvMDIRDFa6zFxTweqDhnTylFqSUGtmHWEeKo3gj6w35GKQryPjWqNYj
DQoIjXIxjjcNL5gnC/hrgbOFoxhciJWYP3ulpaCgzImIc98EQCEnn1A1EcBGcC+j
16dMngFyGGUG38pkCQQfMyNdAoHy/ovUYWyHHdtNZuf2XAtdN04yPQGxlzfEiM55
QbaJkxC4F6r+jPsmrZ2CRGyBya20NK8z3gVKmWZC2qjdzVSs49QsQxSLkrsWnSAV
qEOoqqlqPa4XFWSQQo0ekv5LRJ2044BoWKmT5NKEpG81R6z0/QCjqOYOXbS/w6N4
CBWoAqPyZC2JKLaqtBf/847PSiTIYpHb9DZV7/TapJxfQumP5LZ8aXb8bNIXMdXw
bunzN19pK3c2NPUlcDd3Ez74crDuFOKQneAMpdnfkUaRGFTgbJiN4FOQtZRTD5vn
nnGT0fMTPrNDk/WrdE2t4ACSHGYOIl8NZL/zFT106HHlONc7o3JePOLOYC+HOY7q
bSJC42+BQjAEu8UCBG3lrbFRpfPhzJaSNqjuQWW1PEi6AqC9kUDhDlFfIlihh/mz
xS+6H9kzXNlmSBaaOyi2+8VRztdxT+va4dK6xSooYaghycdNcEvyeTR9XggB8+cd
aNWwciFdzmZic4qjXQO3eeqx9cl9JUk15hd5PvhKA8+5f6D1t63kSQhGJ9SpDUiY
Zklz5xBw4+SAI6au4TQiCyo7SMIjJCetBD1QVSCar62Ub9dxf3rU8jYX0gIAf5DF
gxDAlinmX96J76cdUYzn3BgFCqz9bXTtuvcW84JBTcj2pLpskJ6Qt75NKmqOvvpq
sd/CaNdbWQP/aNNYZAnAKA4TxNxByL4OqgPsBsw4RMBGZsJYYvf9Wmjm04Nh2xSg
TPTmS72zL4JHXgfAHRMMRjWcrxKCnzo4I+XqA4TnsBXZVhPrzNtv6t40pv7iXQE+
XkPehDtkE1zgcEMORRvt5+KeV7aA8dE5ltw0WCic0gB+/FNdjCnarRfY+QjgAzcq
IPLwZrYE8dMmSVs/WmYVTbehsWCrX74B13tGqVE0SCtD8+cDmO7ZHQ8PK+gV9vM8
6DHYg2Tk7BFDzFzSTAZgDW9OfMxUf1fQpcaqk5Z7Fl3Y8b5Nzv64F87AcVdyorme
rJPtTZPxiPcE2G2z5ORaeajs58DrPqeL2nbsVFowvBYXk2be14EazE+q+nnduCLa
ddN77OdC1hZ+YXqwNTqS5OWRTcMaDdvYF3DOd1Jbese9ghBMMoys72rTdKTyX78F
IXfYoEBFgBaiEUF9kp4ukL6gJTeFXQrxfn7LISNmoqydi1h68fY99ASZVZmS8ge/
WOx/JwsJEuphvTadq8E0BKVl5rVG646S2DIp7n/k0tbh6NCvre9xMlT5X0SbJken
oUOUQLE1iXRY2ilMqi6223LKAUqpRowNXsvBeDce2HeJpGlUvMJZUeJkqxjcSy64
nkRJD3zqlaSxyZMdMZWmNFUI43JLrY02QZD5Fr5GFsgEpX+Nuxb38snpZckrMkAH
fCAa/fKzTkKgBIfti5sRV8XY+azVtXpVJ/LWAV6OjmpLkQIN/pNhvuTndSpJ19F/
JXUohXuR6FGzf8Z4xMY0i4BIllN0+HBygH6D+z0mOOohuMpIWBdUT1YsmmxV1Zie
H44pzTbuYgpzEmtGu4tlH1L8WWMBACauepf8O8cz+G7yyTZHs+DEeO+9KuDzskdn
fR7yFORJujxCV0WNJPxK/++Yrm5DBX1/KKYTzy0hNDrcnSk72Hnb3N96CUBZbbrn
ZAg89Go4F6u8WHoEzaiG15zWiOQU8G2qX7YVBFXdW8RPFWRAe5Q/9lHltUYg992I
tZh/RjT0xvnd34v4gPqP7V8BUbeVEZss9zeNMpVfj/Q9AqRRzihgoDKqI2EyXfGL
wdJiXVcnjPqgWQiPPd5+r3bqao5zF3T3LC/i4dG32i2N7SRSspm/zSaikIS4xkzy
O5/Hl+/bNSPz6XVJ4RvgzNbrhyT5ccvbTGaz7UK9fc6JQwyWi95aFbvAzVVtf6Wn
4GL1tvwRtEbv8oWxkJm81O+x3qsnpyUOYExNP+3S1OJw8kwMWwz/zAUnzj2FC+x9
jFkyseAWLjocr+2+ge95YMyjOW15dIM3F+6H/TPYNXAycoEIWy0RsaHUZp0NqAvV
qvInIeM5uD2Zg//E4un4LbIievJ97rbm7Wk4XsrzhnyrBrmFUM/FTJBLhLvJ0p9n
/dUgFM3s19/xO7HCUm9FhmCcJDO6x5J205NEFYMlCGAaXo0Isi4mYtPRiE4OZelv
SDLdxjF1PphWx/ElYoR1E6ww+w8CJHRRW7CR9xh85w2Og8ZP8iUtz+iTMiigrZmW
dtQ9VnpOPFuGw2SiiCS1KME6YNiueS4QtyJP9cxHjmT0cLmCmMk3XMQnCaEGSAcT
3ToMfoOm8XjZJzDyu88AOUqLpbzgoota4G4d4LCKjDIJAHuKODXtd3l6U9mbBpZ1
W3x1hKiHBOCivEdFUWSvOTCYzAZm1Cr2OrTEGJEQE781MEXuXwD3J85ZQjX5NCGq
kG8AFU+ZJWe3//cTP2xXUbz4SOwOxwtpTFhf/g7Sle8RSi7ECLpUi3TCRAdxW00s
nntgz+8GcH/2ohn+rfamvNFD9U9yQLfsLuuFEvYfmMQIuamC367AU3nMguek1NA7
B/BJO6BlfK1qxtBq/c/lsoc4piFXqN4nr7gQyEpjXavPLKmE2lzC5U226TuiAcZc
C+Ar6JoepnCySgeF3Car+wQJ14yonsmiFLNoD2hUP+Cuf0LN5FiKgqRWQtRv4CiY
KdbDWdFiAMeOBxvo0X0zbadOz/uzZ3gz0JTqiu/ej2hDfziT9d072dsX9K0gmCP+
1oQUlwmXD//hSS/RNz198DSo3iNPmxfYqN7V5GS5L6cTIDAaa3juGEk7ZekQLYlL
l3pxQSfBvOuJxpe+8Y/z4PyajwnxVJQ2ZvLKQ7sGdzccSLXdtXZnMnTqndOQRajJ
+W+z5L12nHFERN7b3gjvOQpOJsKhM6Vm1Rhb7uhosMgoNXrQsjIXvJp0TZ8krk9D
3f6ZUXCkfQjmw1pnX+U3ZxVAiAwYJvRpiyis0OZoRBCh0mtP1YAVpmmD6Gt3of5l
CPYWdD3Ka8hIp3YKxo/5mpZOMMltbAyADtWkUVlkYY9USAiwlDj+MRkoELdnalMm
r6ny7GYyLLACl1qwcxEh+CDe2Gyovk9X4fz+8TuBOiXHK/k3cgCWczr0lG5A1K7S
bWEaPC95PBipL07v7Ez/raWQJnWhejcwZlnWSzetRQv5WtN7/4PYMejX8F+R8ZAj
18/tOi5w1z7xLHDYmTBMZm96//DTIfn4HeDGdgQQPETwvJCkoTNVud4nw+zKpSJ/
HMyYI6fKWjFq/ttS4oFBogeXjAe/n5aCDcGbKZH1bjZt4utim/aAqC/bZTutCna/
yCQzkIMglw4dhtMCAR0cE+Trj6H0CdlexEzMWy28gGqVFWVgP7Cliqrs0FzBl5in
yJky7Dgj3zTDD5+GlVBijevoNENiU2x0U9/2wINh9hecZRixqPtJyOwTV3Fab9D7
D3MprshoEIHnQszFb07g79JKtuBTddoKc9+CmrXu9OG7iaEJ9EXByA+3vxlce4NR
rkTDyBjFgf7M1l+q5HoTMbINZ7Q0dZ9ombVLY0s+dLwgKIL7OeJJNT5MMfoY5V+4
UzYnXhbnzC+czp75w9O3lXTXBOBCFbZyyJfRwuQgc3AiYB0tLV/xTyoyOkd1r8d0
nQaSdobiqQBZhDgntzPDFoNhWnrwMiEd/PwDhxPrrYtcNbXnKR+fp0lK1HUUcPeI
Pqyq7fQrqriuAn87bWAAaii6RxW0m7BOvV/1ffcxcaHAMhpdoyJ3xGWDPLkP+lQ5
vH4nwZsC3NwVdM6rqIxS50XdeIrl2TEaI5PEhaVKKUY3KAitrHQKXCw81pxHDP2Y
HLYUesKy0ACNw1VAo4++2qMX8ZkobmOFy29Nr0ffivegBid/SDmd1UfAjXClPGoT
eAb0CJbXGI3EuW3UMnNhi4SGJvmxPSmp1iYSIUKtSDaSUsesQYJbyXRpzzzrNA4P
R27sDYVAbJOY+ipFghFpE3kMHjKD+OOYgKK8nGKEtJywlRgBrui0fShnsqGx1tmf
iZBr6B176qJmOZVrhk95XyDwS2bVXyQG+GJNXXkBx2WLOTMirRrIHbxFuUMC/4NM
6mTiu0UQbedE5b6ZdufxFUXuadxoLW1QSx0pAKzChjCM8QlAPrCWmTVIL9E8sHOv
jhGPzsolTMaBRgokF2deCxHvnVhmrV4lm/LPGfTlM5DmVctPC/5Jt9t1HH/X/SmC
NOIvT7ZIAFQjdVymxdcRReZxplV3JA3E4MwKcZr0gxMNYYQRWpOQp9YBJPS0uRXn
z3EI4r3vuz36t8zT4pOQFNIc6ygYcUyqoyLvbsx4eufEAajhvy3+pbj9kALNUBS1
uNPYLPvCVc1dTh997lmXDRda0jyNm9wNNKgfgeTaOogkikqDLDQ2yXYV2bTfkTDh
VU8ac6StMv+mw2Nc+GBU41zvQTrsnldhVaJ2PE9a7IiB1QQ9wKSIKrFBe1Gbzkzq
unXnjEwrxeIX/G/qOSmfaSR6SSplKVSPbvAoYToWq7IkXvvJjAraf2l+FVz4nJ+W
ps4bbLaJXYEJ1nZR1W7+720aWIm5WVejonDpCkntlCZbwN1kcqFdagoofEDpQFNt
D/prRD7xWDQtqB+DdH+xFWeza4Q+q53lXnF2v7tHdhcW9v5kMv7JoJfskpIXdWJY
pPDNS4jSgl9oI1F9UfFlINeLbU/Kqp8BiR8AYqLF7Wmm2VUUze5ZK4YX1vZGWSHA
bKXAQbQXKs6N9EKa3LHl4kidRR7qzRKVtljGan2HU+jNotwAyZyzJR8ggMZP77F6
w6ycGf7r0fwvhOPdEbFiTXKarR2HpjmMEjNiqNsiU2omwzeDFXEIc6LL81NANvUv
holQDz9/DzaCfKFiBWoYPXW7jRKUiglaFhoo1vneVJ5/buJf7xwNkz5ggYzsrxKD
5XmuAF/w1+4x4LIRJCpqsACaFJaGBukVwVeabGFZf/0CVScppUHPodzAUyEEtNWM
xYfMaxJZ3wpy79daYkzCxu25baJKFjlc9xGIjR7aCjTuY/PYr7ZVzInmUD8ss5nF
AwViQgOJ3YI5rWHC/LZOwM1uLSPsY7X+klKh69kH7nIgSYGvoYrjq77lfjdNvh8x
IIKtpF6T3TE+o6C4C40dGx6OkXq6sHSzdnBBgmXOxRtGXVt6GslZIso3MG8aCAXu
kz1Pf/7z1AcMR2YKLuQGZKabcbFf2K8+fvpPAlU7NcGqPYImOteQnot8n9+VV+Wj
W8utcJYyREZYQcoZpdp2NodaAgJX452mJGv7WWBCTDlLo4pTSw7xNpwTrPBAtiXC
K6wKnjDQUS9YBp/+g8O3mBnJ2ouYuvNAx15HuoMkY73AKysDSG/uubzmwI+ePjhX
tVq1UovPApHZqJaiUo37Fqjq8a5+PYxo281ZAN/3ibFyfcm8hFccgPfNbNNiU9wr
cWrCFV78NltBu+GWalqU9PmjjNabQRStdbKxv/9x/jvLc8Og9JkLaSXIVFWAzYme
B1s8et3ZgRHS/1I40Tt6ckxU1YozEEe3hDgfDpbrF7Mewblyo13KrWodW5np2n9e
9bXiUi1ePcrr21+seySq96i5qIHQwfPIR3ny8tOC4+5IMrOmNRxPtlfW72R7ASEI
DDj/TZaE234pnrLEVKRncYtajcnLDa6bVMlHEWDuagk/Nvltc1JtaIAQFmSqpvZt
+258+V3t+BNQvvKemmvAVma7tsd7vMXfcST4vVwjjHqVNZ5/zYC3uAbwKOqPlD72
jvDT0Uy+11WItj+fz0HH4SCgjBq1RGp4b/ufbTQQTBtk6w0WYusmo2jfn90Aro+q
kGwpVBi4MmDI/kvpLFX6+TXrs+ec9X2zn4qvvxa6ACIxQAm9Xn3/rvsJdOttrGP5
EaIMwjeqrbH9etwSjJn37npRJdyplBwx7xOkCo35jr/42sfttw0abszX5gAz5Jpm
vW3GqFRgndbHN90WYWM9iCtyJUb6ajhfj1dH4b0IL0d/ZvGOZXJoHq6fmAkF6Uxl
317zj0B0NF307bJzavuNz54OMQbdXDWmhw4zn3qcgAJUfnrIWBRMOXEj8zW10cz5
j/L8wDhv/Lb9dPHSdcvgI4IWf+2uvru2ZC4atw2+0DPGDPhoa4r2EqxcPTWULSFQ
uLYjbt35/PvNIV02gySe35sNcm4SChElpVJFmtRngcOsUTlkxQ5YRjvIpwJdUhLV
/CstVfyQN+6uITwqCXDnv/QvoF/oMhYjbGkIPYDc4Wir5iWU7bjg7w1UHRhTWMHJ
Zi99994vCcteIfKgac7RMd4qSXIGlKuluIiDZOQt1uA8vZRJsTbgPmdbPA9tXxMD
VqW82wnK+0kTccng8UZmwI4gJPrslXhvZ4q5y3O0zEgNcaC36IdYVXN0ag5UbZJe
3KxQiWYC1lDFkJl/h1CFMVIYbTE01C86zQyMjzwx0LLC80HxrXmDgRD+9Db8cR5G
3pIDGk9TtlP/wJehSqil3YysNLUN9QUSME+E/aZ0ZSzVx9w139VD1azXVn3Hi65W
3lP8b8fLDTnarAIsrKAMUweh0x/9CNJ6eFyh6kipyn5RRPxOuC0JS1v0CHOwNSmS
Krgu9HR1Jum9Co8pjMdJZGMRwhJ1jvANer7DIF9O0kucAByp8uwQgTZZWm09gAq/
Y/xmrDnLoosL4L4uZeNuqWn2r2fl9Qe2D2Vc4W6eLmnDUj2fRRZJ7VXV7qQHll9E
hImNsjGfRLJuCEeL2BOm23T9F2bgb6uSYjGVf5xdl9eiVb0jEccLfs1WtKqT9fBu
6Mwy7z8a8cRFkqo7Fxx3Lib98uIUftcC/JHtezf/txyRNp6Di6lUPukdy18WwDdS
Jpw5uQIjlGdfzmu0yj/6p+RrmWaU15gyCZpuXbLxtjI76XoxBXuWrbRNR6MWFajj
eiN4phd5PONS9QCb+3eaAlieWP3aq4t2Ky9PaNXvp/cmgCTFC0+sl5igTYxD0I2P
J8931qkIur2jktLCffU+aeBLF3d3XPDO2bHZ96Tc72auCOBBES92eHL1R8SZVv0L
SDgbJ4fIi2zsxF6HgN4bpLVpyM/UrwSeEgHB6I8mZCrS9qlCM8kZSASP8pC4RfiX
r9JTFAfxaYuaVYqGMXB+muh1d4KqfCrGx7QWSV6OXR7tMUz2HvoHPMsAhy/R0iBV
jYjc2p07veEgyQHl9WJkFdm9tHVxqDHqigkOr8V8UYOee4vbm167lJlFDrBcrhge
J9gfpCmOPnrdLUo6ycFgjy5LuLKpvmTAYbYCwBduo7GcYoHp2llj93mN05pBE04t
l3Po30c8q2dIzIwoyhfG5Y7onmGRIgN1zV8iSw6uZDlW6hZxsKvBxH+YrM9H5YuV
4n+nPPGDo+O8wGnxlmBhtCWCoM1mcxeRT8AtrqKPZmU2qO9Vm36/zFYi3+pbypu1
EP1X0mDBZPTIw7K3D1XZc1IzITIIeKFNdmo2i5gK9wZ2CYZSKhYKMCMexqOOR+xZ
zjMyLiegbnOqDn6cR9dqTztO7LUim/9AocIxxXHE6U0es/FKOTubdN2qYGzjiPQz
w/HEzq5JYDGm93BZyn5e3YWWPeNqxZ17Z9pCq8bVPQYcDd42gK42RXkcQVN1bCyh
KrHcCZWwYf7jnZlbqCgcsryE39WkK1IvhiEznvOT9mbUFSxuZ+TSj3tCqqeMaAXz
438FIPC5jxO6s7PhZvEPfiWQ7TVyR1P8HLhTOY2u1Fh6eFm3bq3vLWB8FqIiM1Rj
GPoI7MvYKamW2a7CWlGYZ/SLDs7l5UeQ1U0WRKJUFKGZzgk0m/S+QcciiWkipqO1
bL0T7Fcd8BfVw5gcwjtOKFVxstjN4vOBIgmkZSGPp/t7CbzF580q++MS4cOEEImo
5XK5vyyxkfLXl5tMl+CRKCR/P3LwYf2ul8yUT4pZ9trGU8SOHhHPJzfXf5Jm14WS
ATLObKACDUJzc5apb/zujyCkvuinVPm3QEn8scSfmzTGjd9k996GXtd/crDOhZXk
3vG3aYzoyIdQfpM+E4ENNhp5ZKK4+jh2YPiRo6m4JupwGTGXAdwMPICmeOkymIau
eOpyyFJwnFi7DTavzDYJjEenFykvU+3PoqaMB2pd3A5sfYnc0mZsWooPel+1milV
cu6qEDispjLCI+oGCjXUOUSn+7kI0bajlTHoNs4Al9DW/VamoC/YHXdxKPmxHYnq
aIcV9MMnGxlK44REoIMnW3L3X/aVzMs/KpAAOe1CqaAAKLLXhZjUgcdOcp/pDQrh
qJT60nbmI32/XMe4NAKG9XZpIZKVtr/Biqk+TLeLTj27oB38tufxvd5oohdK8MCu
dRlS4c+qOJ4RMd+HznTVsbmNa/KKly0sEEgem+Olkk6AoVsTHISAaOgmNmrW1kJW
92H3xyxxGX2EJVAiASab6VH7ThazPUSpcllSqt80XI2lDAe8Y0GJioxgh6opB9O8
c21CELJPbdiB6GAkICINKa5YceyAzbCfnfuyBHHt8BqXG4UkQSmCHiC7iP8qzya0
VDiPQ/20TFa8xJbyMqQctxwqXSebZlX9ujbfDKNfa2EiLbiiEWTHDZwcx86RgvzT
OeTlZX4auyiR416/PwAA1LsFrl9fRaLkJO+agRjg6U6jG20Qu5UUuGbuzbG3CSzR
TXLMRI1TuUM7zhdlb9+qXFKQTVkfm6MrqPWmI8g03VqMZ29a5CxYyBfZ5xBC0CSY
ZoXvJV+wEj/6aaoyvpRyJjWmXsa364oI0aBGZGfaOMmXgpKffpDR+csJeMKBZ2T2
ck6K+155pTqmAM/FAbyK/CMD1odvQPzF8OC5PybP0sVWrllcj3bAxvE6AMR3IDzr
pLpz96TPYBQ7cGnyCCl0UTpcYwTC+b6hZMdjDBF/JCUPsfdjh9tAezsTeM5iX2PZ
dXs2xqZJigZ7uxhtojwuGxbJNIzaCAeTn7MQ7vp14tx7gxY1iwjc7JMcmbHrbLKl
TfiujySwpOrwlyYrOaIDCIXwCR4Z0T7hf2DyIRgZrSuYVpPrqXiDxOxMpFl2hu9r
P8FlqJXyIrY+vEup6zPKOCSBfG3cg31QnPyquzHc3LB4dgdMPkNje5q8L254CYWJ
lq+gkLHcRdcd/5CalDz0sd+QkclzQZXSpZuPTLGDu0YHLf4d48t2xGpXYFuwRTNR
2VPuei+XTn45Xi3rs/7YqjIraFEP+x67BCVseS3OnmEfkEQO4oKVgEIXdi1ZmACD
kmzpfBon+/fhynnZjUezBxAhnm+uYVJx7V9QDV0Iu2/43J+QAi7zuFGme098drSn
+cYMBZZBI/lOEb5nIUS/+YUnvfs/r2z+Z5EIyNZng46ZAQ2tvMWjUP/qmdpX7NGH
wKlJJdodtro3cKzAXKPKX/cK9Hvrp88akbXZPw5LNHjmZL8xRTGA+tIhaW+PrUBq
7OhENAxisKfCBVoUQO48Flb7oaW5GCOSCWMFsJV52jZ5yzjwRNWk/+/GJK6dvdQd
Y5YzshWhwLvUWZURtIf5emKiGnWB06UBuP1V1zrcJBXKwfwKONnQMoHvhA81Lj6Y
tZqTnLqUx9gVG3J8tifh2PB5pQ67sLub0NJMLfcqtStRXv2pd9AMVpGeBAmsd7lh
oSeUdXSPCdRDY1DOkZPGKod+TNKLDCgjlKMigwX+sV3Kd5RUbXl9u7JQZ+eBybxR
RO0K6fxhpvWRfGVau6WnyrHZhSKZ5P11c4JP1EOSNDeXmpq81f25wO+bvOPV2mQJ
IHNpUp+CmvU5+onHPpc1rHh+YRyZjYFXgxZ2CA5L9UbsAIcoaaUEVBYFwmN974Q/
G9Z8i/MnGAZgs7izsdyppsLslSGf29HjpXNUGL8P4qQPb85STBiYdiVpWCKLpmFZ
IiuAXNd+VdZZi2K/igi2oEVYF4TzpeOdDCKzTUhmssqrF/ow4sPFoiIPitk5v2vW
5qqJf7B1uHTeMYyDy5qCRt2ic1/n1DCNRKoKIEAEzs8g2S50ZwPue0LKqOcIZCEC
/VQPJGsR47HXleu4i8AyWet1pbBPX6r8Lz1rsxUYwWJdZOWw6Lf2mGgbSfHrOUV+
ywngI2oOWk/u4ej0mRU/RD1tAzmBGdCJgMHGjDd+2YcyVxitB0CChGv1JG5OV5+s
rJl9wpT9YjbF362jyXECtSWKglGLfXJXaGIqRQcKxaCBWFkzx44q85HaZM4IhABj
tmlNF09aPf7mabSjvkqczyQolv0dcIoZN7TnFQeH9NtpE1AzcvZkayQtifbGOBZJ
ouRpMSdMzbw8dG7LPSzOzACdFLrBD7rAh2vP6B63NaCYu/zDm6Jt9b+6b1JMQaQd
rFIvDEmHCt5tW3CBCHg2b+NzY5QgqDQqixb+dXpV7z0Og9ZwB359DY8gjyudY12W
Cots1ApaC7UwFlTDlf2gV/2OxWOqMSZ62RcFlrLPf7r93QA1JiLimPeQkVcN7gE6
WxkJGrXvOO5nZQ3+ZocVoCrt9/wkXP661u94rMel2kodc7uMFgRqytbkJ6C5rztu
grti95PG1ZRqrPELwEgr63K3vbJfUSldAFY7AUZaB0U2h0a2XMF7e+x2bcxwjG78
wtYZ6/F+lIjKpomljQh005TLrbTfzv2hD5Y5T8AsInjSWp4L78VqlwXPbgnwjuaa
eRXvUk+P+Nm7DDWIrIZpzvvPu3lwKUr8GOyLSjWgn+PvPbkyVjQewD4YTPsUlepc
9zRNbLVQUyE1G4C8YJrtqiPdgNZdu/K7ztAkmVoZ6iAsCqOHrASBGnUPz/96HJ5m
kX+yzL4qw8z9hhVNRi0jtnE+wYTVWnn55VXYig0JAWL3cLbdHNEg4OH4xc6F6Oyr
itCsQgN4VPDK9YluekxGT941pHwY8NOUSzMpR7tFmD9z9YqN/UbXqo79pyV/qmD4
jZrqlVe+xu8dTiKpYfmC8Ivv/BQqniKKgPp4wcXxSJnFFQ0FpexRrsVDNh1fzRBr
VxdQloNGEN+GQ0imOCSRVEBxTPwnr5/yQ25M2P3zcboUXDrdhxj3DDgA+2srFpdx
Wq28Xgapb/Itrtmgm3RB4hbhZU2aAMqOOCewFYGGoFMjhEMoU3EgIabxGyFhW/KV
jHwHiB2JekyUhgtc+SE4xSiI0mhu4ezw+6q8w1sIj6wQFJWZGX+ac6XB6DU6cNcs
dgkFifVU0wlS4m+lquLLt1k7XddEr0Un68Gvn1Qdqn6y2SbDl58GaBIz/VpJ/USQ
9l3H3OgcVuLyCJB4hPUaCY8+D9osW/34ncTAIPZHmv8+OrECLWo8IuZR5cyJFP2J
VmDmJPXxfvXnhR0OoNPNcwfYz6a3Bc0s1gRCVVpWNN5N82DZUmgS8gGvdC3vgAcE
8WZ85lvCueTeUXNbzqewjA+0REz4YpsKiOlVtJX5hVBXjSw1UaiGGgZfNe/lLKWG
3S8Plf3cRbkySyRR4uKGWwfYQO41HiMatLQWAzsUGwOcmIelNoFDfDBpFB5iMyoW
lpP5zEDHLWT+m3NaJjl4bQkN6RN0RQ5CH58MdM0Y7l02co1eLDkYONoa1QaG8iWa
SnP0DdP8AQ85Wft2aldjkIPlT4tV0+yKuL7TguVW6DecKdremE/2p6yPT0hN50PY
T/9sLMBPf6kIIW3IG0tV2YSBxZR6PNWMrUtEFlTnNPNaB+38R5RahQrZev1fMYI0
gzcJrMcYOmxK1UdhjE5lqDfT/tEta91Gg25Bajs+5W9/zmWpzpOmeX248l+enjm1
t/FqxIOJIwTbsfaRuO8omKq5smDLFfaqfKVgCmcWgHLNJKQFdC45sgD7+XonnI/+
Uh8zH/+UnB4SJOPJlvCt/pgC4lUagF+jIzroOzO90qDpajJQ6MJIlD8v34RhAbAY
oYVD9gt+FY8K5uJWmAq5Gv3LLyaTGmhUYyzx9GM8VV5c1rxHdpGnKMGyYXA+wQ7c
i1Px1KJGBzpH6vbWTlC2jIP4BuLgJ2Poan7vHPbd5BlJJFrvayPaYvoIDRzTgjKi
xYiw0FPK++oFeluKUMDpZONZj8kJ1XAoo6byR/8fjr29X8VNumMH2lWpNL2YJdkA
Q0Q6hfcHPxGDvka+4G4Ew618LkpwVDz2t+stBL+U3ir2782dcDgeJ0uhqrrdqqp8
/WhfSbdW12bpnXosbWhL0Vk/aCV5pGYmRO/4f54qYpxxF5ARBAjNt0RckfFjxEtR
Wxo72QkbhsbnytIfsX+bO/C8a40SLTF2wCCcbj6coqQjupNm+Gk9XDBTvB36rRQS
KEMH0cSdY4HfJMltkBLPjw8FpGSUKRwImJz3sqz36elI5joYZhb31Hk2ie14qp1q
7zBrBSl14x4QEi2Rc7DdLN+nwGZwVO8qun5H7t+aeaC9opy/IktH8UxrUCJdoA/e
EABHdifWalrrolxqp4TGz4EmOBXz4r2ViADujjFi4agDf21IAOEs3lO1lUeywXkF
KLkHbAx9a/vtjzBRK6aCcHcCObCpgbU4Me89V2wOW/bO9ekBM2v6zFzZdkaAlEZg
lyc+uauJf5scTDxNdL1ZelFyJgfgi+wmfPApNGpK0M8N7/nm9LtoRmOAWZAOII+B
VLZDXFUDuhztsVRc0F8bJZdYA3M+qWGO2Z4MPSQooxkjpHBT2WxtOwhrFUhbtJ7n
+XHKw4LfEYaUrQj1KaP9tbxor9TjM5yTqn8gxcZYSFdnJNaQgLtsJn5Rhi21YOXm
FjfxXEt2RjPB5rhhdv41zJ5KkU5pRo4Nyo52wHWEXCaNoeozQcEEu73GRTlyt4jb
eclGg987qpUq/eWv7zHYenBWmKK0Qa/tPW69YbsL2RQohj9mv3JolYk0leZNq6Cg
HEO0UToLr69RdSDoDZryW59L1tx7+Cx087GeOwoIwK1IF7pfk/7w+pd84pSdn4aK
vgOwKX/dHWrZt3Gv174iTvgqcf5uLKZdUzAS5GQewL89CVIUXVtDfWwvsWoT2wnX
jfdlzHEHBi5/kqurSrrhLFZ/UPsrT3IQppIU0a7n0+TBuQ6yb/09J9gPGRpl90hS
idE45VOW7aIt2gN5tpw3GDPXr5te0y4Ds4zRxILFzrsKcyYyjbli5CPQiPAZAGcb
E4wDsU/Z4jpqRtKR3zd9ojcgpb2NKbPdOdTbakXO+uyzg4jB9FkVCUDrw/fqMHgw
f1KGnyvHHBMtE+8Jr7fy3PK4BowFTk6SuFhohipVweKjKiPSAOptFvVsMCa1kCUb
ckf6HIE5W441QbYNYrhd0DsgXTKanvVe7ySSorBAi2c4TyG4tpCPJ11W7Wl+r/gL
ekB2dbtN/+VU3vr2QfjG21HcPVaBUlKCJfEMpEori0LexLSyt75ng3AaXwByGpKE
IjireX+29zmx9XiVK8Yi5P6lf1UfRZphLY7SGW03xStKAnt5ec4BlSX7jK3XKlN5
Y6MFWECXDDRZKV7k0Rcn4cdCcgg6ilkGnTJaFVBLdB/oZWhaVTfgCaKFtGh9u0mG
yhxSgPRIXKbSZFSa/mMcYdVt4foWYaN8U1HwICRPqIVL+KhPZ54G4rYLN3/U+O0W
L9RQy3VXqeOTamHhohcogtv1pl1tYq/6rpEQ5/2clvhDOfReN5A4/WkowJuRF+Qa
ZTAOt+Ep/3d9xXLdvkydgABM8vcqLUTPMvW4WGSNAEYvwUobwS0c8r4rKhUxJbdx
kiAxtLBa/wT8qEZJ4l6G6o9/kuKAdiCzLyvRWalnQ8sCcnH4l18/q+Ska9WhYpPG
E7gxQNc5cV2YZWJnaUy2BVFHkYyDoP/h1NP76VKu2HMSW62rDT2Ov93c7Utv1NKV
PpYT2N6U36rtnM7WQrzDQGC839Bg0YH6AtAoEYrDTdtCI+V+dfAVUFXfnyqrGRMq
ewHEVf6Rj5OYk3pPZn/wiKXLlnwJT8s48PgODCiro/x722ngAfZJFaO7F4nTebHl
xvYc9X9mW2jgQx42KC51QKXaLOuSycdNnN9/QK+bvBVrDfQ1YttbmuRx2liWe0Mb
E0Xm4VpDJvop/AR9IJqudbIbhViCU1dmsCivwAO/KtrgWv6K5K0GMbPn99QORMo7
poTv04ZTsSS5XsqjSOKe1991E2opMDXOFl+mJYBOGMYfO7KgXA8fm8bc4h2I6qYU
l8vwt1JOEJkcUHjSIbVddw9lFUk7MGdo8txb3N+u/iNldy4bLlEBhaiSl2fQ7wKL
h3MizcNxYezt96wPf9B/2Ip7fx+gZIMWvBNpjEJK6qN0lWP+Tqq9ZGYx5/5CcWLo
wAoEFwxI6VkheHZn+Mpd35x+yYj3U1aIfIH4bgRjNaZW1zcJNDfq6uY6MsUJ6+Go
7bZ33E2t+Pg/MPKVaNzv70+tt0v/ZBEjgtP2RFHKHaasjBUNAJHBPXhTm74nQ9IW
/PViiD8xjsdwqhInqVagEq+pVPD5cUpJMKzQjVC5YCK+nGHuF/neh86bN6GUbGy/
jykBWFR4ieiCg4FFzmjWGRcuEucE+3vAAJ+2EeDbbzYzPJUGF8eNe8lsSRn3D4oK
l6/Y0WTTe+ti1vQMEWB6Bi9iA/Ui+V10FExZW9xJYN+Cg5AH9gO+HUw1tGFCUWZr
JPk0NQ4kPSVfsdV5/VH0QLT/On6P+hVdSSGxqnr9H/4aGpOYSuF1kc2kiZW4kRH9
i4kByFRU962U2Js7ILN4JnDikVhOZaknfIorlbfjDQd/QiHqyyQsDQl2b56XSTiE
/jjrPekMKcNl0Um7sQdObKHkOcAMzvEdH6aFwn1ozsQE6EkGrcHfvq0swRDEAhJ9
RJbkrMb6wXr8XU2bu2cjA8/WwW5sctBshbm+zO09oYOE2zVWEXemArT3zKhOK0vP
bWFcEa9twCKfd1vJnUw1TXfUBdKZsAXvJiRUnylepXVB60I/fzUvukfd2rPn2BOi
URT3jikWs+rI0EfTDge3PQ3PQ/nQPw5nt3q3xO2TbKXjn1wtu55roqS1DjD+laK0
MOsMFr24Wu0F3u8ULT1wV8tQc+LoPDXNSWzHn1i8NTvumwnerOGPcYK4l0bkhSIq
nn8S2+CsjGK9su+z18bDlJzWTEU+C3QUO3lQNkFw1Vv3jveDXUNvM2SZAH3napnE
0sHIkkX63ma31jZZTxgTBtWjGoifaMmJZ6PRjhtoTovnNccq7paOiBNMTDg+5FnB
ti3yEOsNI6BySNPSdHoOfZyuABQcfbiUx7z0DSFGumpk5KwkCa6amlCnsz/KNNSU
Xceqp1BkGBsEWmuyMHPGgyV+BYDKyonszVUgTEUNAqQbl5hZLL1LG2pM6mA6B3bY
pIy9Za375dJ8fh0JkkMSuq097QSIjm+2n1oHA9m/S1aOoJCpyYkUpLWhh2H9Dh70
vBzXXFeswqsThwV4FgcJDzS1Bqw9MHgSLYXNhsTu3+sv17IKJKp2NjXB7vBYfx4E
1l1xeOmhnUoB9II57xF/cBlg7cLjoU2D3Vn1BGULWBYLBSKYzpRVyDF7ypAhLYdy
NWhchTJ9LkJ3AfTbuuPTWXRtUONgrbzQQ2X6OnX7KJYa2y4n2Zc4UuWRY3FrHfsX
uRbpVYA4lutLpyrW+6kKyMJQHDPgdn1452tMZCacCrHuENk6d7Cs0YjgvJNfNaYs
bg4QegHgxWAUW0oztUrc+PXbVAmhbJFQHMvAKqow6+Znt3D1Jg/ycbLSXrh234ki
/0iqWpGtJFel3ilTLupiqKoQD8pL8OnXIwhnMQXqh9AngAbE1BpxkgG6qzzOp4kO
TSIsF04/wG1wqY/kZQ40TBvj8HE+/KlpFO4I+C+tjHAiCqlNlrQrz5BLuquv4qqr
QEz6llik4eNcfsIvXl/w+Sszyz4M51gJoTeAg6gLV3d0l3DiUU3+PcVulPT9jJ4M
e21nPo9dx/uzqDHpEfxCg9VrNipw7ytyr4JaUweb68+RCNEhEPE7uTNoQ1d325z4
3ier2lfRasAjskAyZZC8oNmYBhPAfCEE0U2IoTiPQDgm+xxNP3KjKb5wBV4y2o65
QeAgV60UgVVtQkjg+5z9U27nfaZKflxZpSzAQHQQdvhWgWcmQRhYUQz5hniv4ewF
k4ArwIG47Kz4pDgU8Qc/xRvoHo+QZiW/lOwVIZwIN5h+MJa1rtGGa4F57czwPlTo
nMAaOe2UJLFCANcw9i5D39hpBI3S4GeHEJ6rzmwzxVlHJM7Es7oCm9QQHE2Is3Vl
iQu4EmgntCnbufLMyvoDTk9T+caDnxslDtcKHKkR3AnuvKoaGDzB11qtSmXVyPyy
r+azlCC9kDkOpXuncH67EpM8b7h6DC7CGNZNE/ZrHWSwnxNOkZMnFEHd3LA6APSP
6P34qaB7sbXz6S46R1cD/DG8j27WTQClHtJs+MiTseSYOH1FsBd4dFM8S0vo3llv
D5z1zeiw0u3X9A+yDMd8m3GuppYRqC2K2GPmOujFE3e6jiV3cCyHSxc6KhBB130f
t/AHoO1YZCAC7eYeV+xvLugMZQX5AZZp+Xk5txf+Y1Rt9ZWfpptdsxe58HG6uky/
4Qk63iRT1LH6ttLc5hE86iIRBBqn3QBD77MpLqBlU7/XlU1dKKJztk5m0wE55byp
svScBgSPks2Y8X1zRZAU6uuvIZJviv19wXFUjE+mWMymfxcXhinqWXE7kOlcAAQy
MKi+oF3Kct8tFX/0xblGz7Dwh2hWuZKU9KKAmjjA4sIL9nPD3JjGiNv/UW2L5sqs
IqWzhVCRoj1Sb9MhBMYahCO4HweDHrDkHxuQYMjmVYZlnVyjQXc27+yGq/0Y+3Lu
YP+E1VHKXtQQ3SwZok/8RqY3FAX1o0+j+j9EjwAISorMYFV2s0KGlNJgYHQHqtkQ
UgPruBCA8tF+nGN6LcGeA737T/RnDG4NT6PU4TFCb5tEOeOym4LOim74yLppgCVK
eWT0ERmMmTcWv8NSJS8ths97JfHk5VytnyWd9Lvs3/9LLxO9Bo9YsZFwvEhXnJfJ
wlmtMeymRlBP7L8VThGT9GM5RB40qY3afaTdMqnHFmMdyODwy0F86xpHgjfgS3W7
C/lYZFSsTCDsUi3bacELURPE7LAjU733IpeZjCD2Idlh1FGi2I+5MrFswV60H+CB
frjxI6PkCSm6nVnZUAySJNv88YmwzeSQF7ocXJahH+cYOMtXVMMu6X8K3HjffUu8
Rgs4nflnjvRX4nzNAwYPjmUcWKjJK5mzNBgAZcgmD4vnN30K0kkzR26qN9TSDfXV
Po5Pbpmh5IX24z+ayvf+AgPKflc+nqA3fdUZek2I1IZD1I+y9syp+THrkb+q8/ZD
MO07FICeKBrBkuDB17mPEEHn/SXvdzvUj36JOuHUMEb9X1NMenaSq2YiUDzAOSPr
NmGI75hO48BjGTPGpFqOPnjXbuAiC7CVdmTzwrwSEe6HYcv3lr4FzuWy8wINLuQ8
IwJT9Ab+la/I9uwp/MWgrwICJJAooSsZ3SH7gCnCk/SJ0lGyfqthzyJXL+WtJELW
4zP41hutrc6kBYdwt0YNVcwUYVt9ynlkpEiQsi7mjv7riOxIVyizvoBkP/GX1QL3
HyNxMMX2y4d0Nx7LL9vmqpqvrPVI48vc9hdZm5BrGVJPC1Zw9SAL7T967pThvtp1
eJ587NbTL/RWm9Ji2e/BBk2YLTEP3c3TIQmRhg8aAZrO7DJuDGXdOxG0yycnCrNL
keJ6gNqP2D+NaGxVk42093hoD6A7jk0SVKwqeV01633+FoZIiuZOMd7XWQSeN1RB
IiSfLiaDVJZ9TVA/GNhFPKwuEEjUtEaqLAuh7R3jAYw3etJLK8Y7EBT0LAt2i0st
T1Y9UggBTFRwzIy5Fgb7TMSjOx+3Zwl2seiRQj00FM2AOGKWRYcfKOE1cYT6lWoy
/3+3Vvw7QfcdQSvUMQuAEoQzPXv5kC0ZO9XtKoCVfXawus8hOf40Bf4b5/gb+mdU
7kON1h0biAMl4esejWyiuVg76hldey8kMqFVr8svrMDQCHJej2flkYzuSuBra0iq
UPkOIVPdtvXKDOYxMRVSC+XHMG0GnrnSM+o81eDdqp4qv6vCngeVeKtyIRTXQZLg
qBieJwgPlibABqQ3uSS3l18IztsvJfKghxDe2/2FyPkO7w+iA/JDhMokT0sMUf7W
GtNQtnWvu/7ABa59Ha6pv9Rj6moCsES+Bsrej1O3p/5CYDLRwMvwSYOPHo9mj6sV
nRi8/9X/mnmbwvhEJ1elMrZjauQysmzJvT0l3ysfKUNmgIr89RzkqoQ+Dpw8dFv1
mJWi1DElQOJzmNzZKf1I1KJvjItwMQ8gc29YWe2Id1GyNczPlE6dZcy0dS49hFEu
0CxfGRRO73i6QzrLkgNS94r9T5/z1MXX72zFro0ClMKHINmx3Ig0MSKhok3re7a2
/d8zQVOnMFe04K+FzX0EvPNFo3TyKe1vMZ2iZGaHOXx/gapAfOINc+U4ZqkfEIRo
sc6cg9GpO+Y1w4Wnc3dT2LhVMbNgCpULaPIGfJi1eEGLkAG8NixK/NpznGNrNGNu
RGFuU/23GJwfiUc+2msI0TCTNYxtkiMpJgx6RG/H3a5VvDbt/FXDjJ/Yia2C+csq
lFCr7cby1ncLkRGHAvNF7vLD11/EPHtd6A0oHWwX8Q+sXRRtADjvnqhnpPFb1jww
K9bSnzd5TS71m+By2xYN3WglqhDMJiNxJYfIzQ8qjXfWvCUfp97L5546mXjmXQNI
/g91TkHEDb1Xc+5F1GZORhDp4kS6kY0MCOTYCX52U60HjPSBoIh1sLLW9A0bl6sg
CYQYR+7B6qR6kheznJIMkN1TXi/EQ4P2tOsHprD+yccmpYiK91XMhrYV6JgRttOq
+vkzKu+JtxUxLMsmuhLn3wUHbOuuZiyTP3+nEvCF5XQqekKFDQo8uvCwy0a4p8lT
ZOuw10mCKd5VklqBqz/bv4EZgwNS332W1poUD/MsdAE0FYUKYgIUq9WhCHBnJAJ2
cjWNg/IBqvqOnQRqimX9birRGuZI6ySHHtDai4OBZYiFAKM3EA45VGWm8ya9uSyo
qnRZ6fG7T9JvlYZRg4EWkn6qfSCiX2rFgbQ/ma2UiOL31YoDChwJWLuO8ox9Hf2R
AyEdxv5LsI7jxzKW6cqnDodOzPRC9/PiYmG0QjAP6F1+yNnXEbww8etuoWJChgON
WhRO7rw0ROxwf/7VcK7n1C3+zn/KZ8SsjxBOvGnbBTbPBBq/mqPPH7gzr3KedceM
4ocy5VSv1IP4+3nrxJJ19ZjSGjRBe87Ub7w7dTJembNaVQjParXgBsnReTPtGV4+
qRhIBzzwa50HavHGmPHnnw9upSCm4lAfNQq2VFbMm91nToKFkcu7B3rT+XqqX8Hf
g1rZVgKx30yTFRUnWL5+ft4RCgLyxk7hkGEDrGgIQu8wjoLmPB+iYEkJkeCN4vxi
/oTRJNf6gaxfXwsF6A4ppUC2zIfYujbi3D7DzMR3ioMLWO+q/iFbm5zfXjQoC/Lh
MEMgOtSwcG8cBT/38nWwXYxykKLXD/uq7hjaV/m5/Np+QJzQDi8ypDuw9RL2Csxi
vCmV7HMXbRok7blmAsJoFEP2aFec7nvDCNKtSnMAFXJCEKsjX5eHxA7aiwsK3A6S
4jiwePtSb4wWpo41pRURnMZM8SgKt/B2FbNBbuWDbmaL9v3LitRDloUBVB/8Mntg
IGVdxjVLDvKxTYx6TrT7H+GeRdm4nMDeLOOi3G9JH4RR740VX5s3EuTc8Ly5J6Lo
gv8B1SGfssC6BvIQwl/NPdT0CJxD8KTdxD/k/JOFVUPkOGEu/rzHfi/mohpWihmP
vBCnsMljnhF0z7ivs3p991GOaKNexUZVcGmg5HL9cogULaT88aRx0H+h/aWr4OjN
JAik+JejLu4IkleLrEkfqA22Qk4xcsS6MOEfQP4divbE4lLi5Q3dwrQF2OPqzWYU
eDbxb9OiqsY9rwLjs8VhaAm034nWYjWaUnvqr+7P+Rej0+Qs+RMkLSU17+pZrJMY
wTVvrQTJ0oCzuCAp70sfOpUEIqbo+dk4pQhmKSYAwpcgwOkRPpr0KE14ZvgCLYJt
4P9PW5z5lH/lLpCUQB3Wvg/EynznX1a4u6a3GlLKkmhkoWuFvdsOKQHA8GF+2Iwm
RxC2Oj+P7Mw0j0vbSYL9ee1hiSBvER0dl+J3yBIMqBHb3d7D6LWLasxY/4bLhmYo
cLjnXCGhqDDk0p/xjTllmUS2BuVyYt8ayAihOM+f0JgjUcME4jbzL6ISOufo80rJ
C0jdIf3QwM9e02Kp+S1gy6t5SdveyMnJD7RJgCTQPWZ2U/aJu6MA2dXBe3+988af
YyJVEyhFUWfo62XkscWKPWygjU5ZamilqWb7VXTfjw3K3Cj84zxgluUZ6w21Gsxw
o3xsbNCUlM41ZkD1DeR3bzyPSELMYkknB+GWRBYCJJtSsGITe9ADPt+60QSy7JEI
eXUMclKLNP2tH7YkNFKjaD6j3vzlEt6jWeGr1mZ4ftZv+n+lHJ9QfAzLICZ7/+OD
7FiONhckCWE5T5y90DC0aC/mO4QwwCZLIfqEQOYzF2BUAdWTCSvsoBMZweJZvWDd
tb3oPq4L5jeQ1S6HBkBm3UrluF9hVU/nsJu5S3Gunl3ohtAD8wXayug0aqFJOSzF
oYjzWgkb5P3JpyUxP6Jb/vwa0UEMSzNYwNZLUGtfp8TbISCLgAOdqElYVVKjSDYx
IMsgb1Q2h0CGwuk463xdF6URhTRSaFAZEkt6ZTZixoVqejSTtQq8PuPWBevUK1lZ
SO65nRwa6MbwyStnn2C18yRRX8yO+rWIt9/zBHy7uepmWC4crLngGWpgtyB1+RdL
21qVmt1DVuoLW/C5m0KSiulhL66RUxHTA/Aj9n6k6hefzG1Y7GXrGeOKrC0FsCcw
XEUPeQMm5No45ggC9K9l7p0zHrHhYlzH/xe/5hqkI6rT5k3/YMYMjwqd0NF6YASf
KQxz8tLtIAg73rW4V7l8XlQYx5sBBqp1Zl9w7mKDl5RmvVK42oFHsQ9GpEZ2NiXM
1MweqLgTlsyW6xJnMDU62dI7O7sETpZE+HxpdeChAO6YGI5NdF+62VueICmRPtlN
+tUMbI5Vh+DCDwYg55mYIzjm/5k5CFlMpN2QUHWoQw2wThoevywpXojzb3xcYj7G
PqTKyaVAD3zc1fBOBERoO/ZTL0rvumH7w4VV+MbR7OjNDx0I/S7+uaL9Qj5/93/2
vYdtSk7BEKLpiqE7qksvJGg0mrw/aaIrSSxaNhbBeYeNzxlvBexP3ISjBJdtqpYj
nD9Lw6hoEStQvSkgy3TRJWe5wZBmpr6aXjzGAX946BIgkwGwWTihJnWMobfzUyJa
Smmn9hxu76zyQfflsLMNOaIv6UggPjZ+gigM2n+9hcU2IglMWoVdYP573CFOs/L2
oUa36QVFmP5HuhTfXq+l1dXc2QriVhpOlCBlQvchQVxI0v0bcN1SJcyyfcNXPt+2
Yg59UhXpsrkcJlwOsYegGoRTmVn4L8Sk2K4NCeacQwjZBQSNsw+iSvckpUM2U8Ds
3Y055RybxKRUGm5q0ytxYeLS41BFzF6yZfrteTDkjCKCMchUlx7yieVTQ2wXIeII
XclGMR9uIrZse+N73uJNrhTD86zO2XPmrx7Wk2R49mu2jSmgdG7srrtfmdYgECEF
N5OkYuijx/suPkBeEeJjoFfCS5eqVN5rReYJm1Q9nXdLyvhP0jGUFSxS3XkkrTMh
ZIwutHlotv29MmKYBmvyjKPXsYeTGOXJXmonSa7SlcwB+Ex6c07P1Qz1hdcfaabG
3VyGVVYScJywYKoa/MGWVSs+w5/AB66S4zRgIn00miPIGuhsFh6pepIe8SPbFDwF
yOCuAF11xgid1LaZpxYJw6V+bxb/fT3IUKzYkNEzxXc3kqaVPHI7biJpbUjltl3D
XcPhzWHl0cup+x9fQuC0P4nePOFRLr1JDKvcxHz0MJ1hQjIvPfoWhqQ+/lrgu5hx
smBf6dqacAdT1tFiPucTcB+bZGMVZiLocUfkY18o8RWnbDG3igRrTxMAfRxoqoP9
Hpk1V4WGH2QOGpYE0BV+tCrc1+h6Ttyg9ovw8QD7yFtjWu7KcPHQ2hszEmF1Jqgx
Zbt2kB3MdtU7Xjxllxn2uCYKSjATTENOpovyWD9mmpzU3X1FB6cynpQFZeDeAl2o
4WEsmsUp0BxLBAiiKOHhCC6ncpy1QAZw3ALfWgOO6AmCPtjJv2tqm3JPx5KYDJqb
Yn4A39PZhXf9653vMseevb174PeXlrUxr3jFQL4QCUKul7VkBK1gEdTE9zJC5cpU
K9ofhFXuJJgYj0w6sDV0SN5aLwgo+bpogQxQaZJ5Ryx8FzW/+zimLB/VP62TdXEp
YfamBHV3VIB+6KTR2ASC7qnzpiyapuFXetFpb19K+FMnSSUEmORs2YlZNkg8RAB6
1qhGLS4fbC+8QZX23vady/SU8ijcpKKhjSJcufShynFwQc2YDkCR/jRbI1jzyrAx
Clr0NZ/OmfH1s+1kKJ1qpHq3PZuuZGQ7scTqvm0UsTI42NAU89gXPeSalG14Inan
UJKJ7hbYDoqYE6YBM9jCTOD3CMgrbToqvg5KAxmt6vN8w/hKZOaro0Klw56LE3SO
5wkO9+rCsIJULkn0Q0g6kL+qAlCPs3OedUvRop8b+SrpkeSZva5LH0XZ8FTAnH3U
FeJl+WN3lDIC9eJysnKGK5oQdTcHEn2Q1V/hz/c4NBmF6Xr2goQganThCog+N1aT
Xnic/csMt0RA1xGlNLNIMd3fSmhxulebbiaKDSPqSaIjwCTijaaCUlKkMKTFJOYX
bA1zz5rH9nEVH3/fxO2N5C3hA2V2cemecd2sEFBigPG5t7bCUNmLTQstKx75bWej
ukzqEkICQ5Ddm7GXXnNRlEA4eDUUj9eQFyH1p7RX10hcRkLNqkOB3hQQ6yQlBGh3
bAQT5YvUl0r92VwRSg0REw7yH6Ldagk9Tu0ptoHjM7gRFkwvOXp4MyYHxkVR+AxK
2yVOWjShPwKZeIWcBwOGqoBLOyK++4lLx7wOsaS3g7LjnL/dHeS/QI8M/jF6ROKI
4x5HPyYDfLEMYP5xP5/s/RlOJLaVg4DxpK4pHdkH1jC0DQWP8YvnpY3VJlBYBhAu
SJtlbiSs4ug3s9wbiZmUCnVju8cnQKBQrBD2yxSWOl5RM0Qax0r3BqwlZ4tleo+Y
b3ik27qpX6VWmscjJy7ydvcAncUEYVGixvmmC1x7dn51fCItaXnu0hCUpgwGjPXE
PJLTI9eCZvBecaFziuYAl75xX9gKiiE29+Wtknf2HNSaMyRHg1YN33pbAxssmxoP
AyAmxB/CR7lM9S+PKxauz/32RFA7EvCSE9KM3UQrxW+R11wWlmfZSnumYLf4RnRW
8WFFsA14682vt+qSltAGBsLZoh+LCAkj+17v36VFC/IkYIWsNHtcv4nukyZ1UilV
nps9W5Ae0Azyj7ZDIm3IXIOSizqDI/Upd8/6gJB4W35JQ9r2MYOcqwRyvJGL/eL6
ucKtPE5zewTBsA6qVApSH9Xsvs9jm5rXj0Uaa1jTPtNF38P2DUSWnJ7t5xAS0j8+
swYGEVu2q+WLWLMkDlOCLF5gX+WyD/pUWfdQOprkuGy/ISN2424uqMTyVy5j9xUd
L+eJ8GXkL6HFDCtML6gLqDqOQ7L5b8RYzqWc+dYtnlDR0DAoWUQF5rJ1XUO41G17
aOglYkulH95ty6tfViJQd9rePsRS48H8Ph63QqN45vA43GnPVVokCFPNtgc7OnsY
1jgr6qUPzRhOVJITT9NItGqJzsc9DJ+w5eYLsQytXZbos3uti3MhCpjFevGlPE5y
BkLREPnPoYaraWNrvXcKa0qjSo2dVnDSksGYwWpERuSnZWtJzVMGjXx5EqYWyBQJ
wDp3HNo5pHWoeIsfrCXbvlw6SeT+0AvGpy+AXgj6LcgMiQ6+VH+b8fMu8AfStcmD
7yUFGNrlbI09/NNi88VKRU1L4u6AAvXKUQjXsb9mU/+x0SM2eixTaByx6RRiXjGz
utOS1H+FTXuAzLlQejT/jRxI9wtbg6tV1VKJpKUNVcuKaDuXrVhq4RV1y46PTf7r
oSx8ze4GZNvptRbcTf4k8m2sdM3zhy9TtMupJhuLSW85gm6a8A/lDymvoJZB6xWD
uGhusOJcl9WP0m3RRcglZ6sKzHsGi7VPJKOCys/UaPa04H5uEcCPVAH+49OGlCHr
6jhL2YToqEKCN6h4UtszYtSdm7teX+xVbW1AV4Z6ghk+N6+0Nf2UYJOAqhoJroUh
NtzTgam85Ot3vPS73k33B4BFVDngNIdxmV9F790ULUAurcfKDk2dWPirhwJaNH3j
3Tnt1rnhd9HgQfCdKPhTwpzBFkc1fCZ7tJbw67ZkC+pUFNtNNDLdQmfmvLBLQv2S
mGw2qOxUqnXCsZZ24LfHrjXXz2dYUE9PNpHUa+vVDMJ9YqOctfqToDduSnbGVN8H
AMDrh+JtQtaa8guDG0JBo6GkDy/i1A5g3HVzslaJIgEZPYNUiF2iejlEs/oN0wGc
0CMjbbkQEGCHqrxkMJ9w1VeQLaaXdzFleBcvHlifslcllhLKMJG+cTRSCxSuXhg+
EVBXi/qOOfPf6jjxr9yyO7IdwmcPIVw/175KOch+ep41A1HpC+OJ7AdqvwqGBRrh
MQZpFXDxR9jWryTNlSRJ6JR11e3vn5dOnvRhBuoHJOujA6U6qMrqUkiGs5oLF9AH
+vWYxREAhPhd1KMB+30dUSj9saYnNnJEUo1Lb4k98K7mxLm2ozctEUTwDX6ajyWF
RMSx9NUb4PyRDS2NiPNkD8Jo5wdfzyEItdWZiSdNJr7pZhlUqttXalRNYoGlA1+4
VB/4ZhNqZNxjpnlf5ZO2JsN3cvvXj7coEloUewuytta5g7ILcrEy3SIjctcVJnZv
uu+ebQ/QyHClgDNbwTyfPgvW2bZo1BgMhnJeyLcsaukB8l+4dtxPt6J+McOfZ+XF
v1jq0zcqpShiuCs/hqRAtuH5fyW0o26cO9x6SRGYJG67sidBZUnWbpYIW3LbC3se
G5wodOz+sSbDsaKAKRpeYmf2Vvler/d0TOZUJpe3xdqvRFQdjJu8IGEKotb6pOeP
sd7Ribub1vfOaH2AYmolRfXgfn8az3xXyxNrOcN41XAe6IlBbKl2ZPNW1gQSrrk6
V6Ax0J/7FvySD6X4pm0Vet4eCmFs7S7+qkI+PBlQ5k7goDZsd7InvB2VbUcfRKws
WF3T6cOcenu02una7OXXm+MCo4dmnBh3CyOy37MoKxk9jkqWmye8xqfUf9yztveV
jxY1cVWdAnaqTjRvLTrP4cEqYfiEBJd3EFGfsFcczLg1P6JMlsVXGNtqGSk13FiP
qRMRfCmB+TxkRTEGRaibN6ACEBIg0hTRUiq5mmwqY5TkoHij0akXesRo3nhVTEiS
ZMtgqC6Drl4y6BtQ9qSr6OxWCtEMg6lnRqQxhfDBJr8G+e/TW466S91l/JFj5YnY
WoUbZbQKE3GSLFBSxgKZmdME/kMt0TfB4yMtdLCt0g0Ia3YVv2xtDF0mMPKA9jW6
Xw1x82TQznfTwkfoKiV92es7U1zzTQhJWI4nuSTUWjiLU+bLOoRnhZ2hSd35zC3W
4/Mp5jB0MO6IgoFH+Cv6DxOeUu1+4C6QeGfHinX6YVOQ1s9KOzV6O+3YMfLNeGay
aB1vCeQN5hXJsZy27/c2ZjNFH8erUiQsbz4btKSvUee2CEITQPtfk/0pP/BvyFl1
r3WFw5Goln42i57xzrlwmUuc88WM8O5+Iog4bhwQeXOJdTEDXj4+twt3WbD/ukq/
4akBnufO1COWvIR6xN+uhJsfMotF9OidIQc8NCftnI2h5gKTv/zupvDwc8l8wEBK
et0WcVcxjT7P7AqLXuooJ+vhoTi+PhIs8KNzTn4FuZbuW2o6QyMREPw/HssSG71Y
r4cDkVx3LH3g2N8TETAnud7BQSiQVvjzVOZld3NRg3+pF1XLQhDl6/qO/cnEI53I
empsBJVjdrK4hHYBFS8fpvlrzOib6v3OVul+5IjLY+txphL+vVWXFdEoU9zE8OD0
t3u/UacacOcrtZHzhOCBodZJO0nobSC2SgbSEPrP+WrxQ7SFwoF7gy/K4FcImOLk
oAyPKP2XPr7ps6qK24Lja8k1aXvSldhnxJ8HgQY52IqdvHaqku8LevkOdhQwDUCk
O7AQCAnco1qe2pfQUwHi+UT6twyyI1CBtywLjKo0SohTOwJrsaCNHdBk23GkEXXc
EeocU4nV3HabKLQ/667uoPEIzxk5DufPF2F3aw3fsGmyM9iApCfDhEIdO/ECRW8X
VB/jARuFr3QCtxkZifOyphzOrEC4shdgwGf6wOxfA16hGMJQ7z+vzezgIsI0lMXk
gyAqra9Wlh3HpdbfY3UgYPMIVEKiHWcc/Qiys8tUC6f3zELdG6jLWv9eljUTM7Oh
k5NnUk22rCDacOjg4OcAqjCIuLkYWz/wcVxHxqd1nwuern2Ogem9I1d3KRcf60/O
Vl4GI7ZkPTQQjDkJxb20LIu8f9CaojIozA6hXvVjcPqE0hUhvR2EsW9lldIPunfo
rpwx78UWhHeFM8my9o7f1/x60FUusqpGIpyBdnGI7Wi6Y/iIhKfke+DE7hLKYCDt
GTMgYunbZVALOVIJaQ1KCSWFJ12q6TFBbAnnyzxGua76lC6qlC3xJDCwtd791fAo
pdcbO6AiK36fZtdCBXX9Zc8Xe+qhBkaKVMcIVZGnXvcDVjcjPaBtpG3UDhWxxsP9
WjEAHH/7F3jDjmnBrG4nYzSbsIkCp7gyVLV5Z4VCKALzebbuHsFaQkWqif0xXZGH
I+WhEnNCuW75CD/UXW8Ul2vE5iMSN4veASEkQx3QnVdyC1hfuzp4YBR4fytFiydr
nV3osZvz30lSV+rqk8zKAXURy4kmNYrJmjwlfbr52YzoGHg4IJMPSsucEpf3N3ii
LhZFCvslQp/HQ8YwCZQ2IicKwsSvirtk4f0Tob0qAtNDQTXkl6LDgPaM4BWGbn0f
SL6uUDn1YOnfVbUUZYnvvQgSch4bA6rVKIkO6fiz3OTNi59S3uPUnuyeOJZRI571
9mmZ6OWaA06bzk8cuQ9cPs8Ah+j7SgwOYDYCKbH0zVQYr6Mhlrd5V3RaPkcGDgL0
Nxoq/X/p72Hc9Q0nwc7PEtD8LBi/zvzrWegn+ZJc58DYxf8Ma5xtY00u0D7b4syx
L5ZJyRaucLwM+sUsMylx1Xw/ZZksYmRRYMSLHO2NfG36/ikRggfCHauSYlEhCNuo
2SNFciGjRCiwIXSbUjW98bAESQnE1ZoasMMv7Jo5ZanvYajCc9dp6jWM59+RWQbY
P7e1Y2YE2gxx58g1yHRraHR47oPcYlbhr7L5kq9ncLbMlmIRvjjogz+jg5FMnz/V
ha/OcHLthBqkOGSo2YAF78kn5Q4tXZ2AU7TZI1h7rsiEfVt4aGaxv8+sVY5AHMIb
38hYnxiWa1uypCMfD6w3WJkrquJOnLNKLqe5rBjeaauQJryudF1RVPq9+24BstFe
rUF13oIaohyU/Bqq6GxviYhoWmcLUkWIM5Lr8j5/ak772gEcmmHGTbKOBXfQ6Qve
zxlhRuBWoGfj5uVViET/CWWn0b3lwk7dk/v919h645JtC/2x3RzbArvqG6gjP9Vh
72SdZUa5b9ldCAoEvFYzMrsud6Qt1L/vwnS1FcbdE/ieVSjmxH75tn1NIuh7d0Wr
nVl2muEW+FnoaDL3zrYYhdyu5TQJuZwhoVvvZe8vT8JQoV+N/q45QOQfigmfSVHM
BV69iAJ5E5LhZbtDKTET9vQ/xrONChpJMCxzgC8aRNAy3KeKqoNLhGqhQ2WbLGJL
cXMjsuKJIwNxFaq3CcgWVV1rpa9fsZMk9s+p6gsEkrxMUsd+pFukiqJFbDcpmYv/
4QN7Gv+bSOUd50Vom+9XsYKSx2Bc1hV66NdaTNfF61Sr+WqmdzmY+KaxwutpBWHl
Vg+dsBCQPqOgjxltzGVKkPdijeqvKlHlNAcePVg4tG9wiyC/tJyMTqewV41BxZh0
QlboqaVB65tRkKqMaI6HfdeqTVUWJE4ViI4rokgzuhGQhvAvLCsKZG9fFRH7myAC
Rl36RduyBe1fpMFt6TBMmT6Uo5EOoUGXvAgwx8cJmloiXTQSCh6xolccQSf5OlGJ
nMKxUJf9Ng3seWQYxzqOwDIcTJDYkY4kJeubT/oXf5EmFO2Eb5jJdfj8642gd3jI
bCaGAV28JlK4CPVvrvnW48+rbqBQ868+QfJuBdifX42YSj0YBTD3fWQs2dtz+ZSl
a4wzVDVfEFYxHrD3yfH+H5fFacdx/G4rb6woNX9M/WZfFMzu49eCSM8dIJDNOe52
TY1DY63QHJ77MzhU7UAPuiA6LeechqGzsRP0eQdhODbrAvpMgZ+SA5WKqtSlf+9n
q3/ykqQUuIv+wKNuy8G1X9rUyhIf+x/Ux0MFtN7KT0kgpuqwSAxvdKIbxQWWsgS+
5xM/YjSjc/4ohABvbP4M0KjpVjX9j24dYfujq0DN01qzgXqINejK88TysQoXusW8
Jh/cPXJEsziU0+SEDtlA02AEH4A4KgIRlm9jhY3ujWa+oxuyTGix2w1+PCUgugf7
6AiuuEErpZw26PUSXpscU1ucVSwdQn27VIZXjIUmjQIQs8rBKLidkIfps0ReUHI3
gAA1Fc8g8ZyXKLIzQKG9FMooEE3KmJL1J8ARiU/2f8s/LyAlN7XOrdvJ++INx305
ZxRr5+x5zGYgJdXCApMZ1jqD3JgcU0ZAwzNjNHnXeQ9PN1SIJ4Fs5UMvegx/C1mb
Irv8KjUW9RPS9mawQz1A4TyX1v+Za+tfGR1IlBQACby43mf2Uc7EMaK6Fhf5EXYq
VZSx9+Ckq1QZSXworO60DZdDKmgeWU8KGc5X5S6+yed2fLypeO4v7OJuJuA9NBp5
B0xpTqNi0o/iO0x/Vpf6BxbFNeBVKhu//LpKD2gHqFlOyd02Uy4IGvyCdqUSJwHS
X+FOK4Rdg8cJjfugOMyiCe2H1bZuGTAAeg9BBUbJTg0gVWaYa9xUEnBN9MTpsMJ7
3PrqtvzC93auT9clFirFSQoSumhhjsS6vbmtzFBHQB2nUUnoI5hnNYoUtqlr1SKH
3n0z7QNePbyNyKNMaTt/tXpfVUX04US6v+DDFxl+A1P0zPngAPn9NB9iHwheNP+e
CQxjWmqbGCCl5J1heXBCjUimGVE0yyG/YT76t0533CbiuVNGEP/XqNBBL1kNlU3z
jrvPFWG0tihtwH+kBA5B93qSLnm7O1xXkEljohVbUfVdPt3Gmdn4qKd1Kkem9yD4
Zew041RVcZK5ALy0nX6ZC6wnYH6F39bPu0s3YKpqtwseonOd3ihzxvTP5Cy7FjG4
vh9oapUmLfAbA/cKCnjuDs3O7xFvOXt77ITjryjZcwo33nSHLctYPmcY4EEpip8x
WueXIlKwtUuLV7TnInjNUWGMvppFLILEHtt6nuvniRTplfspC91PtSa+gY2tlUO0
pq/eE2ECmtj2I2N+cwWoG+IyHYC8V6S/3Ig1EnKLFvzbJrTswVk9LiT0Qx1Hkw54
MRDxY7/l6hSCxhN/TY5mjI1CLm+Tk2sZ6qzbbxnZ+PF6/CONFVOgsAG9ogRDS7aB
xbL1JtzcTqOjWlsQYwuhpnIQopnUNWrwYWJs9TyXPW7r+SagOQcyDiRCiM7IEupd
ayBAy43i3wpu5/SQMzKwhpD2GseBxW5PaSzrYjQe3aeTdwETs47r+F1gZafj3c9n
4vFU7GwWZWLWvZbxOGMsoTjOcNH10tURGibbEFIAu5KvljtSUP2LO06vr9YDTIsb
GlrybOpJULZgucVTqW+dFbRQH+ozyvdpwCAEFF6dq3EKigdXHgiJtVhfs4NVxgBj
OaJbe2B7gJHV4rhRQ0heHBajYEKyg9ncSWTrVdJhxpyProCUhCA6MHnD9G4vx34R
LADVtOSepOOgsa7JThtLHZN3h+m6qqvl463ZEIDKRozCLAhUc5np1pee5W0v+c5P
89gxEcJZSqy2huFu/PH1EWA9k9QDl7/huJiPJybQAP2+Dulg/ughG5NnOjNh63C0
3vpRdLW99WVBvKIK4bxIeqedGnOHxZmJBTxkUYysXPtKrh+t/KGbnVxdLp8F+l1H
W95TMNAcgQPcm8R6C/tzPU9bNziLut1HFXUx6hockJldceXx/cFM/WPg0I5pb8Qs
FwT/ur6xnFDW05/jfftzL8/fXZIyr4w7Z7kSiS11G5EPrb3QLmfywd1OvbuupkyQ
wNyK1LbZH82T0qqRvRPKEelL8y2/TPp1rBEFpkgVIgTPoLGhcktZMYChJVym9sYL
2vDrWgvuVG6NrDJENeU+n643SpwkkSmthaRUBiajtecau/EUquB4RGPn5wu/p0YZ
WzumwzhIhot6BIsAt2FmHlds2c717q9MAi0KIWs1MdWwL8Nqxj1jgEv14F80CPB9
+R2hN7Bq3503mypVFZcAgeUvuqgno0IYW0hgB/sKjpCATFlwDtYlQBucPdxGjT6q
dXGgbWNrHZ76QkGScg9jz1IsDeBSQU5g/h7UnM5vT7BuKd3CxIK1PioI73OySj22
vPh1pg+/PpUjQLs5xghtQYiWxEvHXv9f006UwfIhtoXklKTIh2y7PBH1T6Wirl+B
UOQABc4425YCW+YMPRiyzWPdaJI1PH94A8IMwnJELUbF8XzCegQewnpKCpLKSEdF
hUMe/PnPA3tp3El/l01kdVG4EAKWqhqmSHLmS3YX/S2NIaET0hqYYXJND3e6AMz2
XxNHx8xlixewtXt40QNqjRF1XPKnX6B0zGQ/texGGDU5Rr2QiQBe3NuI/BHbDv2F
YxT0Dd7RHT3TsyCz3X/1g1ThKBxCbVn5yV+lt3U1XZfo6zgrmCRdIOrC4kYFt0+9
XvZ/kjQkwL/LqGkjM25V/nbG3HQ8Mj65+lhOUztHXlvfDp2pfFslQ6X0nJC0OjM8
O7ndnMKJmn3/WJlSMVbBCvmfbp+QpBcbLUNRKOgT401oSwLFcBSFJou3lCsEW6Db
mQrAa/Qc0+SOBYDGmMq8AcpCUJc13+H7kn+kz9z/O5PoJHgVjlGc4KXmj/FQ1+9j
jt/WDZZInXTcYgO5LaIf6tNF9YwDbozDBp91hSv6tUYpqcF6IeDggVvTKY7fx3/W
lJGAf+69fOhieaGSTJ0alIwujUKZR3x3ieY5kbLfri1sFKoZDIkKtYCa+LXu4ZqI
MlMK5R6ZRlbqs9wovt5TyJQLc1c3dADX+J+lyLEK//5xqPCowzBHjV6cURhy6ECE
Xugvk+ajYI/b0InSOw0aIda/nh/+oOmFS77vp3pZJ4TNoxXIvlzCrp4dvdZC5RK/
dKIhwB+g9dCrljK3f8hf47UaGNXzVsER2iBPDjdwclVwFYzPQs3ekuuCGZieaj2P
FpSdrh5fxrKl7S+iZm2LhcZCQX5tKIy7I62LHSqxsrSx2gFWLnx4yFQ46fH5UAdN
9oBZfuI9PLSbVcP86kemwQ2Nw2yLpNcFC9YGxXq2bDhGonXwHgFEoWJkK75wsRO7
KaZm1igCRj1dl7nY2C8p/CkL65eK9AD3ZsLKzpeuwohVNXySuEGHn0z0JjJxyxCQ
cyvyj5ACJJ+xm9kTRpvZc5VRcdMcFArqVE3hLdmJ5AA3EF6R3tJ3H/kj9zOOl6g9
jxlRgGk1viB2R2AsDqaXos2WSEA1DZNdb3dtTg/70bYx2irhtZeRaHXsdDRjnPBp
Z8NgfCRPzj6TJgr/9jb5UacDc78CyU/3TnhRSfjyLKS7TYcE2/RZaSuMp0rPKNBy
0p2Ca3tgTVGAMd1MSu1iKpyWDq2rqibRN1GtZD5UdGzKP/OkaHfjPZ74RYZ07cDD
c6VldknfWsNm1tJlUHG84uFLa9P07sSkdhG2QEjxe7Ikftn/oEuo8KjKNcjOClZ1
zX2ecmM97OfrZSy+zF7mo8rvIyJXCLvSZn/eBy8JqO8UNHO1otgmLxcZ4bT2Lu7+
IOO9ZQUm6sdBK45RKQ7sH+br3Vr8sa/TnKndgsG92q1+2cWSSruoaofFIE6r/sxB
VIeBQykjRYEDajG8HZrv1JB7K3qUDCyJUSuzDxehxBkJuoK81Ckvw5pz061gcOlw
eriA/Zp1/qi88LFQ8NrC5I/zVGm0p8tsiRYZFtyBU1sZ1A+lNKczdZAsOJO7ctwx
LtUXceZFeTgl4jr5ZVrB4BzIU966/PXrb6KkdEDNWdKW06V58tFRQxwIqTU41bsj
H3bv0k96bsA7KNLh72JUUuJFbDgEf+isBGeW6nKB23CWc+Qk9TD6+Y2eRUDUPsH2
hK1JfTmEZYhSUhcaNYqQYLoQr6rAY2Pldm7ECgQDB4p9bsTgTn1S3MwK9e/JSOtR
4Z+V8Az8EZkCjhmDCxWDfiALliifqzPxJ08t38taclRbKtmZ6Jr2jcfJ+0utrXM6
xe5lF5ZDFGloJ1JC4xrG9iOo+zzYyIZ6x1RMpD3GoxnkkGRLNsnQaAzgrsJe+lAS
Y7VWYW2DWYv7j0BwXC/mFtBORbnIJRKdqkYQ0Gu9yFnSAoQR3ciDNxtZ3t9u80j6
8EN//BIVG+Jf7ayn+LGlmxZdnv2SlpvGfaqdDUhG60mNatiKkuhNiOpXEFJV/Af0
0awZzcx04Ix+si1vHFRzTjp6En4xXdMfelqpBcxsavpkGjVGf3qM5yDWqOwlhcr4
VZCIG/5xP51tQNUxDMj8LhSbX69ChzLZkS46u1eS4rgdGXPBSyDGxXiRPtFWWuun
70E6lDdr6xtGyxWfMiqFJEmvqt027XD2SrHAsoMYVxX8/InRx4vMWL4AgUVVEwZV
8mmNdMgQ8zDQG9+dBBp4LcPq++NQF9V+QjUhL57t+BjFANItHL0FYx2Yha6e1n0B
EbQn0Ws14/W7qSOsgbrWM/xp8yDrS3uHM0gFG0Vafh3fQOI/o/EZoc7DPBYe6daP
9XX6Cibq1hqaHB/fQ6Eat17cYQrGGAv4pCX24BLAwzEX0zVR4K9rx8zVVcG95c6t
sNP31AsH0DHAo+Bo6p+eJI+A5vzPLWZlcn6fgKM+QDnCOTZysX6aelM24XRv5rBC
tQO4SdSQUrxrpqMyj2RUXv3gwz6RgAa5SKx/WZYjUhU4YGepN6qh4F4tQDIQnwTU
NfxxMhSMSpHMM+XCFiEyKuApJ1u2hENcNn24OBIB2MghvK1rCjg7dLmRwfHaYiJq
jvSvq+iI0uhrz9bdiffKcgsu1MyBG7vl7tn09LcQyZH8sa+s0fA8P8GeNyt8E9Hp
3jsOF5VsJnEv3a6VtRzmi54UThIAy70weDni4eSVRDW+gwbMWPMVWlPme31Hk/kW
i3mLdj/Gg0XNt8sCbMreQaP/pPUjTJpUWlLwqYAV5KjcL0vS7Vhu5DLjG/wKuE0U
NzCyUHqbSC053miKLsvbaeCK7y02DnBItGuAd8EMV9O9e9C2uADrfd7VQs0cvKuc
Y+yYVFtfWZuZJOBMsFGXdxi8mUi/ua5kPhQSc27sh0Dd+yPcfTd7kRBV90z5B5YS
tMkmML4cI2uQfSEncWExHrFzEWGH1piDnOkc7u5jB4o6gSSYp5I16638FhKZ0Y0f
FLHH/IBvs7Hi0WpktLoC3TWIU9pwTOZYfDYB58HNOyxjBDomnQg+ytYf/lyW4W9N
xWZSBAPOz7c107oEJ++38mFBabgoKcX32jjyuS/31n3U583bhx1OlEvRs37jB2Jy
r37dREz7b2nHeYLoXMTWaMXUdslZy4pT2G95DzseT4wMbT16wp14jNMus4l+be7t
IMwCuZOZ64JjFyqD3iB0qizDXiK6AUsksusmd6BOoa+7uT662sX0TMeEpYzJv50F
SpGkbc39mYEQlWNpvnV3VQ4rU73mvE+ybDdgFjhsoPQYa9OeTwH0/1SMOR8GKCVI
+DXZlj+lwUXhcleSBGfisq1QflemZs/hwmmgxYrT/VCi9ZncqA2Wd6eqXH0U4FGi
SdJTJzJU3skxm89eQ4/4mAt/q7ybKigUhwnoOrgnv0H1tikoUEK5jgnXGGiItoeV
MLZenjiPaS+GgTdFLFRZv7mFWYCqKysQHyWhFK7E686/+72ZVJxdD21SKlru43r1
Q2VzGopMTuVld4wiDo1/BSLfzJouNTy4g1xxDO/AcJoPcGMnj7CYQS8m7yl9j8sA
xb4K5fD94nS8SZ6YbpyJYpyA/s/GQzWBg8/Lclb2o1a8FRcb5viWxteTtjVe+rNS
J7HW9f0u6gk8AQd356DzI7gSs/1HSaGllFto1v4EiE9BZzsnPpnuQjneeKzXOAEe
FlzWph7CUgg38DH3QKqk69ArXHt8EZQHFyyN0ZKQylsl83L/A5aIxIzPfZpkFtet
pwHLiczXFG0pFxgttAonAREtHSptR5nwiF0d14UR78eTwT/SMwgzpGbUtjC1QjNT
YOhASgJZe779x0M/CDAuNeKeXjrDinWrLJG4zPvtM0LwUhr8nEoYjwE4duIF1KNS
TRwzkih+PJVcpWcilIKzrExOJg0q+DVdNyZ3tKIbZKy3lPGCWmmT/CS/Nk3ekALM
NVzUQFX+fZxRAEnFkIhkJBi7O/aKTaUCWnBsFyXnHZjelkt0WpRwysWEgwAjsBXE
X2kZYh9+wqncQoB82G0mZWCoKEd4+Y8jpqjwHLzaRkCgC2XIKzdVVKMYIORqOpOp
zf56CyOVt4hex2/SeiG7yg4xkzDoGQSrJIk02TL5cttF+7Z2MowYry2tU1nQjnFn
uC3d/HbNJjQ0zWA3oMinDB1PlyS8460OUdAVwNPIXo4V7v2pCy7nzq/RuAZPfdPE
qXTsDTy8DQ0gujuPZTzv9Z+DQBD+L2iSd29ERMh4w/XDPDMphRAhHx2tbUfgXibH
9aNTqO6Skciy5qya/HJxbK8ilsSX77qsGvJgRX6e4xYIM2t2mA4x7LsA058e9DJq
VlWUXGlupReUq5jQL3hR0QdV22dEpeBav8pFae3A7h3DWmZ6Xt20GtUcXxXJ87W1
jjSUcYL9EXQqOTUneZ/L0oKP824DQsxsTlWb/tlM+l0+fVjyVbVCcMYcNtRUx+ha
/szZ7nE3byqVb+OUeRdJWAkSX2rI21RkMezJEKgp+saGG7KkmB+FzHqCtI1JJMyY
lrQ8dx3v1iA/pJiwPxDN/s7DCwuJk6C5h1ceMAzc8oWXplKfTKZPzXnacf6NHXmd
NapGpcvWUFgQGZFZ2XDES1Mle/ydu7nK9nU40ZMfBkqUycIm7tJFzIvZsJ4HN9fA
OomkO+11hE5lGEMly67NAAeIiocj4kskzCEtb2FpJlcOCpzKlj9N9IRw4VJSghzC
qsKEIcNvVB9jf3QG8DHGOHA/55wYPlYY1PaTgNYEhiHxql5z4aI4VRTWM1ec2jDR
DkDTEOPXOzg/P2SeNH1T/w9GWFSnTNsS5Ok64mmOvF1t+JVVleS4I05Kd1mKr0AB
duToZduSTYWiTXYvZVREnZXhcij9uqgoEK7MowSyZ8YJTO2wh76Q7VfOUQQdEMFP
jUHWwi04A0SLXv7SaJlNrNEjHsU8CeDlHhA1CmXNO1TT6Qo/PoQj7XREmbcRNGuq
6JiPtj8nvcPKJRwzHHyZidcO+4aaRMG3Peb/pye4R/sTagOMmRx6GyGZAbfv/9Vw
zAW/ZFimj+hMZkiQ9U3cuOy1eIpCKyiOKlNJa/pMqVEiCTab6Iz9KoPA0HltTYFv
YCM9o2s+RGyRqcltDbODku6qi8iplPIOgbYII5SsE7xCp1jGRi4mohbp2NXUjePK
yahYeWpTerLR51/9LtHmh+hPGrbUL2sxt0O4Vb0+EZ9SzF5XzZK55XFRAPW9pUN/
dDcquS1KI5V07WyeBB/eGADderWabO2pCMiXHU7SuD8LV/ckdN47BRcTUicbPxb1
WOrn/vrekMj+rbyqJUSwgher4yVYP6xnWDLrEAoZE0paT9JJothNY8C0jqL/yPe6
QkPETTnizr693mDqmYlMrG7LqJa2hznu7u7ksgSpkDQg64Sfbp7cHE0WcClJMwwr
C6gITIJjs98REjVz19vQgdDGC8R9Eh6DtfnSMczSpqTWaN7D+1TQu8eQ6Nvo3bG8
WsApT2hvJEuApoLnY6mMzjO4qt0kdVHgcHvPBR/amt28Dc8qiy3qAulxw9NesSrC
AuVCXmulZYMJCVikkDYkJ23u7kVIlBEvlgslr2GGZ6qcZzIE7J0LkB3HM38kNIfp
Ydijb84eQKejxtw3600ObB+KD9PkyEtBijB+NkkJp//LbLdqwCIwIaEBdlCjmgI6
J+j/4Hu/UALldQaUsGJ4h/il19aSn/EPLe5p4p+7yEFKwKIKPjUy+V8NTgByIuvw
n3jl8fMGiSDEXVLXoXUPP1Yc7da6nU3lG2pz6ULbKsLE7/hKYfySwwuOQRlJgVqF
peahP9AgyIsbqPCF8q96Rvf0Ucx1QcNKNACMRQ2q6lbowxb2FuFEbUhPFALHhTuK
TPSV/ZNCTAletjmvqAIZGjLFa8uiazqgrSL3bOrtvMgaG/+yTPbJURuzsDqu8+ye
cwoCrf8Budn26086YWNoJ7MrDgrXl063KcN1et00kbcOjvfo9uSIfM+Q1zxGjEU6
pTKY5NLzObHWaa+DJdC7j0wqBoEklHJZKPMMD5g3/gT2sAe1id2oxK5WivhAvaC5
TrxLoSV7TtrnYNaBV9zUp4o1KwJpNplH1XQQ3dA3/2NcAmOgR5vHEF83bYPK4xcA
l1g/S/AzL4Uown1EtoFZS/68hNTVi/iw5nC1ve8+S2a8r5c+J8DRIRWNz1oJgyjD
kDnrN3wOI/whdphdzl0RLwLB8TtmWR3vYZ7lRxdSiq3Miub+LF4GImMt+MjXS3TA
ug+id9270amQxx9WMpquL+D9mpMP9vwSDlEsHuolxHATQd/Uh/Y5xXmz+5cegQtK
+uKlEpmz2HyQSup+5dbN6CJCj6xeHQxS60KVvxBSrP1/YoaGr8sjkbkFvUYLfyRx
vG7y4IhXKIoK9vg7tnNesMytBRnUFu3IjTGs1i3Qqydcgy/4I3eaBRF9BJFnMgWG
2pQZb6zD10SFG8h+cJgE7byS42CPJcTtGOUoXjTPD2WvLKo447Tbm1XTua+3G0Nb
2se5e7HCIU0WfxnLnaqDzkL+dcNHqAZZmHBAFK/7ZwxnVdRi+rt8wSkjnjWH4a9L
Nj+lciJMGDaRbwrlhb6NTukF4NRX7VK4UMNfwGYz47RlRjOJNdJ2shrscnBRX/Ym
aI3Lz6GxvRK3S2bpsdEt7Y/PW2BT8rdcYgHphJCRf4OJSESzC/Xze+IWMUE98mtw
U9um0+GFs7nvPQrymUT5i064WH0+GzcKxGzIv9XEQTb00sYls+loDz67iEQZzfHJ
UhutvwJMDwquU4qdGU22QrDOMWUcc4VbNO37umG4vDhhpDcVmQXM2z6nCUpWp3kQ
jHSCwXSFVXbRcOllhak+edNHC1LhaNbW3cOHxD51+LnzY6ixHbo2v9dx+GEHNY2F
YE0CXfj6vvpbdDPWaKVjH/JpDKIoXYVhH6ug7xg/5zmkQd7NHjaphvTcWQbJuXiG
+Fo6mPvIYnUfyW+Aa0LFvfUrBUM//9eLOIYLwjWaitAij8PGg+Zis9lraGmE5W2c
uUXHtwhZVIC4VfCH0Vh2VIlvAG1wHhcRa18nlR7jX+eDor8OkI85U/Q5iqt0P8m3
IcotQJ8cPwhJ6t213Usp+Hi/yJ6Uv54hXp41Gw6W0tLvuNsaidA1iP7rmbq0R5an
3v9z7bDFk9A5q+gcp1ccdvY/bU45/CGPBrjN4Huhsv+tcBqRvPqMUTwTZnDuQJlZ
jp8wWK65vUxSUwwCPthyq+4x7UZ8ow2M6F12qRFFmdftpjQMBZ+JHD2fvwHwJ7AE
QjaBzjuo/J818RkxUg9dpjtbduY08Q9YiEZytDXP8rnGTFQT4WJVuD0To70bpwIx
DcMtqk7A7cTByRGnUUWR0HieYmDt+rKPsXDviQnOjvzN5nusWstXNjetYpaFOVtH
+imcOOh8q/csdI2sqgL66yd6b8WQ+jlknqhYtkwcdxbW4Zt+KPJ8iDcfYgG3Z6Vf
uiKwlUmpy9VkDzXIjH3LU1WfOiSEEnH7CWjpnUq5pOCwDv0EH7agB9ftRI5xPicd
+fd5qCDG9tOQ6L7/KKjwJ1nGQdo0d1WhfOh57UNCULVvd8PzorBO5NC2H6U+BHbP
J4Ag2HIOBpoeR7H3C14oxBMafIWSl64Fh0a4WGVRzenpVo9TP8top2RBFaoNzMfU
H/YgixTw76KZL0c99N3CiPnOK94Pd09S8UEtOP1tKemJAQc1CxeFiiGzH27kGhZs
eOa3zKVfuSbSvf9c8526QyaIXxrfXGVETSEOUXs5HD4Ua3JEQ4SWtnzC94852zE0
y/IJFQ5AVWZfWSgp0rF6EWGUBv2DyiKJabAt6N0A31qOWCceHkljkChjVnJ1NB8T
HMPL2+wNqyCgG6Yplzn/Wn/Lj+qAG4m/6mNfMSCiZAZbvn6NhnIpgatWa0J0DZMA
bPzI3/REAr8iQXxtx/OjQZNdmJ2lnsktV/PynSVCGQ8JtP3AqMcFR74nkJXFWQ5D
ZHlld5mEFURNIaQxaFFRDn+hb+w9gY0CZhhq3F3XhzAeNk90cq+wPH8dgCooU5Az
5EswiiyJiw7eAlWe/JmUQ8uxSebvsLryW16yntPqbQoulGjHTQoNbQL6Ywo396sM
5p4ddpxKXCJQUUJm78q4u216LeeTUW35b5ZQxFr369VUCMglVhjfmnBtXZzEpSOa
aGkKwXx1wttOXqGJBRtrcpQKzkZ3BvN67RitPL3uaHTAfMQ7MqcmXy1pyFN8778J
8k/u4B1PHuHZugNAObywgNxQWSULH3vxj1iG6DVFrR+AnyhKo2Xr/nT2cpwKxAxJ
90ndOrtt0BGusmyXcIEw6BP+UM7UL799vfWZAYmpNQRKZnAdIM/BpLVZJjLcCMAe
skoiImRoTkZrpx6PuBf7YAkLjRqyGi6H492P8/BSTLz8JWv+tMEPTbi+T+gQykF0
aheoE9F+aWMalsRYOYP3eVjzIanzj/9k1aPk7AB5x1bbE1FlyhqOgjML/gx5Qpjw
RiL1jSBzE1eqWwrMTokeULZXRIfjQSjQb1p9kc9Q6Cmme042Kh0WlPWYFPXMoRiP
yQSAVJ5akEIhoBPTatbwjzvpLPVjPzDfDBJWPIENsBl3Y/Y3VZpX89g3q0zYOQV0
InoY54b7c4p8n9Re7SWXotx3h77yhIIMI0jAVp/eXr+dADtoy04hd/MDJm+X6udF
jTMhPWNFpcmM3EoXQPP5Uq+eSwNqInkm6X+TMVOqh97dHoX0kCgsDA6eOOJo/IKh
MTxm1PTrCdnQA6MrwhBfKWXA9w8mUYaknlWzOPp4NR69T49bDhF3KeFBGmEQK7SU
cl2ezZB+us4AD985IYhNFOSKsKBe0pozDVLSckcB8KQkXR537eV8OtT1VIEJENky
Yot5ltaQ6lIZt3wkIZ+kDn6SHqiZ9k4nubYfifdBMLxxyPsk7/tWco71NE0g/jKM
u7GBKyCZpPow7J9Uuav1GCrW2hDzYg5TCPKb3TK33OpZ+JY7c0/BZny/erXu+sYQ
aKLgWV/lV9z7IfAltIrShy0CFhXJiVO5InxtE0P/czD9eQqofik7RgbILz0Yo+fB
TVkchSXcFddB2AEADcyDUntFpbNHOyH5OYWfQGRQ+DOUy6DzBsKB5OGHpjpvj3c0
fEO2qkKCb0bk/OGhe20BCtn6rLt3gsJmba6HFO4mUBL7ILc+gBXToTwNsNAJkKCV
PrRd2nQ7kcJiyERSjod5q3VGEkBs0qDsx4OeECXUgqWH1RWWJgSbVfduUg6rgEP6
TAaYJf15jxbWlGjzZyEBTU83/Ngj9CBB/LO6VtILnPR7QkJ0pHAH3RIxmRRK1dLm
xGxksQkh0jmjeW+EPDedypIiHzulzR/zK4RwUtGEBrJNza3t6VBKAp0pXt/t+tnm
B2gMFwWwh/lYPTBwL49pAPuCpZW6Zl+m9040LTv6WiGg+OL9AEk/t5nz2DmINhSF
rQWJBqaroPFLPPQReQ9A+2PGPism6ZfpJq0AhhibV0RHiAaeaUDQEc3IGy6UXR+9
8L43efkPT0aqVcp0lnlH06GKSWighv7L7bWrOcXhOASiNa/tL3dAk7EGcWgCuRWm
Zq4c7HbxrGq0QDMzqWCgftGcSDJFgElF0HBxXEhXW4q2pl1HsmdZi8/FfGqz3aq9
QZ1fGWAEU5kNGdsNacH0aV0RGad8MjK/7yh74jFylRqVIblON9SeDcXqLVMbQK0a
JsLPKLgrX2mLZW9pTil67Wje5NPfp80EHj+Pi/EGDHU8rkamBIs68kGYvVOS+j/c
XtGsA3eemO7C1Mxo0fsrnLhHWN9rA5E1R+52oGRB0ShWStt0ucveBH+r3Jf0mT4g
P+oY1LxgOZDQpwG7cz/WWsCylPgvw5t+eTF4m65BMetqdwObQzvlRyxW8/Pk8CYP
2ESXIoPYDU5MdKkCAkvQEaS7UPiL+GtooF5F854cr+KnQDl4NR52LAaYA5iS0Teb
lAt+C3is0ChsvuQ+0jCmNCTgWpN1NOnsLksQsiavcZXV/YROzhXaRWcqEEcrIcL2
atpYVOyPQGzF0at4qEgq2vnGLabyg7XkxO4RJOuoHaiczoAmDDP65A46HTM3P8a7
YiUmetdajwha5BEoRkRbtxEAmcUmeV1cV6Gd7p2pNBzUvkAVk9nxrp4TrIiGIGm2
7l41J5Na/POe1yyjAwYIXB0RkxMbNn4HHcRNxmdyuFMHNbdsUqHNPu5R/A2Oryxx
zjBq/Rzy+MYLY7voT9Gc9yb4G3B2AKJHxf/BPaOUdfXiCslvN9qdXOVyJrz93cxB
P6F2xYKq6K2Bl43OYpxt0RSfxpJZpUZAwZeDn0mCIx1CrfJzgphZh7xS0PMWIpjM
Fc6AtVgv3OPUKuNyZR0I7PUXVThn0wjX9uuAE87xfUS3+LEwQC2hy4BRUvY7tQq1
DPSZOU8klW0WUjcYA/ltHQeI+DagiiWQVY8Oc4hswysXnEx7Su/b5Mb6JgLDqDDj
UHc6W5imBEc2L4yzQXcKli6Hw4NuWI69eFzgc2bEF85EM5FkRe4cr8rH3s1ZLgb1
MoZ5BLE0IZMOZo+XDgE5t8pr3n7M4MFXtDn4NJ2NJ0RBh/8zdrZcT1/PvLqYnsV9
4X2VCbsQjbGw0AqBYiqNbCXJyQ/5iBV1bLTgfNgOozTzJwLd81Eu/guD6XLxGgA3
Mht/x3AupNf5dyFZr3dS+R2c48lMMXM31fWikiwNqWoisPxjeD0X7lWoWSex8ume
6OBYDtY7QUxdnuRSLSDj1RHigb6sNSDZKmAHSIfAe6A5GfTnCeeoSlcJm49LFiTj
CxjdvfLK9E+8vWgUOmwqWw4cMdM3z1F4LsLQlbo9imw0LLod32JtbqqUAdHZYG7Z
XW7J0bDG71WOZOJxt/vbi/nMauI0q2PSBNCdsCaWYN2gcJSs83PyNomJjD2gbMkn
pH8UjvwnYmQmihH5xMdpBywA2+GZKRuZE0x53Wpw4G/cFP0Ar1H3ZCh7ZRrKvlfm
KDIFfM/IYvJGANV0L7EAqS/p1cNcnhslgOpv8OFZPaXL+2G/NIwOyKyF155eO7XA
9B0tiwcMtn3pSmmLJwnxzBhIXLDlya9U9zobHyMvSzqK4e1+6mDuh0o3jU7HYurQ
kDcHh/iQ3F0O9dIwGWu/WikokWvPER9Vevybm59Oj56jr/45mG4SgV4s9ehch9DX
oTmHs6rH+dYusVikai1rwAkjxRL5Gdv1mmClHzt2U1acoFDnKJUPiSz0mG/Z4dHj
pJJrNiF2uOfYpa9sczgZzQwIvd01y2PnU2pZkiwLtGtEQXDFx49pmVBeFnW7W0qN
7bFH9ZctLJfLUwZkQ+siO5EW1bx+RFXdXTi5HlgEHdcz6+U7Kyu5QFwW0f8LZo2V
UBkDIgoJTOipAWyaGCk9ylN6eY0/fvxtk3bVEdR/VFIe783D8/H1fm8k2gJh1SCr
17ZfRwDnrlUZTwOwVtOXTKSbvAmlJ1W7o2Ta/iHZNee3sJXMdUincK4oT0AzXBHt
sQiOdXi+jhJPyCSzkozJFF/HYbrCAWPfNbuWbU8g2pgeWLw3eUBXZa7cDHpSWDeL
zZt+f+DiVE/bh43lXOBRLMuPp+GBM2fb7v7a049s3ag6NC12mNybtytAF5J8Jzxk
bSGS6hqhvcTxBSUFE2JynbEV8UCmkP8aTy3sLyif1fCfVMzVumX/hspZW/zJZCKi
45uvWlePTK0sKuhp8/jZ2MqApExwe/LK5o+SVsgPpF5H/pjfnzwsWju0Dm0bWCnf
T7Aty8FDlZ8iUQ9/7aUxLqyqbQaoPQ0YL8vJUOaVnlm2KlLNguyA5704yHuOEj+H
QAh7W94uN6GC9e6QGk3Dk2L5c9hfSVCGZKIyBx4mnsYsSg9i+UVneCpUkdhKVDbf
XSgq49eY4sgeUoQ7oKbbrCO2YEZn5TXuwAO6J5nPVU6MwBIegsk62OiF69aSMFGd
WoLke8rc8W7mAblmiiEZ4osWEfasdBYnVJ8mfmW9berEGds4O8XbvHY2azIGYSSN
rHbv17qMf71/R3SDIoqlBUdQ4OQu8GJ7FmAMitdDA2BTADiGGOGRp9i8HX/zbCXp
AtLTFRsVKH0+Hot9TdOhYZemXADGG+3LaqpMuWACxPS4tsZR37EZ8JA5n8Lf7Uut
cgZPq+qm4+UQvy7A7bIsZeyDmEOepGvS7/YbvAniExwxEQpbvUck29taB3gKOnzc
ajyfqos5bJRVR4uA6nfmKIl1YfpH0lFR1LflTO5Oo1Z6ddyCSJRcjAx64F4ZJyHD
ub7I3DJ+4oE3F0N2MtMAN+nhehqaDhzIoN9CZuaXOSmRAjb/esXWzihvrdMrA3Pt
OCuHgdu2NNfWDzNQJlLbu5eYnr87ErxDhanP2C2aGlf+4V6BGVuLYL5sjJi5m98+
a7hK+Yh88tsr+PeAiCE5bn2Lp3xSi7BLD5M+GaipgbmxMWSFQ1Nzlk/WUb3IO+4m
gERG72Ha9KDGlc26P4JlySlk67/pc8mi/+T5tBymz0a6q6q1mNikg6haXiXsyPTW
aNYcqP36RuCuqawXVzM1sBW7z0IJgDqbBff6cn4CbwZPJLV+7y78Nh0rlKSEgtqD
NpN+1qVA5ibMg52+tAPZqUAPNbhLq9vBCgeQ+xE11pOQEaXCCAJQKMCI4p0Da0we
X9ILReIQ6+5Vj05/wL4iEfffNIngXnDEAjGlOB+EJyDunnH+zjIg9y4kM5DCQz7S
jD7MfNeZImUmYFOMfSV9oRUbluHYkUs/Fe1QA/l29CGfad0vw3LYNglYowOtHTmF
0VFpKLj+WCfW53Vv7F5gC5PK1qJhO30ohwhBvQLTPgT4Rr8Dyns3+ySSj6Vh9073
DzeUl9LjRDpj5Hjo1xOctwDGOZ9N8Tj2Rw8i0wsm7nlHZCWYohOik9bQpXVlUju2
8nE58woeR93XlZQd/kPvqykPaqDssXlsUMU2sa3uPI1QHueFlCyNjk8x1LZL/MEv
ORlarWl/aTyj9X5YbBqzkslwcEDotMUm4b+58Bbvm7ZYCZMoXUXCIeKKEGnqqWFN
e3GBDlH09KfUCZSxfboOXxkXOgjPZr7CYi1onRFjjVBDHrF8FoZbn/gKQr62nnsP
la9IRmOcxto8zPIUyqTqLg4hkKXUwLhl/k2onzp2I0ZfwbveNzxJi5EOPaGUD9NN
sy620/8dipGf+gjspV+8Ft91amGofyFXuT9sD5KU7iDrIAYj62WhwwD0jxIdwJ/0
t7RXrCmb2hzJgosgtUc+qp9EILsCLLJzBuBqoBq/f+Y85f/lmry0FQ8wTiYjVXH3
6s6ch13PXvuhzyMvUfjHpkSjrXmA7QeWEgULmiae3CSZ8IRMf2hXZWue7WRbVgX9
XdqdPmylwD2p38bSqgKmWUrG/DLRyJ9eM7nDK5DbTdLhwSnNlY8TMkOmCB9+auwv
ml7YmK8+DNBqCCUzEiVp3memlcRmTxb7duQuy5jeClfTVJwSjX7/fPpkFpRxW0LQ
nbrKz52W5NolPbTRRUQU2w+8V6TIkxFgXgnXHkdT3u8GXJLERSxFCrqEq1GZ+b/7
QPl49LV/UsT7M5RiZaWMAErQ3OoTt5quEGgXBP8hs4o1wxEzW3wHejs7Oee2tiOs
/9kBGrzAp05NJtaf3Xv+2M4XpUnzPvLqG/rognU0Rp7HdT+im7h+7ToZT8e6cOzg
CC5zTOU+jWDkiQgS+b2VziWaqSdo7Gi+GjVnalh9Fzqvp9YTSlv1asXDcxOXtLtV
e+U7EAsJtIsY8Hr3S7AyfE2t4z7YZijtr9MCkFgGf9C1Y2VRoRA4iksLIwM/z/EI
WHVwGTA4C9HBoDL0iD2Tip+5TAS7TbYJUVYPJ/OzesrNfHIs0uk+USqHFuZjmboT
9qqdlMq40D3xvBE/qA8cx1+Gn8xoQATaI9nadR74MQlSI2xBQdV9WrC7DLI+Xes9
+MaxNtorsp37ZaHatSwJwZiKqVeO4fCeOFkn+aSjqy1O48X/IviKcwkkMMWB9ZMg
ZmqzojNIZbSYAFHAH2nMXrjXzhDAlj2z7wajn02W7gTquUVUikqgv+eZmFwn0Dep
AjFQvVg4SqlT47Z92Elh6AuSolDK0AtcXmuXy5WaoItMbzXhLrqV9eeuj0F6C1yO
K+jnyYQ+1n7TvjG881D+lZbD9ghQ8p+9NHHmuo6dEKNf7WlYt78mech9RQOm9pY5
qMrWYMOSFvPZW0gvKyCxMg3wRIIW6HZUkBHZqdths8OibotvVVzvoOQxXi9ifWG9
E7rEDlGLnlvDHHBfaH70bB9Vo/QeqRrjXfCiclUw48jvzx3X3bZ6g9djxlOwnzs0
VbahvMs/Kb1Q61E9Z9TC9in10VgDX0iDkfufXMAdsXHIU5UPvOb8ahh0uDmTr943
rmWMOGRkFO/h7WmqhTBnxy8802dxZRLdLJ+gxA8ch72M+eCLwHjWVsG91xbkuzjq
63qF6wilY875WvhloutX3BtY8xHI5pGlNlC0cRB+EPxey8O1Qxe5u4sGAVN1PqbC
TOXtYeKf1HCVCplKYvXqsoSO67EiWqNb/m6mTBsanmpiACwA206sEfjxwnn+gxJJ
Ywt/PTBeLo7BPKDgwOI5uVy7W/evTr7Mm2cqXr13Z6d0PaumSHPhi/zBvFq6wrmG
XrbaL3DXAwX6HZk9ZnN97eioOt2WPi1hGEG5CuUmmYGeABTvMNzi8/m2u49PCnWv
AowgLPWJIJcaRBeRkqR25h7DjBpv74Ex8IgqIc96/LFtxGZ0DyNG6LHxnUPdo4KO
iMgUoIqUGV8FcLtlVC6GR5s0/w0mmTOKOxCqC4xPORIPbvkV7OAJvWaaU2FqGcay
4InGpmaZ2SqXDHZSgfNMN6PkNLN/cK9VxE+tGRbjxzIW6Qjuc4fPpuNbV9Vl7t/+
McjpISf9qV/t5Eztn9EwOoFAbZVZGcSoQ90cw+m5Pl02HMHrK5v5uboZuzC6Zb9g
i5F82sr2bTgwICF3U+KEW+RzHejMu7MXBBJLQFwufVD4yBnfAWYFMJtyegDzWtMJ
UJPRs/MYqbfJLdbsbEhcbqAl1pRPCCdu8xxmbQtSpKAkiuIZQfHgJLVjjGnil5L+
WaxrvOyrFlE4U0lxvtcuBPjLlUE4rpP775d/eEe5DqLEfN0LeO5J/5Lod/J7lJSX
3aSp5EVHKeQA5raUHPf2tJN/AJL7Q2h6fEd+IXKNSb8OxUUr07DfZwLiny0OqwXS
0Yo5ZVnu5fv+9ryUC+hVNWAYYR3SpD/7JdIqEChNduB/eqwtmvbyjlqk0olUJu0I
19DiruqTrDkcyAK5/EvRi5hlQmXBIxxSJnOQsRVtLG7ibfG7UG6PaDOuCjE9GQr9
9YOpE8C0+0D30wdMoA4oPV1vAemYPXpqJ7nbP9Szo8+9TyeV2yIUcmBgQycT4cQm
nFpZDJC+X6gF1KREJGNfytSjZdDfE6/ufx+Ou3qkklkQJglk7vkBkNTf7ps5LpJ8
rwTS03N7IsFWY4nUjxIqFzJoR5KE6JfRov5iG3eTQjWwtBKXVWYd594t4sTSfh80
cxIqornC7tKfjL4uqqQi8SOO6yVSXh/WUSX0foUTxasyf5MHIHUKv40KWsTm9ALa
3+nvjtHWi+te4PRJE8QfzrjzVet55HIdhxf3uNoc5OS/k4hom1HFFCBuUZNz07Af
C0ajKp47evqhOAlU6dzYCBYEbuHg2KSUjmBT4Z2IdceN/Ou845BWC+B14Bn+yWP4
+px88JAynIQ8QW0Xz65M8RkE2sKkDrhyaEqzQLQAn1Ffqf6Poq0G5VQ3zzpvx2aG
CLbmHm0HlSe++7u5EKbdkpt/AjHveeigJjE3AwgkroYNu2cZz8TnNR50DAjM8Jsx
0Kg115rmvxdLWDEe/6bEdEl924+0kWcws7IOgv2X4fYmhjJFhWHqW+y9f+agNHSt
i0AgGFFCK491P1QZQgrdA4+5OltQJgYWfH4a1Zr66U7KC6qfEsmfqVU0+e/nTmIR
ZbwGtdlrbZOjv5IzUpxqVfrjnxYL3TBW84lb2s+VuZJRWp8ajA0f17bqCpl/cvdY
duTeN4nMYxqR7sdUrIvqVw6O6sGJ6bRMzz2nDZrxvG07D6O2/+fpXqaNWmGmyVB0
oudJ8J9qp8OwUE1qvXVhzTuUKcdGxpg0DLfU8g/uxyJXghI21V2Myv9ozNBfA5gC
mLzaoKlPjaWuzFZKiViIL6UwCsOL88BCypc7PUhbs7kisqPSX5c/DLdsPVCoeqcX
MHokjRg0zyUGItCqrYtZosbyM5EvrOvbZ9ertK/B9aUwKcdO6DIBlpMBrXvC3waF
XL4zitDGq4tF31vjFkSdGeFYf9G0m0H3suK+turjaoSkdDqfy7/rfTfPzLJoE4V/
j832ZIQxVA7oUuZ7ngHaNhJgEBcQ0FvcbuIUFlJzU2y9eu7uh4WiMFN8hnsiFnmT
GJG436G1EPkdO6RGbYQBR1muQMrWLkK5GySVSgelKBsi3v4fmn2hM3RqicZp3b2s
OT7jEPdT9lHE+cOn/Byo/LuQQMiuTWyezSIFWN3jI0Ktzcl93ulys1mShMoJ71Zv
fgQY9FCAG2+qUkMxieuX0NzmG647G7RoQPuM5WK/5HqUEHQsV6gWE8rVdk9/YKmL
v7FapZn75JV+9NH4iwH+qhlynBVkb7U4YyJwlVNsm5Ce5VQVfo2JZel/zOZXFWM6
nYVXCuaiClyzJjIGNOG0EXpQ8rtPB2/vM/q797LhcCs28dGythog3DQUuPVNyBB3
kp/eDAm1SLDuZ2sZyYVs2EphYh0gfejKjWcz4mOEDTbvdZvvsKj/PaHY2sGWwjT0
poiQ08Huab1GGT/DZSaOlGEeEBdLUx0Kxcz3sz2HN9A8/ZD2tfE/w6J+xwJMjt4t
WaxMcvPWFfxuXm0cTRvv28hXPbZVWWV1O06/qUDmTqyr5HqwlNn/Cz30vq+6RVN2
TpKGAeGuPBa0fMNTT4jlUMnUZa3FQaij4Uu/bibheFPdrLxiTUVyL6f6/LTLigZ4
JIL2QsOg9RE+ilyeBhSxLne2zRZsdF7Mx6rMMjjptNAPU2sRQ5HEfuJZXZZPXTuL
vLbR3rWueVYsJKndHt77fef9jdFQXxFE0ucHruNtkikOXLZea8V1pDAkotR6Paw6
GFM1gYSMp+EH6SR6yxTxoS+q4R1GW0xdCyDMAkJw1Cy9RSm6F0CpnTlw+8EYXdv6
fNW72wJFTGBWCBlMn0svZFj/ugmZoE//Y5XAjyLoOiPdFioXUjNujTzVxa08UPQd
5b7N9w/SmIacrhvPrYzZvs15vIQosnygLl2xeH7EeKzORM7p/3jqLz++jLC1g1eq
zgscIOOJgR3pQtE6gtPZdxb+F/yxWJEuXW97Hv5BDjKFU7hZDk1v5T3KqBBKPmkf
jPIaJEIZ4SZ84Jkw43KJuBl/fvgejvVGTxf7j6SFYYGnsQh34h/iJLkxJ8I55NTr
50ExnqnkKQxrfUsqh8kfJur51XMiI+s6Y4VSNdY0CbhFhZikO8zzU/ovQdpAL5S0
IqkNCX/gIHra+46Pu5wRRSz/5GZdHwPbOItM0aEZ3vVESbzbZPUms2H1744NjDFi
SQzB9UZ8XiLTe8MCxT5mWWBXOL+OLrl/SkANwfzaXdatRMkotvdsHXeCDJ1A97l6
5j9QhOqG/ianVQlGtKBBqEl0+DomyIeuniTB9kSd3+w1A5e8jaK5q8MsSBGGvBPE
Bu2zprAd+28237yKBGsvOwz1KeE1Ma/dJRgmeWhHvEtGj658E6cz6Bq4V+nj5Ntv
ddRsD5rGbhZYvrMuv+rXWD29Yu6l+NgvxwRcSaU4mhJVF7Tfzr32XQKAXLrqXSkq
xc3Vg/eusQr86/vJiW8QJGl56rdfAoxWvCrrBgk1Nf3V9siDebyVMQh6GFjTr0wa
aoajcANncLZ1635G8cwMKClOtoxAjQWd76Fxv1hDsGF7WzzC+BLsDCO235SwCkec
9gw0Wv9Y7Z+vb8Zxz1gLW1ZBrsfZitBXan4yvWeZXxzyvhj5ZK/JNEdddeuklT0Z
cK/TmQwqZTzdmZ18LRjp/WwY1egv3iJ1g1YNAnswDt0Go4FeIsQHLNcbpwVneTQF
AWmU8wTs6m2EEr1PyQxc1NWnRMkLO4zk6H24q6liUiQpqS0z29BIOIxedJyNTTLO
gJzwCB1Su6a4AIbRkSQOFE0YNWlOZvDf4poi5dv+i4X61PjoeULw+2jEYCjNnQxG
EvAMLmtzoIe++8J6c8e7cjqOgjeuQm1eCVI9/FWoikkdoW5PXUIg/Fy6muA6qmTJ
/cd8VYbaJIWfa/5aGBWUjOdrqUF/G1KXUse3QekS+MSR87nFNvuzErWOPrNb7c6n
BpjUsDF6iS7KZ4Jxl97jw5RSG0vaoP310OSXd/Zv9hCpOvKomtfkihKa5cdZcGtB
/zlbuNpgl/JBnxaEZYxdEdsWyLsM9SzvjYeEQuPPU9us3JErVQuV5D7I8NzMYRGS
tIZtZF5RmPjLMz7FAkA6WY7dXcXgjyUTzI44szkQae24ykEDSs+r23TwFt+CmMZH
mTaPhrNjWomPrOImeaa9rQ8nqD4N/R6vzBgLG/5uuCWE8JspgY8+zlPTq+NH7dOx
MaAd+2p26AEuwpeDidwsqE2YEULUvyXX4B2cer941l3qwp+iFPcAQ3DvJHvDpCHX
mHKaUARjfyi/Ti2Fu0elg62qSEVa1yVQ4jEzHRF6q8Aydl6i45RwAUO/lGFjuED2
sx9UwumdK2veDC5wxnMpdT44grrbvqKrYTxftUghYNvKfZCXbVJ4mF21UZ6nEVyr
TMzfdHVVq77aZR2+butKhbDfpXL3HRcftsT0KATt8bp7+khN18tg2wEGdEkQLgF/
zh2RcgtR/jv2ZbUOhXgG2AUXY2Wyz5qRyLXmicGx4xHPKih1OFiLHBN8qBBPTEhC
BnOyjAJyhMoJ6prsGofOZUwnl8YPqhE1FWQjlh01SmvzOf/jiuDDlz34uofyi09S
pMUU9dEbaVOaMpY/gn6B2S7nYg/jOVPueDCP+Ox3Nm+kmu7WIGpLaIbxvgP2k9ls
TrK+v/GZx64tFurfawR7rsLXpjGyhKKvJGmjQfHmrD4rDhQ23z/whOJ5KvbfbWj3
3sjZ6NYNSr2ElcvO25lq1svB0NCd6skcLSQBNXCV2AD8D5O2YPhYMX0OB+pHxCff
pfIF9SVCcj7UaRkdn+j19L6mN6qwFK7HNNUWsjdlrezey5nQgEfgA/bk7TZoZJJB
RQBrZN3Ss4hfnWCK6V/sSI5dVDI7QXfsp3YkT8tmIAd9t+8mDY5tsoL9yCXJ5y3u
FoAPeCiHOfFKfE22RMhd8imB51QzCSt1Ba/AVG5bAksExIJPA1XYfbftAdWJJpY1
+tUP2bhYJLxeNwQPn/9sj459LOnsb+62MvcAVFJORdcdDyEJIy5JyRCCBkmcp8iQ
H+B64XEl5dyd2N1aXfxeuvCa/FjViOY1cD0c/NhDbb1gZzrhOaB7XFaEfzbCZxEb
huPT90lrqubKxkyIeEaRpKNIMPjYdqoYbjQoikmTzFiKtn/rEUaHAOsptYI9RsiM
HbMs9Ki3PfHiBLRGvDWSk+sIQAG1MeHLcNdLwyMaEWsfjweEM/r232V+6oTLKMGC
cbK50Tpp+Qfu8v888QCf4HZuy0lUR59hHpXmJ/YPVg5dx8+R066KXMXwbqV3CTR8
6iVnuFxw+dIYHbMp9/NnId0iVk1pyihbbwxFfhqGCNH1aECPKjt/iX/QFZ97d5Sc
fdbTWxXHu5HThCh0UnGmyiZ41pspsMsWiDzXo5uYkvqdUeCgyDbNZW2qjIfa5w5x
Yw1fz+G9eeIjO72wqJzFi0NSJVBjLOCfn2w97SIJzP7MsfPvqda7sFtzP33OI7t9
gSKQMInBdytMCpdgR9tudLZ+QC4m42G1XOYTz4cmHlGcd+3tfgBivPulSqjmMaXE
Yd8Jg1eQ1KHhflE5Ucr2J1s/zAyLZ2tuySBpXt4bylf4251XnZEAn6bwVmBDtWO3
TZ/SlisovisXKbDJnxEdfyrWmJ/+NCcLZGTy0gAHUnTn8fS5kyoq8t2uu7gQpar4
C1UlRfiyPEveLJMx9svnt7qaCBIkInjVOsmOx3r+zvdnoXGe8kcZYKWL+b1j6vRZ
SynR14eB9O9560hKr+h2OueGXirPv9a7Zy/VBHvt1Xu/AhRYSbJ8lWNL4YyxRQC4
LEABlCKIGEj+oavY/zQV7Rf8hlPouG2qJaSNPrCPTnqCrJ/OZ7pu5KmoAjMcOGSD
rEAh1EVLBXjP6TZQ1N6HX2CT2hZs5MZfSofn3+0PtKB26luu5fiGXmjqraIz00vK
szpngWdpfQN3a5cHLybhYZJwc653mVT7Kax5tlKuDl5XpIsxc60xHGvVOm8CJtKk
iu9dYPWTisaycdQ486In+LM3NR3Gr9+STbC/CblAUsXz7etbT9bip4vezTc9W+Cd
WVWmMB3f/fLN5iaw4FHHt6dB0rz09LqdgNURCe7LB44phjz7rVj+hKuFHIVFIKjE
OYvMp+PbX5qdBDtlMbFiDph7eT1oK5JZoxjx5t7CMzzJNEi9S4Dst3g0Qh7UoGbe
w7Z6mNb+nca+Ln/e2IDvoa5nLrBJ+9w5NYlwAJZ6/0UdP//JOzdpOvORIxQIEbJf
Z5TrDf4YxCKH4OE8ueS2F6sNXl0ouAsE9Ja3KJxXBgSixZe76kQg+DTZ4iZVl3vb
I1JIbRXhN1MDrftZ94/wgogHAMb0tzmXIAGiYNtACfEMWbeX1Y6aeKucJMx38UbK
mHojcvdUqjp3BmK3VpTs8In1F+EZa6fJt0BN9X4grBcJX1YYA3Qr57I8tuo/EnON
yRJVYdK/xFzMA4AVxAlSXSXV0RYOJALyOGLY3LemIGSw1GTsy6dMrvJiRZbRg0X2
SgXqsfLwxGIWaIj+txD1CW/jOu2NuVpSiyIqKhL87doXj4J3drC8oBYE1UC7QOoh
/JKYHa9kGYhfQ1XmQIgfPafEW7uGspy7nrhdjvbSlTetj/345qBuTEpOYKS3QzoE
089YToKlLGtnJ37GzOJvGbzGdWAhOZZXzc+w1rXgYxF1nA3WWWkY11fcvz8FiqzX
LznJg8bogn3TZd781TVmyG3V1TrmbU+jOzQeNjnl13Ri+7FRAVdCRfaeQ+Fpgwat
zwdEkG5pw6PJTd4nM445t6szNyUuZQy391QcGqdRW/a0wXKUjQxa5Fs4by2wkrMd
tMYRjf1qn72s2cWfsPkGmRuEt573YIPNQ9Rwg79NOJzEcDJReSUPhB2t/YIA3XIj
3rNQ0qOVLqbNPOPC7f84DX/r115cJ8odsiNqlAK6YBp35PW9JYyz77UoYvSJ1X7i
ScwYeZ1+nndc2ZgbmRN1Wi3B+PIUAws0LQZI9J/uwHhzcGK75txQlrF91t/nxWSq
D+z55L3nddWP1mySolBdDU1nzYz4d2Ls8Zg6hUcD4NwozuA724np1eBEAIheFcWf
M0rVx9+/JbX0mgkamZcjCHeb6y5ClB2h1kfeavScgvkzSimbvZ5DoyqFgChYP4fC
tRNsqRXCowInWbVSyQWbs7ZCeHuweZaZAkWQbadDkMBhRLHaVU6yNxIm39Kb7OD2
//25Ddh9tFrDrVEHcAlPzJM+5M+OQ/rAb31seayZSGz+yDh/W4DPQvEZE7DrQ13y
Vag5e+7oQQAYqQ7/rnXjRGoTp7q8rH8qXrZmvqsvVO7lsUp+95/c3TO7w+JFHsCD
2qGaZkXHNZJywdiBg42RMOUAJoxlnw/vgwTuZCnsxagi2r23qfu/WxyfZtAzMqpD
4wJkrSAGvXdV2TiqBfawQIlyCwre5c0AV2L+rkP1ILpHz+mQkg8It8VIQtxdE22r
5/5klD18aTSa/rAwD/PNvKKxKPH/GZUByh3BV00WSDpNXJqLO9HMzbKG8NVLTb5H
hqZDXV/71leR2LOMWSXQ6D+xVnZQTGYj1bfJoxPqvm9t6j6X4DPdRVdTaziv7jHo
dIb4Qu+L2sEloVg420hxvzVjuNa1jHz8Zw4uJtZ0pt9qNBHZabGeLrb4lxW3ATx7
q3rFk6eZYJ30MJxKDjGcNyfm/kVeR1lJpZGrh9jVxC1HlP9+TB7G99PWWgVFi4kr
GOv/7ewxvo+gv+VzTILRdJ4lg7gJHmWS+S3MmUEDvd43Oy8XCRTz4sYeN7DbkFYB
7DD46XG5vxg9fPHQwA+INuzf5sPjjSh4jDbqIQsaHVBTZI2wStd5k5lCz5iMKOZu
nyKWK83VmFFsxQq/qQjTWJcgXjgr5K3m2Paj6FxavDSnEzvRlR2CDaQwXuLY8yuo
DAY8Vr1rvVHqeh+8q0sbHxoNMiFz2Sn0Uuz7BcvLNipAXkQqoyfdqN4CceX/ZHoc
Ijic6momOSqxgIHX8N1+zH6b4enu/j30hmTsyIItdxijFTbeStM/WL2qtg7O9u3f
d2mqlm/Lv70eD3pA/tOrWGlSt1ibjTCKgc1AxaXE2TDXYLBd4R8jc6DyzHa/LqGo
IrL8MuBA7xPyZ8jXzVEisA+4G6AgdmsJtSx9MKWE1KYUQfRWpdQzXr7VsB2Biy81
Bty7K2Qx52Yf4RYiSYHQXzG8fTX1akffa5kr+Ku+AApIxoqmwkay1pCGbIsncVcq
I8L1gPN9JI9WMChLCeV3IlqDY/ejWCTcjfNnF9HITdfNGvi2b2O/zkwuUWGvuIrT
yeSZmV0RDVmAYHulIgH2dntwkS5wt8vL3EWOlxW06TaOdSXRgPVU3C7j+GVLM18r
j/9YmThwdNdJI7VgYRtWNt7QN3zgTDEXfkmjYnKoIC7oxcy3iNXOhukeeekoJ0kS
WT6sWtVHQtECVyIpRezIBwTAJPu3dNhB10LHqLR87zWEuxg2mSYWq4lURcXPStbJ
B2TqFMlnbqRj7zF4m2xM/sql7cy3PgpcWCEysmJ057IhB/iP2kMbIRZtaSNukhvn
rkrmjZe0MxtIBCWgfr1RNpeKPyHFZo7Tc0+axtuQc+nRfRmtS1b6ufJvM7BaxavQ
b6zXo5N18QSZwmBLxbI586jDa02M5MwdMooStub5pT1tF9vCP7t2yrfhrBxBZqOR
rjMh5PD4qIrHec/gR5Dsdq6X86BA7M5xjD2PqbxXG0B+mZNCuwsf9EnlQGAeE4rv
tMfLCGabFv7JYi5Va5k8fapq0Wa6hJXo9WU5XIJC0JLbTsdPaBWK3f4MtSqVCwB5
YBhmz6vyn3NrbVnrX0a7kL0Q793VX5eg+6z18tkFgEtLilCJyeWaa/2ZbSMBoOg/
sSi6r1XcQlwlNmTdLQM6g+SUhSUibeP02hZRyPFc71DacoJkx+PXSEq5OdLXdRuO
YjlmYBS2B4qI7Hv+Xgi8uIEvGdOiQsVThV5eWPo3O9ERcQXpNhfhccJKBlLOMZ4q
S/JR/CY3yDfH987Kay0TpVZkQzRMJD8nRy9FY83mMNtI5HzSJEJSdhFp/PjMS6Fl
nSCeerJ9cHUsoNE2ibL+1FyO0k1zzSVu9ngQh8fXA8fsI53WcwieZm1rpMN2ink8
bNW75mBS+oK0Amio1FKv7NXsZI0bZBA1325A6HRh/FNCkMv2Viv8o5Akg3u1cPBR
dBnKyWSzl2SuGSRNA9GACN8hYf2MaAACKg8flyvltgjEXDWhBM06q2UMdkVnk7q8
zduDO6n7irZFk+Uy7vewkY9NPvf953A1qezig4jLw4yolb+MfPjVCMPOhIrGs/mn
AJXfg0nR1fgK+bd41P99gXGXaDtJ6Kj1Q9UO0NZbd5ZJCWkoNAVCpRN9UypqfkFD
Yqx0DR6VY9oH3o3BE6UCTkftIkq39iB3g/J6p28j/57JL0VQf2sf5vlE4aIhqTfr
bK2kMg34+5rwUgHvFMAOpwq59/pwSfO6CNjy0h68wfaLVmyMbbXqSf6d9QNgJva3
IaClR46+AVlEKNBnK9Grjc7dwzsPF7Lg5/q0mNYlhyMvXpPeSlJufamkLyNInUwc
TlZiRHZn0lm0IQq3tbH5l2K4tGtDVwpq+kqK83FXlzxxqyJ4tPwbbPtEk2PNQZcj
B2bwLR2RZ9UHbKNHQV/hGgN6vDUKLw4fz33UJOwW4wAFF/HrdOS5gZXLWCpOOteV
KNZei7x960tbDrh7kW5TUXUI/EBEUMWKEhfpC4h2EjuxM0tl1EYEEIlL4NnjpqTq
WRTKREy3y9ApCupaG/74AV6a4f63PIsxb2eQDxiAJ7kwcco4q+i+Bcc4ZsOV3jL+
bducHJc3Dyed8b2fz+YWpWOPllj0Ihgdq+6DzJglGw16XosAlIIEOqhiX3u2lMjf
TQMWECh01Mso/cXdAtsKHDK3KUXnZB3dFf716AvVCGO1UjQquJCCFYJOfkVdxLRP
pnQ4GHOzEV6iaEEkMa+P2vTC9HT13uL+wrzn+m8ptij1Jndp9lX9AWyhh/w5mD0z
HS3+DTcAuCFfVQzOwJGNqQAlRT3AXpPg3rCxViOCbWMUtK/FFL1IP6Wyx74j7hZf
0FRyQXkQ2f6D9cUVIExfswbZctHOw+/vqNjsAUPKeEUuyzex/D3LRw8vy7vuVJi5
xHvad8F1Mx5qapz1jvyPvFRbujxSaFVoID2R1AIayivZZr4a3fp4yyqYz/eKKEm4
ziX6fv2/ziFYyQYJff63F9svxrGJoG0Ulibzws4eJLla/A2RGnalXby74YJv3MLl
RGAYxZ2kwR05Y0T4W7WfAnG8peAcH9oRQ6Jwek/OnALrIOGPfPrGeHRsYEkk6Cih
Z1EDfTXTAtCZaFvnu0yApPwWw2KhC8IHmAjZNlX6+W+yIi/lKQ8IkRLQkNc05SuI
Ot1MB53Ovz/MX/KB0re04+2tYCQJhetnHU/ryQkFNw6Mqrw+WWgInF4c52rXdwt1
3JZSm9xWDYijjATysUVP2kuH/bXearwjFmK4J5oEePjSb9quZKXJzAbljYuH1BGc
4FvGJxPcZjX3qacitFe7NGWlPRkgmFvOJ6wUgwD+BvXX4OY4J8yrtPaHvSexN2xn
ksi7sPpGTzoPVTyL4GCjgFrM34mOs8vEVGYllf7mvD3lCEy/Wcwl8kEQiFP5KyHT
WfkxNJbTNilDjYm9b/3ctV5h6xCddxgI5oCXvsIFwb23qfWnXgewlUlRm0aYp4jz
qXn0P4+Y7APQjJE0YRVGios42PhU4P7C3F9XTDAa6oeSG9JnFL5ZGGyBn4225tVN
VVodCjdXdU7qtyo+yOk7MAxFR4p5HkK823LW3xORlWD3dOkK+4ZM9R2UeG09DyuX
cjpAvCKE007M6DdfjgvuKI5gsL5RJ4Z4tt2MmNJRiukGm1iC/RbKyLOqTbzEGWyR
TQ/xjA62lm3PaSFLsPzgBgiNUt8EXYC0Xx1wOhdt5aeDED+Bi/HcjMbF0HAIYzYw
NJlfntub+VwqbeekOIq0j5cEckhRxIxDn7pzIIbsQa8Asp3zbCka8qjBG0/kSQ3/
jlRKy+EENRBfWYFATWWNzRDef2EGpZrYfhx8ZJstefWrXU92T/B5bLuVuCa+vgM1
pwDJXLms+1XC+fTJzQdhWdbuRX2noRyMXiK5OjR4V09jOVsryLuxrkfAAPa9KUuG
BClQY4wdlehGSkRD0LPVx6kwgqRoukF34thpuuMnlWmeNIfFfyIgkgDWZoUXGRcA
zXJCxSKU4GEHoWVNzSgK8xx4Uk8SdfnxnhN4npDHTZnAEPX7jUtzHHgSL40jlYlo
G7DdE0cdekmSLp9cDnrV+YMzalfYLLf8hhtMFWJAdDzXnmuqzMAN6DsVX6yGTUhJ
Kf+N0h/IHfp/aVuUkuVsgP+FLPp7vGFFR35bLWk7UTkUZfEKx6SziCEe/RxRrULv
d8uKI5755hCS2rwXZJujFB9rsK8YYHJwoN4V/xmVoqC8RmfuS9NLxX4UnRtDUZNF
QDPyg4oCIpeFBoklx+xBxV/WCDdkMGmRTIuCOAxzSupwfLUWQKPcaVs/wTWaVwlv
Kky30LGnQgemke2wRjZVCSlJGsyrquINEyJp755ck4Uphg6oYBSDA1R0vvGLUuA/
a+dKj2tWJpxTYa1CIcC7jBjfvmDKZ2DqgDSlOyc8kRFI9TrM/bli2cEJi/bID+qB
dUKwKZET74ANhilrc5I3YfLPYxBdZo4qk2LtSOx9BAPuaNCBSEwYWt1vxGN5FClT
LFq3jpPr4GuoAEKToxGepgQn6e9s/7ETQsjv9+o/3jvXzvEyfRh0cAmYxixjTouy
jNO7HP+9Ik5lerns2DKbfVEzwYvY/veZAFZ2HHQTwH3cn+fJCXjGeZyAPj1VKj8s
XSSMJjxsxcpwHVYQZX+kUpRFnBI3zCI5ducLaW7ir9obuKAzsfTLgfzXg4jxlmBT
PesPeObFdbH5fY4a+I7uFmgUWsytURoJ6EyxNNFIR2zxHQEIec1hq1DUCIDMfmxX
60q1jR+1YIThuatoTgxVHVtx/KHYLZ0L7PLFKfgbLrcuoVvqSwiwfeNBCr/9q6IS
CFaEkRpMzdfhrtRF0E1uxV2E5ya67vTadZRa2FSzOMi5pzXg5GaCHdKfJpMig6zP
HprWAAqBLkYJKSuMaZ/cxYQRBWkr1/ruhUcaTvas3cKRXnwLHTlh3BoWepXnHliX
uUtbC0Qov9h/DqCBljLPfbyRkAab/yZIwkD0zKfHoqcQ+lhB2qMyS0rmMed/1NjH
Cl3snf/VpUO61X0pmW1LBTdvKWHIyiJg7JGwCC3k2jXHslxQV7LstwI6ZCLEN84S
T8F6QjkxpLGDSMhRulj4kV1Twot65MWuFqncaXkShOmshJI+gvwEj8t0KAzNQ9JW
9/SbFGJisQJdFG6ar9qbuWAzI+jxp1l5GHdSqehysSQdmpWwIHz30m92rmg6p6kb
6fYzEE/3b2NmDcfdHy3Yiw/RQSpJolKcFc2u+0ryA9lFv2pLjLydCJ+ATUIutH37
uBKhC1e+uo89wJQ2Hg5bkJPejGpvy6kye7D0sAceWUqrBhc5GIE3WPWIWPI1rP5i
KpiTXF4lPnoPZp5rt2WmkIxGLrP6CMfH2EJAWEuDYiNZS51zwo81+2TlBA+709Nh
PBSI3PnFL8BuKqTQBmPXgDs02f6hMp3azyxaEGajpLBWli0GRGcaVK4TWAPDQ1mN
VNKOPTyuKOWI5/fpLQjNGSIiWV0lksHI4mQVYOiZ737M8MgWgy3Huu+lkCiXt9XF
Jw/qgTA9qK9VqCS4S78rWbfgISkxynJDGfhAg5gQ3Z4wmckl2MUygANt+ApfKRcS
DsUvrdXB7srBNKHDobbxTa6lJ5JIgT32kzj8At4GgDU3XNwUz2/QkADB7sJviqpb
t87oW/SWGIkEN5Xmxgyo1wQdO4uZsqX4LCP3It6exromEZzr33p6ombo3To1B87e
/6JFIuWPTstlAfj/Pp8pFPh4PfEwTRrj+aRO9z2aQuPGfhYXdxLA+dXJwLEWQljW
VZaaRb5m8BXugralVyOxR47jR7SLTHvKecqxFjpC9Hn6/8D6rdFb9ZMsvfvXmMkB
Y2IZcL4W09v/S0lDhan7h9xf6vRr1cJE0vgh18cx+KDN6Ja813t6Z4heLCy9iwEJ
56s5oyyNod6ff7qnGKss8RcIKGyynWRj+8zdKRu+Odc8RrKQ06oYwoNCWbLKiITr
Z5GPkAi6pG1pEE9dXRYBPtKP1zwrnsOMirs9eeAfBFmkQWRSO4jhh5ptv057aSYq
ImoYzvTwnfSEFPnnePYa+daIObxvCYMkO9NsTKaiPULonzlw/b7+S+2PkHsI6h1T
tG3eyeKQLy+u0ZpUrFcjOl3xYJwIZcvqqefNn05uW274mSbeAnV8FZXtwm7hqcbN
Kv4k+IkeauJh0NFRT0crk1/EVk03XlunbaZfVhxZPTm9Z2x1EjVYwGQ2mhcSmk1c
TrkNYbSVQ/o5w3ZC7hn2QCXla8p8yFFBIZkKwv2ehvS/bY0/S2rTeIkCqvkOIOOm
HI+KVnXmz2G6OyCMZUnzaYdjuD5c2ZKZNcG84U3btwM6m3Czdm4PP7bp76VtWCeT
kAqEgaVTATNfxPiZ8LOXYtAUg3MgROgUYunTLHCgIlBAJf+UBtYHeKy1Txnt/kxc
a1/ZeVKwcWg7eFYrIS1SuWoUlIO/kY0cnSFs+pQ8eCOUfmjBsxMS5MsMuN7fPU9L
d6moUYbjWFSLsCvjsLTfnBOChIksA8P7qESlX7Ipr3yHJ1TFEuo6xjZRBe8exk4o
UjD1f97w0rVK2W8AX3u+IsaJVnocExThsRQIxBMSSOqCBQudWs7MlKdBC7xkhov+
muPTjj1zJA6wtHVbbWEZ85hTLsWAEoPJ7/NW0PCit+JfE432U5jfNMvYLBYv7GPX
xM8eaZz8i0+H++QgqDwTaYl+OVtiOyEVDGNrtai/d4dcLFzUnpn+NjqJ3l9sGdIl
Kn3FF18f2+KPlRu84afN5In53AyCcCykSsEoz2MigrmLv1DBS2+sDZev7yX74jao
sGWkc86tCLYjOtik3KSpx/Ovz81Rf3Uz9kmq6pBzcg/59x6+E/qyj6Ed4e6JbWsT
l5AwCRAQGUT+C1LQtedpRFpQArTIni5Q5+kGlzsapz6GPOD5TSKRLjHHXxU8ISzH
JEBGbq0rZhcMxn1S3XG5SIskRUDbW1DKmj0Jkj6xVX0Ie0zyWUdgFIyKaCELtDtV
EyGYHh2w+BJDhNuB2aa+cyIi9JYJ9z4o0pKxYdwTEMUKHFIF1BpaMe6VIwdpKUp/
5dVKdAZKf9DcuqRikNuRdQyp7Wn1UQEAZ3JpCZjAtznYjocTmmqTBftXXwwVWtre
HZiINFKNQcYZIxZWkdLbLIxJVazUvbko0NYQJCbisa0UYt1VePoX0AYZTCy/HUsl
+JV8JJ0HFZUX6n392clgO9kNM92B24UOSR8ddv0dftY1WthwN5Yxs4VRYagy0Sqg
9Yjjek1hDKpz3rEmhlGbG7BNDuEVGtQXCPXPgXDP8hKuAi3AQSceAf6TN5qg//rW
JQ18n+jX7TckI2cI7Pbe5XgQx+ihwCE5juGcK5+E4VktNBOGgcz5jZZLbjK9C+u+
+6/2MQ5FlfXFygS5XKVfvNDJKExDG6y+zQPIrRe3Rr3pm5g353AKl6/FhpDCQf8p
ZDv8S34vaWbaFsxbKGAoBjZ4eDNexLNEHf29ZUQ01rO2hDBgdjaQcANJDa8Ljkqg
LsS9Ohz+rQu02mySVYwAANzqlAAXgxEvjj8DTsVZqh/Bo25khWWYVdiWvw22OJLf
At53zXbIspG2nz31LIg+8I8iUvqV+J0j/V9G7JNtpF7Wfbyrw3e9StuUjv+PiRcN
cz6IWhiE4DoO8ZHZORYW4aeihQysxnZBMbQS+IE78LPtewwXP4slG0KComH5YbWS
+0LJNFYXGbpGp9Yo8YDTlbrxPo3Xn3ZLJvRBIJxsYqlajEjYLnQ2DT4k/uQ6OQJT
+l78DfDFGneQPUOToSUtNmwmHvWB4GMWGVgPEwquYsAcQI1cabndL1THkn8y/pFJ
Q8O31F64d3XRGSFuX8FkgB2zA3Kk2Sv1uQLnRsfRDgkBU+Jhqggb3WjDyqBgPsCT
hPBvpS8xNzQTer1ONw21p/6mmxFqOvMLX1SKmpwCVpZ2lV4eAKfWuCtlA60+8o1D
wxsk+gGkavl2XoAliDUBDGdBLm4Wd2FhPKFpSe2wp3/jeU8PQ/Wr/RJyD6DTwiTK
QwPgaCZSWngVeCXKXZ/OC1CZWPRHu6QgTDnfDQaOitAU6/UuduPEBJ25Farn0pRg
j36d0ENE6WiAllzIX0RcjiV9oFb6WtrtwZuHrcTA1hEqPfIHiMkoLUArhyr52tBH
l3oJZ6NoD+CVH5eCjsyUH08oUSn3FKkZc8YpxwHjDkrW1gnkysp9HUECV+Ws8Nm2
EBMlHJqtQVBFhgFqkKCb8ynCcQqlrI4C845j0IirYRbH1uwu/QHuTXDQ8N+3VLxN
FK9P/IIjtAaCxxkfZBw0L8E+1DZHGx3w40qM1LblLv609fgWfVzAY62TC/f8xBKj
CD0AkPbnOK9qcRn9GrnwLNqfYS4VcNH/5vNjm6bToMNHTmKMFva79cK+RyrvqwBk
al72uc/ivWQnNPumbiHJdyhOQyGuwE21PGPLwsMxx3XRmA5s19Muo8oziiWVG4P6
/1ar7Q5a2FLWZsUrQ1HELgqGKP5Cn2UndEQfmKs5PEiKlP8Robq6PBzbF1rrawvi
tpqlvwy1ZCQ63i+2sshgkstiD52j4jJAyTvD4j7RdtIaTlT/5ih1MvRiAzeQgEqe
r8YWfS7MicMcXSHv0oIgFkXYKhAiloZlxT35iv/xqPtFcOSSf5fo0xMQyCv0FFln
ByvPgjVwrQS6jPHCkWI7RZkNZXqsw6pfU9rx7iAQr08H3TSoEqy992/y9W01V/Qo
vMMlyWbT5moe3lhbTWvkHyJS5WcCmYWv8E8zQb4+TUpKo0ywfjTN1ZvDWxJD3ire
D6G8KwG55fEhva4eyzfLLJ2PC8ZbYUW1Fl++XsozxcWKeiCvzbM9GlSwoI51pyTO
5SOe+PNaQqlCTBLqUt8fjJi7QVYrW2fAn1iZKPePaWIWHPqs/dTupQwOF4T1fysM
pGMMJ4dHCGY0DITtJxnJiYf/HKUWANv5xElPWmwLkrPA7hIijAqfl943Td7lfihV
yJLp2mKozym4bSaajsrboT4lv34n1jF3rC7SMEpNG3XjDXNafSdt9Y+uXfyB+P2i
vyt5kxJTxf8p/d/fHojF8TzsD6eHKHSxHrdw6d9/bg2i7E64oInJW/yJPrlq3R9h
DX1WL7p3xFyFRo7iOts07Xs6EC26BSkpUZRSqszYV4lA9JVDrxiLNNv5UNRPmIPR
BDS3R6GLP4uhdkWCvSA9MjDm8x9iH8NmK9sJD4VRVY6ZdoLbGgO33YiWQrsolK5L
Q9hxdnr/uarG1BefIyh14Kmn506deKb7bz5y/KUdE+Oe77+GojrSSAWSdb+U4hpQ
TtM7FD+Rwek8tpIvtfFSEneKHK5OVVHwl2eEwAQbWUKqb+HIs98obsUY6LY0DitD
cEZ/LwEoJ37A4a2aNp5qxsuV2wNYshUFRtmvOBONtZbzGeQU2sMliC8D02ra03yE
Tz5p8kPF6iTWcHKYwVNgi5txHOxBzukJvBIHi80TCnaeRjyn/d9hIYp0dAhbFmVt
ilJU5/7xZyCK42lt0f21p0YaStFxSUjyQZvbyXFdfkd32fwbo28FfccL5W5lrfY9
kvumvz+7vqBvSKYWUXr2an/iRXQmdHlg2UMLHSENKAUWAMsiYO9QsygAt9NCoJ8j
SL1ZLamsyc9ELQguWxM7zyfze6TJ/VcRTKJ4Ity8q+fVgKJBaJPPfCtCDHzoTnsb
NMqaqHJM/L5HDLv5l11vxMkFykcc+ohPVDYldDrL+T5SIC1no8D6QioKlD6/5/Rs
mhmj3/JKshUGxzcNBx7xwtHggwGs0kACe/aRJLUfnsBCofSuC1W1KKmJF0NlDxDy
EWa1zdEObjWXQqjsu5nzOVQnslviih9iN1eebDC58gjF64RWF9spoObvs5S3s0hF
1bKes6PysOlzaHqJrw3os2j73zvdmh2tMfFFEJkD3rNMg2BEE2aj27yNQ4Ga1euo
B1X94Bv0gTuaNaCOYXMdWt4oaVQ5rV7xJTSBQagcse4Djbm2m4zMFIH2jGp2ppzR
N4/Xmi8RVhBv05x1eeyHlbsU5oKNAd3mQyUTlUWCb0g/OFOGxUD9kpPfewr593J5
xiC52WwLbv3zE2ru5yF42SSsJ3bj1YihFV7LasDTsqm32xqRuyepLcgMbIgKyEhZ
oka+sA321WA+9fiLBS7/K7j08wQ+1UtuYXmSmK5l52+hKU/UR3BmJjYhKRw1gq+s
LagRCT47yEv29Z6M9WDy0w8nCtQVU+HqpShcZNdeEzJcpW0/4dis04u4djdYs3G3
EOeiYEyDSJE77/HKlJgHqpnQsynJXwbC68o+OIRh02R29cDJJd/0pTYWmm1folRl
4qHVTRiw095jLoYaFap7+3jHcfQCyOvaq35/RAbKK31O2K2mfGd7FMCdOwpoRF7w
ogFrtI6orgYdPYsSWKP2sAiS9U8jNYR1HcuM3CW6SlP/xksO1MBNOOqg4D8DHJvi
y9+T4I6lS9rqTmLACPvTy2TAt5H15ck3Ta6OsJLNNy5L8LqqNQhmyDabvgrMXuJv
7ZDYBc9eqfd493BeMoXsRcenS/CaSgxr7lbhHCxtCFzTrAum5xoUee0ffRFFQX/Y
gTNFfxjb0r9j3O+A7ZsiNiGKtpkmfxNR96crLt/AHaagvB8P1hsIFqSrqA4lp3+i
ORxkTnqq3r6x2qXo+gjEuRTiXoGiEReg9+YcEx3wBNIEGtSu0b1K+BVjP8JKgfSe
oBGGEbc3HEQtv9IoRMXp+yXmtUcsuya7KnzMRKHp7VPuJv2AvX7U3j0SDEKB0BAb
/k/6JBpQRPRxR9VOLz4upxqo9E8Uw0p/DQkTJ+dBOIRcIMZKPAbQtdHqmJD3GVMy
56+tSgIjkicQ22svXdY3iYr6onLSq8fJtWd87A5hHrzqyGQ7xoA1JTo3X0g1w8xi
Y4VjcgLjTpV9ME7Nh0TmBNEz02dUI6Ai9SHpEDr8bJOSDHLNcM95PckB+NdYwe21
R8wEJ5o0CIgZKAUfIUhKPoyUMgA1+7syI79vVYdkEoDiGjZSIjr8znm0ljmdoRLw
bNXHXC0UbMERU2aKfGCN1SwAPcHsgBoZJmi/xgHCgyNlHsIFskx7SRwwryCsb4dl
lu2h2eUVD6PzGeD2Uk4+Rfa/muP48ILDAFvNXoxcWwnGwmeVSp76LVle+qj3A5yf
KTjZkLSTtDrFXfJz/bwUZlVfswWQY19ZGuKgpFUJ1OVIfZnkMLCA9T9pKo/vFuNT
HEAz2kpdd0P2eyke9xqFr7OnGWoqDAWeAzmxpp58O0Kt0LWv9O9EvLemm//7ci1h
KF4ofstU+Sw30fQG+GuPUly2aQ+e+aAtTQtVs+Fd4yAuZat06eXfWkY7owcjNHTL
XOt5ANYRfn77VWK1W4ALubEVHmtzIN3TktS/Yl/HC8YFSHlFhrtQW65NeqvsQXch
sXeoVEFOO+CotkuS5U7MNbE6ypIUU/FyeL8v3sxw4AgcToGQblfJfyEU/8dozs1n
hSMFJ0dfwO6P87y2qY/f9oQlnG54U/lu2JZQ9cIW76kBXykGvYe4JpnyuaNby8vb
1C1f3yUHeZiub+A+tfa0MQhJ50aFm2fEPRfCeJ1nDLprfBCUzvS65izTgHy3p9sD
J+1Kc8v9DQpKUVBT7kVwkHlXDUTsuRWgMBHAWVGiXSPizu/Hb1XJSXslhg17oZ+Y
HkzZMQGIVhDZ3VacNnRXmd+CwhXkeja3mvVtt6+nVMAt44TWQ/rEZV0TZ5l7e2b7
Uxf9SdINpbLGCQCP0fzvfF9oDeDfWtI959Z3LT5xiUQvwGhb0KQmuwBCfFycwEEN
MIb6MH0/7Amdqc6j8zgbUs6sNCucm2aE9NSAJAjYeDflRUBzLPZZ8QcvA5Mi8WYw
syceGIiWslBNWWyvvIZMDxaWsWqXZJg+t/ux++875T35qPgObu+QXBdfG42S64Mn
FCobP3hGjPAbCT/bpziGbyDwamyjU4j3Jnnsrigf8r9YRn5SeijbOKSlk5B6x1jg
OKRu9P3hbT2/rChlS2tyQX7W+KIEla9fB0kJepVoaHvmCGj450EM3QPooIy70o2c
g5oyCE5LXitJySkDU41NcvhfG9nasiRFKg7JuO5+htR81tqYGB8wXqaaK60S9fVT
Ox3SYykJo3U3YJg2qpNLBt3Nww5/PTsDDcv9Rz7Rz/ZjkifuA8kfd8KxDUY9ldmP
yvo2X0FPx5Us466kCqlMe3xBjQLXyv4zqQ6HlRoSZ0w7V6f71X5DQL2DsM1pdF/P
FaWDv/JZlPfVPv5xeHXFfzfPTNjrFSC/i7iYIFB45mYfFhKLNmN4lYzG9wszM6WJ
Fw4icS3Rn99shXpelx4Z3Zus8/JHgIFiqKr9AfWsEOcP8sYf9hpCMqbPqLFkpIys
TP9pvUelsY+WL9xTQIxcIHjDusLljM3dmVMD8SGpuSJ8YYXaoiFmJktwpWGIR5r1
4R5/CUzvrM9Y4PBfHPgQ4QFA/VoSDshkhccOnr2ueXKYTXn5blPfUais4wLqW/MY
1SRZ1KgTPJpdOEChh9qOARcypTNp3tzDppKJ1U9oMsGq+8dc1I1ko9ifm+c75Y6B
3a+eu5JHSOUWP2pVBnHKCR0ZkbRm/WAR88oAsiARaXAMeB/KfIUl1O0N/2mziUhb
y9jPQyqNRPuBs2ps3SNPZBkoaOkHnPn3T2nbEa26VtPeXGg2sEfGYYXqfKbrJsv5
M1EnpppFhAJ53hWZsC0EcpMCgMFkui3yfiN+56LFW9gw8fNqyWq5MhquGtjZL6Bu
OrdZ8xvGKl+dqpY3NO7voK1F02oaxnKJusZr+vCN7m8kB9oNvbO5J94KMl1MRGot
meqH2nN6N2OlLMmwHTiE1QQUzwWlJkD4nXQd0/Ea4y8UXBMygsJdDsWO2QHNpj1F
MP310dHamOF518bTPdZX+1bNIIN/nJJM7p7l62NaBjWigOL/40p+HBkqKpWmFsFV
1bvAwStZagUCz2IH6MjxBHZZr6VO9EPTx+K0vg6/C/I06Ji/aKo1Z1ROW26HSXiO
Z2p+LxjugjQkKuHazmivSyRDg9S4IGe4+Wc+MrHkwT/B5hRZy9HimoCzJCKnZjZP
njQWjglMv44imnTJavizzHDakHCg9I5+MrbVeAtR61PZ8UE6mu0FTu+x8h/cvCmy
84TJvUZC7lE81+zdYFfIy7V1SQL/sshMgwbH/lbjqoEYuzb/NkwlgO/KeMPgvI1y
7s6rBo8IXJ7Z4y2SHJ8HxhYdTD5a4t95h9A0vQtHgyp7Xx12p6atQYXy/Xzo6FHl
E4c6zOUMU9ZkdqHqh3c9h/DlRPpjg/cZZFT4FONLOfuQ9mZ+Y4NS0Zk1RlmfEd0w
eoHzxqDkuwx4MojuHd2wR+RSpxDRRrPcJvztc7PNOVjBdDeOXN5/dFm6N8EX/XZA
OuqCCiF0Varsr4hWtFWYnSdptLA7d/TpHCCnr2WB8LfqmQeH1dWV3hcmSY4BiPSu
o043r9qpafZZEqVWAtgrEdolp43hmjvJUI0YfmbXEUcN7F8v8Z4v/PoEZMNJGTIo
2cUj+SyCisinKLA5nlpAgHrzhI6yAftIP0OwBfqTXDITy5BJsdPh5i8LCrUoeFYZ
2FnM3P9G2hZL42NAGTt2SMTccw5iZpse9XVvXw7/l7EbezVcNDs/90tKnthqkReT
9B1v/cs5rWVMB+H6ogzR2/KVxvYLHP0b+OLfF0TV2q9DCWlXoKFW/+U28NncOndZ
qwrugkRAdDEsUFquOPzYG1TvNa+pKpv2TYYf+WtzemAriM4uD6yFzRUhbrgqKvDk
d8uJxktepmk2u3AHicc6JArtKZ3IZFvZNjNQoxOs1S6CI/ITEyfNl406igaXjzms
l+HXYJ2IoPY2ARcZ2eiz/tpQ/yfKswrss1/hveIpNrLGxaYsaOIBdqsyommailQc
yd4eB0Qihe7bGGhcFoVMpaaYkv/tA9coFtqCiu6H6FXuJsoIK0WtQMBOpfy6WUf2
kOtT6+VWruQ0vP4vCiOaFMxz7VZkclJnguQt/LQZbkW3VLSK1zahEwJSZQ0slQCw
tTx/JiC8Vn6Xe/8xHrzzvqtcX6keTwTYizzPOUEvyt77bg/oqWNgk0FO+AJfGIaA
wkmKiLUnDg4ML1Qsuk2iwv5NociUB0qnxK3oXtXfHHekBRNVkMUnr4u3+D5V2A/T
RINP8VNnWwHqu6xr8jlJAqZryR8HgL0d5R7yNS3+Hr30H79p6Zn24LVygyd5D2Q/
cw3cUNC2YJB9RY4nYI6Jtzrb1XnoNI8O7grltbymV7It6PMc+0xayNQg6YUXk9+I
2mvxKq3SXgCel3QOjDxiV+ssC2HMr4Eq/+bz91F22EwHRwnSVLH9zLYBRC6xr/PW
IabMtqaBoRXNIXzmfY6LhBeVZP4drbjlhLTnpW9immj0W3EONfT5wW16qxUxQVIm
e5kmSprwkrxxSjxq9D9pDzbeJFDgqTAN+0dkxubnSszbgJptyl8PwgDirT6ELRzo
xDtyz2wuPG+c+nzki6PATUnZXTC8mPARfwlF3Hv2e6mUUIRD4IirxtsGx3bMK6hG
/Xwe/VJ2g4Td+Vp5Z+3GUFKj8UfSFSYvfXh0QqTwDMuDQgJ78TeBbQRiiFGig36d
jdLQZKPuV1DwF5gPvnJ2QJbdcgWQkX8P0EHWbVZ2h+/jw0Rq4wB7PVJ5zQYwxvW9
BTn6sNcDQmRjTX2lcNVQGAOafbvONOjlvx/NkkdRDH6YrAUXeUQGee1C2njnUkjF
KQJU+wZ/C8eoHeXt16RNWP1ENaljfOcd1rqCHkv+J1Noe9CyxoQpDT3QVVv6W0Ao
grQIQZaQF2eHE3bGobMvqH3C9zs/PSsgON0TG2h2yKfAXjH1+Sol/rMEA4uEy+ZL
pB7q9O19KqIRqU1Bya98CoweDLzmD9OVhaxj0l0q4nGqJzKmNNa0E/rCjbd5U+mn
ftxCKwob4DGhgVvon/fwhlia97BavvuzLNMe/hU3Yb54i1AxAlPKCmlkOQAoqKlL
Ydl3MtnDxYXakejUm8HA/t7lZ6eaPoQXhewjQYl7Sku9O8oeWmaRb4GC1KMNyhUd
kdCa6JSKpF4ZNE0fZ0SWZyQFY0SDyZOhCZYfHa6wdssV8nWfXxHjUpUVbSg86Xm4
e1TEnYa4tAFpBovzQPcAgqgE05bw7NVG2+zwD6YGKuBxCinLNP3r+x+4uB503h6t
MRjz7ec96l8TDsuJqJN/GgLO89nGNrflirTCb1BTI/HZF27fgZAsD4MQpV+geQO1
iOHtwc6KIefuDy0S8SBnKHtW0LJGzNoT7FPxVYefLktFRLgd29qC5L9yQ4GnH+R1
ZrsWLcx1rC/AxjKKdglR2O8nFKIAEB3PmVKjLSpZPgG/9TPtK+5DqLn+eHdMXiXx
7kacorYEBlc1WUgY8O3mZ8KnYrWhPlnOpwyh+LqwNzRAiA2uAEBUdB573en3IskD
yaEaEWBKbV3313bOLF/2T++SF4QywMf5BamV6Sv+F/MvMd3tbbZKGK50qlm9+jZg
Yd8T2CyY+n5gmdct+FdWNzTn7WsGgMlPl2spJrgllNoFq+SgbaO+nHBsPllxmUQ8
hQjS0pFVhNUQYi74H1yPGLXv6aLxNF9yYZ5nRrhXkfdWJMW9p9iVLt5kyexY/MNr
OwxD7XA28d7KD75v+RvhZlA3r8Vwgx4N+K/eRe0gyplcxs9nIQdNPi4UAziGnqRK
r3aX5S++EDNfiYaIzK0wPsLxyJq7YZ3WxtvHQNR7gtLr3vNyDenmS5ZRFWIbxDxP
Xyo+gJi2wPLE1DMKuuLRniGSZ96MU70D7oYc2JANrfgW4uWTMalRqZt/Yt/LsW3T
EJjbSwNaSKqkKsSyua4T3oRDQgK6pX8/WY5xXDfZ2qeb2ffMJLwyfa5CzHax1nKO
aZlVB0sURegvERaGYHBtn9WO/9b6ycD9oC84zdiIdkWXq8nTukaoTjduYuh7mkRR
VP1dCBZZkJMC59aDGBY1L3EFlWICN8lTJ6vEbRcXkRwwkTLGpOP8a9yG3DAkf1gJ
77v/ZW8+Fv/mDXrs0eARZfPBhVGoxU2KdkfWLCrB/VIyAkprmI9JN7661JXu0b8n
z2f9eIWXvWMMJrhIRFPiZQxylKvlRe68S+72QpvQIb5+8bEEKVtXit7eua89IYIY
h+HhHezSp3C1KneqEgA8VR10vZu/Sdk/PHvzAifr15jjsP3Ht6ewRJugsmzEi8PS
LJDsjpa5NNUZ/zjzeU/Va8MeTwSMXERv0dIKORs/8zaSqaXMtcSOEGzOUIK0mBub
wBbrT0B9jZYSGFFI8YtNN9V6ouUnsyPHaXopDEOx9O4WEXxZR5e0vdSSbGH2mVyq
Q6iiSMgP2e75qXM4Jbg0d1MDkQOhdSe2rxagjt8lSQK5ueha9vXm+FGEbJNsTlGy
zzWLNHlMc53xtoT7WvNMv+BKST1VhSJ2/wBsMtyZfS0rFCJTp4zklGbiUhw4WJmU
4azHYdIz62kH4s2BUcr0KUXe4K5eUrJdrYigoKpkEAHzzMFASpH5ZznC/AMcFfhF
JEeLm7TkjvjQhKZB0F9b6p2DL/JfzoOJSX381aieg3NcLRQo6OOStB+dfuRMVOzh
DXhyMM2nDQZ1rtctu/rQcN4nVsPidcg+r8oTp+h7/AxruSwy5tUXr8hTgmlvBryT
peTP8oZOpVXptGT/Ru52bWRdCcTLgCaVucL5sMACVtm9l7UkyTzfBKDqfGc2hFzJ
MHdBv4nJE3FKPkKhjHrYSTBlDyh5R4vJHjo0ebL4g5cOmb/zMbF/gZCQ29ADm2OZ
Hh1kmNQCg+EmWZuH20NQ+zfpz/filn5T+Naddy0UsCfoaMrkZBf3tu1FyEeQLolr
Tt4S6dUVlaV54snhZo+l6ZFy+2V9/OCWmGpw8zb/Pa7pHhPH3yU/msBytk14I9ZK
22rO7kZob48QQK2vglwBT1C73a0HuVE9pPX9WkvKP71fhsXrqVDZHvkvy0bGhFoC
ZLR0u6TYJ0OwGw+WW1vtyqrcN+tb2KoKx6kVeZlTHB9W1tG5TEg2P9xO3xLV3LWb
S7fRunvtP5m/huDu4MKsTrlOHRwYNBoCNFFA1k6lGvTxV8y9+ebaKUf0sgenE2sW
PIE+jgNBu+5Rc0cL8P8QSs/rSkNPUIgHqg3Ogf5X5Uv9CM0gMmLi5ToMeRqN35GQ
pw5cdWUwpAWnXSoe/EI16GEVBPKK9TKIeL6tSqFF64b+AosxufKqujPpJlxHoyvE
wJGYcY4k9W/kvKCpARHij5/hWwN85oEyc4ERz42kOjDdkUyp6GKtUMVRzhRZc5ET
K/BE1As6sikK2vV6o3NdSLrD3tUUdbBi7rrlOTanmOszKFCGAkdGYjy6Gqxg1s2T
Id9SGqmuVjW8MChwtI+0priJgXGpT5Bgs0jBW88yq/dzyNpD15bILZMuoDisNUBm
9GHZ3KvvPVN8AzFlIdEOyHmdm4KhyPrvTYZsshblFLj5UBeB4ewx76GxqNjp679t
ls+TAnV4M8+PUKtmIwPxwHnDZVWoFpQhGsQbY0GrXElG/qJTUgLucMBRSg+WlT+Y
plGr9iczTSRS1lA82yW+t0AyqIga99iBNW+xrROAb7XtYztGfuJGh0sY36WX3EED
2NUaVfbXJDwkAmMSjY7kxEbz1HWleVeqpdinvOHBhvv0zqTIqllsNBIk4A8WKnhb
5SYKTUrobIf8+ul2ALWug9fXPXYfWSA4GrF/jSd9ePNVldmBr5GHysSWtK9rrHUZ
FfFrlByVghnBsIsUdju7Rrp1dKY6E2pIJNXgu+eBeMEaLQjTLDjNOoIj/eqWlCha
lTPONQsldjFO8ko1vtzV6iiMa4IRY59d1gjCHauKiJw6q0gjnEH4/6Ogenqq8XWQ
iQUgIr6V7f8IL2IeJvgzx3te3XIvoxG+YAjqO42VwFBO5GAQKcLTdbWO4YPQWmXF
suW7vENlVSWR+hZJaNNhGZcX6oYXhnaGI/BwvsrOWo2VoSrOMz1gYhRLkCKeTtop
rRHy6s9AjlV/mh9ApI34445YXpyuE8G/YyvOYb65bvaqN5wcdmTSaZQJl02a5FtT
3SDOsio/VCI+8E/ftEvCd+AcF4x0wjbzF8KBlTDTsed0c4BEG+WeXxQA3shnuiRE
0YcrsutGmUBp1ZKkQ+tnbhIOtBpKp/tOr3pP0qv8qxYY+GpvdHr43+xjhqv7LycD
JkMRZ9PhH2oeXAK4JgySy24xFD4NUKZm6pxGP+5ls8fnvL//k+OAxNLHVbmkNnz8
wcnSeAEgqQcGEcn9hvyRVJC/xhkH6okdz5aF6bGwdzUqymU5rME1aBNzhXBWgIpx
HMFmsr5hyit9IGF+Bl5qJZ+uPMwNI1bZuhzgQ/VM/fO55vyNEACT3w/SygnN6uGJ
xvK7QWbQnvt8hmLeXhFUS9U1TVKzxkEprEmM/TGS/aPpxNOfqdoqbfM3nYSGN7D+
jHaVXW/YZiQ0BoS6fBqeZ5/c+gdg0YGjUzJAOot2xYmfeE3Iq1dW/68D2v96Z0B2
sD6is09XSuFC5WXffi2CpkvLI18TYlpHYOHaTVN39ughmgVVzAhNZcy0zvC683Zh
N3BcpWBHN9Z8MKKsr68ttVkQAHWcQ0DPal/gbQZSQ4g3q+xZe+0GiVC7QjyoWokH
PamW3vpxRnZerIwCKEhii9/WwZrYeihECBYKfXN34qbKwIuSe3ftkR143TwULTCY
fUU7I3REvbPpLHfUoCsvkAmnmxwGwLIzgCq2w/y5lC88phJQcvzy2h7P8OSEguts
wbeQt9OOrmMG1vPFCoXCa6+mytKtKm+8CANcBr9+8nFadSCQwSibaGL153tO4PdT
CU37hFJ2tAls/IMPmW4vkiS3+dhNYek1/vFzJbgB6o0AypIugSMEfu5ON9Za0sqB
SdvR5IJlQQzxGXscDmcjCNwS4IEj4DrTV+xDzEHzpPtjKgX4QY16nVwp3CqP/WSW
LYcjh6BQaqTLvpKuRLqKe9q3l3MHGIpbLt12JODHuZrLh/Okmu/Hw7KPcec9A75u
79qPcVfXrASYHPeEMfkGGAMp+337Ne3iVH+vfO4eC2W14cpWSWOvMCUDJL6fbSiq
dQWPG+qeft/KR+3DYL2pzsQjSTQ/GoX1g89QWQ3Hiv8vS2NYpPkeB6bhv//8Xy05
gHsbbKqSJQunMDupDMg+J9nNavTr6iQ4S+FEK4u5nBdSUVrq7MMoYS8phJvv1qiZ
C3VHpAYLLn5tM4qboML5u8BF5Ba/4+/imMuyeQfP/cqYT+dbq7s9NNockZQ3R55g
P7ag+X72Yf9vWeApYNPmlhXwDtE4vFc9/iCjs6ESqVd9frViJ622+yzsNAGJ7uRp
uE64aBG3p4Mcrh3Osd/fh+ufUV1ZPorABPgF/g2CpWr9pHKy58zyTLfd5tODkW9x
80Yx7I/nhD/1RTe1BBGdLcRmAgBAleix6eVhkhn8QeD1PNABW2a5uSOnzRKX7jlR
jLomZEZOMUum737ykT0nJMIi0TJVH6KmRMGxKpn4DJWzNgNHvXHWZvfaIJqZiB2z
2pdlyRC/1W2MxkjNXUjIXM2tI6NHY6t1DPaMyN/vYt7wE3yXeBs5rJ6P4WttPY4X
qnM+ogCuVrNFPH/F/I82IFqykpW+VqQso+9DUDGORYh4goKS19s5cpIt+y86o2Lg
PytvXAdRhpvC6M7qSfryw8y/q3BS7OSYwnvaMbK8+kt1pSxW27bz/DehOPIs1Pvz
vb0LHSLcsf5zqabX92F37wAbNWWwFR0/MSAn/Bpu1QzhN5N03OQH2EDvqRG8RlNo
9MpNQLKwvtnAwSX8huJ3FStLOPp4kmk7vPMmFZ3eW83Yz6euvQT3INUt8lGpo4+z
Ql4PiFrDELtigy+dyXBnfUibb+j4PrLSkT6z63gXN85zimdqKJQ1ruBXHsc0yFss
I5v06IncBS4kWZlxp4Kdw0o3yz5MU/aSyk+qarNqfqZivnvXueNCplU9ziMowPFt
uppyjP86xVSameX8rFH+AlfPNpWxQ/X+PKAUyRIknrm8Ia/omqRvn+DSLajtJYPH
XUxy1jyAOG8NR7Gjb5xNOkkxt8cMFzmBHzG9D5z+w8M947RvR2NACIpj7bqGDeb/
OIMAYiukTUQ4rLxCcxOonluc919TOJBjR9pwbuSjl/g5Ja/yzJb8lsBxtFl+BGXD
36DW1ThT/VyMMCxNnT41SOkQd/+meWXwbQMOiw9POgkyiepAIdMNJgbSFik+6F3l
LjkWPChO1tH80SLcy0IXNsWS4Gs7r95slArtsl7CGmj6dSUx8r+5FCU0VUkO5McM
nlEf2dOgY6Db/6F+4svp6p/zSBQI/zbIL9RydeKePS1nF7DAidrK3Fg8FlTyv6rC
3pU7UQiRxSyoW7my33UiMQW1zAnpO32g6nSgqCWZxzt9wKGtNvGKye7HdJa8+m2/
FzSRaSse6hyLKAkQ7tY8m0+7fKgdMNFXJgjg3ePLaMMyeEibnfxK8z/m4Me34BYa
zKJGBcogygXnha6Cp+4WTsYpR6uGghNuZz+09s2FkWuzqLaAvtSQcJNM2r4YdCM8
ENiq6hpIoRgAnJ1LYjEY9WjLN6fysgHT5CymIUU8WlFm2k6DZds3zbFp0ExQHzii
b3uo9Bytnz0ZrWOjsoSV6FNfLyH8bkLBJo1JKlCrrnFO1JUJClxQU2SS1hoH6j4k
uJluwCCgKpEy0F9sXjHP5jY7Keheevo89Ma9cshxd4PTk6aM3GKQt0sCw/418yy/
5tFBikT7jG7iZ8cEWVO1yywopYvumRUhOPkQAmDFqqnx1yoNRi09a4HWPrYiZAvZ
cSH1DJasoKjBDXgDZo7BYrPCUFGcKOrlwmGgeuvYbL0ImqyVOAbImjCjCy8B8kmm
tVLyuVQW/fJyamWTn8JeOw7thXCWYHnqKqVhBWSEbIyeICcwHXlRffoGEL6jbxLI
udflbQx6L3IJxKgzznRybnMN47j9+YR5U9qGtwD/hxjsJKP1G7BnWYu7Fp1PDmvq
gnBWQtw7f92u2L+7WOAEbkl9UzbDiB03H2/+MwF8pC6kxDTkSN14mPs9vQkz7GD0
fhSbQc/kssxC17ecpFkhGmQ8erh61oh0tgwX1qmZEyLB32pdDOiY7VJ4wCx8o321
Y5gGn1GVwCzEcfMX2cCd1W+UdNQJVwsL5XfDdecZVaDZjl+xdxVH/THvM91zBTu6
Yb1se9y4MM3C9/wESBR/lWxLq6vnRhzD8+utODkBSj7vxEjmBMY6RPz6aI4v4Y4M
MYyngfmMcUdR0J6loAhxXhow8iVKRVDm+2iiMCctVbVXUa5mqfGSf2APMqInWpjU
a+uwwMNGRVDuNRHFw+F0VpXqlFGziX9lEoXBtb526lbu4NgXGujBNG0zFgvY+jEw
AeYN80N2ZuBuDXtKtsz3hwtzKXvpPF07KEQD55k60wsdFPvqIIsd/fuNuKamBQp4
q8c/R1+guteqw/PvF/qys6eUumDuxbf2YuMJ/AE1/lqDERoRXukUTh0gQueAo4+5
l0zikVWv8E1kc4ncVnEPX2uacawANMgiowPV/yg6KmndosZghKkZ5PDIZ4aAFoIq
IqPod4ljcjNHEgzcmRuB+lVePyrjAU+odn6UFdqQGJw0++ZgHq+cEaWSv4sZvYpP
dQUvvCxk/HkNEnl3tSoU4JZP3uFRLzH2WYwSjFQz3xP6yTkH5spp8TqdrlqtFS04
cTt7ENmPQL33VTRd7FH/EiX9UW7JEXQJjEAxHwwBLP1YEGRCaGD9msOUxQkn/E/Q
Y4A9THjmRozsbR+lTeiaBebiIQsu6uvkbfnZOajqKyf8jwJQx7xKnzbx08PFCyn6
I6n8Zlbm5aFMPnq/99wEsN+AVXdjK3hkntuUv3sqf3E5hc7lG0AzzGBQAgYmktDy
tYkKTlMb18AxfEf0qqsuNXxiue9ANZ7B+Gh0P1TfDx56x4w6jYsxbxsvYUDCxOat
uitiReXfXCCmX6gYcMZ9+Ni1Q/8Wwpabkm9TnY5fvIT5oD5kXNWdmPmUc+L3UO1c
4xxRCLb25AhicsBogE/CGcim16IYf/QlMgvQ6fkddhxJcRrATwGNI4kkbCezcpEJ
XLVhmOwnMqYoG1LWOOTDVZ++rCJ3hw+sqQGmC8kvlTfpTz+O+CVtcpuU8sD9Cikx
LciI55ikYUywt5z3Jl4/yXql7c/cOgh5qnTa4N8f52Q90TLEs8Pwa27esNHvyakS
pXb6Fm5wnQMrxFWl2zKkBI0USdpNjIpllB9/PURbEtSFSX7PZpn0L0irikYlGTfO
RUrU4Y8oOFXgzdoqeoJ90qAfvx3zmyutC+q/JOw9ZVLUFpk9Hjhq5SnBOCla9bzp
CuQCn4dxUkClMSBTnYEAYi0zKz1ynDPxLHqDvIkE31mzBq3B56mHW8KcsicyUHjZ
bz6Ysr5WMcM0zhmxUZpel1sl4xwlGJx5wswbr+n63krnrDylD/Fnm2aLebXg/52T
K5qex86qHYcLjLfhb+sYBB06Jdsrx7Zv6IxSprS5SJporaUY/vRFyyMZXEFBL1iY
qbZX8Xxuy8/TnN+9CK9Ke2SfeWA0+uV2ZUVrAv19S5q4oLxIhEu5Nmig5CvkyN11
KMMnguzSzKA4eZcLiUzLOzsRwxloHQc0F4bJ2znueP8pmqwCu18YZParDV6cddaP
R35SE60HMQaBWPGDSPVAlbnwX5IO8oVKCpeZqaKVVFItGoYdgDltVHx6McUj8vWR
5uEK1zG+/SElc5z0DtS9GoCtA3I1bk0mEXs6IxnHu2hjF3to62rQ62X5BU72a0aG
85WZKL6LJOAeUJQUAz6Py/g2bP5uGrJmIEyTVBrrXQwKOTAdv2aZ7LQXM55nZ+8f
aYfG7I/hkPh7IBTC5aRJRoohZjclGgshd8pph+pYzhS7q5ijiiw7aWZcFN6ZChOj
Y9Ffg6rW+nQCnoT5ikokv7HPqAG7xNNZl+bpiG0LeAP8yqUsTs1CiNW/D0BKgHZC
z9bj9h8BbMAXaX3mMyZRfz1hMJxG9j/Ci3pqGCoUtcenZ8dUYtJVRuE2La3F59wo
Tj++RD1OYn6SPmlI526nKKJqvEmH1KkFonoPKQWi/8ElG7p34WiOCW8Zlnfu+kJY
d77j/PYeDYXa8id36Z9uGu2K7wXPQzKVI+qlCEk0Ct3Or+zF0wNJAgqOOzYsgbps
qd89G/79+H1sSO8TQeLiSnwBNc5PHZm+9Fz//wXUWw4tHmb63ayigjqWVhGDQvqj
HpHUHk61/I5zrWzOoHDQcZ1nsak7dQWr54PxojrCnLqIOqgkWRK5TumzuUpEZyJp
vAf7+5WtKttyyztuoQLUNBuU9uWUqs1yH+atbGXOzC/Zm8vg3IMvXxEIsKETDXVW
k9Y1Q22U8w3SjeK0YH1vOSAPjpGnyRF5Qa3z3RCJQ9cYDvPm1Z+O0cMAYR3NfJjD
SiyAXCHcZbIiiq4BDQJ8CVgTTUOs81wwoxQwr07+uNVjmtiNWCbtZJXvK16/ZOyf
gp2OinySR63gaEOzruOWGrE7+t2pHFfD/kPTI3Vfoy9DsdhFLROeuSoOS3a0FhBq
XKOJAhTy8MEsfDDZ00s7VhLnUAuGVRNym8R7hRXBdxk8LHPcBbwpbv1+kdmvlkZN
SjhtKbwOX//q30+lPK10Jo7MD5AiphuQGmF6ZmWnGbpqL4kY2aLvyK1NPMwq/GP6
+7XZFh62jKLWhtINVNz9BH7jlj+F+RqR+DTfwLAC1sQ1W0H/MnDoSLTWjdz1B/E+
cPm9G5l14GdYLfl3OEaOyVDja83ANjTHHRO1Qj83Np1d9Kfm6VGoCWpiMOqUjZSZ
qGMLH8UwrFjvG2QMJKClD9uLoUzfUSQZc5LaHJ6Dg58/Vr1xYWxHPMXqF7fqviSA
YqOkv2yHFntNU28Dg3I+ZLuHtZlf8HEpfUBWsloxY4lHpqmjoyPN4/P1364/I5lL
B48431uV6I+3xx1iugxjk5q8ED6t9QOfpyMOm4wYTLaAK76Rbd0l3NBkvrElXSeR
0Lw+zbOuk5Z34tg9xZ08q/B85mdIFmiCOgJTCKYOJoZe1sLz5lsEOyBsipgf1vxa
vbLMzngwHPFd6uf5NjVVCsHEQg41wEE5chE9q2vYrDbwAmjR0Qwvc+QX3x8VBKbS
V6hC5RkrV4vsEkKCp9ZCZQcGGe0NDxz1KsQecR4U4tK9Wl2WUMMTzZVtPoPGrOd8
0xTwvpe4twmPuZBz75wyS8DpatwNxw9Oxn7cXc7ati+0FqWb6FJf5iE3h4E6JTwB
VaKHOiHZxAn+8DBoWoUCwmLVtBh1w+r5tzd6rHTjxkhrAoBy0FQGs2iZp5f6/9IJ
9/gBLVw9FxE/m1QxOe3sOPPO9X2yEgVuD9Hq/DSNOyn5aIipzfTQfdiIcpBkAmOH
ILmKBHD4cgXJlcP7UPGMw9Bo47UfWiac5sfdHZy17DjUchmxuiedNZhico/zmh94
pPw2VL/FXT+YtC7VTWJcHBBuF82Xnup12o6JX1whADqXcrCKxwUhr431qhj7TcKH
FmtPgC0Ovv85KbrdKm9Ovng7NNMTy7VrpTII1zHLqUOzvYo8qnZGsudwYTOxHVtn
sxH/x+1xZvhK0IFHcRJ/eGMCrIxHPp0WGnLzhtOkJzB2QChBmSwgWIxUrIYL4AoV
Otfqk2H4676BP7hlWVsb/zdRxJK3/Q6o4vrFrEeKeaEVpI+D9zJazANVvgrsVhvC
8bsYY8Jiia0Z+HvWgFmcCZgx/1x5qcorh/o6DLvRriZJGE3bhaD3RnNL5+YrY2JD
MCsqTCh4KowSysl1HtJkAIVmAEjMObhrIcz1ga5N3q3wHodOWgwUsASjiMxqOZvd
NLk8pNcaDsPut5abBZ6tSP8yZnQe4He2jQWs9hi2Y5rbVqc44849bk1n4mA+siBH
az1t0aJoh19y7EGEDhfcVg/eBynrAJ8MeCifVKWAMOLYAsJ9LO9zfaL55Ir5hJIH
r4tnynnA4z9clb4YRj4xtUy59WqXNlC/6NZJL37WgfHnxdsgZPrTSww4cimBvWe4
2297Xbg7zM7I7ZqMvacApB92OW3v7n188y/Q60t+L5lpJtsfkIqpqq+uMzqCfv4O
OB0G2PfOiEg4jebKdr99rjlxNbPgnqhzzN24ZP+YB5wqdBI8ZBQGyEBOh7+8ugxN
oeIaR85GSRIDLyL0AGVFnMvRNabZr9PIX/PrOqWQgNtglY7mBcKi42cXgq6vh5TI
5HDWqo/D32uUlN7f/801Cd1ZaFx+5TLfFeyB9O3TI/og6apPTh5uidFqKZMRIKL0
0HnEwixTkHYn2Ogg5DP7h7zQAjq7vCLPLxM6S1+u88ZGzQzyDPzL02jazvG+Nq6A
f9KNErqM46wIkjT/W70i/qOxylHJQ4naLtSQJ/frH7NrGPQiQKuXemHmHaMIsZYc
dd4qMJYcvZxNATrRbhlrZgqCh79/ezfgOQo8li3Tmdvg0rhPqbvYCkxKSNd/Cw/o
tESyLm2UlxZqcvKRghR7G3vQwmBnf7Gzou5yIN4hSWbWqJDrYc2u9hNI2z+NUJwJ
dPzDtmd9LQvQqERuDPTuLATrlh3TYxgMbZ1U4Gv0p3i9EHx7rqOjdJn9P5fPyqTQ
2EP+G26tlsjBkDpiRnyULm5LZ8SXadXoubJ+LtUsYVjRtsPL8WnY7prkU3zmzCY6
f078JM4Kw3A63ezptbwGy4K5pe8EqyX827FdGKYItQ0g850+rGG37ijZgfXeXdqK
jf58lo7LTVtwKIEyt6XLf/hVI+h4wUg3LyfoUNMIfzmloWPBeHm0aaV7t0roKtUy
2ZgMgwpiitJ8fILNCyVNubvrdURNT6yA8TdwNyjdoCzL07G9UxCIRn6kf/X6TI2I
1VqyR+Ki9vl7gNcBZwK/Tefak5zg5VnDoW5ZuW6ar9SP8xXCbLl0YuVDmYGN/Taf
wPVhkifgtfroKEbHJSl4GhErtkSOQQoOUaSxUV7LQyLMTmbWVKs7St1UmVsEHGQo
BJkMxINXTKENmmaGJBMLtqZMLaQWUNRDuC55utfOajsZOBmwOnxRmBO5t4hro8Io
IDL0JYX9pOX4CrmMwKgFZh4WGMex+VOat9yHu3+K3eXCLoJAFFWZcI4wBK4U3OsB
kNtNxLAFzfELmQk2FyL5iLwk86daaX0IOuwLo1FxP8kDt01vNN87PXXn0tdSq3Fr
vn5C0qZTHNDgmMklB2mW2ekTzvMy+9T6TSw96VQ/ONnmToufXyZbjymYu+IX2vpD
OTuUMA0jisOd81EA7Vim+BveaDhAy5NN+qIj579Ckvl0hodOzUR2Jv4VwhlUZiNS
lSset83B2Hjpmim2oZ9oOqF118ckQukbtPA+c2q8DlxMTUC0eiJuuigQqutbi0N4
2PYoTvj45cKxsQRna0aAqJk19zmdGfG3XfJo5Jz52eoPw5RWeqG5w5Z+DUVz6yHB
dEeCtzYsSgVqYEg5T2h3QMqw7hk2YbpwcdkeufaAUkaY/dycGXNv0bpir8qTdAAb
MdbaD3fz7dh5qXeF2Rz1jYhWQyM7Yfuj3BDLTEDC/wXTglEKLux0QiHavh9nMAVD
uD+e15EE9SlY8ihFdHMjnUIGbc94Zh67D+H9O+eieUJ+lX0vyX6h418lWSI5d9OA
p2glLS21sXEP1a4kjD9o9zQ6JE4yRN0M41rr6XRljlbyHaDxu6XI7pPGi2KyWGph
FmWpRS013zF51cXtK99grxLL9p9mE+6mb2BByqcVZvzaRtvGtkvTh1vItXDyq+0W
bJnOQZYM4CauerZqdWi9cFPbF53VtKGnXYhxaGTOtp+kbBQQlqD560T/sQUBN2EI
0y0JTry9M250vTZMLQHVynUF6M1+tqn41zpHGMXCA9aM23WsjdwMk352QjKg9Dy6
dem3cpYkR4341dDtPrKyibfZ+RzRtkwwF9GrNdL8vEjkiNPNNUeKIov8f5nGSqzo
6PLq/W7V18glfpChujuYPCk4lMbsBFLj5WjyQms+ZffNxq42VN4Urpko+E1zR+hU
EUUZzfskJrDGjl8dkLYJzSnlkccFSZYjLoChaFEMBa3uY8Grb4/BEP7HDK62829w
M3edHZVhzY5zjEaVrZ+/8R0QCfLBlihzZaRtcwdxR2rg45QJGyykmk4ei6ovfAFG
FjP3+WJ5SPIGqXdiSvqoUhP5NihJDaQoMQq0MDGGi2QA8PpGXdZdOPrHg904Kg8K
BTKkmvWUUsMSvkF071PvasFCBAoWupo7umIhqMNqJOxznzlfLuZRqiXDGBmSEZtd
mER1Nii+DokfM3cIZRgulQ84Q6nu8vsumeE8PlAoolQCk6JhdfxrneT8B+KcYfCY
CxJ7Z1G+uTDFFRmRrBHYettyK9vuwxIoTO6JyuKk2s3iNBjh2NJsRgZy8r06Zf2I
EC0yIhUPAMI4fa+dP7bGDjm1PntxpmQ7lufM8qigr6QoJm0m0XIifZcyBufwsiiK
za3ZpTwd4j3bqYhEDmnQ4tgT12fDwOgEefxuA2fVoXI5PRLht6EUBs9ABFsmJ7kn
ooy+EBPBbkKgK+OzyS2T58r+O9eVUpMNCf020r8l+xRt82WwRUr/zsZLNczvXAn9
G3wBCiZ5ykIaULAv1opzk59MnigUNJfYEEBHtpeGXP4R9RFJf76ygjzp35CI/1/i
DUivTHxo4D1R0RA6mhorlNYB+MiM/aS7siMQvU+2kZmb7roxBZVlrAfirpKR9CY9
1KGFVwTYdGKhzvF4NN2CbSBdFfO4e9sf+aFA4mORFMgaUW6AkTPIB437IlMffgpr
E3w2tyvTrJkdkF5BL5eKXeU/NAmUb3TRXsZREMW+H3Q/ucmjl3fHk9hw4K1K9/dS
oi7Yb/JZB4PQxU/tMmA8X7xa3NQFSUloTlbyNOckFvuLiJXmosGMssoXtttOzxEB
lYuce8w+l3ngZKFkfNlVUw1l4IB+vEACDOEI7yu5hb77qd2q8qbOH6jNRzVEx9WH
4G8gHSKf5y/BrkDjy/ARkUBYeHw48Aj5eacotAHfw1fkmiCua0XyZ4XbOp6lVLQf
fuBjeR1f0VcAfDfMLCRHeo+Fur7D+NN1rmHnVqASRUs9VbWgoPSpWMbstDcpME8e
6WdOc/HIgRiQV7oARScO1EcK71CYFPjuxqb89G68m2PtxtUc0Rissaoft2A2HmER
NvfoA5ivH3xCJ0vYFyrrB6W9y2HQu3x0QO2KFeF5FxH0qvLpLOjkA/0HsNEc7UeE
L/KdGAJPj9DAu4ofXNmdp5le/qCN10yG0d1xh2rspYQBngQMGmnXWJY6GzT1HwPv
qtGQy8wNePCmm8P2vZBbJkgBHf3GaUaywZcdHu8WOJdOJ88kxWlKK9pEKfiSIiKB
nliXvQXrBpJfI5F/96+D6LlOlrrL8u+BBL57U9nMGjjQEiU1uGQ61Fe5o5Wfyzcb
5gFt1iJCJyXgasJ8Au4HsgXEp/kapIR2pYzDf/5Riaav7a9jSLS19sYw0KXRWw+v
L9Q9FARCL823cuD1zqVNZt6vL4OqsRjVJ4c1K/mHYqEJhtnuz15URfzHn8YmK4lA
oC1DkEwWtkwfNEbD+MKud35EMwayHzRd8zMXk25eb3Ayd1ZMFgsMl46iXr3Th8Ci
3OlT4SyhIBaVgWNjaNfTOodI6npJFxwnTX8hmfkXrrdZ0S2xUDgnpEbVsTcfNbMK
E5N335YykTUXxsiij6E1qyFU+AmEddHV9k+OU/rooshgDQEstJwjIbnFAK8Kn7Fj
wuc8xdLaGr4w8nJFqJQJpwnbzK5+SptvcZCJbKvhJhpbBAqAn+Qew5wh+R03NXUM
4sMKSD+F0Ekujv9+QrL0HVn+J3yRK7J3EPPOACw67etZSk3b3R1SESRC0p9VU+IT
pgovUMNbrQqCHv1Fo/5D+W05iJT1Re9pfPj1Gnm07hKOCFJ6clqXQlXsMUDw7ClG
4dfj8JRaFNShTcngJkVCW55wAM6ac8pS8Y1eue9YkgalRxdmoa/7Jfl+kI9qd5QO
M4rJN+1Xq0UY4b59G8AMZ5CYVmkfzVzeslGMNBcxe5Ccl4smvrFaP6MEGOsvCj3p
RPnhOwDlWc6fWG8qiqvf+Zpqc5ZSS/h3F4/WNcNn+YWESQ+4sdOcLaf6wRF5PKta
xndCh3xxfGNCjD9XFUgRQhfaj8ZF2rlnohI5xoiV6R/jehxMntG3pSdIXPbxSlV1
zr8EyhBDArrPPMBZEKH1JaJHFX6uSRoGrVuqKe42yq5oXvsMJTOYgcEaXVa+J2OG
iS7tsttFjEbxzCuq0Cl0L9msJJ+I4vArH0z2dGJ4u/EBG3h6TYaTDdCO7rmfGrDv
zRqqow/02+b+LrIAwgoDqCuW1LuK3agMSMKoILC7TwWU1N01rhPxitO5HRQOGNvE
ThpvOqVuHgRrHX4OEGWDyDyWbcB2wqOtU0/prW5ItCwu9hkcPh2bfXB+MJYkqZ0+
3MMghGXp0kbQG7Z86SsxmYmK0kQMmAN7XAVpxheQxHdESEVizfRN2POsAzHSVZ42
tPU0KwuhOZOVwvZUa7jPwgVo60jXHWGOHO6y4syyZfDF1xC2x88LNNk7PbKK++pA
avDpDUvysp75wwAZXdHGoAkQjUTVhh/+2RG1bUH+P8Fz27A41k4BpjlYCTA/jWEB
KewovKzSMiJ5ZPmZYh7cGkAPYope1j/ROvjwzcV4uBXqB4Jry0OgEEw70oZz1eAs
KMRKs/gWNQXawsy7vh5fVHPGrPqymOdrNo9CEgBSaYhy1BPbWnh1Hp46NooGj0Ss
le1KB6APR7O434p5fQs71lSOWDFhLbSieS3Ya0cPxZBAZw4taKl6yjxEbKoeC7C2
nm98stetnb8d1s9/NyXvTX3H14iVNIln2HBqRy7Drd4erUUuRWc0G75gPrGLGZDR
4BTCoDpikfFhHb+LYcmq/22KDt6ITOcOGtu2yjwe/+iNNtI/B6sf6DNzJa7muY75
1JDcPtkIh5hH+ujRp5NFgOarKUwMsOUIdmUBTzGmSVBzwqn6lqwzgDlf+YaB53eN
7r/8+NORgRwUahxNNYmxFDAwo8LPPk5qTUxdWnxtYIPmaSdxqk/TtBR942mPFSZi
HYH+GKSjRm2QHLW+WSz5PsRXibMJ0JUhFtbNuIfYzTJvAtqgtN8XiD6HjFmehw/i
0CvXdqKGvUXFX+NxF4u+s0kn5ujA8joAcO8QeuWMZwibPTnibUpimEXdwffzAUGk
ToYjF5WCblM01kSD9FUrYFhMEHu5LXZEWoldaLuFXRVpgdjCu34tyNnpekNuNZNI
Zy69/CZKTxlLS56C0fHAuupow72h4RjgAs66WWLVlW2+IfOvhbjegZoS1kCOkHQG
ANPzF3GtDHDkR8NsHUeBMA4HVihDT56gDLTTHwNUItDxY5vbRRWtH/Hr4a4iYQfh
tboylesN8UVXmonO1PR/0UCpt499UMXistEk3ioYiMsI1fc6A8BgVPUyHoU0FVs0
OG0AGp/rLfp6soYkpBHgdjvt5x3RmYn9OnEfIvfE1bkrja54XJbrbjUlMGSGh/Ox
uUCp4CpPz9sAOhnj4THUU61uQTCabRmrHvNy4DU/sdAhyHvZVzvIYgmgYZKpOArq
jxBHkbRYW5vQUxuc4fj/ZQXbrixnMY1xKdyrnAcnBMstUYkpGBrOgvfDJ7WfiAZ9
byfcSU43pi8yZU8geTnC0+Z6aMxaT5lKEqlilfHDl+M5ioQzigtBse8AMAA8bmaA
h7RIGTxYQSowvDFC9AXMGVhrBOaFrUwnEUFBatQ1gG49iO7Euid0Enzfgjcun/4+
B/gzyxQxIysfzcU/Ve2ELLnGDXJbksRD7e44p/Kc7xBi27cswI+ldEVtp/sofD7Y
w8Oe+ioyt65LyqYo0P61w1gx5N1Hi0bds2lMDck12zB1ehH7dG5iaf4dbow97/Dw
jHOyN6F/Rz6UkhAS0u8OLY7vRbxTMeiFAPmLwpcuy5HYjUbvtTnhMb0x1ISDh8Kp
5DQXvkZcWDuQtokcKwxs4EgDv/bP4E1YaaYqfUqt1aug3cP+4SKwB1nJvPmZFOMk
cI0weX967jTjk8JSzkrziUvvP2BiiNZmNm8lNGz7qrAGF+L6pv92lgx3Tb6+QL6F
Pt/vYzLmBH7NyclmfUbnjoASBOUwj8VE/N33l2Ym+u/k1JYLLE0PdKJWZvXYwVs4
AYZLel8hSjNJddbr3idR6OsCcKTs7W6IS6DG+u816WFYSdylnEoLR0AItRPxbKeR
gHThKghHMDDy3KOlMFyD/fLYe+uWAoeJoEVqjvaPAOmxXCmJAFNIyoJzW6Vo8TTt
FvGqOtz2L+UXWwQTUF9BDJM7IQmg4VK2Y3fcJ+rRAQjv0Vwj3ZwelQ+x9ommIOyg
KW7SpASQ3yDHPUuvN8bRWASKdnqjsL//OZ+W7Sfa1Zkk3dWogcz+LlnWds7lBRs+
vEsu/LkzMj4mupDLY6Rfc82cWkyK/EssSICtKJn+5lk2ghmg+Xsr3sB/VppXeNzD
ywcOJHwqDzfMo0KHI/WsGIh1W2pccVzT2WFRVNRi5R3XtZEDVgokcMfwnXJFkKqS
dromifOVHyrZQTMjMnWBbrQ4lKwuE/hs/79/NApBChEcP9YS2/Ne5VKGH5hoImok
1z5sl8jQDyuCqd6E+PEyXAxb6tT8jbihWZjnQUyoA7doyGNOzllyztX8AT10btWi
iBD+1h2XFrvNr6Ehj05zWIolROEMLVLznqA1//rCS3r+T/xIougpznM1QRB8euR9
tbYlTGxMEWIpYdNBAwwWdF9HXDUz0gLhBcBxNjrBmQFityHSygBHAqVwVgkrSFYr
WK0cCVQqT6b4VHYk5/x8NSLgkLtCmKPF+tjrk0zS5okvezQYhle+lp7d1UcPtJqo
E+fJ8kUCKepIKhWBm8POdZI7iSHwd+4yq0Ghv2xiO22MbU5bowuYzEGIFeB38Sn7
LGYJm5tl2iNMx0x+8zx03ryPg6oIHmXHiyIkVZrgwQkH2eFDbNvgGJlLpILdFp5l
9y+HeJ/aNKhPsh6lQZ4QURzQI2IYZAHu2AiTaZnVHEu9SWQd5rnPipHHU+ReQvuE
cubHCcU2jOXo4Dis8kL/5NrfG+/fc69RVgcExC7/MvzQxSVcIuHOBYFhEp75ahVC
DjLX2jA/QTjCJvjv0ljzHpAGBdPfOZiVGXd1nV2oodfZpqpO7oK0tZwVTi752t/g
H1WM5zzMDv0+xnJV4kMnCaIcGdfsBcflS13PRrMtfxlPwmzpkCdLTmhOsEha12h4
NZrrOzSzFftoES2aG56vXZcYnm3DtkHv7NGS260C/ZKWJPpD03EUIglHbBt1yoKS
OhBTiRk8z0yd+AVsBfpIn301QlGF7ycXxl3CD8yC+b5laZxVURrU4rZA//EXeQj3
HsJCeA9H9bDFXI0yYeUm/9KAdMqa8pY4r1siqPKIVoaTnac2BlKZqrEUkjzhh6kQ
kffGilWmW0Qfsz+mppCgMOtcvKIV+V37UFPn8PigmalrTuoTT+JL+uwuZPt9isS5
NegnSj00iElHAxVqHkggtBQZ5YtiO9xSBJ6I3gSiw7ha3INfm+qtQHUAR9WqYfu/
XZwTx8zV065RLD7irgmUTXxzFtsVDdOtHrnL/LL3JKoNMGhpfC1RytIncDQ+dLie
bS9YSFbz5dKOjRIwWEPnNtAIym3T9ssPcUkmmG0w+wZg5A+PYOFqrdQSQw+RYNzQ
kRCGkEmySjdk6g6tsCoaOM6CEBGt+Bv9uf7l0fWyFdfkVmsV8TRmn66nEnQoHpX0
HFeh4se39p75u7uHQneEo0NU4wJ1BFV38JOfqlpx9mb3GCDLGxq8dzmCs3JtoWCX
3zRNYjtboA29Z20oGgJtTfQRMeBda4BD9Kzp5cMHggIkf0ZYTWUFunwGHa6C6YMP
OGcyTRScHZ8rl7A7l1Cu9OSko04L+GuSFQ2DdU7jlYwEjKdiRhnaR76PB4eRh1sv
Znihk5Vi7LPUfeB6UtZKozSo1g7Y9tZ9/Gz7WLsfV9Cv4fjhzLO4eDNliFUaaJU1
vdG6obmB6sSqnMMxAjkty/qydCXQRaVvy4yaL7soNSMCxindEg/dxvi624rlsICW
nuFL17k06I+LbogvcC5EaY+dCZBtyAJ1isr8vwAZV2Xg/sEKF66LVHsheDmKnWhP
96MZoBpRM7YeOKE1Pzd6a1ym9ZBiYP+py8CoFg+X1NGM9G9sXKsqyX921snYwK6J
/buHTqrQiQhCQYzRNUNRszpbA3JNhzPpojs1h9QzHbzSoN9C/G/u7D7axRMSFXQ1
cXSuOMzQFbEv65aY4I26uR3zU5bkD7Kw8uDXiktO7vNWGgOYGdhIrokmvTQmpEn2
XQ8YvfgBS7OisyNWw+dhfKTzpmeA6AVRkR4cOzKD+krzTPXNgZi4ceseZZlJ8p6Z
99FBAKE8R1D/yWOVgw0m4p7sFO2Se2JfY5GppE99QWvQyvbYc/5LjnO5pRCVP4xa
ILJ612RWH/IWJWr8kPSfI8FQ/drQIwCrOVOTQ64NgqR25Gb1RPgyz05aCsYG96FW
zojIWbC5Ll5OjGM+suA3Kke4kYT1VWcsT16/qxxsg25EPB7aU+uJZayEcgzCteKY
MwPiHmLnqsIjZNvSHE4nw1sDwLpEaqfK+dIneLPucARg0GX9k/AehC8Krvm/e/eV
Ck9ree+V8kJs8M2R3m2E2ZUfFmejueFUOV2Vr9LSyXxa+CLwFT2yZq57U+1AkxAX
bCl5WEUe1j6hBm/XGo5+7yB9Ib+O1Noz/QnmTSj91jZx7vLW2Yi/wFUxDmv5fF4t
5fFdCEM98NWZuvrme+mN62CPEXdj3ZgBaKZw2yEzFZE+Apa4DagDBJ2etOvYKX05
eQfyrWytLrff9EMsFE9wopENInRzgw7gZ9Si/ApEvmfWeqNI2VlJJy0XTk0a3jij
eCn7qX5DwGrZiRnIcxUCAwLvHIVNRwNh+bjrh3aaGXSteAEGOCz/r0swmeNvE+LT
AYiT/XSTs8oRdrtW0HHopzwq03NxzBUq2ePlL+jsvhFey0ERqM5L0We+8hQ+fXcn
YxZIQ4MHwWo3ZtzUduqzNV1dPFQMYQTp+yhFoevIGRCPvJkuWX9bfqj8aGrmHWVN
2Vi2+20YgXfbreXIZShKNz7RvtZnO6uEv5QGGjnAGx2pLAfrYxjImgCDwIMxEKtb
yh+PnG4A37HwDgL0RhBBsfLU8R744w+bFgtwPIR2ymgxWE5Kd6LDww9Qzt0mJ0Iy
Xghm0DMXJTVWDZenoY421pLG6Y+nSHGYrdueuBci+njOzaeAkQsUnQ8nWMidgo6w
U4IOvZJXs6wYfK2FkrX5/WAP2k7PGZfT/X5Cvemlm8+ozn673mQHvyzOvCabwO4y
8QiiGWfUKJUPPWFMjbRYC1hw6y0xg4p6LxKfX0Rr/hystBIPqjjVZvHdVwlxXEwp
FCIrED1crWD+7ydeAflGoRm0HRiOVxrZcgpPLkg2ZYt1FsBPKsPjcz7Rsidr2Oy9
7OTzlartddMBgG6NJXcITkyYbTU9eO6Uw8zHbQ4xTvoIWs9Uf57+jJYHqlPp9q83
e3UyfcCmmcWtGbhLyDndEYhyXc6akx/JH+wveChmB/oamTzzd1SCp+StffpRMv5y
afHHdYP7PfjkDQ9LFV5shLLI41tDRbWeYmJ+j2zbvfXlozWGYE5cp1KYSHlKugmi
rpOqiK1HhrcMqRsGwZ8U5kcmcPK3UFRMixg88x+i7oPotwO1Q4xTjEipwfac7iiR
Icpufzhm86DFDJKloTeC2et094CUF4RnNTsKhqWgcepjBGz5Q3vM/zFSDd+uB6B+
ysih/dS9GGxpaXWutTEuwQ3IhO8Rckq1AfHYmPF5ft/J1qAAkuBKofzhaFxTdNCn
PPm3jt//5RWAsB/yYmdfncdrVZYwODJZzuqYz4aO2eC4mwY6PkzQNAhH1vhCSdPV
w7g/zdwnr8neSCpVLYoCSSI7NTQJz2NY//mHrFsolPjFN2eF5LXX/upr8t/IZnh0
/wMyXJsEym6+ybqx9Lo4vAwZkrNdi0mvw3F+F235b/QuGW4+Cg1a6azP1q0r5z8c
vW8xoWgTs6lrxRdvOAYFZ6NsX7xdH1Jqqws2JrgDVgOLTdzLHuY65t+N9dgOwQu+
RZ7JIo8ZBLtDrunIoNp6DqsOQkeYeWv3mu03WO/nlbzwe/g8o3BEh/jKoxoqItbD
0op3O0FfKsVN87bvJ85+vIJ5KMJg2tn++DEWzp0yONV5rD0HCOdtk00/S0VUiU0X
DQ04Ab2MLKWR20aFdUdaqlRs6zEk4Ib8VK7PVvrYSKuQav8MmcfYKfkxESmsKVUB
0CBMt0fZQesZBkoFNMgW0DyIwq7fRzzc03Y0JBOsB6V7SN+pFCzxvafPJla6F+Qz
PpZ9QFlwqVLbKTGtY0waTcbb4e80OiHSvw1lCzkhyskfAKwN7Vbkg+87vznR5ICj
hSuSl8OuMXVZBVGMFQ5iRZmRoy7Vlt/nUfGWiA0QQbecgHe3Q/haZ9kG80O5Cc0y
25sX7KMP/yF8PhZ0TQJArxeHZKgshACALj/Pyh8Q6EXX5gjZwg4TdHE2KOntwnYX
iPizokPS4kL6yR9Flyj+BWBDsNugiWt+qPJoVRVTGIoxkr96GoeEtnWc3bbKZE6f
wz+zd8lYDDXmw37VzTjTn5cBItHJZOCLPsVGcmJURfLD6MP5mOXUwEl6QVpqeL16
aHDp5yidizaOC3MvPlRE+LAhwCG/QZ9ZGuaT46j9V7Rh0QEqC7V/y+YJC2RnXk4d
iypqn2CMfXxW1DLi/xdL08/hLWHQEKTdpxQHrcpBZqe9XOaydDk/dIKXU8Ce8tqb
o5mI9d67rINb2q0iO9zWTrvwUnP04dhfEapKyOR27Xt1AX8JW4oyzcKiD3bPXW12
g0BQtmpNktmFaqD1vYO5rtZUwAqjwTHMD9V65HskaFyweMjq7HvMP6hA/7w0ZCW/
8gZPzbsBOgTVUuglQuJ+7L65PaYeQ1LssIWxACyZEOdv3iXHUMWMYgX50NKO35CT
auQXqTNF04oE9bQIFD/vxXVtwzFjuqheSDx9ydalbDVHtq+Rx/NVO6HNCQ/NYy4D
34+HvCvFOcYJ3lLE/khKuskeXlrJYI6uoqJbO1lOS3Lb0ibTze8CKO+GlUSVK/dj
XMvuSDB9Uq0vVhLGY+nx3tVqntBO13/PN59sCYNocXH3uWn8P3pUHtrL19GYSlJn
YljXNLre2VG0om7JCD/FcXBmIZHl5qRm9ZKNmnmFKaERUr1QI9SX6SVCe94Uvcon
nHuhu7QibRy7dYBc56dNxlDuyk4yX7vCug2Uy2NywhSMuLlPOxQhP6Bk1BADVXQO
i+xXTNGDNRbjbGAkNWQ95NJR457qiW6ld7jR7mB1C4OTzwd7M5vDNxq9jnyTOcvj
+zLFGA1F7j2bsQK9gmACU6e4ZAw1xW43rr/huRqa9Fq8MHOR6tMnjyhSVbtQNZw1
kTMUROXfEYCuuTs3U5ULV40nfG5sdXL0bkH3vyE3lTehSpNa3wT0gedZb6ZOs/zu
EhP78mUOKKKLberz8kaTS/Mkzx5bgJLdVYBoxzIWDgjwUZFZCNOfoYyBu0WysbYb
waftCEUmFaH5Iqh5kMOA74M+IoXwUkDuu2yETSpLFN0aUAYnbUhTrsGYBhv3q515
muJM0TfsIl282VNJYWN5jFprFI6Tg33t4aY52LEejUQQVCewbBsE/vRa1fh97ia3
kQUgoZgUwhvUEJuPFH92Xai9jPeNUthnEehTGRCXyoCOW3Izi4UJCa6PAiXxq98c
pzRV2yQ3i0Px3/YO5rlZ24P18QfVzfh/ztXQfWZ7dazXxW48/2eTAFV0shy1qQuH
IIwPGpBORX7LCmWuxR6GWFEWfL66ZDBKKO6X/RKzUaiS9knCupFbYFy56IcLtX5K
29WN6txltjDG7cITWrfhCDnRaUJLYNkAwZ/6OMAwyDAytj/wKZLT+LXQ46LYlSx7
NQgU8ODPkKPxk9RjXrI1NvJFIIYc+TFYDUy2PbeSE2Hm1O+vbWcgaO3+XAmFaffA
dygmnTv5keX2oBxLZwLIfWqeBpLv9+xH3bP+uWCwYaeZM1ja/Xw0Os6E7jUhbX3a
fOs84MEg2jJUuETXVnzqDRwpO56+riqNKpujV3H3aAwUzG080PeWOMr6ASPe2woW
+uGRJfRe6wYR7UsqhhpoC1p6qiqE0C6JDmjw8GQmPVZYo7WGXjk8DDDAGCDcLRh6
fMnF2NLHPRWNQbHw8HL1FHIWLGJuXFgQNZgSwlT+u47ivQJKPlSSHrFAXwejiG4Q
TllLHuonKer2Owt6KbCkkGkOvmJGbSXiLwIIlbgXSKzXtdU6/qlEbjzPwAyIXjrD
eSioQVjrskMwcan1oAjDWlTkdVQPRYYe9iaDPjrR1o7GX685mBFdDON13YPdtzfi
0qLuGcPGx2YSymzXo2+EsSz2rxj5MKmxu3eBt+adUsGHRiXv44L7Wsnj6m6hDu2/
h8WeGruroFn14Q0+HG3Un9yP7TnuBl9l5Xw6009mYhQoxLOpxizNiuMWA32kLYY6
NlGkoY1dGT+zwOPMoZ1B6MomUxoKzocHcYC0p8cKl3LEF5NfCMUOv24C4S7wqaXh
mWqXq+XBDoNhHkhmXYr+RhgnVePGMa5VJu217lQA8YdWfIox6FpAsxalyPMORtyd
75pSNxMeVaxiUmrnANLjjVTSVQeyie5vmpog9cOaNkkOCE2++17BNXtQ3s8/GyWg
TRxRIFKkOoo4snth3fIKi1Gv60F5BTKiEzP5xhUoBVUZqNLQy7wG/UE36k+vDI60
WgK0FWkbPnmBvwnYo0Jg3kWFI3r+uTUIPcLM5ORpkGY1dvi2IbcWIsqPiAtc9NB/
JThR6hzzooT39FDpu2Rlgv1EVMugWyE6JVWsnEHHVcmzsfoWaTP9AyVm48/Z9KDI
Od56hm5vAO+PKg244w9HSSE1DW9sQ7CBQ9E6311STArDxUtIkzSmgdWfp/wzwsfT
VwyLvTra2IYJ4Vr4/9mPcOZoF+2FxffKV88Q+3jMTdoEFjhmeDMx4oWja0oF6jS/
r1CUW4sJ5Pk2g1RcNTLZbqlthEsXCuBiJyiMmTHBpmgMSFOj9mutylB/vTZp4m+O
aQMB71Y7mhfQU7olD/QPZN92PH71KpzM71H9yevfE3G7DeGycBAYxrtfCnvXk7r+
eV9suxgzk8/oHbzmQjp054ZAMVOiy+zsPW9SsMoxWz5tJCX9NgnOcrxV9CeEVkLK
fjOKJg1iNOw0XZD8iIv5wl+V+5T5n1AX/ejPVi6RcW6mbg+LhIJLuzLWTrMhLltA
gTjuqY7/EwO+UT8g5qmNreTSPvU92yM2gppUfp2yvYdDHOjk6MX2TDzohZX14Khd
+uBMbpgdtzAcqslacU/QDDIZkynS5iYG7NOWkDP871nU5pfw1SS+9NMo+dPUFYL5
1tu+Nn3KZcdrffVR5+AbuaVkW/hEcEYMSvGBATVbNWNZ9kOWLTlfHXK3Pb1h8kKd
JxWbLCYna7UqV7WDPs+rI2RuCKeAnPRt8weY3b87ZgKUFRcmcD/ITyV4HoOn5Owz
AliMZix6s0hXja4V3YGw4grvUd55BM+MA5V2/wOX2KuBeEQwk6i8BR1wVz6P9ukO
cGsYlWutMOM+CEpDXbn4WCSYBtSmXMRp+7XH1R94iix/lnErzo6KkSMj7JR30Y2e
w+/ATYcnzIbcIHvbdo5oobvua7a8H8yWsFeqD5tTq9S25U+S/Cs5ENJ7fHIgR7e7
FNEigwNeAJb7JyuA4I23Hrkv9MM2DW3MfZQLqaxBx1ZJhcznDTzcv0afiv1jg8G+
cE/mHE4n5N2U8sUiaR1AuwFLM1vG4XoAEqbZVgLHgy0lv9vQW+7O9bFpnyEDcCOM
VVBkyjqNecKI1HcpTfni8/39GcGC/hPM8Di1HxiBLw6Z/VHr9ImV11xHYkLPWSyz
xF1hqcjg/IG1OwcNvjBgVbduD3U9MW6KEXy5sCtoAfMCW/O3H4qrfiInaSeIIJZM
mH92GoXoECBTWEv9aQguT/CshAWjurWfYbXODxKhEpEIJs3QxyROvbBB4UobPt3/
oUolsP9ZUKrxd5ACAHLidABq//qpP0DrDLj4Y62EeZgH5UDurvcYY9OhqKRvXv/t
PKhJ5j+su6rcpVLy9rNwO57GF1g1dubHLbz2C14nzi/km+XPS4YTt67xgPJTmUSK
VsZDJr16QzOGRE7AOCl0v15bSw/DNBpqQKLtQDb0ZIDuenEZMTzpUr8LTnWhfmq6
K9uYPl4eM4AECpJ2wntg5SZ6Ox7oEv29OiNLqSlTmdgaRtFy1PmmHt+tp1VsLs7h
ahplHm59RIEoCKfGvJzVVXrcjlBWlsIwCSYQTUUvyDkekfy6Gs9dVjCfSsdv9bWP
z/yh15edZ9jX6pqiPc32tIpJNh33UgpHdR3NU/3VM9PMbLWsI/nhl6YbQRLKcvFh
D/qinlHBHujKv5SMDJTwSrZuf1crulZw2En2jMdlPOhpJJQxavJWGo7ynSJzgwaM
6mKM71s1xd9PdxCfD/SBogjM+ZgryJEXvY9LS40Noi5FGj9j5/oa5jXMbA/eTlCr
L6TEJLzTAxb1ql1Y4Qu15zuoUvKgp9FFC2QeDT9sCHNQv/kuqczvHBsS9v5SzDb0
Ut6pkVZc8fRgkP3qNgRA7ceps4rhn6aNgCIzVK8Ptwjbc9R+XGC42ubKtmkBGMqV
9CXVSriKcp7xMDKaC2urt7Uv2IONID9eMaeU+7YqszRmxluPgiT+na2J1TJmpYJr
1hU1hqRX+OrX7XAmOGYjfHUqa+BXP717TWyjr8kAuOK9PAIQ3Y4GSzA+YkzYvTAu
oLA1aOupjBm2+SJNJZn7e9ebMD2V7g+rDMAEcRRV2vFkVfMUNrvdTjJUfdrPCNxY
77NcLvEMDlSGOKU8i5Nx9danbtmts2FjvIa891hnFunM9BEsII+LV2ejnMJlFZ/I
mKuNdCU5DgB2D5kMoXfUduux+XQORoLgQPA2d0NPyWhnJLh+ppK1m5P3bW3pYRCs
VvmxCx+i7hqE8H2Qg4edn5crIFLx1jFjLuU7JjVVdkITeAQpUGmvwimF23eXz0Ol
RDSEIU/dchybSi73UFSqwDu4quywr0yyjyrtbb4byBjyGfBfMQrKuYkeW/vE5lnQ
f6PGtSDzb8eXqgUzg1LIzwc0PoNAayvuntGvsVdKqSMJwEBn0iZ2HAW+4/vexCaS
9UszJoeHpKaWwvlo2DyUUPVHLkta03lmERHT4l59oB90eDtIUkcYFVa4H5h4W72B
FLfflF/MGdHYJCcAV/kjni/Z5HZsq2NKg8MdfhqM8jNtr+JNRglo42e/aBKMIuaO
lBzr9jWOjODiSmIow9QZTEvPonhiBugpQYMD0eURkdY4aTcc9HrGCJGbmIXdjtlm
GyQQG9I0rh2A3/H1bGYROUjI3e4BtvCcGkpNcj0fproGe5ttlryvhEWc0E8vF6zm
geuj78XjzAa4q2D8NXAcG87ra5mf/C9t4Hh0/Pq29ffUnLK5rAv/vsccMVRQSt7I
yVsj8SrSKSVkdY/8GroHzGhC9y1rl5CRV0YaGf+oDoYzP4Eh4cX+IcVkssQJ9N1f
apGH6PG+HYVnSusOoSL1pmM8IvZB6tvKbB8VOHX2EQnY68LYZ+kI0skeyNvhjj4B
mNr69b4jb82TU7O20Ia2PrwjUDo5EcIQ9hzH1Lp+zVvOIKleNRneVNnslpuDjHh2
2tnQlzkw1ZSYhJ7WiMH5bicvD2En1DVrazoEXDcMgCmox1IWL4GdINL4C2ve1Bye
+tvsKILcOdXDLH+orhQl8UpU6ciylofs5nno/MFUQlv1vRwI7GvRokeelgLVCJ6i
7zmIILBFRSxY8vyiDDZG41rD5WTuShnJ4vrpmaxMuDU7jFI+A/+TICsT60mBJEHz
tJJjZscwIFA79UjUxk2pBE746AdJnBcT5N1fThz+hXX8x+gH7h8nxCwg/qmZKSEQ
wvEOZMSAiLinfHotonSH2//v6N7jhtnlKkQkra0lXos+hD5J3HHhaoyobdZaY3zl
iFIqy9mnGT+dy/cJupk+wBQFKb+JjDOyAsuGHD2CIbn2QP8dMl8UHv0ayJEHbmiX
3wXqE+HGvHUrvWE78YYj/NdKpG7Mjgw74Ot/GtuzWTZ8BcnZK1wEmS6eOqaO+J1g
kTo2oGvypNxI5p4rldHvga4iSoK70neHaxInHJTvjA0A9ds5x8DiwWcI4h4NFeDg
Kn5znRLf/y3DnYV5jXWmBW9h1K0upzuX5elv5WzTdo1hD0I8Wdm44bUIPioazuV1
3w0N04PPW7W97r/gnn3mIHAP1czVtnor2RiNjoPhwVAXsU03r952EGD1IwKfO2Jl
CUhNIFr6Be7Z7HAF5/QNoFcFRFVjzDT43CLyS76EiqDgT6JY5BiqJeos6lRYPeT4
2WUFYFAyCPy+G0cOvO0lsIXskj+ulmTSom9DYI06TpMCSiLaq7qDKYIUE78d4uOx
0/YCzCzwku2LN2cWuqFCC/n1Rbh6x7sEAv7WsXe0ErX19P/Aw92MlWVAF+86GGjH
Nfe+vF8YeHL0GBemwCE7hUaiVyR3JbCHcm/EabRB0p+tb7B9w5GKH9izOY1AbPus
KtJJJCqdyMxcftYcQJaSY6iB9Xz7PWjkgf400xQps/DRG1wNp4IJ/3KTGj57LUF7
igiIqBBJqyGfxyID0gZgIaG/iZ3xlhug0GfCKhCqr6CuBDbSNgiHtntzVxqy2MXn
PvdqIZikWx4daG/CNueDvnTEuA+Sz9UEgkiwFGVpEyHKX5JQOy1AHkk8NbMWT21d
hM+sADcEyhmiyqfgltdybeCKqdZWPVLZqubg8NmpJvhPhKJtKDWBG9X5+53HG/v5
2qL5qkgwMPgJ2BNuZeGc3F06Zlmq25GKB3HOO3t3D0KoOuKe+LsmzeuqkPS0oYWA
5T7qvGVdV5qUcGObzOZk4D+zePoxxSLbjV6nOx5DwdtFK/6QGTNfzbvr2lbnRWsB
BICPk2Ms197aPzgmcd+gWJcKyrihhB3V9V393QKpj3FI1wv/7BAleZb/0w662vxj
a9VydAylpK+kcHRF4kOIvr8qYAjIiMHsITrZFJo5CGgjLSFZJNZ+BFOM2I/lmwEp
wWlqQnKwDC16djNhBjLYLYC2yWO6ippZva4JyFFZzofD8Veo5TEj1WPfCWXSvYAQ
58Fzpx1eK9QWiTrd59U6kV3RN2Tw9S5KkAYZrzVflfDKQ7AVlEauDYBqtnawGURK
/gTMTTn0unu8s79QkhH8/ul3bhyDXHzC0mPu+qah1P2vI5uFMnSaZIQ66/VPSRyo
l+wJe+lsKMq/SYwkXqFR6uT4vSvCON1Rrfl42OTU7LwpIjoGu0UMHt+JUFxsnHFr
DvsJyTxjSIKEA676nbrS4GcVenPP2xom/mZaExBaemkhKh5Anm016fpZawLx6q9M
ehqRnu36hlfhip9JfkIEluvB1tPuThxJpRaoXp7tt+W7K9kRZ1Z4qxisscUkymDe
oFsDqJwpBXRZg0aCa8hkchiC8QhTGjFajRXD94J7c3BhbacjVtQ9W42sUrLcKEyZ
Ijhmtq0MWuQd+BTYVzOREroqvZprCgV7hvQZ6TMqDFh7mIx4+gesjjppCBxRs6M2
ftd62+7YqV1KLAxnsjr9xO6czw53rENWrbvURT2Vc9NUlMGcAE12JmvPCQJnzXCs
zwRoRUo3O5Y2PAtnXeTBqe4AYA/mTtcVA0l01jADpTpIicyvXdtnCBR5iat24Ddh
ivOIG9EvhsiSbrUXbak6goGHUn6BkElbuCJ0ABvCLzid9iAzmyhh9xY111cCWFk3
7HHT30qd9HnSdJnAeBA6rM5U6cGLMM/4oVpEfeZLUpBI2Zvb7M0cyvW9ABl6ACXT
jezJx7Bzf96Vj2uCDwcM8aU0fZdew3+1o1YS6dYxs5RdJr4XZ3FEpPNefAW0CEdf
1e+8CkS9n/8zJ5zfRDNdrsWxRcAx3/F545AxQlDqF368gBzuVTv3TV8nNqWK40KV
QVv8C0E4QDYnyMzIVw+yIrih7cnICde0zoHIQNybEQthvYPazR43yXNHsXKZgyW9
4C01QSQkwiE46+SglTNqk1jfjTwGsjNiZj4ENqp1ipUj9wzoqpaBgnNaG2/C1zYP
bD/r29/L6/CMwjdSL7+fR6W76fDAxd5Lb4+ZFmRSfSiLdMZ0vSMFMfpc4nUnxetQ
QxZPmWQ0QSOhaJHz3EPBkKM85RDCeNhNPuoYVHTGIHGa5LxiX93Hjq4xykjtQhdj
zBzInmxYDkGio2jjTYNojMgmPdHASUTdWQvNoHmcm/QPkm4BhcwHw+Ou0GZshnkm
aJ8KTdY28UfN4J2Y3bGzI6P0n/zmc39Q0qC08ocKz4fWyHQuxyv8M9UZjMisU6DZ
0lwyVDy8/SvVInOGXVU6OZgPJ4b2xSks7h1eXeqRgiQ2SJiibosjkejWDvP2qDh0
AWe8aqawVV4EUrruTOMvK8llg1e5dUASX+VI8Dl3u1CuOSj8AAodgUphFhQsA8NL
WoAft6bCv6u1caIVJAaGeeeiVfW84XfbL1wimn4ZtH8pyGzLVcSdQVRc889JMOvD
luy14SI9IH9+8np03pcegqpywcII6Fm2kQ6WvMKRBNSTFtyOjvFovI1ZzfgrCKAU
uJS6T5pq0+thNFldRphYzHP3/I2pwgjDdQGyBj5H5yUEoPJ8UvMYP/Pb9HpW0bRu
8FHXKUDT7vDFtqBCKqRkoFc5pz/EKGr4ZcUqtOYf1iroS5Rh7PFlaW1NnbNR7mcn
Bt4WdYDgi1gt+h7UMZem2pwlYyDcxA5zt3dQhVyvGBYVrGquruEeKff76BluJErq
sTgNwZGvHsXAsbV9LlhIYJ5UuDkiqcS8N+qrNPP6rUBoK8zimJyISEbUDWn1NVER
yuot/6fmAvk9kKbCfEFFslhmyQSIejM75J5D2rGSh4jKDJBCf+YOwwMxiM5LGxUn
99F+2OgTFjotDC5ceLcByAE4+ycu1jRvc3vuGf/JPoRjWH3h5czu6wR5o6ByZdSs
lgz6iPxX0PhmaoJUhP79mvb34WHSYmNGPN1MTsg/xlcQifg14cUhR5w/rP8MYz+2
uYp1xvAGSnR6v03HOO26RyBoJQJKcaN3RkiMqMldWSKyX9IsZU2VzMN4+9nuXMov
CO2bxL2MZMFH3LA0tTfq29jByncOoXt82PgBlrI79wU5ulYDIwrG/fip3bBGGIE4
+0V6reJhS3P26aEoiKXKiD186Awmrs1pFw5O/dKWi2KKUfS5fNSoc/0FKyOeJV4i
+pgonsJPp4TC8q1LsZU2N/C677ZnIB6j56kNcaRxIxCUrXyPm+gjJaXEXHUiBsXK
Ve4TZp7+Fs7EdFac5uQBMuyxIGwtl3MMKbc3+6nvJbNmOvi7rUZf6dGNJxNiuPM8
6KWhhA6nGlrNDUG2hAIDaCjEx3fTGOxCN9kSW20bvRZ7I73Fsx88UKfaDU/btEPx
VEnF/HMkb1BfOQma2Fx7OuWME9bruGa17NMHJgH6WVWIq9Kyp+m234lr+1miw562
GeuHsIxsytlF8QD699ak3s3Z0vVw7lofsja45dYLrh52MV2mNRYKocqQJDNrr8dq
yhZt+xTubrEWFjkWEf7nGJTE2hdnTvAT4vrhxMRu/G6hpvI1nPRxpfvUTo949D4F
GrBxX/FBgRqef99JCnqgsV2qMq/eavKgRdP+7adv5oWrIb3vk0gXAH11vieoea2H
B6hG8KRfqkIdfppuyke3Mx+KYPXE+LOu2lpJJM8TRzOGExms7a7aAxuoD1LiRTr8
Qk3obiSHq1VB38BWJfmuaLDT2d0c3W6taKAMHHvZaqfmVGTB+ERa5L5I75DrmAZZ
7c1MO9dq5qC3Li2HfX3EAPEQDXsKf8/I3/UTYVH+E+iB6v3gVwQfAHLg66x9nVlC
R1JI9h0+SUXZaV8gsjvjcOsD8lIzF+7t3QY8qSQXl8grkTh4lmcM9aON6nUzRjfM
k1Six33sNG+dAvTWlA0hvX9YIAjG42C09CSoetBUHXsNbDLXj3QXRrDdj4rmkIGf
+FSVbAI4ZFC9OnBbsOjqqD6VJCdnuy0NRp9u7VBRbj7cBd8Y6DSQzISuROUmEhSY
h+HX1+9UATMkbW8h0XSTN6adxz7EKPoWOAcxv4/dfV0uHMQEMMieYcj3TDCFM5w4
hmWSFxA+gU2FnZ2UZdQV4JvmMMTNZuEJydDFsQ5BW8MeKQQW7nMdNpjUJHOd1tKH
zbRluc5DuCiDBC+BJrNDrqqTmYIlso9px0axhAXU4mZSSXt/NH5WuoVm1X/TsXrO
mibBr4fnjg2A58DzTBoYoqx4Ev7JmvJ1VJ64VqK3UF8NLxPlD/TaoVMTuCGU8rbu
MMwFRSwsx5TCQj1uYr6bT5kiJXR2hs7DwU3lH7eqec8qOz3ziTIM6iwd28frgU6V
as0fVrsF30lt49q9q6BojZrtmSLSToxd8tbvEjsd6GQSRpweCSeLAgUTUhfD1wr6
GKWVb617OVWJM6NFVCxb3p6ors7yqUi4v6Vou2TygfibbXQlciDouxyD9LzHSZ6Z
Az+g5eap/e4E3Pf5+fGRM5o595P/1xD8uiyad72IGWeCFsyHdA9gbBTmRfqZfenB
LVrZ8Bzs1H7cdS3thr+A+wBVdjUWN4ChHL4uRqOzlNaCapmE96Vr1v9DjH1/cmeA
P01cTeut2iNl2kvow9aJTw/PI4es+M1P9hRAVS3P3Harbj/dfq6JmbKqBByxQocR
PXt7jJUo2wXwdrI6m/DsyH0xgXYRXiOhcJqMrXmeXUeGSwMAj1AVyTq9vQESjnF8
F9LOtOxJZqppOZiwESguH/CvYsIX+EsdgbaMc5ZJQ+9xQ2TyLD9f9niAtzvCuDN0
t4nloDC4aAYQ++fmJBAH1/MLgE7dzCDfGK2WKMP1/Pv1wF4E+//R5jyEu4B8rz5/
0fIebgZXPwkr0VldtgF/gdBNVzyn2EHm4ppRkbwDRKEvW4pBPWzR6G2hn5lmcdOs
JqyS5oRSANXUpnqkAlrOrzWCtYl1SfXVJzkP7LRxukADZTKhgrnWWQBJciXEnDnY
HCuSfSIsXG8ELH1mRQQ94AQowo7b6h8i6P6bDl6WgARGfCRFHjFVukG6AEn3hNB9
izBpm5gGqirdWCYPTyOVdqmCYu/W75AYvE2mynIsdH5rKboeiQ+H+2dTk1ilVBX2
bURGjx3LBjzMRvR2o134G1vNKO3Wp70nmLs0QtJedyMR97j04/ENMu1FPWdWXfr7
Ss0dYP3kvAUL72pTkVSHTiTbp0/VKbUEkGR/9mTii3atc2d76jCEAe/fMdQMts4+
05GzjPDiqQD2eTYqXNUVpSoOKOx39iFNYbJW6Ii3oQlIuQi3JCnfz2sLB0rUV80I
ntc5j/DoPIu6zfETt76r9Wdu9ZB+okdWHAI4yKnq1vdZHbwo28GPu6TLS+qHgrZ6
q7YVctQw10PvAyRWx8q1kn6LMxoczGdWuNwl/NHqUpk58zjwgr/bbwqmKjqc85YR
GR1KgjXXQcV3/jq72HfuDWTVASOYk0+XeN/wvTN+qlVJ29eJKyS4wMQfWx6QPOUZ
QorXylFRJdqhupe35fSmsBlYnjjSr8/BxP422GnQNw0XDC7TrjhQ6g2WwVUrHj5c
F656gNr940usI9TeT6FF49muyG/EaMTAQhKp1dn5BC/axYet5DxB1+/vMboFxTrl
XzWUgqVxKmfkwBWTkfbQ8Z7jCcQ3LMx+ioutRqlCMzYpi+JVeBeQQShyapTjqzxD
RD2cO6s+YT+/9pel43K3BCQDso59n2fPmqJSg/PYLDl0hw5mBnoh0foSt42DPvSA
QweQKH0bxgi445Cc7r0zLQK81ccT6JtZcQRrzVlectqFCdlexLHvsytpsLfmGX71
Q7MmQRSSLhNfZ04rOWNe1xtESiXVmu7TzQexGY8rNl0/bf8RtcubzmxIZqeDOdve
HE/rFhPkKzCR+Z5p2tq4ET++PM7iWi01n9ou1Od8gZp/q9Mrqa07BSmgld+anqcR
mG2uWOz8b3IKuTEkaQMZeVLoXvFFfeg2i+ABh+hAhbyGPLFbl1pmnF0qTY9sjpES
hVTSR1cbvZNKs5IkhALPa3jsosIP+EN5cIDlamjY3gwwIvO2ZK7Je91pFmAn/cxI
/qZB+qXxE3mkSi+BLtfWeYzexnF/3u0qS1spim4ruaZunJJyterKk2g9PQtyDcO2
CpD8P0hNAOTIxiVl+/1GVC5JOHm3GbYa3DwqEXhjPFHwYRIIeUe1sPVVywQMKaiG
4sfSwooOFIUVaF/SoyLIw+XLDPlXdCk55m0NQB00id+En9qh7zErq+TEFlD6TO57
vXT5rzpGEhFNu4S6QP/BQBHcbhV/V4hurVnLcIh8lzQnord4WYGRxlFaX/tm6Z+V
2MFVn5mStPh23P5mkc3Xxl1BU5QG2cKeRLBEmhG2WN3zODaV5oScGAA5KDnilun3
t5hjoLcj/BDg/fbYsaV9Mu2Hy7usW3Oav4jD8/3tJCC7op55FNbtmG7qxdCIPd9k
EWjBQo+bGiV/ctQIL9wVazohSe1hGVzQGyR381unrJdeFF6izBVate2vU6GtXaMe
1c+GueCxE914lWAl+TepWQyEzUGiHyErflsZIdLjufSWco4vQowMlybOQQ6wLdY/
iy1X6bERDYXg0IYm9fj3H1x7R7Wq6R7xYkK4zPc9ZhD5u28yJ0WSZjT4EXVoAaTU
zuV7IWpwRPuUx/SAdu2YyMy89IY+WVdVM39ryNoGcrK5Pyfay0TOKbv6nbPleLw3
AFbqyervK8zWQ7fw8lymCE3decq+H2n4vk/pYu5xBzP8mEFdOJ2nENBSNEises/b
Lc++NgtjsrNfeJpDBsgsmsos+X3y3CgZKrCM18UeoecaA+qkF5djxeiTpkGCCLNi
xkkm399DHC24Ch3w9y2ERe8FTG/e3ZuQcJJvmwklyX3YeA+gNG6ZMfJgKGl/MVer
ZhJEydJm+t6m5usgRnX9y09GMXZ3NhJYBvznn2ut8X4GCzWbxbO/OCMT/UYDwVWT
wM/0G5dfiraGgTs1XMZXOHtRaqj9CN8wDxJ3l9/Zeam0jR7rHvB7KJ/myWNlNKDR
6ZpamGPAF551NC0xzjTJs6zDfBgml++8JC0FjZweQ6RDy84gMrO9NRwKolneA7mF
et6Z0rm8O2cj9cMvcgOEnPqQOTj4QAmP3ch1dHZZ5P+YjPVR9fsFyo6rCW9JDMrv
GSsk2r+t8q7x1mNoW4A0KlYuLKPvU7Sc9sI3iiYPozlzG1LlJ36CjP8r1H1oW40d
bGZTIzBiBvKVUlpdmgta1k8XSUTN/Lev5IDqKYmWib5zbqSIP7MNu1P5Gj/Zf4Mm
wDZXg/YygSAV7QgtXVOml0PaIEMKDpiApIx5t1Zdy3On66Js9bm4wjCVXZvLqsWj
pki/b2loK+o96ZgM/ZYSYD/yBt1PRZ/sQCyLC+0oHK3Aqft8loosNMgmRwCur8Jh
LPf08+7n40Vo0qDu8LXBx3G1XudR7wfBwS89FG3dDYNTD0iin3rIklwSPgbT6qhp
JqLxWSa+VJTRI6cnYj/m6oea9wjyB+5lJlOo+NN617K7aEHqwxcoHVPEFDnDh/LN
ZyCQ9NjeGmRXeG0gpVsUPeVDlwRDTvFcJVxI1aoY8d9edm8zhmPlK1B8OMiHgTbO
u/jgsBSWpeiHMeSLNyd+e3o+LOz+3sqUtVCVHFClxKgfK8P6AgCiURcxEVSu4kMv
kKWBJN/LMuqfGwjoF0ia9cT//D8cDwk/AmZ8zZG2Mbofepnd5JlYE+otUNB1+87E
T9TvNAvSqQESuCPpbodrDm2CtnTJqK1Ii6fFZ0T/gkBoz7sQCPQJDHTkSlJiUgE8
fxVvooq/tyrFn4lNjBHSTN0LhC6fm8sEZwRtEr35mamougEs3KiQlRPB6ni8bEqa
Vt3Qy9l29B8aRBqU+++m+JKd/MRgmpFhMp7qPhVmyWXPCVKrVqInErrBE5bipubm
spoiLIFR/V70d85GVFU0izdaZs2VbUwhNyy04GXUK+3bttgIN9/mDQ52rzqhL6lI
vQiXAyyJbBU1sYV7+ByfyemaayAdzo/hp0PHomdNupl55t0Db9Ikvs7EdMTsPIh0
WIjg2SQT+i9p9Lfd7rnhS0EoguMRTAkpO9abF2Q+0+uYdDObXimY9vMK5shSLenP
6DwyEz6UOQgID806uM35dOkkWQQYG8fWEGNm6TNbkg471fIo1MBrKnx1sW9u+RNK
Tc24D8No1IwP5S5UIbDS4Vki1NZbo0D3fsrDP6ABK7zLgPHP4YRs48YrH//n/mZT
PZWFFRPjbuS9oh9kwEE+toRhAwbb8GXWnXQLTNQMgPzzRhZ/VEkE5lPxhKXxk5ys
r4ww+ZQiKx703am5lm1IqYM5SEcxHZsDqYWPi7ORGQrgb3tEYzuUYxTIZyoClORq
SlSpFpiP2VHcIv82FOceblkXZK4PGeBI+lCMGfAiXBDLVrjxe0UZa+b+HqBU378p
VzIYnLTec1IphRdiY5Pm+KfI92BiXgnTu42AxWf2Kpkjb5OOqLana4LtDTfznO2X
8klH90fn/GFrbKceMhfUzz1LdaRbI+fQwcZJ2bdV9kkEQ/ivnv101rns7IO2+WkZ
SISSJDhfeuejFaVAHI/W5/N+pxzEG0u9xD3XPCXEm5oA1SOkZ5DxjeEku+zb0lur
KIctj7rvZfg1NGzSAHPoP7pNkpTUu0UYM0olJ/bl5kSeXqva1vJI/xl328CyHRxC
XmXWomCUBFmvL5H/rRfrHcGZAzIa8j+47nSkLIHH/2qLyt7GXyxfl8jXvXBszw4X
PmJh6nmTILCywVCu9SrFcEHYl2i/CLtIVWBp9+RPw8l2CP4jQNeFYqz595H60aBc
GQD0V7wGM82KjjjdsphZym30+fB3UOhdvM3c7veHDBmPMBkyDOPs+gPK4LYukdr4
XydsFrRKM5OsOi0CztyLBqQ8G5Rm972f4ibxiysVc9lo6qNZ4VNswEqrbQ4MROID
UY58mWYS+8+79Hp8S3eWOF2ZFPSi7dLl7XMwKr90CFJI1LvUexNSrARTuab36pHF
2KEeIUYFBALrLu79HtrlmCM0mvDN0vKS7NecqlnCQCCffmP5Wn4IPfpwUYofuXRy
/UiVqvNqI8dArOlaZ22VNkBmvw/dWQ2KZwhwz5IoWwqctd4U74ZHXWtMbuVMUrir
J6rxjeBHb2npYFyPGYzJlTKM2G4+Yj8JYb35LV0KnD1UgapL78hn9RfwkPnHnW3G
criYcy5regbPvVmIk2jR0RFbFJgXBnzwKC5xJBOi8w3ZtwV4Pk7dI67/6vhmg5Y7
+ybc0IMrpgd+XmcSueJNDPQZ7VdEc1dp2PTV1oYE7LgorAqzFSspvhHLDah9NF/H
F//6wGBP12dRQTTBIaoQ5ceIkvYcoAwPSkW0+zPsRywxyHkYVtZvIwbX2unH82p/
gfktLghJYyu0Vi4lYxTvmbfbvQ0Owzrwx23f7MVV5GILiq1nUDm5qy3k46/m7DRK
bX/Kf3Ief3ILxC+iA53B+NqE5jRYMqglBwY6JVeOZB6WxuyqUQ+Fv52rvDYuHill
Lo97wjJPNcww0aKbrHCYlwPkjhDZasoKHHOrMtT3cQEyJRS7GY29oK4lbyMZAAZ5
/WUufRSC2sYSGrT6UwEmK1v2591h9p+cVfS2dffBMq3LPC/EtNYrELWlrpVd7kL7
afpawZ479HzhbfXynF3mAQ9mr7GMaI6ZQdsdBufXZC2NCcMsSEq0mnxrhkKYmhex
gui12BoOEoLvLxlT3xWc6Q4BKCFgPV0mYONKeZAknE/LB3p/foSzi6fNISS6b98D
+I5dgYoKcqc8I4tFLFrbCMIiPEFcVItUC/GjfWVVKZKBRGf50vD31xrtu71+HaQS
Vf11Dt/eeAShsGKJr+tNt2CnH3jUw/SGW0GZV8uZhvt9qK8lnxl5WSvH8XBla8PM
3WojC+l1inJyWpz4O5QgZsznLPJLx+dPVhiQLJbN15BFm6cLV08T99AsFp6NI5hK
J18DkDhYfMUynVbqVkCEpt+o1+NuSQjzmn0REoF7HChMaE6AFjClreqwHP0M1oJe
hzDDqC/HBhWcckwJIeNOX33B0oQeTYNhBjEFT9qFICcdoqCBKlbx2LmM9hWG39Ym
9NRmsbjV/N2GguT+H1MdJv8ODvRE4dgk/jRNboAIyvuIjMHE5yBKnpVYFEd3LFER
l75VGwJFf3zbizzoUgQTmrer30KX/H4UsQyIsBdQMdDhODpIdXYW5TIzcTYnCMkQ
XKeIYutXdKNVhkkkhGQMiurQ/3BECrWS8+FhpjG5/rUe5KUZ9/U0zsMYqadcflkj
N8WE7tXg2dL0n2jaYqMp+pxe0G9RTPmDT9uVlNVuDPtcG2CuUe4IJdpxp8wx8Em+
GLqQvOzgdOCFD7ibkBdeAjOwJjcdTM9hVDbClYkDZrw1UJNvjKsGGRGXTXkRxZAV
6GlNQk7s2C+03I0vVifLqJXe4hoZnylG8Xx5ZtGv0YhUSIat5acWyZYK8HC9+oIE
6KmPJ8WQ62C23DXymDMnH3s0TuCzxYcyxSsQwe+I7Qmps1K0pfupLeuNpRmNMQEz
x+1SPEryixGUOMCFTGXRYBIOop2CHWsdi2UiSktPg5yiU3bMAVSCYzv2JctvLK66
Rk1lIc3KRYxd/7M4OjYfIcprX1e1NmGswLJV3h/ijHJrctysM10d0TvQnf2wbr8p
6dMvLAJybrgOsy+hCIPcuxFbbwwumtOrf7JCoV6oxvYR3mHL5GJ06JE9DMP69rUc
l7uQ91qs2U31Nj0dpiDvC3JOmwX0jUhJI1ZClgO/2W0H8L1cJi7RDYBxm1wWUx/a
ujzJpo24Km2t6ETwBtTNKce7WWUqn4311jU9N4mXXgginse041Rx6YTXaw25Me98
/d/GiEsUabaGgbR2q+ZVworYnjUWbAC00m/8q2yt8rm+L1mRKMj2EtY5pQkEHpbw
susSo7D4y8OX4oaEueoRnwXeKUvJ4LHP/pB6fMmy8d8KcKbDv4PqfHwsSfwNo+HF
Spf7S704f3dZ2l2SlLib+6wuBDBOgO5LfmdTfz+fEmaW3aWkEMVGKlvby5GA8aKO
EOdUAeJncUWfHpRIuRdQpqLrDKkx4tw6YYAmtJrJpVlkyMPyzbUAW5yPZELIMEJS
kh+o5aQU/26Ihi06HwzV6nUikTvrVD4w8voW/v8xq32zMmRVgfkdSzUrEDdCvL5Y
kzUfAa09CIjcoKpm3KzMh8s7KleKxrGcjsv0WNUq3/gRtxqq0kG2N1w03d3AObjn
/1jDI2RaGg6Z2E4jBQ7v+oZqpRffWznpfl5vwYeMrUl9i5QNU73LgPsEHuPNPYS3
W/oRcmbgWWeM1+BKS0pPRaSm8F7o4dTrB10TElxVuuw8Tx1kG0hSketkXlCjEXRe
yh/CFLKooKbM+Tfg3jaitIT07SMEfF/X5NePaGy97DIgcFLQGNg9tsdQfQ5yhQSe
IDwf9kLsha+cFv4/DMmUIZHbGwpCa8cwLaaZLZbKWsOgQQOSPKeUSUJj/bC7Y3/u
qR/bZnsLnowH0u2aDySD4caihHZQiDP36IbTX8JMNx7Qz6kIz9Ta7VJ/DmCFG/DV
VEQ8YWSRrbWVvMj9aLMNK4oTm0EBB2vsu0x/6DTVpsZa2XE0n6HrQgz8a9AMANSU
RWyycf18uCObH8cUM30iMqNhVwfFiCKthCflWh5QPNx6AGC8pv701RXTyI9fLCWz
QOW/JMGQdy2N04rRE0Lah6GeGaBwmf3CoHYnKEHvdGtavmhLw+JrXhGDSosrz3wu
G0WBiVz/EAzjralbpguJLlI6Cl/6jb8xSkVhtF7dQzYAE5tIkrB2MGwSajsOr75V
nN5Ucb0pyf079vXaUIGmfzvzhPJIprV3+7VSGwn3LMXatf89MtRbZbgCr2U0RJfT
6ZW4DZe0QNNWcFe6IHqkmYrHmKjmhPLVXNlW9MIscnZd7Sr9xt6helPsxNmFg3aI
vyO81fL0TGe1rWDSTSti6KDqy+hbM/mh+wd06N+yr+zg6hVjGin2JQVq+Hbcr75Y
Tk4NXjWdea10GvBw8XGMuhQNAX8hSxYcQRJNI/Zr/SklsOOgXUgmxeRhnFnGHgQj
BTxXN8rxHeJFOaS0evtwQ6HhHp8p4YtICthOrrue6z4UsX036cGGZasWbMOHBFst
xCEw6L6l6E4hEYSHYYI8msnazrZCet1ZeABlYXKwjQJH/ZCPGw4XM76hJfzIeT06
6QvL1Wok8KaLu+dNQF1UaF6513aWNdEKTRxVDThj2UQQ/gX2DyLR+7VlAGCGT4CB
6d1QDjDVuOIXzGJA6zhHDvRoDIHEALT0UZYalEtHvKefO9ZvL8+AWZs2HHIhZdCN
Ko7JDOz+PvlZbEIRr5Gcrda2dIkcPT+Yk7hpsofyyKGKD2XJF+mTlVwnVKRckj+B
anN0ksjkv7wmg+I3Im0wx8b1zJeG/7rGTwoPCpVNVf5NnQV3PWD1slkT2uw4YcaR
vopQqAalKP08pKWHci/1LEWPkok40LyyoRjWriK3WK44pZf5sU7+Ui6/pJeFs+7A
NwsAPTlmYqE92340FIe5abCphGAmJZNyCTNhh49RYu3PWSmXiT2JuTsZE5sumMtx
TRI6beUR4PbqLhxJkSCpffPdm1SlQVAXms7naClZ/p8329N+PvK13WDMaaEb7qL2
wDGAnHZI9LNAyNw1NgN3VPpCcfQm2lcNzKKznCTk/U6tmkCI1fNPP7sbPV0sUFO3
aMZwzIMtTIYmPJjlATAc3gyvObSeYKdkpTtxjB1KZO+WZQ4zN1guxRIa3tOC7Wki
QyUtj9Bnf5LeR7PhrBcKIa4wjHIw2bG6hD1NnbX3c+VBQI0FZs8jC80fcnyXt331
svgtgZJ/J0jFZAj1dtQlniOeUmKGwLOvb/oknFkgSdEAdy6m6SovX+L/IFBfCAh9
IZCSt9+1MJtyrCOVCchZQFrgaKSDhH3OibvAyFZmGqWbiTG8Arkvhl0BEFIgG9a5
AYrvr+YAm5PjRhmVwGzP4eCBSlBu29gX8UpbnL53QgGM3/Rso512RWxH7KyfADnj
eCg5YBOGXlvgdESUJa/5eZCtjWP1Cev4Abmb+TBqp0jV/kqXiZ1eDGSfiLu+n9l3
jYZqXJmI+ChVRsFzi1vCRLHlYkz+6SbKKDJ9/g084OZw56/HUu6WwjhAQEJkgUqb
VcfTO6k+2ZtGzETuVzO/q3HTzwRgeiaXLKo1DuutEya05m+ySFPbVjce9wEzBWh+
jiXK6O66fS5hH/URUBq7MXsCEteBRkQMPYDMWbG6sRTBTxtCRynEpmRHwAEq5Wln
znaly2hdh6tFv8j6QMC8e/0K9qb6LrKP4s93Gj8d0vNkcH2cyP7WLemiX3bT72Ls
JFsYT+BUje1NoOfoOatFWt4Qgtt+kuVpqFI4MazGLiaosWYTfOwq/TMzVTlTmQWo
KBQ6TWiQXLYfF3gqciPW8Lnax8ZQ3IcFxhKxDYrogqVfShKgyw0NEUcdsS8UheBI
dQEhrqlg89ylEXs8/ALDC3hh6RL7AlI27r1pCkGRQBIMO9DgTTkLjAecciIBPYqn
ljt8+u2bVM8sWcCuUFhE1kadd3+c6tk/mKQTUWx4JjtSLI3ypsZFaT7f9oTYd6u9
bh8yQtj+QFFYmE5JeBiu6BprGYpfcis6u+2/lzK7hTObRKIuPd2EH6TJ4lzN2mMi
3OhpBQc1Dc1Qlpqo28WLBRL4OtaAql7vZkRA5GLU/MTnje5l4Ce3NKUJNj/NWVKJ
o7dIV/wTYHeigFYj3B4ULmHsh8d2EAEyv3MdGBbUeBTxWSy6F5LZxKi5Qbk7lupT
3z269VStpiw5s2u+5Nc5nDqjIk4OdCwOKCTIlgMbjB9lPgdSnWPbTzgB/a+p54xF
CdATW1ZIvVmbGqJa+mVEHsu292PnLPEQFgGgQ/PY6y5qFWqZPN74GSb3aDuniqGV
771Qv9H6ZcUqr+M+bh1Q8HlpkaRxzVc5gBbosWQ0ZdRuevgibE/zvhS8S14l4Osm
bw+oT7wR857HQQjmHK2fTGw1rpr0WEZy1KEZr5BTpigjVLP3cDcp+aSi1nh8jOwt
Q/eL9D0mk3kNfkgavKXuCg9wyATOv5dY7VbNYpJKlQXxp/XreKsAmQ8IqOaFG3ni
TSO5rhFDyQaN4sQKFOmShAnHjzfWmOplQ46ZgDwCYtKFzEF0gwyYOQYETIrDIC2L
ezCJuQ8n76eIvwRuMQntKFiCPin+yoG+Ju8kMnKejRrU10md/4LTKtAPC3HYxCev
p9D+JcTFZ0/uYK3nfN8bcDKkE3nSPTfxza/Ghn6keFZ8XqO7E2HYxOO96mv8GndZ
RMEE6utDthvl2D6FhfPtba8YRS1pdMpQ9EVVORCVeQe3UNTtDJMc2XydKJZsHvoK
LP2a2XOnzetSqRtHsskN8qjTkIO+W9IaosdMjK9O+YdwvO9dufDnqUdlVXFqeNEb
L09SUUo7JfOppcPJr0mqrSe+MU1S6S9fwDZLVvVMLMGqVQDdUe/IsM4K5GHhu2gZ
TT0ksth7l4f7zanD76/lBnBh0CHdHvgB0rdk1s3VR2jaiifNiliEeq9jyU4oFg23
85DmV4UMroLYD+GfZMrJhStCFDf0gI16vzEQORBJKO6aBc3fyp/NxRXE9bAS6kBX
LktbOdFtpj3djbhYTYjS5q28zG5uBetBJclxcDuFL7+bSd848pvT6chbEnOeAxgG
BkZyYJ7Sl/B3zLryZ+R2i6F2PxW2SOk0nS3p+f/MrAsxZOfjdI4s7clCxwj8JZGD
zcN5ZD7wGqcboljN93v7Zu9GXnLSyoEwEuhUsnfoe4Cm6vSJGkLnUP373W8upS1Q
9NQEYOCHQxjevCjRqNbjmKM4e4uM0brv7sKhdcpv/XXxpPQnS+p8rCMlTCiKZm4q
Z8/NDArNMYW0WM1fJSqB5pvWnJUm98QSOJBkIYgZN27gFvTBxtrav1vYArAypc6d
Nk7bJeg8Hhd3oghiavHR/YRpvBm9pBtZ/YS9w3a1OItTaLy240XcVYG3n6hX5/3R
Y2IUlYoSJKGr2BIx+xGdNgppjiKaxsJ/7HfaHRm1zU64HVtrh/fjLTry8eH9exWY
trmFPhROXsH7bEeA7VaAJ+pVmRKMY9ixdwo46uTmcnc43u0szl5QzMVfdHGA8s0u
5HIj+YlA9SyguWdGZuZzlJowCyrVV2aHobOJW2SRTUwMRQD4dm7io/atBz3VcdTZ
W+YHgBeRepNiL3YcgqgN8xxTBLQmZ6IishyK8ps31GiR8i4v3736lGn5M+OxF0ae
Q0QwKvBAhAnW4eMsOe9ltv9oM6tJGaA8hpOTZVpy4lz4mnCRmpKoduR7gWeHq0Wi
vZmq1+8u4ZDhZ5D8BPG6ase+cCXrB3zdXFcF1seOP/OweuBe947t9WKQF3EePkP/
zQX8fGW7voSqHWwi7/Kwce8yrGOD2sFa8oS7Q3XML1ylZFmWT0FblkbfNzPI7de4
9kpL1UJkIdAzIUHPQEGqvY7XMh3Y2BoLmRMiEMNU3njbdR0Hs3MIQ4lCUi4weXby
v4ReBWRuiW8ryCalEGkipm4Bg9MIEb7Ihoedop/OulePxP5NQ3lwXG/PbcSg/PnE
jIbwmrvh0uaWcjSKroYSHIPuoyPQDxC7O/ZJzcsWrl0lwmUIu2uq338vrRNrR0RJ
nF7R/1dkTZFESmdV6ZrPleu4vQ/dtlwphS0EbIgEt1Gp/zbSyguzSPjRXt+UDXKd
q2JqD5Pa+K+IdSTWweQaQIxJx6f6MskZbEX3h2okdF4wD4lnhec1lvvpJkCTCScA
aw9v4/EfAU9vs0iiO10iOynWIQWJaDexnap6hrkovPhLWfmoiXe2+gF+kgorkERs
sZ4et20DK75LeF/X9rtflb5872ppK2AhB56r179dBqNhdCk5KtGkU5vrF/+gnxzr
2i0taoiVm5T5vnMxJsX8pnArYBY9vM0ugQ3caSQ5LQsbom6urZ53Q2lKA4BnGaPq
Y+hJCneosNe0zhHwNKr+gG6gtGUUnHlOLIsPxpVa6+pudh4+V5p7UG7nSdrDafpt
aEJJ6ok/hJcxu95MpIbMyl8KPPjpX0aqBBmghVks9VblJUJ5oKRT2PmIy6mwT2fA
CNeslxiRVhPFPT7PM43gTI5uWbqQSsiuajwXKHC/dw/4fn2mzF4eQ60W/crPGfSo
HqYPBdtg9SPmvPC3xJriU7Lj/JvumW98gykrgwOxY7TD0DsyAp3hqSkftRiZJ+yK
4uf0/GOwhxMgEdYHViX+RpuI06f41a7zcapVKh0sAWq97hM7eIUd2qo8MbeMpWaO
aIO4AEJV8xI7KVb2TdP4CEjg2q/yU9Vd3UstL/h0LAnB2mlL6mKWgeT87BvCI88z
/n6TaZ/5WmcDLYCM69jFdv/QTsxMGcvF3l5MDGo1qL0R2sSerVy41tpJ4lw92est
9mAaGu6DOe/fMFZ8NZNm2vFwksw90zk8u1riHmcH0JYoixoH2sN2Q6yUniYGs69b
hzGPDPgJO8k5ksIYG4Df5YM1uhFAUEt8zQAHmFNfSf6Yqq5s6nRadO/lB6nRHsoB
KFBpqzmrH3WCPJ0cF/GB+/zCZcJu30k7SqnbU1Qk+/e74ylndu/8wXKWeqPyj0rZ
BBLIMT+WQY4Ny9rtatf0MC+5OSjfS5ojjxMXnsWlMSFcYDcL++cijH198YbPF9Gw
K3uUDbA5jkQBWewhgx1fwYMM1zLzyfHHgsRLAZ74H6/FEOH8IVyIpZ3XSqkA+Ra5
TG/Z8cFnLVXR07E6qzrSCuRMki1U7OeVKe+W6kHPhGQg6WdMtczORApqU6bUurRX
i9192DO0HoFW4JAC6M7v0McFUD0ygvOWpd/Lt5E5ItagGnBlA0v3WMzy4NN9QpMu
RNxILE2c7Q/jM3hxKvox7BT12uz32I2nBq1E//bO6C4gpVy7lSbZitQVHKTkSeKl
sClPBD1Mby4UTp8+Quf7ofD4hyM/QNUalM4M9vq89/FIn1gpxrVTbVxuQ+xvavOp
Fw4H++SfbK5JBa0yFE/yylMtYqfIblWQA60gvyQmbm+Gfawd3wtJ2S3/rQ3lXgf6
hlTJZ45vKl3CqXNQYx5DH1PsxS8ahzeXRWVe8YygUGn4RUMYmNLuDEDMq6vNmvly
poxjvpdJ7mUnBSLSDwLgFD+cAtW/wsyNsuvPSVf2qUObrkFRP75fwt1Ps1uvYRr3
+nh7iRvwG4ozCsLO+NXCyzmMiGm6FDs51OXvTOgJkflmjruz4+r0JTh3a1rBHuWD
rkiA+ajImJ2APSc9cShSqbbSEP1VLk7+nO0MprMqVL1ghYvTBFFmGgkFcxcbfyi+
5r8Ef9xDk7xkkYYn7BtIXXFs8zApimojYecqS/LeCL0olZN9iXcFi7MGS0C0COuW
HEaKnQ3lTDtsVDtsvWZAp/rV/RrxRdDY8wJdnXRet66SYKy8YXikAS8B2YS3ntcv
RD3PlSon7cV8WI+vBUVtfm46C48yVvXTMW8qKD+sYbjA+I+FyBbJ6ssGLHxuJOUo
76EVizTuxWzYIqgy/Ydp3WHvG//vUap7WLO/x3rH3mvAJtFAicR1NPdsM8PPs8cC
0EEEwl20nizvhBLVOxQoICuc0eTXHPW+UEFpRv0MIB0LscBQiSEb9vJQNjNvOIb8
2GBj/H9+ZCxi2UqIwS0B/o0PBM6mK3RO6cEl09EZ2bfYhVg9+z6FmyOFpsxjWMS1
RQfKGHsvItllIUyqp/zLJWZaGEpE8GxKkp/WpOxH6zfJDBHVJn5DdT3/r+j//jnJ
W9cCs+qHrEQrIXBk5fRreXQccXJ2szQWa2zjrZFNZOc5gRl4FQaSqKLRg4sVKZdx
Q8JfnkH3BWHs0FFZ+8yZmsG6klQM1hbgFUt1zAMKEa/V37lWM8VuFPZTyi5xEEcP
d+ChNvXT2Z9ASSYACvj4CoGEKFo715CYeU/FqGukdb0+b9IMA80CtLSEV7GoBggi
LoRk5t5Z/fAN/ZZKV7GLSVNXpCBYLvk02sTwPvV1Cqt6xl86VvdkKxX9uOJVnuO6
+pQDQRZQ9o/8crOIP0IOnHqv7aFUNlvQC/aL9JFLzUmP9GhdDfDxqhjRXQ0/dQ3n
24nj/GvuvvsMhzhXJ75N6yMyu2dOg+mWuBdsUpXFrZfiSM8SBS2k2VjZJBTABEbW
roqGLPx3T3dkPhg45pDo69H2sBmkpYmvbjkJKya+3z7nt4diCSkzZlVOKbjXg2N0
RwBqKbmKyVDmsaD2NUjBaxzhYlB7TKLNAaJgUtRNAPFwQZlGBk/pEcCg6R56nJzN
+iuyXJzzm59wu47vAeT6OlCCEIdKC/XtCxIPQiRJPaoeNcuqEzE11hUDqG1O9Vdd
SFuCQx0sqCEbH2ghGpapa1eelp/Hh31GmJGaKRZna+Xn+BeX6wpa97f3AaDTKH1l
V20+CJOhkWUOTRJ5B0AyxNZcOPR8m+yfmoqtMMgZZMhPUb4R0c40e0gh4bszhxpf
moIwE/+4vRpQ+a2RKCMBAqctJRuH2mZLSE8dbS/xl6yVF1Y1sSYkAf6rJtX4p3h6
tLIDTvgOXWYL9/8RByuT5wqe6Y0heoRwPzMAwciQw0kTqSY3wmi0yAi+c0TSR7Fo
zOG5XjeuAwK8J0DyObdJU08gKUNxXbiTF7xnP9wtx/sUEkXf4+eEvgSVIV1ddv+d
jI+jF7BdhakeYYaLnm+PYwRtSbVC3P3sckKVYssoKre3+JzEOCCXBKJIROvaux9a
b19mysVtFP8fojFFGOWZaFy/Njg+d1pyNTg0uZB773x/MOqDLPwyypxP4Wk/7cSP
ux5Jl/s1GMDqQDaHo60MEMlRg/ps5QRhRF7Vm8u6Z2AhpJY4QbMaZC07dk5IEqQk
2n1bFhnUQRo2CJgE6/ufMIibsg5RSSWoFwAtTeeBPZJM3I2lIXiz3yuDM6D5VRKQ
hpZ7Vqe3e+SkX9XHAlp5xf5FUp6SnCacTN5FllMb9Hq54sOtTqPjPfroOhypxl1M
jDViu/iXnYTkpepsE1KE5FGq0VPt39mdCaQaU/omjcaXzgdPjRVwfL8cOLvU7Osu
n81o907+xV5Kq1bDe3l3d7vGKdXa2qljQcc4xxCkloiMlCAugp09/YMa2qWDMZNa
vpjN5ZWFiDxzDq03rH8VrK0+vQwquciVSz7keZ0WQWHkMc7Z3J+I8MFzfJDv8LrZ
Qj5PtAbUV9NivVo/11gnGgTnWPFu6mqc+he+IJxqBgZf3q2+vxtZMTb4AcfQIE0s
giNse7e+pSgxHHZ2rs0cEMRN5v0W5tU2vMTkkrrTORF/K8ftuIMjeWXukQuASZer
q4VNnJYJdiIrE4uI0O/4GydWaORFGXqnSYQFjYWjc7qB6k0DTK9tj53zVzRQW8et
FhQTxCE+7akIUjEKal1FhNoeVyrUg3j4qgJ3nRwKDhMf4litkeSvMexpRpn5PfzJ
T+ajcBqpZSD0csKyXrXzP8WSxNBWKfh4Ep9Y3IgmZek176MoUxDEKJD/m0sZHO9Y
ArB6kAxXGcUvGLpd6ljZqPdX4oq6YY2Hym8XJuq83E3YQouFogM/MgmsUvufs58V
AxPdmc5e7zLt7kZ0eCghlwUqjIMc9Yhs4XCaTwrhQThU9HJgaG+OMNgrphRuR1tm
Y+oAeNl/iOatomcC6mjMf3DJiI0JhpoI3MetsnaAa8ZCg3H8/fIBKUoEGe0wDaEA
kKD81oj5JbdFKnmIJFp0RmEr1liKN8QITEwqQtAVroi05wituCOfy2ju6/jSTtQr
axKQI3GILZ68rYG69TUASdfWP4AqRAhtJa/rXxKxW8GUBTggZaEtn8VPD/4iIyUc
FvhqOU+buR0s92kczO/86z4E0ql4cH4yduykRtJPdVAeHqBj3pkULvz0pFmrR5pI
8D+nclVSZYgowwf6fYCDuxoT5Y/W5x7jKpZf3khLqRbAlphOfS6uFQCRtj9fiyaS
Oiu1TMgtDtOnX2xKzUWkf+Xt/QAQeLgZITCijgp0Q35dQR+6FjQW9cyH0dfAImnQ
fszBQw3d5dOS+pPV1ElcPKAgrGgnNObsCbWHdyGUC+OwbryAl9HgjauByXhnNPiB
Js028mawD/KhHMXf6vtHKvdolbJoUzEuNUfXXK3EbuYBubW6K7VJT0iyYzlaYj3n
75zBQugyNwLmfVkJWFS84yBvxuIsoW0toZ7vVmSb+yD/La8voB/6Pt1SQb9g7kR+
WFgoFrPvPmPQMOrA4KOy4N5L/yt4xfrxpJuGU/d1aMtUwxYvMgmfmlqCdkTyW//3
KigRsY08iE6mBRXhEiusySzB+AqH1fGYt/uAsKDds6eBol83GdQ3IK8X2AAySW3J
jptGhxOz3gYTPCfx1XahWqtEosZxDr23Ou2VAgmi0MoBSIDvp7bDAjOjmQR/O6N+
STuI8XeTo4fuu7UdyjYK7X8YidaPKOvmMcN8nNtXsA1+znB3dkaAUTFkzTHIRw7z
JH+NeF2lWLl4CP4imjUu6qvX6x+613uBsD2iHzLYJQTwQiee7ce2IgAKrYPtaumb
tfsbMDDrJtDG5F8oed4n21pksJv9aaTxOg/pOB9mseP54hKOqQ/utKcpM48eYxSq
EUSBsUtltFPbHvaupyRbfqinDQvr/ffJRrCGoW1vY6ERXpAHSmRiunkK6POdH46M
TnsskNqADGXA9sQ6LYpq4sTcJ6xH8BSJTI0xGOtTiun8IVt2UMOn55xa5miiBAxx
8xlxpSDushqZi92WyUsz5r/8dzS/JGU+v5fZfc7TsHOuK8PMa9G6iRH5ixBUeDeW
EIuEhSP0VLTBSyRP6ZVc2Heu2CJ6ajEHRvMpwNcKfwokMx3L2VugkfevOuzA4rrx
/GGtuHvkhrmAiA6yoQLjceeQeRURcBZvKyugtkxlvfvaOvB/jGH5oyalxWLug9s4
mjlDJB1z1Ks4OjzWpJZrl9gA6cCSoaYaXKRwkabOiZ7p8tRt1tJxJuN+6Y5sobq/
Snj4GeoSe2/vgg6trIEbs1U41vRsLADX0+t+O+dTakOGNfTB96Fb9AqLANAKgdMQ
9wRr7bC3aWUq3vHVU7cPtX0bfgEl512sVTPG8inA9cwPlsyZPv+f2wzJQdS21qVY
a+km5/WptF9R7eXdIQh9WIn7BU3lWDHrE0J7Bhpj7VakLG0Wt+qB1X7tWhTLxcqB
nWhFSwuKNHevrZdYN/xYPAtHciggzarxtgPQm8dK2tZI2SyvCal8DRu2siaDdZuE
6Asyo7a3o7OTvJRcBGlOlNdD0eILEcOTnXa9JU2zZZk3oWwngeP1FtacloTFRAk4
STYu1YYJn/28V7/k+7z5WAt4ZX9c2AcI/yuCeTj2wRzvJQrxq9y7O3gFeqTUDZZ+
3bla4N689z6/cAKgf3036A7Kk4xpsdVOjfuUWJzV5Oy6bFVYyZxGAmgi5LhHJaaw
GvZ1NiePZJ0/mnc/xHpxNy7+GwaEugUMTWEY+ljQEdbSVtWjvvYzaSXX5G+PahF6
XX1jKYmfGW9gP0oDfHdVe6Drvpck2aUeSoRrLB1plKyH4bjU23zyTs/5SB5IBSTh
PTx8Fc1WJkLR/iXbqW4kF47Nw2DfiuoYqpO647NXIbuN1rgXxD6XBElGk1deSgpJ
fQhb11D5c0Vl0CXZez993igNJHWVnbx1j3Jssapbxj63jcsAmiS3jdOxP4O1u+yw
tc5y0REg/xs9kYA931/yfSg7y+IOsHSwM7sLn8YzwAU23xbg1OQlp1sFQk91/yKh
oKYDRthDIavBsHe450E3OV2EtAtvVX6gqBPAJ2pzPKW9L9kci8+ZDsyeIbgETp1M
OvRyRHme8CQNacEC8nlgKps9Gc10MVrxQ03oGy/OAPuNgsvk/h7zZ44WHevPgB2E
/Bhn9exaV7P1dF+aLX8f2EXFVE/pgk/MEaLt+uCUuHQDQsqISFEnyBXm0EwWEjTP
OEyQnaE9v7bflruhlvE+RVck4Nb4wk/zLCr6nkkI5lg+S4i1ZK3UGpi8AlaUSBRz
+KLky9nlMc1GP694E50XT6/uUkLmsPKMZ1QVIYY8/w9AiTcg+/0nafd8ns09a8nW
J954x0VnE9USEBZJC8FkrJBi7pwKwSCCdNYvmO3WLjx3jmaGubLmuVcUqK+UlnUc
9r0+Nr9GNSRBDE4eTeO7x+hYVLQMHxwBPSoYdXws6nPskM3H1iGQ39Us+HJe8Rt2
RtoV9R97NflA4g2c4RnB+ERZDynQVI8vq+nnsjIlbjfICNh9FsDbtqtexvkUtsbK
+FRD2btoKhU9XbLSYVmWX9hNOV/DYAEryCk0BQ2BGCvaVqP3V4vSM7aKuIsfnaMM
sV7TAcY8nfnju7wtcU3lp1f08eF4V705Q2T2X6mBmvvgTC/pE+Q72oia7uxLDw5K
pIdajWnogQ1kSo+xCbiL0fTwHvBFa/QzREXL2cvUiA/ac21WFX3HrIfXHJ93FqeZ
BZfrj9Dhi7y/0HM64b91eFsXB8CTduTjnOdv8qvfbKpbfWH3x7NdXwrwvHBC0pG2
bIq6cZ+b8uy2JLTkWRCRgSKLenQhoKp84hgYQjHqzcpuCKR4yT8rV2WOREXRLpx4
r7TTD9DAUi3OQZs8px55sD+GJWfvTAGPENHu20qoFeLOa52FhWKNeZS13sQ8hzgM
6F4jtU0KvArcx+ZBut/EYc8gqilxNVhiz4b9DJMlRhZr5hAztZ+fY/TTyT59rfy6
0d2FAE8cojREQ23a0WaU6hlI7CpEcSleIs+dVF5pmwAOyTiTsxvjDdfMQepyJG9j
jEkc4a5n4S3uznd/5U38HpT4qoOfmLdiiCzOTkHH5WnmSXf/YDGFS8hUhRz7kxjq
VMoYeEEmXSrLvzRSdBdnczQV05yui3RGmoCF9HfAsw7w29apJUHNTCkEl9NREC73
0ugKuBUC7vCptVcgPLaL5gJK8HMDQ3hAnURXMThvvrR6eKyEyE/uQNvy+g5i0f8E
m1ZqwL+JXV3GA9Ih5s19mZSkS0sunbwIIrI79QLW//QNpEqWVm1VeAzGbwijX6Wq
T3bURPQogruyYqHkDqxIt8H2ic1q0hKDfWA6nthsTLeTfm/xWwIA6unPN03GJQVm
UQb4lWS6bZWNddrk0+StBQTzQwPQlo3hSNohU0XpwCxVe/mUZ9N9ORNHIUftFMsb
cn5NP8t4j8kTB+F4uNCS9/2D2SxecGj+0CkLsi7IIZstEk3h7UFOXz/PVOSyTwo3
Fxj37Qsi2mDSz6cSjCk/MHdbj9nNJnCjK4xoRB6M2vrP2SFy0xiwA6TAISwnf4o1
uCjbG/aDbNU8zKvGwOuTkMvHIX+W7H3pZ/CjHXVeAxhKh0EzlP10i0EekwqVdKUp
NtZaGppk5S4LmjS07HvkkP9WzyuDOoYtAWANz/dkecl/+92FJ6xhGtfa1PUq27ha
Mr2whPrpJ3Ad12czU32r3p91Q0R+VqhNFFCNU+mxJ/GRS3ZJ9c9cCXrA0aYkgAfm
SzaatM3Z2vWxEJ/i4VElVTLPkRsF+svGW62SvXQ6ccvzGUbP4581xyarRXnFot5n
sEjvLAxNV0YCSIMtMAg04faMrOA78PJ3QxINMSH8Flb930kxQUJwAMmsiZllMgq6
fPR/6R3/Y8cysCBm7U6UK0mQ7zPVYRBksYmCZjVQ9ycwc2+rQvyUl+njYXL+XNNI
pLHRJddFY+kAU+MPryTCE9CM4RxWeGdwxc2h1WdoarzTJidGvtNOuFxLfs/naf7F
50vkFhsKP2hl9pCGNnGunjByFUv6iUZTnnKLjn9CQRj3I6JGOz7jUh2aDvDGYwLf
fLfXkNlwrY97obNhryizDS2ZLMfqlmupd43AyDQl90BtEnL9+tSlqhs4ooJv1uLo
GF9e8eubyQllWk1tprIwUJmoDm7ed00M5C1noApXPKq3YCLJuUsgRj/KZ3MiYsjf
/HxsJheXmAi3kuJKv7YBSvEhn/7+WeYm4ElZxSWSKmCiA++8slP1CdLmFr1GljC1
814mU0StY8M0HmpoVjP3/ryOV8b/kF1LNhcV0HjK/jICckLYANnLYH3hIZs7gTIW
TnagElOpLjDAvbuSXi1CErICC8LbWScYDbpZcgze1k4q/e6z7CP6SLh4B/Iwtwmk
Pxk4qPTWz548+c7RAPCwVci0Sd8NartwUErjQybdBVvJC0iMAbkwkQ/mgdfRW9/r
BsjLXzvcRUzDw0VToqvtlP86LcdQQnp3fOqPAhJGd+XnpC0Ce4Y02d+0FHKOyaFn
E51IC3/zio1UrNFdDOPXvLJmP8A+Tu35zldBLrRgEiimsZaEh6grlwjjDR7kS4oT
KsLKDC+rnlshvoisW5OozmZIW2qA1cQBjtqTGfH1fvKDWbsqxBuNq2NuZHdgNZlX
v9C8qNbR7VT2WvPH40Ea8qnkK0F9c2NAIHJ5TAWHVcjoM3u7j1PJz4FTCvnszc34
BtL9jeWrU8uI3rO6RMCaR88y9YrTpKHptxvKdN+T9y7B5VyQP+sTGeW30hpLKWAr
uhjPKKzYdpl2GkwCLPNM8jfPBotkTAajAAJsGfUEbjkRGuvoPyFeakzMsegO6fF0
ihslUA2PXOwCQo4kWP3pggxWjyiwMs3mSdAzEfbhqhr4I9pbwns1DWsMiMLufQVr
FZHpMR+2cT1AfSNuljUiMs+229yka/f9GJfpGgrdSwFsB7hwKj/K/uUI2Zeudy2R
q0bfXSY9nldFDARPd6FWmj7yH+0xQHEnl5xEbDf9YrDbzy+MAO8mVF3oJkm0mFwF
dWjXq36YNsVSQiGMpWuPk4fxk5WgG2LMNUvXQHr2qIjSkYC/5s8AKn+fxh0nPe6Y
vMvrEzh6UrWQDGMatrWhhvhsEEbqHzd08A2XZY9LtJySMeksQtOFrs2TH4U++fyB
ARmFdqz/cqkWieyFVdSJyEi3ul8ZRld6oMVcmYbzcNHv5FVM3iZMDGChhR41ievD
M5OoI58mV6eFyyDgkY8SgfvG8aqtt/RIy3yRnHwxP1KuDWt8dsaDW3Mo4p7ogmad
/ul/0w2IO24CCxYeO4zjkOADZYgIbSGMHBuW2FZcoaC+zxdgWwnNthVPIrZVjwcf
rfXI5g50MAksGS4D0uMrUZFpyp6Ve0H+oEoJNqUti2TI0g0a6DvlupO9ivOJpite
DIFLrjhdcaxcYTVXq4cxtabFNc4uJFujUGQBwL5tBPkHGsS+HecahI74Ct0hALjY
ttEklVouNKm+DAL9H2o7ZI5thSHZIHQS98qDKKzwe4GV+plKPqRzZVeezOKVYsu7
xzxlUchK0MXwHc3DXfG0Rz9naR38PVhf5C9xFFXibbnvHh256yNftaKd1x+gb45h
qc8+zf2xbCgSJhco/hPm7LytKSzzzr5OxSDu5YuXuTi5Q/hEEvm4Fwz9ys1SwvDw
4iN5Jj50OVENOJXQRS646CUtZGTRRqOuIIkgK5zlgjWRIeUOoK4E+bNIM/Z/gShw
pXotJo85U+FB2dzkF9j7zBhj/KI6tXOQcflL0paoSU8oM25gFZlCA3Iab3SVhsB3
Ayl9K+pNU3bagcfLhHb2Fa9a3pL2d/sL4X9Tt0MwvXA/+4voGXsYovr0Hgxsgpq/
zy77FTd/yrGZmss/qPMNniGTQca68OkeDO9rmSStLDLmWf2ygevWrR3xXUxNZz24
f7iqcvOY/WN4fF2x+2E6ysbj/nPs6Nli+gD6XBtekeGlrBY6+d0xad/2nCd2Vu4f
iWfd9VrGB6pLHfMxwMO/DrSLDjN5y3/aaDuTEgp8G4Xnl+ww33OesfKEFpRuQ/AL
AP6B09bvAjaGqRiUZA6Udu/+6KG8l1mVOS8K1Lzp+GpKtFp4BAx5fCnjviKpf8Ua
lFwqDcky3zBUTraGlito5guYu2H9zxvkqydWmuIQmn3/U3qUZ3NylOuZnd9VhLuD
rYjdp3v7k3M2Qr57zVSMrTKjwJ9al74t5nXq+NQQs5ZOGoS/0XBhcl2OH8wiNOEK
GKCYAoYZ+QrIqzgVZcnwBav+lhMfUNtIh2Z9plXk4zdJxlE688aEYDC/2dA9dsdQ
P6dt27lvRyms/bSxWSm1xlrFiXeXBGjjiNWRpfpT7wYbtcNQTXEJCth0bLb8KHWL
mF5MDBrgPZgP4qJRSqCzbiRU2nYR6Tiu5Ge/3PsQlmqWZHmJOHd/FglmmeqJHEZX
xq7gkCM9dZ8k21wUtcfDT8b3hMGtY6rNoRVwb2wVeC2HN0in32VERGN1oWbc/Je1
qTJJjYEG4GWOjWrbqz/0S2BrjiBIcZXSlST4TEY4GvPYJ0IFIsoQ5weHYmc0STOQ
3RjN22PS1/Uty1W7yMGa4X3sHWk4oenNdnBaTr3pKS0SqZnt5pOwQro79/5K6mgD
4d2IESlWx9QhNsWsKYtxdhN1n2RdcDUSFbRJDDKfCOqKkem5xncFpKeOvCEG3kON
rKOAM3SEKscGklCnBtspyTK3+mHNL06EZ3v77S+HkNY4CzEgvOpiOSv1W/bAa0+n
sinZB1cYnnse4AsPh6kRpKxp4HjtX16e0M8KaUKbu0LHiJMNrn8QrtsTJ+ErUcEx
glFao5BlLsGKNGINugsiRTCC68T8a35t44LQO5e6fkiFPodGbQ3ppOgjCAqt1Ucr
fd29Q22nlq/te9IiVxBecpxVdo684wzVoF98OL9WdOhkORlugqQbDmj3ZH6q5OwN
3GovZo60fHniOl/ig6b/67KFIQD2mKFZoHpTGIAzQAjEiIUJiz/sUqcl67Zfje34
ROPgsCt/lYz3YQ+tQjidCc8Y81OeQLMwmXOaRzgrehz/xjUwV1+UQ5nQNQCQ3d8j
6GBTodAZecQjuXxpAjJ4+5jxJgPQt5ulT1H/GR1l3UvcVNZHKm/Yae7l7HRoVkgV
PTrT+WcV0ne043VDG98N7B0MCTLw9YhQINlxc1xD9QaQ9Yxi8UIDh7lIuVVZTdj+
AaRrIqzPe4fbEnvVI21hvgzPaJiF6PuRuGd/V5zJMU1k9NxHAs9WzHiK0GpUenUR
EHEFACJpqGw8mhwRjCLxJ/p0v9VqWOjbgZetSSZR0bNQ+dAd2sAdsf3XhbDDbGQ8
CdBMRNGkXfmz22FXtsMlCra22VF6JLKv0Xq5rSx3DTUo8JgT+6pS9lPQNaFkZJ0S
c6dW/MB0oB8DPIn7m1pPE6+XhDZc6ZVj4/sf78IgpddA7mJk4J5N6bQCJAN4NX09
bQtGzj1jHFODBDwj+ZxFEYQ4eMWZ/uPeUJT6uls4PUXNBKW5Q4jyrEGRXQsMN5Zy
Amr2JxCG02jdet/T/03UpLC22iSYSo1OLZIoRoLzUI46FcI4TzwgTF8bhb5ytYoB
33+HSOXbYKHkDYK/fFTWI2n5Ax0X1ObCF35mXkvQ+m9VmvID06pOBKdzeI0gATkD
IejsT1kb55QEpeosnt4UAkUpk424UBhC6luQEpdnxunY7kJSUX3Mrc09UOzSR7N3
zqn0m8muCIUfsi7EWBnumuDO67O5Dqx6k4QEhqIHDUGwPSEPyVg8rE4UuY9t2P0R
mPM4E0c7FRbtumtDJSRPkW8+Ry1XU3Kj4/519w3CPLfnuRbeHPD+/1Vjlh7+sQ4i
7lGcFjZcV/huFD4bBsyvg6h2Fg0RWdw5hzNDimTcBJuYRcjVWOXq7edDpQU+C1UE
8H25a5TbzNEHN8CO3TMF8lFNvZ2bnH80XxYvaGJziTvAnl/vZUOR2g9imvcicjGh
RSYkmF21Fhco6aJEyq4nFoy5Ld9GUmR2g3s6uJjXAOw5Gw+3/AO20m4H/IkAaCJm
TCVIRcrf2xGQKid/HVD43x7mTV+RkAuCfw1doulyTmpTNvUDHrDCjaeq4Kl1eVti
NzGg7I/rt7rzPJYAFClkRwG8XujjAPwT2VNHiL9/NGy+lck4l+s7dnd5IdTKXvlB
FyfhSM2AA8YUut4a8Okn851tG3jHLqIVgpCJnLlTcvvrIVgyJwJHMCiFXQumoDC1
cfzl7127m4QhLEPHKRDcqP35S95wMVt2H/YSbK8x9IadmA67lP7DCGuXlvo0B/2s
Bu3z58h6X3gSuT5EUUMnuX5MkZHPzfJo36MKxiLprn/boUDH6ECCDrbPyY3mSeoL
k5tTVQEcj/d36geGGdSG4CPdkYAgt+VK5rCskmyzM91lgcU73zfFAZYAgMXZow1+
McAWFU3mBXR5vJ3sjYy1vupa9NeEkmjT1RySy0BynB8ioGFjA/yBAPloqDRcKpOF
2DJluTova+ZoJmynWHWJrVbtXpmsOcgYDX2jD0sax1T3d6+Q4nU3HdVs2XK1tauA
gGyUVXYF/PqfBndRaPgJ/H3ZamYxNlEig+MGmElNTU7rg85WV/9Qht8YDKEZqI7o
Vng5N4ODiSLxV6NiNUMK/0nQLNQgiFPanWDurau3eEncAa9CaHzTZhuPpiLhx9Z6
BOEz0A5Q+WqjUPFUjUuj9+xjXX6AKWYNccw5cIQokz9Z7sZzplr7vwrVS2zPrKAU
nBWLvzp9DE58A1RxkeWg6GTV0ql8E0vp+tS0GJvcOiu6Dsq3YoADnNIlAMc1K3By
yi+3Ri40XgycD6u1ZiriBFLqraoRsr++vsibPwSu2NiBj2d4Bygr5k1NVbgE5bok
eD4yi8oK+VpNV5NYLh753BbBzV4QanaxeR0Hm+iosu8R9OOLZN+Q1HJ9mJEFsVOM
mt413yunUTSrYTlivNs2HQA26QcIA1gmEChNFwUwLlfUI6b1xDtemYAYnd3yski5
FBXi8gOHK5B+Rt5Y0LXRVBWYLhhrAWaGGStEWMxwKbtIFeIvxJQQNSJGEvzDhoOK
QK3z9Q5koAuv2mEbkEvo45uiV1INX6NAnTHSXcXXHLm92TmmaHbkyg/KHhG2OBKs
1/WIcREFG1d8PFlOfHQlTTqrjbx9hJksKAaSsT7O9JimbD8awzRoyaiOhCWZqAVr
WQw7i7M9rYkfpF/XhMjC/EKCYPm+ukkBZ8c/+09QnkEGKLmm4b0ScOiF9LIuu93Y
ji9nbWip/mbUEC5KS8PBbaB+YemxM1H5ypYjebccWCUz7M/VD0YfHZ1B1eYvh2SL
F1S4iZtqU5luzUy0KLWmcBKGAfudRb+WWEvty3ITxY/J2mfILBJbpJgnxEsuFWl8
gDvzcSpJyuQCfG9hN2w1baRzJ1X5QJ05z+ZEO2wPGHzFIxzr9YVzhAm5ookzlAKz
N4F/JuUxtfIbDgDrq7ZVUzeXWbv7XqooL93hYZE3lXIsNpARtF8UJVsJVViMt9tB
j4ftbcixddB8i+Zg7vaoC3AzdC77m6oAvfKqUxTxanohutsgJRKiB5JpE5jeWPxs
QAhl6U5kFkBZhcH4HoAIuYMZACXG4RBSaxW0F/nyPhHieJpLaDHHTtk65awVPyT6
NvVsx+luioXRK5Fwgt2R3WK/LQtg9wPbRD12/25KH4vNxwqneMmxfMdMcgWz5FpU
MtNJ/NK/tTgr9sTaqsK83ZMhZtBBjB+XHB+R7fbX+CEOvg7ZnAjz5kUi/34EO5LS
w3ycAm8dGbTv40qnEYSDG7qoEQ0SpbUERNTCPl7G+bNndegUI6kzf+aG1kmAIY/s
TYUQtWPkM8FDQOkyxwmY7NKzMtHn/XhWUran8CcvGrQz9RtY5MeSpKAF6mkzo+6o
ehK+ne+IxdQagNHjl4tMhD4uqSm6t6o55QjqOM9L6aZa1lTnTEx8RZn1EE1A5rVs
U1KvpPVOaJTwwQyFH42KddRpuOyKKQVRhfLzJxSaQFeZLdqY58Pw/N3T42uFWQWU
CVNIadAmIeBX2yFThg5EtbE5bpNvufUXB+MuS93wLrgHablPdQjpPd+qifyRx1Xq
I+45hYTWjLOb3KAUDTz+4O8S09RykJL9loexPsCpv9huZ6wDlEDXGPuWmEG/IyTr
aEAdzLpmReK/bCQd7iyYiBUEukY3GlDbKXDwUUgZK7M0tbLQg1glf1BCLmL+VJAD
SAddpUovfRgeM6RvGyUhK3duozA30xU4b/+QlO7H1JdsQMaJPPchL5oUzEhz2ll0
XEQi103IBh3RH76FtMq1+dWYKwLU4xmNZkBdEMa/7ViJ9HBBfzeJYy5ADkJVhtsb
EXFe6sKJQ/2cHX7dF5Xf5upOgHA5ci62Au7gn5J1pVYrVQFXcDdAvXO7guDDc8LG
ZJ2oJSUaKhNEOvf6ig/zKz/Vhpe0eTesw2ZSCU0AuWdOzx3zJr2+3BBMUgYaVH4I
DmsUWY/0HqNqUQfCU7dyFCvX+L/SZ4ZMb4ncH3mPP3ko4wjz22qIteaOtjDYEgY1
QXejaDcgYVEXfJ5rp1c14XEEe+G4oYXVdZZCky76rVpEBEd8mmy/loZNPlcLwPOe
s4VqICkpyZmQQNEp9tJqDkku+fEef11G1WEatqKRp98/g9QaGt/u/RiK5Bv3RLMX
35eEVaD1EUTxIcmc1k+/dgmQkxH099HwXYqd6OMWmnsqD4pIC2zt9Y0YEq9OcqyZ
XcZdOhBgYVG/VzOXjPCWRnJDzET1HBMY7pyJgnP6pSlmi3LsrRG8TfShCih4dZAI
ik/gs0ZRcSdVligCLiW4xCvze7L6paWoAZAGy6MiQfWsjjxGEqwf8tRAMrShlsk7
nCZV0IRoWGwmQfGKhX5YgX8xxiC/8kQLshSwIUcJAurCnQZ7xqunZR4tqcafXuaI
TQzbtUgPxYVkk2GZ96i4x1erVFlt/JCE1YehUy6XLLdtzXTusTI6TeJxR5vcx055
QNF2GEilR2nymtUC7THKz5OYFOOSu1aFNkIl9WxeAr2K8RetlmcT6xi98342CJrV
GmBL/756mJkwdd/NP+u7XH+BCLNFgZ6Nz0Jzvx/0kRMdeh6sbqY7r9ylm+DZbC7G
TZHt1zuKIDWFZO8timLpUGWtkqcQ3gKJm1t4Uvp50axXWFFzeRA4laRVP6HKjIqi
O2uoxTM4fvsVo0FTxlIgGHAeJNDAX1ESvHGfnH5FkkH50JZmsoXsE3lTmwMC7KF0
t9oYQZwpoiuIHRsqIn5QJ2X4KBOXYJPBOlgSP4MduC0lf9rReizp0B4uHwm/90SH
uPoZDXrQa6vqOWIA6GvkovN1/6dW9FjDwEdnlyKFTnWZWhrpVl+lpOep31/8eC1R
CXD3VJXq3P1UjmBkB8Hc8YeifWJiVF9pJ6i3yRZUf7O+ijUIKjdp0CsfK/Z2pm53
u4t3jYkZBNWlQAUkFYH7QVejdELLQQww3qqIpD8QoVn0v7pspQSy7bfVYIVxSc5F
B0OTtsl8jcXlXY5s/lThcMoTWv7fNnV0UAMp07nyBHeKzBxXYEK/yINysYlJFXjm
lm3cdfQxwYFj35kgl5H4+IJhSoHCsTU0wpUwcnTOni7vxKOKSE04N1/KkYsuA+Kg
SA5m335MnlFNdtK5POzdoZ+B4cPN3RZnf4j7GELYpnkm4QfWY85k+0a45na9z2Az
cT9eb4PrO8xVYK0ld3590rxF9tssyw9/pxt4mwFVcy5erUWLxTfo4//VVa5WvhS7
eHsHWnM3/bnsIV+3sR4ZyofFQQsli2cbcYkqoEhl3++VvANQbsIni755qTNij6SF
8Cuhnv7lZmTlsmjXPL7mlYK7NZf/cBIZ7EACuIm6CvxSuU07cv61dVjzJIsp6WZ1
1i0INcT2d1oFPwDdligLMoG5/hrH0A+l/7TH8SpsNfq2Broi2a8qEBhhDwrlda1U
SnMeyaGY9yz85QxNC7NSbe4cAKYT4k+MkCdfbDc7jjyQ/0Ucu2ywV3Hr5L2iZgq7
D+Dhdegr6OG2k9ErGKtq4KY5epVQGJLe01UtEdPbeHgnnzMi+Faqm0jAWHhSeSpw
gDaTbYNAn4vHWHu5vbb90PmWeVim+W1SeNpnSAUGMwCd3YsjrYq8qkQahZZ4pem5
yfFPXYlGFkx7HvFBLBgNLAQZIVrh6nJKHuiS5sD+ExMoxwi65zu5M1ZXy53so4zm
QJhGhPGgr4weMMXhs+1gjDXljE2RF5IS7VowQ8ezd6JVbd8jWY9X+AI4sFpiS6E8
5lOCSF97jlJDOXWSOl/XCgPLymg7SGFZS/RsPVwOUyZ6PePtk/clIcxWjLYsgl9m
WuLetdCkSv8jGEceKe2WS7WntFFjeZ6/troe7LRKvQNeFZN6YWHh2l5AzpzXIwLR
Pbslk8HkPTKVZdleublpXNW9pWxlDaszM8maRSypgKPKjki8XyyIxFOt60wUCu64
hYJD0qOBMZ+JC+D457Gr2gETvlb7wC1CzLMo5+k92pCF/JxbCNvbr6DqfyMfiSRM
IdHxzoc6ctr/Gl7edYUur/R+bFPtrstCNOvAwkVdUPs3jDwkFB8K08lXIbQrEo/2
1qgiInpd4CLMFsJ0rBRVXAhU3zLNRTZTImxfF2uJDFtztt9swDTaFqjIvJQ/HC+O
rusHq93E8uVFSfH6sotJdfdw/zqOdffDBCIZoskYcJUHMm6WhFWUP6MyrKGYAzvr
OG6iu9h9RMUOUOE37SAhsSQL1Auz7dxWuj4hQDqOxnFrszsnCjQaqC17A25UjgHA
S6dLI4AkFM1CuPc5LnziMWp59QXnEtkGIru4PzzQc1IERlAONlQkQhVIm7A1ql+u
jYe8eoXe+Nqv3EMcq6vnAShus46K2n1XCRFLzRFRi1WQisP+sP0q1YOJRn5VLWa4
X9hjhNnwVhP31Kr74AjVl+oO7gucVh8c47JV3rtvEqIbC88zHrBxB8EACy7sGzAJ
4j12o7whFbWuV2BpR64eB+On7CHyrPIH+DIlwJYDP7s79BdLR9YE8HSxcMd4LvOG
io7rAK22qc3CZA/Esy8Af0DcmDRicG22s1QSEB5qbfzYZvQ2UYRzAHdRs/uuacHy
CxbgkwDuZ0jUGieAcGR80aK8li3/9ZcCppmj0CsHsLyn0gQgVNw9vjHj91c3vZ3E
KqzgRtp5d+9eZ5VpNVE3mX8mmxje3+KC2xZrYku5nrMXfRthh5N2wsvPLzePBM6b
Db/jbhLfXfI5x7BqAnxMnu+CaahJYbqD6V3W6g1YI11MqWkjmeGyD7jFpWcgquZv
vMfpAZjwGt7+rK63SmP9T1LuDeEX3Sj15f3lPwOWAravOgQsEhy2D4ci7Ncp9++z
sFIHXgHcpsVFXELYjWxtKiGZ0PFiRbJONb4VOXTtSiUxl8OyY+pjaXXsyA7QKBDB
2MW7wKSBcGLq1yxaQ2Zy+hYbXiIgtGmlyvN9F/zZBDbkJw4XlB+OZp8Gn6mSzYhI
TxXsPupPhMDf5cjNMN6SNFa7K18Bj+om5c26HiTkBGUbymmd4yaaVRMzbIFjD2jo
5+Anx8CvmiWrTLXCBJYTDLMc/79aZZLMzf4grHNGDW0sdt6MnwiZghbwc9ENNgBO
s03X9ji/GMrhQd3h//0nBrmO4SksBM0bCw8kY13Wjdr0TdBvOK5Q/XIC0qCLKDz9
fKFSfcU0NXjZr3tBkPC5kcbXmHtCxRQwCVfx5YcdLR5MwVKkuhkpmhCShH2ShfFk
ybK6cIvEaoASN3KXsdUgPk0YFgj+ULAaivf2d8+kbakWF/jhLmzV0RIin0UjCmC5
TyYdNRGUvOgOD3jmRB7G3ABuYDdKqiHD+n8QbWAYAnSVBsU7z9pOcxSYcHn9zpD5
cN+796WK+aUkZ4V0umKCSPPREPdfGYetarTWTASCDCrzUZzgjkwtCEHT3yqyUCh3
6OBJ+mtMBBw5oaJHRYQw8yks7pF5zZAFHT8KUbfbb7zqX5dW+pB9OMXFN8+l2I3T
GL7U5hVQ/p12CMmVm11XNzh48hTzLlenv17mhuuAMJVhP68zwVVgjU7tSOc+ioFd
9aDYBvQ3DrsN9iJZerTtux+zKgJM7lzXzrAvDq2lqx4w8BnFN2KM3/GPAapBYke8
s4fDySNRP+Vpdm03iPruQchIXWHlQc+9X6/vb5HBNUWcXm0pJ1MTqAiV/0pPpyPs
jISu3ifhGgaanmGh50FW+MptH6CZx1n05wy+eXpJBSfL3d+7R4REzuWZM3TQNHMn
yrInuHj/o7iObdvvWo4/Ou9o51gSewhXMxdPD9KkSElseaGhJDM0v+qfmOSazw9H
qgakUlcVwSEmgQWqJ+MsRQSY+vQg9VqMUothgqlo54cS7AmUzRjvQxWECPSngEn+
LHhAvGyv8yXO86YZoRQQMwZT2xbCX0B7BouWwTJ83z5IwwswborJJWjQy65rIF5v
9mYO80s347CMJ1LJehpWL+MeYI88XUbOoTL1d8rz8DLGzbTc5qeegLNWxiDuzMLx
Xj911eSwQK9q+GqTbfFJCIpclNlWdKQpNqVV7MwK0C/2GkF8zzXl9oyVNk4RCMj4
mW48Arhq1hRdBN4mjZSz6Gmd5Xnhh0R8P7JlFSwIG8PMNc1H/mIrtmPDVIaAgggp
mn8a3vSAXThvEJskzQJ2WHgeefm3dUuuav7OvAW7blGEmE4/SzotZdWR37C2u0QN
BTebhmmgUTk5BfSH22rgu6LdDyyaNvTruR0D9YbxOSneEs75RUK25QEjKCdjV+jM
uXcyY4+4byCa9zYSJnbOXGIoKJODNCK5CQTIujIu+506/X69nbWgQOrZA2afuSaA
lHqePfwjgWvofACo9CGb5NYiFqLkfTyR3rHPvsRdCgXsFMJmhDPYEhy+21AUUUCE
hDiwpIO6MRW0X0vtuOlXMMk8RqRO+8eOmuCllrYIsNQm0bXoH7FI27rhDC35Yh5h
MxdrmiPEY00crz/AZ/E9DVPVQ4A2+lIUI//IQKU1wctzR2K+DsftOMxxfd/yDqXC
s47RdLMFrnadJbjC4aYKKbSNYVGmi2yUprIrIhsWf3yc5WmZOpcEFYBDE8RoYAoF
5bjGjFxWq02J9au8yuWf3NitM/D/jhE5DL6QBpxnBd3tiXkTJ96QMheMn8Kqmi0x
woVE89lbORfouZalTXAn77DrCpAMyMbWdAezYmVZQtSqTUaU9xl/SGCtqSJrJ5Az
20rjylAiXdfnYU4qg2cKurMk2qorr8qeIaNZSH63YkwKyACOO5gKEJ4PEYEMQeP6
XJ/FofQfornS21LFl6OhhCzs1tZ4N0SPdH0+jfOw6f56XTc7od7Jlp9optGccIhu
K7O1PBuOMjiunziWxZRNQWkZVC6KH3VAF9Fx2DA+xU3XYG+2vLdKabgv8NYGjutU
hFq+CQII9rpV4U8nzyu8A7vMAYnDWneKnedaG2Z3xXQcV3aCmVqquIS+a3IYJg6e
c0hzI1Ij9nsS65BtXH1ooe/FhCRYrbF8ezoIxTxNanheRzc4fevGkotOMRYsTe40
Znk20yUkt7yCviXRm7lm9P9miO43UZES5j8rnv76Xd4x/8RNiQ5O8uPDR+0rVtoA
2e2U+R/23v4FO1EuS3pZuVidsGdPLvlQmr9avs1sTv3oOecDZI13wkD035OTALHo
ygxvvfbnCPzoD/se647c4mtC69X04GzhfpqjeZB77aU5zXJhg0RSM4FWoCLyXHxq
qteOKEtXn7+Gy7wVI1zjm4p7hbAwoFMpAgYFECVoiYb31fOD4aPnAZgk//Ra66Y9
qFU5IMhsVzpWM6mrKunLoW9CFWDXl8PD/HYIO0BT9kRHb2IVNOupLNwZQWfvV+ZA
f6CVVcCoKc46esqa7wfmIRANCviXYlStc7CCtawVV5azzlMwgCL86jiGeOY6zBmS
B0wWd7UlIPPYSXbPmjBmlEf9OUETZJktbb5pOngKhQq9gGm03m4B+ulO97KJ3XTM
AGwyGeVTkWH9mGdJ8I0qsjhrE61euzrts+EW7OJHIt7fGfoUlsqpX5zXbLfkyL3U
si+vczEkUlGIWADsRuKo+dnHAZ9Qr+TYraND+FUZNjoz925N3OeRPCLFOVj/ob1n
v5Lv9V5Mss18nR4ZQpP83TRuMlc2vg4O3+fNUyXSo0SLinI6fwiISJVjQMG4hX1r
GD9/Q4Q4nmqU9Gttobx6E6Q7Af6F5rLvp4+dhYkqqDwZgGEzP/9TOIoVjKNKuwvx
xBJ1PIVvuSZefkYwKHpayaGuXI4x7aF2j+JFE/hGg13iSIK0NVhsMRrsCUZQBYUF
LqMOKfiV9BMP/mp4sZqBM/BPeQ2ThR+C6BOWOXft7fLjT527lxq5yzvQPNj4VNCl
XTEaG09TaKF4HFBiYE2hfqVs3kQpt4k8deAn/RH7E5xIUerJ2U6CG69fg1B1mUTL
B8bpeYb95D+52UupC+Vg1PITZx67jqpqL4N8lAPTdQa+8yc0+ywRv4ORKr8C6U4Z
uVlsYAbXTnJUe6PnGTfUA3fDPo+jNBnm1ZzRFJ/Pd0TTharwPklrZczpXMvJLVgs
J0hMRdKMBSxic5+RRlr7Y9P4B/AQAWMINxN455chg+0a1lgipO9wrQgzpd7ASYyT
QomJNKxZ3f0tnHtk0S6KFvacntPjJwCQ6FA6EZPYkU30J/ACtqi20Qp/DcQb3e0t
ZQv9CaVAFq+QXGQxczM77X2B0QCrTD+IA8jI6ci7BNCXjMXAWSACG/W01ssCTgSF
G2tQzkIdzr06v/xtCjKnLHirGCY72isUp0YWKOoCXyXp1qXQuEda0QVC8m+sOZ+0
i17GwNBrXxVBdt0rZJknkTadxpTqaUJwryuLulQVGu4zRkU3Sh5C6OEXFlGrRqcW
Pdev1p+KzSifsOLcOZ+qjmiFtUc/kzQpIYgh6KqB1RbOUUwKM7JXnS30ahxuJqSq
4Oau8K9tSw72aekdB4R7GDS/cH2z4UzzwFYebZFepSNn4j33HSO4vAEAS0K8jaMh
+P6TMPpTYZknzq0uuDvTDQ1ZGI4IfZKVsYAcrZw24+HoFDDq3mVA6TEzQU2ph8DC
08u/ElzC+od/u4c8VnuxErnObaz/I+jGSaO5EJhoXzlVasULF/HqERNwxNZKo5O7
qLu7tyA0W7SjEYWvlMAZ69veW4dkW92tZJyqG5QlZAHtLei9/runqZ7TeOOrXZJj
ImfNYTUhepwjq8IZS3Vy2UU54xu9DDzTEWNXYyrcROFA5VmiRkkLtdN7HzU07oGr
ibJ1C5ytD9PuOoZ1kLepNAubGPxcGqCx6gBj+O3f143tIlGAqJVyWxSUryZz3fNi
YNxtDN3rHIpbeyogcrjCvu/Xx2jZvUp6ZazHn+mFv96SLvBNP5/HhXk16RHefSdF
c3rxsNxJEloRdJGTX1iX3N+GuIe5w+QYhJY0o1LUjXf0oI/K7nU/Y3du9Ln2u4S0
usBXywD3Ye5qz3574qRqTYoqRxftlkt+2V6HSnbvYymwqyvVZILtJ98twO9Py727
GsJ55zJJF76h2XwKl1UGeeIxxgd1k2DUj8BKQOztjhnimtNIq5rM6GtDiYQCoz3X
L/wNXg20yQ8jt8JIc1Tsl+V3LaQeY0oACzbgvHT2PWJjZxqMw2MX0D5wogRqPNml
44DlVV11xNyZEUp0OV1gJ4h8EdCdeaXRnXKEO1XmgtpABAigHDeUX6vPfynf149e
4X1KC5FfUOFLO4KaJqVhRzWqvNthE9/IzQ4CJ8ayyd7tGms9SO9V+DT+v8CLfShB
ItmcrXy3SYb5f3qH7RXnqutEMSD9/QOXnGsNJHqo2E8X0TaKZTKGZZu9dsN+zQ9F
E4JkFZ+GKIwqiO6piWQi0A4626dNw94ANgJGH1WB/djRpMUk1ezdw9prEl0kHTmg
xzFupK1NgMiQ7nMXXUFCoqRGod+dNbleIq0FyMf6I6uJfQ2k6x7mpAO9Go0FCIA8
V8NqsWYiNT/MPjaVhpUQNsEOalhHdyZ0XiiksZfsa3M2wTd4ljCLQXhpMlqMkelO
b/EUkFusNqfhdD/XR0bwGCMIeCO2QwrXhCGnOWnUqTp2KM0P0WSRdrpuyslmOdMW
B7z0mHxXrHhauyksAvNnX0c2S7u8PG9Fixwim/DbHegbHNLzjV42KmhfWVBvPsX5
hv7unGrUgjKhJfvZIeYZaIk8yUyb1NJzpzhtV7Kh9SPY6FDLYGKUiKoTBGnrAW1p
tuEmKSJ01crMGlLKo2069BkCoVdno0I4lDE+tv5hl8yALToqr5Re9kp82JMb0rSY
pSGGzQOYE3IZ+3Df6ixEk1PwtLnv8GwFWr3grfbqEpFfJjHNXJm5yird7WAc+Ml/
7Kn6xLoqwhixna3F9848HGvo5pakRZx7pgXDZTLmGpWulf4gFzHiYWowwcDxuX0Q
t9tzH3RaJ/hXVZP9MOsqHv8Whfb7UpXlR4DFGjAnGriyUzuaBtOKHSyP1mlk0EqQ
tp9QSAd4QTkN1xoxFchLJyDzTpM9gY+EnIm/7zu3iFUgIIa3gICYHqduKN+U3MVy
mkI7Q0sirJzkwtgva60j09E2qFJMB+IaaLe2EBFqLI2agy0fBemVKObepDAf7mUT
RXMs+CHt3OB6kmkBVoWhX71IFDTjOrAAsWJh7mTNFuPVhq/uxYclA1cBSTLMZFlS
8bxgpLgitIL5Bf+sMBp8eJC1N7/cXu+z26R5B2TmlQnMA5VFikGLW40sJfXTCkmO
J7x5xzj7ZJfnhsxc77p9WNp10V+c3/Ab26x09/uIbjFP5Db4PBfQrNimeF4L7zO3
MgcCr9qTSyB9Wue4jFBYS7hltjMEJzpfCLa7FqkvOYNVgA7j+crmIEhiSGR6EXpb
qgj+D6MXB6tiwjd6xMYPL/vo3/FO2nH3E5/hV1zoGalrqedKwwfAcnZ+Bp5vt5Y3
QhEDkyWeKi5sBbGjzcxTuOFIHo21yP3C+cIOgGXiUNP+lj752fPlpRYMp/JXrVOL
e+AjIoADagEavNtUVi4LFSJVyxZUG7+l7bQsfTYTmZi0qiO97v0aOnZvclFWBTvG
nbiriEUgg9C5hv/HwzBXTYf6lOak2f6Qd7rGAG/DF9zsYui51gwJsl3sPy8goO4h
f+N3jgZwNywUQcjbpVSPuLUV3O0T1r65jEduQsKSmymEdnA8MvQXY7q9+CVxVN4D
yqqaqTYWPDkv5bO07SnOrsS6W2wbM0dTxvl8OZ+py9OBcTIsBf5GkLPDTJXRbufU
pTiWwwna9BYBbpkvxsfCAcUhBpOc4l1AZVeyrqilefGrj8saQgFrtNSjfRjXb1ot
aGPme1md6vdhvw2x2Z4TlVxPaxWDCS7nGXKpXXD8YaLPc7OFQ9BXiOi41uQo+LL5
t8gbDZXFymu+LHKnbJ49PcJC2m5pm/vR4T9j6nHp6De8VNsFrMgCD7NNjKnRmAWt
lVouCoUpUH1ArrF2lW6B1lC4a1vSJThs1irUH/KCYoGOobSll8VZlNgkdRXcRB0l
3C+RV+NBt1mpsr+YaN9O+C4nKLD2X5wAhANCqMzX8Ealcl6ycXhRNTOdNHr2clAF
tvURG5LNsmXhn24rkajo8rjTGIWL6OAav6bFSs22Nhay0bAdSr3tb549wUB863YJ
0euLmGdZwpFxKCwCg2AxjclYDcY64P9k52CBdpviD2uaW/xrEm8pR4qstBohGFTc
/NjJP7qluuewsnD6wl7FFYRMzEZr+M9BO87zcJauVKkqrlTqhVdSMj6Rc1JEa6+S
SbYq14ExQpZnKONXwyxcSIgWTUZe8krbMXEhSngpoXRikD44mpnj2Bk4WwBYf63o
DRBpQQkU21BXNJ+u/mMdwqeNTbab+COpwOZe/0aqWnYvxuMcGpdskySWR1lUz8G0
FWMtS+rUVy/z4C7zVE1787b6mBuwtKGVVMvZ3Kh048sSCmVutvu+Lhpmw2eLAETN
IcPxP1gZDUZf/jpHhLPll0rlMVyxfOkgwhKu+/NAXJJeMzG+eJ2098tllbpSff0i
2zcGthqtQligh1XD5ZiftfhZUwMKSPSMQEdEzAozX1v9fPokv2PhL6IDMReoSObX
zvWR3CjgZK/vshL2sF3POUdh1IkVO7ayQ6hs4BKgeojp1nUzgZ/H1KatZTRh2r1n
ARTU5nAVLw3ugzV6vZPuhfBH6hypO3ZQJeShFe2mvfAET6SIt4gX8VVlGCIhZPsv
tg4zBS7bFck+DBvGx+M92rxzwqO3SHtY3STThBs34Fmo81umq4xzkSh6b5DNiCeF
U83Iy61WI6yOKlL+wy4MnHzvPkPX5jjv71unTSgJcxN+mrq5HqckYy58ztCBHsSW
XJDwPHAjNAuj5f8FoBS10ZBqCXzWpLi8k4Tc8z7KvPSgCSAcAAOtw6zaAvwO0X++
52SEcpTXr9pP4yeDRu0EBvlCZ+CBb536bVwG5yo0sHiHPlpKLC4Vh+388/9tXFSC
szrsT0qgeDSI4DMrBQNk1LkvTaciX0XQd7wXw9lbeInG7uWZjgWEXN0gvpTFWAvS
J6bZdMhHLqDp7jqGfGbOEmOVhjWA42dKqRlH6povcqGsYKW9FgSqYGsJTzS62ev7
qoawJ232O1VpIdN6jLiC+lXPlY/OaQh+mbOHFx4jF31QhHHnO4kP4BXlxlhawdpa
fJGVVzuJ0mqeIeTyZfYEj4TPAKoyqp1lP9okbGdUP8iRR/S5gnmpeJ8TTobcZX9E
/P+ZpcCYLM7i6ZFU7inctHHPPghBk4uKNg2vphGfXerFWB1Zma0AadVVAps7KH0Y
gHBHuwVTcL+B5FhaiQqWWo0yJqfBj9SmekO8uet51aGOmEKFuJ+uTCQeyFD7Btjn
YJaeEnrbMU94WjwSYMfcjh/AFHMwLn3CZ/far8RZ6+pWQrManD5XCq3nHDUEE+Wg
EB3S2VkZJwRWPVecfZ/krXP2bzJDYAQ9CN5DgWnyPhjasuNac2T0YIYhzj229fhO
BPvT/Aqn/4QLiWwR1ARcB3kK4+8uYI4L6P8ybp+by+Qz+erSOqj8vNXPaTobN1tZ
SwY3lSFyBki2+C+Ks6sTHyRao3kdlHbZkH373L30I1uiub/3ZzDNGE+jHPejILbM
Wze8b8mp1lNk6w3vUmNHgPAQlwaYcYEg/v4odd5riYO9zQPnM36O8+7ZNNYt1WnZ
5ng1DsyET4aF8eqrH2qCi6DTL1fFViNUJXDcqgtbxlG+Fck7SHhxk+DUpWvzlzbn
FR+OGoTluzPIWhte5782WNJU3VSCvhFZ9PuzrMB+h3wIdgJdlyYXJCicKR4VE28a
ZUXXocreI7FnoK1yzPxxaHTYQ9MFH9QCnMRv9oQW6FeHwVQysxxAVLAcpXs+59Ha
LMlHYbjEKGxmU9Yaf2hRcN9CAiuVEB/R4Cfvf4Sk+zX5DI1D4BZz7+pTaNAm+k0L
AxSXDzha9qbckWN3HzXhwjHwVS/a8GHSLS8VMgCsUsf0LLF4w2zKKzs3ButnBZAi
H/HKT4vAebORodmdntWvunxR+p1AAPsz3PQRudEsuN946VVZ2wSciAXS2UxXWQY+
Vxv9D5esn3Dgyd+MYkhgN5DkL3/S9BJmj+XPI0cKjLBgYKUiQWWrKOIC4L1P/OLF
f+lMcbVtiZo4u1aLyqn+7F1wUpDC0yk/MFkZIFL9fixDvZ7s1gV+0FF0z+YLsIGL
4In7oCc4lzZAw1SjdYt/0vQTRB5Muq40ccEH3snrLus/KHvtmLmIfDrOWdyfjJBS
zEwe9jSiNZhBAO/Gy7AyrF11fWHG8rWTEfNNCTjyCKVnNfBejiZvwHMRv/urHQuH
EZdVScYbH9tQjLg4GRdzn21tlQCaFHvMaSo5k9/nGLZbQzXgjYoNmRDimeUJLML8
kuAlKIMCgMT2cGj/s5c+KmCqlqcQ+JJWwhk5lABVeFPZO6Cg1gFfDLrZyV4XiS+1
qc5vS0ae5lAR/ti5g4YwH77SETrkWlny32DiD7a2cDKDLQGijejNax1cOAfyth/L
PngDyipo8s8W8mm/Njxt+1BOds/cJpI/ChORHAGtLeNBO9H5YfrpOEIyF4NkbCwB
I6AJR+lD26LKUaP9fCDhsr3Mx1VGXEisOxpW4rHWLQF/NIp/wfj6hHfFNMjiDvHK
J/LdC/R49+njyuWRCMqlTzIfa7Q4CDl3yXVI8LXpsmtRS6NHS70bJdw9+845towE
5buVEq1iUA6m0aClqvsEyrigAVFN3FpCMKhx/NJqyAJFCMO4DIRiaiMtmYQImUXb
6E8g39r9Bj/lADGVg106oZjzruTlTS8qJXvwmCKDnQDSH1HOxuQAhg9YoPBYrgtw
vZMkc1Pf+dJ3DcydME+12iHFbp2fQNvu4CxXTKOqGBmroPPAfGPQISTZ8F/WXttq
kFL1uoEoczzZ1fdwYGNGWsbSyRb+pALVAl4B2EQvKBJXS+bdI+34kyziTbe2r2b6
xsLZzrQ+o2A7mWwznDhtHuNpYDXKaP4alUnTKEJO31WValI8sikvv82+SKNi6LSC
vv+ZuEOC5LHdWW0TRKRRtaOdgMH1j+LPbu4sDtYXqnDjLLAW48Dw0pAkcdCpl4Ty
N8SvBA43ea6lL9/nPwLXjIz2FneaFIhP7dY/JZUAHm1g0VxMzcjYdTekqF5Kjy8W
ajkhddEw1mQiJ5OjC9U5P9XtuphAQWxhuwG6yE4XrVztc4oeXkny961TwnRuMh4u
tpDa5003jJu31aZQULAeIsB3/g5R/MrLEIU76oEDRHey0Da6O0fRcF8kVJphfvZX
3mV6HqmA5ej78LOHZ5etpr65S/Wesik8PROa+QFcHPZLGLUWnpg0GmmoKjOEbZdg
3MqdHOn7y45Z+5etsBWN/Y5cH6HpK0yv5IsR0sL9epd5P1aB8dJx3w4DPuH+AsgS
aVhnSHwZP7FmhhbqTUVmiQyv5B+ua5lHWt7q2tD/XmUpI2IshPjRdnD59EWbPO5G
hDAeqj472ZTIQvMRBdyc8ClbvWK3WftzNvGMLsdnamJaGSK+odNshL+M6fbx5XeQ
PvxKZh9OoaA2niKFfcUdsMq82kGlaE3MNhxOrAXupOFZUtTh9YN5nN4FaKmm9ltZ
Sr/05+vWr+4kMEsuRNu4qLB+jWeFu0nc9ENvUpW8IM/0Cjf5MGnj7+zmiCLzKz5l
fT1nyI+YASazHvp/q4vRUhkTTCmVwqFBIYqChZ1zzdH9HFAq2x0fJ0UywjoBY/77
FULbqrLSGkj+gVmON8r71oxVrjS/V1/agW7Z4gzG0wgcVSMzRdcqhuCaPBGcW5Sj
+sCxwYZHF7xI1IpQXwU5zY8rC3cPtTnr7mu29STozktacUI8C3n0yj4r1A9/WM/w
0HGXYtaT8q7Fk8TkfW8YS+bZNAwb2OM79u7+k6VZYhFzoFI1DQQ82KPLFLJ+taek
WKRfX9x9PBDsrvlAiaD/a8rMkg3DVTXkAzvI6Js6JF/m1EhCzx8RlkI09nXczNpV
Wi4qQ6W3gZ7PdK8+IgeKs2TcfOzH9OBpHbuYZW9r/SmTYwBj5aVRUi6uxicStpsI
GIVft2QNr99DTKWWVz8IL4e4DF0VLrmvdYGMs0/a5eNXCCf6UYl/M6eslpoFVoYS
rQY1HLBGAQves8vEGHYjWI8qPxPPX6XqS3KeAHftMmuRiLxLi6ee9YDPXuT834Ss
Z4pHwMQk6efsxX1NWXhLeB7nHiBLdHF8u/8Ur8U5QluYeFbhyUcn4EhrqkkTI3nC
NYO/bGiGsPjaGFtX3PntdXQrLMl5OKJJ7OBgmkW9+ljTp3dnF3G94+XkyorWxauA
Yhuv0sc0nD29buJtbolc/9uMlrYOG8XBPA25B1wjgpl4m42jjt8WtC/e52MNyX1l
oR3y9VncvAtzjvWUKrzlv3yr49s/4VSJ+kYNGXdY33nLBiCiuAs6W/+XKnbyjmff
pNs48bFBAgt+JSsoMZRWhcS+ClQ7LcpS604iJyk6459kA+aGPUZJr4VwhLtT7BK/
7PI+pU0DIFtd9UwTd3tcuFWd01l5vYH1wE3A+1eJMhqamT3ykATyU2T7UY830Utm
GcimqIg2NWRWD46SK/b21IzYfjuJJ9jUvMRgVzmou3zaj3GmKoiIt3i/GPuH+mxE
p1ZJlvXA7qWvM3McsgUuq2uERVDDgSo7PyP34SNcYpbb8fb2lL54W36iGSvJsgW8
984xMo2Mkl0IcZMrXo9mB7xig6Z6nlzvhxHvxwjQGSVappKfneleicict/2Kh1V3
CUy85xmUvoKv+gzlWkiRwfIKIkLvjd1ABtLb99wxxds3bSgyV7OriJfyCGTQ6jyW
akoxGr2RXmu2NRmqI0cE+YYbXGdja+lffBQmLvk1BLja0ln2sAAGcyzok/5jn/4/
OEgYvb7q/QlVV9DV0lu5y4GZydwO0+iggkuSce9PzeRBzLrTua8t9uIiKGM+eeRn
SokjphGXlXYjGGN/6rJtl0q2vddUN3Vso/MAzsG17UdHngEmcrXjCqkeNK1SZKrA
kKAiXTFQvWeMjAVOubcv3Ez6lJkfvYYb+sYsBmEVCBFhBhmZcf1g5oKYi8gKGQxO
o8hR+l56P+tRo8MSN/blcdNJvSr6gdcGRoJTxe3PdDJK2zC6COdAYfmKjluXTTes
D2q3hMuXKnupQaxjHbWwE4B3ck0CaYQJRt6TvFuGMjVejOZYRng+UC44AWWcSSXA
/8bFVCHabQrP1Bk4GJY/HpUuNDGj0VzjNN+hALaK4NxBUqhgQ3kMRnrBbV9CFk/A
PWJ+DbH7e0yQVidejUXpgUaQHNvE2dkSciDmOBYc+s4qhAr1RdYTJ3v4PKzWX884
b/mmWDfXvtHxRCmukZz/UVh0tWbhIoZcp9T7/ijsMfLXwBt0SrlBbOtp/ZN5Penb
HrOWCBu8mbhB16PAyVXjjtO/K/UMWmpSnLWrXCqmfRWIm8ZFmY64jBplxvPC39ci
pc0E2TOrkO1/sh3pLy2oPxJxavZ0GZQXw57NSpnkkpnW2LnAiLNmgFRqQWHIbx0w
ZwfRZHRp/p+SvO7va5oZwsnffSkfyWXLbk+X+eVBlJPP+1kQHQvCq+sEaw/UUUrY
StYLyFuFioS8HEoCiqByJXl2up+wiilMXNT4r2xYP3GQaYUVgykFGzR5Qz8Cof2/
cDMrHr3Fm7t7OS5XXzUFP1aBF4dOLDZPD2y1B0aH6H+wNvFLd+w4a8xXSixtCJTx
JbCcJkUi4ul0kHKtmZxJbv4VlvZw4pBZlGFG1pB8mLTPk8TfUKLYJlbPRUtfCZzp
He2+qlwUTyvGvG37Dy6eZUgCJFmsW0ERUopWac6DqLq+kxrSN/9lf5kF7zsCq6H3
uTiXVD4naZi+/rMhTLlTUVK6RZLVNuiLweIgAcyssRLiE6WS4kKTX0XMEim+Cbxm
QylwkTNhbYDzb1RIl/Qr7ViIaG6i7D0i0v66S8dY+4Sk4RAGFaceKR7D5B+HNvGi
Yo9CNtyUwcs3m7amFec0Hp62F2FmWyrd16fu6Qelxx/cJ8/A59AQVI5ZkyrKmU0X
eWFfkreu8Ryi0EvEU+/u2QH9zgRXKFMlMQAoj114jMMBnHD8ZfFb8OCfHXwlN/Qk
47AHKOhzx4maa8a+8M8RnVsi+Jt/P2u0V1wtBt2B9pXM28JJtAi4H3q5Om2ctLkr
G+YZTNzWbYXlx4oEZfC+KRk5SUximPI68ox2yXamc1+4j5S+T2sYtwNZKP4RJfHa
9nhOheD4h9/xPHWKkB4E/zbBgrF7KgDgOnrOQybxAE7eRy4e/ysn0nCft3FWd4kf
4gUGpArc1+k7c3Rwg06UDvUv+LQ6TOLUsqp3PnoKZ58G6FV6OQGx7t/4AzBGMoOD
XSsERxDHknLEKjp0PqR1LxAzU5hg0FUJvuNRikvgKEVXXjctaLXIjGjM3FQxhSWG
ZH9EIOjZyxfYHDF/nUzos+2aZXRqqYMoS/A0JXarh0D2s9iLY4PTXtgCdgNuFXpU
Ck2MAHQofwcvkw8snpmQO8YbfMFMnkmEgae+cndS8cqEhcxClmNhBOByiQbceM0D
yXOd1vIoW6sy1hJLGBbSDQ7EJQAsGmvHyqjzToL6eJoelzdy8qp1EmOtgQ4+1UBX
+9IkEjCgZFh0KRId/X+BNIjdhmu6HfCsPO+3JMHwb96miSzjzTPD3HEPtf0HjdwY
SAfbeJdmOiW5cKYsEUepSb+/Irw+TqLb2AjI3LIJBS0uf9fodFeKqHDoIqgOphKA
LBal4ThFWI0ucSNxyJmfq/aBiMkDpH+GD8QNbJeNBoS7xroJEXLZnB3z6Ffe2yvF
aSWzyTbsHFAjh+ivj5M92h31K/yzYgPNaSM+wdb36C8chEwawC3GJEZGcVVeFQhf
QtQbexuTPysG8/Km++lM6HGOlKWpOQ+Kmqmdgj9Oe8QO/ocMNMGmmYM8UrObAhaA
lCQCQTxb/G3hsv+6ArpKP5wRQO/XPgOhKuTK9Wa3RZr3lhxqmOTqlH86duLpA2Px
3jpWNjH/VlQD5Wq/wC3/tqlEWN6lVBmZRcely7OS/5JCupdaHrANoaV45uEF/bJ3
5NlzsY/mPgLkyPKhD8xL0MWEJp0NDD72+X4OoGRXu7V0MmFngWjgs5sQ3ai7AMD2
Nugg0QqNsIr5+Dg3Prf24v0C3TamLzSugpQsKmTUSWIlr+6cOGOdBjiDzwJZcezA
2N6htXB6tBph2nbtD5mOfpPJt0kqXqwRq09AvdB0/Evg8z9ylDWdYPq/RnU0QJ6q
cfAh/gRbD5gJoaqVu87+AXAjNCOnIIHYtHSzImCx9pmHA1mDRzeSLw4IjvrnTAdg
pp4a3ggP94mqutqND8cz1f8sROOSAVJvFRO1wwD3FIaHU2S1jOTz/KMKtlGxsCQF
WQ2gunkAH5uyzYjM4sA5hSAqDHT/cUQtfg9qQSfLBVxxrG5IT1wpwBU/xx8K4uOR
4ejucfNpfwo6kcQawhPKUh58brZMzp2NHrfBnka30c5msYfD9xxZamFLaWeCezk9
xmH15ED8d8anJTzcaWmXxpSn5ihkXENBjsCZnnSZhalHzrLL7f5NSSmiepRXihJc
38gKo90bLjYmGJL7FDMmt1XyRffje2fQJlp1Tg8iYQvC3fsQtBuPrCydpJNT9sJr
XgMz6uqZSUzHfNuqXhC4wcaiwQwq4k/0c9h9o70qacz7Ft087ohbhh74bZ5PcfiF
IyBw6pP753Z/SCuORRob+xJJDbU6q+6KrL2PErOH/Grn8auIPg79eu3dklPRvfOZ
wxeCxUB72QzOKx9fNPkzpspGJsTFvmdLe78AtZBoPRe59VCkTtawPcMkXsXd6mTn
VsMbYQ+j+Wkqj7w/iLsYk3faSX2XlfqJ8PEs5ODWbXY2FalA7ZG98cmA6t6o6kOb
bAC8sDHGaeaZH8t8TPghgxkNXrcwRjC8PCFReMVm3xPkdFU5rOAW85Zqm2yA9oQi
rywwuxH502Q0tIEcnUd/Bb+zGnBlEqOeoU8N+WgtolgU7XYToZYni+Yp3NWOAP7l
sKaOQmzNl+XKdT+BdF6d0MYDuFAWS1y05jxcM1vLmeLi9KYT1DLYzx9h4fXCHLcZ
iFE9OmUvSUA7PWqP0uKuzjiFKDHsKDpGw+C/Wvs0tVZkz7dCVb5plV5/YIPGLEs2
gU786qhE+7YaydprswtrT3au3RGnsHyXJ3YaS8/RuA8uPQXT2I1CVd8PBbKvfKq0
O3AMdJMm6LrMXn3voBeTbt2X7jr1l6TZFxeNqezHbPpY9NEB0SeDLXkoq+pS+6C0
57PUfVnBKoPnQP3VBAt3vOr9pqZuMFqyNshpW8D7aLt7tkwEplsHk2Kyxv6BB119
3cc6zxQIIhYCqOn9CVYltlgDL4KF1WnlvlVg/vPA2YB0yXE/aXKl6/j1Ed4yxYyN
1sjRfitgvypSTt4UHzCpGTPBSnhlMBWtl0weGB5Ai+LyPzX8VaTayPKcWXQqUjyj
nhjpS5yU6+i7vBRBM9YYo/QE7s3NkqJVQMhhO79/iiD0zAKumTwyeg3uPKu+XOBE
mgAA5x1T2GqszkkP0wYXFy4nKzB6fZWwSJQgjsgQmEF+DIpNKvRKJDnVjMo0Dums
uz9dracyGiM9gF5tKflGnO9dOqx9SFkM8zdzHOcxlOMsHeIAgHo27U4ShFQAtrqe
JFEuwcDRNgIqiYj+YCvytdUhf+esAcjNJPKNjhhlYBB67DDOGdcrrFPUvlii9TpZ
nzx5TXKsKXJT5UsZKIy5NY0QkE2mx6JWfDpa1PlWxjF7oPc9aIq1CQPWNC8Tm5VQ
ffRwCb4SqYzIqRFKmaM3k4L2XcRUBFm48AGamTCkApjhEDRMC5mkcFnS//e5aOOf
6aMfTs+3wuS+q142yyx4O44WUvUnZenzpwIqAmawsILUpWYXn//NtLHWLCB+YNyd
G3wbv+8b8XnyEpcrTcKfn18j4JeKjnpuMTAi+XCZQda2TFeOWYq0D/bHE4TnjFlY
d4n3esYiJQkdpC/v9NUH/V6gZCmL/k5xAX7lWCqzlecjDijYOkJH8uM5M+Ifg7Fm
P760Lgeoo+zC8Vl2YFcvRBSeK5qbOSm3wwY7Ak9pW4FL8PemaqZd5ZBdSrILJoCK
GDaVujN+RMegyqifHi76RaoAqOqT13Zb4vkBx1Dyi/8aua1d6ni+iu5Mj5F0X6FH
J3gTfwZ4fPrQHmeFHcpwNgFLt4O5zDyTNHm2/tArHylbOy0tW9192enFeqf65AQK
bvlc1FWCznLBiY3iroL948edXGeHxULUX2Io9dd+IfL0fMY8qbZ+vrs3qfBY8QHS
+h1+hE9qMoIm/4h/l5izr62GTA0lVFnx4KNas62NfYxaeatMYq0G02Pb1pdljKa7
k5LimfU5z7c3YzR0idwUyZG00EHp8vnjRmfw0HT/EZbSuDhPv9fNwmPfWsv2GrnK
PqKpDCPAoicENEdnjqJVk6o+mN/dheVpfJfAqnGDegrAyhsG6qBJjEzNvrW0mIiL
4/m9eGMIgjVH4a1nlvOiLoLzsowxUkn+dXWrXrp95cgWkFur5uYGltJ10lO1Wzpb
jhD5GKD73ibGNwJzc310n7YimRKg9KN6BkMuPFig+/F1kVE5beF4a5Hc1j3w01Qw
zOQQmv3rhqgOgULUM8B4/amJ8ooUDbvRxoxdpJV7afwa38b/NvgEuodMRve9FsMK
A0YPpST9ZjYxCM/kEvXVYAT3/QFF+64qwfy+jzOwIw5ZuXjTZwpJvX73Zx7Q2kwj
dc10Sjzlu8GxyGi2OvaQWvTwJSqnHGxJzXL6Yz9CJsEOhh6zNSkGjOz7Ej0/Pmib
sMWCXYHEQmokffBDDWfI7SdtxGS0TDnkrHIOYBaOfuProGNVvyl25vWdZTfu2jeO
HtIOglzueOMsXw6XDaOQudxQl/Z2c0UCaHURA85UokPXxBJJB+sMuosdkJ3k+EVf
SONFkwMUOh4lsREA8TjuZ9RIWj41/GeRZMnWKHq3nKRcMsa2cF2wxlBgY/jLHsFC
U+7ZDtn1DUokd7XnFzxeDMkQtbuYrrUS3CTFyuyi84qfgYRJpokJsMbNHqy82UKa
HKVhT/6Ul3pvWtHpZXh/3wnD5N3D7Zl6PiEuTlXZwiIrQQflSP20hQ/HsnlsIS4H
2iYAn+H5rIiZjcYQUxbsmHxToRuiYP4VdM2d5Tn9+/MeVtrr2QVOHKKhhIvR4vri
AbexAmFsHv95s82tIBZejSe6y3XTF4mfSfNT6nv8gzkfI/rmrbs2XvU1JH48nqav
z4w1orAFQz2akcWvzf/njUtsc1TzP3U27KOBl9z4UtGCrhfwOtMLIkr7lhRZ5duR
ggP6d29ufDM1sIXqLSHuJF8m7QO5JdNPi/lpALOi7gm/dT3i4rBTyUiH+z8tzwoW
gZXT4sFfuA4e6tBMArxzNmdnJiiIwpHfgGf2jvjTZsffPX/VKYmitq6/k59So1f1
DkCb8UNBd0GcRKcS0xzug+rzogv1JQ8ItJcKtpXCi1eajrfZEXyVJu92QAvXZdYD
Lrt8iARZf/Hp9K/nbh1P3gxsUIUTPb+1Y4N3K77GfWRqUMUfhZN8/tKwPfDfdX1Q
tr1kQWuM98mQ2aYAcwqSp/Z86crLQq/hTZ5CorgeTv5MnkNS1XkkFWFlz620Zm/C
eoA9qT9cC2V7T1UrXbKZkVcAMGMOs/W8mdtqiVfUFOwhqgq9PEOo91CUPGkrFXf+
thPZgA40JxT/H601NK28ryAJYtBoh6T4p3h0U5L0TucYFhZF82X46sL9wbMPgtyD
EYT+xR+9FBYEvbLdQp3Jn8yo3DByaFbBfuBrwGvsYxizVp5h3HQOUJOXG4IWachh
EEk1rAeYmaLm1PXvA8MtHy9ydpOqwmdbsJ/FClop44Y4GVNke1AZlhPFxYNf6o4r
XbzsWUqZHtIAg58Og9HhJfQk4/vrxavczp+v6/Jr4YZ4XacDubV3IknA2rGWB/y0
BUPaUgnaw+uwy3Vq6CF8u6zlSNOaBy421YSeed7gXsI3sY6iezk9XKogAbDEwJfe
b1PR68XoAr24v8cnMTnYvxRMdjPZRHABO4ESpHfHkwue+ul9R3lGCtbATonGHKKq
WwWgOOrIepM7U8SbMbKTJI24oXzVV2N4yl0PwIvCIueVLcBwPT4Fom11uh+zQQj+
sCztJIJnmTNxpySqr2dvgsqsYY8IDKPKXvSgywYxxklBG59nOhqPvJV7qb7ZCpru
sMfzbLc0ckLZBUV38XBXLWVeqbW9WjDnI/MPizJF9OANEs89VBm1U307MSHSacFI
/M00+vyuqHAZMOGSOabu8k8CzjHdVSdEq2nLff2yZ8x+WXIC8yO51kwuOE6Gzvew
2OfgHBBCnQEgSiUOAECTaYDrGo0ay3ufDU8A8pzd4kutr97ioLtpkkbfOHVwloUj
HgqhnyhQfTy1OV3tTMMGO/pjdBug2jEQDvnOOlHGT3SX+5MPDePkzL09LEnitU1p
U4uO73RRwuzDagMlwLuzZgxz0vVFi4wO17xlY0d0elcLzdqQkIJ3ANZ2SuecoymC
VQFUarwPdFzReJijuXTQmhSGSV/a/utEAXjzFGp1I43jBytyKSipT+aKPYxsRQNd
iuVBY1UuAQTLiC6cPusEVIIklF2jH4k5OgMxMZpRkqUyZ13Z1/o08JpMgADol8n1
EQUYcX17N5CKluhUZBLkzS7edxJqqyClwk+SAJp29audgBLLInPpN+iVk4Rzruao
UEagNfRhCVgpev+XTBvo2jENPoOH/A0t41V1SpUR37l54blxH0quYE3Y2m6AWHg7
WThcnhd+3NJcxI9LiKmscA/BExVc+hCrC+zUm50OqhaMGc3LIC+hUpbpEZOr1G6L
UEMv1xVdQ4D3pIzUwfJhKYsYhlZZiIXFofhvyGMWOOfzpi3V1tG5pbgRCTZf6yO8
2p2dxH+pKyGZ7eDdvjxYUV1FuWAHKT/AbVyumGnU5mQpZflEVyXPN6oTqi8DtUu6
sgj5AghEeSuc58vkTVWkmVzkCG6AJ/TcKCL9Mmsu91lXwJTnUvKiQWweqa861g+N
NqmJlVstP4Xnk3zTuQBh5gMJIoae0HhVeO9ReGfAk72Bf9rMxjzpWmZhjqUxGk5q
pCn+/UGoFl18Qdl5euDFhi9iH+cGpuqOI1fLorPBQ8zjkFD+VsYbNMQmCYN5FYG5
bDTVGPT47QgGJD4dZefKLbbWBkfNOXaraAGUw0YtmwU6c47UFwmS4cTYPPWMkL6f
p8RIM4Z+7mnCzj3Rb6wzVsoR3HLbeW/Z31wW2pasXAFKoIDlHIausMHXCoB84Bmx
N+UnFAHp86Y8SL5ah5ICp7x8te/bUdwKPsBISTLof0S23XNtR98wWqgxeh3Ze5tE
AdoFk8s5p/ep1nck4SC05QOzqoDvz6fJIowZzQg70mhq7nMgXjkI2FDcIcOuivaX
Cx40eOBQTEc5HifwNtmYRw5A9Qtm8BxTGiBGj7KIf2KJf9Y9/V28tdqv+TzL8WNX
vMsT2hNC805B7v6dNEQQYfP8AeMI/UOXvu873JObmopAUU7n/xkxBQ4hhJ0ncVzU
8KUzzz50lLutJkFUq9Hxx5VFea0hvVbJbYFIx7Ve91SAVmE9X6Zc5DCQb4fA71Jn
yYYbTYcuRk3IAiHntbeuS1d35kviIqgk2JVq6FVDPCPkFTwIR/mpwmDGRNkGdm5H
CRNk1lLqdJFVVZ4xRgZ47MSss86zWBs+tKCEacgmCP6TQWD7FUzYM22Q5nLcDYft
kb25FcAbkIFhU3jxj7jElzg87qtITTLR+WQzWfNZex4dJ2meL/eBMYFYIRkP/b2v
AEKYwKxwjtFvaN5/0RGlX8OWhY5FYdgtAR8CLKvjl34MDgKw+DvV8m1BSjj8yh0G
xUdpaXUyohC1fFU/bWZXR5JqmDW/A01+NGuhRzRANKMTCBtRsggU3JZNZt5+x5TG
uqebvVdBq7gtWzo/11EYBn2LORypcfl8nJZIbjaRYr22vgRPFcLeq9Xo7iU4gcun
vhz7Ncc3rwkJyYhwvuledK+NtGKln3gi0jH/Q1GlvmS6xbnAWqZ1jRoLsTPVkGgh
kPZkIVJCsIYpXqf48hcp4Jjp85TXyYXKVl5fbfK2rDJDVql37GVPwLz42xUmUkeN
qbACVhhde8QmYtL2Bw8KTtjjnleiF//hncbdp/mawHkT25YyHuf1o8EqR5L8yyLY
eJ/L7HLL71ITfdgv0/nzdp9AkXapqFH27GAgx0Nd8tKPL0EHNprPH60CUS9u9NKX
sylqxrevQ7cY9jF/dLQuRuffXGDYyY6UJYt3ZQ5Xc0YLiWSlMUc3ZA8UsoI6mWux
qTHEMwPry5+O7foPFRbcUdptw1zDSk+S9wkE49BRUoyUnO+HQh2TGr/DlGWwYhmr
NLmaKyqoO1utV0jM3j8AHwmwPq1pcYzHa5M7N/0Dq8qaWcBhmR3YuoK6yFM4OKFP
JW/9lotsKhkxlLbD2T/H0CukhtNUG8ntgIomKdDsiyEiYdNAHrp0dhAJJLN9qGHm
3WTSgmAHMeOOsZccXdshhovFEUQ9r/WRMAu9reXL+zU79PdUG1DVhIaQ5qIgL0Yk
JPXBXjw9XNZlvAaIyeX/YniTUTl0HGV8A7Qyqx6WR181ay0dEcBkD3GnsPGs1Aa9
iJSzHpHGvywcHtfGkyhcflVcgilaj9JTv3CCyoJQ7VPaTSxRvLY1cSYbHZfVWd2g
1BQVUmQ52FGbPkvp1Xej5DAQc4WnrWhTVyYcdRCtnJJEQIIzW6ynIEIg+MsMMtQc
sqzuMIRQgz+AIFOxI/4RYAcNkVF9SZdr/Gnhr+1gDVed7uaQmPIEbriJGjB7W63A
MZn9gts4WhbIUzaTkPg+kmx8joco1UlkYr4+MMgBSrfalJZwsA7Sm7ri7Ay/bfbl
LC+OSC1JnOyIeX23TU9KaITEZBzKsRCNg1TvAPlPlOHLQj3zVLZDfyusdgKs3IZZ
VzJXuzklDR/DRGnF4WXwv31JLhmzkbjunGYlWCf8GYOONo7g7gyWTWiekiHrRJIu
WEmXSYEQ+pGBse4VE5T90H3kZp21BCVCXu3R4SWRtgjCmA9Rw9jK6OjfifUb3b+n
JZRZVvSJGMMgnREPpy05LIvhBZIREPxw/H5q8gYEpwjgzvQhRbB8zHtlkMs45u+9
VYaZy8+jsZ9B/k1MA1CuK9h7/YA45Ddy9VlPtIx1hfioY2hoGYclkApKzNaeL0eY
gY0iLbAdkBXpua2sReOuPzhdkaHZ39nawyyPWFdfWHWKbk2wbdDkAioAI7aqCUHk
QsWP/HOLk7hO0qgxlcqvHPqNKMqmYMh9z6l+9+lxyCWVfKQyimXYrwty+krmlvxd
FyyQU4Dm8o8tQZJT8XFCSH7l84crkoD1FgOrnT5jCTMEDFyHn0n61XW+LVdqWQSu
lFFDqbV3giv9WKEXJ3CLLaZkeygvyj6dp1zYTRolOAsi875Cq31J4mVnp7JTzlxR
aZsiic/ySkyAacGXtzrEoTgsaNjbX0EUtIKB6M8YX9naXPUeW6K8+JXl5MDYM3t5
KIKyw2BHe36rzmjcpcdx5IJ81y29yVgSAU8qO0MCvxHykpZdAjK8HsY+SzOR9YDB
YsctvNkjN0WoSI5KwUoIXTvf73HeeHi6tP/5KFVC6FptWoaPNBrnyIkpEoNY2nb2
XAg79Qiqi9kE43MWSwvzLeDWlFGmh0a6DXYs3bDgxcCcz174YmYK0oxiWK23SAeZ
WfUU2ZGYzNjAG2N8Fj7bXaxDfNP2Rmsia2gPq69AVSVMRnrw6b/lTvNLYlEw0GWk
kW5bRLn85eezxPVOE3gAxWi/H6bSZMBPVGgCWF+v8PXuaEwfDh/fOz/I6+npyD77
mDc8u2CoE0GScwtz6u0YxDobEX+7lhI/RT4ElSy86kM6ssnDxgYPNXqXlbVHltRZ
v5A7hHSRHHE9iEgn5msRSEJ9/kz4gzbgjw9TQarRoz7eTTNWT8HqOfS/zofK5ro5
EY6BqO/RO/cWSyk4oSLVTtb3HrfuAxcfH034PX/y5cPkiM8l9xbSfvlbcmxs+4UX
ISvM7s+M9LqCNmoQeYJJPZjhfOZCse4L+Rg6Vu+WuslqF25UXzBQVuyhtXD++pq0
cXe1JuIFPNVfHvZ4NMw2g8fQiJJuNHzyCEcv/FB6zyqiFphwjlvPKAFaw0LlSwnK
8ufffBLB2JJebM9uewLdNk7lJK1F6VErniwNUm0JcfyaGEIlVkBM4Aps3mn7A3L1
Wwu1Vo3k9STL412eHrEk6YJp/oVMXoj7ZcpocoNjtfOYYFXe5dkMK7e2FAhDqPho
U3gRMd4f4PDB6liQgBPbc0o7sHc5v25GbVrVjYArDIlDvKNqSsXOiGemamEcXeiz
vAzfajslzHjwQLemfXAHTr/VcPuobklTZ+fnRrPtXjqS3utyVqr+qDyZRBkaBHYp
pWQufjYBngMJ+nhb7TmK/NYoTRhqWvamoFzlzuZWocBPozcdevcgY4DMCWiDOE97
7Dg48EfAhDjqnmVjYck+mAmBSlb5c4xfpZKGLGBpnMtijWLRfFikHozwRdTmFPhs
wIsKcOJ7+e3VKxLr8HfsjEdDeM116FdKhK9PYwUHYAm6/jqZ06iEp39QShuV5T9L
a3yp6kqP5k2lO2lMRnsUd8/mGKEcjDd1W6kfcVkNxnELXTBVEMt3IKsfhRh6WGyU
m/4zFVaaNoea8eHqki2GTzTTUR8Um2qux2X8VXRMneYCMAO/eQ2LonM6gAheAzzE
Rj0rftX5WEYGsX+zh1KJROj0+P4h63Y3/ca3IOklmCkR896oCJRD54F3y2YWC4gz
WYzHJVoOuKRJGBeJHLpXQs4zkEQlZdEMAk4KerCVhNDxMKRPFucCFz1sUS7zM3od
9F5NIhnFTfvuv3Ly2ahutwbd8ilJ5WTZSYVD+6e7wISIbTwbqPF/w8Em1+OUTlfO
cIyPkFLQccv6hOPXZzrubVV9FD6rzDlqB2A8X6qktJ2cpmFdHp7LG++ZNs/ifvjJ
0y4BtEjX9x3pfNlB7SP4ErafC4wV8fVFHTQS6dkn5w1yAXlTDVVaFmtHuip3G6o3
7HoXe3s74PfjRBHWolF4vCUcuP5bzYPGHsKk6lGd4iU+6AA62Pry6Upj9hZRysOS
DbXRFx6WiwyKRIR4GdrpeoIjPDgLsrOGsl10sXkuFa1xO6ezEm87FEWQdvHWmpNO
4bHEs6bXYZnPAY2krmQAUhPH5fmM6jwk0LpzF1D+YRMZKo76QyjjE4nzxl702a51
iAaKe/S2ThCU5YMF/1tVvaY/JYd9w6VjoooomeKs/6Nq8XP9nKeAEX4q13fvHFe8
Xi1fLu5sGV+9LO9lbv79eLnqyyZBFKo0zgeqrMhab6aJ6b+OPaRj6Ze5vZfi383E
vV72pzWPRJYmpHRDDX/fQmpF8RbJcfH0y8udbhm0HiewTOcNIP/jvcMRLh75ACGe
5ijWG5XHTT0CKqsXjqppwyZbjwUS5NM1JAxtf89nWSir0OMuiPdA56SjWMupMsXm
frB/FhHKAKNL1NvZTAk3U3CpZRhHKVJ2p38D6RWbUnpC2oLnJ84qcOyfzQv7wpzS
71UJA7MbS6lK2LMFq3DdZG5ItW8SYYxVibmeB6yN7RK98YMmxoPTO8KwHfLxnnH/
c6SMcOzj7bF+5m6tpn233fHRx4+p6LD4cPHqVEvy4wGcki01VekVTiDqYhBzi5qC
p6fhVvbroxY2iXluROHsJ5XjKrfXpQIaWmnPCmetQzKdkRn89mDUIKk/KGnbmy/k
yYny64dGSXfB3V08rbB6+9GvWHPtGFrrdqQkU2s/WGVfQN6yp6O8buJbD0SY12rk
g2bW4oydR664jIqKNjvMJpoJOlogYICxZgBqtEX5GAZeGseMay8nluB1gU+GC7vm
afUmD1Ev+ZC3MQdVys1ljEAwJhyTbPUN11iYF2iHrovms1dHhyA8DuOd4Y1jGRmO
0PdrK921MzQTDhfkdPnj8kcbPZ3LnM0NWqxUNFHtszr3ndP5ir+TvrUT0ej0DBIU
4whChoa14GmDCTglHYyxSbGCQ4NeY3X+U8nJO5VibhCotLxc9FkLk4bqME2V/XHM
UiWtm1sF1L6cwlf3S4lSXB5rvUlQ2KrFjc4Ql08Eoh1DrCOzq1XrtDCvwj8El3Iv
AYCWKRftvXNBJePtc7z72unLZ75YFBgZl3t7qsikPf95b3Wa/BJxv0WApdzlvtGS
Mao700p2UOzcP0QJDD/EbR11nogZtavkZq0U841A2EkNyLamSaUpyV/q+QfKljDC
Fdstx9SlfYonTzJsWV9yZcdch1AkUDL//cWkpAbHcPLFpPQakwPp/zPOcCGhSisn
4kwp36ta0i2YobrfheaHolUo4Mr9QqOZxs7g2jZQgtWex0QyLvnnivDG9ADgwju+
NU+R9Ul0UXWoL5JHSDu3ztDMs60X4HwlpwvNr68GLAQ3rj7oO8/OsXD68GIMXRkU
S5uV2B0MkXbUOHursVP+SAuSll1sADwaDOBwtANKkL142HumWragO3a8v4tQPe2+
Fv4w1EW78fjakEt4Zz7Xafnnwr9ZiH8whUepA5A6k1SUxkK4LkZvgLlCk3Bn1wX0
DBHvTeSSeJEamWYFBYy0W0FLvfHPwyO/FKgnztXdQw+Np4eW7aaYjApzoMhPi2f0
g0R8PvkMJKde8tkfuXdv3t2meUaIeAKamn75sPYiRYlxVv0Vek4GhnOZo8+4BbjW
yvgryJdMjzdkQCg5l3NoWIpNg8bsxzUgY4ewF5MBpnmPx34cKVNHXiV/VjFa2QW3
DZ6Lhcw158tpBYm/xYkrDMMhR0urz1O4BpC8HxtvZwov9qBUDsXB1X6tCuxsdXod
vMh4T3Kod2Ty8o04Ed5gH9L2F2M4F9F3HIX4Pqbk672z5tru+hPjy6osRFjcoYZb
3XYjw6w9zM9h3EJQJbE30UitZzQTY3YjrX7PTikpdTZPevyGqAFcC1QFpOUWLBoP
q+23CvX4lYx+2SwZ4UoM0dhJ9DVamqq2PwtYJOhvC3BPh22+ubhPoBrxJoZREJgV
dgOyhIY7wjrTcgW9RV/JO4a29gIlAMpeL0M0l8jRZlVd/jLEkZzFr/lkRc/bYbLp
z6aqbrN8Hvhthw4gDoUngTSBv6/mypmots0CPlnxvtBIXXjiV6HDk6anFwSVOMWg
PzgHIOwIc1rBR1YO1DDjxunIeXIIanGjEGSpL3JEmg5PFmni1PhfMAV3qRV+/b3S
yU8Bsk5AYI42JOJkEo2o7ievAYH0aj0MJhxSaBexy3Piyp01Bfj4jbW43FvLnHmy
VXtWxqGSfv9NTaK4CqJCN8NcoOYWSraPHRvfiKROHg2l64BsXNn/fE7SbD7CSG4H
2YjYzOORY2qWgbbVy1yEdu+zmDRjqqk2VEZJrSwL8MQokYsspqz/fIvi5LmHJzMz
/mb6OD2pSD8So3snHvmtGPdheK6AiUu5aYlZf1N0ts9PWqrcBAriW9GH+ueRMim3
4XSZ2rBWAgVEpm0DNVNEFF9nrKOxCPwwjlKDSdkZtIF9b2s/y+UBF1sEPWeGtDNl
o3DVXjoLaZWi9sHRpQ8AmDWfEchyApN9956s4aJxsV2R+IPmeeHvHTSUSS9Nu0dV
O9jAvOtzV23xlcirltkcaEUX0fC3iiylNIfYnMnHvX4vDqipA33IuWb8pm8PL36n
xjMaFJgc5BZRpFwAMcLT8LnJd0yPf8yNxoOy1JMLJJWwO4UtgyZ3+RncOWsUobYO
jlL7CTxyoPwvNApy0/D14BTE9k0r7ibpEnySxQwp4NXigeX7TBOe309+Ua3LfQVe
dAVVLOaedb0n0opvTm72MCA/PT02OfGZsfOyCMqlJkyjs5zvekLN/uNfGGJ6PD72
mdZM6lmUQj/WqqTXyLwQptONRF2H42RkqloyMPCjzDvZXoCEFNgpQFo5eOMboMww
eRQG/zfkOhz42C6wmRxMstJht3UywCKi2VSmr6XmleAcBBO5qI9YbZlRQpW5Bxc3
Ygh/ONOhGTg27c1u29/uS0EO75/vJiUkmjNCbzo8xGKWt+zf2JFOqANOSE/Krp4U
omH3P6w60Uxf7uouclOmPHTSUW/ReccfgLmzQOXOUGEDvJH1aYM9WS9xf0xksXeC
9wmCkeI/9k4maJuC5vhPDXzKG77SeUax/qtEpJ1BQ5l954twgZFk3gyqHY3ly8U6
gsWhKS3YQkV4S8hvQ9AaUahFWVlJ8pWjbaVNVV5cjjueUOSyy/Xq4xWbwCGgVvqE
l8RbVPuexSssDh9Xdd8Qpc9t01l6jCfEILF1Cy0urA9FlBIFhDldxxNzuvabsE1F
IpW63xcC5cPzA7Q9bFkT3Ro0OgATQWT7Cyy/k/4dvgSKbz4MaNwOxP5v40kbykEt
3Liq60RSFOPQkg0VLq8x5im3yID9fHt8432fLAPDj3yMXMx0vbOyPg0MM9GSxTkO
xsAm8fjCj/pLp6KTXGgyszVWy79tiM5m33upZMl6P1eY8JRGBcHUwq20wFQqdcMt
PhdKzzfGhJymycSFpD4BSQr+A0W3nGxWpLKAMQabzHFVeuqvzmAfDlNCalWCn9sX
KrzZ9IG923CIxvRSiQ6y+baxulJYdU9S7XcrCCwPnaDP46A3mYJHs3sL8BOOHCdg
ngC0e67ywpQt5Py3ZXeWzoiRsKlrIw72LhrYVTTvN+HnoEOQNIKjwcDKPJ2fS6ge
n679/vIC9VsERlJdZCZgdIXPFSWF5djS2cFxMOS/pM3sVim6CPohYuzpHTHiNpAz
uJhnmzy602TAx71Y8Ims9ztSw73CX8VigvxJsGvH2dngk+0USb17P/HnkQQfA9c8
kIc9mMgQxf9kKXKNo7Xb4MeuQvG1gBBev0K5JOlcpPdrJPQ1LyNsTMY7swI974la
6dm7OPFN+PshGwsPzKW++E6yM4OqDTiFuIH999kYzfqSVdKoGV/lOa5KWbAPRNE/
I6N72RpUnK/DkcH7lXPk2iPn/NQDUhWFYqbj42d1BcJZq6fk7ote8RfM0o3FkjmS
SvO5/tBOTtU5Zj9XBBJ9Sq6vRT6yrsI/bLWCY22XeMINOdEtw6F10cLTd+obEhF7
zyARjWYJCmzCtD8SFkZBgStQcPZyH1KsNLqf70RD6/zlVdgTqAsYqQpnw6HfPdEr
4UHBJefBIkpmjA0CXoJunZfQt2/raflRRZOxPpmMkA2gYgKGsYNp6tADc7Ckc1Jh
l/xvGQi59aOeXH8XUjq0yLCdIXNB8KG1sZguCLj9NO28EPEsjXQHU0qHAmvJrXoU
jGhTUerZt9amXtAb/ZsurncRPXN99/iNDXABJYkmTkHoVgHWUp59XFemFPu8ICBO
PfXQRqvO2e+L4pSTCmGQyfKiVUT+i2jEw3gdkIBtSiGh4i1QjRBxecHyHTs6TjYT
Je5hApgGSnQXUzk2i+nCJH4ff2oidPmB2L81o02vX/Q5U12QcaiTZFkeaICvZG/L
VZNjW6u3ORzYMWznl4bdpVeUdK/py+jP0EjSndV6VQcYJo62e7bXEBzYv31qMhvC
lcpT1mLLdhpkaQNHerAIvJmtKhvqrAOOjNqxIbVwwBKDRTUfIbr+U9F97TXMbK9W
+GG9H+oVeuLuDbUJ+ZVl5CV+A0n01cD0e+lgHeaFy/oCV71tLgrEVTsrMeqSZlvL
HIzvo6OyCAJBOl/xxIH4wpulnOtykWYxISbnHUf/KmNr9hMqi55rU3d1Em9iVZEp
JUCLsQ+02XNBwu9t36vK41VuDUBNt2SK8Fe9AdkvgvFN0IaIOgzBoUyVhW6usQsG
9G/r1k8id8sdiuyBXdQr1BvTxuyVZu3itnovRJzQfDdky8IFcu3rq7Lmzs7w9j1t
z/VY95PVanHptFqrbrhJNbM16vmVJdJ9voBglUBgsTdKXKHtypuKYLmEaocWtWLP
aWw20NZk1KYPZrkfauJGJRGQhelA7B0GYf3qhB0pMypr/Q2wgIAbNx9HZrcDnhi7
eotVDup8Knj8udoSZH4vJcsz+n00F882UuKVk5vBf+QVEMJB2aqq76onh+d4odUi
a/XyBNSxFj4YDRKZ8Cy5+LKhJLlTQVSrWBibJNRi/X6NsYSEOCtmH5uhH6ueUkgJ
dJgSCbpyksuEKao9Jj6pq+j9JLYT9NocoYMYw3w66VEc+eeLWHrWqy6jKXa0rik/
0hJqAnS9gvTgBfoo4jXnt5eSmzXpOovU5T4NH685raj7UyqfVl8w/jE47KTijq65
MaSC79a4ve649sEGfsTzcnl7j1Terf9UtjGSdzrkbL/6nQYtPZ+q8seACurn5RDl
gi1AK/ySJkuILPK2/buMzem9S9EuE8EM0JvR2H+CqUBYEmWljLbi5g/JmBzcqe+L
dT8yCIk/8zi2k20/kZfXXd33MiKzDYQEHOErVqU/4yA2GJuGGYc4WDUyM7gNqCaA
z0Bwc4gcRMTjsE71KyE8hrWIOgkfdEZSiooyRkn5oR9F3Z6K7Z3+dLDl8ldAJswX
AipU2ok295ptgzsH+ITGy5WPUgQGVVlptUMu7JmhUYi8VQ+sx/eikt5SpyaxOgCJ
u1ioO0WiCyQyt9ycgGA1V4R7lanUZai/m/qwfPHiFAqBUiv5glgPxnjZsLN1s7bB
CLV8UnJAKaJf+36auve/fXMm5+lkjwxjCn1CDSY5RaZv8me03VDujHgs/Edl2u1R
5lKo1nC4WlSLE8Hu/7qiaeSWrqzTrJMXBJa9gnHwKBdApmsJRKxkzCydstjBbhIh
MBfsVFznhPiSKGfrE6RPRIFHM8pI4fbq5pf++AdA56xb7gXzgJg56MvwSkbCqfBv
3j+oZjbQiyT8k7xU23hw+ODueEqJnkZZweZ8yXOG9yxYHqJ9Bt1knd2rq0CDOlzk
7Qy2wHvB8KpwHWcM5XIh9iijg2G3SdnILtL5mkibk4609DyTtHmjs4t8ZsPXpPwX
lyBWgeAirRQV+3komb6EQZ4AcGiDjskvsQL7i7tyjJ2VxV0jUnM1Z/1rP/qMofNS
qzn+5Xg446+8H2v8Iqvm+I4tU7n3jsj+YafWpNfzBgnIZ3GCEFBefi1qt4sLwTOS
NfqVsRjStko3VPgMVODMeFgoQT6psa0KqoQUb2sii0MOPxisEcvH7bNIZb6EideH
jQGdvIX8OUGq4eRhdBD77PbqCLpX27t2XE0ue2aVyUL3/wS+CB5N4ceGeAKt7MsG
bpxKanh7qfF+amiLSPXm47bKwdz8sYrtevJzejEHQNCVQNucZyIe0fMdqS/N9OCQ
kIWCriY8bJpO4a3wUwNHz/l07VywciyAmLi9YZSFPj1YKZTz1yyVeafOwsuohg6H
nGuvL7UaEr1jLkyRLtPiSiQCIBf/GQ0lxbxqr4L5PGiqbbXUZld0h5LWyVj8IKv3
kWuI9NpXFGtDvHVQKB4DcUxfREJsldFtLtKX9Qfqna0UxLdXxiFKUWrYHSfCKD11
MHr7wBeAS79FMpvjG29ewbGyPMW/2YSs3Z/BJX6zjQi+MgAzAPO4vJyiHvtTbX+/
Oj+teuHJLOgDsWV3HDXf33jJl6BNMp5y04NC2wRoIERAu6LXs3uiAiMc0Ou4RCE8
v7+0NO1HkTQCrBPWIzDGDZ58HHA57lhXY+yC22Hz3asLEH5EywUChLalevRjkHbP
cdOfMu5cHf5PERQOOFNzfTlLMDL1yj1gUxsoGbZHoWOQN10XmEVdaPbNd11L7Xgl
CbaeH9FuQo1fowWRvh6pRb7qXEBWe4Tgeol9ebrgAzW/OatQzHji6kbyu22/acGX
BYzFtMzCBRg8VZpt3/PRgC/TdcWHOWJ+fKAEGE7xV8G9r3dXoPAx0UhthMg4y7de
zO1vxxnmHqOjB/Okc3ufNcEgcAbYv4Pl4hp7+ibqBgus+A3AuUoyyGZ/Amo8zPAN
jKItmTGaCl4UsoSvaj5cijpgqfd8XI8NKrhUhZ9WXS8dG1NJhdz996EamaQjN1Px
mRMnADk+oe7Q5gaBi8lis70KgXcN9Vjcl/wHZn1+VFudkDBgqZtvjMdIpob3+inj
qS/QiCjjEUmS/cdXvAsINE0GPlQ2CiA22UoUDkzZaMbpLIJuj0BPGPBo26uzqTJu
nRkDdh7TE3pnFg5nzi2S4rGBBX53G96vv6qpPXicFkJRMR0zBBDpHhq8SOHwOcUv
q9thw3g4Kjn5+G7EbYtnvs3mpSSezCSLDOqj0smKagyRk3QlMaPeV3Qw0s3baDfB
KwBmDV6LZqt1kdNiq//s1W4z4oNGXS4wbTcDbypVtvAlyY7va6yfU2I383JSAWbw
WkRvg0xDqIyHdXsJKiFEuk7FoN4p0iL3D563bjIBiMazE1aoRvLgMT87LEmStN0c
ud36lI2YMkCXRnSz441KC8Mxo85Mdj6MKo862q6Ad5b1tSR//lHqKEzoA3G6W8bE
KMmlYLBPq/wek3TdzJkf6HiuxPmNdFf2jJENJyk+pHdtEGEeuVxgZ3+D318BaTrZ
jFYGdHzfyUBYGb9rCJ+MjjQXbOan4/xvGxU1QCL7tKGNFhCElK03pd6Otz63Hmrl
T/9he8n0ntsse8y7PI1qmJ4v/5mMDZHBuqoqRkyc7O56puJepTdop27fmUadH2ps
iNmnkZRYVQikze3zwzgcm/M2qxmmoMiwMJMqYa4ti+WlKfAunvJ0DkhHC8T5oOJ4
aRcIgYbA7mUFKhZzSrFXWHBuprDlr3GYai7ntuaffGF7cJrfd1l/wW3sVy85mCDG
SqOMZJFZa/dB8QyuqZovx/CliOtwZS6em0vXgp65UbAuqodhiPrlHaD1KxGqNFS0
16y5JNLz9ujS8+9nbZPETlimuEBRDAw4eJzgTSHxRokMLTRulPU0Ji0Nqspeyx5/
Kh8efNIU4u1LDP/TYE7fxFBldObw1QYTXXHn/fItvdEjcZwq40qnejF0r24STb9k
LEdkzKgOAYBfMLtQYjJi1OfWyxEGh8KCygZjefjRU22IdS3vA2UrFYKjDMnVkARn
2HJFD8aAGzf7zUupbERKUofqghcr8htCuJEHCLAcwmjqIJ7/0HJ4rFP8XJxb+f22
zViqaAovq1NoCTEmSJHTWsZ4XmHwBbZSurM6d4mGrIP5Dju7IvoqC/v//eRSQpaF
wQbKkATdAuBUjS0RNRVIPcUlgdRKANJ2fjPuZGPsMoSA88vuM6I3mEpuZbZNEK9s
XPpBXiN4sORuAHrGxfY6zhwIAPBRY2/akOs+aW7vPjg+NPueOfefh1tYfyZQXyU8
hlF8yG+M5mLZK4nkoli9J/n6I8jjtiQy2GsU1YNARHTnhtG1FnHZqiXxwRtDfbxo
4yAkHBdRw2O7OOQNg5tX0quRNrvoUxZM7QEI7umu6gTlawEn54r98U7c1Xf+cMmL
CyvmaVdRGSTbwyhVMyz9hm7Sf0ZJTSrHY3AXnqI0sqH0ipTxOW56fUXKPUABZlPa
vnoe6hHMjuifmC8m93zfq75Mp+OULblJuCVSwvufLvLKMteSfY/N3uXyQch737nP
hEDFZZDX6wqV48aqMK6TUYwiuasbHXsgPQX4IG3yOMvqUTqs6AUEsMYpwgBmK2Jx
JNdkcgIQahkcXbEKJkYMjMCsBZ5QkFfLHUT8rrgixlTLsba+8qS60kgrtCSd44yi
zTSdTfphJfWMMvlJaWRK/myj2dAHcDQjIsN2gc9z46XS9EcxLu+3G5twXNHSMBbg
kQCpjYnA2dmuXnOCu2kWMxVTuOczk/qWaGZfjkl3GSAW83xP2l+vUFmYkbwN+mOa
DeusRaZ2SAmn5gW1+LrP4aK7RvHS1glVK+rdCp043qDSzIi7lVY1ew5U/dMDMtzK
VvQ2+3EKD0dJG7U/DR/lGYKU//qdsqVehkXDTbQSWygB14Ih5cf2zLe2BWszz2sE
IupJoCZhNNOSRD/qlubaVTTipttUDiA0/1+n5I7bsMxXnRPm+xi9SZlkBY3duXEC
xOSuiSYHTpNHpfLfslCMVummo1ImkPpBmVz0k3GP44xyJawtjqQJ0fiz4xzlFFwF
jRJbBwYitcYNI5ZRzYnV/CF4eOeHOpxv5jmSy4sXHaT/t2JX7jSSZranMOgaICsw
t6YsbnbS8jYSiezRrkdFvH9VwhAugSeFZcT7eWISALchnfBAppgqMLVxeuXINORL
XmhFuYejNnfAFv1uu8VPGVfOU7tLucCxsYIhWF1mZ7SVU0fagoC7Mt/BcnRwNzm/
nhvOomTH5oWCu1Sbe9IDcUnrDwrR7HTMPkjgg9g85sTEr5HsYYAiVUdENorMB0mV
e6ldJP/YuKN9p/4sdb1tkfyJ47QLvaXirxRBMBRpBHleUVT1b5owDUc+HzPltkwR
zk+D2C2jnfGYe/m15+Z/ghaa0qsycj6peKBkUTejPncPNPT3U3V1i81s70SdsUXl
Ep6h4hyrJaixhf5zg7oivA+eEGe6bwn6+U3w0423bHSHbDj2UK/2HQD2X7dNE/Fa
1nZx9+MpNSRU5OuPqhmRukwKZhnnoMP53qzsjBnrNnp7vXd1JpxBuFqE3l3ZXyYm
FC3F7jZ9Np23KsRMtahmDuO5TKRXWfOgQJvkhKYY9poW969jPWsUwbpADEtpiRWc
w121q0+NfQsgrKNOFOPSNBLqYU9bEFUkLi3C7Cu83RlMPoo8VdDvWrqxIHD8gEZM
Ce5wy9tG2ly1YvECltWRgyKBYAFznKkoJsGeGfR44IWpdqIVX8U9Z8IOIjyA0OAy
7rqa2AKRJ2HkjpawtLTNYxXveG4pzkp8qPd8yQp7BGkgNEWxtcL8+AUeYZZ9AuWw
XZ+ngDUFBotdFy7h2tNSa+nq/uYyrzPTsHaSfmjladUpDjsHr6btCZw/o2ZkgT0Q
9Fjjy70jioATla63PD7tcl7t1Y86pJlBiJWS5kkKEha0DEMV6AZrLCsbWpGv+mu6
3KPZUI1OY678gFe0MI6EmulqKljQXx+o9Ia2X1CdbzhpIibhP3oSypoASa1PleVS
Ke4wfFhwHhD3KleNHg5H9dgTJ7vj2kzDAkqAeWAetkTROOejHh4erGVYUkrxQ3pl
7YSZO83ywq+12mpWc7eCcjFwTYVSxPOiAYaJ4/g56KqPP7wnP96GfSIg9QhqglsE
3IfuauWGx4aoVc0w0ExTPF//JiHsljaNNNLz+0aywpxQBDWw684H0l71khea7xJb
BMVcVXYvTFTUAaHQNwdIdQYtKG0we0o8pOrckJr3XaQQ4njGi2khI7hvcJ8z/7ij
3V6PHx54R/v7oV2VlK1W1SvTH0Ca1DxqLKMVjcR4+5uLTBoMDc81k9lXMn4QxWfZ
wiIHrXvLvhbdlcEJtPDXIfJ/x+zj+sQMYBRYKNP6QHG7VOjs30Y2Op9uZiutRPp5
3Ild10fY2Oip0HZK/ZL9kluzFPo9yizaLwkXFfOBjRKF8el8cSpm/m3VoKMGJZFn
/xulxigE0iGMeSzNO4LEi8pFyo0V7whW1tQ9XgrMgsN4yjGXnD1oJTqCbehuNdzr
KZF6X0UjdiNOHqOhAdp0ZbTm82bmrfoz7r6ez8l7falZL60ZZc1iGokYCEKhz74y
b+xWAvNijAi66fdK8f9ZkJIXo2oyTCkGAdKXjL+Sa3ERO5KRutQf1pjx6FLFnqqa
uz4eCT4PI+IcV2hBd4bBVt2U8ZnN/m32bP4A7JR91Qwi+LTYrFjLnqYZCm8IHFry
9kOUJJtJn5yCiZHM9w3W8W8V8znFjg7n920knUKFEcv5Tmiq8WMyWUMka8ZTqvi0
7TISeSLr0ELTprUmMJKIDJxoIy9XHYvOeOXtaxezpx8itTFrW9H3+wtGoDS3s55x
ptHJk/lVWxujzYQ/ACr7UafM53MDUBxcGnJL7mpqOMw3Q1XtosAj1UgL98dJBHJm
qsjVLmXobjeXfph19UyfkqQnDf+xbdYNhKJl69XodlBFUhN/aTF+TXbkFkzvCJx/
TIq0r0gic6pSCUSGsjdNDHm7ovzOjx0XaZrXlrLNsVOubR8C+wbEhH1pCTeOO3vp
fuhtf9RIbKS9eE6e658P8Iv9GP81WXAtQGHKnn3bZ5XMNn320N1Njf2InLRweWQj
jxZoDayAy5Oib5Ulr7kDxCNQDr8zBmhXC2dzeFIm7njnWLSc7Rr3LC0TmCH+Snhh
XV/OHkC1Ce0vWILvB/rtuRUwsji+t06bE0aMfHNXs1sY5Zp5l1IXB497O2FHECc5
/IaN9nUaz6SQwFfTRoQ1oZDuibsrFgE0W9Sc+0LGNd5OVnMxEqaOmRgq9RtQAnpl
OQiUsU0oVn+NmtFQStxa82lFCbj0zzfe9uyVVBFw9s3Ak3vNltAMvxHLSJuNzmpi
c44bUurCOntpAGO82kxdHyJ8XPysNAc5UWqDK/7578RBYPkqKoFx8theSq/rmXkP
VAUflTbkNIiAZWd1TrzfXiTO6uoa7Iy5UgNUSsxYcA7n365msEy2jIJfj7Y4joks
yZr+sYww2O8zTvWNEYCTFhHaZjhV8Dy4VYV7XvwWVzqkZJHAc95xTXlNUSxWUElb
rUF+6ac+wZweNkdoGcHrLInc0Vdw4NWhchX1qqViklRv+ZvLi9jf/qL+fc9Pwnsd
1AejqLososcBz/8fd4ffpWpMlwaayIt7ja6N0v5KH89GvdRfk5P8z0+JShBV3/9o
do8x/gp3K9nDpn1KFA7Ukuh5GeHOty4umjHAKBxZjjClcQlgcC85RquRR4mkPB3B
N15NfwQ2AoAo7kcsas65RAYPS9hTbYHM89Ah2Tz+YXRFlHyRQTMz4ESnan4RYslT
K5tpwdyLT76IzIxb+7g9kdVSkzYMVSqQMPL9PRRnhdlZbDpglZemua7JZQ6jh3MR
KNEPDhzOzJK7EV6c0oZOcH41H8oDiZjWY1sn6tyr5XFhcfkEGAuCLqd5+AERoS3D
lswjz6RDAPSoVtH7Ot2GpZLhC2F0OMexxZSMIUdTRxIadzqHtTuGWwwhK1usEoMI
PrqNsC32H4LlScTSlMs4sZtLnE2CErpA6Pzwa5bqVGuOBLwVW7RJ9Hp2p+uy8X85
h2qFHqY9PNrz/IRfFT3ClDlU0L/CUsjKAIyotj1AJJ6s8cYNZaAdycFyqCF5cmIT
JF5awFSMGW37B07vge32G/bX8shh29GFLQTqzf1dQCJIGI5NxlLM5wms9+webgsd
KYjQP7hiPL0HjSguVj5yiBByd0dDxhHYaIwrqESWACPPL0IK7gRPjeWoXuZUhELQ
rbVRlq12pxbo/WLKCMF0+Ao+SdWg6WzFOgiAd2U+9XMmUNPoQTA2YKWAzQQOz3b+
4dVZO6xLJ6LLhp+iTybPqnCdX6vQKDP8O292FWzpPfwmu2BlcG8E39FMtAvLLr3T
roYFKwm5v3UltpcwOtHSEgm9XBBIPkCt1Xt7bmzaMRtVLRKLbhU/GLXRV7tr2cZS
HAU2o8p30EkRQUe4+5vw1I22Oa2cA/wcpgsiKta0os4siwAy+02JPCjncAV71f42
pclROU2Ja58ZBUrJ+IvovTv/7ZKbk0W/p0BzPEsyzcdOFRvtnYSptPgddjjEntKS
I08MhtEbCHpd+3D/4CDtqXCOdN6pPxRlCoDxdrKA3lqxBd9gammueDUlZCjfLlnf
EqMr1+4J93F4PKkzKAYqMlLIQUF14dxTZw1jV/F/W9hyJYLrM3uoM8rzKcy/Fl1D
Mm4qaV/U1EBT2W8rLgzweDlnHDfMDP4ZvDs2ZoN7ZfoRgecrb0Mf3GwI4K2EsP/l
Z3oAWRrvAdEGauoir/wKi4IwJTsKd5t5xFyPRqOHAz9TIdjsXi9oqn3HRfZaj9VZ
vwpdlCuSmD1aCwTpJuGL7e7nwZO2cJfhyLKATsokyexLBXlsjtM4tq5Gs9VE5UMN
5YPFTmX7ZGEhYIc/HSc8VcdmngzQsHMmHR+4ZMXuj6JVw3RrSVhyUt/gN9WS9VTN
NJ2Q+CUlLDTBRELnz5NeWi8i3HP0D74RI526h6byX4IVOGu4sNkCmLIc7jgTb2QU
NpKVPmkRRAiaRtc55beY5DaXBjDlV6bUWnOZFLwo6W6RZ/ytSpiNdqJGr0xHRoJb
MZmpM+0ZTSkZPNzSmWSq4HTWVXtl57EpQlIy3zCpzuXMJ0cERy9oep5+1gcDM+tI
BW60FzG501lsa/oTOF9SiZWvZ9I0MHiZrCwLmGvvTYfq3AJhckKLCVPQFfFUteRt
0HtbeUi69gzLLGEX5SmdoPgHA8aE7Z9ildXYPxvtNVXYHFzgswpi3dzmK+8fXxVe
k9NOBlJpFG81fHr05Xf07EKYyvVbtWDFCweQiWehcuNuGz7UAr4t45vZjyHOh3th
y3YNHc//cIDlytEAjwpJH5SkbomBmcbQ+id22JsOMBQdPijbdfTnwGSxPKmQbCHv
BNlmRlpl0CpYgB8oXD3m+kfukH0XOOW62jOz0Mbjk2gZUNAQPbTf+BWwwC9Os+2w
Zgyyo3nP/v+p9fwqi8kDXlSX2zz+sOhMpiSz1eLv5wRdvlKPo+sgAnskQUnM14/i
V+XWqwDrpRz41PLsxmtQYgFIiVB23uckvIL/AUEUgl4MAHlqPziwZ38yvbpDf06+
U/TiTGo9dt8v459Bt+AbR2FSB3j6y2w/bZMo6fOVuibVYr3PqzbfLxkHe2Ognwx7
Mo/pp+pnX0A6MizCp8xQNcStJdJkyF5z3y//B/AH1Yer9RL5pTIXBeKf5qVDAAvH
nVAsU2APVC8dGj08GglO0A81mqx7N5T7S2wzuPrUdSYsOvBUEU+zuD7NT0XxGMay
nuEfGGl0nzmbJrHVG91Yiv59zZIrdQdxHjgeZDOGV+558iNCZDm0O8fQxk+3i4WC
dIYOl/eWYk5tIFoRIv+OqCNCh8NwVKlvEtpRR9gSwyhGHBKDRzWTz/PzedlLVnyC
/bGHPDJe7jTxrbOzoJR0Surh5QZfAGaZCC9aOdK9Kk72AKEOXaDOw7HDKUoSZnUt
MOaimK6IDsxxuYNZa933jZGiasxMV/5woLd88nb23yYF479dbmRLN5iSUfb7yYbL
6O4Jj/NbeVtvbSxLE3eyUyi9ijvzM6LOsfxa/izChD+1FfTrY7Y3/ZHQTtQLDUOl
HoppctZ1AuXhBAYAqigjpY4ruR/yYc6jiZT8wMVYx+rj7ILRV7x/SmMO0pXigSiE
jOrDXg0p3sBO3EA/+krWPvt4WutADoCp1/60O9hlLHwa5Wx6nfFrAOiAAPjINIT1
0eDaoPnErJ/CfVKe4E3cmyEoPfn7fUpfydv4S/S/VmC4T4eDSTSYqhvWKbaVovve
59px7LgBJRTY6IrtGUe/gZ+AiN7TZ9R3uoXmSw+V/c5xCcP1ubxeOBO3ZpIeLATP
Dupaosk4PmpF8BOYP1DcJJ9tJlna/Nep1CmlzAiLSkglyxAUJdvt+jjeyC1t7abB
OiIWuyySJ/2jHjgJnx53XZYcYfb2KifDrMMh36woq+YZTo21ElIjhMjZdWqhTkxN
ljWV03ylp02MDd1OoHjdVJVPkKrW2k8vHWgRJ1mz7IdxFaYAKPZjhVOgsVHgFQOH
ERPqd8Bjr1WCen1MMKn5Fx43A+OpB7NmnTqizQDHDK5bV8pdYVEB4NwqEgc40NjC
l0wdg+NOxIkajoQoB8uEv3KXmW2+nhVjd745d6X8AAj2jP9g1KtuqZDQMFUS0vOg
pp+OpPKrdjA9Jvka4siviA7o+TWuy6zN/8sfgY9UP83OJY2oe2yTWFlRqjtvuChJ
2nDILTQQ1LazL/+rcK6P2XIkaKgryG4K4/xHet4IHUmFBnLOOx48MBSgwE+Yzn3V
2O/C1t0VUtWCsBUMwoTmRTHI4nWuuNadDs23RtvPIVMlGRrcPtAFYgNxxWA9uQcd
3+5MfwNvf9m1BOeSQ9RgxzQsXAMmExPI1k2CNSxZ9ZIp/63Ae8oyHO5qWXQ+LoZ0
fOvae8S8o1dATEc0XwpWFR99b4s1ZFMygAZt5kteoqgcjCgn3n2aKnFSXnEjFoEJ
+28t//pJCSBPaQvVY4372sxHMDHro11Ph5fJYwB8JvhIUrG8zAnSZ4ce8ZFSZVXr
sDR85jAjkVBx9lX6aG/N+5HxrwR0JBo8h+DsXYFOZhg2xRua8syYLmOczJ4cH7Xs
4NJXvYwunGbk6igXeOkhCbJ9krilRpCctOd0/CU5kdfS21NU2Q/nGqsmIUEBMEe/
Y3XCBrnI+ZbIg4qXp0VKhctlMWGtcFEkGmgFk1fTSQ8SPcfkzUCB9CTUr1AcocOX
S9uA3sYHo0SWIIhPzuXtzcwt87Tur7AGT7tfu40Rsf9piuoxWiTRh/ggS07Y47hY
FRzI+T6HDa4x6eNcmSe7wCfbE06UmszMMTX8FtBNadA7Hfhwp4JtS4lOAE+VDfX1
y+OdRG8JPms4nIj1mqBF4emXtM1Uu4K0fJ/qhTh5QkDEeFGlb6EU1fv1NMX/A1Pd
9bd9jiynfe03lcfYcEsmm5zu65uToGp3wcpwod8mBJDQDok/yH3j3nQ71VBDJ9d/
dEcwQS2A5dB5+N8c9xj/Kus6gBZOFbisI8RNi40tCElFchMfYfyo1WZU2xve6AWn
PuDKE47l7DeF3HtEiNIeH2V1aQwYwPDROSrgbv6zi4qfl4rbLklbR7rq+gWlTkr7
QOX60feZyhTQREreWgRGYtXIVGWNRhVYdYT80lu+fgVbFsaOIVl9dH3j9ddj+Mn3
lnyjcAu3Blz+mRahRrbGq4Noy0E94hVnvA+YjP2kgxAweVw5pZDdtVzfFDC4SdwC
3LkFagTQqE4dgjrxwIXlR3j/TDG8rnndPiLFnxjlYIWrjB+EUAyIZJpoC5hOt+DL
2YaPrVQveVv+Q6XTLIt+4p3o2c5TE2AGLk5OYvLcxy0QJ33brPNCEK54nczHV9Ni
ioeGPvDKDJGXxvWyEOAKW6HbI8T6fchM/D4vnqRRVtM2/lWBOpBdiOy4sjFOsCM2
MViXMZHs72cfj1gopRwWxO8zZIFGaKrwavFTE5pilF28xk0SV3hrzWYOUoqz1eG5
mOqTJ4wtZyaJmAv2NuWBx/yAor7+MRIfy5PuWJ/gTIdU8mNKWXT33inZWlOCVPDv
LuPSZhEZY6h+exuju/v+GLWUQyqn5stQCboqRezuwq546qb6UJJAgg++WoU/S9xa
wyd80AgCat+uoVpkhmeUs0Z/DVp43+UW9YkIi7n7Lv5kVDkoFDrbZrF7FhVvYxDr
9gWS2BBYg0Hk7Ca/wmbF0EgCB3shsBDw9b4a6h3p3K3MQf47o1wLAY7r2jQOwqRq
DewbK/rLmUeNMSluPnPF7GxCoyYfKRUi8NyeFfBHc8O0ma83nDg2c0e0//UCOUNR
S/Z9aClzYeT34vkDgoErwr0C5PnTRAoyM5NWNSas6k4kqC+DKeLq0U/BXPCz+O0v
5/LhHj/KdDcdy7p67DriyZPS+W/aQQ6zCpP9IQNmTMefeKQf6YCUM1tsN25Gms/S
g/kXUhL4vzsbX1EnWOh7kixeKYEzChEZMtdsNczJHMXk07YN3CwR0kpT9mDyTI52
kMJB6F4/6me7YDYnt4VVv2dhwzI2vaT50mX8mhFqCQMcA8utsuxNdoZFqF0KY3rG
82KVN9whSk7JNuKyfpfFBCT1af3GSi67JCHDag8EVqcW11phK1yJWKbSu9ypsnuG
iMinp91yBx2M9QF25bCo9eBbV50URauL+vvPEd2S8TfMvumU9MPeY46BORskXEe+
/suZCR4x49MtCsrprn4mF9KUHfqFPj+cpW1KLbin1d0/sVwmXx5e0mrS5ZbD4Icf
j6KjrrK+LEDv5pn/na9NWrbdroseZeC7j1la8appZK6byikgan1eMOTBKkASyXxZ
8nLmx2yEGkadNIcUTLv+3AY/goetDMWt0vm9zzMPq3Epa7B8AFT7gaZBvd4922da
wVas6Js+yNPJYalhoCwwutbHCTRQR4pKVD7VvKB99eLi/PqfVvtU+foyeEIv8488
ELp0NzBDYze3EHQtT6QwKgC3eVF7/Hie/vHViadB4uPUcHyfBCcfNw+q7WPKszO+
Po5C2lCwjpEzJRCQi45FCIFiwkcXzgkIucQ0iWyEhfs+H7Z829S9JyrDqK5lou/R
+jvDIhrXT1ADUW393rvRy0m49SrAkl24vD1p3FmqOQ90TGv9XLtl0o605l6Hn5ZQ
hssuzbMIYJZpuvuz2BEqHbpfwfK8RI88/53rlqXSDY5TKR9t+vabzUuLBozyZDfM
rAdiM96QncqmnysAh5x07tSbwHiRaZM6uw31Qo3LSyBN3rPyot307Id7XWbQMtdD
VZSR7qpJqbicQ+YA4T0lIEhmeY5R4XeTUQv7Er+0KgXWfOkIFL66Q5G/CUeEz+1i
OA1HJnx878O+wfvIMb5okw1N9a5rJaFTVPReLe5LiRqVyn7erzVQZAK0GlI9Q+4M
gEx8b06AB/0RYuh/7/vqLW+Ri/cofrMWjzbiWzM8w0hIGoVkL858ZdnsGJwyk/98
AbRmQ/+LSpKHwPJmjEhjpjeZ9yFoiJ0j3IGye4cFhcCU9B2tkuVRLr6Y1/RncEAM
oEpFxHj4HYBCoYyGPhYGXwm/3knPmHDSs8+SK+U6nnYBnLx84+691z1lTtdxBSR/
nqBeN4vDgtqaW+2mpvvYn9yj3Zv0X5JfFOPPgtAX2SfRlNTRJTDpO9KAu5LRyhoQ
eYtQbeId+j9Aoqr+ZlFYJqXRr5HT5W/ryF6EO80s4x6KsRhbFkH8VKoEfiTitrKP
sWxVYxA2ucOjLwwKfz5o5P+tU2NXNFbF+jV3JnntPIvQDvqvJUYZIBVjEJMIa7Ms
HYHyw005/sHKee//tAEMBWwrfYDgoVkgT/3xCdAfGc8vtDu12F3vRCF0Y9s1+CbM
q7mey7VdTyi/jAp62nPc1G+85FO9iMtxNDQ3frps92JIq9iQPNgSw2FQRsy2r6G6
q9Tt/EGO156dyJdlfa0LYRw5ruf3j+P0nD3xbaVayRFqgzxHmaHInx9txWE2RIZe
a4enNxsvVYoVsuJnQiCrcV0EjsGxVSB63Ra87OjlzTg9xwYkblyAxtkcnNkKft1t
IifIBl5rVD1S7WlSQ7WJfgg4k8mjsiVhOPtEayokwvxFUFlo9bmiG0+rSEQ/vuQQ
Xfb4efPS7JMk6TlVBlcDd/bKEsc26enK1F/21gITPuzsMeENPIHKPmnyhoEAnUUt
YEEqTBY4OqNakPpzO/tqqy0TI49vXo0rqgieKafzVGHs69SlVPuDs00MioaCkVWN
z3womxzviIMctHMs7DSAsCrB163w/+tKNcwxx4VhD84ylL/afBb+PtVSIbq8oZ2M
Dwm/8rTyGYTKZ1SleGjtZZGaXpZf1qOGRVKjr4nvw5d18PmwRMeRcjSPQL7zye1l
UnuZkaq/rAPQw8NgTQWEaZGiNYTnLb7b/2O4VsdLxcKQ7lV4uHq9NwqI2YGjXCrk
YCuX2AvhGhUpIV1xD6YPIs4muQ485vcUxfUxFGJ5NUvQ4IH6EmMUzeR188MDofyP
XORQWqfQjdPQTfDV31gv6He28NMss2HWwoQtcn6/thgksY9pUo1zrVcErkDuTwOp
V1eDVDozAY/IX1yRPHAzGH3cifDz/+z65AcU+SLeprBVX3yjD7mmiF0gO3lrobpz
Az/xMNqENGJ7bhyMIcjka8+F2uI4yo6HZfr84patktIj3fBigTujVM0yWx3Fj8rp
njZR3nEzjO+NZQe6SD7ZRtI/F5Ap/mZxfltZ0sqbqQcyX4TUgCBpL5w53guu6QbP
uiSO5KNLjGskGP7nslUREhLqmxe6tmCGfEu5vPtPPnqKcATK0TDOC/JUn75iG0BA
KMZkWQ7GwSJ/6mf3/XHaXu1nSVVbS5Qx63s0a9ZbIDBfydagHjoA4uOBdboz/yj1
67BbxeZkjJYNRVFAnQjqxvCo7DPufltghoMMzd/HfpeyhtEuW+TuSg93Bva/xT+w
QSrx7KvH6qTseEtV6Zw9nF16bA5li9ClWnRPEkeuXhplvNh2zd93zsAX7XRP2r3K
6uOvQSgZS21dKBa0gByq7bBAVPcuiwQOA6AvjjIRGMSn7u70MDM0H4Wtr9QDwgBK
zK1mF/IjxWrcY8tam6+J5B4YcYu+AvJ7rkeyKCkLX7h8vpGn6QP07kWZ2YtZ0ddv
nPP/EUNGaKQxYCmu1CeHXpSOdvKmnZDMlY4yhBUJTL5SwDWVdOuyqja3sqtAveNm
6bkTl/eOXoqgoTwmTgbRCB6zxPwbf2cK+mT9Ev6ETTRvw8Q0iud5jCJ+XYYZgZL0
rt5x/TK2sJBy9oICW89Jb9MAoqNObU1od/3hIAqKxqSjH3WPWrtAqDeuqniO9xwY
9YBs1OZVtP2g9NELtMCx3bLpD9VK1ZK4lpGqXrSfRRKNc1OIy9RDWbZiEhwIC6si
6/FiOwl7opkoajfU9PEeyxiMrsgZeuqR9uus/ZDokdTyXucmCFGsghaZCU8tS5cX
k9+YXKOhgW8ys2B+k1S83UZNymHOLjfqfXYuEpJQYBFRreTl3KEpRxQHs6QCigQ1
XiYNjSYdHgLcPSfTt5dtTzI7bX9pANmiubYjw3IkS3myEJRcSX1WAEm/OXSH4vkt
Hwa0p0wyVKhcQCSBAAn68a+d47pM5+OZazM5pyMq6Qx0Nu9Gd3a6fX1MzbK7JRfC
s/8iSCzxDuzrvWxRdI4DWBCigJi2QZIde3HserbLUzDybnYkFFvCcJmxRY4KWgqB
41peF9zBZV8842Eg5zAcp4Ir8STVSbSKSllLPJH+7o5g26KAUN1z+F3uCBLWa2iG
yoimuWPOmeOzxd1ffS5SZMyToosYqjTidRjMAIl2vRNC6JXszoMNbq0N0bqBwMZR
fHSQ5VHDdzN4cTaxEQO+QNJOKUuooyO/V4d7YU9FOqyOMvL79qnKyMi7U7HCaD6S
QjHZr3f0CBBUSB8yN5TJ2umQQbSJHTQImO5W3OuBB22DaqX9Kmux6PJitTOrNouS
j6Lo0GNNgR6VJJfSVcifxa9/JGNvagY+wdgYj/H+nGyBNZj6D7s/flXYe6Wy0U5z
pHO4hZ5MLB8SU4CKixaB8vL5ub6+l74f5wQfmyRmpjj6Rb6XuQG8/yTnmFhURyXD
65Bp8b4OJYohGrqH4TisZj0Bkb9KwgutOk9AqamDEzNXjzE86zwsPDjETS+yzYmE
/jEyVj+6cy76bAIQ2ArUBCN/AC1cjU4TMVWgoiOqqkLKxCo61AXbUQHg0fMdup5K
hvgVJDUEy2kBZdmbu9SAja5bHgjAy12DQqykqrx8ovAR4b31mStkmffaH2cbk+I5
kkyi3o2BVZ2qzo4H6H5g0R/EOEnFgcxpXfoeDj/V84bAURU7B/SF2T1ffyV7Q5cV
uf8fKJ3WnB73m/FDM6J7TSe5ooyvnu9zljHiIhmm0LNm8sULNQOnLMt0zP3YRyY8
fGWcjxW32PzEBYpOujVgE8mefXO8eOH8ZEEM4+Bqd015Jiko+WpTxwmphaSE9zPm
ZbHCKR8NB+LVIgHK+LGCQ6BpYrye84AdcR87CaLK6JlnoTCXiGu62WvA5wcBApx/
yZxN/dg7vWBHWu3smNXejNx0zHQ/Q0/jXOiz2B2JIokgEn3lo33IIveaBHlGAa1D
4YR+JfLceuCmlG85ahzPd2oNbJs3LKwip7eqXJkT3RuH78F+fqkDOSNeXjK6Spc3
pE+cSsFvBPFvaiowd11HM5tzENX56n1Yepu47IK9fcD+iP4/WRsUeDq7r0xyCv46
tzTA5/x0L8sfeq43hQhiKCJRKfHvLDuOEghasW6pk08elX0189U/crY5bRVJh7UM
8KZ5vUyuJNkr5tGoO/Hur1lCmLTZzHvdT1SkFgKJHdge3krSINMSzc0XFuIX/yPr
4LGbP0xiVTAlmCRyDKejS5C/AN35J4E3w1LvRmd3qpkAGRJvO+i51kBFImqY3Brj
3fFVa+9EckAiplMb+6KCSEOtmqDEDUn8XjGy5Owr9x2xbXembelyuLE2WfDYWEmT
qMeYaSvkIzY8IL7ztP1CwApKj+zwD5HNAS/QOvcUq08yqDNdiJfc481RG3fz66S/
71rxUzNFvN8xR+/y5VqOBjSa0jqnxFLgr7PgG5EQyXqCieMJvwvq1W1vaNPSRe49
Kk+8TWrwg3NpK9tXixBajjg3ET1HwCF4tPiSyP0QW2ZBmWgiVOUQhg5RrnXiCJwP
8W1xfFA0Q9hw4GSrHMHGVvd84Er3abOP/s97aBptccqcQR9QMoJ9aEnFZXZEvI79
PiO0YkbcjJJZP0FwPzdYivMl4jjawIHnf8S+9fofjWZIeeG6YM8hNvzzYHH78p5m
LrZVIhbUgIhANGElsAroWhRXJ2Uf3xast818hSsp+7wgCAbzt/8Qnah/qCgWOaH2
ccaa5BsZn+JOugM9VQBU7riHwD7qp0AM21rt/yhmCwPWdYOUpz9xRRY0f3Z+pTBL
WanaQGYnZDodRMGOA9N+lObGw20CLUrN6VIC19DCwYngLbmJvSXiwRibM7yan3ix
Zr4exIOSV1eQSx3BKMrsOXL+y2xA+O66l24YqGDkn1ts/G2TLMIvDpD6zKbHsFsG
4ol4PeP27QYPuCq9pCsx8OZaEEq3PoGGd2Z6Wt20hirAYlATDHeq0FySO24qwmNo
Vnl2e+wEcIml74UN+UjERPLIT0tSiDotvyjrRzUITe4gnLKsCjRq0s4rFjMZUdUK
3svnLwxeR7WVputtCe+T/iMo0UCdU1P4tEmuhpG8CwYblbKQyT1TPAD3Yhu4nhWV
rrq0GedmH8Dnp8cuA52mntBMkqWqiuNrXoWoO9KICahh8e99s41FenWHgHNnFaXd
Gy+som9QoOiA0Z4RvEio/DohocGMlJbIU0Gqm9jvxSE9PPgKzzr/+/Onrp8bAqXb
Ri8F3YgTaUEDkY099SbUM4NfxLRZ4xkcSUz74195cjEkWaQKiQEPO7t9hWt1sXw1
VUXxAsF7EQ23Hyzef0/Q98HU9/08LDVpXywmpYAIRP3w/JqUsYude+whFiUhT4Bh
q8vF1yuzK1eV3FAtCPBNFsUhF0ZW1kuLS17/g739KeabEWJNC1dpW2fExI9x+t5/
H7i8Dvs1cEGO2iWw3DKvh8711FRSJRQr5d9/mvBkvFBaf+myoWi7kbbcbU5zuGC4
HXU18hdrSNVCvy3I8hcN+tZrkGS+QM/rOsrpyE+yFwq5/+ESnq0m5V01xB2uoraC
57bLa9pT/S2VtRJc2WiywhD5/xhr7DPen26a+ZqzvxPoBlcXNGKvXCeUfjn+dXc4
9KKq2mROejr0F78HfaOOsexbPONbn0tSk9mjKKp5CcHG/ek8RBETHb8Xd5JOGPBZ
IUGdS5hpCeZ5OI6ytKAnn5YvaApX4MVF0gVW7lW+mXLph23IOUl+nxpwo4zTUvDW
aUlRwjq/xGcTN9qwxbsYg4bJ+hq8sLUjVpD7bmF5+V39UCuUhz3tGnpDjZ6+gmQ4
zysG/cTPfWyban93oXZR/low1Oc1W8t8whHtzF0vkLgO18R0fpy+YGi2ge0GCpmi
rwrYU8xUM+EkwV18k9Ky2GXzWtBLogXVSXOx04hP6TwHr3HW99isS1yW9aGcFFR1
kCEUnuCaqIS6JbKnq5441uWNFHbh+KABYUFXT/epCwpv4WI1/SzT5X0ri0laj2zy
YQP9zfgSgVJ2iWfwiEi1wC/cId8O2URMuc3DvG3kV8T+f+vmM1YF9ZNOVTiZ/4G9
Z0nXVKaMG1uH3HkabI+fitSCMeQY7JUqfQM1YFV1w6eKx2x6iqAzJHNRAIRlDW+c
EwSjeQjZGm97TIAF1H7au8mcJk1aCl37pyrlR9fMC8nEmFxuJAynQiJF3AlazBW0
1TMo9zi4KlMzkuYaOwteczSzZREU9sb+DUlld2IvSw4G2wNuntiZKJDqjS0/chTH
FXH/+cqgYdcULVWRV1LZGf9LBcvcd8PFs2B5RxyReLoUYUAQ2kaeBGwFuhpdlzie
N9ycb+fyEn+USzfe9WHie0XgEF5IEHihc2HdP9v9md8pAUL7DFQT2dQkWUvaNIN2
jEDw85ia5hrgJ6S6+PLfh5J6biiMX1sG8Go+7CO4lKZRK9rUyHwgV2Zhfu/LmmXL
AfmyybyoW3z378UgjLIGropGtJNIyNsK/XcCxs/DY44R+a4NSyg0swNKziwSft7H
YnaMN/22JUKYEygmmpUkXXh/+DBHg054TepIALZpxpvlOxgnsz/bQH86YTzbr1m6
G1d7er6/eZ3msw8i6x13Dqv0H55cYJ68KogOts46xsxzJZFNmQyKtZS0Fv19Bnkt
sYcSrKNDNaPW5vIM2McYK/64g63Iw6FJpTlPAVOQgyetG3PMnFWJfDL1C26nZ6Bm
PbY/iFXiFr1xF/anyA1hHYJo3vzhTM7cYeUBtmjDwLrDure08BoD+SIMgGABESaX
W87ByGKmxd3KWBwWJJ54MU/hLUbHpYLRpmI1Zi7d7fZSrYiDjK9YUFIx5rUYmKhM
PKUV8zdhdyFFrjH+rODHqpN2etpRgayFj24r6iecuX/DxiEc9bi6igyBh0RNr63H
1fJ3a9CFuqipgyf7y6sL1m1xfTrbTd/me7CpPHA7jNvLG9H5PUw2CXZCwGl12xdg
A1Ty2kkmC3iddZ4gQhQlGi/KvyVHiuvTBNtbmR7MiUHt+GZU/lqSmJcVLEQhb0nX
EyoJs2eVG5Vu97arjLv4POp/D3Rc0yz9b6SPgbJ10jr82j7HPruZCAeYiEmP539A
ci+E9pcLIy+idJusDjsWbeeXL3jezHJ5mEbE7UYLye+wmplabfB8khSTZQVFRy5d
9e0HmIi7qNOPy1KyX0fEN8YzcWr4+0RsM49uXG1PGagWIIJWm0v8N0ePTScI1Cm+
sUppCCEUFsGxK0EOFAi2dCjSrpIiCD+L1WN3k0cuDGxX0U2uANXZ6KSgrA0BMR7O
uwQkRsn8yu5SLNWFUxNdKTl1ricS/9TqjrtrGa5W3sb/4QZAYS84GAfV3zPdcTHO
0S0P5dq3vj2doi2HqOsKdHINdFHqs40b61cxc3NM2lmoI57vHAOukoi5GUGc16VG
ukAKwR6Mh/yN96dbTV+Q2wrtry4vIXZlQDgFkfenDYi6ku5tRNSOWe4yzMa9wcvt
AoW5LdHkaKCViRVgUp9QGN0DbIe2Ws7BrrkNvk2pAATbWgopD/q97YF4GG2J8wTp
rhPu6zrW6wx9xwPphctXYjk/9r4tZJPOMNmnA7N/D3iu/V62Qceaq/W/VctkQEEL
fdtz0DriaDyxIkJZkx48ttyzUB1aV4UkAiDH/FArd7xVXwxFmlOILzHOZgKxQpaA
+UVJomFyqzBVFC4ZLcWRkP5Z0aYd16pKT6OBJcrGKz1ecS+Nz6ekq/0/mpT3FxsB
6gGk2HbWxWlb8FmoBQW8lAK5xwvP4BxwrIsXTS3P/YctC0wL8uOpXcLGoejf6CIW
eFWQ6H12bHE0ElH+F9MEQXQu9ZZJk7zj+1Vzw0zguMToN0Z/h2XYTOXr95X/jO5g
vT3zwtS5WpZ6A5vSvfB3aIPvxQjUZ9XYE+iI4iNjXUbF04kYnScCoOswd0Dahiaj
rMZbCPu2JqnKgNEKurKCjQj5qbhrv77IAcnjh5GESLFAxjW6XmckOmXybEIKkUAq
NhC47FuG4sAakF8HBQVsmX+8f0q9j9+ecLCavFc8PJyWr3MlTlxzZnX19otVXpuE
FO1iW6UfrqUlh0SXWB5IdGIZ7ireZ4chzoWYtdwtKgSu3txjydPQdepT8a3Q0A/h
EG/qkTVAtKAk6MNhy5nzn0gWgY6W3tn8+MwKtDmpbCK8sS65wM9qUm1yAW6QxX/W
foKuX0ujjgLN29ZvDWDhmNsCbbrDPpMOaGqKnOYf1JrFHjK5odhS5Fw9PTnV0mh2
aVVX3sOztndK1AoZQxKPDkzKdG0bkR19TeghAiLJgysyP75pT0wrxBRQYau+U7UD
xOhvRMd9vKYXRlCgJKQHH5OK6pUHIj9Yfi5tjEtc8+nEpVhtOn5Ygf9A2ai7oHTN
OKWrkN+3l4RATj198zrb809NT6J51ziQaXf349tNaWPzrm2/PpewBLydSrUbdf1M
z0w6gC/AjPnwUNXnrCZA01qYCSkX6ooIP5Zw5ouUjtIbFrRRsW62rEOGLsbZjNjW
2hUX17IJaNxekYV7cR2O1fQCk0AaiXxJa8vLy2Whgyu9vKfbn5ogq4Up4+lTQgb/
PYvZkSZUXUD87kNKCAF/5RkrOUKtCc9d6xqSJDj3xr/YOa7JDejxeWDj/AeAB3Ef
RiOje5Wgc/J3Ng05e3BhnpvAmTgQG4Qgmp2VlQvOkiS2V/GTQdwqTUyS/Dy2i4zg
YPMWUUTAHrIrzgWWrO4HBEAQx/APr/Kvp9uwKd+Y2YWK2mplxVwqI+RRNh4ZORG/
7M86zDOmCGHSRLnMgOMeBTI3DUanHpeGqUYHNxKjtseCC42mhoies1QQBYKhUMfH
B+7AKNTnB/JGGloswkfAb4QIB8Jz/hGL9VP9Ki4qxb+P7f9GLwSJpNHsHP7RCa84
m9WxCDBKNOBsn8KEy9LeEclQHtgc6141w0t9224sHItahauoqGwgPXhHtin35Ojp
c+Iaq2z31tIp/lWCuYUGEcVoiJxofx4QDKMnK7/WhARqQaX7m9DNjl4km+iESZqJ
nOZLb5NdjKYfxLuoa7dCdy19rzInjooVhgstf9TvBjjnDqukTDCOOpjGslshek0+
9KjTQetYiAapiOI3R+Dut0XMPxm/8Fp2grNJnU1GpVu09NvkGGJOHHo4LKlbYf5y
eApb8/7kl+DtGw5vOX1MxQfwe2Iy9stjXf/yzQPbeG4Drw9ANgLFy3XaQZ8/ewyB
/elrKLhyaSZ0bWSHz+p1mAzgUgPrk/qsT+U5KsIcrlV1xE2uOr5SAtKn6xUJvr9X
O0hUuXPVErz8XEIwI9ybKCJc4NQZnIy5J/xvYnooexLmbHDHWEkA19+8DhVI35ui
8ofDlVa7Rs7y1aEBRUSB0eum9HQ+fdxutaEAL02Tgo4NwKuh/m7EV1FOPLequQqK
HgCpCegHQD4oX8caFf3Rmy0mKBoEXUFtsMuQDcKKCHLTkOMdxOcT3xPV0vRGURip
MDmIbi52UzKD3mGoppr/CPuQmkxjON9Lb/Ez7yRVRY6cHt0YkD2Lxe22A555Ix70
IMhMYfrb9bugklTxcKJrUjg8kfJgO8bSl88IPIDn0wjYGz02aDmXDdP98MDOwGeS
yMb7vaiJGdLdj2PLaRKj1ILWvQtb/osn+gNKwBY4VWOGD62Dx8/2IiVTDvnqckPr
V3In5IktTdRW3ts+gr1WPuq6F9fU/WcWodOAS5kOIwsL9U2r7FNYoPE+ToOaaXIo
D0u8GOzJRQL9AIkVRcBOimH/cA5fqI9PVDNQ+po6jPm+XAVfU8ulhR6p6hRTI30S
88zJwrCYBwv/r31IZJJk/+NxTA35+TepeDKY7+dhesYDECfOtmmr8w9cCuuXJKDS
ZSC5f6m9/hQ3AZ+HX5x9uQILO002gzmOiGgfXADv4EAmu9liNJOZw19aQ5YsNCQx
z3FNhohvS5vqxnznMLqFMkj+LmO/coXD2R8IYHSRHZ1ytyZn7EVCUcpDfiNnAUmV
Sn1Y4Xmz+TLaH0CC4Z4TI9FHZ6x14R5ZtVCt+6QS/T+O3Sa7vGrB5IeGWYrM7h/3
+1ARN9wCOSSCi/iYC72sZKqCSKvLBp7PiXvElYXGWyK/kn+4KtATzL90yX/BcdHs
g9GMm/XCt3EVM8EkvJ6IMamvTOKVZQAs2RL1VMxY83LarZW6O07juSlK8bmSpojM
GzA3NT5WxXrvq+srMYZwT3FEeVzo9JwKdBangyjJguB+WIWSnTWzt34DyN7UP7X0
WQLEa2I2rMYsjOW3SOg03UfnKaupCOxzWpUYpH8vaRtrmqylC50DOBHXs6Jy2KYV
X0kHRwImjAKFEeoTPfLHCvnaelNW+yfxasQzCtmXOx50fCsHZL2g+W6KwcziphXG
m2x7uVMm/oSwWVKWXYf5+aeEzhpqAnq4YuMGhzSW7rJKm5hDKsCrP0rl+nY/5amd
dQtwh/rflqLa7Tj4rByXiTaJ0jNQXnLsdqqYvC6v20ZWtqdPNz/8n54gFmgPYj17
cbvjWYY1uIWpc4G2qFKZj65XuELLKSSMeI1mdHHhmrQ4wSEKP/gQITRKkFjcwu7E
TkcX/6LiyBO4fOnaXIPMBWoaGemLR+ej4kdd6IPQkRJ0KdIwd+RF7zE1YCZKKLzk
dXtVxqX/cWc8/kuh5MGx+9FPbcga1Pe5jn0de9jsUnZpdlshK6t58Unjq5uZMIUv
+I5W6zI748ND05DlrIqNbhOarI/c42SmcRHyrjc0R0c0vuKE7OvQ0KarVRQRJiij
XW4RHZ1bs1ZJXtrGAHJybaQ1o3CcjNqzq1iclr4goxWkSKoZrmgfGlTnGL21Mm0/
7PPuscIm6WPIPpmieNUw/9RF0fMn6o24Q5j1XI5R95I7lGozq53leIg1pVmg2Nbn
x5q5Tjw+K90HJjbvRVfZkozg4qWfjx2+p6FTFDJ3+FRMLK8gwzHv9J63S4N9luC9
PWWGEBDmh1YgNnCMRJ7oP2Z3Bm1zoPnrU8G4H7leUlE7ayUHs5OsSzWWMxBgVxUw
venKtZN8kVDxOQNxxIN8KJqKKe43dCb3KstcQb7oDO7uHnhWPkxTdec/5i/Dp53H
0bAIHp/p8bZfA9pXiXkL8XQ2ls6NdBEcLO7RBjs+aC2Mh5/oSp7MULnoM0eg8g8z
cmkrA9Tq7DnXHCAcp+pJeLhzzwCA+kLZP8jCE3MaJzy657IRz54SVhKdpxVYjLoV
dVLDfBDIeP3v0hHwRvMkLZeWcW4VHKeponBqxbywFUW3Wk3Huwkx1++IcRV8AtTM
bgzl/wPUmbGHIZwWq1SWRULqk6oLm6X3j6PuuiltfuPDpQrACrzcisk2frghYkMU
WCmvwdvSn9gm9InjWoewiE9Y/5Ro4ho6TdOhSDqLFjlHLy3iNLhYkj2weLn8rEoj
unZGPPnj24lwUN7WFgfiVZnptVse1BwDiSh7nzA08wOGJpdO5b/V6sSPdZYKH7Ep
RNJHE94w+aPXZn+KDfD2jA0qdS1UaFfyDZWKdwzIMisQbLHwyXS93B4ZLDtavm1H
s7YLdJtqNYWaY6SEoYLFjDFV/IL9ZOzZ9yx7bsMCBbaSol+5sMoJE2aTPF4xk43W
4JdAJb+z+vMiKXd6vKN9qHSfXaH8Bd/F1sKQ6WWIUNIalx2XVj2q/x9G0W+ITc+P
oIM8J4Cg0XrQgYqE6lsZhBisfCaXkiHoHni32EXfMGI6uxWv/j7spkdZ6jfO/6pW
U3A7jK8XA+evN1EhFmN9f5VTZrsQRiSfrpShjXAI8M2ZQSGjti40AFFugaacu72k
f8nZR20sQpuKr807nBpPDU0i/iqDbRTA/4mv4GW4Unu1uazXix2h1rnUydThH225
1+8cm7LbCD8haR3OCLcgw8lDergq4at8DIGMTGOHNcKAQD69ZEmLDMCQoG0Bdke4
3Y8H9FE81zBMzEei8vmf2feXNJ3KD1ONMXLcBUGozuChfq+jBE9dmjyiiIaJzmaq
zzmKO7R3az62GvqrEA5IbIHm9lYcv/0IowC0rUlZaKBX+qAjj62VbBSPv0uHyW1N
YDA3WwVtwQ9SMuiZCYiyrW6vHV/uyKHV8uVWGzYH7I+U103+/Cde+84uOhOey+FR
W53ZzcmxhXsz3WqBBT/RKHZwqMRmvSwuJX9TETR9ClgcuA0VYDt363Zk5VNxCMci
2T5iFMFVvs3/879Sp3xuYBoZ7KpPwewoD4Ty+oyR846GUpBNuo9i0k2ziw5evQaL
xQjNZ+2h4Mf5qbiC+MTe4GN1SBXVdDGJmusbbGtoE5CxVgMqVka6VhXCavQZEH47
m9H8ExUyd6YNp28CWyny+eJDQjKhymz5C3CRyiVFaJ61KVFdDE66yUEWcPRIlhFd
SdWwCP0hHE2acCeh4PVLE/GUBqKEnEkddgDmtytmJUyFvsf5OYFERHB3SSgR/spj
4TGQxCR7jUfD7AERbsSclXXNX+FrneSeXsvhfHcSkT9Vz3oavHEtqPJsQTpjQ8Oe
kYD7YNTk26lnhe1ubuEo16qlXkGrMILxYBDKhUgg9CE0DbpuktMlCh+ZyCEeo63X
QPEfKIkk9grOtcafXvMuI4CQPcZAYL2EzPhkes37NnBcl22ZxMZD+lQ+6MbPlQjg
vMScz3uoBNB9HRkx7OCe8Le1ghaucQxmAdKRfuprD6C3O8OkbWrWqkDLlCYwR4/l
4c0zmZ67P5M/hWbhs+5HdtRN9ur+UrVfdy90dRifAhUH2AK8XLS2yCiFnJPhboHB
ulkweQwY/62hBn+onHYCDNDW688qwNz41wY3yWHuoHA0B2qxBeIDPduxQkYmZdLi
KniZ37BefXZL/818utcwvx4hINu8hVnaF/vEXv6LoolSYyfbM3MxKPk/KZYS0MFV
cjS3vieD/7Wlo6uK3MSp/FfDVWBWeproOfxYfRdb/sX1vIWPNRLnIwgOXhFIgNxF
3UO5RYBkHxOguYFK/CG1X7LHuTleERBolBeIjroGXndxwIM3+iu5HwGId1mOgylM
pjK4UwF2l0lLtgs/QYp9oD1cAEinNucdf97kxBIb2uJe26HVT+tv4cWMwSDFMwrm
Dhk3z8moFb3PBKarEuwC/oCHPMHVrZ/BYtrlromVidCqZ52T05RdV2AOrRXFjIcO
/MYIQVCg6VIjdk4oYSkxCf1fnimyoGBXtUpxHkJXRt7W4xM69k77/56U5YdVRQ6M
rMqkBil/vWj8001fYs3anaIbaRVOtHmt0qBie8fBf5Quzb1UZBWj5SEpoG63JmxR
1g+cbWJAKcZIDksN2g/G9uba/02Bc0RBpabpHdn1WdBazQ4mNozkuFaFDc7Hq19O
OIFxeNqD2zde/0YjbtXdwT87EpFwMC5clt860h/Bt/g81iKDaapyhEUy295zIk5Q
nvi/W6tSw7ZhmiTiV2SzaYDHilyfTUjOoNjjdBnD0z8tfvu+Dy876p1R3coiOkAO
RIyobNenvreKMVHK5n9tIlKQ18n0u4r13foNHlhco3I31AgQ9j20/oVXILzXEVVu
kJsN+O+eUe46j51MimNQW1qlVE78LOobQDWJ+sqIhdC5urs+jrQm0GZe3pupmcoX
tSi/ZMqcOB4uIsueLAaomUFCJvYqPC4LVBX14znN6CRiYaBlnO2cCHHaKshzfEx3
+bjbI9EAnK41Ak/rbMCPOzM6ug9H79Mj0GknmQVKf5R95J3xfBE2VDhRlX4/7BTo
rnoPOcqAS8IriVQKVwPDHh+QMPzLqtx7Re9u4BJJD+NVgWmcj0pAKpBOLpbXqsbg
no6qoGCxO1Il0LsAUPnbJvgalQbju5M/TMJrWdG9Jn4aSH3GkQsg9pJVW7Qu2WDr
ybEsA+UPp1Wa4TylR1pTUan4EQaVCuvIL8P2Ee+XnOqhDrir5DGMe9qIFisEn8HR
rw5bYqUZ+ltERLG+tKEEt6su1Qhc9z78OJaFLgGuC1LMgSSPy09PEJA0nAAW6YWQ
McF9txCtFcCSfz2DYtAZuimNCQOE46y9pCrY3PCYoGVHRYkx+He35KNl3L6I764D
dsxcXDn7f72ikpVNwNhQ6dhT12QX7EveT0pXyV6pgv6COloWun2d/LYz0iG/gBdz
WNgkz8OLyh/h3fFmJkpmg2AtUHk8XNpjelU8VI/z6OmVR2/cKOK3jtIb1USPdT+W
il20syxeGYrmWSU/UWtpszFFHFTTehYA/GhB/6TnjsOUVVeK+1reEpqhNslRidDx
P73VaD+XCP5wn8gx6FB+BBAH99HEvRrdNedZ4rY/OCGxiQ3BRmc9+ckD38Rha8EX
bEvuHz87OIKhRtW+2v36dye8mNdYWGom6lQSCOgg3QYkeEYWP+JXdazIYocam8BB
LctW99t8SbO/XbGhx8RHbcs48ew7Cs7ddktOrvWTqwI53kH71weXMKC57Skyjs/d
0nq9P7MsPxzgMR1zroejVgf619MRNS6yM5uDZg2xfhudd8QI3/hGVwTH577Y8JVc
v3ZeQclJyUtXR5MbJQSAVGOY+fheZWU16kd4bsFLFpXc8nesMhRaO6SVGxlhdIij
4VCZ7GkG+jCXkO6eKsnsvjdqoG7u/6aBu2i1Cxd2SckEFu2whyXChG/HT2PR/S1i
MHpZ99mrvZongdKf9iZp6WHE/JkjLKPr3yBgeEKPquiv+/mNWObFWYpvPYkGHqIx
IoZlO4jaVQVLsnzsKNm0oh35cg+OR3pI/dvWcKNzFdEDXVZ4NqOig3EpmUJgByYw
aABz+3V/b55xLu6eFxa0xCDJLVrXbSE6D/OpqNVLAlb+r7MwLLWVwgMH28Mv3VHF
DFTnPeMG7DJbeqGeW6MP0qdNgsaF7b8ta5PUEv3V80YU0HLUmJ5YR45c+uDA6lLH
spxDvsZDIJ9MyeAX7PktC62DChCBpYYLcJ2crMVNZ8fGRxoprh/1deZmS+hJNvFy
vXhORXYHWc6jpNXfnHI3DI5uVxxQvcJ/eLVvYXPrz61ko9jJzHbmN82+WgisXYhr
ukqp+Zebno3MKdsfuNr0U5Fo29fbNcZdCHO4Oi7HOfFZeFCfDGEI8gYu3ZhcNupG
rxrBP5BTlhu8o+okyG86o4YdF7GfAAKvoid87iDXLXR34Qsdp8lHVeYr0jvjdM3K
vLPCVDF3xxcIYpsl7iKOqrvTM5YFZFuZatxZX4q2Ab8E9ia6/ZDZhE1+222r0wIM
D2RT62cdW4C0MuUKtkvnp5YajqTxIh/w9f5T2fVr0OWeaU7pdgCrVQJWbJ68ciH1
mZI6XjXzeici9hNR1WQrPHTIpiUmxDeFLe0naGv2fUJlJGSFx3FPElqSJokJbfhE
rtcp03bDmZ58UJCNo37oiqLksqh3h6Cf81sc9NBgw/IBhQrNRWEx1kLQOQRhKoWt
LvQhBp4LirNDCF3JBEHwtu9vc7V86o2oi91h+rL8x3VdByM54r0tAR+N6ltLg70g
MkAo/5DgLwWiTi1PPtnzMWAU03ER7D0liucaJB5Ft8y4qa5exNDT7wQzwx3mp62J
OktXgPdUdat5Z1lZ1tgBvSAuV5mL9hESyv5mR73ylgO5/mR8veU/mB4grtXl9Qfv
5lzzpBzMV8LqiMdE67arlvDxop4z5YitDg2q1xk0U8y3L/gxJHQ5xjWdjVV+DKfg
Y8QEJzSz7TTr7O+l2/OjVidPwUKgAEKLJJZYZJnWatVGRqxe1MvGS7X+5T87sBdW
K470gk90HQE7xk0bJaW6zqtbGGwGDKD6ap4ys0dLJQFRS81/+PeXNG/sL2H+llsG
sIIJfSiyVjsV4wSSc/EA5j6ByPqaYkhDOc1ZkuaPGpGqYCiKrh6ioR8qJfItovI9
NTAxFJghUuVgsrjr70JNjVJVdO1MOeMd8ofshUKt7Iv/nrTAwXX5vynLAe+lXYS7
PUPUFK+tSDQSVRDbOFNHcRJrmLp/HDasSDNbNFtpeybHx7wFMSW9VStu9ljgFJzj
dTaJBMta/dc5p815P+slkkG4zMBHECR82bantiPQkbl/Rz5uCTY/4y5JD/EFGDo7
1MpMFRS26FWQ4w/CaoCyCcFn7vR3Ys/ztxfcvKf6H2dFAixayIKXsE3roJNAsQY9
ickemDJuXwyIvkIYF3B00N6Ikvy64ButGXWUm3k0k4kxaw8deFEGZIVILBGZipUk
drvesGLaSAyDnkpzCYPnOoU6/nd/0BknLG9UwUIZOhQyq2umxJqLz9/FEgp7Jb45
zrus2Jt+UsnJCw6gFMG3qsEnlDej1anQ7/gHQ2ootY9Pmsq7uT6h96VBadQ6CftV
l7q4sBjSFTv4p38XKwCN1qRWHOKrw5g0qIfTU1GhdKf0Ea5by9P9AskC69AVT9HS
p8oYEmXjdYubBgIjcA6StsbGepYsYRJ1b3YUTgLA75vVyvz7aBwgIzozx98gbl2q
Q00yFCEWP0yRtvUDiGhe9CKRMbJsT92pzCo+5xdpkZNuBshmB9brj5x5KBy623C4
I0FFp7qU7lUiBPn1v94KHMKAfpV4vq7ZbBoIKuvj6dyWjwudV752kSJjkeQOBlam
oagK3+tfwHYTyJS7qB391tZ2478MARd3ZvVFuJ5Ucz1AjW00Rlj1Z4CgHg99dgoC
47m5hQGMFE0nTbZ7Lq+AfUMKNBOS3vA07M6TAWsHx3n5jIuIQlMcj7rY4oY843bO
6GyyPT2Ov1NP2R3SP5gRpUMiwxms4KxrWyrrfHooPp8RJRYxuic6gRP8vb8SkeRo
KOZryAyvMl0aU/jT8tN/plW2dA5Ig3OVdZmZSYjopVjM010qQkwMM6i+ZZTiLTNo
DY1rDLxkGlb/rxa+ZP+MNgCM9ud0/OFFrdIdDnRicPy2UfJDeXeu6KPnhbwlNlSW
NlBz9NQWPxkDyAF/w1DASUCWV+H15UtfL5q3Jc7dFlVwJi5SxliQ2gWRoBu1h/Ul
/KCgWrChreoambQduUc/2c3tIcDf4fpLktkAkaKczcR9XpGvj8fYUqodpR9VzA3U
SK8Q/yayyQ1d6RBkUPwUXsX+OHeSVn2Hj0P6eWTZZSn2+C72W0iGL5rQ7E+KHMZF
V+TyuUkWjMVPXOHABu7MyqpSfHHX54DJkj3NNLDytKa+ren6BD+2Owa7vZFrwRyV
qOZIITYyb0sKb4PMjxAChB9oJuX8Uf+ExXNK8wNKYqIRpBL7Al5ydl68BbOY6qHi
o3Ku9TiMtMfZdYzUFi9N0u0bQasoVpZR7D8PAfeP1KIulIPro25JPFLTWQQCYt//
Ok1SThcxPcZl9j1ql38hsdDW+2nzb3TjPHwekEIqzJn3CUq+Rg4SbOiaAcYAZAZ/
tRwH/fCgkVRu5fLNvSPVq5wpsdBeV/w/Qrycm+3rJARfhvvI9bqCDcmcXejxawS0
uawp4WTkKL5P1C5rW8ogERm6XTU3p4aE294YZdWyarvUwroWKJ9lNi/7g/4N1s9l
5gXHGOod9ctJ4aQsmLo2xvBcKERADNW0PbLwdqPQFLzn5dqo0s+nb9UE65olJ9Y9
PtURrR12X31PT+2u0RewITiu6mgQLjGszHnyiNxzxug/bEtsLQOBhRDRKC+qLMv1
Br9AH4ikDX+DhwVDxufbJYejjeFdHbJhOWNq2zp+Y6YmzY38RaSriOhJ0IUxWbIi
C9Yopo4LhIm1rGoabfUjT+VVrMCU8OoALqSdn3pxZhQjS29jJgY5PzjwmcCfz+Ru
wosPgKDqqtrQrqOnjotlI14NzTSYOL/nyGcNkfE9AUKzWVwvWr33TvHDF0/sst5H
6Yh2MbvlqTsDx7F6oWnkQ6BYMtyyc7OE1dv8nCFEDTHmEHZFXZy+ihZSo5yBp+/d
NxzLzS/Kqb7sfzS/kAFNBKM29X8RVaF+ehB+hY1STt0NTDWqRTuZq5vcs+WSUD1W
fERgVO38rEGx9BlaK1WcZ6TrIimmfDxzB4GKuWzmbsM6+XcFgvs5ERPjoE7qgu5O
WiOfcKiZ52FFSrxZVBVf913km7S4Vu3PLRWbeqqPUROXTv/cMGTbmVUKTyZs34Ha
oWQmk3xExbpKXVWa3Z+7byQRPukOd+bXc1AASIwSzDJSXc/dKE0w+0efOg4GbIYi
NkDIVIa6Tbbj68JeT1r2zzSq/4DW7PyWlmd5LAHCN3/mZXWHog31EQjvt55Def/g
rnDTj3bPRdMmgRlYqzFQ7nZktyaRndCotH2wjLTevrJurUBpnoHETrcDmKWj/6VU
gfeLKm5n7LUe7GfMAdMzvCm/WZuG7ehd40+Nd3+6LY6MjL76jw5fq7D0rEmEzzEL
RTGLj5/gyql8iheDPIyIGlqxCFqDT3FDb/FHINmwHkmuyRqCMfQJ4skJ6KyVyNZk
lOtNZy+NJUIrc0kCnlHhtj0ThUvTHuNqQ6qSsfthRsHs5WG+2feVRhhQfua3l1Qs
y7bZyFXn0VxA792Ksd3EzunV5of/nXN/kXgIrwE/VwXFbZMNDo/s7vFTuhfeeVZK
iQdppUWTJz755I+0WhZHURZpCZlw5A9mqjCIEptSsg3/pS2MoXMI4cYvKSgmJVR0
5w764m9z3+zEY4ivAnNyaFoSM0mXAguBHItf395JXfUvLTKn28H+cnzCGVj52uwY
zRcKwAQcs96s+kmEYZmbcAH/OXcUJJKqpmFJtZpXveB3nIK7eGMQzVK8iNL1M3Ae
HtBLMckj4OatP0ig1OcJyQTV/+CYrDbeIl2QwCnRHxj1BGSrz1Dh6Gi1bdDGsPCa
BRzf9pVQk75MYhpldVCVCJPvhPLNv/Rv0dF48io+ryNW68SHyRdm8eB5vKDpy+B3
x6l8U7BmWjNlSevlwKj4Xyb7qlvo+AjsL700e2exHPrpsVNRB0EVwN9VaZe/uGTW
lM931MU4kqXdfhfVyRP+b1b/maw+egS3tatnywwNorjXJnejCUiq/Whoykzspu1j
H0MIZBZJG/zMeX+baLxm6pw3wIov6yeu2Fn+krCPHoZSPlt46p+ASjPFQVKhhIdE
d4XIa29GSucuibCGp8+MqZ+Wit7+jHLzf2sJIFILHuzuhxlucyylT0w4JMcd+BMG
/vUKdZ7T4OEIAxgHrNpgi5jd6rRsoQL5h+FxwKYOwbNqHy64MKcIngz+EIixYGR0
NkRcLEWR5bcVDoh/eSHdYG7JdYrbku33maiowtHtt3tQW4xhLu+Gcw3X7egzS0T2
fUszrhqJVqit9DI3tw6PnOKMk6qXIyPb/8GS1tHcRWD5XNMSc1XuExp+KVA0PNRt
pwGBGtiTbZlWtAwdTiSs2ziSsjwYR/pEVv/0RMZxg4Vc03NcGFaVVoVzPztiPho7
Wcddsl4CNQ9leQIz5qAMnOJ95mGZ3KBGzeOh+fZsbc/WCgximZlIxfqs7K8fT+By
VPnQ3Lnax7X5JRCislxYM2WgODsyH0n+/2g/J3wbSmoo/WWAiTjCWtNd8p7OSjfz
qFRC9Nio+KtvZSGKlgoY5DhYrdrk5IVY8i6CJeD8YkMp3gnANbodr/Ifm8IlDiuQ
VD4flFRHyOlboG8yTT7+o4de2ALJDbYwsjQgdAssvik0Q04pRiMrudRMszDnlE1M
xJYjvwaaNgZ+e9iqruBWPQYpr45OLOI8LCeviw6CFI2OWxT8lyaDQop8FEgjnGMh
qkJ/JRdIDswyKbc0Vo5Vf85vW67K2nzoimwPiGHw0iKJu10d/lKf3wY3SXDV4bbK
t6lQrVBsENMYfBBE0nyforaeqbSf3/NyGYDlOIza8XUPWt0AtiO6wjINPTI6Wu9V
/9TaIIa2Tt/ou+3l79v/vNDleKN4jQbRn3oxVDupRNgzgAsQzU9eMRPKaU41F57a
isGWo3VPgQZ+aDivntgz1FbwbKG0Dt3G9HSpeMuYUNHlceMZN4JWTgKJZPaW75Ky
T4T4R9GPcMRDGpQ2NnMqmUVRI9ulifHJ/PHwu38QNykr0c39DBNkRYVHWlblbsMN
FTv1al8NUNe/wIDxWNC3bZKY8hPhBIe1kXsXo+WUf03xKRR+BNiyZ2JV7DEowBS4
H6g3xpicj/S2Q01iscjCYCEOU2Hmj9+KLu/Yj1BrpAajOH7NdjpHTuaIXJp4svPq
n4u+JEdpLZPdr0xzTMtcpmoiBCeQAghOUMr0b6C6rBzgevNiWeVPnTZ66NxgMh+g
X+9dwmKBdzkyjGZ9+m+qD1sMoH/jg+HDUL7HnZTgjJZoarXB0W1FYalwVi3CEDnx
uZ658SUdVM7fUhzRr9M+DlAF7t8EiTWemvdzOW8qQtdzsX4igo13rszI6rgTBTVW
f+s26eQshNmqMXhVgLtwvZ4qRJ1hqtkiVzbli2//KOwi3phfngYb+baOTfBd5ewH
DuGV8Iay1bOcf9VGC1lTaF3p8joSJChGkqg2i4r/RAaTgtwxCu9nSnUzTJFewqKI
tzDowRrO4kUDK4LN/6ukGBfRqZPut76hc1NRqtcYSQhN+VhqQsl+qCDdU69G0l6N
S6lhOnViuiP3CMHQ3qq+pKsHvoOWzd9ZGSoUwEQ9jFi670v4ruxH5OzxCAU6As1O
Z2yvJDX3/DwoMa7D1A9nXO2rQpZUM6aUHTkQqZlhK+mSqTPwGpYDZ3DicNyjWI3i
MBtg2ldxV52eU+8ychzlb3A3wcvK4A6beAbdSJcqOIJQIJbihYKsfmghZQsGmK4p
R4M0x9XLzEJQnRVX8ann375zoJu2aPz42fZ19OiCzDBob+dXjoD4E73iAftN0JU/
pMCHJw7DvehIYN+e67fLq+sFrqzgqmQBfhT1ctGlhh9K0lj23jJodZPlME3sX/3U
prAFdYZp1w46oDfSB1nciH8nfUYE0GBcEJd5c0T8ObTs8KJcOUXEYgi45gVWzqPm
8ssfLF861v3gyFj+EA7YJ8zDZl5gc3VW8rGrMOQ2JX72dWGsNECxXlVBjJFH18rP
SUpXYjq7YwUUJaGqA2LvCvo1gJq8vk99DoqeWJxiIwhrQ07Zr67n+YMU0NBr54Zp
cRKTwk4cIuc6rBmEmSLYEQk9AZ1ml3VJzAGG9jNar79J4/0VXofDYaA2BXY4udNu
3H/05oZdfq1YWkWmiigZppDhrcT+Xocvrhoo67QuWYd+sQR7aJo6ZmfqVRwqC+o3
HLv3gBeSPY/KD7HOfYmISe9YCkiK+jSOhBHqgDcSpzNL6OIcyzO2bMZ+39Aw5bTl
jxwrkpurmTaEBZjxVOXLThJcqz3wiIOvIcF98cjk41Kn8Gm/k5Xm2VWO8DugtIPb
7nZnGgAZbIv3mOuP+EAu73hnrF5USnDe598QD3ffLm2VY74weLbTEsA64hNGC1SK
8XleHmVwTsN12gw8jXVony14qQnp1XGSQvB9xwNXxyBJk3jf67ctUcUqejOu+1cZ
yV0CM/2Q3WYLxwjLqZKJmx74IsZFdf4q/8H4SwNCIHH/uvE4n+j18MTITfQDScYK
f1LC2nC6G9DGuYGeTo+Fe5Ivlzdfo/BMXACYu5KQkDc1QC6uFq6AyrI/Hd4pqKRc
xamUrYFRA/Ven3sexYEP7wfMaQunqL6jzffja3wYXzhjBl88QcCA1izHcqFKLn4s
wLcg0eQKNxBcBePRDaDpN3XkYSQMWemi70vesnOq4zqAGdogCtMoTPm3V4Fgclb/
O1qducMIe64mLmmROhbv9yCvc1U+T9YxyoiowjrmbWksQAlYA6/MsiViEDDzBEtC
bt6AmHKTV9Nm5OzOFLslWYTGrZlN5Se1m4+1yQnAaBQBqqGOUxBXZrdk0MCcEend
75gSVcXg5qalS9plqhhPpckFQFWmOqG0A5Yigx1cQQgMuHoG0oKz1jjtYYjJGQ3T
A32GBtq0DNH9loXKamAjjmcmsexrZaIC9+oS5zwiDYCIfRAz80d8OHN9vCogXOFO
Ulcmq9PP6Kd4g7sA0v3a03MtJ2/1NZCeXUBACaGeI8BQzvGeJ+m3xTEWR2Z9LqJr
NCY4yHc30MDL0UWLJyhoCzNhKvb0SJSQMpM1sQDNxoU3O1iC/svWwfJbGZ9qwpNm
cm8JcjUOvHrJvJgZiV2QQqeS7jIWys8qZeRnw/cg8Zj7BH2kmGOdwWhvkMl1Z6kO
YjhdZMKDtj60rksCkqIoy/ePxCddnObXIeFYqKC6G0gmnJvOL9muXjmgEYVQJqz/
dc+M7RKZni08fCiMsRCP0xOpxA3CkQA0B+nGoBskjmQhVmx+8+yLs+BCqvWzkpoq
6BaKpCXlqNHCj+ixgSi3WizmvenzKfHjxjcZsseSm1jfKGAHmkdPtiJYzuPhhhTk
/P0iJkZeKUDbYuCSaKtalNsWuJYfnnmyLVmcc+dMsXXZgQxlhv53FqyES3vzzsD0
WHdXHUN2JY4c+OPqJK9dE6pwoGhdsLF0jJXmOMk5nXDV8Aggpvki3PzytSBimFSE
+2bpfcGElv6TvvP0XK5n8lURhgrzjvf/LiWZ9y87Aqz/i90bVV/sGAcU4MfbsC6c
isHQZC7dCeFTfG4763IXoGG7+dZtpUvrT+h5n06DWEZtQ2bwYlH0Z3npWBzLl4fD
B4BxE1ZrFyWfIxgEn02y8bbxseV0lajbeUq/2B9EeF0xFqOFx+qDIgw+aklrt0ZT
Qqeb81puvn9jlwFcjm9XVEcwv99/4nQ5qGSy6kq7OK2ryayFe/mvEws15CwbC0/N
8FgOOlNX7nXTD9RQJGUw7qKzsWRzCLY7VS5OKlVJzCeak+QQ/uNqIcZdH10I+X07
2pqEmkxq7wT2c8d6h0oZqOzRAH2Q40poyAYnp5V8ET963X22PEbPSeJQDocUTStw
O2iBu4LMJTuqAlS0mHsTDoZy7VsdFTkZkE1Ko0s7/uxa4T576aRgnM3d0nfXIT5U
sJm2aRWUVWVrg/b2CRtJ1Do1xikw/QosWjOCMRr2Xry2TYDZpJG1nEaFa1G/d5eK
m9I9OFsp7btPyyu0IkV3VZAuYk3FixKMIaMYAeXy3bZCtImiPRkueJx92FJdC78p
y1hc+Dmm/kSa+hionvklFQDiE0jAzW1Rq1pEbCdefZi/kxhQowazGnQkAELTHahi
KUWMwTfMdoSLRPOw88OupqaEGhJLCs8KYAmOzfs109T3IYNvaoF+4OTjs9RycB7A
v4toF5EJFY06SakJDF3ADQQzl8+CkIqrKQAUy3+NbKjrQ2R5i38Y7ZWgUb/sRqtP
y3C0H4FzLU3iM178sOTM1Lp9oS8d9JE+AhqanH9wRI4IE09ib5NTox3Uchm0T5NQ
yikd/tyxp4GWM7knIaH/zAKanastKDUPApnsK3LFzPff7r/N5SBqpUPTbNzbTyPf
xb84ngNXRHXRIoxajUwhot2VQYBOOOgJYMcvKq4LGjUZj1HKqD+KAUAmL1DY0wh2
nbSrMZu4kNfDkAsXOUNNuMWJ50AA2Q/HZBRTzYv+5S5f8S3TQ3oQkOm3/jObE/9x
eaAQgtvAm+9sG0oOT5wlQ5EWi8FrfXWJ4UoDBPcZoU/qwftiA1yNRnke/jB5MbFO
oQ8Zb4v2XK03u6aht8zR1g/L3F93FESjiZkwlgrR4Ans7TYPOCcb7LwmDIgd6+C5
dTOBjqAQHYqMNUPh6Aor7JL3kzRkVPY7dg+z9sNV/QjT6P1+PLm+cHidKokJ2bg6
wSFGJqK/Q8Pq5Xz9rr1jmmjHtOawFH1UfjWRZi54XgeZsEXg1IuJtVqH1EtwN5uX
XpQNyYon9WMdRj7cHVaoTShqgNZvs7ufJg1/lhzSMLPr+rRWc82Dvt9yUNeDJ6Ng
KxqGzI5TrHNpQ3072fx7fGDda2bNY6/V0AOXYIAVPQ/aTz/zUtzFS73ioz0w+B59
p0wgzpp4IhDprE27nViL7wfboTvM+FtWRysM/wQL6mHynD4AOUGyBnb5Q3DAt0v+
ohx6uuv2QH8/eV0ZkfuJ9ScDNdXhD1yTLT+4WMH+O21SxljTcmwH0RNGxKBZvIse
SMS8lsDIR8jQfSpEsg3695O+3OQwBOvMJwZ2aaBgV4IAxREjsfVO5GGFTvQwewtx
rrEaY1uptNhyK3d79GamhXq8H5kNYvCepE6QEgN+d5z1ingxIpQ9JoPz4pAZzeDH
iJkOIG5vfVU0dVku6/Gof1+PlaxfJek9Yil5OMP6TXR0/DcINGUHsOeiV2h9H7H6
OMBDRMRvKUMYoPWjN07sKbuJVQK6CwRlNTqqsG73KWIrcXvEOJ5oLRITzk9HDGRs
rix3o/MlEBj0EG2Yzzy24ZD2VU0QjH3Fj0MOqPiOsC3bIHSTI821YqW3+EP2hU2a
g0cLmlE6A3vOCTyybx8Khb7mkH4qUOPQVxz9M+1hYV/OV+M4KbAWx0nQtcqvXl40
Ew6RwkhXjRRyVmW9+f/Sw+vJEV5xmbhOkh11dfO8HAReXlYI+br1XPcdr98+Tx4r
i4ZwRtryZtCNpCj7rZ8Bb9NIaLC+FS64zB3LrOffFkHVHWAHHhieXxXhg5m58XfG
uCt5tKAM3UDEfGXAgVDzo04c+1UGnFXX19a6hVgDZZUePF685b2FTQ5SPWtNbMYK
mIpyFZH1B0+QNEvpgLZ0CzccXKNG4MY0/Vby9ZC1AW4WM0629gsZUpH7ybzblErY
VX7A0Lc9/x2ildFgutpx39WcGanf1BqI1uIQY9UKHv2/j+FDehoBGiOnUdySBclF
XyzF0tQ2+ZYwFtG1TcumtujzLr2FjkifBm/G5z5uxdF/fvlcl46fdmSCneykeA8S
rcIbGW5QR7xhtdTXrBm6mZFsZQ40JRdIjaTnNenDP2b33g6V1vTWLSMS4CL06nUD
dEAubbJraqkuMmCSMyKTU3fRWDq+BfhXh7vInvGWXFBp6wInysnkVCE271lQlmwb
6Exc2Yreq4Drq63U8noKLLUHHEebW2w0e9t7pce+5K7KlllKA9slDxNK1rgM3QX+
4WqT+3FVlXnsRjCr8PtV3GPT3tZz//QBlJM2JO7Sq60kanyOB6k2KpInkxxD6GuH
snt68RK86865vGxBt1vuyBncnqHyJluE7VC7/ystvdrEQ6mKqAIJ6niJPiZDkfY8
ciibNkHBMZR7toy8anmpcH3O28dZFi+GkRvkqM7sJn5M1sAgKiceVXMfBrT7UXrD
axOZeuQ6LIxv+rhsAPz0ImvtpYrrDNFY1i7i6lkVaKgKY2Oz7KWs6OJJrne47JxV
ah/PDljXhII/7FZCksOCPJ+GYuXSAhgSOA+zTIJ9nKJq/NxEtokagmOdc3a/nxHE
XthF/Oj2iwHQUj759+4pfkrJ4lYrLn/iyvG9NYxcoecHFP5asEhfTAjwjxuGzgcv
dil/vTyZOVoNVTatsfVUtDvc/vCqAdg4DTG/E0e3Rjk7FIN4kbWs2pS/f+k3m1Jo
Y4JwvNjWKZgb5NlokqL5SYvfeVvNC0Z2RmenCF95C4s+hcLrUV79CRwKZ6vn0HKw
Qgvz0Fta03dEMBnyH3650VB+67K9NeDU1hGL3K3pCyYc2xSIVEUV8D+VRmf+Qkbm
8hlvt03pocpg+kWm7XMXQGlpB+5cStrbxLP39B4N84nGl5NgnK7+AzNSTU4Q9+ci
5CMcRGgs/VXmrLuggjBynN+qMD73Ks0kKGJIoOaCtcsGM1wSzKXohu6DSU99j791
m4+jqMNXT/B3H0BEDYtQQTRI4daF82Ak+XAEsFntrz5AwRBnorynWqfuCqqhUS4N
bxXdc1YZP8Yr4bU4CiAjrHYk4dGZUlM8Fc/kyx9uQrNcJEut8h/b82A5JKYX42jh
roRJpl8IDTFtO964Jd/BOk/3BLjX8wbagZpt+XFzQj2bU5MzYXUAkLimKEQC97cx
3gQu/QdfdqfZbE34QGXUgivJOVZxH0Gq87cmo/PBsz9FcTFWtFzti5WJEhHUkOD4
x3fuNd9BnyeHduZBMObpHeZrr0lbyqk7EsphH9Xyh7dWebfxEh82fTFQqy0un8/p
kRyExXaVlhabXNYO80fpJjKd5b+3NOzfxxqqQObg9Z3j4lcQzfhLE+8swVprKzhb
mrh92joXHeStLMxZwMuIzxkppQniQ311+U2LGmS06Q1HsP6+yvLHCcZoH1ODjmFT
Ha2qNwhi/tNuyL0iQHmZe7sAK8oYcwLSj+wyFnPRvcYEWhDeHdY12SHQGONI8vQC
AMg3fFENyZuGcKOqSFcBxbIXUyRuXcCg0T/xraMJd1Ca9ua26sNiceIEoeVRiJPn
RVeRc9i34T1ktZGf0uC59QV/Zac/l1sg/EGOo25LNvfvpKYjIi+evbA/Vbvns3v0
bMpY7nTxiVnGPla8QM7XpBjbCH+WZsHmwc4Kt4WDUhQpk8WTgisuBK4jMQZp8UiK
H2l49cxVsU1fbWufy8v9PTsH32s43yTnStfzEsk9tOrCjAzvNaOoLLjYjLtqCYlp
ueE7luZGYRJIRzJUxxGLhAbdOVoj3HmoM6Nxymv4KlUp97ZzFujgrfyvHH/k4fw6
O/uF0hSHM+N3kohB6+7waz5i13PhPWB9mNB/Ma6jQ4ZrBUZEotK/veApO62bhhxY
dlRah4pShrTx/AEN7mccgyaw3MEkE6NsBvgYgDilQcmEet9znsSFZpD5XKyi0a6Z
oQpB72sLwHd4oaqkINXrzNGUi667tBrV5o9jeD7sId1d2lf86LDfxrxzs7uqI4pt
gqbDsC4i68xLrR96ShoJZxJWY7dfsgyP1hDqEck6NlVGCXUqKyZBnsSrNnMKfB3e
fdAInidLiiEgeXpwwPtJo2Tc5RDE41h/gcttT+42WGcnZDx8JtTQTFjGrWonuTkm
+rZy1yDCNT5mPQxyKtq/6F9ALfI5QQs4OVI/KW4/CsKejpCuKivEC+lmiaC9vNVW
hzs1EruKSPcrVpJ66OcreNrGpWduupCWcI6G0EWRaTDttxPjti2zEQWlnRfTK19+
6x2xuVXqQIbO9RBJflKncM61Zx86OkGFsEl/DsxoTIANmWsGYuCWdLYesgOiDZJx
kK7Ni1YEjCyIsoM1WO5gb0EwL5q9M55A69Cj7GQ2/HzRjtLtZEq6ihBN10UyxJbK
+WdqK2Og101ivw06WNb7UDuKIA4Juw2mYjZh07N9skdIv0AUnDJ92pzrx0l1nftK
jj0k9JMwZ8nKm5APcuCdbxbbEeKG9ORFr55Aa8mVbLc8nxxF+0N2/89lS8pMzaZ4
gh0KRqU3YJ2PIALhfHGDPugRLMrAivVdOYYA7qX26vmHFv19N85glAT9byc/K7nx
VqBIpnym18xJswdIwvor7H2B+5wzDEL8tnLs8UHLOL+fu4z8O1ckR7FiGAGvq4sw
cDxNMKGOkTl8CSvtZzvUP8uJF9GWvNTmlRti0/TRcGjUvt1+sBfrp3Nn0sjrgobG
s4hJliB6ZhpxHQ+jzmnNJVbMUBUkVtYnogdkq+9wf5yv2iG0jcUwtOO6nrGxaOXR
UcA7h7p759REZMS3s3EU4cVuG9YovTIRfnOimp3jx8d767ek9obEzMTb8ZqO8LZ9
IDROHBEPz2FFq4bN/kKTkU8ls7Mmh4oG3rGtVrKLaDT+RB+/TfM0yEmROHnuDyz0
YhIfyTzm+fc0fKRKr1X9enTnuXtsJzPdOFqi1SSpQKNd38wYwGTjytF08oXb2QeM
MG1ETasV3Coh2kOIrBAMZ9gbMSl0UJ5BiwYRtYrzaUCDB3cc5iG/tNu97mLNfSN5
XcaDFK6Cigw42udADtasC7vCb66XuyfM2BKBn/QHX6gf97pPPBNNhZK90Vc6Ia+C
k7gXlb9GkC1hixta+9QUP9bd+QDlE2BZVaFz/PSXQfYq2D7JRS2xBuG0E+gSVywm
4J7m/+j9fBRlPL3xZVGPQriJhyX5kOpDHYQoTMpQbhaEFGjFldeBSlizfLeS//Gp
vEKZq9Yoglk0h6NIo2viV90RXNGZdvQDWzAeTtwWA5W28MXGIheKETqXIRx8uCFn
b/wYWCjiCkovELPIjMzad1HMWHZW7OeZLDs0IDXfeCqllRjOeO771m2HPUXxgaoZ
D9uod71r9bB+5JTaFnpfjeApAHi4Ywl+Kpakb1ur9ooFybo/ICCwSFP3AOKjRmSc
0qpF9enCvs9NqNqnpapSDEVNHtllGmPZLsR5ZnfZIRe3TpE3HIpGPsq4KdqX1ogy
2CDbxLxYUTviPLFDArt0CvuvQtYvfLqAgGOwqNlUG+VjGYui0K81uFAL0ledws2t
DwKntf8xIN2YQLZVocPBUTikYj/BVOfsovsR3QB90B9hFlXWzFdbhMU+gDYGRPFr
unDox7LY6WsEwZi7kKnj3gFpKp28XJskY7mhfFj53PK5r0jEf7tFogoLfLVu+prP
FgxBrrAM9duDUSTlkRKZh/WlHilMlFeU37yygh0Fe40vadOqzxrjq9B0hEv4M//m
RNKT/II7CUQWBz5VrmBQwfL7I8pWYTfY15cAcYM/mfx4H5qNHRj+uCXQJA5ngXX8
/9jsSEkW3GZGItC2IDI4vSA+Vvci/gZxcnUiH7mM5D3QgxDGXMB5VN0Mi1Lu4OSW
Y8IvEaAlf0yDUN7ev8v9GQGV/mMhWiZiCF4ybg4/NrPnY8zyEMJjHrUnQ1WVsZ9x
uQXTp/Xvyh8nRowZS5TdGDXtXoS+1yAoG7TbTRCCIaj7D0NXeQKbecUvYP01y539
qwQL7zTIEw36FyZMaotQoQLxBMzNcZmRZFlq389Pfae2Sr5QayhVDYKFzbjEZpUA
PG9sTbZZknqa/oEEsNe8YR505uynvph97xbZwR7M3YsPEepJXDZ6nA4y+cRqlAnf
ULmWU4c1Djv+fKKS/zcM8GN+rud/VUt7L8njwpF4pPgu6aOumahCHAxoYpW6zfTe
IY7f4GKPjKoWkz+8qoJbQKgYO/o+8J+BDlDE+Sd97WzjJeuchoN/w4bNpmUvJTSV
RRuyq0/frz0fmufdzwMnfa7Gszh5CN5aOQWDQRFiw85SJA9EiVesnO3SpILU/nur
v3VIxLBN41lcvK/0YVP+IGIw1Hktx9FjtNxAmEAn0mJRQycQXWLEZWm1smacoqt2
V53DL+4xZdTDV9J0yQM1p6rrh/GLMqFj9Xfxjll+YZTGIkwWfNes/FHJx3wje7zF
97Hp6bd7vEprEIOKYV77c9VEe+9zZuwPN8W9Ua/PTqlBshHIDOmPi1aUW8uK6LKJ
O2v3Xqm1vI6WpYAzXklLwP0Q+xqDf27dxO29a7x6JZPLM1AXw7Jdx4oWZmdKK+HK
DdDplGWhWYqssgCfnbh0FQRcSfUGBZQCvPfs+LyRXstUMMVfP2haqi0vGnQGdZqI
gjSD+7AeCtTFhgj6hmjpHl7rgrdjWSfOAv0QbXqMl/S8UCZjutDMKcEn7TVwhyAU
IJLAmV3bwwzmY3Og4CN/OPcIdw4QjBL5p3hJUTJp2Mhd3+ZTliRrQtOFjFWgYSgY
UyugBiGy6+PSO2q+pJzHqnKP7CikhwKqYVwXtOTa224q820b5wuKGELozoA838Mk
7APNa0X9ucl9JMG4mBfuao4zxg7GoTncWJ/0GFo8VyvBWmz50ycGQ89xvbLDHxbb
LX80zxmWOSTWx0I76gKO7ysH/Z5Vgg+BHnzjhNnBPkEHuAhJe0QD2nppOf9W2EDx
7v0A+4Ne+QUnp2FV31qOQ+YQiI9+IEf8FHuL0MEmA7SyqrkTT8G0YoJvX2j4AluE
QnQh+D26jqrvTTSGlfinV7yU4ECx6jWxwCQO54jmwxH9WYDX4iQHvFehO4kaw2XX
c9enIQ/IKbryp3oKQ7YUBTepH/rgI7G9Zy+QqNcNcjyQm/sGnA1UvNebt5Exg5lW
HO14DJg5ZwI0qWM2JXUJWBkcvdinR0ipK40STjKYyvq3VFV2paAOGFxKMdskF0uX
jG1LxubNbRwHAKj7IIWplPL1FzhRuwktuF4pIAAzFu9NeYIVMLWFZHt80T2wWloM
5BX8ex4+l/CBb1K3H8kFtm8njxdYAmM94kEvdZel3CuetXcKBJLlu3OPB7rMkctX
mVDXoTafVxel0fMJCXWfBR9PTMWohYDAba0uwnLVpsJ4j3LQQ9roGV/Fht1eD2FW
IcJ7t9tpVhp9wIZknE6lNUnbuSccawvwukWSI0KfUCuv0zumeFGH8RWn3FT/DOUO
auKe0AnYxEqa57GAPypzU9VMwhGkTvvGVgM0WvFfop2GF8M+EwdmUYImcFQgEgbf
S5ePrwcLjVV89SQyNmZFvpbeLeI2UhRN2dNYXA+6+TkpXgG1v+Lb2Yi83cWm9uLW
oT/rr5oZbCoQTwPxGZjppnPa/UqHjx01WCG5hqjPw0+d4qRn+HTYZPLAquwqj43i
wW0/od6lmyY+IsZ6TtvLkGF8icVhg8bL+SjGtTtdTpDugKSS2AGuIAyD4yiFwh5n
RtdE619vQAgclCOwcxAeiCmpnPwp+yi54fsD7/eb1m8bJB19Up3XC1lSBDzcczjP
NEpGBuZeQrCMuzUWil9zexTPTTbOQQnC+j0x9bj2K7i4gW4hq4IwOOK9zGbiFnva
82im3FdoUTtkMMRQ599FdgrI0ml3YcFrCqoRl+BCLWEHgjkWL1iDyFuj3wmPsTZz
QIPJFl48QyzzuhGR0rmUMgSAsGB1mOnEwgPByg+OGMBp/geX6PSvazrbve9WTKmE
sGMTKFobVtauumf6mmv1cfrtlJneVMISjOEjnbaR02lPkwGD7xB3uvL6ORH1RoBS
CEhVu9MHirao5rRFnC/Kn/S2bweW18tg3q3kU7DucNIORZpy2DeXNjPg2wQXUA3q
EnGO5enulsBBheoFbTvnbAogKWi0K9d1Q+D5icXtpWw+Hkhr3J2a1K97wY7hZ2Ko
UrBHJdL9PmQRGvNKetdE3sAxJMA+F7JJi3O38cB/L3nnDdcyAQaTN8Vn5Svt2w1F
l7fQOFhItNUWI1NGQwryvYHAbBom1BjACsJsoWZ1cFn58y0hmvOSFfdiZ9x0eAWQ
UNpu6IH/09Hh0wFJz+rBERiHa9TZb6WhRgsK2CnnJQHeOmoL4il486BQTuGLtGdl
MuMj8ku682HxBlPbWGM5hiLHzAupNM6Ai67a5n/wpNX+lUur06sUJZ/OPUKvgehx
ZlB12ceeoCFDVcQCC9QWHZitmKQzMGtGjta2vQ0BS1JWXdg90I4jITbl2e5FZTSa
4y3OHRcgDanizuvKf+dniEbtMtrxvRxpACDGVawe1v2I9il1AEMgyY9ma81TlNCA
Pkq3MTUkL0VCpbxFYPWS+ceOC2DFP5VoXPK9LzhQAl+zSm6a/xxG5cCOg1bKKHju
1oVwMCp5huvXCRkGUWaRusZJC8KvOeYkCx4LH5YPUgdx+BABWfHWW8/NG2RjM7OW
ZXgkkMg0oYwe7G2tFT2hzb7+mXG/c7SyAdk/9IK5Nw44wwBvLo3RlfsK1LY6NOiz
HTajlE4lDFHWR/7M+dCGGIevZU9IvG97jjXv7zL4X7qUEoApAXN/oj/1sykfXabe
19Bt1WQHaJfHgUoA8OueWC7fWkzlecwjT8c3wEDNoSwXszb02X7ENcLI0qqp960j
wTT6YF9JJjCvTpdfUGHSNS6spNgwGuxVLGwWKFUpUsiDHRdZDolAWJBrzTBZEFSc
n5ORk437AiJgbusBX4AzxTrl2u04lH54If0dzmjMcKTvReGQDUGiytSV/Atj4OYr
opU/MBIIvONRKXzXj8FONNL29oraxAyXGnAzC7EmLChOEWlU5SNH2jo7KYW1EOkH
+Vso1tdiHYH3g13Gi7iC1Zqu7/xsut09xbSi0tk08KXY/jDaUmXfHaEa3EGFNH5/
mefPtYgsOXyF9LO40ZsHHBjGFqwf5e2ohl7+XLRiYIhM8jx/V7tn4nLcDKSlIpyS
QGidgp72ta3LTC//Lg/tH6Gwo8a3QfmgEhZ/28F0mm07aiQ+XU5YyL3x2OrGHgdC
BkmBEOuIV2alscfEQTeeR3t/z3sMoXlJcy/tsftLJzi5cSsGKiuWu+xuqJ4ICkRc
/vSBVth9LHllur+P10K1b/hl6+SazpYdHvEGkWS4JA7oVwkvNibK4waBiK1nulkh
6GUBtfvbcnxkN77/6aHnAh32TlgHHZw2wfCw2VVpEebetZiBGLGAOj8XIP3DYT6C
OtmeYAbNii1vY2QI56V51o7QNSXo4dACoMWH+UM4eRFMw3e6NOMnen41Ha0y9BC8
5U/iBXUqxX2AmfcYbAyrb6QZLSaUnze43rbhp6Lp4nZADKbeUh70kfS8vF0bnz1+
hUfTi4ht1z8js/O5Od1S+HIZQyd3MMB/7y9nwxIDahgW/J7/oL4u0637LQcFml//
9nlOlsJ8SE9JRXiuaUC5Ce3piGpjRrYt7Ar6MvMGMlPeSeNE4JZ1sTFXugFa99Rb
StYlYiYYP9/uBsyCdCiwNJox53lRN5LB6ttETPGoYSZ34/cOVH/JQ8r8/ML7F3QO
I/thyVu3Ar4DzDgHPCQ8NTONGKYc6FfNk0FWEUTE303S39tvmiUy9hUg/sI1z2fd
klKiz9aUy3oior9/+IwhsrXIBM6ByqNhdhqLAsiXVgF18P/0NVIFB97TdRmuPoN8
0DNYc3Hp53GpdfgDrJrklmILv9S6tTgQVttu3ISdoo29QAZi7H6wnotm7beqQo8q
Rlzn2DDd4LGQVYh7wj+rZjaGHk/IDuF/EzcNMPwVbzu+se8Jnq2sTXM9Rvrg8Mi4
nPGItnaqLyYWSgvx3slGhxVSHQWGINdlPxpAD6RfAz+Owb8V3wqK8lBf85nUcRvt
dr8V9tuZTZckaOjHVU69F2cwYLt6MqOR5L/tOgleGV9BRpMbDKKCBGYi/hl0Nqft
n4nJq06o04wNdvQvRJ+CJ/ZpjIYglqx2NRBniF05jlJd9yzObsKNOdZ1fwAX9gtt
PN3SNak6pb2UXcgPnQu+ZMcpCIgnVBxRZn3Yv95JrstzQSJndZYa6oegrURD+GUC
s00RaxbVxNcoOWXuzRl6TiS51SPGTu4yj+xXtV3OUtfg269ek/sV0jnD/j8eRxIE
CC3HCNPLhqfhSnRCtbRn0LpvHyf3FdSjZNfjYutf+f0/fVabpscoYNxQzUIhg80K
l+EX8sNQM5KX2HYXYTuWbkXZUxsSrfBvtpnHyNvTLyasqvfW5q3kBZMDC7zHxsJy
3K0bSIES3R6cyBi1PuKM8gCiR8qU8MvHpHxNtr5gwZpyuu2++68y7NaFtn7UEvIA
pYW8QJcizFjjdE+iIHQZg1SyHBxPPPZ9187KarGBJeAotur0aSwZdhAGRLTeD7gg
bkXKUNnCb7eaRImH610fWDVGGuQvYNT75Zx5AZYfl6S1fSA+lYwiAdlTyVm0Me4o
Aiu1eEh4KOOP/qd7mlN0kPA6BGNlTUk0qT449tGINqjwxsiinYvu6CSsMwxQdRaq
ljH1fre96LGUyVGirWgNtNIeIdjIaqP4np/E7TCNnfWEXbcHZgfoHhZLNz35U+fI
x0uRK1sp1dTAcCM3nMPS/k6wcFofPIo6Lal2vZ6+gIEWXcEUpaWB07KT4Y0RAK0t
ZbdG9evCGtLX8Ilo+NRSi16zxO1o2+IlANJi92ofDSw1nnFwphUh73NYh1Q+U1Z0
UCWI06JMfs31IRoy906KI3HHIZ5qMO1ogXcgBGBgx5br0Cm3Vb/0gYOp/6vVcnGz
cGURTjcNi+ymx3f/aai72jplUMUuojNqVbdaWu+HiJSyBOv7L2KIVPX/fsS1/nf7
9ymW700FTUE0gTlSIoKyiS5k5pex7ihsG63KbhIVhrsUl1jcmAwU0pRmO/j7CoqD
XG6d7ieDL6RUPZDMypK5wwilIJsKEvtyxiD9rMhnhz0CpPaoUN7l1Xqy+572qWtg
YZk2DnSKRFC3bcp5Morwer4HhHfa7Dm5o4UAOt9jzUfNZi4Mcdia/heismm7JWAV
dRV6/TM7MQ23draK6og/JexB5/+jCtrKqketzDqcgST/lcYnSew2gjaaoBppKXag
KjA5lyeBdMO5tp+hZ9uzjwlPDQX2li2AVG280foJ71+EaqHA5azQ7q1VHfoiKwSt
5CyvRGuUw8PHLqIblUk66dEH5DTHjS+4EOxayjDDFii6Yyl1kZKClcIcR4uVJBk4
/Q9EyCB/6ZhvJRBJ3oB6mybI+w4JvJcvInl4LpgjjVklceF1LUpdtGmvrvqUAmdR
Iv7iqAlRugbXjVpk9/iMmjdTg9/zhUCqLRnK1l0QpOkFq3oC8uWRt+yLiPr82Tcx
6atihiawSqAmC1vfCvaMQICV+/uJVgE/NMUQe342c8UDbk9A8HEGL8Bi+c7cZcOX
p/OPJRZlPIA7G1g2ElOWEtXdAOvsZjtuIOTm53OYS24ESTGou6Xqp/0wgRmcdke7
0jjUb4Oa2kcy8o/MAtTwJs6AfTzB4rTt+jM1pSdT6OptCd3LO+yDHwBFsUfBrtkQ
zODpB16L8s2F5nLh/WkgnIMEuw4TjVHjKrim13CiJD3Uar1zayDsjZfaHEQsy7hx
O0m8c2g+I+kxDZYmcddyexDHUOhRoV2SfgPdkOjrjPqDrjudMXK6FRb2rVS2ZZco
Mn7oT1DMLRdx+1b4qAEh4fY2Qg2BuioqcanIJglFFtpqgvlUYiNuccu82zzbIRtZ
Wtswrg2NaHphKQ2an0gmjkwKcuIaxwUXStHQjCROlIcQCgPgJt3MYgiNcc+lGBin
7brv5MIIAhatIOMmgOqhc3w4IEwVndqyNl5d02hoE0EyVH6hbzn0c8Po/pf49X9s
K2H7gi1OlPLcUC2w6sh76cObr8GI/YTcKnyHW+hH+1q3Yy7cvbS/BUkykue/RdKn
1DZNzruenESIG6xNrke31o4cKYdgdmp+GtuoWSbzXNIV9nhz1kkVFMT7mVJkh6YU
pZuq/X0ra+YCdm9FcHOpR9FtKODFABinnODb2bMwQwP7pyJSIhQxZ0J9M5kIVpg5
WXp6BigIEgN8zH5RywzEFFZ8cEqvcCDfgBVdzghv52hpJ8N8Eft7iR+ssJfGb3hu
ptAN8BzFtOkXg7YIzoUqDO597gE/BIpwDLF0bnc8IznhfiffMwuF8AzSwmXtzyRU
jyOfT49GdwwJ83AowuspxL2e1nTSu1CYn75MNKk8tbI/g+6oZh1SYi2pHJXeCjWF
FBJ8ST1wXJLy8bfhv228CK8XOM4cK5jPE9scGVOWmikSkAesIffJlEAHuzo3aZXQ
rnL9k12XxtGmZpdOKP4HnHXxpzdEnLRnp8AO7NV95gAc/GhJ8Ns24HKJCXkNtxSb
bm4ncMSj5QK4KJCkrmpjvoLnzlisKIVsQ8RCVQXl6AA102jmfKe68orf2lwYFl3T
HkDb494wuKqhiJBScDZ1WhNTS6UA1ujSUAFWeMaUKb7+RUDnkB+P1UE4uKi1VKaG
rly1GzN6Pf5H1INa7q3IlRTwSsrat8NMmfQuw73yZxoiDpnXJT8e1aMV/SmDw02s
p19JWBD/z/oPCo09mazDYIaHovTLg0NvbQ+zvbc7/L4iBD9xixjCyhyIXo5jOUlm
mD66mhTbIcTES9fJ82AHANvEDf4TD5T08U7Ajmh01jnxXRTVqc7GHFEIQOsm/AD3
X16O5vHBzOZovBkC448cz1X84ON2kyGo3kOCZ8y2UuxJtVFDsmkIEm4X5Z26quNE
4KURMAtqPTs/+0ZdVcbvbL5rCdKHU6+/h1JUPSHM35AIvZ3Vq6ZnkRJaMeW9f//A
1Vd0dKK/dLrXs/McDjpUvBBBHiCbQI1jrPqdjggFXLWmMU4e3sOZYN0m9VM30+lj
uS2U90dxmh5VYLoCh7Dk9DfvNMMnJ6FguS7zplt5vHVQ8xemutblG4x9WKMVywOO
70dwg7OqQ3sLnVqM+B4nKRphMIjQlcWEfydOMZK2ln5fNL+5V8ia3AYhKfUKv20U
knC7ZXZLVy6oL3UWLeA4rwsj8Gm/1oQGxJEy/LoD2DbKOhtHBGopaWg5SwWoQLqM
j5q7zFg5xMnmkRtU3H6GN9jWZG9qxSWz2/5hFXxaLlS/QJZ/Al5nWeccBSXRVhAl
lS3BH9bmM3waDE69Y50QXbjY64/D5mObSQv+wrN3VxbBoaXLMHfz0AWuAi5YX7n0
Eqm6pjuA+GaqP+8+59A0L/3ANSdCOSLCTTvLCU4VI1vFwGFkvwfUg6bwGqpp22y4
p66KA0GS7OQ9qVvzqIEWJCMXsNvNo5kWIUFjyaOX6GBNTRsY73W+cur1WDGbJtRd
HL6Aul83siJjsAn40AWKkVbzTXv4hM3CPyN/RglWMNox3I26ruaOE+rU2KyMUvNJ
y9oFv6NRXaSIK1N/V6rt/smMziPsVccSYc9U4YbGxHDZgqERhMa9hvkDiaE1S9Vg
W4Z44RlKkV33152vHFREybGWWhWqQB3vLUeDlS8/BcXu520VH9Ur1QgAREmV2BWx
bZxbyVBHL8U1COK8m6wwAhcG1glkoeGSQGy6zPwV6F41QCkJ2uqDPHZqYraCyZAC
ORfJUZjVIa5YiGOWwyzCR2MnijG9OkpP9Qm9Y//dUrpMxlXmnGyHwKqmwwCfq5cC
E0KHmU6Mcimyq3jN3hiZBch8hTRY2mIcGqmu1Bp8/yjdCW9xscsiN7QZx5kzdPhz
UuxUBdIS3ld4u3npmVnzb1h28uHbPmONmp3XGqsbdHqM5/M8O4NuOg01t1QmeXxA
poy7+vTb6YfqZrcHFfX6+31f5gIjTatuuznM6rs/p/pk8ji/Ra7KrobeJCnvhs9j
eaSJjRkOye+ygggyuhJV1WkSl8Jyzx7S3IE5wEF5dtyzGEFv5zmglvneY1xOLW1D
HRFvib+pV4upaBh84++lSpY+k29xXo8vAMfP9oqnuR1cl/dmrMnDuAWrAnnuGo1R
n1teIr2QXnNqTwiYfy4EtMqZ2ypqbd/MkyykRxlQSFmVVhChuLHN9Gf0CumkfCUs
uvTiha43Bxsk6tRrztUmvdFlx6ZwzAwSxOCkwFgaT62snDAAaUhRakm80c4mTXeW
asDy5CCGnPqL6u0CDbcu/T2jHrNsVp6nnd7TK8Zaox9dyxFcp4YTuvZ094OWQxId
3kAmVs8/6d+OXa8r+Lou4vPUqNpJDQ5cVqwoQyYmnMSwTDxYjKCXNu7EGf0VNOGj
gaCUyCr+I2xmLvSClwsWXWKlK6vD1pKedSE9y7EHZTLcRYqMlkkeSW2Ra9VTOQC7
6oy2T0AGlwpQ6qhEgXBn31cT+vsAyI/NaPJt0X2FLUCC8c9DGunzpki9k7DnIbfc
ot+VEshPSm8YJD0z3cmGJVbD0bXb43AaxzgwqFZJeE2wjg13zZL6AGefGU4dLA5n
JhMzEgymuM+WB0iTi771Y5usgjxbZsBj4whKsTOrFlAckU9G3nIzlae+A4qqC5+Z
azzeEIMgCzef63nykXPjOamOg8CNGF9z5EfdpmqE+r/tuF7AHcyy4/IsuJHvcTOQ
9xYpBRT7lfuIzoiUd44tqxw0DIJYE/r4WOZD+6ckAxgvlh0IguPNX13VtmU2bH5d
lPUockviRi+9ni52JxfTgpcu5pi5GxJ6yOtENyZPJrE/4yront5krBXEbItuB7sM
knsFgikRL/kM9Loq1ZFjR23MLtBReA5saPUokqf2fD1pZG/bmt9/dbD7yXJEBtoK
QZqVWYcltnFQbt0D4K5UCparJHV4/9FSYcYXRoRT8/Rb8VzPBjk2SJEul/bXDIkT
br5O3c4wh88d5EUHSeruTQfFIR9nLF7iOowfGh4bFnoyYCkLUve2M+VYl7byYxkZ
3qU0cAml5wucmeWc+w9LJc90HVB5dHU4cZniIiNI3Xg/adhQZ2VNlsxM7/j1NJsu
S0yoL6fh1sEBY12F8G97hZC9vcHOatDafEdM9oRacqUlv7ArOldoolAtQodMgcAp
qXL5pL4NROLo9IWeJFrw1zxyDdlSelHa0ayqbezgFwIJE97cadloTPrK4nHCUauG
U9jc6lDyZnzWmKe2jji4pNL3yFHsATeG7HadSqWwgbFUvRLYa2akfCgUYZbI2tHK
AxZO1sFjhbSgOaTgYoN1snH+thZ6Z1HCwPGNk1Fi7pnZU/M02+sWR8sTcny5z1F4
5ggglaDABfEuLUpV6XfHJq419hSOhxTQkq9E5+nsXUAIq8QaiU1RJnPH2eaq8QC4
QRF3h52BOiDyP3/GRQC34DQo+Gm4r5NR4raQPY+jBeubv/+5Zfsv+NyPSCyyxRSx
rlJkQEGmLP2bX+aGFVTUERFiregQTDclKclhBYKQ3fznX5X2zT2uOSZZ01SJx5F4
6aSE5w0zw7G6n8B6VB7KVo7KuZuCRkrBVAOOky3m56fP0fOnKKwjejokdKLjkXql
rZzGXcH7LE+RFYx3m5b9qenQTvZqD5KkSuMhRfoXuuh7lVnXwwEaEmzeSmkG8SdS
48PB+Ryl3WfEvxhT/ixvJtSRiv+tu5YQNUgMfMvvIs3TL3VL85dw5LR/DFvheK1N
Q3fsFmPP/1ULomR2GgovbdD2IOhuPTRqHB+XsTHEr1mMajoU54Wiow19o5OMY2sI
ibNMZwmYCv6sS6tOEP69Wvstu0D7VYSmTVDmWAE0U0q++tz7ATV1oUYwUyr56eDZ
MHH/aZKqeye1BhgTKtQ9hN9X/6rCS7lMXNbLrb0qkLjqVkCPfEWeLqau1k5IUqVz
AlT2VqPjIvd7Iid40PmqHZ2hhj9fVa1qmnLHRXgre5jKZ68fLNlBY0q/+v0L+c5k
xSTsOWPTZZUibRHuZE6pUqfbtJuWkd19nlbrXbZnTLJNL64nyJMPlgVmS0ypPm5w
CYA/p8tmNI0XVRhloE/HR3jb0os90dkKFK7qCYxpRs82mDb0Tb/xPlG/N7QTtsHY
b/14BRIsIwnd3q68ejxUYlys1oxqyGR+KVqSGNktlMTX1KdacWVaAR3RPWjLrpSf
CVyazlU2holWMcNB2NQJ8JtODnP2wFtm96HzXZmqoQQ3B0yVhp+VA5JKybv+SMCw
GK1YoJ/6IMObJa3idWA609fJAniMqjQj4BZ0Hj50R+FzysGz1IA7DpwSI1XEJ+7P
uEx0b+6qlRAngF9BzDO/4mRGZDW9KEiJoQk1tHZbKL/75l2vej7laILT0E/bWmAE
9qkgk/0TMEWVGkBTPapvzC2TyyhGiFu9/E3lFMLKs+RMeCeUsLdDn2Z/POfhDlnQ
+s35RAFOa1rXZPArWdp0bTS/QBd2hEUO/rlLx3gsFxHiZK8hzo6pustFsd6T42Ap
60ztECrIrM8fPEOiwc/IbaV6WLQ+xHKYXwThcjG2YpBetF4C5oZ7J8u3tdGBtQ8N
1Xz3noHxSPCD8yNa8fbkYVkGnUgA8uz1R+vkzR2hZIuzOKJWxDsCf0hQ/RCFsXSK
SJQFwKSpiMzWtOKV65xxqifCZRdX4GkAu/L6iiy8+67DJxUmFWVO8ED1nd0kSs3V
EGblqjQQu9otwt1NflpwmOjnNaZsCIlqhDahNnIliN2VXW3HqPxucFCIejLKcP+m
3h0z/tIhLgQGR6DEzFTCo0QNxxEKV+2R+gTsYjQ2cW9CcY+N1B6N06+ElLnmb7JQ
wyF6BIKknmSFH5k6+oUYuCkxEtEaqrY9DxBnyo9Tb0j8fsp8KmB23ofv7ZUxUXNp
r3XNS+yQt6KddrOwzwqPYdRvnKqhlvnFlZ+VUZOmYoXKqUwiBngJ77LC6razVboI
3kJAsjviXZGOA975GsvbSF+dLdQXXUWBE6NEsBAcr9tr29jUpi0FBITHftOy4tET
Yuv2SBzV/3SpFc6KZhWPH3iY/6SoGt/YfKp5fX+RiVT8+RVVWbLKNa9PHr4g45ol
UglvNSKa/5GCHvNJ6AEq89cssr1OZ0J9UzpRLpz1Pf6PSWlR5ykn38WQgkusshmP
dLbSeEWHsFMBGz/qGDShchLg5282f2yp376tE3hJse47djDnbzePJ+J8ZjkeGncI
089vjwRQ5zj+F7CJr/i3Wv1ZloMbLmtUrTyfvso88Epi4xOMvfYegIqRQ7rrDu0u
ogJLUYvjUeABuKSjvsxfMUOs7JaYHDRAONz7sEDGjH1G/hAs33vxmKnVGdd5nqZM
eMP7hWSu3j1sCBUwsj0SwKJKNKCmQfEjWiMt7HuvTJMDGr9Wv+dxZiex1hN81eyx
kXVkgVfsLq5smEPhDs1hHEN7jia0Jge3TO8hDS0ABrEMEsVlGZvWYdM0EShqZ/ZY
ixgggPxxnQeh+9Tp8ib/xKJWU6Du5dqEEULJ2xzJVi2hrcmp/U8O1Hhi4y+F467i
ClXfYL2rp8gvkmgSLY8b+p6fr7Es2CpFdtF+56Tlt9tHnO/CIiN6HmBDq+A8i4rU
l5M3T6w++M/sOj3uyajLoeHfBCrJSIvOqc1bIQav76SGQs2qSP4zd3081LwqgFbO
MJiXtf+N9zDyOI4WPxi26kz2Ht2EH0fCk5QNFBSrh1uA7F5CEXdrhw9MZcD1vkHw
ak2+vCq2Ks3oYrM7PMBKtge0Yo/6KzUu+UA/vwc/J6VA3yv4J12cAtPFwLFuax5t
6JpyayxaNDuoVubUJ1zPvv+DtpRKll7OEQPGl7BWNbIcXsquCCRvKyiyUTeyOF+1
9lmBpFVpPKPZvbFDvfwFUcBnwy6JgJamibBBj3CCUidawsF8N8WdbVSAe7AiMoAg
AgMMjJhcDA5+SCpQ6mTPjIxNHGA7Z2uXoF3YFKyRGlOXL6VHDE2xYLeuC4KIiohF
eIHiEbeIfg0pG2yS3Zy4gEUeoQ48lzkeNlC3blvDMRyJsa6opoZ+si3enp8nND2Q
22v/Vm7d2jAhuNiIIQixDa0Unm81h58B7qR8BCw7uoCH51EDFXm+X7tzdEwyXXFl
CWg29biG9aKVp8EYtXzghCyTkJnqJNunJwpIwFaneRqKPtZKVWLQbWt6nuWoyIt3
hyyLAc3W1z4pTwTJ7xMihOgKWMzBc76SaMrd/W/MZQlRKWd0xJ4eYoHq6I3Eo85G
+331BpnZv1fnWrqhM65C333bmfv2Z6IBg+WkWYcqSugaxUG1pce6xJ7/YNlgAZ3W
rG4pyRTDFJzAnV7FCKqc0libk+iT9EdZ7p4/lBj0z43P7/4xJS3dxLoJRd4exs1s
TIJ5CaNElDFmpb0eMIIuhNW0zSUf32vSyKoq8m39niXrG5ioJWxGye3dwUDSV476
XJyg/Jl+2O3lHyfU51/fFIq+sTMYIinroki9z32twSznQOgjj5lLLyJaTYmjsVpZ
yiK/1agfZbOKPZg0tGAMJwXMhZ/SUDagP+DGo2Uk7UhNSoQoECuu9Hko3FYhurLU
ckKAzvKpen/j2FoHnty/J/hJ9JmfJd+xMG0QmxMbyBi8KeEyQiPR4TLXte7ldeRU
2YP2NEtDsbAaLB1ppSADYOg9dHwDVWeaiadm5enX5pWQyVv0SBhyFVtIy3+YgEkH
0gxClCd2zumj3Adfq31KDzr5OyRIjjX7sOys09EuEq9mjcNhj/0NaSGxns0QzQ2P
U1iLbm85ZN+fWBjOPSjhDaxwAcGNsWMNegfTeBUgQASsQz7dimh6MthuD13fuGKB
DoK09JNe0LQ52WPFVDGpXZXqeObL+wItgHHdXY4mxJL7eYJDF6voWDl0YkR6pEAq
51hnbtAV09sgXYfKF7nZ1F80eN5+vOsAYJMKnoHLJNzW8Tl3yg4sH9f926ArYGq7
WsZWoe2nnlfysdYawde10EyDg0+oJU0qE9tj1VrDJ4grxaAlDCsL/AOaZkgXktEP
uQElJ6ns9acRz5TasgLIBo2BEN1rP4jej3COsHY5oRMqb0i1uXPamNLB5rTyiOCp
bu2XsVZZ4YHawSy8HD3zJLfB/VhLFFI2Meiwsbj9dkEV6em5ifUGsGmuQb/UaGIm
KCKJe7bCGVlOywFmfde6yHWMYDgucH+W+HNKgqxWul2q8ucUqVXeb6tdW6GxUf30
Xz0v6Xr5m8ElqOuwVkXt4umWa7hpW4g0itF+RtIi82D5DUYn2Z9o+4VESudf1rBK
NDdW/dhIczTLpIxCfdOMRFIkir+aNXnYbCtQE5rGJzl+j/N1PTC9+Hg5qWLaVzQ4
HpKxcL77g+VewJOLUM/K5gADkYEOeLGqNSpBAjRtG/jlsqmIqvRxi2CSQ6FLgeh1
Vn8CdYQNVYJACEFSYAyfOat4SMShAQgrwi7lTGnRTNlIcaxuCTByRxirpXb/HEeq
Sw9gRzckJlJr9OKLZHQ7/HfXyzv+8PNN9eMC0/LSf0z63VBK7YJwWkxF5t8LHrtk
VPu/OdSybxwbDQ3vE7p8sc0Dvn7CwEy9VFejhkeXtLB4367dj2NBSzlKYp9g9O2I
eKeKF/2DoqPVE2jikB1tMeNCXzy+X2K13YC4+hcoOOJVhFYQK5oQEGccn5CEoiKE
xLAqyPRAWJJahkybHcejoYV32A/aQY26XZHWMCjd0Y1M4I9bjeKjEJkIuha8rQPN
fStTTz2Rn/f6F7MyJWlMD+ht3QeiLeFRCGqdOwv5L3V0KaFwwdMg4aKamjdNNTtF
4htK2OXj19Q09iWLsUm3bAcGTqvyfUYCsSsOin2VIJ4lVV+UsN+UPETEL1oIW2vY
K+UVPPqf3pDwqSlNj7PPWeBYfb8mmpNXl60Q4hJdGG7vaub4U1TGJl/WViYTYPcq
DLtIyX8VAk1lpMAc3PI390ZWkNlwS/J4bq3/9lwdaP7osXJTJbQO97jkil4o5pfH
9Whk6mQfPGcBhztK9IaxV/dUopTfAOn6MoQLZ+6dyuF05yXEMQyGE4nzQNucT/G3
qULA00ME5Fyfo2Sq0Awk+hjo9D2o3LUc+Ch7OVw/mWTuWO2AuajA7Az1ad3tbnsT
RtFhM+3mX3OkmSCEHviELyccY1oTMtTIfkEZRfAnM3yJR+pzRcqdOZXiFOlGWq2k
rPT2bBtNxJVMwqNRV/0/WRnRXLoLOdQR+kT4Aztx7EulYQ27gM3aS+1CK6uLONKZ
vSuqV1bNs87zEJcEjqMmZcsTFq53fY/nagAjf7jcibssZ61EmG2DCNMw6hxb5bCO
8HILKA8CFSTmwaoiv80DP3J3hTxMGAuk7JTLdvmnJg5Oueg+t/PVnMGyIZqaUNOR
YB0kFaKBvad5FsUugQ7SNXZkfQkI3LyTjpwOL58bXtgzlFNF3FRcqpgAxIdDhK9s
gGqCJyRum5LIuZ9ZevJ/42rDFm3WoNvznIwyCduP7zujwu6BwHmqKpaHrdPlvf6c
TcohGYOvEuDJFBHl6x/TCjFU5ehIj1YKmJcckkifUTq+8VxWU1oM18kCUCp3H+dK
JU9aFzBMgEpn3jHxIfRCnPtfNNc3+oDsh/8bG+NRvpl0AWHK/05vB9PYS5rR/xqK
CGf1bPSaKviO4i8Y3pqvmka6Us6E5eIpYf8uxB9k9pYz9l296KSwnuLJJWHLZPgY
oJFZb4vyXTSkDl58cMaUVtHwUBCxmd6OEPcbroJhy3F/q4NYwuwdvcQkPJaD0gUn
xw1FrPefoh+QMk50JbXEUNU1GnFbTswpNZaEsDJEh8M0tSmY2nRo9vgl4JK3cWJ/
uAZ68KRAeMgbla4yLuXc0aXAdgYjOKtQr3ryTSjyExy7FjJZWW7V05ZtyplOX4k0
dBsSIuowQELFatMIme9Xb4w+uuRDuhzg/b4t1uDG3EkaJyVv0+KzTjUK8CgCT+cL
iJLKjaWghXNSNmrBnl/SFOEUElcQ2mN8bymFficU2WJosokPQmZ2JwpRcez1+JDC
Zcyz0TVYKZwmREIjWgZtrXe8y78TotWyy2DY3Vpvt/z6AWXZaIN1y9i7Y2iSmT3j
bG9VT3OehmyRKQnMIC7slgmwiZqslIFWD7Hc4XZ6FJhVVRnkbLdeF7EIZrX07qkG
mHXPjXdjb2bhzNk5irFV2EoOqwfN+w9afpnxW5jfv2LljoBNo0hvjI6bsi2x339i
WGORVS8Bcq5TqryYDft5XmDIFRakV8IAnwlJzOs22uJt5zOqEEDh2IvZUwlD2JyT
ayg4i0gZFrWVHViTjO4BwmuwBNDTE3BAujzoHw1NE2PA4+7APB/IWpYA3nO/aNF9
uQsFqfpF23PY4UWDwQWLByrbIiV6+fje980Fu/U4gDllCZs/0zcisiumEI1syhgc
znFkjGGqCtKOs/WP4OuJAkbA4rzKXgARGn2C7iT5moeb7g0yd9tNu2FdmXh7CAsT
lBsQNMmXZA6NjRkXEzhJReyLZGz2B3e3leHV8Whs35aYkcFuCoxOiMjep+zo3SFR
fayCPGeRIqR5e9AtDhuykyCHGQbymu/lFRxlTUOWywFAxLXocJrRNPKrJiT76+Km
xssnDqdRkAGETUxFYox8gbKe2UWI5QYkDOPx/knUmuAV5Dc1nsrqZ7d9Fj4B4qo1
PmrZqdUYlsW1e0ZelkUDcqOGVVmxpBLyEnmHMp16W6Orneu1zMshok6RUjYatPYe
iSQPZZMoJIL87+Lklhys6HD+fB6zLVGcDIsFl3VmHa9jd4Q+9qGCWAHypIqJHedp
Dg9YuKjrGZvY2gJ0VZ3B/y7Hac+yNK0KmAnk3zepsZMJsEldhF+fsBZ3RxktUE4h
EXiFFHh2WD9fTC5ow7RRm0JHPdQaDfJWQIU8ygi5wtwEEbM6+kNHC0IowpaSScBE
lpcSbA/O2SQtdvK1/9HCeQ4JVlbAny+ZN8TuMERr18y1/kDN/H9a2emHVwjqUnGn
nCIm+edIK9JiA22l3DCfNJWM98xsEiMTnU6Dat2pyzmosTa6MvKeYYazEC2wKqbP
yLhbWMZwrEGFx3tHy+D7Uai9sVIY6JMhZqdQCrHlnDOWiVmEM5+wUjgKlafTdDx9
OlFrwAPmFqNsUFfmaGEbShq2ceU1sBfcvZOSzhhACGjDlSgrM4luSda29o2UAPx9
R/jv9bbTVDfDlvu9FJWTD3FDfFhXpcwg6GaMbiwdJJ06UrDiNZQm7uTjGFbO0Ip9
9ZbdNMRQklxMTRzAUz22i/cwk/Yh+hgRmuL80G/oQv4eF/uHD7UTkAWCx8nJUM1+
sY2+ra2a1DbGmjo3+wBJLGkltU6a3OjkwZ8N76k6pyaeCCb7RmbKPTMpDKGku5RV
c+jcM/8BxWTP70iN1Zvvuayq+wMSrrPhwehM6h7sg5aZCIRnS1lLd/1wuJMnYi4w
ipt8KUr4tMlPhj66fKUKOy7QUtGXsK1Ov1aCevqogHaKF+n2QLaOYImoiq47ywR1
w7Cn3zwxNBpETT1lS9HM+zPJideb57BFCDDadLne6KzfQ6RrE6kHv+0ov78bZMZX
gtD/4oVCKi8+/n1Y6bDGTUqGl6JvbymZlgLWmxH9bR9I2FhkTdCudJ1yPrnKpwNO
2Nhd3rfCM5ETOhW/SeiD6xLCT433hHhU0so5hnAhqCwb3qih6DRb6FhEy3USaQYf
Xch4Y/JJtT7YxVuA5n3m6YsUo9PW4s1B2nEwnD7j7WsMF57eVUIC/o5PKqibxeSv
gSa61k/FOgxi5V1fsg+PoieTIZZi0HYHfg2FqsFrgrwm1ue3SNZ0W3GY/cS5y/dc
oGmbyDKvrUl9Sxv9TReIa3qcCxGQlhZukptzWh8P6b++uAG+L2gCNcLFKz/oIJ/f
3eDIPh0OOoma2A9R9A12RcjgUWwRxmCQSG7beztp3RJf0g0KVDpgmAtDLovC5nKR
WBjUN38cx+A12B9ukM4ZCq+W6NIMbr5bl00NjSrwnfcGi4v9Etwf2jUlQjxYeeK8
dXnQog0RHwXD28YRojTwWuide3EFpl0DqLAfbUu8oI5PGYmjD2u4oUjLFU6ZQk1j
zOU+dTITnK+956ayJ+ohjNtuaFVCQipuoVm73d6rIP6LvBNUsiCvE5KUgnP7DbQn
MCJMUzHVFBKmubLDgyY+hPk6hMiKFwkYQp8v9MDc5l1Bgu9bQRM2umeaZHkqHQxJ
hhDsIUtJPKOJ+WdZyIe/UT/EHGNyIYa3OqO4wnJTVyiui6Yt99IITkUgRHPQT/aN
lTmxUvyptpm/g8Swa0vw9rvEljdx04v5DwY5dDkCPF+zBGK464GXTUZy5OMyDoeT
5uYEd9+B0lYoExQkrBnJPR6slaFlbmZYMp49abCqtzCnt3nS3qNU3hTwSkqj9L3A
8j96vXa6n3O4gfaKGPKVz2Wxf7CU3vXqv2iwoyQ/AwcL6/YxalL+F4rM5nouvyqP
X4KRjinmIuJ7fmAAiTcdMCQQmQQmPxj05sv6soUPeUqS1BZxIq9Fr8ROuSE3XDBP
gcfoid0SEi2ce21X+/mb/uq7ULrbWSSiBtDiNpbiaUFeGVKD4PDx2DIq6BwT50FC
/u5/FM3EU0+szS5Ak47haowcH3DD436rsgYr+z3fq0r+zi5BZ95VZK1TI6r9oyZy
S4dDuRhPU4ori7+HcGp5xsSmbqW8VzfrqnG+jz1kBCvKMbWhI+HqaVKNQNs0DtYY
+n6mgzat9jYYJRzqyw0tNNq2CX8ZwGYKu5wNHNMhH1KLgSGE0rE2f+3fp4ZULYgd
00+Qpx8LaXHDECwsMcF6s+5KAp48eYFMKQCOiadsQiAjlc8QDFkQGr50b22gE7nE
MoXLIluCgv8QwY8s9tpQAPSzmb1Aj47u+vkufFhGvcvgiU6GMk9tkeNlGlc/KTd2
KMk4m5z1jhYmE/BQWAeT2CqpJ0CcndZ+zQfUAiNUP6FDHAe59veo/YUZDa2/La+Y
i66jyaBdR+0jDa2itl9/gXFTxXH/hZZ+9SfepWJ+Esq5Z4DPDjgv3xwQQguOyAEp
EDQVSCS7yGec2OhZi2hwb17BFvh6GDWLMRhsqOrfnyebe44OvVsbU/nFjcoTjxTe
RL/Ub2biwBKWBF5dbrO7HdWIzXMZM2cEoGqtVkptb6eKC7ajoAxc4viFJoYOkOqn
XXkLhXXMr0gklMX2tYS28VtDGu2vJ5+a4YtbGO1/M/kIfOMAZtES4PhQHSN1jfAO
Ulyl4jmsA+up+wDEO9nWRB98NPvS1U0DMUbQYM2fq9cG2KrqMlGTlkq8pHGo4yn2
r6R2RumlUOW9gdC2YVsfR+62KNsq7i54Mfud59YjBTVw7vVVSjzsAPicz75AqRNJ
PLaO+AKjH/DVDnAlQRi9IFXBY2DQ+Q5age4BIbcJf80vPkqYnfzOUmqRO8Dk1YVR
TwUDLBYOWZ18+J1ZsSyVgrvZ9pZ+P1pjLeVn/ilusUh7wxLcnMHzG7MT74BhppFH
5O+qA6FlrzECNjNowe7Hz4MRLNa0NO2qB9hUynF8lqxsPA4LQyi/cSJKbYxCu2BF
IA05CRafIjTJQq9bKV6i4d11sbw23QlEgDgMGYfKMPXvtzKh9WuxLGrH3Rsi21U9
A2jPajnm3YIAHVUVQCZjtLIRjMscc2IeIOb7raZdS2j31x3DMPDEw7uzOoZG04bs
2KaCbU5Jp3PGJFY50husoicgHJrfEwa0ELp/nhj6cQBCoK45chwgtrR18Mdy1yWn
dS39+b1/PnIejyUdUAzUxK1BmfAicz3Ay3OL4RDNxB59lXW1CgVdY6nwOJPoGOag
8i8HkfzcFjPR9SDQuUjjMNTL0C33YNlXRLBE4JsBoA5tRYULhtxf2iSuHtDDg8af
UxGFjdlsWy667go3ularFfxV1bIlPqZ6OPipXinD54FiBDfcMVUYUPCY9PvtTNJi
bD/gjP3IOSBTxZ0r9CsYjvzObV122xvyi42e9sRlcCBQ71PM5RlSCXkSqgyerRD1
OaYof0j86o6dWjfNP+Se0M6UEkAhC2n9ghFeZR/joT3KRd1RH9turfF+QPrqwdTS
vD8MoACoVd16hEHKpV1sySh0rKMuaaBQxBsfc2DwLEogFyHtfrkgHbqySzFBhyT/
IFIFEC+z4zequPg4wNAhPs9lIBN+n/IOLCSexJv/eUybnoYsl5rsmdhzmQcU1ZrC
WVxeIAbU7jrEiM9J4XRnGmcIk1xCgTm781KjVWHqEEL0Pt9jKYS/ZQ4UB0GB1eA4
Ml8zEnKusPACFY7oDyfBeMjXGFYqw9gi27GX09yrJ6zNkzrofeC84KJ/N07AQ+oD
FZSKHlv+9MzlO3vv9Wd5hS2HrQiFW78S0QpYxSr59uzEF1XnJ5Uqva6W5o/1h3UU
uXk5XF4ccRcG/FWeqE64QkpU5D/x9pN34dxKf6crZ6D5EtGYjfa1EMqsxZ4KnY5i
HG7kZR6+tr3bPfhHm3SNl0Zx0zsGct1QveMOJ7aYEMEXzZqadjAzdp9g5jILJdWR
VPkOc7J5yfersWVelelpPaPxiu747hej770QCc1EwZkIxwnE30VpKCUJH0w2L/vM
qaC7uiN6J33jg4WsFWtqo0Z+EEv+do6MMYpVo3PQx4hx3rzwEPlsbCdNpMFrbFBD
wn1mzchZtWJrqYYeJa/MabFxp/kGsXhFGyu7BO74Fvvn6CPO3wJNCD2RzZOXtOpA
pBAUTuPQTPPDU0EiaDukL0Q/6DT0TzFWX3AgK4/vYQunp2q8JeLX/jmAlIzI54QB
o+guoCIliH6ug7Q18nc/2A4pWuBS37looJxAxCPAUHyQpMUBWOpXi09MnJOQJj15
2A5BLOXugXzSfymFpIkfFVgkjR3gDcHrAJxBdGhvON+zl65dD/41HQcDLqwIKckQ
HEDI12rMQTr4Z9nL8mTXUKDt5gVNcc2HUj2EwAl6FP5nAbtGPdK9Qy3F2mdI5Hjq
EsKTkMln/DQ4XucD+Wh7zm6yshAH2LzazY1AdPiwGJ6j/mnLYWv67rg8rmR2Ixpg
hYP+TIK8YPAX2RIPP24WGgGCqOA/gO7VBAq0V0l9KhQBGzteipYzL043Kh05rH5w
/2FOGUihMFCyYr0gOotPjR65w5J2VYs/qlmk91hVfQOME3FyyMi9reRecn+k8T2l
oZzVTMR+kX5alEG1Oa7a+EpJ8jySi/Z7VFQCA4nunej5AgZmeuE9wc6uNpEyPWe/
ZB0vosKAKqsw30VpNGgM5v8AOLqT0PpydaZ1tvcJyvXpbk+b/z0KlTZT5AhkMJd5
ZT6ICesgBQaaYaNufuxd2RZJ/pXZLDBJ/zObXT6HBm/6GO4DnGikwDMw3KexR0KD
gR3+sxzwW/z8jFjgM3Ps6fej1/rVH043tdoTIEiZzLgRTMl5ljUqAK7snp7ihGTB
hnjOIk2Zs3jj4VjOprVu88mt8uaepUzFTRTWFaJ67uqV5WTNn0wd99DywAkVR1Ov
2o6dE4T2NUvD0V9a3uL3KDPPhatdqBp5v6EaYVbtdbeVIS915q0iAYU/oGsqINf7
0zGtvct7NSeNjHJWucfWBY+ZQ467Wsj0Ems4Lpjhrydi5WXuC+G46N4eWcYdT7ah
BgQns9xzNozcNJVs5RYeACHrCZVq91FnS0R+5/nzjM1QZVcVkNo5VTeCQdWIHIda
0UQtmHQjo3g+aXWEKywV9eaAEsXaox0DZiRkMQbh8gY8ZSrYCzUQ7KpH6BJsNOdY
Wijg/Ui8EqFHOS/8rAPShY/IkXwDE44Prfw/eO1z5XGdyQ+I8rgCdCUf3egrB/5M
y3bLh/FEOdimqc1rlk0+v4WvNx/KF2G1Ixv4vnb6nbg4qz88/P5LA1nZ8EZBCRSr
xRJ27ox+hA8HZHW2geugm+pAxUBT1jv86B5kT4L1vB3+RqitUPshUKaspLMfZDlB
vu8hhthH7UqmFroV1p1Rq01e6To6827rOhgm2oNmb/bJ0G96ryXAUv9cSDG7aUUS
IvJzSWUlAh1KsvtA+z8f4xH0kWXgzqiMV1X08S36lTtFsox8CNt1q+ccjlqlReYB
wsNtvGvZred8WtHKuCHsMPpowu/dS5ZS92XB8Gg2fswkmL+lrWofnuDaGG3tANyy
p0taIUwsX/Xo25TLI7PUDUMzO3JzGbeZ55SWcno8PcBg3s+iRtH7K3X4vgFjJi/z
jCrkm+pZrlQji7A0434/Z1M12dgCm4FkdIbk2ycpilAEiNpp5cTd4AhA2nNI8hpm
DlreP1MGo3AFE20r6oKdrYJwciFK+psooisTIS5+k3tXUeRlRwL46Cjq4lEq8qI8
5Yv/puEJv8FkXu1bJL+rPMDV3XyBSZeffrcSID0yR7qNI+YOflw4LxfEKsJ80Tns
M20ny4/MwQv1u8ZoMtOMetvYvzLXNsYjRRrW2pyDGEmPJwu0lUmyqHOyMQ/x8UoD
2qWwDP8rA0tnMo/ZiIFS3b3ib4RId7tJQyqY0yS1BRnaRcrUCSu+hJR4woF7dzax
EuO+6yYpmSGoksf2QVIeM5OyTQ4gfgF3lh89e+kSVBY/yawsV41/n+eFziovmKhF
Q58qDOayiBlqhLGRNKIMcUF8bzqkyOf6md4nKqFbb3PUdYajpjaAH19F7GuFhmSi
KMta1mYJAotgEWlY2rOmJQv9wG6W7XWYVEVJUaE7+YGwL9tNkIofg2cHPIK0yCmx
lDkCdlCcujR/eOlWZSyjUlvuPM0nSliy8MkKWTbHMgw6dkraeYYYWY0foA8Itxmz
DKUSw6o4u7hWi+AzRmKbQW9WnCM0dWo2tVs60Wh2PnrlCVKX8znt9tXprThDD2i3
e/BfbYT0VJpRs83NrWdu/oiOBTUe8FORfhVxRf7AiWvMwsWQJZfz+3h+dLb+657D
yUkHJlTsv41f4Ez8aQT9LPfi2TEfv2LpOnncwL8m9OizmfFi5DL2RhZ7dtl2bSc0
XYc1scc5Agn5BzKzS1o41ohVEFyD/63jNoSFE3ayk5o+R4iitKTWdQpq952gLiVC
KbgdL+PZaT5MtgdqvxTIguH8ZIC4mA40gVVJQSq2axLpiFKHafPeLTTfjKf2Xn48
a4uD7CoCBV9MjiDEhcJkYiDRE8v3pogMQAeNN7KcM9XZWiABrDtJC+yx4teR3BL2
qFG30ACszRK6s+Mwj4Pfu0qdt0mE16EaoVyAZFo1+knUJWQ1eLpk0wWnkinAcipu
uQO2g8W0jzFu8+90xGzB3CRvtGzwaMNKFS2oLa6w1sxA1eboLP0wkXcV9wDCOdFD
VEVqimsfCugmFW3DscuuhnA1/l4u7ZdMwrOWWzcnVghtNM6HWLPnCuFxaR5QtZbs
bcajaSiRbDMlVGtMEsl5NGCBY48q2EzpbwKoDYCX/UIAM2F2vJRwDKnG5AsYKQac
l8bHuRoudwlIkplD4dJJ8BKs9jobC9xiweN3YATtL267nb07Ub8fMVd1KcvGdYZ6
01ignGPniFH121m0Fzqw12aJm05rq0VDTIc9tTN9m+fA8F6SJOtmbfBVpw7Av+Zx
gk3AVUWDf8FoS1EC7FMRfez35i8iu/PJssJFJ0X1IUhGRs/I3gC6qUlppv4AsPOj
1wabllfOKSKueOb+FoKj+RMfUDDmVkk9bNwSPvUaFBjLz9YYfm/021BT+pEBGt4m
HWaoatwwJaznzmymsdbZjunXgiqZpa4IvYiyUAF9B/aQKK9pcBCbH+jC4EHEnZn+
qdyuGLXgGlYWldXehsks7RNK4ri4iwHQakjAInlu7ObGPZxghedhpghCFkRf4W8d
t23OjJ773kPTEFIw/7hhnnhFFWEDufEnVPrHk+5gUgjE9rP0crqa0DfkdvePEirW
d39isv78U7DZj11NqxtPlZLEos/ys6DIQmZRKjjGxtf/1aAZIuX1HrFqo3kjHBiE
wY8MpAqO+S0x2EPlULew6DG6m29U8wD/REs8ws8RIjI/s8XrEJN9O1MDPffzMDCG
JHD+i8mpdEXD7EbXJ3ky6yO807sbESs6zUhEyqV3EtewTQhCBf9j/h2YrMVzG4br
bfviRcYRtRtYUt6c/RwD1IOE9Nauh0nYjien40WAIyI/7re6MR6FkYZWYnPQSyeh
gwj4CnKjfDfMg1D1JnvX/x6/93dXNUu9zXKGlsh8tyu4iMLmpAJlzKtGE+eAfc5g
AfQOQcjgX0U7RRt5jWrpyVQCPaGDU+CRShDkr6+8m1+I5SMaG5pC705jqhO8TL1Y
bLTdoi1q9Lyr8UDgxzxKo7aF7nXAdQoaDIpostCSdk+4z4SIrvnjHBq2rR0L00hF
SHHYpWwWT/vXSSPxxD3+8UBYqvWM95uJJg5OFRmKslT4Fs/7A4tU7STucVvcF9Cb
Ny9WHgNnvz8Ny/KtP+iu9xCBbjFmHBAAYyHIigGKtyqJu1Yhqqz65tp46eB+Ej+9
h4zOvTyweIFcS7JuDIeqHrpVSItaIoeN5mpJWXv4LNUgc+CrJ7ulQ4UJwkpfr3Hj
szGp0SjjzzlmnX7WACbamKdGaIb5PmTItcep6AN9Zi4CJshYOoQ1YTVGBRRhnsIn
vvtd+sWhI72IS4qh+0kp9rla+aB95ljHwM7h3ez2G3v254XJmxYNzsat9pnHdniV
m0hhVdhNzs9PoA80fn9W4mFAlA5d9focvJ90NtYJuiPo3WSmBQRFXZrNKlRknn7u
iHbmZ3g17/fs/q+Hz8bUn7jngFkO5owxtj0xb4/AVVnS4g2ahx6pVXbr7BVnnGnE
ydfkT09A12twWSDb3tlSXClcz/zEZFkMuyNf+tvBTDU8TaCCtLJ5rmpX/+lPb3ka
OeXwZDvKH6HHtDZmNPMnmDvA1AFKKhg5O9uehGBRuXeykvZMnyQjdOtwZr/bdfDx
dN/dPNRaXm7J+mGSFDUfMNjJnhoP6bbBKfQftmfLwHGgdbIjkMBfbZ7Jc7eSPSu0
9Ks59Y2OoJseOb5amM+d7GdiLjbBRGfSQh35rN1M1+DpfrsB42apGjjsr1Q2Aj4T
sEaK3GT63ryrNtujKxcs3GC85eM944KPd6ZNIG70ToPFM6feKUys6FDJuIL5Re+P
TQlaWAcskyAy7i7kvFPd7qAjNg8KvjavNJAZwZX/Tgdhr2xIvMkb8GOvbaxYt5sz
ocfwhcBF7lsY7TKNAEyOzv9WRyTitjMb/38aDgmqPA17AUyHsmm4jd4P0odcjNyK
ag+5s1tNp2DVMyf6gAoUyXUE9c/XzyrK4MSusc8mADglqCIBiiMDf+v03vAQpIMe
9xOlEghxfHL6pDLN2tiMdDsk8ne66AUWkKDiquLft7vymZUrkPzXvcTDmDMJWl9T
hdDPYkP1ZG5Clw9jZLKwAjMwz9X1TfYadTMdK50vpNStclPmllv2FnsNwAqW3EVG
EXhISfOMrld3t5/sqha00arO2LqYQWy0ZBLI5LvvaSBC27ggRILfTYWLpT8wZLxO
j6jaW5dzZfGgyvXpgpI0U3kbyXLyGSE2zNILFwV0cCnOqhogJqHZFCHdwLqQj9Qo
FCRcgKN2G4V0O/i3HLkaAM5DZumnc5FY46jMXy6wKX79sF5wRYFSeyVXg+bCAfQ2
XeETmqjV4H0smb+SGnW3xZMUwdXoLqoH15aoIdyNM9ON+2vEdsIIzGCLKX8tGat0
u0d7GmrLkglijWf4i6kZb6Dm1Y1FR3RSkJuZhcp4inEV8L+Q9D+SPQ2GHYS291UC
E2XvwXWfTC41tmRF6P7CzfHuSgRTopluwx1AX8OFen/IpQBcDCyxYW8Q4Ke95Qpm
8BYhk3qMFduX4BsFOUZh5hhFHuDojnyNUDeScqucG1IZSLijQOU0FxfQctippu7N
EY5AlrqsxbBXbIvyghscV/ONoRJCvHncfw6uNefu8zTf3CeDcFVsNCP/Yr7RCqvR
7KDEqOp54KQ+2Y/BIU7mV0CnHiXBVrHWIR/0hpz9IxDriYRv1s5KKcvGWJI+2dnB
Qt0K+BwZvOiFEZ9vUX+nHHL7LMi3tCttCJcujsKVyd9I/45rp+JWcGpYD4pcAnvT
JqZPuYrg4KS7nm/nEwpI89dV2imwr08wkye05P/UcRQFkSViigRtm1KTbxvQTVZn
swfunqKSXohDAhBFCVpOl8g88Py6z+R2L0OBdWFGT4wULLvCkOmdN8KXuz/3qO5/
6C1v6B9kcIp3ioy5j0moMwcULXYyUg6/970KwFgSV0kT9mmp41YACDQzdj9yWc26
wxMXSTWsF/nFwI/oJf5nioYhN+tbj3bqhSti1A9bqniTKzd5q7YMQDlasxcGafoB
eKw05CLEu5Avi4VkBaMytxd4mK52uUXI1wa9+AS5mvm7H628caHr7BqAW2zu7USD
cwdrqDHakB+FHOnjggJpomw6x3JIJgQxbYZJWTycEAiYS68zyfw2uv7YL9uQ5lBU
CIS+Mo96WHsluRNbdd/rZfG8yFjRYdJzKEL3HbW5Z+k+EU2sJKIOEV3wzmMNrE9E
X6mJkqzfUPYdbsMfdFC2PwXvP31mwYUmFDIpiQzP0X4z9aokgQQtV/H3WmXzeXvy
TuokGSa6Kt7yOvJoJRpqVYla8CgTu/7McKX7rXZ84LZdSAaVVs/OuaEIi6PILnum
VSUUlWn+9xqQRv39EjtjBX6HcoKYV82HmLRIAY+PJiWn4U4YwHWW6FbLs9rrIMq1
BjzVFz9/xs2K8juCHBbANRd1QOyVkoI9z45feS+12DQnR3HxZGF08FkSn6ELPnNE
4DjluxTCijLBtBJzDLYebWEuHx+TVyi3qpf9vkk6phYJZa2ElTsm0JYkDunwHg2d
zIJWivXet5oB5/mKa/lJ5UdDVSSPcm0++f3FKKhjJzHr7czq7MJDdbTCcjryzSqv
vV2uaBmtoOzCMkZfDTClJzQAn5qVRdl1uSXROL3Nt0FT/9xyhLdYezQs/eOoXe6w
WwjUu4zxOM6VHRYxA+O/8A1mvIkNd16Ut/AuBVs6ZqvHa64y6G8K7E+r3vjFz8jZ
rDkG/yK/2h9F6tS+j9SiOcSGmTqlBoeOnmV7TZZP4zDdp4KM/E1YSQc9qbhDHZuf
FqIr84688Vd8qElOGoLBU/n+pvfutsmdhn530/5PnBiRmWMRA0s0PaZpqVLDXcSY
4RBiiFSSgDMHYTBzs6oOuXRwEckXR0uzf50Pu28eztycpnnx19r3wVEmdvcoGN5j
5RuyCF9htcvhHr/+CDVlgAvNEmoj5w/uGmlR48OvhfSyy7SlQWDBqK/wcEtRLTL1
MyZJFwqWKPyFx0dIJToPtUTYxtAABbHIsJDmnSPfKESwwsxM5zLQgubTzDN3NRSd
cHijssvsDZkh6csLNJK7jDFPMT6TORUGFm9juH35syYoy7XRrnFRdQ7VftCidop9
T66KFghfB+tlu0djHne2Eq91sK6rN3ppDo/3jBlPKVxsWv1FCGriwwAUH6CBboZp
IElTsUwsr0E0DdJB6kWVK2q8W9IVliFrB0k6WdW3aDw8+/Ihis9K6snPH/Eo/mkY
7OiqF3w8GweKEzuIJeMKw3efoCzddm4x28Jg2i8KNKQMgIKmPJ7lgOs7Zg7IOiby
Di/9Jr5avBLuDzv3C0ZjwerjcoiJPre03NNO/oQVjok4Tq8u7+XCkNQ0ZDtCTuAb
Qfz/43M7w4Wf6x5qaKWf81w/t3LVO7S9NGbtx5bctIPCjXT26Y+5sF+ln59/oc9Q
Ts/Qvlr38Th+Sq3JpgqVHauBDn0pfWCPiyROvKIxicNXizsyszTMxQgXRCxVgC4G
x9/Dq1zYy5XPpwvgxG3H0nV1g12DF6CExNAdUjbMoOdzlmvEElOZtsVv5ZG6se8u
mCfufSHQSzCm5JNAtr9bXR1pXljO94Z8AVC8zjeWaIk9Tu4KK14W0dUeE78DiAIj
Y9Jli9RDqJgpEDdF+g378BwxRcajhWqxKMEwRU6owq3wFFTz0UWTvs7ZcmEYW5sL
Ho6zu946I76OAM+1qVgIe069zOQKVkUEUhXPBCEiTWGlXWi7k+/tKpEs62b+aah2
+p6g6stJapbXqbB3LMcz7oo4yDfZ+CxWbaY84d8hFbjmv7J++uTZDfzFzT6y3zBA
DSqtHV0pAfmbf40VRzfy4lWMpST1U74RxVD+/ooDoDOX8nbB9z/4rpPmBfBDdKHC
8I3wFjutmpvG4EHRxifH3+L8Kw3bevDpwmYTssJFzLqwhH9r7jayQ1fpFdWFCNoZ
WGFeSnohDoQMOjM22mqKPZ7b86xOEZDkSdbbTGTUKUgdS8b3YLeOvYqWocMOcmA7
lT8unOLskFTX5fLk4A0JabobdoSHd7v0cxs9VnMYW4P3Puw46j0uD5v/o7oJdL0r
r4OsKTYDl0Aie7BsMtTUwoLIS/LAagPxU3FA6dN+/WAwlS0Oc5ytBMjq+3io8b2o
b6wWLGc8DWZYvhvASxlD9aqRGhZ/PAsBUOeyI4opUMov4kTk+dEuDdTMe/92KoQH
SamUBBdvubmygNAiKgIokaFu5SWuTQaJYnU1jbBXoqqgyqoJKay1SnlhL+fmxDsm
AcWVKl9CK97VObQolpBRKApZ3maaKnWp/Re0nHbX0PPhjWkf4l69djQaLlX8nzDT
af7LeJ6C+Hc4JLx7VgBTvY7W41gK1qrThdE9j4z0c46Rr+HvVW690T8TPNLCWpt3
mLYiy8eN+Pfk4uWiAwhYZp2w5q+GIjYCbhwGrnW97hxeOX/mcoBvdRsBzrc/HtGO
qA1bpkIKei3NBOLRHe/7xQ6o7dkmov8M2REUMKqeP4dYr+evtVSXk5/38GrLx5e2
+kljoNXUjGnqgJde6nINpfqdB0WajkIMoVROFhWH7N7bTdFZCBRh9frsXeCr2ZMh
lnIEQwq3Ze6tsdrSahlxHnXytRNMHWazXI9pj4I2Hwv5oG/Cf/Mi76ieH5FhrFxm
jI1nX4XvDceDayBsa4dEElzt4YKAv+zFX00OVUqyT6uf/6LY7JSJRHqij9coNYZR
qmB1KGzYuiAU7rKJgWy8Dv82/D8fvFvx3y7j1PnDiWbVSKoLD1tEYB1zoZfnReFC
D4UgYAYlNcv7MMMxZlgG/zoxVLNH3vyFeo/ttQfAbo0IBXlK6eY8b5M/LdsS2u6P
hu7cigqNuWj2QSxTSWi5DdiphnaURQxBIqel6tX0pYFxtCKanZUZItSeTEmLLLgK
f17FvUUwXPuZVJahkKqTgegMBN05fXvOJw0bCsvENj2RQHhfjoUZy2CC4j3a50P8
AM327qMTALNBP1K+Zn6ArLr/1SgYOR9IhqHboWPsdw8bJ69nf7QoW1WzDs/5yOc+
8DL5ump3ddV1J+2QHgrTKDTAiaHVH9btWYav+zryPIEp1NEpH+0Y+YtnlTIqS2h+
V/Lw7w7CIaTzFAwcPW0fkFlEaOHD2l65qpYzLDbDlCLi/LTBO8DNLuXTm2L9ij5N
7v44iug3EFmO6g7erlH6Fl0z/rowH+8VbjT84sVi7EajEAcz77T3b8g9adrtq0IG
8O8oYyS/awSRRne714pElFUzuAxfIZ0sfAjj0S3N5NnEpIAvG0/Qeqgko9TozfF7
ecWbI6TffY2Qj8wa9d2A8WCk3RhVPsAaY04OD0orSnLiLEKSsqSUiRGRhReUkOey
8CM4Uo5rWqShQ3vhYF07ZTu5462WCjenzWoiwDxZh6F27gj73SusEQ4j9jJAgDkn
djAvwbtyqvm3W0Kb2cVhr2ke74Tc6e5HV0uvP3umjiW+Ut7Xju6Dj5ZmPOpXJljs
np4QLP1ogwM/Er6Ql11rcBl1yyy95aeeiilVU53FcyhBVVJcGzQcEhhZ3GinvNTo
+o3KHmJbMPjoJW/ukbrzKTap3rB+OZczm/SRf7qeRX84CjvpmpfPIA5w+DEkG7zb
RII487GdqtC+409iqm0W5NZfy7Q8YshevqxvtYeQ6iy9B2CFysoOgV2ULbre1SQL
P0HjyBZ0J+ye9TlHABWGYbkx6RcJVlLdKGAhQ5AswGx4qqxKnH/TOh+qAwOV0jTK
Tf4sETB6Fq57upUzhJ6krzsYXdZ3YVYlSqWs2/4OyLp32+GmjvttZY0WugRjKbRv
Z3qMIVpB0OSd4sTFg3bgm2iffOf1uehet4tqoLzqUjaCbfmiQ19qjcvpa/HjX5bI
7CyE+7UMbRdyu9p//UukLrw6wsyl/ssaUweUfGUWephg8b4pSK5SiggPKJnE2Miv
mN5GEsX+T+J8GocsDr/fEkhGYfxqbvoZ3a4MFDDpQIeawU2Sl6Gb/OLk+5/4bYuc
8CIo7jpN1nExPpmHQ2WF1ahX4tojKT/BoJiT6PnuZQhdqdlY1s7M8YkYJLgZj1dP
u5tyfsMB2Jt8l1rQwYMbKM1gSgDB4YCjmc74PxIPI1kW2d22qamUqX4WbfXIVICK
hX+oHDQ6+D8Yyqpp5hKn0W4O+dUxG4B/p6TFDpG7Xps4K39k9v1ifuFP8nJqMzEC
e0rDUn9fDnDc6UuIJFjjtfL+aBRgWCUQNwyutup7Sjse1kp/Sm4l5kkGXiniZ+SE
HrmEbpb0mng7dkf5EeTHS+8X8E4q0AJ6/u91MFioH8Mb0QYOebqgsYk/mHGgjjx7
LG+pwNYig6zLehPHR8VM2zrzHvEfXnGy9DTeRFPFWjFXtEqp31nDQm6l++EtpmXJ
uP0CFE6+kKTbeKCcdk6yUSpbmwmPw+nzNc4SqLZz8zzRa6nux6RkICrU+JGEa8rX
mITykUek9ZdX4ER741sXi9ICvRRMOOyyinWj0G+Ix5DStoVv9meRh95syQEYX1i6
PVjM7N2Cl3DGNBtljMCSPCoO4u2hwwMrTx7jbsIIEFGKHf90rrHCnPKCDudoYRLU
6j4o6HRZohAY8CbeFXH0NLvywxpacZyRnEMJBbky4EmOumR4MaL+jBCBH40KPY5c
vaCr35QMUa4dwm4AQyM4OPRF7iitXeKjwn9DXN/Iizkwag0VAfwIwawe/OMbRAGX
YCNE1l/ZHHay0DIxsFyR4Km6kJz58wEhPe8onpveM0rNvdTUm9I+UP6kXfjVu/k0
Bq5kfF3597/zMoaPW6A4zcTQoFC60erPUfD0SCRCGDPlhMrjOqFl16vsl12V4PJ9
+oIebyanlN/Z7KCHxyAgmlkFVAejd0Q8XZa/B6V94rnIupcoshPIviwfL49+C4HA
AfwkmZ02bfr2Im7O9bjoavTw47Ap/cYIGttZcuowN91HLHPxDPGgHOeHvcmbYl0Y
kJfxpnhGnK0Pzx03tHOGu/Q8hh5t/s/VRCKpkVIvbwmtBofGlINbrryB9yoyycQt
RwVfGJisGps8qNhbPCM9S6QKl5fa7J0BuFIVaiQixjT3cZiOCqAaB40NCVKiajym
gA41vESPdKTMwmA8aqmA7g2Kx8kqFoN8ejznXMqhgNwJQaFs8yeEexBvEOhfCwok
edLPc6MOH7TJt9QMqAhhpl7+TtVxtZdpA3hb52wZlq4XcRT11yLwwRw/iD6Rjxan
1V9m97f9/UNd7hYWl4vST8Petzc1RSZZyKLEMBTAogwPNJmMoLMFxC3Q1uc5Rzz+
Vh9KcnGvF3MORvCVW5dVndPY5VzzF6zOTpCN7OtzGV/PWEnqxaBfS1hlA1oG+P8R
vZXkrYKeTdAoLAW22JxFsw5/lN4gcStWCAH+aGEFJhx39dw/Byz1kDOm7WTpwnQA
9/6zsrMof+4D46SbZBWxGcLehmCT7d0vplVjwH5S+wDivtfNyI+MjPIHaxLgpAWl
i71/0KfhuZW97Tk+MyNadBkkmZGfoZgnGHf7Nmt4Aku2VDy5nksPNT0OqrgIPqJV
VJ+XCyF3n7nIxyWCRThyjBtQDCEr7avOoW23/WFNNmSTYom/C3yzYmkfATkmqIfX
0Xz8whHygjOkNan0UUeFa0a8MLnxPOptdhv74KQOZ8JPcATYgTLq6Oj4oIGBCa0v
+QSNPraLQhEsusuqa2V7TCcfQ/sSVrn7ude/PJEOhYvEb2ARN0SwGKEWg8DoUEqJ
gPlBwneJKMwnPUdBPYhMYPB0E6wwQadhZNJYcm6fjMTSa8yRDVS9IHHknU8Msumx
beJ0X7RoSbrKFzH24VbCDlyhxOw8Mn7gqciEmjJlDyuVvCr/B07i5Ht/J4h1zaQb
1XBsIcbP5ZhHAmi/mYWHsUaUxr5NNu8W6dsaVcmLl9McFKOOYDh7CqbSVmCaKIlt
BtGCvzIo1slnDRKMT0PqjNriErFbl/zBwPKxSjB+oPbzwHqFuyG0VpAxEigx5f3+
sL8Py3V7xEd/O6ivq9IVwSJ4np2pobhUpBlv5AbjsVZxpcreS09B62aoa7tc3uod
8Afqx/OCsc7IUrw9PkREhoG/ImY533oNqedbKg6xr1Wwhvga+LhuQ4QLA6Ie1TIj
LNbc4/2fnXFaLz3qxmtBnrP6hH3R+ux8moZfBHYE6+HP+0J767Zu6oo53gP7xz+t
VR/VyIxqWM3G4dieWdLDfXEYbQc/3AIFmIuFNQY+fQYTIOucS5JTx2etAMltaYg9
VtIJuz7uxCKx54o5dupecPhCEvxJcbv1tMbw3cR5MsUkjgMQGdwzLqYCmKGHpRAY
8mhJaBrhzmFmxO3CJVb+BNsqD2m2AcY/kqW1bklHUtWQ3uGNK9w/yQzwIZ89HIf9
40XXFYYCDRh+oPwVYO02fWrDQWfBGvqa5aFJdPJMtmAj8iYySa7fUzzXRB0vHNpF
Z9W18b50HCizbPSp5jlJv4qwwu6UXOLwzq1wqNaJmRq85nNhcyLgLu/ZM457jBQR
j0h+ke59xu+iXSlFCJnj6EHprJyXvKpTNnhn8zKimhY8+tq7VlpikZDLLpEBVBe5
epO4rp9iZ7Cdx1tJAv6Vq7yeEYur/Zleb1I9ezZdrk2rCESy1XLCZKT7H6INM6ib
2thPHHdKTaylcOvN1lHTr4h1OZUUHx2ouFZB7T8O/6hUSa6JOEmd9UErgY0VjF7B
EkjkkKOE0lIistvc/aiO5bpv/Vi9qP8DoFr+4W7OKW0JriGFbywacFOBxu//slne
pnFdYK2TEAqbJHMswgJ+yQA6shmS7aj9xNd/fajxjeW7CiGYxUh8iAztMZR6fBx4
TFHWXu9uIfUUF5AhdadU5h6jADabrDPLHGABkvaFErMo8NT6lsLrJMFtrRhfpwPy
cMmkyDk9irkXkbPedVhkVo2cQpAdVT1FkPqzPIFyb77GO5AvLKaA+EOFT/Om8oR+
kZsY9xE2jfLNMUOTNbiUaAv65oen53P+ToGV3Iix0pgiUU1sPmXwusOFRKuf5hF6
lUJa4N5AkxnRMSKSIePiuF0RR5y6TufO4pIcw/xTOlgSqumgaN3UxggiQl4US/ht
iQKEGayFOifrejK+9M/Vn/YsKyt2185JzxzcapHGl4/JOL+mANScZnwhVfmakK0b
4hiXjpatytYK09t3oKQJuNT66jwh0c9LmTLubs43KN5nPqZJWA9NkCmBtFqHyyev
NBeR5zCTayNUbUsmFqPZxddazL6ddlCnlczIYak10PcIaPFBc89RF8dPePmw2Y+q
aaZM4t5SavFOIqX3q8KEEFoiBNT9J7AgzTycRoQbtY9tJgGX03+1YgIjAMa/cMkM
wG07J4AR30DmWmeluXZOuQ+8MFzIJfqjHsUOU19TbxOo84mpPxx9F56rbxRgJKfR
EzP3V8gXfvvBmZi6KSn2+D5YDxwcMIAOO2maACOq8QqqKaJq830rrHA87W98yXwK
t7Ci/UuO9D3F8wO4j/CisBIl+wkYZsJe5CTjBYxjXcC+c+zB2tfRNcYdM73dcCxI
6z0cUJL2hqaS90yWSKmEHudN9qTCWpS1sczOlGAqNjwPwMUZrH2MYiryKgxfQeY/
ohbmekWIz2fiFnKebVL4eFVW9UDvFoGq5se48KmeEZYWCjn94ZnVe67G+xBMC8Tn
2yGdTVv0PQi6PJQTGcTev4Glle5H1AH3UpPJJpVjCHMS/Ckw51BggI8H83UThte2
dWV2U1ZUTevNYTbPTVq1pGeKtTZ0mLTCD8AlD8gBuo/TIYJzBNvsYMG6QF2SkvmA
WX+TkPjnxHExcZEDm/uJ0hYg+kpSyhDHr+xRozPwMdQD2bibUFldw6ZbW3C+u6bZ
fGVVjG2/m1m6UzHeUy/xJeObHFOtyranAj3nK9LAbaJE76u/OV1X4rXtZVAzgL/8
RyVv7ZiqbCKRC9TMVoNNKrtVFvY9Ls/0TdIu7xu8z1jajoVnu/z5cHhyJRc2Tcqp
Gu5YWTUN6flR6z7xUE21Zlks3f7hSfXUfnnMzI06KwZTXzBH5FOIudG8OBXxfMzD
/cWjO/ChuzSmxt3WrbD2oGyIyJfJAZsVkkXgX75qQ8HHoszKMV03n13Kc0gJZsRl
oGD48hXnbQ6iWLyF/exotUQ+aLZTrmRZ0vL6NbeNYxZQWOQGFjp6JMqrlD+QpKJt
koaJ9SH6Iyp0Z3mn+y7t17HoMnhL07Xjsr+AZFOqRHgUrJNQSCVXYyTAcCwq65fe
z6vHkMZ7oDSUw5lLJpGsG0nL/TTYUP+XuzAgXp6Xk2TP5l7S46P3LBN6/OHUgwSU
s9SWLMVP9t3uRQKKjYDYdU7xY0dW12bHJQRRCUU2f1MlBydrX+fxJXzgMtZjjQqh
frHEYK3Gxb/36CJLA/7u7qzw+RvVBPKXP9KWl4Q8UoLOvR89kQxkTAr2WWSNMxVw
xo55X2D5LPI4guIzDYm0WjKe3hinmttlikcb66znwY/7OsV7GJ6/M6gwZ7igeJjI
DSZdcx2eBimzQDVFS7Ou6m8Nii7Qtf0BPevrVJjktDkI2DbpVFoyjhh0ym6Ct1Qf
wzL9So9BbkNd30VmfBmoqIzcZfqZrfV7NGv+sopgLTG1eLBkZ3VjZruVARMJZ9D3
UhXU+LIWkrY1MNHd1hrwINnn/SGzFYnGWG35JJ/dug1a5rs4XmGLmEdjZ3FcdAxV
RS1oucVRIzYojzRk+2qw2pJDHaK/DAtwApA9dhzxp/z9woYHeyKgq3HZnenoLHKf
jJjrlj0hFNONvy/wpE0kuxixiIFDe64GeGBjFwi446+ghuvHpFEPmwzLmYy9CnsN
R4GJk8pPhzD1dJgEtMl/mMllwKa5u1e9R6/C+3W62mUZHnV3IYgPk28in6LsAWIE
+nHyza57gI/bd+XN6aNQaEmgx2qCjrGUh1uzl7I7h+KEyGYNLck/+fQwg5dq8Kq4
9+83eJGI8bnjSk0W0hI75L+zSCIEwv2usAPqm9qzU9HNCg4+lrC67uRBWfHQqnwE
OBUNZuqXR5A4MM1CfP9e/8g9oisf/7awubre5RSlO6iUOisUyFj/E1TScNmKK9Tk
vfK4bp8sRyvWgbD14074f13Vj/nwKYn4sUEmpQbKwBuIfMFPgOCuuF5JZPtkcL/4
T5RFDhJsaYVk4qqly+QCO87uXaZ6vJPscHkHWzIkre4YX87VAQo535jvp3l/WNZe
OxB1VYS/U5QCAnJIZ8i9OlhV2jYuZUhgsdLM/595+jDSo0kxLoPvxfg5ezH48Pj+
NyVJb24aTx4UPKLSscJ9ZeuiLm8S9IF9bMeAljdVb0gsEFyC1fAkLURV1UHcttmg
TlGVlEdQ4NDpZx2pyTg0MUzKHhjM/bF/fDaJ4w6oz73Hq2MkQ6IPaDj0zGMjTJLc
TNrpcy2rdnIE0umQPgsHSeWCbkh6QlNBMDdSVAAIQDT1/Kg2bKfM6FO0p/CaHTYc
IyJU3qMVJfCVAJgcUyPvs5S+d1tQnFTadyL+6BnF26QFxXERXW6YoOUUVpThELmU
kiEzO0CnqauMTA6IbBweR3ro8LVC0KPdcVWG6ZaIUXcVbEXmyMme1RqmXDZEh6Ar
0YTS697ULSAgRLMAuEck1ffF2Ow3Wdh+bKu9w5yR8QOGkP0SjOFgaZettbHCFjy6
4nLwYrD8/zQj/8D0a9zIkVAlKizpsL4v0gfLqZp/tBpM5vqsfBRCbm4E9N704z4M
L9khgEWMNtTcVP6plHTfpaQXhFGCmQCVaNPfg05wYj09+AODw2H+AXm9mgtnH8K0
QdiVRrabkLNQXzMxvOBeUqDwL1DefioPIZX1udS8CRaDJSt3E3LIHnLivm+ifct4
MdV/7zJT1uucVwtNK++Gav2po/NgEJwKUy3VOCl3stX0uoA9iqZCdj4F2jLE3Jt2
EOtXVMB8DOc2CLeO1EcEcfTmKvIQc6B0tICIHxWDddrqJVv1nDzZS6cYIUJnbJ+2
AFWwxQsVrv3cUjQpNJI+AIM/yxb0jXy53LOzsTRi3hLQ9T6vwg+art7HHIq8cnZc
p70/04w6OL8+X/BS4dd1q8HidHjK9RSvnh1KXvJZl54yEyFfDEXNKaKyHUmlWxDd
YstO+oQphMghZXBdNaG6ypx7qWG2reSobvGCCUISynSNu8oZxmAIxjHYhtkAddkh
A0sIFmNkT/C2LtGwsLL29bIb5mJbvkNOSk4tuvSz9D6pQKZO59WOMK9igQBWQqe+
pCj1xMLuh43Tdbo6XcKUeslB4VJuusjGHFX5/cKBz/iZCQgA4urMc7y15fPlIry8
8kBrPlWKoD0/w1EX2ZNt9sulCGSyTuXIB0Ini7Z2ET+avm23bpJirBD0hTL4MEQB
ho0/GZpNYFPW9Gf+JHZqIcRQLYkqpKCYACp44FoFIU4RtvDGht9kIo+JP8ZbXENV
wKDqihAqtlp8PzY+Wy7Cy5JtdHVxnsIJnJRoEGuzrRuxL5LQy+0Ji6TtNaSXicWP
jrQ1MoBxhAofdGW21OB18hjlk5YKbBTAHW41LuhxkHLtu+bAtMR8p27MIfeuSvLC
kafmL3onB/YVfJSsFFwx8THnpF5Lvxi/ijrlLkwnjo0SS6Bn848+4bBU7L/rssU3
7J7ivdqWhKDmFvUvhEqOz8r2Y4flhhLJLgxvKknTJsBhxDLSeCi6F5fPCvhdZlGC
UeZNiNRCbKh6BKoxZGHJ/wKGXOk74h3oT+I+eF2tini1PHJzmUeSw5fyXXuJBP/t
BZnqiaoAqUXEfSFGicS/eotRxU1NKoiqM3lh/HQPVBT8KBSwPIBflp3EcZ0ZSuGj
oQKwyDOx346I4xDC4ovpTrQs48/tBPP/PrePKb7VEjkcADfoxGb6bliTRA34bRNb
DkltCHApQew2/Qj6sbtCtstHH97B+QntdIWujwiXH3sl41h/K2NLTSss/cR2rVB8
0CDH1j8PDVHQs7ECKHL6yMWuJ8q55RASSsxvE2Yaja1ZrmJcklx/CEdB/BqnUkwX
MMDOZ1YAOf6nhvK2XiLxQfpiY74Fe+ujiAx43FRWdDtqjQBMFHG2tl13CRqbzvji
GqUcTZwwlBoVV+iOpeKnCWNbiMJZL9vOq8GePLCn4Vf5ktB85kavY6MhwVT4NEo9
kAroM0hkzHNdNyn+kO0dexWPp+h+vLRX57C4dxoM5yGJyvVSPrRGIzvnepXrF0aC
Ai/jD83fOOQtfjqQzUSLS0+Z3UG2G7q3CHnFEm3uTTPq7ecUPE2VgsC2aZ1TnQfX
vmfEWVKLXnftDjEMrSTcHIC2XZ0yqAK0vIVO55my2NbVpFnX7GXSw+O0xaf7ZNEE
Nvluk8k5UM0kYE7Q0sEBF4WxwflcamizzWiq50a/GU2vCqAHU6PT5i2nwWXa5ux9
9OpNDc4K9QKC/TIhW3CTci4++18xNALy9HeWqOjibM9p5n8nW3IH2xHYvsFrx29Q
Pg+iiu9Fwi4pEIkpR2rSCPsoBzVdYU8RH7XXWSNOymq2VbdI0mfnDwJ0Qjhli6Wa
TZ6KYCXj3lDee/uL/o/dhQWBzc5RvVPNX8vruZ6Zb6uoEo4GELDY8R6evN6jI8n5
y8cmwpp1EUmjb4IRMCNAxuwu/XdV2FSzrOta5P9thwojnBw8ZSJ2GLjnRd2y+C1/
0fN/sW7B/pwA7Ro6+juWZLXE2XK/wgRRsPHdPBItjdcfS+P6HDOd30cxwvrRATNX
lHMa1WzhVuJ8Qt6HBxncLZlNpft8bvNdfrflo/ztfMlJQm6AQ2ES8Tzh1g9aXT9R
8LTY9yfHghsXtNWGGZNEPQf81zOm7QRoE9/SzOusyip5m2qCkIsSrCRMxw+w/M7j
quA9+JFwf/a6W0pbyWuckijiPgNdo2W8rDSGtrrrYbvNPW9VagFJN7NDFDlhrKZX
Xra2W3/PsiYYPy668JVF18TmkYNxVBM7tPVdT++cnO7DFStk6WUiPyvc6dtGYUYq
mYG/++zGtg8kJVk0Xjw9A+AmvxTZwQ0iM5BWisv5kZHVeS7qCUY5stBsOCLtt77f
/gx3FPrgnYLWy94P24IIGlj5M3ONHid4pI0JzJ/d0y2HGYzoxmXRntAcmRFijfMj
QOKa/7uaAaMX1OWpDihGJ+d5h05uguB6jJEsOakuceHdkcvPttVij/d6H560QRD7
ZeTScQ+PfnRm3fd9Zn4NG2fFNxTDd6kjVyoiiF8moByq57qrQokx06xyyavV4zg3
J8CiL7rC/qXayMM0AXDjHrnVCjIe3cPuyPP1Iksf2GKtB/Cv9KOzmzQb85uvIppo
UsJ/oqXjnvCDaJT8hofo/LKyciPlkQ3GLyshlz9vNdIzpzSUwpA4A/3YBWyINdGq
Mp8wq7cxYSoCu/qOWdnzCF7exQ2JSdKgeu5BFNAPa2OgvMhMponbsqqoQ0RBQ3QC
631Opkt7TLA56h8hcyWh2TmV36KR0Be3om7qp6UYrhE+QHWy2bZbVWwJA4RmmFzA
aXdxYkA++6QqRGXmSeK/PMlJdSugfDl2tioQBOiANfsY64Tn/RauUr2qfGl/YcTz
IzolFovlDBpjQhOjKXA1dpC7fPzkyRl4CvW/0ZDqhW1H4yt7oENdq5Nl4Vo+1EvC
cQJ7VO0yzKaBbbjgeFMSSMSimV4ZioWE9v4qRiooPOU40z+8DRvfI5H56oKautcH
37y4r8nwnXsrYQ5EHYZUvC1mWzCldDqi8ESW0cV3SWKX3XO0uCpaSoIRgghLQw3j
otxFZwSrd5TbzKfPhnbkysILU55wLf0cDVFrr/nv71vkCXNYqatZp0z3MtnyIXbD
XEOsyCGknujGpYzbB6SiW+Chq7u3cE3g93/TAPbsQq09GJo+aiAGCL0kz9xzLMSp
2Bo0Aw4htMxPW9mrWz0rqmESiVzodUBhNt/PBkyH6RGCQQx/BZqFOygAprXNCxtN
4bssEdXKsopJ0OU2eEJ1tn81H2fQYpCz3K8DRjCNR2QpxzV1mKNaW9bJAc5Pnlzw
R0jgu3vcynfpBaaeZgsoIYnJUKC06IlFlWACaEemU7FdjHWOiw9uKXO/5sSYd9SR
qdoXlMPP/PUe0UmRj59m0QMdJ4yfy4HPMAvBZIYpJqlr1VxNykPQXyuWA3RZq4dZ
acM7n36lPrSdbui2hYgsHAOHJiGb16uNnr/GbkQQBk753wYXaK9NlCsOrj8QQp8I
St0ZmLGvhMURKOy/cseZ3VYkRa3/ToxoZmujJGJ1eet1PSsgMRLnh9015EqWYdWI
BDiak16+YYbOVw3Ub6+GoooEcdu3sEhRHOB80mTZiXcP2Uu+hOenjlPbxyaKH/2t
geyhi87HHIz/GQPF7YMalFsr1Nns31KPATqxAJCnto2Gac4ZjEvtPU718xdm6VjE
umnXHyourvuwhN/+r1v0y5xfphAFMrgbqjGQSuuq+rhFBiw7qzN2C/FBvQOvvSMM
3S0Jbe5NkSJrVxGprrwmMp7XciuR1hbgqZswurnxu7NI3bOTgBIdkQdWjkDC5Tzh
qK8pLnQjZRo5ketQbX+vytYje0e7FilVGC/JKATRho3UAXzs74R+NQxt6aQaIV6M
cdSBFvEu243eSot/2v5OT7bpJWD/1NIvLf7wBLH5033KThMS267pCHzOURy9py5L
gsWsMWwCaisnlkgpiHdLen1xjJipoWBKjmuHxdNAi1dOonuCjN4rlYMTfzKTp6pa
FPnOh9VSMN2BFfGpzobKiqQ0p+MMTe7LTfhv5jhWL517HJc7c0zmstjosP+Ld39B
xl9UmkWWs2Aie/c/g7iOYZbDkHTy94j9/eIXVApa/PGSU+cWaxOdtY/nPmowFjTd
PdhJrY63sbPWtLaDzv6FrLT3FQYVNf0DBv1vwZT3HgJplKti7a+PZz6KDPtQBPQR
FOj3S8iSdcqPWUxa+V1w9Mb+WHQFmIWeUYP7dgkZgS1bQ0nVDY0qpGSf7tlgYkpY
wshV4I5TDUhAb0nDz25dLerFyoEW/jqv8PXw2O9YW+40ceRug3EH4wUkrf6DFu5m
aIQg2RR9SpBzsN/0GjDK7XzmnAW2XuWIDcmuJ6zufkyVHQT8TN8g+IJoFEPy+bAk
O1wkKDiQH1hqrDAjbpG5wE8/5o/l/qH5eDgWB/3RUiqqhFI9KJgAGkQ8G88ltYk+
jaAdlKJqLpuUPIWzJ8H5IRo6YZR9xufgGNysI/Ic+dOK/Nxe2fT/aFImqjqi7ZYd
Liltx1JgIhN5cvICPmCd+fXA9VCW+7P2vENDq3REPvwxm256eXlHcsi5803Kze4V
n1QOZPO7tnicHjIxSVXdkGsN3L9yJ3CCGlhEtfldNfq0mBnc1JjObAazCV6R0ewE
GVfZ0CFhp+vl7TnirTzwcTC3X9QtEumYCQGTGnhKUZe/eOfbXvnifZthS76bmEHr
kXetmYcGVlafTZ/ajSogcapTSGlZTQAQCcp13DcsAvSQuW7U7kttsIKT8jfknkIZ
gaCjcyQo0Mz7mhsusihp9Se2tAj3rVBMKbn3Hh8V+7QUc0LHYNhYqigYnHAhqLMs
2VKI2zu/QqQUk0DVK8GpKks+NpEGq1eqWovopncZmqMdv82rw4KMq7j9YhS5Qc3O
71AV6goVZ7atZ/SqOYeE6hc+bq/eCHikyJJmYAC2SdBJJD3X4vQL9SGDlJNj4vza
+bHkSPFxKbdPXOiEASAZnaZs5wh/ZDyc3hxj+AkXkAySzbAOgl4PLkaGWewJAqen
PmZBjPM2eIabJ0nGn4ErMaguczm7fJCqY7yN4MR2Y6CuGyptLcLBN40zYWe6uva7
6pV74n6YUeb9bW5uXMmpE+FHxsCmHJpyXixAt42wf8Vp0Wbaxucz6mQm/LwTau7o
H8YT1v1MXEbL5dIH7x1j5dd+orMovCJrufKNi8UD5NvCLX9Rykh76yK/0nxuZKm+
FUClDXINm2ki28vflbO14Fg3S6oALJld30q1k/b6iORR3PxZSAgmq3KexBZdJTjy
lI9gpglrBfjrkjQay08BgcqCGGMuO2TLQTrEf7aVZqo2vTMnUefL5O81LRZ1St0k
Eq0w2S+c03YIwrZogB0ly4hLxuqtB2bp6IhFv33UAXcDJb7oXZRJcUcIpw4CyOZQ
wiIsLe4GGeLNeZhWsmu2pb7xuAeMXszcyZqs6NKmmd51TObC41AU3xcoyIGHat03
k82Mt93ix070GzMLa9yXiCHA4Nj4ObE5u+RQ5uze1U1z/UMgXgqZTKn1/xl6Ypn7
5dxa8c9HbETLjf7EonJpSRdUSwEb/R0lQklWGwuj8LiyTVNuChnMgUAcS6tJHT68
z4PTo80JXtpIL2Ev0iRyhCMvq5zpB3ghhIuSMvSRmaM0XSWZcyPpakfmtKhdBx7o
1klJqHVt2RDBYM+TH06x49hkEkrc1UYKyw2padtF5UxnITiFYEGxlDEluOJpl76x
K3RDv+KuvBaJTSnHzisS0KmjuuiCfPMPlvMuXZzIt3D+h9R5xBlJ3HWtW39nHiS+
c1QITK8+xe4R91SCYYmN4cfnT8NfhMdGHAnAw5VHkXws2ax+XBpD///fZJ7Coh7r
M3mSGNvPwfO/m7zQfKv32HmuLP7As89wVYp5TFFV5ptj3hzfc7k/UP3XkwODlUre
hFV/B7qkf4jWwDcif46fr6yJX4+Se0AqJNdcRRpQNJLB+OP5I6m19qRFnbxubNJZ
AdTJ7XQMRGvQRK+XK5kocKoB/sLZECAOlHbGDCmAlZHvDlDs4lC3wIeE2b1tOvoB
WAVjLC+6eeFtFCcBs3LJT4/6wSMvgZOarjb287hbpQ2b9Bo0CsVjiYn5A1omhhAk
mGg/JPo6CTR4fJLQiUGx4Wp8BsWyq7XW91xOnLXYc9XxWov64hujTqTRaxBfuuzQ
i4AIkzJMN0xkjvX9B+GwrurlbMF+6FIuPgfkR3aA2InmUHPbjp2NjpDtLgsYQ3Gz
hqAl8vzXJECAhrNMRbOPQ60Wf5R2qwkoG2t+BhIs5roEQxA8HI6C8WEItkjRan9E
Mk7UKEYl5fKai5Sy0nqMWdf5cAXd7qMV0ftw85KMuTKC2Uv91iB23iIzq+93JO50
DYoEefEmyajMI1GjBrnsBtDholnLvBtPEUbqhVS4lh0i1CJUVNXJpZICrVXZUQQn
hnRldtk3rk6mDSkqLWmGl5pE4+3NkQ1/iWUTxXIhfjIUZCd3SR1bfoi/JjVwTwLx
CmSqiRIW+n6ojMQj4pYft0A1IA4GQG5p9QsF2bdMwCRrmD2e3blbz6fEw7yxso2k
HKPgJZAyNm7cqJ+xZd9Tx2+sUN09uxrEwrKeC+WRjv+JWIJ0l6oqh/emZ0fiRMz8
Dao9NpQAoR4R/bZM+UvHUExSkmdBjdb7e6AaMJfw/j1zkiXU7gKkeRzBi/29VrXH
WqQ+dIPSUCzGv+r1YAczsccM/rut9Yx9Sc4NibPmNMR0Vvz8NWi+DBlowtNqoWEk
ycszmJhzpo91yIPiE8znsKg7znIGxf48x4BHWwNgRE0jDeIlJP6VaRaA07t2vi/B
Pm4lJCbdj6pDCXN0TT0zIEEJohqPr/XbcWUpD6A78kqN0kQWeTpEXMbj2QMZXrL8
rhJMN3LsOvfKRBRMMZOWR+qaUFxwhXMVBXz7n1TxU4D4Eso+48BDTGRihTI3CQTG
zHLIxpErIC+/UDlGJnSW3CfjHr9BzLLPaqzKvjoc4EEC0v9gxqcXLK02UqJFs1Fp
rNYoWZZgT0mpJ22jyNavWFBWnX5Db6Nu0uTzqur9dZgFovO7t7gUc9TNF9BeM+tO
TkKZ91ODqp5jD4ssmwh2UlS/DXSUvXM2wcFWEdcTU2a/2xyAJTIAGBz3K0socY6q
Ik+Tk2QRo2I7xEa7dd/fyXUs0WtlpKxPYRZX1UuqjiO6MV8i5iDyIMbOpBfGIOYX
m+Cm+3W/TGqmIaY+qTjf9S1cOJ/0kTSAkqpLVWO3qal379rwcKATqzDIjFvE3ev+
rIerQF7fDRFNPQszTu/P0nn29dC7Chys8QjZqoWORb70LY+mX21Yb0u7AqOl61Vc
fgbcW1p5RuxxN4hfA/D1vhyBUeJFfTnbeIls1uRZ3TI9jFJIYACi3CdsBUtz+nLC
dQ4gqOD7xf7pQ/2CNs0hSKG0xLyp40OkdUrdUfYGdaaXcIoq2FfMvO5hmQNGt36z
wfaJ2OWdNgfXzXiQr0clGXtFtMCSHNBNKRDniSPXrZZvwMAob6DBSBh1zvr137CE
j/VcMHYfu6QXWkPE1OKFX4WgXTBxAtuuQWWdVd045S6ZPXVELYqBs37baIs9REeO
/M2O5JasRqwTwHSaLVAN9n6RzD00QWLU/9DS3nQTc84S84ie/tFikCXRXa1b2RQt
q1K+3zVEQxIQUHPNGt6MMufLuzuKpEiFYsW4gkn8onkXtHIGMwFm9ccTit+kzBLd
swLMsbgyWu9vmLdSb2qlVhvkVjQ1n42chB/c6Uwl1F3lPqYHCRRKS4GvmFEjUBjF
F9oGfHOS7kHX+9UG789RNgI+HJw9Sd18HbiVsPvrMXCJZtih9NpiyfAIW32YHZSK
jv5gnMS+u9igoffFYRpq8TLu5beBtoztN463tmeYXaKoeB/wRPLCgyf0y9xMuGAF
pKxf30C+Xr4FpasDWem6MyofWotBM2bUSo2Q3ByNR6zFL5RTU3hbUcI7rBB2+5bm
EVSUyF63EHau8OuCHFXyFMo/3MlHWXLpbNw7iZI5eDYHpL10BOtlSIo4eMuxSgqV
D1u30WaaHlAwu7d3RYG1kPB9vwqu7Q1gRSwwHKi6VbePQHnOBCtahNPI6vjMcgUu
vegzjMOTg31n53qHvZ+fn9/G3u708Gy6YiIpZuo5v7ucAQOVKGnn/2+11JfpsFFe
gG51ybQICJPqygU/SL2Kjm/madEcrYFTfHgg03fzPYT6U+XITqf1Bo2wuVdbmoFX
uUdCC4H6MXH5jhROyAE1wnUwAJXBLPbjziOkZV8tYmYmHNdP9aEpUf9t1pUelNEU
lJXBAeWEluZoUgbHRGpNFkKqcUTZ5Xk7cSV0O5nSCIZvksRg5jVb0zcS0XR9mbWs
fUiXZxj05m6ze2ygXNemrreB53CfxxfrQYhXAd0MdyzeHxpRpD1RgV9dotR2AJPF
VpEpYLCmk+jL7PoIDBRauaDavefVcwTsjO+3QCuyeGbnuw0jhPfICzOrF1qdsxDa
wU+kvOIk2WYlu41yQsiHehW3cCYyhx9/qo8o1j4+qeLYGAS15mNMKnVCC3h0nmaB
F1TrjQGRurBoHPlyUPxS+pPVSDeq6iA0Dp12g1y70S8kkQKOkcytT00TjVJ3oOz4
2yRDqUs5S2XV+zXFQx9cvz4PhAUvFzmRKbPm3iaYy+zSlE7CU5xCj77bQPWO4jq3
s0xWEwl3hCMcUOgRUy7sBwGugN/tiGZZcVS7q5mJ7Y8fzjZK6ndXKSo8QjsrHzM7
MsZskDYYNLmBEYsaXPkUU1A9J79TmLS+5qvYGUDV1QY+MXQhW0fY6T2EFHiH1N75
GxZAQtQ+UqxkDGeLnZgIhanKDGrw3GdftFF950Zbx+6oQ3bFvUQgT8YCqECIU+u0
NED+HHrv20g5RkJBSCRBNcoHkcpD6eaKPowaRHPLHk6RyuF8jalNh6yaygzKyF21
+ZQh6sSVAgtum/Aibg95o5FeHd5NILhdbiynWbjAzZJk+rnbYfzjr6enxKtUVEGQ
Csyj/m+FUv6q4am449V2lcYniga6SnhcAtb5m9eM7rqxhObKo37nzaLHjvB5wNyR
KCl4sOue4q0KMWc7Mw9OMLa+bKTo1zrLlYTP2I+wTe6YUSaLsJgPcpYwhaYmAfdD
eJl/DVtOzwze9pWp0NUzfoYj3twVij0gz7E+N99iT0db6kJpJY7NTng9PES4NPzR
UlRP+82ETX7TojL7VTzv5R6udUXop0tD4rX9nOSR3LE8SAubZ5zfgu9D5meqRzCN
frj4PAVN0EYYXXLRAqfB/J1c3vGiMZjUv1vo4pzLyWQIiItwmon+ujttrn2OIkvX
1C6r1du9xpIeCLGmkhmYXNCDSYSfhlV9e7/ZoFRNBGKDOZPTrF1nigApbIdrxQ5n
wHdB7w4aIuoTnTJ6nNGDTTTU2iXrRdlWngOc2lFQUfy6htlG3YWqnHVXMW2EvOmZ
meJLvMPqY6DQUrjs5fEoPxoO6pnsSZVb/v19Dbe/FZCqYfeNwRQRVqMIZasoO420
MOshDE/k9eU7b5qk/jlaUImXAFTsrF6bWZhTKXpXHNmmCmgX51m90njUk+kFCiBy
Y9eRBGNg/Etb9qW3Aoaao+xNbr2BKONZkW7ZeZ6tiMH3Zq3WRIeEfgi1FdPxjm2s
2Ph6ajv7RfikTP1l2dMmdUbi0G6gg8ejKhJLJ2K3GgCkSN+Kej+FTv3oocvdJKHN
5OPsuBNzN7vaad7V8fy+NWIqtGJGz2b4gmcmgbJfPICBjQUO6WOpdjjE+ZEr44uX
qdf8ifjXkc/EAeCThhygLVyfnVhjc/DmhqDoJAfpNitKRBOEwbB16/+J4ufFjmNt
bNmu9FRk370FC5AB5KARUH2ZRW7MwKg3kVdxe26CoqsVy22YMeH9uyApcsQl0+ik
rpQ3pO3xcICFUu2SffAhSIvn3HQuA5Jtg77kGkPBcT6sU4ZeR5FpqwOsh+kblUHS
kjiz9QhLL0nNPjL11GUO39PwYnMSOxyL2t6KrM81Qun/NI8Wz5QXiLulUWFuF5it
bvhLNaCz9L9zmRc0+dWBIS5jAupy3caAf15Owovj9PJ24T3loVweco9rm3yRJTOj
2iz+u976GWaxdDajr8CLDTnbJA08/cfbfvRgd2JDjM2tKsSz+gAcp+KLeBsVKIrG
IHr/CRGUDtLy3B+jz+haSINvshBtWpYFe/9R5I29EuMplTjZ8G35dHt6xk8KEm3A
QYJi5Ni3NT1VgYF4psIGSQeCbiyn3Hvj7Dbd889WrgeKP6+2uH7PuFxxFvWCvvvm
BR+317Rg7Ve3bN/siGZx0wwq/WWr0KNr946O06EkNGgZdvGMLMzIjWRO6/CeKW3m
vo7IcFqOiES5TBO5nOsZSp1U6b/gV+oo9mEAdcY5RAuvFPyTtjpPT4/7QCXf5B2p
IldhbflFMw2ljbsbktrgqYeUl0nZ85WfWngfY90E+0rTJBlo1og+4m3zcifORixO
jBf/FFoYyStQKZv4fInHtuo6EHY1LN8d1rzKagBTJWpSrEaOMceFuExuKWtiPpmn
o14nMb6IfpbSDWOLn4qHdJsI9cIY+YKo6sspgTwp57C9V9+5lAugAehF9MPG32op
hFp1UMym05Gkzx3pSm0jtQIsycKrNuePvQO/f9LA5NqlyT+CdkI0bH9Cy40Nm4fV
YpeBxxSeYtrx0DN7MNt+B1DvXGympEYrXiPslB3i2fErQLE0nniF1gcJzUAGDGLx
kdGTGFqLvl7DQZ4rXtyZiJzJ+fbZ1eEt9/2kGIgkF+NDbIGNgyl1M56i/MHlbCKB
ZStGr+yMS8Ycdt+NyQWmxBXt9sRUbZkDOZNzSWcf2DJv2TI4DQFKPIZbXhOtq+kg
lPfjCpoari2UBcSuGXZLbfk2OEDpttMweFmsAM12NxNuZMEMc9rxnA6BegKdM5hJ
8KFQjEqAoje2K843BIM+umzZrT3jitvxHzgTOS5/wKKqxxHBCteGXdyTFi3PkOia
yEWogC8hG7OkMnblob08X5p3KyivGAeoKG6YKX1aLkGeUQ+u3gh6oHwVv/0wr/TT
g1G/hpkq0jTnnO1sSlmcTrvFfVnbZlxnmCBWwJ+QAXAeiXeenXuj/CmTgm4hTV6R
tJYzC5Wm8+14tzRgPX1vG0caIWmyXeTB7oCZSjl9XTeuICv5WaSXOr3JIzld0n9n
RdzcKFP7PYilp/4k+oybzNWqAC1Pdb5mmCQfPhA3dvKIaTbKaOAjkszz+QZ9PQTK
0HN7P8IMQqnHPdr7cRKorow71f7m7Zbb4B9U2rnhojeH4C01gOKVV9oy5iTIRt4J
0ghxn2HB0AsmpD7m4zrBg1fXMeC74c59QQTs88yOfxg20mKsImam7yp16wUBu8cx
vshFtD7g+MdrCIutvw8E9xFDFwvBT+te0oLr2u0k1yxmVfDf0CniDeWr+Ygip2uu
9Dz6V8oRHBLQZg81i7/GZXDkZo4y3kj+rharQ4Ccm48ZRrPkwKvPprcjKLzVN2TP
DOIzQdwnFbZ4KBXz2eDcfW8/KMWhGU3U2J4QZDTbr+EbwgFE5g09SK98WwJhfnWY
R6nvV0sX16DryjZai5KAADfIr++/e81H7nGUaWTPsCAKJIG4eibS1DQbemdsrpaZ
7kUZdHNQqMhh9VkNtmVm5ZLjE4Kqg9zI1Ce5+/VDZz45l2J6mzeAuGakz9hu0BR7
orvMNbrCPne9Nkp9CNHmNUjCK7mDjzLCmNNwkIs0pIRGtLOBYyGsPggzJKSFHLdL
AH9ZO4dI/XQs4xSt6xCCwzH3u/YQ5lMr+qmm6bg2Zx+Nw4LCYmFEPvzmycChAh3h
9pbq0cFH8OQBGam8mFuzGO25Le9EbGKW3AB+r/PSHeR1ZtXYMHx+mdkH4j6Td0XH
Ch2kn8f7q8bB+7nSOuN1F7iyYjAqvwS7Huj7VGsKtcNX7uxM46zgEUYi4M1iiaW0
6uXNaFytRXkInuwSwI8nuHltCeIYF9iZYeCTMlxLERlKkktTSY2SkNEejoL5SA14
jp8Ps+ny9suf8TDSJu/0QKHA4wbAkpmaw/59cNl7Wa2J2dXBw/tiIMGK8ixcuYGo
Eq3xjVBAwB2lsDftaQ14NyUpXrKTAPIo9+M2f1Huf0Yme2ALUmWtis8u3wA83yku
m9dTVK+R9mOwlWVTHjkJMVHH/7ZTLswq1eJyI4259M6WjQejw+3vOKMDaieeaaNz
GV6+LGjZol8tAzYkIerPrQSrYmzjfu/oLIEdNkuWDPEnVp/2afL/+KkTSibuDetM
G72SE/IdiNvBu/LSp1iY6l17cM7kiEGSyzp0FIZutpMZMqLdVD/SRV0X76iByO/K
0D2Ed7v4g/j052ZIKPztgeF423LAtzOMEex7kE3QG23Tp78kghea32Jcgt8RD90w
qzcFLMCF/t65wWjEmWp+dtErFfaG9N18Oz1bdaoQG//zegSkPqPjBTv+7fSahJ9X
gSMRtrMYLNVYScW8YmK2cbqZxKImO7RQ3NXpNo/L/YwBXxJkebr3mx+gn9pcKLZt
sfoq44ZZrER/8CY7ss9Cz5TUiuZ0O3lxMrEDyf6VWlSeX3k1DG0/dnK4pxRXnd8Y
TClSYvMIYwK8c/M9cV2+f7yBUCQp4wMIm20vfkBXK1Ql2F9cZEbC5aTVxqfKUsf1
EijhjBlZkGgzzslY42R5MFymOPsqp1LJVnnEVs1nCpikc358oWJNrrGxzOP5qG9/
K3WXM5Og7WLuSgQ5LHvHj0gghOqefM1x4EVQrbhPvYYJIntm2WSU2wsf5KZulsoW
ueJvwtWUEYI3wXNf3xGvWb0PCiLMfdr1+Iwin+3ET7+1o9rxXhVNE5LmvnN7tyw+
WVaTicnTatWQUjNUPilYi9fo3bCipdS1j/OCLEN8Q3XNw81O04yWOwcN93i2CDzX
zzHSXkwpTJlimmY3WVsA3KVdLzT+xCurtDgQIrOS0vR3/NKlc3rO5WgWTQyJlVFY
mKFnojc/o5xTRD8s1w8nrcmwfPndfT/Enkdk8zlnrSCVEI2dHeiQ6uMOGAOhQm2G
QnH0CJgvujbNuDt1MHitsYnUdizvNT6QH9OPa3AtBkwhNRFGfRbYMZCigjaPSu0/
y8s6WrEjO2vnI2s0acsYYgLLUGsl5cyFA9gLUFF/LlkWm0xObioqRqVvkea4puyf
8Rw4TE75m6tEJoqNlePpY6l1KH41H2tK7iML1tp+bETBJiYjrQ0gSSmTFsmiluwh
1l8mKYxB157uaApSEism41N7bG8gY1lqV0dxXGQzCFtIALKEQ7c5LzZOJN/5RxiK
AG1WtHODEui5Pwlx7hXY9nSkN/2jph5wy/60h7JLtBZ5+z94ziF3jPtRJKMcXj/h
y92jHRv8jgoaejAF5+SmiDbqfQxAY1Rc+WUS40Fjl3ijT1PG+e6ous32Cyk9HWV6
M1WYTUUVXLuwnoRYefrd+n4n2gOR47GBYwTt4kWNZuLRYaSUyT/L77SCejno30t+
Dlmwkwg79pIu4Th/8WubhW/+RPikR+VxTd9fyJhjkRyWgAAsjR4blkiJ79V3H9T2
LMjjTO2ua209a3gGdRfmuKj9JBHQ7zD5dhPbcD4A44UhHLI51Ux5hfxLGG/kzTx9
W2EPDkO/N6LGMdYbqhxoB9BBJK3fQeTgRaYZi5kIfmig4e5nDHdz/IxnEvHGG8nU
sGWfzUppPVECaIM9uksDBJcTyjg2ImGk8Faa4U86L6+CuVxsL9YVMDNPMIxhFHkF
QgMlvsWrUUDv60ibaw7AlLxQLeY4OXkI3ziRdrN4yx47O8g3h/ogug98Loz9ApUg
5qVjLWGdYUnmHjXYsPOVAZ2VZPpEWa/rO/YBp5J078vwfpLgd6i2T/XvkDvY8sDE
ZmZ4qbC3bCpP+Z5TV+i96TQtjZ6X4HTvHgN5XMjpqZ/6XPNpdSvuuzU6DPGm8ly6
rEdnxRwHTC9p4iRDcYPiGW+D45evZLkbrkQKIATQcWWMKRpjuivuKuiC6MVo/4G4
M/NoGymi/1X1FFNIsQDiF5NOaajQ8T6eeLc6ozFYDIQg71oqh6kdYHNHZiAl7m7n
NBjz7/sopBHuQQZGKgsvr+H5gUfVP1OvQvbUM4qDsvNfwlu46Oztr0tgyWSREhUs
QKTYJkLj0l6iGLOundbWDPbtF8otFzqocIEmAnPTboTHC+t8IUp6UclxAWI3DajZ
ZcSCqc+L7kTpEJdeYT/TS9Z6vdGDcrc/rd1+aQx2cRG4ZjbMP//auHFMaxGfigOb
5X3vGCbDYeOTFdSKOfRl+DXwvVVL/s5PAJIXl4HSzJhy/6KWlynlQgKaVw0aVjjL
gm3DbFmcB8ySg0hxxrQyN2/UVX/pGSq5ga01pfhQLx/tfmZKuLqufDfNbV6yzEJW
IGJxwRrra5kPBxSi/e76igsvr8PM/4GlQkRDNCkL4xtg4DUMaQIbHW1q7ZTDLXJb
WTK2lBNpMITYtN6bi6XFusNQBwnGPp2F6JYHg5zNPfgpQqmZeDr+tBrIUwqJcDfM
8g8fTuoe2+V1QtaYt/7km1mWxWQ0p+mesboA9vlGEKWFdFaEtgRMJVhyqb6uO6R8
xmg9H4eiHYpGx6TMPIN6Z+A2R+igxbjGfTcJ2qYlj6K3FfgyRMMfYo7bkFHtyNg2
hrgIINk5ipJPUJfICSr52J+jx4rUQJldj18whDib8cqhbO1mQn52v70uGNCOv6A5
IGLjD9Msg5J+tGieB6luf90Uu+P0dPD4AbTlW5ipFFOLd1+GYvGjg0E27mLmBKBu
DfaDBlQ6wlvEQ/6QXzm2rjK4POsNRsBKFrQQySI9CaOLWALHdp7WUAXWT0HruyV8
gtgm1RoDE9j0eVnALykVn50vCdUk4tvJFVBZyqPnW2ujOiEz4ybvCaWCr6Y2avxD
dkPaav0T65PITWAl1ufeWyCDVCTPSDWrzcKrX9nDBVdizn/USwDsgcR19jhe0c9+
JifTawMtCHf+zmBqN9V/TyzJJqvGtutH4vfrQimYw3xgX9xGpGtbahHnFdnDs/Zm
n1IC79GQhWBBn6hzhq3iUJe1su+muxeM3ukSQCqvjAWi8MFZRlxZzcgk3C9Xohgc
uN97S7/mHp+1SEEXcfIRA8N3iXsmsYSHNWEosGDtdSb+Qtk9pjpLhyYI58MZapDn
spoE4biRegcUHEFMmj4rjJByWpVzSWkpjPilBUr3GJ+u6S56PCNbI5qybphC5VRu
1U6nLfRF+h470TP2EcYOEz9kjuW8tPx5sQJPuLzetk+paKxf9khe+K2ZME1NVCJa
zk4L7XVvCQ96zglFxtuzilQ68baHJW7S8AFKDLuPtdBQaKIps7lvMQAgUAa4HcAo
WtLW41/aGmrwDQgMOy926TXt0OFpQiJOXVMZxxyCrXXsYJwL9gPOZ+78uYo26fWC
0E4QCDA6k/IrL1v1uUmXjcaEkL3cuiy94YEbo4EVeEoN9sq6smoYISWaZ5Bt6+de
n77kgff5UWZMgITzCoyJELFvZtKnr1aaFdi4j5cMs7gvkLcjDoolRdsBUKbWhc3B
DV26PcNaE/7eONvjNZj/gsaffIbuwzRhmhiY355idyLmb5wW70LqoThzE6C2a5SX
W+0miiPcvzxmaw61ks5mV8Inqy+sHzsaQi56oFTYgGiL5UWCcY2UOmkrk9gGe+XG
75nf9ZTicAyeaEz3lv/Mt351pL5w6ngVtoNnL1AJiswFmQSbu+2ImjFfQhq3Q1cv
3Sa/AwWev8Vqx+l15vdeGs73Eh/6XLmfemIy0A5dxTUxC67WjHBy8pzezuCFVY3V
z4Snkq7wZd+XGhNa7S+vOq5NF0zlsP0eie7LY/4c7LaKtztHBVtXyR5UnZod1Kq+
cwfulb0XyM3Q7yrVHtyyjHmKuo3LARDF9ZQkSTLCRdtV1EzDN9zSzgwNCp/3BsEO
SvfQyOhsomA3LI63wv4gYSsMcAwt+5/0wqBQqEycyjqHK6PdP8WOWuwi+nL/6OZL
Q125bxNNM4o3oF7hZKZFjmSoVSl0WL5eK6VK+ecEJueQKgmOODP8b91RIEeWhO9X
YCVKXWeyhvsjPLRo+pJ4eo3bj95IZPols3+4s9JpsDwlcXdnAx8fSSvaTvBddGjL
XG9ibluBS6sUnPLdy7KY0Kws8JeUlz0hSTauiRg7mA6BHF77faXNiDSZ8ydFM0kt
egtsqDzbiQZzg5qfwQ4R6X43DvqPrgoRTYZqX2ZuwDYLfAxziUsuB8hCJBkJBVwv
cnJVKA7AE72fIyTJe6wKBp4clZK+A5Mxl2hiUMDgOP7CBnuZfCaaaxVUTsrYLO/q
qK42vIpYeMGqLLnaBvHijsr4vFnT5QXxbLPcCXh98gBljN2nYPQXNH6rQAJMBZ1B
MueEMOdDn13eoAOL4p2Z8Goqrp9saUmX2jCbFVo59meOwp+q8AV2Uv7OxKaQVQ7H
n5LW96Po0ssh3d3+gMnnq3xB1dT1UbgITRqpJ3hEo26k2ia9ApN6WgV/6p1iXRGm
HsopHIoAF3eQNL2UAlEa2q1IbM//jPA75JjrT10Uq405A7L+Lo7SNUUdKYIRL7oL
e2uqoiJriTJy661c0YYnFz5B23KLoQNz8axfPaPh7DjSPXb79AOlcFZbTWHjNYi7
bHyhYb6+iZgeZ9bNBXPTgrRTPmTFnF+ddx1YpOUcsBtCD8sJe6NZRsHEhK2tVTes
05EUClihOCtSMRX+pd0YE1khttM9cGd5w1KvQOP9KNpDEwms2PfSa5zwxVQ+LBjQ
CaQPmq5ejZHutcEdZlFUanp3ObSzh+ICaW5QKj/3IIeSok6SC7ghEPvO3QMM6dAY
zFTAsDjdVdkHwNZlCeiPDKfhT02qCyDPZNTHrScAHZu3z00xA1P95IZU3fHqLoVH
jlu4cnAfLaCud75//q3Jk8aJPXC0lv7htR2mHNtPMeELyK2CR31AdGoWGcB8xDqj
PGbtakRW4pw1nQQnp9bjSUpnOcgxlhw+nj128t+jn9BgZMpfSu7mB5MXf1Vjpbeh
k2tr8LUM9Y5rdHFU440vBMCneVtRjRUPlWtiy4IAHeyv0F/ymqa4FJWeTc2/I2Xh
jYBsng0zEi9Z1QiPw1aCkSoB3h9oQC1914MRvqsqFMORft/R6/PzlsCr8yz2pBCu
9cB96uYyskhlG2hXC/AgTsyWAplwS23f8BadXzm24h5OAI7p8lc8gPZCl5e8/7bd
9iITTmiGLuZYlQD95SAVR0m8wNjXR9uthvinOiVNUXX/iDE+4Fq+EJdeq5+CWw9W
FGstwjukQLqRprlaWQmqnOyIgO+PVtGJrYPBcSYNtH5OTyIbIknX62/R2xPNKuBD
rM11OyTqjsspajV1VkQCI3qpBoiP/5dBaJ7ckfE7PY2BmlUKbnHL6RHY4zl25OVz
KG/k3/8H9e3fTWUhCnIyeu0cYWf1+cAr1gDxaN1Usi8F1MIinfJBYSikvCGz+3C4
97+wYofuOdnLJIdKJ7x/qVmBv6MS5gPInZF4B6m+9wg0KlKHqbD3kDNoNl/t977W
z7rcd0dYAO6u0na3n3zaLK5sOZ5C8n/6xrBKXO9kOvak3gjmSk85/M50cSWLILhh
jmfYiez0iz/KQY91C4R1cpmwQeFgsSgxwT1RPWogqJcQYvTaZuqQh4BCVa7TFfNb
n1nrv4ame4V71iFW1w8stELews3ln/dSm+xW49gujubF4Eaomk9wg6haAgquiRMM
ORYTVCVlI8AldompE023mWe/xcUDjk9kkfqbOjNaKopTQ744xv6OhvPwhe0zQPlw
8Ds54BW32rjcNBwCvlSa19DUapzqTyI2rlzXaejHaQ+1Gdwe9xVrzi3C0iG4LeqA
Upr2JaD/Vi/JJArpsn0CFsmRSZq6W6cVAkEmOJ4jbDM00z2BeOrYzpSCfY9EsWiT
O7UzeCE4UIV/In5EGpwMtjBv2yWY6U0snSBhXtv1HzvC2EYRJCeAUrWhcGZHrqYz
Kxyks1HcN+IhIA5vf7se2ABA8Ma0QO3u8slzgOQ/nyHUl6K6dVuSfF7XNoyAUjIS
QqfnAwTfqPVgUDNep1GwOKAfiAy0IVNGMpEhU+9OJPEhpZc1Ss1sgY19SJJJjOp8
9/GLYb8tj8tHZLduXpqXS/zQYKI/IApfUmYv9YBWaF5qYQ3G0anl58pqrjQTydnc
rs1lmDgAIjdjE9CxqTXeIqbLxkUWTxrAWh3aoUO20XyIs9SW9o9Irx80mL0PKUrx
5M/OahylE+PGYZIH/5rj6sU2NmiqRzI/sS+/MZH+ISHyvcGbQTezKQkh5+ycpAwg
0TzFAma+B/OqNX6E7kLbV7fMy6u2RmTVW0c6va4ZgN4Tt/He2xA+kAkAvMdrfpKr
hG29vnfRfEN5ast7xnfBJcQEuptWKvYjEvLkgFR/82avyx+ftg6a4+Ygd7uYmg6q
MIHoS4CMcdUcq9yQU1FuxTwrPySKj0YcLqcg3Gls7wAEW00ZVGVdT8eqZJ/faXcs
Lh7fWmMiTAGVwNO6P8e3GLyX4agN08B6qt33HQVf/R9NpcpmIHdq/FpkRZL+DiGK
FRhWz9GtR/hWfaXlEuiJ3959ukUMVZWUTuwxuN6NRGJe7grZtCOwYaDWFZFoeyJt
ZiCzLZTMZGzUhRdmCKFED7FhSbRIi/Fvii+Cky0rh0427d34bHzWnG0ezzIFDre2
wxQFveT4g82Ryt65TO8XegMsqwtyA2x0vnnuA/QGHWzonQ6POBJ/q17bjkbI4Pxv
gXd+QzpUjg0tKVfrfJ8OntcE3bQSot+UZM/kL+DYfMaASHGOvkDA/74OSxzo/+rs
ldTlUeiRXW0o105BxPQkoxEE6thWBgNhdYhmW030uywK7q6PYJammjd8yYC+HO96
hHXP2wd/nviq4ZRTlVvkytYOusGgYK5gmZj6cmTE7vQ8ccZoryTKIcesDYOSyBss
LkuIwqoVQjpCCpMvCbxgUa4wWnhwvIOR/MzjEzOvtJ17QaeKQp2OMSKe8UBFw4tL
LAWTtPDi6Y6q92CxPWIeTCSTuyrQdNDq0roK60ob+4o/6yjYDFuvgy2v9syNj+sZ
MnI3KuRAmPcxNMTrd1PZp5pUqI3cEzpwQkNe3TvuxLT1luxECGUr9zvZIAo7WC+4
zLDeC3BhiJD3CTAw7NhwCIorOkkz0qMl7bGxAYAAjFSLzjejtq2Ywt0r+z0wJvn3
95qLQ8V8oSALYjRQtsI9ZL2x5/BTc3fiuvqGX4ZjEf+e2zECZn0XFGSa7301Rw+/
nJ6N5jkC2BXL3LtASp0FDcBGHB+ohFCaR/H5oNCI4zYzf758oDp3PLF6uc70+rh8
1VkoP6NmTJ2yQWCYXYM4ye5ztUZOH3pr0gB27Sm+QrYbWR7M4AUnauHlGh+WDVJ9
x7eG0kfKNkOZnKQKEJLLHyR8+e+hGGxMwRzRWqTxwApJtnhbgbYA5ccr0AtNh9NQ
AnzWh7zI4hBmKySDkbLbkWJ2/VjJ+rri2QJSPztV0O6YKR0o2djnEjjFtIJ5vEzV
806WwLrwdM9bGxsnnyDFFBG0Slmuc/BfhGA1luo/CpP4TDi+TN8PkSElHssdhfWD
sqDFDfmss5lY0PPRNFQtHosjpHQtQUkiF+/FxczqSH0HdypUB9bR3FbmpnaQbBzd
4zhBxO+nWRVOXciuurbAdrWGPHJyxW/TwRWT7q1hKSX/X6ghVT3K3uFND6cauBVJ
XR/gvWCTbkJwWlgYXKRGMxqp3UziU1gLv19oK0U+/6Gtxtrt2bccm7B9roHhMtAf
Pxst1MeVVq9Mp1uD6e7X1UV/ZKkiGjj2rMOgnouRXwm1nA5eKcJNao80b2i8fuD3
R2/YHWMBEZI3Pxbq9gkZ3BIsERzH+oDiZvUEzARPizRrZfvQmU8RUZQN83RjBeQp
mlsyFR/Y/+ZNLDPrkna/PBywcaEM0ycBdNG1E4lejczdHvT7uyaki77h4QtNuIti
E2U1wIJwZWbW6vONVsZ6b2uHwRy+FBPbBvmHt5zQIjFUpEFPEwEqpjw9JntHJG49
2L/dWv7D4VV2P7rQFM7z4+qwlQfG04Z/M4o8OgXc7T0zT1DXgAUgPRntiT2Jcd1L
CluLWWfljlL6dPlANZ87ARmUcMxLN/1lz5EVWG1soPvPdVs6J8PQZTW6v0ddosuw
4fQT706d8LOQlpzPpKMRyZ4TCBSDMm7FttKVDaV33/B0Fpt1hBTiq8yo8AnuVoA/
/ugXglif0YfzKrzGhnJjrC53frUKaWIFf7X70sMJ08XSJYzj+G1JL4lnW17+26/l
sDAgOzjD+Wlt2VAlsvn/mF5dWnSC1R5bqD1cMKVj5PCSS/NRPEZ5PQ6wIuCJnnS6
nXbQathncM5V6wG4g3SedewQhvGBELYkF1rZn08XA8ya0dUA1SPZExVBgcivCIj3
Jk+QgoDqvF5KLJPQBQdHBwAwJcNRO0uCAC0+WsNwsNbQMJE27auou4nbg0GFObTQ
HPQ4YUpRUL/R3GKaz149YenUOZ9iT9x53UeGAuERfqeeelpVJvFVnsfRXxnnvAsJ
9iKqQw9hpmK8xO1CPh4ewaoyq7pjMsg/4ynQX9cWp1aQafm2OmJxzqorkL92HprK
zS6r/slkUvMZFLZdsr+bqxSTrxwUHfbJEtqjSyTz7mFOAdtzppQsk3K8i8EfgNy6
zyZloMiaxMuzuBT4vR1vZPBgQYRw+MEaTmJ8x1AsMb1CJBawYoYagk5SOC/RskES
mtB2tu3DyOflo6XSpcpjPeTe32UfXGMKk4WHblbtotfAo/1dgi3hNN58l6Zq//fJ
htXrkBNDszurC6YHEAWEAkclAhpWauCmQD+busn2jrKNTAbyO38C88J6JD4Em0HT
X56IYW7VbbMR5UAxTf24Ddf1BGEaxetKSLfV4WjQ76jtZaJf91sTzNr+Ba4q8alj
LCCV7MV9+4QDIVzQCrUx39hHimXElJYC3yo/yvO8S+gZB+tuhSgEawR1vo8C4EMe
sI2DesZFhING2p/Mn3JuNc/RilIq70eMFSsHuwqBHH/JjZWvSxE3VTA2n3vAFw6+
7VCVYXC3nPlFpUSDEowcO2ouLY2zQO+AR+93nva38hXHdf3vUeaPXLeKfyuvaiEk
II2sGHLiL5V9sZy4aYq3VmUj8o+atpjih9pJujnyv8rmTkQuIPOpV00zp4ycHZud
t/UzkZjqlD+9jGfgkOfPpkYgTeE19ENkZS/iAz6+x/lmz+/eMJz3VsGimQ3cVnpt
cfohYv+7jQnCq+JsxrMYYboVSZ5MFzBxgz6qZiX31QkdXTkPdcn6CgiyZqre0B6H
Y5BnRfzmo8mKiwyoA/8zLfDl/y3okjO68k5ytGt5SCHGQ030IlFqWNMunIAe/+jt
F58515K1Bw2yicIgq05J98uzxz83IZpJY1mECt0ZEJqpI9lEv/V5XaRWhwnR53Tb
gvVFWyeb12NB0qMvImr5fuB5aRSRbLMLLx2K/EjDgNegWeU+I9H4cXDvprGD8/UE
/sjCkqkE5CdAIZpbNfhFy2qjbacKglCdmC+p5fW6A0YQHBVTHQQ2sLGhKqBiA9Tp
p85QJuJH2+4GPha0XXIoFhhdgNfrS8kjtIT60Uq5Kw0lZCjV/2i4IFaXXSvi3wSL
FrZfh6QQvhtSp6UX3obHTqtNbiAFzHJZWl5axq4UD1pPxD4wDcQWAQXLrZNxE7E7
iM2YGyv6MZJFDMGwLpYQCV0xPKlW045zfkCh+ZJ1HLTZZB9q7RxWQnObOWyPHPAE
Js99OjwGiKGwqsPIOd4h/daX5b0cS5PlcoNlKycpercR/igi3ZPTAw76aMo9x75J
Ggze/vyCB8fA5u8qWjsHcOq/UOmZfGJceZBtVpWSWKfu3G/bhRaaZsk/YVlSYyhq
33b0l8JLm+zNSEhxSzC2oVlVLeSLD1892/hrQK1Iemu+sSYoDBSY815GXUxUUjGC
aDUXUDCfZ9TA0GEtLkkOg5KjJmnRIVUJxPi8HAqGDjYKPwbS++HaXnbt4zLpH33U
W5gMUxikeoABnjfkKwWw8mQSUKQO5XV/K0jP3qBHEnO1MjqUzkboiPgpbnINRGFA
YkbOsd+v4Jv6c5+dZNlIfgjBv/AO3OoQMJyaTvTktdAWBThYkptkXxE93oWglYwk
evMxe/EBweMn3R7XOL0TmA6Eo3kcwmZL8HfW78AuwLXHt4VwpCJcWWl1lvVQagEE
M4DGA83xnm00J/rDui6ADbeJM8Zr6uw5Oe8gPhP0/LsofmuQRPLyrx1rYHhpUCOX
YH3Gz4tDdkd7+6DnwRM84GV2tlphJb7WhGQNN4/4kj1r7qGCKQ2LSjpCYagKt2tz
uwg0+Hg0dmq+8K7N+y4HagPAZiga3wH+paFYPLkX+IdmPjNL7R8+sLN3g29S12H0
u3Un1dmmo9b4uZyNwbengUADTcjHPQbmvmuXz5Pe4YlrCS2xCZiexLYPtia3nXeo
7PpHRoZJBtKFkCRVgQQOuxG3AonSJG3H/PzP4e/6w4TGJcu7H+t7sLCLyHE4rkLg
8VjZnDMRBSfgQC38V5a7lK9SwmhYFLtAVoOp3DXnklvkexNHHMIyXoubGuVJ94Av
kok8m45J885Y4o3VwZKVt16zshrdjpk5CC2XuSwpRBbQ0P2HA769cREQ3a6EbaSl
DBddJaO+kWNlZUt4RmgiiqesiuByXSzTeNxPeMaSPhNiC9eYPe5dJT4UbRZOkzXP
+SeGD0bsKaJ/CHQ0ztWAzmjAfRHDinf72CIixsbH6huXGGlhzqsE/4S3f5EVTU49
ldZyBAp1GLUKt69wZU0CVhSpKgl7LT1qzefrkocRairp2U1MHxoPlBfKmHgqaj9m
89ajf2Eizo24kjfmWb9vR6nhAQoPtFFUWAcDcDqWW3rswvRWq3e4r72IDUi9PHKQ
XIA81qUwINq/Rz021Nuy3ssqyFxg1TLxgSPS+gQt54QqW2gX8sFQmu3Gf4JBstdT
cdbDRyow5AA4aQx0feS94FPyIv0GlJSggLwiXu6YihWCd1I1wEriZmAnhrNIs4lm
OEFBCo1dc4i3yGxgJxGiOLWRaM0f7wewJfk3pM10AJMC7Hv6AxTeyfgsAaEv6xzg
rF5wIddUl2PMolDR03NmVAgx/H/YUAdIxvaednaop4fiWGj0nx239bM4z6sH+/h2
qLDcJUS1LJJrkmrihKMPwhDAe+DBxk1wG9uanCXIS7KpziEEpGoSYK4GaPqsOJJC
GNFtYEmlgxYfsDRTA+QEnkKicILCJ0tgVA9iVf4SwG78r04ih18asS0slLHgD0BJ
kP1xNp8XaFuljpvPxP7pZ4NtEzZB2vsZ74/O4H6ilDT/sTbkqbx34W7Gl5/gxWrK
qCDiBXxSI8yGZ90Ch1xxRxTw8lKMi/9+MsTK06c01qMKgPmwlVsZVl6xcm27+h+W
qwa7yDllgYJ50xXCTFBLI5r53gdWUJ7Ket9D7sx+s0iCt65FYGnjrsUny/SNeOBv
adstssOnyKgr3JoSgCHkbvWOQqNV2RfVW+yhqfbonrLGtIgCPyu/VwAFq1cRhmvi
tsu1hHY3by9G6NxMHgr4NG99BZiBj0QmkNXeWkLK2FWU6L/nK3OZbr0Mprtc9ihB
1tLhAh/nNFg6mtMea/dGixm43Y+HlTklwDHWuJzb9xnO9t593Tqv7bJ1RGKcXLN/
4eiJQanaIP+0RS2e8hhYnWHfbm8S8Zfuppsvw6pwTMKiBoVgkAiiOQYq4IPtH+/W
9uYFk73UEH92jppvBT2fqZstvy7OsxOdT6/40JB5l+5rQwxNu8SSIaLrwbOgosL6
Zj0k11JBzsVmbXC8A/p2uuNK/dqvyxJMchJ1oqNuWpkDt3IreKq7KbqZp67jd3Qi
AiZ7ajeu24kdWHY/fEaB3Yt0NH/bEva+jpPCLaDy+g1xypQULelsbFX26XUu0Lxe
6ju6q/KeVP2w/V5ICMR3BL+As0+qA8YKKR8wyag+cKhVyKy27pT6G1w9z+riLpiF
CWxxizsN9H28BVBuBcHu2Hjl+zzzSSOXie9HLh3HVbWETXnpQj7MnOBvifcGb/fv
9LP0xaGg6HPXMa28e54/b4CSSgIsCcLHMcHKI3zTKpBS4jPe5es7rSRXGJgK+vKM
eA8gDVfBq+D1wwMpE62P68PpNmNiCR4EddWofwi+kqcaf6ogeSmZ4l1hdeA4eajR
tqu0dApOUg9I80UQUursNImhNxfMdqcO/I7K3dhR1hvw+0O5jZz+wSlQqHp1xtpr
b9nd/Rsm9AOGUJE4N7Hpc+smv6GBjSIUW0oJflN6jJ+3nH16uBxLxzVtctOAA0TH
yLlQgW0s2iHct6OGCclhUy7Z21dVZrwSb1jKjINFGYJ8GLXFm30MSjOQhPtOVHR3
aP+CaezidkB8ahBgrppcZ8u6qjTV4zcvzsTltBZyGrVB7ZpnF8WE7OUVTaQJnF5B
a7LaS184uiN0hxt4/3fPH/tr6FUcCqhCTzeE+RO9QYKY9uWajQTZlUeCuDGMJHhj
clY7xvAU6QL8XoRSILCFeCE/sW5lj5Ootiy1zV6t5aFA90svClBFvj9Hc/r7+455
jrEC/U4pIqzh0q6Hs5l8mSxaD9oWH9p5gF5UjOxiM9jtYpLFHNiwszlWwaEfJJLy
2XRjHhyo6bahEcUXj2sxTG+sIS19z8TttcfSYWb0yLrcFU/7W2NiRJI45q29hmxN
gOHs8hyNN7pRu5v9mRvEuARNU/rl08jhtBX6vECk45xaT45YOD9Hzrvfo8tkoA1S
wKfzPyrf3FRuIdz8JNnxDTOqXtBuSWh7u7whqWD6x4Q0QbbPGYx6Nj1WJWZzHMie
t1LmfQsCeuqNqaUVSd3wUpjQyGJMfA5VNp4RGexYpenVKEbVTDhxVWLa6JSbpbWX
Uec5Fa3SC3jMm9M4gTHz+itu0wtt0nU544TVVxBv5LOVK2lsG5ZrCP1gflqZMGNT
8/FGtss7Xu3ATJ5eJt3aFUPagVHDdJ+lUhh7KxMjJNNJsr5/vRNMjW9i6yx0MeqP
2RNe9XZ3TcnTXvIXglRQOBbCDE81TUG6dR3mxmmqPdregub0sFZRSZ/jM4BYdt9c
StwGN7WCVQsB/96XXSrAGQO1Y5C52J8Ad904xJdV+wJ0Po+2R6F1NBoIHflVUYom
BQOOnIGJ2MbCruvKuWMocctkuLrE9MffunI4ZlY4U681u+QXAhG58EateAefp/XW
MaDS85RfFZR3ZCm69mZ1j4NtLtEbfqCji/Y227FzZEdZdGhVsBV/6ngDC+uJcoQP
Pn2kKKjQkvoBuG0PkkGY7zCDvSiAaMF4b8D3QvcYHBiUbs7spJBmAF67gDBlcO9M
KZ94PD1q+qqp6LWaBybKrYB+IjkE2Sjl2ORZfohQbSinER97OIKAu8QNr1cOwERS
fCSI8C5cV0QkCxXUmf2CobaudIL9L0U6vol1BjMO3Be8cq4yVbF60lf4er5Z662a
sbM7HWe0XokW5uH1mv7usSR0s77rdS8x+w0l/oPc7ufwbDHj2T0M423CSdKkEnF/
H0fX5gb//6uK7idTpMIWoO0vuhkrmXOuwMSVm8JfzFfqHZEhph/JwBiQ2qxdQS8G
hmQPct10GPPvVodb3qIeM9mXbccng0bYoPwcomaPda5Ppaa5cuvsB3DJscZ2exMl
OdPNkgtuGTzHJBz7SgZraGX9ucvvPlTebA2T9cX8IX79WkCS5UF5wSTXG1uIaIAm
OAfKkqv4Ndy+ErOJCEKGxqNNGrrTTbFvR4xRcfZQCGR74wTbDWq0uq4KMkSlXoxV
i8DPyemUmxBs1UQUnlUend/3g352NdviieQxTs5zedg4ZbtCcxu5nF1aqDHB13/Z
gVRALCWKtZMCScNr+ti/ULorGDtIkVOQL6a4qdfbLSdLdZppYxdzKyboVEdllbAq
8Pdcz7EYpVzeuFhset64hGpzvgBIzXmahVgVAzJFhPZ9UCdf6BsjvJ2l1UqQRuxT
6ZcVo8qSlwK6T0ZS/dePm5o0OLrxtfSLK6xPITAoW6LCmaEvXjCv2UWXzREFYzYn
IjWSQIyZ2nEzi6K30Wp/v7uR3NepCFzJ9Yy0IWUSwgg6MoTYVnfecHPAL6YdFQI3
ZsybKI/v8qfzBlVHhTE8hQnfHU9vJgi+BOFxp4rg3iUzaTBJRJj7E5bwOeAxvN3m
B8yJpu8cWr72L35EVeb5aohJWllYv8ARIduynRxVLjrdiKIX+RXpfX3dAhJ9BgE1
ti0Tc2IZxBq+ZIve9xgxGk7lfYCNcKYCkQB6UCpddWGM774/i7IpMDKrRj/SO6El
UkEYwQtAarGS3cGwwoBou9jO94UiL3ZvKvPAuj2rNXp4f/mWaB4LXlEOPIUySp9Q
TsJUNmQ5Tylriq8o1wXc0qr7CghSeNeB4Nb7QDTmR/aeRZ+VTzC7fJ1/jYFMlFyA
1XEudf0VISEFPM68+En8ChDWGpqLBO2lwpt7eLCBylPdSNYjviiZKSSrBYHtrB8O
93l3TKXR5H1yD3gcGuHxOLgqakpF+PfAv95VDkNpFqywPB8HWvVPSsdoJDcu656h
OT4ksVk1bCnTXAL6hzqwr6NWuDG5w3upu5HThvP2Xed1iohdWkF5K54kRV7/Dfi8
gIOOIPXuZ73OoiAQ4SjUqNBbcSpSS+nPlF/KY7v2iXBllVi4MVC2IaM2T8SYJrbY
S380x15ZgLLexN1a37nuZrpplm3dTF3ObbCHDznAWg2I+jB6a9G/UFcPdl+bz9X6
TUWArdnSKqWrNgLyXcp/iP3U3ELiIg7nPle59nRuSvQ5GO7XhcKsCjc1KqO78FXn
YLI/uVAP7KGradDJc23gjrI3dFHcKtCzpUSeRYGeihJwDmXEC1EihnBfd9NbOoY4
JANgtFSEwK31t3kRYYz2IhHAVLp6nJ/7MU71cLUuJr16xoDFsO99fBD59xcE3ml+
egqlAAZmlCvfvMJkSI552CmmRd/C+EZhi8bmLeSyXDINBUls5mb/vgwE4tuWCztj
+R2AwRmUp7VDbG87cAFjEgnPUpWrIgsmGSghI1OanTWKRoDbBhZ3auhcpjwPWk5u
mr0Vv7ITYbn5tWKPjeBJ3bw6Y0u/SgXEQ2nkoKsTT4PpnqsNs5RGCTNPyGunUyjY
XJwZYrOTsSRHEsY+Cn7+s4co6zSGHPLA8LPqOagx+b5DudqNgT0jNVMySgpJkL8P
n+lf8RgaA7aZh/8s/S+WvEhUfCEDVS4GqUXkwPJwzcvFdba2VisauXfCiUUElOxd
dvBoyYemPECJze/PkZzESVEC4emhrS7rIkPJNfZGf0M5hb4iTsLy5Q02HY0KSqar
qqmlZEFeDG211bvNtSdYzqyMaZx9X8pScMnx7PFpqY68Aum/wz1z7F7mR5aL93qw
uLpsvE5hf0aPxsAKhYNi7DLmwrlhSY4KgTbfV5rlNhvFxRiabSBeN1ZANGgl1aA0
cxiZWAexCEgXNjUgmHchNNRZgJhiAjVLuGd2QlVI25GqkAfmzVQMxcWYB1BUZ8k3
fHzSPpWypgEQJqxlWaT1vVytRG/Yr40QAKYacPnQ6DTSpTUiQuprGVIcv1KLbxPA
OXezpKQLuBfwadpqfsFgZRupCa9AFdVRt+4fqKimH0K/3tJ1adff5OAbdISYtjvE
wZCnXlaSISWGLATsgasbs5f7+I98K6GWLXNtD7fGXOwLhpRZBcBSbPuY54FkACyd
55J6dAgV6lsDKgJsE4yOvXz9qDQrqqQW/KCe6YGNWGpbsDRtmtSpU5YmhYEhoBE/
Dx9zYKjTcusauVj+AKJC09V/jtVnKGfKS+RHvne8eFsnA+3eyvPGBTULCbki7Tlk
BWdhpLuGQYEsd9BqazFLP+UssrDveI1FNw41lTHf6k0ycmSnOsBj0Q0/oz3RpU0H
nutO3NRwBxfh/ln8nLxCCBLcI22Ua+srVKx19OJzxHONWB/mOmpvEdqgQM6q4IPA
FnAYltEyZ+6kscmzpnC6k7a+p6F8G25SbqnoRXzYbK7JwuBEBpxpR2Wa8oUA8YOd
Qh9YxhNYw0p0aav2v66qLc4pUO1oaZB3h87gQfxtzM1XJ4BUFesYsqQWOsBF32aq
U3rnO8sTuBbfFbtutTLJRs7VRVw8kx5MMi7pS4K11TI0bpXgQI4CtDWP5BTiaEAL
ZV7sk+/M0tkXDa0Z96oq5QjHNYNZ4DGYi/sbM452knY5OJ7l6fYP36YT+ci7SXeH
wMgugH6NXDWsdasjBYCen/WPuRoUBPNZEXDYBLhcAaMj8/o6m6aJ7/BbEP3ar9qQ
rp25KlnwPtdqomWc3Vk+TIH05wTLyTqtxFtx4ZtSA6diZPstM4lGIX9+GMqm9UpH
yBwLnOBZP9FISrOM6UvaSxLwGGBPzXFjOYPLYCMZpOZiT7b0CjOE3c4eTxiIG5ru
k6jNyG0t6YzD6AYELLkucZSm2/6xx5j73p86W/Wq72/KktrdrDvEUU1vL6o8M+4A
hy4BU8MeCjaBW7p14Z5uoFDvk54UFm8Y9FNlQObbV0qoHmPppWiXc5FPNH1pzh+B
C3EeW2DASui3vdyCtuOrlSkkcHneBQSUQBUxM48Hd81ghoTkSHcOaPh1c8l9+utx
24aE/jOjvs1NFi8yry18ivJ/si9dSpIBOvoUH0yUdBK9E6wtYVR939Ki6AQ7YdSb
ReSmDsW2XkU4eoHa4t03wgfAFwRW9dEyD77tQ2nlHS2O7TEEFCnEnsMpXlw+zRz1
Qjd670npD1qsw3MFkywZwRt4JjYcsXT9LtHOxX+3A3Y/RR/Ies+ca517Am9S0ilz
VhDN/RDGO6Gl3sKcqzTmby+4BTpiYlw660iGekfwRBkNdem1+jBgoRDRv/nGAvZ+
Blfa3AEPXo592aGfs/nwX+puOFpFv/gZteMD2krUGOF13gDgG3j96lX5ePqO0mj8
3ueMy7wup+QEBhIcmfoOWZmMrN6rwvfvfkBv6olw8ImDMiY+P6g698KIZl07lzjA
Sv2/gRkWO2gqLS0dQ+YwS0FJPgQ4JTIP+im0K/VIpvJVFwUheM/QEGrno9ev7un2
eWNBSZAMNw5j3PKxNR6KfNzLiEKmQiAfQlguhrtsjwTAUEsVfgyUgwdJzGfXFtky
9Ezgei+FV/YX/9Q+5knObV9OAvXN3Y+6LLUN2xlP/zOSNVBQfLsxFn93AvvBvoRs
D13uIoBlO3EkNQQu1oMWbBm1shQ6+IfitQMazEREuzpoqUdQ3Pkw7NtnFQozNXUP
UnO7IyU3rU7ICcxC9OkZivmpHx14RWptmdt/nUQBM6RxHQIeDSu1jUHP0jxn8K49
xqFFL4Q2IZHhsyTLEX8MqJs/uc8bbQaiAmnuXXEqv+26P2M2i6HC3WayeRjV82K6
Vzn0PQEjAgS1WVST/veP9ghWXkFsvS2ESwudVS4L4N1b2zNpCCO6FLw/PyFOoaAH
LVpKOSjQEh4WWoiSO8ipUnUfCKoNu5F0qmsCV9+aM1H9MN5wR0MVudKx3faaGbct
BF9Aq24FWY++wsfOJKdolDH7o0nGLBYbLZLIwVRXjuD5Yq22aQaZUqx76t7KAYxG
lE0ZynOVCF4/rNCqfeAaFgD0/DB0bbQLKSNTLwVsnSCoKQDmKp3hVTO8n58vgvXp
TD1IVCUmG9OjlIRu7p5sc8y6VmjK1+TJv8Jq3UIwgrpN0/EDdSk1H9te5rN9uWbC
enQdAh1psgGji65nrJN109s5CPRfXuPyj3JaSd/4MbAxN5NxFzzuVkzSi6vdeImF
01hNZmQ2XQTfAovbX9Su8gLmt+a9m0P/xUXoh7tAmQgqPLMEsPImhv/RZFjsbSFU
Lc8yC1Xo38IdSU+m9kxPne6hc6wiHO91RMcih9Wjp17CGmfH6FwYuPpBq4ZC6XyZ
hKLOf8wVZ17NvDEzgiRz6wvrW+3vbAvL9LZWORzHrSUAs9PKYJRS/BUvjmFkQ2rJ
HtPyPku79zCBuuNZxZ12hDGMCYe9BrWjv8Vv4F7j/AgXtGP6dXP+SoQ5/Alg3sew
L9lBXqLN3uKf9XPyjXol185qn4vpeIXIIHwASGghZbSY5g4JHmcynE94AXFukpAm
ETSFKXkUN6UcMlhl1V35xJRGZrZtNopbk2B2E5IHRV4shD48/9b4A97nJ/wjppCP
D34u1KU7QxpNC9v1pGzbhcu3H2tNSRJuj6AJdL3Mxdeb7kCbEsyjfw5H/yK04cC/
zzrgtu2R4PZ07iyw825EEMa+G7R64HRJtZsx/pGN2h71gMzezw/o9FV7hdTXyT7O
3G8cRkycgH2bwqhtmoU3wFOaQwxDxGHfTlc8s6pvW5U7ry5DepdJAR+7FqPFQ2m3
bsA42Epy01kcSqbMLWgJsw9f77r2IIpxqSNkhBs6A6yOjK4oJLwx30syTWa8kx4O
bPrbh3nV0j/ABcF1kNxn2K6aMv8rGWf24PuoECAzpVmr8XNcDXHBbNTrcUBCnM11
2y6Tg7GIAjOayhWmwO/tsgh3nXTC9W1QKD5+93snG5tQCNp8LuDLJkEiWhK/izpN
8mLl8F5JNr92/uAYbY5ipjKjs9nOfWzqOnB57N25x9H25hV6GQ7soI906FkuwNca
bUJLGD6XykifsOfgjw+oGOurA6s6irJWjIKNm1xmMSdJcc9d/+eW3baNEXrCMsy7
OnRi2h7ZunM9hqSg49kfq8SWhLtXOCaHwh9ZO1IwHHi7gm97qTBHKb98s8wqPgjw
s/A7CHf+aOritMXcFtoogASR/osDF4XJ4TTlV9qXJYt+CUGm0K4VMz9F8FBGCNul
1j5U0NdKA1vDzg9i7UqX03lvArkprmjftTTmZLlQIbNZxN/0AYJ9wLHMlPgp6Z2+
yzVYMiV6g4ErzwPTZycBJWFZwuTdL2OzEJbbcP4c2np54zVpP5NZjfC8Qwk4gVFt
AZ39J4N+JG6UOtMzsYrvbCqrK0nRcHPZgHlV0ewMZF8m7Yn+Fo1LnO6wQ8dXZtv1
chVT1VizzXNztyfa03K3Y9korntDdDW3YhRxls/EmVX7halfwGpBi+cX+MUQ9dXb
huvm1rxaiJhXnZDySJJ6dIz+9B1SNUc3OGk6tFW6iTX9BXce99YYL1uq5NDcaOUM
qElBF2oApmqi9wzWNLviZ2xo+OuezFeyZ6bigFdLJu1A3W6jV+rx7BzSD9Gb2oWo
UI/u2Y9QCkn+45i6WjxRjAesaZhrswMbIbuEyqsYQZMEv8a/gtU4VSsokdGzZYuM
PlWque+Jz4nT3eH7/R1Bs85Neq5WevW9Cvkcr52OpBfR1sIcXp9XPDwPbj0avan1
4JmCwGtGu/vnz6n8oZXvlHF0KJ+NnyTtjMEhBMVjxGtPVNp4vnKcpS1DR9EgSyzV
AcqvWj3UcuEEtmR9VCgDyCfWpnr5DUChaN/b/+9pLccfFMQPSAm5KyIcfiE4Hmds
IWqSn7e6yyW87iMbdN2bkon3jPH0v+pvpnKO1aXiF5tS1wQ1ROfUgnaf1NB9S7qs
2Q4peFNrWHzNlu0p6MBsgVgHLT7ImzwMqhVfDx1WlnOCdmh7Yq3L+P4v9FHrRFR6
alol9PhRUrsgssP6ro2uuQA8a6AbFri0FxBfjIIA47fm1wNRLB8uLMWgf0xaq4Uk
syTy1RpcC9oKdQd+UccYy3G/jsc7pGQSnOQkjvV3egPdXjMZ3jk3Woufv9XBmIUh
GZ2U/tx63UvE45sD+p0Ughr7+iPENPbLpWsAa+1jQmg7nwK1NXcQBhSQgYCo+wXx
1wKNfNwzZmaqxXEBkMOkkYgEXNvdRAbe/IJVZwxxP/Wnpmf8sjL6hnMXf8r9rBqy
Z99Bw2hXBt48IQD31/0kBukwPXAmSaQXr9KaPk4+S+sNuDupNaeybK2zVCJT+fLL
TwQwn4jNCN0UO3MXiJB5JRMyOzj1eMl11ptodeqvC09c2tmaB/pnVxb7yITKUX+c
Ojhv9DxmqoAox6aNIM4R5bbUjRPcleNK01NqXCPUrHvMWqA8w7BMBa+PNK+NIFt0
s9zT6emyskPHWxqTTAl9FLxP/gT3hn5EQxY+pc5N1QDw0R/FvnPk0jdar94QgeUA
GcNY8AlUW2HRoli/B/oQVx4S28yQWBT4d1ytbPo8fT1hkdpPrlojZ4rqcN7ittWT
8oTdRlLA/wXN26LA1ElFBIeACZpdp7SomLsl3lrMUQI23n1JIlMW5xXA0jiuSsZg
644a1FhuCW/peurkYevfiJ32keBqKDNk5Y9SAtSweHVzadB60Fr7vhHc+BFu4fOH
01DPcd6DTf1yIERhzA5Ty488/w5VAXXEdO7MPp60ZjeDgt9eNf5IkwlrrHJulyOQ
wz50iKx9Pm+VtmIHg/YMC5A5VinVFu5nzlM9G1xqntq6Xb3hU4nrWs4t/OZH0JSL
dsakS9tVPudUZK6jj0QPW0icOnyiDmvRHuP64dCz0kPjf13vZ3gG7xOqXLyfDqP5
0OGbaliYH8O53Y/+i6S3A7Cs0Lwze0ptbxokceo8G1PiUEVTIRaJoFUOwIcqJXHF
ixwsl+VQrfghu676t+XsTC15zfMIWl93IAlK63fZKHYSBvu6udG8R9DCMh8cRIIw
vddBd0Ud4iM4IPdldBbm6BogZjEoQ8gjoCq8lbXCjhYKqy1etKpPPAr8Fd7HKbzJ
Sjg7RlPokog1gdsrUsDgKmmECYCRBe2y7SVwXe90E8QyYG3o1REH3XQynePG42h5
FGTV5HyhQvjuk89zvk9Kn3uk3gJWW3VwpfpnXWtgPAQYB4P1vvYM+UPubXQ+cbTI
2kG+6mFoFtfqOrcKm3M6x+M57SMSbbu9j5pDrNJKKD5JELDVjHcL1cBbRWPDw0lZ
aYblnIFC9LuRgF1p99BTzsTG44J7obyG2m54hZ6nROLj13H5xULTaTSAH47XbwvK
jm9jpQo08UoqStx5bvmt2olm8AKHscD5m3jEltV4M+ALTgi/tR5z1QQX4WWBN64I
SULzZ0mKvL4hZdsP+hvQASJPjjCYGnmxR4udel2UxKrOUxt5qjvFim0/eDYYzcmu
otcIHyqwTCviN/zp5wTE4NHM4diTTZMSJkM8ja9kYQip8AV11aP58fYZlOUp2tnM
z5ekSmbHIvgc6n7iezi+AX/qjpzWpXz1zEjF2YjcxllmMbdQojip7rwP9DF01Tg0
0sG9RoUcMgZ5GShClmNNRyCXFU60rMWmF+QbJ20gfUtg4B3HXaWqi0EdjBpUzFjq
xJzC6tw5ZZ0CmUy9EKn7REQYwaY6nTpKQ/FXCW84Pm4JIyXIiUByvDOC+cqfnNR6
mwzhoNBRJrNUZK+vBAdpKsz73ufdM/rVn/i9kUlWdg0lqHtze5P+7kaJI4VImBiX
IHmtPtwUMVvKOr68g30AMkpjWdhsa/ROmxHcX0foqtyW/xhbIdBtjpQDrmHRmnTA
fl5uy5FikcCnnFyCQdTrTLnxZbZhNtw1QjOm+1PQLDmJ25bSC0528ObwZ1apQRBl
7OIeZ/UxOw3MVQHvWq0aRnBTFINv8rsvBQf5ZqJTqXZpFLrThMYn/q957XwwoMzc
H/Afr/dIoDjsu0VF06/V0MdHdzADNhYcB2l+HZaPMALvQRcPnbtfwBHui4bdeGeL
mhfKx5Be4JmMKaPZMuwgtrdRDuTcWLUdhA7VPyA0laVDFZASxiaDTh5Ub5zQqIwK
udteqV8fXkJumFcZaRGq3pckhXsnUbtGKRg4LjGtwVvgS1VG/j388ag7jgvWGTmX
LLR1uU7/trSnZkJh2/KXLinQKEtAGwk4iMBiqUNPXq1BBtaC6mqqPDRvaVvb8p3u
vmiIkAzIR3XYkXsecC1SpaH599rI4IolH8OjRqaIEH17GxBMJDS9HhoicRZF9/8L
0A/6E2tbPKa+fWgPz5tYEOq5KsxEZwMomnT1Zfokz/ur048HY1krZ5kxvl9S/Amg
IDmIJVVCetzdRIjOsBME1GGoYLEU46UOVbgV4456jCM1f0mrmKxGFBVcL2/1g60M
EbfWzmlxUbwUdMX9JpE2w6vVvaWEkzYcN/Eq4IUKoCZfRJqxDeF5EYc/RYBOlXEq
ZvLxJFwZiECrjo5PTUlAB3tOraKV2LVT4grlQvWWk9YVN5t4lHBVmqe5slhcBHkB
DKokcQdidjpYzzTpoV1w2N6vK8dOMqoK19yfMu91Eu32w23HiQGzyNiLFkxcx3Jg
ji8Tv63SJScCtz/yt8egFX7yqxRi/aBO59fy8A63djB2sxbbXs1MIejqSfZvXt/b
IMZASiT34sTYIurQggvCvJTLU5MK2utEPcH/NBJCNpFnjxvThSZS16QRFGbm+v3e
a0V2QEDVSzcj1FYTfipqHwaae6yKxkyA0mEaVEQ2GOZxE/SF93o8ykMP7ROZXzHu
LjCjYz2gwizaM5/nlT8tPaGPaKnqnJ67gWi6WSCUsVovDzi0zd2OUDazeQn0BaFK
FYyJJ6/E+QN+YLc9JVaVlhGLJHeBtFiz5fqWoxAr1+S6U9vAxnsZyF4sfO0PA5eD
FiBt/2YsG7rBWtwW6LQqbnLu/Jmzugbb78elSrxgR2IYRVgiuPZs89uodmy4x4MT
1+vGnDmcpKRJy6rz+O2hbnNwSiLUEOfX1OqSJiJ6nNlIZ5PZO80NMgtiGMNRvQfi
kOyEF7UKVYyO9UnOJVxhFpbqoSRS4b9qVeKuqjkpzp1hwNZV9iJopwJshrb5odDo
e2kVqSceuSC3gYK85Z3NGkrl9CNFtJc8HjkHonaIXo9oXXLwHR6PV8q3l9qkpJ0P
z9J7UZcLSDPXKF8KCbqWl9GLX71TiRtZsHTKbDbdsUo0rs/Oc1WsTo+UxEj+SXr5
pCp98OIPZhg7DaZZLjeD8U06c1WTl2bBdW02dQFq6w8lEIJLO0/ZcJ3au0iAjmN5
4H4awOhTYRRfbvNDUw2rP2ZLPnayKQdgWEnmdod25VDmuZzvFQ/f2KS3DeuCB2v7
BgC4uVwDNxeZ516d2qGdUJmSoQ4KIA+llxeMfdhKN9pRUwR5nZ0jPhvFF9f7E7RI
WiStTELiICZmG4/siKzY6MCeM5taz1m/XvAXiDwkveokDKLMTZ75UgYoavam+Y8Q
sKJX0rdiWTgg8yt/IRvliOBs6K3k1yUdWfgyqKot83fFgvMwOfwJ+88IuNf7Un5+
aU4f0PhufTVg4i4cn/NykmDfV7KRmXSWoAPMQ4OztfaJ9VcuqIRqwoOv4SVbb/t+
6mH4lnMJZAxt/5c45fiMbDzt+1KA8B3fIDJt+PDw7b70utm7VOX0rTV1e+1I0Sry
BtotMpKbE/UdChbPyUllHdXqaDYbQjkam9AOw3oYDu9iSO3GjFmToJjCt7iRtlwa
8e9aNEi4PxMqI3awC2HpZEGGIp/3cAbsunf41Q3qit3ZyPj53en11c5/KPQ3ENmv
T29zdWHJlk/ZuS+JOQln/AACUfVq6kwo1xFM1a9EZzTId+NB1v/wX9GXtQJFGmnL
ChcOPGAuulIbKyNxJK55TleE9tO83ewArVRgbaoMSJvmTajYboP5GVTmnzz6866z
iF/DBnaPz7+pDZi47cbgKB+V55Sjy62mb0kcB0SnUHre9dPeq0qTS3jJFV5RtyJv
OAvfXKZGz0eGz95A6xNthPdfhajQNCvjDd0wFSMNovUe7UhQnOtQPGRX0j8V0VWK
fu5nfCMbrnUIsKSCzO1lM/PTOldhEznRCY6jdO5oQvZQZmaazk+jaGT/hB90fPSO
go+6SknnRg54QyPVBq1NeHsbsvBW8f8iHaRmMECjmN1j6o7NjGVhDR8z7W0gcvSt
lgIorYsxKDWM5YEIRl7QjuXJDhyhUAUuaI3mUqSww/jyi0AGfrv9s7hWGA1PPtSw
Q/g9Op+163YFleMlU7dTc7bXasXKyagcaXecUNTN24tKAGQGEsir4tW5Z4z71miy
YdxDjH5Maq/yzWsY7ian+Xk1VE+LRq9kPgIA9kQSXnHZ9mb9zr0Iay/4VmbSWVzL
utieP81+L5AMvS6YeAD7loc/+Bm3IazlPe7sZuM8DgHK3jb9r1X9ytvCkSNweVyk
+BVe5tFZ4WrWhLt0ZicBVrcXDN1/5kKaRhmul4S2vHixF6ErauYvSfTKurDuitRG
kmdvBHL8BEHq9Y5I4CyVCXCGYDcVxGUu+RnyQUruo15UUGtX4R/wLRro60UwhWeU
Y5eGTU2JguJm0yPV+aSu+SpbzFVz7iW9SuSLmFjKRck/RDmZbQqP4DwsnPO/dYGl
TR0NyNTwOshMo4hBuTOV2LXRhzFVP4n4E401s3GZGp9KNkU73kLma1P0+rJ1BxTL
aZJZm3EtnK9nytI75MH2l6B1SCorFstqEaWUKIXHueDMDOm5PzzAig6ByE5urhV8
pdcRLDFR7hnW+t/pfyoW9HZj9Z2wZnPXFi4Mexh5xSdyNlj0TBwnmW3iRpwn53W+
jscMKEzBdrbDP/axG4JPluKfyqeB8fjiK9xCCEmACE8DDZvSMvwgobLNmmJEOsF3
8Lq16CZlXxdb5EmjD9J4kxgu/CAzBr5UTFobBrEpRe+QstIkeZm/pHiqhbEFKs1H
FrE4+kftnvCWbsudw6EoWiCRgiqv7EEBotiY0Rb2PxP1eyHd2FyN1/VRc1RmQUhi
a+Upz2bn9Ca1/KSppTuo+FqmJ12UUEplHWCbFM0IEfwP0w43yN2VaFZmNGUBg+Wb
sGzGr6Q4MUQT4k5VKMNbZA3U3lg2NKA4jx5BbNk7HfqroslBsrt5uz453wvRaREI
VBjAx0IlKQBQ/sH2u2lIYRGxwQbJ2YWwAiOToHmQg1v7eLsV45SL1lGWG2FL5qmP
8qp16UHvhhUsn8Snv1Mh6+IyievoaAGvoKAz2lIoWTh1o5yWwFy9NzEcRDR7uKHy
/6dy5sauKEShw9MKi8M2mo7BoxsqV/qmHeeRgsU46BMz1KNSJfiwKZMQWFyU+ZVM
UUjL92tOqpWqBEfZIE5zI122AOZ/26rShVH7dmr4qpCLp4FdHTF0tgtgNVm6TOEq
O/gQeVxQQgY1uT5WjX4p6BcjEtR1PXe0Da2qO2I/JMaOHm9v8XwfgMZeQ8oWKeJx
uWJjP84JOCjtEFm+W54+4gnoY8H1kkNNy6gvFtCJVNg5RfBepIbjX4nnGt0SFA95
zafl+lHUuUdXSR8IJo6ST/IlY8ibTjKj9ObHKVNjDlxoiOO5QmN7ErwOFlvf9qMO
g7XGTuoNiQQcoEMJ+CrN4uEFiB9jUApINPOYckRC7JLrtFB9kS44y76nNWnXSOdH
akXfRm10EbAUO9a+EGd9febEwg2wR5cObQ3K1+hNhKWqxe70Ws48eJ5gLCiPTDJz
01Z6Fmx1zN4sKEC+rh9/PYX8243fqrZS9t+AYVNojnVbJgGHHiJ/8Q5Nyuj4ClHq
rJaKB1uRAOnHjLbFATA6+wXszDV1V5U6dEAofVRpWgB4ZFLE4vRI1IqOKJOkeY3R
r3qH9bmwFlCXGHh+Bx8x2QrzQ+vkIz6Ie77eXMdS/hRQmPwvaVcCzmV3k8ZIH9Ln
gsu+lDn7QrvGtJPikg2Pjix+El8K6mlxRuInvrLl7qu5XRQEkkmW1rbaoWscJByP
08WwKl4m2MESa6oB3MYq/DEnlov+95267F1Dd2KEZiw4oOZQ4KaoW6i+Ta6sO0Il
woWsxN0Img7IOa1S0+tcIN/TLU5fVCQ0xBQ/kZn+2Rggd9zyihzTfwjzrRMP2F6x
16TuteF7qsB3QvIW4eHTG3DvMQjiyIatDpyZvubA5hV4JICaeXhLGYnSlOGoaYYr
kQL/XN0N2Gz8z57JPkcUS7Pj+XdjESkeQDnIoxXkdyaARLpZg+buZ+hGKAUTpbOR
MCUNySToJTAYi/16u5X7F9DDWNPJa2B7ppw9OtLlGa/E4eh2PeePFDP+rVfFhRx5
mOjenClV3cadF6GdCFwWbhvHGLQMcHhl+8NpnVmgjs8Te7PCbpkjBFDxZTAKNFrS
QS0gBcgsydSGpSPdGasSVJRzEIjZmlkj7GWSBzPPtE/0H6Yiaf6+cM/WZTK8vbNC
PeGJFLTdqxludU7Cq8XDAOqVYyn4vo0xcVY1JUDjUHJ59rvVC+imFjzFdWhG54pj
uKn6Hn8C5q6usvGQLnOHPDZ7z5atTmnG9OleqHju5gUDhh3fIKE4n4zN97xknPZu
p/n2Y0SLsAd7lPnufHoIAF4Ms1iG0t3TBCWhoWKNZWs+qCJe4D3uMIff5cu9o6g6
oZNIFN/kNm7+cyiNB9bPjHZNzLA4vxsIpXrciTETHfl5tAcmmeCDKnV1m3/Otpxt
rNNztPUFCkaZzJN8J4KFoEvRHBcuO5joY+dTBa9Wn7CEycRI6cHnn7O374R9AG17
KVndnLPtGbZsfy0wcMUxVF+QYiwqD+oipkrDfX4j89QJL9BQ+sP/umpdAg3s937f
CJifXUZYONOf/QI2ePX2M5oT8kINijwGhXVplF6CxnRRVNq9KgQdK1LWQzp0Qf6R
U0vhf4bBJi1azNX4rw8q9saJibmBdzGmXz+l8ji5iv1ub9lxQ4Tswo0wisbMs5yi
ZvXAeew+ft5wmcv6GIksgcSIr87LOaUMN0iB9yylJDsRShcLkNqtfWPcNj1HOZqB
dhwOpZnfKVrQ77UU4hGV518ILqizz2S2xr0ddGHaTreGCgQvvIzkosWIpDzUrzkl
o9E/RjrLief3F5f+wX9h4iCjX9D3HV4Xs6iFoATyxa8OZYddgmD5fHnzMrGXtGnP
Purtx5N8HinXMknOFAvOdoEfdEIwR2iGOZ2l78Gd/xYOuLnndwlPVsgXAuwfZ+zu
5Y1vhqM8FUjfuOR+JpL9KQMMZ1s0zp8YZtLEhOaSFPuSrYjTQM26GxHTrGNv6aea
lidtmN2W7PIyuL4NwPIKZS1YWay7HNP0DrRUTLcaFaasylQDorCq40osk3veLueo
c1sfxZRq2d4diaxjvZFbQoZqSu2dbKMD3DLp60BT/qoVsimojHt4vvM/FwvnqjY8
U3TMJvtkGcUrZPfuElohb5nE+8Z2M/a7kj7TzZvdVWazQ+I/we8z4vC7i4wXuNSv
/YRGzfyMCEbdW3icoCX0bgU2HU0wvNk2KS+Xfv7rewOToYjGEIvG48JB2i5P9ERC
ftorJaN9BEr3agLGYpPNFyWtFN5p27SvAMhKfV3oL+eD0AO49XDqhvyqDtbfMRQ5
sluZzruVbNR+YwDDf2xo+Gof9j7Q3oGQznZVTv00V0vFFDLcvNRApBLUXxEAS+UG
AMYOuy/KkhwAN+Ny3oFCDGisdu9CSLaM1PsVa1OsdPOwFRvAeJ73hVblV4WcX5xP
/pjsloIQHHHoHO7cVPikbthkoRNr35tk9XLe4KU0oZ8b7r1lR/6c4pqW+hL6VqPW
Lh76jvwoGB0S7IoXSCBeeMmq9J80nlb+38YPIHi2DHfvQYRbd1jgzyfwvId7HBlr
LyWzpcM9g+xQnpHl64DwM3fSXAjhBsA06dowQu2/mYtHbJwskb7NWC5l05llSNX7
3woTzw490Ac6IlQqUyWqYJKWFer9NPakpJQDYayT70xmyVQQx9xGdhw7RiNkwP/r
PcLkJwU/2NJiMnC3nETo8n89eq9kXWGCpU6Cdn/BiBuG8hrLde037DIsY2qU2YJP
FqlhrkxJ4r/XGHOJcsTGygaXu+No3tcTB4EySDKuLdIcW6U4a6Osg4N9+308z95Y
VjGnFRZOsgUsuUK6uUDE3LxdUlA+O/gkLzfhwHrkQBWdAqn7XOicyChE1LKkKTZ5
hgGbqGVF1ZKb/XgoBJf6PuFqKSh6kPhFeZjRrixQcLnzVjAMDCHCoXyBSxxWTz/3
ELWXS/S3GTS0DcxziIDowfjqb9EIgIE4wSYJ5s0SzZf4hK5GL1ZFD+2udKp94tTf
C0ySpA902/eDsMhTbrABANiG/iLXyU8rQdSKGM7/cpphbWEQ0DqSywLL4cCKps1M
dWuJzMAsisvrFTRAumyy8hvTTJe6U2MDF4HdR5+poO3FqvouNrLZmBFkcSyzJD0L
9YCAkp3YHOUqpA1wT3rwtuitTYiWz10jkQLucEjh44dwW6AUjVJeCogPCC13rnDP
nzs285M1NBIGvOQQJAvyOq4z1c4vgK8vnf7RXtY0H/MzcJkEwXTJtwN0w1+dhuOo
jWHM8e29rC/7o1ofhHajFrBVW5+GJFx7k4E6RaCmqMQA5h9qh6L6xFP61VuXp/ZY
ZCSd6P/5Zyl2wnZUwu0riBsTH+NHT21h1mngXYx6s/KBEgFK7k6F+KAyYJMvj+Lx
2eWBfc18OGN6sqg6jzo7joJE07kqW3n4H3nfKaHxn9DkRXmOSAwp/Jc4WXELgyBl
PnkOpvwEAWhBDKHKxWh4h6mZuyTCSvpgXbIbwHaT1G1sGOle80l0ZSdRTQZGBKkI
XBTgSN/iTQo8zVn5rPQCKQmKWbFCR4c5bWw6puMwdDXJFZvARmkv0tkD3LV7B3XG
go3IgewA02Fw2wyl4P760g7pK454SMpzghGd5UklmpeukLi+fiXs5XjI5+ZbkFh2
MDQyJH/s+Q6WYn3zTrEp0kEnJpU8VoSDoh2N6F3dDjGZzLtCtFTGz16a0F4N/vRl
uq48jW/nOWD9cuca3pZN8wU8uQHrIo/vR26slYl0wTSZ7sGuTEC2gbFt3dEPnwrP
ADyvWx7lDKAXDPMS40iYiGGlkCOX1Vqhv66tsq1a/gDwKR+OIMVH9EFYdBE10pzl
lJvq/H3cghYROzyiQTL2N/r6t06LkPdbJDlP35FdIPp64wsbsaeEqtjHdUKsZ3tI
C3/QWJ/v0Y+0RojT/fRjdd9cBfw+cn7L2L8LejRYDVrXM7tM5llYXiDZLQ30ClaX
6FZohF4u7YPD9NofDppju2ZqUfBshBlVOHAvOzeQwYqpROwaGE6o+idWw/+N5+uO
KDRwZXA6kfRRrSLWlaF5nF/pMMOXprSK47f+u+ErRULOvQdqx79DJyVavepJTH1a
T5eoINmObbErNvZNulHvqPckSwMm96aV7eSr73489paTXh2zsx1hErAEU2nAJYVH
+ge8GLuAYJx4JNPXHogDR3Tm6kinU+mTSxvaW86EqTOlE1dWP0TgxF1pH+fAuIo4
77g33+cHKn+QsqUmJyykP1fmLY0JIp32eYdf3oSgvcgIlSmcHbspm/f1ap9JOhaw
xXVcznEqeWgK0fC8eR5OoJt7S995LT+prMX8NYIMimfss9AtMUeCC8+ZjKdb1rvv
J6y7fBpYz/wpDb794KIMewbQcFsg8XcFelVxCSp9VO1C64n6mXoRhODv65XrGVT4
v3D6i2fGR6USWO2fQeyBGCbGFqNNENSN1A3OBtGB0w2c9VEOxNPRep6i7YkAJoA3
tY5yuGRF7Zf6BPZHw0f/lgStc2N1PhOIJhI1uBL+TY+Ls8aXxmVH7s+NJfrqsp+b
19E6OZS00EEwYMeF8ccBUxS0y28eyv+sURwna5Ywfl+dhEuPQfQ0EbD5b11oeNvd
DTe2JV8ckSKFlhog7I+RqkBh6V6566o6Q53lAKxf2V4a7x/5sCdu4CgHW5cYyx04
gSXUuQtgexWbPhwJunnC7xgkR/THhHI94utUJ0leC+SQXnZvCUkjtWUN62yd0iDA
Ab8D0p3RPv2qhv9olsJvunzVkAqK/bkDIexglHp+CaAJmTpXX0gECePCZn4ImobV
rEUPzRumi2/xSjmWsMN7MOksv6EieHWayVylAAx4mXK/as1K95qMUGJkzJx/bkbT
SqQCLAakv0dX84mkHXU8hh594Pa2xYFZm42Hqr3JMOL3QZg6APWaFR63bWzvzcQZ
TbPjOGRwbYwbgtym0/vngSpYtId+icNdclOvjPdHkokKiJA00AkbYTd+MfOx8iX0
SYZzzA/T0nxMrf6q/IiMt/LoP+Jz32PbqSVms+teltuRCxlGBuI7BV4GWTpliBNr
Q0LGTtg6vyUCQxwdZpl9v6lUuq/0trlJ42IZSb1k+zHFrVg1H0QedPMJIu+VUp5F
niVEm9+byblQaO+iTzDObSw0wm/q4orKq88lzsIcY3v8i10cqHdcxtWU4zJN/yc5
STVQu9VnxHlgvYOTbATMKWgEtRNFW3xyNhws0cmxSD9pA9arGrbnb0S1aZJHYOCg
KYGkYXrxCCbMcNCM7ch+bGd60vqJNJFLJG6RONZdx0ON0khl1RTpUneCYc1byfi2
DmUAQjNAQM7teyv5LIEzO1f1sw+CxzWKNo9sNJg6QU8fv7PVvMIm/8kwRvyOzmg+
GvXs0GTujxCPC7W4nVcgWMabnyKXJLjeAPe9cZq7NUzXxgfjNdG3Ot9c7Z9YAFf/
3uDUrLkWIw3vL2w7LEYAG5pW3dZbmPURqL3M6dia0qgFUDz7wjhtR1lnbg5D2eKz
hDeE5Q3N96DR6aLR0ot2YG1L2vsnPnTyKOF4UBu1llWAjqQI98NuKZNvsRRYdjVa
IJptKGzq9hhmVgVtlgMsvHhrp/i+9k0f3Yd6OcpE57sFon7JMWTHz1EKEWWh4SKP
zWI1GrMeExgpbw1Oek7qu1bWZOr0Dhx/BY7dO0scKAasusDNEA/HI31O0Dr1QeqG
btMv0pF99mNp3IU2nnAHdGghsggHET4PWdWBeC6JOmKfG3d83mjUXLjE+Mux651d
ZR1l3pfo5SQksf+aYRFKE3LNhmeAesCgsDH9xrJhxYkhj0nb7wCNBgFdSPr4XGsZ
u/NUCL3dYKy+0afXrZ578bTXgJt8rfu5vvwIs4g++Adn9m8Su5+8CmIRdcv559W/
4LpUdXh1CcHLG7kq1u4vYfBUW7RewQTeKtnygfZGH+ZUmQIaqX1XwTq517rC1iTe
Q/L/43VwUAAi65J4Naamqy5zTTMeLWD6jrr0IVHy+AbO5FaP8AUOES3vXjnNxUX6
E922BdqqOWiMQTDvNNCCyBLVnYfmgpez0jME85C42wPeDBZELVV3iSFcqtxEXqhc
5vWXplk2yL7fpy1zqsx1C7hlyeb69HO3woVVYsCwzir7XjO7b+w/8lC5+i2fs9ce
Cz2IZxJGM/Dn5o2SbWpdPjPAhUVE2zUZDYq81piqskwjWFja3E7IkXfm90xAUgYt
0452IbY85aCVQquWIeJK8LsoO3f/Yi/ORb53KizAnRMXn8vK1wgYYXkjqxZQh1uR
d72cskjdgQXTgB42poq+qEpwDB3Wk6VsxpReKSNz25OG3WJjIVhSWE4FHGMFcVN7
XO4w/QFiNjZfbCm+szFYgI+qvhUsMtiaMZtP8zcZa5gDbUXVRLou/teQVqxK7XeJ
HK78wNCaEpOE7YMssgD9+qHrf6OWhQmcKoucMv0NZHWU/+vr03v/uXUfJSPsI3kc
YP1lRcNWhmxIGX0Pzh3/sXGwOofNuIiqRfYUzocuZzrvXhZ8GEfbEgB21E0YxVIh
Fu7Ef7hG/vro0k2A547r8daLloEpZielHtWTEcsgKqWfoI4ayFMEzaKVDvi67THu
E4o5bGXr4zfvz+5pFIUhVbFC+XGIAjI/4wn82nVix2o5IMCRcbIovb8y4PBtm5DZ
hj44TrAVfcnTeEPt1aSWTCZ9n8VB6CI931/7aTZAkiUepQF3YwOcXXY3aDMeKVzf
dNjj9z2nKE2lZ3MAS5jUxLDMRZrKhH+prrOwrifJumxurjHR81od67xSvHgL2rK+
VCf/8LQsryny/30R4nvC63gXDMAwgZgS+ZWOw7aBR93HsSU5ym0Fu5WC1vqkGxMH
mcxrvZZtoaPxtGrz0yCiae+rsW/xOdxmLDxlxGEKCG39o5lPfj9IxujJOtQPk0m+
KdI8cgxIklUu/FV/CJODchwid+6WFbfbRHBE5t5IRDjc0D/UehsQjB6iTSgzLZ3f
7a5AC65pJrZrEPBM0haPRuFOBBZmZTMl0FEbPEY/ptmMtm8+UyproDaiLxcF7ifT
Ith1cLGF2mbRgWV10tu4dK0t/Or6MAzyo0kBURaSf4ZjlUOB4lcMX82u715bh60i
zV61swCr1oXGd2Fk+36kEYzUM/fY9tJeUSV35nZF+CGOsB3Drfu79L4yzY1I3XcG
XwcekcKT7olAdGowIBBuvLL75uOh9wbwzrup5J2ob0xzePOt7QI2oQ8fluLB5eiq
h6VL/1IMSNKWybpDeEDgdM1DSW/ySoPZi6ZwdLSWx+5ICahdi6t7S+s5YfLR9S0V
nkMBjD0POt9wST0Xba1uqjUivsAPHP32i9vau6D+WLl3G2O7dB6lMm+mx+w6d+5Q
esVDMfLVsw7/sCkvFp0K4g5y3MsGGcTWusUH7hWfJgynlAyDe+lZ01ozkcNlSllb
LcRaBZYJgG/BwmLuDI2FYafR7BGz7QtDFp8JgM1ev7hsImNe9DgKGoa0HKV5o0TM
r48OGjvmfXyVQl54r8luA9AtyGh3X6HTGAEMYQ4DLe7aSKYy2X9SpzoWzlTJ4VS+
hxd7AzJEadW1xoxTKuf88w4rJeP1HY7RzOPRvokpf822VKKOkj+6LnEyHLHTkX5U
cagL/fMI4P/K/xNk4vYpWTMsvHSFNS/j+vrz3JVjJyxZjVwOQ7p8S8AyodMbMxFt
tHsUEyIrER3aqdT1HnWBsLvd3DJ1EpGRMoKPYJ3pkpCH43UxJMbxjQ1kBRkKnLLR
Y/TAgWwIwajkJag+p67I7ziChty5iZy5szayNNgpLPaXQ4oftLf+ZUmnEc8erKWp
BQp25N3y65lVxotUFz5OPUilhUtRM5/zCFqHwI4KfEbc+etCbvcMRvVm+KUad2Wj
jOxzfXGUb80tY7tJezkyLLgCq+Bq9U2B3dMDtH/pJGVnbKFe8rkO+RCxCLd5Sda5
upsn/QOWj8sx2bl0uYZYF/J95KbOaAkvwvuQo8plqpazdbxPHvP7KGXdkL+55zCi
Ggh93smTbL2TUPBa+ECqNmv72BPBek6Iq2OEbjiEW/2hxaqE1V69k+mg3UmitEzz
1Y1BronRxlygR/FQb7d2zosbG4MxmVMmZZPxGG2Qn1tled4wQcwe4aA3RRzEqvsW
r+canN+omQdhpqwzksz5aK1Fb6mnpLDof98T1waog7FGqs4SreDnDJX4GGg9MSGd
L+RlyPOAg5KFLBtJNzf6JWhAGQ57YnWtuQCFSQKnlWB0Ztyzg3ZSUhs+rVLpzx2J
w0qPjrzMBVYkPyp1vttmLrdWkDAta2brRXU6njjjILSvhHQmBUE2tCmFTbk64Rbx
744FR6aqdUxCrKLOB2XA7AQmbt7dULk8AgZxdSTLAVCTGDWUpUoRLW/TdIL1uFsv
WLZMbAyeIo/H8XkZxhFbyoNw2X689mmkoZ/rfBQfht+zwm5MIq5WVpMMUE/VjhB7
3M1lEtlaHhChSnKLzJ9vZInXTJvd/z/KOa5bjyzb74Nh8m5cwePELNH1wyDtTckF
rQpjHfp27TvJ1HzIz7fBwxHAGS1XruIc6FEtnzZ0wasusvFSCDcThhPX3f2bOAva
/6+yhJ5HbSjhWufhOUgGHU2WjtsdNM059NqRPRJACA85XTHKJY97+L+panc8uo8P
MYS0jjkIjjagcJRzUQmmemXktJH+c7iPRvLsL2LZkVqKwtEDllzVSogcTmZ7fq1V
KEKwFwZ7WvnlQivs/vaCn4VvCe4N0+EVphKPjn8lAz6R4uWO/9HIw/R4+jw7bw0F
QbGi+gzAdI3zlYhfqg0uX2D5ECa09JIsbnl2k+pF3RgvSYAu/jAzVuj/luNupX47
voGY70yTwm5IUGrpcqcs8pzHtzxCJ/yI+e2SQZG4UPlUm5adfXR/3+aJlLjTGpmz
YK4Jc5riHd1/QoOaNTsDqNtbErvlEQly01gcf/FxsbcK7cc/7qoWoAfvzCNIv5J4
e21Q/KBO2F4QBWya7IZWcGuF/27VMlBLSxIZtCOpp0XoNltBaguUvpJFL6BE8kXL
RLFwhUwuG4PGalNqL1bE04PSg9UPy89bW5IQ/IRHonYE/s61viI/0ORMBO0ptcvh
ysONddsMN+TpjU3fTKQAGIp/a5j2mpjfzF4wCQMynKAzj87vZm4PuJv9zVzbgelc
YoJHCQW1gMolUjtW8B/Yeb+ynD5yMxWYFn2i6VfCouOX7gnMsFh91bkDr0/c2Y47
PnnBYAbjISRJlNDRJWAqkFOFWFihrKvj/JyCLjpWj9TOvTcbAouw2WNr0+rO3E0t
hRGB9fdfmLQyNOn+7SNSVoNVc3g769uJ3J7iGM9xs+oP9GzCk1OvL+tkEdufURwj
lgMwUrEz3Gz7RTrMJ9UDBZVbXc4cn86D6SjiXm9JUDX6fwMSxHySL6xPu1BuJoIc
bsQCZV/FZ1y9I/XnVvEXE43qIYjM0Qq8wnsoO3OiltLPti/q3kbQgsWbUaPYRfUs
YpBuNh8Jf53zq7M6vA80O/l6SenOFkdPv7Es/G+8LPYMLVL0C/Wlc8j8kmAiGDXf
yMITX+SFj6IP4B1FdSguxcmjmHWnJUhJy4GaBBN9IEjzUqXut9aAaDRfxxjlwS2E
Xm00B5B3rRQujY7hgbALWbBwcEv0beeNsD2vp1yew4l6I4lRGXaUJDkaVHfjnW88
P6LZXIrFe4qj06aoISIFrRlAYp4H4w/xE9SV/HbcKAWMGys6I/57UugE7DC6alDQ
Z54AJeskMH4p6uR48QU6ZrbwpSav8KHPZ2J/LOsSWly+2Tut4qRQgepBVkj91Z/0
bcB2t2vUFGhL/JgMD1CPvQP8lUzG6Mhwyzyjk9AdVbng5El8EhJy9cIGd2JhU31z
RWKmjGlVtgn6tGc3y9XOeSpoewhlmeURi4XM2RXPLDTtH3kE9eQGcP2HyMK7NdIr
t9R2Vxu5+pGZUEqm/hwjk1Zg964zIExZ9n8hjvTPEujLIKkWeMNrcHRQM+PGbwD3
g9fEI9OErGHnY4nFB1PmYZoPZSP55gHBEvqZ/zWg+2++D3jmxf9s/ESSckwbSChu
j3kEtW0bhP2kSQ1EBFd65y+Tn0HiEIGJ03XyC5BhRIvixOeopHSOFnZFXjpSBMhR
QxSKJ7Q0n+5a1T+7kXeWLS1LyOAXwVu+s9Sa3oVuOvEB/ed6gsbCYh+QUr9OmFkJ
NkdweojufJ7VqAyWus3gcftqVLhfPgAa9wB5GKDUSkUpr9YHojA2idrKfS5pBLfp
CY4oo2t2yfCwOiuKG3p0Kv86nMV2Wsg8xPb8fdQGWqWlC44wM/X08cAphFNXKaFn
hHTReCUB7vKheuPQPKXKqJb26FIGTqtumjTypqkNXmpL/80rFSimbI9AiB3rioLn
k29GWThSc1ZalA8N6BfWhnFcp+mTYAw85CN1/cpDI3BvYJdluCbPZN5IpcR0q4O0
4AsS7iv2FXBSYVSoKHRqHJMn/InMPJ3QanqcmytRVhjsy6qFo31wkWC6JfDMQrWt
dQ/gvq/d6fvcdOf12DdjHYXNiL7oR2oFVrEqwtkSfGZbhXGTtHD4MNKYNUdCtnHm
L0C75An8Q3W24lwVHI64pFPhX8CW4hHb9C/8Ra995yILrYoyFTafscFHBrsADdVV
2NWKGMQcspV4GRw4zzflyAX8Jym85xM93XEMDjLeYV6f6hoQQ4HZTXA1WtZHwTdd
dIDNXbYNIwyrLQze90ndQucLOpYMxmlNY0UC41eOzlOx4H/gwwAi0uGBlLOtxiCQ
6V96MbdC2szwC8qVzHrBzzm55Vwq2xDHUygBjFnYHFpOYQ34kl1uSlvXcF9xh9Rt
D9XMmKwNIcVjPIgWiD/igAAhUyI6lxN7kypxB4K3PX2XL3PYa25helLnr2r9AWd6
oi+T4WVwqfBnNLYl09I1lqdqwQBsNWmIodl5Fb2/xP++rbrkCv/xcYx43rC3zwMa
o8JRlQBmkPi6cLVopFGR1A1Ru/mA+uIARcDaisM7Tm7v5xxhdH6Gqh+V7rQZCTt5
MdgpgwD4kJ/BASxDvHxMr9wkvMMDyMXqKBI/5C49PcH6859Vas1tPb4Bagkr0WH2
W4McP8IwydxMGtIKc6OJUIWB28n89T7BtZ2GczRh8R7nJAcPtceYSSof9U3sJXL1
nC/RdmmulaI9FIU07hg6r5CLxsDfFM93nG416yqwQohfRtK+wXkfJqpVL68b0fWY
p70rRH8H9SHE+zGmqdTLA1GuErDkFYOHBblcH1yMiq5wL4SVZl+cUdg6cwECGIg5
hSe2u1d76CHKKiApUzpyQc4tJV7VLAKHFWguiNRutEVPJuIcb+FxnWDuC3sWYHm7
byjxZzw4jymAhTlAiNaBA95W1xGU/GFV3RAVbmfRDNUP0XXmIhTB+XfACGdIAJXS
Up1+ZMdvloE4fwJQ1/HnlGv//hV3KzEkTpP1pIONwnOxHgduo4fbCBVR50Zux7H1
KbEphgK4zNwmYkX0d9taO76fNIx1AttJJcDbmELhCXjF41qDjiJG2TYytNadgT9P
Qjh0a9lBMjvephM6CM6LArwCBrHJPJmaUakaNCDGWd5Gw9L6QC+kph0wXTdPCZ/S
veETRiR8GIOog3GZayhTRcyvzrXZjRVCM2MbYlkt7gRwXIlPtBezv4qByn2SGNXW
qWjLB7PTqkC4bX3bPfdD7/4MH51FJ1NR/4Vx5z2fJOGpkcZ0KgnD+KTAGe7OI53s
ozGtFde7NGclC+K/zoe3xvJ0XRWS2K8Dc2Ubjvj4tzm+H6ZIM0z3h6RcCOW70b1q
MKIqqXaABvWNqeDRY8YG1NuhPlEvRsfZkKbsnusqmC8DS0HUPm+pvm3/U8/lmCax
QunNYlrOG4rlqZToHDtcgDWemVTJY0Z86C1ZzQY8E/iBf5gyeVrYDg2h+bdw0uYA
zSykWyEuT3noQ2u9Xi8j/OEMU/aaWVapcNJG/cjgk9aSyESmTyoR09vVsMoxUzSy
JAMJOYlQQz0UAwcQV25OuCzacjMFQivQ1/l9jimSdhQIPCi2WXxA/yYR0d8D5N0j
YFmJ7QDhIHjrfoQkdStETImepq7McTr2UMZi9eMMWn5Kj1tcs8A2w/tsf2oZv56c
rrkfCA0qydWyLtICWPFcO+/VsCNcflz2oeqYo94vKRHHeNpa3sa/2QxLyJ8sUzC7
29doAdOKUSluV+TkXQDBZ+6f5FOCcV85MA5IiNKgFeIcW0M6hJ/SlErCRZv+qx70
YCe+DHfJ+3AIPEuvw0S0eD2qQlMYUGSbeKxTtJNDlqyyqSiA5qQEhqAgh+7baimC
E7XdyMZvRpEKz173BvVM/kSMoqoKYvedFRDpuiKr8Y4gO4ARoa4vOlLZCesqOFig
kIhhc5YpJ6iVzX/EXfjlTzaqPhEC1aKTKMD5o54OLphCb7Zh1B6RgY+pNWP5xqRD
Eaj8lbAYGIDWVtRCawQFa0kL6AVSj6nkpothvWAZktxdgH2+TOt3MpHf1x0DUfwa
beRjFs9hiuLzj5Z7q9itiOy5HVzwXY3gzqUX0UxgbuXjZB/BvZLuVj1yiCGRcDG2
xbBRk0raNN7gGD4U1H2ZAyktz0UxBDhawfsXSHM81dAO58q3XEatPmj1Piz8aNQ3
LZuGPHbsOTBg3mCMIv9hRfLTvvkw7B5O9ukV7XrUl3+0KHGgnBX7A61vrA4+FuDj
iQpjlyUkQ07PnJuLhJCvHtTVkyxZ9imstOILnNWhZCeOCAW04aCPMfrmA56/zMMj
Ddfo5iSVwG6arxwoodcZzGixzwOydQ2bqc/MjWNvg20yAHGAWrMlj2UEo4NhDugD
Th/Kp+ledsd1wEXYKNsJcMUjZpyP+thDYJgUpVKer+qjn3kthP0n5T5BvdwCPEbk
QZD8yXd+dWX8dadtWTLlpu4woFgcyp6NIyWr5dQwL63Cdi1DO4e27U32TaC3wtni
B2MnaFwGiXavMoZ3Uw0Hu2QiANViwtM7MSqxk8z5FjKH0z4BQdUYTNwF5ij/YPpF
Nh0lhROVe1T+yXivQWuWYclQU4I54aNHJ3v03G1Z3XRr9MTXp1ZRLpvm7t80pyUY
sqqx6jnFOlK0DHga66Tr7ueJiABfoR0Ztsi4uhqL88ibeVVJTtEx3nvjD9A/q/d4
HBmvsHKE/KlCUtJUp+VCI5r3MWTfDmd0jrdA9n4IUEpV8mdwwxMOvU/jAySXjmXy
AjofPYUgEUsZpRdP9GlolFKDeJMyTUjPwO/d898Ja3nU2T2v9hCPfGtB9GDTyTwr
wwq5l/bkz+BVJEvvxzR4YMQmqLwbo6x8r0yjzy2iBA2KbsD0A2631gXYi8NKDbKi
yDAktWIBTHXBxtznHyz4Ej4aUI04xQ4kdxqY0NdSVvDfTrVuLJNGXKaKUKOhfubs
2Gk6UAAWMEiuiguUdZsaaHCsSjlJovGRCEaQ3SInijxC3uc+TR40nNG1S7XncW1O
DwD5vjYaCGyQsTWacvvJYaVHAQcbhlrVKIYdZS7hyGbjSRW+co2MwZ/ddGi67EsL
QZRoiSXVZ3Br5ec8hYiydYovnSv1tI5WAQrCOmkfX4moToaTfVxJ/HvDBVFQ9NgN
K2G9eYIAP+1LDITaqjd1MjjTNWcINeTCb4KH6raedCL8D0VA/YS/IILdcJR/Wyap
m8ZGCVIQp4jApxXF7cV7C65yZxc79/j9xxLZ3gwMiDeBRdXxpKvubQTJjI9ruRSs
qvVCvqmyUB2Y6enfgKc1rQYICpA2Hm4cE7oANQm2AMlaogYn0CP78Xtzw9OYx7jy
7Q0vs1rBqbyjIUPECqCsmI9kGvsAkB+RHKc9vjCEYM6kx8zhK6DN8s0XKYGLGlTd
a7L4D1hrZfnRLkEbBvaCvabC7lXvUXo3+RbVA21usS1xvtHXdnty+TyxHRjsUEYf
ThCl4brvamBMpe+3P/5nfeju54WFBgFPu/i/rY+Q6VScfOWRtvZooq7Jo1W4Ysan
DZopSH/yj4PL8WuB59Fv26uWnA+wgQ1oZTXhtZc0OvxCyFxKZtzOyY8brJbdCqpM
vEGL50YLdQuX2JoYsrZdHVF4ioNHKA9i6knyZ/8QV3x3b9ykL8oRAMnMQMK7+8yK
V+p5FV9MXOfP6HWkdxXTqbX7iFEgdZdkLGI0Ke8/qrj9/ecbbhVjBaiBxZCLnt6f
GKdAfKDEKVfC3cO0861qh0Y23IoOKnxMSYXSQBbnEEgO2xuspJIPqtMfT+WS/qY9
aVHqfWANuFt1icc/aJ02Fa3eaj9m9Ic2HWnQUPAKC6WjuiRiPWqpO3dRIFxzOB7n
DCWyfjaOLUqA7pQRbc4LYHsaPqujV7BM2sboi+aWNEIOA+WYkW++eNUEpKLJxSRd
HJvWQPX6tHJzZ9aRo5xlovKM5IFb/GSoqV+TuV9c8/ydvJFmxCeBZwmlHl9/wHOW
c7xX4eHkHG7VBnBa5g5RS4naQB33L+oXHXVzHqkPf8Se4Z1n1jFpec95gGJ6FNd2
GAvqCDOQATWggTL+sCxqNGs06dB/z9JjhaqcZUt6P48CqBDAyFu82Qe8pVEX2Zfa
VSiVRiJBZCPf0Q7smjkGvEQOheDqHmbOMooFHYmizDVax0nnF5rn/aG+ejwQhKIl
GsXovv1aoje8oltsbSfgHlIix9KG0lWW3CqEcJwrEz2LjsXpQVbybpHXIJelVF3V
lGrBd48k7fIIQbGEsZGI5JgGNUwPTauUfrnA3V5yZyqyj3n6gNyFAqWUiASQAMOw
IC+HSdpOanA0Ub4XdvORyiZoNFNhQhHA42mNz3TflZ7Fy2BY4QdEzI+Zdw3Yw+Y5
Egeyi+3cFJtauEtlal9Hx6O0og1XlpkvvXgS25hjbQ+FE5XlWNOzVU7nKFqrJg8g
xLjhHtIG7fDY88byfl2DgSj7GWM42qZI1sFATSgqp3ofmexSm3qpAd2RnjFA0lDH
TWBEW+0zr/IEw+EyPhlUL7WgGXvC6N2lxV6tBY2zFLSjXTGmL0bl12wV03cYlhJs
i0M7Hr0RKJ8hSVQUgYJsnqTtLnmqmktLe/eCgWhB47futjNj3YungMb8IHcWBMtx
yjjKr/fEw+rH+5+7XT1vP/9LVcvR1A+2GODqBACaxQCdVMgM4hZV+caABOW2CCIe
x7nDcdStYFrb1Og2iTP3LNN1imlOYdhxgK20qjfC1+OsCMvm83icE1HsUmR/6QWa
NlSc8r3Af1j4i9qu+jmP2u7nXmdhr/6gfIcNKqxZO5XjmWm3fCTcq7nn4qWeXwwe
xwyqW7L86IaWVuoMez2NEgpjQ75dI/wZiVHpIIrZY3VUgUn5oM8dN2v0vtjsaa4A
XVYndGgfWyaE+cLgtHebMlzVlrxOmFMbVK2C418MfuES2i7yp4RnBLbk2f+hqKh1
HGFxl+6xIEDJER9afB84YGUoo7p4Bd3c6GiL1McN8e55WEZBo3NZNm4RctxnOpv1
4KuB08SFv97gQjBDBYjJf9diQwC1PVJ3qyishkjuP8ZnzJPLzrODR7J7xF6FZ9QP
SsGeWGmNy2A6a5gPDiKNusxDMoQSVkMQICaE5obeb7Qf9YE8OD5aSu4KceiksGiZ
BrvP24P6riXN9h6TtwmOMadb/AJon0ThL1FZ8bgYHQyWHtj+zZa6yykXCdCsOx/T
KAfxPfCo05onwgr/n8x/8REroBoQb5tMiEWxHJn/ne2fR6j9mboWrMtYHY93yuoZ
TOu8t22DLhX1gbQueYcF9zy3xMhOy3or7NrYpPp/qSA5jCPapNIg+KZ1b0edP2k1
BGcqBMjwHAl3UOcqI0A6H+cUfos7k8al/HPMxdrNmLygq3ZvvX/Eyn1MpMgcTMLr
JiFi3ahuRSIVvM6qcMA3TdawdIrnVzdha7N78ogllGl95SDMFF2mqHJjb6Zx6T2k
pGQ8bhLK92PUr25CSy6iKx7BPkSBIswVGpB7PEEt1hzzEEGq3UJ7hG5jEbzg1QEf
e5cfHoJhFDcTiOpTNnstLC6ZfG3Iv8eusvbMrRBuCCx2421LMNhqbnRW5Nay5fDz
tO4nk/JZl1r+jcOJ/EvgKRezSv/+nHtoIgGDIy28t1wSzxvPSjzklEr4uW5XP3Ev
W9zzmokDZ7MpkmUgTG02DEBNLvAfzd1CXdJJe3CJBOVjP+T12MaB5DFqEq9/bKTN
mzDYqtHy9Ff9AlZk9MGWbDa3SwC5NTcrhdqsWQYsuMse5Em4CBEx26loyF3qLvSd
R4ohhODSF4xjEcGGeSV5mGJHi40kOgPk3EV3jMt/dxO/X0cxfkEKx44uuLlSyjuY
OmIpGa8+DcwOnYrwjdqf/9JAc7p8eZVz+Hb0rEt34YzMM5HBc/bIzMhijQWeLSNW
fSWlgYaiu4LJUaIcXjjaWVemf9gPU4T/o+xpt/+LbA+WyeQIn6agB6qvwACNGw2B
XWZ1YZmm9D3ZiJ+9I+cp0bdin1W2ISaI2r2Nalaaeay3uGe3lC3+MeXGUfG8Zzm3
/04uuoQrfJIgEVqH8lMa2hVzGJ0TNiALTmiiZ2JwRuJHf9U9fUg8beJ9UMKIiYx1
Y91BzmerGLM+SxVOBq5MGj4HS5hwx3El3KF8VI/btajAfU4M9jG7F5YBgceiMIG+
nap57Ck7xCz+mp5yLfrKqXV6/yWCtET44t0uJyXXQ7agKTHAGYCF+lfr5mkOXgdD
ZJwjkvJxVDQsND7AMiE4iTyo1FzaP1QJEIPDpNCKCMcTWp8DHs/D7IWan+CDN4Q8
uCzBK0YXBBwGndVbqdgY1M/BuJzm0Yp7qsJ97J4UPKFkGcxeiOX1t1Jv4WdcKaIj
6xmqxZdc+xlw8ivSjBIw7cWhZ4tY9ww1M9pxMoA2eCxb6ELOu4pxVXvOF63FfBFn
sI0ibAWuO3SqJJtiHlBGHovvSUNgHFHw6Fblc6KtZXnJQ79dt5seOPOttNTDmQwj
lWTiKdIcPGigtiFFTTm6gWzxHhP94hwBNmRk1LuyR3vuEmy+iL/vXEgSt+YLLyGE
IgpCfqf8coMg1c8qgljrokooaHZNms9fAekgQXws6o6Jo6WrdF9K893Zyntb3TAW
wB7Aekn+4w13cI5p3CITaHThxWHGppKz+4F+LU3eGwzRCMYyqyJxSKz63T2qiN+6
KQII9OR9hifOQXad/3wtXVJzcC7r98AXJS/rSb5Nu3nTdlwmkpNPF9MFa7tjqTQV
lSd/6W6lnLbIDXEqpzdGbrV1WvC7GeNAQmcLHj8AD6TWysvQZ5+ywLQwdxD7H+Dm
PI+aoKKHLtvVOv7MNu/a+ph6Vio56q+3lQpOl/52+CYgvS3u6aV1Iv5N6n4PJY0v
elyXVwghFEK+yl0j/GcAli65wqT7DD9AOYt24Fg5XmCal6P93GzpfJS2iEUeRIQm
hlP4jWEf1UkS1BT7JGH4Rrt2RKCcXto9QMYeMEU6+eAifxDcvQGUhTQH40BZr1Bb
G0e2FwHrovqAGnQqcMqCxpAL5+GJEdOh5N+iQCtDZqFv0pdKBLOlZYQFLNHjAvrX
azEGVjo3VCj920vdgmaOUF/zzrn8AmN7U7ufaymM0A8lYHW/k5vpdnd+MqSjnON2
JNFT/w2ONeDF0Rsh8jW7xweuytt3ZABWRcmyr7ybTIyyzh6he7qdN5PPGcdCZuEt
CwslWVdQX8PaI79IVap9JNmNwe+Rz4mTtrrmZAiMtDWOij54F6Vt74adWWWsVRqL
k++ftQ09hZppwtt4osmZp0AuLWS/Pke/INB98HqTc3I+dvl3KRiUYLVgFH8TC4K3
XrXfrvA94rM3TaaHOU7Ks0goiFa3tEA/ztxaSG7kc5mgDDLctV6S7DUeeuj2PPm2
hQY0zyoKuCHAq4x/H+rM4d+ssZ2P53m/vFE59XOHp22w98BaWGItBlDQr+Bupmv3
Hq5l8H3QClm2iXfDr6YAusLZWwiSrQ/0BGG8wMV+zWXqJ0piYhxgX2l9W1ZI1VJ+
H+sMgLbAIFxf/S/b0/YCExTBRdFfkRCe+Jxp4jGlgeUBdMgSwEWqNfA2Wha+EHfS
NQpZwPK2c2xNZcWu6acDs8zcoT+RPVUQHj9zGEnolsvIZgEUN0PUXq38/6Kmm38f
3I/0yeK1vgYAETCWSdWdC5QIhJcIN2ktf5UEZ4IdRl0IMyw4zuPs0zxebgwl8IL7
q473MRxdLjjAG0Q3d2VP1j46Ilbn8+XT7oTjwadcq8aZ9fJ+Mzzn85QlkPKz9eng
32zTEWK5vjZYcL3zM68Gc2fJuqN1Ur2JVGZa1DiqsSBlwqDh5KXBprjw61rEKs4n
+SUYMYY1cvt7/hlpfdKoMchihiFAFtiLugcGy5204UAqBAtxe7wDU5DsTk3spZ3h
xXur3OP8NAfnwn/oUVwxgQCrU6ToCaOkcf41teA5z3lZrVW4jNHlqv1lzly3uVnc
J7thH1m2n900ffI8IwvjcHQRkUFBTWivIb6JAWtx6CF4htrxYi4zwEAj3/dhwTqM
tJZugubs0wvylUs0gSY7hFujqUk0HWNYiDBHxp9tFfibRhze6e3OhIC9bQINw+IP
fhagdPeLFWrVK3c3unAyKjZefki3kt2hrYMVMKsJGh+sMNGhb6OO0vrZwwB+Eicp
sw3M862YwDXvJpabxHziV5LPMQKi4k4WUCiByT5xspc6XbDeQ5Vf+0S6oNYqyJps
ko+oabtzmsu3msYi3yIrsFC7to257L6RgsBZCFmvbkZTZkydF+9p5VZjrewoVAfK
JA2uc05CRmR6x9IIojwWtNhWNkBge8w3CGi/5pipOjbuc5GUOMlwM62KOBdMVzkP
odejdskGUkXqSCAjDPhQca/FLBZmtk0e7zs8KzFOtdiEr3gO+R8di2H/83g29IQr
KK/mctPpn9GMLcikVUNPpeeJJvD527JdRC6TZZCSy0ADGiVskFmdn0M91KYL6J4g
BLGH5xqMEVquZgkXgrQnrWNQhkDfcciIFy0xmMwDSOLrN2f7T/eeoHNDCPd6eGV8
7BCSuW0zQIlkWuToTMR/CjVPMKOwIY4M6DcyQWDnAWr9QG88MtOwLRNqjFMGQVTy
cYPLT+pznLUVkkKEKZbdvADn5milMUeNQ/Yg6Fc+paBVyb6iSd1uqX/8CUfYMfk3
BjJbVJqhwDD6FbCKtQ/LO0ZW48eAd4vPW0EMLoHNI7vO44yFtGe9TMBPkh+LJ2ta
hNuCLv7tkVrCDuz0MeJ6AEh6VCPW6e2G5Vg6TXrsuOjkdaONQAGd3NOfmkpMVn8O
jlWVpuDPFBd2XW1yMwr7+6SFXEGrQGz1+2N82h4epdptYFMuWvst+mu/tn4Cuc0i
O54bQOGg0cWVlxznQ2FMaqOLfkYVygSnkT3zCuE4M09J7tBGIxHAjJnKASE5hzRk
xVSbNOq+sc3itsjhe6Wav6EGIgcs1ruls3yib7NnUbD+rhcLqrsXFvEwE3R+PYIz
5XXFYJKTg+XGh45bx5khBHD9BKZqG8/JuLJjZNuP39cTURWRlOUguzKC22fUxxJl
4LQnsuv4ozq4HnWraBHE+YhduApxHYgmuIsF4ShUx7u4yAyEuQMy9nqTdnGHjGC4
xLO65+kAUzFVYpDUl97LE7jpufMwU8rfyzBqW4oZY+WQPu0o6j6gNypZVAM1c1ZP
ECBWogCC51aWxIfJ2cfgFoQBSGZ8R+slVrU50up9I/O/pbWTtYFzLpdQvzJLV2a5
c+8fUtzwh8iYVZPugKk4mLDVjrqDTzzXDTtpwDqavKJbbwlGogsesGKThhRdl8x8
ycS6RZ+FL0lCZCfz+NpppCkxNGBSgZRzAAO/1QeaLAdUJh52W6gb+c9vaohRpJgQ
B4XLBELwXx5v4RwhIYiAaaZ9Dj5ccwIOaC9Lr/6mE8TQyOcoL2B2I4HtLaZNDKBU
uaBiszt9Xnmg9QVuyVHU9ZlRwdAdSSuQlkIluzVMpd3rgL7tDXW22FqXfateT7/H
eUMJ/IFZOCGKYnzRh4fyS7wljvOlyAl9mcM6Q5Mc6GqTW3usOT8IjaCGX714f6eP
p5yQJd1R1LenO/3MpE6OHBmStvAFKcl+2o2pug1y/qjYSyUzCitnrGOB0zT2uVHU
JQOmpkbiF1AqgNYqvlgd3iptlWf8B2KjkOgm+f23GiluqVKzk0tT6AZ8Eo2SIYn+
euvuXOKPA1c5xgiafx3TeT/UDxvMmngnpdBXry7xn93N/CtuGW39LT5cMwElN9zz
2IYgSKs5FSBpB5FBNDL2qsKZEYAznY11AxwjFxBA/qt4iJVR9J0Ykjj2Rc6ccA6t
GRoNRSoLaXZoSOJIMTR3OqeX6XxZdV8XK3XBdExEMRMNM1GB2qq7o3LQ5Ykz7Gw8
1a9X6RCCXiBtzg1C6Q+FnSI1ZQ2V5nvFlHtESCCRVqGzdYhOIO0fGUEQdf7avJOV
g7Izp/w5/EZQf2pYSImakCgI/hgwx/oLNBh0s4al2rIEa99SrGIIi70ft+4N98Zg
8wQf2RNXfv8uaQx/juOF58Rf2oX+jgES33xbA4z6g1ZJVy3wcTvZDxBLD/TyvmWe
M4pGl/3K8Jx6P7kanuO3jDFzwx4kkYLrIjREkGtGGZUChixTotQ5z9D2L8Zg1riG
Zh+DiK+Dboz/vGERC0Ma8NwNfLd270ZSyHMrxsukwb1Ra/blfgBG5wl9K6gSJQdH
YHiUpQXAXrZhf58UI/1G5h54ojAo967/5aAVSBEZ5eYZWRo9QxOG9tEGU9kbKmDX
IHtjtfASrB1Qcik3JBLysszY6kMs39PicYJuFybnwTEiE9KNDl/VamyiYMFibXPn
vmec3VhARhkEDBXeUH4Z5HYzsc+mGHEmfxBLS1cmIr5wqVGZYY6oS7ScQJq4WnTe
xA6Zw6BPfzQGCypuUD4yiLYJI6/+AEk9e5z/hcLGr3b+VoxjpTkqj8iJS9QPdK9b
ol8WI5I4cNFAy0qqGvB/mVMch09IoPHchJb46tO1i8ZZ2jtE2T4/QEgg+dM/2fPA
XJQaS5xW5hDMWtxy68RRj0Y/UPboM33O6xSUps3kpJMPe4VNciQAwVDCb+cVafYk
Y3JsdzuIsFpS3T7bx51nJ9/udKou76gvXZk4nBapqraRask8XLRG1AZ7Rl1whiK2
21F7nxrWa97CuPuiEKKpGRAyBJ623yrkKz2j//8yMi4hs6EzwkPvEvSMiOcDlWi2
2ISafhOxtcPDfYQ0xGkLVm5WEaSH0qxC4Ih3BXb+wifE0TI9dtJw36+GKYQWiyoq
2ESOqBzGiEzkF/6Rt/vbHTW3rRQsAO7DXU37rpmYVpRw1Ogg5aBCNBcY/9PoHXJc
XD3jEjy2GhAKP/QnEIM1nIi5meA+e0w2WFpn2/c93Oh5U4YLZVBoHHcs3T0/ujky
o+kcDXYMW0vO4hClGbgqpD7X+2NL1zsbi73drsw1lPlzRlBd4gislTAnnJNBgbAe
vmkh9TZ0UbkCzHj8VhctCNeJWWskFTiqyQ+SHWezAQ3Zo0VaIc0o+w6qJaPwokHv
EXf3xOwcYKPqhkFU0oMg/K+/av7xWlT0zEG+TsBjbCmbkR6tbMsihkjCnYjmeoa0
3jV0rzviPuKjfQFsYOH+MO1p/8R1NNFxDLVb6lepQ5pu7P8cnNrfN93IUeIDYnCR
15Tclq2w+3Fthf5zdPhsQV8E8tx2NC0npVwtpGOXLQUvWCI8ER0e8K1RolhFc8Ep
v3bIMHRyEF8I6VfRG03Svq/i/7vohCBEWpnwW4rXOk+EEnrE00MK0Yx6aE3OdIWI
oTQ6aLuBcOEaOpOswfokdYaBd2sMBQXFihMT/akQ1pFQqDntVoJiXFVi1O6WXFXI
wUXA9U8h1kPl44pIwRtMOQSONUtEsNWZ1c0aFRudM2Oyi+A7OcorCeav0nHx8oQP
WdOIvpKiKJTfOq5cZjRg9ArqWqk3ITdOViMFKMz9yMv7OqOl0iF3ROiUdGHOa0ay
N7nYo0awZwrE6ZZP4xIZa6eMfH1t8Ul84eAAzWEe+CL2E0c4sCFfQMPzECg+2ONP
myFfCBA3E5tkOwJUXfncD5U7tshTAlgoRZfqcO9S9YDtnMsHeKM5AtZxDxFeUY8q
zyLPTY7Noz7We0q5/lnAqh8kCio71mXgk4w7D3v2YhWDM95XQ37b+B+DA3VbKQYb
tX3JlwXP0VEFQqTrsfL21tVgdrOQSdz2Zf6Pk+uyF9luiaDM5mo//ztVZElsbm/c
+9IHUx4LJABvYfNgaQkC/Au1awrNnNIgswGKnC9AWfnP1e/fQeb9ooR2Mq/unr1Z
Xg2KvRTFIeB6w8Q/bWE1el1pgsUFdHOdkQ7SorpPQclTzKkr2W7iB/000iOD9Bmw
nX9grQfa19XjRUYbxViZdEzQIJ9f6WtlaiM5S9ovL634B0XqfdlMMJVlBVStKUGW
CLKpiRqMb9e15FHYlwrJCH6MYsMUvRNbi/VJ7KG3suooOom3ZHJD6SOkWU1UU7X1
99o3n/IoZsxtGWVWIVDLVK+qPRjDurH7tOhe58rp/DX74mjJw7vsmBKv3YUvtKQQ
OXXgCPOcgCMPaXfEP7BYo+o8vPQh9I+sarntnVZ0mWbTy82WS8wkZqKSJTazMCP0
436Q5EjN2i7JVAOgNcVIHIAbddAo01JvW3IOkA6zwd1l6MrMWYJgcJ0o4fJXef9F
hEmdYfi0OyoCd8924mH159WsXvy2h9B5t4dF5+1DXKYR3sa7SaL0+1FDWGsZnUed
+QYC3a3Pdq6HKI31bYw6zGAV0O2t3VPkv2vtOkzqLvLAVe9ySxt49GT2no0L4+R1
NedQbD4/ZXCnxe5O3+FPfVvVQTCCBNWdSOO6BazTd+MtqJVhT/wsmLKhSQ7UOAyH
9cFdLvzWDjeGrsd+D2eSs6/3CVjvP/Q0sutYpZ3AgMigm1Cedz7ZuKaNk7hlvAhm
tI1skIgrmV2tckGCHIQuxu95dP6T/9unKTRsycoBiops04Fe0zCgqoe5w7rIA9B1
owAs/93ruhBThV1fsMRjKG9InUI4No4Xm9mjUfXmSHw9f3vD95BACcwTHrv6ltHh
MlVDI/O/Dv6Z67o0oR+elH18JM0V4ZB0P6H1Tl16G2bZ+H6N33TE4eRDuj7gU2V+
6xfXSNX7jnSGX5t1mn1CzV4xSbejum7Kw9J/73VHvEUBoyENiJOxbu+eSw86NL0q
n+hL1UwEMTs20W+gxrs3TmoXZWkD9388X9fG3IOXHqK8OcvRvvXgyUndeYzmsdKW
oHWejZ4JUo5aTBKI5gXbupatMFGVvvA2TuUrhKOOaWiJb4aWQdWRtmHvdOVTHxqg
fxnzt1NcLWwnumbjN0EDsd3eyZhHqNk8tQ9MHBrnBo2q2/pdQyzzATDbwl80kUN6
YCs+bZH/ezmwlpyW3DoiWudbLjjzBtEr+z75NM/aaZSARRiITwI/y7SeYW7Lyz/5
/3K4I0OQNK0iDwn7OJw3oKz7zNapipaE7AeEmGBUddI9xn8D8mF8uImZ9V0tExxD
xv4esYO8jVHDsi2CqiOa1NE8ErTXRIJii3uz6sMgT4YvyClzaiiC9xZuA0yvg3BG
UyJ7juqGatqY/gIRyODWAk3xq9own7ThkmB4Y57hsRgDAEZETAXiQenmjS0TdXa0
U7GKrmPC2qAItLbzt/32z0VljbdCCBGDi+e3wFiLeSlRE0oInceqMhBFsX/yNbUz
aqyAnQaLje9xC79R6peXVaL2RjC9uNZlt1PYSkmhVYizZisiWZV0hjHX5Rpekhhl
85UZZu9+42ErCaMqbCPozGKwpU9dvM4ISnombZj7gy8tF1fwoVxfRZfIrgXMcDdQ
/MXTlh/n8IrFSCImPr7BV+dy8axbDVHLaenNUUmCahkMYu/jYF54jmc8HBWV9ZtT
7qL/rBtC4EPaonB09HWHoEFJACq//pj3nTYj/NDtIbji8QjrGuANNQ3Ti2z0XKrb
YDZv83Ds4dYiMEsX8q8/nIO5N9NUZGeeaM19DscIod9LWWwr/2Nl6aLW430dP/Y2
6xcvdJWVDuFFaaHA3DGvLs1eCyBvqCxOQ4RZNnW6OMFO4w6N8kmIAo903UL8uyPt
2KE02QFNjzAqEpUdw0o/fskBGwo2t1M3HAjpdwi5R2+zeh3yAhUwDyBCF8dSMTz+
EdJXcp3PF/eJVdIxuW1ZXVNWLdOMXjrCG6YZkRNrmL2zq577B7GJC1i4PWxyNqyd
0OV8sQrJioLTltNO/VGMruMfW5b2KbJ4vyQ17YR6fQe/XSr+XPqfGYRvG8M+M7wR
bCCFLlOT8tJWzSoZ0RXWN4f7N1CyZvMywM3f5a90rHBjqOYb9ZyrKlKPh9uJ4N4Y
mqYGelA9KlYRHISi+p9i4rcBhVShEvh1yt68tNRZCHPn7i1EBkv+yvf9X4rbedPx
zJqHZXNbiBoCVTK1v8bx9PX/GMLimOoTZHcEQ4K+qaCSp5m0WdfGL1edCifQbXT+
p5vSKUZfyDHcjZr3/9Ka3mkp6RQb/c9QtzKKGBYOq8yrwUyUBncpYMC4ge93qzJQ
M+DndeHngV+uWiWXD6nXKWTAXVujonEAizsXGM5NcCKilym22Gt4q4/DFUg8jgEi
3KAvjeXrAafa83eJ1y6qeCvT7e1uIl9lTlKaKtSiJE/eu5M4thV6zsLOBDWm5uJk
PQ4x+mxdK53mR6gDaH6l1/Uuv7lYbHvV6imKZIHQoBMHcw5EUaFybSSPzA7FbiH5
FKsna+cNjrvvMOVr42A1Ph2Rp0eCDTNZV8EpZw/gKWRl5sGHdXf4XeVqCteRRzxI
oFJagytsKj8XSwEQCCgwzKHBcyLNr98YvMnBuLJj5A5eFfeL/d8cixPgkc4AObLd
byKLjFsrlGEmLYoXJjPLMNReCfdr4Y8btXJlCprAJQG/5xPPbNaPiyk9Zka1QsLh
c/IknsYLqOUW6SnRqdJ6Hkqf8r/HkfRaecTp91c9o07IUpS7+PRj/UqT3rQV+/f7
OjBNF4aRv2W7iP/kegdFcxGe1x5gVvpvEEdwJhglqlP0RXbSR7u08pyaLkkse/ZX
Sv6CPynb957MMJjetF01BGuZbOv0bLzGMO6agSg7hB0Nktand/RIIX2Hdgn29s+r
4o1pvqPFj5cbOFtOvolKzZG6vjsFSW9/I5b0G6f1Pcj9KBtkcWM7XuQu2hcAW+vB
lHhH9tYUcv86db9FCbgWnRJnldchmHoN/rORs/gJnB1RqfXXmSIT6laKwaPvyuqQ
XykO4j0mVHpAj+3C5kF/VIgiscJG9iLlGh2v8MffEKmnoBAvjxeyGVRJWrRpDahD
JqsP7K0QoVXIgkjyyo89GaynqzYIumnGIGxmyNzNukSDf+haISYsxE9xQAlEMV1N
9NIUx7sC+Kv1c5BNr19+acL9kObtrG8r9/5hQ17BN/VxHUE/D+LdYhhZVctWKwKU
+Kvg+xSjADKY8nlkwhbIfmpOl0/RGmwLPlU2+mnoxZNLefRK2bRVcHVBLrm1+LVk
VvcmL9nWtiU0n3Y03jHTaHn2UICNh264sx8utVvKuHE85ECZH51L2LuGkqEhApbF
DNOaQIq72sqFVpplgPhFUoCkf7B1iun4lPVPxUKZO6k6xDgxjW6s5k4M2Ge2fQAZ
1FW1pfExYgrL9lj2n98TlZplEnmIY3gD/VTogbFNgB0Vr2NYW+K6WMrbZpMz74J5
HKLWdHWr3cgEffsbuCHQ8KyAW1qiVD6jnc+dpLmkQ1SHIDnDwrvePavVhDBSMVXk
TUfApZyvwXfGJ1Z8AiAhOL+KKTmOehoO91G3LbVBXoUtax/O1rBcB/nK6x09+X5u
YalAj+GwIIMwKx2zuyfpptmepXTxwXUxqDnx6YPvWv2vY6veJ+LOy937KMjcJeGq
LRV56IVdWp9MTisdR2YxLDBYkA+/07h28SrrsXMw7NMa2kXVzG2LY7947TldA45E
/OF2+NHD5HkM8LLmhGk7PV4Wi2u94mpq50d/VaQ/HTDG+HOwH8tr44SoJERQOnl9
fHYwRV0gR06cgPsLfbaWShJh5Vk4RmgVzzdoLLY8cbHfAJESkU+/bebFiv/T7hjI
V2Q8AqqhsCoV2I4icAZrSZ6xrXACw6dv99zViPWtx9ZOk1bM0mPigd8PoFbmgN0H
UROOjj3EWyAkEoVF5mTnxyZERu3qpS+42YpR3jXoja6+YeMe1nQZHOUUoyjJsTb6
gQ+TFvizQ9eouP+OD+9wQmRH8DlGvTZQdVbaroCEKzUDM9a8Grh7Ch+0Pw0kLHFr
as1CDFF06ohbXyNbcynBm3g/+IE6FTyUAk+WtM6BktZQRh7h8sFY8KBwrNkrSiRC
Q7Kp8RTIeeRBTWGzvsFQYaLkQaYkO70DGfXxKUKUOsJ/e4ZhMJ5KQrleLtIMp9jQ
0ZLzuHMLtOcChIfGEQBCLJkRzdB3x50dZGN7dB+/VY6gkDZtR6TJpXVS3BQiWRkr
DB6zAm0qYeRI20+gCJyu/3MvGL/SeRC9WKuLZsGdAEn8Zkvm/z7vyrPFLYYLb4uY
pukIjP4ktUurVIXlUZUhYBm3dNxxVSq4kIvlYmNUKayackYqLUxVrVoFhSe2BkRa
gV3DSeSWZ15UCWXOHMkjcYSdn7WSQ8Rc3BqH++YptDcT/Z6+mTKgBTfFEG76cef6
BoqJqsf+gYjayhPYzi2E36MmkbGwO/hhE2X16gBiD2ijmnJVXoBnfkrFgAEZT5Va
70iqmuGac79s4qm3OxDfVZUUmugJweg/krdG5Qi/LCFPVELu9Ltv/DC5Qz4g6kRx
Yb7NwwIAuMcGVwFktjkRTz1/mz7TKLr3AwKNeD6DLa3sQtQkpU+drOKh6av+t4fm
orkVcu0BkiqW5v9bwJltYNpr8YwrCNxdjaYa2n/1KiYOJyWWGGw3Zn+TW8O+39f/
/0pSClPnHc9JhXDE8RSvcie8Nrhx/CkZz5lui2WFllChu/CNrUMRujmVqZ2+6mSk
l1lZG6aGfF05S9jfGqZGOfvz0iFIRyst/WyraQZDrBRuiP0173tWyOClrXaGlKL2
Znr44C8pTEk/rD1LHht1U7cWzdK+57+ee7Q3D9qHocmIt5RdiEj/H6dk+3pUM9gE
sFYlDwdG3SfgSMaavLz0ilOsdjKCTzoFniiOdyQODBX3mxq8zi0aPI9q2ET8paWR
RP3i0iZlcM/lWFVLMxCPc/FG+S5KBaisJ1n+eqqKhRyPpsri7QocIKww9m/boTKA
QzTgN1UVCwUyJdd19nvJUimFDIwP5WcxuHqOJDf4u+yOjoRLFCKEvVJL+2v11/jC
6wwHSzdGcWD38W0HFTUk8W1KdXMgdPEKv/Mc9+NHnmADWQkfGRJHsGvHRn1RemNt
oN3BsOPpKahlSeJYBbTPvV+kl/zU4pPuOiUmfz17vwpxhjLTC6ocpLHaUrYoybPk
HSxA8y4Od+OrRhbttzyHU0UC09OsrYSw+YAwAD5goDnMPG3ZtvLSgeEIoK0V64sP
EvjQ4+nlToLIz8gVI9onEDdbBjAyuLyHh0t2uqvNn7C92rwNbwRNcxRNxP+dOGgA
IS8CHlSKYOMHYTWOr0oRBnsjJb/89eA5Mtp8nL1qvDT/bEVRYzfwQq5EYKNopLMB
t67IuO2b659ZxRtmU+gYoS5blLWNaFnKXj1+DnsYEiczgyg5PHrvufplMQBVdQtH
Pe5jYtodM3Mq4d3GyHhB1z8ocrjINY6qxtQp6DV4TSm26Im+UlWsMsHKtUZnAvz6
IuOiKbJucaHFWnMcm9100uICA3IkOVIzH+cWN1XQmciej4rd7iZHs6PCrR4nofW1
tBdrRsTqC0X+1YYtg2y3suJLcNLvGkmtFmH/QEONrrArqnsj2OnZLS47aAkqQHfH
WuDE0f+fhqft3VqS/vBQqiZnJrDOENQkxyv6gEXIYUVjpeyMnboYHKO2F1eDpeNZ
Rev7ni8g6JwqKkkD9yCgvADuf0xxTEKbLVYlTElZa1AH477nPrmPlue21Vz8OnaR
Od7FmC8fzlyP5X1E6o5v7LtAF8V94xoELmCx6L/dtqLsDpL8M3rlfrrNjIxqLoLx
pO07qn4bRLoNZ04NFFlK47miuQiibukiaPw7C5bSvu1QSQ8U9qUQzHzQnWTwglsv
CVF/OXeX7cW00DE+T/fK0wwqyR8Rp5p4jeBfajScNTQfU3vRfIaR8TaBnNsclC92
Nr/IDl35YNbSWFQNyeLdgFTeWZmcAZcY2XkSeWD3VX10+Is7TI+aKQNUCCjcL7TP
33Wn7uz/0eCQcKMpBI8NUjycwFtvxIZ5pY5f0fKv+7JeOkuqV2lbTkBahMG1tM+d
lLmkQjbqj86/WXw3T2xofVpVMVx7cuSRLJ+0mD4EdNjQwjyZYNYc/fZh8HvuC+e/
sL5EB8MnWPOLpDjssHaYVrq8ts374tuIfmKtH0frJNqraTkoRS/o/8CCHUqgCgL1
JvZ5lQL1xgbpgBb2iUE5hCa0AkyREttw6sPoPZD9yxJsQTtety1SdaTE5pg+OoGk
Azu+dczDzthZ5crQ3cK2c5nTTMjKtaa0SEEXLhe1KeJ/SVIY+8dyh/1/Gh0e3By0
ksu+lMg6rjeUxDP9Aqv9GnmelniIn/q337FHivRnOd0ados8mX4dK/svklJSAd1G
heFgxHX0xoyBi0X0OF127JClUaPolnVYMXmghhk5mhNxJh3vtQ2toXvYp8RLHRkJ
7GEfkofzU5J878wbf2Ky8CDl8GzqWPQThj+y72spXk2w0W/m3jeIf77AAatHmwfm
/5tPZEFMpAWV0FncNU4ZPEMr0/YfIHzGe0wbq5eRB3hdo/Eq2QzYCfTU8ft58P35
qJBFEE+o/SQlHY3L7WNjo2XpDsh3AaJdN0yu6FlTkdAdjNhtdr8qd9eaZyPJb6Cw
vuwBGTUer1a2x+0hGhbZwSqaKS9kEpZox5iCBM3wv/L8kdSJm0vju4g+JRYpVQV7
8ldbuANnVLvOTeTjEcXY2HeJ3OmyMM/WKWSoGfQ3+J/go5bgQ6pqZpeK5CuBfVpS
p5vp+y6OQkqLJfR2G5ik9wXPJ2+3aYQRWiJl5C1mpY2pIbUvKpqzWZWwsgUD5wyU
BLwDAC/iTd/exGuGcxltRWZXORtTJWLYqBltyqJ4dAvsPhTUDFZRfuwcd/oc8cm8
NWMlVdqGcjDHfq5GDwYEWwb89WPAMZlne6yyYd8Mgpe+ifMq6n06QuxsaZineLJy
CdwPV5GQipkJliNSpt/nB2eUKCT4swJJSVRFiGNvBZCpoQzxqMrpl4Bn8YJUu7Ia
We/v+FCQV1bLhvT6j/OzmhwBijXxErTdKeuo31gJkptvhJvox4xLl2gSBeXA9Udc
WlbOhYKzp+MicPTKQhk6GWQIpgasphoOd28ejZTEQi4nDAyibgxZin4gH5nyJnOn
6+nxjOqZOB5SilLvQJ1GUQ2R+whXPVBmw/dKc5M92eKliXKsDtavluT0m12mF4SR
wbfXSquMSutqCpbAJbZZwSRMQA2dpA1CfQpMI9dSArjevbqQ1sWiYQXIUpYafMEx
5QlwsctUxlG8b2hYLvXLRTVTh/SwnIX0t0CEKZ1SOs6EvliCQXq7M17oFamxy65L
UBNcnuFJhCAI8IW4fncObsO7E40uEXLfOkE0sLdoq/FBPwu9lCAFBxY3hlIRwtWy
PmZOrXuLnC8O605POA9oXsBT+7AMEu0JRwz0IVQ4jBXA/eTBb30APqSZ7uUsauMD
kGqtNPSmIXxcqjsx14DuAKAu1cGSqgRSG5BMz03/JP0wQSVIiaAoejYylhrnydxu
XDNyaT8l0j33fSY4HteCYoXqxVKkXmpurPnnKqhDHbBHkhE2Sqxkf7BDvIJ2MzBm
V7lsiCU36ta1xctsnv+IGnjjtd3m2nb92MmDts0hQId65OeERfRhcx/9iV/smV4i
1/lxfawtpqtkoIlTY0zRWTQijbUe1YVsMzeGSD8nxLosNkGNwV+zHqHKBClJfmd8
cz8IEswCcHYi57cl9X2CkSBYKnGYWy2+suyRidusJFuXK3Wa5qdg8vTJr5bMLixL
NX1kSbfoXGH76sfRXsFORhtnMRko6p1xt8zbs2Zl721558rfcntCAwMzGNPShIqu
Ii2Z55xYCHLVaXLbCiwmInEkFD6EgNaJ43EeHbW4QeTq9THD3Rluy/UHwg8k0wRR
R1c1YUV+tgxiMuD2kXdHrnMIOYyCJNzGZLhojrxVliM8XySSxqtSaN/4a66I1wpY
oyORiFQAQWTBYE5LFgtZJBjAEZSa2XZV4r4IluYzg8hJffV0vJPaYYAZABgpEX9h
K76PoRpoIKNOq2k0TDUt7T+sxW7Ia4CPHpgxszZPlcQlFlEY39UmIpzGDWY5yqcl
I9tKCkwkh8ymfWL24hfoADdfIW9kF5dRYZdYRXspUJ/JNiRSyQqH4qEKeGdHrXLc
ir9FKfEsbZyYq26qvf6vhXHyFaprViUOpiBvNhF1nxgC12id3BuGf9JPRe8IHTIl
Ffx3IQqABA5B6WH9vskLyNLo99Xfk+vVN258bm1635ZzHBYBLZX8+K2DdBT+as+e
bhdQRwtl8tKQFDZGmPtbadEPL2O7t0fEsrslz62VAOxrcnNO0S0pEt83W6UeeSVw
YPflCA1l7L2+khJ3s1DaKmuOYpDyqm+bIzedoLfDxQxwufht3Wui4oTZMHl9+ccR
ciTfZV1xgNco6qOqkfTBVyRNLBTkb8/RV+z8nKrDTBdHy3YFrWr0f94hh/dQelAl
IhHHvFhlK4QguG2ZAXD9rpXoqeEpcIRSKyE/0zdsiFMu7DZg+Ckoe7AZX/j34GUj
ctf4lW7LQO9NBaCL2sY/wjy0ZdjORVgINGPS52Yl5LS/BwJp+wzuJRTxBY1+Brt1
nZAV5qMPnhPtoGNOyhNlWV0n7qITGzgh+IWG03ufaxCu2LNjS8ZWKTYoUpOoJLdZ
hkbg9TK1AhRffP4iU4asgHGE9HHkey1qdntdgpSXW6DZHtgMg+lBqoUS85ZdC+fI
1MfUPQ/kYUOqg0p/0fpi6353t68Fjw2pdO8dTKTcDEUpaD763MFjUhUQDzc/AUXN
IkTMdIjBI8X6PmfYvxCrzsiap1DSvs1p+jREj2K1TG934wSP7Sv+WE1wnqyH3NEB
1PsDQ6/1lVvKWfsuGog0jjAMVj8/4EhC7KUUKICeyaUAwUnDh1f/da260wnvRY4l
e4Bl45OdCUCjwecXWiJm5MVz5IkCskLsv+jTYrcxK+h1PG2QORtLh3MkIvZOH8ht
7B2/oh4g9vXc8OFDTS/NKujRNrhFbhCDPlDaxxUgrInqcTVvDZMFtSa+YFUlKVtL
VBJpdkl8ngYDlB88LF4GXYPPjT9ZYSsKvzNvF/7R/hcXIf665SFicVJYSGULUyAB
NyLdsowIYrSc0QAZgcEbdo9hyrLLTkkCgPRVNjS5ihojyiIdlsoVH1dAdh09t6zh
zyt1EKY9pKiqAU9480WD7sElT73sBdAit5iDROzg6kmPsGxhqrwYDnIw7dhDE7dc
paUZOU1qCY6nxim3lidhEKaj3xq22jYqNXipu5UuDNLBqwFMtDREymH7gbAaMpQC
9fvC92aLlGeroNzc3GQlWzoDAsYg008NBPXn5Lvo8X6Cu+43hSK0i46Rcg35o3w6
QiIGGN8B+ZNI4CEiBZIFNy7O0lP9uhNvXhXfhDTFc4NI1SQA7/Nj/tNLlpeHiRVF
aEU0jb62ywElyH+ugZiNg72g9ooQpgTi27VZLiCdQf5D7w3bpX9OpN66DVEUHV89
pklZB7Q2WyPzry6RyGH8rV04yGYid8Jpyfhwl7MVC+V0QCc6UO0A8dlJHc8rpeHK
ZkKYRb/P8yu8WFa63M0LkqccYo+vQXRo0ROkefc2TBlnO4G+qa7qufsuidjHaooc
jftkOOVvG1Y+onPK7zurnsnjh0cPy6g28NmYrdjgS2512Kv0pZdzUMwjxNKjMC50
mneYkNT2MYqZa9qKUTt/mGT/Uva8+fRIorRWFd09yCHQI8qO3PYuI2/M5u9Qlc9Y
0gXQ6XjvFudGN7/HWndTMP9MBRVikvlZ8b9saSur288dS6uuUKNWS12EWf+z0cx3
FEVE37SqVvoXUhgeumpNz1NngPqK8lzbdLP1C5SaJx+IAWHyDg8JXnpOxQX64zZA
9LFj1GLuzJof3x4zXFHDpNPfV3mNoAh2uzagvTocI+wjn+cIrcNsAnWQpEbvzdef
UnvsQt4bGt8P3DSTgSo8V0kGYlXN0dfxweizZyx/0Z2UqZQV86VfPvL1pXVbvWBm
CXJ/sK4HNQy4j8dZGaWgBgbDIjXi6UpE9tcle9gSgSqK9InT59m7BAFOyX0vli5p
nGRU0/AKo5gHdjDfi8Y4TxD65qYBY8JGu2tl3sozaB7HWK866CNfRTdDxFdYmLVW
Yj1ZAOT/pmFhpffGNmx47s8FqR8yAnt4B7rWiycZsF3LF7NFJ78CfrPYMAOVJBwZ
tU8eFiSW/Q448F/LAdEMqVoTOsUcYiSFkYNgJEAHFZvAIG4s0vN1TsAL2/hncoto
PPJXh+y4+GDEClLFWXjTc/vc3/ufpWjwG6LDmmREvepLLUACcAG/35KiDoisz75Q
K5dyVabWxaj8lUK56DmNi9WQZ2BUiM0yRw4j8gptecwnyoO2AsHQx94JCIdHIoKb
1+ENiXvokpLYqGTMvo8uBOZr8FfYVOAqtIHMFDJ+lJP2ZVOhL/DVHFInrYLTDluE
H/rBCrNVYcoOQRlxDiOzWP5rtJYPUqGXdZo6dpreA+v3JsY7GRKK1BPchNb3O56w
oWBYGaxXm0q5gQcRCTPEmiO9Kut9w2Tz83/ztoYAxsTtwt+6SAHNdskrA1GBOq7U
in+slXB+9mB0aEpwuPHE9Qn7ZaOUHgPRossYxuSIra82EYr6QtZTXC1OEofM/2wz
ETO7RrdlD3+iJd3SW/B/IBJNzTOF/fXc+eRRdB9oItAVwXwi2FAM/5RdShXwigRp
Cr1lkYUpP8c0Nna88gDEDe5J7EhNnZ2bbLmVHJF31bT8vDkYecP2awTRzzmbJGUt
SxbkXLQffdGp9ZlbbhK16vIcu0dbA3/xxxitsK3y50tPtFHBLvTIqZC1PZenuZv3
nURB/7HlvxkZV7LnLrGEy19WyF8Jwgro8sRAaZkvEl1zVy8Y6CbcIkO5Oi+tcRg1
Oam6A/BUcyPEOZrAc4JLc+298ZuMbm45GoRPpOXdJHrY1YwOV5QWDgcxveTMU2Ci
ulq5xEpD6LRRJGWIUhMGl50atLG4Lhw23TbCylHndu1avcFCQJ5B/3N0KXK2LqaC
WmDKUPryM5zzpSm7hymNhWgx8gI57wSUN6Kf2fRDLuPOxi/+SHzscmqEYNOqCWjl
5rbueWEXhpyx7opPXE23LY+IBxnIGc8KPYDA04l8r2Jlyn+9deCnJiV5IYIOWj57
sKA2RMFlFqRl9DJS62Vi4IfiN4KmohjO2Ix11UdcXt53EOsTVirIjvyvC5cYXnHW
/pwQzWXlWSPSu5A3OGtVZOgIg/WmLdfdC3ZRf6I3O4Wjw5KCtyk26KKWmgdb814W
C+AIvidLnjHInvWM/RyJ05JHjHeJYOezMCCeGqamsJO04zJGMjoq8w/aqLncxuL2
uzrR8VjlksYmuxqIXCinNDGFwCAeEYBtVcMqHP9KXuQL0zSvRcQOiIZybls4dXLG
4iCvOY4dIataVPLm8XjIL8tnJ3/+kNYSXS6d2j7/aID469QFgc3mwFMBhHulmrbG
s6njWhMFVvlPjoiG23AZ/6oaHzG+uqom+5bV3euLPImG8lz+/kQj3jzXIypgkDMV
ZoSFPUiaBJ7nrdUGaDlva+dvhKPvcJUTgQBRSIisspcqj09w2AGJExIDw+h8OwS6
YGJQtpovj1O+3k29QToyzyv8f3/q2d3GXomaxCEdXnSCrVo4W9jHc/lwMLF1r9zI
t28fj32ZrYEbGzVj1BCvUrtlb+3Htpm1hHoz3P4LqQgTuDD5p0PwQl1WqQmS9hcy
e3xY29cGdmhULmcetQymXK8InXdAPmzwd4iBX5aP9xWSoGrYQ734OVaPrfEhq3Uo
LyJgzuYHlr+0xR1BtvzPXF0NhwVo06W1VRRGV6VwpZ4RBxjlQGEZGIS0ZzpRAKkb
wiInC/7vIrf2qtpt70Hz99/4pTLzNHk97QUOLrctWVfG0HV1toAWBWJTUvTaq7aN
Rrtc3Pp8wN+5f9q7rSlNezRc6s5tTqb7F6+MXNIlgnzWYnOW/d/Y+z/ZM5EtGJNO
D/m3wRE2qvebVc7xcYM9f066x1je9/JH/WM8wepR63am55Yr4XpOzq+XqHBObEeQ
HGVpldcDQn/hoeDWxTyrvbrSPiY2C//TQ2We8EEK0ZtaloQvtLtDSwvpdu1DC2id
woFwbsoJ3TAPQksoQM14ndCuaFmM1gm2VIqdzTW2s9BUx69wGK1HsEQDqsK766Eb
ke1KvhQ5i9cgrRczZcM4TS/aJE2GKauTrNTeSZ6mo5zWwy7CRT8Jwq04RqCoOJFt
ZT+kmJ+dILnOpFjVKMT5qtsVYoCLHN4Vejngm/gh9CFw6holmjI1t+14y1KeuXDV
zFTzjh2oNH9a37Nm21nmpLcBrHlNBppA6BCFF8N50V+xSlVBX3Wgl2kjR6P82qcw
7XBud4TgJeZrhN40/HQyK2NutrOcNHbEIwfqEMbkntIWve9P8Cp2uPCoXyTZMlVo
JP/fL3D43QAh83B41xtEviZq76QyRbpAw5/qYz1jlIOV8i+Gldcdeohp6/WVvsOi
Aq+CKPfcgWo0Zi10OtZoIANFdemzwg0OCSq+Uget79pk6xZwxK8TH9wEcXYy//s+
0xXRNJt/om6BNthnWIRfLz5Gpa3Wf/WoVM0t+c7SxjQP4XvdAYP8I7fDjsRmeYFn
WTINhIUyZx1Oca75PBlsesfXPo1i7c/C8SiWZCX27iB6313CsDsO35fzJ+c3GnfX
GTTFykAJUUihAtFIXre2F3mD1PdO9CmuBowzKQOiuSBLpPr9sgxuspg3XKr7FTYe
lHZrirPGIcwd+J0QrQrp9vxseyQL30jqkP5tb2OGWl0Wjq6aGfTMp2T3eBCl98Dc
ayDorLnDtF37JjqEQsJfczOlgPMoOUYmHRbBtvvRX5usnTcNs7ZCZp3PyoAjUKls
RfcjjnvoANpe3+nze7SEAlK/GVdrhMJXmeJiV03zd6CUWjlWTdFP7OmdxIdp+OBe
mY+4DJen3KhNlxuWj2jGGPELeIsqQRtygyJf5CkgQ++ergy8rYYlUzEZZqpIKRjz
04vTk3aMsv5HNrhudajCn/e/LWEk5ACzFADpez0bFbkp4CbQH/j+EELvDtAfdh8u
rj7LfRa8EtvjMqs3pegF7Vg5GLFPcyOl9BEJz6NnNti/Edbr6kBvb4WqVTC0ibhe
ABHaR3sQU+f/I0tWYIYKif6Na4PJgLFnAPmuf9XkcV/n+CffT2ZXrTwIchiorl49
SfyfpVhm0b/PihyxM/+4U5OQs8MeY86T4FyZ8/JaAQtALfucfZPa5UHzL+NOn6Oj
tM4R4aC5xSsrwjCfE52Wn5RyINLrYfluHAWW2VnmYGX2p1xPUXyopHJmQTObdOLF
5V/TC9Xp8C/Addncf4EWe0tCzG+FGSYjVXUW7mUuAsPh4k/HNSwcBAitdhQoXUYE
uq/0zNEazpAaPQAmlX8qNn85vAJjV5tu622XN2sFh3Jp3HyjEWEm09MoXTxH/3+G
M7WL7z1SNMh7l4TgXugbA6M81FiA7JcEg69tbPbWjovzoBOdzxjK/cdr0gcC1Hsx
yCBbKUisHqBl4JHy6kA+pDDUfkgr2Y+lS7oVDbufPD8cuo1nBVz6yU/K53LuNafI
gWi9sRwEnahKDI/ZTSdkewaC1vK9DqrAJpvXmheDToyoL5e61M9WLkmZRb+Bl0WL
wW/AEzbeSuPvtM4DJI3C2EJJsCx7fWzt7Y0++zbLygCL3Nq1A/AAK/jODruw9jPG
LzBI0ndc0CqrURVUJrtvXq+A1u//NMNDPf7dMM8UE25btVJPpDTQvwMbNl3+q2wi
A8uYICvG4Acpi60FIMmvlzwhMZZQwOLVcqBigJDq1jl4smeR/m7xNQ74XCSWfo7Y
wA/IG0WTeCHwqcJDvIn0F9ZlHobRSCnDXApkN01Zq4fJC+dxeSTFcKSOz03IgW8z
P4B4C5ouPwmbiq3oJSVdzci+AJnLqk210um7F7vg2y6ppETQj7uqYeUWGWn14lDV
t3VCO1EhksP8UaN1zgLVgWbWQB8gqx9OOrXwulZfl/pBQ33uXX0Xn3HQmTRmC3P6
44WnLTmaCqPC+vUhgGin1eEqYxPsL2a4rPTGkEb/VMBWAMm4gvQkEKVhqh2DuC20
B1aLysrhNVMzbVb9C8J2Ct4pVrX1sR7mLGHPP8rTkuuGhNJHHdieVS9K6qpgs/lD
VdU4Keqznoa/hzESBnIqGbMaBwafIh0BkNFWoiZa9Z5D1pi1CCk+ep4iwFTmRhQl
tnAk3mIssFRVC0zkfyJuS2cxITkZqB4YXesBX4MMvlqCEvuAPSxl2FkOST7b6mqV
OnuHItAtsPqZRhZEw2dx5DA5K/tU4NQCtduKzhmRplXJyx1ZG7ohsNW7taiJDtHF
JTqARXp0STPTPSRvHgv827x0nMMHwWEwt+leLPdaogSqOwnJVcP7d+3UCJMNrwmy
bmn+7ydiCV4KXBMye0HJAZPi3FCdvi4FRFsWVpIsExVEJeuiOAK3mochuKhPkfJP
GyRrOvj+I9A1im6kpljMqizDuWxe2FBOFv6+CJnIUX0VZTBVZ7HFWY3SZROuhMJH
tuTj4BpYonu3HX9ogovLgvpC8IB361Ak/VgVtR/YWwkzzRk7EVD4CCZ1vRH/faOi
I89zxT7uYFSGCdLmcxLClXWC47WXTHkDXyJaMumbNTI132IIwXwK/Te7hNrp0tSQ
a/ZGLv5TwDrhoFevIWnaCdxxN+kUrOZVw1zLHsF6ofska2lKeKESsk7k1M5ZKRJG
RvIGlNvOJ+aT+F7hg0f8jTG46KiKQw9C4xL8jlXv0Eg2DRT4+9NNtaBx5b9bBR+n
MQ9Sg0oVJglWSmDkSaQNpc4aDongIuLf6phfWjGb8UsN6humjDOzkjkRylZLh2XM
zqCxzkc+e9IHcmZrZyKxVBxpwvCgZBh1HpYKYVSLEYIaQYsBysG6AQIrFwnLu3LW
bcDZnrr4MTeiFp/klo824ed96R1tHd1ha4EgBCkqzgXcYjxlF+qe8VoshRIRnq9m
sJQ1FWq13UK9AuDukBWwA0HpK2DxtU+cEdgzGJoz34q1jlQhDR3sIQZ0ZAPQg0Ut
w1kdSs9SFvv46x8MFtSs4dsdEoKgXffjulxX4Aqtg2dHi/c6RdVyHGWmEo5nslS4
jfrhskS4aN0PFYBjToyBH3S3Sco33YV2Jl8bUkE4ueMHLh2oJKFpNuNLUTjgB3CT
E6slHzk5xgjH0WvZQM4/Cc9RuKOrKZlOLEF8vHkaCVVf8OMHEJp9TXvx5PlINyqU
rdQQiat2vd9iPTwm7HpF+NyN3AC+SvfOwAeqPNbCQ9kgju7n148GWQv5+geAmgd+
35ZosRuaPocq2ffKaZSHxTp9OIOOqKBuHqvMJy5JFi+GtiovoWdcMTazBENntfzL
j61zQnb6mzyBtRZGcLxIzsrTOUT1w3IaQTTIMjLcUWg4mmZgrlIgJWZZZhBhWYtH
6Gkkk+Y/hht/6y8sGYL6io824SlRiYYqNphh3SciHz30ryaf7loe/4edcclIYx/F
Jkm+83+11YjmOewpFPKKEa6urfT9FM8iwCc4rMxsRMm+S7K00TcbrJ07sLHMnaHa
fQfsEPkD+tSFSe4Jb1M+LXSVdVhqfMP2asP/m7bUoeZytLN3mN2F6LO3jK/LeXSn
n3sd/m5OUqe9aSOiUcqh1K2K5K2XG4GV0YG4ecWmGtdW04pG1EVn5MWPamEopphM
mz3z1Nom8XEAx+khb4kfl+GQBKqVOg4mELYeeE34LV3o5iaWp0VYXD6wys4EBiYF
clWA2E3lS/Bk6zLDAkdDQUeCP+1wAF01sADR5n0Q4vVyPLBSVo3u16VCUwp19Obq
k6I8Amy+9YShV3zJcK2o+zN/0TsHjNELTQVtaTrE0+g+FdM+wuC9Fl/wsnBjz8if
KkP/PBge0LTOgQib8NaLYfzTsQTZHLwlpUXwtseKTCM51elSh9hMIbxooNZe64aT
/DP1RuKeK0meEZVsfQMWrhqHWxqKT5CxulzW/sN7+fa0IEGkl67/H1r+TsGD8N7i
sPmDxW1bFS0esseVtLoKbz5PTXrIZ7fsZ0UtsT+NtYX9kWnE+L/HRsFvgeueVusn
PkjWEq92VeVKanhybgGdKCwzUlqfrioFsz9xbIbIqb3qcR5YCbDvKUCI3B0Ir925
RhoznUdxkR9JIkh0O5La+mdPWsTqXk0McUMFtdawjkLUclnc8+W7q+Et3IYYYepw
LpUgrcHh3Dbi2yOsCYWk5u4ld1d/ylJo7oUTvR2/A9CukyZuBSuTt70lR8CZaZPp
obJ8025rbURognMLKojth4T0K4o0XibyiqpE7Dsz7i0i6b04tN1PctXTXWky8a04
WSQwZcDeDJQJ9ktHmTaY6biIS11DOqA4gfTuPwfNhJHCGyqCvCuUTwOFuSJ49XSL
0e1Vm7Ib+rGOuEjAcQ3Vy/oxx8JlTw0o1jDT68vfG93N6AUGpBkfpA8bD9gYzoDR
+LJ3G/N28klKNOwixhpjjH26zQoMFSnLtY42VLYbkaEiveYQ1/GvMlMihKX2E1tB
SmO/njDuJUdR/Wsyzz3AaDA9y76aSAMLVIyGJ0kj56r136Pbzg8f8hjuw7nSqMqL
nrh7mSIrv8T3iYUtiX+uKlucl9J77zxlICZKfrpxLhaYXR/5rX6icD7Md/L4byi5
4Bz1z9hRAl1uoHaDYGRzi8nkFnIzjB+i29BW0TeUAxFGkpAG3/xt9xlBgZQO85++
hCiHFFfWPP2peR/Db1FmFKvRTSshs0VxGfaTWscXWoZcISwwCCsC6QarSAQ3c//T
m5IjR8KAR6REkwLemTrVXfkm1sG1Z5RCi9MaBn5gs0ATZfHAl3nazojGzU66D9Ps
EY1l+huBqTyISSZeQ4e9nl8xZwPjkijSYJHULonI2N0I4xJxfP8RP9beWkgwUtpr
7TFvl4VHg6h55A2lo5Z7TMbCLKQqyn7SAeF4+JF/S8oiLNiFFE+34ynrMMSKm2xV
1H3dFJ1rWBbgFqVuHlCJFzJdfbn3wSsRYE1PSSXQHQCn4whgp9A2Pl9Vl+DDYcJ7
2+qfpnOCBjV9F3KnVnXoLjZS7y9v41BKbsxZ9W2L490EKl3ulLQN6oTzE81TuVzX
FPXD3GTuOHSM6oZSn1vlwP5p/jMMxeSKlhgXwvqJ9TWTl8m2cRB1Hn41ANrbT/XL
IJFfU9edPjtOvLMI/Ocjgf8nFACleQ5s0Hf3TXJtBxpOMrfHPV37iEWLBbgvx4gy
NaLtk0DmOE0bmQnzbA17baBI8ovzW/2/2P020ouQMOUhaLtkbZrX8Kq6ApHwyuQQ
rFkfvX1fAHAa5V3BRV42KCTp+8mb2ziDs+ahQnbmNz999CBTKnOlTHBU3C6cdcAv
1hRHE1I8YphoRGQXDMJ2B+4PnQQsxbKc0uA4BIKNSLQzvIORBvcikAwiSvQ4A3+t
PtZvhW3xvS3OsmLv6wnDdZeUXjGZBUotnEgD95Mnbi6SrcCi377MQ5VFQ+8jEAGs
Q/lwurM0FCuJFeN5ces3fILRbBFT2Bg8wiIkroZLYy9EnWlqIpsi7W+HP9KMM8WK
IEzQfa7cPAaxV7tD2Q/bSWFQrupxkfio8DCk+pqYi+fNfNPQUqpTFiU9aAeEErGL
BiZqfNb3sc6zey2U8IIYifBACRY+ihfzG1Hq4ctmiOX0UU9oFMGTMpeWkduDLdsw
WO2RhPGpPjCwmeSwrdGRcWGNKgLEUzNZio9bTDAuwdwWIJM0H/xDrfQB9SknyCTk
6aoQfThXZZc3KtqZkH5gWJyAWHRGhNqfbkfZXVRXc5TwQEvxyjvd8FPyKyrc3L6B
X3xT+QYtT4u5YY77pj8qzgamvNph+p3KRJU6JdMdhqQxTnynRXpJlFEds/yzb/Nk
cfrYzw8YQuWBSR1QCfyjd2FmW3pkKccRZ1HyOeqBgbr10AjRjnUIEW3VWCDx6yCQ
//W95BB/fZJSyOOfsKzYQndxm1lDcXroyvYnFqCpakRhsiNAkU1Iy66C57R6cMvu
85VvFt66wjmJdFmiMVJgiEhdA74r5STS+5pre5zZJa2PPhmdpHn0CkyLnZ8SSk7V
+kPWDjKVYQbDIMif6YOyzSsZyAxG3sOyUfmID2iY5KrcNog487Ye/moQuAx2esu0
86kI6SUPiTKNZkKMV7VmLlDU/6/c709EBKMXOL92rNAmXdpdqadeFPiu6qYo4X4I
PLf7egR2YY+wMnF573Z9dAdHZPqxLrdIcsAlDLOSwtfkQDbcBt84vjn0/Veszn+N
Qzc8RbCh0/3xn2nDtCQ61fpVs5NOMFQY7Zv6+2ujp2n01Frgii8afk5xy76A9cg0
3GQOe6kbRQxSV6PL0pjZ+x8v4jsAo2zgOuvliYgP2fA0kwuLbWcxgpl5HKk6TxpT
s0YI5elYmJQOFy/1LSFg6nw1bvnSBmk9ie+iHOKEe0MMg6eQ2KYncHhj5E/PNkV6
TUid1yo4Kqf3vh1gVRd5S2zkwfO22VjePGa/drDAJFg4PFIhv/c9QStM4s5Z2dDm
RM6AmvbD0dvVlLftxj+r+I46SirXCzT5040xlgZLxGQoQU1s9CST2trGb1UPCuVG
L28PRlw4Ohhh1tv1COmuTipQqsrGABr1UlnwYO4LN9CiY3xjLCK6qOn+pdID7tzJ
RFj4V9YHgGkhGv81b+gA+bEsr75vFMISBFjRxfLXnGA72+aI3DVDHq88Q6Ss09z8
6HLuG25ClCl3L5G/e8LhI3X6x2YIrM8ZF+6Bl2fBbiuSv9xdtv4uh2MbPhIUoO6w
0APSGiNo0jPQJVkrSOmvswbaHhPP/ZIiqGQilpSQ1nnwZI3U+p3h6o7cxjtBIV5d
H5IIWgmfpp+QZVkdBBtuwH2AlDDKKgrVFO/TIgcjcQCLIPylVspmaiCfY8wgsHEf
059qrh6qzr+LOf2Ii3i/i9a3tmywAL+Rtvk6+h12FkWr6l+DVDIlXZpYrFhVeT32
igDCmkN5JE0iUZ4nfX1FgtHzamXsYUSzIc2KNLdF0HRNMti0HAPy1c5yITEJwy3S
oUxSi//cqYhSZBjFnKHPUsG1tBzkga/jb7YX+SgcNMoPJtHssrJXBoKK3QNyKcwN
WEMQVu764dwBRcy3DyOLajzBrimWg5bUk1kpddkF5mfTMQLjlPQa2JevD2HTrheT
seNTP8DCWkrLTWaElbLYMPG+2JEzHCIItOwWldVNoJ51CNz+4NAILKvDjUSqPh9V
RkVlZvHzmRk5x1gqA9aaoxTJq8F1l3WR5WmUcKPDBH2Xra4E5Ry0VxiRQ7Qc1ZjP
HM0Kcvce0++Y7f12zS/fct5mIr5BuBn/JblZt2efWcCaqSuY0nwtgnBox7TFI5iU
QzlqF38LgYuVT2VxNuKpgw3ZOt3nFGbKBrYKtCSK/py9A7jEkHOnjOzrvLzq8dQV
oLb0THgws86rDWMsY4/MVm5s3nzII6eiSKP6J5jleSwiFicLXXYrNvShxX2EoJnG
MpIIkjZVTLWXNHQrW48f/EoQNj9/OZV+GXivH57qLTZe5YtTziyaVMK//teUvjo7
5V8QA/KNwTlnP3oygA+PqKjYFS0r+3tEOJ+58VxAbQW1A5Wb8qEQGRsuksFT9wHE
xvRc+3jlMnvgrosCC2otGJh6H/BDeQVUEja47KXGRTGq8hay0fuxWJeLev0gFrNG
CjVbEjBeWB08nXCdzDzhRri0hU1I+xj/erj6s3KC8iu0LdIQS/Lnv/Y5oQUCJhbq
n8ql5+/uApb2doutLOHZgExoeVbHrMtTH9U1hR1+epfQG9HoyIhGtU09i2yukmvO
5MYFf6N2wCg+bobc3VpiAyv8qoIqXGKLcmzeb4pViq+qSZUvo1MesYGCCMLLezP/
CmTOJQ4yT3yGXI9EZHDUwTne7mSP/CnjczG68kDG7NS7rnFsRq/1rYKMBq0Jr677
872le+O2//ZaKpO3Aa6M7/n14qqSINLLzXFYpVoLv3x5Rr+ZgeTYG6d84sKta532
uA1XT0u/AAPTKKIAITWdMTvxVNWPKf78EGmvUy+vkwVEKvpZ26oHlTqYMtbE3LN1
w05D+X32176ET2XZvarRwFAVCDc0KnDGs6d9EovTsQBL2C8OEATi4TCSL6m5wudU
jPKQgiKTJqR883JeB5sdAXqSzQu6ZsHJ4o3IXepS1cVf9qryvlIo4NDAoI4pJQkq
BXUDZCti1pRh0CIg1Qauin3MhS+zf1If/i/2eHRWMOw/oHut3X82k5Zw/uVdnpDW
8r9TB119QB/SIIHgIZyqXMw2FNxw3CdiQQ768QcIJi4d6CPtCgJczVa7afsJ6qsp
fNs3DRdLM5hLHMxZRMLN2AHbVbkdx0/d6FHcIPP/PDyenXHXHFGjZtmDVycbdn1z
XGW5iZYDdCforlVTEJ/HOyZn7P7WQ4pnJlQaMV4yHuqPeeswcyinSIb27MLUpGft
36kmYvNVm3Yqn/HEOx9qsP+IrQ55QQotqkc5sob57yXYoFMg1D9AIvK01XJHHbG6
L38/NILlgv6+Oq9/dt3GIUOajQbwjw+uAl3q4ihXgVLZG6Za+tzMdt5Sb1q467G6
qGxWkjDdGaNePQhLKFBMeGqXmC8x+i1Uy5Br+UqH7PLwkMl9F4nl9WLVA0ta29fo
krtNxYWXYm+h75Y5QLIcHaLEGGVOj+oFloBBol7NGLZtOk4qPY6ZFWvqsefktxqY
rnI03I1icfjxDkPHt0+4eKUGc2ZspZ0iHepX87UnDkWoT/6JRNzOv8XUlJgVlDuz
V8iopsQk/tAWplXw9HsvnjDkwK1S9rsCnEJgKAP5bmx7RAHH6wYRdFgLa6Cif+u3
hglP3D/U0iEImw0dQlJ4JBE0WvndRzNndhGDQSsya1+RuW1IBipHk9VbVuivqgSY
HoXDFnhFoqOkxFGx/MAsEJyNU4JF0tSLte03dKButQ7mag7l8Z+C0AwKUHej4fTZ
eaHeiK/0dlolbNTjqsZWglosDCQX474yZ9vl9NLX9iZRhaROUuLypSpgylQTjD6U
mNLo9NqNUcSr6sWJ6A6iGk6Okqb0O7MbuRiZ2qemWFxzKUxy8g/XRm/cueanpwQJ
UF4n3tCG+8PiCpCf+BS4eHbyN/0V4wxJPm9ubSghQuqZQtSQXKWHUDNSykWCtUzG
woqVZItKNkWKz19ZSFm+27xOubscvNAFGxFQN4RUzFOhVYvTC/qoa14qlDVrXfYv
WSLmVPPLQYKLiDtlBZ/06PH9njEi1LFwDoyaXNbEaQulDluF34cupxluqGwHl4Z7
bjTtbyZEMaG0l3RUCWLJnqEI/EnjIx6SFUGkvtrG8e0j1jkr8jRhf871Q0lV7KOo
6OLs3ttNrzfFCcyyF38wnIETxh1OFo8RUdqIS4xJ8qP/cJ6QQ4nzm/xsessCmtio
AB9zi1u5RXv1mP1XZg49Fhnx0Ckff3JSksz12ffluohsO9fMSDZxx6abkxqfWrO8
HezdpxtrnvLafP5ih+WAROeshrFGEWKyyXBo12tT89UWELOPoNeIWRwIwIHiL3rg
gSzFaEcBW6B7MlekmuSmtbhpvjGuE6qwzvLOxgwaObYL3EqEJCI7ont6nz9wZgyg
l27sWHKD+qM3XMWG7mOWcPTvUll8VlTe9K1NrUxqKaJMuWx/APfjhG2H2OQNpUfy
rpNF0dKihfP8kVAxCQDqZM+D4AkK0RZW2GiSm2TojDoh9zf5pSxs58Uscfvn7zhO
dZcN+EQdk7R8o3SL/P8HB0EWxlY1yk5dI6foEvYVvLltigAt/tI+Y7O5ro3ttXyj
Vxe+t7K+CXRl7POaz8Feo88qtiN7yykoE38CTIDzRAqa50wa0IWIyzDKu3HBdOPR
q9gdKJ+PwWsTDBhVH8M4B2d5hVf3I2R1XjJzcW9wBY2qOdyakhEHltWXzIECBmi9
XIlRBJk5dEth6mUk/zyj6x9qxrAh+h4+Smi/M0mddeIScFTlF2Lxg04u6WRAcaEb
R1zM13vbzkIFMFX7mxcaWacPqcK1Ql4gIccd5C1kiOwiRfddMli5tu97AcyO7759
F1FvX6vRRMDW22L/6YBVEocvFIwCYiaQBGwov4NuaxXSUJNC5HP/A2vzroKzGgtL
fTo1K0uHIGFcve3JcFkHq+f98X1gBhw0sQS06FejnbQvlnpBZ+fhXzeGGfskUCkY
x/cPnzZSEa4npJip2efvKp6jU9a25/grw+NZkix8I7SPIHjCYGJeFrardEdutD2W
Xjxudd3n4e1CWr10bLq4RdPObJEoh+F3fbq6xmHaXNuET60gOJ3TMSNsnGV4mH/S
ubOBMgCD6XC5wMP4WRgsrw5r9TnSXOuLYV/22xWj9gJiPAvT2qvNwmd86orl6avA
1AAux7xeQdxDWJZWiYTk3qNb6k9svD7+kDzRoAsfO83YbDVbUb16fh+IlYy7YLM2
wHfrxsgoQ7fTHrZAlLgLXDSl/+Pd7gPaiMT1Yu0HDDBbww6ddiZO07qdnIwG2+fd
5BY2fNd/ZxIq/y4BY7CURlxZWCtcaK3w+q9oW2Iee8M9EbhhdLaqfYl2V6y3VzCZ
Cg7Rr/UE+0tSrj69MzDWEG+VQquoefHoQYwZIhqNTeDSNcfcO+5OshT+7WM8Tx1S
Bh8Dvt65QkCCf790MJfazChyMP4nhIwm74c1riR21X4+yjEFM+pO7lUAhSR3XLXh
TCyktj89hlOEfcotiOWijA63uL2/l1sCemmTXffOAjlEMYPDzIuc5Rl3mLUJD9WI
iXGUfK6RJOqCpWelMCdirC5T2Cvw3VkdUu3qEqnZfRO9GALFbiynuU8JfEoByTuo
j9+i0/CuApsmjXaAW7NEWfKIPdCnLy++/GxYrrEnvC8MUETqhMbSUcQDy/v+2OoX
/MD6vP9+98/vdygVypItZAuGf9tCvgLcCQ57M7lCIYDTi/LNQ8SQf4JF9j9zRWcy
G5hbrgGkTk99jiKIaWt0iZ/p0A8GvGBh22joQbLnhpIDX/0MsuaLR8YxwWGyAxx5
rQOJm4pRSA2DMWMdf5K7xktFa2WiAuiDFGw34aX3NzE2s7f+4fuAcYz96O7RnpYU
JZ8pIoSHMsB+YahXab4DtEu0hNKUyX1jGCYaBy8N7re3duA0VYoKJnd0DvFXxcrx
CgJWk6Wrzz6vXftlY3bCTFTRWJwGclStYh6mtvb60Z8b+wX637pf2LEDCh/Yt88+
E1PQPZT8uz7D42Ccal3KoLPUHZgLFoPQuf86/z+cI/+CA+7z5kRSwl/CeiV3ksF6
vbze1wxHSsnOZwD86kMDItweGfWW/8Wpzz1XeBop6BUnm8kv0WLoiXiY3pTC3G0p
0AkmZfQ6e4Bk9trEAsiQ5YId5TYWdCHt1azPIkx1pVvzFZrr71/uSMSp6fQV30JH
1UNWKZ8fNIWfbN7AtJLJz19p7OmEqmE2O/fVg+PHE7CpZqc/j2C1VkYhh9ONbWUS
l8KC0i3gL821WKR06hSDq38zDIs/nvF0JV6j2ysO3A7iROM9JUrgecziEOFCgByd
bqmQYSzx2aqHouH7L09dOz4hnLshLpyOatrbwpIapMLbwLujSgp9SHEYtUY/cjg8
nhhDI64lasoBhGViuP3Nwv09MDlS42E1HY95ToEpT2Y3aLoT8lyAXPZFXU7fE+oT
IHr+AqF1zULdrVgBoRVj37lcVPOgMfWLPvN/90jmwVM2oAmSuCI19nq/XUJUuj/Y
PzOtUdLDBbo+tns+KUlH41SYTkT2zWVOexFxNTge50fpR52qtex8FYqxlR9l7cQo
yY32Yzis66gTCcbi6Sf5PsjMcnSv5CJqTN4nwWWl4O2Fk5zkYXiY718nfFp0GVzA
k46pzL9N/VCiey+OU0wXvGZDnV42ANHy6woxH7KzlOClkKVmkEe3RXM8fF5L2T+s
hII9KmKwz5jKT9nTy5FgQ5NK9bDmpZ5FFs5srLhHFfVroKk5jSsZM8v0Sc716fQC
VfUql9lXPHF4gD5yt7SYTc+9B9AdudLGWscjaU1DZCn7THAyuPnNNFp7Iqemy6iA
TWz2eAfwJMon4A+asPZJydcNL0MyKUHgDZ9voUNjlFlTIoBpISX+O4zubRG+IdgF
Tfb9HrhKZD7EFrBjmZTC3kIeTLyMIs17pCXdS26Q/2HCWXcU4wcyNTvc2vIxd8BA
6yqaOl9BccHeTncLpIFZD4LfVvn1spe28uG5n9SONraH8fBV5dYVdW5EyQbz9q4S
4mpq0LQFhfGrBegNVDbJDmCMMo8WTrA5QTGc0GHZ3ISNMAlPEJBng+EktwdVdhfQ
A4Kx/72QARLmZPR1w3P+BBejm0IXm5a5evvpHRUUDiPGprKCeHyJOR2zp2nECuNv
hv329pQMsz2XKUXO8cYKhEeD7RrHoospPie7tfRPnuGqWBPPbL0KWEDb7anAtVO/
cy+0ZN0L/k5EfVDpp3ZPsyKn2u5dGvqKlYDHzBRXr6JZfB1MRVnJBBrzueSo+GRM
ny9LvtxNluTYni2RoQs0ipH4UYiujeiWGmZpWqrB9E/1d6jcsx6BQGSUQgxWg4cY
cFB/w+SrM6Uty7EbyTZQmlmXm/TUwe7LkN9cBw9oNx95to79z7i0O6rQrHUpXVFU
MZ188chHIp5lCMwAJUJ4xm0m1TtZ2mUVcAcC7tzPPyAKhBpBKuEUVPW/6sChpALQ
M6jSiKqdKjCIxRFgY58KG6ENZI0RSTk/EWjQxNZo7lzV4WTUlc4bkFk1if9SI/SL
4EKpBmlwLj+o8vkPPxPqD43xuNDmpmM/M5ctNYsb9L5/GzabyJzd87rzQzqP3rNy
6rDuGIAuTWQwoHWGX5mRJZ0j6SiyXoxW5nHcEQjWyyIPtk2VYpWU3OK9+YP2Qea8
GRY+9g0V66LEQPJak3hrGhNQzyef/dsej0sRA2ju/mFwrBYUmGgomnQRlJz+jsok
DOYTIq2mkAq20ZFcMa9YhkuelKEQi8rcvH8Quon0ufR2N8C1eKaloOFZsr9asdaQ
tJJox6y4R44bBfcAIDw9kKeRYiP3PX4njWNTAX2uz4c0qTPcs8ZojkgfLraZUe1c
cCKsIlWkM44jpaGanIx6aZbF2hym7Fydor6NRiTmBFniDf/c/+xFV5cdSCmmVuM6
Mrf1lPi7egNn0r539c/olC7YCAJLXXv+3Ju70J30Dnxhu+7Nc5SOhNysgffxsvPk
HWvNbuC8PusgtRj8iQLCI+p+HWtUlOMjTEHM9FxF4HZ44l5l57QsmKE2BDlmzSlq
8r34+Xhseycl1lIlRLX6ady0T7MRIKUwVwroHsnK56RldNd5Ils7s0gMl/lCSEe3
ix7bR2ezyGK670ydA3rU1j0Xqev9c2wyG1+X9QXxdyS6xxjIBLTVYUqBOheL2cva
3O1MepEhVnki1V5QIJAhbmXtcb9z/l5/sfZ9s7wMgDwAlSZoH+vSOOYBrY1X+cUX
KHpAnG+3/DOJVbd2UY6Y5YIyNkz17I1SIAAgbENJOxGHdtmtYXb+g2nfiG6LBFF5
uo1i87s8y6RreOOZvGd/gzIHGVpBs2I5PaJqYPMhYogoVBpRkM0eTqaI8nY+l4t4
qxHAdVVpZXCRER4GI+qO7rzTZZKc5YntwuJWnpaLVgM7EUst/Q1SB3dhH4sNsH1p
WjNdXbOmT8RtAJvzSRMqECbYFW7HQ0KJK+nr9oQCMsvrfja8oaA1X9ljl4QR1PHc
7U6hsQDwfz8uzzDdUeJfGaqGS4d2fo7b3dvoyEwGX2eN+JOipa9aQ6MG7iElb/9S
36oKuXBEXSbqcZIwIP/5ceSprRdmbI5JPjUYLNqPHNPUuKAQ5Xk9wOG4/otQPM5a
7J+vJxRr9zQPx7mRJ3CEj/iGF5vXjOJxyGmdZN7JM2KKTJ/nralcD5nDTRtaQCgT
0JkbOw6vwJoQQ1a6oc2xfvdsOqYdFd5gFWEmBA75jYUOTdRqbpYG1EqaOyIE3hT+
IgG/w4Hdc3l3P1lLZobav3cL14N+WcY9mE77mGxrxg0sFxx9NyqXmnXjoCF0pdME
sf1Pl2royY4h53QJH9HI6+EoR25DpLW83j8LMtB1ZGo+15NoHa7KK9qq2aXxbiII
DIbhCxE/+21T0cGUuPLKlTwjc0kt4ky5RzCggoHcts8GmZBe4WABcOZMDXG1+31r
Vkl5GukXfdcaIqjbuyE1pnmJTLzZtwQAjwgyZqtGT15zGg8KrwWtoyxvMtMmXS70
HxXBm7VcaYCVdnhfCK+6HYnbg63ZX0Vug7st50n5R1Z1uN7rh7zHs+Dx601iYeNg
Tn5VE3jUFDhNeXAGCQF2JWqlM0uGFHfRcMkFar/X3eaBtgTp0L8o3JQrB4WwBFsI
7zWN/pl2JC7mbqG8/NaGR3rgcBUXTFOfa+iXKTupDWiAADgcQE5rMvCvwJaV4icO
Hv0YkDgBTELtRb2+Bs4eLNfwW51TZmhCvkgWwwPVv4hxZoyBrs+Vef/rIKObly/1
K0+xHti3IWjTAFBHLQoXWjTvXWAy3R6cZhJT27RfbQl+2Yi0eejMeevPSWeQbOjV
iOEblbj1a3F4dYVqckoVbhbj1l5SZQzQepFtAtPvQgNQs/veOLfEOw7yrQSiQq6q
cEYhA3JQHqLKI5Q0nkeMTPzVuWBcbyrWygZEUEuyW06ctIQxddmn+zXVlsPw6l8a
nYBZYzKKptTxVKNLGjGZA3a3Nz66IdbK28Qb76yGb4Vixr/i/vUL4NobbzqmPxqz
qPNLZVirQgbIlm9rpmtuSU1lYRHftfFbp+eWx8W5/5I2OPhl9GZ7ukiAYPwt7MG4
HBohEKBwHt8pozAW3E/gXoFrEDdl8GewU0mlkJ80+JFcqaNI8mdw+QwcduJ7Al6X
y3qqqSS+xSL9nQ1DoFHE+c/LD1F/OGwY59clN9HGTc3xQU/1mMXPPr+X66S2QPAx
rHfqR4vw3YYZEOdfagbdm3Xis/nPoOuOXSU4NpHem+j9s9EiIcnug3LvKZGW7gx7
9MUConin7tkoH6H2Zfy9f17N4S5q6aJvg7eD8pW37rVQvZEMYExwZHg+k7pS/lN4
h5RjTO1FHmtWDVcz2Qq3ONu5ZtAuxg+ggVHHWEp18KxNnKtuciKLuOZ427pfpVmj
G0dF/ytKgId/3z9P3t8q8Pt/rckNyKHo0pkUa+IHSeAt8fxXftT0P6e3vf2xnOE9
be1XxLQmqEU1H8l/96PZRMVJ2aO9/QfN57U2kDAQpmHHev5adv09F5s/i4dfZ1AI
CXEC/5Kq8lpkrkvzgepRZqCeN0v+e2jJ7kq2nrxolU+dxq5S05ijuSdpsnxtrUfS
bqA//JAOxT7P/MEalA6B2wNfYKA3TNep4DWhTz65sGQvN3yEE4rC7+DuBS9NRBes
UT8ynuVsivy2hMiqQm0wZ4bmrjHvS2Rr8WcBzZMo3TCp2KFEkAN0ntTQRhBvbPAH
dSPjXzpJr8ZlX+ZsTNg/+VuJtRsUo5U1pFVihO7c4E+Qzq0crmLA3k+rl/dOkA4k
ORzm0AIOGPz6mzwt+qHPU60WEHqJhSM/7k8aaZgFFLol0FZHBeCUc3bXbv0VpZ3k
rFB/H+/9QP04XQmbrbPRSdHU2Tc29+xKqt0QH3C3fMnG076iTS5BhPFwAh+9VteN
MU6JM5zLJBX8TFOfZlMTyhKnExsMw+Xo7x86Z20OCZKGAA8MAWhrEznlFqawUrPE
S0TpGcEpTN/65spWxnE3+LkU0xr8s9T+Te2Ymg6Nv7ugr+yItTaBTKiaLwGQOH++
NM9XqRVQjKAgl5/5RyXO6N1NumGpB+0jqKiG6x9cgThuiHmVAcEbzvMsv5GaDWLK
JBRE5EWwMZS3Cz/zqaZenR3gZ9tS8HThtDgwPYM6/sJjwkucLD5RPlWMzowPS5u2
4QhpLZoKv5D3i/dWFExOvhiSTsn0kxX6+xaV7ZIlQe8vWh/oDpZJX8bYS3NZlT00
U9XyrCOylHGM0AnffKSBpaZcM5yRtAt8qHeIz3RSO0KOWtMd0Q14lnmtrhU/6OiB
ZJ3Wufsp5Qn1gZtpPT893Qoev/VSgrReAteAs4iZCxP5JLEN/7uxldkIyy9Z/sDs
1xQtwNIzboIn6l1JrEYuUCY2bcAubrOx+mlkXgq/R4GY6tTNKa7yoVcgORRWVDRD
ZCtDsSvvcpYZL38ch4oVQuRI8dHi7GioySZsF8TCS5VeuPiYiZnn/UsGlBEAa5Qe
gc3cBYN4IM3uu/BJz/JzgDc9cEDna3xzycX6OKXlzdIkMSWLrgnPUmPP8pEAHe23
1oyxZdeLriyhqql3p/Iq6Y79nroQvXQA8j4s9f7OrAPy91o1J35TUD0ZLvJZ9Wpm
eBCAKb0RVXCcfwO76aa63vRROnI7kIbqsvFNslp2fOsUWLQDhc/UF7DyRaQ5EuPc
lvV+curvXug4NE8GA/5efCIA2WAQOUnqK1sslsCN+EQ2+REDkWqVoJQT2tWW57Ks
ZgrSacUyFFEtestResJu42mZrhYYColvPpe+l3MT609EvUTWNL7B/2xUS0ES0lXK
ngL9pnBuMheDP43PtuU4t9oe7mM/G48RnU6rPQjHzPZkyA32uU+rai7+ngfEGjeQ
q5uI7uYw+L1na2Nc2RNLRbdUmcLBkOf4+mdAfw5rSufkKFKFdmBJKk+zmv4CKEI9
aV3xdga7EAs6HhwSrB6Z7Zf50/VqdFe4tBuxtBU0dHP1Z+9/VzxWgsDKBZRpt5MU
LJ/5+Qwfe0iRHWOvGGCD5pIW5QbeOiMy5RCF+bof6kMSP8sCP4zCNdRZVg4yOV+d
CyxfjaNux7QBG+5GRwKXQ+UWRp1PuUGP2QGaK0T3yefMmmBwSweyYtvT6VXjRYB+
RAZa+2IXo+KGyXpUE+caT6Sjn3+XcvItmePl/lOCSbEB17TVAG3tadUFLAzZ2giM
hW3zgR8ex/XBvrAK0UPkbhNbLt08FkLOo4XiokGfgDouoTtD6Le12fw582yfrmtt
bzrpTL9zpYO8i3bWandmEEorExlLqwjG/KbTsJBKVc73upzYrRzZAwJTZqx0yfl9
1XcdfqkfzsvbOQR+nrkL2Jd+PPLD3yIQCrK+fle1G4FfDPkA9VUVwmpkiHJRC3tN
ZlZ3A/pVinYbSb4w2T37nxrsWfpjyDx52/jBNy8pWNFnca1PpQveB0imh+BcBOiR
j58Tu08fQB0KpnNenzVE+w2UhgySVc/YzmL8ee18cOF5lj03vcOXM9P3/Ucfxoet
5yqg3cf6sytaF4PycYuVoZDEMlfCrbWVxBIFe4741zQsZOSlDkXxeHB6TwxxbWq1
BXc1Nfzzj8r7HEjEoFCM2lse12L41QfuvnCTNp/T3z5X431RiH1I3rtAKS0l67fM
agbzHgxmZTgyzMr2wCHxWH7tjRLA328CdkpNFDH6AjZ2atKc7DyqGhBNpDVQqveF
bgjJvMY4IjOFeZ2izKeC1C3iUWG9ozCAbWFuz6bNXp2zJ7Fp74S5XKTcuNv6nsz0
wCs5kdrJryw5JI5/QFCrtWHTfAnKClyc3KyRqfVP4R8akzGD9QqwCM+Eya8rIJ8i
9Ef6+Iin48hSJmHVWE2EoJM+xRyqPjx0lEJ8ptmhRaObBXFOVwPHKuVTpM7KB4Pm
ImkG+uVTRL/c3gya+hbPeXM+44rKJBJepPRNQmruP6p+UHGo/q5EkMHy0eSaMRpd
gZ+3hFscrpOwbjfYzSqtE+EJSl6c7EIAhkv+oN1mBkjyaxEvfd+J7Kq2UDDljRYR
6pqK5f6E3BDF+gVcNgx9IvRWCf3KsIiUnduO6tOyfMCMfzOdpAYHlDvf61FLBJQf
xLBwwivyQjmcPSrCO0xVO+qIKIM7nVuG89jyE6DB74ZmajuM4MdvzaYntN7Wc0hx
1XaEvRWRbZVXAt7PSExV4XSd9R692mp8J0lP79bOcJho3nHRQLkf2uio4KCvVNUG
xjTHiQyNSfKGtw6IUQu2Te2VHgnKK+TDEDmIamxYJit5ZTpe7BrG01L3qahpN9PZ
jnPU/4bM6v8xiz4sIux9GAEL4bpfBVeCR0AHiEyPC085v9OPDwa2+HYQodjqx5Jg
M4us/wBfTdNgpxLP3LBmJwF2I33zWepzu8gA5ED8kQtQk2H/XKM9GHBB95UtFYC+
LGGXh1TKvtDA85ayAIapQ58dPhHSaw9D0SJafzPrwCrtwVwEkuPhafWirfgty7AR
U6Ze3fGs+mIFqMHNP9KV9SldVeAKC73j4dq+HQ2//3FSdxYwJw4I+5YBIKnElJA3
+GPo/QtUFEab/XTM68FCvaVE3NyCxeV3xoVbtQnWu/pMACLt31XHKo3VhPJD/S9d
NRqm0b47KPpTcY757/lS4nJiYKp0jo+uS54D7pOVLbvwxAXOMzbm7XzhBn8NCad9
UZZ6JXm3gCWqn9YIRctNruE6+V94/gccOxxFUpjkMR108mRBfoUAkZMiXZR3rnBc
dYzAyKRvyxrZMioTfC0FnCo3TNC9NWAXZBiuVCuYTFz7viu/MerjZoSABCVnYxeq
2+MhNwHyaGMnn+keg4X92fW/SHUk7/qZaQsQT+ijMgCl7wHvpmki1mlLD8tRIgkF
p302ucHq4fAYfotYbi1DUN7LtAQkcpxD389kxLoEkmkqcQdm0iPQK9VhTyWFe0hv
heMGCrGbfQydwwZra3KKvGY+nt1vujitfcUrDtC8mvxMBsdOt5ApCYmukqM38Oxr
2JPTUBwNKQH+b+7bRaeHKXyHASTCSfzsdhuysM8fA4TOoq3ilJBEj99cXEUWPl8E
1GDl1F0exKm9DMYlMLo5AcljBLaumi+5AxgD7OxE0GP3vUzV6H3/P29UfVJIK2Vy
8sFcy0JSSmBLj2xQRGLOZ4+Pzl90rL1tFrWtMtOxUv9USTVKy3KRlkZWHRrInfkU
mjaT/A5vJvPGbNokJT6PwqwJ+lKnvX22gK6wqH9oj3zY8D84LtE/7IzW1NNIAJ4y
yMGA3f1D4zpkWYrzNxoccl3jAdyqE9vslvCTJ1jhFHV8sx3WZmcOcqPbRNTfHbRg
Ipj4ESdlZGl9oL3WfjsNxg0/iE7NKjpuA8lgy0k4+J3XqgRZz5ivIsAnSK6qEC6s
VSMHxlJASLVY4j1OJ9/Pw2kSWVwu0SsD2XI7TKyD2c61bJS39kECGaGPmcxJb8qf
G6Z9pubiZEfqXJLGiY/zbS7bR9RlcnCL1WPNf3LgzlyKga7bTJMAY7SCjDmZOXDD
b5HJTsGNuJzykhD/Fn79mIOxEsIG8hNq+Y8/z2cJYvUKbS+hcAbQvdX9GAzTGnKw
C9YCjHkJ7+zV6Z8B1eSNzR0a6eWRHcrcbgljzbd6YdK/hff0+Tkliy5tLxr4UMLg
6O6LT4akDUsklIZswBmDqQny3sSmkyNdt/VVuQscxknlMUpLPt2sh1OKg21ZV/1p
/zm2U+JkpQKd4Y8rtsjUC8KOPWReicXc4wLDhIurfpcrI9Yg9BbC9XErPoRdOJjF
Am8o/0rGiL/FZdIlDA72pGxS5StUYp8kwoA/FNSDv+Gjs7YHpNsF8LZSXAxxS71V
kQasWy2YGW8gZvcWGd/zqLBgACcV5Sla35tf1RrK4fTW1ju6l6ivoXbM7feY6WOJ
8o7AEapwdiQM9h6qPcWXAEqC3N9fG7Tr3w5Ny0E9EcFVO8pSm+7lIHTWjMlO7+EX
6F1bytS3pQAR5MWLYd6Rk3Sffu4j1GZSnJaF5TV68UCjF90Xj4B9cYyozw2MF6FA
XiaIIruLyjCSLlRI7kV1n/ujNJilOEc5zkSbpeXnJJ2VWZeZFHUl7Kg8TEcS90Y+
6Rk3s74MaoNwfq2d9kD2i7z3C8MZPgWvyJN0e7pnJVH5a6UqbnUz96CaVgTsM3M8
nSG99xm4z0KBfXOEAr8V7tWS4okUJ/THZ0zN26sGyS4lmBMDt5+jJra/FtFol/01
0yeLm6ihhvYSqiIpczycX0lhdBgaCguTfymtDUQrKEFiHV51HWb5zbNfX+dcpVNh
1Geyr37oHkGuNVTkgN6MJHkDTmwbSH18Z6LDxXR55Vtg6PMdID2LvssRK6WHwb7m
echoNI6H2A8sakV17dJwx7eeWFQC2HrORD/CXCbAJvB1g3iy0Cmfgzy2jyfLe8P/
9VVzsrRcHB1qoRuxOvy/jZk8m7pXoQqdCBqno9XIK8nhfnnwLI+sCzf0b+ZDpe9p
ZLK936N2TR6atGU6WX+7VjeRyPsrQG2Q682Yw4YX/Ep+CadqvJVowwnJGFVs5W+F
TqRIPNTSYeFVZICeLr8lRUwyqNX+OQKZMnBHc/ylnfN+ah0nPsEqxVqLcpLraytI
zSQ7WnEwq58BFRMQd1dimqwYOBdwHBZ6t+ctcyH6x6lrPeqdiMtKdYvsqZKPUzJN
bF+z4+sOhrYXvX28VNU6Ud0y5888BYgLRqvTBiVnrfJz3YHyAnOza3tffpRTAtIl
5uXeY1eBwuygIVFXFLDdwgfyQTaytgrMfwB9vit9YtV5wkpTO9VFHd+R3NP29tHz
4sq5kd3GTyfp9NpZRnXZwECKyD3yTZE0Thg0TDOMUiAZhJCkDewG3YI6ZQHrBLYE
qzVOn6jG+DN9OVPKdXSocCnsn+lj17+p5zTQe6OUE4UO233RO/Fxj79/+GHdipf6
VbQyDInqLlEBCwI8D1v6gHo/233NWMpkaevastIlixLPfRE932HqVsrKlLpvcPcK
cBvKmHf7BMtbmwrzBDHbwLYBT9jrbphg3RzS4NxpuloD6DoOqIgUTdykPPOJSWsW
FVn11Aq5tKDfXWhBUE6ObwyoOmQ99Zm23J+Ipbk5AHLVwTP0d4XgaCozMuoTuEIt
lqCX/++VBGnBhxQ7uNfo1q1fIDwlGKadGsHf6eSIRkTtdKUMT/GlvEobCy6QeNE6
UG4/M/fN4NMLpus0KWSLHruArebNN+l9mBqhjwL3nZVgDMYlp7hLZas89bk14tfZ
5zt2scKm7bK2BW5R6lQbUbZuO3YlDmzV0p66y08+k3OXs+kyfGb4SHBMoF+byqMu
8mXaSCG9LDqJ9tn1lNu4aURrvWK9I63VyYNBVfdPOvABdQjVwzfBUJXt9/w9oUyH
LiYwwrbEh0PERcIvB+AjUjYeXUzn05haqE9MucMS+JvbIjUZNNk6WAgCA+BnqpE+
9K6b2hN4ETG3AZ0nsCLQmTsgcc0RQSpi/zcV1YwflyKenJFDyBM7TNhTHIUMqdhj
Pq6flsH4IblGbo+k3oX0/gHmRiESnURG7xnFnEFCjffoylARj6AY6hYWiK+0Xu+Q
iMppRHpRrpATsnr7y3rdmpMzapUuOpN4X1QCULsBNv5WjTJHX8tftXE4UwpV2H6V
gPepoCRyyHAEQbufPLgi8c3DflWj+8d7MZTXOmbRwQewNAinXq8GqwjSUFrFCB/C
Hzf0wezTEHa3SbDSBZdrE7mi9ox++ShN7FWIhgHdflGYq8GqMBVkCvERQ28GCE12
V87u1QsFOj8/+HH5YdBgP9KgZNz0P0QR9DbOhqjTtPxcrX04u2quQ4lluPMPhDlK
HAlMa6bGq+DiyH9laH54/RKDl02EdP0cljFABwv6WpjEAZNinEM9V+zBYU+tNusE
3SfaARkNLQrF69G8dcG04iQ9HDmfPLr5nJHJSGBojZUnGQA6N1ZSIpPVYzNMBORV
9Sptf6dV7dtkZ+2/b0y0sl42BqfSAD1jtOvL9qEXIfoeI/xwclLCSKM/qbISDbS6
bAqrnB4fOyUBN6nv3Cb9E7pmVE2alqEyKOCvVlzYvenuYpJRC22XcgKKeD/pehWt
t5CLHnVNv6xeLRNihtlEynyo56OesrmbC96HL8+1pt33wyts8KPkHrojKNQynURE
aFrfG6kGu+ccB0ivvJaw8BpxWrYADpnq+onGLqGQlhJnZK1G9CZr/O/QFrWMruHL
mY9ShRfznOr1l7c8sF3VqKMUNEkXN3XnfOi2uh15sQi7o26MZ8q+by+pAVCgjkHO
+1wdbT1wAE5AZxkd+uBBFnPJdFUQVo8QEEw4XfCZIRDexSzWGXU9GXqQuZSC3Tvm
mHxU6IFmPxC9g+eEj3c6bzr04+nMVVAshzZYC1rn4iO1+akVmr/i09hVqkJmW1kK
VxfGAOQeQGMJAk2WVU306mlWgYDj2C6/hr7AT3dWVtPr0IS/PVwDAd9Rlk2LHeDB
/pFSFulelczOGbVk7YCdcCd/IBoxArGBe8xtyTmXNGqYtQvWnwhU+0FMRVNTUEua
gmjQhNbR5HaAufMOJSD2qol7R0Vtv1z9uFezE1Al52BJ7S3YmHA6KPhWa0CmQ5tf
MuPneJU3+7Bw1xZA84XaSEs32La6Wc+g28qMpo84nO7I+RD78oSi7rUwXdAl064H
Uy01ezEDzR2avvq75bCf5TzS61VJD0NVyy9mtFEhqjXg35RdFQ0Sw9LG4tQWTj3S
pH1AP21k91IZZKKDR53f80E5q8qIxk1U64UaYTgNs8or1/7qSjeJZgF4ktdi2Fba
Aa1KpeTXFpdIxFQatR5i3sppVWfSFUT4PyWeoDzn0qnP7gm1hsvcCPOSa5dSWWlf
FxCtFOzFONxzIJIz8dcCzZah0m2lKkIECpRI6PqOd76jpjBTbErDbswmm/UKLQlj
4Ja8ry8lyvxY3EYtAtgxcW2CDxbzy9hE1cU3DNUo9QcMnYI+TBEF5sMVDlVY9LS3
3kTGM5ctPpr7hDMnuSIz1fMSsgRAScoaH6oPHYXsl7xJIwz3xcFEvVATY0eiv6qF
2b27kS1idOGo/F2VtHEt2XUFJDNhnKvhoVHnW1GfnQmm/4wkWZSbGpB0xKKeHajF
/u4h0AAkmCoZXn4B6X/+I1TxCcDs704E6XCqy3SrZkHATSjibQfmAm9Z4RWT2Nol
USesT6c78mb76MF1oM2Z/1K5MJbWVevJO4gga86SzaaGumZcorPZItUwrNp4esxL
m8lIRocQHHLnUFPLL/z04M7YehFiWDI/phK6421d0/sVJoiD8iWqHDs5Q8wIlKJ1
HF84IyjB+lC2qOTP49ERWM3LjwS97ZGBLbQBjmYy0INIxgUyKlEUzroop7cnb0Oi
PIZkFr4EG5CpSmDbTrLR+UUoUdZC7KipGS7gDse4XwGH2IAcxRiQ99RvC9X0zQGd
uDqf3EYkclD3p4I9HEJOHLY0n0d/7g1H7bfbTD+Jlgf4nZjazowJYdmvOAGuVmQW
48/hX1pAlrh54iLwYF0jGwyNWz7LcQOC5CuRYc5EWPli+JoANCKTZcPZ1/Ej5KHl
tnaydBIJ4b9qvxBdPqARdFD58oPpsansH6olavnhpNABI2n2WKupPgca5YOPLVrt
fHP9vkmH/D6wcgxiEUM2gevn65/itay4vlCDhF5eg6583ZuzFziphci6swM6Mwn7
4ewYDVJuR5dsYFqRbP3dG1MW0LH0yUUjGf3BzOl5eKhUviaG5QAj80+posYpBTat
pyI2eK0X5sd2UBTRenfllF6ck9pO90vlMp+kxnyET7hP3kCkyyIIuMcbxFh/ilFk
EtbOMI2Q2fNpffWZeGM/xgy8egmo/nJNpNCW8CU2VqpGu4/K49J6W6NOO+cwKU2g
cY7Kru39Ha1Cp7QUK1Is0nDA0pYmMJ70pnfXgYyr40rfd7C1lxiKepebThxTNzpq
cyeXfdNT092yNe8NALI9uAxFRg6vOyytid6ts3wpHwe12pp8hc/9/IdHsbudH0Z1
3u3z1gU0io26W0qmPdqjSexUmfeYiDpeTi9n7hAM8KGxfDssj2LYoTrIU4OAylwv
yhPf8UuQJSuxuuFcfWvUVVpqZPPkA4qZnB/VybpBUibc0LTbL48PzSbIfuhBBlKF
y/60ehwI9gx6ziD9zgJMAq1QIu+btdZ8SJmHlIaiSP3IeCNGe0cAJbpG8ZIhH3We
RGALpdfjwnFllGqAr8S8pUtA47mUg22lMiqKFmj0NTEhp2yhvaSTVbwpdbaTuMvd
tLug/f15NcjYhRRxtyua5aya+f9AYRgkp03220HjTe/KaYGCoNFsHpOvazKEehGk
q65N1akn4rjAR6xsKJ87nH13moRHaZoFOLGSNNCyA5w4HsvLF/eQ/0XiT8bBGZDV
fib+1EUUOK4xZxmu3t64yxJlopJoH3x6/gIHLsCaR7ZUq10SjBD5/JlXJF9u5TSe
IQiYzuNUR+LqJ9xILFNix1HuKgFNTFRaEen8XJXTt9J6M+tk/UyMTrgHVyJw59Sm
DsFFkC3h2y7vCgcRihbO65/5/AsuV3HAg+7xCO18hs/fpAZPjfT7aFLbAE+dLiSS
xIbrv90KbYm49JJXLk2U8rJ7iT7tSfzYhRHWrMxkEYY19QqKh9rQ1af14rFudidh
WrkU62aLEfoQ9bR/fRSoM7aKVc6qjfapWXK1Gute6CKOzPbQTrT8pU+kicBSW6o6
VkW/MwESRYj4ihhmPasU9macYKxfEEBP/8cmk6thNso/sIgQtmaiuV7FiXBmc8dM
wmuIpic8fudMxgkbA5h56x5hVNIWkUbFXibT5xq+uM44QDq+WJTgxCb0aOMs7xsn
7WGf7jwb0Lyu7/hE7PFj12hdMpfjq33e5GirfDtQxEVldFQsAy80cqd3KWR98tAm
eVI9RoLjS1vKfHshbVhUZNka5/VI3+4h3fp3mJnyvLe4++KqHdp9b92N4OMKTtFn
w+ciizgl97uAUxm81/hIC7juwJku6JwAhSZ23f0blR+OWntJ7DiLLSIOcCBP1Ht0
v23L//uCfVVa8MgE9YC0WsCzyYGuAL4otdIGdN27TvU/9f/CtmOKLIBQsC2Rj4YP
HD97Bf7aQLWT5OBEWqHnqiVWLhuN8nXzfnOgAR2Ccy2zjYc/jPz/9dkx5QnWJkHF
p5bnXA0MpV65wRDxix9AS+X30kynaA1mJBSI6c5e5dkbB095E80QX+xpVNzWZ8wj
5Q06hyuUnZ0RaPZtBcn9U0nmBcp49EwOJV9DZHkeShY1vDsJoRA6v6yQ/8eU+WdR
KM//iHaLGIQ6n4R9EFff2xB0l+1D1SNSlBsxO7EZ4Ms74Dr/5JbBLlH0AQD2JxG3
jQ/t4Z5SAAugePx2TLYR2Mm7k4WHgk45O7j0MkvjcCMzeLA1/OYbDFj0XLySbC0p
J4HTKMp8xL02pCmyN8WIJZYJj6OqjohydRABNCM8CaWUtYZqPmKG1E4VxIDPXmXd
/FGzG4bEyQZSD1NCu9WdMOpd4aaohEOxt5ZHlddwJG0vJxPjiFFX0U5hVLkWUF4K
s1C+n3nvAQzvTXZ3Toqi7M5l4xBtzJMQCDv3cJXeOrC4o5qDiuNDuvyh6g1XLrkE
YPfqdMCARYPP1gc7HGsnx882O95xQ/grktUAa86kFyVv5TXuOnolf3+De2MiJr7Y
wQLvy9e9aVDp+uDJ6EydCCkuzgZypXfyjmlsisDQFnlELVJ6wa9Nxuoejr+qJhF4
2OmHvxSoyxJc7SlQNo7wgDq5MQCR9ioVVPI3suku9juXiMfIQuvgYOzcsHYgEtBB
+8hOAqKMX+CvsPPjqzihq7IAMsOxDwnu8Hr1QCDIHHGiw+PwyZyiTO4Vs9CQwWwN
PBcLSlfa1K721Qcj2+iFa1izQLQG1bOUtXcPtq5hbm2k2vQKgLDOqpcznER5yMBy
HpMzEoychCGpDeOCrXHHLlxFRTzA6c7GvUtDsII7eVRA2W/aOIOQYoaY90govRVL
GG2At6d3GLm4285MeA1U7DyMx644zVSstn/cFxcfWzr8rb4AD8FLV4uRYQ4yLiwm
l/K3raFAW4bza+4U+MzsJvZ01cBS9Cg7cnJAhUmTb9sfPADkNkCcI8zbEvLY+WrJ
AusGSO63tno4K9OlNt+fiPmZVQGyehelCut0pj3pavFEiIOSzMV/g3tX20R/r5Ej
/6+NpRr02Mbh+vbvGdxe1YZBDXRTkPMxXFSnKU4EL9LPzOKoDi1h6+b3+Y1avibk
DThWCA8/XSQWVwH3SEUho17y5TUwqkN0uJI48G3FY3ayDO5rbAUrsYQ3iGBfWBhm
SZ3oofp5sI201d9V05er6ITTiBWbSdoUsJfVUWGO9cwRMMhPxxta9nVv8zmlGNqd
/Ldr+oNZVWzjTee12BqUsryOPkrkWxJXQ79M7m4ZuuI1aNlkrxNtfnm8CihZXv3L
hB4FJepr0U0PCMTL4J0I2bkZKtc2PRfvj+upvX7O62F31xqP4Af0SI6Ou4Q8gNoa
M3F4X7UXHvT8kMmwORDLb/GcNFJAHeob7MjqxL1XeDRIzmhNWNYcLbzoMbO/LPN+
x/NyBCmwUpLjWnhqDA+E9pdbZ0+2jptEWbajWI5ikV/4cigYc+q/QRXw851ps6xF
SNCq+VWYvFzpU2VbibyQAB11Tot0SmZXqJZFx9CfAf1IDUfWAMVJZGOdMflloeil
53G8zWQ0/XtY7q9CwbPXb9AgeL++s0Ot69EADFxKKyCNJGWuxaP2pvEhVGwb2/Kd
3yoy7Ex5YK8TMnosuQpks7SZzZtC4p17pRyAndDTUeOS5ZfEvxHMzKKM1RI86E5A
VsZ2yFLpdZmfM/Ozmbaws5KeVjyP36SbPMrxfZzg2FG21U+38LbTfO4PLrekQevM
L8iy9oWR9s/G8pFp6kADlTDjGAyhMSW8+5A8QAQOtNZ6pgwsffEEz9RU0XzdZQ9i
9XTzPae08yYRqUCHzMY2zDEoSnFbMiC+NLUQCUMOxUbz1tZHJFcTlhSfrNvlAlHF
Uv8s8cgqY+MWtkSwdiMZvg6iCovRgR29MP1zMfvZopepeFUI4T0tn0bSCBygUpgU
ncyEApazQqwt24kHWPCvNJDyq7pJ6eFp5NE0aRS1q6Dg2kWvwV1hHj5OGLOAY/Am
0YILP2ZE+a/SAkqad/UCytbC9y6QOXqhNp9VuQL6+fHCQR9h7ON3muuH+avKOoAq
dk0Yu2yA+33TZ6Fs/y1hoztE1yGZkdbLPm6xHzEbvIsdmuaVXYEJ7r/zmSMzN6wt
4qQ4bKPHXyeXVpbsTs/BiOLb/igE08BKmWYESBD11NDwZGJrulTe+cYFFsvYpV4I
cVNsbnVHEvOCFAOFtajSUKSs6LHhSbjcIlzCqNuoZTv9KUQIkgYG5Ghv5xVqZ8Am
6HOViKWJhF/RS21tmRyLbkii9H78wCXzoB8tk/bHmGDP5koNq41LmBAI8gXi52NX
52l4kGb1/6waAynOnzY3y6j1YuYXGD19fHT/gAax/r/Pa78ElLGJYZ2rXUqX7Zo4
dFGoILYM7x3UHmFHHj9dMf94CNyv+v41zdO3pkTJbNSaW4P2y93LPSLf0R+eDsHI
jAJ0s7lyWfFQE9qs/mYOjx7X4iwWqGgiqWhCIc9i+ZozAWU85PDeKxDTqLzhprzk
YK5o43a5EqxGU40M/o3zNkdUTtvxp7nVJlddWma5YYy9EteK9NCUXWlOpovPutQb
6z9itng1TiL1dGjHN63s2CDpYeSrEgS6m+dQReuDJLjtLgr4hLVltdSedTyy/HEE
2PSlBZaGudc+5tADuTR3CCl7eAWnXgd8blxnaFB0NQzDOjxTU/rgiKgOpqYnY50M
mg6JTxQmDC8VgIKZ3uOOPqajYX7Nq0ibuD5euW4JJKTDYiHtYwaXUuiIfAPjm3FV
jd5+vJD/vWDDuV4VxbvI7Hb+LHMeS7HLWMuxnTKzQO/Ol6ABOjoPblpXEWY3WbI+
Zvzcuddt4ak87XA2/VqY7AMv6pKJS5YmtKUdQY3lK/PZAw+c6zLHBQnm8S1yJkZ8
LUepDS7xMhZVRibTdDQZzfyLB3mdFsJYgQjN7Rm3NqT2aSMJNCmkNWTf/iTBdvaB
IWvmTdXr5BPByPSnd+L6axzarzfraTlM29Ou+Y9Tx6s06AiBMeuk9bABUBKdNncW
lV5rHhzaJpXkh8rwckE0/186qx1NdXBOLo9gpAAd1Ui8uH8rmXOeQvjpjjV6Gt+k
cstJN/PQ+LhHcROF+pHE54tm9RLpojeE5I6gkIBWI65FTIJPYVTQA5TcPvHNuADM
GrrqFacTaZY3XYjRo7qV0kbJSg4Yz/QtyO6y/yHcE4KgLR/P70rtEzkhb/vVSAB1
o0t2yZwM/BBXQsbSngKd7eXKLC6iiqNTRaES9pFP3mmI6NVafzWI4cAljhKoaEt1
fTJdMMmOV6WORYL8ihwlF/PeyZPN6817KByP4bJYPo/oRXiAx8P7Z/COJEDl9hIY
NolF3TTtI0cxwd8wl5Ula8xFV/Sz0VJCIdJqS86Q0wkFh8ixskpgqF6xk+21MGsO
8CY3Y3f/tu/VIIK74WTcN2bjQF2f8gOY3wIJUQbivPZEIUcdVECz3cyP/hscw9yO
xEvbKoshIbGJeD7Ewt+Ex7w+hgYAyZIn1NF00EltFJT42TUrrRmNLzp1X0/paVqA
IHwXzB2E4o6b2xmxUkDfqlfp11MyS+er4ta1GzpbBnjlkK3vY20mvKJxJtV34Q8f
2eH30Nu56uj6a0Sjpm1on+rbr2okbk66XVhDQQ7IGrgXm2QHCPgRVBOXJiHa4kwk
yVa9s+GKXOTP8c+6Vv5BVaZO8DOuW4k/lbR1AHktgcXUDMKyY6PIRMVBUgjAy4iT
2Gq37fvK3hjQBDzvve10Aoxl2uOCiGyW2uHc5YSKi0PM8aQrSsxBRetsJrawm2Bg
vosSsv1NfxzrkllYvwIH069wF5gS6KctUzqicq9O/ITceFaffQ62QZPCr+MGADCa
Yc9By4pP18SgFqWDFO4KBIE3nH3nOicszBbqzbPk0f69AhPNVPd5dWkdfiJ9DOxQ
DbKR+YAGZnXtojS6L7waenVRKevLxyo8Dw0KFN2dU8ajNc0bXEbZ5wZy6Qx37V86
Xqs94Emg9Z7NRzs4yOmpQALRqDT4476NIHy2xfcIoo5jrIwArUdApTfr8X6U5RIx
Krcy8slOnDGDHsd5tCYZPA4OvfNH7jVAKKgv90+k0uYENUNEtntzBkdWF+03Np4R
RyS/5qr5OFxmI/bWTY6p6Fer1VZ1QhxwGgzkoBC5cl+p0OATUaw38jRhdbrG7LsO
nz2AeJERqwSq6dj4I9JBOkRxGiGZ1BuspvbVVStt5TkPb8z0mEcIjWqxdEk7YyW0
zm8jDWDDNYnaeTSxFUQb0qgCA/5N/KSYw1u7QPU0De5g1SmjAIbs970rwctmcqiM
K0y3Cl5uphMSMpzjap8j4FP1J+R94T/j7USy51LYhn8wHb5R3OVfpCZe2FyZZe2l
fFFhCeTXPJLkb41H3wWf0PTyeHimyB5N+2Tc4AzTtVOTbn6Qnz7QrybhxtoNB9EI
X1NKU8B4a9Fqq54QCiZgGTW90LqCQHRy0K6X+OXJQC6kFZWt670LO1Rmbc+vXYop
RnWRr6smBlWt3QMiNUQv6wo6Z4XaXicj45/0HXvsMfBLiY7QkG+ocggt4Nuy/jjY
iEyDpPWvOWPtccxtjIGDHAk9ahRGL7KTd4ZjkzMnMYYWGUGvM2iTdbqB49MYB9wR
60ddt3Knw0lTWPJxx0XFAHxt2X4ahAGGdGpvGFxnNYaynA3aRp8cm1Wx1dLu5z9m
MmIrC1i7+wq1EHw7yhsmaGAZGVZb1aFn/jVPI4zmENEzhskUpSeDda1fEWBfohqU
gVS+dbOHwW9+JH5V0zEB9I5xakv7uIgqDXhvC3QVQNMQ6/o1+VtvaEkuZiyndpTF
v83d/8m2FhcoiCJkdkILKPv+SCFeeGrb9HR9fL6O5vk3I/CczTpvkYxdHdLmb1FV
2yH1njbwdDuaLe52Ot1Ogjy98LD0cnInXgVmVipNGNFkczqCHZzphhwlyPJi6fYU
EgmwSQeYxTAmLZ90kDt7higiMaWUhkzzCnhHFRZBQ79f4H+zbR8bVohnlObKhzJM
0JasusjgKN40wNUJ5T3OnqZrHO9nsNjQ0H3vgoQCN3qzQ0atiIudqbn+PzpoAb5C
N04fEof1vrmpNuyf+LRJVN3HhT2Hn2HNxmOWvV2mw0yA0G9IrttWq8ZiKBD13+cc
WHnp6qgYj2iDaZqmcgJvc/bk6gPbCAz1y2dZjnQYvHXo3Kjxk5qyw8rjc6HwdxHx
t5u/Sy7amZ2ek+vMoMBAiF2vrRjBO0nzm0FZUIy0T9Fxiuvts+tmHCiPzCHI2lyY
GEoRiIiETpIxPUOMIeLavXzpY8cFQM2pAaLripOUv4tmjP4GpIzwUSrLB517AgIT
GO8RpG9bP4HxDpK++WmUaNKGO29GMHI0QLIl3Lr2pDy1GP3HiWg9o0BmnzRc2tPA
MQpqysugxxXAHmEyTUcZ8sm1/h61YWmona3uFYBBGoX7+DBLWXt7Iljgk6Gewdkn
ApZgtVcMSD8+YfrRxdvuIgKBxeV6H1+2PaG/a/CQAqM9NePbLvcOszogzu8vJoKx
vV/vaBmRo6oRHU/Rt0BU7R/njTEd4sIMAr4/l62JuCIzpe1EXoUmD+IC6MM3Gj5u
TUE1cqEr/6FrtBprUK1nbYIi+cArcrqHRhGQ0azdohJLR8YJZYDjM3XBSbOkNWDN
HwP67uMkcJ1uBwgEfWTtjvxW2Rdsfcaf8ZmptEH+54t0JekCNwBx5UJtlVqq5YzB
OPzLnHAgg1xNuFr67jojgpSN18gm5/pgLSREzumavb1DeIIPGx1H1Uj+xjfAYSDC
2OcvcmkU8tUBKRJNpL32oafodoW9qBe+q/jE1DJOxBKj7TfneugT5ThVyvDI1dCS
t9kGN9hc0XspCvDC22Sk93EjXRgww1BG5xFbGWQkrqEL2OMj3O4zB8oPvxRB/pt0
pS9eHMOH8vlxDx734E1WTLUuxGcSLKlCR0bLYIvyE5Jx0E40haWDMsuylBZwQhF6
p1enDSELxIFnGXBQqs3bwNkcHkungUib0cWzL6klr2mZuBdiEchudI9nPk16h/Ho
E2O1Iw0O/WnbSY9jURBIAr4sdZGQrPRen8knFoZ3E+NR0RzYCxIEpMy0fGC4Hcz5
UUmo/CwGrIkAKtJgUYksEoMIXvuxZFT8MvI5JsrL66dHapACartKlMfSICk1tSBc
EIuSxMkmqXbS6duxXIJKeeIg9hSdn6uRC2mmeP+0wSlV0h3ZMs185kScAtTHLaeJ
+y8KWaK3dRRnTsP2ZqMWx/y+3+SVVTQe64apHHvHFaTtsY3vKdSvMSqHE8i8oYax
nVFYR6wkudviH9oYnlacUdgoR9fW6zKLiuXGlkdTNC5S+UU0iUW3a7Spm2w4EFLr
0ho4of3itOu0id4XN4DkTU40f97eDRgj16NK9Az4b6A0LknnsIdJBjfU+6MD0Di8
k6tKGs3n++h4Aku5baGcVhfR3/+95k3IJdWm4V96uQj4tIgpP95F/QhD1t+d1MaX
UXAAqUeBSS7dwURf1eMsX/fu3c2J+S5igqHfjMCreSKTKoyq17SpcI2rnaoXPdyw
zJAkvHkm0x7BSo/BtuQ9NXgblyXkgewn4gl7XQ6wpUR+PBywL/2QB9CZ99Hw5y4+
/UAKKs6UH3dMTmIb9/vEmXR8p3b+F/DY+Y6ndEUbAtDcEQMrYPlS1EL16DPbSwRT
lBAffdcFYfOmznBOiChKSxhZauvvIFdyesGEotF2KcrM23DSjmiRRf/8vOEV7Xn1
v3vT2N0ovq+GJ6OKX2m4AgADqBIuE2w+CflcOBj7FSEc9Q+Nj2RoPXM8dQIhc3VU
aJkK1Np4Gh0LH1jyJPH0iwWkmUNBB9BuU8tOiVded1UCHuMtf2Cg6rklxT9tpah3
50k9VnnH6Mz2fjY9A6njUhuy4dxweYvoEn7iwg+nk4QWslT8bPTVhFuPrTXhlmk3
ZoxeSvoQqdddC24d+LuhmN3T8ciS2HhE6s+2GtQ6/TdybGrI8VdLzGyipH1cIKBN
iXO9WXZycnW0l9QQFIo9N8hMxJakRJekKnkbyiwfmqcvddpofZSrnMFrYP5XOtKx
IG0c4bgIKpD86FKH4Kd+KPk6TluxKHYBQphUNcVPKIVGSTC3FiqYfdvx/C5KRWjv
/0oYUirR3VNeeR3rI5i2MyLnzqDKO8qkzNM6XuRN+N8XizWfEDR5nY8n5lWUN5G4
Y6LnKq09Df9A0dE0iPFKgaS6F8CXEk4vAeigvP47NezRVwr3NLk5cpuvbldtgF7f
2f9YnBKOcor02CjXvMIJQs846dCwI7D2wFLp/1mYahQnhIol7tqRneRzcsm4ElcI
INfAqg7eo3LbvhVZhxNbsp/Razaea/MKpLfD/fIC1r2oi3rW6HwVq3anj9ERQeqF
Y5cAPWngcQH7pUrSsjgUaziqF+eawt7iXcISC1x+urbesehDl0Y83P0KQv5iWXhy
zhb/yAgWkyQLY6Th8uQmRksbgeKBgzCv53MpaZpWebt3KI49DMgap8eMp+cTHmVZ
tRX525n+IlbzxZrzHYXZ7KJRCefcd7OadKSrQWgm6PXQTB2BYoie51Jc22yQJiKx
nKIwHhO8mws0ccuekTIu04aC6Gi7B+C9i3uLMa1JDTlsiqhUXFbzXkYHYfCxWSTO
A2S4IlFoBGkycjJPRe2PmfqkRSn52m/jJNxCTmJq+Vb5YnLzl3C6PoH66p3rNjhV
dm4iVDY6J5q6fAQdUPXAFCdhzacdi/r+j8jtudEFeWA8l4M7276veFL4ey6vuyRZ
dPfcdLE0tkfATwwX6ovwnUVH5cM9SH2F4FknO8jlvQvjrOzxGOd+dqhpc7pqSEYB
TAuuAYzD+sOzGCCOONNw9x8fBszTL7W+Vi85WYi2QGbFInK4aPlJA57UejSS4rW3
ZBxUEUIqct8DdqGYO31aw7kpQ4/CQETyFlorkzxzqkUlNNPuWGBWS/Wf0MZZpdMz
dxdlzcEYJftgtC6QfDj8/l/9rIWBqFcgRyJxvLQYYBewc/nSuB283tLMWDmndg2X
MqmVDnqXJ0D5uMhhkh5NJClWFfjLl4OLRHlFt3tmtNG5yaKBRawTswc6azU/ggWL
V1vDKSZnMNAIwXG5wNS8aCidi8ifkWXcYF/UsxvS0RX1jvvqVvXFC3GKomIHgsDc
n6cSSAdBMcl3MeI7KTUT2qhkqLafIV7zzO5m7gUwpsYh7kQk6xexjw/6bh8z9+rY
20KUC4eHO+flu5n9EzXH0/E9yTKHDQNl+yE/2khseKF3RvCFBIpOqUyMpgpsX1OH
GAtvhaPVExEjeXIDdWdgWelp9vKZIam8Ayxn8Zu+LgrUqCP8rtoycOsXxiSceptn
7sM9qRSnpfKLt2M78ljROwNXt2ub11YOM/hufmI1RP45j4dywmMsZE9M5noONK4w
6C2JkH5zlZjjuh+k+yKTycbA6i2CiTbMRbbeycp0gM6vRFSGyeFPFrmwg2vXX3AW
dHIw1BgSZ8lSCO7Tr0Q/KrB4TdfusC6RTW4K2yzWzu1CaRtD3uV4TsZI1z96lx8/
2ba/+P0fBBkc0fn5pCOgHiwdKei4/KU9HpyCHCCL2wM3dj26IZwusl7r/7zwozj2
FoJd3X8QIhTnI/9PWqog84JK0T0rmgoE1BD6V+2UDbuBItYn0YuMKYwIdicy0zKC
Kl51tKsdGj8S+A3NdvmIi5aXzBZG+dJ3wRVSk51BMzK4HTStgUrK8cUHmLH1qW7s
ASsbqCBvQpUBjVxBu95tlVuwhY7MRXysxmhe2DmaLGoFsBmtisYTZdiH00+85cS0
3THXwlovlye6yOJZR/pDvU0z/TmiA26pCY8KpcYfIU5BQEB3q7KykNQI/n7dt8oo
5Jims1dC9mD9rYI3etfanjmuLtV+rM3Q0CFte5/HTO1fkV/GIAEDGp4AmSgrV9A+
ZdjpbLIsgEgqwLOk4EWKrAauYwxPN74fy//PaRYTnMRuLRwlEBfiBOzul5IcKr/z
9v5R5VI7d94vINK2X2OynO/wfFVHPW5W2Q2MTK+a42bgFne4h0VJ6+2pz/83zhja
KAsnjxzxQ+RhTnvp/ctqZ7SxSJygX1oUoR0Un4bvbO/qb89T238cEamNZVxZ6Q0N
ke1DbnfplXEt/RfuJOxoNOAeNTpwHU63nY7TTUj5fqBIk7fQZjL9d5R40jiv5qY4
KULGq/DXt0nChR3gDuaQP8GeVc/dp4GnmZ8gIaoP2p+VsrLeuyhgCdESXToIVSXV
I46Kbja7ttpsHah3aS5y+BrjjBz3GrvF/Sfyvkdc1sSmcf22gRk0Ux2ZBSOka4Pf
vsFE29/r48g2cKCSyzgy2IWj+WVWJwdShhDH0ebh5ggdQl4hPB2+fgVDpbW72tQ5
ZXilXgDfBrECejqUliU509DfkiU0DbCWqCHt4p4ru/G4U7+3qYFNIQwz9zkWcyGf
gPN5dWnushqVEZfNyJqFKnT5dopwsXs1bpG9eOg8UqQmVN1XHA/nAMu5Bt80tvtA
zymEGgDDVPdnNidDbgoXnjHph9KGY/BbCD9FbHMQcLJ0EbMMctULIniVwkf038f3
m6LHIA6QCw8MXKVK3KTq3nF/VKwgDOur7F2hV6UY32lYPciJ5JOS8DZEgBqHoBXK
O9WkXSXHUeQtO+JXafuKapQQ3IWvEkYSks99FxSKN9NFyZCzqIAReCRy2Qiw4glb
Fdw3NU4vPDBGYqX87nE7NwyX4vxsYRQz7tFN6K1p1zGm/dnXU9nSezkJZifDlX4J
HyIAC7+DrzjGEOxpQAKyJZPTlQ+qIGnA1a130BjQjOMGE1DUETYbl/otWNiXuuQS
GA6eBIRe9EPawNwQhDB56PJ2uBXSK6g8K6VPnvWY5FAf8ZWL+9HbUrlpIWCAOiSZ
maGIAjpHg3g2Z4HtdQzHOORYqsPtwRmW5Et/bbiQrWev0O8zibf7EZDkUXn62XaB
/ULBExKIrqhqfbEuFXVJC8rXgfEPQckeENCQv02j8u5R0RFhmBDgSxFhraUE0c/B
h80iewa25bk9cPJEo4yHuJfqg2fjqirXvLfX1a8y5k6GDpVYWLnn6NErDJ2mpEoz
ZAaEftM0yJcDlqOxMQ6YGcZZXkP0fkSe0OPrx3womPi5fFRFTYXzjLAopIA3DeKL
WE6mvUdMAVa+AYPMPo0CwcQQlNfCyglyreHgjIb99bR7XnqJATwJKaDG+zaRDyYm
2dGgROsIgGJifJiY7tdBmbYLk5H3Fy5gqq27XZ2F4sQ8jAIi7lhSuEnl+oC1gxVi
G+kCBHHDG8wUTntTnpbhhEuWvaocO9OHf7782pR8Cz6VRC8y0bSw2hSVPnL3kWl7
RxCsHnHYV2LC5VT8+BLcm2z6DvBwh/+9z4o8gETCgmVcIGDbVXdF6rdSi8y+H6ux
FAVS+1MZVnJ35mfoNXRjYnj7+Tm6SVwvzaOh0d3Ytg5Ltvo/qAgvToSfkw/I99qm
suyX/mSqD+tOntTtnUWQmnbAwo7brEsNbzJYPoGeBa21RzTWsQZYGsMT5niFEa4x
i1rdDfYZTCP4u/aXcSMAKzS8EjuM99bx3XVlvhiIdkJjFW4anskeLWMZ6EfMQgws
+nfv9vdmoxA3jWCtcHSAjZX4PppsWMXHrWUl+BfE6LW7X8nhcPfF8IU70mZFvRj6
qT4MJeB0fvyF7POlIfxKNhkdtnz5ERKIELJnVFm2J7UmlV9PJnOUKfU0/leGsRou
NqL7X2l+Q8f+IVqTw6tx7zTo3+cUMJt+tPTARBhAjxkgzTmYtuZ2i3NEnqOePQ+W
Jp/hpMwL/cr5Hr+52Q/JaDlQhWA1anxqByJbaSWYf+N3s5Fa8nof1pByAlZuGBqk
APHDDZTPgomaS5lGczusWjo5FOYUXBeGtHlw0/XaEs9nEFtSzIlHXNI5kPJYeLQt
JJWgQ+DgLhMIAjUObAOlm5OQZDtnZ5rlNna7QCI+8FY75/FSe+rJiYd5vb44jhfk
xVNxqyuzw+Kooyd1woYbVVEwlzA74FBWIgNbt5bcui3/hL81G4FPDZcBSSQ1G0aT
HFIM+frnjPwgeE7+eeMcVGOxmAOdC4P3k0g451QL/0Y7Gd+VdgON4+QGKBba6iU7
YfaWze50HVh+JwNsZiHbBjtFSa/DOKgbvK9tPjoULDbmdlcyPWWDPS/05HeUnAk/
882ogRTpsTD0j7Jh7SFUL95n/Y/FK5KxxKS7ZNxhDfooS6kCHpHI0J/lYssNfRVU
1Fpg2p13CkFNLTU4KJDkcw5mYXede1czfZW3IgWX4ifBYSbZxGrhBTkLrFW3VX/c
mO5bOj8xDhXjbUH9zqG6N5yyhQmbf/jbQv1cFp8Q/XJ6c8se2qEzhp9GZBlAiLBc
07ma4uPiVG5CL9aIqvSv1j8KQeYkwy6LM7HOrnPh8DfR6MPR2z8dnTU6Lmx/whkF
+auKKeYctxDyRqpYEP65Q0tjRW4aWCHIREtnJqeNhzLPWWOrP7k7YV5M2dO+cSf5
PW8sOK+USvztyf3NgOBfRLURtLBPxTQZVekITWu4dhhmEq6guIQw68hHmJ/a56Af
hS5wQ8DOktOB9x+YQZydJuWIP8S1oQuF2/UWJo3OOQP8j+k0Di9BIXo6sxtrCMaf
6MwCiwYzf/VSe9NW4SDNedIlMjjm8Blhf3LDmtXkv1rJiLQAOVlnSAThZgAdsM9s
sY+JLlOTdxmlFz9/oTa2HQAS8+l7CpL++YcoNaP8KuRjxofrmoNuzjmmm66THZvz
IYHXVf7b9L9RD/wujulVNSsS422lrndDeaRfyAM904mUVKegRx4bQg3XUJUCYN3X
icp5hpKZf65JB6rjAstd/xo4WtVng3h5xPu/rDQVRfUpgbKLAIcztPMj8zgjcLKf
dWX4XqMIj4NJD2MG2H4NEXhFabvgFeW5OzXt1+azPNpWpdy7FCGXQVW0iv3RNT4p
+Y3boZXWZZD/UmHGsJpB0B5fBX10jEJSMBXIkw0ipsDxsMpdhgwoHFUz49DjYv+m
GZSagNTFjvX5dtVwdKAafNIJTusiCP43g65+G9m6PYxS25Dd8gZLid1Fltt3Y7Mr
mAwum4Snv6LSSk76/cgm4GvWK1VGcf5SrT8DEQ9MOczqbmWWsehPbw4aQUVNe/+u
PNfh3SLirtQFrC6YqlSrLoLkd1KSxxU8OyhHjJIdsC0XPkH2KFKoBMvC/myk3NaF
X8D9eTvDt0a1Z+8MEANHDbKuhxV4KfJ+ReBV0MlnfuvcgfB8IzShkBbbDLEImoqI
mDvey2PxqblW09TzgjuIm4IHlIZjLiLFbAlQkCwyzD4o5KXugxXQ5+v2XRcFz8rY
k2aXnySrzi8WLK4fQMVpYZxPvhgOEqZrrNiwWKhIToAh8FrbrQ+iImx/AicnYwKj
74JVXF1q1pY+nEhKoMEONzO0rLSlRlF1lTbUHcQcA0jmsQxRIjMa3z71AM7rmDk1
ZcqktbUth0GqJmufXZX+KWoQy31uzbWni/R/tjybKiy1TLfyQtaIcxQK872lyFI0
EqSSZjbYqq74t0q39tzXm+oZO5kVQ2TDXcoO3i7mUqHBGln9ACLZfmwERtNrPA0a
FPPV6bHk6YOdAWO2Kp66dKmWIWprjUMeNwNkrpgxdj3kzTG6mtTZonbsQrcY9eUa
xJwZz6wmimzDDvk795VTPys/1HOIfTRLlvxdGRR5v7mvYE22+ke+9KmYbckMc+sL
iaq1IzKMgniL8VZ0R0gArZ8AjR5Y/akD+rsDzxwMNnTLQFXXH5eI82F/kF8wWRxX
Gw0PBmZ0OsprltVDm3i5yqGAS1GQkg4BDzxsNoNcYMBxxAFlvQ6K8l6TCfelgD9A
l9UgXsnqi5GQiJikXLFY/aulODFEn+xvnwmbsI5u1JPxFojEzuZlC4Z0R62+4fNJ
ijO6xUCcuABY7QQs8Q5OsgwrLZ8FYehmY9CjD/0tsjXUG3wli/Pio7/3IDddJrwq
KCVEvHZeajAkHdsgEDGwZ/XnNIDEQBxrwsgNayKsvI+/2KJ4814i/siXzeS1Ghz1
NU4tX3rPWgk3/QOgj5NM8hJpHdHvlJjJbIZi8+ZJ2JCB8riyZkbO4VR6oEcRQXxl
PD6qgH58KDDpFwDwEQU9cTfLL6JSe3J4Z2ZNDiRFMDmx6ynhf/4FhfNgWH/DjAOa
dPXPtNolRodE4ciuMer9SMRWoco1Wm/Vp0uJTyIjIh0Z3hQ1LSQfbsLMi5LbQM2Y
8aFdBTg89Mr6hekLwZAkVhvgMkbSKBlkgpjNrGt2kKn+OZnnPXdi4nZknHeAxzRf
fcgBpCwOa5XcN4e1YnHja19FxaUbImmYZLvKFvH36ahzm/7ECwvkAsQR9Dn8An7w
/MkRejEwIRm4R6wimxZ9OQT1fqckxMM9t/o7HPCiMs39oeQhHXyMoI8tzkha+m94
ndzI5PAOs3dj+M/UQpv/oXZIf7vJAAyMpcq+Rpgzxe7E1ogUV8P7zuSkd+SuQALT
zHrL939oQdR3BW24Blk2BCsi6uTPjowDafjjqWWbo03n0xt4XItm+pX/KAKPAgNL
VcRVlxtsfLA/M6jWy+7R0GjaAoYxW8oa6tcK1/HB0Z9dNC5e6e15+L70WHAY8LgP
b25ezMnS4Ufs5PIA6hx4RK7E6pKf83bMzSWtv+UFIq4Tbw9prl9f2KAgnK/FZK/o
qByri3F6+egYNo8I5XsBe3IyS55ZncqgXR+I8g69edWnBToMdyMrTTynoiSHSVwU
3NGGlZ7Xi0dluEb1gtafjGUMrna3I0MRi2pD610wRfEZm6ov/5VQHf6GD/6iPg8E
QKFUPbzhrZwFOqDE1FrtMYmDpzlnLtbmctLzL8vGUPGHZQ6QUo2WkXI38zx7tEmh
PPsVC256d+V+2IY0VCrzJK9Q006MyJBvw9o9+U5kpTvUScbk9D+SqfU81YrhGBTB
DGDSja4wtJCZJJZGCn0yPDdSDOmqo34LFw+I0ENazPLhDZ+2TZb6ibgh0YPMfO4m
tq6N+1n4CMX8Js4LsxSAG6qBmdgOMXFMfzgm7S/cYGvqB9T4XZwY78QwlHWphJHO
a+gfO+keysAsLQpsqIHhZXSUMCE7ieMA60TAOwmEt/RSKWT6sk/K0DDNv9dGoOl2
mYBGOS6Hu/5r/dhrEE0FxOfPXHOKnrXIEe7v+WT9w+z9ti+LnoJbu4Pb5Wbk6sc1
mM7nvLVPLrbf1iMhJQkzl8CCfbJ123gQuz6XEgTKVNEJz6KUaU1fV4LJv9Pifo/+
eJg91AZoifGpHeecMl0e6d673ZEw8AHlsenSGtyu/dkXLI9WAVBrxE4eOqlMhlxw
bemmSIwrvP3QCWUTFzMf5G8dUi8uJ2qIlqz1Eoj36Bd2dtAO85hIcxcuH03YmcUE
ZnfmF8mUSGnp/i8aACg/hne0Shf9zYqJZRYm4C0imHnSQ6bJPOFm/Y7815joHc/c
EdM89vP2FvO66Pn8Hq5tFKOtMn7pK8zNxYbHM+e2Wbaxb5GNQ6dUm3FQl31zymXt
Ukid8bpUa+Ya4uFe7yU1BjKBzOrMQbrkxVgD4pFpPaLmZqWQKplEwQYw7myI1tlp
gSZUUNvrqmKDs56wWRVxvzUX+2rV0KySitp3jWBice70hxeNqMygD8v3c1FreH6C
SA8JoRL5ShfCKpF3ZpvfEBPHLYrLM3d6kKAHcW2i0kwPgQK5mrxmiHtSWNtcYX0A
M4GbjdaQQkH3pyCYmKPinsWwJ92Ch5h8To7GQPuKJ3ua/7egRDo2WQ6ZCa20dy93
2mBjVeH2I1hymRcTsnTtBjenEbthPLC65yX+xIR3MCn1/Bwj71YXQGDjJ7MD0T8c
UypOFhtztr5OAjAq2uNziyHd+SvrbmwiYI7b+YjNqQmfZVURZnO/p6nZLE00q6g3
ZQHkv2/t7JjgAXedoRs+IMGL5f4L0wAiykBOzw+wA1DWIIq9w7YiFk2dY8NnYy5X
a3tPnUQxFiiD0zF8xopDIrW4k+AdMqlifcjdpLPjhS2YAbONjJfyUluQMhN4ypns
LzrVSeYTfRm9e8AOETtYhY79bjGtD+6S2ZypzinLFNJCpdmec2VZvKb1sGXlG6sI
ZwLyuayxDi9osBwXuTG93QlgTAmEOL2gFlUq4g8uP924OtHUgMeTOvUou2dWdcpL
vDLhZTe3sOf0P6/9eKpX0TX/ndYeN8lZhoIzrqqzgkKYHFLvK9id2rlQCZIIQHW2
hQSabbzNY5iJ9P9a0xsEcz/lPuYw4A/YKHFgnBvYwxwNZHudHbQPkDnqPoqdJJCW
I6k3K9Na6bRlDCT5hTHGAZVQk7NDbI3AZyBFBujyaLytq2MxhYp7fCtm4Bbfctxt
AFDx/phMmjyw8g1RGMpF5SZvHNB5/T/6Hc+beQ8V21T1M+0Hc4bn8BmBAURYFH21
fctonmYyPhCpLDY9wGH9OqJUxO6ZusXzRf0QwPBSSw9HX7SaT2OBN9C9Y0rpD1BD
5AQzO1DiaF2C5wZhSPf3ef5MZLjZE+Cdra/5T/eoPJLh0YJ+5Vj3QY8VP1/lk6fF
DSfGbG0FojONnvNSVqNgh5W+QVkW7+un2woZZwCZoI2RMkL+9XLl1iJ4DKa6OoKT
iG1PgAd5UmDj87R3l5ESwe4kX4l8zuU0rR8uKaG8VSCb/VGngY/99Paok3TBiL9I
p2ODxqxKNhLRlxH4mlGbJwZJ0RcXtAlLi64n/0VuS0Vxnq2baWbowlo1+yx1wrOO
Bqb//uhzzpaIgYZk2bx+2EheAJTNu0V9P3EFoABnqkW+cZyb+b0VKzHhdvo2JDCc
+TGmLsT5cIxpuXwLGPcIFvg71RFdU884bh/XXK6xZISiwGL8QgxgQPx0jPqkPGIA
I92hzUfQ0Ngzbdnfv1uGkAiVs2vwAGKnDsM40S59B4YAxrDGpMEJo4cyTmB7CStO
4QlzvYHE4OXKFUutB66b2/tOU+uvYPnIjCj31mIhzB9wLd6cn66mHyTski82MSAv
Mw07CaPlj/tEhP/NkdaZLrXhxHryIxgSiZyIfAzsQX38WzxX+yWfGp3SvgpL3hQY
ao/YvrksixPmcj+44n5tl0t0eXpMGTU7gMe/XEPcBqmW260LzXljAkd1kC+P4uKj
xzHWYitLi/5LksJI7qe7I+hBGZPCRu5roPKfTrjlNxg9ARXTAKv1DNKILvkZpWWr
Ri1N5xKxsBa84h2hjP+U5q7HZ7rTzdDgTr30pRZks/8h5Mxi23+dOPpW7MEhvjPA
DW5kzX5L+HSpZ5sE3W+A1zlhTFIWQhjjLXcV5oNfWyHP2k1KTvAGD/IMBUZrsomu
zOd3UtkCEFEa/N4uo6KGRPlDaYuDxCqdgPqbe4NFMcGcVyMi9Xq9d4MpRxVjrrHJ
0U2RvdN+d2VXMBICozR5oeIacej1TQGoqRk1tW9O6SAkPHsJUKRIxQUUzTxfbibo
CN+DoGZl52ZtXEwlyGLfEHn60bbYeXIvJGF+D6qVvPpannKLckrpVLY66uWR/AGo
S/BiiQkPQnmtY40uh+rmYkh69+M1/ZelYOlo4h8g53YtP6J9UfZmD+pZDHfbbNys
VjvMLLCQc05ioWrvE5PEa7LFz1x0ny7o4AnPwas9Tw9EHEqudBld6c09903Im+vS
Da/xV+EuPwyUerBzfBci7VNzsl+TPfhDvIPij69Ee36iVx279W9vtcWaiFmnewKC
f7hNfSxGmdVk1B71+UgClzcW5Emkv8UTvP0+5avk18egHDlohqw546rqiJbpfwvL
FDm9V/YkCrvztO9kI5oaavyTvCTRT4Eu/S/FnxRBY9ZcEe7sXHWf5cg94AwxjHSK
92AB/gd5orowzdjk8P1KAzKoP1i+SEtI3yo/2Ji63l1zYbLyF03RcgYUuQ2634I9
ryLYQStyFhw1bbNavm9rWmCjRKw4SrcX3OWlbPR90tQiU1O5DuFzsv8+AyfXev3z
1jls/KpgpqxAwQdP9Yoe6X793CUY+GA1gujsAwR6AXwymj+V4Msjy8otW0wpfztB
00ZycDYWiaB+xYoAB2eZwWveaNHgfLSp0JqprpAvL+ZjDGOnLLdRYB+txDqsf8JB
4IASpsbRcINC/hOxz935MAxhyH7O+jLdZiMh4gaYeUWc8qLtlIxvmPVlxDIneDwW
BZ9Zda+ZON6DcdddVPiW3bpyYt1WlMMysSmXkWqTUZQ+G5LYaCkF0h3F+6tVOTPd
afhCeJN3vFymOGbfuEscyC3SaABu+8obMojnqCr/+wgpQUNyTYDI3FTn/D2IU+M5
e3xjprq8rwopuBcJ0zi/2KZdDWRI6PQdKm3mqcS5owhEn6+LiorQrA3bsDI3Dd+L
rpX0J5Dw0SkV+xMibmqXQ/LyqGmuSMcRka2VsAwt+WXZmCOR1IIIKIS1wMjD3qvs
q0k8ovEd8Ibk6PV/qkYOgIambTZ5mJK7EDzEtxPw09CvRMnhX6FqdwkbytyO4euq
cAwzV4XhTtQprYyn1SXM7llbdpeatV2k8w98jM6AmvlZr/Y4WO5TQZc3ddpa10WG
wMpjn6OrhHydqM+H7+1zmw2cbQgO7QNjZACTQ7jq5/4S3CCUJMhCwmuRP0b+wK4e
tcrLxT2sqlyRD2ymgbzfeVaE8V7ixJ9htUt8JLU/A+5hdn8qMQyAD5dhMgx5VSsi
7Wsx4R1KO9ZYglISaSUB2DEiUVd4U1f8Cqc1URssISSCp3xQOOFZp+078lGRaXGo
NxT544SUDfefDaQHMAXufmZpNAIFAENBAWzNHt7+VXxmd0Dx5Gf7aGVuIsO2TABF
kvPsg5gNJz1Rx59jn2Mfk6xAIpQfM790aYv3SVZZ62dJgRs/zlIhGnJ4hQLX+Rqb
B3RT9Qz1nC1aQnBcU0h43056QkIad9cgDkAg7eZUQsOllyiKB1TQy4pm//FuYNJ5
GieUYTzyZqCFliIVET39MbGeTh8elMlP+h3Zzt2DoSCpXny2ofUaiPsSJ1xzjg7d
3az29KwR5dqvIVplUwTIrJKqKoALqtG2Vqevzunpt/RJb7Y5Tr4xpNYL80MS8aKA
77DMOGvl3fNeBQmJtQ2uEebtEL1X1301orv3rUJXaE4Yfjc+Mu8SPr/nUeXBnhmS
E2u3EEvlYeFY8qMkvvolTLQrlW29hWb1vrZYKS7H7caIeitO1DGM/Ca3Z8WR+xEK
ultQz6V17AFmn11sq96xdlOmaMqOVKQ1Z5mG2eT4J3gkeVgG3MHaas1m2JKMjoW9
sncLxP/V0YNm5oORhwlF45M5EZJKJndOiiXcZh9zwUSlhyJhJylTscSn9nP/7ZO/
4JFyCIsvhxUNzGBNlhCUz4+vbYzcJEjNLlP67+zEdJuLU3He//DRKvtcrxHvIZoZ
PIHnOCtoFV1298rYbTNjJbc2PxonsOXxmT3Refz4cPlAEtEUWrde12hYiocy6CpH
/R4ybGSo14uZI9mumxpD8wCRNI+CdPZwluuSZ/9/A4BG3HNSK+W9j/o8W8gsE+WF
xQrAB0HdlOAvWwOK2NlSa+TzUG3BaVS5Oit8NNn5EyXlrxKH25r9eoN2RHkYaY4Z
bo+Hpa8WZqtonZc2yDznQZZNWw3yEvYLq+6OlDk4v3uajwDRxG2K2epqT5LExZJ1
jyoUzVqVFRMhTboWyAIMLSWJL294p34RrehMmlpUBLi7DeMRBIolLAH/trMHIsq6
Mj/QP5yPYBVyovYIeIbkLRtSLqOV5lIjC864BK1oO0fliv6mHwGN+y7GPo80dLmW
jc899kOGeMuXluLoCH4DGvKyHwxmbeuaFLd7xhDD/kYpgur3Bthy9L8MJJo/ruak
tHwzyZgFQyrHAlieoCfUrTzeaO5qg+8/PiZ3owDGtUVvSs39j8Jv3E7scDmQe5o/
eXqhe/StFYavjDVuMmYymYrS/R61+1QWqBAQpHW8ebVXpIfuF+ZkBj02zJYDB+9v
Ts2DRBvo3o7VdNFfGBRA80uh3aD397NuxNP3vnMvdYoYmT46QVM3D4wtG2InpntV
nS0O1H28o5RX2ZoUGcto1MF18wpUK6uvViJsOGCCwmXBqZoJ3Hk8ijajyys6LV2p
BzVIwe2eB7CqNomp901fNl31rAciH6zc7qXeuuhUH9LTEQLhQR7ERZOen80XHIr1
BfYJRFY1c4+ihz1kRIpXz5xqvOcJ5pPW3bItd8JBVWAhdxUgXNRQxClmX6fOWipu
Vg+tFGYhShKSJCFl/yqUyMU3jHYdrh9TIYcQovZPLR94Bv6sXpjgRYhiitpIVsuv
92FLK+r2y1d8vXeu7tEHJE7Ovxgp+ygbvemCZrRCcLUAFJi8AlNF2TPzc95nrgjy
BHhvgsh0+b1crQlZRT2wJCYEeYZM1FEX5PVLMrwlyf9zD+eJhU+SiPs2IrtwoROX
fQVAAggKztpcO1RviBSos1imufVFxlULUpiIxJnZK2AmFUJOc7qr1fJBDl4nrZOv
gUZHeQumWo5Sz7cTcc8EK12kYYxRYm7rI2psVhwU76Ur4bxtQOybjkGzYnHSpw05
BdHZcmyNLSKYnxfzCYOlaCdUxml978nUbHrjjUdfB32fG+UOj7GKgZVJkSvKHvMI
gxOdwc/yMEmtXJZVVRylG//A323zUY9SSSxneQHfrbyOGs/AjTokRl1gRPnRC6zN
n91etYHjhjEmqTL62GwNppfJBxhgP4WvcUnaCL3vJnv32ooIfdBCQUBWkJVpUkU4
wqRW+yhZW9TSmPz4QiBLD4m0RobClw93jqr1t+K9CrKDoNuZ3vCFjr7n8aJWN+nu
9jOEWNgSpFvQf0j05B+gMX9nzkDNhvSHbLgGFEn/P9/x0DwgTTZnDfp0w/5jEcJQ
7/tyMPMnSTqiLu/C2cY/YHC8ZPW3zWtnZoWb48J6U8eMtoo+15+wiarjItIL0jx1
6+HMAcT7l5eV8+hyE1bemX1NUcC4ZCvnvwRcdP0qnSX+WVdmClsCgz6J7Yyl12F1
d0JyhgT9jBcAPTJQlqz6NzRvhMMvqp8sdvwryXJEXQk9u0FyHcaeQZQRZeI9fueL
Lpehk41uTjY4F9hDTXs8yiEgqhD8WqEy/Z+xKPuyCtlig548lUGQBiLcXNDVplBO
jcjosbBN0GlL14YbqEchwARebwWQF+7F0v/Hoem3NG8xtz0r8wb02Qi9PSDEhXJ4
o5WlL1thEklaZ7y34WUGO+LDqT3zpfek1j61ZQeQ0yhJzdNxM3ho0I+YT+nJRbfo
8vRrTUfFNcGh/5+4eQm/LMbAES64uxeu/QIl+s9gupmLWJUnVBAe0FL+B/KGxZFT
kx+iJU0cXtAnDXJnyV4HVIlpG17lfIKSjImmlkCrjwN+Lk6N3dvdzHbWTQiRyJo0
AY9pKefEmSZVFU6cnlC9Gl9E6IcQSS0srhmLbVdzD3NntVjbvVcJKqDhjTNHDsXn
cFrfiCkPdmX+huFlObLLXKhK5j+FC79LnpRXtnfxkvzndugBOA5dQxBSFQ0mN6Yf
uhZwPslf85RxtOqaTg1b0MVyGbdlfuer+1r9Uev13CqEWgU/yVMBMoXGMMy1D1Ox
aGiD88iSLGi7J4B4PmQeHsSPynf2lpJZuB0/NCZA2rslptdu+sXglonRq6svo/y9
P5MRU9/TXWhD79hFa73jP40RiHVRlunQDwgYkDeaYOq5GJC0uxLUSMN1+cfXX6Ke
XvxNLs6FeDOOpGs5tIfjVDivA25dDrS1tURXedkBm/HW2t8Rf3JGqydzDnIbV0sm
c87vaRnSYtii7sJnGw5eBw/l5RlRE87mxGKUJNnziaNLQfTAR6+XcCRp2yeVOdtS
8th35lhE47lBrWlR0zA5uo0/dg3NihcRwCToalw1ia/hzgR6mVUTrXbaRE1BNeWb
SRc1DSNqyQVgFUxeAyHfSpmnU+RrmOc9vsNs6aGK3GRP6lgfXNvVrlkAmzg2k3A+
bA3fX+XuLZ2FbaiHKjYARC5xyDeBCsGS5oPJ+6CRbC9tKbEEC4ifNPWEBR7VeKrn
ISJIfZ2EIpnYcTIzJo/rjpat+WHiHi2ZYXuS1kxkedK9FN56/c/KrhBM2lMFlZTm
Ot50h8q3QjMltnlyuX+krxN3H/smjUZgupW2FfRSPxHfWWzGAjemOuvWdYP9xd4Q
xGw1G9+W58ZPLrKsh78divd5cOBv90cpkuEoL+5s6JQxlSQsvi3gseq0nK3L3Y42
Blfti9PhA/OC7Jce8UyuQAHN9aKdDfTaBM2RAQcwDvqd/9CKb06Mt94lI+yMWGFt
KjXX4F1gAk98tLtKLjvLHZN82nAFUFYWRLL/vt5m+puAw8K4pH3+IB5FagIto0Cz
JODWE7a0MiHozMPIRb9Jmt76rEfK/yhVsCNai55NxRw77QtTrqFCALC/t5raje/y
uO6T+X1V7Z263ZyF6f4l+bhMbCKbYqlNn8KENdBMG4PAbCMOuTNV6vao3v/8QuHN
4zEdnKxYs3/sLvX44ZoQj9lJTJCYgl6qLaydximnP6Tg4vCc4sCIQI6vOGuGPIoI
A/7w7u53RfZqKRt//VpgwY15SnPas7jfvUka8PV+JYEF/DLRxQS/KZmEP5ZRiBR/
M7jmsF7YRIphqTDJPmBunSNYDdEnOelju9Baa4zs3qbszlYMZPFrL2F/M6dxYybe
p+OdAjyC5ilNS6TsXkceBx7Z3k2TlWJNDicImlNJRk+3MYJe03FSjOijyBLA9Tdn
U/TE+4EzFtqRVOyTa8lgcle5KdXKtsZaScSIdSIgMovzfzvBN1CLVLoNGLI6rRQ7
GgYwVZixDm8kMrGTZ24JGKXk8oQA9Tg/3QxX6zxv9aOIyT6jW6xZFk+3WP6Z/H9b
5gNxeJMqESzrqhMcfXMV8R8Bmz9E/sZvBCF9BScPTUkCGRgICvPjwj9pN6YUIq5C
h+oitaXvLmy2wcwhuUd6xfill8GjHr745zhJGF9CZ3/JMTaFv884J0woiYT2A6Ko
bKMta4NCxv15pFL9+FmIYVR7BA+Ez50ZgJFa60fn1dNlLgtty2jHuRBTiH4RxaQC
mL+9kk2NDUG/+4QvNo1ST5Okm2B75jLkleEkk+sn1KOMd+EjudFewgNqHOdwUiPg
tJwvEiyyWO2oDRShLRfEOD5HofBq+pHAaKRua3V1gYtpdL15w0lFfoNV9wt2r6gw
iOL5iWTqGtpU0tATfv5bQDsT1v055zuP5LliAqXP+NNHRkM1z7N9VEzoFwGfOaga
7kYvd82I9VC8xxkdaNRo3R7pBOEyHHsja0pZ6eLong7+poQrM1IKhhL/h9DDFZm7
ba0hJg3rQvNeVj7jpi7P3d3RuGEDOvyA92CAz4WB/kIDtl0wh6GQPOzUJuL5YZWh
oa5YMDCNYieJqRsyjuDzZO+8+/6dE6F2w4kQlzzNHVuh2gp86P4UHNznf0GJR7ww
qr/swBpXc7xu+jonVOUFp59Zel9s2jf5+DSJs9REM5rsk+fLqafD+IKx9HMTOIJK
VOJ27PcJKkcu1HOIdw/uV1LPMAnvx1b4TiQIW2ShMPfkmeyRJxfNgAvxLCAuPipM
9sauPmbiCQKn2Y15JfWIdPTEWC5o0asfe7XxEL0ZopDIssxTWOEhNn+jmyv9iXmi
BnVrQtwQnSTg3RynXry/TQyddgejJ4PhpGsv9MIK15JV/pPoH0MV+7bJ06zaIS9g
QsdKT29Y0YWuV9+DKz/mcpYqwBAblsKA+QdxpiOzTBo8ceJPyGnX9bpGL3Pj799E
EI4SI6niPDzOFHOxmXbyvr0wXeioGX1RGjpnalr+giZjvStadAZD2nZ2ONE96wCN
I4vbA4ZyJ4AQBuPfM6InREPHEbM7CEn8dD4l8DLLsgxJHGitnVqRMbpXE9FPODDu
2yRvYcaqPhgTJOOd9ybWLHkFQ+CO/d7g5tNzULsbWgm/jSB++yEfgIFI8PNfJ3Vy
FYAK+QEtyjocrDnycTZt8m3laLva94d19kgJZuQ1VzpCI/Cl6tN4jB+SrUmhkLU3
t38tQKct7dOI6bR/PFjOycKOeuaqwgU3IVS9s1syGahDzFkeuiDn07VzDQSGTh5D
t8PyUVhDey+6jMMKG76o9aXdF2c7ugnCi2jiMMBcoddOu7JybaLZ3MQJrpaKCR9G
ey78zZoZYo1wSxquf8XDhrXL7Newa+OrQGK79e5SXnQh92VZb5ls2AAVHqk1EK+X
3Uq4z1KbIC4E2041EY6G7cbCxDxR4lO3AhS3TvlRn8SgrHDnANtd7t6EGd8LJUPb
064UVi7OyfxSmsYyeX9Ufl7tutFT2bv2UPlYi6NwuJh4LppmcBMbKMVU2n2aCrhI
+csCPifmU+wd8enmCH+sLEa9g2vIsq2CFo8+gUEcYEBFFK3yynYxU5SwlLULFY+R
as7OP7gCKyaYTXLJqsFc6akJp6VoYhQ42Wrzm9sFRAHuztwHmchT/gwPh17o/OKn
cCBViyNMmO5WbGW0VNpOcnYNfiobCfUoz93eGaEv8oG3mhhOdPi91gzzI3s13nIV
9aPQGMONv+2DzNgEzPbBpSfYRA0kGiowoYcfO+ReGc3KiorA169J8YmIuSio5tDP
bM1ds7vnHCXpS0HkCiZ28q8tzYupsvjoiD8H034TkXXD13cQp+Az9E0exhfjrzH/
t8cQqvgdHRMhHom6JwjiflLcSyyShkscHVYaWZY8xTlLTooCMqoREhyhRvVTTNAU
f6CZMtyb+fScRRjUoyjSpgUGnhE63vNYGqDHZVOvP4kSKM0iWbkYtefLUi6HzOZS
6w/MQvIATrAHtFHTjRzWDF1d0QjLC/tCnNQWLwtiFncPKsv2C/Dl9jQ+UsXjgOBw
QmlZZ5tvjZOzb0DzUHQcfUseTXN2J/u1mR8h12sXgH4mv0fkVmI6LIU68xKWsj/a
uWi8Vp771LCjYAoGam3YCe1tNjEewlQS1XTmc5gBQHXejru/4y2MzwoJjyoQ0Pqp
eIK5sR+WGiPVVoKoUNk2TTQLLdU/fBjS5cubSii9tkNiZzuACkFHM8EC6A31v6D/
FqdKFVbo/nZdPAX46v2pWWpuW1Cs5Iyx3YGb0g4LT7j0LE42obNVHoEjFL9h9zMh
v6N1k0Yb+B2TbVKtnulKRIeSQyoAVq7QnWWsyQLUiWfIzgKmMjjgJuCHeNGxrmxF
UUW5qNKTCYl8qXCwNJAqPJAxMJY5aaHZG4t3VR2eL10ysO4PldYwG50K2eGth2p3
H3WecxM72Vso7F+TphS+8f2nJv1G6/8uTgY085K/Ej2eS80xlXZJfURW6CEZc28y
O8jrN7f0qxYnAeqlVEWuXCLYKkYzIsnPGTs4U13BNZx5XmQ+jC48iCJ2yCT/tJlG
ylF1j5qRMz/00lF1wqVUURq+TUW9H0mreJVcQx1Kld5IqW9JANVDGsZ0ZWjxzn+h
wnXC9bEIGhAqvflHhOI+X7s/O/tMqJaYw1CpOLeSPYw50KVKdenzi/w59QYVKuz8
kCuWdMINOB/AqPuxdg6c3cp9lDTR+lLQA3hXqWRuxKcS51Mmu9M/0uhXNcKcihrw
duHkaTrOl7uubSPG9djM1qb5Hh487jb8fyl5mKjSjDOezGOb3+FrYhhd8sl/yUIA
+BEsoN+uvb1vQe+69z+J6g3isNWGZJGKWDkWPXFpLPrBxHDA/9+fYU1CEQ8/6RTK
2iQ3iH0gHPOJhza9be336wbNh7o+8SfdzIR5IlNjxLnIInhjIVOaYDSiIYIrcci7
EEYmGeHxGHAFA8/MnBzXHfdr6W1zR4xc1lF6wI319ZXKtjkISKxl9nXz1/ZYcuF4
qr8Hpzq2hi82V14nkiQ3CDpXE34mahuAwSFYSd7AQyNGxTeYzKSmZZq4/B9Qt44o
35geR13VU5vcZ9Mkbm5VPw23pLDx2FYua1KxAYTRSVl76OH+xLYHRXL9MZIcZZzZ
5wJ0qy3CuX53fW2WKl+yKh7MtaD284pv+/+o2kAJl5o8d5I+RDSCHmV15W8vE2BM
T4jofca7Eodx2PjDFy21yE8xQbMGWQDMCB87bEOjM5bq4NO78TgNYO/GpboNMRKj
WKCO2oO2+6I+ryQ8YGP2PK8e1O0DtUy2XNOvRKyVmXxU9uwGUnbpjVhzdmsGPDKb
i8a+8MODKK6tYJVG3O9MtQcPflLvZxi89OoIf3t8EjrGLwqtDNGC8IDQ6v1u5N8I
cPRz1gFNFnrEwyip5ArwryWB8J72ksHGy5UQhhGJ2bEviOtqC+4ERIPD3Pgf4Dcm
+yK3V0+8g5fMQn9cVWdUO1yj07ALBlPMGoCXBUA1SleUQsypGt/XXSPi3a5FaerD
481eTkz6RLPdJ7C3rmwPDTmC/S2QKbK0D1YIRu0upgvY2cpQosW5MxwRBUS0wIys
8i/9DPWIXoyW+q0nK/OYv1/DG7HyPbNRHzUDmIiO8hAL4RoSZRZ6R8iz+Y84qIro
OYli4oGOQtcKNr7FSXHp4NQ8R+cAspcBtrPAm9fmqY2hWIY5yoIoGzgQvhc0ulKa
5cqZy8SXvm6ULvCcaureLr4/bugDd7bJacYSwtx/6bVKBBEe3VTD1V7iIvH+TbXr
2IGcErQBAPrbvSOzLsMYJA2JGM027kiFygLGaGjbgjz06aLdcp1zUd4CDibqz1xu
oVZwls+tAhj4oWyqaWzT6lW17cliZECVozVkf09KEck7twbRJNO127q6WZOfu/tF
dA1ycFR+PpbD2fvDL8KEV4wSIeNJ8yiOhYfs6k5GGngAucrdA9h61+wWykfjl2td
AxhEnBRWnIeb0sZ3qX+/6GFdDvCtT+9eXj7McOMtzx14VvhNmZC0xX1tdZJvq2TP
6oL9l3EFzvCrkN1sgZshaKJPq36XzivtW1zr7MVipLx+z7cLA5BRutXOoBc0dJiu
RXGwZPPrzDhQyhUu7VBP6Q2rRG1d/lffMFefC3MtNNFyXtq5PGW2gGzJpqsU+ttZ
gYsJS5CrsUHF5Dns+yz4de0/ezoK1r5rJMpW1JjJ8ejXcpLuuW504VX9YPLD6Xez
8AWKvr4WIkXn4o3sR1aPTUEQT+Ykh4fIFBQNRvAluVeUs955td6GtHOYS30qsYew
NrKiH2CSYZtGFXF0ZmaEIYSbNKmk0vZ5dv5fngzNUiGNMn/jwz5qz+BkWxXnaS82
KdJTZRPEalS4RTSVXn1VnQbbk7NOZ6Vqj/YelrAxpqlwlTUU7J9KmGPEJ5bnR9go
Om0yWi2MI90JtU/HeeDz1zdHWCQfsPQW8p9GvHDec3wcNSS8t99juQ9sCBVkLI+m
6q/j0rR6VfheTBhMNR5X8ZsrXa29t+WdKVjxvh1ZY/NXcVOJ+p26i+eP5t3gQqpS
gRIslA2Emj7UuGjGonNxVBF8CVN7+oWm8GcGThU0fP5c2Yz8kiHl5KXpgc8Dq0fN
ohgHa9yAL15QmrFy1HIMcT4goo9HopHSWhWANpWrb9r6N2QjVOgShHDsbbOF3Bqz
5/jQo4et6MCApKCqhRLcr+rYVvexTB4AQRAPn908D9Nzk6rHzJ7fpsb9b+zFCSAn
6f/ode4J7acc5miDf1hE1gx8PtlNCZt30XIVa+YJCkR2yVpr0kMCjVfgVXHwMRhx
24GRx4SMxdC6pAIxIuq47ospeRUTEBbqUFc3rcZXzu4XhdA6wo9mNYwHepcf7BWu
JUP1GlBr7d5J9NE1gI7RRPA/ua4YS7Ivf8zUg9bFUykooBCAl1vAGPlhlT3eEvJB
C012KCRQDddKkpqW5t7332UjgP9bm8n+lpyiFBO/H9ODvkvrTxQT1w3/Go2CUeO5
ZY0p5yiLPH95iryE79PFtsaALST6ifOPro5OD25qXEv+p0dvZC85e4uxUgDW8f/R
GCmsvvEpLhIgygP2+oQbPERViA3D2fz0+bZgz+xpWUxTVMry2MmMqmFug/hxAwtR
IIgolV1qGklZdR0shNg7SrE1BhU7eNpdCulMHrTbUNyVowCXea7Vbdus0IeIe0Lt
w+72V1MAsIe+VOd1xjF84xYrtfIOzK8PexmfbIEHkxENJT1LHfwLIIyRNwwFEJt8
VxRolYpG56Ssi8ztit9pm2BDpvA7Rc83U6zf4VgTye8G1qOymkoC+s45WxTHq01i
TrWws7Vi7Jc2p3pW9ZcGvZeukkhzwNlql6/ffG9i9V62MHHee9DUNLfgqCgy83fl
2VqvYsa8Z1pGlQoJwQEb5m8OUg0y4bT4GE5rm46EantKJ/IjcyL6mXyxCpktZZYX
whcPrDV7tLHfQ1urQE+ASzYNe4GmXRSMKI2L+JZnNJoHEYNcXgEFPBCypXPL98Pd
pXtdOdXnOL9YsnPa2NisUz3giHq3XHmZ178K9PGELtBm58NW5Ax25HFFPC0Gwn9P
b3UxZ0w7eUSxZ+6iFa4k+aia4a1SueWTW7BDwuYRLUDQMSHKO1rMKHh4kd4J86X0
UbtU0nUfD4t1PnbIIFJOIqqhpkNd5ibT27ey/ZeswPLi44zL1p10xmGeAjwAN3Fc
gZT6Jr7TdhVAaSts0wFsCCi54cWWJXwSEpUXLH1y1zPYLmQSh5GtJYAZfBNmBVdp
j17lxWR9Xv/wuqp1bWAQtkq8QQXKaZgiANLx/1+QN2OHsYU4ib5znBryRNh1nqUE
EHYBiN2h2vhDUajKqVa84qXrU0LE4m9dr/+aRvAGjgEgIAtLtOZT3t2BQ1raTaUr
9Gx0xYXOSBIMj2x65hvXHpBVTPxTa9jbbVZjKHp3BSz1/B1O9AFu/y/L/9CE7KZH
V9drvK08RjUqw6I6Yqc99SyQ4RAEZO8s7NWPWg1ArKVqSzE5dQfxt3SxC6ueYsdn
pKomD95zrkrdWtSnseG8aPEY1MHSLYzTztFY8Ym9ftW/QIqR37YJ5GAN92sDl2Ex
i0/+otFyhALwTGpVnLF+Vi1Cc6gRdqrR84rUhZS4aCvoicJIU/Zqq/JXR/4XTa0V
b/zQtFvWuC7D6WzTN/FeJTk3djm9YziI1rHpi52NxCyVuLP4POTDPX7bWr1C9c31
QkxDnJlsIUCV1BKcH/5nxZfHWAKWkbnl4xm2ZG7lk/I5ormuZycCDxDjGerjMpoj
2AX4bByNztxsKadd3pa8OLQYG4cY5O92Sj0imQYQ2e3kH+zdNXFWzZ+aR5I11nZu
wk/ZmsHcbw3PP0V05DmTbu+UEpFCbr2YYpaXf0Siq375P39Y1OEeMmmxPkxSylKM
TVR0tWhsLGT0WLWHXw78ysJHUjS7qXqu03sXzvLOpvuvSvG2yLeiM+hZcWawlsjZ
ksdIRVRUqEsbfx3HW5ERKm0wq7rYQ9ZlawLZJDuvOCfX9Zx2ILRGHbn3lDGw62YJ
pvuSymAlSlBSCWsDYQTVg4iRTDEL8q/o0Uo+b6G2xjwERSvbAGm2NOgZNGv4x2e8
fww40Tk1+uak6At3UWNaFt7Rh6GwcDOyDvy7HnarVgKSJTa1GUbIMxmxUxidKWn4
48lA4jS8w8Q+Ax+AX6SwNT4YjQa8BrmOUOQLzxqSr+bmV6bllt3GgN+5mojem1zK
4PBwPRNOdfvh+cQ++UUKKtY5YrVqAQzZEMj/aysG03RLI/d3caHa8T6ndjMFQX87
3hIIeE2gQPE+LgOgeF+YYyCmLUkXlGGyEes/wrsggjiOiVivXZ6HIcGAAEg4jGDw
1rTA51z9begzcVLC2a1qp4SkxI6ksBXpSPcn9hBBljtHDX8BRHxSikSc9rNTgPT2
NHiVgha060hxePALBWLnDzKlNUnf01JLlTBXF5d0kbhYUh82p9C/f8X6c3h0HAds
nxyn9jgfKds0H3AC2PUovKMycahUEv4c2Mcf1jXIHx1hHfQ8FXZqsgWMrHtHUnoj
5yMMXjHQ3pfAvvLR0mf+wSDEUJqLgQe08IGWPC0QwgJitbanM2LtJElzu5Jj2hfK
ZfHeKx8jUg4Bnez6cPpZtoDMJr6OATxv9Jt1Xw2a5kEPBr5ZjrFVCiQ9hyYHW4Ml
tH2W5IQXUjvrj0oQNAuGTRAzzEmSmarNA1lvdUWpa+mD3k3aD7/Mzu2wDku7skHJ
lLLbRKvhd435IrqJaH7ai+cHd0xiSk0Jp2zMAkDTDhwXcpCeyEd3fzZ/mwqOFcB6
xpnp27T/IqFyjmjOQ8EXn1xb8pOE2GjtlViix0B2JMOEzB0k0aakCIHFSUVzchdg
GKPzpTSKaqn/wnU7gK3UguMFqnmHfNO2SyoyO8xaGqxsvN8DcOBD5/NY/b+2pDrB
F6CKiIH0+Q8leezqosAM7Ohf34SfkGjA5ZZqt3E19+ED+KV1KP3g0nJSc+Ohyh2/
JfNDJulnUPpjbIv6BBeiQvRxl8TFIv97mdPazXJFhOHio1pjqVT1DVjIspRQZXvh
VvSvocRNhnVe4vlivWU/kaEHSzLgCfQMa4F4RtNz9A/hWLtd68U8HJjEyReTybLm
hHmjlRI8nMTw8ypKm3dr7QF9w1mD2T/abYEfb880kAjp+lgRwz5MXaVd8Snyngnh
obCD9XCqOUM/Sd1yBv7EoXUOES/lLWB6Cz91TBAOKX25PUDFhERSS9tfm2mU0i55
0J6+L/r8+GsVh9e17fZrOsKiaR8U4oKnz0sHPtyBbfZABK4KNSs1kcRF//NQVZKh
EQFUpYqh4C+KFxwt5H7VqJUHDLQ/4Dbj5RZC9QwZUJNurOsLYCEshXzNPJtCgcBv
0JP1b36GLS4BaAdpactseI15VFGe1yteF7XyGmvHT+NCwJyOEH6ffmwLKHrl8WDz
+rOlEk5rBZF8jokJsKq2bgilLosJXgRiJqsJbBO5M0fbCLhVfpD466/w4yeYczef
HGsBTH1hfQydBGuIPWtb4b2StcAr4Dfgx7mtlh7mPnnZx/ckoyjqoyt8HxA/tE9p
ZJ0ccyc2MgKeY6PZKbBPYv+NsOUqhaJVmgwwmQEv0Se5B9h9hXoO3M1HwMldXK92
n9kkxuKv2xtDybbEhOgYLowpoQ0DYDeQIY0ZIBKnQdNJB+LG0/7JXh2KiNHKBPkB
AKOT3RCYUo3MlNapMOejQbQREpg51xexB1DWVMmXxII0fHPsqmveLTdTZL52d5Db
Fq52QeA9TnjBgs0eXhK/6ttaoTZrneI0j8GHiHwI85tRbnDfOV12mlt1Z0Pik9MO
tuF+P/N1zKfK30VjU1P6yfWY9Hfcb7jD0HvJS9/+wvgZyfFYfjJf0hhAUCGkm8Bz
ZbtC8atIETIngGyLHIpoUiqQK4vXXvakX5xV62KZQVBQ7ACQ66aXWnN4pAQVcmPX
VD14arVkvAR3bHBOvYerZAEcrnd2tHRLU2Ea8SRCO95EECml5o8vSa39yzWFa9fO
udUlUVNbXoEC4H2k32XdMKx/7bD6ltd1tAO0+uF2xMZEF62GBUkb7/TgHnDwcIGa
gNjQCqExQtLBH6S3DISUkADgkeZOKjQ4bfJqfgu4LaeqXrKwr5c7D7cT68KCXt6c
N6UbmOLvfi7Y51iX1B7M6lofNPkgFQUsEluw/tClK7BAxWPm81mM/iU4s4Eg8zPf
HVnbMRw1h1X5M0r778pqqCiE+fXTZfwIZ1hjsfAhbFqkdVj1PwJGEJm7cwDlXOKE
Y2BvP9+tg/MfSozYjlYN3iCtOY1YP9/+cZgzBUtrb+5SGx6G4JvcM/dgjxkXJq4t
Wpf6gUnniYJqf+i5/Ns9jsn4vX+/l91DAADe4jhaNOg7T6IeCZv4hx5WhyhtIBcE
J+e5hxs24ioRzDZxWchQ5ONT234h6M85JmVr8lZOFjjO2Sw3dW3SXsQ6+2u2UTdH
OW65ck+uqgx71Zfx+P7+9VQiOpSu1ys4JFDWxuO54LuDlG//USs0pG+OtLrY3vzU
p5APAK8Yny/bRekhfZ+bUgR8zLGvLsjlaTqKwQdv9wo7+F33drLpOOO6D7j5O2/m
zaV1/ra5Vpm5WTitrQtJBeh8BKyipN+pUCdlq/+zk8WvOoiGBUafBUexoWwRovG7
b2v7hUE18jX3TiI9AaYUbJXCrldl2qNuF34NktJkGsttkqNtSZhr2bWLipTsoBgx
3Wv8gTkl+hcKE9dqdI0LHpRTZOGqfnKymjwst04IAH6m2wTUzJDMsh4YslMpDar3
5YXZY3I6qaIq8Nu8J5vVI7r8g9bco2NSyP7/tTiD2rnknQky7p8fQWU6/CP2pfxs
qHPCwRuuLfkUCywj2kOV7H/JTZUDRAyeKoJyhW9yXchQ3UgsnutcsIk1gk0Xicnl
QOTa5yLIdQPkIBctUgbpkAjJKC0Qf7La+FyuQGEA6fnWRBTKNU/L1ygMZoRds0Rl
fdhQfNEt0wpbPCVr4Bcjhf5/Cn8LOHnO6ZsddluBHqj/4LZJHZ1VMTSgngngeJAY
IPu0N8PYUHcNkBlnTXJTysJ5lOTHcwG33+YWWpBMdMGokWzEKXo6WiARMLZim1Tb
St+t6wNHZXU73c3mdCQzL2TzoZkp3uorP30V2XDpgqWj0wbpkYunomaw5mAM8UKM
7t//92qJqsLed2vvzi4jTNdlHNXmjlTiI6hMB0PjepFJcGN/b95DLOUeyERymAMB
Fa3lyE2MRxrWWZWYHH1pfL+ORZVHbrtIWGJY4H8lNunw7gvHiUkb6R1IIqI1Og2r
fpSAzZd7dztzp+mwmP8jphfDRmQsGz0nQlHkJFOZK9970qksYvO1hk8a91JwX/yX
6T02zarQcqT68mw6tatL6gWQc8xGvzMqBaKeKo7p+qe146K4TELhLoAiOt1jBCso
QL5U39Y9Otdy6HrLHqBawDeLTI040UR0RckceAUb0QQi34lN1EXZCC066d1w8pQm
ExAu9zolUg5ZXva+AVKhBvCYMehdmi83HPlPDfx26GwwSxgQbjg3cJ87Oi7dK9LO
fU0j+Fn+BIhXnBuDq2KpI9WJK3lxdMSzF810DhNcgPgn+2EYktTRSU+yQA8z9x8E
m3n0fItw2oS4yIpjN95Lex0VapzOj2+QndbJ4S4QPZYnD/1NcEL4ogyEz+DSyuAr
4X8lLUlotxTBbsfgKIlgc2jVzoE6NtlunJqArYK6v6cBvOt6d+PpbD3naG5F8ypd
mEwP2C4xAJTLNilLbnqDk3WfOD3zJ2t24OpeApGa5GbgWBEpPOePmiKyNnY/IHzP
BhR1a9GC+2AqLwSmpmtK8xf2I5I92AhkDy2enlYgI8ZKJ5K9dBZi0SMcv9tAMqvh
t398do4w/2cSFGgOKENcxq48YVJ75QI/xdBB991RS/G034K4IXo8qvlI4DQRHD0b
0P85a+KX09y7p5/4BxAA5YMTdC3fUHvkwu6Gm/NyzvFm1BbAVn4C7lWkO0iYaGMX
VSOOPshCK/N32YTG5ehG0vmP7Qnw0VjIEKiYuVQZPsKrvbpANEPO3ZmETawlWu+s
yVazrqoNf9oKV40V/zl+Fqoc29YTHvdbkA/iRIllhIiBR+2ZYOXXY+C6DRQbEWvo
u7me+LxzDi+05p14hbyNyXRicjjr665Oz57a9fGr8l7Nqw+NGNepGTsUOoKbrdZU
nXPKoVfBBkFNxGTlE1Ab//Sql7/c9yMK27up4IPsdtRmIkLEvpdumBu61XgDjUDX
kMUboOKFT4kvDeimPKEjPwGEPqzOhnR5mKktKgWIXuQ1MI6kV5SbLLFb/iNC+sTH
VfVSuUVqWXvYiIdhLkNNM1dNm1pmDSKJTZD4wJDbAKHg/Adin4NBzCntZBznMFaj
4sHkPJtNap66q8rsubjPRd9WR60DY7rOwAbhq6JGLo4vAaENYvdxd690pqcR6xtd
IMH3i37GMPaGIDvuXZV0MFwglqc1HyhK+Lsk8mGiONUTByP/QGoLdUhzVVpOzLjL
RV5m464pE2ruUVavRpwO8XyXUmKRscB+nHimaVE/jUv4VvuxOysUYjhN22Ayc41n
xGY+z7xBpkrlxr/4JdIe1TWey7Q4qPNudKohpXF8FzaR2+2sITucf1Ux4RyR8uIX
/afyoRecNOLHE+WBfHE+QGcgLCWlvKo437gn2WHt+GXbNRMDsXV0Lilr96MnmIkt
b9PuwHReiJS5mgs4eDbobydBzRSqp3UuCnvPdmp9Sw/Di0FO0VkCNiQGoBf6ezrt
6uFEpV6747DBwkONWgzSFrJDb8KLvVcGjalASXa6iWGhrauTRKhJK0lyHUJ1LLyV
FrFiMTTwCOZyXgMgLIzjDBpSwpyKo/4Vyn+TvfK5C983ayHbcLHLHaR6YqPpST/K
Je14ZUGAC2lzOkgQCfgTY/IoOgquQsV1gorp9VTMdOYDIthL0FxNera2QKobjQlG
mxN3S9+F1peGswSkD/WyzBbJSwaPYOL2Ps7YXdq6ETMWYwwKMm7FhSyA7gCFxvt1
qoVt7O9r/G4ekIMHibo1aMIbXyooWewjlYFW+gQB6J+tUXROT7tN5qWhdzYbSDIO
iD6chd959dFsRf0kmD4YX02Y0saIFgNxsSWMqXLfbm8KRlGb6jcJeazmeS93YmLH
qWVsV3jUWAV9P3WIFBqVrm7EIyFv9CbkXJxtqkHIS+PH98hHsr8E0qquE+JSoe/q
jDRuRH5yEWVXNKMVEVTYFZCr6No/0j4DvfgfweRANGy3hUnPD7QNjVUz8sm7jFMg
TY6LcA+UgydaCUAd4zZZcDiQYZN7dmwUqDUCMqdnDvsWb00wKc2rQ+QGe0acHw1N
OtM6ivsvh4azutA7NjVjfsGsCW2PSEr77DOxUs6rn+xQ30tKjjLGibTAQrqwXV2s
jDXEx5ZupCL0Plcl04jJPh+e4l2LFqQ9ry77STo7Ez2U8v2f/b6e8HR5MgBlZXoU
SCGJ+tsOJVKb2xDFTUy8EWtpiAnQceEHSMrwwX+XE/SH0YeliO8ndgh9RZo3etaZ
+KpQEXyyOlt+K2g89yYi+4Wom8cYgGZofZwk9rYb/R+apFmMyF+Jwub99bXj4hgq
il/J2i24teuJCiYLp3eHJZ7kikRGx5HEk/7Ak1CjxlD0RRUxXiUVhG/X40MBobG6
iRfU1ZEYI29QFCkub4tXeAo0tWrBgmIPoEFQ5SvXS7LrdkKdQNRiYc10wWZxCpy2
o4M3iTfTrFWuNYqPGLQnMhSWsxLIjCuevvDlBFkrsYb0oR6thZCaXY8UtEbB0ZVC
RaHT9lQmhJ7bNnNS3/iHxMP9d34Qfm4ed3KyZY+2N7R7tVi5NKbpLjKEFUMQ5ugs
jjjVun54kaQKn0pDb6mg1zP/RxIrn3dm04OmqC6gYbVQCvgu1PzVGolpwnX61Ebm
eL9JQlcRRuru4owVUsh6ORrKe8ZDyWeQ9edDQuyMMEx4WvcTwKdImb0bQvc0DwaK
O177ERdnh7kC/Zv+sfbialvBG9rS+Z0iQrMkndYQRfUyexAhc/KVN949ppkPPjS4
iMTgScv8SPk+0VlDiFlsTgUA2Uz5cfyFXI2ETWDUVEtTolDjQVlPiSvHee8SuTJk
tEZIiAEV2UBl8zEz3mhPtdSqMmO+1kJoGgmwEhW1sL0eY61QWGES+1p6y4ieQ5BX
sWG0YkMWW7oolhC/VTy3RXXu2H1IK60k8mfoXtTbQrmFUEt+zLZnGIVIIdWTf7/2
wk9V0FsqDVSX5TJQC5WsYYerwPT+gXbjxjUxM2sV/wuSwzuV5yM7akY/2AEgInmw
DsoBqz1OG+GCg8ORSpikooVlAbVXnNUroMxYuF/+l03mY0wnszwAxLozeQVF9Zrd
4Z8Z/ekmVABjCRRtf/IFD2geTUAFHvBzEffVesmxgoFyh7amS6Iq2yPyvGI1sTcZ
YQuAmCArA3i0BrD0xt2c2msejFdE00HGKqeZc4WxBt51ddsGPox252nazLqcI+hJ
H+8VPvBkTfuCUYKx2K6Kj9If9ihic3DcaYDKMkDLPPl/e4IG6iKCwmXyqr2hg+kq
2ncP8p9SohCChLtp6pg9PFXvXDEyG8jL2t84mgn8RvDdSef14QEQnKfqKYLoD+Ot
+8Rudb7lzG46B6sSmkDkjQLUlowD/p8AxUFjrKLJdal5Dth9vypva2Q2Rrr1ltMa
JhjucPosgOVxYvEGFLdgqceD4faHJoqfd3uwv6VayB7DpnPJuBvrBVfVjGrQkIpb
Vk3gSfNW8mXUV4i7hv/9N7RLJ0Q3rxnoahi8hKvOnFJcoF0aU415XMVuJDrouPSX
OGiz45RFrFYHicnGzH3u8yggz2PW6W+2AkcM8XO7OVW90MvUKx1FIqp86zykfAyc
md6dtb74NWH/0o/J/V/OffvqZYHmJFDxYW/MGS0saoUE2E2eugRfw98mBDPyVTRI
KhJi5js1p2MaoyGG9XFY1NYGBYDUK93CD+94iVI/BYB1VqA0U1Zf8d+JOq7E8mYH
PBOZDleLPtBwh9i85lbhEUeFjzP5Nw4LAZw/hDBCbOEfqY7gUoT3J+aG25qV2LJn
bMNd+mpdEkOnbMsEtj04TK3x3Cib2R26/E5yJx+AFU8FHojhD90Vx+mAmI9rxi3A
ma93BevTsKyBiBaJNGM0oZNNBGpjCF2Yy7PgAbgoiXXYiKhh07CYCuFTEgkymvvC
4gLdFP0Aafs9He7MtRzngn7o5VyLcfnwg9MUrGGXNYdoemFqKt7ZBQDxvCoLKo9M
LSId1xH6W5UNwGjvgVhjB3rEJWffo2lfNIALPej2Epl59Z9nzbJMe9DIVPzyoFD7
AmeVyCgue/4lIFp96zl7r7JMFAqpm+jHvhCsvi0ssRiCsAuMRN6PnlR32C+CH1V6
bj2gIVedgUdtFbAWWgUXPZkAQ5pEKZhHRnZKGMcGv1aAod36LUkouHrFp7I4ScuN
LrkJq89G1GIJuTa1UrEcAnvHTnez7Nh+uIu1iqjGgj6YHNM0PAt4QzrXXT58x7Ju
sh12pMsUUDFyMB3m720spabGcufhGwCWClHc1S2ZNrOPYQHT3Tz20izDzJR9Sapz
L1IHSnK372UnIxQXs5/QR5Emu3fht6pp7spMqErV5CQbt6OBse+/TMFMVncNa/ZP
WJt1ZfzzeLx1ANR8klH2HPk9LYvXcA1p8D3xF6mZTHmgolTzxEnuiMtI+Ty3252u
7idNjNcxkgPbGF+5DYMSscbDchPtV//PbD2JHdJMWZCKlpH2crQtBfON5Tkxehyi
znh/yCzXjGrNPHB6LyuZPe3eF3I+nr6SKsGqv/mFq8TMZerqJu1OHlwdOawVFe2w
VkpMHQLvOjZJ2rs09G5jm3GPCSYViPi6TrXdM1YfKXI5jZPHtxWRiizcswm6OvK6
b/w0dYPpqI22UkyTAhkkmA3UbgcOMvdS+/JTEAeElGmV9+w70klGexa8FSMp0krl
8lRu7/l/3NL46IxvJ2zSb8xOiNpqtwA5LGPx7UUbp7ON49gTVQ0ggYHebQi5lQQi
Cf9jsSI045oHWpA4ZZPn3Pf6PhlXSNSsWNcfA6l8cZmQq9EWHae728tG0w+ATiyk
Yk3Nb+RGOfk6ThFmn8WVBJvzOpe6O79nQJo5nxsUz2yI4KSmzMEBUda1A3Po2tej
Ta2JmEShLWldnuIsSduVmURKmTz5IMmJ29oA/7zfIu3l21Qe/Vr4UJWsi6PLhmMc
XCr4yBMcxqzFQrS42dNiInzAa3QgAjirSHQnAlKe8FrPq0/50yonM+6uRUfuiyG7
4Gv4E7XfVpxfoouUQp53pX9fy4CaC2otgAAV9F79+yyIcPqKuwSuKk2ZDuRLoAwB
wHNQGT1tjsnN/YruIGHgima2BzTZ9F013IyI02O0gLfh9yLpeKD5F6z1J9o9TLAf
14tDA/aO2QaskjF5pHxNPHx54ixrpp7aFYYqPqhjWmQ7OSM7PszWLgWOeHixDU81
Xlp6DPLK7je8/5deCyO2vahtyGXjl280aWbtjqXxS+4jHBz5lqrGeR5SOImR/VkP
uTHoQzeGJIRQ4hMsRa9jd5Vtzz6DyKnQACxpUK6TYUOcYis5l9z37g3nCpxrAesA
u3zFzl7y2vo/k/11f0EJUPif0UKs2SM3yIJ39SE0s9lwmFd/imMApanK1yuNOVrg
LN0y302oAjUgCRrVDb4ou3J7BywtmQuSWX4kkcmzTkR9V1cUeMIUl28r87OsscbC
xrprVD4EqFzPe7qSLGpPfSGx+y/n8UkIdjseVNPqeIx1RdlwgltBMoVqYfEhUj+S
xI+6ScmuLfolNc+E5YKaoQ2ZV/yPgTVTM0VLqfDCzX4yY9EPhimhv401/d+y6w3H
me3eKfpXH0hfVMynaYvR8wFWpi5pntDO/B44xq8dfssQ5poJnEqDwgb5Cykqu7YS
ncys8hLC3nAnVYQjDaXGVbDy9becf5hFze1EuOr+KOuw4CauA1wVMzo6Lqq+iczL
9XNcKEe3KK2geLLXKXY317hbTSzKtAKY35naLbC69VXcSo1Jgks/Iu8dmWwJ9wYU
beo2G26JgVde9fJtrBYjVCfTihxZhHqCQwwOqfufrWUzEG8YoEF9Fm4P3QQ4fJJh
2zPa97AkZr+HW5BedEGNg3u6zTL9PR7pDVWbRK3mvA2dEwV9vUZY7vOT20L+m0vs
meV4CSkxhgv1OkINODei8H3mRcZyc2rEp1KWIUNvC984Ut/eL/NK0Wv/Xnr7cfR5
ikN8Xedpyw63b69a0+RxwseeFlA40gBxrl9MzbcFFiJp+IBEiAzWB/xa54PZt22e
+uQqJW0TShtLm7ZU1n+og1mXuVnPM3cl2F9WDkzAImhfHTc12uKwbHWtZFfsYIDM
53qhTaonL1gvgY5dKWK3wriKg1ZmhscoAgbcDy3KNbptqZqo+BDqlksjU/YwQcSO
k/Sx/t+vfWZHWyEhUNDqVwVziMo4C0ASyejQ9ufcoKnX8q+DJr9IiNcxpnmu4LXr
xFs93u5ISwrqtC3L3xmwi4lhiiortJjEhLLLTerd6op8ShHd+BU7xSyGgOgDRjpm
eEHLMvjnu4GpnrB4rVMzQwjtygIXdQypVVW38KIPijf+dZ4Hy0CEko+dRO8mXuBd
78YF6b1Ib7+RuZF/eJWPM0E4sxSqK54VEtq3H+AaDNzSTOBOQ8jLYGjbUzfS0TCX
dT12oAws6kk+QU0ff+3fAaZmfErD2HjCr3PNj1GFmvrXv8K+x52L1T/81u5+N6te
6qdOQbV2cfYK/coUIAY/uoKv9D3iGmwbcK+X54QcYGhYlNTXB4Gl/KyWaetfg8OS
t6cGIVE8/y/nksg5mbHRgSjdmrVzdm2kttzzTzdxvGVBJpAdL63ktH9TQuMUkZ6i
/ATSxzFgSNYzLbPpP5yVJqTx08OqIHz7X57izmdXYu+EC3g1/iPMD0xQgGQPpoSZ
Kgxs/ZSBRcPItcrRhcbehv2KjHXLT9lJSWQQcEHqRVkNTcV6/xb83/gaeK3W/QJg
uaG/oO856yPjdnkhUejntRqjptveTbdiO7o6cHsdJnHfVm6XM+QIY6p4wOi+S0bV
5XwB/XuQ8wPMNK2FvfywxWPx1uFjRx0Pjk6sngn5W9vHh/NSLMHC/XOHhIC+D7xs
QhBaMqR2S7XzD/7YrIAcHxuVS40HLF92yog9Aaqz3h+Az1T38Qg9jRaGsCSABIRQ
ZEZiGJJz3180Rg9UhVjPlPNBQCHvpl/6YVF/ax+7do2z8tHHhSSw6vdqwyAykQQZ
cUKiiQ1DTnsO9xekKkKDbWx/MiGVXJveCDCHjqVjWbXQ0tHJ0lQJ90/FkhVr+sjv
TML1muIrx8GO8CWFJj4X/aQ8YAvEQfRyMwTaTuftYnvKyiLwPAIgM2UddksJNMJc
X5rf+6NXYDhDiVUg5Gy+BL5RJuaZE2SoE9P/C65c8qSVxasczDES2+7ydu3R8R36
CUIvbXa2orKV1ynhFf8+GAwP6c6DSPUf1RTYsB16PigpoaWfhrNM+Lks/X+NR3JZ
sHu+7r5m9Nfi01Na7JNMMnqsA8CtOUX2tB6ItqLKiW4gBfzXNjty+J44DBJQ0gFe
fK+Lq8/7TRLRxS4Gy3UnfErQvxcc6XI5gz6iLYcROVf4GmwXn2YCqI4SLNRfWfrU
z2mzQIuw2ZLoqBh05vFlcPuDWVYcE/IVgQc1Vo4JgKMLNEsKmrPDcVqLX4adDm8g
Llz7HbtNG2j/gECn7roa27R5J4Mho2efdHecehgFeDkaMaHH/NQqp9rWmXtC5wQC
jgENC1WzxDXJIRHWuX9Ay1IM+TpCXSY3cwAyBwqjf/cJNDp4PiVD6MTyD+RaXVc5
jdWl8jhGhvHphk27WxIAwnP7hBjZOXY4Bj/LqsEQeuMpFrEIGCWjfgH9YXQr4FPx
DuaIpfvkQkvzlkBeIHm6qlaCVIW187yi2wTR2iMwY4Ud/9SJu9GKPKSu0VPgDAP0
q2Z9ljL3GhftHjMdbyMeWyubgODC58kW+wtSeZ0SXCpmfSy9tMrilcAqEIB+sHw7
2x5sbWoHVGJaq1adw3GD5o2cWZudjfOXKf5P6Xbvi/g9fTLETp4surwYPGJZiLxJ
QwtMJHhUUw1BZbV7Y37GGKzi/GvfB+HnFdUvP1HeVAFhq97Hb9YRjfreyqXvrfI3
JzrZkpUJa+JlD3v9xAxkZJgdzGjrcvm07to3n/9eLyZUsziHml9ngdA8i9QsezYe
ZWisQnNF7Htxv0VQmdABABsedR3fNtFJ1EVpTc1GmwXYI7lLJRlqtVk85msMTsoO
ZOIh1hzt1FbgKMjfJEpzrrD533Y4NNz4HYOOZAkzU5wIDTgByZQ6XWYvVEFY31EJ
V9ke/Jvh6fzu3nzls1epXgUCbiG6acj+AtKQaYEjZaFX9QwzAJXFhwwUkWMIvsqw
UwdzAu1kl0UGMlF5NV3PuaIFZ75tXy40CV8+CfZRCzg8t/4IfghnQulXYxNnfBcD
3kvmVVfLxGxZtoNmWBreBLEHtq2LPcTxLLrInHguHyoXr9DdNnItYZ8iaDF3l28S
4BTExzJpuZveZglA+MESCp/PC4wy4V8S5jFCaodc/WAZG+WQJDhWUtFE7jmhDcmE
3wRLL6zGrqYwFVd2aXB44PIxJ0trtVYFBGOzY65ndkNzQTyVao5rKjN7c9s4UBTC
rxxPbo1i7Ov5uUwIpkNVFB3dEm5P3pAQSu1n+Go9nt7XWA0PRvTcc5pL1h+bJl52
rdpzALIVU7CyQEZTnWTEd1Mu88g4YZQOvVI/ozwcoSuFHR6ujqxDBPw3RIQJj9yF
HPsElo7W+nu4Jfmveih1R3qaKX7MkhWVUvjp3qZcHV5HxokK1kJuSniyaErHCw8C
oVXgLz9c7Fy7Oo3hIC2GbGC8HvYWm/AIeRKw9GG8al8Xudi27l29KhwZnncLPOlp
fXVkw/7/5c9koB1L5O50pP4pYOq0tXO8P0+mWmTDPCjOKoX+GJ/i2zCyC4sRnYcy
Y2fbcbfpUqRxv9wmKiAfZ63QgFUkpczak3avpuVE+vzOzr5uZEJjo40K+4Whd1gM
TmRMpGDiGPmragyxWAQhjmRRrNcBx3O4DrKDLv3Dvtb7V9+iPNnPf6DrsmPjNVaI
tCTj+Umv08u3gQ8D8JFCLvqJ0EckZGPqopl+SrsJo5/fmdXkEJjRqBUWkZp1yJLS
Lz/t7uKIng640eV1nyDu+C6RhecGby17SX6Vh0VWOmMSrjpEhbG1zUcEQpUu1ieD
vRZSs+EUxR7zPt6gJikoZ+7qUYJmhK13UCovPI1yNQHHEIj2ou3kwvx+qDdRxoHx
g9qzt/In1lzbQu+7NWYR8nDzBvhtGQThmWderh28AvpIH5/rbt4YALeSgCr3eHuQ
e2W8iM6il/0ChSAkd/wehp/Uc8II902YDAU8Fp4wRSB9nwU8iiEaxodYXVnBfUa4
MlWVUuFlOUMFnvXaLsAOsrKgq2Y7q8YO595CDAJfhbPiI9us3DHMrrwJT9ckKe2E
PudNY2TVf/wzSgFzwVCHc9GaSX+X7gefeiKQmPK0iRDwSOIGqdZ7zRqzRYYajyT6
IiV+wpcGtT6eN5fF4SNBK9ifHr2crImBOqgIpno23SuziiNWhry+0WHW+iI1rXv3
u92xk41PwC2xwusGeDDIlm68IFOhFE3dqg/RefABqdrGB3qGUDj+VhMBGCrGhT6t
8FaXdilxvUA9rPB0mjMABndikE3eeHka+g54S99S4jAx1VFu59O2hfLMxd0QakuS
LFcvpUVTwNQmxLZMni4eRxkZyxBTmdN7UvSmCxXIkF0SHllz53grmuJaFphzBNVM
ZuS9zMhUFQcxYH4cvXfixD99v4JvCtvMbrnxyfjeg27wjYiiUREtJ3bEPoiZnO9T
q06o8X+jEEJ3Ry2HTvqsvSHMU7/XPZ7jIbPFv3zATvodQEst1HVrEYOe8mfgx1py
W2+Ni1QAc4X1ekbK2eLrMNJbPYOl1I4NbJbgW62iCSSlvmIeEqiyMJ82mAiTyF67
I11kFI6NEBK6kZ5HRQ9PD1QErPU0CmNZ1r/rGiGgwPKkVZwDCnDL4khEUuOL4D9V
isDp30SAOa7K9UO+hi53DO3B/1KLo+0cek0LQzBD0Nb2AN/kJu+E1aSHvyHXdIDM
6vJj/fOKEQlSjFtoU2nfMhLdRKFSsQfXs6AsPOl73KfQ6ycVl4xaZ6PDVUaVe0h9
JK4oTiU1GAn9xd/mOA2/hpoCKLj1wDw5OYQSBkWzwgMsp6YkjM9HsZV+UQOCDO27
VBMvltAmuTi8qVvM8kHXZ38WDiP1eLJthIFx9U6Vk6RASxTObAsQUmCMXLuIrgFV
9j2aXT6fOo1ag+TEFcTh+cvYV8LMG3amayuBDaIoZlxOgIde/JYa7WB4b57ZJs3T
SD2j9J/NunFjDUFSkQWUG6DKGsN/d1yfwukzs2oYc64zCbv+2K8IZFId0sCQB0U8
PFwQ7F0J4KDHpiqtOj7aEV83+PGGAtUI0ggELtTLEGGuQ61fWRO7vZShGG1jKVci
phY56tUIAKnPssnrmXPVF9luKq4eQtcW/V/SntTYVPturqloAAMBZkH53Rq7l2Rt
rNOkptluQJ9DBAQROGcZiQNlVsvROrD7Qmr13E3X6Y/YMJMVaFCWVWrF9HsD8cRu
ZLPdklV56vck0IK3wMx5QhZzcLsCCeofyeZcyjmFAX6IuGTjhng8hGp7I4qjMGIX
vYTa8jvVNhgaJUl6VFmasTTuIEd5rk3urggkg9LUwonk9UWFLyFeukkGB0MFjduV
Ay1esdRq9uZqJx8yhobpVwrBaxBx8Wvr/sVzRodVG3DGkOXcRPAAMVZ9sEjJ+lpS
vZCrIsSpaQyr+63CIeyTU3/jN3WemHHRpaW5VuQrWj+7dmw7fSvO8iyPgQYEtdyk
7vbHZVAOnjVqmG+/zZdgDla2Wf2LLHje/KyeQCVc2gfHrrzRBbCi04y73ZBzdA8P
8ZFhP9Wwh9p/yeI7wTgdNbJ2nKlFa4Y6gp+Z+Q1/U8lfIPaP42Z/9hFZSgvbTvR4
Y9d/zqcj98+XmuRTszv4YO+V40fyvl2bLTVx5ggkMxQUnvlklnv6sAPj3l9scrZ/
u08wPH9LEg7J2T3K0IBVD40NF1O1mBO13V2HaywLB2RmpjYEa1v+qEO6QM8lw9QI
4pyFH9Ig/zEMWVM7YN1EMegzcoTd5E2lC10vaRCbc933SRc4Wpk21XENUwZMjy6B
lsoEFs3gzvdetsURF3MA7qVMbhS1uFvo3YPxFR+iS2lV6Am26hxHSgN5TNkDVWOD
RoQjFOKqgF/NNF1LvWEIjsuPG32OJOkoC2p3E/qqBkva1IM3zpZvuT6atY9V4JYC
mt/E45vnQPbj8YLt710akKqbism9/PmXuJCnaMatFeAN/D7LJNtbII0xSC9TzEtW
j0PMueTgXtdtoW3VBE2WCdFHHpDIDRTfGv3xISHqqpwtuj80IeYzE4j8qKmXOJpb
1xBUIO329xYNrcHg4Cn6TQbECOBa8aINp30vJuwiPi7LiwEjr72G2IiK3bgZGzAH
1y6JQoQotdTtfvsci/rFaY7RwK/cfobJAThdT3mHKhFGXuqgHoqBU66XMLY88mpU
2Dj/Ar4f5PO/qU4+x8zrVsXe1ZypBR/wBYqdmhuBH/7rTQOGMjSQRuUSp5xIvDhQ
9Az5MmTdwELEecLYE+hVKuklsGXaxRq93gvbf9dKIPz28nAs2AgiNhgIOcmUZSAl
5ff7Xf+EkGJg0OhFxbfKAmjEp7MFk9cCMXOF8/mnMbV/TP/okNNDkNVFxNegTklb
OM2U0rGxLCRDkdIXjNGafEiv1lv6r0ZvYd1Xq+uOXY187PRHKwToF3o23GVRB6ZX
B/5Y8U4d7oGbppgS1eHhD5syP8YoI84+QANySYERSyOPQ9nlBz1anghfmeTfZGfr
aigpaKLarF/E6N0pDID0QegNGYcRjJvJ22z5HD7LUr3b0mEYt3SftNuBBVbG/Qt7
YJbZY5A8I88IGEIhdll3ef93jcv7eip8r7ZcGH5oeGMY/mcNJQE4kUtXeGcG2jeS
qxwYVjfuL5hogBX8NDA8dlvBfQbNhK9nlsyPUqTdbbfWxepnzzGbz7O8c40YCoOV
oA0J22dtFVGJF90o6mH7lRxDOB/CKL4Hm0IpDXSd+GA7/XW8FJ2BUcxq2pxEwKh3
lV3QxHSPqaLbQFmDrDW0nomkuTUp8eeq5VNeYPxp4fS0uJUXHwKzI+khdL6+aB+x
MesRQcz9dEezzya8Ae6XCHxfSU0/LPmGfkoqwiHSh83lo3DSV6/WeHP4MUdDdXtZ
lsQcx3obKG4zsPE8x5OByrnaByG3khsOo+60bKxntTZRaAsR74Ri8WHJAZs27z4h
8NmRzPHqmLYrFJ/cexnHWOZQIHIqC2O1471AL1NfqSUtzKcr7oVuK45qKj3mjrll
uCJ6kCseGeNROEihRi/OmbELACqHzucHEmjFubnOQZh0KvS0p3EMwy1c4siXs/bP
aCL0LohlQbIWvmOFHKq0Y+BOCbujKtQg68zf9BR92AIs7eAEPuIth2YHkRyoipLM
q9NrQe1/Qz2omSjs/M7G3T7YyYj/R3lyno5nW9X0CgAmu31KN+oySBJX/MLAu8/8
lECyIsa7b1It2JAs2mgwsmiUqn8IOdVrQLYgPQzszF5RInnzYkvSKmk0raguRa8J
ul92dDk7z6wd4XJ53ouQJD5dxHqiSovyKIkm5cpWmio5bwoyF3x8OSKgPaBKwjFh
wVXHMnF8Cykbo27FxUB2FokdVxhBlB8zAp6Fe6Bi1NtENk9+cMoKNkDABxbta2lO
BCqMzI1YV8+FOPDYyUKyJOXj744aTjA6oZlWbdO3bLsXHvKimwB9AIElcO1e7Fso
QD8ENBA6X5O5rEdMEWSyM2lY7odX/W5Y4345V7OOLHzWkW0JZ8Y5qJnOikYC+RY2
DAADmvFMASQbF6gLZLxXgDIs4iojdNi5GrxUyUzuZg5Zb5/lA9fA06H0SHpwY4a5
pkwmKp3WR9vxeJx/ZX/FHIIu6xIKDU7vGk7VQMHLLSaIiCqnUICAmWkyogG+GK9F
hScR186JmZfzmwc9OCVUFkMRBTM1/3PFaXZ0Yv35IMuimWH2Rw8+qXh8KwufyhP9
H7t511QjYyLMxVvfQFgUtyZPzwJwvVtj6pTnSKsIP5gD6kcti6Lw7Pulyk2G7JFB
gepAs3eJTIdlciW+8RL7IYV7j1WhC+ZOcVHTyJcda28SRMb4O8XCmHOk6OyZr1PU
m496T8lKLHaf4tcofWIi20rsiyrXEz5FqJsmDAVleUjIAvsvEbNl2BQV1ZYWNrFf
SctXZUneMocJ5v15MDXXUCLFm4q2VtnPox/+Zgml+LXfCWUP1yeceY8G4C4bxVqF
0fV9aPQDbQsCMdJ+McVZYlfOhhsbtJu4H6irH6rVV7MJY6R7vFkEc3yUBaNrQBZI
vxEpjhlyANYl54M8XwVnBsLzXZEaqlvNWVqS9/njpIeEnPO1w7nwQugQ567kG78I
IV8pYDuNtj8y25xFcdro7QeczNEFcOpXe1qHZmLj2MF+4EXpV9JLMTTEchy+/Htg
dLQBSlbBk+lFsHjNrARkuN2dx/+94dJuEonHCQIPvUGEwQW52G0UQYgXsiwWMqcP
Yim45rO4UlenWscTo/gC/3o50c/gpOG6zV+qWI2Kgr9671gs3Zs7RSyp2xWPI914
9osOVrhcp9P3OCQa15WiMk1JNFhACIGfzGBbmncksmUMEv+49nOy1wc7oKboulFe
SZQBT+Nc+oCKCC4c1ziXD1icj2UHgytw9NGz4nmlvwLz6uAYPrq0K8wJy3hIfQu8
eKjxZoLUR4EM1BlIK8ux0tSJWFVNpeF6MrQDN07H6ZfEpq7NBT+OOl0ta+x2iR4a
5jEyWjGdB4zaMx0Y8YsC9itvcV39VMU6WwgiZ30iK+PVpDQBnGL/LuvAJrx9HfjZ
qKN6hMXy0QvuI4J7n0F458GvZvPTukHlmuJjLo4rP+SkYNurW6Rqt6nVUnKx8i8f
TXbG+9m8gfedtF0uKBlNq2NuWVbG50HogrS3QmMtCqfRUidj8UIW8QHTUSqqlCr7
AzBqXP8bExwgAUzd46ggHgSkeFixlvdELLhaC3xpy8HsG5X0V1I8yjWueQYooRFX
YIvlqpTeUqcwwYOYWGunAjPNrXkkrETaJMDnlvUub6y0kTdOr9aZ7ZnKptYuhnIk
oJf7GgVMcZNVgfBn9vfXJbra5OIFiULFcHn2MZDn9UMT1XBnEDS1fGbDRCgiyH9n
72bjDYBc5vgJ8n//AqQ2lNz2RoJkotrw20An0mgg0nVWl2KJoVxY5dR0j5O3qMzD
sEVtWsPOzuaUOtWlUBecCUB8BLtHx+8DgE/vHVy0Uhv6DVW087ToFe1/k8g+DeTs
tybKHJj/ur877vHm+rm9C4LTjGRpXSaFdOE8yYyLgoxzT5nVA5+Awjl7tSFmgnvd
omyEDykj2NmVYlQIMxFzehY89YfZoSdWwVbH3N8A0ZnxjYp5QcAWFYG5FfzMYjwM
llwE7mHkvK4sfHPWfLMP+Uz8pMaB3qlGfyUi8isR1gpJIQfI7NQS1Frq0l6HWriP
9BIuW1WzW5NEPvwx/TnKpY2MU82tmy2X6fF4Tvq4Y4WjOkwwzp66pHyxUfTMzINi
XpLmWe34bgUvZFDetGPgw3bswdvq+Bv3ULGxRduEecTa/F93MybRMVwSKpkjyEfm
rTyZL0j60W3SCmkLwQw0YiMzHAgbDwaXBF9y8Jxw6MZLcj3nBRWCptq45z7cLM8A
oQOPAFORnEatPv5hlyG7XpwDUYcpgyzGETLSYnDvgn48cR/duofvGvDzKRTPFk15
5/nVGuo5Wuf2O5Bfttmv/VKx8IoYCOYslfKXutytr7Mmt7Lq41RLi/6KIg1aVpru
nRuiKTztZ9Nqovb0fNc+rq0pb8XlgnjDeuD1EQdX6RvMDk47UoMTo6Zo86JKhdIm
k7f8h7WbcSO2A/ktVB2pQhRqNl0IBP4I+erraOU1hxefQ8kHxzRJ4Xhteg1qozrI
uLuJ0HExsIeNw2dvOZhD0s5+DH9d0e5Y2ZvQy8cc0rFfKv7FH7XrPCDRtxzac6dl
30z+9IXVVVaN3Q8X/OOwaOUyBB8UYnxSsI001pab2avlBTsl1s/ePLSFNi/wVOTq
pdkP6KLuiczD0NvbAD/KtkpQnfjYaectukHdf93DEYfc+2hlqcarbZ9j9Lm0RsKO
D9s4aynXKlOiIkhumPGEe/ji+7+v0dcugC1o6TXS7MvrgK8kOD4xzxyElgvOJ/k0
OaZcbJ1JS4jyrJ6zmIHeJPGNa9zuYrtJpRiv3XxDFsU10BvHcl9Jqg4RPUREeiGf
GwiFSkcXFMhER3sABgsb6ui1IQcljZ/ur+gqYlBiE09tFuA7dy5gUHoXzS6x7A0C
m0QNJdiQhFnv6FZLL6AZelyGBxVwW19cmN8MoAa9ryjZ5fzox8VctdLAgTcVYC/D
lpXKkdKKfVYu4zBdDykjfeyK0NMOPbIx8ZwCEhwXZPfJ39adA5YAQHdQu7459N20
7EKk9v3VTQsRGJ0P4NvEa5C4o6Sm4qcFqhYeCdEed47qMX015CPB2rmMt88e/Tg9
4650xh601ZZK570vMCvO1X0ypJ3bJR5jp89+PWAs6cJSSEfIqRhaKV9TKSgNIYqt
8fYTuHmaCXnx0ZTtllUPlXrhRHDK96nPwOFyhz3/+k6oR3nIi8z+jilvSPY39XQ0
hZMAxnNZEbscywpBJRcf4wH3iCwCzmmZb3Iz7LFZmIU5KuGysmo3NH6KQfHmfnjE
uBTppvDqns3NVaJU2tTXSbc7/u80BESo0LkY7OM0vS4QE1E2Q8w5iSiIy/QsaO41
+2sretBPY3nFSSE04sPgwSc9IDynDxjCzOvqRecy+YjEhhCYx52BVgjCKaC8EXYP
QPL+t1MgVDZAoU/CytNS38eVsvkt5UjeK/tpXa/DHZAuqzQr3SdALm7GW4+X3BYZ
b1we+N0QAProXFJDZiHyzA9Vo3zo5sLsEbqrxGgILQ71p9TxqeoHM3MisMzRPNbV
+F8HxsPnXRpE31rswdIoTxUlg+QrDfG28ZrSXuvjeIKzRdwvUJTcEeAms0Cal35O
S5lpi0e3QNrqLLZ8//Y8ycfx+mJ1dGhJNTIMo3pTWtEy2luuK1eAiRZUUvzbbu/d
Co8SwEz8o5yLPyYf0o9VEn1Fs08HjRPpaX3AlAAwnYcHfSlrZHfRr0wz67CgMTf5
29NrM0I85DqK6Gy2s/tfgzBPHgbxgeNafVXnQJZz1VdWGKYrzlT0EyT8ODk3ZhL/
pfzUsmsQhlXD7Ro5AP8WDZRwDqHB7V3FquhYkWrPtX/FD2mmbk3xYQYf5aS5uYdd
aCL3p54PC4HOwZxkxsEPi94eIaIjWKmy0WzssCAZfWPNoVJ9WaQSghiHmKdjLzb0
BDD/+V55Kx9i3AYeVvRPnILOT+f3oOySeTnJq09CyZJGWfWaQgfqxTUtZVYz7iIk
8Cr7vg5KW+D0Xv4UChNoPg6zI1cHFd4aDMwr1SDFGuM3DxN6FWvImZ3esSl4Ilhq
csIELyltW555U47MqkcFQ8+qKsfYT+tTkAcHl5Zdu62c8ym2Ai9h7rk8vS5BVqdS
VUHoU3yPs9TjjfTvuELRO28bO2c/r67vUU9sDoZtXZgQju9cen3Xoxau8RY7ZaPQ
2lgfwcT9LGb5MIOu6mSw/9/F762W6fwpOfti2MsUOwKFtfemSHb8JkuTJ/WiBJ6f
c+aWSLEdsPZYmnnobsGa2E5wQT9Aj8bNRyLgmSiZeo2+phFMNeMlMFV53zSLnWXX
859npi888GeEr2CNfRgzplBT2R3IxPUbBmZnvnWN4LTOi27alZFiFpXanQfEVVMf
fP/cfCqfGEevZQ7Y6WvRwBtGDSv9nu3y6uRPuGJq87p9ds0zV5ehokoZPOk2q6h1
pUADalTRbEOYWFjhiv/K60R31MdCUPw4SA7VyxJA8wCWXQd2S6kz1eK5Qs8nUjZ6
kQH5QaAtR0kFM2Scwah1I47YIUBEAhz5q4vXs64y1XZZNiePnplwPFSF55yKGpeI
fvvDsz+/EEnWq9BqUEaFMrgNrsrsJTaEkGv0BRBCmbLD6fKZ6SBs4EyaMEUQVnzd
LlN2f5XYOve+T9mSLa/ZhRgYLO8GD2PH+8HQfc3zQDt5XN/bssS2KseDOJ26qxfG
8xhUrqMs5Q3w+HkEtxmn3yMtlqHU1bm7D4pkMrN67SN3zHW5+QXEo5UcfOC7dmKD
1giZxoA6pdvy+tl/7J6/SE1f4TD6yCeANMQPUL8mMylvKfml3GMzHul6/ecFb0mN
Fsod238tDN7uhTkdQczsWe86eq1Cg0XUPJolYi9ndh8CB71Bqe9UIeLOVqOppIJd
iWLmwOyWBpe5mitfGEIAPuSoXBsF6vePLSeqS8narqcJRss9m0o5PQMoVkjNWbe3
rJ0p8Mhd7TXemQ3y7uJyfl9LlzMjmolq7MX5LOQtDskeq1jF1zWUMNZuSgcUrTU9
p6zIdy3zgZ/2mXKbE7KJOfJJVcVYRIA5oX/OiOe+rgowAxArmyJ0le7D0la9/WTb
8dmm2bCj28fFdNsoMySnP6PWjlb+/wicnOr+QnsZn3AyFlDyGX9k5Q7Y7zJQ5MQ6
JFLDm7B0YVwq+gb94ZGePrvtksU8uytSbDaK6LxAD2is1Tzrww/G6an7gIKWZo4V
6ZTAOfD3J4Nj76+rWsrEGcQtGG5lzUvnfd7FU6FTfzMcZS0bQEO8frQ09Qkc4mDU
ZClO14FHIHO7H2EpVDXlcxFEOiv8NZw10E68CR40NFHB/TI0NSU+iiZ7BKwvYonE
xtWRCZGx6EcHMVUjhFc4md1XDmcOdoeOU0Wuqsc/lcdty6M0jiVlB77b8S02xXWo
ArimvQnXpfIsbHjsxAT47g5leS5Nz4vk6yBAGFxbi1sjqp4w4u52OjfxLjqcgj7v
3PPAsUnZRu3OmIoNKpeeyHlBMscWRphdYyewZOaBr5KOKV542sfayFTGsHnkOa9k
whNs2Y9pVZepgh6oIe/u31qSPByMs73/og5mf4xFy6g/SuZM1fyd3YgGxMGHjP2I
HXoUH3x2ZpatWcdiLCGStq2hqSLlFcWeC1BAIyg3ZLgsISWwohRYXtYRILUGE5tG
PkyUO2NcQzuUXoqAj6d6A4ZC8lomxg1bmdjafFB/PCdBUzw/ZzyltEn8twWpNfya
c1OkCxZc8x7oPXmG+OdVsLeAbPz5vETEeCmYfbTjKIhq5t6yai9IQtQgZuu9HG93
+cJoSyJ1WTFgdy3MjO9RF1h0/cG5iOJGqCeG2l449Q+WW0rAGwEEd3c5AZHdTZz+
Vo8aWP20OqPgFGbHiWyQEl3hi8AMuvwtNz3aBmoEq94T0MLP0pgcgNky2KCCnwRo
Ko6Av8IoIrT5pmZ32qpsoI5Wd0TkgcDrOHCwbrWhkyXX/V3dE+ctDz94ioHN97EZ
ETDdFgPKIikHq62P2VTwfd4tpM03Rw9OE3EzuF0jxTR2QQBALf+R8fEvCFwPu6aB
ALbHbz3H5PYi4kqmFVtchZPXJ86gT2zWEAnGWAG6BtrxeHPgRbY7ThauDslqso6a
+5UOqoLwAyMmi0DBL6sT8buWbTs8UzoOKYCOeNPfny/DKPImJVuvmjbb+Ft9t56u
aZypFpxOoMSXTt3j1dS8kTZ7CO3qXa7baNQpfxPpT47UTorCaUIpPGIHmyq/1cWT
lYE92n2ReYwP8Pzf+WKQA+YbcoXF4HAGhroNLZ8ThKets4lpLnSuylpN8GKCq1y1
5/sAa7t+hsF/JoakQFF1QoTXhH+eTj63fIZi5D6wbIQLWs4l9B6fabssjICVtfcI
IiQCWLl2CVilp5rqQFQXfUAx9thpcoUGKOcz+tmju5jFaAgyxwpWWZQnwUREMZ1S
L8aFiAsTRJqEox1q6vp0zVH4SkwssAuiONN8Ah0P9p6JfRl3qsRJhEYAEn/xIqII
Q5f4+K5ZBidjwUucWHJLGsF4T0Hi12ikg7eCkuViUPHZfy+sWLt/WHiCN+fS28TY
88prcBQWk+Jh2A6L8xdDlX800iVkj888B6HAGadbi3JvWOKAmFJTtpF0H/nka2wE
wJdk8Ro2KvAL+YIiDbFJw0nmUc6dH86IZ7tEZB73xoYJgtbtBeSQ3v06nVEgEQuU
lvSY5bMV96+dbfee4KP9dVDrwh7azj5s6VDRGxJfQR4OHCTg2c/GiwuW98nVLeIo
iDPRy2MbBJ/eBisNes9WsLBVYCFgVgFFTKn7OlRW/OrQVfQnQzQvpSNstBcR5L/D
9OOgXTvLfIVAF196to63A47TCtTBD2J8ZWlRAhLeIDWoq1HsEX2zYkEoGqOmQMDV
lBY4kTf3oPZG4hHU7t3I2wWVJUErQvwdM90f2TpWpC8LrZaHtQKwKhWpG2+Xg/BC
YIh5Ms0/7rh3q2wnyjZdyr6FN2TS8uuRL0opvwbx2WMt6M176/9L0YnTV1hWfFvo
5mYtrgNpHomkGlWBBjfp+Q5RQEevpCwo84QNBLxZ/r1VI5xQD0RyWSF57ogT4ihl
RLZOQURHLocIDWU14ZGrY1iRKhH17WyAS7gzSCjdU0vSWmwb0hrbwtxWgckRT9I/
6gphoLvLhupsxpdiYZOacOXfEfgrXhGx+O/83UULEYs0sGzoBnfyoXm7dzaX5hXf
0XBOuOn1umXOMQAHtvBw/fwkYmpjFrbKn+5kYR0DoeBk1zQI2CnSNvzMenda+jLE
lj7je99IBWUGAdyWq1vER3GMKFGzwB4d3h1e1gKDBXPwi76BX8A/bVUVbtwUPhTe
KU0+OanuEY2NJC8ExPysqR1l/eDvfQLq1HQxDW2ulWE+CSPfdEMg9983sCwXI6hI
dngG7mKKWRdHCHivfI/1BJDYs/DXHFeg1Yxbeu5CssGnSqeX6Na94iIr2Yn26Wr1
28DlR6oCXNGdK3vfPHrKAHgzhW8ZqvdH45BTqwh3xcbmmieW2Tl/mlnqiVZZ5nEu
iAluSMi5+Z/7zLjXa1+M/7zmH6GVsmoVOBPQB7iD92mjvjjMx79CK9tYL/n2QZWc
0jRkcmEF3NMvvmNymI4HKTbWX1XF+K1sGPUN+MY117ku0RGKO3TkI5bTGXyjt6Ch
WfiNLpD/ufVZwNTpJ3W2GQYyjUNpIMv6dconcN+pJ5k11WyvZ4fS0oEZ4UBWe0j4
BKXsjJeejnoAEOU/xP8YhVhCkYcd5dEsdvQKcZ7KCFsSeYb49DhN7payDdQalomH
cyFeQfyC16GCKmQhfW42HstPjIWMVIkgAixRohj9U9DpHY+u3v1OpgHAEC0IDB1a
zXB4DSQHJE4ME8f/xi95rjdAIyzjs6aMELlOZ2oljuYaefrtgpiOLHt/yVTE/ymh
Cfhj04dwJHu0KE6W/P08Q5C88gRX9Pr4cFtuhoJm9HdXHgktS5Fn9yzQqcc4OFY0
4vLhZop212TA8XPCjJ8yCO72ZQMQ7C0Q7n3qv0fvW3EDVKE3J4Jkk/kc083THAGG
6YjwyB5le+dSOYCjua/igGqP2HhJyC7n7UnoIS0yvIduvY1z7g8tZKD24MVlzeeh
vQLymgonyiBc82dX0cCacYjqkRLwm6QM9TG7NV+WKF4S+ztcqd3scuVKLDY/7T9C
b4ff9V5prEax7Q9egLblwI+WclJVlvx5u980urxcM1IFeWNezF9ZLhWWf0IT/XF/
GESQvvQ/tCFybzcVuX2Mie/mw1cu1eTVbNuxQLpqPQLDzZ/IZnQiPCl3vBwQDNd4
/KC1cRLcuScD3iQDjvR3+fsTUSMqwCpkcVyWPzfbY3TmqKEhZC5KTym+EKJ3UgTe
EdWiUhyg2Jk0/b+sqSttB4fP7xBtQa/AbWQnAo6viEw9wX9zWs9aXRVJ7kyI0beS
jITA3zTJvRs9b3cfJRCvSFeUGWWsCHK8qWeIrk9JPHDczGBVqRA7ep4oiXCZyDTC
IZtAaopRLVvghR4wiGXwTAb8Nk9A6u9eIzMpytO8Xuxe+O3+vnlUF6s/K5iacwXl
7XchS6EJ2ROiO7NFs9qXt0G89fgKyN5I57kqFvjtVw8uTBYlPhLA2BHbL2+0uG7P
lSSnPjD4RN8xdA+wbqJeuNIWxKhS+EnqqTwsqPAP/D7FjGT97uUcIBaOCUNXPlK0
cYp9Of7xIsQUeCtH3Msl/sZIjbt+pivIZcr43Mwha1Nfnh0+vYDefKiweh5N0wOJ
hq19NKyzDLW8dsl/XSe5wVB58LEu1hefqv+JM7oDix2yaepSg9aJ3SVtFbFBDr3Z
p+u7W7IZuZ9iGE4cLEHNwIk69eiw/2IxHtNTaNh8Y1cGEENdsREeN0EURNozpHrj
g3/7V+WjzH2fKceLTl49ke8sGGt3whu2WqF5ypS2MKskYNeGLCTUp7pvOsUNnvga
RPXs9PvaeoFu6b/lroZNecTRbzHfQtgxCgumYoWdFO7nu5WEsmQ/zTDuQjcpujQZ
UDd0oASLbcRb/kD06aeJ0Ck1urPeEVYGngIsFWrjgj2uMB68gzEO6pFuI3LcpI5z
FcZKZGiikzHauliWZDgCVJvbfmHHWfcYdQWREKxijEjNVsSLoozk+a4wxAgsSP3N
8WHBhSmeA35kuyhtCJ6LgExJlEdYDvxer664ljNcHqFs7nLjesrUxylN+vXH4gQ+
gOAmYV2rAez0omFWpKdoc3kc9YWL2jyuCfAF8qKxGJcrC0YJFFwQcOrRHflE+tNc
qi9hLRqSQwtfBzU7lpEHYQJDuLjrNIV62lvBESq3uNb0ckjIiFf/jB6lkBqkDfNb
+GLEW/vAqXCeQ5YACUEw3id4rLjd4Vm72B89f47ZGzEpnBscGA9G3ZZfVozubW/M
9XXP/HXJ7jtlIEfX2b/44l+hVZ/qJrXflApS+9oIv3MfnI/YEcrL0MWH+NALyXs3
Gq0//84jbEKgPrTlGNix8khkLcezPaA0f+X2ScqRFVAPrX6ktfvgumzbmDGPekiP
QkTUnNB0UamMA0zpNfxse+FYTKbK90lXPbFl2XOTmTyuEETNg4TOKdZFcQFM60rr
+Ct9TbxFyUwsdDWWy3wIU7WLvY48T+8yPktgnFvGr82QZQnAK6A/JqG9+fo/OrW+
FFYAjpy02XH+sUgjaInJKG68+b08564ahEiAtrvUphgz+noGn16itDk9b4r9OHPL
piBGlRcsvQAna5+hCJ/+hTJed23zjoL0Us0+2O5UixT0qIuuNprmPGmb//oKfnGh
e88WLO9yezqdgjcflF/JbQ0SFUMSX+y/Yx1HEPiTr9pPcJSYNNco5G49W/1TRd6A
FHHlci0Qz44bwx4177ohW8t6ZypHn71BNAbt1QKFkpFwzKNROrShtUCy9+7ZZYyr
dDNSP4fbRTmeQ4axc4CKM2NNdokaGWxujRR9ENmYiMWkfBp22eB2xz/FgSR5LJWe
VrnzbyblOFOHTjE3Ihta518fEMQmbpdx4nawhScNmZS7wnDEygVzJSABI1ZUs7n/
T1a441W6aEEDirGuXLXTdspIR4ULxk5qIEvHrs1n0XbfMwsfqZJmyq+8f6w+QtLg
9xn26DmwRqkGYN9a0Dfwt8+P7zccY/RKhphFn2FK7GMoPN4lHbuwb9aFowHAK56w
8NeaZHlPVUvSX05Y9FXW7Xn45sJb315mst098tQzKqRiihjCG3Jiq8m3pF+tRGhT
FGqL0ekMiNQQqsaHJpFxSCNmhX5z0DvFTTyx8KXIVJNNvo60iLWM1UxPqZSSZMkj
RwW99kPsLMtK/2LIZK8lcnUl3KomDoPolRk7V2Sh6pfzNlMCXFkTMmXa/0A3v3ud
lrI7EHutMT8MdGMkreV7sHI6G6Fr8bjs6ADKFMyShDEo8zPzBgKFnBn52a081mmL
V37QUM5/ZDvYgFr/4edNmx9Wr/fMl9sQhKTXC3i0vC/o49ZVQ1Z6I+YeXaIg9MNf
OTtHbea2QDQ7h2/+ECS6jiDN8n5OtUeDZZFI/DBwK6A9fJKWX2Fy4hcppld7VVNU
F3hPxV7B9qwviOSQZS6WCjBlhdO7L45GiMoPPDB3AGMByahMvJqhRfs8BpMvKKhY
rtHaFtlC3+QbcxSXYaJmtWItLdsWvsioH4nwCHoaZt3ehPwDs11RaBKTSY7UxBXJ
MbtGXHuLlrg5w4oLTv3Rz0+A/sjWUkLv8Li3Ry98IRmp6JBTDAJMyTLZfS4mpUqA
Ky4a7oKtCt6Ye0OveIgy7413x6N3K+E2Wmta+fJAPnW0r59eA7hZGmxZcFmxQAlv
/enFmY/PuKBoyHPibOzclFUVF47BGB0zzdSiQSKX3BzOXEXUJV/y2shTZHGCMPtp
vvnWPKdKK3sGosEpWkLXnUW+VTgW3pZ10RAQc2nRe0Zt9JQdXaTRo1na8BGWCnp5
Uvxy+IWzxB6bo9D12hE7vNj2HMVjmo0RLCNbOMI/QxuTgByshwZHIQCqAyQ54tuM
+Oe/MdlBmx5wQZMEflv6JQ82eiNr79tkqqBDLFzManYsgmo7sUxMqFAOaRMicr/3
cMiqjd63HlAptkFRQq8WXjoLkFBmo871QLGsrzR/Fvj8tfz6+H5O0SmgA4sOozz+
j/Xv9K/puf3c/6RsQJZbtmTldxNVI5ufE+1O0/vP3YRArtWjuA/ML+SZO5/g/4qw
kMGhtLUGVblM+8/fGQhgNNaCswziggOfgRZT5C9WkumIgttHxuc4kELErNu4G5Wy
2Es97dYFardnZCJL31ZggdqoNFT4mjAxIyRzZODhLlCchqzI4iWUS3gSXP/BrNlW
QTaH9zrmIokLjE0fLjXUKTWCWwefcVnj6EtzcwAoDZk6zMp4kPFBIAXUZxNYwHv/
/F61UNEoHrcjAVbHNYqiZzRTisBPe+Wqsy8Qe0u5qVAoyFhoOVf3hIeWjsFmjuwL
cRAJ5Y+mxwxnGqeIxjakentM+e7v85TG7UbJnbMyFFiyYL7M9bPHDUk8EHyJmc8U
fHlaf23lJH5EGM7CxbndmVtAjSdINXo1odrMXN00UO4rTIyxaXDbgOkgG9DG/bfv
fiRr5s/u4/2ecyosTLiN+2z65T2H1o+uyRQ26rm2UuUUt/LZTAFNQIVMcz5p6MZ+
1H+q3tcgX9FeGqae4Ph4h/7DTtvaa2IF75GFtb4IlW1p30YYP4hXQTe8nmaPzjRx
xPFaKiPztnSd+d1cZ+hI3gWjgq1niVW1zWSblBpYDxnjYzEltsfq1zFJeKg/gt4+
VghR9vHd6/MKiPOcATDQxKovC3+xAI03TXjbz3ZS4XdhVYp4vlYNkcG701zQsD4D
c1ybdqgyIFXaoyXF0n5rVO00F7P/1k9Icaaewx/WWqz12zQXxjaEqqByvL5BFziS
1dLn1XfEV2XklIqLynml38Oiv73A+MRzhY2wNgpWNGN5UXAUH1vzG1LqknjviO91
5kaRo+rLefcB8BU2zs715ZV6XXYOoUm6gHZxzTYsYLgmO5zx9BJTE19FpzeCYYM8
hqP6BU3Ruot4pDsK1R4erMWtwOzkAZIFkUKy7WpbyByb18TQ+7/CWssLWG0nvuMQ
6ZJsCv6e2v7RL6a3ewiNwaJKlaEQ2XCvL2geU4ws8X79oLXx6xaRgpVOgVPGV7Jr
UyUnQa6I11g57JAkMoUHpEZAHZvPHeYKXwIPXhuUL0bm9N6iby8q5pUNxgc2EODw
yUVfIFbPHW5ouheKD6cuSHEV/Mn6pznkKz36uOkH7LR2V+0pcHSNi8DZTrP2JtsJ
mWol2EyzWGlZrMnQZ/PG7dAqpv9PYmy91CspqYLqOskIIO6rn6z1N13gUIWWBRG9
kgquHDh32Ot3S3gNcuV0zP8y8fWTbao7UYgQ01zYxfNrDQdiIyVfxyOvc3j7cc9t
n59j5o0V1hwIYkqwpYXPSF5fhqH9uGn/S2W5uykK+MQmUHfVM9XVege7Nsf//734
GR2aLHlx1bb1zEoQRxRo9r4uB6OJ4V1FC2dot+XZ0Kafqc+P05GbecDPMKT2bLpR
QmmruXdWwDIumA6elulxV6U+DLhWMBlcGWTayaxAYH2g+lfSKmSHhIR+5p7wnPLT
oFEWMLP5iHsoJeWA64g2Yrbp575HrGXgGDbPwUSiLnyZj6KtYiDYilbNip1euQWd
m3Kl1v3S464pOtP/EncA/P7L0YTzHNXUz/eV/qf1Xng7GAet0oEC0abQwDVNVINh
2mqIvnlWJii8FsephQAhhKbxRYP445JIqcEm+3+TYnXxGpfvpBNK8CMyBsLxT4gK
JQmQ9PhfgFVCZghR7+VoOuM2/UTd6Z2a3j8qyVL1W8JZJVLVrAmR8mfVgh/YS03y
dGZrXPhRHaAbrGbqZUMflul9YmMrfIol6oD9oFyth+/Ng7SMhR9Uo/Mu9ahZ36T2
zQOlLEyjdaF+vaqgzcwdde9RFg+pp7TC+lxsGwSabmF6y6npzLLsBudtJWklTM4e
IaExbWIKNzmXtgZVP1SQuNTR9Rd9qIc2Lzg5ob3zkJEdEIZgXyoG7/Qcfw/LtU5s
eINQqxIm20Bb9PjpyUqz7nkqCb6k7CUc5BVoKs3Qchca4LBASxPMWb33fhAHs0vx
vz/7bV8I8dPnu77GH9DL1aQWBO7lPXjwP5IeIOD5b7Nexymo5GkpeGpB6hhiGnEY
uoQxtRYkJkCsEm8z/O5LfkRVFZ/QSjfTf8yOu15JJQ3Ujcb6mHbH8+fsJKSL5FkF
i72Nl02OCrmoQkMykbB/VLClIrBYy60vY7lPttASqfxxCx2YaKNk7CfFS+EDechL
zW1+d0EVj1G7QvFio059c9wU/8bVdtOTpHfPmq60hOSIMt4RS1Y06XMEYyvw0puG
6YRxJmUh0ucMLyP9he7b+edeRwpdTEfhPWv7i8hWBc/0GxU8kl8CTec/IJJZX+DM
Dlhc1yZJYoVfT/CjdlkCu84SM0a7z7/W5+kaT+CefyLtzWY6/VqGmig9dgG9E3Fr
FlP4LotaRprGSG8tvT3OnLoFIld4CjZcWvpm97N6Z+b2l0gk2hXaKbMPLcdl/di1
Mzru/n1pyCiUUBseKwCX6H6HnwxEvRa4X235lvRb08w/0Twx0msDhFGk1c7xwkgs
9aQqkRKgi6QYy0oNJlTC/GHyAV/RImH+cJ3nd4J4qTferdIB2c3DR2GeVL1PUz5s
kQaqT+gO8uSZA/1fP9ovR72ZjEC3cl5pMPOp2a0eTQFXImQ3LH99m+UlOUVT3/ua
4EHIC0w19yo3qnyjiHgVDWZKuCishK9Mb69OFYaZ1OSBw6NLdC9Vs9LRCaLJa33q
4mUD7P7679N4D4OXr6WrOc4KC7Qg/l4bTtwlauxAGEM3VQmer8ZVgajyfbK1n7fr
G72XJO30XGWnlOHyV7JP8Kc3nW56/oMK/xHn9U+9uHyxrVI+6cURcdgmjUnBwu+q
5C1r709rGmD+phOqQsUaoGQI7TMnRlpzrcmtMdOUvipV6PLWzgoIDBzCouqwmigP
XbagN9PP4eWCn0W0IdRi/kevbgI82Nc0CPDTrPkIRkY8T4B+oYmf31C5H4PnJjX0
WeIuU7n6AOneU+zjqefMNv1vVd8zKzy9wt1IuiLJ2redHxRw28tVAqfcGx5LhbGv
z4lYTpNpX/WOiu3wgbmR/JKw7gfUTjzFfna3YBrtKj4B2rsO7hLkrkaFzrohLEjm
XjeGTcdk3wqoggSPDefHZVnA4HptyBLQt/u3W5W7AhxSMNF1asTv73dGJLidGBLp
pYRN9FbrN4icFbpdh+0OaV2epb/dITCtbJjY+qTzoJRJOMDiOUtRVhtGiIC4lEcy
vNatrb1pcXrxE4BPrV+dUkIEYyOLx+j0ML8BA5mZkJE7h/IQi1GBYlmI2l3/Rv36
TpPxrcsxTH/qrJyJdJ6Ite7P5q9aREUH8hz2mK9PjazR/iMbjYFXEYZufM+BdvaA
pC4mPRl6mnbpxza8tifqdo04gW7Z7MUwQEjiZKx4E6CIeglvxpE2QmZW437jT63Y
Sccz3f0qeBUwj0jQaOnBUw6lL8Zxn1vEwJPrkvNJhyBoFm3McCHo5uNa+rq1REIU
PbeGXcgv8E64+oQih9EK5Byw/EQXtAmjeaYOUsiOM4Q1lSl1/tvVDy8f4a84ISya
8HIBxXxX0hcJVTzZokjWfGT47ZuUZtA0NqQbL0LOs87MQkhfqaS3QKFqyEb7wVfu
Rn1/J03RfQKEAAQTANwTfHbp8KTBtZm82mSCPLdwWkV1f6FNBoZEKtOg9B33mcGh
4diNK1ehqy+3SmXmWx0BEDdMn5oRt1FECttuhOuw2IPMhFLer82QetZNxt8V5PiP
V5eFx9y6XFqsEKbJ9KBR/+ZidkNaAkI+UbLlIAFj69N/rr4PivtY8EaemDuk5NFt
y5xfpso57eyGxwhZ0GD/RmvJu/TprYev5/7K4ObWSZVNM0ze2vRiaoW3FP25lKOM
xxt6Wl/D+6NgazySjxbWeo+Qv0zcWuAJfR80orPIUoLLNZDc1Eo8XnidZkvaHwby
slmpqZTVlT/fStCXvxDon8El/np4Km+xltguI1W2rdFpsVpLzxaigwhebRMsup3w
rX98wEF0zUXIfxLX3OuW2S/GmDl9AJSwJSXnZvfslbM80HbhNVlHljaVPmuuRkXk
mW1DLZ4o/YGa6XOv97EB4HES2qHiVsPCfdm7uKfdVOo03v/kXAF4PdF2uWtlykNI
PuMVPkeSESuR20b1RQVbHp7QCiJ43nP6BkbAEo2c6CKsT0B9HGqtKfX1pu973Hhr
5dyQY6Qm2qUp6qUh9iBE86SD5i7kB4/9QefM94gUnkdo7HiJw/rlebiTIHsx2Eq1
KNjMN8Fif7X4XxIfiVgeuRwVYHZwgZ//ev/wwM7bcMBdj+gj4zpklzjvEzf/mg1o
/vCNGy4OGNKsKTUkAK64ZgsyJeIybT7Y3tH4zTu7IYuTovYKUwoD0khSRtuGa885
WNmNCp3wALGW1OXMAPEaDk66gdabvDDhFBsU2eMu5Pz0wHAxrE3pVaH83LaoUZVh
YcMQlPeq7RN6OyEc8CAEIgR8xWFMiIrqPIgBMe3+s2ti19ekNNnA0VkHqsb3HRT0
Pk4MGRcVMbmaQrLacGTrm84yRJHV9ytjN5KxdjJDaWDNpuOFCmQwJyQdVrZPTVt+
SqauSbLvsUkaEq8Cn/7pr5KLKrcRD2W5+Opuj89OgV3NnMwAu04biXqDM+eaRdDW
WlyMH6RjQOME2xVzNwxnUCScMx1qx5iIYYAi1RX6T+4S+P3kSJk9bFhlU4P8cuMc
eau0ZybVh6RjRBIDBPI67tww2vDX64WbL9ZBMNHSHUG3M3mG8k+yFr6rWP2WY+4B
/aGn5ZAxmZoFJI9UvtCQs3dY9+J1f5bSUmGPiGJlETNCt216V0WuQdqgAzjEvoxu
4hEMpwcPPvPyfpLJ/eNPvAdvwKfm/2EnTIUKnroktLJ5xni+jZz8/mxbZQSNYOJ4
kTkzBDDWZD2Z+lXGoqI1ObQYd2ZjW7gUWhq8HlLd0NrknCvsoFnFdQsApjN2JR9E
z0o5BvBxolb1URD+3AZZxUAq5n9sz5VNK4MaXZQ8fcaYkYNh1MZWu3EJ9miBeeYg
lrxfZ6VFw0qBsVBMeHeB8DKUEWUp5aoomd5D+8Hv9ohjwivZDT/f0ZOgZbJ+rIbl
evsrPXMZ8j5K+xUamJxBwluTcQegQ5i/oh01RDEBuxpnAAVxAZLJBr4lwrEPX5em
KUXNgavxEUTLhDj3fm13IA11kLIgSiImo82WksIc8vqNOKvto+un5D6FYpnSygy8
8f6LkxcwLu0Li32lGUeMdRQbRO+6catAJy3iGcdYPcamtEQ4DsW49kV4a4x/1bcH
laLZGUr9ehPm2diY2B6Gjd+E0wRW2RwnPXVdlTkIL0X3a05lWbNrMtT5cF4eG0TK
x7L7nHB/lDq7SKW+dXtYN3nvH/eo8lNp+iaSgkUgRIHIx98L2yj2OAUElVBDDMmn
UAMKhBZl7i7aOE9OtjiztrqZ4WuZNvK8d1ggSripBUXSdR/umMAYzPoVdHi4M7eG
ZozB5PExfuquyVOPdEymUBEwuHvyMMk/NznvJVrO/NV76bhct3OwIeNw2Xfi4sP/
vrsgyZZ/3nzry2dYpd7kg6UwEcLczKmGIu8F+1P7kscbzTecowe+bYh+FUXm9T1c
+PbHE/QB1MCPyhLonSA6aBM6m/rNuxRtclWefW2g0VXo0QTqjbkO1ppQ3PVDHIts
FJv/No35Cte3/qPMv2f47jioJofWo4S9f02uwLkREHqUg1fP893hqcqwonLO2iQk
kNNu451SWuUBye2aPe/VdnJSqHxKx+8YUY6KijhRGB6bbUtlwLs/TGofSBLwTYxq
bw9mFUZcXRSD5VVeW3DhoVXh4u+agPn3E9qVphnyw9UXLt9zUCAJHiXF+ny4OP9m
HdgcoyW5e+duHU5p0aufo2pOnucDX9ksYPUhZc/WnmDhY3r+9XclJu7fyZ10i+Rd
t0sSdkg5ziX+PFC2npGVErkbdvUDzIIVDgg3C+smZjuHSA82zUPM7LJPu59XI4a1
2E1tXpzodmfwmuehTmNo89jE8sCn1L+ViAU8Hp6liCa0AIWzN3POvT5ZY97JMhaR
pV4Cn3zZVNioNef/Ar0R5toYMVmRYBZ8Qm1dV5R5OlpIyyZS7qplksq1YZb5TGtk
gvqlr2jwvwEueg2P4mynnnnvuFAxpajcud8PdKBB00DuA4OqCh/2qpZeokwHXjjr
6lGihS+H6qBgEbZY+4vM2/e39yu9n++on5FwNK3ofhTUD3FoQ2xZTPsixrqnbkIe
kkXjRsu/LD1kvz6163h6JtgyMKGRRQgUR2rujDnubKbl6+AlOFNbP23B7CvsneYK
oc03hIzqCVnxmn4alT76FkRHAWAVgJfqYnGdAoE0uQL+sF8ZkkJD4D8peMer90eG
X2ei53eJ2K+hhHLJhmM5QJtk3Ju/b8o2JUpVa4nwi0PFrbtRbcLD2ZKJEkR2L3dG
0WL4OSXnBB65FO65Qlr43iVzJ+3Ij2f71qS5TEWBetXhgOT3gO0kcrmqmoIP4JWT
9AAKAm1Txwn4uKWbWwI+/gX5kBsYMGe8hmJGfrOHcOdgMZswThMumpQO7hdvENTq
/kmiE8peKNkHH9BbgE8rcVEjTmfNoMgbLOyQcUNz96elw9AOik9oNgWI7ecvwUXi
2v9otkAfFNWxCsfjYXOjllDfBbv7sQ1nC9cIQ0GC9J4+Vp+bjCYUZ7/UNIRo41Xw
GhQpPaC+X5KgHqbt2e8qixyLlu3BlqHo77yyx4+oodxeYE/lIXCQJM/cyE6odcTa
p04J99Jk6gim+7UHxcZDxtT3QC22GrMVeqZJhJPc3asVM4UR2d4JMoMplUCbx51p
r92ouyk1rFtEVMJBHxReG5uDZzAK8DBzESvbgaAVuB0gsd/GIJLPKuiPrDp3no2A
h2JxNxpD0hKsEmSv1DLDp1HstD9Oupoyw0CxbDGiUGKRy9U/jE2pgmZSiZlG6+8R
gcoDoA/THOu/Sqhzn8MVwSxllLRdJL2g5xlapaN0W4YQDQeZhSduE0SvEwCY5rJU
MaCZGJE3aIWvn7wtLReOvGPc9X7qhnXoBPudDMfrS1IQqZBsbuIQbh5zsupP+WeC
5EuO3oXduz7WrqswXizkCUpNp3dgRBdIBPMmR9bKqXc/nsqoy7/ezv7+yOq8jO7S
x82+Xy0bZBHkBxFG3gnKfDBXxpacKgLA2bu3lMHSH4qAtWaofap49713heRxugUo
K0zuZ2u483hCY0dgvCgeaKLyyK6tYDcQrgy8qnSjTcvRV+ldAD0T5wVu1i9Hv6Wt
pxgY454NVuYEr6c3YrvT0b7SoJ/TCxoBt+9krlxkSHpF2exbDmnmyykYzBu81xyN
MfGvB6iwv3iKGey3VxoS6Syiwt8pThwjvm6ZQm5ECYCkv+pN5uWSwkPOCcw0nOAC
Pfe6Nr/vTCAW6e6eeUmkhvc9jPAblUcvEPFyelmK1f5jJ7Ue/ACm3SNErgAGy8gB
t6obXken9ppkSi9AR4ij4N0V9Y8WetZulu+pxVOXjxcC6EjH2kZuvu6hHU7FJ5S2
WZtipn5OoSaeBvMzO8x/Tl1bHoWr++MqMmM3YiSuLdTqFonV4BveWVc/WlGd0Knw
d6VkQNOS2NOGvTwDZ5bR/oBIwfFfvmRBRVEp6694JWJgzmLcV/LIH4qvNM1RYl75
YMglsq0LNRnrO8vMFdAi+0kTW0m3ZSaV0sGFP+MeC/cJ5Q+SyvfRfcj8/8JDTN1y
JdyPNIoIcpvdne8ZUY2q59bLB15xuF48PzKXzT4QfWUCRa8ff326kJmiDxClyoox
+/fJnyYjG39C3rZ8aWUcnvQD91NCEFscLZ6xHRA4BnO9bWJoOxKvjEG/sI10/s5y
+l+ciuSKz78Rmm/t0lbxNf9FMIkhbBJArz+mB9nFMfkspyTWX1p54WptCY5mtvE0
ew04zprkr2es7UJ65LlCOI7dp2rM71k0pLsUwRAdAA0pZJoHnZTQxD/NDtfQS4KA
bRjl2U7UG5D4FfXty2+siPrm5kMu8PCYbToCNPlwYgP0QhviIl4PgwH/+F/BPJTb
emkwDqLAfQq0l1eQjbsZbOC5GX2iNwmZDmKIdWATkKm1ld33XcU462EsUOC8AChe
H93VKqIWGdg8bTj8HYXdpJwS8z5/rPExmeVUVwzmKNajmRtpEpLcDfrbc9fPtgnF
HUTzBdlH2Ol4Wj7CpYyg5PpKNt2koob9sYyA0DYPLq0erouZl2QyRGhjWq/6dN5+
paTjIxm/kjhaT/9+j8+JvCON9m7Vf5T0hJklivm+Gjpy23PmQxZH59yF846pT2jK
mTDQ4Y+CzVECKqCJOOcYxGIejOxUGC0Y7Ll3CB9vwZ6WqsZgVER7s28LZgZSMtRo
QBBL4f2vz9cWxFpqeYefAZddeZEqIuyF+s0pHp1+oVbeWwCoj+yKExLGl43jKkfu
Lbl5lmGEdWwT+b8HwgOwVP9msrmeo+cjehwmI9zUKpSZCzgSR+K3sn+d5PdLOPCq
dUig2SgQzAPzw3OzhQ0EXXn1AuLksfHOn2x9rTHtCLsVBhM60ZRL5sV/u5u76iH5
gye9knOnMn8tj9uws09+VRqHpHa2ytuNKwKf3+qPm8WhmBiGxnJgw3q0WdqRXoMm
dfDfNZwjggJ5Ua2ChnvmaCk5KOudozIpPTFfE3qbXEb62L/Sc5hT8oPOKtHtEw2R
xXGG3c3mgBpEb8GkEG2G/FnwuXcnOILhb5iDx0sJ5qblXkIMFGh6zUct4Mh2U4Cw
lIiuAucv3H3b2ijJobBZyXyYQchTut2LkP2rSLMGwh/I7j9zYlVghWrwMyYon3b7
pIXm++pjwSPZ8tMfY9fXYqx++3VP9nx5U6p731S8vnIf493end0ah/ydcUoFKlMY
EqE7YJ0nki9Q/H/WQI0EQUfons3fu3uPG7jQldH9NAeCcu7LktxfdXLqYbNkJ+X5
SOS9iKwEnr6M3JhinUwCRtFAegUUt8Rv057VhKCKYknO/7r4yMMGgATpcWoCqYpe
iwZ6TwhOstkYRTLY1RbUA0R1UnsYPA6N+a3bGbFNSadADltXwNQd5vAWBLs0/6uS
cmVLitpf8rgFI5gn5g40Isjcq7R/DTdNl6cnBLNvhgTrT9Vv/mQsxOOQ+7Olq/Uk
0b54uCV9HaNIPgASSrEdRG/9RQ3emO+gIARsi/acuU5UAH1PvC7D0LjPxBzMcUKC
ITfgIrNp/ErpIbkCg+pQe+d5dLL/6eatvRt/iEOG1FHS2xa3efPhRW+HScvmZsVc
JvE53UsGP7rF2agYItaqIDr7VY/PnU1JWizGGYYuOgF6maab5KOLhHUU3bhZKeIk
Y85P+DxQE3wiwCrXKZn0AnEEia3I7hv1V7Pfjl3Z3fF/V0Yvs6WNH+emhxjiJTWQ
r+upLTyfuFO6aGExCA0Ihpboq1mkpOWcS0oFQ33mZUW7myEjm8YGayGHuJebNn0s
3/RcbIdBABJew0jJni2jyfT7hIQEVmjmlf+RJPhOeC6/GHPV5rRF8iy/L7fc82qQ
VQYB7FkhH5ZpUsZwmT2+FclkCoYYbHSkon5pW6u+wCFCntfR2rNBZmkZsQy7mdk2
xZxDINFYPmN4DsiFsO65vMIdoJ0wQ++ilCuux1ncPP04v9+ldKT7JknG1L9xsYh5
O3E9rBvHeIKJ3hkKMkDByeoIAk8Rad8rLsZRUSGxA+uJhl+JkgqaFxdxgFnewc88
vO2DmUBXXsghJasPgMC9g5+tDpQfMDHBsAEu3GGBz7K7/+QUXeeA2SAKMP09E3R5
tPTql3jTQpN87Ck1XWnREhgMwjWconjzmPMCA2rxBMcpp77hX2PIUihQCO3/P2cr
O6QfnX//Z12Os7BUKn4W2CWD+MnHzWFYlRnwbLrYS1d7S7BkNAsJMjMVCujWl3wM
MLbuqr/tAXrrEmRsrgMFlMCFAu+s6kMe+Ulvg4vFs/BaxIMLnRJshcEgevkdPOG0
U5jSK4Rz6wvxwKu/iJCFf4qxAHTxla3iszH8tkRi7TR8B303UZBaAh/OMH0SCDtT
TKnpb9gE1KD5s3fA1FekB725rEbMsRCH1DWQyIXCZL0xBNDRvpgdADu8MSGrQhtW
mem8voa3GiBeZQfrYYAod0mRXiltwKRN0mTzaTkHVyhzieLUUXg7wHa4oe/VSS6u
1KwjRvD1Y7l0uDsqwxTpyZWVyqbiprr19q+IuqEjbdqQpvzQ8sLmwHOih7z3WMS/
h0BM5taTIBdgPpM6VC4FSJF1Z3FS9lvN3h939ALkpYboaz18WBUCIoN9luA04gGC
icKrWuR150B42HtJZcB1lltn/FXue3rbycgH6RqtZuPnAVvOK/Ys11auQ2kAGDrD
njlvGzIF6/GIuhrvDNPtWlS4+II/a6P1nszP1LIL+ABGV0aI1/yT0oEN8+RV6tdv
HrUrZ5O08Ct8z7kS6T2qVKIffOxNCmo71fgtDTSbzJGB/UXidUE8OuMWrPbhJvud
UC4dlx9eDwNwu29tWgVMliIod/L163aigq0l1Uh0dw+ZAdXVMa9F6T7nqOUuj1Ox
sj9B7jfMmcD0xRLEerclfsoD8IymJ/nZZJs7UHrsVfuLBDKMfHnEUTw7fACyRoCJ
5jQre7+mLLbgHq6Qp4IiX8Yg0n9udvlQ87xGeafpfLLirz3pQWWIsojJim2idcpn
88mu9mxr8Uh26XC9BFE6xD0qRiKr0j2ndzLecX7bkgjAccGFSIinFk+R9mdFFHNL
2rrdMLorESLTQgKyjvQr7+dfgQmhk1VrU2SiNOIMwBKDdT0Epygz1YYlWWacPIlw
dl9A0Mp8lE0zKfRyadNc/iVmx/JEH6BjOFu+/WYmpZ+0EPfqzVGQcR97xKhr79m7
ZGN7Xgvry1cF89pBLs5XsFvnHMlzHCdW4RNGODT+ZksxfheeuPRJu8W1qO0UJBh2
41h6jmEsRvJeRgM5Nv5NdpeSM6m6qETBvnmNWnryOY4N1MJl2jcvG7L47IDud4Ki
1yTvN5CkAPNB2KKWbAhk/Ew94DtLkD3TF8n910f+6qeqnHU1uaKV3ercjEFbGtzp
GgRF/RBknk6dnpAX0ha76eYjItgKgODw/OreW3z6QtVKbIHXf7upa4FztMbaAE48
HjRiSEgQ3HAoGwKmdugrel4KhXBih9nRYydDrlQh164TYrA57df22/RkQr21GwWw
DOSX1VxpbytuJ3dwECn5tL/V9XgYCCZ2xxM5C/HPUZzw8PAIF2soL4mb7UCVact1
occD2V5QGRBwFBohx+EcXIe1FcN9+WMbgot6nPZu7qvW9EwNzE70ZpON/AWPWtRb
gGxoZxXtmCVMUUrkjPGsCgZLjPhLPSWaJkrnnm7Emww75k9Gq2PCacd42OWlz+1+
/R268ZClU/2EebdoyD4ClWhZSSJfICJSluRc8xFzYdqjv438H1FmlAHBgCGAdpOL
zBtjfBXp+ySxWoJ/vd/oFHpxEtvkz4BbIPOaZFLffDN7bEcKIrceW6eJlqHMxLqd
FvNLMKCCjfcv8ueW/KlgwKjhbv/28gd+U08iuQd0LTK2l6b1rA0QHzYDy8cipw9L
qk9HjpJpleJ9YJr4MaXEY2cTl6KzWj41+CxLFjpOyd5oTE+spyXHVj2rjmyLvoS3
QCMnW++lhJ4AIPwOrsb1rlanIyOfqoWOD2aBgxIYBqHDDiYJ5XulI4PkLSUxyXui
5QhdGzhi71WphGq+kLBfJvfFRrHJgKDLB8TfvhIGmfTPZIG1UQFKQx2YM5/4T+Fw
gN1TNw1CswznxD0h+Aw6KV+6s+sUCSYieLeI7QPsiENNohtoFkdkhQ+ZDU+D2HpB
Ypx6czr8OfKSCbbtOMl01nw3IJRLgcGmxmMQC1RXCaFgRFB+7fDXg09Uvoa78wlP
+NzsZXKttsGyE2Wn6uJ6Lah7zgoZOrdsyrcmcOR8sDUaybQoIoXx/+T30UXooL4U
UuxsJeQPZ/Y7K5dL37aYMC6JmK/ICCWhwraNx1LXh8yyKF8r3AWOaXqDU2hYZrYp
KjF3lGS81AACsJVq9NVmff6Qvl7PMUncmJzh8t9PPjaSqXxl/ZGnBOk+Bljmh4Nf
iuPi+c1u/50ectT8S2KnPlp7l2fxGGPR/e+P4L/prSQCpsI3YHLKrraSBggQHUrz
jRg35G/UlmGFRMakpcUIBt1DU22XJQXi/HMXhg7adLHxbDhBFdKqcTkiFu33d4FS
lYI9SArex4PmKdFWEXu4oC0gPJPLSso//OSNBW3ynfnazNlj8H4E6+Jv5x2cOv9E
t/3wE6whk7rACxsxrhaWJQ6afA2UcGS2ofdbw0Yxp5p51D2SuMTgzMXBxjYOjHaO
kiUBQakVmmWf3HcFvQWsEx+O0LMYtZ4sxf1i23XOPPhahhc9EAdBfDoFCsAaz4zs
3J0KNrZgEbwLS6EjTcPJO1pOwWgyzi8rFYDV7n5Ys5nIUy2szc7/ufJ0NosXhdJO
wkq7u9yvr8x3a00h4HbTKfFMlboNijMSZIhl5/7wOZyu0N2doC2YgVzW9wA1eD3s
8iD5J9FWFXwjGmwLT9bq4nHaNuXFeBwhPyD5FUHEbM5RHsLd2b2sQkJaPXX3uPMG
P4y6uQvY0JCMVjwtzXSfXo9+z3R3x4VG0SdWel70dQxAVbF6zGmc/A+kgFz9wUxU
FTXj3L+zMz/Rc8LMZcS4n+6x6WSG4o+L6CH1NePS9E3I1YBeC3mujHoYi4a3p2yv
dLjCrhn8TTE8aS3f4KB8Z+GNolfdx8AnOWEgQuDw8XbjF2dnkQ/Mr/9RTwERMNwb
kKC/C4WQVbOxaRGRPEl6V4s4a7zM7/A2rIrSCgN6hFszlDGcOiRuQsVLjrcGQ193
oBaecuHATvdVd+ivRPEOeVmje2yluideoiRjTH3jM9nYu6fOTFI01TmOxNQ3Ktux
zuts/e90MOaXE5u2RfU+mHSg2wbcrhXHmTEhimuqmKjSPO1ztDL6mSkoqWNbPoBb
icuvbDYtMsEANUnoTJySW7GNMe/IXI0gAk5S5gHYzqLACyCjRgE6vWKzn8v++XKi
ZY9glphJ9qUO1KBrVmF91jF2YMMt64SPvbQ5IWAjtSyvdCuaFvBCm6D+//v03t+b
9i6C4RVLJzMrVszAVCdmPs8NSpQdKdOOFmRCiPRIDt7JFBaaoTmpwl6NTFpzO5gp
hZKoTdpuBsFCL7J6g0frNOHHLXAAwQq8vN4lNmHzbMEMxTLbCbeJDTM7eT7Jsfvn
nP9XJkccKdX0tyblP6Z+WTuOlSriUOMzFfGHnxLqgqDaWtcl02eh/Jfqv/ZByj7w
cULsPpGIeytj+P5aDO4yuEfkvOiFMb8siHZakG2qOJNi0/PoqZZpjPYZGjPfSpn+
PseTvlDXfNlGjppMskrAhEbJgICvQ41hyGE7IRYS8jMLixn305uUBnnTM7v6Pon3
PfosYsZqJ46LnHnz0ehYByFtEWeZZT8QOjxuNW7NN4ImtvV5tTQIAYxozuvzKa5b
+Fx7tDb1bwDR2Nh7XXb4c2njYNlMMzg92xiNklY5K3b57O6IUme1g+ohNsPc0J30
H3gjoWgPhtamriuwltP4E4/zI5cTRQFf9Cr8szCmyMGdz+11nfdWzvDOee+i1/fA
QXUsytcxqX7v2WlYidq+ySPhdYaZ3InYPd+Snky3zO3+LDa00sngW/UezPGOElJA
n0EIAtrlwVjWzcCDUKqFyaPktwFDUh8kMfI3kmGj21Z1xR64lHTRYXH78NFxzqrx
QaVzQxBSvVZUtWsqotOlxkUl+xNd2SpfOSjdC6Zezmml+atafZU263ClQ4LqLzOn
l9fz8wKx5RsLA/58vd+vDcbewru/cQZc+ypCU2Ei+JkO4SGw0x/GGMd12WSnIelw
4quuQz6glXIa3wL6nr+HZrUAvN2OYYjEvLveDzc5LeG62/dwZxhTZIKBmWua3I/1
sx/Qw0ev3Dn+fb/BI709vYoptS9tNEQXziQGgcZ5C0BOffjYJeoPoUdmN2UBzSkK
voRu6aQQ2CZZfj6NokmVwlqOkt0HMWIQ1iKjJ6BDvDTKb0/8O7Qu34zKqGwItpmC
J/vEddV66IcSInrVC+zqLnCN1YgIzajdKojFwK7vekWYDgO/xgcjpL54E++gU+Y9
dy/p1FmAHpohrPk7oiBAu82t7uViuv8tTDi9cgmtH1ZuwDwh90L4b0ybf+deyaeO
sN0suutFXlUfZsMr78YUgFUli4PrmYUZ4rhqj7/nMl6R8NifvvrXzhgQGjoj5CXv
clqChfN5aN+TrkKhYrk0vLjX9GQ2S0bYGtaejbhkhV5VhxZdfx0LnNKFRUfgTgIm
gCr+B9k4XmAHisVgNMRODS99bq8vXYfFxTEcFDfQUv8vy4dO54rWc/eceWYEAmlV
bM7Yg2uRu/np/VTewsXsl8Dx6WF2xBaAUSUjSGwddkJPLrhIwYvEbgmCL+PL3JP0
vhcxusTjIpSpWR8wWq/OEK884zInPMWc9/CjtQU5q13+G/Z6E0TATJRkTtv087O2
UHQihPZagIhe/KBs6n8JDUeo410kMqJKaq7z320QndqGdt8oiKHJgC/uvYIardcY
grZWI6cMZSrGyZJvI6esiHQdghac/YLVKVfEfAF2sCt9O/2qfhchSPDZDv0bEcmo
L1RdTI3o5Jp6YY3Kq+olfj6q/5aahIrCDIYl6rucTjY5jYp2wOM1vU1krvGYMDa0
ECfGgQg40yjGGl1Q3edquTlMJZG3/DOUc9OOoiD5QsJXQlR7kD4hvSP0fihDmCny
CNJUCmxLwJ/PQu0ajk/znpbLlBBeRb5flJ29MA5aM5V3MlNR/NPXTMRhOU4V7crk
HpnHMYhQ+7IbAOYVF2xAbjrXrBk2wradql7n55k6A4Hk+u8eRNF49EhMwCN1bv2R
zBBX4V3uyFJNfky8LM1h2Ys4QV3TL+c2p4X/6lSAY8Sb1U59UvcLG1K8LCMp6EST
mOMTT041pUhJN2VGHkeo40abJaUoo8l5KBIWagQ7yDTjShi+gCrSjoZXBrWDEwd5
fIDZxthgAgXF0vD7+Hohu0G9phMtkH3FfbWEeLhcAKQz/c2j3+EbClaz4sswzWFW
F1rEzA7rBquNFUUYm3MWavNIlnAdqMtSAKv0MUF//Wlq53tBDrpl021s+NgX3YYv
uxx7GM4S8CWu30dBs83UPsOJX3J97FsDSytZLgK03nio3GzvPHgdWMm0vcjJWPib
DXkpCuLlt4UAuPyYUPLw+B8iFelT35UBZqT275eCKsocbHjonkxWNUbBeESnb+2I
zwi5SSz4GehjwU0OOLYuUoMhD9qZW0kkv9JlwMv53U0oteJEklAO6f4q7QlvdfhU
euPvFhoRxwRREW5OuZT7T0tQ+wVEOc4K6WwuwKzUq0zuHR5KEHQ+G788Fnrn2zd7
XyGYfSI001lhU/FHvExnf1/eBeV3US5OWdGIgJSceqxQHQyQe1Gu+YuiTnoUHmBV
qz+mpeXO3juAPevbOTSl4s87JbWpcCdEp1bv8dVXJ46Hz0jBia6XLi64eg7hZu7i
MC42Vc7E/QcTAFpxVcdMRT9Wt7ZN15xJKVYMVezQPPhHGKl3x3YbznSry0EeH+3D
3T9aSsVHpvNhSACy/1JI5zoVrhX2q68loHiup33JmxH4SqCqrpLc9NqRQDf1/TUq
XruSs1SRhZMnLtKh3o3AqjK0DDYxM0zC0f6k74SNJ+o8jhdgh2KXE80hHUqXGY6C
ZvqWawgu+wyujOp2NpMUc60ypoJ247Ga7xel6xUNxctw20CH2Huj+2rA0ruPDgSs
FqJ+fFmRabmSQ5iauOmKMalpfQVvMfRlnJfFM6qIGGckefS53k4Zfu9RcSNYQ/CK
t4sm3nesIbVZfAdSwpza7qF5aenopBB+H730yGQHrSTkGNO+DsdK33EtfkFrTD6p
94xFc4rFrcM1dCadaFq49hInpLHwIa+ab1bTeTrVplmn28rSeJD1nlnffpC2AYGr
oUR9Xo3U7IobOr5/c7e4E4a3Ey/yO2t6AiwNgeKxzAI6ACE6fdLHLEuQlUU2VW4v
9pkajAn0FbKVSUS48OsXrdZlP9gdraSxiLkNBnxhjkopgW23uJlru2DO3Bnku1eF
aztS1XIVgW8FoGjiFgI2VNMp0n8kgt0Lts0Ndqo1uXJ7ZAs+fdOq5CAEa20FLoj5
YGN6QhdBNv/kRZjjSXCAWm7JPabpxIVmOAtTiPKc/PZZY/NvjChdvLyHBTg4MjOb
oOk72a7/ZZT5zWRGW5pEU7z6kZbsNBdIGaoNskd6WNRBIbHsAPIy20+XkbF202rH
F4T0RZ13/G6eLsVZMUkp5YCfAfRIfBnRkuzMs1YTuKaPlk8PgcGLTGHqlfpGD0Zj
2EchqBJqOjjiHb7HCLSTYuwR72uxi4jDe7CSnVwOSC5wkQ7qERcxwQRucFHngSoO
KtEVnzO4WCq83DoiXkM+YftKPchbZXz2MFI1+5YY1SfcGluxEXfcibHlRFg+GUl9
cFdJwNM5u5TY5X27aWA5V0P2/mrM99MXh1LKE0esU4jLTGTNnue3RWNDGDnI2UES
nveV0HvEUS7Zn5QR3e4vvvP9/ZnRznpQuTlDkwH9fzz6T0qeWjqWXfTdhteLlk02
Wg5qfVIPEuU8Ewa6AFlsAeD1LYyheWgy6/fnh4/togOHrYcczLgg4yTTbF8XN9HK
hGUpLVJX3VzqZmAFocyqRMxdua6+ptIwflLexbdtLI2H5yTrRs7tzVUB9H37mKIS
LoqlvgERFKeFcutdM7W3L9774vXmTUSxs6CaHvfdo09l9VdnOcDjIqWGSCvmp+D7
6EZdIPe+TzC2GmTRUjO1SrOvYRJ09DvaLkwoeWBaP5l7x6DmCdYhbtxXsFJOFmoY
8LVP7EZSTITPeWBiC+SL2JS31nH+v3c8WYRMGc+3W7Nd2TaohdnFlJBTTM8Hid7/
MyVlQE3QPK0CdveDsrYvZvDE3BXbfyT0lrjnOT4suKGoH9OkoxcpSlZWnzlZSogQ
wwzXocgzUVAQM/49yQstNH6wZxq2xcAMp41XB0VjycPf4otyspOWV7VOyh5aO4JG
Bg6IamPCKO+gQ4tbWzq9eILf3HE5vS48yx9WWItImmTJUPh4MfgkyYbZ3ksHgRrA
31gOZLB3Ph9ot1GBl9nibyXtWsAe+xZSqm8UxSOZkwRhBxpBhC2se015TL2jGeGr
1/d/vTtpghMW4KyHgOkcQtoyIwG9tVkQwOUPHzULW6cYy3qrGcqpYVLb6ZE0j1HT
EIOHwWtVF2hiLB/mfAG5wmI/KthVDHb+HeKizZEZWrcuwBxCkwhyUCYlYRR7CBxf
3VDY252T6PRaxAEK1T2fjaWQQFnCuwSlaF+58XNCa118UmEeNbxozJGStruLJgIa
T843ZfCmeeLUwZoAzd+hZEHxuECoCymItb0NzQb453qN9EHjvyTuMuPY99WY9zBJ
MFPDEirz8bdiQ0ayaeZxYi1v0AUM63V7Yasu+EAqLSSaztJ1CPpPOMaWkq6y9hSC
MZTHsc7kWrVTXPc9Ofh3UGtghlIVJQIWTMk/pYU+Vqrc0IEiip3LE1/6rpuPGKQ4
iaafzXUcxPRmEnstwL3fQ9WfLHeqEZTS7VFVs8Elvj02W7PHcnm3ZN0nQTO5bzFT
4c7sM+ECEfIdL18CFmKQGBqhTGI3sP8Idp3Wo/T4pMkGoYchfzzmyrUAZdy5cV3h
RG25OAaAmfzsLdItn/P5i6PkhOCY3SKzLRrgs2nkd0iSbats7pKJZbabArMJi8pi
Ma48b68Lhdqj6VdM2hcST6whBuSMQP77EkT4unfmzNpeE1x6IFGqnUTVOyHSXbWY
TGp3AtpBPp6F3SUi6ZWhB6eCwnXBE3WrgLRxW+6V1y7q79MzlgUjpj/BPqUMXprC
CU3PwjZiHrf75ZDg9ohhLpPmgsghaY+TysAHaQ+G7wRKdt6lnUDB6PV9VK3TE/66
cFeTyrMJ/AErYM0Z1l57BWfA+Oek715PUMYTdVjh641xlyVo4QNRYFRhCobdYvAA
1NfEzSV4pKxvDnfnEHs8y6r2DpB2xxA1qw03iwuq2pK/L2Op+pOUoCF8Wj1jlyps
PUHuZWlu4NckEGL5bvS1gGLsXXCy5AKB6ZCrtNrjAlTrg0Dv3N/uw0lA9r03quOw
MuWSRmlOt0GFSm+diJG5RnETJ1IbWGEX9evFvgdtJ12TZFg8UeZRe63zwFR2tFSS
dqBBDUoVaMO9BmhrptVHt6R7JTIXPRG7hYwdCknnOTNj8DJnAYxG4m/CiUr26K5E
RNcYVpnQvkS49lxiUlDXFe4nFbfRhc1q7ebnnZXmiOEWRd2sc+vDN6QM9B9IHntJ
eW2QKXkXYY0V5+d37A3rchjJIvQeahifH7aj24dUtD1YIUwRS5LOoIL61haDLI21
4KJfE1A5ab3KtLjMKZAtrMAkGcUwqN8OTSdA9v69qIZdiNAFm0Mug1JomIPysP1q
DGRcmhSnG3KdPVebaqjnTx7WQWAq2SdaKWytIMoqszorai/gi5SUjJmK9ocyiM8M
pa5nduUZjHmc06wPvHIIxoAE13emWN/pp3FmaCP0SQkq3U42KUcGeznUJH1m9Yxh
cxUhqCVAry0i4IHmU+QbWMG0GXvhF9snSt4xDnZ4RumiAtGUIqh8+PYCmp0BTF8T
2BANb6Z4EnEaIs+y7CKtDVzZa45NSeTzaA9zHpV1z9P2dWQuJQjEqeAFPHQKYSx1
3944MH/Mltj6I2EUkOQT73cjslIN6iYeIwgfLnJvDUC+0EMaA1hW9FqkMDpUKk51
o+ydqo9hJfJLujgyWW7XGXEvdIJJQTHRuDaouhXIf2M4NvIgLvaLB22dgTsrgMe4
aZ57SUnV8gqboaC6l6/qI4AGaWRavIDRrnsZoWVqLxgEypbw1x8SIWYT22oNlW9/
fquUQQmY2dBomuDFb7mLlhNtw+sjcIA0AVmVizQpGDOIqMCymxfY5lOczYY6DPt5
aohKP1y9FdhMb+lkt4K/h2PJnebh9saD8xKWndfhbwLINBJ8VAFdajc6wmYsEcf3
lEitMlp/vFhPh7SbMbWQKCJ6HJcKih41pj8uA0ae0oIf1O2riqdqlM9qEY7NviGg
GlqXGjG7QWMn+7j8O5pBfDCv61K5jM0mZAelu/u9Rewt+MNs2ok4fJrpqChVsn9N
GjI4t2np82e3J30PcB3goUBoYyHd/PuBYhP/anxZFqmI4v2EO+TOmzFulz7ENyxk
chOSh/bjv/mQR9ilMpZxvElVS4cthXVjEBzWrA8OBCmfwL2mcZzMEAmFF77SrRL5
CWnsLeYs4j7ajT873MLB8JVXSJ+PypSwfk55wfNMiOJdaernbA1z/JVs8f6EUs2f
SLtN+OcipiKvodpZsIUufp/2kvr3oBVb25IMKWTyf1cbk7ySVqz2yohgdJDX3eAq
x7y7/lBxCLDl/i20u4UiXAcbZtkqyIqc2pp1+A20kk0qppjgSiORp01VE9fMhcMG
mvnnFylU5OIbL6XTOUbvC6fkCANq1FZOwDqTXIPF5beqra9puD+FPAcny4Qyei6S
2D1VHSCs7Hp+O8RFyIlSLry9XCcyXlrYTlk5/EzQ5mtB2WKVS17dNuBGAkXM8d00
P0LgsyHzhv4MktNiRse99piBALst0wMWv36BfKYAAW4V/68D4DItWdB0x6C8ffRc
sdMDCzzrSwxdfxlTrwVBwa3PQTqdzSKRPQqbXNOH5i/je17YjF1d9znFNCNXx7vj
vJH35WUbyTi0n7whiUb4ib4SF5B1YdUmyN7A8Q9PRRWZtEW2S587VsxQxakWOMij
lRrsAVL3BixRMyQWbudxSP8ZU8tNh9z3q8zA5Mc0FvJeJxyIz1270I2DrL9QcTag
ulGNlIp2YDkTJxMn6pEKoQuc2VWq0RGgiwSf/DEcqwXUqXmyUgcSwXWOZMWfL4Jv
xRHwDiKh7mi9/8bi5yiNu2G5P7fuXF4eiLcIuTPcdgUlBhPOW5bFKmdycOfrn/+F
NKr1iToJRZuJ3dsHbdaIgtNm+epQ90COdmo43cTzTivMkN3WyE/waZIP6Xbn8NYx
iwolh3xz97QegcHXfoAjSSFSvQKuN6d8udJrnDqGuMlDVvlI+rOSMrLPvJNEBZIA
8ZIUIcYWTwI5YRKto/kP5Y4qGwcZRGIbd0lgbuW2Rdr/W0aPs3RZKYclFuSRTHEb
wM7zPvr1SzBob+ovQrMMqZva23pUFoEfLT4jm05/sTyaihaatWIidMJUnNrPniU0
syLkVcTc5ZeyA02qivph44Ns1gH83sPV32hsJe7npGfdvynLzznc+u6HCWmgtLvu
vIYBpHQcQ8RqV4croOtzWYkx1BtLgcowMjlzRX/9VLXZxnvF8tVth2tc3FZ8jlRm
nha2mnfXZcx6KcdbKcauUXse5LaG9lW2NDGD6z+VN1IBPW1CRvk3hOxrfJHzD/QO
Za3j3pJPZkFek2VTi6FRetlLQsaD5OBSeHGMcaFzqcqRTQF9gbq2b8gHUAi9W044
zpLhOXd0IUjfW81Z8BJboGsETai6gskdxB4FOSTJKzs19a+q7IXIL476fIkHU7he
Z+eQ/B3RgzXm3hjIZfAauJOANrDRmAEe8aH2p0LNjCeaF+MGhUmDk6hs3NdzGWKz
RsR5owLnh1GAyX7lyzeqrs6k4YPX6KrQMZU63bhYvXq3ccMPRD1XFvbe66JXY1xz
5q9oMraM31+q9/hdFYQCaVqbv7NNdtKeLEfrX/qXp/UsXgDNPzW9aajwH3VDbjSk
3ZQe3ob2klTN7rv0Ezy6ExFnKrTmIa3PqhLBmEPEV4JUkMgKNXHDhD/ZN9hDERNi
dV473PvBmOJv86h6FB/6Q4sqecxwEKr52U+DmtajGxpOiI9RsyEa78pIf1rn3DjA
YG9QMd0YolohfOdrU4y8ZSB8WJcABr+D6VapCKv6J57JfYxyaQ/Ryesv7iS9dqtE
2hghncYEex4b4YKlnGy1SOYbS+NdrDXijQdPd/chDZ7jY/1LMaGE6lEqbwmZ4BHc
skW8xRIIlOxKNA+gR9Q9alLTDy+S+C6ZexqnSOpsJVi59i0EaxMF4mbfoRcIpZFi
LhAP/pouvKhHeyZMeGAvJdDWd2ub/TdLmxRTqyua74w1bVs24rtqjqoi7XR+xVlo
qnhvHkHNlfNejFAv2FxHcq6BwjUSYQqt+RSndW36fStR/gP9zdQ5mPEDnn3Vhoio
/QEK7QhTwgynYqhphgbsw/eN6I+z4p1k3Yn6928fEe/eozQXr2VnUjlhgktR6kU/
ZEfNjRYSEJw1/0SRi3FaolQUTpvXkW5sjbws0kiDDROVJ4YDchH8VXqPWcH2AyT7
uiWt5hJ56ta5N+uup+zGHcqiPVhjHD+0TIivRg2w4pqOLUWC/oRu4/Q89b1+ZrFU
qY6danT1DMXcZYpJWI27SwCk1Is04J62u5l10C8I8aTFn9h/DN8xir3cTT8EMdSi
5Bbr/2CZh56Jtzo1ZpixpnUfeyZk8RdJh6shEvEsp5nFQjEkRL7Tc+xDMbrQCwm6
lbiFgTOVpKNHbjNV3QuumvPUhSqBaCFP3ow5ptnGABVhquuPiPuJ8mA1LjrPjawS
HyYyqN1Ug1Ow0MoEQRtUYfRW0enMJpO8kUceDTiR6q05zKSxPbH6+ZMqdFg610It
wUn5PyU1jNkFp+2pnkNZH7YvKB1CtqoIKpHdUjIt3y2YfN4qgLU4gDddbq6VFxCd
hucclwzoORf2nvbfcV+Y3BZqG3i6UYvk0f0lx8G4XabBdWJkjmwG/EqWP27Qut60
R+4nRvEFASXAf5cyHkB8MGkrA1JXJcoJfRCRgwuFki9glSUzxe5HwzDkw5f+CwjE
3TofCAC8tQAh1Ywgdr2qIaQa4cO8QMX1+o9HivU80/dI8cUQP/19dmdsaNg1g/vS
zajXV9YlfTCbSP/UCBx8ghkSzf2EH0au51bJs1Z2gxbK+wIhRWYeIs2CPlip1ji7
tRPkr66LnE4NNclw06541fswcPtZTqV/zRfTppWCLTmTCcSlMA/f04A9NRqXkX2z
srN2Qm3giv6rnvC7jkprURV/HZp1akmxB4sHFEdPOQdvBwLF+8+pvK1vp2si4QkF
1pZoIZFni9sXwp18U4SJuN3TdmA5f+FH5hT2+sdKPrT3et2Q9YS5DaT3THXvEgCU
MQk+S6gXBcGW9oYWuRVDcFDEHE+BO+PCZ4KuZi9VG+HI9CpmMocS63RopIMPSrCy
mTuGcJo8xIIvN0c21DQzMv54m6kn2voaQRuv2TxmuJi8pNyHo+XQsOusVdHhNV45
PLyRf+MUbJR+OANbsGPaFdfkvAFFoEwVzjoGUGQfTsnjFIZG7Q3X6KpRJbKlB9bw
w8YClq0EGl/NZsgxfXO0o9gZ5s7tek2HBCgwAEzPr8xqN19Hm+PEi2VP1SoZXndp
KXOWB4MVCIaoHcEypa6U7CT4YfAABVEJrLJlaYe1EXMNs4NglWXCmyEfBp4IavpM
pngLI+FBH5XSyMSsgbb6pJia3UW5Rs5FikDPzbcklJ/7omZIqA96zJNzlbMo7o9j
K5mX75sMCieoF1tVmONjM6gGhldcaGbR72sOJhZg2PuLpxqVqjAOXqrmp0okGID2
lEx5axxcZFPFdDxXejhbYbi/4S6v1Vqlj4/St2OilD6vUibcKdjTrsGN6JiqoVjM
IMvxqoQznvUBiVqY9/vwiI5aRwd0XX7u2NBq9P9wAE+w/xPwM5lbYxK3+tgN3zir
DuLqK/1Z0PopHqaCJukf8ipsA7I3kR3uwLz2oVmelJ6lq098iUevAaEY1828sTtj
NEMFxkyF2sgyId+sHNv/a3+kHYvGazbr841OpviVJLtXubLlHGS6PM+YLQBivhL2
KfJvsvGu6W64lzFUVA4UrrtJkm68q2O3+yLmMh1enjXp2KzAcl5cuG9Yi2iVD6Ki
s8z1iGLSz8JEz6kiaPJ4vR/fCrFmO/LrR99sGPkpxYGtlU4elaSJyGjipOqNjCom
JwXB4kuSAHBGTYIJaBBqtlXojRmT3TjPmZNJ2XqZnDuRFPldBadcs0EK78PUxvgY
25YCG0WYpDBZhjNji2EEjGyhdtzgWwE5j5v67Sg5RUz+r85P/FKKkQalKDLlqSKQ
l+l3wxGtR1AWBMUeTN+OF4vPs39i/X9v1GYlnAY1jmsHEYJxX1+KiY0jEcTP5c9h
3kFKLyClbGtXSw2UQvm4nI8eMbch3MIW+YRFcrzeiCZomZAwoB7Tlh4I9b5Qtz7D
Fwp9+V0HU+jaldU6rgUAZBfRa+XfSzt8XLM6XzP1gPr0f3SStn0EkIPbJFT9WsG7
PMAwsxbCFue28GesrU00t4T7SZ1v6kC9N3ZV3Z9hdnNKHoYuB6iQdk4/RMNuyLBy
CvNeAeMRKa9HV0f3qzO1ENOOnNdqldfZTbxnogtE8IZeNbwsspc/DyKh5z8Jqd8z
1A4IlzrY/uODqegeEf8AazD8Rf/QEzgA83e0oI/kJoud5re3qz2fLZeC/x/LkGzs
tD1hgCZNNEerOUUGcr4rFSpcLy4w4cTBsQhOQB8YCK4pf0MnZlADXfxCqxOW5YPX
nVUhgveA5scMDYIHr+qxt/9/JijLiDvia4GR+079nNpognkEmXAVVYdT3bmsJ+0a
zKLx/GTEpc093zb0wzzXQmHDZjht3AG7bt4CVVRJFlvH/6OwRFBYKrQ31V/H4f0x
O3xS9hAi+AZR/L2H21U/1mv3CFmLekT7MpsXesBUn0q5pwhusFM+T9lfQdfFWOXQ
WSYdRr7xjUS6NJsSgJ+/kOft91pTgUw2N37o5QjT+s9pgMGaVatNsGRtvhtMtKrC
VqwJB8SRzLV7EMry6QfUGdAbBikyqTVs39jJVKr4twT30DIH0ko8GY9c0FaFlnmb
QLzUcli/4IzHWl/Kg+ZVx/k67rhUf+97InDuSGK7Lmic100PnsAk1lUOLnNt7qgV
kaXzO0yZpgBGi0s3WIOj88fFqvXoH/3DVXwvPcAJaKl9Yaqo3Sab96sr73TmCiN7
+LZornvFjG2oqUQHWvqhl6rQm39su3DvkMazppG2BicWgWwn3cRJlThW/+ljVyvq
CY71xKm89L80nt+5/+a2cvKREu27zI7Fbq3dT8rXKFCbKn/xvLzktSYGSD2jX139
LenywGicdQH1B+HaKDIbKjqyW+BnEggQviLql9NXtR0Ifg+cWzIVJWhCjTmQ3Xed
u0Qs94SIEXmqqt2YnnjYwHux+7hhhtr23zll7f4gGvAIYbD1EzJSgJSOw97a+MEY
AsKIk8m7jPZ68XXkE+nqt0G8y7IQnZdlisuhsVQLFkROKprdd9CTJ9BG9gGAYvFG
Y0AlE2jHyfq0UObIya1tU5uF+JjTtx8JqIwX2ct+4Mz5OZWcUd3vOy0hvatmoAEw
Zj91g/l5nPDzs5HKFhGVoHiYPSO6Ohr6DyfTATne8XpcVyTUcvrVVCVAcHQIdzKW
//dlWVe7CWJJw56+7D/qFKIqUaVmW8B9ghNBZA01E3JlHVPqGuxvB3M4lGFCRWhD
oqppiCWIzX87oIoPrKrOcElLL8NrX8IKoCt3z693wyTRmV+87HkZwmjMP0cxuAKU
KaBGoG7M8Mr3omoeDfnVnAHdxRF2eQ46X1xATrnOr3P1iv5sNsldtxLqoIqheSKq
HXKoPrLeQsAobnCA0zJlyvNq1nhnsvuHIfc2pG89b9rtbCxYSB1L1Wdc/t58LOh7
vK9YoBzSFvGrBZMmtw7moD7DIYpj2QxExZ8H3afMItSpqGkSo4zRWP9iSLWSkNI5
SmJxmO/YMbegFhaMl/HW1yXKtFrUJqDXV48nmRT0GBpQW51+HLFm+v8OBjKvI080
hIhHQ1Qp7o+WeloO3h10HJcIWfbp4j0czb5LwWCOurAYYw/Ar+H2+F9V/xokiIwH
7fu/Ff0TkEaVmLsCCsBAip4pCGIiw19KEQnSBAAv2MwGDjXW5zez3OSRIv/AUJrV
qWrSgbnBX8+3w+rEIml756DGe5qfqQUjy5LcqdmUyJmYK/lhfwjJbcch66EJSbq+
SzygCCVc4oGwdZBGnkSKxnnMjF8WxOrN7Dh2q+/18ypFk+J511uCYoFxmzjMN+eh
Th2SaKYQaLZ8XHyki8yIH5b79WZy/H6QPT2226kL4KDbZjQpRC6xrNk/uT2u5KxF
pQbvFH046rQd8n+WsTR7GN+OnGbTRiitzGBaqfZPRjh2NM2+8nMOQ9S6kuYXR57n
D1M4DkBVF8rZlYvQd4FjLsoQTb3PgOWpd/hEO2MmDzxKQfNLK2QCtAZ9nEy/P7VK
4M52ASjjAkISpH8/c9f+nDV2RCm1hUcpNcxuJNcK72CjZA2tbrgxzmmPDkkQWSZ8
gEE6eFzdyXYTIDWTl4PzCoCaiUwhQFznLFSHGcQAEY52jFxjW09vgr8ImXkAE2va
uEz9Y8+q7wdBo9ZwMOVvxvgQnJ69rB786aZz4jwB777147c9vfdrwO8+pD8jgWYJ
X3A61j4MogDzFjHSYJoLIB8jmMEF1LIGQ/RHVsiHVbogxWuu/zkeUWtRYYhuxB4E
VBITOSZ/vb2qay1aqAYuohdVvx8xrQW76WCtkYP2N83AliR/YmzmahXCFiZ30pyf
LW3kNhaaJXJlT1b5KqitH7Fq03oErrvgBJ7KQx1d8qKrGB7vMuMvXeN1pLOHFkNJ
egtoC9DV2FcopMC1SEzq1kScvxdXuR+GcaEWDLZi0ua+RLZYGeOjfhEUgaAO0YZJ
puILqhXDvoAThY5ggljMw+oX7gENk+2IAjA49sBlb22vcrHAuL8TeqGtqSbZUTjy
sxBjD8L5N01hW4rSzMuM/yjgdujoyLuFbzMTK/5Ji+Zt99nyez+eLYRthZbjxg60
iH9oqNZzLufBHfUy5Zuhh84DwAyJJDpab/XByfvHV6ij915Ym8/4QEOQCRmGhjoV
57HNLFlwl+zkCB7O2vfZ22+qOMP6MUZ/80OWlHRRzNHVuFGCxAJmZoRPwJpDyoTD
qlH2Kt4l0hcxe/2bX3FKOn/uDglefEQv2CKOoXHNczu6umoa8jwwKeqYu/xadUrA
DMuvnI0/4D6oN+LgtXdWUZxIcdGOCgw45W+qkkhSs4MTKlaFHhr+QGtkVZULYf6v
iDyNcfcpMoFyP8Wbm1lCpEc4JbNq+EspZrjZy0G6l+Ft1IhjbgQlB2hCfruJeVfs
77dNb+ZSUNzeqgKXmdt9ab5GzJgyu5HcOYdR0Fhp4wovF00uD7d1yZ7wC6x/o3QB
mivFzo297hzCz/Tm9+0m59F+RlV9otiF6VPbFLGnS1fGTt7RihkAncLJbd4vG6gm
9rj9Un9U7UxeLc2ZVoAhO1HcHJzYqX6/M/AfrMXxb0u7ABr02dgtMnQeRwpNBSqO
CFkJnJDWVQMLbjrJqhncNCfaY/Xyt3Y6H19gHvj95/zNVbl4lNGqqUzVJbIObyUX
XndiaI8xoViRtgyxuBgXtRNuFJxWPylFrPG1k7+Pg0HTu/UsNo/mbWzTCeVoJmqq
Xd6b4IOVZ9nuZNuaM+iZEkMV1oUtCLXi0dhi0SreExJfkMGFGoEka3Ubqxfws6SF
tiLgSndWPUAxx5l/JfNMpkptuFYs60A2Bst9lBDU18oMEyuVvEifa1+3vm1iRmMT
ruMmDRO17zhn674HJROESxavgxHEtGqDrJ0i4eUs+0gqYRf+iUT36B3w4s+irb4o
MUO/1HUf74z5s4f0epZUiOp1sDBSC1pgw2wCrMFwfbqESA0MwbEmtCvddKZ8GldB
BuaKOypteVFa0ulrlpRkY/1AzrfgPgJu4lY8C866fFT4e5HMUparaeJ0SsiTkc5K
iku8tHpF+cvdHL4/SKz0ZYN4PLk+roatTmCmJMijWjoxiO/AFAk2lWKJmvAVRLcf
8YqMXiTIXDQASYmMxl2wu5yY4KuG3KM19H/Z+ilZ1iCXy4nCX+i30VnZqn2qCp9M
s6O39HJLMNoegxBJw54czr7684dVAO8FqiX5HWAd/rDOwWCekZ1JKZSLhrhh0iyX
Yxpyqd/iGmVzScCQqVDnhkuvl2oqxlxFQ9LW1T04NBXkjO10RjKcLABmi1bPzxQw
4x9zKDnpWWxMmSi3fct00BafPF4wQrP3HAfK0Pt6RsnHvsVHt9jgBNtyg798O87O
HBEJuwib9lk1v9u4rKmkRzwvHUCuUalhIm+AsndqH7d7aeHErEuXXyrtbQkEuUp0
KzmoXfj+EKBofrX5wwY+4XeNOkyfUYoK/sHdJ3bf82LUTG0LB0HIhOsV3WK3IHPI
aqkVt/McqMZPK4OkVO3IMKblRZ/UeYDknVzvaAbgBDYG71LkrYkRCuoZK7L31vRD
1tQhmKPvJt86n8+UgsfWQqEFcFLvp5cDoRRo7ucRgcYBHJ1hbXQ0JB2eZ7qZNEb1
sgTghGmaGjGOrPqIFi2iV35CjCjxIl8Eqt9YNqMj9HWCObfU/osKCC8p/F9+sr7Z
H+1X7ZOYLgI/vXWNQ9a47frPa1D1TIAghl5Bgd9XdmTTc211Vkj+V1xFDgdZyKtb
sl8daSK0hMHZqH6Oz7lejlHNhWQ6Wq/6PB1qLcTR2oZdZBsOTQsD1jw7145AdLZP
ewoYLs0wQI2Ja+1Hab/QmbvJnG9y3fOfA4J9khleDx2HMvGFnyw/L0ySN9qicf7v
6lQh+5sSC8VN7qcJZ9It9RMCmWLF61bpsSRtaPRrYy7z/gFx/zjJVpTNHoORJ98n
EASWIdTQ6DgCqaYhqGL49e9vmKnaL2ySN0btIc+DFWyZxIkUznpBUHMaDOEot9Dg
6hJQYxcLvABucTzvHQb3rhprfX3oCFlK0j8RW8b3rokCloziQ6uyvy0cfoGA7vfy
3O2VMT0Ah+pf/1rRN4dWOgGI3hkEFzsEvpr94juala+x4eI405leDWPU/nlMpHqp
02nvarNw+sEoAk00miDGmviabtxa6ZQHj8c+Wmizu03Nw/h8fpAk0l06DhiOKBih
o15WUEZfokLEqRQQuxg2oNBti8sv7YZXXu9pHXc/f7zJHThkd7w5dztOr9wi+xYQ
ldF+vhlToAnAxZPc9MHXN2fS+kimXuaburSBxDj4HfYmefkm5zFzHxUfqYzDXzfv
errjYTHxW0w9GQ7neRy92TBTDe69yfDIS4KWFyIApXoEsXKY/8g8/xvS0BBH9mr7
BkfHl7daxvWcU/eoAtQxI7dpsBA+iS+Q72nfoQt0oMGiJtyf4j5qOM1ZrECWUttl
u/qoWxwGO7dJuaJkCZwX/on81rmbwERP3pJDTmzV2li224H9p1WU4BkCABrjPWcH
tcaBsyTJafWs9wDGbXVrb1HrB/Ms5irxf2N9LuFxLF7i6XlmXXasv3ATz7HsEc1A
eerq0tQ6hgAMpoiZmJlyanIjg13OA02CamoG6/8YWTlmBsBFb6M1PEDNIm24OpOk
luqFN8SwobDDuI5CvlIbbK79JgFuvg8eXODA2F9SHniOyD9c7zos/I2aGlzlCLtV
R6X7K1xvvdIsmspilg1rSYJHNnBoiWPDcaPMhgaISKQMz5Vj+p4cy3ObP7o2Rx0K
GFYPQThRZfRYEwHcheV3NaMRO46HrPWPAAdwHoEkGQGG7F/iQSxM74aobIHMshLw
2z8TRuQyaMQ/ux5QyucTuX/lIJm5clBICFr35XcM7xP8FyVS6NfyMDojJEaoICEB
ZUY3DhiU8PmebmtfKGsV8y6j3Gb24vkrMImeZ3NIZ+hy6fzD1irOuz6IXRINv9IU
BtQFH7PYRMLbzAvvmPtVUdSrQJqg8Tg8TIn8OP1mW4Edbp3431vVzTm3Lz2DRdyt
EHVaT3u6zaMAE5ygkFHzMpB93HI0xJp5O8tvWTEof7IZtxmeIDZPEyLV+uwUveP6
OUZlpo2PIlwAs9mLHqYK0U86tMgLevdO5lzyoEiHUcxOQ73TgpafMLBygH+c2TdU
IDkVCOcOoFnWF6XVrYcWpTBuREuvlhx6kM4Y4NMND9h9uaV5seZ52KKiYepnrT+4
RP/UQmzUtdQjasHCr3BjMECyAWOwAnnRIrjesiGwLtHkYNNeZ4Paq5gVcMmf5wKA
pmJhtHVXe1LHj5dzAK9/iYQ/Yk5vl7h7pgVZ1ll5avLExfYA+ohH92tYN/dO1nQQ
yYzbxhLrgijUK2fS8/EDnePh7MEH3+USwarYdSYhXELh/LPdJaXsIdeX3OyckuKt
3FU6FUz2Hqpc0D6U6ObXJCZPTVmBNpFMz4yvEhqyIyTlANweqBv9f0pAsA/99pkc
bR+mQ0sITA/g/r+MlO5UHQ6OOZRU7exKIST5eRbb+xgJAkEjcmeOGBUL/L9TVp8B
itGMh3OeTgP+6u2OYZnByH0yMtlqftQznD1BUtILDMP8YWvjDwE2Q5M+cq3TXKUD
h/MPbg46sgGifL86IcTF/Rn2WEz+lZt/Vq3PlE+AsyDedSUCL98CVo8Q/ebb7E0N
S0XiC6cd05aHalwAPwMFuoncAJtui/vLdrQm5uAOUccpzkStz9urLe2BAGPAFyo0
KsIHk2W612iNCHhz+S1HhxeYCQkw0q/BBH36HFlq6SRpoI1uA3zBC5QI7vS3fHPC
+bZxVXzMehH8Viw73NlpR773wdkl55HrNP60HGH3Z2xf/ZJgKUAbNeW6yKnBpajt
JN5eAj0Q8PAuc7/NujUZeY/h6k/24vkLgHWidRMLkA+/61zikBYeb+2yHj1civHy
xsDJemKEy3Xh1VX/WLzX9mu0idc7pkaQzNiPKvB+5OuMhADpO8nKuJSd9PEx5j7t
a+L+GAiacKSUE71joSVgQlOVHD/ZmJQSdaIi4veIioz3U0osI7LN6q0jWImAPaWS
NyqmQFppRpn10EGG9OgdkANRQOh14ZrH4svQ1EsQFyHzo8AY7tmHJD5mB8Gu2NxP
M6fMn+Kkf7AbVvxVXFHSoBgB9Kx3nPnFnXOPpNLgT43z6sRwbGsJZqNbmt0QPR7A
MzzGydWe/Lvgy84wzEHmOoEutr/8NqHEn2k3pHEVmfy/KTgZj/c6TXyZIDV+t5RM
WBxqbfS8G6d52T4QCrCMeLEuYzzMueHzetDm9GVSg0m12g7Z+cNes6xajDsB5Bqc
B5hY/SMD+RZ+KcIR6y/63H7/hWV7WOFZC5S+1CTmU4XP0W+U7MZQjJBxIbz+NPlr
pZLfTMVAAYOyTbLaY3TQOnPi0BIpJ3kJz4XGnkmPCOEWDQfj+pb9pgvSDhH7CkDw
jqO+SeGA6O4ed3ZG7riCgMFrBSfCaWDyC199zvJ7ziMm/xQ8qcxNoUZ8uWhUyJt4
d2iomlK7SQs9I1p/1SoBmgbuYEyBrxu6Z0l1uJyGos0fHmC81q0CyN4yZ/QOJ6+g
SiAvMIskZi2QjtHTRa0trATPy2WkTix8R/dHsA3KmEsFTEcjJ1jTeriV4a77W9jK
RdPreULHP8BatbOr7LdyQ5R5AumHNSzIHfe/u0phiJCUXzLx/www8qaWUPsWAxHt
xn65Lk7SWPuld0sOd4sI6aaN7tQllM4+Ktzt7M0V0Lw4J7GME/Aasq/3GeSpgwuA
NZEGJe7/JfjoZKIdOWD7LmlZbuYdZ0fpUvikf76Jgws891N+3y1oJSVIv3LXAUQp
EWOgTT48kOaXpKi7+o7YxTWIU16CIYNxmU+PmE5QLAuvc8PfE7rtawhAXoxh5tpE
BUj9uONnp2EXkM5PfyrOiVH/Mxsrt581Bq5haXM/n19NMhKAOjfjTHpTRKxyt44/
IDj5df0p4F277JI5zrTGg8oI4lKmmDBgvTkHc+qujrtULtK4N5tF3l1E9TDBPKop
yHbojSvaod5SDd/RNQdm5qR0yiIxP6mClquryJrCS9iW03oaVyW6Bl6uDNjL5ff4
oC/XeRfSw7EtE4tFQwbtsbF+ryoNvCCPvnDLWRObXDvWnrGpO84kaqJd/UE5AWm/
h0CyqSkumskis4w4HfMZ1Sctjh7M2/dNln5iKbNlLyCDB9q+EUt8K+HBMgtAMD2x
acbmTsvKdAnY4KPmgNEqvji9VGf3RRNbYxv5/BO9brfWzGtcLGFpnJrxcvbfqxgP
VoI6dtfKOqIDg1/TYQOwGCajuq4jjdKLFKuOR1bCpf5QOh60Sa4tw14iqSSTwJfJ
g93kB0A9VoJDybkNuddToza4ynYl87OftwX8Rz04SgaFsYcL25rXX9xzjREqqy+a
nlvn3f85KwC4FqOz13UGiw9FluUlYXyvUW/WXbdT21q1/4nyrChz/Ph7PmfY+o2B
iVVmGx9QM+FTyQXau1XHD7XHelMGYd850S58hibdRrpDpbPF0xtmsI+ssspPbRDG
kBbn64ZioCLzztYqww1iCzXFbKAQZS+wLIxJA+MSk2Q5VvbetNkE2hYJo/3rwrck
tAi/pl3JEHA2UcWkeLlj6/krtnXoB9RbpjVqAyx3Jyq4c+Qie03N1fId1yPGX74r
XE3mHoyp/E0qyr6lQV3qzcFiZ8737inXcWw3uohs22fGicGjG/HPo/nh/7XQKiFV
LEY+C616lZgJDYYIjk7bESPvui3FkBmEP8MoPV7cGJhjLO4wyGlVat9ogE0MZKDm
gU/rVDizel21GNZwWp0iBUVlcCrXU01CuVmKC5jBN1+tdHRMlmj0O0SyP1tplr+H
rCgtNODAbyCmY+dwx0t0KzsHFnba8oLSAmfXdBFMHESwnnW2iowUGYZXUV8/qhpL
gkMtK9Zv8limszaUnzC+0ZZdmFJJB1BrupQmUEqyI45GrFs4RnwFqBn/53AvGNtM
8UzVmOxcUSN7KWnU/4zWIRKYUOK3/aFdEF3isuP87kTQP6y+9uZAbAG+7fGJOz18
CQqlYn0QDQJomAJ9A12US7YiM1hc7HI9P7xQKdktc/kBuqx+jduNk9pFReX9hyOv
hf3kWygxC1BQWwoTqG9+XXPDxGFFtu0c+WyP9xbOZ5KNP8jfknwZeGTXaZJ7whNq
IR9F3LnvR0nJW2LqlrJGlFIo9wdpWVO4FSSGqQvMsRCSG1V2kNue+CW6Uv/fwL2n
gNKTjEMeBYeyzTgKN6Ud2UAOQFrszpVjXNnD+8iOCNujC+yewOKNQKwzRSHDD1jO
wAJPb0fe9q6WxKxCfCwZ/nWuCM9VSg+V0oaLscDCIvHhpAQ7U8s+etWOJ/xDzkZR
JdYXWDRkE9qBm46iixRSxLLdS33GsKzzrkZ9dfid9k5oWBxtAONgnVou1Y/ZPeKa
FHxjOv7R6x/3SWJ642R9qwjtWvl60luAscGl4OeHPwE/01kmYg5Ua99zQEf5960d
M7e7RnQAD/tylz5SI0B3yVUwb5+h/wSQQcaF4yCjC271tWAnyTJ7OA09fKl0tg9c
xmEwbOc8GfXh/K0fFxOKJZ5LclutTys3SgQb687EAlikMcerNCwjXA5F8fzpaEZa
pHExwbBpF3vtLB1i/jG4rzJJcbEN2dEnAIL2/ymfPG3qFOB9wZsfyIDR4OwPj8VM
2covHtfudO+6dMDkhGySsSguApc5saC0bwmfl2EZwZzRhyaOmcTklENMjvpkiRVU
e4F2A8VlQIA1HC930Gij5jH2seU2+QPF1XxE4lcadwdD3n6he4Vn4QpFT+j8ZEVp
XgEHaop6D0zE6PDWluYXGaPlaDYBONVxLG1WpRfRDztHN7zKZPxZxjBs7FQWzRbv
2ex1RvAvBBlplaJIv75D3Z/crlL8h5DKb09I2Nmu1YoAw+i/3Xnb76PyUdHOIXUV
PBn5VL8Vlqn4btG6K/0s0bZeamDwThZzPTFQ19C/lPi9LJ+ptQIPsgPRHUUT0x5f
02430wP7k7782bMCi06bJlgGpGY/8pC0YQ4GYaRAoa59GqBprjAUmwks+bmmTy4i
fyyumO6+9CavQPe1xONszUjW58PW3GoZ/3HPzIS568XHIgubhwguAJlYyTEUaOXf
/MS15tIPwJ1gs1KURz4O/cBogvDXJ1PxWA2Gi0BmDFFFteQMxfh5s3cFXw17rKmp
ejYdX1RNSm2mQA9n9Xgjc1S/uJZSdCxPb8TzSJ7L4cw6JAaQ2AVwBa0TXWk7NdsO
z+rxG8JRW+M37sxZTsBosqAkfqFlDBNVEIEjxWNpCQnoiBV0iydECuMn3CMwrkF/
zsXlbL20G8tldAq6J+FMNgVkWQgyVpRgOlFaC5IvXBUfqz9LF2hk5dYsWzEOTEIV
BasSkOO/ZGJzzO73b9FXNxzfua5eCR0LrW8zic7A22WHiohzdYShQXep+Ka5Enze
q8/jrfcllgkeBJt4+zprWebPVu0fmTaeIVfX3mZoTQLPyOnnpDz9Bl6jYe/sU+pW
Q6Hev8uAOEgkxG8rf1W8JDdds1PcPj4LrNi9MAiTHNSUfAj1hnNe5WIWa7mKp21Q
2FAs3GWkGKc398IeFS7LzGfYwCtvgXo31d722iDCWgo3UhKV2jDcIIJ181Ox9SmH
+wN+iuVQ7jwVCWA91nGY78hQ/EfQuATZaRLJNOmlB01RqqXg/HDfzqbyZZVNloFF
JDcpsNjjATXGKbQWHjWb1h1tCw3Mzu2xmgtzyz2wc86pPyzSy8Yo/205XXSiNVIb
eXhy0wfNBQB9c4LzbuA2jjyATKcBOnh7SqAgmTaC3HSReCYQZZS0Af/0p+haXLPh
K4p/Qh2EH7tOe9qcSNksngJeHddG7E+aI616YLXxYkp83WcnAVSaj75uiToJDbEC
ScpohQK+IcEXucwOJTuwD7DMf7nRj1/93sBM50J8U0siVnyvaA2qHobfovERtcUO
PC8aFWowYVp9/O5BnxnSTY2t5Hr4qY4jYhQoMe2UB7t9NMRLRDTDv7gn3ads3rnB
LSTs/6GdZOzQa1JuRwJhZM5i92WblsN0dqyIrUoz+Q1+0YPpJ9k64HUDMOZjrs/E
s87ASdOuTiEeTK6sIC8t07ls0SJ4X77qh2jmV31oK0K3FMDFCeXCUnMOi7jM52iQ
BL3D2ClsQ34gkfi0lRGv9l2TCT88wDhkloxo3Sx/aMGtz+LEnJg+xuMLCvebES8p
hHnGl+sH0r38bhF2UBElXkl8cGDPxyWdJGnl71gcihDNPNZHfKmzhmysYYaCWavW
E0EYEduQEwztXP3n2WC7TBHWZYKZSq/bRmjRQpxeApbLWk38gYL5Z9UziG0tKMmC
LakPQEdlz7wRFFMyftAlu7F5OpKJZeK31P+Lhr29jirwDNe8XqazlwNUq2z8Hk+Y
OuSgUnKe1J6RvX5k7H+F77j6aCgcX3WhXAYiw5cKex/cxcDGdaCAVY9tSq23/n7l
0XaVQ6MaCtTQIVcQHNEw1XGMqW8pREGgK0w/GeNNJiFTZtaEfCTMyTdKD7kWosGo
gnhkRqrPLL/vpg8o3LVNJd5BgbOmjfdZ15sbbqvT3muRr2+jgGefcu/XB0gE4lUU
2lTeudYg8EeUyAF5cg8eVoSmTkDutA1E2MG1Uf4iW55H2+X9QDvaBXJ9+GTOKPqR
xTw1p0pHEBuQBwRgSDv88QCkI4+JQFGU4jyJEOpDckg8WimpZ8Ow4KFHx12uPnEV
3C8YDc0wAzT5yiIA/NdnDru8qS3SO46+54Jk2xfAnfH2oUYUbU1RzMI4VSRvhXql
jFcd4mVgL0EG9XsCQEyyUpbOjbk7TQQJ0Xpq/GyRwDWHKZijI3yrnR+QWxjLkrJ4
o7IF41Q/srKF0e5LZ1gDe919Zb0NnAgePRwC72sQp8Tych+VzKjvAS2piWhWd2Z4
JuQPMvOln1PzFYGoB2fJbZFb8V5ocPFsJbZZsKyBtSOVsGvwbea7TPVjg9Zrix2R
9G5wBPmAY2rK3tmw94NhChyt+niybywNVv5d6e4nUpXOzl14JMsSPNx6gn60KJow
YO2z6nqUtWtxGl+wqHYH40Khv7s8L7Q4SMm8cM/ZJ1F6i261tcuYQwytNlD8rcaX
4+J/YxuyF21pnLyq2X1UA2SRxY+N3r1VhG9vpvoqqsMgijXVDmwdxVloGGP0jvOY
ulB7fiS+JF/WHcKl8eF6NdYQI21zNB2Sp/eU9ilKs1BmViZn5qObnpjugm5ai8BA
kmYI9j4nkMfIrJb3xz4T+BvkvdGzlSvu+hqIDQXTh2fkmVlL1pGGQIVHoMTRmGJQ
Uk8BOtCrUgEKZcQaXsTQGyyTAcetaHrrPqCKuEGJSLjx6+kfwnLTp9FffsmD8+ak
7WyxN6VJ16E8BB+rQKgkVJgeRj51LIuFGOaOzZeqaTU37pQsroaKCxT0wcsEPJkG
taboaJPoLIHt/yciY+YXfhAA6eNCQ47L5spt8FPJg7wVyISQiZZLODgzin3z7vzX
7pRmiF1itknx3VuhyXH3ah4bCyuE6K7wYI9ZQ38QOpnHTFOuKX//4hAURFiRDpBk
+I1N6Ea9Hw9tPpTYq66hTmsqkMT8adsi5y4uoL5ugRzhlJBXrEXPZQ5yQcwhL+/o
qSO8o0UI1fg2BpyKH1sIPxjtaLOWaSxGxLDaOfwE+czYNjjBwYh25svGTI8P2pF/
fjaNio4KcduOZIrPFh4qBEvwIpAG3pvnTYR2YV+HRLGS3qsyhSM9LYXYW91Avusz
vJfAeg2wzh/WBZU0RZyluREOpTBaBqyIawadEJEvm6OxnWieSbotDTCOoYJ6TGp1
UPgew9c/kwAyyBxSK0QfdinOzR0cwAvwtaYCX794GdOMIaYHRvES+de6BiWPxSXI
0axNSKJFrEibqOUSIn8ansjMfcMFiE3fUNZuU0zDT1jqQ0ZYBPmlAkSSqw7in2Ab
KCtRxmyvoA/sBcrcajDfzSDioyBi87VESPdxlh0hrTJKF9GlQDh9Ol0B1Ra3nwsJ
6wVDPcrXMW9PS94V6Xt+b/c6x7VaHpFO0iYmmp3wll7pcv5SFsxmHmRLLQ9wlAOn
wAsPRA0dCwo9cgeCTtLM+ubGQGVKpSEgIbz+VdOSEsNNSjtn964p7YfUhTmsT0pP
PpyEz9qTE5MCVtPhPwWt2SrsUWfcuT8aTaoC6H9iniE9MLKUWmzj/W8veRt7PklH
EvgYXTS5FIXK8Jp+XGWSZJLMj1c0fd5RBUeE4teFmzDnFe4PSr9XkfgRPsCw+orm
6QQvBCTtU3JtkqYSm3K6SulFrTOajwrmfPfEvCpn3APDaomD+JCkUUWL/ZqwA6Jb
CzLGc0hTsKuMUQQ5HYFgQYH3A6uPm323tqNr9aoFqYirip/2tFlzazGXy19qedBA
2EaFBXckFBKqA/t8eMRKTLAn8eC27EfaTkopl8pK9LapedbUzJ06fIz/yL2xzzpT
XZu+rNkAKQs35ySvl0Mn/JU4H5XiCGcC2m6hmROmAqMqAkYGAe/QJT5Q6m25MmWI
VPgV3zl+jsGoUBn8ZRFVf+F2Dl+NNNi/t4z1WwqzNCAZYDSi2CjfF+MKEj7c4TD+
ixO+sR+K/hmQGFfq2AGCwdRnZoWhxTxH7eit29Jd8eSDFqHGV2/cO1R9RM68Lb7u
snViGCvURx5brVAWCtxocyZdiEX026nfA6KxhLUfAc4Xi6gp224fUCJreDAizFm8
lpsIdJEf4ldy+J50Aekhtav34zyGwOWImpglgil5b6a3ZaJw030r4T3HQ1/67Q0s
JtvUpXJlR35jVnEfSMbBCNGRRLSBXOAbeT1ojYlBOemggt083tz1qWq2iK5BnX/3
w8EUsW5ZnW39mXs0wPxqjvaSFNFdhXQv/Y9As8lZtHylUjtT8WvPQyUvbfg5NIVB
wQgRWdnyW5ZtgNKQMe6UQQMxXTBs53S+Q74f7w4C3qTZFMpLH3tfltJRZ9Qzd57u
UyH/Ne1xAZTPAZ3DloavhQ1lw+4YHzkwZ5BeALbHdu2Bm60tPXa7wBmwBdTqvGYi
XYetWGS8bnqQgIyl2pLQ2aDpIP6Q6weBMNOppWfdXRDaRpjoX2lhGJOh34p7dg7u
TqCEJngyv2LFpeaePOjAR4xa44BeqrBwzIOH663LgaE+XplCSkoSX0fpPAx3wfZH
PitCMnovMioH0mGbM3E2otmKgRaV2e8iN5eQSGv0qyd09T5Dl9RLmlPoAPo2iIHP
TnoWQADDXcIYk8fFE9TYjE+2pfxJ5B56E0qI4i5MJxiZzAM2sYaYmZnBjmneibx+
0+38nI7ZJ8fZg64InFLjfCDuiiggQvAEJyxGK1KLKAhKxkAutEZKTJGr4DTEjYRG
0TQpyzfQAh3DnJ7GZ6FzU1B0GHcVG82cffOcCKeLojOnT86asB86/iwmEWgamSE3
hu1O5qOEpJdGqVZoKQDqbth4WW4CsWdBgPqHnZS8o73YNtn6HuAoOLO557mYJBm1
ETi4S7niRh+27R/ynwPus+ODpe+7t5aqAJkInmsk6HXd9EVbQ4IhlKvrN5efS0UY
iEcISc9qKSsulB/U1WwOsdvfBuAi3plMA0nBeJR3YOjqrhbRiWgZjrGkdGysDNcR
LPkudFR9MsMIsaQoKESxpXXTbu0RCnQ89lVEvDy+o0A35ARuCxGbJU3cCpWNx9jq
SPrvmxQg2rrE8G7qOWD15uE9gi8xFjLS850OggEOqm+0nLXl08DaoC2kz4QC5Mke
Xh9fXEoysU3p3h6BcHYsqftVwMLnlZO8gp9BWpweqnNqzkusqa5revI61adtNhYg
Rfk+BdAMsoBdqGShDUiMbJOMYrgAzm+O8+GGcBInR6CmsEBMPykWVQi5ZuTAArI1
+IDvOPhwFmb1tVWMtC1aAPY+gX/KUENRfM2pRyWaHzwFPcmtdakYc6AUc7A0oX5M
GUMVkjnAWp4LvHR8CQa8ttGeUl1ukWDMXyfXBuR97+/2e+fbUb6UJOIsKeVkpIhL
cwF0IO0Oetw7WnUwt0GeG7pRxAcD3VyYZS5V3KIwq0cV1ohEDtYhuaQC+wmmn2pJ
kRaRpwcdB+tq0EUYlnmiNQB1CgESKFjofcw9i4Nl3A6QOhPPZ4PJjuhieviKfeKb
gSW3pj84Ah3mqi62blk7WraNe0HkcmWDit3/x0pbdQ6+3o3HULXsoNjbRgqGIpP0
Htr7Ag/sOK229CHyY13Zqs1u4ts4qaoPL+2xnAK+DmBBuSVKj+zPdjCBMf2Q3feJ
VrlSDg9ckH8NqgaBnfJFNv/lYKsgpvYFSypQGYVHAelgqe+zXAVbNr02DFI/+h2D
tCQbxnUNwz9rcPgzmlm0KkDo61yQQae6H5vd9XOs9cjalw7s+HmPF4CdrOKVnps/
jXYIkZLteM9b/lrvTTbxwcsgDAdAXzev6Hxo6KWfX6yG1FQeQV/pJyrRO7/W4Mcp
RHbfxR1/BltV9su9PES0wf0StQB6qT8JgJiAuds+26Q2Vyww2cAZUbe5RL7Vgh1o
9jceZ3wGm7L1HqglrWFwOffisr7MgZPGRdrwJ7qjFvFCmBVDNzJkkvXoyapE/54A
ikh/qaAhw+w+4W5OXOnGhJ0tWLzJ/oZaCaOI18yvdXTgkDDkraOtOG8D3LUZP+XK
H5Q870OSnhYglBpXXpGiZbgGsleRfx1220aurWsgblVJOz0U6O+esBUSqAb4yq8T
E22tyaefTExy26CacLYikABi1DGbZ0vHxCX2Qvl0EsTiiY2HdREZK3o1oNbsCMHJ
qiljushlDCSnygpzqUhWWSU+Sw0Clb+xKawRg5L4Uj+AMj1R7UBZo2dhG/yxDePA
x2X0MDJPjjrgUeHGFroow6TcG71aFdUbb4O0z/vihzyE+UBaK9pRC8zeF8pWrgZo
oUNnpuvRQzyNrIfMDhIy8mwUALu4w8jLWQY6GUygWlbzD5QK/tTYwYQatoxchBp7
rvM4KHr8zTjoRjk+b3FVsqp7/gn+LEX+QyAeDoBCJ+MN0BtBWGcPYLbZcOvSlEQB
neEUA9DNbzFFV9+GUiCf/RO+DBysVExM3eDphVmIb0GBuexRyJ7T5yukpU0MKoHK
NLXXBBKyUw78TbFh/NbnrtOFIqo/Wai6QdQ3fld+n3mVM/y7SjjJSL9LPsUUrQEp
6d/iIoL3yJEKzvhT6EI/uE4BaO7P29XQI/xpj27fmnbqE1v4IOznRqHnTDTdDotu
Ai2KOX6/IF7zV8JpOvAWE+LVd9qthludzI8Ei6GY0uRY0WWgBbNm0bsW0uhKvST+
UH5U1bjVjjkM5oDAq/a5x4/pIv0MEo9lSzErV9BKoV4BPBmYvNEf0h414DxFe+RV
QX4M4MoJWCRPPYrsz8zodJS4hvg7+BvwN8yHG+T84l+0uQk8D7TWvyPt+eA6HpkU
Pki+xXGO/8rKuqQsTXqrvzZ8md3oX4h+KEjc4M+wWsR/y2hRrSwAwYnUQUO9i0u6
N6926zVCsy/jSnEHQWv3mTuKyvHdDWap9XDXmN9X3wIGEqOPz8WaxELDU780f6lq
bIuC8HQtfghjnOk2znqpeTP+YCjE6MRXHYM/S2X77pRdqvemjpz7J/qJ2gQ+8GJV
AbbzwWdbfRFP/WVdqD6fxUYa02W5ivTwZ/muDO5gOrvMJ+0lT1KAnsXJ8tgCC+hA
nu6vT5D8YdU2XhoAnHgw9ZKTQek9yaPNTUjMg5hkKmN+1bdPvNwgwJO19W231D8E
80ikoyL2QNMh4jhXzpjyXGU4SMmadEMvDqqzdlW4i68gdFbFi+6BreQf9n2HTG/B
ohWS7gyD5t62bE4hhYfJCOVoSCi0N16Lf6eFPew43aWLct69JNxVETK8Z0KiM2+D
1gvRszCA7fxt9UfLjnqw0GE4RMqcwFn4nnqsTVCs+rHj94duupQlPUaygUpJ757j
IuiUkTc0RniQp7YfqcbOjyH7bT1wA+4olpKpl53zjHV72pZm9qp/Og6S+e9TfLq7
Ino3m4MU0E3jctYH7Kj09Vfvqq/w1veo0yg+y5sV/QyTHCUumfuS1s19DdavvSpA
p9RWJvBqiwYhfweXuJTNhRmNnngVy3lnZmti2b7arS4qlE4cC69qLYptbBm3iiLr
WaNLEBZe2UpW/+OLIo2t5vT42wwJ3Bn7Wqc7TdDNkuZ8u0CpI7gFHCYUwhWF/RM+
orS831jun884RSuEdYvjvq+iJPQuIm8pe071i4Y2Bnbr0Uz1KYjeaCbRUTibVzRt
l68uHrvkjmT4wKt9wEqugr+TUFln7JWL6ga3hhxpw/FaBZ3SO6O7Rsg/g+DLk/l/
0NVYUrEtiftxm5gOtOTTZxVbwMQyhDNRpWTi85S2dyN7tludbkJV3Cmumz9rc1KH
zPPMDoNB5FpWeU07BbshGE58Dt6Q5LgC+RQDlcDcpDSWLcG4Yi4lw7mmlbVJeUGR
Iq6VwBa1cwTpwEcD1NMN7z5TRXNKWsswqFUyJ5Ms8LPZgoJYq6N2zu3AoLihoP8m
RxfSInkcy+5xWub5ceu5B7diQ1glEXzyKei4RvxlxWx8IaIGbzoWKm71CYQSsLOQ
hZxLurLTnCgVg0XkOqq7jh9rKAo2bzyiyvNEm7YLkQxoHeB0at7dWgvFNYjhLC2t
u3L7//oGqdNlpZ2ujUkVGor/VP+N50Of2z8QQSFRLjCJy6Ry07vnHzxsIjBIiTKy
e8Be8PW0NKVJ1bYbpUsQ0n8TxAs8X/a+XZfbdJRwHfSqDFSYL4dDMIHXfJZFaLxv
Ypfla7aGXyo4uifp7o6rgNka5FrojQDbNnAzNKiaf1xQZ8toQ7M87AZ/HAymJefV
vSnZRarsGVxbuxPcE9vLBH2O7lCBprsbMMMmrtqbSRHlMdrJReD+r1VI+cCkOB+L
C98SEjdEC6FmdXaJvsrgC8es7kUSTgTV13IoPxV9E6aPWJ0aQqQYvE40Yj0IMWsP
NPYsSpfWz4pTwL38apJgSLx+phHNb+Oqc7iX6IPQKqiFnhrlzr49m4aAZgRWjb6U
SoE/nO7FdfGFxhuEvwYiJKR9xtliR/bucLbehhHUTpuSKVhAOu3zyNUw66NE4meE
QrZpcRwIN0hjO/Ps8ZOD8TNTgKrNrS0YD5JjqnAtxRryz//kZ6/FOBJ0QcFDbFvt
1o5Mi68/MPz71RCcNHP+ZBLUnh7h1U84oo9SAGzNtbHxbvvdZNP4g7p9hkgg+fZx
VEYdioQsdkGmHztmiMwmobIz9cbXFnVftvGx7agmv2j6ZnirqSvzDgE+DWqVp/CI
IldxMJKXW7j+IuSn65P3he4MJ/NZFfy3PpSDH+0svt7+EQ72AVjHxNndWhpN/oRj
ySHaqZhp69xA3bkP4430RxgWM0lyKSMaIx9BDVc20ZSqWNGHbi1YZyND6pMxB2YP
xFaqUpUiezUyRoZnL8XZ5u+igNgDsUO3n77L8vR8Qwavvb2e2HTm5ksh931WFz+U
hHZqJ/FmDIzrjCOaMLTC+O19EuFYLxaJ5Z0LWn0el2q4g5eChAwzfwSD6r1sdT5u
AcVcw3o6758LqZhPm8hSOIRJ6abfG1PscqB3e58amUubk35fD2iZWZmTxuFyrBsh
hdNa4YfnyEKKCsRBJ3xvTWY8XSkPY7IBllc+bIco9Cs8E+lmv0hfRqtTzDqy2t6y
CSMUjDVzLNwm6CYCvBBGkvkKDft0WzpNujcGy7X53eFb1tbFb7NNpTvqlEKQRukY
OTq6HawfvN9smRyBwx1/Dimu+moiVSdDXF/G0ZFddXl9vajVAam9sOpZtCVC7RF6
YG8+uDT/n13amucF43gNE+jvaR7aBpj9eHu2kHoCWhUvF+FhVkTUXwjgH4VkmENp
qQtB8Rh4qTbWaDHB9S4KjwjgOek0qdRMPKcBPde2gWr9u+GxxXAdN0V4g+R3gKhi
0yIgw3e2ZR1HLDDt12r0hteFF+Y/FE0vDa5xf1Vbn79vWxhOsXpcVFoXubTlXXjJ
/OFT+0YKjZ4I7v151Q4IgZAmKxtSvtNoQZLu+qVbTfCS1d0jhiEfJDbAfb07HyyP
fwRJ9Sfyf2RE+kz/w8wIBEsMEH5c35EyRN0hwSOMPz2JodIIVG20U9a6z3xFODpi
64xdjqnMGLBlT4kre0LtP2U2+rzYqBRonfNvVVtyUPaUnJzF1NZJDgasiWYjhoF9
C7lYoqCzB8V77pXXDNTnAduYVMmCHOahM68Py+5QlD6vnKV5t0yhjnwu2J1i/DGO
Mc2Y2zc7NyDmTjU5tU00Awd533Zc+2C1N30xeFRcUQlEaNW5Ih4hc332/nzTcE8C
Ad/mdk3aTdEV2UPhdYae0szvjbsNl9wjXRE05ltD+++jMrj8mglRKIaiFThrOnVq
sknGdPwkCOcSKNDDwXzTFcw/w1QP9pvQ+1lh1FTVcPhg4/lvKopwhi/ldbyXetfJ
cuKyh9bE6habSE1jc1df2ncPR+pcrtu+8DbyPCExVgh2HUG9UqMwnfizzoYQqy9z
3jv1TP7vzlMDa2ooyTq3QIdNv+KOlt0SQ6ucJEltg0O/tx3upfM+6vWOcnXVpqTx
IIAEPXuj6/S6bARU46m53fj4u5k0GjJ29WR4aodofgdkyf7hY/7SXta36Wp9V7CB
dCcYKtKo128i1INWaWJhz3QFdD+f9ZkylPCKGczd0NrYHVZzrcyHQyAgQVM48pCD
ptvKSfqZKwdqAUYBqvJ/bxuEl6jtmqzjYVqkxq8/X31nqYfkHnTViyaPylgmPv2y
2pMyBAkh6sx8Pb7ATao+p3fdDyt/dXROb88aJoW+8tTffT8VeptvgHAg4nVEqdJQ
WTIIcJnytTRQnNasFskCZf7Bp/Q41NdAfCD75D7rh0D+cvSiw99nqKqnNYk8yDnl
e185ih7VNlBIba7SNBWGauSDFkN9A3mB2qmnPcZL+kH4O6ayV4jSHPSwWu07H2wD
lyfM/eWIUZr6fwkr/zn+Ngfi49nB9KUK6flgZZoHYhKGXHpAOlJPyKFFmaAtUTlp
f8eWb83Kf6yJsxW5pNYMZ6aeslFJ8NMeyQACfmtu4Jn9dfR4wBBJDPWS5TDpgrhf
RlTtpW+k44/7gUcpeq+T5cYHSnous0cOp74+6T5+RcP2Mm/mzvO2rV8Kk2oi4gJM
Y8JfQLhosQhQ8WFTaaWxUBfespQGzQj0o80AqMy1k5ddISREp8fC4LrfDVrWAu9B
BhDLCRXCzTWcBij+Rg1urCI74xZUEfw/lWS3F7kuidhXeVORNf39KYdxaeOAWDHK
kLYWT8I3SMyznC2amKEGMJHvcIWsIseS4TW9bGuyrXdA/GzWonDDaq1voYUvkc/b
IXaIXbMfH4ZShJNL+WV510U6W3uSSSki8aYQiMj+Rid/6SMsq+pwvrP/RTGY/8NN
P2tZXh+qi+3NjXiJ56g8xLgKF6eEvdH8+s3/OpyG4ccV0PI55ahL/48HGaNuxskt
uiDyaDgN8P78ldPNUiO96CJH7qwloAmviYEtclJZhSMM3qIMv+ONU8ZIhujxwu/o
79nNU3O8yb3/v3WlH0iP1iODZ9eNUiAyEQJ9zuvS75kyIpfVM8jJf/s2tunCrZof
qbHlImYgHke8A1eXnx3MkAhhBre1/MOuxDGEmk7LGJDuIMAOaZu7xjGlUi0I7mRR
u1XoVBcuHdMBEDsgAMOpieRL2JAvngm0u+C/wiP9US4zyfRTjYS5liWaAJ1fwWYd
jlIkL9h56fP8MD80i6r1IqgJrX90GktylZeHvdoUZKrILipgXVDMmiV2FiyIeh/C
rmOf91HzIe+gfAgQxgkv48XvdzqiH4DNKgkm/Ub8ZCDmG+u+SbCTXkYxu7lH4IQC
dpoWdRC6kMsBxLleMuiIw3goe6PYhmBmroDEoszy9dLmsJbZiv5T/n8i5mv9Ure4
nHAZIDSAblSyiyymmYx3ZDHZHQ20rbRySWywAbVGoqJobpiPMxWcWTDfDdLWOPV8
EW4eQwF5HkpFZ84c3EiMqSGxScY1rpJhdArwnviFd24w6I+5mh/Up3igv3CHPylb
xsE2sUkEjoYwjn44/u5xWlmnz3tj24dg2SUeIB82aDBiCW6UfRePUKpgb+h7tyO+
q/Umb1GdmPE85hBZFi3TnxoIRJusy91fYFW3AK5ZHjgmQ4lPbzBB0prrxEeO9AHA
fZ+yjo32r4ljyoDgWERIY1O87xSK/Vfr2EwLK2DypX6RqG3VW57dh/+Ijc7IL3gx
unlgeijZgIaVyoud0SQB90SQWeW614AGOOnlWd50eXheUsQbyS+28h6gSpXOkrpW
ITAqYo65xigDjgKOT9BHazjFhlJutYHFMQekzdtf6iW6gNkwc/w1YdtsSiL40O7V
5ndBczXVnHwCjVlz7kiIxTs7Brx1mJkES99JPbONWcq/RcsssO6L5A8GY1vxUXN1
dugtU+Eh5KJeIW3bdsUWzcwFBsiu/AQO5ughfBLjVwFDNtJgqwGlF15dAQF3+yCV
YTB7pjLi3ZkQ6h/PgsYxb12dyJFeZ1eRh64BzgvIuh930lG7eWaa08ndELbXI6w5
ElCWn8YCnAKjgCzCseVWdnmndo/IJvvbDlfZxrijsozFvtXpRJzMAwmxHNh2L+PM
0uYYWuDjiyxtYQY5TxM0UEt5oo2FKfWOeXp9/Ezgf1SLtOUxIPqZMdX15GnA1q7H
LTHy5+zqt4QmwMn31I9uhZs7ZFbATcvaOpXyNvdMaR9I+fudigvrzQVhxgVqjHIN
VxcAmrSC8LAmXlUjCn9GysL3SfVOvyAnqMO0Gyk76TiE6CQLMQCf0rt1rzm06BAN
v+jdoSaUZ2Kb/aMSh+gQ0thw7k8dOYNCwmCsYujfUFTf8Rj9Y5Vyyd3y4PxRlTdo
Q2aP7nl7Z38Fadbsqvl6xC/KJdZYv7Ia8EJ+XgWWFlK0UArdf0dZVYqhJbHYLNJ0
OC+Zef1ug4smgxG39lhigvq/oIhk9Yg6xky1Rwwgg0n3cAdgwafgJJ+GnTn6rt8i
HoRstjkAh9NMMiz9aEPoBv1XdsVWBBXM5Wst8cwLQjfD7JEcIQzVOUdJCRvrDnXs
r+dPYqFWpnEV/XjTFWFMKM3rezGSwgP6LIFBBDVK2dx7dnMo972pJzuGRVJlVlPC
JZlhqdUTDfD9ZtIIR76x0L5s5vAKH36163p+UkrCoq/KWF/g64k0AcT+Xk0HItRR
TAeDEQ/Vn2VpJ1OHK656Cqo/8N7ap7les7DIHZGqL3YX9OoLFnOdkmK0+MHxgzz+
HPTWC7udUfm8nXEXEx5+rr4RRvPYBTkvf3PZ3MrLwNOYzgC9g7xQxmdl1rbQ72hV
pLG9xIa3sc64BpBFZP+op2vdmKNlxEnRJ5fgFM6U4SfThuuwWKrjCxQAneyiY9pH
/rCSLNMgfjp61liSZRfAaqpvTCsxLT9BuHZJYW2YJ+9z1SaFCwXNS3czN95ZwVz5
W8M/zp6dPjQmLGo4+yGUJc3EbQjukoWE1NLFGpUZTisA1k8SEnf4p0xrSsiJTCOq
8YZB9IcpBQt7ZJ0bxjRgYjylbbyBaAtSkNIp2piqHKt816/C7GFCiOV8VrQmh3Ok
6yTwBVs1Xi8WdjPAnZxXogtpI8r32+e/bCIZYreeRkm+3ku9T+bXeNxS0+42iNGg
nWnnTe4iOJY0/3gAoMp+cSfhkQiSwXgHX1C1j5jCsSANkXquKZ2QUn8PpebY0NNK
HfRbRXHue9OF0geoAxoorMrr7U1RM8vFpmjuEY8rHxNDziHAdpqM1NOgkgQlflSD
U+fLffJXDL2UkAmooNaF/z5iZqdZnhjqTUcAeFvufJH5P69gdLav6zK4jL9VAjC0
J51phQEuCo2DrtqoPnSfQyDGjshBfFkQI4WDJspEkg0D6axn8+1xiHSn0TC22JEP
qv8Qxws2Re1bvfw3VfNgui2GOGP78zOktpEcPVGr7seiKzMCWGu05COCYC3ryeF+
9Db1Y5hk83q73KNhV6PviN6f+4dTg4fD7xBFBSbCqcq4HcmYc6RYyxPRbNS5dA95
N6UXY7Sh3gbRBJGRZIFJtPQt+XZLRudohS+34S+fezjtGeviMoWGcOdbMqLgRr4D
+Uv4IFNS64uY8X9Ew+bRvcy8UxyyZizXWycfz9w/cjHZeXERyvsxpLpl4san4kfp
5MlluXKo2vvEG0lu0DHMjrUxKCTIWNJFy8CMM+/MDV9P+T+F9NSPTmUcMYz67m4C
rUCVsIzSzneF2v/s5FxfH42FDq7o2qlWiXJ/N9b7+6Tlv/n4XshHRUAJNM3UX6J4
VU7W2gKECGVVfBf4LuyPNWhTcV35mqelg7vuyHuJ1ehFuwzKIuEu5qKn35YobYST
p8jY7i0YDTAa/p3Bktxmtv821+b/kYBEwevUU5YZjtb4+kz8rF6CkwPmmq93mSCz
NIOXgyNbrwll2kHfikeLF2T1bsXt9ZJnvCg0E+V//b+inBpn5U1e/w6MBJ4qIbth
/j0TWqmi8PN8klAAvJd4Lo2UI9AuOtpElm/3Ixf39kViubctq5vCWZ+iczuZldLw
JlCai17eJ9Fv908SsD2LlecJNGlGVIptpJ+Wyhwl7H7V7Dok1sgesSg+8K5h+xKE
6w+yQF3YVMsutlhw7lnyXKqd/93e46i3hDVDk60mjCu5ui2KnnpP3iIPlYwqYAEc
1KbCzO32kqwGGMuhmh1iuYi7RNvW35L1j0LZL/flIlTBHrc3gMWBw7qDWqbMyVSs
I4XjsdJ9YvJsyq3NENpzhhXSLeDBHhDHmfhMUaSssv2SiF2J9yzpALkvEsZ1Bfpo
FuC4QdnQDKYncCJfwhSefdLdQQmo3aWOyzKme+dFP6CNBZaP6Jo5Ojo87i6yIzdQ
cuLg634ICP//0dS80KqDB1CqysNlolbYZrUyCV9NBexl2qCVQaThjZO7hrsENRM1
23GRy1FOnyXaX4Vat0Q6I+CGCUFsEctorDHdJS32GJX2+LtVVMLxu2ZgiG684/aQ
9mQsikIPuH067fRy0uFRn5pcvyTeoCN8l81sEGlyF7CLoMy8tuWGlkEOZ3E9WOB0
7kqJBTW6pR0bvSXnCfKjEr7x1sFcJz90Fdlr+HJJDhnUQVcoBnRc52XeONIW7Sva
M8SWLkefmdw0nkWAHB9y0ZdnDcyE5QN81l6SI34jR/WUY99XP8YlzwWZKOaxEUDX
R0aZ/M/r0pOxInWYd5wyHSdJD0P5d9qp/2YECTZDkBOYWPz3er5AGKFi4Tx4uX/J
ME00Im+lWQMuTFaAfmi5+g7/B0ZryTNIpZtlBi0v3ORqcu7OmsTHQ6fM3rU+8oCy
dAyFbtjYiFasSirL2gH69cZqIAPCuu9ZcYTT3wC2idCf09RkfUNyifggZDe86xS9
crIunx3KE7p8d/jBOBJAT076QDsni7XrXUc5A4lt9iySMavgdUElNCtEstXRL8qt
21BUKCRTNiWT/UbBURu2woqR1MrZ7yaUF9NCMt+RbcFdvpxW2Bdci9hmdmIiGs6L
DnpEBQhW+psQ2nZjFr+F9poiNFhLcuXXscICvseKK2ldlEZwq8fUfeYVSTClN9qQ
ovayYJq4q4eYAGkPlVyvyztZTU6dg6/k5TZucx6IyTw4eHFnGay8ta7+chhCpdOM
SS7shVGQON+hAvHmq4jP/VcNs2QDe6S09ubiA5iWmPpVN2DraquooETGJKoXnLMQ
fX8A14NmJx99sUUAUYoeKGTsCN/5ob+9I7UNWTYgX/6VX/a8Lk4OuCf/Q7Ctcb4i
L5xwruabSgTm3O/HI5441mIzWiftSs7cwCvLGileFkI97G4A6klGk0dcxN2NrlWQ
JheinOkAKujAA2x+O2ZsQs05X+VihyIH5v3eYqzVu9pFpKGfEwaBNUe/BEfjKWWy
IHZUxydJbFxLMqHLShn1CtfIaxX9FBo/5H20K538Sh+1mJCUDfyrdhGOMRG3BDmG
W7VfecXEgj7CLNX0LYQseKEjVHZn2zHR0xzaIZ6kjG279Cl8ea+r31g7qpWj0at5
63OEfoRcYiyBLKKAIt7uNIsN9adssGm0hKjVDdc8XvWS7uMCtOK0+Im6dFPr6fzz
G9/OHk3GacftJVvd6wQuItHEfCsHtOIadjrqpBVWzO3cZDvsXJFxv53OO12U0sVH
i4nN1HSVf4uv029d28n8G56KhUDJX0HHZ3QKsl0vbF1s5dkx7fYFkO3Zm9a4XG4D
VKOyhOB/kWuFVnbpwHAd8hbGTrm/fhjJutBn6DgJeoCuY22ZKjH6XVIGWpqSCgeU
bYonVftrF4/hADx9vAh3tLe3DdGlrUaQQvFrtpr9iB9y1fU0uCv0+aNWk4w2OYvq
7HrTxuuA6E0dWqo5WUrKF466FaqzjqLLg7IMdkyMlSIf7vlpcOm5tdFi2D7XB9CP
HuKrd7O7cp8HU5zgY75zmUUO/5UvUnne2UblQ6Hr5KEQNBekVbpiZETBWrAVXQpa
JKEY8f7XDRnfJxcmXUsmDop+TfQqgRFJdQEmC4epIYaZ8+8D3swNvB+257Gw1wqE
NyXQ33cl2VntxW6HaPWFuncbUiHDOkcYTbJ9m2EW84KTZ2SIA739hBtpoYf2e0Wq
qqoOw23T7IMJXrAKyrME/rR2vpqHRFGsVh0c27BG5ZHC9gVncYX2T2UutYtwZcn2
/eounCyFlbJNxGM97MHgof45liZJQ8Q3x765lMJhHkd727tT9Ez4PiLGXypwoPdW
u6rkxv5LjSOzWWNG5DHFMvJ/Zbtd94FHxJKWRcezaojpWgJLpXYmk10LTLTh5zKH
Be1nWAXf2CoVZUK+146EGDvDqD4wuwaHi+xpFjxrAoc+FCaJtUaEI+LqLawrhb+X
7Gg+zNrk/xgM/V/mwoZ5mGdKeD7LIftfRWueCnkhwHddkuhjtep7+OL7SnWw2Q8s
46KIUJhCiObw6dv35GADVBALeD53VYo2XoLCIsrLETsWahCqmEl78qvZhJm3ivvN
1aSBXhuDoJpM0haUv7ZFaqHR1QvUjtZgyi8nZtfJ2SGuRufZveadMQT8SjDp9pdz
oMdsUb1rPaC/FsJ2BYhkH7ZO4qsnY5WwQy4VYcxkr70FUs8ekwG4KrSDcG5DuDbq
hCGSXA7mypPCDxDLcNTDF3W/vwghvU89j3QPGnLPGBFkcZOXTgqICA0Uqicrjiw6
pmrFHCBrnO7cEUlFH6SgIgoX1XKskmjfuqHLm1OGoCbX2UiRhM43h/IdDRY86mXD
Ud/F3bIqeaWq8FSKKy7HDmtYoGWta81qmAupM3Da0FaCaov9tvWYqMIXXlVBoAZr
rE9SHuqncSwzvfc7Q6GlIIbA817QMTPB4U2IRzPOxZ0CCNWklvwHfUYqD4FrPl83
B5AD8YthUGbapgXJswnZvC8rmh48NSErJdPnqZqPUbTE+LcqZRbjZxF/rk5ADMjR
LSrWZtBivqNtimZERDfTjE8p0BlQPAfhXRNPaVzTvZJNnbl9if1sRBS1U6NOpfXj
0PioS8DjJcfldBSWm7oc8TPIm8pvUyUA2+q4lkpfXZcjpWnUO/P7+aMmZmTL4bKg
RFI9HyecWDYk2fL3bOslSuv9Z4Ek378Ea9pMX71fYc+nszQsKzY3DpbAk3OBoukU
+CKlk/CJYCFUEcw6+d7BvKF3nSfDUCV+RR6yPTO8G33Yf5DC37LqehYkWKtjSGSz
sVPAVJMXNj7bPiXfzVGrcCzY6cf2RZo3D58iRMEkvMNHEdoTzofK8YdBhr7/Zytl
PW7imWgfKZdddN3AmRbi3nYl4dJRefDLwSHekDnz4otOW9WqGOgIjhOZO9zCBLOG
DVZb1CHCT91i7D7o/YFZ1pfLMwpBnfELkYH4hNInN013PbfRJfnCg+v5oxfTHM1O
awJ8yR1uzh3wnAx+EKPxLe7vDhy3srz25awcbEq4UCyDK4jM0jJ3NDyR55vLndZR
fgppBEbYsdI9uYW4G1R7kqJRt1fJjqm7mf0Xeg6Dd/6jvjZmn7nirBqBkxnarcCu
5Jx/nW2BC9RDQ5L6lHGSjo9QNUzQYifyRMBRLqQ3NomqV/j1W8+41wBx9NsDb9WB
MYApH5J9iEpvfA5c8qEZi2wexlZ+JHz4XTogL2+ImYLyWsbeDLeQ5y1ewPMMdTHV
ICGWQic4p7xrXev/9v2DkEUfDfaCbLCbeLtw0N6XZgvgrolhukYQFps3HlZdX/TI
t4giyhvKUjaFvY/eAKAlKaa63RqOtB29ot608xjvWS0zXo+nZaJQF1BDs/ew2ftG
BZrsC2SsU+TD3eqbvOQKP5ipkQH/4hOhcFNmUonn8U7JVibCu1StOS1MZHGQIpcb
IErBY2Sr2so7wX2hgEIXXiXmgiLzt8BPk9GBq3KjV3iiIZDOkT4z91XqO5PwomeZ
lIqMim2qVTLQ5MWowVHFKeEevpMGqqAwxFELSX7h/53GJp20CxBqAE/XVv8Wff31
bYDvQBEZSA7N0g9LLOxLBlQU95YBssjSHsPCJSBekIegrV4DBomoErKbEQ5ZAmyF
IJB8K+X12hXdWWZTKswIhQmj6XCdqs33Y2ZfezrXpXwVnKkCf1nqJ+pOo3kcnSWy
35GGbhGRlNAx/80uLDMAZYVhNue90g839gILfMEef80yfmVmtc7XsgEP+GI00jyv
IbfTAlA5E/zSOW2za2HPXeY1iXCh9DAz2FEXzKo2GXK0fiGKS8MioxtRci33EwcC
VzD1oUepJBRdi5MmE7X38w8JH2JMG9TEviEbUA+edEHpRmWALLbKXssCUmmGq/42
ABrU5zJ6d3tAi6hVcC9jVx7OBsvIvde5dmMYwElBJ/LDGjnOM48JUuIoQ2n+8Mn1
AQdev6UF8b3RG36DE59B7k+juipuJJk6hZbcu2G1bTMVwv1rHJhx1JNIp3WAi3M8
p7ExibKPRKWP9c9H3XCDu5cj5wNkF4ttLGp5FV7YjSi32SpQ0jnRF25p/dfp+QL1
n8HDhA7h9mYbAFg2DkVlxxueTQxOVjiUyE3Jg+tJs7NC8CxLqXmBG88AqQz0v/Uo
fxODveR9L9mwB7pkkftM0zbMvwnZ0AQTmprL3XxyObOUmoDOam85ltGeT24Q7p+v
18p7IUtieW0UkloV0MZF5I0aOnAVyzZUXK9rDr2BArXEB2X5fdKKZEHfbwipZ4Pf
zY0XyPrJwxlTlSGgv858bV9pn5ePTHWyucME8UL20Tj4MMQdWdV0PotX2zC3YEoh
H8JxbYDti3BN7voncq/aVTdZe8WkBb8fWkdoL2k6ZILj5EP362fhzfAsaN8XbdTF
83wH3YuReLuY0bzc9tUxN8gIkz2HG13EZqzeG+6l7Dw+uvVzH4DulOJWRdEP81jM
dOcOZd0vk5rtl2xbl8tNnGn0uRo9imi3ZohJvJmRqmdzI4/iKY2iztvFboKJFJOj
/g0wVHRZhxjt898h1Mv7YGsiwUeS1eWHMJsDzevZ29ePU0Akp8stULC3se90nNNe
VJ9YdoUQ3s5fxlxgFemGFIOZ5SwGHaEY+hqC5qGDHfuXJd7Jzm4fmN1XViurTWjo
hxLHv1Pz1ANbiybFxYyYHkbmiCLCnnJvQ2HWekegpgBYG6ROyuN9JK7Ftm/iOCOi
2VH/8rdSbkhh0t6NlqdVJ/45ZgJ+GR2nsrkMnO+2vXHDS8+yC6s5rd/I+rXJZGgP
hE2nRG7/oJC4yHKo4IAhoUNgX9VIDerworiiLQW/7iI2mi3gANZMTDdTB2c/i9Xl
q7CkuZMIhZ+7QMxCPreFX+BuUGMocC+qGhigGl120B9cTeJxUDyoN6NgWzhzJhLP
e5QZf2KcGfiiwtQGh4ks3JUlCNVD1n5qZaJDyuosilgIZXBz5omgn/euaScpYnww
9CvYa37bbWM64cqcOXT2aNS4HmRr3lMyOoegMxZiPySt7nqvFLRwSZ1/lED2uQmK
V/evR5ZIqALgjXOnWZJl1z7KTbt1TNf7qtqkBrsyI6k53M7b3yeSn+P8dw/HGjAt
Uix+bUOekLBbv7pthcJ+0u7FCmoVmTvNk/Y3/LQGmvE00GZ86vX+EZ7JPYLXBeB3
5sm6i2IAjfpx/I+h1whyAil8LdGCTf1yKGN9cTKWj5kAej65SnE6yzRpaKNPBRwD
q72AdwXagOtM8GosE71BvvdZY66FHB05OdHJ5zjF4fLvTO2WBi6micW1JYa7AIcu
PDGttz78WvF/lCuGDsSENv/vZP6AgblMXLFCh49v3Djx0++lQ6Fm8FXfonJ7sSNP
zcvGsopJgFHUsdo3Nv6WN/d6v1EhJNSgFImZzTOYA6ktxucROV6y4EZ/asyFiO69
RgXEduZb+IDLir2KL8E1z2o6uWpGTWlavk8p+Ch6sXFTRkBL8ubH83dp4Is8/1t1
SlmbLcYJ5kGpHgPfapywVUAIVhC/ilGkzW+kdi2UJO75k8ma4Q1t17tszDbIMDjK
4u8hODfAHGgcHnWhiIV+6uEQI96UJVLYr61s/wQu5b4vuUPezUu3f8dNOGGwsPrD
BJnhpMQ5agVe0oWr/BUDq/x/563Yx5bO35RKaJPlhPrXAopSahbx7pImQIqs6zRi
TI8hT+hZrVZr9Cht9rKmOc8zzC9FtNh50IrzQn8GATSgGtSz8SSSl+sVr52IwggC
ZRwVPWnsT7ocvjoeeQFeCrJbJ+hfGbBW3xoSJMQd/fCTkwkg58HsZ3D+aY/QqK2E
Cd5CmOAIzU5dIjHEL4bZ+mf0UJiaG40zYS7OrRKoKzHvjuEtn9AqCCUVddVlDY3a
aMsf9tBxYDV9QMu4EE33XHqY1ujd4N4RLlpEuDE9g3+peyQk63DUiJ1d7hIJtuCh
AhoJ7yxGk+iJRXekMSR94WktJVOBtFcSBx3g9+YDNhtG/6uTVeNj99YuBz+C+Ll4
DbkEIrG/3n5DA/oaRF4HWdH7Mr6c64eegigZxjh4PeQMiRaoAwKgz8yYkm/2BJUw
JWQ8O/X2NG9r0S8VJGJ2sk35S+MMdKgD1KfED/XDAgzZo196dKc9kiVDSiEqaCKN
MbyKAiWYxjbsLu5t/YIo3W2xY5S6FFm8ROedg5/jRFJHEpOdonUjamniNWMFHovY
AcYpPBgwZXM8gxGJyYoR3uvNDlS1FVfox9Yw4vfJawSPhPNgMYk97DofE5oorpuH
G4OzVdg5zUjQnYnt5vkGjuB84DgPwzGNhpVc6tNQLB2Q9HKm+MyOXYyNZdZm6xue
tZj0KORaMi8i6EqovmKgX6muJjy5KzGjbv4MthdFoncyrLDifqTPJ7WmIhFvkOPQ
Zg5073T/0FksF/wkq9htTC0VX1STF3LA2pbgjjdGTR4MwfjMUl9lrY1+d2oTVzl8
sK6chWbdmGT4iWPI/n7UKetbOv0Aip7ARBm7rUDDTzGEje0UhKccynanAu64+TKK
4gX/F1+Pgop3HNhEanB7BPPg3wYPZCb/MZ6SHK39S5jYdF4cjLvOPfb2nji6ZF8V
TsJS7z0mI9mnIhLktnaCVhLZ4X1f81oOn3hK6XY02RWNofAtaj/XFNO9kHoPlNu4
W/YLiydRGH1297U0y74mfGHjNSEy//iU0L7zqN7i2uqXh4b1Xs17yhhtbOFrR9cN
GECB+YwFB+Xh/153Y9x9XtMGOfdpLqwzZiehc2nYAVBkAds9B9HaU+hWXzz/lARr
GXtHvwCvi97BivlCYJhLWG+IhH/axWgwJYv8h6wVGbsbu0Wrvxw1Op2VszQEDQv3
AhCvIqSlbOmqhKfDSerE3eSNW/hIdrRXDfEUVM//1vspHHKbs1P3d3k+y1CayYh7
CLB7a7Imr7do/pYNbNGlvRMC9fEmg0NS+APIsZbwslKB4NthcvR0j9JslnZQqg/O
fctw5rcLICbLwYqPQ8YLkTS+MLZTU8RBVOoAS5jhjzAm4kuwD1JqZPrDtryOz67n
i2QktfThmGwfpcmHkH3Q/wD1eRwAjqLGAvuY286tChmSHlQaQsNViO6ddp2fYYga
YoK0TU1oK+CaAk/U9+6OwAJpLxCWFaDHB4C+Ayc1bThMzrfDejdTGR/cpCruvMKX
No+nIxNUIdk5dfc0JwA8h7jj+dtD2KNHuuIy2ooRIzb06t445OderCNAeXjDumZQ
wuG8dCs/Rs9BgSjcQJVKcXpmWK5SySwUi2Sj5O2UroPLBHpXt2pHYpXvJTu1Sb+5
OgcTJPTSQapirJlVQv62vx8cml5zdyQSQHkuI2Bi6VnOO5ktX54gzF1Grnmg0ttx
mwqhmGuYajYTzBu7uLVsSms3kuDEhOZDPFiB62SOqRbxGKIabxx9Agap8VeH3908
feSZNN/sdOHkD6RW711OqM5krVf6a+Arge3s3nVqwFNDP5WDKgNXCJjhrgDZVUsm
cNWmnjrICsd4pAvzttcEfht7N5kTP1pqLl98CHZKtkFmZDwXquvb8ASvpLDeNOok
L4+vb/aWE6i0+EJPMzIYaZQCD6DMTgU4g8BU6bMhAYZ1Qyzf3t1jrA6GPnuXGogd
tHEx36PclyB956nPv0uk/81UVz2xbn1sgh7Kle/8YL8kdo16r3I9J1apRafzUZTr
9Nt8bNt93HuTLmLtrLv8LWoQUgIgOLbxNDJYu1DPLftIFZBFlY2GhPhVCOZNAlO+
zO4ljmfEzPh9auTiwZrErkI9edsh9N98cvB8Gg6n0Tivdu10DPj/NKKP3uZsP4UZ
JUfitjjynZpil6Bk6uLaIj3o6TVQz7uYwk0xKF6oXFWMDEDCWAPX69c6UgOBNhoV
OfikcfcMw7ZoVePDdEzweuQ4kYefNJEA8G7vhYPOkXbGAQMK2m6wq+r7OuKZIh9g
R4JV3cZHX4qP4aMMZ4+lsycfT9ig+TNXZkck/t1mARzVk4vNBlNC9S1OOzAzuFZ+
uQaTY5ol3nRM6HTZKNWHED7nj8LFJW4W1gAAyoCYigZJ5lZ9mvWW0YbYV7Sq9Bnu
E8Wep0GHNqZBot4miRxO3aiYmxwFVmdcP6vuQK2fodiKCLrCEcdTBLHlRMDEycQr
jRZF1/2eeEU4DhUqCUP5ClJjjJgQFffCG91UUpGdC22+jqZ57OuReygYVOqYVlPN
rAKtxsUAyN3vXM2INZoNETuDMn/d0+zi9aZ+zTr992gThj+od9O00xfrOzIhEPnR
lVYwo1C6Q3hEwwNlrx1Djx4M0UEobxyC5dHfS0MmGZgg7m8SwZWs8U6iA3Qe87UV
1qg80sVZeoldozzej4M9dZkDI/j2FqJAS8Q2F9cW5cB1v31qjQG0SJo7/8UcQ/7J
NAqU1EZDCVjQbbdKyM5FgYtJqSucPpDXurIheVJiFAYthdVHCV3NMbnzQFTDUGu4
b7l5E0v6J2rMtimZo/n6FRnii5JzDQWKGZyr4fOnZTgOy3BURKw3qt080mQGG2cX
BBUMgVbsDk8DiU9zHI902koeyG5sNup5SkBgJ0dyj9N9JeqbhheMX4B+PzJ9WWno
mVPggG3sWx7vwwOm5ySrunNthnnx7cmIZQNzJ6S1Ve51yxjjSLOa23ZJkiPTX/70
yzLveOr83XUWBYyFM8ScjcGiGOiKw7ElLxPaQ/WdwSOs3Nk2XmNNoYzPl34uqxub
cJASaYbYFCloTV0gvZ0Bgw20SiEc8Rv5Tdi6sHaLRDkjhYvrjqZnSapZaoQ/X63s
faE2A/eNbkfvs8FQWiAByH6svdP0ft4IAnKev+ibUJ4TFqnUWrEwwhCC2DEbhpoC
bDzKI2pKKv01A1QVhzoN2hQIkwnnYWZbyx3V2PUJohymFDhh9HfsX3OwIkHD9q5T
gGcDg8T2Cvt8kcloTaHqbKUxKjh/1HKjsEBP3gMwxEptKvL7cs4SNh2UwxV5qsUe
e+OY73zfGg+Xk/Hl98LBi91Z7iZ2ECzTxAI1bplTCBmKCdg1+cUhuHK4sqkB0FYa
KjkuFzLJDebKhS0HPICcTjfEjna206hH/FzuDN31/MVYX7RvboNYw5wv2LXhjBus
6lED8ISdkhTaBv0C567vs/53YJD5hTT1dBvcYlJgyB4yH/SK9UFt8hI97t1K3vWL
VUqTASoePt9uTq+Zj0220Cmk3194rVn2q9UFEI48tu9fL96DrSJXW9Je5TqwvMm1
DYAvz+CmsGsHRFjrzQBR2SgS/px2ZH/MKmE3YY6pwJR74K6bOARgQxR2sBmpObLR
1g0s9K2WhDrEtCGZSPxDbxSjceuKXrHm8OComSJa3KYUQRkdI+sxDcZTf1bzph5X
zYYH08gjaaFcxG+Shb4nrJ3TDBz4Rg43jn3dPVaY6lTn6wHEui+3iWAoM2iW4kS7
aQB8+a7DBfRNFwW/TkJmsXEhzIqAayCrObSumiZezb6VVwNZcTTkj5rrYybVoJAy
wNPYf1i2Q4Ny8eNVhQD7lQraPZf7naIxo2CfWH8txFarCvz6+aE0P3/pMTjiuw29
+zMFJPyHBPsn3cjeR7VWLY/TAf11ql9SzA/bVnO01pTBw9+dZ5mkQXFmpIRnelgl
f7pxYkOS4vC1MpgVwjek9CK+dbcuMlwovHO1jED9gjfMrokJqc0uIP1zJWodc/R0
Bn/7jVd+/ODjdIjyFbE7HHHGYal7nGqglnd3lGltoeGp31t0cbHwxjd7Vmmt/Egg
iAq1nk+kqLZ9x1TdftE4xz399oK5YSNpS+JwdYvBZTZzKrMt+B27Dacq+soW4kz8
PGjF7SaHTgbeTq3spSEkJOTb9yoyguvwKcVlBxXuYXRYIReV3QgbYkHR8JHR+Flw
aHqQvxUQNh3N1mkGaH77D32Pha79w1B4x0wwthhmb9bcJ3Tp60gycjGTj1rKjnVi
nPbClbJBjnZBl17arZJ7WNHt1yviYEx/1T9P9m9uSjSZapbBtdxHQYNkWohmQm2z
t6d7ph0AdsmvqM4EzaJ7hKD43vdhlmCwCFUjn/vAvSw2lHHnHePBlsYo8pXU/39w
96yF3fqlHZOAhvYytp02HsR0bB1cIvwmH6dyDbxlxh2MIcJT0G3aIw3NSur4Gjnw
9dWrhaXC0FMnKpczYIMoo4+WR8oYP0Xpt3Im5gqGFIpeBKJQSg1TluWGY6X72Gp2
Xcbx7YEHx+x+fthtrdZunJxNAoyE41OcCQFUVMw1ke8ow7Z0rPyko2IC8UWZjgwR
R1d8U/lc5hhruJY9iOOXO0y2aqIBvjDgturD8F4iYid5ly4DvVfOfcfCfR6vAJWh
kY2BWMRLZ10eyt2COo7Ko2Qb/X5Ykf623uhMl65WjhOOivaxLBK7GVKW2Z10I81x
M2O830M1W68kkEX8/5jydU1X6WWfFfsUAeVALqyZinn4JDWTUFc86tSnCGl+oKTr
o59mlEu1xwj6Eeb7KJ0ivNUOUxUdVma2Ua25+Iw9WKtPDEpP8c9/Km9xIbG5R9Jl
VBSqeNZRrrIHSbliPXdc9AkN7ZOHk/FVaOLrNefXm0RLUmH4E4ohe22vEKqnkDP+
DRwVMxgGog5t3Hxc5FJC5hD+iZt6MwDRrJTBL4/9DIrunedUcTLuuhAijqcjjhv6
IqEFFl2IZUa5nxzN5zgqnhHQisHI0L+35piFQ9OLFQAMXeGmxCQFmWkRqTQlYNd6
YB8s8k1Cc1vywYbaMIpPUV4FdRyPszA1gG72lOy3PTaygZdVb8Gbj/65WEix6nQ0
YPrX0REzQp1b2Yb0huKoarYj3IItzuu9GK/FHoaw3NU7wAdKAtht3WGP9QRO8MWD
IWhGjH1rZeLIRJ6DCV0evl71HttPiUJf1lzlonlajZOAvUxh0znXYKD1k3X8zqxo
PyyRe+XQU2pN38+nZmLL17VS8C/La7snPtbGfQdMDtEbxcQ5bRuJErZgziOaze8u
X/FHYUrka/Og+RXHwfpeV3589CUcHRrPv6p/X4BrBxO6CcVhcR6yjrtsm0F4O2H4
VYnM+IDgoDtIBW79E+KyeXV17HseM7LqGj+8gULW7jXHYveD09M3dLds4m8NbFnv
xRVdiEcxmXRN+FTixB+UHYOdpUX+RY5SZwXuDMjqVaNMF0kMw5VreXvy+2pQ3fVc
O+MuAM27Cu8VLj/Z+OjhNs0a48Z4jQjvki5x6qLpb2VDj/1wEEP2s2dElzIuHfLt
MmsshGk3gcOO8M7OdJpIS5WHHq1LmUyNmPdaAmejlOyVyN8GP3gLfj6T+lNOiEyH
ZK76VPvtvdy8fLFyub1rlUtEkrCC0VwX3s6mHUbEQRZP3XTWQjTR+VHMH64luShH
FgH6vmgvF1e9wwmt78xbLUM/3lGaULGa2bpRyivdlBWhRbTeLX9iolWPck0i8nrQ
X6bSzSkofRIaBX4ItZ9pUzvGTzQi2Zs+OyhZ/hUdiGaFyFl/RSgfHWDGre5kMEYt
FmPs1ql8Dpuz48JE1CmDX8XpHZgiWt19gioTL62fuHguJ2uPvzm+OGWROREBR/x5
NMHifx94aMbHqcVmPQxd9dxtcN4xCfRyHzX8ub96Waew0vXvNvbcNgZuCdACeljk
5unyqkMO/xfpMyL9o1EoXR/cKsLIlSGOINPRebmft5qLoMhvjj1z9/0yn/R+L7K7
mS+Owl17Q1jSeYsAmhjdnSlugQ9yO1QBw2lbEjOpXbM4Kw079wEetcrdCoiHCuNR
NL2YMj7CbOcf6CfQoUaq3VE5OqHkqjW12q8JUsCt5wxa3+gkvDlJLE6u/5oPZ/eg
p6yyGsr75mN0OFBQcDaLrem9o5U33w7ZEGxBWrwtrA/Hhwn+KByW22EwzhVlrnjz
bsTV8/WmlZ2+fsIsJPjeShtYyd5DXyLN/2HeO/r0sCxebo3hlf21YNVsV9LsF615
UilIWdcnscEkNUgWC4UbKnCcX9j8pxzK9Xqj/dNNwmEMLkimA3pu28kfCJBnuI1T
gg2QhAbPyrglrFcDCRkoYzea8Bnw4Geivqkn/76Bq0++2xNfDIAu4IbJMLD5Fbo6
fCS94hf1BGZ+qIAHFWdILOhR1TeeBk/yDPM5hrngUbg1Yq2YYO3bOzsTAIw6surc
t69PbN6mhxeacBC31Tl0NT7K6T2a/zjwC/8FGKqhx7PFKSPevHJmgmJWEEPlA2Ap
tJMBJHpns+Pw5jJaJQfQqxi1IqR4XsCx7Iki8VmDj3l7KnT/MqoZY39neLh8TwU4
LVhBetfDghBh0fm3p7k0RXK/e7OWP56lIPD37bu/ABQHObmu5zWByWk9xj02zMkr
VrJy9d4Yc9aO+9sPN5DBOFkd1kNr+/yXtLoLzAn12u1WW5WEN0FSCFoYrKUOJ/D2
EZqNIC1xefLSpjkS8G3Xz+kNGnbKYxOK4m48wnIBsNTDifPqnQ87E02HUj4mdoA4
eXL3eZS6/PHv8jlmKu8ei/0On0mmKiqj7TAZGpR5uJBsFOxYrQkO+SRWuDusHCST
c8miXkgTqbyB/Vf5hPqKTnWKf8PK7tkPp1IwNTia1sMf9vmRm5dBsB/zX7q4YBY2
/eflfLGFwb+RBhdgPYBNpKoxVPGH5MfoBtgQv8Y+CJCsyLdds8JmTXpDPmy4K+O4
4mU/P9a1j2Iut4L6QN0N5XtTWY5kr9/cdd5VAOuSBQrWBMWuEcxQIQEgav947/je
Bvv/KLvH1pT/7gUNibDSO5q0yeOklPo8+qO7/RnM/PMWpCVMZwzNftQT1WQ+LxbX
dXkpSsfQA2IpgDnB/lFr+doFlP9y9TM+pdd+KSFodZR0QMX7iKELLa97owi4KvGb
4eC3ZymWAspjnfMjWGQ8nN3ezTz+EyDK3NZmDRWUcr0r3bjitOcDVrCRrDCji818
2TK8ciSWSKp57aGoboxbeFkM28pZywP74KjH9Gx484K0g+X0LDyGpcG8d6xnGLHH
j7VK3+tfaUgN0lucI6AzYA4zSdQniOrdo3GnKu4+Y/zk4mqvsGCwSs9yVbpHqWmL
5rKPxpnYc9DYJ60fbGXPT6I8SITHQHtUK8ZgMmbql0fKb25dTYeISyE9TmrIJdxS
ofVrj85qqaTIkGSJp4ER6HpCmkHbrB0f0cLw1hZHJpLo5mihdxbhX+sE6qb+odrl
iL3nzBzKAb3yKEYoEROAtuiyg0cylw2SEaGQMvUCgJQZaRhX0SaDBtDYGtOqzhM1
79WWjjPEH6oCFKduaxLCUS6vIIioxIVzjXRXrlDSy1cakKVFupoubqceIefE2nfp
jwMjhNmtuvz2UdShikj7ilg3d9WIDCmpNfZ86OAlpcQdWhxYpUQkuj/6+Gvhe9O5
35OJ6yhHdeb0/yOL51NpGGKOfrzuhxOKjLv9+JasyGcp5Z9YXyvnDWS+fLyjfiwH
Jb9dmGg/VPwdfCXxTGIs8udswVgtIzkW5pEPMA6HUwwU6bP64i3fGfcZuMCvSSex
NFJZNnSpkYYH66iQcuPK34So7MT0q0DG85/6TB2PLtaY9dT4VcGYZFfPNx5vIdw6
JNm3n2UjhzBfqRJQ3kf7pJKWBJLNr+h4Op9GgcQzh11/L73XQ7v+wNUghQYQUsap
Lf/PTukVnJTpcMRQU6rePkKyJTZJ2DINUeZHPrWRlwgJwgoueEfO9S3V72k6c1WQ
9XG9qchzgnjmF+9ju4OruZ7jSjVIKt6oArb3SOthRN9qKhCc1NDSo1v/JoFHk4YZ
Yq88Df3lb++d9IkjctNOoMq3ma0RXt+FgF8eCPMxYse5jDFCRGVGS21shryd0nky
4kypBPrO7fDCJmgie3fJrBwq2Dl/hiGhsXlz7SNIME4qFy+nKdAblD4c+MUgxStr
ITt7eY+NdTAQzfxcFw3sXLvrvLIZjAkkf7xlukn09uSqY5prNUt5D7c27aT0gw0d
39LDMschpsRaBcUpu9E+U794qslW1me9NiAsOh/n3AT3SBZ9RRaCJl/BT+IQZ1h/
BO+HHNDOjvknZ1UMAlDf6DM5lcgtbLC7e3TJjtyHZgJZZOayA62vuMeVz6qEbYMM
PC+HHvc4gWrc2+o+7WreNkzMJ4DptZogji7xLLc1w3YEQwCvHfcTgzc8eCHXX/BU
CNNVjq8gZdKkNVr+ZxBTGtqg9V8/97Dswymo8HK0L1kU+bgUVvPmFGIajSbdWa2g
UBGbngAdH3lYp6FbhNPS/lvGvgZiFVQ9Pydhr4M4t6ymWzavBJqU8wogLINQVRi1
11vbTfwlNshlGqd+OjRnVauyjMSGTGimDuzj2FBVM99KvvrfX8K+9vwWeepDhWMu
lewmT5tFgnNdtEnK2voC2mk0a4NeyRwMMYCc7/CQzw8482RbpsHdi8ytFcNGTtAV
S/B6YfJKRr4osrJgm6sW1/JvJvGoocEEgxKrY+IE7d7wXiAkGXeeLKALV/oEqlNi
LDq+Z3Pg66GKh/ZDX7qavciny3GHUWz6GKne8xYoUEG4ggAxJvcFsI85d3IfeKqs
aiR7+15rW6+h+OOyBbH2s0qn5Yf71KFd1z+gZ9iJ4M1AMgLrxqhGXtEtrUXjqrlU
jv8oA39rz8Gtdbe+cd6rAV3rcX+0aI6i5t5wy24KltggaSJJznFBWvwLa2TbV7Xo
RWHXuXH57t3kvSxU9Q+xX1SXwOID8XZ+RrrzpKAfeW8nqRKFwGClxpbjHvpkw2Kl
ZyIqkUZpVj6yqzAwjLNfSwMQEG8/q5lHmNXcqZvA/1MzDO+/zI6ZJX7zCnyIT0FH
ds9ldEJ54ViFJAptVbpLi53TfoegwxXj0sWBxjmvcCsShgeNabWuUJNqkc7EVE+2
od/7vtq1Nrxrkz3Gdq5+FZA1HI4UgDuRvgxCLouSzCokRbUkVBZzBYymcc4jydTP
yCDYyPHxL+APonab3x8+OwRptx2F0xjktJHrunpg5qrOT1EOvabFtpPccwzez0iP
UwCd2cfaWtnRNyR04tfJYDqUpqOdcg7BEbXMj2eBetIr4Lp4P+2uGpZBYstrG5vW
U0s1VesJhWnvCULQq5kvWTcea4qi0F0VDy/XdQcUWX02Y4adA11MUm2Tnw6fR7p+
cPU1769FISA8HoqnnSOi22SGyTT9IpmQV7opQq3iZ6Lof0nvW+WLcU2edyqNI2QZ
OfEYTBY1je7NPyWyyErI9eAkInmBIjq7Zb6KXNuB8wXutlW4RD+rL/1y5DkSWcuJ
akMhpRV/MqVrAMalRkYRDkDlf7Ys0I6hHCab53W5E8XGbKrj9mzJhk/cnBVtaO/9
qoxwplMvKZ5TT1TZ0HFuUAQlAWOVvfiGnjJywRAZQTUHq2UZKYBBcbAorvQrjaTe
eBWky7M2LGdLZu/bF23v7rKinaQin8Ave+fBoNeiGb2Cy8jdY1XlRpcrVR/BtAQL
AE1onozIsWvWAnX6uj3c0fyKES7Pz5mWtLB5TCysyw5YZ3dOk+hTM2eZe/CLOu46
z4Cc/GM6gpfQEO08V4kTSibywDeM3tviK9zGvp5rQ66AVvc/jEuQr4tem/OtrASi
Nc8PKxHTtCrFk+84KN0NuG77pPUHotJdrHHEGf3RTJADoHc8SbCJjiTQnAfgULDT
tPggk4k3rOfwJM71xmG5dZbss1YEFpX8aA3HWuRGx+9uSBhsqEIfB30MR7MMmFSi
FqctA4GXywVu9NwIKGmekBrWzVAcvLEmIB4jAWeyA3UaAp9IiDR8UTUxxS0s87rG
9Uj0m68fsChF463gQhLFVbDpcxYCa09Pya9llp1U18zLbsVAL4T27jtI1l3AgRPS
GVTMzL33QcJ5Q+JW0EWYeNJyGxoOyXk+FNpFUNfquznYaUk9PbvhxRZNUSYsRKoc
Bdj1s2C2D9iebxccn0iR5pi4e5O3IMaNWdrEz8VBwZGmzYMU0JezTKHQQAT27avB
JRr6/MI8uccohgcJ3OYh/qpwDVEBPOfryVmQTf10YIIj35V/D+/Oje2LcORmSD3a
lg44yA1+/SixTLqZvC4gyGb8VFh7sjpQ3w/V5EGkYYeWwB2j6fXaRgb/q30quRR4
TJuh6G2a6XFB4cofYaBVTdQXHL2gOqOrcmMGcZgDPU0nnLn1kYndr6v1OkxC5MSE
UXJhY9u2lwQfPWXhGVhL+J+pq4vLxtLSkuIgz7hZcT6BJsGinTvVgS6df5oUrRvd
6GLibOezxo72DejLee//tY2pod6TMtrWw5kHvOtgnZHgAasztwyK0fl9c/hwqkOJ
YojGrmgovBpkmbPjO040WP5LEAXGlj4aQCsSKQ3W0eMceEhg0Tm/4GgY1R/8Q73Z
+g6bib8eeIRZ1zox7ZV3gBZkAQtJdUcP1k3ivkq3ZdSROJUJ4odYl1uj0kdgX12F
vwe7KVD0hXAZ2MNswpvYiKUCsdRJAPHJFloeEkC27T+PP9Llp9CpvNqTnig1cfaT
BV0SNkTR4i6EqTfvruf6AXmjbJy7ZYYld0Qz15IvlaopY4JI1RJzXfsgazk9CZOf
v9wvxIZH6a8c6/FTyKrmlU94kJ/Ujf13c/4EOkzIxF+2R45l7R3fhnD9q8rbeFFD
msL/eihvy8c7Zo/bbRXTqnyDEd+M2qBcuXZq5Iy8FBltCRld/M8mW6LqOre7f+PV
ak+n1FBJHPmYSZ3Gf2KpE3tLxieJBsNoaVR7pBt6zJvYrmiSU+/Yw22jmLgcyt49
pwKu9nOZ4D/8B/bysKa546LxzSl8vcZNx7TUD50cMTJfPu4WdJ93pjX6RfK2ia45
aAiumR2RQNdpNgH8rIjH5oN6MX6IbJI4Msj/CKNuxu2Du7FSYlNvGSm8ZS6LqwfE
q0xMsCEkQW++aZPBC1PzHdWTYghrNwO4lbvBVkd7aWP7yjqB3wKa53i+orxiJjaG
nTg8QZirB3GDUaAwPkRZIYUKUc9aQHjKL5A5EgnFG7S0uQT9ap1lSqmUt7xgW0Ra
OVUx74tk76THIrc+6vgl+sa8L4QSLSHFlbbiE3aI5kWGZxKgl6EPZDE5qXSkKJEj
TrJTKFSMCgOfMESCFTs2ddgAclayhgFiM96H17Vj9SAQgpgcmhOiLXTI1TOO1qCY
ygDZjN0OtOR9uuy9yVpsCE+ukj3MMdURfuGevWtv7qD4B6EvnKQ+T9XWYOON+MFd
GeO8HUO2LEVGxn9nRAzvtG+QR4g05aiqS8yZc1tz8KiWyouFIzEbI0tlDymeM4ck
5Cuo8LIlvxer+ieI1H9HHbgz8k510nU5GphHYP1BYva9YgiLDlrM5VzRs35CuQkD
nvV/8PAIRSKGiz3jaNRODq2g6y/gESDw7UeAYxCpXH1KdfzgBxmw15aA44TT9eln
PsOrTMo6RMa8102iu72g5LvD866Z09VGGOg3YlOsiDIm6t1ofEzDu93Kvvry4Hwg
rRPFvtZqKGMoTrn9cKLXr/bhQdcuRFDAAr+5P4Bqe2gHw8aGytPfqoaIwtrJH6ig
ZoOPL+LzwpoqgEfVp0WiMYpbbO6dzZJpGMVQXSkbid1tN2L2FRA8i/Xf9jz4/gU2
rxzb426bCBXyE21BxF8LeeIaOheJ5ZxHOnnyLTsp2bD6kLY0XmPpcQ4A0+DGIG8g
5BNR9lmElWYVK3K2FTeVIJ2kFvh5F7c+OoZrXFqHiWCKEtoQsDBhhhphjfQGk8QR
cnrid8w54Ghy9j9R9cYA0jr7/BdS4ksL7Xm1OHO2CTIiKOo5leQNK7tgQ/0eDfof
TD5SViOxd2L2fq9vU5hLqtK2WCVNsV6VfUq4/+vMeCFxZbZh6y7PNYMDUEdakANx
REmPNRJLmk5uXjb3Zwg1MxwtWGyucDocZWUiMCWr/ePilyQ4TEcA8QK2eG1nwx9w
+HU0RWgEf8tLMm+owXh9QmQ+gFjoLlkpWPSe7LbJM5IpVvzkpq7C8dOtih5fJOHd
wj38WVmxpZdkwgrfiqPWhHQyoiXHbponb6JG73lcgniB0k0jf6Z8x0G4Nc4Kp45r
PtD6qK/ZraJp20rU+TFV/kTvdP5vT53YLZOVk5UW/4/AMs0RRM3fA6eo/EijJ2sN
8xw/8qAem6xBG0PgRrW+iSuJrM7GOPYCy2rRmAtTqWv24zv4H6M3Xt8zeY+ir/B3
twkezKXz8QK8JMGJG8jVyo5ndE1OZzyvVcJbj7XcRaWC+sfAFC3sTeYunMtTdjIi
An4ERV5dWgrP2ekZmshnUDQ0JxuXLymVcTepTSF/bIqbspvotvtlWFDsO6wNF+BJ
qITEgyYpychvm/vcN19HXrDFG9WBACbgnmH6rWA3dLnp6nY72FCy0ds3BmYafeY/
k2F5Ise9AksYv7+MbVSggoyEhrR72hVjYL7gwMV+9MVnz+SJi0DKkWpMw3eHmAUw
NO5VU6k5lzxecj4QNqVDOOQSqnOcVWVAxV/BjmWQv1AfsrNqAV2S02QSeprSHoUh
9HEgaVyhsOB59QcNQt0cOLJMJkRxZAzCaUxvK23/hG51s+Zj174+SLQLcGKanlPe
SwFmvgrVH4lT5/hetC03XiYG8nKoa0vr++TFFX5TDbHkNtc0lzUwSZydhmc9OlwL
FsWdWEW58tjk+W27ov/9i34bmj8K9jCO4ogfN087wGJA3RuYe3RaOkXuolka2fbJ
yc5A090qkgfHCser5V2+kNgYjjFtDLik3wLLVFZRVyN8aWr3KVrkT5GpJayhT6LF
ab/x9Ocykc7mRvvWwDI0Y06EIDb6yVWYPrZY9+FBuZXWOqb57/tkJpFhI7QjJcGj
psFZpdZUg9Wc1EICUq6awgjCPboEREhqpX19PEZsgKSep9Uh9q/cN4soK3zx0yD6
gypfx2zG7C79EAMxScLLC7usBTOiN7dIrrFCV1VMgQJrwINZA5PEtl7rFLBV2o8O
E2akwDGloHtgEZxsTYI5clhxa9eVygiADvxAjaO2qfTfGEgOAe84Zt2JRXFO5N1Z
Kb7eCtgoIkN1g25itu6qKlT6mwD8f1AZTzDaprQ6xTBm4Yw6Hj/Uq0HuQw2MhY9l
Cr3kI40GY+OLQbcwS62Vx+vTG0vsUJ/ey661iRJ54W7JmN+ISV51jgDqtUgmQP7f
SgWgYNwkkOsya5FSTPBOCoklipE+pSH5qyf1azVRYkpqIWdDOi7nfUuzHptfPAZg
aXLQvuTKLHG/K/VCIW7SWAd70DRrcH68JY6NZ3E5SHJLyLMbiN/IoccScvWW7PeJ
gPg5P5GSJDXqN2xMHqNsP1mY/qY3qmSCN7z6ELONjO0kaM2IUcO4UFf0Shxzf6ay
1DVHkUGIFQFAwRsYQ5CWJ1MRjJKMZkgBrHPXTDEMxIenqgFasFWCyydyBXp9qEva
hIUIdbdiWTakKq2K4TNBHB+qDzgx8gecK4KRSav9ewnNrwhy+UOP/skZPHP2ocx5
pbShyu9E44iyalR3nCG9zrnm7q98Cn9kAx1OhMo3KLxDJf+2Q6N+/PK0fZWUhPTp
JTFdYe03ufLVNtY4uAzJMkNu/3DmcBkmUYGpQv5DhoeLPrSfK/c9AACgtWJt3giR
BHLtN4RLYcCMYjgBnOgdp2LSCf5nTGH+IDLrnxqI3+Z4rsSZBZe5uYOVPtLIZ0Si
9KeJH4QrLvInyRufKV8WNWVCSQ4sbwVF9keJFwoL5Mx0qew+HwXCyEA94Un8QHOL
7+BSI59LEuWWDn2QsAbz+JWNL4oZ2vitFZjgzW3U6IFu/aB+rOexOO2dHnPkGDYQ
CMrmAGOln9tWrZDLCvt7aLMH14BsoTs3G4/BMTMuqVJglQq1sg+05nAaZXBJva1Q
ziiYUXmt4/99Z2gnMqbuNZtif+BPgvsuv+sdp/29nDMKcDOHHYOF6GX8n81Exe4f
Qmx4qbLzDTFcI3nSDQQ1UW+Ie+S8YX9t927l6E738itEYA5k2gZGCZPWBxysDcxL
BzjxBQaqJCrYVGnzeonfjmXXvS+gXV4Y5Ydj/99A26d9pP4CT5gW+OwUztxOJ9ac
pXS912xiwowRNc85OZ1fgiQolHzvCKGIs8v8oscl06rSHbVxUBVsymO8dExchXWi
sloke31tTZ84Gt6M/lmADPdKy5nfFRGAUjmQsOOTNIokPcAJT8wADSzGe6ZQGTcQ
cva8b6yxbogwLfutjjDtpL2S5JO3JA95f7IxmROsfg7ThuHaIXOpFOt2Bc5b0g+m
xWRF5Oyu9CXXXl6aih/OjhJC+j9LQQrJVc8vsEu4j4wYH6+CMUJOCB5cAS7pj6iU
YrGFkhRH8VspYnhCufp4/q7cllfoYq4nuJZLNytQFUlg1uKyGg2/pzbtbnhW4DXs
/7uNyaOXDXub0CIuYprr/ni0Q1fm2nkKR3ngNARXIhC81gH+QTRB7LLy3zj2hHv4
SEN5TuorPvC8gS26TXk7sHOnkBbO4WZbQ/1UMGAExmH7d9zJs7SVxU1QvuVSDYBv
8ufielrNn3pyre3ic9JBOVwa0Qtm1U4meIbebroXk54w49p/k7AlTn8MSnwf/zsC
U+EAQ6oYNqc1MfxLwG92/mjyMKx95xNvcPpiw9on9/PjAjuoWqai2MJEoGvDUBdq
OSmUl9dW0os1exHmWbpQmhpeknOcAYEMHXYOrQf6Ud7NalCfo7Dbat90kY6euTIO
FA4Y8b82NlMsc61hY3dsbbNrvKxH2AFHE3IGjTbXfJGg0P0HJdzi7BJkXUlZTabp
NBgfL6RlvgpLWzEXVOB0Oj5ozKTSUpYkvBRUhEN2IjQg6i+dnt6b1C28Ss3akoLy
akURuybU6+k3xR9ASzDa9jH4o3OsexcUKttYauv3zYZ+LpgYDqx7pSEZeh8aJ0io
6pzGGpSB3P+YKi4oM+V1eY8c8zmM33EOIGwkV03q/DrZCRXqw37ga54wgwsw41y4
eReXolQRg2Tl144fTDcsKpk7D0A8dZ6Rz3o4t0IFy2ai0s0kfyHuDbbfbN0UPYJx
T0dQO12zhUTvrPIF5uRqZvnn6+s5md/sB0kzUL1izoBr0nsCHgtws4Qyb7sOs/Om
nrpPox1q5zq53dXGkz7AH5Sc4rY8QlCJSRXXi8HogHiVnh+o+dZnFUVdMiewWgTZ
Ld5PT51jbHCz/QxVVOxxGpuf1ESi9Ab20eNpGJI2umZCRxLYtZeZN1krINIyRet4
yz1EcR7E5p5uwQMgqmlxLMuw4mYfB87RDHfBhUYBPCtsZoRO/DaPAQu+rWbynCJK
0Ux3zsCIPjyaFR8b+PzN7pfRCFKDF33YKBAdxMqZ73UXWbmbvoeQYjwrKsycyKQt
PjgeCiGAR5QjS+ryli68ilyRiSRMtHlG9lnIIYVChJK40Ba70rGZNDNDhkvf95zH
VzpO9tmBkwKTe00oBpIi1Ow+JZ7lsxbMXrTDT4EpLWANENzs3Wb6BKAAIthkFapk
rPlhjTvhkEYOLMALjvkLHZwZg+ZauTW9DgGdh4B3n5/Z/dWD0CJLj+DurjVP0o7M
B0jaN+bWKOXsUPkjARBOzS8uooQrykP+etxQD/KXAdBAFPbIM5TPwjO+byU/LpPR
0X67ho4ed1BxfKbhAUIDlKL6hF5eRmTlNdfKb3bb/vr3NGflyxINtxDheR+Iasod
5ThxlIFq8i9VBrYiil2Eq6F0iKGiG9bETI+aOB8FyvL87eS3EJ4V7NquxlvWoP7n
obb32I++ztNpA+r3PMlA12gvUMDlVBSSIluidHtrTIYQMWFqY/RG8tnccc9WZgA0
zpO1wJ6+TZ/Wr9JKglTpFVMfx7EKFflGGOo0vbQAbjfEYwxYRq8k0RGcOFhmJxp7
wPXHhG3FDDu82ITv8+ywfk7Z0qM5hXfKhX7Ha67LM5IX93P089HJawb8OqvGaXiQ
d4vx6HS1HgLR/kTB9/HnSkE7SxD73eJFw7qC8wPluD2Iii8WKAkNsQUZSxmSmCq0
/nU1CfCFZ1Uifm31VKJqwLvdJEeFBLI0yPnJspbF09Q4t/abb7EefyVUTj8PXRcY
1GNEdPDApp4aVjrgCIMFuGFyicXotkkjCJdE2miyJ/IUDYqeQYbI3OUceOMa0CJU
Xqv36/L+PbWzdPkCB4k0h4j1FwyFKT5tskok/dmxcu4Zoak4PCiKB+R/nK5S3I5z
rU+mu2p4qIcIGGge7wu1Qv2I3JHRHFQf2qzPncH4G1YIOwyIQxLwLYKLh922GGI9
nIKVHMf42zUwBrm2LJ0yBwQhx5ivi9xzhUPEJf/cOGEnyZdr0hPr4rqQYw1hFD21
2U8zvNuCWEGY0g0lOic7/bDx/2PFOckFpfHv7t344CrqktcczZA5hMALVPZjYDgC
882if1OPhVYee7FzuaapOymbEPQCFfY5MIaDNhilxy+2ikYxib/alhoMltVBPFhz
gJYG2hGZH9MVBZDAGNTM9z8ugZYH6hPNgTEOMjG8b7dbE1OGyoSp4R3CsC+SdKOr
tcs+pUBv98MDJzZSjlc56IuBNlhi27UuR2ksx0BhCbrZmnWOcV2EOA8OBCoxMBtU
PZdBJ1aKdzwFI9iYPnHDk4hQXYqMbsvmriXOhy25KzAce68L7rfpPb80NvQXMUN6
vmkENOrmLzewRIkLkBfvtUBXy8nyICJsLqXk8EGM5Ore9if+XprLF32Jues+UJLk
kAXQwsj6PDH/Yn6HfrweUb2LcD/QAxWOkOhTzJsXUdFsXUGr5hXoc4bGi/+7WDQS
XhZwWFg9o/jbBj770dTp2bbZGpg6kdnIgKTUsVUgMfhwkVEWpvGH513G7ho2w+gV
xr1aBK9FiIUXHEm2BR6gqk8F/9Odw4fLhkgCgpqgoBEcxmOSLTSlFsdo9A7oimSz
W17lEeXG7rvYfxAHJZJNqugpfzoBWRqggRrHNF2ozn2JQSd/w1Ax1vvfdD3ER7OJ
gILjJCaCiA81WcAkdLt3nF+YVv1ooCT+aoacM1Wg8ghqjz2IryaqUFn59pIxyr6r
aor1hlzzfbpizsAsZJebBqu5idmv95i4Jd/FOeQqF/UxKLbmxjkS7Nf71eNgpD/x
VtSdaiA+hZM5KFdIeJQbEcwfZmMT6tAEOLYLQKY8atjBC3+cugbwRF1MourHFN41
4SvPb6nK/1gwKZgOi6UTgyPyLSBhz46NpZhXjGC5qO+gGigfOUgxfWOr51gE3mHQ
un+m8U7LB3TvWWATUqFtjtqRBJ+b1rFZA76JhSKvXs/gNcHBkZRxWhiIrC4+5mT5
2yz1DCOEaqjaGrIB2Y/YqZMyfruOs7zb2cq/eCbUrkRBsUe9H6SZ726+crsN0ZMT
Wa02pBw917yOQcnsyjACeRrOIOm+Bhy4pEhWatstZdB+s2GLewn6/aYgPae0fJjL
oupFBNEEjv9MnKr2NrM8BdksMC2pVJg7MHbyTJhoeZb7fRemP5qZBwG4xN+yBUkx
Tssm452PRk1gJbr+K4NpWg8FnXXyFP1IkdNjRb1/vdmXJDYxNvQMp3xdINXmQvT/
ooq14OeYNaVbjj+X2EITqORjUl8XWyonRrvZpAYjw3/3Usf0DhTaMxghQYZdPRmR
pVOe7ftvb583k1JujPzQ9a6Awo10d3CzBk6TCH/YV9EY24ykyTUyMTqVhmcFdWIt
WFLDSEI5m4TPfvvzkvbgfmyDpETrwYkZnQmB4146fvfcpcYFxtlAy/SQ7z+T37Vf
0HMcZ3XH1iBxF7tOHEaNXZvLTICcIrGM6A/8JdggZzAVrlLAd9lQQ7NoFYLIb8uR
84UYtDlAEyLqwe1bLAvkZR+7EEIT0GykLXKBkFs4QY9p5vIxNROK0JaxnN7HAOu8
skA2/SNysjBE1S4g3F9ks5XBPaC749saoBGfG6Cn4MzhjI+5Cbja00E/SzkgFkoC
/6dGnTwuq21mOsJPXmQxNhEmXh4ZP3+4DfnkbFZDpKDbpwgWfhn1BRSQDnZWLORO
Jc+iXemqQehL2bNnzhvq3494rFlK612B9yZ1j5iA7tE3qeZmDmvgkjjl3Ttzpl0B
mxFiSCfOPVLe9nJNOT6h267YE8CjolvXKUIa3AUeN4iblKf8Oa6fAqe7J6x2SC9s
zdHhDvsRUpyneDIEc8TrWT9bVjHmd0Vf7J8VLcpHcZp6sRk8AdCzOW+NkCdJ1C+k
YO7gmaGXx2uwy2u1oLAqszlqRm+6/TqvVsfikZPPtb55J1J++VBa8Yv8DuaK0YIU
C/Vaivl5o+GSIQGBVL4GuJn02aGCd/9Yrq/db79n6AxxJdg7ZFQmLor/jBP0hc3F
VQalttdeFMRl6Kv9mWOyYXdtjgi34I/KKew4l5yiFZAxpvQyEh8KimhZOdq0HjAo
r7vv0D5mLKGRtuP5ave7IHDtMTsqzS4fFGd/UrRRezj5IEfMflOV52Swd7tpaU8x
oRQ0ds/R91HwodVyapmE9D663JyJgCslKjvAx93X+mPn6w0au3YAmlN/J1YWO+ED
6Lq4iZ+4XqRP2Nxf5KSJiaxke6o7I+9m9ELaH4S/l2O++RzZuW5cQXLlh7vCfw9H
kqNwc0FVLLOCi+XQP8wcs7iLrVl03NjM7E7k4lHjZw6+P7IB/4y5bMdx2KPtCOk3
dAAPVOpvSRNYaIdi44RDnSVNfrDyaybwXUpHJ85gZZGrkLlhUvOlzfDx0i0hk8wF
BGN70gY/oQ73DrP8GEQHMVbQPhnEBunpCcU3qM1AHFwIE1GZcjMlCl9ejBrV3wKF
VPUDlrR40ggftCUw+meD4DT9OnXeH0PYTJfVmSSaXcQF714wo0XtCMNHhfAZWO5D
yt8N3cmhNP0c+GklUiho94i5325B0Q27WAt3Z31obZfD6jCVTTLtBh/Bs/3F33vr
GQCFhREXKge1lHrGfY4WbMP1PBzeq2MOkWs+yzadMkS7vynrlMVnxM+Fub0XiyX2
yNGU8ojmahmt5g3NJ1YWm24ZE/2veeC9SyEef9nN6A+MSww0jZC0Gvx2e/c0ImeE
QMzg91ghaFD+Kibchurbs7RjcK1pMhFBUhBUX7n5ry26BeH/wJnNub3LriZc6nGn
3wBDNR9dMqQ7KIJAm0iu+y9kGS6J6w0VDNLNo0oAl5rwsIFTWJYHR5xfESWbVUGm
HyEJMMP4vX1px0VvcVbUKXwFNr6fGG8CMGTuZ4GVIzGKvpIPTt4qVw6hO3nuH/f6
4HdxtU0Daj6V4IyA1mIpARvZLJvl8lJPW+5vHWVBaXYo6fXjgMlNfcgFKiD4eCfa
ObRSIdaCD+B8JEIDD9G9id7duQGrXwkXcw2wPQ79RTeVAVKraEpp5XZaGniYsmdE
Dv53XjPVcM1aNugOEK8GpqUW3PkJdzqsdRfpp0ghWbwzm6BpSsRRV5CUIPbjQw/E
nUyCojDnxMfGFlLBL1Go967ekSNdffH/fImsqrc2zbuR9jVmvY5JtyO/uC+t8++E
Ys6jkQ0nXwwniqYPCuVIw6/x2saL3Gq0tjOv1AUrxg0PA6VoPfJmneEvhOnbIBpE
0/PMDmc3y9o4D0CFxATrB/JeTAtT4v9N61hcmgQFVYUCVtBU07Iay4jd/54X6QDi
HRl6Ze++qGQIGoP9ufURIIKXJeCPiql6CTpu5U1RI3z2plgQ/V6eeqx/D7dXv/S1
wHZ/XsdzADrG0H3BQYUFj+IIxAjcw2FuqXjP67Su1oj4ydnBVKUedmRem86so0A3
PNn7rX5Tle3UqBZ0ccJy8xTZ0NAZF/U5FslYYm9BqrmK6ugZEM9js906QtP9DE8h
3Cls8Oo/Vmo16ttu/6qQ4pqWTBkmO1hSC2BTQ+0MHOGTzI4Vac8kbOsoBqJ7pBve
gADspLZxFou6XEp1Tjo1NjcDf0tmag0BfZCc/t7TVomlNGEBfG2uaqHQaVoZb6cV
tOqY6Km5ok5YSa6iQhgHyDGTjSUImOlqz/g0PpsQRIJ1ykRsjH3tKDT3xDYem12p
ZGDIPjaXHxceN7lNO6cvPACvTwPdEBYZ9SvABfsGzh/7scJbVIEMjJ/cu8tdzmlj
rnO4z4g/l8Lu0bhdC8ultQPADcaWKZtDB00ren1tF7803+L0GidR6F+KdwG8BTYS
q5sATBDrnrbHwxXD/GcD8sivCbYkx4nWajxsFBtdmDMOi92o/+q7OaMeV7X/Jpat
fOtkHl+bb7uOkCWNQgTg1bmhSXyzTjzXrTkGNF2ywLlQVTwITz+d9nmnjzxgXrjC
JANW3UY8XH7TQEjs1uyaqy9+G693lplVtp1oE/UJ5CIPvaC38I31pAy8mO4KS4nL
rTS93cAUWyP4JCT/wF5d61qXahCvvCVUgCKWOVRY1y7thmARNLlc0gSzMPV6+Mio
0rJSEFEGse4BSEMIXON0URTAItbh8DYinh5A79Llt62MY/IB7JBPKWIrroU5WkKB
ejKeqclGZjbqFgFIoMpEtmm5BOAH89nTcxTKNAB5j/sxmidCKYNbSsUxnx/g1IVt
l0VwgelJDr5IY/wRqFfOBPXF6eEydrHBVomMkizIEFoSOJKCD5jCGkWk8sPAcS2O
W31sgwmaz+tx3NqqSvpVlvRR/jQFI0BHvrsqNdLA/StlVALaaxU2ka6LGYIOa3fw
z9gjEppbbg9qzPXkvt9nRsXtrK1eKTZT9jPUyLYkqTF7O8uv9jJR0sCddyiRvt67
roT9vKqIZTjlC8RjWwgriBb2aoWQHmxMwuEICu5FKtdN33cMCRNZeqqFvhHoAlWq
8vNV5OCGHrK/D9L7NBZHpw20TpUgjczgAWpg+wKUPQn+10std3GhWTxEp/wSYDz5
CKd+iWq2vbELYa7Qvg4MHo7joeq8r5bg9du+Y40GIZsD5LixVj9JOL5K/jRl1jRI
AwVOaua3pxE7Qj0UZk6+nPUeBTF51V7yEzXhKLZy8PtyaQofYjCToqNflZbWQh4a
3jW+lxW19+uqSiOdxEK4HolL+4lqLq/OBUjHXZFZ6lU6GO8n6L2phcUFGmVPWKLv
jcB8bGattC/jgVhPqXseRnMogJgy+tuurkXvCi0NWNhyDfjmvxXglk+/3mgw8XZc
+vZC8K8TT1cUizrFer4y3jljKvoZNFG5YIXQlSQIfu+/G8CpOmxGRLWUFMNrsRr7
IoYHMisSU5UY0qX7Rq4WsMkGVNnJuMxq+kw4isTAygzZtwQNMWvUjI1/vy7dP7rK
0/eng6OAjkTKiGF/eqhA7lNvnsqgqIcxbU7UhK1eUjQe1bIdlbTDJLsAiP4bJpnA
oEkzN3uk4gMVB2W6dKGesA6KGlh+pwKjMSLyJL31AtfYfgNoboZcWaghz0m91XhQ
hfN6O43X2X4vdPTSUyL0My5BsvFFwVONCmVMq3qi+SDkxxenVftBEmexbX+5DqHy
Zb6K9X6ONhYxzyFA6AI+6oBHXmfnvxQ0GMuoNdMPq0ogKo50dTdOcKNfYY2zlTZ3
Gy9J7xQRW4Ta82UtW0aGGWAX2YrEwOBr+8tuHICBD6Zhp0cihtrWybwFFlwHs5iE
MmJrLW6BRZScSV+prY7ctEytq1RLzoW6hfYVrK8WDYSQo8Jkp8bEsU0zUVfzIsRS
X7XY+9Fcy3tJoWBz9a2BrNN4IQELJNfW9EH5+BxGLvUsatvfh2X+YZ24bhpG60iS
5whwxtLv+bqLe1sz01WQrXRoRAjQiTAlX4JQKCMY4NlXog875t3C6/TCumjo0GRF
/TvDuo5HAyLtRCjIQXi0Xk3C1B+YWWUDZVJDbE3iBsTxjsc9uIB5dz2i/l1k8E/b
RoNjNqcpsoAxRYkbX9c79dEW1VTkG2OaPXiloDMGWjqMD5LyJbiKMB5J7jVssLMQ
VZDVLIZg50alG1byjCNwSvnKILTImWXuHEUJM+7El+/fPPptroJcbSteGwDo/4bZ
rQXLAY41ETyxVW6RPax5OwZjcgvHYX7EGLWhDjw/65KxHbhzByd3FME07B8Ia2t/
pLtVM3BACqwSBMQTp37eQEsFeoR7xNbRHi27TJd4PrV8geO3rWBs8+udF5MhCPcn
C6o3KajC8ofXb0+sJIa0nYZbDZOKtkMi9FYOepAGzyqHuLcHhoxryMqSwLLTqcAA
CI6DKUd4p7XhvQXf2jkckxfMz2txjfrBhQezJ0BsXsxYKQEPPE2dePqMX38UabvH
t3RSgmoWsbCKgEh3pogDHYgk7Fot3/dCt15XaBvunzS//E9qVpM958OlgC9GmE5v
gqNJcLxG50VZk5QG4SbXvBSMgY9/8n2c/4m5qQujj16gsUhjj2/GJNUn+kZLqrUr
dPQUGmOevOLRyv+L0mgosCS3FPzRqXzgs5Y00pMmnsMsI01IxL7uqN4x4V9M5XFZ
b7h+m+JonmzIkL/PD5+sU9EmhKOW5UEwhHz31cbu4C2WP72uv+IGrJXzg+EQxyKH
htEW9qXTgw6AipNjLB+3ZvwH+wiY+BqDr3I1TFc2ACaOT3MUSfvvKK5g+iqo9qOS
01PNYUL9RnHwLM4hs4IEl8wXOo0DwwNIyczLjYuW/OkbQFL7alql01gboTvUj4ot
szAeFAK6ucT0UTrCuG0T1aVBKARZ9dLMZjN4ms2mh7LJ0zIb65PHgkWXonAF8J7R
G7fE/tHkKnoEoYqEbcK5RD2JwAjbys2ceCO9MP9N6KS2iZgQUmqiAKKpqmHPHa85
FOOzTQztpX9eEZZtmpQAVTQYJOxIHvDJl2JXyUjd8HM5XiYdPmvEQJ1HE/FPz+H6
q86jAeSRp2JauOhDisF4ItRSKgILATLkvycOsxSiFrZV9+a2R0lMOv/gfhPUBKyE
j5pl6hl+dNTXvAIXnjfbCwTnUuQ2BF82jd7w0F8pfz5fe020dfVVta5r6OxgUIwk
OTeujQRoaJMlEX1DaG1LfoxT7hRepGdsIaU2qFgqrze+yh/OJn/hknjXMdq+YQQD
qrPCAb85n/4RJCuFoLD3fb3MbhAvuLhkvEeGfdlUuCJKCiC6Nx1zBBmjJRjks4Xu
gZcRNXBV0XKyUxbVYY03re8ivIEL2CvyrhzcKGYt1b1cRkPWWDV/SwfUIbnkdwN5
RZMmpSILwWwnAZCno9zhQKFxR7yfD2tfPBJFRa689D6qh6IKSejXCkR786agwgYv
jn/7pEIJUqBemAqjKL0VDIidvtzQIFCDB++y4tzX2HUwAISmRnlKNvzQfpYySuXi
BE+9P2rBrLAezycgBT3V7zra62M6qhaxMsLXCTA74rxYsEJe2jUI/5KUhIyziVxT
giq5p8zGqmvD69XN2HkQV75YG5t5iwHAJYArCga5JNA/qn8Dq0q2K1zFHMM3u8yI
s09aT/DyspyYmR0sryZzUhjHmdSXy5saLcptfcWlsWNhf0rFjBbbbAK/w4nz4A/d
loKTtd7nmAS3a4mjFj3D7LniyzNTgQfdG3U3DxtVFW2pmVue3LNotx0NGDQHB2y5
RspeT0MxYuPpNPk99CwoA2NesPhv+fkaQlrl5KAxZCPkefYGXk9B0B4k1SiuUfjj
l+PGHVnhBupFiViUDkNxYKq4JcjpNUNbx+rdvouRTfyXrRdAo/i6I5xT5fMPregx
PQEk7KHYSbhGoEQUBYfhAYW2+y4eK0lHXYADkKI+A4HCvti/ac/xsBn6lPLlCD7X
qFYmXvqXnzgQXnNRhfVUvby+QK/ZZG+BOsZmTSr6knmCv/v7sn6h3Kps5CWZP4e0
K/k9jsVF2WsdF9/K6mopcDFnym5PMXh8MqDqih36X0WA+KOLC+gQD6MJToU1MyKe
+wfB9gXfLGBh3DZ1QliaureXn4Fm5UsRS6C5Ej45wkNwnRBMDUqnCWqadNZ5HfSi
/01ymwW4SyF4bFpzCAS7ie9tN3yMMb7v/pAiuVO7m7fnzD4j09O9vLZwBRJJs5Sp
PQgNz3updwHbkiHSXos1MFBUa9wLkrAo1pHhOic/xBwF1SgnQEwenUi5BGdHEQIa
E3xF6jqhmfN/WM7pOEhxgrNDJDsAloilqusCJpErjRyyYNuKhdLKuQwhU/yJt8bS
VnE6TT5VkQP5uZ+yfiq1SDIkjfflHUPyU1LLI7sHCAKWH6kXNoaWQuvTKtVGZ/Nc
Zk2nKQT3r36492O8wcd0bfIXg8WjHoUz4/wKdt4LDHJL1i7v1rLDtDi+K0dFCdAr
9DF05NsPeA8w0BrDEq21KPE0QmEXy1DbyskXVXGzpvEK4wXjr8eQNQXA3bUBbcdH
qBhp6ebjKdCi2jlipk74GVQrFguqmbjb0LkIFfa2ENwjSkAbL01xQiN4udmgFKJe
8Uf7gOxzCKiXAZt54i7+hVOcVtoPJ3lenacDtiwzuFezMoDPTlvGFB+zm9cikD+F
t485kz+TlXTbQ5+d9+C8JSxhIUkfqrWerTNHxXaTkQs9yxHU6vxYE+1UwJbtbuIY
sgyULTeM5WOSFsSQD2rbJsx/XS4zWzU3vcFF1Jq91vS/a4rMBdKh9rklfbDAFeYV
0C8NKK+sCOObLO/rwvN5FNyn1eEVOjtUWAE95lC2TlqM4CEQbgl7juWuU8zdapZm
20zcnrS0pDRJSMpOAOE+AykSPoC2VDPnH/1Z7+SsxAbJ8EIq5/DmwyB9mlTRK4KV
GYa0cqSSHqaqwg+gtomIdi19p6g7ms6JkL/1zWP9S0/LnqWD3CfWQTdUFSOlOp5L
f2dR3eWBQ8KY+fnTeRZlX5N7AI5Lud1HLizkC8JDEqK0+C0xAkmsQwS65/wkoB+5
cgKGFdvqarfFvpn1UIAjXRMENxrnGsHo86LzmRGIydnmpdK7/05KsE99cP8tSiu7
Zo1zObLQsTJgYMESMVVzzxj1bG9TWhYFNXcj6bh5y4UA+pElHGuJSdlIo/AFqDAw
lXgDOCq/UF+rz6R0ey5siZiVosgxdkrusbYtS71dzNDuwP7nR76Q45xAUbhcWDTo
Jwm0yBCJinupO3ho07UG8I/eQR8/gGMRKhFLyJBrWRe2FPrmmEunk+dGJ/60lz+z
fVBTCBLcmzxGiDdwOnFEen4ab8JyqIEnvuCT5oLCX2qntvDEm9iTCDWxXJZc/mcY
+I4hiYa8bA8gR35j3tqc3EKX8pZiB8g9zyXTHuLJnbaMn0TQ3gsto4hkD1Dg0CRn
tuWOcbV2k2t/Lmc4t9pZPBwu0uNCp+++CfjOKpl0A7Q9fl9khcokaJYI2fujpKZT
O0D6G2YVlZNUdkHoDTYofGr9PQlMpJiEzXNJMBCAYlN5FK6w283jsGs9tlm/QSGd
VQsC1fnF04RSd9P1slf/9LMC01HhMMdquxiA4PY/ibhOjfwu0dlly9wRQLZcKm1R
NpExtkb3fKg29/eTb33Cdpr2j2VCdNbugMy6F9qE6JWp4pkRRoVpLOoW3k0L+wCx
OOlSdvbF0GEwVs7aCcXCTrl3K7S86n8K5VT78O5XNBKBFBJR/0m1IBTQuKGtau60
0186JW/FaMa0CD8c1c/LXyTfyWWp8B42YV4H03C55klfCmtCXoZrIK6WOpEl5DSF
omX9Ob2LQ626JiXHwtjbhhoppsJ6POI8Sa51fM7mRZYPZcWzwsLUHY0zfVWJeEvb
geYNr4kBQ3ikFPn4qIOPPutvuYcZ33I75DRpuzNYEwkHkvAPw/uM6M8KSqZKhS8u
u40ZkZBiHnnz/Xd0r2cCHAEGbGeJR347XYzLJfmD/feqHFCLS8q0BOmPH3X8t7LY
uDlPx8mzszkVl8yjq8I5REJnvIlR4Xw2sxdRDx3Xd4/aL/L7XFxSOZt6m/x3MPS+
TnL/wLbAMNPgsLyIrqrqxRcaZMmTEaIf7D03hEHmUgQEQLXb60YADgIeazY0h7jG
5NTxq9lM8lqBfWTdm5UV+O6m3uq+8mOJSNNA/VTU9A/eGvHBSkQXwroM40bQi8bl
/1Twhquq2WkWy182Pp24qgXvEmvn/wQUT0MVCCSJRIe40EbegnIsTFIdOdpm2taB
Gs97BC4UOXFu+LIfrUTVsTjvzeUAByM20h7/gn0eg2azlmzVwmuLf515c5I71sLQ
fhsc5DO5LGSSEPTleen0Ccym+McW+Knj2UroDlUqqldEsnBhyd6UEPUebdP3HzsO
VpDqwlidhIf9VAUP9whTFQeDnu66IALtOV6FX9a47amQfi65lJomHR/a/YTd1TMd
0n6pliHUeuVtpQ4ECr8as64hmfPXMM0bsWVVAh1i6PKat9myCMAhTExR4qhEP+wv
QPc/T0m26oDJCcV7pBqLoNtI1VFavZJBH+fKalrHV6TxbrXz2q7gBVtVCsdbUzma
vAh/Xdmm+kP6nh9qsMNTFBbVgB469LlE5O1zz8J67Otf9IDDS8rxO1ULZ1ZEbBAX
BybyAt+z7Nu/ho8+lo0xXd1z9CiMfbqfUf+g+hSsdYeaDon/qXwPiPGehR5INRq6
Xak9e9xkaM/7XBdarNkmSTr+kOVxwO6btueacFtFVkCM7mDw1Cq7unv5Tg/SqnYS
XjXGXwDfmX4jhh8a5rtJfr7kNKe5OpjGNUsE1fVG/MiQ3lVaeHlReZgfJT64OC9g
2M6MNN+f9t8bRmIvkAzv71QpWA9D2BAOtxAxN6lb0aBYKn2yEcIhbIeMcWYuXp+1
9i0zw1WOiuqrZm/zdSI0S19+ORqpsXj4V2TVB23XC/DFJ14Ct1gWG79y0TNWXxaf
NYlzCUrrZYtnV2/XaPRnSIbQ70tzbyIXsNDEd/sMp20HZ5eaplKF9Lt6apIx+PHL
3CR0iYI6KC8cWsRPXl/m7S/g6yoRv1Pohqjk29XUtpGpfzQKhgeykNYBj6e6pjAN
dBnY+jVNl1kwLrL70jvc6WNtYw0TzCPWNcODbLtm77TFGpf6+GWGp45nIVzuX+yk
ax8bohNJYd+lHUvlTNGKIwrd5izXtaIauoFkbOPPpSdRRp84dJxRL9TJF44uNy0T
sRGzbQp1Clk4hGGUQ6BtUknIO+TzhHY+2TbQJUo72DaAOTInp6O4giyDukk48814
0xLYwrWInP+0sn96t4pyYwHdhGcnhHbTvczPo0fYKFeAtLh8l25NC5o8f0oyrWXW
3ixGrEHDU7BYjggvuCajX30AOvrV/uiVVAXeVmRbpl57xJA1y0d14c2gMbx1RMvH
tbehrfpaAY2WP5BI/S0xcs065BXNNomFjQHNJ5iISPF1HPrsJZjlSP0//lG3vfO5
zjFGq6CTCuNO/gULSmYzDvv5ApYMTyXHDU5xNGML8hTLkByUGMESt/+28ac1mZ6v
rQunxCBisy26WuXfUe8bfunVO16hyMRxCbfD+F3igtHF/0g0jxL9dQH4jcnR+k9c
Dk8aDzfaUi+N/fCQkOl87toeADnHnSaHPLTG5TEnDcRC5ogpOwuGOQ3+xUJaeFlx
6uv4k6nslPQu8egyRDHzpU9zGFskr54pM3TGgwrTiHs97m3b2gdM++HbiSUi+hKG
qpw/u2//YN6lMU8/U6bVAe6TxfqmWpvvr08dytL74TsaS7/MtXLm2bCJDs6pL5x/
BHcknyrDSrg/liQbttFvaywGqTTDxk7CBg7VQUBDqi+4/UfPfeZRgWsNAzb72KBt
9npgNJ4pKRlnRBhxdrIvbPEYu6PliBLCdXvEC6aj28a7pVSOzoJNTKkLuSjUzaII
jDAcaNohrkt61dsn7NoLveZHlYGYaRcv+tzWSQV06lLAOOD9xeab7msmjCh7qBoP
dk+4bX7FuLFK0WlyDJufsLSUFL73BaesqIFand6x2QHWHdI61lIwnQr+i5AcWtYJ
lHxLG8YB7cKRRWleKi286yoy4FZ+OE5N/XG6spsKbHQqpsNmn1HOEjBjZXT9Q6LS
msHthxUjMvhlaSib4uffzSRHqqFpTitcNyZNttUnbObNRQ17Ertu5wGWjXuPO7W9
fLfjnB5fKFF+nMu4a4Rs1d9p2lYo7AB4U4+Sxxjzb33XcclW32pdQwu2Poua70JM
PyIdVv06vCN1yof3WhtWfIR2Y0Yb4RSBe2rM5jUEbVLBpavDScGyJ+FI0W2/K+bi
Sb6skXGub8Swn0fXhh3cxn9U5kQWjYjpSvkbq2ctHsY8iQnyasvfpR++zJbFzuoM
XpzIv1tlx8KXkcXHMcTmvf0WK0EX8a7/SnshlnF5nDtnHumiK2b8aBjNCFGhe+nb
NScPQe5hqpNj9DeidjbWByR2f/V6ZbiFF0wCl09ip0vJ11Y+XXjZDAmWMVdWysqr
O09JBo8FcIZylut4c49nMOHIJoJWnrZEgCqnU5iXp6jtlXeKrd2VEjCl8BiZ5Ris
C4kjYnGd+rQCB8DSWzEM+/n5bUL2wBbQRAkimWqDUtKij1utawyK4A/NNr3zQDSd
uUTtked7eznCF/Q2sIfKafWhJTd9g0LQ0lH1ydrlgAbHYHw0BjNg3NmgLNTI9qIe
MTniDoMJbDxmqD82L51me3WH2rJyKr9NyVPgZcz4ZHKTjJZ1ND2JIHSVsvGZWwDF
B67d1dX0rgdccYwDYP191mJ3LxCsBNEBZcgWIi3TkFTPMQzMn8JNq5gIdTagZfIY
aU+zzWQI9oPPUM7UC41zwsDWhPitFYIQO/evl1/tA/vpgNQImPfb1PYVROmiZb/e
zwi4aTLAunyr8kGWL4w2TrAiMx2aVkymKnZ0UAPffxrKtaPWAWS75RLgR2kRe2hU
nvln3nTqkLP7nUdTDdgUPx246FHv1JqrUvJZjUxkmNVrQxexWodvPVEVM9v58fOF
Dzm6JIcrah8IqiKe2krwT7wbHjkpwJR4f1xm3EBq4366dqOwpdXPicgUWTGYyr2j
aHSnT0MPH6V231bFtxeU92OMvB2qtxulMk55Sp2TvYsQX47GUQ95RXiiH+K2rSB0
KvaVOxLlnawg8WszqgJuAiCYRj8ITxZhdJxBzNxD0lMqVIEozml6MM4LRIqoiVQ4
uxGX+GibhLsnPFk08Ea3YzjS5Kv/uaSk4qHVyusnNpkiiHX9AuLWR0nFq8EtYWDv
Cnyth7rzDCSYHEPGrXdNuvABZgFMAl3uQ/NvSyEH88GeYw42ai/ER3WAHKtS2r+q
ZvkmVjzB+SDHUUEVJ2qHoupp1qnvqtlnsnCRp3+t4ANQbf9+dR0pFZ6e2RBpV/j2
hswmDmAyW0nUnFSpG+26XL+FhzYxMtE7BN3V+Zw1sDDKAby/1gleP2Ok6dDHzz44
322VuNGX0Zv9rrAoyQ2IbvlKdsfdl+ET4uIVooVyPI5xWbRasMtUoBSZNg1ljWE9
//NXD3s45nTlrNNb/2X5su2ChGJU+8hVtv9WEq3Eql+oIBk8wR5SVKjesrIDMpYv
InRopBOmd+dUVg3X7Do0KRystxnOWGG5nzmsNEqBIJx6UGAJ05fo5wa/eB15VnYq
rYhWZb/UX5ksaROwHXYS2pKGoBC6T//E5abOwQV9cRk7WRYKOAVziO+q6HAR3QOn
P51SITOZi7g0AoNom/JZUsMtX3dvB9OKBCkflRLCragT3srVSXwKDroUID9uluXy
hAtFo27tftn3yjVefB5h81dXC1UqPZVGDUNDPAOLMUni8R5KgtJJ0nfjshCKSdJ9
Pq0U/uG2eEdV9scpQOg/+nx6SvA9NHswOBjCRyZu+VeN4JzaDGO4TmlC7TzIQWA0
n85DRckuClfive5cGIzLfpzt3oQe1qszjMvy4a38vj7qMBHZt7bR/ruSu6vNod+t
Y0uGC4ZHQJnBhR/3z1ObUEfyASduz1Gfn7MXcZW/7uBYUHJYWBaKuMuwnnKPcRon
EYoFm7u3k+6DmndKapuSnKBXFfc7CPTsPZ3RD2tzVLq/AE6RZi4V+nmej3/E0SV5
uxY9B6IkGnL+q2hLLxxR8ZRaKnKshKw8gv2opLz1UF9drhGFJrX/SnCIrVUqAos9
BQzS+jr0xNEyZ7AxHP59CyuXiSNlTWJsrGh742Il7KH7Jt5ytIN6H9Ev2Fegwd6H
MOPsuwKTD5mMrZDQt0voYfLm7c+Wg33btSJQQaBScU+r/yNjKB8tfq1sCiQIYvyv
gnsw/uwj6NMcdhRaO2Sny/BALZXFBD1qmq0Xvkif4XWLaqK2KF/bENluc7C0nO/7
YslMlJUEEy3oH6qBvblyxJpgf9z2tzWoychj6SnNuN9gdLCW/ViKf6CC63P/Z0nN
V2Q1hv0GChzaYLflD7fEFzwlwedXC9+lXgD2Fa2Jd3BmTSXqJQ4lkeYiKYjZWrvI
bwabg9DSvpPxIQ3gzMphC/5JZcp+pkIMtuf3h+gbz7Zt+b+Zm5bRidES4XGku2Pl
2e66f/eA+SDUHr5eKD7HiastxvG6U29v3K2R2PlI65LPfsGt2XWnq4YpUenkqsI3
Xs0WO0YxCDLNv6MMdahK6UMT/Pb1B8rOUDB608w/BUqQ2PqOtG8TJnlGo/v1oB/b
RWcwzFWXdmdzCyg1zSnumex+n4VK19sXIbqu6Q8SKaVZZHB3gFgNlJHTASBxZSdP
p2g26qDzp+lWeloffYZug0kSwkb74WBgzOEaqOsFQ2p7OJMKI5lyrXcuSUs8qA+e
H5uTqzKm+Yk8in2v29j/5jEfUeGR1Xos2o5D7S+3fh9MTRYmpOd6TkMcdF96sFsO
1nJR62cNjzhZhCaAZj66RHZzu45ft1TFvml17sp5fZJnIfin5sGDiab0SXpM3feh
ouWdnJ4zJe/t8uAfhMmVNW9huFmJu3/1Kr+Q7zO880610B7AITHskJhQ4/OH9Rh5
1TAlWYMNNbfdQKeQ+ekOm2jUWOQaXmnwpXIadwY49ws8+6cFJtNnthfanK2S6BV4
/3PaVV3sha4rCIKMDzt3NdVns1iQy4DlvS7MmsjQs3yKd7rAGTH9MA0HuBdXcQYU
kvM8UoxOct18iV+gAySlBSxYZKOSQ7tHT/0NsEMHEHO4fArgv/qP1gHs5APcX4ls
iOO1Mm+LEAHMSn+dPpLacH7ORXi7pcYhQxAFpslfPMeTrrfcs1Ei5w2WhKNXhB9P
gX//3n4wUUcBaXaM/SOCDrenPwD8urHTAI0QlnMpZFcgzqLC/MbMF8Fj7z+T0Fza
opDYHztzMGBepm6W0IW+CEtHfrl2DF4rfACvUrbNJMWS01SW6lInfbT7xH9E2PRk
zRtlvsQxMzRsAZLqeKUtDCBPphliygRn3sSWkT8k/G3fkxZnnYAghG1mi0GH2ctl
S7s06xQhcXcmhFFnTZfJvnpoxlKxAGulZladoQZPM5j/435d7Sqzl7k55hWQSiP0
SqtrV68nHOeDGCu2mOHIrLOk2fyVQ8y5QlS7NxydYo3AKluJE9NZzS1pdqhS2bVG
zJZsJPdh0QpS4eCdu33rbvR3ggm4emf5X7MCTzylVbRrk+0hZSVqgyqH9XV3G6zK
R28cshliXzWnkk6emf4Jth8+68FiR/SDNP/9EM3FxauXYYmu1hxE4qkcqIk2jIs9
hEkNMwOOPm3fPVP1ACsLkeZugE421FtsFSN4fHS4CNX3zI6PPmcxDfic/6+Tta0S
uhO8/Ljelgcuo29GtaVgWdfCDrVliXmBvZr1vRsW0R8t7NWdmJoDCR6Ua0OYtxM/
Cx/J6ZQhrpxPwfGsMajFUVw6O2QwtYK7Cv9LruojwthImZKKlO+alx9IKT5HNZwu
j1SyAA+8IEvWTW3KJ2mBstXFg21/r9kmDJwCuT7FLTJ6e/FdM1EEhZMThIvvwGXM
MIPoERCD87AV30f7uYQoUkRpnGAmSFV0oQwzM/aHCNwpABiEBBCTvcQ7BxEe5xJG
60LXEAfNukN46VXWvH2ogHaDpshSZX/GLpm5KlZ0o6PLKrXMEuoRTILcDaFlJ0GC
/vI7HIYHDGwjSIEWCPBjnp5iCD5DZHCe0HhN7K7Bz2nGq612CmWqQNmmmaa+yFCi
zgdOhxFGb9aC4sIIBW2IdyLiq9Jx0ym9Dle565lgpeKcnglQfzzoOCJVIk0Yl+MT
s98ulUUHOnELle/DczCYwIrlhLzIwj2RucBzHoLXv6cBK5+m6AjlJIWukLFeplnq
g1PcBhn7JciBImsA4r8ACBZVHvCD2s6qu5kSXqkj2CziPSKKzO9uvFxxmk4gNQa9
r4I8x5QVX74folUiboCwZ43m4+QwqHtqmn8MKNebCeW2EPIXFueQMIe38ki+ds0e
xdxpgOvQyhUurtpzKDDRjaT0RR2lhx9lO7hstp/OgF2pU+mck50YaTG868vbEnzB
Sr6cL+huIfyrbQO8E0JwrATocbfGljO+EVHufU+spn8fzxX25JNqtLlIbKwGlSgO
VtNDc0micl++HULgDYHHd3JYMktfGZK5oYJD+8AhIC0EhdxUdGgj7ZYzfShlgM0a
nnAfO8QfSgFmsP1TTLbXqApBHy4IQDmqIBjKmiJdXNyszAffvDicdFIe+gVjsWZP
tig2AWf2q7Cw+KA6McuLbzqHIjdUA1wrxDjGPfr+O7p4OqQNiGoxEetlRpLlRvXM
jApXhr5qZ+G18E+75gTAKGkZ1N5CUcyTOKQ8yrnnWF/DgSBOQmJYkvxHEQ3720Z3
taIx3IOIc9nRfuTaYNf+UwXB6zffthO5bM+rp04WMXfdbzuDRsxH8lQXiXzxcZaQ
yshQAl/2Zz0+ybzX2zbx9mOOfQbtaNuQCerd5pAA4ZpxvUCaNxLjdtmS/KvXZ38N
QoL0adbrAJFPC6PoWn0FkqkPJ32IM0Y4Aq8g5pBsbvoZZZJ/OMpDoNGTKK8t+bgk
PvTBjhTIwYYgHcDpVwsdfDiJkRxT3r7HW2rh/am/Y5JYonWOXX3TapfNsORmjuYr
fq+VTcZ35w37Gwys77q91X5OEGvT/7MWm2uUnKGZlXyy85AnMiMvbGFbi5CsB5/R
JxVRMN2ussyx8Ypn2R40x6rBx0YsofQ5+GiJGSSU2VTbUfw5VVbq4P4bA90LHgKx
SCrYCbrBriUmiqy7UdwoDmWa90xXsLaxq0UYkxyX3L7d4Tzni74R7CkExjZWp++p
n9lx6TP3JHQAwiB/BD3RVpak1tZki31jtU9vneW9hhXDq1iEq7rwxMUAKeLRlAKk
bW0+ssQfrlNEGkaFnRtuhAjkHFR74PPlPYRe4XhC13iH5LwKV8rLQD/xngbWaQsd
ceTAvimIAAdD9GdY8QtPbql4RAakV8Ffm6BzPX0oFg2zerfxr/V0l0qEHhIAhyOY
qwe1y6vAEW3I/9tRLbuIw5ZhckBuBDurUBr3UTNEZOpCMSte4SiCAi7qcu4QBPGN
uZMW0gicPgBBmtyq1sgBUX4GFx0U4CIfocx0cXzaMDqbVb7sR6itfpdpWUQX+woV
CV9eAgf44h4REXGTO0XIlQ7Fh46vv2ykDD6SDExjhXPAiB1w2vyo4gkEzx1xJCue
gVhOhI+P4TFoXYR92V33cnLTDqQeTXg8M/rM0WJx++tZ/bsPANev8Jl59Ez1KpZZ
H80WXvjLGLCJRAJR5/fSa/lbr94sDJkf91LhjauMlTjJ1dq6Bk5XQb/dOAzHvmXF
gV1NLcmTPk4soHkRPG2dBJuMbslHjZ3JJ6tQVxJJolctZKmiXz6CDpMjrF2aiEh2
vJJWEl25Eu77SzfK2rCamOh14waZonReX8SaulA1/qc108Rkj+gW2eV77SInoria
uonnAhe3kifNsfsz70Z/vhkLAXKnqFj8LX+AW8IpYc75O/P3nUVxEvlCc8uoht/g
PKopkT1LYSOGXSzE8RMRcFrfRkXC7fYgm2QKLvYCJAVZGEENykQgE6jq4kOJPei0
5/fwvCXAlP+d6h3Jcm9oxjhd/19MPstHL3qKrWcIqRlRGxGlxQ8DMeAa5fcwkoAT
CxssMd1X2BldKwc6Q0fVZEqN58ArggNdhSCwKZPRIhef9IuQnbfUOVJlIAO5jSvG
+RMU/hxWDmRdqMiXxhjZFDX7SdT9e4ArYK7jARYUlgNyOmVbQ8Dht2Zzj/fgO7Hn
O5sz808vnJ2KH9e1pGZgzHCyMd6eFsBkUJjVQMxNC/LJXKXNt6d6ayQDQ8IgclEV
OUKTfWla+TvGk+7fRT8S7PeGvYCFr75skD65AIeX5fqXWIiHwepsfGqj3PGtkWfr
G8K0WTCCbGvjJhEjionnwOg8k3f518PPJ5FzsY2Z84Rz8TZx10Au6kBopQfjJaGI
M4rZlbe7bQmUxPyaSzep+Rb3afiEtx/Bi9pHjblflDKo9AboNu+vvC1uJpBhZDE4
kyqWSORX3p6/N86nGUwTgVXM+CooFWKyvwLLDVFWlbi7Go1vGaPgmdmvyP9qeqcA
t6jusREC1n25oAkzS0WDW3wxAJO/mQuUiukwC2eDfdnmuz58V3NXJuv5WJ04Rshk
urCjFkaaGnGL/cPMWCVq1H0qHS16gpkc+TPtrB0Dj8BSi1WhGBUxh9gTYfZAljuf
cYptn6dv3OCdN+VBu/zPBhzD8rQNBVdClLr7WFBtA5ETvcQgJc633dUsA9WgMCJM
d5esQFIaJ0wfyocejh4VoPSk2f2W4NDS1Aq/HxbZdJzbmNWP+JMAciIRnB07xJqJ
SZVp8U5tRuqQis6vHmw4G2+soLBgcPs/N1a5wW5rxbDs6FcGBqCg0LwJHgUWqEeb
ihk1x2hUzZuRDz2VNdRo0o1VKnWjSMYDguu3CHW4K7XEYIUU1KXaYp+KECBonKu6
VYBBfcxZQ2px9ns+zwiHJiKkG8lJZxrJn71y+M4P+5uxy4nvkTnSDO5gHMrGWsQy
penjVgOgrsVeke66Ujy4QMGrz3mfXWlNl+xHzDfxAt3f2eNorMIbMGzSeXfxh2+Z
r/yG6pUcSAVzQmcg02XJUIwYXeKjtgvh4XUklJFDz1e1Lb8sIAv6ylgD3GzTm/FZ
seJ2gW8Uef1kOpp0Kr+LFJiTov6uKGkmiReYwlXgvjFuwhsy5983EpTEG47815yI
AdWZ8bVBsjkqbN5xIFqgOu/88yRreDEuG4gq/qozWBDm7/orSTVFT6qsbpjcJ+70
kN/tJgbfpUX04xITG7SjZmpiQH16Z3NUTHGoMBpOHtQ8TmjL5zXY1CnVp9gAIjOA
7YBtsNCqc+/IpuTw5C5YM0uIJahXX1X+NdgzUEv9E4F99OtvqDtkNJJo/VU5EOgO
ytL0QZpqHpkTwsqEk+6NRIl4s+ta71LSDZRapuaO29ZiRv9oHcBtviEIEUXjdmHR
lSnXO+9XsEf5OCaKzpRqfm6r72EuRqELyQ1yXQDJVlnbaFUZZn4V3CMjbMYNws+t
iKx8/+70lkrbUtjnAQ9kx51Xzx6F/+w/dMFtiz4L5BkW5ROGurFxebra0qxzqbV+
x7/ZHR+/sQFu2NAndGGLdpmG3X+4lOCnCH7jtVdVGODPRQCkGq5Vzcx2J8bBW2ry
OqghMCl54kQp9oR/1rOlG1ZAjnavdch7ndBiXw3j50WrFc5VK6h1YpCHGbwZX3uC
tGJhbYAQqj4YK7AaKFJlXaRXvAe5u7B0GbYP0yUbrRVFo9YkaaYKoQJYxU8edfWi
j1HfDwqaPHBeOUC/iD0HZDPV7lNitsL6l2mwTOJq+o17vx1I1pER0n3ULxUV/yZn
H0/ztBmxZ9lT6BTnoy+GVjhGgQbmlW7AwEO/A1sH+7URD2/Ir7IVxqVEPltsrEE5
rzbxMHtiFWD35NzzgLrZ8Y+PAjugJJhN0ZYO2085aWKjPkPSJLIzU/ng5gH1UzTO
2/lKuF66++cqSkA+c04UX3FX6AiyfI90b/C3YpU+bNkGbwTPB38KrfbVG/7N0J0G
IfZwfTeI76uSQhMsuBmNEf5uaAoW0v/+hFih6XcJEU16nGE9flr3Aizv4B9AwMXp
lABaLS6cX31n0lbieFJXxj0HB2MYGJB+p2HNeNyuOFPgaHZXy0ZukY3x2ZOohhJ+
E84MfJVcPJv+rNkYoNByASwdB2DTVhr7+KJvFqVg2jOjB4D00jViifi/UDaZsW08
y2W5nMR7Bm4185Mw5lus5Xn/6W3ZmyhfQYqRw2hc90GygeZPj9z37+tKQ0SkLZtq
dsrg+moyeMXHLs1hAvrcXkzKxVLNg+th1QWRz9zlDkHoBljtcdIQdX0wmjVq4jIv
OSDpMgFI5feOf414PeLOm7BgVeCireyMdR3t/NCAQlh53gXg5CjBzrxkN33n2wSU
Ut9pQ1Fp0NIR38QiIhkL9RTcDbKfALnhHITxFfNY2bSnFP3hY47X0yVVM4IEE1Qf
uKDoBJJnQS+j4b/Q9ataYyFJbXch1oXAmGOfVep86gwHU1l8Xaq5UyTQTPdq5O4Z
D9PwLOsB9jaSlEjgLc+8ki1mXOLjE0ma6xLeL6ZcHyav7xgL9IvVabRElB4i0dKX
dm68ZUN/Q+zvpUq0amf9FHRUI6Bm42KG2qC8nMpkahJ5w0qyR14Vr/TegMU+LzaL
kHRtpgVYT1u169j2OnxSxfbAAMxpo2Ace9/3p9dgExqcWMTKm/TK4F0U0IYvUaae
G61F4hPMgnbzgDJN2HvV1YTI+MCYjG126TyUgfQaqKo4m+3YHmKzm4aSjPKoRgDS
UL5ceznwsDa3S7aUjaXfoVkXG/AkxTURtNZp8n3OvBekxPgSmsDjXzGXWJ2tbLgQ
NvkC3/L5ugErsIdczf7Px9ksaf/uiS7vL4/liosC1i7cHFgEgdBWnScZ81loCSHx
aYLgTpCdeVYPghO945wwr182j2JAQwkp06m5lD6ui63TPMTE7Lu/0H2OWRme8k9a
PSe2x6Eguv3gDybMDkduLOMmGEGPTilbdFvIF6cC1TgFPP7FhMtTeE0zLZJFtWYA
5Xdk78hiqo+vVUVtjsfrA5DnaYeeRopqNaIGz/eBJTlNfj9FX4XAa6meSoz0+ftf
A+ZYQkbGrO+qPFPniiS9vFs2aBRom0WzhHxRq2kflHRRSB0vP7Q185DcuSMAJ3zf
CLg5iAaq2dIEEHL2o8ZdgqKb9ImQOlzacSTNwDR7Ap5peFSQ2K13fwiJqCOMCqXR
tJAPO07LN0uEVv74sRxhvIZ1mN3JsadnTNUdKEAt8Ydh8l/0bFGCWB93XOfpt0TP
b9oPr/zQnFN4hI8sl8Q6HfYNhzQs1uEGZFYaAfagxRQkzdatFQh11vRh3tKQr3RY
IrqYWpe4Ey2NtVud8l6xqMlfMSy+JicG9jaoeixPHtz33zqRL9Lg6Jqullr8eOGl
i5YN7xn7XD3gD+qktHVmSyESHjfJ2vK3HFKzm5FSPcOqkS/w6VkFP22EflV4vbrD
QWYz+UOlB9Ht3WBlqsldPiGFTjCNqrAdEsftyQDyPRqmXFfeY5vxPRLoAu+nrabR
T/NTYhGsyQE1WrDx1ePbw9ShJdK5E6OYypYaesQrv/PVxhVSd5wJd4zpaUVBhvXE
pVHU+ZbXncH/X2YEV3ZsxeBWRYcZtKVuPZZJnlav7nLVzD0H/KGN5AgB9Hk+t/L0
pVQYbY0ReUeOboF2y5Rwyy7XClwqlpZRiISC/kuJAsS5+cO64Qs48/ozU+gv6mIt
5MW4afvyu7UmDnsj+jgM5XNT6bB9Xs8vyGzdFdUUf5R77FVjBtdvdZnHbesGeA0T
goOjNoJSFelPVMu/FwgxAQX0GKdof6Ogu3R7AkMWpq9hDJ0rjtMBW4JxEpXQzOYV
U79ctRZWL/wE6fYHZjmtjGmDSjqVLGcQ11c7VXnVCBDMzImx/v6ay7vRfqne7oat
smamVGdoFjhFI9BUr/hu2COgWfnxgia2mw8ODIqTMDQ+jXc5sREDbW+LduRlrJEh
yzMwq4UC8/67cAP+HY2a8JPQNtzSxy8t7Mh476vZscej5/i/lL8Q7jrS85hCkkxK
NRb5c8d08p176GOfkQkAPVFjvJxY6PC8xb0CodP/o8bY2zXQDyUAQbUk/HIh9g5K
MWc58fTePNjVMGxbCMTZ18HKs1gFREYgRxyGb+t3J4JBvMoZcmAzpCdmHTYgn8zQ
Uh4Y8HSN58YNlA0lZIpcKTpV/Z165k5VuRPrkyAmhGX5bgF8NdJJTBJvhW72GMVH
/MhOOESw6B27URUV+X1DFaJjBgdc7k4VfnwHJcgGs6rLA2aw5V7A6NwdM8WFr0Oj
ulEWMWd6GhnKMGpfT/WBuFxF2B0fM44Fpb8s4waazkRNEG8Nc/Wws94WHG1uurqh
94HWLPlj8HJS93ICbqrG/pygj0NCWAFLOuKXI9BlJdYAob2l2PG2u4H84dKlyFwd
TxAJDteJBRybP28nWB5empV4OVRGcv1svoaw3w/ZWAE5XfP7Poj+zLjTomjR6ZiZ
iTiv27mC9SmCT2XXG/j7uGEQjeeSDBcUEosI70780zkzJdZVC4pDX+xoIAH3h4Op
+yhNIi+sZuiTHpCSr/o7ygpiEUJ/yXXBn2T0KFokVEPtqGCO/M7bEgVB4GTIYQVH
8TwpytBKGW7BNmWa2jQnOaiu6uTEBkJjBI986DHtfNI+Lx8k28dHR1KObXjQWaA4
0xa5/CzUX/oJ5x4U2klZTsVGKho81zt5JvzLioyq+t33oW4zj83SSXnn/IjWO0WR
s0J6OE2DQJo8OnRZGzY/4mcBLqknt1fxMKclidslP31+LTl1OCPRnOlN+51/PbyO
iJKShCE98qmRUHH156RRFwDVXYbhJBqbFau+p+sDrdeyNGACiA3asgW4gIbsGBrt
wrcp/6onIm3ftxpp8AIN3LEPi7b+qMq7mD99f+umu5cjcuRtFnkDppRuNza2BjB4
JoZzolon4CCLhy+L/eyix5SYCUjR3NhAxv4ziXqU96aCHsUN0fAfI5KBosweidtU
PhwOYYDMz8+JcwAnPgUdNC+E1lltttjjbyASK6oGtia5ow6G2Z0bE5zlUv+5WS/g
SOpvkSQZE75vf1ZYlBq0UtN6CS90qXKel3p9G4rpiyQhChnXqknEz7f+ObzKYz6N
/L9oTUvjDimK10W4J4Q3G6wO2Wk2bVBewejXUxbxVCtwV4761ZTE8SOsZb6Xzub3
NrvauAaxOkkYUgUohbBPnEY9DcGd2T7/EHQojvk/Cx+/ami+8v6PworIfEebdok5
qCFHm5JjNVOoVfQn0tCHqia5Ie2j+WMNTChuY7Vj2QOq0FUj138/6A/jQKd5H0sF
BpFIaIajtNVYRr2XKxmaGI/MRudMUf+quqbZUe+X24LFH9SlvgKMlWnM4XMVAORB
6OrXP/81QTP1xniVhIKMIE4fUuehi+JlqcssaRLasOERlXi/guF+E7sMVHuFsxzS
/gBl7imF8HSTwEIBky4akrC4xq5RCPB1v/rJHiGQ/Fu2gr/ESj/Y9UXk4DNCoTt5
+zOqBUMpK4rd6IomcAK8+8M2baqLoNd6Fb6yDB0JyrfR/A1gaAQuPiE3OL5SSRkC
g2EDZ97RdlVzkf5/L8LAUdIrvRgTeyAPiww0p3ZJc89AvKdiAeuvE9fSI+ZDJQZA
izSjlmiBm4vqj4UX/qVBqNL9eoK5w0FDQphK/9EEipYkSlXjok2mLC/Bxgwnkz9/
46T5msluYRovy3wDSa/S1KmuEYD4r7JLNH/1RxMgKiX58RSaqOq59CI0hX4wRtIj
TKVFNbi5c+QAR9TrMpz9WIhPDPqHtJOpRQUHJP2PZMIh6AZyqc3IyJEth7/916an
mu8zJpXgjMfasFfSAleSkdjmMuqyGziOXfPVUOR/Paa4omami0c7NBD4lrx3e6FO
E/goVcqIvMpu/PTrDqzdLFL+NYxGtJtrZD54kmAXJts0x0vmyOPvJQZpq9r/Nitp
pujx/IKrbK/Di7rdyKXGiTXU4K932swf1LdSsy20jyrxR/jryCtIBFbBJv1FXgPy
bZkWP4uCfdDNYRxnJdpCEYuWMLIQsY23oLfcHLWU+7CEKR9nOXkNnot6zT/nQIna
K2NIht7wSZZ+e1bAaege1NU+rJWqONBU8wCqi/8R8St/eWZpWsDVObqGtWZC5LxB
/ZHiBNKrFLk/IZromccN3WQDgTN6MSnR2gS5LLFExC/a6pOeFVoQpF/srksnc3hZ
6xfTXRWV4M71XzmBOknVQTcG3ZVuTcrJLHU8lp9pxwLFy1xGkjpwYsXEVyVZyq6o
lJc/8h89606/yZaa2dw45PdPSGmjqj1LHQnQu/hjaNcLdTfCrHPzJkclHV9OtfcU
9H5jYbrpW6sZu8hFU7r5gWZPmUtgpRp4GRoPvOvGJlDKDy7Ojk0SVhruEvcrdQYW
SquS8EXKm3oCGgBI63Q/SRX2Fo56cj8q1O1ZBCYqFSZNpIDRZjeavAfiEkJiJqvw
UePUPXYUrSMk1ps+Nf5LeH7PbV7xMo7E+FT6vIyN1b6Rvt7bg/gZQfHg5caXYwS2
UMdMrwuqg0kQOvWFYEN1QK8hk1gDUsK3V/8lFbRvEsD1mUnVMv7ixjNx5NEvxaZt
JDCfgGXHON492r1K4I3U9EzNtNGw2iWoVxD/Id8H/AEiusk9GiZCqioUGMfKpg9W
Iv+l/jA/kFX5IuDHPrc4FRvhqc9cXN9um8xxvFKLs5N0lL77ebjfGXdZCC3RmrZM
mdwxro3M7teMuna52kOFpw75mvh6krCqSvNGE99cd18ZyEJHpzSNIhEvL5AzALeK
ctpLigD3VXWRUa5322JDgjW9KrLrUSlYlYkKuRDmlepBcBDeSJGZmTWWJSBKluh4
Y3BZ950KrYYIAoHTWcpn7ve6PEkGFYj0LPG2m3XYJNM32JviOjWeOdOGLtatmlLV
BtBXal9QTlzJ0BZJ4+j4dr/QZnkKeaMRgd329T39v7JnKWmaAjhqq41Q3e8T3wpf
fZLZ/vkOtTTpBqwkrcjOJoZ2K+9Xc+uBGkD5uAn2mXPn3jRUQgMNwh0wlhZUUiVS
9WvHazP2lJRxCrr6sXpIhB3AFAm1+zwYgOq2XIpFXR+e1YoIMr7qljsNWEF88XG6
xQ+zdVkj9NDcvsIHlVO0N7fz1XUTRw5arQ29hDNG9MJ8H5y0CLEsOVhGXYKEMCeN
73ZV1W0Au+Cj45BueJ5RMEUjw3dhXWRs5Cej0ogkROUAdT0oBlvkKpHhUrMODnuD
zm8h+rX1nIwiyktkgMEYj/hkJlcNwvHqxmYQEKpUZM4/Dioe8FCLd9xYUp8hNUET
ctaDdJLJCeyRb7ZYt9TMQdhsteKwy1tt59jSBeqjYWQEL8tYse7FZcHpJitbXmvu
Q3G/oHKAg0CYQ51maO7no+zpCSj/AWAIhR88jGs9FGJPNryowYOxUKBNI9kRv91b
yA7a1TikTaR2LMGKI5BGWUOp7cYSfEwEhMBhjyquRVFT6LsJL/rj5D9ZRsxVT8w/
Nliz7oIUSc/OMSrT4aJjeIDUQsdOGd+P3PJ1Wz9s1s4RH3k9vkrTMUdLfBzIVeB1
RPt9a6Kx91en5zcZuIs4dTm8Gpoc5FHUWt2dbePBYbpzwlLz6hQifDRo5Fo6fOLq
2b5XEvtlMmJsnppiEWthFJoircoDJa5bGyptx0rRyJZ0Uiz5YFD9o0s3rJj9zKVA
bs3JHEi2Oqh2YRaSNMgSDNsEoVye7jYe7DatPw6JGj6Tff3+FyH/Ztmrc3ZIn9Hc
JHEFUEJ8tDjlSyeBo05aVm7v21VxWdIIYkFzjpspJdWmzQr2DMIngdJyiCFIbBRq
IIDVBjVCw6U1tv8dgREw7J+/omeS610wH5qoP+onvM51XCwzZroATxzngFie6CAs
Pwcqx9eoeTDhl19JZyd75CW+HLw/FAC56VcS7Z+SOcHJA79q7rCnPJyNVcBcmkSP
ReAT6ahDe7CeyKZ9xUKp2MG9/1B6DP7hCdSjicuV5NLjI3zBSX9rmyo44GyDZqvo
XY3WAggnXSreS9tEen6n6UZLGMeECpSSEszlmkU4GZh6RefLhgNIvqrTG1dvT0i+
a2kK3sLvJ7Kyna2akGnr0nGq7nysNeRkOpsOjSlXf1oiW4GSKV6KcLm+lNdDTpY5
DwQ5K2WsPk6rSLOSwfQoDLTlAmV5gkEdPwBgYOqmQ0bsOK4nencwcNlbY4G1H3U1
KFQ9KKxRLGxQbq96YBg4P1cfms21XRut2ginV1gcV78/Onxt3WM+EFKS8ctJl1hi
KnXZtuypgHTfc4G8lS9vFSR7JhcmKh7pYPlSgWKWNJdt3/w7RlfYi65WL3nvsZ9R
nSVYTwt5giiiUf57mwm4F4D3pAHZEiUAjoDMAdDmmy82ITNTEZndDnGyiWtWO0IE
Mbo3YAjIrrQ/b97eO6RWB7L+LNIiCNlGLQNYksMZAp/xLW1sGMoBCwmp/lfsHnMD
GeywjDnag3LgDuRaf0BCS3t2WY0oujmbuWBy74L6mK0XfcS762iiNnTAPp4Wyx+A
xIZi7JeMGBSDf0UMh+tXHt/NI0NMFr4OvqljaOah6gpIvPudBg9d3cJuPAQdj434
9/Edebss0f58gMD1QxPRCODXNVng2p9AfcmO/tAa/b3oq94tomYWzoFHHq0W1+7E
iZQTAbtqJ08YIK2ck+elWcZXNYq5b4E3UzrswELyAUtfY6YyVDOVL6UBViE72L9t
ENXXTcW8KIEfJwJSRv3PK5yCoiQooVtQL+O++kiK17xbYEkrPZe0/iKNS5G9z7PV
/s4oNbPSgSJJ1TXvk9WvqZAmhKkvAiikgBVi0mF4r+gkmS59S4+1yelf8kJzimx1
B6MYKVCABNcnEhVFuLIFlrTKhGr/rXj3aLeliuMP79JEYdI/xYKoUqJ+uI/WG9od
W4WQSGCp3XPiuuLU61VxfmEKff+LCuLk4CfgvZXf9qj98H7ET+K5xGKuEupOeSoe
71BWzH5WzVROJhAoMY9QWeO3wOkLuW4bVhE3JXWMqWbk+CYQeHQJoMi+h4Y1QTsf
lNTGw61105Iw6Wovpx3Bidqs4lOAYx9VEn4InDw8SPpwpPqLxL39FkpTaQCf3y6a
vMkUkMyBmlM0P5Pn2jrFNNUbevzBFIkdH6kDUanzKq1wde6f0+0U6ZtzVr2xb8QC
WQknDCcvZlXvh1pKqDeuUXAJsDHzbkNU8Ee2DUXClZxXFhgvd6wspefki9vxhIzI
baH3Rvz2C4QIJZq7027m7gjM+4vrYFvb7EmXCmt6ij0Bz0PfdEmNHzi71yLMJ8tL
BRR/o2TwOheOS1LZ2+vWW5o0VnPRzXewey5EUitZNJB83MJ+TYITYGAnBy5GLFI5
7lWzWISbMfCgM9hX6gasMKVZKbbnuhSIjOxWQkQeu/WTOuZJF+dAniR5/tSzt7nV
oTwWy844pNqJ0lDtn9kIox/dFcH05xod4OymKUW1yV22SdXSieP2n3jLyFy6BoZ3
Ehm7Elk3gAA72PjprncuDDkAuA690Y3ArFdMpZ4naTxpJMFtYRJSz8iTHEHxLM8D
1GEeYv784UXnMUI7zNQuXuaGrhuWtgZ88nZ869qDxJQNwRZySp0KcwObFi4CS/Zu
Rwj61ikuSUOWGxxBMq9zOdQq00KpR8Asowt3IzQrzvHq8EmSKbOd234LkZkZx+z/
OqzxCEm1Jpsgjf+gVqeCeRYy+uizm0G7PNvzo4owIEf1nmtfDj3ZVTsEfovDmJQl
OlVqDDkGf1DKJ9z6mmL3ll2wljpCQIpebmQFh9mRvAiPOxkk48K8RzKz3weUmxfZ
X1GuJ7wXgG5JFDi+7jbD9xaVFTvLGl4npfh+CaR0BxwJk5Iwy490MwBZGguYSjPb
HOt0/k3jgPfqGaYjAGxWMtNlb/LoSGvLM8xMQmIvx38ch3QC/kq/x9VpS69sYVFi
oBsGpYkY8mdIrLiOj4pqjjVbPCiHh3x7j22ZZica6W1rEgBsfB8V6xNgR6Wb6ETW
8ft0JBcR84kbKcoqS0hla6SqhjqRPAmTDYSnORadgTJPXHLvF4Al6JwlORZQwenD
MsAcBE6O6JcBYecuiFFWH3Buq38cYKva/vfBSnD9FT9xwg50H74kyA6Suh/qsIZi
JGvqRQlvloIbpsGXhnUbE8FdVW6CLlrMigdYpDM4bOScJXpGl8UX/PMhY7UqNFnt
xO2VhFa11NHxna/TKD76/WgV2Kf/gDDdI8mJ7EVzvAhum9IlYo52d+0hHwvEKhTX
V9U7FA2PhXVNf5nxyrxnmx+n44t66mICKv2AUgR4YpkxH/8wvsh9HuOpa4V4Sgo8
wWNGJ1ssWIkzHemXHmtOUFs4U6d08jPO7EzLylRfHmUeDqFSWkwSztxjsxoCOBS1
bybW7hsBGsCeAYWg2zNFmvZaHh4pz8XFVOeRxEMk+vw7/RDqKrExST/rKg7BkH+j
D3c4ebFUq8vCrfIyxRIrYhtMRP5X1jKV5zkcSodVMFz9RNkmvV6VNGf6uyW6cNSS
e4NYvbzKTMwoZ2WUO3u8kvr1r0vVWiRClRaJpjqT+/I3hkV0/YwNgwZtmDbkQQtI
nUhTaNLb8oo+ZsNMhgETuLYCv3iDM0ojPMXSZUO20DRlqEuY5tobdVY1mK9zaojU
ggkm8SjWCB+N6abtZZz0fR5ox75uDux1aKvP5lWsnXOwP5vK7LVroe/cc8oix5Zp
RN0BrwZuSAMTdAMoMB81IJ77Meu2HxOUMlHf0ORXAYnNPG27kACpxgrpX+CPYzta
wuXNzUWo1d0cHgUiVIlUnD0O6Nlu9IqCqJH8Mnbhptd/Yruuc/Tzh0ub1iOH6tNh
seNVTMEu6PGy/JW2YgYtz0OCY15oqvGTHnpTwFo2LCiwLMU2TzGCSsmUJJTq51Pg
bCVUW8JAFWroljNJY0hEp4+KnKBH8n8uKLObCKIsvs6V5+hDTb/X7HN4xcWughIv
FT2bP7Lx1KmI4cn81rQVJlLEtx47a3idYRZlnucUuSJg90SboLKJkCzuwbN2k8uZ
lfELU7GUbTnctmI7Njr803vdd0Glo/uvcw81ZU6S9106EQ5d/rP2PGB+w2mQZIcI
sgTakc8IMaPWDFl6GTmvSF2oysDCfnZV+fK9phoUT+rkzNjBa7Pzto1UEWYdx9PC
QKizk9lT8iKHeOJHPJiqyaGVLQXSCQW70Rg7xndB58oShqNtu1gVMIiy75/8W5nz
h5pCUq2zk7VE9Y4wsibWpowK6xxeDPzfXG8/ez1pM4TlYU/XVFKwbYsP3TLZRPCb
dYl/4TxYYGyRbBizUWhurz9xraBRk/Rg0mjyKydYjntCbCmMxeRvEklwm//tLtqW
PMV7MsSWCt9ih/f+T3g2aTzPjIR3CLwyiDMfRHPX+MNeyjxkQkfLzn9LHe6ZuKLb
geV4gzk2QXXTtaMdxERZbK0PBno3tBjSCqfB/y8nHaH+GZ6jLDl4jxpclxV3UOtt
gQRbKYVwOh+FrkhGLdCSNhTqGjOs9D4Mbg2RpXPMzJrH5Fxf4dplaMRLC51RBYva
98Eo7fU1h1JbMwlu4b2B06pzeCR9IXbwJI24NtMoPm72IJiHiscu+0hU+VYRJR1Q
i+VOIOcAmpI6hbc6gmDyiEkenlcsG5q0F9UPorT8AmZXqaUPpUuBm9W0veHT4Del
QluegmOfie/mw2FeGwYli2vTaGRhLZl0NJ/f5NPgB5hSD7WKobhgqZbvrDM4bJwb
ZVISOqjx1pctqXiMvigXbARDM7nPns2wcr/oqb9m9EZrRpyMUUZm+K8Fwj/ijuES
pHhoMUd4yutXv2zwka+4jJ1xMHUU4Ohh/t1LJ8eRa1rFkW85uL1MvYI1GgLT2Oaf
WFNHc+CfyljM5cMRo9wslA2NjJF/kvs9j9GSG7aUcLtcZNlmryLL+rUXjtDH+WdG
0OhfHSupkwYVKZ+BiLPwmi+2jD/1J8G3Oj3pJI+j0IWhT0ARFO9T8iQNTLHJGS1S
CIupt2TLIdy2bmp85dMtTCankzdSQj2OPnOdazkzC8HUQ5tTFVXSkdbHuSTmsYVc
FCoiAPbP8qKrZ8rhpSycihsF4tMUhO909ZNKRdYZXPi9CmgucDv/E0Dft73N9F01
ECMjelU3W0YDJsLzaqv1cvkxrkRldzYPwGf2CdahkEyTK9ioKzoJS6KKPFYkDpNU
12h9V9CwKoQjr6H3bjjzIArP+6CRGF9636thq+BwPnNoLBiwP0ybNPQPP+JTDoU4
ieq+2cgTdjbTtqwicmHjQ7woouqX3LpA19XmKFTg8lIdDNJp/+DzMPzRXVt+uxi+
hUucScxXf/syhelNrJKwrfF+yzwtqQ66iMynkm6OmxtqgeoNqfxaoa4JSiZF/17Z
u28Hmhre63XCQrasyjI9CLqLAKYg3PHoqYaobjgEvjSHYdUdW5NoycE0JKQ6m4iL
xHtlzIBnSPm0VoEjs428UNrfTkev6MYzN6mKUoS9tSb1p+qU9HLmERyqtu1ptWP9
5nCva8XZkOjz9pBVB50vDsTly6p6meIKTv5goqk6xzOENkXWqBHIOmRl4JYOsLg/
7Rc2qfTGoZxtWPVHZQ15Qqi/jI9f57eqWRR2g7xtuqsYCsx1WoVH0TTqrnOutUT8
DkLOVwwLJEgPatF8KtxXfVKHDaSAuw9/rYDZfXs19mmMJvg+pDBWdJ2VMjAZySd4
9C2JD0XhSy9FDKpH7LLeOUKp1AANQDyHTQk0w54o3h4F4UojHGuuq46NTmjKNEwk
THmrvK6DxdI3W6oivbbCSQS2Nf+G4iY0Mj0jdNRFzvlmcNyJGyLchI0aWVFGfFct
dJbnvtFwVw3eK8Gqk0HrmakD/77RXjDzlqzFFLdnIcz/hyOR7ls95eAC86lhA7cH
JW1MU8NkvbPF/dqgUkL5IlPYUbub4k6UNrxfLW9kLsxzg6CbChO8BqoaqHHa5BLG
CjJQo9Zt6csLzFtRdf+Ptkfs5f6BTCTHw2dp2Q6fhae6yVsYd7W4U5nzjvNpo4q5
oVe64UyH7FRwcmaz0D3QAH8DvNT/dKnoBpUSbR4I11dlhmpRh4ziX38b5Z/WlbH1
zuIKJfftkiHNXOHKB7X8oPD9WwgOAvlmOGCDWvfuVx/BKiF2H3sWGLsjxALhETS2
ftT1L8Bt4goUmH5rsIS+VFlJm2+qyge+6fLfI5C1pEFXE/033tE8GlN5rdVr7uuq
Hc8INuVb7/rDioLYOttuJFhgYvckmwkNV730oNnzcw4HdwIIQkjSmhkX1JNUxUYU
H2TZXxQiY44AwZM8oze9ifbfKCocTr+h5d9bMQIYGNpD8sDCi7vUR0S1T9Mdvxg/
R9bzIoQmB0mg9fFXFAXghH/ZZqkMWBDfbtWd8w0RABzs99mAmspjQr2Klh6gu3pM
jJtRKBxC2IY6cuiVydYSndELgapp4UHTjrGq/G+60IR9Yl6RkUNnJEaoQ2kvb7Uy
DnlISBRsQzv8PIxyylsy37EDssn1g/rHqFWK5gHJ13h/Xy79KfOwHn2rE+fJSsji
rDw6SwOsNs06UkTL9TV3g8NkemmSA5JmB4g5kNsKC5LXnqiKyw8CvRpxLw/aDRrP
+Wji61ESUgpN13tCOS/eiW9yyRryGurAhpAYweIkAaOSI9HE1IrTmgA+Q6wc7u4c
0CC0q3uogPmf0n9jljif3GZuCf58b+rlEpuqFBUXwBA8mrTIZ9PvWSlMLXcmYnph
tNOn+9+pO0RUOPbXsApNNWtqWzFG9DL2f2PJHMlIb8TYHKYgBZYY0dxhEoxpHce5
n0/EVea254cngUrg6UnZSZk62O/Vq2h26IrDIHnz/rcYgBFscGv0FZTLVL/slpZU
Om35495MeZDUlNGkBKhxc6o86M7T2KnceBoW1aTWQhZmBroEvi5T3sjatxVw5+fW
rI7q0j91nE790GZzrWjxblaYpxldeXOseDaT2vY6LjT3hPMIBUHIMymBMqy0eOMs
D01aQSHwtJJ6gt4On8pdaMFXypgL9yP8MGSBSgzBEx+kBFF1BlAvHkPXSfYHfwkB
M8WQ++wlGyF7MhUHsObtxXfasYdLTIHgBHbfns27UyEWYtaljah6DKcpSbJhqcwN
g7g7FPcVHVGvoBh5+lqILzm9SulX41lrZPYxMx7tonbSpoHu5s0VSOUtEmY8cMgk
0fNouK1gHP4htkCpSgvih0pDS/0Gsc0vE8LG0Mdbh28qws7SJmWuMJfXYVvnFELg
W86HlX2p57w6qI5l6G4VlLdvJcrozH6Mm3F1AKmmrKonMWgeDnRcT/SWPdaB7cwd
JnHLu3ZTr7ZyWuR4rRkO2un0dufqp4P6tXnJRIOcHK870L0DTTCmEhAXK4z8/G2A
IwJ/S9Rxu9nC2PF0Lgmz01R8NGiLZAjO9BUQ2I2i4vmy2f4VORLMKbT/14vbNHKN
NCgL6IOYqSwRnL8EO8O79G5p+dRZCzeHSO86tqD3l/q9Ggws0qdAt2JAHSeW3CBT
/A6JA32pD2N2c+Xweh3LotslsKxH4IEBb80ywxrnA+zC1UmvrQujapo8rPkeqh3O
4NKX91vkKgwal0fIvSHJMbcysJyC7XRN1OZUErhiuC6EkVoQLmN8one/GTz7iHfx
HZisOiNzNlHA1MLOpdh3hNLMPLxhIZ1G12D0U74v9P/jlN4LOeS7ui/OJfhDfdyu
yAKtdQf2G2gyzCd/FZIbHL6ZF09sIkL4ZNpul4mig9h3d5WYzTaO5EoLkhSMKwqR
JU6kIgvESyeFFtj6hf8DzKjFRayTfEYzp3Cm1p23I7RLEtSqjR4j42kEOTY4WKBd
dcOMATlAfVC8NE1w0am1lwjkkhrHlTwXSp0efZeOT07Y5eeUsXxoNNbCClJ63uty
vikkpo/HNm8rSO+rba1z6CuwTNGTgQlLBkuhWlO9A9tkpd3PZiPpNwYYBKj0tD5j
bhDGNz8mMgizGB6+UhVbAx/FrrvZH3DWzSQRQSJWjHIHXbm3kmqdS7h7Y/Ekuk3T
Jc7TYiXc/V0LsRElhci8+fFlzto+b3nCKRbqnujK9p/cFAh8iULmwaXfkNHo3/HN
QgNo/JoqQcitzx4WbbnNZQXIUrZ6Gf4K8OY6acKxZaXoX5xhrEfW19+1l3L35jh0
K3A2kzqp4aHQu0C20ytqjE8NPne1oSEe+pWthK/oDygg60JPmBciqHc9woEVs/F1
eh2lXxGkS0tbLYbJZbB3OShKnUDp/hk9/a7d7/rhu1IYxgTiQJOtCM+lUKI1RZUD
VYmLdQogCxj7mqnUj8e/eE98glBl+3wlZMCplDunaAkBBCn37jklx/7/OQu10rLt
nTwcWQDFwsJbDHuC06WKL2nOOb+YZtVIwOoCF2v2VoQ6COpCaqUV5Mv3eMXxPul1
daCLj6EJ79TeKSkDacP4lqGICUtinvki4z6JV8Z/exPlsLUTk8fzGzd+tpIBahQP
udLoYXTqH3eBnLRJyFBTedd6p0m8JDEX6/1g+OTb98rl3M0P1i3rJIITwg7iEfAW
h5GRcDzzoP2AGEyrxerJF6F75PA6Bxn7hzymD2MsiAx7qcRd96ghczRG+rdx+Cc2
0tTrP6yxNhgywDotB7ZXLNePFqdorluK2h5QkLoMEeaa5gpIBS8wPqSxWC+NRaI9
9Mr0p7eeH354E3MRcatO92N0a5aIExV33Wt1tFpcMlXofwZUkzpFnArj3s2LH9Ig
6uYyO33wr+FzknRiKAnurVFHhAGmlVtmEG5ZNoygcPFV1z3qqUQrjOOJLha+m5FJ
OWCWlJpGdc79GD7xtx7Hjk44SgV+43Shb4aYGSJ9DI6g/3ezKdrvm5ZnOzZm/ENh
AXzEluAEg/pN6qhR2CRtetlsMab9hjWJVWO3Xmkx5qK0ONYwvcCViPxpwpv+/enW
/dfQQknMhdOCQZtzTywIOPc5O7qDgXnsyAKYajY4KS1jQvZxXEX+7WpC6/2/1di1
G2NPeOliJ2Z40KZWmNo08awkh1Xol6gGP90rhGwCFYQyhe7mmPd6+WzxRkF74+tp
Fs8tam+/ifxDk9OCiUEheisLoC23RmUf4bU9FUfIsBElhIFUTVshuDzoGvlRw4pw
25+CNFCPktLiplWHvfHMJmjaS8KfMGksz0XlkG2nxpd+rYwIjigkucZCyGInoRH3
LasVpVdHTvDCtYBkXonRyQGk3Z2/b9HNv9Ey2LVGz474CbKbQHx56UMGnyLgcSrJ
Cp37GQkVH0UC9lk/hh+ZundKmlT11PxBVTS8chzdwvT3F/J82MX4iXctgQqRKhpJ
Ej7Wl1Sh4oWMitsOAklZtqrVradHnrSDDvo26Huv66ILmvhT+ngvGueZHjR8zzGJ
IP4jTmMtXPlW4vYQpL/JaxQDcxHt4Np3M7KJc5uFAZoYX0Wj6DmyrvUTEwJCGEoM
NgVa8n3PGhfDqDKwU73aY4+NbllrzFx+yQ/VdDBy8kwON1orYnwiFt69ahroMU8t
cAo7uvc3wapEHtoZ6sfolXqKJ0wOdVgP7Dlbg6SF1UV1gVDLAIN9TqMqZtBsUvT/
nrtlkOJ7PXw8mNoYdvoeDcBRt3ClgXdaaD9W3s1khJ/azmjE7+ryCZlSWHOgC4p4
w4Nc9pmjYn571LAXSONiuK1WbQXXdeNV8S9cezkQrwdKKpMc8yIZk8SLJwcLpvYa
mS2kvs6pzvx3M5Ozda9WK+9KDkcE+n8Qn3KUUYvViFHLdxuVikO45X5QYjybouy4
rpu7ahLSEbugR9wpn3HS5dvQLJfe0E8nAu0LBYP/SPoUxBqZBZZEa6abJNOrJfWX
ZLQfT0TNKdBOdRFVkoEvDJb3tpUoMHv/cH6Vo1xC6HjS2i7JDFPMkaotnN+3VMmr
gMj+S8wCaRS3MI0O1vJ02DJO4GAmIGwg7OKjJPUmDqPLweZVy2VyU1BtlwmjrxW5
SbNGPj1yCoytt74d4ldnrc9bP0oxoC0kvjQBx80jX94Zo1nN7d0JmcjGnwHgHlmY
CC0WP7j7HGORmq0+9YsZQJERCjZ9RlTiUr5FRWqcSHjRZLd9ML6aEm2MFjpomjhn
IIrJOPLszCRtzbWxIt01twY/eDKZ0vV2IufLH/qGgsNwVqH/KHT+5r42nJIpfnuy
2TV20RyuF46ONz+ei6ML9gcfMl5jn0aTlRAjUaTkRR3PLrgy+8nS8zTb4kxD2VBa
JwOluXjLIAwpa1vw3x487iwPBspLoK6qnMZjZdMwx/uPlxxBV3FdPh4hvbGg2pU8
9GayZ1xZX6V74TTZzmDxfylBcXkEaOnf49kH9q+XiNdAsI4FGSDxKU7Ul8FpG4Ap
Aehl2ImOFLzeZXAeg7dT8uSZF0W/3l0J8NVqig7fyF1b/norOHC8js+ROxRIgdbJ
+SbSuuemvzh9CqH1WX5+FefJP7aHqZlq4ploINGwnFaZDIeMf5HLTmdQYDYzAJ1C
K/RxYH1gLcrNQ+FbAb38SbNww8k0yWf4TL4x39P8miBDtbIn7VVUmbnEMM2ze4sN
yro4V1WSyHRuY3RSFLDE+kQ6F0b/LUREpCpJnUMsh8MzppGU/TjZ4aLsYmE+6JBD
4nbAelbPEgmScfztpqVih7UlB22tbSQOZF6RQwK6YQdMscuU+yTc2LEtEySxhtZM
g0NyJ1sH7MxjKeBhMWTU4gi6/inXQzoAxgZa8uMWg4I+ppqP8eArplovC4A7lXy/
Pkx0wWlyvihUtnk2p+HXkbKJ+0e7rqjPZ4sNXQ3XoIAcAHUsh1hoE7g9CUI24w76
0kpWfxmqfPc+B6vuk+l8bISpoFPGV8QI9GAOjvxoYdcH6SrwMl9bHHUD5L/nyxza
ZqHYhZrLJ4VsBIWQwwdbU2tVbeeVyCa4JA3p8f3APRHefmIfIAkeyt0re38yOYq9
jUHiODY73h0I/dLCzOaxTrVW+3rIR1RvTs/+AjlvYL2HMggtUE7FCJtr123QsrM2
2XgKTe1ZI6hIpiyKdpL0dBZznrLyqSXzG+HO74MXkwiboSklA2b4RyOFrFp8h3lQ
2chgQXR8MmIpDPMKWTywInn9/OU0NjjhcBrOl8ODzMN41gRbDzqgIRw4p/RLNO6U
jZwOBUEP1sOJ4vyTDNIxp35huNdtToJ2KKmr6iOl4ucwJaKI/FOeh1IzPwsaJ6UF
8LA1mZ6oSlzw3x9uDIPRzGlWAMtfBE8Dn2dp0kYmuVgsLwM5RVSpAeOptGEbXC4M
cQVAy8CXaWPHLThBpyAPF7HWHdHsiNUpH1fC91/c74ebO3aD+v34viEIuwLvRLoO
sl9/A/FhGFxmmtNEh5L2gqYkiewDuxZUYlv+sZgmPZYaTHukKwJdXInG3Ym0MPW9
pJ4QewUAtwksSuvYcZDa4DP6kp5p1/dHZV0zcvES0Smo3FzXdracwAyu7snA9xIl
coeSh3rcxVfpaqMvEu8JZwU7fcZ4UsyUYk07fDmGUmKaiS4zFWQUjZ6ehseScnmc
wQwvrxRLNcdg2rm0QdLzmoJsv2dPU4KjwkI00LzrSGtJvprxkwQ5xnqiDBZXXupE
4NIneaIm4vLBB6csXkqspb2jMzIpEEWvI2AtSZ10IzduMbRKK/6aPM+bP3P+hpTu
sXRJpuXQIF6UcCfvyQWbn0eo0x3GQ2KQrxnrruvmQ/DLfyLF6aMMgsO0zrRX+adY
HPAtsWIeUBVofJ7zsWz3CmlcqE8AWtUvh2uLfqh0VK8J+sgarTmz9TdYexpbaRs6
Qc1FLLH82+sCPqYRyMU5VyL57YnUjcOKsPb4JD9dAAX0Mtuh6MFEMa1u+HcPsstB
Cl4do8K5hSdrwQeEdykd6CQrB1AghsNjtIe3yqmlWpR+hf/aWrKh/dIGZtWtZMzP
/oRz6KRCHfJnVyiFHUNM07AoFshrZ2eArcXBFZnEFjPe5Vg26cA2G0ZXRjN8T3Ya
RkP/if6ptl19zdzoMe7ttoC4hY/7nZUEWZ9MIAR79d17D4F8MdUqWOq1KDL3P1kl
hM0edHW93dVYkUVZVciotls4I1Sxosc2XTV8joTVGeVnhfx5fNFGsn9k1Xm12ram
45lvXPQbomBh/x6cm02PPK1OTBT909OOX4l9GgeOBxWkTMVBSaHU1Lqz5P1eXD0p
fh65nRJMGXU4sE2ZYJx6+J0p3SjCNFwGfebCXseFmlk+gNBY3dZZ6n/gGxZq4oaa
eqB2JF+QRt+LTL+QLgyk5fqG1OOS2IAflUsahSmGUU851V4FxX4OQJkvvn40X0Ep
M26iykci5Kf57IpfETHOe15aHTxcIquo/JXWnPN6Nr3jE0CvkW4mEBpgPbQayhT7
086i1heL37e7rE/1+pKO2buLQwI7R4t9+hW5hsqdhYoVTvPH8lgQ/P1prvPCE5D3
n/L1P9HGZ4YM3+NV4XU5g6zf+jp4t/pi6VO3qKdcAdzE4h3t1KDyUoZazkntDRPO
W762wFAgCZlnncb4EXtYJl/bUyd7tvfcmk8L+NjPAX9dhMa6BWvWXD49QZDGKaEJ
HIiP9u03a9w335O6rJoSliGJg958RHGJFXxuqk8dZD1euWBIG+jdPBUmbCJR08o8
I4oPl5+LXjNBEaBGDgXBfnKM9AIBVrTPvgraryY1LTb3ZnDx12UWqio8G2dzxfTO
0IUf9lsTSI4pCHVkTb4ri/GaZzX3riM3GuaA1SD1rbkuWejH0H4x9nsld1gYWTqj
qlOlvW1CuRhYfc1JIdGzA8gO5KowufysGZuKg+B4CmS6g6tyEsaHOjl2StrLycOL
xHrU3DbB2PEXfyPHGgnFZSszCx6ONMJpIQA0+vLwXzWcE+Yu/ym2HjvbreJmpeyx
TF9FQoDcqqxXPcD22d+3CItHD/k7c7WR69CewV3C2HyKIW2HXITgvMNIIK0DOfMJ
vdAAF8FrR9bzDfYdBigee/geNJIBAtoVecFEjUOn1WTVQOT0tZ4rYYyYYGOYjEDe
NNQNrM7AgVndmW6Uhu/ev/rRdrH63XAFVNpXGdHBiDtoQiRgzstS9cUzALnluSoT
UQhV8raQbFRGMJC59AzTKNBsguMp/LDywQwA8up0rX1g7GUo1tFpAq+9Fwp5HPni
cQRRTOrflTM4M42+q2NEyMWNif88VtWO0gXXeQMxoypMRnW6h+L6iU/LBq/RFlA7
/y6EJ5zjLuun2D98yt0m2ROKrH85k5vy8jqbjsnPERRLmystBZlZseG0zFkSRIGX
9Qow9q0FhRtQwJs4na+bw1C6be1ClueFK2zkEduDUwTQFMRTLq/+dac6sRlscSIY
loe42ksD70k8eRYa50GoyVNMbp7oP15VqXe5WAO81j4uHFZKLWassGp6YvwOUZiA
/QYi46U5sQmv42dPHwtvDEm2MjWW1WwcbVJ6yyx8wkxPyXt5ZG0LEWO0XU18Q374
EVmRnGvGsY/Mn7KJ/MWTCK39naYW8l1f9BtPV9RM2b4cxWVHjoC9LVdNmdHqTiMc
psmdKQVwHtBGXth/MpE7Z6yr9ek1PncgryWONiZ19oh89/bmOw19plYZXkxjzstb
4At19aSaXsvTWNyxAqUI5S93NnLTm3FyhIUpxaJBu+OuhqjQbAcOLgryrrNAxIpZ
7oM+8fYaVg2taWlNxU3hQkvLu7eFzVO3HElq9Puifsi6+r8r2xhQ3UIavbDJDK7+
UQeJzoGVkYFgDATHzC2YUvS752ANTSOuyiU9Gley7g7ug04XkORB4bXn38rX03/P
yb0akuSdws5h91aBU1C0hIOtJtXU0oWSl9XmyArznOuFsZyk86/MAIlzcnfilY74
8tqRqICp3XH3/bSXWHc75Oj37Do3QzArlKNP/LH5sESYp71ufR+enDqKml+8RHtM
WZGTp7zJQE/vsAJYmCr2ubvUVqCyMH2n+6swxol0onyXLoMd79jK/wZxxuN5nL7D
10M9E2LpF48ajH2RUTh05Ne9cLkSfjcgt2fzA8FCeh0i6bXisGKXG3ZFH7kior2u
8kAJV4QlZ2CHSlj4TvyXgKVmshImh97VyyBZKTfZ53LAFo3SvdgwFTBkVWV+ei5R
4P4N/i5r/+ENVytJBSZZdYyLzgrPo6tL46jUnc9XxtbBK2DkUwuMQ2mOhRfP454Q
rKz2WUh0SYRX/gpGrjwraw7E0v28Y3Z5UTK/zxx+Ri2cAlCHzqxT7ttSUBOyHI1/
mso1u5Cx3ARRHcfTQBS15G1HWEsrtDJmECQ9P9wNTDJU5y9Yp/VC4BuFHdEYnH2w
lV7pwY7XfZxrDC085iA+AwT+JcV5HaRp5TXcHSE3BV13aX7NoRveGAlC67ADDVb/
pVfV9nQOf7LsY5+ehKtS424LtePZnFlfQyd7WV62e2tKY3U+BmxV9EseRQzcxspn
8qhq94WBWXCaDO1C57wawSiu1n7iH5LE1PhQY011vetAcsAsLa8uuhpbZQieQgZo
ZqN9V9C4m1viqgEXrta0UOaVEXjkpKryRd4Dkgtck0k6q4KhzbtLsY4bNlQQH5Ti
tAUnaGlWUdSOdcqxyn0wECVhO4x86SepPT8mRNn66He+mnDsk9xx+LNyqIcbPvLK
SU1STOXkdXUbnpyrJDxnhNiy7YH/tXL/jyu0/NTk42+fuxwIC+KH7iRZyjIZrwdO
nGQnGkIiACnodulRuu7DbfCDj/6+66klfTYafz/7FhyYlDWyxV+IDrFJv26pe7v3
YonrCZhHlAO4QemXKIa9kupmjRsx2/MGkDOrfHf/EwZgviDHmkLl57XQAeRgLoxT
2WJ2J3DlbllQoJBWvHOTdxW41mNEBRuNavWyNA2MC16TCIf/pQHP/KaRV/fiFBc5
BLotSQ4VVBXxV+1xRqiTtSoAMPJ4v61KfJuBgRIDIOk/1dhMZyLYAYKeK8ICm3SV
AUcMrqGTjcXs90EoqO6YeZ4zptL+bGiHHwpoApPLxUoFF2zHm+Wm6/ptVsA7rqCC
x9yaSIwhv+Qx99kPLXZxntlf/9kcdlAh+oH8vMcAtQkJ56ArVfaV47Fo9+WvWq5h
RVvmbCtc/Ltut0pJwH/BrSL0ETDGwzQloD7fwg3Uz+2X0FpNGTMQObrjyD9KtJSR
CyTTTR9Zreor0SDhaRgD88ZlzkdHxKUNd69LJi9pX39dwD/RslJ685/lMOSxm092
IQbsdTJa6S4O2OIvJXQP1B4yK8iJm5QQ5lLOozXFiQFReke4wLyNRKtbGPprcEHi
2kwMb8SodsU++lzJw4rZlrwHJPa8HsGDvft78/hA8mlgRAtEWP6o9WCLRqCNf1zL
DiO/wo5Lo1q5eRd+qrYIjJDzVtMwa2oWA8jd0h648d693gnPpGO/bBNa+Alof1YW
KoxmeeC9LwXM9K1JfJOg4wlh/su7WXtcFhNs0e2OPkvtXcGT+5/x1sp5VY18ZyDB
E0B9if1Icta9vq1V3pfrycP6g0JfsXEVg5foPyGUWrAI6c4ADQIgob+tQE7LMhPE
A6eWZEEDKAwx78ETvbv90xHdWRoHOANaZsNLz3VdztRac7yXTle17CyKIIUDcM5W
wrMGTtYS1+a9LmxM60Rk/etqF+CFEv0DEaVRvxXWZCn9tElTPAOTZWe7QJWKfuUH
tsxVMXK5IB4VnrRelCeV08poFHAqRZrZiGYZ1DS1+oq1MSbBUtAwJFDrKE67YMDM
1rGmtmn1WNs305AIEu+CFf++BydG9iHcsOrm8dRD+wgGZRsXBGZQVjkPDW/tLs8S
BooAU3YWjlCrp+0PbSWieh8yKy8+/yHJ9i01X4aKkI6XE0bdd5Fb1sxjJu4yE7q4
O1IvU3aX2FveRf88P+rNMak4j8b0ObzXOsDZgCkJ9RKYa0tplb/FXDphhkNeoDOJ
XqrpY75xl+ol9m/lDGyzKta+uq7rZqgaB4Rhr+Z/Qit1RlzGpxtA86WHPp+m0hKw
vZmYfz3rln6wfHAlPh9TxX86QgqJMH+WABXh79bShZG3o934WSDDn+18tvYMQBEa
vSWs1GOVw/zuvZb34r4la6mVh0nLWbuE+orZmoNJkCaQ0IIOzaSz2LOg2Oo/ck68
lqGizgeEh7qSf1fEI4MPu+jqw6Ao0jmy5b2p+Zr63EEc0gBcMngv3/6znWW4pjfv
wEXNnwnwz8l+LDC+5OZpaXmpQI4SPhgPku9WE6Nk4wnWBL9CiTiU62+Ddpf0VDyo
oWrwltnb/G27U20R6WHJR/81bzZ7aKJui0WIGYX47QOe/c2jMgbYitRmWipALaCR
3oT2hWiTxa15gBn4kT9mVAbhIubhOQC1MtfyXtxO1X8eUFTsid5c0EVoVSqNjCvG
PxrXjghsGkp5O5TU9g2c/d0SLm4FexsrTWHeYQA6+SLQT8u4ORjA5ZFuV902dkzu
g1rlYUspWvN2a8OVDxhtQYIw2ktaRtdwXY+17fKHSWiCenwGVu6+SSNlL+B2Eh2g
gablfnGdKyHPUIP4DIg1ADwLO3kzUErKH3V1HAivmyTWZGZYkxf1p9Ab2/JPR1ZB
fq+IYqjm8dkW55xVd94LhERwk+jekjSKH0LcfPUgkpmYhFGtGXmBNdgx0u9raynH
NJZ5Dz9DoiXDvQLuehKQV9goP+SBfu8CxgQtdtX4xnVWyfsP7z2ye0JGcoE3pSUi
Ig/v0eQTVMOIjC0B6JqtNY4SMDPcx3Cr7gwGhv1E8mVB6vqPpH5W59AgMD96LpwX
Nmymn8iS/2P8oqsfJitV/AhCWQ11v0wacxXtGE0bY7yZPV3AqS4ro7rV1Xs2YBv+
o37F5NXNnIZjXJhQ3QgKDsYn6qi5bJKMZZKTEW+Mdqfp8yFMZJrSzltFX9pdkus5
0xdjfBKyLiwUiGXfmgDRLvcPZpy3nKKL0ztYec0iFq/CbxWIoHQolS4Qw8EO5gVY
oHPRtUO7Iyu1jrlmRaUgT0sURhxSeK/WdhK3zujXxHPgyssdWXqv9HGxpQ8mWiKI
2YRuCrs1I/GpIAsTYPbZQmtA//cfNwbHbsUflIr1k45+0F+nVN8eAtcCIPu+YGeJ
Ma2hgSQpHM5RGRczyov6hRZrGt5A85Uq3v5Ofkg5kk4iZiWuwtilMv+24oefAczz
Yk2aw+slaojki7szJ0kOmIulC1c1B1MPGR9X23BlijU7ojMMxSSF8tpvPOQV+1h7
k+RPFHwyjz3F1XTbttavDoXCTblN03vlb4+fY/f/geqmUp4pfQnIXy4YYyLi+zhr
o41itCAxBigGvwxt8KJW4PFiAZkrFv6xmlCNQEtzIxZ06UVbFhw02rPO+mg5gJJH
kHj2O3+SK5N5uSnPCLGRQVbqBN4B7TbyM3eWqkMz8d+4xcMGJwihAFfR8gKLXjKJ
9U/gsihs7fQwZ8MZPLvbTtPHZf5aVSWCnCmcVF+NdsPkq8P0GcDDGYGr+TwAUlbP
a6NaXUaU7Qvq9H6hWlfBaOC2cWnpGozvNJaPyO48ORUCq504/G15WNcDiFbgbBgE
9XRUMfLKxGLvKk3Mzlq5RDILi9Yh9ThRF3DLF/uMN40TCuux3pV0gl1IcSSCTGUq
zRJrm0N6VZ6AskhkFwfTfsQ8AuTslbTEfWkYM39FrBV6F665Z8ajP/vl4LweJvHI
YE5KaWRsNKqAP+efW5u469q/z1RH0/YE9N5f7m/9GGc93F4VXHy284QhpMxxo9hJ
GbIqKoOug8dkh0Ka/QCYa0PR3Oky9O6m4gGZ1jT9RMJ08u94eGHPm/xEIzdLWklM
lL30dWKZFlwnOaxwJdBK/USzpUDGptaK3ezJyI5pHnSEqAlBEZ9kSwifx2Z6uN4p
48KjMBgMlSA3/9ZhZx6tkWt3baTpEohVSUAK/BATu5adqlw8dI+CwCoMTmKq3w2e
DtqGaAmJz/u9VDPjFPWcjUDg2r9cUc/GvkYgyKJEzxJ18Px2nglElvbme2fneSY9
uvoReRyS70d6gIeiX5bBNBakFOarN3xrwDUWSoNepENjvBjf83mFsgWK8Eh1CddG
QNpL2z2p153LsCkee8lpqPJxhqH781sqYiiQRD3Y2t6YXh0OZ5B1vYlCndXCfVkn
E6V4zk+xfOhIbq4cWCDmr2xK7olu7PkWeGpHQcbMnwYWrN3guVoRwSp/Wpr9e6Eq
qolw1JavdQZug9C3F2c5wasAfUoetiCU28+fpyaoSwFx9dlkmmpxh7rjhHGNgROk
6CHUfASq6824s1gU3Dgbj2HN88LSrz0jr6CrdZuNRG4zZ/DM9LBSM63OkHL7UE+0
jo7LITiQTCDEEbpLbGyMtH+/Ney6rdjfCycxDHdBNjObFLEgs1rvwjwb8uisT1as
qyPJN+1ojh2HffuUKDvl65FCilwAabSltVl0MyWIs7eTAGcsrQsRk+UdprNn3tPv
61qJDiW4U9oHnuCkK7EdzHt4JHLw76Ia7S3Ei8edRbD0Kodu5KNbeoLpEMt41ZAD
4DThVji/71tyokW6cIihEHRAeGd50XXjtvOpRgGmhVHJbcKQQhstsutcn8xnclC2
rj83Wrrv18+CcBWAp9mu/sUivtsuk++2ioWmNGIyZaRvExT1uVaR8MHmPT/MjBBM
cwLfBiPd+UwEwXCzYFAN1495/bpM/RLFwL06CbT7iDiljWndjEHzrb09lzlFBj+K
sHwrzBZ8Z3PDmaVnLgoRVunZO5x2eiPCnAI2kalMfmsplu7fy5LSVjTpkezM24HW
gOZ3KDdVcjPRoPcS3+ASJSzyrc7+J0OLBDmE00pFUmHoKQPH4+5Feo+x2V05dgIW
+roSVfZNq9nOSnzDx6QQKQwKGbjWJuX091MHz3z36awQx3UoQX+5kQ4M6mSffCAa
8Lg/wnmtLM192nRORnxoNNmwZChuEhQgkDfkaJdTveZGhcUH4JW2U5n1YoIVEhfo
+cZl+o6Lu5iri18THQOQ+lMVTa3g57tEc2k2YPxlJ7VWstUMeTjrbof3UIlKAwcS
/26SWGCuzpzioGHZUAVLtSJyraHW516bM2zXwsSHgi38DB9vfafbG6TJsdVvC6re
CBhqjWDUXjbOe/CbO4hoOZSVOKD1KWNOyFGAZcP2DxIybIW0stuQcfogkwN5p6sl
5Vc8DxFCUNNIyHdwC39taGV50Q6dzQ3O8VeteQ6syt+CwL3IZLbKSj5MZNwRJi3X
IASq4/UvRmDox6U6zw6xrVWsrL5nE+JpcJxOkjd+to1a6froY5MiLV+WbZOMMxpn
igXOX3iBQEeSlpykq59/tAn9SrGzJ4mYQC34sBA/lZ9BH9/mnY8xwi91WZ08Neng
x8BN4Dy4EpzPrIs7QBnuRB5hJwfIQERu9Xwat9ReBhVne9YzstMepKc+5wUNeGWG
GheSiBnXlHfWpWO/wm0KO1cDbvDaZIMBnKdr7aQApJZoqnholXrpXEgA0Q2W5krQ
lw0xyCMdxVY42RciSUO3DEa5n+oVan6ls/9NzOtxPfEkvPkktgJF+GCyb4JCh7AT
3MchRS8xfmGfRlM582XUnfVUdyGzHU0dhQW/VsxXBWn/NrAjxDkHEwAXWYiAINxv
qZhtOjJ5OCZgSI3R7XYXpv4hkPeJWquoStTzsfWrzrUWE1lDUslSD9lX0YtseDZ7
BWITNo+0AglQPct3MEHdDdDIB+9fmaRUHVXkzXoRasWb3mXDkyWj2eofGpZ+Hnt+
JH8vBez2a7Y95aNCho26UmLqMAwjSq0UAQxj4eCN78G3zme03dJ/O28kcK4qtzjV
snK7KGBFVMIKwtTXaYQTMlMpN+pE1nU/TZlQCboy3SkTltJFJ76Z17DgSqRugCJt
+k7tPiIjg62RO3o7gU77w5cvRvA3gvwvQRlQ3FgwUiShBwN2Kge0zZcfSJTBKC/8
Awtl4h6Re8NGXAjOj4UsEdz79tmMdSCc+EYcFqrQQxQsDdIGdXEW35TYgW40PJyd
OouF6SSIWo4cPFSriYs516Mog9SHkYvkRtGkraaLxFsygUwHR18XCBwEao2LLtUN
B1Fof2a3fTb+UHuV6UQK3I8p8zeHfCRbg/ILd50Arms5klXxQZsNhSHO2gllu96f
3gjM9wBE2aj88XRGEUDv42hBeXrgbYRrgaAPn/xeAKnnRz/XC3UiHTbJ6q1wkMgO
fXRKWpwfntXBEcs0cDcavY6Y3k8+DJcBRLme8peei/SQGReoF8Vd6CX7DKNAEtvV
4K9ve2MT8sAgsJywikwrgQFbpxTXpRWa/Nm3wiDXQicxpNoPyw2MM8n3ztu0xDBf
09CVISGKYpzciBCC0XwsBcV8nH8Ukh+zf6wuvw0Iuo/lt3vWAdbyJKDqeZauS+Kc
hFcMWtubkyAQj2hrnSDqIZunkg0S6aV9A6dGLrCvNRQZvtuXUwm5MiWlhN5PxHX2
GovU+HV6k5RKmiOeR/NTRvaj/tG4Qe/jwa/wHoXjon9dTP27+fEBMrLtVzdk2bFt
KQ+ZmOSdSwYomQqzPaXuXqxSyKwMi8t7tJ3DS6i22fCPeF2j7Or8R5DgL/uPNAR+
1vTrULr9k+lfHKYCKqrY8YX6Z4eaWQhH7H7RpJvZBimAxUl5+12t+AyvZjUu68r5
s9N7zSoAmiWAMTdYWnuuJf076SMl6F73NIxqMowsK1COLX4GWEwxrLuo5gYTYgcn
0MCatJUz9PEcj9wkHoLqz1GusR1c9iZwc835G6z+xGiZIURubDwIPsgRmwjFTM6q
YNK3m48xgAlE7AXDo27OWRj4DkHw7+0e2CvmowcGbou7n1GezCPqbyzGTyrMXrXB
S4AVaQeB5gmmyCmWHvJJz5xrBwdN1XQzrW10LbbTeVp+qRogatD6hjdQiNMMpJH+
qepf4kpcvry0KXKSkoogBOYCk0Kq1n/4yEMbAzJdDCyKfW+++KqFEgQzfXhUXnfn
T7qT+YcWfEAEf4dDc0xXhqe12JfksUy8Qu9tfaRoLs8b2MfYV/rgyISQVjd7Lpnj
3HNWmdZuR7z3Tbzvb6/QhjdPOlcqSX4+eCIK4rsQKKgNRxaDTmlNrYSJTuIhalTx
jsaLM1VKI5wiM6EcSKT66Qx+bCmU4gMfOly7Al8UEjeidoqVMYRN5vw3bDcgGrIX
chyA7PUG2aJiAr28iqUz0T85zME6PUEBJj9UYKKiPFCSJ44tm/KJ8X/lf2rugRir
fKjsDRMGFgHcPwB0ayrdO840KZRW+9l9qfIof471pook5/wNJwSNZz6Vvf8GUZM0
1iBz6u6kkBDjk1dJCezorUiOkZx/Gvwghr8xbxHA8kSdGtd8WSBAYYFX9qdUwtz1
lsOiNFzaDKhLoXl1vEg9CY3rBp52iRKB3jJQ7fNzPGq6S2pKWzjgHYw3R8wPY/RG
+o4ZvMffjyDLADc/OrXCvDEdzvMROQFJh80autnSHJPE5VGgjaj1qe2GhybXK9JR
vMi+EG6vSkZ2GSHD4k7TK4O1Q5yvSESCcxlC3rEG9eK6UlfD2j79kGNfusWGQAof
ZR0nvCdR4ZdEwbL/n/tJBfah40+InO1WaDSI9TrUQNZPjXobg8gpUCLLD9TQhWSr
f3JeLzCgYS2jS9/5RqwWppumNlDmN+yLG7r0LBvTeoY4X3r4vmaPuJQlWzAeN0cx
c6oWogLWPHiD76e08AvKyGU1wmZw48ZULa/wTNOko5LrdgIqMDZoJQTVJjALJBoP
kWkTgxtODnynyr38WzxwmMbV8F3V1jxIBCNi4KreDZjw5Klwe95Z+lVDKhzzAFQr
lBOb1pXehHGgW7wlTnJgran3NK1PNPQZE71TMzqMc59K6HRpRe1Txej/7ZfgrPrK
ED6ktj0WTnPtHYOY0JUJ9mJSedkLfguZbp002WIg1ndZxbTvkF7vcywNA+Yuw1m0
F78nSgaP7SGhgNyN3VoHML2tse+ClhsoAU36bCs2NZpfYtIOhNeAeIneKL60+tMS
ArY0Wt5rHTqH3Ms+e4PoRm4poNSvn/yxf3ln79Rb/uRWhv7BDg+lv9FF2MSWVng1
x0/1o0zdKGv8bD+ZXV8iLnoYNN6db63lFLHoOewKvbtioKynlrpPNBXDgw3ghsE2
7WjHbM35klfREMhU2HahTerBk/omnEkfQWKks+aYVrjA0NAtTDKNucNNAvd9au9T
fabsNNKM8M+qlhvdwCGvt+74pfX5juY6XBqq+cQwKh13/SIxqj5Gd4xdYzGH3mLd
C1ee7bXQ95VToKrB4wOjrWDbNhiT02l43uymsdHFc99TX+GrTWcIu0Ai2mud20sg
tNzXi1isIP1S78tLysZU4OMeooTK0cBfIUhYRchW22ey3YuYMUpCzniKkO/PNTMM
4t8dEl3wrWeRrHb2maG0B/cpnLdwzW2GEZX1FLdtkgqfVaWyZG4nRVuoJJKFSiez
Q4JXMU+r5SLxhcFmwciCxy6HkJksZIV5f4tTl31pzrrTGC/nma5gqkXKwdGOSVc1
OVzpymwfpx8Ko0Ywq5PSiGx57ORaAE35BnhDgSKt2nQ7IzjGQ8ge6KHp2PBrRjWX
RxVwaL4Dy8qH1/Bjwd88gWNdbKYjAMzFs2guRMKYf6/m4au6sagJIqptgglRxxG+
J1/7udFm06SGb6K1RRW8viO8J7P40n7JjeR49qMsDPL69s27kPn68Qz9jtPL99Qc
VDA1xqeLGLX4X1P/PB7MvtrSuqkDwE8CRu1g5goiAhWWX3S0qgOYFfclOKvsZT+9
Z5nmTCkdXKWqRccoSs11K2m5087YISaE7uNxOZF1jAHe50L9mSoS0CrolzEL97A9
OqrvPkDC8NtPWN5qOfl+Ja8jQE30msVlSx9q3GM+7izeB3X/IkAdIckWpiHbYzK1
nJh+gXS+0Jrg2SqbX27d2RZZxvza/tSZu+is5GsKC9X9g6QiR5J/6ZqFaNpedrcS
e3ICo/A3MoflGsOkMHois3dNJbUz/+LPnNY+DbzDdxHfjdf9u1Emk/bneYlYo6oc
78zb164wwG2PqzNyJxEugkaBN15kaRZ/azV0tdpQHbkZXzEr0OgCDJ0rM5jI0XLQ
+VVGBTpy6uicAk9Q+YnhkYbEnuHKR2dyqmJpwKxfrQCiiYfdpi40jZCv4MPKeJ1O
PhwRIWjawIvWbwfoOUqZQkj/A6cgED4DuNlNJi5O+G2/F5ZEisuBfnNqccefd+YJ
8se+nr9MomiJfOoDcLKtkW1UH4lUKKjL9LJiFAbtCQ7jam5lyvy9gXQhmlHyM4ud
f79ZdZCTjX9Y4UPeTpNtWyU9L4I1N/C7LTSJ+ECCxGqWhLX5SDmE5491oXpwyxXW
X27kcMsJ3JNCj2zFhfTsD9jjjn+QYkyn6UKZdVYr0tPkFqSKZHvis8Wip3XVcIOG
9Uy2wYzzIF1mnWFbEFr45zE/buvrHD/fFiL7nvzk1gySKIWWPIiJUJ/Rqix/ZPnr
nHiVXBUBj+FMeBG76RMAnZmHnrEKqBrSYfn3HsxAjoNsvT2AZSApFfM50m0rKaL3
EUl9Xp44Q4k7DJDJnaSI97+9MKb6DhzNH4HO5LxGoBup2IC+RmYBz4s4lsjcc9G6
UJQRcSBrbw8dFmCR0HHqiDX5+VfT/wlau/zt2OMWiWiTffNXRIu4VndX/VcuFbkz
rZ3YIOT8nJaO8326VTIz00S7zYcTzOc890HKpqxc5oPq99gFuSjWnbtgccR+02e6
srl0CupaMUK6I/tB1nHK7fvyUmz2G8XQhlSS4fNkk/4Zy4kxfxKdRf6alLL1QRVe
s0fRauua0cGE22iw2WU/L7e9NJ8/+UPdMx8RStbT4oshXq1r4fo0e/SGt4x61Lkc
gP7EPIBaSQXrW1i5qgr2v2wr6ISYOh1cWR160VEkpU3EqC07TofveHvrPmErHLtx
G0kEHLBS7n/lIVMlg5KGl6aTKYrR2MicqpmhmIWCA4QuBk3VhdCufqUCc2baQiPE
Yk8NSgIBdnKM/0XZKNoCOK1+PSJOB8kaxe9g8IsMv2ln3oYjRaE2U7YDb8ZFmZJ6
dwTIUQ1mpezygb80WwWaxM9W+GbC8a/wCtDXopUAV4mpJoFnm/N6HUMaknCEEf0W
h9G3QP7h+JcIMLtUwQMqHjd4c1cNeupqWGcif8dUEuBzwU2C5VJHDzhFM4GuWIj7
d+SqBI0dpsC6g8SQQpraajabvwOfhrme3/FusMQcaiZHcNpiFwbPQO4Y5ps7oqSa
kIRQ+g7953iW9N9d8MMLqpfZRm+GLxc03/gmkZ1fEPtkSk0iyOEkXRbuMYBfBWMW
um8LHqOxGP47q7t0zBhX2bL0prNTubF3feaI6bRqMkR5qVw4VUIpjgFwqawZFOHM
3FcjdM8wfw3A3ZZpPg3nspA/prbO5tC+X3GMBqkoDebi4dlmKV0CIkdd66VopRVT
/+PV54M0ZyXmNlaOsflIDJtnvtv6lj91nAsHa4571bUmAyUUMtNrck67GgZdY3j7
gzYgAakzLlQ/Nn/JqcgaQhCfPMmontqWVFbStl3fFuMVHc/YHKaH6DWZI4CeZuuv
74AOaS7mYwgWl299MyswiMQXGR+blTg8srD3vnUN4sXXaW7I6BtpKn4I1ZWyAfic
Gf4GCGg2gR84ZMTadpYILRu3Ya57Kcq2245R0nnacRudYOwiJ4gRYu+W3KOHTx1r
vfWW4K8vOlWUo0kHe3RVqO84CWu8lVu5vkX3F21+6nv7NRAAHuZM/f0HYWCq3h2g
3hOZDX+Te+kzDJMX9fp3n3Ge/LldkOjkBahV7KDJNtRRz0461Jb2A7QlmmBWaoqY
mZILTJBqPo1HWubVw84H6/3DJkfd0KpOBs9ab0o17WC4ukiTir33jw6P2TSudaMk
JqaCkkCt/BHg9ZKLH5RUQHixcop5CW0Sp/P5sdZaSEiQVbVb3xCQ66VnxrMYE2zo
d61qq1UjP0TVjXid27C8lAMByfB0ScPc8UUf4pxoSC3Tm2zF5IFM05dMSN81ptjU
92SEB+TijzLpSn7ft1qLn46TiI//r5gNoCtxaL7spqHSV+AZ/Yrmc1z2aHwxnWyC
G6yLHnd9Kqy6Zmwl1nxb6jhZjxxBEeLkRQPmuhWfQ7DE1VphelNBSsbL066Um6O6
CG1n2CWmxpSdCfN+SYrDG9r/I7xqhH4xhZa+X/4FQ2FPdYoJX1RvY6U7Hc/NSizH
ILpYtkaG4YlrGStm1kog7CAe37wXml4aFX7lWYGx5/CrUjwrepI8eO3CRDAFtZET
QBC79JeAm6hP2DyGswUqv4I1jL7frsILKwcUuIBcldNw0UUrhviULKBDerjP/mqw
EwD81sdD7OLx1l2hc6DICFDbAMYlzPruKzYHzuBkrkK8a0br/+VoQs1oF5GqHPKK
p1v6gBrbtHASo/nQQCEX21zHOA7bqFIcjAD74YAuvjjRaIzFMi5AylFhZFT5ZmHf
nOMlvaX6zs2CkTSj//fvS5ODpjyvAIn401Jti7fh0SSOl4RIUd7PzLGdpgITjMkn
M8jC56ODZC1UV0K25lwzoUnnzXtpiPSuRyUmQ1aESghtMhIrCwqTwh/XBYiDDqS9
TWshBWU/t9CcLuWfUBdNI2ZAVfTaEvl0QY7tK4NOkBN3PYlS9twVyzmocdYzkuG2
eDqzDA+Q7MwJbWQSq5cpiczv4f8FFQ17y+IsRcqN/ltPFNsLAMLwh94TUeJFDQsu
uGHcbU/IPjWT6ku/VKGeoJNXak0kZ59Wt/BvkFDMbaghbRH6fN9A6yD/VxWJ2Dba
VFWQZvLRpLO6vIbTcNVS4/BBnETGktMdujgTI51hmLqNnTbaviQeg+vxxDBDG90B
Od28TZJZJ18oHjns3slhTU9yWQwqVvQHU+uZOhqJq+PqIKQFOoMvFsv1oLhZoqFV
BWH3u7djqz72Wy7KndOSurPaffIkVq35kj0i7cNQw0wnwswGUWGTIl0bFJmk0xNZ
97dFLj5sDg6CPr05KYZID8GnxRYqLGAHIkodCZqc1mw4fdDK3lVyKAZrvjeWreKr
dSYTsCOHH67KRheQk/1vFEtTxyPLvijXZhcQ985xNqst0eMAhPJxlDGAqBgXp7xl
D5aJEN3RqYE0NMqalGeIkiL1CZWncfi8ORqic5i33N+6zaXlyqiumYu+jChJkRBk
lMVYnuqzg9maAG8DxD18BQNib9i/eHJcCXJHhmUNN03CXSuCTKPN/3EN2UrBaAyz
6ZTMvNH+162HhlDxMLyJ7uC7T1xHA6mWHkI5PBfuiqAxnN4XFreSWIf7Enth/STe
cHUxsxlyPECIN9s78SPk/VEXyZVWPybwt/4nGo++EYjruHqM/Uniin/fe8mcGBa2
35eCPotzC5lge7Egd5Pw8NyH78jwjDSUBFbni8F0ESaaoJ7tXYuiKtmu2Gw7RlRv
f9/Ntyf7wsSskpn8NSq4S3P45ugcUIRg7t5b2pCEKFuwA6HXPoM+NfQ80D4+srPu
jyH4hF9NeqTsuO+tMwY4yjlx3YWSdETZ3GR+RDUxuKz3RNdEbG8iziw2THgaWmNL
Zw8l5MGCD7etMvJBh6RPUAEFtNXb98EP3lH1E4AcuCAyh8Cv2r9jmXwh8o54KdMa
ZmvpCWLBu4YjIjOSZ0YftBkhfzGdOMAEohqI35AhLnFpSwWuBKyGhFZq/ApBpoi0
wbAB8TfxRqCEf8w93sRyk5jfKGYQEcuuCGlUCyxIKx+oVcaV/DI9KiyoBDTsj2vi
G1hodIjn5wmFCh5AtTXjUPixq4qDSQhDCNbkuMy5Og/V65s2aqVh45Ta1P5elAxH
K3u2+nQj5suVRXD+TAVwYwGYTg9cazTAjB0Aj/tAp6AQJ3qv50DSUj4rLkaCrRf7
Aq6BEnfJHvEdDATzPy/vzEb+QwJCo0Zog/+ElA0PPJxUeYMyoA4PKhncidKU4VmR
OQYiDuWKJw6gLZVyKDHXlRDGqEKjKIKbeni1+DNQTi1YiOJPlKG+YLAjTEeLautB
OEnh31WZzzl1iFiwLglzBEnOEZYaA5jmMNiJWSNZ/FhDsYILcLmvP5TRSEV7XieK
igjnDGhbND1TPB4Anp17Ee9gpnHcDlaT5sLBQeLs20pR+6kNsJmo2Fid35Q2Hfoj
K5UiWZuT1ClI3hozljDx66DeOAYTOliINYP09A1CRGc+c/YRtr0osRxv76XPdLSR
eX6EyCmVLWMxctmjdjHVuWJwxia7xlE39YNESCCcsrHJL3vMYMqSxsCZqqRPdNYk
dP9gE61MAgIS2TTOTBlD6/yJGgdCygBuJg9Q7GCtuEV+hGvHwRED7qRaoHTmmCv0
//uTHM91vvipF1qR7aJH6C5RttgZQXRI7vDeLtgr8lMEccfd4URo/HJJ9XdWqZgc
cLIQeUenDfScZ9DnYrU8gI9LQJtsqRSixJDfCwIdzNfvedQBq4Q1FNuW5PMNjG8q
pPyxmzT+WC6guISAAgrMSvZaJ77Gm94kQZhw8IEHC/32Vez3FkGWxQnHHoOidZ3r
CQ4Qo34B8HEiJkOEe8VE4ZahtJMppsRYHb1PfqYQRxbzQDK/ijgAPcDfkBYXsNd2
0WkjnPEJBgpT8LcpWt20Rsb6uQ99a9pbikkZ2/5HtgtH3CvCIdBCpZ9UI7o9WXJf
95ZxRpULHrJD8Y4Cbz55PfNDynrB0WS5WBjJEDlOt73th/r9NmXba89vMkOHz1sh
VDImvBD2S/2hieQ5zl7p35lLXoDZiof592qA9N7FRJccSNsDupOZUcu9ffggFiFQ
3eFKQ+pipooGLYJ3yAhGMzA3LB9QCj/EVmQG3XHJlVDrg4uiG41Ig+0Dvu4y7Ln3
+aljKwcx5kBWZJjvE5g9KijWkcHPWvPDM2sZy9IckoqhzjSHGxcwO2p9q8Kjo1GR
dw6tNuv0E13rG4YxBLHi1rcOVqtnUJv/FAtu0HlvK8ixH9x4lQs7TY8IL9x6D/o3
kLupWyobqyd/hxWLSmPh6bw2AcwQ6K5luEuB+SIHS9rLtNxeyAHQV5tGBH0t72KN
p30BFwyprupr397OTYeKNjevrynJdVjqwkvUQIM33iSQkCMQL6mfevFgvwr3TUJV
fdeOsCC0y1Lq9pj3hE5AAVC+Tz5p9Ay7Qd4k7S+KQ1vIERRXqHFUc1d6q0HBjlCg
sG9/bNTjz9z9nNWyCglrv/xnBQqgqKDXaOSIfPAYX4p3Ynd3s+yIIBmzpY8oiuWO
GeMM5KHP9vq81jJvD2efLaMcj2aLsVHUSrAT/900BY2Sp9ztEZsXAFv38FeSMgQX
MMhuSqxjrhQWNWNY2u8AyWIWlyfdHPafA+TDcgvvRGr+I6wItJcRJwbAzop+op3C
ZwHmnF95C68McvASOmmHKWdH1Rg3tU7Qlm19PVcgLF2v32zToGSnHk/8cWjcwvTL
teIUJ5QGuG28J0SjieCxD53BsIV+63AyT1h+E6wneHOHxbfLXwa+s0bsI20EldrR
k3pBO29vTi9xpcUoRhsvw2b75YLbfgQshn/E6jxr4IAddAXskUgz1P/potM9Fzdd
OeeJQ7YlZ9dFQs209FYl6GfyxtPsAmuXIDZO6cksqC7812y/SRwd9SAQnWS6s2Kb
tiJtD57744mTX899fW/N3A0AC2uNCOf2GAsUlLn7fwjVWtYoLo+ajFXcAQ44ihll
IC9sm/wotakFolzUrqxnKiL73sFKxOljYXynFkfmDYUQJosBVXn/CY6X8UXECyfB
g/oS1b3e+v8c7Jsr2+BPnI2QDVihZZj8bcwt4KjX1alGsh+tp//2sg1STpWsDXbh
hm/bdD4PSpk/jy4LAYM/6aYnJZ6VHJAIJ/FZXYNdqJb6vhdt39ApR6QIHcAnAu4i
ytuNslWqOTF4mUPEc6TN+tDfaA5vVpqBhQ9igrJfsFSqO0/yKBTZrRAusPOCcxFR
a24/1rRkLo73PlEuMHNOZrRYhFuogSxuhMqOhXVzyGYIH0aWAXS7r/D2lIQ1FbBp
JdV2KZUvK+04Q2FEblJHnSksfVi0SMTytU6T3I7UXxcrA/emm4MZ66Q3ilUZdHsG
MTyknJ6sAPc+wuYQgMK8bqDYSHT61a9tnbOYsdjVBAAwWUwiFiW88QKzl7xhxBhN
LFTwoKWdSbuszrbeo80osj8mCDFPt7nZeGjV5zVJRf9JCF13cwvbVbIRxkLuEdPO
lx735V5oNU9R02BPmpLixYBtqCQNKK/cKYmBgaxbC/sJ2/4D076ghhrvVH1KS1/Y
uQ4tvrzjKQIXasXRTytmcz6G3dUo9M0ryR872mL9hxrOwmDu/uGh674mV/Lx0w3l
pEQgV4/Nz+K9q/t0rx2s3tfmBwdu1C8yn7zHtYgyo6AxjjkrNwO2FJFs4/1I35Gs
OZRMOrMkKeDy/IAKg3HCXWIfhyX4yJg9VDI164D7JJ9tvl/pPtRlZ9bUnUafiSSY
lC2HPegCrnM2VQi6kcWc9tu5Lwzvfgkfh2YQcgLkyaJeQ5D16Yz1BlTs7osAAlNY
no6lgfWAN9MuB6qEhbvgCu3q6t+97oPmDDQXjiR5crJ7WtdN0nUjdPgaO78VDy00
3NT3lhWHeDAhaoO1DyQQ/CSHKwzAtr78/nOAzes52F/ewqQgmuofG976hTFqIsnl
c06mB2fBdwytRTSsiS7870WhrmiemGILOtuUkj6hrVI3WE1AWkr6DIDFO2aKDYEA
rMmv1LgQbMCuptgW6Sqh3Dgv3jjv68r0/O+HCXVDorj9mRoLdFH1VH/BGaRPc2le
ULzhtq+rqxtw8x2LqDnhtScBrl5nfLI+3PoSnhdDT0w0DtwhkbxOXT9keb15VqPA
r7/id9wY/gWEcDfIsD9uxlRFHa1fvL++mo3jqcPgio4hQ1CjY4gR4kR4wl29T5sJ
WhLvQOlsMMPoXXOtGyVYDpdqPPyRPsdLz5jaLNQyCIfyXoD8ghd5PsL7HM54WiXK
kk2pOGOfL5Yl7K4ZEu9Xy1+VWP6Y16QswW48DMwyBz5GZrck31C1ZbOpUj8as40p
CUHE2OJWbVrNb9vFn4hWEdYX2NOKSnTtYipHVKYkNFBzPR2qTrFFDEXQUNDcoWQ/
HLTRqaL0nl0Jfq9gkS2hGmAunGvdWvfHWRpPoYHguXwxSBZvdJstHCsVLmWODTXt
hHtOxM2xsWdHjb95kbaPPprKXzr3wJ9tPeKknV0ol/yEMOsSU0yHDbiUtDOxjczp
bs/j5FqdcCF8Vo0r04eLMWxiqg0uqm59etEf0aH4xodz21NfzAhIwzdoennwGaRn
7ftFzPTmFJLrOSU+16b/C21R/pQbW9J5mbzRVwivt4DELIcUcBRqINUR/ZhvM4S9
L3wzvOXEwueCzikRWYDTMpMf0gE4qIPvwT0kMUdZ8IeFc+jfHGQImnXuQoPwhVQe
dU7RyN+ump42JR9iQBEbM27PTodBHfp8DTjNQoVBvHiBlLj5d5IfGQGW9V5zO902
jXnmd2HotaF9NHgu6RBpFrBtb/zBBYoyWcUSdjNRAdU9QR/oGyFtV08U5tr3Vmh+
1smNFCvwuT2bWsW6roiWkT+K1zYr8+HIwV3rcSWq59DPyY/5LAMiPXiJ/FV/iGbs
zfHzrbZ140dnsKU5JmGVmkPF1u7xSq3Ra5gJHcdgFPjLd66FmAMTQTuAfUYDMy9x
fTJOh6VbRN1Jpy7+1jOAN5qdEUCa0PRUpgPvDSRugUm4h8bgt2Ta60FyTg986YVz
Uj0NbaJ7j5014TsUkmLEGB6E+y87IafzcL+IxexylWH4awjnod4HtXDeXZxy54R7
X2jsPPLEj1aZ8RvVIRIPFB5ogbqrmiK8BQovDGx7trdKg69kYD4QyuVckh2jAijN
y304LpunMGG219NnbGLUiQReUnosb2+QilcqwZ0PcYo5uwtFZU+MK0u0kU8mdjlY
inKh7SPzP8k0qVkUs68rngFbkw+k4nDQt01gimyZnWfwsnNINSP9W/S+UyeEFFzT
FLS7KnLtNrRTBlj+rghTF8ipkTuGnm6JWCllO0TLAk56yh4w1RcTjrmqvV+z1NNp
feaQRVEh0LnZHOHg9kVRK+LpJbeiomAreAZ7NNx1Yk3phpLagdXok8cqKb22pKaW
hyhHr2XwAIVHZM3l63lbrSxlCo7k4FtohtPeX8BjRQOewF5PPRb9xz0bQoqYgP/R
gkpu7EEz4Vdy0P6tjer9m/6tk2zJ9mamnOsI45d+6uenZCdwW0xS8u3p/scnKL9f
GIHpPQLBaswvJD9N29O5SFzEt8md7QDxcMRmFGgpLH190EsfPZ5kJpfF0vBGT+eC
P0kMzY1e06JjyDE6j0xuBt87p3szvdrrh0A6F+tTvu4wgHZQv4qH3LYq0VYTdKXi
0uaHM+ODB6MjbOp1kSJVncBYDi2i41UFaTRS+5lhDmJEXvIlWFXnGrbbsPbdKREN
yrM66KMHbwd7ALYClnixz0B6aLNxfKQUzzrv4g2ysGuiOx0celooc+X1ksdpaq1m
42NH26l+DzyVaBQXA04K84OgNY6QnKH/5tM66MBeEhl4hmtqiyJfCduI6VqzOzLI
YsT7AS7C6x+GbBqNytFYZA5odzUUA8KEV7R9XOys16dR/Xv+cIBq5f7pRCzqBEEX
rUYQvIiObrx4bSCHbNTQHxBmaQgPt50ZqUZExw5v75JUwyShun9Lz+o2FLSX90OD
LnSlLn90iyx643NL5m+J9Kv1zEZW+773Xnj1oCnvp/YoxNrNp4I43/Lyn77yid8m
zahSThmrU4//iTy+gWB9QJhmvl8nyP8WSPQQrauPnb02JR3Fs8actBRnoIOyyRYi
xWcQciPlK/HwJZo8I38efIRKSoje/tW8I8duWrOWQYrdWwPbWeXCBEwkBS7L0Jd4
V34IrUiyvvsNvcqjGztLL0t/UgeOmmhYn8MI5AXcFeflmQOoimJ7X+byqNArRn6m
XMqzDPEa0EIa7t14naiYE6yR8S4XZ4kjkxn7MkLwfJsX1JoiCusBA+21zmF3lAfT
plk13fnp90K5budVJ8mbWkZxG5L8s89rsXCly3IMszA9JnOg/5viKXzr8l4yHKDW
Ttzqyq6S1tHTZMwZeZrOpy5W/T4EN+/nHq+r4NMMh1y3ImaS3X+NK+UsGFLx+DQu
nI7n5oH4GKDovcdFb1TBr6ZP0ogIDDatfIWpm2Tng06wcJPM8wiFjPoTVtgDvqyP
ES0G+HhIizK1enw9kDP8Ypjfk30+hiJOI4BloChkeFNRrXJD9hx87r/DvFRjVMWm
ygzQkCcLICao+KxtAtotf9ia44fTY1ul+yReqkRphRxxcIYd7hdSr27BNqmVk/tm
AAn6PmQKfy44YHvSvCpqWqbwJLNcK8wJKNv24SegfyscuVaZseKcxz0mnt67nAub
8Zj+wi+Tri2aeDYT2D7lfKOJuTsfzBOcZldatfa46HZA3tJZifqBGU9KsRhU0RCn
dABauXIuq+XtbpjPFqcs3SZU60VzyZ3obJFOnahIeNO/yLqeUw5aXU9WRfC5rZ5Y
gwpS0U8lAve5iFMBy25lIO3VSXAD8yJa2aQnyfozNtbMsJc63Nf6GkoyFeHkd8O1
7drfl+hvOQAVjP+IouccYlp30Cg/bpJEBbK6ztnrGnFqyS6JZhkKegvkQvIFcdXU
ddtUD7/06y7Gtm3CtX0UP/v/GuD7uYcqCN5sKbPqyIDcJ5eNuhdXx9K8O/YeZipL
YmO+rmTmWSeetU9wIHKpoIdcfSnH7Qb5u7vPnB1wfplj+PYIVTgk7k4uYuwiyiMx
3SR/Pz9ezyGbto8xm9PF0G7UgFstkWOb5d+0fd856ly18RqDp7WxtaJYbouIggCa
z0va5AdacstSuBuFA++1kUk6THtMvCfQgvKbI8l6/zIFIlEbcdrH8O1HsN2C8H+Z
QbvbApRkjFhAEy2zRR/Iv5PFkhknFlnFj5Idb0GWahzRJyNOGDJnoeQ0uspMgDW7
DVQa+J+LJDTXBIe/aXDcx0Ot0ofcktuDvvU55mDYYmnlODNKwOTAumcLptc+wD6v
5E3pUtTbLIgbIK3xgeb32i3cy6TjGgqmwdpnW8kdoJAiuq8359XShZ8AgeuVWKP5
kXs7t7Mr/1qRKmgPf4ln9rSyniKvw3RYNbN8/GXkI8exzZfP1hkCtJSWOMlFiJhy
PwQBpOBLVoplLMeFfCw3ziSpv3bf+K29WjfA4Jk11q2BfxzFOsFkIAdDfCCeyDqR
ev1NWTaZrxaX+fuIUEC+bjHVW4lZQc7JaZfoM7k2CLSHuqz0q2HGzepwNVV6fFIo
yat8FSrtv3uVBdZrQuRLbaHd/5VCYTuHgGHk9x/psC2rHQaRkODq0/OEOUmcPpme
CGET7kTU0Ybpn0Xyou+I/RmK+7KOD/+f3xExdG/qQqxnmHld9I16ovVYR5eagRmJ
976gJlzKrTBsDLPlUGRb+gt2vu9oqU7AiGYVRjzJtJ8Ghx2CtmPA7p1e8Ltoycti
YeoD6QbwS0VMM9c/Y6kz/v8QBu4xjkguS5CWZIVaYEpaPnz4UXJPD/zZSIyEBh9h
VBpeeSs6aKOf1ApSLWoQTDXdxlnXrCt+TfdbXgvh9ns25eD286eeCoMnOFKGpbbu
rz3r1sqUcdSIqbKlRr0B5sySmoUr4GlsVN9sbh4TsLep+H3/nQ45otaDvKDOC/Tz
WOPWIhJU2in9PpBd5NbyucGhDghKM77MMzBszXY23u3IHSY8lxV0YUswPEZSnM8V
rsx3u+qBZVNhmDnjzb57Mas8RjSnCzqy5OlB6fdYIth+zV9Wan8UMoEyUJKKVxOW
iORQyLxLHnF7IeY7dtIsK4XAIbsVzcidMqM0iAW6Qs7Nz9TdT0v0wlTTx5/QggVW
SichQPAY42PFOSzK3qYTh3HNN3zONxLnie2QhkQx/xPUnKrQTjsOZ9dqyARyYHi9
gJtJ2g3eU504z+G8M/22u+Ft92P800RN9ree3XRpvU2RmFPj0ukBG27lCwZTMlxS
58sIiGL0L/igDcAxcPFVlJXaLp06cEbiZcVdbI84QzlGF5+duaYkaTGHY+ph+ESe
cQr++Vd2oQieMKmxUYzO4xe66chrPabkoR+ZecY5JAdnlfVigDANKauanexpOaHA
E2ahKoLLRr8VAnS/3eD/7iHl5XpaN0j+m3IoTn5d0OTNbJeNl6ldbBz0SBxB5td3
DTRsR6MyHd35enzb9jHvWlFIO9ZpxISU1KO4SEWjLdtPYhZZ56NQgGejxnWlOBjY
sSrX6cY8t0kh/LP7Pinv5ATx3Gvo2//f3LrtldWMgsv5t5RJ6ndl2cNaG3F2bCeW
zWxWHA4FbDiMdrEnTOePDuPQCDVsTLSGN9YY4fpl8DgP3I5Fe6ST0Or6HEf+X5tl
N6OYEkWfaNc44lRlFDHNnefKT3Rkup1hkWn8XThOlCjG90GiLvgxsRLmGnPT5Yls
runQyzWVZAL6AMfaScgtD4fhJrEE45GsfdL88JPmeIQI2AXbXg7uI9cfUIgKCvnO
+enb5/nUtuXM1RKPWM/I/EI3bhDM7pTjMnpv0DAdmRHkvptmcbRMsUMqrCS/+G7H
8VZY8EKFa0SIKcoYqEHz/RZozNaSlJOb38yJ+wrH4xhtMm6KI8sxVmdJSslITXkd
7a1oDBJfXnDaYsw5QGKIBPH1wenI8ZvTV+yVyzF8MxlkKRfCBxwQYHKAmPJxwomo
YwW3qSKQxmbhVHpaVMAVbblU4Faj7I6Tm7ZZ2HAz1YXL09ERiUg7trUPEpK0N4wH
5Iihi8GvEw/kYkjY+pJZeBZZq+0A9XdSorWDkdsJQGQhshc0SuP5nfGchkE7Tvb9
UwpOfoF6BSoaSNEUSj5YntvM5O4TxTn19P4+hvkeL2sz1oHT1/rRbipnVBCgTGoK
RclOZVIAL5iqYes08SaqbTIw0mHINnax01uJRsfqi5XaepYzSrv7pJ604AHXtL4G
pylxnyLH40PYfYnZ4JnrbeeEqqAL0HDZEnOujDfACh4DoDixAaB4W7Uzh7/ifTDy
e/n90fo923LCOZxWy+BmSx/TK4Q+2q5YTZuk/bZzm3rwuiHj7R12uwUzqnlmbECD
r+vC+4fDzyO847tXkjBz+iZFBz5EkJigKjlWGHDLku+9xKTR1s7aL8gK8wIU1BgL
vF4Zx1hFY7hZfj9tY8is88/hoKj+V4Gc2PdkWQBSnX7KCX4823d1kFZC3ASBk2cD
tjrYsEe4GUYqkKibjVQbDiLl0WQqv7kzPypd9e92+nYjBjI1RLzUvjYifbSezrrE
calFPhtPHrI5ujmlADJ/YRleOtESEDhJdE3tgkxgmrrZJYiOAx3QNlP+3e5KdaWS
jc2yxbhum8JEak15SIDh/QlB9LcRpIi+2NlFUx2JzcFFlvc5hTvsQIVGcawVfrXl
s6ftJgo5VOsiG9hzzBgfkfEKAFWTNSLMA+NqV7pgpb7VZ9jl5bvBkN2PnX1pV1mQ
3ucfcBsoT/6REjptaBdjTJXbZoR3hlVB0R/NwRljuIN4um5zLc/DMfdWm0CW5q23
auvcEFoaRDoEWzDbXhKmsU30o6+e8ZZCVcJEGNPYIFsPrwH9zrfxdmkmglO9cucp
+tzBpUyCzLa+1DllD56ypMUr5U3UGkZSXmvmv081D8mB0Kq5TVXd/cfV1ffWWm96
nvl6VuX4W/7c2moHv/JoPucYlc9KBMXyUjSNMa4/eDWC6vQILvUvIJtPzU5ekqNs
2Zntq5gyM7rWk5SZCZRE4iN32U/0HwCJsvPrCkEOW/L511OB8AB+Vt0hiwZC5qpV
GKz3GvZWTudUzYIJus8nh6e00v4QdK0nM7Kx4BkO8j05U0lhUNvCmknSx7QnDwwW
AbIq/Tw9lyUa1+b4q/ZaMxUybRsKFNUlWHF7HdzYjin+vgD+JK2WYa2T9TBlOQZ/
6gg63lDv5MqNJLmXRUV0nAuboCyJpEHkssjVlJajiu4RjN9+vODmzTgxazJ/0uyR
5pF4ZUN3FuqTl10FsNqgfcrrXHV8uSFUpC7HZSVhbc9Gma7zbikD1M+IOJ0LsY/y
DoaegdwXWWab1jsm2cIwFIn8BspH3jpapHMTTdHMwpBjl/fGJGQ3aazKx5MD5an7
DOUVVCf9ZMFGXeOUCJQHuYOwS6B9FZRg8du7dJSW+xC95NiWe+4Nz4+9sVp2QcK4
fsMUS4/k2a+MVUpFL6HpKlJeL55szWA3r6+X86wbgESj/B7vXXJWD1p1JlPEPDT2
99KgAbQvT3653mai6Hd1zZL1d8nm9bP1qeUbkgfetyUYCXgpkJf5qnGFSln+jZje
bqy45OirBd1/mIcjt/TBchg0G33FyYKJHJJIsuohf7/YCD0f9LsN4DJYsjQ1Z2qs
vHPFF3cAFUzkICOoia4SPmgXOe4/JQugbPd8gJvpqCMJygsTFdLBOejyO1t1iHQ5
ayLLDRtF+bdTH+hRE+e0yj6Rn6l5iKRYQdqC4dmIPKIv75E/ttfs/gW4QUnJW27t
Gq0d+Ng5jL1lN+Ieonm9jg88hMI5SgyPiB4Wc69JBOMVYfiPLr+tktyBa3SlS+JA
OyR/wQBoLvDBWEk245dD71GDvu/eTq7S099M1Znz8keOeahHckS04SLY8eUPukK0
GUj70Wvy+mpP9jOKB0fVgEZtiwWs/fvjqyA5DmUfv9Sujkd60n0DbrnQqf77iA6z
Ow7DcBnazDp9RAHiMfGrsty8+Uro8KlxcpxBHPASw+/4rP0+k1+xQwk1Bfg4kQz0
zgTGvjMuYTs8m+slSgCKFCsDu/Hl/gYtS3LxSDli37BHTG8OiP4UVySgnChUoICf
/SXBKVMzrevSD/P4YRAXuKPUbgNZ9imbXKJZOmYgBb9Rb9ZFld8upnEFwRqRZiqr
SWQMbzQ0VOWGkdwiKFc/d9/GpLXQqXjAWYNlWREmTuU+3l5FnwgmA/MtqiLXnvY+
WtPkPjoFU+B8Jmv5OVEmCNfIOC25XQKZfMboKbCj0bw1SZhpdo3Dxkcx5yW7zGaZ
r16Nf4ZpDKMceCDMv0qm8OMM+b0igC8aRZS6rR0js3r9QD0HuDp1Udw2+YaYtg7M
dlw1K2mEmd2WSmbzbL0+hu5R1ec7rDqVofboCHNtF0ebJE6Xm8yjZTbR0sQwkidd
HWp7DRBCmurOdKu+ZKtPL26FGOG1FGfIHZvUFH4kPcpchJm8oyX6KvRiuS45gMqD
Ggs2IAneQEVQlmSFmpMx9pnKFyJ5L41xvencGUZi4UEs/YmwTRJ+xrxoo7kJzfry
NtmmCvrMrIPF8Co2YdxEF3VF6Ut5CV2gLlBtapX0QT9N6VfVj5lj9Py+tz90Z5I9
WOGaRrYUsz3HM0btbHWIy7cmGlefK5o4JGaV6ESaiEzrx5/9/cGgvFDD1Yn1+0qA
pIWgbJxEXfZzsIwyBJgVJIbSLf3xGO4JrFEuCTMxutMrAgF78XN5WWoc/LGbkeXf
9XmhXPztN8ek6jrFmgp8pK7h6RVedSeeeYHCqf3w4GWQPkYJOiwSDBTyHyDTheAZ
DfRrtgNd38d9P9TQgumXzNLdwrwyuuh9ri4yqxQg1bzWvc8eS3oKVNONhUuWKXqL
psAFnf5R+rDMWoy38cBNLOGAhujPHXjHF2IsdSaaFc4biggzPRgbTp7QOG+tt9oS
M7G+20BPz6qUA5P3VZNiTTx3Kzbyt6Ri8jzOydVVVTJeNcSjTRM8kT7KuMVTgP+J
pBMeTqwSXkIn4N5G1mWlrb5n3i4BGiZqVDAA7by7nZ1xfvqOBqs8VE3cTAjDHizT
6QDai5qS+cQclV8DZxbBYcTd0cc56tqlM1/M02rdWXn4g0uncJkoZZSmxzzCXC9z
tuvSELzgrxT/X3QqPEVvvL8cFnmdHGlW0AvVHyvbK8fBvCplX1132C0s6efPjaK7
6PZKGmEChCXOAT80ITDtG/dsGdBHZPDVMxkRt2uA08SIUZDTXLo+a35BwfuVfmqB
dbbR8M6t47vulQ6kngZ0LVTRmdZRdA3MfGIC6vks2lCWOIDGgwCW6fEASLQ9hPUk
6fo5UNSFPBAwJAOWgY6++5xg9V87eD1dfnnP8IgfQyUSmZUtHjizcM/QDiPWa2rn
68fqpxTQpZVAfrZ2ND6mANgzq71odrSAEVeaR5QYcGm2B7YB0V025NfsIYhcH+5I
/5brcQm4T2/aUTC7mCpcHAU1qb2QkihY8U63FlEvBJKNZ0KotTSEVIiCQo9iBsok
Eo+zfoIk9LsGkJiEUlAZKytP0p2bV4yrPOWftbP6F4Rwul3pQGca29jpfKlwJx0B
GsGkHAN9Ro+7QK6L65ESKlPtDVWRJzoGOp0lc2oSTTJQDS6QjK4GceNKsIGYUqJ+
qJlqit3P/XLOps5jJnE7xOLaOXe4hwHoa9DD0+/Tc30kW3IYYQwsppiNBo9vxm4Q
6fpHGwsvn3CtI63puik52i3X11/Cl5cpRY2F7WJyKyKK1S1yE8fazmhubcdkcjN0
HloUgDTX5bZ2A+hYi13BIXg8Z14bqvdF/geKFogMhRlWDyUIm6PJ50fbpyMdouCh
CbXAJZpYeXswfHGfyN/HgouGxGvyRdUB+1kvZ8UJSKmFDCe/clFqNB5RiqMKKAgH
wQQbintwsV7KTc+ruCi2elWUtm8Z/W7gs7CEYnlcU4E9en3f/cms6yUmt/Bxv5Ew
nhYGnYNpawo4sUshU2O2ONDKO3hMhmSgk0MQQWXTj0CWgmIrefJbYCKLcUzgNrpb
bNz6CDg0fTyzlpNCYXc1BmHJ92LZHOy2+9Andjto6nSJTV8ZPIC9pP1JVKg7KY6E
KLajDIZ38NPnFp0iCXI2ms78Nu8NKuBUqmm7OJQuOKiXvh2IM70m4YWkI+tCqIfZ
0+55av2MyDkJ29quw27GdW/Ka5ZqMv3bVTNN8dk4v/7kAfE09hZVeFSkQXygCinF
fZ60PUqi74ydasbNS+dBa3k8LBHxNJ0pXGbCCoFww4CkizRU2iq4+ejuGtBOB5tT
hKROQZy0Q5eIW+xtqAvAG0zITi6gL/Vyp9gtpNb1J6trnWD31mP5czqryHJDCATa
xncwgKruHgVQg2MvqR/MVX2JfPnOWMQ/wWCxpZ9j8ps7Of+AbWLujKxteE1ilCvP
Z2LMX4GejQfu43Hj5phXfMi6YhmXnzX4Pj6THuotUfnJXXVsV+Vr6aJ96J+ufh3/
ZzOToBQdZkQpqqW5if6gn2+XM7TXeQdEwAFdM+paZVPFgiN+QDtqhwLbJX30EPOC
vW2vybki4UsiPydPDWVtn3goF+GR58DqBy7MiOpeuSGcXgqRuXo2eSFM6lZwbTGr
n8xBBqMfJnslrGqoS20Qq6r4G6+FMJdBkW9iKFhAnJEj1JNC/4Rk78o5FvsqEfy2
88mXfulkkP11ouQcDSbBoeBl3reiNP9gPG0+VzwEjjd29Dj/NZEWZZiSmlyfZ/iH
65fYH0DPU+wH0fkIdvb4Z/NocBkg7yOYlHDPpAASK62qsg9uQsNsZDJ6uu/Bic0I
2XLB7SPRXGi35QysYnc/N4ibXdKshSD42OR0syaGEHdUJbz2FVnoLK+G5hPcCfOa
/IxUJ1TH9uvtAsm+3jH7Tf5WC8+qGESSf/8WKl9cvKiuFY5CY+2x7xywXNq6vZB/
U6VIGubMMaWiljHxaf1x3Vq+ubmQi6Gp1EL5NU3w/8pr9MY2IDYVVST7s8Rgdczc
B1apCWONGrhQn7HWeXCfDNti8LqyNMR0aHkNeUP7baHh9cfEnYoRvl17r7Qr5onB
Jx7VI/aZOQ5fEwbf7lxI8Sdps1tLEeqoFdqQRDNlfRGfdGy/4unsV0Nc4if9cRs0
Yl0evDmnbOTw+XBnCLD6lnyX3rV/z9yFjZJUaQsgYyOJM3GaLoxmtBpVDa7XKEGA
toB6YrxhcS9VXeWcp167wkKbOPA5tKuha1+Z9CHUWDN8E+Pql/djNiyVB4l3REAW
mInygk2T9EI2wV2KmUFHHlB8qa6UX9AQuVIgWJxguRDWZUdnK5iLgPXX1OmQtnyf
570PlOcX0DZSvz3hZZe1ibROG7QNlMDa/MaR8kOBpHcxqOH9GhhO/E7SBUh6GDOd
ruI0gC3H4OsQ8PGBqC2qVZOlTXT0BX7mxn7Y8S61/ohI9RJNr2Sdvu3UBDIV51Eu
OTFKxXODpemJUXDi+ceX4po7EARFqLj5jwRdZ1Vi31yA2Y221LpdeuL229L2YCAa
2KuqYz2TXg66c+pM7pZ+iSSfMM0tCEnC+Kj1ZJXWtq/bTVgXOm4Qcgh2ZVpaxXzN
4pnQcMfCiCwz6elKog54QyZLnHv+tJoZ2xx0v53hrZOvqmyJklGfWZs/M5WFafZn
ROYG72Vt9Zh6A5kR3E/+k2+BGkob41Ja1uzAVZebo8zCNqRq6qyVT6y5E4ZB/GSt
TqdDcW0Ka7vTEwJ22cpezrdPGH8UPwqZMBbGn1O3lx81n4F9PmzhQ25ZysXEFSgf
5h6/KFMqEwFfEzkFW1bkeXwo9YOfJwFG7nIjBD6wTAm4K5E/Wp5oItG4qcAZdp9C
Xo8oJKYMn65kl6nQ/7QDbd8ZI+xB8qSFWhIAfkpyhyDUNOQeAtbtgOP475hb+KYA
1FIkVkQncHkHOFyDlj8ePzOnFlKs3vPVu1/7EPKoHZduvc8UPcvNxYO7tfBR9CBu
QSDJ9iZ0nfVosmYmU02uiutadhgfcYt/7EnZGRnGRWkLrsSKl8ELlMpC1f1Tpc04
90coucRSGaWS31siEzBbDcL6Zwu+U8FUfyF0X9bgMQxcCTTr7BCz4zkV2HlOxrJm
8YK8nvIvq88jMD0DRRru5TPhzy2KdwgvdYOdx6hQJqQxGsJT+zr0WBNOdzhTSOh0
FMCuPuGvO7yWTw463ppM9lFU7AJE4sE6K/CksyIVfFdjI1whvfZlTM7ckKA64a0v
e9Hmj88uHgNw2BQU5QLO2ThtEMWG416LkFJHPLtEJe9qYUJtuGvll3511mnP9yKK
Ygtgp/qxWf+SxFyDCavcXFThzmBa0k0j55uXKQVIhfvWk/xvvNzirZmzEJdPjbw8
bSvSAN02lkdyre0haJMAS94ylBqBRH6zbusFaiD4KmYhi+jaqQmB8GsJGxUfmDqY
AOCud9RW0dPZbSHWGcOYShpjilLkHgHfxyLA99f3aIQMnbyJEImdIxVHErlXuKYS
sTh3wPQQet6DvdN1euIUY41VBcaEiJUxEFUzoHFSpxNFzZhUa+45cu311RIPpXxF
uuWc6vn2z/l3Lcxw6HePKEcElDpDMKl+O4rjxd5pYGtJ2ElbV9zzF5IW2m8WD/2r
UMue0TOaHEJy+a+0hiBklcMG0v9ktpODJnx6tflpztRfFuWVgXht2q4cxkXk4ZbM
qtIWIKB5e5SJgXUlLL8WRz3/0o9XpMbNNWU9JsjGOB7QF5vP2M0vWA64w5PiEZZg
/l5PXxOeg/3V+pxHXHj8NfMKEjNymfvDEPAdV7g2ap4r0jYUduAydh1OjnnpBWBn
vc4XPvci6RKdAEXea4MkS6sWGQXhc17P2LV2Lh01cXKyYmKwL3xf5JKeLfFIPN2z
ZpJ/UBsCJRlU26slKQ6VxHozWQ2pychL7sPL/lTe0NZptL8FfPie5yhQYXb95qO8
qI17ofK1d6i/h8r93Mejlp+DGxdU0+hrfDPSwnf/5/cdB8OCdJ5cMrgEDcxxpADl
0j8hznmq1y4XGInUcKru9IPOe6D9G6TZ/kpmVbo0zlDfEW0hEONe3e0pgO9xDjIh
LNSMBfFrW87Uh0hnLzjYbHqQCB1lRV/cowuG3vFobSwOPMx7BAWKkLt7Qs6gvo6N
qnGXhkkxW8DHdshGR7lmWaXFcdUw0jZqzn2SULvm4jDu4ZrJVbgmNqS8rOFEPkyg
kmlqW5qZAGoDu8V1B3uIO9Y9PiX2JNVnD2BMNmSr4ntP958wYF8wgRdUYn1RbSYG
YWVvu8vGZAkVm+/wI6Auxvaex2UHc+7LdUPsy2aM+y+FX+L0Am29YjWtMIM19OYX
QVqiilxf4Y0NbuAvGl6rnttSUKNrcQni2SzifQcbdBRO3+BxZ40KyH/BI6DEA5YN
iyor+oM4tlYAx8n5c5B0ON0SRMdfZE7NTe9ud3l7WDEszGAe+th/ad9ysXjFyhUm
jcm5qKaSdecRtvOIlY7Z992M6GPu61XaC0GJtY5ofk4QIXH4gVR82FAcKlmKK2Hk
lrlgA33Nnp49O6Zll/X7O/nXnFVTCankBmsmL/b5StoaejLbSe1n1nnCoGk1lC47
jg3kWXuEFfgpSEVCBxqUQ9ObEd/j+SQ3eCQCjWXkKnrpTIh3X8U0bQSY/sMpD5eF
XXKXDI++8jVKtFlhmsE1Ihs6CATcoldv43h7BnBHaUkFmhr2O2/wGwRnUCXLGm6h
6JtNXY3gI/BjNKZ6/kmGibpsD7eP6XJAt0VGGpgdzb4o5te8SnaEBMBNj+NN4h0J
WjQtTt+ei4b2YpNYCqtVAVrNb89aaBHSGKJ5gVtEdEgMG7KdzCqnHB4dL1gW2lGo
8jMWcWCmw/pjJZB5fkeXlap1p9Gsco/ZKiye5J34NqaWcaUYhaPBWO+WsCinNmpr
AGcn/DudIxzVAQcvmXiVXklTQ5HMern/fLjJPzMS7ES96tnDRO2hswLyXbF5g0e5
yYcsncsbBG6c5SSYy8tdwDf0+Iq9o7e7kuQj/+WkhxlramBk/K7L/YSZ/+WrFwYm
iaPSg+JNvdHYgBcZW4hiHYW4OmRKLA6V2gD29PI+rpvd1k6NvbCNezEzEdw7rv3b
pJVhwNMjFAzJmYRS7dALkkEo72aVuNVimquDU9CWjTwGh91WnEEGOx6ob7wn67ZJ
uFfDEfQgm9IYBpaG5mA1HZuNytS8BZcIf8uM0EdcgZ791F03jq0ItYiUDk5yO7tL
Z55zYTTqhnQNxW95ukCluBtrCgEyvZY7Z74/3pC3tyJJ4pO8JuOLjVTyJtIXqedU
JLwQBYhxcC26Rs3ISCzjUQKIceVyfliOMI+q38Ia3v0E1JDKHw7+TSfIamed6aXO
vXOa375hDikxBZzAfsnhDwfUdKCTs/dzEJU5G0AH6KOyeA1hf4zKggMOq6+mT65c
RnClbDEcYSEWx3T+PtcNYOASZr5JDk7GE+wTkk/HzX4Ttapc5HCGvig9nHUVYUxN
41Z6htKNMHQHpov8tPJIV5wQ/VJbW+OQtcYd+7kQ9kJaAzEe4iWBRUZZyifhb8Pl
fVKV8RySxMR4chY+v2zXORrx5xj7WHa96wne7K4rEHOqpgvecbYwIHgYo7OhpDiW
t9QENkeyU5lMOzVGrcgpye4lwQFQuT4j98yIeYCnfGInFmvrxfI3L2FV7gQF2EDs
e7lTwBEG36oSRQnbXnGRb1cP49gugOS4L/cIgiDrM8yuKvl/mG6vgKTHil6OUqct
/cDhMr9rT107A2EEgB10OprC4hHzyKZ/ieKq5v4Xeeia0BAnh4yCYr16Vw42weG8
S3B2tJhR3/xhcjGCZEe6rJ0IkkA4fdeRR2XC7t487WYvV3d6R7D111xfnVkx6B93
5ar1JiUiigJcYb7YUZKEmiG0fmnwqh97tQEAQOuMkuUYd6Tr4MkiEtSxZH4PNo/d
8Ay3ep8R491J0Sg9pyX4v2UBet8D9Jzsjo8gNejKl0X2li/a3J1r1NZHjBm3hA2S
72JtG3Q5My70QDcvenJoDPEqtdHBqjyBJggp2ikEl3gyo04Rou+kWsPsCCYE0vO3
X5KRk7/e4PGREx0w+XBEMzY7AeogOauD76b3Tk31b+4/mnYALu4utziAmZMruRzK
zj1uUgWzDSl5XRX87Nihs2Wl/b9rHB/RvdYEt/0Zjqk4y/d+AFtVH6sazzUjhC1I
QrLTdPeObdO2a8nelkCLpTtw+m3Kdl+TIHLFd3KdHbVXUjjuksUhho2+dnaYQEQ6
qxZtYYoY+I1vfwaI+n1ComnR9PXiMpWWTLj1pVq6DNWK4Tci+oirmBjp0/tUY2gi
bhPXZmLfmKIXcdQJETWB9NtC7r4airTHeJY9Ir07k3x+VgpJTUmvsUF50kJo5UsL
sts3PLPUOzdh70KtZMmbsAM4lxISP7YG2iEMTuz11UsZCj3Z/biT+nKGEU5pMIvy
s+wG9FWucw4WJUZHZFn7c62WvujAOK+9JWb1VpVzhysGG7bl0QS2RRyOo8H9LJhS
0u7wgINbVw1+64ewxGOrVJAxSI9HQDexZYXTZgmORGGKcpJGq/TjP6lpmMYq0/9o
mTSoZNmUtdbaPCXLc+UfTcDG7I+hdMCtDT/OPAr4mI28yKLDUcUGSlj70iE9pOY/
N9G1naGb67fXz1qpdqN6s7lfhxcI67sV3aEMKbk+Z0lCvKhaANrHipanaTv9xP5f
q1ygeA+sygw1bS0BVMQTUg72+0cjkhCBWru1omMdYdhAkkISX4CJGcgmd95gc0kh
x/THyysFVC2XnrZkr/PZ0pxsiAvPUNiMS2ps1L0vxHHimxccCeRoFWeShaDjPNVy
9eSOkyPMVwMz/0kqcNIpDBUYT40phfzcGCJTrLKjkri+fXFcSgL41C1Q/KhcQEw4
21VFf8dC9boPKLGtkDowPjGV6Xw3/sLPEz0+0UHgCWOTNtN35MvOygCrZUMZ+7V2
2mQAp/dIsPH6fcnrCzSB5SfHbBh/Ir79/EHVUR7O9Z1uNyTfznSzwJ7hiuoMLdzw
qqJe0TTLVu7HwVY9I7yfZL5f0d3AMYBT8/4FexqiXN5yicfQQLCFU1Uf07up+p7y
yU/npm260uMtt6km3b5uvbMEX99PZYkZ/QIIU8Y9HFjGQQ5hksJawQb6UZv8x4+e
uL8Z0jHmHjwAmTddwX6blqgUluDjAxf+0X0NjE5kvIvWPlZ7ShHYw8kCCnrzv4/D
/b8zAV7e8+tauIpnULvQv43Dq2I2p0VMHU1oEskxBFW0dRO+b1WyVBDnfMHa95Gf
nteVMEUiuBF33Z27yIuphvjP0TuOukFfuiUoQ111399XjV5zyQQAi3eU+GQnNYIr
/yU/NpKtEnWbddZheB8OMU0vrjCtr+yWDPo/JWluowhqAx+fm1wd33Cw1mhU0MSO
zSS+KXjLVYeBrGvgOVh6nupMFQEGOOnsMzBUa46XDOBMxtjVyaLUtvaJDcufHwcJ
aVOgz7wfhwhgRwBAFwZWzx7HntXoZMrwNDyehw8cBC6Q9tBn9AE8PxPI/C4gvBbL
JFLK7iYtik3NT0couAkcptKqAs9L7jUo81ISDDCATf6bDBBZY4Xbkgx9Dbtsiaq6
aUH1yE1YIeayhmJNzddkQGM5nsEYov4GNdJg7Ycubrs2PiXo09LhtSP28dvuD3Ir
+EHQUfk9MHp7XkI9yqF0A1xEOuS8Tn42fdjUP8Bb34W+c4nJ9gYCltOglzXODecM
fvOF6SJWYs5Yb0davdqN3dkn8woRsabYZpEVxyO14Ny4femn+G2bQEC4OIJsIG1K
2axpQ9YcVdAu4M6YFjYhA8m9Jyaflf6iwUULaUFMnl1un+uPNwgvw/L9w5AmdLh3
txfRz0mcKbTsawo0YFA0RkxP4jl2gwhwKtMPqTUex628WOd+tHZxzu5NlrhsKltV
OD/GQa1MVWLCwqQTh3dqIGLdlmP5SIK+uGs6SiiNkTlf/Ea4dHVUqWyazUQXjQFL
zOh/YY7GO6TbgSC7T2MtHKLBPsvENBFLUFGSqd4cSz+hJ/rY5YIV2/4QLGXYx5Nf
VL0pEFIueVXq/H1lfyhZ1qC1IVBAr58rOLJCIpKatYZvQ2HNjnaOeNdpP3aGRHab
MwbW7qzuAfw8FfKBdXEepcLdOaGBYVTVOxtW3GVUkJWu0fTXa5u/kL8+OinL3RvX
fB7JjehKnYG+/UJAgY7lYeZF7zeKKqurJ7MlU6ScjV8yppJtWFWYtWz2jJKd4Eld
GDKlR3/EMdPDSglQJOeOL3rb6qGZnvEyzzENWbN7dedgX85wrBadcT09KXSQmvI+
PBPGAGuFHYY+7HGeNG0fF5/Fg9C1xm7obfPO4zo5eXWA5b8gZlH7kwQc6Ewxnlxz
q+k0A3iOJKykd1yUr1HwcaUSW3n19lxZhCmjbIHEUfbZWxgQLnIIWQvZKhdBODx+
3wFs119FGIGXdemCEu+EaEt/e2D1WxdY7dQJyNR2wRzVKJmGe4N2nYNPtWpiyD7b
dxR+Owbkt3oc9SF2XyjXy+TqTyVe56CQtLTFFxzwTSErpUsg2koII+2Wrw6JN6z5
uOkhEc6NGXaAComBjnqt0OMKyIqNh2cf0log5MJ4SrhR8PEpVxB0XcklAm29fUHZ
1cof5WjFhrim68FLlndLu0a1itRTa1gZ5+rAd3ViChTtAyjTNxF9WCYtPt5s/uxM
+AN9rd4e4STh6cYyNNTDpQfJ4jLFCiq2SVmEYIlCdBBqw7OCuO9ks1YppNqZ33jJ
svduXRk+8ESGN1CjR8Bnbu3741HSE4dAqQ2bzzy3hAkiYCaW3prQPuA7QmZIBL14
myM3s09ZRKMhA5SaVnZYVrvqnxoKLkqzNBa7dlEoTatunJcn92eX+Cc2h1zOZ4AV
K4N64B+D486Zd4oPs8vvpOZ/IfmZoebR1iympUGoYwCBWjVMY2boQhlCTUXE4bTl
MIjVomaQVWkQNKXite0JsGAYAMmgRDoJoDmayB0fZB6DvrmGKc+I9AGA0Ot3jjGP
PfANT3QY+rGVKmlSFibhT9p8/dNZqzqrvI3ZIOyjaAHAuQfsKnQ+eXUSqK9bj8UU
1VJcVJ4GUxjJZc/woihgISnhYfPFKWdcVlpSiUvxzmYKrbgijdWppiDRYJdNMiwX
LhzzwEp7WPECfCrU91jkcEY0ibrUfy40zyywXvtSS9tbbIi57A5MyjY5XfmHXSjL
y3mcWQjU0z9pv/2DaCXTAV4rK8WJMoT/ZFKIy1SWxxJEjReZu9uyQdVvIbKr9g8e
VaTAew6sHRfUGCj6O/Sd1+dHPM2ChTZql7ODzKBMZ1YkhkfD5ja/sY2oymN5LGB7
QO4VjGfGKttYy5jaYGEYv1+lvbo/YzJO0avYhXRlWGNFGfw2rPUWAmzaB6u8qJ2N
Wy4YGpTcGBNg1tlepICKrvi3sFyjiBb04VZWT3RaX55/eq9qUYwrrAM4N75EBxO9
O8P4zvJMtuMFtZghhZX9NxYS+JbnU5t2X6kURtDcmN1pN6BXxn/n7XQiUKOskTLm
Sco3WjecsE38pkGdLL1K2eMx3cJplaP5xyGqWDa1d4XlrilKYXZWArl0UBAXgIeH
g/kzPOr9zg0CdcDhPk1HnTrQ+PVZyeqvnVrh2XYRGoJj1Dx89O7qbKPBczV4Iwfn
0Wtl85Wa+C7AGcg3QEOBLzlCUMbuFpsADeRMnE1Xs1rCHzV0nfuo+mDTnyzJWCTP
KQb9j6MvA4ohQCqHNVPpl71HszEaubO10LIp4QuGa4O4mawd+5IkZ93p6RR8QeYA
6/WbObxIvkw6eOy7YoAl1C1WTENE1PmcRRC5X4a1LRmlTTyIiDT4UN0jtdx2UY9i
ICtBOihhPwAj56SxlSrWcOb469V5linfIGXOOKI6WxviLW2rl0JwTbGE9YN9oWuS
XU2JnbQvelQAmAWr2qWwPHUDOLO1UQzGEuts8VGvuMKysMpQtcIvLo2NrMizYEz0
L1hoBa5BcG9ni+SL1GnE0/JCpBlxsXPeHC/DCZddFB0zldFYad82kfdud5SzflZd
TXo32roTqrN3JODNq0NAK7Y65OBpW10vdN6VgUT6k3w/6MhPSpY5fA8rtAvlL9lD
RnlBLfxe3xp0AYtDtgZ2A0deCUi8Zd5CAYMgxxJZ7NnM2J97P2DgupP6C5l5qT45
rgARv4JgVHsRyMIFokmDzae/P35kXQMCupcY3eK+VMEdOy9w1avcoQMhahagl9dh
grU987B9eeOvJmMNmb05k82uUCstSv5eoYp/CdWl9o1e75k87qAYUekAG/P0Hwlm
G3VKnoWgffOpTquHw1m00FbT9grxYpcB6g5V/OjuJfrsMu0YbB9IYLgK1Sv9Bdh6
Zydigum2ve3v8pVBOK5G/08cSTSYYVcD0q59rirbDRwqAnCb/s9KbwPqV7OMYYMZ
ePI4rJ25DGDb+wQk9EQQD3lzYG59CNXuGmTWZzWAsTWTalkRUX6Tyd1MzbaNUUy4
VKKY11C5yjiNr0te+JIXE3gFoZ1vWPOwmnbUQkEEpoZH6q90SA1eWSWiJcvvdo/l
zVe5CHpwG+r8yry66z+RFU7Q3Ud59DAYtN67qRkYMCW2jav7uC+woxNYg73PiF8r
N4iUyADM8yLV70wh+2A1t5Qj6c2q3R8DHrjxSseM4iOacA9ZhVC+eAs8hz/0Dar/
zcNHfGn2Nk1bozEg/iI1SmhPF4fiIzXmygnoqDAmU6yOknDsQpbBWUYMar7ifa1X
mWvfiOm0vVtdaBfdMwvRnKSkNbMRni5PYsMnEkS4pFn+7A7/GDgLr9f6myHt4Ssw
lN5qzj63wp1S14DWOw8JS1AKKbMuJ+6wajyixvO3YyT3l6bhofCsFnPaCvRTGtJV
fGaUOxjiN+fVZ0hvVh9b32ZNctxX4w4iUhdcxn3Qq2qMEMrNegYCs+lHQoGqcWN9
V6Azm/TlpAuQ3l3Xx2IiyfKpT3XnNyNkvsdySRyA2zgQ03hulX0dNQ0cjQF4FOkE
m0kHuqbey3EPE8hmtsoPo221uddgbHuK1WLcE1UlEo/51TbAt0TqNzYC3xFiUqIa
Zi26MhTR6Hfa2wJLD3qaztq9FHOLhbgyTi9EcwLaLTPLP/WHmStiY9AM0fbuD2DF
F0znGv+xLNVVDi6x3CWizGPRErkYfoO5LKQblhkCM4EeVWmbYsiDjwP9zGCTqUUT
KbrBp5lDg2vzOtgOSyVIfWPJ48uyM3nm6VmXdtMqK7ZvGj4G/X8NM2UNIBbW9CZm
RigwgWs/8ZuI9h8SA8O4RqfRupx8oymRmWYDrMPu9/KfhpxafZJB7s3ERsZF+x55
UXy1J/tEj6/KscE84IjqdUeVLYvH55ZfTPFfmKGj/lMZo6afvCwKgX0eujubDfCO
heN1d/ml7x/jYflP4jisQJHRdW1tb0nDbbYMKYePdgEPakKPtahwT718lteiR87Y
SDwGZ7R3mylvezE5h3a8+rrkWwdX4JDLkILq/fFq3ZmmJ/LgVQtU8vgVzgZp+jOe
JiWNvkDYIqP0gMYEDgpq+tojlatmbDxzbPfeMuReQm70mFcmtFlkQcgT/Aiu1O+W
JJEqCEM2onJt/a00vtR8n0Rb67iFdRu/NCJA4ldQZbr87kRL4N4YbZvfyBxe7HA1
ZnW60w/t/weL7N4AHzKm1kxnRRDnPmfhV3Y2i/0FEuvRRIphBzPAZ45qL/tEc5ys
JWq2cNI8hrYXZnofdnaKHuZ+op2AR0OGm8VwhRP9aqmcqe4NBx4r0SUmIMGoxbxp
eurYDwcO/8ALSaYDzI5mihpM1Uits4a9YYZC8+UgeAV3NjcZuwfS3XWiYFWqxMS0
Gy8u0RggAJYGavdkjq3MipQVAjoE+ZJMItq50c3BTJiqX0gZZ+1GynrPInlCtt7p
xHFuQ1sHW2sjAAs5BRG7WL5J7SO9rM5N0f7pH05CmEAMw1uH2TwAylL1EDj4hRG6
CGJuxgW3GJ1kQS6bPL3lt+MUU/6JjrT1qyc0mD32fGS1V8AS1chd+2SiXiqPDJGP
GFQYcfzSVvjkgEz1GyI/6373pX8ieExLhgKUSm6FNG9KQWxMmZBJJU9RywcmTqF4
5eKxGuj5Fb/dUUY7iMfglAodFH35rUZZAKxlaTI+7XJcwzXrv6l3fay0CKpNMiOu
25/rcliBKz+Ac1IGffw34ewb06IPMC4jCVnMQL4PLUl2GwVDavoynowF508tDXJi
c9DJmCpfO4I3Nzqanbq3xvpHzKYAMY/6leSKmfZwDMu//UuVi7BaGiLntVqc5sD7
voCMSpzvF8P7wu8bCKA1d2jHZxAinVY5RngUWZokrHnJSVprMKjg48DCeb1AzdWJ
1Txn+w9qEOQnHKnxySSBuGX4s5fiw9VJRu2vPwiFkP4XDrMN59PQIdWfa7YvFro8
vVNiq1c6resgihyJkNdzFIXRwvkxX+ZQN+/uBPz9CPMxUiK2Jj2WS4/vaZ6kXWJn
1zTrpU/EgN2+9oezEPUkq+5FikULx1G40GwvM2KrAjbDvFYiQ03asndUwjbXsY5o
8sgWKHqHuvS6Vs5SKtvi5h6BEzOiShusUBglu/OyiT6MxOmLku+qrsbigiHzD3FI
wt2JKl9Vps9n1TsjQ3xF9FhMMfN4eLf0wGUKg0VxSrtrzjcEa2xxDLwGPKT9JcO4
BekNgOMCNfG1rwqXi2jiW6alyMdENDeynOdrVbwuUebik8XsAschi90PQ1OCv0AE
82Gdt8CB2GfDkTUGXHXoKvcIndgWXnceZ/gwoEib/vUjrI4dtLWpkHkM2s5dOulD
2lthLe9oWrLu/GABHDBkVq1lGnz2iP0ML8+GCglKHR8jAEMasowm/YHTh594Drn/
qOJMIQ7l6AWGs+t9O9+CgEHW4kgf9xzJjZIOH30mmBVwXVqnoB+8howZZBKl5z2c
rNvzYLs6rplET2bhxNi7N06BtBGAnveAh3I1Df/nkYXYPUvLOG5zwAI8IqvI9IKv
mU8nR2GXY9uW9LzsB9R9XdEauk7CDLfMOPJPxtf/sw3I8ov9UmRs8ynmxiW95Hs2
tBDvfI7BXkAYz52BPuT4eGi7P7W017oEXu82oaQA3z3LRniiKMH+yMIHQV3U3j0t
MKWXTpORE2FdKBJFl/dlEiq3zI52O4MlYCIeCfsl/Ry9U/BnOo9qqVDKChFWCCaC
zQrK8axAW4+sJltHXMpKFUDHfz6UcUJ9X+DEe/SklEh1ac1TuqaPWRU2wplohj/l
q9fAe5OJszxdmzx0ffUakx4fY7P8seZnA1O8LdFJ+hm2kmzQLvv+9ghQ+mt7Sz/a
0c5mBg43MKHVFt13RdA00hUqNIoNooB1JpoLomHtKwQ/8+86AzNbDI7f0BxLa34g
ef7jV3ZoKuLWFYGIhh6EK1W5eoftQQLRg9zIZlZYAizwBh7maK7ZIw3bN16Vvou3
N4lAeEAixjXbw6ebY+CIzYhxISNyZDohFvQa/a1fTnElPB94QatTEVAf5lopayNQ
eI+3/uoPspu0BsxEysw5I6za+EYJCUeFesY8MU2HD1400p1LkwfotG2E6nmBLyjp
R6SMtZN4ST0NQEY8TU77j4aRrg7lRo0zI6/71x3CI49cCNx4N5XlMTbWY75+LPp5
wyeoDAxT+OrSOjUevNfRNhX2HBCC7y1q2DmX0tbDo6SvdXJjIMPA/kUlvsqJNAq9
O2A/PDisopmf0irPLEhiGpaA+g5q1Q17kmmfcXBCaEhprFhqWYgFUjQkxFSIg44Y
5nVPjsw4KDpwIcdiCZSDmqTzDwbwlpl9c2w9lX4qvswzAYX+f0VZ1MnxGJxL6RIj
dipcDUuxDvGGSFKIEapf6J4sMI8+ta5EG70liryAS8vsVNT5BJZPfBcfn4yOQNRh
bSXKBh0hFyxFjfmwSzXbXKW5li0MBW6wxHfLgOz2GwThiEbTZc5ure3i7tjGCkcH
dxcEAdsivkRlZTE5UZqef4hc1uOcLZipJ8lLyAdVifADXMd2ZTietL4a7W17NamP
vTa2BJxAr71MzSxMrGzN8+itPT3E+nonXWgqTMTENCcCqoolpXy6y6l2TjV58G9g
wL/Cj802WoPStpyPHZHKpmcsSMvWOoOzvzJdinJiTF31Haozuxz1W+neAAQ3dYCv
FO4rPCCtd/sWAFapG0x4hoQUI1o6eA8Vsu0TdgeYBJ/jfCqyqG8eadw2+kUMJ1II
VjQL6Tuc2bmXesBrLDJST6ZUfDDLA/RP+cvrOVWzFSyyLK4NpQfBLwZTDlQI4g1e
/iRD4VAbI2RijQ/cSEbhAOd5mVIlT0QfdGgeyMwZ7rLlYXE1xS5+Ho6fwr2reslC
els7EoLxu+omSwhwDhPCafLJr9v/HeYNPGojsvr4AXYo2ga8Lot2aUbbpTnEC8kV
OTLN1/sz+MXaf6iMUk/onFMdZbA6cvUhZPjoMXLNRnM+LqQ9ynZClCThSw/D0P2h
D11/etM4CYalknn889ciaNlL3UBIWP0t9mABS57auwvdeOJ5yLIPtBrc5uivfrk+
G1YbObNZLopjRRm6jQdtCOGMddJFthieLtcm0X57INj530lMSxCLfTIRvGFPkaBH
ImuGGUUiKZUi0Hld6dTxvI3yQSU9A0+sseRs+lsamgaxEz3x+MV5lwC8YWaFYZe+
W2VASygAyJlkeLSz+7aFKlrzRPn40CF/UplBkPDl3A1q3psPYInyS27tyqHa80s+
KEimg/Mc9d3NPutWa2MNDqPaO01yxqK4GWoQLI0bfzrIlX6cMhNzBojJlasR6Fp6
0R15LRXFq+dYOy0D31QifWjId6ubxAN0iyi+gLQcC+RZbLiuEkYFKApm1AQE7nMU
pUHwzYkO3zqoXVK2d1/5/bcFeCaCCJfcPXJpBA+SgJLfmQhAa5VcmoVjT5UBqi/E
y+P58ZBihbJ1s/AScnSaQOrdO1r0kWWrKiewwtS5t7chy5E+5Kbx0Jcm1aHzLFNO
XUo5vKKjEb1M6nDxIlO9ZK2VOX+9fdRDqQqbYkLgw2qPsr+BQrcfSil+690NScD8
aVR6wpW9Is2VEMdFOHEhZjF81GZvtUGjiKlct2HYaKOQ6Ds87AhvQOlvXA2KAlIS
2HS0vvnnKo78PeiXYVfmplosbMPGSgoQbi0pAihrJm8NyzDKulDI3CnbMnqP53iT
LttiAb21DaHVBN37Xf44LfcnVY95vUKupTnEWjBiO/MLI2L+EFU2E/in2aMeWsQL
eDoCFAHG/A4g5kVe+CCwUgRGvQf+WhzRZZ3HYuq46RsRv3qHsvoxDL24BkQBDfTm
NKlUoEIf/00OukDbuXPZmrftbrKBY3y574fRIeXLEBXd7s/nsF9uuHjhbQ3WTgk+
S1vGWQ0aTnvUtRQ1gfXWI3IPJr5KiwdWFa3MVX5epnWEXyHBGyoP1RxTkd3OcuBy
xhhA3UxCLfF0qsVqsk/u1BxoOF70uo7K9TvzsRZHtcbWIoHqiFisIp6a02i5zs0N
WPAVTOD+LozVGkkDV6iDZTjwO/8YicSah8sVKdsOGYRD+Gc8nJwTBKQbM0GQfOV4
L2AX0E0VZFySPaf2ZzVsLJ2hjC+Nyr8nyCO3nysBItrICxyVMHOByuXKbf+EQewu
hpC8J8aOSyWnrq1XS5Sbv2n8eRSCoWmHsxyQ8Fw0jOBYFQkqRBiVbIdX2JMcR/M7
qOJYo3jRLKZUViR7P81/5WWpnNURDOSqBoDpck4Q/YnYubi/jCQaSb1dHqwRCwJW
mFq82+DGr+YHvAtJRx4msoACMr/r17f533UP3yB/x8uR33iKgwr7B4hxCDFHoUgq
zMgdmLY0L3G6r+N/CTIlgbSQr7yjmN08ln3QSxjvbYhSHveH8sTliTAhb+X+f0YX
+6TXj/INKTplV63HMuMWc9Tw57S3BJv8Zys5ZL6BiQDtIPg2PoAKtW0Vk8D2BckK
s2oDsjHCsh8EHUas84dVD1f8ghx/u8N6yIvTMN9Llukga8MP6a3BwcmsM/5idesJ
1G9Qqt00mBAIwomsZJTNZGpNomNUxl8feyIO/CQXsPOOLep4lRR0J4Tn+3yzHiUE
s7y/P9T99gad5UB8cgWEAh6QfuusJoLCEN78otm5FfJPS+YmXqypOXtKjsH18k3R
Kn4wGiuc/W1QwNlEqDqJYHy9NLll9e/iFtjZ/9LkqlML3gVxOYoQiQI/8/AmYhh8
MAmHiHq0f6mTjsLsNliOX8JDL6g8TEayHmNyqAgLee7GQeZ43tLDjZCwdi34sukb
As4QTklCil9J3kSvy33u4VRFJruwHN6DlXbQtHDHYpBQHpRgrPf8qnkzYiBiBZp8
ntPeQhh/Kzv6rji8t8wk3AUdZak7xqW7yzeHFTyQ6hBHsQw4zoxYqlRe47owr9Rx
dZ6Seh60URBTRYLEKZX3SavQOnBkB4RD/Rkl8HYl1RjLyaDvyAriizel/qwir3aF
l5YVVHEG+hDhCQeHDwU9MDpGwUFj42KrNvg2l6Jpt3Oky9f0KNU2m36ofsdmgNPa
qooSAkxL8I/kz15R+G+BOfdqteRJ+7mmTmYjErrKqnEjBIorQHIoW4j2EThdOAKm
dQjlrSQdBTc+eEZIoM4CiIaYy3Q9rByICiXHmM+XNmB7FMsiHP/hor8qQ4Q8KP3W
+OPBxR9Gr6H7hXF53B8yrzWR4Oiz9/yVhhcZQtqnYv8jgYHuMP0DrEs9/QyBnVAg
QS/Ocqeuk9UnbLx/5z+xMOt80rD59GjEz5Lsru9OVJ/acLBq1jm6NVVWYJnQX38Z
WjnBG4fghfZxh7JiOXD3R1X0rr9KjW/jlChEbxNylq43UQmCNQgEESiVbrVMqAYh
y7iIzSlYrf2o7NxM2kNsSIJZ838E2mA5UcWrJsNbkCYABag9aq3erkL18ENlBO12
CN7X9JOqC+Ra7flS1RTZQBgBHQh4SxNOVljpktaNTrw6o63URKHFBZ6405pmK+TR
KhXBiaGwBwT/n0lRA8HiHEABmY8mohIHk2U1H1olt1yCNFCsbTU2ODmJW3eC8Hef
6kvchCjCuqnPCywFbmbJxsYiZjieeTpun3fPunPQLFBGGjh6IYac8rJTOsnd+H3m
v7VPx0eVfKkLMEELVNJNqraWtjlt686NCJLp3xIj05svu8hcLgbms4CdmjRB7wrI
GLKiwXt0t0bFgTTsERMDKTJI7FrZB8qMsoTWHj1MSNYhaZc0TFwCE/JAfIEu6qzm
d3yXLOuVCRfBDWjfPr+BPftgcqxU72BM8y2yBQW3E3I1PRXunfPdXwS8siHOw+JX
6PBes251D02s1MM3Yi3RH0zV7w5FC8PVzWWdy6ySGGzpccPxLr8f7q49tYKRY375
6+2Dd2bwCQW7CNOZN8wHQxB5oSiRhs4SXfkpPkTtu40j+WJUQrIqQP3di8OAe+FY
QJpAjXmByEjOJOFpBELVT0H/ycczRZKWbISw/cPnE4ibOvaUKc04IR51U+iJJ3zO
NiS2v1WEh6s9R3MNGpvnP5unXYAxJFTvTx6QmTZM75/kS9Lj9+AwXIarMmHwt2Qz
jh+anW2ymV0uUt2AOPMUPQaEZedks/PZEeL2vesfRP2Nkkj9P6tclHPp4aXz8QG+
SGHK5y8dGqycXQu/Qf2p8a4Qu6snTwn5yKBMGSVz5oMUGg6TDHaA5l6ijChUe3tH
HmhGUyJ7eRTR3lXalx0kAh3DxE+QHtXXcGSrLv0QhOti2OO6MoVSk2NJLPaJWCUf
K9KkAQnwe8GQCTz6ogUuCX4eFEpLqywnIxDdQb70oRntG3tEsXpNbUr6CgTxyFyE
0tqVQ57DNTE8uJBKsK5UNF9AGBYTBvS8Sm1AJXahYeEM7jiFUPUuIb/OvyZUgbbk
2B+rFfP0yduX3fBbvFI7sa6G5a9H70Htzkm7JgB64E5ujU+qxCSTOSe1rnBZf8O9
Xv+VTM/qgbddkQuz3TYCrLs3mXWeLeVJ7N8NFRIAOHO07RkE2mAiZIdyZc12y+b9
D0suGjtPNz+tPJCWHcxD2QyLCU8EC+fDJE7x/nZstBF+dBN0/q4tfzz300EeDini
VpOhn1beqYOUl/jkH0xfZEyTS/goDE/svFCctaXXUgVy1r4fVAYaMn7OcRbVllNo
2YpX0J3NE15F58oT8r9ri7gFhbnsBCODn1J4cdWC6V2uNVT6On9LFdbpzDvWZw9W
BNU3sJ/RtmW80ZpEPdJquOYW8VRUAlZDMh1j3uxh7HkICa+AZiTBtTrlmtPQmHxX
P1SUmHDLWamELFWYUtPsVVLdcmAuwT1ABNHS1+UU2MfBXfkxlhG9ygGM+tH1iH/U
QANCWCu6blmtnLpwSXTtFpStcrqGa0+h7yRQ4GSwchjGSXVpltMlI8VIjobWmBQp
w3MaU5sU8XDCD+YHuyfACCRcDg9umf3D+X0n+ykOL57VQIGFc2vfHEWBPLFWQElD
wRa5zNcndnMKu1JFXvoCi6B7mrvINL5/cnKhnMXMb80bgYDJFd178ElYDXw/kUuM
cw8vQIKoXAxG7FDSoajro69lkNBVE9HRL2EppnUSZjOP6MUJcxnS8jcsefQwwbJ+
G7F6SGZvDz2rgsJE9g1x7V0TX4NHaTXdFeC+4U+SEgc6o9Bf+97EceyCk7lJnWal
Szd35nyhN7cTaDCCTR6Lk/RcqB7MKCiJFhRZ3GF36Ip3HR7A/6hayNBRjxuHhc0k
o97Kd9Tg3U5HcwiChZk5Z73ruKkti6pCc18QUYls6ws5H6PQtRW6/Z01M5Uqh71+
IEQVjTU5iIg3IN72mRYK1KA6G83L3VDzUlxuaMVGAnjUyVa/kAQGgk+NUieTYYOF
BithfC4UT8pUqH1rliwuAh53VTm3aMHj41nqKNAjf44Wl8hllgAorWV4q4+0Oy9/
kFIEmyDDLWzoqg5KYd5mO+WC9+bOEpJkSJ3hfogHYfU7ge63DbKtm2SkBUBWzoEb
eZZaOQpYtgSEoj2N19W4Wxna9q7ipsLVN7PXG35lc0I0gNEPq2OvsqMEhERlpsK/
C7Bt5gdMUywiC6GtRA/kw8FDymDjPwmGq4oTWka2itYsqzXdrQwVXyPY1vkzIicq
JkczW2HqgMtMmLmxthQcVxU3EmTRHGsTp1vknstcYtLYBbdn/IemKUADHiuc8Vx3
C0pBbjuHCaEAiLJjbBAxU+uwSNy+ilcz7HOMwFU0/dqlm+yBByGDxqdzV9bgXIXR
rDDyJpaGSgKnVMya+5grOxroJT6yM94uaYj9jk8tBMVmEest/kqqjYdpSO1Vgqp9
4aJAghfYZbEuueUYrLJbc6ee5fEyZxm+mfIRWmtELCEDw7VgnZu/+t/gC5RNi5PS
rZdzWJeNbPQQPwsQJAhtfCuOyYwe7lEf3niNKOF3YLff3EsC7nGzur/wwKxL++R+
Bpxh5WNzXeBzmwGgxjxWPQV1hZozp7aIO4M9vqvYdax+NW+PWi/sZTDf2/kS2PcN
Sbt03qCx3n9mXAvEQaI681ko/AwnVF85vFjVkh7PHkbVBwT3CN5JVUiIAzx9gUip
rx0bs/Z1tW9N2rWMUSFevA/3TkIkRovVya4aGd/mTCBAQscpG9Xzhl9ql5xgk5oL
OLLULkvXZGr9EIjd0uzQB8wOtMMngrqdD0OcyZN+WdJQZApEMgge8wS+c6U7t5tK
wP9A/4vAt6GzSKUkSbhxvu1beCWMq6KwC56oERR/zkqXzQ16k0FHYszLtmpRGiWj
tCZYedBk6fvn9mQnzyozl3OHJpfzgxbdQtX0I65uOSm9q9yRgTZANeobdrsvp3gT
FbyTWbMcY+c5B02HQ20aTDI83x4MsBbszMWCr2/U+KvcEiEaWcsZHh4wJ9UkLLio
to0ndaoKcL8/dgGgXalQGkpqmnuJ9HJg+9AtACUvcezZD3jt2jqpCcMsCFzWGidh
AtLyM/lVZ8FqTurk6+7ZmL3VIvt/S5aMINXnZp7easy7KQco8PaUNlgSg9NWO2iE
JccaWX/67MJlupopVc4P0dIzgWHgtTwfeY58KxOZgK01L+0yOx4QadKrUBjhDN8t
ZWJ4uNZjKCEVWRKNa48IH9e4PybDqnf1kr/Sd0b4LA+zOwlj4lS/danC0MWiJ7u1
OS94kJF9whkoQCgebRbxzZX+nDjLJrRawW7Y8HuZYwZzNY0A28J+CDHCj0ZosZx3
bkcJmh4t2Uw0L+BpvnjcLNx1UagTkboTud6DEiEkQMTIBdZbTVrCedjmrVjcme+o
LoQdSo7ngKb2rurCiaFwstpIev89mSz6vmZZW6eoGVhCoUkRh8jg6LUXkK9jFZvM
M3utjVu2UWj6IyY7zrmxkQhErSSUGSXO6/J1AvUCO/XoWpcI9cAyZ8wyr3UALck5
54Fy9CmBP1cwQ4BgERmDIp6cZswAbvE0g3mKmy5muVc699NU/dGJ7IZXHSKcJrP7
PRvfDaGao+ZO4DmDhQRW1hfUKf+AsQP1Mv1epjrGPr5VW1lh7UAcoxiBgWLMFEJg
uWvZo0aqRf3Z7ZNJg7tHQAqXHEOsUmejjIM2iwrLDOI6rYSSlhOJ2QXjmgRTYJE2
zNgtdMcm5V4PGMqyP5vWxO+1Lr1pdHarSzR3WERQWSibZevx2ePDp5pM5ZRtj9kZ
LIevgF3WCHz/3UJJRc+tjhPI/Oubn26X0KG8HNnqL4CCVaGmgHF7O7/jYpEE4SlZ
x8LrJg6g94gKUvLIwZqviS6hlf4RZMRw3GlbIq4Jh73nnAUyIph+8j5zLl0E7+Px
k3HZEalFg4YcFEnYav94H5iMOcekv8nS9qacV+u6eeFyEtwIJrC6OcQdGzcgPqxO
BOZBjwxoi693fQSVyHxvZhnl7rYNPzJl9mR5JAEXqW9p6HuR8CP0BZ60pEdIxJko
2iLKoOjD/RTyLvjREkikGH1LbH704d7T0+Px/blkidjmAjGP9f5LcWuidj688jnM
JGJExNKI+B5RX0aWKlSy/fTM+nmjCab1v1GWgQemuy9lpOmrpO1oSUV3o1/yrIwl
EU4PiPnaNCrxUT3XDkyp/pOBTgG0xSyRDVI6XP+GZXOyNqME3wv4VpykuHev58/Z
3EFIXTLgYGNkaOdmkFECb82cfywHrJygQoif1rCwquygSYJPNg1S1yILFhSKKbjT
Lh9pXq/ezVz05hb6f3kDu1UoYt0zr0m3DjhnHRRL8jjUxEUdKvFe5D504EVxHDm9
YfBd+x2nH6foMaIK9NqUskARzESi+OG9EgYueCi7lqmziVda4wqnB4ZlcAhotmHa
wZllxK/0wuL3htImfjuQxAyLjVvYbQ1vIiEmWT2FDy9UYOWGH2L2qj4Yy/2i4ILW
wy84PWza7rF007lwAOmDXrpuEppAR7K1J9G2z3tjUptLYfJe63T5+QmZBuxNzlS/
r2WUDF2SQEtVJePAFYuKJPCX30Mx2MrjmYi9H8wy7gKqNvOcMGuO/A1S/OlnSy71
HgUZ42JrpAiQBS9qNHVsTDASKB0VlYbGX85Hc6zJooX/WzHlcpD4X370DYQoZzgK
6eToxXxWPPbh0kCM1PcYw8fUWxDRGDvjkQC06LVOLXFUFwSL8/tNqKAETCs7PPYI
FYasKQfj6zJrzANPDPDgbfvk+eJW4ChGajDF4So5NK3j3lB/wRTb0sJLKauxSqEO
40+V+4aOYPuPr/DZ3/2NE3Dfj/QhPHaqE5LUy1S/oj9MurXOMutFGBdTlMAFE8Z/
TDB31BjomT36jhHsfjmQf09wcIBGGdh6JMElUkT1l7EWdXE+3frIudfYN2dhN9xt
KWx/qn5MX3e538IoPCi6ki0p/DMbxrBDDNGoX6Db9nWYlhEBzUR3EVahsrB5+n6k
E6QmNoTp0wvkg6RL8Ti+biaDRkQbIkJVLv9KCG/w4ugJ1tpm3e1ay5nXuE7LKKrZ
pb/ESiTV4kvUou3ygua/kmk+jD+wbxt0dAy5S57itsuJTlHDNLleOCcPqEU3/HO8
EKRg9nVP05Niz47knTo7MTaLESa5wWQyxWezfGNDSw548rBOApDmqj3NsK7Aehu2
RXK3mjdJoA8VAWzxZk/mNAhkHP1+aggP0pOfkjHUWeZ5EWCnEnyiW/2bdb3wnQSh
NXqx6Eflym0+reoAzjnMN02tJo5Y03kBzZGdyd+2a5/EVfikH5DseIbLozEQxzQj
FULZYLsiG0v0MMzsUR7xwahvWNfmoXVHd4biJSbk63dTNHLwvQak7/VtOdiR4npL
Kya7pI3WX9jtg0rTuMFcTJJUsb3GAbtYcrVy4aOy3a1eHMm3ZFooipIbl2b9m+V4
ZqTtXRZKnxhHM6jqhVgLbaf2BlCbN1df5FCu9MW7PxbJmBj5MG0Lfsehtmrovi2/
3bTAQYgbuF15nle0abpUUjH84iwTzVF+NhkUc+DOjt1lJitG1UXb27+wRFd1S9Mb
tijI9Rag9Twdk/oP2iVLNPfInjAAuFsUdUL9pUP5SXO6yEP5fazCkejrHt/liXav
hXp+c/DF9zcl3iHNHWcppi4HQosuhH5ytU8d11RsK2feu37h9TY8OLOn+wejwp8D
IzmOKPv+P9fphLX60Rv8WkhWYwYe1iHhdFvdQz5vQ5192VS728uh3bzLkUSLjtgu
HBVLrJUwfyKhorjMUFaAp0vgk7HQ3Rckob0QpNw5B68wpKin+nrGFAGNe9GzpkZk
hOJAYJOeHaSOithDAdBY9gZFgJ2kR6RKTpC0qZAxM1IJxb/cmIGK+S9NBvgiK8aj
xK7kxxHK5s6KyZ2NkOZyytK1YHIOlBcZwgBDhja3TquyWd18CvtaW0uVYRuSjjy9
McOO2DmpOzQt9lrERST8NbW3eUaxubWRlrzRj1N9eD4FZ2lQq9kuFB9noI9g36la
LcmmAaaQIVQMitNJ93EEGFT4Cawsmd18wK6tt/va54RNe/aza4owlIEyzeEdcC3i
Jll2nigcA287Gyto/FJrjGFzuzlZuO069/HEtQYTKh69Oh+4CNC7x7HPeB+DG3qg
e8uqOuzij9/3jv9VJsdoBPwKaaHs/WasD1h3WeFljn4xNDVSKXWWup8ufntSm+Ew
GYUTadKjV0ANZfyUqYJcmLlOWgrqSkHND9hgWInvjP8qIxBQE3n8p4yNA82dxq08
kfxQfjatUw0mwRnX+NNXVnn+eEp36vUjsLjjvYstaqCLJtlAFRWGSeBI7Oc0iSFj
6JSyIjrKyfXbvR+H/dcXSjHT0ouMTF/Tdx1L1Nvi+dw5gHFrl9mCmCn89bbOqGZZ
rhxapmpBr8k3WInXacQIaFNp1U/Gz7BAXP++dIw+HbSgCmVydB47qu19zJymDJjL
1LsxVGtSEsLtp5b5kfWjwLtn/75HBrmu/rjwJ9sy9FyFjI0Kj1SrPR8p4bC9O6Z6
3ze6G81C9UjxK1KY35ntYo6OYW+SLEnjGN8d3xV3qBgtglHL4RnCEoyTqRF31rOc
wyemKWhezMf/IBt+zwyePk0V97N45QsgX6AmoIhkj43hiI1tfysfXwMy/XaA5xup
gwAV+mxKlwFobtS62O7NFvDdMkfCHhfmRgnhuYjQK7ljTbYrHh6Rti9DOUW16GSb
ZOcgoeXx4XDxepfBoJwHeMKN0K8rAiWevvRkxQ9mzf5xShUZLVQavQCW5abB9tUg
PdBbzau3NQemA56tn+AcVEjGdrM6IbfRyNPLbNUldv+/zSjR7lrGB9wJsjrnFWCi
Ab0NZsLygKD8Z+MREV/xAYNAT5QGDZJYeUVjdXbRPnCGAahvlpZPBXWtfDIhimsw
XQGj7i9gYP9YtijpD0zTUY0b6zG7zg1TqbuhztnzsEN7BuIua09fYIz8jxDib9xd
L/7eJ1oI6kMIOiA4C0snsEb1AYNkh9vXx3QWChRImeyXx/n1WMG/Jygdl4Ln7rOT
S1NbQXyd7NF3dXeG6xoaWLnwjuaFcYqr26g1px4cxyQCTLF8laTB/vLfqf1ID5rr
TcIdO9hUejuHIcHrjSGQsQf/+y9F89wIhfS9Wb9t1tfLt5XNw6LJh9GpjtFGIBpr
CxBhrqNSiSuAG/JU+vnvhuyMuXs8FyvYbBEenDWrC7VPW9H8UM49vRimF0omgl7Q
aPt9zQrpSyV7yjnbxQJbmB0z9s7mYO7vW+7sSxLowhZT9+Ix2pm1gCFJX8AeVZi+
c121KWRpqdGxHNjnRE2svOUkc7NXF1nxqO8HkiMAYNq7frODGC8gEiDQ62oW19AH
AVRdnvBcBocL0Px16OZHBqhHcoLsNFp7ok77Psj0D2K6HBzT+nHMB49ZeTgCnUVJ
v2T0xZE2Lg3JO9wodX1ty+0VX4nif8dJrfPPFTzMqYla6I2zbbeqONZbtOQhjne1
O20sL7DTOGJkLXc6ArOh8Wbul/ptbWCVFfs9ceFDw+1ubCleRMUVAW5ju2iwyP9w
Y+bl5bT/jFEBEqxrNW2iCqHmqnbgjogqmbZVjUcQ17EXyqomRSLlsZa6JON5DNri
v28F++7MPESJeP/T5z0z9QdcdR/XkUa7BVP1+r8rtX01XSAK66r2B7Ap1l4jA5aY
Bg13+u14XhxNVK3BZvTmPU4RgKJrMMQ8B7NKGINsX+cjamP/5iAn3ILiceE8zlZ5
/UkxenuCq2+a7kXXirgZj4vPhiKj5W0EmaESpv6sGni4ONP2bvgH9lztbSfWBJL+
AeByyCoWtxxVVDH0XFuWfBOaB0umhfX4fkBOC8/Wi5XK4PCzpccOibX/W3RZBNEF
NG1/r2nsg+Og+HBGQJ0ZAZRSidL3d1+2QY+wg7OCgEs6iMW97/L3zwh2CP+0FtNM
WUFCbkkGCY+PE2NG/pnwYQTe81+qHilPWPet6quYBKbtl9C/2sZB+FYlh/AvgdTm
LoluhOmFog8KCo6sf3KM4b9/rfx9p1q4n0ubaBbsl1Tstbm07Rs01Flmk9+N8K7f
jliRDg++KS6ETY+rsHOs23ud3vyErP1Q/wubRwCNABctIkqtZo9cMGv51R/WY76u
lRnFilUU3kSmpuG+lS9afs9mIhbjDu9nKad2Ckuv1/nGjMKNlvm8shyBMwNytdMN
LuZuwdlWwFr8mtVzeTeM8GOeFKUfXd5xvkO3XZDgNOUYFvQlE4MXGOt4s1zN7XPi
9CWfi8A9yVh1QlzYd0twA+P3wsGmkLWtw5QLxm5+C3fKJVL2mJMLPR/qy7XeAoJw
yS6vRiwcg7BoJ9KEWykpv9XaJ3HNnbAphedX818oIu4TOsVGImalPfntN1ROSbLs
7ON0Rkd8N/w5sD/M5VEf8eitC0iHsmb28IXpVN0nD1pgr8D0U7X2GcQQ50uHQT4O
OXI3hqwpNwDK8V4Eg3LO4sWj/hd1MJjsEP+mfGsTe0QYY9sCvkT0HLeq9JEtl4bD
LhdzaZMyKpJOpaRnYLly9m0ySK6q3GoL2wihXs6FPS1GdKGOhFQdMN1AvhMP9HGl
joLSuXAuRWetMpAz3IrkkE24Hf0kluoDRuAK1DU/TMQvknALV6/Bix6SXxfVI0yP
nVt6PIqKiJSJO6cZinmEnRkTMrCplRRkJTqNfvAyGPMsic/l0BNdMtaxWJxg5EI0
4x3/JlepqoFVL4qF3/7PLU8rnuM6zvE4mBLYyYK7QKm/9e1mvl1NodCi3i7NySp6
9YOMU+ZGRz9CIk0+3DzkGb0P2xW0bhmNo3HeHGL6uYW9a31/DoAoscDLIV/OVTZ4
xQQzHZrmfRnJvT0T2W69p8DbXkFEMZCxua7KwuGpQvh2154finqj8QQaDUvI4yvD
1pWhaT2kEpfKrhVIlND+UiZfDokELi8XNn8zL/ZApM70+yHJouCGT20TkUhTL3mP
iWulTBk1gChHvh4hFaOuLXzSf9NVAlGvjS68lSDcAvqkd67INM9HJkNef2mUuBf5
rz5BX++xm/ohbjcbmXK7KbdCd+WMPqF12FCrxjEi+ZLsfyhOxrn0mKbWTDUNEtUk
MsAk4HYhzEdUB4ApsduVi0Vq1AKBavfYKI9S/Yk1liU3fiauT6JiTyQZIb0u8e15
ruzsJXG/CLwuS9b9WU6fB2f0c41/DrE6JWQvPAiSV5FSdMvodz27402cNRdIlRxG
2rTKq2k/aBsDraB/UiDPHxXDD6Ov1wB6Wsh1uUL6fRswqRwzXBKvh3VUX4JvF0zv
Pm2xIa/FGxQppau13+soP9o+8I5vDpYzv4fOxMQz6g/INCyYSLMksqEJ7tuCSuF1
k0zfw+WfC1NaHGk+qtG5PwJbLZDONSzND6cCzSeF6sDxUotBNQkVw8U8XYt5BngF
F0HbivyHXKucNpxTonLoZkDA842s7joDs6glld93bK8qHEfBC4gtTN34a2Lyl/UD
ueauQMOscRkjlMv/ca4/mnlcFwyFHRagKNxKsSNShUdBzvkoAcXvojTyBJGVD7iH
F9qjKI2PD9r7PyisoCzM4ZeQpkSIPlan98QH9IQFy50y7j54NHXD+MvJQE08umZR
3Hfm7T5TupxmoD+2+GE5f4qFMKkFHzUhpD/jzMELUbTDnwgCNZYoxvjObHPuCBFh
38vse5fSXfNrmHe2aLS/e/LA8b1gFptfC4duAiKNK1kG+mS5XU+LdzDxvYiuR9t1
+5P9spmbuEgAD3bMYOfG5ZD87zVx9QK4PbVo7v+/RdlxRqE6skdCEIpWZuhYxwHF
0rD7Wy931tHxmUuTtMALW/gIvfTKgXUPIMgH5NA9wo6kV6fheixl7zhQNZ5rYVnF
NZUJV1LXzNXGi1oPTCv8PgEhGaBRwVQBEhNE8hTejvVQm6YU+z7Nl6Ly7iOXif4R
ot3jE1XYury4JnnmcybT0bpeWC6V8VxGQp19KLoxURE1+mQT2x58rOmC7QQJovIP
pBIrwUm2dHEwswZ26/tbWI7tg6uBDU403NU3N5vsJYdM2zm3OTOHnXtaNxOl3zCF
mvh+UGmlf+lQsJzqSct4uPaX/14Vyy3kGItYhqwGfhhmiA/fhi8T18O040KJpexO
Ra2DzdrGmbixTg6061YbWfSV/TmCBJtIlB3PsYp9zWhzoada7TNhvuce1LkTSdhD
qgLaSw0sMKjEB4NNscjVq1W5uh7TJSlXe1lQHBWHhlXdNn/Eu3ut42uX6THgdgv+
nlRsrrSRG4h06a+fJP6YW4bxu6tKsSq0JYI//6+fHgXWjQrpqIqDcEjSmpAQp340
qq169mi6SVMU/MYwMREl4r0lNqvn/14LnaD/GCWSz1EzCv0X7s4NUawF8+7rvv6U
f04bTkW0XNb5fFiio8eLd4/NTCbz6qIGF7k/t1Gu1z6E2r+10q8dhfbDO6f9/G9p
C40rN3zvTBoRTmxiZXw2oSMmzm/2Gblb6NR4rKtSRUIIh6CIzIQrvKjQ1vVz0cZq
GYHGMTGLLx2u1pbr53hJwx2DiiJVfwHeVQK1g10ybFSnnBzJXTGaVfD4F2s5yx50
+Jba/4iKXMRKVahqVpgB3nVIObqUQ3yiINg1OS1bVJggQskFUDiwVa96A6apR8I6
llNVLlL/TPxnvnMPbwRIbeI/fUIcx6yxT8o62nSi5CUel7KLnsg2CCNhGhoxl8Jr
5mKODFjA5NSKcKCX7a+EQqvAEgPsjnOg8+cFYaf1SuF2y+5BZUN6ROClxz11GBlT
VySyq5dBwD9NqqwkII0aNUDGyPJZBJac/BoJmeVDC6lIXeQYcjfAorRjDwNVLFVk
ofsuZhGkuFB8sN2VhmmVjmG7qC+KfJGDc4oV9cOLbTzOkqRKW39Uds76IEEvx4aE
xh9ZGcDcmUKStZm5+iLhUoCE9hjaaRLqMRqa/zaPedQKc8m5spnixRIvh/IMwWQT
XmVm1dCEbpAqqRT24c7T5HEDCmZfYlMfOyi70qvLCkbqGjpXf2FKflgTLqUnFGiE
A1jfY7TahbE09noBz6v+umyIGDUkKaAKC5QNFEZ7YTDEEozQGFNuWoYG7r29Urh2
/Q2H9O21wW+UqnUmbUDsEKHW4kLqB0cCUzMGPD5rJ9tXK0L1cWFdUdqAuAghquIB
sGKub1c8CeduwIcI2lLzjur24lKToEd5VD23jsB1IX6rO1VzRANcDCl+2BxP/Lwb
A0LbZoJRjWMNIIPG9YL8n+PfsMAhvcaSpwzoOgJuaZSzt2adgyuf/wWxRimmJPBq
CIfZ1MPpPvk+5YkGxI628BFjXw0KriLtboUXKXRntMdlCBQVedHXrmQT3xr3x9BD
SR3I0VAmij/dqdRSp7GyeFrmUl39H6Gv+pR/nJeJ+qNB7gnj0XEg8iaAdYlfRRKv
s9Li4rRueAuRnMABpiz8RxRgxtIBTxEL/JukoBNJhVGtxjdmF36GaZQ6Vc1YjQca
9rZL9Sgg+ag6z9pXNIrcq2DVixvh0mz9nYaIOBV46fkyos+Zs426hVqyb0kLW2bN
uqmPthU6ikgr3CH3CPMO1YBMQJjp3/OAwuUkwEVOkI6cGBH7gi3lyjhwFHIczY7y
5ZsfYCO+iw5wf+SkhxJwTIzXHmnEadQymr8nH29ogS/jRDR4qYNI+o/61c09bEbw
PFBhHL8lVJDMDzbZ9k2P5TIeBv9ZPYbC96QsAVj4zVSDQLECrwlhSRK7TBEjWuUv
DaqWD/CVIt9BmyaOBex33Xl+5egt4X3hVBs30ZkWALalbyyGRbfBdZauTDg97m8K
M/f+SWoucBYatl3+lfXT4p8r1hz5GtSfYY3CYRa6vm57iC/NXHGrUcaQ6tYVSiri
K7B8F/WQ5fVHGQs9mzmLvm3H7wxwlhe+8A4OtX6PPlK6Qnypq9XocTu1NFsbRMJp
Qfz7M/cjErasqcGxLP+45D0YbQH0nLgi3P+WfiT3yf28/dwh/MeGKBzFAWgBMYeR
7SJ3Sp0aVWHIufSzZZ967GRZoMXawfJ4VGDe1DXC5soh9kEkdva6oDYOw0pKcCZv
Xm/E4Wee9SK62KjxqVQUmh7enPpr2U9ZWpe6dtlYZgJBCSNomPShK4uj1/BIC2ee
vahGnZgSC098O5GfrmWkq4ywYM9Y7UeHu/37DmiViHeraVRre3F1NlhYYO3mCdXg
h+EMjXqQnQB8vtn7FXdHJBNjr3rgdFVUpAdkqrj716K3hp2RsN//nw5PwQJl+1bV
hY0RfKkeUvXkooLpeR5e7gY5geVRMcySKkqlkGt+8mCwQ5ryfHV20/Sjp5wK04Xp
Eu83+opORMSCf+uja4gblvkS9jNzDGin/xH/94T6I8kAcoQRLQMjBBehTpFn9KVj
Dlrnpj/+qvVotNMk+WSdHNDFD0wnmBRWDJ2EIoyS+x7SX6q59pkr/qdjT1VhWlj/
3iJljpozcTOErqMagI42+C0g99RsKocW9VJGPJ3Z2BxLZnDqFO5n5U/BhN/A8KYP
hoHZ/nNO5p0Pzy2z7PekTcT/hraL1Uh8ND/FqUYJTmW/WMumN2cPInIA+flPgLgs
xxyBhLTb+TiRxQt46pB5l+piv6Hfxv/BrfILtkVYQoPe4EqQVJMYlpmwvTPd9gDQ
AGUmu+Dv8CResBaVS7lrN5aZzC1XP5hEAsklks2qNH24lBhbUxnMFicxTJrxYVUm
r6rEpR16WjD0RAlDlgOxSo/Hr7rmJElfCgZeuln7QCahEQkG5JLZ9KTaFnivcShU
IghEMV9563M/AbZ2KK4ZKd/8m+8KZ3yIqyhiStj0gRLDONc6s6dzL0PVcnajGFB3
RclOKTmSh5OA5CF2lUBzjIZxdHySDK7HTQhrmbE+L/GLo1z+qVh0h/2/7B9QxBiu
uTGzmX56xWO0+ljdiKH2hSrRxa9atcU8L7U7p25BKg2FzZ6BMxFPZnp9r+flqHzb
rN94WaY7Gg+WDH2aYPQ4vA1vY205Tz/AF8jGjnRL5fdx6s+rOclE87FdOB0g7WqJ
NIUxarpeHd4DiiYWrDjyUeSKkl1VJd1511zm4eIj2m5X7inaHguRNLwuAkW2Hybh
Pt3qwP5ZkqB73w1rOAD5zOrTr/ZGExhYgnFNxDgTkG14vxqM7hvoniLYBNS+Epbf
k6M7oqC2/MOYMKbveoHmao1DIrRK6gQFxVnJ/UO5V+Ls+TBtcqbHFSEh2nwyHTja
dNmjKWOeX6NlKNFzGcRB+f5ins98k9ySWyW797SPvwf1sVCkNk/NCAhWP8eG1GU5
g917ZHqTX2S5Lk4irEBvqN2nzj54HNY0M2GdNp845tu/bn4hJ2N8QegpSricITBV
txaFejui6OKgXCHxVBrWH4BoILBgbgISgjDx8RePy8Nj5HzsAgdpjrueYkHXv66p
3ZWlBBUeG+8m3L/FHPr12TmopfvFyBTdigI30TuP8Pf5yzolLIO8A9LpTDZKPmvi
T9zpWQFUGY5M5D32YIZK9LUoiSmhPl0/DUypg/gkvW4hDivLSWr8afw/v1b82J76
PfJQAlt86yjAWRyVN6xnzderIdRJuVDThbqJgIEc94IvwAxBaxkySp1lwK0jM/ii
VeJ3V8BMsUaOIdunpDMrLiWa1uUjhGWLEozQq8+xYKaGA8qtn6fF1QAYC6dRlZq9
rn8UVVbzHB3bvZRm4B3xHzFCNbMsomBjW68Y7aztcoidtKZZ8nA7ihBWRlKG9ONt
ngY8g/Ryxn+Tbd240uoSYsLPJIKELbDNFObvfYmBlOI3OP9gaAaT5g1jBnB9+b0q
Ajmzsg5aYEIGu2GH/o7USx0E7pmuM3brWZiN/8+jMozGDTKQ4KonALrfipDFomIZ
aGPbqEsx2If2GD1as+XykG3UCghAcCTZ7sMYu/khtanN08dPBFcK4aApG5LAXEYo
8p2ZeEiKQzqImqQCemN2s3rBdIOVvzcqMH4QH6NlCpPn43eye1VCeNG5Cpo5L1Dw
XZbQ+wf1HBjIU/x/6uFSNYFrbzzuYelSgQ9qd+nqihp6SIbQppTbnrD5idkZ5ivR
STjpaL8u9VCBFNwJuUD1FeJhta2TChRzBAyEbAWkQ87OCXYDqgszz5pqZj1E+7Pl
4f0ynSiXwUJnBcAPP2Jwj652EveAQEd3SCHoZujzJST+ei1RXK7xyHz5QNDd4TQQ
E7+6CNHHV/G/AwYbKsRKebLgIdeC47SqqYqJ9hjMXOyHt6jN1QDly1UoI1K7Ff+n
f1Z/2y/I2K1L/gA0yGHwd74HvfMHNVVW0ISIImO3emjYtJadotN8q6hEow1WixTF
v/RlQ3fUKmK4H7AUvmBaqXWvHlUNbvDGl+cb3bhjsnNyXxB6CWtPf6amQCx86Ug+
m+obRDm33/muITG4lxI/6uci4nnFfEFBGlzVsFYiH1OGiUAjVNoDJqi2jGoDhkaf
HhJG4svnaVfqIm63BL0KItk9jGP1mNHAEYwL/FObckKkcCOJi197TNC/r3nf6qBQ
zEl1ikFffLP/rphlmYPCCMY6yAAcFmg+nqXTs4Gt7sWLJ3KpeOcC72+pwsvGsiJt
reNHTxI6LoeYbohGC33hNjZGVZ4J1iYQHGhlOyQ0mD5CcAIbDgGEClA3uEV3iSYy
H+3TCVA+PUYRDMXEN1aeNa00DnN3EHbyEAMRsdAUVTlw/bcYaAelNcmeEX06Tqxn
OMWnZMuPrTmRHqDX12bPZGtpAp1IBC8dGbQyKwZGpDhizDi1q4M9kSUJjE0U4a2H
bwTR0CSoVEtrTT+XN2qMEOzdYjs47oD9ebxdOx/Yirl8+jsavjGAccdFd9BMoj0H
YS9gckJj1/L5E0YS3Rf4fEtIRAAqHeIlDflkdd6+WvdLtAGgdmE5nAv7SXjIjLQn
+RuFTgzDV22cLKoLD1v96F1NlIumEyX+mXIyWYuamdoEU5cZhFYsl0q6hdBbYYd+
g0RG48jInJZtfvpIC03EUEeF48Pzkig9TFkO1F9NFX4UJBFffxpwqd1zMmSF2bQe
dti1OL4Ebfa/T5pJXKoZJBpezR48y6G46p0m7tYhGhkTk/FnGW7OpBtRfLpZObva
98T30pktid7L0amXu7Ax3wyz5AbGMdzOABq2z3HlJRtyNXiC9NMSYgDdkeV4rR1L
uEIyBg9vnAhfxrHcVYf6y1MApBFcchYhal8BqGt5nfq/dJ71C01x+D/PknlZ5on1
wmMJgIZgGoCo7te2MGytK7iGiKyAkPwIxAVU9s32jMZeXCOTSOK5peV52kd6jk6/
EpOI4KnnoXj57EUVX66TX0XnGO5TLc5MdvMtY6fPMVKmN03i8Klkh7PMQZgE2pLl
g+baRZg+hiWYsRCmfsAi4AxD2IukWoh+L/u1sdRziTM9TVb2Xpyq7OOd5T1H0Fn/
cnK3M40+xV3HvrRnVcRin3ptMZDQWwy4foE4i5DIYD+mIfaSWTkrS3t0dGV0W/gd
1xuuv+09x4Wye3qpeJV8oiBcNsGlGaD7BCdTdkEoV1pd1SDAwd/D0IrUNdpVUVTc
RZ72sVMrBlkJ2sf7G2rxXHMOKgbOVBWtOQnjwPY45HGhmXo1MA5C4GdSWquof2rB
hYpnWgEplYXFUhBIRSaMwhKTr49LqT6d5QA+eYLn95EjhvSjUKz+gHVb3RJSKw83
Oga8GHmZ0YellC5RsqD5rga35knWaOqdpga2cmyYk2oXlTLC0VIQMTaBK/1clViR
VuzIIFlNOy6kLPIMgEO5qxoqJroTln1Q0SEyGLgNEzzLTKwwDf9BL8RQym+Rlpmu
v3i208rhPhDe9EOLiC+q118lMFfhLr5R27bKi8kfPMOXDmCyemkZYPP5ti9YZFls
EYkr4dQi2fLx/PLtoVPx987/EKlu0RgkAgTcaZESufVAy0V8YDBypm+6E9e7MYvr
pK5m2ejwetOjuET/dGWKx0sNgaoRI7Pxun0D3PUU27XaPkrL21ve8/S6AIU7Q984
3+HiB+u7zXVRnR+yZoc8pgLKIxX3FoDsey6xOUmIQCirKbHY8pRA0+iQDicWFoNm
5GNXwEVM7Ji9N7CMhbMf6OaGn2qebRxPE5MuWfIFuIcUCjdm/Jw91J0pKOZzh/1P
XgJAMltuOD3x20I013Y8SRHA/JVKPcsgf2n2HlmwRMf4+SVHMR8gilq4uJFUXt9/
mhlE3ZyIDo0zVQTQ6WaEvIMNGVbcIMu77iChH7jtC0aMPZ+mzBfHebhYPS4suT8M
lQAVi5eZaSYGwEfxwYTIQ19KFFNC+YMKzu0dvmQ23aMTSjbuX8Cr0R9X69oIZCaC
Y4E1H+w+3/KBl8yAT+ap+n1AfXIdm57gX2W6PJR4No4q+DS5LIip0a5B3V0enLHv
peuhoCdkIfpu9K5GdJNiRILUIVTSCGD2+43zMu7mjR8BzQA4zBG4joLPWILQxbsL
OFLDQRMXMevaYck+3+VBeBBFFtYwSvuXMRMyb4AzNU7sfVGmQcnWR/qDVoxpn9Zy
G5bFBxkj49IsJ6llapt0y3Dqu6E6f17/Z37eOAXerg0Tf+kVeDNx7+aHhQgoix1m
IT0cnPCY40Nif2lVaIj7LQCjs3YEbl6aT4T9QaZqiFOVtT8/NwQ2YWIoTA4QoPIN
lRDhLe75Vt/RjYHi8b1dkDS/oUVD7PI+Ly73OQ6YmehuZXRQPzs8vENDccpr0D8X
5cVBL1U7hYC/fTnld8SzPEo+3EW022FgKQgeyAiv2MUkdXBrO6iVK0DK6Xm5X0ll
9b1wTppHJ2sgp8IZ8kb8mQkG4mjpIlyaDgRP+KYS25BA+YBmNrk7URhkEN0HQOoz
okQm43qs/kBvSL5O+igXiIBUMQTtLhcmUzMYj//hXWp845pgxTrd06dGCFFVJ6DA
KpR5H00lS4elPh7HaSvBkFqWE5d25ifWPo0xj/sKLlH2hXWbcQCsuz9MbTY3SPsh
mqyF32f7XwUM/f1sVwTvS11KZ9hz+c1jGLLlliP0A63+KNHtyWw1IaNU7bxD/bY3
dbeOtFX0vjvWcSMcdZqVFQbuKHrouRv9IZqStJNH8q+OII6RbW1J98fM72w3JkCH
vkP4sQvd6A946gwgIjb1EW2u7flX9/SVR/6iKLBAmJMyA4gsbklTDCHKKruG5Ssf
kzFovou2O/57b6oYqanDt4tNU5LwkQg+zvX7GZr2VMMoYdve4wnl1BpD3sojf48k
zuU12NGgOmaRrrFwxaNQWoXjgwb7uWJ/u44nzSDxWp1RYhPu7/0TolU+5waGN99w
s/cnQdMJDWvY9FKGknZ7Le1dKc+QHj9Ivs0I+FHk8AF/BScMKCyHF3GQm2o5jcUS
wRWFzEPmV3qa2HuY32I1KM2MogCOUa59VoYuBTqU6jXLoNEJeT+WazictPLQSh5W
HBDujqGJTSVevlW7mru2ZPT+jRrdDTGweo2Tnvr5seayzoQqyZubLmariFo9q+gK
D1zNBUkcZqYE5TtkBaqPszubkbVb9SRhiPR0yncFVGP5wdBuRsG1ZnaKwK6zMEs8
tIDdMBrcaoX2jfQjgF4YDPisnrb0IGZZ7Z/rJdj8cfXTTI22HWTpbh5GxQEKs3pP
zphBzQIJCbO0uxPpOoRixgB4/IsqX0We8k9F+fEim6tq8T7/M5M9jPNhuNx/wglk
nehoFqaD11m2EPhMQgVR+9A/f8XOxXelTu9mB8sHzRUmncuK8fUmkqcYu8Hz8Ud3
lpWowkUdIWUsMD5NPHom2zeZekkeMKb/B0MJQz3KaQftI3vBBWFpmWUlTdDgagd2
DLx4Jt/vPbQOaNFvQzzoPox231J81o+4OAAEnL7fsWTsYphOm3NW+MP28khR/x48
Sk3fP+eYHwpcf4PEq5zqKZj9LEg0QAX7gk4CVHSA86sYsw5DcnpU+lvF3Y+HpHyR
qv/HQUACl8hECfUcjqCQJiyZbgE+BtogvaNoDVZCqKCgYrLtGBiUE4uCUF8gf5Sg
LQ1QfnQ4udWheEBNW8sr3sccUcAegf89HQjHatykdD9n9Q2fsK6i18EKz8lRgF0+
v+5kzXus5/M7d9QH7uZeOBQLNCJA6wDV5/kwb6njGP4+gzCY9kfGmEFhSEcuIsCi
MVjEkyHeQ4wgNCaNRShe3iVJxCCFczbm9odgyZHcFWE28uY++PpHeU4+XqAqvTPK
lNHKvEuyn9Goz+Wgp75fyMdJBcm+kJTTcjdX2vEndqfFhTKvgQMFGYxup2e1zUlI
ari7lvyv5s0hN4H/Q1A/SCaTfAWC9VrBaJI2+DilcPnEV0gRtAwiz2pUOib2k9TM
BQysO++9Sx4oF40CFUYL+czrdsIpG8IukxaHBtr5hiySRC60MCYfxoTTxJNQDK6F
aguw58vuLaJxEf0DFjhXoSV7JyDrQzhV1NUc5cEk58z8/aUS5LBYb0J3ifG7Dyn7
84nm+9gCkE+TGyQQwZplXSaPItqgH8DU8f/kADWUyrQb5ByC9jZwoB1qRJAQrU/l
SrJ3lxqABdM0COpSC9wlRjKw2cx8gCLF3BpPZpLviyn7+FL5c6MP/BTkgwbjCxY+
oI5UArsSX8GMQi342Rn78sipkqNnHwGdq1bizTX8byj93xcQ9hd7B85E+RmzhTDe
1acgL0pGQTIlZcoy3dG3NStkgoYo9ALpN1HGGSiXGsrB2MENIMATMC/sQ1c6TgVL
2ZGHtGxHYUs9b7Yrh+kEh4kXJZphUrfo5qDX41CaajGV3/dA10j+D5bZHZ1D0sOE
2qoE039XwQE7WoZ3cpSyz8g8hydu5hgQ2dP7G4aE3U6mD6Pp2a5w19yVsASzfzla
N1mavLc3BP8xUMWQAu7vdVCEuh/pCPRQudeblT/xxAe+fEHALbkGO++L0Y+TrZtC
uF/r2PafW9DRwSDDO24xWYnBKamLfx3NCKibFMPOooyq4qlyMlP3C5MuOwGuLhrr
tQGoUvp0bnKxH8kFa583m/O3rYvceJWAJbviBqU5xSAl2F86MIDFATan+RQ0SNPO
p9hFbuPcnc53iH9ccqKpVf44VDgjzvKhjnJ1Ccbb7AEquRMcbQ7GVHLndyv33UxX
O2Rkf5ccJRflx1YnW7VAvqt5vsO+Byx88idMd7VB1wLFyoGiBSG2ugMnPKjJoLHG
9pBMyFDqtFP7A1o5WdcpOgpipYUyY5ctL0xRymbxTLr1gEioZLYbj3pOxtXYTnGF
qS3D4FM+E2v0DTvmUSimJkiHfdTDgZooLj3HjDTD2rAfrD8aDFhNw5Tjtxo7FhEZ
IrCyyz2TP//rem/bGXrKv1jOgkfhmFGT5gYem4Vq6VKc9gillI0U1vwQJ8m/w+0p
Ri0zhpGRU+IZuJDL7eKMFG3nlFzdd/FlepJnEOeIz0/vYaA9KaD4NSkFCHDwkVB7
j4tgPgAKSQ3b4e7aAWWHD76scHYjhM9gWVDU2gx7JYYT1+JcqqegriJc5C4bcI4n
hWFeGlaf0TqJI784JI0/5XKYCKXznpBfF4Wdqnsi5V5FiG6UCVjg6gogIr36jnSL
ykKbzvE+6fZxNrJmH8r7jGLgPKMddAs0eF1WU9n3JEqGP5JrxugD5lhPL24XQg9T
SZg66nZYylbxgc1YzSwFIUT7eLy26WK81FYRL0xmPwXlvLlXmBxX+3+pyIcDEugL
lZ/T4UlKap9YMG09/wosa1BMyfY8kd3OmcN5e4hHRsC7ankS1zsZ5shESP3Rn+od
MJVKR2IcL1PyemKYHIcfw51fgzCFhxVIfKD002zfDibv1ArtIWu/DLwDdzsFwbQz
aUzbVupEhsICO5g7Tmxjp9I8CN8SM5HQEXJMUvTUSsb2xTQ4WU4iR5/MxluICDbv
sV42orqMRoKDe336X7r/pQObWUVgT462YHdrwtmvN2x2J7Hfju4bdRX7i34KmjNB
0el5JC1bewQ8ucjHsZ++LZbJHaoaPrImYa0kDZJB02ZFQW3LX1Nd5qcmZVG4x52i
kx3kuMLwXY9SIr2Wo52c69u2Z0NIPnElaTGpUct7wQUYnUtA5a++zrsCJNV0uOoI
yPWvJB6JIqpzdB/+ohe+cikPrSDF47VciDbfmZh5mmHolLX4vwXh4+23JDxX3BTd
cWKIuLiR9Vuof7taIVZ/ZJxMpk1AvIiVYKHbhlQg8GmqvOBBg0RLKpKOirfTVSBe
IsALEWYSWmyTT+9NNKodeVNGW2YRmPEFFhtwy18fc07FEfdeJelMT4ZP4JC1HhPL
73+IrNOQi94FxQbpjgwphqfNZkqAqw5wfwW1iLZGEeffOfe8X5VzLsNyjvRb8jgJ
+bxqJAWrn3XobSd2TeNor04ns3H1tu22gSYHJxQH3hyt8PsZHZi0wsAeBDItbsJ2
ulWcNu+lACqo7/rhqZQqBF5L5w+eUGWx7s93I96X1x0LWsCgIBq1N5zk5w/cxTvp
Nrf2uVlLEk5zaTrbknqGq9DBN6AqjVUIh+HDfyKlm1BWiEaQ3seOs1t4s4YudKoT
0T0JI9AYh9jE6r44+8tkwNgiKe6N+AUeBf4XcewZE+lsomoDn62fXRQv22pQSCYk
JuFFx5xkiLVPHeXDonh6RQxCa8qidsiRo2j2y3kCqYnlTIRMDJydcxpIVDB0NUQ3
Y5/S04tm5LcP0HoHOSZMF3IfSsczXWwQY4GGNYJakBwA2h1M7uGlqzdhXQY23UVq
WTMVczKLOEtiXthVcmp533R7i/rfdVggYd0gymLtPkqXps8EFaXRSTA2D6cJs0u7
Tnf5oiDEBQcnDxb/cO+15x0drmL4V5Yg4hxZskXms7pZd46eDa9VDQw5noWIbU5T
OhjOb02+qhc1wqWPYgEFZtYkAISi584wcLp63g6copHY5ciEsR3poKEsEtV5genY
0y+88OoqTPVenLLYhfGgEFU74wF6bHxzGW5PIQ+WABBdiIhxG1YVBin1Gbo8YC5a
Ygi/tDxBoqRaouhZgemmQOKN+Eo9o+jvvSEPUSXCQqSiXzuyk6NtGF8keUZk430O
aAyTs3BBlc8YzSxjLJH2FnqzYS9bx/cH2yfWcFfosywJjkKAOHZHHY3AKz/+YMgC
tFP/JO88Q9/ch7JNxC7QPaegy6XghYDYYRnIdptNVMobOOrHNJqpa701mk5qEw8h
wDevXbqeiuFXOzu5g4d/r+/xwRr/RINxdAzzL/fXJqMsuZ9lVzhGKYb/8dh8kTjO
82TblqUBsa3q4M5w7zcF/lHusz7THHxZzwFMLdzLWir1k/YYoQYjYKdFFQB3rmWE
Kgm1PK7mc9bxSzj4/LwRx7Z7yhfNpPk+r8Leowx47ZJ9la563uW1/V9sdXs06XU3
He28/VNVmIdJRI0EYAbEsdNW6Too+jPUNFx0b5Mw1aVxVKntWJHE0q5XX2ZeMXJ0
8M5npPxEMCNWHGXKxNmk/AhB8BufgdU4U4CGTPQWgRCzuW2X6w/D0GJiSmFHSbtp
nXwh8g+jwLu9fsK/qo3IJq7H+DiARuwuR/J+4n3RZO+Ip1BfDWpGz2HgEdqMDCmC
6yEjZpmdd0UOrBVM74kiyPDQTcfT3rJ1Gbb6qF21jPH7DZq2+bQPLuOgYXPOIg8E
NlTGd7v8ljAXnhSC8nkyxXhVL4j7Uk71rV2m6JjCnsajyklt8Mibz6PYXr8t/8Uf
8Q0eLh0Uk4F8Asa1TFyyMxIY2DtTyTouxjBjrUhpk67MQF5jpDjAwDPvh4nEAqPB
58fOVOaAHdLCye9onTgLEPJURObYZoLUcPo64Lq/KWE3Dz6SfwJ1IWkIXy1Utb0l
EycKQX95yCmu18mjGUyTCYvfibNcNJPz9XRqQXf7TKi8dAlinsttRdopJthdHDRI
9OMGH5MAUL7qHTPnnXjCoE3qCwlY1yJJGOyqlIiutJ2UUCocwdz7G1eXf+bVVlTl
Sz+QnEGBInW0ccUGKr1nh8srQUepS/5gmjGmS/nP+xBh2j8oYnbwr/4+uZtgyBoa
UC/L146y+t6+3PNZu+vYQIwtj+AuRmHolVFfpgj6V0S0DJlAauOCqrqPcRLlZGsH
oDHE9GfoHAh47iW9yJ3ZoZC74tPKGhQi3werjbIghB3YavJIxYYBD9vdmY/6tsqc
HkgASqrKSI303aQgh2zPGFFqeph6i4bBd69aVHoinMgE7OMQc7FNxy3ex0B01mbi
mDncIuqfFAg8y4kY0xsTlI4RoQkHCgoO/nRJvkT01D5Ta5R+DmjatfWicR2P3GlF
gzEaRz/EFH5d6fjrsOU6t7je5OpB9pTqD7I++pk+JziPxGqAyvLHuzUWtfJQ1xqR
2q/NLlPf/SFGzLxbq2r2dVHSnpSzdhqqEKvmHQIuwNfwFe3+0dHoG1cPKJW9D0dH
L9GHuAiODU+izqCOxPEVZvWiIf7i+O6ZXzy7yJ2B/IbuYD3J/N2lgPxFqS1wxF+q
tjEJWl5S9omtXwqXiXTq6VcJQCS6InT2mgToch/s4giXuF0YaseoHFr00MyA1OOK
yEJeFpIQn5wMwG8RA2k8xjqVJTxOTtocuNny2smLdyF2+P2U3kBi+l1aGiJUD6nV
50rvFke+MW686TlvCHZECM7Sae3rP1NVbQi4PhWJfTnuJ6d40qxms3k5Om6daQT6
A7DnjTOeYGd30T2EAQtrxN2F3Urs0yNu8WJzCZ2lJlzdB0jJl3m7Ysmyiz/bz1bE
Dq926ebjUI96Y2K8QsNz7GsJYdHmgI+ywzeXEDrqdrNRYFwWJ0WVErNLVG7dojU+
wExIANiPux9u1tMbNqHK3Zc9mO10Y50kdSQddxjBsyU2IQ9i9HPe7wCZSW63TckM
DVVgEnIodIhdHbtFs48eIEKyFIE8B0vKjIEXd02aDbkwVNHDqQD3HIAsOoaVP4OZ
FZixSA7lgj0/9xsWy1ZjgJ7o+LD7p6CqCkRK7DPF6Ph1zGDxOHW8YavvEr+AlubG
cp959a8d9DzXcOhzaLmPdJqK0UolvozZZ9eufxfSf8qUA7nt6mXE4v6K5ww5NYjd
epfBMx5S5xHwqZDFW81PEw5hdDppMU4Vn17hIr8Mptti7amgOj0utUAtOhJjJfCW
1LhL998pWJ0pu4DEZxO7gljjw+47biVZJyyz5oPEIJ7BXXf+8pn8gXuS7pTrCRrN
F18XCBjtuubJm9lrjfMqIhl8KvSo5mjC1KMkXmDYJZlTHJvQTiNAxigVhbu8G0B5
BfxY187tDVNHZ4MUcB/62PqqudmATUO2JJ2glmglfnBdqSqkbcRCCIUWmMHZRAWz
46knMprSPcZ7dDyKlxVLKca3cerKJeydtZ7J8s6vWcTPwnItiII3gYLCPIeLlHWr
NSCPvrJrqgTpAZUwgpNI87aU61SY6plFmXgfIrB0SxBtb6d2PafA7JdMlZ3kige8
WenztvQgLBfYLZ2QYFGM1H4TQLKJ4NYpIwfpvq3Hbn1PNLbc2KgoCMFadQx6NDTD
Uwngeww5Fxgza44E9qqti0Hn1aX4Ec888zD0GCt7HMOadBMuVA/TOjUbfqBo3M84
DzvelMAtaBngmvIzFN0A7hvzD0gX5jeyD9VnJnZxTf9fvTsfnU6NrqD9m0aWwLbW
v5XJRMnReFo2EqkdBMeVsclvDhD0JW7Q/bg1SLezxTbUsYEfLTAB3OHQX8N5Q4dM
681ip7LlFFQNB7j7qLVad8Xu9sGeEOrWdRlvCWk+1FdYlYvXLBZhFMf5uZ0ZFPx0
JBQkJakd5B2W547nKs7mm7ZK8yNmfb4LkM9frj3fRmnApFFmdxuP0R+voHaThPgm
iDNR7iT3To7mX+4jteJBD3BKX7QI5VuqUFh1qF0PyUIX+iBHTpOVBiJJ9nUOZ3gK
QfveJ1yjH5hczK2EyamSY+vMaCxQYqXTKAV9ZsTWbNL5qNpngKOmU4Ed5vL2Kzrv
pJzb4W0P6jyg9agMmAbrY7lAlh71SWGsci87TwgHajW4tQX4zLFRU11oFe9KDHXA
+pX02PGV/HYvUueC5ggpaQDE6emcGgAUaFCha/MELTuKsKlSL1ytSAyL7OzXzDRK
0Cid5v3tm9f28lg9bNeZukIUyHvLWy9zl7Xkjs/xlUmkstN+ULuUQoCJ1zKzzid1
JCH+mZd21o/m6CBjSvOG7UkzaHShF7KOfx268mF0Mh+KTzjsFfUg+CWQX13jG8XW
j/+1EhSvPOtGT5T8ahl8OJou+waVOdjjFPfdxoB9VZTRup3pYw+Vx/lIyWAEd2kK
ZLXKciGrBfNYS5RcEuieMmLtRDB9119kfi3mz7fGmqj3hKTh8TVrSoS/HTntcRCy
SU2FMbssg9qT3SBPnF5sTMBEXfbhwCqT0BBhEYi596JTDzIH4fhhAJDqRvbe32wT
efXZSC9bSNTAMQChQiBGMmS0ByB2P95Ke5atNpqOe3XU4m9Idj91PQ6j0WcTZ35k
YE0YlLjeDxrpdY9C03ioPCA22v8k6FgDP7dCBnS6z8licHMzF8yMXQKPLDXxRsQZ
Gb1D15MOr+JzG0eJODSudvV1wR4nICTaKZ3L4+/C3HKNMH1xv4esFRPoXvI0RCTG
7Ujh2C7LhZ6mSQ9HHDm3gTz1gBUHtTTGe8xw0wWRqCyyVFvLAjHAYaLDM46JObKJ
x7UK2xXErlNSD6xDbLYXNp59lFKH1Zl64I7gAahoeU0i41W+OI58y81r2ooNtH8L
del8necyyTcbt9xH9A/WfaAtdlxQfu3s1TixFiLxDgXoKGe3zDeAbAHuz77VgkVP
JBn7eLjKGdXOWpvc7jjiAkSAoOfwMCLbhl+7s14M2M5FdKFBOtkNk0vtSg2hIAgs
R6R2ZCJHgUYvJRnU37OIeUsPG6AyyvAJZGwYfepYK3WkpxYYqQfuSNPuZXh8ag+U
kP8D1lsgaJ35Pub8aKOV/9vMKh7sJ0vHbjtdOoyDdqYg3q5dkrdekuONUwJUgWGP
26UEJelh3hYtGBEBRgXSFA5tEPYJtEz6YRjjRumD3Y1rtTUKmlTvnMA/tx5KmdNt
MyDJRhnxbfaD03Zw8qtO/f/wqv9CGnQ40BQUeRu4nAvU5Ou40Qkj30tspPMQnqEG
KSjSi+/eooQF8vAR6JsnXjRb7k2t6VkWpe0OYnCtDIJ70wxvwW6QGtV5fkpii4Mv
BeZ65aTJCntGfE8lMpL3G762AwkLIVH94SW1a0PjEBEG2Pj+AYyp9EFTSWpuWmgf
51ZWldJj6aCq1Kn1jrdV1Wy5Ll81C3Z4uKqf3u90Mmg10aSSmUVJr2biFiY6Uu9W
P/XbVtR1ig/VR7nZltFR9h2OITYXtcRT6rgIp/Yo0kYwCMpq42IKJwUZ26VOzDFo
U/sx1eoY6BGtMoozhyE20wUnEcr5EP3HbPyKKUsEQd+M+Hcnj9hbHWoLVNac/WJw
NyhCgOmMpDfdaKdMW+Ud/V9R1m10RescmuoBKSR/TFYeqqQ4kFblce8XwddtVcjL
55Sq/B2Egp5rpMDyf5EZKRLNPCfE6v9loognJTEhQJNg3jH2DuIMUFs6yCXdQvq5
ciSt9A5Xrp3R7z2WUrMxnKBkNvmLhuVbjYspwD9qrNxK/1MTe6HKk0yzF6jUcRy4
UE/Nkdj6Y7Ru6n2Gru3KSOjbxTdA38fKe1m+F38ltbHBNRpChT9CZpbl+lAydfg1
vg9oCTtYatb+8AJTpso7+ejQbLyxDmp+Yekb1PmMhiMQTRdAwS3N6fAAmiWBmCkf
7EqlRnA4Fy53fDWz7dLyfBZRSefBKNcCL2dNtuuP9muH/RqmnWrzaNjTZQjOpzML
IQ062AI4lbIhIKOsIbJzyqh++tdEqo6avL2KQwzlk9y98c/UXQE0bSdCPm0TyOLy
CHrOptyuyjs5kX5W87M2kuAJZyr8xMsDMJedhmRJplTQUwYKCOp4UEY+XfYZZ7KU
YUmxPG7qVTiFU2P7TPRp654f6aFnIzbL2NQzE+HMd0Urg6/5wrjsvIlqS8RiJK0Y
Mmh/NDFgajF4PY+NaBt+4kZy6w9mBWzwrTmS9fvu2+QZCsqSI6uKL1doF3m6k72m
Pvu54i/Yq2sWCSWeaon6qbpLhMsIYDlk5NxxwM4vk7jO/RYp3xlYebZJrr0W8Anp
oW3VXs/yyhPVzRFCP5Qh8ltbs9MPdRModMkkbvk76D7dKLXTdJFfVOKOtVw9BNhM
MhkFBQ3cECioz7whcZjhxLbzAqDuH0xkT6sc8Esr6EYMUyLcEv6rdfUyiEBU+Guw
2G+fKXZgeaxC4EtLlvDPtL4AQHQVDBA0MLfB2RUYNPGcg+BGxJkSeNqAJbwhj2On
CrXQfTNTXqHgjba0BCOagYX2HtI8IzO7yCUsiOLVKhcZLX1IIv/rzo6lT11RTXf4
Ln8GLcVWT4IjZe3oguBeNzSLEVZKq5qU5fkHImDIHQ+IHneT5ejhe2LmyutbITzu
jymadW2E/Rg0nky23VdTMteH6K2mJB1corgJG8ZRZZmKtYmGaPi13010WrFpsveS
efPI6/DTNzRg99hm0aEci4tns/qknwFzx3jIh0LnGXZHJ3Gyy52a4FCoPV+b1LFR
mCn+PssSAzxcwvyOzvoWMDIdZs4RhU/CTKDYJiX0o1XwIIJx/TX0+57qY3I6/TPu
MC3HHvLOuYXoljo4NXouSCjgnlcqSsmt1eTnFaCpKo9NAcMy+whaBMSrt7+sPhHA
SsPQ6zq7o7vewujCFYWi8CfR41ph9r6Nqp91NNXqNlbTri+CUkZi80Nifv7B5rOR
nLzy0IyVzsEc2qlkyk1DXwYWKqpXHlUIQSaSV1Srwv9brtI4ITniC0RnK4eso3/u
hz4vEsDP/J9btwtOfSn+h7V1Lh/jzA0huiOAC3piXav8pfYBpI3cRvaMLszxnhC3
BUw7ck+yj/wYfBPlPvvaBfGzkhsGmxHdvxa8I1ZEbyzGV0+/e1cqHFo2bXZRViwL
BUSlxGYDRpyjsmVx0i0xvnWC/iBHD4Yqe/ewg8MJHG9lNHXIupqFwXuDaoh3ozof
n1Wn0jdWD8p2f4qbXNm2lt9d/swfkiQCHzRfIfWDHP52nZvwNKXKJwMlz8fPD0pb
gARzKiL08xpr+if7tV7wcnDmzh65QdNeGqLiMNLtLr4wZaap98hSn7JR3ylyZk6g
h/30cFn7+Dgz89gOuNt/u9U3UgroBc8Hz6nKLsSOygFURDPDZoiKwS1Jt65xaoFc
53bKFVm6CGyR4RMVBDxMtVNc4L5WBGNi+nT0OpDIifGpsBxgGrfEAc8ii9Q3nf9i
0Kx3FfE3aVxiJ9h2uqeHLN0Dm2SNX9k0hXuYMccFWl1zomdOAXNDockEZlFfWQiR
33xpU7PQ3ugqn7SxaYdXPjXWuUm+sT7MS+iWeMOyM1PSwhXVbrHmgyriBU8kuG0S
qh1t5ZI0Pg6+2AKeKkqgWhXwfws2XZZKzw+h0tzsN7zvZtMdv9efnVvECkeHi07D
U3SQlcNYpQofnxqoNsAhgKuxHR3yQKnkrl7eaR0m0kpmS9piLYusPbWJr3enFmnW
/2jB/P1TbJa5GWZHGnHfQQpGb4ITS40KKAr04MebYpbfd7WT0oduO2Gmlggoqhr/
/UyTtKYwRm7ai9b7o8VvoDuVVeHqlNXzzSGhpspKjJJXa5GnnTtLFGE2TXSK35xr
TuY9wfkE4aYJIdvWkGqrMPagVNRzUj0+Hga3PyG5EraN7L3E7I9zLLKlRVuxDzaL
IEKHCSVPatcbFZkx22aW+pgl4lbgoNRYuShMr9/4CxzqvtZwfPzmP17DKXMhjZyx
/cepK8iafo0Ybc3rv5CS58QFcunCTr0jRMEjLGo+m1TbJpR5zLNDKCO9WkDYO0t/
W1nIBb/seCqDGg1y8k9G5ugkHByyy4yHpLRppsWacI5VgUjTRY6JAx4+NYDnhzTc
icwKEs06qO/2SiJFxzMcDC6vneaK22+nJ4j0b+9ipgj+Wg5c/4XP9KNlegMcwtZD
U8TIOg69LQr+bnE6RJsok0wy2qLETQxTmUVKVk3L08NF7hCoAhiZNlgxwDEUidSs
w2j+R24nVbLOHVJU7KdtBXMDhrsWCAtmHV+Pgd8ORu9RXZ8/SV7owklz08BISlSz
qZWw/I4wcTcMlB6MvzsCHvB85xrHfSuLicjyTtVosCNddl8RkJTipEczUPc4xAnU
Rojc/XsB1/5wIigPWgpZGOa0VDj+zx/3oQhABOLIcEAu9uj0ixwKuK9rLeMqtlkt
9RuQEko00O5P9CfjS1rxGOE3bEv3tYe265Gev5M3IPXj+VRLRCLyKZEmu4QVnRQv
Ta8VGvq2EpW5vleOZ3BEzVrGKr00YfBizCBg37M5rwf5Pt9ovLQdXlzggFAQ3Oy+
oLD8WGJEF7jyKYg6RDdJnI3cv7xJHxLewF1bcmmuyfVX39BEtBsHBcj90oIdnN8u
4b1ZOszgipzaAWa/+0R3vQlkLDXwuAsNnwlF7mW3u7e5+Odn2jeZbqUViza6HjuX
yWqp0hUtjKsa4dRxAUqUnaylkMYrmnlBczGhtHzLT8UnDRLiUuJ3x3n3f/Gzf1zZ
OSZZSNUrkaiXRpI9xFaZ0dqc8wzsmCqaBIoGvQfX8+r11cFINhg9eKGi6Fz+vitS
lXORX/jzXcQVclaKvNVSlG2oxtWalL566kwyxntF1LoAOS0zxf1eeynJiP3YKylC
baqYLfs0vzy4ZPZo03H//Vne66vyxhpZKkc1q2N8Rj6KX+VuYZW/r0AudwmUXVQk
fqiumlYRE6aNw7DbrCCr0tgtAadk3DNHWxYqTTxOKqgWBBxGMHwJWKsuxd0of5qX
YlgiMausv1tDMEh4b2+zGkI0WWQO/PM1jbfMy8rXeVNsPrloK+KF2Cl1bwJZVGCN
6sJyu/+Ia01kzGZMkARBJimhXfDtXJ+v9wFUIk9FpgijufbPGJk+4g9uO1GhXhr/
vTkpcrIXMIC0EzXnKvxZ3QMNqhKbiSn5QDnSrfUejfYZEeKKwj3voJeh5LddPa0N
IiCeKLhf92Lu8Itonh1Ixuk997/a2Hbt9uztHjuQ4M9mPbphsktGbL7Xwx0Xt0Xh
1V9GVt8MRMyrSrVjqdP+x//PiV3D52Z9+Bg1+DqjwJ9RaRAzteQGwthU9DXstFr2
G9W4X8yg/XJUM/HNEkdKG7IXql/OqGvvsuIOQ5W4YVpgGcDILovnQmnigTqCdrLB
uUCA8AmbWjk8FeUM+ItKlgA5W9Hw9IitEdibqT3Q06lkO0ZoAcQ27PDARcuhQTD+
xmzUP91tDQAhFkJqfqZbQRZu6t+5je1MXYznmwIBYgd0GEO6k0wMnNSw1QDy6su0
WpT52Nf1mq5yuds5FNZUns/HbXId4Zc6oL4w/KBjPEknsQeoyaoBfQ23DHiMzleT
ymqwob+zGZimyM7pftPBH13KTyl/Cy7k2LfnmTBSAMEfSTpC0wKESRM+0sDeWbdJ
P3Nc8WeEAX7fGlAD2uh8dRUXZ7ao2qo3RQxqIEHV02DBbrYDuvZxDY50RGUABbI1
AY3s2hfy+1DfD6JJR8qHbxc7tkciMkst4k10KG1GkewDybl+SSCVgEToImUTvw5c
KKcsB+0nKuNkc9ndw4tF5fQxPdf2K+h7xhABqh5bE/rj31js/9EctpeffZDJ3BD1
9R6APAZrfs9KG9fKh61xu8GVJYgcu0iE10VXjT9ENDqHgM00Hwpcn2/njRQhtPm3
F40JuHDA0pGOdJXB6Pu3mCje0YwdBMn8lOntDQ6z6mbK75X56UG7hK1DZCybQ/wn
ewsge6sBYP5f3bvPXcSLSVmUHwoLsQqy9A51On1Evhr73rpFrT0Tk6BZlSRAIPrD
p7vyyS67ElAGLFr8XVV2a1+7ugfA2wP6sWZhY4jp8Mhs6LFHAzIi6klvbEBjYbsH
X/sQSBnR2wg3GwZ+T3JDV8/4uHJIX1u3h0uzmm0RRdwibS9GDXIF5K4lBvUL09+Q
Vp8BqKE16XhIz43NSjxYHgB6cJi6JPJdlwg2FHcUC6cSvM+fNXFVWX0bGzIldxHm
gZiLQDQKmcixzUJYw42QduPdQT/jgU+PuWHIIJBHIkwqB1oz6QqbE/WcYZIzR+hc
y7t2J4k3xFPMDrhRkcNpEsa3d99zuEhnRL84v3ESiyogXLE31xDdUA8/vko9tafL
AhK1gUAyCDVg4U+P7hPedAoqhhTO4DpMjmIcV4dym81tWQ3BNot2Z84MPH2EkVHW
x61ruD9PQaI40jrsHZ+qrTpYKxOBvKcsmws9xdDTsOUhH1byBrxpUXGVZswf8m+1
kJS63Le2nSbEs461nT2UPRS5qB5qH0Va6xG+j2dlnyZbqGnvCFd2slUOkHjXLkiT
MET/1y95fHCgk7L04HDLDzHsVD1V9aMfsTaueS9erIxP5p0KTNvL7yERLoH4Op7w
fS/qJCmqlp/6xKfHfusX2Vgt9Hp4ChejzuJk1m+vir3JrwzXqjvNfsWnOoZLO1wo
6nilrzgv/LoyueyuNd/fEfmxoBw1XUZYygeBydP7ON8AhTKXLZnyCDuGQVWbzrEV
ojfCaeM4vwRV+OZBsO0aQwMvSbVFYUEZhMKrz1uvsxBzjyv67jyTyoZ7JBRNkAA1
GVk8PFwavHLIQK8n73RiAD61bQ5qo/AWl2C1kvCw5CKC0pWPmKYfJYJx2CdDbRkD
kWBbMu8ffP+bvgIyHxx9GT6QQ7+F7AGJ8LD2M3OlH+9pBlC6d5+5cm0Ff1rB3/Sf
ZGqEmXL69SQLi9S9yEOOMmjxbYsBJIYFTFPeFXWpbdUKhyt0SO2q+MdGii3LmmnQ
eV4ncChPYPE0L6xTN4QgmbKg10WwBQSFCAWaqDA3OtrGW+yafcjVXAWdGQJ4H8Er
Rq123YBUSBrszf/4HQU9WqWntqV5cd7ZMP0P5xe0L6xl7KwxdLHmygQwQIPyoplG
ujxh1GDbilb0k+HnT3PWxkswrXpejFeaBmB25H2UgAXrcDX1c+LcKh4tLrdjU7k1
BidmtxT51GCAyGxXxrMiIbhOtVcjFaSVfe7/zrNwWpzQj8Xqd+ntA79y0RkxI994
nH5X06N4h1HBvjn/YQM7//eVkNknLOFBVMEXXU6DDzEq8joJ57oxkgTcr1eJRKcL
mN+Sl9zyTaWiK3Y9dIbDIAGva/NlE//ZVjfNZWHQjYBCimcL0to7i5/05Hg3XdTp
EF7UvWDKeAB9ILv3mBd5kE6CKWmjsfCwH4jOEz9QBWGxGOdcPsNUvtshrhGui/0e
d8e/hC/39lB1UM1emNT9Y/5Nf1aAqCx71g8J75Ok9dD1WOkQNQVaqNeD5mg8IzhQ
QW+KETYGGrjO6LG+euoilpmLpJk/aKYoNQMjLoywNZA+z8jML4zX29BFIjG6VeXn
LwXp/UIdcp0gxxh7H/qDFuqhz+jOMtUKFVGj0p45nZSKHv0s2TCUDj4ETQGiOqaU
PJip1Zx+L8MCwValYk0Kx5gkpGI7eSw6cbeV4SjngeRLfOzFS8tFK4PJU+oLLALV
7yNegsrWXS3Hmsb1Ez0E3oBmedwzFHqAyAAjBAyqRBjDLnm8uy6aisAODbZiw3pC
T/naaJaFmMSz25w3Kq309Np46Nim+xxHThKDcez1f9pAGHn0WOTRLXpJq+CQ49/l
P0TewUFRYsga+o/GH9ZbGj8MZdQprwObD4mjF6pCtCBijDd+wYBxmSzoJEvksn49
Hv6ULXy92XxTl5UDipAe+kUyyQGj4v8ro5ZLeEHMS4X1FpYqGKaOulX2UuiiWRUA
gCJs8+SQoMVCvHNJq2euLa/eEicUtM/voohEV/oGO2Ggj5fj6sSBLZcTdYyCkwPh
SGVq0efwFj1vXfJr5xTn1ijk8ZLlz6GoR2Gd4CFfb64Ul16fLqT3FyNFcZLxx1fs
ZUbM2v/CygG+VkUOfY/cRDT5v9QRmNFuFvjW0dErc1z6PV8d2qa4JUf8DXMexvNJ
g0XhLm8vVLpLy0qBOUcodIJ4x+ySiCyK18ZOKVashdEOlK8/r4AtIWQjFIWy8P6X
mLQ+B0cB+G4dKzVIBH8W2vFOg5nV+o1UFp6D51IHJ44K86/stFfT06vDpw22DiMk
17oAoApU4d8VUz+OcWT39FZ0Lgh8OKBj9ym6RNz59DwAN2WOVzzhBb+KwApoiQLT
99TFVYt1vv3TlbQVjRqGbmMgV+iYAUue5mpcrycjcK7qm+9FtM9VdzM4V1PlEdW2
NACCjBX4N3m7/Ht/oostaNMSRzWFUsxpLeZISVmpAgL3hv6b3Jh45k0WWHvGVK04
plmsk7wOovmJ+WRBaBHn4KBa5B8BRzLj5vBJfQhUIkqex6L/JSR5UBVKZwrntOhd
EaWKASRqor2H+GVO9tNNT8SvUlf4iM7L2G28M8uObi7RHCQBOIflEWd8jrplrAIx
jp7OIaO8AdxmWf6zlUzE/a5Q/xTuxaegG4hpGDZFUp/XsDOTc76LrHGaaNUHC13K
hmopXZAm4Bk31eWfKj5JtIC7/9P/0YZbfgTCjFQsoRtjmKdzUnhFutYsE8Eai68k
XC1vOAjtupRTzv4pJu6yKduYDEORrhVI+SYp+k7JRn+E3znGvE1awFQMtQQvYz7L
4M7zZuMyhs1F4r3sTocOMBVyyEHdrXGj74HmcccC4tQPAvoAKpCS3yC8IMCFVT4A
SeWsdoKtrEM11W8l8BJZB9uadTZEWbiz3Y2mQfnAC9PYpE6U4RjNbXzf6VBObWfG
BlxQG/UaAePfRvMhICpUInow8gq9wCdlMJzyjVKvhm/WVU4f6DZkxl4HZibKe4Ts
9c551J5gBhOgNlxXTIEVT1bm0hyrddATyXMEFF0oqcerCMAPW/vk99ouaCr0kQL8
av4BbIbWzPrm0HptE45KLRqMMKttAo7h9kRqweqL1BG4YIPy5SKLbKlIOMOJPzwq
SdJiibHNX06gD5wWcQARsWW2rX3UgC5DCqIJ9h1LYLAK3BPcqMqvkQTacXpHDF1D
Y+XlMIF4/gCJo+1bv/BKqF/5B7VWMSuqBvDTcv0kw63FH6wuU0s79NUUf6rEQGp3
+WZ0tXeJG0K/8vPsLC+wlf+vlSyWYvVg6GqBIh5YKxFHJV6AspWTs4waC2QCNOmY
29pVYh+tXo+vir98Etmx/uAYQR8BGNUakoSIA4MBtyD6RWfFJKEqewq1EedBIPLS
teSTM9VmbTnvMNbs8qPQNwYRC6JZf9Bm9Inpk/5pHzPQdm7kTaVkMTEwtBdbXhVK
wPHmkBrFAPt/h3NLmWtOm0HjRRnlYr3ENgIAkNHYxZBvAuy4Th3gk84x3kO8d89r
kF5qpbet9wLdZuw/zpdJiCGjFqim3zgpGkUcQxd97l2ekus0xdbpyIORfXi5nWoU
/NrDaIHMLqbH8DrVDNDClZi74FPiuW2AMKVkf0lMRkYA/62Y9Ia37gvD9G70xHHB
qpJNxtsgFnPh0ZNfHbi0HPPThNtaKrMCTuYRQkYlK5R/7EV6Wgym6cjC71AaZLln
kCg/R9jBcFJ9qIdPWXUM1if1+sezi5htDbUKX8ia2UyrXNXOX/Rv+YKoMtP1eH0P
qXToovaiYXIjAyhqzG/TUW0SFDNF6ZeKSAn5tRp6o6jjtwfz/qlglL2LcElTiI3w
ewbqrESHMsFOUVH96u90kFDFyTVTGSdkSeLYmT5qEbUsWHgIcrxv9Ih9fpbelMMt
Uv5/2XaS9BNr6ZuvnmULcVnCKNdIvBDP0j2ZlqzMH9ULbYTYv22VjjK0GJvlX4a5
C/NgsF+SRAhf7zQt97x5lqkDfdCISutH4/n0+ecC9uN4oplKllKmvOGypkMw1SH6
8K6SnzzXxs1CNVpkPXN0kUqo+aRwMhv37H1BhYSgo98G1oSweccETSfKx4Fwt8oz
wRM1mh7h0+vuyvEoRPHdD4+1+sXW2Nyxfs2HD8NMIJm34J67NQQcrGZ1EEf6hACS
ngbS9iffFb0jic7dGlUSYzOXfkDnIRk4WShz3fwBnW1PFb5L61ZwSjPCHEq2YyB1
m8y6I0YnpbCDSnES5iEZo0/rfGd0fjIz6Qvo2ImQgS7X0pUf9XVLbIuTQXKsx/fH
7CM6SCLluIcIxZ614bAhtZXKh3T197wqBKQ6hW+c4Oh83pT0m8QFLQ1MFlyB4kIo
G5g+rTOjbJes/geqTWj8WIAUKafillGmZCyKH7N2Zl8rviYu5Rh0ZKvG9bSa4xuX
PmrDzY60Th6RNFSdnFTTfoGncFmAOq0en/bs1XLN29WEtKFHifMH4hdMPw9oLIsX
O4xWKWFEAnuPqa41qSKhVxewrz2g1YgbKlPMQdbg5j19FDUa3G4meXZIjtzBG+qc
OTNkbL8wvwpxlTY5NOnscZRMYl15amDpGToCmwsnAFSVRF9P+1kmWsOi/nEFUqEg
SyW5QyWaJIggwFyDl1PS/O4Q08S2Fka8mDnMytvufQZ+au1DcKU5k4LZCKo0UNvQ
N4DE4ct3H4w9+B16w9IsLxtQCvl9Hx9dap7ftkWxUdwOAqZ3v32Ovv5fY2GZnueF
2zDLSj0HvdyHj7IgA1Eev55U+zeoHYTDjNmgP7X2u+9ALqNDoB+3WSdFsvVgzsYF
pBHcAH7OtatiXTdmXSbq+AdDKbmhIJI0GGE2ZHVjj5CsJgtqLIVYLqX3piLazB0I
hIkxPVJZ5r3HK/wlJc6J2AN3xb8VBl7d3hDV/89X9f3j1t1wz9onUsTfhBTdpRE8
fNc0AzVSxzFxyNH7U+bpH+JX7H913pCUeliwFgGEA1Ei0Y0Px4Hvlxbjp+DVFZ9t
QChUKoSFigHdufpZNcRVR/BIWcWQjDb+0o/qlgUK23z3s2Edn5p1rKfJ4Pzt/DuR
w0q3lDaYkmrrrXc2tSkTBMVJCkfpIFp0wHvCKkt5R1TbkxijyRnsJs1sK+9HPw3T
qvpmCqR/t1kBkWewGFyo7HnnRjcXEhtCu19cydUFfK0EvL4cVDDdSuBTmgvX+N1a
XbsjVVEepXeyO+JnDnyq32Do+Ao5ni6Kh9nAY63pfh0YmymbyJttUVzosaZvEtSe
hQyVCEMRmpZBb7+vIARqnBDuXL3JOCN2Nt7L9XMOojHOj/pTmpSyhcp2BocvdKfY
W/Ysokm1VNQzXtb/9IXw3nUs6qCs2qPE37VeuuNQXSe9hha0qGCys7YEBQeM0NsT
9Q3+O+3QXFi6oueIsBX3MYjV4Pp1bZuJWt5YyvimRAf1lybReW4bd7qQUB922DuX
rtYVn1ZPjXdrXBCgQiBQRKVXNgLGRCBohrAIRo/Y1/M6gHpR5Wxgpdw3HlH2NVpd
y29gLdXe6girzvMevJwk17KRiJ7yf0DY2PMq0bn7AN4p4Pv2U/fV6UkA2XiLN0Zf
IHiXIcqQ/PaF6dMkfDUbtD7dLtMSGfvH85WYljOyjOqwXf1O5c9jQMxv3Ifw0Aix
5O6jtij5rp7CCfuGxMv9V+6tV3SaV4VmEPZkvFEOXmHxzQnu18kDQd1wH90uQU+y
IraJqSJ+hwPxAtokyvohTnN95sowrC5lGSJw1GGrGiq77HzNrux3Pd2o63SC2vW0
Gj65B9ryoL5rkvoB1P41cx3RyZDJ6yYgAvXdcgDJApG3wcutpnryB6xmZrrFiSoJ
hn+N2RN+lfM3qYm6TYg1rpV3scB/oX1rt1JWPUwTcCLSq5DiAKLfickCv7ZH9dWe
gzF9XJLgAAuta9YkSXSvAd5XgkF70FMtrBLfYCqU0jex95hFXX3DJaq7WSEEJ5mX
NBZctIieZG9+EpjO9ZQtHhfpU5jIgC1JTg/Bcqd7npBb9jKLQmevQls5YtAijGVE
x/vi4gPtzTPDgn13eBzRP0S7LMo9Cb8vyHE1BmXpwUdeXk/P63PEoeK1MP7aFchJ
5V0t2o+u/nEK4hegwXEOO9KA4W6IvrZJfboCCjiaK/NImtxtQKHtahhJ54D/67MJ
Oe6ysTeYWKWZ7X6AHH/7FYTKgSFNl6gSBTcoXBzaDXLTpx/169eP6h7kUV6dKR9Z
xDB5IRMHvV6m7ohR2O9MvTxOfwATlrHViOYVT5reboLt+wNR/z6EwqKCrl+2Fo7+
Qb0QCU21fAyjlQBjlO2U7PiGe1sRtxHrSBX7JpEZT8l2/NNIzHKE3I544fZbG1v8
fiGHLswdkdVvyITiWzqjbdKwAnflMgcVPRurAl2hrtHyMkDGvr0Zly4M1JBTVMzV
7oj/kKC0Eh8hLstbDWmzCA1l2BJZDX4FaWDI/iiQ90DMpwsvUvWcbiORtDy+48fG
uUyXXujXZQGENYN8+iSRBIyHhhhYOCNDHr43Xrqe0+5HgwQ+8TH8hefyj/vNW4eq
SDLEFyy5HEf5/j1Ek1toZ81g3AlC44mEuVzCnZ+Q9CtX30wz+rJJQrGRHH3UWk1l
9NDTtY7AoqaCZRwz8yti3QKoT0xxRN35U1i9/3ygFZzNlFbiAs8jXaCjVTj7N3xD
hRJeZ26U3/a5WD/lwNFl6RFuhvIwj0AoM+17+JIaL38YQVHl/nLcT3CO7YABp4bm
6L1yUK6Gu9+oeKFBqi/Ik7WwLowi+9y1F6G3aKNjFbnxH9CaibDrT/3BjuocQPAq
7atFoodHxKMqZHxqsC3Wl7h+wFYBOqjYdiv83aMUnzS5UsCHLlhiwACTyRR58HF9
ap8V+m8nfCgLZdF+FfT3qIbnB/MTVFGEwFOQ8wmsz6jMiW/HTIvTamZ41cBSe+K9
Ge2gBxFOHttO4xxY3/iTFINZAQ5o2aOz6QgeegZ62gV+uAuFBJsuKyTt9tw1se3T
LPRwunxDYexoGh01Nzdr/sDeEw00GVLCVqeBF6c5S0RpJqiQU7nkfgHoi622zbSy
ad+Szg+4GZ8Wx21V8dA9EWKxtAHu7iJfqLQYezfNAUp2+b1gUwmUuCmsPK5yN2X+
fCeW8hwHBUkgYG9oMa9I3is9wesl5RjPrJNncUGjSqinLaM31dOHZdzsf7vWdnKB
FgCnANTZVHcS8shoj99Vg0TW9bfbOKQoSoBKF0qw2aunIzJiE7PQ8kNLiYEEbDhN
EPqBumNKQBDzQqv5Sk0N8PUz1f0Qzn0TC2x1jUmX3VPwSTlSi64ZaqA+aCmhie0D
jQyxoR++MSb6TkwQ3MC2G/Z8FTYUgwngfP4KLn+QwhzAtHDHVN/MRhUBEdsjtMG2
1HS4xwRO8xYs8suT2x5L0MCGb+S3hDyS8oO7U39Vt9asO6JXq/Sjsl7uByccxYZH
Om0rntTL4JsLKIULySma8dZ9KJ3OiMrZuvGWmD5dSoMwrB9e0CFTx79CdrbeMBVk
qGj4Dru2UAx847V65rh6BbxFr7zpYkxMCzagbvdIP1Z0PsaGtKVH0wZx76mE8ZuI
oB5ll6uySXO2VdI1MGkuZNatXKBlXD+eQZ+iFpjElfjCK0p8MsrNQj4tYmhyt/T7
9ulaItEDvT4KqaTulDKZgrLPYoXDLg5odQeV4rDHRv0bjTbaqyFG4Te/m4z3kny+
zHXyVte3P5wdSyJ4ez7KPpSmgxrHr/hwrm+anqAHFJcsddn5oKpkd3ExMmSrLO/n
rnNU14hSOYIxAmCHISvHjLkMI6IIQQEDARchFlB7BozMibEvbZQFN3DvVeJWSTtM
J9+rZaw+aBoAex91P0S0cDc1J1y6mD6AoyqdsvJs8ULb9SaZfTk+2VjjJ8KWSwoJ
+LYzKbDWhkv26hzucZtgTUcfhKsDodWn9pw/u6elsR9hHq+Z5nhzN/Q6RDkro3H7
AGKO2de2+jT95sCbOEhstVqagR4VoiZ3oKjc22gDC216URs/x95uWbppCz+ML3Xf
k+RY9qdXRHv5uZth1lk0e9HIWjxVpmQ97CE9bwff8ohAeVU42hdfRhGKBYagt7xg
eZ/Eqn5eFXnIbFcOkaVGNIG2PJSOavcv/LiNkpTsT/N/5lSRNSJH+cO6TrWLKbSv
yfsAvWlZL7AewS+WEx+Ps1h8HAeXelq3iItxxec+z4Gtl7qghPsJ6XlXfM5ISfCX
G3wiCgwBIZ7AhDHg56uTQIZgwXdrqvGZVGCXos5Kd94ZsffYhYxNH5pJatsk8ZyJ
qrb4hbh0XfiTGyILyhgDYp7169tZALE0z6QyH+l6GuR+o+JV43Dn4T7w2YR4fPh6
tzdTl+cFp4BoVNIrEGqsGanHtHnk7reUn52wmIrSWRM6eAN7X/aMYOv3veZdvnUc
KFSQAmK9xNCOq0D/hgj7AM+0/Zcbp5isA/rzWgRnvHscDJvHMCInN+CmLisaNzF4
0sXeG9UoOLmTG52sDK93hrnYRL9pXef7XxtRVz91Cd0DfdIgjm9O2HR/Xav6jvbN
r371CnJTVng4PJyR8GVcpB/bVICguQixznG5deaIyeDY1w7RqciCjWVR9SyFRwuq
2W5C/JEPDE1bCB1xjT6SOzYyC7mb74YYgIpqXZH/ZygYUOpzuckwRRYFb9y/kGzW
pRpfEceSCEW0jIIQ991hwRWp2piTZsdxkzaPwdhLMMkPRU538wDD9/4J5US//rJ1
AGn1WTz1NF4H/6Dfalh9eqW8me4svpW9+KlFt5nlupLG/1ok9UoJPhfkR4Ix3vaD
g7f+n/N1iwWZXxl8ZmqSLjGrIrW9ZXfxTb3+p8DtfoD/UVxiIRBAqgK0tmeoSir6
vtGnWdQJCt2vZA6+oNuu3aqqxTLRCFsYHEc9vIqkW4J854EffBXkeePggeiO+d6H
2BmfTN1PhBWK3dSD2zozm3OaJwC0nUnUtMIvqmOg+P86rUmJNYYYWblsED6TB/Ib
nk2+H9CDtyHW6kn8RF51JTVASiLSZEEiUgBklJO/fKFXrstaQG/9fdfHgFEE1zq3
dWxTvsvurqdeYQZUKM02ywM/4d96FaF4nCGQyCMKVX+UahbiWkG6esze/43S+3l/
KirVBD3wTb39ijJNdxGcvd/xomybWFT5g3A7ZkKE5alyiUbROQLDRkPI0qo7RsOt
a8eh/qOKFt88/PD0ycLQZtL/87AhuznnnheykOapfO2NEULm1L4g9MxbbIcUUV0f
EawIU3VWMhjreNkWAvn7u8lN5h/S9A+NXxv78+fNEze9iOqMVSf15ghR/xTNi0iE
3I/DIf1nasensoubpah1EoTX8Uj+HQdZWFYu5JkXPoKTdT4PLwZbaJOIFGyG2SOx
mK+y2DHQPxY60WHKOdrQ4+IfuwyuMHda3/76welxOa9Hn0s59I0QZBQJLqpAUgUc
RYPphrDINx3rpN61DFkj1T68qZho5e6D87JR6VjrvDa886m8uqJGWvzLrKjxM2HO
e51L2QjQE41z+z9TkgdLpcQ1FZD+UCPKDN8BQFzWAxzNhA+XVtzLbO9lmoeljmvK
ZMlsGQNty60Hf1WaE8V+cRB1Hd4aGTiR3ea4EihRSiK5A60juD/s86vxZkErIsrM
+nMOFP7r2IjKtTxckRZAp3Nr6MGZOgokm1iCNuoZfcGa5rCXecnsF2wU7D+QGwuN
YzpP2c1sPAF0uQAtr3MhNNWiL9T9vZ52dT2ud74Bg0Lo1YmqZDcQzm1ennoAngmW
4aQCum2HCeP/yID2YI1GuLQFNVKVMIIlWN236RXS/iShxZfenM3+p4b2iGCUJfg4
IB5TWIfk7SVGlbMXDlYOWP4D2zoLKf4SJgR74ClybHHbgq9vWe3yWQzxNBZJ7kH5
/fBOQkxAyJxzocaOecQqVBLR6+g55WJ4/l6Xfcoz1ToED9AclYmGsjmMx/kB3fkO
NSL33O/ydHNSysq5Z0cWn/7KomY8Fp4HknH8UpNyfCLjD2zcGO+xCs8U0swEYZ0w
okgz48A3vGWrbKB2ars4ECla4RWuo3ucqe0uloy4L6cuxAlPwNAug/Kt53mYfBCQ
Y7C09No2moQBF41g3qWQ035uuUhA1ThjwvWAzX7kACHYLH2q/kU2I3ZLbMXr1tkZ
M7kXJURNn4bvnuFKcU9OSKaaZs8uoJLXcfRP+Gddhw60ScjNvnr31LhaJDrv6Wb6
ybPBjOXOz3xQqZNI/l8gCEhBstCKcWu8hPS+CbT3Sv6m17qiicw0yOtcw5DHox6h
aoYUyUAqWbLWu+gca+YsQBsga6AMG+kLLZvVLSOUMEaqcurzmWkv8fsIEnfA/LhH
SOION7YyjNpNoQW9TCIw8ZpRuWhJ0d3Dd65YDq5FTaLL/E+e7mTpHUH8z57Xm8Zz
6T7NGjT73TmpUAJVApJuqg7sf7JPbXpZLp0CDYeIox7aXFdbFxJw5/4jC/2t4laI
KMgoV9H0J1SAnFUeX7POw6IvMfJcO1GYaq4IDQCm/i0XkOFJuPpk3AdpSAfh7D9r
hn1ur+PLdrmPRz3T6v6aDAq9yK1HLxmruN0MBttnT0ejkIjDJVNMtVzv6N0vPLwx
xnRWBZMYT3futmTRuPeT4enshLPRiWNoNkPZGm9TLmsDtWF/oxK6GdXqnClyOVYc
YS79WKbKD2MYClJz/ao8jIPM8V/d4I2+yGgJcnNpQoqkx+ByxrBe4RK8Eu/szyLA
kioaTHknG1EbiMg0Z2inBYl9RiWGNTu3SVTCdLWwaq3dBV3b9rbp1nO6tF5hRcpP
zzcwcxPjgCBPlMiDS2u8igqbR8PknkHzK9DIjES5W9tGlvf58XZbJNxXQAMVLv9k
X0DWtSCXb2ZJAO1sjV/TVwZcooyOSqT7Hbcts76FL4YmtoLqY3naxRRsG/AZEWRP
y7CUduR0cHItOde33So3XVA5hDOLJByVA5i7IHEjteB7STNzuuvi9Pbb5YnnrCZU
c4eYjyvP+ducE7yXjXVFi+Nzptuc7QvxeT6jB4Hja6AMPz3SebJPXqhbLrU7/j86
GEYhf6ybnrb0A3+wzS27pHoZWzMtrVsaE7XKI4NmpS+KfYNA6nnTslUeV6vXFykZ
wNlozz1RFgSYmW3cILs75ccN59T3fA39hCZdHu5RTXn+RhteoavaVepKqyyP5Aug
Nrd/I/kB4hVOQyedlGwiQPo4/0VOQ3z782++6/SMuGHmpYPObbu0DyoUFd0z5YWO
xxU8I6uz7M0b/iWOwV0/t0SPSj2QLCPP9/0yRikUJxsq3mbu2x1omnB/Yx4ws7q2
WdwP0I6HPd0c/YJNRI15GmJ8/aLF0+z6d45mlRB9e2z374uUoUMAZbjBj5BJFnkB
HoZznb0s7+5hG0xtVNA2akcQUZuGYOww7HCkO7qDAijBgNUcSTU6Xw/9GYKidxHE
sWi5mzwqZeAEryO+zS4046+uI4U4oCsx50TVcuHpat/RGARuhG91TcTcc/2YGe2E
gOV2pty7X0UvA2oWbNfwUvm8SGg3kbJu3aevwkT5oaazC4llbl17PD4KEa4wFX5P
uhFftUY1REDRezo8Zidd5y75QyRPDaFDh+kShmj0kjAOvO+3qp4k6/TRR8OPIO/u
uMNVWU7a/bLjFiuSd7x8ZtXw9KZVPG+M0u4GC1vOeVRWvSNQxE8M6BXEOiI8HP7p
HX4bjWHKbgpvHL/wsARH0+1+yN0jZwe9cRs2m0QWykmf2++hnFfqi3dgIi/GsuzY
wVss2NoZAHh2tjLIa/xOMVsnCx0TRRYarEtt6rkWqId0BolzXVwR1UaQzMRMcKqj
+/rwi3UQP8LYX07fChAaY3AfoRRxIxQKnk4LrfECs3t486SxAJQ49bQTl9KxPorm
s2SQ9qHSkPuQBF67mTwJHL7wmPQ7HZtbWBMXpmmQ5+s1An15VUSBZSPVDndpR3OS
mArkHs2RZuv7O9QpTB2J/47wt8wDKBUgLfVsPjm1r0LHBKQEMy97yyZWiAOdxoo2
3XGoTscEAnRmjg1pU90ypns7BNbrjl+fu1QMImVDsK5eH+O0ObrAEkS1LasQ3JFE
RqdZfc4Ufvgx6q/nmT8yFcDlBmaZPI1JBk4pzf1VehN5vowaSoGLgyDOXzK2YyuP
4Wjv0SI2n108AbxBBlAVG1N339ZDHhi4YSsfGqaN0qCl/oiYcns/yYrB3CR31I1q
DfGxBDniwydmetncLF4DLBtaR8PIogkswC1ayHiAnl12EJl7Tbvq0PHgIJTIWm9R
RuufNsUmqF+TijkDkylrHN0aG8jk8a4RcNHvaBkLOf6srK8s7GOecYeXM2TiJX3I
vVo1xc8ZqHsiMw9kwoij1hsXnOxQQ76h2DqUvYKRYwQWSrZZGYdPsJVRd3m3N3Vk
ov7qxdu7Hg1Exxvke8+CROh6832nEDAVWeJr3kd2JcN0JHME5mmNeLBt8KTTEesx
WHy46Mf2vbpwx3mDkRCzvmIBpD/Woc1wmRGstJIs3hUoSb/jRQIhA3ZWcOEHtErZ
zYgs/pYZAcA1BEHbuGA13i/NdAjlJ/w/Hk7Ze3J378JUkm6zferIqsJPI+9q61VR
AI65lyRZ969NBBL6pQ3xrhYfTVMVG5K9iEVnpOM3oYHYy0KA201AoxtpzeoA8DWN
S2qUVac1VNR+64bkhr3/dz73Bu8sRTp1oI9zOqAZ9O3ciIB1h8v4xABkwGNkBSpD
AREqWNae6BOra3uSU0HcoZYYWw9tpN5ziiOkoe6l6bPjJInD/FAqUZ8UVuurSYJF
+/4ehVyd9k1olLT8mLAIuXptUlTSEuAL2ixPwAx4fmcFvoLTtMhOTX+gi+s2Ch2Q
srhgfF/RQIkua88FbMeb83x76vBDxYTHa+wMymwFc+U3tszwc8LKC13RB34aaFv3
Mc5b886wiJ5oIm1Q1ZduZdW6vxdE8VZWR960R9TuXDqTV/Gi5QmIycZHm6bTRD15
ubyGgyVm6sr89cr7rnIW2qRDWJkcSjtDNppS2JsrVDLLorPave0AUgFllnShB91n
fWYLRGiKWSsss33hgGdl1CNPk8+wSS2wb8YGkGTED4EONnGtR5sW2xck2R4ZpjBA
6Tem5l1L1lYlNOh8ivKQhMX8weV/aeXcapEMsqwcFTM7wkg/JHrIPi3OdrqBs0Z1
NO9NeZfSGsJ++bfHjdbe72iVUCCN+mFWUxsIxLehUnjn6NyISoF9BtPXfbIqF7yn
Ye4ROIHKGc5X/2Z5r3llH0i6zWLB98l99QhXAH0C+SgxbjakvM2FcI/xSS420mbR
/zHcQcZqAVt4m6DQRcjQArf0G3ARiZYgWyM0ls3jj/mAYXcoqeIkv43CICsdB/VB
7tWTr4ur2l7lj41oTV0xIsEKapeFXq2VTLmQXiWcdDhj2CcC2IJ/R0/ZFBHUFYRE
JIvy7IP3B6SB0nc6u85zawouT7W/N3l9sxKuiydAmVwsZy484RhEBcIDDtJS4p1P
ye+ncZ9VRjgCm5UJ9jUd4BTBpMoELWVmuUdooh1jDzqHq+bDV/4tnAXnrWqxNLiO
K8ouLGWyayzL2A7bPTa4jZnGzx8nhYGWpKxCHADz9D4LEOPqG40c8pHuZ4/V0Bc0
1/RqDTjx+783dCkYSwLbB9MESUsuuJ2WMVueouBbGY8pPHAvpP/VnHH+Ify/KKvX
BXwZjUOxGouifKYkF/hzCIfvJWNzzXPI2x3VbrwJDQQXtUhJBQM5QCH4ZNODmZuu
a2MZTnx1lXHDNmRv3jr2LkYFfua6c+42KRgntY7n47pH60BCAbtlDu+N+jvW3I61
D/moPQgT4eoWZqPo31yFcaUYE3c83sT9UN61GrdCzJmeKr4UJFnKQVWWTVeDYiwT
D5tZoAjbqpX+QpAvfk3HXvZ1cbFnBffVvn13i77mkE35Z6podyGz0S6KG8nXn/gl
MFfjed2zBT9okj+tcPgWUNWRW7MOdUzqLtjqxwf/xcXyOGwk8jqgB/0++MPzCYDD
FMlsEDfz8WC5QBm1vNorbJ3PKZPcIY344Mx45lLphfaOfkmkeUcY5EHsjHtAlTTJ
3h0dnkgslavHWu2rhmAf3lgfisOjLd3w4RvuCnbOHrXhN28foVTfjQSuMG7Z20zP
Cj9fd+tJ/t/EXhDrO0Y0I9IisZG5gsYw6UKgHrTTb9+GrGh1u+/uAP37xafgx6z3
fdSK7qH6HykIn1fgO0Gru5Xth4OEXxtGGr6xS+grTJAYbXiLaGdhl2d/50uh37Q3
8v2dqJqNrPpru2C/yk8J8yeqWXaomtRytQhLkbAgTdSid7eP0chH9eSmYcbAP3lL
AYv9DnQXSrys6SVElP2FzuPeGD15cALckNqLGFgGfRgRTgxIlKp5xmPrtJO2AxKs
s7huIjAt3fyOIX06dnppyYfWBLCtl7xA5kWaf4jobYQhv+GcBuPNPVH5BpfObRkS
t2tRgSDQMYCulwxxZuvGpPa0m0mV/ItHkJUQF8UJwT8DWWLq0HX0ojmJiUcEWJ7t
PMebcwSmhy96VpIuF+nNXtCInvCvKQzl/3A0WCzeb5fqyRB18mwV6wUa2K845Yp/
5nNYMxqvPt5d9TmcMJwbWNtj7YGAmvZKYUIco9OThp20ZsG3bs21CGsX2QFfXlbw
F0Rc1+5X4rFMHsn4/hSaLb+kFokv2khXYt8TU6V/2Gyq4gCQIY2P+o36w3pPjrj9
1QKX5IzZ112k0GITtq5uHt2m4PXumnYNl85gjRnIXdtDCGEKKZBQH2CGkUGTx6uE
u/4bDDbI9HNpTMYYxOr5+J3R6wBHEbWALW34FiiSevUkrhyA2w0AehNXuVlCSICA
O6Cz+XYPNVSDFlDXD/feUQc7krg798St7fHkXHqConr+B7wfmoOZJBnw1MMpj76M
HBhCchKUWdGmCty1HRLNbyNZNfafdqsJ6UlyRi5Ssy46TFzaCoMtam8U+AKCBGAw
3LX8D3cCX7D9mtngn9CGaxDFq3TGn5vZSKZ/6TlSXWfoAk+NMZVFnCUxTLfMO0ZD
O5HWX+2Ij7hySVJBdgWG2p6rF9BjGVqLtduj15Mv8lvDYeODjP2lomLCNZPjV1OD
aTY2fHwaPGI4Re8BT2AaySuwgLdrJ7bCS4AEUjoQOt9xetnFFO+tWRi07d8akDl5
u28L27F3RrHQajZHkGROIDSHDrVg9GA1xKub2QQnXRDxj8T2PiVzqHZR9wWa3B58
IZzTWRLIZjfpR3tmY8mTbRXsSMbOikgEouQDN+u7se0OUMEH2WnCAfsvnFLC+ztZ
hUHimk3Gu60EqlUkKQYXQZ0ChzBRWrIYWpMBSCmPD+F5+180a8gKzGrAOvWv/G3n
K8q7AQVQFHeOQ8KV6wkMhiOTfnkVcdbxhjFUaYMJCKJo5meVB+bHtQIkN7S9Fprq
WbApugGPYIVQHaBdbwbC35wFIEVMUhmlA/iUnm/6cpB9WIsybiEebCVl3+pCpM76
aQxWmQJrYGHdzjkyqgXwVK/mx35uGtOUDUQRLhFqF7ybazuPE9iOxlFCqQ+HZjOi
1uv0uwG5AWHQI2YIM11d45mi6kfcpYqKf86XpJjpndJe+B2L0jVtVkSvuzjns9ov
ll6O33MU6fkE3G2Y8m5sc5wyleiqnpkoY0vRbj/KMgpwnq4bZl8PyiCPHWmcG0q+
282EDCAMMslnOutazfcnU0pqodfcTktJN1m0oI7FE35lYqo/xfZ/393HGYAPfXKO
42Ip/34uTNQBipxiONr4g053vqe3cfvDh0nMGWofw9eh9mb4ysFJ0JGTlNgeazJd
87S1mOrKfsfJAbs/+lAqiChtQ0cV2+oJIrXCvmCR8Brxo38GZ8AEsMQFPssX3oIB
lhXfTHZulViXSWTKYyJcHIzH8E1vEq9/rZAyD9kdgslRrD/k+p0O7KJbbSq64EoJ
zWFtTs23xs/8wBVr9r0u+PjDol0PlJfw3hJ8ulsMu9m+rMTEzQOZ5m49i3Bj1dnr
q2o3fx2jISS13p+0QpNDKZ1GD1jbBdTm2F3w8FboQoYTaoKIOAwZv6JwaOTjGkzh
W4Gz26xo65YfsAqUZFGL+cB4Wqapbq30XA1X1w4U504BgCqAlDTCXd6MpW97hK5s
lM/GLRFXhA34Ty1rp0m+HC1Reu5BTBCIBfSJX32E1pbouUbfxtb+/aKs99EdSjLP
Tfuu6kVGXFEqrXzYtKobsLxaqI1Daf51OOa67UIf+RXjtBXrC3KD0N+9lg+R1s6p
OaiMGR0/MWkkoq6po2GQzIMrbqEtipCbn6mKyXVTcSAq9OzjlCIJXqK2HkJdTBtu
Di0GUqbYLQpY1jVgewg1lyD4x94PQct8i3CcPkWAo0vr9WqqPqOeyas8oPl/Jn3b
GPjk1rTu07vA2bqxPwrtIke7oyaYZMAqs2lQL3/5tpq5gnk9u8fSqB4BPly0+Wlz
C+iCNEDZ54E6GQN2c2+FVxcml3cUXu1eqRuXJdQbO+dCVEc9YUUela6eJklaNKap
iOW9eCnHk3temrWC8lm0CXdhsESqRT7TfnDXgamFAfAKKy4arFFVfp3OlTBboSeP
L78saOA8/5EW7rk75xjaPK1BSEY/XsXD0gKYrycDBHojKDv0ETOjRuITxBJWPJPP
RefGGVg86rK7yk8xU7ofoGroaiH6xyobr83nQ8x16c+OZbwBpuyMsKh22H6Se3+N
raypvfjRU7yJsHxsQbbtlVNOllRC9eeF1XI8bRQxnG3AB24ovyQOlUFXj9smALF+
JocsbzBTTBloktOrE59aCF6GNE53VcGff4TL5upSCNmtMO8vfappQHNuWIF+2WPJ
ps2Deckw6CwXveOnCoDrMV0zfWDPIMFYl/sDMBNbNGxHCz7lS6pSSp0mFsP6fg0X
+6Lp0gd+/+H56ooNvo4+5pKz+BycERZV2kYNq/u2vqeUkUatR2VMSmXv+nfmuS33
6SJ/sDVR4140l3JwJUI98sd3m17Uez4ycR70nS4a4qhhT+kbasdicFvujzmhE0H0
lBqEDP8UTena32rXY1t72MkGpnjZTSTwzuwR6S8QH90Blbm3yY6Ob48CbEKqByyU
OuYmYYQ/DGfVXUfQ82ONNElybkkAXqQLFY9Yhw4q0IazV5C5WPHvgfQ7CPPDZSA+
umNk61qI/zQQv768Q9vKmPXPxMJYGNBZaF0XFqo2BergIoAe/C+Ery4a+GnI61UP
35UAUHUK9Me/o5i0QNIWnjhm8WOK1MaCa4AJ0/KzJYJQWenoDVn94CTi2r4xtdI0
haKYp7ajm8TWnuY90hRIzi6N4NRa1M0gGwoKIwxHCtdUe/MtTlqFHtv8zE/AXnLL
kpqXlV6w5kVUjHgUWLzIOQTs8k9RUYY5hOYmGrBhfy5966Vj1Z4a/jTy7p8HwTxK
ZPIjeEw0n0ToozXL7HrcBVHKTFy4te1tXqnxNePuexjYnfVRZV9ndavBY9JbM12I
EsgDU9REtdZ+ddcJ/Fi6M2CTtuXQ3WfjMonIudnbMRDxYcxtD3gG7b649zgUq2Bo
AZ/ZidEi58YwaeRI7pLJV5/FUyRozA+l2ajIWf5xWdl4xM0k3D+3l0SLRwc+5RGb
fxxCW+Lai0L/b3VuZA2hp8CNX2R++RqNCjBHolF/lngQLMh8ZhJ+h7+bGJJOEp4F
j+08Efo018Bnyo+M3fEPbx7I1sXJRT+GXWdrr1hraRsG6no90I7SCOz+V1dQfpsz
3yxwCQEChb/MC2LNQ57NUYKyGryPTzM0gAATKyzIHeNN3cd6mpdiyDzdOb3p7XEC
WhUBCQ4dB/Zo/tLVSdCHrbzRi2IUcEfs1HrgE1CrOuTvuKEvrTrzBvJBK39ewB3W
gaKGpwqid25lZmeTE5bC17FIbLx/nJ29ey2wFgTrjgSl3psDqYH97Yo2puZrY5pU
nqMJpBfr2PVwPfvoQmn0Lc0xl1uTRwmPra/JJjMJn6Pfg+aTiCdkfTrGEFFbL64T
aLgizjh0tcf0HYGp8nvbACGcPNFXFzTknVa+abHlzR+KD+cX3LZVXbVpGegaAevx
JXv3sHC04Bfl6HxyqC6EoV6e0eTszhWiqZn5bS7f+TjbQOPyq5jBaNtKQRLbeHEW
8mKHqJ/8cHd19tEDpqJzFn4SkQAEnp9CDCWphyCmYwUYEiu6xhkJfqJctul3ljBo
Mx4DW06ELoFztRdimIDrp4UFnT3mjpP34BvEqA0gn3TpP9ty8w7ptRnnRqhqqiiw
6lciazZbd3jMZbFuv4HQF5ch66kCAnc8w6l16fFBG8FWF9rEOSVt8EIgIeksZgJa
wsL57UEo7u3RgaYH7oMdxtAKMoNQECDsMAoZ/4DY6NUUyohCSrqgvw7ngduGzR8V
MmEhWoSCEbYU1n9hoxBfxi7oaAqX/k/rt3/o+yKslBBR4KJaDzmCmqkK11OonY4w
2B01KqFUUbGjSpnDRldI2BAiWlXbLzC0oi8Z7HchFiIdZLsQhrpZmU/+3cntx22K
XmTgtX1R3SzkWvxa7RAsM2Uo0vXxoAkRAwQpNisca4sayWnzg04kdJUNSWlrTzBU
WVUzEbjMviY89l6KvJav5oOQAOSgIJIK43rKu3kHnyfvpp30lz5sGZFeeWY97Tne
KhemWtIbupaBo7vLdXsNOVEMhwXYgRM8LPs+Qr9Pqe8HT+RSJSF5eSAWV1LZkT/X
t/G78+Qy5sUW5oVKOJZsFvY5XFVGfttG9PS4re8pseahFGRhucJW4TS8/zjLRzbZ
NaE9cw93kKVqDhNNzXJzuz0Po4Ci5UXa5fXXiVjl9g3z7aO+DZmc3uzB25eoLSIs
iKDh8WeBTUSJrASQypVu61GgY8jYaurAmSOzUay/VH9loK8Lb647nKe+guAAlIGd
pXuHo0ehkVrCw0kDnnrGb5NnTf3Hiy4zM6hvtKLV76DEEOiJqNvMXopUbz1Gl1Xk
6oOQXVAwaX7ypdWOwHtiz1ANGyZBxxgIO61z7SIm9csXiTXSA2G/0Ouw3ZOXwAJ/
2RQ+b4SkbjBpyqD9iX6/iyS8LjpOCuggbAuMACFuACl2/ZToqqatcPK6ejm5AqkA
2dJUYyA+MYa3720V8ElekuRSenKiV54WDxszEZkUIWXiHHngu9DmAFnFR0ebVcW1
bS8K1+QBvq2NBrEtnIoG51n9OClKPG/Fptrztz8NRkJWoWj9FubZBTyyLoUpQfVl
V9VsnuRVEcGvalgyAJ+kl53BDjxG52NLENmB9FoxBFnQbER9nqaJPN7gfkk7iosn
E+SB8pPjWpS5UDACqB/aX9mSSqzJ6NVN/h/+EsL4HARbyaQMj/sRh3lUv7yE2guy
pHl6UH3LRenIyDpbGk+uAaeW5uYUx6hjSH4hlJfYCv0Sql9VaaalMXaObO9caQk9
Pj746qux2NVvC1q7q6pun5TBEJeqM5oGDgbmWVrrW+mBKoQn5S+B0AmhBFY+w9ep
qqmexYsk3XAsTWWIw5iDGtnWSafzGa8EbxUEqthgYjwwg7awPm5isxODLzi3WM8k
n1He6Hv70zGt3h0IfSktxlG8oqzuhMB4ah1DZs+G4IQNnosD+KVAwXohQuvdv15T
dyOd+AYK2Wgc5uHY6QmemX9L4sWquE0vdAuUKoiNHwkwHW4koM28dY2Hu7gsGt9s
p4IthJDA35w5Zl6uW8uehX7SaqSaqj1qy0FcdK8f+2zsCA25oYUhWs4xXMWGpVF1
CvRvMVpVRtpPEV496UMfk0VC78jAgIK+XngTf2XvESbEbh+F0O2IFkVzSNEs4kkh
7H9t88GQpRYxkFbIq0vvZCMUxrwT7O7Ru7CavyCeBGsmb9jrhgRWNPsW9thcc7Xz
Vb0CMxIL1wjzjb0DsYmJFGa/iV5hO0gnpzV2odzEuXAO8cfrQdhDF53ovvU578Gt
tFK3omnNByvl2qLcMYA7BW/CCLf2QwlI/4enuTZaUxSYWUI4UWin0+HdbJqTR2u6
xzguDp1XJ2oXVUN+gNnGtqyAk0ZPw8ex81gMlEro5iogNFF7ZFpY6Q5b4jGLe6lb
kqa+HByYbtIkvVefnE3y6MhHYBBsApCYZZHdMjy00MvIDJIaBtOPySPxWji38SNq
XUWrtRjNY8SyJbJFBb+oKpUfOdPt9k92hhYpbBDrVYCyqMP1UUdHWZbqJi3B54HN
dA3u5gI42Kwvo5WINcnEwzBpR+6IAow2SKXfYfY+R1/DlwJ//qcFsf25drJRXb48
LmueJV3LOXGasX6/kueivN52f01iyvauoDqlsULiy/QTZ+En0LsYYOwQEJIbXasG
52BuDP8pwwxeTeFXlbRR3gNMqjgKlLp2UXk5de3LQLFRofRuJGyIU4SP04z/fT/B
f44uprZqRjMmMb+w0BDK5KrQjQ262eiGEEJ6zPPIQ280P+cDibAs54pWMosN4kyB
HshMZSDixn4ZCEdqBxh47808vrLSTu4FXYTKzLngJ8Zo0VIy/n+5UGliELdzrRDz
HSr/9NdoLVAvCxJuKRK+GTE5M90NofaxD4BNgcDrqstnEopeziNw4DxLu0jF7dtS
NNP77DXhPNoNY4EwGPMi0dvhYa83hLCPI5wuiESZpquh8yDBGnTtQH65sTBjDpdZ
TOUsrl06I/hM1H3MWzebOf4M09GAg0ps946Qa47lSkKQTDbWewIPtIAl3LN6GV9z
ov/pSOV/n04EM9ZINHUYvKd0KtKJl+BF0tfGn+qq9HmiLw8KdT7VgeAlFlOyDoGu
xH+4LtdxocKEgumyp517PCETTiBF2qnYtGuqMPzDqOHr12DyGyJqIlzKT4jQQBFZ
erYb4MCrjMPMpLb1qj7j8mR5KtTxSmkoClNz53gp6Ml+noHdgGV0RqCuIhCwLvK/
gi9fSUvVAZ8sRGtgPXzk6CKnRw8u6szI7YarLNEQwHGHUZ4ekQ2aQNfwXLaz91gj
UTkFIzCunjiYzNvXxVWWdT4zbrzXMiXtmNwtmNtnZkqEX8zBFFA/xvHTkIlDZup4
QdwCrurVvfx0SuLJGIq60KlUL6FAeFr8h7Uw6B/UIqlBIiUTr31eO8msfm7Vb59N
KftysNLWmRsT2MpfN6Zoo/KTVQw3BdSroLu1pbbhqsYpGJnXFIoYciMM3NdmT3w9
NeRGhE61gSJ13FWaddw0LpagVDJYYrVV37KTHdUpJ52naz7iQvY2zlDChItPxzlZ
u2+RjLQt5Dyc2Pj/WMq4aV3aiVjv/3+UlaFjVmPa9hrqDct0HRC2X/9/aKpsxaLC
KCzAf5SL2QVqu4ajluDf3e/fhNi/lI6qHtgv9tZKmm0qIDeSfctB4lkr9eDtevZh
LcK1dDM9M7wunhSg4biFhtJPfe98AiIAdPmtyKO5rXoVMkmqmBfkTd0pMktVoSOp
vbaYOHBZcbONkM8I34jn9zovwzCk+laFTIzimS9AYgmGLtkfyrNn3zlI86hOoK6O
etFaPiCIz5XliWovDgQpFcGZHh4pjyd47DKanOVlhk3wWghBwIoQV0ypS9RVw3QI
41xKK84MBI5TNAFKmBzQ7kEKl9NOHF+vHD19QtNx2mdvFuKQEEdZdQZMG8teqSw6
Am1PNE1VNpCV6tXmIgyNUWVPHEosd6QXUgVsyZwkgHYN3qB1YGIDTzjb3OiOWUsm
0k01sjYKT5E8dpSJqg9wQxJgpqEWOrPUQt6AXuie2bLJWAkHMbVXSZY8nbtkN2Em
7AUTN3TaA0TwaMM8ELpRMvXSDRSOb400dGUIAOLzmw61ASgxbFhlOru6Q9Eox5UB
OHhqq7C9YFzoI3Oe1KsjIHu/mikqKGVQIJeNvoUVWr/boCxusUU9mEJOZPG8jTi2
lKdfnFie9ysi9zyvKZn5JuiVfxENoqZtRtIG56ypErIBSSuSZpBo1VPR/AWNZcaH
X23VkwMp4vEnwiOEfd7sl4bTKQ6zwR1us6gxbGlOPW1ZmreL/37dnVtBqo/JQQg/
WA9+F7+K6MdE7VbtG9SSpcWA5WorRZWd6wZrKE/aVlTzKfflkc98/vVUZjIDV4pS
BZ2tqKL32QWlKC0FkHqHFoW3BPR7hrMv0ehEy4VkPPDCegGEBoTS4nwq8PR1530Y
m2Sc62ZU7r28vBn3Dl6cLkgZLvPWIQwZKo2m0RL2TVopqFb0Xba5ih+TlETbngkk
IEpElMB1g69DRZl8PotQ68wYSYNnfXSKHx3IPJjPe2VmgRzMa0yo87B3dkEptEj2
kh3Oc3rt0a06/gmFC5p4n6nv+ttaj8y3feYQyegVDnVHxD6hI8hS7EYVlFboernF
oOzt/6RtmPLTemyA/g1P2DGifszqHHyIzC9fRKqh6VtjWkCaCIkpc9AvXOTIoe7g
rfRWCRRORbh87LA8ECDXdu/t1CBTBSGWxLLVLEsOVLsRQkvIQGpbTKHmwTVWK+/0
SNAKnxJ0iM0THo4bZ+CGMR5pJyDKradrOtmWDIIt/ZQlQ7nw5rlNJn5n15M7+OLD
JCvUFXFxldi7aS7RaZGd1QEm0YDs5viB7g/POIknQjkKXPCs5ydsku2UcjA+78Bc
dQUE9ep4/FMUNl/wGworcUAW3NisqXJBxuzfuIL52ub5lI1uBnFxa/mWDjdzQN9z
nVMiA5/OoYsjT2L3hCDYafVaydPeIO3ePwZL8cZNWqJAdGOMc2NGM4FmEGOHZGr3
Tv+flwmQAhA0LzSyTJ/5xqfyc0YF+Dbv8k6RPKcVn/lgndBw6ubZSGcl2CUPM+b2
/5nOHgHhm5/A38PQDkMBy79ijrCIz0Pgx9Je7uj2Zcd6qWANWHFTV2NH/58leCcP
7UNzLrl+0WwkTSbCvnUJw2s1mUYVMVkeJzO9Wf83VlRBMc5l+QuK4+UOvMdRs0qV
9xLkbDC2YSW6Erio3XZ6eukTXl1ZiSwABB8MnkhOJ4FYjqD3kME4IlIQ55hqL8Cj
0JGHsL2FrihOsD7pO9xX6VnH+5z5w1Jh7fGMMWeGTzFAGD64dGxbgh758SPuZ8/J
rL8ykvi9uRrfJSf7mYwzBEuzowPc+RZGIhZhU3dWDc27O4fXPF5erDPDyhNhnD8s
n1Mv/nf1BKbdxSNbjc+svJ3iRNhQg4IBIBd+1QR2IZ/Z4UUjDYZBUfcpHCJeieL0
dOitmcdof60OGPsmqIzKTx4Eeuj7gUlZuuULx9Vx9o33YE5ej2oNGbD1CQ7jbnfw
mczg28EvW7B5rxR9U/sk5LVg0L7actO7jxee51uWk+iax96k49qNxK0eNY7x0JvH
8kKzc2k8lCauYynaRCvCVMbrxZhZt732rSYzAyCiy+I/v1fzT2VD5gSuDLKD0KaM
bNk7GfMvoUfz9OrYwdLIVFlwENSeVB7Xk/dgTZ+R/Zc/dpkx04YdD+DKlXn2jwqZ
cY25u3Ug9J4KmlxfF1GK0J2OTOwsxLNyWwK3NABq6ywtku2CEUMjFVSNmrJnPiMc
z1oTENb3VO5TFTvdzveUfv4jDjXWiZkGu/Fd4/be21yozlsec4oNyEclSKUPd8Rb
F+vA/2QIYjusdf3SLIPXBu05c4ovZaxnOBZEnuGD9SwKS9wqHODofzgyd5ZT4Dms
6RpoWZivPZnyU7IQJkrdO3y/f6UJ73keKRlD1W38oaXKz/CidF3taCAR3ToUOudk
rAJ+rxQME7nwhOEL/8pXRso9Y7dSptpi6hfFQjriOrKrEpVfH3exmJL4X2SLH5Op
+rKW0DpKcqA5EIqxOXkhbEWSiU2w8ylKq1owlbpDGKbRPa6AcDXCs4YWKc4RK0fk
a5CRTceB6pBpQis7Zy8Am9Iu7wdMgZF+fpO3OmImbUTU+rxFNw/o+Gbfi8hoQj4x
r6C4bYzC1jHkFYIma9ChhWZRV7+cDYeHnveA6ZNHJTl4xFpk6/vH+SHe/xRnvJ+b
yju2omPXjIDsBj6qPmypQbH8bARW+Q+9hUD79v4KLKEar9WsJqWQJ05UIx5vyApG
3Xblmc/FpOm9fDg5tPB6ERaKkrDcWjdIxjMsc8Wdq7QHKD3fpoiojTjd0zacLNJP
Yu97bea3EsgjGcaVHISZOaPhrM5gQbazHu9bJJ51Rj3a9nftgnDgRIY0G32En64p
6aM1gbB7ipucaPO4HZhkmRTTLGKtyzn3naxJD9xrfN5xv+u1GgqmA9h4zcacrutH
fVCCEzkmnqrt17hCMgtd2mjvbaBNUp4caJ4VqweQXHIzjiPXlV9WJaO8laLp96IW
ocSHVh4I4/ZlM8X7Wn+p5r++qKNPjQ7ApN+dkQzoivz/bISnt3k1sbca/sN/7SQp
X0QPqQYHml7650SyFlIzAs3DM+VGJuR3Xyw+Zo7YGTRF7SBQwWB4nvx0DPNRgZQ9
h2TPYUaYDEaxjfwagbfq5XvawI8epOB7Gmf0BG8QKKJVIh2aP3CdDqCztgB5ze1b
lg37x3n6BBi+0rtHzPheKXklPgnMnAk9HnIJmfxFxFiNqUWn1mhsjUZDe5OpeVxY
F7S7LEoZoB78sgnQxAm3HemLS50AbTC7YIw4VDWav+tnVHD+4pIoNaLCB2TcNqhh
GB5zpQpLQXuUdDezhPxsxyjPQ49Iw15iJ7SS19GNYEA9+kdY+cMRVfbQUtrgBV7r
GgJkvuhprFlJ3Hy8SIlM63js/BmxT+fFHBuSNoQfn1aAmE8GwvBvrrbrmeV8SDK6
bJPVYVHkapGjouw3GJDZ9yNnc9SnzU0CnYGtB4Zdpp+qHAsvgpksMW33mNlGb7mN
TDGZBDZN9EZLFbbrmgIqj9ebsnNbMpsk1xsny4KImbMmvT9USJ8Pn4fwBX6TD+1o
9GB+vpm7xxD4Ls2WYTOFejJC2vLACIaxI07Sx+LfOLFacsuK+grbUjk84MdBNlDu
Lhw1zVam5Pc6kJzbShHfJu1bcz+/sicdDH6bKk8mgAUYvj4L174Icq8rA7h3+jp6
QgXHdWZgBqdo5Jw4ygYd5jwN6Mh88D5Fzkl/az/GynLMibguotJMOPh8JzrX1/+O
wINUvDgZBGOVWaW2hHQBAnlNzZJvHSXFn4dhkgOMvLF6MeE7vDG/65OxuCg8HZJI
awYa3zu1ZLZG59sS/dz5WyO6i38lFdVh7ErJaQfWejU/xz77JOHzH6xfTpO2lHZy
+HJQM/V8gA0Du4enO2izAJFFYqAGVbnlQzl4NvW4H3RMDBxaaoex9+PNJ6YyfC2G
ttQrjotb52sDkGco53gWLXRJGDr8pj03J17FooPlcZL9QM93YiAKiH4zVs5jmwDu
lXGqBj57p0xTF6nqGKWzB5USdIBqOSwD4LT7aT0Ht+MvXAcZhu1d3Ijg12Ux718g
c3EgPk5MRJtkkXD0joAVuGpE2b5AKpbuLUhrFJK+wePLJy/nHSk95Wso883xRKNl
UB83rr30d/V6+PyATIGpr2Rp56EZdpBfoG0ElJqL0Hh9RNMH3hFPCdSALTeLcrIm
OQFuL5rlngyV2FQgggO/aWp1hehgco4pB4PO0H3Iw/WDU6VAEZN3kTv9EOUW089S
TfIIG6SPLlMKMM5q3fTW3u5bHk5+CGyxorBs3Ett2dd0eqrK6FbWJxNigPvqRvL8
5sEHdRWZeru7XqTYZ5oe1syNCSThBLL5dQ3t+Or2ybOeXWsTNIaNJGfIZFpLncLf
+hNeyh0oVOMMGXu5/VvrAMn2hE4l/1FGBMrYFu3WN69B5G0r7IGArvxq4O3yjU/V
U1jugi7BWqg88bRqXVDRS7szWMYFrmO+MOSKdv7ylhcve9b2HGlymu5G8b4N2gC3
T9hNIE4pi6MQFXjaFKriObVg7IK/eWtri68hjtfhFsgqCCY2GvVxUYRY079zGn2r
VTFMRzFbOL/XDdVVXyOsNd8HrwowrWZ9xHZggPmaTh9Nas6+XaSoBMxyMrHh4HqM
PudSJmRyzE7f7XX+SwVqNjFrG/gvFcyKbid9xpTjyIA26zMvoQj3QaKZP1eSZKsk
QBBl/5JWuKFh/OmKikeDp5bNosK9gL+8j9OzJigWbF1M1MY4XO2PB3ATrr8oUQcB
Yu8vMF+nThkbNTKbmlLZLwOfYE42QGhRD/JKPLsBSTw8dCc2HvaAKFtYHZTOnbIf
nS46HdnmXkfRZKXUBPRxUoqvk+H5RKOrxhy5l4h4Ype/GavX3qjtCWV0eKAOwdcP
egQE7ZhoKPGXUMz4+cCE7K7wcA2DQhq89qBqGW/V5CC5u2IKBd27dMu1mm6dWZc3
RMadQS+F+xjuvt+8XgBbYSxR8fIh/yi/29Xuc6+drTNdujEZcJvmek8B6NN3LS6G
Y3M5lYuqAiURYqMTXy05b7nxNiQlCZkBTITJV0fGP2uccMkuQR2hFokp32NL07wi
QFx/sq4TgzWlG6pxMrQR3VezG5/p40nBSsEkoUNJ5T0+g6yaNLGMiQRfqbamDFPN
g4Ni/czLt33+1hipzBxI0rSzs2MnBg0JXrRGRtjnW9t+XXfzSPypHUZs+Z7jW/75
h3h+Z+oy2MslZMDun0dYazkc/qXx6fsw4Aw/mTKt5GZkNtVX+O+nyo3Rkk5Mw0+I
nUgsWWTo1+52dWa1AcKjTQ1lOGhjMUzBTboeRVRanf/IsNfAmJDFa1fpR5lFtAhI
bbaY4LRuxnY+SWWbxuygnVFONWqYL6wfBRUgnpllw9DlIMYhu0I+Kq/yZ+lkbXDJ
JXypCV5XhuhxmO7VCSC2TnokaID4G2vhe+joKmL1bulmqGR2yqWPYfOYf6aVHmFw
sdzjb4/UAhkkayO75/TYRgmOUUX2XYOk3U86uEB50zIezCi/wZ+CI/Zq4gmOXzD/
VyI3TR1edVQ2ervMY4P+7ZucQLk8/pSCUlilv8fvFyvnBhgadWr2zQ8Qvfn5rS6M
tasRyQu5eicEqbxbm7THBGkFiXps4Lbc+F2s3ShcVPw9r/yn7eHweSFiC4GfN2BR
SIWhhWZZGXrCqlS70mV9N8dPg2+xVJ4jL+W1YOONHB54DMrscFsYELkjwYzaO18H
m0Po3OjCg0pddENGkbgsgX683/FUZjfm3nQn+ltnmJiQwF0MQ1fuFBWEs/aXzepG
cIdTZtE5kMhWnJqqHrlu7SsYCjeqlpcy6QFZnhSCVgpubE1VSvPekhUEm/nYVSvg
2KSoOPlDOfe8VHpM+GtgC8laNJ5aQbzRNflJBPoetHiCs2QfE7OegORwUmsvYnto
YsnNskmuVeThJ5AvGjh3ne+82U0YlSGvc6eiZkTHFdFfvL7YlI1nEnirTZHw7JcF
mDh1Infeticul7hGnwSrl+KBtxrhnAD9puw7oI3OdJKJREYpczb6ArqGe8HMdbo/
ayqQi91/rU8Hfrf5cacyZbS2GdeWnhbA0TlXrcK4Dn/4Yd2FbitowYayjTp7ZXf9
AQNmcEJPrxreJ5XqsRDhglLUeGIjre31eshJHeK6hJl4pYWB52M79dtinmwbutDv
MQ303w4a4B/DlnVaNQ1DkUe/UkT4sa0MWiFvprG2jTR6KYj//N+XIEt+Sj8eNIBJ
817twkQitepYNqBc9EZRVyCOrkD/1VcrsdQcNCeuVUrpJnVV6FRXRUtun+t/1XuI
dDQE8pvC1D6qUWRJP1OAhNsHeAKvXFTysv8igU2U56W1y5XGfK02CC6oVRyRIcQK
2mij2obB+USC04ZnxAFLWbGBZyLilTBSpmVFZnqjsXDX/kImUgzPPaarCeUQ5GdU
aM8X57vOTwhojDVw9k7dWRiLw9qFAK/qngzX4H2jExfQsMMhaqgXjZMie/rBhQHi
dfUJ4egOqbMXzSEJS9y1vg2G0GUhkxx20RArK2TsAnF5awazQ4bvzuGcRJAEhHWO
6kjT/0Uw4XO13HL3Ql4DqupCdl9qC4wqHllpj7OCmgVAUADhusykkO3vm9HQFjc8
5m2+l/HUdJwCUHF62asEE6DQ04MfuNfMfskl1lwAlecvuc7+CEPi0HB6f9r0t0kn
8xPMzzjVMyofQ/Q82iOQMo8RQtDQeZT+aKsWGxwjkjIRJLVjoqYx3bfsQ+4CsVLO
EA1aeWBpd20ohLA95jJ/j0QGeY6NCD0DahyjeexN26h+WPJZPrC8qBV+W4Y5j4FS
ylLEopbN0erV8QJXFaBSGvguIF4Suws68FO65sP9fpz8XGvFvCw6p6N2gdGzXTVF
9Sao75NSp8mf6AfTLSg60vhzUT6fWEgKp/iGPkUeaakTNJ327E5tsonnj9YrC8KJ
6esBj5+yZqstJA9dLZT34QydtwquqZ4V1LLT6b3vyHQ4lNKmgFYsuZ45Hv2KoaVB
C1bIS4gbQ3ROemZsfH3BSz6eRIwVWMiRdjcOTUNCdsb0vscxcahcDBqieRDrWVHX
XhlWwNlhMyzaCrzC0SjO6xXDv1aHtSCYqJIb4JzDwYlBfxWQhlGZyVWVQWTYlC1I
LPUzV8zSCoAnIwUr47utlH1r1aDHlVIwh2j7NfuBcAsanoI+bktXlICytDUVsaZq
TKhfSqfaJ4oHxl96hrAFTOH0TSCZmQUEmvl7gpdmgCcd4gO3P//+7eD0b8q9fe07
wxzFM9I3y7ZHOeUkqpMbO/Vftcpdde30u78FeTDJa5nazKNSawngXATOamHskami
JqStmtKLiuKomlTqz7sc62NqY6bUwkQamet5IicPSie9+UdAMcegfStfq9sunQdy
krrrTu1MjrpWQIsTRGDAd/qXbFrRCXYntIWsQn4SIIKhnkoS1tMl/YXL27kOMfUS
FnlkCan9UJ+sRLz7xikEzl86SyLOhIcJtBDrCrPwB0DeZIeazTpiPc7Ya7V7xJqB
opJ5+Mp9BxaW/olhS8X6w4B4ATrByHe2OLzHpNfV+RNM2xq+bW6JpDNuccAac5sX
WiR3H+tjzpJrPOTyAycWnlvxHl+bBXHHEa0uIYPjSmt61+mTY9UZdkcVfozHQhMe
5vxtJkUIEeCuqW0gY9NXkhazTleTq9uFItzujgD9vEqp3Gj4q9y0xMGwEdTEHNwv
MT4qR0pv/Kxz2LCKZKK1Mpb/0KcBRWDWiPUhZwwsizN5lxyppGcQMRvda9FTG7Gr
MCjIdH8aqwWC/hsVU+RiaJ+rLlgebfuvSUuH2+6uhg2yWmpsDi1iAj5oFgMAlDyf
vszoWujjBTsybewgyRzvDmHHQVgsjOt8ts1OLVoT50+YbnAoYafpvTZ0cxZCgrT8
Pl32mXPGJE0D8xqd7f10kLV4z8M1JcP5hT6U7d9pHCi9bV4REvHWG/H9RxuPQrVX
VWAHfFBp0GEnKanFKxGIkSGl3TmQCPI+PSHw6ReNsmhIFKvDgDLcygRCSQLcZnCT
Yjo9FROqTGZDFKzOEIeDXPMhobe9FuRxcFWAejtB8PX7BJb8KAusr0vZmOPUAwSs
7z0Ik0yQHqgMWryVm8+j/wDEnVKjASdo5xwTWS8QYtf0qUqm4yqSwe0YWRCx2Ihe
AJhXaVjVRnwwwC30QDR5MsLwrzg0tfizO63s7MA99vWEnTtU/XtAKDP+VYN822YO
FMd3aNS+hjw0v6WVGFh5So2MnUOHksaUMiD3JDwiFIcWbuTrnA5zVoH4pN/+HAxf
dEFEimqv2XVn1Wqfl8wXZxMruIJd4bWjtLVswzGEYR7CmTAvEq539nOHuqxu4TU+
SnVfxydmPKDNCwVDlHbpYV6D25Oi7AnsuhyOqPI5QG1h5E/acJzMcAAj4JsvvHDB
s8v6mw9VcZBe0wC7D1lY5JtucxaJBmtlm72UlWnV+jd1R5COejHs8ZYhKscsTiZB
QKmHymkbX/BmJ2kAF0LWXGsZgKfsrJ/E+ooGo6SIjABZNm5NwzkqPhd77iPX+H+C
aDJ+0ON6SNK4jirSgkcTlatMz/PrSNGAmlSawjDl8I2gbF60K/8qlAIfX+Hdf0/V
VDo8b/KF3gJsniZuPHF9vfCVL7nV9A1SMmARlqyiXgv3T7VQQluORh9VW8+Q52rF
jqhDNNEPDXlPEIkjswrY8qfR8RMwjVBqC8SCbGB7HzW+bQmaoYOUAsOIiwbnU4S7
c1YVnHO07vmtFBk1RT9nP8+2CI6k1hmHlKSQv6jgWxsXGnnQw1MJ+5MLHtIF273d
kI2RHtQxXCbnbHyCGLy2uwawyWgPUGd9TWDBKrVt7E/gFU7I71ZoKsLZU2wK5C63
5VQC3/q1ZXNq8VojkdL4COruSoQf8FMNOXP4gx6cFMgUewrZAWCRBAocRX/3oatR
FE7IBdKHaRPc2prpaAZiG7ZQmtt0+7m2TxkRxYyC1mFtWGTQkqug/yo1HWyFlIrN
Hvj3rYs0vr6zkDAbF1lnUwSzideuG+yYvalFVPf73muab9nHNFw86GP8Mk/6XCow
Tf1EEL37t96cjYFTxtixJfMN1IwLUmfzQoXy9aAlyNpS42B/mqy6Pvh4piA1q6GP
4t+wCOiT47fZszcm9xVNDF3x1GTQky4u91UUH5ydnfa6eUCwsyLKu9xGCwgjNkwZ
PQkG8RpYnojrpfFgkUgxImTPkngnIl2G0f0sZawiVEU9XbzMcsd/tuWmMDdvwkeU
4WKZ5TSixhPsW8vfVyaZLld61BvwHlPrthmHhe/zVtbPe/AQL7YPWmciWHmo2mHn
TK8rH8TbI9xZkvFOlSFkJt6W/h+q4H5LvFlcsnQ/japhKLlEvyapoiIdXYSNZmcA
iP/Cr6TPDgHPXUYONB93NfV86nn6+AtgDE6R3+LjcDAnKGMzlfP+fOZOdL6Wd0mr
oSMsGd7hZpr4pSPoDUn3zkDbO7cXWuJEs28VYzSFeoAyiPQZc1BB+3UxwO8QNKqJ
nOilLz6Y0+8vKjTqnzoEfUdbC85RDXmOt+QnDo7en0BxqbzBNw+rxkLqM8+yis2K
cxMwHRT5QTUO8zrKXDyWCcOt1th40k6WuYsuoODn7QcNgWAd+lpXi8FQxR1BQWXe
dchaZd/gMdM7w8IjfV3Qukhc7UJ6cmPbr6Eh69ksrrpf19AbrZU3uJHINff2+aCF
WTKZ0bZuIsmVM+oVt7hRe5H1hTfgmlMxys3NKAEnM66gFwmcvDHOuQSXuyfbrMQB
LnJqF0N7z2bZI6FTi4sXfSWAIR+w1l1n1fsEhSTVLQ0tkyeE+2KkzikBx9lyQm9x
wI760OyEpmdzFEY6mxG7mcKLUH6/uZyYf7LCbaUoj1hsUSfk0B9t4cNSM1d2wtLS
ZqyeXqT6820hCpvngN1SYQM0oiDRlOO3MB4MXia76E1tKGIYXZSkq48fgn63Q6g5
+B2xpiPJ3TQFSDcanOLMBWtiFIzqjDg4++tkW0of5iAEWfoGdm91XanfA2fj8/34
AZ30spDJwRXeESDD9iOczyup973Z8NeXzu8Ayar7REJV5ZhrCm3yj5FGtuQ2RtJW
3vrg+fY7i2uAK2E2OTFbyZrBkLYjVd+C5JSpYpw3aZEmg0VzwppoEu8NSxuCdsWo
nFnars6bGtzvxCZuZhwAfl424UmvZmsjhcggT+fnfy0JgaNdmfJx/dFCB8QyGMg0
iQ6Yd/rJtbrMlHND/tLbPefb9qCu5RBfTxWWlpF+lVJEp9Gineo5xCouCjJ/RXSL
fL0VDweKGxQsecwgMSb+URTkgqcNjAXr5QZoWrKJAfWFpasFNRr54XF6TRtP7vNm
HfpgGclAjIDBtsM+pXipHZkT+btDwyYFkc9f7HUDARuXg6ZliegpB3Yca2DL7i+G
d2UjxlqdWKXqSiEkZioDBgnG28tMhqutlO4qfRX+VohkUnvwS07KbCs96LTAcJNt
+6eXKW8yR6IzytI+kSMrw4AlStbTOckK9YMpxPudNFGUiXxtRQQlqRmMA4W9aWGW
vWhANLt+WnBE+ZNXBvIoL/KgSuV+/9CAC3rsLiuFpHInVY5+YYZ32Y08/D+xuMsT
3Tk8/qzatsAIr7cY9JrsBYjduO00eEbnqdTqN/+5vMMdFpN51k9t2NzNulBq8cQS
EHihUSSLN2+xvxSBqA+nu5GULzGU/b2goGux9UJiQ6frAkEoYJ91RvIKLtl8UfEK
X6uG9Lcv67K2lbMwRDZVVMNRXdf+U7101jNlBphMqbU1WV5Qxk5GcAdXk1wwuKfH
87u5cG4Kg8S6NMLs+Rc2mnwvHa3V8JpiOZCWHV6E+h8lqyIFNfn6Ikqt7UlLnENA
ZBnAKRXwFMlsHnREtbMJN5bK/ueZ/suwMoeyInP9f0IJG8Rp32OBxt4FbiK9rE2T
AvPU+z+9vJ4PQpnivzUKnBh1UjNdH4tJcY+iJkPH/VVJER36KA44EkipfLUi2KE/
kXdRlfgVp3n1NNli1B2HxWpS6eTRJ0hiAlG+kRbpRyT9Ot8fvGACOy4I0MpQCUbM
0VBqgNyL34Xo1lu8FXIW7YrXpv8Un+cOli4qgj5LUS4Cl4YAdjGUlRkHh975Z9dc
Phfi0ni4sknxG86V8+yiWDMiRl4PUImhRuiYe/2aCM4KUfU0qBc6FEt6V5p253oS
doX2xgztYO3hWwgbSicp2fFD4PzF1jhTqVTXbAnnNpQhKJSJkpOckuM+DtZfVIFh
UZClq+iJjmIXlFnina4vrZDZPEaRkyylwu8I1CtFZQJEeki6OIAbfKk/6qFfFsFs
ou7KULo8cUfnnE+9uv6pEQLJp/E920clzNOa/fyfCtEMF6W5t8vazVTagz8W5ShL
4X8OeX31FbTIoAxAklQcr2ttGdXEA3tdLYMRmarNooDXNN/lmRhdMCLb5zdvQR8l
DTtLTzCtLU1Gi/4ODzmA6WeoTwVCn5spFwU4BVhqmpHUkUxeagRG3Db8UHuWS1yS
yJL/GoCA943ejGXe++x5MOP8oflG3y6mo8IheakdgrSlkXbKaBmpvcg5u5ajcPf4
+gHlUzYY+Cf3P34q5tm42CG8gxUhP+O+45xremizFfgZBABKmP3osAjnbD0J4ylY
iaAiOP8iz80sUdsg+JADQrcv4adfgFZ0roo4qTxN3n/uRBCizfDxt6Y7H0OTKsIU
ReY6LWqFqSLDuFeyg6WLzc9tfRKOOEvxzRpdE6dpA+g+CJAdpAzKoKkmbuFH+LDH
UvO99yzHn1+gsTYPwr/N0yywu5+gVjyHu2yemmkr3OmBSsAhbvsBYqOosiG3cS6n
f+be1zJe8YXd9hvKCX+3jZvbH4GwtK3Fz6EFRRMPQBXBqd1sQLbqMjeXEzGcEkGR
fCTn1kx/1745nylfyLuKwHsf+7Zue37gpdwccc2Mtmj+/Be+U0h79rcClQju6ydE
5/B3CdNXDInWHeFrqj1Cj40UwE29qilRnR9TAqpKb3ZDEhGpufe4cJ7/KGdk9gQO
fZgs7emZ64g1XAkn2utAckiUO/hNRF2U/Zww3mWWuRDfrSX20z2FRxQFrgY8805e
OS6HYmRVOCBr9rWlDHacBaN9C0z6Fe5GASWiG09PbaZpNJHAp82bMVyhEbs+9ct0
5rX9c0hyHSQ/f+m8FMbwH/ze442YW7/iDHEHPZM+95o7LaxZ7TFT6BaoRmF+hInu
6/QKLNHUJMRSf87hf0hoTO/bjnzVi2mRIi8fS4LheiMnr2Xza6LCeMf7L1bv8rDU
xQskYRQfLx+IJ5QXShcPZ9XlNx84D7HmgQ46M/HAAQX8yKoxEGAT9TKaxQF6xDQ3
3nIt36NWJ3yvvSI20V48NJ2F+2tEfkBIbNdF2kgbhcaNAHUgXEG8SDavZhG89jeT
3huiQ5HeFivDwHDcbsFkBFXUyhN3ydKfr2o5HIh6UpOjjc3exdEWT5j138SOvdGm
AotEmPH3vaGGxlLDS+k1qseat9DtmbNpOaWaOLoAOBh2ibVOZn7yyI4VZ31DnCC8
j0vb0vPf79000WIeDSvjBaqVAsVPN3cmVqNcURJswBIaLfs3c63NnOcDBMvtT62A
xVKBccMVNdupmv4XF+HXREdJtqoqUKgs2QLzsY9WwdwvIZIfXTbGopQbWZxMTfMo
6k0R1UKsBpLTQR+Hu2SKdUB6T5zxd+o4ZIugMHM4Lh7MimuFYBFYpaELJfuBVMjV
aXWQY9LK9zT5Xq8O2ML70TPiniZ+DJsX1W4PpGPHNrd7M1Bv/F5kLyBWVT68NviG
ZLRcNa3diNymoYrN8lzbFb7InRO0CMgkmztrHVAzyP76LsmcuGW9IqL0j1bIy0z3
uTgZHU3fJ8Kky28q+d/xPUqnfkAirCXLwVrzQFLuAKZy+8+0HRQVzaZ6W2f90oXD
b3cEN5fAfgsxlRFzR2Xts6ENldl5KUfF1XIUW9Q/+p4Imj0PuKc/Cj6lKlFfmrj9
PquTj6wlIdGbc3xIiWnJbjB5ur8gZ66QR6Rnd89DYORv+UhkfhkgpG04xTpi4/xV
/tPzYfVoU0rTKcYmNW14i3xvFhQOEfsxAKV937FqV3dlNJgVJqwak3SuTmj/DqTp
Y41xeL7Cw1Lhkq4eAL5mUN7haVPJXx44pAO6Ru8mfqvlmCVJHMQQbFex3hZgH3+k
lVfEnxZEEtWP9vyfpCva8LySDxgdHWAblvBLGeFIAyqSGc4i3eH3pkQ3I8PnF1nm
VwLnItJd0KeREDwn5JKAWDGle5yO/mYXwWCdEh5cfsutDjBogNcZD1T72Cr4/xjT
vd77+fV+u2FaIdZvsYN253QuBL/7QmHJCVIZyB4VCgOPLkWse53ERgyOoRtrvS6O
jFjYs5qCJ9Y6+xQop+LK+dr3yi0KhXUlr9+SwOqf0Afeak1H09eJu6KM1vfvVwJi
E9MntOdtFDViJT/wCr+u+d2ACm+mtPizuwvWA1f1dxlQNUW+D8NQV/C63huhzyUE
qhLlZHL/+tjxe+5avd69BTKPE+EYbaS77xmjuSN30ZQv27W91Q5JraC+aLA/u7K/
fCuNw6c4ORwHzoaY6074S6TpugkXxT8s8RI5w+DWv71uN7U5VgvWQeHQEN2KTrK1
6iYc4QXQzLsN5HRWg/Lnjk2IQGPz1lDXpn1uO1HCRCg6zeiq83UIFo4tKop5KY+s
hSVN0+OKEqDj0saG75x+0TNwLq6jh+atEK+6jGM093hV+IXERuB1zx6BNbV7BJN5
c3kqjpPtaf6NZbH/ftmzwaolVJLohXT10OciT4HuU7GsXLb315auZC7jl6Gy8uY1
0dgp03fbdOMz3IuJihS+Ml4nmxwoS2waYw/bMHBpO5ZAyInZnhWcYQzXogT26R8Q
oZ4PdmUnQrs62lxzncU/7q2Y5Qp42dQbbKqU6btr3tz6ShPqM2ccgGB0gPuo2xst
CVCKgntKo/94i74QrHLOuOHGt/xrYjD2PARFDWKmvElbTLJZ0aJqdByjCdwJq6Fg
Yk9jJ238EqqRw11hEEEOdpgoF3XXU4chNM9xWzOgavpOd3hesVHoSdnXHrrJ9TVH
I9749vCwlwiBWIf1jSU0zB3HYc30H78n+OFZHCJ9TK4mR7ei2cIx/WhrD/ektEXr
l97VXTI74SRHt5CxjRmSphL0fX0UcXq+AI5ofhRdt28FxCDmJyQCpD912yXpAdAG
aA5LYqO3mrbD+Xf4SsZs3bC3CFjArf+FjiN5CpXwzZ0xKMqJirDYMt3ST7Qv9io1
NNpoIIEPyZicv5qzttwTDLSJIWjhz26aDrogs09fDfR+yu8ts8kJFceYAMrbb+1N
3DWBxRh4swH9wuhxzrogKSErlhuUkIljIOpjPazSHTpL+owM/1d6Y4Gzh29m6K+p
jvdzutqsv83B3jhZRdOyh3mLiahmLc1KarxuBD8PSfW3MTEhO6yPCUd4iCxj7IRK
j8N3gEU4SRr5Ei+g1lE2MV0t566LTVY/D2ruzrGVOJ5IiWse1cyCm8OLeo2Bnrd6
n7fAkGN+6ibN94oHJLh5O2iggLPNg5d90EMygmaWIm2VoMla2XnTdGHPJZbmbUix
MRekqV/3o2MN4xn0vqeDugiqrwFcOvN89A5hf5iT6tqij7pupDuiCr9pqzsBcCbB
QVQSDVcP9diqUd2JVmRXSk2Xp1wSay2ni/hKEnX3Z6TGaFja/u+Ef+YTXO0tAwbh
npqcKMyVGpMSOVAcee1TDl2zHSyuRRYTHduzrr7o9blRr0MVYZrdWnIt4SRoZ8kC
X2w70HKQIqKzatWTEzLegm1/iE9LGlaE/z+8Cy9Hu8ece2OH2QzbG4sdftuxyp6X
Luh28P9w/GUw+mQilqackBVOkQW7PTgcbs4/WitXhjCGKraMqFTbq5GKD6NcJgRP
kg7142jI1eQ2NvkpHiDq9RvH9Gb6HY3I+oJrIGXKAf5R7fgmYhon6fRbJLtaDp9Q
yh/ipmk1mY6SxnTF8C+5pJHbtRnSlxxjTn76MQ0p6NeLjRUJFuu8V3G8NpK7HoAE
c8bQcwBhj2RAMMVCNiieGuZNBP7aiDPPeWptIhWSaQOOjFDVn2ofqZ7+oqBxoUjB
bDP/2O+OWo8CUBZ3twUGElsxGA9YT/mWK3IL+O71fD5sdZuHqYGcONvgGl4DmX64
v1SdRGv6UVqeyZcY0M8K/BUqs+dA8AQcCS1gMQIxCvfjqyDodyPjaekC5jt2Yjd3
+HMLtf/UzVIz9z/jGTQkJj40WPictNoWRJ3caLNmkWzonck63ybjZHC7Y65XG/Pj
vsdhd86Mfdro4Gx4a2JbepYZABFb6OUc7mU1e/6bCDyslR4u2pIRsbJSB8tHk/ae
6DTwB6sKwP1odszjYsWWQDMJMY8hmANeEi5P5nhYgtEJ6Gii/rj4apE5C43xmWC7
FLtFkHjzBmFyWzp/sMYfc9FrVf93HhPx4b3bkRWFYqT5WI0gYm0UxrCCQRzEPiSo
4AICcqNTXEVsHCFYr8AGlIJ2OcyXuW/uMUQQXMvhlIZWC1uX0FvKHTyJ33PEdGEv
0K/zXHCKXXvR655WYJKZa4EpCJFiKNAzSLgvqJQnnpRxcwWGEhUPEsRV8TYAQx3/
xIOZqq0Xv8y+cU0hJKzeWY2nJIFQPG1aT2pqp5nYKQqFtGfZzyqiOZCn6Ao6lmxc
PlorIcpJAfqe/FR5lRjs/JDMpe6wovXHso/8dDLkUg/xUE2NBlfD37/rdiN1jy9Y
HoDngzmSEhzkpb27eEmv5NjZNwK5cplIyXj6U3QFuaUn/6EPaAsZIQ3GlKJo1vLQ
4+LxH4RdA0mHOmajkqameoATCreG/kEDQlN2lNLOUPWtHdiYTkbgujDPwpii5GEu
gwP6Pbjjq4E/bAWQqGuTQu7c8L9uDcoM4k0d0cyvt6gbEqjX2IdrbYGj/hREOQUh
navZ4RXUcjvoRF5tvDsvzgfw2jIEr+/iB1RUXq/xH1e6t1eo3fMKOGVeTr1ZPCLD
9RFf9spaxicGBUHV87X+rpn7zreXT+2OXzUbAwfNk8VUs9m64crd22heeStJozjk
qd7kpWNLIBpmGlfJHSWPgHHuyDZGfcm2qIVxGtAoZk4N5dl11c+bRuUsjmm6NXdi
wjrKc8SZLMqv5nTW3DZoeZEg3M29+Gz+0eQR/vGNM8Jpg1gDBZENs5jliZ/+D93o
dMPyD2Y6r/ZPq3Iw4tLANhf/Evz1fZZpGHpx69N4Ecfu4VwXi4x3fqZaslcgeSDL
W2m376e0x/3vrke3qfkyKvmDJ24WlRi66BtkCvbbOSMG1Vtwn2ZJWgx9BgGZugjf
9umt2jSTL3leetyuEYLXC8uvNXyZP8jMr2ueHUuC5koIJQpyA5kDtNU/mvaopdEL
PcfS+Hvuzy05ukwdzUsPWRRr4GoER7EX/4UfqAkkcQN+x8VBf7FdBiAfw0GhyjZ9
wt+q95N9PY+ARSCE48lHtuEm1zq5LcnlKCf0CVnkslOPgINHvIWo2LkJb59H2XKt
7qg9O2UqvDq7fDIzz8eyRekHZN+UtVsBZSyFTzU82HbtIvDyQTgL1Ppf1bJohOwq
hcLgL8+ch/c4YLDVb5u0zAUSGjPJ+V+qo1QW1ZG1UcWAwHCAUK8S4NHGvmBxx6ga
T3qjeu6k6JcTze009Oh5uH+XGyJnqHmzTkHb0cHy9iP8XdfyhB7zCa3jEyksbbjZ
8uCif+II4zv92RfvcBaCwFG/sBl3xLCkh/6gyVz9t8SBvTH+GivuAPcU/zFgKEKu
PJOdsXXe80LdFERB5OGMIHi7LuXD5Ce2+NdfIaYMua7eOWTjKUFFyGlLu5PIwhm7
TPAlX5+KJejUlp8pHpk66KvzoYb2V00jeMkHc2s4yRrxbt3cB3deyUufD+5x2LmW
1uJzp+og5zg/LJYOuEmwxPOz0wvfvRYaqVV4dYi1pJ5xQgBbbKP6TKCa3fnRZP2L
7OXCpd+p0nAOdqEUP6vmgu892INVNxKx7bmFgultFfr9B38eTfao6xppa7+uldRV
lKc4s10V/cxYhKB+2T7qnXBDNEN1jv5JgXVDu2CaWIHrZvyG81AVCF3H4EhqBUaQ
SVk7RZyItdzSKaCwwfPcD0SyX9JcgTp/tbgc+gBFyWIROUc1gghXhnRyDB4ojpHk
DuTzmTQXykNsSNfPv/cqcFi2A1NI+i64g5Ma5JCatCFbBQoojOdHxUYjpa97WUEl
EcT9rp6688nNWQor7NMQVfSrnxrDg2AYpvSXCMn6eygFUNHpfCj638IaY77ishYo
VGe6bXBYOr+orSIdOa3Rdl82LD99rsZ5H0IWjm5mFDyQf1hQ2DEywqU2ucHuyP2p
rs+YrUTIDIICbOnivMDuYAGXZzVOi771Dv/fr8tG3r7jk7ljAty51O6N+6V2Hl0X
wF1tGpazz5n92zI7BMiiI3f/lq34S4DDcdMRKGoA3pz4rH0/1c0HGyGtjGeD7uZe
omp2zWilRMOAxyU4QOhJG40eXHd4/R+5DwFNsRh3or/Wjb3RI6NbzdgdofGn0P33
bEKj7ezUDKYb0NxKeY0Vpo6+MQvs1N+OQP5q/PJNerSBdosNRqQOjmljwCDa7B6M
EMUqR2WTK+6iUU1Pw/km6bVmYJQQLVTKrFYWzoivyHD+ros2Y11Xlz50wbg/+/tH
OQ4iiDJR41kZQry60SDhEnnKjhY7ercDQxXzE+uZuFh0L2eWaOZ6OCGVkSfwzEgF
Z5UxjCoY9cfXA63hOS4cH7/F0pCB3HN7N63qNl2pguQVlPXuz26o1nqCt+iVx/3l
WSgadhl7gxm6vg8AcSMw2BuJ0t9PJEFyHqSlvrrKCB7ZEbeISBHiBbhSm76JOeYg
3UvSXLCmcIhaCSdwBpQ52v50c+RR7evCayhjTym8w+rjUSvZ0WZVEBfDNuTwfK2K
10DMLx9GtepK0IZpDltnkc/nXPy38zD72FQmh4XwAOITuyKr9u4f+61dozL1IiHM
kpsx2blY3nDqH72+ROGph+hVOUwueObb5qKXIlHWSAHCNPqdNXPLQTF32oZYPXH+
9crq/C9rJr+0rALFcNfU+Jm+qzKnnkPLGqXFvKvtNroz+Qcq4tuxJPiHNs68o/ev
lAk3m9YVEPWt1wVzCJjxgY6dgkY0oae8ReQm1brXSydyOF8dtDI2+qufFVFwO4AY
rytxgV6nD1X4opzvNQv+hOw0x9lOhTjIeZb/qitAXMTuGHUd6VzizNT41S6isIdl
9Rt7a6fH0eYOqRwW6E89Sut8gL0lHXnXSWSkm6GMTY9tPJ36TpWn1U0WaCB31XYQ
J7nqvBxc0lBPjCmVne3NusVmtC1II6Jh19Rnz5BLEcBrlpO0El2jQgHJkXhOSxrT
ZpHAx5ly3cXATO7zT/X6DLUF6vkjU5Ev/5eLUS660Mq7O68ycMyUoSxZJtuGDKOJ
NjOARBHqgIIxOSI4SJVUuc1uwISlEL0e7cpQovRE8MgUYZSg99xPeZXHiPRnsneK
7fYwdlYcjt6DC3wm6lWs+g3fzTyRwPbWFn8IPaUIlu0sCv6UT1cKa2C7XGQTNr+A
r4svuvax3nFOhBlDmWiZP++hub+RJ58CJSYWrPTckSjI7Ly+qJu3dZcqzXfgPxTd
oz3fOBkGGjBFX2keDjpwyD7OwyFwnXeNx91prdsmcrhu7BW2zpLZfAcecJU7ortA
ZBWGLLZkLOnHz4/XGVoajyK3PoQTem8UwpLLFQyyrGKMRzCQgGTYKXgNSTJiugeP
bJkNc3//EMDIWpXNOYLL1wOn1OTZUkQghGSWxIkEzyNR9JGDc+S49MFMmxaclM52
SGBPa00VfWxU3Du1mXCGXi76nymIyANuYONdu7p+qG/oLCg6L9aA/w2GVM7wmrae
/GJfuGn45UjRtJg6yXJro6CVlUooMVlju6+vgZwvL7gsZOECSjiE0ghVx3VBGSom
JGGwO2O0MRBfFo5m9WdPZuJfs/xf7cuyBesiJcNJZ4z30vBgWc0Jui54qqz2LJTj
+8B66TCsYTv/fZNGJ/e4NAZPm+O5XtItsYSOqeelch183JTBIGGSggWxGBht/3fg
3cv830zZmkkKE8pHH3Fj+2GtNJG6RFSPPaBzcfAWgb3XxHskNoxAwRu89qOH7U+v
VbJOzkMGr1ouR8O+7RJYvh5N2qXkN4rKEkS20gdQqlPtxvdGS8it0fwJNR7CE9yC
ILPqRGFOaZp0EuNhJ4nW7bSMAIzp/0/XxrYeFSRhujQo6i1Gbovnp1wwgF2P8vut
WNcTC3/avBXjVeQCrFqqUGoNvS/WpES/quk2xblBsFWKw2S28Ct1bJGEqsm9mhEO
cz5Nh7yXRPEx46Vyz6sz80x9QYY1u3C8DhfOXw6blVfWG9sWRS5NN7RAQ7+WkN0/
j4Z6nXpg3dgGvKiOUAfaclll1/GDRor1+RmxYFkqVcGfv1Q73x9qRzrtH8wmJX0E
0ti2xmZp/34AL5jb9EW1Aa+4yDiVG1AqnDKZbbNguyRWejdDlqnPO30STDHCFAlI
p1vUFrqIhkiKloeE/JcOakKlSjAQScxpA1BApr1x1QI2bvW13Pg5yPiwjMs+EpMx
s71X2FtbF7vocRv8eNWRGLgXnhQo472D0mwrGtlsTaY1TZCPt+F5E3gMJRuustpO
tpOvp6WpQbZiNWoPoGBULpg5PFx5OFTrq6nPWEnfzgU20bLCxEG5orlOl50zRSgY
zWwV+fPEn94GJdvfQJZuDMKbNA/0uNVXo0KauLFlmbq0YsjnxV5bTunMu4aSUGeX
oLBmGqr2FbyFy4w1B4MbfjX9X+iNlKrFG8evebPdM8luFJyi7pRvgF4GCaDJ5MRs
xQGzYeS/CbYkesrj6qVVRegdXNR/xlMFGtQB5W5OvyYM4bG04gff7qWhEPEnGVj1
ABuznYoZ2qSmGYnvWcLwmFiir2to4R+rVJzYRAwfGc+mZ/QOvaqxBV4Uu6YcvUS0
weOo++wcJmG9XbSzArE+/hExRVMkdTJ9kGdtnDtJGQrI+IUyYKpQCAW5bVEn8xko
R3teDgPdgKlZ+QE+Vak5y0WnfJ4F4Ym9Q3YbC4DfNZFWpFxPsMJZLBz0tzjNQ/P5
EpEkAFvFX9kWU9QyuzhSI9bKP3gFB9Rbzm3F8qni+7b+mO94jiEiUeGHJMXbek1r
NK/ICfDLGEv7XnDlczr4eyrrJVJG90esQLr9G4aQKdyWU4L6dL4uyf/zDXjBVNi4
S/vAqo7Q40uH1rMm6v7waIQwP0hcJpV3ZcOwGta/h3ssyBugmyNUafX7b7TB38tA
D9Us0z/afGxYmW+kwvl3f6hXqzAmfILmHCjKPDJ3HYDTkTjytvZwU21uUOVffLJn
KWLCxLq5LhKS+3w3Kdjh8ayIS5ukgwG/kjDmn5Hvi1+PmgU6SRaYzKREowbNSSBI
Hu0R5EisbqWS8OyF46C3iU4W5shGFWSoSuxZsm6x0OR/me4H343I3r7HOi6h4aCS
syOZJ8fbeh1LIpSv/XG/GaciKIUZ/XVCqymSu3xiV3yLPoueGLqp67XH1CjYvnYs
O9dQYPnLW7e1o/a7WX6kl5dutN+x4kSGq7jmdclwhcKsYxU6VtPfD1aRdzBOoH0A
Gzp/f7ib5O4PQxf8Th2J2P/My5ZE8mZlGUHlGqi72FVcO1TrTF0u1lCdGTNKTw5N
3Ls1jxAW1Yhci+xpepzD6cV5MDszlWTueJkR2EbBDeXWcO0nY12SyrU/EQQ7YWDz
ag2FM8nep0Ab9N0WlLCVqbt4rtidwdrPqfMbge4EVeucH/4TW0MGCkhLUzTTihpL
jMqe+m3DAHtjllPo8o3zWUW/4DBCKn6iq3V9IIsJXQoWP900WsGPgtHkBbs2zM5i
Xlckyp3nAICoEG9Fzmu9hHHzjZc1iakFsCC9VEA9MUDTq8ZjigDg5FdA6wtJpuWI
A6UBw0huhkY62ts3XBgPJcuAJLh/RgF1qYOhRl3aWLR25ErfgvdI5xiQCCCm0hcC
R94F8a5/GbOVJFeXW5siDBih2kcCwPsg0PdWugw0tbCFt3X40AgQMDJlRXlZkzlC
Kax9RHPAlzTJnxJaOpV8S1boB4snOql3Rrdp517oI60gwrM/CWMSFFwqJDC+T7Fy
tmlB+6AuC1LjivQilvE0ytZuQ6IsQ/ekJSC1xjBhdCMHVthiG6OOEb8jmdowzTrV
Z8vlNHhnqObbRxdKTdopzfsU8LIzJjMrLmQo/wtfaKeNY6HcJ7Dm8Q41vSxdOOEs
kjzMzPe+wlH4cpQ48rrTrOHYjuzodrVRrHkVWoJtTZZKBBSDzPp4ZIpAWXcVVy5c
U1RC4MOAn2bS4COo5HeBIbi18l1LuDdL6F1JfJTV+J7R3fILShyDc/ef9xKtsfPz
2GJC73j76O8A1w6y79uNBFUUriUZS7wz0lIuHePy6CvPE9bx/p3ZJPQAR1GnBpCC
wBTtGh2OIpVgFHuoblAj0Tx/cxJkcUkxTVDSwK1fUtsBesBM5p8R/mGkXk/SLLWr
2iJfKyju0tRyhWTiPRwN9cGUaNn8/TuxGHvj0+NJdBRG49LSqc4hB8lHimI8MOum
aWjkuGKc/7KwAjSBMioe7dFObR+AEx+Sd5NYWFneWggvjxAEqreCeERh9Wz21Sh1
kOvvzIg1EG0IYMNnDk6NgHIdoHCdXVxHCNkb0W8PLe0/KBQnQWeSM4uux7ItkKAC
uHBgIiWs0ivSv/AUmA5sCj8v6Ay5a7gy2babNLDOKXjO1GS9xOCtYtWDllSDXbnd
96rdyeeuAmBu4FtKh/xuDLZCO0kUV50wX/5eh1Oxv/gcMwOEMuCHz+nJKLwZnAft
fpfuCS8kadN74MlU9e4ZJIGYmqcZ+gmGp1HwjTPByEVRPLCrDZnLwWU+hAdzXb7Y
ROrCMA+Ytm8KoPI5smfMZmNGIW3Kjw+7taZc5dgRogPu7hAwxbHsN8uFPsfbTB5C
S5FntauqkwDz9jwo5HHIGbSIOy+caHYUomWBRJc1A0uS5QeWDH/1Oh0v1VE2i0bY
gAJdP2mQezkriycu28DdRNKnK2YWjK0RXXeue1bMdXtaMqVM0fmoT0zrZ+8O8pDc
7KgznmDvhUh7LGpZA1Jn5/tSwj6Y+H8pgkTlccU4fhXYNaWS3wPY868wRjkH2ySu
G5YsWo7zL8ynL2xWuS7YJJlCc2BaFQ+eqSUz2NGuT1+eQ0/ygHXUpmg5X4Ds9RV1
wkd4ufa0oOCKb1gNrpqP8fGw55D7oxyMA5FFkSvLd4/HkggPQIMSmHij9pTSlzeG
de3PSIyNWkQZv2kwSzgZueazsPebTkhIpSGFlJxCZwl79cfelvU2glKHTVcs9P5L
TAQF8lUySdOkaWZYNiqjfGoBQQR6sj0ldWTvBK8jY5ayymidqpirpzOBzbuiqjRJ
LIh3lH4Z/4Q0GEVJ6/+8Dw0T1TE5KTyOLCQ6dTSykSrEcX7bFd8WfrYmh/1uSNvS
SZnUp07YsN7uaSF3nCAcjjS2x609R791EZfG5Bw8ERGlhkUsTw88e81anFFObmYH
fwDWlEfHGC6f2NSrHmyaXOOlI7BkCLyxcuRT5BP16rFsLQeLw04wD62/gpzQUpbu
AhYwfI/7tnqgsQr0vU/HX8Hu4t0/OvCWN/tSsH99yJKA67p6t4manCP2t2xsI7kq
8cgTfJRmKLEBjkg6aCo0wjXCMie6sqbt6pjmzvYG5CxmjHtzyAYIL5TFRMtinPPc
x9G8vzXng4+zmJLIJYOExxT0kf80gRSJDcWaKW5iX56HAEZY90K1uiM9TtUX6ptT
eJXGxpGmngIRxEJlBrm0GrmNP8Q7pMYGXN6l9Ycrrdi7gsouBSYlsb0NSC7DtSO4
R57/hMqPVMFtksRTU14gEXaoaPyqh4jwyOl6HhGeHYCsQYTv5drN9/LgNi0RlfZ/
8G/ALeWLBpHGbKq4eC8ltuCMM+7P2O/alGl8Ls/WiVcdr2hrkeLB1QGrx8xnonYo
0RfGAoXPQhPWc5Z6l+JUiHLXk3Vb8TUgLqz4dO/6umRkKeqV9uUzF0F7H9an6Q2p
UNdTforbDj3B5mJ3/VoaFSkN0a4/UM+Ey7i20PA8/TcVHqYuQbpBaOXuo/47RBu8
XNrt0LBe4ZG8L97kt6Hawsf9aa+t2Bu4IBuqgpeMAbIVMJcMvrd8Y8PQimPuslMf
Md9BHv0Wry/NBdgGdS+FK35QgqihQVnRKO8eOtzauO1XcJ5auj3MuRH9fp3FA7w8
+3MXchk7gdS6ziWObxSEyxyxUAEiPe+9IjSarUUzjmN2eU0yGocavGpZpY4E8FOA
Pu0AhZ7mIdD/x57vbKbnG/tUsMKSQ+30kCEg3xXU+VIv5qlPmaAXPROSn1io2CYm
dP6Fnr3Sel01s0xbUlMVYlEtwNIotEWGXiOge3kpQ6YKyOv/k7X1JY86Vl7DIRjL
hZ9if2GE02HOBgfEXFY7e95HBgaKPQtJy1HcLa3F3z6oFb9dg0q6Ey6v6/EHSzZm
BITpjKd2cqrs2sAb3nQUg7uU9t4SfTqNVeprsAuvtMGig++ReYyQCIrtZvrTgUl9
3uBBXOqsXRGSKXHq5BWs3KFzX0dN1Z47OifbuT+0ojCmiCzYQg7Sbz1uPgrnzgyi
rTTyNaiC/PgDj4HcFsk594ypp1EnBYWaY8BlFo48dCR/b6vYW7VdpHZRw4lILLeF
LoPyxtSve7ecs/eW/SOP6EYaZ9Ly9D0GwslawI5XYYpvVlOsZV1awB4PV+PvDE64
MxO20TkTF5YBiPqP5XTsUVnYp4AyxOTMaFc/wxgawSz258FZwnzqW496DKb25OyA
CSjNkV5/BJvnYzJpgRNerhXs//aNfOSnTI6ZMohqRJDXMxJ9sLew5hRIVXUaA/t7
mAsrdGqu39tJzto1/xEjzVMCwUjaP7QWvJD+Tkd3q1VbXpnQ0ZW6ed806Zu387RT
MbWF2+AbSWpHGHQHQKSYBshOW48v4TvTg7F7PEHOmVsIxAKSQ3BpKG6vormxG9/v
dYkyoEd5Wuefx8easWdeF7Acq/q1pf34Tt4hWpPs10YT/9+52KGSqKe9w2Io8QMf
Sk/dmgS9iwOruUv01K+nZoNxCU8wMPW2doVdFCpsY++aC/jrVLUJHicszAwwQRW1
T05QKiQjjclJ7brViT/Buuayz1rfmAC6dhH0LLWjnGyhvnk9bMbwEQc7yI/0o3ld
cxsSyxaaKu1+0l4AXO+47LA1Ab5d9ZYOcLQbDTrLxEU8vJSpBNIh1CjWyXLPizRp
rV9pC9IKAMgx6uxvq0hHlbwd9CvAhr7enkG72HI1d5czWtSC3B370A/u1pr+A6ju
axjEexJQ/hVmhnvDZXXuThjQJ7vpHagkl1B4FGA9yNrunyVFN4a4lsrvUzxklgHZ
jFnhyeU9UdKPoBHnkHaX/1FZd2lC2N5zK8dluLLwvxbfP3TKBQfCstXo+u2IfQZS
wmo1qhnlKRv46Jj0OSU9L1hFYme4PnOgCiwLy04TAKCgzCIr48aIP8pKq+J0Etf0
8T0Uw6ItPMogcuixIgIngf4Lu7Bj9y6kz9V8zgiH6N0eKOYNR70c9XIcz7j5rEPI
PsGza/CWRpxla3EMJ/pVtCpAFzbCk/uh4Nxz1dDZFrXjcsYF/qXaDHbYWPGOGNcG
V5UZw8MgVZozSpms+RhDdjJ14qNBeSirbUkY85vd2l46q+AkMBAbBnIhv/QLccIZ
dVRlv7m7DH8/Rx01HHsucWJeM2aKHH4gSNeE2tgS0AubzkT/9eCmRgHF+o+DTkDe
BbSyR8cNzg35waKHG/rrD3vo7aDuMjKnsmlArn+dOsBus2copH7eXLbWX6ZC+MeW
ajGurQ6uv0GudXor2XHtcm4RWtZaro/JpZTWqjI5iGh1dMZuUEjpU2a8u3RZ7vwL
+JPBv91DrGYocJKyczXWiTjPC9o72lzydImqD1rlSY1lXOgGgvIewniuJXvrocwU
WWf0c6caQ8c8z2unULOVyROwhV6nb0/JG6QRjEX7mguc4RUxi4YfDWlknZqOCGRg
Q/b4MS7iifs8R1HpfBMiCDjiN4HnGxPrlz1SXTsYbOjl8PNPpAh5JkGf61aaHaOp
QR//QebULgBAsRHeCbwxXYUnQdpZdPV5373dP0krYom1TArEWnVmcW+4AA0mDFuk
9N2g0Vh+ZdPXn+wjBZ2hHum8ZnzUfS9e+kJUSCEQBBEUg3XD2zetGwQ0HfEzEJLO
vN9cSMqzl7g3teKfRFTU20i0qF4AmzkoXtnZifZxzzZRFwBGBAQKPw6ElnKa6KoU
jUzFostbzLWEgogNccbKI2I7zIzsDcuXJM8mwpYxGbmzjLr1Y4LtR2N9GP1Sle0b
p5RXq5DptpDFR/N8NywcTe6SmpUPFFYSmymSwUFNk+F3J3/MKjWD0+2wgwvU8pnt
FxmG/p/9XY6kp7tLvl1IgeVxWBDv5ymr9+sEukWAqsg5wMmqjCyPdszCIj/jwGZM
6Xm+pXo9Ft/a0cQ7hS+8aHVD+xLt6PXa6DPWeIeO4qmL4PXe2vIYrHOIyBIRrLYo
STF19fZSzaXoyLAH9Z1ZHbKM11UwYhq4kv/6tMsfZT7ShkrK5dbRNt5JFhPWyOQT
vUBecoOjIkMeK3bWNzaUmYki5hjrLKzafXkZTTx8XWm48PsS+8FGe6XJPfbwc8oP
JGUlU/VLF7ZtL+w5IACnxpE3IT+uYfdHCT9kMyj479wbE8N67m+N/odxs5/PGl0F
h/0MbAWKz6qAsOXKlVSWdjmfSuIgQ3TB7yUfkJ2uhMgVu54W8GuFdNBL6pANSe+3
YAKsWqve+IL1Y4jfwDlQagRVupFvTXktDFFRogN+2Zbfw0dhrlKo3DDWhMLBFO2E
zepoZDIoeA3q98l/wEp+2pF++yI6DGvFmO9xl7AMBoBLrSGvBtfqlNygg8UCmHq5
eCB0AByYEZIc0odauPeaY92Kr22OkMYA0FVkzTCsdi2bvKllVYY5ifY07opmhV5H
s4gJuBUVKTeijL/s1AUxKwC+HvsGtFLyIgJ579s0dgltARfal5BUYLWjnOn394bo
mz8xtwrkamgwSJnK+HfiMN2Nilw4tWNAhB+0jTEOWTS6EPvaXx7Bt/LX9684Qpfo
hOLt6hjI0QJw2JeVUz5yiugjiCR1Q82omFMblkERTX4b0EFK5fdmEYnNnHnpL3uU
j2CnT3iD1Joq33uTm4Vmd47j9UH16402CH1ouSJsh1pkeXaLEh2Al9XmF1r+W3xX
exFViwIRtuR4INc6mSA5z1KiSO8YxeOqb/GOJ5pytQ1KovBWR58DC7DBWRTgMH4m
WB6blwXrM495o7R6pMQi/Rm5ic0vy30xpx/6e19wvKXd3d9JW6vXe6xJvgH/iNH0
KO20S28Z+lUeVguW0JnScBnJvGIB4LvedycZdbrg+bQ9glmHROEUN9ujpbztvb3v
kbsxiHWl9Th6jX9+iH3jyMbNoxuCNb7pFYMS7TRtEy77Ajp5M9Gij1jnQRkyILli
TjAOARPd1Q2wSffy4nsTwS0WcKyPNh4XkNVsQeu/gKdtXWCutKNwi3r2DQjOJjm9
PFt7X/8OVD47JhDGzvek9XueqpvkZd552AiGs0OYbxA7x5Tn5N438IkPxKVRfnwL
foOoRVb3ivIs+nKp7JU5BDNxrkjo3Y7BthW9a22mkpMvb1WWkvz/yvnB2MyhrXPc
tMg1Vek554GnwnFCa28FnaqMo7X5HMuBJqMRxHy2bzCkHvq65q+MVAHMV9VLVO0n
ZDrCQBnwCGnKeKxsW43EGqnvMx7FeLNEKlvemIigaTY5dT+Sy8Ru4uI4NAsaGHCJ
Pu/Xpm0EiMq2YXi2tvQkmXcijtdwBvJBgXqJQQPXre3qT7e+RSxr3vkz8yW2x4r9
PDsHvFNGBCzjKlvjsha5eadCG1/C8AdNk2sQyadY2E6YdsCZaURwG3ICcPk5ZAf0
tng84Dz/aR6R9GBffi4VKepaGpweYbN8E35ZrvdbU6Uz3Ta1f2yXi0/XwQgf4hUh
3xN2paYNEbbCA7zkLktsri6pRHqv2vCMB9F0V6obi2BxFvhczcnbyojXLJduG5KR
B4dtXdQCWWb4f7Sqk76AmDMwhORFPu5JHYXwOVW2La1JJ2evzoFgYIUfg22s2BKU
RddCBaC1sulnWl0JuFt32hjUPEES+rc9us7+NgiaGGiwmcutemBoz+r81pc5KffN
R5KcgfBP+et97Y74JtPDNwwuApKskxrnxwpdLPXVnKY+eR4OlrQR7bCiGitHxc8Q
ogJVWxN72munI7Fa711v4h8muxzP6SEo9QRb4a99g5aCwluRfJhcbSpMaous1+PK
L5xb1MsrRH7haHPPUuQ2YN4sJvQE0WmKaCjAjoZiHRhYUynbkyTKWaYoY+25wWov
F2jUXgnlznZ5g7+wdRLN1vpA/OXTolk0oNjsPtRGBYzAQP8un5yHCE73iAx8oW3X
6pyXR3w9epxEp8P1dfYOnFDC/75o3r/IuIhxIBFi2vqaW0c8c9jDe0UzF5OWr9ss
a2LAQ7IO00bt9LfLFL/bYl1vu/e5fBYaXo8L8FGj0XZbdxTObepBwuh0akKsiAhg
RRCEYjYB780k5DcNnTT8na0nUJv97CQsda/qX/yupzGhrYXpRPejKPTCDKH0jzoD
h6a3HfnfR0aLVK7v5yC93muUpjHD7PiaPRO6yOsFT3j6uN9GTp5wyCn4Y/9et36V
X9DWLXO2r/QF5zN/G1JPvZe2x6yvbHAEGiMIS40J13hq6RNO/VJFtxjhcS7WaEml
i3NprJwagn8AL2/hvnXHySnolHu9Wwg9eSqSmPV9dYneewwiLznkhAgClvUe0aL9
CCtW7hxNomyJjnwrOkRP54r5kaR0troYLXlu9tXgoutFXLHY+9+DoSA9EYy3uGkQ
Z02PTvKti5yrqZ8Z9OlY/CEUeRWBdcm3LerIw6WrQrPX9EqWZlreIDp6z6D96UFT
bUVUifGXa3U89ifQeT70KDi3uk4hrwow7hlrrx+ZgGBMFXKg4956HrcskNjU/Yjh
AC1Pz9GRj3PvVc9wPpBO60JO3VhozTcN7syu4auuAa2tHUOP1UVjh5I9Rztni6xa
TC+qLAuIflXSJ03IRB2udQRLHBxbzc4hNlDyyiRAokK004yXdG2r0PnAAfMNafDI
GlOseWiaiAZDgOyl5zriCqC80UYF/vmv/QHjSwDcOXWy/C4CJtk6abJexI5XDWyv
8HC21p4Oam+38XdNa2vX/ErnswBJUEZ1djEyh+GiNrXtx26LTRIdsRAW0Rkqhbfs
EcRPtTra7ZzXjICAKADTo2dwqO4oQqEFkyJiBVs8TZGs/9QOuLkfqaLnZbGj4MLD
WEy2QQ7/8g5kjUoc7uszeULGZaKUIv+04b5pA0kBYCS77awCMvAeGa8dbDArrVkm
4f5ooduDi9qVmRuy1o7rzRQE1u0K4BBfR4gUnqhzH8vsrIleg8HQTACkSkA/HSr8
POsK8vi9yzg+HGFtfr04QwdyAg8Rxswiqy/Trqp80EYHAtEn+JT+K43BhZMKcPUL
RLzT3Xb//PAVrGXAGaDdsbKysS7vWJf01+NL+X1X11BPuZfqxybgiJ1K5f6OOujv
i4pMn7Rb56mHkvocXDO2bHFFIFu2lYS9mOWNH2/GIKqOXAttrxvZprmXu3SwRwmC
Hy138LJXJ82OhnOSo6PmEvdS73GM/y+PM1kSEn6j61vHRC3l+pWcZUgp8XDpngHv
HLXRiiEYEzO2KLoUVhixhn+kss3xNZONsh20QfIR9LmEmEzdbJiM+gsFzcjHqO6T
PmBzBbK30sipr1F3HSRUuJH71CSrlaOh2ts1ADC6CBo1oEdeacDMYxRClU/kK5NI
8XmzcfekXqygSe7WHpojjWp1OLlgpFmjq/x6jG+fw+7Yk+2RA3MaWPI4ju2Sje3b
wa351yY45kPF8QVp4pAuKOolRFisqb6lTNnI1rR6kJUTlhkj0EwiTWTi1H+T1+77
iyOuKuKsN6SGQZRCjliNlrutQKrxXd4z2yxTbsN6Ff7u0dqD1ylA9AGVFdIa7kV0
ItnOMBrrpFGPop79dGrT/QnG8Gc1+oixTY2TVa8HZlAPpwimcym9wcojKNbzoulX
fZNIdJtSFigJSf2UzOJrLMhomE1CiBCj3V9BxaoESzMuETP0wQtnVO3QAfE8TQLi
XQIyh2VzE0FU3KBCfK8fJ/Fba1t2D4TW82qauvD1OofWve2c8WKMbv8R2KWbqbT1
vYKg2b8sCwrIMzLWBkfM8mX56le9wrhpbYe8a2Z4CblNCc4pJo2ZSU/2OjvZPF0h
1TrmqIRY2PcYt7wzbyiw51Gc86xcqel6HfWmXUX9fQq07izzI4xuWDVd0gPzgoyr
2cgiCnw8VMceSQ6Y73ax3sQQU+84rza66hgJRqYBjTuYihe0xRf1Ewr4USyKBOjG
8aZkBe8jq8qYHm7jFww3xD+oPGkeK2d69ke7muVLM+MZhuSnKW7tC8gkg8CSUaMx
YG7uqB17ZrkOrdMHyrotbOtH0n+WJ86hnMXDElV5aZqoc5/0AD0dolFFEQE0OKme
lXc253ASdDnsEnMIw1/W0rHvJwzUYU9LXEHZpcT9OlJjxbHwqfRYc14MUQe+1D+1
MosJkzrsYnQzPGaPMn4l3rl0o3+ndDIGG41RQsL8XpWe+Xhv832S0s09xiC7OY+A
4N/Am9U2YebijgJkByQHsncrlKh3CrnDBlpIrFkio5/Yn4o2kCtNvrYeKCAwyO0v
HT2PlLBWKnMSnNUQQ8qQKm5eJeX7yujArPiQf+Cgqm8nt0K2KcYjfpGeuzKMkaXB
7sqUl5D7BThSUyec73DQBlaWq+HK8pqpHJHSFWNav6oNU5fOwK6KnPLbGU4IFQR2
0xi+qxSMuV6Qwkhy8xyZVheR1KI6UK3YKQ+3BTjBsZcFdOuee+MwucY72OHi1ksu
Wnl8AcRcmPMRPP+TZ6XqF9/WlUR3i7C77qI0i0YStlW3eegdiXnvUCPf4457z5Aq
89gCQmQNkQNPqr1iqd0UCaq8qg1w+JbpmJEyp+DWlZs6YVzsezBXoFmiQgtq06xL
UJ+y2PvYIpEVjx4P5MZfiwTc9aQ8jS84XV0PtTpZ2kO7OJK/QfkgbPOv2XsfX+sj
4fFW4sQb6wHOV8yIYjW+I+Q0NSiuS5VvlI6M8tXgwMypsWgOCHaGx6ZcvcAqUpke
kaY9rkkNFXjB1rAWWEpQYeQawvCHZk4Fwp3iJjqLMxj/An8cr4pddVxkwL1KiVTp
sYZeJmLZb5C6ZMG9yMzE0d4wFvgpWvQHqrOu3S3lFlliF6AL8MJgR7HMY3QYv5g+
br2rtQtoq/jP7Z0gUWO/AGnrBagZmiM5nmHCMjWDNhVF/Xesv+rGIubgdBgC4U0j
vVGDOVUdc8bu0wIgqhX8mnTNcUkr7vim3Iz/ZKQuWDts88icqF0rPOEEpfYXkxel
bNCO3PC5HCRC8SdjpI+jmO8Oe0iufDYmHrPGwP+kmcpu7f9yEHGhLh0HUYruoyrm
AKONFMd0sxbbwxJ6kjNDaMdM1UiIvgtpwoI/xi7Bdb3Rmd2BAL3paKszx/lIL6Rg
aU0zmzDOX9DyJfel0bRbljlO9QW+B4y1okjHn3X2pKTifN+tqZ0pEyYI6G2lVEXw
4VTlqjnXlrNUyQE9wFJ7p0ETp+uREcje2uq5yeveytv//0dMcH8nrExvkVl8BNoi
b184lVY/STJnmL6MMeDtCUecVsJm6EK49t097X5zysI3cMpob/yrt6gLGek8qdAE
ztIRf6ZcFJ1Zr2k77jOG+QowBW4cHYyfyp3iTiKHGo7B1bWBxeasfffvVJp4DRlg
Yr7KkbUwkZUKxvpyOSYVJFUbpZgggtHbfI1Y3mVDx8bPLWmcpkbQ2Ec+X/gULyTM
mNPrRNl8HYj2KUR9du9sFOYqHqGFNYPW/h8Cek4jTa7MsD0nQPemw/xTNVHRePLX
S7VeYvaRFp2suBngXCTCrnTs83HxGZLuJth1W4dgloxRh3EkfaX/bk20JIbwxUoY
nhh6IoAtu8/y0VRh5qdxdUjy3FDFRvamsZYFwacAkQoTskpRCUqVJRKiMsGVqjjM
8yGvzGpXmJiBM1IAvbMP87FRxFrrnUR/1DVCjS3cydLzTZh+S8NBZvgrvn+wSttI
MiK6nu6SIZzHoNrfVnnWqGrzMUfeIQPEOpkfVq2W3Kdsy8L/y/MNEAuDYCxmnOQX
npuOjJMJG7u7IMdO2s2K8FkP1rRjHvh3UBu15U6c9tc9iAlozvUKQU1oitIM2mWS
RT57PMZ+UYgRpbFwBcS8lihF86Gb4XksgME/oEht32fkXt7oppdeHZKnnZ0ACpj1
YCbK10/URvNjg2RJVY9FTSflc6Ftew/bNP6XST0zvF/3+ugfT68T+m6/qbYJ1+dh
NuuwbHo+Y6K3EZGXX9J9P1sG5QvSdCRfD4nWJg5Uz8sBGNeRwR1uJ5BzZsa4T86T
G/4i47gmDkZiJHY1vB/f3cqKFPpkUWXXcOU20RugqqoeQLw1LC8cPKUvI8xcCDI9
z3lcKBWlxHX0PU68v2H567tUtVpeEmyAEWhlpb4KEdao/XnodwacnzFFbqDxiog6
8BTZdIjfAw1gTvlIZKGPr25XX/p5oHddVUqWcncevQEqjj/dBJ7Pq/Q6OtIgVvq7
fr5xS0DpJCM5CFg/RFxb3bOGeRX8V4lInyfiJrFq64aqPRG58LMQDuhXAob4H6w+
rn2y9c2+nvhtWl0roKlxobc2KOJ96w/oyGy0XLYO1vr3Ie8KmAAlCJcC8EuDXROZ
n6udPyjtLB/JshfocKGUPtdeg7DZ/hSqbQW7nnz0HYG2Lg5IHlq1OqT0baTlc0FA
/LZlVbgu56EmwQK9PrsgmiqSLlOcNxu6H26KXAERBhjIQ70L3h+PhbBmzQ0eE198
5ps9bRYSWH2RtdvTFsFRbVV8+9oko2pfuo2sI74LNwUMQBEdLnD4ziXFyX35GMeQ
Ty1OFRgCXeWOyJVzoQdM9iiYeIYU5lrlLF2v8+I/UxB5JPj4641LaNGzBBqkM4PT
A9O8qyRMPxO4dVszdm+A7smV80Nfj9cMGaayl2LchKBcfstuFMiwaPoGOrkhzSwd
zPA8m+kUQTrU5henzJb1RiuUTp5wcbYPuFQJ0BCUulautGlckOkZns4sztdtrwEo
gTptfkeZLDzce/0Mi5p4N7REUc97JFQLycp2/oP1h2kqtV16wr7YKS7ygb2+UDW3
VOImrUcjDkM8ILj14UDYu4Ragb+g1V9L0suiTu65XfaM3MzA4rpgDRYKOSJNRk5a
3AxT8xltXsyUEbvBMUtu/n7Jvz3nWJM1dj/v5HotnC3Ta53GzomHp1ftgG5x6+bt
dO6bpmnQN1SdXN9xy66y36vww4X4agcNNRDlDUZrTWsjYm8i+YNkiBL2z1GNsFnP
AvHhNwwOLOD9aYYg4gRPU9Xb2JozRT1FwXp+TMMX1hi3hrUR7DDXrzHogKbN2JkV
ZpSzQQWDYkP+6RXJzJVLnL8QZjBqimKDGf7Lj8/+edlsOtlJXjl+AGOpoOkgI4pe
TlvM0LSXBbxoDjyml8eA5+1z2kLHCNMZ7irrlC4dWmKJgfUct91vkEU0yigoOX42
c+WkrkccDT+754VD1GP+39UrfPjUZ6WPAdA66yUVf+X7GEevRMGIf5V99TKdqe7M
fu57q9QyAT3gdvmlUh9n+PrulkwhtNrAIkJ/nV2/6TKz0s/k4RF+dnxsbHGMvNrM
SAEhy7+SRxhOfuSdj01/Yk9CrYvTG8dZ2Dx2a4/bJTDTLQNmtSg0HopU8GxbmHsd
BndZVnFXtt/nSZRv91yUck1RaI64GE9Ia/uNww43bg8kAjLHChKKCqpsQhN544Nr
d9bXZvxwu9nkK78GFWvHMZ6ZfFjUN/sCZXUsoOAS5LWInIRNYTR3mqAq0irIpi6E
99gHzu+ROpAXMs7YT4rcidSaMFxZVEcUnGaLV0/CIBgzk2IdXFw2Vr0qlozu8hWY
L65/tx18E/GGq6NaQDshwSEzU+2gQIm7Y0ApkfgeJIapbZ7IBP3VD99HRBXAskuL
Uvd7vzPsc2c3HX9Dqrg2Orl9aH7LUroWeG8DnZUhbW++ZRJeAFqt77ADtpaF1ZM+
1bm7cZ7R3BpA21nYJq2uCns0DUQCvGcr3xChBV8jjm/yCLt96BXFkd1St75OLt8l
CbWVwKmEAH3PLgMLdwGQd4OuXP+kx9LRh7NIeuPDFiNTA9yGnczAGWaYUWljN1vy
jvbMuFbl2m25F088pSSikYseIXU6VZTVfBLu7gdbth34p56NINHhGD7oneCAvJef
xV8UF3aYkgDEe+87fa5+JIViuCadAuOKastI3nZmTcx+X5eQuX0hKnh66oeu1PeA
FRbRwT/NgyVWb0Nda5zEc9iAwOo21mnfeHw5l4NdQ2WmHlhtuuHI+T7qB/GmGbu1
kbxKLKWIYemTw+EPoeL1shb+GL+VlShFnepZWfKWDWDqcZyAFyeW8RDq8dOIQLKq
XB3zGCg5K5fcjQoRnmzVWZP3Ytd14jmxE3QmRaXwS4+Utj9FAjNO4CTWHgn67d1X
VykdDj9sbN/0S0pgMzEzXW+CVMrZHk+Ni7Rm2kaqR+Eo9IMHyUi54ZfkB51T7TxX
otFXsxWxGXQ9uCxr9fexUykvn61kqBq6Yg2REtpmQrpdY+nClLWulXTjroONWdNh
kEx8iWztRFghpkZSyt8KA5aP8OcZ27yxhcyDhBC5BvCi5Gv8UcstlnPhD5hfIMYh
og9lwViVGzISKpJk+MptLGHoXHesldvvKSplOv/MkXqTRMHrQO7pULo/Zir/6g38
3c4cMkp9ZUfFkbFg6OpSqCDXatnoWLV/T59EzHmky3m/0ujVKnDKM9AnMKaz+/0P
8QqW+PRgIW/YXMts0tBB/KlZKBX+Vde+kbsu6SzBhZsh229N141ETggvUvI1JtPh
fexFCQRX+Cuw+l4qP4JG7F+TidBgH3tnI2BeK2hCn+1HN/6H+sfVyYERxv5kIM9T
gQ9IE4LMywFP162r2eRaangtDh3lem4AM1qzWS5ioj63tEfyaG8XwjrfAfrv/2uK
UIJ1kJ1AE23kXRdg0ezZWvrFyh3Go2ra7Q1+scvx9e7BFQ7mmU4tIYCSgjtnKCOK
Y201a9upWo9TpSCgStqadMD9wJpCi+8o2Prr9BE7vIE2Q68oiv5+OBci5/a5b4pI
FHNIWWx2+18eDS+M03Yn9UG8YCDf5B1gBHo/YO4y1eEVWF0I1ZwRE50kr37QaCiU
mXBcw7Pvlt+YNHvL0YYawq9MBly0tmhXTo/ANKEXenNuPFAbUFDB3Lk7Mr1nm1cI
zYCKL2FGRhvSXf/J93AzuJG4gIJh3qnLgg7JdaqOuwfx62oX2ztYmyp1n3fJo68Q
+tqvlaCqm8ZqVYrZehW/7RWEslMd8XCD+RTArPXBwwakztPGXdyzRzLRQQcxS3q7
1JqX/hexECjgvvF9JmZ9MAi+THKWgjt3HyHbNiDUjjCC53pDc7GHvfV7dXLNVcrw
1jkRUhNrcq+rGptPZvaSd1fJM2nrO9YITZ1eDHlTPo97zdrD4S/jSm6NymeNUcUz
jTngRoFd9kz4TGiQbGLJeuJyR3qRzB1rHcBLvB8wJJjvDxhh3Sp3GJu7cMyxIsmA
W2eUwZzUxe2hs6iuB8y1XNeTyyw8XNWO/A3xSdpxnpZtwQjyv4FlYjfnEffx9h8k
8HxnRpYZ5kYsuFRvWRaVFK8zcM4oiTdOp263IB9jVt5QuIPedth/Iid36iRCGlTC
ZwwqtxxomeTCKoBaI6Y40WMzVghQ/z+j+IR0YbJXMO5uiudm5qEFua27SuF61xRG
ss43bOIiNIRyNclXWrnrEDnZlVHvtsZ6+HiNyALS1am39TcO9nxWRzWXTS4pQ3Cy
ARHsmWt0fCk2XZQPcaI+ji5wcZtkXbJnx9bewwmzgwv/hA2FkSfCK8peWZlaygA+
XBzmA9f+CpAtInjHjKvJFsSNuJzodGiyJXeGdrL4788bZe/n5td/MBhtfO/rjkWC
R4Jzisyr9iyeDK3Z+gJqwAvyMsxUKSq6AKwAQQgQOP9BpRRV6N5JX0up6D75PJgg
m/t96ufM7Wizf1Mdwf8V/SVGuAo6M3IHVQizllbYILCdTLTo6mRcx9uhRiel2EsD
QcAKs3eVkPDnU5v3xbYJSpuk7UMHK5E+2iP0aDz8VTYbdbCs4aBXRLgkWa7agr08
yS9bWmAP0k0rYoaN8UljRgzdeZCf/UQW9fgx+TyMJbi8vWGgFDGqFS9iJh8TKr9v
xICtyHscfdMpGuZEUcsuPZ+vDcUbIr2kuqxem6O/O4vcX4RfQ4bAP61Hu/kkDjaz
uF8zNIvOmIcC/IoyC38frshnMJZMpTe74/mrjfQvbvHPlZmPM4j5drEoGyarSRhp
strUVa/LB2wBpwgjK3prp2swy1ZxWlHbLPFzGi14W/QXvkniG+R08+Ftc+PwbgG1
8NzwvZUBzsXdvgmjlJG9yNRB/3uP/qN6KSERjUb6g6+WsFNIaoNJZ329Vklz10Zn
LwrWnxv+gNuUrILA7mK4FLmTBPxzKX6wrSxT6x1uojftqGHNjnjnOwsCo9B/GsSN
FnIekSy29xlBfGeYe+M8WBINk6mU0KKoJ+XpWBayXtaEEUyjk3T69zFMxlhzDoc9
LqUEJ5xbDrUl8K1XzaEzY1MTmZRAr6MWxSJzF03kEZD0FBk76mNUJTtMt6perH26
6aVVNE5SxGYCUPbzeiMCVZ5nN6vnFDLlMwZwHThzbTIGA3U7oiKA1oI34O2h7GUT
frrgCXLSguTBK3RwkKSd45aNractl3CkN/a7QVI1u3TzfW3C4Hy3dwM7Ugl3CJCi
fmNubS+ocR+Y3IF1tEyvms/816KChZTTQIDCHpRqdOaeN0Klnevi/lD/FfvWddcq
23vuzpCqaBtrp+Ait0D7m0QpXV9vIvhBAd6iL92n8Oxtxm+JMBRkZIswhYa7VN3z
0r1npMcNRZ3L307EmxG+M32Mmr1Sp11wzotb2OYR+1O6r3lW8es9QttSbYxkYLnK
qUfZEZ7r0EcO+y2B7jAGzIQj6+ZRlh1c6HAQkYuWWrvqJo1j4hqkGAmSpHj+/Uga
ytVWRKQ7xWj3l0Qa/P/3oBDAN7wiflQyZmpsVUjzfCWOx15bLGgZ8hilNza2yUcX
vyqSkp4zxrisUj/nYKx/8z2bSZW1EwBk+8e8Munzudm9fBHQ7YL7t4mVNBNNr2DC
U5qdzHn4ud3821KwQeHRvfpFluVdO2auwQxN0Rpu0kzMh5RgBLhRvnV04aeYQvyO
GP9m5DxVYVvRdClT6fra1cHD1XsqGcfFLhyPmfFa5ywPLyiyoh2wjHIL5gvnTTkp
e5OGpss40QH5aPzMhDDVXS8Og/ZlLL/qIC3M6wSt5f1Au0wxI97R7iiVXvl6mAn5
N23HdJseSZywZiXbPxn3a8BqR/D2+zR9r8zAPkZ084Y9Or7yCJzBzgJasfzBTdsl
r0Ntv4F+WXyt0lrcB/gdmJkcG1+rEkMuB9U1ZMin8AHdafaDTHeHZncOeujOuFab
i3JzpsYYCdWfE5FYO8IIqstL3/ekU7ZXbmzELG2aSe7oSdaTT/SCIFFJJcvEjqiL
VgMz7jrNMzbtMOod/Ge8/m6N45+Qc7dJDrL9uZjoDwFL/faonbU7dAs+UrARzBlw
aBRozMc5LKnN3yBz5XXPVzKZyjbU1EAR1vsJ7WRiarp+JpDkzjfGu3yFV++IC8ul
o6JEVD+w6lEObnCjr/vyg71wIxgBYFOdGYJH8QtFSx5zaFZVJ/BJcgJAAU930l0F
E4YQSDiOCX+w7E/Mn2sWnpapen2ZmanePnJJ+ZICjBRKbAPgA/Of5gK0HMjl7HEq
8DwnqbZRwyrb2ZirdKcS/7bd0fNyr9VeW0WRp72zuAJDax2YfLfh1MxbZiv0LS4l
f7I7+jr8OiDzP2WrRHN52u8PvAkBb9CKAQsLmc8+BJF9ZQo3KUQBcUhKjf5Jo2uO
XtLInejdiMw27RrPkR0MrQHzgS+riZuD2Tv7/OTLZMJEKOCI+U0WOsz63VywrUrO
sqUv2UjoQ6S4d1q6XWDyswlV1qfJ9Lhb84/T4VPXA2lJ4SstyOK48oT7gE3e37kW
dQuI+zbA3bAD1hjCSkKDcjJmKH38Hu+0qGHkDg8v3I7qMIMFH9gSsQZZDwV6/eJW
hq3sMSDT4TnfrDcxBCwePrYATi9ba8da/E5gbzDtxvHUXRYqlDxHLTqPrJ+9gM2S
VQ4ip6XhRFcRuihUazlJkigaps70ZVMpC21rzQSFDdkiV3EuvT9Z5orapwYqEKdx
yWlmz+7F4Fd41L873aRDapw628jugNAFD6NeB2bZamSFMAtsErf4PJgUPfebI8qF
zGgutns+FDIEPryXwnhH+cAX3HXSv3CmkAuUoidlX9A5pgpI9D2sjfU0NCdoDduu
E6VXtrjU3iryz9QaPRy7pRdv/2ottWQXeg2DRjWUXPTx/r+s6hLJ5MOHZwW54o6M
sJN0ZajbDkpoFGrzomU9RKNLBOLOzoRdJfcqGydJLMDt48k/tpggACho3HHUydfV
mFzp8M+QN6bv6fNJlLb/Jjm7EUd0BFme7fU8IgDGAwS8th7ngssKPq5PKlikxGCs
BX/KotC9TeOfeAQu8kMHK/L/cZD0KT1qADaVFw4+qp1rhTD4ujBokxv0Fo4ZqqAI
lcROqKm2S1gLmf1Y9qyYIiDIm2rzldkj8SvSW8rs5Q3hbBluMVKp613mbi0VNw8L
DL607vzTCWzgrSrVxfKKDu2+7adSGSoKPEBldPQs9TvvA4c8nMMCMqn4yGYsto5a
aeyvEqdY5nqFr8U6P5hw/lWUlsh2Lkz4REWOf2ZHPHDFOCjivjy49HQV08EfULvM
o7T/dys7gCCpL8Z78V2EpBMMA7f9YVtJ5hqwbzriW8oQvyiVbeKMDLq2LGLfkTwL
KC/teMRiJ2AoZomFc+8B2UXyhoHhm63QxVotyr7oL/T6bt9kQ5zjwdVOgBfYFzR5
F5YiuuLnhWl5btW3izF8JX8TQiAo1g/9M0LjZNUtXfg2IzIaC2bkG4InCT7bNHSb
NxBfUOSo+qevhq2NeDgGbpgF5/QQQ2ZgMnaOag7lyhrpLS8jof88+eweK2aRkHcf
lb0ZVMXpp3MCKC01TGaNMQmESjbM0pZWSX+Zsi7VtDCJaanEagyJadEtqfviC55e
qiNyCztbXm+BAbxL17TjNo9gyczBHORnj1sA8oJb+Gs+0u4gjYCwmaSGCYOJAuAl
CCo6wIDpOzB5gcn23hvyd0Qs3d5BrSLRM+EPW5h/CAdmXjrvefEQQYKMwQ4+Sobq
3+Qrgw+5vjTw2vazJSSukPlln2Zf1rhPs3Ic0OgZBuwzP/xdjU7XJR6UtKFg3vX0
csL8/u/TvO3vPm4hzbh7KhVW9Us0xCo+RrXEdTb2aBYOZdCS+IIHrJBIKSRFGB2g
62wqhZXjsT4BzcedwVvxieoqx7n0nuRdltP9HbWvuwnUAB1gSiDIXG6GRODEmmA3
lqphF44KJ20Qrgt3KDDRVOIDgTMeoaWob6JrinkZB0iHEvae5ofgJCtyqX3AQEDp
c3m/3hosmlWRroBBL1sRwwo2NJkQAQw425M6BDqSnM9zC0RYeRtZDy0xfXhKGJx+
ovk+LBEiXSf2d0H8sLwUli0a7+kOtfcA+RcNPF6NQFftLCWEP3ugmNXvFBgHrv/h
XgKMHDcyxbAb+hSusMZ8R6eXhJ9K0zgZS8B9nJvPtxrUtJni+NfCPEg5JeqNT4DK
ZTkkMNo5gI4j5CLjikw60T1uU8/BeZIpGgFaFJ9/oiIMwhRgd/O7P1c1+cYKiHtg
JYbGLyCjIHejQRcVrbdLSKwUsoXgDVWMv1M6atfOFGtBWmRR1odRs+LWQR9k3bie
Iykf5PtqkPveNG2b2WgB7rmd7Lx/PLfl6fwHTuT38IE8J2gt2EYEGTtkPS8vU3SE
5GLKWlLUDliKsBnM55xuo2RSvtvAAyICgPIqJQO7O/idFCjCEhC+tZjM/nLjkNVh
GzPggqabLOeP59CpWmpdDVqEb/O3v6Pg0TwwE9p+WjZHzrnzqCZHG5ftTu3F0TTG
lrV4dAm1efemjAeV5YXVVr7004n1c+lMovTTVc1fcpWL/lkMGPpKCl3jfCihIya7
7dc+cw3kFGZfbWQPZGhEcCSHzJF+IOSjZnRzDHfJYBMbP8bc2AXTMEV07SgC/l3s
3qJKEAZVrgKITVkvZDj6hya24VsxxtA/E9rABKSLpFk1Tn5L82JBV+KmbblRmbnB
d0jO2iQxkq3cFOaxXcHvArValooSpBbF2qGMjDJdES00Kjd9zDe34SknGBuxKMdD
295y26IaFqCTDSwLgy9GY+tBJqoAA0I3txoEieX5FmmpX3NFWwbnEJL8E19NqmwE
UDfyj1191RAz0Hf+JTov4zMcxbrsNLOuuq+g+CxSVgI4FiCTaQl9Ikml2s+Q14Yv
3HNmEdeEHbGVe3ZZ6iC7gj9EMH5NvX29fNDtPiXwQswI9ydnjr0S9zD6yV2B3/sf
9tlGCF/PNVWQ3ER9PYX1QpwWjKp00S9Q8TKnvq8qt/pmmNveWrrnh7BqFhI6MkJ7
ciGiKmRPbNqlWOHjpW+49q3ibFQL+0fyT+JgvZZLMjkFEygjK1SKAICad8kB4eHo
8iz0+i0kQscdqWtFJYuV0kf5G5d1us4Xr4UrRFD8BGpb14GEr+LtTULYjGWI0BFa
1ObRK7LV9Gh5Gyqh4/2ckVHfZ3q0vpx3OIDgPGFRwgYg3qLkjq409gUDMxli3ejd
YxOKPF2WbwoZXnIbyo/TcT+nT72sVUgbAcgIeM0ZM4Rrw+JgvCZXrDclO5/Sgzho
d7UuybH/Zm32+1H/Pd8Tj/I+1RVzzFwY2o6YK6qAry5BMNUV+nyVfT5veoD6Suww
EqwsuvPNOOjEtPuXLRWbCPnuxTGvpqjQYV7IVSYwFftpsHhMd72xgzCDbdbYTFqD
PIvqNPlmG7l/mWKh5XVZUom6ovyWzvhI+Zgm3MVs04kxBRIjaedpNZiA+1+JjX60
HEnqUP+AIfsDjqugBJndIEf3FecLMeWush4qzYPwkfpz140R5lFwC2E/F+fbiznC
8Gggm/EUtJMhNZQ3Fa+5tKI7z9UfAQ2ofbqRYL8dNMJoKdIUijjE8E1wKTo3QiMa
GvxBzsBQl3HTt7d/CrjGpP45tBXI1eHlvWMkG86ImfUDOkVIb6jVCxgPR8hAH+qR
pZHKN9opnt06oQtfwEbkZ+JbzzGtHraQtZfrp44EBM70OBCc+AFp3TTJ4nprm+1G
rptR++PR1OnBFNA9qgUZi2k+9PVeMmL2oibH0L+htuf5InE0edEYUZXk1OQUFGzt
6OpKE/7roVkWcoT+3yyZxEAQDKRW9oeRxbj25N21D3h5IWmPHkK+1AK1DSqi4b9T
ZMctaAmDtPuHKSHXenuLfc7ip3Bz8PTlWsngVhdxCbFBsQEK3b+dEfcTgaBIMuVr
CWFoxSGOl2oEKEjINvZFSx9XTylQKHqoOQg+wYGrEqAbxJ8dEpiBTWiICg5YhisL
QqzO6nTJdHsu6fy7UOMdijZOxZ5x5rt/5JpRw+gZAQCT9B8uz+F8UQ7wc1FDyoy/
0nimVyHiXNKqEZ1S3GQasMPPzB+db42WE/YIbH6CpmUd4jYTFrwOOT39gUlR6aYo
mUC5BBaDqU3ozDtl4xR0+KAH1B4EZd8in83cvf+dVnLXknk8Yn9LJ9j5gvXLj27I
R+L5mYKHzIWqJgHOD/yQBAXooIL3gcdbFsPJ7caA02KebAwxZIumS2BVeiQLiLlg
d8GzYZgxuRRLic72IYR+gsIVYYqU6/9qsZCk4YmZymoCl2KhLbGImygFPR7oigOx
WFHlD7/fSK4qPJ6aY6meDIaSUXCSPz8DnZ8jkTuv0Ofkui1Eik3I3Ps1FqdsVRWA
PaMJZyW+rDpjohcTvOfwErQfnBSZnnhjbrmK9k7sd5GZJiJVADo6CpTjJISMoGdx
aDTAGHsTO04RPVJUznE5dFV5J+X88P+kym/6SLiwWKkKQBuLdugiUD5AuYtdtk6c
CJgdg8XSxOyeSKnXQqMeU2ycZNpDgO95Tn7hOpIYX+YOyP4hFGP++uBGBINMExFe
we8OPEbeEfMCYMyJaSZXNyakyExd79mIf9xC5zfF8tOhUzDU2Bg7QWRIS/BLJLBa
eYoXDFZnxCQsTGxI0SpCgQI1hymRHahtot6yNT30YmNekEC0joIzK3+WC8f7XPhs
vENXp8IN4Hj3QcfIFzdfn2+NVk+nKYH0R9fLOa3DF7L8HgdRSSIxDg4n/vzfMV3f
E1FT32IGCg+9a/NyAdf6RKmz3EpYPASb+EKYDlhfP3FEQ7ugy+M1GKoYXgnCFEXn
WIhuoUZKVFY3RFh0gBp4zBxz+pfay5kqntuvkwGMySij84SFPTGk4GAMQCa9xWCS
4qN+hKudw8xuiWZKwJQXBOc6kgVFbn33UJa8vxCYz0MT8EJDdL/3GfcZacEm/reR
xufGOaIK7dES4McEbu+PSisz3akRg6kf4E11pDXM3FPtw8TtL1UOgWbwON3LsbmB
6Hh11bp8RiLVPKQluyipCwy5NHc8t7zmwdUmmXETBCldqU4mSc95HaBSiaJ183sH
x8uXiKiDckjPRJCP9GTqtR0UGTT4SwRf0A8pbSUWurttFYC6d2Ag4C67n9OjBnDx
d1c6GrM5E22k/aZ3U37LyKTQoD8eOsWTWnFE0+wDz+Jmcxob4e8pHkJyyQgU+Gc8
Uc5Cei2ZjMs3Fl272tblMy+uCYM8wTOVu2HpJVRvikqgSsMD4h5FjkEeXDajC/nr
15OhqHcag/tGjCjXeS7qUUq0FhxhZwSF7uVNm946SuWk/+AT/dtNkB5STJQMbl+u
B3J8s44dHustMo5GqjhoBOSWPKsepu5T+Pk42Zduuo8ERxLHO/PLTbxPYo/Ijzge
0Ou3H4Fd67qUsY/bCANMEnhzlH2sbt6lWSetrk0gm6FUDNfkjRQkT7Jz9wPU6P7D
3/yswBXQm0pBfZJhETq1TWYEvrsp8KUHS+E8ZbQJdbwjYppohEbxY2i18Y48E1aJ
ng/18qccHJMYyfdxfR1snQXidsxxH6Zxu5F/pJI3FyWizKi3qCAyeKXl2qkE6AM9
B5frUrnASFQ4HtFM0Igt2JLbgab+k9reSR76ds4XDm3/jJd1t6UZOCcYvpZ3+qJy
BUVfEpD9NDxTWRYqEy0hC17hAzXJ66wCcnNYuSddMDscFoPXskUUiYkM/8J4mmmW
UqgkOd++LPpBR+tbeBmBY8DLzV9kFJjysrQGlNGiGSQKCZjCT+BJrZfJ8pkc6inU
QC6IfEGLD33OwFiWsKOBncCTv0S2YiTo9NQDCBYNl0dxpRbtFUPIQA/RCC3iVs4j
sZtuNUSEYUJPRwjr/MH9jPTvM+VgTTD/9SgxzjXzVLoXPIItrN0T7vqKy1QCI6S8
SKq/Itt716u0+yTyJVCoiKSRNOLfGGve++ayhQe9EsLED/bNDUOWXDSSVYRfaGcU
tKHxYqZx+1948NlnlXz7QmHh9bbBrghzlUd8VUw+gitGNsylUC+jA2uVO3rRAYsX
cRjzPAskLD13PUCbJ68JcZtjpR2cipU0LwYRk8YCAEghebGO2trX7/+xxevdFmcq
1HwAkBq/5OijiScLGVJP4gVxnCjzlQpEWXZNBtwCKwtZEnh3htD5lXuZmBTX7ILC
aoWzbMdPkUXA6ZeZ2XKMPh+kfGZtv2zhpmi1vQ7qp1rOjdmWDy9sJqpEpSjP1H9L
LnrhCfqSKMqKTY9MSq9jpz1SNEIFDjRA12PbTkj+DW5gT+/B2fmBVkDZ/hRZaHmH
01fqYVMG2ydLskBDHTq13cqaQQFi75V/EcwCXeikMmr6gnUChI8YFACPwY3iWRyX
MWrK45yn3/WD4i68TJOJFli+vjCRVyLe6k48KQvE0jWhrNbMc1cFXfFqoKPOTRwS
Vpm5f7qD7EZgUShYaZaHKPKwztO6zVq58R+p2Pf5C+57ZxEdJFhw1BPga4JqGcO9
7tPMqeY4TUGhi1uTXWGbHtuS0fvta0L3biu9nSg1YgaNDeViVDaTUCoktI8+uRKz
Xd2LKmYi8Um9IaL3KyCe4VUZ3goVBu83Sy7UPdCVsgLuPPIwPeEBoxZf+qIedr2R
7nTW4MzTkgE/YzVfYHQBXs7he4Ii7E35gcXQ8Vke+hHRyjZ6MaRLI5j8xf0atueB
FIZvntqB7+wqcaobClp744192nryHNW+ZmKZL4VtAsQsr0GMEmZ9s6YGnXL46yBr
I5Zh/UfVlY7GB2u4XDptodkfHVCNM5io6y7VdWj/zXBQB1u3Zl/BmNccLk+QKhvU
PEmMBMByXfVR9smFz9q3b81fBr9xcMSzxMR25ebUklU9aW9F09OUEA+VlVbayn0C
NvzT91wwLdx9GZND4VjiCWIvLuQrotd0ynLRigxR2WljkqjOaFUQa+niYKS7yHvl
cP8yWADSeD1zLriA36MPlzqS9QMgNCOkyLM5o6rP4c1uRhHelRdvQqLiRbhRS7sz
FyYNxlFQl0j+CvIm/mr/TE/M0rVV8XcD1ZQ/XBHb5S08JWqGrEacwKfq3GyEtLxR
efIn+07YdWfjle84igmHGgo0ideWHy5XL7wm7KrswcwbaylQUtLehWcK2sfxQZwH
mlgRCzDumfBeLeWkjh/bqLNkKgqVIptRksrjwb9fRnkxPP91ogfQCiYXaGxuhg3r
4Y17gwY7hg2yuoq6ox/WZk8EC48kJ0qeCYRw/fbErJMQ38OjwzWcf4A7FrRc83MR
cDYX/nlW8GPEGyLdeoUMj7e7NEZaAkTRRJ2wj4Y1nPwERj2GyRE6PDqU7+72vRZ8
6Zv5WAoAbtJJ9wCJgcpr4OX5lgKNh5L2urhx5xOIH8l1NqOWS2IKdZKXoOLxPQZ2
5vLEL43J06KX9ySurlicPTVWw5PxudPqysXnbg+K9L8f3YTx+0ZxRBjUYt1eOo0U
J89AVJ+oDfpaK1DSMvXVa/VLY9N5429vswdLQsHbx8NAhwzIel68PSBW/VBkir+0
AvC5lS8jv98Wz6c2bAA+ugRUnc5w2VoQd05X1qff/3tKdoU/VbMGMUjfn2gKJ+Dk
QfNk7TouZD5ZV94pmZR9QpHP7jkWWQdnpS7CDOw4fUvDaq462e8qs6R7+jieSRZq
6rME9+VtLcGG8I5qVvimX/JFECTx6BvWAwFUjElNXMxVo0A5mfHFheYeWqMzGsxS
ngkwE4auCChYxttf5CCxo589HLbo8XJEFhGjQJbXtgzMLYa5zQilg7rrHX3XkO1S
9vBBdXePuPqfXaqvuK8TuEQtSwPzgxZ/Nb6bXZMZJHfHt0/rpamYaBcBgqgqICNx
Ojt2q1pkdJP/VqBx40snElJI3OiYg44jgpvB8odgen7jCzscaekTxT9FADd9esSx
hGhKdjJN6yq2GySXTEbtVTPva3tnzpDRCuQlG/w90/r99Uk1RXdpeSAD1z6QxOeV
RBsgIASqlvmK5lMv5EZ9P9PXF093x6e72uJO7yx7/6Ael6XDTkVy62NuPfraSHZ5
6EO5ISLphvsZZ8htkPkEOeRhwqGnBi0ROLCcgXbn3Yg6uJuJY1jWEfYuRAN40FdT
47czKptuIhsMHZmY7yiUF7cMw80vqXE7EtZhb32ZR4XV2Y9z8HRzReREj/ghBwF3
gur4Fz8qQtuT3md9M3qNOd6LDs8KxfTdyetOoCTHy2Naf0IBSuoskAaDofo374cZ
hrySda4z6HxD6Jokz33WAJSdTLixq5cpwDIOmwvjXz6m2JOzNMmulzrZ2+j0FS01
obdIVvwSOC50j+8Tm8MzGbVw3sM5Xzk00mvi+gexGUHNfmzgjBI9uvAJaASGb9N/
jkHWNflGWYp9JXc5v+3VQvb4hOIuVLzUTN4J6QgANuBQNTsVUoaRnhstgUdz8DGq
XXdHO3q77gix+phc2O65+tQfCp7/EWATQqX4kEO5xZtLWQNWVAEoJmd2p2DUrR5a
PRKQBZP6Uo43bzQbStxtaj9HQtbJlLo9X8rSx2i7VWRY9YxmX2LEPemIVH4UgqIi
sj3k5iVlM3OjbqsOsIjhufyplMmybPjyX1lQaHE9U0A6wMImJ1M6iQU8MQp25m1Z
j0fwzoUUzykf9cbS5blnXHXYu7N+XtfeTCSiwF6lYEA2/HECHuL9au7Cet6FXD9j
rIyWZco/zi3DN9qMKZXtPv6f7PqbIdBtepMTPr9JZJX74QJTnSvZK/ExJC6MeG46
ZNOt/G6q0rE6flpVof37M+5cryE0TWcJPECfZLtk1i31lEYcWGFEZWgfsBF3UsVK
LsQ6S15Db/vx9j8PefvCIZ0gPx9OkvxgWXKfyFrcHM8H6Oz0Zz3ZedtGpamH0Ovs
KNAKwOimbOCvrL7khUxIzd6eaYeJhWKef+iUL5wXSyWJGTc8A1aF01gtplj0iAWt
aSOCVMjMXD+5WeFWLRjdW6Eion+VBdfowdYP4ylkwtQ9NcFl43VJr+XhO3Qb+Jn0
nEoXNET0UKHEEamJ+MsLD+ATQ8IwXOWr9lxoHlaTACfBOGSj0jOZgUSibqHMYZxX
oJ+jE0TkuLxGij192mi6ZOvUekEf26VYRBNg8I+FbFGVJ6BfUMKgFzyov2xQ2xIb
2/WTUP1eWUrKNgvjEm2IK4HHnwRVcFPRlL0TnuGYiuJ03FEkV9CzBqtsfF40fJ0L
aoBuZR5umVFu6mMfeSSsu8778pvDe1+BFFceNFZTTjAgC/cdZzl4+rKSZSwKgR5H
qYCP5BNJZd1FvkSiwyOELPpUqXQigPyAC/wf9Q/76XVRS8S3FefQZblVjewu5oZP
O1c4MKd0RaEhyTcmulHlqBcJdnfwCBH+3+jv4vRTJ4aOfARKNeTurHFd2/JiP5CD
gN1d6YDWiwn/XUJIiUHCCR8XYqJDhHDrYglZx2I3R34Y3wfUgMdL0gROyuIp7pFZ
8t9bfO0Wjx/vEEZE6I4uhif+qECXsVXAmRp3L0gOhCq76FCzLxVFk5PF+rttGkgG
N7dhIKzbk5MMyqNp3+B3XklSfXxFLkUe1xzmAMHlBrJYFBbE4eRM+Eyxqiuxs7d/
Pp3SeyNopgjPPYs99UQFX88ksBFjGwdN0b8BCzi7YwyJVF9tymk4xl4Q3+Dgx2HK
CqBrTRoWIyQl0u8JxdTcDfK9C35AOQK5qirx37pGCFOzDQYwXY93sUH+jdGzhBiN
0DBMXzaYVBlir8T96cnT3yuJnlIYJuV/JDdG9toB1wJi0B/Yzd2xBHFD88zpSnTu
hWDlYBj1xv5F99gC3Z0bJ+gCg6m5R53QwvhQ95oLF34iOYrxta4QRRBxfNVGR2rT
OS8Wq9kpD6kK9a9trD2Vyb78DIlPVMcnkWM+EQJQP2eWLYIdZyYsW+J8+3AeS1V3
Vd8bLBJu4ObcePA9INu+tYl0dwyEfsr3K6kIp4TlYd/537JiKzny0qO48gijo02I
//YRbQoxb0mOBSguo1qjwapqiw2sc3ERJG3lPUzU3FGWS11VE8AOZR3n6nl5eMRv
aopas0tBR2pW545X63v6489Z0Wlu202ryHAMVa3LUMgvLSlROQAapvnp6ILsLXvR
liK2byBIZrPISNwKFlymPvNcRacqu3+lc7uOffFIktg0revVTjVelsUsjsb37Y/Q
kFkmUdGBNwq3IBug2ls3U0IFM7oov76yGdJmVPKXqA6qQWTE/uF/CuuBETb4ax5G
DxzUz/GzJOrgkQtrxO4RNKExewjFx0c3WioZkWuDaUdE8vEdSdvz4xg8Y3CRprZC
/gztVc0ly24+kDE5QulV5VUqKCD6rU1Ndy4jYz9+LHIEQa9p3ZBn5OmSsUPXSPYk
8wYOiA1CV23EKn4dBAGGeRz69IXxsycJp+NYUUwJK7AMFYsITLFz6tc+go8F/N3l
/ababyBLEKapjjfzwmLu4Qw0Ki2SzeAZcL0jURvdxW/6/1VUXUb3aoFP60dcHDHb
tsLkshSgPMRg85uQMIawzafGa6rmpO9Ywe7yqEfZj70xNuaMH0mQT1a2mGDxTbeA
hp+r8gTwAyjLPrBl0UeGXy4gPZ5ZLBcWqvgs7UNM+TGGLIVHkZrXxypWMmcooe9N
vtcqALXqKzEG+xL2/Nqrx0Qi7dWu8YHLUw3TJ9UKwRly2tktTe3Zs3YBKhyBvWZh
qR5GcMLmP24lQel/NlUT31h6J3rR0HqzwEfyUFbK9BCrlKAei6eQmJqpDI/CtITY
b+QvKiYzlMWwNHc5fdVSG7+N6ZpXh+ZoGOJW6NKGeG2Ig2CksLfHoOYVIrmzYfSd
mfWqPRp3h87Uf8MdVydWiKYIdKN3wIcdf8ZAgAsgJMl9yZVi4RSUKN8HhkP0FgVB
lC3ko+SbGbNbIDC1Tn2luEL8mxSTEBaAAVLQ25K3Ls/BFMWfIMH8g2laR812Agcj
hT99cMQonR9GynTqlaEGQpoaCBgfmwANPDROLJCBcRTWE7myaE0WPkyf+r8ZvooU
8oZLbQ9IexZ3DOgmH0dsNnRNQ7Lu7Mv+m9S8rRpciacfCc/DNR4jXxjWFSfwiG4r
tX1T4yAZPZsfvli9Xq6Nq5qe1Z0CzgDZJCqV5uZczlMNKOozn1jWfKyMCHy4YSfX
TUqQj2+OYXYKiFG/RvJH4XkGi0ht11pqIBBKRRmK/44PyvSlZmpBM5aw5GVj5k0X
tqNaJOlqzZGENvRvMFyMlTOZioQp//H3VsATmTZuX7vuO8p1XkPgwRxVIYjW011C
fhhR8tqjvl9a4BwGL1atjt2j+yh3pnRqLYe7LrYQtenDO+7fcAVGjPTzdFoZPfmE
hijGTTVgizdwAXj64a4knnQqDw+zeghZQbcuBvZ8/bF7JgoivgZseccFYHiK5FPv
X39NdjkXus3RGuGSnEkDCEh16x+PC+yj6xr9HQC36EnrUyNb4VmTR3iePPCouZPg
5DCZu1ELLTnxRfwslX86gL6iRgnBPr67t2NLTICKuvi8dhK1EggyEuRCQAvzveUG
ilz588dWpumBf9dfX708aDcULlQBoxv7mPQJL8y8PfTDxb7RBfRQbjGIxssUUnad
QZS6bFOcAMZCcfgU/fIC1kM/HeIEz3nh9HS5xUyK+OpKWbUCcpX94RT0yno/d32b
CifauQ0yr+t0BWWv8xVzggplVXtetn3dmuQqBlCkd01TnchRaO6NkDVcdaQDLFeF
BNf6uL2p/7KBXTP3We1sFH3+Q7GWBHO/BGo+J3sjNIZ5ryh+pXLyHSorXPu8Ur42
q9WT2hYBiIjY7Z5LP/fimL1kIe8bYREqBI3zzxrlL0BciJfroBUUjTSzoqd7KpkF
7ASbvB/0gql/zhqXvQWj8FWyDH7IPAiFTv9hIVrbnGoMYtrmr7GGQDwfihZL03qP
DZqcuO1FUZeAKVcV8K8Mj82IHFvGRRSlsCYIHhPTSd5FXaAZnOEstIk3WbyiiNBy
PH7nWyX5zZvC3WAttQj9XISOv2jlFsZhTwY0rOMNraB8Yirii2Rv2J9ezwSamHxB
uDAc90O2cA391X1YsUsz+NHVbSw9nvRkmRtTScytD5oQCh5L8z/M9bzZg4DYmBCj
samA9M7VXAPZbIZpcQOJzNWdyegBuAcIQm2bVuWnnh72krne/itS+ts2BvDGWG6f
cDMqez7kZYzbJxIhBdwIZu6ErULtbrYrpcN+/Qoq0Xh1/VORgV8hwAxCGz1cANwk
W2fFnNRLeKhYy1KvNLpla8OkkZzLzGSe7jQVt9jRdgusuitr28tZ2YJ0hWHlecrN
nV/ohr0QYj+i5vmTw6I7+zv2QSBm9UUw3jMWbfZGhcSExIM917ZqSxIQzoVnxXla
n5hdyjE1jX6VFmfepR36O7l9EY5O4zo6QrfhG1Zs9hqBACV2LbZP+sEqQ3M6HhvV
iAUB7unSTwbcVnA89ybRf450pNpT66VLrALJOnDWsLPtNOiakFTJu2kJNz+wEdXt
h+gx0RBStht40rerzZYJUimshvm2SrrJ73VP2bslPGXbMx0CB6S5MJuhxYq9e/xo
0cic8aufTdyPZXvMlnee6j74AuEDyNXXdvPF5hYT6KLmcrj3sWZC46AAH/0/SL5D
YO7nhYV32KCLSBWCUAcjm9ijSmjl1VZh+Q7HOn5lHdU9WXD57gzuDYa0iehzTRZj
U+AldDJrvglXauqrGLjE06v3RuLE0vjc4KvuRn4hVJ/ztWWa1ZbouyuI1TcXiV7f
1lGZ7BnCVMdbHdkVstzgnTmJGXyZqrjY2V3pljlGPLOHY4s5Pk14y9T9mgNO7unw
YoDB1EF9CxVGJ4wyvk/Aix8YVtBGh4nKIEvgohCnkAcZITaeLiBG9dFSCtRIWt5q
4zsxlAbTzw9aDPdARoE9IAPiketn0YqbsVY4U7Tl6wTUnvgZ37kKD4iku0uwcOTZ
qwsijNcIb8Bgy4tVGNvULHcbsbJ47BYsZu7RZ27i4pg/w3KSigOhfjXEsnAiHUk7
mKvQpq8GS9Vkeww/V/yPQUc9+7uhWFsUhXzXfRtdUlsoeooZWQYQn7aEJ1kqdO7Q
CV2i9LNP5h20ma3RJZvWGG0G+nRnDu2q4MJueLRVOShU4L4GnYMFiQD7L0WRlrJu
LQKccQPP3BAzOXc9Sd6LvS5Ks0VckWh0Rds8XFk46KV6TJegT/Ph0Rgf9/4uAxah
mG+8yVvbsVtu4h5qsIa8aH5TQYYorXyWnceOH6uihOLO4wDNBDOBGq0chaxbWswg
bDO3P3GjUEmbuZSYwAHiYhHZHGlI2dXyaBapmQQZT3s/P9npWKsvYhdLZtYHwD88
gqxql2ykeekXquzuOur2d2v1DZrVnP+i4dr5Ysxs/WjU93zvJeY8F1XhwRv0e2Pq
QUU1jH4zK3RJIUbdGkyVI6r8O9K9BuRoiEQH6oYZLUJBq6bM9goJ/8J6lvxANMvg
OVgMZJoUNqnCGA0qHbYdoMKGNvCYC0qInmNj9OVxLDkbS6hMTC0C35LWvdEAm85R
nxFncegl4q8ij/dP3iHxPr19fSx28tj8eZisHQymjcr8lCn7aHWt4/wCCu4bGG0I
1Xyaw+aljP8fzqEjrBbGmLTtT+83n0LMfZ4ZaLcVnpkzLY9N2LyTufDIX+vGM9PW
TURtWxbATr9/aC49WNZwD3tTthmqdMyJoNgDZfz0r96DpttaofksBR+eOF2PtoK5
Van5u9MBiGBfK2tpmAzN6e7e1bg8O1Su9lThJA/72Axfu7gkAKm/iCQvvin2zZLK
V8drQeCesiNlxUDFoN6e9z0QkXuEPqGAURzLC7dCrWApRjbODl7MEuR1qAJPEK+E
qlMGXZbmqmJCSRYiKU+rMdYyU5hiunudLgymE1QtQhsBaTyAmqOWZyWYSJzJt9mi
Q/JDkRQXHBwdW/DBZIGe21DqtV7NSTzMjFmMQz05S5HhdAkhiCxlgC6E6rOqEUpb
lfI4+b/M2aTmMXQ0DfO1ScAebG7qwOzSEoaP5itdvfjJFJ6sDxA5Ud8StlDSyPdD
eq2EbL2f93Qd9BljsB4t6YVqzFSOUTOoSbuPKo0gQbUB/DQNJ1QkffHw8ldUhAZ9
RGQ4/WFODo9qwVTxTMMgNaRt9ldTZwGW2KtP0HQusPqqWiwSqV2fCDeq2OxfhjN/
M0jsHKl62UkwmFTHeMj2ZSxlQDM3ZM4n5kfiPwNtPgiQJhzJ5RCDnK2d6aeee7/V
AEcEg/AEh2f8RLdPHtA1zgGDVr4hpydAXi6bOxd/QCgBEpATUquZisBJq+aNkl50
6ZG8lYMupHGXH1D4ZlDQZOGrgGgYRb3PM8lhRDzZgep+Qyvd43TgRKhW0AT/xv49
1NMw2Xnwh9so/vFTKAZMZqOnrAKhqMbUeMcLDsiWLRAHlf42Y/sXLNRBjXkBzZ3v
5asWMwfmwU14yBF0hceFMLGdMvkQy8nZJ9oRd4xds65jVkt6W/1M8ljV9sWGwfRM
wjHPd6bAXM9ypw+laa4+yhEUDZ/GhB6HTpTU1qnPSSoBBQ3oKBIX7ZfjQ7tMZ9MA
hXN0XQ3uW9GJLGBgHnJH0YD0uVyGRm8iHLbzJrQaCRVY/CdGtY0Yh3MyM3eCA+bz
ltN3jvz3/AEeJffDmbfrZrzrCCStXEN+kZDZfqHgEA88IYIfmOxrHMk3klrMsG1h
CGwC0D7hP3li2Q0Jc8ihDdaFMVtUMpHTsdjTellWUeFwFqWKkgXBA+VLaqtUbfry
23F28fvhe4l2E0ln04p+dCWvc9wSV5kfPJurGlM0XnC9kXuq8qGeVy4HKgOJYXe3
P9mif0jQZ2g7da9Lb/LfXFv1ASA5tOGZDwIqJMBZ3bngInYMgGwzzjgclKAjb+Qj
HCwSnJWIjtFZiHu+nlqkYHv+kP+keB0Yvra5PTd2riltIeUEMeq021t1rcw/CaIT
EAv+x5NpIvmm+8YY3MsCGn03aQT11/OB6iI9k4Hm6ny8QcUBoalZj3dkWrMGAApw
8xPkT1LhzjcnlnNEZK+4iGpktP5svNYBb5yKaaPB6P9eaY3gMFazz9KmKDgU9go6
Op2xsk6EiSYucd+ZT7cL3YLGWswS4CNg0t2WjIEVp6j7+0bIJzg9VHtb7lfeqmQU
SXQT99p2a/SqE68fv4+wwVA3BOvotNZFkpPT4garRK8JyOak7959OHnNpY73vW60
K/OkAQ/kU8vz6CkJ1+1+j08y86pWmlAEc+q2QANF3SRSZ/AT8/Z+IJpcfGBW1kp4
WX/nryzrjvS79zVVNuNcuC+X/7fO/EDvpUjaa7fE/S4tm8dHdTNx24qjkaXttVUD
c0jFHBRNICSAX3LMcbepcTJ+QPswec4L5fT7F7UJITN91KHYf13yNl+n6v1nhLLj
/xPZwA7SvX9Zry/AXkgWnkBhkyHs0KwAihQp16bTnhgy4GCAbttK8KEEsx2Jx9oV
aXoBZiYLYLqJsLbi+K6J9DdPCjXgZmPHW+8iG0+Uira7hx4CG37AXjyt7CCKeqQm
2rwgbvYEbtIbGL23X4a+35stSHqPX2U+uIIzynjcVF4NGxdErrKmrHyUysVMIpPG
dntNGs0UmvuwGXMTgJIUS18vhH2BY1/PdBeEFLivgDA8kSmQ/Oq8pI2FYsc8LmQ5
v2lrD0/9buLSBMW1cGF+qR2f74GvwunMM/zuIgvz11d2PW9azxSe1fTqbjxGLix3
UH8NEtxLoWs3LxYwmQ7Mf9tcgZDAePxoO9MmyqZT3t674NORVDydomsAwpSoe2rq
VL68PmeMY6Bk+wEgQmwwMlzJXvURJiYaCjPOxJ4CNDVI34gCVxg26nUx83cSckcR
VSb118ZCWmPL6UU4b11038Ffac/uQJj0RijZJQxa/uNhg2yN+D38ICo1rzpcgzAw
Nal3KQtt4ZSC91jY0wO0CCV9Bvog8LmjeL3RqIKbyt5EUy4Z6J5z1DI64GQ9v9ZW
5tJr9bjl93PtE/u0OIcAszqR5I5pmu/d4z0w2wwStd2DRwxLtGGlFzEBJ93jFbQa
npuvJMFUrSrFuLtN+KxuleOZhnfPG5sEepxPdVYPMTCVdnGXHF36Xd8gyRH9KL+t
QipA1aHJL9okFT/UfIpvayt/x6MbRnY74QMBe5Y55HMgFQOuAXJa85ibaRRNGenh
KDE1VZfNbZDYiksHC8rMAhD6igJbTSF6s8Fz5c0VS+SZYf4Ulbox2Jk1QofhWKFy
gTVK/De8OPAgxkyWLJIEneQWWVv4Yezwo9P3MTBHQ15JYyDLopP49J3I2JCQJy7N
uVIgc5+crT4huf54nCVAifukE74yZvqp/sljYLUZoy8exMRYpJzYDTOLVoq48O7j
Z/kjSzarUGzXhTxxL6jlS8KBWZCxjF81CBDZ90vh35MEctA3q/X5DBr1w6c03H1D
j+JO0m3ZX9q+H878HrpWpdZI1z02AcfoqVvj3dPbDXzbDuOzSZHtfmY0rWUseEzg
KI+nVVmy3JfMyQUSYSCuYJHWApDKXWbjjlG4G9RFBKUJKLLf9ig/LJaWci15UzO1
X9lffBFciquO28gWphRpoMV1kbCpmIBO1T62cL+2oipZuGWHGbM903sxMTrj2GdX
MVI+XcemyBeI5SI5p0MqfNjsIJyUmwxkG6x0XTnoFOuTkGpu6IZunpJCz+kJhcn2
9SYXuq20yvR0zc0CMD9JPjm4BH2gOUO4TfWA+pbpfeLcIwrmT41zh6hpuGL3GpL+
NKUZF9Odxk4KRWmolh0RvdshOYdKla5pKyw+rEtNR0gSdM/gfJN4um61wLoqDT8W
i0V65M1xgH26kecB06tDNo0LRnsNQ0B5jNxycY+Tfpq1AemIyHMBODxa78FA6sAP
PzkICjt0ZW7nai8TtGkxOwDge7evq0Nks7knHxMNYqlGm5MbLhHTP6SULspsbvot
btkhR70wSgxegPxKxQ8b3U1tJy6fTohQd8ZOwLwvmQiV6hWQWgFf+7LPf388lrpj
LQValQm+WzzpKcKzc3IO9XI8wtUpOGx6xLoLl63w//nFBr9TVklQCzL1DiiDvR67
0qI21t23Cb/j+dfte31xHZiOhmuZ9oBx4mFUndKh6PLrATbteojITlEkGKotAZKO
TyS1cySuaRc6B6H7F4VXu7a7uTMK0KDCFwTONctFzHAWrRJ+uPhaiJU4h1hUc/p3
ETSD4nK24wo/mXdQJC47m6tUovWIM3x5dLa9DGg4qtc2hM0w7YHD1G4YLFqF7Gll
/C+K1iDQsaDc0uxQP4FV/M+1Pf0tiJHAgeqeSHqzISd1X0i4jQ6TmWyB9Zb1K0u6
3/C0TKgZrZibTD4P+oF7et6ucEET6qgE6I/tSYuNWEOjtYfmKoMZ5hBVD/wXQMJL
uYQOk1nFWttgrhtMYDrRwxF54HhBQjwA6r9hXRfg4gR1u2e4+jIVesNgne/7g0Z9
aF0Q4l6WdppyJsuVQARGeuyON22U2xGDl+jals31+uAPLqTXXCpM4+IodfFCTvfF
sYqHkaKV9GPiT23O9IprfPhAklyNk591L4bdJY/Cp5y7ZlWfmZW2mbkfy6LnVQiE
aTb3TQqIrWtzNuzDbqzrVDA2yBXfTK9nyf8xlRQQuI+7vjVlHsgRgdT5wUUAiqCV
mOCpfWLNzeb65DPYiP/T12AzaVxTVxSL4OTwZxjiTBvXTnFFTkO15IwAPMsGF/ze
EaI3ChFAOTz4m9QFlMigY6c13tf6dJ/Ko2ceObj5jUJixBhFdIvJOWkx50YkuyNN
4S4nZCW9VUjSq1jBCKhnW2kEJYrnFfTnSxMVkIJddN0zNlgVTrd/D7J+py3vekrH
+8RZwwdipIvDEV1sMdvaMl/zY311Av1HVgLzjNCedWFOGR/LHq3GCYyXvPJKS2Cb
n0OqePjy0UaRi6PZFBvXTIcoG3SxmK70HSJrefWf3DAcG2ggwnohi7Q7vy+pNEXk
l1ZLcTWN5wH/N39m/ZRJgbvSYks8Rc1guCbGgmXltXfzFbsKad7pM0sGXdt6hH6R
X+4LVu7t0ShCuSWSgsaulMiufJlehR03VD3Df3vyDLCFbcuocZWyOhfZ25cghFVt
ik+0huXMQX+CvAzERl1LrtbJA7G63VU06vC9HhJeTRWVgm3ys8QS0fq7LectMHHr
Cgaihh4gD82DMDbqJhsk9v0Y2Z+Tu5Uo+1o8EX1VR5fsUyQDDlj6MZpAJ3apq58t
GKCNroxo6Z7J92bPTQ49KJ3lcEmgqtCwmaptKR4xXVbG/pm9lkHjpikBdlcT+v8R
F42m+l9KLhUgg71B9nfs6BdHRhvy35Eu4xuZalxFQuLncumHMxzuXmPg3FFM0VJl
LF3qxO/ZhHyajtuccHfKKQ7hzYOOOfjByg383i7FzeyaTuJAHS0AK8uINMqqJl5/
S3+hb1RK2DdWv0XzNuziLlaEZBl7e/hgGjHBt2c9/3EVfPQKfqrJeiP+Kq1m6332
gRqXNCJTpWBHZyOychPo6UOdVG1hsPvfOAryfwf/cZNm77pEMExyQlzdrrYPVSc2
vGJx3BMy3nIzZODKHSAVl6sbENlvonw1ExRPgMmrpmyRTdGYJ5KaoyMFW8LRen7G
+lRYlANMyYJGVPd0U7Y2VePDPAcfJFNP6UyOtLhpOvAlJxIMGQSQvBCJowJszc4E
KgVylEszLvHs3Gf0fZZ/ZV89lPV25I55H7MjHY5LXhDduGbh2QctiuYvAgIFiBOi
AtzRL8hz1RTAB9+AmvVcr/yQU7Q9Zd5FhHs0KrfIVeqhdCDH8fBFuxe+X5FXAiry
aQ+s8vC4OPZLElpLL957RtnFjSwNb5Jp3lD6Y/AifEExMHvRSAXkvsp5Rh38O7MB
gpSvZL78uEEOAy04yQo+ZAGfWDLxxigFLUJljkamJEhFbRAuzJN1lN/tj6vSdt8Y
+vIj6dGZiDCosePuRjAH3bLkkqRWMnXuZkJCdpjOEBtcOkiuqUCnXnEi3DRzjMDA
ji7cRts89fLD0r6pkDvzHoWOoNy/bLyQiU+51cgn8XyZ8k/jEHpUVNWVL+vDFHXp
JMlQF6k45uW0kcblY7ZUEceNdiCwC85lo9Z1LPbQjR5kvRLLokyCl84otcdge5XX
9zCv5w/IJ+0+ld5IEIn1XRaDt2achmGMxgaZ6EGHEMwCoaLdhV28GrQXU39OV0eA
52tno9HFb5hxjmd+gPR/WBlAjtTC7Dan+GTio2Z1FPfbPc+29yPZcmDwGWTz7GXD
1mc5ZfiuDIakorLmvHIldRvTEQVDJfDaE/x7XOEZNt9H4SpYIClfwM9o3NKwNnXZ
Ryoul3ncE4kHlxjsEhzKcoqAJqXyKqV9cm+ivt065r9U9pqHF2Y3cE0rLYlAUevq
oY7JSsRqZ2uLiSjeb8dolvPH5SYdwFkuvpuE+GenovHaYopZOwUtDQbecinLpa2w
4YCsl/wllm1XrznNKnLvXyUulGWoxqDUDSaQWLIp5dZ0kEKDevlGdCn8iasZFqhd
BNbNr6oqrs19bxo9ijE53K81xGNqKSwzWz8y70+UXGafCZFWe0DT5QCaXBva5Md9
Vcl6OFyufEhqTauFDtBKeGy1apHe2unMtzRIdH0W6x3JMuoWOXkWVZ6CeTAcPuSh
E2AhOpkRF+2cVA4tNsA87IoBn1EUMvwinLwYnXtkkVp8TGO8S0T5N8F5ks/nwyoZ
NCZF52ygCSVVQWjJKs3C89ar4Kybj7DM/toT/OEwKUfpm/S5FIwUcm7ObkNVvjjW
c2kaHGWoHfe61kpNIWj0Jh1usL1yqCVLdx0q/AM8mFOrraPEeMYUBt55jUYs4bEL
BNjRDj4BZVc25Vnszo5ow3gpfN8jeeMCovdapq5RgO1goD2oW+e4r3iwb2wVC99y
ILocIv1psYWd5AwVt1wqs4PkcMpMSCBL4KZ7SpEwOXdtqyKebJkBaUhQ55+wAFK5
z7V8EO13kn0UOgAWOpvJUGY1aL1xdB+/iAbo4+3gFZVy6wPA5J19n7PNq8raK46y
0VX8lvxBjknLsgm2ecDES1+Zo5SJm5WyxNgN9ibZ9cjrtYZQRgq9yrSgpCNB12On
+KXeOng0xtFV7YwI21nRKXBvdjaFrxI2xGqyli4n6hkPPSKhjPelcc21S5vJ4piH
KWLllQQJBVWEexPZGHIhu38l0vVS06KsZnMghqgWMY8Qc81V3C9kVyNwqwMYBwuU
ZAYcfa1oKg01DZaed81Kftj67nntVcXuIoEaO0OqAa//paxPp4tYOro/qGg/I5RM
itQ/do2SOUiYwlgkU3s4c10xP2bG+nAS5RIMRCSvSB2GFgazLmWX4qOmTB4bJx7z
KdVsmEls/ZOjZ0GTiaA3ZIGfKVbs/O4XcuNS43vsdoi6v/6oWPlEhu1yrGybmiFh
EzjiN6W8FkHt27HAju/w1RaHgG4aNVQarW4yITbFwq18tv58xp4eH3u7B+1cBJxE
6tsknEWeMGmNZthkVuFftTLODQEGvyraYEahGUlA+9HECeh0aDUKaKhPkFxBzZG1
wPLVcHfMRGv/yKHI70ryf6q3Wg1WDLooN8BUrm3bRtD+TRxTbG/jQKOGf8yj3Eco
V2RX943PnzkuoS0IDUCIZPwMRh2xfG4JWK0AtE86etoplsQnqlWSgvN93xQkRKdP
FYNpFjomtQ7G9XBNT3e8odVOatXt5+oxTta35tVM+oBj/GDq1LDqAOfQF9GmMG2u
MqF/nai4wpiTxb7ycpSTcyC/1ntG2nv4bYcq8QyfYIajhhfizQCJiJGZfUMN4uTi
mnoi9NrkzRIKKexUowZ0lOwkrJSn8S8UrSXRtsJ9/8l3F9aTM2SaoMvfie0CpRZw
f9/blq2ZNfZRQ4NhTSLkblUuUd+71N+AGMDpXj7cMXaPr1BQev/M3tk31M5BWi+q
yMZpruaFc2cu78N5XfYk29SGjHUMoWy11IrwpA9/aEvxLtrKYwZDf1eXMhh7SF/C
G6bbJmFluUZ2ZjdphL4GjAwqQuMg1kfyghlvxvx4sd6PK/kKDAuAjA6Dfi5RZ3s+
FJqrAv6ZKTESB/LUS+pEiVfJOidJ6cq1NTfowDw44f2uFn0kEZEI9lDKS0aGD2rK
LaX9+nmcqBMlbIQxfVw3P4TRBjHFv/hf+EosJzG64MpB5EDkMhDDWM3ocyqPKUxq
HZU21ZWh9jvJtVNxJ22gjbjuTGVI9uSS3Li/q2LEFf7BdbXhoqo6TJuV+XcdKguv
vL80ShayFLybAe5dlj8SoAtzs0apokj9DmjT+nWlz/pWvhVCxEFoMsCV+iBAbOdx
0BjMrIERFkZtTGTPyT22H3F+cJ1Qh38zUXeftkLV0d4TS8mlQBTy5QS+jf5vThLI
2fm7kM6UgbMXGsywdGs+fdAPFATskenVXRSNTXDOyv9Q2gALK4gUNWgepIkwZEMU
RZ6EVLgR19O3r22490IPEeYAOi1Wt4N2LbTjMY0aXd/l4/EM9Y7vKc3Ln92jWV/Y
IewafgA8zWV30rNBgD/Qmb5qXzoEfQOoNJD8RJ9vny16QdEEX4+QdT2qdUEd4p4b
Mg0gefBw0C+Astpo5lS9U8UnkmuCsgJovvV13NO/chOk+Z36fVSeMecDmqyEpBov
yfNVLJyH5Rt9VSXBxTmpGomzetaoB3jVzT9TRwBgfkXD0E5a8/d1ZbybLtS7C//6
GIbi2sMGSNtdvbivQEAYBtd4z5PX3ePqa/wE4zouTvZcNVMjZ7ZJqCN2FGfXN3xO
t6aMRhuUnjHNo1I0XEvrbgWj7Bla05pwIyv+bYjES4ZWFgFz5ZGrtpCNxInKG83C
FOU9bWL4yIY64HB4fdQ/bPRT0U5w10+MluC1isoTMTZtMDmeSuX7HECxJrBkhOjd
zwZgGcMAhjLc90qxUGL9K0Qa8TyeqdVsf+t1XGVHJjDBgbZzHM9ck0X4J23Nw8oq
FuFevH35uJXYkxQ+hikGU3mduLY/Zo35gYZXdt3fPxTsroNmU2Uu6x9ddjGYrhrV
eK6SfL4CS5N9eabtDmEXdnIFv9yXxPCn+WtIs1dRvp0/2v87xbNvrkWTqgdQVlKp
UHlz0KhhooLBpOV5VlMM1lifiiYPCs2ghWQ3A2Rnsr8RACdyxBplEdMsOGMKSkP/
4WTEyI/urgIRKD4LnafvqsjasWb9+BVAa1zRzScBCEMHLmlZTN8ngGGLFwyd6KCB
SgNLp4wTd/Pgk9NKLl9RJ7yyGWaos+CJ5dGdXum/G/ssgFfssA5DPzJ3GvGYiRPt
KXAR86jNtj4qjUiiPKVv988nGv0Wz2WHpkJqIQvSmPNE2SpAK03XTGzpEervSKWz
PCnNxsy7SvT0gSYUH4B1SqLk3d3hURkSp+C/vXpH0xj1uXFtMRmPD6RVV1YWvG0f
S11rCXkg0Diqa+K/qR9TFdrTFG6dJn+qwVAtr2D7LJNd2c1nHbwjR1YCc+ijWPZT
cIfcpFV8ACwQRTEaWtHRb5j2bznWSB8bJwhVxt1+2rJAaiWIW1valojC966rhMtq
xWRZtazLrVsyQd5qXdO+7hpZ96RQd90Xuxx4lkbdsaJqjWEb9K2f1LesdpHgRYsw
j8eXGBSYXRUUyKa7y4yKh/B80+fpSyBOqrqmW2v8F/+wT0aSfPziWQA8TCXcOhXY
KE42HOd3cf3DjqViwejgJRXMo22GBmCREszCCUWNYv7zobAbxFSx6CWoP64x5NE3
+k1lVbGgsDadmhSmK9eZ0Yck7mUOFlWeX9yTknksv9By7YU2S+EJqBHYZLdVQI1Y
NeDAaAZ4HRL3sJOl59q3y2GL5dbUo+FfRREyc8UsWwDx8I7IuTnlwr/yzx31CPz6
wzqGkZsOzgTUHfhcf+UOAyPfCPMjLdpQqWLkmcicpPiYPOI9p1GvdajQGUmS7bLn
cfbVZDaSgXsyDj2UTV3UgFanYPE1D52OEzMbzJNE7dy0dhAxnHBfjmQA+NkBlu/u
qajvkXA93uVZjPK3fDL+pjBtbaaK4Jwsp4h2FPN3UrASjMHE8jNIqHHL+M6ZbKGW
6KIY/MzRPkFAnXfzGb8a8Vkb310JNJ8fLutKdVQmHxH8tnGMrJyLHrTZTMKsZvNp
tno5XagUJ7tLIDrvnjbypXwA9smKOBGCwdc/a4iLGfbsFbAmZvKJmNhrKc+HtJ3r
qZcXEvtfxVNBODnc1OPIrmMgSq2XUnesmjTG20o6u9Jqi6whd5CeMFwOlOe/mGFf
30xLTWwHXVs9f1nf6C7/KjpH2mNrATUMAq9e1K2UlDDLyDQpOpd3raK0xRxTSrhf
ogoUGOmLb3DrJyPk1y2QiOyR45RlbA3HnwTwOBZFrcaG9ISiqwtzjYDZYY1KUi3B
1NyJxRTbB5yacYNlO7OA6rkB3h/hFjTndgoyhySxYzI//fy+uV8Xbbo6x6GrJBI5
cHv2wEM6n8uf9dMrJshxkuhfJ8IyBOO//esSBiLcPdRUsWYdk6QJjNErCRiTbb/V
xn0hFwJRrV0wyEW4PM0WFv89YGVWnPJeJ/QLx9AUVxPW0SZVkEf1oEQVwX5IcAww
y7EHOlqY02NG0M6EEYK5waeScRuPw2P2pRYxlaXOqelpKRwBq65qFa4/TThSOr1H
3cy+NP6oK/eAyNn7uOIkarsNqyYic1/jCd9Ga1pnH218sfmDpa89TvMJ0QASf3Gk
0rO5I/qhjtAR1KbyAI6QKdLrNEgYvd6vuJ7wXtoL8cI3OQYO+R7+VfLJamm7/lh9
tAlfHN7BTUoPFz6FYDFaYU85qJc69uBt7VXaM6qx5nzvpK2LRIpcY3E0m4bZ2UHg
7B4ypnX2h9TZx4/XbtWWTqIuTjBhAW8kjY0HZ3Wcq5l8IieE9GxCq8QZhV2ddRaX
JY0/VjkY9LjFvBC3s5yoVM8rl6/yEGgpBRcI+qpdT0kSpJIj0/V/d5hfbbhr5/wX
dTKw+teWSc7G2nt+pmkeHRRDFdtJjyMEwlMlGXa6r+usncKhJpGa2XkzjJdG8roF
DxS2cMX0lJiVVl/UOINWwhgq2xtxa+BPYllE21/VAX7MYzh60Hkqc0n5fybMbimi
KOgdK6+jtXcDYLeIcIR8c045dmxZDHtgPfw9P4EWxnV8FhgqfOkMmUAV/Q8Bc+rV
nttL75GK3FtVuezo2VceAWrtlNAc5ihstP1p/K1Az08TdCeL7TUl6Ny4BzE0uq1c
5XxyPvREgWJJFkiQNVvUQRkM2noG+Uw95UfR4VJNC+4AMzIZO4pIm0JcSKvGu4sE
hQ7ONbmEWmq872IkbSlaBzk1Rqu7JJ1RtQ/bmcInqgi4vZeJAduaWOxIxJdRFzYN
X2GLIK9opu9iLQ0fg09Nmt6oOy8jmKL2Iwv9P1gTr5axKs3xH/2/g/NcS7lh2GY9
x5NYCcQMWJpX+qVYNWfguZjUSwLYleJjuOshBgyq1rciF1Kg68BnDm/C8+45hMoM
x0uwuelUs1TWqYe6jqMrs7h+v/u58HILxILiDvvBgSIP3wH44zpGnZqkRf7Aeo9k
xVT82D5QWc8esbmLSZ3oBLgLGyBInw2c0QolnOha0fi0NSFXJ3riuQ3CdiBTxkOV
sLI2f3rHhgr6yE/ec54GkBLlwDc8rpnRsF/rXOg1XbhM6MG8RMlmwquEdQKdSCK3
btIUbe8iJA8elpkMXEHWtZ8TWVDkVzspcGNnIQm50DEyc3JKDDT8LH/uJNjowdIy
cM7iUa/JBfsiYWAhS0oYqWcZROOKiCeOdtS8Dn7Vc31Avm32u6BSZJnSEIXHZeu5
mXlUHeNLjffJaq3DcL9IhQ486NV83ksd01/Dx3X2lDvDyEMRgkTu2Iy+4hqkH3HI
PC8FjBaoz8L/h6iynez7M/9XV+bFayfK05x0Zi7+lxZMt/nW9P3MzBXJ8sc1TbdG
u10olRXc+XxfR/EUx3XeS2pBGgoDqUmO87mYMTCGlIf94ipdXSoRTUO6lx7A2V3v
WJTa7QxlA0yPhzMeqJMrF9f564tCCKG5AahE+mcP7UFfOi/iJebEe+ps7xhu/oWw
2K+m2O6GL4EVdzhAVgtGMrupjfE6Uiiqq0vOPO72S9G6m8X0sU4Kyci+l/krtc4Y
+bzE+KrdLfRqHcklQt7GArZevMfXRfkzJbR2+AgTG3ohcOt3SmFoLUSRR0vNe+iP
FDcfPZrou/D09vDw+PqZ2e5UJsjqsBW1Z/W3m/mjNJSI5SR8ibnb4tOx4bfqM5JS
ZYopGrnus8L7nhSJ16SLmYE3R8ftGdR6r0V+fQ4yhKhOMdNybPsew6VUqpz1Y1J7
YabRGX6PyHMY1oQsLZ26ASvKmjFWnjmcmIbG8jYx8/mSoJb5Kb5OJHnbRXIf2klx
NZ+sv8Kboj19tQ2bf/7jKlWeKk0RggMSodDEZ2jWAocWVPtl0lqc65TW6MPToAms
Ev6/Ic4kFvaZgZmTRo9iDcuv/XreZT5Yaappf8gx8mVpfmQ1jU8XcfjoKj43UMJA
GsH9p6ZRUTs1/KYS/RFlaQ2TYOimxMe68u11lTK9LypI1kd1zHixqcXU5Bm8avFe
wT6hH0qCA+NpG42r5QTPDb+WEjj2MQL5B+SqGfhCL+BGy9aY+hqpmDMiBZdt2yDd
6GXWLFkwM374qOfxnvyRz4WKMDi4W+1B8hl/fy98XVkLh/QyLi22CC8sOqvi/aCQ
7qZyFlvnucJx+WnFB7zivp8mUyFp/n+AamvIV4Pfr1KljsdVkp6oNjek1aW6PznE
3/+1gadLZlMDeR46CjoIrzP44vekdKyELtq75Ktp7GEptD6N5s9Bu6I2Rok8n3sH
H4fCJ2XO4owJg9J+j18eyDdWAa+ySkSIYnBcODkAYDxiZMvXmEMFqDsHANrpeZOl
2nCzfoWZYdJsO7lFfoe4dcZmq7kHMqDkdh/87tvOGSoE2ea5drTwywJG9nDYf/Sd
1ufw5ZoJSxrVTV10pwqATNQRda5h4Rkgnd9mWlOjOlovmvKzuz8qCJIwLpkT0pKb
bIS/+BH30C/h6exmyFeLQKKIqUWLH1edj3wtLM2syfltl9gdPCon5LitvBAs9o4q
ZrTVqmdgLhCN3FZmJmYUGetF1OG/3T+ue80ONd5YYWYvw8g+bLr8nWEfnbMMb3Sk
vS9qfxncXD70zjixRlt0+YKV/VAOMGT0vwAmJQpfPfsYaGYgD/f0FVb0EG2K86a7
79ndQ+cyrsYCUjci8p6yAl/oe6Sl7W7kqjGIZ3Vnh8QgnuEZKHbRajKrqVt+tEIr
68MwcXbD1eBJ8OFqAiRE+egxPZULDXSjW9a/O47KXElOZ5QFDLzOgEXed4rLe/Vi
gEmerGm/HTmajtRz00EAzvSYFgzipgJUitRcxZxsVzoARNQqv6Ivzmu0DzjlsdNL
c5I0gJHOIpcl4ksxFZmq1Cf+fP+84HebjX2qzKllNyf+R3EDHfO/EgkRp1ije+lN
otwtOMP3ereDigoftMKy+oSyxA3Ah5dHmHcQ8T6HCsdn8PrzcDaV/UZ0Y6LhR5zA
pl3BQLXbbFrK0U3CysZPenqJfjz/DMmafjbrjiXvr18Fr0nolrsFYaZ+HfTNqKsb
8+uuolrnmaA3g8KUtdmYBWh52QcLiT9v3WrTbAHFNvYdd44u4lFeLdetf9LRr45D
a5YVvtYBoIEwL7XcD1bwqpxG5LxAoyJq9tgY/UYSYLiyKd2a0PYQSkRKhF+EUZBR
+zYFW7ag36m/KjGkAPXMj+r/oVM5EhrLkpiewXuuQKLH1/FATznq7qQ1/rjofR76
vterGbqIvA76LA2eDtS4dFVRas2xrYilqoZCfR7oat15yWAKDxZMNL3gEdEBy351
+k3jXHn7Yw08eF6ARYAkm8xUnF3Nv+/zkjw/uF49uw1/70eEeTMxtj/ufkrp3DG2
4bhvup2AJMKh4Op18GOttA4cYXT2VlsiTcQIkCLEOtnP0yZciDL1FHyiiX86IEmp
LqDQxHW/qV+ISaezQIhrij+rcxJQlgM4UkYIG4a5K8jSnkX5qt0wSkyau57s0xe3
93+tJyaKJjWtDhHjCbWhiZEJAzNhchs3oE+DkuTsPNSW9cMtCxwbQ+0PJKD8JBrv
UGMcwtUX7YLW9X/D42RkiuNpUWUjJnkeKtFIMiZhK+vsDQ5CC9nqtz5z0MW9dgEx
9s+H0Bsqm5VULYGHQ8lxQirGeGZwf0YNEscyxYQzG1SR32wmZCSyKKJLtmhzsYlJ
bfnfjkpgbot4hsCsvM3i83NQho7+66gPnIPqQxIeVRdU9QwgCHKv6GbD3b528l+k
e9rntXog58Odh5X1yEvhf25qZ/S9B+4S4bEuhjFLuaOI2QqnIUtFlznZhsrDSAfU
cX4opLDt5DMadEaSrf4Ztm0t8O0Oy5ZVLy/rkS3vV3uEsEfVeBTnydOdEqeeVZ2G
ihkWx8GSflZ8hTbcDeuujaGjZi2CAR8aeFuRHzmcrt/PQ7MV16pcydRyEvVKiHV/
DrBSxNz+k9CAJA95tpeb9pXEsiKDvtiWOaiz9n5Lm6/RSCg99g1g+MIS2nf1mBdZ
nolmw/GwnFiLbax3UusUJIfO1p/mlIN7389//PXBF5OGYI4KWoIuKm75z4LH84eL
PawJM87Idc8bunyYLWKbRFtpNL/9hO5fv5rSTM3qfFXi7ddIVZUfkGBaJO4vgLYF
sOmiixUVn0/cdTFMzNOKTNFaRJf/+0b65ZiQ2cLU7Y+0vh3nG/PQ02lobrw9agin
vHOPIeh0ojfhVsFFnxRZ2Dlw/2Xqgdy6dT/HxqZrhcBL5pgvu4zzRnnSjDpJBdES
HE3GGoKY1GekUyfjn1HnMaspiQnWo1H6djACGfnIGLo8t5IsbfmyhTvbbSgnB+Dl
mJeJrQUIhOu8u76kv4S/OJFkl1LE8zcPreGslcFcH5bkDpdG6dEAOu/zNmwrwptb
1OhAVKYwum5iqbAQwqMicEr74/8GH9MdmLnQwizdXOiBK9FCVroN8SilbjxeL47w
nhFHLdHlf030tFdosnTvnlPFG3nFab0z3+mth7/Z1DN3g9vx8vsrp5sXtvSMA163
Fn01j9nmDv3r8AT9zHZ2J+ABBDoFsjA3uU+5eXRuXyaSbG+fobtBP/cFy6fOHb9/
S4js0k3N7QiP+8iPX4iDDh94XB6tk7R/l2jSl7Ezn3xmznCvyvIOsR80y1sTXFgi
QbLBsT74phi9HrU+G31AvjFWL906NwM/byyWGIdEk5NvY5gHxHZ3Iu5uSd1YFAvQ
RBO6WFOiWaEwNe5hkXasfRErlt7d+RwqVhV/8uAPl9xP0K6e2nqlQJfE2FWGSKup
gzENed4+kJ5ukURZmGQXLlRvW9yZmv7yLjdd6N5I6SBeZK34wGL957nvtwBwwUwN
aag8n0vGYljUe5GqmCB10zi7vi7t/PPoF2C0nwRXdbGAp8i1nPUKK8yRbKv9Tvkv
HR784a+UOh5QV6qLgvVhauB4r74pbBILEesupfagjJDIjVh8KFuqeiqGQsY337tL
UWzJV//rIOCyFxEkkRxkHjjuZzfpbqYrqzXRqFuuOwn2MGOYkDITIcgN1MFdRzy9
BpHxGGprqQyTkYG9OyOuTO92X0puXHn0gZlwb+P663AmOT1C+8fqNXgyIgushryN
rvdXk5eQvyIcL7kuZQw3wAIyXeaOmT08OxIwgA69oLMB80AavJ2Is2Hq0r+mVgfP
/boxleNufJo61AsHJ62AzMfdgrCQuYA10YgBzAEmj+l+yPDjJa/c90eOM0KY/w+a
9rVcrQ6HuuwFKBb3aFplWFLZ55zxhghtGQR9jAzEgO0oopeYp3srtgQlFzjkXmjH
rh+v16xAS2klyH5ZH+ImZ9m3aTWn/CsnETtBg0CPCzV+yqX9lOWC7yzrrmwV71Ry
YHMOBrRtiWqZqnapWTYSoGhEvvrFNNRZmnLLUtp9Ai+6A2JSJH+MY3NLsESrqTQC
Lf9e72HrlEJL25v+rvUCMZHtcacMgbYBIToxjCJJEo5aurVY2QRcVS19STpsol+K
gokoS5p89L8EDtkHUcL1KKpABMznIVDfNup3aUCS0Axxk7qO4PTIyBqVbuobBn/O
Kz38OdxaSK7DCrwPy1Ffr9A7wAVdWdMOTrrYULa9x5oGxWCoW9x9sUM3wXPSOxzU
QEy9OZsH6gI3b0NVNUd+Mb4EpH8sqN+3NlbFMEWzto9EUJb2MXkPfi1Rsfqqs7QM
IUcTUbE/RtLnRMacLQhfY0cUXtAxJbaqeC4SevoXqSKd1nQqt+MpiRfmP541a0wY
mgQ0WoLsN7F7FCQ5b14e0yfm3B9nOzPshrRTOqkvtI+xNIrRwPOuLYTGEpGbR00j
OCwK1w91quzbHuLPkNeM5zLPKy2AvubzCYuTjSeq+D+9LWag8q7wFHkt3UNFUUNo
kdOgpjOIvMnoe8cmEAzl3QMwzHDscZfrzUDoLT34ou142CJJDk/vsTez5jgHq/PX
4oOy7tAQGp7jSqswCUyOUjgkBaQ3Jc/mptcqQA217mtopP9AnlRRtfYzvymAyN2t
PPtlkMBWaQp38OHKLnBwJefDF0CRqeezbvazKKCGbDugqu4J4gaKSgDfPHLkIHst
5SQmNM2L2y6CHnbkO0NNi7cJacAA9WoxOEJsduBZxNztFoy8c/FYS+//7hNg3Ry3
uSWJ8MK0QAFsoEHy1rHek9EiER4on7HVb6iX8yOwbgcW1tga/LZkcDm1Uiq2Qf07
6Gx6R4x+rrpzjWoCmvPEKG00p9V5cCIn+/Xf5K7thk4LjnJZPMML0B+9LHrDFLQK
47lPeMTJmYjeCpwY6igcKE8kj3WWcQ9E7ptx82YJ4563fCrz0by7tq6AkNmAo0CD
dVy+mmyZPtkFPFcL+lZ3SpkQFJVX0+dNm7mGwqZrhnWiRIVccu184kSA9F0afCeY
q56Om/2VQ9Tp5GVupgDJ42dWA9aZRt6/qLlJx8RGmDYEQmHuw053tnR1wn3qZ2Wv
Su7aLttdaM7W6e5VTULq/bHQ3KwC2UHFiEGhYhTQ2QiQAv/fFCHxKC0Ijxlz3KsJ
J52EYZsGWfta4Qt4PkzEMjeY8klA7W5kGEI29Rj7ctc9Fzzhf6s5tUK+A/UfRo9C
uLevFWysRM7hwkoq/UiL8P08x2N2zJ4RcncuSBZNq5C+NCAuS9n3WhzQmnPP3WUF
somrXKmLtfBIVKxRLzAvaUkvFJ/jFv1M7l1LR9JqDA/2EGRTjbrx6pruHX80VFbB
Iw1ED8wdhrs5D5bX94Cr81lWfogHupT1kN7v4tV5OmxaS0Rb23H1FJL4kRgCXWv8
VJFsCMSfmCycm3KVvTO3UEJmH7n0oBEmOrfpHwS/GAxVnMzNuuQb9kImK9DXWl3M
rfAwjx1hz04imb2Z191l4eWv2kHHCJFvY8plesO0xP92OL2pAwf24s3CFS+ZHr08
nP5z4MkSAB583PrG9PO24YQ15opfv/yb2WJClTIC4+gx3wC5fHQcXtFs4fivpH0K
IAs2LfBkvNOqeQ4sNTKRrdrDn3rn+FOxg/OdscXjOHUQwnqD9homdDeAoH2hqKsW
h/knMs4yzaHpivCbHFv7LQPHD03agQosVfTcpJadgbC8uH8f78vsrPk2Jj1pccPM
g7DXbTj0pZh/kHI7SopKnmtFAY4KyJnuGDgnojotY24gQ6jqqGoDldo/JmQ7idmC
8zBWWnIGeUmR5RP80e97LvPCbPZxg8k7sSerHsZbENhXFNjYG2z3WZ5OQ2JF/RUf
WvJS05b6wNdFcDgtklmDe3bhWraF54uPYKAsXjvVyMoYrqSdyCiOgQF8OxhvQBQh
pAkw3YoVCU0olAWJIGpq7ur/0humdNvuoNlbOWblc7vKWvc50/5C0ZV66Wk01ZC3
ZqAQxBtQhbUoBUMigIQgiB8MNg8D3l5jEK3trRbiWoxBqTPoFr8OWBbcU01nZR2H
/Uk+2FFKMudZsppOUWyKhw2E3ew1hMhsMfUWCg2KSffhNNI/2KU+Igf686xjfAxL
8+XoPLqBp6ztnPeOmBn7RAAI6IRRmmnT7634clTTkzLkZao6GKOkCM7M5/zo4nui
hUzKlJ2kEGua+44n7sA6BPAfrpADynh6kbADl9GJMwBioNbQXIIi4vdRXMGTUPoq
TcHemkPhULoZMLGK+sUUQdMIzSeTs5O8pcSntR9lwx5hJa0kBo9JN7LSEIPTEeB+
EOO6zEtYAwcYkq0LY8z+HTaQ09lnaqSzy0tQYODL5OrwxJfG/glBgIG4Om/ZvR1o
sYy2t1V/UrY/xt/tDPWvn2vToka+9KYvT8jaNDdZggqMvRtijoTJHIucs64cV1Ci
HzrmuVjhJs0QkCiEZkKSH/5oQJRLuESOMSQygFijLdn1K6z+eb7Oa6d4hzhA3/9/
GGixXMVXkSPjY/nDxubE+byL+aBmEE4QQfIrb8oGPxtbbC/QYiWsEYfsw/x9PT4w
XGLIvFuDrHQH0jt3xOTchZw2DJuF/N0Smo2iLJUxSwpkFO77LNRLrSzvPF3aJlrR
9izL9i8iQikR17f7L7DomP0XpkQF9Y5wRn1G9djQjX/gd1hIExLXzINIjypPdEjT
GqZNUw3vh6pNyxrpDKaqpERIEw1f8jBfhKBabuBAgXdd0ymGTOjCDNOCIEPpgb4A
565t6/cs4pSakYKCTJZ7e/he+U3lcgZxBcMwrLapNdquahKgKxZKPv0KeII4VL6e
sQ712lLoFYOknElMXs2W21yqS7/bCHRQ05FqQ3P0zNIQoCa+VbWAudzR3hGUfikr
uHd6GpDDSLOo+JBVXbVvaTJ/bOjk0Ailp67kZswnKI4ja4EwTFaOyKqBivH/1QBn
tlgPxY5xHmEoUNowQ9ed2zrhadTuWpVs09D5yP1+mfbG5zVjo7D20oXk4zm/vcg+
t/32pC2A38sN1FNGbweYaXI7opofZaTDP04oymvj60N69H89a99Q/enehQtzx1yN
OWiKaPAEEC3gSFNFRF3zCprxEU/l1Y7o29dn/6t7wm6Rv1Za3p6r00wieoSjd3Xp
7qMnDSsw8fbr6fO8RMY35s7jkAjXw4bcb387TWaBRd2LCMGRkA18YT7a03OXSHmN
jy8sJ5UL9mYK9BY0d5syAqglBDy7F9ItWSV1c5Xubjm5MBLvk2LPu1P9EETOEaBD
y7JpkG0FOxbdsSQDWkGuY785yAV8bo3/0sRfwO7gSTQ2MAoWcrnNVtqGVmbdqkgK
ovfryfA7J3RNiBbUTsNm3bkHD/OL5NP+tUWgzQyGPSM4TPimeLrT7YIwB+m5trDY
otsPM1TaKttwGpJ9SdWxICcmvpAB29C0rJjAofhzh36R2a3NPnxihcTy6uSA5VzZ
gnkG8dciu2Nt8VYn0UyS/poPFVPdE+NHfSCgFDCCr1nsUYpETUKg60n9faIbZcbE
BxRqFmdxQEeko0lAaCZDo4+NgikmgViUa0P5UBlpEfsub/nr4pcx7s1Bb+55nY6x
ClqXV+xr9+InIoUPTca3pJLK2wlwFdczk/SEBKJsqPaIfxvDDdJzIhEfxT5NWEob
qB7ZXAsCfYGBGS7z1iJsCZTg9K6IRuR0idazhjLXB1DtrWAqp9TTE4CeIKxR8fIa
a38Og23PPS0x9qr/PUJ0bqwc2evELJiEls5AsJSlKRtJ6LH23tkJilqYBtiTVVIq
z67bOaCDWn6Asc91WcgtQrZXvN0pJUXfHK/xd6+cZLh50zJeq3VIZKac+pY6Xc9/
L9QSdFblUAu1YRN7Xz9jrPZdPFUH6nIzgzESb5JQk/jKelntqjDs6XHQrlFYj0ki
Yc3i/V4vriwRbMgLASgUolwPa4mYCmw5yHIdMiQq4O1bYLjIzEzI2fv1Oh/Oi/HM
2TwtUKrve2A0sZ/3AaYbQLMRU1vDaEsgaD3OnG8nWNbk0w1rcg0mbooJ2B9hDFwt
/6kNJW+3OrOQRAPxKqvih0aPO1W0TgxbKndkY4Le14x+RANDuOrAZ766Fk3VAofh
x+s6csgEz9KQ2Z4yUW5hbqvTnrkrlLQtBG+s5miwzkbWbcH3O5FuR+opc0ISTe9u
ZP43DbhcjHV86FTLA1rhX8p0pXE9uAs5s6NKOGKMPEolSFPmvQujbKI6F7m3A//y
Qoyud4bAAKyAA+asFdyKuUcAllCxpinmmSSsWmMhfEu3elB2cELo1taHch7Cu1d4
vrM7vVLAeTdC1V/lAFWFPV1mUkc9axfx+GG7HWRvxpEaKOlAnkjDZLa9JAJXN2wG
+EwX/m+qazwOWx/2ERDnF32vOPjvRUIcnGksiWA7NUKeCwG/DzkwXNyatgQB/VCY
Rc1troZloiFweOicvv1FIwIcdb0zWxQmT6CLvwKPYTC1L8eCBJaTWTXIHRCuNkJr
XHzQzGtT/9d/Gxpp5ElRmrNvheAnBI9XR/DTztcIahJ8C4JV/rhV88uhoTXDkRGA
maaVrL5hEgo0WIA5PbmIWUSSIN8d3YngxSNmXaAgR3MikqpoY+xGJG0/eZP7CWWw
4W28qLis4PbE/qmxkdilB80shtqwBfuTFEekpErKyVDEiW9viED86hPTl9sGO3oY
v9FOd6+GHDw1pjpPmoG4jGS1PLBPFPmNPkgQUoNCk7lx2LBIG4X9it28g8QDoxEn
4QW0ciGJJS1R6yZT3OY3EvBsjQCpjDbb28Hyuh/ezVwuhGEN7odxtI/bxoPmrLtN
5l7irhTHB0iAUGFHWL6hOvWdmDlgVfj/XmskuYmYV+88EGgtjb/l1+K8X5BnB9lw
knClCO1Fm8NtCNIcy8xy/LvMafg2xpc9vqu6lNaUGCqZP4wzvJbtxFJGwis50ulu
KxYM93w0JMbyY9x62EST3w/HRotTRqlyuSZhZpMzXqt5wWSsRx77rdafhcmKiW/5
2e+tJ6apJHK3WJYddP135dbNJSDRB/int83DDqxLL4haEtxNdoEjjCKeLHNhbzz6
m4bY4hd9ep6GypDDNlIdHZlKiM6pVD3dC5/mqIo34P9VwOEbxtUe2fg01Qk11/sc
qaaw4P8MQiguQfdjGdoArK4HMi7k9YFg8itPWtrjCgMzOvpPOzgDXkqKdJ6461ZE
bwF1CfEcYksUzLzi7Kw628qktnWVbZ/Ci39Va4mzGXwr+P2ud+cagehrbfLKb6W6
BbElPkE58D2D0UFzqs4x3ddxBegwdv/pKQk+n8/83uxBd2WfBwZzNxXpfXy2kTQa
s02BKSPvl/R9IwSF62FHgkbILUz08JstViuqQ2N1hkp8IjnSRwTnVzlKw9yv7/+N
tIJ6UCfoq0PwixcfEcFvSUpdgJRyVXyNKdlaEBz93D2i/c6J3gxRE3v/Rrozg+KB
7oIVElw9ogZD7UR/HYPKnk1LMO/mC1MZUpCtopaU1VWsZhNf1S9GyPENLGnqq6jQ
1r7KJRT4THRsDCnb0GpqsZUr7YxDwndq20OlUEzu8aLIqOYVdhKvsmBouaVvVx5v
GT75OdYtQkv+C2u2SSYPHoUhzqrYl9bvaExBMGjQJymLF9l3QMQZdXm+iFjlLINe
30eJs/HmQhLZa9QEED8l7R/Sc5oZwwRJnQLFe+pGzTFWvB6s8igobj67bfYOL9he
M8w56h8qDqMdXLLjAiiB37nGwRMIoSjYl/QFn5bUQasQ1vDS0uMRx3vN6fTxmZIw
oX8A61NiEFGsbX6W0PDMVWE5gXsR2A9AN0pet0JIJx3jvfzO9SYBMdP1UgnMelh9
d9ux5hW7qJ1cykf+a0uPAgIWkvhLvNl+igNQUTvtn9hjBi1Wnp9elllJ89k2fxsF
ZdNhHRkT3HnSHNwLoWTkgiFy1QzPWOiMlByIA7I0lxqPb3T1leHzDZk0wGUB6gml
O4L55I6j9+3xo+WshhxSxxQ67LdAlms9q4II34JK2lH1qLD6be1xMFRaUaRP+9LG
E3xNAUxGPc911dYRxl8cKmFAQm2hUevZ/17xi7WYhlbK62nnriWV8Y8pD9DYY81G
LHEqD0STovSGDGwxSwt74So4iQP4dHmWXEy3Yn2vUOTymWRBBt04IqkNFxf+jpIX
eKXwjq8Z/lp2jpSozwM9dG6eG1sxRGtR6s78fYE2cI8NIrSzgLFarc+E09pJpkx7
Am9aW3xXOw6GHXsLvfYVFXq8PKUFnWxqyHwF+n0hJvPKmtDexEmzWHIYnrDQ/B1n
sPcUpAlAR7zIjvO8MZcKaTVlkwKuG4aHODuwZWe3Iv9doOTLcIMvsPeZ7aVdQLY8
NFrE6XmfSeUS8bXRX3OOHkD+x4pns4Z5XQDoY14VpF13R7sToxdoVGvQhYw/+fYe
L0JFy1RE9+lBwmFME/y1sBDvWy9WBc1mNYyiT+vVzcxB4lPQg8C6OSTi9XHqqvKn
8oxjdxIEwtzqGPbX3LUZNQWmGJurFZRCupXp20tkGzhaSB/2RGUS4c47y8cB3fT5
F0I8F/ga7HIZ/ZPczXngo5vrKvKXTr2S4pvWMVpMhMxcE1IBW3GmDKDmf6JLTVNt
Ya9/uxlnJ7ubBhkpMOMROaC0ECLtXO9lBtSa0h4w+oSEBNQZWRljLSXcadpUM3Bv
JOa0Lk356vAFvwHV6stW09VRlMdcjOAb3NPC/9mm1TUIUTutIKHbH1uIwO2BKpFA
O1Jm+GJg1WLhS1hJFVmPs+vh6YtHN4OQjDHBPQji2UcL4tdj/w6LNvyU6etd2TEI
vZDuFrdFSupIhhGRR0IyIEi7hmYdmZR1h4L1fWPvqQEkfIHsfzWP45TMoaL4/reR
CDEkDE+mFhmbVdYBiIEe2EbDxxCV1mh7B0bGlpkyYWwczDLSJVOOVG5yicyf8+Q1
ex6DHH1EMQly/MyhC+qkWkRrgrnnRQ3cVFevk+bOPY3SRKI5UhkMChM7H88gaEpZ
vdVecjIMdU/ru82r4USJexHJqDSPRiZrNC32rG+BXr1/+eLlQgaZM3S5zhgecPKk
5cmECDWwjhaQpVKk8rHsCjejSIhEodl8Tcrhs7P7vUr+JRZyyCXKW0wMhsRlNo41
u8tAvTMKXIdHWIqXisus9mxaYI4bd68zMjQeMqJbNyQuz6Y4bJDkKzAUrLPZ7x66
DDdesACrwSasKaZLqzsJ8hnIrm5AH2lCZvopxCfWa0GaVKD05Gp+gg+fvnPfvZnu
vss3OWIqZg1Jsf06f/A4T1I3E7Ia5E7P/BP68rrsCp6L8Dkdj1vzHJkLeUmJJi+X
lIFZON42ToVyI5Uq7cUZKNAK0Q0hBxjultM5czZQYCkOVfxTLj3h09CC6xlKaXo0
nQjZnzqxI6GgDTGFLjzTUDGON3mL6pMFUnhoFGFVvEh3sNMR9MRNNA3KQrCt6AkL
ySNshPW9FCu84xuSu4abEUbFTIIZ58Qb5Yv01lqbivBurT8Lqks32Yu6TXcyIOmA
4jjZju+7ZvypOR0gZEk0MxBecz1xPgGEeXPOODoZd6+W3PC76OuiN0eC/KZ2OLK+
OtScdw9u90PI+iFihWPQKaWU8aWnGtaqi1a0O7IKuuqIGdat6F7N49k9yzKiAWEe
6Kagy9DCI+sEaDSnYbIOBudNXqNVG98Z/bjSNfvw9TT/QI3v43gFCwx+XuIS1CEr
b6AHZNvQVNbbMIAbpwllp8Bb3weJQgjFd85HwxN3ciQ3dxFp7Npzk2zGZGyIayRh
CdVaEf+scEhCsr0x1ZdNy4UHLfKOjuSH6VfUUV9Fzi1TJ7yUfy8j7RSzbfOIN2+C
rvOosasGoPu21H1AEnWkCqZ/Tkl5ACf0IActMWkFdlZAPWIUz8RqDHih5jIExQ+O
I1O9COF18zJQjQRDSV72bg2kAokr5XoZVMyTTnnlGDGtnyMkifp151Qci3Xkmykb
B5sgv51zS1ypf2kgNLsBhTKHr+l8V3yrpUTqCagCzoEdO3gGT3hGppDe9C/3UQZ3
q2Q6Vi/VCuvcM/4WwPIWKnYEM99lxVN4uNv8d0ySvTM2V5o+DlgDr1LCa0JquBKH
Ouj0B/stzwc3g+lefPaAUN3qWFMO9LKJXln6CRIa4QNso+PO2yLPL6oaOUgn/a2t
MmELQj6RpvBn8r6Bqyc6XRnb6UYFuw2mn/M1nXRelZ2SypIBHbsiMm4PaKxxQ1uy
t2n3qZBVU612JrTP//JINZPilVyosfuFSTjdTBuItSUfDRPISdR0EnZ6yfEKInjR
z7WqwTLzy9zYwv+6bJYciRSjSi1O5b2jBSpxkx954KbBXlnTapZ95gzuA0LFh1gF
Rdq+yRWE1X8rmwr1CwPr9DOWuv8Y7GdUMJ5QHg4Uj1FJ09eYd3dGh1YEC/4eQES9
0MULrGrZ7VBwel87ElPVg5TzPJS+VkUBw6/pAXsHpLdLEAqbQvGon2f0s0ap2WFn
H8gIrXUvrEeLsmqUDu1mG5cwWGh7ZKAuPGmA36DsgwUxZLN4ROS2hSma80+PeHL0
p1y2WmxWfaS49llWzGZH0b2zDCvOlOX+Nb8GnEh8CJa7odWBOUSI3LynoUVChxBv
lqZ95UmoOWhV5zajmlJOnK8qT5CzBr3m+aIWLmwZ1TQxxkh+ilee7EwuyBgHTwEb
FunJ5eynWIWhZLxLajjABMAthv28zTIY3CX8wnxvBVtMIK2DGbFVm78S/yDm8LAj
vzYEdrfKD+j98rhLe+6ScIQFubCdN/YxyewFczwlxv4v8+Fkj/4R8ha+j1G5jTD+
1VpcrJffza4CCyKdEsP44v5o1c3dY+g5ztE/1FX6/fo5bHnl9tNnVELhaFmOjcAh
6dY4GLPO5PHhpRkO3xiyBu7L2FpAcI+OYaDUiNrUZ1G+1wNH28QZJiU/JXCMZ/7P
XVnbm1KxG1339uquA3CGvT7Q9tqc0srdyVS1VdzkWlnku/x4kUizCuFQQegWhBV/
CZPy3RliEko02+sDUQf+6Drbtxw8TSzPx34k2+56voqAGvQ9O5tahyTTbaObrEvv
L4zdLC6ovv6mwdmBzMVZfJFncJJJZ3HBl44HFsOIqn2cJI28V6QfURmSbMq2fRIL
sNtYCdfHnWhDS7njkLUG/SEmj59cgqQoUvRJNOr/fn9AhfZjNxwTAF0FNPtpd29m
dVnvSQVuKd3JpQQUKGgQYCaCz6iBzrKBoupckq5WFAzZG6v/0JvUxy0D7WVsREhK
YgvCxp+ObpxR8lzUQ0EM0rDl6d9RjrAeB5EBrvg7UoH13nG7rTGUcl+16q6eFqBQ
in6RnD/RaN+UnaTZ/GKclUjTsbzkShV0+A1meq+Y/lrB4fid5BjuAxtx4LqHU7Dt
zU0CowbuVhM7kYGnv/XXqEV7FheP2C9YRfjvGuEzaHwE0gaAwfgPUINr8M/PgTkc
WN5QcF/iZJ2+RNe6yvFzGqBrUmZ2vUg9Lm7KjHuEktFoinuHHNRRT5iS77eSCIgN
RDf2xKN4zKgdtOfUuw5JBe3YADBI89WpK7kCGwR6p+xufoj6Y1fvsDeQxCDNVwuR
areEqKhEgH+jb0jCEae2HwVcDygkjnAcMgWVOqYRk0eF1SWrbv4ps4ShQ8oJIVxf
FKvLsb32YKZlWCRSwbNRlM+lUfX8krDGrbpGyMuPTACorrvdR36scfcn7XGm0SQB
ypNmqMa21fb5JGaRrCzrBH1gNN2w7wQKmoevpWcnhsw4+vuIQl7PIYn9kZnM6IFE
6uJT5HMdJLkSHEjHLhHKunG+pTOa6cQrPn610KFYE4NCXBJilyyVAmEjTIm6Mp0e
1rA/wJC+B7PrPY2kK4RO0KglEz1nqy7C7Mn4Pn7AH5SfO6ZKiUVEP8vP1VgjMDJs
GBamJxk+EBmBOL4v3457uxbLKy4j7g7IpcphdFWcAs6aZ9nY8J2FKiBFw0Y5xUa4
hXY4pS5PM//LT/BqsnuDLRf/2hWYeIAz8kCgHAgaLtbP3B2YoC/3PCSoHccBQqCk
Xhv71VaBV1ZVMYMUbbaigxbPEFf/s688uMqhIOkaFSGle4Q94kJ0ifcy/w5luZmG
+vO10ZlbRVBNmSFr6bZUM254HKCo2Irsc4EUYqWaFLVWZK5G5dB1aD+W+ad+ZzyE
D/Pz7+OPNPXs5gpK8hlfgkm00n1sor1BVChRSpPQKIZrXK2vIs0+zFBhWgP9lYoi
8kM4+PaUbxVnsVAzOQBmyp1krlmPv6YDL0SFsRIhOM/OmTcK5Ce41DcNo8mL/HVs
q/vGAnYbqXeAdlt0e54UyESTbr0wgLrrxiOQQUhBUOKda2H5WgQb+ryEjt31UyJN
xVNKkVC/V3sDZpP3p4o91pkSHABAZ307p+fyHtopZ9EpQMIlSW/OLXOrw8d5g8VC
9KHOKSvti7etkpk5DhkBeYmveAizvB8qS4v3Hu3uHbIc3lb1TfrDmr4uZGZTVFXw
RUnDzMiTEKl0bIadkpSpgAc5Sn7mGB8bwZNg9fdqVye4uhfuVjMJ4b/TBXxCZpkl
UAHJ+fw5lhK3Y4G0GxV1CyZIm1SKbp26noT8rWzWhLNwPAcD4aVg5SjQmAe/Xj1M
2XTeI2gS0QQ4HQiqfIz/bJF+QM3vyRvxzt8gGy8CEsZ6cRtYPrFRlBOhkR7xos0o
woSGK2hfH4a3ejkEytcWr7Lm+JeOnSSybArz6V0BvA4NvLqf1FktHOZQzIt6Pn3x
mdLcevEqOsEiQVjZyJ5wHq/k0Q2YkGVa4U3wPS5ekP9OF4YI6L+b6Yo4DmyXqOoU
4apF9k2SZbGjjeE0Bgvb6SjsC6z2vRzu9oDnK/c/Zq1PgMBLmap2oleE/DQVTquO
nMqwL3xZoi5WQ80t0mbTWQNvsT1/yf4HbzSUHRuy+OWhHOIwzd46nF3DXDsSDTxG
c6MHi3Zxtm/T3PJW5n553/vgEhrdytutrOtrFLlJSULM7Orqf5q8v2/N58UDNoYm
BXpUwBi/IKxMlKkm3uZH8wffreorcNe/d25/lpfGHPriPRGDq+A6pElnNMoC9uyB
08PzkZlHEp76MrF7AI5ja2C1ydu9lskYXs7A4sGgMRWOQo1rrIWRMc46vrSaO5Ed
qdQDE4cP2FGaLYYscvzY71E/g1UDsy1ZK6aIVn3m3D8yAbaL99/RJ6OcD3r7kstl
gAam4EMoCSMBou36JI0PwVjNTImzBJuiLwGcCQdrSFbUBxYojl1z1CjgSpsh9yTE
SsnnIIcDI3D5l74XxtIF4iNgo7gTrQfZGUtyDoMe6G6XELc/Fpu4B5Y4qduh4VpB
RikcJXoO+cdx6Z6ogOFGS97jalJMJLXPb/ubykz4ojFFPcR7ZJH0rKaxUe8bx31/
6shWimLvpUQ8zmjlRjdDthjBceqt747SX7ZF9SL9IpVUfO54TC/fgqngN68h12SA
Q6o9C2jKJq1KYHzQJ9pdWG/VD9RecBtoMVkcJyQHv+txBlnXp3TqoTb4nRrJD6sW
WMENzkBEKVXdYKf3RdL5gnmdjSsEZYrzyWLDHnr//hkot13864ChncyKO7q2ZjFH
swFjh2EY6sDKGVA06SU4iT0DECNwrcCm4Jj2vKe3IVTR+m1vQ324DMvJoVlK7DbR
9vQAEyHWUAOx2Uvhq1YJS7ZCyNHf/2Z3iSTOAjlW5ttwLvtwdzR0SsMogDGVcAGe
00gc0ZNZZHQC8b9qUdKZuCP4Tgf0e/bewXOzHF7+dyf3cVQxUSL2ZB2fBzoz/cHu
ejypzTZ//JaRSQqLNQSrqvMzrdoWSuZAtkL+DkFR3mkEXU6JJB5YXQGhcZ7XJY6Q
gqLVOODLc45Zv9qmp7yjF4DA5l8DABlzpC8LndnHjeimmQ0rthxERGULW1QfaT8k
fTF5YUk8SZgxnKm60FHEL4XBqbq1adaUb+/MT1SzjOPrYzrvrbKlrGzuk1VA/pv2
qtYdWmcOVaiaOkewgrmzEY6bCHxdOqavoYkymZkUkWnXmjtNrjLpzTyQCtLc9Xfi
UzWpvNJ/guQ3pHoTcM8/ITxAAmRujhtR/vqJENYDo2k+XeWjFhVGRfruvdFniC7P
a1DRIHAioDB1EzEAgdBNALfVQpw1OZsgtJ/X8FHDudJ+OJKxMOROaU44TVK5jmFn
ZctitrcBx12K5g10AJ7p7prvCybBpcG3drBoDUBXPzMoWgOTybXLIPTWGxeV3nMF
ca8TDzcYhyUpGsexct/wfYGH7qhGDxq0Pjm8IlUoMp/qckpNb6JUn3/G5O5gfw6a
s9uxPIqLCrFhlCYjfSDQq6c0qxe8YyZy7BH9vhobKMY0XqRDdOb+GXb8jjvneh/c
PLkbwYLrVeRA4hswZcXaHpGeMjDW2wrG7r3pgdXeMBgai2HOjFYxb7LY/ZpKtMtm
a5BDihBsg2fq9rGU/a1aplGBC4mY3NG01whIfdAPkQ9NDNH8GBEAmAJIkOCjIKBN
EBj//UyIgt7ou5bNW6GIgBL10zkNes5AEO3Q5ixX3bLf3ByISBRSUvhTSr607z54
RbCnF+bHYnDZ/BULuauj+tLGk9qAqdp2HKir9e6gzSRhYjf1ZcOBWHLLVbeQJEyw
u9DF2BeEMtvmObMcDB6ize7zsClg9/pq2Qk2jRVHPTCB0ElRcoq7pnWlCsTwnPmr
rl+ASe/kV/+IBqcMQDz3hvgVUow8DuCKSInxabNsFEyUOxKtzv7TWjPy0BL1NCrl
A00DJh4Df2vPfL+FRBqef6UasT8JP1EXjhBYSzgRb4mY1Z9q4b2pynajlYd5Lk3b
51SA8kXYvUScX2uElNfKbm7BqiMdLxTul/lY0r7NL9gh/0itS80B22TaN+PBHmjc
1Ms6HooBKsKurJfq6i5CsbVLoUFr47WZQHCzhObFb4lvrys3V3H9LuKiVYGz7Kr8
tiZ8vZQ2ka5HizvU4k2g0fQZjhXy+6Gnum/B9Gj4JyMRF5Mo6qqqOp/cDuLWLkUk
vmN+J1ONsv+iwk0VBqFM6BPjiUhrYvozxREEco+kD4WtbJla4q0nmsqp7AQWa4xN
9PkM9A93GQsqxdawf/dmP8K6IhFhG6cTvwTAkAlmkvKZdYJh5TlDasl9qqDTKW1g
8hX1+T7H6BL9je3icpUMumiH4rSy2I03BYEXFu4Y5MeQDPeVPIlql53BBwfvEIRH
4CmJIvTEZFBN5yF8Dj6sDCEc7KfH7XAvm3NgJSTZcZ2g/eGygmzVWBWSmgYYg8Po
LrARqUJPuAzo0MnncM26ZW4prefHuL/m+/WA6SMJBapSPQqDfOoz6+nFq+wZcARA
wqzBEHX4ybZBZSk5V95Byv/gQcDAjCao6EYVOOkTkheI6HFOA6eS4l0L4BEO5bHg
KtN1OCJFl79LbzGMPPrZE5ya19neeMKKB2neOp8Y51Pqs5aXpubyuWKcaUE0Vp01
qUwO/eZwacbkwG3a3LOdCrQw02MhR2piCJiLuD5Ewe8lht8SMEzccM2yRU7L0te2
/VCnlj4rLTPVf8hFADzqLb0tCc5AyXHLl2BnqsO6h8VreAfae6lst3Gdz7TxLH/q
hM5/qJ9mlo6ApM0dN7g0/tu3uUcd9SjZ2q/r3d+HSlGIJGSIax2zz9nx9YhG9a9U
bI+ijgcnWy38SKPdejo4/9kPUbZdNVbsf348XcXr3Zz3SUapum9YwS4ylg2Nulle
Z3W4G5KfvpoQhk+hce/4fc+DGWw2apVq4XAZeXq7HWZYHCe9HnalrwC6hR28Ne5T
zj/CY0AECbQuw6T6FvLyj3P3yu4yYhypmFSdpoR5QaIoqpdsea5JrwBhwmxggLNx
QcSsE4sVu16u15c+8aaUofHz1MuGBOdanXi72f/yHkVvaM5T60dOuJde1/RU1ola
s4/+8M36VOLVQt8epqFunymeP9Ohl9pF9GnrWPdD679Rkd9YhqQp+GNoaYed0hqj
iOw1PH9NxNJ/MYnQXBhOWAU5HZnyBX1a24cpIrGhlzAwl08GKrjFngFppGqrChai
2l2BapRpM0mAmt1BARH4ue//OIFOZC0caQDkOXaQV0fkJWojZdWoKuDWY1VKDIkx
H35Sag0P3Kt1moIM21LN+Ft8CphuVqCTkglKGyJG8Yuc2WT3/JZ4C51rZMb5+e9n
trtGaNeaaGZplZ5Mc/MxOD8Wz/rjdVI3XlcDsLXPy8D4sOjPRrheL9yIn27pjTT6
qfuJw7/Wvi3QilgQmhLC0/u2eSRLyXsb1tWZjkMNOEO93MrlOcsnn6saf6URnO5D
jOuIac4aOZ6/DcYfnq+3xyiXBffnQVTGz8YE4El6qTk8pbLAUpDrQULQKyHknLdT
DoGMAt8mq1QBX6HjmyiIMBce46l57X4dypCMn9tBZMqsxov/Tqg9gaPVPQ+MYj87
PsY26AC2r6lvlomLWhGEVTQ2nARnsYDFdZUbRLITGx8AoOR0T68828i6lc/XXGXk
acAEHJOm97t/EkwR+32nNzv6UH8eY2zHgcBUUFQJfkwfWqPyIXFhWqNjMTxVFrpL
kvUICHcPv1g4dISE49KNFY4PbgmqECMC6dH4AjHvF8nwjrnIP21qUu40Vu0/pANS
v6sc8tgq3vG2hNPF7qMUuIpyvdzj5u4bWo5V6NupWk1MkGyIIy4AA0GmddzO8/9m
DF597gTGINV/RkwA8VgmJsg7xIjSq2ftiV9kucrsN71AYclWr31RwN6ocV0sBNFt
yL9jnndmgv+Xw9k9kan64/TX2LWE/Gqv9Hos87+byl9vmCIP3i4iG4GktcWJoUAX
YcoxmXm8XK63+agGRG9uNJ97JeM+mZfMqXkwJ1KwYJJ2R8u21JzFb8TP3N7jSdra
icO9p5qy0bu21gggfutdMHCBqCLFe/jGz2hFdHVZ0zz8SVisGh0S/yOHVvuavVLW
e/gKRoyQuPfatcIYBbaYGqaH8TIJK3eeqRzGAe618pNpHG4R7p6EOzyfyWTs7jXf
t1vFBK3vaWOgwMV0CWApjxo4p56+olepyDW4VtF8PIYEJsvxi8mv5bUNuCKP/vfg
b0k/Ebo7zuMM6pyvUh2b1WTb5ulX3V90zoqMvzvrq+TGWiZxm530iYsFgoKSfPyR
enAKA1WV69PEov3sgUR8TkG9Iid+ACBFeQ94MurXoaUfrvD28yxllS+nzm8nlVGh
qvGswwS/PBc/ZH4xSU1d8xbladzOdvg+Vreooc2EKdYTfO2DPbcatFolHyYUJXW4
gu+Ku2VmJ16LoDZPat0wf4bZeEKjs9ZHEHVICJX830l/hRyNbm6f4TJ0YkA7CJea
psY/U0ca3fPhaVhiQ3KjFBmiwA0J6yOJCWPZNDQaz3uZ5c/Xp9WJB3LAThJ5mAdm
zqrwLQYYF6WBx9CjIegt4bpPCkQHQDIm2p13viVvcU4tcMi/RRfOJdgC49t5AfFh
00QIYMgBu46skqIRGAn//hE7LpEiUMULBnKLzSfzXXpTf6SucQilhupSTeOU35nE
72oYRJCnQ1PGbx2ky3zw9yx2K78CZ16BGrpaZXx2by9DiC3838n2tLX/V9U9iKMi
nIeWhU3sE6y9KOXxSMz2YOnYEQc0GowgSRVsmnhARM26JWpoFC6y7ynlryBJI2I4
jfm0H8nTFzf3sGsWGMxz20EqNSq49epKMbpz2e8QJY5YpXjjpeIZOWeMf5u3n4h2
XfB3o6R+XuJJKta8jdSLZhJb2cxNJ+MSKIRSKPhR/SU/b4C8nsX6V2j9T4srEXby
DV4Pv4bAxJk+WF2a3ZPcYYibWA/KSnQhlWvqSmF+vaQUk2iRceJZPjhqZGrbQQxW
UzrQkM42JNgrOYCqa+pw3dEuNbCEOLGFQYEuJvr9vNC1tF/pQ4Y23I4xDr1azyoY
Bf7SOTXDNVKhcEfClBTNDCU58pSgMJ8W4tM1npnBCoqCLy+a1w4KzfeEaLnl0UQT
+Q7gsPV7Pt/O2iNNEpyeIUCLwgvNn5hLFuInjh6GteVU62KvjmnsLAMyFbiEJDhf
19S4yGOnXBF356Gbe1bR//tJf9t7QpxQMB5V6DemNiMT23VtnkQ4nko/p9iZk5BK
vvj/CgGASXq+mjSgVcjJxETVAEml8DfPzlcf41FgUbTrHm04xXyClfQ4AggOXMrr
37G+m9Ndzc5IKi3vseDy85XfMaIEB6QpfFx+JivsnVTexQl/Syr4aJ1MjLR3cW7J
zyCmSmmgiErrsk05v3gDXVPt4tH7Qbsufj9NcmhOkG94SPmdil76fauMjMpfLomz
8ZKUbzY1s+Lc7HIMT8j7l5ZqJmO3yjXxghC4Eaei2cOIBcF7GsWxXTk3mfcXNiLS
tqoV0DKm7sXwy4o7zr/8UNU+oHZsdi2n0s376py+p/Zm76DFPs0asJdvBlegMpAR
S0NhXjQNDEW+Cdq9m7OFrcHi34Zb+y5CosJrMf24xj0trp2Fpw8bRqBAksRgbndS
shMQAGdPlsiSrV6IEoLpaWXnUNATMMoxerZ4VujrfgD7o/DzxAVr9qLDxCgvPkan
8No4GAGKP5fjrpmbbJkKExMgSuaahU41iZpG6XlYg7ANb+OrR6Rj8mP2Nrx614l4
e+OvjyT45rAvTMUtrAS7p7kY3PSpcuJXyDoWTnBwkw82ApFD3JBLEzyg/kD3FnK/
xIsuBMFmQRbv+CtAh0WN05No7zD0q269SHeGgUZ99Kv4HiI/8ch/i6deJVTn+Bhs
TAepjF1rFnZTmsJ9p05shEbwIgEAhv5Im5z9gMxcgG7ByOktxcVUzPuivB0DTgiD
yW2eB7j29x92E9D4r2UkB96VV6t1Iv74watDsvWfHHYn/A3TWRZIWjbIDGpRRXcL
z12ayIU4F2OJ+OnlEDn1uRHcJEZdwCCZjhmgkH1z9zMudcmnf/N7aTfu0BIGky66
5s//VX9pHSx/70MS9kCYUanU9YN9ST0y/iUimY0+3nCu6FILwYA0nfEZ1iu57Okt
FfHDp7aXoGk0O0ToVLRgstOJiVPMQ9GIgpoLzXUuLIH3h9mTMipHWBZAhLT04Dol
QWvPKWg6QkI7VWLxerDsaGnhekCdlLP2nT/Qiw2hgKmNfgi+tkAA5Av1q/0OHo5l
fxzsq39/Qup0NovjefLp/HnQBnnjM0HKty5Xgl8ef23dh7ire4piLrsY3ikjrmDt
dxn2cQdLgpH8oFsTbx9023Hp2JPggXN6t1M5wB4+aO5FK6MN284HzAaABdFcNBwI
ET5XY8ALxiTMw1rjSW/lYT8pSets3JN58kfohEKc+KejsmWf6HhPxS6h1wHsEiph
05sBmpaV73QR8MoPt9pt6UPGZHzmnXad2v4rfceHBVLvfaOS6Os1q+xoR0ALn2Cb
tQ1TtOpDtXiaC2bv0TvzGFKmVqnuwG+Z+Pu+Y2c3rYdHN8+/YoPscIFop+aNRX7K
8fOjCQYR8x61ztGwkYOjdJcK6JGNLtKJ8HL4AUtKpUG/PftdaikkiT8QnI/q9xAL
x8KnSY16WSDxP61EJMhaHK4yPZRU1PIn3rXsE1jvczBuAhJd6Ov9iUzISbi5Sx77
vZvr/1ml4Ng/e2qBIkNl0l1IQI3goq6fcXUT8NpRexkImDmvXbe4uHQ4AUjTiUe2
8zivIqzMZVNrrHSwzJtGZOnktndHxg/DhRh9RQrwRiR3L19sShETXx/UDMEcxnci
i+EYQcjrXp5/BVwPY0O7HAZh82hdOf202TG2ApT7a9favlxq0cLlyBR5PSZaSeOP
PcGqFnXzOlVB+Et/7Nl3IhD6o3Saq8hdmHssiIfk+U523AMBgnMmriNmq/+yh/Ow
GYypkW9Ks6cwIYWulek5dqyFQXpAK8Kyr85zO2Yu68iyjtiPPkPmO4/HjrwmXYRP
SQwHPHIG067O2Btymtfj4cl2vxi9n1zPuNVQ8LwR/Q3JDXBVWE/ALtjm0NixbO8N
nlt50CvwngGQDHanrn0oG6NYidP6AbmraJUWCboOXCGBJS1rN1ne2XuHV86MvOzd
qwK2BZLb6pMYsXqkARYhZ1Ej/mSTsNHFpgaAjwogzF7Zc7HcaIRPLlCTmiKK/eJp
TKIGvmcOFDBHyIfo5uglXVPDr5Jvh9nnLt70o3Px9OCxXqvmCoDF4PkZNaYlIGKW
mB0F/Vtm1f7fW0taXV4vDgoE6FgUQxJWviKx79R1eCyfXW+OB/jwz3+CT+hmqF7M
LnAissAi+en3AVNik3S559jT/Rw890YmUpVEz8iLEuBkTMaorvJhYlgfmSOLjdDV
hGlC8/Vvw1OksKq2FSucqzwk3TenJTjvAaIMU3TS0aSOCcaCFxbhrwSDB1b1PkU3
YgbSg+38m83e1dwPMBLoDEUmeTj47mm78KBE3/OWXFsLi/1xnxCpzEtLcfsleOx2
3CbWE+YoQ4cok7G699O3twX+v1KhC+/ZkkhtaFtwobSaeVax4uTETBCmDYn82eoS
ngDXElNHpKiu0x7GVxfOUyBfHYx4cxRQBy6bK/W7GpPjj9MQbvmVTEBVf+kFHbDA
Yf28SbQpn1zPYNx8Dr6bCVxApbfxPiO9RTxHiLaUb3lCcPdRwv2QpicZ113Jho7a
5Qn5vvuZQazKIHlqctvgzwZQGgcfxVsfVVhfzpDY8zysahXKU0Hb17+j5f0ZprSy
Jg1YksDe/bZxXiXm3HM144BHYKk9IIXLbR0FGILHPxnGwhMC7rofqpQVTRsbRfJr
H8exDqiucfs5tWVrYiGzVcCh1SZmqtBgEgyQWf+l+R/RvT2XachfqGYT0Dq1yWqy
pbc8wCou8r+/htXkfGUWyXSO/SIV8oUT109uVrRBT9BUMT6BMcxFPCOwNzKrw+js
y638auFdqw11oAKKqSRWd67DRd/F2JstfbcU3wNfiJ+T9PitucryFu8R6q7zG20f
4wJ8f+jXQyU75VbzEJyINIq1FajeCKftrV8Errh1PeT3qNU9gp0lnR5z85KQk2Eo
2WbVpTXkJ8kfnFuej0+AB4DkjxgCyB+gJT+9DXHLQ+HeXd/lhsqECwMsKTfZoBIg
gfUmHOxty+f2gPaff4KFUGdmdPQdGmG47nW/HNidkox37iYaysBa0mVk9MSDHpVj
s52faE5Kq7vPSG76gxFqOqCgfWKlH3XmQ50ZNztNDScvPtEWpsbeNnHVePw8NYeh
HfPaYz/nmFzBBQ1oV64DFEgSwe8p/tQfwlnHt7uiSgtz0K+VGz4vM6XmRiYvHRBE
nNeKgyhotrLbEFWb1ryP6ppZ65oy+xprYAAOvd/WRbEn5glwWzKEqVeAUXvsjUV7
gnSMx5yoD5HGy2DVClnVtWDucWF1yIUnNqpOIQkifr8lEMs+z+qK3648JVJSQVts
s/7dCblsJ8QYu2QvUDslM1CzMJ/6czTfBFD/F5iiwBnXxPPoK82WSxoPxoZJ40E2
uhKnQX/goIHohGUAQl9DcIyyp2uP33S2vxcwxUdHQcqgxNTp8f/GbnxJE/4JuEjV
q58udqEGK/6Q6vVClh3FayHLaZOxiKFYloeFFWbSF+mgaylilHD2ocaK5lcMQDwI
971AAZtGjFnp8LTl1Dn077/i35QC71RTeIcRnaMincaJ2Ffuk4i34h2EOVJlBcHg
7/XhVDbA+aN10fuWF1ypZJucOXKHhLmwrd+Jh1uCjL7GdIK+MFNZiBVySzsqzSj0
Zc6AiQIrXpWBQDPuExXHkRzmuvkVumhFVS9ofxJGMQLD73Oi4sA+pTYbroFSDQWU
2Nbr/ilI/smOKZdrQwEpUdleeXhstsT3CuQ1oEpNG4B40Hvpo3BkJ88cEa8ul/la
nZMF0YbTH4/OfwOGOIlDHYw03OxmWQofj/KngpzKkIqFM7OgK/5d9GtzZKWzk+ea
0AUyBD0K2bwG04lY6MdqiaAubTGCezarx0MYzXakYWH53lq1Hhotk9+IrmRXU+HT
pNzaIqacXyrw7X9nhYHI9FzA0CrfZ1V+ln8xn2Nc6vgeqxS9VjIZOwgse4R7RlJ+
ux8HWHqDnGZL4UKhc+HcSkZtM0v4php0hRJAJ80oyblxu5f4+zbfrd5hqRfDFwnX
6YQpQCTCKkksH3lf+Oijw5wATz7Ih0eBXDnr7y8mVPmGLObLoh36MH7ODH73EJGs
YFK6FdeacVkNL+Y5J3852mQQAYxVCCYowyVr7ZVV9ZqTwN0Y/UFciuhgRr4hwKSy
GcjgjV4krUluxkQBAIpPkG1by02MhryQAvtcPnXpoNVuaSHEfetMKGsjIado0O7o
HrXCbDEwMDCQdRavchhE/Hf16rfb663d3qL4jK18zxWmYPQEW2r41NLm56LM/PZX
y1lcMqORGnCs2q0w+eziiMnW6cIfkRDe+ceyw3c7GM0QBChUx3+ohFPL2siGgNIr
520SYmh/+Xm2EI5f/zZ+0+rzJ9t8v8AD5Ujos0Lvdi/jjkSL19ey1/GOx1/FgbnO
vzcDWWWD76irHU4pn+ZmogzOyOCR7f+5dI11FyhcCQHp1L4Jy9YCaRgnib64CGeE
JCZ58AEDZKp93NKEYkovTxBF6TACGyVYCCMNvSy6JYqqsjgBw7lYS2uVSiQasVxG
oOhahpZybuyg0+2swOq/KyGBUhKvQ4zeq1z3SLL0w5CTGmhBvGL2SwEaYNf401DT
wrZRmcgnRdeYKGXDMSPWbA8FJcX3xvUC0T+RUL7I0CB3usd8bznV2zM1+xRYcC9P
15sdkj7KNAUdRHeeJ7SQKtRzH45otnnPXglCNYMiUXZIrdPDmhJ6XMktqp+b59Zs
Ba7fupGwq87cG1uuRyOynWVwxrl6NcLpCw4CBfYAcrdYXFPeC9rxlJqqcMX9LzTJ
wt//kdb/b4KKCi0XxQxCMSGQYEZlT/wTLYMH4A1fdVEs7CLFUqXPBl+YqXlaru0J
zQ5rT+siyrDzdpG6f+/AXB3cDJ4bRyc9E7pzcPAeKNK8blT5+iCby/bY1yaA2A2p
mi0Z47S5liZOeSEEx8TKd6xeo0IZhSrdnTC14c2/jnpExzs+88JjawhfqNv1YnUN
MPFH1RC0+vypfNn7VIvw4nM27ckvczpxTVs9anTG5obhCOMsupubdGiPII0m+BLM
7mN7rtrjzJQz6e1pvSNTGRKNFXdQV2v2vFw5xHYOhI/gv+TcX10/4QsXXn/eGLt6
nfJxJ8EMDyCAA6ndqDJqxNmh5c2NyXZYrhavzVrQqzzl7vrZNyzeA88U0xYKCV9+
6lU8Bqoj/4IvO0SwNWt+HIKsFA/mMUCaP1nX4Uf/7l/BzgVbzTRLH2WmOfQNxl4l
LZ5JsiYpCUJAwrMIaV36BQvk5d1lfw4Lk5J49RSgl9UJztQVcLu2lhCHaFsl/UDQ
L8uadvp9ixfIXnL8TYBVDPypjEVfDwGm09qlZf2TIz5yuACEssaHGew9ZT7vJZbD
HZV3i6rvzJk2OIMSDapb2u5biI9OkSkF/DKrwnLdl5tO+IMdDSdeljr1G6m15L8P
BseoCY+CpBJ/mnC5gVAshOBrlR6LnlMKr67zWQOFNLJochyOvv0ggIocUjrXOHMl
bY/0MhBUtEhyuxplTR/GyIUaE78mIzdM5qJXQ4LOG5kLLirGdJ4LC5nNOCwKqI2D
/cxF+4rIbGN6IhNEgR7XlIcvGr3zhaHILBkoB7TAl1XWUqIyuxW1TktKLHP1AGW0
mFvGxIK62W/Vtqpe7gKfuKa06CZOeVluo8gPbmBPZ8VgmHRXyNoBbHX5REAq+Opd
idkYcRLrJYg6aupTXY68nwShfPTCb9V1XLBTsFBYABz9vreURhN592ZU6H1io/k/
Rg2slsMJSES0omrhS6faMxfdv2k4aLMBfq/5c1A0i4c6KSHkKSybrxCahEojwMWR
felsjBEUVskq4rG1Zj4NiPvz8rtI1COM96+a7PrB9xrU717xzmKSpPgncBRVdt81
ChIdhPPU0C/Ot172sCrDA6/KzfP20bhEXq1/nlKoKyJjiQK6B8N+BgWyjT/ImJBO
Gdd3tqye2HXMLYCnMXBPtKvS5/mVlyy3KSxwIfsLR/75vEm6XRbIcqz5y4j63WrD
Tv/3pJNmqpnH/p9E+yMczW1mOGWSxjqzuwvw8OZ3Jry+5oPQl4Mx/gHXtu3f4I0T
W/yqQTfBlZdfhAiUwGmm7ndlOfC6IXcIVTdlGT61IJ7B2mI+Qt6Wj5II3sgEbLv+
wKg/xT4/++tm6JG+q3J0UqPt+Y3ZAWE7kZqFTeSPJBxVy9Fypjpj+Nd3kUhtHx8z
SKDuVl+Pt98A0BKJDXgGmFNYp2b/tgDijDZxaYL7LT7KTs7T4j1IrbVqWYtDogUu
xEtOJzw4+hezdAq7SLR5ihYlR8LfZNV3VbsZmdqqqg47BA0jzL6M1ARe6fcOM9Xe
hyO1LvxdoG3KMx/Np9+s8dEDBtLtD+pYC8oelxgsJsLGKPFNVdxn/qrTIqYYcIZ0
8oUjRSkU9qIgqD6uRcN9XCTuiLUlxAcreOhN+ki1p4jOlVWqux/jJQduooZExrW5
oIWkpkI4fG7wSDjC2TIsGN0N8egq+dayIlTX3NO0RHTt81RcJyaKyT1GZLvWfQCe
9BpIZ2As6oT9mBV7+lkXQvVV3683ubCh1te0cDEyCjgWiNxukrxIlEt0LQ2K8QzI
dNqArNuueAngDB2eWAIu2WcPNSAkA4/AgALARGTSdnZrIOGf3fFxzGMLQVC7b2u4
/eUimqo767nJxJ4gRJkvpKacLXrd1Tp6gKzbDtKIN4/fSSAJeg89nz9kDEYcSr7R
qcU1kufwbtw0xxq4RRR49BLH2i/ARCyhFR5nHQ++OTk7BDqNndhaklm7kMySeodm
i4USQcf+2/zADqOaAzEpBVwjEqUymr8cvNBAL31pMNdWuots0QPO8swxYvTqzC1A
MGuTj134few0ulSWLo1nY8Yr3WbEfUydkm2bWtBhm/P9gCKN8n+B8Z8zYli2oUve
pEEJ4+ANOAvOGJ+jpJAsfy7hj3eNa0coSIvHf0MkKQ5vZNR4IgCWyALtdmWsZ8yS
8Og26Xj4VrypTW9ktCfsksfSwPq8kS49pEsk9BqRFCqVBL7BGO21OZCTzY6ZEnqU
vy9SKEPrBXi+ts0MgV7cerLXaR6i9G/hLvNDHsc/YIirz3gd6MG6CKIBGnrfmj4+
H45YAnUblLABxOgV5oMWHANnCxrm/bu/UxPFr0Z4nTo1vC2/unwhkWMP+gICBo4N
s3kw+b0SxsbNBMpNP2hkCfNSvww3/UDVGsP+O6zdzbiCLCQykeuEV5adpDYlUko4
3jMiPH127avJ9/1NM8zEWmOqDQuPm8Prfg+XSYE/6ed2ldRUkrX5uGWnWy91W1ty
BiyyhM+iLPzU2MjJjJyX261O2oS4CrGn52Dbsd/b7yMjCg5TL9BGk7P5UItrqmqX
VtwSIg3dE5Ukqpl7H2UhCTYoSPzcWyzgD50li1Vd31hdeAEv6Kcj/plvEq2QzV5k
rebNeYi2zQ3f3DGlExkks/x7a4oirSIsYlW4f1qVVAHLTZv1C3q1U7KHU6IOrewJ
1fTubJRvkP4n7qvBDHAAMpaUfJiN90R0UZXoJMzuVMDriL91KqcWFITRCE++ae/l
T6NjVrfTqfdGdEwGgkIgarJwtHYN/dRtgZSL1gcAdHYI89RBoRomiA7UixwJuIxa
TfjbcZCZg4cgu7WcOsX30A+ZvRVOxtPzM4qDNbtTiGfi+zHhdKycmFpnJ5+q/o1g
Q5a2D4urW2MGVGVPHPimMippeB7IwoIvA0LDZz+9T34dyEZEp1mBH857XTllW+1Q
B6baeiWEysFFugX5lgVfRiIjnBKjfmzlSLPkqhUCrEnbfwMV2lnfjYbsfpCp2M6F
mEJR3mRKyCkn1mm1Yx0oIuUzsh68+iOy3QhGqjTQYV22Mub8nnByhRDRhYdlcTU6
YzWmv4+c56AxfFHW9MR4kzXHidY2fuvvioXDao0JboKF4vG3wQDTRjWVyg3aNEvq
86kOsmxEgfmkZs891YDN/UHYmuz1jL76M0uJ1iy396BsSX4uJaq7QVFw1wuHdoy6
kbqNUmc0MArfAVVYix/dUSpTrxjpb6ZoFOSpAVN5GSdhENn2Y0VKp3cxwq6RX7L5
VdhRBfMYyMD/mYkuWCCQYjU02uN0gAf+4woHlpQosAl8RZyBqUAQxXKiBdsX+ObJ
pb0rogBSuKJUc3zHD0tCBg/tq3TvgTl+QJUsCzUTp9zT0n9vLa1VO20tsKmHlOtj
sofne4vhuocAv526tvLV4XhcF+aiiYWKJaAyPZfHJGBlzZqKMnQXxcpNptQLr6/C
4ARDB3Ad0hkqckUBSRty+RJiXWjV0qs+510MJ3zUiKwQMiG5P76Lkv13Ml672suT
72+wOb+ApA5HenfdUfgk5Gp/1AR6RBrU08k2lbS6WYBGwAEXcKDdqsefvgh+VhoT
us4RzDlrtsYj/llFOUMkcB1KLA1OdeWLC2hIu8l53tE59cDXMiIc7L02AJSakxtg
tV2u7n7rb2CNdDMiqZQ4AjzksEa5O9MvlzND/acPoeFz1LzmmsBp4G/VTiyrrUXd
V0Iys/ROOtlKs55IAjp/wn0pJbb7jmFYsEH81002Kw/z922ZOTSCeHomhVzQPvc8
5SsTiZuTruwHGsPSgiAw7JY1AVThR167BFdtOAnzSPDbEclo4IXGfuVIAZa2dE5l
kJy9Swp7/Ed4nWP2PPiQNbJ5c2yFjo4xEuTUDcMA6JJ7W5tQIprlaWCttj7ns2Y0
TvX/VnzwLBhiPDQDA8peX+ooEEtrmLOT8QHaU2zXaL2A5K6L27OxXVL4wBbHnEVj
ajUSzdvy9qAi5KauWIdY4u/KlwGC4R8BqaPm+VATyqx5muTG4p4mrHDOYRxX3K3w
pGjeC1pJju7D7hgeghTPouRFwmFh9wiNRAg0IEhuwj62R9CXDtO3aPy2D86ZGGoT
qWO3eWBs+UDXteLwuAlCeuVWVwpQUeai0aR+BQP9ML6y61H/xiwn3ShtG6toCPxO
HhRNcw6TaBTuxDgRJraM+QSYhyPaE5rKHDVVbwS0i7g7GCTEO9RIHNVc/G5rEzX3
ounSpyC0cDaoP9VPguGJmhe0TBTg2KJmJ+MCiqk4QKTiznvKG9tFX6YJs6t65S2l
1A75tCgYDZ5hkDw2Keaqwpx0BoOOq8FbrNxCWnvl86o7u7DEMrpajS8id3nPG/hk
FHSVpymPJ0lmFtxwSH+EYWH1t5msI4tLOa7PpnQo5gzw3tP8JWgTyVKACyb8LFac
l+iD+e1It6O2VPeyNyCgUj6Ca7oXgJFv4twYN5PZra2zL3tG+0awUykO/sT/xsaJ
qmWqczAZpwl55QwWwGmtq5+GNeWLpXFhCbWpQbLUYGsWph9fC4HvQnndSdzO9ZH5
5CdpFslYw/GVM7AOx8GJ+wM+0vqgX5E/bHklccB050Y1UsPDirLry3YDj6j4yBYd
iI4zskg0M433KPAelwZtSGKzzpFDgKRmI3v187wI/BkGqCDB91GgDXUGl91nVXUR
VbOSwZaoUPyQrQ7BUR8HjRKHunCbF87bwa4xhtjxYCDQ8UR6wKKgnTgrVgBTuurl
BaiSAD/53BWfRUDh4l63KZxUwovEPFcHYEqGrPXRAmc7/mLnJ9Nx81pOGYo4PIb3
vHscD1nU48wL91Vdsf0IQASxSwzl4cbVfenZ7OruENsDnQtoLimVhcWFhh3CSGVU
LbJ2mM0Qbjz5nSVPmlWEYxyevoKe1IqdpmVuMgiNK+fIdXCQwNk5k7EKWDebGaxI
zBBr+Yhbnwi1kpkK8xUXah4xYfbeIFS+eh4qenNiugsR9eeeQFn2demNLrsYqn2v
ucqzLtEE58uGh6AS+joO7HrK+TxTx7TzkLcNzSmWNS7sxVgf+FaYyU2FahAOY5Oe
SS7YnT+4FY/2/bOKJ5B6mBrpHF8NcLJW3JxW4Wi0PEISJ/jhNFUj3lzatMcymGxc
tRl7HwQZsygDcdRUfxI1Xm42WJGUg4CC/iOju8k8E8Ceot4xvAH4N3zPQGLj16y+
AaTF5q1O4D2XPqwlMwg5bxt+dRkT7itx0Qordmf/kpnlG1F4jImIxQ/asVssnibM
ouaGbBXUDY6Ck3Zsax3ojSryoGzY/6xrO+0HGfhGRrKBfSfpX0dH1XWeX7eoOokv
NO2lpHh3QGW7GCu4o9B2ySDq2oIM+XqwdUzPyAoIMVdTmH3i+6ido9MMD3EpqyB3
lf/O5n7ZUL6flXjt65rJhSiWj3sBJUHY4gWs7u3DNZPFYTHQ/+m3IIxHsewwLzzy
dinzNmOczNAzGUx/J6ri8JfhSwIhaliZ5L2zTU7V/m5ayfZ9sSOUzNYmnRloDXxY
5ODr20TKS/RFDwsYDOPWas9LTouwZALSohXvuYtmbKDGUs7mlHjNI/GW3i1b7s4B
4zryzPCDYlDNo7Ncepm5M1/jUGMYxoj+oUNPrrrk47ZmhFAWla57RycU8U684sFo
H1+aRKV9w2Ejw8fJbEOXZ5kuB0Tzhz6w7DZPLR+ES9zPd2puaeYQfvtDbKrJvnKg
MdNM1aPPXi7LiM/h9HeH/l2oqystVMDwN/UKIImtGyXyBTBJOida1ioabxjhN7kp
n6bUhw1Pxx4Xc0YkulTvtxF3/y2aiUKY/8bMKpWJ22R4P2v/dai3VK8fXVCcl8P+
3ALa+vgQQDqYZz9Ey89du+UxX50zR8q6fVFV7AUCnPcZXDt+b8VMsnjTgbresgtT
6H0JMI9lm8q4OIwVdjMyPbznKH6FfyMhGso9tSGwZeKmChaL++Wa3djCrdq1RHHQ
k8EZ1jL9bjx58StuPMui85ZO9ytl9TVcGWLAW3wRT2gh7gmNz+sNS6jItd0Oqka6
XfCh1g0AN3RqUc8VLlZO0xRsqXNDbn2eZ+Q6dKgZy0b8OMeMOQzH1cgNoHMHzxUJ
JKdJJO08S+XQthQqkCmG1afKsOTc0jC/X4OD8V0PZBbSHXC8+PNpwdJpUQnGjicA
FhNlr0ZLCFIVQvZiEjHQD0wWsLAwSYdOCC/16ZvLTUgv5Ya85v0EgGVsLV+TKfW0
kWOiO1V+6ayMwRv3Preye4XMZOkEf/p32Cv3we2PpurzOOK67xEe4O3AdsgFbKdA
b8oARglNc/DzHo9514KcjbVVgNwwkAuZEc1nqG4LOHDcqczYGbwtMvPamCj+T9Wc
eSXfYCZD9exexdN7+RwJ++xyJgQVfODMsCvFSfs6r+tDhZDFivoPONyAv6bLOtCv
ko4wsyhfLQJuxGbLa4ZU2sq8u9rz6EhjwTmtohMynvu9OVyxXkerl/xz2g4NjIVl
K6khNN3AFo8RR9Pu2GLm70OTX6ikX03I0vZM09ZcG1DJhJ68oyYwxewGweoRwf4w
6Fe5qI/MRjn/2n78OE3FVj9ZdlL6K500GuA/CCG1E3zNcCaqqw9reXZRXh2hEnx1
2SoWHtQl/Kd/b/vBoWwcGitO/adZHY8jr6qfuXx7y/+0A1Ia3y1Rgb+3J/OAWlT3
L8F/8EXW53ylWmrhfzyGlh0dR/FvMJtYRZpLtmdCTLzmWXVNTN3nNsan7VnkDlSA
M7MjRBJv9/fTmMJFwLa/ynOgsd8SqI7hWkVpMrnXirZeSApkfSPlT6hePPhXQdpZ
zLxlg8NoQGwE1YRfULSsWNkwJh6OV1L1m17Ct7QGQdcCgcnRUA+XAhRJRckrRDhd
Gm+KPlzmDFL//ljBzErmJ+5xzOGYHQYBOcYGgfEJx4xPhqVO09YZlmynGRb/fHXb
7Z9YREV68z1DVUkf51zfnWv4WPjC+RPSPoES2PXuWUSmWCE+9oNlxkr/aEgynaq6
V1I+WtlHDLLQA0SOCPpkXzKuwxuKzprxVlYgZ4r/vUTL8/vrh4JnpbshcfgCfIEo
cKvpwrRsBh14Q9NQ44U+e1kyEMubKk7rh8YPXiQNUFreXQIXro6mFvg7eArIb0TQ
SeN7Z7eoWMd6czkSR882eZSFd5kgvY+sbVmcTnXt+a94mrU/1yQ/2EbF4fQrxM5B
7p8DD5jbtjhja0pU1kRPQXhV8udFj9iDBqaIc8wuIpRGluLArQvcYVLlirEd3OXL
L3xrlJb6U+e1xrJAs4rXu3Wr1sc3XVoLmNX18k0sKn2YDWxufxuVDX1YTtjjus58
kXLC0RaAqvzWQbbV8v+ypn2WXmZ91XpVSoshSpzdzixRa6SrA8ZR+EVqz0vOxyDk
1nhYIxSKbBXWpmh2pSzPYFyT3tX6WBDrnlqwFfHDIgx7m7LDQVPZEa3JZkI50Zd7
8W2MVQU6GpbtCEyWt5jdQ9hQ75llA/3jmn/xCBWE9eXGpbgoRSaj4aUoV+Ijoecd
qR6YTxA2yU2plL8A4V9pnJCW2JrJOwxZBge53oOz38cBrrIzLBWH1tC5J9i2yQIx
kN5VlmGhF89pgGH3LNKvdeiSE2E00x+D0NKJkFS2t7cJ6UvxbLhlxd6E389HYz53
4oKt8IVWGiph15Y3FWQBV1BO75Qv6kKPGQeZn3GsqjPDsWEA8+MiSu3RR5LSGw+I
TYCRSOPFB5ayQBLcJl5BasRzlIXjVgxnmrSD/M8PnlG67ZfZ/NISqX4WTHvzNHst
gOketKYY95v/hqhGQ3JQK5Rsezvs7wIcc1QU2RXblvR5AeVKSS/yRM1kRHIF4fNE
fNzeo5P8F76EWJM9Hd1cNrWii7ynerCZib9zqXsW2AKkM2NzvX+s79aaHtT675I6
x7THvoomfRRwkOZYfZETpoHzhWZeuYrsR4MddbsKVGNw/n/mXMaXU5OAsWMvqCfz
AHjTJU3uLQhmyNsddLYDL79gdCce7BH+qWwzmfQOV9+FEEBYc1ORDL6j69dHJFBY
NmNfmwhOVBYF2x4X2s2IU5zbcvE7LK+0O+FMjJe+vep5t2l2L5b9Q55avdFcoeRr
z9PcbHzUGQ0AmH9SphHXr3GFYheLk8W4ug5Ve9p3E9qiIXky+KW6J6Hu7N0123fh
CPnEzLehHG3lHSHo8/DhOC35jhow32pnDNdAHJZApKQ/2XN4Yu7q8DLht2pqkeEJ
P/pOMyhxUvvxcL9qNP4c2cDHEzr91vz30iAQYbOS6RBIwu/9nCM+fRFuejd6Wpup
Ca5PKFTK1E6VEwgUXaIxzqAvQKPRzGWlremnlVnQJu8RnztdjoWsh11YkkkYe5OA
PAmUgiGXMUL4faJTkRp5T4XEKpuQdmS8/4FpFwufKvt10xSxiZWsYVzJf9GuS2Nl
hN9I9Oa9zb0xtI0c7Cfu6jrU6REbAO57Km6R9Zh7kwEjhrqYwtjjA2Q4b6uVA5ub
fQshEY6cDEPB+SOtrngWb0Iel+nbInH1yqBrKVg51GJavu53izPnoVhDAizF1loK
lfB3FIo51kJJ+JJxYkctpv4ygz/IShSecZgN6GdiuSPuMQ1T2t00QlWT1EAdQyuW
cZQcS5kQ269cHqGfpYJFkShv9LwGW1V2Rk3KRjLCqhPExR8vEwqopCcDLCIwx2JG
jceKXYvI9l7HBJ+jkFpsm3k9umZaveALE/r9sSBXyg49kZnetwHx4Bk6oP60E+++
mwNK9QUB9MtC+z3oRK/+H+oUCDcPCtTeu0hsgTDfNXkg28xyHtPAgw0DasyEzYMu
zqCHoOqKbN4RufHJLrI3u5eCTOOtEKiJeRogvMM6JhlJ/THwrbbb1PWJys40MhWZ
Xe2dq69BFttHVxQXQjsBUwO0/KT56l/afXc6wSz93XsA1lhmSkxjDGyouEQKeDLW
lAGqCgZqgSnUnD7cpt0Zxh6V7b0QJEkV6GTJ+BNEoESY8MACcEeLEOyUpO1a9nys
RGB5QbK1k7id1ZoXKpzpiNuXcLltpl+cqdp029h/3xbXdsKH4qZWxwVBlvbUCcP1
J0t/PFdHx6TkYjO0oNcxVkfHc+35gZXsBgVXOK3r+5SR4Ss9S7URkF0eMLD2/q8N
Qm1soccHfjz0af08FTkP8jwpE/1Hd9W3z8OgempWTE74gX9dUt6nIgmkrr+33qga
WE0EUF+EY8EvZMpuX7ssK/9QP9ioqpSrze5IARzgsdTI6B3RWWiuSSSpvqmo3x2M
iNAUbrMLcfvIl4k94DtcCJlGMnnE+sHYVKBnPNuB32INgS4ovagSuocTuMtsAHuf
jcmSg3E0lNBV1OIVMl/d8V2FRBtfmTkqat1jRA3yZqG3Ip5WwH03dg2ekjmjRbqI
1mjB+Cs5WfitP+cOvbLmgf6u0Fj8aE64rAT6rO2F+H3z5I3J8Gud/fBi0W9ktOuw
oGJyoHAjrR8e/XZ6Ai0lq1PKuhaU2Ux71B9MPsmfSr6znrUpCXxT86s/ZLP88uMr
qaghEx57pjC9PTioatp/Jeg0XNXoY6mKvLB5P2MJ/ag0oGDzIqRKtz5j4T7ZPR1Y
XjhnVURAljoMIlmrtyDgGNUZvbYBWMLJEP7nmzV75Gcv443a3Ew3cSJNPPFpJtOX
3yQUMazucaWpLtLDOyCGp7qAH7HY3krITKXIIL4bNO/Irs9kOSEIgY53J4TQK8u4
QxIaday1/mmdFbhMJt+sP+vvglHX8FDJy9LGXOrG7mnBfQUp2QwBYXoyNDmhNN7Y
MShJ6lzFQ3ODSRNtNIgxPXOIMbyMgBUo7PVsJ5WE864oFPSyNjUeeGnjuzARnJ5G
P9qb2CK3nKxJypX2sdFhu+uAa7+pFI3BqBFZN1B7J/q+9Evdyst4kIHS21F9+FBY
MLHY7dSkiemTcUGuHNDsjIyD3Dc9BC/8V/rTSdOUNjqC0yI+Zwm6go134Zz4fzPL
Yb0Vh6UUC2CzcPJYkAK5Z4EiH2D/LeJlL8t0pzMXT7w4tNX+S/0z43segHFRdl+C
ZSh8Htt1LmDKRKYGNt2Nl9VESRYXMHBX7pMTPPR8Izjs4PqqWJebqNo4NP5Vjd2I
ifC/a6g0U+Yqh/c7pym+kZojYGr6FG1wmLVuMXD0DKfEyDoD7A51gbJ7Xl5nmvnK
823zyuABbyKj1ONkApC0olcn+sifgFcH0JhlTxIs+iuH24fwPr7ZpYYJllBpELt7
JZR/ZGeCG5c2GfvQ/H4sD/+aYE4F5Qaxa5cIjnHkP8OVVjHNWRGV20q0S07/KjPG
A5GszyEjbEsdpx413e/1UEVVypAHfsjY3ubujNfqB7fAVEYSOXD6RnLYprbozyvV
0cXsEdgdS2dLR4y1vKXLyvM/lTCmfL8/xbe5KyKLA04o5K2x641Y8Om0mchOAcLv
r0THs35/sNcy1jE+M6xpSb+5gnp9mwy+4zOfKf6C8rj5BOBx/Qd1++EIgfhMC7Z0
Rzjr6esyTviE1SlKBqPpjErqJPIMoIWmHsotW8egT6pmp/TS2NBsnR2pwxUEJe6/
I01SVmIAT1cvZw5W6LZJdvFuwRujo5FpxQUSgdspkFivRrwCBzSbxN7DC6FSLgd3
8pmcEKuvY0jHtgAvULQuxOQ7lSaNqnTD9YAOh6bX+AFvXGlrX96QMNB0kUolsKBT
r+IuOTnl7fgDVQnzs93rnDpOYH+OJbGXSQhvFiCy2ary8e4rZmX2KQyjNIwx9BD5
G1p+jI+Yqb/OrZqPnIvzo3Y22Vj/tNXqKER35UC5Nz8wk4r6Xm53QIDxCWDTEIxa
GdsrZsf4qmw+hv0ay98GlbLI7Wiwokz+v/0zARKGbsZ8JmSOLSJnlYufeOMF6N50
kyew5LclEzrXrH+WFMwwPtB+xy5fTECIX0Umedhn/b9qZWjty9Xl/dW6irgoi3q1
wo+HM3/bO4vRlqp/nvI+wlv/M6wXIZK4UcP3zlAsWouCiwMSTqlQsbkPTx1XKEUh
JZmOn26V8eJFotH9YxpRfezYf02V5P4GUiYHdwLLTtiMLXjrptkTPHDDaeO6HmVZ
Ls0atgcE3SzsnWQO0jE7FvSdrSD80V8gmNNtdXTrf+hVIIJzBI7/8k2EaVqZ2cEu
qDMV/JXIRlSc8HfCXpmxeQm+LJJaBpmjh9f66ajxfEmMDYEzroKrFBD2SGqx6Yy6
glbTpTyrDznNm80Z16o2gVxCHVBBnUA8lHO/daU1ViemZnfZFUrEd1SEysZ8WMlh
eGjYrGHEJLYM755ipWEFCE0h4TNa4bS/JRs1gOpINrjLeoo2I+fqF+HBarmSUDi/
01ebB6+xVz8wU4QzyopDSs+17mGQcKrAkBVSLPFaTfq3lrHvuuAJGkI5v36S28mX
3zK/Jfu0WqKvnJGlh6XR0upHlOv/uXfBha/gRAYuMFZ9BG0MRnRIn/jibhzFY+Gm
aSnMPOWesNI18F5tK8sfMseIabXjIs2n3DAxyWWPbhbNNeNwXGEeWT/h20uDi47c
Vi8Vq2Xek57d876N7M3gZlyQdj8G/mhn+JQ2FOnyhZeBDu1ekKsImRSUzH6nb668
iFdxIc3PaFKmaZCdgT1mHt8trISP37dfZu16SrvR7R4VeANTBQLJaHTFrN8e0N6H
pxDJJvjO+N1RQzbNZZ/ddaewDrLuqaeET9n8Qe4dbq2MaNsOyeQRpDvNLGHNsYz0
7aVMA7yOoDAZkveqnP3OQAaSDXlY8BRagHnVYVmPWI0poRwSUwdk8gAjGiz1xAAS
V2IkVkyvp3bib72NJMxLzsLb98o/y4omfW2xLgRRMKRppVUuOnZLnl6RusKSMMUL
jlB98DX0MGpgzDHmvK2iN10x2dSCoM+OhUYHHuhAOeAVzVjm8tESDGxG5eeGcuRA
Z+pUyN4FVHAm7fbsvtvR4Ur7jwGaIOdZeOx9G1+Fkoq4NxcpMROQPk5hK23wGIp8
tpW+kJ9NBaj0vlGnhYVkoJAKXrIqByvqSiJtS6UcUAtaS5ZsDETq2NAaP2yZltO+
l5lCdqd2UmwLoPX/ddFOjk+sB627eVIGv/uw4m+UOZL5oTS1Zw07cuMMz1yrfK38
1nhsSba5DmimoFPwiZ4GpGvInEJc/0PGpsfYRdRFoLtmFmCMZemJ6IWK/zFtgzZB
NPS+KUfI2ZG2Y/tUAog/VZe5SMnHl6+LXrL+OQYm5hjmjcA4lpZVFuSuIM31Iwmo
va1topwQGSNxPrUb3LzHxq1rFvUWVNbsckYIqU6dZRGOsBlgdPx5sCAOSudwUEUA
RsWJioOAvZgk2xokRBSqNBmTJyBKW5EQd/8Ks21JXeC7DORCMQPh7I64vGxvhidi
mKZqCk5kmnC+9pmk77XUsuD1yq7eZy7iQWSY9n8Xyy2hIPh9O34kHHMbWpCAZfL0
2/eGy2zYuQMDsLyPUlmNthwgTz4yRQzLMRa8d3MdFtnIueZsOJbeWJKfHV02Yf82
pPBb2KIoeel8swYh+EAjO1Pb0T4fB0+FigHDpSIZ/nakkiRNRfKKWOjjYrNqAfoG
5iaIbfrC/z8hxj4seCNvQnAMfgv2SJPSYcg5PNFbSNo4uWm5zL9blhTE3ug3CI5E
j/F150AL7Drqj2gUaE7ZYdipri5krhM7+xvLvWuDZi5xLbk2PoRZnUrrxpbTg3Tr
Wr/DL52UR2VOis4Qy93s6uYzq4DwVh8Jti6i9LZHCnl0HvxwOhMxUySwgCg6ac2L
aSnA45zJtq9QjeuwsuoedE15zXLZGWS4KO4KZn2ojMBYx3ZBQIdKZ/FJOp13Lj4p
nXQX/w9m01PBxwQs5dmKaSEcoT+0YE3T2oiMqPcC2DhwDernAlZqh9ZwahBmOZC3
jt3s/qFAGMKWqCBiLrXFFY/7Nb5d67vJuB+GNogfZwFFuaOvAm/tWBO3XzwAkh7Q
B4nkoYMMgP8tjm2qiv0LeVWw63swkoV6elHX2bg8UgAPf0+bYtXwrfcNVbgGiP0F
X18YSitOyeMacox4EnYgJLMKjm1h1LssVnr5o4k9MnNmBkLrjpxO7yjdGJ9mcbpY
oLfRFKJjicTY/WdAntNHNMQht+aX/dR75RjpeNRH0EPAdoFAtfYtwXEZtIYnJHjs
4Z+Ip3XU/5z6UbrCuYlRVty4e3IS7idlIKSL/RLnFdRHH/hVmhtnYujn1z61sx9n
Ykkx/vzdWByY7Mu/pVVlACVfLg4RAxIS3RCjkWi4JoRnEUD5hP9qwL41q8+M5Bxj
gc30OWtsuuX3jCKUTsNbC71Bc4kZWxBrdIXF8oRY/ChVzGkVbpLOxjqmQEibGknK
Yvvkb291IEfb1smYVB72VoCQgE5H7zJszwYRBx5RhxzN4cwOx8UcCozEYDIGuRca
rg9h2cwIuPv8p9k+HkG4X5GhLjZI++ejAKI1o64AM78sJ5di5U4y6ikHsAX0rhcM
bkR1lHz6I2Q5YbU4/GlJ5SRp0c3WLG2CiLk4JxXCqEpexkSMYN6GVyV8K4exJEec
bfAeZoen9pjGujkwh0f/Emv5s8IAcrr7SHMR8fOGrPsjXzMDZ/0HSl9z5r9fRlzF
8jZBnNzTrO5+T629cOgDHqbnEnYMgYx+YifEcehIOLqFBPpUes5OB8XykCH/KwvE
ZAAuJXbWlVOq4yzvqyE6PX9Ukus/jgneHMsThkwjvrDgSxRWafd2SBiVsTihac9C
kGCkqaJNAnmJG2bXzO04WKFA5PGBBoSc5r7H0MSNmHbo/CvLiYzozaYPtk8Jox5C
0Xf+6lUYIBMbsz+PKost7I3yqxKw1HERTQA2M61k8Bz7D1XRWFQqz+XK4drm2CRU
XE/d3oKxfNwkjCKpB7CE6sFXpHVs7JShUreK0LO85UYAI7nNlfm1jRdIBiPX/7Q2
7ZBoSKrm2nx/8owO/vGs/HZ6OP3mX7kor9X88PXSK3O+WxL8iBAWvhD/+XvCSO8F
uLYEt+Y2GBlv3vSca7vBgRBYeNlSuHjWp3dwkDPsbePr5alQ74ktSCKQzIqEiiBm
OKKdIyRAG+uhN3/pJ1UFt+f31B4st7LMTGn4t/jruEZ2fXB3v/WyOO6BvVBb/rK5
vuUL5z2IbIlWnrQ+2hcL43dKiCclqv8RipGYQZo/pyzPN13XuV2xmcVpJ3t7xbxi
EZgS5ZOTQjkL6d5Dr+ZcdlzXrjlAWA3/fe5FXuOdCXG1ZyCIhwKhwJGCpoZfJY0k
VKBP0TU1dmENfPuD8RaRG4X2o797WpHzKUU+lReMZhMhNs9cotk4r3sGLjoEmPGS
RQi3yctGdVzXHoVd8jCznighoau7c3UL/j0AMDH1IbhRGHBvwj8TGj4V9QY3l494
IH6DomdMhhKu3CpY2i+TubrUXzgUwnCAgYTK6dmipjjH9z+fba7kDqhnmXMpBuDg
y8fFIDXpDQE1aHPEjZ58K2DCaAxJ/yals8S7KaPXmSZvtqSuR0Ahq0DjWv6VWHsF
bFE7jFvVw/xXt441w+ATkBwMutaMQrjhA43oPBdprK+fMGY7rGwXiiVk+OOdn5X/
nKsChnltTDwNvP5oJRUCN66aXtnTSxS761BNbaIQmaZXjmEa6h6zulUAhsh5IiEO
W5GadzcPRahBJZV18MLTyq8+SHGXqMVKWp1qOXDiayahMupC6x27jEp2iYLDqNJI
wpzydgTL5Ti/V44UOGDgUjDPNVOWbfBEsRaxIT41kohuwANyZzMvgA65kUzSFpwS
iHmH3rvy1BH5aN0fM54IsaMD0X6GRDUTFIq9h4F65YW7fFRbz6wFHwDv36Ny5YXG
ANEjvyUgHm9YysSJQ7kE35CxDBbwXyZrVtlHZc4K/EA+F2KdVTqIKd0Zxb+YG8DO
U/ProxsE/TIiCkClMWVl/eRq1CSZiu6+Zqr0P1wqIb5H1TNbOMreNaLJTZlIypc9
YjVPIy+283GFogk8V88rgjkoqeYp0IIyE75yfi2AfVHxS/DP2yyxQzny6E9J6vvq
Gmrz4t9zBZPYNF1kBcGesBDBpBwQf6alaHPYE3wASBWlSMEoz1R8Nfa9O67X+Wyv
tELiisobr8TVtjbJVny3nb1XApKFtvzMc/v1UjqgQX01Aa84MHWbGCRGGh5X1u0m
zYQ0UCFUMG+CKnExdzZSBNLmRJ3HfPYnoKOERlWVv72ghCF4QdVZalEmCm+7JmPj
UBkYVypkCpOuXyLJ0EpBZq8qhu4GwLhSqZBH6j9oYfHZkmQI5NE5jvadP99VRCcl
yFsXuw6UXPpoTUwRmvB8Hu1ta+1qclboNemDhoXTHLAbh0GrjivsHFVmJjnNiCZM
OjRSYZxS0pPTdrK6b9wQRFa6Fz5GBymmEiWAHqsB9y8IDxxMASvNbMDmLbDGIkuq
e8xWEcYjwz/VI9IqRqqdjxk+qHtb85jvevGGMU52T1ioayrTiaaXLhWkFPhfZpO5
4xa9+B2j1r5Qkjs4Mv+O//wpbQI58xoNXcRW02WQ8+AXwJwsv9b+QvSizd7L2WE5
bg1GXauDjXpb9LlyMgyBipw1BaSMEL0OSYpu50sKBTKtawZbY2KTfJcSTLLBjH2r
gW9rqvg/C4hUNLUHfI9rSvdy855uxZP2Q4RT6R9JeJ4AOQ5Fza6Qjw4D0BStEh13
z0ElikZSaEqLV2PLlu3TIgFVm6AwdXlutaAtCRN4AQjchjE/35xcV19WRVaOKauU
S/ddIJZgt5gh8Y8CeI3Q51f+P4JjYQJh3NKGR3oRSHXi+yv/Qa1O/aK7ttpwodEH
fdnBtCiFXJbUB0pewu+RVvm/XQsExmpftOwcAc4PubdiHoQtD6eRdHcwtEnAGr75
WoVCCj3nsycQwQ44Jv5UpW5iSUGlwk0Rhj2LdnIwGNHaIj6Yl35VpxYT+gC3ZA21
R+No6lWMW/nFcPcESiyHoxVfLrH+r50WR9RgFyZBmuwrxAAaJZIRNdDats0IpfKG
yP6/QboQOMq0lRVXr65vXPL8RBgRHGmjUp8d3C4x1C3TJdk63/6dBZogLU40ajKI
akQg1+58QT/U7Pken7qilroRSzHMWBuVFjdZxs/xJBbc5o12B+AkheiRz5jkTc+I
dUXf/E0v5GXY03TrfBRpFVm/Nf3GyPyB3zIS/5RWP/2NuDzkqvM38i2Dusg0DVxJ
X+GHR5FToG3/JfMtcFG+AfCZrHZvbe/YBH4cBzMxWtjEI/wzBT+z+9DfrXN3q9ti
+KDTmtxaU79OSzOAvBNwUUTPPep0jZU4fsKOTL/cjE4XzLYfNXbmzsfaYiWnE0om
VNiMdZzJ3tr/SeWSLZNuag6OzcF4e4cR5cZh99KvgAWyBxk5200/xcUTqoWg0OhM
fKhB3+zsNLzqpOs2Vznsv0XwK2NPflKoY6tfkK4F70Wgfc8Oqqv/Rlfb2CGElHlD
Xwm5MtUeohJn0OmR2vIYoCv8q1LnI5qgk9O4Dac2YdQKgn3o68eFnriha6DXQYg6
6bfEWSm0MNwI18k35my1+13Ju5jJfGlwlQmknXMGKXrg5VyDfHqywA+1lknImXK4
R6OYYf3n6j4ChnRQNAqmexhGVoKX5nG/svzA1F3rEHqeO+JhZahf+aXCNy1Xptab
k2Nn2L4mnbK07bk3XqpISDBaVBr4839f/hKQ1HGbwQqdoy/rdEajzyE8BT1Mgcyi
CsOE6UWuP89yvvgagDHNu1eWV0XVO8RQvce+WOoCNAUfnozx2JUf+uv9VN8G1Fci
e8Esvpp+DEKnq+RsXHiTZ7ENaetdFAP3VvA8+wkhegWOSWd4K7a91UB1o+gh1ojL
bIZVD5hvCETA+CxA78uPBduRYlecatYLwqTsl7Y4EZ7mhAmhlFxA5UmzFILJrtNX
z54ef7YotJc6JI+g23K173kOM6GnazjV5m/fYFf5RDj7DAHyscIxujVRzYcU8b2G
ur5WE/J6h5MwjL/d2RlYn5Avs3xpm1wBxlsUB1zxLjWTCFgEMRtxYgnh8kiHz84U
hKhSveCkVEvtT7VmBOfLeHylg5K55+GVnNOW2hiY+zYfopV26GfF7qf7Xc/b/Uai
9a2wrdvHyPDBx6k4JvsUicBLu5nDH5s1590RQNY/jKCsQjy8eAAsVziAlAUa0Vla
ct/VJbKfOdb7x7ox/WwP/ROyelXm3EbUlVaqbiQsjkdQPEeQyRPbF9i0YXSWFD4u
0msf3Heb0d1ulQpZb+wsDleQqkFj4XUbehRJP4gBjZiCAvDrKqSPLNtdsl9x326s
JPgR47+TkCIHcRVbU9zzpM61+PQzu1QUOZ3Jg6c6S+675eDl82SzwP6lXW67rz8V
sfzGN1Wp+PESfjUFjGz8w44ZqALBUtKR70m8ismmYApYDcp+dFVgoC0babrKBoom
Tw9w/gbnaRRsdN9FkKRaIH5XJ4G9u4m1Vu8gzFQ8R8Gj8lJoJQ4EfJFhLA0upSuS
AoaE/1F/tg6JoGfrzSs45k3oivoOdATlp4+pTmhOogGxseC1lGsmQzNHtdI3wVoI
f/5WXHdKFq+fugcQiauw/ZJJ5Sl4TtVUlf5P5J3tCZuE+24bZXJcBuV8he/ywxKb
oEVkG4mNmIL6yssQ1Z+n2pWrfQG0igrZolJU+h1pJbubFDZ6YMpznsI4MHFtE1OT
0GZGM9LinE2KVhxZyf6epzvZvPzbDDNkiKHq05GbtVOL8uwCKYFOD8Vvhq6U7J4H
pzdEq4Ms28NeKj5OXqHcpg8+5pR46VYV2WTaoi2xj+CoOzBf7bfFIXGRjZl16d/0
Ri9FVrO/SC1+QgctjD+vbQzzfVKegHdLpwuw9eFMhJbwyZYre4pukntWgyHzoDIT
haerRTHkRpTObC0ZHQEHRbkTuxy3wQZJVZkmVhUKxT13bRsJO1PuH3cZj+wp7Jbp
A6w6JT2ZYWMsdv40Q0Jx2Xc2ZjR5Pa1ritwIoQOyQl9kaBDz3RqtheLzGwvVCp0m
9lJeNqR8su5OIRW5QdZC+tgedAK/7VxU1cv3E8714S4PhDgC19ee6/hapLNM0cXx
Wdkpp3nYvM5T6jQTyx3QKO5yz2FAbjh+uvnKznJPrYOIMWtA9BY3yB5KyHzrMhQg
yzC4q3qLv7fI1fmjFiebc7z/Svot2Xi9Zybeqj2YJgqro6ea96kq5TghJZoHzGZC
+TFsp/IcM3jmlLDs2UU46Vk9SXLBPMHKGVcVKvEpOhoC74vE956jPG89U3f1LD2K
bzK8lmi+kCSxx9n94j2TjDpQxtnvTG9hCbwbUsiVEQ7H6bUxPiN0xg+fpgNhoaEM
jaXUVAbHXwBdPFNiQ7Pe33rpAsag/ESZY7wgL+l5SEryLHuuv3ynt/GDzKC/C7Ot
JcUNCOtMRCBkxfAKq11lIUgU+y59g42PJ76BI9kNsGl+zpbiMzBsJNEzhVrg/8CF
KjG6IYOSb94RR2sExp8rkZJPZnDA4kiR9bz867LXG0/Ek5aDSSPVLXaJoWLMcfAR
jrhpmVcjVcSLgtdMMF/2GWo7GotkVhZMW41l7wouKIeMp0rei6IroR7UFzObDbNY
IxqyG3A4MsSzfM4TlozCpWDYu7+X34FMLEU1l5TMrDYKCc34XOCaRVqw1j0Rhq/R
DwC44UNwwFEogcu3sAmAc4Jabc9tBcdKi3CX8sfMRqp8iArAruRufEfOu35DVAul
2Afj4PHKVoXAb2wZlhVsxs5tehPb2yPA9vuCdWOdLh+qgcoW4pSpE+Ww1daBO0HR
VBda1aYXLr6BuyGP8xWSSkkOMx2txMNqW2dx8MST8rgofBoIuB+516wZiCw6y2JU
e8WF4cL7NNe4ICt2shPC7+3fe2bNmu/Ys3RVp3Y57l+T1wzyII7NI39y/sCrc/JH
WNOKqV1+hI9v7a6owf8eGGPc/Jutg4wym73vYKRKv32AHJtJkuBDDiYshXV+RByG
mmDrU1JENal/aDNxr3w8UV+IxTvCt80j4xfy6mWpFnzPZFabKsSTWW29vYOx4QLf
SelrHbTqe7fZrqrBnxLZ2liWyLgDRU6HrEZnO7KYfa2taSzSmaqEyOAQsquJVP6E
ZX3kO/8gCX5BsIOdQRmKYKWqaiFIPYQg1ARavOWumLJK2ilXK9Cph3wNn13Xo4bA
Omh3hCrMxdimqjw0uZQLkQVh3zsrb+lqtxaeb33hl8YaUUoiR6AvNd7SbRdKZaFg
vVeymSJOXQCibddygGto8Req6bV1S7AV0jul0p3fqRt5TNZPLrHTvMPaweHG7vyb
/dtalIB1tCJm4yHCtT1U9SZ6q/sm8TJK0xy4ENrkifxaUqQPZJBUjsUs3wtp0ZK+
vw0RyP3u1M/IsnJJj3NxjmRz/6XDSbMdd2GYIxiCvpSdKVjFewlihsgLX0aSdrhN
LaultMCFvwMDtvsLkrlm3mPrTFuQHcJTKlYLzPsI4vh/n2pzilikg8fmAecwdc9d
NwEaUd60U45//SnQRCgu8R4ckZ3yqjLswRLrSRDHYJvg8dwIn0VHLmVGitprih6R
p0T07EVR+hdyFO6LMmh6b8LwV9QklusDdWBb5b7hW4+fgcD+7+Y+/XwOMCJXW4cb
5nmamcptkQnra9k35fRdStAvMIjNSR0Zm0s8jcDBvKQGt+zdZvsLj0BPWSU7e6yF
gnR8GGc7TkIZAg+RddZQeFBwQUoR/GO4qPz40qNr2jLQa2Dm+Q5lO57kq8sXmEzo
ly0OBihE/+qwyEpzViDs2/VvPnPOa3Xz8ml0TWTeFlz4GeiDkecs/h/jQueGLWDB
CCSWuzB87IG5jYfvlu2iXuj1r+xM1hueoSFmFV3uWekhnKUvXmCc1N3GtJCgY6SF
XA5Q8xBsLN+cgGmjewPgk18PXw/hsrtaoJeje0CA+prkPVptkqu89/KPLQxoaMJE
bS0XxhsFqL+rTbbi6B4p2LNvwH9JvrE2aaX+/cf1QAhC10g7CSoU5dpMZ861WyMb
/DKwWCEQDxwyG33pdYgM2tlTF1tXqOaB7/QPjBSXCdRjriw3nu8Y3E7GKS5O7gBe
Hk6QmOuwsOla4wRWQgOHwrfpiWFF/K99Rlzi52obfavpmlDukpfMH/FMfdRTzekG
JSMk46m1zYd1ItBVwxdOjlNE0f5zkEWLrmSGa+OK4EUUd4crNl/hHEUwql3CSDDy
CtekELxKWgaJa/cuwubaLUFJdhETC/zw4j5EO2CAiHWPiB2V+EXZOoWbI0+bB8nw
8eP/U4DMSRplJMbwgmfuLy68fHPJR3854oMrYbFmYctWm8BX2DBV8s5VTw5vHnQy
F1h5IVTpkGtlegraIr3YyoZA5eaPemNLdS05Jgzig6Y0JUo4S2jDwRJzsnid9Ogj
Mo/MJa8S1KXWRCf6VMKvLoDuHpeiSTogFNHrN3Q/ka218ceIKGp+wK9SGMW2tRC1
jht60xS7o+Rvuzu8d+QzwdHVfpFsHeOJZb34+J2j5qQZXFo919Nl6abJfv7Pnv5M
2XLkqkTxsu89mMxoYhOm9DyitO3jNDIx+Odvj3jIAr+o32rcBySM/6sswVXwzMT8
cC/7QVMyCIcDUA+U25TJR2myZhGie83mmQvl8q6+AluxjGI6EUBkKD8eaN12E/gt
xRybSK1XwJ6oOsl2Ep+PLtzIiy5H7FTkOZ+8kx8uNC5H5WSSk86fk5fz5h5dkcvV
DyCMB5XDZZFEADXyifxXr1EU81aexXeI9b9kOgn6RrcYwfCBNnI+QvPRq2kCBDMg
S0idJhIb7yCjWt0DwhXdXGUY30kkJBDwGEEHGsbIXrp8wfPBp57Nrbuisj5eyFzl
Wxiq4Unpc9J93i297Tf6JqGcoQgn14xY6m9sk9+scPzcgt9QP7RtxVJmt3OTIqS0
MtAVNwEfoMYXqTo7H8qb9b6opMY0YryNKmdS8ukFhL/0amB+dT4mON+lDv+YTVBJ
n9lKGNe+uPQsSUW7l2beOGVlliH19JGqEl6Jr7mJSx58IvG8ak8UQ5LS9+Ep/+Nb
suNQsb4E3Hv0FWmAep326ZxX9HEn/JFjELb7h/4Ea38r6Xe37mPNxKGXcwwyzyKP
sgBa67lNp/g1Wqju9Imnxo6o4qOTNvhVJzS25Ga/zD9uRfUMP4w4hDD+tpQFupaq
vs0chAGZcfrUPKNJhBF2aEywVMzCsQCPfE9z0R6EGZnrVPD+x5T0ljJI8d4Hq3YS
bXvk8rOCIgjLb9Uzv4T3vQefBsVI0HjA7lvbj2ep1WR8Vet07njDRjTcIt1Hj8E9
8fuWSjeAAL92JhqT10xU2GctrQGdWkM9+cjc9KigcdpC81SRPPoxDDgy2NuDet8r
PeS3PN0sdOni0Dztns8dVNnBkI02zIrCoyvirDz9LoMQVydYL9c0n9o1NZYCgOKG
z65qtCnbIK4B5L2JQHeB9Cw8oO4L4oiaiGvFzcm2+AyFEIQRdIHFMg2D/uJErW2w
wDxssS2M+QI1ZkzN645Dx+O6jHISUy/4l6BL2nJEHJx0oIe9NvTPqHen0gwbwHwh
VCeA7K0gGH0E07f9czSQRchgzTNNXJSSLursGkuAjl5L4c6xoQkv2SdD4uw6SeiS
HKB6ZsKgzh9p7h6oD9You0OfBck28Ebp0saBKv2gXNvRTR+jr+dnwetnWezFeQk7
lIQcUzYhFUBeyObywdzQL72E0jBQ5Fx+rZJHiv3eecJSaIIXq/75ELBxJXNmJPqJ
sSCGm7nwfTuYM5Gp0ynH3bKtxRc+RoVmaOrKKoUfiHhjuHNgJsISZq5uYDZ25q0F
nou+BlxH3aC2ObkD0xxp7t+tYSMvCiXRr73uJrCSFTght4YGRDuXdxt7O4xT7ITa
uxAyqwB/C4wKA9lvZW3St8lNNBhTL78fLyrpJqxUXIjSlUn76O1CjDADmGN3vVQB
4NX5jvIC7DNyJ8PoDG5L8a0OgW49nt/lfUxhtPFOREnWko+o5QuGappNg3vU9tJ/
/a/hB1S7Z7IgRsrblP3rvROos5B6YJlg1rIqMVxmpf6zWYtDxcylZB2GXjfWsAwA
Py/+JdR7IBZSgSYNrm7vpatLF+VqyyzwZviJTuwh+1M8syU5kSHJ9wa5hq75UMfT
rE4yayEGFqbZ/OWwN2shkI7ha2NpH68Tt55jKQOqd4VO0qd/GDjdWf3VDdzF9684
3FVVte686cV9CNIOwE9U4DTbixEesgwhtC/QIJsca4Gt6lZ32bUHQQqoUQKl+r+1
MU+y/Bs/CJuoz+/I5dZkDG7kteyORmI8NP9i5D3Ul5EvGOydOS+DRpa5dkD3V5jj
iNe/qMbI6c9kRskrrTsOmD7HeFbEGZ9RVBbDUf+7OEuvXZj2Pu+PYK04FDEuT8JC
EEEfkNQguX0HHXye4hvVaHEjgbuDYxm1rWCTLcQDRyKHG+AIA3UCxMNw52zeFdqM
3DEeu25iGfxBp9cCnqh8QbtT+xCfBOUVzheyHdT9ae95WCFTGhCTqh+q84dfydUO
EOvzFiMoYvhuHYGTxRNcUAn2YE8db2v1mPK/Vd0rbKzS5/ipxJ7qY1xh60tzUBWY
e0OoS4dCGcRUsN2KIZD8ZaHYk/35EVL8V6dcpuou3O3d27ZrhIiX8x1SANfyzEOQ
qAI0OQph2w/DnPZZY6BSbXVBngHUBlDXpWBk0yaRZfckcfmgawuhrmUHcmmM9lBl
4fXscmK4QBEyGt+wch9SEu0L5CJtqzkODZIio91tkKpyF6hkiXYs/FH6ECj2Ogwy
mgeKasaTbbGDd4UXvpt/Ylq4HyLg/h3kTs2LaRAYnP5KSCBJUgwo7fpPzshVm0fN
VC/xR74utvnHFH7hwDwbxGqjPtKiHpU+lFJtMtTftE34ByLi6c0P9uKA8ApmwIlf
leJwWfaDOibqEQHocd2nkmGGEN5xbCduN4mpBd4/V+EElAZRJh+j/+nFHggh+Z72
j1B7C4Z1uxPQsHWdP4OXyxBEVfkuEEO1b3qkG4jGDNZWJr0Sp6Tuym4EINNpQAI4
OtzeB+3f7Wk57dQ5BdDLJyMZ3ipwr7BLgxZrQ+kS7+MgXgoJ5EusX8epa5XBkIin
phqlv6fm1GWUsEE+AzUwGNarnkofZZlxU5RXB4lcNJtZDVWRZe1ZA4yebBNwrAwZ
hb/fQKF+5z4HbRl2Gs71OtsZ54HrJPv8hDwQCQkfoodrzZuijgWJxoirZGQYzTwo
6gQPp862j0gHic8zkd/gk3J+q0jm+tfXkHt5wPv2u2ybL0Ur+faR3/lvbhsmgRPU
cNBKnB+rmyhW57Vqrf006FLWKJzVg80HdGLGjYfT4qb3KkcPK99rK1srbvDCxoOU
KYovJratUltBTFlCB0xcz19L5NoZ9w8ugyPQWC3NHyNuH8cndnXRkzqpXCR+BzfA
RMPT1rgHmord2G9FQmlvAm3o5oq2fpG5T/hITgHSiNMpb7lCvnIBSmzE2NW2WJwN
PlR/IYjchS08vl8pTMD6c4JlZe7EvxY+bjJsnlswJrSSjmIbgLpQeuRaaSLrCgLe
9bXu4OsQMn0YN4o3YXScFrZSZu1lLGYieUHc2FDSuuZ0ijR4ngGvIRywP/0H+x7P
Q68Q3ae7PiLYj3xGV31ZOcAyjPL3uiamwWGkfdJrFgi607jRj6T7WlXt8ZKmRk83
JBaIvQqGIMhVqx9r+bUH+p/rpeqbpzuGgkrBF5Nl569kHmqTDEy+njS6/hQxsU61
+1iNbCedZnQowy5S00tMbzCjKH+zCP5S7Rh185qYGHcXH6SfTjU8WWGHz1sHQNgu
Cmtq5Y8yGSrnyN28xshT5NdMFtvW4PPVGE19YqQXh8002DooVcPlMqhk9nGK5wJl
GuJZi1RyVAi7OvYQBINp1i3xZVLNCXzE6VDAhIhK0ApPumLUExyLlGtpZiHuO0Z/
+f6B6HkrbhZM/xmXnsmg/4IZUC6Zn1OtfTZG9YHs+Z4LBLxvfBKDJulbyU0iyLO6
8Rmpc40c7w0U8KSsjgec0CpaFJ6z8BpKyy7xnV+x9lAEgYNFJLbpSRj6gSoS7pYn
SaVH6adXcnQYpVcc6OuYYmIsqFZbqvmVUwV7+zx5eGMIqw3ZlUH8mhCIAFb+0z7I
AKROLG+6r/o2Uwexru6pmQYCgfT7GkG/UgCqIbk4mK4woybToIgGccLJpD1ZdERv
CeWin+Z1k+S4az+yo44swpI0gqK6myN0zLuN+VOhiNBS3GE6gp/3jgeF29CrnAe9
1TrtBK12wl51Os257h8hcJPnivE7LUwkAhmtoXOfCyzX8F/RvH8rrVIufNW8JnGq
mn5UJBBNuzsNSd4Q+LeMnNk0RvbQqz5Rv28/sgQdx1rikAjPgMG/i3S6N8xuMP5S
q44tilg91yPpmHeBy4J+7uoFD1D/g58VF/oThc2STLGRHherXVRWLE0aaBQVrGR6
KhosWvIb1S3Mzt4+1MLxDBPgK6MIPQMR+Oam8IIOKI0sGxExOu5Kf5rCjI0ZgyDx
33mFabJFkyTKsYaF/aTUzrqGCks82i2XS1RDXiV62M01ylHWcNZOVHrQ2T/d7/ec
7XPCrziwlcfHhQ3uTqHe7xb1zFuKYyLAxl6dhkIobaZXLdVlqt7OUVHMljsZ0qh2
w3PXympq3y+d4j3Ge9EpS0u4TdUmrHRw19+g3H9tNNn3x6E51AM3IGmGODgndTc5
u3bGfTn7ghERclM8u6KDkF5DXTYoMS0GlXy6n9pwqmQEkEeLOqT14gYPekIMQWyl
rJuYXArLU4gF9103QUIrt84/Jo8AHM0LlJ1IvPArZGc9zzOBtolb/txolMSrZ7SS
7mPGPsv4S7nOEzLVaPCpbFz0E4orp9RgKlRm4202XQTFqGbPBFV7VZTKZV84+9aY
6K4jvRkH24vYf3xtRHcK9s45m1rZIHH3hnVkVRF3cWntB6YW91gQj1WNyWw50iZg
nX+GPlwkHfNiGbmdGGKdLZczLYqrMjE3xSSakFaCeq4mB+8rhKSAdk/2KFwlT7hp
qB/sPMj8SP/NlHhUFzNjcBgHpN6EhZAHu77QK41i46kU1CKU+ZnzFQ2Ehn/3oQmF
9kRe5WjwDA4oDlfcKYktXnad6YPBMaoftC8wTUCDIonRce8NVT6o8ubtLSBEDvvJ
tc4yzmXw2X6LCfiwo4SimAWIUwRid7FQDeWS+iWM9WXgtlwz7SEgbGdTS1iJFvsd
rU7g5Fhfl9cjCrFPSvUVG/3di+HPBqcNxTGxWaIESrUjU+oLfvx0Y3v4ZG+/t2cZ
SCPbWbUrz9Gqoi5CIkPMGPXULNdCXdCwP2jIAB3rRXtOomt8Yly7zlFNVsGZ9AmV
XVHr5alo0cv35E0xbs5Z9UToAHj4oVCxti6HyBX1HRGIaPRHEY/4ZwrU1w95u0zu
5Hww2rndhIHw5g1AHTmLqWPbdjV4++rDH7JiC3aKo2+fzp2MhIqmN2Rw6bb297T6
ZCu5qefNeS4fdNVw+p0XxpIFaV4E9j0xw5BU/36PIKpbViD7xDxbnqGtoXBu6Gu5
BtlenTVuX7kTQW2cz1ZZ/JQ9uq18d8rMkuil2rVdbQA7k7VElWZl4uKMtPdYjg02
aAotneOipoWLC+85/V2edXWQnmlX2A11yiiTcwgwWzBSzgFbnzmySo/0MCQbDGPj
PGu3qbd+C77V+YpmKSnLLd9H/I4FMyl3m5GNM5AYvi9WXTTRSBsog2qmpbA6MzP5
3KH6Y/nh66+tm0Z3bRCOeN1vcLO2dfV3uQETboY3b2ya2EeWwpB8n9Mjcmwirzj+
Ne8Zd3Kv+N+NsLwomjK6ba9lSIDrFi8HvFQItC9xKmn5eFsemMQsnFqLH+Mm8qb+
wkhFadEDfLZ9WKxsz3l56sV1asbxTNNjjgNcsz0M3Dbbn1l90pr5qKrAcCTACtZN
VfVXWEQXFr5DcjWCJd95C4+jb0vCgG+MOm5lxzJFQNSQroW8tGwcxCebv14VUy9N
PZKhk69hXjdtH0fuoy3FG6hgrk3W7MHsKvulHtYqsfeqdqy435YSWS7gjCqg03JQ
XchBWUuPoBo/Q6eJs+2DzwhubYpoVSFzAYiCO2EyDtlrIRARQik78WJJUPZlbhd6
l5GKnW9/CpZP4y1N24IY1ZbmMEVyOVlGliBhkuIuU5ywkkhWtWK0VENaAhVXIe8W
2MSRdQea84o/jGyWH+Sz2Nx+/IeK28oZ2z4Lah0ZaxiTX08jpHZjkS4VcveC72rY
fQQfk3cYidesfEflaSAX1YpaA6+n0rO7Wlloq5xznGYc/MMRQS0Opl1/NJkgXGRp
rdU35c1pfrBzxEiIz52cLTbngLn7RivvugS03+1AWu6Ns2jSLG4hhAvBbEfIEgwu
IC50HAugbeef9nBGE/dhkcPPGIXbZTfp73Oujv+q8+VVQ3IBwRFjGUnlIeN7F+1f
UgyTrPmeqnkVZ445SKIETVHNjb12jfEjYEtTkwS0o/gRl42rk8dmRRVXYXWRzpSc
Qc1bY1UlbLNGU0kbJngj7ihukwLUTkFrFkMpMDdyRnDb0aP6MNvsiNjo2RcKT9B4
l7heT7mzBVF2Z2xMg7y1LVdgAYIgdZpsqzNuv74imqOVbW4cPW3QbuH6MLRwVc+K
9WHNuDE4eVt2QoqHI+wfglzKnqZA7dY0yXooPVl/L3eDXBAgxl2EUzjUpc+iAf4o
7odC/vxtfZA9ypdTd/yMtUDrkg6OPUt59Bs0tDEOzwUctwtPxk7oR+kPYE8k7G/9
FT1xBilyEqkIzsvQsuuym41nMwlcoLc1x0QG8vEDsA6Mm+fXSwMPRA+RGxf5hbay
+/nKtmd3TaQF5W4ohMG9QOKPx6FGno8DHfbzeLmZGVzNCScRusSOq3EW1CmcrsdA
+88vA+fiGzvvrjoA6I+rwgJ3WlWpSVNokmPcXFXlt+sGiaJoo1q4XkIgmqtB3cjC
IiEBaVrb9hM+k3rbDffkQVzocfRY3NWzIn8TYJ24k6fydljeM2Bvp4FejT7QWI2a
XZNuVDkTlJMDCNVs0KiPYJOj89A7BZkX7THc+yEdkOzgHA7fNy5BVeal8wfO70Ht
xvAqRk2sYtkEAsvPit+2qyaR7wrVNgJ+EtSLa32UVP2KQM45eb1vTkTYZd/HKlgp
9tn1GnpUfCpX04VOftcjF5hgvt+DH7irQDy9sVtkQ5p1FmSBStpppvTWw7GB/8X2
FAhMpHP+tlRkU3n8RyJ30ENTf+BpgWhaH3EdMzZqaFEeP8d3uwv4poEKXCtsCGzO
lpW3wuYB6h1+31nhMYTS3LnU7swfg3pNPWIXWTue8fzAKGZ4L8eR1dM7nM+o9Nkh
BukAZbGcdlmXdczyvThFtJwFOdTo4BchQjBFkXbURRM4yMjbphbfAD8AeYBHSaYB
IpRlf3MW1OQwAsowSVmpKqwuYfDG8JXga9/JSHy30rI1TrgmIMezxLz8o5jWiEPo
5752i2l9uMaxyokAQrfDDyenqZrNG+mWxAnUbVKNbek4DY3pgTnvyPnP7ikjOtbH
itwuv4DLwpZGzLJNSUXojE7DH3eUiLQ9W5PKg4mo7FMB27UVmdgzK+ciJdkmiizz
HtLQ6mI10y+CfE7YCN9Buof4c3Ip2QvrnnoTgCPfpSxfAa++OXpcwt5f2zEVAblf
S6oidC99aeZdzu1Pm9Aid5P43NLv95FP77vp6VcbYBWLyEnkMMy59PNccsF+eT3J
Quv6Kg0t7Bb+tMoF5SUs8ntZ7JPI/h/z2sWzGzyjw7ptaGzyuUn3FxZRmNcSLQdh
a1A2ACDvq+5JFxXFhoVKC24cohUJGSZuzHYvtFX5w85c3LyboYNbHe2ySBWSizUf
k+Qm08q988PnSO5iHgZ2mYG3a2GWyeORPQVo2SvIbbRTpZyy21MJyPzI/x+VgX2j
sTgMQOXuBfgu542oIzAL+PNtbWhtB5DKWX/lGmzOYIbu0LxoGtEIrGTZtJCUN+jC
ncG1YuTC2+yXhdUH9q7tKO1yqsnqMpDfNl5TjIys5C01MUxPasRNCwlGMzuDZOdh
S4NhV3DbNm2CTqOqOEHahrLx/3qeu1c+bdydefqeqMrB03QMR2L0qOoH9MnSHagt
JlTjlzHoTuFT4tyxZ0ipsg1Q35n3QEiHlwAwXwPlvDbgXAMlqxAL1kfBWejyIri4
GPWdQujNRkprVJ7cl/bjQsfeQlFiFiAQV1WtcWe+36wXcIBam+M0oB+xHXu1b3EP
PSMfYMgu7NwQ/vcY99K7H7K83AA4tfgx2UTOHzfdySzxA9kM6Sf0RHU1alXD7hYV
lIOWsg/CiW+7YjiW6vZcrbNhnxsEzR0oM45AF/cVvBbr4aMDG1a2s/co1kb7BFHz
ch9LjN0X1vfUOTSEYHe2DvqpusmNJfWraMxvM/BXLfELF7SLLqHloB0r9/DK17ph
Xkdyple5sHVKCq5UJ89JtCwRtIu21MN32AV6Q/AYmz0dhFX/XvW4Y/U+uOw7AfmA
jWTXmHjvbPMErdhaaB8HTFnmHgDXl0cOr5zL5KG0jed6vwoz5eY3/TZ8DOl57XmA
rdATsTbzgqxQIJwXUAT/ww0gYaYykvsE1PHDzuajWTqZ0wTocFvgX8tzhipft6kf
xB3rHSF9jZiOn2FEskDgr5AJwtOO1IULGb7OoNbqL8jj27N+h8KeHQNzs5Oa0l60
5UJQc9XgAp3BRRwiWN+7K8UvF4boiXKX+co3LAfWw40WAOZ57b+m1VTkxI6n4aih
oc55abZzakONsXqJiX+34kGuyGiD79w+PzZgoZ4YRXzvJCwLjsGOL9Qr3tvdDNEF
Z2sG36Xs9oPXHT/Kl9YIiYZ+36Dpt6m+ccYGlZseM+ppns8Q0/SO1Bphmfs370Cd
Nd1DUHH6a4sCOzUzylBg2AprU2mQkdaECTje3KtG3JAzyOyFqIq/VJ8IFuqZYUkS
ahv4J+lJt5IFsjfGoHrmULNW6wqRak6vsYT2HW6MG/HgkG2U9NMG8Uy0jvcAJ7sR
lld0vszJsJPhQjFo9GVKhufnHsh2vI9dEdAlZyBba9de0FbmUCJlipwsETWfzWv9
S65eNmM06YTMgM7bC5ga6ZWz+d9Hjn36zwyVc4rnpnRSqCRHHL9kkaOmMyuFmaal
BDWFsTdUKm2JO0QK3kKFU8xnlvQHmKmzzy7VSODOO+cGQCapOM7TPbppZeLdBPUT
9SlEfxcuEFzHvaEyPyL7zEaAQIwRM7YbVdgzIt75jDU/0e+Z2MVHzRNbEilNLGFM
vRwS2+vzX8eWygcCAilqUJBpbwYEr/t7Q9TCayYtk80uJ5PV9jNqJifIzWrfQJzl
WOIGpKwL3oX9KvJgk+vGpo5grNEkci1U8nGOo4aLhKctdzOALoIumNx9tFj9sKTf
TpWTWaih1AwYv38x+oBeHUbYDvyczQF/KW6KzGj42Idw2tl3eKS/B7vWa10Qo6oH
Y68Hgt2qZ6llQGs34k1vdq0fDavW09I1OwSmDtdN4tPBV5sRcBpJkXnGyJ3ylN2S
G/JBjqD/FLKR1uPP1nGjdxofJ7Qs8Y8XHI+sbC4FFbzLPkIqJ5XxZH5BQdrX1abz
/COZJbjBxaerH2Y1tqy8leQzfmljFzsl5ExBa3bqV39W4UeIdRwcmOgNaMoGL33E
CEXFYXGgoedTJl/0Hm0BGMBpSrvx/7Q6C2VzFEHKXt1GKA9Ll5+Z/zQa1zpw6ks2
a8wYcK+vnEdTeawUVUzGg/mTpkDyfrv/kJTkzY97Vop+bVwvgA5NKUqU47Dm4LaC
GUf16qaQ5sSa+6vVLL/CoKgqO+hMow+Fn3/BCDXxsKmRVXgL3sEO42tdAwNTarTr
+6t0CbWG3KWdJmS6IB2wLJuahsPE1Seb426UxnfmPFuOVYfF1LN/vWjPpJ7mIKqR
o16q7jAFSMYocR/Z01zqkweGYacM/mOid8JIeINOmEAshCZOeufq6pY3fNqAxXO/
qH9HTtUo43rfa1prUW7o7ODb9ngU4+6BWVFTGIixV9lFH2c8QIqdenpOcxjVjx4u
QfpHXlrweDAcLcnJAm/Ba8ckCMqwlzWmGmCWOhSSCPn6/zOMGnBfn5k2U6Azt+aL
VKJFuWeAXK4YxvDLpQZvuQSn0eZeBf2wDtCXg6Iwh9lwwr5K11dqeUQEMbEinEc/
ktgqrVqZrO0tqpgXdjPTxHHb0aMW55RrEv/byhrHY8uCa2uNyfSdxTSxvfiXNq1d
Px30xgVBcNPbcWwRi+5E05/BoWbpVw/7oEuQaNF3uy/GO7av0ZIkmmVgwUe2uuBV
I57Zxy79zPphIt7DK7vFywTUsKjb6MJ9WgTpiyg+yjbAq8eGdiYJP5JpABlLtED+
n1MvZnIsAvFw6k7DZCpKM0lJcCVUKOePwf8qzY3zU0MYwFgOMvyfCqHg6NNkjone
Kb/Fil0I7Gg/yB2GT8oBeJQPKGmrfcGNBZnfDDRgaP0qEOyZeP6OkRYC1HNo9Zdc
bs8m4GvdH5ash6ToU+c2Flk57y86S5pveHjqyIxjOiaD26TZW/XfHSk+4MnqCPi1
iZTCNZ1BcYhOllEsuU+iYrnKCbjsDUqd0ftSLoEQP3GYfwpslNYX6XEdMxqSqh4c
B5agJLppqGrHvlvq8HJ4/0Y1VxRo06JIYl6v/2HSX0aCTgkZ2iKB48tvqHno3K9X
6WVItSP/AjW8UCr3NOhJ2YKWnWAXmJKFdCdylfIWwyWY3/6MIvR+M7gQ8iInEpOw
QWFqm6xCsUqf6r9i5HOJALYR/akwe0efih7QhFQRud3hr4Tyor81zcrGGfXJ23nn
Aw/F0lkHMstW2JZSsojcl5uDy8gQqzOFZ0WAFeUp4CJ4Ls5KQWCvtp1dWlP145tw
bHG/NYejgRGM/zDdmpuMRmvmFtpgUKKMa3W/EiLJczX2RQQI8Msi/8UCwGFc9K6h
QOqi+hcIHftLaWPBI6SFmk5s5PqSZzak/himEUtlGkcFwUoK5POjguCE7JcdCCHh
YMy+gYun+Edsp2FfFKr2gGpGbfFbEVoC3iY9YXOH9ItEu/9SvncF16jwZHLI4Uji
lijaLkGM7s0ZiK4PjROsZIJBWCgKpspjCVeapzeeY3G4qlx9nxgPtNYBdFDuvhgm
2JVpmAFdruNYCIl1LvYj3SAoyp8vb5OkM3lmtnG92uFXGpP6kWRL1py5KnhLzowi
EihZsOoadZjrgIpjd0GSua7vWmqrjA3+hJMeaCr9/bZ9BTOwKtXdJ7LpVnGmxToO
7lXofG96vIcQXkfdOfqDuiCWuAPWJ34ZmE5L/tvP2W3Xycz0vpAFelqbGdKCBS/0
fAz3D19xmStuXVnaVUHL+zdqtI8tqz3VAci2DDSIYXrsbgul1wk02CxrQ5vPa9/I
joUdXC2seOnAk8NBKrnJPXQlP2QDGAsxN2pm3cjYUAEJJITRl2OD2ZVUZ9pVHp2j
N5N175OkjxMJU93++fQV7Vguwn08jBV3V1qDFs3Mj2+4YmDUXXmL0XpAPEMsz+am
/+b/swtZTsXUD7j7xBAMehde9gUsIK0FYlsErZNXJU+2pg1HRc2XXpqX86ho8RcS
z4Hi1qGYDVbZWMncM0PHVj14FeVk47PjuD6hPxOiOX209v1MeuWzaDXcTdUdK1eV
QtxuYXzP1676hjbKDa9VXQDyo4tG+nF9pKn5sF0ubAOJgv4eNU5UDkbyor+Gj5UX
qWmDu7Cnm0+j5xHvFh9n590nAZdAcfnAtzip5/jksBQcrypFN3oGRQj2FMRl7/6v
LQfnYxhwfDHi/31ouu2oXQcy3mTaH4t7FvcWBy5rsYm8cZ4Tv7/nVu2/BCypde0E
XUU5UI7TcQqE0y6Cq1DJ00tlQzjpFJILJObkfl4cgXijR6a0iRla2NjW7s9gN12c
zlF4XripCP1isSIF7KE8AdccxuS6MRw0rA018tG5kgJhSGiS2IrZODpRQ/CJyTa1
DvcMXc5H5fTaMXUhlu2Pxp9Z2QXO01d8aDPeuxKHD7Kz9nYRXOfIkOUHFzQoD8y3
+Tlf331N80B4Pa808XYLXlyCOwxiCxuRgSsDDMSGyk6NEtEd5xzy2u+soa0GmfWG
jEzCPepTPBHSPtIqcZAIDznJv8KntRRQ/NpRkog3FcrVejFJg+/nFuxoZhI22Ulp
t6hbIKb/xu3j30OMvwXWlsrpjkypH8GudFFH1IPYQeZ9ug9+5Ux6kHWkyrJpWA0r
/iJtQAdoe1I62VyYOvxmp60i1tk4azBCk0Ds7crQfscWDV8EpxuA7QJWQf5NvXii
+rqc+CFK+xtoUesH2V4ZWPsYCeEzKXidsLHEnfHMUrYScvnSn92uPcw6D2C7SiR/
zlP9cXZAyGpZskuI7ExMZu7qADLUWO0Zg9RrAjaqBsVpXxjcS4LisgvgnRQ/6z3j
Yl5Yqar0U9k4MRytLXBAeAGw3yO6lNY5MDPhsVEnee85S99Ce1r5vEoqvIn0fWGS
ISRqSmMzR4xi6/5MCssHhmNgFgbXm/rGnUx30KfUJe+LZAPeTvFM/NwSvM8I9g4g
WLmwGB0gmPH17NWkFe0glb9NQ8qw02YlZISHJviQXihid4r/GMMve1osXnIjnaYX
533+UzAmLzy3D1qTtvAdllA0g0VvzQCUFdK5WzXuCBw6bNzUEnHneOcibaRWsW80
yofrulC8In/UO1I4S60oCzjqrnMF/jdH4QA4gvBKUrabZtBkZd352KL9AZoBDVh4
9mQZdywRyb5LjH/bG8C+lSj3t+J4lK68vugkQxPzddrwmqJs5sAOadX0D4smdNys
3qGx8dvcs0wyv4GvkJFA+FJNi0I/+YjZLTJzVG1miINYqdL4Yn+roZ2BXPg5h4tU
1EiuM7By534wa/4P2LoswzsiI0p5TXL2cMwEDral3j/qrD2YRrmBvL2XQ1ev9yFW
z7ksaP/mlOVNGxkAfwdfd945Yq6FyIQ88vbhK4wo4I3+aNbx4zcYTzKQuSzIhPN8
q3JP5Qc8k8T4mLzWn6AcYhzDWKfj7x1S+T2kUexg2taHenIof3kSyWjJuY5JrLXP
jpslvVO8ykspfLkt3fya3jW+0tzKY0Mslzos+n7xu+sSU28w8OLuLXfM7jqncHCp
BW3WKGGrnz79stXkd3eSLcLDUFUc2h0ss1Dm7bfq4QNheJSPDsu6ymp+CcH0rh0m
7A84V3CDewV1eTiQFJ7gk40N4peYJP33rF7Ef+ZJorcsEX8jor06jfQpD8qq1snr
1QOIAiEfgwK1IvJi7OUbYpQ9meS/SnAKQnvTyK48I18GItAAV+dQNPj7ZsMQTduv
2kOXqPZrEcHM0hxuNFd6u9P+bazbnQ6ZzsWx72M9X+MaJK6EiL6Yf1jCPDrhFMJx
NN4kud6v0cbYd5zu35O9qegxOxPZ+cfKX4xxgrbJbwEjc+jUdgsWid6xPVt4kcwx
RyffJJeNTotbRBsj7ybozKnYP2+criUitUW2WQ8tlsTJC+gKsJRk9xt51v/8L4nF
49k8vCyYGvnNla74tj4+sjDnQ4LMfIGY+rheunAXS3KxI1oj+W+BR55GICwh8X4B
6215OnVs/SZS2NWZRS6r29ZgeAyzpEMZkfbwWZMNMpgOlYZ+R0mzid1Osd2k1+Bh
4cBuj0kZeis7XJmRDwDVBM2gqkBasu+zhAMAaMcU/wga62mPDddXrbvQOiOoaiR3
S6ai4OGOBBRQL74ilpaJYyYXx1U+aKVfrj873TZK3Qta3+vxWNSMBeMQW39GhPF/
r1pGX/CwxUnjAHocXGCLt1LrWttTODx6S9e1OLxK2qMelgeafpqV6Yv+mHBzGfKj
baLJ5r2qmxVMtEgTpYIvFZiwG05bRqFfxPNoiuLCc4ZGHEU6iCdLAkp1nGnTlW+A
T/2JeeOJZPgsCAP+j+5fYyVlN+UMz9mI321BLPglh90PKFXiqNlWxE7gwiOBV/df
s9DF5swxST9oOrXkS4TZgL16Sp9UVECt1uePyxgZM2Gf3MpOPvJARLCsoaLl3jCg
+nvDzlYkR6sOuLqcHPGNCJ61sribnxtzxeYOZLwcv51aQ8QA67Q625aYVhBVP3ne
wQ/rv2DPHRnBFyIIGs+/jYyz7L613WYfF5ISCNb60lTEIMq2u4kD6poJBJtPXNBb
IrnNwaVEuUunhGlIOcuby9GOqzvkIrxhuBR6sY2msC41cHKFFYMTCUNNIzz3lKAa
4DwpRQA9602LMXAAk0j/q+6yjkpb3Vrz6DYWE81+78S0rMnPQNxaXeDbkZ1ZuONU
cRc1Q0FCswb4lzsnm3d/eU8n6/kbuk+nvjdGTXORidWdVKpjLrDSZfzg08v8uq/O
zFkBIdZn6GR1kMEg472mAaXlJag0Y5K9xRiAe5OvyY/Fjd7iJ34YRznFniNVDvrc
dx81sU0uTO+V5EUIBRa+q4DI+0Jfbz8r39pySw5r2WSJJE2T4UrByfwnkUNkdFLE
mXvzG+LabKt3dcL68MQ9trlOqsRUWQSxAPIZJyEW9sZilbZ6/2vp+Pz2X+fgMvnt
GbMGOzxT8LaegLwPavb4ksvmuabSfWD/PAU9ggaDAoSpxETtrCFgf27c51wRP9ct
3l1Z5a5nWGai8TKvFEzHXMaUlbQ/xVZ88R1sJiLPMa8ppfGD1wb2fClTNIFhqWlp
pomCm+cZrtD3oMGJhMsSFLeaM6qS9uT138Inw5CzH1dcqS/NdlZzA3YmjafpQMLL
HkHhISwhUKss1xuXsDf3f8n/LdxOw0aZgesMlZ7L0/vYcgknaiLSC7sa7DebKac9
hUF0x4ts5Cjww4Ke7roFyde9+jTDYQoS8+mYHeOnCcQlBwRonzeMkSdIUYuwq+7a
VxL6Wc21sLZcMn3We0lJmQvXY/yHnKQOMS+KxB5jIAbDViQuwlFWOqSYfDQYRKu/
3yBG4yNKLodJ227qFTKTJuF57a7K3cLBFVzuJY6lTafX6Dz+khpRvylFZYswkyxy
mmFhttrrV6JCy8hSEYf8J8lCR5+11BRRxdnK5nOAPLfYMQKY8AuE7x6PY2tn9t72
7poRza+JORvkzEwPMkDyrYvu00jNjY1+TgM4TySrS9T5zJQ1zbznXJWXa381IVk0
L9U+fhFyslrQBiX057S8fvhMX3EjTRwLDdFqQJ2IUBdLhpVOk/S+ShviM2I+2/2E
e3H+7nLwS8JccJgujavs1cU16+iEu5PD+1CxnlJTPpDK0sPrdkFXVqFwPconvyGP
CizYJUEr1VUqOMGGEd2XVkK/2n7uXMAUPd2tedcNTKlx/waRitxiCdrI3xV5ynPN
jui/jjdMGO7DPOS5xnUD20yY8fWgNnd7aXF6p84VTtFt+9fj8xv5aFR9XEdm4XhQ
KoDmFOCpIqk6fo7WSmY2ZNziTlClxE1zkbWGneFQGgfF/+M7gaoG/h2q0X/Sjb2x
zg9NVFngEnZ9lK8sEpHn1MS5KQeSL68G8TCjAQaK0uRD5sAxWPeiwuTgFU5Frc5w
0qXeS9ZHY6Zk0jam6tJlmvZOpV9NrqEFvU9g8mMkKCMPqLEiWJehdk10fxF0Vede
crfXQzh9srAzJC0nSZnxN7SkuPbtXIv0Z7XYaP89njyDwk9NHhL4V8lDtHWPZHMT
luUtAggF8eGjWNl7ktC9Vc0O5H7V4hM8rxPAhNUNkOZ5Ss6OtiPvHbVAeyqGwjut
tqHKDb9llreXtzLd0Kp2Ga2lHSPkFbUBwsSBrzng1EDW4xm1ZfgQk/iWnmxrjcmI
bk/N8GfGqDrspPaH3i1P4JXc5L8Ht883yNqTP8pD84yOWhq/8Xsz9gO5K9mo3KEW
saE1A9yh8IDzw+cc1Sl0UJzgpku+nFVjFwrflrhVGeelKQIAOT61pBo7qiSG/3lZ
EQXyv7veFgrRCKWjcgnsgKa8dmi/nL10PZunGWzDiS1AfkaNTtjipP5FLBvGtGdZ
0GlqNfgB04SmFZBEryXVO/MNiMTNgNSLPuI3MGH7m6ga2LGZcaFa/8h4FDCIh6Gr
jmUtpbFPwkR40e+mwnHceVoDTzCY5XgC+scNFy7ql859/LHUewgf6065xd2jmRdE
R6VfkLqQjWaUPzi6pynMWHVtesiAKELzYX6gtZs1DQAp9HsJy7pL1Z7C2D+jMu4u
eNGCPqiAtT4ZhN8tJfBGCRTTdNvUTB+5kUBimRiJ+sJHOiotH7sBc90UDDs4CQBM
Jii+QCw7OndxXlDMvy2/abL2ZAeFp9xBarMylaSv1CzpQ4o/DugDhBsKLc2LhzZW
dBHjiQU30+eWkonTAkemk25f3100kcWl5FIuExbdepmWut1de/TCiolLwCr6BFgF
gKwmt/JCKEYJ2XTEXOWXA/jUnmUGn0ltqTMC7ItU4MzTMkZuZ/GUO++CguU9ZyuB
8nCJDzjWBi+Vr0hTnKdf0K9IkW3ZNrpcW3fWdJSGgVl246cHk+u2zaRpTjYc144p
xtW+A2IsBBoTIeWaePC6Wv2xF4LFJaW7wI0CT6BGAuZNIgN/K27NAI9MewHqFveh
MmfO111EHO0tY8NW3FFYvscvQ5sii78iB5J5G2gx2osjjDZdILeUbIaePwpksiry
N5+poy5kYPeXHOx2xXWWK9sD2sIA72HQQV0VkUdPWd3KpUUzRrpPopxxwX2fONCG
LrhPEbyiUQmlRIK/4MwpcUq/2RzesKYF/Rz8wObaX4sG4i7mZW8h9bKmYT2Hg41A
fT1WoluwhKFCPJ2P8VX2/aE0t5ndYGdBhYKldxxMjzMXatj148YJccOzB0P9YuwP
GiUsOg7n6Uo15RvFqVk33V1B0nj/uIFu9tmEltXFp0GLLkrKOrSQhQernIPGzxKr
uphaXq+gNBj5lCnrYclLa7aDoOjzHDKO2xQxz3yksK+xGeIblMh2wR655JxY5wcE
FPMdhH0txuBqnzZcHMDnQqWf+HEErTWqCPqdGC+NehWa7akE7N/CR8XNLCUijkFN
O8hKnSDGuRYZJMxKR+et6fGLiexr8StcjEFYbRoENQQtCu0xoFFj+G1XCZ7ZErtA
TWZmB7L11QnoFQ5iMxX3Ik4Nst3SBbWYmd1NgM32SUr+hVUklJmx5OtQSwUgk4jr
Drmg7LaLNwFUIhi6cdB6l6B0Xw2k+4Jgk45Xus5wk/qYMW1qpxltVMlCmdKcZ0am
VuP3aP1AyEHov7leHicobXuoyGhoh1XfHa3Pl6NMC2QhBGOvdQpQWUR+AOM3sIkk
/FU9ZW7U+ThuX1hUiYq22+Cm/+07/qA4kBPsU2U2qS/CrHzzC8+nBuZpHBa2BraU
2vCR2lk/L7HjVXSmQ6SM/Nu/ONkXdOVUhTQCOTac8VHZo/oUSYk24rBqwFwyG5FN
xW5kz+npEAqaxembkkkFP9Z0wBfchgIfkI6MC15yz6NkbA0nckoDUMOaRX4QhYXe
C+Rk7VQRKNGsNvOuaJi4W4MI1rAxVAoWktKtPMt73pWEKOxWOrTmD71kbZgZ+iMa
s1QjSQmDuuSYx4SAhSG5BDppIJ84w5deM6VYiDeCD5wIkfXkh7InM0WqurZzNYpS
Cfe9J7NXAuMhijHqNUTWuVLB6WXnfWA/QK+gQPk9Qgv8rP285/qKFfPmaP/FjJqS
zppDfJWuw7UE8nHybTLXl1XoE21qj8EHeNsr1/GiBiL2ScIJyWpcbBJfvmyKL/EV
JenVwMrnCg6nQaX1kfRxG06yTC3DuSzAOQ2mEuF0XCJ2lmS4zP4vyft8Dc8yKvSO
7MomA9vEppjlgZSKIasNx6dAx+XrGTY1Vx1PgDi0R1Rs03RGt1bfmLHuXhWYCrj1
pFz9whd/C/VoFkOyUoEi+KYyKhIHv98dZL79qgjErvALA57QI8lVdSX/HgvHqmMa
FVhjmOqrsNCLImzXZAt4XQ6TdIDsH/qKA4+sXcj6Vm+saVEp4mDo4jhChfob3yPB
U11kNda5MMFDtF/Zmr6WmPwwiGJj2uOuWtAPduPENoAKElWeYZ08Q9z52VrNpT6H
bvzD9dfVv/Vt2y0ax4WOjPk/Xdjk5/txfBOLMVMAVg9w9ylR8E5Z6L5ckzpKyxaY
+jZozagl0rI6dN8mH0RzCkIgn3Kr1sq30DiDUFNJ59Ffzt+BtnwaS6A5gBpO+kvj
Sr4eC02Ou7OIFrbrk7HDkseHAM+OLdHrG0X3b3qX1at4VCAwxVFmTKSnFmqtEVsI
QLAV0A4QfW81MxqSjNviEnokFA1/Pe+lFARbkYZVtbgMDJA20/C60o1oR2UOOgbV
6JQ0RmYG9dbCA43dpJXEWPUWurF5vPDp94DAiO7trGRy76uv8whEUWXBZ6wRvwxt
H4BG2uMe/sjxE9uKtjo5cYUEcDznx4UUY9pAvHoVsCxzWXjNXX9io0uJUHdKdJpb
u4nslk20ajBDqj2v202bHjC7i0lfPEqPCGIuLAJtjCfF+EoMpsK6xGlS+MFjRf/K
5TyuDlidUwUwmGp28XsQs5OefJbr+hpXH7aFzliPHnX7idk96bf3wNo9KPNBSnAm
T5YZslp4m5+4xuVzb1ZsnsuvTSPca1KecZxBjBsCnQNgHtW7WWHqH+E2ejobzBAu
Yv6hdQwZ661mSt3Tryc3Zo683QbMFClEZFxajl2lEn4R9XfpEI5jGSZcMQDqeVC4
3M8Jt4v1KaPmRKCzsxE7QaQbIyGeAzhDTMOhJU0187KJYwuB7TDsJMnwnikLUa6Q
ceQoN6dtaT61VU9FMad6n65g6pLBTLpFT/rUtS9bBwiev4dME9+xfZtaJL7m6Jha
VaBGSOS6TC5x3lQmhU1rxnkJCojL/AeAjZVITFYoz4fwPO3kH4OA84Y4fIcBDPMm
8SmAoM4yAIz7mLO/TF3f8Supo/x8SpH5CFV1jzEy6amHVaPpylJUlv5PaEjGvcGe
PY0JEO7xWynOt83JoTHm+HNcA1nY1ITL2YYl0xIe1QbAp9a/hE3SF/TajN0Zkk5U
tpDieYVOiAJ6B0/RbI5qQtIG0Sbnrz2eBX2/TvC23qq+YMsEuMsohT2aV6Cjh7et
GKPDRnmrYv4SbFMyjlnvYzdGOHvJFZNSfs2fusLqMc0/JCe66N6TmIs6lXLWHUbi
nOmFZPXfh4GTCQY5cm0eWUqI9qso69NVJkjyf6nxSbFTCMv2olwKngGRxDL4yUzg
OC6zacOFb0dNP7WvUUzNZBqpriRwt4Ralyxh/YYT/zaHR0LGnGHpUQrSMcXNfCW5
6TMc/MVeLdN3i7oJsRRjA7Sg+Bu14EqWFG/5ZvSoG1z/o6Ex9Y5LA7mVOXi52x1g
ceSE0ffV2Ly1xloT5bDGhA+QwoLxRAUwDD3cnxHRgT7+uYVD55+zW/8NnQN2DGiE
8KWUW6IsdUuK5GnpUU9biHMnZeQVgw6vHmxReLOC7Ll4M1lWK+0AiluryDHOP1da
AL4FbsJQd0XqJRq11wP+fs2ZDGIIhAV+LoXxZHWwtieiNNMmMJyQX+0FVsi7+mrw
yRNVASC5rYUnQunEzIHi7uFKm+og9l5T+SO9BhGU6xR+ZdJiE/IGcX34gA1Mog+N
tzoPyE7bHsbGjdvPMeMAtFdwXW/c2ABIyNCCoKpXcC6cIFlsUhKgqtPqAHXIu1R0
xkba1XNxXdTbKsLMQ0t4f97kz3dW8KiD6HdXsVBT6vu0oXgN3qivCHtEhBnU2ZgU
5hTYAlVvhJI2Vg6asSdhB1e304LtAh2HOecdYgU5KXRnD5Q8HDpBbz1khUs/cHsk
/e3PYiOWwelZUiCpBr9LjdcTHXsNlpvc+uwI6dvMU9N8Kd4IK7BYfQRH8mpRKbaj
G/TsMPHsH7UsyqwTkX/M5MhXAQRQdsCgq4OJx2hoJJ6Ilan6fjcpaH3xg628/VFn
d8Lmx2eS5WH77EDMoZASkczBnngdFvC46sPBWoPAPEsUzv51Lbs69pTGNaWkmaTe
bsEuoAP0ZDsOjSXWyv+63XucJvK584ahrlwbEjpc51O9fnmaKZO7n9zyGwYSA4Ne
OLq2boU2usTc4R98QUxoDrv/jZqqhRoXNLdEXhmPJdDZHFBCDxnD15vrX+GdHhGF
RxXPPwlXaWMYAai1fneEGp4xPiTOWRw7CpQyN2/nxw55yQ67WGVR3X5lp0J5hpYP
nVwFevFksp7uTSouX8mDyLKN98iO9KIVXtrBdS65TOnu5i9qaMXGaORS0QTyp6sv
jyXbckCydWeL47ZQnq2YXxI2Xmg1b6vQFRlylIVtOc5Mn6bqkixWtt3AehQhp1dQ
NZO+KlESeyNqPqadIFetbw/BrhyIyKAFBMMPUZ3IE8pN6g8bBNUExqZdZeO7icvO
Gr1JQB+DKTTB3ZfFeW2QuwI6d1+MqqH8o44J7HMqKQY2oi8soQbrawo70KoCDd4Z
rfy7OTMMzkUkG6NGsQ/fDQ+7t+nO2LTEhppIpTDubdPi1kC5b37mbooUL2rjb0LW
4uW4TpiPaOcZOQ+vngWnPhNhKibv2+qAKaQf6pN0whc9K4G6avv+umooPFsm8t2S
UsuMS06VOR6zUyEWxfRBW3qOLnFAEt3TJ/asqsulZsF7PZGUDANkgbHXxirFI95J
J7GT85pkfQYAe+o9v5+6t6ndLWr8Y+fGngrEXuEXg6mV9XbkibG+r7na3MS1PCbn
Cw/z3hy8Eqd6P22lTauRmPgQ04rcwFLznEjMFAAhgZ7QjzrSpO/ubk6nS9UIulvi
mDmW0Oj+AOgN/nCBhAz1oV5d1nd5P3Js8wt/J50ijNwOBm4x6P5D2eoN+TPgPdnu
Vfs9X8MoNhHc0ogSb1eTRiDsm0VNs7RGjlR6cQAYKiLJcLE6N3iMBB+Axn5DJlQS
MHcTsdzlePIkF+4HmioPhMMw9hu8r+L4SxJGfPaR/7hA0An+wPtWwjTfe3OuCNjG
nBCpnvCShrdAjGhbr47xUX3zg9zaxyItGbtt1m6mdg3V9H1Z8E3dUX6z+lCxbnUz
X9dCue1t8Whgy2levsRs2br1GLzh9iJgDJWbYfuuLin3f1eoIKUsffqWy+cYkrMo
s/61yFY73Pikjzj1/2IMRyrIV/bldcggvSwWXmGmtJEGvPSrWBlaL2Lxy5VcQG7v
6ExR0hkc/Am2CZYFHC5JeyzF3f/zshVZEWAXc8bg0G3Z0qhuF5p4YRqucLG8dF9y
pdG/WsyEjVtmAFvux+CeHdkZrdqHm2C/P3MPhadW7/d49GhUQxx7Ghqv0R44yK1f
SVcibWZht+bGlO9AWyQXEau0nx7cbrClksefN8vjf3xmGSkjhOy1gaLmRCtNohAy
zJexWpWVrkWQu9d4CaaOhZgxvhiXr2T0GYkKKfSAGsfp+wEp3kPiXR9zB+vlZK6l
dP5tbQyIogNot/c5acZai6Li2C+FXRABSab0Cv/iRXPoPxb4IRVUcY1S6kcj/VLs
JbmTa1DpNJCbLApxvwW3KzG8np2oIzSEkP+v+MGCEbl7PCM+gck25hhxhhAmLI/j
c9AUYZpt3QbQ4EnXo6uy7XImhXrPRV/k6tP95EYXFOoDPvoet9KvKK16WbbIHgk3
KRNBN0mTO9AvEXnD+1d1BSNfB7mr8cfpTQttGr9jDA3t4RH8SSQOjxDHOkZ7cS3d
VZaDWlxoKswA23LCwFSJiy7HKQBT0Hz0AbgKtmdgefd41st7H2y/ofUsTGWEnm1H
rJ8hjliZEJYb6cgIVnDg+y+Mc27aSSgeJz9evJGoFOlHEKya+9jjn+niK+TPXk12
ObY6WR7YtcdT+sHj6Lp09+ix0BoTSwjkcvaRIimLzct5lUyskHmXy/jmS8CUhUZN
SyidGJ4ZIp/6eDPdHZZ0BlkUWuEZWZzJmA+GY4kMl+PGJ42KTgI4Iu9IxMYNpNx1
2cXO2Epr53Wz5jZJqHZn9VNZJYMYT/b0xkTACd0R54TXxbz3BpWZEsKi2SfKU9Em
Bt02XEWnwicRVKKkQHPMQM/InUEdBRm+p4DMj0umnPSZ2ZnutOZ5MWfnQIcrLlZ4
KLT01XYcwv5XDuD8L+xaEmDCZfgIjk+a0u/RwnLji4yB+XJGbTLiNeK2jVDy7HFM
IFYBcewpV6y+6vwUAzFtPxT0R31agS6o128FEsqhmwiA6OnIkpBQ+8WyFYC3n0qY
OLFsb/31aF1hwMSH6UWt6w0ByrpB4Lqy4N03h7PQBL2vCGNXqjm+pSyhbHxCOMu8
hpCkb/iNKbW3dzGb5051Xa2zVYN5AS9vtrIPp+bCwMINQADIojBXmCt1FjrzrsvW
3LcqtvF8nrgtdNIww0c79lPG1t0GJCZxktqr4q1m52wSzB6akFVkPucA0dLWMZYx
2BZ4U/ZBx1htZ+erEA22vqjaBOnclJUuWivmxJnFIjL76dBrdi+skTJnkhZG0gRh
OOeELoPSGmIC8GQPjQGhx5Wf9f3wDyXS/gZn3iqDs9lRw3psKxvBUWHNJjMEWWin
B1Ra/bU05vbTFGo5dBHg2E35Hr2APo5HuP0WcZPDSvMyROYkGfsS5IOMVwmM3REy
j6fzBv49QTlEpXcFrIZDaqWqSLAXneE0Oysq7y7wNoOOEQvXNwgWuqZ2B6z47Gbf
8OswBNFC6t+GUIKuLLeJW6oF//4wQpV2HeCetqw5pOG45IzHjnK8Jcov9bWpZUpQ
1rNnQ2B2Lc/C1uB7e1Wx3iA9tXqr6S0d4r0Hg1OFQ7P3z3T5s/1aTrU3WTF89WX9
7dfLVePMBO5bqdP6yo8VmrzFCjoLvZu0gEhfs0X/+laQWS1k7GGk6G+RSG2O81fO
JvA0ch7d66IWO5sDl44ME7bJlQBY+OFvGBgPeGIqtPLGbPMSVbQcmmTGc3OMOusO
Qq+neYL4M17+gtT6M5kBFHQoMaoeDy7ESQ3BjdQL37GWHKbntn3XLY7bIm4dgndb
jOH+XXjVzzl3F6aV6WA2EnUu6rTv4g10AzaKwNx/97xeS+SAgK5RPhOy+7E4vgre
+X93yquTbZ+ZegzgeLLZBzeNt+Jyn39ZNJxKPva4tpkLyYl1t/j/WPLQy3KVVCb9
73HTaowM2NN5CNq/AFs4YZKle3RoAkP14PAS8X0k8w3Z4XTDiqdRqELAb9G3hNG5
1q/Z8Ep35j++70X87Pok4Kjctu7rVFVWYY4R8Twm32VFqI22+oDaoLPqVmsUfNAu
8tXPNc7ui+DGv3ctu7WhVmDOJzXx3Q8gduOyAI6ldduGboMWOP4oWxrYAW06jC1D
LIhftBZAPczAj7PLfRk6A1RItyJYYJB9gKnMijuF2BXygRmgKQ3kIWChql3JDUMO
rrNSQ0vUnrpzYgInkwS6T/lBuDMSeBO/sBqIcno8gGwjJYL27j+AS1jkk0MNVHzI
ZZ1wWd/sKdrXze4bQOMt7+c1uqQFvzIcxJ7oVjNfP1SFDS7hwx5VtdTwK5EY3bxT
6mB4dYA4aalgTWW/07Z11eXMAsAw0sYxcOK7f6xDYbM4FPQXycGOKPKPOzX6Xk7z
9vodKPSToDzJXqva6uXbfwhkTDi8L8srC82upUF/mxHnJyMo4J6JFwQl09CKyfQE
oYbJUvhLdpuk3gm+dx6JJslFTCpelUkTzXmJae8uR20h4I9QjSGyLMpPte+zvXvD
5s0kMQtAHESRCdszDdFEp4vyqOKohzk7R/Ie+VOl5MFJLEodkUfj5Hr8fcNV4KLi
1otyzRRJAd+NaXh08B7ppOsn74x2O9J4VpgGIm4PCDlk8zdLQL8Qz2++yrfEuNAx
+ucsidgqxGdaAJXUeRZjhryQTVrZTCfSAgz8Pas86ZILNWBfgCO01OEFzBlN1HfT
xT9wsa3Mmj/187JtEGCOvJzssIxFJFpjkUl9oeXf1nmB1F0ohVnE1nglfVomOnaq
bPlT2+CR9c6LK9Fz6oVt/Hz0Css+ujxDqbt0dvYZ9Tlrt55lV0rYBQnY0sy+Gzuh
PMrXyL2bROco09DSq2aWZwPsXB/1Fe86CP7yrnFo+F/h1zRKPMxFLOHYqe6hdADc
v3JZovX5PRJo4RDf9vztAa2226aHjzFbvGhDU3hxW/ND87yH/5RHpY8ZYHq1feCO
6brA87MIDBqrX8+2HruFvPPtRNnE859ohmr+zVVUMTcDfX0AnWhRtj4SWjgW8Auk
sXI6DHX+NIoLRXqArRsejW7u+fO7xks0MSZjxlKkNxdYYxhf94jdSeFhlVn3yiGs
o7uPnIc1oTG/z9p6bXZBQtON4oGl0wBCF3gYOm7rcqiCuTDqo19rjS2a3zGNogEv
LT1rUt50hKT02IL0HIH44V46Y8hxWXEmkVc4n3FwLSqCtmbDNr9GK/SOddy0AKWf
dkkrqNQHDs9C7Xx7uEORJZ55GXp+uF5+JO4CGEcSZErbYsNa9eLM847TxJU8HDSk
FlfmyxloEtBWAQEH8qvBbANHSVkorcJ1pBFlIQcChXgbHeRQK5cVTeA5Aqonv7Ww
PeGoP4M8ouvbyAr+XjSjheoUveQVWqswRJVa+O81j8Z1y1hGcAWNLrDEyvi0+1Pc
eobRWHs9zRS0AFohQ6cGbj4Tlghb3qfwAzYVF72q9GVEjnJu6UQzzqmLP4J7fd91
0iVyhCizXjQJq8Pt3Uc0JnYtBmMj8wilqrNLgf8XbN5mfM24Mx049yZs0EXoDMK2
WJeF+wmBas7vumU8jaJDv0r42InRlcNtGtbSxAIAmltgx1CDOtW9Rir2+WGrPi4L
NBEpQN0GvHn2tZxzJsQ/IZ3VMT5t3aVDbwywDsc23Q6/QhKw63L3vO0gqi4/JFMQ
T9fdJxVaXetvju6okq6FKh5mujPHEvCVbBEt24ofCvaJZlJyWVq7qs1UstXRJmXp
HZk7lKQRqq1xkNiHiOASCadi7x3KG4gDEXSGhSUKZkijYTKeRxW69nq7jgX6plJo
3a2+bdgNFZvLfG9P8yOQ+kO0HjqwuThAMMCiP02lcRHpatXOE9jGdS6oNy2f89Ak
yPo92Dk6IkdUexw/7gdpqIHzxSHqa1yjH539izlENmAVCYIV2UeBrZ+y6zt7KV5t
pfmgrtAlPtsGlgaUHb7yPuVaDJgIUSPOJvGvixLJO7GTt9GDqy0+ffdAHSLuenKs
e1hhZz690j9X2md7jaPyHbHWfC7n3p+pp4s5jOs4VI2WhM9jMW5gcKRszKBCRAKa
SFrVMLlhNdlAM7abaYAtopqMhXweRGxaRAt2vn+E4S9I/z9k635td4a7iSGaXNzB
8DgkWS0CUlBdvg02ykRYRNtUAk0IgXuEnTEHxzcdhnM4LX1mfSRqNfMnmru06CBP
IgOSFza+pnER6yw6sWBbQwCq8IocuTHBG1UCibqlhUbtpzYqqjDqiItmifM46K4O
qzi2QBe6yOW3b82emwn+ub19pn759Kl/MoT5uS3WXIYUrxri6UtcokNBjHguC4d8
xy3h9TnsDKJCpiluxVY4I/76I5q1DeGWNIbLxQewuKNARc1lTpUTLk97JF0yijCv
zd4EGkCCZI6R3t5+t6l2CKod+pgjvvQ6mJxxfUpeWLWG8/sNZWXAEbR6TqRLH51w
do27B0o5Ti6pTKHTDcCac9F3SzEZvLQiz4kTWrKJgPja/SM4QjsRRgDAi7kISW8v
Z1yBlus2e8o/8AXmWcz0AQ+uUNhnaPcoHQG/ABVm4AKZ7alAUTgf8mOBdHt06tQ6
q3sjvIK22NtjeTg9r5xI+36Hi08qdczlbMlhoBPp8hpk2TO0R4U9YuEy/ZOK7qfH
EPg5nuAlyp2UGBQ8FKOTLkcqcLuJogNJMJGnp80G7N0xwkCFvjKD/mDAHcyo2G79
HHas+Ug0wk+Hza3tWf1eK6NNJkDHvbku0M+tXuxYaA84Dan3aK8nVaERFjMhlZkg
wCT2zgwhFX6jJ54Ccyvge65D4wXzqsH2CXsygR4tw2PrUtRjFpceQ7Bwn/TDKOPt
TYK5lQW58V1xbuDMQ+fw1MBvSgP4HKsY87nngqiL71kwxvVOtotv03GHGkVQQeMH
UKGKZnF6BwqqJIHXTeveX8iycpxwftquh2VDJDJufpngBZs/cZRDjT0zgIRdvGrX
BcLe3A9uKoJwWLiRQH6a9H/npxJAIcjaCgnRgIALS5Y3qc3oSrJZ+ms7gRhAT7zs
jENoR6r1tD7sDU7JxN+v6vlK75xsypB/7xkFGMs7a1fuL6DzJ1D9PkIlWJwHM4lH
KCPmjFx01ihG6Gpv2hfhZfxAjIVdhzTo76KsHmZOW+0m4mKC0ZuqE4qRFxPg6TAp
hIgPtx/+am5r6H/MOwaykMolElgxUvvMMb/Z/Ncp1EFE4jCDTyLKyglXV1STSZH1
bU17JvxP9KWoJFw4LfKEGns6YFajwkvyqTNJ8er2gYz3vrn7ja/7xW8hA91TUeKt
lxfyyTg94ADt0wVIRsTuPIOwWJfxNRu7rhoIbGVYv1JHudzyw0d4un3p7xopVEJo
CtVoBsjuV0hTxMoloKZrGwYzJ9TW6hTsj+jlchrRh3DDyJlnhGS9cKnWLwHpIWa7
lIY6hOMMavUp8LijGAUK5IAcKlMTHDUm5+tzZ+bxwvX6fzpBlA1HXy6oKRZ1Vlda
WICX7nwA1+NhsH6DGp3vf0QHSAmrOWoJ7iuy+TfuXn9ljbaPyT433WNlVEeujniV
kz5xLvrIedwPKU7MmQBj+v5TD6VhVIzyqvDkRlXjTFsMawA0sgU2kre2u0LpVoCT
GD8XwtrrnbigDaOqATMN4r7uhpBKPk2tOWpkvWBFUHtV7aQiIIK4C61SiToZNmBa
3cZxmEs9vbWSaIRdtSnLGnEMuzh9aGDZwsZVcy9XpXRX3+7TKuM3gIy4nQxHLEWV
bnwJ/a0DThNzzFpg2hJIk/QPUVIWpmKi/zHRDDshHI7/o7cQGkdHHmVS4lsF3FAo
D/OEkFRKFzXYIEUMrEGXk6w04f72BedaP3Psfwpc2d54V4YXp+rCoFLCX38AVDWV
FRktx/c13hUK5H3VNe01q6pBtDwD7655wMnkUXTFuP4aoR4Pvz8+kTD4IfaO7yEp
P0uKwXnyo09cF+0d9dvXA98ravX2C++dSBBBqlYKG53V++M8ioLV0xNLClI5dI4j
fp5ZINneX+WL7cq7bZDDKuIwkwLD/Z+ZerL5OSGRNpqCKatnLDsxkwYMAYBzA+Iv
1C01jJ4h2uw4S9TOZOvwIS1e2ARLbCrRceuu1BMgukQVSaDgjO+iUwEjevA4l5RV
DHRGQecxruagBzZuIkN70kUTAXadfx1uLePUcTCbsQnwBPDYwYeCa3XyAA1UpZaF
ZaCqA5f6TMyibNPkutyXgkgHS3MCw2NqvyX4uQ55ZcMUFUaIzcGJN0Ukak+6krjA
txUZkyyEXfjwBfqH2RFAncd7SpYkIpH+4b5JKmJMyT214Qvmmhzmkido1Oqapuvu
P5dw8lUCdULwbq0bb+tlkIFodzZaV+rdPbPj25Gj68Ru6bd5DTsCT9M/KJQhbsJ6
KY2DPifHduJt9dBvyGZMa4uC7LtZgeAtvEiKDIib0CEhTYuFyyRv3n0OjrTKWOMd
UeAlgCca+o6rqWsI9yGGx2EtBUWFj1GB1IYXwQ5nvXRbN1o6WF6HIM63RwnxcjYJ
JDFFPSTU0npBWMs7jnTmS8uEPjniDN/WBwADqPDiXb5/UqZfcVSVnuZjOoXSGKAG
JF49Tc9nrBsZ/tfj/xroqLLzI53B1WW413Gcmis74OEuENJRgTJbGrkz9vPybiFX
F3bAx2+vYdSAv4J+fFWtHyEz4OnAIR3WdaWDCvSSPblooF1HK1cYW0+hh9ZeLn1a
CYHTY1MTvfRBXO8oxguPHht1Ofpn8DoINqGyqMpg8SXOFTbd1LVJ56faSjmcyRpZ
KW5ykRUaiwLhCNUJ5KtXn8LSdUXJUQ3AqJO5FsUKKtxUTWheq5O/ahGdX71Bxlv/
P6/olu913+vOTMh3i9DrabbqFfYdnOqLSMW1q2W6oPbQILLYd+l6HVAuL8mJgtgx
KlorcazWnzXIKHsocHzKT88sTSQWi0p4FLgK98Sv95m8RkuCvykSTC9K15SO9irf
RgPvyMFPPjl+QsggPBjfmY4t71JELQXTaXK8Dco6yRFZzsnyznAbpZSt8AqECTEh
4a5pXi151jgvVWj+LcZ4GS/RjoxwdiPeI3MgCN0Pk47DTjo2sSRIN5V5iG2GewSe
9zdlRVPvQ5s6xlZFWBGdWZd2usTBQYCyk7YTrrwyjUPlnVeiP3aH9Jncq67K2LhY
BlgzBUsKJrYnbiMvO4CbvYJHpO6BJyd2SB24Mf6TV6iB0DF10rn3LUBkrM/sjK9X
ja/bDMibhAojL4ERtSCmZ3HzLKBmPas2MNc2YdMdQhjKbw/Sr04hKVfIKXZ4766a
h3otBUCD3zHTpMMyQrfM2DVVP13jtrHwniERoEBAsXWJfOapcY46nUWNTIJ9IR3k
xbm8zi6/HogEnS9O/kiRa43OwT0NdzvpfTjeMwSTomJqila32U1zX2jHublKoxgC
1yLCvaChV3083Rnxca36UyQzmfu+sUxiJS61OBdqFKXI3DEbfjVGy5hfYns1Rm9h
/wg5PbYelZs6SU+dWgCMYlWjCJYW5Yk3Q3/6Ij7WTC28EV8Lj18H2ioMGgTjTfy/
sPrL37+PyIhsCed60fN5TEMBnczYqlxeCh8xH7VUbChgmg1UgyZX+8+/EhQj4ihR
WYvf1Hp2ejSJV4yt9MQO/hwyeI99MmL00ynSHvZsZpuXsYuCvP3oMensZd+qDd0A
aKFF1JgNX1/9AfIlC4S+BbWtkcQQR22QPRL9KhWlcSeWE6Q1FSkG7Zt/U5c/iBHt
DZ+sZ/oQciM7q8Cg30LHgOgphDDEQgcntqpruhdRX7nq2zvw1nQL3bgDg/+ofX/0
5nRIaVg/jR2NgSY9oPVIgxndZj43qPrNugvjEZkUNpz4HbKFHJ0ywKW8lAEZQOjd
5W9YA4yBdDifAHJZ/OY1CZ1Vrk3oTTtgIpRjaCFn1hMHwwo6rI3GI6UUDD/ZHDk7
o10+S3P6bKyyLTO50zavTKXMI6B0cqjy+nAX3wV188ooR39PHgROd0Y34/yiCNuZ
OVeUeelXGnvg1hJFS3m+YHzuz0jvltUC/k/0CO+SoRBq/iSxrCCVp8jBzJlKT/7T
7Cxl/n5tp+fAAw8zpBoX8EFBSn1v4TFlJKjZVYGUAKVqsDqmrqDGFPyFfBchoq8e
MB5+FEIWOplt9orRcGrwm4nzPUeoLHdnzfVS9r7S7OJNCPRkMpdF5TlGooAMBbrk
Vprn+u0BB1Zxwwk98HGwhCYr4+iz844tN5jt9kaXAnbFzKG3a0LvykRbhdYQR9iF
tWg6Xsaz82LWSeg0+ab0dWXF0+DQouIqLAtbRWTHIqukIIxiMxu3Oxg/zC2ChnQc
peCUW/fciwkqmU+z6mIANyezkEuWfx7IzdrJ38byy1gQ4BmHxuSRoiPocO4dzhTj
gagdqFShh35ebNkbOYuDs2Nr3OD1RAHEli3CYd232nvgKL+y70EVWs7w0VvvbtfM
iW8Brtx5tlWrDPQWy3UtT+NgfMXkQvzle4gGwBZrv1fBmfeCFDfIQVmRK/b5au+2
TeXSOIOTh71/oEuWwTvyEqX4OOZPDMuOyy4I3EovDFs53JO0fqd2cYPw9PsAgjQB
ERSbroj87RBeAWwCc6Ji5TUmzERyj2RrjteMYIanZnbTOkJD//2SuQ9lVptXM5mi
JCa4gKNekbEUJ+UyiINn+ZDx7pzGYmcZ+dx/88P4rNC+u0wQQX7p+ZwEfDLT3vqy
SbFmX2fbv7EPK9PGKHoLKjgt1CD8bubUjZ3V+Kq89jbEeNmShNjJEmTiqfHW4Lsy
/qJqSLEjJrFtTMbNAOTcbnqMw8OqadipDTHiwtVPrFME4MB2tI1KaPTaideS3fLX
BPysPHnC6cZPaWCCGUv8vR3yq8tvspP8N1qCWpkUrtR0J3xBcr7XPR8M39dqMWnD
4UmORa+JK6ja63t5+La/mUwQLQRmbF0koiygTbrbQn+FGHOHWFZ+VbOtqjX8S8UD
jYpC2DjML2a7e6+ZW7B4zz2KcUXc2FzS1OM7X1B5Kg5ccNPWmS/sIY9WfEbedCu6
bGb0YgWB+Kacf6P/HBjbyQmcFPm3fAm4lvHe6EAGWYwF1kibssPx9wVLk5DtJ61+
4Wy4ozKB5NgM9MVlVor+nx3cdA7ARI3eVBXGgjtSV0JPxH5+UryiNT5PEa8nrhfw
bCPt01SD01vnongzru+/axHykzTKQjFrR4TXTwHVcxXIVj5ej4H66LIyuSLszj0L
DB+fNiY9GKiwiOmJQ1ezUANIQ4zWFoA55FIx38dzFQnxKXQh1kBESPwzBE2cFTie
HhttSeqr2JYaC4gBkvNc/IvhX8IJBVA/loGcXcyFwHlZCw5SE/1I/LYvu1uPpKAc
PoSCKKHBicTuoNTNVx3/PQHI98vdzFV87sbZ7d09+IUfPBtvaxxt3a6q1G8OLx/2
t6wcDeCOlmfJ/ziJVKDOSV1gtk4SIfyPWoLnQvxiMTJKmVF3sGmg3+oqUAFNxpDm
hbtYnFVpRKFPhCg0t/3jnhQ7BpGeQjYkWpmXNJgAXWWxdjhHMj8NbmaryqyXevq5
QQEnXeWd4xMl1oy1tf9CS7KY8cfZ5QSDvva9/fQ3QYecDMDU3yfshx8d3ywbYTJ5
jfAtpOxJFXgqhvHT3Ci9JDMs2H5tN3BLNsLzLow/w4IxxzSOUpZEUc29pJBXj6DU
KO+CjguS4h3bOOirk5F3bjo05SD+qE05eEIgn5XnRRaFyx/LBCoyfPuG64cXN3zn
/qiinE9kwJL1Va2RCztX5C6nB+HAJOJZEHuGxOzbvfyphqaQBpmxch+cZ+NHwECg
n5tE7M745Areua35FZ14Bc1iUc+ZmQjR7zKYBIcdz821qeHfA4KtLg5l5BuLacKe
EK+WoW7V/LubnhA4YsARQZV8r+rK/tHYIeQCLi6FQhJ6oxCGhirRWhx5ExxBijye
bv/wUQLiovl5DjZc3WX5ctEP/sapg04xGOQObXwUfR8am5hXxl7vOJVuPplafI7p
4lAzVyO4/Vlvt2VA5OfQN0leGL4csO+a45+UT6WX8vSxskgOq5+FWvw7LnwP58LA
Vw1GVUz2E6oIwezT+R9ILvAmwq1xQGfGltTYrjQlRuvd9pr5aqmH156iZBN9MMnO
pBkqnKANtORgh17XuzbDZJezY6OvQ43IIe+NrzFtykJN/3dTrOdSTtszjzq9h7Th
EI8ibhIbTwfvF6+lqslv7CnK9PoJXLZJRdyU81fHQqorYqX6CcbYhEQ55FUnnHq0
KMhk8K0PKcb/9gVNHW28GsegOL3aX86ffoGCRjVpLciE7pgr+Ij9Y0h1GuvEgK4q
qBuRXiZ8Yim8eycli40aXdYHiPdHJhaQbLBXM6hZXRjL7+3SvqTQMWmI7QzTRCJn
cIOF3PJVazMM+hnDktNwhC1CTXaf08lawjhcyTKwQGCQc0+JWZdfWS940x/OsDBG
XX7+KGPpG2LsXyBOSuj3b87cmZViFlQlnyRJRaw8lM8O+hJwDQC5d/jIs9hJGnKQ
aV5UBxxIf4PnbK9sQZbGhQsGeI7VtBYFcHaCJX54B/MprZyJR47IYtFSaXbomSZM
G92vVG4U36pWrLz2QLeGp8GQ1f07RRbWEcgjE0Lbe/g75UUTsdhpzovQnXOnREDc
1zNjw4nElMYwv3jUNkZmBzrz3Jj3P1aIwKnxsMqjE3SOXezEr28nlv0SVtbLWWCm
RttzmjmkR1ZIh5lbtBt6DvT+UmHjPb1sr9lXHGAB8a5YaCVeyhSs3UMsJErVxrxd
aznE83G/KMrmivZxp/BuW1IJJMElbsUyL73PO9ZNoKnFj7W6LUr1rmZ0Q2Ci6sG7
iz7PN3gtEjfE3hgfLj/E+Ug+XcAgX01naVzL6IoqZzHDuCi02xhher2dkwPx2ne/
2P2A9bwTJvA5EPPbgA74iknBA0T5zVwNdJAxIuHSmz/b0c8BsOJ3Sjz0N+BPGs1A
V18W+gi69StOXvJ5/AQzXVU89qWXRpUZyPYFAf8hh7yydZn0dgehN7A1ZHCmb8qD
20Ts3BHctAO2cRu+bE4xtC075CYwZjjDEBQLt0TXHju5JBu2O6f0Hz9YWhWmelh7
sPUZQ/Xfoqx5alPQ1WMQqO5sgVfsVpiiRwYFM8Fux2Abd+lSU2ZoZotoL+t+X+1R
FhHOeo6fKaHfIwvA3lkcZ9HNztj9MzChZ13fI/PcGjopk64BdCcbI6oAstlULNG7
QQyTRHDKybS1nTBsPk+V6AEyjQRbV+fVxl4p0hxEn3WGGZ+ZXHmJHEww7tmdCwH8
YfHVOI5jiRrfBjBYQT/XSVYI63+AjC3fPpTgKEHUVrhU6VvySfprPnIBTi4GXbwl
GMp62PLJRbWwjkBg3vScPvOYIabreVLIRIzqyuMeSGayValw8fEyJ0TjHGXhpX8w
ccLbPOR64p1SXIMehOY2TjH99cm3wjhNdMQUG+4MQESBO5F37VUDhF6Nc1C6anQX
ZKDA9SpUeLUE9SsaFwFgD+XvtoMJi86ark+6IBv2hs92XRywLrTN1ls1X0RZ+1W0
mD1IFd0gPHl5G/XUp+GNhFIuiFIvGJENSuKiTpu5xnHZ77lfhU4whRxqA53PaPue
QKcLOxczkl4WautN4vyuGWty2IPhjwvZaR9vWdtpvR2Hl+U1vNHXklPPJrI2ukf2
WYtisxRG4t9MGPhLEmkk3o51Y6K1b6YpOaH4Jk6Uloz4I4I8CZr1M965pjzlTOAK
ynupocZIEW7ZzvuX8nVT648Cd/ir2A78vpgqarTqeLJ/XI5ud2MwhBunBXPTHhcq
nhxteULImsaIpNFInp39jxEbPb8/+FxmXqFknzftu4PZq7GXqo6JFKiViw5nGPPV
nX9VV0q5JmL/By467PunAPWyHRlK+bNjzb1p8iiMYUGm/SXNNE5pPs30Ac2HPcya
rgKLA8kM56nfuDM9isf9NSttZILfYQp+W2kHY8rlACNipaTuQHjoUZ8Mzwzw69wK
0ydFyR84HgJZTclQKLL1dU2L6kgh9pCgztlG49acO/fsu1bk8R2GEiioeJ+tAbPN
pkKP3ByBDYk40pmhypPVHtNU7OIwttA5kXHeROnqivBmvr3Ct4VqrQyXWGRn2wr+
GwkFW2O3sarvdJXHq4aYClrjglcgBsZWDPBEdOC5V6wt5qPrRKQTAMQbCaNo0eep
sP5gAfwedUbgwDcpO7Uq8oahJddGGiul/t4uFX9DqBta0gRps0g119s1/0mePcBx
aCETYDe97xpNcoHR+hwh9JOLEQCkVsRTQL2F50l1y8s+hXj2G9qu2A/K8exNr4R7
dPQTxHLI1KYT/Yme9NPQ1dw0qx2yg859Sh3Wf3guFKz+fNCqUrNVT/N9KadEzhm4
RHvEiIfqY+kvtQmhpHud32cAARTkvgbOEZQybQ0MU+EgYa2i/ySQ0ghIlLsI+J4n
iwTIWqCAFNSjCda8gFqMsKt3ZEQkVB8J3bdLDBjifIfMThRvHc7ThhJYKBo0zwPN
Wmx7NMuU47L2gATf1/n8eO2OiUbCkTb15MVutWwbcx0N/C4hVvPhSw1+kJdWctTf
zLqQbtUjQA/oc1M6fqR9wOMGyDZWyi3MYpuMmAKejgiAX+EFqm5B/eRjevV6ZR0c
qiuGBPWQDbmsnWxuo2RzADbsfG6S2ONW5qtD+Zlq/QKfByM1V/ijgHzYCEEmmpji
sjllCfYx4pPNoN/sYyxfjuD/HjMHhtDEL2pTku8llhgdvaUiUXWpjN05Wdlmmvn/
iGuBmiUvAOB6xkqq8m7So1Hq1FJRbZAVG3diEPS1wnT4Bcn3m9BO2EiqpikA/myP
CLKQWnJjFFUAat8a9wq8vET6WFTHV/Hqebcy5HP3g+Tl9zhfnLiHQPlW/IP1Dp38
l+e70cZbPZ788D3GMME6cANHDeYp4qU9xe/ZkFvgmPtXaBSblneJmUOqDmWS0sx+
nZVBqLHCtaNEFV953Xjn02A0xxYQHQ6E84RKF2u4uogzilUSO02OD6WnU11O1t4s
pnZK9JBsG61InfSTU6KNTeeSXAD+s5R21Uu7U2Bn017/nVPla8HtxBzazUoqEhcm
MNOME9zR5IFGpg8TxKakYFh9Qref/lijU6FrVNUsZ8YmC3VFZblGfsmyn8BxJU6y
rOW6BsLYQCenMT37Cj6qU0OhX392Acs+Tph9vKAu7bj/zZQBM2+5evXspLjku/93
GFVD3XGrcp5P6YT/Gt/Z0a4TPu1mj4uF3BiYvHJp2fLXF6pGFfRkCF6RR6cc5iFP
jdATcB5BpCWgfv5LW8cBGxgfLcsI9cauuD+7meqJLvD+m4AWw3oV9LsuHWHslGoK
9csJeyqIAfn4qlRX2KqPioWql0ZItBapvEANLog5WdAobzM9NHy9DhviwZ8wcUP7
4TLpkYDQ9UGSg4GAmDI5IIic4RkHrX8uVvpuxzHB7ufQxQ865QM7HvGJFM1B46Kj
WHN2NeaC0lTncxPO8UoS/KU6npKSqWPzagGb9ULpUZIVOtlqTdiLPS7W6UQFtiL3
cTNokIZUm9dO9jDO/iwoKtrHQ3BE2XcMFUeRvX/iLIVND993Z/KyQHl0BD/JXFsl
ptoiQ+sAvZSA16+BZ7aPcJhG5YCqCrBPJHKAFe8AE5WgG8HIS76ABd4FElPiS2uV
j4YTvS9K4l3WfuJGVz0r1Sdo4BJ0j8o+0pmNlJSMjj5UuyIKllaA0e43aHfBdvZs
rV6y97fFCSMOQm8wRVyU0mdUnO4GC3WsgJll62oVhCLxHaQaGdQ6HNEQ9+3+V1XS
FPfZaAGgeGppd4MyN+f2Z9FpCZ0x9ztvBOiP2P0Pqe+qlLb4vvyY9/1o9xlyzkn1
dT2u15JhKGD7b1sMBIJ0zOdiwDRy8cpn3nUGOgMWzK2ZLdDqUVBSmPdjpj7e4Uvl
r3a4D25d6p4TWfTgzZQq+hLJmIrVrqzJ8VKt4LELCXRzIx3LwUTb19gALnMp6TOg
XOx1l7WNklST7nqMaFf2PZZ/P8Jn69ZiPn6GiC5SLd9WtSSJH5/UVZm9Pi59lBwm
nHAg0eMAR8UhA5T1HQ7nk5mfvT9wnZPlH1xe3JgbnPSssTmrEhN0LTHrwQfgQGlj
WDHJfFLorxrKWNq93dc58YbWATpTCVHWbicYHe/PeFo5dyAvbtnrFYZ+jlA3brGK
xoIJpBMKGC3q8Gfmv6ROf2T4UhwkZvZlBpblK2W1Mc4cKwLhf3FlbQ0xZmc5yYRJ
ptSnKD2CrDBGgQtvRSmlciAGgJco//2t+DLmCpGpV4VW1WR+4FV2nn+nKCjHTgnm
1MGCyZT+GhhQ4iQ7Ho1s51awO9qu0ccI/XWBls86JIw2psfgkTUOAjUpLfnOp1qi
e4OkJxLqKY9IvJx3ejiqGjxR0kDqG/tqA+HVRBggY+7TZ+i3t1LCouH9LMVnLhkK
r4wn0lFBm5BcIJb49B6dGBTzPPS2mnPq5KfdAXk/KPFqI6PiFKKjVABJAqba8L0V
TdnEm5z9rXfHDG65b28fRcSeeTf6iqW3qviPCjvxSFAkldTRETogPcRKHqnYFCxv
xcsM8jyLBrsCiI+cvPWCS9+IvgEgx5/0Y+XO1/hhPtpIUzMSDYqgaI5QRrwGNuxy
5KrJkPyXNVhalnZsXXOCWUH2R7uoPTR6mMLSV2Xl2P+9WAI4dENdyjcLAnuNjVAS
axU2t/mDmJC+5J5/8PGdklAVYvPO3MJynbRkwHO88tP9rGjv9SEgqrwPQxVsV6r4
zYalOgQ52o3TdHpHGmWQriESkAWwqTnirb6z5zeDxWoXk5KD/VNDMYALd6bdkET+
OVj9uW2N1fhYl2xHz8wvKpx+6FK7NtO0STHEY5e8WssHEk5LvoqeBtGA8MSEZ4Qb
55O7Bb+y2PmnP3tLtetx/zyKBBvHjbSzRpxAzJeTsLBgjM6zzsknUPcmwHNf4CAa
Ce/ZCbdYMUpG2rudfSia0gkkg6yuG55bcuCPLRM1ulF+VX8tJUPVIGQgceUyqggc
p0njETb4RfXk16se+D34lUuLgOMzpqFKbo6NqVpsg0aSw3m9M8u2UzVfPXHvF0iJ
dtD4gqTBN6xrA3D0TMXsnEx1A2U9JSO3q6UfzdICzzKO6HcLoWewGbdVNQyj5tCa
xbrf7H/6fxkYYo3gXwA4G6Z5iwQKWiu3ci08eoCXXdWXjAk4nK5Nt9wqB6ZfrnzF
kpQEQaPu7JKTiY+r+u5tgBRYXIJmUH53x/33Mb42W2542qQ/Tdd9UI+DNmJZVkmJ
KFsHjHSHiiaqjb2MqNMXvXBJyhQCq6b6NkXbY5XNX8PwGcJ0G6b5EazzOx1PssrJ
3+i5kwK/bIvsXjtujcwg3q4nzHX1/HW16DFGlJw1xyyOs4BiQVd+lUMOp0zJb4PF
rjRwBhYk44eOAsaUxa1WMANgb81oXnFm4QHzR34YgBdM/q+8/nHTTMpAYQxIovfw
Ou2+Hz6jrSTXSL1+qm6MWgVVNLyVfo7Xwk3UyByFtSbom77a7WV6T+M6U9ZHy04N
Uk0p7lufy+iXWKKi+MDnDnIn1YEHp8KXY9ig4tB8MncK5OuIA647leMjnVQ0Kp5T
jb4ewCd/e6ARRrUxwgBPj1ZbtrP6ZtEiyy+8fIPHEUNF/i4Z3smaEKMH3N53rejc
v+3EvYfzkT6CYEvh31DjopRhJY40V+RlPtiS/6DcuAnE/duT2PGJTuwe8X2YC6vp
FsrjDeXkiNmz+c/VuGJ2SM/0znfKYC7OXyJLH9aRBNEAl+1wIMge9bQpOZMTyOzs
Pd3/R1amr4SFTnQC/PyNOd3ASJEtSqjzOGu8R+mnmE+UkGn3LAOVSt0hDCuIclMp
dEGZRic9JKcDyhZB1BxPRfPl/lcpAD7C9WApZ6BEh7r44l7PhglK44kQvLzoRNcM
eFJzl99SgmKy1hk4GXzex/SJimoumbX2s/wvMUYrvapTbVOWItd0zoKzuqcgCqcy
wBdba/cS/NwsuMY7KpeDX40eIl3QI1NoolMkPnbQaQt0zBqQJA/BuIlp153G1js8
w5MasiTNhKBowuff6NyE/+vDVCpqZuBQHjy/sNoXrcxjcrmtGn/JPHVpP55mTwJC
Qj9J4DQ9e0nRINOmTejLjGGO+E/S79E0n/57uDVadeQG1aJvvVj9rhSSVtHNF77r
qrf6+UiSwRZQ7UnQnecUBs50Cb94gleygUecAJ7lUJjBu2B7wpUjG/rI1zTsaFMM
Ngf8K06XZ3Fnxks3d/qbUOgIamgoEQ3USiefWtD2sdFIZehMSz43cwxe8jPeP7/s
i0KYXUV3vZtLLSkvBtALK1cKixF276qxUcrsDLvYIv3JVmMEc1LkWkNl8OJmAZcE
16dRdcY45MpZ04KxXxfVKBJGn3+jyv0wyflO1SWxdbEoIFGmzBkmWXOOWRwekZyR
N3B/qpFK/FqHqEVFXMk1yYL82QEFCkItzvJV3OrzXPcJE5xstown8IwOo71ltTgd
SwazaF9p+APxBCagWYEhckyGAZ3Bnj5sa01ZGBnr/3JH7Pjg6qr/JUOJFEte1uuP
Hc8/sHqfzI6BERJk0Koo0UCt68U7i5rpUOyyavlZHF+ttUqyGBg7SunyGviDuj2F
1W6iC0XufjynSnGTTB522CJcX5b4PBFbr/AHVEGu8J1OUQnYOwOqMhjFFwVRFZXX
dbksQWdhvhLd6hJVzteIqrL9s5sKavnS3ItRVNBWcl+vxyJj5/EC5BcO62rGRpJu
yc7/BThSqSUxoAgF8bHTOt+ozg0VD4BZFcD7fPfMiINbdPp7aWR4PhsoyDwvluf5
iIGXKNCnyiJSwHwFZPbkFuujAorVHLtUhp3KPjZEP2jkTQJ7sUIA2jg1OK7LqRxx
d7c/D8MVUifeibKAKhNQYHv+OLCa+8BsOv0Q8/dRFjD8xN5W3FGelUGevxb+rB1o
ZrCmTr1VnKY5hvXv1W35QLjXd9/LlF1TmCfBwcoNMk7AzIofkfdMQ9md/bNFedvM
ZahsuSj+SBiI49nOViJI8yla09ERjaVwxwY0U1QMSpyc4DWXOFku1vwKG8mEVnkF
WaDZg3QmsdFpy/uAAGc2K6PZRyU5ku64nm3PGLEGv8HF52SkkONBXHq3d9kXvNBZ
VPs4Hs5AUqxdwKp5EFQw97lxW3wDa3uwGc9gcyMGIzN9yypkkrTIGr0nprld4ZN3
6cs5YCKhDMBg6JUNZxQWks2TU+6VCln2r5f9iGTA74zGCiQrCX4pQgoOyER7v/4t
zOBpimBN9Q143CguvZcJEPL0Z6v+LuN6AhwYahE+8QfwQKJJDbJe1zOVywRC6cCZ
o7uFpIMDyCS2mc4wDT8WQebYqYSbYfGajwIbnUIuZhxvRLf0B4FOg0PNNmXaHcc3
z2hwkSGZ5nHSBV9D1TQEr3tugF7gZj87D2fLL7VWVxvs/Pel5ruV6fk0tsG74ppS
D5XpcFCtbBCQPkeT4m6BGbytGC7zRdVCCJYfuAK31bHNkAMttY+lGex5ilnycQLF
//qaIiD5WOIXB7FFAYpz/uFKcAlOgX1WkvDljlrfWq3R2jQqHm9x7dEbjwZAgOU0
3WTvkLBKJ5j4WHPCGcaBUGCNCEOPYbSZYt4+w16LuIyz4/Y6meBIWAKE4zzHYCBV
7gumxLp/XF2ckzpFtLi5asSphSiFoEXUS9EJzddoPzN1Ft7rkSBdejpk1cMVwL4c
/gSJF7c+z8MZ8DiGK/cVXK4LTCyrhAkaTUz3WiAS/MuNjd7Xk/ULU1LqMNXm8NW1
QOodzSEz5tS8S9qXafCcriBSfZwLnMNc1kmeEb3HdaEVPRwfPRgtyYuDfU4IjQR/
x3myQ5RzE96AEJki4l3BZUvxZN1JZ9Ko/9F0BIvOUNmrHCVyJ53vFq1cf1oSOnWZ
bfxIepnoljKBEsgX1l4JMeUlIBj6GO/QkL5lFhcpr8XDqruwLLMTjorb6zepPZ0i
T9xJE9ZN2VzGiHjsEDMLeZZPpXQVsd7pJnbPWT249MGkNOGJiUeENFNxq1NkheiP
7OFOFdQqonOSRWhBLyZ17EvSiVyYnoxqhWVeQ8JgbjHNzuLEH9NmAgoTjxnqZhPE
VxoxlcaKcjMUNbZtxNfuZJzL7Kk5lC1fmdX7N2+andeZheOza64FPxmuFtzT6PK5
/dJ8EdCsSiui3Yk7PE2GQrabvw2csCm65cxcde6ymqvExsj2K1ollzsZpUUqkkdG
JXg3/20h8LU057SY7pemfOtPBiwXk4LklVUO3UKoJsOSTDXuDMObJX111qvIdEav
pyrKnxuO1LyVDA9EGpn85h1WhsDVxlzCXqFeZYInQh6b9mrS5jahOFi+sMvrbN5h
Nk7+F79lmeNdLodISFCsyJJmg8464INgqZhbQ8Tgc5d+2KqOrSu58Q0RhOBNJlMR
AKlWjfHsH1vh7qvEYq5Ajb/DCMW5oIoa668P/wJBodzQxZCMPS2dqopB3xNVbqgq
Q+Fe1nFvS83bk6mFlkGMHadgNxXy6N5uF0BEy4VeNvuGt567c/qo6EsYYya/Zb/i
Bx26GClt7Q1MwJQCdHfuKBidDopayL5w0I1eBXDnWCuF+T19AHWw4JMCwfcyZU6k
iywXY6hw/z8YrqFxYOXd+1t9XO+1x9l57FwZOwuWtfmzereyvHo7KovSNG4yzJe1
upDWwEJOJQ3k7tVfZ1RQyoyqS1C+Rd4UU9N+Ya9ukYriROGUSAKD8d3vR+rDmy1U
aNrwy1/eVKxb7und6IkEXHwN98IuWCDzJKElijXhQ4tRwhPfiMwxKY4aELYSgPDl
Pco0leLZjC9Hhmu1r/htBhz7Rm1UQQBmccJ8b4yEI83kW/QPtWwC1z4YBrnCnp1C
KFdzPu9RFHqqrKCzm9b9iAjGZ/3JJR5MywdCqZs9U1Iy3gN7RUxSZC0GdUo8orva
ddm6RwcSmNBfuMu4m4VRzpu8e05HzqDS3gfehVxBVLeDS0e5J3jt1PiHMtrdHCnV
v2Hh8BhtjQfRaCnr4RV7SBTHBmUhb+Hlxqhd0vL1Ss54o2h4h485D9wnZuaLr4xK
PPYmNK0QA0CUqWxK3zLyq9RN5gRRsBS86DzGH9hGiooNu/qoYRs6+g86dqcQBIRK
XKAC3Fu74EmzN4ntXsTyOxZCsHItNWDrKP1JQ+y/bptXRISVHh7/Bmsa7AK0xq6i
VqUb8ASFfuwnX+XFpK5I81GT5bAYUiIKaDkph2cjm7YszferGxw8MkxLsJANkxR6
rHVRbQQb70dJ79GpV/7TwagRl79WBmwVs5CsdgFvsrCElfq1+XO5g19+t5GnSBPD
aTkh8Wf+0q4gZuuQjtuxMGGiTMygv72Lp2atBmGnOubCbVNsi6roCgfbkSYCf6f5
ZtCZBsx7tUY7F7e0Tb7M/vHflW3Xdfg4s5/YNbREGS+oFmw9D+RJjq0Biyvc13LT
sRLVfyR2oOhUv3EkRzO0j65IXfcUirP0VwfYj4+mnvyet4eVgJlJR8kkYlZ/AK3E
W9NHvC5yF1M7/Bhey1EENBzl5KiLVvj6NatL5GmZP3T6VIBUft+itVCleV2fawcc
D4fj/LSQBaFE/rG+7EShZnELKfVawbB8J7Jc/ceiUEmdZ1c+CerwzUFvoeiQNAxj
UqYWqAMkHIIDr1uSTAQ8z7qiDQXt/kfTGdRUmlvWMJs72gm8w4gigDIf62EqTksq
/CXp/0k6E82Cwcory3Rfun/ct3XVVETp4ER5HLxYaKz7CYKgs1YURJs9pgoFjLYr
VFMUMh+AKz3qy5SkYUY/v9NN/j8y+CYrvUNgPEC5b3mqea7BuAbFjZMfGiQl26/l
Esuhc9MLwYog7qC3l0H2grOXlW17acVQbS3ISOFJGFze/e2NdyYXfhoxjPkgBqeO
Qfok/OrgU8706WuVBWvGXZeGFWl5aFGlr43vBLmGVrVHdiLVaNH6DFxezEOQfU+a
V9vRYM2S3tdE9MWFLHtydti4ElLhjvz29NHsPWJicZGQWfwCwlZJbXkAwRiYAudu
AaN08/yJUYN7uXkB93q553Nl8HtliC4yaVVazGKv5K1OQ50rAzviDE1fqtRHyqja
vabvlcBiJ2O9jeyouCMnxbMI8IGmslrlcwsF8ei44NkZ9v8qdlbtDQ2FCXAn6odC
SC67KO/fpHRvhQugq0slF2FSDZn8J+1lrn7Yb5oVeZea0kqxRKlrAH7A/oFhXlWr
hAGTgYUumNNiCGOk9Q1obmazojLmAzTh2vdwZNgAXW9YhwkQBCdiUB28o6/tTuXM
2IMrf0r4ZoPvUJaWjf+uGjecT6Ufx8yDYwryBU6DYHb6y39HuVwQtoScdTXDTgJR
VDO2a6En3kk1KKM82wk8CKt4ysfcIE87hxdDtXnUb1UMy2S5+4eiEAF16GVMPQhH
aL0MsxjPde9eLkoHdP9i+x80364L9sddOrZOgbV0ipeOvx01PQOqQPClUYnH1akx
gTbAKj0EeHe8DQfE86YmM9QbYCYa7Uv3Q9aVGcIwN4/W9qG0dHSZpgbbjr+kt9iv
DjuGSIcbJQ6htA2AWX56KjfKZ2c5sgIK4mVPWLpK9vKX7j9MSLoWK4Rsd2uzC2Vs
uqjqHAy2qRUr62Us5f+WNtkGCP07Sw+aouE5g5wrp/Tj2xVnw5dzj3+PoEbvc5uP
6cY+ij5dU08ESoflotdeN5REYrCPYZj8unPTuSMICjtynd8Lkte8Tb3CSLlqQ7Uw
vTUwD6ILMknrGe5mzeAqFX87/Clfe5I/8bjJQWcTUG/ZJpUqnKiFGzWCjwjTfYV4
7dtGmNbeCb6ADAPsRsWSjehNjzSeVo010VrXL9mn3+B8ceecfqVPpshiTlgrothE
+3lW0Z8f7k4M6PJJRvJZY+YmOzOl4ZIcqJA80wXpTWZZwrHjk8OTpGKMRyqb5Tul
71V/Q+ieaWZKKu4c+SrFVihqfADCsw822d/wcbD9oG584SHWtNd/cbfbALGnVSHa
kDxH7evRTguSkqeP3xj/FWW3L8draBCOBcot7zzo5zAWuudURldohTfAdEuN5k07
cxrHw/ezPKK2zOuhdLS8IksC0ESyNY5taEBRU6QN6hhYc6AsdvVyi0ZATdKrua5R
eUHU8afRuoFo12nZ52UMncx/TqDbwE8pqoFTMMTW4d2iPykOoWyh0fGoHvv+5g1p
x+Rg+okFnGg9rhlihmQoJWIaZZ+YK3UTHX1UuqCT3Y3c70w+gZN5j7bt34iNmRX2
afJ+ZNybuJssJ/JpduwjjdJRCfsGwCMYCn0s7u6czcPehfjEilguc8XR5kkIhVmO
HaazWmX2HAF2e8C/8P0/POapLW/I/qsq3XHRRvSkxc3cSEnIYq6EHhWxoQXdbQlE
86nW1u/PRYNW9g2fUcnt9/8c2eAGb6tmHhA5gRcJawArZdSu59MLJ6HcEsUiMWuK
ik/TKQz/q56/wOcDCT7epTsvWgvk9EEDQT2AdJSYevnAxYoqpI6NOR2nHYp6HCE3
nSCjs62vP1rWmn+XyjF51vJUlshm37LwjlOVhqWQq3a472LPR4M+t7Q6//kQZBiH
liKRtlWl/VRc1HI7en2FXpgpFJH7QfukrOQzhlDt/AzSCvQd3zuRj9thrVkk6J8u
++K7+k7yG0f6jAPw9tf3s8fEGH4k4ZS9V6QAGWEhUTRPpX37XyJQ/Hdzxija5jvV
EwZCjbTd7FVp6ET6+6tiUimAM97YOWXEayrQAJJkNqZiKufRm0ntLqIhEiaF0dlq
N1bW/tYjlaTIFuJqh539AU60o/jk+CwWOkTTA92l/Q3PS48LOFSqTFUBCdOshZCm
RpFl0k9Jv9fCxWxFhEGIN2MtrCwzXU74g4G2W8lYKCHkdlK3CG+fTFBJ46iQcr+Q
tbeD4kOXNqmqpbS6WIdVl44mBxJfPLXCCN2zqQamk+CLkQLquUWNBmwZcU0kA922
USs5zkz40PqRKCY4XACfwFYKGcT9Z6/4MGgBpWzofabNjYv+yYy9ieN2eA4QDfke
3/QBNC1Ix0OgjjqNOs7gGf3fQuWVTTs25BLOPsb+i4InyoG1JgHf36PFixZVuy44
qU8gUmNhe0VFQ2ffKt1qM/XYDx8uyvKVbIdwfo0GJFeWhqUkuitA8FRv1jvuk7SU
cdbtHJuAQo8mQYN0mLiHwNq3kk+bAamNRJw9VCtgWGstl7hpk/8+dqMVwsA9so+a
LPuTk+XylpJwwQ+N72YbnyKTLfPhGg1Pj1jkz1BJXpnGUT6NvxTPCE+l6sHfulxj
5TVwyVljtRe/XX3+rfEyg0BVgIdEhtHD5ub9nw9S23iNlcA8Apwh0nMBBudZMHwF
62no3tbucJv6AjXDoEpLuO7wfGYYYawvdUmVS6EKDBrz2oKygKtbd2PpilBjaiuO
fKKCqyr97SIMkfyp46fuxlM8OoXjhR8F9vgtHQI7KtnBWi/jAEvcVN6w1rzRybju
CwuX+tMk2Zhtxed8ycPPHmAG5QYeZXTOqOwptXQotom4HibzsZRzm6fmDl+5dugw
m5l6xgzsscblKVVDOn9gfjXGczoWpPBbLJcnM1jNp5Q45ysLLYFqPGOKSd0yrvQc
pIKjb245xyZei6uiixWk8xVg8fUwktHxuAb7vJNRPA/SwyKESeTDpXz/zWNpt0jH
MkI73oRwdB7NHOtmLTLQg2hlwivYErbIqvffF5q55KWVyoRUJxdHaER4YORtG1cI
Duh3y7OhLEM3BGL73gJBy2gD/t8acgGdf+ig22fJsB6cU++rqaI9oXKAa3xlHeA3
5f3+P5utSECwlpmhwIEZ5yRWhx5kp9KHY01UeT0d8aA/MUD0YRJuVKTjsxJTaaa+
W5cJZs+/XHfhb5Hx6VL4bV8lJUhFWbga2xLVWX0P9BpaM1YjVFN6pVvd01wkSrn1
mCLrThaPPdTMXivMhSR36UHqxbSZ9VJtjru+mLcs5IFxDkBCByNAbU5al6rvBDuT
3YsCy/dLJoedcQkhdKCiPja5m67HbKVsGVsan2mJuKiqzDMryxyFhI4qsHm9mWZl
7Y3gn8RpkxwaY7jLdvc7jL3HMghF1ApS1C+vL09j1ALM6iMV/MtM5SIuySf+1OwO
R5avUhNqFArTKahxWdefVhy36yVxTYehKQpZQFJXVFB1ZzxAlPGAnXY8gAphm15h
32s4myIWoT94JP1NrijkG5ACYXlLMAlccCZt3OM74TFgjNPbvFejrqqyLCG54ntB
jK/0bQrdsyWirq7VHT9GX+Dgv2/18/ruwDJ9FCcvVn4Noem11m7i/9ngEmQ3aFM6
pBupn+eR/k4u4ut/moCqvse7oSIxK/9l9M56jIRFas6y68jlbajPVP+8/v0K9hSX
JZjio1NN79BmiWR5Strtiw5HdfsgWnMbpHFWvixXJtzlsbstOmARES8qzYZm5hBy
w53k0+h07GjdJuyF4lXCGKoLGCvGK+ps4czmq37lhwCOX4UPMOjN4IOsa6bke4uC
Wy5xsROklY7qt24aTSk933UVhKo3gNjNLbGQ4+dNJb81/D0pD2AK9FSvq6w5QqpA
H0+mOKEYMfLI0BY6NeyU8ODQXNAZeCrXaVf2iyBiPGchYWycfa+Z8KUTqIkn6pin
DibHGQyZf4HtyODOD7iUbLsRbo52VtKEytIFb0CdoJmbVmnVTiRVAhktFuEZox3y
tOdOHPfh9aRbTCQJQDx1pG2PzMyo4coMeYCOfM+SKNnXlRoeP2xrMaPt697VGJWw
C/XTm06S0b0Btj8xUd/PRJm1zTXRYcqkZZsIWiPUiB8GOZCxbT0GxzKtekjGOd7X
H492lZeV+D5ZopmnNbe/57kv2frTuCsBOb7FKD3d1L2OhZgvY+wGbywv39ROu3qx
XSr2fMjcWjNIkER2I4xWl2TjUraxHOKdluB4oQ6BI/1hY9he+GId9VpweufbmQIx
IjeZDYyS4WGuaqgd1gGd8WZV75iaqXX2gtlnMBug3CVOC/v2/meIYR9mRMjtcikH
QZMMNSOXsBy/Ad4LOcRA5fbvblhqWtpTjnBXriB4HSv/4ANM1NXQ+yo/3xvs3EJW
v7PPBM9jbDfhAIcZlTA7xEw9i35UVPmn/O2MKtA+IS5ldl7hZBIOsfwQj3vF6TAm
tar0jtqX4wEuGk5nMM03UBM97ImO6UMPwRqcVa2dDzDTmBEMjXmdwj7MFB7pYC8b
PQkMhqGtBqLAnaKo9Yqhwt+D/Vjee6UOHZ4umINyEbotCC2HQ763FcTgsvvot+5c
CNn2A6yw7XG2/CuqTGuPWFpyioF35dJitqKilUrB2Cu0ZUYAL7SAXj9geo/9kfx3
Q+ChGqFoYg4Gurv0bX7+GJDb4qMfVwnp8qaoZlNKqu7mjDgM9obfzQwxAb/cCqe9
BR6V2u0qK9FGif8kl++9DPA3FeZzt55KNH6BsFTURxW+3j/iZheTlbdly5nSV8af
9aldM6TMp4PgpFusP9DSUEzlyORX6VyoM6tWw35NGIktYZoRCoLITTeIgXEHcwIm
wBmErsIW6hCxICGeDudXWutU2xV846Zr6j9QgqQ4+cFOJE6Sao/6VJUIIDVJzZzE
BMivMH2XhwXILioDR6Mstu3QbSSUAJNLdV0IMgcAKsVcdhG9hqXcMXR0AiMmoCQc
E9xYokViG8/kUEsTKmBxkOJbfDdL8DNVzyy9qbv8a/deJlfZs0Zp/uIE4CXZKDAx
ksLXIWGnAyXbZnN+LOz8TGqeA9n/fm/4Uj+vz/IYoinn52BFa1wJ1mx9b45ucpAW
nun/1bSrGHP/LYKEUevIKUDHInkLJJov9twnPTSsjEhtPtL0qmu7/YlQPrYIIsfZ
+hYW0CcVCMZe7OmZtMBF8lCNNyjwhk1wn47BSQqZA4nn3H2wkGDhf11oKNiPkSwP
X1KWxJg8+hcBSvoHwqLZcLZi/W+bjbTSnlRAzk6LT9sFs5MSVpQMQ/w9TZpJQNbS
vv29oz7tXa3ypq1YWRLoxtEtnDh+tKCT0sGQazM08FIsjrc3SzrO5CW+bqE/a8KL
NlJGLz0/MwP/KEyQeRZr8UPRxuRfBw9/xXksLaEs4TiQEIdiQCL6E41AFq8U4d1D
f7jsvGiTLIqiIwb8IPhMfzDqEyD+fQWr4PClRtB/BZR0RfTQMEiqp7UbC49cE4h7
QRJrWZ77QELtTAXH1VUX5hqZ+sHCmH87w5qPUhs4z1tgbeL8LBfd8o7aqIqHKj5l
6dbCh5AYsvvsQ3clpOHDpH1S+u5oxAXW72uGYd5tHQNMrBfA9OrZ92Ed14YrM9Hu
K9onXWRDqhQjNC7MOgG9BXj0T3ydITBU3wLPGLVP9z0+/FFkgMMFzybHvAFEDD73
cnLFog13X+nSGNHwtqbslFiqEqUiBEK+dHM4Pr5X6LlomV1pNyetswUtDyNZRDnI
NT3C7K8D7NpCiXBQM8jvfUgPCf50t1eQSQq3BQW6WY/PB1ZbVCpdrlAg8Ct5FBS5
h2LRKSKQQIk1c5C1m1LUMpLT9TXhTy5gn9rasfaEz8F/Cgi/YDFiBuNkru4mxFos
dNmqyoiMFJpRXYpFoUlMXj5B1Qgl0pYDS8FuBT59OYm9I+EclF09YUJ+7QJqJLUv
KVgJ+8Ms9VJ2gzLEaCgtJcWBbUy7PiOQ05FgznxqxawNWLeOsN++OQ3KNjkBL9HG
dZSjenDb7POm2opKEFf1QODFQ0hC/OFJMDS6VhGMKyok3NuDjSViEPcZrTJ3MBEf
l/abLDSXjsQKbV2fhtHpEmsYy0oLU7mnbSBhWcwmJAUYKXHfDleU/9gAoFIAd3SD
g7p7Us9l0623a4l6vsw+cULZOsv06gNL4LtVc6ozG8NZORhWPfNz+2roRF/+B9JY
EpjG0uS8GhP81UX0A49B9wVDcUESxtxbTKkFTZY6OMbEdpQhMOfKNsTirs5aflTQ
uy0WdX/9PYp+4YgKqEwlc+zKx60Blvr5gVfpKuVKGdTTwPOCFhBAWCjkgbKx99wc
2WmwCDgXzOwPHCF8plpvYYlACQ1XCFfPL7wvY7t0VdmDosGrd5p7RQU1JcukkFBe
RO1WV4xBVMRRJRJXvGSvVQ9WHGJKHTUivWv4WDARybowqXMJomlCvFAjmQcQlven
Ajvv4kK+tjdDEucyGZaio+GZhuqmabczBksH/497tyhmflNY0k/SRX+lc3cZ0RJj
Ttr6TfaJj93gwEz2CztdcEIL8scp2QN54XtB1H+0IY5MXuozkiQ7mXp5u9BgP4Cx
oCCpo32bEFSMzjOmShRcvyKAAcKPNc1x5XJPpaL3BDxXIrtRQtXgIH9gjmIOOAa8
48u2va2w8WsMM4RwKirh+SbvjYeX6Zg+eLUcbBM/ECL48AS3cCAPUVlwpWM8OwG1
64QeSGi0AKB9gIQlJP9FEizssiq+O+UmT1CFHJazswXsQyNF0ZhRxysshJ0dV9ww
4Hzp7amuisDjX/5qO6xBlZTgYgfKZ3H1en2sQKwDuIToFoFUZjQMqCALzmRAKt/i
/CVM13tJR1ei40dx2gtmuATkwTVe1FbNZ0FU4badT+2ZOXQ6LlzZOfL38NAkI9sR
iQUI2w+T78XGSVT6yxzFzh58Pbs6LEdbNjIfcowYkjX/gP+rY6DneUhTLtw15FCA
EocplrfKqCOFtliMZgJyYV6IxZjEqExvypduQzjRJilVHDTtnUFr0v0wfp3R5U+l
wYAXIuIm5IO1PgWI9NeYStTGi6bVKg8bcj+Mz4NFKJovdoma2bO64QW0MD7l/W9I
g5S4hVa4r3VcKecIkznDEp9jt323NE521xEt7pODac/sGrHN9Ml46cSsi3I/ZTz8
gn0ZytxHGA436eAHXO4gy4HIrG2r3jdT63zwrxPpvz0Ta3pHS+Q2tukj3LohJrEM
bqTgc2KJrBY0pi7cy64Qk0TBaDUuBlQSlIcPlVe6YT5Kg1FonU1d78+jYRUYvvS/
q1rFoBKkM+m+wbQr94xAovV3L0aSkzdWZInnziEX2SvRx8x1whQ8wYQv+PZGjRaB
AEZQDu4XmDn8WHmo6EwUy9V8iHXg1V/ZbG+NsTHvE2Y6UfOt3Bauv7Y/IBM1wOWn
YlOS0beaERnf2V8BBxqXEvVC3oopbgLwvVX9+AzN4Ggwh8phlj8daLv07W5QPNJ6
MPp0gVrmhzo/fbYeDUfYYjDJIqQuc2KfkG8aVgQnULKJAWJNjZeeiUWtgko9LYJN
HRNQgrNes93K/81Y1lJ2NrnDoulZtcTOc/UlG4ZNvPXybj0910S7UkJj65cbejqB
8Ugdz7NwOemnrnBEKWKzQaMeoVrdZBJTdgm2nHHcHOzoR1PCXKURwftE4+dQZ4pC
lh4T+nSfiUt3H4nnZ5e5HrbFF9Gkr2Djf+PqYYjDFk9kDS8ItKXyxY2zx80omGNL
L2Nqp4DWRZYseDIa4KCkIxJmuSM76E+66+nPxU6XbVc/P3XYNhLev2xyfE8J16mP
umNPLcoA/H2+bKgc9fUD6sVqYxFNaQ7vqpjUr9y1XVeO+tQSR9dyh4CQAttiHH+O
91idmWOzh4OEJd2QvW0vwiLdfOE4IrppVPYDN/5eDdgeczjJo7oSGnZi5X5gMrDd
5XeqVDpdICkIjavxmfOX2NLjkp8zGIwUZGCRugs3A3HJuOwT+SMRMoaoZq78fp0i
tAh/0TXRtYeS6D3w9+3p1wLARRUfr+Nn76EaLD9L5T/7RDmnYQcl0YCvRnnycHm7
HN0kYRYVRNJ5YSZYpq/pJR+3hoGRF/lF8+TimyETxpnBzeJ2Ae7L3xQTL3aG9+48
S2wGCu3g45WE6GURKoMy7V8fO7hIWedJNM0J47L4dW7YL3XpNNGqS1sl/Bra3gco
zNkWOMmoW/4YGeQWIP0oxPG2QyXEexHNu3D4NlO5FUGpR1h4gIoj493ln46FW8x/
MWriVjV9I2epAOIeVLDKh7tQHAM2yN8bH8yjJrEpHRdrf50BADIiFXGgpMY1pmpK
hNj8T++PA2i3bCmhlU+K+qdYoI/znNohVMfmjNYof53k0I90k/II2fjnSWsTfEuo
LWYXTM+Z1PrzSz43HNOWz32wRCJ8FNrQemVAmu9z91UezaeEgh9PTG5DKuJPlome
W2azu7eeXOxBwiq6D2rZ88OSqJoo4CDy1krVE8Oqg6lU7cBQeDiZjEahoFZCIu7v
wNPefuDQ/4dszWtA1MOkIjfLZcgrZGhOAuiupivo16UHjAHalzJ5OrgS/sVe6vkY
uSmXbWjwR9TT3TFMoFXZ/JBbt23loHHQZnBG8sFzjXrDk4lbMtmR4Xgkyfw7yMwG
AB/oLjyUqOFMio0AxsubYm+hIrgb2zSZtGOqX0ctiPkPOZsekfOJt+uHiq+Yf8Bk
p1SWF55jnM5NgYY/0+J6X7Z05VCxHoVKrw9CAR4XW2IrQNQeL2AEH0yR2t7SL7oj
7vrIHpjeI/y4mKKzeqvL4f2unJXeyFJodVm/rilf78ETEKUvfxpGSGLYjR7G9YW5
hnhYvROKyk6oTikibg9Nxg/hucDGw1tc8M7JitHyyQjdq5QwnZcjd1bJVtK+gRvc
8xiVVAUsGAfMNmiCMXOzZ+BwuEswO7isq8PbAEuRYqFMMoONGpvH3lDyan+YPVDI
/cz4EBlqX2A/nB+eI5+XucpVUDHL8ukg1NIXyGDYKeJtPo1TnKt4DobrtqK3FJw4
sfguck1c4rVAaFB4T9Ix14lRD4ExX3xBRggKi8+3IVrIO9uUCTfz6KulHkxgp8ZV
vXytpyArUI+BnJuzIKoD9Gz0yIpLxWzTy/R2JnFr6arr8nrrhLQFfLBSybXXWGlG
x5QLrR2aznvrGgX88LhUWz/ScTr6m1c5Ux1jUePQty/Er1o2cladf+IKd4EGLWbc
LmJGrpsFWlrhSJUjpabUEstdPY/G3c3vhuSbfYvjrM8CbapFQS0Y0tupKWqjxXFE
9iUnUd6OVxoTjdpf8qSz6Se0Rl2znIiC6isAVRGQQxW+Ksnh2uARiFKE4PFInOZZ
NeSEjmbKvVyVpce6vrKEmlPPbXo+B68lWtozDsE/YetZIif7Zg6SXG4M+7LNiIyI
5VFe/qAob5LjHb1Q3TQVIZpaO7a6XESkkPJfW3aOls2x+2TyImm/80xIhAKMqVSJ
QTzCWxcjRxPLiShp7FJoODDD57wQC7wsTcnF1rv/oHjndr4UYzr3BbRwywVCjSRf
zJPWIOrxHKNppc/3JcmMQg0zlPOZol3ZSaLZshtLc8+9CrQ18IgIvHyarvWPepF6
KKowdbej9nLk7axK3IG2ixFS2O8uwS7VgNC5NhFmhAWemPG1JkwV5yKHujtKfcxb
bO1Sm7MHX2kBcCqpRAaCv1iMXmQiN1xVtHtWvUenunN3SPM7kYqKhFqoKEOXJEug
w+EqL9Je2BV5GycTWsnDuzxonXgTKrmKF8jPUnz8slYwmphNKrV0/KKMStr2JbwE
EjSxc3fENEvtf3sNgsLP6QTAxDoZ6fZ9A55MaIyHJMYXiNOQ0SRqYlZVkCtOpg85
z5w65TC4jeTkypHQ+CcB1bnhGqynZj0heds1YmSPSlJRBqXu6eauiQGtEqFeKMpi
4+9v4KlHbH17L4r8MBldODoSwq4yryyD5PpUlHWpb5JLc23JY4/lf37t3BIK+Hrh
g14IMKVEiZkV5IIys64tU6/tEiqt2EhDdytGz3nncxReLtWPl58Tgwg60iFPFIPj
hSYT+q7CM5Pg9LLyT1gJRR8D/qVo71SnhOu8hc11N9bnbHFOnLg16Duh4ROYBDi8
D8hHi2PVLXTapOLUmynTpzPqa4+n+r+0w2U+K328HDp5HcNX3ZPArM2RLwEETmqI
EOagOIuduOX2Di9vKx5sACoeRW4wD+t3HkBvKZTj8v1Sk0sJ1v9nrm6kOXYWgUJe
00kj8LwF+O9Km7U95oC0E63qsYc0zcNhQ6HULoAq+c/ilyv38/Exc2g6zQ5Iq0I9
7oGxwM1lE3RKE58tEs4uoGu75iyv9VKFOXprQidthrgULxMpPiHWksDm2r3CqHne
4T5KdQN7LlfS0Z3CPtOd8jmua/uNXr3T7ElnC2vGuhYKNlXCDFYvjQCblztDwvSR
xRkP6bs9YjbO9XVqMKfAJkL33nUOdwmCsgtBEIbv3rA2gjGT+x9Hm8hqJp0xCh0g
YaYT0+ezqakWB0g52iKwHhq86Wg+CMFcrJgM6JYSfnl+SXKv6JAVz335oroppk47
89yy/VdBO8Yvmy9vDpPGMGKFsjDs0cyevy/OqA8yfc5txr1VmyjSIfCuW8ud4PhT
A07CWbCm2AzvIKOkKSRmGys3INPd/3YT7ycRN23BpUpkxqSTk1oIAJrd5KhCPlpY
Ih6ZcbxAzCB+xJXU7FWWnpNLLLMi+GJhxBnebgOKEBOS+W7BoT6k6e4MSg0KFBrx
MTRa3FSEquZ/8/ePmxpQDbGn/ikj6FdO7hMOF60rde7Rja5KwlfAodjkQXIPP0Js
D/woUQsjiKKNJCFNWXb1OCeVDBSZmBq97Wd6R5fL6jIkwV12lWShgwciy4RFBplA
IakH3w1RUp58z3y1keJKoDACQFSxx7ZncCgP2bB4MuGkUeeMxbOPKO5kMHa5JVEk
p8SoDox0ECVb95yYudF0eHefNTCtSWUc8hl3tIDjdgrua/hHR7uVYuEOJHEl0H0a
fDJ5ZQqw61DqrPLXQSGXfh4wrGOvw/RPXLC8zAPhDGc8VG25FVZWMhmzkpXMxTRm
NtLKorv7iq/K57gBsMe8JndKHoL47onc4R2d/0gBmjlAQbQx7JDw3x9NWy3DrDDm
UtDQhchosmaAQIUOksp5CktWe9CWGhUldmtHzYdzDeG2R84xFIVROI3rmqkvhJA0
EfLMC2SADEot1zIkEVfkHXojmjdrOqS7+VkDGKzzTgVU4bExVuIM6lr+Y1LVqCqz
GyZZuHLT+IznI19fMUUGiopFFqdBrjMZUhxEHPifuybAtuBt9FMXrBuJwT83W5oi
viS4zaxHyo2/3gfyy/3T016OLrUrqXp2KbRNPUvhapTUCU2nudx3L9n5YMbQN3XH
WOdh3uhHFR/6DMWd08E0tHxxGS3yC3mbEIRnho05hEAieOjCNCb9PqG4AswwXQ5Z
g/s9Pp1CShlInnQlc414Lfbb+WY/LAY8S8ZaZfAnolPPbBRMdIJn1l3BtmP42+0+
F+p9xrQHjXb1z8hvKDlgnr8DDKQwS2Jok8Gg7o+QQr7A41CLi8pjX5w6q0gm9XjY
k6cXWrKU5e60Ggh2T6LS67Q07Q7+0MJovAqiFRzDwM+OuYueeakRIMm+oFkzybmk
fZXxJCaFnFf1sgieG+pilRZSa6nLo9ZwmtnPK7+HP/b7cjezyqyZ24HI9rbBnez0
nVhhPQhBTkUASSrITnlRLz50mtrDr0uGZuuOFQ3+hi0MMF73VodB2BgFHSnHjcY/
KTgUOSjXPpAsKKKt3DPQwhKoWgjSFQm6+CYCXfsYJxI/eMpb7WkDaenmQ6Kena/a
+SLunkP1ktV7/0A7PpOU5nKCL9EQTTBnGSqjCqylxV8GT9AmPQ6M7Y1I22gXSaJf
oc35Ulr5QweVPkvl282O5sR3xXfvJRpzwa0lGQOFSdtqs6rjHGTkgU0b120Npfg9
8xsin87CA80s67aMRuv8Wq/FVHQe3fvxu7aUb0UtYr4+emGH2Aom+n1d4y4ZIq83
NbIvv5mu8/HDUD9E/gtZq/r8p02HOYSujKjmWS4kNzwaPOSwZAufR4gW2tJzhfjp
F6v2zbDid9j64uHf8qUQa/C84JmOm5WcPD3b/O7G1bWDH0ySf4mUwM48BbpwysG+
SDQfS642FeAP8SiMQE+X6FuF3I3zF0L0xa6eb3sB+iIL2ZDRLThGaKt8vkRJer+P
YFpX9BBqtT0ZYUn+hYoONCmMpNrGTvsT5M6Jc7WL1LU1RikdHi3VT0e013omS/Qx
kCHjmDo2xPm8WNEahYM5gn+9wIauAop0hHDF0bselVa09MLoDtd3vuLwp5c+nFyy
4MoHkCrcU/fd5YsPWf08H+hZKOha6O1LOTap+GfzsIs0dZTKnu18v+xHVgnmiFCF
c5M1pDmZU4hS61LIJD3KhhNImzEbfC6Tu1VcZYNB/WVhBe+ioIxeSjbJMpGSj0Ao
okLyFo0XiRcaSqnYxtI2j9Q0y3RXJwHShhE3M9TbzCobmArLZx8vUrd9nLkD6pdd
iiwmKCjsS+QfRswXDEZhWuvIghR13CcqldrHbfp8BdOo69/YbHFYWt83iFK9OdEn
gGo22VbYxcCk5Y/JIRUaYhad8OqPceonU9+A9xUME1kWcvIdG9HWSXlD0zFVQKrL
19mFaA9lt5s2lt3ZF3z/ElIrObXR6JCfn4VNIPj8XbW5TRGf38HegX002B1MUbnK
WDm0PsCWGtfWrRZpo+Qjj1TT0thuvTDg2KneuwfXkJsXrEaQhInhw4l0l/XjHqM9
tbuL/yt2vCuWWZainFoz/9cd2HKn0ocpzhltqdIxOINh/RLsxm3l6IqVQ/HSwg0v
sxcLq0wBAtny+cJVWUGfdF3ZNWJWqshygGwgDwo2b1KfDUTd6XaYdvvqcqHeQql/
bzAByW847cggKhfpveuRsDfEdQvqype8i5+LEcr/XfWHgIjijDPUdbg3v4DQhvkJ
GVUKnr9oMxUABqJzfBh1W1q6blZHxtqIhlPbD7aUhTftK+rGF31El/BdM3+jtTct
4T2nykUEwkyZ96bjcPyt3GKsBTXWinJtYEabmbOOtY6DTvv8DbmcqEIrpwXU/V9e
yD4VUY5lmBT6sjmUlBJNBcAbu2po2Rq3j5XIJEO6b+YpWnXTY0T8U5wAWjLF9w+i
neFHn7/b3UXasStTnQokZ6Olm/4xsSkpv1QII0/4v3oFoQcIfg+JoXPFuyeQm/0o
2MyEZ7N/j60GqtjLbbL+GSej/HUSTH1VuA7AUMlsSNatwg/tPj/+58+dC0k2Om8O
tAb4HZ6JBMXtK8Ia+Gnv4k7hGDbU23ZNUXOkd5MHa5lA6GSLp4MBtO967lOQTHuk
ht+8J5SoZkIMs9lfcgKphZpz9bi4bCSYpnXg6S13oTpdt/gvyFoSPZizFT+ReR/y
widx5ohbLsLWONAinq+OCtTvupQsg7EoCvGflqV38Kp3qL0lfcmUxyL0Ap0T4uzW
Y84/C7lX2EIII34ExOdV4Z+M9xZPugxEXn5ZmCpS2HHGwobye/urccdkhhS/nSPg
n8Eu/qyX6PhKh1M4/6mq1dVDVVjO3cHKtJS+vPiMgeSFSff47jTrQO32bh2a35U/
2Zg/f5LsK4UHq6GosJvQnWSLOkykPvgUpu2xoItWQlAZ2YzdyK9/oYcVsw15S3eb
vmmg55RXXYHS1Y10xYfgBlH6aCGa/gGSonp1zCpTzRW7Yq6aykEkkySKdsk3dGH7
zLTSQ1Gw76UuHdqncf7UO1RfyJQM30H+dtgSv06LVIw9uF4dzsvpCQlser1t8lna
ZufGfR+qNa28CnWjTy6JDN4fauxUHkAemDPl9iSHMcnwH/fKyn+KwQX14gs4xOvO
EGS27uphCeVM0SwJ/g6NPHwGJIWy1nxUo28DRoBF2hd7xcVw1OAgvxYWqAcUhpL0
yxZesJL5wCwBgDP2K2AmVlRi5HTC0XO9v0dmQf5PexRbjw9T0zPB0WjXGiv2hNIf
Bwr+9XQ6lvBKY8d6zNJ5rTCYOAHFxbYcTBZV+nsj6kQf07yLCouk+lEu3OU9yi8q
NN/d/vAzay4eolxUSc8mTWSx8Yw5hDuGWF2uwOHAKfpuSDgKWXuORMoo8o5pxleY
I9AUlSxGO2yxXVhT665gmN2ZAbk6zLQjUjYFWF9Il+jKB5FBkNTjifoJRPjo0v/t
/7/dRQT7o9YenQa5IZj6dBpURAc1b+UFvO1Ie1gztdFof/uRbHfhH+/Pcy74nt/g
0tRlEjTNROX7vx/vdULePaIXcA+aUcWQPapsNorHlnz2ZMwnssOv/vMM8YytAIH+
nnoCCCeUtUgdQ3/JzPm5wQT/FIk8QuZsOn780pXa9ArV6bW+2kJC2+J4H8elQM+G
Zr1R/NfyBi9PDI2uDqU892XwAi9KkGvLtjRYiw3++pIfwLwJJLU54f7qlTfhBM1c
pcQaPWn1C9O+1pBPGulSl1Su9EKXZvwz7mKspwPbxkner5e7BvoVgIlWOz/pdk55
qXYnHZkfXW55w7mqW+cCw+jAm+/3MyLSsqF5JTWOMC8ge/quT8CoDZhWlR/8U9Z5
sBGabwIqERnnEl7mgXKaaAzm/Gk7EQToBdzATKVwvuVd5h+0m2lhlkYUmihRH2ss
IOFDGXayh6pJ1unY6FaHnxjrQ4SdMJiuC173QM+Sxym9mKR8CV5YQIbo5wamgMLf
cIzCLex1y+Ry69pphVQCJI0Ss4bF47yxcf6aZo5MNfTQ6dBnoYu4wa6qF+uLGm3o
/HVt8SUgwhyBi4uaGmDcCJgA2tGcXzTKm45OiQzW5I71iYf3VZ4kIYJvFPHgpsuH
sjP0fY1tw/NuaeYpGKx4o+yqNav5Ua910/Min4J3YynH7w1lmpD9ZbDK9q0EHxLF
T0CdEbYPd+7QgdplQ6QHsVQApWiCiLwXgCd0n5KcJpUje4aVan4pQNqQkUPQZ8ud
ZryHlWZxzVaK7WDUYMzrnK5mvluM8itwht0NuZ3MkKj3latG53qS6C6DR5spQ5qS
hiqcykHloDLpRwdWTekIPpqrlziqPCrB59cFt/3EQE5DTlbGUwJERAbM9/ZMcAVw
25DfdDIRetjeJbUfU2XB3Io0MX023q7NZJqBb+tvRSsNBSm3UfCAjxm3dyfPHlJL
NYUm90EgXwvQBKeNvif1n4QXQSIbwS1HIR1k4w5dycLwZcIDjB/eHT6z4lhuhevm
/4I5k7WoyxkMXzgcDCcXNYPNVdQXlHUZLW8CGZkbONs5rDdwe0QTkS2Esu4fOdce
z+7icVBYRMqvZBHB+y2h+VrpNfoPgAkXjBC6wFiutP7M8Wqeo0WwPYE+ZGyWjYKS
eWxUTP6Vdzr4zJU+I8rRAXlwQmUQABtLP/dD0jGHv8LZAB9QVjhmOmUsu1xwKDuC
geeQ+d2457bsv3Su4S1nalNVVJ1IFbGt/cYGqtmAnlZ8cOXScOSxhX0rN++qrZDp
wKlsGAECkYdaRnV54wJi0dUIyXcI3ktgFZJLgzUKdSgCFk6HuDw6oQXgfPdm+0yt
cSz7Z38Zmwi04QmtfoHmJtduicZF7VPuQPbSNmmxoOgS+H4o++HsEyXwsTc9KYP0
2BydmoufwuNQJftHFyrXdU0RVo/4gFwfvZ65i39r57Y10vyBxByA1PVvLCL6hyRD
Ek/oZqEksIRj+9oXUr8b0w4l4arDyvNcLIlOBY3dFEKYlJ59UoglEN6rkf0QLuhP
BWrHD0Xe0Hf1J/4NUR/N5dtm+WvP8RzkXSfE9gNTMg0b3BJRIGrKT6YgE1j6s1Y5
2etntcALMTOCOyGL58iAui3QqE7ch6IYT/VFgowEt/arlBuA1aC9n/TH6+ilqgCe
mF/EWG+lOGDy9BhMLYr72wEFjX14Wl8U23/yw2+P7V0ApdhWrogiPd/3GH6k4sVe
SvGz/DsmgBDjZq0tDNRpVTZ6aNeeyC0/uiLi5NGaEzDkIKx85lonSpAm7iW7SAHR
iCdpcsR2qDyzhzc7CCIPDr0H0DwGVktGoj10By9aqyPB2WFjmqiz5ImtmFnupEj0
qt+wIaaAcQ26/YQCFjAG/XNkPwS/A6pPni2/IodS4335tYfp+IEAdNGH+V3U2uKg
WxxyvuJYT5EJPxxs6BMxX7MEYld/URTw92asbi0ZJzNYb5EQemGvBNOmTiPAwTXa
bXABQtjrvlXNpkLlmxfi2zEmmWqvCxsGcnYe0jwmpN0AzjNb6jgbXkX3CPMegy4h
JrfxQHH3SCiBHErUwGujYDQ2Gyy+6Oi/ySHiMgiWA0TSGJVtklg8PZpNXJyc3sCm
nqJHWqr5XTOp4kz5niM50Zb7M3KrhMvshq1hTBeU5HgYkvW66t2tq3YkSywwoDvi
rV+2sI5NIrHaoqMC7uUC3H25QWO5w0RiiWJu1006N696M3PrQHr917bse24s/mSC
GjbHCCn4maGEChtcEFahqx33f0b86MZdh2DR//PkwRTxlDgDzse5i9hSFSYEdiue
rxO9kcauWi58YgxVexWWIGb0cIrp+ojpRFqW9EEj46MN6VRMdQuLYf9gmp/USUs4
ryGFnyvsLvO/aFOsl4w0mF59R53Ag1Jh0es4K/d1m9IDCwGKnhQddhq2X0J9cuLw
tzBcEjop8/jIYv+14WwmmmweYT1KNw1vnsr1zNkCTHin4FrgINtWFMEze2ImVuYt
48gxb6WOC0a1B2v6CAKVQAFFwlapajgD2ZGsBH0yiP7FNs8wBBps9KzA4+R0mq5w
B/WV6Vsf/wRkPLvosFTtBB481kzHYfYLsZ9vfBHV0g6uS69FrtmiOHfcD9lIjGIU
486BFBKUmB6alU5yi/Wr6y8JQj4r4vMUNPqSq5dmW7gNBHcRpe5uerwHF/ZOCQW1
R0t5GOkYPU1F3PpE2S72lrDx59IXiMc9pJseiuZGBvAVMd8nfA55dMFoQl+tPbz0
7oTs5gnRJVOoCiAe8KIkL7h1e0CH83W8zlQIS5LM8zQI0Nq45LKlDhVoiw9ry+ik
qzEr4n2MHkvJPsIMiAHz/lqaKLdP14Lnhm+a8nHEHiWBI031ML9YsaqKobGqLAc+
Y+bbxPRlSn3V3KKgQ1CeLme+Z5Edt6XgOzcz5cFh31dlgETL0y2TVlduO+YInmJS
8yazSYRgn2bj8VBMuQvR32lNTfzn60cJ7mFy6V47SnaRSiXjDo+lt1uKHAP/az0T
evJBpyxoHCSqym0xwwIXSj8I+WxlIzCYiSJb/YD5TsJYPS8jxQhT//8OiSEVJy3d
iFvR7JZi6B0Uv3YB3zL/HVcy3tYMVJpMFotEYVn7VeqVx5cObtdDD4u3Y+y7NIgu
y8fNaJxWPShSQYRQnmwyPltHQdoUF1VNt9f0OKlDZSXD8N6R8zVbFYzMmhd8BaFO
7hVml/Tn+IlwyAZyfbRqsXljsxsLcQjeo1HKjSdxP5XidEYGj5pr8iATnMEk/VlF
JSaWpkNH6PD9OfmYKg3/sieAZ+f01+OSZjjdTjxCf7jUBYzd4pmgPGG5Fj/RCsRI
n+MrFwmaL/SbXda6STe2lhUi49XdWGrBkJl8KXitSAj7DgibJVYyE99jdSw78qzj
XrIiC0ILdkuttAmfdb+WYkyINqY7oW4231Yx5T8Cvk3v7Y+49sJZEbjdUYUSb2gO
3Apzuj/+iDnypD65K/7f5J3R/Wbxmxpz+Twh3ir8D8cb+LbJ74Vvs2j9Oa9/vHlr
wZ23OLWop9GWVt8fm1owXOliN1TpkK90g+tpUG6w6NpV35yP+KA4muKFKueOuEyM
4tBBLDa5ngIxxiHvI9VQgaSJNhxv7qBI10GqW6ZQ+63mjJgBQa/8sSQrwd8hcRQ5
nnRRefuSiSBCwCv4EO7Pa++TPBY4/bvCDgKuSWMVZW5Vc/DihtFQWOhUJqYA4/3P
XHb3ItaWpZ3xLvm2pkxQcI2DAHvt8ObKvlDSkMALmbpOv5eEjuUTfrZpsgtpJKb7
LYi2xMuZDFUwrHceZDOFpVgIc7DL5ewDqmVatVpRRm2jNzvoBT3O2jot0xWgfiXe
yETMKq9HzOQusmXitQYSq1RsCtIw6OxoO/VetF7wCXuB15mwUBgirnhatadBf/rE
LMs8NiS7zN8xOgPC6sdrfLnssR77UMy7c42ja2YlXW/jRsptOPFD5U1C9d04XBek
AbDwmM0PJAQOrE8hnWJhgV8rX6MCyzg/qLLaoQtLXhjO3R79kHnmkB6NOGw0ODjJ
3jB+b4Il9eBe33b0aXw2iug0I2A3kIBAv0tsYbP2nUPU9npsMgBgskQCH9fRAzyv
BFqKVXd7Hr793ixbjpazZKJdPv5pe1/Pzo/8tXJBCszcIfgKcu7NfVvOw0jwyqIa
YD9vvACbVzYrfWPbnzQNbWsT4Mp3LSYtYtAqjiHgErY2e1qX+JoOueJTnZI7wg3n
xzAWWvqfRxYQoqXj3b0WjZe4Ik7poxGUAuwjJPx/lOcPaKEevnY8I4TmI05WJQ+P
gQB9NRXi1Y9qr9ww8vov8ak/u7Aw7yokESlseM1D+L35bCz9UINjYrOElmS7gAoq
c+yf/lQ98JBUfqNsF1ZGUIy84Q6t5dGkKnwmNae+RgVtR+z4WPsiQQ8meebKyzp5
shdxREfKfpLCYYHRb5x8X3pDsnE+LenxvPpwWCwOwbytSfF3HbvJqNIzhjiI4Rwn
FbxmdfEYupvT/rRDara1h99ZQVN07xRr8oEijXPs/UvpoCxM/28nCKzMjxv1+QFa
2HXhf+ZDssF5lOc6lvJ96zzczu1q3zJmfG+CWgbqCAjcoShob8Q1Yj0SmJSSXkwz
eXd6x5XAFA99g+C101GR0wun2ZzTmgvkpzuCq1TGdxMkzx4BnJ5C664OrcgkrhoF
KvFdc6X8PNxHsruzwL0wNTRxAofPondFEEE1iJfIrQItpyds48zQtERkkXWWPlf6
hpIjJBKH8RxltyZLUZC3dUQW7ZTaTTxn+Y2oar5aLYhNdjWlUJfEP+rVK8XDo9QR
1znB2foVAA3Pva26UKVmvWf2xTNEySZFK8JEETJdvG3SRY9ch0G6VCUyoKPXaIBv
BzmVGLh33l69Rdy+B///oZDN+CiqHuqQS1hhmiXTquL6+9FykKqnLgPBfWCPg8qa
a8eukRsaGtqVITWw/KZ3kh02eooUxs6jGVmBHjzFOIdk8KYOLZSDWQxuS/mtQhwO
FQI+fE9kUDiY9J1eMkLFDgnvD6r0L1kF9lRY+8fOnqJ6GWGNJaLEIY9adFjGQGby
YyAfmshOmwpNYHkKe6eOdu78wqFWvyzyHIl31ogaMBtJuweDh98QYQ8nGf82pW9I
RuBBF9MkVMiy2ek6prGt+39zq+OQqU+Xk5IVpLwyxazxNewmLQDZwZlfxjl3HqGd
H+doC8T7BGJ+y7G6L6CtqiD/MaE84k+dk6GsfYV7Pm37LEYFyfYXRjTTOLhZoQE6
tKqsOc1JZjX+E3fRYdQiA7UBhHkQDIaLjVDWSecg8A1uxZ2oApbf4wqvzpw//QCa
E0vVqvSukUOG6WxLMo0LmcNZYJIf2UqEvnrMXkC0XFMpbZUMPuIdPaK59Qd5kshp
5Ys5Ggl0LjjjBHSlxrhq7p5HcSDEQbyiZF4OKVLNSD7F8KVgBvwd2QL742IoIIdR
w9dQTtTM4P3+k41CmcmYCeUuYOG3krqszBL7rsfgHIIIDktzQusQU86THlsc7od3
sQeUHdl+xljqy0jEMTdsMRDiGCd3ua3OIVmhT5es1LtAEFWc/WSyFH5YL2xJiyyK
04BQgINNOn/qsgjOk90bTt+wKSJlXvmmne5fnJmKD5C9s+pj7q7zc0CDJ6Ixq8uC
6OjyPJhCHrxbxzeA0ytBrE3wqk9JjmzUSODQMPcotIXfXN7wnh8xWY4mQueY1KIs
DSNtyb4EcAEkdYugEr9Qo877bBFd6I3Ii5hqLkBmtOPE+65JRhSrk9SM+Gl71bEP
G/FfdD8HLAyirQD/WTcxUpOwcZwrDlSpG37RJuC+WW2xSzMri/UoY5z3Xu7iY1xZ
EJOSTW7fWQMSVj0qwl4y/hF4/fGRoNHpcdcKrOEJcLMaX/rBG0vQrauW6to26wVI
rFbs3Zc+SluLbsJTAEyTr3AQxT17uBHXakgOgDO4WZ+frohK/UHyIJQvYEsnyY0j
+vNISF8VGzsJ6EBoBebbSEX56oJaSxjjjsIwAL9RlYdz6IOg3yq9HGu3CJ7ohFqg
z56oXMZrgibA0EIgMOTc4HzRB/ugvA1Kg76FvMsWrIcQ3MrWNQG0w2ObsRHW8mpn
4SUvDTTej6Iha9AgxLcE1tvdmpd1eBySTv7dQjyPf6E1DZjCSzBXxDaZlIvh0lku
1Ess/GPQuFBFcdSMA6oqN/H5xDWpjeLfl+gliDLdwj5UGOL/nVvD+CS1d8nCIK8n
+wwppRRO+NZEtoJ3qz9DS9/wJIZbc5ihHOLkqSSNYn/mQ5ukKQY70tUb4vC+viyC
gB3ssYJMSApozfI2Ws8JAoQY+zaKo+ciQQJ9TizDIqiWaRCLnSM/IYGQR6xffWLP
ANl0i+fyk0l5Pc3iD7Mygzjzro3Q5HUBqhET9vOQVN+BBKUT1yWeYiJSAc8zMFNp
JwdZQU51gyeYcqwBBdqtEXDjZZAmm9geGUM2a4Hliazk+eLhL3GTXzDpNvjwQkjD
acebKWZY1cYMlLZoWoZ90PY8GYx6q/fQD3pa0wcnlHOElbLsI8W/Nmwe/kFvaUoZ
6xVC4nDv6Dr0QbvA0E2Hsv1zQO9NsAwyistfFfP7TylJsp8bPv8CbfoB8TxknieS
b4gftvj6oC7SfBPtaRDDdHoODfSGTJU4mYO+HCwvg3pOvC25QrPMm6zFaby02ZNM
iXQtbCRn+GvSmR1sNV9vGQiqwaKvW2GgdkYUuIT2M/YhGUxVlkr2JT/I8kjcZu15
NiELnFXd9ozbmWpViHMi0WqHSWRc9KZEYn6wmk/GFnCPD9XugELSC4W/pVWKlMcH
36vxnOp0dPA+1Smxh84UHKLGscKFLchQ+43ho0K6n+BC7V/aG41/0to/0JLNnEgk
F74Wi36/8Xeb4tihQYqDn4ECi+Y7F1eF0zhc4aRaLWOPzO1kLINle7Vv7IkgKoU8
sV/0wW4BYmSv1+QGHeXKdrM8gl+r7WkgQ06zHqIW9agmUbFgKz4RxqIbHUy4Txdz
R2sb/6yuD9lT3pEdxwPczXs3x2TdqxL8EEVCX2tLZ1QNDU7bKW1vEdN5kU79BJX/
lrigME77mwoPbzOOhjDybc5Ce3ve6h3Pkg7Y3fFQyjo15wfuRVXl5yneG2lUYAJu
XObwSDN6YOgtDw8GYICHFhSwjVxXBQHpKXD7POPd2rub3weP+CjfoEcPFsNsYpxZ
oVyUz2uK5w89kcyPqy0E+u8IMUwfqYTEqWb+QpByAOUS1OMV6HD6KSkAbyiUwE11
vCvz+lKjIjcVARvqaUwT9BeSiZKK3hq0qG4Pc9Nzs0lzwOUj5Zvfvn9Y5TBmhu7U
kqMrYIJturqUhXmA9RS4wnlDuFAsPMxI+kd5n4dErl1gS7JU0OJdnvzQ5qZ9DNih
pVU8DNtqW1Zklr/CJDh0rAG79PwYp6aPs4kJ18dO466k6KdFvUmC9H72fYbhIc4J
AoraBPIjs3rs6D3bD7WLElsLkF9VB1OyRwyUiq54dMr/8V+QbXUKcb+zDyc7ZU0z
CWfi240NDXadKYXWknZxZENhIQvYmoMPfT8FRgKqCqf/2m0DUEk19mwxbzVSoxsR
jzhmKNlEalKdU88VxUdLx/WqCY0rYharm3NR2rZlKlK6phC2kXvfo0qqnMlGujsC
5jbW2FU4IxE9n/Hgor3TxjPlPWVP5rG8x9Sq07FIEg11p02x/k9KtFDpaUfFcrVz
3ZAzfih0yT91MZXa8q06nZkeikQlVYGKHohu3PcUDBqKLqKe+d/DvAaOe/MA0On8
jGlZbaO+QVXWXBmipOialgq6qTluyibPIp+bLORoGKa5g830oAmdLvYhnmQZFtW3
amKvhyvZmDB0kSuswV00Vq9DVtAyMNopyUl9ceLhzl3Y6tuiVG3rgCC2micM07cg
IahnQoV2apu9Hg/NgAGSoOE4SgbmvynnOlwb4xt6hNu8DnSly13ORL8zu+TPcXXJ
pTXmpdKy78w6WQpDmjIzHy7oe6JyCWF54Qgv92RVcaUWrM3zcNNFH3PdkxNnO/ay
Wtk174W4nljKvS9Kl4sAYJyy6FZcUZmRCI1qTxZP5GtaxEbBDkw9JDqCP9OQTXlQ
o1oMJcEDFMVxlniT3t6cZTDeBVMVIPcuhkCcI0RWXOw4kubvGOPoSKqrAmL1WyiP
KJcQXzJ22gTkC09KpUZ17rwSxQoN0t43HStuzBPEj1C6VcjJwxiZ5Uh1PFeI1w5P
V2T6sjKBvDcd6qDswySJhOMbjObO+IQN6ixYwz+dJioC2tN40p/szwa0939qhzHX
afVYxiROFuZ9PoVJ/twZdFGTIFaBdLTWg1sP2JNVebYJ181di5/R7QgxcPuWbkA9
n9dyUKJmJeVgzMKM6qYBEzNANWbuXSAfk+grZKPhAOKc/5urvqJyF+agnT+PRbYc
jPUUO/zMouiwOykWbfJwbYXIlhtvOdGHUEixHcjNMdf1jXqLTdyMNVR59OSDGA4k
LhQzONS3e93EE/sxvlLCublyefnO/aBUrovbDkY6CS1BWGgNJ3PEikG8z09NLE2n
IikRaY40zYheeeO+bcyuxxVi6FWIWNFrwrql2XC3KvIe7nCUMr07eaxkGHTxdX2h
/RAw4arQKRBIt1Xa1c1stHibc1GJtigl/ZkYNgFgI1FGdLTWKO9jPS8LE4OryG9j
SabA4AReRtiGQD5GV7nOjuP9iekINNFy7mjifPO1rReT3np4wyoeClV32TWLPNMR
qU7w5HP5jhuvGzXI0AL1/KmEd4qs+4j2yYKVcAfTW1znBQMCoGG5+uE0tY7nOiP7
XxYX7NIH9G8oRWpOUxwyK+if+nlxLB+iACnp9npbIzD4IgBqyUfCypUzh8DnYRzF
ADVV3emaEFXJ4x7wh5xR3YVTPmT+FF1BsRz8gEl60BoWfvuHUw5z6M4rBMtb1pch
frL6kB8gKCbrM7sLQiCOMB57jMXDd5lqfjLyU5s8WXTj3YtLG3cbo5tJKIB7Rt62
ds4LwzHiy1srIu0JkbGJmsV82IXsuD7IklaixQdBOZT87vB/3XeFr1yAShqOnhDz
8p9ZkZdX7dkTAk7IoGQtCSkDTn4Q46bhUDo7iEQ/ZYG+iHPl2akx9VW3jr5a7HUh
/dwkF+OGVtqiciSc0PNK9gO1yJmwiM5aZo5PoEAUWH1OpdQQGGSGkU3t28lv55XM
MeSBuaPUiam2BcuwpWmp8GYu8Y7n41pcTALKV/r/zWAXax7k4Yo66mDJ2xNll0dQ
EOxoVRYLH7pQuFdMup/sYAKVDI2Gft/WD+oDUTwHTER3bmhdprGsyj0eklZN3BvR
08quy1U+91BLRCxsQDBf8m9t0nlEWCnTxVOHPOzQSRMZxJmZtGkkoO8C1fae8nQB
Uv2opZx1BIb1hzO8NPgpap4IChQEX6kCcgEq4PGYp/8o2rVyHfDx1IL4DjaG043b
N7edvxnPGtoPggaSlZ8j8PC6BUe1qEdp0nwhypHFFu4LrftMJ4Fl4vNHP+9VtZz7
bupepKaFK3N9OhZeTGotrspBOYqvzUdgGHWfaO3Y7Y/j0anWYhLJrBj0RkV7O+Du
1eRHF/P4hrcg/EcW7ZHsMz20WKkHJfykteoG+BAYz0eH1UIr3jhscqsrpPX0aIen
6Kx0BmBWBdK//S0XY1+7Ur7YNETi7L/ZgaXlibLNS0d1WA1e9wB83EZ4I6CksM5v
tD2VpqXjTKvWVSfE1zTCFzv74PQ+nAhbZUjmE959gTDZT+FyisHP6Ij62ZxdHHmT
36jsdRx1GCZiVXEsU5PB9Bdu7Snz0NAlmO20wNOYw+VX4l3GTBgs9L5RfioXWNmr
BwlqjIM3k+GIJZh2wS8VbMPRedlvbTJ8lBEB7S8+astef3t6s9IeNfxonKK3cK0n
ECupwPrBZ+qmHMrXfy/TAWZ7+cYwuQNzEsYBZI9VODv70/AI3pTKuE8tSMvRF4gs
7yyeXatTI0LNm0v3Xg5NBRAwbX5/RQJ11y3VV3u7eYcs7ds/srz0qT2jMQ4F5GLw
mgBShe9IKM5JnTJHSdgE1jUcExjTd1rkjWBZ0mgnyFlTyul6E0QlZU6vJoFIYifS
U/inyw8puMg5d/gu66Tzo2R4iWk63VJx3n/vGfyHUWImcn98ANcKsTwup0OQ86Gv
WqSmAEN6aOhz0nv9UpXQVDlS7sPp+6MSuoa3raI9e7M6EcZ4ckhYipy9V4itiRut
/F8CxOqmmY0kICG1lvyxp2EuDjjie7fZNRB/cklwwwFMGi2P4HDmvUVbgmsDNmye
RSCoZ86VU766DwoFer9DXt+DLocvOp1aWaGd61FaiWtb06oZnB5sy1q4tigMiRW7
9JT2QBavOk+qg8t3AFaL07n5zDDPXQEww7sNDM3Yswb+BMMZh85arN/OFDVux9Ys
KKpGK1gn4hbxlwRJjzEdONihfkT4p+3p5iz5Vi1ho0g+qzmjpBLq7zISiK5QuAGp
GuQ7qpjmuZWiLxgXIWifW/m4piiaOfrA8h/Qn1mrw8gFkBYqOqxJgTi4KL/JiExr
Qpf6bOZmTn2DKcSXFsbocZMPv87L9kzLyDpaX0vmMAHk016reUcSc/XHQ9jJvn8o
ueBwDcBs1lD0Y31AolONyY3ZnZ3qN6fYHp+71lzMvXWACVGlUTBpm7plpsl1h9CY
a0e5a0gNm8AtU5m63YjS9h+VkdsfItJ00lETN++mytKFJP0LWHr5uhHzADIBc3AG
pcu93uSvRld0XYeWsO+zwEDG1ohR3OBZk82u9ceUwnCYyu+q4SOMbNYek+49sxZ7
lvxGtyYgXK7zufYqKqlRtBPdkzMQYo0HHlVljCVehxi2hwAvEhzfa9O4VmROXAcQ
N/jZ2hCuy6XAVMZhtvRyNaLpntCLE4iM/FTkI6vKMOL5wmRJrWhSCNYWIF4mY9T3
lIDEmWiNqwYMwzuBPqhKns9CsJccU7ZsXLQVNVTsY/SXaOXpfUI5bKcUrUDoXy7K
Z621T0fNsTP4vQWTGhUeB70nXjYPEDIpvkGmRLZLladqzGrIWBY01UmzGxbcLIXQ
DTna9oFOI8r03z/BWcEbQEqX4f1I6nJGBhvDA3prqOFM/FotA/gTZiSHdnN4G2gR
G7ktl41kQhZz5+naN2lXLGKQ8XE19wxBc+auMT9TFWtDTPDjHai9rLCfq/eKq4nq
nuxgH9yZBjcXuEx/NRN7GWcNVWJ+VzHDNvjSFfdDLrHcV1FaREsddA/yNNP8hy2O
EjPMyveDO1SLeaT2kGgFvCzanN9Xb15oOzgjTn8Mgikc4j6KW1EdSTambJ9vLZOu
2Op+WXvRquS8Bmok4CtBBd9KgXvnxDI9UBMO20VzxOBJc6Y7NDygk+niVgDiSqtf
0Spf0J8Rflb6FPixGl90Bj1jVu2aqW75mFLcOqxrOqyDjarZi8cT+PGuwk1f7Kwk
A942YcseCEFO6A1p9f6VwjCI+iXaE6aldgvKHFjf5Qnu1rOs8Txvn1MMHK+ELctC
DwstAvpMmJo4cV/MxHZGGzuKoNkjq1gu0xEhpMgmZB+vKs333E7VoZ8JS/Lddl4L
Jge45oWM39EsV9/b+3iGmuWSEW0gi0MNb5/0mA3FYbmqVzRMmW7pOzU5RZ2eoYH5
3yVBA4lh/5cFxik1uU0L61o2Ye7r9iRuxilWhQEHSf3lzqABpRYtkimrUWpO7CRm
yVNaf78gp6KUliSGoS9BQFn5VR5FlCnTHSSm66mWqqTVGMFo7avkCWb9UmcGBLgI
c83K7onJ5LYnHcf0PMvdZoRXco67DGl0S2AG45QtCXJVZOzZFWSMMlq4gmu7Trkb
+wtlFqgVcNz9Wwm3K0WQ1kEELPxm2h5ziF+mMWcMJNXFDREfB5EX0ehKiYWCvsTe
EY46eb24L99D6d1x0v1zzdZXKmNZmhuRyVOilVLmav2jR/YEGsgIjEsS8Fm9ReLS
oDX54og5JY/N3vqEMnMb8NGtRKPjt3gWU3VvadEIm3EYXbvDhB5BayHkCHfk/dP8
7vyNv4nHdcBJXNo/59d4l1Wb5KUrDJGE4QdDpNOEqWqSnRCYFg/09cNtnvBlD+uG
A4YCbFX3k0hnKx85RKm89/p2xYvoSAnDFuYr39Y2ISwvQW3i7xDkMngnCLihyCv8
zjN7icq6/MAGerCe/J78MOEN93OassFt9NNoAH2cd2WEne1zW4Vwz8ur2tj8v7ra
Ynss/Z7DSB+UGGdzDoZGz+8s4GMFoXbQvXP2djqGX3OQ5ANKdL+AVrjcgflHG4bB
ZP6tv5++iPLrPPT1So6GfJswcqRARaY7qzCagnHzWF+hiRHoAUBHYWo01zrVDpdY
DEHAMBBtFiACId23MWu8ZvhSO+O1MC/rCvU2dMR/aO1MehP9lQmJO63fJzNNI575
Kx0dgs8ngbnfwsqNd70bsg+9G7VsDDJNhxi6WIK3qf/s5vy8aKo9eRGY5NLdImx3
ubkEnREb1RYeVijD7Rt7JvZcpH3hKzX/2efo1ZYX61ddZs2C9tGIDHpvw5WQomZF
g9QqVHAX+DESTPQv1qTQvaMAVN25/6cSL+dr0/Lq1VtQhIIqqdR5BaxLBS9GCX5m
S2lJU7oyKiuS80kiaWNQLVqTJUatBhDKE16/WB7aYUXH+YFJ8A90gz/LZ3oAlY/v
8rYY5ezLAOXssGLArUAJwj30suAW1XWn8O9NUr4YnO4yQCstwVpIhs1oNMEZGcEq
GK+1PxaHpIISkyDy4cH2EuOfL9OBo6QW7BoauuaMFNsLb0dEWpdBs3tskizUsSBE
Q7ljvkgAyisqQF3p5gKEnB3iBq8fSMmk0fsz0kPvHQ6g03Mv4RtG31k7lWx/Mox7
apHynJ8EC2ZCcHiG9PKm2j0sf+ZuTOnarYys6ayzTZu3hppJ6x+BU5KdbIWcr0x0
VppdPAv9hOSIRdnOnvqzUo80WUaRpI+AcK59G09Xo+hItCNvfs360ZIsXUQg21zl
0PBfXgn+sFRenNrUQJdgxsEy94amRERdtRuuL6ftSIpfThhhDyb+hy/X0jLMlRlr
nDxJ0PENGo7F/zAYAYDI6qA/JB6rR7ymCI7/Fh9FUi2dJNt5cBNfQKZzg1Brl90w
cJimKLBhj69XUjr0CBAbLAWe/6YCU+zqyxeKUE4+E863FIxwUJIeC0nFGvBrbQCq
IgFsK8u19hX07+CvwB8Z8Nk7MRvzpijLEcT9ovwCxJJimAPKCybP07n6n0KsVZW2
U0IIgfFlK+pGMzW8x1gVQfGbQqlAPwlbal4hKkt3YI4YMsgs9FHFoFF/IdyiEADS
w+dpi47hBJofIJx3UPUpleRpO4nssrLtiT97bDeTtW3qNucSpsvKJ+TgOpSUaHHK
2lMaz2W+leGYwI36AXVkNfKjINw7GFcoOSMiKk6EbGA61AxdvMenQMlCG9P/TVNk
hP1GdjBNrbI2LbinIKm+PxQ+AJvk84K3Jl6XUX9KeCxuYvq1q/bpJWWiWapMRzQJ
oDTsTXJ7FVkkZE98dPHgxdXdBNhVFD20nSEwbe+uRpf4M7py19fGJkymtEcUkQ97
QlQl8iCG/XYyk7vRR6u10FdQA2O/5GIPib5szotZcmkaAM/ZNbytYoJL+e1Afto/
+cUqTTOo3fkyPm2m22NLWtrLLrfYCeuv89juZWKUiKgf1gycpElji3kSNPfI1X4R
eMs13xwEdnPNBO2J8R6ZBJRMT/aX41Nk8N6jPIp8/41YFPYpOwHhFu+fxRUhWrn+
3wci6mP6Aefxm6nNA7QFOJVth/3QgQb1wt/MGsibHAZe4qcHYIKRxpcNi/Q3Oj+F
sLOwiSz94qdSOqXmtjFH8qkTOX/vYKiXzOjNwZlxwzMHdVP7kP3xtzxlPRYpPbnk
sCG1AfUyTpT8fb5cmErX1xsQd5f7HTV7ClI4hwsFt5e3zHmZ1OB0rkfmxd0EMCG5
usfXmLFUnpoq+QNbntacjwq6s2TNdgUeYpK5Z/tg8d2brfTnqqsjr3Nrunb82y9d
FZGHD97M3Z+d2UwuGasZxIgGSQ7zgi91Z2oD4hL+G5vov1XBkpPEPJJKT2Uemm1f
S1Qo1GDEmYY3XrR5ozTvAxiJxkFi8YSCnkov592zsQMguqru6nGJZoUNUNsk826R
ibXbMdM2zNQCQgcBk/Wswb/wiMrIPCAKxQOB4qIf+1qjdjlHN0/Mm/2BvRjlJSVw
N4pHdjBMvTwVOOTU/CJ9bg+m9o60yxE0MGLgZq2mNLnSAPFNUgtM3EQ4DFdI4fFH
KFsrlzjQOTM+4QsSRZsbeAY6QUNorN/mJi53sTzgkizXqAPHTlDB/DXpVdwxpC6E
Jh5gztmqmIUWisaqytzc2RIl7ACJ3P5szrLZ1jIjyc8lZI/ks2jmXZj0grxBRSqF
XpDry4S5lBPJaUTq6SNO4rXXCnBnnKMeL5P44sI/oAH4l9NGlrKqeraI18QCcGx/
I7eo+QcFDNLNoP/JWUXNU18vOu+svKgBVPcXNg1GTLhL7YvlgSLbRyMbFYURrS6A
3SKcLVxSAFZpbcwHbMO6xflPN8/k7tGYEbNc94BIWiQNCcJdh0gLZRVMpBwtZvAH
/dKMJRq+70hjoBmclCNo7QS6uViyA7RnCPelCwTUl+dF1mpxyjLu7kC8dJ/uCKqd
sFbv504V7ZPVTgtll/TDNe4lwH8MNHuSMQpZmWB/4JMmwBeaUuyPN3TusBdJvS4k
7AYP2s7W/Bpic6weUykPMqPdi8BbalWTRKNUg/6wkPYe1880iOCJYea/CB9TO5MB
seAwKu80xb7Bw2GYsZWLMFo1O7tDBXtHy0KeeD277LdOXDqcb9ftLncHvk9kdOKr
NN5V2d2ijm9cI10fM7YVir1aF8Zc4mNGAgW+2SqH2W8hDmx4SkzLsjn6fkwxj1Ym
loTHKi/ugAMYKb7WuMWWKvZSDbUt8uHsbHb6jkNQLwGcho0AVnXn9VSKse2U4yfh
nZQxiJ3M9cuYaVXueUSM+K8nPLw5vGkH1TnbtuiS5YOxDDl/e1yl2z/oNIq2Dee0
K4EpOulDm7BAuIVOd5QkSK4ZqrAbkJ7g6UnHrWCNc3Jg5+BKrHd2KZ+bi1sasRm3
C4Z2b6HT0XpvkXGKDXl7LssGi8tjuUuKthc9hKL5XWucfc+YZFgaJcbM+xnkokaH
SFei0kBhoKE2AzTxYW5/9RFwQi0yXZnYFmHI7ko9Yy8trqv0L72COCGRsYqMaK/0
AtwvEVMZt8rS2mXdQJJWSKRpNU4odSVVkeMtb2AOirMGqljJIXWTT+c4qqWnaE+p
T+oVlbbnKTjIXdxXe4C1WzFfpC/EnQPRC3YpIQfOsRAcsVCjSYhvUchsxSkdXUlQ
iSCpSVADl/h6gri7T/x3/hMu1Xm7XKs64HfZ4ypLbk2eHE7i6Tc41RLWwZyUNRmT
98+oDT4APqt4kA3zqMSo4BNPFwfPARTLtw/a2dMXI1kHPBtvLm19VDcaQCizpg1W
VTOUxzX1+lQ4hsfyg9T3SlBwo+MpWWDJHW83lXCSm4smLmG6utSTqwmKv+U6/H7r
/FwWnR3qbQ5TG6UaQ2FwllMZcSN0tdErQMb/aA62RuRS8oQWUtOQsgULCdCX4gcE
TRyK5dhjf0zvBX5k+jTufnT/RkFrjfxri31o8JjSCEiUiRJ2/WJJ6WE+sTgtnQsn
im4JoMqitN1RpmiI1K5ck7Ff5NUE+ArHb/kIW0y6HkJpxSlmD1xblD6REDAlzRLS
34pfd/z+nhJAnosujK20AKS652MEUHiWDB6oNsDaXJt+O8uJioj4HDy3PYTMfM9m
y8cu2t8jbZ3WUtqm2Uo1fbePhhOswhA3DQ1b36V6mT9sY2aocNTDm+QKUjO4gzkk
usHSUoKDZdM2FbjmTE6ZGjXPewtmLlN9MuhsdueZgUav/5UeOZ5qd5REyfEzAjTY
IALXePCS8VifH9Ucdy9qkLlL2trEz/6Wr94pn9N5z7l4i4MQmusjMTgAno/J8Gga
GDvp+bN4S1CvOEcsCIMXTNRipg5rVlZh6Xm12BzTL56qvg1iCbUg/qRVO+OqG9Ys
eFljU1z4T/UAmizrG58sBCvGPQ8oefyFcowNXb2uqQhzvStSF53s1QPMfHh52/It
7tBPOzsoxBRdRmxTacROPu40XnCiii7fcxOeE5YL/Knj5mVNwS82CDv07i+vE1Pt
Iwt4MWgOEJ+Boi+frPiBnsL3Bzeb4lSLNENjh5ZR20JdKB4uCs1mbxdlBGjsLPQA
4L4ncxh6HFVHdHX3rnF9DLR7O583ihhNPPaxhmV52x/w/wH/uwg9/3xYyTvff6i5
gm3l7dSLk2Fr8Hs6OGGMWnDbGFFzOu2Tn5scmOa3lR2hywZQKsOK7Sihhq7o7FpF
EuRCg3qj1SS1LeBKvtT7/NqbeQfk6gCCaPtrIflF49oJKseZOD7+B6WmmsnanvYh
d4aQDTuraBAnkAOr2PqpPTZDG9bSfJdEmAFwTgmsmyn9tTKVn/2VXxzlca0GER6r
c+tK7kuq0wvp+Hk7kHxfsgN/wGA+w/eSkyU3DUDlnUJBW1OQzzGknhYaur0sYkvv
EQbgGPZcd3yLt6VIV5EBLSNn4iz/mE61UeKFxfdrcLJqd1fZFmMkEc+VWS+m3omw
D4mGrDMfD5fv2adspenO15mAjwe4aKkW/47R48tzeKjJ1knFm/NAtpY5c1E9ecJ1
WOHyvEU1xGyQz/W2t5gfKb1qlnb8WvNmrx6SSTvZfoSopDM+XaOUYyeqbVvhhV/W
wYlLs6vghWKcKBk0NZRR9E3RvfDR1hQMB6nNMn7rlOrzR+HkmWkCz8e0gzy02eye
svGD0SSsMEIkD4L+8VnQoH6qIfrMM6zcxqv4YwadEKLhtmJvim6/NM8QppvivYJ1
YqNuMvyflgAJC5S8EW+oGHk48Tq+QVctTjcJRrA9i5py6YcYGBbv+NEEVJf2ljWw
FO9Xa9WCuDts2VoqSAUmoSoMJvuqDqpCSshlbJVkIzTSmBSfKJYzZUlV+ixeATcE
ln+2h3jJNKcHsBifSduyg5NpKMNPFZO6vL75yXpkTawzGCNdwnGDYZ6ij4Yd+nGS
b7kwV4PGlNXVCtOrYghJ+r0W7BtGpHZPRtLsLOcbf0XNAYN83AZBwnKgbcsmAWWi
4Jzgcbymw9UVWN7IgmxFgcSr5pmrEMZhdV8+HX6k/eo34nyGmfC3J17JhhNNU7Jl
RPnWS9N4EleTOqWvPXx8Yrapr3q2v4MVx4jnipkwIgDk61opDndxnI7g3ah+/kqy
qCe+lOgEIxR7ctvZMSPL/fwW8AJrF3HCgbfgpUYqxUkabR6IVr3acqZlwC0apKxm
XHwR5Q2bU8nu6PkO6rHrsWhh1EFgF95u9KW4EDOrWaRmh2CDKFt24heTR+FM9T2P
4iFR1gf93ovHspkpQGSl79Sc+3iPJlcrqWQpAqjTGjZi/2SehQeqBLpLvF1fQfn1
zvJgjRCOuGvmTGALVL+8AnpM4tEUy8Z05NVD5feM/NucP1nYOHWIZsGsl4osMTb3
/LXYKVZSAKa2B9xpb6JLYKa4kpKs+uykxehEwzJdTYRfxdsTE9mrGpndMZtJj9qc
LX/4Y8ArH3KEW7s/LaUMyAUyskEMd6Y6quKUw+Lg0d5pYhBbtbayuXAvHtXr2PvJ
fYLAMCyoeEITbtdNwXxzDxA17vmCgH8SikAUxJ7l28yHMoRdIPpbAwJJ/JdDxiTp
YkjGkSCI9Srvh+6JPg3CYdx76raG4nxz1bSuq47Z4/vHyzYKffAp093JW7kYSsPB
Lj7FAXhhTCfvaZ9ok98Ez22XLLgyTpwWioHShbwoP6eI1htUpZuGBILQDsxW7FsU
cCRMwQFLVUxrR4KI3wbAdSm646mrKklE+2auj6zvdg7Q8oFQudShGuLa/oBNnu8t
/Y6hqhiCgeE8+WuXwnbtwJvgBBoj3n04yy3Vhh6P+m1CeGlskAW931Vx8VKQbiVY
AdkOg3bSJobc5jMcUAz1tsRGhCBn6j8eAqoEDROa1juiUSo8tnCZNSqarJx5A6bF
rJ3acET8yMx3zlr7NTJJNhMUpuWpBWhWI9hKZyFC/q67vU4iZ8ISdSgccjeojBaT
42cneg1kLGgoRSFWfVNeGxCMVNkbLl8SqiOGSHJN7UHsf5M6SkEcjC3cQLH+Tyfe
p8TUp+xcBwiILrNL061p7G2TyMmh3HjIf0F3wu4pBNAIOimEUi9doHIQx3O5bRLJ
uxbpcxb6Vh+y+16ApHnkLsQGfoOTpVJ/lc4uuSlp7PWPTLMzd8EJB6YJR66yGZ1z
ObM1HldXdun9ZG8byC03phSEDaMnQgVP/Q1MlS9HT+wURbKALHiyFHNtte4Oz0pg
JeNkJ+jU0QdO5FOtCqdhRMVpU0KWWvlLzI3blM4Z7bIOrjhopB3KtUb5V6rp8Org
/eDZ2zsqVHBQe4sE1NlOqxvGOGwcL1/VZWrgADKGwcljp7rvrYEUJzE1R/A77amT
gd0fc4ErmmJ0OWaAupaI25DJf6eB9QQ5scS89Ui+FQdbfzCHcZx6H8hC5OOsVpa4
PRfRLkhMqXlKqZEIhfN0pkEKMV7ZMzKNzyMzFmhF1xrs0NZ5U1besCy3DaLjkaNc
4h1plMfPCy1Cleg31ON/q2AdpBqq565QbCb7NUHMk7zRgVHs/qnhSrs0Ek/yDt0U
pgC6JYaoP12WQgt9109PwrQWRypa89JNjgtGR+T1jTMNQsi6qjC+P3AlWZdHd2Ty
Ssjz4Qb9NjsluUlo3HPlNB57u1GLjTc20TzecVZrKQzCWlu9ZqUHA8DhFTDrzywt
H/0NvOKsPpMjYayhhIESMMPN+fANT+OAuezxslPjdfAye/wA6sDJ89GGtWIlZ3Nl
wZuRhCoRB0dw50nJUIV8cRkys3E4MXhl6PjJhWrMJEN0em48UaNyHUN3iCiNWQXc
AUfwpBPOlwbWWDVIk6den/j06ZTONF+PbUE9RBRwCB5LPi6CIMk9UV+NC5jmN+se
6WpC2HkS23LR9+xFlxDE8YB9eeRDoiGDMkcKCEgyjE9IW/scOfXas+bPqMfF8x3E
Bw+VftpvGL4Plw/KK39HBvCZkZ++/yhusTCs8HVSZ4WUevKgFNDX/v0fT23bWoB7
3HK0fevEQUrpihnBUytEYgaLHrdD7rAKSxDfD+BqJXqZi5IGQIS2PO2piwTpX49F
75CdSJEhklO9vqclpFIgDjdpHnVg7Uh9W/RD7SECaLgdE1GSbWyHOmeA6Ag3k7F+
xPtpiv9AUVgqouVgJxr3m+VhIUqPShfflhssgVk+SeFdRmCWa+DIzJ7X+2xod7CH
gXWOi6/QxPNV5gl/zXn5fMV9hNFqgaOwLyQ35l5htSFsa/yQTn1WMdi/ydP9j+KA
aDbrWbnsBU++qlCHTk5Nwd2yo2YAhpiu1N3eJ1rQFgYtdexIRNJJf+BKXooQuCuC
S2Qq9GOJIE0BoJ22SG1xx8fuK86q2WX5KUqExTSx10WLFuuxdtg69yUqoJj1JqhX
vJL3+7rhv42q8FG0AWCcjfV/+JzfL20F8I6a7zLWrCdwhL5ixJXoF12BwMCqLCle
Cc8MaWw2ePwM2uVsURhjokv2ZVi53oleVc+IxsVUDlNy+5D/GkMYlt2VpGXWhCYf
Kx5WKf1p+2Wo/2RSc2hRM6M2DsB/goFezsFm4JLFRI326yXpPpoigj/Pyyg7z/Rt
GBJPA+C7g+rFJul/tGn/9MoS9ngrbK27AEoVCswf96zz40sz+T//riAfS9Gmg7MZ
fKh8T0emDOMUesSMm3qucG1RutA0UhNT1Rw4m/hsnfB88hVkHivrhNuFisYrbKxt
850M9vv6ckBbNBaNJsUpGluBgcdtoM4W1CazayoYKNnNO4yUW3pWiDnOHjOgxiN7
kgHBWUf5+k2O8NxrEEXbDBDn5TqoN9ASQk2SJZhy/pbhPOMGLcWmi4pR8L6Hfpfd
GpuocJZDEqC2eZqTRzksK1NSkQsbTmqKKpRSMu5vknPgHmmNQ+aLdN695RDMpHbP
s6ySrviKDThwSOlIox0k/ZCpE2C7R3PCndh/GXCsxV3YEuNPyaexZZL992444Sdg
DjSdSXruZ2QcT6DA7meuzWsw2P4S7rrZQFLz+dVALjzu/XF6iPQRaqjhB73hcuuW
l9iXZvln++WtPzFRN48iwO6xGEOUpZSpK5UY7z1jFk9miVpZKdN3670KQdu9tG3q
pwPQV0//JM5VMjSgHKbhWUoYPBbeDOKEWeEB3fCpX29Uzrz/Rd8PsHIFfMmOmQFM
kUfU70AHb2yAQlo5GXPb6KNv+qMPGFTxjCZ72mvjuCulmb5Mb5HZLw2ZjULuWS0n
PCLdPZ7PST+WrznEo7aMmUE2xtbq5kMhhuIBqPRVjZaZ5s+mf+XHqGQF0klN8h7P
NFMCeuXFU1C2bW7qK3PV3VAnODF7RkUnxh2kYSc2hoyIyOl7uJTt0zQVipmJMROy
KdJFJJbQf8I7qIhEMKVQ06N3n8+O0GO/QhhJivNeERNH3Vl+xIsthZARsMwtfcqY
aUeq/wAZi/7I/zfgBgCmd53HX8z/azRjzP/jqR7TC9le+Bkol3MhhK5svK7NNa4M
gVRDjVVXbwiT4TyRN7XvFz4Q1GbH1eWmRy8+NjHhGOAWDsXv0P39PpV2ol8vQOiy
V+qLlAOYQ/Zhn4O5k203shpAMaeLLdFaFfSf9nTod6QI8PISkqU2Rm51dBkC8EJG
ocXOC5xkkroaCnDLPMdzEMoHYHc9fxQwaVMhB4OnzAWmByplyzKYqSXONVYm+2xe
REWO4xwgwveras7xTyNf0Px7nZT3zZeRixZjGYrjvvGGj+epB4PQNf0MJ53zSiVr
7OL97MQNkSqMyoiPdN89mOp35Mxaj43XjLsUymAp4GylGhRW+aEDyl1bgSjJnkvC
Uk7VYYKXyo8R/U2ubNsilVtHSMricNtTio60/a1f807Sj6oa/8QjtF2NwxuUQUY/
Huxw3PlFSpr1gCkyXJs3nZkymATjYrgQQESjg0M70xlPR73fLlLP2cpWB7wXOBrJ
Ov+6gLxR8AcAB9TWwTIkVdmg1jkVigNEh2DHMkTy2kKyQy+oOVgrZEgZ1i5ItbV8
JgP+JkdaKc87LjZ8Fc54+KFn0OG+ky+1ezQZAGYgwGmYkp1AeDZzvA3669NHsRWe
iszunO7PgNIpZTFnfQZkY75SbJ6mqekUCwkjgTl+a1EYypstRZLEtRTmnSUCHRS4
LWGWI5bBpp/kYNwV8fRchWFovcUPaVZ+nGYcc/9G7tC6Qxp4W+7mA4kLcZS90Cxr
EwAdhLpOgqyWXw1ar6AZlKXGttBVAJYu/ImmDa1a7MxHMKtj9rWBtXzWNer8p2BM
iJi4by5dCYC39DkHZRFRCCVgOoWT+PLjAL3ZEp9amm60pMUy5CFK4vnO3dE/iMDo
WxzVcqSQyOA7ceQ8dACg+A0+c27AsHue4kiEWYvHL90kCeBrg1IQSxV5ySa1DREX
hpMpP9xPtF6ONLjCt8J1HdPi1VY721ET4AHcA23vdzr+gPrJCqe3o7c6UVSsN3dP
CfllEjUKdRehlLesQAMt8t7bSGPYrhbfX0gY42YuKnx1kceGAvVQGWA56Il0Wn1k
2d3tWD3vIcmTei1EsexjTDNSCi+K78H4G/sfaMBG9NdWpWNWaq+cL9rPLMa8kxF5
WucMzd5icQpn76dASeAn8TMH/HKT7bvRzLq7wKp9OX37J/HJPgJiMFNmJ3/ip6TW
NU9oxe7qLOAUm8v2/E4SjRH1k6N/Vgepal60sZYC01iq5dXD/puZQ8T8eTmcc5pW
aZLbge0c06MvdBymgeNBpxq7qSJiEWob7OPZBhWlPVkHUBLTBfjPVrKSAVZdaOoY
b2/3mgNLnW7T3UwkZ7qFufYn2XXOCadbemWYAYlEn/neeL9PpwPixaoQSBTgX1HZ
UArI/tiZ6sjOfDfQ4AcqNnXODK99lno2IYwYWKzr9imAzx3JaQCngZN4eVL97bGI
qrGJ6iMa2qGd4aFZ+EkEVqXWBrKkKwqT5dOicVLAG2cRWcOAmnxzaFNBifxAAafV
kE4Vsk2IDQ38iYlGRPMJK0pPjG4Qi/jq0JhA17G17H9cs2oauhrPrueudXsWBZwH
zz32UFJSYrhwL9nAt0/l/2Q62cEqdjW0fnHro20Qdm8Gv59CIsi4fe9mxiNPsBz6
wXdHMsxjhxwvygqrSQ/as2siH1psMM7lAdTSQHEsT04NpWL3bom8Cs01HoOvjNk1
s/l5KRp47GaeSWfIXgyBLlVgqJjhkLbpGhijSE5Qq1hpJXiFr6kAV3n0MGlPL/cJ
RmH8VpUffGBxWm1ywB5nOZUBZEBRi09EcFEliwKQG/cAUvcOiEtuan5jCorzvJWg
QQPI3hHLNen8HRk+jwuioosNj5iJk0ZRywhl7LiaBkF47ZV+JYzFdMK7A0aLZ+YV
BjMbf8YXWCo49sJC/TvFlsMRuKBUvsqJso+tDKwVugAI0FGG+qVaz7mxopfG4U62
vn87uXN42VwaY0tlSTrJjrbadQgPlVWnPE55zkgCujifLNgGMIJQE/E+aZaxus5e
Lhs1zyy6pmsPWbKJUIE9whhlOUBaUlOUKd70zcNmnz3mY1HgLZDfc1rJGAgLVlus
t+FDgihzCgUWKm5syCJ0zXhxKVpaVjS70VRogvffmRsHP2QaqlCJb1wZdBgyBxJK
NssFjSRD8ThOhKQYbHUVp5IXviRDUwaLldSWGaX1XXYTN+LqhetzxGmQl+ZLLvit
t/SEsdfS/2o58reLwD53Ti7h6NGSkkK26KI61C/rElnosj5wcS+WO57hpdaVDRHb
erWPRAbi+SAGnLikx88D21h5goPvgj6eely7A+g9qqT0WXxKNUC5PkLyJGY/9SJw
xb6d4xOOhO2ktt7b3vuPayJ1oa/lcs5O76Y/6m2H9fg+zl+UkK7TZDEUGMa7xNEJ
DuzLfsgljMMzuHypPAus/OdR27fFLH1FsEYzQ1jKSmteEteCw6Zk349U26NlMVrb
XT3onZ9RWcKhrd5A/ssDG0SlCxZUOp67lxYMC/aX7i4ViPp6cJyFpOcGQmOWjVSN
jUJUpjojjWtKZ8JqGHYke81emoK632y4ItJzamENYrJRrgAg72rTPXkKaGObN+/s
UkcLAxMQglsaqN27EeYwAZOlDvNm4ZRRmndzlFhExwp4091BJ4W2WR0mMsAc8nVl
G21zybm8wsjgVfbmSjihI0bo4c887ujwL2ZVZxJnoFUL4Nr4XtxCks6wh5yOqj0K
ViJoiOL0inuxnJeQwFrTiktTRckZ6u67e1X3VgWJSk9XABY4TzgfwyEVCo6b9bvW
fI08kzArGzynpegspqoVz2+16wShHOfaiTyZbUe7ICf1U2dWZpNNo8qWPMEpki1v
FAQoV88W3ru36D934v1pbjxWNT91DfMhZ+fJE5YgIYoThCpEfZeE7knxOqeFLDwB
AlgOak3BwEhzC7PYtWUcJWDKN0ZuFnINdqWwuLuMJgW3Exb75lqpvdIS6+Su2YiC
K/sGv9nlpWFzqT1Qi5sjRpLIyst7CVizaJo/ala0ZatjXkKd36L9kcrg3ukBpOZa
IkVAOTLMzvRiUhkTEa/DEmkdzsomWmtkhzPjBV1d1RorPWoc3ZOziQihCMRMpa1j
jjZC8Jfkap/7rWfQ0r2lE+NgFThoH46/6gOEjkTsDolOm2jqfm62brqddVTIRyB1
s35uf5TDrbP9x8N2e6OtcsEorBWxnH5ZDsDKlkBrr8UUqfCqQhLYCdADBF9f/3p3
FYvEdHWHyILlZlXc4yC8/Oba8/AuaHcygGaUM9wgwurIIOW+P0eqhKEMUTf8SG+z
Xop3jiBRTTWP4TWDfxMt+98Zp9wwKIKbvfHOQkMJ4FEX/N69KvVbMZYbXiVYVR2r
uaaX95Mj1tAk3LYW42AKD/8AO3Qg+oQ8gyXYjFSvASscdwHUFfRyOEX7DB7Urrt2
hFK6mgnzRB0O5v15W2KqfOmCQIWmM0FQaVhqPLJyo61P5td1EzAIsNb5z76kqopd
FYBeCJ6e8eNfoR1axIfdrOvBmPyT7OAXQtpSgw4xYBt9e3i5p2kDGXG3nWLJ/0sC
ZApBRSrHxC6oQkKb9B0Hr/2CctqrzBVsd3C2SMwFo9Cfcra09fLhy72CbNwks9Uj
V8UeJUSq1a+QS0DyfrHbhHv7RThy5L0ucVV3mebSr2TFfO8HFbfJr2ElBbcTEigV
3ifWEPhyTcovvjNa40m6khUTm8dEhmbVR2gv6eR/MVfB8f20QooDt3OQPyTOeQRC
/iJtFd3iZkzn2oBERm3+LdYHPvK5/KpyYLXmhKeuD9jgn4+ja3i5hfNomC6BMBHW
yZjBMwjg+HZv9RvzNSQAmxM2AcGCTcAb7tKNKnXJIAFxdvDpkgvNeyRGv+3HG4C6
n1wfdffwIQqfYeDknK0DTwJ7yvcHHA5WSgVJkl6z+ZvNBpgGqg9qvMLK6/xT0ZNg
2fVoXr84bgSfcyO7PibLqrzf/HCflcVC7MEZN/UXVDEOhHqzespp0Kwg53/XFD9Y
JN/I7trzRrXhaPjRjqNLFz+KVrXCA9Supb/WlMTSuqNme5Vl4FkwtaMiWHVLYkIW
pCIwbt0VkwlugNmMqpUhkkWT9/8xZI/V0biyAdRJmPrpHecq20BlEYu/dRPWhaql
5+vWt/LPtbtJ+T4c9Tr1QPg6CX7C/6v68eR96iyRt7XBHBzMmI0lhjIRCVa4Q33g
ogX6TUH/itOQnD3I+vTRZr+xX+/BAEqIqdmBQ1/tZN8HbRYLU/6xks/KCMyILruY
Rm7zzT2XPUwHCPL1kWUGqojmrbxRaC2TtihbNdZgBfT5GmDZgIQOmvfW9IBxO0dM
bq+USGeROzyrPIG0ZJvKuXKwGgtUk8lctkRHx/PN/UKeEmZQtl7ocrwfF5FEkp8i
gFu+S6E+uxHyV6cJm33XPRkJXMbT1Ult1Eub9SZlPo0IxbV2ZKV/wwdz63Hhn4mc
4/S2cEsRsgVhbfJAPtDts2AIvq0bd2RLYhGlXvU3pzutjDg899k2SvimEXRjpDRN
McwEwIWoXTuFHsmb2LvRgo8Tdp6JoZaYSCYDOw4hLmXacJQHJFrG67n3VqltiZiE
jowe+89a7OMIbgzqf/pHW+KRBsU+wwqrwGtA1zHnA2ZfKQavCe07OYTa/OoCnYaA
mcmvUjCR9WduVA/8EYNDvnAuvKro2HEiJYmN/ZnPfNDCjzsPDM4ll2w/NRFEtaAC
yQzT+ZpeE8LetjtkeXhXiBdctWdgcIJwVWMeMk266WLBuuHH2C47unGN9Ky7OLuk
E2jqRu/exH6EDYMtlQATwq9eoWjQr498fSEJ1J7H8NPPI4Jle8XrbdnBBkBZiTSl
+VdjuHE+sOfoIum8uOQj3cQWLayFAUmQND7n2nEcfslzpJtfasQip3n92yev3Z9W
bY7SF4HpGmz1SyJJvSNqUy4LWzc3UkfObNJunDDIpLlDDsqulZbRr9keyZpb8dpv
H+lSGPSwWWm8YJbDydt+kJRCcVv73aWSf5HkWlvOmF4Szxl9JmJiFQujPIPL/RPi
dnHeurfwUDAjpqjmBy3tdChtZC1btbO2E4wucBYQQANilR3lMMPG3M1xnATNy9dD
pY3dfUIs09kdHIoLHyPVanyKTdG0V/NVQeavcGH+7ceShIPJXi/6IWMOw7LsCa5H
qSOeCEGU5quM6hu3ghOLhuLLSX+lQpumiMjKlWZEFv4ouedODtu26nd8bOcMQFfs
d4wKm9YG1oOtRi8MmJOSYu6ldx7gIJ7/vky+rqgWYjecgYKQSkXh0TqWNJ7IjesG
Yneykbk3oGZuaFRhtnhebtbJ2sV5U0cEOON7gn63pffhV77FJJVp8Z9mqi0Xjkl7
tbhoQVJ7l4w0e9vI3H78MX4/CizQL/atRVCw3WrN6BQkn/Dbloc3IOwE5iNxmqdd
EWRI/r5a96vhXUJLBRUEfryB11EwcOY4TX+fWBrCjI8020q/Fb06oOtF8NuPbz+m
LK+rHtucipGagSZs2ph74DbD+yT2BaMkVZmdsWfeewdtuGhh8oMdixs7U2Ed3ZuO
WL6Bxr7+TsLj2EdLkUUSjQmEnGsd4VWbAOKGjYqNgSuaB3iwMyY/ljC5YRUK6A7Q
8Ehe3GD1B2wc9wzbxBPdnnf0B6AERdyiKIXQV5Uom4fFdSjST1POFmfSlPX6s+zY
7h07yvukx59jn5R1T9oFVX3ElGPygcXjeiG5kDYFOwjFHcDeFzxv+xEnq2JSlMhG
FvjSdvvNsobHNW+OrJY/Gp2l1LS6YsmO16ojBy0zGs0Z9jcPAyV/Av47BygK8noP
14NpSZdp2iJ43CaZoNWvkJ4sWkzIyomHvFOX+8ljCIOG6SoLtGNiW4UFcWWhC3/+
sEXfbRpPzGbH/xHq2DT2rWDJum1112QF7jr1/SE2uQsJGOS6GZI98H4cNKKXedEB
FNM9UGAovhcYHRy4MZC89YLknDAQ6CQukFCt5zy+x+O37aH+U/g7W+oODsBOKbC5
dS7+9vQTChEC8cnEcjAejIT/Bya+kaBP1r/TjKxmrOwz4+wy8WWXlBP92FBLY1iS
TRcc6vjepJ7mdZCyKyxdOY2KPVAxmc5VhjbS7f03gBDd4YGc8PY69U9PR50HNsdJ
SfgcT9+T2Y5yi9E3b0dRgFn/OjzABVxU0zjSOR6xpgEfToXkvYYWMui268wRl1UD
eWObOzIHCgTx5E8FnN8B0QU1iJUtRksW/YNLHpjXxanVeF0dIfO15xlPZUM/sMnv
0TccuVUldEL5XmseWRor/A6b80fL5LqJ1rLrQxOW+pxToCsGhSfiTI66wO7nXOZl
aqKrPt4RQO2I11vxj3JcsLW+pAJWh9FYBJQkTmS7qocxql3/sPBD29jvMECpIwzA
IxUQKVxA1PGspBeyO52qwiOb82ICVE7DLb8maamigMqZw3w7f2XD5vZ3jJbl6En7
+s5hm1kvrfM6JObcf7NLc8WPna3z0zNg/qu0IPujRFKR1KzlNa4N0zOs3qO3wUA+
mZUxBI0WJ2uXI11Q/QjzZERIjrxZFYJg/Az9OXZ4Ns2CUprraNiIeqFvXE/a8qkW
divbYxBLmfll30JEpsHKLBEqjKvGpjeAz50oPdsNY3DZgUTybmDsx/dpAtLhqdTL
8thyLEaudDtXpUk+8pIQLTlR4azBfaSOGM3RwfUUn4q9WG3+g23MhK3ZrDoZ6ce/
By4xjwGjvwqmantJLS4/8epckw9SAodqfUc+cwU4ayH3rX6ocAwzu0SwOKvTGkrD
7HZBlz5J++mnfJmJ2PagvTNAiPXkyrooGRbUAxzA/Cguz+KofNOmZCwts4UFEmOc
uEiJQ0Sz95WtxQtKr9s1/g37YSJF2d9sMo2/GBSFsh1i5dMImYXtZ9tFKO84pVHa
yeAy0aiU+872kUhob0jeY049CTxVLC0mdLcb17GFWnYWLISzPAbGrV/+yVxAr7IB
ZBUZk6+uOokFcuZpeUHjKTKl9q/gQrIB9p7X8t82RQ+8e1igzqVlGhdWgqIAfNLH
UiZ3dhMqsVl+cj8QQNaC6zG/gFrBBdRCbPA1wOJUk+duI4zAkvysQp+7UWK4wuXR
eg90nmPWn4HeYrc5QyBkOEhg/I35QrmKc/7NB3/jwoqa6Gl99uTp6U5fl6aHMd2Q
taTi8wdl8qtNuppsBYr0yBPADTZLuUGUD0FuAMUkrE/6cg2mnZRpGT5WtZV6SpHG
cQYtSwFr6H/B4+ZV2NEytZF/AlAHJWqkoSvRn/vGe+yAxGPZTZugWgST6JNCt6V7
NRloTi7bDfoBezYjqV5bJvKtYgONDVN/41b5MCIhbjpPVMjaoWw8F8+U54786jqf
YjcoGRV2lJR4maSDm7swDHsHo9qvMpk5fGaqrk+2G5XQaGXTPezuUWVC7LAWWNDA
GtwETkvece4aCIbJb5GHdtGyaIiCAYZRCcGZ6h1DWtIAwV4xOEmwO89qu5nTRGlN
ZWDImVAlTmR4682+2US862R+VI0+i7YLGMg4oVjY7fc94AfqpONI2SQctuZqLbYg
/fMLwhacq/gtUyxyPVfJC8kHu0Lle0bTSge/3u0MgU3sA074LBidR7XEqZ7KhvPs
hiiXyoxqip1168FYXCVHigZfgsqq87EeWERCeyVukO7VsSFnCeVXcxDb9jYSLWzI
fDwP+quVtmS0NnRB1dNan0IVg4kKTBHuUlCu+NUD6PqjOLAFtuNcly9Q5eU2qLBo
TX9Umc4ExjlmhajhCGObwZ8CdxjSauC4Fu3+O/usA9LrwREUBiqcZbzcSUnb/K+O
ckil5oaenDcISjBs6tf8XoFa70yfFWM+IDeZWRGUe5Sx98GWzCGX4JsQOCeYn6Bd
ss42YU6kjvJMoqbXkFKCBOPDkT7jDDj5goOSJuZwLpkZAg986Xq7P5JLGhmpZnaP
kHYGYeXEVy1TXP7DLUW9aqBVXGnjA1CINjQ50gnrirmzkNxx7WX7nER6gkC9dD1q
fEUvXmP8byvSIY/wtGkokvYQ0dklXq49mo6OqDx7MEdd+6cAETx1k3/wv+pUCI1V
ZnQl3yXNp0CZ81Kgp0nbHBAl6k6ruQAVwmq7P2RJ+6cUyYo6+hHjERSRs6OR+/aZ
wA01vcehKZAP2Q2Y7xzoC7LWaGitO0+OYSYCqYySr11rqYbHHAMlHLGI6EGf/oHn
F1ogoK1jB5hOksEM8zg+FCpWy5jTeXdarPzRE9cz2mnWvTzEVCebIv2am/baHUcN
CTn5uBXH6dmdsWV3/fIzFAdKf8JVeCtn05V+1ufnfBxE16oQBHpj2IFl7GQq+jQg
RJTuQeTMwa6DHy8yFzukXVuGdXUUruoMx1wR6NDlX8tXRIi9ocVGXS8Znbpp1Brq
VJ8j6/EwH12zLC++9WEf5b+DUMqLUvQsnrSlaENkUA8w288aThGyxgIjrSjlZW4u
cqKUlZur0Fi1KMI4J2ygGRyT8PXNHFDtk7V8j6SOmaaQ/AbwUb0yT6+PCgTs1Dt+
kUrAjG0sKaDu5NVe2D4W6KE67wfq+TnfC2ly8n4zohRzt0UBpfAulaG29aYyzQmq
gSNt/Yk/Y0bgI2WEmq46Bp3A2sNeImCA8YwyFDDzX/QD5L3TIcP6Wx9B4vvnHqSY
d4YA1r97f9WWuaLEuFf7mZzzYvlmbeDh3IOO0lVuZAYcG07o3/0I/UHzikpYPhwi
YfP/Ce6JIgkHUn8IPWVovV6faz8S/cu1BEH1cNsMidc4RFrr2+/Fe/u6PexOiqJ0
z05mCY7E+RCYMo6Vygu4V3xmTtz1glR/MsfG5COfsOFRqk96b9RSd1EhME03ievd
HKD6ZXCVfJokntJ7t+dyiRuULJkxiPjIUnZ9bCGOuUFrp9sUMa3OEb25vnHP22DK
eLZX0wcjEr/NkgD0y/Y+E2oDe7CbSMmzlnff32cBb2W2nPaOo7QwxVihiD7OZNOW
Nru8/ayMJqxC9jS/A2PdgQPDuGQb98t7zDNtF48w7/Q7wdvwmLkBTb/HUsWnvVS6
0BPAOvPfGqas/G1Z59TDmNsdK1NeV14HmUsAXvw7eAdxMuxE9Jqf3as6JtvExbAp
kXg12pcMMfdSAFku/tG76q5fB56OV82IqMFk3QBolJwxbNrSEkdK9GvufMlaQ1fG
BrYnP+WXZJNxhp9NeOwRamPCG9H7tMP5p94SYyi/K3msTtZnhGNvQS3XmEscS/kC
jiPCVG2ivhOJxcjwYrux6rkeRPeUX8rzYViYQVEInQYZSDFM0FdZcuNWwuCtytNI
YSNdXeT0jExNdmwg05yISn2zLwZA1N01uw/MCy/kzqEK07jRePoowmGGojHW9X+E
VeaYcBa+Jq+rJCf2l+jC64SNRQAPXQb8pcAuClYkBOMsCCCCGIHMTE+5jyfDEKPJ
wrDeug32P//W7N6ZDyOcLg3NFyaWDvnaxeQrY5CvkWppcDm18rTkLY5mgoafl3PI
TjtrkR5uNj1sGQ++fGWS7Q5oIeIUHQaSdLlaU0foGCRsYCeQlyymR5fMFv870JZ1
PFplLpNkVp2okmr4rMjkocfKHmtiCrDywLg63g7u8JJStEMi5EVei+UtToBRGMnF
Bi7wL4yr2gbOlUttC7dkbPxV2bigq+FxLg/acx6j5G3UBgKBJdBof/7LZfWE5vsM
YWmL2TzK+hSqApDvLyfjm04k/53zQkwoOyvLyVEnFnq7/MLdtI3GcCJXeht6Ymyd
1FUK9zhHgmiotewZMr8FfRX4BVjVECLe10CKjbIot7z2yJ2ymHakKMmA/mDpmp9N
d6+4QarB4zUn4gf7QGC0Nwoysd4iD3BCpPYF0XogwC+qqWFeWlguuPepQYMSbHbF
Y+TpWO06NURD0iW7Mxod22vpG8uHveErpe8zVGkFleDkxjH9kl+UwFlOWbZYCCSW
ToG4s9GdwvS7xd+/6fz0ZZzabyZXWT8WZU6Ciu+Ay7wrOxHcIpUMwRui3dO4UMmB
bwls4FWFScceLyP3DUQqjsO5PnRo0PwTLIe9xm8GIW7D/hmG2Hj5k/llgmJjwao0
P6EdpffttnG/ClpKtyaOmYP/0Yon9LaCRko8UZGqV4jhxGy0ju0/F58FqSeiNybn
5wx4SZiPMwkAkHwgklUQGhrS/ka42a+3aKrlmp9EVHs/j9w9ErgDOiZCcH4GWDjy
WHJArw7G2ZYxePmCGycqOnuUeyNTFZk5XK17d7UuKecSus3hXDEM0MBzgip3nVtn
GTYhTzsMqpswmeg14Y9lPS1uOeqdbYIc9l6E4EzuDLJodvJ4PgCfa77S1zoJ1izD
48/gGQBe4Rk8xXwCnp9BSUVR4kINqT24rREZ26iW6rJKM5w0PtrA+k0mPv33anh9
D9fy5irvV2/Cj0FZbLkAuEx7ceUA4Z3+HlSRzmWnhIl8FX65EvOCpwaPii2WtA9R
FDO1bThUa1cM7i3+2ncHNvZcAAWcTgwmQlqga0WvGdnOHL04Hlyj40b70gGyo3sX
re9XekTGMGjiKaxxAAdXDuH+UgKIThiJLCDLlmoPti2zpgnryjZxp1MTqKfg83IT
jsJ4LjRXv7dfUFPvlivpl5XTjV9GfT5Wt/xYYZ6obCj95e+pztSM2i+xtcLC8IWV
mLQ0vuI/XnveG9NSCHiwVwcqhtGd3jF7b0WlpQmaM3mkAPhG5zGIfNAZ+VZKKVGb
YK81KgB1MLiJiV8IQS/jPKveZGKfILAxX10cQmD1A2rUizO8OWBDCewvftdWHp6H
vRmqlApFGy7qQQ/6FuI28l2JIlTqZb6f3RSm7X0DBTxrltfNFsH0vfkco6Dmmaa7
Hzjhzog31eF6GdM9KybT+o9HLFESctRum71CrDelKcExwPnSAz4dRsybIbcr8h9I
0aDcACTvh9wT+qyiLoKDqJrt3YMdtnQcwb5/TvOE3BYbRGtC7eVtRxksjH7D+Fag
I7nR2DLrJsuEJ+oEeVEzh6iTSpyy/e+m7NcCabzM+JVXP4AfUFMoqwufGYHjNsIG
p++ZmfXiw9Zp/3CyGHQ0ZS0zcweAgVrFsNQSiAGWLqYXaHY1qHeqbodkA192Syr4
LO8jsiioxRWThAyCa1TRK0Xr2OThS/msKTlnczM/odxwi5iuuYZ3/yE7VEtRdiIG
DbVjH47dyybJEsG5RumFaNXXfmiCwLCcbbce8Habv+5BkCuKY3MoY2BYb0+ChOj5
HCPvDws4+HiMQI8qlKLd6AU9sNzQRd00mgkFPFYyvhen+4RaWoCYcmR20DI/pEaw
uSDqSc7j7UmwA2/htkp1fMjvDnUi8V98ofZiSStVQZ+1Wj23qwTFgqBxTiPytL7B
KZclyLUnRSDJI1Z3PU/ok0joCHWuhnrTMqUL1KnT9h6+3mWG+cQ+e99VQNAAWXFD
JNO+eQMJti2C1cOFZ2OVAsahM9aqqslk69DZzYzg/yy6tC5692JH9EHKUcGXvOmU
BdmPrbZslfqwClxre3ZuEVgGYUn0eHKcZmSEcdOAv7tEXnn/X9dRAiofZfIcPw07
yFt0/27uaYhclKv31/ZmdTcZPduzB2ORPXUVye65RiPsGJjQOIcR6/tmuJao21+9
PVmjmt0JHY7pd1x6FKCVwINbNSjBzGKxyUp4ZLDMqjEuIqQEh6bKseTfIzJpUGeR
/06Fnhj3KjI81JE9a8X2CCmvgMO5h5nAEakN9ZGGVMgA5OEX/mEJ8XSJpzcNubTl
XbErL2R7EuKGsCu1sq9FXNCCZhOGm473n0G3M1J9gDw1m5tgenFFsNHEfLCAB2Df
DBy+kj63tp7goYUrj21mYRonRj1X53iX0rFkMgV1qQPENVGfZ+R8j6zNJIUiOVo3
R/qKMvgh3XdHomn6PimwuOKEYWG2OHnIiX82y6vWBOgZ3/m4U6Zgz6HE7ui1JwQ4
FTfL+qrj/iCqBWwaBP/NwrbVY2EGpcUxeg+5fzvuGaU/83N8qtgkjHLCRh9kdyhe
8qqRHWddYC67x/9nko9AAyGNGZDf32KlsTbj/Qfd9LgZWGru+CEeqyJLqBUDAQRq
+8cAKwsMWUsmgCsdCyT+FZbdG061LfqF4AROLnfzP7tgdmYhGhriU8znNPhZAxzK
J3F53EttkXc9nu+Rhv77LWRo09piXNmUY62/CtrWJu9SesBfT/aLuZOrYEBaa4k7
BKHtfqMOlqinonN5eHyQ44H7a8c9eTw6X+wcajJ0ZcJFwT60uv7nwI63BAkO9wSa
4kmLivaGzoh96r6l4n7cmsxLBWaB9ysykZagof8TU6EvuhWSeFlhxGhR0VMAe80S
olyt95VoF22pwM4Dx+QOiJl65h6Lb3DQXoNR0fQm+dNk5DrejIJuYtawrpJvaZHf
i/J5lVBeS4c5c3iJPUGdOPg0hklZKhtOZvz8CKNS4UaJZhexhEuBkT5SX8OpXnNM
90+WOuJLG5CVxRNVetiX5KQyP3cDeKulGF8M11D4+bajFlAiqkr+SZm61aN539C3
62a8AZv3b1kon99l4Q1BWkJ/gtNwjiyEMa6aZHbeFLeF3/tnMaZY+QQ7uDJZ2FQu
KB7HT3XXVpiSWf0t2uxNbsnzAWg8ue9eWuVLNkCfq4xU/NYFKVKx9NpRr5GHE39H
EeZIaQFEOfRW1G1bj+DZNU8yiD6g9XRKKSIWtbI0+Xg/EeEoR8/XItY4BU4dJTvS
nlchztuR3JRjcJn1tGs3egcsAqhHSgmuGoyUH6YJsbOJmzEMaNds+V6N/NoQ/ukY
ikp6nUc+47baE5NX5AMI5GDjoSfXMTFf7lhwMfvfuIPmoty8NGkWKpF3ODqprRse
/0cg94Bev94+yDrm/ovVM5SAv8wPsJt34CZoerToxHOHjAr5luMZZtVADKz4glmw
eUn7pIfowExax8q9gg/UKFcLY/sBiy1H/M4OM7SPpy4BuP5mArX5oZTH+iahUkou
qi3oPzOAeYG3NMkf7fE3g5yqxk/EzC6gwjxGHr0G54TYpg19oKvYG7QBfs0sy/yv
1WoFbJrOhazcGg7UCTMVaGSomQBDT1PHq4HkKX80JJxzmxThfpJhoL4OEFIC2kJj
9upck/Ml7tx0RqczOvlmstEupfLjqzApkPvEWAMJHOLns85c0dajdL9tyq7h6QZS
ume89q7GbVHNryd+XXE4J7X3/lfFIPaBSl4gMvQr2Fey6V0fIQ4PRb0MD2m2mvds
Flqf8w/7lDbx8/xByaTLqqCeyp4n9eteS96KicOb4QHRjBLJUxry1p6pZTq4EMX7
w65ZdyndR5GsIjm9NIKWmTt99cXJW9EzmVZ+DyzzE3dX5ROLHtmgLYKBkMnU05y6
O5qEEU18U8K4Qq2/ti7zIDQD5EjZakDsH7uybj/OFhHdxe3wIj/mZnMEW/kHcprO
lYUczM84YwUdwTOtMam+CfWlIFeEgBuvZqp+nQLwqDIYthWpT2kXiw6E2eX2Xss0
+PcKZoF+yWBQRwU4E94Lm79OyQ0IHJFxoiwAIAEM1NYEfLlQ2vMq/YG84DL+NMoa
A4sftT7+qyMmyUHt+KKnJQytSheWnjDrflKx/HV9q1R34/yM7wH3JGNNYq/cs4Xa
weSNnAbrBhdW8XKqy2hS1Hi+9uYU4RF4/rHTAV7XG7Ul6J8nnceWoesHsdBuD/LG
tL/jCEQcKsBB0OccDS0/diAB6ZOPvlZcxSEpqYOtKsKT20HY2BUsjZjyiH/G5MMi
zEVGlNz1eNJuccmJsvymnz6RGefyWAebr6rwmKVSYBFq6HJpW637y2k1AIXYo0/j
maoFQbWLcN9OD6YKhRbh6eoVZ9fyJE8JHMYeAS1OiUEW4RjFiZlX9B6we5+Rx4rC
3NrO7lCLa+TYCKpjBOiwGktMOq+1AWjR+o98sZ8YIaS698lCmQ3xItDDodZkl+WU
b8gWFDQ4uiin49MnSRY3qLUFVEykiErygVjbW0l0fRcfwrynhSXYav16wMwSqVw6
IKtTFKDLtFquUUnLH35RXLYwO0C9e7JdELylMAIvETCD5P/sKLAR0n2x1zqPgd8E
zkP4BrAsa9x9nkS9azxWfVBAnROSy1UMUQoF3SJvXoXpRZocqrpKMhEKbSkXZlzC
Lo1p1Res0/6uUvq4qtObTGovyHUTs+YQkXFS/fxJWrzNsMW6g20As2gxj4XyyhAK
rYYuvDb5SsU3M0Vk0wLcwPwuC/CLydplaiUXm3vAmJN+dQTQbQBhFxPZf6hPgD0p
MwAFAv/CFJ5kWt1jNySu6zKZnqGWhEzVmmVR48Z0BUe21XXeHiitoQ4olf+MyNUr
Pf49KNxp4fEQBfGDsQb0RWBQvblFUQ9pvA9MoCiDCIRPd7t+DX5GYNWLBKdd0Xit
mPNHuGTig94fIe4gIHAXLK4/UyzLyfJjhIcMoHSLNNVwXnQjqG0X6igWHfDoh8C3
HodLHD63+zJkcFSbsPpEsg8jEwifqbCkOtGQzOVTRMCRYq4cVX3lGvYGZiBkt9ra
J20OKBrfDFV6AH76ksO0ei5cVnPyw+OkELCHjLTqz1FgBaeWbZsHAkPPhZB/NZ1C
7pksggDQBgEyZA6+pjNH8AhHX+ODY9YGsBZPxxrvbHPOjeR4Pd9i2jCrCsO8+n4e
NVw5iJAbLAvmDwJyrPk/xVHcyGx0XsZhYkGhBo/95Ezrb/lM3gPu7VtgsYC44RAq
5k1l4nsm93+1JqmohEDC+Wq99VxAGZtPmj9YE5HfHnRPp+IvD6yH3avtybQleAYU
9tKL/nGUEbnrHuO6hxB7zfeoIkxrkEM1wSb/R8EvElJbi+pehhRSWg3Z+dghwy4v
Rva648GyP3Szs5RoWBMeAs7N2DYrJ+GtjADtUQNzTNLsE39l3SF89rJjjH3XPstp
hOHunshp/69Up6Ajc//nvMGzSQ0H7sF6SVj8d5XY0PGRDPh/gPzu/C6e25M1pEro
H9I1Fsb742SJxsVkZcUnM5L27M9bVTA3YjM1VOF5iYcgw+MaZP7EXiYzi8l/M+w7
MnZ9Lo+jXQk3+014P34FMD9ZysNYFR0sXYYxw/7EsrTJwbdYzH+/i32aiIFmL7nI
Zy9lT7NhNzwLNHynNLvzgcwBAStQedGOgUnvgCaWV1EjIi/x8hD6SiVMHU3mK0Ff
hXp2FnbsASn8T5jdDIE9qYFyXTqmeyIRugqMtNyZuMf1D92T7E5GY7lbEFMJrnpT
uaobzqfxEqLHgQ6YwhHAah7JLBd3L2I2iqcP5YMs7nPq9NWdDJcdBySplrStRYY6
zpCrryFgzOeYSxDjUp8tqbcz5lZeQlV5D3ImuExP9NDG9zzDX7S/Yk41E5JLkSav
PrYqiH31jhMe2zVHhOXDq/rYHQY0qyoF+CIdLT+8HIOVPnFtzHMdSdgvjPwPAXv1
04xFCB7zaLfW9aXqvU61gtk9cTECFV6asHM1S37sWHd2AD0uFLDBR3G2c0/v7jap
2PBG2QTPHeiHLl9pJik6KN+DWJJ2VYdFlMU8at3xC37crIB5RbSWqZ7tBn7se7Wp
NasZdFSwNU/whzQ2fRK0PObF2k8VS0Lo67Hm236Hhayesx1TKa9YR9Opxxh4zGK+
zVgoTbRInE3lY2CVBmiIBO8KE/An1DY9o5Kl3Qvt9lJJXnqeO8YporZgW+9HGGEv
O1rdNQlgW7ny4KSqOKcnNcz40FPfsKXSKhugZBmSOB6CmgSk7n3iS3+sGTG5JXF+
HG+2Wz2DghcwecQGRwhhauiliQR4lTcAahUQDtPUvobvNir9qwwG3I4MTQUz9/Ox
XczaXd3U6DSk8XeWgbR5oskCCqtTeHTcKkgtXqMgZ63xgGsYj6xV29ax43Wk1jNu
zbmAAwxbsjsX6py2h383DB0f8qDh0eXPBguWP8S9hYzaXDDGX4wGvpxmTCMWs5iW
QkdQwq0DEMmCS4+AE9fbQ6/L3y3lAvySJJD54ai90n+M7EqRGJ2uWxbCxCjGu+95
R4uminlsTeIi0fdBG+y4BohB7pzANe2ZtsZ8jxu0EvGtTWTSWSPT2h2bD9J3ZhLe
aVo9qt4DyrL6X0wUZh8TZUkyf1zVfFiC9tO1AQtUqyzPL/nsLVLvvrAs/eex+Qx4
8Ou8+maGCCA72thvROLq7Bw5kJvJiNKrAyrEfCIwlzHj8VbMSYCv2qRlk9KOaZwn
vmrGB5s3enmY3DyX5ntTf0cBvNHCbdLKkWem7Vx50+dQeYHPM0Hx0RQbSsImmGDO
xEDcwvaKu+e/geLwC5GUo8BUsZcF2Year0XmnOiuiRzzFgfbVg1o0DwK51+Xho9B
kujkbw6R6Ilc7bpJYKZa4zDUMo+8ZoNThm8E7ByIbE8AkpntiY+znt2FYtapck17
KAXg+RM29V0lhyNTlHWM6Vyn380a9BBwoA3SnyEsjyErFaDUJT2xl7PCxKxjUZRc
fCxHN1WwF6ieAJHlr25/HqTTqD5h2PPzzoOsjP9rV82cUKTTBLCtA8kLHUuWAGNK
r6B8Uky/utuJiUV50olg9gHev3WaF5WmKyjhtWKhMaCcrksBUkPVGBhqFxzGGZwI
BE2O5f+Pb62Z3CWUPEcvKuK8v6jcEqW6you6811AzH5VlAlElJG+6tX7yqetMllz
px+1NaMLaaTVw0ie6XHorXxT+NIFUwDUnTjb7Vc4BP+yBnBC9Ryt3JUgOG190Few
ASdALM7OZoYoHeVWEVtJ/d0PK4Q3szCWZBAfNl8BccUPSV7r3hXtziWTRgmhS/yf
Nw0w6d5HZ0Q4e4colUgr1/l5wunm/Twijtr8bs7CACbqVvbZSKOy2BC0iPVE/GI6
iiWYiGjCPHU+vVVPNeD1OW68vwLr0hjaKosWWyZbo0Xr7R9jv6ePbEg97r5OBwku
bFVbT9zWGaQ5AmTq/2pKTmMn6oi2u90x7DKalQwu0MwFPxcryMdSLFQ9nhuL5tSk
DCenIDCW73qxXc9Kxb02UiDYPSBNzMp3F8OxOjUfdE1K/2s6+nfamt9RQrtaFlr0
kkyVEDXzaTMAYjZcLs6kcJZ7OR9efUFUoWUcDVEO6eE61+C3SdFntT0St+OoYrgq
+t76es+AR6rWhHI/V1Agvf0aHo4YJAUCfYB0WQVDE51IY3q+MlyZ65Q56Oqo9VKx
7OGwlQT4cfqakGaNzOjLul96DwOvXM7jLkbmQRmmWZyqjdipJr2ZUxiPd71kYylU
mMOgtuU0A3K02soTP7Y7eFQB9RHkLnAF5N1EhF18A13K725xDBrvKQGT3g8ZWVA+
AnA5vCz42cA91v5U5WG2aXDXc+b8AmTVJ7u2sZDt5xH5nGpzLCgHQlLzysgtvZ7t
b9PmFeB7EiOcl8dtlg4y4n/4AAa0Hc1fzVDhNbuVlLIhwcdXre3JnJtoaCwkEsy+
E+/x7Y55doy1b6BIL+cur28y7lrP4vDpMrx5u6KAA7+h6bbXNfbn39aCThiM5WQf
Z2babKayFrsvlS4AgkwNY337VwIyF0q9VeOCzYLuZZr/AEPRG2Nvic5KRwyewL8j
LpfkfezWuNOoWKvDVXQiUDlHHSnaz+cw++8G853bWcVf8XaxjscbxI8e2EWWsVvh
gU7cdtVXyy4IKD+sKo/nYaahWL9aALz78UxH4dWJs+Y9DB8AmOUVnEMincjb32W1
W74zit6TzMdzWLmAdwrUKITyS0BZykBUFfhi3NWtDwzkC73l1A7ZNIRPZmr6hDjD
B40dP/Q97MypoYL998+kY4K1Vcxmq4l6vW3zdJ1HMs2lS166JbrO34NKn+2YdZwF
7fFdlPjYe4Ut35WfQiz56FdT/q/3cIDEilwVVZS95NE7AdU7wexg0lomwwfutLhv
DDAjI0ah2GLPjUSncM4TN5gV6fwNcEWHbPsDRIQMMN9gq76d+RkVJShoEq6ZR6QW
1DF8U+bgr8B7ameCo9YNfYFYxDpTP7w1TqOsWZiHV4lsv8H3m3XC8alseuE1eorB
onblQQv4NUOXlB46/lR09oVoAoOWJV3Sr/gg2KxoQ0jn4vnwLoz5YoVyRheAzUDj
Lu8DOtr2TV2YYMdiCDf7+pXf7KLGaQIY+nNnTwcphiScfTt73E4x+K11QJ0IC2uF
mBwauPL3CHYZ/5PEjW4qP+/asplG8D9E2xGGICsknf2h896Q5GOsX03bSRpJ5QM/
R7EVyprJomHcnFlM1FL9T0S+gf7HJJAN6qksPA8+XmwljSjhSshx+0ivIVPVGXp4
KXw0ViFVrcrEvldpiVPhr3BXCRl6/twW0QPFUotZEdL39DwUzXWYJ0pmtpv1qUNe
CxtOSzY3BI2iPvgjzzeqTJNPBhur0WTp+XstE23QxjjP8lQFFEdJ1x8fH5CXEQTO
cxCFZHGyLQ04avlcm0COgQDT0Ff2cnNXMLpINNE8sbk7ILajClcvzGYa+Jj8Eh/Y
cRQIMH3vYQ2lWjkfsQp8tQ2CnlXQSwsj6BptBKOSaqo+8hHvEdCUlQckVOtZm4uL
5HGFiDJt1eE8ldrc14LElmbgLfbZ7PJOFR2B6dEHa2bsaUzkLyAXEmyUS+w45D1V
lAIlGsxwokq8+P+dH8awVvkzEb02eWh+DnFImv30oAuQ7dSKsILBOLmqRevIgM7y
mfaXJQKw17m+ztjjsQSVF24JB8RVrN0J1IovOyajhKm5aJK2R0EaZtO+bripVaXk
gtcE1ELKq36JBpdQ5NQfgXpK4pxoIXA7m6AQD8cY4xhhdF0Wde6oLW8EFj7ZIGDF
gTZ+D+6jYXBJXMducr3aLng8qEWggLjrWo4iGLEgGf8KIrk2UGVzGc9BQmd6+Zsx
Wi3JF5IiFauNcb+p4jwZOKaM5HBtBqDyJCJ7HB5AFcEMQJUOXpIJfte20HN4P9e/
qnONUL/vLTVP4KFBVkxp+erCwD/04Td1JhyNLE+ShQ16B/r146P83NPPLZt/1315
U4c7PrvbH2qAYRUlFZD0jJIbuQb4RBgz23FSQ24Z3+GjHg6yntGLqTyLUvf4bkp2
hA/65xWhJ0NYGQE599sPWkexRBDvW+ifZwUcuP0keSHv3N4r/GoGaeMYekQazg57
MkgPOlrOIzFnoRv6CPFeea9qho5IrE0HCLhTd7VqJrRL0pAV90+yUUcLYh/3jddn
VCtoVwts/HFAz+l2lEIAPV02PTTX7UzX39WFfNTuCEGP2iBU/qAopfTHj73iAznQ
X3WT21nD+LZWQe4CCbwbcDLZsSzwnDg4YVhECpmRz15FcNOc24jsfo9rrcCHMJgQ
+JuKMcQKgdFj0VKNuef8EsysMRNgLHeeu/Lh0sx0D5y36jAjc5ia+QCjgODPUzgQ
9Jjn1SX24hrTq4iegwLblHjSaNrrrnK3f9Zsj7llOIun1XIsCWfDfWrQ0sF4MrMo
h4nfeMVJpfwpv0LWANlgKZ8MsD3qE5Af8Z2Lhzl9ySis1x9KkXk3ry5MlyE0rski
eI0dO6rHfXFgCJ7knIUUvmxrSXFKiQnZsbJ4/61Ln3eVolv7H1NcXmG04lWJyRUz
lgVthbTh6GmWR2oMQi1rJfRz5nSVJGptuytWFFFR7TnGZaaBgl3NUBT/Y9qONzn7
aq7OC6F1fVgMCi0OrRecx804I5dtTdShy3ZWcI3Ie7dYSvG5NlgrDse9znpHdiRI
HucEqqc/bhO5LddB8dCy8cBRaW+oatTwMo+tDtnStuGobYA3HX4+m6s4lI74liVZ
jeCBnXr0NYz+Mm1OhCi6N221x7SeOLcXKWGM6feTQRLERGdq1weokQxb/wyib86K
uQ0fI407U+1aXcmVLYMTohU8NyPQTB+CEZK6lFaIKJzzDFC4ap1R3ejvvPPTWe/b
TFKma0Df7aILLBiZb1lpJwovG/g2B68BxrcQ07tGJ8GmtC01NAiRhnFALjxSX0o+
lSPshNdZcP8QopFZEg60GLv12s0LlOVos1XL0dUGdZcbuRpQqMuv7ZrgQQSYwcWC
px+0JJD6q9Q1I0PcfuSCJU+ir8Nqke1xjKK5K/wdHtaeiHA+pVZc4QJLWLwPuuKl
eWmEbZ8IzBtGyljdmYeggCARjdOD+B6E3B6t9bZRiDp8p2og2d9k9Gl4pmSm7MG3
2fm5hqjaa6FjpU+6N+1SWmaokWg81imauATQXp35fh+lIDhITlKqJpOjBladQCK/
Sik4DO+GzDqMZI1W3ghkFU2Yf0WVD94tp58OokTCXF/NM1ukVkkYsPL0pr/IId/3
ZzspS/8jJx5rCdFNZ4ua61bMXXx2IZpdOeiEjA8XoXerGuvIwIzunrKTWE3DTFU3
I5wXEF55JkBWQ50lv8p+vxywKrqc1pLm0uJxYMNDpQu6Eroi5qedabX58V/NGBA6
z9d/72j1fd2nil42LfGzYYslOwGJ7Tm+ZmBJiB3voNeROpZhJhL4bVTbtNwuy6hf
OmbSpvGIfK9pGmVjUJut/Xc01kJJYfdayyDp811NheV+pCpB+6XvyYLUcG1QT9x3
H7OvfwlNnTd6Dl1IsKvJdmDxk11/KI9ppkncgdaWspY0piBF3udVCaZO4oOEPHGF
R0P8vDgh9rRdglo3lFq/3eJ++Z+ofHD+fSD/OpxfG5V5MH9OK7TvH0HL5Wy1H5n1
YbjiF58/MdxTM9A+NJQPrBJGxyTyU3pVaCnSr1enZ+CKmTtWquxvTaC01H9cgOiG
OxXwDpbJySDF5FjvmRvKnmA2s2dZq3D9a+BL8ml18Jq0ZTjuu8qn9zOE7czWEGOZ
edxdMdE03TCGa3jxgcbVOx7PG+2pkC2leBswPDFwBYptUEfoVHZkDN7Mu4Dwi/qU
zxVjebCLGkNub1cddQ6MH6batit6iiHaEYPtGXZ/E3+5i16maW6zcn2X430XUC87
un9UIV1gtQrnxJMTKt4/6VLYo+kT056Q6DVQJhoQvGglBVI/xTUEqPLvDX7stQCN
lB0WRusnkN8Gmg+Ik0NX0QaApGq5YGDYQf1wOBx7OCDhv8t7t0APoaPAgCIsLtfF
FPOHYPmTsSuxhBgKNMNfM87jKhj6JlaneY4POXbzUpMDf+BYWe7Or3s4/0Qlgyoy
wdsYhfBauyTdy8tGGetygn7ooXnt/XIOC/BOsL4L+yIf9/wpTLUI6BWtXogVTtkd
irssm2Yng3cQlsdKF57ENOIPPkvwQzfdY2IPM/GfB4NViu7NvJVf+FV9T9pNZeJc
gZgq48p+ctvoxRJ1h6xF9wT2RM8tYCXK5zZ0PC1zzcGz3ODzYT6eaXYy37UZZ4k+
f+bdWqHIzRK+J2IphhFvHf6GLRFi2KRbvB4z5B3eul6Zq8WIMBnEs8qqaMrcobIg
VwMRvR7LHUnzf/zNjbB1I0O8gBlkHvnVlu6Exjt4mYVk+Coi4ahZLoDviGrk2Epf
Dv/O0v9y/dnwrbdSQ2iX4kME8aeef5e+F+USoEIBm7QC+Fpgos5vL6dvaImnU6it
GoQl8rTwwHkwiaOXNmF6P+njwy/nt2dejhN0j1zDRNFPLxHRJoJMtUyDORJSsJSU
TQXz8Gkf7YZGMBVNb0wk/6nqw164Ct4Y/QpFpyNs/Keq5jgiz9HH6FK/XenNb/K2
zNXf1OR1jyaikQUbnHWbyy0aZxoyAXUKMY2kehi4JuHArecmMVr2GOaGlJ+lg9lO
gSB1imZFZOkIhXDgqxuorTpN/Jnd98KA11xY0sYkPxZiZLYPj3Jv+/A3sGbKQNz6
zVTw8SavDE47yPeP+Zam5DYqkF9GZosHQXRZESzrNzQ2yZxBySC2q7bmEOVN8Tz8
TNgA8TepGdvK27O7RJ0rojN0BsELfjjD+2K4czNgnDq9WTnqFkIVl3JaEoTEpjYe
92xeG7XdqrGBjvoTWfi7N8Zoqleq2duLyNls5mEXnsZb4XaTI/4mzKuDCyiJYKWG
Tb30FceZIBIQOZnS4LJPCFhWrAvEEwaBTOAIb+6U6tklg+L/tZfGtV3YwdRBc1Kg
1rv70lJABn2+VrzbByFvXnIReYngimROtDzPNI9ps1JKRIzYNRJupalEQf9jKS67
0ca5OHpW3Fh4IREgEVkKa3QSFbFBonaaCwtxJSWrigjsjVk63wJgsbEqeChEnl3o
wMFzHuHWyB9n+ANB9t7zX65I+kKt9EMLQcItSj2LbogR7NN3V8C/QEAoc4SR2D9F
5i7H6M+Jb9/A7mU6ITG07UOJsNUdxcrbkofZu4of0g14eIhQPsDhFrYxF41FOO8l
50Au+mjtV36BAFEPiEgJrEckCReJH/Zm9LK2Zqknmgxvm6UOgriF/uKLEn3eeE6I
P+PkaiT3yXHcQmzatXIGBWMbRvGnfSW7fQUq2JsDf72LRnsY88Edec1fzDEqqsUF
rlBI76I/Y5xJmojNKdSvv6U9fR19a8xTJLTEhW2V3CQucLyNnCCgVV8UiYKIA1HA
acK72EvI02C2gEonURQHkSsJRk7R6WZlb9q0f8OmjHvEPpxjV4E/9rgrWitMDy0n
1nXVQ46Yq1YyF9Zrnbp/stU65I2g/wGqjIYJDuwofewdaSlWTNc6pdQKgtOkuS0b
E87f/ES+YIkpWYgavM/T3O2UujGz8/5jvKt09SbHDQAeNFhad1oB3NXavsXu7EKj
NjF4myqa6VKPz4UeFeVlCqs1+0VS3HG1IYH6aBwldJwFRA/d+wUSnDIalU/xU0xq
oFD53FTwTVG6NtMzSX1nIgBBcuZlVSdNEj/FHrsDHq2+L67kNrGN4CQ274QmnqNk
2wNl378hUzvZipK+TaulF2kZ1R/RdIrGgCGXZez4jAj6KPgW634HDOJXM1q62OsA
Ki5E65XPRxAvrdv4XJ4LEphQZPBwhrTeYPwoVYbUzUPQWvI9mc+Rv2TXT/mMS+eu
1BkEAVbYcHwxt8hrOEtGm/MBe4WySexawHtIWhbf4UgvvxDR3GRm1ZPDZloZJmmu
BeRmAITAKeczwHsnWzox4BXgP2A+kP5T7IcNYpKrBpJx0jpNWSrnNxz4xg2fT3AH
wliDNvSV8M3gY3Bd6qkx5dW0JwABE97WMnifDG/n/F5RP8Xpt250HWlDLgEXIXPw
HqiwDY9rFAbVNsRaADVsS9zocRTwk1POepApRBUAAAC0rbbago9ZeepHIOTO0OD8
OUW8VgFLxnZCIuzEhesdN7WMEK7jivYk8gSvtIFVr4Wqz4vhEp/dDfFwXdiUcp3I
5loflrIUHiAw3S9nwfUVQ3kF7I3QNlkeTvTb4VVQ7spa8p+1rkPtZ8clIsqd1RI6
w7nsNU+MrZyoH6BrnxP19yuj1LKIbFriXepRX6nm1mD2lakaCodiuXbrt7s+DXHF
FAw/i4q2KUSgi/j7hXHJf3zzynfOA/Ho4HCGxlJulOsiuI7KBau8a2cypbd5Mlzb
yNWWjrRgLfwlSfwkfgcEck+tOllY726ImazciVfcA6lagpDQ6pSc4yp4Wvuxo464
QMTwPCJ+MuWoB173KXXSVluhF2YgzI9BTICH6qEeN2gCps8WJMyTqmYLBSzgupZP
vHiZ8fBhXk/0QBHVtMCwnCTmzMGfuQpFLX/WcQLduUfo1o795q8PC4+ar2YO7HnQ
wBSC16/5olAIAvRwCZfFlTWMxf1PqUwo6eyeWGM2hp1m5AnN7HkVhc69bZZA7hOa
HTorddLJz9uvf0INpgB+rXeZ3QxuvOmE+EWAE1IyDSKD/VxKIibA8sNvK+JzpRfu
sf9glxNJmtI9VV5JVxfZE+aC4s8rZaDFh17J/k0ESCW9ecQeQj6nOWTnDdejvv2k
0e0UDtTdOO7KFEZA/uYEzgFm+1THi0jGPJx05GFH+nkBrxkhlustyg8Rk9Bi5txQ
8bnEvCK7HPDKTGQztFMLI95G584j0Wwo9sI/7YV1R3BaDA4TFBFNK9/0SxSLG1Wy
Jz3fcUwQ9q2p9SOePNrQUj2VFLMXecViSs0GJISUs0rVrPtGXk3WtljcvXk8wYKf
UCQuojM+ERgLIup4VPj3vaIYexe+CCbmfAGFHa4JG9WWtRfpiVzZ2FOhP3xQ+PMm
FTqdak/4aYTx2F6sGQjAYxS129ZeDe+uxlCrYssrhjVFzmJFTS1IdDlfVZZbwIlI
DJJOfU6yg1jswHvf5OwVyQ1lgx7QXXSzL6+sSH0BADiQjW+lfFsUvFauA9ZbQLZf
4eUUUG8XN6NBrxW4txRI9CKdKdlcgD82+Ojr58OyCvo03rKTJcSLQWO5lCxyv9gH
ilT4y+tx3DCF4iHpfUT4aI/K6AzQVNKxZUhMn4vIZuiJV9tdeMpQUy6YiAn3udhy
2pCCOTq+CTZxfRtmlT1Qyo8dcZ1SRVEUHJIQd6J8Ugc6hwDiOBW8tkF5hJolfXlv
VBnkF6+rfoniyy0yI6hFmxPisTn4Lii/CCsTnH0wDrwJAtpU/QFkF17IWlL9mMBt
KwWjaiK+Nc1kWSSFFplYtxvu3vD4F7LP7RW8V8lbjsYKVAruQN43cROb3/se4qNm
X6E4LizQoga37gZbiMvDsC0OQV2j7Opd7yJprCCgt9nHEmAbK6BUk7v1+ts11iCK
VazObDs0Oy17Ra273eoXwM059cQVkuPgzk1qQIVpdfXF7k43p0b9P15bDaRfUMyv
tL8AvDifWDkLfFVBBzeHWRKF8qmxKuNUlgj1YVh/aRn1GZkc4ancZgZnHpmV1hnh
yR6nT5fbFIECYi8GJsFNMkgiLxvSN5c7Qizw7QxY+TA5Ma+1Dcheul7DnZK8asCR
fWsQ5Qwg611fb8YnqSnKRKoETOVSgORBHyTJ/3tGGCZyBDCwH9UeMjFd7UyvZqFL
au93wPjCOFBZ9FH3F1+nAsv9RGtwg2jopvcKF6z9WKr4PKEy7DfaUrtn954PwHjP
TwhfPLubscbtfQHgAxuGTyy5RbL/S7haBBLY1ymCau8CU2xgPcg4tQXESo7c05a9
OonBaJyfiwCPOMGLm1440jTE78iKD71X7svYWjfA6cfppDGZEx9WJP7Qh4n9TzMj
7NzwipDohCuoogLV2UCq+dVq7uMMT2s5aRy2If6glHj3W5doDUSDljwYqmnOQYS5
C9QVx/jpWMoDBC4oi1jI025Adq9eE5DUCkcg1ROAOj0ZntTo9JlG7KQ8uyj+oU4+
ghEeg0tLkZCeWzkzKtpVPJ00d81h925fisPzgxe/UpITJlr1xPVSOeOtJ1VHPKL1
cCDsV3oHOR4vAABq9IyGRitWT9AaHoH0oz9kbOhqBCM/gGJs86ogEFLqEKT0rAaj
nd96JHwx1amCi6EuOEZq5rL9gv7Dy4Ev5EiWr0lhrA+fdJsspXKPFAeuMTif5AEx
UlkZAbYfFaK4ip/5/z87ytKN1GY7V/1BM0h9qb40WVJ7ViVVDOB/90gcC6MXCIH4
APs0tma5Ii5qGVgH9YlIzUZhOKd2h4/LQTJVgP82k0Ud1WXAee4UBgb6yHif8fB1
dlR6uMJQybPXb0uwWI0FI937iT++l/GDYrqv4i6qTreqkIIrE4OxS6hBHl6JsXF2
GiHGciEa0xwN77UVXEsnANOCtzHFs8BpPuhTlLkxR3MrJC4+vfP2F9aWuTnPwq+f
Gwlk6UEXrCNKwoPRkVZm3KeX5kU04v+/Tm22+ImthncC+IaR1pYDakPAi3ntagxt
qLrSKQygNqw/J2ztGZsKjKFtHe7n86v0mJaHV3NbHfvd4gmRilS91yHE7wrVbRNk
VpvoCA/s8Rm0GM0TcLVS8j/w1EdAGuvkK/b/1uZgduIHyD+7IBIaquBk1EWBOQck
pElgvgKRyaMPGgfKiVW8HsLpg9Os0ClBkEObpR4yrCZtF+HwkKlAsRT60g/EKHpr
bf/BwXEKPOul3vRmFbZXyvRYFgObn7T32LoApTa+O8Bb4g1YZajEA9165OqQSQtE
vrQGRtlnwP21DYNZ9/weh2QMDBKELzJHPd5CK8jhX7v24GtgLZArmms6vey+mUXp
mX27JWfWXvdagm+QJwi88lWpdQFwZTgqiT2F4EvLWa6Qsth66BsL3GCUUOOUED2I
JEiMLdKZoG6zBiFiawXB7kvEjXGAsT5KJibXgGzuDqWBjVRvLNMwBrdUJK+d3vnd
X1PiGlpqK9uUGZruceDHphTLZq56H0IaTsllWetQLAYwt3CdTTCf9wlGuNUu5qQQ
S3zpoWFVgzU7xZIlVgRKXloVVHbeSUCP3iHa/3OVHOPa2542WkIh98shqpglHu44
vA61730DHQ1hOonpWTh0nRgJNgDandldt9ov+HhUyxf4eIPAguDApL58aFGfMHra
jrw0AnHJcZ2M19Fooj0E7HT6oV8bHMY+YNqeb5MxXAHQqVUnPxsFcZrAxlc/yb/M
ynyEef9jpdIBxa1oN9tpq7ZFptuviwUyDsy4wcu2FL58Zv9qL995lg5VEp2QduGy
j877xAAtFOF94Ge1zWsALeNoEX3a36EPfQFJLAdBN9zCwT2R7f4yl6s0wQGdceXB
jsXtKuM84smFPSwBTVZXWoSUxO4TBaL1TWRfqe1KgqFf0QvUJh7cQ7bli89BaVkl
ualbsGctc1O5JEfWXwe2laqUky3O21C/wS9N3ZkWsGpjD/a1MkOmJ9WFYNJlFG4R
dsLj+S4y1LGbvIMPkRHBxhIP9Xj1M7G72xdf90y6Ngw0cu2Va9oPc5qgBeeMOCPI
bRVx1JU0xZiZPC8yo6KMMkYiw53A+uxYTj00MO7oTMKULRfxvOsU856mN+qAhUEf
WGbBMHmmBGHcZMY3MB8/FJWuO84ThPRqKu77QlbTlTOWa1tDL/pZBfq6O08AakKq
XKbJO8Z2T9xCXk8mpAzZZvv7X/cmnoF4xVaH1f2gZMtlBNCC71vRt4nWZU0by9hx
b2TVrB0CNfS8O5kj48Roo8tcY68Cuh+B/Y4ya63JSxbuKBfBOpD8AW5lFVQBEKXh
KgZkuQ0rcKiGpHFJnWry5by7vOVjg2rAYw70XCz7r5Xdv28+wbiGOc6NCRW+g+ub
PExelsUnDoe2p3up1SvSBuW+hEZ0pdYLve930yAwA3Ucq0H5uhUxrSMh+kPTh6U+
IqsCBhbAAQPX3iVti5J8g+ieeuWnta9kBb3qXQkZZXvTHR760a9DeUmH03wJk8uK
m6Lv/oDDjN+9JPfIiaNPWwb6YmKeRp/LdQ3RANurKlVqvxBz0byVjIFEbmB01rW4
Di01go0L9njKmwbuNxsyy7l/v89CbgX1BdKtTKjs0oZOypb7BihL9pmq3FdDSb4k
i46NjC3i4Y32pzd9VpDkO7KNfGSyOUAgmoV19UG/g8+2KiMPMfoI49yh+Aw0pD8u
Kh9gA+sHx1us+jDNvGOQe9Vx0rPlCtkELuxTlU4eKuPOG+Su7rCLTCZfdnswWn1K
UUpH/RwtOODbZxOchumBeD6PogQZtAHZrlzuti645tkbdJFzf+qeOvRuXAHV7fs6
lC6kOzPiXT6mJiZSMUsnUSnXasElA+FxQfgBdNEQLL7hgZ08ACaOgFawad6FANbm
SRRLMFEPiAI6q41MJ61pJvp3fdO5RpxB6FhqeXhABDAkdWPnc0SU/jPdjbzd6Uhr
LjIDk+2pvrL+Yq1JGkvbX74bDkaeILBKOfAAwPNPVHpVURid5EguAZiWdMqvIVib
/WhAGCIDVvDn7bupVmYOa4GJvEjzCauGLGYEyZs5gyrbUasmAnnuEPQYk4HIErqZ
54MXT3G9mim+8oUZ7LhmhA8UmFQkfBQNejm4hE0UtPoOEyzhwNkx+9yegpxputxG
8wWpkYCNMaVb8lhWTTbNXJ/tg+hDtb7LHBFqzst9vplcLyeO4C7iu3nug8RsdIrt
bZthG4jAOd4SLxfhmAW2G9QVIKtw2v8toVEwtH0ITgbF3p5l7sslmmf7VtsrhhdH
SJfxtWEymJ89mBdlBwkcAjceDM3KZTEJWWoRqUVbDpLVpp6mizufGPu6FoMc1MAW
fix1bdysIEwUe4TE9+lNsmqSwYI1ebiXQJEZZz/D0I3ctu3HaCD0wfFjaIBezP3h
/5nR7HPhc5oFTbeZvy6rDZxSN4tNJrGQHf3rjyllRuwdV8wtgUl7Si4hOdaX0q15
R7Z37RU2z0xamOxLDoygwm2+qheISc/Q+q+Ah4unPUOvqyimOERzRPS2gQpml9N0
inPw1JChpRrfqjTcvrY+N/WSaj+ZE8uYVkOIZxJ3R8l3TFkDhvR1p7w9gCypWW2A
JI6uaWAs+1y4IlJXLADy67t3B7TXHgV9jTx7D2tQIf+JG3cByJG81BL+t0a4SF9n
vvKBYymQvE7lkQ2xsoGLPV6fUgx4iuG1jsLvH/h12rx1EQcgZdOQMPNMCUuP0rS3
O0JK9roPHJwZnBlrjImSoPrEDAzgCK4Tw9QzUZA5Ch6UgeKvgaaqf5m9K6mYGipC
k/ZaFgzaaj0pD9xTQe4A0wzPwXo37KyIBvqbzQEdbgv9coID+dGqZmkijLUBeDmf
lUlLJOOTYJOn5Lyy6geuI9SSlK9BuDc0SAG4vG0L9QMMXSLe0jLQlmHOoeVm3hv3
nX9QoavVZRuEaVsBc6aack4OLhjLjdtEkkKw/Zqu+EmZ0kZf1TZbUqit2tbtWv3+
fXJtviNBLyg3bFoDay8MTmLZfEhW1bspluPHHJBJu5IWfBxM7wAJC9QO8vFeUgxM
w8aIpwu0Q8nVOQE6T2zk2poA+uOYr8EkhIo9e1NrxwcpC3K285HrBPIb+9Z8nfjH
VnLAlCLjFbgBItJ5WNc3Nifcg0W5rK38pqe/DwOMOSiU+pE3N7zhweeVFSdwjnlx
iE9bMcWasp0vh0Mwkiu4GU9bnGDtShnbSQ6C3D9YCmlLm5RalsFzmqv1TVFdfgMu
CnFNr3u9YcdsrnCsBJyKXuEfFmMNI5Y5n12Q0h9NOmJ9DL1qD3PME1pniZnF6hKY
zcU+l1C+KF9PDSv9ytrwjQTvvQS4QcsLPFpYmDl+9i7nLFpIel1yxW32rDfn4Vwo
r55vzO4zrgZEBvXFTpkXR+OtOSi7kW/vehPJVHysG361FZfU4ABtdbNTZlAE6kq7
uhlpBE5K6/bjKe4aN1mtW7yumWPFVO+SxqewXKkRpezBfsIDMDfJ3Y7T0CyBwYj2
j4jNDtR2Y/FxRtX3wNcP08SdbbgUOHl/bhwQ78eZmM8M26rMie8MzUbNJwELzQbi
D3cHHTW8NJN/JgL4wDlnwMQgtnXzt18fONWBU087E2uyhkVvzbrGNOcGKk3wh8Nw
Xi/ZxAVyMwgNHfSorqGlM/NjYouy+EAmE2cucE+tRRt27KEbQEkjP0zG/p+zvc2/
p7PimXITjDnGVPwRsMluLBgxm1FM5eeXcGz/hxoOqGzcHre/aR2vhu7dp76Fg2Pc
4mKK6h69u7hbRWfmsqAlyQFxvV1BNpuzD2sPtGLHv5FfzPw34ngmxa9szPPmS12p
B1/O0glnsecgg3DO2gtrgLID75jcPH3kyQoS+Or9wd5kp/cBg4cFmo7OnlP2L9zp
k5w5S3m3odbTpaPx8QE09Ia7l6K+S0q1HPRk3qDsJDdf7EWgd07EiK59RjSv4xf2
XteCL+TyFENqe+hrgyNny+o98/4QtjJHiq68tXT50B58WBKkvSoHvuDEaXqDLqhR
cjpCVYB3JzfNFxMArm6+JnpCdqp0mPGLhtzSmijUVzhJwv1+4MtG2XMwvotxzY49
dTWJplQrBrqYKtLXxLWfKxJFcadgMDMTA+CHZtrV1Nv23STE50kdHXOwIqkirh0R
NQyMlgv8IH/hdn7WUQfNAHNOOvzscTtKaGS7tA1gWF+xuDgy3HuF3U09E2dsIn0K
P9sbL94VWxIpx3upn428N1HiP/rQvMHTuNGFCdUZziRipMes9KZCuDRX9STzz42u
ORrFyoNwFQS6VPFXeu88ammawCC2MZrPkGj5ndFHceEXTGW/ETIi16aHcQRPYuHI
MCeqBxivIvEmvCwN9xaTlQyaVZRA8z1CaTZ04QWRuIkTAiOBZKr4p6wk3IUi7AC5
JjGl4wABIB/qF192cuSENnPnajUfsB9L0a/5pRHUv1fF9iG2UCDZQWjsokI1gAFO
9TDUtK6mc8U8tksgACTUvdyo84ZuOnwqTKe+WQ+4vY/ADoNQaqUVmcfx1uDVim+l
ZxjJGLISbTC2nrhoVXLu9nVv13zYERIDGq5qihMu+IzmZDE92VTQ4JjDEZux10aN
wPW1YHl6UiV/u/NItsDGksabpFd0Re6WuMgGMNmp050WECf8cHe192ZV6d3gJBwM
q6hL0WxmX7Tr65bzPoBC56DdDAAU+nDhvhMRIKGunNoUlxw7l0Uok0nMPf8ghG5s
tOlVJx+Lx/zyoOVMJZxgI5Nyxsc4txjTT00H0Qh6/w+q6KmwE5Rfl/fuyrNuZDtZ
8oX1tAeuDb7jLaRGaHa//yXVIH7Fq9xxnjgmCT7MC3K5bBer8Xs51Vo96L3G273m
Kb5kX1FUfnFjvyXmjkJtoyrR7kGEZquuNjzyJjdPijksCr1/6EYjFi8gbWx9Sztt
BxbX5822uyXB6hPLM7J/oLMZSLpea/iCFEPgwK4nM0KZ1FCmRiZdsGY5f75KotDm
UQmpjXPlXyWMoMywiiyVmE0s69jJdNF18TqLRUhIDF/FTiBK1qFThzSar/SEXDVW
4CS8dEZ8ehkd4CrjWTO2FWa1ceL9pNFUPxlsiMr/4IM7KxqhEbhYFflJKtsG4y+6
kVNLxbY7vtLNTLE6yp/AWGytfdUtnisYX3rI73EyTbk3fMnOeDYG5nlr/bfbfBkc
0XiGu12Iz/RRwEyLqZeflKBQIVjQ1ggrfW9DPa1jtFG5O4oGcNjAX/ZQVZ81XSE/
2hc5e7SZpPr5FzaMOq/ltiGkhIm7YPPSX3JbvZEk1CjKBMR30Uzd/8a/puIRn5wO
AjLQ40uKujf3uPPbrbxhsWLPn0VQOkf6HHEGjf8JuiJqWnlu7zBKHZX+C+Z5E4jw
nRSXegQmZFEZMeYsv8cIZLZhn46b195vy6DFHdE4Ac9j0fMwDMqFcevp8ELwFzi5
a+oiVKchleFYuhphjKdKwCjca0i4Hl+QzrJ5cVWgJ4s3z8R/6NJo9GQ5d7lBeYyG
5lYP82Ouwn2qVttQwoQwoH43jpiT+onWcy9EdqCimOsZb9cDs6PMye2rcGLynZA5
m5kAiVqchyRGWroQhAmWgn9j7KzbU5mgSIqmPIcktXpDz62MNK7ZBv5UdBKvmUJk
7ulkMIE3Pe22dtgFQ1flgNuMpZDCWywgbe7spKvBf1ZsGx/NKhB7Cp3q55xUDzzR
vtgSwBPeOt9La6cLWSCcY+9k3RzoaGkJNMPOQcpjUZ9891nuqyDSL7WiQ/ySAONO
xDqtG3g34SGr+mTlNVAmfVoJmOxykMBbOJ9SFl1roWaf5ELbZresW1AeHazLM66n
t84Kbx6+xsrM6rtS5VB8RNqf1Wp232f/Ywcyti0mDXHLbg13vM+LMjzoc74lEmIZ
Swh9JyxB/+lBuNw/I1kk//OjqSP4PZleBddeG7q0XHCrZbd9b4+NzRLTcVWi39X5
I1xvQk2SBLQ1MGXSMDhlHCSP4Hvu36nfFhwIk1tP2YBe5OpH9oD50joFZ9sKTJ4e
EARFJSKGpDsu8KaQt/ezfxu73YygOVc0mPA54zXmTY2b45hSy8BULW9AM6XE1QVB
gmK31WWwaAW6o878WfeO/dDLp4SV2Ff3NuwZC+QAo7XCmsqh6hKCTXL2iwCrvKb3
4IYskJJwMvg/O1VE+xJ2T/ZGLZ2P39Hzw6QDn3Tc0Vione4PpSCYhs92EAxxEAnX
06+2mFgCAiQYiA3gux2y160GwpA/kqubNrzqv+vcsri+cTlJzehjV7X+xg14nrEH
byuJeBzq/YqX0G/9wwT2BL+VuRbDTQIfnkMLws0e62JS57dsSWSrw8F0p9tXyjnn
ovvFChhb5gAvKVXCPbQNiKxrl7Yr2ohYnMH31Dgu7wDmLHM+ebE+hrqb1pu/TeLC
9Tk8ziYYwaHd1fergkL7+RrXa0kHANz79TwxritFRkNcMhCmHS6TrlSem9fmrIXI
aJ6ZIAb7LC0jl1yTQgOS7i4IkLtvsp/rRlm6+f1YB8CVbAJUSlrexv33nXIuWqYn
wtPsDro3TzE6eeoymIRt8z3bNmGacf0sTnj78iWxItqLUQm9RgwhfFx56HXmu5AZ
+SJ2b16E16OdeA5S2GRibK5n2H4weDg5WmTodeBkdsPXOxzkjPi30S6Nt53JHPN4
1iftAyF1cJdFDATS4MDnM6O6hfUB4FByB1Cu20DdobI34MjZW+od9tF0JJCAjV5K
cZFvehNwWF+2k8U4OrHqOKKfkPaRD/XM8E0g1evGecixYNdOBlW36gr8Y+imPdAb
yRNelq51mop6tSq3fMiWOw8w/KPjTghiGl5a9MjSPipEDIY1+Y71fpZaLVmCdSvw
9nNj6SEszSnkQx6uT+80ELG9zUDRFKp6IQWijsnNaOM8WkeTzR91RuRL/vnzqyhf
bWGNDzHpoujyvrzWKVwvf0G57fDhtIRXVB1FdQAa9rLRinQZsdzA8GKkebvqLsIu
TXtbEzCW/dQfSl/W/TI5FxYMA/S2cbYWGurGvCvsIVIPm3y78ctUy09NCoLsCWAX
4gA9z1twFIaxnGIgEXj7VOrJxwTOQ7up2yNNnyqPx/plPtjVmtKb3F553/RZEBvt
6Lsmqjq9RJOV+uzBr1BSbp/CBtuZwP66EGDGtJoftyf/U5p+F3x81tXB6Msg4kFF
+f0JAEomZSGrwhEq+PbgQbliDAO0FpHxa4R3e0xj95xwzBvg0DVtNnMPuxW4AtQ2
xhkK8T1hD7CbUIZ70yXc4JHQD44jOd+hRZU3M6eW2lfaINXfj3imB8xRAim6JxVC
S9lG+VqzsooIIlfQrdhp+nEm+3D7d1WhVCzQXZhxDQQKsNYJOSnn7fLXhHNGAAOT
RSjB5FKaHQyKv4tnD26q17VpDBsRIw6iR2qkmh3yw0NZJaXXEo3rMwnXCwyih6tB
RXjPhfUXAZa0wCKikTAdO6uTE5qP0Tf8tq4rUEL6OeYxKzZnEZpax9tPbIUfsUCg
cEet7qc/ebxkakBzFXfkU4QqG7NZXDKbOTctwJkAftK18FbfVc1RV8YR31GdhaGn
hKbK8jCFsN1ogDR9Zqkb9Z0d1xWGBS/kkBg1JB0GOec18zlsyuj+1c5lQ7GAHiEl
9uwONGt2ewqw/rtuwGOOzmbCotJ3lzHCOWDFTnn0LW/QFNvrjfpbPTmsH7eedEjS
8YAX0C7tMOrHrVCw9s+4+GmwL08UFOxu+stSkv/1OHTP483hG2lLYiVxo2kXDHqq
PEtO/3NHSsLG5MoEEF/I5uR3gIUL130aZ+pTue6cbXyc8I+RN9TEEOXdJPuScWPD
N+Do4Oa50EnI7PtooxZidn/mr46Vw6Qoer6FKvLjrI9rFIimGOuz1a4zrX2OuUNo
3RAtHN3M06n6IT3pai60eq+l035MtwGm34n0qj3pnl5VGhyp6lAwWV6vPvxhe8gM
RPRUW8XBcxnAbnFTtKRr7SI9I/rcyru/4KrV47WgUf+tERrpbRYO5+Us51EtcFaj
W5B7yvWaBkXwH/YhxWks2iEcs1K0kWG/OwOnVKfXbsdf6UI355hG8Khzcnt6Q8S6
9DjCydz01vzzvKQOCFs3Lz5bRqxr41U/VnYV5y3To7ADdJsk+ueGiiJ80MUMlutR
PsKcMyIiRsHChxV9fpOmaHI9IbHghyjYrc/Wmu1OLE6RplDk9kA65/TD8xepRaR+
HaKDpTXkKn6z8No6EwAjip7QrYYFfOi0dHITBemlmkekYlUVVq+s90DewNjApgig
ScrX0teSZF6vU6+FXn3oI3G0kBcYo0IxPz3grsjdAvfZvWY9DfO/A5aRoDvdFTnX
AI+lKZLrOv1YbyeDVLZ4RSzoVoZiciiTOV5jRfkf6sfIV8eG/dxsGPIMcnxEU/gO
2/4TUBK0vgOTFZqs7p9cwauSSn3W0BZIbtiSI4EY9zoLB+UmzzRppimES4BJiC0y
D9r3H4VwfKAOEVRU4fIyJvKDkodGezMaNMSYdkaTPyX1IUpoJBbSi0LeMnPDz6mi
ygX3ZEvYrZKAO0oJILz1g2oNhixr8yl5Im81dtNSHXUgIWnw4fFSFLOtisjV48ug
mjSeeZ9xI+aUfwVRwVVrewALK3myj3nEljDXvmpmo2cSJXrUgWs7xVDLF6sQ6vTP
8nzrTaOybcqWZOmqxMo5KKAC4V37rLmpbnSfHyMCAkzNG6EBRd3ejYB3S9AfPgfU
fN+15H+XnlETtIFad7wxIgmou8hpNe+lk0Eam9vMnFk3rGDIXgi7b8QHdzuK2tzo
xdDVSUy6GymEvLy/BD34SnGbFyyNNvJUqGKJLdPrIffDoqZtPbeML6BXAFBGGz8Q
GIcW8FTCjNWg3AANjrmLnTWXrp54ivpuvXJJkS+zS0Ev7ppT5/Eqj8G5dski/Ir9
zVRA+U8iqKFqE7W82VpyOdhWB1naJjF3o5IIbbB7fUAxMIYmdaVQK59xxpJ0sf6i
ao0gApBEsaHHdV5gpCPFrS5aiVdGyrIvvPdsVZ5gr3U+E0JlXAZ3OcxTSOl+UKoc
xLqE6Dlia46mGUxOXn8zKN5IXONUhKFb+7T+v3U0JxiJiij2rIuZjrINm0Vlbysd
hEum/lk1dTsvBw16HUA6jYhHLpDaNVTDAvJgeMp8Teasq0nVtoYYrK/tGi7n1mzc
coSjyMyA5i49U30s0dprLm6nUFZpaIxK2ibnEF9OCp+yEJ7o+eM1CesRlrXZqWjQ
/pYyq4C4Q4MxjpT/YcEUB4rJqroX5ki9SlP7ZTNZtRp2HYjUOU4v+6joSE0dNBWh
paN2Kz2HlyDbJfC0qkGEdbpSJlzdggiEyKLCl+2mf6j+gI9WOHoOqPBr80eTLmF5
drSr2Nk4zkk6a9gQ8qIIVaZ3ct/20sbnuxWttLAUV2lD4bFihKMUtmYZuXTbv9Y3
xooD4MUH77sy+ni3O3zyvkA/ykqHwrmvirOsvdHhO8qtmP4zsVTOj7cgC7Ktz3xP
JHr0HKWGt81Jw4BafM6yeQkT/dlaQOiBepPmZl3cxq3ukkn/pfCQjETZQEGKzITQ
VtMbyf5DDgQqswQdoLjC1vrG5zmehruJ4CdOOv6VHyWBElycBAI5dkI36QfZiRGb
6SH/XzkLqnf33RScNr3wXsHZEDeB2048NFkOCcPiWET8enFGez/kgUTj4biUq8sp
MRr+3Mi3wU/lqQYiNj/XvpjIfj+lNqXZ4dxCC5pIzUMkviI5OL3pUS4dlTcb8CgE
liwT1pZH5sU+ZiNlVN50N5aQ4fX5jgVCHpVRDxWzAEsyryI7gsgd4heSwuyrgu8d
W/oD+hpl1p3/LbH+VLvNhuKgcg1BNdQANg0T7+K38QGCXKoFtuPx+D1kjhRC0yKt
zVIFtjSaDo0sRdbGe2qY9JK54FPvaQxaWEbcgZnFpC2MIHrne0nrSudDlqpfE3GE
g1A6fcYlZkwzGKHR0uzX8MUwNtfFvJfNf9s1jfGJTEQjZ5nvT7QTYPFxpCO0bA77
q+rjO/YOqIOWV0hvV/Jb9uyJTbDuGw83y7QfWfY2xMMXDRr3W8TJPEJR92eXoPAR
k6ERIQDPpzHCZ0sE3WdiAC/HMQna/mFr4ffQwvzNhRPDSgFcjFLLEaz5dHzzWWIh
CghOrFhBHh+KNJ4rwjiotVE56sy3zVa7EvgTo02FBUTJdqD3/8FrjXMG439WgyIN
jqxVNKHxoL8bL5a4nkvvCNpPUqaAwzGKKbAp1SmNFO6Zl8sZzkM3rJphlK14zsBc
gJhOZbdBYmPZMJRrjrJNAxkfFSNYTcMjGt3RXScTzJ9h8Kq5EEehgMWVnhS2m7Xr
vRSMVGG5XsQLJvEYtT8ukNp9btNQE+Sawf3CGmaA7OweW/FwCGmAF/XqvQ8xpWgd
jF0mYRuUins5SNIrZe26UsByYodb2CT2nPXGkIIQt4RvybBqkcMtnUg67ZzE6cnW
4+v2xLN+YY9J77TUacxp5w1qjOHqYoi0afZzayqwy01cposvNumZG8VtRUpvtpSo
V0b4iSPc7QTHfkeBcWCWCAEtknMqIB+ZUMQUCaL4/NC1h1uIHj3O++yfb+AunKN6
y5cSojeE+4csgRj88QHIb7nKf0REB32D4coYq6tzz1bZ+YC1840i7O75SJcsjd6m
HZ3Zr2PUuKpcTQDY4Gx/047S71tFfxf9vOicjTleTFIgq5QoUiXOuIJsX6RWofRl
rC5jnBP1+K1TYHzYvCZbkR2oaF71LCVebWu0g0XY7dDfxSGcdceZBJUjo7TreLqj
vmhxIBndR/Z1bR32fZjMoLKl/zphFBnoBxGxX+q3r2YJ+CIf8oUN7lQ241+ToM7I
LehwqgIihDRC8278BAI7x17ousZaMDJFbC/v9CdTAHqP9EkIpXdzPJ+mLU+/Yu02
16CY4mC6KaeAF4/Shgxbo1tcVO61yGt5KcJF5c4wZWSg6aO3Y7c9cXBXaHdnSBcD
vGnqDVS5VWqAFu7kGA6w4S3AogqpuOU0yxCIQ3QJINrcVvtoDiMipeiL5x1uMlPk
T4j4NlRs4+zCLX6KY6NYBM1YYzX8j4S41Xayum501j3NNxLjKmx+/fB964q6Ub0O
KPYgKeOMijEnr+nUQjnC/Oqt6p6K/Fj39K4wc5c73+tSxLeiPqMB/oek9Q42wxfa
vEeO4ID5ZZnIFvJyZqXeJisjXiyB4CuQoJ0MKP4BeKRSndjIFzTERSqPVv6TA+JB
ERI1W+kpKdGTQPOHU2Mgdj1YnSSi0SYVX1xkuukQIWAj+DdA7MAmyg9D9/nhYHAF
7aPHbaMPqDDtfl8BOXebbTZEdezqBlwLUCOuWIPlavSuJ2j66ZU1WtEYj/WCwpqf
BCg5Dog+gyTm+lpZPVUmXme818kBdciyKvxZ9VOYGplwpSipe3Mq3uOQadv40Ytf
/BP4kd9o+nvrj3YKOa2xKx3Xa7lvc3zWCgbPtKn3kScj86BFntkJzSYUj3D3GNHO
LxovXylPJ3vMvTQYiqSFA2uCm7I3eZ7zSeQPwFicrFKu3LZjW3t4Ovyuj9CsCJWN
86rM1zFZvqSt874gBjrPsKz7qLW0Ny+Q1n29jH7C3vHHvfqH+XNpPua3plVJnDrB
xgCYV20gMFLtRepp5DnpeZcecWeeKTqxetjVWdsvCtLIIeiLMCTFmUW8L6WBTv98
ai2+xiq8MxKsOyWVE+ob4Z69b3SZhAJ1TIz7jCKIi3F6ojB7HAyXJtMif7rWZZzK
WPhaDp//kY/8WU7Oz4mknGNekwj/Y8O2MpdswNu4B3aqDgF5BLpNkbPT1gQrNmBR
z+86yb9GC9Ee+JZ5o8stjE2+SsocN/Yn9i8ZnYp+OyShXoQXFOfrTYTxn7zypoSn
z8d3iz8VaWLl0g7HsNvxLhPW/2tHQbhFJ3eMx6955xiVaQWma0yQX4zGXHqwxeCN
vUtKl43Io3z8UjgK+IadrCTABUTLFMZ+pFqw1rXpBMqZAqA7ytH5N6LKaRGFtljz
2xFNMlt4LLSClvPsFhgJQqiihXU5ACrIS7OFbDk5eDqwYgKNzc5udVGqmxr92cS6
bSIYsi1GijXq7qyGc2fe5ePyo2MjNn4bgKnMZQEbpyYQ+Ov7KmxS2MNtV+omE1oJ
vsRtUDWvHT+OpB9dN2vEfz9IDyKJ1EInesdQfO/YhORmarkz7hO2ZC2eLcod5EK7
EpR5o3UEv7R3d7YTRssdGsoMX7pTMjVAL17xAODyIkPK+YUzZVLdxRwJIISsfHUd
+Z4jhcEtEVz1ZSJvIGIMT8HSokncEbG0XKIsbImX+Mq/XtTHpDx6Rubpt0pJu7w1
L0iA6Iywyv/x+Lh/IOEyCEzZMwudhCQpMuhqiamDGaJSibbtPhG0k/6+MwXQtSFd
93LtbEfFi58I8tgeHc+Snui74g3GvP0/yvIes49lViC8TeqnW0J0oOWAFAgly11R
LWXgkn5Qd40yM4ptoORzAxJ1EdEsjuATKeCbh2J4WisbZ+FhH2Ou0ogvr6OgmZH+
qnKZvFvDFr40+Cz5E/ehzPpIHRp83EX6DlT2MRLfri9wM0gnctcrDU2mBZ3z/O3d
OGtd7YTOA+muW50POgzw/EhXjSC/chYQKw0ZFuUsQR37uAYr+Q/o09oFgoK+dY35
xAXwuxKP5PlrID3/VmgR1fQxox/d4YOdoWWEisXm43byRyye2adOYQmNeIhoSTC2
muGj1LX1YsLrtCQG0hR6bM6KVpnCkQgTfUw2EltyIjkDZh1JJWjjZUh3vB/XqbTY
jW81CaZVv7ATxlJ5jdpm8UaQUt+VESTe6lpIeQce41eZZaAeiE86AOZlEBaNNo+w
jUNnpXQZ0q6VR3YiiyOn2WsgSKhlYBDfRmASAkFU54AYETq6CIhSE+15RQBHUrCN
p8FofSoOQgxpMrLErMmW06LyhnVUqClmdlEh5eVN6VgMwkBreozn4+N8ZimuMOGq
tLmTcVqEfelnlI7BvZPU4SXnxn1AGqpLYb2CinAuMLqr6cghCoWYOhlkoxUVHHVR
pBX9ieObvEs5zvMyyoMxXDZSopfEXCkfpKZb+bYS7URiXcFT439XQ2Cc76i9/ssi
7ZfADf7BXibRJtHOUW8ylrrn/15iVe+8MZGQLXxwtFpKhZROKBgVBvuC6r6RvFt8
AEkiDB+KZA7FfgPVfCEGaVLNQhT/9tE8oFgFK4kcnLh2veyy212d7flGdrqQd/fy
vsVp2CYJF41ppACpQK8LLmHMduY5F3YBJcdWe+SNsSX+x4BbTH1PeOSBLWD+LgOE
91UOtrY90aokjj/GSCTxuwrbNtQjR6UI9ZClgP+oSroAogCsUdONzzC2xLNeHB/T
OSyLp/quPSKmIfZF2v2B8lzIFs4Xoc0IpaAHFZuvigaeYoC1bqAXWplda4ZT7WyV
tVhsDg8a/itk3oeChyhi9sPUkQHKdnaDWQ8TqJ5dMlis8p2svqNMD21mIY/lB4mt
N1ePCTriDG0dwYzE40a6pMhmKsYxJzZHej79b7CPJ56clOMzUEiyexAl5Bd6A6bG
bRDQ0ahvqkL6GCafLAKxJlHK4DyQOiHT2dgUHK7aXIYc7myyiPQgTS3AcbygWsIS
TOegux0ujh/529xmv94ss9o4+k37NuYqdfp34KiuaRyW+uhr0hrkwzS6KgTHFf5M
6qxzyX5Js5mxemAIIE/jYGXN8J+0DtBz2b9tMiTJ3JlU+wefz34N0oHEWD235Xw9
j66mFjzYtCP34P6K+aD+DaZzycXKw6gyyjAvB+BorjM1QlEESDqtsyQE9N1ZG0JC
L8mMgCkV/y99iXaSOX7/H0DHuoySuyel/kr2chENrCFQ0SMsEhY6Y6AGV2CDPm83
0PvMLI+ENkEv8TXHhAKvqRezAGoaFQ9Mloa5rFnjxxJ8SJXJaQCxyAdlei12FPTO
KnbBfKI5zmEuUxHnrUZ1fkHQX1cYS0FZuoG4jY8nfiOOjyj3z6Ma8HIehC8NcJqZ
nKDCYwu878gYFL+6o7w5AA0ymM3T/jEErm+xkNAHrieTQCr7ts2kURseA73eX15N
CeP6sI0YP5Q0uADTUzk0ZgsiRC4oZEM9Bcuab+nvrvweWfFNNzKNcYqIlgsYHs80
u5j4lpEZdLo+/5D+U9u9S7UY+80juijGEk4A3X1stTlFTitMIH2qxLKrHs3ShyX6
2T8daTfLISLoX7aECDX3t7UgCm9stH1HMpdco8uIXDP/i+RPOtzZOUF6hO3MCXM5
bWzIpftzsvL7m1EFU1+a9WNFvVrybn+DU74CZhNhlmsNcQJ5Huo1blb4NPbSXeCY
hs4vYe/+1As6uHNgjZW/wRc7IJtZrH5xJSGYGja4OUeKJAM7ivDcO0yh5WRhiuGP
DXWRR5egIXkxF7h2zWpWWYNsF2ABeUaDpYYEpiB/mc4RA1zUTWjG7voyW6Bya7kE
6yVFF6EnpyO6G/DHlT0vEtS7bVOToy2OJLLmsLxhIMNi8a2pmPFls/wxdWwxlib3
NtZzR12/ikT5ZZsr8+JAXl1xJJo8lZIZdSofhfxZ8V/lWVXsfwmKfwWkDkwX7/AF
dzGCexuLJtAqB3J8VxebOHEjiKa1vcjrikgIMCtYQ2skbw58ktEDQzUdiO3IN6oJ
ZzKnZH7r/zEaCVhTM8vZDnjIeyVbYiPPqoGzbc6y21fBXZzqNAsP0smIlYizj4bO
SA+nlRXt+ZtdcdvXfQ+FuKUcdBGIzLAZ67PosOKtFWJS3Rzw6BIFWx12oqMQ8XeJ
S/pS41YlDJ/2GGgB+9Vqiq6mQyFMCpA755PTCdcmHo8Vbuk6d/NFiuow8R+1qkAP
3wmw5ixwaoXXAasve5DS0YLvwWYf7XwIiiX2cdYJmyIFvrlGzZtXg+e2Y+GCYSYq
UnwA2Bv8hhnpioHsao77JITHDNbSZ8mmrV+v8mOUr97JRAuOcNFxmxbcbSWyqjRN
dfxkRPpk28YhaQcbiRph7Xl0W2ykNyX3iRh8sdAROCrL5NKJ/1ruUUy2TMTn4M+d
tgh0GBXQbOIZbReHvmEwaGGibAJihYkBNWjItSEHaacqwUV2QP7V5c7oL7Jhs/iG
EjPxb8u4GLk1JPcYyAuGSwrRAf2K2upK1MYf3uYmeLTvHmCemVq9tg+/qH1Sf3Fc
6aLZJhPC6AmBQbQFMPu4Z4+PeQsSpYxrRt1Gw6etrsuksykvmknHgLQtpxl7nDBn
Twt7zNkwZj5be5DrwGI5CDqOYN/76WMKnOl0YuAW37k8vSGVi4TGn6q4OumTfZ2o
PRAkbQr0Kley/V+OrMc+PoM9Xq70gwaHRuZp0Z4XzXXf1xFcRvU6Vd7n6FqOdEPC
Loz2dEsHII/II8OQSd/cQzVr7jJ4xtcagcn2DFc3BXJ9gzoIrgruuuIqJRx0w7bn
v+52gM8QKDJbhQa2FeVDGLjibNKZDWgGYr0VXxjkPn2eGAzuClq9tENkJL+MFQn2
yKtAHkk7ZM+LzT1rSzpvPnkBOmCizEO+Wi39UA7Wl7bkjucvW+kTHzydp3aD/RTO
VedzdDljySxnmegt3FSmoUIzlcHVJbV1hLs1YZzy78IxYpqZxMvBfCl35nY6VPak
6G3+SqZZvNiyeRB31Nw04OQwv9IbbAd8vhH9AGxDwYcR07XmiG8sT0jsNNFqizH/
pBkmunjVatbAXoLHrqj962rrchZdFw3REnrAbXAp4c8ZUqZe4bQrRrNKzeiJvJas
0dKVtps8elo4oHHfS8htRosxZiLoB1jeOWwroiMD449TeGCX7dwc24W5qMDc73gs
pSzzPP4rAl4B8RCpnWOAoMdv234SWIOCNWM0XtssrTw/lWsRVIV3t+WOLxMrZetR
MnGHRy/WAZV66B2Vol4ikH2OPIspC5Q4ziqbHTaO0smNIeTuZzmqbjlYOBLvYAZH
xy/Z1Mt6WjbrM5XVMD64ZSxvx4hZZXZ1Sbr+aS6FnDCwJXy5d8rCEe7CZVI4ZmSr
4Y4p2R5QplkHefURo0RTsv1GAiB3/cu168pjpFtFbRgkIXDs5K4Hnbbc12RQH6yF
T2BdcIBEu8jkIxj5fyqgZRJJRBbzv+H3oo/0TQR80CfKcVntjSpbmvvCzBNufef2
Y20iU5pnaKADUY/U/bITuyXcoj3iV3Fjh7H4OSx//X9GvZR5oKcwIjX9dkwdzoSO
RhGlNnrq7vKxHx0YTGxfWmS9eBSWND4xjiNjSYE8euEA8/RHJuj2PYlnmCVitqiL
Ef2GjS27+UhmyOBx4hAYHcdfFdvzrXjiEdPLBTbGP4SZknC3odRpMjQztgZRHf7I
PXFN+MQeyG3FlH29gge4Qfk4F5J2g1A/xLquR43Y268G9jjDMGjuOEGbaB+k1xgl
k79goUlIBMWi7NZK3fgbVRIq+RY4O1QcdU2zYBVTJLiBzSDLsjk9h6F9oeQq9NUf
L+7D8DMcBlhoTEnHNMnD66sOc21kzKxSet0ANHLiTz7y2KKOrpV88TW3cPT8QcPJ
VPk25nc1n3WpfLbWdWIynvUhFJLYo7U5isfY/+hD5ulYP56YigtmH2zlxWHoQrAN
NZ4Z1L6izpBtqgvI1FYSM9Wd5tkPAgg0Yog1X28rolB0FkH/FKM+K365veLPJVKf
yW2BRQp3zV0N7BTGFNhvCqfLqLs7OEAfNccoFcVrtaXB6tvCvHbA+Mxw+S9C5Xbn
Zfa9BIlnn+U2adu0GhX5V0WRYJee6ls8oYYnyCit5PBaNvvQu9uQXefHmdKGIetP
FDng8my8KYJgSRiJQ54zu0fH959Ti+/DlRrhZSjfQcBeb6yX/bgZ9g050ktsGeav
DQHhM5ahILtFPAo5SKlJkTgSSlN3i4tEDUNHCGa0iCUVDqubs3fwus8bzoQe1z4B
DJCLwAoW3UAm9GVWaMWVZnWJDjsmmJHCvK9rmie9m1izvkr/x5o3XvmXchl5Mh6j
nXT9zEGxzAsfZXnYTlyeIm5afegMIVpKkA4tTODQJ/HwVoczrqwA7W/+2w+IvhdV
UkBjf2Eshg8V3h6dmNumaMY9bAhXSksni0L1/wuh+CMTE2+6VUokbqdlo5usPkqq
MZIEKVFuh0Vi/daTC5JNyEXeXPtArmmpV8t1MD4zOR6FtU41LlgTo2QUEtXw6G5r
5Xm/ilnjabGVqWIq33Dxtcnqs1Bh8aQ3AX9IGpY8cVN6uY+zqhtG88sNXNU3sXte
G7Tw0ghNqlNuejym00fzm9OAbkXLHpoZWpMM3gTWByg5N6nKS5razS/bT1Fgo1l7
8Zae4FckqbQ9jmW+lLEc6/YywQpsOhzX3GZT1B1eL75XaQRY5h2G+YnS3SASRAON
It9ZGi6dMuQdKav6/1HXSp9gRzsEGmdfrjNMSbtJFreg0J9CGxDIM3qCqArEr7o0
BtuKRbQE7JQzXaDBj5xDVH+7Qd0WFVbZeGoFiubElxYWm5sfruODXJVZ513OxMJH
2xrhsoHVpOvuoJkEhWL+zF3vA+Wg0KCy3Gt+OxCRFlopjUCggBZRCq3TMdeoHjCX
OsDUKkSINRgne1HUtZyc9WG7sB6FFm2AMJHgQTVU7hfIBHkcf1E436PZQ7GP0zC+
w/SGVHhpOr/Mwouy4QUEMtYRsYw2CCVZlpdRsD+OhenY1R64+KckLvE+sz/w8FOr
a8IVBwOqaVnoz4vnKsw3j9mmFN11Ld+Ce0Rw/lVJXVxI/N7Hgflvz+G305m2QA/B
k7NWOnF1U9cQAFsn/aIcJbQ6U3VT5+6iwS7ZlwShDzY1EL3Z0LPhNCLFeCN12xg7
5/cv8KDAlc+sXCDcRneoimeUcr/xVmMD1gVck5fphJcTZkCbpgE0EE8qUd8eVfiP
NqryLjrZshZoJ1mEDRCN4GnqUW5263CpwNEmSVrUBwyrVXCgMxryMSsx2hNAJnWa
Ch8GAw6I87eE/k/y57ODOIWTYa98iqTUoFhitMrk2n/904WD63sXva3mIbHPpOZO
IZ4MI5HODt10Qutyw9H1FHv7moAcLFDi37TnmH+surK9LWctbJNhg2r5t91uoi0q
cYl8DypsXdaUNwt0JayPVIVCmak+4zeeZnz+CWqOaSNEdSyu0q3csn3B2Div96yN
SRW+nFWjlff+dF5JJNTv2JlnVnYzwPBHd/RBGjOVwkkeJiOsG1EdN2TomHYn/MuG
33XNMlQrG+XyOHTK/jFI5rHEz2DYhTNcTBDovZjAnMgf+aI49GSOBWdLSzPaQYjf
x3FuHOfy4I8ZmRbF6D05GIQ5YH+z4s/JBFnr7Wgfarly50vki/QKvpq3RKhhv+vR
jWcDhBu00RvHsiRx45I00AszdtXHyQFC2/zxMouEH5rLs+k/DR6r7fkIZseeaIKv
5u/uHq3ESz8i5DitBb2Dj70D+wgwaj/X3XqScq6Z9lENHf4JldiYiN+qFiYqKOpm
5sQ4QVwC1KvswjFcb/BMRf5heHe2feVsWQi9ZH5JzCKxsrIaRGj/c8eSIWbZveHq
fxkQC1F8RlD5M36ZqGQNoax4Yn4x0yZlDjZsI8RaR+XbzukOl3WMVEn8V4wo4StC
/VGctkod3y44Dam2h0UBIZT2Tr6CPysH9tth2yIedFkICsVkM5zwWT1SQPVWsDr2
iOySi6UbDUl4Iont7VvThvczAaMsEAF1GyQY8cdTpkyI2y1IjVuShfap3MWoOlvL
UxpPYGP7xmjKppJhQM23Z0bep6Be3VDa6oZKSfB+6fKbTWmK0Im1q7VQp3yC1W5D
rqo/UU7qa5zK7r4HX11tKJXDhdyFedpsv6V/o7f61kI+7wf4Ntgy30WJmEu6Jdka
NpUmvNxzvwUqu3Z5dCruhmZ7BuxFl3dL3UaqSKIcXZCzEcOtGFQ2LKKZ0rqyURjC
xsQOCxKZHKnLjXyBilJpWTujvN+QDOju3aQP+3Hd42ksAymSyVEX3yTOfWxtFAfx
UBARgPvOaJBX2jXkdP66fnFFPZuvcFr7AYvyIM2HWN+NhydbwWSBwarUwLbxlw7q
2gqDl+OtO82ECeZ8PKOh+S+Kgo4wJnpEyJ4K5EdK00sRaj+JsYcyiYUR8wygGzfR
+vmywP58tfZHDRZHP37QfM+VJ7TKYT1Uk6UODJNArzVJXJf2JhH+1FNWbJz/YIuq
FPvWmDMEYS0c4snVFHUL/HXflhQZvRcX8uaNQCULWuulCRaRLoXTzqNWRx85y41v
ULAezwr5GvuO0TMzNc/G28O6axC5o30OZllj4gxxs+gkPBgDeXx+5EC9lA07j/W3
T+hUqBCM7nv3oFWTQLMjz0FcJMNP+T1vWdkoiWV7CilpVeoZWknVwSTTAdmV+YGP
/z0UZWm75kevAvdwoDJ1rSvFkud1ZwQNjXf6/AJuckwINaRe3EMIxtojipZa/8+J
ywVsYMvH4LnUP/avM3Gps6BR7mGLcQivyzsde6dS6XeRyc+B0Hf2w4QeeuCKpxXF
7mBW33uT1cSb3Nma8vsUs43cBFjBsGWn2esLqM9NPu+8+8HxtAL3krrqoqxUTlgo
s0EC80f5cQkrTp+qp273QghDY7AXi5zKKGDfVHQCY7J0b9crFtnQ/oIn66LTymLr
XIvYeDNWW5meM7lKPU9cjR2A0IX1E9eIj4DCDEWeyB85dCztrnaCequH8Kak6hx2
DX9I2XDKAnrzw89VYQmPFVzxXq8946TS26o8OxAu4Scacke9TjPRkZFB9WabXZDU
tXQA/1KcfUihiAQuYgJCktA/4Fnc9aXnSvVkqOak54uKIxTL2VfnNDcp9iHHZ1ee
TtKF1J0JKKFrm66Mv10xi0p0t33CPZzNTYLNf64NU59KjiKRCUqh5FFZIOlYhbeR
7XFnloX1/8JAgdD+Tg949WNguEH8EOxglbXhABXmBcYJMfYRyEwap+I6A0L7gK6x
+xlQhZXVvDOzxk5mZa7EkV3pSGy4OwF6zSz+FTueRI2vMQvA78hBRGh6p+ciHM01
f1raWmvHwGj/qqpN4M36dnQ6AymokN1QsI/hc+nINOK5mK4ChBW8ATB3bCVoBgnO
Od6O4PVlPRsNsg1l0Lhi6sBxfEf8rjWTJHxrc6APPmNRaOSWxKMv0jfI22znPDxT
1mAl161dOahQvhAzoXp4tKhTYkyTekIkLqPqIY2E7D6gpn/+jbVb1upnKZFvJb6t
VZXaphJyQKpY4C4e9sC73HDE6xupJlXsi+IpG/SNcgedR1TrM1D+k/sjtSWL7f/g
JiEPmkieOlWI7LwvFRFgrm2b4hCUNM9eml2sCC28c38gToBx+VTZvz3MIS/IRQaK
Vy7y/6zckp+2pibQcgm67lUv+010CWfUHxSNzqZLQVIY6oSMSjRnx0Zn29SOYsJ2
8DhreG9G1kjd4eV9KyhRz2JLf0lYStpqg8k0fd/IvjRdix8QG8sYEoxc+OGrBHT3
AmpgGW0M4kE/Q92FM1ItTZSFQQt5EnllfQ3Lcdy7G2YR24C37Arit8556fPGvJbE
0F0GQz6sPI59mNHRpYR+iq58DunIn6Lg3aEEhnc2X9BSuAX+1rCtqqflH62Ns/u/
lMlEihTeFwvshGKdrgubiCu344u1ihqjuMLesxTD3hijW/L+ZicsgPDCuV0qQdMe
o4iuY5MPB35ksgIR/CkHkmxwC/DSJBe0Z31BUedFRKct0zsTZjb96aX0KoXxqe5Y
zYR1VOUWc4C+nWTAWIETvJumAOuppKgcsv3j92EdZy1NGgTCEh0MqHYde18jjtGj
FATw8A0ea1BaH/84HPpfJswpVzSWnwrnUq45DDaWjP7OKH0N/IbIK4U7NGpiy1Qo
NBVriYkdFuKPFe8xnWfBdT0hyBxNOFP74bV+EqEmcAseXRi/DcL6m18FoBX2MFlT
wFsiE3HgbcATTBD4tW13eWK+9MI9UEtN6MhTv0aeMUk90rfYT+PVePhVGZeaMgcZ
dNFvV1Jj0KY5Ey3DhF2PURNfAmElKZ+fTDKJ+xcuSZad9Ai1bWCxW1nKK0JByT+Q
ij32S0uQkcNjf9eMjg3a/tk1q/T5ZDZmnL+opSuP6wgkArc4IeNjpq6VP7DyfnA3
U17AEa3uquvma0gCs2EsCebaeeLxRNTgBMIBDz2E6tKqNAlU1bLwb3EpPNIjaUMs
5mo9cIbuG2fNHGH724HSyCKpi7HKTXKPuqywPzEGrBRJf8wWbG5cisDN3Wv8S9Df
GmoNocztoVo8hVmhsVfEBOBvWx/q6yzEsdCzoi8lC3ee5ggGd1siR3TV+3om8rNe
S66I/m0D6+i+/Wl2bRCWgrCQ0ki6Kgx2BQmDL9vx/1klmSn83/noWN0395JUTpYt
zKVRyKAVzLd18iZByT+jYOoMNQV7Y6M3oUVmS2XVXeJamobYIev9S8bd25Gjc9oh
ppEyN5vb61fa3gEEd4hZ7W7IOOuqkguYmMY6yMcVuwjHZu719lz1PkWt23I0ynsZ
QDfqbgCmZNfiz7eshQ3N/XU2vImJzcFCx7Gp4qsZCUqnj2VVXqbhFawmtSEKy5yZ
ZgxZmv5abMjW6pGZnJYOHdX2ykLtbl2Nkq7Ui3MqUPJPsOdxAF/NNzpO3Nt2REAb
umFo4NpAAno0H967qF9c1axjs8hyeVyevojmbc5eXMWzWCuFPyPWmdtpn52ArLFU
ZaHvjPNxC2rPxW2WhpWLtEmu+REl1qSpoeToVPSwJzIc9L5u8xdSdySVMLfHLUXE
yii1NFJyCsiKZc5Tqlc8AftIISTqzbbHWcVXVBftMjuCWLlN0RXTfKq95UMBXsp9
Y3YRfE01B3SWAp3VEEveAy6RPXpHWxiwcMiAPqaMVt9IvFZXaCI2KuX1L82t4Jq3
5kNME0p6j5Xazv09DmVYIzAyxc3XNoqmWsLevRtTe28UP9YZKytGP2T2PrfbaF+U
cGLmd14DjC9JkYaUZZ33D6w9brivMOMavzJICC4HNcyC98+6D4J5HCR/KQDiOg2V
7/+kg0DD0ydF1JsjU13feiklKp/GaOBFOvC1HFCxnqhNX1S0NhxgYPSdduME4nBr
qw23df/fSZcHiO17YlTenbsrCa952bywHurT2QB/YEiXHLnseiwGTedWfBVSEo2J
JdlT3euWVERjQjewQpxmGqPYpZya4+X9ed7hBT86IFqMMfOnIPo9/Q3podjomBrU
EyfpFi2s54cXgRiiDfjKswz9oCmh5NhH0wwI9zk3oUzzSl3V+pPd4WnFgo9o1Vlu
voRS5MN7jkyT17D5tOKK+za3Z4Y7tP763eXeREC6WWVtabmlwRA0yA/X7kRXZ7ws
WQwCYhMzBnhgOCtm+yF1IxZjiNeN3SpzUMvJDImbKWKKhI0YrCGqwHqVEZI9QY8m
meUHGNOQf6dAhWqV/zPTNe/RZjaHcZWIELEc6GLG6jh2hAQipBifFxk5OFQQrzAW
OqirJ8BuuEM9daCVvDEj51nP3xZNbI+U3Dv3hwqc+P75bnsvUBjCzKnFYS+UAPlk
2k/C16S91iiBokVXn6FtTnK0Wl+6ZwK8LlSJmWynXdbmCvN8xN6ualxcPVww+J2r
B3/a1po0zdDXMLPlvJ7IrLL6TyrKuUiZZyLQZ0i/J12NH17js7ZqM+y5Sz4bRMIx
t7T+E770XJmn3j617HZUC6e4gYmoh/SkjWYfXWaSj48wgVib6rQ4r28qjYR17SEq
yYtW6tTkSSz6D/GP1U4xMjntSU8/xYY6ONHhg8sPaey90pKrfGrPz5xpflo6q43U
3xbdRfYQpkStC6rb8u2YMq5t9dcrT59Ep+jp81pLE45yy3pDiFrHP70BeIRKsvp/
GhVCP/Z8FQiY35juDRY+w+xjLi8KnNFi7utgSgHnHmaEq46HUmw0ypEX6XydnsUb
ttKUEQ1PB6tMOaf1Wj1YZ/xXa9biU72SyqblVHQzVv5VF7RBK7SMggAGbCiD+GRl
WRm5QXsSw7Y7Y1atcbR/bZ7iNe2UMIQuDfDGPt6w/3UNuWUYkLGzhwgCdwL2gqq8
YKrb2IG28GJbTP+liNmt7LMWPDtRPMAAc9ZHVO414Zm+hcRJgbFaxexGYx0Mr843
ocb2oNyMDzIFu8UtPQUAlZ05TAIuJamKLxFTqbS8rO77KMlu38+Gx/AEDl7cSHc7
ugvCxzDyciP2Ib+elto847lNLzu996Wwdb6dZsMo6zfOkeGZClDjlR4SIl2NTBRd
bTshfjCQwcLz0Ml4T89+Ssih34iaRAM7I57giWUkWG/L1BNIBClvDw1JSwl8Mtsj
dMvmg3ddRhJLbxK95rDmIWaN7RHnXMaWrv0Er7cdR46Ie25jOOwGTBNT7XCeDGPC
Fzm5SrbjIsgpg7VTLKFFqqIA9e1leBpoa0zt/Yv5lXGupHkNIHmOUdagkOT60sKF
WT9cC7xKmaC+t7AqQ8MEtZS2aP39aPb/2dD/br30A1ocFOs0s57ZrwAvGUtoft+i
U8lnJ6Uoc65W+8zUtkRyf53wrTufq59pA1DJvtPnFijjCDtgJW+b7rNGw8H6DRde
9HFoVb8IPpFm2+VOhukv+9tv047ZH8DwPgi/gFhzcrEWkfAi2OoiHlZS+lJ7gdRy
fVzfJYlPhp/67CMSy+AMwmEgDsOW+Sni2dTDuBBPmb3y8BqvESFRIUxoUHAWBh20
b3GE5h48CSBgRCql09znIWMcDOJ/7CHd3n/7wfoVlaa/s1YDQQ791GWcCsDz4Lns
W84WBFt6Qste+XLJXRxLSPj9SfOPlx2Ii5wfqYqLdn40XlbEen8705saw8TgIEnU
E7yZaYwUIbnSwFBEKtcHdVKDZpYFSmcJCFDVDJCSIEJVFkNDfedzHLDG3DcIQDWH
9fGLQ7WKSL0Jmd1L1NqmJDDqnlIBWVj3W030QUTFTQYxH3wviDKDck1MtosWJnKa
iR67UTAeqIJIjcb4n2bw8SdW5h/LfYTk6p3PXn5vo8v8qjhbdzpc2yz2qDsnXLl6
8S8UBBW1SK2SFCOYBTOwllo5v8FQfRoonOp/YFO9GLuAMVMq4Ulz3EmGbqgPopSb
YSDmfwc+Z9+znrYyPh2FuhNsLTna3x72CU2rU5e7mK1IFvxORQeNiG1AgRH9UtSY
DaalxljmXqON90S/gVS0fuf2MzwxW2ef/NNgwsYaE3blQT8i+x3ed42U8LMihnzs
qXDOoZPzAkplUmAVQSEZSO9yN142+K+bO5I1GSG5WxRJ+f6Mcw3/rJgKHZMnktle
EgSlgSkjbxsv4a1rtBuUgD98ieqfJcWRV97yDgOT2C1Ccc3sBZ+6bFJcv8mcB+Jj
OH7AvMCFjYBkOUkXitLQTVpsysjOmZpnpg6po77VQMVkCgAQywdCAOruqOiM2oW0
GR3FQCtKSmviW/ofUKrzdHdJUdws/IOfvoO4nHjrZ6lVDqW7IBee33qxVZ6HosYc
QP1ffCCpnMqoxXC5azbK7rzTypLWXr0bRZv8g2EnKf3ituY3nsBrV328fJtmrINu
tEJ7Yh9S28nZGpfY5E+A9uHPiNG6Tk+EstfX5bleXns5T2sPu1LH92xVjNnVlS0N
vuCqxr6KtELlMOTYrHTv+FWW5WR2EgUNVuD1IyBc9wE/onzHgZ9PB+SvbVl52LmF
Y5ynh04KOjUr755BEx6xly34g+Jr5lT5ipN5ZRueiXRy2vYS3NngZm7ao1HG7Nar
4GN6n7vJD0QDw7z5TkjynpjYO8ULe0XM6adqq7UaU523o8MaosNuHyF36oPP5QOs
ewnoUV8Zqv0fSkCXVfbq9FY82wPa8yOwM9PlBPj8vcMNq84o1QcOhcdkUgK0xfph
GLahLb0AakwSFUMqqcayTjhu6+quv8sRGiozrDRbDt50DIxKzqRfmP19sOlufso3
wupad3UolEZl1y02q0daTm8aYT+9un5lMcATv506Hp8MLhcf7ogW55iFb5r+/zpJ
jfr+B4qvePgLTjqax/ou8RpX1alRrFGbFs9trvj8u49ybVJ1PyCJEvSJb62yT6mj
ojZ8apiyU/h1Oj5lPFhl8eaAe8x6munUaXOGYLZAQlYQfczfkzDo7/4nVy3rB7Gh
HTv0R4ybdK2jP1jRfbu+8Lzf3JXo9HXlEc294nLNVySY9rsh3IWC+fKV4HbC1Xeo
w4WgK2FTtdGtDbYRwtLKdJgJQkvcdwvblRaneRtcCDYXDKht+TkQAV/5PAXlEyRK
t4HwXxMRGjEAvJmWNe3gcCRXeJRR+BgSYzVOlNrV+dlgu8c/tJf6jWQX/t/o5fLt
Gq7SLqU8sAfSS5okQ/pHMRSu9wkZA9s7UI9bbUTijcy437fM0jsNcui/VjxnNGCN
YutVWXxHc4GrSKPiQAQSr9KnySaf/dY8Ti4rnmBSHePZYq/BIvQXoSkLjqQOERpI
PbgQ6Ov85UVdc3GIASHRtqYJ7+CUM0lQNtExQ9yKLK5V3MG9I2jmXuRcXgAoV7e+
ZEv9AG8TWkZh4svRfLrBl29tc2l6KGabeU22m5Z9OfD7M98jfOWoG1etYmEIBJQj
xCgsFpQIsIMUhcdBAHoPIUrPX1gsBrvJHOXPi3v8XpoCqyZhiB5RnmDrFiFiWqkA
PUd0ADHpkcMali9QAvyw4+p5UXgp8OcgEmXY5HCcxmBjbltk5R1imgHDDQeFgxsb
mOvfjHEQXYvJP2dszmJP0SpjP+VJxdJrcJnu6MXXbOoNuq++XgOgc5nVgsxGGSyC
G4cmyO/LN33EdCt9uVAaWwXlDzCwbOLxR2gPbPJhymrv2vHoKsZU4U4eCod2vDG2
k86BU6NNS9PtXlPnjSTlsJevyLkUrukotqtlHOqPFigb8qn0l0zaxNiW2wEygIdt
6uAtj3dyDktcbpmED32hi5sxGF8YW21ZqFgbbJeqFMAJdCKpPSl/rKd2uTQIBxJ3
l/pqsQ2YQAMPas2IwvKI68H0qcXB0mMJRnxrFxKT4Ey3Mzr9kA0JypEl8zPw8hfv
q7xcivZPNOAPqf+HjVI3R8x5OiMpDkMShDWF/+wFsHosM3Ai2tMcJZtbyA0WA3ZT
9y9Ce9zoyn84ygEC2EhVLHhcj//xeuQ6awWagxcZTGqbQjM9JFwSnSvTuBR4AMSO
YtVTBA++ORz3wCVbVr7rWDPdxigsWu51ZMF7AQv75MJJEHvFkqhCtFUzV42kzrkr
zvjoBZIWPJkPB+LZWwIYXHi8I2IX8pDN9ZVaI4sCPoMCawrrSLKQt6KJoWovGNYM
vuxqC8Guad6cHH9KayYEZYv1YnzkstlAi9Ti8zpqruWEt9U1/FvNFcnsmd7MfP/h
wxDkqnfs5t+MSru73pUoIvG8NZ834K/fBPm6XeBT7SBVDNLUslX1RXvMexcwd7E6
a1Ik0rKTzXAghy8xH0yXWWbXPgiPAd9TB7DXhCmJf0m4PT3nz3MdEJCFcWLVuWds
X5dcMJ58o3WuSCLBreYPX2dQbwaaQPWncnENLHkFNyuqEs5cqd9mGj93rjV4pcWK
Od2LGS05kP4OUSn/+ewFflC/eGLvw4KrMlCbM4tWnyvx3KQGkAy0hzcQZm1RhE/0
EmTLZLtK5vs+NrJxJU2TBqcRs8SD2Lp3hJJFRGKwMsEESr1hRQb0Dg3xsut83NZs
6CGwt/bF8iPNckLgXn5kahWfarL2BIaVL81suU8roDHzG/TwwArF9rtNRxJIgdZ+
V2XH57KxBvVjw9UpZlQ/LZAVajYo2yVGaQm9D+4Ev3lMY07DrhvH5UueajtaoxwR
esyO4uelXZOZkn7fD36TD2fpNN0KM8Cx4KvvciNcmOSMoY/49nRcxz7jJCaiW93R
AT0Cl0d6ndDwarP76MI2OriIzsc5DYenrvvg+BaeLg1D5vqbr/aJ2Fyh6L/F2H1d
LhzcgvnjgPIFCHVz0WFCXza/cCyDe7/T8hX9KZO/apZrsDIB9zVTKWFxh6M9aWDT
+LPSjAyF/Mqg+tFHb5hn0sJ59NY+0E/O6ELyoK1n5NEQnGPXB9IpFTZ7HCxsWggX
kgG/VcWxNtBvknk3PWBd08ooPoi2FFCKsOK6Oell8/PaOeaZjCNOtkc1feDnE/fD
RzCQpHk5NoUU2qyZbl4WZKGhF/hhMZr4tgty+YIQbN8wCUN8qnOYcReV9x/zqJV/
uTLxRaJy/+kuXRWcbs1FUYiu+80Ja3jYxKNJzzpsr8iFrt1FrfbM4zjr31ZecCqp
XqbxM6P7SpmQADTv8qs1tENZqQARlmp8drLfonmK5UtfUesC6agfEt5uLtzvnmNI
2wZ/czPQMc71B670P3xzFJHaT7rwMIfGyghPgWueuAyyUmU14OnmCMP2jqUeVBu6
QOOlvWMaxso/1d+zMdenuhCVeh1pziZ34Sc70MY9AVsatZ88VHOytwEiSWfTAqoV
sL4Lqx+2AB5o4OEvcx4VFfo44sHxIIclnpvEwaMHzX6nP9NIEvZvFigw0ENDycYz
C59m6y/quSqftOAkmMBNUoO7DfdEj8itm91TLxWvFAEM3WaxETZZR0nxVUroWhdG
pR1uGPQuVkgIeVtVRn+lFUEvuusjftnKtokAZdW1p3Pz+S481djhJgcDA7YtTi20
6izFENIS+7CrsTz182pNkDVXTq0GzgB6Q+TJnV1/HvolZxdJ7VcPGFJaR7ejOe3m
/yOt06sUXNAI6q7ecMPPmEEsNC+nngc/w42yc88DVK+9o6kmOpVN5z4ElfYpHBFJ
XYe+FI4FttozHx9p4Q+1o18vr2Olj9dbbMwJBx+RrUz4JY+GOvcyphiQtyfcL834
RmPQrFgOXi9LFC0FlPo1JGPSUkqVzi8ybEErwOCNi35o5mCjsgP7+PNoxTyt1SzF
jw9D8Gxt5LVIfY6gzW3i1Tu/37LFz8LTVyIdxC/VBKs0aSBvExPoNMIQKJLb2llC
KtBmWwCB4Eoi6lmw8nAH2RWh5BG1W6Ex4WoOJ2/m7LlZIjA/AWJaDB74p1m0Rap+
A1tZLl3u57zfBFXMC0bDIaxUX4InJFLGnKsZsGYcAudtj5RtvxUxtuy2Fe4GVern
s6q0ij8VfK6/6OMNv658GP9CazEho1tquIWCzOPNGnqIKt8gStXfZjPP0xA4B1Ly
DVilSXDeE5G0vinKpelCPIr/kr1dL6BxOo3ojjvXvSIt9TSMjdRkPzJMWpU1ctnO
16zWL9cK+RAQ3Wer7RX7O2f8uoVtlTIKR4asKj3Nlo/l130P+tLoN8joGji1IgnO
/6tKfacGK4vUv7toxmp43b43XZw1eWOnlkugRaABAFQqfFNlMM8aG6nPgZqkMM8z
MJ56XJj+0zL6CNNvPGxNZ5ut7rfptOuA/SA4Z5N/kB+hsuQWVKP4sh+BOmOqlSK1
qMvOduHIdPJqBJfR19Z6dmNtuiOlh0z+QtkJjXldi9sSbdGcNUrB2SbNmp3tHWdX
xCGdpuKqzikR1a9IVZOcUWAQH0JhgJuo2WEIJrQ2wTM/ztCQ0GjccNCUgSYUEg0e
EnFhri3YOmxM3kMe0XZbU3U3v+iO01kibzktJ/GhhC1BFGAVP9atAbcevBCO2B+f
SvgpwqJHKtnXWuUalB4G/5lG/RbHxlQatC/1uK8kdsqkrgIy3MSqrebK6RKOwv6V
1iiWL4XzoxapMfHXV9yAYWaeFsLCXkwVS21PT5Y4PX0xU36kLiqulUqIbvvqYBaw
QHNq6i+iHy2o0H4FouKp7t+9K2ghnjEWajUzQWgm19LfZyScPv2Ogb9aXXDFyZpC
d+v0WzirCjhLuhp2rB5GmZgz+X6MlV0JDYgKXBKJdywlRGmbdTCIeS186Tzu2E+a
l98h8gnW8QLw6xuyQpJMbnHuagm2+d9NwECMqwXNq01staO1F1d1efemJH0MLvHM
7ZgK2knUWzDrvYIQAxzSFQLy71+jL/7hyWRi0eB5Xx8jk/GKY5yXZuvoHabOtLVj
KPjZocpMYdMQ9b2PCLqrWaChuH4aqdRq2awYGmMuxMojMfCOahPrYyM0yhr7ac3Z
xtPt0wsJaYKncrpoRav0TZ+kITK4JgDSBX4i/ull3Lv6bkPqnSubwjxBlJ0giH0r
9Wm8l/kWV6tu2txfrj3uxjjWxE5slBcF1/0LXTXO19YsIoGGrXrwT69xMQOHurTD
Xon5HAvr7Nt8N59ecbhwHb+DNv9ug6ZZIRHjOVLVbZ0VNfgQRbmbri1B8Qr1uOSL
0kmXO1ZXfrDsOL53aGaHPr0+gvIqKwEVszVmtKX32qtIw8SVl0ACKa9QcsDxtUCx
gE5qU8xaCaYyZ//YPpPjQ++X/aQPdI6hidkQ4TmPXetDzPNNn7zZDf1a0P6f659B
TPQtTQ+G3QQBe/FlCSdY1rGC4kO3lxrmQGWRUkjnCTSJB0NJcn1eokLWwUue6MkO
75e7rVj4zjcjmWBTOG4pubDa2U+rSTebFB0J6lmfZyaRBNf8sfrUm+UKNtLfOeHJ
Vc39U5Xr8qZpX9OR1lkhpUkHIT4EHLoxZbiJNDrwBMrBcD5O0J3FmpW9l4FLAel8
nlC8MqLT0oVCK26F+h5olTfe7eOcLQyUUvgNIxDPijgUdwyTDOer2W1OB8DjPTVl
CRIiveWYs7VyhF1acf+GBuJQaGR5SkFVap/KHG/CHeIpjRul/NknS7KHRImVWbMe
DMhnyr0j8oCmkEgddYoZPIVdiouyiyfd+uQF6Jjdm1Jzq4EmHWe98EKhvlzGccam
qTBrLBZTCdrFxsyOpApqUpseQHh4f2wpkVd08+6ub6P5sZd2IsauiAIg70qcGPN8
TvcWoKayNkulkwoXR+eWhRo+KaNXeHA/cQilW89kwNUpAbSbV8ae9z/WPaByihqN
iRHZxbjA8+o0O1PhIQqXEg1aLHyr1RkFYxXAw3rVbEUo/feSHybmeu3Q082RuVAL
cUIL68Rmvb3LVw1upGoa6iPjpcJfAfluiPdCiYWj3BJ0d7SHyGOH5Aa5phSK8npQ
HNzvACjQYhXV/RHVC3PLDaCGZHW9p5SfdF9pUn3K2aZJfSMJxFWIRQbfQMzfLsNU
99lARZCamXouTuMi9nNP538U9wfb46GU8yJn8DVO4C4ZlCNcG5CfCMJycR4irlY/
Jsqvkx3gdmvI7hcOqAM43gEostOb85i3g4zzFke2wHLj86CD5M7+X4XHgK5dfn18
aTwJk/uaRIWjJkmaSP3nDedFk99XDQAOI9zEcBOUumekOeHgnBbLNPSIFLHt69PZ
Ur+yh/2uN/vHDu6ECtri0SHPoyOLUUrUJRWNy71UQ4PUuh+qZOnf5GdcepRbUef5
7E5U6LyLXgzP7XY6uUanCwZrQ9HC8Fnj8DbkLhG3SS3PILZme9QWodOCI4jbKCTX
wiCjncLbKIG9cud3+Pw8klEBFehwm7u2mOQUFdf6IdwfFDNNNJdiSfzhK4obO9SJ
D24EyWgL7fHnuIF1C3I0XjwDdeq3FaCNoiliS4ftqjaz1QNyRpYnGyKWSyrvGaWK
4Vj0FVF5yTVPkGzQ59fO5Gf6VejQYsznz/aLLl/OdmZaag3dsZ1IGH/bRTEVpPXY
WKMPqq5dX4aY7upvz1hqYj6L6TSrXxCq9RJRhSDveYqtpHj5ulGYrG3tgIHtZLMl
1N4ZeLn05h2V/9xVXtMCwHrz5FXeTU2qjJsB6xtnmLH/lZ4cG1BReiT0SUxDOm3F
DEPdMeoJYGW/MiQGwloOLuS4JHPbihMvkgemj0pjJozfdS9WrXpiD8PbVYkJj7qr
pfOznKkyZh6YnyB42N3AUu4MZRUws92dccD2Hv2xByh9GyZaaTvlPFfMr3JOH9tz
BU8maJy1WD12eR3ZROurEqUs8vyE+HDy8MhZbhm+Nypl64nTH/SGiTBxGZISwe91
8IyuYeCGqHyPNhl+sJ9SXVGIGQbZEPelkdY6rJUIirWpNWAHlyEXYS/yTozfLDdM
qoUQdBfTfDWG++Znh/dmD/vhU/543US/K4uBuQd9CUn1ePnu3p1UTO7MpJJ0OFt6
fjdNXiyuUP/wMnGZBhD+uIgpC/K/Pu1gqurmM5HkBwn+KwXRVY2CGxV+SQyzrXD9
AmboVDjX249jK5xxGNP2Sh3CXkqff9kmdHYgUCXa9xPycQZdJqKgZqFbJdky+haQ
JdwnK8t9p5XzwiUbmXU7iHyBcDy4p3j5JjfiDHJ2G01iQ15l0x3JPA5c5PxR49hz
emdWsDd8KXCY97Ff836HwkGV2twCrIW7rJUvPlztGbhQZ+sZtZxdTGdcOxYvfxJ4
c/+MgvutcsnIYuv0iIgkHRU1UOXwWSyidx5axQaVYGbTNlI5RYYgj7h0PSIp1gL5
95YPGzPsUNsXVTxAWmZ/you/ttxNCOxj3QYn/xWdZTXG/Yv+MVObgHJJyDFY9Q4p
NjZmmj67jZgxE+kH2wI3e2xzqrgvk5D6P2PAWsXucSIslWkPjarYgKWXiM+pMFGj
RlMSTfE3RRDVGStz6CSouyirKsDql1EPuRQp7u/O0Rfoe3nR52WrP/v/82deWzcx
FECUUfmu+AnkQUH2ild5JYnRbp4iuQ6XqogLeWA89c9TARBqE0ZmLe+qdfc47kr1
E33JXd28oBG4/jdraJ4H2Qzm8aFztELnfCV9EGfikWiOwrVk4BC+23oWVGS7Q/OJ
jRh8IhH5sDHt6cDauZLVA5DYnycW3SYuMYWc8KuZ8JbWSUOltQ8Ogq7QQWUqFuqI
U5M9y8GGoQbLKF62gxybc3eryNSUaNXuSX6066r2a9k8nYmX1P5UbucC9RcPMjrO
91KQKI3T+RralxXvKEmcvEb9iAuvZFQFQ4ObwamsYevXBs2v2uwyEOZZ0I3CVqf3
HgHTsd5RuTyG+Zlqa1aQGK6vZdeEhd7YI4/DlRkx1wAAlo/R0KcPnmPuU2mOX3Mu
SM3gii8VjBS1VFP9u07X80k8aEGlR6cS88YftmxKRIfTgtplvZBZbZbp/YxOpBQP
a8HAgD60aDeJgzaXaCzdlR/iERg+dO+xx7MezD2tMbGX6r+4K1r4/6zuYnqpJAAw
ESbOppwK1z21CXcADXZc31KWdKEXRUJHh16SCbN2b8iQqrNywoKQ/TJMdzh62cce
7h+iokddYZ0XPhB6KGrrvbg0bTT2Z48iCLWsUzp3Tg/kwzZdRQYDnTpEvkkaSw1N
OaPjEjQ0cYpMR864WUP+AjuwZhFqwuURw0mj6U/nqqb+Z8eEEznUPtL8/mIEiAja
vvRbnIPv6gW7m3HdGfSONpjiCt+WtESan4vmZm3K8oxUJIMJdsLEKRD9xsEFys/a
YNAJFuNGosLUmzoVpoxpJqmzNQwpv5r71hDg48fLGcYTBZqe7IXxUOa0hD+bIotP
J0A7iti8BCsuZSjWxAG9wJqBg3baHE+LfXSPLFYtZq9sn41rWGyC2ecOwKVTUjOP
RU3kD14QCTg7MtFts3LwaktGuAYTw9O81Jgg1idbMsQ1cUzm8w35yfmPc2Pllt+Z
kUGQIIy12v35XnFFj+VhKx33y3l963Kvfib/6QMPSUwEZMCsXpVFmGd7kmK6aVEi
kcTLuqPPemGPh0iqhB7MPh2Kgv7vcPMZxuPYLGVjJFX0VRFt5gBmOZ8M8CIf6m1N
JN2o4wlqTr6sqslE3yHNZPzsCje5lqyV0Ixon1Xep4iDzN3uvltcQgOZUR4yp3Ir
c3IsABIfXL9UQeOmqZCna0m/qMhD9kEivF3vDINqjGMOh2a/Q11kwNmj1RBn5u6+
OjbwfL2pTVywpLeS1bcEZf4PCu+xNX6xY2kzIc/UzyikAjKQOBQ6reN0SyvkUYBS
AxoIYJomr4XKs9cr6pmKsz7o6FMe5ZfNM6Sm6ljMu7j+65+M23SGcnrSx2JoQLC/
Lc7NNC6jd2cvQrI5MwhjVajOvV5/ypKHEXT2jY0BKZ1zG/D4TDNhPlxqFmyPBBd8
xgtR9mieWk8lSnt24E2OEzibxydVDer/0G71OyW1WUNwC6emut9COA9MA2ca+5q0
sJ8lKEJ0PCJfmPKB2+VLwFB3f5mMiELfhTpU/Pr6FazTxepwJAyHiXhm9JJ4D83f
u10dmr0pk1f+AMyC70WZ+Y6lFgIu5VVGVsgZYY88Pe31lofahJr/q4/9ZJrf30Bx
ts/jWcC5h0aX5p9Z/4ZL7rrtg8rQcjpSF0ozTavDiChDDqzsaxhCVRU/9cgwJ3j4
DoAM3R4diEi5TUgxAsJEpgUZpuuPtuv3B6Vf5hbR2t+tUVX7B34IWQ7x3lXrD/Ny
3+f7JJQktCrx/d6ziGjp/Ck7dFO3L8WOiBlQijkdjYsRRs6HqL/kK0qntjwY0+Dh
0tZ2RE2i1tTsBrWkU5IFO0QXDOA1TRixiKw4F7J+WXF7DScrU7bLdGcATI6VL8eq
CQSMdtQbOCS3HbLUJI3RXd7kE+4J/aGsFUisyDJAGlycG2/ZMm7K5qY9KlZ0F3WN
idqzVM87GnfQNZoivmgntqqqJ60ESe77YF7YwMVItSVeSOzt9OZWj/phzedFqr2/
wF+rwffx+OHYEOML/ugkHEkKKBlmQ8mUoXHMQyCnLELYWhuG+k9gyikC9Tw2h/+g
UFruILyYmpp4BarIaRW6F//eFh96of3X7NvdEIdeuIztumEi2+wizTTqXGtcs8/P
zraIu37UXW7hBRwBnQT0wEErhrMe/MBkK6XEqfvX5/OjTNQbaG3lLH+qwx2mPxbt
gncqx6B0L8FJMT+4onCJr6yzOF47z4rgxcoR22j2CHS3qiJC96YzUIyWl/QtG40d
ZcJssUKEyHKls6LiiJSXIKPRMLOkXWUh2w8Is/H4UMDGh8YHxI3n+P2QqRWOjESU
dpLVf8dMk+BJdS3C23Lat/vn3Gu163nb2TRQdXlq7smKVrfaNUpcsGHPIZelxnUd
goPw/ItVLavhvnoUEZEYVaapDtM0Q80tEkv9U7vu32UQTh+hd6ye9S/ot6nS5P3/
GPW+1cL3WjOarB+pW2syA83HASdRZ/OXd2KzHBFhzoJiQHSxB9gKsCzAYz/SJNkO
N0vF8ijbUxop+dWIKMIvhZSLPS2RbJccXfs9msZJwG+qAN90Pom56NeE/5VI8IkR
TwFSUzT067PyxQZ+hm8DL0Rp8aGkRzBoA1677BTfX9ikcxVJ7L9nAa4So6lndy5O
52vL45uXcSv19TmrbdJ38Fyky8+tqp5BPIguzsb+lnHOOehY2QZQDv/JcT08VTIr
5uNtu71O2ACeKi8I+FIZa+/F4rcxtPUFwEr8OQsH30AzVPiiZF2cBihuVRc9skt7
WbQYXBZ5hEpyinlBKSEaJwQ7QXa8NjU9xwQHz25a+4Rpt/MYxCMUL2ckB86rVIXG
6e82MPNw1Oq1T58GzqIViMxHIC+eerOVRl+hqS44uyVJT6BLr6A8HDpLtpj5gqhF
1pD/A2FB6Ht2HekwJgBNJk0XtRADhwqV2cUD71zs8NiYUx7tCNV7077a9fp028FP
g8jGLTuKuqyzYBAUvcKqlIcIAfESreSQcGKGodshj89j35IHk7IAT3Vf0QPuB3Og
DH1jln+fp8QTqQvTP1co0ZakhJsYMqThMC6btXwpLc4swnJPNTwQk8yOsDeJmhYO
MSqrgoE42Zj/ls3jiX/T1QSTsQ24/7njr8kBinmhFRdcPfRt1EaICUQTU85Dslsu
7SxqY3RlALnCIQQUcMaHQK0p0IN7vdUYbC8IaxJkIpWqs9mOPFxplgUAv/M5FHh2
2gi+8uXX2P8royverNzBnnhTLd7AKrl4a/4shYWrC7ZX6ac4qo9n0AziwnXS65LU
PWWJlZUdYsmF1FfzkhLCqevFzIRW3OjKUPEK6uoWNFHykDh5DsXHXcFWG0FScpCs
kL3vQCu66MdS2/39ygRZgJfWfeJhwryEMHb9JWFz20742vF9rIwB6Bgqc8+oYFCx
pK1aYCJtk4nVIufBGol31hRpQwUeXjncBd8OQyTc6fifn0i/dyMtzlt0wnb15Xv7
bdjFgWPouGfwTsZB3q3ye+IhX4S2E11VQd4wsOWs8asbUCizsZQ0L9HCrg3hTE0B
LumT6JONDesg3cwA+0av9kOXQEY8ybzBOUOdQppCCgcEuL3uTfdjQ2E1BmRb4KAc
2kK4k3olR99eAP+wcDeBbvjWesXI8FbZwyTMkTJYGPj0Nrt4fNW4J62faqdJZ/sP
DL5aJFQnmcUAz0mrJz2Aj5V/8Nk0h0YnsiFGo743XBulUHsDbI4nSIMyaYdGUW07
uCVY+V2jh5gG/jMw1AItUfPQPvVdslWMezstKNfc5P1Z51SzY2Nls7S0nJjR7G6M
auNFRJ8OR1PbZ1h93B9idYlbN0mfiyUx5o6106/H60j9Tj0rOSVL9K6q5NvMRVXD
Cm4k1gr8pyRXEvnjJ84UMxRPfi1A+ZF/m+NyrFcmg1SL2K4t2lgOIBuyWYM7Hdty
dhVgP1G+uYb0/2g703O5upcHiC/38ujxR1b9xnBaWHx3/mdySBoADiy5nwyfNE4K
RydqKXOd3ZKy2zUbicI6EyrJINiw8yJA11EHesKnD64fDZfr9jPXV5HM1zGUkXUN
OAHL95ZJo8sSqJjgiPgg1tWIgNi/PT59S5ZfHTiZmw+n/YHocJ0qKUZcgwmxogxc
y1LeUdEZ2iYai0pC6QDtMhnppOb061GkJC4L641PWMT0KeXLMix6A/T0T0OwgZJm
3PoDTm9zXH5REalIDTRhFeuinvMt0wpFZzpMuZHAKhBu+pEUl+cIZyuFJz1Ao/vg
VHiD6INzdW3/oLJP4ueJjo3GUGvpD3NJ/b1sSyXjlqEDqwW4cCPPStT726AMVyOg
b19qxClmhAj2WR5tXVXdHDx01R2oBbDujAxmhyQulLIBu1+pQxheWQUMsiXgYWwR
TONdelH9G6xqFCP/pbqGKwpO8H7rvRkuG+AvJ1pbMCU+59wRdxAh3/h5soeSkYOC
0lT3stGrpX5PNYIBqUnrJfDicVaKM2PeAgGnh+3jzUJJYYcL1BC3XvDpY5uOJxJk
JPlZpgHhbqqIciSvR+ACwv5DGYO6nDIxYLTBEh0QHbU6BBon+LlDZ7S853tlZ6C4
5SAbHAqNZKh8451IXxJq24Wsu9iM4F5QlJmZ1jP6VpwDxGWOPJKF0pa5kVVENIh9
ZZnYS41/4usyaZdwCsbsKuOpBpdRImdWePlEUPCpXKTrVrSjYom9S9R3z3r5sjBK
wm+3VtgtJ/D2QmSJ9EGya4wZmzumGSj8P0+pSmf/T6Q+CB0YATjcsSWxjwAMhDv2
BSiWlDX7ynUaPxjab3NkCjdbxaoo90qXqr1t4xZCPDkWM5GslY+3IaUUoU63yGVh
AHMolgUZ6ZX+7Z5IEeFS60f4EWcaGaoJCcp8bDXL7jykWQGVqi91h/JgrLiGQtF6
XlH4blRFeFVYQPNLJiATytVrqmdbdwg8otbosw6moVDzGeHeSDORBztoHUpKfv2h
5ZswgiWo28eko6KIwEGs3+DNeklyk3QbrUyBXppoQxV8QVhbgZT3f3mLzlWcSHL3
HeCwNVob9j8nUFcvjKiUkCCTENVUOT/rs0+LasW5wYTwd2OQYPsGIq4B5c41F2ys
4x77YBLaZy6yQYhU494/mb61hjkj59D3+4IiAA6MLtFKyY94RxtuIpclJ7lfL9V4
ml6BGxWnbwqxTTvxkOOaHHyS3TAQhYOFbo0mKX1YwS481/p0usd6zyZBHmyo/TY3
fHHNKjmB5luYUPbwTbQ3qrTQD5afSNOQbvm/nAkwp6ZaRXHSNkXiduQoZ6skcqvq
rQWe/ZTJQulYJQFBPku/i4S47vOg1I+0/UrDKTPRNr4sbI45d8tDDL7wUoGEC18z
B9zJC6nnJnn2voAm8ka66DylOteQZy1NSXLbsKckGZlJTOR8ehxgU+tPzff5eTc+
0KudSITAXa1TIsIvyvr5+W5D0uQPIQsjt1Hz+vcP6F6SS52dhM7Gs+BDIoebPznL
x+XvfSBs7GzCHgFZp1drLVbhOE8fnTIE7j6hdXpJ7q68eEXNPaDIoRLFYozyx1wz
8XRCaR6+UDBIohJvN/eSnQQf6gMaq+rNUR4+7Z7RrllgcF+P7ovWMQxBm/KZ0I3B
J84QGsm3CpXvkUOp2OlYeJK8yh/jqh2FYsDgaRDJweKpcxeb8Ofhlp/NB4WXaRpP
x07tNKQUbdvT9wA0LUA5qIwn+Mz+UAeYfmCB/SurM5OHR68ejFy1GtvgnQRwxHaQ
Cgw2OK8sMgWZD7GBJz+w1k/9wk4et0MfrFfiLV0XRjmkWB2QtMcwaO/cAjxnczwC
fMD9ncxWJtf1WEvqgDGqCofuCXiOi3USCNuScCFYGG5HGmRAM09A23i4nxWghNcZ
HpXC/ZLMZ/am0AySDowmL3MMmTfKzlPrzzwFNZ0teE02Uu9k5PM7McTm7gMPmb0r
Z3ziT12nMuy/MEk4t/GfXD8fw7FnNfqhaFItxam0xEqhYAkAybRceyvtBwGKDmuL
UxVeUOnUMh2S/sjAxTJyY37IKB2w0DsqhOge69FZgxHuPgyqhY9qI3V+wWGuOb3Y
NAzIZJnD+LrGmlK8ccEVpcANftYaUttoOAGWjuvLT5Y3c0OlcO6wgTmljDw3u9KO
+2DqvV8vB0FTiYVhYKUjwDjhP+AUlfjEuL8j7JABr7RlCGmGF7dL48s7aaGgUnVw
MaKP3s3B96D7/mMwQ1gTVTLseaHYZPnOtdCP9+OQOtt3i3oSXfnH5f9bJasQ79uZ
k61iVOim5gDCYvUQruANtALJZJRxuFcJrL0bxCpM6iptPjPUhh8E7ZLkZNJkk9CP
F+1jVF3+7AGOX5xHTnsuwUj4x77DPzSm7rXhNa94Pn1QV1dTXGayaT/giM4CyWzu
NQYQuKO4ObEmvJ7Zuomg+8SJ+sQ1WZXhccZaTiZfDBhdlhzaxoeWe5h20cJWEIvc
USWkV6vtHXyL6COUWqaI8RnDj+FJC7ovxs1Upj+05DFeJuwnA9c2DjOEZCmsriE6
Q9X5cPFkBqCwLBDxkXwn8ZJbV2OZbAXp/CBffA0PiLEglr+ORzw6uGciDQ5WS2Do
tfdnsvzk12PHSVRUW+QEnXOeTdt5Q6Jq2v0r5Wx8W2p03OVD4ChigDC742DHxSwy
83Uan7AI6xZhKKyX0FZXR1ZucAK1ULfmAaS1f7/jPTvbfXNbQpzkHMNiHyWHu6+5
E02RQjUNe9R1NMAtRxkivkStO6pF/zMCHS0dVi5TCEwBVtI5gBZcx3k2xEC93BI0
EPI5JxszLabYxP69oTUbpMwjc2e++OOyh3ZKPAHXkRy7PJE4uL16vR6JYv9ZYgo/
Zo7WVyT4y6E79mE2YmiLdvHklBMMi6qBWzJ78O/bTnX7iFX470nKYqfEJt1lUVkV
U3uqb6oZr0HFFmh2/VIouKhyENmrS3yguVC3uvEey0u2Lpvv9VqdngPld0BmvnYF
fe7WpGHY39j2et1VK4GWzlqMFmYNbqIaV/fsiD3uJtlQUddqqR4Z8by01YlsnOu5
D6AQFbNei9LjRV2at5jIb6yI4BeOzVMTEMNNLi1MaUgrepk2QNK+AY+jkTkpFngM
WViVRd7yh9RYarvV6nvOFbFY0GtSd/aCYg/Goxbj7UEFHM/19v4tqVjo6rVdXB7u
rWvRVvPr3mLgL5KR3MoQ/pdCiP2uPTpWAAoviUxsCTD0D/K9YGW9QMNcDuGk0/Br
/bGqPZKoFM3iim8hIVBsi4yHzWAK7yWRXJ2Ch7rv32B5RgRO3O4dzHORg4IfwIUj
A+ZTQpDLBCvMHEPYRyd1LGhL4abUS6SWyewyJlLHZxZi51lUcbryZjkMs7HB8g0S
6OOjE0gJ9VUNU8ouUMU1kNztNZG0V1bjfIltDJpfBPduumdH6CpbfzEdGIF0DTUF
+GhCU7HYv5KoWYr6VtoZwJxx708kDsr6AeQdDyP2Z7zGLjd4clzwjyd+N//4M+jW
eD7u/YJcrayQmeZpVBd0pJm+Skkr/eLYkg2TsgpiA1F/nc3z2k9/4LM/QCcDt47n
KFAwC3h+K08vnffgfWZ6V/lE0M+XUMz058a84XqGVD28/FuCxWggy853PFfw/1p/
CG80I9kVVCa5Pm2U+C28RubZTpLnR+B3IziaAr8dieVzbIEtuqi0sTB99/QjT0sN
QxDR6p22lw877b3LFLed4sAzArnvhDCpyXIIwsscuKaPW0KabliwVbUy9mDlQ0cm
Vg5fKg4nEIBYp0qkJQiQow8zxdUlFfhO/Re76FuQD27KPsT7wwHO2MXCUC5706KW
x7dssVhP1s9il+Q7aE9ZVPJVQXolzcay/AhNje1yxUElPis1ApyMnxg2cIwE+xq6
lyRj23Jh7w1eZbm7T+p5H7hcAIELS0pLaLbC0P4/GP8exYdj3TpIvsPX9g4g+tmT
d1dk9Xj3ucQfaontU8ZBb136LhuNIrgtqMzIiGh210MH6kYpoSriko2CdCZ9h6f+
QZjeGmOZ8LcslRhfg1VNYIamaee8+8WwHTJdAks5cMgM87ALCgMqVNKH3Wpf2+Bn
dVK5Lg4hvrhuq5RdW0cWrlx9SYuRx59n7pwEae/HuYbBQaVaw3aRFZ1glREFr5mu
HE22OTSbFMNwC5pfP+dphTxw33LhZonfTbpmkE2fzVvrGRyAHLrQbcmC6D1DjnK0
JeM8cQ5tTpc6FuT4xB+l34RHeFB9+ZK/1LyI0Az9vN58lxJXp6+R1YYHb5TQYXkr
zUSYAfmvggUS0Lr64Ci+gG/dEQ4SfGYh7vIarUxamdUZ/i1lZdazqjkBypD4YfK+
v02m2Ng+5cEGD1v8nWcphmhIpWb5HgTOAyYgvO6/VY6iw6KeZKblSl/PSFhuLjOX
+KWBQPvEUozpAUMY8t+mpyXxwJ0oxRw9iOc5urZyTS8kX023KLGx2OhHMOVpuTDn
mETG3Hs5lKq2Ky1Yicu8h+xeuY5nvfLoLXvY9oYs9GKNskWyJcez/HjzkR0G2uj9
12G1n6JJ+rAF7EXkYY3GZEH5wgzzq9/hoILY0rtG2+jFOypG4W9Z3bhy1WmKfVlx
XL1pHCDSecUVYg9vDmSpmdNBBR8Z18hFxwUaddqPtA7aiWS32OE53QxCKanAxn/u
49fX2HtK+i/IH6WUDCWY/Ueh1aLGJ+Na+dX607ePvmZalf7esjRgTwft4YS1OVkd
59wfZthLwyGuOK1MFjQbHkKH2Dpn1KmMF9j/ahtYUjIoZKxb8Tn/cBY+U1Cfj/6J
6x34UqN5P9Fk3St1laZFaevp2AksNTVdF1+jflymB0XrDRnLMu7WHkSfF+Qq/xI+
K6cj1UmtgKXnD4jm9uCHcG8bnlZ0XUQ5wnxH2uxVE2RBVrCcXwzh7VVRkLFqhuC+
BcR2SPh34kN1R2iqNYjk5tSLTEgpiSgRJbtWsTucDJx80e8m/0m6mInLFkEu1NAv
Vb920t8F3gux3nxzI07xsZanrbisK33bOulpwfXmJU9rNyesohHmfPQ7yaQCCg17
5FwhyisJZXU3CY3vPYC+v1vl4Yp1Q/qDeo51pl6GWjHe0xZHuTvqbdIg0SAR80XV
uKQjroe322RfHBvOu0/1Sjida57hQyPuguRt4UsqZrGfj5eBFkhZRjj6SAUg1uzf
IEve+a86y1tRTzZyOgV7NMZ/Xj3DGII6NAT4iUazeTEOeo9SxcmbfQOy1UKj1c0i
voZvLEQH2Zh8Mbx2WjCzrEDURCZYziT0ltlZVWsXLgrnXhSRnwywScIb3evO8owb
+S5KG41ibJAcc57oQLGTdlnD6BO5x3uN2r9ycnKtA96FWJwxXfLJwvXsyJvrURa+
Uk6TsHQPbVpznpqCIH9IYbPesxHAl2pcimRPl009Wzyi6ur3RkvTOFVZaXaXGmVu
/pM1wM1uxR3N+MbXtWRT4nVoLe2gTMHgBmJvTTOVJDlX6W16SZO1UllZNKLAP2ev
62CVrB02a3mF1lMAWMSjSXRCDy7/iwD0J852YDzSLKlztK1DYqwHZqfVZyALL4+i
dO1UiqwnkTPZsq/kVSCB6TrWV1iKOe8m5cYcJ+XD2py1mqE8yqYpL5Z8l2778da+
hPRVBq25V6Mf/mkSxsMF06G6Z3p3uI5NJLeeBL3A0ty71W6xnjFKCH8vFO2M//Zh
khYB997M2K4zaaAgiPhndeTfLqoOmYv+YJTcm6arbCzi3z1WPyYHrfhhx2cVYQug
soyPzFW4MGDgunYsfhbSn54zlzAplipH52QULvTr9K2CVinjUS3ZqDax9lGCi7Bb
PJ3ozzO5MwFn28/NqF0dIni5JzmfUCFJQXEvIX6zxxTqKC1qpNJpXrYMiWwsG1hf
48BCPeiT1HtDAioXB1zo6eSEULK6Y8lJBpQy33o1shhrC9HIUmAYK/C7iuQE9clP
fNI1/Vwp6CDa2fHGbcze1tHM0/JllJTiWweUyqSO3ktoFfpTA9vlN+eBcr5bFXir
X4JGFQaxOC38/ynubmSwsbN4G96/x7RBPHTtQNVt6QOCa5Vj6efStv9AFwtarioS
jQA9typcOmKhVarlZU1EqjfTPL/BwDdTmOf9aoi7M+ygIqTITuZRwPWNkeGhuBGC
uGUEFxXBwEJfJquIwgXg/dOxj4BRFcl0wdOiR72hsO/7OPW7a/cVxAKkNxU1WD32
LAROY1NCz8+oFtE/hL2N5wvT4YwTH/6Sf7JmfqAc0HLr2ED0VeaV95l4miyadIcd
Zr2iK4xBcZP7wmXS5aur7Zq0HrRJu1y0iLmHE4iJ4jLg+Rnwl5Dbk9WBnZ5A4tJA
S9uH+DKex6Sg6BD1zPRFuGrM7d5vVbGuCxWRwBJFC7Uwv+7dxO1sfh8YYMI0oeHW
OAU1QM2BYlXqT6mla37GgZtlo6RLdyV6iWaapDjlVBHyXfGEl9C5+AYf4JUW1U6h
RqKB/e7q52pdROZZHop7tVHTuX5sUZ3lGKyjDtFItpTHMpJiidZr5oqGY6qHzqzq
sRps7hHVMdIIgIFB6GO8O5JFoIdmriJFBOvqghPdfEUMSL4TceneWw127EHhCypF
AQ6pQvpCnbcEEwfy3a7rvORRnT7ACq6Zo6YoezC9Fl5rHP3gcZm7fVCowJud/0/x
DALs0q5Maoem4d+TIh08T6hoL3jSWCDyaGjZnFDhAmweq1POV/gO6TP8syRm1QXN
p1YubJJDtcwQxMoJ2duSXK6QaN8DF2ceGCZGRUxAzKp84EjbDzUMEBj9TZbYEbKn
Vn3DEZT2XFKQTGN6lsg6QWajrwWanx6UyriBNzLYX7iI8GXVqQ+2OGzUDdxtMJB7
71Wykf0NDwTmJ6/lKWHmWJCD4rzKjMDcOHsvAKqHSbVOlUBsVLpj8ICxLxgMbVGa
LKoxtA5jUdrwZRNtrguUiIEVpbI+8oLPnGS/v7SzK30hNFXRSgBA7HoucY4ne3nV
yvGCFaY9iMwQo2iIh9pBnrR7ml7BnQ5+P2KmHEVb9Aokic/XQyhaMZl8WGbLyiik
TxnkOJeK4+jCKcnEG3TCh7MpdNmzaaPAz67qJ0wlVoLBaRNZIesA/B4zZes7MWUT
S8MnDlh9b438FI3XgmrEjtDpRVJmjBnRg5oOWhwbcAvc9dZotdhUG5tk+e2R4fB6
Xor4dkBBQI0rROEya8LyIRldZzOjQCIvZZLaNyO7N7WgowGF5jxYSE11sm+PeMvn
GoPMBra1nsrVy/hfNtZ0ehyb5pqYAeuLBcngNMiGiiLDw+BELX0pF5TSFYv93e7h
lQertUk1MTR8QNgOif5j5DqjzlpDNhcfiaZzHNR287yDMMIYiptjTVDZ09IunZ7m
VWBK58IQFGIdxT72H0uPb7Sv/FjrToP5coNFUM1tFAy8x+/lced1Fic/McyOwCjQ
G9B1XJd7I7/e0eoVxvcmqDlnv6lYkZgKrnyrnVxnjMTF4zn6ZuU2ZvRIOqmO7OHj
Vyhrbg6WeN79nxa/cfkLDcF6x5fIdVW5O8wTZkiNC/nY4bu6OyZ+kpjOpQJ8Ud7b
Ua+iSkvIBiOb4dLrGRz2/yEofrPJZ+SKsCUO+AUn33J1sFJ18SsfMkQH9d8JvAtY
XXiU1owNg7eX1LTocjFCqMsHmREQagr/+uzAGboEAgMY1m++3KVm7VUxbe2Qloiu
cW8RS8gJmllrQ9fOPYyy8EZKYgk8BqzFw79z+1emfxsG3A0NOriqE5vG81hCA8zS
XYRVE44dQrO9kHRIPnO1mDOSvuBXSiOKYBBRn4OI02qOaeK6gneDwLTq7+J801IC
GlOn+BIKIBml7Fbuu2ZIzUtPxooEEkvs+wVWsydIFz7enZFmSKUBVzv5EqRR9HPx
tlNxtm33cSK55crvkxt5cWvnGqlb+UL6wXEx/JokBx97r/p3s/ORB0/Wh+qODYHI
xmqzn6EoDGmheaAYCsZAJqDXBMLnIp+maG8hkOEZY+Nz2wKCLtSAo7m8kKNw12cs
XUOjECCgqFlVw07nh8kP/VhirxJNkqwxu2E2FEH1kBrDv5EpxFxf/dUhkMvb+h/w
NMYtEChGW894G4J8lX199UcYHGKMKgLMsouiVnjND9TmcLWxxYXUlsjfdC2v9lKN
tstujgASM06BCofWDu+u31fP3yXTxZknOKvu7kJ2imabBouXU48VVb3xU04KaGdS
cd2AzYyJEF4mk/LUX23qlswADvoU3Cm+XcJxd8Vkr3BF+QA/e/Pwfm9D9GThZycb
mAonYyi1U3VL0D75Dq8EfMoxzFOA8+9/7aIjamh9fTLj8kmwl28Zd6PqxeNczOuJ
yDtZB7/LryqhU2QuwpPRliSuiE6VeY61IGqk6xOD1s4dhWW96QcR1NK8O0kcrfHb
mH/3Drc36rOvyjWYqMmYQbk0WJ1CO5FkPKH6vheVOKtiXNxpbpXLc66doZSBo6pe
MrX6menjIKLZzjcWyAPmYR+mqqmUfiQaHpOW7OKmNkBTplAwue8vnlWYGQVfrm/A
oyObLKr9OTQbcAmOLatB4A9PF0SgRpoIqyGDFdvtos+9jHRT5AUxBmlkUoUdCYue
3P0syibMmAfHL/keHN9oiJ/O1BreeEInhG1SuqhPIXPqo8H8c2ymdo+PHF1v/Z3N
04Mz37gf2WtjX404+LrjJMWt6TVmUvUfQSKONlmx2JdGj3DTTqPoAoBFIBUZmXCv
EsewmN9BjwnSiEHgIeynHMNM7HdTUAj9nT+DxP/DEKIgwXk/CO5FF7sBX0Zg/Z7v
Uue5XpXItuXY1K1ATXNM30ikuQ6g9O/H5dp/a915o2wCqS03OswnFgyDE/v3XRjT
90YDrYdJfdoUXVRlKyKaHnRboEMbWGAYfKSmY7eFCQ9bCdWG0RoEyymeWga/d8v6
fx1q6hxC7GMoHMAJkOpb54sDQ4qa1Nkm1pbc4QXA1YwwBIRGLVNwrolz7RlpMNaD
KcbmAWtNC63CzILvuE39AJBFt7Jgm+798nKTwFw52VEN5gJpMcI/UYhifRA38WAr
O7jpx/y1G7QmaMWNEaAJZUHsrvlJO5EhCDsLVpwy/onDumi7HDOUnw5lMjj11TRb
FgM07swa2cw6xHPAkCVIvbCyIWg68lUyUClGqhHhckn+v60NT84kmkchmmkUSQPu
YmqLkBixHNYLJ8T8mJRbHOXwhaeVO+gNOsJtSHsqa2abLXfuZDyKpELBY1umrNeG
Y8vf++SKP8D1h0ajd6C/g/qiglW5O3MCq2tp2qFA08V4Z90U7nMJJRpgtovIBS76
J6stjMebI0DRaQ3ZGD+NGJfIio8mqUiJ4Wx42fIqxJk4pc2VdJUo9kfls31k1iN7
meryn+1WUOj1ifSy6BCNEeSlc3WkhDBWoXhL/O1SuM2K6XI5S4W5OiC3xeNrSjQy
kbxGGcIANPaLDE3Ct+OzVc3g3idRu9QZck77nmeTo2tqyZsrAXzAxv+oV6hgyvR1
Y80w+Cxy7G+sxNOTzBVaFPDG7q2iThIPiCLIITn6U4AdzOA4Ui+snb7f8w79WIwi
1E18TZuYfFpaUl8YlLycyT5fwUekKN2+P3ClzZ/E9NCe5yWMsEHzNBzCTYVUi2Kz
S59x2F5tS59590IvjKYAUcSuDgl/PRarWTsIKdjuHqi23Hpvr3mHxnHwykXDKlh0
HDmmyKXQKRjNPDuU0lk/dWxspfAH05pgJ+Z0Rvq9cmkcQcfyxY7MSWP0jCPHwMb8
PNNnjzWV2CL+UtlYGUwUuITrby9uq+FuBdPncTCVlio12qUCA1vRFqTQl1rkGlvb
cgG/zPxLnmkhqWwpYuRoezmySG3Od6KkBzi9L8gpsaFah1gM49/0HqT/2lhAYM1E
vOg6vzp9n+jlu9GeXzLsosQBl3Xg8WCofTur4oP/gHMEFh+zA/xz+id/erihNoVb
Nq4KFrkQOR74NhB+3J9OyxEPoc+ZBDbttfAoJ+5sAIZp5eM6lnCySPny7HuSIOYk
0zYW5UJZhWDfSHpX2zXO0fqeywLfFiHuoHzE68EnqRni38qAiGOOqNa4rGzI3TZ3
6jsWlyFA4jNn320+Sj/R4wMBP0OLImDw50OTLqTEmeR10El+/pE/bvO5zTAHBRoK
pU0RsyvOkKGSrNfJ84IDfEMqtoe+fFC+JHD5VSEggfSA3bfot7uSfd16unMbjTCN
m5A2WtcJ04vuNZUZDDdn5R3X74AzutBM617al2nporOJkUNv14ZAKFbooBuGcBC8
r46M9sMBTwNfX6DXQvbyGVDQsEhKNp0Zsu+kqODhdl1wNctQrXWuZOSU8LdP+CIk
pfo+Gmumyp1mtM1LvNSUp3eDrl9FL160trxdAF7VtT6COiiVHUGGzFU4XPBmd+sv
oZUPax6/CrePK2RS/Nb1bdtNJIL6nPsEOzSNPqGSorrlWqP72cijtJFZXk2lveMu
XsPbQYjIw6X18KPHzqu9YShvmbVa0QxIIVOaUNCng7Sdb/wYz65VT5EZmd6PWgsp
R9EBuxT+K+AddD8dUztmJLqfgEd9ijr8DuDBewDgo5RiRN4nmcd4uQG9NzPOjnaU
zfpGm3MMwkd4BjMYpkh2pjE236SAZZv+3FRhQW754vyjtaOjiuIarNQdVG79aSuV
3x/ZtO/hrifOKYURGZRflQ2JnrT+8KVb7u+ZhVVa8hmNoZUx2LGRjSkSIE0lAGIP
Xm9ltpQMhy5zpxFh+OFaGSmwft9p2SewM+JgFvaXFnwnSxgW1hUR+jNMpUxnlMD4
4zVff0gP6AaG53iiS7iL5eeYgjX64AqoW/ke0eX48IYMXlkZvA3LojUvyqqbBy33
BOYSRX54z6cQ8sYA3I9I8LOpRpQ5tzZZfZLLlxsDyZwpeR4lR8l86e1BdU1jpk7u
7A3myYjmgrp6DmRFT9tgmcXCxxuRgYkRLvfDzQDBKLWIx4FQDXhD9iCKp5+lzJbE
qpCc0jTAAxG9C665QpgCbgFPD6r5zMcU2yhE8KM2DJlyx9+UwyJ1Ycvjonont9Bx
duwZvToHq+1OkCp+zkZe0QtSECReRUDQCWWxwvLS1y2w/v2M5N9u6Zyf/QnR//NF
OyFmai2mO7JDiX5LjYajRuNEmojKgTN60vll5n+zNciH6phCmTCa32AyRLm/TJs3
PBv8denqRjyVe/eS5oZdqi1XjuXCR+u8BLUNwQlzK+1LNimu/fm1KxWbl3xl/UOp
lfjk8mrNiMaiK+DDIZy3B8Nb+Wajt3MkJ5f7LdmycBr3mRK5DSEwZpbTpGdZaFpF
jroAnFRwd3064lp6iRr7pnAT2rewVUjcdhTi380HY+AnT00ll7KhcRpLMCqe9XhR
cPP+SDDFIqWyqJoRZxcpDSJKrJNvilj3nkj+rXYZsZ5QQaylyZNksdxLfqgl4AKL
onzUivNi/27/AVfUhCNb83aJK0HCzZIjwpmBioeflcFJvikExDePPAWXfumAOpOC
Kii0la9ts/fyyDLAvqUFB9J4gWtEnSPc+dh9RxYrXZk5vh68s5+CkSK8uJ8f600z
Zc2RaI8uDjnukqJVu6Hvf5MApm0SzcYd8Ym43tBW8qUfNqZjK/ejgWGN+PYe/9su
XC49EEXdtT0Ap5DFKwkTASEoDChx8cGKL0+TveRXjMTW1xO/DtWUtZH1/MEMlnVN
76Xx1FkQpLq2QBnAoNPRW3athxDWK+80mYl2kkRevXej2k0wlW4n1Jr53n99dWJ2
OxOPa7YQ4Ab5CfrbSWeZPU0r7GFz47HTswDWs4w3nKpcVT69Bgn0qhbunK6HB+Sv
nNFt3zq6PlPrqgY3bTj+jTe6Q+YWB7tP7HL5ht0NuxTm4wB4xOC2/2ONnAxNWITL
MefFuLTHEi4ByW8dNl3uubIpDg4b0db0UgPFT+/RU09XciMbwecu7Nw6+qrOFeg3
oqTKxbq2mzjW6ReFBJbF3MnMV37Dv7fTEzDGDy/styTG75ozMm9tsu4YZeHnaI+9
y7aMjqaj4UFi0Mbe/TfCQYxaX/HTEIRaFRqk8tJYH5TdJzwWvo6LdSjvYSel5YtG
p0INVZkQhj0AFpUiepjTO6HsVS+OOsCGu23nyBW2JYzwhXNvxsRLDG+2cdPGxSmU
TmhZ3xyt+l8dc31imRi/xyglCiQN1lDzuZOSmAI2KwsSR2wNpILU/DdF+qnVz1Q9
CxXmHlqqP6de/YVjxmdgBgOp10gsmJtdWrGEVZa7B0bbiOhbaHA4fchUgWBkShvz
k+DMCiEgkv2VKiJyxexWwD/MUN+yfb5li2LLh6+dOfdqgO4fhqigG6wjXfPFjY9P
0BtUoBbHwmM+Ce6E5RoEHNpNAPg/mKAhNoKLZbTPadetIVOtteaglGvbVK+9R+b4
Rh/PDvXNWvAjGBAlP3UIlspmylBBCSl6I8sD9zkrU5MtlSq20qakJHy2yW/bn3QB
MH50nepTJGGwGTIc1MwVtQM7Z2e+x69OI3AKEfDlkOAKcRHFE694cdM+HMzblEs9
JEIbmF2CB56yg/iUFO/VvOPoHBWFmruZGlyH/Tpw7TZGOYKiivhuB3wUvoNm0CiU
vFMyXpY6X8cMu5uzYcZU+s7mbnvhQvHY2oNfODqJERK1hl7sAJTQ8y3fibkNq2aQ
Vl4Ka4WgPEGYkMeTlayifhh22Y5MU3v1FIk2HwGkm469q270rPzoojFzqYAMwznb
QNkyKAkYudYla7dPW8tNVDTyitWc/PbkpQhvkuOnph3SNrhV0t3NX5cz963jcEds
blCMw3Cc1txy+qzco/pU1z/scyC1+ZH4RMJFIHjWCj3GbmGzvSJomVkKR7bvl59s
8ufunOZZfNpB3xp089yq3EFYh+Kt6lZj/TsqG3XMX/DPQvLBKuPRliyF8+EqrhTp
g/v1P8QlXsNTsDZebVkD/9/zJaCXDfiKkyEHzsjEiXEh1r4FrGGcEVNji2idj5FO
b43Ir224h+D9Akujqo6tG/lhW/B02XsZruWYHZyt/zymby6vR4V/TXBn6kmrgQCE
+ysBaitY8z8O9GaXaJZK3m+D2oWPqvbaLhGgKG5sSUHWvozuCLyIPSjB2FXz4fXs
aamF7pmiXDX59638135auQ+PLpMn6Uz6yszbID4v3yBBY4tBESjg6CcgRewT/jy6
NDr1so8wtdX7XztLTaYL5X8xlfrLlIX5mJk86ZBA59EjBf6v/WlCRPdpz2soW7St
1aDiFqN8SE0/qrXLyQwaYvHXd+uQe3pxBTH8ERpwIPDCEp71BkJ/rNTzrpz0hZWN
cEbZvQ2CLscTYeSYeEa1N8u42IN4KwWLS244Qkve1kXEIBMCaJwtjBJuy9SSw9dd
9/57B1YcS5VDtsJFPzLW4wTphCzpLuBh/8EO6DCSdMIjicSoc4d6PILYmT5sMSsp
vIwDEThwVxjCvPMjrrogvDpm2pL/zRhjSpS9rSCiQoEp6KXSdi+cLrg0xnCuB59u
DYALEUms7+pR1wfHtl6/4CcPo7fSaBZN1wqJttDAxPPtDF4cTMcwQrWL4WaBFv6y
KaRrQgVbndxIG+nTrmoT0lsVSewnjBEwf32J6KWWRzEtQgGcvjo1e0/04usIH8Md
g82Urc+Qq04OrH5hVzotAEhHp69xRN88N6EeEPEm3oTrgtlEM0n4NCnU/VXJbTAB
1T0WOjxB6zo954RWQle5vxt1D+e903oV78GjD+iFOAKMU63xoAjNOVPRC7Zx7Mp+
vBgEkmJ3+NMqagpijM8O9Si9ktekHdoPIU3RNhrRlmGOFCW/zKESvrGFkVPExxnx
lwux+PwicZnxX0nc7WO0TW2Rh8wzyC89+WvQxdbOcxhWcUQer7OX7kl2Hfh3nA+O
hD2lsxWjkc8burkOl02vpNjgn2zqonjB/1mtA5bk6sulsnWCU10uNYwsH22iUnmD
B3k/VuQIA7mmU1uHq0xVdTT0kTRUyLi46rpn5OfeCMTSRDZErcqUokfmkXYRwED5
5is4imIz9qhfRyziFwb5y9SdKM9o4aEUZpb2mheck8zwtFAV83PfghNt909BZQIV
5kY29xxMjRbv6mGIkqWWhLjPN/AadfNnqyQdWxnY7KEsi+cm5tLrlShvOAc6s0BF
u3WhyGnzKAsfJnq1HRbp2QjCDCmyAcf8J2uRlsRRL7bluRyjG142ZpBTl5F5ec3b
guWy5zc2acrC9HYAEItCgbxxbSkz03ZfLbg5DeW3Pe1bRLmNzx0lNnULUDRZVnz5
QKAeC7VNBiinEhibhjOdNHenZXdINQCi7k8Hue4Raah6aqlCkZpG6SLVMW0+TNyp
bNRfLfvenaOi41sIM4F3Rh7Ecuo65+nky2oZPCzCy89KVxvzSinA/y3JqNKrSS/v
6lszLyWjcn4CylFUfAoX/HDWyneoW3ZjvnDlY5Vayowt+0Pp7zRzi+ounG8mV+ey
tL/P4dXFSAQU9V7G2h2PnUnvwFkRAXI889QiuwyG3Lm+bG1DwQA3cPa/GF3jTrD4
Tc0eBTD51sh73ipSrxI8pDtZ3PsYJtC2GbJUP12Y+U/GmI/aLTdFcn8+Xhipbvo8
P5Bznl9cEKgklHQGoQ6vxl1qPMwFCKkr9nHZRlxm67FZDtukwzJqSPgumvarkePc
YS6B0Hom7BLJj+zqcyDDNm+LWpSx5ZshFX1mcWA1k1ZMv+PL1nuRMZE1ORjjJnWD
2TUPU8DxGUgFHCIv+ozL74oaxXQWVZkKWPWjG+OF8ZtmBlZ5j8f0mc+5U5o6SIak
XaBEDUIIf2F94E7X9ALBJAPGdEr8o1dgOz2sLOgm71dGkKSe5AWwpOoI20k+oYTW
9Pgp75AZnGlonJqS4sykDzIAIX2HD9dDnRT+WAMTOpw4/sL88tEEd/afF1eUQxBr
RA6y0bbZlWh/r5gBKnsIR7gmbBGLsSIudGIISjSeEJPmI8XvvnPfHGdTWBhaEkU/
IzZNRHmjjGGLrgJdCKkq1PvxvqL6vQwLDtNYKywKaXMu5UJYR14Q6U4ZyxGGaUJH
fZ3OACy6zt5yQ4LrnqoEHk4nFja5Wk8sypBp9zZZaTI1BC0yuKJQQhdov56umW70
tBTYufDwCujvlERh4JLIaQyaYX/Ob/Woem33+Hrl4ylHD9PbCOYq3yfKDTzcMNBw
iITUFaU0V+CIeMUzA45oU22LkuHOhhp7+sKZCYVi8Oe/5jaGgQxv5U35SjA78N2D
zD8zOJqwH5/wSspbBTN+mzFQqxEGfCbLLVy8fTrsg5vW7dQxH4JglG1OILT0KhCJ
oc7kPlO0TCrqOYqYao8BYF/OE8FOf6dx6jXYyxAPpOzaCm/D9lmNUQ38N1wUPtx/
0+PoOQVtUCb9XqpHS5NiIMM0zh3OFTi4bx93W72Cd3YXvMW6l7vqM90ELQM9zFMn
QAx11EqwBYmwNKaBiJBd/DOMxEOXMzEnxNHWzrZKmm83xjKjNv4hmtKXUJ3LuIOg
FcK20Bh0PW4QHww5oMk6iNi0+bgV7VAfFw7rrSLDJFYsHWAN/6fOT3ndYdcg+8Dk
IdxZv9O0pHUgpX46Bldv17kz2MppqbVHz2bV6ktMdkNz90trXVMicS+ruS9W9V+r
FpX0aLBdyCspQ90S/aGIJKn4ZE2UAyFe7UnymdwhQiKbBqktzEQxZ1FF8ueVT3pA
CMQhXQDohbutJB37mpM7CyMISNrtyT1ow1magpPpcWCyv8D9KD4QvbZbJyLDz06W
zfBqob+7m1iYEcP3O4jHeIILb3cZ8TjuGcZqLh+Zcu9DO+Hee3lKlTt5VNsvHQAs
0mK+O5BOteDZpHST6SsjSgonwsHKkATZtShMETJPit0ERd8F9VK0VMWb3dBLpf8w
w2LsxSar0TKczJx48A2R6DJuFkEyi2TwRQNIHc7I7SKczsz1X+7sCz18yZHqOcL0
Uh2KXZXE2/ppqgMZo5HAUUHZIPtZ4X+7ZSO0Vv1k0xMqSxFYaRm7XkFdKAEKvYaZ
nxfR/MFzdX+EZcHFPo46J5MZl5AAv6JJ239JlXvVoEpbfUH7pjcA5oxkFosz7+qb
r7YAqLHm3l6b0fwEZUtEL9AkCtdYk6AA7FCjLVvV0zQ/LrvrxEmrXS8OgBVPdNOu
ITkSLIQzOITBgucP9OLN/kNUYdV+jeRQUQgRl5GxUnh6baISsgMft7YvDtanvk6n
5ZwTWEhGHYeWdnnSXM35OgakH7YZGnqtwvbquYurJFe4jd7xF++NTsWYZdX01Qld
sQVdwU8zHr5Yn15k/VwI6PyBXaZJcj5uEjn8G8uUpA6dP6vFkkH70F0TeZl3ei22
S3xS1+n4qPRW2QBu7exNSj+Tme67g1Hhtt3FOYY6Mwkt67XJvwxyh9BJG3Njb4rC
dm+rzpJYvcjZxYg5vEOchXi5fuC1huOpGl0A5NVk4jFcNux7Foxg9G6NpqQCHKhM
P+z9UMkHyKa7EPnb6c5nzj5orMEeN5ih2XnCX+bA5FUfDebGXeAZTtQzrXq3ZaME
x6tWaJ1WNr5I7p2zgbTHoDdRg6Lx4my9SOAmXP8jFcR3l6eq44hMckKMd3sQDLbT
gIxYuZZtBI951tT2xtkmsUaOol3WHNM3wEL6AZ81BFcVvRDFkCn/DLlsgJw/nvv3
86j8bTCmXVT2vx1Z3zTmtIGh0SwVe9CzCbTHtdkpmhxAFuTw9Bf3QdGaVVvzVfj6
NZTRgCnKCQuk7ALulIpjbOzMb12KFJJp+MrZxpNdSkUl0gjfxCOOVXc4MJnV5Fwh
4FRXdBOoGUJSZkwvuNvqbGqF+/0jr3salGX/Rk/oTmfVAh9WZ5jR2O3P5bCsHeDq
WNurE/GhaDjLi2xT/QP9obz0rQSu1VrfJWw4PBpAowfk3ByrkqEzj3Ck+XFsrW7Y
4S8oHHQWfr8zxJDNrDz68Kugcem/LSLuuDST0OaivpE0tsQjlDkRsTjvkIyWs75K
tFUFkAhPyXEAT7IEuSCNoOju/GCQpadrMenBSNK+3Fzg8zy/lLUp9obHaIxTxhT4
QW944B9fpqWc8yjExP/uc/JxZrIsHCNf3DbwZgiHmTEAV+XfsYqaRQJk4ab14yvD
qcdyjrf7TkN6zcmmOHMmp0ReyrGCN62Q00QHA/RB0KprCuX1+CIvSxS0kXeljLu5
aWdxk7m5U4HCK/WJXph9ddvWojfZe+ised3las2eXMY6zoLbTBYLlTFO1httmrPF
GOqPTMTxhkyOitoTDl5sCmi5ovoMgWN8LXAIHuwRmpjw4T2I42bGg5rEfwnec3pb
35/6STuhkzXvFdkjPTYQs2ZEQ+8FV06vu4uvoFpIW71vHz1bKIbHg0u96SSP5uBz
ash+k1fcolk5lfLK/wlW8rIjidf6vVCbGAne6jKoSsXcrYBTCshy0VR2dohlZUzi
JWYg+ZTQaagkmX+B/8N+AuLsz40tXmsc5iOunS7i/pSkuQqrpH8Ztu//tiLGoWic
l7jNZINxxUX0H6Vb2RplgJ1LTTUOTGe44AIX6hcdzOhf7m5dF7m8S0rEw5hRLt7f
UbGVwgfflWBuVSv52FBh0N7vHA0CbCV7IcKVwHech12NDORLDTcZ4BAvpU/BjLFE
rcI7MznOT9ceLiA99Y9GvBoTlB7gG82iM3lN66Th2ymWl5I+aes3L2q18a9WFZ6j
/YRUeKGdhHKxu7gTaVFI9JGTcRx2+vAA+5lVTM39pk/dx8ZpvCgq8sAPn1iky/H5
n8iijXXugxy5RedccTJKtFTutilyjL61rVMYqRxJN1pMDsH8oLX2n6elKy5jDSSW
Lzjzrx2JHnz/NteVdeLNoWGWaGGncUjqeY67EZPqtxi7fezewvkIPaHuZA/bSdYg
2MxbCIqhFQF4XFd+5OgrZx/SVPQX8Pd0knowT5JyzZP+Qpd6Er9huzX09V4xVKUk
+V+BbHFsv1k5SrG9l5qvppIn0pDQlyneXJKNqL6SXJuB4xOZNI58VuWQI8kcTBb3
aoU2K+Y/D5CiKpcw1E1PB0cZdf+hsg6bpGJRmrWWLp7r4ilo2eB+j7WUby0Pcrqn
wnMQTYpVnO40FNGY0IGPpuEWCNLtAfQOucij1OCQxMyC/Nq3SBYT6ePM3i1pshHR
11lI1SEisSTkbegpXGvK1fKu7PmwBhIEZz4181yhsafNVMpUHOY+npj9dYBck9yD
VQk//D25qPVU3sRCk9NdTSQAVOWHxsTrohBVQ8zMQ/w/So16eDgTdspIk5+I9C8s
ACs0txV3o9G8pyBWgpYS4dpS7rPwadKrNCYPwELdNR2fojtI+7lOvGBuRh5OZabd
sy5mIAE2GMEIrezp1mWRZB3UGMTqu+wUbfmg4vNtlwQOhaYUHVWymrgP6ys1M0E4
Z7FNHJsESsZ8ubMnG3hB2NJMpQg7Rxo4yuqIhLkTTDFarTSiJ24M/B7UxVyY7EDt
pAQ752R4fFEzGCvm8gwX2YYcQiy/sbE25uXJR0ESCk488hv9VMs/vYDrpx0OlYFL
nliVnFLmEh1+SKXuzNCQc0nctFjwJyus5cCFo2VQ2S9dLRFA3FLb5/TcY/ZLDa9e
MVGhqH2gwcSpr7TPFen2DPsxPgmPkNWwZmCN0Svn3NTarzDROBUpNwseQ1WribUF
SRM2IWCtWy3IUDskgrirW+ev5Ae/OXlI82GQ+a3xEiYLTx4r6UKmVqVDt3eG9aRu
YjkmzhJq3/whLhOvU+vPMa9C/Tkpg2uoMdg9Tvz9Gm0ZWSzQVy+UnqstgxeXVXK4
ZVWlche+u6j+IQjsNEyvkQaBFss9+YlWlSZZ67B0HjN8hcySKTCHImOwLTeu9Cew
OaYZTeB7pzc7gLc6V3iv63wDEr2xLK2/zKbVwaPCa8LOnn4rzRtzNpp56Jhcsdt7
1nARCBqN28MDJsgowa7k+3DGsMiuSx1IJ2CywcOU6LuasaI/2om1H7beb4i8XW5C
g8iJxC39L/0bjN7wZ+Kxw0giPKXDnOCZAKA2b93UQO9ecoO1QoHFHwXKe6tzO3mC
+LmYJE2SiNUZ0XKYWm6W6ShswhweFVWJHI9iaKXrv30V4sWojYfZjXCywy99MTzq
01IO5g3dNg06VTKmVG+PtX9h2u+9iA3hzQexJfzCyvx4fGZbUCx8RxI9QvmWLM5T
WAXCtvHGswLOeoeQZCLlLNERvhe/9UdjgPnWu/brj5G2opvfJd08YNF157c0RgYo
0ES0D/gbKTYWsv5glLT7ozSrGPLGnzXfcXXHlBxFmwG6dOVxaajMRudX5qlXy4a1
fFv0XzLNgqjmlbr7ZQMFueiLfG9CiPVWT0EKSx31B0dJoXdu+CPxmFESFt85MTM8
DlgthjKneFJ2dhcCoqX6pUaPUxn+nKdYC5lL8pR7ykpEWREmn8z61lEKVtRyT69e
/oKUuFNsyYHYnMv2POvUKWKGVySU/oPD9hAscRoyL4qjPVBIwvAWyE+MoT1lZppj
QeMf8YjGhCpeBqKz4k9QqytZO1y35vjKgMH1w25BZP84wfeXjkV9ois4D75pTnfT
qRwq/yD/sjAqfHI2hC4kf/FTuV9gjfsOB9jFuoGJylvCrsboJpwajodEhS9+fqRP
z5xYGwAAzNai9SRJ1LA2QlJOpI7Ltdm6QqadgTJLv0v88DqPBmAkoDIbF02pLuyJ
qQcMWSbQhb3uL6GuIozruaXC12AmvWOwX4wX9CC1M3Ij1vUkT1IjvPBB2k74NgrA
MN8vsAONAZ6x8gSUGsL3gpgTBpDMX3S48Yn+PFEFRnFrKzW8J9/lVxLVW8FlaSSD
W0a4uU9mN3fHEXedpP3/6X0tFnA/UtaZhOjeppPdjMtAWOfNqVQY0glvxegHLmHS
FaEnhX9IJYH7PJsqItO1TqHJTlQUMg3Pgw1fdThP8Nlod+pr0yZ4e8gNtI0LdZm2
cg/TDNaZHVnXQ4Ekze5yEy+++L9vr1kjN9ZlcrG2WChcMBfoqYHzJiIQIxccoQkN
i7JfDqbGCMarEioLAKnANyEfMXKGKVfKAEZL5bS4A5cGTOyYtl+9WNCc+25UJMtd
MXfY74ZF1KQOVaXKEanz+DOTst2TA7Fm0lex5lby7XK0+VlyEjKjPd/WAhyzf4OX
GKDXqaw2//DlWHQqYenjVv4M1QzchP6s6juhqWOi2ocC8YMo36LULmbGZS7s1YWL
VQ10CyFnZxD1OpU4oW2r46pR8o/Zuzj15UlG8j5sRF/J6tvDPHqyVWlNfBeU2vPN
0+u8edclgfZx4fxoDVqDxGoaM6NrdODM/62d3nBKYw01V5Ersekfwg0wI+cUrQtl
3nKkaurkfMEE98hRWLTG5KiMXTV9YWfYtclAbgQmn0kCmYl0gOPBr1NLW2N4UG+I
nDZc7mD7xqOnNmB/Tws4B1RfY8VUEpbR1O1iHm+J9t6cc1qBWyer1yF/gkDTB/GQ
Q69/ZKbpRwPGEnpwj6GMtBEgjweAaNQ9V8DGHkDE3mpIalvBP2AsfDXI6s03edCp
81WaQr4geES8pefNKHIZZx3Ttk5w7zyoSA9DeWNvB1Muq02oFpQWMc8L3uyVuNhv
jcWztKuzVrdJ6FP/Tf30ODpuFbag7uJfpkgjSHXoEptZi7+DesBD/8KtEMRmoO/j
pIJEGSEYiHB7+MhK5z0w4rHXArWnxl/XIU17u13DvjKB6UCzixizwTp3oalWaLX2
ghlzWVkW7e3Rl4bVCtB2oDPtQHyk2COaMkwu8GFtnUr4YokobHo2oGfYrwG4Qyt7
/KX7Re2nieWg5XRPAsFci1VqmoBkftUUS8kRS2nbYvxyzCOYH3e9OmuCOxUbrtaK
JoFiwOpdLjI/z/291NKyhzdl/xyWX8fn8xbxJ8I8JVhoJPDzKPdWuPA3L6qBezw8
lDNnMcZnyCczqMJCs43/Kvn57PYO9KMgTRpALGFKAyefpzeGqeImO2RUJsvVN2IC
FYWJ5RnjO1emJCPYFZ09VYhokJwI3AcDo+0BNg1kXOWzQknhky+AhmROQ7CaB2zB
GjLgpSCF5K1O40B/+SKmvWyc1HEFEDWB17q3CHD2B/i6c+N2VadgCa7QsfFdGowB
3C/+v6+9k6rwrOxGUCHpU9CpmvyIF92DrDDfoGrqe7bnGxdJq7v90HfVd4Q/+f8Y
DcYtl0yKtwI99/XCVyIbdr5cKCxTiyj/XLStb/zmWlE4DXOFR8Oo++GKtKUc4eN4
ZW/dpFLzzFPmPiWGfE4rUDwFgJEoM6tfwHGs6eA8VG69rDsgnGcr5XKxxw/3ZnKE
/PMTujXWRjq4NXh/Xkr1zX4LXbgSSRQZ6tubD5Gr7PiUZKYWtDQRxwxtxK2oh+/C
x2H2Gj8/jyHVX2BMMYNo6P5LJiDQb3bH/xtWSM+8xA0QSowCIKVdERtN3gfivs0Y
wqXD/Jdhh0cYT088Ajiyh1qSBUD2aLm03xTjS3N5MkY29Pv+cOTm82vfntCWFy8o
A8d3zYP9bRnN0/g0gcssOCQ24j+mmzPAwRSB9Q7+/FdLBtWTBtE/jySgU81iR/wG
GowyGfPNtYHslWIa/p/BxUIfbKMNHzU45mmnmjIAewO3wdCD947gQz/h0ko4zOEb
ovOjDHbpfB4MYtgiVFTJF7WZurw+L7uL3YHtX0v2J576O/KU34Q/lRJCrXnzwPOn
0hcLC6hXYOdUjmx29SNklnoM/jWK0wfkSVgJp/XUOZu/yuZ36+J2tUxVau+0j9S4
ZAP8H5AQ2u1BNS+wEKt5tHwh5UzsfAHX273Eh2NsLlnUw5+nBR3VRgu+r9wesYvX
N5wga174eQ7aDfIl9TCD0mNxcy8znP30GUEgPzIdG3j3YxvBWcFx2QG3FsPTcz3C
dTYGYM0B+8luKO7/3cZWFa+QXukrn8hrpam35MtxGJd4cRN6Gfs6QTh20xLloybj
77PneVuk3j48WDVdpzBmyvRl1C0joMCZhWbV2+gPDJOat0SIiS/CzbflCk1TPvw0
p5viez9s2IIQuplpAkQvjv14e4/fSE20P3frKvZJqfFMBcup0tJq0Fe4AYJF5SkF
oKsm9K4G08fUwMyEEZNIiMRnEd+rSWlMKXeMh6J8VG5F3zLtlydZQElzA6JXoozd
mSdD0RJ126oWRyEfhbINyDG3d0k4PsARCJsQY378CMtadgLQUUb0D9ObYo19swre
1DA7U+8+BvwTeblIvVmQaTo6geUwQvc6TAPTpsO5WxUfg4Zw7j9zUpQdivQEowl3
ZlNMVARbkYA9N+FPDpZJj/kxQ9fzVIw+elVAO2pwfxg4WYM6RIZibgMCPhSgdRTp
VwbjMQs64tAcE5WB2bVYdjxfw3VYHnhthR/82saQr74UfMM95vexxI2E+wT2yO15
UYGPU593mHIJN1dsy//ohWDSlXC1sqFPGIvlp292H4KHJphqhHQ5XFm/xZVYcNni
b7qtUR7ho0AY+6IA+RheXAHm+LaTEN3NpaDOTAMMPcMmyOs9aReVMOvzzGj/y+V9
IO092qyfbW61eip+aNgrR4PNhHd7D7sLXKEDBuMkPj/q+UWS8MRVUuWbOwhkM5tN
v7nwLNGV3dqN9+5DPSmYQfJlg8TPjIg+ET0BM6qyAY2xc8ncvhyeVaE2HIKsE0Oe
AINvdeMlgrHC92fkddW2ACS48oAvfAm6Zg3DwTrDJTHJm+8gtCrA+OlFZZChmdlQ
NwYE5RzzLbYaV4t+T3mWB58uH/N/rXJHgGFQ0ZeEcHVSUVaivMD+99nYBg0rEd5+
D1CHW3dGGOlyGLx6WwmzvS1PHuPGXlvwvEK88Fch1Y7O4A8HBts0VzvKm7N3NVGQ
IBMxmS0zD6wEBX0408vowuf1oPQaP0leyt6h3H4lUzxMxvxLXCRFRyGMIC3eYe1f
ySe+3LA7ksWLJyHZqzffmoPfddNpPxduKVjGtXU32KGpn5iOVIyHK1CbdVL0Llwk
PZetKDQX28VQBoiM7How1cS24ZfSmqxaeM4ucU6OtM/hwh/EYtSgZofbcsAHCvc1
4BFSZrkUPShqk0vN8nEWWcZ4/7r14lGp+/6+4w9rXKhsy8/2oWX2Sp8B0nR1eukT
S1WjF15c6vjZzslI0mt9ogMcJovkvBukZBkpl5zbHCkV7473c2qVf1gIdkhnqoxU
Ez67nNMo2xX7II3w9s2K+NTXpqUQEVwRkF8xGashrNRIGXCl+hiF3UKfjyan4rr0
5LxjONPW2Oniz5fehOu7nL33GRMItVMONqEZsrSDYd4Bu3ubG/WkIQS+nF96+0Ds
hinKDEFMsabr2kKpPbuY7PYGVjkdSnISCOuYZ4LIh3tIpyqpM5IND9za6hIKCSNO
DC2ctgb0N1aQ7bUWMldHKrsbjIazUGhjVZtWGmGtWkbQLWBya9rG0XPhjdAIaMpU
OQnjmA9Z8ii1s5HCBenHhc6JqPnNnxuWnO3XZuKHHeCblm4y0SEfWNJBJms443To
j3dX/PMKaPygTGgDkK9GLy93K0DYlBjIUmg263Fxu6KHMSP9z73B/Wy0lc5siyR2
I194FjNxY/7vDgwmm2bfu1IpN0rzY/WmJs/a9PXpKYYLarQmbL3LAF0UHeS0RK00
A4pOmQ1ddcsQ7krqczINgoLZxUBEzVuvi5b4QgohMa4m9v2lrDUjUHI8pM5kJzO3
8GYwotwB5nksTAnS8GK0oR6GSTd134I1Wd2sBjAnE0ES31acLLZgIg7iqewK57Le
mYskXavEDfM+tn7KhNapbZvpwwgR8aGu5GiaFpU8dLt86d/gciiLJ9Lu/njCvSd1
XIt2gApr93TUmxKNtIGsPtFLMVmS9SxN42W3PIbHF2ak1nCLmBVr6nQvn0NA8HaT
JzU00f90aRZjN3cokUX6wH9bGynn5M2dBXuJxdzPakSMabze9FPMWmsrLCKKa158
v9jhDP66nwqSRLmQkaouOx0ChsiMvkZNaO5qcNSm1SqDx5PomOC6R0mQ1xZgo4f5
IJ33jvLEEcAQtTSGrZbhvC23EdF8W4oqT2rxbO+1saFT7Oj//IB5uZ01Johpv48s
/t+QtyXjVnldFEgxFta2KYqJZPuuR0MvoEcYlPBCX1EdKo6eyruUjbAqqiJ55el2
2NCAdKR+mbdGsQFen4dFwn0liYV/NQjHYRP8GJQLc9Q8WaXw2DSRbAsArBTc57oQ
rloMc/OtM8J3g+qX52bUtpQrtKIlg3pz8DjdlWhTQh5LAKCgLe0klnLfz5twBM2j
POx0rsE2YPOvSdLcZbDc2MNduoWayTdQKig721f1JjlDz5wWfraLybVw4KJgTvB4
IVPhndttZzwODgeU08Lf0GWxUgyZtvqTxmo2jOkjNccQIp42p66Pq1JNY9Sk9S3V
WXR3rxhGA9dJh2L960vF9csVIn1a8V8A1PV2Qwb3/Hzn76likE+X37xrXvJFLwFP
r4o5oAG1xT426kweeTRaVmqcsU8KIunGJUFruWZP1b4rN+pqSlvvzH0rEqbTcECI
srySTL1ztnQA7OmZ2cvCDkItJ0SKK2/qNvHWwrtrda+xGQYlJ1iJhfj0MSg2WhiW
7M/kWh8Zha0IoI6+7c6lB6Iyh3kOfcb0uA7Y2OnVBeG8IL0Jk973y/ni9cjSYdC1
tUH7uSyjiMZ/syOVeLQ3qUI4/hlxCai1GLIz0VB1nep7aZBQlXPeoMWD8pL0wTZw
MXmEwTsYkMTuag/BDDgHYG7kCEmxYYYvIylameo5Mo1k+vaZuDEliGnFroUsZ8Lx
dR6tbgyqcxBByJtsnRxbQoZpC+ff11jTFlhHpQSDy19jIxCKnwX+CJ96kUlrVTe3
cWYyVv+QPuF4EfHpcZLnZXSJ0nPv6kQEjD3ujQ8hxfBGkBBnzP6W3zMfeLEPjkQL
ZVhnUbbmUWvyfItbiMoj0PnBQItyH1XBoS2z4ZHejuV2wqo4YzxSKqrJ3IkynESm
ghDVoAzd43U8cAN/WxIgJsAuwv37isLMe/Z85AZ2hXnx0LQAIGLYD4shd9zuXVN8
xNsNDslIRaAiMzaP/MhIog4/Fp0Kh32SUhb6SNESdLx8j43D3W9m4Gcs347DYNgA
hsBAgryvsJ1Eiv0UyKCMnvaYljNrKQb3OV39UncAWCDfcn9ZBILKxMDhRbHk/q7I
GPo6SFaa+wFy8wt82aBBvEUrHtcaTvaENhUaua7JgbaTQckYE1xS8iKUZn09LrEE
XdR31DMLogDffcaWJZEPZSyAlZuN66rUGZl5JxptJSC1+FtJkCk2o1zPBysoq2dr
v5f9KzBGckTN2LsInrtB38srfdtm5xk4Kav2mWDi1MCypUg37B29MKX7cUXd6fJ3
O8qFmDrZN4k+2SV18LAtoBD6gw2lkq79DxaHPBxA4ZAqC4d8kQPds5r2JhZMyQ4H
vy/4y5rqcux+9luXasAQwLYb8DOf8jFNTE2Cn0s6k6FjXfWc/yVkuu//QKuAAeMu
aubGg7lzsyH8DtpTSCv1/ut5FjPu/F0PgWRzYD8V72LSELfRJhNujl4A+M0y++fK
1dfqPENYUGV55tBANziQzj9G0sn/vYg+ziWRRpGnvmsDpdU5GKqs2SzNXAwteGve
HIMAcGZBtkVOANhQNgFuFFiTuZgVcST5LupF7leMuzLdbgxN7qFfe/mdlxlFdI6u
AdzSk0Z20O9Qca4rrq8RiJOkzc3jwsJ2buu26r2rfrfpZF7XlB5s5OV6rj8f1Pbi
7jYxBLGN1++YXDJNQvEXM1XzKDYJ6xB+t9KYscmKRWfFJn/UbSPOKWqNJg8uZd2d
woHxagEJLd8yrzUIDaiE81PCUVrp8TI21580Z/dJdAu5pUPXXyf/xFntfMW8vT77
+FnjYxA8D04VVDJkI9oypbbEHttzbntJW6GtkTH5XWUYhOrL0lxLyk2BZcYue7eh
Ql1UE6DcoRtbZuxPsCzSm6P2q014CnhIGYm0lqeE8PXMqko4kZCs902YNsLsmDBL
fgS5aWg5XZNZIWgdV8tVQGnYrx5rt+noTOJv5uMKL52Ey1fFlmQdDg6rTZNHngZH
etXw6FOgEYIcrarb/iZ48sKWdVUgZE7PoIR/LJBerZoOgCrW3Ww0GEXiPU09nsBh
YpPNqSAtVFYKaI1MksgEDr0jgZVvhlK1ofTPTh3jY82RVKvE/xV5gsoAO+Cd/wtU
97UcpLicKZsC5m6aQzOQDfE36kCKeMxGBiMkirlZ3nkPVhzY2SysqtdzWzINnlpu
wGZb+YwPZWMD0uA3sqsHKT9XPSy8XmR4pTyRgy5xHFQhAwrK5BgmPLOTUrYfz/hy
cefVUzuadWbIXUs2GHKh15d276kvn6fs+Iu3WEqQRwbqF8Xm8oUoSEyc9hkgoMxS
FVtlaiysm0nsfj3IOZNjl6mx3DAwo0OTCAZ4TS0Uc5IMkOigFWq4BsT6PmQr2dw9
vZRZf5jMJy9vu39PtHJ3caryyHQTyXpn9iOTKdJr9qOOwJsHci4rds8+BBAYU6+Q
47Bsic3i4auBEdK4YVYXVz+epz/VDMQ4oBlwQoyHy8B4GbbdrdUqIP56Yzv25kRc
l5ylpEAoDVSzZdRTPick2wLoEOEbscXn5FdPR0mdUO/3QzZpoE6odRddONyjQSiE
kge/IQTbAAzW8jBPNfyvjjl0gfckS/X4M3WrpZiX08RbxSYL4O5bwUYAXPbdtbQD
cZQGZjVia4zQK8lgmbNtMUAKPHe4kyMW1DJNtW9tPE/O/2LO3ItZc3CegYoqADpW
fPpaQSHsU7uviunT8yz0o8i7nYbKsrdlMiPhjUktpk745AMNi6TPwtNrWUmrUNZS
7Ef2p9ImPQZ1AwrKBt1qu5SML1P+AMHxjV2/AtJcJ/lTiQx8TxhYgYatQiW7tEci
5BCteUPBp4h85+j/8wiRkZflrkFDkWBsL42gINhJnwJG9gHfbvdf0xhkiO/0Nthe
+J3yRH750LmSePps6Zx/fGnYUVgc/WHcT3Uo275Z726E1qz0YAQ4OzpjTCdL0Y2b
Bw6BQcZvZkbyE0uwLk1MYRQHlx0cRPgIW3iF0HYAcnOu5aMKDT17eTPKwlonkk6L
NGpneXdrSpOzd+ivBl8cHE1RpkZikxKOz4MaYPDjnB7NOQpZHAN84It6SiRQAnkY
9nbUQQNjDtCEGqejhwS9EKIeUwQETVZ1WYVJlANU+pU93SZ+THKqNCwytn5XR91h
eM11NykUYdN9HLBYPCNyybAUveKHo/oo15DVG9RaQOTkk6C7vOwhdzZrbRhUefhZ
+Copx+bm5GdRIwZ+IlY/RJmO2UB0NJjMYnfOoqsoxdHK/KsuWLTMlLwWWG1G5LPr
zlQKbBMoPpSfFguNEXpOlyNm2QC9rAWTC49p8VlgJVf5kOlhicIPLL7WM75OY5KB
U7HJliVm9KUL8oMeXMOQGCSJ8F1ldJaEr8JdjsAL94EWaKvn4erJepRltRPWWwpQ
phQ4aIJDrvNt1vOO2AY+AC+HQAJidfu7iboNylmrFJk5O/5zgAuy4l/AYIjUjj9n
/UrkNNdHQwevQVj7f6o6fU4FaMRcwZmKJix7koNo2fsXs3UwH+1y+I88EnGZYWrv
p19YGtIot3UWFpq4eIhntRE/AnSDZONDeFqFb3B72RqEEJJ1NewWI3RlcI1rXmUB
LloXB5Egwh7P2C502ckRiwo2b17ThNPxS8uuM4PRut3gg1noo1nEKcNrQElBhznv
qeIIYXs0vA4Vr/9V4LLYFiQAWDnXag7KcrLOM5HJDO7O/tl6MZy+1uLYuS4BOFzY
b+t4oRyixvmIzw/O9nCdGGIkbGwbMoYtLFySg5mrAv2ujbpbCYWuKEsVuDk7wHpv
qABO7gQ+eXrFxzzWp0tDKosRm+FsPl3p249FVke0O+yJOaSufL5R53OulpptzBrG
MQluJd2X01UfJV6xJWtgdzh/gzNcnNaiw3e7MjBiU0BLYe+gD+9ohOO7A9uMU6bH
HVxG3zZvQq+4nuJuu2AN9sRrPtNvbTq/sAcOdGCuworrbZi6ouX9XZ0qxet02cn/
5sJkpMXxE2IPoY7pSiqAOdzFQuIX5ug+cT0gzWO4KLXpgm1X8jKpiHKsGbnHmuUw
kKpEP0JjCbfBCan+Q3eJhrUzE4fzuHHyUpiaJYBHPC3d6jvrTTgKv+1bAV77qP4b
dooIGjjp/mCWPtRJ8bts9RuntRvaf5QCJAA0+bBbvvlhFC+eUfR1HTQdHfofZ5uA
E3OuDT/1wURHnYznoAUfy74kfYSvdV4SJyHw1DoPDLHqcY+/XlF/5vZax7wYMg50
Eixu0miSsnffxbQf9b0XUW4PG+FP8k9jw+YXu1Y+ei5sJjo/vd0/v6it/loR9u8t
1gBVZzDEwo472SOVb/8Mtf+TLQYjvfAhHIBJBapAoQtTUUqxuNHX0fd5vyQxR/Ku
eCLyqtjJrug6ZyaWqgAl1VThbDyRiFYHp+DjfiCmv15Iij2XNu9PSeeYlSo2VfQm
HTUBqaIErOfwwK/0PPKZ5sonzmxt6B838YmvIxSy3TaIDD2eUxra8QRHh3WYCixs
u7x71JKJquASHYeLikxNK4+o2jArRge8vqiwOYsAzTjawMCgG1RKUYZbW5OmktPS
C3XE1vAsRvmbzH9P5qMHpwDk8QRF91rGb4MTdkU3z3TrwQDUuVWCVN4fJy4afsHk
1DFxoYnRCG9eeBOf7R073XZc0YhxXpF2eGX1iXXcIhJQ7d2zQHctnR9Ai7/Ig1Op
6OacPG968kUW+f9G0qmyMZLL0YihrHtNzseG87EmO6k2Vcgyr9PBCWuMeWmHTsq2
T0xH0mKeJaFPBD58g/J/2yYGyLxtIRhpEMNPH62uGtcugiIbA+hcGVug2T2+bk6L
Ba0HmUhxUEBgYPb+n5JdUx/o3u4EZ+bibR0agyGkEVXhcHrNF//u+8OPI/8ZObcT
Q55CEpKtzl/+oRQ3kZ5f2UXhwlFkTRgb2j96SucQztQILfkYDcS+7HKeRMjsi/JC
afCMj+ULC+PYprI6uX7F3MUZd/P9ZPwZu3ZDpff8inWX2G1/xm0MvI2a5v1duz2a
m/Ty7Oh8I74iLnkT5tOThY9Bi1G8cRiZPaN9MP4+6WGra5yEYEhErMmHvMobYTIW
XPIIqF5P4OIGq8dgI3RITqbpUHrzzxSbmQmTeZgu9ta/IrtaoXYTt8A+TCqbJLaF
h1vf3/eGsZ94VdhvSnffTt86SEKiveDhG3jkn8vFmQzJ+T1YTZMn2QvF664m7S2G
kFFpL4/LklKG0HBj7UipC15UevmXRPJopqDJyZdajpHfQxzc5nbAt/Npun3YeErf
1ry87IZk2oRcthBwX8h2P+TFfVykhhVwn/6vjQKDXAUQJynvow8LQe+edEKJ7uTk
f+VQpAqwn2fX2gvKAtaeBF/6LclYzPgqVprez8Yd1/+Bdtkiea7JB3T/EVtNxWDc
QPEwKdJT4901a21DgPlCldw28rALvwiEAHcODvhrThAW2aHd2zq9E1d0sRdCChps
1JylAyp3sI1tPHTdLB9cf++1H4HnugsxFSJ8eEBRlHOF0OKIzKeMsJCxA9sP8Ca+
5TqgFto6uppZlz0E4qszkhgj30lgEfwE+bO4Q31/uhBmv7Upn21Fej4tZ3xKHN0r
iDJGT7Bme53JjumoIQZxkeiaHVXBF+PX7e/WP9hXeHcezhiwt9hcpE4VhEcqzvrY
hK9mKISrF45qYsz8ARuEbENvv03ch2oKuJVunx1xKQ30/IsErZuzQlWzBz47NfZU
sa9OXBjhqsOpz6B7q37tjry8AFISO0yrb1QbjuAYJYlb5MaTcAt3+3J/bwawcr48
xJd5NT79g5bsWZMWpVElOSCxtyFf2jPFz5DbN5OpXDw1M4aPoYGxLB0+epyLUuJ6
suzSxVWKptRHe/GesIzq6HMIiNSWRJea3ithT72wL3/TjGwUrIsQAqk4qpYLT7Ea
X6wX60wLGsc1w43G6WBigIyKmOJ5nQZqurTLGeugiw3VaBHuWKlKqTxhmn517DTb
F+ZZXokWfUf0QUFlErRU3TjwBZAj2wsT8N/SlkGUVrD+zP0OovTf6StQjlC/bjMl
p+Er7oJR/APMj8xNA3nuVY8UrmoO9tokD1k4snWZ6vlMHatDOiXaaNL2FHG0pVkx
6+gXFmwmnmZopsJ189j51P6eNm19kXrPNsNw8YIOHglepFexZ+nqzBakPIXTMgvL
OpbvtgJ6kfdftWmRTEpGC1QcAmIgGn581DiyFk3dja2yppAsnAm+MWCYFlv/dE6P
pm6wppSw94C+XAHqiJsyJphTzJE+9lq7CCpuvIpSCW0h8/qWqLKwQ5n9FkxE1be+
6vZoCikOwmIWnmHmpr1WXeAxrZIawyohp5LzlmH4QX9ne0nwC1kh0g1Y+a6eNo8N
LlKoynIzG27HKEdaZP0tzt3jzEurZY6egPOllIE4wwVHyUo1T6GESEqGbx0/AX/M
btA9Gw7KrqZX6ZTo9PWK1KwFBsx3YDSwThBQbbRRqaKJLpqwxujIHGqtBz0qT5Eu
crD2p0/tEtSsQAdN0ChbYrzEEwJR1IRSi9MYxbAd6En9F2PFAmy8NmAlz1gYILMc
RZR2idXN7yataKJOWYZy/tZZQ5CVYAOy3iBpS9Uy1QhldT/WnxUp43djqjqVhoOs
HhnWB7Wy/p95nOKZa0xcVqkldzSNziofiq1/kepHqlbl86xal8bShs30eTgvJn1n
qO9cMfAT0Ma/+Z1lRi9pcPO4QxiOJcbGufFp2T7p+MHRFtddWkMxTuwFvVLLm0mP
REmcbwAYdv/AdZehXBPbGtILx4zVwT0Qv/FlMu67EQy/niOolHLGwFISKrzELse1
ORE78Q56ql+mjxDkAyfanC7D7wuMJT/u3Lw8CILd0LyRoOmbrjNcpZE55RjjoqxK
RS3idxeRO8vx2L4EKZADkJsAnvl5Uh5ub5vYDJGOWN6rOVCqKRrvhzXHS4a+QZij
z0YrEGSINRIjPuGm5YPy4ss8R484dK5Pj24Efu+pcJxsT9QozcyxE2W4lPezmRkB
UTXwqojUn1+EJK78617YICIIwXEbV4A0Sa8qzaZNtiByWRsokIego3Jt0PXhKnYt
E5xMRztUXRmz2NyYG9Q6kRqJ8w7steioD4NOf7FOybFu9hGbwgS3dlUsv+ErZ1EF
5N62y9PG3Af/ehWgeNbfy6QIlBZaA5eHHKwwIiXPYuWhm+i8fMyo/wJYfeqFN60u
tLNmwL8Qf/Jyqg1wGNqUtm7lOPLWjaH0BqoTvQlvqakduvGInWzcl/dnlRd4tMFP
bxyzF8++w9eXcEKgg0LUQKllOozac/wSrmonf6OFglRv0eD4kQipgAHieY8TZ+45
wjwqCf3VUsAt3XKVXRU/F9Y0hy65KC6KlAESduYo7531fN3t4SvI83N+GTkb2fF3
eJbzCP8i1ULAI9DpqfgQDetYbVep/Eiox0Sp8zIVDct8tv1BBwsL11H6S81Z5360
3k5mn3jHYbdjweH1pyATA5PFNgyVyXroutIgUYDj3CVWhUvnGLcrHyVx9M2AVV1y
L2AK5zMMN2CqqP4WaayOrlHQQZ6rm0UWVW4oHAWsoIQBuwRLJHBYTDVubFZwUpCj
cQPICKScHZYJqDSbIerFzSXq47RT023CackB+wII46hXB45R7rKdmqlE6yW1E/9d
BDVyrE+H/I0R1gmMfoatQoByvQUkb7U7n5YKH5DmW22C+a81qICndPKDlNSEE4m7
jCy0QMmRlhRWRbsAnl5ZK1kmObv3xWmWDfGyt5dpWhebwgHmH2BAFF/pivfMgQoa
rOUtqUGs8us3zLf/Ajg6zbfKyq6KMxthD9LU0oPEQW0mNat/qA32I/3KyZd2BmBz
u6zadBpIvf37PrZ6IvWr+hiXMMM7gUdvmOKjrftaykKOw3iTnnwVpvGzAZYI9NB8
kD8y8pX9c6GPTIJ8wwih4b7VsZSwkfOuOkUzuDBYUZWncqBHpKH3vfcoHJDTkJCg
kpvQC5RSRUWrVIF6sG9xz9wOEcIBmtzg8Bfmd9c241ZJOZmpz0IWCpUyW3D4pikT
yfvZL/QTv+3y5l9Ix0SA+LVmVoVMG5OGGlJV8BduZzhi4DFw2wlzsG7MqkZ+jXeY
V2ZkZUB/oIiK7b8i5RK7BQnQvquSHKeqCKEnQSFKGt+PoKnak481n6n6I4/djU+n
CfJArWZpshx7EFyDNfwGxMmU8TJdaEnURGWYa4yMFhkRGOiHmrmfmW5+bHA+egut
bXbaFpmUHUu9DcKEzAgz/fHRDwc6tpLb6c9QT6gdS1+T/7zOvcZt0UsV9M+WGH6k
9CG7na/bvV/lO1JvOE1EQ0vM2QIHOaz3pr/BHs7NVE6szHrZ9QsE6NzpBMDvFeqR
aSGN2URcPuMUgP4pYHYN7mwiOYkyk2IBN8GhERRiCaGp70fhNcCsuOMolcZkSsBW
wNqw1FrKE9PYxmY2OYfDwQgULXJpGlt9wrCzZ9JpG8Iot4+S8NROXfpdHuAiijDc
+1Ek8OwWNOvqWsytZIwgXh4ApuFoj/Cg6fSakm5tpdRZS+vXY7V03vyc5pm8Eqn8
y2Na9NcHlkcgwXiygR5RqCJZZftAeEYXC9q9lKjdTMcaZRRS2HFyr9HyXNv8qZjl
T2gD06pVSJVkMu9t+1o3TJrU+rcT4cBvL/JI6XCWqhkBI9x2IyaO1NuE3Y14KMPJ
Dt/LNB5SrMCnsh6qkFpy4qzRlRDsE9+Sv4FBMTpN1ZsHQaaMEzXoWHkOLyeHI1RX
MIBEu47VeWSZ8Ws/gspDnoGJtplbIrJpmxNfTykF7lGl37wvmSyYhDF+u0E1sDor
qZdwE2DZzDqtkkxb2go3anRMlUwpAvxrEzseSvFRIX/ads5BwEQpHUwD4xhdZX/+
I13DXSZ79oUdLKdCzzGDvI1qnJE+64bl0aGV5GgG98jmDs5ls8XjHFNVZJmQHddg
gWQd8H3YyHZasICabynoMBRxxn/i3breu13UBFg+wDQKm2tqIwrT8UWn6h4Stpfc
0/DEVwNR2UQSugDSe8BvNrq3k6r+3FUc/6Z7+vm5DSpxM7ik5z1WRwyGAHhEOyKH
axNnMl1nQQ47HnJ2buTddDB3xYHOl3/4Gi8ti3MBigh7IvZIlJ8a+i7MX9GQ+He1
O95EUUlrJhzxZgLm/PVrCPVuREoOoIIzRYPN93cQkI2OsH6/0sjI5MXkIDJos0xF
XB4zTIKO20Xv3cUgJFrRfR96m+b6AJruTQC/pKVYT8s4/eFtYXq/LeTWHRROvt6K
Jd+tutOCdj5U6OVtbDfWBaH6KJ4GDxefR2EfeznrKv16+YlyIZivNr3LR58h1i6y
krQ33HDO6cQ8088WH3vpcVvZzFgoiZ3tB2iNEzZDRT+Jo065gWZiANzFT/NDlKd4
/O99FWMqbhnASkuGp6beJrNcfVFH39vSccT8qv9jAHw1DaEWYdX9fiAS8yhgiN/v
FdDHwDOyVva3a0xzqvkWlF8YAdsQjqd2st2K8XEpwUB4KUb6Y+GwZwYQS5gGMqyi
LRs55pCES38Y4ypgJCIuKmW5QRP+ExXQ70Hh1T9EIKzVAcaf8/Cx2MwrFxjI+Dg3
jwBHsGDN2RxTK59JX0PS4Np2Z8XC9qehSrMduUKCe4SfSJXGmRRev3xFNS9S0n5E
yVDWEH4Uv+LSj+C+GMBjkCrKBOf/Wq1CLG7gK14e3LLmsv3DlLwXqLXztq8S5FLU
2/JTPiRp7k3cHePHqgqyMKxOK4PFPWT2rpqcdvlpuW7kTbLR7ZMX7dnF9OSHZDRw
+TTtWQZ1uyFui1d79XB7U7fT4b7FjaSQIlYIEH0Juxs5kF4803u5bhokZ/qiieU2
51pXlw/Zve4PpqzvHoEEoLfJ2oHnmJmp66yQLE/AErOxr6wUTVb8knJ/XkfSfnGv
xAS2oLjMYmZbN0T2GUtOuXUr2OkeIDfJ2DpCw1Y8jNYbq2VFd0zUZrI/vHebo6kw
8U2nRAhzjchqMVXGUEoP5Zde0zMr1VR2XubjpsY2fRH4Hq/oQEv6ZlthQD1P8bpS
b6DiS9k14UzY6DJZu29G6X5U3AKSuc/huaE9VSuLaL5bTjVF93NYgA39NQc6wz4q
hXPJ4r7YYqWC+FOMDPefK/oFLsaQHy5KN2Z/bkMOinnE7e6QHWaaL4QuFpMv4TGq
jdc6w++nLeeHBJCoVAR4+Bd/hgbxQZqK0SHkw27P+h29jNf/3U1Ku/TnURvn1/7s
XSUNWmny823EluGDmIJRPcJsueWFPX20N6G9u/wTKLJ2sEedrv2zvnGodvkaPv43
iQyhG++DPnW5MU/S/Fw21iQmCw7CRyMdLn+M2gl7gapNijpiDBQLWpHbr/kHclOb
Dz3+XCFa3/M8NOnLTU3EkMw/oc+rlLfP15w2f+0XC6+HEyV2agmVDXSx+oChtGgi
AFKIfVuP40YvE3qR8w2uSBZa4a1pVaoSJC5O0afumu1oyzaGxEAJtOP5HEzDKjDI
EC1pKTIsF0n6REgectjK7JirCtnvvWEWoZMVvy+068GQXn5ylrpX86mS3625jdQD
x02Z+hMp4agEkpyB5DjnLKiDq8TTWkiTjY1kTaxk8qzv4aTAZf97h7795mxfE0EJ
EM4Wq4umVcnWebyP9bzyi+zklL6xkLQC3HyVa+mKwNsgDlCPOB+edNRXJpo5VGLv
KvzWlGVYiam/mhB21se2F6rDxXTEbUuaNOYTtgXH33+rEhabuSsDlrE2BCU5rTZg
XRiHxK+drX2tkS0k/H9ijRyEC58dxCSHf4CpyazTcs6U8jYBnyMh+yccf30GvHQO
lpJ6ir2gm0d1ROZ/Z+qs0GpHXgH+4P+qaf5BEC7a1zF+K5G/MAQ7jcO0L56IrXge
HBvMuoCYbOMN/07qvb71JNd3o/TDvrz2o29wrbZksgSFI3oM+30YFv5dIj8322LU
uBqGCZFVuHXTLLdNZK6OOUJfcB4Sh/4u/Fc1G7X40T5zA3yaLhwyk/g1AlUCrJar
NvCllKasYCcqtIhe3gf42BJx10IuGk8Od/YsaR2Nu1aWL4JwygDXkDt6zHsAzcVs
AWuQMCtI6E7O3Agt94w76uAUSpIsZMb8RAJltPD0onudxmUws9ZQ60OyhHhpcr06
z2sKYRGWlvkKYXAUZ8Shoe6iBgtmY0yNSFsiENixpnFrHJl+wcazGgn6ZDPIfclG
IVT6+y6lmrngROqootqPhyiH7xOBsugrO0+ZE9YkMR3OI6GXMcjTd4ih6WZaVVLr
juu+5XaRHhFUQYLO16VAZXI5Tb4EvwY4YNahfFtPlDYKcwYuqIz0a3QGYPLDbseh
HVRbn+hKgCEU45j5JHIY974rN60ErzBAHsoZTW4Sxv6H8DzvXzWzgMb3uqwDsRGY
JNP9+b8tPiLtRh+qx1PNWexCbB84fWYot/J9hgixCD0bWZRQfqGaaErhc0QOQ6R7
81fXVHxU0vI2ftjA2t87k7ATE0ce+9VxE4F0EgOJ9TG9RyIQwWmtt24GaWXb41gp
dV9bqMHHY5rzFPAS9PBs1zOLMubLWSg1WzXfj2U8xgfZn6r+qocqhJWEOVs/2TDJ
pCJB6FbcErj+H+R3WSKti0kADTgpHhOA9Ugf/1ljJqnFY90MMmZVBWd0E9qOZ/wq
F06RdVpdsZeul9wOjuYlHK6tHwDmXueGJ7qTcYWZSWY6kxpSQ6QiCTTWIIEM6BeY
6JcnNAsuL+o2dap138WPJeRDkDWO9J6VyiN+cZG5j98zvtw/8q5hZNo+CH6qOEYT
cgsbUK9Mxu3EioG0wDu89/3HPYxFu80IfcsV4T+fTVoW+ycxRfDVbUO02z4KEqAx
NP1Il1AFhaw/K+xMS6BsGvfaX5cqoCkuqQjHta5ZB7kOch+7M5Bty6E4Ml3zhkdE
rGRpLUenArh8tR2cJJH1J7G6LAeIsLjel7hT7XWZUN6X/mJ0b4XkAnGDTHNLTVYw
RAz3U3tMBYbOVXv15VPTYe1yZkLoz0+I8/hmwWDQZjUpTO4zklGAYApJy2ikqFJ7
+s1d/m+zTTAhPHqWnRRAC3eTInHhN7pztCuCLYsZzrKEvUj/zJzwyU74ZqQAeAXo
Ez3ar3Ah8auL/zqEP+ZqIZGPzlKE4BHUAe1nc3OyIbObv+2cZbIKP8VijvOJsb+x
5XCCN0FtlXj60hknBuSyNVhJTgCGEOjpNI9jXwGvJh+sJTPzpao7+bOTY3Bo3Ma+
FXjep8yDu+HJnANHYVO09pUSLW/PHIdhF3AA/6PVnY+m6sJzM7kl+wINyxPSB5ip
7I8lI4gKcU7ReZdluaIVN6GUxPqV+FblxhcNgzRR/VFH/IYSwUQQJpiuY6ll0wRq
iYfMb/HECLsHePgQztn8FhdzWzYmXr8afHMB0pbCxUtsUe738KxvxaIQpNgit9N8
eY5a1Q6SUhC7a/V/oZDM/7nVesJ/jCK3+QmjT1CxrFRq0to+m+5YG4jE7i+Mekxh
olmDGsbwKcjxGwoDkAQ9WuWZf7orOJ1Gdl9ILwrXaZfyw97LIrbGynyPFxGp1yXq
rIhVgQz3vFJue5MCB9hyeHJkjh2WSU8xiOtB4W3altTW1AVlAeS7c5xVr+7N4yFn
MtfAwQFmCcnKPPiSBBGSGAZqtJ5HrElgNOr3GMCfBTLojfkGDrLr458UVo5wzo3T
ClaP56isiZHbH3TXL5rfnf6y8Cs9Pq4bonJOT2MFRccNNE1HrYqfTyGjCPctC4+d
Z4vXQGFapIDdpQygNXBtetNw+hCvHoCPJt1l1BO5WsRf735Lk9scyR7WiYtJw4+e
b12ws09BSeb6eTDvXwcxEKjzSF+pgiSFCQ0xS0qGDSyUnfTp6kGO0mS3fgk2n4OR
rsPnuu4rksP7pfoiY+9UMugjjHgX2zsJtBoEzyB/bp17vcRaVDAVndX5TyVR/qMv
vVYJDjzs5Hd57yCC1PoWvxovpbf6LlsGkDmQJ5teHVCpUCJX1u11EwQjz3AzseFw
hR9hfCcE6G+o0wNMqePoXvgVaoqApzAPkI0yLz2txpEmxT4yoeCTU+jDR06LX/ga
kaDxlnupZRMkuJiN0owyEe5Wcg/IV0LUnEl5r+zfSMhxy9/vES08EDSnJGgGE7uC
skWI0r40f286+h2MAbjWXPJDkAg3lb8R9XYaDHggnXAqh+53Dz/eTT4PrJ5xUhwn
9a+L8v5ZF3tYsWoQzggdOjeYoYcFFR69H4aGcYhwG9N07IitQUWXiO0KY5YTDiR9
UyWO+OdCnN7FoIK+/K0nTM5rbmIYMHaZVdCqF6LNRsKcY7b0HPri+Mzz0RmC6APv
aPfDQJsW+wM5mWqaI6IAJLLY7s4fkKgFj6ne1uM5jIfqBJuLfYVRbOyS7s7wJutj
w/swMnvWNOW0YpdoXm9coF8G2l7i9OQyQ7fefK1M/IwoKDBdRQPbesmzARgZC0So
BsW919qhiRGnrzB1LICQ9769ppxncs8u99xOyHXXb4WKYs/MYMDU7buaYMaOkiJP
4LpJUvmITJOuBz9nWGI39alM1DmYlgT/3FmOgdEC5SlG3ayXgK6U9vjWS0kxezY4
FLmU+K1ch0nt+D2FiR9lZNtCho0HxptNPVbV/H7Zw1niBQzUz5ZdOZWJzr+vTIJU
86qeO67lyJE2fPb5/GpSBtQU70NbDucCZ57FAswdm7e+hBmhAJa36N47kn+1WiN7
rEKZznC/YD2AmjRI5kLcqFiJccstoy6aVvl9hhHKEpRGH0qXtcZXScPRo2In45ME
L0IiBUJ+AWb1GLZpFky4fZ275kHLSYVKRB4uMVrKYiQ3+xlQEtxU/3a0RJLiIvGU
3uKTOR0eervCiaIoBuEt4A/N9jITFofH3Vm3L7WDG1wcMcZUsZk0u+BSYugFj6hd
O00yy/r8lR53so7YNIQ3n2WUz6C0g4FhlznR3rvllusyIhknKpV7U6gWGjUcqs0n
odm8Mz891HlpbWvlbMbkCDCPq73CwgnqvS1cKHll8+9U5811Ut/mTLJP2anyCCPI
X2wtLpOLkc0T+SodU1dW4XcEtvThFJCu4uqaSZc6hovLzBsJLTxoeqRVtvUOd8A0
HY0qfZXVmYh8kNnMu2NE/C3zxwM/PPcftTjw2qXls84WFRCNy0GAy8UClgS6kxBn
hF8Wih1OxeCCtVZwx8MiVYdMZiF4QS8GsM3ZTXTd3eyrxC2kUHmqEVtKZtC8op6y
zVQ1WR8iTfIXZFXOn0y54WDMzq0GeuAVx/yXXen9aKLiMo/pfPm/3RTIh7eQ1OJ1
8H1oXoj42alC3vi2POFMAkI3PblfeJTSYr1uxPfqxJ1GVG3W7LT2YsAIg1g++9rS
s8X9zU5Jbx3tpocbnvSINpYIBTM2TYbJqQ3PXUOkBCaK4LDY6IcTy3M9MH4rvyoW
0/esYDh3E0pFqV81iUZ3tFEytwb9J6kqrgmm4Mg5HsIaCitHkb9UNnnscYUOuYcK
aJPbo9MfILL2UEvFKwy2gJtRtNmn9o7SvLBJNeuQ55r9kMbvwlYIaBCyqkZ01HdZ
9YfuifP1f4SkkNs74ojV1rgS5Hz4G4TUAsw7hPiICHicMilogKkv8nP5GMyFctqa
gNuyvT0iju9wFoHStxzlO9zB50BVMyB+WGlOGIE2eEc7sj6NZGJaFq9Fob+AG4JC
zztLPZkNBVTVxM0BRl7L38leuaasuCKMXln0a7WuM1bFWtjZF+aQJcQZmwDuIsP1
ImuLNVq+NwHF70hUA7jtxeea9mParl9LDbppFDcCLVgeNw0eS+Phv5C2j5DGpfLm
FB0dPgYbdsS3QV7XmqmDpIi0isqVXIhtFDiQ2vpRtx5oxyweB0oZIMftZS3ueaL5
cJjYjB/RU7Y/WQyXn4BE8LRXrLLLd0EAKaWTcJipCAIEPDi4EWqUxxs8Dx2sfjhI
Xv7KJuKOim0YgweD/W5R29UcKCfiDTqc/3ahVYSvl5bj/KPsFkE6Dlgp/jIrHHi6
qlrfcHiv571JLDTxTrqE1QRtAGyt9Is6kFulSG7iI7E5EqskjYCQYfnAs6HDkrSz
JqYwVjwptD2itN9Cp+O0XrOxWcFcNlTmwHA3qmSa/owmC+b8Cfon6Wd0KK8RxnVJ
P/84JGO8Kor1yrn03eLRZ8e7CUbE1RWp5xeVDJ3TlIC3f4p/+cSE8ddvkEwDp3TK
AnMUVr5oudf/2v4khmDD3aECCe3KakQKXfYrUqfm26wHjrS3HOfdChvVr/Xw/P94
bOAtmh5Boxomvu9zbehiofD8bEkGVXbQ24pDr1k6IXqJMwL/hszxPc9VSMtlFnk5
j/pv2rDCq54fwjHoq7eNgpYEc7cWWKZsXQnIubEncRkKss0RW+BEkW4dKwPOk+w5
IF2D2qWpE8Jqgq8QCBTTBkEU7OVRpTLctVoF+kEX1O+G8ceC2bYVpC6LJR+YXEuI
uIju8itSjojE+/EQgIMi3YLTQR/fuQVXPnwz0LOW5UA2qCq9G53Aj2R2IH4t0gT+
9P3OnLNCHZYFHr3iyGg/9xuMA6fckKnI/fKJN0wdJrpyUPydLh+WUZf6tzImtleM
ATdG9NtEppNGMYq/Gaq0qJqi/SSPk+wGGqsRoGPhkryBJN//Z8qVR2EXxoDngqUx
QhLNCJcd5XcrjDegqIYziEGHIBLqkvjGdxj0+G9SuXPj9R7ET6l8H4uI0uaY6R34
+gOpEfZxqn8Nf7FcriqvCRU4V7ITcx8N/US/pfbFFHMg3a3CLh/EET0Y/x1ktnuu
iC9/cmgPzGecS9h2ehgAAmLE9gagnxHBaTd/RfqFbfFZ49EhfdU9By4K7pPbyK31
cXXWrqP7ENdmuG/got7lcCubFp32Qp2hkgT0ULnZjMGq55y58/8lDLnEa17zDSP7
DAFb+cT+fD6YFSGd3eM9Bk7ERojj78ag5kz66W9WCNdLYIwPRrMf3/NNKLaj8Zqa
9+lK6ET0Z4QEfU/4tO2N4J80aGvnLa3J2vcLDCOGLlKArW5/DrFwV7opYnOdJ6gS
mIPmOS7tLnJdtUDrAkmDMijqYrW6uPazv5O0/mO0osiiRWk0Bl2/hY1QL6MmkqWA
oJBZlbQNLvOSaohcq8G/hvEB2gCoDsRq1idmDUDc3SgcyoqpJ3eroGaNOPGLzNTa
b758I5aCJd3vZ3i929FwsS7RV/n5vtrEIyelDxGKtUZoFe9tjKrkSVB58/0raWou
TG3wthQWseO9IOIbUruQVeCT+9PsxQF/5203HHeTVta4PTTW51YTPsDRUr9Iml31
I22HHoeNuo3YVFXkuAKTRAG4Z3q/nOTFRIZb4tFf3DGHuvuBKI8++HBnMsIfrful
MP5/RQ64X5i0UgyhhAm14e2P6zr/p8fVs7706sIpLDLl+lgRQGZ/e4xEB36TN329
iBTpxFK/0tU6/LF3dJSyhYB/GyEDtDJ3hXScecP2MsQsCHu3VHs8rRnOKLXsz960
f6nQXPuaHy6Rfi6hCq2JQySvw0oQqMmvxaDzUxVlYGm9Sn2F28ozHCZyyEXTwvw9
51SNb8MzkvmwYnjJcozS4ipyngYigjzmWVZxlDfRz/7gTF+nmnpqS57YHD8jLyMT
xfigDfxJXSYRIOjySBaQE/JPQ7Sxh2omeDow17DhxDhfjC9oZ/uDepJpr7Ob71YJ
JA0etxWm7jr9GqAKkCJorrP2Iw+9sesJh44swe70knaT7j60k7FpTSft37uLkJjT
2NOfQRNxT6/YSu/Oj2BT+LbuHX5Hd2KPadR5ao+uA+LvpTYeiWYhb4qq7DN/Sd0H
y2aduvO0kgWLIQ1gbREprz1EuWMRB5Yio3pqby2MdiIMqKkFZtQyBzuIiKO5v5IY
NgdyTYyc86OgbxQTl77kcLVBxOgQnpm5oehlNcx/me136dAjTPAsev8YtGlF5iPF
WoXZUeml4eLU0eiwt3ao9D/XaqTXx/TtyvUI5lkqhaiqeftQbEzpvnFx+O0mZe91
eG6HLHGgU0Vsm8dED8wsvRCuNouugNsZYfM6+QbpJ7xkHyJk3Vy/9II2iiwAitBT
FKWB/kKddoGntGRcpGph8OtZdWmueCtoqMKIqOqyaULyqRQHyQ+4al+iNiehbn1C
q+fkW9a5si3BrJJokUwCPeGZ7AtZK6PqaTN/f/IeeDLI0jhK4icjGjuBsLMIZ1GS
snllDABuC8K51uJ9ULsHu9l33BCes9xTPxrxlbrqADhtwfqMghRBvZDOKaaQ7zwg
vj6NNim2/x1QlulSfqPVbUpTNk/U2O2UvUKJtNExCtcSrHSLBbtQJGF75xs2wXne
X99VkGGrN6TypH/aDyWtyQSK+DOLxbTA86+KvvhJvq7qPQhp+mkZHS8GKhYLemcx
err0v5PutYf3qM/kdrtV/Ae+r34S8No7039F7vprtGiR5/f1SsgPCPS6BqG2KlMG
ccgArPGRufhNZqO1G/cjR17HX+RDXm98OEVgyh0aH9X/5553RHMdKtfsV4atljfu
1AuZMo6qmu9Vwsla2Fai/cAPbh/vBJNjBeLTU239NrnBVsQh0E2SEQx1HzXy3iLg
hTtI42uu3fEJbfiy58hNJp0I17UrrQlbic++cK2GHC+eMzP9/+Hbv/YZyD+KU3k+
jgzVoRYl7vR427mDhpx2T/P5j9mzB6sZrEfNJ0cCHT651mYeBiyYCujURvEcwbqA
wDelj5I4h5TP/IqZUXyzoxmDImdggYlInWFnHleBGIfkt0WvxqN52GPkUrBRZnNM
z9j2/a9TKyYW/TQvJIjjZb5zPq5vRoDE6qiDBBELTDA9PI0E/guN6Ue2g33QqabU
jelk3nWUnVdSyGkBIeI8CpJaSJjdwSUQpdoG3Uv7m6MtlXXVH5Xep1g/TcPBb8gb
jGXqLNs5FjTco3fsEMlyOe/PGg06l+Famu7A74i6KeVM3Xgadi/O4tisemfvbjkc
+f/QbYgGxy+G3RHWjlY54FC5G8aiFjJWa+WBppF/rDHZ6PTLKs4M3khjlPF3gdO1
H9/tPy+juU6lPujaMy0gAymTkdvpP/jxspamkp2H9AGFUv/G+nphO4vu1og8WKgT
LoFdopxAIGcAd66L4kl2AZnUhox8bLzWfqfixNAmjPUlpmz9SSiVHAn5HdoNDcj6
N3OeKig900hZ2Ur5qnoOGhcssJChhx0W6MYnd6iRREYhtfTbRs+e5OsLAibA13GQ
AUl2nXnrRBPeyKrDQXH0h3cKuWFLwkPHW3/EU1pxkEIoXdbqojWz/RdZ7f8Wa/NY
uNgz28HH7j6kPmyn22BSZxnaW5sbKJKFWPvqLS+OTMJ3wDrW2WE6Bj31r1ap6045
uD3/IzmZCIJKeUWE134sIhLw/k68DVB05GZDRFBqA39Hk97a+16iFaBBwyLSgsAa
kfmY78jLTH3T3EGRVRIDRGUjljpq8gVE+o3zboJm4ytJbXToupFABDrwf8dBRcOm
nYq1jo5mgq+wjYirhE9B+BtE54778mXHV46FbHJjs7RRct0Br6LTe05LKhADt68e
cJ4stJzhS/rNQE0q0Sn//hwbPO+2rebPw5zauLWVUJt4a/kYeZ4qobssWKj9NwOe
Rbcu6NEl7gwjB4b/v+xW4YujSdRC/uyWv0/1BTa6vYKdCYgHXCMQUKWffaBNhGWo
P8QTQeBmqtUh0RNP29Vttf0NSfrQdXQb3KRWYWkryKa13DPWbtQjMEwGzXJ+6FjG
hy+3dA75p7Gvzi5Za42uQRJjIhl+xFQJuISWMNp8dEnCcXvjLGmOsmyzio9eubJf
gFKAywP8auiV0vpvM9diUjTbM9Xb0C8oS8qz2uZorAYneZe5/URYDBvZisuhwYbR
/wBt6Q2TdfATk2vnTc6vkiCLtWPRnHan3DOzG9ysvckh66uaMuBPzUs/OGmVOTFA
EtmNHU69knmwUrDDvM6aG9Qx4p0d5RtkFQSvOHpGyv90Pd7kN/jhlJQXETfX4Ozj
2L56q2GW7RKUQI75SV5ZWDOW3n8uuMvbZmqQHn87h9tjjHaB9ts9DarUOxRbE1EU
Dc5inn2YFKwQ8d9rUDX+e+2Vq4+HZgBpbHIt6D03IWhL0hLcKbVfPinwKXj+ye3D
vRoeCuKO3Rq6B/bx2I9zCv0R2Z92+66Qw7Caqq+3qPZWGWgKzDjsIsvfLxeew3Jk
yyWOzGSLnZIQ7KocGvNoD+ZypxrKcv0c35Nige06v0PqJV4yQP6rR0+djiywIAeJ
Bj14wUCvFr+rNpsdvjBtZZzxVKMOTEZyr4tCe8Kat4Kn5gzVcaZ3Cdy4GYcwrWKq
dsABDmYe8bcE9EFcGdx/xxDP8RdgMcWYsPzE+OhNbCc66yMIMESuMdk6/9gvLnmq
e1Iw3vb0XQtsYJ7IBGDq3Rmxb0a50lRW10qGySf5OUI6kk79c+bELAP2fHwxfmLs
YzNCUcJDu5OGFIDMITJFbMrEsCKSpaw82H91/ErSFCUODtqfognLLhplKlJ1FvUF
Wz8J7TbhCZurB5J1nH1MLVHSFQvKrEtBi5l7ftQzdKDQB8Ea59oXEc6ppyG+FV7R
VnztI3IeLdUj7ZhsybV2g3ug6eWwhzgRCb23792OOrMKFQwfum8tUvD84YmI+rXo
6/Rv3Zl/ycjCT3BtAz0+xqlYd2ctRPcKLQ1Ba/F4KWvmSok2hHL0LOWl0TF/REvQ
II7MqOo1XQR2xXFMl9wupO1RI20mfjvKincm/9vDQXo6n9CMwl/3fTkfRN8yQE8m
EPcSSOftxvW5Hpbc6DCFqn3kCHcq8jaEf5+LbFTd3QvjyrR1n2W0slm2B00YXurd
4FgC2AnoRNrSTFNWLylCizrcsVdB79n75y1Sp6LEI634/HghhvM0gXaqGYmJzJFH
NH1ENbcfeY296w6f8BtOrHG63GdGzAkNqvuGxY0E5rISkbpgGaPz0C8zDhgCJBUz
nvyBzxvh2u3E8Ao0143pslGgUT3Ki4EEEd3dyL6emKAkx6km9/YXPMt1oxaCLFPn
RIv1UKul+etgPOgngDnsygjWgL8nvPGaEoNVk0tiESGqKmFjTS2eBvUUrnIveBTE
X29aqbyom96/1qF3JpTANU3do2hWYM5AfayZfrb1HALskJNK7pgSWAHkJYNp433F
gWl0fs7l9o+BBdRuk/CSPFPhaGhU9T2ZjSNWgph0CUGBoTQKL4GvP49PDauK4vF7
dpHe8rWqmoed9RnxDYx1B3nwD13aEQAo47GrpEJUcmjGRa/rE42HNY9c4hHdDhff
Jg7uoOaJiT9E6UR7vqzWIVLq1kuusrIxMa+Sk6iZpIqZ6Z5ZwYrCtdVkjA/e/rje
GlQnalm97T6NmikMT1clHfcU63MWpfSbYoO9tyTOQkTpapVx/ZcQTw7hooFx/rLa
6g9V2Sg2jaxStuTr7A3APpOD7s45Xyv0v/VoiAGuVV5QBroOMz65jc0tXC94EZ3r
CLONJnl0/GSgobJxN5wnEDKdPUippksRV3Vi1Vf4LhQqhrlm1AFjkUMyX06ZTFdr
+j6LwuFnaOctrimqPg1NpfeQOlz2bm9Z4wXTqh8IoLgUenmAaTJ1ecJjOtZnjWCA
sns1EOrNhMl+obGy/siXg6Blq8W9xLRYPQTwWzsh/xoIudSyM5ncpXCrTajnApQ5
DWGp8lfLUA3l4KwYxjAyN9rGiYQhCGZ/jUJmQ/OAtUrYGxNOtcyxCya/bUJLIEVH
+3otqWUy3sK1U2Uw7Qgg3XafkJ4s2CLF1rqyDkxubOylIOyX+oVCQcqr8Qd84Ggn
8LPSx8Gjbk9gSoIoZ9DSeKjkS2Zi7CapXRXC2zhT7giT5NRZh42wwLZTC5aspTjd
4mBl9KeXuxyFnsVDccB1+EDRRev8OY1un5CK6/Gjx4mz+29z1IPmA801MQ69sH5Z
MJXhJVeniYlsO7npkZJLBnprk9s6xvMoOdiO7X8GXRhbh4mZGzyr8P0lCFpQcSBF
7AbhQkf5Zj0nj5KKxVL8+f08DHZPYlosXkt5KtEA8T/jX9OJDZC1KbQCAQw11z7N
17uxgBK/JPiZAQTY68rwMSaFFUi5kjVqrJAX4ERXkfGAUfXqny8Sygd3iSoj1YUy
Zp2SBwX1PBfgq0jjMKDnepoDUVW8cvR7xeQDZ2T75xig1IoyUHDyVys8XXEwo/2F
43nbMOf7/8TBaFRtRpwzjhdAUWoXxK7/bWdm+sTLAJ1frdjmpSS1AEx/L9LqWUHw
t+KdKhrx/2Ttl92TUA/3aPqp54nmFQQA4MSKsbG/1LCcaAaYOy0NAn9+F4/mOoRE
LYYJlNwqUQDhkaQgQz0TK6mczras607m9wwcQtHH1Ck4jt6nFvXX3ZVKf1k2RDqS
9QQFpRMGzWWpjHNeMccdfifGg9XbJoahy7kiwKczDC8CfD28l6g3ACfhv9T8Jkt5
8cjmfpVSNYBzxBPzI72X+S1dUvLlpSxacD9Fm3eE30H6nwEkhmWgkU73SxPDpjOJ
y9qEWPf78p/2e6v9esIsSetmQxke4ujhzLx/DbyZrnOm7qef+0wTHL3OVwzYcpWH
rlw0SL41+rWrO6OEsuAd+DwFQgPhQZyvtFwn+STM9L8WXuu7f8kJav35jbBdreSe
zTfj27vL2Nsdrz+KftjXQkWQ54fZG18m5TT+ncI1kbLUykI4GvCXtvgyUGzhD9RQ
iftq653NLGEmE5uVG9jNj1caRY0sOC1JKiIctBnMExhfsN+0BvLD/jC2Hqe+WpRx
HsghP7gSYEKCX8SwHAjZjbI6onIMeLJwR1SwIMgi8mAumMEnxzh9e6PwyN9ybj+Q
wnZI80QhjKd9BEX5nZSE70TW0J7Cu2NxMN40RwL5FLvYK4s4ZJyAkPOoByxOHUqA
NVWsEOwfCXZHi6DZEr9CxsV68pZqvFsEUS9crTt+IIokttz538l6560xax1FFIs8
3KUDekRt3cfl6ZJW1JMN836ljGAxki36tFH4ldQFBQOVBXp8lgqtTViyjh76QlNJ
opUb99wUg6G/OSjVKclLSERNinzbENGdLbMuNVkziPZUVTdnpKi8NuM7iihruaba
k5+QFRvYGsh7EBP/ls2fE1duOYUZKeAK3nA3NDbY9ZigW3HYrrtZgKs5wPl7zezn
ZNAon6F0fyjmFtp7Sdxba/veSNASV6yUBgUVrxb1QLjAgtGeVadQtuS88Yz6Lo4z
bnWzYEikENuRJ+j0a97uZlPXsVU2bR7AbEOUi9g1Wdpn574x4q/GKDzpFAozz3YR
JExbyrMyEw50BKvJ7GsKWVQn9YnNoa2utgzzPI8xo14xLrU5YNGJ5mfd5V0gL/cC
pw0FzbKaC/qiEZ1SJLz+O7b8Yjhi8gO11J+ebXj1e2P4Tr185yeBlY09x18twg32
A5xBWw/8N9IV+Zp1zE4VlbOSTmD66JYZSGofbXVw77u0t9BAd/oD+265UNsh3qZG
8j/aB6hN0NJCraK3b/n1IyynJo4aFs2E4z8yK5FvqyGvvS4QUcpirh/dUq9qn37F
qQYymf52IhZD/xHPPdqHrxeGXVeyd0lmt28eUlUlnjtkELLF27vOzU2h8zWrYdJk
5lw52xnVHAzvYLc4ar4Fb82m04t79UiQ/FBntgXQXDsasPO02EIGjEZogEG+s4bL
hKqyrLPWdlqEr9BRKHKeAJqrBdA4QrER0XalUBs7Y5B3PME/glNGU15KurjONi2Z
s9GdtADtUltbiuM7ERrn2JRENg3YlWOIvsF3CWYplBcyeFyGKsyLgRkLc19stbLA
o2ClFN0845QUnVOryZFhB3tyyvFsMjqirsH0ibHx43tCFxS0X02Pl3y3TIHYl3zy
eUi+pQriQM6htiboUXoyVko7CykIpCoTXmaDhUNdqeT8ss9pNmXpreelYsPS4Iae
ImJ/hw8NrQ6DpTN/nyhDoql91V9wH8//rIGzNoohHo5cxuRltvLXMDO8ezV2kY4i
WxMf5+R7Mcnn/0XYq0vPhnyX9+hS4+OLHJUWR4acGty28+Rk6aGbSFW4sYlmvlkU
yRo5ql3iWU8wb5Oxzm+DZ0GOrUgwptFI7Sa9Tw/dfFu/GWciCER7MigaWk+LyPJ8
IUN3Op2UHCkWwR8KTrLnn7nxOuU1ccMe0v4hT4sWEIfcOjUKM/YKNT+IMM4X7XKD
pYKDMl3EgQOFFHse52lDifLzVlFN7tDrZPKyzentxEM1uMCvON6SoldcEi0yqDMi
zQqXAV/vcY6XmJ9/51qaFfytOIjx83cApfiqEzzzjvVsD0DH0dodgIx4VcVZdPJ3
A4tWG3uLp7+i1m1h+UeHiPdEHwwcxQFxdEKA9xKcO2dZgRhPMixTYYwrJVnHVOWM
OjoVZAGpBX9lbf8uQCwfr8mg4mgZ0iu6Yl8Gl9uq8OvEAfhE2DvUdNI3mjXHqRmu
iKMSHuW7VsMEokOLPGftzYxLrROs5NY7yw2MMQGTKSPsJ1haNJpZ5WTgrSiizyDJ
sFOvbn1pdvbqBa4///3i9gKXO2vznygyKXQvslUdRW2U6Nw5o7DOzLeeUHS/RXi/
w83bHo4s3pe1ECaAwHrDxtj7rdOsA82NBijmxjTJdjrcYIw+CUh5sXIW4n74bfO7
V0lSwfOQsA6N9QS4c4K5eGuY0bHxal5DD9JGY8ui3j6yqevWvBDtaStpPPMrQVTh
qq4En84RMfCL5Z+HaVY1HXV/CSAoyYkTEtAxSTUCXaJo/vAX1+8u6yUTPtPa++Nx
lTCn6KKfqjG583a89I90IWel5IEjw1avtmnVdDWfIkM9nu8FGL8MLjLIQ1N8rsPG
O9/qYtBI4PyQY+Cgdt+ysZk2F6t3tvVVqfR84sly8ppS5sqx4FMQRTWecNfaiNrY
K5czx3LtjJWt0jFrKQI88rXZWni//dg39QP6Eb9KVZ6NrEYxhmbC+Yf1JrCEd+jr
jJBXGJwHfpiK3TzM8Du9TSYlN9MuJIIKhKfuVfS+3OVWT11jg/fOHsS3y6DaE683
xgeHUf+4Mvjm4xzTee30vlnf0ZF0CtWYO53/soQyaXDTiu7PgQlR8lmEQqGfPuVi
YdNJEcwk6V/2tyil2pl10xdU3fkoou5rmvXGtdWiWDW4Rua6v4XaRSnlwijiHdCO
AFe34cSwVI9dLfRMz4UA5ZEfqYvSMX6FvrG3cTtO5jrcuhCtMAJu1sOBYApfLvIF
RKkQtKdmGpkrtYuwaUr/Q9ZyMfgt0hlTZr+DNwqoqTbvrP7xoxoxriFr6Qb+r684
xziJhgOQwwdJ7dKLmfaLLGJTX+ni8KkEOfyVBEInXfXIjnaxuOIKhVLNICXFQe5p
/UUI9GZSw9CCMjHRkas0FQa3JyTgn8/4u50s7gfJK1K0CVYP4iJw9jp0SI+ua2yb
vrC40EtJvyWUxjnJMI8dXb+rqDHZpGB6UoESfFyuBVhpUpBv505XIaK7M6Ys4+R+
DZ+WQIqjPVxZseG6qDGqS2JQJb5hyAi+OAixGxjxMUmdYt8ax5R0oG1BQDFDMuLy
iRFES0VXWfXexxvqWQkv2E1djW9CqPc6UI9MCUB1jJq5MB0IiqtELKHzlMsCR+Pw
1Z99j2hE5kl16wy6w4ZR4pChqZNDvJ2uoWEcOBv8+HbUoLA8eoemelm8ejKUlbm2
QJhpI3w0TgNIqNkBcmUKYW9HSQIDNLv7zwiuok0HZaSOVaAkfvVMMHpY+5p4mMnr
Rowy4MTD9A0GnkoF3/XRHadsafgtkA7td3dNFdOI00Rx0SVlN6psO+LmT05qkwU8
E7j0N2ZFdqmYYF6PuUB66hp0V5eNhKc0tFHuCn0L8pyf3orzLYSdTO0TPpS/U821
RBpT6UZJVk/2+U4s5nw09vrWPwokIW+xODUEl6o87VL75fzi9HruWJOafp9VEuoD
SfN0sH0kjveJxt/Vy3EGq0ODgnFdFzJ5En6JX6LaW7lxByBFCWQsU6xGA8JElAJj
2Wtp343us41xU/vuyuw/+bx+TR/IJz0dz4wRrgB5E0TCTBpPUgZhYUpc21MdDj/Y
MlnbS9NjkLiO8RDleKA59DLz0BkZuUCiftyMUecC9NF9TfA5y6ITcht3swMQy4vx
a4adUcSp9h3zgfvgvgxm+ZxyAoxw37AJEdnE/S3cnyXaEGJtZ3CAxdoPO87aw57j
/Xk8XkKaVILf8969/CxceYSwARhbCXVn0OzGSWbiOy59yC2tp/lVEysHTN/4jN6j
IdFiRNK4s0CJarTs9IBLXF9Ag2aaO/gtzvDHuwzv/yT2Lumj3349edTsU9qM4nJl
fTk+4t+EuJKP+anrGN07CtrhbucLE8amvDhNtCaL4GzwqeZM9JouuzJ9lf6S0uZ7
fH0sfB9gsjC/bJ4Ix8vagd+RcLQKYND86HkyBGCecfXkXBg7U/pTR1FQ9/U+tt6Z
fW0HAvcs66JA1pKdwnUZKINc+TcRFqxm/TU7fqUayK5HZ00Egf3s2v0CsB6w0MT0
dp+Be5bgWv2s4Q/aeQiB8sXBjr34vFaBU49b4Poy+Gv6qpqwS/jp2ayxCHCVq2M1
1ch5c2mvWZu56rsMkK65lztBqfs+grOutm4ZzBbRb6cP4VJO2tJNYTEcBGYa7+4s
sXFH1jAC8lazEfLAd+aRwNyi+pCeGrToNyDYC7RtPtRqIgQVdzBR/6kGhachfnam
pE8xfyIWLBMZ/o0oPUJZAfjarZ5SxA7CSOJ/oCHY5RvR7BWA8xwbmm1rkIrdSPYM
GX20Kq8OyW1pJTKqK/ZTd1iRAUQUHf80Yyx6ATAjOQb+f5nLTguDwrg10qj2/coP
zn9QYvrDjnyTYborHktxn7v08ynLMDFjV9hr2+4m2fnObvvNCPfSi6mA82A7n7hY
L/M+YaGH0BqjwoyK7es/tVSeba5GhXdgI8jDO2BMdxlVc38etg1eWdXTztlzDF41
AmKe99+B6+1ZSaAOFdATRRradhH0f0DgpxceZJgWLF6WgMO6y1Vx8W8mZgbLJlVP
5C21t38Jccy6LTu4MujNR/PY9WAplJmp1rpxt8qI6EVvWH9HN6lXNTY/le21jHds
RMBoGs8zHbg5+mkgnBzHMCSY4qQ2/FZG7KkrLlLszuxnJiTH+NPWZkA8GOZ22tKf
STcGaOUduL6o/lW3KT0pwpg2sud+bWyQnqIXFadCpuhALXY9ymImeon/TM3btiV/
JXFk+g9idDYK5yzq1tCfTG9G5w+qBGV3VqmUlVWRkcwiUlwY9QgS6YxZAHVZxPHe
PLDRaPQ1bMuPDjcl1HbyvIGpSxnbfh/t5LaNsc5vDQVUvMvrPWkvIP2TNtAqMyTR
lVr2aLY4lKowaQpGNR4pWsgXy2qrwjHIRuqBc8YQLKK3Wlzzue69oNvp+J7Y+WHn
0cKxy7OROzff6S2WakHg3p+17/YiVOTD0BcqbFnHFlEUBQgoTn/fIzKtknTj0Er+
8gt1NvyLl4SnGPdoueSJV48a4donWdi99NwFa9jTeZoFkbJJupqudP0yvD6TVjta
0AWhWhtuFB2oV+mQ6MTKoi0CRg4JT/TPRg8meQVP1DXhJbkbgw53cnQ746pciDsB
w9lV3o5iL+ccOdf21DOplm7+VQ0VIWgV6v+7Nmr6ROZ257s70tY9FnFbxNVCoU40
df5L1DTQoisV2SOXOF0QG1cz38OQ31j6NEoViohO8uJ0wXjU9Rd7MIpwq605OogY
i1flk5pe2xxNaooEZbUmAB1LTRGXyd12sRcIrOF5VTP9VHQnqoavZdEquIYdcvPm
2/SICDGmRBBSMAd/GHu9DQbJJ8q8P3XbhljxnJxfxP7+sjYhcJWzAGUkf2nsRG3Q
JcZuEzc68a7f91Bnvd8Y0GRwbvsl0BpsEREPHcXqBfqKDuMwwCckqtz5rfRiPp6D
5SSzdIC7GV4K3GnESiNcl6cKfwqCMWlEewbOpnQ5nXFXTH21kVPt/uuHXl6Q8Xc7
Sg39eRDqjgfuD5MMcx6o1TiBxIO6Lq0S/10P5wbo5IhewnoNRAjpO/fIYceD7891
/zi3SWjpQ7zFTfd/p5Azcx9eqe+8bIo7n1AOyqsiOST+GTwv1rPtGkGTLIrfk/Vd
VWoH28hknvZd/CJMVv1ZemjufNrGc78v9c52LW29MaCD1HGK1SWtaNlmPU0smOqj
cquzNGXJeeO09rwvXoKKF1OTuspIKfoaCRr96V5zk5MeC/vn4FdGy8x12qvHsvBt
Xkm8abutqflC69DhnuGMoPOd541g9+CEsTGl1oJDhisyeSj5dmhTGcVt74IGXRYI
IgvJg2ZuPfFM6zDw3v1hax9a4I+4PE5yVASB6FG4mvyJjR+hv2RI+qwnkA895cIe
Mq51BkmfTS6fzrO7xznZhboOY2cv6/U4/v2Q+r+Y0rhKp5ZerGrjeGqCJRE6P8MO
joup/GZrxGea7d27wdpS8v6m9Nc5LqIMsgjribPx0KnNPUXEwjx1Q3C3H7gMLDI0
+Cbx/Jf5IzkR6ygRMlRC98r1o2jLVFcdZixXIF9mt1KOLgVgGyYFuRRWAadb5Kt2
Kmvu80VC8lG72QLsyHYM27HntjbsSNCNzTMKjlpOcpHtSXKAtKGgRer7dQT8gcfB
0wzXkvbhq7S3E47v/M6X2QlmpYHMkczzaO/6XrtWC2+a59oLg0Ah0+O6vvcp/UwV
T4IkUKp9a/ghbTQ3qolhB5V3JQ1/KgqASVRUWc0fcqyQNSnGpFhTAPw85dQcP4lU
CyXjVUSepEwvU5HlSIpDJrBEMadqLBo7bnOBQTXIsiigx1t1bl0yecjjX6Gnb13U
kv4uDEms9qnb/K5fwK6FM5u0Yur+1XVmIca+jHnQfr+8op/gDTgtYu5fS84hhX97
oz2FKIOnRsjPUC2iPO7d9xgrVVmnXsq1FZ1qydfUc7FixYAr+3Ex/i6lWdXIELYj
APPgVVd+hUeKPLz0++iXPfV4KRretQetd0s3snx5XmjIGxdpi3NHhl66aHqmpKDN
JDWRTrVITxIEK8/sMgfcc9u8nAbQEgSEw0KClrMBhXFSTfqYQk1Q+D1SBjf/vNge
cj/GY8SrfcJlRs+2eoU/SJqN90nzufCdvB0cApfuixW03Hp8DmA3z96CkvO1n/DE
52qoPdYhptI/Cjg+G0cR6ExEU8iNDapSwgAwid56EMtmBoILIHF/F3e7kxJNpgCM
YLQaENdHuEcGBjFnaYnq8yqjO/FhKcZQsVeyqyubCI/hBegJx4qEFQs43IYcAWcV
vzIPymtw+hgOqOgBtk0MP36qKgGV6SWSVGzTCN1zxeog9XA4UNK4DjxvKJQT7326
nsPkRi90oMNFozEQ9jhdXBeW4qt96gf56haVU3/ze373Yh4hD6hQW8ujv1mkrG1w
suYHxCQRTuuL6F9dGMRTLtOeVk+pIhJErDErA3vd1Fxo2/ry27A9VBBKXzdSRtFN
v20/itR8xjlbJ1DOvUG7Xs/O1mzlFr+COY3Q7HYjDR8qth3v4KiWNG7DGcushG1e
Qj710SdQ52Gegr7ThkcDYuBhkmKYHSNEqd38Nl/DKGc9jRKSHA0lS59dkJS7lPZ4
XoBZU1YQZzLYjdcLcjgSItV3OvlymSSCtklRz7gBuhTuJdg7qi+2R3x3ksbQh5s8
dW1ASOXdvqaDEI8T8c5PaoLPY0Gybnj8PhsrAvF2iMG2aZceacB3JXyte4CgYIpO
QTBt/2i9m5lFzjYCFawhxPmktgDaazC95VdMEelTfwLSiMbK/yma+3WsAppxXUhp
rr1Dc5LRNbk+/s6/lUsUPm2O/+Womu3Wnt32j3cezao/mRYZnGn8wkQj9XrgQ9hK
nUeWGIeE9fPqUDi6PnA7+kQs2KQUCyKVzrJqlYZQcEDFaA983AxLTlDhNtRJfuJk
cDdfpY/HSbvse8JhHrhqGpsGhWlWu2R1fisR2RpImw5y1hZ1ZumsQQ6lNvIdcIbg
Tkcj/+vvwe7GgXZVXWpa6baox77MViW66nwfAa6N0Fj16v55AK1+XV5P88ozKqrr
qCFT3vvWr9VY5XNUaNoWiG4DgJqLA2xFw9hiJxdpS4ehOKsn6F+lQd49Ucqafn+P
5QwGS2izla5G1aYAPbeMVmr7/gr33W/HuDo1pEVcvjSVtTUKZnRQYv+ykh71hpBe
CSQHMdeKxx50WOtiYs+GZRWW10xZ8L6fV/efNa/35T9yZzCLwFgF5mSgoTMFgzkQ
ZSqNZPqjWnyFS6hugybXxXNK/wWZ/tm3m2BJXadog17S8dLVH3p9DcldEx2E1F4f
5GqTdbW1TJrCBx8XTywDkfBDipHTzHfN2hzyFlr9CYTbn7v8myF0WaSedbI4MTU4
pW1X10ogeBwRhUMKVIaJDQo5798Ur1pZwYi87Hbl4O7Payge0N35mvZ5yWI1Qdhn
x8UihXKCbWUeARgP5FK7SWBhvVeI9YkT+ZJ2wGlcn1tOHC983A2HVTchKkSohJVC
0arYWjSIUU7+x70PaDk5aRWvY+Eiqy086S2VLyLJ0j+0KGU3uqF73rigB+c//Mhm
mEFZKe6lT3H5UGBfK2xW+fzsODrMSd3si+1UzrZ/REsFl337FUBAHlRWIzZ12aI1
e9p+ENYcDeRkReAetPIcm021gdm+FGebWRSu1gzo03+Rk8vd0VbPnAeKLPnqaYPY
ZYMaIhUQI88n94bj/Dvp6FTSqos2oRngH+j2nL3W7kgDSd6xDEnconLhVFbjwKAR
y3MSDwydlSMdijSGY7dmvcsh9+LTq1tRkVQkBCj/XysCBuIfiseWrfXb+tZlOoCQ
4pGxwUtUZu7GTJu7qPiwpqNR4qxncfDuLooI2a3M8DHUtPJ0rz6Q3e1VMhpCUB+S
j+nCqrf5g/PF7Or5aGpKSTQKPxaVb6LltglA5R46aZxbvaDLINRDhON4ojbsainS
BLar2IaKl4aXEkTLR2gfWDQG4zuiVvU1oIn/a8Vpn8zZnWIBeDPePNnfAkSv2K/I
cWBk5ncu5f/No2qG8IMZlyMa6cHi07Qz/pRxkF1zuvIzJ2MATNjGuq0x3FCLXey+
g+a4k3hgOCn6NUnK8YUuy+DS9rvswEDlVFQbnCRccPGCD+okbcrb/ShAVaWa7mPt
gt92oIvJjI41TVexTIsG5ID862Zi/uglRla7xSxoFcOcu2C8qSMokERh2HQRbaO2
EY2kK/vSuM61/7q/f5bUGDUP97Iwl0/XWDQuq4ZLSxLYEy2L77o6xi8DOENumnih
8FUlyXS+CdWis2SjmicWbKDC1lJCW8CAUufznR2lpXFHnwn/L2+7eG3ooeMxIMNw
kRbFlGHGd3UCVWDISVMy7jr60atdM9B2IcX1RuFHB8OpJ/iuZr8eAr3CyoOKxVh1
u496veW4DYclhg+ex0IS0LcQDn1wyvyr0xra/Ec2e3Oe5qivwD4d43NsX9BkIaPc
niYicN9DJe01o8P2TyXl3Pb+y4aRwmjYTZOxhfuXcOmXlQJLY3k76QTQHVOGFDfq
2J2PnO8oVarHyC1FcaqU1vXSfn4XbUJi1+Xf87loNL2hF0XZueGS14Tu6CpYLnjU
Bp/hUqqmhUSJkGee24hH98zy3UUovpi9uiT/dPwmtHFBXR7Sq1EMP3SeyOGVLW6H
murf9Ghk9+67gYVv/QQiCrBAzCwjZ3Y0TAokhFRIPCMsLwGQpu5QHpa9wHPjQyJT
LXTGHAufvaEbRNJnfSgyQ0oPfWxZtG2Htko/JaSd8ZNwruB/tGPFcFzp1zSiJ73g
HrPqnMN3pSIr8/5/EeVLUXkPlUtFvIUPXtsB8OYLL/+fYHchYsi+35131BP2OIEy
jZ7KLkC9BjP0SuunyDz93013op0jIfL1Ulf/cEf3lnyT3jvu9OYLvMnixwWsKg6H
HlJ5J+Ct/gSPbEDN9IGsuODqALgVkhHDR0oMgCo0Ha5YEEe8Hej/uTdkOQIzuA0h
IwsSozEbntwklouSitcYmW1HDGz/NOGWRSYoxrA28uVwsauvmdou/YTG356hWe+O
jhqyAjSKuILUxIO/HMEDnjHfjntlh8vrF5xDrfCcZsBjPj4C0twNDpvU1IWPP0gI
jyoLEQEE+8tp0uggCX7E6mcZcqgqbGUIyKB5VGRZswk42yWLhuROeuhwj5j23eq0
RSH2ENg2D1XkaLAMhLUuJ4AueQef7F72Nm2CUrn2X5NY13lcPk8T5avFu7XRp5q2
yRbyXrESwUOvjqvgfybv3L4zNVuuYFCOYDrh6gJH/pBbzwVb0AGwuVrdWP+KeB0j
NyhC0Tl/aDogEcpc+9YvDLOEnKs27772SxS0UqbevWDwZ7MX7vJlcpi4hla0EmML
8GH5/7+AOfpvmRTbaKC7+qnB47vaHVpFAN7SX2BzNOUVBBc7ODwqPm+RoGxiFBSu
Uw8JdEjbwF3mduk0HA5U5EsMqQ0brPeRXoZmh1zuwehz/1cFDMxWxx6YrS9ITAKx
Itu1Z+xt2iNVTqeumeTu9JQ0Tub1xalstAVC1fwXLMW9y/c8bP8pSqSKa/6J7S6V
uMWI+jhKadYZcTGPuyxRZ3UdFqhyrAJAkP+MeL4LPXNN8YOij6ACB7alKvzHu1Zb
s7ev3Zk4WpplKqjpXRuTZWaD5BE0gZrA85ZAu740hVkuaBE7vSaQTyAge/LbDpv/
MEtJHBBZI5qGKEzCkC2cqOiVL/PwVOChBucRY+jT/rIrOjS72kQQGD0fTCKBs1xN
2DtuoXmtzPLPT66x6VJN4mGV5KJcbehNSMeEG0f2r/kx86HOqmIPcVXS1uIdASUH
cFpAFmDoTxdGzQ3eqhZeRaMk5S3NtdyOxmF/kbOkrNObAx9NAsKmKqK5c1Oe+8m6
UPYZqxa5hFBKhv+al5hkvQHFFoZ0D8AeJpq+J0cqljjoTiLfXbR8sEi+cVlzgQML
gbAmicxTSjlLnoGJ2IVSEN93+qci9ZiDslfcAwy7VByftlQoDzoDMc/zBmU5YX8p
fxfeh45i/Db70u8vnOw1ti3uil+/+u6/EBXO6kghPc8ljFuTkH8lAnap2cBG9CCJ
WNermKgd/eJuFJkGkJZum+sgsR0cNVkRucLIqs8JWP4R/ceZONoV0ZPDBuXu/GZM
jEL5AAQFFYnLZrHis9ToZ6Dqyobc+R0MxFpdy/NLzPBmwDguA2W5j3xZexoUWRob
1iCFfbKnQGB1yj9LY1T8KEpcJNRsebr5l1jHgz3ujS7cNXYMjZXC1xyCZzsOWW/n
k/PdONWYjiUWTTdmxAa5rZsE2xlhf8Ir1DhtoWBf8o6OKeOsqBnnj09WrS/dsfQ+
+Xah8UDZK9OvQX/zakj3AHZmEozm1NZnL9hlhrHTu/pQSna9/KwUJDgzkUg0OAQl
keYzrYis0bUl7CxoGgTHgxFxvaywAASYGdHB3MK2l3a/8PL40CcIM1MU7EGR4a2j
03CEIAgIrEEtXSF4ANygAC1MGQK9ewdA8F6IeQhBR0pVfYpnxp1IhuN4BJAFXIT0
ANzjWpPC/OKSijxLngUZXuMyKkMSdvVQYC9TjiGDqhCZM01ijSWuJBeBLQ9IeZLS
qZ6qj9/38TRHBnmpR/+veqIETFMvez+b3fxaUMcmiDJO32u1p/ABZKXdSc/AKpjP
9Z5g2GK+yItNmU1fanD/ePOq53eBb4501WzgxotichR4ezl0hoX4Ev+fsisOmiON
5JaIaQxskVPhBlwZIGmD8X7N6mqB+D15Y68r8DDPDADjcS6zz8BqoTW5ywgSqZKc
aPbkmNG/Fg9mH3lXgkrUuLHqVWVc1Ao/PM70XqelgOqaTHxdyh5y2s7A2TDeQ45I
bPPk7hhEjQR9/jmOQAcFR7THNGTDwtFeioi0xh3lJgs0g4/2FtXFtZW3wBk38fyd
htTkzbcLrQJj9OBNyxc91sUVpgph5XQfpOu5xnrAxkq+ChCFsloLns86sjGEr8HI
z85/5aQh3rwkgBJEhKZeoe9cmcKnrT2LOzqyyIXlAVymt2nmcfyZVCS2cLHzQCG1
uC49M36QkqKTOpi5aKye6/HhX7wVYwE8wWmAV+opNTRHG87NBxTJ4Y6Pl+GPT0T4
8hGveCVEBVKXFJ0GBlSNDMvNrKZo0bVZYWULNeL0lxTi9eBubaiBoWHwSdlmy+1E
LaIvYj8IBeyLFrpbsfCvmOUHephCraqbbkOgOPzCpzQpBtW2xMZSrL86BPwh17CA
tXWCAjZNeA+yBhT6TmA4wVe0woppqUoDsNOgr9rkXM9FhVOWj9+wEJ/0zGWuAvFg
gg28v6G6JrpNqIbLJse68PsHPflyjjsu2nwOXzrrIinkFFloJwpQPWvkSRVtNOmb
ogSc6n0CmDG/VUfdCEQJrENiXNVOLjiMHgIylQO3EYNUQLKDXq7lKVz0K7B5GMtS
PgDOADNbPiL7Fgag3B/H/er890mPRB4Y8rP+GVewXUVf8rn0HZ3msTiSjbki73ju
HDn/wX3bRl7/h6mZ0NqlnTFBeSmRNCfOdgjvul8SJTgtl+fd9i63kMvKB6iJ94fz
rBZUBYZPDuJPGq/BSKhxcfc/nyLvmjUT+kjliPJoxpE6wnF7e6b7CxpEVk/EfbrM
ir4Sd5veoxBVAsWixolAPX6WldirKnhpOV5SOzDP0vkp6zqBNjtUnuH5dqEQtr+i
bNTGFJLQ1ZUubo4CmloU9cGhFA7OOjsZR6ovk0TE7I0cmSPj8JKOlvu5zjp00TSO
iRH25o/Gg4U09L4WC6BLYQSfjRuFEvv1rIc/LoKW9kwCwQ/RDofc9eirzzUIpHuH
gIMFFA5e8hZVU/BNp3stAsh+ivJwJ8N+NsqhotxLXkIsVaZibhLowegzdQ7gLDJY
X1n8lV7QoUH+96IKmA94FlgO9gfb+rEm5Y36JAfTtIoB+3Wtxf3bkOpEtOYrh2qL
BA4WyBbXt3UsRdYeUuzzwuzbL/+S326oHcuAkzPlahjzpofrPGWjoM+Ue4GuQZRF
vqGzSs7yFgh0vE8ciHm1hQyUPWR+ySZd7rs8/ArjoXS8dmAQwUsZBVlpDn8joTRz
Xa7aNduKxURB6u28ovUMdITFbix1pVELfPQUd3YP31v6hAYDSrpwqgkdU61ZBWVt
MpfGqQs8UI5WPcaqk0EKVvLiFS9O/U3+6myJSThtI3LoUBtwos4ok4XjK8VxURZa
R6q0n9MR99kJjVsXpEbye/MRo8CYlowRB82phl55ehG5QToy93UKiTkhDGYPuJyj
iDrJn1oAL7HqU1Tu7Gj8l9FQYgkvId4mR2k8fq/qQVT9Jo28xRJcp1SH/djElxrQ
DjEh8T3OGgWen63VsFOmrtVM7j3CJLMpBqaT7rtp354ITkCN9XzuM48Ip8La8aqG
GFO3G4DfIby6Zv/ojVi28Z+JAz8n6RcOryxh0BJyjttEx27ILv1SZ93tmoD3sO+V
r330IevX6XuJddmywhxIEhYtROCAWJmsbyjdhE6bJ3jZBaGa64mbibewLtlE5v40
bN6BSjrcaD2wktKdc9Sq1/1AmShjkD4lICryYd1mJJWmg0vik9wgoOv30UnQi5ol
g/mhyW3gqXHg+8p4CmyvSOwFxBz/Ceo9UgifXG2+N6Qx8JLNJKeBMuHVNqyn/AvW
pog3Qimkkuv0Z1kPBrFPHuoQO2AlY9cYtsh95IwTKey6/IeeWkSezSNP1QvvVala
tVIcu0Vd6wKgIVpbETywv5ELScwBXOEHosADJKSOldBC3v5Ahw87FqhURvikROOU
euAeqhBEDML27JnxE9VP3T51FjP7GKn7KbjT7FyJKAQ0RlrJVcyluV36m77hYv3x
Xl7JmwBn/vrsRHe2EamjCYNJPswv67SI1WH5o1QOpbwWAhGAH8zHQzB3oM5GMNbj
5YhHKq/msFlSLrRj8O18F1PBQDk8LyRZ8eDxtsv95xlwYNx5ck2n2zYXibEto4au
GwFkuu9ADukxvOBWtFAbYRQLYw4M7hRZv38niaboy7essE3eB05oQJVf+c5YpxSN
p4VATgwbiJmrzHkcOYzGStRO++qV1MKFyAIaiTjCEvh4YhwhKHeYitjkqv568Rhj
HlqsN+1MrU1lRbaUBCPQvYkkj8BQ2efDjPZl2jLDD8f75wqI6aFGUBdmraMMKb27
aNUG5YWNYgdxhR8aYXymXawSRpW8IJs8+t8LZwahGVZx3niHbnfm45XRV2w80PO6
vmgobEqkpRw2Rw73UdkPe2+1Ey/Z2dxFnyTFZStr0wfo5pyusEpGVa8bgeF74AMh
xMc7xU1AZ0yGWr+BCEre6XdtDenLrItynsdTPb102uDldXIg7P/ACHSKl9gLxP29
z6DS1Vsq6sO/HVRwvH6I8SzdX0bg5RVsz0qYwVkvUG2ApK5654F1u0AjJAosrufA
c2M7KBO59efwk1fWQKK1kEIx3uCplxHoo6GMFRCL02jnYGJqKF11A/mvENJ/lo8K
0LS5lXF8n/bRyCPTnoeKFbwIBcbphgCLMNkHqivkzE7FFfPrm5jl4dJmSkZE+uiK
gabP7cI6rehZoo6GEmrz59C8kFlru+udZsQcsLI3Zu66GSlYHb0/Zl8JxsP7BTMt
QMIRlb43pdPC9fTQJr7T95a+xyCrz1cohtlEEWGmwc2FL9r7ZvFtPGZBl4zG5MDP
/n7xWXTlAU1zxdHIB70GSbWDVdH32zWcVta7O66UZY8pGqKbIoGZA+rHSae69KDn
Dr5sznKx3PMR/UrltnjX5l0h0PFRYm4Y3bNLkAGbFT1p7AHIB4jNK6DX5CIV4WHT
XznbSmy1TUKwhFhoksTibwmX8yp90M7cm+rBeL0xkbHHVBPxkqjgIBPcwtRhcnT4
8lXvzSdRsRF7LXaDfhT7LSMCf7SYuVJpvUGvobt40UInsBeY/e0N31900aJ+2h/V
MXMnQpRzp64HWcVS+0Fod91xv48Qbtm14WdeE1cm0X+FwAMMDSzBCTeqhK4hzHVf
4Sm4HLeMi2e7weTkPy4VLJMbwqjqO576pBAX1gxs+sDRtrkOE7sWrD4h0+iM5TG5
xs3u9tIApJBn2TqRxw8mTP4hubUTvAIS7YKCHVFs+gskf3nNp0aQy0laeHc0WIfU
7vvdl7flXXUo8wKZyA0KGqQNC3aah6T1q1wwuQgutMRNLqi+ZQACGnOcowCaMfgC
8nfJCam3LNzKBnuQHPXQTWgb98l+XKsXNJRN1UmocDc8YtJBRhxSFuycFnNaSzRc
zCCOFzwNSbde6n7TRaTUma2Mj2Gy1Vz0I0oYwyIqR28FdlX//5dFCOHqt0bBZW1n
LGPXcJb2r+fMfeZnm5sav6C+xRFW5KjXXKlzFxOoJ3M+1P6r66zZqDiXvlIC4GrX
IR7hq9LpAvTmeSWRsE/HbsMfFtbltX2/hO7rGjb+xU8G0friGK0WdKPlC8RB2H5c
xKya2dhoiIV7GmZaRcZkhWXPgX1VE1866pgoUnhSe0xFO+DJSSTeqT18koH5UxY2
aTcsY4dfO0ezAwwpmn/Y1WW6ua2iyolcsuOcYI8s81ow3VeOs6rRYK7gFN3X0b1+
yNuk8tyufUbCN5Cc3V81GfMkFdv9d2rkFJGaCaf7ar35a3sv6u/6P3i1dn8Gz24o
+l5DByHzfRgmAopdp5PHX/3YP1/U3NjApAmdhB8h5qJH3cRymzIrQrJKOR/KTJbM
bHrcmV0KbN1al9UMFbBpd5eiF2nG4rnPoM+8hHKqEgd7fx0GhElbA9ngdfiVY1mv
tkTlp8Qkt3tqY+0x/V0aFgTETwPfZkHYrwJoC8qAVJGqclVvwRtvwuGc65AvLHYr
ohU0lDXeE0WKcRMD7bKvybGOAXLFqCrPIzZ+VMxr/rc4Q6yGAt6McrVcRK04552M
WNB71KDe/KDmo2KImlg7pOGTitzFcyIZREoVvki+ZGJrEc+BBHU7CnXJ1RCPZW4P
nJ7MymABhU1aeip3N3asnqXHywGUrnWRBBGbwIzTusD+MpOSaiJ6+H79QxvnOVco
xXKsD2j+WsWG8a1rarz5Y06+cuuMAJc8svpJVKrT9nY8KB1/9MTCWTipVZyOYDQp
5Iez3Jfxc5iXb4cixK3SexCbtDe1Xegutr9JkzKX8PfewcSonK8StzxutyeLhzxG
ir+HwsKCZCxl07ntSFC2cpqzxY+9NmLoPuND/dUv2H1gdyr5TjXYyYKe8wTvJ3/K
NtcjBrZBEeKCGgY+puFrN33GCLXgphd7zmnFvfa5cpx+jfDfzBsyWwQvXdrmRpDv
yADbDe+KxxfjAnDS1Hd7BNpeBjLH8dtGXF0AWY6t9ueWquKB9Ew/nwHa01aByYZa
881JAwSiPp5M/SkSH4B6piUXSmDd+cUcCAjwPrqutx6lAXQu5W6I/3qv1EezyPPo
NhRJ0uwuKj3JJGPjFyUuVKB4tgFjiblUDTKVB4xeO4V6mV8JQ5PrAzRoMAnU6VSN
iPwRV9H37VBqGkLb/BvIz8n5na6mIm2DYYTlZWZr+NGo/m06uL4Sel0G/DFZ7W+7
7AWOUzvZWbzuXj519SLqZYJxd7I1jMCbVuQCzBvl4sPeEPwRF8Afj80u9XTckx0V
KGxDM+OUhJ5yfk9ldFE+x4KXWbnqW5uG6AZa1X9HwodXxVQVJ+qlX+F25gAmIVOx
r2ubVrtKGXW3jb9tBFWNdXRei79oj171P4MkVKXtqVcSjQzch6kGUtpa03rNWDGK
gJ2KTzpX+oztOkW6VmLVEW//KXbHFpyImpc3KlyTCbmRlMFMpYOx4L8X5/Jl4vb9
OmItGiVd77FuGGoErR/Yh52x0Mmn94DsWDMm+hQw6QoeTgFI+a7YXQFgV3fCsfWA
sRTbvENRZWsUHpFtZONAg9kwASTVl3qFWKVKaB/g1jA4+EjUawNbc9HcZeskEKpr
4UGBDPmZtTn7OhDl23sz9XHQuPj516bHWD4W3P2VZ2bhu/AN+78w8LWAyErA3EFx
pyqUDk59jsA/cAj2dZ8B73m5ZQUVudsg75nEAjpsAv3RrK8okfqTcuVu7sojJcaU
iUEqp8FypU9JLwdPcfTbeAFWznnVbk/khrc4Evtkqrp9GtL1JfdPvbOHx1NmsnpI
vAXfmR0kblzdOGffAscSHSDx7CW25TG7BjsGdU4LJcy6+fMrheav1EkApcbBMlef
EqVrgALco/RqOM8qNk6FQzCRk3LtfyDBVs0NszIr/qmdgbExpHpedzObk/ERardA
3hiEDNgAKKq7DezlMJXej3w2lVAAUmwU82GFpSu2Uv++iwlt50CMoDiMsouYPcLb
fETQ1e1uBIEB+KUo1chgyiK4jqOWMRHv4VDp1xGLPooDPe8CQ8KNlGB5SBnprui3
kXooUolKxGg6fCCbiGSDfoVkX/lvsxhDIJ03f2tHwQ7/19hzEHyHUJTPIiegfBNx
JGQN5G/4HR6TFx0mISAEurkBXC38SsCsXrnKAqXwTSGrHiRUf7jXwTQsh+vxTfy8
3gT2/U3U7Cc7zTLUXP3+2pLt5SsOZ8mcR4VKcJdAKS55SEzVVQdI40BhsEsPwWWG
OkcYLqL2MhHKtiWAfwd1cve3RC1Mc2ZFB0TcHQZ8hucZvGwls34EQjn0Y+Y+8gUv
D3hi/DnYPYW0jFTavaSVuQ59XSZAg72WLFta6cg0B9g7MsloOWq1HQUscW+Ijrw3
VIZ9U267T3JNh5BcF0KL6E9l18zKIYlcaNz9crby78bRrCtGmcqx6Jt6K/iNv14y
oCqbERnuaF7TJZ0m+x5OsZAUKOt8fFWTAT/CNFz8MW+fGZ3ki3+yVte5+/OliHgW
o6XnUdZiLeI8yHn6xJ2m6lwoalaMsb3dc8indQQGr9ImXRUyYYzc0ZX5Zb4tunc4
QLu+m+fYazc+chpBiq6mFAAR9Fjzgbk6pBrk/5OPDik+ziiIrE1Y+aEeiWmf5Uk6
lN3YQwFXxwR7pBjb/EQ8xG78AnuP/zhro+F0+TsfNRSnpjN4DCS9jR5JuZnpD2Ph
84hISKO/zZJ5qO9FIUSVlMWmfThJP5RMs/6FOJQZCzO1xvjzSoyFKBW7Nvs/zHwU
VvMTD+AleIWJ1Ayw1MgWDJqOgNOcxoDM3X/RNvn8UIFEzQOrL5sHG/KyjSWzqvCq
4ff5++gzcjgLDyIPlBHlNT38AAPU6C+KRn+0KxiQ/ycZMUvYgQcJykWI0DEuhjVh
KcUNPWSsoyNs6BDbwgRw3TDYl/mjA3EY73p85aQkaCXNBzCI36ahnQb9Ss/Azkpg
tGXp/62gp3dxrDscv8Ob1cgGx88cPrp8TbBGcM/6dt7wECCSW0HtDGGeYcWV/DV4
RMFyXT7WmxGOuQQLi3SadYaf4aoH8iouyDuAbE+d2WHxhiSag6yEGUfvnrj/fQoJ
2jkwz4oqQxIIHUPqDXtSOvcPRTqk5bEbhfDrTnrP+QkpGbq4b14c8g2VY3vLROq2
8NebjcQ5A14vVz1VuwqHFPoZcqtVy4sK+3KHuAhnNsYa3kk5f5ZZPk8neyG9Jj0w
nCjd4K1rMopu11KzdFpMfO8zNhu3ppDYSG032mKVryEYDK4wnvpldssY+/3Qv2JE
QHWGZ0sVX4PHTVSS2YB/Y6tFkuM1wPo+TehavR2PypHAAS7Ir93T48KRRz/izRBl
EiLhZv/uMsLRl/EyFD08BzAI3kfWj4KuYargyeCsiIHbeab0YPG4wYOTtRqDz95f
dtPQMRbAGKS+Dbe+pU7elomufelyCp8R8midWWvwVx7l6y4i8JeEVMCaNjpQznN9
gNLaRyeNSjHRep//0ow+CzOGZoVE/7x8j/3uodqB4r/Ou4rRT1fmVVHt9QZOMrt1
t/Cu29uTozdD8Iic+rNuNFn1otE3DIZeqC47f4GIBZmrB24FEcRON3UZoyqKhuQX
C3rIyvmHjMX2Y+F2fYMahNSjvw2hCF9fKpq01n6shSl/Oe65YtXFKET0Kzcjfjzq
cFMe9iVucNfQ5r8yLIDB5veQYm/zxLDHfZEFsAPfaptKEgkaDDKDblSzyk4bMbji
+NnuMMApSvk+C4JbLEbnPvB+AsJu2OJz0XoFr3X9dKMWU6nXWLJGYkVScllbKIOY
TyLRYRLEJVk8ukqTRyZes+VdqPdMoi5yCKvsU69uakJE5FlZPd4l0Cn31xX/63gu
oNKdu0+4Gmw6JNXnkPDJe9RV7XMiMS2jfhk5U4R2zFmaT4vNHOjMn26Xmqd8L5Dn
4SlBJzOYAHJDviTKlJEuEkxe4w+giiM0H4gLMpcP9b+BnqmZH9Uc5JSlcRwfpPAl
J85GKMmnTXFuDnVrU4LBEWH8VPs/ySO7z7dty7FRcTY/p8FzkpEMvXxoZ3sWbKWI
3S9ZYmMGt2FqK7DtAGU+P7Onb63WOaaDzZTfjNEKYSnu19lv4Vk6KvOHrwOIxgcg
lNNX3pgZv42QYvtaWoYpBRlGpxTL/AITDrcOUVOk5fnvR8TfzTzNk2LNtDIz5Xd8
0D+G7QWmsJ+XhV6qLeWApdiO9z1DGJNABq60xNNP9fHbSSe7R9QvCX4h+S4wn6vm
GMUjpTYRMn1f2dLeE+meHcP02sCGz+sEcThnHMrEsG0jum9rIC2DVgLQlGt8Ozwc
EA6uLrvzfjWHqRH6ElDFywI9PRG1qJbiZcJkAFnpiHDTx/+wJXMSJsL14eH8U3ov
//Lp5jYQnfwhkF/jZoX8Un6kUWBpNrVfQzqmKmkQJprbFf3J8mbomU9Ji0zFVCeF
t8tMqADLhSlU1682R74+2RlYoZRkW82458KapbOR8gHKmsrQld4uQZ1+MnkXS/L2
E9kDZAljlIcU/4AnJQgRlXwP8Z18Npay0HgYVC0Gaw4jC9OiITErHA2hF+q9iiCY
HJOIAvz/aY1vic5xH7xfyNDmaGBlSyBTLrA5l6eVpLd/gFJXqwQrjBX75/SCQANB
bqaSS8HloOMSHziASNXGT9tG9sl8/5Rq/LbFjdCm1DrxhwAAzIzsNVb45jZ0YWmx
DZLKjcMBRTrCqy2w8VFTI6zQCcUEsuPL2/8nJqF0jbCN4BoOpRxnQ8Ji7wBK2Ny8
G3dugQXXsmPOXhjR+75ZwTYitLq8ERje8qTkkxFkmQOSL3tCjJIhMIIOxNrGXzZ8
H4fDi9PLQxjHRPzRhNOZaTc7UyAkRZANSM7WO9WUBtZpsLtWDCRxSxdExJ1dXlAr
caUu7aiqm5tN0BT5OhbqR5pWlCro7D+zc6UaG/6aj4D1hflEx0VZwn5r7/1mYTju
ekA9juZmK+nxnnyOQGxE0BVAtEdNi4fmUVKOMJOTTFa8bbUNU7parAqoXk9MGRJx
RKyQ9+WIZn/EjTpTLYdKcory9yKWUlGlGKwTaPLIS3KHFn6BzCygNyeX//bs48tJ
5X5HoQvFj85nYvr3f0+4+tp4+itvzr/lOErWgD3iKlpTsfeCxSBmrib6x9J8J6BR
Idf99reD35vvK4+GljcQwKqYhb3ZmGEHAvjPNPcwgw367l3QFUB4XDqAYCOb00+R
5BO74cGXTFq6HRA3YMSyoWg+63OWoIgLS7JuMp508C5zMKTQsbkZ32keBDDBcpOy
XzJmMcVfYd42l2zOlrc2aEzkcmW42An6qJpSHxt1UX5iuhfwIW8TI7MlHEoufcQr
UIG/FSR0ngQjAMf3V6pFy5Gj6dpHRMcoGCK7YUdCxXu+eJJMOm7dWGEqkjhbQw0Q
3PmbPPqvgFLhDwJjTeYiWcg1LCDxJ0QxSrklgoelND61Ihmbc3e2G14zUDHGe32E
/LMAa/lkDiwAeYKvh6538cT6tpMuBjTOoZd6F8XmF9S2pn5Utl7jVTmGa/3CArqI
UvsoiRt8ymbIuvO0Vth8XBf0k9fepr+hZ9IdDxB7kW/32boyHdAYuy6UvlcMR6rM
UAO0ezZL/og38C1fcxdLZzMoTJLuCYvauNthLA1ai+fQsjusU7uiGbq49CaGhtmd
l3frSYAixrLo7mln70Ag/oJ0wTULVA8ozypEj2sV6ubDSLCWyDFC3u8n616VLCdT
SB80i0xHN5QBQVW0i8swGnZWzjNmU24NWeN9Lpw8Q9aX10emNiOv12EdJ7c8RvZn
l8peIZUH0KdevJwnv22h+PQUKWk0p/YQn421mVbCwXgrSAxWUQ3ekeHCBRFqKemd
t5rOmY+85Xqbw+NI3F9J1d2onWpaCnKlBHJuLuNmdXsxPZucQWAqejqHmDa2G+Cl
01SydDTpNrZdE4c88PcAgiiQ/8P+qf5KQWc03WAzB+q46mgiVDy80pM/3tleCzFm
25msREJWCvho8Stws6nT+UvuBoudz6e5AWdAlpo4eCXCqWuXO9cj0/auui7Ri473
iHI7wGUed2/m/L5AEr6gI4XhtOMvkXncZ5nA+xdGHbCcY2evNNLEt6bI1FdG/fde
OcBJDDEnvTEInoyRjppyIyY4+71HcQ9VknWji5hVTXu5nSrsUPx/mETEmjCjYQow
pAfcB3DQU7MsCca8MnvK4iDRfomeCoBPge6ZSxTU1blAiS2O0zBQFZg5yrm0C5vF
UBOIG/0q8duNxjQhKiRgN3fULASoxXav3oGMIGz1zyfnvpJloWvBsKDtx4SNmGYG
h100ormsHaSDqZ2rRur6J7aUVvAIFt0ywRpSKExCB/bhh3kVcxqx8vQtPMRayBhA
JEIHqMLptEA04UChv8bgOu/50MUrybGtWHKN8zU+edcarXza2bJstfvl7E9/ChSm
koLc+IX8iw3KvaJQXLJI9sow6P4gzjlDTqnm9e6+UP1Q0QFvRGHqzD5bhrtexfHz
OgLcFE9XzHKzTEDfHbLUNtXVpITIKZsZn264mGtttV8L/xVBXzS7Snsw7aLx/f44
xBPD4py4fPWpROWmaRU3AV/6sA4QHN27QT/orTA9ELWcCRQQQtmERx+iC8UQuU1X
st1gP7TPaiWVQWrtwhBBRn/joHuEE7dTnDggnb0fnVJVirdyG9y0T2Xh0HzUUWI2
6JVY5ruAR6YsUciFBUMZh7Mf6E3demR/ztnxswLxQZEcjDRh8hF1Q2m0zGqkKh5p
QyHNkssbbj/L+mTLC7QSkndnPE7bMQrfd0Ijfj2Nwm+XGXm7K8SkPnyewipSKtOE
C6uroyArE8gaYomz0wTNf/xgBpsDI3KkA25VotjCcr6GgwAG+92bmzhLQnnVkOuq
hqjyDvh+waiZpZqpBA7lDqhZLOzGMH2svpyelsE13hTAs7NHC1wViKoHekVB/AZE
PGr4azr4tkWFT5DwdbFZnv+Rj6UDpLHEx29X2j0sj/KQNZEuEnaqkvunFriVkwB+
7+6uPvXdM1MIhIwRA/Ebg0bWWX4VEUBnmuxzpZkgV77SHmkkOUXrJD5a3xDFDkou
1jery9THPCJpkxh2u2fBtxdFGbqJhmiB2T8H1cC1d1aFjZJsg92XtUBxr+okuLNB
GrB+LNN1c0ZuQVEJRMhAwduWN0imVR4lTCoSRIkR/71rl4JRUU4O7ReadVVtNCgM
bY3DsB6nPMRoOUZFqpo7i5isGaAFWkw8btFGGX5VqOZO4fsb38XONXA7ftvgdWTx
TWhNIwjr47q8BprhZXwoDsmCZR/5byaoFSs4jJUSLE5Iz0oLKJjFqjOE+VuW0xGw
WLr0pbah7DCD4iN4vZ1ybGs2ToX5KXB8PaTgX+/ItxIvNU0UmXvLHk5Zx2OaQUdS
ATAjHqMKEp07yLHZl/FZwhOfv3erY7GBVGLQu/PgIcwnzwcVTe9ia/PX9DZ47yCk
bv6v5eBsJflHZRAWWKg/2BAMZQYcabk9IFh/bN6JThAZ67EACiSIyDOUGpDwBBSK
CTCqWsiZGlHBQTSYdx2PNjMUwtt6T/qOYWMuhkPQSKed2dHz9g8FjvVJqVtctxFK
oMnSwbTEkqMdNb9hZ/r6FknGd3du4975fhyO3bnWUAm3mNq75QY7DQW7/Dl+mh3l
w2V39WqYGLkH3olntY4AqbhbAU/prCJP0KkUxyJ5nO2IFsIxsYLNKbp5vkHByEEj
nSEj2oh2bGT90Cdi3CvEzToci4SlrqT42C0sW74NWWKLgs9zHX1IDsdBnU/P4f2v
4XrsAZlVBoOQTGHKaBOn64NR24Kth0g96N8jmsqinrTspbnr6AGzK45BgwFIbDwv
1adP/B4DQzQDux1khTRoC5r/qNBFiluWpubZdCgsOf2w9n2QTRxTnXQFFfGDVoI7
mXbyjfXteOb9Wd26LC9TgObJVLVmGJl1a/DkdWFk1MgmKCu4yMT2qg+AXOhr9Oc9
mUj/GJz18fuzg/MFMjTQ8xM3LV+dYwIhMQ20MjJpzB5G/khVsUXmIELoKF/p9AJo
yWFOGnYnEPK713eIh6bdar7zkZOfsWAxiP971A8s4K6P7dVp1hvkSoU0aR+WKUZp
sd40xBRSYowCFkla0Al++6kFz2IWvw91mAMZjKSYZKjTWnBU1c61/tV+L8KNWyKH
sRtcBUODHhjuEb/FKojP3tuuk8K7ca6O2Ldrhri8CNlFWUFxyqRrAVGZ4jcNHKq3
98g4LQpixSdryzZIdSbofEgDFKRNkqNpPiTQ3HGdYnlkSMYERszOzFpyKaP/gQJx
Rh3PITHLqqbWQHJ7s52+g7nJgYUU+qRGhNixkEKHuLmuzxYCtFrwh2rBCvDw9hLS
+Mol77Fo2PdywMipbHc9hte2VtnHfu57LQLL0JcXfut2FJTBCKWBO8I91vfWwi/9
7lyn/LIPBOagQaU2BmbCPAQ5GwItQTHOyHTIW1dW8hZns4KRjcznWk1M3yE+IIOV
NbWUzRuNVPIWEuisqI0LPmRAbnqVyMZ1x9s19GATCT6veP2fCSS2mvbhVh0hPBn3
8Sq7ATGLRmHiycPUlMJvA1n5gtK4s0DQivHtk4nzN7q5sDGCmeuOV7UnxOw+QP6i
NUJ/RB9aM5iRv7i7ehj2y+Jdu8oMIIkoYDfkcR9mb8XysjY2wuybRY1TOez17aKj
nYKASC1C+HsG2bMDQviKwAIJz4uG+FY16v9urankz3s0kWbO9LPrSkWO8lvk+2Gj
bh3ycyKrNIShPYZ6dCivBwi6RLolzBhN6F+K6wM96n119JNlH1V0UuHjGPv4Paxv
iOQ2BICspqkABn1iV/N06I/2fOrCMJSYCXhRNYWH1OUslk3072BkWzdAzB84Yh4Z
MfEe/J8weghGF48me4EmMoyv7ggiXDxXX1ESQ+a7y6pZF2fQH9t9KXwUxrNC5fE6
qhoOdAABH2AOJLwPJVWFemxu/NQnhzANLGUqNAc7svyqXqEw0Gn1paIZ9NvCRNAD
jVoTHyXdAvnMc6BqlHPKHvHQ8vOPL9MosW+SVkHXwCEZbxp1Jfzp4Q92fpI4FxvK
L7itSWvbDxt2WlmlRiyiI4VlPOjb3eLvnDvlHm4N7EIwsWlGDWu0WYgby0GyU2IV
G+EtATVNded36u5oL31BMB0J2UE8+IaScVm6oGTDi9DgEmXmEfediMcckke0eETP
C2Y37wVBYEbNjhqhutbVR/ry6TEBkej2nVDvhW7PA3ZqLPOtvUFucf4aY5VaMyjR
VzVBWRuDmidx1UPx6QOykkpEY7CxABGzyEcmllXNPDlYyvygW3BWjuoqzQnl0NSj
9NKX841umIfcNJL0mNZLAMKFxU0WMQmKyzREPSj1RIUVfttVB2dmp8o9B9Alzgm6
KLAFEEEsrd3wbT7zZBCvHWTrKiNNdorv6fl7qjXTT0DVsHoe2cq/Cq9+givLFHzT
uauCbFjbtQPGVTU5DN431HR5StwzmbNYe5LXHvQGkDf96steQdA1fbX5JpG6csAY
szNG+4q1uq1Rjk3jQwSAbKzNz4fCRaB4K7/iwcBwltWTmt9M/jWqsfMwreOXQ+wd
z2fZecOKktGk2JxLGxe2hP/X0cfrUwi+MDOVRSJT701q8Zmj13+n68ZhDc/eD8ZA
jCCWkA5DnUDkWq0mw53hg90QwFm1KtejWrJoNMtyii4eCZgH0+22rqnwMti4PXtx
nTsSakF0eDFHWOp9Ix5huj6Z+jeC7jDYP+uVgRmWgvTKOytYS6GoXdNackqYmd/N
/c4uCoDXwN+tJc/wgyBjSIqGn3nl9TzR114kgxcW1sazm9unljdhL+TwGPnKwiwv
FrJMkq9xOH2cldWLQodxJGCYqfq5E7M4fJkohErKn8aYW/jiRdCVfgWyWBGcB4QA
nV92D86L/GPZv0q0MNmWTLeh52QANhHKuuuqBuKA4ECkTkzo5ttLTldeNrml9ggm
DitGq3opTpR2xWK+QnEaorHxtFdNwcQU8h2oJL+XBfxtcsafcwOEL5VKQV/dcUFD
DrM7EiRX/Db4ZfLQlmQ+fq6EFs1C/LIV9qTnen7+ndnD0N0c0lL7LMbFvKxaAp02
1NahTgtg225hjHhg6ET/o6Nhbw3KMp7hIsmwM/n6FS1qwyfDQT3u0FDJDt3kJ4B+
hFgiVLvQUFSEU42KzQFawQCo3AXAnwivssz5atWiWS1ZI/n7Uh5/C+BnUK05i26Z
0dVDwZl0/XinJcGxrk6BdDMrL1a8WhJCCVvhYSnxbAvJt53bTU9seftvc2HX1k+o
AGn9zy3PnA5r5uM6mCmIHHTFgTbIiKKPtoL7OuuWBUfZlR0EU+44lncnExkS231s
I1vKdg+rzqh3dxUYvWKkziYavpDCqjJoUnsDlITEfGZRBI59kGv94B44rD7ksZrz
UoFS/nbBNgGaGiKSTgFNpIBmYVHKbJEBVckEC4wKRfcqkQ/+nRQLTddbfBpcUr5j
AkAZHDYWJnXTabdcEy+WIafa72UTP6fsl7wzBsSyKPvCzqut6DsxiYYC24egiRkM
y2g8cKHmpO2pWBWzpKg7jEfZWb5rAjs0mak7gHvCz95/lgJGw5klk3p2VWjNQBWQ
9u4Zs7f3oyHmRTwM5ZrnrOXH5o3whFHcGVDymBjZGgxbMzXGlwtuRxArreeJzaEK
hjGNEwLT51wXrdT9PEBo6uNiegY2btHwZhs2qH4YGYuE13gI59Y2dBDh3jajPzNk
mbAnuXu/ociA8IeoaBw4lxW8g8NKQlf/ZVoh23heAFSujIA0H1XcoPr/uemHGuyv
KdL/TNkAcNEdLqrCraWSMsx5bHcPkSpk+3FMGIDLZA+ptDPEF9jWOAtvuB2RG6PZ
givDfHXlOARbDLZBj7sEE2VKXH/yW0THrGeuB7SZZrAC10ShatjKDMXI9gXgRb24
WH67rTZkRb5ZKb/jkOE3k1IZ3JH6tmS2nqP10Clb8SaTQZigpaJnwH0AzQ2ZFzWC
K2TGr5RmrrAe/GNf7FroNrCORM8fG59qeViared9fAbd76fYZ7SrtFbX20cTmk61
l63Ko6COsoTxwOpoQ7rJbjF/Jny4Uvmaz9Z890WjlRwPg/qmsRSkLIVYw0Dy8Nym
giAEx6W21pzza7N/oNto1SjzUX3k9vfW9PV6b6mR3q32HnHePg8VtPfiQrHxwL6U
IsJkzyENfpC39D7o7dxUFiG3x8dRuKfT6WS9Lgy783Y2gVMnHxigTh0Ak89XBJDb
TpTucEBYEhimNAZ5vrATyXj/aaMzkdpRtdGnNtKcKlV3Rn+JAXyHNYmBbHGTzBPF
CM+E/SS079/b70y5jr0oUNaBLKA4uYlrr8x3YJG2p8oZkV8QbMhA7xWcEges6s5G
LmwVNRMj0tEVK8f21J84sfX5Go/RD5Xwq0xKsKwEyHg2KInfMAtc9ldlNBoLmTTO
PstIVlghT1omkUT3DnN9AOCf0tXFi4a4/UvasM5i1GtNpQ6jfI91JRmH/UMJrTV1
aW7+2BtD8jIwo0fW7AAAybYEjgE9OGPoOz8FtnHaoQQzR+UlWNRa+l60rkGbkpYr
rV+dmFQe6el8APx+qrOlE2mpFPLP+JXIjRmo7fiHQjTUgS20BEGUd5EKcWOnnVN2
dj2ty+oFRcjSf9TpGIlGDQPdKqDwnBVl5qDXb2mzUJm7gLzbcrIleZSSpv1mMHdp
6oCoMA9NBimoFK6Ex2ds6tfSHpFvZzvGe0x80p74mJDTo7ZHGQ1bo0a5/1/kdU7D
reYlypzdQOs4NHI8v6Z26y9gkd24qJqcMT58/n9tjfY37cXqGk1xYwmA5OPv9TpF
GCw/l9Fz8/9XdTUir6kycpJ4OoLTNv9EbFZS16cpSFBIzxNHwTilbsbqAdjLeYBF
rzh5QKwcyNPSUgjjMUYXNux17jugNOx4EYPAPzp8WRY4Jz2k9M3DEb+XsBnR1f+v
dLepQoTdWlyaBWhsSnCiRNX2prZpcZM63Y3CpquHVIqetDX1fWKSFzkfQKHSMwVG
yiHcPZG6OJ08EQ9jq2LE+Cft34G7CNGZfMB8evp4HSXdePu8v0bsNquzetvE561B
WzotW7TUlUmlmkjEs9dB2APsJjsi9YpcQI2QdS1RlLZhrcv6Hugd+IJnCoLlEIf6
cFRKHZcU0TzfaS0QOHWkS94vboBXeWhBaoR2q0OYma/d/nm6RXZ11pddo0nBDqQF
DpTf5HriOUx5UHsg/vPoGgs9g9+4iP/xNDxRAvey+HoOFtLzyHYyFIL5ZG8L1+1S
8kx2wDmS2U8xhbplSYGWiAHWAzhmtKBNFoS3szNH2Xw5mTVdFq3teSKym811hjPF
0q2+7jd8yfmF9Q8aeYhxP4uCheJwJtwQZpEMQebkQS1BKz9a7608BPoJZdLb7Z0c
ZLBg9xp0h+1EmE8+8K6YYOM5HyL7rYSMx73C6qLVNeQatJt9xzNIIs8kzQgglzhg
nOwCN0Q6VdZR+McUk+An7i1oavoCJHxumbi+hFNH85xZIed5JhnSY+QexuAUHJ8S
aGGhT/WpJpjm4NzjYoGf5Ksv+PqhzcOF9qqEVSI7HxUefGafKnqT9d3wosgWU5JQ
StCyVkUwMemsePfoFQ0qQIQBbYM6O94af6GzSD89HrZJcw5+0CZAFbSHEqAkoDMd
s+GxDRVwOx2Zjw8K3wZuKLXWzGZREGFJGCaMWiJW7dSUiH2q0UDi75Qi756DOB4v
k8JQbhn9yIE69X6oK9PhvsvXoGs6+y6nFh/jD9aqu4mpD1un6H+JEf122mgkNoQV
etToiBCWCq4OtbXKSEoAgpZDnAAZkZHEqQg2qessOAhp6esxBOIUOPmtDcAHoLMg
Hs0wI31hLpeW1W2hu1CZWUu4uG/pTpAJRiUbF883oYUSwjNcDnFYv5/5H0mqAhni
JuFZCygT19f3V5a2lskYM9BXHP0IXE5ZzbgOoZ2y+5g4ERWgbl4Fz/wVgE/5LcyE
ZEzgtjik0VmufGYkWkglTG/0WPkU58hfW1bqSY5pjk9q8qdfEld37M7Q5WALUtwO
QplQ9qRqu3v+uuvclu6Hk+1iZuNz9QQ0YK7KxGnfO7acMDbP7DhkABc8skNREdI1
xji15YZhePzSYliyMMqJjvl673Nk0GISd/SXP5c90kx0y6o1hxLxYAeecRaptKah
e0EdMvwAzR/kZchGH1NM2HrBmS7Hmw03NVSAgOQNolz4/zwVHevQ82/Ibabk9tr/
kyKKd2Ku/JEntLZ9idBI6rt5DmoKXrlTUO76xWxJmFWBq371bFUQGc4zqiC23e8L
6DF5ryyuOuss2HUnRSknpvb1aq0M3RCf/HvHgP5ella/PUhyOr/TMKas05ZiZJv3
ZLHBoJ3bUJZ8jro7yN0e2yMcEKX0C6JQRgokuF6Hf92o72Z0KBel21UTsqQczxke
VWj4NfUL6R/tqrHga9QhTWaaJsquDzIZH4WMz2FOj77X1LJryaTrYhgqBWulw7Qz
xft4tJaVFckr0QSFKgJ8IxeR3HFOf7RoZWr6TFGXhPzomf1SVmZ7v2UZj+a/XzDD
zTnoWqa8xiC9JoM/XXZbbn8QV9dFcPK6toI8WpgDSMSQRcEBB6gcgdGm6tAj7XCF
2jxXs3L3COA9/WRfAShgjASSHiO+wsJcaOUlwxLWJJBAmVuKvQP43QEJwrR1BBF0
27V+Sa6klIdwM0F5gWcfI212aCqEWFCKPu/iYiZbmMJeSIX9OfhOM7G3kgTrTI4m
9xTDq2GVn//to7I8LbQqILGaLzDtLLu0V5ATpxaS2IveAE1+nbvzjqOxPFrbWE8x
b5ElPRamMKrGxOqblKSjEkyPyO15uaMdqMnsW/oDro4nBVQP00ivHuldpMnx6V1S
NLK/2XPF9nWpQwaRMN9zTr5ZJwbUnqcI3jlLp5ObV3NZIxbmWZJ2Sr7pBMcxAMlD
vOQq6bkOebA8wJe2wBLYWQSMzxQunHTKwIBXOjszHOkhyi3jeeefP+qCLmTPX6b/
eZyIJjcC6Oi1pOc4w3afSme3IuxTxrlt/dq5BbMalf+6Qn7QSxLSUlIvVa/Uel9C
+hJo7wyLU86xM2R/mbsZMJdCbNleQ4rN15/WLEsi1na86Krw1u25lavl8QBv1Khr
XLIQF91sBW+HG5thtBDg5jPljCeko4f83TQJGjPbAlxdh8R4Iz4iYgW8PmTZYrP7
JJkDzMbQyR86h9OY1cI3mQxlUoDvoIganrRkhtzL6hL8RprXlzgH6BU3ukuNadOa
EZyJjB6a7/XKwi+X766TDD+LvQGwCJjv5cLviP1NO8jWEtoOHXM1P23RLxe9ZOIA
ZU+eqUsT5Q/qKQpFKHJxUnlW6P2OIR671IEKCuOz5pgbk71uAdQWL9K+/zY2ERGW
xvgrEtm2kqYly4QFKAKQqOEjmTjJCkkci9xp75x4SBrKPDDcJJGbD9BEcgAGzSOg
jUZzoEhbJCfDcSW/JPBW2x5oU9F0PvosRyUsUUQZcievQr1FSNjk9QwMvEuo/Hbz
ZBUCQjtn53GEsTtKXlXO41FpcALcAHf7XFi/YLcNut6fB3M4Y2FWKFisCAvNTAFU
oSZ1jbqjeRRXLtqB+6TnZfI2sK5d5fngX6qXbdWYPkBUmSmQ7ahRKmY+ZYMKOC33
hlviFCBGJdx39cTE/JV85gSywLtKaSl7JqvOvkdENgptcCZr08HVF2LTAqovxKTt
VpO3h04DrZ5m8XiMmknO3ylJzRysAcQ+LrXMmFXo29rUVVNIFcQIFWcr0UDE0vQk
2UfFajv+LGcWYMp/GSUT7a3cqgxgMkhStSu+h4Xmzhwj05SEZ9QcIJQ/6A+s4tvA
iZ00AQpl0B6rHao98hzsM738Lpf4FN6DE25l6tMIWW+I4kVZrH/9YLpnho4brW1x
lV0tNzS1PjkGi5ks1qeG2RyLh7bJBunBQX/C39gUmGGTSdvPRNi+X4AhlG27BM0B
EGJfyoBAE90G5QQoBm3KZeMPRb3/nIOTUGDN+ghReLNNnfr8aW3C62K66whhio2N
g0yeHaT+DjMzdNVBf9GzrI3YSh4Jbg0RbhFmc595GOB8F0+tRN7sbiWYqbFkv3Dh
i+oFSNHG0vgp5e9/U1T4vrXW13JtZ3dvbhu+y3R5DuOmZOtCUK15P8/X9xV7jDCm
irjIk+htzQPs18Tkhm5CgL3ydUgsInWaZoayV4jS5Do6igRqDsaREd4RffWMCXIa
7/sLikYUMNZcxuxs8/MO47jFo45HrkICI0rAxA7w3QwpziRwgfwyfaPH86BmWWSW
MDgrBMXleI3j8bPJ+Di34+9oci4YgwN21UAEUtSyAAeLy5/i811KJuJBxjD6K+Dh
GVRZtoNNORbKfr9mMrLZ1eRkTJqnE5I3goduMYmd6iw7PhMchne7ieahc8g5ihZr
C1V9O5Kh/wdsgLPDyxNRj7YcsEJorYPR0/bs+ERQ8VSMXa8l4yAl6Nv0+YPdGBkb
83SNH/dAbt1kliXvJF9atsG26jwbJ/XfB+ihf1P78pfHiDd42znuZ9vICUzQmfJN
AK9fL/H+nuuT3QEDOMw7sdRa7K66b4F1bsfqNlsEG3UdiRHzSTPU/bXQggPStEGi
MhypheCrZNQh2rVOi7cSRkcvc5Gn0vUIM5nY3GyX5NAC7cgHlUIm0PF24sUS6koT
3/rwtUGezH7LUav1wMjndyRlMtkStNplbyH3MirS3e6U/3GMJlH0sw4fUMs68Hws
74ZofolRoz1CEezudGJhyED4G6klZyMfn8mEhyUUVZ8eR2xlkNNqiBEIIuilA9cM
iB+iGKU8BDa8GG7QJQl65havl/vmuwR010J0pjEgC0MhRAAfDfWjrxJipY8q1EN7
3G6zLLrGoXBnDkwMFJCtFRjSLv/HVfXBQqf+yl6nuMsWYByNvYuiQ7eCHLISsT07
xuzmGN1iizuu97TGJMCedH5rjT4Kx5kkmqHFFHY3aaxLGGyiPcTBWmoL7vG99Bai
eB0JMkFAO3lOR1N/rWMOLlekN7YUEwEVyt9LTpj5YZ7rf5R4cgpdyNY+GmGuIgtS
UftmZ9dz1g9VfqaDQtasEHCrxCaG5iDZ6vt6dWuwDmkwTiENiv+mnuCvxqKpzuMh
00rejZupfL8QyA6T9DWpb9qS4oBwUqftDF7WGUl4WTu/oMrVlymf0PgL/74jmw7t
eWe6IR5qnfyF75qze1XkhezkJTYfYAa4c+kH9SEsE4uDs/p4xSbc74N9txsH2QRS
HMT9wO5SU46eeiiHjg0okTeaOhvmewCtDuA8BdiU64iozR117h6D2xK2l0AmGefK
4PjESbUWYmg/InSzsR0CTLPMJQCZKL7oBLcbKS9gUhHdel088PrdcWdT/CLM2q/E
h8BQUFEXjyktSNkB38OfxSPusXnpS9sG03y/ybPz8CHVHKBIc5TEwgtNdimQ7+8+
nDsSfD+mpTkNvZXbjaa3lc+pix2yaxVLixF6FR0L6wxkvlnlU4K+O2qkTjrTZ8VL
Yx+ELubBijh4tZ0zhX3AjOUK1CZb6MGiQK0vn/A7wyVpj9h1tcD+a42zOGEZjfhX
E8XvWuS5tajc3q4l2dFPvrG1yXjoqWuELdw1dK0rAnU1ibUN5vKPKHzBq7O5+wdJ
HKx0cI0ce0qTFsyqSfHg46unwMHloC8CN/Ej4dpgTX6fFpGM+hCZn0ezs3Hn0cPQ
iaQm3nIi7YmoMuUMTmKCqgJhw9WA7/Xis4iHSNJStpU1XG3Z8dmZ3O0tNHF9UKqY
wOE2GxVtvoZEUopyfmjg2xPwuOPY6nJ9eCGBpr0R418SeRuM7fbOXuKtKnvGpnVd
6uPJL5cH7UYX26tyiDZJa0RK0eRoQveSw4F9jBov/kZ3nezhnwYjq9qksM6BV/vL
FAFRwqN7yGQZcer5NVXnF2BdfhqRMzov/zjbjc1F70BGMwTlRFcCBd4yxcEJfnUr
iIGkkCe1SldCCsiFYYqu8A630LgRLHyzs7n3H+QUgKI0zKpDC4boYBVTdEOZl7Xb
Aj6A+eV1npNNRNyPN9ovVE1BOrjHRDpzJoU4tfSrMh933OyciGIbdAxnH15htNUh
UE/8/0xZdfs+v7pYYY+ru9F4K4zsNscEhc2/xRIuHTrwdpAQTIjoWIwHoQGXET9l
1nj2a5UEjG12jfQB+0dMbamMltnonOkyvQ8U/WK/um8FS5GiZpWyWDxmCS/fuUHc
rd/ZYFcBguN/2wrTbcgsVmSVDvHLYdLziRx4IdK2HQkbGcw/1u71OJmtUOJ91YSZ
nTgd0fSnyDXEoQjXYyW7LqN/djZLq6wPjFcjXuKo0EcoArHuFvUwC/uX4krPmJH0
Ufw47ry4uRu1BtyLdoDhMcUD2TPRWbJmwrUvQbRzlaMCmwmZioB+gxBxndawJCfG
ZjsH2rYwZepN8gO6fzUrd7NMX+3dRRAWWbnbhvia0RsWw9MvrZA7XXW9dUEbqJnx
zJXJnWuNku3CUqojCROTsFo7TmjGooW/kJ9azABWCTy1f1oWUe3d17acOTGeYrJx
PlNCcj+wbbyoT1O2/JFaTdg9Pi12wb7mBAwc92Hd8fsF+1VDb/aFMz6hV6eqntxw
Cgi6ohvWljVCmyy7lvpSOTWv3uFRW0+I1YSDFiHVXBS/GIC7Uy9XwyFUQZsrCyNS
0LH7QW2fSRkgXHF8AVlBwh4qjVWNnwzD3oGcK3NQSUUGDugCbKq4NaNXfJJyihzB
HBbIuuYENGxmNwscWT4pNhpo3JJNkTORumciusTGtU9wm9dQ5adSBZ82E1+0homf
YuxqGxs8X75Y4OOEP8eHsKkld5PAlzKh9mQ+nxz/nONUCCeJ5A2tplT4oE5njSq3
ZQ2zXKMVLsxsvoyj6rD/xzVRD79Vc76pvtmHMQZpPNPOQi1WlPplNjVhSe5a0KTj
itGjSfeOxtoxuQNKEJRdzylHkUZNNovkNawzF1D4cqRQwF9qWTqkZLLDjoZIqHEu
D6DVl0uViAXKgBSlNKrl8ah6z0Pr6HXFBG0nEYZWr4MsZdttsUif+TL+WonXCuPX
HlxPY0v1wlILuXnwcKJVpJfjb3RVs2kFWAiNqX8ahKwBhPKP/SqmGGIOSWZHphpd
KRA49fFcWRx+rhJQYFHnW27B+aENoVNgTJi/WgnhnJ7PXKoA/ZgKI+B3GaWqvvKz
547ZhSqfyqeOqpP0JXOjAFFbHirOMgzkhTx3/kfhN7uxe8s7U66hGCXhXxaVETNM
GVGM5RrwpnAD3ltikX4wfyCTJ846LTp8DnSASD5gZnKTdIDkbI2pps8W43DKcIQ9
Pm5nHfCo55eZIu4/Rbv6tJuGt9XfJrbHECEb41Esw9g/P1xEHqJ/uETBFoLL476z
IhMmKOb3+7Jr4HI4iEzAWw4vWuXhFP/7r8fnIJ9V9URzaw5se77uMSco5cwxShFX
ot1bPaY8GEri6i9NkD1sGmWk0Vkfqwd/y6QUawSzDOcjxnMtstFabSV0edbdBJDG
IHZYBX0cwlchtheQwT1/uz36rIVPljS3QO9kEbbrab4cLt1Hkx6gWlwlUZERMfos
71Q2ZSLk7rSF/04l0NkMDBM7Uko4jRYVGW4v3nfRqfh+agHIdn7Mvktv8gxHos71
x/TATyPX47Tgdw7ZNbY5zq3DymbVrU1Ak41bkqfxjDGo6Q2l7vDUkWeERdN7gMr2
GWbGi7XztL+g9mboouwHpsJqhiBxoanQhJKnMtr9P2aDtGrR/tsUlTsD01fHj1aA
Efc9D3maVO5bQ+A4+YDlM7E6/VEWah9iqQJEKSpeoocOpR3sjqF48bIUWaKEVzxa
8vPryESttQbBpCorbbuixikZLNzh8+VpJnF8DZ6TpeAATPgyCfEc3Zv4ieDzx+04
bqXgdbBtif7PXWDrjdiYCYUlh2VuwFZ2PY/744i4N8z42xPqZxjb0Y1FfnXKwO+c
ifaQtHC5ng7jULMkQZJj0o7xOOeoN/2hzaZiqItG+tEx4/+0LIS77gL1gagL2laU
UZDqe9Gm7BcdUoLXUrvV5E7ohJH88I/LAxrvvzaMuMhslBu3OYGCKh5h7Uu0uTm0
BVgXWOqqlCHgPWSzFl3SPnh/gpcR6Q6zZZzZiSe+vsuvMyjjN8vNpD/VXOnx9Z/O
8St0JmSLJH7BTjmVHw1fQCmxa+m9oVVTuTM9Ur8OeTcHJHjURc1dxA1KkbauD3Pl
VJOGDdSclEmBFaG8JuOR2MvCn+IXxbVJACijbhxsdQvzr1TMkw5iD2b4ixQzXbmY
MnPKiGe1Q0jRiSdCt2jmPT9qeFLVSme/74ys6yTnpphVJaq0DCi5zkQ6zC2Mew4T
p4Uv/7hpCIho/kSDCZ85WekWNNcwOm7lGPO2YcKAJZ2GR/BWqmwC6RVQww9iNfb5
HIVKHml8yJ82dda+zcDT+RDjA4fxP40swhoFJCDd9aUHIlBh+pvqY0Gu6wtZfEB8
8MsaJXcCisZtl3G2RIIpVq7H5kg/Dog29m31NLlO2vG+mlDhfXhYKK8GuiVRPmH+
UHLGEPBiuhEz9Rp1aRm9NS9i1NH2Y/u+72Gga4XDiZR0Z8+Jo55vGVqr+wLIJWvq
PgF/ZyiwMsiH6Axs2qQXdoO2TCSRgdO2l+swBO+pdLhTtZk5T/wirULSe2Sonig/
OE82W5wT1rheu5GDMIBPid5VIslJgoTaGWPkL5Vp0Cgo47mxeHBO+YyQhjW1J4EC
ei60umapO66u+HL2UPq82aqjYIFjywpiVvKvM2nhXpZCPSXLsCaA/yV9lkNbfdxS
YU2B3zJNZbeQUXvBraPTKXClbfq2yqG9cPXncylTYl4TfcfepPOEybbjbCKWMcd1
fHu7t5dp/gdrUEqf31ZEjl2+/QQDt+GfZll2g5wfNGoJfUXioGCv/fqnboDBK088
csIGspuGG6nl9aU8i87XQ/9q8pJExD9Z80jWearCIQo+zc+GsKPLZx4R94LA+WbN
2Ysd+DUNHKWvyHPLrEV+0w9iwnkrAYSN1xIjq6PZnjbQOiFxuSFls8d+vVLLCPZb
obHEdxl7kzoCMGrvO8m4V43cN5+u4Qyw1OAupKFRVEug4lOmDpzfMUXkLORQY5dI
TDOp2fZnDJVa+sqzAK4d6MqG+wgXthnFopLkmYL3xw5RmEQm2pjaETCqj3rngWcR
9GCqKjgfKZWlUcumjRXnHXl/uVU0Esj0bKlVnMNRlMSbyJgtDeg/AwMVMxdfKvQg
AhFZb5Qju8wGuXof4JoDH3EP1vz8gU8FQ1tWfNYL08Dur/ZOxtl1Px3uBn/Ai5Zi
WcNGN3kPP3WorbahLYD764rHvKgGPi+OqTiSS450y7P79U+vR9i6nBCIa7+PRdWI
g/K/+p0cuHFT4vK9to9xWqRdRCGT/ujyYuwW8LEdUxaOmVh0nzxsZpgrtYHd0/ry
ntcBVUhB1yJybIY9ZUJmpLiMUaThkYkmUO1kN1o07sf58/qbCDuK6rFqEjIzoxEe
RsODuxW84ziTT+FenFbtAM/gLunvYNAFEA43jJA0iZyka16mdk9hDfbUOarZr9po
Uui49Ymd1MngsxSyyOHl/PCroPQ8RURFDGTdxtOJGR22LIWz6FBpHhFhNbC2Penn
21Wo1Of5aNqeQW/VZEU3v9kymfODud/6IfrzS477N7Eo2pFQcR6JrAO9YC+BZ2id
gGMXl2Y8/FtGzJyHARvRqbtXBEdyGLEu+JE9yqDfKkc/oFdXMsUR0gazpveYtNMH
/2Ha+ldtApTsPLOfSYR3rqTGcyXI8RHYtR7MXs6YFXZ1e1ZsUT5E/hJ2Ieh30h5s
5PkxAPQDbrwMDL+FSzY/kzkt/8UnoTxIRckzS0UdmLJFNDI8poXmf4Z0DpmUeaLp
nKOTd0sLF+SGBxBd1TWwz4zfVgXsLhK3THZfb941EXG+80ujWXkSy39qnCfPiTTS
Od2+bzTwitvnbiymogjR0akq0XK5FpweYW9X0VeywMXtq0m3tTCB7N4xxx4/b3ny
/VePvqQQcH2Vl3Jr7WW5gFHduMejDF/8C8P3cWlYWDGeQDk3WvNVXkvUC4C5bH5U
4wVMxezQOBXvfyEhXidPziaikDFEQgOrT2BF/vpwjghXfvKAIiKdGtPsnHTxvtug
U0Be/kb2C7g/KUel+PWVFce0gAhVWCfzEGbheGlpRG+6K11yW0AiBmUnVRYc2qin
+/LiVl3LG4NpwPoZkmxAYDBAVcO4ynhJCSq8ziIXlDsiDEqW9Dj3JcrzYIKfB5yJ
jrWMVCSXUECTX4AQzmKfr8Dk4ru2tUURQFK240rTwSI+sFBFg2H3Zy5lN7FvpATR
kGasn3skS6qBPdO/yM88JY+7ya00OBwyHt1CNoDxqUNdX/NcgA90md6+d1KACVzp
EU/dZH0HrLTgT4/AOIPNfUW+8PtuNeYPAq19pEq85QwAioSPdri0SPgVLy1d5D0e
71Ej+nZOMUC5pvn85zcnnppSISQ68ptd8A/tw44zCBjGBO5OHs4Chmix22KvsCFC
68fzqq0/U5le5xV5b0g3/Vs1zM9carmUpA+Uu0Vavz4LGfL9DwoP1VqOZM0heZJM
IvjpoAGhLE4NhgmkErF/mWYZuq9tQd1mdyWnis+yVVc0Od8jo01ikbCrVoVkhMs2
XTv6Z8hq1h2JxxSRBv04GP4wjW7mWmjwzqhALHju68VJYkUM/F/pPNMkeFpJjQKE
NwQdGITR0JivcUmeum6SxGUZsToIUv++elIYxI9mQ5AkCnHVo3paDOtWsRG4GfxH
J/EilRpUMYXHC5/NTVfyCEo3l+qM1yWQvt9K+QzxR7gqhT3xubIa3KHRiX0k56fm
VYcq4iUMmSJoaRs1toodNZnGAf8VYZViNe5ZaHejOX8oNkoHxUe4d8Yj6jieQowu
joTrpPwce3k+RylG+ogxk3X3y83y2V+MTypMl+m7GzBkoK+oo2kgZJs3bdy2L8pW
DqJFVO06XWixy3Z+EHiPL/NW+Aj5GNrR4E4VbLeRY2LBVEQh5zxpksOj4atdzfYg
kxbZqzIOU1doKoUglSNYq8GjrfcdpMNwKLJ68D+IoyfJWLUhXpvfA6SNdyhB/pOX
6MJ2/EbeRpF8XAAQKRPHlhNZGOdYcQbkAOxmhqMJYff6y8RYV9g2ayl6EOnbVPdq
SaF2khTsVPl2ng49/s0Pl79cqegL5WDNTkHs7iPtsm8KdW3cbx/WbbYxS+O4kEHT
0FvEAzV3KfGLzKTDmM/ZZQV52WHjz9D8K8D91sxf9p5aGt5zYFkddEC1/xvPku4X
vXEcAZa7H77YEujQfiD+k8nC6nhtGft1FfktvrCeqGyL2QfXAWd9HeTtaAqY5wyI
Py0ERTksWB6XaFUpdA5IVxLFp7BX2oJIJwmnL9RnK+FYEVo7YNx++qs/gBpCAyxh
a/TSrv6x3DD+eJ2lwmpOJePccgssOYLmVT+Lh+8zGC4vHlqBj+jsQlQW7ddOjeQV
NYCx/IaA3cSuyeLxlR0sfpS9vLTW+HzQCoPnSmBISSAukNFtVx14a9wwJHkxkK6V
YyHesKhhiJaGQny4ybAbFJZRDAaKjXUjz4kBQLrTYhUKN7WtYhVvxR25t+TDlFyk
cMXhMvktxgZi4IGrpvQdY2/cUZ28+tcrN+3XWPdWL80i1FonDKnArJWNDuCEiyhE
ebqBqBnSOCR2+2L6mj6piavDMMpGAUToL0uuriz7nzP403QYJrodAGYk/T5cMn6g
pSXa2LbkHJpHcvK/6v33BiH/q2tXiXsSiBeM/6cBv3xAIHKMLfUYi2jef402BZou
/Qb+8hu1jBRMxBOLu/SbpyUC5Dx48ZyZFFh6/nqX6fIRaQYMkW0UgZZicfidTtDm
YIYGMFqZZkpH6fZ+OBjv7Jr0V4ZM6lqYWQY38nsGcM0x/pJIFS/SlbM3a57oQ/SS
cSlY17cIVbL9wTo3vYcdU+Zuy7gNNfwFKxYUJfYjt1qhW+iO1iJYVX2kaCvYOpNd
auNCJo/aGTJi9YFA8Ms0x8q+zf0T6VmQhOle7BDnf6/ozuYqb2Z0i+i+h5pprVuy
ryV27oNOBp4DKDpLJN2Kk9RT+U812pmAHxeAKa/p+gU0UML8gzVPxea5ZqhVtBFD
Uq40d9NP/xIer62/U5uKuofqiO7nLqev73csjBzjA+DZ5pNZZpY3lqM2nfnTw1S5
Hg2lnn+EvfhjpvkjUJsr2kyWnK2i3CCxxKimxxyoiaXTxutkGv0bzUW2QO4jRjUP
cLekHrnN6DdWgurwVKA/dt/20zdIC9HqEp3YCSSyO2cbIxgNG9nAvtSzDA3D/dTM
MdQjj1rwWwf8AU0jD+Auc0JJqYbgo2cyIKJ+tMRAfAWCOe48Pk3q7tNY3Ard9JbD
q/wSoaNstohgAsep7S+JuSh3S1o/uHCp9EoaABFZ9/2+CEYx5Pnuqa/r0ZtRyAXl
o3y6Lz6JN704R6o4XAMjYvkNgWkSvjZw5CRjV0IN7Kedm0TGdJoFcFFnWwMUqS7C
aMz8F2dBqzVa0G96ggHQF7Xp2GkJyFNEgh7JwbBhMO0IxjtnvfbIeJVDJfoESCPE
RniN/kMYM4AyIclUzTyMZecTgO8DysYPk9v4nS8ZQ+mUfllySJDu6JhC8RNWRSBt
iw0xui8aTPwFUXXgzDEuCp1UwARFJvhOWzxDWn3r7YyTlwvKkKnF02PF5Hwa+uPN
oMWNkmu/Pu0ltc41EGEDbAf89lZSLYRpxUAVonnt2pCZlHmrzGD/FnMXu3NleCIk
pqKMqsmTuWssR7Tkw4d87ZXZjlfWjyNLc25yzDUUdfXLs/A6EsbQmIcvfgVlpYVa
F7Pz/t83OX7oUQkLG5mmjSrGye+R1xTOvjk9PBdMIvvvGBdWV6Cm156mImwFgxYK
0cnSOBbvm8jMA+WDDl2uaz7Ehwqv8Fjv0CDYQuiC7lH5K+OBkCtf76Vrwf4P9PZZ
4SDlx/jGFqEFAlFMpfFT5L3LDRLWMFMyV180JAyXEgf9AG8WNX0Q6j3r2Qi5xIiT
E1Qgasnyg81c3eK7SGgPjopLvMFbEWNBwREUH/2xMbZKI22dFqB194fzdp5EvlNg
33gR/L6e3wyD+Nw+KUHIWB95P7ZUbNnkLYEUDsRqqSocDXVs9tmde47xxaJ6lE/W
YVPtx+/0XduO9dsNmus+ryhnGmVviZKUwlzvp1Oj0vJsOoMQ9CDHLNP8AELriDUC
9rz0ANH6gkdk0fXEAAQxKKx2mGpRT+mbXz+J5nD4EQNHzwbYtqk7u34Ga5Sn4SmT
Ijyd50asW3FcnQ1ALHpQqA5W37S9qYqqcHmRblaPiiUShp+nuTNUl2CsbpvEpB7J
wMgIbBAa0ZZXtrzCc7IzYMCZhxAFm9e1ecMtqlO6s78hkpbTautGEoeoNDtx10sn
dr+VRn/kXc+soeVzYsRPpleoyUZl0jFOZ4TS8+ZtRTlwenFhcNwsTHsvIZB18JQa
SZlTi1QJzBfwjbYDnUrg5uXO+7MRCfsZ1dTwOkOtaBZg6fB5HWOa1DsrfJuqfDtN
dgkT+mqo+AjskPg+h6xRU737KHg5KSgsbDkc9aZ09ugqzecTD0nlYZMG5QUPkbbU
8Nj15eHyRRXcvsmcSXQzNLyNlUfPgz0DYWtJEUlpKsR2nGf+TQPhsr2/WUNXNjjW
PVrWzCjpZ+SUTjAwAgvtL3aYJzbTjts+uoV3/IMAKsTsbM/V2kchlp3ESrH/hdzl
KHCUzoevfuMYVRe22rq0+5gVdN+B85tL339f+iKEokUh4PCmzUG+ceHsci7IGW3S
F8FVZUYkfEyBfuUjmWDuz9bIC9kdAtppX74J+Xds5na1v6kDMQDQgICMc3jiEfHO
TrezKMf+levwlJozp3bZJqD05jJFbM9QdW4yT5OzM+ICHSdwk7VCUswo4u+euphB
mTs++rDrU+cBVkQAagzsZ2vAka48jRRJTllQQL95gtCNCfUy6P5o4VV6lHD4cc3i
8/NZUGuK85FfMvJ/8TqJOk4RpD0aQpWMTjQJhjKSGrgdmYmBZkqvrf/QzdFmg6ST
+quSKYElmdQIt+9cX/oJzisrgECYz07pcRFyq21LzyjBrbGIYEYzjdkFmlbXbboo
lH6fP11cBKtbQaVq62/h0qRY8L3Rnb/ujX1lcgSWGlGEhd+0MEMwKB7HWzWp0Nqn
2HSQW5UTDiAjEO/6nV5pE9OgMPWnKst2nQwcu3OP6MFA+cB+RmwH6pGOSTl5crZC
3AMs162XST1ZP71WupyU3suad9MsDk7q7GYkCx4yc6ffpy4tBOkRX9ImT4pJQRzQ
8BqsTh8sjAbu39XCsjSCmgeziZ0ebZuhFJS8o0V2OEGYuxsedCRom/8b2sHQeQqg
D8GpJ93aeJPRR2jPQS58EdtCZLYEcRWPyzZvYziRXubZlzijoQdDFarGxbUPKbDt
6LT/x3Ip8QsSgo3I/hmfE4adCxEeFvWZ5TZZbqrlCkVx1xELXMfVg7T0Iap1qnDv
Ns2MTubGeOyzmxYlaIPc6WcMyzT67lP3/Sgp9RBYt8bp6qXeF/xNam5Ruu+A/UIs
nS1h+vRHq1aZFkDtYl4rB3Chm5XK2joMzDwLADqerYuKscJx7mQdFMOMpcwMN6m9
Z+t7Y2U6Pw+31t3oJ0GLCOIsq2d1DUfbuJ9RDEOaDyWBUJxC6XhLpWBKxvqlouRj
6QppT9F9g6UzujAECDzQSHB9xKfS7jDFZk0swLJbO/UcqZYoZ7kJtNjf4irhRqdg
tYPhmPaQFLYf5K156dLVMJjSkdZCtKUGyXQrL1WRaZpDWnwNtqjAIzlMamHX4PJw
RDX5/uV8aKyhznvb3si/7czvMZnXSVUtqalPCto71zVs9dNxzt7MwY3R/pF4Eikp
z8sihVBH+lv9Uk8exSLC2Mrw1RiQcQ7i7KIDiytf8ru6S0vpY0vpiM7uR1D7nXKr
X2HSTBMQyAM6YmINLPKOGrRiPrZXofVRc/2HoLwieIpULqYHWWMQ2TEOs+Ihh5gc
+6oolCldZXvqguLpRvKDaTL7Q1k/CD5NuovRLbElstCGIa+ysYhKXQqUXHYf2cDK
fWdVkPmojAMOJwrRBffs1Aun7ILkb1mgPuxVjTNhJbM+SzcV2fbrxT/3SjN/3TL4
pi5xWvndKEnOkvYtn8CB/+c3SygirM0EKnKxguDXvdqAw4v0wfepvTzORw+Gy5Or
Agy9yvRWMiF5tnKndP9C4JrMvcwLsmJ4pg4SE35dycdFYTB3qADl1CFtC0u1fP9z
fBKm0/tIUjc4KMW7dIhtp9u4mj+7nR7AOmBPrM1r2hNzpfn+P6wQltoSZUttpBZu
bgpsEXHcQRHgS93P/FiJl+DTyIbH3ugAAV6ds+o8NdoXZ79jwXn4oUVva8MQmP1y
gu1PHEckpG6Aa2G9P/7CAL6Nskf0AhMML+cbCKqJUG/PDXy8aEA/xS4dLlvfzFgy
QUFFdf56poyG0F6g1VLsgJJucvk49rjsztAOdY/Cg8frqi+cXaTVf5DDmxqXQAXV
EnpcK8i7wXKLM7zPic651HU+slcG+wT09uTBhyP5XJoBZtNCtynNEzkT9IGBeDCe
JpXwyRm4kgvsA6+EJuIUKYkYJTrNbiekb0EL7kpdV7JH/Pd93lAEmUXm5oiDoKq0
3+G+inKB5gKO9Bso85j3oNM7R4SY4+jrlMIua8FUeW5P4hm2oAGIpO/C7DxOl5cG
aQCHfQsJR0WGg29w+byR5B5oN9AqVrz5w9HwOtCDyUt1oo9voHGrT/H7CzdJAGA4
JB7mGrX5ZqJ3r9EMgrDSzTduPfvaZ/vwrdwejrDmtrwjAsVEdHkvN0H0ailmQpnJ
b5xdP+ULVexHK83tkTnZrw/5IRbXGrJVhzicT5E+dp63nYRLDIOJOAvnkasxPzXZ
1BKoXXQVOS3cWr1HsuDxkXawkeqWeqikp9Uk2AoyF/R5l48iCR7kq+aa3Uk+5Nk0
/XS3BYAkCqfCj27rCoNY5/TN9ALsU9tNiKUjQbA62uJ6LPJ2KM8sTkDW/ixp6KWK
9yLvQeAlgSTRtgBdWdDdvBxXWPzDHmASNnIcZWNIXvShK5+6P8Mt8DvGuTgYBjl1
+uN5fx4Vcvn5sTJlPDf30gbbYDtXfv4VUcg3f3Ra5kn6to65JyjucKr9wsL9j6gh
hBbNjUqASmd2ON7HbkiVmwb3Aph4rk8YZ37Ds6iv5TrgzK3LhdW4Ovoo5/M41q6u
wrl8irbzYdWOmWSwfCZkRZGJZ249837QPWgp8hKBGO6DVYXmGeJYEj0yP0YMABDw
RY6uPSsSAY7ub8NM+G1m9HEcpE9tiekUQqkKzwds38GdB0VBy3ok2spk0nxXRaKU
kvouiV59QBK05WKQtM3mA2DKNYcIpstUug9hZ1t4eDE11friOBNEU7xLSzuKm7+x
aq5i4eCIA4ZdPX301iLmgTu/IpySOWNImBtaMQaG6R+qnVBWamwANsal87+S/3N0
HCwKOhCBaCXfEVUuJLUiUEqvnwPqIKw/rZWe+24QUG9Lg9IZu5TUA1jMy+jWsWr9
EzAdyW0l82x/T283c1O8SEP7eRPb2cl1+KG9bC6gqCfE02iEyel0Gtnram59blZe
GpKvLY6QEY0ipLxVAEDbo0VECVQor0lFAADi8GJzQ54CR+80jxA5FGZaIeTxYU3v
OAHq4dYGt1fRS6p1FIZmo5K9XRCDc3kiddmrP/Bo6LBZexMes92xmBnd+zaW6MQL
7A5erD/e1C6wYhc8OOwsHMAqAgMNy4Rb+C/rZazqZbBJjcPAHrdbtlRlFkZwcFN7
TrWZbsysny3jNQ5ficEAMGwSzvoZZbBYMixs7Y8ZwVX5Vk4SC26mLpvWwU+h87e6
Hta0lu6TAGR6ZJicwBjHJfOlx8UQHuBjTcXVPf6BIhXV1oUtz80ovDIDT0UswWQu
SzpuIlnXouuqtpxuWMo32eavri9I0i8ixkJf/RrsW/06ZKmiuhPJBwFmAtAkGhtj
0m8IXsyn75niSTceGYz+9kCjfKItJLWQ4FdJIUbpyIhUiMH9h3Chke990i1y08PF
GZDEDEWb3hL1xPIReczV5/bk4EznTZ8Kj844nQFjonQMvXTtFNs/mTTFxhDd5zho
YtEHKufyGdtb/+cjJhVD0YS6oiCC/JpV++KnxPQ8+KhwYMe2qhaO8fCbc/Xyz+ED
TpwibjQtYBPOp2gOI9aqxMsmispsVmyW4uL66w5/0lmeySXykUbN/14aMH159Q6e
pUn1luL9ZsfAXWPzeUwPmLOtMDQyMXqDSZF8lC1WG91Gv1oLGKLwO58W15GCSXnt
FhSj+p8cvRhyGhT7ekof9/JSnvyjINjPu8fkYNi9tfeu0zi1AbOIx7f5dQj1gbFm
3qnUM7Peg9rlBMNP4Mgcrly5YbwVZN6i55AlX2WZChpzcjMl2e5MFg2gx+n+de4e
9QHYtPMjx2uNAFo8JkEMxiqVGN7A478yQrVxB8KpjJIpCbw/6Q35dKpwpG2njwmL
1Vh+P/ysAohS31ZjkIv7AoOxqvRVX4dXeePgdE6o4a9o2HQtayHHQbLM6HCX2I4U
Ohn+AR1dsKxx07j7BRnKgyTgEx9X4g2p5fsVMw6qO3ziER0ps9TlibZyyN4JvTe9
QBPpH+LVI5WdMtcET3fAMZOdHEiqHEK2k5GezuyUjaysewSzLIxg2XM9SBpRJ0Xz
jFnqvFBDEMLVQmb4K7zyP/9W2WefEc5f06lOclpPuQYpClcgVpCvd09TwJ0q4a+W
sXBRDot7odRMC13tkSo8uWqGrK2It7mphF66Q/mO6/9ss83+Zb1QR0ihtjMaWGD/
Admixl1nb0qY4IT+jG9jou3ugrOvsodAQOk45QP9hvEABOT9uGPXP7Kx262U4Dtx
r/S6A2uRXXHllrYVGK/hPxJpHLOWQL4lWLXfNljqCPknM+jRy+GmcsnjMGV5wGd6
HhP9km7NWAvsRDxBgtFQ9AEXcwqdhFMl/AqDIcpUttZGHUGoAnIPZfQb8tEVyHUo
e1FXq/zrZA5eySRPJao+4hRo9xWnqcX+cbJAehYW1L44vTvT7Aa8xr4QBTxsJwo9
LrmnOGBEQLVFUKSMjAuzFztLhegnN9cqD5y9JnEQV30N29dwaEjYb9v7dKEVXnSK
AIJ3VxpEe/1zmq5C6OpA8pHjb5lZuhyjiAfc4bhqL4ds/xMRHovTZLY8nTx55mfr
PJjsUVvTAxKn5dcof+HEsF8icCmiOTOLsOeZAYXqddYysKsJ25n/0UAg2pC2YhAl
zy8eE9orGWe+mUL/PGF8LB6QQL72VRq8sMnVUJA3S4Oa8KmHxwA72lTv/aVBA0+Z
SleF3G1tncI69SfF6PqREfyZUwBLJqdl16V4hyeADAD+/IHnZ/C12mujqPKTXhIH
kzevaiVin83KG8fFBLAMNMzvQ8drwr7K1th5GHN3TEbBaSh2NAhraIbsSpmNxI4q
vrRdGwOWDq01hjzvXtdNWEdYdDtk/0JJXOJHSvhrXifgr4bZNHSWW8LXwY8Sn011
48C23eacRVftzl7MwkrDvWyBe6gtdUbmpXRE7Kpdtr6oGe64vzwA54aQhRMKVtlH
3L75CtLh+WMx41URdp0RiNpkE+yKHI5BU0YX3+j+WC2URVNYm2co8BqKYaFLCl1/
V/CDXqMxePuPwxDAO8i0y7JgJRVVT9a1QXL+niI5HiR63FzSd0/C6/5Dsav/PYdS
gnG9ctVaMeqdKrIFDBS27eixN+Fwt2N0UDI4B3gLSF/F+wzo3oqvLpNbEGMkgbVM
LmAIbTaBKM0fC0gr7DvPWNJXD+050uimrbn8FRhzUEMj95DILn2rgVcVRp8vpU6l
8t7SyRUJ8CQXRjIyg9f8/AAG+K7Gq2boDHYRZ87+FTRT0jxCw78UAGIbFSGoq8Yi
gr/KaDEaVt0hVrXjeJNEGF/wwP3LJuhL6rqmjFYEUFRIO54FRfkwJsY1oWEfWjIP
HQVEx4YiWyqn/D4gB4KWImgMoTUe2ASDUwaWeKARvjxxLkyAbyeD21OsGfOFok0E
3cUAhxeErePC/3jkLbIInbbTkji+9a+S8OyKtPcyvx2tGK2eMRMPEJlT4+XaVC7d
Pk1d+Nv3HjSL3nY7fmOHzNRbl1kVmk0uZPK1zc0bWZKO9vKtXsw1NKWjUYsfake5
X7eDFQmBH+kbbRKThpg63U/Gvsn9yDkKUK2OAf1k8YpsB1fi3oaP/72WvG0rp4Z5
RnfAbY42ZYoTvE5Q6EUGLZOpKzB7pZQ3IEgFd9KUgAMCe8ZSHFwevnIrwHO7ULM4
rka/z4dRygFw/AR6OplgkB1liKSW31XXseUd61DKwv1tzVxTSNm8OYmz9+I+Iho0
hH4DNPzekx9wL/UvCYwkHu2uQbj4DsD2qvoD4FrekV84BVpSlqasxImlbUfeY7IA
gi7GWKWm4/uTAetnPUTuEBA05K+xI/RoI4zz2kAoFhfw6/tZLLP+GUb7YFA9o46c
Wr0lGqXHfzyc1/16YOoqRPjYclPBQcGb6BmoXUa1zvcqiK9zNqXzuc+eyWZnz0Gv
Q9b+uUC9iLSgXr2gqwVOsGRE+m8aVQ8UHvx0xCnbsi0NzC3RmTWOHgfxxxl+093h
Ue42m91qBTjREAi8GsyCpRYbZnHEpzUCdEeq68bRAPVdVfXimrE9KbdbuIPm74fi
NXofp4DjlxDBRktzCqIKFHYb0uCVmvnyah7vMkdk0YVo7ClE2mQx5lhm6bj8zyxN
/L+yrh5RNu1i1hldkc+LUP4bBUCLH71qkZLNjg8aF+w+p0W3GshiK7T8lvnod+7k
tGAK/4tZPZLpgn2SIMd0FRcQE9ncLpe+7lTLNcmyFuyO0oPaI4QzGJ3f18t6gNlF
Qu/Gbl8Rd10r+UrMuHtTmVxHDq965zz2WYeGf1Re5V3fAnuGbnaB+qnrWIiK8L3M
oVHzk0yBfXAxP3XUyJAYyIS6aJt8B399J8ExDGSGTQioz8amhQVPdzDJkovicZCB
tXUk/Q+/D9OrWNAzdw3JuYrFh8d1bZ/jiID2PNjx/CCV2XricTcMo62h6nRWwS+p
Og8u35aNUyN33LCMAMr0KzDTn+AbClbk3K6GetMkp//1J8wKRkYhDQgRemE+Elpt
WiOY9lIL5H1DHyn8FB/IXm1gBOSvp0/F25r/JJQfuGkgKfS4WqvkkvqPovzvTb3J
B0UNWkDSkPhHqiU3TlVl4bk3VoMyuWM6z2mtAZTZU3B7yA1OhwaZiUvd8XGUmb6M
k1LiBOamI1jbYL8lBFgsDCkWLmcVY4Jrt4vrBufd+FIRXHNJYvJKBkXlnc6k+TAy
xrg+qpNii7b4zomx90RPYQoEM6XuBeE1DnGWcG3IZiDXu4M04/cQjkpUXFWh7zow
RYzPCbjS097B2sdfMnzyU+NeZzYsKsiwOOo/1hbaAMAg7qPN6j7Ro9mxtskUwuIp
f1oEt65ei1PIIuhO634I9M1pIgJs5qq1YPAKJ5YT3uS3nkpXBOoReFhm8RvnV2/+
wJO6aQBD3vRAT/KZ90OadxN89KVqVWoB2nSWb7D1JHjzLS4uHaWu+/LsfOe89OvH
D3JU26+kvR7D8T17OsdzP2BfFIA+5Nx/knU+mzEEi1OzKQ4DW93ouQc/zSwlrwjo
AsDogiOG9Tfz76NSj+AQ8lO4sFVU79BJDajHJ3ymishfPvtexuzw3ygi2gFy9q2d
14MAPpqTl+6lEsF+gy0J49hiSykreL3R1j+8Gn7IgslEN8E1jE37BJWVTCtWeCbr
BQLFm8Wey4C2FeY4pxXE6Gts2mXtvSC5H+J5+a+1oUA1UkoLkSgFe5cAoskTIePy
yLjKtvXxCHoiUijYgaliHow+x/9QwNgAUoiA3Y/YZE15MkMfu4xHOenwXMyMZv9c
BvaNv33Q4IDI0wFU1gJ97AwiA2ZhIbTRbaWRmMXo5+CoyJY4RI7aKRGS2lSfBd6w
kPE/yM7ZfP81vF34NCDTlWIyaEGRT5ANfRBz+5iOvhcGxwYrhwM4/h3RMboV7phM
MYSYAQFuecVUF5KkYbFtmXyMklSArR8u4CVmQN5ufX3jLGcPTauJYs5dqid4Ue/h
rzJwPpkuuWy3WGKEe0MS7LM2tTOsWwkccS3DjeejL66EMSl/JpIxc5sTb2AWE/0N
nmQkT35GROabG+T7sMXtlsC6wrhJCWZOsaghKtFfbo4wJUSGqIP4mw7g+sIfFPYn
2XRad5GVWf77rDOqorJlzB7Ipf3QB4IN0QOVjOeIdtVJb79xI1yGpODcC4/Vcqmt
MAacAU4GHbniUWV/PTBHvuK52cFFQuIVbHDPt3VirL8RaDrcxJVNnX8oNl16SGp1
rtT7SCavYusfaJgZg718cdc34ZQ6gGPw+07hn46DGbdISpOHzLT0HqiOBLerTOzH
1On1VQJXZNiD817s/Qu5KO//l6emQYcESfr4PBGudQnkFNMWaxfHp2Sr5ael60gv
VYqrBgbqJhxSKkJ7vYKSgyWzoLQwpS7j75vChRhGjL/bZTFul6kxzKevsETfuY34
oF4IK5Q5QGvRbf0QIxe8h67mZE+7g/mj+TbP7spwK9pgMa+QNJdWVEO7vKO/+Z6S
vMCFB5P80/gj7Qchl6uee6j7eaqMkFarSI7OznAghyiYnMINnux0RyyktAQE6ZBI
rbc/o6ifZ8v3JhMEFh7eDM67beRJerh+1M72dvGEc5YpAT16kfyLy/zHnMHSnWY/
HDHPCtvqI9Ecks1VvC2FXTXviMp0yaHFztsncxdFgloiMxonPnOndMKohdV3ew25
gzoLUm1lo9oigbJY6x/fvFuGFgSxe90hfEkHAHbc3jxRMf8F8JOv5bsMctCNwvFi
fByisLgOhXZRIVR0jwekd4JkBt5htsRWc1OfVQE0QdZ4qtvWJv9RHgDRBMIkjFj6
JzvRHboEOWtpU65+irgVFRzJEzlLxl0zi6k7ZGOQ0Kv9Bg7w7EfXlxdbmz2K/0Po
14ZRw02bL1LX91fwtCLKvC5A31fvszVvgTEoI5+HqyO+V4YDmB31FOQPzQK5cwS1
8qjwkMC4Wt2mfQOmFMFZ1dj6Q+lSiQ/YGAUSvMC6CRZuILMbp3OVDQsJRR5zZbPq
rVaWqYPuLhd2e2QmDkrwuYytNBPa5mgAwicmFC0oOf0ajfncCvF6M+C6Ha4HraU0
jyQxIxu7LCzbcGXb16buzexG+CmDo/2xcoh/M1D8EDvopubIuBx4C8iVaKncqyA+
Xp9sFKm1juBX+7RLmgC7rBAUykpQSPv372nbgjJccf/f6Jq0vXhyEasuMNFN+HbB
gjU8F2BfpkR3J0xS6iULqO5xvridlT7hzDy0vZogKLUuPeny7mraTAPgs3Th47cF
rmI22RGdn4ucyZyND6NWCoxCE+MdAEMfBZbJc7VJSUGR2hcI8hF4KTkxjasGYkr3
u3DHhAnqbAgU6sQz1bOsS2b4JJ7/Kc4NVKAms21YhNebX/nNJTSg84P1SKBp/ldL
P3LMsO/jvIpaLZsOVcGY/tQtxuh6X/GdyYrcq9yBwHFsw43E9pkhJRHKf3+8yueh
lsMlBwuvS9PYy31wMGzdl3JKDkDoq2xLVEM0I782mYnMtxKrWbfrs0LKKTwaFTTh
VuV8Xx+8Uva2FYWOPd60ozDul3prlVOOj/9re3hyw790/9+Bx6bgATAPvz7N4XmL
lU1fh9oqvtiWavP4kPRCjMLKNbOd2mGqc/PxMr/j3dRHWi2AgEFLKiWihE/5slWq
pJuYtPpCCDsD0BOPRGna+L1x7ayEo9XBKDg5ENtwtVT4a4XKt+TwzDii6ctvFqo7
/Y5wQyvOcc1N2skUAWmeC4xPeII7jTXjw/ewhpYDAXc8jIGwbpdCJ5ag1mzqiqT3
nVckK8I6ST6MxYsn2k8t5sa1wClWLhzbqnIiZuMjZxlhIyGmJND6hFZjmN7Qo1ZM
qQaW7TuDZDG54HMoIDK74d5kXjKjJdj2Nq8wZ8Gqln2Tv5pGbUWYTmnVcEObbpJq
D7Qco3jyQdTqtr/fC0rjS7fH1PvsY7RGH9cVdZndEkZMIo1f7q7oBYRqjjTNPCpI
8gn5WHkxGTwN5xVM6j8FMEBNBif35UGUzJp41vl8ypTNXsByUZ57Rbdmb2Bb+Eng
1704hPLErj8mvs6YO0D+Fk4FkadeeQGuIkoazzCO2Y+xEhEPjMMZEncbPASFGjt0
A+EIDLVAEnTG2I9K/V4u0A0Mt0ayI+e/TBEXo/pHkMP52/Mfz1K/R7sIVhNecUSJ
4QgCFgZbedcLA9A08vZt0f8Datx8a9sNLImKM1SoRMEMscqY1Uvt6D48fiHJDwW9
2rHDbdOu4EKN81H4MNtVV5FmQ/DVvF2y+hheB+k3xTC6zgu6rwCVVSdVEAQMKfKB
TZNPdY6EhleZ7Az/qyVtgr9ea6zBO5lJCj9Xx6HY6spL7L/ba6I2rBVmrnhQBmJz
u59RwqLlQpV6BEa4EdUaLibaO8c6k2loDZVDOJmuiW20L08fAnesiAbZlOGNCzqJ
Y1dry4lShPAlnJvKZRzL0WNQyvOgw/w6TlgUAXuXyf8DkLDZeKAxy+LCVl5meqqR
Q1qlsJkHoQ1ShNPhYjYNwQ++93v0W69tKcwdotuC2VfJO/CXZ4dbW3tjg23lgmTT
7KnadK9yplwZjxJ9oQiVL0A//44M0t/5ZXicut7fsYcUfjlk+uECaFxEloY6CJ+s
HkVRGKeaKNSlXF60GqvQyY9EkVvZf/+G0iJMc5OyRswwVpqYvmDEnHtTK9/Gk2X6
R5VrKMV1vIyQY9jJPVVZfDKVaQhcUwxRw07PqIIM/1lJCewHtw5eLoAeFJ5oI9Yw
RuCJ92UtroV84c0veDLyoQcBm++GPOtCMzqkTY5AHHdClKN25pacyAL+LKktiTVY
aWooEjXvk296h1L5qJSvFXqevexmgYdir768754FgFEGSf9XwaO4ynD2nLCNJP3S
4uQLzHpptGtP75TdskdyLmnraeWq3hR4p5EjlujB3tkTSZ+dxGTZRWEt0Iql17FQ
EPNlporJ9RaLWTbrnA3iOuK6B62mZTKEqtYigoJ+5NTvMSsGGfKdQoJYRAOJmpTf
6Xn0YrJmo/fQ/INQENOynddEOyrCZxJLt1OauR5tGrnOS3piA1B0Grb5WGoaOZsg
GloZwXm0avh5sWrkpN2L+gywWPry9VUuG26z1IEzd457xNyUT3cL2oX5z04XETw/
USUS9l1Pu5NkLlxHuum/DWuy4lzmBtlhAn7sAaFPUXDVFLWXqJNxr4Rg79iQf1vt
jY6+CkXepKsRq6BC2kCcbgitxhjnPs/iFApOSde02lhNdYHm17zB27N7gtw5Fe3L
mva7wluPu9fB1RNz8k4VVrOtrOcz5ohfXZXCE5Q1+ULRSJf2qIh/VkRKuBXnioLz
Bu/egazSK4QPNx4YyH33tvzDGR+rdlGw5gsU+VX8tJ7P4LboqNlessKhyS6s5ULB
xTlO5BoztKGmECrkflbcRVhBaSoP1L3TL8VasYyQV8JeDfqe5X/160AfkTBFGxQl
XpdauKdXvGvVLJrWnw7XQ5UNy/Zp228L7QnBnmGpfHWosxpwlxZsXv5WU/gpiS39
ikyMIwKpQLkN6w8f0W+an7DTKKVdKOqCyVDu69Wda/odMrCoh6NIHWIAbLxijtHW
c2NUpBiyF8BvBcHvxYCPtiIClWfK4Tj01A5TaWrIdoN25DaP42VR6IMsOR5SB6If
ntq8U4mIOVy5Z12cduUCp3LnyIV05RnsFpxIt6jzfjTRiLVRtBrvTqCUcxQ3ZOkz
cXyDxEUvo9iFFPhexoWs0qPHdutRBokUxuAbM/m6jOqHWQGw/OYsmN2fEYCuJMcq
5yptGRDoJ0s2kq9F+koXBSz2xa/YkxR3noFZhoc4RZ56le0Q3bBfcqjbzreHAjg+
98mg1zfSEpf/cayEbFh/u5OxxLMpKhBfxRJM563HlnzdTXGNiPfJjoTIV8GUVl1q
SS9PfyStbPsMWRBUK05w2d1Vb0l0sp1/RcuGd0nYfa0wPyRcaFnlSomlDYrM04eu
cJ+kPKFKmB+So0bfPPGhdUKfp4/V84MN6ACNA/lkftSkPMnIokUsRkLUPuFa+60l
YZnzrgxtwx2SRXox7cDcpupvgOz9qDyfJwaDPkN1V1Nzu6SwhAPegFXE5ffr3H0E
EjsF1bt8iJGyET6bds8lXx/MAKJuQRvHWfiJ3Ra4Rgg+I+ervd/TvAocf+kHI1fH
vyb2HnNXlV6HJ9MMW+FF0CIwriKiak5m/nPu1UuTgJMJhlOOfNaB6BKme0YZsa8J
w0nZ/H8coEJeQEU8yqpFJ7epk4cAWjbyvyb0Jr8A846bLpKanR3dbgjkNZtMFsC6
dZxysMNnPBxR3VG8Mn9Lcn7OkZuZiirOTApjbm7GJt+flzWEO5QNdTlyw8d7FOqt
MeQLVaerc6PePZskCktwjsRXmsJ5AgRjKJlviYbT8KvMN71CjIHDMq1bxLR1nkKv
AMzQdzUbtSFDrwzqwbAOLr07iBFfFTiuA8d4r4cRloJUob42n+lp8kEf19LXSaNo
pow2BZS7WCICIo5ZrEbqVnA23tLKYCIj+qykTaDo+DShu+ph5Hxtxjk7aoB+rS3+
FXM/DJtVyjUobGddr89Rie9R0H89106L5X9Q1CZZZa0eKDNCLiPamyZGgyFBLdl4
fJlIG4wciVzxF2XyrPa5gKO8DvByxt74XI+dhFPnzFGPRtPb+ZSs1wrsfnUtQmgT
/QkEtGPIkFnNzq4L/si72KMjMK+M8gnyw+ItOuNNOmNtALvyF2UiW+Zce9LFauOS
sxeCR4zNBJOqbbHJqbvaPZRObfVZNjTh94NwJ/y7qTIve+QMl/uV/pZv27HsHZwX
A79q1R7WSSvGJLR0h/buL5564V6cXxP4Yo0I4xXgnukxtr693Pvj8cmy13st+qGy
03ju9DE/WkNANr3qj4yrnMXLEvL5zBFSFOW2ve5JZ6c6on8JnHUvRA9eRPgETHjX
vFTtP9sX2jFO4/Id5NtpnqT4UUr6gWoHVdrA7ytFOVJRpA1Q2auybViX7ujJu/gb
c/ugYoE58LSm59ZXn277F9hGrxCiwd3tSOuS/VoJF8n2MWa+iDRKBlUuMdSDqZdW
2eoqHwZhYUWTRFDQSS/BV82J36nJs90rpGYrYn4akt14sTcHiQ067aM554RgaT3o
Si151wiMDiKS79F0HmeTr39KJrxncfI+wDSqCnFYHajmveBKExdqA5Pdgd1kf0Xr
iUtYaQJxkjg8Dq6u//HIRfJr82slJgxDhM58ugmK+ZgbMtXvhte5NEL6is6GUqAZ
u92g9rPNxUyp7SJUZ8g3XKS2q8zNGcNYzMW6pbJO4ysj+AreSqM2D7pLWazSH75s
QjtpUvrTWifueoOWjZiUvqTUYLNJFVlaMJQapFByKJ1tlCZqY5VE4izMtrO2EAqy
cJnbjZQRyQNdnRUpUJk0cFO+8pIKgoRfwkFsMF0DdG6lxK510KjCw+u8wE5gy7sU
IIYSfYsyn4poO2kNoi8AnktLulZBVQ5GQRRbS1DX0gftOTCCVwTH7yfsBu1xTw2M
XNtxnVy0tBSCEdrZrjHyboRXobkjs3IUC2gWSnO5m/Pu/EhlObf69IpPqgSFxQYn
8SG6ZFtK2TAPTbqOnkraYUfPS5X/LffdpUjST7dOs0DAMnGwuLNT91YqidbgAWlH
xzb7JS21Vn8bVNkNtmoB5hjRx8fbbsJ2Hul1SpwOzU9OUdHRdCZcM+E1ZmhCkNxy
25DwV9LkBrqtr0u6sIsVEe9h7vJUx8/bZbwNXz9wKtSneo+qQabtSwAMCv+YXRcM
FO4UcL9+Tgijkv2Sn1s4eNZjee2mnitBsP4Kf+tdWLiomNuzQC4l4nHPaSbCdNdn
rOu07m1vgYPu8meFP44/AKav7hl7Em/mxPVkAcppTZgSqGb83MC8mnmYYjeUvsWp
5VWWuFbuIOY7J1c/5Nc1uSqbWsFn+Yp36dGaZej0bFnMQlR7AiijejRxC35R+ndC
ukWpmZJUT+Jf4EU3W9AUFzb6wHPrtEkYmKRVt8DElcAA/rSRjd+pN4nc1qRQsXCP
/l1OAkZLIz8boWlHeRZSnPpu+dVmki4Jr4AmhdJGri48JKstqm+GjPYoB28JsqV9
DCpursq3skHINiPDVyH7+/+2HA/BdL9vchDYw4ufIZfXYthh//jiNPls7VSceG6x
tTF68WHEI9UmM3WbRuQ8ys7A3qcufJ1JNDkdz4XOaEGbPHbaMb/7N/dv47PxX3Nk
rIwJmIKvvIDPDF2H/YeLq0QlZGSAEdiRR+eUqIxdTvhHy9R60wS07rYLZjwpS9EN
3kLdf+U2+H7RmZCe8+HmW7oO1140Xy5eD5x6aBXMpwJqy8yj7CIH6Xulh7xUYYRV
F48O1pR+3CELL6pU/dYpgtq4ivIqkgeCJdw14zJ83f2lZFDHHNBD1cU7+9V9bgk2
2ygWoSXYs7emeH7EBENJptqaVc0wk0pvPvh/aFu0/R8pXnoFV6UUKKn4m78MiHTR
OkJeU/TBSrOK9dOJT/2pKr2HdmKLGGXk/z7MwWGqzxEeL/igBOwW0GO2GWstLhog
a1dpRXvQswkAW1rOP0smCKsYelIR6aLs9G08CkR8w426FaoMHWBvSuE8cBiwg7bo
YYQkxi8Q06mUKnqrBbLB4h7NGd4rFSIbv7zVh6oJ9G6CGYEJUhtvaGZfYehj2ref
4ztm0+d2z5HclKwTbbJluVtVNKJm03uAkan71EH+fa2noT7D84VP25jvoGORojnC
Ey+a0Tn2wUHl1Cs3jUHW6/JVa3dSP/l/xUVGLtrtHoclNtcxhRi3c+ljc61DDR89
Gt1LWODR/7R70CG4sls5cRoikgeifHaY3mkTsfnzJ2f4iGlaMS2Enn0hT47IMs3m
VlMYPIBvWMOVaJXSwWanDa3wDcIpyfe+DSLJIybLYDe4mg8PrKbbBJ8DGoPh2t11
3nkO1etzMKugqz6+8j8QFguBtpQEd8viDOJfZOUWSxmy1PtT39SfjQpLQ8u0x5K+
azF16/pOF4r7OKeA5RDT0af5Ct6vvU4ruDR+s8MZLmwEknoGqnNhD5JV1jqzugOQ
J/6lah+PVJdHDQab5pYDW4GbN7tUefqogNBGZYkdC44NXKWTa6aJ9AqeMEqwD/k8
2IZifbdl5ocwaR/miD2i4cWxJZNaxnrg09npkakN3LPruYn4L3eYASY+mr7Xkc3X
JusxpQrgbnxNrQJ3NTyyn3q8EA9gYEugGqB2iqNssoFwFmUAhiMVzOdqlkOctDfW
f6XheqLQFV4N/O+ps3ViY8nvDNS6oANCOo1yki5BeR8Z1YWFnc09del5bX2VEoet
ypGeaSPK9BZkt9d+1sL3NHKk7ftLqeyGi6XY/4eR0cCmXMvSjaM5qneyxaUeiYDt
elcv6qYDBFibV55b3eCN4kik+ymT34uWfrossUVEPhmTZ5iJATmSz6TyS4tl3f0V
76wAyrSAGcXFHtYN2fg8hvGNJhpn8fsZhQhUydr5VtVjgxbcZ/OPGnJU+BV2q53U
Fj5tHCWU8hS4sMSCKgOjbwSJ/exa3zOlKS+V1MOXmF/mLh2U1oNPNPSVp7+fClnJ
mDj2QI3LUYiA2XzfZeZDiX/9riDJj7iEJe65Orp2Xf90VJpvvILeK+XfgceMxw9f
43dOyhtxRS3UcVU+dty1xrHkfinTMpqYaQrS/+HH63fkzuRmJEm8XnyhIs1ZuOsX
j5ucp9JL471h1BSzP0lmLKFkmkb3nQDIJoBVdb3gBNXxyj0FjeNeF6vuADdME9At
gB5QWCxwRyFVhu+G/Uy0Hta/upC3I7fNWi9pwTAo08CxoQDpMMpl5ky/+3eiT/rX
PNbpc5d7KzZKnyLpCDPvyvZK28mweJTHYbp9NXHcv0l7xs3kRAFyCZOo5My2/h/I
FhpqiQopp82YShsyjWqjex7IS9usQIh0C52gxguaUKfosNv8GG3LypXKOI8mpMh4
E+uW+aO8+vQ47TLdFYTFVYXNGPJASz7ac7/uWrx/qiajIV+7iY48JiuSXXDnr085
lXWx6DbmVH8gkeddE8A+RmLuC0rpBsDyx66+ezrVIIyq4GKNePReOFEdvmHpgRs2
ohiXa6Sz5kTBO6KUkMeMp7sRQJbh+Pnamf9JAZcE+pIFchx5PNwy1tDNa6YMRfH4
A4+IosvbmCeaE7n8vApmvjw7QVry3U9tWflhJipFRHfwDruY2DqWda4QyZIu+NFo
UNGptpFjs2AvjVyW/7JRxTIS1i+add7Ns6t0b/HtvbC4yGnilOdtuJF4qr46jfuL
aBGxkfArz2VVBxq9w3sEt9Y1ydaReRn8epYje/MeO08YY2hLlyF7QwzAlFRE4Bw0
wGP0kbzdy8Rv3eFQobk+omEAwr9dbKrHvFPrWOXrLRfDgvisorflZx60jRpqoXeN
2Lcmpeuky6MByBHPvH7vJUhZo5HlMvWxsTY7rCAm5zFp/jwdx4o+bSrHLOnoX4+f
lKt02C+J/bF4pl6lsJNJiq1qVJJTQZSZ9nu8HIlWBOGyknGjF6OJn36x0ILCdUR3
0MXgpqknCsX3YXvH6jhIYI2gVPRGfn2BFcRueImjueZi+jkFzvhJqikuql+6vz31
vn83cqTdF7Qnh/+vxcMgwjjX/uue6U6G+sWoyvuC+nzOFpbgHD1qFR8tUh8iz52B
QDk5TBg0dCKstYDWsfp5+7etRcjbzQioGy6qdPyDJ1iNDBHwdLsGxyyRa9CmtYnk
UPDLdHXS5scVU0xsLyctJdsoQwh3TYup3Vs/S0vuA1KIerV67ZMS+NRAOorn6Aoa
pvLcvY0KlE6xSt31WJ/GnUHNpugz9dnaPVJOs9OuSB0MNc7rhYGMpJDvqjImyoyf
5IEm8ztbKiyS47ZBBnJYDWJaWW84Hu1rj35Ok7ljs8+Efr2O1Gv0+KpN9UM7VQRt
Ym1ePQ4FiJ6J3WKexlg+AEQ/Z8g6qn6NvahudGcya6T9O4cSPnIOK5ZYcj9roCBm
llnnDQqpSA6A3f873CxLORDejDmJWyj3MO2PQhE6ITrSI1exaVBY6I0JROS9W8JA
qWSDNZv0Jt5lp9Tub4cTEjop847dv4KRGBQhHQ5ZDBRFp2K5ITfsFXimlOBLvRgo
4G3MRc2zsacKzq2uhdNnChKuG1aCS/QDXHtejIQADPRW605VDU2OxiQxfm1Iwdiy
AX/BaXQsc8zgysJ6bzFHJWYL1GGMdQiFwiXbEGVMQC3xy5EsWgeqnnBOG7vkVfu+
qiI984gFNa/7yBioO/1LDz3yhQH1BZo/NBVD1VBOr8cDzzp67KwdqngtRadpr2Ok
WhiesJsHKu2s6xD8fiaoCgLRWEmA6J3tGg5BhqZ/K/GKHuVj7T9VJTvLbJb8DGmp
6vEAi1GZV1x0cyPr+qWozHaCDrpY2bSMNbujylbiLVH+54dNiWk4hGrvV2k9zk9z
QH0rNs3hGOhg6XI2r+S/fqpb8e9W8PQB8v6qaeuPZjfyorZeXUVP//l9a13OyucA
YpxJcaOVKgBZX0FIwh8F4VlTodbVAzZgN/oI0MruoJDoev5hwRZliaDX59QTbDai
AN/B8rkfwwhtpZLKAXODS7X3NBUYL/5xjWQ8l8sN/S/hCI+1E4oXzTlOP2D5ySB/
8j14W99LxCK4oSz5PuLiUzF/2yKb0Vspzu/x4R0SNCE1gOUxwnLQa0gRF76F/tk9
KRe3pXtUJqPFrPsjPF618RIUmDVRWoZQW2+Nz06NLe6lDWOIoSW4CG3/cpW8GD2Z
m7erunoPkNtaqERPdiX8rfuXvNIUgwgYny+MphRpxVIgG3URpw1syREm/MCoOBrd
gzWfB3Du/Uki8KfkZZ4kfAOQH6aqf0FGyYT+Q0hijprpco4Dq82RnFeraVyZldvU
H4OOVE5dB7048W8mGgN0iIFpxauUNi9nEX58o65v2NgEtB9Za8ZkEeH8lujyfzel
ckYmCSuIwC0DdmICJFNUePGJ42QDG9jBk0DwU60QgIgWqjZ9WnJPNe1WoQdohlTS
ImQuKEMQO5Vz84r8d8GULMjjVrMdcb4lg8hmtJGBFLpffJm91hwg1vlwasyv7SXj
v847+iTg/y8rguwzIZqgI3E4WN6xs8mxpeQ1++4zAxi7ycFWcj3d9cUGBczN3/g7
Ltd37Dp+CLW/snHKszuDI6PgqewUzR3IBiduASFlThXSZuRZvyUHIx7CYPj/7MUX
/Eade3jTk6MVdxyqDPwdzfWQNQJx6yMSeqY6tAYYaRS6F+nZAqiJLybEEvb4qMVS
URISOBlGO7q6ppJnAEA0Pnd7Dp3H0dROj8IKBWm56A/+t7ICr5QHQtXKywNoRBKm
Zr0vCVuR04LTbm88JfBSEJXKBOrpDr8onpH1HFX0UvgaL3hApJ9yYOrp1Kb16ihX
wejuqxkSl//ObPVkqDoHrIXCcdmPK1vvIcUyD/YOAxAn5D4Ly47Pnfprpt8PcjN0
fWxbF+JSodTipyHgXlDkvyhM/R8PEyUnAv4ncCj/lDUuS1c+/wGVi4z3sqABtziD
O1LJgNXPT+pKXiK3trzRZLFr7FbMy3F5lm32gT8SBRyzx/IXrI9D9u0IMm0fei5p
Bhc2Vqrohx9I9rWJU2aMAS21t/pdO+CxYCvwzV+s6X813nUh78Zvf7BS17HlcjgS
Na0iq7M7/AOeqXHnjPKeaTWbJZ3142E0SLwYGtvfbgXpAHE0H8QYye3rEY8wCgpw
aLqjKMeqwKupGw3wGEzJYUWdkStGgn5qax2Au85daiEZg/Mtlusw9grsoeXuAn3B
ljSvnd/O5UC7KWy686lRleZ0OPRPyoysDKOANMmiHAgpNbuvQM5kwxjIv7Jn+jhi
PzoIIkfF6jJ8RxFTNgS2rx+UWGMKA1QfP1uVHiaFIBfFCE5vVpEbGjd68CNya6hP
fAXtN2kfTFvRDdfkhuhdC3opr/SBv4Uzp7Per86ZAEXUUOzHR0XlCQj5XQTYvgk6
2sRSDB9giVANIq3YzoT+3ydsazFMY1Z7q5r1jWTDnW4AJxPieH/9MggLU7WVF8vp
T9Vg9MLkafEWS5nOR+q294kr8jT1GbLIiYgD1ctlOz7NrmtpWPn0MQZiRs6pIH4L
JdhOm0K8wGH+uTy2o4QnEaWFQlqE3HE35UMcHI4fBE1gL2yjQCOZCCMLHQCgKWb0
CCqQJ5PJRP9ZSuK6b6hLEyzO/OXC37NuJqicHRn+vYnLfkIHr1qCCcO7zea+xPwA
CLLpv2GRLuPcTlZhVr7Gwub2DFWNHI93+3QecwKKImdHNmBh9iCpDj2RFvcJY7BM
VD7Susia8mhTJCZGcQ9y6k9HR/O4IG0xvjPBnOXoYrsfxLo/fsgcxd3SUxaAriJz
yVZjzFP5M4rbO37G0VCHndgwQxE4OQqtGQp+Vqc85NeWMz4MRNxxpnJ0ZTJklDrz
U0L+w6emdXWsdLAemBPu5qvY0YVUHwXtqSAs+Zi1OefQp9q00tgX7P6W1z1CvCt5
tAvazhycKY8fi9LPbefjLCsvFtFDlG2Hs83HuxO12hspyw4QYy4ZCoP9qlgxGAsD
XUPunsaQ5ud040kwTN6piFLP6EkOO/XssR8LjXHtJrNFt60z2pHjJYgpVPpsum3N
CCISf5+f4QMTBB6BGe+5R0/eCzb4ZS3wHCZkJR36hsWcX6aPvbp6hBp8w2R9WQyC
liAeCBjIFo8Xp0329rBEFqYcibKyuLSUyxS6NyGWHa4q+X1JBnWT81lldRscaY1c
eZZiUphgRm2g3jd8TLnrLVVyBRL8NycA9JzDRrnIC//sGQ52DtJnblcJBfGYpX8U
I6ZalE2SLCLWb3wSbuPSIEBl7XD5YRPiMyV/dCTWR7BfSxgTEq2M4hv1StHhZ7Bt
PW/B3iUhLkNid+DHhpRJd1K5RQ4B8jR6YrW70UQ4N8LsWBj4d7/bZRoNydFwqOqu
1eOszq2daRsUu6aOf4Ej8KaKagSUedVjsueE4LUtpdQFvVfjLtXf63dDfuHmX7g9
9XbeQlyn1TqtPSQNn2gFNtKLUCz4sushS6QF3giVhSjNYl9ks8i1vDeAx/bDgT+4
81LKWDTHAW44fj9JiAanyMzDzPRBPaP0bKjjACSFRzvg75zYSOJ6xfinchDXCz9w
xON/19Jqk+YRu5xtoDBuD/EcHtC7OF+6fQx3B+SViU5ktuf+YXkbq2QA+LZFpry9
mzvsbnKMiAGnnZOMnG/yD1eFiVMk/kZspxtJkFWAaxL5+WGpXrc4qw9X+FM9YOwO
fO16Ywgn+jVC/WYrDsqrREUj0KVh9L7W3Mtd5EfEHVJCPQ5u1ebTl7YyRntkiWcC
uFQKQNpuzkauRgqvHh3PKs2IY8Q3SR7W0yJjYvxz6FX/eI0SKrRlZTX5Xn7zX6k/
xgnnNv0QNhNbixDEufY30kRkKrnltcRBObFIq/4k+Mn2N5aVHeBDOXOiSL1niFn9
V1YV+mvpMxRF7T36NVn9WW9QaaUnDpVK46hMlIaonaTE7pka7+rXIgDGY19BEbjp
EQhc7Njo0SQQYuIfoRtFmVq/cYh5O6Dt82AGB9W9215b+NqdDBzTnHBRGi7mGKS/
J+GwmUCAG/tMrcXJqFMjCaZOEWxZ8fje18NmCU/N5XEsInAMQi8Q9b5YlSaq7+gH
8pnEerzzTIZaG51to5UFrXCKfgQcITSPF1/Ab0yk5mfS2NkrmTkZQpADJ+CVHk+I
4mbw6DCjWImjQkyqs2QzWQvLzH6nqHMAPS00N+g29oSLqOUrlEotzBIFEEzG0AWt
ugCCDgCnYQx+GFhpgGIY520X6URpDZVtSXWHxNKb59CCHuOo1is/wzTJo8MgsDFa
bd7lRiUb1RrodIdxo+XSVWqnMunxAiyI2LS3HcNs9F4MWiqxWQRsHe7ujZ8KajOk
WAXfbaXl+YX7px97BDBZmvC+1+vHmni0WUdQxLRpLKv83g2jmc73aiLAfpfoqDlZ
b3nhf6YDrnYG2DFDAc3sQeJTsljKEqtg7d9Pkp/u9qreC19peX70vD89hcOUxlxh
tHUJpcP7Z3VchsrrJMTdyLw/m5Sx2hCve55pXIv3zs8jp4CDJrVChDR4ezgrroKj
4Mc/Um4aQlqfdcwTh6IBWfqC/OxZfu1X03ZToPmWrc9coREBCSXKA5eesO5ggsuc
Ea/cwVo1dAgMbZPtRT1UspukCakGNvDfDTCJ0dYYkKqf6VkQ6Hhs+zt35JSc7emf
NtkDvVSJvPytW/ESBFRfieOM3dcgUevE7y3STbz3dEXJlpzt3zpYK2GRHf/rZHia
vLzQ3HV3SDWnOMGJ43q4pWVbjB2lhDpXZcnmgl3NDn5Rvtpu73pIeRG1cxIhC1fK
6TDhwH9SMGNrSoGA26wM5ekk+6Jhdv8+bfzHSjI6MoNWpmIDFTRx/4rIOY7LjMsN
b5qEc2Q7FsrsSRGLvgja9C4Dv78R7VBS+Z1VBSdrl3J9JJQ5Iqrm4+Xn/H8y7Lov
axH4DVMpQF0SyYgLsKS/K5KcreI3KF5H44mXmTOQRw8Qsc5ecHn5vKpJtS/rnsxC
BgE8/BdlfMHfPcKLtHwaYkwW/cf0f0Z7BXu1l4WqpfeSn8+K70drBAkeIVZHOGoS
5L6+Lvn9N5u3nOrXhQ1oA0g9vGPiEqhMifGoM8hWAjUWfsyu9XKi1iLnwXVGdVpH
97iiVL+VdCyYEROlkBZVfSULN6CeBuHh3r1JryPNW7CVt2apwpSlULyVmYemSbo8
Hf3Ub5qIHaNOV+t3+EpBCIClXYiHmI8jEMI6xFGRNhjATNsdLz8vyJXJEnB7x/CS
vLArqaHIjwr8XlaPyUqe0dyIqyDIkSDqy2cPpB4BpMj20g1cmGGJlMXriw+lZ7OG
13iDpG7wkQlOyPxcM4LXR7FEETn9N80lHub6MGWq6a3Za2Ck/rhz6FzbEWeCFYgI
i6gw9j+v6MD0TMuqz9hNXtz8CT87hZCQgpEPRsrdTAiwY5Sjn8n+z3uV5Tmeyua3
WBkccmMDRxal6y3Y1Ry2COw/jHxKUIjet9cMB5KdeJVQMr6ShGL19aj0uSZui+/3
cIukQGKrexMQlIopqhtlioee81Ti4JdO2C1MxUTCdieoew0YY4t8xpUxIc840m50
MhBrqOg4pqGykHlsk8SwmVycH58J4LPxTVFI6v+QvBEOxQaM4bNUgn8+TE8LTTAE
pi0ZgkmeXKxHgn6QXEkWSGmtDhIooSzGA9QJ4t2OEIiC2cGJ7k5oLAYY7ReQpiZ/
8OPi8YT2EKJDIzWNxM1da5FH67jdOHhf+JN4VhMndhxQfNj5YqWts1hVoSZllfQW
CuWicnYs2/7xaUS3YmuSMGMValuzyq2aPAyLPmZWzzB6uCAkwLNbKxb+tVGa1sOb
vwpYNGaevhIVe2N8UN7xCcCeB/bPJG2DPgPJ76+2PHYkMPeirSveMXrtbhwyZ/Kc
JaB9nI5HfFt7CCb9+rUTLfKZThdcJNVoRiTlFA/hZak4J6IFDjvgn/eG3btOCAjb
r0PJIGVUB6ks2zku/0t/kGcZu93we/Bx7rFGZWArW1mazPkYajUn5hU2OUaaQnbA
fN2JACknlANFhOFQASRKSscy8ztJl1qV/aZFU7NIEmK2d86ECujwjZwDnOG5nLWw
F99s5o5tHpC81BCJ1ZtbAkuCBfPBTMDPyfShZylmKHMfagrVWM2qVf1iuS6w8rWn
mhwvfaZOMwB/zKL2fYBQKZFr+dr/g0YKhyG4xdwc+pOJ1rr0Gg+PQoinvetzcV1V
wBtcZEEMxQF6AA3LYp6HdcDIOaulX/Kw1IM3eXVgBvRUv/KLgvUHzfHYlFCx51H7
Lw6/u9qac9pSFEJXlNssuzO/sthuZU5N0jm2WoABXpmSDHr5DdQ1vWv3Q7vhPN7L
as4PzUEyQdh1Kkqd2R9YVeGVmQvy8/659w40J05VGSzfAgFhA7xVSWQE9AVuancg
SdFL+Xji9FI0LnH248+CBH1+BsTaDpiU/+bCKTrp4ZXybMih0YJrQvdhNE66iVw+
y+Kv8AdS8JXJWhAeHOIasu3tav/wMKbrASBIMeSsWR46T04GIXrkjHTT+FYL27+M
uHOhmjbhnHhvCrOCu5DnkffXRgKddL2jUB1KFlchWUgZxF04PcA4TgEyYhCruIDI
PQtaZcALhIEuedawp19gRWgrPGOH1yRdd4zAWQ4ozDCYKq4UeEaG/I3nV+iec4P9
RzS4hw/d1hw/MkZ465DGWmGM4DPtI882FDxf0yJ/DENoAJauOzlMo+Dw7ltiiAWp
cnlP6y4smh/G9NvKxsS9XZ7A0C06ac+ayhdKkz/qpUrjplEPOdlpjtHWRJ83e5pR
ybCO9X6y8PfT+nq2PUNprpmSZNwLghxSSofZ93vL9sWgIVLn70Zr2yyO7OeI4ZdZ
DBRh0KK4hQjWocQuIgyoxclrASDHOPb2SZbK2mwPGxbiZR2q4IjgDLyqdcIkq1wi
9PJeOpJJmForzHVLUMEQUq79U4E/MB3hJT4l1NRqraIopUDb0CTu3MyGzXVyr+gZ
hRM6H7TWS6Wr5i0emlS5RByTvtRaQGEPYDnFPbu0cYVzFDrm0vgdgudNSTQ5eTIS
IoL8Df/+fAXQrpJSiUr8OvAeqpCylEw60MVrLMYHstFNtyJSfI1lDtkLcXe0laAS
a4EeakzynM/vPeDPIv9TYNzEyjbP438T4iCmXfE5sns5+fSpiRVp5np61ikEvOnA
X1cOot39ZLXxRyGcpbn3wvUAfob6Z7DiyGImeOljUOwAIShCCXlQrWpUofLdawlz
1b2h7/MZWEVNEqP7N9whAGeaFC/7Rp93BnCMcTmC4/xeDe34da03vnFvNY/smyqY
t0URfg7yc99LXZJnnT9STP7k6gCUMtfp9EplLqWjkFuGNWKC+uAtegb1hUddfhuv
0rS0RTsDCGD3JaQW90bZ8Xd4ZrXlm4Mr7lwCVrOBzbB8ill+H+Dyde5SuZfbwQ5L
hQqnRMg2uSiQBHstrzVKv5O5J5qbT20FQvFo7YsckK2kkvLEupEmeS/BI5M4EMCw
3L3stZVkbTQO42+jbLlirUAFLh5gCTEzoV+Xm6wMqDKG2n7fbjf5HQicJJzisvz2
BdCRxZssulUpF365qFmjWldxm1l7zKVwHPyoEofXnWzqcnb4U6+ijz9NhUn5wl8d
b8IRIuEVZ8ZIhqYrkV/2hlK+uKTqBRX+/TBVWTsycWI2mB5fV9F11BKyyWl91hp+
07gfQRkD8B37hwmuNl5h7cT4FYsN1ckVRrxXq9h7MQaYtTNn8N2TXZd4DkfgljeY
REMnV+d2x1SsRpXdtIvV43CuqQVY//uaEIZBaDA/39DgCWLSkZm6VwQJfhqNpudE
dMFGqxUWemNlTpbc8SsThYgJqj3JDza90aIHZ+8a2Lm1RYZQDfQCSFeWItM9iv8p
qvYSGPajAhNLiFKjIvLZaUjiFt1h2hWx/iMgtGP77ipBOWYewMLmk6Strb1p5pEM
OUni2X+l7LJQzL6LqORESGxmRjZhn4VQ0jNIL3uuKXQd4tXJXUwISrFt4oHXzDJF
KU6fk9SuMSO+E9NYjRJdEaUpseD2Oc2aOtCG/R3qiizEJkw1/OtQVwIjHJKSC/dG
AM7M4mICVJju7ft/BKvXfWEHvXkZvkqOklHriCDsi4AL5h27K86MiU0w2eePQEBf
CtVoI1gotMSmFXDNMC7chkCwp2EGxkWNhEskIWOGOKBsGb+k2GtONYf69l62m8os
dJvlhJ6j1Jyn33S8oOBtOl+Ks7u2TrrymXiEdsI9P+ngOtRqSrKoht2+4q0E+DNT
qEJaljeYfwVFDWseFbwRwB2zmkOgnssd4XiyAxhTOgZcyXTr6i8dGB2xSY9F289x
2kru07CmGSsQ4UpCQ5El9x9WJ/D9TZGq0vfR4Nz2JD8yQtIY1o77DKGxctUfDudo
VQPmKe2e4ATDUM3Glla5R2bxz3sodQfuTkRaIx3IF2wcM/5FTuZK1Ab1MZGk5vkw
bSdXI4Hvy3FpsRAaK/+KUDMpss9UmFsrIIuYj5uHMnubagJuPFvRaXu+AmcBUQFh
DZvqvo+phZyzPIMB91otT4JEG9SSSAurLINSeenqOWiN8IKsotvpClc242FfkulB
A+2s4xSyiyCa/iGH7DQJ49I6n4Lm2rkqC7AfIcq9cASzcDYkNyxURqqoNqr5/Job
mxmKPALlOoTyeWv1x7stRWoO3/CiLO+amqH4UFGvk6x16hwiDd1GE0DbhuhtVmRf
zib16X8+YE2oaqIm/Cp4RxCrz4n32rem8PncbFdunANUzgrn8A0lSKgbJis7r8P1
6x2i8g2vwj/geMcnuaJRJS4TsjzWDF17gNKuFTxRVUZbv70fgQ7ujuzYKbI5lV+k
kjcuUo2Mm4rVQMyJcP7LllCUNbmq0RjRBxQbmcfjGXM2iQhtPj0bAKWHty9J4shx
YhAgKA9ZGJiev3OBzWhBu26ssHCcw7VmiwavmM2hbkDoG7yuWTF5UyH8FFdT+feg
uHw8aoShLoqKTHCFposvyTPWd7BFmAL9/nv2JBq2zo/DYa0977+t+PwzOphwrLoG
f6nlpcaD8dD2XFM2WoM343d7XKeeriCM6al7siDsqiaAcTj/ikz5KS9w3v4RgYrl
c+9CfZ4AA/EXrB/WJdVTGWLmS0FvW4lTBXihj8+o3OIy8c0T1/MlDmwTRygP11n5
7JIrX+hP6fAH9e1MeSY674haSjgjEvE5nCouI0Wc0lIQikCSY6OI4dXK+djAnS9h
DJ7Dc/m5GKwWtDVA9DZBz8gYNU3F3b/RzI6rRCtDGPJYRdw5+Jmp+UHBXyXTu/sa
4ud2cSkX0fGduB+6lAlW3TWR7WQN4nEhaC7pKYQ2Hvo/54aDTXFiS6pyzZsdaetL
mBQ5WoZm772tanvLTkJcEpNumthnqwVBZkzKqnhEvbBCUv9+zSXliBX/c52JFv3F
TaTCbrXCXxaY5yGv78YcM6fPzGHFFcqr1BelevZN8WGGtBu2Y9AlCJmupmrmb4WY
+qmDzj0WrUWYfn5R/A+P5IqqNb4OGKsaM8rQim//9UlSkACvisQFtpEyBZefUc4y
c9BnEFson9cuZZL0gPbHvl0ZuPeLh8WZzPKHJrd/wuHMbXPuM7vWP8gMCXdcWATo
aNh2yvDvXcMIU174so5r47mEFxe548+YzAXNo0Klz7BzYPxSIqwwoixQmn8FV2+7
2nx09r3BgY4mpMah8lqUuaX+9rLK9QSSTSCjGtOkF372zb1I/+Hc3o95VVsvucds
0aZYqvCc7ZQOX5jl3sDIegLA2+5umqZI2eDoU/kpv2bN4HY/sY9Tc6H6zCHOL85B
JadTyTgXs+J05wm/Pfe6/9b1AocvW4EV+yyy6Toj6D4ZH52NKQKi4OrsP8OgAoIv
6jaZ3W+5+kUcBHCfG6iA7eX3k+X3X7TSW4fJ8wr0lLjoht539IPLVbN13M9C2Cm9
D23gB5OHBvPUbOZu/BvG1ahYnI/E4Ox2cfgQgpOf55we5/W3TEdrWfSDmrzRGc0K
MO1Bimwq+csbBL72EO5/CwGOd9OZiGzWCA1RH6c1ZVuX2Z+CJK4iUFiq0VttWjj6
J57tdIBmgqzy++/w88Tq+6oJ6CsjEkf+YElc8dOQKVdmPmWELtxCXwxNG2bsBYdA
zlHnwKukv2eLUH1nFicYo8LDYDKm6ZmD1gGaXEaOnqBqDSKN4FNWTponO8cZlIU+
F+GFJOEbbTB8+HnA4d/Jyg+qcx0hxdqzLGy3aN01jTXsxd9aazZpF85B2dOeXTuS
SSiwsx7gUJW4OLtSuouCBcuCZ5iPwrDPNlyyPGin+hNklj3e+oRzGNXq0nqYd9iX
uPCNzNtdV07LFcolQolVto986+39JPlF+mwJueAlQNzM4ORkAMHacHXEe7rU4vui
xGNLTI+i9wmwA58Q1n9i6TTacu3Usk9rXgsKHNOvOBznCb1lBxpLY/wuaELDwX82
FzqwYUs+UsFuFmq/vauWSMBLgaPl1tdEVSXeEKCOcqT6icIr4aScDOKGtaRDsmr9
a6oGxZ/rt26Tr0niohHVvyIqwiBcEAWDAC7QEkgu2pfPE8+lG4HvYUgz6cRF88dH
pyX+Ms9XDnUufdO0LqPbCjy4IbiZH7UGmtx6oBP0aEgOtSD8z1WrzffznAsndv96
4JoWNfnVhiEH/CjvaLhk5mXTg+UIbFDjDkHf+jgX01vG28Rfs4XE9GhZUYuBbWzI
HanOaNuf5WYetwnkHm7j2p40v70R78UGj2JdzcOO64iE3VqwKKq6pPXqjNd68bpf
Me/U2vNBh6Uih2XbhDWCrJl/XX//rAKMcuc8hFR1zyTPP1jad9g9myXSm5+v1xGn
KqRNk0nmndhem2+gvDnj/XawAi/hMpG3x449TR3WRNYg1kfB35H+nF0sybuHnUWR
wgEsv7A/69UrMj8X6ktjVLwCkZtovTvvYjIphckxzbJi+5Zijau3dncUvEAYuGAI
lbbXcM6wSXe7b8ZZYrepZ0+peG+XvBAnCrzsc+TGNNssTeSZksL2skkvLKc6/btZ
kN7i4/pCnaHHsD86juxxMyqycwLgusF9GQAuOSFcJRqiX5IEI8a3LhJX5djcZ/WT
i9fRcaSPGnNrLj3A08R3lY6QaeVtW9WrEtN0svSBk4XpMfrLjjTjZ6EyOG7EoII+
yLf65uA90mO5Qb98qyoH3fZ7J6WlkAnW+B3OhW1gDP5bkWytLhLnh6Jmo/yQIBha
tfKhFsF1xwRJAoowu9QlHDMf3SeuaeXxNOC1K+owcVxHlbAlGmFi0My1t3syM9aI
2OdbwuomXAVIYTHvxpZyvDYpdV9ilETLaXaSw4IW/58md35Q7f+y/00J4h3fTf/s
9NY5xFYfGFuOICYqHrYXn353TzetVhQlHnACKJGxEjvF3rewQ4u78D7WJ0TMM4QZ
Nle6eF5ZLhJtvT7dMagzY2Uv6qQo8mQ22iZUSghVThNTUpC0azgiPh8tfL8gRC5u
sE8HIeMNyyM3CiCdPDrdIqfKZhRdGiogfst9JvlEo3PS1fMijjSKFgFpOErjuyIl
T8gUL9eEJZKmR6acygipeF81mkdwxCOqAXqVsiwzqGIGr5g/nyEV4KDR6lxGbypP
k+TivJABppg8sKAW9LmgiTgKdE4BFMLTP+xEnf9DMoU9lQqif0dz8Jw2Bs70kJci
T48TQM5v2cHJRqGyQr3aLrwNFTPgZCUSNbIKVWCrPbL63PnIk6jQYoifuOc0dKbo
WwiBejgHWTpNHYmvWVFTArM12B41bAS0pDLkVa4eapZbO55fh8J1r67M5JkccNN/
RsoWzpxHJdcgFeykahkFk9Mr6uWsGBPu8GdXaahFryCKSnKe7CnSI4hsHCqwRnHa
AtKdKWyawqpOV7LAlAfokyaAfaze0Bz//mGpko5qjVzsRt1o4htXNgO5eNkCabBR
9TXLKU+zMTXH4DV184eoLd86TD/fu8Sfpn1IpfjXyXoPnrqo9021LmxsY7Gu706V
uJa9ZURERn+qkm7bYv+5XGZar9jJA64TfEEFONLNV9buRWYcAg7SE2Hidy2cwWIE
j5ryqkbg5MDc9fugpwiS5QiaBXPoq2geHtKuTz0mj/YcexE1DrabmwIXLGx1bJFb
u9Q2eUPp/qmJHZ8bO20OeGee9m9cTWv+/3j3n2kcWCFp+E8trKULWIszi0bwSG6K
V+W115gmAVd65xI8OOp08t5B9OMt79eYP5+0EcvjSpINfUzH02M8YlmgCJnpOaY0
vkYuAVOy+omVbLWfZuk/aW1tnQS+sD9mcO+E6rd0u9GmEQC6oe9S5MyvuxfNtPBn
B0UlxwQ2BlPw5iAS8hs1bIyKiCSe96rv8O51QtiOdqUkgs4COCY8/H0HKw9Km4Et
fNP26sVOHO11J+gSGGyc/RhRWvWs4g/1xz5gvl0Re854Sq63gNGcTvsiCxfBH4SH
zlBum+en+etn4jf6R3/pK+R8uXkWeWhxXWEC89VUrz5xVeuzkOoGmGQ4mkFZ7T2C
RmXZIaO53ZmioOGV9hPQJQHPFjSTWoeSRtoY//dRUV78J0htFXVrge+KUjFoMGDj
nZU7NQgJPqnIoCwevbU8vqtiPWjFAxvbdTIX+DfAi20ep5NXqXVUbidx6AjALENO
1/NqkEY6Pb5ZVWJacGqleMwzKv2G5SBhvfK2Ncve1g2EyUN3AUzMrMeEdbHkhGsf
76Aa/xwvJdZ7KxGbbWSCSD14ny9pOrY9xBlntWCPhrkMNzI/FiWfhB3eNeF6N89p
2DRda1AHx3oAKgaOAMkUx2CHc1+y0vCFj5lqA1P3HXEpLnVH/HjZmU4RjNPW6tqj
S9NIeB/ArlgmnGljWsmOkpSVbqkLqT+nWhphz6KfuyFZx4MUWZ1Vj+ebiKS5QabQ
ot/LZ9bLjc1HTLfsrqD/deiRau8+nqLNoUvKw3yZb3Xv9xGwCGDuMkbNUCtrUc9K
6JLxHQ6MeH2hRWeNTCrBDOhHse2Q7OqEWT/rKtmIFOYYSE6PYY3P+kM+yrWeth1b
jU5FL3mWfX343nyzH9iGmpznxxHjIsUr7/hAnR7xETW+EsD/POzNxzTNmQHzE9Gn
sJWd0rQ7KMx+Qq+gueSjwmqsVkD0vYHn6QbfbscTEhDWvZuyHjMAYlVwUMiDUoxy
Y+VMg4/pUo9zZ3HaUNWAgJCKj3HMF1ZaT6Y1VdiAvXHJWDZ+a6o1HsH4J8G/meeE
ENHdKOyk/pTrobe9cavZWEQ6Jgtikmpiopmnmbj0adJJTQbSKTj6E4dHQ2IOmKLS
QiFFpirhRY61FtJsMN2mKuQR/hlGLG0T91Flp6lz9ndX6DZ6WD1nWd7z6JziApjh
MIb1R/ufrHjeVBzoYSDmyX/L9OgNIJ2WOaU+H/MBp0+zd6zrYLQIjghd0NOIrX1D
fwhIcMcN5clwQpVjb4dYBdj1oLARZq3zCzze/Ja4KeiEPBhcpmEQLRBdt4cZlZWH
4n/Z+A1QlZmDJZAf9CpW5Y6cMZfl0HU9mNzVozCOocdMNRN9Dm91wXTlOLk8UiD4
8ar+NDaxF8ByyLMZ1m3Yd/x3Qr6h8Mrc4apue0NTSzk3zhiHmgrRUi46B8I1ovX6
aC2NpIqkzW0/JYxI9zDAZglkg3mt6n29B+xJHnvWOPq7Rb0QyAYQVviF6KUJR8uq
1YrD/FJalCWyEegePyFin3G12Lm5sX3+KKp5dFC0HxU9C8FCCkj0U34X/USgb6vq
7OkGFs5cFN2ZqngDDZOuGI6Fy/DebqUKJbxNeaZgB3HIlZn6Cq2TRNz/m1A7025u
g/5IMEeRNdxUTHeXHBhajzgPGVJqb5/q1fI+UtLy04yLW+/ObRQk9sw3SLL1TIGA
6HUs0NQ5h7RlZdkoVSJFY3x4xr8tRXzwxVb2m5TqvKCVKI/NTsDzvDiS+weWhKFj
3GdrBkhSbj+jwTiY6J6gU3bQkr3oQwdGJT8d6vmVMAFTtXDZ51CpAA6KHofIYEgx
YUKT7LVOnOvKstRGmMvS7cs5xG/1A5omkcUo799mw6fS0opgwLhlk8WQ0jqeBPqm
AMsAgGOmJlN78yKG3HNc0rcKUdu7OXcYZxJIdNIdSQM8C3am3QYxrGZ5BOD319fO
2ScXTySxThO3/u5HxdMZtR+yE4alEn3DFikUVW9nngnZNISqQtd0PCbXneX+hNGI
+LG4sucPDHPIKqEtMgEgEvEmgPHLNoFe3h4m/YEWcWdfjFoR7mqSTFSpk8UVuW2B
xz7S0ot2+9khdbsKqCl0LNxTITrRtWzZACf6cUch7SEfmAztjGtIFxh7WuxSZrZv
Y+4SMWPnceUAr7w32C/JHNgOLhEQjJE3rl2ovRPCpbZH4vCFJtYzeO6fFLipGG3C
hynaZ80EHlLss4aF8ScyT1A0Q5bTqrGtsANdvZJfzwvcPY3P3+ygpILvAmM3HFdd
vZGQXPWnCvgjxTGH6a9GwEqTzouQGVCcWePbcxIEBF2wcraFi8+QXMJ5N+P0cSXF
XZ1lEkfIpIglSeUYa28E+57wu812Nrr7mJfXnTB2YfBVuh3GT7ghmuJCfw7F0VNl
D/1PWaxWZ8AKAPD8DJhyNbFxDm5u54judSAn0ML2RQa6eVb/uUYoLCsVveZJF4JS
FllX9mXvOs5rWK6fLimm8cgYrvTVvMYPIcEXuiBwpjPy3zAiwZn0wxtf653fNeWb
j1i9P46Du7xzjqmlreSTTh4frDUw94HUyJNbA6fHifbI2CB79JPn0tzN1tBzWkEX
KiNvtgRFT9Al0wqrG3yNhQznO+W2NPggNOk39Y0ej+kjgVHIT0Sh38FM+gDd2EVi
rKjP5lD7L/Y+uynr+YHA3EYAVIYhHC6LupJCi4DD5KJPweSy6f41HxFN6Dum50JW
N0Rw6fKPY6PywQ/fbRu5zXKtjGOaWvZgyTgC1YfgMqbN+hh52BB2RxXDy2tW0aeN
KSN/xJx5cZKlPrATj7B8OmYQ+yC5RGs/wn2O615GhoshWzUMx2V7JKObYdNfXlcZ
LSLPyXPUZbVOhCfPwP0ZkA/zjLRjVIi2qqhLCq7b1Ske8ItMSWIkHspejPJ0G5Nw
PYMg4ioS/TIh3R4YxwxAdJMc1whIIyBhpaZ9uyUjugFUImO2cGspsykWjYRPLbg3
WzJW4MM7JxnNlWCa92MGswmf2lIN8FwHiDw/oACo6pzWuKjp8koCi9jS7d2Pwhwl
WvgNBmALpfTQXTybFgXf9jVyub5PGMGLZNm+pmKKlLUVu6Qy/31qMq4vpm0Zf8FG
B6yx518ZJksU3/UfT9A3hfsW/774dPmvGNecmwKhwRw0bPOOXeOn5XZDZv4ivz43
8twIHQFf9/VU2kC9yvlTG/cnbdJe7KxE1RetAOe7jZp/T8RzNyygzNTFxWb69RyH
asfL0RiZqqUGVEHTIYUo5dMYUZHX4a7D3ddn9tc1F7cZZoIcUHVGilEj/sXAMcsQ
zzcH+x8hBKdIS+UF2ct3q+UHxT2Kk9LC6pFewrcfQraPxyno3o8IF0ueVrPWwcq5
OvH7ia5Kjcu+aTlkAFYp1bILBSZipJ76H8lsTML36wuwNZBIx7S06Z2D6swpkYi4
8/qjXZ7RttBhYWwssoag7Vq7uzdm9dndPZT95UtNC1gd0dvfxrBXmv5rbNRFyeUw
GfUroQKLwc44XByYElOF01pcNkYd0WF4DidMFmOsopqV/ygq0xLkAbjG44kEcxGJ
WE70tBQgxhKLdNPOrPCqIvrm4+X0yj4PSV+Yzg09FEbFmK4HfKKB8Ys96qo3Kw1S
Rf/QTnQcz2Sj2wTPNxb0ocTQsh0oF8KysSx9QflYqcAz44dgsh3a8nicyFbtJ/sJ
y1T5oHiIX6Y05KV6THuUrAfeXXSzXmghVfEGpV/oz/ey635rW1kR0+cyX6Fsgylv
y36VuN2npu0vX03XbTuXoNsrtUnu0Wp0KGXztb9zFR5ljJCJdodPJrSp5ZWCc0io
1Y2CPCB8ozdLeo/yYMnFmPrtt84J9vAUYuimJVDFaU0rUZCQBOqS1qlm3JPzExAU
4AE63pA0Bl/5b8PnhMbMONh9Ps+rbi/JaIK4TbeaILnWvK9Ofjr/gmlqLMgGUQ++
r6Ty1zWm62eQLFYdvIOpQq5Q/u071Z6eD44TePcnlLl+6/vEFX0nycYuOmd9x5E/
B7uT5cChpMyZhviE2GTyPF1fI1NoIDKeCK6yIDNM1PzspWof0IdT65l7DTLGMLtK
8SbVs86TBMh4kcAmk8KdapddW6zTAKmw4hH85/iGT3GdhjiVLgxM6VUCMk0I2GpC
XKCOeGQdbckZGUTYhDra0PYpNhh9F7/iQ5c+FFP88sSJz2vB6NJVVRgNU91mBMcr
b/O45L7sNfteNlFCI67E0viJ9slTUUuTqzeFwFL9mn3OipJFewY3i++DQKrT+Kpo
u95GQKyErf8ne6jUO7Hx6D+gEMeUdlvdUJ9D0vH7RsQAVYmOIpLCwfYOrGiXHj+U
gyvmCkW6+uwqXU7WKsck6uqph6l5tJPDdBeuWsIXf6UaYSV9ZcIpCVKlyLE3zWHo
2O6r73PapqsIIBWBZ7MtlcuQpajoj2Axmamutji8CyM3wDBMvYJ8nRL9f515YJFS
CnYHsIVp0BuLxdnP5DIYnN9Z8UqKcFBL4Ym1hEKQJ40knj2fozV4MZ/+7G0mmRJL
dpX58f3SQL4gcNuvfLMi3odqjOPbNjpJ7E4w39OrbNDnjiBCCtG6zaoaAd2r9ELC
OnASg2JI+sZq66oxh9GiOfhEnXyQTo0elT8MC5wTiPGsmwjRw/gdr7Vnz8TWZ0L4
Ttus40PR6H96KS3/4yUpB/M5Qh4Ay4l0OOlvm4n3kWXJREEa8KVFotjR0BHhQ4uG
kY82jGWFRjDNCIsFjxqBq1yWRr7MtjxTS4uyOuf1W1oaYOf1Sd0r66F2PGnKve4K
09KiT7XJ2BhPET9uV/xIHi7/n0oGKRL5MfqmdbnpUjjYJz2/4Km4hd9NH56m/pRL
yK52soE/lUC0zIKdsPOjY2pfO/t7rIi1UqOcLQ6IAlNAVQCZpuRwNk8J1j3T7eCY
2/ygpHeQbl/yPbju5KNtVHB6wqWHO3Uy2KRGqenU3Vn00NfIUY71oiyzYqZBinUd
qUUB7kZIgMBCIhrLUsLaWUcUiLVgR8msYMpsdchzWRIANPL4Oq/Wvz1rvE1DUamb
6UmfccLzsyxohm1U7CWDEr6hYE84VwyHgy/E3x26xvEWPexlKws1t7rIJa7FumMm
a5kimvXkvHG4uNlvEX4oIQZ9NvoEKICExpVoGtMsl/HhZyl5vDyWlanULuekVQAD
O3ir/l3E/VD0g6kuC/QfAQBOuNb3WgPYbzQds7Q8cdQozqLiVeRqGODfg3rkntKE
icnWPMxwqujqfEUCorQXdBHjGZtDaf6sZ1p0qvuK49lf591eCUnNZ3TA1QUrhBPa
FYCnSoH4mHS+XBLg8bkY3yvIAAqx+S857R2ZYydnt6h1nbFxPUPuOEDtjxS8CfnS
zjc0Ko+bR47i60qT8+XYGFL+2IFiZjA/UZBp5a0uYU3Zq+m0Z1eQxEyYVtSGjNBA
1rV2lYzaG+HFE1PAgtkCUxHnYRDHKIe/Nat4Vb2WgChaxn4nDqpR4hjC+78K0CtT
Fro6vLl1OFTipYcVqbhAdjSMqkweJEt/BUfkCCanogG7R2WDIP71nKcKlGA9a2yD
DJfICYn7k4mcPe3WA2FY6J7T+177iV6qEzafPMj16d2k6uQxf1A7l33+/+X9Az7h
s78jyU9IkXPup8Uq4osQrX9EwljfWpcE3epTCYoGNJEjDDeGWYzkbucg6Uy+pSNf
0JGBvSYRHlj/jwmcwCXLpdhezsEft93RdTXpyqD9LvhXTYwrDUOvnRDYOPjQyR2g
QvpKKsnOAIWYeOjNyRQAh+fml/wvw0l8MEmgzTgxlDZm0tp9fVuDEe9H5DvwSM5S
f8qmBR/jywBeF/w38n3yhOwjNi4Gq8w1svRGwb6Ih7J4TNcedeMYyPyxNc1Avjoj
EhD8QMJPnXDPGgBg8p7xvyJtBMm0ORRcTn1LpEUK6XJ0ijlMuDWUTJ7uq0OMzj47
Wudsh3bb5aKKKovKlMtBLWUKvqpLd/BXWqgr1A/XI1Zfm6RwQkmBp1r+toY6Ecu1
ZhwDkLQEl/prk4DUWgSa1Q3v4aPEaAFiIHr0/R5YisCyVkX6VpR3F0bx46N586fj
HeEhv80ttxOlYnvONfinb2VGD0ovoK50FmO3pCEdx50oe0wCch6HoMJ6nlIpt7/Z
Y4bRw3GMe5z7qsbHynfAM9R+Pi8kxOnoivv87DfeLNL9b6VjcC0v0d92Lmpt9GZn
ZFYODPMbjoGdrSgvBIpVw8qjLmEFD75r/H4Afrw/GVyU0kOLKSgPnn3WrKPO82dg
GPHzxAgC/eLhM8iBqtTokR5IcspLiLmvlayCz0gQlDzIZwkicIFtjVfiN5y1eJUH
VI9QpoNd1sDWptRugL9HUxm1pWyzQC93LdmWpCDAfGrHgO91Dp+R8jB1RtgdPjSc
hRY08bxsipXdN/+qrnXWNT1uyMPhYgUA6R44KMaWZifZwAiv0mDtkvdKgPtwKyac
6TGdWIPY6UkL9tssHrOgdo/oZ24Z5N5XEU3DTODnB6m/X5KuT5MDkBUecIqQFAMT
eF4sn3Z/a8gSYVBSRSOxNbCXA5Za89ukKycNwrb5QnzB34YlytfXFVeOIgkC0Rkt
8/6mrprm+W7HbRgDqeCV+kNA6DL5ev3L9cUvJMrqPlYe6ZYkmqDbMTiIUZJrYf6c
z+oSHw/Xth0KNQrVvAX3jZtXkMCnjZPZPA4FYcw0Ksrvcck4vQvDVmyaiyoxOqx9
dYPPEBm7CC31dgedcSzH0rhSU3D6EFUekxKxmVt/g9+2qljZqag31y+GnTYo+rtK
Ta4Y4QwThLqwehNuZiah881uPO5KWXigWwLXr8K+YrL/S8/EB9t7308onYPX0Dwf
OFd63kYT5AWpf11JudFJNErrWXBNk00DV91qDvYs34Qe4ex8Z04F8L8kQ/t3KXH6
52np2BcRFzOrKS/Gk07awkLsjVwkxaosV5ZmYeSZfXT+u4USv6bbAs1qVWMX2thW
Iv+j2pvnzgXBlCGRnPfPD78cyDTP2tRaX3BrvkEevcC6doo4en0IN+7W0dGcyEit
Sx6XThXpmo6FR8YXzc2kBvKKVZeXpypWRhgcV+4WduYgEUXbjJLkQROaFRYF4735
Msrbw9yTb/15I+HS+ONJzF12uXBLbeiPt2dE14IRE03efx4v4YudmPqIfdXoShHo
0eWTP8euRDC37c53Zz9EheK/AYkrMJXERIo32JzRwbcZ7C7ccBaDHe9Dxu7+mBF6
zv8rLlR9fZcpBn8BH+g2taXP8yf7yIoapr4aLBVgPQl96WotKpHlOqaqzwpJHm0T
plXWv5EFC+DuhYSIkMnqWmowmlXxLfGW3gERybDlP6g110emYU7k5i7fZoYprd2o
zLglMMS3zOdcH8PDAMOBKnEY6az1LsIHlx1ve344OJbLvp0q+P5BQL9PuJ6fE1n1
PcT5Rm2iyRLOW51wqM/tTk8Ge5DKpJoQFy0Qkjt1lmJ2DDeJHkvHFHot+DLbh4KE
kAAQCg8LSW/2l4Phwh/FcBiCVtn1cJ78rfoOYiAkEJe2uco+ejHCBRSyEnF+ZQPP
iP7eruZbmqngTPfDmSXouBVUJfAsF7u8kp33Z9CKQjJ5ZB4W0Zf822BDsF/yWr3s
EQMMAlrZa5H1edUxy/d+XCKgo6n+kh6V9prTUlVWNV7uRpfv2JLwSMxJ2Xl0uUkm
yQ70EAxmhkbBQjDFdCsuNM8IlMkYD7uwCg7raN0zn8e57sL36S5aK3hnOtQ1vuRC
fBHT+xXxhuyXJNq8c6VmWTAx1hwdYCT+UN90AGHUbK+AZSM1zscXaFh0mjZV7gc4
nPMGXySKu1U3eAI4enLG8VWyxEyW/wa+R9jBawGnOQG8ulOx38FyS/qjonESRwIs
sVNuqIRzQAc4pikfa/cm6PPmeTJ2/aYXETfO3Hx+fKkNb+wJu/TscjayDHey4AKT
mNaKYjJTafTASb+NydeA/RV0c4mewvR4BlIjyNyehJFWlnSPc3acaAFoyyXkEMas
r5VcJk3IHyDHMi1uvaMuyculbzQvzbVlsV1NB/KL8rvK4x3Awn3qytyTM73ZN7yt
4WBTUUJEx2fxM8nC2U1GBV5BUEMAl/NUsZW7w7xDHP17dbnbJKlKVhkwt97+QixN
66HFM1fq5y5yAOIuZ3CoMV1iRjiV0e2fIje33UPzuUUd3odG59tjTuVecXUsTGrs
peSosy5ItTB7CwI5R6DhbGwDcuZm2rQf0cjgIoNeNwDwsDnNZzpLKoVJWOPHWusj
oFzLj4e3xF8KsvZtur3lOb8+2sfCarVkLsc/MF62+Tfgo2f9LCN0elYaHSor7B1T
LQ3y1vBhG8L+OVaDzhHlE/y3+azEpvC0bKJ8pJRSBUiEhS8G77BetXs2rHaXDhkU
AGO+GsntwdG4pYGeV8FDn3ZErhU/htCvc46y0ZvX69jJ9auvUI7Yn+6xEpJZLHyd
NkBmnF5eykQbut5xCA0fe6oLCshPHWU14PBXwYC5irObWLiSOw+XfKOH/GO0Y6Bn
Nht2iR8BT+4iKYuhnbxlJr/cUWyhh+c3pvKKVbgOE5CArQiFS5g6gLwfay1JTseY
ezQEevOjqH+WTCyaJtoe3J1mpYd3TGua4e5lERuuZ+UrfsS2SEHEzuh69NQV2rr5
7Xa227T4AI87trSHdmZrh7VXD4VV7AupnfbXgNodosNGzRkDRbpLnoeQzSIGzUPF
1rFGlWQDlyYw7r4HKbElIKK1wr62d1Ta7BS1/o4X1AiFWiXjs/W3rOilbNXYs2Dm
VYYHdvck8EB8LGeogH4vbFo8S9Erac4tCqDtXqR+ujA15xvenKUkDKJN1wini1eR
5kbwdeu/7roOdYq3NdbXvKyIJhhvgan3zK/1Dbp/chuJ5B6bjERdJrbcJid7JyyZ
w8+RgR/Ygzb6TBy/iTjvIWLiDjBAjFnJTPNCM3WxOcq3uk/KB6qW3MVvrGXxLut3
8cVBViNvrrCkCPwU5jV4f3y61R05uk+ipkTGX7vjXrKHLEeehZxY+YJ551gdofsp
xyg+Q7mtRNut91TjRdB7RbETX0EV9eUprBPe7yJk5usnFv4BsrkrdU8iAngKsp3T
NKEX+UVWyoO+KOtPiFtSDhVZ5W2y15FiBtTEdslvMQZmkvicKtiFN0Hqt4qJfWWf
xRnz71aIzl70swE/8WxEZMLd0M1Ye9kuPcCSkBb+IaUgRT44gOvw0/KvvhD825JB
Lz/onH8xJc4sp+aHlVWADErcRR1B8jYZ7i/CluP0r1yYfQHbQarB5zCzvGKLEqj2
z12ZLpIiz5ev9oZ2TDYB4c6rVJSlX74TLaccwQKijLHzqj5EqsciPfpexFIG1elw
Bw36538WarKODWJWdVADc2AIN0NyiAnHLzO6q/SMufmDiYpQ8NCOKiylm0Qm2qBa
ObjegpGkob/6jmtVBipTzKE/NrLtA6p34ox0QHRBabv0YDdTr/GOJzIfpEXsPIPc
rOLqIjaTWuArZlyDjsAA38asa+jAG/utzevcRXLrd6evTClIqTicqr9bqTtAomyg
wLsyhi9FF85C9gegaNGRPZWcjZbK9lmK1THH9orNQZ0g4ajABsFcjaoGgjaFzy0H
tziWl6QwOnPBuMQRTaoNPbQUNR98y9j7yn8qyIFh5qxEO5bTDQ10uxfzKvinLWsd
2ehMuM6fDN7fSQxuYG5X3MHszxyIr20hbbieb7hgd/J58SXbYayNDdyw1VWgLEG6
lwga+d/yfopkDApoDyORR0NbzKE7qUHJ1Kjq5Go+tByhyTxksYxIyTCheHQpQWZG
eQ6eBv/YxaVzb2+Nsfn7KDffwYwMx7boGSJSdTiNJdQUPsfXTPjHB6FlEd/nxviA
8BIvttjUHmDP6D10hZaJpAas84FhlPfqFvNh4X5rq2L7b2wkH4RjTrR9B0U27CVz
/ngPJSfl3rD8KZiFRus5OPrfM7tNpGPDLHr/4N3f4kdfW/ZhU5doaB4YIFEfd4lG
l646LwhyTKVS6fAEHfxqzc5nW4mphNE2eh0r0Nbce4Wirx/kPZ4b5/6h97Ftbauu
2LQNzOxoK1iSPPT+WxKBfm/sA34Qvt1ciZt+G8kVW5xbPFcn1gT19KijHyZRV7sB
4zDwzzePZNPbHMTZ9+iVxQ9DAgLGPzjrdt60Rw84Kb10B4M8+pEEUJNUH5jFNd8X
+9ewffRmuF4bGMBs79vInh/oS07F/jEI0AVQ4wD3hOaN5mxyrilplRhZa15ehVt5
y4EPkbZFbQ2QgP5oX3fHfqxvt4avqJEB34FfrgnU7tquwIy15cCWFt4/tT1qTOOA
8dAVrcvzIdN2VNviHmsrKzQVmDhzWHrC5r2+ZcYIrVAZoY0NPgL8xRZS8Bcur/vE
HgBSfhRicd6Uf23nGrCIgUpkOz8D0T22y5z3VRV77XXcmha9qP1vOUbRnuTJ/mE8
yy0VdKEPtNfopyXgqX/KDCWHKAeu1D+geWxWe7bTbxsAGhdkW2EWcNst9aUhOl1u
DK/nCqq5pC+8zDTPvk8jGTVn/xMAqfnScvTm7LQXI4zB81/sify4RJX2SNLK1ZSh
pT7KHOGnt1q+kB4QQjujIbRTzCwJeelve3Kdb+0py+aCfpBbYD2YaERgkccWTOlA
ekaknrtM45ZMWXYoINar7vHCOVPtu4Q6a2m93p7ZfWe7syQAj7azIouVYaYgHOvX
cGk2DFi7Y5ATDmra8Gk3cnPMNIqzCjibZV+mmWbdA7SuKbCRhcXzBoe6beRbJT8B
nB7Eyq8LHpp5DqnY5fRnryfN9ntYSDye5kSoFPejm5C2I3pApF4GZsMOyuRK+GMc
xGRhh+qPstk6yaGqr3clfbcc9BShruNdnMSBoQ3E9UJczi+Pn5+YCf540iYY000z
ROKCIuv05g41KSSpa0XYkXzqTDT+7lPEIa2iXHWN2rob+uf7FXkieoLfj5zDvPTR
mJZJZNC4ZlWbSAvBlekWXrAahPfrcsmkXtwYYmwXuMr6pvOo0UeTX/15SLBnEGe7
gGFLwm3yBZx3fLfee4tPYrkbnFvMv32iOQxAhgzp49dBn4xDYsQdyjiCMUXUx395
38bTI1I2MEMTfDG58epnmordh9Uc1U1x90NdfSuZr4Mv3nMvD1sVYfjHUHZeUALb
UAoaVGGzr1PUbEh12f0A0kJfwO8zXVC+zwA9hO47KLS3IHg+7FVQNyedYub+QA/t
B1+JywRkt54KRxGMpiBDFFZjmYJnvCP7TNO+WPMvy+v2koMO3p3wS8LUuqoxCEuo
RV6yt10oPvaKhBvF8Wz+3p2WRS0Dz6sVjFW+7mgg6dk5uRT+PJDE/QMhMjMm3ZGu
9WJZ+r90sBf0KGxgo5sL72Hlu6XpvBllyfOQHHc4k0Fy9vf9VnSfjNe16gx95hUY
WCZZ+XjccTMWF9lv8vf5uzAI+YFQRKriRwJ3unHbpWGFK2FM66wHkueI2nFICqWs
XaLBAzYiWnARw3Z8/noF/iznz9fVcKSTxxChhTKHTSU+R/ixxxwQEI8N/wJsQEab
BQ5k/ZSsYwdzwkCFH8AAjW7GOkNOdGFGgxAwl92t0lYyJ/m5oLImQFg/Iz8uw6Fk
XKRP4YkZCyHnIa5pO60i8wh/3J/5uT0gYcuy98ZPzgVEaQEDkUdgI8j8ZFrMwLsS
H/EZITLemV0EoA9nvd4f6h81m8wkqQ/oUZDlU1IPP5UCQVbbgnL1K/YvxTQKTBCK
DLXZ1tlPPNsXJ9NfYD3ni4JTv2EAyuSJsRO8hltQJR2Gh5o9PJ28q1Hx0CZoljb5
HQpdzyAbXh8Q3GvwE5O0VS6+27VRksUCzB82BnbatuBZbdAFHHNd8lXvqsp2ITZA
I8JLtBvn03toxbKYlztsz6ztKYR/pB9aI1/5JyVMTcFlJqUVjKzoaE2lR83hz/ZA
ovJQ1rge3eq6+Szh+k7cUWnMB5qe8GO5MoOCoT9AtHIB1q64M2m6J+X1cdCiPsZu
cszFkjDY2lvXnPqMPPcHNDtUuHoI6HUCDHePQThEKZ0d47iWLYtF+fzckzCjErGq
9pptNOvGklXNCZYh+u1ea7nBbiCwMT52DUvZoTY9fph+yTrf5pbNVfcNziDf4zUc
Lw7++cPnAnZIiOEz5OM329JBSf6SNdmBE9f9m6krm9O0Dedw6w6NBzXk4JiaolmE
szDX0PlXRRzZ/spLcFOmRk+jnzne/irgKQxRePyPPldowqE7bw5oBsvRabkNFT5P
DvjO3ZvuIi1suB7FgIsKRfFmfCYv+2hYnJvop6l1lWC7YKp6MajOaXWaIpoluKoG
yf8rUYWq3eEIkcjb65SDwG3Iwjd4n4CI7VKUgLHuNX6Cvt06X7c+efbRqPn6dk1M
c9EGlyxwnViwq+erH5dgGh6+c85zSqwmUPIwQcjX2JYJikSc78Zm4Hghq/lx7oDL
r7tL7/6nP+PqtT8aBjkBta3silcNxGnYxE6ztUoU3v43cXbBKCiVA7bgkCGA25Gb
MvtHXUzZMv6kM0YoJ5zcImXODnqmkl8YWBa098h/arQWSwE1xrGJBNrAuEuBA8zL
mrHJowHoZueG68MKMe3I6SgSgYP+EYCKJTdmipbNbb6SIEm88lIF1v9N9hNGXcKH
KFEHzJxn7d2xLSAXuWpEizNkdN7eAlkxT5lQqre2y4VOI1K2UFaTKEMrEvxrdycg
10yqJqDJjp/nVzfhtYv/LszHatFjnPI8o1gXmiG+spjkR+RM7q/bNPqD2OHnG2ny
zaAnClzqYtFc9cdX8tE14GGneSnfYReDamVMVGpv1vtE4g0ckPaopZ26uvuFt+WT
HgzAikLRoT2EAyaymQEM16A+p+957b/fgJXTzXmmxfgKxJyT11eFpV921aL0vyxb
RAb27Lc1+cZ6NLI6H90xCkrkIaJlAABt7IKCBqCpXGAEKkYk9M/CNrxxqZKCVHKW
jCCSMatrhelzuxhwmQz0so2ORCJwEhFKFZUwCwFQ0M/3fBwk6GwWrH9NvyQfb2fN
VdY+Zey5TfPuzANvBn7jL6kkF9zN/wylxXnW2LVz6CNhvAW+P0oUuVzaW1x4R5IG
gv7JPGB9BdcLVTPGhHxftuHbTNtRYuAStOXzxfJ3Y5lYiCBM2MkIv0xDWGsBHtJm
sxdaqal/lo8lUp7Aoc6pqvDNKFNHD2J4yztRdE9Sq4gkGp/wbd0h/rll1m/I1pho
1Bg5FGlygOsRjbawUCOkexNEFPXTf7QucSaCEmsQEyLJ9Z5Cor0iq8Lokjl1SD2g
7n854WYmvEip7icBT3I8jpbSVt9UcX1s9BJYAri45kT33V5WNTHqdY6/4DMrMEHI
IIwSvZf1wtBodX6hnQC6sXpDqgDz2pf/TjYtwYMlr2hvlCy/e5an0baPLSwCPUml
d7J6o7eA97dWRJileJsLe2+A/+mCL6Vuyg4Pd10RD94DYZ6iExZDNavzFoOgSPVR
pHiqiqWgEyG68D/sNyh+0Gw968ZEpGqBi8m8vjOi55QDGhjqLAapE1eU+enjFjId
rtsxnRfl8CmPuxAfcwkYQ1VxOUEp5rKhozOGCENCvu/chkvtbKfxQEa13g/nYl2S
pPGRii4L65RnFRVwYhmpN4SNCUqcOfqJvnygr8IrGvqjfpLFizVTrOzht0yY3QFD
+awNFvRmqJrms19YIjfJBu8r8M5+562A6yu5k12k0CgnZvrmUcPe2++jriHrYiJb
3+Dftd5s1q+zI1YyHHBwIRilMO83VBJuuT5Jo+doIVK0jFWzc7d+BSIdCBRVepnm
tO97Y4A5ChMHGjy1QOgsNuoeXLcXlfC8Vp3qZkESdSWCbVPkByu+90eZNyoOOCyQ
pvc64z6ETxeF9p+FZSWkZJ4g5QFeUOkxwFaZhwl9dzPO/cwph90UizR2NI7WqHyD
LWu7gBNO6U8M3BZLIjLp6CsygYIW3Pj8Vi6udpWu2X8s+qfb0+XTGKVKY/nbDrab
+U1+e0FArtzErZEXJHBCdgv+phYQheXuMpP6imRy1lTL8OK35x9sLZV/Xuax0bYQ
mY6yJvjOn0jW7ETN/h0uqekqxKPVJP+8x4a2l7EPaKd7ZtDV72oo+Xt+qj/4bDd9
FEwEmUkrX1YdTp/XdKparo4QxyzsPXF2BVuFxLQgRnfQWJAEr5WRSkCnrKfcBh5w
LNO7MTCiaqzc58Dwz2cPMkt9OaEW/c4Gwbbot0b/H+dM8l/flRWqldrClJL8VEVa
gdAJ2MPvTV+0lv6wwPyGmdsLtyewPm15cToaYp6ix9aBwG9+cjSad8KqEof//90C
wrB05iNXsuHjvxwj9ZqXYH8E4Raoj9TgvBkX2TIauOaKU/YzPiTvqekI+v3PxtNy
GhCh+QeZM80OQ3KuNGHGhrF9+hGitLMl1WpFfOYvl2BwN75JmJfrxVbydBcQ4zum
R5g5ta1VTYrD6ztImcOyJii5RWmnzwStQIWet8jy2V470IZMAoRHu8Z19ZH83/R9
U9MepYVuJDwBboT8nxfbMP3ZwjV3KlPlgMbcL7CzvSFs2Jl7N6IcVUMWqtZD4di/
jMOihnh48Z6atJs+0yeebRbWutFtwM1G4ymVQQwM1Gg+pqatHXYyJpAF/22m7Jsg
smkbuP36a7KPPfofB68MMJZHVKx2eszFiocdDm3gxeYtC9dn/KtsHn6Y2xb/mRKS
WKvpob3tcV8YoTjMrm34ayYiZo6me4lYgLoOaI+1TmIJvuXoJCSCglLHzEJTku6B
jE371fAe44xD+M/wJyZAyaCWxsaSik9MN6BCjQZRmfxmd1F+AR0sMoxiuMzyt22T
uLKWutAsI9rZ4NXuJVk9ySqGKzwgVXhvwqu1ltwlYgRCHvKI6BK46MxGHV4wqcB0
51gk5C/GG3S7lWudCJU2z5t3ORpl0+EvbXQYQq0M19XXMSacMUJeZRJJrtXHhXS1
3ch/od2F0HMB6/LQnmje8HKvLq83y2qWO9vo751rUL4cD4Zc8T9xuF0adrTwulWy
gRydd4BxUfz9s4WeC0kfxbOaEXAhPoVr8Cg7dNtP038bwoooKCvTDl8FXLSCwcPK
7594fBbM9/zeAtDrV5L0/7i4jdE5kXAZquaiX0YbI94mG/iuYN1M2HVJckXesCKA
F5FVTSf+sROVkfx7usCbHGeY1702KsFFezsT0ANCsCSlOCha/A7iM2sE/voGKkAa
reu0P+pk624pg/gr10dFmA4XKaKasfZZ9sxaTHvyujoTHepdUL9hzvzFbop4BjK3
pRcxYChSCLqKZU0O038j+/2RgBBqmbjaEHLRdntAEzaro5ahKGj5yEscu3b9fpdb
AYrPcVzywt7YRGQcNx996qLWgAezeO3G73qwiqjuQ7dRJrxOtX26Ygqc3nEkqfwb
hkTyZ4UsvQOgrVm1VDRglvGmFaexOkegQMgzA6brG2+o5GKW391/IxIaBMDDWgaz
3LHkNS2jja4JC+xhmfX9BmppYMF1Z56asBXf3F6LPvNf0YOHtSZzilv7Jr+WoWU4
KzkTs5PnJlfwrrrNO2QPIameIs5WfiRYEYohDb4uqy0SuDqCr/2RLUlEBfIGy1xe
DkIj2jdd3wMmuLHAGQReiLs3zuyfpDp0rhdHW3qSDqkgnAP8RQEnVrg7j8j4P63G
A2qpG/j4ONRlQwTk4PQTtVySMAuEogNiJbj5MekxMiFXevIB2fpBNBQYSVgysTpu
ZDMK3PbZseFvgQADf55/H9/eOt22b7ZLy9bfFyBRch1LQtFUHEAElTNLY8pWaAKf
YbxS3vn5eSvkhrX0W7uCxljv4IMCwylXyDnBf44J/4AexnGQNtRK0n61GTj8vO0/
14fZobZ6LAtVK1kIkYPgU8awgeWv1Nw4PHwq8uShBq+JNjX+A4beqU1YhsBV6ruK
NAPmgajvzhn0ABZTFkF3fwUipiFWpMdsl4F7RiZ5nPc2Q4mpezUnHUvwQV76B2NP
sKWLuj7VNoUxFwKJkquB/7WN+njh0ho99IH+eVbjAyCuiRD5/lWfu4ZjYJB24YZA
Eafa1BJS9MXaYo+ANlJLn3+jenC80OX0XATkeHArrHsXnSRuJPo1MNqRNk+lHs7f
/5awHfnatVv50aTA5AR4hV2MTyLcYRccUyVLjl/nVq/cOEvj3jtXopSG6AQRro/p
LCN6ama4bJ0UvZWiIeOAYx9LLvO+ElxJvNqUq5rSrFO0TnFFajse9OtCPlbclbqL
nPmf1k3EBQokDTxC1mcWkwRdZilmQO65ojQNQpWpfE7jawks7yPszqJgoyXL/pAr
z5hv3KHk9+dQg3AqrA3fK9dW3wKzncdU9LBhDaiR74kDSCOrH7KZMkZR4AWDFlCp
aaQtMXqK0+WkiWeKgQVeKem0dqhK7kMJ6J3p4rxoFrWhVF1uWzhhjuo/WZ3b8E5f
4EVdAnVYALdSsfYrD1HRdJLTkAz6sjIdX9DKc+9BaG2mPV1J26JWMwoLF9Men/LW
kZaOVUwr0CGyNcOb2uzqhPmGmNmWaom+8+vdFw3I0dbQ6jtGqrB4ICzUsOxH6u9J
vlshLMtd+fp/dLKthkssVhpvEc0HPfaTc+UT/oQh8iY8ztxsGODcXI4StODb3G9a
dgo7313DAfOJbQY/gbavnhxvai2HEJW7KXL9w3dJAF91Eqmftei8+KbnHidE8Jsx
F4zO8ExrsY+J+C1irTrqUcKzCVK4F+gCXZl7QK3bd8nz4EAQyb4qwDTyl29rHlxD
W/bjtzNa9oICJxMC2Zxe41pyTDOP8pgfST3ai/BzTbvs86ddYRMjd/9pKKi9jjDz
OwTu9UQXWjENihlXJ4+abL0CF0+PNGgw25kQwY3AOtGJdq1iPHKNYZYKUiMKRdVq
DIRQTrmE1/exfOcelDto8x+sTuAgbFhuGLL4fw2k6jEo1WmGZq/PE7HVPgCHuO95
WzTz76769kBmiRC2QWzh3epao0a2YV3FJlS13wadpTUI37ftN4BWg2Xzku8poh0X
E84YogMOrw3KouJ5YU/wT8HbjsjGm6oYkTzbrlfqcyNh8TfDyolnRY8Q9oQoKu7Z
7/lWLyy4V/fdL8tGVR/K0A1ubBNPQ5o3+P99uwj8Rs4eGffUukOKhm6R6B1vvfqR
DRhORInc41fnKvGhah1i2oc7f2rvtZt6/qeBVUHE+dt8uR1t6Yipx7Iwrl+jgdaQ
Zzq7VYGBiha4Gei4eAjSkCwzETHSguYKDBL5LI0BIfB1KBh+NHYI6DGvm5ot9uBk
tbsPml++S12CQte3PsMlkQmlQQmeHzY/kTlnVvc8v/036kIZBcqUkK83VXFaFplY
zhJragWqokdou5jHdfxUKlKs7ZwewSZYi0TvcoPULjhm2J8p8kYkq7ThczqclAt2
00ymq/qFDTiBmR/eIr5y8Ivu+5P0T5A5Q/HMNp7bp8Lmxca3zfHzKjX3JDJ4MPZa
slDSpB+yXuBgim1zJZl5EK1PSdJxAY96ZyED9NUlvR92Hg5vfeBiZpxDF21+7bN/
U5BoFiCjLeZZE7nWp+gZMjemB+q2Ueglsodba+hPt5qGmcvEPx3B/6O0SOhGSJJ6
0c0gg724UBq6lGjluDTahnaANVauBwWTEoJn47rc61gEySbdAujA/2o5VmAUe6Oo
zJbJk9/wX/OsgIMn8+BsOFyrzoGp6rxdwMH3fv69P4UdpBY+4eSVrFoJUvg2qBGT
pBISqUfxejkUYmMayNLhlWJmVXGrN1/D8UOT1qeDio886+w2Ed8bZoD2NIRAHZ3p
jC6ZL1ob+MakHA3IzyT2xKRTC/8+Qe98CJqwQQZMHCUjn4RkR+TmzXRRt243if/0
fTvCEz4s/3Vv1xDHQmix8mtJqQGxqdW+yYf9+GUD33Kcbfhp6txKh74qDeyBoJdP
ivyjSjPBl6XTrf9pKrhOOJWZ4AqGZ23b9BG4GwIN+a4egCS+Siec3TA6LwryOTyc
/RWN23a8qdOcaezRNy+ad2fy+PkqIKoQhK1SfXQklH7vrMvGpBVRWn04bE8PQabP
9q9HKZA5QzmKAbQNpDDrDVI4+Brrs0i52yVQzD3+dYdSVlFjGLaCyY2+xeIBDhfn
22jdqDh5yk1afXq9lL79eeKkD5HkbRb87ya4ib15lX3aovuiJp5lWuNY9l1kfEIi
2mDjzXVsdpmmfYbBEYweUzwA/2+/TpM9y7WLKCgHfRt/94jMzMtyRp4i9ol9K+RA
HgfpPHTYGYyqcIy6cZVjL71jJ9ckHr1pSxFy2e9qymFQGyy7Rwk/1LSndfVAYhAv
aQTI6xXchZC4fFtNQlUn9txldq9jNonBYvBgeyZzbG8ZENEu1XVIZTBvdYa78/x/
7WRak/2C6AbSXFLZ5chTXbAje3A4ql127QTmhnKnaW1rQsbj0dNFeVxAHMZIf5zK
jZMf+G4SR+M2BABKmtKldWDkEigHOGEAKw/np0ZflXU8/UWcmHiytqa1v21K1TRD
HUKEO1kXKtxZcP1oHXxJbh9V7Uce2jQxtu/2fcxPW3i90txUA9qVqNI3Q17bpOuD
M5GnlwsdmqfAHL5l8V5icunXuXhvkDX97gM0S5cGt7J5c/5qrjH0Ryp1KMfgZ9mH
brMsjfuo7Nq3yswL4MCuV8BgBM1duknFUaBfXNSJicbYzza9aZ6JJb9oNSOaS595
XPlWUpR9p+m36nQMRxs7C7BFxN1mTx+St5Dr7f7Pigx8LrTpizCdHCukfT/lHUNv
Y5DhfnPyYwNN2+rIoZtiQcvBGv0kcM9tkGhM++KhMU4q7KvQwdBDvMS3hnjw45NZ
RZHjwM9lLw5AraOc5IZ+IdnJfXG0d3mGay22HoZw592g2qCyGjS1hx5tCVi8YIm1
K2d+aFQYjLVrRs9K5srMHnw1QdW9JqZkA65Nru556YjHYF06aSHEXSTFOP8AnTqj
3R7wPnnkrMBcwJE9ETCnYAQBsLTyP6k/LUKRGNWuSqxnKXeEJxapq6Yd2fjU/2Zn
7wAqiUfypBDsglKY4w6HlCdKk7S0PlC2B+IYI9jjWyY1GCmm406DV3T/onXSyAnv
jyDtUOIATSZ3ftySgFnKPFvOnTMv+lkXdfJ6+c5m69gK8Q9UGU2Y2Ygjc9hYs9z4
js00aBlekA9AQbHV4cIctOeqKv6heMgrzkxgupN9vD4K/Uays9FxH/BRZGp+OyiE
+54b/La4wQLsYtQp5tt3mCPn/jnLEmuUHJ+6eW+h/efX2ksRcw2uTCErs3+i2mW1
4m3EGgisglzJWCZAa4y5ba1C4HJLrdMHGi2PuO5WWty7zTANEg2muj8vmDM6QpzH
Ej+WBG/Rw8ZvRPSvE4nzr4r+VbhVACc4I1ft3SPDG6g8tHZQVaXwCdxuxN7X3l+b
Mzz8tBVY689QBB+sSTU5a7cgTyYMlStnyMSxm2AZsKp+Lf+TGIAfaKcJ6Q6vxzGD
WsnNBt8ltJ/kTkqjZSB3zUhWys8a5w33/88VfXQp9jLz+5YNVNuNsSWlxwLdN5OC
HasDu5kown6B5d5d9zQdoZIzKmuBx3mONllyH1MeVBJfRH9aDeB56OTpN4ndHZGR
FBDKedUx59H3fz7DWjps/dFAJGXhwOpYKheB2ozlu0u0lq5OQYTc+FhLI2m72Psh
3sLoUDWBE66/gmB2NI6SDHnRaK1qD2k+aVnpNyzWKYX6n5s4wWuzgrLLxyl7BlsQ
Cjwce7jXHs7D9T7EHF8nz4fd+0kiD/4xzG8sgM9ABmpWQCbJsGQ/mBIMAvrvwAhZ
MURyFr452beHc7shlbsb2gN7OT4aZv9dhNNVkdXyl6I/YY1tT5EBggq+Ub7Gtpbh
qfFisB7wd+c9Vc6fxEotLMer9D+0ipDONOkhgdYC6ymn1SH+m9JHuyph21Jlh1yw
wH3RLnqHJ90+fINlyfi7cjV0Yz5S9OgoD50WNGTSzuQwo2eg7T2jo5YZ3nXB4Sbq
cV9a6wDFEQwXP7/aWY0XvyntUYwkrUyLtvgcjo8i5TA+w7lHO502zY1v/qWQ9jQP
NFOu3kEsZpkOynidn+vZ5205oF94na6h6cClyUdli9kf7J5tkg/SmmDazRzNTVwM
DJnQ4AwIFXnox1qFQwUBZrdIkE5AsBUqHhBBHTFlFyUF27/MgrR83KPpNEJWviMq
Bbdi36xghhIN5rJAUOKwPtvBMF7810iDjRfZgcmD0TQgGx2n+6GQ2Ct7IujJgKqP
uS2lNwSKIYDfY08LHKyFxMs5FQT4yr/DmPRWu78J7aJoTKihfkqMe828htF1vZZi
4DzcgxRS2NM5IWcCpqSRm47qx14TQyEX0CToUR8sq216EdvevtPi7zd+VlqPHYUF
mMI0ZbHiERHUsHzRqZpNCEq/UXpRYXUc/hFLkop7bcivs1s/Ow0x2duXVyAY5LwJ
Amxo1Hrz4489BJbqR/1H685DbGU1Wr77b9cIibDsCByKf2kNJHdHWdTy4YSHCKxw
LDcFIP/H0GoTrzJNmxR3A4tuRxHj2Qiqnhn6Zynm/rlaBpfFSsZwg/YKqpCE1VYA
FJMfTq0jtH75G5j6UXDU+DCOjzSAUKOGWRyz5kiuFHVGbBT+BWOv3HBf7u+/GmGb
jFi247F0ko35q5qKKn9m/cGXkFEhe0QoV3XvJrICZ63f0LwVSSPGw9mSQ1uG5rWf
jXwcXmtbNOR+oXh9y/QaZrUVMRNzS/dMII734W69t75tkHrSnwi+yRcMxqaDBJLm
GTcS4GVy2lCJXh/ERrDT5NsTBmfeTeVk4kb2qHCoc+dhg8XTFtOqq2LFHz9wvbSL
HivVd9P4Wvxox594AddVWHwcgcZc63Au7ojNQnr/RMP1JykPgtZ/LQ9V//j7RPsz
F0bVOa6cYo6BUvmvsGjZtJqbQETV+AefHivQKvYvOFevBF0b8iSOuPvPJOp02aTh
wc83fBgarqraTB53Cbqkh2rczI56TLx5X1tfNsrPLip61VMHH1/0115Qi+UdXLY/
y2Eiz6ytCrKC8ry7+ETNy8UFfDi11oJXSl+2jJ+KSZThi8g+TIGhx2quHGjLVwYF
7l9X6A0K4Q1TvNcLjUyf17s1HJ9x1nkRoMIChPSsuAb4Cbyg0Tq/mOK17uU9UICj
gxEE4ELch6J4KisTvlu4x2FAjaQW6iiecMo/UBt3OAaK5Z3l0HXfkXP8bxoi1Qzz
8438pmYQk2N5Cl3HTXSXm+5mkML1TMgz2yo+ImUTgz+0kmPutLOOBE6IIpa1GTRz
Kdb45GRk/4XlpY2SRs48vCcXcWl7Kzhd6/i7JE2BWD6EdiLOJFFi7CWi6RkZdDWM
EW/h9hWe/UA1Sx27mDvkCh3dqbotp+NudezBkUaq+HLD6SotLnPVrAb4o4efv7n1
96is7B+ekMkoxHsFozT4UVBqXLJ3TUV0R8p9PuKJsJ4DGxkWIggvrDgjNRomhoqA
5pRwHT2M6PY4cS8aEcOAwExdPiqW2gmFcYUyI2JUv4Xxeu6DQ6rG5J+M85/bSIPL
expAvKyOhbkzTPVOjRGFy5imkhsyzV7fwqpEb1AV1yl/UJTCoeM29JjayZSN1YZ2
zYx2vCOuoJUr5Tvsm8aP+H4T2FmH9qkvMSq6+gw16nDI1FLVkMHgp/VXHxGSBJzb
StQ0CelVa3BTrw8Pgl0WNDKh3JcvO6ocYJtk/J1gAYi5mabQcjqvuNsjAY4omQim
4XwBv70GyoFAfTL6S025KGueGjDS4z7GYYgqY6qM4wYni1GEFN0pzbHQgmcu5cfY
uhm13cZVM+Ldv3MZOwHpf0LQMkYIOQ7F7RKeutX0K7de4VsgHwjJAp9qdgtZcVpU
ob2/AkWz0Jk5TMOLpJBrx2ml6QjAYNc0q9VHOLQ1aobTpD4+ahzO4QyqGjAkPlSU
w0ZbLfMlTLTLotK/80jEXiz8NyRlCj9VljftT6/oXuslWFkbczCan+29wSDF08gn
cqPLklsuBbg/vqucQApH3H6BKjl25NazAne923ykTNHiw5WLaUMVPAE/acNLII+V
CuVPAu7tXwtKhvkQr6y6J1Za7IyM5bdbS193Uc1iNctroo/RrNv53XPoRyp/MLpy
bVJ5FzPZ+DgarDqWncukBMOFwKkMf4J2q5e1iuPhxFOEkQ+AJxkbDLQG0RPPrpCN
fEGJYpsTEa8p8OrTX/Fq/NdW9JGUBHAwcvD0h+0a6rDl1hszZPXpDXv2zzKk2lTT
K+ky62Ze40j8ood7BAL1udkXJ0BPag2U+ieNXEBK4ECtQGslgKnvBpPGk5AWE9kc
6Rh5+Sc171/bq0GkeRIGHGldeqSG4SAqP8nuOemJZ/rGOGTdxJV+XwyvkBPea80z
DchLIffRg+zRYlyB6wd46p39vN+sNiqlxu/dVxdfgTCOhoxBZ/cBitNaCU6SzplX
olTHmVQU9zgFXaEySRkBCjYlP01HHOhqD6sJTAitds0jrx1QxJ+o7GDgqfReQqpe
wGQ7OQLVWUgKRXcyxKVLCVwZp/kGVWzK7/aGKpQMctmVCDTjq/Qvwx2QnJvSW5h+
ee4cIkwHMTr7BijkHedN5j3bd2U6qWzR284cwL9UkU220EYyewZi1Bx5aUKuseC3
lu4dtgUhyUwIKbve0GfyBpMMG3m+hIO+Qq6XOqhozAkcRtci6KQ6JLyW5pjlVRCK
ds1SzpNElKPDZpNycS8/bAwYxPcMZzweUDnK1Y8YSRdUC6sfBxctItTeLKI+/v4E
a/NhqEktXd3FDJmGyjn+EF3UzGW155Mr3FmClFXYqaRX5tu88kJhi2fN5nE7wZ84
6Q8IM1uaHzGYHBEeuizIiHKT3N3334qwwgPAzbFB0D1GTUMjzu3WNLRuIQEFWkqZ
+RP6osOcYgiEpIbKpwohQeDK11/UBU7HoJu2KtGUvv9gQCB7gL02aYKwTuUe5PQk
bVQbkoiN88Uolt7sAcgrEbxzvmItkJy3h45+jwV5C4GMwSaQgll2GhaeVSy/MTsM
YRD9xkRgi+BMAhILOGogAt9LxgUleOu8cUbZN5AreZXHdt6qNF0qwVA6JGVLRkgw
vLnQ6syL9wlamjzc3CiL5Pm9ZpttAtqtKvJIANfyvoxwHKSAiotiRWmO/X7KP0hG
1OSMY8ehqmTqx35XGiLiS1JHL9FeoejfnFaBX8tY4+eaHY0EOadvhqxh6fo8/a7k
fzsr/SMLgwkvFiau74BzYKwL4t+Z2m/t0TtIzdmVm7N0NtaweK/Sz+cw0WapX5O5
Re+lWlkhnmQqrM2eH+dV8xFWNn9NAb3OEQnaCXjsq/F0UjFUCtsGEEOiHpzxr6HV
VAczEpufqGgIochilBcFft0bqsic8bgj+/39l+948hle524NtV9geObODH7yF/IR
hvnXlE6kmDtK43YgNl1oesLI1DIPmvIkLNJ6DClWJmCu5Tcbb+thPikhcDcCgNOX
LwdwgO0hiaN30iNU/L8VzxAZYmS0jsxy0pfaPTkL8B545FUObFUZzdjKBD13tunf
K/PLTz6BxLuywYVKUN1Ky9Ua/SocAFrqy2+EBwY9F5gEX5JIHpAc+X+cJ/beWfb9
fVC4BGxe3RiP7xs09Et95UB8XbviCln1pr4ob9gnmyfjnU0KoY7JxC1xDSVrOp+z
j4hcbls7T0M6fr0GHV5lzoOWfGQL5YQUL1vvhBnAdPOwdauX03vpZ0/KKJ9KgfBh
FxvCbHoyITIumyrwyxCP1H0vAdhSFmSJHsY1oRjKqywWFizg5QsEWg8xq8njI8AH
vGj/FV/JQTOOSdqFaqWOhUKriLOKCYeRCaIjsmiDof6Il4X1y1aAkRlJ6+rzZRF9
lcwwvAtmZujqbcHB817KVhiAsrk9aX2v4ixpfxSsyLPqwWlhzS461853rh1dlcDw
c7SPbJ0MfGEcLnSs7X15NIKYF05A5X4uGOqdPe3o+cD60bS50RiGU7G0bDuslGUK
xr6Oi4T1usiSvbE3StYtKXHFh+85ezQ+COtg1b+rTtuD4i6weyxxb1kXO8q7iEfU
iIMV8ACuMQ7jz4Mw5l8PRs3cdZY0r2HUgzy0qYYu3+WWpn8Dx4KUrNkmOFfkB1L+
d5gwVZfiBe/3W1bJZqGwjgN58rbjnP4QEsmF39xxcCP5pY8vJgpcseBY3L6V/9uQ
Q+ArJhkUdQLIc7GOEbg0Sf0JkNYYjy2L/TOjpg/Fs7rkYJAstpHJKDQ4xlTiuvdX
BtWXP21GgOMMvt+eh82FlqqK5b1XXGnQyqmTsCuMdSISNvtZ+Y5P8Zq+hwYha/q9
7vOtZm1IF9jgrWo26zN5kA1WYKd9bO6UMOvKrxb7p1Y8nc7yuwRNYCAY4Y5DLMww
prAFninuAiWx9cGbSIMP2VLaLFbSvqWUKOtKjRNHTKzLXLgcVGaXvpjvoi7Cis71
EH5abqrQzdkergNzUY6PtV410SrcsqSvZuVakyU6YKmi83TgiQuSdTv+xzmrsZHz
Wmx8dSyVSebVOB2BlDjW2a4Eqy+PJlt45eSwTeq0nhuN+/qIiB0e7G7injQquxOz
xBPUrtPD/LPnVERWmYLL1E73ibuyZoABsxkH4XaOvW/ezZVnO3jruxrTmx8feXaR
D7DWByOhs9NhkDvU3c6wfq8E0SyaIKyQa9aS8S9nYgP27Na7Sd91xCW0CTvm9uXF
kAUxc5YqCgofp95HlaV1LxcJoZV7FDoaVKBXCPys3HueT5ZwvtK8Qr03kYWWlb7X
u44Z19AuhuPSHZ1dKMMjJ6SW/2f+xZ9mIrT5zYqFKzo0Pm87rP4jGwvNS7DLVYFQ
nZzkqKEtBG6fBVYxYzsw05tAWoTD6fK/rsH2DgszVbG1UovrLzyNg1uRSTegKM5S
dUafojMEHMNGCAxDDsxRVHjBrdat8GhsF7EefuNbgV2+cqRnxEhqCV9J9bKfyf6Z
yyTuOSrZaf6e4c5oNzEj9sp7SVNYM17l+VzRmoOxRhponNk4HGHS70UdB7ZtkkgJ
w+tzGKSgOQN9UqbckdS2A1AH3+Cdt107keJDjuyMWebCJX/YrafECH2QAGLuKhHR
2mNv86FAEeUIR0pr9VRnsHAM23fS0pKPMpbCy9jUm5aNmhNi+wPvb1ka425A8d04
MGpXZmDdNyA+gUBuzANofV/+f795CZGLc+IDGuf4myXltLgBDmtBT+p+ttDsBTcd
K7vqDnX5t2ALkTCxXN/y5m+UxKsxpLeIluC3OQFzGA65/FmcW8LxtWFVPp1x9yfb
zbc1ROfi2SBFAaxr6FcFOjvmeR3HLySTmnF7qjmy4aQP8JwbKJ7zDWI2/qew4XP4
kRU+DoUOuF11h2Uc6Po1x63V0zIr76a3jfE7PT+KfpCwGryJgS9B3BQz9bmEaiVE
f+VOvapH66sEhOMnnWKprcH8+I8fR28LGHF8+dB/aBCQR6+IQRy/T2o9IVqrCP5D
UKe54wZQJfC2jq9F32KOu09Ys9o9rQsR8iGLhy6CkCgY3NTd3F2evmlx3R4Tpyj8
GO0kJlpNxp5ZPJvInUi1IG7bw6vpjZiJLxWkckpKwefi+qXaOaRXjm0sRBW7GX0y
8i0kPWP/JS1wurnvQrykBMF7kWnNTQLBanwgh2gGAw4BE/3kHEJJu8X74w7znwXR
whUPCB+hR4CWir/lfY/nX6FWsK2QeYBL13OEIe+iNgawoFeY1ZGGyLptY9O0f/3u
u2QaQ43ZQBmN4mUfkD8E0A3MmntQ6gFJd6Hn9HuhfXIzjAGH35S19SNVpti8kpPx
JAXr0DEeEjNXNLCmuvtMNlHkwMs5lJsOXUEDp1Wv7tA7sCGns4LODszvlBpkkcob
JQgL6md2s9TTWELu4stc58i+pM0+tDPMkVojRt82uu7Iz+cmHh2taVqrhAvCu4m3
4YPfAlGpkqC2AGHu+KEcv5fvLxiEqAbUlKPCT2CyaA5XNdWNF0Xeeea8op/yDkZ/
QpinmOHF4m+Ps9bF6FSgiE28hOU0tHAnXVtZov/YUqs+/uv+5mI7Cb5AkPhlC5xP
T3qRbPTznn4003YE91MwQj2HJFYxS1mwxlUAN1wre+HEaRiegeskZRCXxQyeoZlI
6qjYUhAxrPSYIEE5ZiLHyBE6Vm1s6LoRmo/HGX0aiwJ+tNAxW0HnIOnwNL2gwYj7
H07FpMBGCqnOMEnNFqxiIibcUiNILDAByyHFnEr19oyjrby6BC9ItUtCP0/CVw3v
/R4ZVo0PhIJDOtJ6sP80jp/Aqd0YFdJfdB2jaBSdEGCIhxQ3G/Hqhhu1tA267ghj
My9K+eow/ulfOnpAMkuRCSoTVy3p2toMgJV6yc9v5YO1urrQRT2Xba8EkaQdREgh
naqFWPQF+paz/3otYqs9qb5qu+nVPdjSAopN1pjXfoV30899y+aauDlkNaN9lalb
K9EVeSylzVsdQ4iYc265G3tlkwkJHqB/6lfkhrVAaSawOIi/J912crqYZRAaQNRf
n4X+220y7TW/MaLD82LQp+r4yFl/II4c/ImRvHldaEzlvu4GJsLtnwXW4DBDkx7U
2CvLFW5X3d+whb87JVn+7q42dh2MCzII01U6WdBmEtI7f4fN2D90LVdmARZL+0vM
Ed/DDGBigBvZudbYy4VxJo1G3lpHDpZ+L/v8oOJhJv/7vz751J+54PaojK79UznW
peZZwFIis8WeV7isedTf5ZfnKvPVsYwEioaQoswC2ZYb/FQ7WqHcVmqP58GG/obg
f0dNEE3GKb7wL/9jzEI0MedzFhmJutkuoxZ1OkLDNeohJk5Wl5SbRBt9cuiWcxTA
b3DLo3Q/xVg/Asx3Si49CluyC2vw9sMLPjnHhZs3Y3X771i+DrHnG5/m4cs9graU
74zNn0PawdoF6LDikHaJSXqDC2slb9E76rLIyRnpE5a1Sqme6IyVuEBV2vIQnK4O
cj4aGOUq/NGZI+G31Kj32q/V2F/nCMSPZf8s/gGQY0nxxkBB4fYDZP2H0QP/gUBO
4+0o964/vFYGnAwudC3z0gdy05/20HREn3F98rLN2mVKG1PFV34F06rKgc8ukzuN
pjG/F6IHEEaWlRxtHy1wIABzjcBoCSBy5zeqnZ/2tzU9V3GLDz63clsPgQa260Ov
Wk7Lapq1SovFTGz8bwoXsxPF/0TdcWLfYU6fZIKq5w+5nzkcfEruYR3NwttenMYV
HoY+QUwCjgQSvwDno7deEd8t+7+4ypLFwhPc8s8KA5EvCxyMisuSZ7WIvVK9eQ6c
eo8JHIyHwvG1kpvYfKfUwS4BywJjYBbPydFQsaIEoXrAIe9PpYgWEbgppVhOysxG
cVul3zKt6sX6tUAYWWpN/BSeLBceGDPkd1oljZP9Lek9LQQbtiVFKYg4o/gxV1mE
cCH1phL1nE/Bfh3iFKHjEUaYi2WMHhnYnoTLQlAbV2P+NLnkPaSEo37aoj09EsEH
GhIXGHNMgn8RWnaPEcVPK+18mQP3u/fObVgBVBeOHSJwAuOoOSskV1LkZcqo8pr6
ZhoxpxYPFsU92VqxaPW4uxM6NXDj99+Tv1nYah5qEBzFYe4uRsyKwpa0xVvrKm04
tk1jiaeBFN6rD7/PZOB/a5ZdPDlI8JQYNg2Elg3EgVohc1dPnwysFgt78rxrGCOM
8TaAcT+nDLCmtHqFXJQFwsaGzpapvJJwd/eDnoiCAXKvqGCN2LN6g/U1RWNTFwLR
tBrWE2HxBJivO7UPi7/Rxy43JBSCkF2sokn69ZMFKfLr/Qxd+Mx47Two7JROvtF4
BasYP60RDYr6EY+8JM7kIvDae8B3pyZ3B2iN6dOVBqqM4aS5BCffSwfH6Bh51tGM
cJLaBvm78fCt+GYnUb04ap6HhGjt9W57FlwAJZHbYzUjPf8R5csj/vsTb4fSfmaN
CzgF1W8KfgbRtLSNtFauIpfb/0kZOiuqRJrGelk4RmC8YlND2eB/KE2DdoD7EfwX
3iwKfteugdZ02z3XzU0GZahXoi5mXfvj7y/HwAVtJVKW6eSiCBTzwskqEdPQKyBl
6DqCucZErirJCNcdrxpmXI5GVKgE7Qi3xpt3OeYISakzUxLLys5E72I67a/h1UEJ
BwTlKBJDsF++mY7jURk5PJ9hW37FMJ1TtNI57Z0sjalVlViixFOqBKyvGMIItQJD
uTCfY5eQkJ7fuQhllA9JWkwW3kMLvdEgZgehiqP0rnAbn/zAbnFudzUS0bVlOzIK
wpNYiBGp610RDEj+nSeRQAEZHi9/WTQsELd+FWG9t2hNIdIcpJOtlSpIpGE6AIkd
AEE2sQzKZedHU4bwLYhTyO00M+V9Nat0+9v3KM48y4qBnfv36tI//yi65XS087i9
mcjNsIvVBYbB9NC5WGzQK2RBgttFD71vNwtoKxJxIxbksC/09+FEkytiiYDmftsD
onZLpDGrxON8PQvl8wyiCAN7BdDXVmygIIfKfFX1l5tZhKa9cotZmpNWJWddLxoz
neg0T69AGmwzOLk93UUP8bqHK8f45zIZsq/jRaODrlcaCazQbnpW/HQgQh6lii9M
Ovr5H2IiKb5WnqdC9ZxGCQ+6TbZSjTZ/8SiwMlYndPHd6NXwD68ak3Xs0iM7mwId
Qq6cvRet68c/sghkYn4DMR0D6ORCByF9WLDxkC7yo/tVihM+H71Ue3BanRvPIx9N
IV/2KgD1XYG6e0gowFFrt7GcQtfoZGYvTpZX4l+2hGzTvsFkKTe5ExxOFW2Wq8iM
y/IepPvQie6Ry7LOnb7kcSquMaXkoKUJunI94FKDxMQ2kjrAjN8jbPD1VLDOxL0y
LfOgTE8ng7+AJa+TbiJmvuc8/0DMGqmsyZXWlnGMxhWL8XuZ/9vpQJYpSHOwp0PL
ck/BqGJGqDVSskXnTP5nbvjPd1dzp54jmJKEE0DsPBTpdGUrKIt9euE4lqZ1C3Ic
H3mpQR9EHyg3P0gM9cNMMvmtEmZcG+yZIFk7oz82RmvxfDDQ0zmvT1LZQCJHHlX9
Dy9w+nX3Gc6/Pix5HElFqL7G80usilHdQ48TBJt3v8gZoVMSehJSIwRAHhMhYTMV
NEcTTWLnurOurCEraKBkzvhd3e6LbuXqduo+gHXAYxxZP6QFX2dnX8kC8vzVowhW
g7tTl5pi2524V68xu6osjTF93F2wojL7QuAzInGeR0uHvlRNTLuWnEFMmCqyjQfc
7vjhL+d/XJwPXnRlzFVBkhJoZkAV574aywoChIVc+8TVts1cV7TPWuSahO55Pn/0
d4xZCepDDSecum9x7mR+b+NMdoSqbl9ABcRrD9qaKCvUpUEaa5vsKT7pKHTdJSSe
OqoiItrTbcTf3cGoYxQCvcaVTo84GlTp2TqdDLq3DGPrc+MP2kgQd7cCrXYVRMTe
Od6L1ZVF404zjdaNRacLvubWqNLcs+oduvmzJzjTil/mIF8xiPnBFiaXSq1/TUpx
7f1vjw6ickMBsL67KzC87J0qtFLKDcw88/HEsa/raIH4GkduW6WIm8Et6XfQxzBO
1+xUSTakfP4lhhZFpAeLGpldbDx5NfusfkZ3lWTZRqu6y/gj/WkCGRJADZXggaur
jrFvtVNpvo0hodxuBYA8IDzW/BISY9gcab1Imqisow0e2Ctse1+nMsCLtx8eLxtn
Ui2ZcWn2AzQT+V1fn1VcPgsSFQTqDe8h77E73en6euNpXMBaROY4AL0XgnY5JNgB
bFuC1faXWlQijP/JGTpLWaTIE1Mc6WtW0UYlaz3DU8Wlf2Zu9LbEdettW3ZWLw4U
1H3u7DrDe8uu5JwbIbOnRzT6mqdrr79e3HB/T/I250Z7stmN9LYa/3t6/6t1GJ1s
asCKN52NymP8VLGNnTjgsCp0X7xHS4EDMwwRTGvuZ9uTAYh97ParwpFfybwwsCB1
FeRc8Zcuit77j0oXd+fyEQsQ5E9y2/qRYFikkexJ0EMNWVT308fkh0Zk41VYh2Eh
ejk/oByG+HmZuwkSk1KNbELDmRy7vZbMrGbyyrAGva4LfctdhpNq9fRrRi3yHiZB
NLUeQ5Tz1Avm+Hgl0EFkbWL0SPQzI17sxQvP1Xlqdz/AFzHsz3IP0KvbykjhnraA
r6Jbu958Vm3eM0mDaDTmsTcpWV4/HUSz/fv73f3qL9NWjx6LNHootPLFoOuZ0Spl
/TNG1MyAK+HOZrz7yhfeWwtuESMqSlFpje1I/9Kt9rNFie5LuVKb9y3JGT01HHXB
hIL5g2iCwHy1N0PFtulWSE6F10h7LOn0kxl+50CL37h6W91TiR7M8IbDxG6T4nkS
bWyAjuz7V5sNrOxlNIwu5l/WI5uXryhJeywNp2iRs8y1pjDUBuYyirPy7wJt3Th4
pxHPijnlHQtRUK/FZVIMfr87UU203AiLU8jeSY8wenPYIcChv1SmLDVNGFFKPcST
KGYZH8UjE0f24OWzil5r/JTBiwMvc/40WF+B+ojYhW8Win9VefyWOCRPgLeKfDwP
RsdL0ftzR515sYRGFHRZqUUZbfanff194IGLm4Ghhz0lVlcNtUfoDtahj64eZE/O
SBEC+lai2Hs2puMbr6wxawTjlV2n5l0egKu/+NX+RT2phMD/n9RVcjxO5jQKMnIN
itN0pNKAZcDdVUYNvgZvdu/qWbb2asUEfPbm5CQrWMAK6B0ZRiANA8kssLlNKK9f
mwXAJwisGnxlDSJx3NHpnr/PbHI/bETIxRLH9MdFyBeVWKWWpZfQkU6X3kAkN6dM
VoQBmnfiwWgssjns91Cv5FrPq2LoKQTX58AkSOIE522YyLET0Va+YWrS4TAIGtbu
x1nbyU9MBdHR6nbyMmijtL9bDhSzDxd/L7iQ95ZNfjuRbDzLHK0RJxfXzXSdeo9Y
tUKRPT+V5qAuSSa++fIxxwmhBYDMzslXp4niNxsl/fE0ek/b5XzpY+kFEBneYqKr
HyXKiQmgYw6gGspIOoAOpHI5q3WDyn9oGpmfH+qFcbDAoOTmfRwWJS3sZhzPoFS+
3DrKuB4ZBtj+QSeccEfZsKcXIJGhC4n33ap027TjxeN62JpnniNjn6+aGw4wWuj4
yMgF2JAm54gUKjuvQTw86R+NMb1G/lVab4c86znHjrHgxsdVG51eUGKtEd+FqSdl
dYzRqpZtpnqwhO5DLzjp8B4RShLKTT4eyONAF0Dq9v0dzTJridc9F+CgubWbghRu
rcRxQUTqqeJTkRNqL3mLP3eJQ77GEu8nWC1uCLVA4slxK5ImhoaN0QafTmh5c+gM
nXO3MZrVvR03mmwtDBdWsBrtQDCmTPpa/eJ67EcrflnxJ2Cj/nKS7nSJDUMIlHb4
uWCMDJ1HyDRcB7MGjlYOzftXBjz2wToBYnlGVGRRDlc02P8i0+LJQI9uDowKEI4r
/92jsxPYXf311e8ExnmsDjbEW58IGyROm7k5/dwV9V51089Z9K3DzAuegSSL2ke9
Ln8JjOrzF/w/m3FpwRt8Ho6UyeVJ1xVYT+117VsIRsMdAfY3HcZ7NJrXjfv1pqkP
bokYPaPgWRIWsp6jm0J3Ybyc3QxeJDWKjdVKx3lAY3YHC1Ls1Y6b79Uu9vjftX+p
RFcUxWeM+DOqFZzqRZgZDPI1AXK5kijxLSGnDrNi1HRT3orwyjd5nnm7/JqMrmIr
8m7DEaSkOw1Hn2C1ub7rMKRCpgaQJLz4TwB8OholaknXYnX782cHt4NjRBNMCk+c
HWRKHoaiSFohQemt1VMWaw51sZWlumgOxd/NRrJQiq+gOPia17gu64JBFNSEzhao
lZGjYvcKcxgogCgfDo0SS0O9ofmNxsobr3HFGDKec2cNUdUhPXxJgoaP+BcL9vtu
mspN+vRAZ4x1oGw8hxOiTaMapH7FRPYWfbHA9IUcMnf+lwLLZKUcIwo+rtoCRwWv
niapvm9IpCi8hoiLKu5ebsXv4Sp6NktgoAbDVJnCytaOR6yonooUiKwfQ3xfbXPj
I8zP8AEZS9mueNJOg1gtuV9uEjWAwKFi1skyLMvfsYgiYYakig/fOgFeM6PbmYSk
2ZWvZUKlQFzbSGFEPZRNluz/kFNLfP85HjY5DTsbORpX7naxzn/S6Ft5pA6hJfUm
LGwGNfYZU3EiJ1NjP4L9oTHMgjuBkFgy5O1nXvq3o6gDDsEV+ywpAY6sQ+xdOSdy
ETNzdmm5LbQCbkkvFhfoaeJqkUE7ZFelyc22iND9SgxpFyf0fU/v/SWa3J8hjOGl
u44fu592hkGCge2tkX7toDHggof6JhwYyafcd6bj/wqhzlCxk71n8mq+oE0X+aKe
zQERUnPUpSMgeLQvVU+cTaS5VpmdI+cAiAfmlJEvSTXsBbVXPWnp4joGFtUvoPrY
EICEeQpPp/eueOHUcVgTRsDiyLBkM/niDbmMqSFG0YPmDhlFBSCx4Zcq7DteS/AB
VzgTN4HeXGhC8dz7z2wOSdpL9R4MM3ghgvNUZ2unWInFEuMNbh+YJpf8wvXZ7e7l
rQa8Vbakn4ni4IeEqP3LeE+EqdzypqChzl7KEe21H0OmMWkSiAyls6aoMr0Izkgq
BYvktYBJ38UdtEIfVncwJlsX6UvjC9e4l1A177xtbYPorEwsa0fY9g3Ex5xuSQJ7
9zkC+iYjAndwi3pFRFZ4hbXnbVjrHzEZ7L5DbDlhjfl5SVYJJt1bJk3EGEnNjnWm
ANlhOMvQ0RI61oTX9F55N+g0nCV8FYziA/6lbsGexKmtlYzUOsgREIgJGQxFgMNW
eZbtfy23yja09ys+vqGWDd+IaGGTh/kL2DcDgvSpJB2lZEo7mQD/D0x9jKSu72P/
C3WDytBnM5oj2Z9XNinlIv3vn4tDW7S2d0AvvKQwcb7rP5CXmeKbHYAiR0g9nB7c
ApPEcZ3SJF6BIt4dbgoIk47V5ceyKEZ+G4Co2iJUGFcvM/FfJJd9KmKtF8QDrq2M
CUTh30PtnLL3XtKNRoYC4NtjP6Vqi0Z9GhApBkWgvMbeSL+WrdrPQ/t6AG665rhv
lNO2w/MK1FBcI4cYYlkDTCW3tObuFjqtmm+r+727Xyx7ZnDN2sOP2NyDqMRIjOJ4
3SzkTJ6fk9OQd0fUdYBPilagdCrAUAq5Cf9Ww8eWoi9eMNFH3+E0VcVQZQBefc7A
ZmLybcKNhGY14Q751VDi6pvKCbsOM74/PppritwT+ImXu2fpN4xOaaBW7bE72uob
Nn5JortvLTYV0bumWsOxxpJrF4BhEhyQMqVD2U88oU3BeEsXnXax9y77yPR16Bg0
jrprUkYqjZJLC85zd4sPebcZ4y0p4SAloMJ1QQIyibmZFJdH/Stnb4YdTwTYnWJn
eTBsEA/9+YSpsEGINhapN/GFWfjSYMQfUMEb8t1thqPeaOJ6h6FuPusYlhljn71y
xCBYaWGHkEjnm8/7X1DXtdEMKkGONk6isaQyjkdesV5H/VVJhtcm2aci/eSAyp0O
fv7M6mqsjskZWpTc0575nwuEyn4mqy8JSIMaYQ1dI0mF590o6ddKbIrcc+oxTOrp
W2yYmqAbf7QabsSuFoFVuOuSLnW3Nb2LGMcyHL04BSJ5H5AXCE8WCDi8zjnES+Cg
JHTXdQq/h9vD3PU13Puok8fRZU4xMgHDRrPPcgPcpjKbVLvWMpF+ipR9mbZGJmvV
tB/BG5joesCFmapykHXDvup6jhRoN4a0t5n4YhUQ+ua7nlHMPEtY+kC3Jk2mYZri
UZdVIby9KbcqftJXibCh9XKLqzBUopCxzNXG1APpw7ff9CyjxpLYGD53aag5G8l0
6QfL9ia83v7czDNMDbttmkV6eXRRXZwtcqWnGEMpFt2SLIklth/12ouOTmPri72z
X7A7mZbPcN0qdZZ0+mNMCHQIX9D1WMVNBVgSFF1k6C71DKGsZZO3da7BUC8S300e
sZm/ulxleRGjSk0n145i7tmGR8ohHeVHjHVtNhWGXhKfpHx1rW7n3iXY8z0+FI1h
MDJlMnbu1g9v2XvMb7JqjRuvvQ9aoo+NmTYYXXLlQSJvqDbpX41hxlhn/O6+Bfsx
22XWlbudMhp9lKDtr/V0hSfasWzRNiru8M2LxYXIEPWM0+LwwrgaZ2uOh6hMkqy3
S46naCd59x7ZrYeIT6Zwy+VvC9Mar1HP1EfIjVBQ9gxHzMctql8quFKgN3InmTNg
Vj+3LTDaPNftgkkKLBb3enZ01+LppmZL3drywCyrFaC+tfkGlOWxo7ghPLhpbpmR
QJX9EeAJlT5xCBWSVMANZt2/BjdW3uzqAs0q/PIqB8lTXIQeFYK/Sq6m90RPFoT+
F8UtBYesjIZ3iHU5Wqel7qQLnrvqRdKpART4EOOhtAO2q9veJeTTHOKzEFBHjeWj
80CN7fMfz5m4K7anwgqeQvnkvaOgFi1MFHXFhyocNDW1iCyDyNqYP+LxLJzAmmVY
+VnaJWiWG5dXg09cIdY+Bw0mMWIoVyGYFE7WQpxUGq2O/+I25s1TdzMftJxF/BhU
cZLFLVMwJBCcF4Av7Q0v8iZsnO0jGzc590RNSqIhSNUbC33qgA44cF/OqKynTekU
O/PJpiRjjOTSSgHdSDw2aghjOmiChNcNKqdFxjnFCBcus8lZJMHXVI64dMGllnZE
N7xbpAMYv9weHwsO++33uPAkC2aJxunQdkUzyBo7cffciGV4e4SHS+i4BGliK6Bi
/WRWngEwlXflk9QxV4uN0ckcHIllgDbltVnU5e7i264BGxcZJ0l45n16gaW0ok/L
cxLzZMtvUeMiWYWln0SV4HeCnQGqCbTXGneJVb0BIkTGIhxJesJf3bVdmm+kIfKb
vFOrOf4WlbEyQYWomHcNqW3I1zkAHlMOcnh5D5vi2aXKszZJzzQgEaEOCGITbUQ4
u4vbvkBcXJVuj6pZFPnY99jjg+SbGZlt0d21CAVoV61UggS6xilYF3DlnVQ1a/pZ
7ob2JbT+CAMNBr0J2g143azN1z6o7+CbneXbnWbx0QbAVTCuFTkc1WYVkJELflo5
ZVFep+1TU5FowiCgXJ0WP9kjJVWsqL+n5JLKwJg5Dy6BWuJfoL1tp0V0YZVK5iZb
etM88piFtPW9qR3sGrpPzIainNcSdy4wX0q8iwlCura32g2lIPod202Pm6ZbvYcP
ImHFrNYPGcKN5Lvtqz53iD1aore33x3d3uDdV7DUCyTkasEp2v9poG4Weyw7e3L5
HDboeJSZQMFWTFBSmUH3okPXiHeiQu0JJXxHP4H7ZEZ16HPcTjwFinqMN/KhnSH5
Jqgk61sw43IcUJyz7TUsatwz1gn5Vr+rS+hEBLoyALgri0kixYAmiUyD8fjt6Vy3
i3L+13dXLuXx3Ok9ee4W/wo3brMbyqHunEF/eyxrNrlB6lqUn0uNAcziL3J5sqQ7
1BcHX0c93GqBTdA/nrEC+t5XGQUL7wkcB16/tBFpcjqJazlMzPjNmIDRlGMHbFRQ
zGd30vAMSn4DUhRmVDq/qYhwN23l9REqKA0BvOAo7ptqbeclD2K1x3LT8thdqrln
Rl7vcF/3NrJo5j1J72v/Cyj42QVKYML7m8i5NrpG1lFrxZontzIuqMRYVBa35Szp
De0DHkFlKMLrLqzX3dbaE5k8nPF8oXd9kALlMtcBMCfhKIau5Q8F5+o1M65F4sPw
kaUT2vBB7LFO/zAOmCdpOSu7t1qgdE28LjITuhefdCyQ4QTOBfD1+bNSsRdCCITr
OYbJ4+6Jz5TihbUDIp4KL8eW3q8B7VdQZcsGA+tSC8DOnaOYC9EDVDDJd6cvtCus
nxmw63YZi8k7NXvr3r7ef5D146US3wpwko9IttH+ua6BcGrnSo5YGBgvDQOnT0ug
Wxl3dFCCxLK67oyhtrafxcXKW7VTvkrdehcLnvruP6K3hPWwS/aGzJmoT7qfAxcN
Itm+9IJBBolXPzZGX0PtNk5RlHajQtzNfTJ/wa6S5YjKNU5RPowI/tmMkJemqwK2
ox6qyFWL0iYSoxb3aKThHVV1Vm9ZENWFQ+zCT9sh7aCVxcYDyMfIr/niI4XVHv3D
PKA8GJJFEujmtvrRElDis+q2wwXiw+YjnjTZA/eKkO/mz31ttRfsqO1hNItMwzod
WVO9mtHs+zt+xXKo+EaAaNLa9XFnySTWLLk9EABJzfwWJHGu/DDjxTQvIxA48kHu
FefHKiHJ6z5keJXF1I7V1CLdTu7EKjbitoyxnzlM2+h3AUkkvuGXElnM/6ZDO+kX
msk6aJhe7tkjvbiSokCmc3+MrMcYyEEVSt1I8CFZLGssF8awDOVS9YudRfOEgCHz
HcxE635/PCdIK2nuIZT8mpk/PHFxr1Aw8dIgJRp8K+jgKEQZcApWJnEsKFpwWAoc
KGnoBdGavNQjINXNhKX1aUvj1U7KwKmJ9bsknsw2by/tgIvsulAx+kL9mM0pcXJP
UsaGjZx4Yee4i+ubJhfTNgakL9Cd136rvQ8LtWM4HWrxRa99TnwX5g0FsGaYPZ/a
qm2XcPH8fg7RMAsUcaD5qFbkoQV7LU6m8GFAJrQBFLYS/iQtP41sYWPVBEo2Z/qS
O2Uodh8ZHqS/IGSJEYBqaYtAixE9vOf8TX45DsXKMYzviJH0vKjwLGzsZ6O3OkKo
bR9X9Rh3z0/TQ4e+4/rLpgNxZfjtAGD6FEaN0h51cD2VD42Qnf3JpI1c1Bx1y4Qv
UkjegNkE5EY8MEdvkO9PcJbIj9mKYhC/nu3D+pGqtBWtOWV6uHD5q4+q//uj+WmA
/et7NrUUh3e8G5SJSBzVmzUr59buUlRRDqDpNbzqcyx+YmDmZOuGJQF0+NRdZz3H
nTLMFMewP0Ts4/3QPuWQdnh3zSOhTsIG+jhl3FsHjsD3hKksuxPmZ8d0k+7rTNHG
Y8GfaSGr9p/2hTo4a4t50VYkmM8URW3yKQt60KN9o3CdWbO+8T/BPPleNpi5jC8B
Fce0FLsit5WU1RBPiv94y9oMp6UDC7O4cNfWZjiEpMGNqcGcFkeWcfKx08CwifXa
+UNvsO66gWub6KTdTZCcOkZ3UODbhRQbKJsQaiRJI1Uo59XyYY3HDG+jPqQUYHe+
q42IOnwxqNDLwchGxe0FiyZLUI+1Z4pAmK63WxJw41Uf4QkIAr1oopP3MvOaGP5i
YalnvWU15kBKhwQILy12eTHhzRRqmLmp4PkEdseziNdLk0vT7vG8h7wRbLCadH2w
4YlZZyAKhJndIm2bUQUeZhMlxbJ8vy1Oq/GKvpahlEQYO/LOCrTBPHph+f+aPlZh
acsG0+ktxm73Vd79s9FoEa2lGSX+Fhc2Dn5PF36DUKkDcap/zWotciKcxLbzQvut
9M+A6pCEV6CV/L3wYrWiHHywK0AX+TVSy/bN/X/dc5HaZo+EjcKDR1gLKWG/UPTA
tjkAvq8R1DYHFCmLGoRkn6dFh3+Ew1nV9fSTl+Lj/jtrdFmi253xgoZa5kvJoNxS
rk+pVUYukliFFTpUov1JCyB+fOiRlYdwmFpPPY6uUILxjve3fetO1VQJrQQPGbTH
Ts/FmJyYffMs7Foi+Ny6VuxpaZDdIwFRqISVS+WC2e0IRY8fHwwVfe16oPxmxHs9
X5LOmCgGItgRz5EWMKYiJswkNG+KOeueNiqEq7cNE80mNtbZ/zj5EVYL3Psud8Lh
OOEr9Uq1ThYCc6+OLZoKun0m2/+VgdyzW1xsBomE2L7klsHzNXGmHqAiKBhysXxU
V1HWSbFOC5SnsRdqrYCQ2EI9OkDyDN1VUsLo8db9ircfxGIL3NgwHRu75AwsGIzT
ONnkFbb0HWnH29LR9YUWLMDcEcGBTPQJd84DCWuocwBHtMW3m+gyJeWkrYQpbV4s
F9zLaXxl9HqzCP+2dG/3JrXUHytMxJkoizOR3KQHT6dXDpnQ7HtmXrlb5cB22M8Y
6C0Kk04fHwGXcH+Y6IZTbwgZOr3j6Pg8mvAGhUnEpkJCe9249RDOYII/IfJux+Sn
bbw0UXdqbPdjR9QQtX+LlwE37cBU2i3iB++X/2C9eD2raCq9NreN4DA1v8Ev+vEr
CY3ddIJ56wmZsji2+zdZROO0ezuheVhBbZBkgWqajwOg9IKuoJVhhnsutY9VHNDr
xTdsUAaM0vOY+BMv9OE+/iCXr/keORzEtkSJaH41QWojGl2rBZ0eWPIf5epgrU7o
pyYhGTVNL4mXls7R7EUX+VGSsuCgsPZ1v1XiwJTV3WQ1Yn85B2OmDPp4kxw0Men1
ehRzJJDuXRTY76ugkVOozVzJtfvHrn+PpDIZ1SP1wR0kADAZYKWlRhkWdOP8p3Ls
Dp65+nSIx2UztnmD724mkhaE8XGS89jhYl0LsKFLULHfF4yXClY0YHdXrleAFC1P
DNfQP0ojPnTBP4jPpArBYJ2DfITHuN7143cVKD7ltaNb4K5ilNH7j/8IwTXkEDNs
sf2Sg7rKGfvz//Ayj6r1OlGd2n1hNhSK++CiydQklP71wENV+Z8lop9DGnkGwVZ5
yBSiyVlj5/Y6lueHJr1LEAxPdadya1CCL3BMwS1LhyblDxrTbSA2G9GPiXgb9dJ0
S9y+isf9+v7G0S0YMCaZVcqlgLLslZ9/9OdwfgU070iBpA90erxG8Nl5V/MSWzZM
TZ85bbf7Jsn2KsgyLJ93BLkIwMTqExkdRYsZbmRGGhYbMtAtdEeyXEbcwISHeuys
qV5kQD1C+eN+WU31nQmEVgY3c9LEBqN/WBiFsm8v1lSzsQTwUOzSk+xy99gzA2Bz
CEDQg9egk54dgxqEnucTLE+i5ulac4d3wpEyQIabEzmBoYpTrxj070+5KD9U8nAx
PaEBmSKYh1Dz0u4JCdDdPmaMG36pKNG52dUmWx4nMgx0X4JL9pbUUonYtgY0tfYz
P9Jb93YIiu1u8tGtCZEyaqpaMvcIPg7L3YHyveKxCEx8g53IRwRnD+qYjxclgkYC
2BR978ORWIgWcE3B7FzmpQs+aVMnU5+exjvkhd7Undz6AMdPHnb6i+HU1EhRnYzM
YuDHBr+dt5VwZHL4aSct14NxBMLfJf9pBJ0B/YtRaebJphVHMU1BFfEM/wTp6Dka
MZ6PorGApi3lQO5O+OG3D6YgqnsonuFXGFgCZHl0VPLqAh2KkDtlID1QBaCD54b9
Oo2fxA6iOEWNSbsSPm9+ZDITa8Izd2ipPHpXt/t4MAzRKwT/T/M8v2dUBYkkAhXl
qPwyqk+RYcSnTH+86k/6l4rRHLC2tQ+5qvJmnMKbtknDRrilKhBRLQs7rVF11RW1
ijOjNZ3CvWBfzjxTSejBV3rY2nLM7ZlaY5L/gGgKrQJFW7NkX4p+AUeM1nP3bAsZ
bAS3kqrbmDiWatz/jQYu+81ptJXo+W2d2jkXe+494nHk9E6gNTbvA+AkX7l0SdUX
2boTIjO8fZp7li0oMsvOAuY2XDveV3uaLJSrzTjNp5PawSa9XvId2pGWrRtJ4K+b
/te2xfqzwDeynb5UzNcQ02QRHqwwA3FjeYFBrwg9Z7enGL0GJnKcixbeAdWkwgD4
7wXYR8Wchcr5s5NpOLUWQ00CAyLo0IhwcfxFBzgDspEggPnueYc1IDI3MsdkZNPE
3IIFIFEp0fUMKpF7tEh0u15ZHOW92E0vdwnLDbF8m5RhWc9J80eIdhNFbcqKPguS
8/235aZwtUunPUHCIwb9yqZihYHYq7KuQFN4CvN6JOg2ICY5Eck0tpY1ORvA/eSZ
mIGN/9FN0EuIw4TzF7pW9Rw5OaZfxV3Sn3oXh0XmE9TJO96Q4IjRIL1mvvUrQTac
Fvd5J/Bu9ts+0F8poDGWJDpnnzTfbDukUA5JYkqiqSaOlPJ2+k303FwufKh0ACMr
AfLCAmmz8/zrkZy+/6keooDfaIHKZplmpv0pIynZhvSOmWYvnoNRUinPFvq4Cb9z
7IDYoRTTrGc3fh1kWbwc1aKYT9BrWy5vc+uEwedg5fCdDPMG8pe2j7JzEJuB/ilJ
a8lnW9cKlV8JAf/V9RaW1l3uxkCXg1qNhtCIP8gg4YWfPQkXHLrbhyXirvsglNaU
T/yQT9Hvjv3S9QMaf9WRlfYqlGnz4pwh+OOUWEXJSYd9d5FLv5PpNDygOfPAHLZ0
K+JJxR8+NK7X1Qk90cRDnI/Uxk4AbBRb8BSDEyYXGZQ0tpashtn8f8PCVsIMWPOT
PscsDmGT/oL5GYxzPVUptMwwAgw49I/W/avgalbRHRkvhOzfYfjlZFi+veA0Lz9P
adZB8039vkI4iBhLlio3mfkvs+S97vEn6Ml5FPDMVkl4MV5FvDCaDBMG1A/X9mEn
Vh6opAxZUohnR4TN8s/T7ATRMmZCLKi7qFqa9y5cxSHlLSeCnvIqqVRBKQdr+Lsc
OdmUBrFD7rpbvN7CAyBsQTcZo3+GvPOQ1OZVzVG/rkLI4Lb2+JtpS2zgamJOfdgl
MEJK0XfcRDVRO2DGcDWnS4SFwD405CkKpxw4dvxjrjhtpin/ormk6sfeYLdJOBAy
dry+5GictJPM5cTFKx9F+PsseGsdAgQ+FYUcV4CHLG5ZgkxaZcSrdXzzPsxhpoXa
3eL8lp1fGAt2p6GXHLVMYlIma4znuR3fMD4Hc9rKcK2mRTclwboBIXWw4bnmsE6a
ROhudh6VJTrRi9U4khhKEKkWcr6sxSuIzxz0hFAESFEIG/B3Umu+BIbP3EYOr38X
CkYMUeUatHL2prAYTk1MaAmGv7d6pg/0V87MMmjCrM/GK72CBMxqcbBsUmg6YQD+
0uulTySG/sclcWt9hh3ZAj8EsiJc4UFjINxuvPxQWFJyZL1xFDMZ0+qY4k4nk17I
g8Xyajz1kDou+xqiPbVhY1XggFRzV71bd0diJAg9KbUJ4ny5KXrBm4WR+6oejfWa
eyg8/SMC6REqi+DV4xDwc52c1XeJLXJOdbMs6+rlvBY5j0Wq2njhypWBJDAQKDn6
mdrSz0WcPGZw8WT7WQIhPz2nsHekt/8juRw7txAZQ0P/Ro6ak/msjog8xBxsH8pC
d5oJacVB9P/KrtEYUq5uRJkN41l0nzWyW4SxmI2/cSn6XSC7VrWmwgOjD8DF+yUw
6I5/LI3nlp8uOmw9AgFmDEkPodr5zn3McNuHSQDha7RX08qbxEkKl2ISwYMxuZXk
dV/v4RRk7E1O+5sVlJZ6cOA34chQNW2Mcbky8LRFlElnHsDOPrPvmfIzBRyevySu
aVsrQ78tY/rzZUmvJsjjkfQ5TExWLXgugHhhqLeaeyOUSOsVt28AulY+ZGm01I5b
0Gn5K3oW2wxkG3vRlVb6KuaFpWQCjapNgBphB4+NkvJ9nCco2omjT0QqvFaIyOt1
Ly8htkOlMWX8UlnZoXzz7cYByNOjxqznOFC5DfgcJ6entTOAGRNOZuXSO17qfFXf
KJx9IasB0/gL5AApmTZwDpq2FE6WSqOexDfkTKJb0Ceil3wZtTFOQY574s8Qzmo1
cvynuYS01xKKDZdYxK/Gd2hWLnCXNFEQHUTp5rX3RHkpapSdH+422nVtwmeuXaRX
1FojMBem5x+gURLxQxIiiBXlqm8m+VBTia+kglheRUerpRO+8ep7qVgd5ILAX8vX
OVkZ7nXNwvrUNvCkCTRNnI85pNptmRoqmiTXiFv/S595Fg4on48dQi/BUWqYgG2n
sEO1vhWFTNqqh84i9PqCDvlROTeAhxfwHbUyrbKDUSM49Y1BaaW+hnbLrEkwzgN0
G3WThJDqYXP276PNyDbvP1hoJacZOaXpD3ihEic2x6Lxws0gms9+yWobinfBf9YJ
3tYIGsWar262ohbi2B0kIGM1ME6bJaIV8UeVXhFPQXl8yIQPgB/iTVWy13UDCvn2
uqsTyOt+LuT1uGrYhujH1+CgcMItG7LUn9QkqQe13KahFAr/vv1rH9OTOi2zEN3V
pImW7YIjOinXa3e7u8gKU+tLvpJtsEqQNqMQnu5G8tpHWBz5+zbu/iGYwjCUmtb4
LV87/vwtHA8vXwEa+gyi5ozdkqeiaL6Tu+6Uh7xMcu63BAYhHK+lAHTOYDBmqO4a
xA0gQ+zW4FRdBPDkAne3+Sr+tyQLJmXVli2aE8YwV4CcNjltiayAcO9iUfdWFgGK
KvNnK+5Jfcf5MuNQr0yMiXj/pMD/Xn/emAG2rd0wbAnnBNhu+ow0JiF8lCIJPEbk
cbusgd8G/l8qDB4CKl1g3XsxNVFu+vDlNiOncLe6ywgGdQNkowe3/Fl4lultbB7O
KIIZHuJ8HuizpsqothT7E2x6iBsqcW7ztysFqkKWtpnkFHk7PkCd64D8+5oyqCFa
afeWXX81iYKFfttf/oXlot+sRyRjaH/tdKCQh9BWtJaVnd4ob1aBiM++8EBJB4WF
jsv3sk+RmOuldSAgd2h6BGsHHZtQZQOlBvJrP8OMmw+AH6mNAoogFMoati4GjzIY
2IgrZZFuMFSumqTx8VkNMC9rbUsOwxemp/NZmGrndhkL2ZEqvVkkw+eE4HIIRcfT
mzWehgA8iIBglwUUpRVGuqvX3hOLn2lHvS369PKGuf5PUjfX5Pqs6xN/kojV+YPV
Sh6h12BrSL0OCWrnQ51MAUXemlzZ5MCvAj3oaq8OP5HzlhBxLFxFYYJ2TeYbYVN3
hLcmGbQqNCk1oskb/sdvWtcxA1xas2qah/fvpI8UKW7e/6isUzSfROUBk9C2bhUK
RZzfqIMqdNRCAHRxDIOgIk3j0PNoBcZWXILcTdLQwCjK75Sp80or0rmpfPJZZPdS
c3sTvaqrYiAwy5/PBrzG6B7jhFbCaeareshuUwj5lrZ3oC+Lb3VY+ZRVAyADGTGn
n+lgQ3lqzl7vx4cbklswLMNQXhOa8hx+Hqx3zg0tY7Vo/Y0+EqrImfSRblZT2iEt
HxUoWpagnR78Ma5JxvPhNh30VD2bf3VGt2PjO3VAmw5gYQm+qff/w0kPjwURUu5n
y6eC4qTFhdasnEhr4gcZxCfkc7QJRFsMpp6wBUYWAB6ksNBCBYJztbvYAH5W+oGF
8pPidifKW6uIFJv+//o2f8aLPCO1HJxH0Kv8QZjNRL6DPVMPO6KJaEvh3sBRJ8K8
0Zg/se+4o6Jkvl1E8Pw0a6iI3nJtpOt2T5JQPYk9eKLYfghrrBvBIUXevcdhko5a
yoFy5u591RKPw/s9s2lE7tnxMWtEgxacBs4Ihf2L5ajjVvglvHBwA3jNhwTfbrtR
b6M7C4+diOrPdV6+Yo5TXs6Ipg/PNNFFwSwuB/e9ljpkjsmOwEnR/5HcNcrOvhKQ
TGKJCGGdp6P1KuEN7FiIOlOW/O1YhzOQZDANRfDbZWDM6UkYDdozWKtCyEfHfyPE
msiScxcshkYcESs5tWRQ+HHfOh3AvfdukxU3VoPdFDKsaqwaGm/i+PN9Tujgi+dG
l69prMczb7QjtrlPDt+UDKkVfYVADChk9r5qAVX3PhVQyCRdPqCUt4QoruobeD/n
IDXen3bPR52dG9kwAT9rAvd1hpJwquSeXkwFAj9K4H2YR9ggfhWOB6qTU98DW6QP
gRUiB3GdTajAfOoBb0hNI9iq5YMnal8DQqDoqE9wqJIeuFvOTFyBRUVJ9av8Ifp5
9gL/wbQqAXjX+ezMjEM7HYezfuURVYJe1tgXGHH/RHU9gumkrM/xAqiAm6HkVh7X
MPoAx70Jg56inpH4F16drkQlUb6Cp/qge3TL+OHaVuN2WvFAk9WQlGCyxUhJGEk1
09p8FaXMxWiOJDHXeQzwjF4JV/bJ/2qeaY2XhenkolcSr87TU5fS6ZSRUMWUNR4Z
53n+nxMdNpzUCdzUF2z+DzNThnUmQlyLeOdwjkYjw/PZkXpP4tqWWkfJtZy0ReA3
sxVQG6c65JWqYsmSf8jr3H+JlPUbpe3QENl2X7EL5CLh8QktUGLWro/eVZCnrZQc
ycAUlr5E1Be/28f9pdQhFt0t8g4tYcQktdUaXxl8Ozxji0d0beS63yhmr6AnlO3q
7rklpaQ2gvUXPCinptniIPaiqubLANrKhOCUuLRCtcLoJgulE2EINC4DYFt0vIV8
UsIn9li16+QD3R47OAomTR0h/QqCKA82mHIp8S7IfHm2PupY3M1BjsGaExpaFd8K
gHEbfMbc2eIzvZpOMTem+oDsjGTFXjOUrGVUxuW4n5DmBhbhJQeRtZibnMsBJ4GW
ALMN+zVNMLoJajKDrGiYPeqrPQVNiRk7dx0F3RdUYSNBDrCJqIRnSdxapwckksj2
ovNq0rhs5JY+/tF9Uw/H1KdmpHLWiCPgZNJAr8TmoA+MUwkE87HxQ5lluisHQJ7k
H1AbkXqjdkRCSOlx8Ftn3lnMQUjEcrY0cDaDaz13QbPEdVyO0gH6jdLjy125Mb/m
oNJMDMcVlkwQOtLppsg1szMXe/WTVQdc4OZqP3c784Mp2IRgn5NcWiDnAXDkoVNS
p4qhyj6JWrds7H5z5AfNckcfQu+rtiLc9y+amcg2h223bULb/A5qzM3M5u0Kp6Em
vL0+gqHGZ8PRtlWR2HfwSTMB7cuh+UOyPxdTKuHR+f8UrykZJ0jB3Ii9eK3uipCX
bj7TlkwSMr1Sv4JSYbAwPm1UzDB4DM8jaEc2NUIY2/5n8kv+SypQOp8+KthEZo4p
G0fBNP1q+R60RijTUNj/QGNFL0+MI+l94qaxESgxcZ/tA1/tHvy4BZAaHjjGrbbs
BXo5uiStv9Mw6q/etVowVQS+p+aT4+u6hubQQASJf98x0dgDs9QYPOvNaZfzLTPj
8wpWAP8VFdxGbtsQAvOyxERyEjeKhFpMOuTp4jUxB/Np0UR6o3fnD3Oy/Uxcouy8
ws3fVQUk23efcq2csSIyqiRuH74uk15rycHNHSvf5+hqgfX7i14bRFPIm0+EF2Lb
EMOEhunucMik1d0Kkjq/Uz/5BcFnqOQkzaA8TN+iSTPTZJwpL0OGthwTIjnbxRGA
faYpekGNtYyLcNNsfcdaZ/0aPEvc/hPowOk7SmMQA+H86ZNxdjsYwW7UkcapYaj3
qEZmtY6iDLO1tM6ygzaUJCpMk3OgGhHi2X0v4M71FWOGYEubFOXymm0POS71hRRR
ETQES5g34PQoz3JdYomtNS12WGVjyFg0yoL07q6kjOcB3XVXeG0nAVMuJEUo73K1
0kEKyzgHEewNq4iSUFuGnjMICW0E0oz4doHD5XdzpcuE5/GcK2knA2//iieGtGTH
qubDMqHzrfnjdQPRcpjPDwY7tQN/XR4ejFUU6/6PORMS/17LbM8bI3lzpXehJMxK
yszKNn/HXwDs7TjwO+rz4zlAuh9/Zyq0uXG21zunt21CbWlleiZW6TWikhGUPU1Q
ebk9PyRK84eIAusALUe9yYoPtS/4g4fmpfVy1xYyhtv7Lw/F7bbulO2c5Zdrk1ar
52rxM5gXlVqayXPK/IklWLAAh2lAFFYJUMrfxDRj5C1EASw8Mm/hO4x5sVIaGGp4
u+B2VWgD2w8D9OR4J+N+LSZTkiRmD4m/lM6WwsQf5T/1EW+NRX8Wr+uu9OOdYtmP
SHYkJPh8D0jTOpK9YtBvdASXITn095pp82FJuMPQs69K68GE1WJD5UJAPiSw8Fuf
jh1msgsIf/QylRGr2MxKL1TnSZlpo2gxUFX5hn1edcaW7hHo4APl1SDpLOmQLtrt
8488ko4COfaeO1orJbuDB+9xUh7E+jDy5W0CzauXyDEL9HARRF3aSN9JJYOUqdRd
p68JAbBtZ7nVVQ6Ek3LfRkcWd9WLu+8STjxgJd3y8NlJXQydSHcShB1qXkylQvcd
rKx70TjYLQQha0rTGGAY6Y/SjKdp0IbawGCpsxNtAg7FsNZFgPQ3IiIhnK1qOQbV
4vNKCBi+aoiDi25gQOFf14xp1kXZa26+1e4iXITxPBWLu7FXEpcWELXbas4KI800
EZkxmN9Vu3RWUn3aESYLNqaF5SW1iJkfKhRgwU3HBpNs4T3Lw3CuwRrpImf2eFu9
IkhcQCILMZtzTG2HsDz4LwMYPqNxY9fEB7S0BHTRnA4YUEwm6+FDOhxlLvmPqS8V
xOKn/PM62VwduPUqFUEh7Oooh3mLc58Tqglya+QLIBeMQ5FweU2m/QuyUHsWYJri
EjKtHv9eB10dFGLmGTiPv/zuXuBAEtDxEEfKvsJYMUjrr/AXjLZ8nr1cgzC0IJB+
kvMpyrHPEyhN4lFVg4peWBN0P0huUoekTb18Dm0P1eltA4tKrA4wYRiDXZhBBnML
fBHb8czACEQzPqaroJ8Brc+pSUxMvnh5Uh80GhQAen6m51TCLWR+Hse4LFJJHU7K
bC5fcmS8gKQkFuQpcdbMLx6ja0oKZsflWyUIvOxbg2mcFJ98KZPl+dA899vi+CEP
c1kdmGOv7bhIQPNX68RLbAw4hQWJ1ZRQojyJekcI7eMaiD9o79FiduCIRcUM7e2r
jyX3w7SaqK12u7vCYnSnIIMOySLK//v7ZHLQBdQQ3dCE7VKAi+dcjlsGTdis2MGy
RvX5MlE0e7wEIa00n/ZO2ktYOwoTAF/r/IWxiN0v8yiaIyyimoC2PxtP+zHvOavZ
czCmQHAwe/1ZluIONYX00S2a8M1lL7u9vGMdPBrQGx4XgE0Q8fOUoOJ8VZv/Xzg8
usR5OKDTE6c1iBl9fsjbW8NCUqVP8fsAwUcJ/E0+v+mEk9P8UgnmTZetbSawqWhd
FiblAFG1yq1PI65ZOhvWpDKyC0dZMCD984ZjkXFLG+lD89f5Tk7kvL/JblUDY1TZ
bMRKiVUurTQ/R7wHxJsHd9lgy9OPxPkxLCN4MfSAF2USLf1Hwo9weEVIKvwzE5F6
S3elLBGyIAREsK5WCfWLW5DwwhDRMnNplK2oaIJhtKg0MwCQW2cZ4ehOCL3XLSsq
eIbvo2k3i3pAQff/QQwLBBfl+Y04QGxHLcbY7Cf7KF2zwFzS40iOmCEiUhMo8pN6
pbl6IEaBnyHRGvlzL6jMP+lRFjXPKgndNZNB0C3F2s6rS8T/DyvICTlz75Sof4AZ
T9gOW/6yp/voF/8ShSBIxVuhCgDkq/jGUaj6L576D4j7W8Fnk3e4rv78V176O/cv
1kADxkfmS6MgX0e7yj63Ts8FiMVSt1Wn6DB1YUiXRgdqewFoeBccW6Wm+zVfZMxq
EDg0CCy+j6qSjHzCPIii6M1z1VjBosWw7sQ1potcyuyrM6ZHWdrU2Y17cyJCnhdn
E8WluR/3qAcYU1QUKchy13C0P0mbIbFFwVzngALRdhBtmwMMfdkQlCbscrqj+COX
ZcP97rvaUkTY2WKBvw1BPtEl6uI/c8Q3bVmj7bb3l4rgL8raL+EmdHWXBFoxwc4C
ST+9j6VAN1MhsfqsZI34EySgs6HvvWUQB181QZMTwj8bxG1pNczT/hQlyw2v6Mz0
fAds/d9nAXjD7e0Ogvc4hhGHGIuLeCfKNfTBR+eno2MzapjjABtLPrB63olvzSVt
uZmoTWk8Mh+Pok33oXnrRTfEEcra2IsO45ydd1tdb6k57ZL8bHtKStJnvm0rO+BY
N0dU2JJE5i8sgo/bHwO9y4H/p/iW5jKsETkU7TGJM7k6nBEAIYv00XINIjLeVFNh
3BHJpzk8iGiKYEeWmvTiwd+xwBjzFBFbvd29ih7MSWMTmk9jY/YVMhA27PO4b/eB
atEGMAUQUzcVNJx5LoHbH775PtRjxTLbyHtpV66qJj2ZoSGycJvW2VTUgnhWGFzZ
IjBbcWfbkwPyuTjGXsgyKbZe/fumZqXLnvQ2ogaPs9+r3tK3Nfp5K7/EwMLnrgUv
UeyXqw8q990gGRWiXO+z//O7is94hwYY+3CmSV+uPqe78fIQZvN9k0lMGTzsfdf3
g/5GXhoEUftKU0VK9bXJC0lpl5mx65ugSelx5/P+9/sms9ZV3UcrXousFOadIOjK
bjMUsEW6jSyXO7+LcDYstrjyc/SQZiyGeG6v91y95FfiLojgPW1t+to1hZ9Lkhsh
9/0CxOHFq9zznAAXEqmkCEooWb7unEPdC3iiq05BKEJeET5jFKTmvPs0jwNUX0rT
jvCl2MDJx2hRoMmLzNoeDc5QUg6qKryBIrCfBUEItV59Q1msF6X6f4PSU8wzzqoR
BV4qcomWL6hdZMmn4FAvAsP5cNkEU+JgV9WYbcfJG1213F66XEdkKVuXUKq8Q4Zj
cEEsZ+sa1lP17MFbQwbSe95wD+339HYu8wrBDh2qHWv7HQgtTYeu+TfYLSJPi4Yf
1M/zd221Tj+9n8sXD3Wa6n7drxhovGvVACbtiYmGhGaiYRtKVAFysW7BGCXeF9cp
nC6N/kBuJGwFipmQ0SdXVPT1ycgUSDo2Loxp8BqtYqiZLyymDGd2C+2wWlEkap1t
Bk/2lnJQE6C+4DUpUuT3dh4OLOxoM63YlPTJrZeDaOayzVFDtd5zAaZQTi7284gC
uLAs98yV5wysLEcV/95ZPj5VSdw8N+3rnORdtUdYmXd3ngsDSPIDB7oYHWBn8JA9
b42o380rHVgSGwoyJCQS2TpHX7T0h6fXi6Y5ZAAcjA5mJfzvDFgT3TIvtZoKzCvd
Tod89KoXvQaErc7PZqYgQBSiP8qICKLVxgqa4DoJF8Ph7REb9yNky0W73FxkaT/8
gi0bWPuiTxtVaz8n59lSjf6JimZKTD+klXGYGMJAiJMLZuG1eBIza33o2gjiATwO
93KUxmao7ojA0G+F9l12ic0ct7Ql9ims5S4+UQAd6uTqgNkKcyTgU+Q/hQhjQoiO
6G/45EvnL8h3SoZ0U2qsTsGEQG/lb/5NVc+qwUfitc6V70Wa5nA8cOpi1iN0fEJb
N5PUIniFhhDseKLWfrZKjy5JSWWmVnBVE5X9JpouSukXfyLvCNWz433DyqnjZU7h
1xyWXoKsAuRngmuy/U7B1+H8hBIIXoG4i7vEUk5yPC+LamTO04eXRClkNl21eiBY
wtt49rDEcX2PgnkxRZ793DyjQOaUYmdjK0KwJvg03IJGznLnG9irMBEf40ehi566
LHUjK1LBFz669s9ZRrTctVprlPsYXc4JkfCI+PHpwnZFGxCsiUc7KRYsnguEWVwE
kn74gT9nnBCBIXaKsBhGFUWDrZP0yVgiXuR1BSSb9ddP6q+Ls/2FyMmHX25VheUr
zJSWbDlqQkykQ8sQoqb5CQDe+fDO9USgnPE1z1XA8kGaQqpWxYzXekL9RKujjTfi
Qz1hfs9c1CIjyenePYS+0x+fNrzXJlpMwqXFtvNot6VKaL2ER4JSaIrLOJYPtXJE
1ZrszZifFB+8Y8SHU2FMkkPB2G0fRee1T/+jP7AQSSeFXaPUM2A3jf54Uxt1/TsK
8X2l04dTOXRvORzRnr1FJKuCsTi9Trr4NNOINBXZd0aQYaf4UEXwkz/dXDRk9ouD
Rji5XkxOrhsAOqp81JdwGKOTlepweYBQi1rLuBxox8/bNb0/kqSU9juG3XhvpdMt
6XmVkbtNZ5bKJAosu/jDCkRhslQtEbnvnIf6uGycndAHOHHNKbrwIBroyTG+NyCP
OByQUxCY4aZNcNuPYpJqpwrSvsgoOYqcMSPsqkZ7qa5tj0BpRotQPZwltu5n7kqK
YhcLGFLfrPlz/WYdSjv085yJUVlRfX+n+PQoNkQ2zxbEaqiLGWtcXUysIJnnhb8Y
BXxbdViihiXHXMQk1Kf2+YU7Oefr0rUX/iCsYu+diWQHSG9UiEQ3V4+UsKIYjqCF
tDEK7mJ5zAfj1QzQIpjfyl/xfyuad/qNEhmx1wd2NrLgIS87Oilotb+oxE7xfsnc
AxLm1t3Z1bKMsVP8gtV+07ecBQf8YxQB0rwoTfOk0vMTTRcqvUlJM65hyw96n20m
sGT3W65+fE4c/oVXXAVFTrKr3yCmf1fHR4u460lma3ct/s6Zu3ToVhVIWI0zVBoN
aJQNFiEoZoGQV41nsYS6EV0YUG8e3G4nB0EskgYB5Mwu6Onc4HwyhRmJzHv0kqw9
3+UHPAMrM48JxKvXUfEt8xbHKi8IX/f0ZMlhco2sljojZ24JCRagRrfW2av4qQcH
S97hdtlJ5x7Y7SSxvvC8FfnIprmaQKmU1KxE0fqkGI7ZT5rg4YfH5S91l27ajf6l
zqiTXjWgCHnANlzw+erRhy9y2gXvrZx5gqWa0RackUMG/Jmo8o4aoEYU3ySyKfrL
zIkHJP5HytPfnnnep4kWMkq8tssoNv+9CDjpOD674AU0VjIxWl04ry65G55+R6GO
RmzrL4T68miZhe0kv7M5vnOMO2BkN7ZXkLznuCRybwE8oZW4wJH7ICTSwgHLIs8s
v58DhkzV0ptBiIAUNVZUcE3KOoCV7EfHRWAZHNQZcZGRXcL7NZrI0alyG6WyILTG
s3OeTXitiOspxNSXVbBMc8dPkP2XuVcMRAWEh1hwm+ELRh56PqBCb7/gDarYlKLT
jR8lhQxKrSxK4vLoxXMlByM8xHi2XYBrjfZ/2lSYj+u/yb6lBgu8RmREFQMxoWJC
GdP01YlQ6h+w2MIFhR83N7vu/7xfY+xOINqRrJeg3424P1mg0Jb2oyNGrShS+Npl
ym2KVygcJkW12NwW8LDuEQNnYGBCak0xmFx7BcdwHdTjMlIz2nVnx5WhkJNToh9J
12H+rT8NxWP4KwJze8G1pnkK0oj//hxeifz514IZUHlw42cW1fAQh9agWALqi6a1
uSVHEECa6yQRIaowPd1DOHKnDEDWZSi/udL51z3X3HMzMiwp6hqG77tJmZmSeOS3
wI4WhZJeHk/pxrHwYor1PBNkVV9mqIKHoPenvBCG95kWpZuxzmQN18vq86+6/j61
gkEn9Wd+RzvEWcWFAyqnNy1xHtZjAGQF2aQeMsVTU45vnLfKk6IwuxLsAmxbjyYM
+yDnCvf3DGTVAeKydBR/x20d1WJ21Matt2xi/TOgaP3NfJMD5wKKs9nPsPsPaB6+
YPJ064LZtxw8AwWNna5sdu5ozGEDvYjqZBLQTB8IzGuh9WsRVoR/bEqBSreSAAj8
CwCkJWHtI8lP6e14Xxlp2siETXC3IBNoWYEIq+lIkx4r5bSmSZBkBi4C5tuyOBRf
/qvmpaELLTqK9Ls9nICFdto8N0LVSWWbQF/oRFPNhr8zBJd6kYLjwEU0w91I1ECp
IDOcJDiBBv6NqSCEZ36CTtybmlVzamq1uZ91rxVT5QRYNvaI4wD+OOjkj2edvEQr
2nK9+AuPhxnFSXQtCb9eS7KWTJpL2RUIeRQYVV6xRSs1t8QHTeHmyeH26a4bYioh
VpGRkUhEWBY1almaccvgqK17LIrjUKA/rTGVLq2fXZ7ude0T6VokaGBvwgvdWo2m
hBoeK/Y7euDnIVySExA6BYMjwpIYD7xAHA1SOmKy7roibiVDn2X65++2g8MMk+CY
Nq8otEK8yoZqZKtNmlAj6vQGuCsWO8NJCrpnDZY2/whXof9gqdQC1+JQu7TgjXab
5aNTJ9gExJgaalppDX2sbGLBcs96cpKTExEP40x0Bmsrg9LJbByRMQmkoDMSPAof
kWAed3A+G/4WuZd0LrdA0rU2/lNmk1tz8BUeV3Zz6/u7R2fy7Fll8WdJp7k+yn9s
CCOjqCZDoPL61dXreDgEW5jIY8mVXHIJtqnV8BxE1acuwbI5MH8j9n31/fcUlkNU
VC/fymgAdtDRgt4/eWQQ2tB15oIWWFvTUP68f0aVSrN6858Un/IYbqMBuD0RZ9fM
xSlJDj4DRPJsjFKk6VwyGtHP5QIMXkkuiyDZIXM2MBWfMRtkDyi77GthZ5GFahh1
PAoQju4i6zfX8p5uF/ZYIeTmXC00MFLsewG+k/x3aADvEy5elVLZizXgPvkrtTjs
4WnSynrhWSaY3u32vqUFRZ1Yv2DVRnhcp0pB38iQnXXVndeL/CV/B5mHUrBvX3W2
UhCUzhVfWSo0m+BobZC9UU/0vaNzrBj0kTh+VXZVNqvuO33xQwcNllSZrqEPpg9O
cR5r7mWC/CjQXZmxjKzpGsEdHZS3LkXww9IREXdWgcTo8JB9VrTFglVXs16Y0GtO
QV6ohamBJdzGjjurJ5RPc6Qskz2X+EEL8MQzs7lRI1S8SACwKKQ1EKSNYl/tvc3E
JIVTgxno7sM7mzMR2MxbnyPu//p1o4YeXmzx1UkTkFSfeabth6RVBDx59ID56E1q
wWbPy7XagTr19rxZ2PV/+xyQOcXiD5b1wiNY+MOFBcik/tBcAbeaQb9vL0qD2psf
8EIwTJtyjVE3Yt3i9LDBhugB6rBIEuopnZVw9E3FYjcfghpaCGRtEZ+MHwyLzU5a
gI6fnttyGaPwzO+qHMJpIPUOD7rS7aX4cXFwkOZRmb6SCfuhw1K7Dsaicd01t2Y+
J5KM8xEiSct0z7WYMI3mgOXGv9a6pNAQ8jTrjoSQvsu2TNQBNi+ARAaKOq5xl22y
Kn89Yje3DrfUcY86NL0IjU00TAJZYMtrXIMZxmRHZmlGBWFkdZqo+O4OCCZ1hKLc
ROtqpV4Irp9FxJgPR7ZdYYlYDl3qLGaGv+WvtDWuenrcG95WeKPuMEA1AlgwCGGI
WjHDp3I/hdisjySsk5W4J8+/bzlAntPXr9baZZYSlvZwS4UuxHv6cUyTbgvuaCfX
aQ8upafp6MJ+OAN95l3jlaIK7F8rNiCQFKNzrtss0Fq3c6Jv9Jme4bVx3k5sS0R/
yF9O3jxbk4zxq4GarejmO0OJrqfwyXr6L11neIwW/JzpZzhuwXJSC3VqdJeChXD3
7PwE0P0LRrXQ5EJaKVrOpKo+mTR8qnZoywTMmEqCBmZ1RZEoOEfAgjXFTB6fcTDr
xRMqrZ4p5hH5PlglUyeExlesYDpo6Ky/+ZTXgYxTe5Py+gOSozZ4c1CAH6KUZD4P
V3bvFABy7bxliOsHFFs42Xm43eBOmhhkjfI99SxZDID8L5XX58PHm+LWIhGGFdv1
meuIoCtto5esscCe8OLRK2/zjMSMfuLwbLLs7uHkqzveuaNNDSzwgjecSqq31VAv
CXOBU/lpahSgQlUL+4Ehy3B1xd/55PTxHEk4ToYu3+0rWfvpWHWbGA+G/nYGPa5i
xFhLoYhFxlTYWdp+qGp1RYm9ZclRIwHSHt3ICELFgK68bySzocKgNvU6/by8IsF5
9PtRux390b4Uz/Cd6gtqtLOlKxJoWIbXnuDiPw1PJC0ayYIpvSuHM2r5+KFgNlfp
lzFz0S+e+iIX36PMsONdRAmzh3GnS2h08OVgVa3oEWsJewKLhOaDRO4HHW907On9
dFdTnGUatPdx7z1ESdqxHwo2zJJLiND7E/IHxGQdGiMIfiXYVyrEEmabYldWC4zZ
g3YupEeO62mqGV0ub3Ortz9rj4mjhDBiz5bO3O3qh6Vj1IP3DAOZoH2vsidQTw03
y3kkqUntsD/f9gBigoapDMe6VdNjPknhqYug9utOS5LSTCwmCWhVOb7ZtcLCc+tT
iwHBwntvFkr8TrximDemKty6BkP3vWgGJqrcsTeEIHJHugkGEb12LKyXMDEG9QZx
KNn9ELzmnU8xVtz9NPUjlyHSoTuT/XH3zFD95E3j8tpKydIV2Bwr4K8kF3dWWyMY
/5aIZdEnEttJP+JbNCOiQaBUDqnhtoQbUrjzAJFciSVrtH5kokaMbGU1nIASNoRS
9r5uhf89hv7hE9WGOVEQrewGfQyIehxbFU97Hv4qt33J9YKv/U543mCXX7CNTBHs
ap1tWKgCylbWo+RBFafqvWVv84VneS7cDTOsiUrzNmhKaK7zIjR1noJeAc8pCR+u
xM+TW0oTmKG2dGQshlzZ57gZ0Wus74JvJB2Di4yazI66CXgnUBSE+8sKA3n1JE3H
xOIr6dg/fHJhvbcC0JaDIPTGz38yus21T8Fy9wDs5ig8+zmAnjbkq3ObKgSnab8A
8hQc/8L+lf9bDrMNXGW9szcfI3KydXAPz492TRBEyAf0tx4loOteI+KFUcb8zg3u
Hz0PIQ4NeCYGRgWqdB6Y/WHKDFg2Tx4Vh16vCn7TmP/Zfp6h5KbvUE9VU6vlGm+0
uChgZPAiikdUwNhe+0s1rb58xd3Ng+LTcFSiUgzuk9DNBmfkD0MZiQtPIZ+Ba1x5
xzXhgODZIENRcx7Eo70RsEc7asBBvHtZYweely1CAHYPUHTagwfFSunpBfR75D5P
rCA7tRVEqZSuUV9umuz2M8WtidbccEi+lZlY5H+lnFkwphMlUaN2qsFi9nIynt5B
Bt0089+WNsuAN+WDhr1dokITud5jev1kDocSNq/PSCk2Zo7T5WRoAaRuZbE3dP8L
VvpqKHWHOAQIBrIjZJJCfakdvM4Y6UlqqxBkW37qE2VDr+aaTTvEWMN1OwH3uqWY
3MgebOymfMt2ZpTwiDW0eMyh9x+p2N6Ed9q9x8daAa00tA1KO2NkCvXbm2d4fdou
oafEIWSgWzLPtjHgvKNV1BUuQWiRf9fqokSZ3CKbHdOgdFQNncycCFr5Rf9YZK30
XOcE1xPY2k047ZsJuil4XP+n4OmD9dTJpx9C+VQvwrVDh29QByRh34/Bt6FUvrSb
iBWStpkJK8IBN+g5fo6felVM65mDzyxbGrkadpfm1Xgy2smUcIbRazvIphDp7uMa
NkzjpmR5t7baUIj8d5tbBx+9k84WJJQyjX5VTo+S4BYVTEX27ABGK7v3cKLrRqGY
Eql78UfNfPqcZbZC1QCwlDxwhM67KKTrHS4ZZmUiH7aVmW0vW+YGghNi0z3AaMsq
RGQK80eTkv32B2HnlJmoZVUXdWml4bMHOL7qVMS/gEreIlhqfVlFV75D7SiMyreU
uuWcXR6UykXc/W8ibuNUN7rPmzobG0YFKbND/UZVC2/1SAtt+8DghyOrWpru9CUt
tdUTneiI/2JF3KUPdm6Aqd7dbZKTlK4VWuPe2d4vIF0as2tOLbEVGnxZFJpKLWuN
JgQkKocNmB5L0Kj9mBfrwoPIFC6EtaUBhMeNNSxSpXG0Ue+owkp1Pn+7NZE5lsYM
D0MTfG3bmiBznBCqQr4CI5l1oQzSViKHwnniICtRsMN+vkh9/4Bzjrlv874SlTYG
+VlWW6LX2Dc6Fjtd1xX8ZGZIGL4ooRTTytxwV21qZVBcJ768v/blXzfFkuqpF3QB
a55q27V0gI/4SmtbV/NfnhoDgfIl5FV8eZI9w2i4ZNMEfiiyI6H8AbPty7fkgnjl
ie6rufnDiiA+fBTgquEgECrHhN3sUvhT/nTvP0HyPrzvIPAzeQxhjdj8CHODEz13
NB5+MlA9KAc2T2hLq7xeghozpi+lCeODtCuA+gGuNt+rB7M1junJlH1/3CMJWkz1
oLJzbdM+ExqGOrZ4mgXb5vLUHw9KvQdqPBi3S47MMuYQvJeZ+eeP5afCQTzobUl0
n5AbJZ5BYi97ODzyEnQV51AjWPRyNs7b6Bq/cE+cvWb8ASSFI6oJdcAMeL3qZGKE
KVkdHBU2AdkCnrhcwmDI38vgyjXBMuYY/FJPf9QYesZ1WD9P6FjPXuOgskn+6P+n
8CRD0rzpJflOQT4zCMye/ehG6c+7G0tx/1GoseR/S2Y2usgrF6FHQY73Xi4YLHL/
rmBmzluh+4I09BkRcpRzkSyS57oygZgLWv540K17QpQXKKi50lhZEYWMA9Yj4Vsx
pDFTqJ82drtIrOfYSYK+oswyncSfUmmYrteLKiWHmWi9UE1+ptpClljcSoxkEbzg
PELiQtaHuV0LmG5+CrZj/aexvEUo4AXSsNTqtb94ANkAz52iks4CA8DExoBvHTeO
s/WeLEt1ZMQFXtaGMRBCZnJVWRCJIe3GiRYGeFmpVdbJaXZL2+vbxlHF3tQvsW3k
RyNRmE2OgeU2E1nMv0yZ65WTEjXc8dww5jfdP9G9fb27cAXwcJ6pTCrOt8IA/hxB
bUpRNlusbtfPXvxGoATu5nKcy8u8kUryc2bk9WJe6VakmMr90nniYH+hCIpBSQc9
gsHKNTZcfZ1ZgqsCPIR2vWhXBOcpK7HKCL63KZ6nLhP0Z8QYxB7a4Zfs+O4bXqyk
XkxoRRbUE3S1IHhfcJH3Jjk6G+Ho89n1p071nCjRkutPSBU9tpqa9gxiHy2vUrZC
4j5tvMbxTeP4gP1mJpDVbMNeZPCNpTj0wZnIsd7QjdEcye1jiePZKloYcXtI8Md6
P2d197O7CVhQz+QfkBWvs2UrNWRX6nklOrxElZ9RRf+0L5ICJWQlDxUoFV7nJ45s
hZ+V5NZxjmgNoaHS5MWuLKpYE1qKV9i22GJQcdpBN/iGQlgAj+N6NGfsSpRS4w19
+wmX7gVrTzyfQGZ6VB+S5BbQA/0I5rgANE9PlnYdVnHRdxGvFhLtRD+vUWgo00LW
JacCrIKB6oBu6DGKOoCYWM6/96MI8N12hw0rji9tvT1if9HDahc380je7wZCubPc
w5Zhqq1z5FsuCAVNWipMN8wmlcZ/VqLxc57WCTeMihWRCRd/BXfvttl04pRWbsJW
IlbZiT9l0bw7S7OO6Leeg4F9/5Uhw8zO1UTdwPBWfZuvUX6licCm51b+NCAFKLDW
IMwv09nIhVPN0aBX9wOBDYhkLcgS6tXQh/BY1EtB5J51YjzFblX+lyhQElhq+gZ2
fkxbe1mIEZmEmfKhsomlTnuvov3xlpoX55q6wt3dxPAfF5fNwQeabY4fZW5oth/p
vAptTqYYoh5VSOlOlQIVdLP+L6HGGSh47OInPikK5vCuzvsPApR/M6GfP5TfaOkk
XCTt+B/N2wZOfouj9vw0VFQmFRLCA5G4Mul0NbuJqNDDP8es8eYm25x67ED9k7HD
eekxQzJrLVZFhE2aFQuNuIXhkPoIG/41Z09PNRE/Wl5grGaRiI0Q3A4NHoH2y7Ht
0+Dz9HDPAjUjXftgbzR+VzmnvsdYTW+iFZbiyGymg4R1WOIiNtX78T2jXqtfhsAR
QZ349t8TN2ZfdxNYWo8bMHK5byS2nBJlZlr2lUAVmXQAXUJlEf5pRACdEm+r20A9
vcPXt8WMhRnUE04PwBi/9qYz6W1juq42R2dCtbWP0o6YS6+LCTXwMpGe2Rph4v33
HPT9u2ZWWvmHuYJRdtl8+X4V2CPK8XrJPVPGcMpeOkbUDS0+7zbTgmBCdofX6s4J
h/kKfVaPr2nSlH++RJHqwz5Os3jQJmaxcPQ34YOxA7o3X+ztB5f/OhxTMSy66X0V
A4NLg3pHf7QN2HnqvE6Y8tas31yBrR1Zbk+8HUWbIvi6F0DfOBpFYDJe05JyOmn3
ignBiCGb2Gzs8prhllrDT8S6CdDq02anPHVGQE27nl1p/JP6Po0Z8xpupLzv1U26
y6hVm5P/Y0DPXf0FcH7JnScmhwtybFrpY/Ie+c9C115aupQNOFMEFKjqGzEpNHsB
Q68xHeQK/MSDkf81jPjAuRd+HUuhYGHOQYCpWufaCnxPj/mV76n9k0MQpltcGKEO
tLjHzpa9dNqCzZHNrqkYlfxPe16IIUINvz2xnXRkfV4uAfRKcS4usrLbzD62KP9S
oQq+56/kFH2POmqAn3GSoEqubtxyp+zRvkyEyOfRDMZNDTrsbkGrTZyJ9P8AkySQ
zYe91lFARabXio0fP8KFmYPPFOtfO6VgYniVgkSPWMtXYaVK54zmMDGDGlpHoqLA
wnJJXha76iSyPPIAjerexe/hNxwqH/Tua1WH5bcoo8Z0dqK2ifvnzVipQ9Wq56LV
DPSkExfMu53zv/FBIUNeq+AW5Auamg7q3xonFCqwpJirMV4eTvfPUWgYsKsVxpyP
UuZLXU5DZZgWlZPdY5olt9udSsWJNS5CTfPzLohk33ZCTtt+C2qw+ZBbqXg7jMXV
+Ws3boY3fevvPf4GnX7afn6f1mDJXvRFb/hbnHjg+9/GX1aQQQ9ntQO1yDXYNW3c
J0Arpt4k97CWCdCK7It6ad+tRJF7/Y8FhIG5aAmyLy2mJXUHsBJ/BwGirZ1/34tH
QXrg/569fhaswQP6CmtXFE6JlmOSUBRgDaWK6OFi0GBSScp73eyOV3Z6B52AX2VF
oTMUNy3lnEEjGH9U7iUNyEJe10oEV3kK6D9Y6q+RvVpPQXZGyHLAbFXuWfYxRIQZ
PBd86zHZV/D9H9CUWQYuv80KS7Qpiq0Dt4ROzkDJtvRMygy+StArjKFOJbr7xuYt
YRftNBgd1pdyPmtpcil8ZF411QmccjoYUrESMmAaPFo7Tpn7CmSwCuTKw8TCcNKB
xmQMSo3j9eWlx+kJRHe9fKPmU/Ihwm7fIqOR8jTrv5mTcPW6qq6fWhDBU2rh/260
s7irHzocespV7Mu/MomI41Bkscg/mA5yVvJF6us6Qk/RB1JSC1HQA8IKvJGYZm9h
fqX/cJOihwJ6Ad4ajYw+rYIgg4I3kIt7/UvLVo91vGykh6SkK/HQiYTBBQjbE4t8
YPg85gmegbB8YKp8wX7N6ZFBb/H2oD3HNemBHMVlMMgVfmt1mXBYkfrNVz3FB7AO
brGCRke8GCXLZgFF7g+zF2B5O7oDbECZxTVa7RxPrRCU6rH1JwFucH0oi46Z3Eau
spzvs/LBnd47lOzqbihujUzy7FpJshDBkD51F1qjCBkSc7khDZVYBh6csaVrQjW4
F+t6pC+mWDd5vorAmBhY9Usb7E2G+CBUaWgIR+KQr4TUZlhCqzx1Yahr3D1QHftg
hmrQdiI8JuvsKZUf2aZzyJSPGXnd+ODVMYuS9diCY7JqdQ4bNiYw6r+NfwH9W3e/
sFFufIVWSCXuBnptPxfY52QVcah80Q37H2Wl9R/I7SdzUib2FmRSv+iHUhRtRED0
xG7pK9X0QlX7W05wTE8dT2giAiLOg29mM9VH1qkHh0mwDwolLHOxZdz+rM7+Zh+p
IYJ8+tFOMoR/2GqvALsBB7uw7qqV3XS1nqmgTZmgIGQl1dFr9RFOFgUUzAnEWuTb
RXaewQybNomF7Wt/b4y1eN5cf/W1VCLwQQ4K+FHG21ywLaiUSjM0/QMPpUIftOSr
Z74HPrkRdNzWNpjq7cJy3mknGoA0cgPzd+fVlVo/ojQmYo4iil267x0E4VEO9ZqW
zdoHEpgY9XqKH0biPjwkNDVqRlf7oM78jJgd7lnVxh7X2wKpqotckMzK/hDjqH/F
wh1vOOq18KG7ATZVwQGwEEYBgaCXNDTUAzFDNEFdLpjr42W/XWhsY12wfbW1qTgY
GwO5UcfMOCu4E9kJauk3r4exoK7fVXDQllsEyB+9pw94r2HVWUwJIAIU8tLTZwGs
W9QCK2QYisha/NnGHzuZVo+Ho1A8iRC2siIAjHqozdh5vhhGiK4JVrZ17yQI3v9T
5ElIZaMU59WueICW585oRlBJJwP7TGC68LJWB96fMKfWwjRIDXJUckMBD4ldDgGc
VzDK4jB1HjpLlK6j1UXNDSFCutd+g9c74nSGWJdrvOVQ8GoB+ghXcSuh/tWMWrYh
orlF+/kiwiXX/WhrhY3rkIoCt28hD+LqL/bZufGkTEpBPo9iz+iI8llQJezTW7Ap
OlSDqePptFD2ZFVWEGWEql6KuM9J01Bc6A8LfsYpp1yTbhgj3PcBESIRnf4U8EIN
nVj5CReavU+ItkZh9aFAVAp19NDB0ikfyohaKY0ZIknzvCDPXlAp1/mdCEiXnutR
FxH6wL68fVvE5uxMfNoDawmIbc3Hu3UjdAIImh/dKtAcOPue9rLH/uASmyYoB1ll
MyVygXFjeAoF5Cn8Ke1tvzJs7nkESYECzZKaRDxAI8f2ggJoHPBWG0m4FDf2ncyI
wqv7VFnlUmSdoin+Mju/EvK5DNRJbIUC3lqW/jMRrawpd99Gn/RsthK5MzPxBhWY
gIoO8SRHBlYn1Y+5jF83u1MyKoMX8TMoQ7wRcss/NiHWjRnvKdWB/NXWfK7dOfo4
6FJdBOX00ZGTpf95Ropo8W38fuVCpNWBWdHHFZPR54ptSc+xmwD64WEn7MseXpy2
85fdgh0aPl3m4dOwVY6T5gBOJkTRVC4xEQYW4O6BoA+c8oWRhQXOMUHAxzrWSFJ2
xBWr0OWh4h0WdlJ/13pjnUpnw8DBJPFJQpvKtvFesRFe+4jHrwKLgN34iIsWgfL3
hIHYzHovbR0r8iGefeHBOaU0FYo4MPyb/0Cn0dARmJTtFA/NDrVzatANvZaXHsGC
0KcDcGXhbMV99KcZd0N0XpuT3PBna8YEmcToObm9SPkafH/0+QVLdMOzvFSLXgPV
LHVsaN+Bdk9vCcmFbVcMhaMTgIZCLXPPO/0fCgin5CL992Eugyx8TinppiicJB+i
bBwMFfkNYuyRWi10lL0PTD5aZG1zMWzlI/nsh7ocYMRUuIQ9Bzfu1ZUO9aTWHbsV
TDQYEgpc7u41vR5XWrWp94tC8icjzAUyHYo+zsWaiPDB43VYDDitLeJQbPMTCJl5
e21BEGS3Ats8MdT8es3FIPdgSX2DbiscKf+C/g/3jw7+17S0es2lDkRkxTqRkfM5
cgkRV7s2tcV49Mdl3Ih1QfTpQtDqZIMK6YBDeuTyQRi75AilHljGGeSXe/HXpPWx
Lqb2SUAFYsqjEx7UNPJ87dTySRmVhVKXtrBNJQQMjWPYoKt0SBWqedDGvembh3Ga
Rb6wuOb0rgsEJ5K6uK3L08nOeoof//H8y8Z7ZC1PK8jIuhC9v7Gc1EqlPMOhro0w
oknTUonDQa4Sre+iv3B/WofXIDYT+k6wTcn7ERQFHhid62VuQnW3XxptuBLyrJTl
G70myBFeujX+GyXldUF4Ny7WYUkBOdnjmiJiOCGSPLr8mHHGZokYDkOtFJvtaE7g
16xCugaXUwm1LKJvbC9vhY8FtzRjN7eB8ZgeOTOTuWP/9CsJkzv0RYDQpiiy589s
IsPCNm7NI6cVOpAw8vxUn2QnyE/Ap2oDRW1Up2awmvZ3SbH4Uszn4Pbtyve1g52G
2yi4EiePdFms1iMtnD4+AuOy0P3cdi2qpv9goU2pJ+st6u6CQ2BNLs5jqEq3mSrN
3KPUwDVYQXMuNaXSA3KzvwbC9RncD/rB3Xtjj57nJ8lB6vZ5JdcaYUAig2bz54Au
W+z+dPWX8zZeb225ErFtT4/OuPcIuo+23ww2P0X1j3w2646xrMBUgMEb6TE29x4s
dEXMVzyNTzvWGFLZQpF16gLrl0yPOz1Y6ZxdxgKR4NYBsLOmsIdXjVrXsN3A4Brb
dG5hlm+1nMMGI6B8W6UVcMByaRTRa6uThDlyU1wuI68U4yTojOAhWCs1kJfIgvjN
/PmYgc1wKP2c9CfMwWw1ZP7HbAHHNY9Ym2hiLmn2/8S0qw0KxPhHbpLY+Z6LFptL
pNA7fPidRuktvAMl7r/nZAg/434cEjCcyMX+58UB9/FfXF4Pf6jncdqGs9RDhU3M
8MS9l5Ls6dn243mcr8DdwR6NdAHi9kC3s/JFYIr+l09+MA1DkK76JmDE2EPzdawh
2ffm9NTn3/Q3/b+R//uE13pxpG4hYHIaU5Z8amO2b+1tqlkA2/nhRxdGdbMxIWHk
j7jqUFEz3J8zH4hHZGIWVtKRpRMguwbGYkyJp14tmMs7DwN3rYpjFayucez6Vslh
D8sC0Bwdmx7qn5R8ce6CU7FXJRtsXYxZdh8BzcLlFOWnjZa0TcUG1ZbUU3rXposQ
T6DjQl85RQ/ztWA6eCUOb0eyvVz0Q7JyM8yy9ESJVRePoBkdaskmux9/UuIo6av6
FMJ3cD0JzYSjCcoib7/zFW9MVN8+QbXYyWfxaFJwSsM/8mWuaA1LdiCgop21MeDU
eMJO/XFoAyX5WOOk0z+j6Kb3RHLJ1kVbUDkFRHvZpezwFwSb/skmAha3weeJhrSN
gl6pkJLa8XhwxWZeJWoSp7uoGSVk31avw81C0JD3egUBAf8DOvwvjDs3z5Svqb/E
qTUDVQXqGBOkmdZqtMjVCO2XC0K3MXecGfOqeIAFT8Pi56fOAPY9PJMXmCpH+Svp
f/NLk9V+J4hWlfVb5bXKhiqPAyqP1mb59HJrdSv4HdAsUxu753L25JEFCkvzZyXg
1q8/cHXU3IIW/MCYpmzirKd6OKEh/0HiiIAWGPKV3QloUYk/AytY61oudtdrgikE
RH6rACIartbXjWEyoNsdcIndb0jOrR5WdO8/AS+YDIop4x1alf13PqWitYBIlJsw
tn4DwoKV4s7+4jN2B0Ca9GiV9X2ceoi9qdYs5CR2ok6xV2rOMnGPi2lDSJ90jMEp
g904p4rFni1ZJdksm2e435kasYfDzGrutVGCPQKA+hu3AHvWLs2+1+BnEw1Me3oc
vnNGqAG7GljJbIOnULBXs8gMoQbKJyW2167W260t48ogi55ENkvTgperYBHK/EoQ
v3xEXgK1xHDuBDhFj4GJD2fZCdRkbdGdBCDSXvQ/o3CvOLoawxFomumlvQ/XLQiI
xQ5fU5MXR8e1KdwzUbxIkbI5LRpa0Bhzh+pvw7KFciMrT9BvHjc0IS12UQU048db
fX5n6qMXBCxd1+nA8t6ZOulKZKpfnlVvYD7dg69AK5m4W6hUl4TvjgL6ZDh1Wom8
/TOXfE07Ntne4UVol4h4tgwT/VUYPI9AXYVuw0UA6KXSTBj2HSsUC/igwyZm8GHw
o3flzsc0mSay6Rsd7a1X/X4P0pV3vCHm4ExTtq/s0Zz1OSL3DwgP674gwVUgtkVm
OuXeJlvq4DvZJF3qa7v7j/7exI/Xe45+3PQhU5LKMSolcY5KB3ttbsqU9UhUYOo8
bxVSsrikZLfaJP/8bprdgDww07mKxXvO4f6mQboQBiebe6a0dr6KYq1Z+Y356BO9
pqXpkl6gLl+riN6EzUgYf7lWmVicX1uFdwOWlJzeIxpnMDCEyEwKDfoqqZKlZoZN
MKVdAK0f11Z4b1QZt3IKd2eho12jbwmYqTTDamZJgauy9I0lPJxAqmJSRNJ8X3vh
si/YHA7knPMMsaTE+1s1UakcPnfZVFbBl+uLZ9b5d9gtf7vEE0cb0u0NRuROPjLm
VQNOoW1LpiKgQr+78yDpGO7JOsjps7ElDtaRdpB4qyZp4C7DOj3DXYB06JHZCdIT
ZbZ5XTuAHFjs1cxymfY5ojc5OZH/PNT2/WZAD19twI4Gf8eJSzBssD1VK3YcYdOw
sHh/G3XWVRydkCbgHvWfxuRjykEKw6+vz7mWQzrMWtiZx03sjCEMM8FfJ7iw67pu
K7bngniorbPTSeSmjV/X1ThDmKDqa2ooNhDLGgBEJvDVA+3ZpVB6agX3XWPWP4Mt
NL69cYOEb/l7BbzHo55D0fH7TKwc8ebmfiFQ6oeT3ak2jK+TUTbBqzbz3AErS037
daOONMUfzMG1PdY1EsUG/DKoQd9YioQhClIMC5N0PcrQgnV4ABjgasZyulnm3pSy
pBqPBmA6oy3U4g+dD8clGXOKSwOf00fPcPF7wkMZ98V9qpyEBSgREmvOcvbnlUSI
npbwNeHNao3aD00BR4obeRG6zY+ytnyLl73yQIYNM3/hVOPuRWeLnmXC2RzpPcHd
ntN4p6VReW0DAKxepzFaJCoF3Pn0kmeEC10APg7PEEdGaIj2+7QA6jfgPYyJ7MRJ
NjpRgVjHHROkcZGRfxqyDG2aI+LhOJcT8RiJXkFgGilW8jJs6Dq+dcVdCgE1datQ
N6Kf+Ol6MSlLCmfzDcCHrG2vMFgqebQ1I58ATRqp63CgbZNp/VdrpV7yU6FqXwDn
RcIGfBuDEF8k8aXeML12q61zO2V+toKikKpxMq+4IXJ4poMlNIFRsoT2DS93u2ML
tSuqGAkBw8M1oOGVi6ah90J2lSqC5FqWWACc8IPzsxbd/oL7s4vcmlm4bI4zIhWH
trPq2Pjm/JC9AxpWcZ5Bq+/NvZ9FSLF6ohK2k130WU7cXWG1Vpnb5biWzuCpv8Iz
4T6OYQb/bXAt9NDzdTyLmK1KFv+MgOf3D2cN44IYTU3nLXru73IGAzws5Ftcwk4i
VcTKolwnh62bn99+l1ONV87ltz2gqdGycre2AdJrfZRmx4qrNMRfPlTjBPdCUpbh
Wj1vop4bUTsGCq4GUSYdbl0+xFwFP6Eiu5foWCNAojRIMniUAiqAP2cgA4MKuCdB
RQ7I1yFDeuVWsNLDNdFr8i1NoLbStm1E1jOgk85VmEmuLHofuu8iTLbXYzmD5r1g
BDoVURywFTczY7ZCmlmYVL3AESZqtt/D2H5iBjQ8gFmajVzuTWTnfbiTA0ZPzohE
hE4uUKT/u/QRimui3rCDmuxiw0pzv3ulhThC7an60Wk9FI1yCCZBd8MWe2UAmcdH
i5tPBTEmSD2Yu3IXXMfsX/G/IWFeXGWo/Xj3WdR8YprrVrtwmu9uT+1X3uzcO+xB
HBbFSXtNIvpqdZzgiZ1ui2ACZ6csrEKm6SfroTHZ/9TSp4o/nmO5cF5hHQkST81y
31gh9hSuYQfT4+4PMZCkZw6JM4yIJ2dRQuugK5NziW2+SS4c+O37rGJ0ONVFM15d
O840U3XIeM+R6yjQSIfMRuyN2aZ77aq6897nU9HPO3DXjzVtuXVipqg0C6SXj9fH
YyQDAATDk8acC3YQTZtdGn0zwbP3sNZNkx5SM3xWpN9ziPhBqE7MIRR10VaMQivZ
DlzKzOSVv7FXFcJbuxf0tE7E35VjftgdmJE+XAsmzpl07v/O6zxLvDwS5AFDKUqu
yyuPiDxBItHrudymi4YZkOqCJJ3BAqhKWGp2al16Q+w/H8uLjrUv2n9NykdQBMSU
N+7V9/7mwzvu9I544qHO3LO7sTNj+wPwHiZgMmFw1nsTrlid/bMOiOrBiYGu9hhe
ce7ncjUI8lalue5LCRfNRop6Mp2YxE1M6BZgCGys/TISfsq6a7oIth+n4W8KWPWK
mMHws1MiLAXYgMbg/a995nJMAjFQUCI1OP3Cvh7f+pdwkg9FrAL31AwvhK6RfrUN
ph7m1oGFDiTdKrSW8MniLEWDjKFNYeIFs1X7scIdfxSV0zMNNXc0ICbHioGK+R2Z
hiWamE6kPhw31n2nLB2Reqm+xZem4f21vmj6WTDkuABfrSYK/AUTsPQIZBYjLs4n
j6vi1Y0ohwLrf/PIwyg1WiDVYT7+OKyy9NrAcloeAl8f364sPxQV0CPRFWpMfFZ7
/6+xwbnJkSRizq7BKpRMDvS+uHJM0/DKcpZ7g4KxyRUhaWbrk3YPoiTBC59qLU/A
HIJfDbMe867qViqQ4UITu7Qz7s7mCB4FNiEBqn8waxSl+8we5qVGLkchY3Ji6s3A
7oNVLVYpj4fUIBzXYRi4i3ydNes8YXnTy5iaIz5U10DPSWTk/sbaRWQBkPzWXb8o
hsT/xvwHPD3m1AVCTCYir6UJDXi7IdTYxPba50beMYO9FH5bq4anyCJIiy44IR2P
dgmPc3FkgRr5pbMB1UtvIgihhRfu+QS8NhOSxgUzwdGo/7XlEJEpf2KhARKeba41
uWNRDm/r7AX1Jj/62JT8AyFumUifq9dFkG5IV2U3U4WqUOHUjaiygUo8arYF1B5U
SQ2LvN7dnCcV2k5ZJRQ+xhfHT88t4Pl8qILE7b37iUMi7BlRDoqU8IDt0KEZkQeh
V9TF/rEqbmcEB+9fa1VNlpk/WENGJYRL2dkX/vYEYTjWz8IvFZiSOrKVQhhJ0bCm
Goafr3n8n8oEkTjlB4cy7toLh8Hjs55Ihz+atUaNj9/nLKy2rlONTaqtAkcDVGv4
3B4hxnGbkkfWekeZFgfnBcmlW8BIkXqY41eyaJ61tVODE24EWygpWHF/mC668fKZ
4kwfD2OFtZwmnd6E7U7pQahvldrfZhdYn3dzG26lOgeTTIOm5U6Sw7SGD0LhXwss
Mz6JHxnEt/le9DvhU7H5VZjIR3yYMMOE0NmAciEAkQJsWH1NGpJRBpuUQsHbYxeX
nLQNY8RSJF+NbxPiJjT5zv2YQZCmUiuR8omoSVx/pQbnPf6J5FW++T2PWxoSBB+5
j5QAszc+ruYgivSeSGcx3VniXp3QECM5e5vZTgYNiH9HgzNIFJ++AY7WRU+5N40y
57gIEhv511khwppncNeGKrAz4IGUqS5FfbNi8YEw8JAW3eNGoFrx2A4cgsucTvZl
SBIxoVisEXiWWEeqkPjr9ptoH/snLLWFDa8Y+itwaqSHwSzDv606255RJsJY7A73
0pMo4AfzO4Cp4r8EAX1yOfYvHQAo0So/5/kABvELpFieripSoDNvHS8jpLkVrjLp
4ZdjK5wzD818wdkBSfbPBDWS7oylsKyJmicxp43wt3bVOpvcvwOIYhOwhRKnsOZK
8u99g1pIk1yDNzUbTEUbFqub+vVQEHb89/KFwT6B2H9CxwVHtf6nbweviiu7kprn
0fOHP50FXIDYp2r3J/obun4P7HU4KScvY1Hv0XyHIn+8PX320KXEOORbT/vd3p24
Nxhuy6H75AXqQ9wTamkwUoAFlycHYBDkYtvb2cmukCW23a2FfwluRvTSRWQeFFsM
tUbDcO1vxiGZBM67TagHvMroxwHaUtz0s9kWv26clA0SD3oPynb5x05IrionizIY
BnQbnMDAYcBFGVoDgbfb7FzLNiEnIhylZLpPr2GS6vhz7QIex9ZkweXxn0cWHUGZ
aji3+vHmyYut4CAuFvC/9hNPj+CXzgU/U+Ik3MtPDBjR7XDOrH+F5OyOil4WmNM2
JoyemxdNXAsH9yZBKYamabCVVdklH07ml+rN4zoTL27lTdc2JzqAy0ABLkmkinNX
dsJbL1o7iHkl3+F24R5QN1LUY424lMx8dHcbbjCfyZkUVe3pmsv4fAerC0zbjmBC
U0oYk8FwcwbpN1Iztn6VZ9ENMktH4HmgkXDRCgR04U1e7GSg6lWHUJ1I5XxsTOtV
yyRT6R/8SWsv6586MO5KlrG5GNobIXAwlNk/vLCCYl245PgQMAlncN285e2aS1mQ
mzfW7gasOlrx+1uZYyFqd39EeJ5cUix3LTTJafQIJpy6xso2gg8/Ys5kqSuOOkUt
T7bF2aw21VQbLNqV3qMNtyWKLXnjwONcM9vMljxrQi0W/N1STnf0VON2pZhCSlY6
+bTXZuMla1THqS4Q2TjflCgRIPFyPA1vVXxNB/ZhFEABp6CJ8WQAgmT6Q59SU8pK
OjPuZ2Rrc9zpxUhpLidutP7Cjk9KPetylN/abQJ1u0NGNLjb/9BWC+fC45wqw34a
IAryjNDtwQ9SZ0KuKZ9KmaqSOEUTosofHdl4/BpzscTX9D/7cU41I70slYkQs9ap
S+7GOEO6o0Ig/p5hiFjkzQHpIeJ/eMr0H0CD8gG4R1mFop03LCwv1TYmdD57zF6Z
Vdrjn1/q7ikMF3LjPq+0fcVheeunTvPQ8/ns8lggmzLsUWGq9ghAdQYIkVPQv6JA
PltQoNfdwMgAW21V/uhxXn0XyPuHGxL76+Lc9jVyj55Hm7hS5EVRAf2GbO9b+9Av
IfWAoaanLHm2CiAmcvnaZZTFHumr7mhSHN8+qHpvp8M7Yx2cTjo3FRuRJIiIH74/
EWQ9QOmdr1BPRP9+ssymoO8QmcqiQFrOYMgaaTbl4rrNg91okMzJBfrS1r1XPF7J
jFAbVP+OFtF3IoUaxygag38xj7ZtcFDb0jDWOVY9auoRwlb8EpW7dgG9kyPrTt17
kDVbP1nDDQK/hd/S+TDQf5SyjaNZryhfLDhwh+QBFMxE2jmhSxt/R6GgjG0r4fAW
fV1F2ND+QX4oYPyM9C6T5seoG96AoCspLK1LK8NMMGvzT3U6YBvo+R0PjF1DWeFS
G1GpTTiJ7WHmfqGbXwB/kONKG4PIOT/EqWxmvzHXJTZYGTFIpBJVcRi/EUA2+GM2
9NdeUxfO5G5cyIoaxu5NAGUyFYNupzO1roJRpJSrpqGJ4d1W87om1JvMb6MS1tZG
naDN7mXmvm/6jiU/yryJ9fGquukNLk1kGfBjjz/ZzwS6dlzCtXl33U3I+rrVeItj
Oqc6/A0Hy6lFt/03DGltoBhQKdQjWHHnT+VNK1mfJFeR01YcF/BlZ7hAeK2lF5tJ
eUzuY44NKfVDn3AB/8xP00uyD2CPgAIOFMxooFFv66Ro8CN7QESwkO0f5PHQkdMu
l2H+SPhTKjnBP6iG1mlb5mDWbhqW1JpufHh+7qC9SSNlJj4rkWY9abTsiDdd/iGM
pOKeZe6Ynm+vQzVl10qjNPMQY0ICjI2Ld//SpMTTbq/5io8NsNyqXqwGSYt4SyoF
WQfvGty+bX7+QIzpTWVHDQNL8Lf9L6El2vvR9xbQ/LwdRSCkLx2ET5YV/JVSvBVk
5NAkWWjbZnHkR+cMqYoeJM/gC/bzgmk8aPUoZDwQUoJa3Le8A73xzaJObOL+36DA
UqwwGiDReDj7GzDPfMVcyYKHw52AqpsCyLDDQEa6/sMdn5UZUbAqCECMu4qV/D+D
dcQ1YszvwvZJgEjwhACluUoNt2tgB3S49rKgWagr/15KFgavoJXnWZzyNP5/UHtc
hh6/7GdeMAe45ojuu6SWBdRMQ0FJylJQM6/LkA0Sw4eGJN1UEKpQUHCYi0PBvMla
QUvLo2lUgLgzCqheCzuyEe7RB0Jmrfd118BJMQiMCpnX503LQVAMfsz7tjPYYMD9
UUFDVAGJNjE0j4532HabR3QUgkL/RiNLdFtCAydy/nxVVl0kdOC9M8enthm7/56f
ori4z4zurLiVaXPmeEz8mhp0kLA7dze6XfmMmbgRG7kxktjVO9YBSrHGr9RjuGxH
pgwxICdm7bXzH41G4sJ8SZHrmc6XCHDtD2p8xHDWY9adfXGpP0WkmMNhJwFGl1vo
fNLhMCH5jRMhxT1/u7JzOmpnzVafzuVVjdwthZJdGLKx12s0nEsTz/n5aaMylx/+
+M/PHqTGRymf9Ia6H6z/XnrEBmegMKqfzIpdUNGu9FfRtk1M5zDRkJj1YL5RBcaX
ImF2svI/stbtoLo4ijTjI+Pb5DkR5DweIgS7FbEOydDCaMrb5xJrZT7AQhqlZ1d1
G2lblQnhvzfZZWfme3nr1qHjtUpI/jE6JvV2TBYV/1MkLfcDEUoCEfqosyg5WmIS
KxNQqkfB6QwgYHmsONPKNQtoMqFByqOaj06zV8Gj2KaHkM/Ir0PUbFvcrHQR5Bbh
GlLM5O1b+2zR1sdw1YK2uOng7ybstj1l8kdkcXVghq6x2h+TzM/KcMYiAZ1eCo/c
9MmGxG8ZhU0LkZQMRVWZ+HzJ+ygtv/kGgsjKTvUQsgfx48odogoqEzQS1PftSq6+
I2rNSnN8VfNLaEYf0E9/5c9FWEOm1eEVoFO1ikTJtuMy9UOl/a86ye1jfNoWC86f
OeKEnZdujK4tYlORjMBGgMXKFS1DWldJYF1FB8XzOq7+byUTWYwOevl+0MEjnF8m
Zz+dGN27eZ59nA+LPTa22kSBgWOi5GNOlWmaidEVfI8Wbi6ljsfB9S3p3IRAk7Fe
bsdl4dJrWakl3KBpmuhbtbTGhIzX+O7He3fbrIDUYppXZVSTNtxDlTHEX18tRJou
bjbIlTmHoJS8YUUOXKMGfcIh+Ek40+rIMZjFJ5vvO8kt7zB/XAAKEPQuSFmnxDX1
CejzdIXvo2cyU5XmSOV6Yl7LGsLZFX4zOObG/riG260Msyhs3jiaJQSsKeq7iAiS
ZYOb8LGLeHkFGNfHyWSRT1LqajxKPR3PCg1QsY+5B9lrlN4lY/m4X1Ro6yPyl8AX
sn0PFmQd0JQsXNeg+4tWQ2ZTENPWG30SU2VXoZPXxmCqPSeZgym6Tjr4s0auf+YP
j0+RpeIeqLRt3NcN/oCJdRuelO7lrqqz/SmJQXcbGVmj32xk+ypRupCTE73EkqQ8
Vobs2IiGV7tzL/wqUpNdSGFPib2N5U94LYJnjm5Ju7O3N9e6PwwgOKqUabBv14Hn
YiTzpGeAM00ZJJw4BNMcusFwLC7YLY5LAdySh0H/Rz0972XFt8XLmoAJ/dLWxaw4
lvZJBEUchlZ3fYUF6W7/0LADMiAvEQEAnGze6kVliDPwhnaQzELnT+QVH3Fy3lR7
1nNtnKbmGNHFFa/BVub78VUCOgNQSYdegrwA+Fy/YmEL2r2EJLu3BEJ2q+xjS3IG
eA12dxkZ2zf9azB8CmT9HX0SwFXkx512w97ZAn+qufYQp6NcaScBM+Zu39K+guYz
OY22dfKsKnKRebyAlM0WNKQ+wsvmQ9bYOq7BpNvOwbXEIzCzqFRFHKZ1Z6K3+PqQ
evlZ62MuEAMRRWcOUhAXOaJfb1X47gxhVTz6Y7ghZiEdySr4PY19hzqQMXSzLYzr
81idQ3s25tkqYSYlgvAxYvDbTe6OBxqHS1MPU7G3vkO5IaXl+cWHhbgHINjuSb+I
cZRs5dNOlnrC44l4HtyPe7Q/hkQjtROXZj7/P5mUjgbI7IBwSTK1pvfCdRkfg5uM
9BjnCuNHF2zNY6E/wsNKDa8Oj80KCm73jrPznDTfBMujs55D2s3u4eQrhB2ewbLT
cJk6D1O66moG31hEicMAH7Gi7vI3DlskT1xWpm0kyj6ZLsNkmRwBbWvN7vJQoOKR
5VxiCSmvPBDk5+1rfBoZDwZbm1YRwgA9nFvIjLZwk8XBAZVkXWYrfA/ZogsXBLpZ
YpdFZ9DPifQqg41uayxCPG1+cMKqlQM8lOPT92z+zJf5iqpXFuY/mM48S4dDbJg1
g2BTdc4E88XcvIHQCMMzZKiCqfI9SfJBUTvaf/zaemA4VlmQtO4U3W5QONH51/L+
FPmoPsbOHNU1yAkEEuCzzV3P75W8HLtqmqH++8E7SfscydLVxWTSrvwb+jz0bFU/
UlPpsHxCkMTQwzHFLaupKl8w66omYpFZxVieCuJmgZ4Zy7bnIFf0HB5gmwSgqDIL
QtPxAzio6guSc8GS3I3d4aPHV1UX13kZeRTZ2xO+FTFw0jwdY24EwJaI3Si/AWdu
2mRg/MDn+lQjyLuth5Qn8jyHnzrbj9YryXEzZ6CTHVC7FP+mEWM7zhZA5Vzm076R
WC2RT6/ev4VH6iEQUgt3UlsymmhxUbx3cwHRHrX/uvz3d5ckPLn1mwZif1TzmCEL
56P7MVZLOqoJ/UElzU89XIKIAibIePeGhv+ITgEywGtgZrhBIr6xCyzKDLDQYHr/
0+XElJNXOI6PYaT6/tadQFo424yKJ9bHb13SaP3yrHXlUpSfcFRfJrT9uwE796Y5
mjiWbD8qjDzzwbP/SI/N695vYagPElqMowIAbokQbe1d7ULxWRFkmaNolYmlDF6i
zEnqnlWC14woZlHfZWGtcTKnAjtXet7ulY3kJT7FdKGfCMthdVYknOqK4WmAXEHs
2utztCwmkHu9ugAd/3ya95K3VuxZ5gcpDw9s/TfLoeRKTvsDiwSKMH8Yzo7V/gLa
kd/KKznBHQ226Vc/pqMxoEcvHQ3jMtst29tGhRMcGaIWqmfRQf5Awj0eymkqJfn5
u8UvoE9WvUJoHZVk/NQwnO/6IUaGf79NrjWKYG/aoJ5acaTmhYmVBpIrkgD+m462
W1vSh/WoV3zuDBPuaTFXsRZCTjCgmW19Hxw6fkgGOCk5/XqJFdjJtmiO4JYPs819
61VYVaclIuhkOEHBiSPnqzoB0lKpps4wYM9+/I8sPl7A3qG3mPajynHX7Zbq1Vme
Uf/antv56tQ+UUrlFfmt/2ZM/cn50fBetFy4XHGOw1/boHVKi2LmwlqiMymEceg6
tsDAyzI0b2OAclrY9+RKpxbrbviRCOe7Nw9wblG7Zd07ogNsaXBLD0sBGQaM5huZ
AbfrmnR2DbzmoYOJn552+Dka6YX1JSyFieoiGkoLRYt8yTA5wYy5ADSokq+8EFY2
Z+wsgNaWiWVHSy0Kd2e2JNpNQWTOVM2KbKEK5xRIn1JFuToWzL7XsoOoSc7exi5w
dLcUikc0UX5tA86GEKYKrOwKXi+qfNZZ1lpl+ApJLdv1qfvUK1LjhrZO6P0Z0YA+
68e5KgCDGrhbDtzmASisSI/PLeWytsLWB9OvXTmvv36CD9YVj3f3rhRZrUdFBSQg
tIUjy2nqA7SPLP/CKMC864l0oNJ2BJsPnvduPy9bzflYN1WE4U+/paTboD8pWa5k
Jey8xTcZt4GGE1S/EKnnPoP/XhczAynj/5u8foF17oa0MC/jqSsoyxzKb5nNpS16
radA2DIf029WKXNjWh2MDt8JB8CYMpR5oUF9/5u6c2rIUGVpLToOqB5hY2X1V91N
L/1mchmUu5pT2sp+Lm/ECVkAp6f7tT0DsVbJE/JiFyJGRUrkVkyG6+Ru1V7fa0H4
Kbb5Xro7yGKCSjKvmvcQVvCHXXgHS1UpP9EGxoGTtEdJ9Sei5ODbpyZlv+roxXki
dDwH82b/adiZxgNcwf8ZzmDT8jJPzA0eWtcnbFwdFtwLolkuH++bLBasdNNIivlT
XbppaBOGbpj4gfwfe2Py0OnhZwfQRceVHxTTYG0sv5q3CDAkffrnsHmmdY3ipUtW
Z1Mkva4VQdNIwvSSPNkQfcktU02J7JOxLK6qfPJXeyrx1uwaMuOQsH+7yHY9z/AJ
ahlokuwbj0Ux/E8Owmzpyo234TN0QnyzbKJlL1pKMWdW/bqHYtniWfNMQ3Q+5ZAC
ijyudt20mE3Gs3l1ly6Rd8acg+KEz1mEcKiWl+6Lhhp5YcO4neClL/1IupZLCt4K
2nSZHnDGdYe+9uoljFxnzERt3JwO4IAuJhXKyS8sCLZER5vYHnBfC9BGPS76UUpM
ahsCJzL8PeojKUn1ysUumAOVcmBSTfVdJGaO43EvIWTSax5P5xX9AmsZvSdRvARL
sFvFAq3vrpx/dMtW+gQRO22s7NgL8hNJVUuBHp+rnJCsLZppl+DaGNB0tA9zxoW9
mhdkuQyNwlLjz6CYATTJu9Iv1XFpHajCkRK94pdF+4fb/tpGC8DAx8dqSOFAECpE
VP/Ce2XST4IjJiHq5VYMn1K84Rnc57CQjY4yw7152ahxkbFDw6D5bT2DaHhTsAn+
zWPWcCirrOPorfyPlDSsJ8b3Kwrsi1Wf1OU0BQ4Vuvie0iwXQSWzx0XkmfVVMU1/
tgEXNwnWi4GeDPnlWuT9Btbl1kFUTAui/9tiEgCpLx+ijGswwQZc/qqXB4KR7A+2
gdJ52pYgAz41s8bWTguxc8DI5yn76AUnkyfR7LUjyUJ3zMkw7KPyg2tRhcTX09rW
tjS3FFdAHzN3CoydSORJlJKWPJIjFF6eM2flSljXujATVzDyEeMtRLDlBUf8CdFb
7F9lIcaHFsiwn0sp/dsgJeQD6w0MttzARSgBCxLD8Uyc+NXEMNrjhR1KMm724A2I
OUmK8CNe97sqQs3DgyjO6UMBbD9yUqUybZcW0FM1NNgTgaleTeoYYOI0hugHOGWM
7Y9MDfVtN/EAk1EFn15prhSxr2Irdvsxe1gEUr0va6RQII3tLNqXmDPApN9/C2fc
Gxqsc86agxkgdmEd+fakkj0VteWWG9x2x5Lyv0bY/BAtR8wchybDCPA18Yiw4qbk
51JIlUs3m/TV1T+oAui9nZ1nYmKg82vYSpKbuQR6FDtKoMLm9gggPr/DNM1XwdX7
ohfFiahZOLwn+voN+hTbjKDEydsgrlJ09Gc6BZd1KxrfAGWLBfQNzOKuW6kdDXQd
9LuMhBoM/ruQpJrH3JiJJTuvosF6Z4CbWFFh2nAb2WFnjjsVExfWGek1MBkmk7bM
qOM94LXn10tn2H7Uz6WfZYpNo25W6T/LDKI879YbEAj1COjvkGbF13fWGvxhNn8D
XXINeurx3KRKngs39U5X+NXmvW03MaQRJvEIBzAvUcBCM4flhgTV7MoGJG4Fr+je
wi4ZwamyHAFb6CwZnIEw1Zo7enkeQwxxL0ieSQZtdb/92Gvrc6kuic9Bla2wWtVf
6+E07cFDEiDJEK5cjx4+zxyUSwZuMCnQDAtxC1jT78PIRT5+aXs3F3lwerQH3aq+
pvOET/jNKW8qCp6oRbBcZR77FX8gfZKcVACtNURCU3Z8CYCTDz1M/rXJSKwMCsfX
6fbcoIm/mvlfPPVvo7ze25JKtzRlVYKUvI2FEhzqqWr0yTschYP6u4g+6NSlFlzj
zWQOfb58NfP8kvWscpmiK7BySAkAt84wsw8iLwgPrrJ4HBrqvVqV0YPC/HZ9JFEi
oe6DCdnZmKxTZzfuKpchOWxH3mW8YCgKPAnohoilwYQf63MdGKFctf/hnNAazA9O
0+yLwoTLceJlbnyIuFe7bCD5YTymAOIk3iRKjvIbaDz1SRWnRLnnbdn60SEG6HIb
ctoytnAror9I+pv7PBUu+0UYlxU6A/QtIDibSBdfbRc+zXY4GnZDzn1jqk0FM3mw
59FbLW1pbFiCKe+w4455LKonEfGIbpjlS+4ECwqJgapkVCZJ6PVNseNyNpcYpvxU
vFzhxC2kdUiZrOVWAtAIMRDdqPdPOWhhvWtoHyn1f3MnXNdtHLSQPu8o0WQylEN+
6M+BzHIhN+im4BcSfLJKfOjIDe9jgVA/sbuJisWLIi17NdJFdfPl6XM2tSjW/oxg
UIoFWqCcnPlvsJfaE8bHXEkNg0ZEuPnsF8oEGIV/Ng/EvhYZPxwRUDvU3hoU208c
pTNqt6D8YrI3ATXzC7LgDlWoRVPAi5WajYOcxoxjdhw7GQJHPNYSVOFqjf/xqKq9
GLFt/AONNX6O2rZycqwLysVbbgk41a0RxnQCkydbAu+9XU9MEbZUbh1eJqUstIKt
hRKYFgKd9X8DSk3/2uOZ81jlg/22tJxLN+bRnikAhnievkU6j/mPG0aQC/VMqTig
Nbrygb534pCgl5LpXvccUFDwOPxRjmMG1mQ2hz8T2tGxAvu7uLXGRz6+QbeLYdOV
RGUUzcD/4ETpbsBHB6UmWW3H0paxhyi4Ss4H5hon+A0OT+JUXKzYqGzreA7Cl1Mf
6RQZRizPDUOKBWF4CIfe9matKGilZRk3sF3+BwfovGHNwtjQsr9KWeqjuyQUiNy/
Sw96RKudk2F43j3yK8wbWFK56/UxRgDwFZWYum4TC9z2lCG2iaGacO++/mS8WwhF
z20R6u4Ikj93pPGYh3NC1vdOKuZShYNz7DDbE3HwXPIxGhSYywhOahyfo7aUxGQq
XC377SjWATUqiHkCZWylAW7kBiww0tCyOLDgPcWz1dF2bvpXhOL6UqzHFpKIXvaN
dF9kfPKn9WoyVa97IJWn3egPKThqZpfQUD16yf2l6vgAn8tF5AmxSeLU+9rtO7lo
0B3z/plSBYUdmQRryrCS14L6jTkU8jjNc8EbgpKQFcKLEaBbj8PpSQEFg4O3lMx2
1HdnL2cKp22rDjNb9LJ+tslgNH3pmA8cpKNLa4DzzEnBdda/dDjhQ1tg22gye7+m
yZMKWU8xQ+fRaEsM5s0zKMsAfd6V7Gyh9sYtZx0Xjh0L62v/TVaNh/sjHXYiN4Wi
XCImOg/lCWgm6ji7/o66vCRXcM9iG5p81uf5NxuwPiPxwE9ES7nwzG2RKiEx4VIX
36mPSruulQMT/hTc99uUn8UsKvkANAwKWsFcPkYHKEMQoTIw420eookSxpXNPF4W
1r/Kj8nGeaPRwKM5jGoEAWDXE9vOkEJIfNNikKCLybwGQRwuv2YtSz4GJKsfyRgR
ciii4oy9gmbdh4TJlUsxjrokigVDZ8eaxk5sSPu+TklmDq9GJSO+DNTuE4sSY041
Z5OTXWgYbHZr/goLkRdL0M5M9QA0yjnC8GWpc5s74YvGMabu9C79Vr8PxLW8Yejm
uOUYNU/fBGETG5QxNhWwkYzF+ZsMhgwpd2hZbSnnHcMfRtRM8AbSDMHKKEFgi79G
qyObCEEH6iTVtKu3Cv/xE49eT0RmkrraXzRsf/tu+axNXyXCSPMP8lzeqJLt0juj
CD9QVFPEnOOEgQmGAbXVMhkMgQje5jOKCE2kRgkPGL2Sq1f8eM+hrbaFLB4DUtwx
gqbgMDOzXAbE/j9lxtP9tcXd9hGx57zBzYGRxt61/Kw1ClrFgRq+pi99+FmgEkOH
af124rBvLZDXkeHmNmXF7xsDk1/u4Eg8gD4fSAJ/RVpjus43fZWtWPXFuWmkBdlW
irC6Du252O+jdJ81YjfvEs5sgrBX5b7x4p2pene0FsJDNdamKK7evELiBrIO0FhT
zEXVsRJ2dx8bNQ6aQfOUZuJupAruC3TnnQRYaEfLJhWsOwNK+vOR3yCcbWPpmsAO
kS20gb/YfOBhUwom5CmHgyALhxW9sjey4GPmZOfMWYDFYiI8nknrAyzPzIcxr9tF
Rl9GydUmeU5oXKzmPtYVhAaE5n+tYgjdflMqA1x3EvZumhp7OfcD+dIQOioTg3Rl
/tgWlaBDTmWJceif2xZNs1mZzHUSXa7nL+u/uvaHTtgb7gxzxWjJImWNcgVAJXDh
K0qKwSfFWo2AziPHmLk9Xv5pUy6QRUs4GVsvEjE6Jc/r4ncO1lL2YrizJ7cLD2Jx
rXDIuKurpLnmuE6XqGvvkrSDrKG9TH5Fx7NazKy+11vHTgtQPHBImj24/0M5KonU
LIAGjZKnu8vqOk0zFWlrzgrA4Qsgt234N19JRTiqpHs4PDTLU/eUvC7AjkTjcrB2
w6+PntuiSDUxr/zkib3nZobtnxpGidV8FtsDCHO5Xd/+gUNtcRBTzTwnbv49U06k
dUcJIxL616wBUKHqsJ6YNywfKPxVCA+b7TTpxqJ3skJBQSL/QYGDZHO4GlzUgy73
BFQlikqzG06Mq3blaSr9xULeNZZZ03cyT2s4pn17jcSq9oKjt9dFJxfoduNGo3+B
0MV6ATTkcoUIBHqndRRHiHtvOneZYN+IWO/5KR0jbgalqUC255eBMt8kE6TChs3X
hWfXEzcKJV/2TvcQhJAB+3mCCixluMDBJMIH/N5C1bbtSQiDFGeLzFuhj2424ZSF
gRYoaNEdajtbOp8CD2OvsoJD+kzAkgP+Tv6EevhDx69FMyEBjlCOBXuIn5Aw4uY5
yGlh2PhrwnzlGG6TvXK2dZ1ov6kMCph6UH9fXNu0Ildr0rNKr/o05AgaSX27sw+e
nzi4u7VhzzMBRbcfQmSIw3jgamv+d2JIANP5CzFTONoD6wMN+RWJp0s4LRY/iOC5
+9Dxv+kAVbGD7nrKQzUHmi6DHKX0WCDizZlotc47UlVHqjN8B1KrBak0lTPZwcTg
aBmF6NrSk0GwMBsWPAWrwwXn9PUPW/api1I1HpGyhVO8GORczGfP2y76D7pBfT55
DGQPXJ4uN6KcX4yQtlkCQJVkVgbmmCVd1HmMaQIKwNp7rD9a2+VGgwDF04E6Q4y9
xXy0iIKIOt013n6aLl486r1inyJOkcLE/dB76ZDluRJWoAFQcscCZ9QmlmLu7rbr
IoM5t4h15Imsns4BhhIb1z8kN7xsXLqyGnnm9UZUBuYy1ZIRq0Ye4/QY0XIR2Jps
x+B2U5E8E6CKmhptcvZzfWX0Q4uxkvvZPJIU1aBrRfkGzOD2VZ0D5j3ClaI8NXsk
BqUdwj1VyCKI4WFheVDnn26IWIBMgvH0sQOOxPAItLHxcyoG9GOsYczuqEX0V02W
Q/5uMtQntRDpNGwtbwkRqeuCyjyTIN51jwSwjYC+/AQ97qrREr28NJ7/h/5Hkrhb
HU/Puxh+VOTRa6w/cGSBAN9cuudCG1VEwu3cHMDS/OLvsVKjyogXREj2sbfdgWsN
pIfXZzV539cTd6DQLMvAk8UXKYIXv0wd/hxeK5hlmGtHMHKAd2SANDylMyWA9Rbv
NDVGnjbISpp6UCWlq180uk/m1lWDBwvJBijSaxSn+t9KYW1pCLcd3WJcS78tvpgH
KJSWsavFTAGj+8HJ7M0Sqiy78mFAb/KyfDBg5r1JwYMEvswVu7caUf3ayn5xER6/
YCkP4eXtDrKnN8ZifAAwRjz0Y5xJb0V2OFhIphesw6N1pDyatndf4BuhMW3GvpUc
JVTdZOKKfcQO5T51UDLkJ+rLXE2Nvp0c/24CRE78gh70/k1Bk5jhxdhdQii/AFqQ
s6ueNnuUbSIgFvYAjudb7bt277+8/joOhN7oC8Bn/pgi0XsauZBWunoUhWMkpSuB
5LEHZ9PPs0WgZK+I2EliO9Yqbt01rdjbDLVzyFBwCnjwahx4uTnhSYtS+uUHoIj6
Ync93IfTj+9RullV3DKQpL3NDvN4eLE1H5kCBpM3m+GqPTQQXTT9IWFW1NqaMmBz
kOiKqRxbQdoyQgXTCEgR2qahoS3/ItQjGqUAHiR8m3jWQ8RuBqkdr2aAjjB09yeh
bEEtqUmDCMtQ47Q5q26DAz0cE53FQCwS5I6t4loMDHY36ZmpLLMjwOvyFQx3yPJk
AEg6SlJmVDvFvLOc3NA5jGuflkno93z1WlMf5ObpsGfDYIGQdG8hMFxE6gLS+TyC
/Yrnuu2ij1EfdZDJxI+myB8pLYQhrpwz0VoXjIY+DSNrD3qCe0vocim7luLke/7y
zrnGHvDn7F41oCqgL413rgbqcExps+5MKUjsGrUj7JPjQgmBVjCZXTvDa/F0K5xl
1aUqKXopLExF0J4SSwN/IXNHud81kJYiyUjtdIT3vnNYOV7MAJIYzKVl8J0dizCX
Zkk53oTmMnX6mJ7LJuGQS5zMzMkEWJW38npqF25LKuZ10O7Yvo2kqb5gie2wByzI
oq/fFq7JaOzRL1RFYG0vlejs8L83R0ak1n8i7J4ENEP38J+OGLxbVbFv61p6OZr7
S+jFRv5k0rG8NuXfMQd07CgB7sdeZpswGohSXbqKW87Xm8C4u+iKXmXRHBMy03w1
ugG3OfSHZvtWHgPwKs6HBmMAntopIUHgzAiq7q63ipsNp2GZAs0PWztKuJd8WnyQ
Md9DEj44tGRugIGrhO1EjffVJALWsHp0nHqiDzM4S4JnZthohJGIuJ3asJ9owF9g
HLzr+KfGhnnPpJugZOkHPE9rKJ8lzWWHkI/rpXwwN7y3V50AcVycuPfBlD168B5i
+fsqIJvh8BuPmbgDz//vo6Um1l6UEeS5VAZf6GEoEVBwdRQak2PxEXnHU0qCD+pj
dVQMk4u/M5kgotbwraWb1PSO+SgwyDG3UdGtetqJufR5sg7BShprufah3db2PiXx
ez25kdK+RkL8LJAZ3Yg85Z9V/lh1t0gJ+YQtPQ5ACicgS3M7DYmF6hSHsrDc1XaO
B2TMmj9ok7J9T4sWeSa7SNLEgNqcOzz+t3RdldRqm7RUoTEYrCE7EQIW7sJLBoDb
Dv1XFs598lvu0bvF20OLlZdwfKiOLtxvRMzwZqeMirHTHGu71ywNq8TGNYJz+Q5p
lg3vcaUv2LX3dE3w1cxAewQHTfTM1kMn9Uo9Vt8a1HiwY2/xlWaa1JT75sN8j14r
JgNH3iVxNJI32yDW/IBhMAPJGavKkZmHluwtykqSO3UEqfLHCB8UJk3Z2juEyXre
vfzuHXYrs3QNQXPc/eJTX5hRn7YU5H3HWUeXnXnKpPEpF6y+/myl2/eXjpdv4uJX
Cp3EzM4fn0+sxJSrWRFXgrFMB3ejLIkeI45F9FcNZ1fNFKiaWHw32ByTGdiWLFfR
hUIvZJ5vGdBX5VK2yOeGtsZafR4vQwseT9xCXnz0M88xFLyw3PjUffQv6QPzwOHe
B6x34OGXDcOskTcyY4JPpyI6lISlpN3tKP4UK0SC0oHW0dwD3pKdEw+Rcpn2ImPP
rLBiV5xKnC93Oxvf05TaUdUYEMwQ5b5SOnGbhEEE0x3rhftTYvWWvtQIGCcqYnlX
6jCZL71PhyMZVkPYuZRpl087mrcLrGm0V55DbD2BusTH6T3MD6KycvqVGvrI/zIL
XhUEFSihi1p6jt8jTJUCvd+007pblILuUJYnGQdpbswrWvBLQh3sPb6g92Eg6t1L
9GzcTe+Xy2uBJnhIdzRe+UD+Zx3K5crGT+0h6+GBu5Ls0CbDZ2mbU+rmmwRvXgEM
WynCjFUnNmnnNjkYTIcZHXLMs7WJ7DLFc6Q794b9gMf2z/XwZbMfXoCkMzumCqG8
772hsesO27FxPCS36Z1wsKoJTiitE+HQKvrTTQQO30U2XAhhm8fb7ndE/nZ4CI+Y
AENfVYB3Rne+KofqahAu8ymHmgm5Wr/Qj5UgFz+yDU7SUP6RRuIpaAMhvJq8Vor8
1obbOkLiEFMsPFVuFKd5NBWCxuu734ZWnRiMP0P0GGb2tLp96zr84VDS1+rCUW9M
IOSP0hW7sjFaszQegjuS5RRA4KA7jaa7njGovtqqis+jotolZtLuQCnPlUBMKi/V
JMGAFOpkyjwbz1ClqU/jRB+M682F5ay2/TxOgLE4b364a0Ln9Njo5pUauq+nnWp9
8na3Pdv56JWI8BApWUkgRCPclGkucjlP/urbhXJLXepGGlokgBsgSagDvrOwXtWb
3G9sieDt6aBsy3PXLcy+hnqfvFvPBzLy/Mi5wtdmVAIxLlKQRJgwY+tgq0Ku0cgN
WBj+0iXFNxJMM8BXBRMpYvsNoIgqEAFF4PE9+XsiuvBp28yL5IlZHW+tEK6ohEEg
ycOPqqEqkLrFqKQ1YLMcbtKzxwMs/z9vKIsqOJRKjAJSw4bInJjnFk+3/TdsaPUY
vQG0camwXlMCZe9pzWr0D1FV9yTj00FVqZkKPxifi9QSoDFLo8NVDs1Xj3k3PUZ5
EBUiDUAM7wo57ydeQGMZ0pI1DRil4rFgyKtGBjx/hNGhRm2ciRQHFJVQPW55FNy5
jQlGqRHCFEtmGaCxpECBt3/Fc4GylUEkQb4FsCgOG5KQdh5enyjwi5LNGyZJBRO/
SYcDDJKm04er89zpZs8OirCv1nisY1rAN1l3YMRSOJy2ReB6oBPutnHBfpUGefUb
znGI23tPp3hp5/ZQNVACUz1DXRmtcFOCKthC8wxBA4uu0ic3RzlJ+IkdYTuEzD9c
S1x+mK8P7kfuHpJW6c5rgwibxox0aksmtDTl00WMVucG4aZAF4n92f70jqWvI0Te
Z/zXA1XOY6BJOYnXf7KtIYttDn9sAX5mCkFE/t7yeWOf927T6qU6cDMqsc+H63dT
OdItOnY05s9+bZiKrdmHxhrrVWw2+uASOamN4o+8gsRWSu8kxCmemYpugkU6xpUl
McFuMRYk5S2vIyCRbIPS1gEHGSGTP5nJlKp+JyGy4osWy4Xi9kPecy158RfQVO8S
TqWSDIYMkTEekWXAu2N3qAS53lEzkMyu5gBTwdTHYn56dBcueLSK1b3uYtFHhYn3
HczNmkfXpMwVqR93VNvXFRT9flye/dTRecTM/lCCCEurIuLTRapJFEDs2KnwtGey
quVSy4lHS+/zK2A7CSKUQ6SGNN8JOn0XT+wHZWj2gbq4p84p5PVzUczNhdaXA+lR
WljZRK5AVDW44FRBfEWhLiIhG50vtQjbWKkNQifhTgzA/scrgQlUi2ifwkJ9nOrT
ndT1pbO9KhZZfHIKlx8mxqAPSK0rk5xxzqw+pZ+amOG8N1V+aQXUxFThmV9MigXw
n3Yfjg/vaPbOBwQEvfllw3E33eeR4Xkhx8VCrhUGSjT94sKRIdLObeY0IoAdxmKZ
PxmjwDwPTlP74FuO2Jh5KFEMe41NzN9Y+KBTZY8cmcfhKZqeSoZ0DhOJ9W2BTew1
g1DAdg8ssm8Pm/1+lFMaEeIvGTowHg/F++Wy+gw3cXOBVoieM6S+d2ET8e25Ot1I
psi5sJJ6fJkhkkTFYqKntYT+V71pt7i8McAZuCXa20vU47hYTO5gM75yfGEBKsS/
wD2zbeV6oavVq+zlLFLU3GtbblJjbGsG4lD9e6uXx7Skn4LE0+7I7/btc//uFVBR
X2jTVJqQ+lvv2CrBYl/HrMMKuzKxbKEhzHNQ0KBQwVGS7V0pZ6u+ojNxKrooSTTM
BirreJzt0AP2B3yP7DvNK8c1GNmHVqoggxW1j6y5CXZD2fV5AN6SGkDVrhbE2F82
tFwmivO4gj1BrgB7XNaKUdsL3QVseXwGz3Q8rDf7l14lTXAxD9BDZbPr8AkGAdWE
wXeGNr/2XxzkWFvHcVkXP6TtReKJOKzVltBHMFvxXDLfdRHeCjrI6TXrx0WVCF7o
rBj9yQrlau4wWRvNg68wDl5zu4I9R+cM9Lkf11+iTtUb/S3Ayu+YibzjoC0iO243
KcuonTa8ZxECeQR3i1FfnBzzDdw85iQDtNoWKhCBJbwrSSKyFHmfZpKhF2wt+a/w
BxWLiCCDZVIo7yJ4Xmhvdz5180e7uKtZCTNjKirIOuWg/iGlge98aZAePeu50JlH
JcRwYEs3cImJubw71rZnx+kgsyVIZGd5yC1uXcQKDCDmlSWdkyaZfDIriM9kwoK9
lLwwet5bbTOR8HZ7345RX5s8n98O0Dn3qetUUvG0NOqvzR6I6lBsILajE4RSrhsU
QRrZmFMCf+jockwzsN4K7CLjDzeTLVNbK1hOlB8fJt+tr2DQwDnz4Cp7/2ARMz5U
8v5iQZuDHBkStdntt3/0ydJ2Np/WwKgJuuTegxaA78bMUjcQwQLqoEtq5M3keyM4
XB00KPT6w6EpnXInQmGwpUhpUWa5sg2nYP193hL3A5ZrDlwO2p6cKeFjYMQD6SNd
LW3ioQM+/WzD77U5lKmWCsqe1f55Y/4Iw19jsKIHTzAu5Z61qXyAmYad4Q0rfEow
lOUBrA2SYHt9OvM8ypfcbfZtTo/dMikQQqvU3SI5G+6lSVRRONXqUJu+FGSmiKeF
V2R5y2geu4HChnd1NMEaSD5epUKz4gvLs/vVmayZ1qYzW+GWSi2d+8J7qnItOXay
T7M9SQGSWTWLupQuBjkaUCgUe5N7XGtDUzoU4nMuZcIAX+syrGyhmm2ONZufYi/f
lbb1WBqqNndmAnBivIEgav/VOB0d0Km/ZhmvQaMmRKvzmEER+/9Xn8VRrgCFuwMz
nMnTXktPIIgleRzP3uGDtwqRMvHcl6W5ijbiDw4yS/ju6DVrdPCpvJMfa01VE+RV
BQ70sE5wmkxxLNRLgwEoXi8PoGdBijXWLKChQDzKoZuu7YYna1o4XWB2IurSHfqz
v/A4vpPlwWlZaHl1DFhPI+PlJOasuNBVh0WqOcm2PH6lpPftnX5QAoqueOqAdI39
zeGX9lGPasLmTMfjZaaFUkhy533lKAVpAiMIixQhXnTSI4aNp8Oi2s8+sozDGyMf
CDKof8rRpIEwWzVXF6Kd7kMwkRaBsuYlEMlec2i7CttLkHg0UDT5wA+FVmr1Zfxy
1gcWQxWiwAw8WrtLmJb+Vfu0RyYGhIu1G/50ML1l+A7sW9NdVADH6CShQ8WJOz1Z
WK6S1vkv6C4aJpZNJKriIlF4OTNLsBwjkwticTb2aykI2q/JERogyKIXXbHx9lk0
4spgOrvsZbFjySqDRIHn9rvOEimCFQvhmTdUALQ1sMhudnNUIE/J0PwdUKR2fZZs
uXfc7SeroLD3DFStl19shgXgRV+qCjGe9Cl0Gy7SHolQNmQv79U3Dp21JTlBeMpJ
N9PNT1s323fjqHDoJcJht2oOZWKzhUQHi7rtKHDdBDIuM/9qoQVbfeRlWdLm1GVT
sdza9OKsoP/6iO7bbSnjW+UAfZxtk3rPA1J72yO/ZTYjO1GT/1xPXVdKE1BdqHNs
1oIRVXpKwjv4ebDBoi9PNjlg2a2dM5hFzA4ko4NNnIw4VgwRTVSNMPAZwI+8tBOX
6/IwvFiItuzeHL6st0im7R3u6o/JxDAyPR5R/V0rd7NcLFjnk32BzFuMGZ+zuZHK
7YOfxXJWOELJz2Nhb9+bsKdJNvM7eDNSbXJQqzOhueWM3Bl04VUXlDS2yZkG7tbv
5lsmswV70RiZmaSj3eHfPQmu4W5bHQhOHurbBi69qn1XqJZBB3LdfxpOvd1jONbA
76E/0RODzPoUB6wlAPk+Y6QRuJ5gpwx8kYazhFWWTlcwJtcQr33QUCXv1ZJ4/vvd
S8TVe9dEo7Jg+Fpw/WuC/93xsFPUzU8qu2N+5CImH+OhNFRmjwrF8KzDnQNOIuE8
zKDyyfYHfMyIObuMVI4ZGsCdwKQWmUz7hSdSKLZ5Qmlvme0rudZGDMLT+RdvDhri
6O1xyxv8WtMoFpWwkk3Da95IgXry6eGu7lb8sDyd1K1yNEKYjYuekbiCYa3SUdld
RqjU7ipSik57bp1bdDRPlSAb1SDuFchjK1Zjhgib8aDhmhcQWFBh5n70kRKeyliO
xz7mNuL/oFm/33QQF4EDAjgENrUdihiMFOxtNej5eoVuDRF57n85152ZLdrf2ROi
5a8qeS52M56vTSJQx8UNkZH3XbG8fuWWowqS029h6mZfypF/9cbhOzY4p5GmgdRs
RP8uABP2wStWwk4wMdRVj2h+DfyGx1unYOBz89NadoP6s4U4+NuL9IentfZ14hlB
Os4qpgGXQAAuAZ4MzZ+QbJqmIorgRv9qd5qyx3wjOvZLrcWCXJc9k2wBCn2gsF3T
7vA6Z7Z/oPAPlxNru4S6bmcYbMDcyPpvCpBSItz+APEeaIFAcesNLmrVjUi+0p1k
MBpUSdMVcv7zjIeZ/UbuEvi8lIykuWwyvs2XYVufROuJlZpNxIdCA+F0Fs9/y1v9
6504lhM7R5XJajkCHw2Wji5k53joPV+L3mGSox6/Z57H+Ym/X5OBCTBwCFd1dO03
xw3B/9EpTevmLM4CF0w6ZOkGU76bQT06Dtn2xzaSrGkJymTR6TI2W6xwYBtqYGD7
84yNhaNcZdAlMiZNyQMoiAMQygvo6nPQ0CBrIe2Xdj5dx58SlPWcmVI8Rtig21OH
EtwQJ36O1TP1c0VmCseQ+lKFnS7auegChTM1Bi94hMvhzwsceA8hBePKO7AGe8Oh
ubiFDityOeL253x7cYOH6QcA4t9hhwg4xtWDbanbJut+r7QIz+oNNt/WwtYPNx9W
i4DzMPw1AR/9D7K8dJxc7kxnqg0icJLs9v0r/cT8N8bfLQn8Z87VYjh+i2iNPf8h
aa03SeWa438TG7jQC+/50ONCLIUvqsfPA2kteAB9o1QUtniD0byoYqEArPGZcLuW
Zz6Y9edszD+qMEy/xf7rF5gWbYhwXeVe0V4pMm6NLdNYLEF6C0HFDAOR0+Zf4RB8
kYrQvSMefMh5Lw0pftsXL/N89LYCT7XW7sMHH43P9HVjQS6d/JtY3lIHQxxR6vL7
ehTIdnVNHoR+gLdhZa6riDZ5DMpCwERLkr0ePKGVn+KVdw7dimeM8EeVyCtOfLJT
t6ZFs6DOxNzVOExcXqWRUhfv5WPm2vpnSigs97+8N5sgGunmzCr3KO8WpAJ9mkUg
1PB/fMLLxVBPCNiP9OPY4h6RpHtZ95fCnz6b7ubVN5R5M5iz9FF9Di60vFvwHhkn
dGRZKLQOlFFZ6n98+5XvwST+ewxrqVlcnt/yOEQUEbBp9LCRSV8ohakyO9FHA5qZ
2Tkuvv4ac+q1EyS0W9tv4x154KhSEHeEegI//jjBQs7K3HXJ7xo/RAUHmPY3cn3c
kH6bF+LFl9nNbV57tUKR/mqDsHfOog4NvJUPnXFCdBwxeTqxLKq+M7Mmfn8lJ73d
YO2HhHqVavnuVocbBs/mFFYD2SF9s8kz37pU2+8zxxrfCMgf3O7dMzAUUbMPpAyE
dWNBjo6kTALmW45q6F2sAOO0+/C6LsIkV0CL0Tx2yGjUR7MTKviMrcUoaNM+Pd6V
oTYGC1JgA6C5N5BAI0QlT3QfKoD5DHE2WoE2DQL2CsOZaBcrN9BBTavlPaTbMw4d
CiSP1zbTVVxnszwXoxjwjL926bzVuNVf9+T96eG5778hotBUKgpV2JELVPP8/tls
5eyyS+iXYOhqsUSwBE09kQ==

`pragma protect end_protected
