// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
j1eyTRh6lGT6yZI93uHp01/L2RXI7+A2p/6p/LbdSjtVMFN9Tl9bIW6J3JoqDVvl
+sLEHQosvxpZIUo6GXvk0m/V3L+EOPHkeu8vkm3Sd5VD0kUpnZMtClMwC3b5kAAr
QI03LmUsEK7vslIigLYNkvEpwS1Yu+rbS6hqSykQUKo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 13248 )
`pragma protect data_block
EThUWvEaEnd7dGVcidTeUWqXxMN9V1cA5BJmHImlTnQM7FPrqhHz2gZj4OGKqHcR
G8SjYbupN+CH1tEmZ4m1tQM/mccNKqRUDesbAGUn1CyULf3AVOzn6Lk9JnxakG5n
tW2KHDlJNnGVgFdDHpxCwzhvH7xD9RMrVcEf8uOFmblKeiofeDaospakdSA+AMJ7
EzQnq2jKD0Jq9n60Cq+TSaeoBZC3Egt6pMWLIkJBv6ZNYGUTr0r9h5iRuO+gxT6K
HJYonMSL3Qi/D2HaSkCRyLhXQ/Za+ij9SRezSsc9tBX2U/wJj/Ruwhpsmtv+6gEw
LEAGTTpzQK0TY3pnu7VigWJw2+R7DiapL84+qJ0ofOH1ThKvYvqIoAyxONtiivrO
URxdne5Og7dIKsoThu37aeErD8e9otzEyQeZfbHcxwm7LLhdypnqtTeL0//uJaw2
EXk5Le88FxXpD5T7Wub0ZUQrXVM48r+Wqxn3AeHEXEiUDPhy/vRRqD8WeBALp2FZ
pAWhnFWCyUyqYRBFKpzOvg97lopjAd1nQ2vNjLfkUoiWireHVrX44UMcozkA8Wiw
0ZhVdMTvwLhAhCcZIV7oTzIdK7zSSHE6G584OhwMWnzh+JSFHnbz5EGannACFRlh
bYthbLBkKprNYP1zJoy6d3w6bMyilwgTVTzUaBABL4oYhX9CvdsOfIHxJNkx54bK
HMII/OJoV7TQshvZGcLCfizEGsR4J4wbFZopGmipCqNUBqGBnZoeOWdDiLd2Yg02
1Ygv0Dvco1hUQgb9k3El+aF4z1P77Zacwmh8EEbpZ64rzkT8ZtWgtgGoJ8T4a2gu
3S6uFWgpvclXLf9zFltjTdiZJ2x0ixLr2qkzkn/8WGdEOCBw8BlUU23htBa4opBH
3qjVc+KIQzQf1HLESM5AmtFNkEyKMq2wzAoh4oL/PAL7SZKiU6xXU3FcqxzftE5G
wgUfbmut6bd3YZgeRZ8GcL5/cewDp/4oFYnz4xlGVbJcyjcXnUYI8ELo8RgK0VeK
iAqQt48xtG07UhSwJuyp/J0uaalypAsFIoPKsyjnjdcRj5/Jvm7M3bjBcqoRbYde
kQlFG0oQ99WoVt3/Y1ubb9xGUhql8OHlSJIOb2FmIIctPuXO7JyFwfw+gw7D/nZ4
tDwLidiVl4ItYgBnRdmj+VitUI9Ct9215jCujDa/JHSZBXnIUn66zAjid0yECCFN
hj7GsBlJurPYA6mtuST2IOcmt0k4vSeQx4xmacqVfZmPnMas1eUK+ZDUTTbsKGqn
awUhJTJKDInk4V6g2Zpp5DYI1NQApYLM1UgQKRAQ41yZkPNJ3DN/eZR7mnGoo4ME
LayNVEHqZxZ2t7pZWRBp4wu4p6n7CsKMDajDT6+icdCcp1ZVfGGskB9FL/vusyRh
sGf5aLkfJnQ7kDa0lG/ORd/SQJfrAH8Cp3ZdepwpuxwlnSSitCdSunI5ipef4Uip
SSgIbKGxJHnJImZtEylQaHDAyjLOM0rc9AQaNZm9ggmZiE2QXd5tNx42CPIp9OwQ
UKGM5nZ7Wi2QCsO4ajwXYjG85DKil1v3HAZunEq96anWIqYIowRg3V51xJqKRyVj
uotgMF+ZBRWoYmHkzAy7oVz6kMk3G5oqhER082ZjUo93j4/a1VFmKstfUcDhh4rk
bwt2NKkG5DhPtxLfEZxhePR+mjR+IUJ2S40ROCYjBmzOAmDj90qPZM4NvmHTM/fM
dGuES26OPI5FWpJissYCIZFWP5hvOOsYSnZ7oVSiWPvTGGabiAeuFQqDUvRAWsIk
kYOWg56vyF5c9LA2ohh53Fohx45646J+/9mGXPIdKaiBXK2se/saJWWRFXQ/LFmH
U+8XlfPebAzSEiXfvaOoriJEvtXtGJnGTJvPiu/WyVWv7zS9qS0jkTL/xtYDmrTz
kygIzN5/kXXsCkDLlSb756NIY42Ajwrj0cYaIK1cdI34LhP8j0s64H+V8DhyoUIV
A3k44J8KnTgadrRQEp+gkUylCrIbDwoOuLnX/7zf73ql8Ae9ptVB8rD1d4UB2CzQ
V++0mxiWeDdrI8VTPCRw5M+pLYvvFusL75jNmBSuBsQC/gpppIWYNKo5HegJEBHC
GNUlTyFk5Ehwdx3sXv2S0p8lbjlsJTCITwnOZxyeiNPtXY7/7fvv8hOgjmSGqFh5
VUORsSgmXm35/7MEx3jZUUh2klvbrCnBo8E6yz1NWWB5hKVKBDs7yvHg9Jkfn4Mg
/KyyaGhOsq4eEgYVlCsp5RXM1Y1GOd3AHnwea0yCBdssTzgGBR45AG6x5zmMhpir
OVKEXGb0TNOHx3QcMsKD2gSuh65Ls3NLx5CexGL2fzB7yhcnECF82Rnzi+kOEqb0
i5SvtDotN7OkN8qVQ1HS4xN0WZ4jWH96P1N87E5PJeTVCs4/O7ijwCWTZBtOVlgD
RHz6HINOX8KdpfPT9By+NUIKMMJnw+6st0DbUrGcQ3/y6O8yv2Sux5bwarfHsymZ
hlJ6S1dx11RL9/8MMzzteoiUZutyNbdah71PpuAERRT8pnEoxsYVBN55S0puzLa0
nnCOQVqO9qBwdZ9PSXF63v9+S0EU1czwrGjBDf4tgXojgvbL7KGeR9Qb59W27cu2
J2PSbSDWOsFOOtAOTafR5cOpri0ofc8Orlrp1WsgQsT/Sz1gmEXyMmQaVUxaRoCc
ggIKCi3PNBkXIA7W+SzkRWSPRLmR6OmGABsAzjc1VtKB4cCptw8WZKVB51eN7DHd
20YSYUgAwMJFdLNYf3B7XY9AnYPHXgFYpaXfEVvxZABGhYrb6bpCarD0pTC79Q4D
6Ft72NSKwLEhm+yn3uwHdyI2xTydGEDv+vA3lBgKjSFFiYIzG2sjRLx0n5San2zQ
7hWC73fm6n3o1dmTEs6dC+v7cH7tTjoSt1ghrihyvFLY2R5pd3EgVNpAKMz8IATR
ABpjd3ipd29EwI0+EiacZfCw7h4whddEAfV4yutxstrdYrrZlKW49h6ZMyQCJ77k
pJATrkKYkl+Z9eUqrTAPkwOn2EmACXn7LDCyRP7IatHjRmxYmhC62jYQ584fL4nk
hNorqP1KzEza9dALVpu2pvDlmuftB/HTSsd8+fPgJ4MfOCLDGyD5aZgfFH/3Kbzf
eKF1xTyzj2JxIENPjZ559OT++Egkp5dDQpDdrxAgsJaTFwVclqsWUxII/pf2/RUV
sUcJbI4INXyBR/NeGmWPeo/7/ddemlsYZWD0+qW8ELURRkgkRrO11w2GUxTBm5+P
YwXxUCR4nlK47x3mZgoEiiM9RuJYdRiYO1eCUDnpIXcDdn1easkr+gRCNo1aGTcQ
f7220X3hu6gxnilNf3BoT4N/TjUV9UEER9aWydEvnWtNPc6bd4SdMIMhN1AOIxVs
+z5Jbi+f2xm/2qUkbshLTQrvwgkFSP+mvxT0SI2ZGZfdx7O4eBw7vR3akTvL4ltG
jyT9oSjQ9YcRHoAs897YU921CHP510uhTqhP4YYSFUjlwFv5ILtNL5MgL2p/KpSE
f0dWvZy8O47U9SBhPat7JfC6EH8xdldH8MtFUW6i94o44gRdnzeCmD4TeM5FWCu3
8fG/YhQgIOatged6mp963TCKsyT6d8YnRzlmFuNwThrbxd9qie7HW4i1N7L3Y/oZ
MTUIy+SBsFueSOVYgpFY9PG9lBdD6BsvpmW2WUawx+dSr4B66fyA3C/2igBmNeUU
v2uQAgft11Zo66YfNJ8dpyLLoOys6aJ3/xgrPlAOzEb0HxIj2Brq1rFmRGoEbisP
HGUDcqwWkoocjqqhb7gBJltcFWhVRdDQC+x7vn5BG345syTo2sHqKEHqRNVNV5ps
S0zDQs/PjWG/kyIBiGw79wnRMWkiiarzxVkbc4zqtV3R+8ZkISxsEl2XuE//19xC
16EQHVBQzsi2DcdtT2YKy+HcA3os9x+WBLpRQAADOMdB6lTn6SPrG4i2ecl1dVOM
OXhvo7QQ9rat8kNyKWykAtPsSWrN9Snx8zfVJtIwxVNovNbzbnrkLQH3cutXm6Jg
+jMy3p7KKIoAh3DBnQvs+aLUD7l9usRpunhZ5b3u20Cyo2+jH+4+Zfb8qMsa4SlO
oHCoeKAWNkhwNUSsWa2bxKwS1XACDrtaCDCywpgox9BmfZlKK3OjmYCsukrGH6JV
/q3AMhqBhm7Y66MNQYoCqVMz4ZYRdHBfh1vhQp1JjkdWL0DakKaWMtaqR/bKVSnJ
80u3qbfcba/d0rqQKP2RrM0ZnYXObRH0I3kG7kfgSX4JDqVMv0ZoHOVH6DWQpYo+
AYN2I0FoBUNL6ciorUBUAIE9FmMJ3U8R7HvzM6oNUPzfaPYcmz+gzgZmIbLX109G
4lU4ipBwmtqbdV3jjcKWN5+WV75o8Kp3Grt/264nBQi8mRvR7MoGVBpHP4jJpHD/
+JL6Wy4kYewQfSsgtsiJiMMW1rSdUv78TtjxROFhbXzw0j2C9rAiM3AjyFI4lCO9
5QM8Ibs5OECLlVd2tq9yLvXbkJFUkFpYMK2aQIAF1oYEH/ynbZuIeU+OktgtczSD
4sJaFRAMst/zbATLYKcTPvuKNdQqxFaGEcgmlzhl2Es6NuN9T+UVx2A+aIfeOZW8
hM9toxQnptg3AI2UNBXWUkmL8LyS8ocw5C8pan0sOT2D1nibYHpmjTHUKu9O5yha
n7J4aivLPRYV3qUU++/OlLIvOt+mv/6wy9jdxpbfTaFYsX39yTEV6TbWz+bzq8rt
MykhiYIp0Ww+57/svc/n5VR8mPt3Ioo3WujO5BWJtZzIECg3K48HDgr34+zR1unW
0qYVt4VuMkPhbKDimrgm8PacdWlZhh+AV7Qau4bUiwdwA29dtkGJZLQKyIYPkfj4
AQPzk7gB5pOS5yx3LXsvFuLZSkv+XnNijMpVzosOd0kgbLBV3UU0HQqWBGe4PFJM
zkkwaZtiM9Dgg4W02Ap/OOJTvG+4hKusOIEdUat8L16SfJHIYjXf/J2L7WL9Ll4P
nc/jjhTC+WT5bC3v3q1sx6lCOId7oRuCXWLjtA5Antgil6Ja/3pipJKhPFhoJhFS
pOrvo0kz4o1zehvMl8mlFDAQSakWPkO7JvaoyOncjqvlboNg3aQO7w7XnOWwksDA
HdLQdweIMnA+yjkzSUiNVlxmKtgvCCHQWfG5PrskaRTtDEtuUrpDnGlYzySUbr90
yM0uaQvgbo7EM1xIms9RrnJ/x2IeF35u9/hKXopgSDgjB0ouk8swPIQ2rkSYWuhF
ZLQeaGtPDcQBKdlgH1gnV/WGlD78mAmHxqGArfGClGP9bLeouAtLTpMdS/SotK0w
SkbYCIUiF3SGqe4q7EE/MzaTqBOQk3klAJDVVPl2grm/uMz/YxIR59Rbjw3Q+dC8
WH6KLhG3uGCxFufugCYFA0EyNIMgy2SnkG1Rgj1S7CERBr5amSzHrWiQ9aKqZ5Gu
eTgxlIrkRz08EUP3VN4zfjrqt9jETfJBRXAml2nrJQLlacjAl3sZwGO/xMVH5WOK
p0vXnMAfI/yQH9k92egkqcjJ3k4De3uAgIygfeJPWZxPi06fBTaVSuxF/HAYzK1z
6dWE8sHBC3wC7NFdP/+jF9eQ42RrAWl6xKCRkYxqE1fYG67R1WgWV2teu5U2/N4b
MmUvuqQyzChWWAarwRs/DZvw3RhxRwtAXZoA7aq1+6/NiJ9DmqGwF2ZqTGzTAAVd
2Oht6EIyEmes3DID5bK2Ta3+0UHNnKS28pJcH6787Yr6M+jv3XZ5G5m53zTocATs
8gqWjqewHcHpRl5kGnm+qq64yFaaZlV1iXnuX4jD9Tfc6kX9XAjOihG1DkVCt21q
T28K7yfgLcqEgS1q93NT7nOaNcZ5ebxLCwzRX1ahT1+3L87Y3fD/zq0IBRHutIWQ
6MQR3t1j5mziTf606MikGVXfdQHmTkCtsqZkHXWwPsHAItp+E8RnZoP2/RxkklRQ
H7Re6TRWa3MBZhlTynTu9w1n93gQfPeNKOEenR1bq9DXb2zCIazPhuKXV14cidfP
0EeBbRFc1sldI2Vmsh5pdbybv4N9yAsxaQYvgvw/vWbdtbypZ5pbpERNj6oeC8qb
44Li+5P7DfgcymfdlRNxraZnWhB2vnF3e77yB6ESJBKV9X/0TTh9vNCpA9JrO9FQ
8n7qhskcsy3ol3X+QMJobnO64pCMda8aMFsa3MiPaYf5fG8cvfbAWuZp3enZvnib
Gt/viWmEtOosb5g92t35oF4VEcIJmDQEkXtk3BHsAgCyz42h74LP2vINHLeHr/Ez
M2R5dlGJ58qBTy9KGAmB6VZfXsBVhOz42eSLYyElFFFKCWk0YdOu7sFhpoR1LPI9
+oGEavaTx0muw9NX2W5oYcJ+o0hsP1EFW1YRbaUknefyRNsqyTkmJ2HS32mYjRW7
6W4mEWhl73O1219MlRYkqn9o1SeibdKxFc3ebyUUpgUhUxh5ZiWaqWntB+K+gU9U
oWTrc86NNJHSgdkpFvDaPph+oTwSGyDWjJY2A2PMrtn0WjwzZA0vo2q/+5uYB5PP
nUf8UPISUAD7lCj/bSAOCaum+t2wptgz02mNhXlPzI88To19gODMXUrqqGUq7XeF
YeZ+GfF2TA/dqjA4swPWag+NLaRIxjYxAttleazttRZ+5vI+yTuyUEvOC1oMnCZq
a76NdgFqZhzboifQdFQZ09P7BC2IcskWmV3/naTtHAlcl4D4FOc8Hqj/5yV7nj7/
TCii8YaOq9yCV/Geh56cORWRw44kXCiFLN0khL7qPqS6KBMYb0d4p/Mr2O2cqhAh
XF24kTPSld0TRpEYhEOAJ5N+C/DUMrRmtArxLN4EI2X+ABCz3BoSuZuB4osxz+9G
yKuo//PceonuERxc07tyN30yeApQ8ZuyeC3NlZFFWAQaYgPyfEKhWpxwZD9loH0R
Av/Qrzd5wMg81P41oKfjFaPIy50JFchQK59pp9lHkFa/PQ6lZGvCShYeF/ADlSR3
dXFeFxVjljdaXmyERyd7mv5iLL2ykMrLrT7kCna8HTK96KRxCEISC3YT5JjqC3ub
1VJdkxmrr82jSDtEzSRpOOlnlbtn+XfJlEgi931Acuk68bWJ755/Y7yf+YlXlA9f
ArHafkRO+1cMXFKtzLiWd7xTYDSzgEZxvRGzNJEmW2WxZGVQikIOFfJ2w2YGmn51
R6VV/Yh737XKcM+bFnDBbWHVva9pJW195LZHr49+KuJHGD5s6PSzHmlto1OCeRdC
qCQch4ezoR48b5o7KXDSvtzFwuhAEq+MufxOOiQINkHFUxAer2PzpcZXP62cBrmU
47sk+Rd+AHZNhw1L0e+L+lQ58zamW+pYIQc2DeVCJc3YK5Eh7vIppUhIowl696y2
pCdiezMAmZgUZ+9XXiNOdUEfxcE79aR2HYimZSiGA0O2qH2CgeD6vasX5FtPtImO
20ycudIN8pohPlM2pZWawWeREksi9jOBczbyY/f3pMQ7mXoYvjKEjALZhBNXYSJV
7causPBiVC90sZ4nMhGVdtDCUqWHSo0BHS9VsyvqY5ZGdJ/rJr+TaK9BT1RIk444
IGGr+1PrEWnWqTOPgez+lmA2NtRTjQqr4IJkpsGe7FUaYq4IGFmjMprio8TeMk0v
sw1i+PiaFNUvyn1lJkFSHJabZkujAQ2EINQeNuCK3UZB95Erl4Xabi2f3FXoyrwz
vmirWezjcdzmfAPvundDMOr96xhLN8GCfmA7qDwQDTJbZo0oSSneMungBvYOIrvm
8NJWx7YaaMStRubgkRmQuO3zrd7Q7Baa/S1F0qHrnMfXUUESdIvVft87cI0M04+G
ampp9bHr8zoQ5HBHyYOcvTwHRFLiKKTeQZctKEdi1S8ObGfz94M+36cothjnOvXh
NIlbr3lP0TNsa6xYcu570Snmsyhqwgi3vghNofs/zmtNL598pgg1Hg8s0iUAZ+mV
NLjsSoHb3N5bpRp7F+48wWBh3eEGTYjWHqsrLhXw3JoWUmj9FxxWxKm1OiJRXdue
lHoXzjiJxxwNTMmBI6JDWGHGFsPUfknKMgN0bA0AcpDaWWvphW11Z9Z+kFxO08gR
mn96ZjEhG6dFMlpN0/BtpwiWNlcJg/GSzYuvMqCl1ztbhNTsDfKordR2E/rswyYh
6o3fx2EaFFS4RkxQBRq0AQd+zf0npUDsdJI2NgfYxiNT8MBxxFkHd54sFcJgglN5
NaQ4TIlMhXDHO51lRihWQ1bJ0CgN+sQWmuO8oPo3HFraxQ2v3FFC8Gq0HqQheWcF
73K1I0600j+1VKTANY3535zMNiQV2fAvX3Kcm8HoeGLymkBMhI1O09pL4FHfVq7u
IDGRoxKV1AwNGRj7O1L/wsRp4nvc1larnqbgf+vjb9DuAU3kDY2VEwdh+fyc0ncQ
Gs/6Qlp9fqGOSUjVmbpZLmb6QG5eQU3KncDKm/XYdlR7wxuCm0vuNolPY9kNjPSm
L05fapajBHktYMhOJY7B2RV9xDdG9H85vAPyef1aRQV35vHqvJCLEnIH8kH2CwGA
xPK8RDNjxJXwkAVVYDfHl4r96rdl0g8p8I2otvNy/2laQqoO1+rN871zXc1xKdvO
t6AV+eaU9ytnEoZ8f6lgCLhwAEk3v9m0r3conUswLwzgo8y1Q5kUrZVEZRoUj1lN
EOYn7+YSC+EO90Lzcelkv8UaB0e5kG6ZTlL18ShIhOwXKEKP0fh7rhXJGhlWDjlc
8DbdF+jf+ji/Rjo+9hbhmpmWLO+CUSL6U7uOfdrDGj3t43vw+lJNXPPfHfu14yE0
XeoVII9qHMt6hneWEnSutLAN1OzqzhdRDRz+7J68cPH/37VLqcxTMyU1+5M4B+nF
e4gwMeSLu6QiFjvOvbwpg79FOKDfXUwaBCevuRCBiKS3qMNVGGc9wyNcBVM8xqOp
UmrmqCPxcGYFTOLjN3zPpFkYGyMwSJIFFEwxXY+xGUa7DSkUFA3V3mtjFSXXKTKe
/cqVZ8fBbbQcSRFiM8ioRaLDX6byjkfpBdEDLf/2akHSyGV/+H8aQeN+EV7Dx/PJ
QozOM8hEY2zhr61mMIVNWRF9Ac103UwMh5w1otX/NAVfisbxBTCuyvXwTcjftxqW
wY0/II+tvhEuu6lT5cu77vXvxuJ/TwqP/cQX/mGO5HkNkaiZwBFK07D0wM4oz3o9
w0+SW3txGGKQx224DUvJJg1t8yaOa0iG30Om9E2utXFL9dS/QZgraw+dobf9/vf3
Z8CVo4rCqfvupc9vsdIu8yi9CtYr4PvXViD62At/JSHk1u+iLXmRjReVKFy8tUC4
npalBXqaHKs3Qvdr19iTp49RMbKImSxgiueJf1TAmZveuBR361RqUq0Z/YOtoVfy
vr0WugDWlwKG1Dh/eZJeTpvc7UHufJmnMnZ+9WQ293NXqfmKmDKyxzmOReVzIXz3
qMuGGdw0wo9V/L4f2Kv+IKPxYgKRnpSc6NUlEAPdLkyeZQvY6bICs05rNoC9EkDU
sWDdXBhiNVb3N7qGlM6D9ktnGMwAONXgiV5oadn1cGClL9o0uqr9SYq2H72KpiNo
QrImSUxBOAljkjuUDfHcBK3+Sukf9Vv9+3frqJWh1ajlUG1lTqntRteOxsswHk/T
JT+gCqxCAboin85ogyQhmuOECUDZZyI8AhoVWXY/eolfeEqX4Oi3CAPRIP2w7YMa
hsVCCu9hsHjmUdxSzgy6ePmBqpqq3skDcpfzDgVW+ayq6ENF+dpG1UUXI6oCuldS
ECIVMkF9D5o+kJhFwClVSdzpkuNmAOKOLnkm98EjquEljIWjS9ZyPMIf6chMkIHd
5meQsvU7P/LpZxcoZ1APQGO0x2YrbDtHMIea1nojprqTwhgDdEuMeJXvcOYkh6KY
uQiLq7Bizg9E9juPeMhDybF6WNk1dSAYZR36MDDq9tZaG8j3h5C+KuwiUGHGlxrt
EMJXWgiP1qpD8Dh3oftGr/J5uG6D3QCOn+3Y9JbmNTwaMqrDpQqQlCMTeNASinmI
KswKGSFZF5Prz48MDX3e2vE6nlRn0Zx6tMai95k4FjbziloD0vkB8XTPrLxglL9d
cUhqYxBPDK0qBMn/9IVxJbIDwlSZFQfZuLw3T7bi9Y6Dsml7WQxaGYAKFIJUtImM
XmtdjX9NA0LGKMslMKSi9fB9mUj0DWqsSRcF51iJPF44UZptHm/wo/CMwwl+wfhX
ZE+td1GKYeTttD/nkyQx5fhBadjuId2EuJaqMBZnaRUIy78ExII3XDGfHt7sXNyA
R5bJhlZgTMsOCjEV5TFcg/yGFWaIJXf5BCOKhdhcIBBDLU96jNc5J7w3jMJEnstN
mqhdtOGCANXdfYNHD3YX7Ja49Y5BuO7dTSGFNc5aC1253TuDg+L7BgCIbwB7rC1Y
Ah8bMkNLCllbU7Vb5CHqSKEMJYAZQutxDVYaK0OzQ9wb/xMJb753ZLgRmZLUs99d
z96k1h2rXbeWd4C+patnc8orZHgA5NCvk9IXz8smfaKh/JGSkmak+dTPkY+kxzm5
ZNXDo/MdgE4j8HJq5QO6lG5fgaRbEXk2tD/5UxDETn/zJmL+5ie1kjvmUQQOjG0m
APX6SdxQfxoBLwYX79Ux5nFaGQ2UqKv+OufkaKtjTbztaByBNhizmWXPPVEBg20d
h3KZ6Y66/qNnvdsax53C53RrGKBerCkN+pzYOXlWLtIjqXiooQEb+BgXZ4zw6Fuf
JsOVvG9yH7BTLNvJJEi1SYSEM3RwrKevzS6P2Rp2tWv0b3ODJXbJmbHlrVGa/7+x
g9mbQL1rBWFiatgwaa77GwTiQR77Njkvk0FR8nZNEr1k4k1UGBeY/9sQyqKytGgB
8+p++u1AnNuGBUg1+Q76tTO3F+q0N+GnQ/dae8HtBMuMYaH+aXPkhugCYsvFNlCX
90DLO9LTdGQyE7Zg80/U6T8Xo+j3c0rrTk+dzCLcEJ3+KTDYSXfhD6l6VrEiyffZ
x5pKIuYWbHzwKknY5YzHApWTEOShbyDTP4aF7p9COUt4BjHQdJjOHhVhbXyYE/f+
lcADlR7MjeU2FUjTmcoG6Ilo9+ddkjlWyxAAH+YWTTGthwWPcuapO0x8brWrqZ2R
5lLilaYGufYObBdDEVPeWbyiYRjXCPrx06rt151QY/jCtl4teVf8i/KcWOlMAjlU
ob3CtqaxlPKfnfQI2eh2xUAyQx77eVH8tX/aBz91nH8oFb0CNy28pzDJKJl0+ggi
sEzd4zkPdSDu4lCmLWw3C9YZuZWtC52QL2Km6rhlp0jB14fp5Dg6kGUJAzl6zD6g
02ux83j88kppOjupJUDwB8QNoPFSQglPPMQ2Q/t1kW05d39Wno8++eSOTh1e2Kpa
IHEVnMmlVpAYLNd9RSbLBLB7cCt6Htg1eFIsDpUPC7J9eaEof6yciuNhwkp8WFV6
BNtWoXKfjYnGFqb2SP/fytUHiI/7Wll3VfR9sQItOvIQ4ZQLXvi276cHEOwb7E9Q
ryhKDy6VAeYI3VFvJgvbNhXchj0r7DkVH9AluqHnHugbui+3S29nrXLvc8kR+RiU
ZfFwA5tSSKPE/kGgsepmV2XrwxLqfQhZH7K5bgOCjIlPW+4c+k2My4eu4A/rWtXT
qp1mqTtd7RBX+Ny22x/Ve5/kHXrh2gUkj4U5RY+iT50SJBhcVVsbN3iFDloGMZsc
X1c5iSZXiNxMMEOC3paEVw6Sm/7GDt8BmyFRsY+3sbaROXP/HkZ9CCmEVaNnHrbS
Am0Wy+yq0nSYbEMt8u8+U3V9DUYypr7yHLtRJs8a54MbtHWdVzSEJGIJ4Nvd0Saz
eZ0BP3W9kHQT7kjNwljeWDg1/UQuSsueVZ8peAkxpUn0TjoZsZ5Ok5Cz8fOZcsme
4j3dhmwVcmqcTChJck8yM5z1RuW4VGy3H63V1BsSAK9nBskISDAmxx4kmXHQ+9CE
jjg/r6M5N7JVzWHcwdhoBB8OgIwlGhCRhRMPu+9DMD3F15Nwci/G8GAZzihshm6P
saXt2yOcWXYyWjofEf2XqXlCJ1dllCpHNP2h7NwiOGyyZklyOYWCzJtdDyR/TGcX
nvxCsT6r8BDKcpVpe6E5rwrQc1d+QaGc50fiDJveNOz/No4rHORYBPNo89JcyVKP
4BkSW5ZVd11rZGfZhmmRkEhU2N4IhiX93E/k2L6uPz+N/RiG9OqNC/WSFPrkbSzE
kMyio6/pilppUJBNICwArBNRnr3Bq/vz+wr39TbsACAaeXuyVxkoiTANpPP6GDXl
4Q3L1o63qcwwZe46drC4KrebCD/HLMxSXcwFL6JJ9yLPLSKNyASPl4tNqtSL/s+F
nEaXQje6sAQRKHT2uNw3VyUsVELj90yWIZ3655OFni6Nz/uFMiqhOKE+EIGOhKp/
0zZgVbFAR96S+k6wJPtZaiYTS6xT+8uB8Sqq7LJ2m3cDb1fRpP9qSRj5XdEFIffR
XpO6QgbGKJPliasmF7KJuEI5/sNb/F4tKrRU+QW67rxo/FVyF35rikP7hhi3IQtG
6R/AjVyLxUcNLqd5NaajbRS3mdvbX3SI6UxeEjhn3kDItP4v6R5P8SAC2OHKB4zO
Z7rYcZD4i304Y2jspssSN1lIQdMzN+y6yQOz77P8pXjID+GwBuBbOq0lIGlA/nc6
UuJDtVitDvjwMg51A6gDEaSTVeub7KNTpejaNPbOvVLdSZCV3hTikRz+TTSPnTs8
2JwxSM+m3rV+tXWW4z4zHzX5X+ZYIonn2V8m/PAzP6/MARVBmwMArEx4kt6kZkXv
jGOWogBTpoLejS8JdvVw6R1FTmmeOlhTBikw2hcJ/DErMJkl5HaoY0o56UlG68Mn
1bpen20je0VbxvhiCCWbMJb3KQQJyXKmQSXh0sbA5Vn8u3HtEGVPBnlPzPi5DMeZ
7kZUkf5n47oZ1LWYPVQckhOiWQoX6Mfqz4k73w8P8LOFQN3rZeuz1Y02iwlcbIxJ
EfsbDZyxU3KIVEDX51HzfSGwfYcZNNuEUhmKGbgD7u5+ZnNXB0fUfr/agnOMa7Z/
wq5cCFHcAQW9JpTEQwslYTx1TDmjsFwKTJtXDIPbobiHqZ0ELw2fWEXApeaWKQSR
KlETYSlZIKMY78WgufgsTt5tZqaXleARXOUxUb1M9Id7WL0ltdajKTAyekH49Z0r
pTgtUM1SA7BDxqVSR5u+lg04DYZFG1osduf4O8OlGA7WBRxuRETZgUkpPit6+cOK
0xveXH+09EojhUwHYqRg7MU5kWfT4FmjfcC1DDbGvg5RCAJCGe/qMKlgVOHme2gJ
GPn6CS9gWnheULEz3LQBAUSi5choO3ci5ub9v8npsFy+pD1Bk9FraJYp6gK9ctEK
mhnDrhBt8740zX8x1Ef861f2J01glXEMQgFDAIk351d2lHdFxBshTZiizQlb65zo
7N/7Z/otqu0a4mUnGHOLI3orzrTTv8jmu7K/xhfJ2wG3STfFmyHfkf4EYLHjApvo
W7JVE4wNr4S0QbBfnMPClq2XtTenloH4MNojrC2hK15jQ7JjgfnHXM5fdZQrwKWO
smK7e748DyAIQKg+judIkgDBdvgr8EJ/jnsss/ALDKNiky+njMft6NdFB7WjoqtY
gG9klTFbDACHnlESPJqeh12d3knxWIxiobwKOnwaCluuUSktYZ1/FoUCcJd6ziFf
GLBBdYl5xpJfttwS+QKv/vO/uFqSxsi+Dhlr/lc6Iq9o796QxGGfeBwpBzT0AcXh
Sex8fAVLwSNvAWOgquFKPeEM/l2c/Apqs/UJzk2WI+bjNz7TST3d6yRcT4isW3GL
RuDSwBNRPnPDUrk4LjwMPMcEMQX3texk/+crJ1mHm1jn5zArRvmG7etzEp78vAZy
owJteqE5m6sIcxcTDco0CBvjqY/2LcDw3f/23JSlI4djoRxBr3ExE+YFH/cexwHF
QH2+GbK944A3lo2tKzHQhljUsqIIyFVdQv3CB2HQf2X51R2S3SPJRY7WXm4uFRjB
j0WO8Kv09mdsLmqd0A7qOAGgjqRndhf4Wtj3edcHNiTTtAmR1BF4iAvMPkKjftsN
V8wJ2d/Mf9rTMepKYVDlGct3yId6U4GM1vzSbl1w8j/4iIKjG8xpHDEHRAou/1Ne
ticZ0+qF11Kcc1+82BJAZ5Dmk2Mjj6mh8x2FCI2q9zszX9aYQtMZfLds5L1eEsU4
pTDn7OUfwObibdSk7brqqXdcL7ks8b6oz3mgnlRajcVW4MT2ANbOOuXGZy3VnqzB
Ouq4zzqLOVAqVC6VMFFZE9Pg6ug8+ixz/bCGB/LLyGSdCQ+F5IczeL8TzR/rAFlO
wuDXTsZ+/FOkRxkEBssCLhACEHlCIEhJiWmiQXYWa3aP6VczBvunoWXAJHl3O1w3
aJNtifix3sNK+j1bWIcqINe0odSkepk+WuhOPtPGL3V7/nEuK3KOj7FdGK2WNIHC
kM0RGSNzzYQ5whwbJs3OFiBGkWabErKXMrGBt6KFaj7TrLXYl5CMbBvDJnlxnF5a
M7Skj7QojmmEFGNJpEyuEZnnXQ7QmJ/nKNKaPxeh7bXP3IDS1o/CblSlSDJe77AM
TA/2VyY2liJXWXT8QI4yTwRC6MdBc2ovIMAhqAc2HUb6hEiHC5VmdXQ5MoNPQ6ZD
KZbAcjpEGOPSiyacoUqFeNmyyzBtlLY6WV23CFLLkAtbg+VTP0atBqvNI+cX5oIw
u4XDkqp2fYk8eSC176XWeV2ftJ+5bBsi5ec7VA6s63FYHgs02HemVnM5QswEa41i
tff4vPz+bzeXNLxXodKbCZNBrX0iSJ1U/mUf9dcQu6TCb1PIXoqi3g/5guxVf/1b
+TEe9BtVftinSLTvJNLYZUbfYUfSpgC54iiXiwxQi4r0l0HN5iyE4zh/Muo4wEbH
wp/sx3uVw0trrEIKTjt0XoFHC7yUbL2aHbva65WV7kDFJhpJ7ixNtRF7kA4BRS4N
qwL9Uu71qMW4PZvA5Ei10BJKYn/t4N7POQd5fxEY9GChH/rRzPoiEjxfdKdQ9nSd
oqkusRo9upIEi/cZBdQhkIAp1virJnrvIjDtCN/g10ty4uc0ID3WiZ3Eh9kGh+hX
zhQkjgSUCNPh3JOW7yYAxPcksu1qeKfVNp1A9EI6Fxkkq6HaMOWHLdTmhA/VG39w
OBQtEvkSk8OsZ1kUNsyHcWkWh2fo/JBPAE6P6zXEar+EdkeCY+9mfKYA7vwuq/Xi
5e+5vqBT4TtnHvkksp9bfukRRwoalm8veW0KgXPIl2s0fiXXE9JnYcjRgacnZ6QL
RYzuV3xCNMwyp/PhDtHw9GB3RM2csgylK9/9eYnndgY1OEoMe1tGrBi5z8F7AuCI
ml2b8KZ1cGvHKbedSV1gS/rQHhzZdT3ufDLx/A8dP/6S2ZDntJHGGR1jDf2BjSHj
Q85em/GlwBGwPvXrWXjp2MthKBxj0a56stk4Za2WcCQs9BGJW9l4bSKJy7MzreOX
GgDaiI8fpjDD1JVaAbYLFd+0bZ7dKhRCrsdMszwY9OC9EEaKuSMPMVJR1gDmQBit
DNipwWuESCufjmoD0K7bqcNZ+j5Pgkh7MIq+1qogPjQjcVV51cj76abVSk2E5q+J
CQCPstiXhvj+uMKqkpy1Ven9gwhq3AjXgKjiqs+nLKT0pHG75gvnYYOjQWJOdpn9
61s5l73NSQcKXXIfxgV9t511gz0zkQfkqihnW3EsQ5s9nTeJsOXhcexuH3feS7By
jLdilitXsoUG9PBZP1R83rajRlfyRUAZWffCVFDzluBXvLePbP6iPd4j9sWsk0XX
mADfEkyGjYWUV+RLNMPxPG2Sk23CAELCReH62HAil1MfF24hxIR8jRg3ajumrxAD
eQEdLHiaE70gFsiLtUUU+5sN0b03hzJ+4tcLYnPHsc1xBxn2sEN0mNHy8d59gdl4
8e4uIyGICz4clT/MpikEFVGEXOnpUdUeEgCAdpXQXtwgDDBDzlAXV4lpD8qAqUNM
oW9luyBgwQx9ZcaqeTk7Q4e889NI4YcmCpfAA6K/qRhZufL5Uclv03yZ3bIBOmoA
RuU/AW67qQqc2HeFHum0I6PrZjquf8+dQvV0W/04hMvDFJ11qRfOvco1Bxqd9dP3
fHf3v+LERmUb3EQJZv4R5zCe881eVLvB57OJOnbN/HsciwhYFoRu6SX8zEhD0t+p
lA+qED3+lZZzelyI9DIOiYOpZzMuTh7GbntSjgdOB0YCeG4CZTIflXIW+Ql/Y83u
CegXMMCNBkv8ik7b+IrLKeAEUrgs2WVozqB6mErAbO9se8tZ+wbZDmt8HCUWntQ/
Rpig6lhjKp7aW6G/k+YLLePsg/eOv01DhIFdlRTMozlwvAVNRBBPbUkSH9tKUEhN
UxC24JQRlc+h8CpRMSPFmD06dJ9uzZXWIwLqUiJlt5F5bwXB6AFusWwFrEaKfvEf
nqVs+RfOYXuaAryypRb3kxPwZLWT6dB+137/gMuDmUGAjfMx+1RiHt8F+UoPKJ6m
K1QXTSWy3AiscKd3JmOLQB+oLAsYtN2oyOKHvaB1mCwQSnr6RadRMQQKpO9sQ2eF
8No/p2QeBzuBFVq6qNbw87cvR9sAyEbPItAsRYQKL6YuBvfpFzhDKW8wqqPK6M0m
oPTOqvToa6x8As1Yzzm+bFhEeJN+2rqsLQVpTsNrT33/DG2ZzaTC4AHNNqkIGQ+R
c8S0uI55UOcVKtZFMkMKbWGrKG8WIeNqecbEfW3EcfdRuprrDdpAORu+a04vcx7h
1YjlJYIso6i+uvfr9Tk4V9YnXvduUU9Wl/3YaoGXxx4mC7jcY9KuiX+REItj/yJC
IJfDGuMj3RC0cr5pxirLCwzf3q+r4U+V3HFKystGybTHvI6lBCYfo2gE7V4LBsQ+
mDP+v+ZHARbqePFMc60XbyywryvzAn1r/RkzHPP1azh0PKg993HgIfMwwcWAvw5c
1oNmIk9tFkSgmhta9KFNL6G/CxaSNxvjjr+6gSKaf7ZwMiZbMbq9/hZ6fikMUxB3
zxx7a+mqex8/mnBCdM+7fOB4yZIG1yfmPX4fx03gGFGipUOecTpstrAu7lwpN/9L
Lc60gV0NQacwpeX9oThb/WE/Qt7vm8yJ1+McHw7yuMVfph/7ZCNvxKjYrlPKp0i6
Vegol1rfHToL4ChZQiVYvuT27yGsmzzidu4JTlX/zWvD9kcMnlOMrIH5hCMgevJV
2ebHXlUur+TEFWIbZ995ypRD+oPAq8W0xk385yS6DQTw0svMzmrm+nZVDT+uUf7c
Oi+7DoXhO50Bv/5IRNTRDGdo12I826UN9jMCspoHfMb6m5cGNaRKm2Yq2aI9CRHe
uaSuwHm5wXDU7me3EJ4epcIzGCTl43j/i0rrtxuyTvN/L6p2ksBSc0R/9TMGOctu
Y+YqnIQ3qR3QW7J5ABAedBDhaQdTR+6iZr9yQMxtWm+dIAK+uZ5/Gp4i8ZLr/QqR
mpmkqo7L9xiFpBKzuljLSsu1G4bwAimabHwB/XBUqM8UEEW6KCUAbS5DZfvU0Nnu
AifGeUt3CPzVDEywtI1J/jTHDjm4R6h6fMyJ48oOJb2QaFmIt/bW5eNmTqs8uI/a
VrljAOOT3cKY8U9ROPeGH8T+cXVonxobzG4Uk2VPA8EouhUADaiaMiLFu5BRmeIx
jgqYmbFoPToJB9kS5WFUPcX50gs3rkq8q6wP87BORtJ3PJYjagMg0bM8oUffQd91

`pragma protect end_protected
