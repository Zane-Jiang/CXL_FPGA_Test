// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H6sZq3pjKG+KQ0I/BirMvAchlCOCKxbJ1kgA5k8JekzB7nii3/hYd3oAoLKJ
Yeqe9FkCCnarhzgAta/VV07g3ujDT7b+daN71TEYhC2YFfh6AmUY+bR3ddS5
guTPiBbT/cYwitcVbO85Oj/hroLz+kEfSuX4wTLoQj16DUMyR3gSJK8e3n59
OYM1zY6N0atwC8anYrikeJHzh2lS9xRNGooOyriXEPjCmnzx7vAxMre2D31/
Tu+6jIfZ0yFCNOlrct7PyHrL5P4YM0XGbeuWmRY0tteyO2/zpV3tYpzj1JRy
sCO6Ke5uTFGuk+ZenVpSX5sy1B9ae7pJMrxRjUy6Og==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PrtP+fcQfqPeW7HxMVxJ9f6/L0WV9ZXTWjIyFqvn+cR8rYK4eoa/jwQZ0hA7
A7G8+eQiPyYttCPyfG3ny3KOWNEvPfRtQHX1ymfmB4DXlglfw2lP5WynfGWP
YhAbDaWiiTmB6DA0KBlnkDoPt4Qybm/ch4eWPeaQclX3COcH8m4VZTFn76MQ
yk2zP++nOWK4qD5mSTOBtp5+Me3kZTuGGmbxyAJT2Ld7f7xJnkPAHh2A1DRT
0CpuxH6JOLPqonKDgmpwqc6iwa0uPoJHHNWd5x0OTt1Z1pS3TyBDTl2Xve+n
MTjJc1rwUCpc2nIeGtuFjDDNVqQRqXH+0HI1L2ggEg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lirdBFXwWPMk75aZZd1mDbj7wnGsOhlsAzoSTWf5MpJSWIFcGOCvo0we+AMC
BnKGy4WI3bX6kLLBU/Hf9gikvG4D+k2wvNWwWRQluVsfs7yqj7+nNGArwQTe
EVG1M19qUQHmnCCD1a5EcLdRSn03UxkSETOsF95PgEWNXr9Jzxn/beXNyl9a
566ktJJH3T7U3InKKBHfBhOmQpN1oC6MSU2MYcXBObuomadBNtIegTeS7WH4
3yZnI5hreapFpNWs+aHGif31HxThVgLJKBy+JGGMyNdQjF3RYplqVHlf+Ctl
41JL0/kQ0nJ9pPg9TDUTCnaCkejJoK4ufuRc2SMvzw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cAGYqdsOk+oGZOPVtovagHcfi3sCBjFQDSlS9FbcWMsCSPyz9JoYbH4TPxd6
TBM4hzRZIyjZ8aKwc6IJSDBpoc7FjVIafN9INU8OKq3IUJ4eyXrbvI3yM2Zt
spszpnMgrtYLfTuwF8O2AwJn7y4dU8q7iEgd5RDvAUl0NUSNed0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
C/AxXQj9kSP4T0X1/xiTLSlxLSkl6z4EbJuoapl1mNXX8NL7r8JT/6wiUt+b
VUalH3MrbDun9j6O2A9KQPcy3FIozSuTkBQXo4F8946sOnabXx7Wi+vzKKGN
C+WOWn1SIWZRm8Njcmu7zgGHk87d7o4/kppleeWMk6D8ooE95bR/zdpY/K+u
SnzC6u43n7hKMzbVsLRXJGuex/2xTSF8VN3nSk1xM8kjDTmuPexPNdzKb6Wo
Rdt5nIxTJFW9HqXYkQz8e/xSfrdC9AFaEg4kkUSW6cv9dpTIc5QAICLZZpp/
QVwbWl5v4XaXNgP+nXMTGD90cWpW1WNqPea09E8sArLJP5n1WLm+k0YOOkI6
SwrvJFJQTuyKr3c+xpfqVzyX0GZxp+vAYaBjUcglSjg+TuE0YuSSuUmrsble
hVbqeeT5N/z93jQKktUXzYXeFRMuqjJL/IVkcRft8iqltrNIXLzct+YspfA5
DmgsDvCDMsO4dvDA8VwRVpJgGJ00CM2/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NOkqksOfyy2R/5+bZzAH6RdsCVv0hXvb/LSvT/6nS20oM8yhQDnymWqjbmwH
/+i3bK7XtHoepfwtziwZEY7sy/ZaRgArbi7/gHJRR9bXO/HZEKt7atQ+HHVX
3bzl/nM1o097DrulqDPTjyqUXqs9lO6+6mwCgJ6vGSTm+ob4spE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kQIkk8eu4PWHMOFnB94rESGBqFL7qhK6OdzH8psiVuHosh410ZwgjQr5VyYR
Ihpr+r+rI4U6RbAh0pW8kzZKro6FqFaiF/6viKAu1QQA4V7oLDYW/wjnEDaQ
ksbUT5rT7UV1ydxcU5eNPGveux/uOtAG1Krv2KFYFjS4EWN+7tQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 91936)
`pragma protect data_block
fXEMrRvf3mLpS13NTS1H+6MwbuanvXk076dS3CWFNp5usxMg0yvHJ/G2euXj
Ng9UGr9ax06T9QSVQeVf8yznlHEXDWtt8u/PA2RXxxqrBynWL6zrZPwvum8S
Kmi3CoMDUGX1sRZDM2Jmbmay/SWqno3XiIswouwjKbpHmMqfG6jRT02IGzkc
MYL9Mg3+C3yPfCZL39MT63/B5bJ2jD89IzxXKGLhAtaKBnHDS7EVhY+ETlWS
NbIrPerII9yp0B1WpQMXjPwRiPVqWUaI9K4wkHtA85Pp9J24rgl2hZ4QuPiR
WoDLDXg5W07psLhD4i0gSaAe2PM1GZ6qI9ftK34Rxu8chBb7oz0O5krtpTsu
HfGIzjHSUSG7CQUUEvhKIy0RIJpIYpS04JJo8Qc0jkq6hCASBHaEUQ0h1nyP
H9DZpHkKKsDKMIbTeP3q5OWLyENdn+lQjs1bEJy6qhpNovF4C3cnACCLlirV
YvwepiTbN+Qk4SB/DVViVsZzKxFnzL76UIXAbwmOkidZW3K1hE69i/hVJ9wh
KMxBV2I79TpU4JOuxtSU0XiozmbKkR3dF6ePfCtqxPE6XyYhxUiVpvjLxaio
rTWFgYryv3LrTbM1MiPXO74jeNd0Fs/TZ15sOoBBKyV6VeKh95o88b8w/5Z6
LSGqmSwe7bUM65baluwZ02u3MDQkeIJkTb/+4abEgomCiZ+mS54kkM5WRQcv
zUbS2sQ1rc0L56valrgzsZQd8BZcxOJh6xkYV4FulDXrFOqJ0v+LDJ/KLaVH
H2q5X+pF9ad0hcpRPIJasvRD+H2pe78FnhIV+QKbhlmJWbqrrPFizRZ6YUBV
deYjkKtJyt5v80ghs3c5/JdH7s/lbIvr4qO/sEZrAplnwUH9AhOpOak82jcz
bDoQJtqORz5DLUqSP2vhXPAS8nRdjiktV2GYIAKcKwYwegn9umeUNrU/xYX6
c0EFNzT/Y0wgNRjxY/1HJcDp709r3FfBSxFuN/8L6/dXGXfGBPo83a9G6EQD
i9kjls+fo2VHxdShikINr9ktgY1v84Kqk+gyALq53ca81Dz5MPOjbmOMKU6K
pI92Awa5CWs9v9bZyJwj9Sutq1X/b/oh93woAo8RZYyT0DLlXT5/ASXmvodn
NqXknrPHyP1qe877zR2d5g5I2qEAGm/S5lx56SQd36FoD3TyVFAUFrZxxiMN
AAeUVkVrx/YPDgFVFuCDt9hlt7mFPza8SsbaF2GW9fFt8/keQFdVAbeRm8cS
VqMjrfoHlCRzjchzcIPPNbjMzdAnVsHsFnnfWmShwaAYuIexlp/VZPzn2EiK
ZfvHRb07xMXz6qyLA3YUC4K0L9Bx5Btds5ZsYKD0g/7K0LCDS/I49TdwAead
9Exkj8nRJmIYigogtNElNdn1dKGxzmpV+Io9pp2r8FVgOkTVaODWrXtHjdz3
521CX8lYZDHAlsVVdad1AmUIYJ4A+vlWp1pqa+UqXz3trhg7pTny+4mBqr+L
1rdE9S7je6kdHR3tIuWeLhlDKc6bczn6d9vkVL5D/FbzkpUNJg+lNlsETIyI
exRa9JvXIkIYVbcDjNDMG74OVsEUlOX9204QEHsOt0GmeYuZfj2S0/bX7SQh
fCYgT6EEIYrSix1tr9LYXIWH5hYINITzGKCVeGqindFuMjknv3/krdRmUYJU
WdWvoy1GCqXvJ/qYpQVc/AIEqsH0S2JcbgzzwHD3j8X2jmVgkxH7Sfk8u2TV
zU3JTcyQraepif6inQ2naaLkkx9VOKdmXiDS27KQBmBxMdK6HdVvE0QBAlv/
1AC9hUHwNRhqpv+4uwbuieaVgpXcKxD5abQiH1pRx3xTLH1mwXF/HpMUxQU+
DNF5zKQc0adtFdFQ+N35oMOVIryITHGqlssTtYpqjBdPFs9br1SZ3v8w2sdi
erELrq1gcylZp8DdZ2t0euhKIJScZd3StkhTNUOijVEuGGgeRSoMlBgeAe7V
8aUqb95OWpehX8gCKTQj5expiCOnEuHPuEEIwOqpKffbM5gDFwaZu1GoPqWo
ov5Yody0WvCJ6kpgpPfPyvYgkIUFMOrwYYsUf+nGS+Gn+Wb11h5QP4RCV+TT
3zrrpfar7z4T3X/FXGIfrz2Bg6OzgCtMfwsauvMacaqsI2v7Qr5wfszMuiab
/6OXtkPomhBmICWtkzzXmELh3Lq4cvG2roFBKuuVPLfG0xvkJrw3Kf+ReGHJ
Fy8s7VJ81Rs4fcTjDCVTUX0SEtdZO0anDmi0ZDOCkHzKGbWVV4l4gTsFAb3V
yRbbRMaSRluvmT05cWLj2CwH0uBbyEdKtdgi0YO85wcNwRSdh2zBj+5HxNCh
90TbiJT2Mblto+bK7HZz0nhFY2OuYK2GXGHL976azprAFVOb9JX6cbFtycA4
STrvjkDtpwWZMuhh4WIULoqHY7f7GrAEdGXy0C3WKGdRswIIt2i2cP8Njkj8
ChAq2IXBY+UpgiEe6yFUsQbMqJFp+Bt2VbtpSvbyN5+G6822c6xhFZZ73cse
gBXgyjSLU1fo5TsWGfN6iPwDUUzLsBxkt9lBM4WFI6+s2eO0pM0l152DTW0H
oaaN5NuNQ8SmzvlbamZzlw0XR/aP7HT0ukfbzqzxZ7eZuKRac5Fslz74BlJL
XzWiCE93mfOlaeiv988meMk44GxHv1QT+4h/XxutUvwk+l1ylkR5sTeFOAwV
qq0zEDhMsoIrlXEz1vgn58sr5zLaJq8oumy0snDfttpL7PUGCkQKUh/8YhlP
RJDN8msHs2nEnrN9LbayNhuMUrzzYHNHPN/CjVLe/F3kDVieyxHai8EZggGj
g3eb/aKPCWEuIaBdDojOdeu+dDwDpBUXy1gnTC+DI8aojdml5Jcoc6CZQuEg
YEe7XkhGJwLP4jKpJ5/ceXohOVASZlNXSFPYE39Xzc7AKMXS8EsRad0AuLac
3E3YyxZlTGIGdqgzHJeZAmUYW8oGpXUfV2+D7faKglQEf5b9i8Bkttf7Yl1+
UbTu9AhH2j5+d1DSG3efnLBvlGSoatbZgeYsSrDF8R/eXxPwm2waPlbwmsmC
gg43Bm+DihxEspq7CUlqtu8r4KyksPQKLU1KddJgqErgHA4nlBBz4LF6cK1q
B/ynDEDbBliirTjxPnJgmvyYVxwfMBnqO4eVC8UNR4KRItsJsDtm5YtgnHL5
IxqdSjPHxEftvxLqpnndf1dXa2SgCO5QKo18BIa/LC1COpH6AhdrKo3SGqHc
vNbgMPEuHBgKAMWeblCZQrTUP12Yx2xqVgzEMKrx6dki6uIzb5OTnEEWpiSx
ns5Gm1iefbMIMqVGNXOeQS6VH72f6Hq52AJYMf8xoHRipMKAmUfAf1X292O1
nE8f5SKD8/0sVwhL5JmCbNKagm6SBj8Zb6R2vTew7BJ4+TDHh1t9WugEiBc6
ijtcV1EtPBCl1wRfbaAYpQwD9AT9HwxE2hRR9rS/GLpL2I4Jv636bHIymHKg
THizG2/jycWXVV+t63U4x2MFwMiMxCEvAu6LjNyBKx9OqAuVlm/83EarWAYg
k7zOMHvmzBzH2I3NNeOUoAvhMlIziqr+xYfAaiI0WRWIYG5bTpsESK3Kam93
L21MjktSQ95bnqyH2zBy0XiJoSCvzSCeFBwTZ0y69RErPSLCHgC2mCHSlTqj
9epyfY6RqLktzZ/ZyPL8bGKM38yxcMb/pc8NOKMj7X28gN01ZYs3+FFBceju
8qtOG6Bkm5ImfcLP1NiUk5l/PnxTczLENi4ZztgY2GMUcWs7Z4mAmX7qybra
5RJhiIWXihqFTjwW1AiVXpyki8mLPDqAOFM9/jj/upFt/Iiy29VGTqsvLHOL
JA1z6Qx/CEV6PqiHxOuB/GgkWqreXAFS8PErwcRWEmJ/MjZ8hf8vW3YsxT4W
/YUZMBVOTS5G63+mb9V4dxY/ERXRKZLPqznCyEAxtre+4BF27FdExlCTtz7x
nw8Tkf0M28Zk82uQ2PDOZCvh6qfA4Bwn+8oaE0zPJtzc0jnhAUlcO/TIxAfj
fY+RbfHuF8SWSCvlnCUFNNbfM7h5NBbyN9BXdO6cTxqRYSV1PS+3EhXcydiV
ipIcq/HizXtKpbW5c0DJkYEVW8BOixC2ZlZAOLqAwaG+A4wyNkaoxFeQ81Zr
FAQZcP7x8RR/o/Zm6dtaqz18bqkUU4DIGUVLRthJGJtA3sVpj8EeqTAwuhgO
2jqfBL6feoIm+m5GTUEMNEK3D+1pIGnvF25a0bbm8/smyPGBQz1nzqIQko/q
HMt4FEYMCUk7y2xVvCrOFJoNkVGWpeXdtkxkG2gYxgFqz7Sbe0xmTHBT27RE
I18yT40IUns0PaFQRluDut2WEtest1AJ3NfYlSbRbm+VticZ6QY9/CQoJuKK
ygKAs8Dm/zuT1Ca/zNQtUO8rl6nV1Mowwdw2W5ko6O9ulPaT6Tyl41dWnsWt
UiRALQKiYYNghS8wOJLbencISmVBzOSKDkDOdkCSknO9MuToOxyBuWm2+i9C
0wrz6s8EmiqfDXprz2QHRoDK4cXqkIiOx4AuDf/Xf2V6Vyx1hwYmZ1BQSUb/
/NjrOVS6Fi9aUuS9bATIIuZDc13+uwIcQdv1DsjAPsgVj8RXgsTTP1P3Sd6x
XzWwg9yJYS7KRlUEmVavRC7NkUZM0vtS6xo1+l6ED5UiP5tae5Xk87oaNMpJ
faCoN1hz8psgQXBuxME4loquyiiPVA/JL8D69oM7IROgrYkFIn6A+2vTFRew
d0DJUPulxTUiMSstKB/VjcxJ+jpBnSX265b3KCKkk+Z5TY1W/ejDEKBp/feT
SGBUTggv87ruL+XoaMCDyZu4JhZKVW0zqKiu398okNxrvYmpcoSg3Oqm99Om
ZLH1NWKHhpbs9uDKVMIWGMcJTkdpxE71ng7uhXC1/W/NfiKqaxLUDaqRwKmF
ytEXZXV45Dx7gop8TH0I51+N3kq145oxGD254beND0fg58mLQ0A2fEHlSGEc
Rdh+bqyfKirsLweoGatuazRie4AzmZvjd+LpkN8sKqgiaYaCO7x8DsIM/Pwa
Y2ZDVqsJhj3fKNmiLvy8a27Evi1YwD7VMATlvHQQ+ZWvvK+/mqsYF30O6URm
n4OOAkmk65Am4N/SmL/m2LGdzd3uy36TqQHSViRuhNG492ufrVOtNtCNW8YF
Cu2j5C0NIaqPXQ48Xlxpwiodrem+IkPGytBVkyqP58cTYpXyL++T0TrfcWSr
dOVQGgLSrHJeWwhtdH4qyCdYmsXK3i3TXZJsb+bLXW9erGFQC2KC1uskyO0y
/23ooFm5QZbfC8IdcH3YmwYiSuP86AVDv+4mj/OYHG3beQ1NiSA2jJ2ehDLC
Ppit/nbXkKIHmbyUgYWyGD+uoXBTMO62aUlVMTHB4eGoaBFN9cPaAn/sL5zU
kbL0skJZ4+cscYPtXImC5XdP5mWQdH4kzJgQiYf37O9z2Chkf3O6duxTzXKn
gTgIXLEQ0QgfBrNo5kcEZdU5ETNoK4yzcudOLR7HCkTISvivd7ypc+ErFYpy
1uRc62eE9b9POC2Rp1lSb87bWn9NhOD47LgUV9myYxPKCqn45MIV+XgSfcTk
ZDqlkclXNfp7mT/n740dHPe5CB8EZy3zHqfYANwRy12QWR1vYiUNn4M9zZgP
f8zmaQMwH+jZ1Pb+vwg+bd7PkTbVO5NYDEPmvjHFPAkQmDfaLb0dQhQBWlTT
1v2Ey3TzrENLUtS0QMo2acXzHB7LQikdsDDWrXbUdhMeH+GAYryEN3BEPOOr
VwEDumIwp/vf24Xghnf0iJuoHQiKx781t9o5kUHZljbPBxBleDxWVuyt3kZk
k6uhEpO85nJ1byhSihHqjcOdryIt4A0Djmmq26bM/sEd86uIj/lxqOMNbqWa
B0yJnPadPScrNFYV3/ia5SFCbJtC2LysZrSJfp6zus4ZEC3n6dsoAMyoQIs3
d89lH2FRNNriZ+xJnIwAa1gRT4Qz2H6+eC1tN36GTYsF9f6CjvLYAkfCVrX5
PbOU3Rq1qKdTHUxDhJfEHOf/y0X6OYatZ49w9tf/wj0OnBT5SINj6wmMz/Bw
/oyT5TZq2xYYSQBk+f5f0x12GWhpBQBl8hn8lYQ0bbQIX4OJu3cRSJBz+QJ2
8vu5N64Ba/riiZp5rLKpxlUORMxPLwpf2b6A3xAqf/+cWBx4ityKoH7+AZWN
unLE35JeAbW2CQdpegsb7CU+oqXXwvki4HFXwzfDg6AGzPeDCcEbiEeOassB
2o2d1zgIMNNEMRPfuvM6vnzRcZDVQzCD5/nAMUxqvU8ShU1xXIANCG4I9/ru
cC9Jn6K1Si/XIJQLDGsgYrJJAX3YUXz9PbE5Bbih0oGHyi1/xEL2GeoRYomL
RtTpD7NtMv/SSBtqh7xcBGU4YnCYb/EE7f16uMLzXBEVh+0RtWS9jlZ1Vbx3
+vu19dsE5LGKZSGCrwlJNzGJk+BzRxATo8/9KglvVK/aB/jDU5feNl+jZWXQ
gaNMC8rVjUVu9SQJIc0qctdiiepc3nsGeLhXF1oaymHjHoETgJwHsKjhk7cu
6p7pHQp8jpNkYEH+W3QJto8aN20s0JzX6bGDkXZ44b9+hMqen7cIeDEJfUFy
VMcSOY/MjUVldSql6SG7WHpymQ+poy5Y4egD2iP22EpBEdGnVCfTUjKdKFD9
W/HsxVGP568AW67ii6wl8a/n1Z301SzR3vaGBNAWxXJGK9kEGc1ymuShbjji
Ae2H6pmNIONycIq4GxvAglRNB/vRRoGE7//4OIzYvJQ79EtKHbdIkvA8qkGQ
36Bg0+SWb1xQoauO8EfkdQKxLiFbuUh90KI0eoxPtRfESezFz77VSArC9gLv
i4e13ScvX6R1EwSJK9NC3ums8jsE2VKiL2UjyJY1Sv0CnLUyeAlrvCQ4fAjG
GQ3sSFnSneoppxyLxjZeMUzofmWJ3nDjC5i8kyV0ojLyUg3dNTIz5WORZ73t
rTxBReaAuF5b3Cjp5allpY3VTJc1wBHMLdzjWd9pFvgw4T5iO0lQUY6B4paX
jl3sCt3MKt8B3n6Asq2KTkIMAVYUdF26o4O1TWXwazRvS3z9HF68ALxKYkST
GC3H572kvEF40JgsglmQbaOcss4OqIz2NW4QXTeV1PyV+PT7v9zusO0adj5k
zEBpHXmP3OX8FUZnINdZ4VLiGNJ8a4uqavh/bLC8rG2g1X978Xe+yxAo9Fmd
+r+ED0UqzNVylqz1QELR7tQ/G7sK5lauqWdKUiTYvrgvN+sF4AoAb6T2eYM9
Jb7H6lPExw+BZdXtgIiF1789NANrInDT0ldfazeiAE6+hhCDkscLa/peB2Dp
OR43GTBei3/iTJyFyVVa1uNhNzklXDxi83POHT80CUHxSWbr+UxqzLEeROcM
4BurHRaK2FmRBUsMTE976sGHkq4hKPYpLIckBtp6DdmSbtivb3foH+b/c3Xn
+75QTvgMqE1q+w2Sp//kjaPZpZ34qLkaXscLO5PEnimXzBImhaejnRu+r/Vt
lt5n8GDWjCOZp09s4p1mInAJYK9WbWSEPaM8ARmGaT/pUneWrAShnK8YIuHj
8qEIVju3ypbT5Qd+Iknyi8snKt4U9ZSQEICv6YcBugbtWXPXAYYJYusMzf+z
Lq9S/Yesus5mI5A7K307Abq0JZO16isRG12CLYCuscyyE0ahwS+zPKfb7EHR
ZsQUqRHKbq4uTYNXQwL5OYr/FlUCcSbJBmK5UmhRdmNTSRCGjoeMhnXRfFan
XUixOFOBHBfyc7OkklpoyG5Dn7v/iyyKlsfh8xOh2ryB9HSg3kDCcsDSjFaf
uBhDyNUeqA4kkXZSOpn0xrMdk7R317/pRPQUIeNrE4hfjbsc1WnKqbP0t7yd
gua2jFtMgUINEGLgKROsd3k/YFvgXLuygFzIxLacBj1DQpvP0mmXXhZw7E88
Uxa+o6JFNpsBe/l7Qi0K40LvUygZ8iEC1pfyuXGm9Jq6K9krzsur0L6Ae978
/mhRXWCAzoEBxcmLwu4Yana0NGf08bqxGJ/l7S6/oGpEWmauHLpsne1bYgg2
DhM8BbEuAhYFBuNDlnYLtTgpH7+REWiEGnEwzGAkoixBkQ/S+9oK/ChV0wcq
UOfQeFfdjYL6MEigTRlYHv/26U6xCsDOrADuQ8kMOMEbEghrEioBPfRXmcOl
mWJBwRfD8f5kKFFWUOWbLpg7HbdM8deU6x9P8wePlTYOHyQEkmummNhK+wBB
8sSNvlwGNeWhM1hbYfZWMNRioBqJGVpd7+6krLbsNlzDwPqAagUvAltP6qO9
pgJIlmSBmM+3jn/FIYdtgyrOQusR3+ZaMwox8hdfsh37u32SNFUv/u2aZ6Oc
ijtjOX94QBoQe/M/xjh7myAbxUhQNWtcikWZdInairX4wHrCzheSmaqTpvJ2
0h7zLzFHQCHgJ2qJnE0EMMqsWcx46psop6ExpijIsPLoUfVuIyCBnnPMHTK3
f5YtWMCJp+Zb3Q6v2Cqc2AU9qBzomEdRk249YLaZxBfgZOcwesOQJ/MZBHqo
u7bhk+bH4yZzEx8DYL15CWFv0wvryPYbqlgiDLC3URWVo15QEniVTreXAqnU
q4CY6w7o5MCnzlmqd4wsaKy+K3dpSmuMqdvmNEPNzPqRuna8ncaZ8J4YNz4s
mAnGbgFFGI8NWgii7bepc20JWytEssDB1LRk2ukxuu4WWTiLA82Jz9Eg20lI
csaA66z4k7TFT7bqh1O4TB4xguC5C3Tj9gOdMMrgOcFl8r8vMtdBv6XXq0x2
4V5kk1dnY8qumdVNpnHahO5s8wvlsz14GKQZfKohdpJT/8J4BKAXzqfQpxxE
oud54wbD1wHzZyWWWiP07puX/I8aubnRf8fJvwI/+o4cUtNxgMCRWQiTlHyU
jFtnebX6hfVQa/RMgyg1dBfr6/3U5t+195JNsrny2GT3WCSGosueA2mAxouf
QzOrmOue84B/Mx/mfFOCAFz4kUKDLYxAc6R6mpUa9wJrl/tLsjrTuY+BWiUn
kUB51TkLQ5mlWMBh0X+NNDqeAlnoNG3mh2N/qqqP0cHtO4cAYoGVMIvAntoL
ARLe2HbcRZmHqsr83zJ5k7+mvxKvWqNzDtgxcUHxMOdg9ne4RQMB+arZnR7r
pR0Z3981ZBegGy7Sd0GaHtKlmLbl4d9zcx7xhBkTvq9EfAkpZKQirCkl8BtP
4I7xS/h2e9Y9K8k9NEpE2oin1ewTINnbQY8hwBABUHnSKEnaYf6yusoDOl6U
eVO+HQUNsz2zJMaHzEpUvGucGRTOckMOcNGWxWjugc5ZgHVMvGHuFup/A4jI
u56tI3SloN+xfBKmK29HYn+FcaWoa+PlN5G6Rw8nA7hB0FXDRd9+DpoohNxS
3GWc/8vstA+TuC3eATHYwKIYfQ7zZMrVxNTyiP0oWM1TWaovYubiWZ+5eiaL
pTEfwsJfeU4Ne64VBxcHQf7m4rSMCIAEibEFJR7sTU4sef5kRjFw9jX9O5Vt
s1ORfV+baSz/Khf+73mszVdpA2ub0QdQZOeU6UgVjQp3HigLeBXBXyyMDQxa
hZux1zGRexTxxasP3Ierud4m4jrt+/mVXCnvjW7vZvbfCE2wx5zuMRrkrAw2
yNu0QDZDN3W/jcekjp19s9T88+x74cg6XYz6UotHku2Uj4TMZ64CyYyPH/Qr
ujk7Tz8wGFbJhp/My53b5h8RUBYwoHJpZHNdrc2wIZ5N8by/RPl4VKLoX+qn
ih7bKIMuh3sDVIT1oPEwisr5cNNthFOF77OtZqCs7XR5vVIcv0Nst1Kb6peu
et6vzdGzOcEZMBJpN9bayh+UpFmkA5ZPy4NcbUoEn6EIVwfzSlhgY9ajYOqo
T7zM/87aKqa/icRd54YzPnyDSi/LNP5LKQM0XACF24Jc9NPjT3uP47d+tIdu
ir2wgouArqRTGlMvGY7goMhqoCnySCJChI19W5e4vNPYseYt5QNVHqfKhr3D
ECirSMg4/Ql6kGGLDFQuLSNEo0mGtJi2LL9MROq1mDGszDuPX1boxW8LodND
USAa46pMm5yDg+Mm+Bz3g0Mjeh5NNzHdrHauMWxcuzKR1vs00SS9pnFQxTwX
uODwrf0BNVzqez4/w8Ei8EM1jQem0BMM4ZfoYbw2QdKeSly1odP8xLoBHxXY
66+YXwJoSYBENtioy9LIplCm+dbvuUAbMmAa8eiRm844LE0cIpI4aEF6k+Ss
j0zlwLFDw5hgyH+otFXjZx9mkFQFF/XEtg25ZU1kTYiKITcN0pFy5T27U309
kghwOAKZg8MdKvtJRXgioO+ACQfEN1rR7pINkh9tP5FGXrZn+o9lPsxVft53
qpdYzHkg3zyxT9BN+d0z6fxkDJmH8l0j1oMmifiZk/UinNFWrI1HkHOGA6X6
DYV3jmeJnH8saJ1K5IUCjkniKM+tuLLj7jMrEywICLy2mG5uaPiXWJoGH3xo
8Cdl0/83kN0nskEFQXefLzKqTVzPnY8In6cgZeMAGM6Ru3aSmFHJOre/uYwG
eHrr8Mf4EQrcpq10O4rgULKJN8X6QhFlHDsCPJmRxAl7Xqrqxo/dFtnV05yp
EkGRS3kY5X0lyXMsTvA5Sn1xz7cAOTywAGzyt73srP4jCdvMiQ9Hgu8ugYri
aHwRsQiP7akV0aj4pcIHQ13yhBvRrQZKGLOM2SZ0SFWOEwSaxx0kIWz7MEe1
Anj9GE+UY/GYZED77U2eSOTtxekPbCziydEWZn61gPk5MxP2knaje5FZs0Sj
TTpghRBy4Wb00ZrdZg/U0VPi4G+xuCvZwvKi93o5iX6oVd3GoxrVM+bLCL6g
OVbbIS7nSBAR0ZnvnQ6PtOFv9iFloI1i/OjBfK0by3dmEGoFCDLpB0BecdLS
iZh+lP2WBsbR4ZwxdYMhdZgTLPs5/8MIWdnmCeco5OfImyFZdtDAMqAscC0a
1fXp+lfTkszs4Jgb3yvZCRrqf9D/Tpblk66fWogYiAhfYlCh0cqNIE1yUEBi
a1dKWEkRluLm63jXakjjoXN0Dz/lpOF5JdrIpgj2chfKFaRuy2a66/YZrqg1
bX5AYc/YQ2HqG61+azaNX1Kl9SAZihGj6Rvc2HclYI3iEHyErYcog6h/biCJ
iYzFgMBvKLY06ocCNxIKQaAsAbSc0r6GpyyJVC/Z1L+mO+KXFrxddvIP9M8Z
B3ImpEbH2DO3PiCGoJqUKMQPgnZLHql3W35hNmJ/pLFqe5N8Kpd2cttxo56Z
A9BqmNo3XT5AIw2yR/oycz4myXancIwMUd/2TGGUaSuJpu3K/IvqpxwjLa4z
AB1Yr2GpEQlRSsNBBRC5/O8OvN1heFBTP6VIpTrWxS9vrMBMBZ9iw2y0ycVv
l+VSi05GeEaIVNQW29gn42NkuR78yJGGwnCFFnLhWZWKH7oOdIVa+vCwwWvI
KY0HBM1vbSVvLB+8mPabqjuJBbPokCOkOqOT/whRrZ/sfxYkuIvxUyXRBnC7
ZFoTN9PFw2RKLBvMbWaWnhk1fI5zME9NY3xUnNyw+ovbk1PST6xfIYrS4b6O
5plW90atqU2MXPcZQfwU7A6oWkrhBOqZqWm3Hz7FVNDE8caNXUngdXyN9rT/
T8ShtnpNkzVxXsHHIWyvfm4zBmR1wLd1xt/7/7mkIPVlwOzZ3gQHHNwAvW/B
C2MFNA3r9tnF1xTWuQ/Ag1LcoE53CiAkI9NjPyLYoMq+A2T+r6JlrmGFpcTE
4t8Cgg14psn2rgnS9wTZDmpB7aLKa17cw35hvMOIGYWX1QxeYkUHK/Z/hrkM
HbLdQoj/DsA3npuiIlrzDdSorRZAdWq9zpBKDxulBD79h7sIpPGiu6ztl82k
IuZoCnoLzN60tBYLEiH4cS3aXztOnnDjfetus8H4+7Eu9p6urrnnU51JeGsz
5LFExW3Qe1cDVRu06RJMglF43qXCiy0C7MmMfHoWKQOyGNurIfNzPIe6xztA
dH2S4cL+/oG7rxc1WjyLoQAAdqLV0inzuJAfT/nfFZ0U6zZcRBYzp74Owzcj
Q7/EEQbfM5fB22F4u2EUoYEeQSGZzTfLo+k0vnHs/bANfYl6S6TIlAdntuIj
wyyyvq04MtjV3y3ZihuMQGByAztNGjaxN0vv1gVh+u5YD0eWmQAq5+hZEnIw
cRth32CV/2Ecwd6T7j5RoWdBbKFQKH39j8bSlMrNVYex7GhMccCicruJ2WCY
R8FS606Phquk+tNhnkEcb99BwuaFgFlCOg/Xd3+2VK+SMere9dRBBOj/jxX1
IJ6IT8s3qpYqoJfU98qVPyVoa60KPNYpgl/j7JWY2168oUDcwxRv77nqEn87
2K9jjU7kYsWTuVIOldH6ratT3qx2rfXClReYKCwQanX4PH4F0VpaDlNdm7yF
YimURXNg6WrE+k87UiN9rD2T4JE/K/bWMYnVqPe2SDApGLcdPqtlGShLpvTH
DpUUYn3JpnTX4ExrwRjRa9bDYywa9Sxwx7yTAwMGT0geKzHllhaI8jtTgjab
ZA+XEm6gFQyi0JIN77oM6AtN2mbyG4uwixobr5w18xuFFd8g1Hyu6bLhvnn4
S/AYsC9Olhd+dvvPtppzOe0NGB3Sdf14ah8C4rmpJ72PQA1bXBj0NU/jxw6+
j49w8nalDgVHH+5JNjSfIj+PVRNxrAdoWaKeDCXsAiTJz/OkbrfFUoR4QXHQ
asLVAO4UPxSZlw7lkKlEE7sxNdFBoQYNyT1k1NrUs/vk0D8RcVmCCiQwYhyy
Y2eokm3bs1OInt82Jo+EZ2S7zYfIIpQeCnGboj2EZGjc6EnUCqLfz3oouzNj
/hZ9aXRUwJ6i+tcn4+yrDbrYJznMszKRbXoR5v0pyXvjyR3Du1xor68tQqJA
YYzbhalh/Nj/A1tOgQXmF3anu1oOXjf8Mj3VRGsYvMCyLZn2116XLSyjHDie
anW1Y7LKtGJXcUDHxvRkN74KA0gWKwh73gG446cjvnTn+ObkP5q78PFUvip9
YPh8lZ53AEezHF2YPO+O8dItQCM26brHpfNQgCkyDuk+X1tIQ88+y1NUKdWg
6AoRYBdAIFrmLotlydij2XNo4QSwGB7ok2ZsT5oLrzBzGTA22aKM9l9SuU4d
bf91pJiNjdT5kUbsggQzm04xm7dIeRVzG7eFup75JOC0Q3EK85lfBPmHG7d/
DMeNbo6IDfBrctMD176yTuIDawnUxAGry/FA1OdDloxODfMXXS7/9WQCmh+E
NWOVsuCToSPNDZtF8qQzSznN7UND6/c/mUMIFv5mKr5WwfHunZd/3Q1oK25P
5HCCLmQkxrnJAtgwiuWTMmvAGnnmu60dXwnJXyZW2aXv3EGbxIMrriDtHC+k
gFt5/MjTXpHKw9OJchE5tb0+RcDwRG4LJsWyHuhVPoNK1lOIM6JosrwB6Pia
vPwUHMOerhtNFhbA44+Gq9wx9srQOiHkZdOpzHBmmUgUDt1WdbQFyoSe6kug
k6PnaTXs4eeSSq53AopR4ST3COlsKcxp2b+ukM8IRUrqhh1Fa52QZ6ulbKlr
8LfX4ymkl/IPMFHe6mvU3Bx4iq5KOBR0BbdKLpJD6nogeSWz9IkChGb9fk1a
/Ud4eHXuP/7CSeTLWl1MOQb88FVE18XuVfDQ5wblBt+0BeSrdj1TOdgkAwf/
GnhMZo6bkqMjMAGe2Vt1nCw9nfE58mTGpU4+g7hrPewx+shIdzFmheFeWcoz
mYxO7WmCXgfYmlibCWG39jolyiKoJiy9UDeXu67VK3c0eVQ8cV9qCjYeYhmc
Z6hlJxd5uVkgZmdY1Pv7fH38yD/msJgM43Eg8AOR1Ldq6ETxZZjYcVzppPRN
/UudWXI6Vxxs4KzFsCBi+FzIWg2X0lHuSrWE3drge1+ZO6f2o6UxjhMqb8ex
/iu9vFjt6s8to7IkVM+IH9RH/e6KvlfM31yEmmsW3NdGtoqnJwa+bu3PArCC
U/l1yEzwu3MHFz380ElGtLhPPZibJKNHcCj3EPDUIjU8r1XiWqDLxvWo+ilT
OQn4vyOq+eXLf0RZGd5qZrcOmQjiNWq2VZ3yKObebILUnzf0OWI1ljuJW8YW
Z58Phcya9wUnLtymyzUeXVp8/csxCNlxkF4pB4WCxtpPpxm4BEcSeke7dMhD
pkayb4EJRGgwuhgGes8vUKrBzofVxtdi3pL1sQc1mXF+mVeCXTxXWV1T2VBB
IjPX7N0oVHYkyttgxsH12Ch4zeWCavVHaKd/VQfGNw/LcBeGVGK7y7gJVAGs
QW17qSoeQ0ZBmcZkOqdf3B+wcKEmShglxASc347L3ffkgSJXdyllaBSkAf1P
vyxJjgdZ3dObGcaiQHr2aGNMw8EpVvNBhN2fDcWGnL8eFKgupbe2Cz3120zf
63fSI5amG0dPVhwitpLqF9SjxZY5cYxlhgyZ9jzRPtDcgbi/QhMA4QFHr08z
958Eq+3TOvKZj30kgTiBajKlPiIgCyATdZjymL3BWZ6kbtAjq8kl/+tFxXTE
mlUA1lt+KSu1Ju9IGiDYMnfSBYmuCXAC+fonu1PAp19lPxqijb7/5WBDUK/7
MtUGQDt4+fNUUKrUgwXYW5S1LzB0BEZ5QbYNqyYEKzXOvRO/daCWcX0zwYD9
RDhBh7FfZzHD91UdvfEBJzrQnkbHpcgr0pwSR51xcXrlCMoomqtsKwvwjpxz
6OK+zGRMUAQX4UFGo9xUs8NBmGGc0NTHRg9ECa0Uk8BpDUOveTYnS/BCuOnw
xcDFZduK3mDH2nbRyK/DdsHTkyV+BE3SxWENfQcUYICZwT0iTjth7UxGhPpm
LL6Q62KOOkeGw8d9BSdr9miJ5xdLVZlN0EMuZTvFydGfVVEw7B1BaF9Ddjx/
wtzpfbL2/kzZEpsU6uKPe/7VZUw1jju+kDsOSp4GT+yl4iJXIv52uRavWcVx
FsBbjsNQXeCF/4Sbm0IaC0eiU39FH/EGMZsbgO9oWpoxerAN6vRwEltFG0Yj
mGbI27q9jklgamkesyo2lqgyQYX3uYeB+UUpjubO3JfJHTR+e8KcGhOG91V9
pFxTzZkMU6783PlIHlYnb0URUrOl7rn8G1/vTn7JGdVkkB4DyyRRvI5b4WOz
BiP+X//QtaxSPeR0fUjhBJ7y+1PFf+Xd8M5RP5QuMUbw5mKtR6BT8qWfzfIG
Be1MM6+DmgoFTaIMD+dQrZ6i5w1L6p7Ss4LrZWHdPcOC/yXeLAqh/HNoYMGh
B7iL8346YSMiAhGfpvmZFPvAHnst+02sUCc2jSUCHHqnaO2xsqd7JgtJW+Fv
LcL7SEB1WzwhR+8k2XC3a5S4Vk2urfLgpwQRUrifsu4VSVPf6lq9DmvCJT13
An6bgOw1NaLq3ILuBQKgZryrpz5AqK7T+Ho0Rj9M6yFIThl7kcQJUZ9xRfvm
+OQ9LnDcwYPAXrP0KdDpY5285gt7UKw92cMwdQwtqv4PwtyOPnmbPuNnfbtt
CRM3HIvDFjswr0x8YUy/B2fsuWj2g0khOgxXVfynlI16uCj4KJZ80oaFq+uO
4nyI4QTzEcwOEyTtB8tEe49Nky5o8/sxLV+F1qyIRpvdDkqPlRhx5LiPGfpk
+4KeNQtQRqoaxsP/O4yAfH26dEn11jUJ1cKU9vaCzzW/NpeP+B0zGQgSUAfu
RqV8qhZaK6ad93AB82oInRPpdNQkjPH/64t1QXF/BVAj8+i+C/3nvH101wMk
bkf0DpdPGaf8pk4aFuygI3qBr3CrVt4Y6qSv0KfkDT1UEi7xIMWEEVtZSXD5
3jIw9abAv1Mf11lER9UW8n9lE8Lpyt5xRPvbnROBTV+KhZHLcbzGHwnprmlt
rgQhOaQyfAwOv+T6x3FI7qNJuifj6Sd+FPtwrzdWeNs2dR9LtjxDgTODMyqm
bV0UmMMZojviqjn7qI1XSyQdtMsonsio7toSO2GneSmXg1KWktmYhuRDLqWf
upfB2pp6t0DtNxY6KnRcB0Amtgrovzr4seAlJKjjz2ThZCI4bmduxwjUTR2Y
l5XwMqr+X6GgSkA7WhCqclXELKXhmjnK/Pv2kBICwDv/dOI9q8Ikod2u4NUW
WVYkDDD6xnItKPagVcrLyleQDYKUGIIG9TExgghqn5+pIqfMneb87pks23nN
82PuOyAAb3CC/U5KVYa1/x6/6VYZjfloi0Rfz0OqPQTY+Rg9Fa4leezN7vAE
cyYQzLy2m+gEqD7iQDbuDNSYCyVfwSwnzOFJ2osu7m7/1EgS0qsPMYFDPkX+
Sw0ABWH7k02xp5ZzQy4w3ji+A1VtLvdA81VCAn3FjDtEcgXNqyCBN/BPGhg6
Wkhj5oIOKJtzJJfvrIyx5eTvj988IDkDSCsqjPKi7fc0qbl8JJSX5Uv5mrQr
clrkgxHhRl+G93qowo1v2anV1YklSWDuyck8hj986cFRu7/yJxJBhajpc1+6
fkJdxwqoG37nxvniMWskA8jpp2KVBKSN//R6lkduwOM9sp2QaDnskkYQqmRu
oft99prAQCzLv9kBrBRc3k/msGNU0PRhoVG8AQqxXUBVLLIGPbfM804dN18f
9No3/ID/yGF4Fc5M+q/1AoBD6EhjhoMnvVTmbNPwzhhW6Y9IGWAqsglxG3vZ
9LtMeaQCwBd2F9quALh9wDx9dZOg39GYgKb/kvNE83J825radZPVRWWJLmNk
wVh5X8nvBsSgDvFtBnkUiBIcatscj7y9qOD19CZvFx1xTPpBPHKqr1ff9m8K
IgqMe1YWsOgFb8O1q4pGnBA0m3xSb0sHYymBTk6txG1h5fUFc0Rb9xuUTy3C
AWlVg+sThYrmSgBBd5Z03ifNO4dPAzvEpIddN8tjmR4CMv/sDht1jeaz9hCP
zNefCeWkGwCuNHvXPD2n9V0DegxcKMcTnu7RXmV78AdSGlU0pZlhnLXS13nu
tBlhr6DUa+/pZxJm1UMq4oA7zwzCKmfQw4S2gsGUP0OwmzuKrHkphd1OZh9Z
rmTN3usOym1q1ZrzbdQebuZG/VvDC4OrtrQvIGHubD/3iPCTkLEy/vC0acR/
JKzK3OuUMIRkn+AiM0HZ0EgZdtFsRgyRwQ5waSAoPuegt/H/Y5LZJU6YhQ+S
yfXB3pF2C2vlhuX+XD1hD36NQezxeNCXiwmZJ2kLDOZCKIuGwoih7FnENL1C
2CpN8YgRs0lyo1P83auHEPgAgsbEz1xb3XI1BPpuTVJLNGQKlRGpkoYwWvcm
rmScAdfNYYYDRV9yyVGAN0gvxCY79/c2DMnFx9PWUNEeFrRwA49V4ztzRTcH
rTxFfXMiohqIkcgJpOGaiy1OaCQ45kD4hQl7IXASfyxyGS8XHu4dYeu6/YI4
ZA34DyBSHqlw9w9eoN3acD+fKwXJJ1t9M1ubBscbSergEEX6O6ua59lO1CiA
gxrHRiCqNM81+kxcn53sMq0x4ZCfT8osVk5hkAjW6OeCOEaJHBrukyK84BXp
6kT9KocHIwV9XIVp9X7P7URLcTr+pj0bFAbWQlexWiy+g0Z3IiZZcbLRzbXs
Kx6nO9CzMju+3TRWOvbJaQOAvX0p5/2kFtljyT4/QJOsWosCiybaoAJRKLmB
xcDKBhKyg7fBlkMjTLUWFbGA4QDoGvZKHvrkkjLXB0R+JmgWsveEsHJ1DTbb
mVNwcwUbYzIG0ukqJiFIP1V2K4wD8BYVR/PSXUKjyIc/j+mbavtfs2xqt795
CJHeb126uI2ziUSXsBE3LFk2iaUKfbT5jEWHzG6ThItavMnAHi/VeojKNdU7
dW+qPPdp6KlvVwd7n6Ud+MLs2IQKwml6yJ76SaDFbkdkmCGbgJ+2XLUlkNCg
25zkiSfFwoNDXViPXECb4CCCQZJfx192Gib662eJI2HREZSv/BRhPEnJkGZI
6iLZ87INq8iK5yVpbCGy9yNT2AkZuewu3ZJFVO0Q8ZHHbd5QLx4JS2vhGt8H
fWHQIw+QVPRkRU1GK/vHa26FbQuzIB2SefA50QdboxwpR+0aU8OziHg7PkLc
bTuDiyX1k772V/I/3JOSkB7sMgyChNVwnQ0Wbvu6z7++yCNn2chQlo4JfSiG
K8vf+1kTRFbyNy+J23QcOJo1vmsQvFEfafu1+Okf/wQbvFW+aPlIQIkd89qR
D9EG254JT/op7ZULdoREqb1iYrBYayo4U+Fb1cmvezqPtAFIv3/bMp1WruCl
VbKBBrO/TOfQHEu3NUG54HVeMo2HlVlrRcdOSzzMCCioy2P7lXbdVB0JyPU3
hqzldGMYR2vpoBve7kvIkn7LpBKtR7iL4DQ6Mch0FsOccTfUa2wxysk6FEmI
mw8r9OwS39H2A9cRX+beKeBpCZbqVrUmT7yxGLOqnrYY03+eY5J9HoAblEuN
FXSdgvUQBSEnr7kMZHZQ6pOuidH9I04tWmQLAfnznhvS4VxvtYDnO9loUPrF
FcAQTbmpO4G4WB+bdukXjkAiaAzO8ZAb9nBut4guH4rsYBwXctArYnabWtNX
EObbA8u9B+KhEZ9mFXBz+DEPYclAIpnvO5OGvikdu5ir0Y/7tDynKDvJqG8t
nJZtjGPmMHI1b6oOPSsZqx7u3nRD2iNwS47xMS9AU7PpvLMkgTHc/0W6T5tu
aD0Wi1VKXmHWlNwwJxreyoosPFOB92YdMIpK4ElE8w71XfeXgOIkoEOexySH
sH6+13iMTLzGYZzSNllO0Hpj+aCVJfQEOc7hTGYrpBPHNDDpUFcL8/xkgZOV
NLon9UB+ekV5uDaExUM5eT0fT02SWiVtcxwn/nr0qixddKePSI2HI0E4kSbv
7iblLmkqEmDnBt86cZpZlx1Ia7gxeaT5DUEtrrA6ykRAYfFvL+vLwK1KEDee
5mYmVFnHtGNiE50fWNKDjnq8+9HRG3Tzy07HKB9y6U3VJiU6sPkISqJOB1Oa
bPW+UelhGj5IDhiTQXndrFh7wvl32zvDABKTX5CR1kQlXTbh5g04AGBCvsvf
jT5V27NY3piiUIOYzf6omD8qfUHgb07Pf17/sxquGvieqqAm1UuVhE3glohf
THs4HxpP5B3RIeKNc4SxD2e2DVb5/j7Xb/mlZvryYRuf+1SHXRHSmckO0rnK
dS2MKMSHYb9ob+jwOsIsv3/K4gUc5C4l0mr3DQRC1tCYoKJSnIA8u5gI4GZ8
5HnpD4XeAbV/M/SiA208VKY3omfqLW2LMLlfGArUVqD58FsAYCKrweuYMvbe
6NNydZUU5ltLeg0+9i9nVXd2aCm9COUwTKlxfGZQ7sXYzUmwNtdkRFkwV4om
fVAxjnAngmD+quDbPuIuiHd6Oqg5cAoWpLaZp7kLohMg0cTiG1AQwZ5ELYc5
kotUyltQ4+F546nxWumHQ7WEmwE/fMYuL2ibML0ePtciFmTfWhry1h0jiy6O
N+nvr6ECUSw5BEQ9ssuNgINjhJ+DNHfcfw+nLTwhkDfXntPl//8klovq0Mny
6hCthyipJMvv1+9YZzba4TO45AwSJD2VwWsUZjQ4Y5Tf5eH2/pR/wnxuvU+p
b8cd5VWNF++CHqdV5dwbo+wsJMZlMueDuctofdWdNY9uk0sYTVLCcFe4+Hp1
x8O1ka9i3RsFMGnYsk6hmUHnDBzPKDMcXAWh0J3q0IJjYc4zSogRh3eNx2s8
2yK97lI1jO9wfmLgJew5S5bfgtv4OWi6vHopcpKYwmhKZGdCsYTTrGhWhBoW
Oa7uKLV6aYQ1uSJbge4nHEsVjnTor0OBG4jTPe2zcHWBh9+UJaTB4vXRe9jf
rWK70UVbPhAauziGB3TmyGkBDZyMqN3ErA1ykIol2RHmiLZUQR4g/ZP6f61M
9gtfBbRXW/Og9+1l6rKw5W8GF0RaTSG0xvjY2TX5czsq4nczPBA+YYyNqi20
CJC6udIKvJvh63qNF3SrJH5mO3BZVhTPnRv/UCSEuS/p8LSeiLhvHu3+A+i7
cAiuzCWiWl2G9aI0mRMZvePqvSYrNFskRaAWHneU82Q6k1fEpnA0MJ7dM9Oz
/j2hz2RQWBdiz7WlU0RxkqW3FFfKkaxTwZMzM1Ql4dGl4WpQVwO3Tz77OrYr
FuyPbPznlJvfzEanMTJMP9xW6egNxQf5j1TZjlE0W2kipby1YbpJPAt/syA1
0zzywooZt0nB8gWbVbRgu9i6AdO3WShcWTRAxPOl6bLR+dabse2pyOCJrX3u
gT3Wf2Qkbp134c2zPPXriowMBrXCxWFNtevG1RdoSBfb3+dod4OVDTRiH8+K
wLlaS4lxzj6zh9fFk3cTAm/wDCLC4DcaQIYv6gRF47HwMNHMe2pMow9ZGcM9
ugil7/yuQZT7+LC/WDhrkswe+nzePpMvdEZ+OnF4MsPX8XWByHuJS+8/mj2h
XkJ4N1+mhnlYc1Fa+PtpRyDtSmNjmE5D4jHrmkC3vOu7zgkkjWLVkg+ES2X7
wjB4HpQvqVrO3YZVt7WPw42Qpa70cYVnP/O5z3l8wEIvVaPOASgZUN1k58qu
6HEnxNXnBXKqNebgbj5bhL4yDy77CRAWLPqbHkQJhVMKGZqwukVmJvNYrppZ
OGEFWbRW+mih15Jw50xiynfVOBRXkI8n/W1QxsSIwClxQyyWOLgfGmWz/jgR
nq0i4Pvzbxz9IM6lYMLA8OdUFGvPHE/SQLcMugUx92w9L9EvpC/833MVe7SI
zlpnekiGaORrYhSkfFRRzpPYstmRCKm3HvHS/p8SZ3ZaANbFa0YapAD5dnAD
iGppF+TQrcBdsOuLcytiP8uj7v3wrThg7tLb8zswdVohT6MWL6bhrK2IiNn5
QaUFHWotX+DTP1ki242vKAwPJNSLXs/ydAXeorwODzAylMLGoR/gULeHnjzB
1lwJSXgNBwNJK9A/55WU09HV3/AjBieITMMV1TzjKRYZ18rOYYEcrLnrvupq
kf6KEiCMDcuCIIR3Lpbpxxw9eTalnWWhTsxkqMlvgVIXYLdqH4WndT7V8+Td
42DoMbj13LdW3hCW/TSOcoX/mztJROQ1Aa6lCgtAK4OaT64RcRX2wSY0NTWl
5AQ3cYPTNxQseTTnKYlFRDo5P7+euEtrbV+9RXhzoTLy6AIn8SY5T//uH4Sb
fCKvyOj/BHGvzHWVsj6LdEPoP4+EnfT1jslHyTt8RalNYW6ZfczYD5AFq14f
1oYQzJFMNxbczSIkI9cS7KFJ3jNDVC5YeYYttiv6u/gJ8CXmGgNZBNlqef6C
1eU7Lgx5YzaGj+5Eb6l0DulQhYzIbmShVb2XAUwy6rqUwQXslVrMbEZpHieN
V59FHH7wZwBqkwG7tULxK6YhcxgXl/Ar8i5xBh6q2LwpINgidcUHH/L0Pwy5
N6pgE1wDanCF8oq+cdlVcwnRlQ946LnclHjiUc7r0WFTk7ml2Ifs4GIDrWOD
zgLK9c+ulCD9bnWvCQ2tG8Neyb+2d7L4/Vv05sMKQxUfkkoruDqZnkEqOHYR
Lb+iFkYhpj++vVqwsYBkbXc/DoFQCB1NByVPoUPKNj5rxk9l6u3xCE2Eil+9
d4HyPzQFIt3Hr2VKVvdeSgdC0E/m9dV10ra7eK7rKcCuJ6ctiMXLJd9D7Hdt
0vfihEuVVxRkTGXFFF320i1J+EUahV7DnP2Q/6JR3d24Ux416bJisZC+IQkU
rpkFRZqlfrBO4fFJ2AR1OduS6qtf0L5Vr8JA9ARujCRdDfNJXGW7LBFHboJ0
alPcfwxZiKFYuzkQ3Q74nP/5T+cYUwS8oxRIVh8lgDiSykMXd3JErv9UhBrZ
g8lc8iWV9z0DRmcDNaV/qVhM86O2kryg3gBGvJcjRUrWtswD4ha1fBvDDNzK
q7uRrUP9f+S8nDWg3q8zELOCE3TMcczh/0lV7v5gqerd5F2uWFeBK9lPNMw1
yZZdjBdk3KUJYvjk6HEiuC6HldRCJwJMdRCVJvySdnoJ3p/SQ4UNvYjse+bT
6DuwzOAQK9pvvqh6GCS+ago1HNYoBdzcE1fC8noiddnLnEi5Jk2vllbrhRF0
y2LFfP6AUqi1b/4XoQ4TOLs6eMa8DsS2H5fW5C8g5RZiiEq0QEonMOSzqbW8
Cd8k8lA2Wfo/aNMsD5nHON74GY2KBvzcYPRKXzZBrWMqX4giGT6ERhxq9h8J
Jk40xKRwmItRSAhICRSup2MpLQi4h5YjuB092wzMhNjYIckt5iz3txMSmefE
MMMS7F6IMbyr4P7V1oEXGgfv96cifaEZKL+R5yLBMX4UgTxejOAPFwUdEesq
NkHn8ag4U7NK7oKLdb7OAMNP4BBhj8Uv1+gWKg2IEfVS0EM3vBZcWr8Ca0sW
I/L1PzWYNyoSRdLTILiZkXybmRG3CAFR20kfqcw5Np2zDoyo/lYCBlCvpsNf
KWXuMkfiJpuOmopZsO3Yi+/YAnY6LAozr1onKLhjUx3lJkbgHi+JxhQ6S+oN
z0EHflVoOS5ZQtEXRglf2FPb32gEXKwPOjm/mUTi7WgRXzCA0Pcq/peEv5qV
wyp9bdiNL6ud+ufVkOfBISb7b1QvfY2IrwwefXOvT8nEoyJmpxCFy2bb7St3
GNmGtH35iFd14vC6Z8FvM1MaD0nm0R3RI5RRWUCDzJeDIXVbB5s9tCtva0vx
lhfD+T0WuGaqoYstlUHoTWaVW6xdG86OTcVnEPZekqg7bwlnc+r9tN4nwkCR
vZ3mg4/bYNzcu4I78/rriG6D7SRTCi4DPcANjPuvB3iTee+Tqpb1s9N9Mmr4
oyBJAZV7beSf9PjOQS4gJYQ2QGOyeJKORBZoIPSnkO/CEN3WRTZOwPq5cQjN
cDGroFXgSZukfNmq7COAyOSzKJ9hlXq6i/loOjSYjUTOqv+ebrDHvVFz30DB
foN46jNDdxJcJ24fVzCsYEafYf1FNhO7NGhiPcIMfUwbfhG37sTXNUpz6dZz
rcRz8bEEtfp6CxJaDPRWrfMS/49BUKWDk7LXFEHGgNJr45mshdnmaNl0ov77
ATfmmOxSZeuMjUhwH+h01VOMuSY9DBQoOkgrNx9Op5UmK0hI0T+uZiEmFqIP
HPOzqfgA1kWEyIjX3iehoYhKkTfVJ9cxFnZ4NuLLqztwPeF2FNkcxzZLlWYv
YwpDKmb3vGXntYGpmMJ4BpFrbWf/o2hNpKfllfS9+QPTMePaqDGAb6QwJscQ
BuCDvIZvx9DSk8CvV+D81Dq/+MzEEKNZl2FaxqO3hlBeRPRbPtqZbofmMvBX
LRrKDZAyp554OBebO4tVzHqxZaqvAaohnjYJAlYS2tYF3+o2Mg1JKdvZuvvY
Iqa4Hw0nrjCVPCieESYTCHdkI2YyL07EM7G4WN6jdXGYRvd9KNu8q0Oh1JV8
+qsRYALMgQJhjCKr2HyEkEYwsTGdIgT/IYNlyF0tmzbVdh3mLF7T5VWeWeDI
Yk+jtkkHKJ+9w5C5czC2VyRTRwkpbPzLJpUWYyapO90gyxKkg8R+ccQU4W95
DDoTt+PUesqPoDaqSKmVZew3c2h6uZWYyyd0tNtWQDnjtfx3mwmcEDW+p0wW
v1DMkJLS5JnoulN1BBnqpe0C3tE9RF2LIpB+gJbIGAzWhH2ST4T7RDyZ8TPh
FHEuHuWX5jmxxpK3o9/f1A67nD3irWph785+YKMmVC7deXp0K0hTqJSy0QLR
cdNFMrLh0eiePBrTU+lPLZaMd8DbRzD3L3rKDQbZZ8lceTKQ8gMF1cN/V8Ho
schehU9R+N9lBtdsWcbPdQYG5MqfQ+41FhgTYZScHYvODuImiUicMBNVtgnC
RoBsKAiL4D5UAAArhe8+K23B24nw2vf+XceOpzxFO5eFwCp4a2ACzbnFcNYb
HYwd0sxyeMYjzbzl8FbV3QxDxaMvVeJjg6aauGjaEWsdWFypcbejbfoAUhQR
a9/4nuZtcJY51bOeRn9RkdcyiclQXsltFWD3+lu8Geta21owwijnhrqvGCah
46jJP5+eqiOaJzNRXFs9ChFWdtvZpkEYv3lXVLcX167DD4trblD+UIWwFP4R
6oLH9EimV8yi3xJdI3mlQ8/PihisBlvTX1cMXR5q5zzd3UiBOJpmZFG7ZGTy
TS+61+X5f/zVGv/DlSi+EsdfIJERk7RW199KZCLyEI1PdAWrQh0n6jVYGycB
Z2aIDzmSY7bSgvZBUxzqnFFSdMvlXzMxbCdCwZR/38maOBWOjy+u4B/HFqct
CzLcX4gyT1j/wZRZE2HEtOcvXQNNUzfx687F0O5moBCmMUko5t4JVaIY955f
4y7A3stLqJMUvv7iV1G29y6vX9b6BwxXUEODzxyA7qwPwOuRFHda9VBi0I7V
PACFlEjWQeWF6e8xB6pFCsL297PZHWoW/tmpt7BuA62F7oUnx8VpDkbm4Jmw
QzLHZ1fjnund2yVHoxbUp5M8erqzLo85JgiyoBC1YCSPGYSABveoVNy/nmHg
4aQc/kOAzWEbUb9VyBgK8CGn84qHT3JtuQk2KKV1grpfmd0sgrr6hpn6st8F
sr8Cme/vVx0En07PKYkTQfHGepeM3cPb22ErpFIostvX6sndl36b3R77MdL0
ltnafktcInow2/YTGxyRWYs+MddpQTcgHPww/jE61KBe507DJXC7AY3G5qH0
rSQaSLbneX7T6RG60KjdZ0hep4HNNd7RnHfm+Ju6pfjs3pqAPoQncel28o6q
ca1eD+OokhjjvBiL32yLXhyKfJ8g+b+fUNgT91sRbdPYnlwKnMeeKxojmcm/
oQWu02v/tjArRbm6zkUmNy2hKAbCWlx3E/GtWw2c19fjLp1/jMYCnM0SCL+L
QLlgNBmzOtMlu9QxQKwfBWPpqIeQigarZLpnEpjs8ppDIMxRcqXyMnnZbUBx
6H2gvaxGebseRwyuEfsFF4eSxY1XNlmBvvGnrfLnDNorKbLKF40czjxpsxB5
kx7fnZc781FY2Zw1y8hngIpcdpE5FAtsPqOWMXjlB9GHT53SymrLYBMTJ+UP
+foi0p43I+stQuj8zmpx1q1XpJDqDxBAB4tqYWNyE93e9zHFRyzAVh0NWDBF
UlZ7IkAxn7ciq/4/Fm6Wx6UbEIu5w3f+5zHzQ8b9sCV3lHuRwMeBXS4mx6lk
XLFkmwwlRMU+M2QfPlP7Vgg3V1o7Q/kNnc5p6vcJETA1g0xMpoP5q4af9s0N
EgR07IaGcFVqu/amsUjQsK22SWRpxnG0cDqydAuZEPuXAFMpKr3hCR/HnHdF
uE/f0SL1Q4k3asAKkLHz7zLgEe3w1VB7S+uECM0kgnNqXyGjLGN/icsid6bR
f7ALiFk9D7T0xQUYyLkYwkUODW/0/7gIEkSGaMp4Zf6zwmnEQk6UQQ8Wf9Ed
6gPT9KtwgkLVBro9Lq4qHXHnzJjhwmJc7m6IVp8oAY6KVAODcCkklH4aW2RL
XIOiiA4WxFv10rako3fLapPHsURyVqfwZZ/PyrAaSgyoC9+zS+6afYdsfhfm
AtB0PAJ5FKknq/Ol60UTwpMcSbbk5xYoB//Qb0X8edSKHB1Ao54Fok1ifc29
+vSp1Pql0vqtxSkk/I6elmGuSx5AkcCk7vtGOR0lRplRkSa1K4Ns112y/5+a
dsnDCK2Mr14zw+z4zn0a/3dSq6XHnYMQoIOeCVA7n7P78xufEhI7k02P+09w
zMPtBMyz11b81VUoKgDcxAmG8LFv5RpBbudszl6WyFNhc5TZFN8KXdOvlb6U
dPI1yi7n9kMM6O8Jk1M6WAmt+AMHT3lngdTkPOtp5sztQTdUtkUplWtSyD4z
9NTikzi7C3FDxQ83Jy/vzDtw7ifWxRaxYxGTYrohWrHD9kO5WLFuL+LtF84t
DDmTGiqvDfTOmXpT6dfIDu9Z0vTaRZjPg0rhFwLDr+kSabvpLAvv53aowU17
kfv4LPQRP0lFRSgiJ11J/8SuRqzPtRuJQjKKoYPqLtkpETpxN/5t6StfasgR
+k+qcAduv62/m9oOHn32t0OjbOOJa32/h2r6NIpguh5/Lu4e+unaymCmIlk/
j5i6JIXPm0f3LCDhrkrHLHJriLC3/Hg3VPBlzbCOVJEnEksW7Nmjedn1R4Lb
olqxcbT53PVr0YyZzTMObTl4fvSG6jXchaFlWBG1OjjW6vSc4rW/scFFK/qa
bVIGe6muUlYYiomdScmnMX1uzzoJlb8lsxCCMDOiepOfGo4/pvRSdsd2FGJN
+ryhm+kd/aJTUMl1OxLfocQPY65oSFxrMc4Uipfha7fvoFNfAGB4kppLyUUJ
NjANCvtHP3osxgLWjv2uVnuZ0MY48jpJSoX1Z40NqHmgkNX4u2acCZtC1vVm
HwXXK+LdYttfbYrJNymBRmRGtCziVh2PU1Kb4jLXO2Qzy1B8tGU6ePZBL+CL
cB7Z1AuvcinlkVYaGV30/rdOHvfoizb0KxVfYrLNHKr3R4owpn/bmpv81Rdc
HZF7V9gR+g7yBXJUobHTweViOsNp+/twaCRtBRch//bAEsTOUpXdd5JPNSkJ
Z7PmlUHqciJR0AoQiYBsOLFBsv4CKwhBXM0pRH2aCFVOcYy62SryPw6CeTwh
JpRFEwrdTpwj86vFX88Q80dhl1NaZKGrW3yqizw8Xi1tZpVY2zwORnILPY4w
TzT1jFDQwC+k3YwgpZTdBEvm7m2CBnLQOJpM29Eoh4b0if5yQdKgdT5+7jir
sCThyBbH/zzG0+GbhCkVgPx/UQPrnetlBrKpk4A0uMFvq15BeT5ilAJKVNSD
8gng/T942f435mj5DG1RSurVT/cX0NbNrqoyqErgLmsiaBp5PWvHUUxlsw0k
aU/y0EYj0UFIsJML0XiJ2jcJgVlYNgkN6/S91PLbFZ2FQUw08/15x5EAOQqA
vYiTAaNWfmdsytL5NtFKguYAw7BLXp7LLmnyTIkdde+NOMwWiuv+TWBG9SqC
cvPjhEUVcaVNjMS0bVgZYbCCWxd4Nb16g7Fd+cdzgqkHttRXM34BuAtQcdMZ
XjoZ58mrFHWZ01Fo9EXJ/8neoinK6s1GY18H0jNpFsukUGfBwQDVeF0C9Hv/
6mSjUuO7Wm3u6ZPSoZEaTnv1BvOFo0yH77qiDIiPeZK07O8SvwdmitXMBvaV
jFDuqewkzdLbq1ydq7ndUtYcQRiR7ScrDH0Qef8qQN51BsVN1DyWO3a7DHw0
kR25/HtCnil6X0Dl88w16j3vZreH7qA/S3wYVoPB20oV8UxEt8XQQOZNs7jl
BAZUOg5csVUC+QIqUmLboI9DZhG50ORaOno4eg7V7VOoOPJ0bjHm+g2iF4mC
0CVJKRg5sov36Vj2CHEcTxup3RiqFYaIVPK88IzeW2IxTvdvNMA+nveyVGeV
YVSA4RfqIx0JDS5dPF+dw/VM2bJTzcHdmEbPs8+LTAahBLBp6SJWk039YWRu
xcU8CM2RpczrjvY870yfsXCU1xaiG1uoqbRwXR2/59BIY34kV3HY7Zm1/YcM
yZDUtD8cY6ING5TIhy8QPZYwgYcm0wMo3vh5e3FmaD2+xEBRWp/vXm2WfnfN
p5Dm4G6E/nWU9r2ovumIV8F5TjEklfDaOR5xXBjYBuNzdQaSisleEvhfh+Gk
pwKvrqZ0o/tohpLT/aoUjw+bTMzpvqjLhycnhFfUASUBJUihyYlnK7i129PX
KVfi+wyrgJ5V3dBcuH2PoQVy1gGdIMfD05sHDwT0/S/k0Ye8pjy1NGxP23rh
dGnuIsXB1J0TqYBstpseeddXXL5dIHv03QA1dPuBz5+mJBd1tV1VSjETUw5T
6MIj9uNugJsdSe+xrZTxanl5DscOmBGMrpzBumtiaSm0eP/l5vj4IqK0Dt2B
WjVNttcc4bbcUz3BKTiOQNrtkmJiSu9Hee+uFf2XO6KYUXiKucU6VFDsklep
r9CF9fJfzvj8RHF3a8HrYEPfLqhB8yMV1cRc7MuU7JH48APCptwXTC88m76K
bQr0WtW0+rzMNHeae0rh3x7C2T626+oQ7UPaqA5hJmhHqXjpeT3816yMHnUT
NoYe3xcBCct8meF0jq0Z/l1TWG5g9MGjxeQZ846EViG9bn6r3causcU2vYPu
7DQeVVKJxHILKd2jcKxHB8ONf/3R+Ayu3WylBB6QA1iO+QsHI7qcV3KQe3yD
fF5xxzMdgPEZfTo95le4zOi266nrldhZ06F2PWbV1SCr55deXd+khFpv4J9X
He+/Q+NL/kQVWVEcc8yqp/fZPuo/NnlL3eDgN3wY6/EqxxxfPw+WjeV9Ws91
EmkXPySpA91jIzK8ZytQUx3Zn/sq9NCPrkoNyAuaoWTe87SWZt5GFG6XTxrX
YsJf/aDdQWf+rRVnACJ3Ki4ABE2q17CmolT+jVhVRean5mqmYx1nPVNiXDYW
jxnnJbEED7c0a4MBTNeP9AoPBr8eWu/wAP9uDUcPD/pyRJbCh3Q7QkGPn708
MLa2dhnz5UkvZabSii5pEHOEnaP3remEqdlWdjmBwNn2+F/GTnD5Pmfld1vU
A7pYMMDhbzmQ+BSjxIL6qGM4pQWjPRzL3fz9QWB1PYv9+f9gtG5qU4lPHMVa
OCUPgxmy4kkhoHWRJFgIpEpw8H4Grmd9hqlAGCu+h1bG2L+02TfITffOG8Au
C4MQkDHHhTBV1Xso6AkpTYpmejbS0rm+lNM4Rh7MxeFFttHTUAO2ZIre+ipR
7Wl+BDAZELVmZ/dXPaALBq2TU/M2XnirrPEVdX/4zd+uXiS0YbK7O///hyTX
WzvdMkCRA0p8GIN1k0EVV5dZ3gmMjuemHRJ9HNuIZV9POLeqpCH6yRX8EGiu
12Y9UYIUH70bhyDNxlrUk5fZ6DMVs4NhvEvNKnsogTZbQh6nBUQmx8y4DKSw
nfs24Pe/eMrKpkP2Bb9YR/+z1bVo+vdTuBFYLS+GB8RB+X8zVY4ahDJ8JP3H
NYravirRTY87LydVSXKwjDAgVpXTaRRPexWtwwbzbM/pk1cwnotGAXvoBc9a
15ueuTaaaUBtAJqGH8viS4hxvbyXPGneckeHP+eTw53r6oaioejy0490++mB
aakNV1k7oW56WpR+LWHfv4AmJfDbW57yHS9ZBBLSTbK179rRZo2sPgzZgFu4
rOQSf4f/7/YAmUgMYMtKOt/2/n4Oe0vzVVmY2UoF18/MGXTIV/amwHXALCe8
nXeYIb1U6JWhwaXLKoYBF3G5aun3vmyq3gbDJr8L3JILcXJCj7IGqePUUj1F
MO13FI20dALWt0/+GvSTbXIUaiNQhrfnGk9xidOSJ6tbPeTrSu3RllHYpn/D
qnuW6B7to1yWyT2LffMBN3bUZesRI3LfDSP41F/Kw+Lo3vLG/zOU1l+I3QnC
BQECsu1WiTy/2LfaHYQiuR6b/kEjj8TGcMMT3oQWBWBaodYotmye7BMkifyl
mURUXIjVAUcn5QebF3+0BBpasIKtL758wsu1+FBjS2YUd64N1usWARwJzQpo
Ar8bCbYuE/EElcvZBKpIWHWn6dT7SYZxc49HdUcdsad4yx+FDpKGNohg3js0
9GqPneCP0DVBDOd+q3cQen2I9bqk0slWF4ciG8EWgTyzqNVTMe7fvH6g73vA
Z06oTKy2pXFMxQv2Adw2rWCT6pJm6RQ13UWm+Bf1DCCYcBJoOi5bPUczjoNh
WEfH+Z3wHvHZRoPlF/RvMcLlZ2o8+eJ5xY8+V0aezlhd0VULM2pDGU2OQ9pM
mBgsdetcQp4vKsoKLAiNZjgvmUiMb3V5T4zu8HDv4isJyLc8KAGrr7HpO7Ya
XberBvzhqMAPuPyq6Mf9DOFjeptvXIPw9/oJEr42Xou9fkTjyEFI37KrnSAr
SND4qUS+7cmdEr6Vw5V7B+FVUL/z/MhZDe0CfZ7VDBAH6+gUjNoMD+tWcFN7
OLhSEwdvQWRjVO2COUeegiyRLYOWOIsKxWf0bhQAa0iPrPdoM3klqTQWcYp7
OR9z1giLs56J0GafJQ8ZqL10zJT9vRvqMHg86lmH+/NvK64S+nl/YJC/CXr2
j8qT3pplX5uy9GsWdEv3SqTN3W29JAIDe13KyxvgshOOg5g21EtQde8Ik7xa
XWpyuDRh3PbQKvUvQnXmqs2Lk4q+Wh9Y2c20pfctUfkKes2A96cc6D/bNzun
jhKWUNe77vCIDayRzcTiDkWTC4PFyhqRHKeL5f0Fqo7a4/KDB+qDOoiu7DA6
QrYt5/s7n95BzAcl78OdcnvUMRlRwvgqUoQHGllUJsMoEaWLyZQrn9vwpE7X
YyEhq/nN5WJQi1toIErnmk8uvFTAex7GJmnXfyssuQS7ORw5qTmyKvBNgt6x
vAmvyPxB6EaK+Bftnb7IIcIIFloeQITW0bA8lFQV08cdQ8VGSUCAIH66hOA+
pkMmbNZ9kMg2bMuURYVYDw8VoNbGYT6ralx2spSLO54McEfy8+Q6YAY0fFZi
zd/cBYEnS0I3z47eQz0K+FR9chKf2Fl/UIN+I3H17fK18toLdQtmpvFDYFUG
QOdAiGwy77q5S+X2ONh6lHAit74LIGXyo7p6DMJb1wRugoXAbEqQJNk1wWi5
inn2SiiiTkNnnwtZa6oAd2i9BTBnu3MwAFmWIys1QyapwZL0Y1slgJrgEstY
nIbKmp/wuKGfCuSgu+JjS6NsnV5Bry3qx6GXohKYVTscd8F6+vFOqei9S9Q3
Hl0HE3ogaZUj42nFJk4kF5cwi1LL882pNafOZwEAERiPh+VFrk7pmgjfBhbB
eYU5E/axlFjarN1J2lNdzKB6DArcbgg0oWp5M/9ZACD+LY4l02FLc1BkeiKW
eF5G/0AWYAkVChgkKVTFJ3Z9CwsDQE8d2q4Mc6zOHc+W9s7fekPafdXU56pT
6/a9XEJSKeAK/xH6lGDa+oJITQ4kYYm5A3cmAZKfa0pOGO01qyFsMhvIKOE/
tPwK1fYv77GL4JfCypFhGABJ0JQExPs7XGGiSP72FCLOOLxDVo6IW6Gr90f9
F+AsouZwM0iXoIBiLqegjETc58IbkdDPwAjzgwF1UX7GrXUy8qnpqzrmFsZq
7OCaIgVm3WFuISPXPXINoM6SJud7t1B7jC7DJMiN18AbyyiOmjC7b9nPruHp
kaZ1LTAywvtWqpQFd6qxJQv4dxu7qBaR151/ojcLWaMBYvOFq6cogWXRjYkX
IItDtHYxOAATeAgLPaLH+s6nTdt+55d+Jp34o4qeh2sqF07d4urcFxMGQsV9
cemkF+My3wAMLmCFFNadxzanVe7K4o/wAkpXL6cYVVj5HrKqR7MplopHvA4s
mfeH109+YdZXcwxuigZ3R+l86ZMIt+tUSfj8yArM0RFKWmpyGMcWRf8sUPaB
7gZILwxCzi+iRW52AHC1hT8fb/ZTtCYs/q/VlnvK/Wp6xmXx5H+tUQ6kxdLJ
xu1xL/727Qozqv90N6nKhAvEVZod9zjCV7ZsLrbwaNAqIVTFXYvkil/vZQAx
20rmVvaPfX7yANDi4Db3+mMzcb3vYHiW24yah55d4gRsqMLfzmW6BLS1bWqa
tyZesdyJcTB7GIP8dJXzR9HttVHh/8jfWxA2DSGjgAIEB5EaCQ+E6t5Asti+
wKbWJEq9WV4SacC8v3AFI1sdlWo+9/XTvN2f13hhvp+G2IGi3GaqIIW7PCNI
ZqxYLx3luNGcFN8bWpCDaQMCXUOG2viVpQHFXN0tYMOVBSiR2ny9bm+MC1aW
cRszqRCIoRR/ODVgwtAi/eqxrPFwaGHyGgpfsqgfnbz/fIGvZyc4RTlF9dne
9GhmbUzL7nHKvt6VeAJ2qhOexzG1H6TAFaz49KAdk9963ksyYX9xmFCF5Rj5
HxqI1mboVwCS6UfcQk+8d0Fv15GinF58PjYfI5MxKFVmH43guTVsHNVzRrbw
9lLTG3yGmUkLZp8AK8Pi7W4N7Xj5zHZftZ0u+DHWMk0PUhvChxBAdQX/mbmw
2mNPADcqNTlWCUUkB58a+PXKd8VVlUO6EYLQ8qOxPmYpVX+yKi8gnPFg2+mQ
0Ore11psaGhIQIA9AN98GkmqoYZJM1QyjOPekKIo9rxJ0cAkB1S6gPQVkMjh
ZEu52Pjqot4oRIf1apUCDa/2EHwW7grvTMmnJARuPNCi90Gm9BZBuG79hG8/
NoD6N3xS7YP3PxCngC4CBDMFk0aMShLEHH6pp7nBV8CYF2+GrVvU76pQiGvB
NVwknFdbqxJ3ZA+ad287ny8mUI1ZBLARvHXJtPOnnVJxW2JUsZDFXZNktx61
6QO473wTCyRIyr3zdbrdO+QWx2rC+RpbSaKOY8PMRIvpwDjqW/K2vkISmonl
b7umLH5bm7+4uUmo+T+fRxsLopHJJqixxKqv0RFtzlQ7/NRDNwIr/fQBYioC
UoBxMPjeIO3hoUd7OqD5fOvCDWE0byv4wBL00Mnn0ybHwKGtMlAeLfihkucy
kfI7sXZd5iLd2iul+a7WpVNXzrN6QXN3UX0zgTbruQMEbQlDZ+QBgEjIVkf1
6nM8QPgMurHkLSDxl3f/NwHYcmtHo159lEqyfHbJz48b4ZNs1uvdwaKHi4jg
BKCgVzPlxW0H8bfgJsZMLm+jmGEkuDNkntQEnnhMyR1ds/6e9SF6BAZJ5HI0
CV0YNnFhI8PTANkMWLvVSTvQddiCsygm+IPqXlN+ar7oBxQQRkdqrKf5dyRX
ls1DogoVPziMjXrTReBFbn7f5xMm4ISwj8hwLPLUyBNYzDBZi9PnNEv5HfMf
nrc/Gnh8lhsraZtxlg7p4v9DstmQxX7dW8w2yxXb3F3sFXy8lxIkCZiNUocC
+CXGn0yxa3v0/81UNz0J3CZLs7dTW/tgLp+L4g37FfCkzclYrSrQM65ln5kw
pdRo7nufBQUHF1qU+bZbiyWEMxk1T+RzLJ6UOGdBp3KwacxckhSiGmdfKhnf
7CALdKGu7CP6uNBLxB624UvgEESfncrykcQVG4hHaKQWBd6M+kRL5ByXoBl/
N3F6iH1U4BFXHWl9YAkeJMgDPSjpV4QixCyG1lK7PP9rZeX1qv5xG0oooQi/
HxigoyxMwBKBVLc/2mRj5fgoOEqhWIvn+RGbzOiKixzX02X0dA9eynNxoiiq
nIMM67mtljlTFg+Hz4g4yy4u9tZvZP8cAf9sVCdOf+/mooMITA3dc8UM77Sg
oy2iROSO+diMykODXdpukuEdMBjoeEiz+8axlzJTcf6WB5kuVdWGTVh28qcQ
L7V9hlnG1A1wtIEKOECoLgmKcSNbTZbDLpAH3Br3aau7jnpHhuh6R26qbI+1
OnBB8O+Y3FZG3tGpZ8ZC8E6Rtl7iiY0it2dDu3SZ/qGLXRR9+7cZL/t5pzJg
SrDlIQ99KAhrCLzm3eZVxHuE9hJbRKsbqAhmZR+cNO+3IBQtxXnrE2bbuBhW
UN8O2kxgohNBVXGLDyo4aJhAEhbskxA74BHcsktZuMjvhV6DudZbxoC+CPWH
DK9+O2LsuuJBKnfFlPP3XGQKXOky52FK/WcXpY3hmPSR76UnHIJetwhybw+l
RrCxG+bQJP/ycVb8+I9G4eQixKwteSlsW2m4ZU/mfIHrchrnLmT5MiP/CsJL
+OeXQEustdGMxZIePD6nDVDyB7vDsuIznCAIMO7NJJsBPYak7pTP3SW5gjni
1Sq32Y2jDo9Wqro3JIemKdIxutKAn9RjPr1T6TygxfmGgKDlfQRLXBHdTH+R
SGpei7DsDgL9g0++Og9c0OQFTxFD/afWLiRTR0XyN/MhCMhwbkOuCLs0S7gT
z8icu7kbkD6y4SttZiLSL/cNPNaWoZWRwwhm24sS9TFalLdxOSaHodEeTNbI
vIKRvZ64vY6PmxzApsIB725eQkNsqyqJJEvVdERRgCnLOBBLYl4PL63jtVcz
Sf08BhP/6OR6tj6u7PjCmIdHMAWod3ws7JjDI+Z52YxqJNrxwEwEO/SmL/5x
1CegWhHtBN7eO2FtOC3cxTs+4ZPHjQrP9enOXfa2J/zrVQW50V2GgTk23K0R
q5FzH2I2oQh84W3SpmLG96OvO2sPnZyRFoSD9aoi0hJ1KM/mssqRMJkz29Oc
cFD7bZLZk2SZvzhltX6LF8PV2r3Y12A4X5rDOAjyoqv3hcEEhqo/oR6vxj+m
sNc/lHj4PPebfBL/4GqTHADbGbRcU7d/TDqs3sSvpqvQxyhTy6Ettw6Vflg7
te7EvupMVeAA7n0oULvj8Cxn6uU97UZpNDUQ/h6Lo9jvt3qIvQ/giDwalhSV
8GbOPmQmJJkFMn8Gp6KQ1bFsii3EDcUjWxICzoSoQ7HJ0nmeaNStNSa1Oeh1
jM24gf5JOl5w63RkuOSizEJsRqb1jCioInFUEMoH41OktLlvnVBQr9tNhpUa
NwYnLUXEmfwpUK8pCmEG8+XE4+2Cv8i6ASCa/ItsRdtYsecqeJ9uDSECby3s
Ey0t4rUbII0nEkSg8cqtOPMfSYZB/wMNgmp4ZO7PV6xUw2oYmrR3FIl7HmCx
wgtMfLM3eerBrP2OuBkmY0LTvrQ443cIfujq3mC5rUO7NtaTyP0s12kiyXmG
0x5i63DBrGIOSEkY3LS3MXtrv3LpEigLN/Kt2cXwOW1ml5Q4LmxQNtAIbK8t
nGTy60Jw9hmaX5fJeH9Tj+Jsw1KUONP7BCbEjvTv0xR9bodmAJQMY5dLAgvM
xZsBmGD4dTtcZcdzTFwwL67dBCbCYh1JZBY6O8Sa9TjSvjfyrV8t07iD1b+0
g+q0hb41NVqH417pnJT/dya/aUmda2MfOu6+2odyF1lMMO6o4+s/18QE5NjM
g1XThjeBKf5+NDdiZ61r1SaigCk6Ruf4IE07qJrcqtuFNmdgPXjiF5RDhsw+
qWbcsiRaWs4oemmHddPnm8cGln0+8GuMky2SdP8uFbQaRHlnNgAuZUMdFZ+J
pJ2703k4lOCHxYjHpgqzYpSLU4vieMWZMd/+jqd646xoOweymzfgWFc9KAhC
KtYrcCY2A4kafuya2C7XVvKQqQrKPXndiqYct55/R4kTixGOLJ+MMOeAzte4
+g68fC9KhpAe0gCAc/3NUj9G47SGfeAeyq+ibq5PQ9q5c9eqiYKPeha9Rmvv
tlc9nhMm0grrAFacf3ITErJPSDpAE3aqUdcBlcy6BU/1j9LIc6eVHC3aUbYk
y3iNh35qBW5ACs74KMiF4IZgr4PENHzrG48wGw6iacH0qwr6ZnDxeciwc6j1
lahl4jOZwTM4P2GJqfFtoq7u5gZ5jmJx03wob/U7ooI2eoVXHGXQ8DqWy1Nw
RTsLVf7P8a4tJ45Fn25dCTxcCaTlIND48suXftKx+qDKDJUGwzxwCQR9awod
uLI5nR2mkNFmaYg9GFXYqhv8ei5tW157XCGGUQ7GOwH6W/rHxMo0Ll/IvDdX
kGk0zP7rqH4Zr7Un2WKrz9fqpnQylChq7laECByuOsBAoHv5mDLZvO1p/gHu
YxNwPlet0vr2v+MqET22ek7JLs3lzUzcxKMKNqbokesUv9VIAlo6k1hK9MnR
QuL916fXFg367YHaRNNCqOr8Fuf6nuUrMFn9bmxoPuoh3WygbiwUXn29HCeU
C4YgNpg0vmZmCG6SBPsTZuaJ5w5Gv3LPEtWIH276E/7EKoJr9G44VKx6ZBl3
VqpxsdTt7i4oYZgFmKH6BgSXMoz/ssRzfwWzV4UPTm6VRLZZMSSQ79qJ2PnN
zQJbEbYRlZvcBcTupTxpa0njZJDb6DMSv2NjrR0OMuIOcHVxwZZsYtWxTjMf
p0JqYGjaR+OJW3yTDg35r4MH0PwL2VWo73jQLsZB5ycvdnwTwNPo+DmhPGja
nceT0mnKU4mpDXaGJJ77VCqHHW5Uc3XZPra6mIgo75W2f6tdZE/Y6gAvcXjL
A78mla11fNpUJ94fCxh4EJrWRNeppAqhW7mQS/lyEK0p8JZrq9xEqBspY0tf
1HKvTyzjBDVrVLV3OjNozBZJTB8+qWVXFiLplPK/nsqR9OOxX2xhSh5wJ8jL
Co+LIq9wsgzcElXUWJL8pdQRSsXmPHgRS+AM4hXtyqVsTLD3eBV4ZpSy4k+h
DT1d5hafUWqNSK/to3paNy28dcMjNukwv+uDLVyCCX/wYl8wAa/YUQGbZnzI
888HoaFm5ciPWMnJhAsi7TOD6giioRxaIY1IxGomWfAfi3ADysNKRbmTVlo6
KF7fyyhXkFMUvkLOeLMw9dzESONxxrfKB2bgCm653JR9mKVg0iOJeY0BTeBg
unJwr4LCBPHgxhfHcJ6MCXbRuFqUdJAEyhnVQtg2VNqGSpRZ0JH+dmBti3bh
SiX1GW+R9z0YGNooT4P03gZvf5GYA9P8atKsO/Cd1tZm3kr/2G6PrIe03EM6
7ALCa6BoLFvBONdzWI0yZPdotX1y8wCez0f0xEop4InS6huc8eTtj+y1+Ns3
YKUVdDtse1L1KDJWkxKJaEDnu/Z5SD0NyfUilljkXwCn+jHdHyG/zPgZ8rKw
VdzD5G8zUNkOiq1Q8VoCDrWsm5xnpG9XkI5evrfG9oEcxabF7Ht3qw4sbojj
Odpd1vCBF7TvX21YMEhETTtFtKgUb3wN+A406UuqJ5f72zk7KtsRs4odFDN+
HEBm5ndugFDKQyyDqi1Edaygqok0Xn9vMEPU51CTxQ9Kig6vPKUb0NSRpeHO
V6XhhJ3FKd+NTa+ThacG15krMvPaqtKjjWCfYLMoCtHLTbDxzHo7aty+wnGd
ZCF9JllteU4BR7GlESQ2cztGJeYzrG5bj9hVk+I03LpUF5Sq6WrPnXplcy9f
D8HLeXtWFRHe0k/CDqXlebihNubYkipzIsD7IgHlRl+FwoFmM03YUkQSMpbe
AJAjmUeCcNDkPgsQ+d+xpPNmySEZqHUgsNQMX7lyUzfojZZdPPRE7gLpiDom
jy1pZUJ6wYmn0gOQt99stTJf4Z7fiRqnTskMQTd5fuDxRq4oy2DD/ezK+H9G
ZPs1vJ0HiLl34Ui6RyMsb870qUPtD92e0rYp5eHf/sFdKv7nLSsLIvMhqrwx
W17DP6DpGTaMF3IOky9uLJDVMBvG29W/+cfikV26aXh62e4Nx+jb9qHLC0Ke
HHJStf8ftb5mXijtuuTFyMuj1tUdOIALBtLXZDRmAr3DjjB9SWNf4sczvc7O
XUaOJuYb3Ij/uUstqUAwsSjDF3DiI3TNxJsBllZcA6JdqemUXvvXF6p/D49K
e9zPFfnIimPK3NeiMgPdI9FNR88PuDhgGqec1pVoEgUZfFiMkjchNxXBdaqm
8Gu4djidUo4XYwuLXPZKSNibp245uYnvWZbhUnXVq1k2PA17MUGil6nLJzQs
aoIuymuIbB0ZwRV0faf2YDTV4eZkt2wDzCGPpXHJkbRLN8drIqHi3U+iZh5R
Ucu2lT6l/q7fNPtg8nezaPk+6N2BmW+13fRUrZQQyGg2Nbn3pS0LKxLWIgxm
KFiaNGxFktjPPhHZnAU5VhI3JvRPjblmXrl+v/Dzn96+5E1FK1Fp8cH0Exyk
9pedR0/Zs6lD92raWlJGkCwj5yVsNqhoWZqgR9lbrnWEdk6/o/GjjvT8Lz5z
M0yJOqKHeOtRrN/AQniwDK+bjmu7n/3A+5j8lg78jekjlS5xvjtztm7A9f/y
1LLklA2beHucdhqqw7BHs2YCEyTF8JC4fxKoJMkj9JMfpRVipZzHceuD+Cqo
8TFtNQoFFQYVNUhqYB4Wr0CHLnP9x0YvHNm3oDcJKnCfomGWi6xy97MS+uL0
5ik1iYKTrh8R9JTnRfREbRLdckQhsSGnimMlliRVq2AVAZFks1jo/zo0Elyl
5G0QDhhamy2c7xSD9J0CDqGPowDW9cIKDer1IIt8myJhBAHQGsHDHV9ozon8
jBevyu3/NPX2EMBWKbuNK2wBprfA/RytE4eHjjvAtj7Odrb9rxrg7VwcnJ6j
EShWmNxijmBgh9Obu+Q55ZGox21V5QFN3xkpbRDNbv8nwOVB8AmWmQYCHYcx
KtWI4izIxZq/gFKPJu9RHWT8wQLw0kr5IEvTnj41jAZ9P8kjKXwl26Ecft6w
LBWwBICFU6ceUYPiLSetsr362GTwtIjZVtlTVPNH0QhmTV0/BGkiQ3cLk41v
fzL3XGcS5yA4nQBEfdMck8FVfi32aDc+GiX/VLCtKLUhz6QCVnaH8K/7WJhD
fD+oIolNzETCsRMJlaFO8OKlIIH9AhOrD3S8MQfAaJxm8g1FcUWCiYOaGfYe
jzaMD2ELTWCHrHBgV5Zozv5/8bFkS3R7uY6nnMpoIWSvnMCUUYjKB79qxOJb
duk67XfvIYpLinlJwpi0a8Cj24FBTNWITg2z2P3wbGPge0mbuzDyElEyQtGk
pyxsia7nk9xRErIwQ0MGlqjgFYLknOjl3IyOiQ7vhDDKtixLETXZRbnqiuFC
8mEOWnR8fMiADh6CJrwMySabgf+kMQ4mRHpdFQfeNuiq8M5J8f6Ew/SeuAYe
T3w9w57xvrsMWhjHbpzro36LU9ULlCGBYlPYggmVfaZQN7jIkLSQlqUBEOOD
NuLT4Cfr4PYGwZNnQPIgsaFHSSdAHAHU7R8ujtujr5lAoJx+KH2kN2Zv1lAI
Pdm+DnNveT6N2uqhZL6iRFhAd2UX6xgnmed7m8jKgLCmWElo1OrU80UmkTpX
EqX8PFQdL4hmEsz+PpYwOhSgjVOhdX63EJGdGO+EImBCPp+BBItjQ8EKN6Pi
FgPGmfTDv3dFJ5bIx8L/KX46Nx4535Mo54tCTcI1UWAx2IypU/7XiRg3VglO
kSOuMv3WaJV1sFoJWIMg8MJEV9pinKEZEG5wDegAkARgifcjPNL9xmshA7p2
SF/hThDJhmu36HOdBOp4DOoU7BiTCTDtnInrJIKFKJIZOMA7cUIX1ME5f9J2
/WlKaFH61a8Vog1a/DzNbiWFeZ6hs7xnoDeM9ypoLrrxnBiBnDab87r+wz4T
kdnJM7LUhlatYNbdC3cSEI5bI8bqVwuVXXnCZDaFLjtnBtusfsI/gfaM2Gow
vf6JYPqsaZqZCPkz2+CNnPdXma1/Zx1Pu0Z4XyzlXqShrqlN9c8EWuu8YmxR
lDtBnc3HtsKlW5MAtVo+j4HN2CmajP5w/21NmGJwkGr8Iu/M65h4Nzwpsw0U
wesfDBqQwb+r6BamGfFDS+R1i1wAj2mbbXjT0YOMS9eTJQCVZUwpd0tr24tW
9mzwYu4cUQsW2MFAvl5vgqMekEkOBHT/TlRj4LEG2z6Qu2tzNssnAyWT3yRK
ElvI74BQ4HIYWOCqo7nboHuLSqAnOobAsItj2Wv8+OX7qo84fO2BbF2MGNAg
3FjcJRVOYitpD/QtYXgLBwJw73M4SO7TesINzgJ562u5YXwE6v7RLVZROJxF
as8kcCm81nFLCzEN7YX3/BzdBxWAqVejdWoS27Z8iwxRYFRaB/Ta7HfmKvHm
QwQxkq7JpCc4zvG5gXdu/m5Yb6MUWGrhnnBTHPvNkSoaYQIpn6Yu1HnpXbcz
PXhUmVRSfJcMT4LFDvjSu+ZdD3SI48Mh8/iXSttaOK5QUC0kCcOQ6lr1xLhd
mAMOTniQuD/qzDGcpbTZ4MdI6+043jm9c5aAXAEJHZdQaWqpuDpbqDcJRoqn
/GyvYd+0hPHn38QQnxqrYgLETs8VP3FddcJiJbFyTQEseZ8Fp1YHToQM1Jo3
UW5I9i0jcYOC5Y2pyjZZBZH1zJxf5fXIzfTlb5XshXOA0QTh1wnOYPt5wUsI
ycFj/V6OLWfMVszJing7+CqFVD6Jj4V438ql8/8wjjJKtktOe0CZRh41DGGx
4lMy+Kh4e/BoOR51ZpFTihP4G1F7djDpRsrKslp4638+6LDouj0aZ0Iz+C2R
WEwlfJgk8UmsH910Gzb4A0X+roly81Ckr6k+7tnpj1tu8IQz7Nqi1zjTKya0
J6HNf5mzYS4drmgO1maNEupmXVQsYyL3ZQHC7GRQbpM/d9EJDxg8IgWa41aK
rdxPO/yi2CnZgV5ejewk2gaRIzpP06+fYQq3cQZxp84i0LYIPDMwm7T4TawH
jtmA4/Vmoy2cSzzsHrhZomgDViIBm+IQoI1+agTN490FBQqnbLgYujizv5ma
k3xwK2a3YuqGti5G6ghZ3LqIMccU/tBMSsUxgsTP/aKxsW6akIovVws0+ZiU
0VjzKK0/qyq0Bro9Y63XtWEvcrbKq4RqjIxI3gcvaYvjeNZZUnnjBVhSRfsa
NqpIJ7s34h2Qz2tzCUd5PDy3zk9l0/QTrqnR+C075sjQSjirPlJG9myHbBJw
T75F2h1CYIE0236VD2ErWYV3E9DbDgRizFcwyKFmDUQDKt0GSiza1PNGGAaz
SfBd731iajVxUmgF/wvdfEjSjLoV+lELrGH1eYLgJN1dnkBg8vgw0uS4S7cs
gU97vcFQsYgTkVxk+1iLfWV1NsrIRMko+5e97bx1cfa2GUyYkKfhRWxnZ9Hz
dIBCsWd7D9pI+Aut3eRMJf8UKG8ZBBOo6EcbyjwguBC100tXAoF2BsJvNJq7
jpdC5+RKVyFhgF/G+UAwss7SmnK7/klTPE8YRtrM8oVcerpt+TqJvz8oIDXk
3WoJqw74Iz+1FJDN6JcQGkmK/tnoS4crRl+sNBLjC3Xbm7Fhq0bXsX2GNwYf
6kvMDCoeXwX+z+urQq6/qOSeiS+HAdph1z3QJlXQ0/OMj0Q8uGQCuo7nyl2z
N97SKirccVuz2tSrg4+bRd+KysLzWrknq81NFuyTE+kjA+CwzndbAkKDDVCH
/0tRMwCJZkwqOPvNSL5EQjvMthm7Gz6yd4R5muqVRzHGsm/LLM6Bzx0hZ9H0
RSpSUrY/xr7UTyphwa1PBhAXAjMawAcdG/QKbb3Fj0hid+prN3RzwRUEETIn
BnAOE+iw17GJUuhj7tw8+kCBy7nGpiSez9hsYxUi1odp9rRryj0euLFIkxgw
0nQf7/0XJfheJdj/w/XYWZKRnf0gL/TiPdCsiE43dsH2UUgnNhRmOO/K04XC
lG+lq5bwaVZ8tmvFjRp7BqWBTSnvWUuNDbicFSxxsEAen24WXyDqouSzebt+
PLzBNmZ5DKmn9K+7p4cYNJJgQZnvF44bI6Ukw9poT/iYdGALVn3O0B/hHDHC
xmSHAAUbEVN57eMVZZuxQCxt5YBC1gHC2lEcr4DH/MxEQM1m1Oj8qQSU5R4p
0qa88O+8Mrd5Uwk/I2PeG3tl3YKMJoN/MIOsBIcbaKgYVkT6V07HeTN8gxbl
W9esh+RpLx/D/emonFWsn8ucPxQGmxEr7qtMH66kV4p3xH69LV/TiKQNX5kj
H0Y6nHY6I04n5yQu+ANhSk/y8q/mZTiK0xizLms+8ytzx0w+A8VkZ8byNYLy
KtTT21fcpXbTUKjyhblTEFMp+5h+un8PL80vzyQtbOHYFTArPuiXissrOein
zKEuoRf73NFQ49aZ1Ysusnb/grHmy/R78NIVNdbuhUo0cJNKhhjK445Dh9/N
yQ6Uiz0SWwE2TL6qOEE8nYiYDlrONn55tgXvQ0OUR/eaoR2GD5p2Qq5UdDLY
kSUavEs9pDeOJMAnRb9KNvazzwPUYK0xCu7qFyFuZ2RC7X9fJea5/0JDsv5b
Qn67QbVT9V9tTB06guqwkYiDWpJdRUzLQ0v2HBT9MTh30dgDmrQu1EhpfvsZ
Y5+53Yrrkz93DVRLjsAEmb93xyn39KoaI2s9xnMz3+HvGeWmjnIeo3cxfA7F
UIRXzwzwagIfkh2gdNqqIhOVbXj5B+2FCtEj1VVx0sIFCY/CfwPB2QNbFD0d
T7NH/87PrAisQyTaqMoXqNnOEPISmWyMW0xsXniZU6IkX22TtsN3WcbfrINN
pi4348Hn6AQnGFSdujuhF2BUi1uEDXQgoIcsgkv2h7zFZi2zMK1fzZUMriWa
hKHGouixuB/rmjzsf/KNe+r4xUvUeYtBu6l+TEcDM8Kt1dkbAh1HVA2R0TsP
Xnoq8WMnSZKSNUwzBbmkqoECdUKbRGXpsnXvUi08g+cyUD2nAkvi+q4v9ofP
FaFwL6qy++rdvPxN2OSzeI11ypl88bL/c0Ro9d9AdBk3fGLQLilzQAkC/6Oi
8RFxpApUSO7OGm1PztpEJ2A2iVVdwzIOL9X9m0uONI5Ue3kFCaeh5OrUkU3H
bx79OFvUXfqr8x1PcKvXOwbV9C8nAosB6ngesnJnxPwkkWn8uE1VwYIyOUQ7
JZRGFXJT9YJBI1Cu2C9clTMm3G9u4wwRCWeDV9FtinUUVb3nE+uIjPmkE7mD
+wWy6kSisJK1PPBarnX4vL7F5ocE6F4pZIb9dGNdszQq0d8A8lZM6yZwb0vG
dCPT0f+xCu4bjxOotnMKTNHTBmA8+h37y5gg01StyI/8MbnaChXXAMeLty2+
4gXCva3dUeNT0tMhfpxGd9Zbdxx1pcOuoeExwa7Rt5rMDKsMepoW8XgxPlAL
t9w6NEgS6X3r/ybNVDJ6+g7p0EXlKjE863nGOXmVOFt0a0lWXryYp/RbN2zu
BvaEhgpuyBcAB1HmyNVeO6kKuhOb/GEyQbpq+0cIOcPKRqXzyRV87ZX83mjC
R8p9Jw4mS9rEok3OxVJ7EJwIB/KIgx6lOkmwX/oQkWsftVLpnaR3dcOy5wal
a1qc9U5iCVSpq6A8J05gyLWniADYP2WifyijdiXRwR7G7A38aP9+QocJshn8
/TFPkNOh60ccC/qTtT8Q0AiqcHNwbn/tPkfalhVRUNfsfMKrd4nMKhKK4vKn
J8LBCJ4/2n/OYgCa4qgcQXYjiSi/VJmJuc9/yKZHyt03Z+qxt17HyvPQRtYu
BaTbMtrC4e1vFRTgwNQvMQEUK+O+Ox97ctEEvoa+wrZSzG1CV7102tKESK4C
LlMbgLFOz6istcUCIpQ3FA4vXKCjjwM+KcZrqSYk4TwO90QDHhBwZw1nlgSm
1D6SZrlX5sYea+iDlb66LDsfP2w2x6yL96MlOdRzsMBe4U3Ea0U99/Hd9ypK
YDiSXCE7HfFUI57XyR0z0ktMY+gj6VWsAijVAHX/M6K9UI65AE47dEVjVv9X
Uz7v6mHLUKAKeO6JyargFV5LCl8yBM+VxPVbi4ZQqWjnOgVtQhtGNNDQHuor
pxJDAKKwEC8phJ6beN/nTGsM3qRAMV+0ik9GL7+oBzSnYhvhlpWFYhPyiHk7
CZtLWrkV6Vog7dTpHFQ5t8uWJwkbj/VS9rAuKS7r8JW8oMtBtSOBbcn+HHYe
Q+6yL15/zo9GWnxL734FFbnfRYMK4rJWFE6NVXVS4aCzCXCFGxBZMpnequbH
LFR3DWgVus3nzKVmDJyfq5zA8P9Kv5+xtewP03YGCx+jaEknUWEOxWDsOLwk
aBaEgbYOMsqzVUFG5YUKWUPZEZFhBnSawxTJncuoruDIyeOkjciGIXzj9jSR
ZD8e9Fl1ZfIzLDXUHWRtn/d+Az6RORGwCoSFhFj2WKbQStuyOwWnKNf+h20j
2Sjg1v9eQe0IXpWKZQBYlNt7eAeZ33kWGQiLC/xouAuHsm+tXiPbd9u9C1Q5
bjjvxCV5DdbhdDc3Q8gS21BKkAuIKMKdM7D8SYGQHr5FqiKxXayITR9WdGWs
5xMkTDbozYFHVJcV7Qkam28td1H3n0cxa4r7pD1ZWxlvMdj0PKppYhjmWrpg
zKuMZQ9UJPA6ki6zSSMMj22CLM/KVvrdVE5+GL8nglj/H/qpK3IilPsP0qPL
JOPCg7/MIQUItMLKTPyYhm75rdlXCn9Y5SrqmnqFnR9iAQLiS1A/EzA5dt+t
ndKno8bg4FB1u5b4SzYofRmykBT7RXKvfHjfq9ntMrW6GSSoPEGjcvzLXy+R
k/Vw/iLCLAbrp/7JUpAoB2PnBPfA4rOowiRrHr97mw+sZuNg0+qKTycFwS/4
eevSy1U/072PgGzgpRGnufFzYIBMBAXrAr9XPyshfLWnn16v4lhB2UI9inJT
Uk8l0iR6ENeJfaloUoVB+etaMLD3kJH/JedKJlTaHjcLKO4El5+8U0pJj/6w
pF9PdzhMt6kY5I/Eh05YShBt1Gvd1NlIj0p6W6dthf3fyH/A66LHqb5iklSb
6SP+DqkWEh9N09KOq/451b4eKUzxK4n/ehsqDiTKfKvcMy5liX6q2CajHJhq
uY6d5TzBDnQybuuiyIa4W+8HnZBrExiUKSrr0keIK7r5iwgJdEfAsbMnbJsZ
Rrzqp0b7YyML27c10ewrBRv45c4OrDKyVpLNUULsRJY3WU6YiOGXelcaQzc/
rQNFViDeys7pR6e9lelJ4x26dmDA2gI5AlmS+qUGVOZpnayrMZMc1+QQj6Fz
U4SOQ7G7XCnnxuEWYvWE3u6gSmArscR8P/KduML4pQLkycziaaTdXFdM1pMh
doj+t69iv7m0fHhI37wnTKssOQmnoVPRUobOwWRVMRAqqysYkgcqE3PnEQH0
4gU7l01XPWS3bEif5POQOSJv4SWLf0Vk12l/kpWzIAUxyw80JVWXdHNviGgO
rUr7CklFEP+o+bQKeG8pfiv1ENkca0uz0NExvx/0obqWS6Ne+Syes864P1Lg
dGuHnBGGz7aL/hVXB+0F5TXDOwzJLMbM7r7boOqlRd8XieazWkk9d8ecKjXl
2hmDFpobiC6vetypd2+b4l+xw2x0y75lKrK3OObSH5MdGucgYX8FQkSh/s5F
9tll0cfDyNKSO+/iuxAK4M8sUMX2drfbtg/LLgL/RmVvaHDypYUSchnmKbhP
qVOQxYEdhq9+ii2S8Baiyc0zHfghiSVTSv0fCrHZEhKSIgAHHRsRlYMcCq1H
v9XJQ3SCTUx1dNyvM041kM9QzUVvppEgG6Vu2XDDfrF1scPzsw29DHJEIj0s
cmb3IW92NB8BZ6MYbLBP5nEEGR8NqFc4QaIHkxVUowvzZOCyW1L7r9RmYWF5
zJfSketha9Zp6raF8ASxfPwbWSq5cy5bmWQeNBJuMywia5bnEl/YOJGWo/uL
cHpFf4lZK8MgDqnfsEoJQtVrrbcyNvkFoYbEmPsNqFhJHor9hNySyVzH1mTS
oiXn0NSdTmtR1UNqJCPn4fJd5wL+ThcULwXxuYq4vw+rAc9VAvsBLx7Zu/gP
03Ok/yOix0tkwiGfe4JIL8Naw1onBQYGqxxKOdyUmvrFAU0iEJZKS2WgEJGN
Bd8GYso9e4bLyQOu2RpY9TxhnTwnPTfWNVd01jD15VtJd0GQPqcC3KQmEPza
dYyZGAOIA+MlO3kwJKdRr3shkqhVuUKo1IF0sKTQp7K8Skc6z6yzTo2QwjNE
p2k7yvarn2RITcVdl0glwS0v4uMkf8FF/KiUm2CQHTR2FMhjZSOOwy64Qh3o
5N0Q1bay2aau2+5VduZ9rRzo+GLutZW/b3BX6oFCm76punyV6RRaVKpMtZMe
mYB4vUrVKvxaSg3wIa6aUEDfNHOkUTuEY3rdiaqLmbv47jdVoODWLQNw61+j
IjbX27TM9xVNqrh9glZY6Dmk789KEtUbwRP+piZDuQRy++ELNAC1vvjWbj/F
xke8hikhY7N5g1LUgrOlGxKwh/FTpxNdPGXHYa2zxOm49LgJaabhaQco6SUy
7mxHDjeYcfKpYqsXOfQ4lap1kyHJ/xqe1GMYQphppRUWy78Htl94nTbEuhje
LJ1OOfWQBG7KvjLktLPmd/7laI4Utf70SeVTPz1MK7CVW+s0RQUQrNzuphaG
b4jdYLdQxfoQvcVHRsynCk0sveweqvklJrrnIphovnS9hoE/bDzlRVN5xB7o
cC0UrKpa88x1wHHDwDhXD6CyRO6u7Z5H5cBdSdju6a4/0lu6rvkrZhUcRXzv
KwD875S566uUnRlIilE7jfMtWiBhEHDFswxx62sUwfldILjmPsa4z1MAeb5O
OQIGAXBPRf2/tPktk1ng/3AOVAP/ZZuA0NppApM7zHuBjZSPNsNI3FD4gtlX
ex7eyNPdB0EroXmDsA9W9j+9YhQoUEh+3SIrZm4NwilZmGZa0QP39fPJ5ysK
d9kMyi/EyYj0vW1vMURXVm2xXJbkKBlmXkH9nQkvLk/bDKwd+VsAYTKwM2pn
xWvRp/NJ1eY++JSdwf7Q8UeWX3rM9dNMhCRvN2M5HtR/I0qKoVRroXg5bjWU
tfIkYV6eKQ67MbGsJUhgwkBX7BTfD6B+A2yvbmOTm7ub9Nikgse6ootAlZST
ihZ+VMhc8S4p9QnXa/VIGT/uGo59qD/+lLfhYfhd1KvkDBIb2cMhL+J2lKNB
O+7YrM611JX4o3gfZ+a7cCVIv4qS+sh64YQFU/LsorNk5Q/cLWCWQPLCEyVb
YGtYm9w6IIbvihHeNTcRREm7TLe6J4rbDtiHkVRNWY8aeLM5vBAX3Tv67sfE
0K82M78CB5aeuqJgKkQSvO0zRmRq7UQkptRVHqRCbHoyirBWqPF7B9DS3hfH
2V748rMSoJdccdJzNfv8rll2/ls+NWsOrJ/bzmCJProDMcVCelqndoCCP/Lw
2qzWlhbKANcrDltmaP8Ry1KkiYNHn87ri4yB/CMBBjvUYwLFxVzkazJg5zyx
i8VS4BtU5oPEu6qDEMfkNY0l6SlizSx6KQCW5ykc3TDdxOz7zXMOYl/oEILZ
Uhmyi1oyKbRon/m2IVVzCT78Y2s8Tq+p7eMHbNsO8PIhZb/dGmqlD0FyhVom
AuwGYUZ3eUycgzZQaf8GQZqBv7MsUhap4FCXa4ztw0hdLgBTR7vcpluC9qZQ
Y9ObhfsyVFtBvyjrXWoMpcCq0VvCr4ECtfl4ctEz7qwqtd/hLbi02AdZDlLc
wQBbh2ptimdvjSz5LkLWu92u7eGjTx2N7E9e7vuDsE77tMrJz6LYCm9CRz1+
JXQZMfimLByK1/NTriTvaqZ/RYUcGQ7lHQQC+EcXJpkyzePROPEQOdeTS3fr
MHHfUrjV5xK0dAspSP6JMI0+5vEbX0MvqgtB0PysJDeJjsK/ckLsqU+BnzT3
YAaeAF/npFGAbqy8RiAMLnl2sadwU0b/j3slZ0t6RMcx5ijshjquyg3D+su9
RgGWq2kapXgsswVvH48LGmWzxEhjdHFvwJBIHOcX4KOnkgxatCFWi02+K1Mg
q89oBesHmpA/Fs8hs8Q2Inrn1lrGm4HnvJy5YK8SsAwuX8pMeR3/SymiGjbT
YwgmenlOYv+INe4njDHk6iPEXI5zAgcVL0Npjo815D5DxXnzzq3KKP8NLvPI
nVIv8F1zq79fGY1XpXTnhoXfLhW4y72uATpzkTAP0VzJaEuPZlAKnb5nRhJc
wcdg+eGUHlqjOwEEPf/jjPvuAk/XlZCPothU4G1Qp6q8wqF9SVDCby0LNpgm
k7vBSxiyBeb8qVtpp6AKlWPIdVnubqZm/GRZKF8OFDz3aY6alY1zUIBbnKnk
R1RIzCNBo30RyPRJOcVmA2PYu1zCsnoJkLJjBYIx7ikHF7+mLD8W4OCxOAnX
J6nECIbtffC/rPIsX775Qe3MmBVqVCLD7YVbhdK5gEZ9GGL4F2yylrHXOXO2
SMd+0CAm0iCBdJKYpnjFjaS9YhxdoMZIc2Jvg8lD8h1S4hxbLk2zVTQICajr
0Tbea0JR8Fbr6IsDIiiUuy5X+DeSkqAV3sgSUbBq2cxxncQw34tm8Zt0HFkS
ApAfKN4jnzuFPoVazeab3tAaSqpadclmGQ02K61c0LauetDaBZHTQ+iGIyVq
JCbhnh4f8RzlrZDJJOo2JBomFhfeXDvkZnRbfncaV+gEJypZjYC5/6l7HkGN
YWT5gKtf3D7TrsZHflyEtjdV3VHHKlMKzBgIVDR0+3+JBpOxnBfUjoXsJl+y
PDZ/zD5rzBYZTZL5s7meR0C/T5TBi+wJ8sjhCyIUuu8cDXW0OaBY447PLG53
9fLDCzmj4vP1C9i0zDwkEj4J0gytNBO791iyVgGRrsw5KieHIW47xiuj8okR
1klt+cvmwBdtsg9GcoMYTcR77h8365e8NoDRHOov+nK1S8pzDjOJX4MGIjeQ
JoDByqgbITs7yqwBrnmWI42jIz+DDv058xwvtZBTSpfOVx5zuwEsR9cOcTRY
E6VRtV/VKWhNXh6XRo3wppyWWlOW1WDhgGZVT0Y6TtPdcIHUeq+s3JbPjQP5
mq7283dYv0+hu9UJjjVhyuBRXk/VX7Cu5f0FEPaYJwyj73vhPEzdAr+QxOWj
HQJ37K4nCPuGpSKNeRlo4W84PBEp8YhzqtyLHDrF4R3ylMxLqfPS/BLm/kLz
Avz4k/65s15dMU/v1waUk+MF25sr06+pX/MnWj0s6gPbI0rp8442PVeuCoC6
H5TQVl9Vd8dQ6wjbJJsGydLIHhTd75k7KLSrM616W2IwbSD4AD4ZB2l/W7EA
OYBPLeLdHHXSHqJLtIZWMySveoTikZfrrQIBbZaXZXS0fSfC6PQtJEPBhLmR
ntIYn/z6ubc/jzllVtOGSbeiDmeGeunsrTc0chu69FMf2CAl99iHgo6OjSHG
qbrL5DSBrMusVA/1hqpVYfSdM2u8bR81EPA3tWB3p7A920O9wkH+3QjDDRQL
xO1q9GsCii5Wrw3NozYsgOnupUmI5SqGaqf4kWAR+9y6MXpcXPQ8C6DkDLFB
zXjNxu/bLyk1a3muepV7eHXnkE631fJHybcL3B28UQEzUKkZAjyDCp0qIw4K
BQ3iI4sYW2IdMJbJTZmQiOTvF0wAgg3gJ5amUvS0t4aZ1R+olxTnxrh+Pth8
F+Ijrg8vsyvMwFiwW7qfHApSZYoAXmzaWpjlb8ZMZI+7/5GVL4YYnXG6k6D7
lcZEN+8dil18Fu5L/DEHcnTDbx+CVhhQWzCa2uAny6M9U5S4t0GQlwKXvORK
FHeVTAn+Wb7ZxC5sEfQ9Hci0uAA84cy0TL+8LOB5l4TdTBO84C6mKE+wjcdY
h4NAmbthK6ZpdBD0g4x4v3AZjbysNO1+f7VEiOOnoxypndpElbq8SjKgtATt
9UHCKuNnrVatmN/d4AiHL4+CGF1x+1Eml6xVgQec7l1O0wAPoViBzEWM3kun
BvgYc5cek9wgNLwxWwxhdbNZQw4OxwtE/sb6s7J+74EkhcE3R3OWxpMF9HEM
GPrOhptlTAeTkR+ihHB2IP1iKloUQ5J6afoVEc5nrvtV9jiTTOewtygBRgp+
qskZUPkGPFH2OWRNLykGSHDDk5FBaDO/kqLP5FWtJEDfp8psk/9ynV1rmb9P
q9b7Flb0xr8M6JQXAzcYvUL4j/Elntu5Uxa97MDfZllmTdNKX9GLM8aoELbK
YC6nUp4NGEJUPhwAgxXxYYqNxLCOv9uhnqEVlusPX4DS6YRyQIVhpvmJy0o+
kCbogQiRwKYduPicxU9xpeq4dzxQCcpLOCYvMjkWP6QPbSMqY+AlmYtnVfvc
9hOXFu+Cs0pmqyekadp+lyzahhmKYfXKnD1CYmaEUhIKYRwnD6bjZQ802Y35
VwxkrLILW4/LYsGdmthaDBJ4KGinIceXfN8CPHXyMJnOIXcVwTutfvtziFG7
JzEYCbEgrKS1cvlTPC4hgCSY2fc48g62W5QV+9JuScowA66mokTAo8Y3poL1
D0enRw2UboCaqq6KZ73rnycZMRCc1sEur82diTZh69jujfHDfoybONycPaUz
KjpDami8M+/U9pWgCp52RbvlnPdsBilhZzmDE2gk/Gmo8iHtJBuZCWyuVkTe
bJ3L+BBieKi9fMKnnQaUXM9HTQTYk52TJgtVKDnOd+lSjyYq5+7O9VPMoKCH
O7aXzrgZrY7RD/BlJaWDFh0SwhZsFKD9K/epiaMVS5wuzomh7S7j7SWXlX/z
0bSP6dSqKIWRpF/k1GocHYyeavQBCV1I6Cn/dB6Wia1lgGfwPmE/GoBKZB3K
KFI4dfIVKrWIuw5JXvrDSkx6Hd+n/kp4Tn/Gr29882YxPsbMRdn4CBFp0QOK
VSI3Tm6ZSGatqQrEIWU64/hdiNa2ZOe0kxNJNuYqxqL0JIHAiFtsQxLbyHer
IFU96OFjxlb21hg3x82YRX0upufOowezsqCw+vjylv6tiVVYj0Ja3+eZiFK8
NLLm+xySraTaDt6EdZkwploBQ/dUi7YLf08xAYnCmluYjgxKPKKIy6OY+F/c
ywoPbgYliIWV5URafNDzO1Bsa6gGJFSzSh38a0JuFqu2E/rGhKEO2nU3sfLk
VxqcPBDVgROvB5coNUJo3jonV6QqNmZCqK7pd/DbSUyDVe2kLc66LAGs5gZU
af4SVFFTxp2iEWhPX9u9AyKXw2OoNBd6FnzlKPoUPSXJSRkbAzK+vIHXybWr
Is0h8L5niXqiyf6Gv/Z6d6e8HZeu852B9iHC0uRtOMzcz4odFaZGgvWMxbC6
N72y38kF6UhyyO8xC5G3FweIayeDz+98V2ktT5s2pS6PfYq2vSDhs4jUqnm9
uhHpuNb75xR9zUC6Um3tTAa9Qai9UO3R/nLtztYtNvohhzOe6yXcth4ME4UA
G3tHZcd1Hq0XoAkvvd0jKl7V8WjnasNIMCYZz+HwPNOqeN1RYjPr49G20DoY
6Z2AAaJot2Ti7dMR/imI9pEX/L4ixdK21dG182ycZv17nVlJWmsnunKHWyyC
czltnrfsre5uMlp5TM4VFY2z0xSAa16CDrinfTh1riUNFaSx/V4Ag0n+Ttoe
37NHTrDLjSsXD33cC4XA3PB6v8uvslCX2AEgSF3x+L8U+1gNCi9BJsrulXZT
FO1DLNTYbhx7AS4ieDuwXwAXcCIDq7f1vydoIIpCg7RYPm/PkXPgockHO8UL
mf62981NzUGLSQcaXNf/qIAiKjoT7CKINLk9LE9LshtQqnYnLYbhpOCtFVY/
5S11y+Pi4DqapyDYmik4zdQTnTyTKDxyYAM07sy3jQSeu9VaFGmE7t6Fa98Z
Zioqc8Twxoo4Fob2XtXYhZMd42IKB+fr75GrABlzm9doJaFiEWU35MqaH5HO
OmuQj6f094lpnKAVm/KA+8WZFP1JEkRfb6q0sOzFnuFRotThvaMWYq52twMG
LaOIZ0kgd7R8VJfLGubtMQ+BoQIRjPjjKhb3DlYCbGjILyBkGj+r6mBbgloX
QcQeiW1kiGjpgO4IXOl0CoY31ehNBmq4/zLbY+YdPZAV+5yp8ReOlp+pkgAQ
bn/WI4YZAvRWIYNwAVsMW7KdBFP4Nqx5Hb77/5ei3zeQ/L6o9hRcUIdkgrHt
ySg9hd+w0/mU4npSTSL393xvNDGwFE3fgHsDHdi6h6HdM08mV4TJ3irrvrRR
rUKq4WzK/A8nzDxxYvClOWIkvyAg4H3pKl0KrpoJVU0TjoMVLmNSWYT6iSsd
vighY8N6gUo7kv4W6Dzem3nT1vN/2p2jBiG1Nx8BJIUaBGNjTngKH68oCOyj
fsqy36+Fn+9I/ffieqAZrWOu+468gFasUntGQl2pOI3pcA7XkI3Xq0ZzoMEH
Ba0JZgeQRloSiW89iSwMf18Mcs0v5dwI4Yo9MJkj5wDxvdHYwtT29ge0xslP
lBl7K/tZ0Xq97R0r9tRCZL6GFUvpYQoZOwMfWAcLQEa0B7Uk9SUlVQP5XxmI
XMw/2hfz/6pg/oUmmtN0EmR6LtsiJ1sKKwrqpm0XgLdkjbD1F6jkqo97g623
LSrjJkiPH5XQd/GwzZJshYqt7bSBxt+V1i98vWrDf63NmbZeE0qYv2HE8/G+
pcTuOQTNBXkm5D1c5Jps2w5udLbOgaMa5SuaA7hoMvUsiaT5MiqQ7kPHEAIa
lx/O71gBEPTrau4Y8OtXt96J9gDFRUJT9svTJkLbFXNBwqGiWlKoH5Yqdd/C
FhPGRPtP8gLyrJr+qtl1ScT4ZW4pMcjcEeIeJQHf8RBwDMi7u9pCXHhEyI+Y
dai0u8FhiikhKS4165S0PqQgxjlEgUl+wtd7zR35Y9z2Nj60FVFi14Nz7KId
1T0AwIohL4ajCvf/NX7M6irXQdhPsYzlX+ZZ3kYbqaTuyWPCcw5HyYiXeQma
9RomfIxmBFt26UM4CUWyi8Dz2DUUvXnKkyAQ1cjXTMaVNTyRvrNmaBXQbceq
pCR2kDvJrHxoTwdRoJ9CnI0rogFQayUHhXSgJOslTK7y/mewKAezta9/oQiP
1ZO5CoOsHoXVs2fjKhPgicYlCLoX8X7v2/t3hunLAbRCH4xM8Hv1M5r6awlq
GmMNXVaUW+O0uJ8CPwHd4w7Nztl0JUhHm1kge71+qvZ/kpJkTei7KE5YL7i9
5/rgG712zo08ho/vJrlpqd6856tiCsLdroig/thQEljZp6Lljfa4azdpuW6j
ns23+b4k9/CLQwZnZGTEnXYQsSnG526fbKkE/QK6SMHiAZRjs6C/GhjEVYyp
jD9He/D6u/gnGt2THtVjB40g0k26dNFMoa84yLl8PPOcRjnwMNoYEDw4mrny
9tUDq8X3Ch6um47E2bNYFAq+8jl0Zu02cMz89aNt8AE9pc3LY5pBMJ3Aw8PP
eCLxns9agTF0+i+5dARxOpeWrqeuh07PcJA0nLSTv/+euyhG/4GXCzZYKkKv
mpjLkIshl066rNHwygtRc+7nd3tGWenk3vm/s7yE9pauLbhFql9Zphb5SIHZ
ioxBi7EcfseMN2mi2SW1jreGUn+J4wBl1/sCqIR2m6CkqxD56FKgHMlQaOiu
TGMPRKPV+6ZxI5vN3iLuOQCeSOar08kC1CaC3cJEMqtyEhA+ncw9h969yGRp
/Po6ImtpA1wLllpCsgyE1EdrGl+qv57x6y2bCMvoi+p72WTXdlpXFF9+bKZt
MFnDWe+YoPQ6SuhxwGURJ3g4g7NrZDZmVhhMYDRwp6jk2mGuGxANe3xfl6Uc
o2Q3rclkVL2DksS5CVL3FZbtMtrOuXq4aJfk/K2loZJmzH0VSIji10IZQwri
B+6+K2CyL9UPR4sxeTA0xqpnvRm4z4BMOHspXEQ1jjhZiUefAqfuMXtydEOE
kCNmP7ubjnGN/Flv/QChyAbdGE7H9iO2ZCheUnV21Em1dK642mXSr/tt8O3a
hbR591aFa/NIT957fAcWzonT+DP3TyB11M/TmKB/4MVqP1RslFxcUPoPfl/M
QsVGgsxfHOLrB3T8zkyCJN+LItYdEyPti9PWCcGtYregOlhqmHKCqufXGqyH
QR+VaOb0WbU6tANWfn1cfVzp2RJ/lLaZPUY+2hLrRQKZFBFBhajecIboWwHg
8g9q7GqBquPQRe4EdMWktpmP4pWCeUr5SiiDZ190rii00RqB+nYCpj2JefAy
1++2Yed5WO2HOxjTufhtK4NO1bM9QnxIXFaij9u/nVs+Ii61IXX5FUN8AsK9
t937zrlof8KtkAWa0Br91d0roDTCtTlkkJ4ekhmygxM/+evm49u2yFyqcwBO
jr3gcDWzyNC2C3tCNsWLHrpy0yZEJHizZbWfFRgaYjvHFD77quufLFXrYa9N
4bS4EoawSzF9nXgqcwpbbQ/wkJxL7g8imhCIVj00kWMNhdgQLT9ecQ4CYgK/
qvUOhb/os9csjPrGje8W8rIA95GmH6qDB/+vD+Ya3bd/2+swQ7Hfcq5S3eP+
TPlbzrje1fANgmFy+v93tSui6vJ1c3S+ZwTnCsoZP2QqQK6iZ6AV3kVzdKpk
3s9Z/UINDGhWBsU+3Fin/I8Yf53sjkbY443qjf9FJNcE3MAVgayLWXgmDA47
nIeNA/I5m9hWzdavzrdQBUohl4P3l2z65lPEV/eIcW/Ko0Wqr4+X0iAdNrTS
mdH8vxjCCMgd2med0uxL8JUpRVxMKs313hqPIkIYHa8dAMoWrJFPt2g4V2jG
PD8DlgMtHadWXy+J1FPt5gSutmJsiqeDm2No0ytHQXrmjnSCT+bqLOc4qdbN
3ODl92DOvZO0GHNO5WvIXuPkhO3aZZSgUmrd2npzXxvgOUqVurMZZ2DXOfLv
qxLTIzUsvcJGuDr/lN/d8iVqRrbE3yLSGEvnU44JqjaVW1Snmg6Schqt+S5p
OnGN7kZiw4sJ/q/7Xlk/Kn7TRfBylnOE234ipg1mpxqud6uGWrX73VokygZw
V10S2CweLhSOgmC0ajxmUEBm8ZpzPHnWEP6XccM0Uo6r1te3r8CPepBJzx7E
Qbvfx+JvfZJVQprWWfKhG3RBMP5BdYFluR6MG3Ljcrz26RkZyguIi+S0Rj1K
G/+Lm1b+ZTi4yNKXVNwlavg6tq9vSxxKT9KNUbuQt93O5TYzFt6yNg6gbXQs
bNZPGD54FaeVYT6KIR/9GdZZg01pFt1cLkn5LDf5BgDmMFiQYiZO/SDszuAY
arEfVb2ITroeWItLIkfO6GDlvz9eJ2R5I4JfaacZhNvsH3aGIxopZXz/sIJ6
u3C6mH6ulZ5MJc9MCYQJ1Y317EChQO2yklcQHe208IETz2GfoZESftO7SnAt
DKDk0YArlcT5O5hCE3/5fN0f+U8OtTs8B5pcbtwKW9OUL3q5U5UhWha6Trc8
WUtsB6kCw0m6IB//erk0Ji8S9LJEx0a5+BYiNeH7uNo4pymZBzJkgAePW2Qv
nsxZleivr0VTUyEd6EJCkjydNKzOgQlcE9gOTDD0+AFJRVFCv4RhlkInjBE/
wS6NehFKqT7jlqaGbcHFUQQE621y9u4Hdj/LU9KRDtFCljqhydnir6HRiPE3
FuqXwTcgm/o1Cumx9OUwwLGDt+f9RrsGnk4dXX7B9xKHRqXGQQ6m7WqdFKjX
OoB4YV3o5SZgDqQALykAr4QbcKoy+8irFhu/f8YwY8FkRoyHDcVHhBA33s7v
ViNJMAT1hbHIQHLR69ONR1R1mGrNumy8dJpVxj/OK4001u1O5t2lZtO760tV
WEcXRp3Rc0Y93/KnRQIgURrXbNLA55PEXpfQ/RhoRq/L0Ee8kDDaFhWaQnuf
498BCivTLmGrr4cg2QoIr4SIF84qTrInzcbdMFP3tu7Ke2LgiojYA9KwPtp7
oG4E1PSSnI44jZ/8Y2hAE9ohbD/QlBJWi+HG82mSpRltybptJnKFTxmAU7Ad
tD+EcvTOBp5nJloNXcsCK2DPlyqQ4Kcl5BaIR0FXf0XbB287ZQ0QNI1tTFSA
Fryrhv8Crv6bTGYMpy0Ko1uKpvuNNLMrsxMQnThp9DeV9WaT2uh7CJSoE6Tf
hfVvtAcihRtt3hIhg6vW7bg34/GcU2zXOD/6Uvz+bztQgw1UDCxdLgtiB67k
Q6RTFsKyITQiyzPnKTT7L9vbfsoudgZRNill/mHRK/r0XdP9CeV8nFrsWh8V
gIXGc/vJa1FouYwhs6G7QMNCGj9XPFWFDd0DOU9b9N7c/ckfDCM9FDWyWiS8
E7EkNUiPhbLEXVbWsd2f4IgALfX7YJx0VqBsAAMU5CTkdvVuuSg0HajLvAjS
WniWIk4QfSRe/s4feKRgQm+Bz6SgxTNNZsPZxSEDOZ+LWm0YtkYMy0BIqrfS
fJY17oWwMzyA3Fh0KbYNRVVT9HLwqNWc3u/UfJ2DloHy7I5tClGKRN9sXUEZ
MUTsWnlqcToq0NQgKTNPJm6EOIiKAIPvaT8516OlU2xoKFTYeHNv5944PfiP
0yi0hejuhOkjwnj9RWbjXpxRd60QVq3Qn6OtVFmDQsSFp5FyYeRvSkTPl+pO
QstvjAYIG5NKEWu/bsPJVvLhj9a08K2OqD5vJc6eUpH31YbiXiFTojTFtojT
Z9jb0LWoWFhHClJtzK4+sy0t7Q/1Jhfvd/ZlyNfBIiWrdr84Io0ao88BYd2n
b+q43m8PntUkal9ytolFpLtwY5HlJSO7J3qPhRONOIemRWY7mAJ6yN4RyjAN
0AAdd3iV2Qn7uW/JJ4iJP8YDvbbvfphqWTbXXrSEzBkxq4wZVe4xnEZWG4Bs
KnQXfjbq98K0gyCN2sEVFN5p6AGX8Ai+6KFfJMt9qZ91FoRC8L+GWbtxLHLY
SYsy60XJ3a10BTrQSvzG1y67h+s3axlz9+b8ifxD+y9yywTC27qqscfT73sl
M9ALFiOCQCGhHGxw//238D5p4Tpq+PuqRltMJdStiXAfQJ+fOlQ0DQ+X1614
FtjyV2fkjAq/wyhaWlPW/3LOi0yQaNMMhfF4i+3mVaK6VlxTiU73g5xW422G
bolxsJuXsSTWWKVkczX6wvyhxfQvRMesWELbqxGhU9ySllxGANrOZ+ybl3ei
Vf0c6+TJs1XFOTJ58JDHAhHshkBPq4sYXUCOt3XuARG0VD/yf2wfrG0Lt/n6
NSzuop0D8d/b4L3RLdxoat0ooq8LhuVNtxzdqH1HMLKdvCF88Q2REGjXljNl
/3g9iau6jnpPbipy1A4/ceIw+AP8CmFw9BYuAquf8AGgtUcN5zHTxJXhpIW9
vCHC2L0YjuxzEA+nxZAeFG+BbwxDpgPiZSpmvg68fNg+jtg3RLKhsA3lHGcm
E3XOsi5rjLIcke3t6oFPWj6/TJZKXHFnLUvx/UdUBrmruZTnN1nCjv6GsL4f
YjNPE6KxWsin+sj2tygvexkKRqlosWWuTbNXgXFM14kivTaCKJWOz8a5O0j8
VVThVRGhoazLCIMGtg1ny6ks5vaODZwCpYTt5WJqqhmL2sIv0RVTWC3XbL7Z
cAoriRVh5VCZ/3NN3ZrwjRVBk5TxFW29AcJ2kRdN/vHdAHWKNd1Sryoo8MyM
dje211J+G7vPINPFjNzBUcsIVQruUGoGp5JHTpG6+cyXfAeeFc+v2mH1+H+l
HuM+zZIggseWBje64v5iaxcCcgZJ0e7QyM3huxp1qbeBsFsLTuPrQYnMMYBH
izMsPHpnXZN2LrsA+m/8982lzmHESfkMuNz5DUsodUZT9kHUEXu3Z3N2LZ9g
tAEQEaUkypeSty8zaVYySRdnvJ05HFtejNqm5GNjKQtyiGtVi2RIaxLkr5in
cyjL4BQE0hOpKarvw58znGnU0M4x618dWYVQfkUQ1Cbp0rSuhDUrmGQ1L0wM
J1F+wBW/Sqt7YmZReJQ37LG18p0kYrnfvEZ9rEdiPQmGUd3XmAPUBpMSVWmU
u/pkmNL1ZW6vux66YAmNgk7Yh8XyR453PgUqUxpw/3w3vYh3rueSBaHFb0d7
TJawGERmHE6wCMqjKRMzf+PMRfiSmAvHPYnVffrgi3IlR5p583rDlaTzC056
iB264XKNzTf5xv3FtYbeZu3tdCJvnMGiyYkayUYxhkq5ho8c5X+tH85WhXYH
U8HCQrKIZrf84TVe8pxFiDEC/4kJ9K7XubYnxIwdD1xmmkZakangvJ935thK
uVdYGzDH2C4d0Mq2wv1/WIMkLzMuFUG+Kkf/qFjPuoSPFC7RraM+O2i3nr1F
GeaKo3N23sFvnlQXOKJr7OjgMejPoPYid7Q8tLCXIIyvpIh6wlx30T1CYnVN
U5yzg1V1CJbmwChv9RD1VD1K0nb7MW6dKMjarwA5kcpqRj++dPncaa83IuiJ
7DKU/wDkpImJMpBnQWuFaf62swqfMlO63XNzhP8yuD10bJp2bjSuObBnfWeW
jmCC4A+6iZNId+nVurEgWl3sYvudz1b2fzmNT81DHG9M5MseqHxYAyLft5fz
3FdaaQdGSXH5uyZnrTr2+tlJNQlSZxl66RdJrdWc0oftfEyLyA4EpnN062eJ
4arYgE8mqM5UlDz2jvO+SE07vAkU5tRnHwq5aEKHDtjtATAIRrNTA3+jeUxf
F3t/69hJDv/RrhBasKug5FNZf9siRuB3nQkiOvDPnNw10Cc9+mEIK51hTISZ
JC65j26uGwO3ldjHlldeCBc/VmKClqgO/lOyBkzza47G48luQqzgyHT/lwH/
46Qb5if/wjgQC28hmL3ZqpIoUnTi6gmwwJkQ04P15WaVmEag6P8CPiNggmzJ
Wi+UfvZk9WE14NxwVOovM5d3VUQN9HJNG0Kjhf8s7RViGq/eDpbn9FtN9vVs
GJD4pxSVbP8dU9FHWA1FoNyFnpXyD24DUHmGyheZbKOfYOrOHIT4iWLPXion
/2nfDD8W5mA4159o6ilCThhshG3R428hI4R590tmZ/qLk51c+UciFpjFHoQS
KFSWYSiSulriibX6VEQ2RWL+fO+frQ9P/r1loQhHCfy4lw1W7NU9wRhIpk9C
zCuJEJ+rQEcHjm6ZxLcqj+jHNPkFvWjQSjOXwnEIuIOT8xkJImqcXb0MuEiY
4AFNNdJgBs8OR67tSMl1JAPe/Higt7YP6CqJ0c6uJZdZQr7nQRgn1Htc8U3W
omjQIkUtufWkyCFDaDI+uOuAa0LwpvRyY754OzOtEt9WD78MsBBpAsM91ONA
v3sjJXNb76jOxGAh5CnR6+HSMeLn4wj3ntKoD9ea0e7M1fIuPTiOnRIIfqwN
swcZj7eTIUPApDTKzLdffuuV1A4GoZcnwCcEzBCCpWC7rjxmWv+jlRyrz0WM
KwZE3CV71qbbvpisvTZrAT/4SbjPG/RvcBYoXe5LXhzMo0Cl/9g1QfS9A4El
qvecGiwskJ95flaFg3QfKtRQBmAc+v0zM9LYlAmoJubrAElbMUg2vGGVtoAz
Hk9tlxeKHK1cjBrqeapzvWd21+Ig8nWgXBoj4mTtDJctonutQZVHYWrNCaGQ
JNbdgQo/Oph6hK9TsNVC4fDj8uS+UtFltQuune0nPBIl0pt/o8wZbbTsC3I5
WlU1wxtY/SWGJqDzmPEl68oOXhiZ7wtpmKaGIXziPS2cbbJtfd2qSaqR5P8A
6xm5oz2LuGj7NdfXV1iWaaJBxjUelep3IyOlEZ2J5Am4hYSHfjN20v/pRuLE
fvJr2LzyEXfAbpPu7QuFJk7xt7sjDohwnMpCCdwHKcvPqFKcw1T3c/O2XchW
8sDfhqlH3WZhMz+AAWxo796BkJez9AYfXXmD0VbRUGRjWFqtoGaSjisMQ/lU
ub1hKx/hzrEj4RqjGYdJ8sQW72wSves99MqU9vPdPQWM4kDvzm418JPjArcE
HDNeGCDZ37XPCrIxsDSerL0fT2Dh8nxXKyODG1/gM0y6r+m5Mf5YiLyn7VS/
ByZKszkZGn5YGI6d58aQW+6frZj6Z/yist2YagWvcekC4+l/oF9oqvS+EK0z
j/+Y4LsCyG4JQgrpJTH0rz6vkwxcAmlHDyKWQSoXu7Tk4cHA0T0F+0JS6MBX
VbD9kG8ovoTeX5vFZtgMZ3Nk8DHMZZiMFLXr2QRwHWeYwjl0Z6rIq/GxVsah
FXxd0X0Ph4p1faJooSyi7DIGRfH2YSSdzXVCVIll3tVq9buY22i+axKGfaxr
WDBcPj+6trVsd9RcrWrt2W4LcRXsjkuHnCrpgs0IDPAaaPFELCVy6+nShcZE
nZhPi1h98rscFvNeQyE2N6OZmGTv4QKPwwoWql8WPZN3a5Kbse0R86cUq0Ud
IBoVWcC7SDAN8+4GRwE0e8lpvW5dtcZuQXXnj9oldwHXOzsSeB2/cjtY20T0
Fv3b1Dd8+9Q5F5VAqOQwRszWWGDY0gJQIRgivpnj4oPmHAgF7SJvZGjq7H+L
p6KtrQ7xBnLiuktjXCqi5MLepEOIZ/8a3dKo5MiVA9U1GPYdFxZwH0+0pn1w
ZeK/APEPNUhbuSYkwpbnQTKB5YUj+3/MA7HGzSNtag0n3hr6PcISiXvcLaqU
TH9Qyl+rxZl1a8aFs0BKuEgvOVYnXebIzp5bit2HVXEDmVsLtOYa7bdA5auk
b5v6yaIwmQGz9Dy+cnbOQN58G4P18R1RihcbRw0MFITkgoX71/M8lA4a+6WT
XBYx1GjZJ9PaVfFuSQKBGx/C4GUMHyXH9uttara4mWzgRew9JvepSZpNrf01
bQMdUvzEZMOdQ063WQHjzvgm07N7nvm0U4zFDk0/694j65HD03UHoLO+JQr/
jT2uU+7Z5BE4yZopR2aM4Au7L44PChQHU33iQBISXwDBIKwrfzAtRQtR8Frv
Nz/o1Ym3JTprieX1vA2LZJPm023B6u/Oh9lviOaNz0n9tLPgns9gdqRJqMU6
lRqX2QOpRtkB0GANVqXXtyjecvte+zFiLCCTThTtUSaBgMtLwezTCa0E5QFJ
dOvyMS5hzXbgl+TlBwodvLmNoGNrfQsMESbn2tQlIkorJ0tFgkjBB6tdl6VP
47D/i+Ore6qtqKXCwLSH/6A31DG8r+ZQebyrFanhhQvodm6U4fKbc2O9z2ld
zafMwKNKSuGNE7VI6sDqqN0AxBCwJFwU2q3IEpgK6oMIme4hmm4E/iGNnNUF
QPkNqCGOg0JKSXocKc7+6rVgQVOfQcv7Dc9HuRahjSHncA7TKF5EqDzWFliu
yltp4/z2TlJoilGqgU/N1EvC4tth3v5wegCFnAZH0v8oZI4JuqWnSP/jZ8Iv
SfZUh956abFwgS7AZn7ZxOmtGBtut7Mmr67vE0lCWV3Pc2wpBTuKIBU4josV
KeD3GChh8uI4Rm4txQiC7WZA3Nq7QwTd2zGneAxTExpwQNUU02MZCgrKgMT5
FJ7yAHzh+freoInwfmCYfz2fXNrd8kauXE0ynsf1HPM6E6D/u9RF5tm6h9Ra
H8/n/Wd7WBDiEbp/fvBdMikzL2d8MQQ5oOnX3uE9VwDXvnomR5c35HUFWJq7
xv34ygLkBjzynPfhch/okTNvV4fjCjds7sPfA8B4u8WRstvo38KR1lVYdP/r
K1cySTbRe9qsHR71dmKgN4Edr6wGojXjeYWCHs5iBkf99BIECaJQgAifthlj
TQnLfPkxL81dS4LXF1dRpToJz0tTLQhtzSgJTqFbXD5YVaPc3Um1X3vpLVBe
jt/XKXYH2/YPIbn6IK/SwSja6Jkq9oe1cagoJGp3Z6XldE/1fnEtkg3DGY9/
ploxcw3NlGTqUn04+TZQKGGOjaMiLyKAozP/vaBVAYaJxdKdknxoFUMdJEBD
NgJzCkBEMxt040QWgvFJ2XTVSKIGsszv8NE3R/oG2RiANI+yksPDy+brMzUg
P92Mt9EpqFHFQSjv9sxZtsEc+I1XIzR+w5YL73KGBwRlcaDgVirCTIIe8Gcx
437ArEDBGpdbcY3SDhid/PRs0EFC35gmw0rNBuoXzBICzPQ+7Fj2oubhTkkM
pgFsXET9MQOzBNUGL4UZ5q/bDSvLi2t2rDc3nXySLig5krHPnvCVirLAEsUG
WIE2Vq91gFGeMcFOGOKvtNvwlb5ZuwqJuS7L71fFVgCA6ek2bxlKArTDKQDW
PUt8Ja1MNGD98YbwitqMDYaZkStSlsE8WWOAQFqaVNF1grMabg6LyJ+Z62Y1
TaBswuE6CKLVBN63GfP9epG8tuvJAWcu+yvM+5TmLBA2bfGDsC3GZbEe9P71
SIxvR329ajNV0quE9QoJQ1+fKLnwq78+ZrADLoyZiGul8lcEZg8KfvEtG53v
PD6mTVzPO2NRbg4mw4/Aoh53YHS1ojPEBOducKRAshbp+ys4/JCP9d6+NKmT
rqiOeXYfSxS1QMKbMLKfa7E2gR+D/C9qtRFTIz+qvZ8wKx5Xop85grNAWLJd
MWywwH/pk44tIFnEUvGM13BWFttz9fGFp2r1TJKPWA6AJ24Vt1s3r5GXhVYr
QrIZbssHZHaeeBYKchmdy20UKzvSE7kGFr7y1er320W5GlGgcnyANNA8ZYZm
4k+ZiAziGpkfQAutpGmWceEi1jd/8vEcxuCeZUOMelzUwWQOAuN5BzmJtW3C
mVAhVcgbzrAY44KY80TYGIHq6T9cJnM5+10Q32qL6WAgvuW/ZVvOlzGfzfhu
lDXBhAUDwHmUqk3lcM+ziC6Ue1uw3RNpeE7jArnyJg+MSxuE4AApon4/ESWl
TUjZ1tZ5B7a4mSstH5JxRMmzB6hDdA533zKIcNl22qQ5OYrGvRmnnzVgGymd
pxvqumk12LuspDVYzbxA4LmkY97pzvnzFO6xVaoNMDMt5FyqNM2PI1tNWGU6
bLsjHJ4oRbH6C8nDVmVOz0WJufy6rp7z9szxDOt3l9Yy0kivP5ToL6c5s4o6
seLkohgqKNZhhPUQ25sBPBhVx/ewHvh2NH1cTAvBs8YIL6Q5533Dfu3D0z1o
biqdQB9GSVvpuSEdDZtGpxhWjt1iH/vC8TntAxjl+3GzQ+pPFUtJ8HbD126f
fRt8IRNp4GzFjv51jwaBCZcxQyXoNozr8iiwn9lkejOKWkklW2o6FhNFLKgR
rVdOT30RGMlOQaa1pqcNB8QSHrg/1LRU1g6qHo6SwHc0aNqE3yKxgA1szD4b
imgxI5HMtZ7jrmmcKumBBQjWDk4f4zHd3X/4Y9y7UtPSRkX8bcoL19ozU3Wb
7u+3+ywtaBzjzvkG1c1uZIiCuhUHWoS6RwSxeSpbRwATMurr+QZ/FM2opGcK
HZ/1dcy5m9yw/+om5JP/K5WT/pxXDm8T90WxT0Sh7TfTo4a+Bm9sxuPJBaDH
ZvdWiMUtpzXXvUVUojhOJ5y2WJg8LlNe4knwBA1boNFmigond9R3D1oKMFpo
W1ynBch7dcyiZbtiyVazxrFBfN8NJGABwf7UERTXZZ6cmI0ozXrx0X9aBoTE
hTni38rlGzONYKeqTpK8NFX93HVbtohHUweMJ9W8JI6pQuymVZl5ZW5RcdWa
GSMh1HZwE2Gs/poR4mLcqBoGKZFxRN7zV1vDfbBgP/5rnFIbqa6UdUaDUs9D
50swXRjZwu5x/ta0QbZYZ+GV2/Zzyfdu3b3hIrXViWsTZsO7Bt/O77Uqkfue
1HEPf1VE3BZW8cdLEqa4Xu3RgzbzXtwcMBQi5f3NpNbwNEdAm2C86oCyGV0z
uhmIhqCy1WjGMoKynb+0cjOZhfBDjCIpHOoNcIC36K+nl+10A8TFrwLwqwRD
HaeQBGDc8WDHDYraKefAtay6J9+Fyh+WKdsJRbpZgrmVXmBCo3x1MKWQlnuD
rVX6ABJ5mqFvuTl7kJmrGinaL1rXEfySAfeswiyn4+hUYNPC0NDQZuhDfPPF
mrna0NoXfS9CCQ5qMV/JeBFlBkhF4hcQLY6+VuX3veJp3rjleyGxu4UFKxwO
Qx73cuSdXX3WUH58dMQ3iNUmmMFJT9PNDAZIu8qejrG5whaEgj8QWV82EvUb
XHmEVI+hjy9hReBu+4OOYlIH6VQsaAOBTdBx2QLbSnNTRGhuaRJwPadRk34l
3rLcbvObjPai6FLYXZyv1N+DCeTrtqkh9IJhFYlp9anJtJk+bnYZrc3ClhEi
jHcw42SAHA3T7rozK6mBvXuy9jQR8zyZVvY6sdBVhe57/1Fa9AaoCXASKQ4h
4v2+H1PdwjGMibMJUrg+dULJP2f1xj+xKgvIbOi4PNLTZc1YljTpBL0ruwfW
Fex4V0doR3/IvsJ8PemVXOE4BDSlEE6TuIzPDrE8tYs8Nx6LCd2QXT5n8622
PJetgUpH6JZkalPKp6L5IKNXuwe3HLxMboQK+SpWjbaIzvowsHYdvKzv5S5K
W394FUFQe7r42J9ZU1d4vVJybHvQQCXOShjBTEUzo3Vl8qb/i/wKKyQhi9mX
lAZHAV8+/3y+ewsSQl/tYxL7mU+FkZUfaK7LHWgnlhCf2e295I38P9VDu2Cl
3WZJrkQ3kdWvQsiprsY5IjDjk/qAdlnzQWC2YKVBi7QjnJSBekyWsjeEIP9V
/U7JVV0jaLeyY4DlllbVNKpyDFYal2sCFohM1wEsofZ+6lbKJWKFOzTRybri
2hfZZ29oOWeQk0K/6ZU+Qqew0SjjTBHsfo5CFYmgBrrhvHif7LmH2zWCJXQ0
ugyCzYDR+sPZPqPO/UGLt5lpddZTQitSbcSOKTJO4jzCG5ANqLmZThCTtv6H
IW8ZslYLH6W3qMauJRvYGHMnFJlj6jgwI/WzErpz2DGar4E1HPOxbIPVBbTg
peADGttjJsP1s6kxKqUlEQq/SuP97YWEvsgXI78MakBREK5y06GjdnKXTDh8
zl4REAQvKBqfoyTMfEnePn0qe4z35hcKykrv4gkwNy++8s5sqghn971R//ka
rD4eIdOeg6Jd+CdNcIsGMX8PImwbD53LUw/Po+x6ovQjPnTZnbBxhDotvK4v
LByONZ1EFnmTIJ+/kIzAUaYkNTMPMa3ZJEPVqd0NMGAiJDI/CjuExvL8sJW3
gt8/5OlBP4ASepbq9zfQrEaKmgE9wA8IEuTXd4MddiPyaUjF7QfSz/1Lkf4n
YyzhGQAxGgQC8Ej0GsiwWIXNxj5S5HtF6k3U65YGFY8OICNZDL7cRPo4yoEX
d8AVJQEE6W6Gvn3UpaaIgp9+zose8rNAmR8T4dMqyplovuXxr/dGhBOEjl7x
NQcwxkJXz2FtWRSbw/AvuQ66Lq9OE962rdiTRZ69ZdBNMs3ac8sujpTUyTEC
qCDEELgNZmNGUlVDETkl3VDK2aYfVlVzUbvnz5rEEJJR/gxX8n+nzht5tMJh
FyO04XtBApMYQCXtuuKs9KApDxvamPDKrQmlDJFjI802Pl6un4otzNOzUUTp
QoBkW4fHCYhZhHA2d7Z5xq5FfgqQCgwqipDftsngMYyjgZkO1OIducCnQsgw
g9YzaI2kfNiyZSKp4946+zoXXrSKYQDApxYEmbz8P/MI2C5gUm622QUUnK7s
tW+vfiq6/3DqG3xa+M5wJk1BogtnqMo12OCfGZRi6i0ukmnok7XVfweOEerH
w1mAlaPFmnTcFHYhsLxvlKZ/vPvl9uFi2aP55PWApvgMjw6aerwFIWe65SsH
VdKuXEp1IrGYaNxO8aVX0GLIn6PkCy69S/Nfg0Zh408bMf3N2rGlYxKfNLAz
rydL7xhfwFcCwZ+TyZEPzlN4G2Grra+LzGmWnvXe/3e7PXGJqU4amBfilz0T
5Xc0zcz7NeaXQ+ofuLYE19lNTTXTI0hqSWCh2w9erIvPhMwMWLnrTnjsZleJ
pJ1Ob2satdtu0eqLEzJ8CLAn7y7Y9kKiwp22prDROR/G3tBD+RGpIhwka/pm
FSTijkJzzT+XXP7Zj7rgsUlMyOLUbhgt1k2SN5rXwATuV42A6+sKFwHkTqcb
uOeumQMz9BKrGPBgfLqa0/mUgN2Zw9DsH2Q7DYUwijIVpw1b003QOGYzQLuu
ruH8v4soTJ643qIjuaV3/SwSsMbDy+ETJddlLHVtl2INo+ub8oTkIpgwraHD
PU10jhONuEFyspXq6yY4SP4PGVF5xBDlfKh6/aUdmaFhzsu0uwn6Ai/HTSHj
B52rEvMeyO2poFOXPPIXuzsp98Ai3vBaLzqI3fVWGqnojxecAZF1AeIAo7Oy
eSIhHHy//iGZm4JB2B5PD+U5YVhSADd72DPRUElCGD6/VtVUk95Bf/sK+ULn
hv/PAZB022BtNyWcaGavO2yGe+WzuxGpUM/ZZF+E6fjL0WZ0gzj7W2OSk5bT
cQjMZLz50yv+ZBsivyP8LivnU2hw/Gv5/ni1sfKwtRT3S3IF5iLZDBlnC/G1
8njNYTNG9ZMOsRYhth+Vb5Uealf2g0VPbSO+mJV+H6FcygPEKDIxBUI7jWYv
I22DdNwKldb7QFeqEMoxzgAyqx/r2gxsFH/WvsamDHxMu8U0YB28fujGTHmo
jFkuUmwuM6uYaExJyRABJ+zAlD0w5z9mQT3BCY1pnEsZ7kFB3IyOas+lcvHh
T8dMXec289znUnX7MZC31vo+y6cmK3jXzje1JOM8Pdyvv1tAaDgV+ubQcwjb
T6OWe1XN+kScvrEXjCxYAhzC7T9v8MhbPW30rAs2GjpXE5l/GMzzNbDsuXBy
8D1Ex7wPzH6h2NjdenRgBBop+Oug+MW2g7npzdaU/p+QdA5OFSFWbCw8/pB1
Yt8+hOiGQ/FoNIgpdyMLWQBmPjllMTM7wodm3ZfCDzdojZACwqkcr59CGjga
0ZItys0YGnLNNaLQZB7bTm3AS9sAoLYnWZAeqRf6ox3qkQEi2NbqFyt64QRF
yQTgQ0Y13JQ2083ahNYsni+NdlOjIL8srLByKMVpICfgO/U96fskFzISgHlX
KpZM2heuPPYhErcoT7Uzen942lmPKNeCqzfPQSSPJTDkiKtH5NnGN7V9ewuC
DyOBnnEUO0V2ZodnbAMglwnMu/hjpX8eoqsxBmugtijrnsIa51823izLqX2d
VjVh3yiQ2Np7xUiaRgPsDu9Ax4/nnNQGzDDo1JgyUqYm+qsHH7FfGVvG6v+9
71Z3qaAESabjcBRnHrKoNB8rxCYiAS7z/sW5AWUYvkaSpFgL67jOtnfQ7vRv
WCBKA18Mf1JcckEzeAi7wEf2j+tslO0vQ29FUeGi6UMjVluUiCBA/0hPTLZh
2yLXk2moWvbcSH3LExr1AxUdCH9to3GSrb04hw4Shgg8F4imq1R603JQQClb
qd4yOr2Sci+zzQh4JMNUhL2kNcR8V8EdLLxPZd3ygUImc3LHSX8xZwlY0V4Q
BsSJ9cdoguyC7xoGJSb9IGKun/xmjxsYU7xQ6F2FBPpn3WYKkB4l3yf9N+Gi
pYRv3gMaQ9grDAAAg28dspIKqXbdAoAEcOVsfV7nZCT73zvh6PtymXSQ9Hnw
dXPpxu4eWp6StzBNK46aeuxk36sgjdSwCMRhMzL1Ht/+bxrN+aJ65IOcSnTT
HuN+X+c2Uv7qMaSPx+4s/NWLmQZtZo9Ly0MIpJGdITDeRayu/njSweDbrrC4
Z+VaMNggkAKQD2+7TzAtWZ/Uhg5hs5A3AWXFN6KqpQsFH429fZkwL6Qu4Boy
wnlYRK1Sm1huQs94MaKK9SAPjk/EgJ3h3dw0jHMcYximrDevdKPHDl+odW/A
kLP67eBwzGrFxIjlx73JGSMrLlyktaDoS0ZPcPuZ85wS/sY4UphfK0v4YHsj
AuqU51UhXSzXet1RkN99CmxCMPHtNsSG3p8Eda6vTo2d1YPiGeZLDFxRSs5z
ALQcGEFq7AasSMRn1UcCwFy3KzFw8UXNwLhSnHq5/8KmnF6RYrj926ScQGIo
tLpxEoqGJFXrbJZemCaJr3jjqsQ+5kT0xuJI0uVr0JaI8X7h+qJOXyBA+MUH
0/ffzcHAra4mSahfGhKRPxNUqT1DlFJSOOSYBGro+hR5JEK9Ht4Nx2MJ3uS+
n7T+dFiXpxJi0LPqBsu1el3Qdbono2w9bhkDf9XK+yaKHXQsXjGV1L041WJl
E0teRN2K/gSlvrQBacSfetcecpFlXjuVg/KhDIyNzMfFq+Tel2LUukjnz6An
dCCMzJlQmybBRACjJDThLO2fZ2+CNc98hsJ61DSbfSShHRoWxpCL5HzAK0Yz
18RP6rLKBIiaO6lE3iBWOXE2EE0DHUfAqLeSH3qHYEvCTBcnXu+7k8gLrUw0
Th9cyXQVhuQO4rB2LrW+9UmcIPqaPzpBoaPIZqaQoI93mf2bB5PrmKBgbieW
8iJ7OtUu2BqPKDzIa/abaHjLXl3ncmIF3I+5q2ybKk+45hwX0r+iBMUYaTjW
9PWW09MILf+mSMFz5k908HCc5XgOErUhBs876kNLO+e/xfug9dsnmnGaijJp
35Q4pb2ZF4NemZxVp1TtkUqmRFurJ6mppUHJ7aNn2pHLooYuPN4E/W/OekjC
HmgB2brPN9an1qV8OVILfzu71xgFSeYSsVMtKm9/ZqYm3m+BfPsHeLsbKJjX
edqFsSF2KNrTM1jVSywifSozVKyyyuTzcjeVKG17Q6ndcp0690twIMSiWSgl
7VQ2SVyh7RqxNq27OqkxUQ2LjI9bVk6WzxpReXxKgb1ImiNycDId6Jq82eS0
FPqpI5xRMDRLAXsYfbLBgoCbRTXL9tNj6JMPLbaoQYXtryd+byvhJQaqGeMe
wGUh3npBgMg+tNgKuol+4mZO0Vz9ZdaWbfVxSdUkuK1tFxaTy/Mso5Y9bG4m
9M8ZvfVMeShqsT3jW6fPn1oIAdw5vqxpt5HFZJWSS2q06OW27iOsrqku2ap5
a2uBn7ZolxSpHPsHA7i2GWZex4XRJCePuXkDVBigQrlZMwkUnHO0NElZzGpd
UigrcutZyU3XFB9a3Rzne9WrYORJvkHKLyRiMlQis2euKU6eK2Yck+Bag3C3
8JhkfFc7Yskjy0f1zalm2Ofu289/wR79UA45XYs/O92am9+exDqBIQSN4JKf
YniIJqwBIS+5zxmAbot0W8G3Eeoiv3mvqmK+OUcfQvykDuTg5qLMaU5XTwPi
WG19u4DmuYNBhIYFWeRThy5xunRZ8rvONVqJ47zIMbw0h+5EapmH50AINdtx
YnPYkzlb5WhdoerK5YErs+t3QS10+CBkS2U9UyCFwybQwsZ0FB4RoQ3jyR1r
yyhlkagrAiddoeAWYhB8FhY0t7mo3wGLLNLl++NH9+8iCPTFeCNYthw7b9Wj
F3qwPD8ZuT4ZxlQXBfdVDDfRLfTn3YGFpz3WzjmTCwJySaDOupD6TCmKZN29
e6gpSey39rUpmbdnqtb/6V7UzbnxWAx+CdlDsa0NDsA6PrcOQUN/1ozupx5s
gw/49GkwfTliBOLPCdiZOueLotRN1s0wBWLi74GSzemvuBrtUc6+upSHfk2n
n4mSFDYBTNDOgWmMPke8D2GyXLEv9gaQ/SZJDKOyAlCoqspH/bttPdfrFZCR
67AFTeSbyvJNVcMKkhhVfd//IH1ZwzRCrJUbm+cLGQTWBj7gYGFVfi4Hp6XA
l4ckhSA4EfD/qOW7T2nMyccWENaTYsD8x+ttci2H3JiJ+pfGsodrXNFGIxx0
P0/+iPYFfINGziPiwB7dRbCsBHAqKL5XmJXBkKYdOa4rxoHFTRbZn7+azhYy
2vfAyMkx3LSZUQpvNqZ5vAqjBgGHiJdhmPQzxOVmno2edTez8bH5rwXPaPxn
yWJcn5PGuPKIEPG0eV5NwgMh0fDhqUtKEIwKBpVYY5x7UdlJUVK77foRUHrc
IuGGUJMU1Uc+b2D03zi+08mOVbQcrMElOz3RFmdalvJ0Jytm8yQE298b7Z2Z
hYyKgB1azj97DdPaYWGwegV48ufReX6n3WMGO1chQKOCJuYVqBwdnPYSbDzA
kRlmUORovbI4/X9TsIgKd6efh8JV7MehFDyCaQ589+aIOCMv+4T8k2cKM5rm
wHA9tcU6S/Dg0HnUsLS8vhbFqbWriN+O2OJWUmKua5XxwqSXBFWa2ylPj2cT
c0pPJTmT+EE4N8m9+ZruYRoNeG0pDgcPhXALy5VmE8rvlwRm6fmPQcccNXjD
f7eYWyxhIL5UmR9uT1vPwf51BZei8eFBkOvas+riMRZw/jOfsZvEAs4QnmFo
5mrnZpwp1m7UTyg6FDupAhIM9gwtFxH0rKrQ6geAl7y8JZ5wbzersRiR201F
EVRIYEQ61ATy4P+an9PguwSEoC2d8g4Ahb28UyEkqculIlO/ttJx1cyBA5CU
Q9UYqLkUZIBzEgqFZISvp8Ol4jxXVh2RuiRGXjhHU1EaycPxqCSw3p4z26eH
VLHb5N3BpSz9ifnYpgURu7R1xWeMv+v7y8NDzyllsggDin2woC9TGB6N9JPn
WgjVLHVfI2Ccvm9/v/gs90XbGqIuOSurYoCtunKkABfxfM0bPG5R4vNjIn+z
iEaFX+FJy9vrrF7CPpxkl4zO/iqXZji71XGNXPFk8DjlcfJBi8ulHZIh/D7C
FBVag4TQraCSY+9pnBupW+hCA9rLUbszUrbk/AWkpYDTIX9eDCz2oQCbA7PD
Bg2a2oMKHAJ4Z6msRkviK/9XYsXOi9wqek1m7FwoteUYKuJsMCukfzMqaSfs
izICcnDveZ9uwNVKscZ/qDB2+91jlHb2T6j6ppRdrLqgZpBGw8sM0iaCfZSW
C8YMsy6GlC9lKWufAEdmPztRk5l8iE74wq9j2SzaZqA0WlCFJVKrIX+k25ik
i6/ZcauB3loRglHQtmpXbM0iudx/rO3XyUUGHA8q5zts09HujeQLJf/jyENU
ZBJVJUucjOcj/0mWIsRj5p/iuNw5kmjh585VVMuHus5sn4xIhXgalKw6MGqN
JUrmi8ITHGc98e6+kbLGnuVA6BHcFwCJYOeIpDpPSlFJDGZk4sLLbCnStlWu
n6CB01N9sWirYVgeGx7Pi6wwHwQTfqWjltPTVMvMBLPmMJBGDKTs5e+cnu+F
V3qUUsMK1DGUVo0/ePABJwTA1LIg9AzWl9I10RzjvdcOS0OSZJQTgpUyisE+
2f99xahHg6O7sa2WzOHYvOui5ir84akkBRoSrCCb54nRPmQj3OgP0Sxf8kn3
22OCKyj5T6gkuILIfDssMZ7w9MtxelT1uu2OUXCwhFzHltgJeBuPD99oS41i
m00C9ffqVtmXXkdWj4TG60Cyk0T2ePVeB1pvOmpFlvVdty4g5VvAjuC6fKNu
tFWHDeUfNRhtAdGSxH/c0Iendx+Jqf1S8UNQxf8F0y014RecW9pLg9G75gDh
AeXaw5SF6WfgxREgOnlrmsHBOElBz1FT6HNFPMuiVhuSICfv5A9W3kGB07Pw
hWp12eSztHzmI7mQ87q9+DBlXvV3kM8Qp1J7p6/xOvodnvO0ekCL3wh+y9Ly
SXZgjO04FaAG8m4oba4JGc32qvjYRk3jymMBOQovs01URi4rfj8SCI1GclyZ
rD3K0lcVAKxO6kxZPHdIDJ/u4DXKBLPylSW0H05fDVCX90oHGzUOQuFOOcMI
8WcmqpZprvCyA4tn4JqAZzKhB19ImDOOOeUKseBnnhRDkOKlsQ/Gnpk1ki8s
qW3iSqGo5Oc23l1Q3xWzIxz+NMraBRyB/k5rQBoJTyaJVq05bNr5fd/ofS/m
vVlaL3Ax/IwdZgJi8X75cJG/6qkC/1X1pSyUiSpYE0DCp4PJsSxhW6vNS7lj
9Tt7up/ImOqbxX0BOSB+e7VI780FX+cWHUTBbYgTKSwXKLPVWgtYZhyHputG
jlMJNyLxoDVKVS42lIWMoFGZ7kXjRGN7Om51jx7RwB0IFOvDP+8ru9S3/h42
yx8W0Hs6g0+TQ+ntjkk1f/vzCMBPRCY/dYpJwJk0npaYoFJZZ3AimICdDXZC
guKb2KqA1JYl1nzpqXANGWvR9fGe0f2aG3oMMKURYL71qEbg/RK2k0WyvwPz
W2l3wm0PFf94ulnJpn9IOUD7pSM4yP0wx8030TkHuAveUE0/52uJFTXHS64R
xtSPmS+uSgINUbIWSzgRxESkHf1KW2dV4lVGoynauttlugbKRr7NGf9QwY9A
8rmRWKcCq9I0S9SxZLjkI2pe+y2Rj3ESjsVbsAPyvWQASjSbTWP6BX6cRvKS
GHfO+XI5NLr/6gGRFJFtMIanR6FZa+Bxwht+0Ty4gJpBFN6Ps/bZ4PINDhWw
ULMt5+mUXiBUYcHcqR9iUTkavnuDHh8nOxY/z9I/lqCUJGOcO9j167C6OkN/
MNByZ+F4bUYuDzWER9EX0L4/cJaGs9uhC8OCL+1fCGRFXhyGKsWj0hvVjlU/
ne9N9Pxl+bfiTGUuVr+zF9yc131ZD28dZsB/d6sbfB37yBgmpiOR072WIT+z
Y6bS4/tEt6J9xGsh+mgUrXndWTV6yFHEU5qaG5rFcydcdtDIPN/cbys6SbIX
tuXZMXcqXm21xKCwijrj5CZVou6Bvaeo2oIL031I5PyEgku7P7NJ0YDNj/OM
M5JqthvFnjN6yVjedcD8QaGERhHb1Js3QyypuC3zYqdJrgJMv2uyIFksdgtC
A5cUdtgnKvp9qHtEn4CqnLwTJ/gGz+xuJenhfzP70wjsy4KfgLVctV+IBxJK
sIUsofRkGA8OFYUny2zfA7n8keT6e4qwPvbOiyVmxXC3iCX0zSykg7LXrsR+
EcTVhncZ/ejEpERE739ZrqZQIpXtG+dIv3YHM6Ojy4Sv2YrhDK0vRgJv6tlg
Yg2PKcsUSBDP9uR6tM0D4LVkVn7rQiTYLHALGHLKaeJ3miYvoSjUdkNR6v07
puO4HZqq3A3ucx8G9FuwOR/PDZIDkThZTt8iZSKYLRgqa879Yh4RKuPWnlgH
7l+6mtwQyB+aDE4g4lRqnc1Fs26JWlHJyg8BMeT9Di1DFM/nE6hyIXRn9Qva
LRVRwNydiHHU4rcUM0Z8h0Lf2ClYJh6go7YF9LCowOyCjGgy7tNWBkTo3+fR
0FAmAMsxcighB7j8SB2ZpBmC2Pz+6EdooAwlpI0OoYrGu+FQrpRBaJaqdOob
PMyGmJqC4F5zfEZWTu2L9TKOGzDaY40LqsFtdsxC6pogDc4mS0z6yG3JniWm
EruyEkqFLfE8xaDZCZGo0+IDQpPl6xInFtHtOaFOblN9Kp+bT8/fnMOXNPRx
DuuWSSTQDv/lbFBtck9+sm5GBlN9K/0oFx9rEhlXKtRFb0rerNgHZnSeA8sn
6sjAVf+gol4+im6YNQSfd8ZnXq5JgnoDF3b2rDJE9Tm8VKzte6fKD1PLHEMo
D34m1MIqLwLMAd70z3od3zbaoiqLlH5a7PkWTEFq7jukaCvaieWuMTOLbIB7
B//RSq46dynbHRMEu6Xt3+kLv/mP64mnYI8IfVo9E+uKe61QXTdzmRtVN8sx
8tPzPI6vabxdx8x/R0WAVR2vdU03Mk2mb31e+o0CDQkAGvprtlPmS+C5xvaU
JxuT7R48GGvZ5+npFoAErFJCUi0m/G30fVIvmXiVrMNXY66Rn7Zvz5XlXmHb
qdGBQM0KrQ7nWG3TI7yQbNR6z/uBbblJm75uKFTA2uCHmbcvsAvdbf+HhmJc
B9lQ++v1ng7FZk14SxwYZ6+wnofIQPgyLapuvcPeihThoeZoU3lGxRkUi3BY
apzaAyoc3QF736qtq62bfNVK+ok3irlgpdOwT7NKEi7xy1WsSN6oaINSqtaP
lvmrfiyTXEQC8fxnh+yFPTcTfr/HW8Rzd6db7rKrV9AMSIHvxF+//EMdqiqa
eAdt4gcRr6waEQhJJZlYEmEtoFDugAtWhxYqGhAHX58tR7o9w6BWmfwoWO6y
ndNw+LzS2Hlzg8tJeyEGhI8vpq7uG7PYK/QzDTtQh1eVK8nEFZhBZhB3P5et
SllLkWb5rk8DrGufK8lPWBpq3SPY78FNsbDyxIqle0WR82uVBFMBkJjCf68C
pKJIjPa1A32yHWMC+pG05Pu+NW9z0ZS1ASIQTRZfxm27i5Q2yN1rnW32fXc8
bdfAx0GWQkGHe85FhHqxUAHHITOQXfGi95Tok8BoTGIkfJmkZLyQrAQYO+Ne
tnOhBUlV+26T2Gew7jPcJdm5YVbF8+CQNrwhlwXYq28hmf9Vkt2htyNHwfXm
A/3mKJ74TpesOdbbbdTF03zMVmoYtQjb1uljt9kC2KuqRWSbkoaEkH8xa4Qq
XGu/thsl9jFeKGwcwtSnDW/cvjKw6dP18i1tsFGEmSQ+OnFZtQmv1RZXWmab
aEsHx553b2+8tGOecgZN/VDL3r2scATj7490cuqbXyAkIcPDqmdeXDk3JqM6
EXaHPqtsSM+86XrYINycOgOKSbuf1xODMeT+ukcICsgMNirK3R5iabMRMrAK
NvTHnxtNqfisfglOrT59ILKAQdUEzVOyDmK0HsOThAPaREONJPKjYeU4+PAp
Q/syIT8bFUa+UOTxdfZ9qdsypKLUstj7V0kXQpWOPa1+Abb472Z9Rnnfvl0o
u5fWFc5hbykz1+FFLPPw8AtDOLYVxsbmbg82klfGyXPxNxIUkMnRp6H+r1E2
Z0AUlHQ6T5vwCW+lspzmgL20d4wc+45dDkhUJ0kXFajVV7uNkxsaoyET5isw
5Qg16ke/wk2JFrzbxYIPGEmeBp/douSleHyiC0MOpfYviFz1BQrAq7f5Hy8x
kjvHc1LNo5CkWg/LNS25NMgd3gDkcPDDQkAZcPiDoZr0Ka2idpLo1VonAF9X
ikBin7jL4j5Hjpkdt9nDOMlfFhwzW9lO8NYVBJvWs7tkdqVa1IRiEcVDATHl
7HLzo2+/ZeICuom9NlQHjERwLCSGAVXmoiTV5VL3t40UfQlFCuygakBHyCoD
0SBj23NMjclvXw3/GFEXO9RGSh5d8/1oVUDhFWYOFQ99WJjVpXeT/DhjnDt4
GYre2CyPtWi7vZ0xPuDtGU0944k2Yus0OKlrT1verXi3pZPKsQ0LLmugtfvG
Fw0yMfvsDWGH0TZrV3iFuY2cCCgNTp/rvPDPKkiuEaVuUD4AdZYRukTNorQD
f6re9CSYtDEiL3hAZ6OU6pobQ0aYJBTkk0Yx7uq0bQMdjBuFF50WjhfLwqMS
pXZ6dJraC6gKoQu99NNp45HdA9CUU3eUCLb1ZeIEadVL1u7o+o4e518f/g7A
DeLBZQMbxIw1N/WVt9x5oHsSjSXioLTEJkDEOTWNThH/rOWThyYAmRq2rL1J
X01H3QkPshUUR95GEsj6pzi/TUCTUobBGg2L2ww3NogHagaUbSqUdJlhn3yH
3MoZ62spsDRysbNRm3p4mK7oSH1O7D8/EODRgeNEXHF0OpkmCRXkPDNNPGKS
8tGco9PcyEc/3bYPeYeOXTBKdv+fwX+OOQCixwCCvzmZIPQWVqd+ctLd15G9
cUD0eDwP72R7OMXPKZoHn+V0yuPCxPThtiQsqU0CLOhqIuzGTEHjMy5NiJDJ
aYLYK8sSx3ySw3HJlwvtKjmb/Qe2laRXfvkrACgc8VR54dl11hyTfeWOZn2z
74kw31NZbr2rilb0Nie18dKenLvStFsmii32d2UzYZPEgMwQnRLb7C9rYGPE
M+7odze4gJBWfcuFqULmUY0yMNJvy6vImzdvkMfES4DUrOjYaRzjwnZ+bb2G
3MW95UI6b6ULKUMYvhij27Ah8VQtIIKLxTq/YM7X0Xjfvklzkndx1sNsPCZ9
GIP+jOEqwwwpOeVGGvuNYHSaYCTO6a9C/27XE6AMMDUVPB93Smd4dyPClud4
AcFZA3/OuNxvWGnxd416gqTnVKbUVqm7YMmiELpDn6ARjetlhnLpf7u3MXus
rY7sdQmgz3eGaSd5mc7w5Z4bHcirGFK+sPCtnpc2ZYpt8FYmIKvCRE6mGjI5
JOHDoMzTKas2NYwyW58NLv3ZNhfXH/LNaF9LFTVDTfYpyMz9JwrKLtL6E5Rp
0dxTDnhxY6vGyHP/YU6fvLZHbHItShHtaBfrnuFvmQvD5PI9YMcK7lrSpLKl
bYMagZ7oBTpRzEQxfuoIzRocttkkLPVFy4g1lHnmG1UziSlBZ9wrN8YtW4EP
2zjnvYjPVGE7BVGRSnbuZrZTKdImWpmejE+orSe5mBdQ7SCwDMhiehf8xK8G
sfUsEJSESuNt2ubudhLqpnNvqjGfbH/U3w45vIXkCSJVaKAdAHc5O8cBwu5k
CHLHmv77l0jD+NfHQkRF+h5lK5iTbQe18AQPAk5E1S+VMSbHguCZpCTLQMVT
vcXY6g1V/mOcq1QTRCTaey0yevWoHr0B7IcyZKqCC1Li3Bmz+RdaIOnK2mlT
htAL0rBpCxDsF/H77ifi6YsxnHCZZSlJ8yooPDLYcui6yBLIVvVyuYk3BJhe
Pkf3loi4V+C9uJjVnWt/kujgrnYwTtGlf8we5ocXFXLMhU34cXsmFGCYwhlx
k41mpy5u+uRIdkj/fh0CSWtsRPRYMJAZnGsL3wo8+LdFPHlPMF6hgw4lCnvs
pKTl904xWPURdjn65Xr/2qmGWnhlLrGaZO2vMcdrObQxeLpmUaEMNJUSwP8F
3y2saHLVw5dWkPfmjRg7//dEKHrIIbke1pBBwg3wofd/a0zIx3218r2HdshJ
ZoegcNDwmiX8CvqPZOhJPxgwiWbqe4PIiPuodbVw9cnpJ+cFMt3G9Pip8OGA
kRnjhCxY2UOKG2HFmjigmHIeqQsr3aJM2jMy5rim7lNXUjguNXnR/njBNJEP
ToKRQspAEk1EnM4QbIh+Unm0Ml46JtzXz9C4UjQsM7fCZXzdqrSj7tEW6kyG
SqzH87xeGzkI8L23C2kEEdOD0a+Cug7EfNpzaH30STG4dWmfrf7GX7lGFyeb
1F2w8PAdUw3lJk1Zni1DGI3tMOUMPZK2JUgjFKloX5vpKh/cDtB2M6ruXxF8
L8KNKyCTudMwptOhrzrpPWPM1SlNGgktkPLt2utJf0YAKU7p0obx0AVI7kB/
xvp+TnsPVr70AIkvt7zjpW6gaegEfDwHMVqWEQHvK8VOobp07uBG0qtW48La
8UIN8uGY8o0zL588Cqf1axPhKcm8zKqq9ULgr2iJwpgM+LpEoqa8foyJ3mwQ
ejWc9gI3CXcTb0iKGoz+RfDjzUiglnPusV6oMS+2Yp+OUVC/USY6iAkE84gx
YSkAvCdzYDPCN5gfH4dmei7XNuJvWDMAGB71JAda3BMvZ7Iq7AvT3hZsI09+
pqTURBQP2htc2p4MaVd0fDyrbijZetk0+HMw8CehemEICiLLagppi7ZQU+df
mbqMn6p7A8qYQO9IweSaELE98PnBbVZKeig4cdl6njdmtVhYNBQdhfbCDFfT
nRpFSU82XB/GtGh5ITe3EkLenfHLvVlYUV6zE/w5ceuMoPkPrP8/mzASyLtZ
ghUT1RGZtQwbqkS42KJJukPhZG0gj1x2wZfn36h9ASU8fooXdxvVIRGugoxP
at/dezsjnZS051nZgmbLhM1JX08N4qPr8MEA2mBUfAu1mWAehimlbgaJbsk1
lESg1koQQbrefSboRqvTVp/xvWjEibK8tYCR9K29MKaRnSKFR9i+wJcj2GlL
pIiyv/OvvkmxA0102kE8zJIav8rYAzgt8UEwAOhskX6Ta/P0DPfWVPGs01Kt
Xd30850yLfKAC1zvasDbnR1YtZe+jB+Ir7YVXrhoerea8Tw77T+y81vJbf9q
Euyy4MYJA6vzZu2kihhJgDHRS2TUNo1AsLS4a0xc50qIbnel5pj1IKmLBjwA
uJVKcCZnLdff4/Lroa/+wbEU3i2TdWiVthXPlbIKQjciwMzfnxfbE5+BuITH
XNYulCRVyH63LE/jCJI/f59jRwXy3+mGp8mfcXAW892921aDksprX7O55a/1
UNzMgltBJITxMUuuvmEZs32SwNPMGlpsjdnCGB4A/iPiHdbf1l5uPseYiug0
d72A7NsE5czWhuEv7Gac50/DlDp3yRrjSW8E95Tvf2SEBfAZs9BL3bnKI9xD
ceaZAFE9U/HFrNCSgvYVsBpfwPm+AhdEGb6+aO2HutSBOExlie6exXHfMnBT
Nc0Ejy2CqA1Q3dyXKV6nxv6lij1v0Y/FnnX0tBkdTkqSb14f5HCvosr4Flx1
V/7BGc1RM9BxlabfLuTixklm9Qgw/zkiMApjXq5pOBsM2XL1txgKhxE0X7nH
WLs1Ugk+/L9aNA7pUmnzJBeDNRthKjEy/YlIOgLRrfZ8REh0TJjDZY4r3e5Q
zdCyi1zkj+qE/6OjmFVkQjRhrVXgOG8qYysWohNRXzY3Gb0MZtXFSLrIuFeN
cBg5RwwfnSKsdkFwwxlJsL0fqexV4kBFQhVQnH1h0CQ2kLH+1l+VhlXHUFXK
emRWia9UMGibh6k0V6n4ESVjJfzojhXMVcLizSi9Meh4YI8g/z1VDJ6yJnVO
dtSLX/HTvrsil+WVPrcAHnqO2Q6P9lAmBweTPzVnJsZ02oknlTxShTuUgWYR
9aq8rp9uaTY0VozaltoHQu4OtTUlXJB1wg2XYFl8ZdmNdu+xF9otzCfdEF+/
WS7c/1peMMNb8oTjVA7xyfZfeNRFXqnVtO2iIXwiwSbpnhYDLSSvjJr+wUgf
DdlvCtZLGkWZCy9psSSMiKuoKK1Zz+CZ3hqiMdhV/F7dJGAnC6e20e3/ohJ7
pQgv3ymM47gGR21aSt2pee0znsQBCbPiRYpL7HYj6KLjwlVEaQQNTfIvkAvN
N/g41gLf1FOV9nAFqGCRPqiJBwo/ea8+nlBxE8Q5OlExpoEPKA2PfNqC4j8S
uVchcwQVeOmoE5GDztIWIOWPixdjOOyc/J6lPGaSFCpl/dwPsC9jrpcnPh3A
mSL3jdkVVA9q7nfE6yt2UFI8jhHXj2qKlsgDOc7VJc/spVRTV/UYvrRHei36
232YZHLAwm6yce1fTsnq1fVatvk6B1/uGENu1BWW/bF6kLhPl2b/HdM2IdoS
J/qbSnwBaMuowOqnkWDei0hSO/QayOvYoTgpoWOfLC7L/R1QKBQKniaw2Scm
xa1ie0iEL7XH8KdlzEeazxtmzsDaOSt8aDQdjOWQb0xe3lLPUFF94g4gDBrm
m+a1LgkeEbDag8ity0c4xMK4lgrIpe5Ju09i8Ujz5mdrjaOVo+LTLhyR3R1D
/C5UCFFQXTGHANfjvPEBzISVaD+jtz3eZVr152OoVLLG5oFSYRxP9450oBzh
t7AxUpcOaznuoA2KUY0ER59/TWDQENFjd6KI0zzyEu6hrBWH1EhBIxWOBzLW
hTtoMPBIMaFi/a3yDF0Y0cidmbuQ8zTefXt7FkLLWGfuLNJu7AJm9cdImhTH
T7QjWnYk4aPxqax1AiZ+hEJBaA1/g7fVUlwA5GnLOBIY6jNkoTt7NH9siCzO
7LcQYhCLjY0Pt34TS08C/8tAKU11QhldIv4Jko8njz+8hAuJ6x1IlMjVOWZg
exrkjp1Wl7mqAwvpHriS7jTAxielu0sQw3CfQp9xzXzHUSgtpTYwZjrJKbi9
1EAMrcSB/0MyleImZIblaKmSIFyBk9hHnuU2v3BqxXh8Uu6DHZ85JDfRnSC5
K6Y1hDLdwpoQNRsH+uAWQf/qhEfNS8rwtfqI3hGj1ZJmDGtagulVI2CUVcf1
O0JRexlFgmgFyyZ68gm5Eiy5tQkicmH8vWGKlEgj/MooZv+V/RNhKEiinOnw
BQ0RlPo0gQFhpzRQ+x8pjndXitGPNFdW3GB7v4p9hP4m43sBUrpQKD+E3pBW
j+s7hIuXMwQ88lB+YGBKtXAvg6KiymunT+zS33mJe5D++EULiZP3IBITR1kR
kvkmBAaeMCauxoKGf1tqQk5S1QBBpcks8AUzBuyI3YgsRgPR8jQhd5+hjgMk
KHnfslwcqWDj87ZhXmhJvYVhjctP9hrXZxIrRv6ROpqvyp8oK/ppxGhPokZC
t7U6uXDHjfBL6WWyVNxbvJrXOS7TQDaJPxja62e0V8vzqDUh04wG5rh738F4
1dOnIUFV+IZo8LIlvCFqhEPtxoNRMTvXxkPwTCmt8xO91q6fnBMkDtKHLh3f
39lZA8DRWeLN5pkorge6/sSEriPvaEx76wilQdtXF6aWq+nA+itz8JJOtuKz
ESW5R8N5C1277o8YsTzhwVvTlYBevnCPhuxjGlMPP+Ar3JY5wLZofnaLreeG
28N6ChFJL7Z6ykMJ/C26g00322Bz9i16m77HxRsEDCYVTxFUK5u1/lFwqEgU
Dlkcz4GIquyocUKAWygeH5TeSJhELueOL9jjZutJLpYa6D2O6M16aWEo4/Xk
Wa+PlblKEGmwFX0PtF2R8fuyg2blOIqqAYqvXTMSasgdyW9po61dEjwnktoe
U3eTtyoX6aIydzBsYYiE5hSwjdDVv+Ctn+qjOQLcrXqGCVgSN2Lc1VeX3lC8
roM5iS4B+wMRcGEw3HkuimshL4usMqbvY1LQSUbZk+GDr0li9M3Oz6sYPfA/
9fIoQtnbVs2fS+I83V48fdf4QaPfCm56biRqFbryG82Yh+GN0fW3BJWJ0rnp
PGcCdBgG7FqYxM3rcOMM6G1/9X78pspdvTrOWwsytlAO3rf7JUUUHMafGfLt
7zwh3Db2yN16Rvv2uOEoo+f3FtclzsSjtStCB/3yOnOUdwcllCA7H8bet5xV
CCpLwh9ecMRJpKy95KqP+2KMLCWzu0Hr3zll546AIo0ee1jeWruyKyO3d3st
YtGqrnvPKEcnpi+2t/kZRjJOI7MFaUEmXdTWqXNJ2wR3XT3TVByz7fFJHo2H
ocYfmym/JqLOmrCUH5NW/IrKfi38YfHPh/dr9+kSL5KMhpJzIuzL2oujxwTA
xjNWPc8C6sXft6yl31nzOzxmW+Y3aPZVZi5ywc1+Pzj0Zn4UnI0ad32pg3c7
Tm0/gxuLgORXqIayRsYZQ/JxstTZGo4D5FEmbcU8C/e+e5wDD96JJBco/FGO
T8JOAJlmO7Vow9flWSZxSV2okUfNKFrS+71T46U/1EV+bQyo7FeXR5EGZVtO
f9iURKJlklvizYh+rr7bdwr9WGKtbEVyzAPRDQ8lIOHOQJiY9HN/CA3RqApi
jF7SKl73pSGq3KsHdWvF6PJoQd6CYZ68wZeVTjfFu9vcEpgK8UFPBbHOYAaN
HSwowybapfJOdoPd8KiPFFNNQrbveRbOA3ebxFc+w9/IaWXa2vyy3jcezW6Z
9G/lnt4QG0xY5yMsVWoMkFkMa0JY8zgGJI+AxC995BkjYMvVuWFnxPeI5UxJ
LFxwCgZze7HGLIIF0rKwf5NobtgrCxQVoqcFpbTojXD+5k0UfbzpawZQKjMs
xTKB+fssbcvSQ/bEPxCbMP+AliP8DSELtUUokeEmrlX1RMskY3ukGDbUktUv
U9KOs6xlbd3xPXtXv4NGaX+FNgHrvRaFyFGy5BiqJIl7Wh6+svr/Xu5uMVaj
jeYXzLC3hUcuk4Ni/jI5YAYYT4VJCHH/cj2ZtFbVdwtXC9qQ/rj132k1VsFa
4njW69L6WN7iaGazrElLzTjRREYmAiHWquW2g4MUkf752X0KEP6/vvayVcB0
oPtXE1mD6tpaKqbpQlvuSElluzvThHwSd6g1YPsnex8oTSMDzvdAsTjVWNB7
0GahVY8pKSz3/sBFvHVRhgUnmjlOJ6avN9lGUm0HzlSiGPlc6HoZe5AGpRwF
Pg7b8jLy6CSBKcRmJkpmVLhEKveztIXPMld/S4X44eLMA0bAlbmg5XBz1AJm
5PHcw46FsqgSyp3Q5lfnHu99zZYof4Q7ykuvEvg+x0f4cZeW81XAa4CxNocZ
/1egWUuEmcKd/QfDDx8DKo7gx9Lrp9PX1OmgvbQ1rn5kbWuqW/5egY+uq2d6
1H4RrRlyalASUp5QNn4m63tJ+MGwBj78PO+l6sEutgqCPP1aqa8cNrw8UQ2W
v7H0v0gOsmlTIK9NGlU9eiIGZLS9RngViI/4RN/f7sLSMrjAekI2ZEgFCYf2
Qllt6hb8GLPAxGgKBEAfyxFXAESzsltCprdBbutn0iBDqp/5CJNiAlhEFuCT
m796IiDqgl2Ehx1njJtu/cMSBpYVyw0VDlkG6ctqgf2WjgUx7/6v9i7TUVed
5u5O//8ZQ3toCKChMdfpexBvACmLkbQDqRRx2XaR/y2TOGkTCxitDefX34Vd
iIlCcjBu9J+4Xz1stVNsVYh/tC5VmsciX+6wUzmh7x37Db3TdLGosGHKAIUz
9H8P9efBGNA/8cvqC9MjbmCUZnxT4QGjzTARw7W/rQrshJFR+FtJJtrLo4g6
htm2jMOBlTGDp/+fPMPUims9KlddW1MR7uhAZnyCQ4iKx7dIwZb9Az+6d7eq
7OScer4s5w/3HjQGCes66bo32RNEfUZnosawJ4anG7WA5Tvl/MQ0JRP5oQuU
817OsZ6UtzuCXxf0Y8cub/nWEvOTsrN8zYeT9WP+Bh+Zc/crdiTYVxUbGtLe
fTjmd/adknSGdZVV2e7neqi6VnN0NTfq91mnbPGAHPaL6zAaL/y4tZ2TTbnE
AkiTwIQmQYF6LWOYzP6Oj8+GzknHTcIJM76mv4gODkYhoihoqZr5aIy8G2om
KJBQ6wkvc8Y4tN5R6qxIQ+DsxQXazEQ2MC8lDlEltZgpmx6zQu5rThUVvg6Q
RNYJugvsPY+pd0SM31R9dqVwng+YgPKYItRmhuT8mUjhdQ5rmOZ87drUt2Ou
bWZIi26yt/kGHoF/7TaBDBtaDVY2I3RQtNOgUBLD31lx54ChEyXDrhSUz7K6
Q9ymVnsy6SAU6i7QQ3PwSYk55CBYo+wtHljR3QnLo4oha6ADCyt+JgyUxn8s
NkbcL2zMy+iLMbCE2UWINuE/kZD+wLT5vMbIBCtYjsRedIAcTuCKGXK3npJc
yM3eEXUEqUE8YvPjYlEttwjiji32a91IeT9D/dWAKYMYDR6FWBJnmJ+FYmqx
qEiJBu1saomfdFOGQ2PtSuRmEbVUWJbfse/rDbAEaiNrmlz9zu64LlELMLTe
AYg4V6DTMO+9Ma2GFOIOYUoQAGASByiHFpMmnZJkZDfMhOtL9fT3HwjnZVAR
IiL3mvuwYAVQuK48ZITl6w8U9UKYxkVM14EIma8zDax2IIl/mowSON8XXbo4
H2gZy2pBujcJZWo4bE9X5kneT9QKmsvBdyhA1hmoj3M8R1w9PT2ambbO09+p
ikkIdOOP2GRTkIYA5lmQDJoWbV23dORdZVryZelH1VoGYAdoUHCL90Le6rag
LsqKlnwcxZ0YidFcO6wbAaTeueq5VSDJJq82WB6MHf8S/pX8gRqmAsyAkyNY
SF139uSyPmREt4o2zTvlF3gljvRMZjtHLHk05CCAa/HmG9jlX8Acg60vffmt
R0tugdkTl8p4nsaUXwNhyEiNIekn2i/9OXu5zypTRSjuhEFWmVqnpv6Mh9Tr
mEJDH8+VtWujI2SBwAntrJp5GiJn9TJ6WjKAc/NZl65OSSXHfMOGg2yRwbTN
zCVeYs8Lwgatm6xxfAyM755atEHRFLv/bxRR59P40D2qtFdpuEZxe7qncPla
mhXIFX1OYpwdeeKnpbi8IWVG1/E/b/IRPo/JL3u+Qk/Dyn2+IwQ6/1HPayNl
gpWnNAKfYzc1CPRgVfq4h4jrkX9eCUxaXTlEbGiiH1SDCsbBZX/Stm8UspMh
4k7o4XpB1ZUhcd43O0ohzLKYE8xw3KC1NExQywd6BsIco4zYN7XkoXpnBtQY
qDn9tORrMAEo4zXFQStiBr/jRZaN8ftWEjKXCVNw9MNby02a4i8mR54NYNIb
UFlDYNd2ekuNCJ+rzSTVySlKeJWPAvM7LqieuJvtQIV7Mc/zuL3jKCcSTDcy
2OZLpbPkioaXhjB18FjwVddZshF9WFSTzcvbn8IsK/QSvJqto6uSgDgh7dff
sPGywlm1uOb0F3vJiH4aXyUj8ssdwFhQ+iIZlqNKwRvwOj0pKBNc0PLt+gmF
uV5EOmZghsP+ntP50FRXYHgDoGlgs4CSf/ZGWZFmSqdaGpQMVSlemOK3Ng5F
XSmFMAQ3ySe9KWPAPAI0L/99Pge/YrwbFn/Hu30LN8t5WOkZqrfis9riZ9K5
20L7UiRHmKQNMpyo7w2sKgBaKOzBdKQbmnRrc6bu7AtEch4xExlHqfbMGk3E
9gD1ng7zTYOr05bZhshCwQ6T6f9m2p23stOpAm2fAX3hs8/13BuXvofBpC/+
6S8eJunVumYG0hsXyy0UXoNEvOCy6C6QLN+X3cxlA103fflv74S0/fEzXOcS
Bk0rIqwb3+6thC7mZtWkD4BKiwl3HgyWU250JESncQYT4aJmxCye8/N+GoUK
MI2yrBY2IlHLxA80xhL39g5T0LFvZ6v+dOXYGXCCHBwjztO8rRxjrmr4sekz
T9L7de8ta1uaNlT+FUvr/NYFCxqWqU1AhiaYQds2/CQiJOLpHlPCtZorQvu2
Pzs4gPGSUaSp8As6LqQOe8kknohHxy7HXSiZF5QRw0Q0NYYdAgX6W6Hz2yjH
8Q8qfUyB1k7E85torFNNfAYl/+cTpd0sjTxFnPbXWS8NnXxkXrvLFJmBVFt+
Aw51m+Kqsr/BAfeO4+Q+lnL4zxEz+kc3D7vmGoZdqFhpF2ziSRhZhOBKK7TU
n5FWZp4VZv7ck3tU6M+cNwij1W+KM/pRx9QSJf+ghWzZe72hr5nN+0X0Uefc
Gox2jnod9aN5YgR8ZlU/jAxPV/DpJ1x0O8Da8ZNhlyUI/lpC/r1N3h9F3RBX
+GT+yMrxEPwuurc6Ze2KFxRYT9U0zVi9KRTeiXVFB6t4i+yb3ttGnv/0h5z4
YEnuUvCPY/FL6mDfaIR592kqcXa08Zm27tpbQL8HF1A38Dov4HdkvnnOnDpJ
PXXVxLbmb24/mpJDf18+QqVwmdt40n5j0u54TJI5rE3LHZtKd/PF147D1fkK
qmXNdLsk4OkDSqnUwhSqn9xSXGZ/rBv5Xcc4YuCNF10Ko75nMnt2GdRcFxYW
OOxOGDvm3/X6geWs0pGiHpHMSreiCOVLmLG5Ft47cdQZoVydLDKUzA8h/Lwy
nmXbyF4z9Q6fEXbd6Kt4cFLDXErkNV9ugYrNg5OZDRTQnyMaSLB76Nz5JUy+
r2l/ZT/VSZI0GTJp9Jqfd2XrEcEABApX24QOeQczQssM2LHHptIlVYW1KXeS
jmf3tZssN9fRkPlnyxlLjTiiWVfHDXWI+jmvwfFYtdX8ZQIUfCtaRb7f0rYm
UloA4071XwUjmd/C3g3A3pyfPaxb2QRDVlvABW7K9M3wOlq53/8yV+pdAr3w
ROrRidTyR8Nw/58wM4dKS2x1QKYIc8uqQgKb2wgsfoXLPRxN1m6isynwIxKv
ezYAHUmrIk+elcb36f1VSyDdnkN3Ci62/LlMdxiiuZl9e7jwbLLQLqr4zGTZ
EFO7Ol6rBtaVy4dmbIxuE8Vryim8oo/yGLUTaP7vpKgLooqztUl8iiqSwa2h
EgMTjNSwVR4dVV1kzGqTW1awnMuVd/V4zALZaf7IJfD65ENX2tD88PTr2So0
6bTL5VzsU5R0Bc2q1NUculiXqhPEvl9+v/wfADgvFvxXJ5QqHKNhiNX333Bf
L2Oj5eF2Fd1S+r30yYMZZT0S0klvB34Pvqeazzk3w9eNrQO982t2xc8PW9X4
La0MVPdk1JPal6/kvQ8HkB5fUWMGJdxLX2ZaDC2+rF6FyNan0txH5I98wh0T
jteJVVN1A2Rifgjii5Ma43IjEjObHrSJlb1vFtIxvzeIRO5mNnJLlfywbHE8
iOQxB74liUl81udAyPDbLpn/Ntkold15KcV35rug4A4grviZ0b2WbtFffNhQ
EgK6S91GBER6I6/ZFKXKC5Xntn3WuD026yBF6dVQ0qWnc8sHJKn/D5G1EgI9
iZGgFGP1DgPzGU6TjoX3z6nZglc0pZ9msp7WSNqwORNgCxvM1o3n3nZKhC/z
7zm7+RKBNqv4+taSO79st2VPCk/S9+fQthjRySH6Ee9lAxhZQ/FiqMiAWXcY
RDnDvRHpivOOp0aCAMgLF8zmUvpysgRPFgWT6OU5eNw+ioTOpREj8nTJVea4
lfGL4YNv2rFuO3AyWw5B3nu4bJkuWXcdwgD0att+JtIUBPVmwe4Wumtn2Cka
COaepppdnGxRqKSI3rzAAeSGbUtDIi5kpMmlkJ4kszaba8DKsiFgpS6yhpwn
8aKWTie8OIaDv9Fl2hDLF7rI5t8YQc1+JFE9mdPA6nCwWBwVz6hijkaL30cv
uiQU339v1a7i0ulX/fsBu5TAeIMiwQIVIfqFVktr4j179+3Fe0DaEYvqPYXX
PHyShfKGtBRnapXxf67r/QJK5CHph+4XxTBOi6qIdjQKU0r5t53d7AEdrM9q
PP26PTMmkOR8QGZuuW3N6S7gI3EcxXK0kYKrW7DFFIjCnCsywbbkYVBfsGCj
/bINm068WWDpE3uUnFOCveTYJQ2WUNoUkRyj5piZNt0etU6NeZ2fq889Z/wQ
oRatzjzsXy2Ja2AWAK8icSUL3bxT2QrSxnM28Fqk9WZFxd0lVUPUOP3P+W5D
Jx5CRk52a3h7WnUQrNLfNwN7prAE9qEhwZ+kyBF5Fg1iJUHh12OYECfoLcGF
PoerYYbCxMO32CqvnNFetrRECHWlj3Y0U3VTwnYQf3MwEgIK7qWhtGcAZEzu
sj2L6BcFbQ6UkBxE+ZFdqmRIskLd4YIk2A7pgknB7hIc7duU3a8uSeebqe5C
byekU0Idwbgi4iAIZHbgq+CVnju01KmoORPMoXG8UyaBAdY11W1RRlBp5z0r
q8REx3Cz+e0npvDA2GJCcomxUbUw4ADAcLt105ZMd1qb9yvoPPxEFXu1Vel9
FwtyJP2vw7NCfOEURKmNboAiUi52nZa7nMVvArsuo6xiXo+R0z/Uunbf1Znn
69w70fbWlnrnHIWzY+GxR7pb2qN2mkwXNwUVUbyYTMHsCv05ylFTzyVH/Wa3
fS2piHhhcEu7FevNcC5xl0pov0M7wxw51XBQj8XRTxh4jfxuvzQw8Mh2w7RB
u2x4YoB2juFbaSEn4d1y5bj9DQ8IUZVVvBMfSiMf5K9t5aoYVR+fmrXJ+ypX
1qOLJ2MfAOVuvD8Vo9c/NytR8yeS/EDPji/Zy+V3Si8Ft8Ew5i5SgBEqP5bn
xYsp7KNTwiWffm51V2AWs+h/9kLiWGxS/cpI0V6DHNwmbXmJHx2c5QXYSzY6
BXjLDXSHabOgGRPQpaAi6JFzFwjXd5moppGmMh4et+A39RIRcUw5ageMKWpd
sCo6S9njYroq1AtHV6VzLt5K93L0lOJ2ScaFHnP0FzoFfmmBsL6nLhFAMy4w
wvfYge1tjFqum9+gM8vbjytTQyF29Vd8AFBgM0Y55soVve9tgaKbd/+YCdxJ
y2aw2U/o1TQ76jPt539Xa6NEBsLcjTVSubk+/YrrG+MCyvGLa1d91zpSp4+9
ZAIb96aMVewMIiQpPNzvmw30fZJvxtZcfdNB87RW5CpoUDgpYiZlYJ03SRNF
RLZnMGkhrqcaLosSp9YbfFR2PxH5zPHnx3QqnyE3W80ImEjlekRUZIWpeGtk
JFc4bO8dDVQKZazizYOWB03dYtuuEp6EU4n8e4m2tCSsMLm7954TwaSgLCkK
/SXo26WbGooCHraBNXIEWxEwrM2nEvF2+5sWMS71v4HBUOU9TAhinCUpYaxY
L9FnpG7fzveXEoqLKMELoy4AxVW3qAYw/0ec5m21+kGH36YddHkNfNLupkPH
e7yY6qXX3pfC2sBUcGrSV+2t36rhDZZf4axSi2L0iS9p2ylIFCcgcJvUwXMn
/xYVt76KLfyVz+9YQrraOXd/rZDytn1fHKA4bLQqZz+zH6FTP7biLGLD+V3N
nUhKi10YZQb3rNhw3UesXBnmPiwp2PmSrX1y0yveOUcpjfQ5rvA3u6OPEouN
dit3mJVbNYrykCuLfXHJ48n39hc3juDG/JJwQzrkW4ILYVJQOJZB+UaebNLL
L0yUDv3Cc9nTU2N5+glA42UpY9B/+8/ORFZdEDtmNhqcWrkoJO3vDOjFg3ys
eh+GPgGfKbbp9/dZxZgdF3u6zksz/SXExCUOtkP3JKmoF30I0j0YWNSPUv4v
S8S8XrKqGZu1ru7kzsbUIatX8JtXXezBcoW924eyWER+dQMfvmq3mi0wOeRa
rsI52ssys0semM2Gogkh2DXJVP3IdjeZOOEcHNEpFhsk3VAnxFzu+5V1iAhp
06/OlMIwUTC3JlGqSnHQiIyKSYp5BbkTEf+PvMJltPcUXMw4Qr1z0eyRRKZn
9Db8JvArfOg+C3/ogoNrwzGPLxVGqCQHLA7frR8mfpOgS2OL0igeDKIZdv4V
BtOPAzozZXXRsbvKdAnu9CwLvLEE2VY/Vj4LAYYuNZ25KfLFYBDVCVD5lc3g
vMRuKMPBMUbUPfVTPkNqJertTh0JUF94xN/BnYuASaKID1KeL4aQCEG/VD6X
jtAkFjYwU1Kxg54sFX7wFz/z1HYV5nmbEIKz2NMGhBJcsF1Cljut8BK91K7b
uhgaWRhmQwvCBJ1nQmEBEUiaJDcVW2foAdeyqa4DPKEdoeNp0wbiwUMClCfK
z2pWxxLlkoNbQcMCvT3BRQ+I9TH5tEey8StfIANWtrepTkczxInAFJqn0mRn
nx9K5xbNh5bRiZobjI7ivPPbAj1REoC31tI5cNc8RTyNFYfr9RrLB3pDqzZ+
uPw0EwLlq78HDo7BXGYwlGR0xQ52JGa1PIfXfQZKEoCrecUO/6EtKRL8onep
1rasEde4NoByt/09+sIzmXxQ4OtawJHYtF0ASA4SqXJWzXAzni3FtS9/lwx0
P8bPjQR4P0sTKvpQa1stQSDuXc+mjQK2NxsBq5Zk/JxH2AFn24oFQ0j2TnaC
AyUvt1eRAsannDFz5D3c/XLJYXfDfSUErGD+2wpBWFhlg87AlMFgO8A7Rktp
ur/a7Y49UxAPIek7n1nIL9CCBi3SmR9dT1Ojv6r47B050CT9B5PeXKDMTg/q
SGC9jmhzM0W/pzkVu6bR71uN2AjYSxzmsIfYj40NVIjkNLjslb6e6Z7fbt05
/wKgBmC0mgrIVwEfQVr6qKS3efz51NZxWyTjdWAE8I/lGnaJCCo3wIzQZCDX
ib1t/moSbseWwhjCC+CVyybjASrViKl+pEQfXcI6ASVO+HAOgpdl0HGb2nXu
SSlJM8GTL8eHRpNGa4YTUD+M3WIv3Jte+1aSuE6BKcIgqlNxxgtLjvBBEnbA
tsiGjSMJJIbeKYUVkx5/zEo9EemqKqD5GF6F51uOnaG69SpaV8z6j3Vs+Xv9
ewfZHEPjkVOk1B5UW3Nz4fZGSBt1sLfmZEV+ORNQcAJcrWIlcZOjuzoK7+Nu
i2WXx0WQyJslAgWaOi9voORdUVADyuwMzwMGvlXiQzQiMzWZXV4M+/gHgzyr
dUqJoHp+JUE+CEIakUNSQn3Ako6SnXgcM/IKTcMyZbNXkGyzzh7su2faLKnL
bgziEmAQzmu8kFOqqXFwWHiL3IQ9x/wXWCtAiFhoh8VFuaDcPAKhTsMy0S2p
jz/+Kmt8Lb0iLdPCn4qfTdVbNGsCER/S2R0USE8cchE5T1PENCsJsis7eVnW
DL0rHDJF9M04PjHi8FvpPa2cHeO6GgXL3hTF/t2rjvw/pCIjcKKyMqsKMCYi
C3f1n2bN19owT4FK7OWKxVeeKeu6rCBuOi+bYYZS00Oz+QrsU+wFNvk4DpnI
EEZ7zz4naLTQ/+7/3DJUmqjRr98LAsfazEOUyH1HhDllmrDFcNYWvDChodlj
O1M0qEaAUpOF0If8M9onMRZ3H5ZAfxDPmC6G/X9nXwXf1dDQsFd/hhYTuAUI
Avn9zPU9rzK68gBzFs4PLXbrIzUDnVEcEN4W2Db8FhXwrxWV4Ds7aNvtENko
y1AVjBZqOF78j+nzawxzOQvouoOL8QjVnse+qnTemQdi7TCaF4iraS07t0Aq
+1LOqHIMsN2FX8ZUSIzdqF1pPPy6YXP/6scntGdYmsJbQ5s9sE7y/TYg/XqL
ZwEsoUO417sIelg3kXqUtXpSTIVvyhx9Esh5fZOV0JW3lRWpzHqonDbZd0L9
9Lsuk9ucFKH5Tqsn6mwZs8CR38O9OnQzYamyoONWFAt7tvu7vq37bToZpasm
cRru6OPW0vQbFl7ojHE1/u/ZlPLigRX3jHS7+SaSt9yIFetx4TJEdcF+IuKh
XWOBtXSBXmxvDVZ0IN+PwhOey8dtzt/p8Bc7YtAojrj481BOLXLpB4NzPLtD
z82vUQ4rRV0vNK2NW1DgoDbjEIfuBqaNV/WaYWeBdA8qyPQ4U8lxhI0skaH8
JKpizPzQX7H+cDYYuAgUeg/mM2KQcDnAFcNU9RZ+YzVr10nc7DQGmcwywN88
IrXW9JeiHhlv2dCkkEa1undCM1yA8H0GLQiQOfi8o59coqZJjeloLSsXQtRl
o7ip0NfEPflxI+aKtLcz1HFFprQPPcr5vLmH1BXEIEGibA/iB4jsqf/j9Eba
g9eGUSYWYj1kc8UZYUgeegqjX07bG0cuCoXEQIM54WriIO9GxSN1hqcMGVbL
ox7FGc4b6wZskIY/MrbDGzRSO616k9hASwIizs4LskGy15o1Xa/Ez8ENvjfi
oscnWMa/x0/5RvKpGDKWGCD9AciYqNx7TKBWRu6r+78pXOT0GaH4MHRl323Y
fYR0gUc2Ewph0dw9+hb/bDPL//au6cjutd7Fnd/HBhrgXCVjTx5lHO+5kkaq
rR/bWBjPiYYjn8ARxspPVGZjvtH81kIWOVTds25gaG9iEwaThcRIF0/Z5fOt
PmjiTE+MtxTsoiFlGn0IK6KbrGA7r4lJhygzSP2SRLLgrYzsPONlrowKqKGG
//Q+WN8gk28ToXeC7pfCuoP0w3eWc208q50BFXc/Z4oRRaBbLk2dHwlOP0yl
+2Bv9D4CWaLgOZa1izZld5BV66nKSXDHyNZo108MmEYU2Te0irlVUMPLsMND
ymL0tM+cfckkjEaZBPqM8qI8+xiUDsnaaoslim4CXvqx4FRC7d0WY26yzZVZ
CGKNksdOrn5KQmGgFsMZ0S4gZkrwN6JXlmJ4I0AT5+Q9gXiNU0de2MVDSXYG
ww8g6Xp+l2MkHQtnxkrPKK7lIwbLG2wUjOFb1G7wq6+1etg49+3Hf2qSWaRX
pxhOxLgRSunwZRePLcewUlsCG2sT7iZyVUOabv1RIY6ygitalDHf8ZlP22NJ
9IwrKkMJiXu1ZBNnavlCB3Veefc+SdsKzzx0KJaJQ5Qnu30uD/BXsrnms7Ei
Umk/f+whSSAVmLm1qvUBWCUY0gKNY1xFf1+Q2Mz8NftxNdmdwxH9lLJeSsJW
EUtp2WZE1fkoCFOL3y6tkzeosMawQK9aXhHCU8zao4OmYviedK5RGMTc8Ywn
rdJZI9Ur7rwIIlJJfOsFpsoM12ADDAzc7A0w7hswL4nzb0IQDUwuY4+9V2s7
p58DFjdJOpDcn0iTdXukyLP2XAuI+q5JLQbQDzZhfdoYPKzfJe0diKnrxtyR
c/eIF+6tqXtR0WLKuttRKAW2pEtP/cUvJ0R/jMe+5M91rTXdRYpEigSBc+9q
s0jiRsZploTkVq+0lygE49VzFwJzZsQWcp0Fah1Fpw34mPVCdfFU6y+lKbbk
MEvGbWbpJzbJuw4OIfYyUNjHB6Jzajf0kpBNBy2Zktopnxr3zLt0r336a2AS
/XxO4HAl9fAvutZSWbHKKHSWXS1r1Fx5ygC4ExOvfPgPMdWKODDd+Bs7k4wA
/WihPjNIUumhfV0/hZ95I3z1eM0fnfhfbvZfnfDZpGxGztyLhmr9RDGNsirS
siQzHAMEPBsVUYo9MAvjUuP6iGjgqwsIWgtck7hLpbj+K+znh1OOYpgsIiYy
8Je+S3kbM+TsZZKbZp8WAp3BXDfaX8ffkk7ytOdg+mFq7lktxd3C4Bbc0MPv
8vEsOL8iAGYP5PLmsMpGZoBGkVtDCfa+XZZpkPgZv73R9SqM1vXosyCRonUC
ROiW7kaT2ugbGfi33i7q5RfurK+U9BQsHeCFVuFPKWeHrHIiUJhEUGW8LzV5
WViQl4eW8N6InlD9N/+RFf+mYunIhmU5LsOnpWRkq/okguQRoM49V70RSo1s
brLggOBypLzERo94jt11MOCXdrPAFK7qN97vCPoYMjUm4yERJ0htPpe/o+ly
+aSSc/2xzcCrRJQ1Kh2te/sXaby7ZR74PlhzIYIhL72CzEKkxaW5I/CRFVs5
Fai8/E7fu2NVKMitrUgTK/jT79Sl5J8zEMTUMRIl7w/lGEBE43ApwZMUhVlM
5jJAghCRoeQ5IHmOtRSZ7GqBARW18ZiDKAaKmfYDBY320JAJaddDC652/yoV
Cm/gx9Yl2L5R2EmBebwRfceGqUQnDjkzq2gQZrmlLylQBBkD5Sojjohcz1/m
hJ2eEYOnHUc4wf5zi5FpxXmpHD/HcWXUMZLa45O3wMtpIqxp/GZX6gVrOVzv
KcjYcdJiHRDXXdh5fqsIzpLIQYT0J/Y4HslED+K4LmlxvvMKHE2Z0JCyYbto
Nt5QbfLjdSws26mNnqpneOd2jkq0ErWX2CHUF7j5HTXlRDWkIXZ6rl7R77N5
a9k8cxd4PhIpB02NoukhWVYbvzqY/tGaAEktYrVKe62tIYzPkAqld7T54Hmw
O7n2KFqs8KOcrDItWMNy2eS8uY+jmg9uOvX9YX48GKw3jhmmMXgrbiriO4ka
fZk4qOWjaNuMd4DFJ1c34JhMw9tb3xz9CKGhfxTaJCV6LjcZWcyNE1vYWDUb
gRyTdvmSk3pcjb8iFA740CQ77dnNjFHSDNEyJd4yOgLNOJVfhQyM6qw6g4af
fYCUZSzN/kXYzQAab99N2snoAs6IPjHvKIMcGMEp8KY+v4PVqUsA8sCuAb+L
LmLp5wlzTQ0EgIkUykIAtDvXAEkL+qOzGN2BhE8+3r+ppuCvbVkGikvHSywu
NQWn+Bm70V4aFAJmSbU+BSY0JkE2Crnh02PuRzMWfAMyiFhEXQN61q6ne7GH
/LsL+kKBS31dbzMzlPkqTBQjvHeWSOlbS9MSC+vtr7amtGtKyL9DTK1mGfix
I0a8BEHNZiXUeexokIGL5l+OsBCs8KaQqThTJUfD1KbCAajgqxw5yEQ19ryw
rG7/utm96F/+xg4pKFULmczba6zut6AZiMhOFXzna+7R1bQ0S9YZXmix0Glc
YAeIf6pW+59Ax1xSMqPtq/Ts6oePZd878R9qnH4umVb0ryQdNGMdeSCkl4EX
urNqVe/zxyTgGztebc3mo3tQSuJbRdQL++ZdPAFKHTb5kiGTZLpEVXYK6CyX
iQ16IGiQ/taQlg9+CNdKQJWQuwy/f6rQC/3XPOTOsqoP6YZwOuoA3cTM89fL
qdlxvvJV4Z/HB2FFcEY2vE12y0aTA7BYz1LIoR5tIbM6dnbbGXZs9RWY2D/E
UDUkjXOndCBMog9hzmC8BgE6Q9QXXO97CqYJNyg4V5Oewhnm+ESxHRuSw9Zf
eu4FRRvBTRsqSqxlBcWP2D78IXGzkrQj1dcOpCAKzflsLMH+7mvXxp2XfD15
VdJ1lDgrVXNERoxiDGP+Eco3SunRw1OprxLOKDoppL7n+SlNh16Ws+ykDfKs
taJdVtwcpKaOFXky+nN9EoInuOe/1/qY5G6VErenBf1puCkmUCQcUIdhmbiB
TW97moGnOkbH3rw1kxdQG3dcSBn5jW48Vyuw2ku2iFD4Kko0oQXjndEt3kxd
GEhPNnZZC687iuNzu08BDoTG+aJ+KmwHMrjf1ZGR2Gs1whvSPeZisdkm6HmE
WHZc0YexMmzsRTH+SJebBvNLnAtOVDXeSpt6ZJeSKtW9qzfYa0TyxmqNHjQc
wuWA4Q5UGuhUXtITBgidutAdNtDDEYM1O1/fSaGDho5e7DgCTMd7Su1nQ3lx
gc/g49JX9V0DN6xx5HiuqI2reehSrc0Q7rZGrIjgdTnaG2rWVs7k3ouII+Ty
2ejbqDb26SK9F8tv0WHnDrb7cd92PAKsiXjihFvGDLjArY5tYHTM3itvvumM
RrVFq0f27weXot3hEhj/vNAXbyVbpUEJ2hnREEeEiBtGIqZ9m5HX3KdTOh9g
fmyGpPPu5vQGWmHwM6JMy8ze5vZ76omuFP1mevDwNoTFbawc4Z0E1hmD8Vm2
brPPwXfCsA2u1zz+RAYtloucijT/J02fH/8nBF4MuCGS93o9UDjNAY2tyX29
vTtPAb/ds8ysgBAkbC+asLXldGa2riVw3u+Sa7iHP0Kn4kuFu3Kan7rlyT18
1PAInVSGRVyxqYAAY2z88pO9G6f0RyX+Nusf1vtVOBYXHfwKIXMnzNBKQ1JX
WABIgi8EvdWACQvIasIZPUYzONoqXEm0GjFGqqDMR48/VS02eK/wQNIfMWuF
4rHGLCbay3Z+vPXQuVNOPB04oXoC8Sx5s8/lPIGxsszr+wgALQdWZp/ip8Wd
l+rRs7zcll7v6bEBASlScgWHONAdbNiV7dhkGEi40RtQNmYztLF5yCyGa2BR
ao3J7XD2ED2e5Mks0oSwUpoD2fc7myeOYNOLzK4xkX7LNy6FuglIXZADH4LY
Ng1LL+NHjLliGQSlzEHFiQQ6a/4kamgovQenXmuYkxXg4JUO2EHMEeGaP3Se
gQhqW7QDvx79+QuLRBzdWnN9mMdhDxynNrm4bGbIgmMe4OTu9PeIqfqqkxyu
0vzNVqX0uN5HyykADL4QWcdrQdgMjf3OOOQHsa6apjQLD5SatJL9Xulj31Xo
DQFRxewkMIwWyvMQxmkf/HZEEz0Y8eyaJoaAhMSgJhzPto+wZdUhlkFIsVSc
BtxtUQgtVeEAwTSD2NZoV6bV0sFC6G5WBoV7j1OG017flx850DBuyCqnSCYS
r1w51NXF+8ee7HZGwRBAfU6V4veJluZGNDkkSI4XcPIACVrjsWBx4ZSLyIvt
bXoVK1M1khqzyJePyogN727UTaSPzSf+T3KMs+2ok18Po/cjckibZDdt3R4b
lDrRZaPTON2HKR/6SJakWL+XFNoqty56OwD43DaSSMClxFBUfrFZSPw+NcvH
X60liFEm/X3FB70HYNW+gYBi5Ok8ixb5L0OERGLYCNoP5BZQoGDR91OPUojh
c0vP5eTTiY+XpHF4QyoXsnm6CQ2jjyr7g+TBofDjF8glfkM3Llyc07OjEqVs
Rbnl1QRUWCaUdFJqAgIa4MKX//aObaDNDkKrqaEfROFEKXb42Uy60kkdsV7n
OTN7RgAxy3tZ1INsiHoUTbub7obbrCUpfayPQCCd+A2Bygy9BhogAGWPzflZ
VBVAw325ZmRZ6LyIPiBRON8dGaS0s5oI9dBWhyt+XjTcgNy6q9IQEVsXpk8R
7eBUJJRlMZemqGUF0dsdm3YAXStucNcmycoAdNabYG/+FWyxBd30zKH0nlft
X+EyvkLb9VNdJ2I40ULjUlChhR0TOY1R0GiWixJqjBWxiB5pxqEepv3FNbSz
Im5nWIs7yHCdwfVOFcInyuVRUuVgEm0KzerM3mfJj5+ghemfLt+oS7bGn+ka
G29Zr2iKfGcuYr7stGWuC9zRm+FeL+sMdoo6VYBsY4Xt9HxTrTeUF90jdJmY
/bThUPCvVtjAFh2gwc4g3cN60b4j0SNC7QNJOi2Y8NSyQ5H0ZNSBijT4Xsu5
ZfHQlIfbyT2oKamK1dnxIopyVjKpO+5NNRAtZNqcl8iDD4UUtIFwZZv9TerZ
LBuNvdaz3Pv1iSqy+GH4OWdVGvVd0pnqQ1C/FGfe1BNeOv1mveUdCaRzho7w
6LfIG981FTgeoXPSJWZdFMvn6+ys+byeMyBrqTNihdOJM2P2Mq5m1Ryn1tVQ
YgnqhbWyNAYzC/detvVUbl0Ynb1/StLCFr0GOuSkxC1uHP5z2UBZ032ED0Ei
iQTB0L8SVbZDb9UypvnpR5MYXWsrA9gYbps7d2/PkZ27XEOA77lVmHO1mDYA
zIyRNrCHqqxhwRl3zVkt/vmblJcC7MGJiM7m+wv5whLgAY02hKc5cVJrB+op
1tFFFZ5vb6XpYjzjDCbc+GRFZdGLjl5LVYpBiw87d2Tk1sgQtii2BF/rf1rH
hoLGCE1P1HZDRDiQ2sF9GnPNf5WiveOrLzbImjUZKe+Ur8mjfYdwnpBgexD5
iAk/EGGsKKu2RxDhwTnHRkUyNM9ox7exgIPi30u189HU5cSuRpUCmxDU4lw5
amvO5uQnrctZxgl310gpaPbv9aDrKtV5eSChU24RecLv3YncnKSxQ6X0lUtx
sEC5FqzLviP+v5i2BMSXozHOUimw/5geopd5unP1zveB+b6JdVAxMEx0pNDY
roHfOvue/AHELpeaNnrxSud3lIRcJgyaEuToFHd5EpcOMXhT5pMB/wBWUg4I
eGGRzDETBsM1EPT7JhXQhEJ9dJQUKDyNGxD6/YicLCIKqu6c+ocDKuRcmFr1
n+2qNnuixXAl0X1LmFythrIRwKK5ABZ6npXzP++8dPVFeLvdhCR2FlQh1QfM
TCKtR3UpmuV9fXWiN1JC4Mx5uEIECoYs8u4fsHXmMnHcJcUTtDLxkxeyZmci
OHCwQOuTlgPnHg0YKxCKBYYUdXy5Zb6iCvF2k9sxDUdwovvyy+0dpPoSm1Yv
i8M3oAWk7+hQeQakkcM5PfEUHiGMsV65CeUMSb7kkkficbNYgoBYdvabaegJ
gWwolUhcR1vXIXhQZpLjrqenKeJsviFcKQhz1n3NV0O9d9a2o3mKG1cHiGzX
JVb1G7wRItc7HcUvSPP2KVczD8ihpQHVFezKlyRr34g+Ht77JMTM6jbjo8m/
rIbHcqfZ7AioGKF4a87E58MitLYczVZZjBNPDp2DxdcWgqJL/7FbBoO0OY91
ZORnmP2n+X3S7FprgNXSoUqQlIaPqr44AoWwrMdYVNLG/y7066xwsfJCqRai
YzNSCe1OvSlCmtMVR2IWTeFCCDBu3RLaXA/VVfB8reHEHgJxmYk9WEuh+5Hy
RusPcOZmwmI551ssFIjTAxWdzpJT7wIZAyW6Ft0LC9MduWEQ0Hbmh/Z07L3x
b/yxp4GzkU7Cers8QMPtZHb0ZA8A06zGCypcgnggcoNACtgAfqEay4FhXe79
6CmkNzlcmoHMQBS7EY2Uo7x0uvnhXg95d8pBJ1I/RIMjoFUJym+RwTCW5Ou0
mMuZY4MBixdjocBsb7wqIlZC5EtkALji3G2LXFPd2SnaSVKn6coTiF9Ym12y
+PrD5CHGZHJOdgugMWY/AuUbLojhnUQ3uigYSrl1Jc6ZDdFDl012BE+Y7CkJ
eWRN+T+0K6Hrx/Jois092IjnsXnzO10BFEL/ZR4QlISx5QHnxK7hZoKXvpTT
3WBxyq3sr2zL/8vvheIYO+1F7Hu1qjvEOvpHanlbjK/j5MwhIrQuxKzwIH9C
HVGQMADrV7kGlO3ohXhmNUacRpM18UTIRU8J+09yUU6rjhWNu5+oG2inuq/m
cM8vWkbRKO0dtkPzfAQhie3GU1WfjwBfRlh6CsU6Y2qahF+uT/1YInnr2yE9
uSjQflIVkkTcZuK5uPY+PbcD3YCTAAyklpy2HtKj9XwLKE89ZG3pmWOkC5ne
a7n5u22Wnk2grRwZGSa+9bUHnn8Bk5nHsi5FQE+2FExjElH4f3NuE+9Np332
yEQDb0VIrJ/eZK2QWKvAlMbsCk0e66Z2+f44XKT9lqQbmH5neji64SYnPDmK
2nsuRfC4kqC5TAyzHCKytASrGElIKhAE5ancg20xUK/Tr2//4IMfKQNx9+d3
ZNNMO1ZgWYWu11qk1uHlFB4Sd7y7T5boz1n8tkHSObC6nfjWXa54sEQkX/rG
Dl5Tu5TUOUl8ElUY453dPUjYVd+qt3CsvWQRbSXDVS7ubd8ACPks1zjvEKdN
v1uUrVKkKyNPbDKxY6rRoKn7j16Qj56/2VaIlj1pTPKYn7hMDZOzcCDu+F5V
70cvRXmuiVl/QItli5GlLuZHXHuN2gbDPggxKLkhooy7kwO/NvXmCgyzWLze
CScjncFzaqto7LTKlt6rxrIUTbtnKOHMkfh0M0kSv21rGFulV5WAiWia94cK
qSe2QPh0w6rF5aYL0Bwma1GluT8qAK543HxRLQ54Yfk7GBGt2WzE3sABGzJ4
hPYZR0jcbQUbftBcHo8wHErnZJFPJACh4BCJzzmFfPNF35inVGsOOQjSuYtH
GOzMqpanCxLC3KAL5Aekj/DOG/+V0Wz7eBu4Jm22F5649a3iw1mJbbQn/dR2
YBEJKkVmQq8JGrf5LmLc1+qCwo1XShciX49plUqqCS2KhgClPPuKWVCfMWBe
GmoUU31PRfm8wEUOZ++ha4nlcL7rCyepYmhIqhbRobqU8fu30qyn63+zdRF2
oCtIOl8Ak0biSYGRwyJ3f6jcbK1ugIGRUUb1qmqDVdR7wQkk3jzYZublp3z/
k2WnrApkcrxeVV3MlZWCo8XJQlW46j+XiyGIr5iWbvbdAl3d4hObrjKQ90eu
JY/yLLIjoZCfJnzOHFjcEE8F+sPgZXtyxyyEL2rRVYhHsomtSXO5labPqYkr
DXcaj9g0+afQhtdh3jQr69oHm5YUwRPBkyN+aZO306yOGwOMwH2Hxjyc4Jox
8jGQAne2ORXHIPGsXxhR8y27MUnoZ2A6uL6VAYd/gsrGRIVxsIwXj85pNlnu
BwfsvLBJeqaP2maM2WC/h2RzfH4FfrwPVEUSZoCedEUYM2SB0YyChlhx61rV
usmgA+ta4VPr1hZ3W/4vFd26tjkX26lGDvH5RxVMWS1twKcgF97BjLqaJDh8
ekzQwQgMwVmmB4O6MNJBvQyuEwZV/Jdm85IzPy9Moebwu1uk74bijDeO1iIT
M6QPMhwh3afZ9Y5LEuItPp6Rg2eRfJfCiNfXDUcAO2In2gMCEJ3278HT5teL
7JhmuFFyXzd4nBhgHJWTOlT3DuwOIt6q4qWY+/s0OJbUE07jnukpBZlxtAs0
+dlYvp60tKEI2mj1yYZDeePf249If1/uNklsigKZBf5Hs7vtymsDZae9976C
0xt0+d1zlIAzpwUKY1L2pSulYlYfhCfmGDrqznX4V90VIv1HvpbhDVI2/lLT
xk/FZVYxpuWsJFYPCs1+IcPIecgtnEaf3yK0ZubjHQ077H1m0iVlP9G8jIdg
G0teSdc0aexJsEcZecY+sOrf9nUPAf8QWskGvUNe+ak7jn4D40c9XUf3pS2S
XUELT+zdeswp4AMkPJTd03MYtb+6yFDW6OngBiop9Az+v+89gnPyWLWYOPeo
/5PBaRvUKJVQd/JhFMYV0o3I/7KQ5ZIcsEWT5eRri7ZYdwzeb8PLuJFw0AIK
kvIGKuZciFZJOsM+08FVL78tI7LC2D8lr9mI6ErwUzOcIdYuvgVEeqhUIDgj
eHS2TtnSjZa4JaGkmRo6O/uJ3xXGWm0JhjUYrcBb83eKL1F/vR0/8AwTs3II
4OfO06XAZHtzt4+HwvNG00X+CuGOmiksDpuQ180AFa6yVBTQ8tfBciJ7WfdU
Qcf1lToaVJL0gav0BSkZjXvdvTswiY4qZh/BayO2Yw7qMq+nUqhwy/pjURS7
3jzdzHqgHfTY9+Y8iPiaY3BS0JcTr0hqtQ03QwxQbtm6RYarp3iInSRGJHUy
Tbzbo6MEtS+0IiQe60IzDl/BV2N70gZb/4VNjXJr2XbyObHhzU9Dw5zi0SaH
I69H4SERT+8vPOhhBmLSMx06Rtp+D4pvIzMxdDjiqaUO1v4RtDkICMuRLAKK
IsgiYjbohsI3UXe7I/cxchDOmZ9OUyW27w5OnHdwn/0EpPKf5USLY9QB4GKD
pWvwoXt4h0ua8sQvhyzONmWScoDGuHsjiPd35fY0TSc3AVmNcWv0dtJDl6a7
GTnU+ye7syPnGRH9TFD0XTIcX7GJhxaK7elgdc1LFFMPCkpfckj7eHB8aR6E
kcqlvfMtNcvlZfKhYR4kZ8cfVVUlf0BCeknpzgNQ2t+tN4ljL/KPmy1bndoY
tAsRpeEM9rzNnjiKoYO1rADOyh5QxiFIgTNl61TTjPmG8AwmGbnfryHSAVf5
BK+FrpFiRDdkQ8ftb8xUU6XahEaTRtdQgigiYDuWfHjX8MnkiDq/NFsVy5EO
Q9FnOzgWChIfjUGrhb2rN0K8B34h/W4lOFJTD2+/UtGTuBSHTDd4KNaHhHH4
fkfVZivtgc66ygxgDaWD6BayqYWK3N8RD464iwzyCGyUCD4MD+/M0JC3EuQA
U2NHHzSQhafpOsiEjcJsG3pWM1lGQQLg0tmWWyFPASQrEng1qjRRjotgKkzK
tcBSiCcZNJzl3rfnz+ykzPyHoD3wJYwPfePW35yU+Prqem5pXkstqpckj1ut
2V1yCtKF32pq4Ap6Z07TUdkmtSXceOG2HAIfqZ+n52Xvq4wlQyioeEzanxgJ
CQYErNPIcVOxhjjp8hqU2DOuAQQG4/N6qccEad6Hhj4f6/DG6LE1sg09kpSi
7bfGBWITkalzr2rqWUELTmH/jrbhAlYbTOQW9ubjkO8BpTelTIcuEwTtyF4I
cpSN1TKoY9JmGgqHGaqnQNqnPhliUhdpiDjxIqtJCIXYIvaK6nKQNfdcPZm5
OE2fR9Q9FmgnhDuhkXUUZAC1xYPgVViwyylXmm10jQJ1BvcxrN9EGOtqUpQ5
vcsmVcn2rcZ3rsVKiLLEODKLYELEWnwPZ9uLc4RNl6e1UM5quY0R8tk7vn4p
tBUYAYWdV/XyDVC6XsAapuIodmAvOcPlMUCD5qtccBLYfvdQX6U+m6A1wRBA
hFWZJvAHxiiWIWHGWxIrj6fyOuTFZXGB6RHDQEddbQyA6yrkyGs5DROYoUa5
I+qgl0gFvhb/p2V6rSVxkHHAu9bqAwbu0TZ1wpJkWEUqanC002qeLOmBOc6f
P9ZIluNaAcmqU5GUtHF+OWU1VMvrp3HGzWVU3tlO+0WeHGWgvh94LBesr15J
rKJ/EzMGlAuSvu784IFRYHRrtWp5gANxMZnJG+D6pH15TH0IHBx9wQ3SNmLC
ZRUJTmDPBd9wdNwUswXoHigiiVdBF0Nai//70C3ZXM4STweM7LnnPKsp8Nyo
HH49IcAy7Xy0UBY2vU+GQvSMd13ZmUe4dMCd/w8QZuvSQ3c7MV3MgXrfVJnL
9xgVye+3RslwFOWMaZTvcI35mwhZGIbM6B8AKBC8ZaG6BrnDOnAQsqGwRmNn
vnGmNwGlTInrriZGcojv/ZvypbMNWeSH02of/RzIEo5Hze5z/KQuneV35Kh5
vbY+XgY5P9JaFgz4Zf0AiAflenHPXAWuu5z3suIUyujWcCunAf2WJaoBW8+6
X1K73SJW6mF+E3S1XYlmX8cRvVrWnVIVvFqmKwxT0PE9RMIeruODZ3OoHCA+
P9d2ceVnsY4b95GYRJaR+7ybfw/5/F7HHkbjx4sZVx3lK6xKDCwhdwkiXHIz
hj3AVRs8WgL0BTYqHMRHN7GgABlZH7sriWFNNMprJV7kAt2g8TA5HBHrJliH
8JJreitWLZswpG7HpHcqbsJKit+REzNmiIH5WHjuwQrkV3LN/grExirCOpkC
PEMLZ58YVNiOijSf18igEuaNYgmPmM74eDNhMp0gyRFAAvoCqdQxhwWsQRjQ
GMoQmLHLk0C0bgkocFg4C6320kAplg1i81yJ48ImhTdDPWRLCleys0iXc7k0
4yOVMaYCWtMjhibnGaA2/Na24H1B5k5kciJG00GF+sTuqgP6+yWDo4x7jqTu
hvPLLIkTpGzhwHeZ/h9IjckefQN3kvKPRdeB/b+KNKWkLgUrI5uLC90vrtCM
4O4Q6816ZD5hyGUKCoT1MRZPVzSYfqLNvdY8V5k0dl89po0twkABfR7B1eip
pjgcOJziHstre7R/eyFU3Mes7kzdHkFicVl81AqQtUzF5xhkrReGxyFICUdu
14XsqL7V2lROUpAyaErRqg3I3VQ5ItbBPSHxls5ZXeu9UEv1epO324hMLtIi
Bl6Y2LZpXnXZQD+TN4OhjfgLoLbQkCBO5MqZtScYQLSAdXeDyD0ymmbThiTt
QpIwOatWWhdF7XKWvc5bxCyVJp0At1rSaeCXZgP0iSlW+GR/wAMKHx7SElQC
CYry6x1sewQDcabIHqLTks7b7u9m5uoR6dfcgLnd63WHSkAXg6B2FVkYPfc+
4FLWM98NDfawhI0zyITFu22tw5aj/UklMWCjKnjFge3j/dsViYzE8lcJINL0
KOUJCbHPXvrbQ6Dr5Qb/otPOQQaiJPsfS4W8yC7PaXyMZcz6Wkb2dyGhNZLT
NgwsDV3cnLwUyB1sBshh+sC6G7qh5W6Q7RXJt8yepYEbI39sFB9Dv2Dupzr5
NCyicwim6CjWJab6kJgrHapELGEL4y/LSxM3hDBMo4TuYXwantjQ/5fw59Ji
Hsr7I/iRYqv3p0evhL17caF0M6qg8sYN0SOwNByOLDcKU//syjb1OanouC+4
GQzcbrN5HIhOQpwpb4MPNKfq95aVYVZ9KTzXgXvoWGobqyWKpUgUPjjxvcv9
RV/G3WlM3XwKiLfN4NoJCFyyXCYavA9DbefP9JJLdyjfOiIuCkcEnWfqyxjX
FDIqKI5Pi8JZtDtKSk0LScahqOG7U7kyS6CXam1TEFALFraIEGdrwEFfRsNE
8ZffadU/CpVW+yqhS5Eowxorr7lq+po5QBdiXL6T0jePAw3vPc2Txc/Enb54
GJpveY+0qf7TmP79izfuEhkEc/WdAAdwV90aW0HgynjGZRZ7T5HxaGSR5lWY
vZ6sSyQ6EHv8v+oZpj59lYWCHjisdVC7+3aq8rE4ZAAYItKwFO6LVnZU1IT4
tMMGiDS7hx6m2AM87OfiW4bCuBMFwqNeMst46W7oVj0vnJ4lVD8+XwsB2But
EL1hkXAcw4trMgDtQ5kN+oW2Qq5Vh3Qhq3Fsqe2Q0NIPsBoMaJJZyHx5vKed
ELtiBs1Oj7JR5+sDw/N4QgRHBOAuAZoaZMOJMvOmaR5Q5O1nJDyTLOgtg1vl
f5rVY+YdcmRgw6XaXMKDbU4qGUddBX4JUIz964N13eLpVf8rsZb1K42DVdL0
QXIRO0DVcqYZtWIauelnxnK39kMd4x2i/uO8Rg0e8i9l38xyjAH9fowqJp6Y
LKFISI7FqQ7gwMQvrrYE49HL/ILME6Vb/62cAopvlaXkeMTVzbjBKkgFrJlv
98P6AOpY7wQIVKp4KJ4mXVGmV8ve2q8EcPLq92hwYeZGqceJK14myRc6esFI
BvFP0tRZNVJTkJcWixD4i9JyyzpUwHGU/7mpSJQ1nGG2eykBPf9ugyDdT39Z
WFmDe6iztJI9dFqieQXVQPaXFmDoS2zrP5P4L2TJGmfggsYgaNm1qPs+ihwy
PVZ4wM+YCZAG07i9kT6mbr0XbNl9Fleyc6M8G0FPuOVZgGS//8bGK5Y9ks6j
wgTmmq1aYInakmCLz3mNobpa6YBlfSbCCo4/5s+Bv2ljIMnY/gSISoAjYSqf
57/f363fWlYX/bKvu5yf8HXbyuENtpGyBDu2z0r/Sp7HhbhOR0kxLYUnWt6A
HWTE4wffSmpZWsMnvHwQcf7fMPLLi2bW5RgEeWquGmBowCiFNlAmqCqNBt7w
MYWpGjqAC1mLyrug2FHnGCJYBs6CWq8MSMtIKBOG6t5cjYzZqkBx+5fN/9Wx
WFDs7tbvJc+qjvmLs75WNDeGyk9N2tHRe+mjgBZXbaraQ+61dnxTwoEfNlJc
lRE2rNu/uxJGatC90eOC+DcO7Q9odqUG4qqmzEVsK3WVYfJ2Yzv0Ffuo6Hw9
SoX7qUbpbbO2ubV/iGUeFJ1sQRyS1x+qPCGWLz99A0QUT7hdRor2XRVfcd6e
vjM2oqJsDV/u0Du1jfLFrQe7V2Lca1fiUc7wAMy0QL4Wbrs5wAaH45YKj853
hBENkJyjguCHCFnciPERelG2mvFLxXhm8nqlQ+GSHTGPJNrBMc6Mo/aMNJQc
oXq5FpvephjpJaz6pISU5346bG5KK8GHZpU6gV/aEy0Mmm5yY8V50Pz2hOfg
6BVJs6QHk9wDU78aPndxO17VVAIUkSePa6yQfDeqscz2XMSmrOV3NE8LFzdA
oQumcb7/5k3liDPNKGrFEcfevr2nLxHgx1Gw9D3hsmAthqexaNxX7yzKw+n9
P8zJhc8g1zZlw4E7kann/ams6JPOysRVkoOGaGFiEbD10Qeg+LY3ibWxgibI
5Zd/mO62LtziQGBiT8+xYZrUoQNIHp24dbH/L/SY2Yqmgk9UK0NcoR7IQnSq
6Ki0QyMhdkJC/E1n0lRqYoyLAR7XYtx9nW08QfQCTqzov+uuWsUjaWKCcuo3
STmD9W0vf07K6HKCzbk23AVo67m4i+pPK9iAWU3/H7tPmMgVKGaeKDN7DDLr
nbNNGaPWN9xTFz5gvHDlBn6a0VKx4GWmxKhcoxYWTvX5Ta3EtXofsNZxtB5v
k61973ciTWIT8YwtJ3sUm0V99pn103Q2qSRlss7RVyAWt3lmfxYycDXFLpcR
KDspA2UEKqoupKBx3UIv1h3d1GL75x7ag2LcTIUovmLDFt00/RAfe6DrrEXI
WZ613ckFM0C4K72B9txhDek7fXhyRQB0Hqp1hiAe75SOQG3DId1SBvtlwX/r
y4g2e5JSgZtCcWoV/jYz0jczn0OQeH4u5oxcc8A+14wpi04Gq4/Bc8qTRNDL
QpaKPzkbUJJ6Hghw2uDPUHj+DVpupTvDD+5bYPuDlEpIgJ6Ko8ksoeG9bkYE
wUqhjGmZGOMxIazrZwOoNw2Af/DwQu9j7psiTHsM1uFcbikEvOPWOhP1f4WE
xoyehKp3qci52AyWwkWpxOxC7Ek54IjIlWdnG+nX0Gfd/47VXWW5AVT33INw
4Je89Yaxxp05Io7TVouhQWKLSrFWHWmc4Oru/5L3S90VWQi5zAL0LPodgE7v
iBDWHCmeFLyMQwi8iH9XGXtp3wfGUnKyHW63BHrbiS6BSIxIu5ZOfa41Sa+e
FBtkpy/JBKbwxYZKQ3J1F4KSEe6jAYRJltbBUguLqACnb2BQm2sueJL+uXqQ
xjnQziqJqYwiT8vuaJYW6Ct2gsNVhUaAz0WpBoAtOmJeF0YAGuHWyjiWRimv
JW8r6QfQMm3EFr228SIxslpmElEu/x75Un3xobO1geG3Id0yfSxw36HsQ5ec
9DPb4FETJlewsmqCysNLOIhcv+sl730xNUPcpcldbSxKp6cdendJOtT8ZTjy
j1DkMdrzR9SzdWsanJ9sJItgs8tkOOfhoXGjiPJ2QWuO+G0fzDlN86ZrUOy3
FvV1s4TYpvogg5E2Rdk1LL+LRzu2OtasRDKDJVoFfrQDuCY7LtqfGXVRCepI
brgLwGvWNTiJzAYSTjueSY1Nlh1PBW3A7jtJRRtR2jeNBawv/TZiwSJ9zLE8
hNr5UnTD+pR2vjWAXCyrumZP3YSo/PHuS2xetAXH0Ir8L3obYW1GY95Ifexr
vHq3aA1TVZrYgbh8kywIKmwR7V6eMnmH1tLBDcrkq2IDRUXeO88u2mviiSC8
1ajewUBFtJrkMzHZYYWaUuiyBXPr+q469rM0KWQ3gYZt8HlUFStWefVFkPtm
TYZP6tX8PnBYWBCAHK+7/py7A0VCi5Qk40p8nbF894GijVivvKM9FoOnjDOu
jfp6eBVZXrAtY+BA6pJkoHEwNtPMdwdBESmSQZGvTb7M8Vsm7+pgDBdBK2h/
Gy/oCDLEhP00Yl+UTeYnUrO+G1b2MxufYKHHK/sXBgooIvRxlhdhONHOADMj
emoc6mto7NMtBZmlh+YV8opOIyT++RDGmlZ63p57HvAMg1Ix8fJv2ij2McMk
T1c/jfJFetzVxrDw79NJ2RaPqSwLtxvLP1GFl2xW3YUD3Ubl81ES0btiFGvB
LDwSIBcNqam/c/RcHySzGsDGRLmkWQWAkLPo7A7FKZgL5iP0AfIrixK4EwMX
SPOIIXj7uAYbn2qmYstFn7RazN6qwLKU78nZw1KizU8Gy0RGavPI+aayP7dA
htDs6zklvS7RhWa/qm4OjufrPAS7/Ph/9x+avY2mvwam+sMcMjxl51v6o79j
ujaEGRrWsL/L2kDUBzT+J77B4hSRnK59+iHA00x+oecgXMltBp9somVG2LUG
ENejlJojai7OeYdOKjlA4kElMxHmZefsQbvB3XSsDrHp04p39F2V5K5PeQJa
WIQmKToofpESJJgxHL51xWxIs8CkLyz2Put+0P81sdm6GF4g9yoifpJyYN2x
560Vs6biZKN9lhCYG+rBJpcrChiGYmyQKYQPVn9nZBmHamxaJroqiAfb+YiN
jaX4EWrJBNshZ6HUqvMikmCVcHPwnXzqRmjLiDw4O8pjLLJktqi1iImn8S+H
cHaFpLmzvFvai0QHBGsEPw5wb9OAs6HwsBcDCxR0kV9L557eTErbwrf+3cnr
xwXD1R3ZLZ42jo0aF0EvpxpuXlbPeyIw3nzuyajlxANKUvdsYiPP9ezqtF2X
n5fQ/x53CcGL2K1vMAfPn94Vnzns8VdhDOzL6O6h90T3gsk1bLiXIvybugtn
SIqIgUe6UY0m+vJaw4MwZ3Wvq62H1Mr01t03D520RlMWAnlyygPPZ09mGimo
aKQ08ePcAe0lUc1idgB0K1L5hiQBKDUr42V+gDdghOH/IPTNh6pUfDzABPQ7
sBMEmAPcd2FIqwFEvftgXogK+tszGAj5LqY2+MxPhE2vZDFpRMgctI8yo/Oy
xB8EVdNJij4uAnSRz8K7UWJ+O+2WMFzjpFZCqyHS3j8g7+dFrMs9H/9Omjr2
HdXD1iH27ioR/yslO18yJ27kWqEFYACUNKoehk07s6Z+GEjokwxkgJZYhUv0
akBHkAODRhEjAex5eY/crQtfk5HDMSp/YcdWMtY7wKGEASB6eOLEF245H4An
fdGrKW0JI4JwB3+SUCaZsAOTePg/JbqA4YPrRXoxqX7n+tjZu5Nj2icku4z3
b1+n16D1bQXfQUPlVbQB4PT7Qef9fQBX9zRXtAahgXFFjbrnS/28DidmQasb
pEN2+vMHJxE22rv7pNU8JbuSyA1JuIriVuofJj9FN1ewa7QpDhsIzB2c0tq/
6FyrcQ9Yso/riFuFTq2E2DPEH8V0PaEMPD5eLLy64KM8XbMpy3AXyd48qIUe
OsNpJZQJmu/YWsgWzy5o4bzgngwvcl24bIxY4jtqsKWaiPALlanFaxGva1DR
Vg4WeREEXkVkeqpHGHzqmoaAWBhIorMfZJMuYbpYt1C1KjX1RgtS5ceYSMQ5
3XeYFzuNM23wpmWmBS218u/AkJEVBzYfgzXlDMs9rYlfgtGrJcoMu/Pd2GOv
lNsjA/jm+z0h7fwGG8CFgsZEd0tTM3btqbadi17n0o8eYp6wsOEUtvepzSR0
ogYPilPdcIlPTN0rr3yZ8evRU+mf2St7DbC9LMaeEGh1cxldWj+S8wFj75Ti
5mBwYPVixAt6qX1wYx/xC/Jgw6SGfgNlKBrPv6xfw4Et2z7P2g4cRKhk8lhi
EMcukIMZUHWlNg6Glof8oAL5cQDQs+auRMUtZo8AeUQ9YEscfBgFmextdDSC
S77RYWvmtDhOZntdUCvBhblbqdTS6/1K6EnPMNO+YM+ltsNUOlk1QOES6cN/
DEnS3QMASZwlNFT8USMik/l1tJ8ivO3qmRtGb07krg44NHazsSFoD3KEicd7
X4TbrZT6xR5Mu5H3BIMyJq++TQwmhJWp+9lc9Nl4BIuDBgx6ePGTjXS2hq5x
3m0BeHpbF455ptBqiDaAa+KufC9WRp5XyIeEEjOVY/TH2yWt0Sz7R2fSE60r
HI8nTE+8s39i31R5sMp+1OV6hshte81elU6wsI9viT09rzuCR98nAw3m+K/Z
eIqanPaZGV6Z9xzvxlWMjVBnahdH+gmupkCmk2Oy84JgPX+6dAP+cw+qC4V/
ehwWXdboc2WDFVJ3HFPzlprsQmKsEV5ULyWbYWQhaj3uczq5bJhUsnDMJ+pV
gfeVacSg5/NDZPL/wasGNWDCKlima6a4Wc9K0q/lRt7OoEBkVUvLTzBY9zc+
4Fxv4Lpze+omJEGGoqQIVWccD8JpIz+lmro+qj++Vrg/i7Nyom7wkJ550hzZ
/NE95CWqPUG/vhmGnAIewcWvPoupzy26lG0DHPYgCjhvaXf9V5XI9/GVM2Sk
AyHJs/ntEcGg7skhDLNQWfZjtM2Pu5a8WFg1j+5EedKxHeMnAsVM4unGqrtD
X8XAnGn4lyBDoEtMNab0FUUxDbZaIn/s5eq6Dbm6UBlvNNjqgXxuxx1Em0Ai
OZr/oA657MGB5p8ASngQ1Tq/L0RG9vAKOi12bHrHgn0a/o87ZZXAO6SmICIm
RjoTHRNQQUEwKAW09HKMoUYGvLPl6/CpNzne/liZRpOXDLutm0nznKYgGQPh
17EngxYQnhPowgkS0CZht8d4Ms0j4mzSsSe0VnS2c5PkS8VtREkCosMyiqgT
mpA3VLowVE+RkkfCa0JCFUjDVV7Cclfmft7LfzunYB+S/gq10kKi8tUqIRes
PaJ7RBj+TvGViW0GjBOPzpKDwFmsGivkfgLYcjLnGwtqEpn8zUxWjVQTMzpW
rP0RiMY/vgAdKX0ahSCvQn9/xQuAnMjlD5Z5T8j8+p0V2Tx73mg45gzXhfh/
Q2eclZju93UX4K2CVSju9JCJZc9ZBnGIeJ83RdEHkN+HZhFP+uGNlJ15Wofo
Qvh3oKRaFgi5o+a9+rt+TbXLIVMJqpXOhgeziThB8wt0OzPXU13KfFQbYcD1
650a8WnIkNoMMSkms1X163s2k0JSi0ORUP816lj/9EltKB/j0I604GFBkQcY
wMcxMfWQCydVy1bL3XWlxnfyqMjMIq5YffnAKTU96Zu469nUzbe47ZzARIGQ
t74x3Ef7X1TwEQQHBwyRz85ds7ZsaIzGeRQXJe8IHMfgyHAMO8XurUY58iTk
CdR2vZoSN4bOaO4KlI7pXfGhYHVO2JE03YH69gDM21DjW/xublyULZDPxITP
nRB1HBGICtVnW2z43V+Uh4guhrGjce7Ir41yKCfVITYwEixe9dFrtanBGFVw
X8s8u7rBu43pEep/fh3JEAI+xREkw+I2S+6Ew95L3CJZ00EX1tbLwUB7IUhP
OMm6GJ3gvRWEB1H9HwYZ0ogVW8VAPGfA4GWDwD4FCXOA2xqPVymMUoLX9Vqx
OwoBXe0tRzHSx50SgbvDXVftkQ3NRcPBR0yeZUTXv2vODcaTXTxW5Y7D5WL6
mIz361MdnrzjqDQLTQHcI/1V9slmNA4QN4f98JCORZIXm0faL+IZSnQUqxpL
IG4415c7hH9TDmFylk+U4EkZ8iy36GtNQWKGq/nNtCZWwYRDTfPSX4bhgs7/
lwsjANm4H3Qay9NkVoYQ0ngQeUVgURgpXb+ODGE1F45f+RTTqfiXZypWLAYq
Ll2+bxjZJpmhhx69HwhFUca04sakCf74TPa1knaib5wlBEPBsdX5wc/rxVV8
j8H0w3isuTVaXxM3oxt7hBAu668fb83s0bHHO1Ia+hXoJri8upN83B0aL+LO
jCGurpdwQ//PU9uJUbv/aaRlPx9BvBjPpFIKeVs054dSFDhUjjap6LqO++Fv
cAeTwfFIaTgLgF1ToPMzqDhynbNnBgmXKaqIF3NIIbbLXs1kxtTqfpaLt2GF
8Alxb2JIVIoDhsVuOCtApTKH+vcNV27yEssgGg6/JWRtGut54e0LGNqAFjwy
zjl1PN6m8LBD2s6+dZT7HbC74FtIuZeh8s6yF+3EH1p/vhbVnKSimBI7hW1c
Qi0LSrOIXKZ4ZbwMwIoza/DulCpvFzXXjsiO4Hyi00H6oSLzePdVCz2c2+wA
gHeXp4WM+2r+6ISpmat+vscX3tFRwOred3dVtcfy9qLdEZpglqX5bTKoUhfO
5Qh3in9K1ZQa6bmadHEN0ZasB6qPzdYWH5QpqX6yGO3Uyiz021FsrtgH8mzy
TXaYsdW0Cw/XNarueowZfsnLeABCJ9uE3/h4E7PUCYk45bYytbRbUFusSI/z
druJlKfbOA0jhcAQbPpHQd7qORi+YmVl7JIfL+rIUbZP1fXc6uoVnP00D1er
530Z3WPQdGf7aksPTlzV2jf7he093o06Rd5ajSlQNkvlR4hoWIF3mRnkeCB1
FAzOR27jJU5kNPWvprpyZe0XQNDpRdM5QoOEBANATnxeNvhQ51SkLVQQN8BH
AdcymNNEHI2PQhjuu+rc9S9AOwPBUwfI8QnzERhbKhi/KE5msZoDE4ANNPvG
RqVsd4RXAf2dzS1P8c5u2LRgE0ItVOc/+qbLrCptbczpj35A/8hBoJSkVvkh
7sMZhDUBFb7sQ4vPEvUrQ7T7x6rpkwCiCIBii1GWCupC+dKdHWSCNCiELLpF
0L0v/uKoH7pbENvqz5kFtXVUIUVmE/WCSpUEYHkO4kmAE8D2kJU0JXLaUEvr
1cuxtyBTRXrMUBuHBUWw//O8AltWT9EcQqRhXalLBNU/FaOJ5VnYX10Y9nUg
AOjOmyxaUrAEFJ0qoJKF5nkGXiICCWEnSjljuU38aS06i1B8E+Nzkf3dNpSF
ltjnEqcFL989nFC811k31fIpvy1fz1kJehycKZF7l50FTJOf3BUqThD3eoX2
cmMLGjzWLXgg8E17J3y3No1VO5+DZkkGw/ZhtTt1IE2hpiTE+1RS9EZG4e8u
yUjpqRIxnLTea/lGgemjl9v9zAH0M/OQGp84HNaHzepilBJWQsjpKRdfZqf2
uzDKXf2cSDId6BXWRMhh+XYa3Kg/JT3gAcjX0aaulMiy6zvlFj3BsVIMAIwz
Najwfr2JLyeTkb6JCwS1m4xp0Vh3SibN/tbU464ZX8rmytJTMt4uWmV7Z8Hy
gW87PjIu6Wg0AOmd6NjmXo91t5+G1N8W8AmLdzKJYgvZem0C60KAoB9RHFo8
VTFoZHBgMfVkIpgIk3GgKIzQnH8J78u0+KQPECeRLhmu+MV/KlEu9ljES48N
w6MoPKFxXRMi3h11eLuWv3ZK+bNUuhznFoMyCnMJ8W0czf1lWYHcDHTta777
FgiWgHwQC8jBSgjhfqIXWYIpJP2pWaMmM/Jg1B6WSHsU6tpoxQLrElsh0Zhv
DKmWYAVJnfqH6V3qRnOW6Ugz6ZjTxaVPOmCgcrI6e9pgq70zAFMdq3DeZ1Gk
YMT4qs5IHcMGBH7Ewx7WtZd58Xe9X3myIJ6F02ziuy2Y9hZf99ISbRYIX749
sDl9HDKoGs5Y55UG2yzihdP2n+YvNXNTLKHnpPG9zEmNs4iUKbndheRAUeP9
jx1jPsuD6XOqNDH46ZbCcQSiiQU75Ld+bxL40eswDgLmvree5iii5L4FuXFE
Hs6K0BB8UILWMVGuvWDaZlWvRQNZtKckcW3hxT3HFYYZSp6oos4258vjNLzQ
eVKmLhXESTtc7T3wVFoz8QBsAllKXvMjow3ZuW0ri+syD1RO3xDS5UDAZNGp
3qWGYIwFVr52cY6ja+0vnZPYnuwUnmXOf6XSY6UYhkkUD5+6x5etNH2imzP8
lpgJJETHMsRGrqCd1VjSwUQ0Aj2yzMSFeXf1Y2F0GCvqNkNOxQoJtpV/SsZ9
UGgQX0IYi7+bdekN+n27H5ji7j/6QpSsOt0xTSgK2dR3SXNUJer8pgkKkqI+
GgnGwN3q+Mqnv+Lem9r5xi+um3/NX1scU88I5vYl1H+U30PC808y0+0qSpIF
V3shKTvQ/ezBhzIVvohLVEytHEs6d7C3uioP4ZFX9WsOATSWujxF3ZUDQ232
6fRrf5opH7gLV3+xU8H0uIlvmpqWvRbbUNmqb9Ga2+o6RZkMaxyCTJLzwWfA
GjNU3cVm7vSQ8C8VtDQbo/QRxyG1IZeBalBtMxGqfiD0ZPFEm8EzAVAZ5ZJj
3TmPkPCt3UlKxQXc2SZp6sGFW1JmizW5ng9dINPCi9/8vxGv373qLT+gW5j+
0WY8hjiS8ek8Dhwz52wnbs3ZIkZ0SqmBKjR0B+rky1yWE0k4at7v45nVOfzr
eG0lSAB2cIOWlFhYRmkUsnQvtSP/M0a8s04PUbJ5BfrdaLAgamYU4rKOouXA
Hz+9jpBo8TG8ufBmrbvM4qxAkFvpp2D8YwLgFsGWK4FYpZXatOWzoRnCyW1L
BGnzZr/xtM0a/krrWw1aDfaw1iMdjKhDgny1FCph1urfuOrAs6PswREGV+Zg
9bjqIY/1dOLLbFfAiyR1cR7V8JoV2yDQogvMYQL2abBe9fGXB7LQMCgWzd7J
q8pLmvFjiowmxHrxKP3xCOdROpcLPWAlDabpwEfeZMN6mQ4kvcXmkD7qGswk
gXuIdFiWzY/W/ojeo17B1AiG3L0lZ/0eZZWQw5MqhQRV/4sstxqofK1BgPW1
5kouwb07Up6Re9pjqiJtQC/TiEMmYwJcUvq/D2rQP777McOBx6LNMad8m21C
u4nOSEMocmBy+jpUSlSnHQCkGTBcEDdJxaImZEOPDeezzQixO7WgQcvYqEmt
S0ISKnrGEyLw+KbzIXSMg5/wxDmKIRhZd1N2cgf0nAmQE9K2pWdz3IsVdSm3
wibTeQD0U8GG/K9mfsXr4rMvhkueOVCjWu5p7sLA6E0g0sSVsfBmNH4WFE4O
k3jT7K/2uQ6uq5BuDcdYVfKzpPfNryKfbOY9nBHtULwWJ6rajfpW80MSTJwU
/o16m5zqbQeV+3As6qGItjFI0lmnPEyy230r6lb+hge0iMGuAjctJtFg66/c
nKTG4O9JCWefok4yFENUn9miVmSp7dP7jrAG/RcuIcn+m4Fxn8t8olvOhW4Q
zqH98no8ZZW/8ebBWoylQb8KO2r1xWGlv03L0UqJy2X5epKCnLjzJq9ix5iu
BCt/siumce2hBxrDnsBmpEukxexOq7ng640j1skn+FWHa9FsLrI2UW6XTqNO
dvEE4wvpn6OPPBMQbUXd5+a0HBvF3Sd4UdCKEv9M4o8B32hVgMt9tf/WYKIp
gV+9nP+u6OZ6w2djXHAZ7iMmS9qrgVPFyK3mpqqnHNPYzBRScFpRdNrYbXhA
xPINHu9DNqSoCXs78BC5AizIn/Y82TNcJxsr/RO/xwphx3cZlNYecSXUDXvL
h2U0uTiZf3F3e/BX8mIKj0JdoXAJ3YeYmUy1MKCExxBRn1FLGiSOlMGLsZRt
kHty9Ee/CI7y7p/mnIaoAIRGHMUBtLblXi+0EdWFfFEhXP/lvQLgpTB1V2vg
yfjOoqfK7pz2BeV8Juv+JBVQzS6Ix6fcw25YEZL6quwDHaH47M3kFBWH+6kf
Kb7d+mDvknNxGoQHvw0C48YfI6mR+7zs+uPzeWEx9E30qYc4dDs2eRYwmS6f
IItP5QiDrq7JfK7fgjz7OlHPLWJJ2hr4HIntoV3kRh5SoEYYZMnKLMfQtXBa
7QMtKo6eCH6sDScQqOJYD7m9XHGpCwmcPqXkI5CvC+98ciOM4uYoc2t7IovJ
VELS1lBTCfrZKW2b4mRl/FxfueS0xhCRJX+jzTcs7ROgIL7dVEh6KD+rOn+2
+IgRgpQ29LFd7d2ddUD2T1EijU//Iw50afeWeuoTfW79FEuJL/Eo63h0GORy
/S/GaBfwBP0krNHim4iv/1on6Z7jEzgizigQMkTg1iebNyGRyBuCF7YqdJve
mfWD8ja+FEnjKE2rNrXhE/Mtp5fa+sRKupC0mK4eScqwYI4fxiIExw9izu/9
bhXc8AKah17lyhB7laOKD3ER2ME5UBcMAiqoEfWDnvdaQLjBG03HC7T0EAWX
Gr2gxrQM4eD0JS8jHLyHXT1fHrBJpUslYQX+8U61xxDS99W5GhRl5TqQUwdb
pPFn7RJVpTMQtiXXz9S5Fg83Zsi4RT8TT++tNc92bMTX1iHP9jXzEHOwhW3V
aR6En5JbcS+jStEuij75P2HCgyiuJhjLLPtwwBdg+b8lB1Tr1tnOf4aoMxqi
HDcp0JcJGXJuC+J5vJiwgT0oVt6df7cbhzTQ4x57Y5ZYraEZcMBbL1LrHjK5
M0hMpVP8+1Ejz8l1GjxlCAZR1+XZ2C/1RsM4h+hhJ+7LwL6HdInHZcfQZxTB
E3P5haIA73f8Y5wXZ+JnoaVr2LRu//vHU9JGWxtuzERYW0Lkytx/GpwH8x0A
gr25PvSQCPDZ9qq4D5yZnx1d7frXy3q0M/fZSTYHbrWjNgyso8GW+xhHUpvX
GRivtPSl34FkStl42m1hN8xPIOWZFKr+ZulsVVXZ3ni5Wcqdgrpn+ve4NlQf
9jeLei/Dt6bGX+8oIqtPgV3g3j0nosuKBz7HdqSVF4bbhJD/MfmbYsfXc3iT
CZK+fX29I8Ly6WRaNCb/ftrqCBSKnu6bRl4HmGqt4M1cfoXe242XxBVuxuM5
QfVnxHCZDMHaikM1RxBvLa5EZR+gS0bXNddc+3xafxNe0ZuDpBfYi4UDcZQm
lQnHSSvnm9ogAZU6zr8Ertu3/S9yVKve9m0vU/KEPx0vEBBJ0xstTO6oxe37
fNamFR4s9fWYNzAkHszSQKQYBmTFzmNFU3vIT+Ei6zSmPFebZIjh4BErZGkj
ga6yoyPWWanEaxwX8gIC4lNWzgXdloEmXF9SK9S35SkK+OFc0m5FMO0/c18g
PSn27OfUP1bBzWZVABIwWHBnHxlhpTsZa88eZvWof9/PWN46AiNLIKM+d2Q/
jzTqqMa6wqnG3PrgCB8/M1pe0ebmPipovZ8OP6Gm4yypNO+WvWn/D/yt2JD6
9H3Xk99Kqf50DqmSCafTux0/c9tcyyowVRCnBSNsxVeGyV4gNlGwMyU7FdZR
M14KCPSJXOUk+RDIWIsxN9WiwLOTF+ANTVjGYtitYUB69ZX+HX+D0qmpCznh
xePYVxEkuvr0peFSlyjYGFLcy+/pkrkRLOX43OTPLGAeaVr9CLcJf8AuMTC3
xT6fhh4OCklV9m7bsLvETDCGH4G9kb/J24UWNN14u0K7Fh9MUxkPs4CPl55+
eldRxJX/PhynP0Ad/eqRvTdxa2ln/7ZBgXbmDO38VmbbeGGvUDMTO601mEVR
vYnINoIybvBMTVKkekqGupKe2OrzUZaCtwB8/VyPorhoUyRClsvKz/f/Wl/I
iHGh41tl+E4vlsPvqofIA+3nwD9bqDDAtV6N6hqfrgWz4Lq2sHSpIdpJwi43
+BirfoDvebPVD74L3LWnfHmQbeuGC07qJABL9V9yBMOUyVX9s6eB9q78ddB5
gs8hRlk8LRZJZL+C5PRSy7clHg0odNB6++cn0yC0Bgpwkk7vhJYBpN/xsFgL
u/mQIGmAFmFvvEMQeR5gXCBeV24XRdfGCa2lErQZuoVz9lBunrz1HJ5a9g/7
yHj7L1t0jz+vYiaBcj90I8OorcPgphO0ym4snr0Z2rwdPzu47+OSmf2ey3xW
tpMZLYshOgeQl3ts9dkFN/KEWMIWJcPBxczlNMZVh9/SsTSO5YM2C3heaZ0r
XW9BpjCx/GlXuu7KsQzjch9xOeiHECxjKtKM9Fgz85YM2Qi2nwEwBzWgW1fx
DfZnNg/AUKra36Pjsq+aW9zcSXUtaP12PwB9TeAuWmNsVW0/womQN9OggtKo
1YnkKwEM6y5rtS6md3rXndMCMm6O0OhV90+f3aLavAJq5K6Tw0SLy2RCsVNm
QrcUPzSBxuuxSjg5RgA/yBFay9czrYbEWRpAxBh0CFAivw+c0cEs4qUTa8eG
nSJflZwtnOereg3SoNBNKHeyHtH+qbuF4xgvgCj21/cXJC3wVrKOH0ecxTfM
XPch2xqsWvId+ZWjxnKiJkdNlAB9a077wIIVgmnuD/V8UzF+kd2LFGmhmPBC
pNEF3RsWeIj+m6at45a65UmfRXjIE5ju1DAQznxc00UokLnkHIqFm/pXAr7X
jNMyyD+baZzddOVoSwdzYQjeoi94D7aKWLSJl1Pjziw1IVXCIEa0U8L6m05C
UYdMhO0DyDbgKEI9e7dUIpIJxTWR9JG1+9LbhB7GuDacLitXeme9dFbTwkSF
0fO5i2733VdADE5bh5nNhbLqmmApMjSuKNGomCa2a3W6IVGQm2ffaCVMQHCV
39XpsVg1QSZcR8YBqpzIjfdYSInZSiRvPThwUxPZQE6m9CaOeC7SPN4gqUIU
mR4tjXkABuqfQegQbIsHyEgpWIUDgHejp2tTPJ2tPwODXsLXq7tx6649MSlw
TW3rjxuLZzInk/S2Fh+klNos/UL/+N9JkHL5ZLKZRKK7ZaXZr4ZA7XXA3TvI
CYjbnj/OYQRr6ba7f5ve6ZIvtpyZL3OeYqe/eSsfojSr7bbVaLinwhiChcNY
WB3vvhtESl88HNQV2/NwqXOoI4+0YkatHXG5K7kflXNmDBa9bxNgeGr+o5ib
GbjpKQF26Na6r0WZkXt4ssHvel8qmw2W8a5i+cIZJGwhv0UVkshSdnmsqhHJ
1vXLYvQG/F5bH5h7S9Foijl8+Zcbpe7ZpLrEqIXWoWCeizntG+dmhY80P3xy
DP7jv+Z9FMkHzA0Ze/nwa+wEsnchUXQgmGeJdSl/kRCtJDoJTSpoQBC03VJb
5ini5pWtRu7Sb5WyAWstWnKxRduf/kmrFVH/NBAtC17jdCvLfnldh0uLArar
RdWx1Mebqn+JP/GSBb2rtaka/lFxktefg0fMWIbQOp/jZ8ea/XrrG2qKXG9a
Z1EG/GtiJImTGm0+yTEjvhacz2SAs+oQgNvZTJlwUs8rhMEVi5I4SiU5JsWj
p99cjGF2ctQdpv9w+EbU0bEJBGkt0voy8vdTXiUpg3H/1Id4pPdxdRHl7WNT
uOSiUeoPR6zAli7EZfNSVTRjiy3eAcPUjkBMe0GLuaLgp5zIETTLoPdQzXD5
HlBcBrZRpJpkuMQl7pgVq0kYk72kNWJaCQPr2pdMjgxBj1g9aLeXksz8Ochi
AbupEAjtb0NJ/DioPlpO6Yb5yOPR2ZeEkVmS/7LDzLV4CT+NanoHcBX2+ICd
3O0MkusIoCHHSEEnr20GqS4Nn7JZ6/NOQ4Wkd7foysrqpKvTgEcK0SD1nlPm
FzCyAwbgL8NHNKUUvQU/oyAtvNPdjMc7MD7hfM4cBmfSXZ7TzfxjchWsNQZP
aVHtoQorinJpWcCf1tp/4yjpPPT2wU8wW4E5ruTUeQNjFbMVKPJXH+CwNbiK
2xPf3OvZJkcHrzS3ZIEn0wPddCxyzV2kNts/S8+G9liVzU1cwTqM+8A915Ja
Hs9GWTmtynmMJmjWkGfB3aCwRhfeVTExyAVLKoLuI7lJZLkf4o4BHX0d2+2K
Lgvv96sRiJhA5/dIUSQR0u2WQY5NzNLOODw8C++7bFeL60C2diGCYepJrXSe
XOJyZZUzcRLiUcqkoKG12oeaQWgOWpOMsP4qRoxLg8avfI771jGZd/S0MjsO
2PN3EIOhLk6aDoiCbwN5Or3dyGQKjPpesSJZUFtfpK7vFK5e5YUUk4axUtUC
atuk9CK9Ptoy9gFQkH/G3wtydKiXx+uB0GEFHhrozD9XzKMYdlyZrv21pDf0
qonvKhCrvSX+pFha8zv3yMoXTWheCg5lyZvq6E96cfD7kJgZ2LsWLSp3NPZj
C6yZKv6rAblhXSDR66lBZChu1Zn0zsGEjWbi+HJr3WDjy0Hs5zOHKxm8ne3j
bBdM4j+rJaUxdCgTnuSYHcLrKMnj8PxmliH9MTOKVFkfnBrdvqhGD4Slt5X+
/jZsuXMSqrhBGBeOyBryTVXaawYnXhg0xvcwGj1MgV6TbndgsaFD3ikQfvDV
J/lBvmhjCTpU4XT+IHTZnH36DFGEf30LJaVsHOonKqtQYCGfJHslcvBV3RVF
AsEvkqVfFeKqW/bTyWiMd0cYI9SQlkXm7JaP7KkfLwZ9TrG1bujmU7r2oRLC
lyKv5qNLyN9MCq/M1JQU4v3rseqz2pdUq49l8NEpJw7SemT5ksE812yiUc5B
bk39wiUPx4yb7kII+v2WdPvWnHGbjLPBblnC022VvubJOWDdXKvzB6FVyf4o
tuodin8GUUAztGtLrmnlZde0aMu0De+hUekngYVWmI+yUWnRwqq4SiQn667V
trG0LneoTvQUlxa2LJfiPgq5xantZIkVrF5VjsAC9Txg+zOts5qK7pJJBS59
aKlsKgwBo4X3vgJmVZ88f954l0jmkP8Ar7RtGalyo1ICMGTuw1T6zFm2vo6n
ed5d+ShG0ioyCOSx0CUMdpDtXlDmf979S3lsivJVSJcM4KEBeolSfMaKxNda
p5Ox7bJcayHRjlgKqa3zqKAyJGTihgO2TZN0QGpRZOaOtkPt9Kmqil0kaUWN
13ApiVqAiLps+yQOo+02ilCaei6PJIM4c0apUHjG2FeH9vp/UuFjeWGOmF39
IV1genFwXJd8tZ+MS19QP69Qq6PUcV7prbtMHqU1fHD3XFdPZ356Ebi+Nr77
U4K1J7AypiTS7XB6AnmxPx1vyM7MKrqAxRKtNR4ipgMnuW9GSGIqeHb3XkVI
Kfz72OC9kgX5jbtC6EUKy9ZTPU04L24GoALbQloljoSvxq6bkB9vIwD10nVJ
kk4MLiAxs2+adE7toyZ4Fn+iM4Vh0sjf5hSPA84Pu5UOIDNrMnMOXD3wzOrF
xIcxuexnUJontOll54e4dr1Gi7ctRhl65qFpAPcx38tr+6FIpmj/8dnljI7s
HC347EPzEsUjr0uNYesYiLuLxZTtDlrh9s/+UBCybzlrLrWUpaJALiv+zCvI
56aAlnmk7Tq6kA+JXXT+Z7VScS685HCoipUEJobCZT8a7rgzp/pAEeimWETn
pN1WOPI318GA2O+6aqFhuP9JNiQRl1bMe/7s2bR63mi1q6fkVWDxKbb187q2
gWfcqMRUp39ot4M+X92dfNltvj0C9zGcG8h8PwqnPqBDarCh2ajAysp95hqt
vmB139tl7lehiin8/BlzLJ3eumfb9b2tO1kJOWcN7oDEXQMHMMKXTXI2mqab
y7PZx/KCtnB72Gf9V0ZN79y7cnAXuMzcUlzHj/BZErZPD2vWAE2G2azfwpFD
RSvtQFDMCkCfXugqzNQEwddfcLK+6DgyAY+6dYPe273PfcBU7j+74Fgbf1IL
IsY/WjkzhHvrHMmdaR2VD48Zz8cqQEEL5DnejKzL55vLqL4DfYmF3tSzLYzw
U5As5y3qs1Z1MoVmDBDNZWkwb7xPxIN/Aauyri3Czg4t4ikby0MdTHNm5FDn
+FVpS4vHIuftEtdL8cmwQkYcHEncN+KdSJu7vwH5gkP4lnNZ3NGIAi8JJGWN
gcffW8G5j0glzYKnDTEVLQov34INSkiJoNFHNqj3Hfupb3o2aPL7HKKpf1NV
aTtBSzDNw5UEav714UvSoQEM3Rf5+JBWuOO/I8J7PD7VGve8AdznFZQKxDxc
PohGP0Z3q5YCLM9wnN5orCNQCtag6hdEAaA1mF5cTM93/B/1WpnNit6/RQm+
Cqjlqu+eTjJTCxA6wSjbKZxNpVdyFz5f6HLh7StxSj04bNQXn/X5lX3As0GM
ZNFSdD59caYtAlcUUdFHYMwd3NLtR5Zf0YdLOWYVdyG4nHFOAAJntdxp0J+a
CzbkR9359JkKuBJCSZcyN+C+fxYjXCOuucQtPMB2DUyWwsRGTjbMzlXHPHLe
Y3O55JqVZpK7F0c/8vaJs5sUMEVWeVZhim0rffpqGdWsWvM+1mGk3eec3O/V
SBwHJi83dTo2p4NdmfuxcihJQqWluozqZcyA054/R007nx71kTMqtxmt90p+
TubYYs4/4wKiAGnuk/p0fVCIJYWQrqH/4kSu7Qviuwdh7lr14Y61bwGXXc31
pjLN81spyJjduNTtWhwcWwPQrhYuodO3/4oz12y/Grfb5UxZvvkniXyG7gbT
dn5U0UVtP3OkBMK6TzhA/F3nl2NwX7CSNBXUDeY6tSUWyGBosiNJK9NUpKnH
Vqk2h94dZJx3/vgl5SntXHAlUTe3joVRQ8GYGFaxRlvdc0wsL/P7+yQg01LI
/wbYHzDTNs/WdwFV/tq0DmWR7pxb75dsas7ZxAh2SjsJfJUPt53S9Q3DzcS/
c0gUDWlV2Q6ocybKnO6fZa0cB1P8Pk723ccxBeyPLW5jYgmgSXTC7Wh2KiXi
nCVc0r+BPlStrKfaZNt6WvelZWUyqfVFgAAjXKVFopm5corpfxT29X1yVLuq
dFXfQjKGI/vXQGys/f7hYpHc9NNZUUYFBMmKvPShoCq0MKpYrkIjKkUYZX3I
xyGJE2plLoB0yc/WZKvFhgtRkCQvMRJ4K+ScsEtyL/JrtpWanpw0upziRu52
ql1ycNz5NiNhW7aJWCYi1w9RFu4T2CsTsdWyygieAW/YmSX2M7v52fzltX8Q
pudeykFCEqVXS8wFqiLTo9krJqsJgCjv6XwNXiSpgA2G6aDSb1RHjQIzu+gp
fHy78yJ1Fkc1rKu22tFHdrcdqh9cy9VVMvvjgJcxYSc9Zpvgo6MpbxIFlguJ
TYB5GCPuRr/JpBGlhnmv7JMF9avG1/hC6SNVC4nkOarve0XPU6tUu0sNZ0ym
RLcL0BJPtdqAGh1MhvPkFN83kK2zsEUZ9dlDlV2NZF4nTZqXznqQMl+vMLBp
Y1bRAUeVAABh7amj182Wm7IeHWbThaY5l8ZR7x/AEZLwMyEzT/Jo9+w7StTs
jbqQmmgN6S12tUaaxaAUIqv/MxGUG/lzRU9nNZganwwYxOMatcXIxWy/gn6T
249z4eSFHmLzuTwb+k+inuTS8Kc09sBh2mcptJ3A+EV+QgDqMTrVdYUgzmF5
iUD11zhtL4V5t6TycucPvBpOx+Emhbu9N77bc/3g7GdhpeXSAFg678YebrQj
jziGvWa+N3bJygUmqJ3U33ofW64bYKHSTyvHjb6oA4hIthAiKmLaz3iH/JLF
Q7zMmuGpZ0bZ6veHTfEPT+PQpQvxq+rJiRqQh3NiQjzoKO3N2rlr2xeeIf/7
l/PlFn2ZtWVxRa3NuObxHMCBIbeNbe4cNttF9/PisrTzSZ+K9Pgdngs2ReTe
r6a/RgwLxDSPt1w31ijJj2Ji4egXBG0Q5rXpvmABYtm3tx3Oy+txIm6oRoUI
4VjyM4f2z/sttynFdccdnH1lflLXsuiB0jKMHD+/PNfD3sAe7FsbMUhkHYL2
jcBud/HkyYuRiX5VMDGIVWJI2AlhhieoQM3d8GjBMu9Oi4T3KHqvPM8dA+rC
VJ2ZLIgLpQJO0NOPAUmNI8B1oouJtBLnFnOzorH6bI6WAOMbW7MFAHPEUgLm
88mnmxIK0aCTETzgRmCgbrDE9jJxUE4czEpYC4PWnde/tcL01+qtu77408m+
ZlWmPx3zbn+1LfzM85gSwppgcjwuwWG+4gaeFXtf3tN61/8DW/CIhxKoW5Dj
djWTt4ZlDBv0k4E9ttcJVs+SDSob+JuBJxq01yC7O92PtDveVDrynAZE7Un2
1fQErObN8rpZUUiOrRQg6tvnm5DtyAEOeA7pXKCSoHZeslyZfe4zkMitEnUM
ZTYhqZFpaqmsSA2LoML4RUYujlXT6Whh5wr5V5pvvBqcyAJHkW5/MPFO0WeN
xRLF3ktyvd6ZfUObE2esd/9rGNRVL150jbWpj4z1OR9TzIeFfcM8E6uScqd3
ay1ZJo3UgJu3XrW38Rh/ZUqw9+zF4UhGxpnBqJXRjh6MIL5GR2u+oMj9QHxN
ttmXlKZ6BsvNblJjCzqmcfUM6WxOoyHIhmFECogvJ2ZGCKpLEmCpH2Ypns/0
qIM0gMCq6Vkz+USQ4XcRzcPIoG3b0FqGmc19qo5VNGfYuFn9TjNBz48GmOh4
XmzVkrwhCsBPoYE5dEkyRvpHYyi8kRloqabi0T/yrcAcc6O+1sUp/CV+CO88
KrVQbUZDclX2B3ykf3VdHhwlJQIu4YlS9hXbHNqVlz2jfHSw5YxLzunrWjix
/yk8Ou7TuGhoQtvn4ApTWoHLPDDVE9Lu7bTadJE4uSUpe+kGrL+uiBJQ7+fM
t5USkjxSH0aDHS1qRj3PLk6+ntgIlTwlR88RF/aBubb7IOx0WSckmmPPPtOD
uPXcKTCyuOo4RNVHwVNdlMoOCgGBoTb9Jr66JdjIMZTC+rNZvRhjHlMKyZMP
O04x/53/bp3npIMav7p6QKw/ozsrcu0TI5IapMprBt7uU7cE7ROZLv0CNxL9
vRnMZMwKzFyuNbZnSGbOT0zl0JM7hmRAMzG0YjNVl35QsIacF2QawiUvkPDa
p35BsZhMzU275xcz7nv8lW6RWRjXL4r0+k+D0a6ZwLIj0riPt8lTvH83XK6+
iviTzU9+7AvQbqySuUBL/G1lXoUo4r8pf5m9UmoLuaHB9mhllUStG/qfKJBq
s2m7EVhD7JulrKj39/FId6AvTTLtX0jtERj7iL3ni2W3W+Oxo2I+4ay2+hJb
tbfEIla97FVFGdBvm+c6pD5UE79iGmNbmEcdq0G/FFzZc0mqUAr1W2vguxc+
pM7nOfaJndHA2mAkDGXmars2SVEwkoKDiOu36Du7xYNfBG30Qeq6Hgma2die
yZlxy9purqV3rnQ1zuTsRBgyJ0KgY02eIyUsEOO61pIhTsviy6qwOLEoQlQ+
jHz5haNI8GwKOjk1YSoB24gnN47n8SPyl/5Lg08IiqOCF39pQUAeF3xGRFkg
z6X6lsJTkbsm+C6BXPaddFFTYSDsCUra2GsBAELGy5tnoil3hj0IboVOtEwE
NJZWe8e2qjRIkOZI/OaaLJ13gga96YxvAA+RaD1K1dgNoQKUxqzuVk18QBeo
taJfvsqUGnhsSm4L2Pex0uL2/jjsXJHn7JbmD56aSyPMr2lPVOEghjxNTDZq
Xj0BTS0ylBluZLGT5tPBBx6A9nb8xiGIprKvchJgcrlMFDTAMKtEXN8tjOd3
FM1UazE9MA7y3jdl2m7KRP45dlsl1hcTuxVC/XvEOuZJhRo+W23w87UZpa4E
Er3p+0GPO4JEArvKtXKuyutGU/PLc1si+HvRe7ThLR56FEOOSfPnhDoXtj18
uc5karSTHVlllxaFX2Unf0EgO2R04Rc+yjM/VMjHb7p2iWKMWcHLzqaFG9Ch
37jcUhsjl5eyqf2wZ9VOkx9xq4dlVppm8tQuprjv4smbTwWveRjUSMrVOeEM
skpbCZhwCTBWuI8qj0feWz8/WLBG+RByxIqZESrLRniXLYB/495o23Y9Q/Po
lK9Cv7kYAJxU9F4XT09rgd3upWjJq7ar1/KzItZDxJuHyEOQ17WTY1xQ0Pw9
jQwf5T9Ly2sCmGDE5FHEHufVJKruW2W5Rj3kQk1WRFBm1hJFrKg3YV731KXQ
IIUwKKS0IcTfrqtEWIsdzMBUmYPRL4tafOg0UkIMq132G4UZNKW0IwgLh+xO
pBADCreXub9abaUyx7zyI4gGqLdRG8OKU8VDC1vbw/u3GoiPNep/H4Kqdoo7
tpGYeif4/TWSkbeo+/SJPqlqq6YfdYRTQGkbPuCk7t1GBybT53bSCgR6mD0l
1TqwC2OsgI0v2fF/o/n+oE8PV7kAkILQ81/dix1oUe36mH1iP7oyO/HDdW/9
3EesFZnlyTIAXtipEQydwKU228JDV9RKdxal8hQp5GZE5nWqLRbjixmaPqZF
pcj45rddNdvCYrvGX9KPmPjnJIBE2geQPRPS5555mxLeBEyrSG0lJdmKbExX
kIC/XWHMXoYT/Wqov4l0SR6EA/97HmoW4xPggJite+L7lnSvRc5fWJm1iHDe
yoOYyjgVDpKBjKrSo40bm+4AZ7VxWqrIRKeKsip7DT4UPoy7S4aNmgN+N7KL
0g09lfeeJ5fSTGjXSiLQOTXod5zCLMUTXvqrNyoTp3CAIatLNAXLOmaPa1vd
IopyKlF/bY9EtXglXKCCPmyV2jVuUN+TDfqE97b0Rlvl8ZMHD5LdVche8V2z
TwMs6ZFvHC5WtsovBJURtrCj86K0tGyBvXiqzu1twkxR3Tmc/alNdAwNg31g
f2MyZ+0iBasSkhohcrEbURtB6bv8J9SQxIHwVUTzpwc4YA50GFE0Q44Jm+EQ
SuYohJU0ndoxcW7nnMkGupKsi5XAgtSYVMAC7ugIjJMMhtQSwYsAIL6XS/IO
7xC/7Afw4jE8K4/QWujO3V4iydfag7/hR7XKVYIBj5ITvsvehRhH18cl52WH
ug==

`pragma protect end_protected
