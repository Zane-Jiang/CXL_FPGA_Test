// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
FUjWTnCt7A4Ntlarb1Xk98dUg16aC1jKNyRMhxBLlqe09803282dcL/CEm8bUCixbGUP/8BUydRj
JjLqV+OwL8IWCW/DVFAoOpXolem1TZWN2BvNdCvLTVRyZcSfjFsNvOTFa+yf2upTzEeIFBihak+q
OzO7/aC82b+V6RZ4BPGurGhEgMESRmxff1d9dINlwiPwTNeza7uXG6mHbIpMr2gCFqKkLeVN6AWE
/HJPw6vZWD5oWuPz1iArr+YNBjH5tkeimKLyadKZgHIuRRPNZE0vRPxeeLcWUPSRudArlXoNnok1
4p2WoPggRDF0+BQFpi/4LxbGLDLenW66J8Bi8w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4608)
wVnU+V82QpLcrY5FVKCsz0n6514r5k8XzH1h2UtMLlK0IKNl/WeD0Dt4NgDjKgIyqkUXgEogPRGq
pV7M5gSgjOaT7iwX/LWgA5IKUnEYdNB5QQ5gTaj5TdJl04JKvOuhLmhcR4Z0f6ExhKmvcmVo0b3h
NTT82RxajwQWPP3cmH1osvkFJSbQm7RilpIheLEEa6rKFhFBqG5XnZg113UdfHcEiiL3aErTtKei
4l/ZaTzBQcJEn1AuuMCz5HiVsnlzgJ0MrTgL8b2X0VGeRBV0Sb/D/U91neXL6OA4lnR+um6v4zJW
io6hhvFqGfmnwtyIzS3rbAniL3d4+ghbEomzhWMgxDL6ZfMvybXZYI7Fw7TPX7Hn5gWMh+TQxhBU
9/9aEyozpNIRoaec8kEX7uKwK0zq2V3bmJEZhLSjs6B9lJBZ5fx3AM2K95uIw08zTPbqd85QZ1Qi
WmzU/I/EDGupLy69N3lLxHqGeysXdKhoO4YxMLm1OYEqFXmJHlpLO3UqRDGqA3R09Qo8pZ65/23f
mHh8lIj2bj76nHpvey/h2eCXMDHldqzYtuPe9q+FH1np5DzNJrgwoxei+QivZGDn31RqJfN1QjsZ
c0NNkZCefdY93YWqYrk31AIOQDNVoDGX+RklImJbuw5IY7WshzQvHQPdpPf2QegoNFM+2Yx4xySH
Bz65b7hV/ZTXc94p0c7XXI+NO6PGHBcfmGhWl4Z/fXoNDxw/NtGroXznzsXWZElR3/uZQbUvUdnQ
j+z5X37n1Inc5217kEOAhnxTRW9pPlhzSKqfS8+bzi/49jGke9v7vThUgVLNjZLa/klBVodsxEZl
MyUTX9oPE/OvenbbHoFW9hlG6FjBGcL09mey9cS7/lKGVZk0/PY4lHlJA25p/39EM3+nK4BqHgws
seK3/4dgnZsjZzNL8zQJmfXSlVhUqULvKL3NaToxiLcUWTlSc8gvsKcHJ6OyDcqVwFjjWBDfwb4N
4bd7v2vggih6/UZbQ4abNGt5KzkkaM9CWhbakK2TrK47Uf2Rs74N3qgDX2kIayRH/kYcpJhXS6JX
TUW7tzd2nr0gamRd2N7uZbCSGILKcPuLSatLf36xi0pTsX0Exj2ESpC2irpl0rI4qqzLyMEngzyH
cbNq1R/apZcyKnI7W/ky6UYahkTLy5ZYeXTcWwQN4fnKfLmxORZBpLdsf+K8vFfo6fftqh2yUvtY
j39JwLQS3KEwNRuKl1eQZ90WHVEp7iXB5iWP8l4VQ9f8GMdky+MQhDb1NKsCt/zKg0aE2XrvLLNn
bqxyYKmK1W+Tz8UNtNdJ+HNrsfO/R4JV+pBV9LTvSdfDAQgX9sujWzuw2rQOIpD6dFvLwo0U8r3Z
ISOshK0Z/lUwdcHZSWYywk5bbcW/7kEFu5+G/1nHxq2+wjGKbNGWigP6jQYX+i/ycaYcpppCBQLh
VYUlffU3VURmXCjci9M3e7OVH3tEITfl5DF1THBEh951DZHSVpwr40jX/MlP35mRHVaDrVs+RIC3
W158bWUeUmuEVVMy2Pk+nPN0Gc6NIfVWYM36AKAgcHeGHLbivqGUgogRacf5jgXcmgLJJyuchDla
6XnKT1LriygbmFJoysJmTZ3i2nXC4DGGmG5WPgV1K11VdnPw4BZhh/VwxY1dGuzZMxawMlNOb6nC
8vcpk6kid9LiUO/ryWlmCzy7apwHX8ytQAn8syO/qyaL9OIC4GpbvIDF64snG+5K0dA2COJ9eO62
udEVscOaXGSee/7Xusd84C41JyfP2iETnOYtoFAx3bucPKH4zbXZHbPr/Q4wZZc40d38OWYNoG5M
lSJihT7M0ZtWXmhZMSpgXgq8HTaanWHo5umGNYpZWxC/Vo3ncfnVj7Lx0LRGXvUUmRQqdpjpUFqn
LPeJQOo/PgRKEU1HrZ0HulHLhPLMYEvFO/REroko3iyw7JrftzKxLBSCn8MHvPzyA8etcJtqk0hA
U6maMcWScsBdB3jXCXpB4MJ9DxqzXlF7hyLZmR/WT+wGgfT3TF34ApLU24+7J9nHgylW24klCZN3
GDimmkIheCFER5oy65gnB0igXDensy7ZKWML47+8cTWAFR3jv7fIr2NNxNI6dAwY3y2OizPd606r
VfWKr/ykluKHOE3XSCccnGUsTdpS7Ots2wcnxy3N2k3VUza+Q4YH931bESb7HDxEceH3nWkk//qZ
dQr1zSKXUB23YT3zYjBwrj4dG7yEA4qX+u4iSekyxQ+uZCYbsLbG1Ty+VdzB34TSKomUSph6TJXh
vz0NghpxtRy1+uWVICnKrJn+rQGk/RAWJ6YcFB45e2D60N87t6fxQqAoz5tdbI2zCrAukZUsoK81
HRmCIb2vRXcVH9ZhaZIuTOUj+OgJeDd636a1LrlO5gZQ8b7xT3ygmvnswvXrJILDacXXGFtqq0KK
cRPInrp5/FTBxeXW5ePrlhUEE7hQ5vldcugFOnV/CU5RuWO5QNy1acuFBFFbQObHgLORNQfDSaRR
SlE+KJ97pvlKljgQHovJ2Cpo3Xtfllm2ZxR/FDkxg/+dDWCpx6LO3tbt50qBfpzgNIHA//e018co
125vBmukVP2nl+5B1dUujs1GnX0U2oHtyseNWVICZeK6/Fv9LixY0UXrd5Zpo4t20uAx9RekKQ3Z
17ITkv/9B32ZCCafDX+/oZIG80gIH+zsdSpnh60I3xQJNclWSVEh/3SJfr7wGTUjstj612EnADFq
gNGv1ooVLWK06YqizilVv7+4CxNrN+WyfFAmioxraplP4nzmp7XprS61Pi7ovgXCaqy7VII1KfWX
7WNkAezK3xQSs3lpajd83/ETt8sr4NPhd1kREBUMoF8pVn1rUFW0GRJwCRQOu0BFxX+IgwLFxnEe
DRDvF4yl+l1sc8/ku4LP4MRRD97H1RU01fAoHQiJdU+wizgBuURP/zy7kkgTiqlle1V76soDcszC
JwYBIU2N+KehhraaPzHvF7NHS3qwWORQuDMOFsSPqTS6n9f2NiXzwBUb10beXqnSAGkYPxOHD8Xp
OCJUrF+HYXOxdgXLZ19Ybo2nBEuFqeod0iihpj0XU9qwYD6x9Jp6xtkQyaKFYWyeY3Ke+FqDxrBl
8XCZxRFvZFlaD2ekYKwGqEQ3J10kDZGFO0TGC43bnAlKKNWrH8mx+A3yAiIHK6Vm7dzijaK+3Cui
moA6SpB6ox2TY8AqCtMgmHeVGLjFmHt5DXU2YnKVQWNDuJlIpEUV6psF8+oGeAzWhkOFBqGH4pyx
LQJz+qzCyRA4cJK6Augq/Bz2z8RXUhOX6XC4/6+JrLwWe+0uggAh8pAfZ7nnCudcIgfOA6gHYwL9
ieCsCPZAFc63kdcv2ZRR5ybDQI7UjjFMxiaGjVhyvKcaIGlqgdDI93uTZxWUk6oyu2gVcEexBehJ
HXesyC8XtvLMf1hRRKVlzMRIsPpbDudbbaxPUuMbvFRKvpXn/Td5pY/ejHJiYwIXeGLXDD6lVqss
71cC2nY32L36+lbnoeutv77nV60ixD78rTGFistR+A2oRGqhrqOsQoKbxdk43gyNMkfroxo/s3Cs
eHDVKVb+yMFxdmxfSzQnidz9QKaFdyr8dLtNLZSFeAFGZX2CeNE7Aj+4R+moXFWV1V7X4AW5tc9b
05Z8Xxydls4a+HtcZoDbtBz7GXZ1u9d7M+frT8Wb0nUnMFEycEzg6rMO7F06M+k33Uw+0tdbODAv
p4eCB8ubwyvxa8se11z4L3cHezGrQ3ta6tEGNVT10PKiRG/5CEYUPgoUWfDV6wGI2nQCMqh1NvO5
6v4XljnJJBKU0J1pm+hcAFAMhEKkrOdvT0VMt+BByj75hyWotCAGx8cj399Q5kcgYhxZbxmehwmP
WOW9RGH44qyZLWzQgndWt24c1bKubdL7s2qp7P7Y9xYOhN6IXdSRMInATHjzKT40UQu2FwwZfewl
t0CrOFpkh4trQ9hBj6oVgFZCbiOWIBG0QfaWyfnBMyTjlgEDInQD7YaUBzT/BzzzkUXec6rsGBEg
ws+W6aOMxaR23nsROT9cL/Bj+uTdgjOWbeSrU83xOaMpvQbtrY3Ytd689hWKxU7MLzX6lWl14r9U
/odsnZcvEPfFDkcsQbPTDGg0pKid/R1Wk+m0tO6XuJPSiG+Wj1xFVGm3fP5pZdfon50FHOJ3X79O
C0TzCfxdHab37s5SRXOhFYZIbIGD/wGssQs3aUlr8lpVzrNSNJCytgRALaiu9fmjX6/ZSdgCHs8h
UhrakSnReNDmC6jLHmjwTVrWDm6f0/Q9/IsUfxg+q+rIzo+dXIxEg/gJdw2AZlnDaV0Kt+4B0GiQ
8EVGu+XnjCfq86Ob+1gRpsBwK4oyYLsLC3Y/KN7VoXfwbx1rctNXpmW0T0lpowPr/06fqJLG8bW0
70Yn5tDNpIs+qaPvRLa8uV3Cg4JmWZDh4SS9KRz4rJRNLH1Z7NwTTasWchbIXVVGJSIYsVHH+AZI
vH8y6dFB7yHXPalr09s/CKQxM6B8UsDJDpfRkqv0heMvo6hVwPYwLw+qsDjyX+03yowgSJxggzC2
pTQLqMoiLuVx8dJhQRgDkHnTcG4skn+9yBhhrlCnqH76P59cNb9C8yrffOJLT8+xuP7eLmHwzVjN
KI/ZZYNoJ5f/cIcmbSO1zjVDpu/WeRJBbyIrh9JCC4I0Ku011Jw1f5eeI1O2R3y3EXC4liMMtYoP
mg8IFBBNuKmBB2YUFbCvVqilv82XPXGTni0baID0ghjSuLZrRWBbhxlxHlqg3CcNYhZYstAjScYh
uY/mVv+35nU5cqqd4a1orJqnHJQrHNsFueg3vgHELUeZUYtMamhgSQPCZdVOcJ8TNQSUZPFpZNYX
4oh+zMtVzNz2cSIJGbkBtjjIRnOxWlkKycsH4gYv1ser01bkrJtN8+nClCHoUKhnLBzJzvLZBsFE
zypi4UjUxmzjfFvZUqnSv3qeuMPCLlQGQlbrAERPhMNZLNQ/mb2LYJbaYykyO9nIE2u0DT29Cqsk
ny3+dTT4qxgrarpyj23MmOfozskeq0cOsjmFcTO+7quauajv91myGHj6Pzh1Il52YgV+riNAI8xa
IuayVmXTKUGyWkYzdagPF5j1YHfFGVUys/auUkayczEog8BMcEUlDb2AWAMSIMkZPWH46ccm9Wr9
WrrIhSPfIf4zZD2IlycdpFYbgcWJbF7aZacD6TwWEVYYMKXUiHqd/2EDrCCwhXqBVoUOmfzYRwRh
7NogEjWYRdGaAc0nZZ3RcvVcI25dQ2imQAHQGF2XeHKRFQSJ9EkjdovaFAi1khtiCZ25hGJ6V6rC
qRFTLHNzlTtYzR1gDIaRUWQN1TUXyR+qsPwQcMesf3Ov8hifwLgI/ohp8YdPXYRAaMLvgFQUBABa
EbJX+7V8GnIj1o1FvsvUSxnPEotMvV0v4K5ppN7YpS/PJTWIhhO+w59GRbi/P60/0CL7xnVUlGFd
alCgBUlLCDJCWACYPLFxB1ReydG4f0fqXe4oCZmT3T2M1EMh99VYmDMKFjVeKT5Tmkmk9AYbiC4Q
N8mNHXP0m8YxSaFmJIPKJm20L0h5bwxUIGqdQgsOlZMuro6p3tKz4cNzC/mnzB7KAN05RYi5958L
usAnMJ9wlS9AQi4rvrnGaB8H/LS32P/FosfSQD2uyzqpmEL93j93Q/DBTLN8pvvIjzS0HcVZa+3H
5Q5gW7XR3QVJ3xS8A5QZH9VjhBMq2xj2KnVkFnVr5vrb3hmQ5Ol/R89SrG3xSauakHiMqv8IDYaF
fRFWhvILrpw/pTipExWbzU0VFHN40LtGwogghVyGkRLUX+wuyPC371T6I4Bnfk3RRoGxTAAzO/Ic
+UYS6aW9dND8TnKIAftqZfmoEXNEg+en42+CZcCNSB60IN/+RdcglQAIkAkXFbCLW78jSNYU0LkU
B1gE5p1PFWxYALYb3oAtwqAXl4aMam57KtFtbJkgqxRpf4co7xAK04uTAPOm+ztoAFysvV1XqutA
NOFmfQNtOuX3KHiQI1avD1A1diK3gndbgRIwfLxtPJtY5g8vvYgL5oQmqUf4/P0cCQh8qVPppj7K
gdcmvQ9gm7VvlzcvwifHoz/OrGF/0Ozz9x3nyXwclZR6bv+pdou73l4SZi/IhVpd
`pragma protect end_protected
