// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
CWROTi7RDU+4KAanRvt6WPsY0N5SYd5/D8hF5dd3oC/HXQUmpgLYMVHy0FfXSrBqr/ANe9CB82bS
QT5Bu2S8FpOVEgpIkhGzTI4OCmYDqdhR3hyq73afIdOgclPFgCdN81VaN4Imrc+wgF6Py+jCED5o
MVdcbe+KIq+re9pyvfC73rxlOMAyUyMn7XXVshcjdRNKKuqWijlADLv8fdbjyEvYY9gRIjbU4JtL
9sUbH+b7HzMmyqIFort3Ulh/fdlasO1b1968kx2sMFcyCTTtcdv8kR0Q3iDOTl4Z7pQ7llAp6PNS
5LFfJM6K/0VIqL3iGj9Pei8F5NCCN9nwLoFByA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 91088)
5KW+Y1+H3KQ7TCPlqoFeFic4ExaQkIWIZlsbQYA1qB6kmwByyhxQlSalAhUVdjd/tonNVBc1MNZr
grHM72yd9fJUgtYF+N59D/33XtGKqC1IUS6HpxAney4qMh60VTkHoiBkrLdN7LPm3HnpQwVfNuWh
lxQkEulY0SeWbMAqNC5vDobQpG8qCIf++Ef7pPsuswxYZFpNkoUUEMUGAvz5yzko4UtTutL+5Ir6
D28btMhhfMMCpP3izu4DqlcS5iwNtxSvxeD7y6dBnt1V2kWm+JgYSod4kS8rQPIWQwlYTBjx3SYn
DQh2y1HBFHN5Fh7YzCJcQMT8CaCOIlqcsFM98pG3cXTmPsECcOrPPfl6qEdva1mhttKMP+i+BgAV
nO6REtwR6ODbUDuzvmSooDeZL0J5U50aB3IK58VfdGtrVnbCe5HVWnK68MY4Z3Fd4XT2J2XoIX22
2q2O7iSVEXpBy+hQCtZC6n5ZBE9KX1LFygw86GMLl85d414OdJiFvIvm7RWSrBGWUqPG4aJMRCwJ
oMuGVOQc8hK4Gmtsj0M9Eky5LmTNSK435xaEWUoFaG7VzFf/FqsjeObF94dwgYvX3QeBTHyT4Rda
fE2YvesBmyWTg1cbnawGTgd9gyEMi+1mmxmwRb/SYNAQkRSrdPyHEj7kf22yTR2XIEOjOhuGpkf6
PUPRT0ly2XMoexM/nwVaCU0sxMLMwIacuPfLre7XpWadifcbA0YP9y7enY29rLRS7C8aHfNTuz7c
ktOFeJNnrSzK1Hy+ZGgjaFR6fwPHFOLzjm+x93dK3wlO4mm8rvIwzIneCCVM4zt057MgytGYJxEg
PstqMTZu8x8DvyXfsgHK2Ul3v84mHzgPDfHJS9szSe8/R2yXE3zX+qHuKxBBo5zUPYVoAAPkPIr0
JYJtbI3GMgFCh/VRhyqqt+gvNquiHlqSVggIXxha44PtBR0pGZc/24Yp3zG0Xn+sldSmhjlNw5ed
CxFQwcdnQUgswqfKi0A7VhK9D9u2CXUGy59U14B33vOTrKF3y0W5hx/CrQQOTzvyYALrf7yj3H3Q
4N+NQVHgACRFQqM/LpuHLRpX8+4BiiQp3QHH+IVb0RFO4rkilR03HjM2H+4xNTUcVf9GmSrYsKXT
RHwneJ3PVkuPegSIT23o4fipIVo5k5DhZndDUc7ukLwXlLk6GbdCpHcJRkzNqdTfpLmZGiLTtTzn
XZot4treyv0npUTZhrsA2dPNMBGBSTi0CNmntbYmE/8d4m+zJSb7R3AdlnPh6F/dka+OWkS4zVRG
tavtrSuQYQkQM/67CQ3fkMUn2nCY04zmQn46Oek/W0UfRHBK0BL57N/AI8HtB9nho9vb6nuHfqi2
6l/UIBnxKd5NtDBpDLuiOs9AaqESzmRXP5qPKT0gWxp70UX6p5UkV4LpYLB4qfroneGTEHvIdgWE
MpheVAUNv2HUcfuJMGj8RJX1fOPvvAuZoyUD0ve184rLYTrfOOEpUglGhrzJzs0Jz+OSaq23iZvO
LZwnkDLzAKsqg2lnKkq/BF+0bcCkzD+INrSpe2wlcT3k6wJb4keG8VjQIzmbIhgk1heI3cpaLRhW
fFYVTLmgTZb8qor/iVWv6TMjZNTZuavVV9HbRJ9srqYkNSzKgtKe8A9HloH6nyzeh4zaCgNggef/
SlOG4EbAtwwg4WvDuBONNzijuT+CAP+cxeYBUd7fgBwxD2DER1Jt1nSZQ86aiF1WwMP5r+q14aZm
x4WosQ9XOEV8zuYb2MPZGCi5q6qTjdPabkuGkajFz6+lOHiDECVP8hXdLrU0EQ7UkVyTGa6p7REq
IiEgJ5UwPh9heS2Wf/sAR5X9IW9SJt65sSa4MW/+BRk+EbpSl9yKzLplAcg14b9ydHQ2LjxAvvJx
fJkeFmVSZtzvqUGiltpi/OLAbY4PgEZuwRtFqj7gCtaZ+xygd+iBnURBplujYF6X5ZCmgfneT9l/
QrD30Ap/E+eo/YraRkFFyGVlaMaKEnasF5KV265SQjh70BjZu0gAdX2sFmey+UdzUtAV+3KSzta4
yGj98vIhCOzOrbRMEcAyHQbdewH9CJC8LbiZBAPnhMHL8542UQjEEzxuMIxKaEfExIgwT5Whi1wF
xf6gaWC7wdBWlixVdPhKKdf+Ro/DNYMSALfcNtOOisB2Dd3ruQ0n0/BMTu/x79P1XBoQOwY2daK4
mt+css9MOfCGLH2TwfcW2Ka3GTRCcbXI+jE4y8M+Y8x7lT82djH701ur+QKdC3HLvOPSbSFBnHHp
08ZHem1oXjCCQFZtBOa70jBDG0cU5YGeG26jSskPFNMNSqIADbkdkNBohBtiU0GIL7vDK7sYDBJ6
j8M3v9vrhwtp/sK6WYnYlQerde/cHX4xWETqAIEbQgQlaet77YKPZUVu5EqNNrj46/N/Qsr6gt3j
qjyTEW3mVWkn0PFbN46nz8JZhFlWUgbcCpxxuG7+XLIb8NGZpUiv+18vTBcYu/OLXssdWoVdZ0z2
d5VGA+rdX5H1Idh7CoDKBiBaPkRh4N+S38BWPOl5yy8vkcUMDMTNvl+RGae0p3nqf+rbQaQl7HCP
A0fqZl77k8HxWTubZZwf5Awu+zryTb0q6sVzLGOIXEY//01qmphey+VyI8sB02njibFA+bIdgLos
QUVvBB5DXv+0fAXtwrOb910gCY/PAu6hgi4dv+y5t03dLRU+PAJfnfhjd1SlqSecgTq/8fHvh6fE
LJhnwlsKDaVwKp5bQG6uwnSG1KFOzRtsiHtUJ6LCVeDdcER81UGS82RdkUu8zbaPyuHaB3oWIh6t
+wvn3ZC854BAAFb9obJ3aLQzYqf3Bd/Fv5Fuyyln1ioQRSCTR4tzEeNWB+9NzA4giKgMio3QPH2L
IquFTzDO2u8fLQ4jm4a4ZDhk60aQf0zxhWifo+dm/W1Wfq7q/mguWlnDbKUmZ6zilj2Nt5P4klE+
nemUTG6p3ZzYOGmeXvyWRY/Qk74eYJcW8u6zKR5mUpu6uuo5mjOg6zABPXUHZjaAtxzqo6cYVtIu
7L8EmW2+BB4fMkdngeOhV1FQXr2Io78zbGbqJpvNJpdCFvrRW19n5X4NyQ3FmexHRIx83rwJcaXK
UVnaiWFcSa3/Q673c2RostRdMV0wzhihwYFm7WR2dTmuYW6BFDVBTHOXul5nNOxrQIemG+Ga/iHb
iecPGHvhQpccJBI9+ixyFsZmdgixH1xxa4d4nl6zIBsVbHXL/1VocnNPxkBYP2KfmNmzNTav3C60
W0vpqlxkJ5efTfLHekmbitvGQYqB7RT7KqMYVYNzywM+ZWrXcHIa750gFj+m1fwH2mBZpQDdoOT7
jFkizn1HoM2oR+rt3lFFIaSlTCYH1n7fkWdYdHYh1gArWHuIDwbfDd1d6/wxjwAhsRQQYUAbPgXZ
rRhkYCrb0MFdazt/7N853bxSVkp7ZVajFC6WQmuL0E4ezXeucjVTTO88G1Td41Cs2mZhgyiwknsY
1BYtikoCBsUpi6WzrwSCBZT22WX1xJ5vu7uT1f2MTq7eEs8QVo+cp0PsMg4KGJ+1YOHMfFlg8viQ
8s9RiNcOQUIw88DiOK0CxSZswULAc2t0Aj2K3lzJyPhJ1vgSpf7SPIAC2ZFuqZemG8NO8W9g2y9a
jEFFaUiFzZghJvXdYzOihv2QmFPOXZJTuzxUgWsKU22rrR0dm10liJifGAqkLTSz1x7bDaaZEmrW
hwye1bb7yNudk8XFAbUq+qu1LRx3yReJblu+9EcV9Rl8yBCanD0RcpuLKr+E+SVgLsfI4D4Zd2Wj
EQsXfYgl/CYSSnQU+1I98YdIt3DMnnFTU98b+1pkzPinOQZ1u9HGm106EYCGK5Qs578CRZZHJCgc
bDHmympwplSXizrMsfZYdrhjDRsEm7pNrHGPZk3qMIlQf5UMHKbl1EX6Wxr+/Oz0M7QTjlx1806q
GiA3VTA6ewkmQv5cljkI5RPS+xlLknyAb0spmGVbiH0iAZNpS+rDiGZ+SSqSBSRkN5bacBkYO6un
l59/NitYRGt4LSL9+E7TKlNk3HGuCLS1sLvVs8Ui9sj9tiegU7M3zzs4WK20gy6sTaZVGs11U9vq
doGkDUmV3umq2tgGSNpcObI557o/vzSlPqOX09DEgvD3CqffQjIeWm0znhh7qt/3+r8Zj3JOBNiW
cUiFjObXn6PSk8VtuvqnR/N/DppdAfzJ9pCMXAdBRr/4RtpdIGrxoJDQNIT3K3FvK9s79Ng8zGrT
8Q4HYiEhKPt6tQc/JbHw8dPOECak0ASJObyDC9+6yovUR9bAiGIB8AfqNptoQdBJxzze8kwAIFxi
zIOg9Gzu+KM5SFaf9R7rkasXeGsCq8RDIfGBEQwxdjnJPG//tB7LNkp2UcD0iuIVcsq2JPDKC6Yl
xLhCJDSzhTViW8x6sL2XooGtMFCviAKKqKk+6nqOEjqNS9I2GobUo//YCn+CxPYUmm4585TNMezO
Ui0GzHg6gSdLamPCZcINJtsdmWWYS4PwrKTQq2qG4r7S3auH9RTFijRyRZsUtH6LuL/YZhukvqiG
el/D/aEf3MntUhTAbWNf5B9NbZqFtvNXOsZvVmo/a8a0HvhE+rlkybY/UfSwOBAcfcC8sBoHQZKx
6bASaRRjo/afzYnEn62zfdKbV7oSFngEZEES2Om2k8hXIMnmR9G4K1pFWeBGjAQ8vPVc56T5X8QR
Bnm46r1QLngkZTHz7eQJOzFr9eGcIRc2/MUvmUUehcnYXqeIJLt7cyOgkWGp2WH/vRKo2uaBEbNa
GY7a6HlvzemCcgeXBuQmNmuDoddGcRTRTBCwmeFc4aDcZcMsbeIHm122R5i0orPD2VYCvxrPtXVu
xNZGpy7buZy9XhMWR0y8EGRVQqaO1F4MkWgLm7wm4B2u739M/lzbJRhk6fHagslmShxSP3X5opma
bTfd3AUQUSUibZZ+1Vxs/txVYGjumLCNdeXZDCpHjNcYDCEfeS9WGsW12ZMhEeqYUjKV00f2UjKO
ncrpMvdPOiGKOx1NiZtpAYqcuUE6OYvid3IhXxtabRLSgz259+lhSyfWeiAQBGEi5AvbD1MfTLfu
snQxC+wTal2Y484mCLouzPSo0HGOZvqpC6hQR0Uwmv3gSBtu/ySVjgFjd0ius5OK5OUed7g5d4Tb
13ftKjC1KKhxPchf8iJGHwy/VHp8VGD98Sr99eBly0uy5p8h5w3Dab5qXnYl3hgfE0j7v+mGbc15
7GdFu7bkN+QVSx95ANujOZFN1QFYH8Q006jRzSB2BCtO1mr7FiVlPioHdRdY3SP7Kgfqw+jPA9Do
Gp87YrwFXST7kyJZgCBw9Bq7tpCfTwGKFloG1f3UPHGz0SyMa154bQckXJAh/xoay/4s72IKJZRc
EsUasWpYljRFcxJPhBZiMi6CT069Uwd3xIIW8GYnBXte2V0Pdy2vlzpM/ARXYbC0euLpo1FwFKMm
pPTukOkR/T7ClqMHf1yNRHcRiw9yaFbaRaaJMCr14I5sREnGhYm9U2SSSTd8Wh/8+7nw8cv36fzB
eRlUAd0PbaM1FJGAle8SLEcrFZXRxMCSdsOlcMUG7GSn2IKAZneaC9hnTW5KNO/b9D5IBr0siH1n
nnfUIqYM1DklrzoqfFkyZWsZgU0VLbBE909FNtX82HqRrtF6YAZHfKAmdgTIY6I9lVjtBF+unpyK
WrpYiELnwSKwy3NzLAtl1vaMw54qzr0Si3LWXvrsDE/qEop8fUV92IwVHbb3OKPI4Zqr4sP7jCOf
81yONXV9kOlS/4PVxFJKsDWSuL8h3PjtMqcnL+U5FJ5iAly6s9kBz2bZ8NOvlmCf9MkLZ9d5xxy3
vK/t31temrmNvMv1AZa8BYkYjPDnR/DbLQ/I+Mx1l0q+/suGSBoONiSPSJTruUraB10y2moZ8e0L
5XaEYK10eMq/Ab/YG/0UYHCb/kdOfOgjMxkbJPSlGcTe9waToS9eAXk55T4wnO62F3UQ99km2+yT
5PDyFmtLJ0yNcVQ2dGz9mCusBEz/B78EcEdgt3JWccQ++cwZwq2GkbStXK8Xyp9Zg+DnMOr8A71G
/9fu7G1STdWah85Tw2k7HtfXxSNF4jvvM+SIs+qiJ7BGpIMdY43kMHeZw1PxlqiTpRD47UQ3QxuX
JNtWq3CYDVYz2Jeg47Vt3UN5SIlFDHquFckRWFJ2apJ3p5iYlIza344Izi2YMxQLRbSjGQ/3bb4Q
qNffh9Ra6EtuuTcXJM69a6yAptEaNN5HzTwxWUzLcu9UbrCF496LfuWczH20Q5PBrpFiulhT21cc
9x+ZH4xnoCNRChBzITUAOtK5QiDgG3a269X8BGxqNtdS4H2WkLCDLam+ezX0P6zOG771C2BLnoiZ
IWSpMTSAOMwUF5/cdGCkPMbvrI05cng9FW/w8ytduuYr59YiDJse8aJZovVNTB6G9TCgA2Lg9ovy
XdskNODggAT4Jv48nlNSnwtL0M/XvyMWlCZUPaQKEZ2U1rc49RgQBJGalBPGp0ubwMrYC65NHTu/
Ec2tL/OpD/+3yHc3QRG4PqQ4d/A9Q93gbfEFzLeJ6HWTZXoI5fr69BHOkjkFl9QPFzLtBr5UrzZN
/3Ehy3+B/9iBO/r99rItAz28/UVfrl5EfWpuC38z+SIcHJYjrx73w4W1o3esbpI1BRhkrlOYtGkB
9fizHaR0gehEthgHmPb2jHg5Qf+1AIFyXKQz7jYyS1uJ725qRw27ckzOXikjlp03zjFYvvEl3j4b
ZXKY4naLK9KfvBMJ4yA6lXVhM5vnUU5C0FApoZdJpI4PkqLaH8ZlPTo81itgDfxd/SLLAx2wlH70
0RgENRCipJq+ginbEYagLW78tns6JauS8YXOU0QYfKojpxc71IcnQ8+30b7tg9X01H8ZAD5pel+N
HjnfIMigs9WT5nEQEFLDQ+lBMGXxc6DWKuISCMYlQeORTMmNKr4dQ3da/Fqj2Gn5zIY7IvehPPZh
MUmRne5ljXpUCPnGU+cifPwdyp0JIRpg1gn4h/QLI7yie6NVvRWi3oVekITGpcW5G70Q3bgGQCzf
61xgdn1IAV0JQqnKlOjr3Cokc4JE6V/QmmjBzB7zuC4DB+AWOOuLho0yHAw/Te8ASywlyGXb+6Ne
Su+6am2Lnd6lsq9N8nMHofsty95VTpgFN/lRr10wFgNE4JDApGWruLoijxf3VW+Xlik25lsKwePT
phnPKvxAAG7IWDOvpjYe2iHI1By4MeuHajKAtrYYR0+XqyvNwuBF72Lr8OGOqol/TuVhY2SE44Nz
x2HjN86WZfNRpLWhjUst1Y9rXeCYOkydNEn0dL1kgg/5Yjuf2Os4Ye7CzRPuSY4FpVHxteMOj12o
0eQijbS7QBnIBFGi9M2HvnTM/P9W7zFD14eFuiq3W4EmxrXdAFrY/hkqG8bJAlGV0Nyut93O0WmD
coDDQSxFovk9eoRNOufailXb8k83CKgFuosdcyCACFepEpvrFRIDtBG6noZre5bjxA2l+Glc0tpX
2M4YRrzfHHN9lwvxnQlY/uBSA8zyvmw0gwCC2Pz+rP8YdaW4Z4t3GcoaSi1m1P+2cPCoEO5mrqz3
aIT/r/wFQ2ijTCPC4e7+wvLgDqF4nRfm6tEnWETZlaw6MPvUJywLpcoXolfHTkN6Nhq9QVxZUVDm
N8jdlUjrxXzrTtGTkSMlnyxDABCZKsknEVMLVtqlij3PAQoYQK6M1vWCF12hhBHfA21Qkg3NJCQD
R9F8uwBadpS92BGkMX1S//3RK/s3SjBe327E7p9obHU0yMAg+d+uKibxxhLeNABDo4wnzgEthRHN
WKe+qSLHhKrGsLAxDgj80V7k1uPTkvIM/gQWpkf9i9y5bni1FU95mdG7YY8d1m7gDtVW5o1TNfgj
PoODuTA/iCt2EB2+qQFkXslZPUqWL8cKEzjlf7ZKWSPxjucWbteBD72+Rf0dEXfV8h1HGBZ6swx8
+fe+I4kNsKCa0bxVUehVK+WjofXxbCYuFtAZs7b/adYJDJi6Rsb0LMkCdWaNMTxNnyfm5/URAf77
mRI/t+AVeIDGOYprbD0oPAE9QppdCt46xBzXjmavxVHY0QYX4k9WU9coomxP0f0zY+hRXcK67JeK
5mEeAuKNdqPJ6wXEUy0btl1ycmXvRzNz1ou9r7SkB0jFNOwLwXwAQDfxJ3wnkxXK6qGlBJht1n8A
F2t4ZYa6P0k3u5ADNn37zo9fPwD+rwZyEhT8SKyhw7ZMY4Xyn1o1ABKknp25cuZKWmEQKIEuU1p6
Tnhd4uzCCKLUdbUzR5wA5w+mcGNo3jh/GvegytU75K0ZKvv/b0DROMFJllIMtpbZnPJO1nMAk3gw
r7VQSpD+7m1dujG6xezsH/ak1l/Pf4zFImlijyxcK6+GMUUYmXVN2ZtuqxoX9SOivkkLW7fygYvZ
iVMQWgAnAeyeqv+XDPyh7VKn9DetuLQLlWkwKRJTkr3f5UfG5VK6tWuZGtXZaQLsN9oNqzcSR6VN
tmIVK5m6mLZwt/DHk0ZjlEad4lgF26hSjS8/FynSsljslVMiAoyxQhy4rRkWHCgE/yrLSVPYVVYm
rXwKR+Q6AnDtBLYP+3BSgv0Qj6zxLPT4iafTwmqSYFITZFeM54KI2mM64fWsf9Gc0gKpDhWNB0c+
XtvWuNzuBWao1Jehceo8gBZAmNcZF47Y/o0FHGSwM3yP50s9dtDqyY9A0FT8hzovTekvB+lknsrC
xhQf0dH5bBUhacmLcapqy1x38zTTUx0hEPyauft55K1wEXyb4wo8YyuHL3rxo63avqB/i5qi3lCr
IuEqJ/G+5JZdvvF2TB23L2Fi51T22X0ZmwttxEC6Wqh7xW2I6Fe4XaoKEgjtd2QPvnsvrG88doJI
qxwaZxkt0nxtF67c+PDnlVjrwQt1jZoroffLbxdGqvco5o39W8wvEfLgIXhDcQDSHP/rQg0uMX7t
wUAjU4Ny3b9mQH/zt7qD8dWppUyXyqgM2VxWJVbtFFp6vxrTxFSAQda5IE+kOrrsUIYKUUur+pbl
yUE+XmnhM7rktjxRXCpXvjdUPDospwR1tkZUlsrblQEQMnEkioV6BzB6WlVleLJPOVACq99Sh6me
+OvYlFAuLCAysoq05onUVo6ZVlbvwEfPlTPfDiJ4XJ/uuZ6bSE5vBrfIlA708P3w44in1JADodsn
fMzE2z9IiLfbmADodxJUvvdvZ8satcvizOQT7PmttVZ6TWqqalsYyHO9yYrXtcogVz83vZoUCpwy
CEmIiacl51vl52bQwq+oK3sy+El7Wk9Pkl0Wl+zSg8wz61RxwkLREN92HWa+aUTzlE8NRr+30x1Z
pa6JhMgI7h5g0lmcj0v5ITEH/Mt1ntoeEoJYNLNm1/uaWEyIm4wcHmZgpI5CG4Cqd9ho2hu6hxAm
1OZGbsHhqt54GoLOeylLoSQqoyXlRMR3oEdOMfURsFownx/+zXYp35ZZBfc8VDnqqUV5ZiC0I6aa
M94PElPbFF1g/ThsKeOfnGVlFb/yvnRIZlhjuAb1Y0AADAALjhERvW3Jlsj2YPDkpeUJyAeje7gm
KNMl0icgkfv9DphhuXO/LIfFe2sWro3GNWpDqR/SiF0s9oLmUxaxQ3dz9x6eMSZ/b7ulIWlPM/Po
k6pmP6JrHy4cFR58wuzCFmgujmksbnmmC97I/8Ox9DdwTryFMW8edHP3IvzI0aSS44I3KWXFqBn7
zcVvVuHdwKjp00k8W3cmwY3+gLlWKZzcNWa3jbOh3sg8GrQeQRbOS5NMsQU0A9rDIdlhXArLo9Mf
t8xJRz1rvj0iYyntsrJ2o8ahcMKkWnG2hma4pj28aQqfbIrw9njRLftXolJw1XP3y95zJfn1HROA
qUDx7Cmk91uqAOPwVIjKQpO53FXohXMyEeLWfRBFaGrcwnkrhBT72nH0XwN//mKAOpYNm8ogy8E2
nJ52704MkBgACFM4EytXZ9RqHQC3kMZFn0UQG829+tBIpl3kEjXHl0Dd16pHUBFCMjIWh1W6uyim
ywWTWhdkCwoTfbaI6AbfxyTmh2x9za3CTR5aB2n+OMhHRofmHVFfLCXsIer4tNoqxchHADiUFvIj
BBcLCqVY5ekxaR7E+TFmGcvdg6umpo+rdaxVIgA3KUjE30WKuvW/haNT00uSphUZZ4FpRa4R/vGy
3aZUbxRo4IqNqbDqHuoC7HOpZ7om2j77IH8K/cOb3NQsfEHAo/2JQ82GTUTKuAdpbyAOdr+pvg20
/mOsMxjqXWiqmyDu0Gri7XqD9VNmPzMcPt0d5iqDFSRaAOdxt6qDQ0kURpH3A3mwofmUgEiJxUSO
fBN7hGTp8OBCL//7JHALWdo8dpCKcs06uo2tAnkHCA7AIXuGN7J8ypi3yUQlSIeMsff8DtyeUL4q
+xZ2RzCLUBUG8Tr/kAsf7nX49DQKnoDrqyBNCtSJ1pxlqK/dPYcfMc4FfivBXhNP++W6PaGdrupk
ffYCkAu7rfFeBI80uEarzMMdKJBlA+chTzfpRA6vcqrwgzzhmNcgKjPHLauAjAylQU54O8mHixzn
Kno8f9WlYf1VbERU7JCWOBpvSwnDNbxI3i2si1a2zxm0bjF858jrX5CJY4dRsnpMEbkweU7YAvFh
TxWFj3dTR+PKX20cD5mKDAYOFB1gEC11jMzllzVhifDR5PnOACbED11+7UiH6P+G26z3XH+EpEwA
mLeoF/42QH368c9bJ6hyr1GToTuxPyNMRjQmCkojAsXzxUJDMwzQqyWrR47ryNHF+RICMTiL05T9
fFzs5YfId5X4T3rLI27EY2kfQC4jn27+7kZjXlVNhTeNW8RZJ614RILP34ls6H/jX0ApBnwjFOwg
McQtnN71m6bKTDSGlv3tH0r7UxKkgLdMJxRvN8z2RNQBZzY2JRkjp+y3fHZ8DMKdsgkyVzYfBAfH
gsZ0XTwSTwOrXIeTcwbF7AqIisXeKHCcGmNnkf+aKS113LhhX7xgIB5ji70NGTsbzUXmAQ23c2N0
7sLEF5xFC4XC1ZQoABKVf+/6RzbXV+LIlAKtEUSgbusLtAyLUIFiZZ+zoGNXm/B9JBHQzUFdgJvM
pPOTXpBr7Q7NYuUA64QoXva4ZQIPWkPChhK462z6oQdwjtHehOxZ1GKFnsCbMp7/2684mZ1i4x3L
HJvnJ+bGXdtKz387LEESoaOrOQofbXoZC8f4Oimr5PDvoRFs4sA0RxZB3Xu0nvRooUWS6JQGXpx6
PgxJKEJa85VClOG59Tx4iFd1L4ek3bS2aRjrLTXQW7CF28DEM8iAvZsC+nMe9Jt4AnblVitUS+Uh
t33B45kV6NeatPsZYjC5iVS0zBENMGSYJ8IzGW/hJtVLKR8R8efYL7gFvvwyPf+goWObf6x+4OEb
weL+RZ1oajXodHhBVgLt5AM+OQwssisSIwY7FFLhMbGtT0CJg1iG98A385rPtqp8dtZRArJbr83B
U/KxfVXKYBTsOjuNS+A9uOQBfX4E9xAFz9VAuO5yO01R8MtqP/JpxhGuO1RPGMqEy3/MoMLgny1S
1iWzk9MhUyEQu+WoUYMRKJ40TiuF6IVenF2KfGTL8AcU2fOQIRuzMQoHXkUgBhyA8C6W9qOMGvDI
8XEfqdwmUTlzKoH5CgYZNclVF0uGV0as+7a3XTDmKTVWae7zsqKLioTFXT5g9dQ/CIvdvxP14u7C
Dq5tHcsNgcsCzcWYBkrRSTV8HJ+GmT8CjSN2XMPcDSd01vqqcOJFmsr+bzPEEyq/HOg6u8w7FLvJ
VcsTrElY0ARY1g1a5CictgUk/Ca633ZpDp0d67Ea86gL3gaV3GIF06S6ffxUdSc6KBtVa+C1/kIS
kIcwFMqTUMYw+fuJjptX0m6iXtv7oDh4mdKtbhnnQtviwT02U2lgudxG9QmoN9ZxDhSgKMnh6du7
OPwUZKoWvzGxv5bIYD48pCUVTXyCHmfsEjJE9J2spSkv49RmYYEsyaVtfzxuUr7GxwfpAH2tR/lZ
zbs94QOeRA2+Ru9p4Nu1ijZK94Lm6SSaqzKBIbNetqS1u8rJ/W6MNicd9JnyiDsdr+Zy0cUiXq7j
wfmBhK2orKAXrDm17P32Ffbj2k7VcK0e6TJxVVQvERPF7aKLhfheskArzdtXPfjJmP8D+v+dDwy+
d4RN1omO/7VOBTrPRtkNNGjYXmxPnZCEaGJR2qp+jgmu9JwXtZWEkWvK70/reuYy0E1QDcRdjnA6
f+iJmEPLEuajQDnNes3ayBlWLj36N3yVFCOhiy+oNAmL+r9inESDNp99Cwu5+mhjmpGpVacJMOlZ
p78hLZRktcpXZgIpKKu2vhj6dBCnN60jSPZVjoItuXhYr0j8S0dj9yWRHY3ek0gkDCDSb8pF6pgY
Hu8BuH++d17JqQ4ymyHBOkrYnzn/oWDOiKumopfPr4DTgPfOnLTS/jq8lmJ0OdOcnFLaWjjPW9zW
vr5/OpB/e7qlBr22gEifmziGhS5cf9O9u+KdRfE01DeULgFkuKl7bTE9uj3Ls58u3e6VmgXYzJNk
J9IVtH0r+X8opdaD/JsYRQzmGnrgViRh2aBg96V/8/j1dxY+3LiJAFsKhbdkt9xCGmXWoLCmomie
NAGsCvjw13BZFB2KmaiRDHknP4Ae4fntXb6mFL4Yf5bgYE0xE0DvWFEU9sgngfYibhagRQOX0lTI
oGWNcpzGyfG9WoKdGLJmmIw0kpRy7MmcrGFdYN0F3XVsPc8iWUFNZqXRqBwP5m0dkDDycgAqe6fP
KGPM4L07GmhwfhkvlJTGzNe7obV9mkTOe09Dt0cRLWtIihPHkARjah9+YuZAFbXJrjrmqIo5jmIv
oBVnMhqVgE89pSPswolVyqypxXeLvCg/wUJM78cGSOnYtNppIxphvRR2qajHapgG5uwhds/IA6QD
PbeNUWQmDozQIdCEKlU7QHWSdv09CowKca81KhENCzyZg7Pe3tgQCA3SHeEXhxWxqtk04U4Nosf+
zRV9d6+K4YwiyrbRGYu7hZ0vliGT/k5fjYpDh/Z1dMd0cNe90ONjsSMqFRGK9nsLafPkS17KrK+A
SHIFEOvE8yy39w2MUhRe/u0vTpuk82ulO/27FGJbcpgnnT02M7Fe6RN1gVooaqL4lmw7wdwhd6My
ZGezqXLC1VLpc8flqvCb61ImeN47CaJX5RGdEBVPcC7W9zlG1GbbGpDDZbZfz6upeJ7GGdbMzIv9
1SSBSt1uVWs3ctGb9m63rfbrMh7jlpS7FgnqpaSMriHTlj4CvVTuXf4U2lgsWVKCw/J7tch933tS
cx+1ZN/TboTIq5S8zuOllw++q0obi4M6SrAdVanDKl2VRL+iXQ2+xpHXegAYXOg0nwor6sNbRECW
LeNCZHPYrCS49XZnmd8I23KzYFEvo9aV5y7zJrPzQ+RJfWm4YqGPPYYBizdtMSU7828XjRGUfghU
H3kODbJiLDsBZdjghKv8hro/sAbFHrsvxB7AbgdOICsvPctx5a8VpIMAOcs4ET5N3TFyPnhhqxE0
eUq9zvUiIU0YDWQTRDVvETl8H/9SwBcGPaP1RVidHQssBfyFhWYwbfT8H8oiLxu2HBFOodVAUyFe
hCk9QVIVKzEXWIdpoHIN1vQe8fKtzhuLexmcbJLvWYHid0Mw7SAMuUuf9dwVcxQ4Kmc8HNz2DPnt
uBIGSepVy6Ar7TouPhyLi9YQ2yUSIt2ePToq8p6RwdP1pdtNocoOjENsigS+b4Wq4sdDRVNscY/3
Bde794hFM87kTk1qvgf2JCapoQrbd1eBp+ScDspJhab7EdBd3+nZtbtSNJl5SPiX8MTPA5V3d/uN
Za0nMFnTj1XjaWH7qjmG4udMv8HfVwIm7ni4/sNaJTQIfqppkbQkTfmV1036e4p0WxwFY1tFH8L2
lmWLCVa35wKh+xSliM4CDTdixSiO8/NUQrdW8d3n6HWAJKE8wdmg1I4K9DW/05e37F3WFRs+Ul/3
/8suJpBqu2vbIm9Yj06Fi/hx5rvWOLBra431eqBZgHADaWeysV759yoz/vMtYD0QH0PwRuSUJQ+3
aq59He8hEQYNy5kdir9Oi0nW1aMufWdenCqPyPlwNq3faVz/p5pxyQHTm1Qtfe6kRCkFCa04+ZMR
DlO3sVUD3TLqoS09dvfl7ANwsgQQ9LMc+SoL2cnfct5HPbhT18FfZc7e0KEwR1YRT5/BDEpLxDE0
fiD7PIL8UNkloZi4p5gsrhj3pXXAHtYOKIvyJcDklkq1yOKuaqAuTZT8P3gBIOWWJ+m9+6XU/rnQ
8n7jfoV+WrG9ivYjN6rldLHF9ovcS9ZRBBYj/pAjV3GvDD1pS70J8LZUWRclQ312EnDi8pnTGIis
fT3ZX/LIWBLfrrOq9f2R1sDwLG+ll2NMFInyFzbe3xwCpze8NCEfupr8kE5zbV2a1yHtoe5On9hK
qJ3Oqi9RaKKJhAMwIWxzeZpKlHOa3Vh3Vi9WirI1SpiVmEsnyzmIbDZ3pVqCao4SzDEExwSYs99i
I8QjcCJIWvqqKDHJe3tgN/sVWHM08Yqt2eex7MVE7eSAO/apY2+NhhMeFD0d//PIUI3qfqTiJWgZ
dqv6Zpv2AmIA5PuwcBPsks1YZDPxvw0NlwIw2AnrbpErcuMVQc+3n5FkTMrbXWxVJeLOsI0hLJZZ
iJPcrQOWjtb6dbbnX4PjbX8Nie4f11Lbv66Snut4sABOjcHPCShSOrh3LUO+Tx+v7fEY8YPMDQwH
MZwYTwioYInCsgQNkRVMAcj1IGiK6suA/y4DyPgAgwJVWjn4AFcOu2gEG93Bx46BA5QBNeeDPK4L
qKEGirphzw7fdypjreN5R/n5O6jHVGWf9uw/IMmjclq9yY/cSUdqXfgC5WhSRDwaeo9EnIgyCgnp
BYZbKy35Sj6hn8VedwbCfymPcWRGvIqPHbQzbdIrmM8rqRP54cHyAfKgPSniCtdqXMI0QZi1bUqk
8blrJ8tHdikgdHNNlq6cjdisRJt6LSuAu4x64r+urtiVZapMvnaIQwdvZYRhucMgdljMrC1Q9Mo2
4pjRGXeiJb3XPNxyry6BP4LFVW6enF82wNOaoUhrAB4S3birQbkjawTXPYVX+MVvoXbX6SIrCBmG
0SB5DZHZJKRjoci40O6IB3AFRvNm+c40/ykN6sv4DRRVY1W2i5nyupzJbneEVi3swfNvYPj2qcpO
2NOoj7lH3FTx+7yM870Q/ybTWY46mwnkzE6KvYS5P+67cmt8/UcXhJvgqLEXZYAttmVGb87thbR1
DaccLbrP7KtI5wNzyd/AXcRcdTSPNOmSbDSm1wGpbBwwLmXBu5PMT1QdKqSzPUJ+OKmcWMhMtqcp
IV9l/DPDUrADFTuLErr4QFFZzPJn2QEcxHbZNVLIlkBWH2N5Yzcd/2qbqktmjax1J4UvEBUHFlvj
vSy49Yu6dmqW1/XXwS0teyqZI+iEyiM8GfCGuXCbZ8GMHd3qhjLhI87FNtE5V4US2vaSkByreYLR
pMLfJvfDGyWdFIn+ffzX2uQwCS7eUPYTyG2RLAZ3XaT0LQFCO96R7weM86mZp7SYyJYoLegeZyDs
3G7k0rmGow8C9x4t2/+MzSnH6VMk4kKy2mFbXlGSQeTOnc974Pr+cCDVxFc/5aAJ6dCuk/3Pa2tO
jZjYkf1yh7bGdeZdxbTaqekw7pAXV0HuBUJTupyYocnq5QQTgLFP3glrV3FAD6h+o0kq66lJhqXE
i80ZZCrxM94DVESrQaWf6U6KhqCTZ7hJkFdC7wCkDFTJ8JSpuP/eMHnYDWlVSg0e3Is88UPd5GkC
wE8hEKNC6tRtSfodg23ikfMR/9p/+fDyL553OeHDiWBFKt2TbtjGEQ9g5N6WNc0GvlUYOqKO8dxM
tNLgek/a/QNnj6SPVQ5ppw9ogCT/VBNAiB+SEVp6eoKU5s+5G2A/ge9KBNtatJro6k/JyUHQ00q2
Eh7yPGa+0RHEB4KmsKyCSqNbzqhkk3QVNNR+QdRz+R1w7C/OJiX6aUwM2PkIPABgHlO8KRR2SIfK
2lL+ZgA+DEwHXHSW4uzVP62Xf22MgZr5uv1dshAvauELQxtpc4dQTpmU5Xc51S2L35c0g4SwCiLT
aHtFnJvQ1t6WgoKwrZSDOYqQbm28ULhJjfCxUTMI+25GyHc10ITCBK5tbGxvq1U2ynXcrX8ypQQJ
SpAbSD1rd2f++t5jmtn0pem2Xp6pBo2cK5ywq3NwJC+jjGwQiV4SIU40J/jWzKxrPv0wXPeoFDrG
7j2MKDc7LsFE1Zj3B9R8pa9bq7fDIdihybfB1rBfzk7dfyOaS8+tMJ1XAizqWTXblVk5fPOC6i0E
WGpI+JpZRMTL2tAlIRrFKu5tj+/e4aF1TYThZ2pPz8N+IJjZsJF+ScU4ydLR2M/oWbf7KIxRAv3X
QUZ2Eqc9Ln4K/YIuOuweyAp1sEQxdqzUXODYapcalHfNw2J0xVpUK4P3irJNn92+bIU/K79TjDM7
6qlNsykf1IyLVsZDy2ONUA7AlDc2I6fHRK+VyzhMG1E4nYCU+lqDr/D0zPs0zovYRkYqBcKbeoAl
hPljHBmxDRmvdD7tFvviE83+kgCwvvAJ9K71W/DMClmBvuLs2mAgiBFtZ/pIpt+EtiG5wJFLRT3T
bQ+qyMWuTxyvMDreU4/TNuPjtvlffs21C3R1rTva2Q0lrLjR9ZGLT4fVTS8yrdXF8YTUY4X+7Sxx
B0GhMvEJe9YOsExYivf8yFQb+9TfZjKJO7nPKVP6T97uChnpuyIDVetoCJjQu/XVO+I2jGGxhamK
RTmee8kUvOMdce7rcd6jdJuhkN6UU8OoO04CZwH9NFyTPbTlWZbm5wrOCkdtNNFw9rwGBZ4sB1Q+
9Q+JTUfFGg58+/mlfeyfy8P5m5AfYUdRKD2eJ1yjHkjWwfClEpdhqFthwG8NiE4qMfsqU9RFTJpx
SFCBG7pOwttgvymWeKjHeaB7NeiH3YvHw7GM/3dZO+lCGyieR4niT9xWjme7q0sASHGm8k6swpyo
2bIdemsRPg1En6TIybxZbreFYHNUI/Q8U1wKT+AB4ZoFHKbn+PPdZONCJQ4l0duABXXVa4ExYtSw
YDVOrU4CIK+aGakqsmNHKZV6UHXzlZFdBoSNHdbnQ7RTb1GOC9b+PEz41dCN+KW/q3uBMxbc1J9V
X7euPsTeYXAIl3141hlclNFwPPYUxDxO90kTqar8etQS0HLe+jX0r37AiukslTaryUCOwDVzzFPh
ZfxPT40nreFCMPRJpXN90jHfHScdtymXCSquJZhsnqrqcTVwPMA/1OZR5mx2knmJxXwsJIKoc1hS
yPRJZps5u3YwS0uAlC6a3/eMr8ons5NRmFGvwD9K1KRWplqL9rkNGebjr4H3rl0JcPUXIUPmLuqQ
JZCOUan8tiU5ri7TUGgNK9qMqJWrr88lCa8D7fGhJF86Ai8Z77cdGao5fpHeQ/VFbJONhlhjT3Bk
f+zkN6ywHC6BALjlRheJs1HpzdjbuoIGEtWGxU0mIOUFqnEoOT1R40KS5+lIFiOtiG8mBS3FFQWO
dGscZFkzWspe7kOt0HZPQoFrVNc9NXroB/4bphJTPKPzn54HA19NkPWmiIUE8EJOqxmxvXyf2lYa
2FuvkICKhfrxPez0W9y0Q6a/ORbFA+Lgn540dVXO44kE26zLdKoGlik0GjrTV2N/d2BQ9wuHbEa0
ozSs9Dq+IEAOI8vkQcE+khIDNRJBAjGh21UQpTkYZ9gV+5BboTZ9UaPziewCH6LHlo+/vqNv/QMp
ciqH04ThJBzDC/QSVoaAayd3ASOGIs4Ko3bmm5HlQxWMmPWNNSKwzCSnbuPpjFNVSsD3ZOfWc6IF
ML0Xc0fEWsEONDLeXaegpvvRxgQ4uTxyG8gXeTWs+G1H9fvWqTlRuxmcSjGm/KLo+v2id9Y341ZK
NDGVrXotP0XqnNMXtntocUNIZGxOsS4P8wCSV6aVNmZZxxI9HMK1LZq8EZ+Wc5tb6LIXO2zHeWmr
0nJC6/DXt/e47ZHEA5+E9z21EOgUjSNZhwScQ3srZCU11I2odU8n5Ve+yFVnWVYbV+c+3Zl77Jjg
GmiTvZoP1cOhdwwipIrOI1W1wlOuQX4TRdLaASK1PM1H8eFN/zN+71uuWxHwPAycta4EvDsaS75y
YuistY+cXp90qiqbVyupyquAx8whykOn0vDlrE7/c311AVSK95SqqZxkRHSibc/8LXi/rt/JUsKu
B8JhgSZo85LYLay03qXlXFpAAjelipkFmkNjN7GgS5mREzlrMDSf12g5ETqqcV+0a2qvZ1afcpor
qj73bgQssEdzn9r48COucZa7DtZtNkaSxQHJUL/wll3k0qEtFBT1yrEq+lWN2YD7J+GkoyN3/vMz
s1kML2WGJnrr3CgpvN74faLm7yV91PcBQghWOUBD1vcUJ4zJbe+rIJhb/4Gfq1WajSA4mwMRRMdY
fGdemziT/D407/khx5IxSOM/CgjosGc6nKJmgrHj8an2OS4gnmgtBuUNsVEsI8/6d4Wg8NpKf3Ry
1hFtswgU5aCKkZN1EBo0b5QZo5PNRLmgiS2dNSkYt19RRn0r+CBYKdlBMGWnaCmhFDQntBr8XMx4
2y4Cr8ygw4YJXvRT0yUqwwuT7w/goqohTASwy33idqDeNsRS/Kj5jwIcbLsWClzJY/yZC0Y54E8V
LRFwa4hnV4mzFEqAusSfn0AY/9SBb8CN5xW3EgIBWI0jNfZeGt+Gpz/TweQefwYUkhs57/2n+9ca
uT3EemiXkTGkexvb+My5mP51TpjfXlpDMT+hjlfg6IXhzPLJIBDDPiTqUXWUAdLP7s7EZUudFVBA
rIRbWvEjl11l+mUclUnQVIGg386PolPkeXm30iAFCLYjpiCe7VP0GfGPGd9lsD4r/bFCYPvHFTch
0is2A/l8yr0brezCnYvZV6eJNUUxZL0omDb7YySc7I+t+oYsaYlfM0LpatrQ83T1Rdy6HbUAVqNg
XHdm5++cw/9odIrJPjwofQVOlNhlPeUM9aQiUvQtxslFEtTjA4FfK+wTDi6+D2m4jUmlxha2/btD
hFPfbCYKpR5hLiA1TN1jCmZvvnFXKQEgixURyG8TBGa1AfWPAMyzdh3SoQf8zKreEvc0qGcMIObx
LY5sDwb09ZdKSRYs86pEhQV+KC4iolFCP3hIkZvft7qZVCeIhNi4/C/Cm2virkFIhSXsgq8KrQeM
eRcmQazlQsWhLdPO/ZpOEOh9lWz8goGD+widdFtVUx8prlP9DSrw6cmGAtdmr4SUfdHXJvev8vzw
QbVMnlAOF/U4qQK0vo6FDn8MuZOX2DUCbzFwt5OK9NKiZotqGhSCzkZajajTNJxHji73Vk9cOc/+
1hPNGZ1VT8xavCb/i2HNIlHuR7ytJN6DAzWKLyrBa4OVNc9i7bRdiZaZd+GKVzHoKJx6udztzK2Y
z/hx5zg+NnNGAI1OzQ6OVRz1jXch3tiH3TakdwwXSggqbgeoDmJ5Kk/aG22y7e5Lt7EqXrcgPewb
k67WWQd2ArDqhgRY8cMm/Ai643XtsPWMQVttziy6bYw/T6n+xppDMe+DrBKQ9fiXL2tFqmpP+Isp
WegIIiagoclqF+H35xb2sPylZ7kcE0RXDM7NtC9RRp6sigN6oRD69Vt74HsYavT0kVJGvRtBQ4hD
83PyFWnRmI0KPhLlcRMpQ891sUKaTxbz/xdZyqWXiuC7A8lyJScXzlqw42BLyLOes7C2az4J1hE+
QomGPbgQD8ccAfjUaTbe4ZPOBtK63bn2UNk8fH2vaH9hP4Iq41hVVA64Kl4pzwyWj+r0r+K1ey/W
Wbvdgnz9F8XI2y4Mv2VKx+JqOIMRpSqBq5+a9orq1a1SMf6s0vu9YxpnA/tcfsiJvR2mjzd6hDqG
edNoyOsILfu7D0mVneLO+wFeX9MIEi/lgvt0D2As8JQdxes4iMqTeCXE5hhNxrcq87yn2UgNQzkt
5p3W9NO+LGxmtpr/58GtCrUIPSjO2pTeHIaXJ8yO4Q4KhS/dKMhU+JyBrXF2WcCknBlNawGp0EpR
XyeR8PR4bDkS7+Rs1x/xlbLrwFoi6dMvuIYEYgeoPqmXxYr+gwNMP50gUjrjqbWkRIt2hjgR/QYR
0Am53T4Q9CGHxSmg957+xaMQaDmUxsLs36lVDidNOekYPAZZWTTCYSu2WRTvXNNjmZbxAtNDiCUq
qPZ7DdE39WHEnl8+h7+bxWv55M73fkyABLHcK9kU7pDPAtlFlPez0dXEvQQu3b4AHGjCkMJAYuFP
eRvGGE6Wi6xUGr7wbQvUmO9HI4NN3wkW5OA9pGh7BMcKD3b/2dpGnaEMJjgJvjz5cTCsx7byeWVn
cm2Asl8Azzkaiaop72kQdFiuce9MaRrqteG27fbyExvtYfhetl24exwkMAg8i0CXLRC07cDIeRao
AcwgytBTkzxahyZZPi9d4FYFgRlhRnDidtTsUhY1DhInjyPwW70IVG0EmexGIo4LikZJedE6i2Qt
yGZM3Zo+llBwStRmvIs9Ul/cpRZCpKo9UnliXKh/Kd3Z9ujbDEm9FILH7B7OpMZVnEK2dyWjLiFv
0yqaWPKs02+fJ8sJs8DMOVMgBDYWbDGTbmUYPKjP4c6Jd7HC2SZ8V8JxD9l0t1yfgZC1W/Z43mw1
ClIC/Y0BfCPbnSxlT+tVyixIh9xYtL3PPUWhcSHSyZAwGRtPCwMGc9fLrvMcVwvIID0nbd0R5r3d
eUcz93Gj9E2JnzLGkhi1/SEibvUS5leHbjI9+Of/RdlLKK8eSGP+QZf2lAvnXA3JkBStCW93eHAq
+SAqa4gyd0PI61mN8fxm5wnaP4nujhyyiXr7xhm/EEgFL2FD2zExd8Uav1YRfSrBF/JsQNcC/KeS
wSd69nEbXqvbUchcXQmpswj12tRPzktIvhgMos3v2N86WQMzev9sdA3a0ZL9guJ+ZI/pXGyuqmF5
1oM/fi0Alu/kszeuMM0j/559LAA7/hCwYdah84GsoTJhMt8zqnRtNMGkw/Px44JLlqiYQa/krlKa
qZGmaBWNBznGzGRfcW5/s91ceNHWozmgDnhM2W+s8bnZMaViHNn6Hg1tb2eA5D7bqgy8DDT2BAIk
YL7zPZ+59yrjO8uAVMu2nL+8XqVBc+LEis0aErKc1K2z0ybjhnOCBTZBKVq/O0L3nGRMPshpMCIH
GKTOcQuMSG8bE/apeBoT2k/LQ61dhyr2z3as82m5BVFv//oBr0WRRkCy1f8HrZFsgDHBTEThhkcD
9ionW3gFTq4UrTTKUbWY1DeBgH+oEM8czh+ySvMEGnvX3lQpQISoVS2ZD6YNyZXrRG8WMj8sQ11Y
I2rrvTv1GEErJxnkiWRpARj50p19bJY3xRLs7GVlDaLkNOHhcFT4HURRweOQfaqEHuRuSRpkgxEO
D7R/W3cuLTdl1E7YcFAAVhIthL6MAUm/a8qJgvsybzvwYkxk2PvDnc7YaS6eN8l9/03Y8ohLxzND
3fAe8hpHg2rP8iz3d/WibDb66O6gMwM5oBWXuzxf0brIJVwUPo8yPi9ZU/yKWSKYZ6Qu7zusHkDg
nYb3u8VOAVi6ryvEGCLhc7GhDL9JYernMG5GMe4B7vcCK8hsEf0QPBaylDFUqgATFAkAJdSNESRg
SOUQCOG/g3nbhHuLf6Os+C6QhI8jphET4Su5LlG5uCIwnvvxUeoPNNB3SxvpFWTAkbVI/1hQxrTT
FAYpvNXKtSxuzm0l59V+FHXB47VS4RhDnyxaA6iYgv1nNxkf0Tm0PZ96kuHSLX6SImX7tYqSfS/I
dqUvjwP7kCh4VkbpZsG2R4/pPTSfmC4EoId8AUT/OzkK5tcBBupTqI0hASfy1FfZo9qKEaJZEfbo
TRHBoROlStzelyNk+xjByJpg2MnElvx8Kd+c8MRn1n0QL5lrWQKWc62Sj3rjK9/jQ9vs6+QdcFAw
qzFXXADtX6TQBOhWtdcrc2RdBx9uYtbLZE/uROBiuwGxTVi92RfgOGZCG30HSlJ6wWoKlbV1Rn5R
FFCx83pbb3UEUlUkkq4mJxRvhbSDy4x4Dv54j6xODY0Vh6KtB2fsq/Fcuvqn9yCjb2cZJobcF4rR
2nGvp5AxhDR4RQI1QXNJXHWMkFq4m7Q+oTFbwDXs6aaAHyx9hsGkK+xweyuDaaK8DJdIayzGYXMN
vSx/y7y3+jIz8OuKIsEped7obtibS+JO100xn9o/sPn3DAag4gJJO4QiKzx6ZKg9Ao3Rj7zA1oCU
pivyb2MHLPn2cEWIKugtnJ8FwVilQAT3OH65MYqFBzNk7J53JxU8cn7N71epgcOE5Tqi8spLzTv3
S1Nkn14T1rAZZbSKhhAcEnHaTTtBDVEFLJpeuHvhg9eI69VyIUdQy6155ggPapfprdP3emiVujrY
zZZ8ZvfSbpA/+7beNXBJwLI8lLgtJ1AhLq5VFA4cBvn6q/o3dig0gMVlEB10qU8nAdaD83LbIjMl
vjdwd1XJSa3cy3HTlGhJoWuvZQkGtYCerfriqkIhWWedVi8HcwBwAGSri6q3PSfFg7VAEo7hV+h2
z9yPhdMvGuoBPIgqw5WOCswmVlQQVcy5wx/EoI3icZYqsmUgnK/N+GwMMaU65YPhMA3TBHF6zGMC
upGbt2i2/PawYherF7iQmsNnGwkstx5WY6HRFCjOv6gdseJ9xSz5r/ymiG0wrbLaBr1Dn8B7Z1fZ
vfW+vloVBcMSOcgdakCRCk/epiBqEPyoy+n8ulDEUT368eLzElKCfgtfHeY8lC2X2Fu6bEjW/4o6
lZ6DC12DzbOGbEV4zXRfWew0nq4bKsPnPY5uOEqglcm5cIILl3HqGnq1vfoINbArVWPgiXWwquNw
JrfJmY471vxnhkonyl6Ae9H8LAp5E++bcpgoorxl0Y6SesxNrHTe7sjprnJ0lfpL/DXTRL9G7VTH
/oon1WAUgLGNkxVGSYAkqQPjzvBTy4CO7poJ9sVkqkb7pINPlaKZ9UCEFuKJ15PkPy1zd2IOI3tl
8JX5APU/FUVJa7uvQ2UwBGEYz0/YVfnpoUH2eYnWndeRnUaN5J6R+SZ0WAA8uDDsgG57AHiFJLvm
Q4VPisN/jS880wGj0eT7w+6kGegPFfjjdOSrLunMqddUzwVdd6ZaMuOO6p8xF9gGmoU3M0GiGKyb
8VARbkboXKoLb1R0vQrQAMQFwhHZ9t/nbf08hLU11A9DZe5Z02zcBjZUiJN4Yd8GQOvpNzPBBQqJ
AUdAKXuztGKUfQ+xLdP6G2jwi7G6uxpxNFto6bfUjdfZqZ2gnz15v8pvkfBjxPjq5wsUnGUGaMlD
OFcHFlufBLy3StUmdGfDuuettVayDx5QuoAxvHRlgUG48k10kXku6xVhSN2/QxGm509aURqoRECs
jfhThDjNn4Zf3AazZr9DusYfpmf+CF3GL0tv7QqN1FSRhRjHbQxZxDJ5gg42f47Wdpx8AZ7v57pb
2c0UiYdD9fozCuyjo4mGPSDErorYVJ6KfoG9pEHUPTxWqbnb2XJDPHlV/qNij5CZKRean1M3eNWu
J6eIhxflpdD5L4yb9VVKuBUjHUJkwsj3BRi+/zepEfOH0L6ZFS2bqi4vryYLtjBOGpYdEvcGdQz2
aD65c54fI6OBYrOV1F/RwTieFqxoOUQ/zhTVbQ2bgW7z42qxP8HJhgHs8AutZnvNR++a4vTDnWaA
BUN3oEhgBRqKNQFnNWel68wDX4uVH5AsFvDCp1v0skiakooS8ZVoniGPCtZXPR/lJyg93ECRFjg3
ta73ioVhAT8BkJQ4J3ZVqMwNezGZ3lRG/IN7amGOQfAbAZzPtKvw7HT8/33DZM02yA3NExq7Rru/
ZX5gVdBXg0sifldY/EAP4BQF0glAizZd4SFRRHD4GHdijHE+gf5Rvr7Y/cm4oIFVHSSSWXlgooYR
NKVdIV7iUE7mbtsqP7ySzACQOGRcQwXbM23LQcbAn1O9Ee1fYK5y37hFcUlf/wQNeFTcvu5/nDQc
M3HLAdUW/UtkjDC83FV4MzjB6TkyhldCNFHnfOT6BRAT6VtfVLD6JDP+009WJVFXywyqHKS9KXug
FIlFlfZdo3wSytzuLUXNmf6/NEk7hQYyg1jzEY4JqZ3JIKTuqxM78pGH2ot8LLHOhquVFyS2ZwUF
g545n5FJiBgp14xARc6ZCIN/BdmQSH20CLw6yb64kFhOTPJvYrJGJx+TJXLP1AfS/bSTYSESPlWV
AlMAGYm5ieSd0S2en9gIL2xoCY6CvAyt3LexSnIoUbqtNWxhDTwn82w6m6UNy6JJb0PMZZJDxyZZ
SuIY/vcq/2n7tLlGKodEELS6rpaR5scUXSVF1Mva5nGrhQXC9tFjL6Ou419HoGi80ngixbCaYkOa
0ns62MFMZQ+oo8r7RZu/oBOwRAgq78cVfePtlZzoAlt6lsEyYPWoZyIy+Pd3KuS64lfM4DsM9EHr
ap6ZeVCpds+hgkqa+g7t14oz9u+cDpuO3gemi/CLRXZzed4edzeHnymaKP9+dOxqRiMIkcLVi8yX
nFAE487VLDKGpoEgD4xF+mKaecRqVOEqnpp7KZW7huiCqnOWorxNO8Rrb+iQpDirTx9imce8EQUD
xT+0x593WFTZs1ju/HC7izj7OBRsLWzU1Px1ZHN8H18chytDPu+uhN7OZ5BELyqwmjdUJI3cz0rV
HX+ND5dmda0rCI9V9eBQ84EYKHq4KvzpGp+LZHX8fErZK/SHU48t+iz1tDs4qQb8ke+/BGkzm+XU
FsjFhdtwNTh4M2JL0Y4ruxOAUyIfk2YU+LYKCukuxIXZRP/aprnceATAx/6StJj3FKLMfqEIWAAi
bPnYmc0mhXduu58u1Dk8sQ2WWHh188gkazeWBd3kSdCxJVgfmW5U88dl9E8tU3Gf44ai6Q17Wftc
e3nKFvPLxZSEoX2s3WPQ08wT8Q5PLYS0WxBCS9w/LRQdmnBfLT3IxcCe0tqMzsgM6m13TjQqBxR5
+ABu2wHimMPqnxb9hi6R/9JCfSHCz6euup6FSDua5Yb5q6SnQW6Z2n7BvnZf5/7VXFaeQ9kgQMQP
Pt6pfPHX9y3yLPeGjMbn8djfNIFGbH91O5akTxi2Gkjpovm3bUySRvpw1FPCrajS9Mwc7AM+AuF9
Mnja84L9uOSmXj78bxpBWu4pKZyvz+pj0vvilwJChUsuldo3QMGRNDQM4TXAs8myzZ0tbUYhPQlp
WTWcPoiBrwOof/PUjHTaUkA88jq287ieDiR5P9tOOKgYaC7uLljtdLuH9LvVJbbDu11b0AMU/gTN
lMTrmyF7d5tT1+fuwNC26jG5vAMTr7CefUTgk3XHMTStGjZdq72N+W67zxkUZjFYrUILn+QLuAqZ
cgrcTtP/0UBxUPcfgEkxRMBws/x2PRTBDZ9iI5Ko375UPirM9LNfW6uBJBchfviPrKKIxlAYz3zv
nSQc7m15xnmre82iXUolvMOMmlQ/eBReSMHqSHnLeDm18HH7+YV/lnBRnP1zpZNC6tPyOcSoLQ1c
ynND3VYyVQkdDb6ncCWWaA1B5s8xwdB+i3dB8wojHyekOtnlgFq6Yi7Ixffvj9M00ZM8LvkpgXfP
pqubw/pjQSOcBAYIsLhHfxxwK2buXRiRcGeB1fAMZvLw6OyKt3s/QkUBCSJB+aLC/BSAN5FfT777
1oYsNC/7SwnkyMWr9psCAnmfHS0vjWpMRpq8tUcMlCgtDKIoZcrHRcY/+JdwcHYTnAREq4DFVPPY
cxJNu6vDpXOpXqJ6VBdWB0YN4uR8BRncalPE60+VN/laDm+rV1DFbM7LzHvxU2MPIlTjdzE0GKC+
zbq0kbnoA1dwazAUpXdqknaOPZ1DCck0bKK/yuL+TIgmva2jBAu2Zl3OyuBQggsJhetMjeb0PCYr
gCpt/IcYW7m9xcBsx2YjoeWijcSyoC4VRWdfQkf9W/N123kSOoh/Hq8qlG54L4rpsfKgna8FskeR
VLiE0Rsu7ggLz0MzXRpz5JmFFIbOjTXubKLAS8+k3IytYzrGpblihSojWnYcQrB8X/I6YZQ5GKt8
w5D43cn6JqZYvdf9XDYYZapD2jN1/sG6npzlfbeFMDewnFzUQGOmRJSqTVmbMitzjzcQbJ+/O3Ai
vFjVzoccay1BQgJeheavM6taBwShLSlywfAyFXFwkOVv6sAbIQM1Tu398gDgM1XZNtX5pcLAL+tu
ntOtUMQcKTK9Adzq6MEhhBhABvy/LjhHoz24944YE6+ta0xfIPvtE6ySGMx2dGCtGGlWcp8kQz82
+L+ghxE91eB/nAvxvTl1DHXEK9+FNv3lSo9wMLJrZB+kt1UILKgUa7EB1cYNilFT27f8tZVFvcSE
dSgQQRf9lRdMiqdUUIq861akboDmaWWQfjF6xnbN91tWduYhuEMjQNXnDWBh9MkuQJNuF2Kkbm8H
kib3e7QDgKEb8t49x0aSg2CC/jolATi8Gmi1YsrNSs5v+B70vyWBJf3Ki9l4Da0PgxJIrHteRSdY
QzUaOczyrMPOzz8sK4tDX8ZsZaEtRFbjLdSIgZB3+OSwLVpcLlEAqj5FHSGNOsu5vV3RZqyULz79
MXWwhy26je/SAYSE8ougR1qvOCtTlD1U+aX8kFPatcUYFGQl7qPoZjknm/xxTJ+wIS3ZDUNpf6rC
mbwMpZLnaPe27opbTL713CHPV4FnZhknt0hhJdQDqWMLobi22BpuKOUswvdzIvXPWuEV5CG34jol
F5yehWPBzwWy3nUoN3zd94VC5plWqX9Y4CS8SQDi/F55NnSudNR8AcqwXlA8jvaCqs2Qqg2qxsUy
Wasz2kzw/f8knyju0IVR5iYkgyYwFg9RM0M1fXoT1oEAnCMJM0VazXX85TFFh/kKEzjfbJ/MrCIp
XAqnUmKt0LOmYoITvfwEpXIrcZH3jT43/i3ewGboU9QpLsVwPGBJhxTwT4bwVyw2BzxXtRhPeBMl
5+h4FWCCZOhkPcy9yy3IjcoeV9EXUqQ6KXnhkpyRexZk29FaneH+F0NO2yXvYbB6lHYBZq9lZkog
C+7Vp2txUmyMGS5T1VXEqvk2NYL0/ZXg204/r4FQFP/S0RaA73snGDZgWa8Z96YiTjmL6MlnhZMI
9eu3j7Qtv1LOKcXZYK4T0GTvBTRe1iIK3ccKuEBOHVVlD9RNuVN2hkgmgJ8VMBN4nBRBQTPX+imD
XaJ4u+OxxVPGscYRICnsdRTo80JLzTYoXFXoMJJ7Q9dYlm6/8k1WlNnPrQnouH6oNjnpVT/RSPJD
6uUa0SBGv5+RK0GbBW3CtncvruZ9HBVGZviUEY2ommjBMnRSGNCWsVTofXGH6A2hae88j8sG0GCr
MWuyYUyQsHZHU+Mok30Oe6jjozzMUcLEIYafyRM4gXfEXK87Al1d1GU6F85/Ft1lomgmxutK/+gT
F2az3QbACi/INL/9AwE9wKUoiDPmalbf45Ul08SxDNC02cUYK0/vc9WpHt3ukzyWQAxzJj934b1W
obDZ8YA+fuXp7n8W4q5OLvBz2SB8YFTtxCUl1b1fak/NNF751r6eNbLVtTblrdre9FurTXf3ja1a
oUCQN/t01E4cAmlDHqA0hHAXfWjvmLJNw3iK5u52BmdU7hwyhHJwqsWrxMGTq7V/t44F/OFzF3qO
9rmz+NqXJ0/fPBHxxrhy/h5bmWUpg/OgkmfcCubqhDhF81fwRv0RZ7Sza8WsYT32uyiCR9PpRC6m
T90By/QOYRJOcMJpX+YiZAF6y5DTUIrXpsJQL+M6rJAZrt9/0NaQtAtIGp7VwWl7JLl5jdJ0USHI
xhSm9NXDU+Gkm/iMp2L+DSJHBAeT254ifrhnpkjcpXDGnxpWyg8PAyCLWMoSRlFvB5e6mIVeaG9F
rfJJJJhF1kH+rKiKfqrtxNqKwA6TInXJd3VRMV/eamfGWjYzp6WWXyRH7D2SDRSWM2xhirwmeofD
/HyQFHFivtfSTE3TCFH9gVbX6CETD5pq4BUgaUkpJtTFxiycC3bl7w4cFVtoZ/QibTsz5swAJqIC
5M/ZH64+U3pY7TEkY+4K0G378slUEsUMz25PEWhZ0Yd4U45sdZ+xQkpwcKllG5JvLz2lf1KRKkl+
/1WujGcHKkm7kaxfQfm5AtafiE1qrK1gUH8Yj9Qsd/y6r4Paz3f5wk4LeOz+d7vkOLlxE1yFjFyV
+M63jstSS46x1dDowFG8HzX5pGR7ezHxo+bnEPmL60y7+x2NKoDMvokvqWky7MCl4BxPxSaVS3e7
M5Fd7/2ICfGy9YhuJeDdTnpCkdK7g3sUUv6TvPSch0/jD9myCcZ74u2PR9LbHcv2PF/Jmeeddq29
Gcs+fvPEFSls9FPDoTKfKAyHK1eemKpbWsUUdC5SmTMvuRNdl+g8ujJ0d5wDD8LveRbZ/Q+34xcj
DicLQGfTVxHuiM6AK4aAUApS0YF/ZeiBfHEEZmv928ZgIv8ibEH+Va+ubssO8JOq8+5oGA+t/CfE
GuDTcKf5Mz48gbeXuelxAEMZM1f9AoqrscFkv5eOdiwfQJWt96TK3044zu0vgIUyh8unRl0y8lT8
izKGU90Bt/sWIkDi0QT0WyJrtXPanqEcWK1tj53wtBelxy3/AH1ZoA+bkeuxb5uBugl+s/kbDvBB
BxDSB9Groj8L/+p0tcOxyaze9ZVsgFKaVMWDucBhmyU9xYI8IRQzaHen0nCDcLKM6QGr3VZQ9vh+
9Qm6Xlau3a4YOH74ZTNLge3ADI0aOKVuN+Oeca/3IHgnsC71L1+tKFia+ocGBcT4S9nf9wez8ff1
EbK+8U4LwqY8M1E2CPLATDbQmg4wddi1ZGqrl5L57b2WwizuRreFKn8fwTc//MU4vVBh0w0s0EaT
hs168fCQe8XPIIDZJpDiTuQIYnU4x8XyZTe4mB5o+6RJhKCT2tX97NyBIHmmOygvr56YfdJ2NFrO
F84QxSwdAW6zxZZjkMMfS+Hf0HsFM0IROLeZlNuh+gwnZR74c5fUFmOOslQFD5kHoLV7FV94oRD8
BDUCZUWvchvLO3Zpzdx4dI9HbGWOGOmmAk54hV/uKjOLAnv3ur0ErTfK7bd+IrdJwqrm4QRxiDzW
BaUuHD3g5h2oljuE3Q14AZ1PjAqJIIIfsM56e+RgNChBgAGMkpgVIYKuG3jN1B+LgwW6aWopSCMy
znX/VjwQNSU6WQUdYeEvbghH+i0/24aKBqEzIQeBuYtzE/mDUOQlji6eh7NjbW2rTKWLJ7yvri/j
CgvNJCO+/TdGqbZmFjDO71+qcWKuGIF2SoiwfPioEWw9pGSVm1f0CgjmPmNUydQjdolEsunU/XNE
BQhw+DV9kCwJv4glCsp51Fi+CAR1VqiKFBLR+i8dPvpu6LcsUkmGR9cz8Qg8fI8WKXDPA0stYwEj
tGRNWEhgNiAE0culcqsH+MuayJ1giTWU6EsiFuveDCnzM7yeAr84oLRw31OKfmEbY0XyKxop87Y6
1Q7eNISh8R7UGdffAAYnnXV2pD/tzHKMrGE4yOKce1U3WM5jL56AzFug6P27fNdbRxzA001nluk8
69X3J+JIcmwAuY1plyP/nQ21yP7D8aRXNePN8ZzLSKdNW+fEwfDBeACI0KevRvh4byDuve6EoxmE
FuHpHR+YKpHNkUYIOFkjfD4LdvKuBGCpwWNNbBldQ0bBbbJnzKaFxDP4h7rKXJgol9q9FcgpJlQj
AOKObW74FR9BS7cbGmbEmglECk7Ss6KjgyddYWfBZSNxw0bwRMgfPfiuoOhhdQL4O6tFmIazdWiv
dpAGu6F3ORmbHj6KOOxMoefHjf/vZGY68BZx0P2UXt/zxF5qXDs2DMuA1crdhsjezQPdSMBbOGEE
3FaSYetoNXU3eKdScPtcos28DoLy9kDv7Ghxf2AnkS9N0vQFe1h9F+B8h3qtDPKbLq7VifClB/nR
j5NyqEzT9y23XCHlRI0HMtgCz/kIO1XWDAEznVYZ+0u2k2IXP8RBnFn7MKGySAQX01g26ydLKKm7
QjsQMYA+p4mLXb6SDXi3orUoc4eYOveA7vkDSsTBnA6kShxmSVfOze4F/s1ktp/bXMYH2iOVT3Rx
SQ6cbKzbXKR326ia6I61JDF5S+Fx9fcSX4aDiivZD0XwamIYV+88+E35N91xPnWpd057QXgBIoHW
HfCJ/k5/adg5FyPxUD4CG45cW7bdg7JxdbJ6edEh/fF4AXEwGQ7tcKhM04l2omC5XrIavk7zoyg2
cf/6f3pjg49Z+aKgdLR5AiGnBwX/d1gQMLeF4d4FzZFCVgRhx/p0uwsovDvL8leC/OuxPFvkYACy
C09AK+MrGPnB29DNNuzQhO0A5lhnmDS2o0i87YKjXrbvpWImolY+GS1mDlP2J+k+YeGt9ZEwHGp5
419SG9IRAtxMlvk5r1+18u8OblreQ25vds/136eq/ojWvIrDNFvmlA0Aul0pnpzX9UHb5ubsdhRc
5jU8xvVGWKt0ltpretN15QDJ6Q5/dI2p6FS1lnafIcbTNSE6KLYPDPK03Ij3h5S6Cg1/vANT3PEo
wE66ne21aQyrPU0XLPbVIFGJJurcIRFuDhpdh66F5r5yDI4FDa7V/+B0X083ji41wRuMDxZRYo9A
OFxtWxzu02n9DoZeJIQBx6fHV++n6S4Sn4X7mqdiIWdosE6l0/sEeoNENns0wW0TEkMTtopQGBc0
vVhEfmjgj7JFRV2viMo15TZSwFm/84E0+vcWdUuV1s/6Rrmg309Qn5jB/Yh5O5yPui9wBPFYtpD0
i5Bkh6sPNrUsW0VBmK7c4BMTpp1AZ999xol8nyQVFQcTfTG7LsWF3dCq9A0F7xKO2bwBhFhFv77m
eRy2ecbXv9cKtyQidubr8MeFFQqNB4MlFi90/0MlrXPzI+7IL+QutAQSjNVu/pCsWGho3TWTp+Bv
uAgK6upbOpDJNJiR0qU7Fm3lMibRz+3WPWd3ugC7k5f0mSr2GKx0Pk2bs43h5iTtXwCtf7TcSIAz
tVQCWl4To7b6glFHD1XQiLA+LwN33wHJjtF60TojHqIfh8E2wN7x/HS+Ify+h6zWK0eb7zr6TkNr
WeHYJKDIA9u6nQRhJ3L5NEQzwsVSLXetqhHT9sVpDFWn5MV1z3F/MKeIlANP3JC9ob6F4LM8QRyh
3FK24fklqmQQ3lthz1FfdNGuetGeSdkwRuunRFRDOG6xfuyYYU7yxwCE3K/kQWeL3zm898VvCjEE
qh2kxNZGIxaRzWNvRpV6KzeQ2uNlzBtwiQwa8HkZ3LdCpDgbBBbrQLVws7xFRI1buoHcv8c/oIqJ
yveAfSQm/fOJgsLMSCEao1uHsqcOz2tp/MzjGxKXJ3ifShTIJWD7dIwBeytMFpbQ3K/csuKm+EAv
Ju3+7WyT1Qbxcr5F59B8MzK1s3HRIF1MJaAXJNjjV5P9h03Z4ZBfNbDsuhr4ubRuPZHXngTkv+6o
7jtpI4xVHdbsK4dcB03IIcr3kovVDvRjfPJ6k9ARwBflqS9ehWjgKS5c7q2oQbrBpQ1XKPH9uW4/
FMK5Cm/OTN1hoFvLRvK/ptJuaXc5OQ5rz0woCSFV/SZ1QYHldal3JgD/D9vBNRaWSmVIPq3CoKOh
2QqolerdcVw5AYhh9aUjPdvKCgeheEKTBcjdCgl+M151otL4Wv/WwnylkXeCbnqPC3StbdE+8nJf
v/kvRWh888+sG7FIughO6ZfHYoeZaiVKYlPOA87vMM/DCnXy/2Scefs7OD1QyFjBnKeIPXBN6Wer
DdRQovhmj2CjFVWFZDxDB5n62WZYOkBA7mcybtVDWWcjEZihPqnqQPymxXt+jnKqgjMxCRdeLI/i
RofWqtNHd107MT9lEQvHLAMxUGjqW//c+Zi5Qcyo3Z/awZN7ieqbC+Kt4dfvPi3nMI6hW2Pue8AD
IfcDu0KlgHgrR4URNdHMPqsBwiiAI2oa/cVooItOQKQ5AfI8Xsrl48CwJbmRMcATf7t1Qdd3Olhc
GURNDzhryFHvjd/lYGqjg8lrSFZJ46aesVRl+i8Q9YBluqivF8AaWJwoPbjua+vQHh80ATeBzTjs
q47tw3zr3/ihtBqzXVwSxVC2XezTHGi8I751ZEgu16lam8MnVgX4wTa4/91cxGHfsRK2deGlAR1C
zg/BN0nPbI5KtShp+yY5xkCiB7sXvAblVdF2gfXLX0ML9FWRcQ5ejr2nzsk5G7qPAkkHrudggMDq
1SLOE9UZFKj/a19aVC4N1yaPtWVWHVNCrdNl2YZRUfhJJon/6ijexPuZmdFWIcG+uLuR00RDbNWL
VAwFk3gljYVN6yK9FBwXJUPc9EsRYzK0RnlGWT6dti3S+o1QqH5gu/o1IzV1cvQ8g9glkr5TJ2Bp
xBoqDEnOgmKWNQXRGhD/pmWqZaquRJDYF53aAe2zEjyP10ouAj0n1lLdmO75q43PdDrhsU7WnJG3
9QDcjpSmbdsXS16RaitI/LUTc1t6FpUVvts0RKRylqa07bQh+D3fJCdfKSTofjZYd3rGOgflhxAm
hBfHsL3MOwD6HdOxQd9xRj9ej4yDas+gPKBQ5eSXx8RL/cT2o4XajVjd3HdV/b18FY2/ZuISf0T/
GJ5HKXNJdpRWTGyRpyuvYXgR4AAKn1QGuyPvYLp8qZqZlsbL70xZP9rg/5fuHOcjvMDmqz4tspnS
daPq73lauPkEOsJNR4ivNCMX2aqXqVeLHuS3vEzwQ+8urraXiB8o7AIaCY6vsWCFcP2nfhAO4nxQ
Z9bY2jtGP7y7DTtDNYW0PP8gkXjDY/dK/66Z70DS9cbG8KNwFncmIkF493hoqufFzOIYxPfebmRf
PjQUvnr0lP+VYn1lzEePeXGty5sSPOwNpd3Oj/biySz2S7qZ52irz9C03lNST+AGRnOwjqmIvXMs
E8kNgikAy5ZKmYUg1Le3C3yCeItnNHKKEfX+2vpY79b1WXUp5fDbU+lNW6ugbm+p0DZTLiC4h4T/
ic1mEE9KkQX7wbomAkGbiuK4rzAXLToGy3p/3/HqLd1fAJYgSLzJmcMDV6zLc1oKjPPx4OjMX0gz
ku1Bb2AWvHwkitnCnnIrCInQIQda2O+sZ+hgk69DKymUSMXmywNnRkCdsbfdYmCitm1F6zurQThp
oJ//zlORn5cvTMycRPrLKs5WXJeZ3TO6PnCwe/FYWBko0rPnfQFJp/0ABoMbMnhZBpbsbDcKm9NR
kAhb12rvrhJQL7ecbIVKk16NKfhST8mFEzGpGFEkhAno4M7OGKjJRt4GodM1Q/1Kr1RS+MfiBz3q
VicoHK50cFqiz85IRs42gZpdVC+5XumkiHqrWB0SgJiA2asSxWc9el0K19I5naBWnmqBXS727zhj
PNVEWjCA+bELDVmwVuy9hjenbHmCejyOuZELS38TaRYXvTP00Ewz0EMyGzsx00/odzdlHGBO936J
dmde9EwJkcNQeeIRCS7g6XzsVOe79xHzSrdKhgFfPBJCvLJwvyOZbFQm+bw4xT9ATAC3vvIWGU0y
jHfB2aQ3uoxZMGoZecc4FHyxi1x5jwUv3XNpAxTsdhlmiA2+64+xkYqEygiufAzT21V0R//Lp/Jd
pwdbqorukrF8ki3XEQgonk1xTJOm+gDg1VCNKGe4+rW2aYi55A626uxQdj6kcumjjghJnm+0b9c7
AIapsP10nez7BGxUwbtFEBAoMzolOxoum1kyFajoRnk2Tcy2ywh4aEvp+l3/LJSHZM8il9SUwG87
67R+9mn3PYuB5TQjg0kVd/l9d+RBNZWE15yXFetJhU//IKcY73XL1JV1gqVNyiHAOJWD10NGOlA9
L/cAVKZPJkNyva+3f6oBTA0vKlk41L0OjjQyXBiSJ4+zogdAlsYUhNhSQJjqykr3ljIOYPcYiA1M
muKtEXR15kN+Ps7yW+er5Thbjwv5ivWUPU1JIam5VRXc8xxwB/4R4QuP4vhTNmDsTTHMWnT8ZuBD
6yqlzaaULNCrfa101RE3BQmTCw7yqkp0SqpaqJAwUJ4M3WwKxdcD9LgDXZks1Lu9WgFWok+y72sj
dXNEhAl6gyxWz6w0r76lAmtMITcwqTd35LQbUKRP7L8n6Yf10QQxp3mb2d03FoPuvZMANz7FZJJg
StRX0FAV9tnY2rInXCPQYVX3AZXDDhM4FGEgjjq8nAEJDnDWwRGZhbWKQf2VTQDtOXeg4ha+n43/
T0rkYdJPP+STGMwle2WEoJNhTXJkVVI+GMvvs2FuiaE98YNE6bUaKshVse5giHM9gohP3q6lPui+
XsxqsnxpBHa14KJtUq3lkyfigUbYgFA3H6ZK7KmOEuskBzFlZMwwu1L2+sowZ6QvTuvUPAAC4Zgg
Wjg3F5OkyOMSiM3VXq9HnfMBBxPtCA6LqVm25ErwTWcHR7dSfi0IJdujlvkYtca+rw8hdPtcfg7F
2XmatcrbgizJpTxp4i3XAEkdt4V5R/BYWgpx6FFrd7wuswNjHJVwMXGrrUj0thwfCdTOHk4zk0EZ
nOJvFrtC0CalankSRyvlJ6jjK1OizayvLfERu0ckpDBiyaxrUesqIMeEKv/XHuv4G//KT/fdBKnc
DF+hNmL4GQCNH+Tu1Vz3QRUD1DY5c4cFQKniyH/GTNojyL8ble+eWGh6A7VamjJl/gqr/1Ge/Q0R
A78UVM9lWBQkOho+g82zroivIfGDj9fb+/zA2UNEx96qKxexkXiqMgOWASXKg0UGXp9TiOjKM+6D
Sr+UnjEF56OgadpBLGk1qABDdIjE0GJG6xgZ7O9watwGRc0moz0vKC99s3FODScsUCZT1Ke5j7RB
VXuVv4CSmH03cCQ7qA6ZsIWrVSloKPup6iopWZS6DndDv492ruyb7Qaoq9AQkn4OG1ZU+a7tTuNi
sB3AaWj4aCrVEN4whOzMuwbEmTfAvQpuoZmfcxP+gzRm+VtUvXIjgbEqIgSMkeBjdFL1Kfp8Hbev
O4+6UzEqgn6WD32+LPw+zTiJyRBczMWrbyfsH4G/v40pVApvAdjxfD+q9Uu15wTI2MdpAPt7oKxT
FPM8Jtp9d1+PsYj2JkwWfLrTbBJfDlqewVMwOPy6Gt4U+bMhWGxqrlLQRAQFxfHBoiVV1NiKKMqA
3l4WDKAEaPjhmLTvTVcqXiuU51rxz7txUqznNV40YXZ5hgYENqejxDCEdoJOGc2xiLPDGUAMSra+
sM/UTjYC6CMPdqfI2wm4foMpHrDPgOou2Ofls4TYOHgUFO0d1Vzk6XNunTeC+pkswyL5e3wbX0jM
LbEh8wfkdUUQJ9f5SuEvQwvZnNmzRh9ca9HCkIrY9ZGG7cKoM7mQci9NKLW4p3wP7yROErMneiGy
JTAzi3bWLcU5D3j9eth7j9pvkNe7/aVnwSgoStSDi3cRvAW5jtHMyjrJ4KNqv40NDy/FL1V8phKi
W0rNOHo+6gshMxJLh4JNJ+kkozOEbYY3ZW0CdqZ6yen106KOpHMbtiSHoZ/U8BB7GFnTBCT/jea8
JD44Vvcf0ANoOj86Z2BKMHGd4u5Y/jHzpl7XRNnO5sYhxlRRupag20znREStlyo/CtEuQLAQ8Y90
V/oeyZHJtQJlChDKW4cCvRYek1gzxurK3Bv4kfuHAZEVJaT1HBw0624/Yg+6Cc34PDw/CjmVSnZQ
mtr3msWuGfn2Hz4i/a5vxe7wvveHaZz7oDKdEzQyPdFFUGCW/Krl4BO+W1Bs/z74WUY3EpVQW3Ic
KXspt1m0m9WaPuQ9jEuaFTgkBt+gnLYAoJ7p1/vulj2488xaZwbdjB9278nM6uuzBo53rSk3v6n2
1DTW4mB34RM0K7q3O7lYLi6hqucq8sw3P7/ImPQCPVUVDjGYAg3WoBhBZGqnwASt4BhhfvOxWize
wr9YtxEja9SqygS5C2lCZ4L6zr3ZiPLR/MzLjRzxIREcSLkK2MbfrCaP8s5VDvC+xhYxpFDlYRdS
oz4D9UFyI0cyN65Cngz6xXtpvO/HxbfsvtTLEnqyJkxVw0aM0aqpu6eGZxO5y3vOnca3X4GY6ZmK
r/k0chB4V3wXWvrlMw7SHWE35Rzon8TGdkaTDq0FWRAco/FnKLAtiYwzlS+6xqdFvQg35Z62gygK
nucne0MXSX8qM8LUxIbjU0gKL9bA4Eeg8uCkV2aVGMNGs5DFrbIZPsJEMMIdPHOgL5Jf0q2YiUOU
S4yWljOAVjIZPxBE1MottykS/ytQHRkPCe8mWTEmarmm7X6KRGGuATSRntT+nb57PKhMx4eJMPbu
Afz8GeM9ai29T2apP4djoiseGkiz9FALdl3y1ZifUuuoqSiC92/AvlS2MnGJYhESCJpL/BypHqLJ
fSkDeGu3AqqB+Sb7UbxalDnXyKU0QalP/IXeY1Y1qQVWUSO7AuZlphU4J8w6yNvDsTgQ8E26y/fA
149Z960vM3hgEvE+Cvfhpm9/EYpxZbcefOVxroESdfacih0LaH1BxOj0tNliO8ggFQvMkjhj15E3
UEtTWKr8V1K+38yUjoOppPNzhG0OHRsjjqH5EHNKZPIXgi2ilNWGf6b4Ie/+EmDIz+7Ja6tKiqX7
ceSL72kO8KnTyM7FPj4wote2AQ6Ak4CuF3u+wBKg3nYwpg81Lf8WOSGDDh4mihfZbkgu/Nf1ZH8I
fFVLUyjEHcjYH/BiQ+9u7IwnVMG6VtvFyDA71yO5k2crgVDsNPncg/Rlcs1Wk1fEq8tWojzpQ5Jx
xPW5pOFfkzENqHvNpQ+hjxgcEWISiqUV3i/8lEIa67t7XN4s/s09byW3/P5aJYe1KL8dc8iFJjLp
UbbM1lm9EJHzMGeZ/BvMMcM5QQXr9PZvbtmfdqGpsBGakWUXz6muMuKLoYE/3d/EqMRlTy6VypWS
ATjRx4hrvSEXdW3OAn4ONzZvWaIrY8AVH82MfvPuiO4oSkjKH/3yO1KdKXK1AwkLzlGXmz23oBhH
JeUk+VaAW1q82TlIWAX2eUaEqJelsGaVQAUY0ycRwAro737rW+82T5wfcsc1aMENRTx8gESYGNyZ
P+Gcqou+Wc+BaxzxH4iPE7T+y6Ej/be6sucjkdot12OH8KVeFvHIy/5k/SbewLrGpgQVvFyVbky4
EOAOtD8U7qnkXzvrms7og0ndNMpBDkLNjPMBmvYpdVcxlGE1WexEEwz8/mLAgAdgjRP5FzLOKS3Q
1I/Sptzqhh6R/RpvhIh1xflUb4wvFtw2kTEUM1Q9bWtMXg1iHQba/OEG8BVw+ssaRUoc8thynhTE
Z9EnP51sNuCGZvyOwY7o+ibOAT/J19r6ISo3xdNfuIEHW4YDcWHVPdgc8eVKRf97vYZFGYkHIQoj
oqWQNS6NYtkm3FmJ2NG6fg/IhGa70vLGQhEQYUG1E12x2qoxSXE78kjlTCsBN9ivIliTgk357grr
nBdq4SXfXDd0n5sy/5leCt46Myg7qOCjyWMZvns+/q4UW1xSjT/91Diz5XlPQ8YL3QRcEu/K7NA7
kg5OUryXkJXDyyx2RZt3h68FB00ZwuLuFYpqNdzs5b2Jn/sKNHzYtlbTMJQvaj9Vsi+tdTe1Cn5b
1ULHrCTDAL3lxhEeUo2i7EeTzLKc01gXbCbviOaPdsPnSkY8Ut56cnSd3sN6HSbBgMPivfDxSqlU
v7v7PSrnF8YSVjatqpxGqcw+P9DKSuFNbysd+zTB9wWfsYSw1PywurtJsYMLZKOgktMtmQDsfuMp
wmaNz599nfCUUVdJ/rfGZv+CubVsb5IAHgTbOoqnmQs4UFnbccQpcpbML0B9i2+8WV8Vs7jQau2f
90Dvm4EGs61nYPSwTCedcqRi+vPBVzb4ApFeXhBva6uoZOaMipD1bXTQ3Q4ofq+Kb6yJdxEIj0RJ
MDh/dul+xFB+kkZRhdAwrEufsp3g4GInHQ5nv6rYkwe4wuj7r2VXNuVG3BDft9ugwl+GqcUWC2EM
M6uwqwvW8UBKUqOAc3icbG1+1+I1o1ONbUFwTJSWtVIFDroIaKHlLubcd+ipRBtbOSuj9FMmsnjm
lItpHZm6tP5BDC5vtxqU2qQzYLOMAdopl95jQhwmI4GWzdtncCwqGhlPdMIaW0pOYy448kojOoZP
++bUjdBrpkY95K5T8YAI59dTdMSzY5nKbGrBLNyOfYkX9doM+XDWZ5+fFuPGuT+//7CN1HJYD8Wa
4TOczGXFONdUHFtFZksGGqHB57HwdGWfGQLmHX+DVlrVaDaID4xe3EwfR+/m3SFun+zoPVWdKXF7
4xeqlCY+bpZXXnyH1LVUUbn/VYk8GbCc7NrmLjMin1FTto87pESnbPmh6/TLrSiogFlc13Q9XoK4
AskQwKJGOAiyp031k8lgZY7YqFvRzjn3NOU06wHX0CrVG35+9AOsDhLOUfRVeWKBExE9rjH2e8oK
sKimcAHv3Mn4mMRMT0X89j5RNGgX1mrL/05aTGGnnkZXdFkRL9sZifqXvUI+a+j+49NOmyWBt/ah
XcvVJSK05VtqX1TdgR1fe7AcJmPtQJ+rFkRHfpKSsPYs+wti3ciFI8510dh078tCmaWQKlZmO4uz
FtAwc2EtuWrsUUNTJdS9lxuX4EeUE1hL5iZvmEylNurHkRc828hGSAaDAl2Z06fU8RcqKA/oB5zD
ogsijJsqLnc5W2FudiPjQbRG8ZXm3JT38RwrVKHAYfFdvb0vm0bsBwKbLPatEUUCDGEVgcigOiZy
0jKQeMfWltpg6CAHsL0MrFKRcshowpScRqJ+UY+ZmvJ/6VMjUX3wF0aEzwOMhOayXr6N7/9v9oI7
AiILvky1O/IOKcsyABudJBfavPeuzvMScWYavRICdz1GCJhekHCfoIaomsuivCm3NklOM2MxY4Fq
ASmiJa9xG2EOTS7q7GFMKOasj0POjSNch3Hewru9IlGl2Ks20xUJL8pd66ruA5npkv7NQ8ScAqTQ
XZC/fXFhXjiHWK0LVsmeDt5/aJbMCiMhXrL4XFMIcbTt5A0NAuLxsAs23kcs2vQnUkxm8ptOz9t8
ISJD0LphVUUpzaeF4N2s2LJ1PccstODLvUG/JEzGwmZKnRsfwOkbtGhTlRHuRIk8QxWInqXDfg0r
VsQeitulV1xnYgf42zRPYP+eZsjakepjYdxbpsVk69sMm3wgErEg4z1yz8QHR0Q4GaUK4Kx5qFRD
+woUfpmWDGPwZGTfkRKNHY9eQaqZJHO8M0dP36B+mU3790O/5QAq5jidU7YYmWu+IGUYMVr5ksD/
NqdrsU0eyeiP2qD8Wo83SbY/bFzsMXE3EqVrk7MSVlMgWZN/uSGcivzY+vaWIt+JbeTiV6Hykme2
iqMJoZ1D8t8Rv3PT2v+W3nfb/eIEcNSLkaxWG9+P1mn6LWGUBgHQdqrDTidSEHBAMe5rt5TiIEcj
rJJvpKy2uoZ4/zln7s8Oc/t04wqmr862rzzYdIfRnHWoKSJv/tS53hlZueb4tRuAkE4V0021jqS0
yblUPZxMsJDLsP4aX5ajBlkFtutvAOgemZKqEN0PcUh9FREX1hYGrYZ6uTmCIT2T0exy39ZoXC+A
1FEZqmNoDMlIrvaSX9jv96k/TrHzbCfAhbVPhtGXg1tmqc8i/dghgjEvBPEMguaXNWd7C+4cXrXX
o0FDdMm7P5Q9VK98X9ygUBHf/vZrqm8VCMwt9k9dZt80CMkM3G0vFcktClk1RyLvMjH2eTEW3vPs
Zl74KzEJWXC247rGLXxehH5e8pbV1wy1EnafwUHN4Q9CKhppUDAmjL7hGdAWiUdmTAhdy49aLtLy
QN7RlTs+BtsgMd04o1m/G3cfmlnLguTMVf9TK47tHHiizdlJm8gQ5FzRVzf6WEbVloCgm2Is720K
Q3RnitPhCZJpLYa5LSjSXY96XwNyt9t7gLaXZnm7Lt7Abcvuzb/G50FuDuIfovxGrZ2SpFqn5Kxy
g0WTp/JpoW1qmP/voJYFNQilVFbfORr4Tzibsd42amPIPAq5/5/AMszxxBdot9FsnTfvjPBOd2gy
aM9HNcVr/5MnqzFKOkzF4u+orpmCKD1Wux2dX62UHXwo1nix3QQgFZ3slVYew+tTn+V5SQtjz3XC
NvwJCgRY4FSyhdorY9yMEWgo24Hfo9ghhO6Az8dnZwQ/14Cq3ElCqy2xuV4yOdVczKouFqlRpJkP
EmhImjQJ+Yo91Nwz+xUdz0OpcYili8EnjfwLhE1UIN4vJGX7ce8XMfErJVIw2pE5Sig6N0qQfsq8
baUMrzBn24lh3Y1ktBLrNh9cBtpAV8XK5Jw2s4uB8oju7Op/9L09QhJRT4IW4SpZXfGI7YQ16R7p
8bJTao8f/01h9Q3v4waRG/sShl1MXnhCgpqFFMLA6ivNMv7Ka1mbN8cRYHXrZltb+xMPfaGNAUCd
m8LxKAnbHywSyXP666yR6V/lXXf+ZTEI3vFFHG9RfoCUWBlSr63SmuUt+NRMa9CsQFMhUgKV+1J9
QWyEHfiCJBKooY3LdPl4u3GWou6RDamLrwvxu5cFmxeptAxz6qkEB6U4ccSD2xapOX+40c3Pp3n9
z5NfIknHgdc0lT9D7p7myqvw9aTApFuk6cpOyfHMkVaWt4ZWXlUTiD8hZ2dXNRbWQMw+ykVGHmCK
rOORDzhH8HCLuz+txV8ol7YlLpR7GUIk8lYsZWhtDm0aaTciW3fUjQM0LlWAbKQIKh4UbKWCv3Uw
62sPm3j0Qml/zAU8r8Kx+/GZkQ+FQUfJb5DaDOVylbzX/zdoVjf1cpUbTrWvD/gS59MtOVdkzSvX
hTHhnW/n3JqEOZPEot6QOibMlC9aAve5asMYHzAfCHN1BX6IGmS0AQSMkZZJasjWc5SLJdPmkoRe
w0KOkC55g0q/e160xlHL2XFHltjj/Xmh+25OSSRJC0xsWKhzXJI/vLkLi6XjvOM4S3d+9O9YMpQK
DXsmzZp/BfCe5o7iRNymqJT1bA9QAvUdP1nb78DpXernlgUQZMDiyU4vxv2V/0VR6OT4oJr4nYrQ
msGnsgkG888eqUQrjdOzNlXyRJOzY8NdFtxDPO7zY6IOnAu+MTEAatObx+LdYDgrH8qJNVhnlB2E
nTOfua3BTvTpyfDdwX+/aNtHftfYfXDaKdFQ3uX/oTRMI8uQ7cmd3QgwBh4kUfMnJDXh8f3+vGl+
U25tHNWcnnZ5GA7TYPFSfCr9ypUsX501k5E7bSNgw8ahC4qjx9JxhY/tf5hmv9CktaxJz9/yRCMf
woVQZOZfbGt55v6002PChvao9Boarr0M5vYuPuV5pHi2THLuNYxwYNLuy9tTwBpzZ6N2doQqu9Y3
L9EWLelUi4qdYR5zdJXAGzPAtig/G1w82EdBjYzHTQmjekxBpe4fELzt3iMRKmUryQXXROKD2QLk
vlpA08+NRf3GZChuklYT7hBRkBM1mXYbDR1wknlIFYEFmUSlXs5OonR2riaQY9rmPkpFXHAREl6Y
vIwfHVz8QFcnz//yS8fiFH3ECAXEGOhDCFpr9caZ/CxyEOw+orYGtnpUCOCicv6aiUkW89TM4cw5
G5OtKYMB/dcS6t+MA0qNOZHajAAS7wnMAW6/CJBbciQF+faq8CwjfUaFIzhdpsuj709b6SH81u0Y
dpr3wCMA12du9wrneJ3Y3ehyW0/eY7vuB1yUG7G+AfBpi2c9ycacOGH4f+39e4+Qm1lfp4hq+l+0
vTyU1hoc16S5llO6PR5R77jbI0B9QlAFWfG5iZuFB1M6dmzLR2CgY/ZM2UsIKOTYI9T9h3V8ACgj
MR+VcIxaXUdXFJDvcLJ8qgr929oLhZl2F37PYi35Z67micZjyZHfwoAI6SV8L6ocuHhsDq82jGws
jBn0ByqOhhEVg6I/PYFePamJOHQ31rFzZonPRRhu4aboQOY3xonzqrP0IeO8uv22/feeRaPS2SUF
6fOhOxjsiaE6rXfPKpEh/oyscec3Tp4tAUmsx2I4TzYMQ4VXVDFM2XTlyNiVnepZRjIVxsfNABjT
53iewnZpRsBK8Ptw8qlvSy7qFPR2d2zbTMuUQb+AUeT7RheTiWsTMxIzFzQGievW+NI/Dywsf/Fm
lsDhSCp6V41TwQJQDyycLzJ4PfrZN6TSIztjPAoz5aDJEd2Y+25WGYoNWbHl+Negv1zZipyrGJD+
SZo+NzIvSW3hljpHOXPbuz5bqgXi1EQ2RSDeXRr0q5+I7VFaW36bD+xqIpJoGKoyaE6VfguvIKKB
SIb4x8HUtbQ65Az4vnvRWAYjXaOTDoBtOHF5hq4TKFGfyTx50XXAahlFavDT4wAKz4UzBywBTG1b
OY/6C5ItqvffSBWTjgBKMbJb351YvQDEM0byQRIxZ/10L82VxMbh3gBpyoCeVWTr9Pw8wxOf+hya
2k+RY/5liJs9WC+Z1ZEGON4JnFFHLMgsr8MHloC6GmPGuhOXNx5vlq1Dv8BNqcfPDP4JvanfaCpf
UrVg1RAANegQZtqoctCAoW6dB6BThXajTeubX2CjYQN7jKlhVqlCPvMekXI+DKYcnqFrcezc/GLU
GNJpEh0mGhv60GLTkKaVvUOlE+uU6m7IUJWAUBo8yXgR7LrXSrl9QkVvBWddbMPRPVQmClnbD8lt
b6jH77r0SSKx5ojrhkCbo9fRT3JNwfVkr2/GdMwUAru7ASTuh3F/0EdZSueH26wLlE4gOv7jOaPV
nB+e4biuBiwlXZj7mkFgR6SVN78u2sd1v7Mm96FUPYe5ZtwPeO3+frn9o7vvhZ1FcDbmc7VdTX6i
YLtS/Cs/5CP0mR45Wtt3cO8w1EztDZIe8w6msDKSoWTFNDgFqt3/PlykoODOL7b92Nh2Om8jWFRg
2UwoE5VtYprhsBaGRUAL3Y8I2hnzjLqAIqCJkytgCBJ76VSGIYTjHLP++Rz/+WvvQ1VaZoPp4EKM
aIPjns7n6fPczaNzm9EvnS3agWb4UDBx27MOunNO/1fpqKvwsqoD8q6ed+BZQ0WhkApFkWZbaZkW
Dfw2uyR6B4FZqkyfkRMIs48UsZ5wh8k/MTK9hf6GSkO+KH7hAAw1gtIWfXQmFuUOpxW+MEwdTEm/
OxPqVt0LGBWkpr1vKjbOp1quj/ZqNr1qLkW3rDlB9wVeg20/xAaxOm+snqd/OKKwfjls8jaj7MDa
uPVGxnCqCRC6ZKac869t1dFlcTggLZAfHTz1DX/KchqgGH94SbIqa7QxnW3BKtgVhs1tYYYmpWsc
OWkYJe6G7YlRSN6QEQkHe1Ky5d8E3IRQmY0mRWSALp9KEZCmyA6/ZgEf9edBy8rVSBVR1qr2zg5P
Bdjo35aC9THQ/fSluYnxi+2dECCPSwrxp9zV2JPiz+UbFcxBq7SXZ1/6ym/VdoGjbAds9XjdFA14
Iwk2Olv6ibfnXY3XlJtxFwRUt/VdINZhi1e3+VRHyn/pDvLRzwTW9i0l56AaBkbBL5XZUvm0bH+T
PI01ZEU60t42Xk/jZrEL/yzoT/tSyHf3FfXfiAK0dN7c6/goMq2onudb79BYxJxlv35qO6L5Rg47
nzyg0EpbdjLxTgh7mXwiHDOK59diVkWFLPNQUHawduPbllJc9+FMykUS8hWeMuKk4q+M6gcTGJli
bcxeF9BHTKyXwKx27ZG5qrLqhNgeceaImq5l4JKqlORIz5RUkroPGBQ5qEcK7vrXRfE+UK/b8/YZ
fwsIGUGoNgiX51eL+aBV3CNsaCoKUTd2jm483pp8uJ6XUtkZiNO6UW5K8mF0qmIIItfVhz9egpkB
gXLKfEk2Rs1SpNO5Ml1+gfTbov3qL16xJfPZNVrTIm+Z/33i9Opz7dGZaMm1eL2UQBIMLDw/P755
dJbVVCVoI/neACBpV+5Ueb+uuFl/EqTZ6KWqjfo+9aZuOtfIKiScq+GY5O2K5XvTtDOZTqeRA+wL
kiBTcKtrN+80OCpTI0GBlBZgZFRu9w6r/duMYqW8zIUdIlBpmB5jPwxbmLLlj89jK+j0vmuH/vpo
Wa4EaGodKTM5HzJJDjE/HPjYFqqJDnVAX3pIPWkwBurmKNygJZCcG2SKpofSO13hCktSfeozzsdR
/xQCYBYoyj6xa+H6xkBZtj+vdNp8BMvuI4vZl9ADqRb+J5l56Z+d3L61p0JZCAIcDzdisZ5RK7AZ
KYMsyVFmdDP8NYVJMPmyIIcI1Fgs2//NpJYhOiEWBh7tQ2EACZGFZXV1O/JnbgPYbEi75515sInP
W7fk5m/Yyn11xKBL1h0qMeHq86kn7paSeYnhCqFBHXauSfArmtBJO7C/4NdWsE1RzwydljCw/KCO
KsymT7QTn3XEyTnJ9P/JcAw8bGt9S0CFqnoXswF3jriQhh7C0pUWCYnei1aTB5/C8sFEuQPESnrC
uUTxSsbnEWw4otpXDRhCghAta/eLRzEH37p38yuAU93UHj8wrFG2Lyk1QcubP7ZY78VnykbG0ANR
ONufKLOOhR8oYoBCCwPNcnMTJGFODh1qSLKgF38ictJK4IS1PNA53iw9w1CjMMUOwuE41Icau0R9
pbBEcBrZO+XYc3DbY1uFvqwimoODDeweo6mzRIG96uK4H6kLbUo29gpYeMcLywjeIJ1dqlLFxvWY
UMLDGLY4MpxuqNj18gUWkTQExez4rCw3GYvCwMAkMaWCxCCpmtXvGbRdB7SuoKa24lrqMEselo5j
110fDdKws9JCJNyQjbpuV/CV5L3mfVp585TI3w1Az0bm4nt/zp0GPrgoOWBldR8thBHVyvlqPRJz
I7I6hlhiVvWSe+bqkD8yjCvAvbGZN7EDhd5A3RRppuEYppvX4uQ3NzW9d/+NTyUg7bqHaPXIuirj
KoEW9XgeP6lihDXDPQkVxwPkym9IJmHHRvDvvak0wLg6AB8dl5NbaV5wx622OXYIZpljyXcFm2kR
51oxuzMuHsGNSL5Nr0ytve46ytJ5CxSo76pmniebzsdTkRpQXzQwXHi8jx3WItxEaiSxdyp8z5VI
9ncJXwLV8jsIOil7Rlklchxcm/HWkMiLuXDMdICEZnKZpnq7nQbQgRUXSmvuktXuy78JtreVaVcJ
bZbycZvotRpzZz2MylCbRiKBRNsaQSixyiF8JFdrGYwk5Gt83YMVdT7Gnqv70SmBD7fC72VRmoeS
fp75dMGJajFSi47BFj9lXLOx1cV2lO6LML1tPbQnTLlPwQ4C1rjFKoIKQgzj4rFiEqqjD8lyMMV/
T5FbiFx+k+nQ5EFIAxaqjT5QiI/HT6V1eKEloK7jrhNOiwqynUHw9sEaDvUyXdIClXEIeNXqO6h5
m+0Ogn0sYXTEUxkWguYQ0rdcpQOPT9Xh7mXwzLuD005Zyl6/Gw4ZwsgzEIJELJlZPpGH3jhR0Wfb
rosDp1x4sc3F+XPOqOtq2ucXts7IJsE6AfFt8rG3us6KB5LnT5Kp1yxtzvLsxohFSEFu01UIL8Xf
vU5H/JAQsF1Yg4I2VSVldTyiypwUU5aftAhaKmXIgDRvCrOrD8rhXZY7HCaq4HbLFcECMY8U/46a
SUAwfT5WU1S0WvvZIHGjn8E5zLVC1yFsCto9ELiiD4F2/1861ghbpowrtLRcK0dYm4qRxpUYNCXE
YKCtm1ee1xm35pfEsKW73g9lnA215Y6CejldXfLVFyrNHQDF32sXQEPOHEls2sdKfZAup9aqLjwh
FAJYflkaJcUuNgfnCRNBPyDMgrrbTEW5hXN86BngngA8ulanJFl9uvoQMFLm1tGj6syImn/vNRjf
JXhkSBYdHRH3IVDB1NY6Xb7sGGOyT1WwTY1gGlE610qUPSwtqtfFtCsYRD6lCA7Br7eChDlh+27K
AU2sqyObk8L+XUxRNOgWOCxOk+N3d/r9qoLwA5RwOLrEFOYEifx6CidLIXg/DfWFrq5FM2yR0Hr6
+Nv/rGiWffdB6XnwsisRLlpRqoFctiu9VdlwYQdnckR4OXPkhFFC/Mr/V+2982I7bUq8uRISvzGZ
0MBuaSOR5U5qh8AZkvYchmZr3JMD92i+Y6pNduYehyZ9t3H4JOTxVhZOX1V1MngMZEBnN7fvJnS0
t4P5dVQJx7mXw9yWJyuWyKBFA8julq9FkV7T4NmXA4yIJLGIT1Wmj/jYz2Hdit4SF8ZHhJHueRDA
jx81459bEoy7sKdYXoA5UJkCZqwkMlk5tpzgvMEifioY/sd6Y9ajMiCwwxXfVndiLdZtJgUuZcOa
LmnbZ3gOcMefgX6Gl8WSWV88M3yASk6smogsxNfOnVjwAggkIUTZ9HDL9D9kea+/0wLL+Wrxkg+T
BuEdbTQCbdHG/bBRNn82bPzabMjWnFYk+OlDJzR9Mpb4ic+LJJPyC7XLEVQeyv3VDyK6q+mTg3U/
XoB0RJZoWYAbtAN/JLnIyV2M/R4I9Gd35AxhPYIFrvCfKM+CPWMomMBQsmqzs67EPqQI0UK+RxNR
7yKAjyTpWnflmFdEBTD/pnCu4CQfKxR4wn+AQPhFqTMPgvxtVD1gja89TmluZ2hQCyjJW5Rsx9eC
m612r6gtevpLDFrRaODVp7udVnKD1Gt3TXxAdZJ4pmPnMKnYisF9FMgxcYgGztOg5Ej0tw2mA7yF
+F/6rwKnvEYOcBvC1dteowTuR1DGD1ESOpDd1fSGQDP8nq15yKHhNr/M2FoKdjYOee+g/1ski6FP
J+pZqYHglY75qp5WtAwAZeQpkiE2CpjJZ/N3zArBi+CT1432jHwG/VV42kEFM3VtG1QQd0/FCHjQ
Ry7V1TrKdK8a/4qrhO0ndYAjpuV4sZpBo2PqreqvqFx9ZRm0FGoAi2OMTWzIe3YWaeSlYv3QGKBU
O/VqkHZArC+KWKig+PMDU59ecK5LQ7cnpvw1GHCtEZgWgyteCBxfYFdGNGlEWSlzh/A7pDzuV+xC
k+LucBaNf23zrQNzos+I4lQs4+xsRXj7AXQZMEzuUhz2iyVgZRzgNoAFvZf1TkgKHqycmh0inEqD
hq9QaxbgQo6laAlvePEsjZJaDfAcT9mFZ5KjL/sgheN+SI0Gm/HeV6Wpj4U2RzUsT0iqFuCjqosx
+dyA/o6zglS12w5umPFSSQfbMeKD8ATK9zxdf3tbGgGKjUjySBnbrjIycCiUP7aQSjH7b5uKlkDA
fDeNq0HqLyoR9RxQZfvh3v68fDaOAceoOwORx4M2q9RaA2HwH81k+jwM7dGo7din4ohDqLGcAsnv
lHBDljivAMImul/Mexn4FIDJ3u48sqRpSrEJSkEVFtsQJDme8NkhYL6RWe8wnVmLtEtBbqOD8klT
1Y6TyNJzQwgyoZ1X1YHINPUdh33ElEgFgP98j/XdAHq1blBE+odcPz/UN8MbhvbuVPU94u629Hxe
4fjJQLnPIx70Qt5TmEXEF5FWIeIOUOV9YyEuRXcu3axd/ETYWROpzAQzlQoMi0SCTu1qAUcJLGnj
UKeA0I7eN7FsXjprAw4/KD7FqrSj91mhc/9auqQ/ii47pfRNh1xXeIkOjHolw0Od5tSm/I2+PlSB
mqOfytUgRKfe3F0kkqsazYXCEU6HHyqMR7d9R+nsgasYIWHHEALcdD3ndUSi6pvCwOw8xOknKVrg
zoQLm985Epz+VGEw6Nvki0B8BysL/7nG4NAH71slB5ojvlsVanST9FMPxAUBCbzSZVzDE4GcEAHs
YmVjUZTF9+bZQIDeKqeqlP2ioMTQXmGL+PebdyvL5awOZZLC6HYB68wAtYmTv9Q0HFQM3n7RkX3K
hC634IaTXHdvEVF4O+7+41D8Avh+pdAonUv2vMDNFCYTcJGBdGatvJHOCkuWuHo8A+TG7/ObZLr6
0WncJUCky10ZFn7B7/bPF8ytwT4LHXk+97GZT596SLR2m0ZblBCTcAZreVLuo7ot+lmvGwZ6bcYt
iCnoKjtH3GXpuI9gpkwN/K1M3m13/KMD4JRXbTQRP39rO7tDcBn5ft3y7PxzfWdNK+U4QCtSurfp
a3Msv0Lbop/Vw0q2+HGqWgz5SNoKOdMfYY09L85rx6bktt0ZiA/SbbnSyFFiU498pHZmB2wix+Kw
oAxz1dhb3aGpiurvuVEvbkVFEjSdUTEkZBkBPZFtf5Dj1rk124e82FmqumwByt4rkMpmbAIv9MP6
5kZZ9RbV1JlCnhFPoWbGeoV9h2wzLW5p6b9UfcLLXblC4tUiq6XjBIMANmXHfnt0XN9dS5/i0gcu
zD9hOvP3wUYchOO4ZYo0QTtpwRkU4xdyv1ix5Ue+PA54Y+rhV5KISMBSqCLVskFoTimLuLkvryAk
k+xXkwcNMx8S2Q5fjN/zlbo7O6HKmQgBrJNAB3vE7nHZLm25Z+uBNgBBHsbva77CeqPhzTqG2bzC
/azBn74kTEepvKNXL0MWfdLpr1nDEZOiE8hiVUlH670oa4hez4oCvakTnH7b3U5OwLfxpQ1CVRKw
JGXZzd8fIZ7uhxIIhiUjMnfnNr0eLpEhSqSpf8IIQfr73szLgUUk42fmS29RpiSA3D5wpsT4Aj6Z
dn4XxFv6Xzf/RsFdOe2DNywAWbMOANnM/NUF3oBee3kqNFp4J6jfi21vuEjvgqne97IpF8LaJFGx
nKLg+d0v4/Lq437cwjgnUCiiV5d4o3fVAmY2N4hZNjTYeYgXqwTbUn/0hnVHorhNO2cH3yqG7uwX
1By1H8++HpcF7BiaJ1x1Ej9rfSLfGDnBft9uAgu7JkwqB2AQwUPSBrX2xh/cnlhVyjK4nEbxzPXl
KqwYFCAG1QaMoIEsKRTOetK2P3bLTkmvWbojbH2pQGanYlAy6ecsLilsKNbg67YXwMAQzHlVyilS
DfzdeLVD/UufhA8dBPLgeCzuu1pwacrH7kKg1V4gVzmb9xbCbZLWS+veQGgao2dCn84XhoHdY9u+
Nl+va3/NOVfCnS9odZa9Tr4ah2IEhoRKNoZmEeTYAswdz1R+mB9YgWRYIyePnKiOiMU4b5ZgVlx0
3tjR/ErrBxv2Gr1iP9lqedTO63U0laiOWiUHlRn/LK7YBV2gMS5rlD7NeF/Bu2wY+Uisg34PvHbB
K5G5072uiIYCmVqfMxYElJUmy5oM69MWwUqfv2icLhalE7kDuM4i3qG8reZIGrcH6i3Jp2n/2ivz
prKW7HZfyK0QT6yy7ezqrRZvk49VOlOKuDsJQP4610uoh3cR7V+FOmoK1xUnIlHWY7Vy32ZotYZK
MASt8RcCPaODjv/XiqHqMfGBxZzHgDAKOWyx6b1U41dWRTL2sCamHVxrq5lbmQlliQAiTys8BbPm
kTCM2FO5HsEm6pgPY9/TwekA/Sh+OvMdFtzpKVcQL511atdbz50VsQC0WGvSXHwiGOTFcspXOLna
KGDo/cWJyU5VEO3Fj6eFLteXA/dgdvGTrZYmRPBMT9asw+jQhFbDUuJntPiSuL4TIACAKYNVXNZZ
e8cPANSokwrZilopNASPSUTPZjGpiahhNm+H8ygN6Qfr/TCrXe/G2Wu4W8czaQuZa7wr84XSrob5
80m9+z5YDD7/A0iwMWDBt690rJrKLKw/2LZIXqWigx5wd73VnVWSj/qhZX1idSbq7aPP8z8WXKip
pBh3QmJ2MIoTFubCaBF3+BIG0Kbk0QHkVUbEpba4+QlouZm8aurG6aqJNRNcypraMv8x92ggKIgE
WbKsUupljJaQkv/SL53iVIQgNQKcuoGX6pc2yWbyFXB5UMtBM+d761+XWVldvt1x6gcDqPJkIAda
fXu4OWHfF/2OYzcVIGZ+fDskMfaN6WX9uIqqikiPZlLlUvXqNwq0hQei2K+pajHOZAcHXj1tyrXr
SKTXDH09Pv032eBWCbJp7W+EQA6KXzeGD1psA8TaWYlVfxTLo+Hl/nUMz2ZEscWYucW0mgcGW5KJ
LEjqAvvWWlUHtNLzBB6YOYNZNEuCtTLrkRcNrTcE9bgr1OiktO9XcPWUmpzoP13kx69RkejsDTGW
fFkiRKtul6O+M9xBKsK2LDsDdpJuSk1sUi8H4GNx0XiUT0OL4+QoBwH/6xbTOVX4/i7ddoSOwsc/
79AQDPUZLOLmzSBqYW8wOB8lpCwtQX5JMzQdft0k/mKj1u0SJMVwFbB0xq3ffL7B3V54OVD2mPcB
+ZkdkJ4GBhQwNT0hVfPQoKqzDzX1KmmBXuaMkyWtG216Y4ZCLppHaRtmHNoYUM4FS41M4ko/zW/F
0P5VvaVxihu8f4Wn82FUZPDKXP7XtxqbHTD/R1G18RFKBK+5eeSFPt0CnvmLfKMOkID9LSDq62t0
47xNJS1bb5ZtF4EqgGBHnheoQ3AvyuqYR+mr4hni5CoGGUdpK+LfeRUf844vCi3N2TpqYGtQm1Ie
bsxlJ0R2p3DJQ+9026fmW4/tvsAF7AitSF1Wmk7A9jRpML1FcL/YCOv4v+XoH8PbhUgqZCM46k00
VRqPAeuq6NbPCjkMb5J1uLsoMV16zWTmudt2jNhyfEm5yr4XYnBoHVQ83U8xhbGLGTSIzJaCsxtz
0v3nGbPxMQDfpX4T7jPV2ydMZ+U8BO50/IVh0DzADoVeQTD3IP+QMWUQihplB2gmB3EVZW8VdrMB
xf+FPZ+P0yUZes5VRjnB0CR6vgeilH7YFqtg0fXZA5654VbMJAfVkcD9ge6y8Qpi2ziI/JCEW+Nr
SHe2TNqz2W+NaKpyTxGKLAQkPW0BO9pCzLPlL+SDHMwHmsRWaLeOMgtgWy3z0ZmufcT+dj8YVRLw
Fi0c+d2kpsymmlyD28CBKEb5lEeSQN4XrnalxxS6w5I2tX6zin4EPUP+taq3RmPiXYndgOEny5lQ
3RMCaYXSKa/4/BLEsMK7hWbda5F3xPgUJpfKj91kwRdan30NwyrA/4nJHVjx80jDy0mDGKWnl58b
OHOZp3S8ZfgeLnpYOCFnTZwaX6lbd59MM1vOwISXRI75xlcJr/x0tK2M41Nd4HCOA+qacTQEVcCg
dhsHdE9QHK6LDPuvDT/VPTf7jXRzcGAFMY3uyCOrrhzjR1hBa8BJB3S7a7CypUA//ZNh5h+Dk0JO
b+q0gyJz3F/6khehBRojqQYcPQL4T2fz8dDFJxbWph9kd01xGfWdZQCfJwJpn2k2HBxmPyzL+zC1
nuI/DxBszCzjL5TzJAi9XFwyg7udBnFz8vKaig91ErCTS1bQflsKUyD6twexbqGSixJNt10fAdF4
hDuZBH6k6r7gshJBwF/USgc7yyu5GUb41SrVdIvMeRgLMK7VfPAuRXFhK/7IlPPgsC1scdq8QQWi
0uXbcinpVUgAX/5rVsRzW0ruD8z/gfEoRdrspr1dm2W7Do4FEk7zqa5IljtRJesx0/DKszPNZm6w
GgK+DzjG6XFuYlUDs9JKEYK/qu3r0HMr9ucoNH33+4vsRVNk756fYwx5BZ0uC7v+DyiQXI9DbjX7
buYqeJk7ZpjuN/p1VtTqE25Qejj17QKzJIe2ZMv4wrvduZxIqSi+dOQr7HmUBbPML8I9zTHJrulT
lYKYgZ4DkSLGijbvBb77nHD8rXAWbfOAh8qaA9+ntYD1eDqNBGSVb/xtGzuQkSnYgzlwk+Acj/C/
q8faUJwT3W6tgU1jEMhL3WcFGzxLB79+/oDi9O6MXzb9T8E+a8fA1obRTeMAroYNXQQF/9VFH+2A
iQ3GgInYsBJH0KrPPvH6wSahvHTFstEe2GORFYYY/zPTVnm4snBF4Pf3b12k9+bXDp0/0HQbcN9z
Supp5CkZjHtDNbM0lpSWBlZnNx4W2S3AgKqj5h6Ma1qsAYbLHvXunMfOpAjLaDuUR9n9omlU/Mf4
3FpaGBxljQmKog1u3D0/kfB4oZh8OgvvEQb+bMXhgIaYDxM/NKKocGM9jNQZhatUOcay0fE4IrAh
+1oTYmq0Nut3cqj4hVmA79O6t6EsP1e8ws2EHWN3blGYiWxIro4+xv9bEpY//tZmq/Fzg8d18HwO
pxTZOQkYWl2wpPoK5772jw9WbFU8rH/8GxeqUQBK4NUfgEl5Fm2tnAGwPzDXWvQt/TfK4sCoHDHW
VAdQ8By7zs12VKquWTmhYTW5etV4DQCBl0UD75W92oENlNXxo4RMoswW9Hwvo0AnXBFTzT6+NXio
TtqyKGOU/d7Zq0eOosTv4IwoThB2FmEnvJlgCW6E5rf8cJStlMqvKLk555TBNmuDUXs/mYabEDuJ
K1BrwgQL8MGe+TAYJ00JeCYJQC05z5FdlxO51sgQ+QmRp6ArcQLtP1Q9LVfU7zR5Jfpc9BrrPRLr
7hnSuggpRzQ3Cttay7giXGiC+It0mvD648d7ddQoB0N5WofODbkUOIq8Ps/MuctxPpN4G14ZuRWT
ylg2X7SO9N0oOTZglrM1jlA3fjCXjG09biF3CHg6MMnq8NIY3AnBVG9zRS+UYyznE1o9KMfCuHsx
QQ+N+fCcJluV3ee99T5QZgXxfeIfHdCueD4ulKw3DE2Nlzh8hdD10iPONKi7Acx45tS/owJ3p+jZ
BWZMgUkjTc+Duj0UUK8lPcTfP4zlLOEZ8Vr+aqVyrVBcgOAR3dfbntBKSTwjnVccPWfVyZIl7T9c
Z7uZ9MjJ9vP3EgGNgrL7mZysvBJbQGHe0Kb+OtkFbeuoVxjGfjyzFkbs+2f/ZJ/nl0enPRWhpjqU
4fAyQTNzaDUzDKoeUug5+IyId2+3c9Uye9sRo76pxQpcIUxZdQXZHiA/JrmMGLH61fRcX5ZOUOKy
lI7sB2TH+Ku2Mq2UueunQEOsHf/R48YpUFSWJvyJY4ud0h1/s2xAQ0Ea9dRyDRfq9beOrB4XEJz8
lPIjPL1EpOfRdcJW7wOfPiwUa+4DWetrS5uM4iyaqplhbT0D8c0rHWk4RUlar91QTs6lye2YIbeY
2z4KKJQud3YFsWkA2YQcpdrFX6Tc0uwnXKM11nbmGFRfiMdFEjgPu6F+1rDKtZ3yTums5wBVli/E
8hV3yYmzYZvhqWGA3N34xgp4XZI0RNHc90xAiugED7WKPRnOySPNq60cOV1/CTvfFPV+zSTbW5Jc
3GjzKm1vLJRSNDWsSGrxwgbxBglZAt/D5PLW2YE32553xtcfKOlj0cEFV67+ShIfliXlZoL9GIIA
2hMnbV8pzUnSQgzrvGb/PrWPvSrjMZBJsX54iQtdUwMTDh33NSmxX8OUIq1A4DQA6zSaE+0vW0T+
IBkO237wlj2BeBelFsyNmB6bvXGT8KeNFFmiecg3S3vmoWNRQPXHlukNno1/MeeM5YQ6Hb0TcpG7
/Key2+XyEF9ly+Uo2ihzWAdkaMdFqb2MWjgTnGTCzpbhkAyMggXOFLLP7+s/E2kL3MNodjSWYzfx
tBm6pTm1ErcILLo2Ae97+XX6xh+O2QdJE0x1hH5FPFk0CDA12QDh4+HSmRj9NGECF8LEy+0iSSxt
BUxUg1nR265Dl3jJJ+vBUxUgF0n8vq6eO9qJSDjmKEosMMq3Bgzj3OsFKnJ1JPXwq0hPVV7eHUe4
oBIqD0GBV4a7R8mpEr4rxzC2Ria6yQoWJiPP8LP9PvPEcTWLdL2LI9CyHsyPaE8p8KSz77ZqwCxF
Som78eRvKohO76fLwv2I3QGivuoS59wSxdbLdjCMQw93ZYT2TmS+uavxzwYTAYm3ITBPZ6VCZNYO
h6pA7b3QNH+d6SBidXG52Rt6UVccxDobpP7nuplUKMB8Fm5Ar/ipU47HL7lHNey8GZlt/xhh06MB
04REAB/62JZPAqWXWHy+WmJ9Iv7gpr5f2VR886S8y0267uCnLT00SuABqRvgZ1Cg3EC2UnWjqhIC
VpHZ0NFVrCM8NkIypsTISsv+P7M9wVTo7wixy2QwW2AmVbKzBEi0pfzuF0P+/0yS5+oPmUn561eo
pEvRcfkuCTVERMBVJv4pyuvHi+3+c4vpU6sh2l+FZylWkenxwRc5E8Q4dTq6yfYUSwigq5H5cKZx
bbaZ0Z61vuo9Bu5kVMMrnnJr4RlMqV/V7j/6LS1F4RQXodKrVNpC7uiaxvSgmTiGVOyOkd1hboml
OKD67ujOI63sy9OnOpJw7RVQSrFdvGogJ4JR9RGWKpQVkUReWwxvbr5jw+3vJxz20vgXuU/QXlCD
afwRevbiEOzoY1OC+Js2EGC2n3nEohxp5K4pb2RadjdVreJy5BYHYddd1WGdFfNMSOvJYrfWy2gH
Zew/aXZF3F4UMHz0WdnYSBHAb2NBAB7s5a/XyMpGuBcxmEXQl4gFf8r5CA0YdeJSXOuUgqYhsarR
gz0t5wVzLFvtkGC5CC0IdJ7P1jxEJIETsdB4BqDj9I3XwPrrObe926uWBl2yF7gArkx8Q7TIeQYN
NnZqHO6wB+AbicbQi94yo3dClST7KAXPQlIo5PTaGoHpKibMDMAtYd3rVHK+A2LCBNN8mOa/fQR5
F2REqyKZS9OAoFWHJYAC2NjkjNPs5W3dGOSB6vwbYU3wkeVMBn2/qk/cs/mHfyX1rPd0GoNTD+cy
N2bS77IKpNWuXilZGtCfnPiXpO5g0SB7SFEo0d+FFRmK0It1T3uPfSEagL7sGR/DtXvEmNPENQHH
8dBdyG5ZBc6Ee27w14QJW3tIaUgqfpT8nd1+fyPD+HsROUbAhcciN+8o6AkgjSkHFYvcfPdG7QAC
6nVfxX5Oo6t1woXGvR5s03YJnmVNNGfCVb0ULKM0XxWXXfEz45dAzcqpi91Ib2I0gxVLRpFZec3J
uXaf84oynQuXCSJFBlJD9WlT4hDLXpTqbOcC8knKevQ+TTiD6Jprr1gK1WkEyZVE/RkNIo6RrFOY
WRsFfj65uq1mEzxBPxF98NlepaiGVbdWRy2Ly7qz7tXB1ONWMrrSN1pPB/zRzL8AF7iF0TFheSAD
0AxlVoPnXO6gZbN0r8cAKO450Eg3QuozDyWjZO16IQc2wRBaw+ZkkAB6aaQjIrhXj7acKMeK+lHr
GBMD+OiKq/Qekus2cRlllFRzcXLx6DBpZplQNtp/rqAjj4ZhvU+GzH6/TrvRCLQmXR/tmtUv32p8
0XvZhvCG6lYmTcl7KLNmJOmbAY0hLq1rbT7uuRzSP3CI+cEIFtSCD588kg7Oh1jbgTHmSG0sxZBL
G3E6jUzf5ovx5esg4S14DKbgx8RcsqE5DluX6vO37FgaigQLzY9x5WKyB3mF1J9ybfogx2VfkL54
zayHPC//aIIIC2EuTUrcBKOd+xkiI/K5dhqF4R2rCW6oPoOoGt//Am6rq0SHnLmnTv3JrDobYRrK
WAu3CESiQ3fY838SCMreqajyVonXMWgRyGJXT5QAtKMUGQD0MS8jdtvEsnME0HKsrAANBms2m0dW
qfvpYOJejc2t1NWRv4AgO9cy0dMVNq3XpDzhwxQDzuVhna1IZFIjoSV+JjPldKCA6BMYdp9751Tj
6UW/+By511RXLn6eTVieuRaJMpaMrTpTHYyS3oisXy+uBVhtQB9dqxeBMnD1XXqlC32xn18Gt6t0
eW4njE9Vvs2sNrmTmVLd6s5XzPrR4yiEJ5MOh2wSxwg1uHtC0Cw4Y1rKsl7As+3A6jFvzSfn8Wwp
/lOpNCh147EnUqcYY8kVlBrAzUB4jeMn6dC4J6EaMtD1m9Tx4uZyJsckbR+0KJfsGSjeDf0gIDpJ
H2pNPeTR6JqFHKuB+zgLwm8Z2zlXw/dd/1PM5dfGBZp6P5YEthnSEanVosK6quiqa7b6sOvVy9fi
PN9CjD65hesePNBWLolHQWiBXhmweo1CWNzlPdbUxbRBIecQUvYzbTWPXoUE/Fx1WXZv5ciXf5FM
PlDP+gm3spIiX2ECyuHQipw8bYXsuywroXF9HDi4VGV8nqpQZGfSAARc25QWeyPPK4ohmPLOyB1Y
qbupcolZtDBIfCE1I0otLUuD28WxC1BqKmi79vhfqpvgw/+FculR0yKDT77BwQx45QJ3awx7pjWT
cumLix+ZdspFQ99ntY88Fg05OzWdTMEuJxGSGAEpEX/arsA3S049iravAKtXoHBBhK713Sw0dIYP
25cv0WtjI2kih67rtiwt59uHaKQiXUDLDvTuTB1Vl3qYphSI1bumLWbBkfHvoRRmcC4hoFfTrUEa
0zP+4JcTVgd+6EwkpGrbJVrMgxPa1JIhrVJk4Sj76GNQc9JJkR1aZ6svZkDW/p1boFrcwKQjWv8p
+0P1xTK7KWBgzj+PAMEKMYDQvDQP5of0lSbXIOo4nneaRawlsFXuGWgTuSD40h1TQ9DcL9y0BTKB
2vfNhQb0luBu9MEuLukRoVv1dgHFNW9v04+gbdFQue/QBOrbU69s7+v5+iz9Uk84tbQH2unLfFdp
vz/yJpI/mX8t4NKd+cRaqsvlDIObju+DdHQklHcxMMNXcmpYEP9asFqrMIndKqVBhKnF6yEu8B2w
eDGEUQ/Sej8Ho29YAxVsJwGi2c7q38iIWCMQ/c/WY11pnoK/keix+XsmRdQ+lvLSv/s2naZaPlPr
GLsM5b/hVejwshO9KUXroLRAEhbuUoe+VQMsEsho4DTnr7rxefNBgj8WCkUZbnr49mj4ZUu304FO
Oogw5faZDJBQHtArRLJF8zG95psXmlliAVAD1jFUf2yJ73BL3AiJeIn2FXw72vtYkCluM9L8CTdi
GFRXjWRYpFGqtXoXW/ipA7LqFgDQUK/+MQFLZ0qxeiHZrR0a3kMI5o/4vTQf+QLuuh8hNmtC09hu
eqSklMAnsRIuGvcAQ65513u6bSj3r8FbXSJJ+U0yIrqFmDFghi9fJgD7lXcC2N285VFaFRScChQ3
DQrCwWEFivmKRZBxB2q/Tno84q8l/cr0LqcKasY5tKStu6M3iTlhh1QcM5pux/DOQKIPm3WWTizZ
t+Sdmhbl2SFNK7xsudVYhF78ePglpAmioguagzy/Ooe1V4EBZKu1/yCuqjzge6KiCdsaP6gbgRla
ziaBUTeH7Q5Hg0qG6YiUmdR5vztX0nfa222zUzEUfsnn6llU1IoiXBjv6kW9vS+IGZljV1AHndvR
ytliLh1b4zyBh7TtlutlwgfRXDGvdYaIeAdnghh0yYbz559I5rpGDCC7jdDoQMmXnqyo8n+/NXl2
Mekn9wh7QYPwKXUGAWzzNsg4wv2Ry1G9V4uy1ZWuTi95trcO0z2WhvkiNRcalIcfN3NOxTPqNBks
soMouJ17TogB6P6Ahy2kFkUbUrlDuogqosoNrypaSP/pJYD8qe1xjeNjwYMbwEnBgAGm5eyRyJZ3
cnHFV7D67QLAFsuoiXwg6G6zf6VnuR9uUzSEee6LQRyVqFTVtJko/BIEBvuTMIlVdDldTh+TqQlE
3IGNhDqSL2cwj5aDBNIyP24gvUogJ4Y0IHVon9Haa/712xrhj2u4yq1L+aaHnxKjPYcD/jRx2DWX
3cRYTt0dqLryb9Rhoj+WWhtppH5/6Q5IAaHTqeaTkhsRjDzwmrPWQhkfcFP+oA5IT2aL3iZdvFWa
m5rKjaRMcfrEDu/aLYzaumNpFeLphxabxrZDqXw7ccj2iUoNVy3leaSCowINhdiOoaU1/Uk6r/yj
i5TVatvgPGcpH2DytlwnwlkUkkWPnna7a3+AyYNS0TuaRixpHKrcVhs/tUCn6hUkQfrwnuoeIw6Q
creCFb3UuB6BTW57hr2n4p8W7pDzy3ufzbf4fK3H+3xyko3bukxWl7dR+pV9vvCaD4rrpN+FgKo7
ij5LS54llxAVKA/3T9zcwEvc5Q/VqtVTP4Qc47eaoyjggM62oeDcw5rvJNWqy8RCs08uMdi+qGIt
OpxfE/MYtyFynxNm+tncp9ZZMuCA4CZhOzvX7wiPwd4955aU/14PyL0EkpR3BGW3qjacdqG8XwMO
OR8uTQ06VKEVTCenxWuOIhE4ZqVdVzTDQgD/pAr/03yb1eO0dvx6ZeJqgDdUrOg69P2Ll/XdnQmB
ar9ChnbY2Z1LqaXte3Y1uq9JyidRhTjIlSCwP0ReaJoK87jYr0iC/3RJmohUjbwDlI5yGAADGxF3
hobrCJCeyLDGo7l01SIyjl21rEMAISmzp9529zboDMbG+6+aMvzLtQircB1o+ZL7uZ8J2AIiQAwT
3i+dBi7cSKeRlIX4puHwwZqLJrzn/dLAmeeRgV6uSmjLElTlduz2CQjx/nwXqzf0Tv40OODJ0RUk
D3EFiKzQ7T3fohKgGZvDYnl0xVdsFoNZSNuJM9mSwonuKGHNxjAFHxMB7P0utE6D3yFpbhbKqnOP
uJU+WD6igvwqAHkPN+t1cM7aYxWEI6/Aay7L+7/2glKu4HUlPOvW+F7d0u6fUczXTLFwrQwUNtfj
yiT6c1Q4MSQRfLd0X/7sed8N7udTVI1ZtxlfZt0iryStHI5Dia/8L3zRKeZh9OytLqpcTEAZ95lH
Umgs8TmbUJ2Ztdlt1gZEDsp9RId0vKy+FjavATl9E5wA2CROOCiADuMebcTpKCRXpEE4TGYlPane
ZsjTkbTPrrP8rfx0t4Agm3g2PJt8wnDt8tuqke2KuUTdS+X1BeoGDqyK4hyLTNiic/RS1z4kXXtz
ZOh4rVdNmhmNasLVIcwX8pk9RDZk8gzBvgvGTsHgyDR/KbdRCi5qj4lGGpARv2dyXNnHC8jswZRR
xBT1TXTgVwTLpAXlCHfVPVleuW/mGqlviXkWCO/j6exzEMdK9fAZ/IiyAFYEz6oF77YhTnTsdrF8
ZFNxqzQjnWJUvUsgk7xUCo4lHKCDN/cSwl5L8WmDbAcQQCLlS4Qa2tZlusjw+MyXfjR9/iD/amtt
hk3+8PbkHHPHkOXPQb6ss8bKDv9noefBxgySnlzlpXUXQQtFC+ElOfXMFOuh7OOVE3pvgRF5h77K
rwBOipIhYDE1ysv0Fn7P8uDWUWHYO90V7btKCbeA+3sOixZ1j4xR7AhUUQmUv5BjfYDzOd1uyOPn
CYqubrbMXV07X7AI1QmOEvyDcR01DxvEpjUY2gefNiOwWcBpIcY4Scgo1Rp6No/i/HXBjoRljn6A
r7CIvsChbX9Yc2f2fm6ewYigiQ37nPOYkeFFxG9bTimwpiKx2hy87A8Mh+nxZZ5+KVbyqWw+icyO
/hp9c0VzXA5cx/gtDpP+0roorkldZyulLGvDZxPCOMZXyrQWOXAv/b9hkfX3agSEWfi7XS47jY6N
htBwP/IewMM65IMNUaWfRn5GOxudlc7EPInJYLImp9LhOOUPK1gUyGZUBWVvLxduRklknp4nMVAt
7UMcB3t3dmAvGpOhw1pHtgJJYJ2hbhFdbJr5ZoeahQRzbQmonepI8Pi6jthnW37Ux4Zqk+J7Rzmf
+HAfSWzBI/kw+GKH2MPmZtv1ub27cht2T5rQBXOSR3EGHooLbkQZZ0yk7kSHem5DC6eXhGsbOIRc
sjjGzsdLLXy1AG98yvCMi/UbzdzHeOh3AMwzwwLllOaGlyUiI4SFiEQJuNBPOF6uESefcLagD4zQ
EMM6QR/CPmut1sBDYrEe4C7puRh40jcjwCkhjeja2FBO5rH0/D3D1bWmlSj2y+9ABGVasGAdTaoZ
jxJgUEVnhFd9rDbyxSbV3IZtj4iO9aBKWvM3p9N7m5mgj9cWDbVJNEkjSf5PaqbfRfsKzjemQjcB
ukdEDAmF5MzHxpXtLVtjOllhu7VLib+D+Al0W5W9l+OtiE9Qmay6bAQgdrTwAf6D++fQsSCGttuU
bwo7OeU6Tgc8sYzFHiqu71nHGuZOj9CU8miVD/+t7w8I6LAWxgMicW6r7I/NuMu4kHw3WW0v6CBY
UtjMd9ZYYEOrTXc7kizHdU9Joii7ZQOQHN9/cOd5CPIOk8AJ1W72jglZB+ph+8LD6v9RIB3Tgaax
m8H8vaSaE+lmiOjRa2DAQmmrQC6Br+QJyDhbjaNflr9aRH+NFJZ3t8Cy0z2VZnHIks7AZk3s9lo4
hW+wuelk31b/lWDLQi8qp0V9YeJPfgKgAQAcv8kmB8XCo0gLPPr/mQZlLwOBiuY+4In4EzokqsUq
k9IXxtt4cUnn38Mgq769OzlbPG5Wc7x6yRoTiw0AuW+lpI7CCfN9gabxCy1Nhk+45AydI3g0yMrc
7+cgphogPJ0BZHXGiKDDNZQxOKOQE++PPKftk0DWWV9Q7UWhmtIDgJPoVpdzW7d7L9jqj601Z49F
YRE0Nsr9qjDXvzq3eKV5uq1inmtYHYNe+TsE1EcUCO08aCNoQzm1M4S92ytpPlaqy+FjH0BdU7d/
zFziWQ8kp3xdkVAJ2ctfTqk5r/FouY26tHCovG3VCy8qrpt9I9aatCkLnh61HCu6KxBtB3P9z+b8
7/0Ni9DXMMtQ2+x0nGJ34y8PKPiPT0hn95bVxY67uW+uTUG0x3cWFLwdT4afPhMOeeiHOTthWw2w
0GaRs1mTcEhMnwY26/PZ0ZWiK3KQA0v0qhEg4IwZGIhPMpK61wiCJchNv68DZX6yjRhLWmvqS+R2
UUyR3EKzXz5VBDQIH7QandIJA7IkMx/9omolmtYSS1zRH0czZnAelle+q+751aP58Xit05uMGDeg
iw8UywWJMMlaC0EMnDVJ8UrkeAx+dOUqpaUGmQsQB29r3EZklSwi4HQ5jYBOM2dGjVIC978ogAX7
rFTC8insTvf+YiYM7WdLj517xFSM7LGypMNaOSqRj3wA5SijPF7+lCbgHokV+kPckCiW8qMML0sY
Eo12EX/82FqN7eIMxLtocYyk98LiArO9xx4YcHwqN2IPoVAcbkMDhg/mMo2HwrOMPPXXKIk7tBNC
oV4vSbVW5g7PbADqjsyeuLBkMPlEXd7APbVLLZuvKLK/S9QUFAFEdTuSHlqjmLhyvYkxSQ8gUgr9
NutdBkompD95lO/sWg9puEk6SLTzSuMeAekaDP0GDReJMQHYCBuvZf7Yn7Rl3fU4lvhZM43Omrno
XMLYcR75LttK5Pam4k4KJVg7Do8Dw0YfTLeEVL4wtFz/OpHV/IwGaiS4HmBnQdzvw8gFFSfqbvk2
Wt1geWP0jFCKEII0pMwsaKFy8AV09+GN/FbjOKK4tUR+QXDDMeajmFv9rouKI7ooYaGeZlB9fmTP
qny/orSAuSpVRtDpy0Lby+CcdX3UEdulMYOCSJtGfkOUqz4z4LG4oLxcQedf6cRi7i98RwWt1QG0
FhqipD/qu48lIc2gtGgANrBf6zXbKxGzOieyGopb9jeQNrwklGKPD0L7WYEG9cs71VKdUbNFU3L3
tPjnqL/U7pflNKQEPNGMTlj8q2Z1j+Zt+m8Bkayq5J0L6YDEQj7S47NvQqGDHA/25nsaKfmN1ILp
BDHJzXtG9NzipKhvEW7WWCOdCE5x/ODVBEWzkOlOz4ias/SZlHa/D2VLT5DJ3hgPUdva23OpFYGa
1sxRFk+wMlqjA6LW6xUVuYudnHmKXTDAQJaWFefWGmXwnnT/WKoOUhSO2pMm7byBB0a0SYljEySi
Q6akBlylZ0V0HtL6YSBgiKYIgoT0137vZ26BWJJnZ/kabMQNENu515Xwba3+SB46L5y10LA15ILP
ugRPPMbg+7gIZAjxx/J/iWUPENM4BzFePrBW0br/4bqKXMVrBCjQJk3Wb/rLhdSO0Kox9r7+C1gv
1TSN7OpAc9qksYSbzhjGFnVRKtgjjdCP9NmfLS335PXyj/Hh7cmsem9he0XrOYs4FNOvYIG6M9wg
URQmgHl2H2k8C+yDGkPjpXYkqmniypuC2g1WEUCaxUjzCtYor5Lmm6WlV3Tqz37MU7KrrSUw0vuh
Z7UFuTDkNrKajRJEmTjCVUHJaro8MiFu9xZImrxR52WmZ7KmxUHiR11n6O/9dPGAO3nD5NW2Dh4j
JV7UK31BGOuySgOFB7lPGku5MjyoryHL/bfo6HKqlkQVWK5N3Ox+PohZEAvbeEmUrvy4q8xfhSpN
rUGXnwJnYobtkSvtz+yXW7BUTQv1y1Ey1t4TGka6EhLpxrhZHKo52sCnu+SK5TBKxdK9ltW9brdQ
YdMdkJZQHqq2keWCFREoEB24ch0lLEydMI3liskd2phRL87EbpW7h8Y05cSGvjtrTSc7Pm2s8hjm
AbvSqqCsgNmA1dyBOoPV8rjddfKlORXlMGx+WA8m6YyJHTZROf/ssvMpIo2joS5Sa1iXIXTvsshT
2gKPKP78ueEBGr587frbCR0YHPAkwPJKks9B6ph/be9EuWc8++QCVGMOHVROJ24L7mAJ7lQAI/pu
pSnVuSPVdEuaySS40n5oe148DWB2PNUuBPKvo8xbEAOqyA1sHhxAGIR8pUBNCcgIXV+67og/PB5Q
aRFhno6JXYHWjl9KJhlHxDGdwRuvBfOsjlGmpyU5YE3kBWjn4TxSEGIGD30q48L6oVaGiyq5ot+h
3mj28GDPNADOKJfShc1lvd9z0VqxSiSWmjjmuKoQRuKrLENAYKVHJ5Cf2QlRIb0CZb8+7kfqIw8e
605UGA5ZpsTRwFtW1rhW3cVzQm6d9Nd0MJdHL2INp9qWb9St5ivs6+aPSoM99kgo7z411QSsmKGG
iGU0aqw1c0sr5Cj0tG0bVQYwFLlVIhXMfbY7zaHdAYjXcQ814+7K5CScfPkTgDlDpvjBqpQOl32k
ZMMUJnZ+Bxgxnd7lRxNp3DUV/yJbCgPfK0U0h3lEmQ+PRueYCOOxOMP5zh901knIQtlSfXF2hHBC
BMFUSr9LtrMVNcBef8pb0WZ9wDRlEPpMM9GUJ3PjnB8BD7zoDtcS15SJRYySQjHs+CGCY6jAA/rA
ebYFNEXSPDXfMpBBt7rh5ZX7KO3ZMCfU/cIwcSLcVVeMdyXTkhVpAPxBBlU02Wej0Jnm0dI2BzCb
zf3CH//NuntCbo9t7ylvmNoyjZxV8riczFRA3ndUnKV3CFRvlehupvf1Yw4tcH49DAwNx+t9jIXm
zzhWbpKaMIcxhsKw5BeNOY257rrWJ0sAcT0pmNUttad5XZgqxx4zSZ5Kkro+uyL6q1klgXMdw+35
qiz9wCtooFhI09t6MyLOuC2dBc7aZHQI/cghWRUwoQplnKw5Co2Z4rJSsFh7Nz627hIkp8Wzm86S
pudTUPxGGL1u+IZYHs+WljA/BvaZiwN8jBBP3zoopikTZb10fOjL5CSI9QMaBofS+wJmkvStHPW1
fk26cftDU5MCfKtfWujN00Wjyoc4Yue+MPeFf5GWJrVdgdK0maF51pBfXc4IwjGJ2hlutDiZy+vJ
Hf4wvyDSMzBqIlCYLR4CGK/SVqNsy/H0b2AhOFL9aT/o/TpTP7AMYPxVnbhaWjo07aiElGLBc5h0
A7hTnziAaAgiPVaDkGVfjhN8DqNHZcx295DohfkC/W/sU20BJ1KC5hJVdSOg/BvEYOVtE7GDrT8d
iKrLfZ05bLWzI7X2VeoZt2iQpz41MUSs/E3dERZKKkKmMf2dDlcCQcONR1iJK0E+nkDCktrNpOJZ
d+y5zdAgTMfd7FW4KhoP8k2DU0lRPNZqLcAX1kneHD/TiFZE4uL/deOoSPHwjCFgi5y9+tTlSJVH
XAy3Fgk9mRfKGSJoaf08kz5S+iiymzNTnhG/ySqdJtJioLGIiZDUSnAbhq43/parvX5f2PjxU/LR
c3UZAcyW3pmojQDVLsLfHzxbdIpHOM80bPQDcQ7KbTUVKjLLPTLFfShvA3CnZx50M/mewYheJUC1
SWUZrrJx9YtIAZ7wZZz6Bh7avc2J5vupfEEit7qyW8Zx4iYPuo00axFmt5y/dIPmGor/bgVg0B0C
j/QTNgWrjUksofN4tjhzlk+fVyR6RnGe3LQgI2o0HeboAcD8gOMv7X3ro5sD8WAbGJ8dboKOZonK
3ZW/+Xdz+sTOeB6WX0bwbGR5VGRzVVUr4y9diBg+HXpf4BaL3Q2LTXPjrJ1H2x286wvlQe18e1sA
KExT9znqsrpKFyhbXipJAGFY/KxD7rFSThESdEfTyu0XsjJwrZJlC5Vel0I1fAFDXJJuUCK3wPlA
474GPY8Zf0I25tlA7DAdHZthrmNA5yTWeTbApasEms6lBaogCs6qHt2dXv8DJRq3wbsHkk8RkM+R
g8039VKo0HMY8L7/B+TpODzKX1kWm4Ko0vGQDW3TfB1X0DwnsfkSuExKupqxQFELuHN/LA0BjbnF
Lpfmr3BaQKEJs14awuF7M9QjgiRSMkv7xvi94CbD6fY4F6CPpPx1QcR5TC8+xm28wWLsM0Nvv6Rq
7tZmKvhvNmFEbLoU0urG3NWPbizaILmBosWC0j3440weNp4yvaTUnzn7pPhBuQPL53I7EXclbS9A
hyCCw0OevZ8uPAk4BPzkBm71JHBPqHo9xHl45/y0rVO8XsGajDXqA7RLD2uG2H1ziRVvxx52xSNA
9ZXFa1a7IlF7eRDZinMM8glAYrbNDZoKXHvOEIMYcxLf2qkvP9k2mRLe88LHdLgZiBB4plxRJ0we
rWIkU5qKU7zIqZNlmNYmpo94bBUgVSL3Osivg/2bzCj2aSVj8EfUYxhhYrfwjEjyEEDDSTDHWzh7
8XRbAmv80uELQrw83jPSrwU4u95kbVU9WtqFb/ykN4lp+IIDx3AKiCIcpvqkuHL9btGI48AIyQRm
8LtRvF/Mk+BpXA934nOn2xGCeg95rHe/jKu5l3ud0QmUGtBRFXzZLAywbDjD/aEkQ3P7bLTyCAFd
W2do3CmCsIycXK6zMaW0vM1dpF4f2my3A/LIE4pmwmgRewX6TR6xhw5rtQxg340hOq5vZJ3ZnAGD
w1/utF8h/iDrfOwlY+zgSMSDcwmp3k1lleTq/hV30p7F7aQiyYCE9HVJIz+LGJ/UeJK7m28tBUIO
Ypt8Vnsw4o7/tW5GdtjrV3FBKqM0rqaB+rsMrPzR7EYuzrBepB2yYGoaMl+5YDkVLbKse07/dNKc
Insm2l0ewprkcrV6S/48GSvjoeIjruC0MTZ/QKtVcrY1Fo6I4jWlV3Wyl3n55Tb2vXb0VGBcCAxX
W+sdUfi3ozbbdaR3+/LFDvGI0jECDoJ2Lovd0Pd66ur+D3oivbZs9vnPB/za0puV90nGOD+VAof/
88l81AI+P27tQ9aaiaWEjXB+dzF19JIfzm7Xu7ag9rRzr8WRPQiQLmRP1zPowUbVtwOsZSx5GvW9
to9kXV3xXa/f6pr78WXU2Bha8Hntwk4Sn7zJIc4uATsrNuPO4frSEIxSnun9pe2J8YdTW0kY0FI8
Ba/g3xDmu8BJB2U6kf/KWSsPDgkrNcPrxAKnRy3MHVJDVp3ZuyNDb16NYjAxGCndqV02y2MDAizF
ScRjy5iJjZAemTfoi1LCufgV9QCG701aZS54zvAjEWPIKqd1iX2b2H4VLTRJK8Q1IeUXfkdCCDfa
LYjY2YvG0Pnf6K/h4paf71xfdJHjtjufUOl+lF/NFT4BoKZcpu8gkIQEjVG0V7QRvWtnunlKa5b4
clbtBnis4lgyXAsmkTcHBiyamUX01Uu3bILfOhYhWdToxb3FNzgydbjbHalUz+14IF02aK7l000b
NQeipogOMMYgn3tYzrfeTT+tFSgq20cmTS3wrU6jHOzg96ytpDY6hFtt++8+WjF9sUUnR3HhQcEz
yfV97CY9UaTdp1z92NYMsHTNshLoiasidzYbJkY6UBaJQ7Jdv38jl1K93Eou6p8b91xXH08gryvB
+0WV5IAYlH88UWSfC5AKz6PSC7ZaC1uyUBsMG++aw/qzND3unGz9laSv3RA/K/sB+lUNPcL8voOW
RnJGixaq/3bJ4qYxaPvSdPQQe/+HrCgw8uCQKk9tHQg9EbTISjpgbuqtm6k3RDJvJ2xpBo4xQLMa
iJdpMb3cSWtX8/+2SIqrNuM/ySubVsao4rf3qUMSL7DAI9FpBJTjlaeqGbiby9Qxkgdg0ndGZGOs
s/VZrg3wqBP/cBEdN602yFnM2D6HHI6H7q+lDGOXm/pCGpAOyhPn1eEdQ/ES5G+iBpal1no63q3w
Yj3rtEehG80S3ZtIdeS4YWlvoTuHBZlLPZBvNPlSyT44u5glecT1PA3s674nOkBbAgn2MgMReXBi
1AP28+hWxLZm4P/WTYaEuJr4uEprKb1jM/Mm3RJmOaqJ4UiEZjdwOtZMMMIXBWe1952BGn83sNRL
sPZZ6BngFq4XiZFzf7XO5k47iAfUedsuMkzHfTQhCGqgIqQmdW/FlLV+dqd9l4Zf/SoSIt4OlGjU
e7/HSfkuuOBCaPpsgouBGT+L2mH5bcmbWrZOneAVvprQ4U7kK3Q3xmA2hTm2IHnM6zD/gueot3Zj
leNj3vcFc2QGUC78Ao5QPTj7fYcfKC8jGKqzTArJtHgUL5/0gXwJMRMxmuoekvN5X5OV1KgKxgMx
G3pWqN9+N3u5Av10BEvIGnZo+erCf00Wx/vnq/NKoZ5wwGsCzqBA0vkTTdK6di/n/egEl7kbH6fX
5ENN38cvJVQ/m7U/pepCObhKTyU12SfxOqFO/aHHQsXHFMu+v6pc6l+X6cQ22+bHpUiC7FQVHROE
yY4wHzBCow/d/8INqDACBG//5kK4h+J3lPTImAqZqAcrgcPoc+8uNrDnIh/W12dkPw7gGmCOfa7u
s9fpqAakaa6P0hC7QJLlUyG7NytlqyiN9IkWGMcWQng4csz8QZnwxKxFG6+FKbqEPQ9TWwFJb9Dm
c5lRRf7x8C913zoAdIBu/ew+oD+DV8+lS24rfnLZ//i7SXL5dHtR6QfIs5AkBhkA5898AQ1q84jM
yFgOYt1fenDUCclJ6TnxEZjJsHD4ueHpUsGh63WKaeXXLy9nA/Ak023s9zuZjeFjbNHhXGL654CD
hMAaNUAOidZ2IQ5o74iExP1AzTWvAIKf7Hz/rftx8P9bE/z/+piK8FYsC7ES/SflF9n/59Iz8+Jh
fm9AivCwld7iFy1mtf/RFzfo0lO1h2w7ZLv4TjBhYt+A4YzicPQeokGgmWbEG/ENDcBsLHKbWdnX
M0jm6ORpV90uojt3nFhuVmJn/tW2htIYflp1NcCLqSO74ZdXUAyMKZEr2jaaG0XgaxH94BBEvR29
K7aAcTc94wGy9yOtdTEjvFL5ptxVdvlvbeP0G0LLtaFpU3qnkHHmxM9s9OjgmvkgF/lXIcOXBNFF
TyQu0zzfRs9r2ZRJDpW2tF21rBcaAPs3lRWFOBSGrBy7zZU093ubTL+wXG4MIaeFZGgdbGPejnvZ
p6VXMDRvunroxev6ZwPhYr/4w/ZPfTtvvIEokzrO8EQO3H2ekVL7meYWcpSYuIKT5d/j1nRwPvU8
37kpZKF9fhZotF/7m/i9cbqNRNk/7hBLBh36Hw31OnJ+CsuRVWkkDkl+DiAQPWsIX/GWughR6MkX
j0/ATuWzGam+dgkZbHxO7fziW47w1mrvodC/06nIMvDFAgQLTzem1rO7vcuXF6izlrkrCcLk2lvP
GNZ5cMpUds9Yq9hNQj3DykHbnDaNfDVOcU4u3efo/QlpO5ft0XqMpuvJGflUg/MvxBF4bb1uuy/q
Rtw4eLHKwSOAEEGzOaOf7bZhxEgeTPWmj9YNGdcF1OCtNyhMX0VKwfx8z3eQc65D0UmrKJw2CrbI
CFNtVY8Fn9mcGP06FedgVUwBso+/O03kCm3NhKcUVg9VU1cTw9mmNwdWwr17pYGDNoqGkowkFnSw
IBymCwX2U7TXvBfdOnse5y3yrF0G7jA+G1ZOfBnNq7cg1Edw0HyHFq+cBBkewZCQ8obTCtLJoJ9O
XCfKwQYUQfJ521PyowW2qYQn+J7JMcdGOYlG8MZaHbSC95WBVeo7iR+JPvw9Ug4ZWxz7fu+azLeR
9ItZNk5CHYAqOJvYFIqo6Q9JxXqEJWNQJ3JXwZojSdbi3AkRPxO1gcD6XMbWwR1Oe4tao6V3vCLW
2S4UiLojKFCaQ6h+guqvf7GZUuNKKmUQpUMTMPR23OghK7bjzXHYEXdkkcj/a+l9vGArJmEFHWBd
xHcrl7EzJBM/wRTFkpMrZUSz7ygioOx7bHcD8ocsQ65EW/md3aZBpWsDDpWTsg781ikDG7wNWOrd
F7SPdACmN2dHRg5nuvTZxvs4Hmx31GSRmcWQHhbafK1A+ESOLm66GGfGCVtH9n33+HjYlefev8Dn
gRSUZihArINj18VX/hiGQyQHtLWVba+JURz+vbDBF0BW11qUJvPuI1/1x8kjrAoMN40aRPouQtpB
/uCWR6MoHbCeFAVvNdAR6huCFI3KNyoyoBMmgrYk19VXLhlyzEYKXkqa4cD6p0+knozTYoJbH38d
rrDlSQ6v0/V2TQ2RxKXJYxbHcd/uIcDkMFjFBuWupP8wY6rA5zqe7TE4rpOdXbQbDqVNyApB2h11
bfXlKpY5R1CEqM+ZDYVatu1qO9p/oMtJ0KVOtE0xHT1PSOa+zpSusNkwo/Lixlgw2jgrTWa21vP7
ZKRDvkk4SlKDoHa5jwsYDa5X4B21nOkVT/j/XdEIBEIv/0IhvfNdk9rfiS/XsJWBgRB8nVeZFUkE
Xt+ORnqpURenVad384k8Bb0cuxJh6zQprpmf8YpgcTl5HrLqX+w82dsYO6HgrnWCWvzHmsfhLtnB
PdijRcuv3zDFFkfOqff3VFDSWod+SlfLRWUht6aE0Qwp9oOAjiyHcAEoqnQiDgnbald2HmkPIERQ
geutMJGhRk/9tNuVfQ6DXpuZm5fYfpUvC6ZGF7no7Z8Y5YJw7zFG7owZrR+sK9jeKxUsePYbwHv9
5qVkSI1edBg0jNym1Q/PXJQZfexOBTnkIvsAQxIFdKov4R8z3RdPL4sFyaVNHIPXSfrxfJeQ6s/h
5TnqygCyIP/wsT/UCRD4Qjx4zBuy2t9FMfVAhwKSc9MmkpKR73gHGeXq1znxGHGYXFf2/robq5iA
WPL8Nw3EFWHPFhf32j73rNg+/Gegi6Ik/Y+Bsvh1VEOuA5RXStRItBEZjpTMccOStqhVcmaLhCy5
BK/JaVYexYPZSjrtWPQLmV+k/cTmbRY+0af4NACS4s/Ht8aCQ1zx42JuGklMbBbaHr6kExgv9oNe
i7cfq/oOxdPBZNnRg8zOfBB0Cyo72dj9mO9uo10RmQ/3d1lxGobydDFFK1GvEKXW+yi3UiZijRKm
IY/KPabMNt78P+2moxxZZLPyo8Z1uDMOSTQbtvrv6LjLS3VVxMAsAcT95OoFCCH+jx3+c7Vohli7
2PWH8ptxMnjvOYtndsgXTTAJRXkMEmfNjO6saxbSrG1HtIfMsLdTU5X1QQ0UryIo6CC6fBwMCdMV
QRwJlBndy2kv2f+pX/XICGztC228+cUweoNMieZMbr+f5HdconzVduKuIvR5myt/V8a5uYXJAYG7
IAxZYsnlVV0syIVEDJm9xzWGGncQZYoKrjEqR6OC4zEdCfEvwHUDmQgcQbCilJgiYNc1DlAIgMxZ
BbD0fthZV2lVMJ9Q2CnG8ipz9WdkxSbrxmcNZHGr6aycimqntzAtyvvnA3xE8H+0NUThZS9rwN/x
a6qeDweYmK9s/MoBwb+e2EZsGoPz6oaDfDHyoal/NACdSo/5mgKj+OsMP9eShiZhaQHSf7zD8bqp
1717lFs4ySHcIsqaUBXd3M8zqFVHunkUCm7ogwb1RX3MdL73vHOQ36YN8+/RWU7k68s9lxqj4yzu
yhBLi/PxU+j1lpIpKvMwNrZfVawcuRJhS+PSomB33D7f4jtfu1MHQj6wwpZIpQCFsaQYUGnQdy4k
4Bhys/TFoSwckrHlxUvECgINPY23t4Y4oLgpLGvr5DTxwUJHuA0uQcr2R6tI3rp359vrnE/FNhSA
oA6+VVhJs0QYAQw1Z2+XYKvtEnar2WeApPJ2vizoC01vq81DsJjcJbCZnCRgjRu6BySZo3rJPHnb
91BcQXlakocWB05CuFZEdpyHULPaP94b6qZxM79qN6V0Tixt2pJqHxLf246heRhEaOzr+F0onDpF
+JeG3uLpS8Jh4X1i6Fiix+VPzfGGp9EMhXmpdH1LLJ68B4/wVlakYdONkmjzq5YOMdy0pv3Hat+q
OMFd8+0fJBhHkkSQb/8QGjezti46f39HciwAPH4DiB9D1LQvV4wmCoPMx5xTPnLEaKxwSwLoWFvR
Ppebg2lmlIAX9ZaOCU5lFafri70QgA1SGBFYOHUWcOMhEJjDpKBYaewwtZrXO6QThWsZodMRXeEW
/hiqBRGlKFVhckRqDZ9/M6rHQ+unMsPj4lBTX/WvZPQG4uxH4wlhH1ZfRnrFzYA50FAyR+VS6OpM
wpbMIhnqRUxzUoABbZKe8f/xYBj2Levv+1m5opgn4SuJfT+GRmGB/x0gyHGdUfukf9OOoXWNb4iM
gQq690CoQwpSA2BAwHkALA02pnosW4chBY60AN93z+2KO7S3lFjTjAW3jWBhxznQQK1lltxT6vHQ
/n+1Cgiw5yvJomCAs9zflZaYKZzd4MYnmOCiP5C5RRK/WAstfTCxulrOhl745GMrpxSeakhNo3WG
hMEG6BCJ9rZiPKrRZ3VXmLiFh9wu+ntIqviqmwgUe/XTkrq2MSoOOOsYVQqoNIhSKgHFD+bZb/yV
A8GyatdANK/N9/5+m2zQjW2IsCcHk914m07NGUrCINuOeIeHX4EM69eGzHdu2niIePs7nZzhe8dJ
KizWhXR5GJLsZ7g9w/Nth8tAlHZERCLu/2YXBd0FSoYYcOBPwj116ZmmbH+tisX+ZSPyde2PESPH
28jR8o+HdpYJNKwRKO0lmB0Ub7mh9E3QdRGA6m6TdKIAtOajqfqgXyA7PBmJ9pUcDY9z3pfKMIKx
Fqh0FsggnuMP2s2c/I9cVtRjm/fbPtefxmDqiQZIFjJS62jkWtVKfKPRxtw2sITCe6Z+dJrSSZD/
XnmzSYiS4l7VVfBF58E9YMhOLfTg9yjizgk/wZdQRCFfwMCIGcgQ7kvPWUysg9/57rfaoSWFt6Az
Lb8csZ3u6gcdcXxVRRTznUGRNtyjSOmdOYvUqUmJh8jPTjKBKlwa2gnFHDVxtuCISHiF4S0mbrSL
opJ8I8QSfmFyiEYzqPpMF4OU3Dd8r9r8JhSJEr2kPGPpUj+JumSvoLE44It9J7SvbkCnC2ypYNRg
omuPBNSo9J2ADSyn3vsBTJpKMUjqHIfsO+CKi9L2CK9Ttq0R9Wv6Kn4e3Nn131JEtPG/G57kTpsE
ojmY2zOXBDJriDN0qIKR042uLNoUAmTlHaWAVkgQhi3dRsg4WNhzhZuyNnMJ619cYkgribgO79Xe
gkedfUCUjHz+lf/ytKh5fu3VIx67jBMSHyDkp8pLpXLfdqnp1WKYETBDQqf6LmPOZeQZmgS9D8Bf
XL3txSQChc5jqj+Dube7TJd8RP236lPAuQJCZMftZ6yEIZeCBbk2hbNSdUeU9/3Ti0+HdUUCKX+/
a1fxyMA4c5JJ2yt9yYYpLjXhmWV3ReI3cPLE9IhkfwWlPjhsA8IhA482iKhKjvXXWWVcxyn/YAly
/Q1KBLXfLSD/GTES0lEqPquPKOBK5i4sds5xmMW6qIIMOckRL1ES/6ERtA7V7Q1h3UqBw6DpA6CN
tIQs1xN69kI8TWeUk5lON9Hjq6aUTPq2nU79PES3nlI4upDcQYo4akjNI6VIdW/DDggqtREEmNI/
akLdwbi0IQBV8rRIUyaioKvVJ1R+YpwnOyoipwYRGtLJWwD5qvVs3xotEUvEIDBN6B/M6ZWaQqxd
iMhTg1Jw3/Tx94AiCCGmkVyR19FD/1HHZXf5AEBDxP1c7iFBQO1rlQx3pr0gv13/pJuBCblKvQW7
ehlJ3fI1+Ok2dizoLvipXMR8pCzpRinm6L+DtUB3AX6z0+10qxNlFM+8iTOmlE0RJppiJxci3RRl
sP+atUJOWVyCdqzadp4TNF3HrRbWHCfz25EcmvovCfdCcBvBxsHu1J44B8PvPTwlmDwDlqp89oN9
c7WYkhazxkUp0glAjemGTmkTAUcWzkbVJfctvL8iSMxeQ1j+L020q1ozsGIegtjx8P9ZpR6HMByN
hvS/MH6LDRP2QmG0Te5a7hCDE65PCdjvk5JypHaIhv8wLtNFNCTsjOKbKgJtYlxp6zfwlIrLXrx0
/TE1BuqLnNamtTMeOMDvDHjPifiPZqTqtsUo2qJqgACeFYH6XtvTPr1du0NHTHdqYVj1dQvHFoay
YreejlDsUp5AWogIl/OEu1e7sY2VI55eykPIjG6tWeDwMAy7i+XLkqAYg5Iazga4xi6Xixo01ksD
zqynftD+BLkjpGkrVNwH5b6dGFpQEICpYq7ONyyWtMyecvfS7dlOgCznpyktLn6m9NjXo03Zujqm
5Sl8fewkK2PHX+37YaGKsSViTDeLooUp9PaKUzTnUCqZWK8iHvtIS0ru0GG77MGOMvnfkP7afsla
YmQwNC5SzZjzESk/bpU3jBYG0kMvPOIdQf3dFjoqJH7h9FO+8HPAf9VXZ0uxP/EA3vB4eiZDqBCk
LVSM0bTgcwYgCiMs1DmcLxfZHaM9fWZ5sazhBy+FMfEQAlhwnplWKvi+mFBHVciSNtftBq36ORl/
bSKXdPjQ4QZTZN8wr4RfDGg4XsqYa2akdFygPlROTtspGjH8KNbGwiZRIJK/Dwj5rwtcxjQ7gb3r
NzAv3KO49NqR0diJuCxxPqzNNyVAAXFvHSTk3XejvYfXYtkGekJxs37PgDkA19YVJu5GaAG9FObf
+TZAjgNOztVsf2IkDeOWBT8+M2f7X+thJVVWR45OKTAk6I+ZTzQUqBd7G/46ydBedzM4MyzHBGi4
YWj/Usb3yPgnbmT4BowsgVApHtVE7WT5EmH3BkNxf09C2VVeZdfUfX84OFv3yPA6lAggWaK9msUk
DAR2Q+gcE2pdgDB2SNnEDqGaRMjYpvPq1hl8KeXBcIp6WOm5neD++UKwE8bxG9opZ3i9J8NtIOee
ZPVkaWnlTow2ywCn9o115OR1vW9SWAMpBqX4R4/l8KY5Fsh1g5lU4zHfrBidcM5GzcUJiFApm+PD
jIQXmXCaBeSS3jlTRpt15f7TYQayqdsHoT1aTutKT3jpkPq9BFxM1tIuheryFgBsmQX/GPxRf6k3
/fJmbyJn0UU2y1WA01s3gGB3swM2LCJItaEiIlg/8Pdc4dWB4XGNoenj3dD/9tz6dn6JRfyZrlzY
Gm3XLCC9VMl7AqOvCoJpJA84u2ZtNfbwbJyQo90KqUNyQ5FLevhk1dEywpLCjpTbx3gxRuZMcvsa
oyhxKJf37pCT7c2tdzvlDgJkQDG6uTaG89XZuYAopSdfJTmLJUZxhTpImjIzVy+t3q7HaQgNF95H
UhCp6bsC7u65Kt0VCTIIXVi2X0P+fGfvanODN+GU2N6lIwNjlMcF6OeDZ8vAGJv6RhmU1ZqA4H/G
25CM0mBv8UlUxyPbZynJ/TEBKOD29jKwXpMUIrwX1EbjO6HEuYf7PPIfZOSYsfc9d2KfO1i1uM5S
dImzvdMLlZWyJoKDCcp1tuQyvAJKOUoFkMd4I+LiCc5p1fENHCA4nor09S59hVd8X3Q+JWzyOUTS
LLCwduBe/WW9xMpqZ9auL9t7ZbA6GLhrRZk3ICiiSCCtTAPHC4TmT+fgMxooyy8FMeFwwLK6qRy9
spRRhrnCPq0hIZwdbizr0mN24Sf4RYoAvLhM23KvahY9qPu5IVNQmtI7z9CbfV5bJQ/iZ3Ocm2DZ
uFvhtbwNwGDV1E36zkE1UFjYkZLjDZWqCTAMFH7VDFQFEcGFsKijoe73/0qpYzf6k9ZetCN8DrQA
AHr9MuE60YNEq+2eNCfPWtaGt0LfHO+ueElcwv5J4tULY0F5F40C+X0sVGoEWqeu3LE6HY16p5Mn
XGpZLnyLSiDdM/rZ40nuH+C7KKqD1EcYP+HWM4ZInmLlnMQV+PgxWghKkMVIei9W6hsuvCzbwbGe
HktrwYuyZBhMV4tg6OjV3/AjutrF36P72/R+IFJVarV/Y9n+HON/XnV2Cg5F9ylvnq9Us2u5+lrx
iEewurUoN+VXjIGhWka/JBKD+Vsd2ZwDWG/KA0bAAvqB6UPrtRM9oIBCYV/KwmZA/QyBBQjVDScC
DWL49BleoGSY24QUmXlXJcb0CScS8JKPSYVsdbEDbObEkmm25iCFTchhZ9z40I4lNybkWArUBdv5
T/WAMx66p3EzX5Xp4p82YfwxWNY9lpKjtA0ABJ3NdNCvoqSgR/EMFzJJRLXc+4Y3kEox9n+OGZ4h
vyvIERZpJ/vZiuTbqnDSK92pO2tGoUXpkZ52OB36VqzJCOjNuo0vhPRNiraUYatVO/b+ts+Dp8rs
YDSGfA+Ch2D1VhbQ0K4I1R/qnjoLOKd+XuILy60Od7It/zqLhHS09f00xBUFzFlPYcloobGdxEKX
fiREIiA6VoePODT2JQzY0MzzvbMXPZfzTjv7YvjFZU+5kwpBRaIkGT9hoB9zSZ2dvtCojTNKJB3w
7a1iSd2rE/0Lfo+URZ38VMhuBv6yam/djZasgoU2CTdodr6SDeDlCgyy9eoxMGGisQv4SzciZmGo
xv9Phq6M0UqTaF7F2pCtBra0esu/mHx7NEObsDDRDoVW6z8ZuunXTE9Iq5z0Y+ZPnrp8qehgtKO5
n/D0SRZp44Db82vzKj1NDZcr1RPZVwbhNpQrQo/HmNE5YudUO47sjmEzoRj69rVkBgUbrF1x+wHz
l1h8Gj77NyB6lsjvSX2bnroG5KFZIM3NWj3JenzWarDBfAquCriq7rxKVCdZ52KPOBRQZAlTjsP9
CiC+/MO31Yu0CHEKPYrrXsMDvekUODlDxHo/m0vdRHVe1uJ9gdahZ8DrxRxi2TIsz352U8V5h+JA
zdzEbN1cgbGnQSTs4Xr7D3+dFjLxv+RaW5RnCGzSSoJOMEHAA6oNhDYHGdgA69krCRQ7txnfOOkO
qA/Nj2vw1lsF0SZbbopUpQBTnpj4D6ghhjlCP5MHf0Gv4E1U7z0QlN+P2r8y0oqYoqrgWDJfl/HK
9zeS2foPNkDeC10NFz5x/PKBh1SpAIlGt+3YEf2mUOu6D/cPc8vie9o6bRxG/DpeaNYsRoWKdFvy
5fxtA0RJ7/9wAro/diEPA6GU0AEAWwVJlM5XRGI6jy/gNU8HN6xPQWB4r9BvNOLt25DhYtUp+2Hp
V/q9bmAD8NQLVs7L6+dTIc8NZ2fZjaNeiSyN/a307AsIO7jmJ3xrc2NRvLJjq48RVFV/+/iRBRmF
XATQKqzw+Eo/8G8IoeWgAunIhsXVWqg97cA3LkkHvOoKYSfo7TygPFfFAtyCMw4T74DK2GCWt2mr
KODe/g4b3GO7JxrApmKLQE6C/0p0ORyQIsp2bJUZiAyVwtNj1kp98WYlWoNvGKjBxcArn1hhWc1d
DYBVXz427PeJVNJCJYYfcEs+F5TE9KdsCwUo7C9VW58XSUSC0jod3GLsz2pKBhJxfxdMVn4Ljkpx
cVYm+RPvHJ3WAyh1Z0RaMEZQByt9GmCZjhAS7vBuCbXm3fGTUBzxuKnZbufz4YyZ4DF3q1cEfsLF
Sr+4qlLjRdNvVQz3rD02g1p/GD+rvHie418wxCCNmi5uZyns1HN8RwrGmJVx2vdvPD51/iR0zLoP
tFKJoy6KM/fbV/7rqOXyfiA1rDNK4jIDHE+KJwF/4hI2Cl6ZcJNvafvFW8OjafJcQYycDmVlCLJM
mKBQzB/Smf10tu3g++1QxbDySFh+AH3rDv4HOx6lUYAfvRleqCmzcCBxw1go4luboYPDRfbTeh6s
8rKLmY/ooN/Tmz4MwZxCpjVy6GpCbU5iD5oNzjZXGHLTMzSOc/0jMbIn8ltNtfx24uaaNUZVB8V6
NLBahyvZRVi+I70nsc6f4XxtRY3Pq+YiVeyd5vGsmVQt98R6ZP5VTmdDr7BwZilqVyp4PhQ9Edey
Hg7PVZaylRPLe2JITkCoRdXrCEyxQvTlvniv+M3naeTsgUUYgeTmG+ah2XN2LZjZlA4XXCLUX8Pd
fwUYjRuz3Any01FalZfGf3/IS5mU/Nkm5VHSUAu0rrHtwRSve5E55Y/M60Ar/kBJ8cvj/6NScZMA
wfnHzhKlhIhy5uS3QfUt+8zMsabHFoD7EejyOrZ8Y+P8H/0EZKJDTvdMvumCH1Fi8e97xGa1+7M6
XSjBHB0vSN3zAWz9QtCApR/zYbwYOz7ITTSJ7t/Y6597+pV/CoVOu5v4nNTKaV8aeV5Y/+1HHDzY
yC9Vi3VXeP9QwRmHlxC08kkGyhN10mG8FSslFe2YNTvmJFEVXehZR0VhJCgblf4Jc+x3ebEomn52
fQjYrczRGh5irxoUgsptglJt8UmwMJPIPKWVoz3DUPk/rJyvcmAE20IHb7NCvS24wnJ/FaVqipLt
d1e8gCvPY0IOKn2pmTkxBWhJH3g4ad1R4Xa6fCSM2rJMGiRa44D5kI7c94wmkvBzt5bRTNS8MuSj
Sz0lVlG3BkQxoXICoyb2jdoNYyJ+kNNovILqbxrh37eJ4GT6bZGQPLW83QOcrAPZ2zD7WFXLjVSB
bpm33MgfiZOQEFqmyM7HXtjTS2mn/CHsWPDDhEh4h/rK9zX4NrzUR1flj6KkbBFljP4CLCc7eRaG
5GZpANLGhPFMq1kUZDtREebR9kkYL7TXhwrKmHMPyqSnJZYTzKFZKQ9lFvoPSWMn4l38W45G0kCQ
0NZGqkh6qvIfkslOUWU3DUBy8ZOGmpSTYxy+nTcoFpuodr+nT6pnHEn/LgL/T2NpOaNR7NIrl9lr
wlRPrr+uDtQvTDe/8ghgxXhSSwqGXmUfmEGGfKD8WsyAg3tX63Ci7V/lIeC4AzqXi8PW/tafPu7u
yXXic/hyP5dpwPQZG00Jr6xKddBkADpPi9mea6Eb82tDl8fCUoIBugaSf81kwR9EzaiwmQJRoC9S
7yvSV9b2dAH81pysp7z5/DDpURfMCAuG/KUXF5RR2PMIOpEqDvTNROyt7iGsC2xCXxi8wvu0ncWC
UwKJFcs6joO9VNYfsGU1ZF8OcbbBt+wNXWVsdWmdMETnhI/buFEIyASos8c7KDM5uxvRGxnf1Lqh
fth0AYqYlmEyrH7zGFjPwCsrUNl5PJZ9whpLvhoyXLDjbntAERRDgVC++dKweMVzFj1SIGNfoxwE
GToVlV7UIAWv01YCvWQtb5c6ckQhJRe2+ZGRB6OB+B9PUjH91scUxMbmYeAo4HKtHkK31JW6GXWk
NhvFC6NVulKQaaRJAtQTgNoXbxz39QcOku/LANJ7uJldGe/5kKayT/zaRqhUvj8JV/pSi5Tfk+yb
XMtEGijT4vALdBnQIQ2jgQwp3PijsHRrD+JsDVmAcUnVrx+h46eDvztl3+A5jOdi7bI8cB6jEVjU
+bIVHK/h5kaNNqeNxPzv5ieW4YlG+KcbKGU496kgb6vuhF7Fuh0CRs8m9luKtT3qycXIr/fLDQcm
guy159LWMBQm3Yt5ccUxR6b3MsO7g/vywzvSmLdoYB4SEWQuHquHQ3wCmbUmxJxbaXCJSdH8NROo
3BY9MiPYenWI3afP5HFCL3+lK/YPtSL3+DvyPEOsCcksymVdZNjx6mNGbYW3ic4DCEYf5Z8dGG3G
fjjHiWwF+HPxPezxLOLPgDA5wZgSoseHMHWwg3xNYubZgcMhz7e0FE5+7KfYbC4LidHhjk51bRPK
vzA8veql8ESm/ZqMntvlTyIGhnYN+yUji7wvoNO4x5E04GBzvehFoK1/y3ms45ij1F7hix8nKK8T
vbKAlboGY5Xoep3VGpkC71xMFv43jGuw7j2VGGngRkRk2aaMjmPOQLZMrouA5R4atqbk44iNZwVQ
DwwhZAR7ULVnmU4RZLrKnN6G5lTVv0svRllsh7diXdELNtNCDYuNwmC2gPTydjWTIuDv253W7Qsr
/v+5zR1ynT1fxXnb0iob9hamZwyiNmAEahysT8H7vzy+GX5n4foUBNqAheRQjsWzAQUQOGxAxSAK
0LQewwUGm69VPZaYgF7sL9JvSEndS3yPVwJ7ruREuY80k4NtUk4GmaMXb5WH1tb+CrpKIN+BPse2
Jj1E3keWLjMOHkrWDMgRFpsy8GFEgTSRRwTP1l4haUyjYSpDm9HTkTo0vvZaUl5ESuigQm9WwkDV
HzGj+UA6MQfgAkDUe6JfyqeI2Lhk3vv2XIj+k7P0vTWFZFbuvUeooxgdAvpk8CxEbphBqBnT/9NM
LBZTrqa1Yw4RMENFjzm8hyqZKW1jR0HuV4Zn9oh1bxcLsfCpyQXHscPKDPI0RA9Yt48heFeI9J20
Xwv8mNgd3D2DLzR/SWxS7KMZTNL/LsVqFQK5Qu73HfMr+kMYKcM6nzZBYBy/KzTjwJ6n8Aa9xk7f
RrCapAKKcQ9pJfn9p93e5GvU4jqmu5sIhqXo/MWqQM7x4wHr+9so00VWY8gPnvRo8KaPv6+XArlX
7kl0Av5Jn4pTMp1mAKHW3qfi0CSm4JH+0lj3BJY3HfuEZMLGSODhIZJmnPnSDD/BYh8Sj7bzNHtQ
RrVlfZECv8HOliZPLfAugCuyw1VVtQ0ju55eNy1OgNhCyH6ALCUUGlGFUdN++RIIz+FD5QFEq4FC
pTjpHabUa+FYq1maw1W0Zf6CMGZFVDC0pb6zSFlk+WzYqu6DSwaF38khOrnEEaJgcgecqaQSd5zr
/KtXxHTMxZAZvSy02WSdDPems4rO3M0IHgWo8JUQmCcUHM0B2EPWioNS+NgadTo3cdWcHY4AeCaa
tS38cD/Z9B3IWxm+kLJbULNqs/gElXDBrwM6Q2GqPfNQMUPEbinqXcdyYNuVebdFgKILh3ll4Ss7
f/K5DNk3k8OMdzFbUXjiUcFMfVhWSef9iHAyXGhSoJ4glxBmHh7E6Y04PSivzm6KLDWne8TgJlVk
HDHbiY/phL2uB2clMb0FHbWouSqz7ooTaL+E7w9aH05oAkHhZz5dRcfV23EMin5yr3Cbzis0xCpg
HqgmGxd78TC6AZF0CbyPz3u7xyWlpWxLxWyGrTWFmixdeFf0BOd9IP5TbWM3X8YU5I83z/u2UtOT
VobyMLL0q2XEHbCrRpzmjWqtcmYuwPamEvhWmOdLBFsFsrfJhVup0Bc5essKGBGddZh8OEzlaKhG
PmYPXpm+P4r1v25t6L64ngET1+1E+GO3LDHL5BpHtGSfTp/bjVr5fpY6nu//Q0HJuGqKC3ywuBAi
nl71sJoIx6OBbslX/D9HzaC0Th8aEoPaWur8rj+0EMt3Wk37/8VbGL8WlNz+XLKQdPqz9kffBwSd
lleFlgzxeNXX7MOyG9Y3Wud/E0O0/+Ju4LTqadOF5GV6JtZ27hhNc0OYWZBSpqR6djdfEhnIVmLY
Hes4U9Lt0evfM8npZVFa7Y9ciDleZEw5XNbrLYk9FCpDqA9AHK2mNAE8MQucEX4tdwVNe91KSItw
QWccU6ZEYl7l/+tO7t/GWEbfxtd2gMCh1p6iu0dw2nQ8a1pk4oqyBr8BzrMN8aXu3/hs2qoPlU9k
Ij69tPZDcItNjsFXKU0PNdhUIbvFww4RQS+JXBpv71jaUbtTZQpaK0hDWjFtPInyGSSMtCyHf36a
nm0sOKMmUtBeYJXz77/0+AuEhc6IOvYj+hFL19GVFChY+/h1JZ8MB207tw0gjYVcFXuLwSAvYMUg
qQh+PA+PPtlvS19i4lPeqk0ViUGL7fLGmNKpjFqV8GQJowfJXboTzeiPopJaaCnN2KtxmmVNA6hE
RBGOlM9/vA9dhVF+P4IlUeGgszSEx76HRh46DgXwtdP28ytvuKVH+xgJi4EaFPnieMot8sIxpsce
BaIgeFPggUYD9Oope+U1jzCNfMtmOBpkg6g6wXRPq3iahQCGGm0wTon4Lb3r4Mu1gmOm5y1WHOho
5J/XpB7UwQuropCg3dciCWg/PvoQAEmPt4uLBznvUcWrswWBNEChD6xNbg5HLrtfUg9hHac5NKnW
gzcCjkafzGpQvT/R+a9FyfLDHS+2j2eTOWOPzmSw+PAz8kRgldSAmXSwYyu9mwER8gsd1xeM737d
/v4ltyexKwHxMt+9J0ZLc3ydxfKkfit18LaQTrp+PswAEEjPdrC7Q7zVhuEyYJneyYt9fLUHI+8R
ePVQc0U3LYBtOgcNz2P1/5eMTJh/HOzFodwuCPdRybH25vHNRHwJ4XUR17JB2RNpAz1gBNTgOCgI
NO7cqfWYurDV8nhYItIewYyKBJhU6SwfYHyuIn+JfEH/Io+gFeDLb5Dr/s8BNi8GNOG6h7jRadID
Q3fsoPUIhqHN2u/juUvzZ4PFyRn3kl31ZmgpkH1whfzaRYAe5WBaNpgSnXt39qlicYUX5BwbUiSR
FF9LVj07BUuYKTRgD0DmZOmbghVbpSns4l7QvQtM5Wznxj3Qi3ufUyfuhCz+V2R6t/X54NaNU13a
L50s1m2x1jg68hcPybbFquYHIRMuYCN725rEQ1mL9X/+HM7F1aEE1Z/uU1oFkvd2w8OgrPATWNH7
kJstgEHF1VifoaWRhsz2Kyfjtiw321+vrtrCHNMGxaH1o40BaKQ7wW8axsA10M7wdq/OpcNNqM18
hmtqam0jOTkiM+CObUQUqGH85ecPUWIICLCi5dO6yELklhLWBTAFZcdiPh7ERqT/Y7sJu+fbcKV3
hOamV6wd1oxWgLZF3NhWVwrslNlRTlWFZMMoHqCoj1N82wMXdm0kWTr0aXd/Buga8y6U6z6Z30lc
z8wx81bloPi387SgjefWW7IYgay1+xWdPSABK4AAdHpTWYugt/VbBX1fVH8hahLFPr0+Iv7fhCSw
8duUvLM4co3p9Ei5JTF8Iv2juu4iGqBc5zb0O8iTiBXk8vgOVqW6aMsaKlLxRRPLlMK2zH3nL6Uo
jKpHBl04GIJBwSlEqqEDe51svdm7eayyBy5tyrzo6aVRKWmshEhpb4oesH8NGbiMVpytgYAYx1ft
0efTB6oqJ4q/ypLvO7jjvfmZTFNtGzCFlDmDmADVQ3ue6MM0lsuJIvqRENZ/BHmybAEAL1+Ub9KG
VCDf4H3AqL4JHK7sruWX2OWGeJMsHdKsIbLwLkIqIF03susPkIBTAdli89jZjFMZVpyXf9o3PV4f
GUzBb23ZFCal0qipOK0RhlPxwQr9zELvDrkAQ8IkabM67QJa3DjT9OqRsVSw5TDWirNrp0jsXXAf
TcA6HuAJnmR09Qh/wB+ghuVOUUk0P6j57bREgk0BMxITGl0mLlG5ee1O5Ia8/HFtcpW7TW5x4Sjj
C3XVcRH5sfagIoeUFEgOxk6+nEngSKLIeqsGOzwngxhyhzj2xm4HQrb2DWQ7OcuXpN2r4mUeV6Di
+fROpFFZKnitiibWQqc9G5nLJCAhL4+4jpNWeDh+WSaQVx1znpf8a38KTyUp2LoHWysiK5YJ0Oul
gkFm7Q4DygehX+XIj/dqUNxs7AKpXn24rbgYjruZ9abreeTjDrM1EnK8YsPYHh8To7l2EJv1zjGa
10Z0Rcjaz8494jRMnMUuZudPaXdNXe6fShru/F+PjLsY1tl+ZJqWAwt7KHxeHtLI6qlyZRKuH7sK
hoWL8yVP90sGoyOV4sn5M+V+ji9LCr8ALCQ379/LhFMZYd7cDMAIiUYvbx29fc6j1neZYL90GYC4
f7Rtz3cdzuSn48ip6nWbDDrx62g8yduuT/id8S8iXWwJra/ZTwWjoYE7O8qBHKzGwpltJwm3cRaU
+AoG+Qk0/gmXfZ5GYz9a67uOBIQ47lq+b7YqLjXud3SV3UbUF0C4KjHsilg4x8Yh7JKrN2K9OvnC
o1VIzRTLgjckPs4BBgv2f4rUA5Bp/dgjeAOoC7f23vRuhdfH6AzjBOjb48F2bKYl4LjxWEP3dSGE
8znwvGtQfjWYi6VZwPcVzmuOol4vOqssxtI+HoEe+d8nOvBlS2knkKW5WSnM8vXHJW7M7Ta7CkqS
Dn6t/of9Z91lHDVrBs3ZdSA0M7v5jJHdiZ1nhVucDQHZM8mb/jA50BzZ2WYqZH7gXZBJA9Cq4PlV
lqhWvM6OxXToKYO6g3anBujLxw6IsS5ZiJC5AzO2PWgSgdK6YGYoj6+BQsPP+UG1F2qfGN9aTZgu
F1HScsDcZ6G34u3pWpIGiBJLK8NOUslK9vSqPhvCNWMl5XXjSj3qEC5b/0/q/1OzJFwf+6BGBgJf
F8a2FV+PhIAr00kqvlcoSmmfVFT9u5ryyKyxUSY/Gi2QFMYk5iPgIGNA30TLnpJtKijMwxQ742gC
JaCUtKJBJAhEccvosnskS9iF2CdCjsHV9ujBg/VB46iWa+kQdapKhlomUIaWJzBHmapy33wZEqMh
o5WO438ehi/yx3oXc9QZD2ehGysAT4uldXiFO0tRRH+mp+tf6zNAFZXwfssAMVmtlhK4y424iMiq
p04rYCF4HOPGO7SDv7Y8IK1tO19uFCKqB3e95Ozolah+fpiR67USbQvuSIDOVnddHCf94ICuikKn
dyioDagNoYNC4P5RJJNsIrzhITwUk3OZlGrU1ypzrGby2/y2vSQ3/vO9EuljmUXM15/mdFHiy2HW
0SDzZ90HlS8sp/m+MsOw5+ZFDfCHKM94/reCdetxz7qhP2HUUSDthjNbep7WKMRV5Qql0/f8Kv0e
m5QWbANFc5s+4CCjtu4DAzfETfNMxOPTa4wTJ1eGqHaOKDAROL9Fzk3dm1NasdIxPgtWHrYTOLPa
hrHl0aE6XnlUoNH7PfIXPO6zK48aJEJuRTrJtJfuqOnpznMrmoXk1mPrk2PX+8BaqAE8V4bO9BLO
URtkjwwpPJ82LWV83hUpFZYSGFI60cB/alhgnnQ/bg7xtWlgb8TNUENw1HrKHE3wtP/e6mYvuJS3
T8MqH06VoO5kGfaMA2b6K5TKcyJAP9MoTfzliGJDBV5rW5jV1ukY47KELJ99/y1vchdNqxaxhrjG
I9iZSYG7MXS6j0NvDjAZxVtbl4C1YoF5U1Mdd7S5n+wKhogBLQlKXHdbSg4EAwijtFJPLqIOnfnF
ZM11vBrwuqa2NGaDNhYzYQgsLT3KdU+2JkcIYiCbnkb2uqbphJjaC8wNznTASkZkw2Naz+rKAVhr
HiAp4AAiJmrVdo/j2YyG+UTd8/yyS+0KJwbKWwMkLhkfzyUZdHnTV9O4MTkB96lFD1+7DoY68DLN
RO44Uh/RG1zlUrBsmJb/jFbVfKu7ZNOXSJtc+dLRe9TR8b7s+3wgYezhUfV9whqpGaIEnp31zAih
jAd11lKdmeJXxQ5NUqu0mnaE77zORlW6Y5+2GjI9nyi0cmad8ZWyFuJ6MC32lLG0yyf/YsC8CVyQ
D3jLES4zr8Fp0/8X3EtBWsWHYakQ/2lwQ4jSOUMGbjhq9HzUZ1jEf68RrxPXBdc1pS1rltQ5U33w
tKucs9J+4lCMIWfoWOUF2vTdQqxZWFvgO4rkq5o+NP7rC3HA686gr8+icdYUYiSjF/nSELqzTgMf
gxX9jsgUFk88uHqR/K4RtDnIzebsrymuFG6M60zuwwMZtSsEp+tXqBQ1zCK10WrBCgQM7JgxtS/U
4R/CVleVR0aCJnF9MgRWHheICsWJGjTEV/2QuDOjlkL4+vOSpkxWV6IWEZmQA2MUA4sFku0vTaW8
YuQClhruB+OovE94mFWjrkzSrBEpCByWJbmDhiRcjD1/8Ex0FON/xukY21oy7DAt7uYM+lW0p7pb
3gmY2jSNZLGODodPNedWBF9hVHkpQglrj5Zwgkq1qZp/pkO4pfQAWsUWm39XsvDtfKSFOLJZGczA
7P9naAjpx4U6nTQcnxkcUfFFRj6WpsWkTc89lu+BK0VlMVyRLXuhuG5BvNFP8eYIwPHecOCxph6L
gMTMRKazvHXOuRkw5rGmgtvPZR+oPt3ieCgBnmYtwiVvcsscgWVLjJUaaQ3o+uF6YE79pIVXSGaD
Q1Y7/mnh+7aHl+TgZ6ucdtMrcscwqhuKeQqY3vFo1wz2R8xr07ajlvG97BbttnI5GvQC45iBQ3E/
DOvzdK7v0MNJBu5F0VIyCRdLL0Xan1FHLEasdNfZU2903inbY05W5yd7U19aTMfDnRjNWpm8vnsk
Q6Zlm3FUaTHelbzU31AXcJOQEFli9wuxyUUkQ8/HQaOZSi5MSrN2IOQr9l9SHC3faVBGTD2B80vm
DNk70E8WKrnSQ43ueBPyEEQ+0l2/BpOWASN3+9POfhsOzPRQfcVAO1TwbG7Ge60bJoQosIR944BL
iXpolWtl4GbVRZw1rsxR+cSrTcLxoaNIqfaElqOYLMDN9ercna2ux10362Qgs/sZ5grNo3HQehye
o3u0Q9VCzkJ8t7M/QbhyGXMAfqFQfLRA7hLx/FDUAvsIlNVztHcd2EWqeKdGBwlKyJt0DT1HH1xy
4ffC9HYTV0f/zx7Nkq114fKf3Gne16nstXPVyN43I05e3niJv1sJBPBMrUTLvv/A5m1dKX37n0xk
HRgvBuYIW9XCanm3B1F/vldCx5hXc21+Oe87O/12IttfSkINKMS25DInnlSzfuxBXs/d/5uSPRSS
yLFqNMP21potl1sV8erEIODqVeQtNullypH3vxN78SS10zqvvgpnUNqt7usNMvAssbv6KHOkChMe
//SC1v0vaE9d0Ayrt1Br0yPSzDvmRRIKrecGMJbjYhn0PndGhhKtSRUfqEznuA4rQIytvWs2/HH2
7VUuoJe8yyBEO82Dpyk+TkR8g73rjL7rYpvOHOCdXNXEIeC6iYG7WkNRPBB2t4th9iNFeJRYLbLj
14WQf9im0/2OYP/CA7NJ28unabcHoXuFtAohZnXroCoMdafHIhu32GsqGF8WCewtddwlvzIdEKxk
V1trGWSdlvsTIcw0yG7ZIUJsfFehHgv09ZC/BvaFFihzIsM5eSC/b//87AW0dicS/FfZy+uBPgjC
HQxrrfWugMviEUGC+A3fOT06jo4A08E/7ec9gBgwFkaWH4Y5xHWBxELmBw4O1+NjAxnu9UJk+Xxg
gShHTuVngXZhOJH94Zzo4bqCmtuhiHyD+strHmMLgagx3r4jzdiRHv0WBrHnAW21wi00Y+EOWWME
MqR1TBJCjQwZpfKi9aFqWbPjCznm8qLawb5wnMgd8jDXLXdsLhusO3qhMmLmiMxQ+NDvxaTeE7cM
CAIE/MwIFRPkubF58uY9pLKCCceSbC+nk1kXuHxvZUVuYu8ciubC/v8OKiZRA0mPHz9ZmPXnE+w8
zNWmQfFu2kFsFhiViZ99GKu6aIpJRhGaKklSN3XJ+3gUCZiIAmf0j0a6ZKnm79wJZegG2ubCv1un
iRDCg9ToSq7lwvYDAnYhr8xwrNy1ptRoW6KmkQu8sua1a7AFKMSHuz+n6kWaJtqWdPWbk+YTS4v3
Y15G0M0MQVnMnAQN9e63YAvH5fHU+Zktb/dIN9TRZ63r9CmBB+fGfqjKF882OxvZjT2mzFnZZgUC
aptyVEzYxYMIeNr72iVvR52UMSbW+m8N0O33gBtIr43igN1BuEevKVgoPs13SzhmwIa14n9iy/Vx
SvlgB3T3i1G67tunzcfOw0acvTyUrmeHORadSDxtezivUIT1TtD+LTf0LNqfCMMQYmBazlDbJUbU
xwy83df1gNxAHYx2f+xgMhpSS2RTHQRzO172yMsITNkRbdPe8h95GESIRW5A+om65hg4KZegVRS4
YpBOHwTlnzxkSa+ADPqI06tykTS2DA68N9t3oEDtjFdaxEdD/QfCpyOGVe9rChFc0PidJcFgjlvY
uY85g5XpSp4DuFJtSnAxX936A+hzvCJdngB9gNEmtO2RdzgNs0T03IOVJdk9vO7QvZJ0V3kupJlZ
U37fo6Wm3IKfXre2Q9wcOUnBVKiYoliBIPvG+yimHKmFOjk+NauKmFv3B8dPzlwvN/9iVxHtGLv3
SQ/zEVvRlAyHCcKzCoDx7zlGzf3qt35gmdfTCbRIlL17Yf3dxC5LiSlIlXmER2qBmCtuNGBz6fCn
bvz33mipc/zpFRBc8e6JJxT0T3kYFB+IOCWeqk0EJa2U6tPNvBW05t5ARhu2yHzjZGqoqirjdsnl
NOz6L/imvkGDF5pcePd7OGVd6mMepZ1ztjKOJHujpDbOiCYx54ALCm1txOhnPtsAr8RNkUrV3mgV
DJe29XU/C2TpfT+jHsCXr8lbk6okZ/zJG8dWpigl6FIvgzFCLWGAstbruDBZgZqJVmirVRTwBC1s
LlbMK6+WiMYhUYCgpTedNIUHwTx7QHk9GWx1BxeMVquQsAiQ9d8sIV3vUIqxH31IhpTDAT2vSIR5
1RrllG/EYlomv98Usw/EiCUR7sXuzK71TIXz1GsdgUV8P7H9RrgR4OmOHKfndxhVfdVJ8uN9LI1L
EIhCE+jxsWLFQF1ASBXPzf6CcWLazcwj4KnnUsOkTWCEbi4en9gIxQO4V39es1jFFNSZ01wW8Nn2
Kfg2/RQtHpLjY86W0MNQraLi6DU8EuDpk49vGbWI1v3AYPLtDrcbK6f6+Ttcupic8hCKad0wnV4I
t2xsQ0RArZrhpOZn2t+r9LXgPPSVlRll4Sas2rFoYd20UbR6NB7wX8o5phAasRNa/BqdFdV6pTIt
ezDrmnXk1ba+7gXfw2hlNMnvLwHZnDp7TgmYy8J6MTSQPR2fVVAjmu6Z6t9YNcein1LxGeKIIvEr
QZkzeZOKBxd3YLNeF6St2j8y5PN2z572pE0B3K+sN6vkp4TqEtKsmzKCkgPYcwyZY5I6PSx4BRnq
lVeWn9TiyLEfWlWHeQF0mHkSeS/kb6+2Q44LyrlcWWQFqK3w/MwH5AXfwJYiQsQozeWZw0QSWX9d
vrVAtmLhS/uBiaCrsFUTKfaEGd9f59mDubTUYNogkZPpqm8C9ax7WerPuEDoEtqokC4T9d7gHB3k
lxRX3aWHi+6jQYaZRbjnJNa2r0aaXSiH4Vt23c8eR0Zu6gT/cIG+k7/79/1DudY3I/gsbnc48bxQ
SSHgh0UFpJ8i7dfEGelpLErOzchNmFcumSxFDa0vyjcu6IyQkUzyGKGS02XmDcxwXGMnX2h8hDQM
ZhA/0X1Fumi2zELLxOnq3RpB1IsmabWOAbW/Wca7JCBq2g89iT3KSpgGy8VsYc8m1egbyjYt7Brw
9ItQWC63xfLTUctezX/145fT6lcqMBWJmk3XtwRztR8hukIMtNDfG2HM9794G4vADnEknq5phe4p
xOppMa4C4ynJp26e+FbN/O8uvuHSTgOxmYklpJbzoPpPcnOvxQo8/ByQAClGg06zwbSltrhdD7BV
qjwwFIYHytt+Q6G4o30KQ5dnzKhbxFwOaTWfOnSXT4Tt4eYb1HI7OV6Cwz/EaEy4JlwVr1iCj2Lp
Bnd3uAlrRnCDkfw+szPn+Wt2crnnEwKsMmdvBY5r9c9lvDJWL5T6iGJwkFGy7KsYZH0IIrTE1tvF
RuJaibSSaBzPmA3pZHoiSC/WkqAmuCq65BnADXGU3pCYV2mNZ9HKjxHdmVsihuURHC5JI3CEesVy
3avX+QFA64aUbi5Il+m6o/pLn0pJxOmv05dDxddwA55qgA1XrnUsNnhHf6fjE+eMaUQb+5HuiApJ
wKvnSi4PLtJFngo4yEN+480UUu817oY3J1+td27WVrBa0WrVkegY1gVI975bkbfJuJEXNYA3FS/Z
u9F2jO63T+Xb+Mf0JwUgKd2DL+Ug/qYZMuYKIYLZNTJF9y+ZqZEhxFAgZiL4Ck80ettdhWECAUHQ
0GFq+vZwVUQW4pIHcd/iqKJUbZJuhYs6Yduqm6Bwe+DIhHOrcrQWwiRwJGpUp8Zm8+gTivgpFh3A
V5b6L9TQj7GK1nJechdulBcYsrYHz67o+SI/nShAUobXO/pP2xziFwH7WuGpY0TFDtJHQq0SvcEW
GPC+YeZbSZDaQKhzNHghFNqpnDEwEFvaoKhBjOPO6WYLbVJu9FSP/tkx1bSArRl6b+2C9CmYGOQz
YcwVGVYEZyO/+K6coDDuHdqVhM6FCJr9cZOzg+0OK6FAA796wbR/nGXm0xbyyCCheBpMjKOLudwg
/C4Vt9s/m+3eRXTVlIuFJQosES7uuWg3p2BlzxADU4j28BvVcWvzYyhN7AOP5knLg+e1vq3FTMk5
XPKZBqtluOxBuXbXETTLvFSZpZDKEHfPUV9jlktKD2l/iqA1yrJxCb1wE1mkpdyjE05y8yqkakSB
nWRDoaE8R7yUHj6MJdhpa6lXPAqhbL5pCjURTgTh574jKl4EWp1PYEwueCCQcusF8g1kFSgBmU1y
m9Cq/BBFGzHkJZ25aU9BAonVPREN5fG2rWNTZqwljf1iS23DSxuR7ef06/OOnCxzMV7K0jJEJWcV
wwx3t6vyv0IsaVJc6H9pUsVOgzxJW/mvCBKHcyG7J8cbEg6xL/YroRjwlpoWT5BdyIiLOMgrsuRd
KXGDdPALq4lUtega/Fs3IP19aVe4V+YU6eCapG8ERd3CX5YU2Pa/oFz1i1PExxh8l2KVlL32jVbf
ibP9MhPeZdPMBwQS14I2TkIYZiMflvRwadeP9rSEgG2tHHD8BRfs/HkQpVIBdgS1Kg4vRZs2Qoxa
gz8bR74Ho8ChaR+qTssJjRiSeUleQmmQMcZYAscZJ3srO6K5G5yVt+0yV5F8p4Vqc/fE7rOBubHk
oAQe1CzVjaHjbDsNZJIKsaaNCBppmidKs+Dmdehoa/QsNcVlRlkh4oNrxObS9aVF+jE2LX2P1D46
NY7kJWdJdu75b07rmPnO+Wi3ZhySuF0fZmgBWWOwyBUUzw8Hbm8T4dp8SFEmLzt13aVaTVY3CKwE
wVhg2IqUzNmqiKwnmHb/pjncigHKHE4cuGAcaoktoZ0ISI5IJ9KlVbmt63ksoTT2kxcQ1vty7wAd
KnCh/jLWejTtRBdPDonNJ62/U3xRAszJP58Uk+PeeKNnHXSErTyNDBg2TREoO3ZAd9tkZSBwS2hU
ZSe92D2g6f+qka4b7uH8NsbyOocYEquZZZzkgXTryedlfKNF65heapvvHgn2VFWGDPW2RHusivWD
TA42kYzP4MFfvhTrzYh3YQdX2UCJiGs7VcuGSVVGMJ/QzbvvEM3hkgaoAUAVuKaddjXYp7eaGTOQ
akBWnbgaLvQ618VeYqyQXcGknU0fxUi5/pDD6RUI1gm/S7eektWxOpmmsLkePbe4nM8SYIvODIKu
043E9h5JoYeGyNSbNO1vgoBNB8P1fTr1/ntOQKd7qCAnUfzwjAikPUh9zPf+IxtfRJVqoaqda3O7
PiAyl2dotIarAv8/mNxuTq1mpHmTJuBaQ3vrrHwOUmKxY9cnSKPxotM7qGus5XTe7kFEqg20AIG8
VnwtCGKzaIU/7vy4MeGnZ1DLmU5lH6D+I5qp71eGks0g5ls0rB+LBtXefagahDc/1BzxlHPcBJm9
GjRmGi9uJVeR6oKn56j+/81vm+xM2IdHYduYWFiwSPM7Xb5ndzSpT8jrJrlPxWFTFdy0CRU9rp3O
lkoai/MGMOzTswsp+TDFBNUYUf2t1q6AuDcq0wGwnbgvAETTEp6PjUeqIjPxhFHm4IDfrCSZcbFk
75t4kN6Xydo82QKKQ4VpfDQ/PtR395/hDy/c0o+PvY7rCZTM2hleokZIGx0NkJNUkCs9sufJZGkQ
WqDeRLR/StgaSxR4u6XJ6EJKno+mVUI81g912CmL66xRnJhsUUbDbGFhEJaZDEfbQ5ZcaYgHymmk
ALSgEeMYb4hsD5USOgInqVJk27ILvMEeoSgbx3UseqzInBguWXPc7ADKaBYOGL5Kzddjo0t4ia6q
K6nW/zqQ5uEdbN3/GVmsMKHaOS/QN5qhBI5XUfr1zMY79ABVDZ1gdYPME1DchTjD5gK0etZ+qbiX
Hr4z2eHUmQCmDVYfAqzOL7Aa7gNiTYPMPhMepnjU1WgmPYh2F0AUUebZVkZ+FeaB8LMfRZ/Jo9Qt
NIY59FtFgLqD29/CQyZCo5EUyh9qyOlAdxkyhfy0L+jop8hy7TeLxqmBRHSDDzOJW/7Ti4BZgsex
TpMS75m8n4kueNh4VBOdpCxJOu9abRO2ykIYlOpG0YN7vu0ax82+qbkjm1aI7YdkMMuFlOboAQ01
86JX8Gyfp/6WVfzXx90jjNsfxpgb+kCKflm3QGvTWKkExgL1+PnrSxaL0k34vUpCLizlgEbuVUAZ
5Imfk+LBJHTe74TAxDITjvThPKA44QUo0O0BdMaOAkxQzlgaH/yDVeToOg5mihVBG3fj7FK409ix
CtaxpTF4fw/NL+cj8/cDA+Vlfm85PlClqWueyo2+4KOhTG60nD/oEPmww50ibFbFmdWfVzIDKojl
1H1nK+cWmVT/ey+F9gY4oT41jQvEsYDuO741+KRnRbi5BIGLnSXTbvqK2IsZgEdPgjem5TRa5QNS
z/dvJUyohFn+d7Oy0tJEbJuIQj8Kv5Wm2ZoP9+9ZUoBfqHU3SeQ0gwqbBQBzT3IxlmYUswXziPxq
GFNmTUsXqFayAbe/ChCV6VvhU3xFmh07giO5AJ8C4jf94M02lQqvkxfYD3DUDNaz/NMwqRVqhf72
tzeOKHZyls4O2WXCrcIJvsU0gS5tARyQZ1pcqNfGeaEL9o2rNt7ujIP3TYDLRgdnsL6PkFWzOZH+
GPsDco8kCv9O7CZro1mo74/aqQbr22TO4w5QsFSkjxyfyyeYqo4vIrzgCE6lgLHAEDflV9BCN8gI
Sk10/fepd2pM1fsUxSLoTHIVF9wcPZN5F0y0/kVfgUY/RK0Jr83yHAcVcxHfMDhMQhE3LaprlZbZ
U9wQA1DcUOjc1xUpkim7haUb3aRlZOPcPCzntmmk2Pg7onaBXpy9i2zvwrWzmbVAVOqWezaBiCAf
6Lf+CUg4SKPEhYzx+dkSlcXxllkrqrtN9400aWR4YiC5I7aGu2cWX+kyPMkDuOKcC1Cd2o1x5TNk
3TochNTR+Z0p/AZD8OSzejMTD5oyFQnuLpOaihChrFzlews8pMLL/oGnSgemHP2lGo/zixCkWCt7
WtmY14dFHls9FuBhHeAW39nMpTXGaM3uGpyh5c8BHuL4TI8ysOzKwHbQfEycrFwGRcuzAQWDss+k
7RCnxJ03r4P3sG944Og5oXpjpRdjOgiPMequl2hM/zPFqLZGMEWAy8mJghjuhDYQkKA1aNfUP/Fd
irapd5Rw5za9Pp79ou5qawM1ueXveEpzR1Ttb6bBN4cg7sNOsRyaPN6eyjg09dI5mvD7PO4pUS+Q
2SqDLYSNOx3SyyfT0nI/TOAvZzro1XTQXvPa9DVhdPHauFhjx+iZo8SQZ7JeG9BH7f+t3ncgXi1b
kw7l3+JSe8VJiRJ3AsgVMb8VixkyUbWlSuMvOmIlSxk1XVJx2ZxeY4bNjosnWNAyN67zGQR16Tgj
HIR9Xjk/af1ErD/YHXolavQM99AYb8/Ba9zMq83x1KjJ7WKaTuO9itEwIPGZcyKXVwIDzV2LxGJA
sVLZo8Do80DxDP0q0Fcz07Mno/8bYL1+RcAQlEJzXNucjYYCX42YgY+wBIbaurCLOekbztZsQePf
B4zi6GavFqFfDEOODtTOswltz72hAbCVYjGPTf66muXUpVl10iGxXs83xcQBHXgsXu/1Pl7dOEUn
cO22jMObxn5Eou1K/xCtgr0nqyCOZSLl1TgPgD14dGiBEfDjGbYNO3W2XHeXhhHjoMYpjMpdKwVr
BF8KW1DzvsiAQ5ylF28vNtEvv1kx0pEk4iFkIA0XSisEkcTNj+3Nq/nYN07biiai+qd1H+RK1ux3
KgoCeWI1SHgW0tpCVRky/SuNhUXV7I89wwnoCrd7+opCdsIyi0lplS8MzZ0JktO39oEMw4+mSuoS
kA4dRVX9MI1vExWNP0cuONMWf1IreW6VH72hHjtPsqCEIwTYeN9A0Ncq5LI/tkKwGaZubrqcJGJZ
4SIG28/E8TsPyJ3F22xXw0Nz9KwxD/atDVGTBTsCq6Qt4d/WaL4e4dsZuDGeLzJA4pHDeYGilxv4
GsLPldfVaem8YkSTLT1mnnulSNLcPc1m8F8MDB8L9abpHnKbncbQxcpLqE65kpxuh3ZUTTg1ylGx
xsqj04FvGCDmqB52YsmDDwL2saWCG/cyUJZDoNmLG6PHK4QUMmIVNOYwe9BHxkO/DEqoATNK09/x
wS0/lp3gBtVqFfFRu5fHpxAHqi6UoM/muKk/M/6wn9c/AJhuXoqia70QlFkdxdKo64PBwWTV+MOv
K2ImJr7t69ckOesQw5nGbYVDSRgZfgv09Wt5SCntREeJvJw7aOuUK8Z+igjHQ2i17k+LVBcLIzW4
ioxleolpQoNJVOJD6Vcp8qjnnKWF70jNfQTmZaux6MpRCpWbKzx8fwKvo+4xxjHqItjjCPWZ/xRv
Io0ErKnxxsSRDyEY8HEIIFI/CJ7M8jmfZ3L/grGquT8TvaSYu9tu79l+op5vTtCFpKbD6JlOq4Fi
FG21JZV5uuLrgy67+Qqtr7DBBzUmRiobri4fS6b+aWAA+JUo+nh6Ya0Dynw9GmZovTWDlQtjQx4q
YUVDTi2gyB+Ap8ragjB1+I+l6g8dOtwNz2DQ0oxRN9qsuQZ2jrzqMocyBCdpBt6f64RWdvDIVack
iflVOwXMh1dLkmG/sq6i9k5/K733mvuh8RXL7TVaDZzNISMsxFbZhTfnByhe1QLQBzop5ghgxGeo
XJYPG7xr1d8R4nPgnOk7DE2BwsTLfldUgaF1uBroMM/A5zj5jrW8s3BOXq25xYYxpBd809pgfq0s
0/Gj49QnDuMjJhpRqyzD4qDA5wtrAI0yxnnaBkZnAp4c/aDB5dNQ2mQkl4yilyyYBp6pYRCntcfC
ZYp8nqgKF3myK0hVygpUxhvqzLkWxqdKh0wdXrnF2lD0bFmi1k+dwhPjp0ZwjrVFz4EVtSe+d2Xw
RaWhRQhU+c0H8xAOoGkjH4q9XLO92+V6j0qH5AeVMOel6XvjhsAIN3qHT+/YD+q26Gz/57R3vCCL
GjScUaL9ZMtq3dPIO6fXPf0fYkLgW3pM3VaM/SEHM43cfbCTNerA5f8M9/5RjsjvPHxQ9hh4W/80
X8E2tDMQo/eUZsZTYgFQxMFPvvFF/lQwPTFW+4ZNmvOQGW3inC1Y/6PugUvEQGVqcelh0f2plK8L
SGRibsbK49Rchh0Rog1S+L+APi4q27BPaHdlkUuE8lLp2EmgEurELsWjJ4vQ7pGHdsbGiSHQPZ3W
Wj5hIUkbTHYUraXcPAitv4FJSuOhVCEXNPpZf6dw1mFNA73Ul0e4gi43owh1I9SsgnGMwSlgd5TH
vs5JjpqiPw6971ke2D59K7bM9AitgJ1jl4dFl82qtLss2c9fVgtw2H+e6ZlloaIfVusWijVvFiCN
isPY38170Q5PzOgeRoTjsDGt/tduValdwoUIjtpTJngb1zV8JKTSFFjwlvLQxmEFNgw4Gx3p4iC4
OOKYAqR1R2bHpJNQiow6iUgplc3p2yXFVMRYeEXV36JyJKc0OBbetDese012eADhdvzY6ZYSZxdT
NYsOReL7Bgm7tehfgfLMtuyc3x9AGMhYu10IRc3QYLkDqduo0ePYB2pbxtl6qsj73cUOAHYoS6vH
YETtQIytpmmwo/rxWY7j97/YFKzZ/Pmsbo8ABeFq6Nydt4KOhnEdmLEX+VxSt2IhkKLfFDZL790u
DT/KBgguBe4DTt1n473F1ZJBEYE79KEbfYsOSAyPg+Jx+I2DFeerQP01gy5wilU7flvdNTarFQY5
wAVIqIRk/gcz25XJEBQOHMoSpt24xMMw2AS/hR6RaW/Fh7+E5/D0Q/TqyHEbw+ijC5WL+ualhuUZ
URyw+bUXK9wbGrDyMULNYH+kiOme0SAbkIHlhkEVnd2cQqd2wQqpL2TI9hs9IgcHTJw0hqvG5ggM
48j9QQDIYrmm5CN18Yi5D55WSgTtNHmjFcHTqXryMALL2y1Dkhe7yBVUyIGvk9E9abNW3efRT+mt
IeMrLfMXVyzeHQoYkMlNui1XkaWbvVwCOyOcQn+sojQuheIZwvtY0Gbj9N2ebLDrcEcJYt/wUBuf
MD12SfOyZFgrXKiy9FNfVgf35tZOe5lwvnEd12oN0AyoYWrpivsEnkzL/PqqBHyaM99LmlZ/gEGO
f8sUzGw5Jt37cN5sUjIdYMEZ2sTcbGkkeLaYR4fwmi8TmUj7rmsnwcQESRBzSheT/2y6NVEpRCf0
6KhCe5a04xTJAtfy3i/vQMtDkTv05UdaojtAhGm+2vj6XpG3DxKXVe3hVioqOieqlgCll8DV7iHU
Gi/+DS0ZG+1HPjTKAwaYU+xSWCnqDXApNeZkPb+q2jhCV5nYLJ/g9rRd1W8V199E+Vos9VXanO2a
fHzw+A6yyQWryOOXv6+lLz+0rmLQMHflbMI4I9B7iGenpwem+esCHv+N2yN7ypfHDYWJPJZ56oR+
oh+sgK+x1g0ce5aibms9ZS/75GgUtH5D5Dnyf1Bk5PznsHkmlTE6NBMTk18l/HsDrRkocwbwkwb0
siyWUNfdcwvQKrXfBIEh4MSphl2Tqc372FFoPnb5h8XC3KbEqpS5JbCItdEKUaOzSyQw6oAitPp6
+vl3q8BSE8Zc4muc0dqMHG3SpfZVt4veXTXHPhq3qao0+slOeN0gMgr2ciyGwCmJJsfXxLdz/JOl
IScyufHJqEQ0wQJ1mMAJZdxlpDoxooxrrypVWzQyNeD0npa8IBabgJwOpwNErOgds/86QGS3/aoE
nf6sTdido1qMEtj01jIx0R8YIVr2aqLjWavnmMNff9tkRTBCX+PbMJe8MekI5j8SlwsRGVSXXy4/
mbJDe5JF2bA7gkw40XP39eLf2s2Q2assqz7Z40nqHkv4eYEelT5bsa5jNtDSprNr9KW1tgwvnloN
eRcSq1OslMpxbd06Wem0YjqJmMhSUh2EDjDyKdCfhFY6VLrBvjcO34qn2IW4AnNwESOzadzfGarw
51RWsT148YsjsXJc1si5/sVBiumAwAL2kymuZ5GFEIcv5kd9giwzFRXYDS6TihGEM1eejjf6lRJ0
Et8JNlPtW9soWn65CqlOwSCJ8fgtt35GKlrCKqYD4+j/1oZkN8yV+5sLSvFjEeqOB9z0u1zwEnRj
aFHap58mkM1yXmXmKzYrDzxfZ7ZViSKG/OzyJK7SnHU+kcyd2y/GXOO3HfohfPdMN1X6t1eU3DDb
kyOzg/hGT/N0PG/o0ORLRRZ9kKwFchUp1lz5si553+ld13rr9puZh/85+mOe+0Z/W5EpSJNQjq15
sJ8REoSWZYiqGlxmtfXpyiS0x4cmP1Oq2U6OtmQjKyg5mxkm9OB3u4tGubRAKTzbNH+BjD8yY/KK
/JQVYj7SsJSUFAg+mEjrc8VyPj6vcXRe1CIgFz8ldKJHj3Cvl3azpGHgf+SYd6rWMQ4z0P5EdAuQ
NEgcJTFQ0Hilv3Ew4Q0nac+rdApTcAJlmepc1xXEUkXZVqjyprnj6OC6baDFSH2R26zHoY/nxtfc
g92440P3ScS0bZRWthLHCFh3HAgUibS+PR8DTNACDKavI+A2cP35Y0FGMAx7ls3NjxynRdMdtM8b
mm8sWV27lYDIMMVQFHKxluCi17i/XHf7tNe2DLbzpgAQfcAXS2MqxeiCkkFj4GiJ5O7Fo6zF+1bu
/qhfE2uR53e0fJMuGhH/7sPxVlOc7k8Yz0g4U5oK623snxrq3kffUPfdDbmxD9yQ1KZXEO0o4Ex9
LQPZYVKtF89e8yaPeWXeWcYhazdAI7N46wloqiK9N58P52OQ4dkrT2ONeEjgI2HbyusRawP+jURM
1bVxB3Hcyyoe3JLCXShQqKO03WT7kGyXwRepiOFjDiJSl90Kh/aHw0uqp2Dtdak616OldXASu2XB
WDK3UTQi6nONddG5D7dxB3Dhc60a94cJcxPB8nIRWIRywWH1xz2F6etUV83Tf3tOG8VoTv6JcovC
ZJ6rEDXkzYSfXsXkfEWdapeivUVLzNoO2LjOJZ/pHX0PdW2gnSrs50dbG78XvnhwpcbTPyXDR0du
aaxvqR8pr+OJyDT5jKQbnm2bOmnMEuneu4cbROHvyYsUJIJ4bgRqfjWcUCNgwfm4pf+C3GpBGG7M
kPJ2gB1NaCaKVoG/PWV99vnH05ueAeMmihIY0IycYgOFoyLYMtHiQ+h5C6NMWBCf9iCErZTI+sV+
pnFLgvxZCxfsrMBI5ci+GI+j5ZnoiF/WRHOvwA8EAYJuBlP9/8/puMZKl5FQ0A4mScGwBkTttBQe
3alEjbwA8fYbRb6rik7D6qD0COyk38eQyPCb+qJ6FidfdFWbCO9hYt1QU5CumxMXMzXQn3Q/1n2y
y1GALY01CeW6rPKkXLxaF7iXlZqe4GK8f2KWN5fmtLAe8kAXIKnoNb/uXIktyG992tnqk8176U0n
qg+s7UsojdaVPJdyydBp8qUFLeWpZK2NIZbs9gxjAP1eNGlMPGd5+F2YQG4g47Lur361zXMzr9FS
PNk/ljqUjeuYlUVXJExwxryJrRjtGbtIMlomhVjkvhHV1OATYkJ5gBzdWiDi3lqNhIHO3wfRrv9M
sDHwStbVBxH8kgvlBcA5FDWoiQ7OGDLwMskbI+CT8sZ+NDa1uqNQXUDD79d8R54ONdXEmBW6c9AQ
xErhS/1YfiwfWR/FS1sWsN5Yi2dRzVl2d2OE2jhgKkBHnkq3GFvuh0yug0cS0TA62iX3ArHe2vQ1
JbxbAF2VyZFXMyW0EEzYZauze/oYAS9q3s0IyblnbeSJVnZh1Je9sUyulVW5/Mg47pyxn/cR9Z5/
HczCF3Dt9KaBmvDFjopFzgKOw3+CEWUpVubRwQ66DMyb1t8zZWTmcRuuIBQchdAb5l2O8uZdFM7h
bqf5sv0a3t9iD0iuavs8gKXHM0/q41KEIYe+5yTyooc66vLFoPSKDgL1J1hjPzRYpKF5/gJ921Zm
1dRCbL4y2ZI/IMdJonxZC32RVrYgw2JofAe//j87RzgmEeMRvshBI1A89VROmXLYcARetTQuljHk
ebzGWii1pYCGpAVRys8yI+3lGrpuwnV/c9nnEIwxEqEUwQOWVW4uKFDoivo4CS1CRPOBiyoLSJ2f
A3gLXsYS92VgkEvLBzLb4ZkaRjQbmbzkAOgsfInx2MBUH3WRkcI73IuxfphD6vHS4oysigxfAJ6R
ETARjkc9EVEktlSu/CZbYXNNDdgUkHx+gMcGJBpqasmysDt59LcTqfaUW4sxbYQkjOKaaivCzh+Z
KLetdTIFD4nMw0cMtDc+YTzcYF6gnKNLxzqQdqreq0w/JPM1GmVfcYyZg9Vrz+tDQt6SKX7xp6eb
gAFpzkgUzkuPUURPmkm0wy9m/OJAUhPCMAG6DYelAo1hazw95cJ8gGqJdE9BNcxEdEcaY51BaZqs
1zkiV7tZXHYzMvTEGhzngVRK7l92y8GHYd6gCiEiJ0Kte7/K+BxVZye/Ug0zMTuLQalDU6dJC+uh
GVKAwbalJz7hdzW+USGuCXrn/k3Un3Bv9/p15XnkXQOug7CpNm86wXcvrF4K/Ob3nHvvGPnhwV6i
5SHDD+OUvcaJ5duNoIY5ZfNkrMxJR9uBCMjs5+FuPdgb3IJBQwLTt9kTsYLvNme3eAlfx/g1eVyo
JT2FvLE2npuxN07glA4xsnIQ+nwOGCJaHSijlJRhZ+ckrYGEbDFzoTbkW1ZApzPQwBbQcasW/aJM
zcjEb05x6cKjf6BkPuu/M44C+vVbp3L1Es9M7dEnpWuNBHtTqiVugrQ0Io9tUSVb2ytVHa5h5NrK
WpP/jQVJvqz7hJT6I2iP0coE9+jfVMUqXBdag3QARQFpfasdg/YMozHwoYOGy9eGkHy079m4ngSX
eDIALc0o3tLYr+l9TbuVfCV97i3jSCZkIz3xA9q85L+Gc6E+KLb0QqQimOHqlzKLS+F142OBmQWn
cvxscmJnHqkKoE94bYjiMx8pmBQeeelU55ZGhiEvG5guqR/dHAf6D/G73QkTUYDMO04SSlXsPmED
0GOSWBv/10DIEpHUyPKRi+zlP+udADiYbMsf75H4Jx1u92ialwChPXw8WdQPaNmnXR7HPwHk31hv
h2ITex47xgSeG1e4zdqePgig5eFsyMRfhEW+z5zP7zhke7T54PCmXWvtZCS5k6WpwVHbL2YcH9I2
SoB8T2gCg8oMOh5j+LNUi0ypCPZQq6W3o7N8cLJJ/4U3QTNvm4ErXt8Mf+S4uZLwgpk8ZErIKzAV
IdigwXUTL8Gkey0OlTdCbWJ/zlBbY9PtHxHNxcDqO9GwteOfKLmBUBwGo0yT04F5Sw1WHtWx6oUD
gM9AiWhFI3a1c/bWvGi1JzlQtOi3kQUvMZ05gTCgZbCIZwAJTEWi1iJtj3VebmQGIGrVC/TQs8Tp
eODtvDDGfasOwSIsQdmKb9AB2EjGSefUNenBx8c3gvyY2RtS7FcLCm2/Rfppkk176PBTdYUe03q0
xMfYe2JOW18MQk4kcj3y+n016g8dz6U7YHXHJX/9Tm1LGsQatS6gqY6RYpyHyrhHpez3TFhIPKow
rCS4rS8B8Y8de9td8CkTK3ZM3QalvSCy4ZKGj6kTPVyoWr9J2GZYlleuZtu7uBC9kfegrjP1w7TF
D7FrFS7Yx16/5gtApOQcBHjZfLboGV/981Vsv5OhNqaIjs1f8k+TYe7fCC6d2qyqfHejozLZTzso
uEyr+KgCOdbrs/NHIxMkn2DPJptLKM3gkrG8HPIhn9q2+6fM2XozmfDmVJr6rmLaueYjOxBy0T94
aIUpYZ7JNpJ1y+6qTP+jT9KwJ4sLOq3g0aKaIZviIQdSR2OYlol/Ng0vSEkmW3g0ZHWxMDsTC/jS
th7Nn4yZ+eWLCwhPwB81xyE9BBLpylxcb82U/4OhbdajSSWUY+j+3+kKpSvHp7/PY/gwTneDbSpK
i2WZ/cHkdGdbX7Q1v2ZZnI1KFya2DHdijMf7DCDunjp/Lzrx078rofmho+LdityJWPzWqDS/wruO
hFq/wjniVEUmtdNupFfhNKDCAPk4diXv2s00FeqEUH20FMV09UfDmawwMLPlw0C8uvh0yerDXibd
hIo2lUKCe3P36hfQzbpfFo9Di3SDUmSrALYDkwMbFHOvDN5p9k2sSCnOT0uF8DUzJRmgKWPu1gd3
yBN5XREpORlZHwy+xfbZScGT1bYFRdCF+wdkXQBoX6vGdkRJyWStBsW5bC9Bx4lb96/5P4PUEY57
mCcxcDJwlUJw+sWCfG66Cd9ZZcE6f4w5nFXM8hb6vS1/dtf4hOAC37lswweunnCyThW1nwACj9ua
ygq72j8tY8fKvmFEY79sSQLWQsGJQlwwCLUXZFX5YwFv2Das7LBUCm3K3+ISIS/UJ7l91sk2p4U7
MqIyErBKWt0+H+OCGYF6CJl1OPF8RQfuBrk6JQmjXvL/ay+o4PHQZmC2uObV7sKuuVz28iH4xKSP
8nlDvjnltkMebPADvxI7N/vHjkEqdbLXP7bcoT8WbEa47jKP5+SyNOxA35QVIybPggEAw21/C0h0
bS/nTNY42pYynXJumY8bPA162YRJpRqDs+P8oLY4fxE+S1Vfq1okGLLymbc68f/3wMH7lzgsuL6H
3awOFg4CF+46+p9YhIVgWG8lmidTv4lpv7/LvkLD4/9tTRWxwbgD5GI4k2tuzW6zXkl0+D9eHa09
mxZMjX3z4bX4wxI27b7JRbA1B8pwjU9SJn1Zyv5v4qW//Llc6G8v1UIBbFG/pSCGTJUajryZoGVv
IwMyRC0cfyad+nV4R9aOAZjsKSZz19/2ftmSiuU6fhs+O3tSgI0/ajYSlLgCn1Myqrrdj+kjWW+/
LXgfxqRpYglMQFHnb5eGIOhw0YACiArhs5wk5g41CU1ovXYNoTNyTK9nFvoMEkZyKIIGmXWptwYK
nlX8EKyjsK+hGTlgfJmuUYch9Mhu2DMmqHt5XLHHgHIc743YpJ9tlKjBLzOMum9RhJ3rdIG7e2Ds
UCujOBl6Un2Lxr1cTyUn/+U5VXfP0wLy43GVxToMb6nSqgsBAOo63/JrkFomjf/RX78zmMFjMdZP
gUbt2+CABV4U70mpq9dxF8hNAppivM7mmDBKA7EcpJagxcoW8d44jzsl1OIW6FgOITYjH/MX39VS
P6hfKODwF13O6aaGpzZ3OS/bNCuCqoqJ3BhiBYF8Ncf8EzcrAKqDQDX5x4frqNYXqqJsp2jzEpfD
lELCQoEAkkK0I+z0WAXzAe4zQYetMnSgH/YmVUUNS3MEmK3HieWsV8mGyBW67utuN/BaFFrEgmSM
TcFyUqLXewvDLAyhE+Tr8Nm6MmeFaLXM25hPP2kYbKXH0RyiDyJExUVfa7gLUhGfOTqcy4l70461
mvhW3lfjgOovQ83Gsw1RiWyjVnnvlmReUrgGHziUWtCXGXaxYcYbF2D3Kj3dsvEYqXFnQjcK9oPw
NOwI+CeuPBuhTX7T42+ZfnPMJ3WJ8QzmnVxcxpe+Wf0gEt9gJuIDSq4uYVkxXUMrJjjdQ31VrYOL
qIcfeU/Pojmo1lhHeWp8Ue8SDM+/n6+yOFqeq4ekCE2vNkraCZz+Raz/tg+iOiUPCRTFrostxyn7
erlKaEAirovOaPPKA95xzhYt2pDSb4bPer7Ejp3UCvR1jmsunKRnIuKMefGqWTKQhzh4FTiV7pBD
/Chgt+iLC/bQmh31T++o45g/dvbjC3vnRzNN365HQ1tJ/23zfpBXic5sXMsBBqAtqEGU8dCvOif0
fj1hGJiyHQ3TsLI6e9inSIuli0htlY1WlHIZm85iCPh6MqgCR/Fag+Kx17mYhMws65UqYJYWWQpw
8m0r8qfsY1xQ98bf/ms1QL+EdK/ROuMFulraMnBtRMROPMqdz9GLARxm+5QYP4K5BSBXEW1U+pEw
Lna0n4AJyMxzVJh2br2xPFTRvCKjHTOeHCemZX2xwzgH3Pn9GIrPc0k9vVzrs/SgRJY9pgbUeRrM
BCkbQDucKfvj09CYSJsn786/rExnHmXzVFztJ8v5ryV4wS1BdNnf0EcC8WnP8y4s6KnS9BnYw+aC
LcOj1k1lEKDSvxHt2PVPeBwxGtGnZgmP0/GmjJpotctD+0+BfhgoAinc4gPSeujAkCg9Jz9lJzqK
1teH/h1e5EvmEgKGZMyw46N9ZR6RVJrqMYCArE2if+d61jhL0Ioeaf+lQkvMUTRTjJCtYzVAUYNX
hoyHmTCXt/2BblC5I4q34PksrKp2ovbvSAHaXxxz90yQ26uiLc9qjcrvFVe6XM68pYN+teY47KQw
nYQKXP7my3Ne6awtR3q8y5+WhiPsfo7xlOPMbbzMwmVFPoYPbQs7QPTaB3AZd89c+M/vdIyJSOVR
uFrJovjYZlm11qHJD3ZAGgyM8wtlMBiZ1RVGKd1XVT9+LOJEBkWIZcwtMPiDZ9K8w0ML8qMCjcMO
jBcBg6i8TfzRhe88DZXGaOzSqvJuGqQImuz/FRlEYlXtmnweJR8e70dxi4ObUv32mULdTLEl8u2Y
hTU7oDjEXz2Xkxs1qV2E9+RxtbVWGGMFuvRQhUh0EqsKQS6uYxfUGa1hHhKpOvSRhY9qZueEW0bJ
c/qAapz+w9rOZYi0kNFAEfXBOOB/VOGdGX7ps0446nNLrd2miH2QNxmJVXuUMzgcu/JH/OSQIwO/
tV/faPIoG6FWkyixeOMmm5NeCSAjMdw9QP6Uec9rADVZgBG4P/oUYuAl2D+MmH567aQtWxIBLGTL
RlSS3nvricZ0W40UcXncu24CwGE9I/AicXtstQU5kJxSKXpYduAaQt6M8068E4XDYH5RxIMsM5hh
DJrTWtZ31X9CHxejnXbrZP1TVAH2VPCCZ2ndUo60L6uCwXBAY8BQDgn7r+XTRqV16VwgqTxKujgQ
3fu8c/7Y8f5XCa15P71bnqTBtueaFYmvICBpzaWcQxwoB6o4NF2DA55KzSkwbVhG0riEcLobmpWq
2KCWsPeFr0l+FHEIdSk6rkhb+f9NBNJ1wYuWKRNGk7yjPd1c03cNYMMh66D2f8fWdjL5wyKJ5n2g
kyMirUFXcSuA1oWLJHgVaPnBfXun+Hh2A192vZuclVYzh93M+GH9P7f6QvSYSr38EqNPpdEolzHb
6sHpN3b+7nzhkiAUP6BPY42z4RYw3mr/GM0Xgjd2rTKViU2j15zZtHrTcg7htE/0X5YAJJ9gd1DO
ZnrkwYxjcqjb+QQyZ70Buq+7Lwx6+4nN4j4Eu2UClLOnLi7k+S5XhtR84xb7hD7a5FK+FtF04gOe
FhgE1OvBXOTUP49LaEn2P+gg63SP9cfc9JvV8Uuseni7zf1krn0JUIgiyNPNL8OIXYkjy2+OYpe9
Nx+f4kpWwT1ojNAfdF6dw8WWqwZLPoY/cHznosXqTuexvb5UKz8K5SntpstePQFIW54YfgXJYCh+
VZsusyLB3HlMvnXN6Z36vvPu39koQt9nYYRJYSEyTAi3pva6olNkUZhx+E/NKoZMojg+w1G17cmD
7kNH9f32aowvvpRTwIckMFgkCC8vrKp7PlQKr2S4dIoDPmHJbOIwjldvRZMlusGHCSCnpVB9BepZ
0rlbPbE2Hb2fFj5g8UKD7Mbj6kd77/kp9zNas61CkHejkZf3XC8mHs3pmcUdtLkJGaMwM9Th0NWC
d29F9LQeLNq7co0qPR1pgJSZD2xkAeTL1hFbKcJfTKGW06i0nq9euuBPUebXE8fAJBW/lwWIPI11
GLk99Fa4JI4Kg2ByUpcUXDBGUpOhRE3EYrv3Mfw6IB4ppse+pYN+r42a60C7F+NozVjW+s9ZlpsU
W9or69BSy8zuXrOZhVP/i4MCW1KswFhHYB3jmn7x031vtuET6fcn2fjjBW8ssBsL8iYqEcZob+UN
T5uRfhl97vlrsBOUJJGicuJeyvsV/pf8W8aZ52wdYTr40dPHX+IfzVx2PFRjVrBBiXJ9oAXET3Od
kn51X5VjIMdb+gYePYTydLlHpvIOHjC2VZ+bHdufXqPr10R3Dy7awFkdIM7Pzm9zqdz9itFcQKw0
r/Ps/5YcWT1qIwyEzX7clt4svx8TYS7OJnDXpR51v5Jh4V4ocBqNI/twxpMaoOg0uV8ZVhRpahfo
2tm1JqXDQoofUtEb0E2sbNSxbZE2WuBtOtDtPTJinM4KpoIh9lr9TCZxHLWz/JDhi2MtzhT7IrgZ
S3UQIdHOtcFzNaUIHxRwB43IzHYm3eSOREBUTxycDrmJX5uRaI4B/cw1aEVr9BOw6mzX9l/Hmjhs
SAWp6Ih94vhURT1GXVRmfqo+ArhXm1L8eZCFr4i3YOjeE3X31WgF9SwHTkdcvA4aIx+W5cPq90em
kR1zshH6YVSfhDhFTEmIFV1mkONq4pFwd0tnBPtFdN7gLRaVbki+/yycDfuRLiavR4IW0TnZ0n57
ghAzbWnlL8nzzFD9sWNoVfwl/kSPdqCs8BPzGMg65SI2sO7nmAVJHi7xoDdCHwdvW37F3zXn4sUL
vMTWW8l48j8SrwPiHO7w1EkKNslMcKMyGeRlaGd63mfhqliQIj+3VJ31UUxB6TFjr0aOT4wxdZme
agJhqvNAl5BbnwAyOzBQglRT28vDwIs4Es4HFV/GZeHzpdPuZUmiduvakiR5qQHIjgtxaj3D6FKW
9Ic00bl5O5dmLrraZo4RAPh/WV3JsFDH1kRB7Fx8/kywMfpg3qbNLd1FBh6Es6KZtrAnDOgoLIFJ
QcG8i+ElN/e8zXz0E4ChFp6GsWNF4Oe7385vfHzDC/rvqpQPPMNri4iEWfKnAAUtlLSlL1iCwXtS
ve/2W2OZDTgsWYINAMeKVf+vZxQBK8c0AJ/xLDCoVn7w6Mgm2O67KPmWmQ10t+K7j43mbIZif6OZ
GY9X5NUYT0Pyk6wU8gZsDNXP2uCDBGKS7lUMdi2eh4yzbqqf8mk84zGsMzqDUYk65w/yDVwVgJuX
zrhxzyMBhxAXM+hYELQTZrKohPM4mw5URvFzu+brhm+rUbqO0k6eqrshJ0gnBRMv1Oxh9GcKx2DQ
+8bc753yr7Fh73nxAI6CWaUGBijJMxMa8w9i+BAnemdwTTSb6Or6ucoPktQuAYK7oAYasHCdw/gU
kzDw03rCqLB6PNEPKtvv0PS2iw4qBfkbksST3q7NN2NsWGHvUms5f57OEP8HGZtHI5rUK4RN1/6R
nu0eIJm3Rz1VOD+FsO2qMNieJjPbGgXWIC2qFOzPuHyREi3mU2hq8KVJ/FbhiJPjUO2BBBkZzpVE
48bjqzGgegaz8YbkW54ADLX9B3tTnchA1V+bcr9jqKK1BPJmhO2iCeIUzlDjTUElir0LXtFc0A61
1jD0JlPgFvEgcceXH+IPGjxxaP6l8V4JfO2EI1K6koPhpJKU/3w8EdfoiyF7IzeQtq93pG9nITXt
PXczPFVs6GBv2u8wGXuuaXLmFg3MV7xqPYzRKf75VE2Rq0wSPcC2JWb2ZXKBWPEngABVqBHrXpbW
UtRiv5mKgOYB7u1WK3WtS0No0LTgFQZy8MXUKFjjl/qkk2hh0dasPOnczY44QKkoKhHXBLn3DJ98
2/S6kC1fLj8xD8HYcXgoxPO4t464+giQ3g0BoWIcRwe6/gn8Gt6qqHqRkeLrcosEuZyGX7BdQgf4
PgALPG8XTw4ea06IPRyxd2rFiMK0XnbZf2na6BR/LE+Sbr90KNTvUxlJK2lvOrgmA6SK1TF5iYlf
rDWTywhrjxj3UwxrZxn4rnHAxy8INIAi93E6uGwdYKF8KLieF+HuNnA2NMf8bJRhmQINLjDtFh96
5wiknkU3jitE/42kehBvgnD7MqV9+XXHDlJFrJwJhki5sb+UEtXT+qBqaiRIa/J7T8mDq12NY8+D
u1yv9qbWKcFflJYdJaEo9KhG6Q8wJ4zxRlGGVKQLEOGkdl8Pk8xXc1ne5qEnqYsYOzi5uSwXiUkY
if+9YkYw//mjegnQeqbUTbqpO1/1NB4y9a5L/MuFSfzYy5/akqC+bRLP5Se9p4Iw8K6r9J3d6ajh
YZgt1mDPvOdnvoKpyqroRlacJsFe0L5etNFecP0Yrzr6JsF/SyqvY9Nt4mpsG45yKJhb3+3kbJkz
cZwUjTR2zDf84jI8p8RSjPcLJld3yUp671P65wnNMnwTJvYgriZ9bcdpmUKiuPX32IywBbCVn715
Nr/j8hMu6ZjdiTqnYfyYjTmwTub7ncNSAnJBQxyiRrKgHCDMqNUxBGHhALS/fQxt7Tda42IFwjrT
YoGg/a4NyV4qCMk2xpG25/7nS2ZaQKgaJpQWHuCahtR+cINT7W5IoTUBUYRfShJLluFYlmVigCdJ
+w01Vm9wH+NPuzbWpA7jrSqgtmWhPeKn0uwkVzSN+sdffNX8UuTjYTdppNi6r5rxx8ii1oIeGZkt
TQyWaQwNCyGxLVY4wIEMlAO42PGVGmLiIuiBsKD01FJjNI1N3HIAneSDQkD4jXGY7bqBWkGvCKGE
CJCJePI6y9kiJiUU/tgIPbFH3Sfnp+1D9NGFqVLiAgY8N+upZ8/ljmYF54+ubDdpQ6R8dSaAqNDN
Kh6jgTGxmDr+RX9chDEK4UvljjyFi/aT43I9qX9/+1n+SybLieCI8ZKicdgx20Gx4Tx8gJqy65F1
d0sssIEPgsBU5x14pY5t3fQBKlvSXeqOlN0/IJOCR6MJ5+NVpByR0NdVbECX+nnR1wes71M/gj3D
ccgQcBWLyUIJXnUZCGXqlp9+Y+N5JgEe5N/gB741rgf77Jm1uWr1UVsuWqiMrYw6UW1V4ysVbojz
UreDMJuHV0RzwWs/s/c/hIc1gcgyk6pe6uYNgPjgWgJ56v5azT1j1rZDiSIqibAn/69cEgoIn7wj
9bZUYuRIgwEK8N+TwdJImeULFAZxLMzrm0agQZI2ZqoEfWmrWNZ/822eTkQpA869dlQG+/oC+5KN
SlPtgmsC/4w88IwrMiQx/ATUnyIXlxSCwaJFvpsCObP7jFlfO1r4NsTko6qrfSiRQS787/ooiwcA
k//LxHc4EdcLSnV6ahByd/8ZSxaZdjaYuKroG+IQKDgoEk+GnQ/rYCKjfLzvuoa/EJ4BHAdxql07
ngOiEMUSXz+UOvQMseevLuI8rYMaDh2+zjfHqFmAP3kxnm7ni3vAB5tpEqqQ58jhderG0nBvTMuO
5n8y8fCiVFbkZmePbY/tpmAR1AzHTOCW5NCURg2VvWToNVa5xguxd4QHIJi1C7/rp32yQNysXILU
GkfZ3yIHOxEQzAVywwlO2srv+4oblHq+ZnVkA5+26YDMsJMZ2LbnPSlhu3Wc7UOa2BNlY9jKYigu
/YLS4Di7ibwJDA0FOzFrNMfailMZbsHwbC6QF7DEuQ79HK1yaBUc7mhzA/Bv1LwE0AhM1bFoe838
LJeyMcFLcpl6hEzwoBEPaEbpTozm2X5k6rjKAny00btsrPj+9erg5Jd4YQtgl2DFzblpMxh475g5
S5pP8uLuZPGsTjnsfx+SggwoP9KuEfdgKtXuL7eQjh5praTRzNCsQYMnCFzRmf9VRvM3zbCDgWnD
7CDyd6sF0kyX+ya6y3B1oadJfR7QiSo7JlGXh3q8CRtriTF/dNQoL4jy053sqfkiSKBgsA7gJEMD
mZnFSS9rwNc4/9+rqbjV/5DqDhykkPOtu4X0fN8fo7ho1hRl8l7pndMXY7Gw3pMOr2+056gsvsIz
h7tXzD3BvcLriRaiFb5hJVgmiGt55A/XsYo1AnKhE8oo593knUT/q2RbCyrZvybiQ8oM9ml6rNGs
S2/ZUvzyTRYS5MrK8E+vwzv2E0j7o9dX53BTeAgbj3ICv+rjIgo9YpELEBLjaoQ6w14m+K9tnyAL
lXbX4ZZE+eJ84ZzlAEXF3r1j+Yy8QENRUEoszo2fZhQcRGGzGVVflcsJZYXVZ2uLVQA3fqK1KLnB
eRXoJmcX+zSew/+nkku1Vd3WdprJ5A2aT4ZZCtgt9786AAh0My7+2TbXe64pQXUXZRhK9mqeLW2a
ySBwzHbwOFfXKxrfhTGuyWJb5CTfVhsWArR4auHzn6WBo7AIlKM11pfqS5KjfutCQVJ8FlGygvu8
KL1t320eqWnq6kHAyhRHhEusGqm+F2lVeZNpIa76XfEdXRgtdajIY+A4psch9q3OjvaLZs6Ozyax
Uj2HEUi6nPlciCbQ9caOZ4uQo37KeAQZFkZAMMOxgUme0jNV4yJ+JwznkEN6qRtz4xKmnsKJDlxk
+KPtPSBlHaooK3fxRZoG5VhqSyxAB3ULI9PnSXgJZ7bZxMLJVWr4w52VxwnGE5rd6oBsR4ksngE6
GRiR7McuGOuU8gHz3AiSHnVp/2xiUHlY8kzsNT72oNKo+GUU3ipb5n51Pu81g8UbuRD6xQH/EKqn
868oZ4kPJMrHgwNpelU+X4ktfVdS7DPiRKnXiUGaHyTQ1YyaBu4KCJdAJNiJ0wlxc6rx3JqwmsSy
QmG5yFq+XPlNAOqm7orRTSTEltffKRV6/Ak6Zx5C/51LbzPV33l9ytt2bWQuySIeLCW7Y/Nh0d83
4WN7z/XBOnF3ExddyJQ7rQyCRxPL/xXXAsi14GBvg4b6JDYx+00F6080q1HsEdjOXXvotNoupnuH
fALQyS1ux0dWXD0VL1FmtIofzZv7ymx3Utvb5Ee3HCXcqyUNK1+LWWqehLHmO57TnRMXABcgFdNG
eHrobm8XFLVQ6QpP8riJlZO2WAO6p81L4BOrugqfAQClVq4a6tLDukqOM7gUJcuJr3aHWwDDPfZW
vZm3BJuz48A7JBx2yIy1/B/BgxXWjJNH5UyEV0cIG1ojWk1jrYP0HAW14od6YXjMFQ+ay9nM0xtv
VUDxxNqsnu4gEsLM5Vm3xJP9J+1vE8QEw8F0N6unAEYWls7T210c5GAD8elr3fFzMKeNT22eKK9u
FISVzv+5Znfyt6WmZxSaNN3KsbcY4jmOdj5wjEqt/wyDlZI2mtdUmAoBTp+M+/F349kfPip2HKhL
XmO0O4jOYL3qI+Ot/kx+lyjzh8l2BlrDLch+eMzMUUc8Xl3XS3Ukc/axLxhNlco0d4md08gjyAvz
TdJVqDud0dg871Je7bG9GsH15lNzQENTjCTdn7V6jcnZ2znNDRsjjex9BkIJ1xJFV8UxH0GDcKua
Hga/J6mGkTY2zqrhpGIFW+8uTdCbEuAUJFZCtcupL6HTvgER2oOoaYz5o5jARMAgn4vUpHGzFU6w
CozAy+akfgI4PUGoq9pV5IUFL3EwHXkLxrixcbPsktLcIsHnBg7lSk+UtdyFhy+RBRa1Fk4YKow1
lOUXoaHEMBLICwEbZBJUxwHby4mPAf/IjJYC6Q8JBCt6fjhttnAXN+ndl0KBJr07v5aXZGK9woNI
WgHuup2ZGasVq375YpCDj+rtoQX37YYCLZLksMa21aJErwbOTT/nuQtm/3vmiRDu4HUAnYVTefYZ
yrjttORfe2Fz1T2Kqjuk8yFLWJPvPt4azTpgZn7kxf00NFnWgqbpSVUm2dlV9L/D86Gqh16YUW5Y
EdbVfKMaJik+zRc3xqlOAhy0TpJSPVtIbV3Yt3gngs89uAhVfMotPq7u/UPvpURTf6NPZS4I1r8e
RzJ3TNgTE+w1VyuKqdm7jXNa04kw7kzmpM4fjXmQunoQUvoaK2QKzAZm3jPtIgrdldhnZcWg3edZ
KKtSw4a6i7B7EKEWJGb6Lqe4K+rUB8mZXBoh8u0l8m1/iG8ZaFykHDHotKu7hThvdLpyL8iK1SCu
mfM1lgdHdIjLn/lPw4w+FWiKcoMAttxCIEbZNq1toxXlKjUWn471kcqm37cYY/7Cte4yHEkELlMy
K6bVPX7cQ6uOc2+wiwo8R5BDlee6JVty5Mb8h2O7wAi/F10jCYGOVlfG9IX8KtFaZgR4gHydmw4j
viaxWlml8cHC1/eEz29H6Eukn67g2D3BZyyneigMw4OeFn0n+gmMnrw1io8C1G/DTRCB053KhH7W
NLsnXTK71mpZe1x7MPQ7v+9TzsV4ijipfOPUmsgiPlaog+0nKSegA9KN9MM4LnZ6mxLasy8Q3GtZ
AhbC4KWtrnAeXB/0g5d6VzfQ6aUYa/JrWhiYpxVs7NDpNlowcibrQaAsUz0eEeYzMw/UaVqtmG5D
ynGXNheSGFrHqrvqIvEZFCzTyLIwtpeqj2SuRC5XcDUuUbk1rsEPUiIWxVLD6uVCUuXAicb9xJgR
FfpP62ZgxJ52eC97pnapiPOVHE6Qe1puwctwx/Myc7EmzvDjJ+QnnVtq/o6eRz7ucMizips2sukJ
Rl0P08uGHXEZvtAQ/TlP+4SpMCwsEKUCqnEbdH3wrnuu3aAFG12e/HEQ4ywqpp4lO/cnHu6hY/Ug
qzS+sEJT23r5SC8jLjQIV8W6Krzy71Nuq7lQdADipXHfYn62xAAlqgcNeYpAGU5vSL6jWSRtEgmr
FF9xdjNHLUOn9D5o4uNGHpH8auXgKngSWR/ynxUjLvHseIE6dOOOLNkO5781DyQrtrzjHsGZlTMi
Ngfc5UZ5VF3I4cvW5oVzYLdCN0ugvUq/aOQw1h+7DPBygcjU5U7I+cenBAPrO+jSgusaCxruK0F1
vHFZa9PXbvEW/ySHBL8q/+pUS2taMpGH6thwiaZpI0nk8jGoebUWnOAEjGHwhZRkTCuI1kGKdMgt
d5JyS3uUpYUBOmvI+GWhRoAAFS10E6o2h52bpQBOfA0pfTelFLR+ICZY2gvX9aNokgJ9i72cRJcF
Qy2GIxYbHLYspv0Lu/L/VjFAhFk4CoPaJa4hCrCl9a0cUcTpg/P9nEVXPvRhexAondoXjTMG7JeG
3REbPJRF/Qeq4GQa8y8UE4mh9OI5rN9NF6yhy9wJyVLM6os7vw298ho31czx7fjEU9VYYYwXOb9c
cQexVtw7M/EFZ2LRz3g0mt9YUjLgijiqV9dIYS78r/gbMbMLDoe+3u0nudoASJpg/0b3P3Hif6Qn
vg6OlxnIt61PzweJJuvTiXUeNcV06F4lPU+0EjrqPfH3xFsZrL41516+VwKOps43wUvMLl9pu6Kr
TCTdmsmdxjem1IhqbCAtJLqX0TKvm6iuMDEVPyFKfCyZtpi/S4eQEin8s1Y7gqV3tfX8YvEMtI7U
tnSaMBDMA8EOEEBS2RW5kQJt5v0GuCc99wy+8N1Lt8fYkol5wK4UEi2tTkG4g926D72wKJ96Pd9G
E27ds0Jpms2oWoflN4BunK8gvhLN1y45N6+jsvNAXW+wWyFpAGGpLWALWuXxyCOyUwlZcpgdj8Rc
qlPFcilTWkWAWDlCpHBx2wOemneYcPeQiss6gG8lbI70WRGVOy8riLdUqzDoVFQv7FfEVTaE6VPc
wPwRhillwdLvANkJQdqUO9a4tljs3qMaPp4fwOqAbaxtEzQvSs284jf6e1k9Ld064h7jx6OzK+iG
G0K99rc5Q48zje7CO6DB2HE/NDcc4pxrypQsgp6YEQ4+/orC2r5P35MwU0AK2bRd1zd3XflSrY+c
x5THaDyNF3RpF0+580PRRNg7louG97AP5ME1YOdgCUf1AuWXEiELiIDQ0CjAg+/lYDX3yUoHXf+B
DlmaPlytGJDnbfPNx+sLcRVK99NOCQbHVqpfLhtG4HiRYdJ1w5rFd7aPNyFBLhl1XHpkW4IXZk08
m9JEdfgKqlr4JdGZOPof5CPHY+epG+Owol+b3O72yRKZVzq5NOcvXN/sdTlbMhh8R3NVdEmBLXtD
P6Gbk/6GO1QQATg6otXnwTnrkS/V+TrZO9zEQKzkqRxrA01qYZWOXv346zzrChrybJEjtfnF6uox
GxfYnwe0+FxubEtHEPtqVScxXt6Qe/XQ/She7fC4ESm3PGOouhbKpMNuZQ0pyg9hVUQOeAtq1KDO
zd3jg9qtNcKsYLDPpWvWL+C8yjyYKsf508i6fbMFszVTOG760WOzRFxNVL2jUu+V6k4zB9s3qCp1
Q1aRW0HfVzCHbquCUUc9Cyv/zoheKfVZ+DVz1fy728LTkAtGt/FkDhhpOWAYrJpGFzO/i7DM82vZ
p6qah5u1J1X+VJJBxubKxn+2KFCKdnrTFHu8MSSSFyse/hCLA98vrBoSMIsv6rbEsPYqN+Wl3Dko
PifGQzqt2B2lw9zYVhf/rYSYKZZQXDZ5A3oSunMsIvMmizwEIwuA/kJGsVRfHTCybjmy7XPnLIwP
ahOKZByu0ICqdt9D27LX7jWFqYP3234fei1xBYr+g6OmMfEtahXOq4St6I4J2Q/TbRqEVFgUr9qA
V7YUOpyz4befQoeEgudn21OgrZdJPxfsdaS0HphnI1yma+a243lPuUiRsbgwaapnt0awOMpoa8oQ
hxNS6kzE3ZBF/74f6UM+IFbJuX9/VlqE+T8sT549r9qcU4koiLBGczq3EC7BRVlnMyLWtEOCP6xT
Jxw0P3yk+8B2ioCvAvy2ER1r8kCYK5VPBLJXporMfcvAtt7w+/3/KBpyUvZoy4ulkKxmin473oer
RJOrYo8evpBEy5mmKgODgNa1jC7+2hht4OOSU7/tP8xM1Ez1tTyB/SHjpwk7So6U/OP8aDPktatM
WlMYdfqbyOylUUsVxeS5YpUdNBh/kgvzxXoDVLRDLFKbQQ5iI2YJ7dSwSPwpSypVc85olodNYgwA
8vs8p0oIAk5nfxp00P5s7lDobCWO+JgoSr7YyJSFtDsWniVdxkugsChTX7AyEkn1VFz2purG9Izw
vr3GQvtb/2sSmLO0KtHQJB0lbDyQcoTEYoVO5FBxsOu/T/3xTwPaKwOgyE2yZZ//pWlcetYsE17j
Z9OHtU5nPWJYMHXEaUpdpc4RiGClcJAqjmga5lIzceHCy7ViohDHpa1Dx58ynTfSjOdZBUEBiu06
u9vUkPGgaYILLVL/qPqFhSfolnBBpzi/v723FFN5jX96X/4brgH/ZKs20WrfR2SN8AQS0j7NpDyF
IT3ARBRxawp6Gf3rrUkvRuZv1XxjSCXRbp7YcnQ5ssU3rBgQjV0qU3rE35ojabmBcF1GhT/rfn2Z
yiB0CohOoE+8wuOVZPS7K1dCsj9IZxkfiaU5xeXSfGmHBNsyHzunGcSb+6k5rjyE3tI5n8j7aaLM
OktPNjhG5T2gfKrXUAQ1gLjwc5x3On2nfWGzzgiixnfkSOUSwbcCNFQozC8IM9EFDNHVxV+U/2PE
Ua5RpazjJB28h7towydrhYPSlHqAEdPCFkS7W9y+HnaSZO2oq/FzbVoEsSf08Z2grI6U2ju9cQF7
uXF5gtfyCUV4h2HrQ5nlPyJESPzA78K+yVS2EQG+Dd99Tyw6WCeHoz/bB8h2haogt9BkPWb3K75d
ZVBrOUBUmZf4mtdJmTA+19VYCGTOawCHUg1HbXdu7OkkdKMSf1RVHz7iN/RnUvL3juzFeNw24dEu
XYWxLek2NoVYwSoDbcE8KamDBxk6ZjCqx+gfhj7m3aytWY/lkcLUE0VvPOYc+mLbF3Kt0ewrTBb/
J7Ecg3OxSfnY4lQrRUulfwETPwhiTuHfF6GwuCRAnAeuMklxJE/m7cabX0oz4S8smtafN8vfOA5s
FcFnzKTwm7I9YVBV1sjQWAwrR5JiO1xvwZdb3gAldMoIAPvxnOOgrMSFcm1gihOCkvpXbAgbJ3Hd
RPZONqsQ4VJAb0jpH83RE8WYSQhIOYKiBs9ubiH4Iw+Bz90OATCELBwQtH3yCVB9hcSCcqVglR4j
MMXL5LPg/gYxPoB2d5wlAEYKzFG5wIgCawWwR5yuM4sofRKcQWzNwVqPKXK6avQ92irpL1TfB3HL
lhmZmCJFap383y3wiXF2oy6Jz2k2hvX6hyxi2AJ+kpq8s7eiVhj0OWeP2lvcjAR49xKGYK5nrkfW
8hXpQcP0v4/Kkhblo98CGpeNFvl5NU23XWvNO6gOUZj3SMQtz78eqkz3UInmJSW4s+k6wac3U0Ya
RDKsXqlZwqOQfIZnP/lZ54m+iQ5HQXKJfDNzTXbLg8vo+KXOh6AW0VpjhVfTGC8LYNFvjvCuOJ84
yg8VVq/tXGdf0mQkdR0biv6OAxtX751UKqhjDwrt7eNB6fioDCJiix2M4CzNHQAmOAvt4jlHVIEK
JT49kklWpB5w4oMNrkFjV0/WZrV27bKzV2Dj12NFS2fNveAUuST400bYQBEnT5lj1xoSqjWSIccP
9RYR3ocEQm52CnpKbDFySwE/wuV4Y80HgDMAea0HtBvbbnWChtxasujXm36QeRIsZmwdrYFVmV4m
4uLWXDorsno6xdwjL1JZLUJ1qzAOg9uGPBVl1pGxNfAUVxHx56QndN8dK4p9mL8iUScecwXfTBUr
xA9sw36R1cB0CIu8sx3bXCQJkze9rGC0Si5MfS9sWN+nUPbt6Pwl/YY5PlW3ckL/LRkcag4A5rAe
+4xTMX3gZzO7+eHnCXi4fZKN/z6is8n82GYPUQ9OvoLfDpDyQm5QIjz22nX/Mx7EQreLxPRald5Z
CsmGkVvv2cGOvEMrutatwMwsmkyKqREbTr+Df7ApTaziodzL2NAd2s+iwG4nGGW5ADmS9wX2aR4Y
b0sA0oIY5GI9evLho0piGJTWlT5WRHQYvhXk1ClhejNzR/nSlU/zLpS0DPTKvcZOvbL8yBn/KOS0
JklYm2n+gkThQZGhlV8bs4sQbmibBxN+JLpxStEgRG6Lqyy0RNl3SXFfSD7tmSJsrRTR86/I0xTO
31anh5QWZxPnVxBJMlIiRoOoFlkerEyM9aMPs/tNBmXTKUPv5OdNTyCOFb29EGS0kVA7hvOYSKPn
JvO1cd1B+VCy4mJgJCFNp96ZxXyIOfDZepZx0ZtdzfcYLHMSNJJ5Se8Kwfrjuh9YekKqf+2oGZjN
ogVBZ0zGFuP4BWj40bTNYQIzsmO5UbY7pMpgjesXWEiWu0n37X2apq81ojYWiyqw8UGRwzuf05nQ
HWabp+91xZHiv7paydiNj6iB5d9fIHenatUK17yhYuTeIdhJaojnC3k8Wi0Wx6pYOu2DaDZwJXeF
j4LL3txdQ79iGPzZySGuAjkAaxBFShQV+ctP6Og5YyI2xTjZoPNS3PVGDJXX4ydi7SOAXQnGvStc
Kh8q5AupwjkjD+UsVPcyjysSHiJLcZYMOj1V16l/cBpzrr8jgtc2z2xg9ZyvEmugUWoyjgs53/bO
74tR9u5fNvhzIUHP2cGvJexmXNTPmp/koDZdnlutG09CktxyMR5/2SqVItVAgWlN6gcrutO2y8+r
IEG50kHuuIhGleBjsEKQh14Iu3mB3c4JMxjSVqQHHm9PMxXhGtMV5O+zX5OfK4svbO3ZD6/gfSwY
WWVkqgTVNYuebhddlQHjOCdNcU4q6KbIReUoUf1Ydz0Jm7XxmkRPv0ubs3XReWBzlWSfpALLPgTq
T9Re7RwrJYnamXsoS2bMbObzYdne2VG1fZtK9aPJQR88Ewl0iPU2s3EEUlntsR8gLU7hJguk4f+o
H5Onm9Ch7uhsFB3530ubXhIwa44qedVJmtzvgZP365vqnqY3TVWHPeM8rdUbUmnd0TP56knKxDZE
9Zx+wBhlPI5mB1DPHfB0ecooswZAq4cpoi5zdlaFm4/Y17YJ0t2jAs6AdJTvW49uguoTwk1PBx/f
HPBztCIkW8UqEPGRX/xx21/4ltMzq+DkvzRpfovVLtiFrl7blSunCtr6whSMOpgazLXcrXoMyuIS
jlMNwNGkTIQqbaXEw60TRz3w5tV++XpafdaUe83LJaeiUE5eoMyEVa/z+MNGPNf6H9o4g+DjDNCd
SPwg7PAKF9qi1rhNzTrCkNQKG2QmOpweVJg1B5c/sXp5tQS0XV/BvSaLEvGrHZMdn5qbSpxZDg8L
SK9bqJZicmqIxBZA+LvEKbOOWia1BIuPU7KMkyl/I9RxiN/2oNTi4PZiCVnezichRZIylOLHPSH4
3SOmjtaQRV7tBqoepmnXvDuCoi10U1WDEaxpPpQqPYfdBroTGKFgIDu55QJSk0z//gPbn/D+l1ol
8E3XbLt4yBKKsuiHCe7NU6r1tJv7r5Kz+JWul4aW0leZhhLxBVJeaOZOibd1lZuo8350PRUStQai
QAvNAPumMYD7bO7By5As7AmjgBc1tPACDx5PjuQyMhnhTqzNXtnSwmnrWGvA9u3ZoYbnsePz4uGv
v2UpiT/F4hAIB+Kf6TnO44PiHYSvISZurWHl4y1izYNbZ0tQVQKwNZhfYkorfac5mKkewSeHD2Wu
fNIZhR21sB+9Kh8IQvCru6Yy/zROzIcQKHoOlSO96ULJa01GpK/jTwv3A3Q1ctzoSC3ThIfXY0V/
5aw385EQW1TldMLvA/3cXTmeZP18ksSmOeFG10gmKaFeE6fe1IEOzFplbrJUpYNeL5cUhG4Bqlo/
G5dLMhMESJSQLeAfKFNPack/8OFratV6K9+4ru8JfH0mNfih6wvRdB60jFUOhpD05lv3CWG/4dIh
VXg/rGg8ZJaw12TxdKCKfuFWajH/LyEifaSF3YaexSTEJC8hq7w6NYbcCIOb0ETabXZLxWtRW7Q+
UT3jefiWi30D5KwKkj/zzOohfZ2KZlyD7veAiYCOooqxHWaDxLtLa8EWdyz8lH+BjY/+bEPEoW9W
3zXN99r3P/PEzLnC4evQFWrCpO+VQbhoEDBzpi8yNZcBrdihmqdfaJyjPHNwkkhHGYi6OO7sbFCt
r44+7WHwVlyj9q3mL9EiVsiSWxHemTKkbSZovCJCC2V10q8kvym1z+CHNUgsZoJFTdy7dWnGb4VK
lovSPoYPqkrz0lJpa1625+vAV5ygpwdeiDDWd1+zgn6qUiTAi5CTMshY1ceNtRuCn7YLvs0XnLff
GhvcbXMdLuV2CDjdufDs6hNDOzllLtdK0/DKdIVHDARFaM20g/tmPQKoC6uccVkZk9H2Se5gsxlG
uXEi9if17FEA2xWUX9/I898XNI8HL75WBE4nzo0sVOxcc2yN+4KeKe1gJwY/OLWHDwL2h8R1X35/
kCLSpqdT9qzgEoTdhg0yDAyGy2IE7Plu7SLI7LTaz0NkdEzz2pCQGeniAxKaGuXykMk9blPdMv3d
BeJZ4QZBcbTOsM9+eJ8U0vh5cNTo1aYN8Pd0ng8vb724tyyErqfc1wghLIsbY3xBYvmnOQrejnlD
LsORzMcFd3LwnKjQ3yyLLsQVpiz5UzjjyMllgoCmh0nEzn6mYJLhcpDDp2e11pZ/pDYG1MmCIFJG
+w6q1hSLyE3umK63LVFGIqidtZWAVdcXlDOL0HRlS9DUZHf4X40d9SuZvDIMY+ys4G1AcINWwRnf
i8IyJA6j7Uh8D+MQuC2Ms9AT/9E3lI/lNJHPBMNuQ0DsLtYrapwSsEZ++nJnFS94CvMd1KWqE+y6
w1714NThfPtDldOZ6bxB1LhHKI3tf7jTdZPYlLoGnO+gSy045ZX5of1rBcMgwFj8uf6W65OYUJht
Ozq0hkrl5goxpI7M7KKfOwA7wIciSrKnTMRsvhu6zUnIf6/llkQEOADCxML3ti722UnZEZyKSeHP
9vojEDcwfT8/YANSSbi/SCuVhJ2/QRk3hkdwzvZTUDf+RJ5bfBa4gSa8byTF3lYqr6TQacGmxcFi
LGJWhPhumkNkE7FNmMMr/BS+0hOc2GhZFbodgO4dIeB9YVaA/HoYl8ewe5G1gF/wKRm1aNai+En5
KtLqeudHszN6mOviyp8qxNaRsvJd5lvLrYWqMN6nU+COzbeTNZ3cuhYgPOE4JitijRLiuP2FD11W
28Ck+R5xN3n8vugTv50p2NN1pZxA6LGXEauQf01TNhh6j3h5n/5DXpMtBm97oY5qi0qR1sgOFm7i
tj3Q4a6LmtgKx0OIxxqOiX2GczrqcgY3GGieYB7NeZU87ri+5KxSkGssgQmnFOWa5JOha7WPimP9
BwBelnyR43Yip0b9QtJeYKEWrnjnC/b0hQlrra60ylHNE4W7MlGI45HiBN/Wr046cjjgytOqcbvS
5RxibzdbkGl3Mt5Ts2UNg5KjO3xqkJQPN++yiOARl+Ty6XiRWlKdUyzlt3w6seQnWj9fsm2MwBdB
TfwLB97FwlIw31bl1vkWgNT6jRf+mEZphA3fLWLOGQWkZ5T4kIfmU/8RapZjqoY0NY80mc9yGpFT
XjRUiNvGJzOk5XNTf62d9NC0WyKqwILZKdhk+1jxHMdpVJQD2a5WwKu5nG1/+sgW4DDLNk5iN6IR
9ERqIdCdFHJwxZBNodWu7YNJTPRN2sKu5zTjsees45q4+4c9CHRnpV3oE4FYzlLnvaT+ndklmDOT
wPX+kfOrzU/PNQConnmOkB2tcigXUwoSa7ZvpsA62X35tCeA0MFdLmptaN8O1GPX2G/v8cmwkEvR
cRoRIPdXpfDV3AZcour+DX7tsn2p+32s0IAlH6y/Sj03e+awAX8W7NLZ7zgQx97H9PTt7EwOMTYu
SpAix/nycUWlDzJC31y/KXmoaa7zEeywq+C/k6Ewo2ixH3XK9OnQ1LW/grv1Vp/k4+VRGHZCizeZ
Uin2Eon0/XBiE09VLyTvW21ELnGsTX/u4vU0nzYF+Iqk2vHx+IMc4gt6bDbeHm1YtTu0gRN+X1jU
aR1T+Zah30LtP57KgsrZ1CLLCDNLCmDSz5ozblG9lqrAm6LDiCP9JCF2G0Wpl6XZ44c48QbkJEEo
hVHUlZPhYDlehu5V0jIYlrXGhj8rbNu7KIekXFzVUUBYXwQSjLjSC8vY4wX+PzN3iVdurGy3HTT1
vB7v96B2EkE5Kno1LR3dywef/vHq6fDY6wN6XG0xTMvYT7F6D+HIyONvqSVC9OT+8utlR880c6Ud
vTAXEnFe2rcl7YcQ6GA5JnzA1xxl9b+QNGapyAcCRXZ6iXFZTMpsCBpfJNhK2DNIlh59bMQOqg+X
sKbtRUjT8Sdpc2xryS+K6WNcfl/L5EbKnm2FT/XwkN2RJcp2VF41+cSqx5ckSebZ/RhKM9Vleigx
aoq0WscmP2UVy2vpogGpuZVB69Z75QHmkRmwwjK/SaGUaVYm+v8ceGjb0dFbo7YIbtFQH0ND02Sb
o8ExgM+Rn4v6D1xE+e594c02KbtLNBIDwZSbfn4wypWEaWUK+8Nd7X5QzdVN3IJUhQ4aoN4z5lBF
SjQ0u6foyNKLBrKsdpZk9t4eYXq0K8wuA2ldxXBKVfab6bf0HuW+hz5f92rL8GkRxOdWO+7+LqBj
JtPeVLSrqa6vCzws1hriikPccF/2xXzyzndueEQ3vpf76T1hCj0zpHBcAxvcgORYObv1oOP7hxtm
GNE9BO//qk3avekephXIr22CBxArPuMN/ZfTVaAd2MdD9Tw7fz9miRo3Nrx2k/7GUIMk37JVL/tV
orfNJpcwtoH/8TebmdH+cflqp6MxuhGhqJRoiLgwQf3/UKcOlXFIV5GN53Z35ali/+UQieKvPumJ
0mgBjJIC2kDUPvI871m874W7iHkaxinwBV+xPhM4tQwcPdVEjsPanUneWporBCa4h/9fEY0AqZ0d
3AxdR1yLOp0uKXEvEGnkXHQpfA6UzsE1cuQi8Iv5OtIlL+Vx5iDiga0j5msmQBn+7vkWpfM9uAQh
JHb/VD5CM67P9bMtiIFNt6AJbmqUv+HJX2zBQcqsU+JVDEt4hJgdIARAxAojE8cS2iBAnrHJrW6Y
0mHndz/l1HUw2Dqu2HGzUblKvj0dA0gKjBz99v6HPIOCqVWxktdCeXWqPuHWOqULc3z3Jw19OJ7r
ENQFxj7Mjl9loNZgp4yRUcFlF3SalYcu4DWtX5Hz/REqQxFDnI/OTPGrKj9yx2WcXavT9qxMs0Aj
cNNImO4ZDKE97rtPulfg1gbq+DWIxG508JarBS6UhO6hEgHSHI7kGK7cnDZRQu0kXOo6VcKpm6vy
31ZnMMlvMmo9W4N14xO1LALxscoRpMvVwG7j406/SxgB0g7/Vh056ilPKdZALmX9PjyhmK7Ctogl
5xq/8ohlj1Yq8+lwKxidaryAEypRaCzyqqpr5v4xFd3Y2HSugJDmDHcZ/+8UWHFFT2iy8shsPYFJ
zguGS4O2Zr587wHED7WP4E1XbT1/y4SnGdGL1mkMkn9AVWGcAX0cLkK0IgjT2PwtoCuY6WYfTsVX
yvPmDGYYMfl7oS+q2AvMW4Gkq5tSI5b29xbBj9/yjDEF5pmJ5R07cSmOTAizm/mitxj4ZfxMUYg0
RCbQzOQS/Tq1whNFBDS8Z7nuxapm6D/4ZlxR9P9Fm2cm15xElpJT3GGPUyd0h1WI00ZSiLAmQxIZ
U6AAbGl2PpxiE48IHQYiO/XTnmSmxKLblBX037JWkfTaHo8Uc50asOYjoyT81w5qbpn/yu6fnmS1
FafK9KxPURZspeQ4kqs1BZv+TRUJmlpqqLd0iq/MPXDAgjBBUh2StBq3A/E9h6Hppx5JBPdP/L5l
//RupBAU62dDsOHF6y7KW7DXc0BcJ4yHCD1DkF9j/H7XXDC0dAo+WpvntPCFIOcgqS5q9x523VP5
swMEBP8NsTAO7j8F+xMJOyGQg/qbjqZ4sQc5clSNb9yrrD6ijF14789TjjpIxKWQ/ihU8ts/Yhe+
iPl85oz/zN1PhTpQSFAF/bNeHnnbAA+au5wcklHvw/5sL36cnDLKNbUmLzjiNH8K7jZXZW9SmjED
NtKqEcIn3tgQVJvbAwSHFAjTmW2wn1EqVeMGw/yBWk9CIcGtvOwMob0C1T2zmw/sed1X7s36nZGM
WMnl7MI7L4eHeSdxQfXB5e1XJHNIT3GR03yY0wC5srqSQXGLX9Pkz8DzbslbC6rBNCaJjKf2pqdU
gtYTHOSXoPDPjwL07t8hnHT+CijKz9I8wivVvssEOCZym4o9AgmeD82psL95Y6em1YiqCwxA6tDl
Ph26qi8DFfp6UNmAl5pHrWiE9xga1mdsFUJjDaucYaY6FUPmM0bVdVfaW1mtcSAX2OOsdc+N1yiN
bcXs3kv7K/CFlKMHGpa1r9gWqZEPsA92UaOmORTJG0hrJKGskplYf+YdwDhKZNdJW2x1M7WXup/y
j8ujy9CUWfsZJf5NJS3VgIvdR6suG8+FXVnPVmmcZlcNiTtaeOuQL7tElM7x4EoPxFTFseKvn1NL
cudLBxxj05NbGFutre1DAwdmScCRSGwEjTjKVergJnR6ByNZP088rC3NItYZnDn5DV8DQifwSCMW
9xjCZ2wXirkm429IV1xoJrINpV8n2Nvu3BQoieVuF7WJH32FdVrRkdL8jUqU6Z/3gDYRh4BYDKPd
b0CYCqYQD1GoBXaXGCK2+/CPZgK/m47wERs5T5ltBGSqKCEoi1KWFq/45rFzLDzofWa28ru230/k
o4NSB+DD4TuTStkNXlggESQjQQF6NzwoU0zUWc55a5viQIykPM8TOPVVIA3vJqxG/PVXsYtikXXu
56AI4AuxQ9bt5pr7PatDHpFxafkmJr70DlJVsw1DL1DSrvci0XH7p/65e+pHYHXXcHu6FXLL13xE
1UZXsgyfDqxTlKdWqO+tEwfzkks5sZOWs7xnFG75ObY45iVkV5HviqjdeBPiL81LA9V/YcQB944j
mqIcGlmNrp/OqMZdMPTHapPVKYvButiFh/RyAaKnClTJcD+2wR/f+22v9DuWY59zuihZAoKdcarh
AVoLAqGorRxo10K0U5PuvjCc4CndknhUq6DUSCMONCX6sbUMdaWHIkKuK++eajreO4nyOlBdibCP
GUbNzWa1DsX7J4ui1gtjhL9typN4bN74fDjVi6lxloewRtAC7DU5ySMN4+BrXEwDJHWDJMuTZHx0
vUMDDnqut0SQzpic15p8kKonF4DrXszGUZEkjF4Zv6zAcWNOuNjoWEkBym6+1znXN0a9EPBb9q/l
mKVCmerlsOzScaKlinj5+89NrrauNsdlByNYKK9mqnc48XJ34mrR/cshqiSHTeqodxp4f3I2HyAi
obVuCZ244ZGuc/9c8w3MMt8DlQeKyU5nYQ1KMJFEXp4mYx4qALklMkXwPemB9IJE+KiSXpq5o9jB
K5M7Jk/uTY9zDRA2mOsIFniC97hkCSEPDiPMrGCDGVbtdt8NaTOKI7XMf77n8hE7vPYbcCsYa14B
uuw98IiTC8PWoZsfhEF3tdfgiee6azBbcDxEtB6PDu9UV3zPq5bedQTq3RU9/T5aKXNky0rogaiu
clpCNf5MzGINHaH9Nonax5M42lkU2Lq6lLyn/tzbk+DtJH4TyX8SDVaW6ZDTQ2tu/ksfv2f0WU+R
BPeUXGw/Gqpc8HlJBY7S3JnMZIDkxEo/G3xZzWqNKoKxt6oobpi6Ev/cwB1sVWHg8o4ICoDA08Iy
3Y6Gvpwwr+0/0Yd693r1u+8ms8H8kLas2JFRfTUn1MtR2hzl8szFn3Z5rm+/K4zy9tRlvqwtJusW
IZBKE2pV+J2uH0J1wETSORxDvt788E5lrk/w9OJzSB+gbiSqR5b6P2oVtc8XOlD+6Spa30yCa7f8
PZh6V+hNZnH4swXUOpkQqFhVzLTLwa0afNTkXLlDQP2qpcA+i/mIWeoKd9rfK5Wj3uqqgDQ/jst2
4Ed51WKlb4QZPxWOqZb4j3Gmlzj54qFuFZfj0muUWwLIoRBrm4scvZxuh9q7kUzNy4vkDnwHfJGn
Biea3taHsge5gboCFwukZf3IQIVPjR/cfT9A5falMWh0OFIcSdeFXPzfHFNF4Gapp+jUQeV5XmPd
8aXvs8Yv2ZEYUvkBsxyVfAehBFAyUfw1sWYeS1dtZSdwQaXGez+yQlXQnATVSzsYs2vK1WWC5GNC
WoXrde4sLy5PaeGxhCP/3ZHikByZiDYDBjNvqYj6nmW7W28xga64WBrLWPmpKireBQsurgtL6zuO
Uiw=
`pragma protect end_protected
