// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hmklI1w2z0TCHfkQ7yMtj73H9zAslP3RjQLYqosW4M6WQ3nyOXUoMFaaddyd
FS+2CYs2bEafXqOEIo/FpRDCFiG4aYX8iqVoeTZVrk40njE9rojqRMEFbuxH
35V/wTvb/hPj9C5AFPYkauToHdu1JI9s8lcbmefZwWQMkosTSnAwzY/x1CN9
fo1vmx3ai0noK6OTdV6R8RBUqu48KP0ZRn1iftPWRYujmEVqEvVQMPuNpxvs
6UYtc/c0VFRwQd5J1G88jXTQLT3D+m5ItY/HWeC/7+amzLeDFXug7sJeFsAv
0vmOHSCntNTCRoJHjOtl2uQmKKGlvuYwKhHJF5Ee6w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JdFZ9nypFILbCXzdcC7kR0bgxzPSDFHcISOeRsU9lx8iwYbFeJCOXLsYQEvi
QdjkfHEkcD7qQ82LdF7LpN7IvD3+WBTZVsRBKDcnbCN3/4SLPjnzRrvV1azU
ZoxgvucbOkFDG+N9Urvfvu+MK2uu1nK5+YLrKYpJiO68wxZZ7Dnr16k61oCd
zaC/FlAu/48kF4RE9uv8ZzMYS46YmiOcgxW75Li+enoPUO1dTZmBWph9tQyp
XVLUz9/LgvPGAhSNTb/prtcUwq/QsI8ylnBbyWVHetx5jvh7hwmfjQfvpZbj
FAGKPxo+4qzjbHbzXZNik9BjWjotAb3dOcg4C2/OQA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lnA3ccK1KZN50g7QROTbycFqcsHy2i53nLSC1hdqPXttky6Qa2fwKW3C8CvU
SMoR1eAiwlbCT3Dt6YvSCtcHXyqrIrovPFnrJb8cciAm+fTwtZoH5VCnfnrs
Oovd7GFLQYU5xEv8Db4KbYXaw9qZoHEEKvnLwtBbDho7pDHJ8IjQ3whIhw7U
OBFkuqQcRpRCxU+kgGX0AolocTtea1HBH6BCQnWzqY74P/YoREEkBhr1AgM6
5fFFYjK7ClSgHKV5z6WDf9qj14JyIOi7/GOHfIFJYhaJ5F8KwMa+I+1xBpW3
C4LaXihm0YpWNc5QtinMa+rQfMvNfKnuh5ls+y57Kg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
j6S6uzpljmj1Pc6xn/3rGCeoi1UzX+FG7CL+863pujRGtmdnUahqZ2x0Dx5c
Vm5+Gixo0FCMV4M6Dl2bsFSUjl2cdsHl3F0GWgvi2RhznRXt4wfJr+uDsFQg
N63iXEG6phLa2istKlZD2P4NxjUDcgsP6tjTpmh10u9qzICiqms=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
AMt/YG9DDgGsunCxUfiM5upb6SakYMVBQYtBCQKJwlwXccwutYOkqB3ftCTR
VvBr3dLCH1ll9icUnIIOfCKUMfhdoAmG+KqxVI31WaaVQubvhqjT+KsazuRm
Tlq+sg1Opa7QTA9o/DSXV6pGP6thsT1sc9b/BbtjWkq5GIRGl7dwQUYm3N7f
Rd6FwiEtHU5Cg4zM0p5OreLcRg/jOxBFE9aOkIjAEXvdmSImbkTA5C9qI8bA
XOAuROEUBe7PiKinVNfQNlXnOeI4hxb5JUYMLC+6Wg0N0H+DapzoWvTDPsY0
ohaLZHy0RMv9HYi4x6w15mrfzgvIVaHcuJrNN3tq7lNrn3FwK/UrvpUKXFQZ
ZWyIdpqmoTZRCl6IKNlGU6TmSysvTWFBgh6jOzMep3CTEWkWh3MxDRcsdegB
dZ7lqLJH3YPLrvrk7fc9djbfZFDn28j+yW4aGVUV1qCH5Vro7z96p9rzu3ep
biV8og3aAZV7cuHuI3n/uqz68kQRaUil


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hJgjN6MwNdbSIRbmc+d+2vSG6wcVWq9/SEZ+Tzs2PcZFU5EpuLA0jPI87zTz
ETLszjmdc6pb3pLGB2/82/0UXekG7kNcM6PzxVQsTFls9d1xFHGhwAJbCzEy
vH3oq/4Tmi3uV2yeZdmiOVjXndjjkC5Pgb/jKJ55/yXKpPDVOMg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RMzhBbTawwHZvIdEZAvoOikz063e6sqbaQi5Tof6+B85xcPmI5dLrGidPkrj
bxXtKoEnEzyyrUuC96QfvEfyd7GRh5svp83Jgq3+DCenuHK+Q8/yuFODcBxV
8BDoU/8zUYGzhEfVzouJxrV9f9B+tdWrWi7/rq57P8bucLpPKIg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1264)
`pragma protect data_block
vrYAD/8lUJa4KUvz2DP3QLdidMMmA2wJRZF0Rgs6gs1KZ+X/ixHYKhXAi1Uk
/koz4bmd78sEC7yRAcxFuylcV4GPvlHwqqG496ZUxqyqsIp8XJqmMY1SlIFP
s8Mt08/Ed9t9/WYhie3JCXv5u4SO2cD31ZewzQ7xmSyUXmmDHzG5UXk5hT2q
uK2nce3uhNBQrP0sXDHY6JO8BTFBQ82FHfYAqoPs0/JqH0VTxX4LbFynitbb
MgWyP1/0rED+vxqTbDNIlIkhjgw2eoNeyLtzAJ2FVLs/wXjqWprpU8v1ngzp
Ty4j6qN+NyawApJcBouhfpSKGQqm8yuNkY/K+YU88kIjPjQ5aMSy3NTEfwip
iqJr9uH8fWyltN5xTdciVJZ5J1czvaSkB339bTgCSDD/uF01CRQ5r+Fb0W5f
eR7rK71bazuJGXjdBNii3m+89fJYOrRZ1QEsXIrz++8FGO3NB0NMqmCOun1l
F2yy4ioJE55jK30FbtxVpFGTwGwWq1d4nrLL2ydbzhZp2ar8s87MO/5mv0nn
peQ313IQ/ckf8CaAVpynT5zzi0PbUu4q6orO4veJz9AA44kaa24dXxPyprr9
bP/OUbFE6erLxugChNK13WGUUYEdrGggbi9zVLFA/QedffuE9o8Y1g0ZiGKX
Y3WyFl984K3E7JUBGa50dvRVtwyws/nzUe/vIQABp4gj+0D/5jGFbWQ+7vJY
6xZxMfj2V1tFiwJDmXx2ieRPLzr+FR/1L11JXcr8bIigqR2wjeMA9wF6RQMf
maLTo6UbOt+AFXPvM81Ko12sWMtHM9acyuHQRC4JjqewwAiZhP8cQjBYIRD+
qYGcqotvSIJRPwGEjGhFUdEHcR7WczIyvpzRBRUncf9p56UOjkOOfvUw+aZn
LUuOGU2in3TMw3Nu4vkn0zCY6WZ9o/RV4JSzpxf6wcQ+19IQ9Hfc0cNJE1gr
u17hANW+vsn20zMYDMjQybeSVTGyIgeYoffggxAp6c4qBf/wgwj2v7MVm/OZ
s4J2BgjqQFGaRUDLUCylwBw50SxHgCNRqZv01qkFZqaHH+5xaJ+MM/+/FuF+
nVzVLCGwgNH+ii5HYbJu0kn5AR4X3Dd8XD+/A+6SQvZq/A6QDSFfrLbaEehr
CjERUDbaDYNDYqbpPKLfsSw/Zx5mz+RCeHoHZuAkJS32OAYg2MRMLdVtbCtI
NdjE8DSXibvEz72v7j07UDinXfkDQjyKI1p2ldSDmZmyG3S49Nw6vYqG6+iz
Iq026ordDqclSO5VZtJZoiVZUdM2nH5tXUf6fUG9UMm2V5HHw5giK11YE+e9
++rVz6vfjqNRScAZhL11fkN1R8wi1RgppTtVpA2EIkMaHjeAOJDJxDHGcIP3
KEt8mrWyNel+cF+EbZ/CUGGVaRi5CNP/FJRXoq1BlkzFZJb6NPJY57/tU/Ro
0K40G2i/T8kubbzj3Z01qOCAICVVJVAChK8MX+8lgr/iwnkk5WKCxj4TXVvR
WmjSvVt8gfakWbVG7sFAV1c0sqPt12MuO+JfTvac3JfjMbA6bxxP6Jqzq4xD
TY+lG+PYerj4g3m3FJlTPR4aYeqmW1OgN5tgFBCI/7vZ5XfSU9JuhhENdIww
88XYIFDE6m5GywhGO2eQSaWW5fAeX2OLwCPHDmSOvB2xIZz5EXJVGw+dy5O9
A/Gxxg==

`pragma protect end_protected
