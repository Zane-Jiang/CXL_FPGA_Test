// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EkDgazufSNtrOR7zoqlH1UK4A0gY/lf6TqcsTIY88acD4WES1nc6lQqiD8I+
avOCF/EJAlvqBjEgcGDEEtvmSedPLWElknmFhT619JKW3UpjbLgDjjfZkC9P
ucCeiW+FcnJ/Y6BSRfp6pklpzk6ikJW2iXqe7lvpEcyotIEww2xB7wLnKVCP
PepDZCicmzJ/6cVBhP+apYqfWhhOgpUCHU3vBe53kr5z44HkBUiMpEmgidco
eFY/sxivnp2w8ipl3H56f9wbEfGEobTlcC7koxn+x8M72KT72tcMiJcCawEx
63vLw8FqopKgxeuIkYxnVq27W3NQo9TGKXyvqVaDhw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pdqne31cYz1nOR3MCDaLd7rEShASOZK+3C3sy3YpUJXgCyk37ouVMBfNFkyZ
xGTddey8F56vOtEn0BtvhZHY0UGjt8VGuVA7Jdz35eV/cFWZ0HeLt/WgMsxW
1R7enoOUaVbvbJpesSkrJACV3GYJEtAw15B+M+VJ0Q83qIkCDRbEndBERvwz
KxTTZMw2Z2u2VKDMPg5ppUeMC56aznMTTAOnCJ5oBI1TnMDoKrqTVsuWv7o/
yB6K1GHMbfqKt9WpVid1d6IRJtd8AmktYkcf1fa2PT3nyIeus2u45K/8Nq5A
mhMPp/KtraeGBL8ajwY+ZNyiAdSrWl/HFA0ykcl/lA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J+DAfIewX1Vm0lXtWj5uvmziZXsZZbgv6tILiDTO8Gk7A9mHYLPej9qWfbqL
+JwB+I/x1Vt7aZxd3MuWhf15UixPQudGkyBouK80EXupf2LXct620CF8Nbxj
ZKCJNcpTkR2eKleHS6Qt5/CSI2aw3InxpB6dsRmPb4QjXszyvqz4iwqD16TL
UU80Nnd93mgG82qG6TSnXviM89HLZ/JS3Zu3cBebdSdNX5neg40GpLBQ8Mbp
KJvTDOTVr0snpmkIieWIN1yHu6Ckjt3lTJkXfpk85N7af1Sm5/Uoi+MSAqsW
J5UhiIS2qCqYjSYGin8VmfQuPaYDUBqaPpyb8fQJ8w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WM/csh+gGOlH1jPUFNfBe6xG1q0KhhMZv+6oWA4qKn3HWuHAM9BJO4aBPFdd
FxikZSB4SNjm2+nBbndwoCotwl5fdNTxZMObd6e/Tzvv4VcizNsiOEdoAJ+2
fFtIhyD4WapKxC94fplq4q8d/EjGaBACSCHGrXCuIKuHA203Cjs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
f7KnDaK7IZyCpCm3alfqZlOCEX/9PfPLvregz+nxyOotD+LJEYv6NikCUGPO
T0wt94vnVumTvkT54DOrpQb4gRvSvN6qGIapRWd73DdaSfaT8gnL+Dy5vQxf
vb3DmTabMmQjcXzRA3bLnT42wux/lzhDSPMgs3T3FHAWszog4h4URY8VtSYk
iRd1o8gjWwKPs9HxOvtBzSK6KcNS9+ABEP0LyOeFE7oYXEmH1fPLGxBooq9Y
TWMpnqQaCzI26eKnICfRCDLRKWjvtF9TWL1faLpOuMjJxbIxvg/eoPfGY0P0
2hBdXIs+1m4Kg1H4zYvD3gXDsJfvpZ4IGVOv5/osLrT4c5/F1c9KK6lgOAvv
oiLxdPrVk+rVS6u49nFWg1cXs9n9mCHy1Qxmap6cwWvAm3byYUovlDqHzctY
gixC+HSdaEtRd4hjGgi2cPSpHqegV6aTtyL7y6V1J67IAkjjyp3Bg/rIzGj3
/qUql9lVV7ccAmDYAQ8Pq3vvXM/JEBSk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cU8n1/K8Y6ApoGDCrWC+P6naJJh1BgYFaR8uVVbfezRRxzdBCqBwcByY5Djd
qz1Ni+8QylFSOR/22sVAU06l34GUJjPRcEomi5auq5aeljsAU2cndfeusn/B
0lNpYN+sn7uhxOhW2vMOd9ECx5G0rETp1dlAQHhUx+89ou1tmbQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ri3voukTLyZfa31OMe2IabYp8mHOaMOM2xt+tmCMPZg4aivRnu1fPsl4J4wK
zrDBTrS8Iy1wsn9na6tjEmEgwrUeiKTS8LHr9Yj4MeiZehjPqXyArBbT/N1Z
AfVnbXHz/HUICzkA1Ke8Yxg0JaNiuHzFhZBrUvWJ27nOPXiFgjI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13040)
`pragma protect data_block
Pq3iJPskNPlQC9ZwN2JO28zcd395JdnYsiF0MPaqIXOb3+f45nr85nfkYzCN
RjnT4p0ppcs66ABDjhn9yVkfOtSrKX9GpX/sA0QwkAxolmhyuJhH1huejr2m
HCwitDzXAVqlzzI7SQhnBA3cVLFvM/Li/4OaKVc+8y1A5WPXyCHnteio+hUs
TrDl2tXGxMpeCrd0xD7n10tq64Hzgap3ik539RaMXDIm3z7K/hQc5VXirnCo
LNwTSVH/iOy2Y8PlWLwDpq04/toHo+iOIHKrGuE+JyWnBrDSwGc/0/yoTJxu
OSGkTATHzq4i/5Drq7Ajllda33qu51oM5bZzyryWDeMmJBOrLCVHXqD3bgrz
GgjD9nGLYkaD+TVcgXj2H33ABazG5F6d+1y0lSDUv5fEQWf9kF298qYARezR
nqmI/g5n5vuxPvLtSSMtG7zGm7NwF3Fi7zcuLmJdTbgMl0K4EcbPVWQEO/PU
0efaC/RmoiZ5+jG2t63INcyRxftYGladu/tyRh+L9sXTyypUYy/VZa7Xesev
7NwM8kW/xQdTBQdeixKHcFpq9xWVsMsqpTgEKCq3q8YGoKCNBCiGGDe2FOYA
bLQL+izq+AO+3ZxSxlNOSzqxG1zWxNFQwwgRKqdKhqbeT6JsU9zoprwkDmgV
3FunW6pYrj3/v8wfDY1NBwMkQISwJq6v/RXxOLjZTFa+A3rzzU3DPG/N7SM3
8D0c36gDAdLN62/KH2ZhM7nF9lLa7xunUdBN82UYzQJGKCWzWLPGX2WdddHa
Dykk2IAD/TrE4sPeUbbWM1f1HbNwDwPzR1t8zJuYH7UJDMBV32J2uEirDssz
BK/JRJ72OJxCX+dEv13O3c+Y8AM9Yh8wKJ3mdBm63hfo1iagOcYUwxWEeK1A
P8X/MMVWB3NyVnIqW5yMRhom5JY+de3OE/IK1JxEJd4nO2g9Sp96vlvdmHqe
RH9ZwgCh+UpI/udBIfRSoFBMuCoMSWLZ4ePtaxfcCNnjOarUzoxS3InXrPOO
8VJJ7E90/Bf95kM0Mikqkt7xyvP/TecL1Acjs4gttjAGLf/4sJUTcaphrnhi
TlwmBGDdUgebwKdr5yc1whcUkbO4DVxlH+QBVkvnwr83ZCyH+QUEccjUgLfM
nePYUtSMLxMVFfXjGjSJRynr481x2RO38NbaXNpPAcb65EjMsVaFcjjQCNW2
Aosx0d6IdQfUyVbqw19jwEDjP5GoQIKiNpNZ7uMGrGMsmoz49e+uHUVJ2DL5
XwLOMudgJp9WdnlVYpFsubvbfEfSAKLj+YdgcK80GSrGSwH1IJkAccmfeUtA
LvnwxUVFo/xdPrJ1HN7VJnOwZLiAq2NUCUZsAqsLmF1rrOO/Cg/XozNaN+pv
f/YrGCEGmnIcVVOAwM1QoKqSOcSPCcssMgJ+oQRgTooVLSQ+nnajOeKfDP9i
l24cwNjcuPt7fd0DP0Qnmbn8E3AzDYmjSZlyPqgpX6vUFWrGYf8yG0vzFmOB
n0JMYs9ZbbI+laqSPv4K3YzljS1uT1rLrEMM38yz4qgKoN0DLikBTnwtzDcM
qAz7aBgD1LQ3VaT1uzGocrjtNmFuY+MUiTLWdE5r/F6ekIDMQH9hduexD6da
k2DLyUChMxdFN4tXcV0nmsgWkZtd8bJYuQvS1Ynh42vnd2Yl239Hpjm/X8Ci
hMynPLUGj0vYayuMzFp1yUq4Y4OvjqARr+fm90J4MdOgFl8sk5izAArVKxH3
iZte/Cn2JsoH/nuRS5ROHuQYQKJeno3ZnqwqRUtFqCX3wY0XMCSDR+Ic+AUn
4sW7aX1FnM0MllL3k0izX9THRLBIa3ZS3PJUDkbcR9E/pu742B0dXhkKKD/c
IaBJY98vv64QErKwZ3nSLgenori1dC1bGk7+VC/oi/7X51WNs+d1s6b6GYmt
tUxx/BFO6mqi0InY45iSS0CPA4Bn7wUFoEWCPwU+F6cnpCHqU2vNoVoQWUcr
dhTnAGh2tWgbrdIADmxFsVsmaFYvmcU0AWyDZQsDdiGdsxlIeEtu2xETlOIQ
9hN4Uv1KNVnFo+EQ/ePriBu/QeQ4HNSxFL0F6ocOTtsJSkgLa1DuVeE8ukLn
fDI/F6dMIH2ZQ4xKNpH+V2eAW7L7us9ZmE9WliVgzwcE23MCE4/nmBnpyrAW
81CGwgKgB+q1McrB8ctC/dl5FTTgCSj4UxY8v6wK6FRz+XNLBmZlYALdeVOt
zyQtf1zLERBzmOZxOh9AkpMDQ1unNEYWZY3q0WC2aSKEOfvXuIBQLobIHhJ1
IVCTmrStcBQUYRkLwJRg14U9BJbIDRDodNyCotLb8c0gVKkz6rKfLGhNa2Br
0j4wlU24IZXXa6+20Df0wMHsp3bMjw2Fk8TkZXMMNIGQj4Ductl1rPm6E8KS
W7+lOZCF4FdNI15pVyCrZRrbMeAyKdZUkr47fmHPhgwNXctAPatHNIXhPr9m
BXyzPyFLXx0aAHJK4Cdj5rKYdbRT7m4kuggK/6ixms5GJJc8hDA6R7BuEAmH
7GujVo30p55AP8qAMsJyN6Ja0bkYsgZg+9ps6nE0slgx9cOjppATUvXb5CsH
F+buV+pyTvPHCTr2XCbvzc7kE2XjC13RaUMdTcfXGsm915sHdbvWd9e9Foe6
/lrbrShODTG9Pu7tDu1wpJr9NR7y1/O5z6lO5GX5s8iMXxuq0M/I2C+8LErH
9Y8x+Ww/ijNu3CSEF5yE6s0ckcEs9e7OfXMaUSagPAmUJhePpF+YlTw0M4GK
khLv9hMU0bk838k0o3eWjlicvHYBEz0U2KT66Uh70QAAcdA4KSZKjJiMgvOZ
coQxvyKx6wTysuYNDwM4S12GRu/6sPVZU/z37Rmggd1wizfgISG6xOcEUW2/
oSp/uSvtMCjeMTeBb7cweyCJpWN7Qs29AVOYT9r+cYqRfyfr72w1gS2tM3lj
PxB7uQnT+6b0mv1ViJYYQahrg4eQisZtaNKQpLqDcxD2W9WGx5vVgWEcqIJJ
11sSursT3S1OOxyXDa2LjBUhhuvBG/WQb0aKBCMifAeLAwSg4mh9YnhQNs9L
qYDOhQtKhwT4d2ITvbKYTkdnm5KGI+yZQ6LuePkvvWUgiG1bWsz88+m4EqxI
aYJQkm+ggg3ABfEHd2wXIPC+a0hiMeGr2maUnk2loOwQ9rhxhyG48ZW9XNRg
hq7PJpSPLw+rANRgYbBaddRQBly8SiS+zxlpsjoWVXYEQ3Jqv32vIaAMYROC
drmmx18801Rs+ONJ1wA6eXympReDGRxTVk0iWUMqivu8HR+9tO7wlioXpvMx
z+BLCJpWT10AqSVCMJTfVU7utEaGQn42l57fbQYSvmjzZ2d2yccLW8rdsYFg
E5BFNhEuqcnvMuqPLdRd/GQf/sSZ94Njs791ZCICGfiyiTKkT2G6UMvxmj9c
oOHTWNm0SL8dPz/G+eytWreh2kRkQ6+V75BaZoT1ozLEXzpI2Duea3Nmq7Ic
8L61bNf+vGf4MSHYXcLet4xSC9VxyTpjIYxsmwoOX9dKChmgo2cKLDQKE4Sc
QagVmzRYrfx3+GQaOSdxDAKwCZQHADBxpdO7rGRR8Qo6AGvVrJ8Az4ws+dMQ
Io0zf1Y+JAoo9ALWa9UaZNQeUtvH6WGZlcwq1x9mi2PQvOl3NhWxqHaKcWVh
9KkqJmiyYR8GNnf6l1kR4jMZ9XgZIOxtUJ+e7qg0lhSCxvnFnnUyMXKbfPcS
JA2KvjDmngh8HJ8Y0PjP+r34RAb0Z53zkzs1wBsy5PwahZUDUjviX8wX8eoW
++ipwhP+ZECB5hhUcwd9OxHtECqS8YMGlvK1RqBe5rJZ9DRPp3ZLvM8eIXFv
sGaCll7LLZZKaQpevo7YfEpg0bCjyXzQBT3wRzPmIMHeB+66IVbL4VFAddSB
n9gZmkN+9BFsImSTiNKV84Bg3D+b8L84BKo3lEJtuCvsDyfKaIoeYeJ+4MRB
wqqKRDVXeX3vMRokiPYheMIZ+RNY21CCRDX08hchwd7UciMvA2NWBcaMZDaH
fTUTWs1PiABlFTUY+Zcm+IdGrPyQFLSNrZhcWz7HuF6lLZPbejDGEA3Hbh2V
K0wRIlcAPQm/h+MWdQGU8autKbaWeHd3psxWLdCdtYwKax8knRFpth5h1uB+
6BtvD+Uv6SSCuKXLnrjSBaG3k1Swi0fGmbrtT3wUgS5CLBh8ccRPnhHLPGyu
pz6zUa9B/S+nILsYVneoy1ovysQYQEejb8y5TFKJlX2sc+ZiARc8V5heKlb6
+0tPrQ3rkzvLYIb+ZeJnr3P9h8eZFhPx4sGofE0caKbIdAkaTfedpAD5+34L
RUUmsD2gZU1qHU4JW3Sn7kdnpPmV0RvSWwvFqaf4nmO+SnTaqK6vlxhYaXU5
SH+Te3l5bkcCG4OzCCMz2AdWqHMJxAnf8rG1trXs2SgLXBFAraqr3F/Aicw0
YONSbAFq7jJHl7ClcdjTgPvSW3WdxJOuDmvJRqz+jGRWME6e4WY/qCRtOdGp
JVxqoGSHCGVJY9wsQLJVNZenWLrgWUH8dRY7ilPNylF4YczGiAUVNAp+gz8/
uKWkHalBQ9jem0wkDmtQu8uyUFjFmyFQeNltoNwe0jKSWSDXQuEv1ElUeNTU
XvMk8z3OSffO8zbM+Q2smJv7Wp3FWonW8G4gm59bgTbwmp4R2PUbZYWzST14
49YWj+6KWDJrplrhHD1EJnItmOb0gAUphsRuF4pdQ7m/OUBqRD4P6gTBLjk+
hbXCdcq4LTQU/PLRZQY7WIijWd4j3F04PdUD9ebcrjs9jfVGNT8MABmn3gPi
Cr/4K/rWXIDE5qJxDMAN5BJtJL2y4Hl31URIdcdCZEK4ANHiJKObcx7nqjH4
cLQrNAwaoilDvqC0lg3+Z76At+5Dx3u85S6x7vr42AkUdK+ZQ3dn5bDAyb3/
XasQiEAG/YM26No3wyP32NuLAB7oBT68OtgnU+RybLyLwnftnAtZ8Hhb8Bae
eCWD7F0BpMRU2O51RhbqOwR7MbtvXwNMYYZzAy996xC64XUpC2NYB51MghA/
9qHGwnBH8geRD5oShPJQCnO8KeZhIXWU/bEYoiRnXbb/qwLoBaCMZ56MXZI7
DX+cH+seIZncxOneatI8XCjwd8qJJh3Vz7C3GethBY4JmckIrf+w25Rgal7I
vwXCqX58OVXR6KLWK2NhsG8l2O/U9d/t/d05E6pwwM4Eyt2pK6oK7LXijufj
hE8YxJS+6VO4dLQwp+oF72+XTJ0UHwinotZj8FgAPbsrVNJk4LkoojqmikUn
lkFYMU+p0I2JZjU5VWHIvzq19RnwrVnnWYgunfuEjzIkkyO25ntiAP+Q4B4f
aEpJcz7VTsduXNb8M6gXI2ZCJUrWsNnMwPsDNUyGTWVjoqXMbrn5cZRXyR1R
qcdyK33TzQxw305XCaFwZPUg3IY02HehjjiS6V34orvGuKPqXWF+pM7YPbDV
T4zIdcjrWn9qX2GT1FYbXohu/EvciV9vRahvSiOi/hTaxruxS8FFPyPkLEAN
FYjIEVwW5K9YeH3V4xIkzDPZub2Xo9QZeglqWfBIgnFR36NkVkvctTYgh4VI
2PUqzChjhtVAJiI42vVq59BAXoRtZZGdeVQrqVClaeaIF2lXKKub1F09BXIa
Gc78TWWIOP7itE8gDJT16wmvCc3iVYSOTMpfsSMfMX9sxdAZDeymBCKzmAEH
jWQXSaVb8FR1TaSDEwO8T1fvMHJ36cIizIDMhROTNbdKQvqN/Z9zucN/78Vw
dsW5UjgNOfs2TB1fAvqlsePpDjf/00SJRMttbqNxqnCVIezMywWHif+flU7c
AhPE/jwcKpE2Dkjlk7e6Kfdx7kCZKku4QvOvmVAWbqvY0hJ3Nbc7zqXRoeUE
/gkdsQbzja9W3z7oHa1DolHlAUnUMf40BpAuexjvdcdHZs8dm2zjIcymgh0d
lJgTQWeNvgY4Bq9vORiqU4fQI4RGrKOSBPBpuHdRBbxBjdMmzozDB5B4kBrI
r7HaTJ8qCjoJqfjK0xs767TEyLmrJcgSpTBJ2XfrZM6Zpv4cbmu+EJPvm5j4
fa6aERQSB4ay65wLpStb8k5MOfo6+P4u6iuFM3dBEOHagHYdxQ1vfAdV9h0z
GTppBqjk0CRalGcIVxCAWeA6XcO0F2JtwVx37NVhkGAX8FTXrMg2KH/Gh+0p
gVzA8ZUYrlAAci6WEeFFG2H3Fzuc7/D6k/vwroIxh92Gwui5sXoBRJwpc8ST
n1Sr1QnJSK4OxQxcCThfoaVtPqBsf/KGAindbDDOmInAa2EozPtHli73hw0A
2gKbyvW1MZElkm0IB5k311XqrINi45I9MnHD19XYlgulEAnDOQ5iHlsF9iS/
BkeVIPSVbjwfXqdcGrjFzFH9f5eMlPgpS/ZEYogHIptAwrYqeSAsylrNGBpV
2hxZyx5nyc0nEZVqjLsTnU1csMM5AJmnlGBsTFlpd+JPApuRIRdeEkBeBle4
1Gwcwof2cpRSiQoID5sTggJwm7/UBEMCTetW3Op5rKtXgmK7CvkBtNcOeMu/
qe+gpOkJyK/Xrmxu/kw8KdeL/H1f9xJFtjEucemRuqxQWszsFaG4BswL2bgY
KpLWBtxbahs4Xdwh//xe89Mtx7FBfa1yonTmJeKbD7FtwaVdYCX1JiJYBZgw
d8k6zYKeEuUK1/H5IS7ZVDxQ2JN9l7pV4qCTxUIfIdqvOIM0vqxtgDPDoe96
khZ3abpEQQJs1D4fpjQx8v5ueppfcHgzmb+FCXbduHyD0fTQ08aS67OuWGgJ
tK0N4E+tIo5L2BhNGgbRk5rKggTMIZhggrhlzehrnf2dm2sTFZiM/MqutwEY
i7zlD43rfBn4uPh0J58+3YxFLmiQT+R9AilNSjHDptaEn2PCXLewHNVK3o2v
XaNwDF4i6pCIgd+cXNM6eg7NidlAuuGaHRRp4uifRvUBD4IpufIHf3aDL+u3
GquUizHSnP9IFptosFXc72mlq46A3pvuCdKkr84awPWhsw1pwBGp79xYGZoy
66Ppnd2ezLq3xCEuDwxSSQ+eybF3EBWTJncttfUrjhIcAczZi99r9l/eErZ/
bFHFkk/wtJk+JlA63fVZWCtUPHvbAKpykCdstXJV1usRna/Qx02jbUrrvvF3
EWEl5Wb1cGJeoGfzePt2C0JCNNGaTAB89t1RPDK5YhI1BJ3wq4P07H3jC/tO
xLNQNyR/tjLKg9/drsdLx415UjCyHFVSo9l4FRO6XtPs54XXKXwPggIoGSDZ
6+3ErxfenT5CoFoDuBnbu7O/suF8UC2vvyEZ77hPSCGmPMaCbpmCy98EAVSw
089f4TJoagkGdF2lPdjjFXPb+m78krEk2iaU6jHhCmfurAeCoh8xkZaB6fXJ
/y6L0g/uGn4cnLx/rxP/0NgDoCUcBhD4iRHiDsfVazDqXB9A7QyVl8u1VZS2
l1+Yo+KWEaHkBmtpIY3SX+nhY8qzQtisnkfDwQK0vCZN2FCoTQGg09cTPf2y
W7uf5eseqD2HA7EGmvg2xHhToEfhoRxJci6h1OxaapcQd232ou/SrVX0gtmR
BEGe2qzoFO2eV1tihiFY29CipN+Qq0xzPpLGdMtSySOXoA1arCH06ec+5dGz
eGM9XWEypsU3jsaTgCZeBSZK1cAqCyoeHzaqlD4ygYpeYk4WqJjjwFPV9byl
Wfe39Q6jVfZnvad8ggNtJy8MYJcRUlMdqXMzKpZeVYgWJ5KIXlrSfUsFKXqi
BMO9fw13PRXBPV7b9QjBQ3+2No+VnWU5SqwAhYc7gwoa9p1HGsiBw6I4BzWb
DrNUuxZ0WrOYRcurGClLmT1hhnrJxwtdbrwaib2tRfCGSqCNT399A49h2COt
oue9un1vfaGU14h6ineRAMnaED2DAd5A/5hj36riH5FmDJN12LNpSyIfODMj
42HdHn5cDjewymAmnwhxoXGkI9VdVP+NYsfICCkluRCodUwBsNswGLcn67mk
QGGYqsm9M1iUvujO3TMfs/vZ5D+vAyf0QHAUwgcy/RU9SdpmvV9K7m6OpMM0
5/6wfV3dXc9tpWjDsHmKCAUYVC36dI905V/rJqkdcTrbMCni+fVAcMuvVrSL
RBqhFp8L4LOxugAdyBZH50Hf5GB/7bIzf4yaNfq2AGO/LL0Qy7HaSFYuqWG4
t0x71tGdPFqznIbVcXRLLlBnO1GzG7kd0pUQkKYjdaAo8me9QCPe5dBXNlmD
eSzYRZ8b3/+zPKcuJW5K4C2I8tZX/I/LRg9HKIEWvUb36TjRsOK0C8p8FZTz
b5akWFJxIJUriUuYi0jX94GTs3l/uB4OAhNv+h+skyNhwFKpHsfdTzQxaXNT
T6rCJE4imk74VLiEs37AOBFYDSvHeB0jS1ZR6Jf8pP/9wdwd7IzMfqUyTEPQ
GoP2KMLpNHfz9OS9FEUcPIAytHj77Rr80Xl6Tvyk/PDdWz7+e0ZNLgXSleWg
AuzVyAialLlVhKXyvNg/fM6dZ5wscihoWlqcFHGS7GWenlrPCNmhkY0XbhXP
ws1nDL5qjzi2BcfGlKcpIP7jy2A2DwsEfG30PQVmwbM5lF3fm3BtHXLYGPVD
m+iDhP1Xp67xyXuM751JQgohb4UWff0VnaEr6xvpnJxWC2g4kvrG2fVjxcoK
k4X4oiMw25RXKknhmVrW04uZeD9prK+HHrOpXJJwgRjAD73KlreS1tzA/lKi
Ba/adVlPUpysFZF2Rsmp+qnqS0kUYxIs2/ae+DlZ/9bf5gIZ6l9z7rKMaLg1
PZcTo5t1e5VyvglL78MGF/u+ALswsUxRx8bBOL2Z9nbq/03At75f5OWR1JS2
hsIpjsEJBBtjA1ezij8EGi7YSRgHWCayUzDgJmDOkMyVjlesD7acIt8YeY6d
GU9kwReijf/ZfQmRBiCPZ/QiJ3wyCmlP6fEKlzzhbzscjJfqHpJhR7dd4h1D
s4lnRi0U8zT9d6qeqgnzg3DUc55wGGj1rZDZCRdlNnGqmY9A+Pi8VzLOeYSx
oqTm62WR89iB7BOcTbPmRd7mOv9og9K+SLIwQ+YYdGk/BLz5v9ZUpSmxjiTF
EH/j0I373P+l9GeVIJ7FGas4crW0I0WNDHPyTHjJb94Fm436YFODkGz87zG+
YwmtA1PeRCs3UWHI8IN6mpEYkyLrnaYxuvCjhdaYlP0H6o50RgruiH5Dsu1j
kO21chz1PzDotGirsg8u2i/Ykg560TzjNDvdXSEs3IYUA7+bFjX3I2/2q4lq
q8+Daz0kvT7PjE4KSsDZ8OItvOBrYHilt5m4xk1t6ulxH6Fzfro9GfVU1CLg
YCips/9LjJvs0Xlrkyh6Uwz//UBIbnqS1YIcxsh08apR01kSGaJryuv5WKAc
7/FX8kICDMe1/Ki78UNKtIVl6Yb/dSARlCB/Pps5HkGa0UmOCU5nVZ3EWgE5
JWGf+d2AKcrr+xd2KXw35e4Ne6ZoJZUE2t9fGq5rs4X3PGCgDgXuiDpj8Qvx
fAx674pDhFhJfr9R1lhjzzV+uyoNUdbpQBQjaezHEvweyU0SFzmTjNI/OE6U
+PaQGMkYVO2IF7ZXwHEFb5ahdzahXqBtJUWevqS/RDCNw87tIy4N+LTY++y1
KObVxwtgXITjhAfmeP+8w8Neu93YS3ClMH4sET1XVGSK3ETfG8jjL3XgvT4q
DB4OX5Ca1KdX3S+uYOIkMGAQJcNiFF/a4ReEM9F68bJZwquo6gzCcu7HFFIQ
G1KFxmeGpH32eDVhljVHFndyX0KRkSn6tAsY1M+wqe1gkJLVA7umro5rlVlT
vCRMFUXovUuT76xMca/eFihtkqVtUwy8qx7kOKMCmorhJFv9DYK7GFmTEOgc
X/PjPLR6w89eAN9JB3pYlPEMr6alPXmLLsXcjdVXcL6rxNVmRt3bi+dwbBQm
BAAJVDgHQJTodavF33JOwS9vBg1Pan+p71Xof9dhYHmjT93ZC//Lr3XRmqXr
C972vpUV/FTeztorf1PeCfUXlXjPmF7CV7pRS8chgp/2CddsdyF3UdNSi9ep
VArp/XCxvOj14eM9hKhsAI6HjmFeVQn6jDVPoaeTEHSOa9BYGBdFxguEOEXA
c4Hliz+sFwhM49OXuat4TOZ95rwapvtSsxcloUOQ9TURKPBw38raAHp827HB
gZC+P5ZdNbCj8n4bnWrgczpTE2R3w+xfQiPlBJQapPeUMHLsXanhEVYCIpv3
Hg9uGJn/XOCIpaQKU/RzNX0JnqbEe8fagmQXXdg70q6BCm4ZcvQXyDsm5KSr
/5/lg77s8VU91uXHfXZJ+5no7axT6lxGmtdV561h0BCb4SfRb8ViQLf52yCM
L8zqEI0b1e+8BhJavUFl0g6KjXtjOjZJPG2FlMcbPv+KWFDXzmRO20gaKz0E
CNl3ePYVfTUqkxOSSfeaYD/zMz4K+D4khQSF3aArfiuJr1jDaG8SW2Ln6i7F
75MguZvhb5vjxKHRE6iAwIH0mCVJ9egeZiLzGDPqI5fnJ52xmXnLA862ePO5
v4mWsDMLeL3DiDDXzd2hJ2Mw/fobniQ9Hse3FAyS7m62CRuIgnDbp1mJR3+t
K1Sv4wQToTsjjPfUZPNJZzHS2cT+n1Mj3mft3rNVCtfq+yFEhkMkheqn1abz
29fqBiY5gRcEyIHN5jJnZAE8xcXqS5uK6XZKgTqR1qMyTXH8tF+dSfI8rEut
wqGc5zFtjbjQSeJN+OLK0vJNaERM1/UsV1JzZAF/0Q0vuRg3EpsHScB6hRCA
w86ywm0xicM29GZKa9ycsJfi0E0PtP/7TWPsMFJ60eoFOSvioH1kDdIazNJT
1ZXMoe/y3a8L69UypP9J+vQA6znHdJYzXPHSu3EzEzcOOUCcvuonCdsrw0BF
fjGLUBV3x7qzsEUcfZoKCzWSZMmexrrYJm9Rib6jXPbhpwbpo7kVP1/brNAl
9OYCGjHitR1z5dH/QO0dVA5DBGqfY+cWVNiwZEiGrnjBaNPD4oGy8HpiJv67
fpVQ7TLypKs/Ta75U9O/CFpD9GymHTn3BcCCQeOXX6GjZVUhbJ2ianDRUoIF
MFbLAvpWjxnnPHbKUiusWJCMg4edWpFUMCCdzgxf1HIpcrAWHCpIsKrbS1dy
B9f0Bw4EcMILU99RqjegcEtYaEHmznsnCeXFvQHWHhi26HrPgyUnUG0rzOau
I5UrqQrwYmouuvhqmbU1NYzRzB+KxKkxPAy7bq06KgPx40KTONpBFAr3nMF4
fOgzfRe9TVc9IEW3SQ5tTNI3DnGvoPeyi6Ej7OLJui6nv63zpcKtpbArO5CG
29GYgcNpbPtG7o7ZQsrLCYhsj1J4vd3xAp6MVkPHyrgMFh1gN5Mb5uCiiOV4
bP7LXip7vbOZ6jusSx5rMyaSgenFppiZycDha0JZiPriKOhPQMptUjwR7qSL
YRdaanwuYgQPBmFOaSsnFQjHeCDqeOzOL6ZIoelXDszse6M57pUgu5/fwzWt
9NHPE3WkTOGEOy6zkBYD2wBaZj3IactJ8hAGDKOh2fr5HCUmyhiqzGfIdahI
pwBgntw4TuTOkOryHp9iCmah7+Yv0ujzI8WSMTIZSrAU7kuq0+hZ4w1ftNQD
uqcPVtU9D8w6uBwo7lt3XzuU0IDmyP9QBu5kBSm/Cq4sahEAvxdSB8VQ55OD
lhIC6m8Cl/iibO0dhTkYVA5AQTvmlZ4HtLFL5lZZr9otiURvxsELOPty2QK1
ZcpXhnkNadZB0r7ljLbo1F/85LN062wyRHA3zAqcYMTFTe9vjwLdF4GF1We6
QglDTFjp2qEGK5qmFHbhaRMjmTTrfQxb/wsVQrRryajn/Ptyb+WeUxPW/Zly
3k2hNusd77baeWbgVaJuTiy3OVd5E5H2GJ1dxGyRPYnZOFzl4PdE1hb9Ubyv
aRYt6eFilqhe6jMNs7iqsFXrROB/JMavid4HRQMn5kpMTKQZllVy+DThl9ql
e2l7FkKBAEAnukcvRlVDN4/1/Ev9Y9+bbo4UsOnLjfhZwVBks6lf1SnJN5Y/
/kWgZLA1X2ixb0bh7UT+S3Llpb5xxHF9iTwSdy60uUFnD3SYJJCZ85KF76/B
tGuL9HYHVSX2PKjWV8VxKaWQwpXzNReh8rjFIZw7RB9yWeqBmI/lv4z5SDf8
6y+IZKuz44WjQVEJGtC9H11ysbucMDwstiNUOd3HZOKXkkTAyByQf2j/Y2ff
Vas8TQDKSu+yGgYHa3DveDCk13PawwowVfobG4SJoxAbD/VYxu2a8XFqeIue
VTxWTsV3RuZUSbr6IKo+LIczpIx9VKcMXDKXvIAMmzZCoovDb+5uFEf+cMsG
grgLBuTFukW6OfruKrfFsMeHDZ5qCZi+/IGqsxiFCmJnFFLuNrcPfeOGN3x2
8Rsg4B7T86nkHlkzAijGXAa+v6+LAaP53mGwT1W2R9sNNq2AnStNZZps3+Ws
1o2VlwRqAvcBnwr2BAX5c39VRZT6dMOBc6x08HuWHaP9hSyB/6dFINZOErQZ
EQanH1n3WkaTWmAJqSpXrvVOTKbCJHfMixrVnTfvi+rgNz//Z6b7dw63GQ07
CFW1QlCdz4xjyD8Mk5SJ0qra4lknZPdOe+zpixi4y8KsZJn+1AARwJuevmbu
dvwY0Ff/ysCp2ptNuz0uH/A4N1xOnOCC1vlpMVdJrniMK1juZQvmtBJ1pNeJ
Lpr7RWAvn+uzhHLBAAxm71PmWxQCzxCFW4JXZjfXXu0ISfFP+B/rk09YSz1k
0NIX61pBbRDg9vyLz9UZVFlMNRyG6YzIZpAgt+zoHYng18/wjlaMFz/pG5HD
2fcdoZQ4dMUPAWvcA6BQxro3edFuerGYFRJlg0Qbjs7c3ogVclh3wLLsrAwH
lxqsrLDOIU7GwtGOpiQCr+eYUYljfcTauHOCDJkDxG8AAQR1IuOYhJHbsIIT
7zwRq+4NPYJKvFzKXVwzEBKMjQ9sud6IhrcILNi+Rfn27C9i+ABQBXNDyvRQ
0y1fDFN+WmPgQOnu4BlvmVixJNDD0/j5oiT6VSmqukuPkI928TlQoFe+MIgJ
JHa0RKdgz/CYz1wt33obIzcOLBDUiAFSTRbX3bR3flbFuFIqrjvQQWzor/HC
JDQ6rRRLHVovEi/QclEeGp9cqgpJ0y0bzLdiB8DtkNoWKhG5xD6Z5oYWGdJM
2EZfBzsWrgL1Hy9r1CpaEdNzMN76jobV3gBQJOeUdm7DRh8eWQMfkJb/YRFh
iD0NVKp5wImHouw52nuKzvwFhACbXwXNCw9U6nvCBUFL3+9bOEpF+WAsORSS
KXPRBeVRqyYXmv6GujO3ya2Z36t0j01TDocf7OSz4W8yuP3qpJxLWwMxQU/b
NT+Zbn0GLHSlEYZcEMYKx0MB8b1nUei15UEFfghsknPYvPCkV8HHiQTWDf/N
ZJe7JfHE0xN/4VAuR/nbGspsmB8R/qhJJ/1tRD7YMUOBW7sy5M1wjF3eYqh9
x38amkAka1cqG3gQV6WhZlJPLKYHnWoOEAfmqw7HwfdPqF49sw2++VLqL8Mn
HDfIDHXpanDQ6A89Ez9vHbOr9XgNr0w6tsuRx3nGPHPj7fOaFl+zIIb3jzcA
OTMm5dL1urE6FZm5Tc9N2mj8AxrEnKD7fqdIuxYZveMHtTp86ne0ndYLSJlQ
ZLnVb//EFLlo1LViHFw+VEzLXf2Zp/32onm1KgAWZrKGpyOJYlREfNxvjWnJ
M0ms0vN+nR4rAWs04/zGy2BOy9P1EQ4KPzoy3JFJuvTaCKBEWsPJ7luecBm2
h3IDeyu3Ed4uKDZ5DGGoZ/Gp0D8a4n1UjJb3bAkxtR5Pqzc2BBXs8zZ4eh3q
2aDPOM1v+r/zKUgx3XO/0gtssO/0PeuLxKvwL0PXK2wwgQ7XFsMtsbLMOtjy
w73b0p3mvW9GhmPExqCvjSC3UBce/P6eCdil1ILfMd5oYsVVFad2gt028A6m
SwfVxttt0AHf8/ijKF3uWQcixBlwUSsR4t61kpUUGUqFdL5k8zJDeLdPDFpv
qS+2mq2C/0LijRgfArN3FZatMzfdsmMo7uuvWDHyNVTQyM4twVd2okDhWnH/
U5xvCjokDTKuf9u8YVSSCl6ZAQNUdWOg5oqVXpEaYKkVJnm1Ez9reUYqGoYq
4tv+vOqRzfXld2PjocVwQJH38+/goQRLoYHIHWlClyLZJ6FiyFf96iJBioyx
l3nqEJdm5Plf0f3DZiTSbQtEaFvVS9HD+6BklFmM6SZAF03/OPhdNbT9Mwt6
ZKmQQlkLQmdyXc/EK7TTrh3iQxXOPTI/4/EfUy3mKHbRkl80xgffiz6KUtC3
iMklnbNHnEw7pLYXFsSyuMzRMJ9fzDk7S4dTRCbhEavKx6uCVExaJODpPkvU
aEkTUmrZSi8D6f5oB4qxSjRX8Z3ccgs93BWxebGvfbfypvbywP1fzyJK/Rht
5fI9eyaD/yJHaHrH9i2ZCmNPMNQ80d+JkVbtl+Sh24V6wRj/yGEEifolOuXS
7nz+ir5Q2IpQSuivcuzZB16qfx9G2q1eGhznfUAj+Eqp/lfy7VapO/qOaNSe
OgCmfnYqBMDUzgaPQ7mF+aKK6WUIJrqnRfC/Z9CEtrW1iERNj6PSZImyGwiM
fI0ijuBdsVeopzbpkPXMEznQ/OPVJdmHJIwnRk2PRFVMTppbcYCeZjMZo2Hu
F4KOxS1hv0V014TLlbbRl6RvoJxHsdB3/Ccg81xaMHYNcoJpHPGrid19y1br
8O6SSpdTaSoajw25GJPP3HS9oVjZDy4WYEiZDK9ObZEV6vRzAkZZpA7u0/UM
q3MwZY4m3mdzGlgSL+6dJyvCMjhWfrwKL9wvL+b91Coj/u7my4ID2DkAz0tK
EyRg1Xqlp8Z20MiOhQRGglO/pcaxY404az7PgqbniiS4haAdl8YKcxe4wZ0o
AxBT+6UjPXjqkpNBN5M29VgTNwf8HPWMFqWl68DMl2aqLE6/octw09Ngt75V
PvZ97BETJnnaVmewyvWz418NNFnZ7GfIzwMX6ZCgXwcMoyRkUI3MvwWGgUZp
+x9RLzd/UEPtV7SIiEvT1GUox+Y5o6FFwHfdfm/G/TNCVC7LnWZkR1gCEsiI
Uawcz80ITUmd1iCu6B+cp2I01np+dpzCG1LdNZOcaOOMdRkzyPxRH7mWasAw
vejhgfJjhxk3pLs42eoTFQNm4CMNNYFd5AzfFtX28Iwpdjgi4SPfa4RUv9Mm
n6ANrby+xHXk8dW3M4Iw4t8FWUZMeo9hrihfrcitk199ZwBJxPaqeXWUcksq
DDd+0jKz1RoKZaPxS0jimPA9WbJoyPB8MCWjHHiiw7QSX9BGfBaWvd5YCbAq
bIpORYy9a21EhTjlSvxwo+Elqo1z/eA7Zuc0sRtyL52FS2aFJ2l0txZes2/y
jaL7lMzIgLJJkMHXYGPkSQTtX7FjDG330HMkJ4ta27A4d2HUEjmJ2B6cImri
X2uBNYDVs0MErannS7aNKpep81sv5UPZ/k1+d+hJ/c8kOcL52YfzU4Z8pt95
2TFOJ9mg2VM4QmsvXU+TR1SJTbWzSJhcaNqpsMSwGgvqRbgbs6UKzzLppn3F
ngklmuSmLPunjcLIhSSJHt0QtaN1lccNB1Fp920vkURXGwUGQpl9e4xqWdYh
2QILTs4SoUE6rbfQ7n0/3BISBsYvtfSvbB2dIZj7Qyr5oL62AUGubBSiddLu
Q6RYGRpfBU3BO8Dt1zTDyPVi13cJXqEQQvBXirNVSDs4OQRw7zeUuEI02YLg
oUMy7YrU/FB0DfMjtekpI8R/BJaxvHtBOt0a00B2l/eaZZLimbg/4zfeSeeZ
bPnwNvOy5oApo74nHDmwr8uMsQKmAVeW5cma84UZkj7P/M2hdt/tB/Vl6KEA
/bpzhP8uu5o2HDBuwyD6Td46Wu4HCTAzIfG97bhB7OoD3W04HVQEnwNX+cPy
sdjuz2F+mJBTw039McxEUnQBx5qqbKtyv4VEE9wHAwYC5pCgEwshHiC8txiG
RaxiBrNwxPNd9z7g34ugboIk8WWLPU63MWGcNQnVwSZMgjlhMkugNfaUgum2
QEq8UtXfqIYgGhau+tNE423x6eAR6F1Nv6VMyVpkuf2oVQUSKVPYCTDzKSiy
A2UFYEfB0rGYJcDwhL5O2SEWn5HcqH/4mH2GYIw63O63q77uX8bNldkHV3Eb
Vpc1eFN3Cd0YfK0FDiRZzPqUl10F4hzxMvpzBl4VwS6wNlIhLWLaxEwlPKlr
XiCJPWRPSU8PUQ2wD1P2lpekYzjp+r+9yvk1GzOzdUKaD7Yz3pLOa0TuxnfR
XbZHWLIQkeqHa9a2I5Z0mTfdbQy9JeMe0Q3LRRY1QEyTG0u7rXn9kvAucSlb
Em3kQjRPOK73fD44egXLqdHQqRogxVKBEW+ZF5l8OBs8ndj6Xh4AmpHFgL74
XSsWf6JVpakDCJCGQs/bzHe7aR998ab+dVQxoB+us8guCYDp0QJhKDXTK3k2
0lqhmEGI8FjlBbWmOG7Pt7yDgmVz7WbLclsAJUBJ+i4Upquq92pZYLHAf8vu
/EVKkH/adcHFgF2Pj7t1IwfiRBJ+1burqWj3pcxHnu4k/K7ZbbHbX5yFbQPs
imqDvaB++Bb1rYNmmEDVqRHFCvr5Sw+TfjAWg5RaCCi/EfwdZRz5CxAy437B
azljHuMVJ/ZvVTdSN8VqBz/LXB8MBfJtkIFHeXCY7+AUX78MceVBclYGKfdB
HtjwTG5wes345tOdW3IA+s1uGBOW0p1hjZydmtqZ2o1gTmu0VPryf4v/qVs8
sqhd8YYh7etkmkVd6Ili7ErJS9+nAizgG76zDL0V2QjZXZiEWTwYsLG+ZQ/M
J3x0mnZBZ1wyOTL6BXHr6xt6MkJFrKaJAlk3nA5VvtvQDWUVSi1/xj2Wp5FL
JjBBcLYNJ8JzlZ385R2AWWxDKlOy+6/5Q2X6mOB16QiJ6xFPSa7WPOd+HYQc
4uprLpqm0KnjybMfC+b3vzUVJCxv+ZiH+ZDg4bjsqPFdnHXtfqqASRt4qi9D
CGByn2l1GqEc5jvGSvwlScrmLp/YtG43c34XyFYXHkqjiFB7+060PLMWzq85
7DYAx4fszr8bObUF3Woo+8WazfuTzPFpYR6TuQ+wgJjksuEicnM+hwMmbp4w
KFhKcwU4LyQJ8HHKPv7iXLfxCKllXe1iAivYrdFZFPpTI87kDRg8pr2fZGRJ
Pud98EEMqXIJd5FjHt667aglhuemS7HX14yYnYzCw+2+H4BKgNyYE/phvfoY
ip69k5pGAcDBV9TxUxe+FwXxi91AEiSWWHdzFe0TFYZsCPy+pWwiATneDe/2
eKfe+q+CvY9ZImh+rXhaSHxST8rhCuNK9Q1yUpF4t1KGUO8pck2zYDRfGGcy
MrL9Ud6byQHIkBIfjR69GUm2cZWpQicI3z8TgFcAbqAnUSc=

`pragma protect end_protected
