// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KaYMElux+9kMlbpEN2ta1I/2n5ATVs7xB6DMAL/JiFVna6DNtR91LM+RGvR5
ZXUjdogfPQJfYk60o/u91F3S2FvIMU1IZLN7qm8n64ici/6/zzl9Lt7UHGU8
J7fn7XFpQuv4OPS7c4Q4Elyc5CQZC1RkpNzp+5P5701nZUJUqHuWql4WoNeG
VwfaaTzCiTFBeUdeT3WNENBf7/vEHBANyuynyaCBRlCgV0MFCEe1+tNrByNn
DJe0c8gI6Nuwg1Ox/H3bR2a4hWGuXA/A//i1PKn73fQFWz26UDobq2BILh48
SW3jNRswOj96W2KqTIOnYMWSY+60WyOM+0gghe+wsA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VfUo+7FKEaz2oiHfCuG6FeN97VPv4rwpnB39XhY8V7mOSyd3RwrrlyHCXdjE
6Csu/8qLQVldiNsZezjO/Qz+DI5/bW2ckueH22Gbw7pPFTlfcN965MOib5+A
Jyg0MwHKD7KJMt8l27BJnGLBY6sPCygDo5BM1gUU0W4doNdC/zI3YJSgZtDd
vn3PFdzqLQd13pU4J191BBo1ZPZiILkXk9bXyt99M28caffROu9O0c0NInyK
8gmV4a4y0W5P+X1ICq7dz/opK2a0IeXatmkbR4oc8OuJ6ppj6GT236k62AmM
zil+pWKTtM0tQXPoyYczuNlOMocLigk9jdonSfa0xQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iNRknznEAOQn4lCEt88pOTYKg6C8ESeHvI05jzsOw6+8pWIJ++128blFhJD4
sYoRJbn5QqjVmwLj2QO6zdXcyKnXIrNL5/qJKP4YHdbp1KTeJhBjSclpXJPG
sazbNA405YEo0NaohEWdjp1KsF+HHzlyomLxhj0LJLg6AxtKWLiMuh4ob84W
wXSAFaPPDxGjws6ZIVeMJ1bEWPtZ05lO2cWhU9qFEI2HbH1dKFdQqsE2XmPq
yCKtVtHKTXBy+w3M++3/hkNvMDsG201hMcMF/xkfBds+LBWRknEjNYchvDhi
+IyjP8E2GuTzLzcJW1oEwtYxpVPfd4A/DyIYWTg0fQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Yz20hvAt+U2ZRz3+b/tirl73wESCXhlCiOvm+imCwx1WTCuNnKT1C0BvlwDc
3ilSfchsJiji/tRch1BORShQQWprkAGYvbgbaADplDEmLJuas7H4UrV+SxTQ
Dp6/qcJ14QaxJEEKZRpsspR8n+gBomHnNa22Nsvnv09CS7voz90=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VZOwV9X24ynfselVKIrI7i3t5n3Qy+D+pLNrLnwzw0R0D/vl8iDbSGzrIy0D
ymCzlrpCMmjvpRjNlNWzG8RjssEqxswl1cZkO2kRL+9444bo2WtTihSEmoIV
3sbDBalw2ZebToFJcSPRgQpm2dp9v6+fVUNr+D5/GmfsBiTiFnZvb0Gt7l06
Z7La6A70iOuOoQYSiwpLwz4ZA5BdF1noY/f9lSjzEMDnlqUKwVrUBUYFAOUy
n+Bd/NosjqAshksSWimAH2kLXXkoNlh08ruJ1eulb+bB6GIgTHe+elQopNuY
FUEbABY3wy+RnOVkH/wChQGV+exDQ6VlTJBoRWHTaL7e0yuBlhbFF+P6tofN
iiiwoUSt35puXyFXqtt1JRA5Q8gY5anGhTbgYBvSOp/SWq1CSqE6DCB4gBYl
gBl9f/xeYAsvEU5bWasxxuG5Pb6ecgPgsCcgntqds3H1fmbGaCZvllzdQbtX
zT015/SIJOnXPpiU59bjR2xQpSwL/cKP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
j1mLZYQXQ/2w8Mn+ybpy9bTAV/5Yl7a6ombhrR1zLAz7bb+mthDlsVeVNxiz
zYXivhNSWokmBdHhE5mmuGHLwJuNcCJD0nhMimh0r//ATy7Xe+w4q6ZKd7FN
GnVxrhqcmtdvra5vFNg2tR/3GsF76TaPPnNt5rrnqI/RQeSWYjA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WtswoD+hYJDp22dei3lSu6gSgapgVskx34B+bUH8FNdmtzxWk2aNb+5GlWpn
Ct0FVIwzsVsRzhKYYoWuJNjBePahD9oYdixCRaSHmDNeI3IGXgYkHnURQM8X
fAsw0A3PpZ6ZsvfsP2CqDH7x9y13rk7d9vQ8kuWSB0fqiZleGFE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15088)
`pragma protect data_block
01C95lRebTQDN4c1Rc1LraUKB2K6Ec7GRDAV8VeG08V/LySt7ZGY3+bXl21Z
7vewxOBjaEkOn+h6nxsIxtP9Zgr/tNUlEr62kkuhFNthcnRiCr0H9FwoGyMZ
Fu767zCmsVCixnwlC1O9dbOQSoDNmb0oDN/eyjMmcCdZ+sO2fFYvpKyV/KEs
LwcDTjrmjLb6CnF5NMTctTsABQU4/XFMVco8krjNVk9Ka2oJnE3ieMe5rc08
Cm7L9SGrqc92YPFEpHhcOAnPoCER7IM7+qcTzLyjkEotmfuEtv8cRWNm15Cx
igc6bjdc2Ygj6siA1N7cnBuoOSz4L/CpqH6ADRnyf39dJB+5HF3u6dkz/HYA
mAjkeibpdAbV5dsdurBlU4z3ExYXE/0zIHTE8q3iVGnEUrQIdXGsterUrKxs
Ja0e1MuZW7i3fDTS9kZYm8PCvI3SJFV8gXy3q2kBWmNF/Vmj7mPQjX5vJEbi
QxYLggjFOQcMxA9X/DTr9RJ81xkMjdqTc/SL9wcl8KxfVBKkNZTWcg0Wk5tR
7YG2rAA/mi8U46oe46DWDnlcnsLLF6YdVuyerW+F/hOs3w1IHiM9/ytClsua
V5LM2NEG98K173FWXvrSHDbclypSWOgMee71n5A0DIBecubKOUqHDGvUvoII
fU6PzZOebXMl5VmepmOt33STWFdkDUT+iHDSbmnEBB8mAd/Ws27bHiGn6kGQ
nTwGnFhY8yZJpoLaFpwdx5HTJVqNxwRWPcldrm5gwQn21/lvknGfI0r/Eikr
q44jHfLsNZUUNMWCW8DfqMwMecrrvZf8jAgCvtiXG1mjxtuo0902rOXzgGXt
vH8aJq15XhSsDjR6Pklhbm9oKMGavyo4UTtBiTsvNIm29uxGPjqkPFObxx5I
h+W3X1hqh9WmEJ6w7N2Amw0YUwF7DvTiCQDTDR82q4gGq4bZMvbOgjq28OZU
F3PzsilUP/le798AmsXILwOF0OdRv/cHWjrWXH8h/4UZ2G8tneLKUwsHMN+k
mXcp9UFQPbEiwcJN0ma2wNthkm4kkWTXL9oymE9VzMABxFYTEOrfbH6bJuoj
PSuIRey8d+cydRN8FQxOdetpDgKTfb4qLZMHZ2GUsGDqMsRHBnYLIhzdSdbn
cxD4Yqjs242nroxwduhl/GS7fvmYGWyOuFz/4f2i4XjO6r6Om3bZlLNxjyOA
kgi6ssQHrcMjxaf53HopT3Dk0Qa4FBMMC2XGLGt9k+GA7jzpIhoNYB3x0WSa
UViszU/GSciEyQ8+UprytKCGDn39q0lKI9dMhR48YIijob1psW5JJGvr1QHm
AkjKT7exav43joDgJifN39H87E6A1FJf5+RLrAZnmQpRmvqawhrRA05uKFH3
rwcH2gl8N1MSq3CKVI5SsOndh1OzrD1Q+t5E6Pq6xXNiAFYt0x+eR/dwE37a
iPHMHSrM42RPnr7Kb7VsrTYb5mP4ukSOccS7cwzsFi5gMqL9z4n6FJNmK4zk
nAdGek7YB6FYBJ+dz0sioYRVcH968xNLeCIxXjaMIR9LoPRLzvRSYPmAP532
2nIJUDaesVc1YGv7TNPmHQi9vughcoNSOlMxe99Ji365ztkN0CanR00ew+3C
SopsiceJb0FQd2itIxK2oPlykhYmjVw6KTdVW9Z3EKcTAeb21W66ncouMYhs
lCOswkApUbfB1p6g2lPa7B7LogZNU8c0xmSrdmIkNIaypJ4OSqmbHx+NHd+o
/Chu/40ZvileN4jrESB1YyBprhKdZpGWp04C1Bx46Cnpiz52RHnzlS7/x+/9
G+/GK2k9Ue18seTvFv6CLuy4gV1XwHUNbLbMZU1t09DhQFRqgM0+tScUyGN3
Zr8kxhCQ+WxnV7p5AzE+hsuxI3bHsQ4nxyHBKVsYwT27FE0H927srTscJjN4
TwuPb+YaIsgArEBNU0ns7mCQ19PPiNmQgZ062S6lMMYWu5AR4dYULmvrG2dx
RlEkpmie0GZcom2tVGPWC3OKcMuxoyKxZCvI/xEDwe1IiyGeQfo5hpPDLqdk
blyR/3E5sGncvSoEN2DtUf3oJTmoQqKlYbxjGWFjDtu1PCp/cjJjwXZtkAJi
pp1sLQJaDJW7DUu+4bTSqOWQFHKl2nJXEomU4R00jKUJy7Ncji9Ubx1+3Agv
FAi2VdKk5dpdHy5o62sPLuPmMRkxXPMHMYRzkMWqBV54scH3XvNJiLkVSfCr
ToYfhMq/u11SOGG9v8SMq80+fi8+iSRVXvo0x0mCTdlS0lcGFXPJZqADwVa3
sgKiAqQ1p+5GNIVm95N0oSFQdJP7iylT0piqWfjg9IRYndBLVQkj1TmC4HT2
6cge1RicBeluWBKFefnh/9zxqDnL4G0bJMNYPrzEyp6ZsfUcFUX34Wdeyk7w
+CACmH6gaBhttybsYTV5SIbTyP1uk0dKw1QteXPsTJwkT//tA8aTsXX/D8ay
Gg6OpNfqYJSCKRkcmiQCl45Ij2zs7/o167YLMRr3RRziDfq3+/izxE4aJ5pD
GpZg7ppO/c/O65pEvx1tyV76B9GXegg0FelDbMMkx8ptZ0QWGaEp1Jvr0R0p
ctsLRp/TOTwTwfi4zbuS/3XBwGMrma6BU5p+jmoYwskV2jC8aekm/UN18Sy3
/W/dTQN3L6PJ4Vq9m7U8KJJ3qe+wgefRCXBDjSzd/JUwNzQpCs8MzVYTZw/T
tz9tubTKg37tb0ZtqV1NnK6YFnASvL/YuzlsHWxsLxw62xEMhWq75lcJ8U0V
Hg2++6ubv3DfisaX59JzeXPT6nP7oS3hCpvUMeAUiX7WFBAL0biAVIkqtxQ1
mYIgznC7na8mlY2UJ9jGiX0exbjCH/PZOI3F3zhvjIQCSkaPDXL7ly3NK36d
oU3wcAJ4Nd7xWnYhQje0tGRg55TlqpbfWnMLgWkp1O60HpTZSGNAscrJxnIB
khn+HP+XDvuRv8whV6HyZwZYdomVxWZqaoMPBz2Qi4cxgQnkGaDEOpFwHz+r
MxdO2Eve2cuUYJ3awRKazD0sZO1CvU25BY/PDj23BUk3c5PGqOd/kd+JuDkq
J2G9z25I/PpSffvjGydZSBRtFzprLu222zynE3fXkjvy4USxVEDYTAWDTJuD
6nxA+JpIeNXBaatsbCPf+wjkaggJHdw3wy36lNAuTNufkI66RspsRcFJL4BN
2KblP6MD8pYgr2BMZ1+k4LsG1Bdco7QxooJK+oUBh14tvlx/O8mivOFNzAgQ
VPyT5SaNF15HN6V3pTNdiT1m4i09dLtYVqGY9WXdHVTbaDL+SG3iw/2PZkpJ
rn28l7iy0bXgM4uVoIBFsj1pH0HRpKBT7ErxiL0hZHmY5lbm39luzM/HI/IG
EpCuWtm8+z8htHGRkXLT4p4z5lylPNyfrGPN79ryGlA0mmpnOXWr2lLFOe5v
LFd8D4e9QDrwZE9wuAlF3BkTGol8+TTZWVj16egb9hSRISBb+Wz1KyFrvWhX
V/rYO32vU729tXZBKpWJHcw9RQ2YViDUp2H0aG1o4hts7XDDYRB+5S9oPDiK
bLV42HUOt2eMYpFFYrJdz/2LzmmTcI0UnJWhnTpxZ2cMtKMGfHixDS5TGbrJ
ZOcQ4aJAne95it22XNlVxwoE28EBcAALTFogBiCB14i7QB1rFkLKkpbk2LO/
mDnWfKOwwmwQr6euu2tGvkBkHx9mx69utKq7N3TMppH//hI8tzFQWhrUoWC/
pv+Xo6SW9frW4MLp8ZW6W58uq1NFxrsHQnzsjALA8survMExc9lHxDue7+G6
U4EyUkR/cm3Rzf93i9iGWa0j5qsq5jRtJZ9iih7WzMD8O3oig6xwckeqMdSb
FGZavNKA8KN52QSxsX0RjHUz4pq/1aL/MAnLJbKs6UpRG9SZzmM9zzFidhh6
0GQq9AjUraTqNp2QfDcSzA8lfrspnQgjLkqEg532Jpyf72ULBx1Ddk9uG0As
vg63unhfye+WeXfVG/V6W7zaEKFYWDanCpw8ugxiYtwrYXJd+9yY0y4dLJ6h
gWsZKD5lZYik8XllGYQdsi3NXJSDETbWvJv5IyKsyRx04ZoNWnvc1A+kWyIN
O9kxOV0xq0W9WOkrLcwlaqC8nZrGESf4Yf+UcLicLWw+yWm4OerZrq3zsINI
p+uR+NMaxAIg3CSqcO/p7MFf0wQZVqIo7i6QEhcA/Rth77wcDL5qjbmc6GpR
u9GYX64B2ObLjE//adX9HHN8EdLhVco/eO2FzU4Z2RBVhpWWZ35Q4fAKjUm/
wH0vWb1xMFU8wqGQDjx7BOlYSAmz4je1sJiox1OQ9IDp3MHjB3TnyFdJOGgz
gkrMskXbYTZZot3XAKL2tRRbNFm0qCovjumUiHOwRND64Kq0fqREo9KMcm5q
0NZATwkkwUBpn3uBIvAV/Wv+xe4Ps4kdotnJ+X8fUGI75MLqPU/FoMLJubx5
lBHrQyk/OB+Hk0SCWTlZZRJUDpKdtFVwsW+tgkz4yLmkijwsQ03yJklq1dzC
lYLjxvnl46K/oTJ8d6NUoPJTFbFenxpD/k+MbVFVrOW6lMvpptb9Khoy7kFL
lrwSxMk7BMKJTE1S045tUp7fGe7195Eob4ht4+AePHStmVUbTz/WzJIMYnDC
KhG7OUBq5QAfpWgKMif0tx7wsujKvRrDHK9/bad8ZfxMVgsK6vkieYl2wyMi
pySxTt8meba9ADbMlozqUBnSoG8ee9XHcM2uPN/JE6IMg2PCljlPaAGgmGo2
nwDYpi/7ouw6joYXT6M5AC7yRZy3D7Cs+VifIXIYeVS5PuYMmElIsXGHZ/Wv
WBY/Y0Wrivd+2DBjNn4sl0Y6tIIVCdSYSGjMuvCvvgZSbAkzh74PKEaDz6BI
+5knhCpD8eLwO9PsI8UwYR58kf0thTea3m/QmhOscJYN83X8UoZQ/xgWuG5Q
6n1hEr9yrxFN4eVDrSqJnQ7Ad1fIy1Hqp/fHIDL4DXJQg01dj4jV4/1EiCLv
ybpjSztDfAmathUvB307OZst3iJpSiU0S4dut1TYA8SFbnMD1RMgayGIHCw0
+wLIUxhatJrrvfrlGDRVAr1FanXvOOKQopwlzG24Q5rKS1mgFTfbpGINsnNu
V4JBxkasaSNkR6TVU1MSwI91LW33gS9QsP5BXVG7N5mSMARMA7W/yq2Ur+OM
btGqIhqM3qHnnSfkOLE1gPyBAL587z4UbuZuUaBL/TWQH30Ofld7XdIfCtt6
NzqwtXML6NM59Yd26ugvfV5iVDfbubNuVXZNCLYfC931zh1x4R7sdj3RGl1h
Eki4EoEUA/SdjP1Yq8qx8pnxJrewOJ57al771wA4ZfJopMhqCfJZ9xYIQwjE
b068AhWb1QiobrLZGMy1abB7JXvXUDgiKQgfTp5cNHhrGS806e8PDhsJ0EEz
fduYxPcTvHsu/+ISyWBTyf9go32baCDbKQwyNZsdfh25xPOHiuAzuE7SZjV5
8T666KUWsgRnldePStUe4TRt8xoEebMAodDYnUZabpW9r27/pe6VDgfQZksz
B619fVgrSaORgfTyft3P+9CDwopbzyOQK4YHcP5PiCcqxXr1b+YjVmpvQDFx
24KE3+w78YEJkhkHtgKmB83FbCbtFRE1s/oN0VxB8uMg4Vk8KUdkt1QCs3g0
yIhxw2hXFBFc3qCdNFTG6KhPsUKoM3r4UfWVsLwxOEYGPkopTQoNqy5JCPiz
NhUZOy0UwtfHKKxRdsGYPowxcb7tN4W/7OghklFmvobKShPFLFavfc4TC4+d
3zQCv8jwq3I9QfUZ6d89+oZfX4c30huUnUW6pKlsA+M9RrvQeOF1PjBTQsMB
nDMFXApgpoinQeYcXA1D5l5HsCJ7qfNyMujGdW9inRNvzBgpyBuEbGDUe4Nq
GbMN1LTw1c0jVYG6LS38g1osv9aIamgcv8dppspdgLQ1+MFSvX5VEvwHpeza
vDsQkqBg40M48TU9KvGY7R/NY5ZIXIu3y/MSrMEO1M0pDvmFPGDjTDYWVvhW
LuDlHt1uQ/M+VaY9BieFSdawjNWuDTSFuCPVZnQVnWy83Fh44QuyFDB9M71V
etnb0d6+XtxizwgqREQVhw5s6vDml+9L/74IK25KCN5AozeB5+CWBd32E4HH
sOl7xRChE/Q6m3io4GjpwcEJt2lLJd3GYslD9/pON5kA5JI4C0KwjdCacILf
5YHOogdU1NBj9tkYeT0EeE3skSZyaZ8gPMoksy8ITTh6ZGJJtbUGqHv4RMxM
eIR9QWM9m9JJY35cxpvlMOenwBmHv8smStXst5LJ3cSYn/S1YCU5LHQ622hM
4wZT3RgcBkNObj7zkAY/6cEpeQMqs+pEGt7tsk1PJUUAMWH0UKNOEIIKI9bM
Gmm7hL4EWqMhmC82qM0rHTDZJGPqahT0BagkVf8KM6LmKPtipD62HjvDIz/U
BDEW1DmDuhmE4/yVel+JxLy4Vz5Wa6l9vKiph360bPoQnI3KoASzxKQOMrEK
UZTfAw5bXPnWvQ+dhZjkgFJXwFnGakPF8S/DIv7u7A23IKRBNcWX2vYZNSRH
/7f4+lJrTYRI/UmeCg5u8gjZ8wOMOp3zGAE5zBvCI9Mf5W5v5vhZe7QsBeF5
WgGi/CVmVhCNCMS6JlwLaNlZ6a82Tk2lQekTkDdo+KujXDAJ1p2XOrFAMhIi
1bH9MbrNe074veC7j+zdOzahucb9+XsYve3CefQFUdyGG86KwCSzakbpLH1I
oxisr5xGhnpbApBUxKuwQDyNuYUIpQcuoZ8aX7WvKhvf6IexMfrk20QuC74L
27qzhoho6KnR7rv1/nZEZJa0h3lwiCu0AArVXFAED+mtFQg34gfxKGQGZefv
VMFXCcsLK1CdKZChkwBwS4RAW7SbZMVa+YAlfgwWJfTJIex50efYxG6GGnu+
lqAOIjQCLq9IMCG17eA4K5lkoIXTgMIjAd2/4Emp01KbDTt/hqRjohx00GUD
tM3s1+OprrWotBW4imWFrwJgNCeuOTuQzaCluGxeQKres45PWe336ggGt8wP
Bual0VGpMk4xqUPJnAqSJqT1059tGnH7UD5DfB3TkvutyCfdsKu1HhjzpNd1
HlA26suT5FiGWY+duvh9sLVcxsCvDOdR0gMZ7eDDZGHWC1ygYmvVcWSD5UOb
kpmiO8i5UJ5zflE5zpRlZHY6gxerZ5L8RYfUemi1ugir9G3BGqaCwJvpmjyu
6Dnqev+aqbRhhPuZfGZJfsk4lIAsVH5xmTC5E24hWTBVHvgMVOldeuyyo+hw
feGETeFTexTOpjzUffoK40TUEPWMpWbuHswT1p4ix/yxTZVo2U0I29w9lWI1
j1RkW13mtCneNt0hrjR74TLws1myyvlh57S+PBT6Lnqv+/fTM2yA8nfafDdd
HcBlJL0aLmIXXDSmQysYgO+nQDjMUblvxfdSbfVo7aHRLH+N95Il6YmQPt5T
lo2hfzA8/+4JtGIKSC/nEB+yHBYKGPjDqdRmPZStp7VulaFBz4UZI682KNgh
i5Bg1zMWRdDGRs/VaRU6F/NZpK6US1vycUnqzrlwK6ml9sOBtrjcGHuf7Wao
PAZB6XhFw9YcOr2r54tnttx8f6ABZgUGaSO/PF/rIjsyK1Nugtg6jlE636Vw
kcli+V4/XDtHBV4lgljK6R+yeXPbiRl6gPDIM9krICGLm3RceligjGkMckFy
4QAxbAY2Ilh1G6yBmWj/dPeUdGRE9JUsmtnI2Wh7Qk/nusB9d8QELEf2eJfO
+7lJ3T5sCj3xd8vzn+GKvrd8Nvhb1qXsxAVRRiSSFD+Fjn21WX83k40ESJOx
VtRItGZTy6ejfi2zC62QpWL/tGme8G9uwh03MXCU33Ku6NsyuV5aUT0vLZr/
n5kkP50tjofVrj4AuFSA9zmh42jt9PAtfLvOa/VCxVyz3AtngyEm8ELQa7dh
b9PgZJ8pTj/mwfqs7e9fr/JM5XMmdGW4czsehNI5Q0t8Ih38Eo76HbIIxtbD
0tOdcZSFzHXD38zCoW9vaXjqX46wz8OjGlZAw84sISPWwa3rw5mFwOGKxfRp
84t94gKN+F16uFYH4x4u59Xukd77LXt4ULLZkOi/zUljT2okuU7aZI+eMam0
72nZ2y7l7Gh6KU3dDqzDNa4N6fjLviZLOIbgD40w8P7smaATT4lmtF/KNr8E
OI3VBKzSjUgN05d0LBB0Qv9AzR3VrJEArGbNyeko4RH1fZArA8SZeiFDZAts
WArTFSeKEEazR/3r3o//9o06oZIz3ngJRE9+YWr5RMvlnbX+/2lD+UTVEkbt
ULgOMI/CGdiwDOJRaDcp93OvRO3hQDcM9pbmwAW+xEGJSvn5kSCLiViRizOr
D1BUQhL5ZIlDpwkGInfFuInW47qNGJOpk9XgSOE9X1d+aImE+vjhnLf5l7AY
saldbGLMpu3JyjOK2HfdlWVAE9tjoW6B7rngtvkemjGccL3U55eiERIhG6do
jAvrrx9l2IpbLtgyRRAnN0JPIVqnR6lSsE/QFGurz84ZU3ffXCG1Xjx42DYq
uJu87N4smvBWFylc6z5mQHmKcsjdgJSpDhd0Rvuv+Itw4s2NkEaQK0mOKHFS
MffbUgJtqM3o/pzVA0mcucTTxiYQKis1efElVm6fUiy1jmGV4L7cltjC1Cdx
RQ84XcPtZM2HC2z7e/HGn3AxL+wGn/tQ7kXvXeTCOPegqhsfwrLuksrc4qq8
JhwZyq5s7HO9ZLzGh5PRldHRv97CQEsFbtECHaUcKBynz/yEzXWZN/S9qVe/
+5xJJyCkqGVRwxqUrGrHXmijnF20pvWRnqVPY2qbK/rSsz2eU/qTx/reY7Ac
FCocLj8DP+vPbFeB78beU2OdsCa6aTJN6nY6pcNECZVIjihhjNXmUUwQMjyD
eiMCb2fOLoDomrOGmNkBw1UH5Ya0bMwAJmv55EbpF5iveG+KticCz7YMMaZ2
qMUD4IIvK2aY41GWBRrMoy6k6/tc/pkU62DfW9VghuIXN7r6fcCsdRdhrM0B
hWwYo5z9DdbyaF40rWYGm0ExZtkakINIUi0n+fcz14fU+Ci1HI/Jin7Z9v+j
Q3LjcZjYkXTRzfEv8g0grKCzLQgbdO4OabCEuCJ+Td+OUFdtirXWcW/UMnZZ
0xvSlH+FVItL5AnwG6cX4OBWcd6nVu8Qmph2DlWucjxQmBlvR59v/APM7L7l
5mGfHU1901Mset8GRGk1otLOUnExbbx5e2IslU0/WvTJQHqWfcsp8MFv0PJC
ap8eAYwBmu7MyAhRS1BMdeGtt/E+uU9D1tmcQanYkp+ZNA3XUcjGylA3ueW5
sYc0H//2scf83Kex/L+S0gi3buTlFVaIdkUjB3lKfSPuTak2pBZr5TLFGA2q
Apeec1h65hsE2mbNZuofF4smrO5uxyzPcQZ/B2lBhCo7AbPDe894vnqV00+N
qQeM7p2FL5rzAREXdXxUXnKmT5iI1RCJCkGlz3cSWe2pbNkdAKEEjjSr5b72
8YepEf0VuTGAovAsN4y4ClUBbECpYtCV1X0Q0cFP2QJoJHOMUsN6hdcygjKs
LikWDuX/jiYLooZfUozcvJySeHjEOMtjwWn/1Nf4WwQgzOCxn3b89orLPiRd
jHbXuiuwmvuYRj4PNPnYgX8RGVlKTroG1+H+u8N9JgI/ezOUwOabRBwlOrY9
n/J0xsFQMBp4Y7qJodyZuu6hdz3tRnNL/mDLfJF/UnFygabiqx/02hf8AayW
YMNLVodLVq1O41vPTVCuQH/tnBW/cCspNaM8f+szGP/nWMhsFW8xpAOKxrB5
paJVsQzT0VMl4HqjFuKdiJmJXw+WIeqkK0KxXmOWE9aJcj2gsHGkYiGHQmZ6
K7xIt+cXsfrSXIQbTIjh2RrhbEoxET3HmA1F9fRJxAbpAKAtbCfX7rSBuGtr
dGVeED8Uult2J0QqgLalHkrHkCwvjx7C4YSBsZ2feWLQ1pkhwkDjkr7zdnkM
GVHxyl4gtLcpAG546zjnId9SvOx5VWLDXEflWsHQ0kihip2VwfZ8oxFmlaiS
BnoRGUBrgnVkZJJvlb0YZ/uf/aDZM1Oi9XBk18c7dPitho14PZ5GE6msgFE6
Z1ewo6X1XrXXU51mJo1BxLVKOYV82UK4F8MGXRp3XEayEDUFVz9xudKazGDC
slRIXW5VAvkbJBj1YXr5M1XZ1q23U1kbNtOJeewD4oIu3PK5zveQv4O9rQru
MftNodlJCawLFov4ADa6DilZPQqHSJ3cbA99+hUTY0yIOtpzkvdykbg5b+IF
H14HuOffPdYn77FTOCEfqhBaIj2VfyJ8Yw5qsPouzGlJZAkYf9W7TrjbcIz6
kjtDofLI86n0P6mIFbf/LAOWOZpL5Owf0ZjbGuwPdsHKXBGVjG/C6pdFNp95
uXFHp6cbikgZdE4lNHbc8QyBM9xaiZd2pyhhpwL+wtNp4tEr2iDTYB9wuE9y
YBBM6JaeqXLMfSUD8rgy0VyVh2pwfv2Blan1TLcnxOIc6MFoiRZWHp8q7/lk
+7Ef5hp0IOBqQYGYzCzTbZa8XWnMoU1u29XiNfJ7+IfqPcLKu8kevKegljiH
GHSwzK3aMhf3/z/VCLesmnDe+OKmjHb7C6GCKoMKJ2MkFp0e0JZ2o7aOmX1m
MKQ085WBQnYQvdN3da/SM/PTvW5DVtfIbrthowXhuUCkp1aEhcrCUbXxzfFS
6Bo9uUxYwkV+l1VGjmtLDs09l2bKlYIC6XuOrF9wOTV7ntNHeNV8wSs9g9yY
A3MQbOrRMsKjKWVk3Pro174B0HGiPCFw5fjyI8T5kNY47VICYoQQ3mbYj6XD
Y+39umnzplDME+5+y0KbaUe4kWM3GU01NJsAgpDi9W+y10RARP4GaPTUVqzc
5wM77Vli9StSjG2B7/bZXeC8U0BmjkaNhj0FuHgV44cruiIkL14r0zmimZ0P
lxtIIU6yWWslMCFzmnKB/kNtD9YGT+ZdxJjssJwXXpUvpR4e3Jg/mb84mJY2
UbS2uUFxAE1a0hT6hyD1vWRa+BnWh635hL8NUuvLqN9gtwXdhf+UGY2XLM7c
7dazv50V9Xn4jqor4ty7dRDTOI6997UUB3+Y5iOzwddko20vZ7sM4tOCevjW
iC3BgQZ83yGlEXVa5sPQ9iRsrjK88I5xjJ4iLt5ha3t8Q7DKYgJ4S7Rlw0Ro
KbP9TtsHblv16dk99wHCf+hS4Vyg5hkjpK5wvsJlPs0SzirxssDc0olZnh8S
hbSWqvelJs9xMeZq2R85Sk4ri89BQMhNyqkrYeTKNHk3ONbZ6Q5g8tq2hU5J
Xq7rKQTsRb4ko8jtmL0HxXoIJFSZBaSTaMLLoZ0acykQmj6pUwnFpAkGdw7I
pR1WbnNbCBU40zvcFTTQ2WOG5mgc/OKBLRbbYKr9N4Q2rJrYaNA3E3U/kvqo
BTK87fGechEJ8xfgVh+soj+R+y8gkZ430i5vz6gWspF0moSo8F/YnccdKPVK
XMJDwDqqJmBPW0uPOMQog2TVaDFx/aleAPjkOh6fc7vZrkOjeJQxd++YMfPF
gE0KZlDMZDx8LsxTKZK02EJsXQQQVjPMfFBPhZpmRcj7al0Gq+vPx/4h4+f/
y1s8sUwW/2ZF9LFmMWn+rP7q1P0MixcpHMq7rGZCyjdoe99j1vXY5ILa63bt
Qf12d20U2SWMKB/79Hl2QGC+uFoHCYJPZbdzox6bW9wnSEAy7JIdDEZsq/Ho
mYC9i2zv6H23LgQQ/XUncAicKHeFD+1AVCNm0kV6mElX8Tyqf9rAJB2Wx8Cy
jmq0wJR3m96s0sBvbH49s16Rtww4SZpSdwGMKTHzCw5Kw9g3/KS/HJQNWHBE
Mxz/6PIwkiV6hC/mSAFMu3IipNqD9m3Cb3QDuw2BAd0xWKON9Tia4R/doQMh
TLpNi5Bkrq+wYcxfLF5cC44B1oyPSSTr+ioKJBphM4ZVXWGWtE5LU7wF1GDv
Xi9sDodLcCus6fieuoaNC6mhhVwyvKfowlmnx1zjvDYfInpkopsEmZYXbRBQ
J4HTz/iRdg8Q/FWQ9LGZ+nFaJuMBmEqiQ9Mq3mI84eS6BQ5bhOu2zvDTRODy
ARCxC3oAmQADMjAhOEe7RTCPJ774TVdSpW5oRpd8VBKMc2qwhnbiZTy09il9
CaqFhDwQmAeZjUCac5IQ8eFlQ7+klpan8tu41/wDBKib6ixqeauaTbgwI5yN
Aw5sdvLLyzeAFVIhEGHcc4xEf5A1Y9EApLJs84KnpeqnhzIXxVjJ2xmOjf0X
K7cp2ncoxczcxhQchFSFltdFl4dCqk7JC3Sjs0rVItse2fVxMweop80zX9Zh
uxeGh5miOsoL1CmKzix5/lcXVsb15WM1bAyUfl+oWW/BtOotg5mZPUUGKx6V
me3feV0EzsY+jnjFAcZknmY01FXpeg7/IhH4fwJQY0fMJ9iDnerKzCPKOiAm
Uzo2yjZ5TcU+qvMF1X3my86R6uQIoSkaJQs10IPDR9qmMH1Rd8uw/3Rc37l+
kZl7XkAICxaZcIsRUbEDVZU8Wzop+rDhXZhx/JPbGqY4jxMeXA9qnDnh1G4t
t9zvgiWKXT++GkCWqvXL3DjICdgmq+W0PN0kpcG3CCgOyhw4LUEF7IrbNLlw
CUSgSt86UsLnTa6EZb5Wo4Jp5KgiSgKLw/DeuP39vvCvFKDN7cgmyHq243IF
IXkM2lF9K8MTBD6TT9+rHRikBCUuzGxW8VwHdN5imdX0YqBaaYe1Rrp1DwuX
AKOEw+QUYNoaCnvjlJGc3rOKu+V8wMdtEeubLMT5be2rDV7NOA859Ux3USxt
U0ACkzNCN2yg/xBTwW5HqIgAls5VSzGVVwqXlh0zL5cXyBu9iFSIUUpyobvg
mjOxYzvtqVQ0ZwQikc8jwESrgXwH62Uak95/DztpdBTo8wtc3YsILvSmdfe8
Jg06v/LXA5ifd6YESDxL/fmQpgOaM9puGxNFVPhoSmjNdtP/R78i/BOMMKEM
zuW63JFzpWiSnOzoFU1LYXZPuT7sdNP3V7XIA9RdDpjtse57uBN13N/OHSpK
pCeUbBzGcMcv1rZftKPZ9C/+DLgMkxsoLvXIxMSZJplF7iZIoseoqYMHO0iq
wwVrW/wtqn4Q0WfYd8XAi927qTsCNcWwRWK/KU0qAuxIwIOWf7BoxIQOqTJ6
xSLVNscmQooLzXgUTcmUcywcHd30dP7VaN0sK9L4637BPWK+GjdXW+QcUP81
51r4nQG1YgOoyjVSCkKrQheTBMmdr7FiLnrPD/l2of0tUFbdFosBDJj940pV
8uY7d+tuttQX5aa6UOpzpsKFdBTTmej1ecwuSkZ9HTLHPupmqVQ9DFnQKXL9
2065Or4N8qtlYlBjTPjWOfIgQDJHnSClH7GQEffSyJgqo/Fk7p6XcdtsnZoE
w7eYcgAwzQ7PXzYft1tTRf+b1NoQqESRPnRWsabraPIECcFtpCXoxIw3rWzb
ki+pgTqN031yQfLn02AG0ysS0BArhIwe5BMNUX0m+qx6ofiu0am6CG4oaBM4
6F2F7jj1JWdECzL/1ht79pyWo4DEVOJX3X0h+inEGxTWe6UJ3eT0b8Hd7u/8
uFfkHQ/MHi88xe7U9et3I28qAMM8pg+oF6FGPMlTFhik7UzCQRfIRmFYQRYs
ulF3UErjRT4ILXsLNXltYUW9sfgReXOJmPUPLUt6fL0HZ1EwEr5YopnmSG9A
Bj3u+hQqaeQRF4IHyAZNwMpGTsYwB21H8cpOS7b66wpivHZvu5TGJrxMGiVr
o2h4YEzXlat+/6Qlm7K/R+Mxrr3lV2xiat7W2ZQwfjkzXBB8u0ikoryIgKXK
oaWT3wTneu8WHZYmZf4rbDsN8UyhVPA3M5s1wSc4zttyiS52zmDdSvV4yzoB
h7J76ehHqx4KUny0mDnySqUIh3xFu+wlc0eAug0+kxdeUuQNNiiBuNSAAvhU
fqBrCy0FsMB4SrlEqdpRWCjP6bBa+cJgEIe54WsI3WOLSlglnSdogrAT7Eez
Oiol4odXAtvx80LHLnlJtq0uEjktAy/YUih0g9EBjCC8P878fe8PQrE/jC9J
3Wpuisek9xhx5VvXEEp8gmCJyNb6EgbPF3jSb4fJjxzE1OYxsMOavMP2Si24
7v+CAv1e7ouW4u5pbmX+S6im3NlKAEix8gB1TWFVg3tpwAjNNvqMvAODTSVX
Yx+ziJ5vG6YaVEXXiw1I8k5F8vFrwmYrPVT0dxW67OlcIGsyf1u3QKvtzen6
MNMwAtYBJlILym/ol3O1NJpy4lIdtEnf2vGXuxdBOvRx0moSkcS7p63XLTPd
twYm1OpsOBOk4gOPwRuv8BrjyXrNSIYBo31WRMVbUjWOsRdr8OiBCC5nVbeH
jgGbZBA2N4fdZmtNHHGaqtltWYMj6XKHDqm3SVZZmpIEngEeu/JweBbUiC7P
mhcNhM/llz67KHndDM3PgSMGyL0M1zialr56/E/qBFTw1jPcxEHRnJvAuHOC
Bmv77ZWi1ETzNXd1FvBJjO/yTyNodGp5A3XGy0OrZSraFSKLGZnGWH5XoR6z
7I3JHDbhvlX0bzzIYvukdyU/xFLJrW6awyT0Zhl8MCuzIfLDmCw7Z+nSwbdn
XRq1TjTSYqP77X4DDsy48y/wIMgRk248vEn0pK1NCFdnM1V166TRu9AQIwmo
HkXsqk6gd9uG6hUy94DZCuL5W5WiGuMVDYyS17SaDPa+hwjCBbaIhFqUPnAV
KwbIqtfI9Krc89rPw73soHYmyd8g779V6T+6iBXY2dhlgF47FvOyHIlT52f5
hmSmDl880PG/kOmPijhmji2ANrxeTGJpuZpa9nlBPzZz4i7BxDG8qUn5oxk2
NZ3elHsaKdadK0UjOlEACK8mHNKJ3zDntma1ij+Aj8SFHsZrBNGRLhoOXlwT
HhfU3YgAewZaFh7heWiOSbKWmG4qbgUZKKYd9EPBZgjw9QfzOfdlZEWNtWdN
ydNWVyYZaoeXUL8wxoM7Va5Cu2GLsY/OJ8lP5el4feqheN5tFBFkB09I1NzO
irwrNXQuT1CphzSOXmOEoCtwFO2fYsK0fLPhd1YivaQ/qfqkpMdnlZBsQdfh
g3gBEMe9mO/Yov8w0AJxOBM9YSpHCOqRtUrFG5BRTTIfV1IOv3IWMc3TLkX1
auQjR5DCeOhIH8+otjfWzwn94Xn50cn+HXWgSCtshBPgc9srN/7ufGDHgGRz
uleRTSexIy5tDjOVaqB61wboTXRNZjHBJWqEVnuotoel+jdO7WZnlz1iYueF
S5L6vz1EJuMlRRrm/oXkh9G2evD+zJ2hU10MhKvavwLCFdCDs0NNRLwsrWjG
GMqnV40MVy44kofqJjr8EN7hNErRmfbsBT36C/A7U6Xss3yEiZMX17GMfGgO
zojytSiAxYy3ji24N/2EYYOsPhheDO1cAP2ITAURM1zbkbql4Cu9jtzeyq1n
bevMMlNhKYxZfVgYyPgbMih3XNtFHoLQTey2HvyhvZ5abnd3Euo4r3QU+y1z
3oU42H8q1eUAf6GUDTNiaOQknZuY9UNvJWHLoO1oMNQ8qK/oxnW44hHPfm5E
InvpH/Y3L1Y5dP+4OdkqI9c+/5OHDDWdg2FNkt0fDKWQM8ewiMqvGtfLx/3W
/YyJFDOkoTKAOt1H/AxbGcYpVAXHOgWMsocRwkyd4+SMPnScMUZAJ8WniUb/
7gwm+1MSkdL+alq3Q+IBEDhikpNXUUAO0nxo2Uck8cK46HUaaR+lHUSNOkY5
Uzj4GHDnoPMyyGx2xdld5iZceS3LxqaIIrEIZgEdNFcRiT6SiavTMYgmvTu5
OmNatjNvZfHfVBbui3V5zoRlf+qZNL5UHVypLkiSfayXFFKY9zoioz/O9D9N
lTuXT6N5KETcSkhsx8NBnWC5OrmJTC9MXJGuA5ux0lCgSwGRash7ybrTtBZA
nkE1wTtQMqxrxXpjBLd72ZggTMnpNgDSOP6bi8WiwmLNRo0vSNM2kxz+x951
rEvEp3fHMR9WEI/F3HI7V5gHwpZiPDtOzG0OKt7Sf/lJYVMfSNAHIfwxU8EM
wyzIsR8r5H1C5U1OmRcpgM3axnSIU4hWYzkcJ3UmsZyqAc4aCYY5X/vD83G1
lsuQUERHnJnaZDkhOspJi2SyKDaxLQEhLH+ewu3/1mlKb+Awr52MgdHyXOzs
HA7EAEJfNnV7Q7lJKzz96mHOydguqsz96o0anhkqMoWORwDanPbc2vkiiS7Z
EkA33rwFhlV+Nfb5q0kEE9cBuptyaShXS21Kj4Je8j+7q/dYIzGDA0oP476X
1ZWSguY+SGZTj2Uc8qAqBtMfUlB9Iz1M0i8RFgLyO4x+7PpUKtiaYZrmMc09
KPTQUFsgEwGJDzRFxbROyUlveox/yOFy5/NTy48NQd1F6NR4q1sBU8dHaqZs
lW7UaFnb9dEJNDpShHcrwD+bjwz7RL0W1cSOuleAc5ITYAnB00smjc1DsGr0
L+xdrbvvRKSNc6mUdxdsfE6eN7x6QJogkf1wdT5lRI8afKukYPxOfyAzB5bn
aZHEJiIvR7YRh6OTMxupe1VcPwSLpUqco3kwhVDdP3P64A2hSKfiK+MSSEDa
F1l8jAelgo8pA43dCxdmGaIQpoyqHGdnXxSXtstAYtq5/wE4OKYUsHJIXKoE
cZ/qTCCKmmWAxn3CtWOVKh8ztRE4x2iaKUi3w+k4EiN7GK9wh3ClwQsk224h
q4nPPE6awypoXwzgyWHMlyBoiGi1dlXcakJI8ccx+bj+JI1b1LNMM+vyK6BX
2s3pDaNxV7R60JHaO6hHXaxbBdV5b9Q+91XFpjl+X6GcjlVM7eM7PDAHX6LW
SPeJ9b+CLrYUFEmgzUneKiz534FB6WZ7DXvFr7xHG4H7a/3jqelV95S0fhE1
Qa5v/axO/Q5HvyZ+hRXxGhwfHlQj/D+bK1JWmXZ+WSDPVzB4yBN8GBCSkfm1
oUxPEpV24KnaWrxMyG2KqHJpTAfUwBug1LSjiK0Oo+DVQfCdW7EuLOVcD9if
kjxMFrNbKeOC3dEAnvphigla+r2QBtdMm+PUshz9F710VHnqIHdoy/g0wUyD
RwxE5tnWMiXkKpTmzUTuLNl9vKNRCKYZBa9FLgDDxreMJbBnH67zFx1MML33
Dc2kjGliuc24u6gSiOagsFm/fp+52VN4ZpJ5g/gvHZ/mrJ/8WvrcsJm1adCJ
U1A082yWPGLvsSPuNMsM8eRSk405wiyC8flrRXCFELoZ7zcZ6COnsaKKoTHA
JYBUPEYaLSGWYjsVj/Quff55Q0WuJLX7AxAkdUSM8sZ5uMn/nYFefyvdAuRN
8U7hHYmTPWf4vsHuq6DDmx5vtO9iqHWVwMYAZ8saBXEvrJZOO8Sa0cmD92pt
Pd6skNntQTfe/owyBHAf4Ra3MrcDW/ck3S1uqNyOuGS9ZUUYIBV2SLTPzFE/
6z7rFRuW8Z26b+AaLU844ZPwPBwlygqMFj9VwIp8ufLG4BlaNT2vEQl7+kgI
qkrUZdRzeWr6LOC+gM6N2ayYe2DhxCRRyxL+tbTJbPryoinpFFhTY8E4nWdA
8n0URGQJmS7Priz5rxWq6G/i1eFRmVerxwYDyj9tyXYbm0GHaN78MwFVxPEy
gsAYegrLc++ZOLacegko1ho/DuwXR9eCwSnp7qVaz4KdKpjRZPs4DDy2hmH/
2Wb3axc/DmWIpThEASVi3cP8Tc7mTDOGhIV4Jp/dMvOgjsHZCd/sIa7ONv/6
dSnvHaAO1W4gSDhKTmttOYCd2pMHrX/TLnJLoFTMSpmhh31yse658roczM3B
PK6Z74SlQzSh26R1UBFPXZF41WD6UFFFNUgz5zGcURdLlNi8VFxDQ0pHvkXv
0xoEgC1RF1ysqzFr3k7J5Jzy6BE7hzGCi/VSjxHYG+VBxCTGJ2oUVn+4aYRk
A3DuuIy7teDjvFEFxzKqXVm/vsQEqYCBcn8k7dXdcI1wreSucbcM4Vpl+SBo
tBCjbTB5xqo8vgRUn9cyvHjV19mkSXX2Ugn8TLy2HWfsguKuM+tHlaQijGmw
b3pgxQoLl50T8lsSqublWBUKjVDs9N7G1wJEuKXHctjCmrr+M08n7OsF/2vW
3CuvE6nmwd5myPCeDCfaXMuwEHkc7M8nKgITJLg6NvRBpgqhBqHLdAoXbbay
YxPYD1qaOsXhYpeFCFswdcWueqmKUwZe9BQyYkeM9mOuMifw7GeqMJEhT+sG
dZXmjnnW7bt3ipIg1eDg5Mk6fF+3JGIlq4MF149960khN4aGNbBkfWKqJ8SN
GnfbWXMHV9CLITuOqN1+sdj1q42h5UzMDiaP6zgqQi/Blik3SR23XeikRBBi
PTVxNkpTvKrxywRLqLJJicuHPf8z+3ADgl4lo6CT8VWw3mGmEUvbAqqYojon
sfyfXL6qgSw5FRHjXyliG1B9/3ar1737kTI0qsB7wpZ9RiCTQ1ailxWKp+n4
tk4q43VdOeAJXFx1TNp2dEJ/7UDjpYL/cclWxBpbGqNrSc5LnXb+hojrtzgY
Ak0PjnOTddIF/kBu6G9/qTLkGdUITc9FnyaQ+rLOE26VJ92VE82c6IEXS/ty
CYo/1faMAJVjzmVnytmKB4IySpRX2hNFeRlFtjTq44gCuFyyn9G+g0WP7DPj
w5jUqfW9E4COlCNv02VKxdsZP26j9YTIBG8EldqT9/iXxvNWL2QdrmvJxKk0
aIK8i/s3VozVAwg/bBskewZ6OraSGjCr5Drap4weFwNT0tvVhHPCIC+OVzhb
8cfNzeEay7OryHbDD44tZg1WSzeCyz1DnmCwv1nyzNk+JL0QBjg3RwkHuo2n
jj/bq4I8guS6kKRtEr9lcjHSS7tw7zBA5LAFQ1aAvMCoQe7Jg6kb3NqAcqmE
PIsP0HRgcNoyXq3HPZBL0jzOTOekYN7pn+tQIzFGpBWJLELM6793Lw+kLA2/
zutuj+A6y19UVK+s0kTwVufL5sGK+q03i/NAcEv+pdtBFqi069ytPq6OCL91
Ijq14I7/0YG9LfQFeB4b6rkqdq3kZfzMnhb6kDre2Wp2OigMz3Gc6GtjuICk
Yvlvnnr5+DKkCB5i+B5OR6axl/NDzlXXzrA5XCEtdrNsBKuOd8o7aKn6wYKf
V533tWVGnXu7BPyS6DJ00VXDU3RNwjjnlOaXCb1EmxZDwheMd6R5rFS5UZOW
Yem+OCAsRm6riP7VgZvPtjwJchy1iWkW8+TiDRCNQdPF4g5SA6G4KQOHDdbQ
huqgT+uSo3ZU2GkmhaVbo+T1x9+mP/mFaa5CM/52ScOTsMYQH/SdqKCBf4vQ
9ke/NLrQ3Cbn93eHGeETr+O3/Yg48n0ddCIIZIALhAhn+lOF/90liaEkst/M
mfYB+j4dvulhrlIgmgRieTNR0KI9vMlw98bAl5RLF6e/u/TTJu+GtoxUxdrq
+mUzRIwB5kAcGe/JOT83XkORSxfSBjqofXOTPPp+f9fBk9yGc2l91KngDK0o
R2un2HBaySDbpN0V+OkBd7ji7Qj9CzWPHVXIb+J4nUzw6DoBQS+4w6tzYde0
OrXnSX8xdw+Roo9VJxen0HIkggfAhhyWvBPsPgMz0gNieb5NUpU1jtB4wISr
QAoHSWv3BjoPLAQ4as2rGJjMN4Xqdwbixg/CZdqfZXvdafN4gI4MZGzaZkpL
cLpdHh2U5cdST79WdnBc5fW1+ozrQRaqx3tYG3RgGxPdk8SPCkNbqoo1FG9E
mVqoX0r4xCcefHo+R6wED5bFAOr7mMSO+Nni1c+Dm/I22tVxgssavBlKcwDJ
kHTbk1QgbpjjclnNQG/+MsTOI2WgC0FR36GQ2s7Cm0dF4gH2lFNyq3hceRr3
pr777/hf0bwGQgY1pXK2W/su3rhCB8uQyldotwHfPYcjalVdaj/sbKMr0S9o
7KB3w8GbGKCCnokkdJKlFm/57Vl7r9TtUwZ/vtysYOtA0I+rP0EYWMdGMS7W
obRR8TuRZYd1TNkdmQEgdmAlkvSOkvwdS8/dNA5oMl66YGVAtQcN2aqYAZKN
q8Qa/9OvWkXiHPqtTaDna+nW3Fy2YBMAKokSnf+jYk4EUWBk71GLoHVX67Pk
ET6D57EncQe34umy63eLKTxS7Do2r2mnjmvvEr9FtweAHtNNagmWTmYT4jtR
fl2LkOiTIxTAdAqgFA==

`pragma protect end_protected
