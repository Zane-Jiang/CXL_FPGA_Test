// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0KUBpH+s9ka0EeCLHr7XcNfBl4AcQju6QnIqbNuj6wkCBaUGPqNgO3MFY/dn
5COEaNKMndqXqva4pPpuEVv/5LZD55TZpIVs4I4pYSbcajZui9ycmPzh+Vf4
lgGltPeC25oPiMIQ/LtAbIhumGumTylZzkjDIGR0RpUd0JuWcIvswj2sJcGG
8SfEM1S+0k8oclDo7gWPz8Le5Rg45u7r7mnmr+6szCqjVZ0rMJJKpmkWNnh9
dA/TphBSIRfYMyYmzs2nkwXLLcZ9jx0+dJYuG6s8Q1Rq+UBpC9FV5YjOxuAj
ebdlCfW58mjDhNm0UkMBPpEPr1iRTZFQAOIkx+GqvA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I/h5zIQYOcn0joV175xVC6llCV3yWPTxzgbt6IbyVJwzOuz8CC/MEQNayEPy
KeVGKhmdNy4JST/UwZxLgVW3NuhahKmy4Ghpaor0E/dTg6yL+oLY8aO/CUr6
IAK0GT8v9XxCZ/Li89Tix2uigVR1kAIXX6JWMCtF8e2BReNksGzmmfOIlpu2
FBosuOxmAe3TPq/ZR5pjRFmAOXSa8GDs1xXqCLt1Sl6NG+dP/Lh1JnC9074+
UBjbjKL/5m9gIigUcStRt4p2O8sKQSOsZhW+7chg+Zb9HiLiKfUoS/ul68tw
KF5hs3YKZ2BQe+GKVBolpvSbr0zA156vRHa6Zo+LuQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IjJV31t5qRvaVtn9osU4XDUCTzSQF1swZR+IfAn8x9pCeWzpCA4ns+FtOzbd
k19sSpFf+TAWHWIIRN0T384tz7l0neCIyjRauVic75IN068JVECVHxuR6FtB
pXZKpYvFlt3miNCIKU/H8iXMuCk8BcgQiSe8OoZlG/uUPeYN7pcvfm4dhdcS
O63gEe6l8q8vOiE9wWs4w0COsYLP4WHCvZnqBxCIhkFuDdHEt0VkcZNEWKUP
RSmOf3YfcHRZwcFoLibsNa/dZA1zllZb4Qp+YUzjG5qxoiuznyNW0618Djsq
TNAtlSE20grvI9bNXabLAvGUEoA3lsOynlylpivxiA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tIzj9F/xpaXc2m3E49LL12uhrZSGC9x0sj4LhNF4qmhe7uSdcGOAQ5RmypFM
tpBBxXIvnmYtj5fQdsY9qs+ZHeiQ9+lglKqj1OqGh+cBuq6anLnu42ABJugQ
ZxP/zddkGHe8SmaYH/f2vG4C3ddFITqY5IEro/OlaMwnJttZaJM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
CLGwR73RgAKrk+F4o6RgiBZPFObb0IAkboAPYvh0uGREOP+HR29iRBDCwpp3
1eAdWFE9Ye+Vr2oXE7q++Rv7ElAfWPb2YBvKcdrGFxRxGLQS9GoxA1b1EWF4
SCaH/ELpB5XuqecRMaSa5y/l4S5a6+XggAPWehStyMkCVCHi2dtPLVvakld3
9zaXZZxCgSFpdoqsaskKwoc4pexiwhFAIsRlpSbOXCzu9ls1gNq6ql0bqwyo
NBz7Q6w4lw5C/WLVR5pAfhbWZXxZw2toi+lSM7l/hQDblJHSPFQkSEM67lv1
qwjIJIs6J5ezk78WqrsEjFO9G/3t8Pb0CHiEncreaXOYu7JS6NzYlDGS0zbi
8vL+23gCANT1ZTGozGU+4ccAKG9nMxoROHIQwSl/UwqPByyLpU2e6YctLmS2
w7gGlKiqXnYyXTUNYfU74sP7UhiXqtcVmxzpDie6/LBRpcwFNQma0fLTy4xZ
G43f3mqyAtxkzZn1oWIceJ97xGf5IWQo


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
C6RIDwW8mqMmgfhZqpqWKzSkV72sAu3ODQEI3FzFSB6CHJG5CwnrVtvRKcu5
Wqwr+a0G6JvTBrsZE6aWGPQkHw1g0HKprcnap5e/wGHpiaYgFFXrikCci3pO
uuGCEYEXunXbhAsQxqliIL3d/xb7INSP3IrePV8LUB9W7OmmqVU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OHZTnruqKOhpdF8esfCynRvAb33x49t3QYpK/xc4l6VCUt6TpJdPvx6MiTSw
c5nUKKzID2OL8C7+GfCz3JY8Mw5XWmIIXQ0J46IYLs3Igf/3RW3sMwU6xaGk
r+N6mkhmvzhG4ncvnPdqrZxpeHYG6ndOH4FiFz1F3UiiImCbwxo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 56928)
`pragma protect data_block
+NJiU7iNi9oXEAztuw/dTjdG/tQ2hD1m/2YyacyS4lQFXW/4MQZ/AloqDWH9
C9aAaE0A4iH/18f7uZv3a8jl8lOiwPXuVjHhUSpMSHWbpPwbiOkbz74iqw02
8qB2/M/sgDF++ZVSBWttPXztIwgWuYVGY7nR1r08vLY7XhnINLyyv2n9bTHa
xps/kLT1s8h1q5IbyHb56Zxwr7APgPKcY74nwUV5fii2XOm9oDUOHX9mel2K
NywCbJdukWebi9pdV1MM0CqYTtAHLjCoK9dyPcTq0hfrNQIecsA8e2dRi9Fm
mVoRM3EBB5hjCqA9bq1azh53Ah84AmNWHoRxH/iM4tG68Ph2ZJuZ+wbNMEbI
1dCWbyZ4xL4QFBwllyMqt6RpCHbPxR8mvsgKlD7Xq+dKK6DQgvEMnsmpGLK0
Ff6Cs5yu3Cso4X5HeaM4OglB9B21nFY/5fsCg4xHisXFRsfTFHWKI2U5QBGx
J0Mn97uuvOM2Oya5BkQ+kDhCujqj49jINNp9LKd3UJtstQ63DxINLXhGZQH1
5kSTcArtSTxaR6W+OmqAbEXpNYcrVTTUvavbPu55B2vG4LHuvEB0DyI07r9W
Zi221zim76tHBpc0U5ZalfcIdoh34GG2mTkXWvrqL45wuEWv4a6bZb2o7Gbg
0SH+/ThN3i4pHf/5FTO3ISjpkxH/Kn2kEvaxrSxPpkdNJhBut0mpSBUhHuia
Q0L9ZeC/8hukgszRTj5dQioN8Y1PQOZIccF/NkJQanzL3gwH95TgiqPQ6+G5
5386iSE3erjnMP07kJrD3oP1qjVr4kupsNxYdBySBMCSUDvhrB2BaQZnFTbb
hafVBi3u2ccCD1c6FRo4V111MsoJzO9Cx/u9uvG3zuctO9z99AUkB5f4A/hM
j9y+qcr3TvpRuFLR3KVJJI2x8gzAzzxmFQrUWtRWFAwXHTUlrRQ1Z/MXBDYE
IZt/pmvVIF79mSsdD/Vq4MFZQZgntilzvWj/+DesOf3ykjAH+ZyiEH9Z18Az
0lMnK+NnagbPKofrtnDiA/GP+34xaoHciyC/B/sZLfwjHtPz+LqGOfFs7Z2c
F8sj9QOj3eEAcUVtdnx+CfDUlRcD2oCPsK3xNnvVwuzS8LLykL53PxU84Uro
mRqNkW7ruXScC1Zux1RjyzXVgiXUc5896zxjxSCcqVAaKTwzC07dM7o/pEOa
taBW9p/QbGgeqEabk2dWw6d4jASZgA92IyiLCTH9F+tzB1nGekBw1aSI2IDB
pW3zda3P00qTzp5QrpoI6mqHytXfP7cHjlObl8SRPoyiQy3hnOfn3AnYcJmg
hyAs1b/lWSEOg+ei+R+0P52aDjx0KxR8rW2eLGAQ5/R8w+t19IbItWMeunVN
5Jk4QHi9xjPNrHfQSWcrkk4AmZ5PIqcPDPaGAtXRPlW4i3q6RxBgrpHUFSgN
rVz4qOWW+5iOUCQ5RSLcdkaMYzxCLt25SppvuTR9zLQ8zaBYx1zbRVaENXPP
KXq7YIyQ7d8adD5hFlJwnvOJlxsEJX1RgERXOKsyLQ+J5A6AmTzQMn2HxpTd
DLGmEpJ1Y/rLV6D4u7S1HuEoEgSSlcVLg3lpOUuBBB0K2IICZNzQ+mQJNeFN
/qxxdZy3eOtJZFB0eB3T09aQ2BcgAabBm5EFKDu6SUhje69qUIa7e41ixTXK
fT8+XkdcjmuoRcQEnK/epQGWMf3GXZi9+LRqtGj+GYrZZsHu9QFPk8CvbUPo
s/fJCircsAbH5tpGR8razkN7uQqrlmeVsZJTTFC/ikdkKA9NfsOewaRZ3Czi
PhJykChyh4Ajn42gkTVuioMgBSyymMyK9C9qDyGtDIwDXibQECAo4Su8bOz8
Fitivn2LTmo0JUEZnFUrq1/jvP5t6S1rmI7p3eTYyiA9my+ZnTss0hhqmhRJ
lJkT+KxZxdrzjJqhF1QqNr4TTkgfX3PKFo1O7iKFo5JEn2RJ16Uv+3gB55U0
DnAu/g74Y4bYcbzddgYsAAVc9OucuFW+ApOdogwdZP3Yiv3/HPfz5sK4ctjf
DUQU1vPh1UHRKfzU/CivPQCCKhQ+klITKu4eGsUVKnrEkhw+5mcEsMXDnkwm
31O33Ev8VDJ4F5oCuy7kapFo7nFtxcNi9lWcyGmbO3m3rPGr2t3EKe4BceTn
bjenignshhiMXhb+iVn0hvoy2BNLm2mr2d4JZgl8z81RabhD33Tqo48RxQZ4
7N0kdqKd0oKPnC3shobEwR4WVVwaq1lqRh0RJ8W4EgHYaF57JGJbMfRLc5k6
RJPl5tzpcq1SFAjLvpb4Tm0rbbsi+zmMQvhObTdYUnYoQ8yTF9nFX3MkJZXV
GCEmLdHBVSCuLmNV853qwskYJEN4fEu5/4eiP9+IwazSBX/xy7zOiQnU6wF4
dxLfb8PhJuCSSNKTI4IrFcJQKNntYiNjd/0HRkTmbXl6B4dVkRNdaNftdQAA
RCPFI/5vFeVmmM7H5/9U8V3SvJPSwVXomriIGSfqqJMaBVLtQR1NvQ5U969Z
+1TNLLXiHJKu0OogvOxB6wXsY6Ft0lFsJPiZRsATKTxGX8feaY5ytZcW0cz1
BY1AAxSb5I0w7v44dlW8ahRN/wwRyJ5OCwUqjnDiRknoQXXO2XjBxWAdobFu
MlEB78o4Xn2hsYZvQxPA+eee1MskbtLUnb+QwPrNVvd+a8/6F/SwFemPVdkZ
wyFqD1WjnKQZn1hMiuqw//Lvf7X2lySi3BD8WoZavMW61yU42IfQObaU6ulk
0cT6zGnef5aXlywKbGkl+tn+l5Qoz/ZLg+YMGPG408bDpXY5XCevKCne8Xmf
pzUZN1bfv5nfH60DN48rVmRXSjqZxyqL43mpaTAc3388yffSdFyb4y4Mwzks
GQ8f02tZ89b62FHob2Uh6jcn0njID+dyKWRoklhU9SMjXPfdcmSofnw5aO4d
Kfd07ZCWFBdUrwdUyBXtDIOTmPPEXI2jfHJ9+Pbsv3jsMFeBtJUC/8ENIVwO
dM5KaMudHFdy5wJmGu8JKgPEyiPrkXUGx9EwAYpgEkLsNoADHhB/eRALl9dd
ZXvUROSzqrLgQ1iq4bT/iuH3L834jefRXhHgqei69k/+WlSzfgXwgZT+V5Hh
j6SkKcQZ1IMClvL6A2hd2ywxrfHO7KByx4sjwbn0+mprZUPj4K5kdWYODxCJ
6GQQEiXOVmobptVbg+Cb8asbkAFhyg79bDgAryk9HczrFHVnTqe1+uKIsVve
7F/H9l7LuTi95pJzIDhWtQXcvL/F0vfCDy1iISq0n7HOp+AVWVb6xYifIf3p
iZBrdsuPZwi0A3C58bvUVQT9ChHqwqoPdTrFAHm0k4/nK/2YOAqBAdX/WK+u
HcGiCelbS0zl+PIu7ckfZvYJOs2zJFcAkgGKXHDJRl949+JcfPM5UaDo197Z
eOYDC+hvCjpKGDghFK+h6TGvaQBQwf3EpudoEIWgkeQVrwkA4jLw3OUx9jI0
zT/qONaHt86e1A4csdvUmKiLD6W0ugfg8Rrh8Gt/hLKUQo4eZvCK1nLoK7C8
yPXAj4KyvgCDj70jtydJfHd91lUt33BDhChbjzxkNDIuHuQFIDbVAghnwPOb
U/SzBKF1O9Bm/JhkdS5qJXMkjE8VNTp3PM/ZH6v4jbeapRuPyaZ3FutOtjK5
nmd9hGQnYCG+hDJnttcNlHsTm7HXFpgrlWwmRIZKH1rV0xOWBDpTR1KeffEk
sNzPkHMUvuOYQ8IlEAs4rQ5vEFUWY5braph914sQgdjXxtxbsmYgviYEwPqF
Vk/g0y1UB1QHv+pEukHcSfdjNvMG3WxlFWUVbGpvgToxpBW3C19JSzvApNcg
H/uTaFQg1X9GLEn3ZeBZggmhJSufUuLEk5nQsfAzEs0AcMSoWT8WpC5FvmYS
kjwbNgb+kBYmKD1eHw0xnp/rsSXpMiTfDpulOlG46ego7wmigNVXSA3kg4n6
XtJUOmsXlTrGqvSoeoUV9Lz5IwpppN8lUEeBhoy3KU7ypXrvt3sEs2N3Wv+A
0tW2I840ti0q5IYUEZJlOXzbVk5I4wwk35BsuZBeZSW3fS6S80q3cO2sb9/r
+w8sr0NsXcn7IUUPmZAWdc1lCrVCKFjqqDfh21tLRm3etf3ei5QuHCXi3d0h
gupO+ActbdgSMvTizJ35220Cht2ONYtr9aMedWQyvr7I7zlA2G+sSw2Ugqhk
x3/+rVOCZoXbePCz6pnNCmKyVm0Yrjn3wtPxY/4pPkRkjqMEEQWLIyQ5KOJM
pFPjce99Ej9ebDlZ+n8gY4bS59X7opbsOVIYNXLRKzQBrmmoGXHpCcazkzg8
TgMITD72wVG42RmGZOYHuRQpzyWHZ0I8puKyC//w/PeOPtmXlTvV9gdSC7AZ
sMDSA7jjsfFDV7hHQUU+z5wZq6y0QMwCd+CQtTpyVz3AYVnnOq9r1vL7Uckr
okuhPnbauAq3TUaUk8qETlcttImYKNOSv6WXejz/NWAU4uKYVQVfDMtBV/9y
QxSeNzGOIcc53YHWSU5OyhozLf3SqMoyQAqPB1VmK9pMfrPTpf8gB+pP0eJ7
oLDKz9JQ2OyPxmZgt6JbJdYXsC2ywa22qIHqPZ1VJvxqOvWAAGJJScBLAQiZ
rvHP2+8L5YaiTbUgMrjhVFO0PBoyBiw6jLpQDIDEqbV833FFJ8G/tcdyK0Ni
MVA5cB8kZfhKTbxVH68eOwg0PKeE7DuQzJ4yIXILWW6NOSPn66eKnQO2MBPU
NHz7RBhHMket5/0BWF5AwhzkggVNhvteeCy0gE950+1gOFpUiUVeqPT414gO
hLLZwaYDFYyMrygnN4MXztZuntwXxIeS+5K9Y8/ipx2tWqLIFJ8YVX/zJ+kR
OO/IbKxMfABYtwiRisw7oI3f5SaVrSk2KaAFN4YUy2OQQaMM2cMIQ/uUXPBL
+QpAxCHNhuPY7LFbpQYkMJJdmBEg+76CaNjRstDPDUqnCu7fnzpXRYervX8s
ddjNmKw1JTMxhXq3dRFQiZW+ZKcvxYE3k//k3Zmjw8fRmxMym3f9saRNBlQJ
ie+HwlyqaeE6liJWbnzlz2dbqtdJrVcmnwdxxht+z7tkwR3MxcgRuqj97xOd
oPfL39vQ06E9sK5DDb/XHB0E0M3ylf6tOgfl7u9EFOR4YfHmPJmSX+JwVmEU
O//2cPnU4ajyoGdacCGZBWfwOgN5teJ+2GgBRA6B9HjlHRED7MRNL+N42Ut8
E7GENF0DBrhZPy1Tp/YftOZRxKJsM1s/ghE5ZWzWhCT8bG5L7ZKMox1qCUhc
gwO7e525j3GYRvJT2GFu9VxNgN8xF+qgknvIdnEAGV+1JwCg8FG0vr+5TZP3
buPB88sUi2vd1Shk0lhsLSvqlUnb8l22B6x8EdB1Xx+2D8mzow6aJy2O+jpU
Euv1VZvpN3ICn4qfDkycGWBIW0FOu2B1+udK/TDy7zVh5J9gXk4OLZ4HpuAd
NVpi0Zm2BEviV3R5gt+t3bkOcYYsUlMffe/rdt29azaBbmXeCZpJvmnDUpm6
7RpPNqNifQxtlX+r0FKGNZTt35dbxt6L8kn77KfdTYrTQrSy9Q93y8UG55yS
9u61bz7Dr1rLbYluelbg8u9qSwHX3yrHRFICtBlcRwnByM5HKyOeBp/sQHlm
5P+dRhK6bEFzZEAsACIlf0O/p2CvoWis/CaY6LR6FnihmdXNZs9kvldt4d9g
8gfMy2cr3Ela/Guhk72ij1EucBNdLFQ3FR2KGZuGo3ZmSyK47rq0cl9HAYP7
WFsfx9K3bPPabo49RB3klyzN9XmUVH6osawVdRK2pbqmwkNy9pOimfZ67AdR
P4umVfQMOAnB0BVmyTcL/4BSwG8ny1hYr3vynZmMt1mnh0JKKeQSF3IPokf6
N8cjwWV/U0+4n1S2vwiI20KlRHsxy34kTaQtJGLdJigeEWHZqLyKoLAxDWXQ
Mk5SU3uhypZaVnto1dfL8+T+0prTDNJMFOyAWVyVNuAgBMWzqDbhx+cmP8ND
QfXrA80mQCsvl/L9H4SlBlJWbcFaYS5NkqT+IAZPxzU9Tvx2aCHCPtqzXTr9
3TPov2HPMw6nYbh5L+wxafLFTiGcuQaQsjTqHG0ODxPv1fFdz159W0Owyn4S
xkzTzEWRl2cnSVxEHXKZdHRg+yPDmgw7QRI5RtgV8bwYNR0biBbDy07uWbJb
0x4SopAOTzOyl88Ne76AcKgN01K5E8fNWIZRxDaXj+8OOvA+p+6C7Zk3kcGD
ClGkfw0+9sXZ8CMZb/uOMkR6T4Xm5jItVISr0c5lvSIqZ0phLUbK/tVelHRb
EoR5B4fcUdCIcq1OYgO3jXQFjDjelZCQ6VIFwuvrKd/SKJNw0BJ4Of8h5n/y
dIADSP5kxAN0xrfFT/oUcXhxkAxFYoVM9Vj1fVNPKxo3H0rTsT+IhL8Pikxz
CYsknp9iq6vmALB1RqBG420zDdtB/+ymCkG1M5kaqAJN/enSz7Ph0yrJLU8c
+BQy/t7WeS59VDDykVQc/3fL8cQQIUp9RhvE+ENNERXwCL9nruCifrHBuzV5
NhxpHx6HcDuZTSAAPlxusqT5ozhPXpoe6EusrOlvZvVmE2EgQ1vVyYHw3D1M
wcQ/8HU3Ys9ASzwyy9CQPhn592BhhGyi4MRp+tO0oAhro6or4Yvhb1Bt4LDz
z7FrIOW1zPdrVlY9iqAu9gRatB8WcdzfaUepcv2ENFxunq4kHdCOohe1DHQW
lwJZwqBorulpJ+lkdl96YcaC1zRJAGzVXHWMYIX0IFGkaglj9iyxHc3GgcBJ
CyuD/t4xROG3UFTk4U1eI1yQiprWhzXTlsQCgdeWx9rAlFo9SC8C9MfUjvag
MfiWBvhXDZScWMeJmNIrI2977OKevMtAEld3wW8hjyMG1eR1PKZI66sEkb5v
jFFWi6/AJ2mQH51ZHxF3M+u9/qdyQUUGUK4voLqZK87vuLdHzZwsteg0XVdE
BDBCC3hPOCPO6XfxywnPk9zvv0ogeMlhywO4n6P2mh0vo3/B1uFpesjkRSEI
YyZAczvojwDzpBOOwOo8GRSAy0c28d+kHi6HfMBtkq78M5FU7D2R3XVZ1y+B
9PGvyH5iImn0e8zaYa7DIg3FK3REeP+tQp+LeDa0tc/7NnQYYRH4RLtOB3QI
CM5QYzDb+Xq4ueVvV0BTa6yPErWR8geeWtSxfeHXRS/t5RfcpbF97VWMsW1C
JncUz++7Q2ovNJmBK3A9ofeaCBKo68efme2bFmbmx0sWLnMuwZtdeKKsqcwO
R4uipaJcDL+Zwqb2h1awX8avT8238iXwBTvp7EXhmhvC0trtavR1NcxDbJxQ
ohi9XbmBHwrowYXECj9VMKAWMQ99axrmseSlBOZ55JXh+SurjjmXP5PRL48t
26aJhDMFqfiznT2iGY+gDrX9/kjWy9I3EZZ+jxG7aeQdNqYyEtXjQsj4ESJA
cVUfP+ZlduXjgHgd01z+K3As41HmpHqZJngymmVma7+pvhLUwdTVYaxMKY03
uqKbONyeIMH06nT10vZMSd7zFveZwtXCOpkl7+NzGzWdUwzkr5r482VPxnPD
j8Oc7NrocWou85JElPuxjZZBSUd90WWxuQ7PTqtkCbNsk5o/B1qIh+E6twX0
t6w8lAlu1LJTor/t8JtQ/dL9ine8l1C0mbgA1VaTdW0B3Q2HRvgprBO8zqti
1MRih5sLYM0ydVZt2rqUGdZqD8uA+Cwk8BlzOa4VH6nKMW3LOl9TSg9N+dZa
lant6FO8U/cVTI5nuG1X/LRQGxcI+izArJ0CrJXjx2OSBzhvOHneIXQG46Xj
yvU7y7eNGWg/mkvkRRVWWw6US1lfHQEF+mnI79WMJnQExzYaCzOGHMBedG3y
KTXmofKAKuWBZvyImhFVbfkrO16G24Di3s5X1gyv9DtPGOcR52vhMa45D2qA
xfip4/zsNC0HInYQZh5p9xRbRYoCn4mxPR7y7pSAfD3zxdIQjcKGvzWOrx95
YNfP2Wxoc9G9de5i5dHTheWkXWyh80tbQtr/dSyomwbLItQIMB/iPiSV+3dE
P9HzbOuYO3x8pbkCOkFmt8Sa+z9Qs4a9nsx/e0jy+VwgCP3CQkDmPwoxm/a/
nmcLnnDSLKNvmj3v2aWM3d4GrNYu4XqegUKlISSp8H6b9fH488FUxTk+Qq5M
nhngffd4/hRa2JlT+dKXWSAUsyT/97JYAxBhdWrK0m1Ezj27s20hNpymYRHI
aVJ7/JH2dBY70ecgm7RVSvV5cBLTXD26AiH/W+lF0dzBQaldl7nhhTUepQB0
wdAorS0FoZcKaS7DNkKpDBgIQkMP6miX9tREd1rg84FTLe7semhXrlOM5NuL
IXadxkZ5Mu2m3JgrM69hCgIERWL4i+W0/Iwes6kgQhZLQ9Ro1r3sXAr3vfoR
Hu+rqdZCo83cFq0M29HkCgx7WbyIaHpJDzlgX7krHeJR9XPMRdiXiJE96hIZ
t+kAyiJNYWmom4AOt3T6K3tQoUYK3ZDizIOfP+Gd7JrjD+/lJph/nHFPATR/
TRYUdc3IR6DvR1tYbyK2lsL8gNkS6HdBuq3kgBWRnf22WK86sfs/i1wggdDb
0taIkwkqOqmdwfNduu36A93z2bhBGVWSEPddjHdWNU2FNQ6GDeifpiobhu7H
bMVBw2jRfnp2d5bLKroR6u0D82qjIjJFiL/h1ShrE4P3UBJXPO34NnBgZ0fr
kZUz3VnmX5OE64Q70Ye1u8q7664dHHkAcrgKw2j0humVyghOb9WgC/gwzp2c
L1XXQtXWBuDi4XZgo4PxvBsQRBS7We14nee0MPQ/NBI9SwHulA6GVKJEcAPt
G4LroqN39Pn+YAwP6sSuWpjjwRI8CzrAbQoxeSjXGA3AXcj5JdXk35lmSG81
4tp75vac5PHGjoNrArI+dnb72494Ze4lLYU6f/ktDqyAUl3dU9odWANSdMCd
wvibaS/FaNQTI8lnop4wSEnpwiiiXodflRchvXgTiiTEgNwWhbX0o+fuZBOb
KWrNnUpoYtQDQMLojTRDVbeKdNp6wI4Aulsn7zWfzrJ1Z/HrzPazisbG7lFd
p73Gg0RkWtFB6R67gQDuvuMFGzIvq0LjlbCLJsjEEtJgpm3qhVI8G820MRaU
W8Gmvh6Wq/kMB69d0INKuNZaUngiDLN2SXEtISOIX3bztqJS0IKyBSe0hdfJ
OooVkkXjNquZOi+936eiC/XBObNPNo8eG50J4PlYos8fzBVBvityu/ggzG39
x34m3r5arYdCBH3UpITEt12GlCi6qtEoI3YQ5GmhZRLYRsXpo+IIbhDza2f0
iNAC+xGt0MBhE0vn1gz+A/XV42UthCj9YgsJHsB5p8a53+a+bD0VxTqkvwL4
0/PI8lPA7FT2ijMsH+wxRIelGDazUktg25loFfJBQMbrdXPkkW3UxI2WUzaD
/6ulftaL0teYCdPRsebbO0ZSsNMtguTVV2v6YpsT1vEdWgMt7vcTYoAJ0ZTg
RT0/wE7oqLScZljkDQleGhkUDxdTdBYCod4rF6UvsOEjmlBt2cKAuNDHbvrw
NrEdbjRVmTcLYLmrKJxSPrZSJ5mZK/wRRbqP1j3bP39/P5j5Uv0pkRH8ueG6
yw1GmcRb3TedrHklXqui8yVaMT9ewP1aWd9nezVBFkADz3mRljkCn3oJijQR
72P8fH1e1MTkMcENQFc4QfJvzcfuTKSvEUi6AyaLMLJHJCKRClZkSNL9fDpX
WcdlO/Nj6REyAYmd7uU5GDWx7+yYyF2zwQGy81nKCTA2M+N4kEapFt1Cl0WJ
EhXVdQJH7vkGAFB03oqqgMh5LTt+ZDS6YEw3upsEHOcWMdjdpXD/hrL/8IFL
hioOKewbu4MOtc+edcLqwe0a0jq2glpXCpztxQhgcBy7GHq09+8C/sq/exK+
oheZI8jmCH9nVLAYJH2wKPHC8NNxnR5Wy8BAN4NGmxxizCe7qz+RJUKcSlZi
0FEABNYEah5i+pLQlklCBvLPwgjqWqo3Ojl0l3DKNcxDLFjPrSXbIpp4mmRr
oKB9YfEcU3KFmlJaMiTAC1y4fCp8ym58SDrSRecy5VBrYmGZzIJxOzkaO0VV
xt8EMWiOkpZrK0i3TcQ/etTfkL/DLd9g5uDe31MhDYfrBWWsKWzprJekOwTF
KpfyP3l/oilRpOqT1q4/GRdAFUsZP9Fg3KYR1d+Z79BFLuoUnls1PCJriKnb
DE1+cndw2lRHg/uLisgSzdtVc8BoZfNwSV1xsYgdgPdjjvB2nAj35jEAe/7/
hQmhw6aIPP/67LrNXmoMHu52TxtBK8pNqhvEugFLtVUwmarMd5arRWgEJF/+
v/Far5qfP+4vk98J1iEkJMTXtPlj1Ci31EYIqQ9rhkkB8Y1KkbpeqPVMtutD
eajhy27ELQ9H5QAIdX69Q6vxKJi+vb2adhfGDBs8azocyxsDUCBGIm73Up8k
we/epQ6C1tN/GxC1JjxYy3DbS94aKK/HLRhSEYSqpcx0oAKbS+oTktWH6WNU
EBDaD/UptZHpfHWP2NUVTpF5c1JA+QdjFtTCro0dn0Lr1O+4PVYtwa0x3Hk3
5tC/SM8YjPlVBBm/lIqZaSAR5auZoP0FUhXKYCYSsSQYO9diGQPZvTWaOF/X
6atxUkHxKi8yea0rjXVXfFkWxpAsT0esxxj64CZ3xK2aEH/PTZtNm09moUS+
NeajfSnjueyC3EtcKxWujor8wztT36T0a8exQq37mJzHW0+SRZ7E1UIhhrNn
P6eTN2oMBbQKidvyCV9o3Hgi8a3xrEd38xVmiexGEQtZzC2Ls9QBCgyFJ+Ox
yjWuogvNC+YSc1oVXsIP33BFbM9wJrKDRUkaqd4mSxJhZtZj86t+XhEWQL1K
gdpQEASrMPvPCM9q4lN5Eo6mZGIz3NyWTdh9jxA0NPjgJdJVAY4Z/PCJ5gUP
ZaozpUPHjauSRGRVGuqf/tz/sOO6Ccgm9leqC4Xz23g3bCF669JM+YCa7Ek9
IZXabu8Nd5QqzmwlJWgr3S1Wwt1WQJ3RqK7XYLJxPfar0HvOFJ7GMecYALzu
SN0RCin/ysW+8vsxWDzACRrwnLgREx/KBTrMTp6RDUI9wDIWLDwPKy8csOon
EZ5k3rOxzb9V9iMsBSqI+JXZZAXFed5WedAFaJUNTpkMPoJhOcT7Qmogb3gY
SNa7rbmnhuB8mjTVzrp1b2mDjQsualjOAHSp5RysRiMWNuqldzashE3AY0CD
+nzpNt0n71/OFNFojKjg7mobX+w0xJ4I/xAKlJ2Zd5aa/FT474ltDkc+sP5R
ljxrEFsYjElloDm1upigbXlKr5mFzYk3qhZ+m6zeVFyOklC5B25UDEXQxPyE
URNu/MkHJRDInEE/L2quow9H5FpW95rxROArjYNZ5HlzK+ZunwEOvDMmzfCJ
T5pib/ktFD02iiZZAuKlqystFjuRQG4lUZIQS7uTR7hB5TkTpHevKsmrKKtz
POTmsWMnE+Qztg54uaxZpYXkUE9HEpQSU4p9iwc/1jUiWRvQTiCvvPEFcorx
bv3FsShOkM2hL0H6jselo/kzsC/EgZucUSgS4IvWX68ciCRmrcgq3/U+KwPv
mUrLq3RB7QsM9fLcK09nq4rK0NUQjJX96LB3gjGunAegnB1yziUTMwI87nkz
Ud4l5qvdYO2BwCCcvGMbc2MV/hMG4NJe/HeH71IT/nNDiLL+1QtvSwqjVAy2
djN7ime0zKQ9cnOic5bHlcKH24yVfmK4zzCsi+vzgYv1cBhqY2A/KYqhUCmm
Jqvn03FxKCt6/jvAvSdHSSk/ATh2BTGoFDHA5Y+8cCVq95yLpjCdmGiMqbJ6
vnPeKRZPzZHXA3evZ6J3Mw5CALFOScZ+on+mhmXn6XdeN4u/kwVmGwKQlVdW
pZoQJ06wlJ9CBYoX/otJxgzWiCkq/H+hfXC/KsXg5WKFILuWxMX+mC8fCrDw
3MLnVe4wmsMAAayE0SmRloOpPnVOI0uMfU3FWzCcLbFR/DgUdrfcVNKeqK+n
zqG4Kc0KjnzOLJY3muQySAFSj00RV31VlDkkROmw+liH8En05SfAhjYsCs1K
3XZFbUmjiRh440uDQ2JlkRvjbb8s8tranR+XkiZTO4V292RjT9JFTHNvyym8
b8BZxzu6ZioeAOmarsWvNVBNxBexv0GOhJ4TuSVYLJH2T2xwwrYpwuV4gdrp
graf84Idk4TNsrMSMzL6nN64sWlRUO8URYybzrOrzNKtRgU75mATOWKKktU5
DojgKUMYxCLPYDhXmF0momnp2QBPYgCZMsVtwdWolWfPh1ylV+kpsbxrsG/h
PDKeC28AQKi83P1yqGwjMhk798brV6rb3d5SMp6cTUeDTi7KiFmb1joEyPZF
iVuMxVO1WkZcnvPZa1SvNwt+gj/2fcbUkM/PwoeLJUtyJ17+5lXEMM34D0pF
IGjlsJNcM563KsQZSn26XVbGErJc8JFsUnbHXnWAn6WZN+c8DoVYuvr4tDvS
nE4aUoTZoeE3JYoetAMKdtV9B14QSpn2akYITWxkVt5Y+NmxQAEq1F0glf66
VsH52IGXcRFLUyohWBPAJdvUgkLVP2Dfbe/RA91DKbltYbZ1KQWvqn9yXVoM
winmScBPHG7RVKfjo6B8q7WdBrXwgzX0BwIxDxy6eNDW8yBELKJnjlmRiERX
4Ve14fsP35KTG/96klpvhyd1FwGLsqOnrrHbe3qvEuMmtznVQnW6tUlohrSM
1OaxrapuivYJeMlY3AH/y/FtVVOnr9EJO8LgicfaNkLtaAA26oa7tkdG0kjF
BnzgBW8s2VfdeuqIVUwUi4/3URAyfNPVDxU+cye5aV4IALVB+8Q0kjBa74TP
E1ImRoJaonBsm5TtNk+mr1hw0VgGLio9jDtBuDXLNgTLE4orGKcnrf4IK40e
eTRCoGfadso5MQHxd/KG7RALjqQ9ImFXLVcycModNoGV0LJr/5Jhw7S9EQ8V
zIYAjOUOl5Yso8bQCCpJg09i1+1cfLaHg+fOxDuZ1pPjp9Jon8Aif7uil9NS
39ils2q4NBtrp513JaV1DC+vamAJTK4XdgIZvuUmo0imQEN445iVKHdLCn3U
N52VVszYbTXVG44d/hJvVSJriByAr0nr57rZMWWZ/i5kxwAuNSup6RxTipTp
driVrIOmHts9b8B29lzl2+NxoQtddILIFdNBt085qQcnY2mgVPsZcvXHB585
nKbaIP7/Dtf4glSMz2oNwcR6mzVjBy3vmmjO9OCr0vxWoJCVCWwxxuh5YHTS
6J9iD612bWLMkFDkkO/oHJ364THyUK7weEW8AoIUfSPMTigOmUuik2esHv15
46CClVfLCkhB72w00EPozL08RLjptZ5mmi/X/X75bgMRNrxu6xoedUl4x6Hr
i4OsylHNuF/H3DacmvO8LzxLwdYFZofF7rEwOdQi7ST1tQMu4qMfMCUxRGMv
6ie7Lz9M3Vw/1auPVpfUJ+idZhjjesObRpgMd5VrEhqwNUlKWxTaY0qwjZIL
fT6FV/NzPBWPC1pXGcjwwhC761cvb7gEMuiHhSpSrZusedsddxq8qR3lDU/e
id+1MCE/8GZOQ7h5HwlhsJf4NrlNFyYIqUTM21de0UcVZEDLyRnmryxxmrJU
Jc4HakQ9BYC7yjDPweoaAC9LGSlGbZnde7IT0P5VeSXOg92Ba4F4pR9/UQzn
66+WhU8nfOcXC2PXhTPmoFzE0BSCHHPsoj1NNZ0SfRilHyMOOmKI39a3Arvg
ZXPgQBFt519enBxY9K6t/uiP095Kk+rZmjpRLioPSzFk7PUU60cNr0olgqui
LAD3j2C2uQc7yDYGPPhD5izqMy31xW76NY9dNBhQ1GpjscKtN12R9iQMm78M
GhzNiXO/9okDQcTLhhnZaG6o21cA+6ud1okYIqIyUyLi3MGZTbovuqioJMaI
t8n/PUojqpzDfjfNyXLt/Cqj6xSsrGMEm1GV8+xSnjdTRItgW5MKsCQx3Eep
0xU5+n/BTL3ijpUrsGAonJzpPismcAGwVxW0GEJa0TtEFHWhDUk9SrTPWaxK
7Pra8hN4vMaGu3b9lrRGLhXtaV17qWYUiJQhIz1KloEBh5HoSyoWGt++Fm/o
diCr0TZAM7FvcyXyaa4EMBEuCCM4pCygZd1aVIw4zR/RVqZFChNPDuyV+lih
s7H5MOqtOhsFsUM30kRVxoASRve2XucWRC0GQ+ejBj4L84O+9V9YJFlF+Pgh
EC2bgRRmqmzhZBcGnHrwR19gNc1RiEBqUzjBxVxsdD2DRig/ZJgjfoCTCXUv
9betZ3fbxxqig6/FWdE/Ga2vhArqMgKAga7PTAcFpP9JXax0Y5rkUq8vIWEN
BTRoG+WCD+lPGVUWHKnWj30+1KWgFWyyuzcow9upHpTRIeka13k7bM+wE0Qo
uAx5lBSyVkBvEUoAqIRm2m2LtdEkRDpjbDdPIsaZw9+dJYu8VNxOBz1Q5ARb
4jWWR5PjsOb+n3Wg04pzppDqpWCGIV0ijBLsLlvAzwItXRptf7Jvk81p1flh
VZ/7z5E4O9MAWuB7LeXggZgESo0acN7LRXhcsHKe7KTBT8CMmZ9mXgBJFWTA
/RzTrL6jfjw+RvA7FezCYkToDxjpCNNZxADFLrVvIubaBme9mQPE/b/q0CYj
GEnJ+4LLCMlDS2kuqJFub3NAEpBUo96NUIy8WgLqIOig53gJs6DzCqtzF3b5
o6oLFfZVL3uN4LWWCVvxIWKoaYb/R3YsckPKpOyydRdgXRnPNOEUR6AKyNZY
oZqbwW/h79eVSB7t12EZPsrOhuMnBJ3lbZfri8yqcrcmkLI329LLk7/5x/2l
ZIFkosSMLzA4utzn1VBHB/sI2zepjP9AUDQR5j5ntKeCmS92ixLvhxJ+O5Xt
mmztSdGD3x7y3xbAl9YrgfVJz0xUCESC4IX8rfpuH7PMU4S4SsoGvul0qZ3Q
XbnV8yK+FPzo8Aci+OD957vECK44R+0HixHj83NBvihK8hQigafUBq3bKDd5
bdkIARfpsk6XcA+I1gGqkdCeXy01LCG8jwM6yE3g5GDOb4WKYpYBCIk90OnV
dtF8fWTAwzU2Y1s0yf/ivyVCXyT66y3Gd8dXkBXmsyUibB2yQoFMhhx4CJkE
MUHTv+kaRyGmVIpVUri2kMyJ/q9dS6leDwf3lYsYObaSMhwA34otvCYW4oXk
WRLalygOGHG6rGgaf2TY/DSha/V4Z1nn3c2KAI2xzbfDrAZnL2rktCH7R/Ix
OLhtK3D7h5rJziv469grVm6pe5FuZkFZBiSBDYTIiSgwXEMf6cKpj08NPiID
im6thOtPglSjjpb3N+mOCqyQevhQFZrXkcRy+kw246Vk3I306HWSdpe++bwj
GR1xCfqCmVx1Dqjja9ODlNlek+0kU1tzdFIpMqVRM4D/aVubCVYziZZcLhUb
9I90Pvk4gZOYnSHzYN4I0ggXYgEDGQ5Ji2GX8kfQJIL/w5U58fSpRhHPUkLu
qq++oGqYV8DEeYy4xehBa7SbMpJJK84dqeVA8vIoSU1hpUOn5dhptaF2AbwP
Whudassuej8V2rJMF7T0SoXFKw0re/h/J9JDLLDqXvrC9ZRQMlKESMrCS4gO
ka+p8n7cYj0l5njg8pQDgfuYU2TS0OpFGvdCdltpuUs+MOdhi735434yASY7
bXdddt7B0r/PTFAwmx9JLND8ArwjvX7Tp1h4RZfB9xxzACBpSlYtfkCdc4TY
3uClv9dv8x8Aneb96lKuLosjx8M9xuNXOyYXKck78bkWuOw/bYCGME5xCdFE
IQbRC0Vwo0+y+27FmhGBXvDnVzSb+dSgi2RZPkG7WQouSd8bWFzXvQwtDBrT
e8fmZ0Fxzm6piRAxtAMHPyad8TWbPFtXooqK230jJUIHmWANiLWWqUUAp5DO
LD6TyA8FDQkJxlhb9CQtoFRKk8CCvKF6h/Lc4wAwYHgf8x136FdctF4wincR
inXQOjerPHClwXkPluKFh8FxgrVNtttZ+LwYfIufqFz28XIAsCUCktZ0YFii
9yn8YFmRqOw7qIItZ+T6u1Ptc/x/rihDbTAqQyrj8UPnIjXzexResfydGWJl
AAhb+7/QguIKUQfYgrsS/JRHx4WQG7jV2sUyXx0n73SbiLrYBmr4RZCVyUsW
8/Z30MjKRAQfpa+ct+Vlpu3r13GBtxiLWRhZy5XDTyIMR4xLj6Rv4WyMGCM6
KXdvv4lPEDo5J8tomX1mMFLE3n1O+kXyMAWRFrprjTX/yvfgm5O17li99dhL
EJGD6X6xAV+675gc1n6wcOVYykrumycotIkER1Zgdsy/BsK61P9CYK4jrCWe
QAw5SLnBGaIG9JF/SAMaaiyapjggLuxmpUJwuSSjSJT9oPQUj2ij+m6/PwEF
otOts5VebXR78fnq2zNO98PIKiS96dTHuC7Yu3myunvt8+C7+XDmIsB+sybZ
bcFzKthj0pBjVAiFUQFtxiF4pr247MOwWufnvc2sYRkpYQ6vhx4wt/gDiU5j
w6u6p3pe1mnT0Wxf/yHa9YEX6/ldD8kP8q5aZSQ/y97XLaeA5EV+Yb4QQNOy
k7TvDInQQv9DIj8d5g1XWab9J1f4vvHUD2zke95l5yygMIuXJE2G7SSooYCY
Gn7/gXUptHssZWoz12+xVPdxnSMr9KF8W9w8gfSPEs6pRobTeDGm5PloTE0s
xqngvs3K0j2rCwbR/zJqx0nEoo73T6fNjfPTWQ33uEZbepZVQHvAHHD7mPKw
KFvXR5TUOiE09NAnah2MPVx9DIablML4R/L6+4uI6J1F3QY4650GejdWtOLk
rqW8RyXxbMYLmar3dw19Zyoe1xIK14QEg7r84dHmhkeU7NDXW0gtJ3bGcnBp
faK0QxtNuFNATS0TdPLubGEX5J+xa9ihcEkgWiOi58dyiXgU1QwxyE3hlrNB
RltapQsNnMlh83yK2jwTfZUZdGIMzzxzn4c7uSJyovhf0pLSZGJeIqcV6cP2
Y31MtTs/VTb0nrVRlBbKGY45O6GJY7LKNKy713MVY0BN91KajNkGyNK6jcIP
a+c9Sulg8+s53AeN8EbOJtWFGdq+58gxVttNjUVBVHf+NQYbCtsOG5degyTV
3wvwSlCIXMnsOnqCzq5hf6va6NYPwgg1xIPGIAkzhZHlTgH/J3SdwZO1L/jJ
s6GHJqU7y2zkU4cjUieC6ZmbBlx8hkL4nWnRzI/WOJggPjzqxfgdCbd4q/rG
ms9i3Dhf5YrQo8CIupthQDappKfhrggCQdCezGsTjRNUBMHv99AwxC486jBP
Y/7IqJiC7v7tNbcuzdaQAyavhR5abG3pKNh7KkEyiKXjXhu7Dj8s3WUD3qkM
paFMUHe8R1JmVQ7h5lCAm3ekQJicAMJLf3odgub3asHJQFutnZs1R1Kvzs2n
rHF8Osa7znpFujFfZ3Yma6Az7oLoWEaqyUcljrZb/4y9VcnraOLZWpy8XTb5
BIhttHhKuE31bf6Yf4RnhzIeeMNGcOoU0xrqAdxGjXLjcZ6qY7Ex43LeZtfn
AK4NJ72OHYYqOTnLMnkSVJSUGNtYWs1UW7gHAX3uF+mp+3DhO50eorKZ76W+
akFvsdHUDNJ+wWZ1JN8J1+3bWVnvCSg1rq4Rte3EFjv4ZCeDy8siZ2LhB4vs
8+bEs6uWumu3RYkN90qxz4eABbVA2saFUJDlTrFP0l7dGxty3ce3ucNw1Rk9
RmTE+ltOuPRCt0nJS1zd/CS8pKxf0kXn8397VXSFqX165mFNbav6kKJS5hVw
t4xg9pXJRKynXUdGNLZy1vLpU7dHStt9miVO+E98b70WzUrHSxDNXpOVKVNy
VK5GOJ2qNHtlBZgXeMuRN9+oA/zf3Ygtdd4evjVCQFaNit4RjXsck8BloKJC
ctt/ZmwL52ejNzZn9p38Qf/LvsNuLUFxG/sPVFXPeWGr4hlI/AZbe7xq0zlf
xOHjrTNCI7x0RX64NroJFhfZiulLJOgOhL3QzDJ6EV8DdJ7Co0uEAUxr5c18
CYQ2gU8nt7iHADtaklJR2b/UNq5NRNI6BS6BAnj1E8eHQdWkZQI9gTJWHXNg
vP2OmlnjG9c3mAIL18ENFwpHHMeqUXVB6w2xOgAOCC6IwKGOnFyN+GUIy1il
Aynm/Zol6E2Kiudmoe/SMzR/nP2aJTLS8WloVtoAGzn7wncfL3G4bGTL7p4X
vAQzNRPU5W+kltgEeAxdsfN3e245ig32u3vMzw3fQrapoUoaoVVB/Kf0rucj
GK4lZIEzQ9as73nvcsPBMcfDMiG+Mkw8krICI/Fl/YirEP9imwqn7JdsZzYJ
7XVXa7H8Oiho3UQZJQQ0O3vSdmlm8gG5tIo5J1oARFAHMUeC3+8fETzr9P+E
l/2UbqvfWYSAdTdPEVu2LR300STWN+Q5CeshkVwTUpw6nBELQuczwoXVPjtq
QpaEM+slymKc/rS11GHNKAqGSpCRkb013NeanG1zHrOIY+HsjgB3t6tYrTql
dgCl0vZEhTkJ960O/SV7EfH31fUQneEpA2ckofpZBlwxz2VbJ6zGXMLcprZQ
JPqP4Rf3UUaO7rwH9XcnG3O6Ebz6edkR+nANImyvsbp5m1AbrRBslUdqTB0k
8GVFfiCrZiI/Pxx52hYBN8eRZADIZTlDGziSbUzBuJQXwA+8fmXSi9YB3hqQ
SZPV047U+Qbb4VjfXIyYqQszs0czbiobsEt0SvUWJwMngyHXp7csgZWkt+rx
nZI/vzeaBgn5N2PRc+XWzxEJ1DJ8StP528SJi0UrbZprHf+Oq+/rYghA3a+w
WFi/dukG/m0kmHnxeKJHd3jn9to9IDxSnAJdbbgg9L2cZM2Xhuw07jlOSiAW
X/EjwjHurS/VB+GiHy09ItNt0S17ZaWykZtBZrTqnbbVjxg+EWb0mBm6R0Ar
OASzQG46lVdyS8qFcp+J5Q9MpmKdc0aSqH2zpqNZVkYjfa/r8II0GAFrxtef
0RW3v3rLh2ILAhV13HEsYgXADqXo+BpfCpCgiCk+JocZjB/Y51vcDJ723Bf/
man0ZCsoYl1Wl79LbFEqKdlMXpgCFoSKW4BpIkL0dPs6lGvpO9K4x6KItj+G
dtG78ceRoe1XJiLIo+gTggmnz7Llen6TyqAfFNaoS9UIfZTSV4Khq9xXOXjo
GWGh+DTvHyyT5Z6dEKO5zoQdaAj0Ecrf3Ed+4HoqQeOt6J7PLCH2YwyZH8P/
cVFIle8yGcd2oUUuj69ebdxVdkVY4U9etuVKmdRKC8ubmGDZ5ORlbTPzdPXR
gS5lFTMmz/eCWIhs1t/oTxo0mCct+95qYJXWjPSmYKYDJV5ufdCynHtr5zlz
BDz5H4NkgVd32vWofFPW1kKl5xmPWfHV7ZNxRHML/t1uMYLPVaORtBnPQHCk
iwVD3v1G7yyNyekh0HGxxYGsSRrfcPML58SQShUwN5VIJRrRr7Nb8AWH7mZ0
xlzxJekqxTaNtoNCapG8Pp3U58Bm46pb9cIKPyuiDnxskvpyFb5flLjZ/lfT
/JQSwio1VAzxG9lEJ6LVpCxEzdzqloFqLM8rZzyZyPsdVL0s6NzBIwUhkKzn
HJSB3GR8a/vhJkcFE/S/VSVza7+AC1Ld6bpJtVc8rjhaKd1kRCfLf/WZZDwa
A6iPMbd/n/IMlMyUAmtZvh7FKL86Pp7iQE4bjUK0ciD8sYU6bLqYYh8MH5dt
31agyrF+kPw/TzEg+K546yuQLoViNsAdIRAaSj5jmvNg/1ytYZtu6DTBpohm
7/6V4QIVDIaUQP0pzor6LbQ+4y6j3/7xr0xwdkLf1DtEdqf1VCqDcMUVGdWx
vHAv0R2OeYsyoYMOZbG+63XHH+BlnlxvjVOa//N1FcVADC6uaYTENOU/Mjdl
FkxTE9HpxMjN75NdDOOGpHmWd764v4UVVoKiUly1rAN/xkSDpm0yq6r8/rYc
ssZIh9OSORWic/F5SVh0CLK81y0UsJmlHlZpCU5OduvEWJoePzDk+xAIAgo5
XanF2JAnTErrocINlvj/0AY6/q+xY4lWXmFoNDd8qO1nz5KqgqZPrK/vsKdJ
Eagrd1grfSi5IYvCVTL3n1QTkfMaON7UoAGqaTZDuS+vs+MMUTliZFlQQVOd
RPzQuwGdNS2Bm3YLiAcG4uepPHs8Ox2fRho31FnkEU3JGv3K84fbqSIPtclt
4uGQlqhCZ/C8CT8iWAve3XXVctFPPm7HS7pQT3rwLo+/KN+gZD/Chu/bFPhj
3SwMXO9yDKLhY6MA82ZbitsjWjoxw8fnYJfMPRweXl3lPFc7vNIlQ9CdPz1I
zRJjJj9Uqw+xC6NCcPdj4kvVsAt3tY0wvgoYUUXAFG0d9oWdcUvp8MHV3R9U
GYoAKrw3IzcbLlbcILOTxVjKB+6eX0Nuq5XbPpqAtJ3UEueNqvKmmYpae/T1
uAsTbATxZeVsgqZoC5pEuN+UTvzW2hDIT+zLMVo8mQIj9xp8Gu4ikRnIGFDx
OSFITS7+6ooEqXCpYajulefh28XfnYXulEIZfaeHge7QIYpEd1WYUCb2CSwl
+Oiny6XGOCvF18m+WrtxpZMFkU+oouzj+gnodB8mWfzNQqkQZix4dYHzxfes
J5C33NMYQ8WCuCeqjxtGEt/hqApZnMjAVsNmNSCkQ5tAkpiUuUS1QO2em4z/
qazQoBiO+LXxQSikQkFz3DFtKn6XECBA0N/AlQDBEGcm8teiTDju9AWae6uY
s9bUvQPOek5IjzDI0WO/LP4Dud2TWGukURBODfpUg9G80lOohcuPRff84mAJ
rm6oqDK7tnpVGqEcGLVkBCf0+GSwGphDZ+VRSOQ9tRfT9I+uLbp7i7OPzF5L
hmuxQSMakZhynYGQIO05j6FW2YeWiQs/XYHpMpdnXJuSc4ketRIC9Ng5l9W+
5p747pGg9ADN9PYF9Hmw4PEpfoX0HqNqkWyqyW3zFBnUxQBBd2Pw01MQ1ixM
nBNGrRKR3vsm4Eg3DjByzJUiYV6TqDsJipW0ts8hdEH0yX0Ub6d08gbnkYAJ
f7omWqpE1WaRLzYT1qb01+8Pi5rT3KGn7ug5NiFQ1eBSoH5ZDwWaIBx5VZ8s
+AarUPmgIS9EL1Vjk2hNn7vVDTSCXqhd1VDpEbcqETlKL1CJNriS9qUkS0iu
t0qO8Apw9CiMyYCM9LLxRhKr+VTRLRHFmZxLyqXMhRwDzSF0wXFgcZmhdK/6
ZQZws/KaXCOasRe1uyaW5tOfAi0CBQABSAcJmGxYCa3VUEe1wzmfLohvveaN
0GU8+zdHaBOmzXYUbg8kQjnT/HobNBRJ74sgR2PUjeRKK2z0BSxqJQItPTMB
eWs0AJIwCnibBSgMy8VnV77J/SAVw9f2HESidDtGFQmt/9rzIPWLPCSYBgjX
loRuyJtOR1UgAFzQRCuok62+oeqX6WYXIbAgacUTOwp3ohSbvEomSfVbgLNn
GOeWDsa2f3ZAmgZD7nine644dSUGlRlKlptHwBGYbg2HRCwjkgE5FVZadh8c
PLkjYaGDuuIky2ZPnb4x5M0somsSGFI++x1CKGb/l++boapMvGxhl1vQX55p
aMXDhAHADvUgU4bGhMJgJN/YdlWHJ+ss6XNGkJIObKJhP6rTnYDYQh/ICz52
i3fN5TA35WXFM4k8zR7EwMgutIGRE6hK7q12+NrEvVKNtfASJ/9hbjCGzVp/
UfcWugyd1gIusQrvimb5Y/TGd9+HAnV5xWRq+BXNEbKqG33b1XNUHSxJ1DBj
3IkYC+okYGFurUA5ZtsTIWNYNPRn8TUCj/M9R9ziKJYnrfkdzFr+/HZoQrin
N2aloKiF9wXvYqTzNHRA8OCFrVzhk3T+4GZ4XDRYxfPX3pPztmvIsixfN/5V
9MZgz6oav1lf5S+oZIEsd1J9B2YEPZRl1U6CoI/rmjbH+bNk08NRNBciGe/y
l1CUcjGMOlNYadUyB8cymfLftuaoTBemF26uvwfISGhf0r4RDT6d9iixQHie
Znb8gOI03M/iqhUzo25V6KAPUBWJfLioZk+pgTAdqg/OyWrlFiFweVGg3yL6
0mVDAaS/PX9rSn1ZpW96fWBx6eg+/YuMPOmuNQ926+08KbTXYuer+AvS/MId
qBGWXfrwgel7pjtXDnt18/a5fHdxWgjC8Lwk9jgwkzzUP4dxCOjCp4/WPlPA
j0UV36Tce2K4uo/ydoLw1gim13vjIwHE+5wi1PZiiYXq2wsj57Gg7rkgfrlQ
STtJNeSSJ+xxsEVi/lYyYM5NOT7ImQL6bN8OFjzpobDVi3/Stk10lzAkPivD
0K8IjDvlPKBYmkKEsaS4N4FH1uJ6h2GTWxfCSlLRlSave/sUjbMgH2Nua6EO
d2QKbkN2ZfZbUTSvzxsMDaSTKJGj5Gr2Pspc9A96Y1H7dEAu0bj/3iNlOnM2
i4qeAUzwrIy9PnicGn2R1lsd7Pv1pX6YYmJ73lK8siLxO7F6xtESxTyBo6FC
m2mw/bIgEz0ElrjQQ06hCtWV0MLjXzR4tmsqb/MKD/EXynanNp+v8TiO17bf
mXGSt6VsGJnVdCCr8FH2HPavviCeLQMwkvixuPQB4JX1iTGYElDsetcfacqj
+XKgJcVnVAcuG56kN+9jyVnOXihKRYLU5l7vJ3g8TNc7yEL3rBtr3ldxm+S2
tGnJH8oyWWro6lse6Ss6xWkUqfz22cOJZSL9aySV607toB+ScIyvhwjLJVm7
9TE/CSoQVgopxzfhKf5gndiPV+NCam89e84IBsP4lCAJpTAYDKFGgMXzMiH0
LHuL6PMrIOkFHj0BG9keRs12NavPnCeupYu2VVFRjusPzigSypB1ESfXUuoq
dgXrj1JIh7SbmxDRW4IwvI7PkkrVTErwRs2GfySuCzKFH0R1lP1WyyhpRkcI
ruZa6/mwWkBaCWCk1ZXiX7rg0nQRPvEb7tFJteRgQEXUKY0TkNzAZyr2Y+no
tCdez9NC7wOkW4W8JlUwWxAnhba9KdLQu2RoJlJBy8SCoPFMBKkuwZIVIoYn
wVmVNoHSrS2NUyijkJ8kKvLujXrbktEoQ/2xlRX2NmvILPgdi9QdcoM9QUjG
yokn5PJhEF8TRoSE/kaUqVul3CBlzFEkQ01J2xL8AmAnyYcejzbkDmlwHNLx
jfiQ1c2jduZSBH1UNlHbLop2rkbpLzR1DVLvefmsVYPxsc4jdV8FTFszIOPI
1gO9hdHmiMLHoXqfWm617x00whSecZtAUjT5ZrT2uyS8D6ztZsaP6UVdkdpl
edATUY+K4T48U707hXMvA8cNmOoI8Fhkac2jQHNuu/lIWhU8Vy8k1nl5ncHu
6jXWfETLaAvxxc6BQ0OqmcXQv5YcgYu5oUysUPdPbe3MLuhm5VqqSA3qWnxk
1kPaAViOnSCyxtQdyPOKENfHg/ufyatMIR49KvUfHzAGOpbhrVsTJ1jeHCrQ
+3yc5PaMOshkg4KBCGvNkytZ8XxqSbVfM3VMxcoZjame4CBz36hYWGEisbGz
d+9YWFkwp8sHBHe1UQUdMEw9ArgASknUY5b3MS+uCI5WYxyFaE71Lm1eI6hF
Ewa3Ml5/rPlL48MNZY6mQ1vOTn4YW77K7tiLEWbTAqmb8F4tTTb7gsFUeF9J
7Pxbt8mkx4uxyIvGJbxwFhIe1Uh0FnZ2Yq2hxvijIY8X76wr4HkrXMboBtN/
OhY8R0b8fxh572aLkvijq8amTeFxa5uqddyZWXU1w6uQzjrWdC1eWT8Ds/bM
hgBZcw1vR43InU1BcoOBKFByHUAfKWJA2zvBsD/m4KU/+cEMaJ0kEQD6NoW1
UYCtCJ+Q0oK81z3bouH6UloDzdNXbsn8DyqAOFEH5V8yNxuKE0JRwNhj5rZQ
k5SSV8NH3oHgKmHbASzIEXFkMBCM2bJlHUCrtGqa1zLkg61L0c65CjDNuQrH
qU1+ZXQPmZ6s7h0ka1611awMMMo3EoUCKt2Io7GDd+FisA3/XXmGUXA8DCpT
NGUURO8CcvDPpdsfGzpiOT3QxdhKg5w3IlamotUEmKrlepQvJQNnAIBGE3fx
zMZl0SgGbGyIamjo++gCz3MkxyL1PymIIMhEQqCNkqiTN9khfNpbeccJmY97
7iXV6NkS+x4uI2wRsPTCOa55LEXylXt/WfeCdbGLr2dnHVKEnNGRvCl/Qm27
eo6QmFbWNKrGzKLlWiiKkHomAooetRjySiLYHdcvGMJ2FP42KnI+mkzbaec5
vBXr0ayqUWQM9qEdfL7pt7jp7wnZhHNX5+YtGvSuR6eWWxnyhFztNw54tbXI
O3KOMyRgCgJ1VS53CymZPIP9HrZ2xF3V+kTWXnaJV/pbLjhOVen9vU+2UD9L
lCtdhXPW9lVWa9beeVTBwrVy/tMXKDLRYkNveCwoTrDywF9NP+sdFYPAeHNo
UHgblPPSTfwJaHbFvoB+5tHgILZrNUGIttfVa0eXNUCy5jiqUJuv3w5s9KsH
eLs9/dvdNl85aGyvU5cwnvwKuGRbZvwqYv1nf4aonQ9JGSKkKr9auKnd7Zgy
19KF1KUS/FyfHvMO/zdkBy+K6j42AP3Aq2a8EcVhCj1pN172eETl58oFHdsG
P50oJSSB5bSdZ7v3uhR66K+gWdkm6wCNa8Y6uU02MDxNLTXqEtc4By8eDhYK
WQNLgjf6OmmKiAyfxKC5jENJjUmXv7sE0aqWQ4mQI5+QTdbxmCj60JVenrDT
j+PvBBxnHEDNnjhuGuqbFB9ccLB4Filepe+2WXsGBKLsepS6YjLJ5z8pXtn+
ZW+mnGSIxRmBWQsIofgXBaIUzB/MW9URV7eW35rPP2v6qC79jePg3LiI/c92
eiTGlZTTVV1naobCzi+b697F9LbWCg7AtpBkitCc/iaoQ1YX94H/qpdJ0NFy
sxjh50VJOmX08PhCNOsCT2STusmdYf/jNEPNEKdBKajyfXjTfDKumLobJ83L
VITUPFOFatD8sex/EaD0SJBntIEy44Qjc5btQEKVWrcGC/VnXzmRvsQneP7v
JxFAe35rm+InRD4I1U7VXzhT7SnbKfEaZrfBxKTM85VnNMig8Mh9DlYfc2Uo
EtMgjoniboV65YXPbpcZcqo54NeYb2cVNVsHdXlr5L0AjOsGcqET+I/LwYEo
4CxBGWrm/wDcioX5E1lOKqzQ0hWVJj0P6w03n3JelrZRk2CqvcIqMYHqq+11
21J9NwqCKn8OPhEijxuMu5EpmOwxx16hXOkzwtyHBrFhMJYewCUV7FqCiyJj
+7fcpPK1BcMy21CAddo3JK5Jg+gCtfHO0+rYPm+QyasNhKJn6ZyyQRj+954e
0ZpZdlrCWAPtiiHiWILcqMxAbixocq0I7bpDjDSyg6fRNMGa0vJWRnW50zYw
krRogY8XtgUmbbiUBJVsi5YliPH1dqXgGd8foVHu6YF5GhYyAhCpZEh5CKJO
5oK9ivEY1ZuzXvalhQKNajhLWDyDuxRhL9VqW3jxF8iSUvM2hDSmfA3mViZN
MBuIRGnoy2qM87M5uUUROV3ksdUoTamjbTt9cO0U6vAt85XGySA1Zwbic0iv
HndjLYQ6W26pgY2L20JE/1YPjDZErUcPeHR89EmqE5fQ61is32kgxZumiJUU
ezdgyFRzCOw8A7Jr5fRTiJp66THMFq6RlFP/NMjR/UrHtdwoFn58LOyUKHS3
dArEWcQi9qLItvjBfK5m8zROzFLFNPPGCFK/5lyqy/3PCyP00OdHSaBN9MHk
w3WU7kuXWlmKCGgcQf9JsTs2YYSBt35x4ElFPqSzb1WZrd+XKZBz1R6zhqZc
i4femq/cz44Fy+zdNC+PYC8ukg7f4oarmt1FTK3uzbI2fVG4sCr7xPPLjUDR
lBat6z4DsJ835v12AxbgT5VjLxOmyFKL636Um7KltOR0eyAyl7M9e1V3qR/W
mQsgS25aWyr0wxEs+qAxhTD0lUyDxQaRzc2JfLwhWWILmsgNwWi4mTc7xnL8
VYIKV2KTsZLkllgvbWilxKQcg0E8w2zH2u6xMCbgFMRLH6EnRZJnDDWDdP9s
b+fEnoIaIL4H1aFpRcxV86TDAuGErqJJPxyC1O/QfX7sY2u6dvbNwD5FR1F8
IwJ6nnc8vzn7Lo2TzJXHrTouoCbzQRKL0hZ7ZbiClllO/A8YO/Q4sGGU54qc
a2DU/pzaZHebzDeKkbmy/CmYHgI9wTvKU7/CFou+SR6nqACfYSBgmKMVS4NH
HhvE/m2ZB8G5NPCtnwEQQxmZGVxLxadPnsjEeg9LdO759V/vRSR1YcRDGMN7
xsFr+iQZjJbQfi2+Jh+oQO6KvISQGOghMoaqOZXeKg0WuDMcOa2CDgJQhZIc
BcdDvpPUr9j64OL+GsQKGQ5sI2MhtUDJKsA9/CAmCgimq5b2b27UrDikicoS
wl4wzhODQB+OoQXcoJTxad52Jr6jtQsCwX/gPjIhQyM3EX6E3aDm6dO84af+
+1jCQMascoQTdwN6oZh/BACLsE5aSkufim56qYL0CNewHHWSyAvABxVfIWLT
hBMlpQLGVnuDXRiArG16yJ4YFq6oRziQbVJaxSCYtGyYo6ivBkiJXvUMlZcS
QEiQg24dBLLiepzvpqilLaxxea4OACVfhyuTRKP9+nXEs5Hq5yHwtNcP4n1z
o25SQVFPWYliPS/EGWl3R8JII8OfWu59hho5oII3YzsKKvoF64RkY6/xJpcE
triDQn2DV44sU8ng5smSJkTc0kZ6Kgo90giwGtSEj1582Qkx4/CzjzO2AP85
j+UTXRCDZO90pOyHkGXsYISBH+E3Am2RDLQ0nNzJQnLPBqNm2lIFH8tALn6m
BaY7g0BRmsLZkBV1dIAIpWkqyUERtz8I8uuW4T7qNNDpwT4J9mMaDDZqmXtn
GyjqpE4NB1jNEUH3ebYxrvo0asl54/cL+8VJ68hAlRG5Pw5SsS8pwm4RgMh3
xmVc6jrs0Px/k+5TZaLOQSVatIlEPOA8eZc0/FLwUavE6CVeuVAh2cIVnCOI
Nc7NJ5FLZJQ30IX3Yj1IqaeSoPO+DkuNdjtc36aJbgC9HE+slMSrDYHmStGr
hzl39bgGg1QPGQOHgrRETF7WnpVx0Pdi4Xl8lJimv0oZTihbDh3TRFXFV8M5
rJf+W6BIOA9v7//Y0zt7KXunSHsuELEbSDChvPuqrJ9aFNqr2ArgHcFRB6au
J38JdUrFj9uYCLvUbdTo8xIkIhA3nNnphQOtqQuc07I+tIv7ARXzSDbl19Og
EgEkHo4RFxwmoWKc7XE2nr9yVEklHZB6vToNoAHzTq47XB7v9I6htvk+KzlQ
0uApELmISlej/AqGQz4YDYZd9LwhNFct1NM00X5owL6vDiXjL5+U/5Tcuw/W
3N4zKWghoRGgrewE9TxicaFMz+oAB3KsWsE2rnT7es2VXoWT0tsZ5EPChOZh
7KVPJUu+chu1u40eT/M7PJPl2ag3sCe+jT5e+br2kj78SofSFPdIYuKiERTG
cy9sRntswmPZJjtcsHf6MoFmOkBxWFb9ieHd2cgx+ofdYdjGHx5zWDXFia1I
aJoFq3H5gUKUoxCnr5lXIH3I4sL+T07pUy+p+I+PH9jyy5IuSjja9JbCufy8
mmFQY2WMpA+mFTsRbu1WY8YSXvg1EKt/SGuj16GwxuanRk0S/Mm7JU0OdhQN
ITM2pbVZAhkuVAbhOGXbgCeCAJsjJJHCj8Wp9vfA8JzVLT75KcAx7i/Ud+Cs
x4rguX/1d5sOQ0au/DAo+cZn9YQDalVrNnyhpUjUfEdNwPiBW7XqKZI+NawT
9cZx4076wOge19k/ohp2Fe7Iw99OtK7M5yWi7WteHkKGbRmiCVowLOi06/A0
XexewKmkSg2/1nZWl9Zg5NQKBHGhUWxVqUboK6rU+1DpNo7fqnaLzCfZK/GU
GcfeAE6bOTJqVpHiUY+I6N1Gzu01aDKiFLBK7VnET86rrum6Dsav+eNAWWeT
3DFLt+AGz3rV/LqTjDAVmOn9XBWh+Xuk1+9kqhUGyU/Dj+16oGYAEHgnFhzM
+/guMWoI/XNb/RTJ9U9xD/VlrT1VY1cfP6yKWfDlRowSKeGcmeGBIphOEreF
6oyJSuVWCcawY4LfMYcj07lMozoHgK/qKUCRGMo9d/IIGhVcipARSJPwaE18
fNy02mtbs/WF1e8bOxssl+NWvgySx2zQKg/XX+j93KG067xMWBBHvXC8abnV
6hwWeFFAmZ+kF8BGbGQc/l0c2nuBFJQpCnpbz3hkDRgqTTMiQLnpHb5hPxXe
077y8fHaU5g/PlKuiVsY+bLpRILr7wuX8EQXqy3xpvgVbeIq+tVo3aJ6rT/2
WobrFsbxGZPyBiQp7h0Et7cU2hmn6Wdk92VzU4NOMABOGktQv1VRcC0NEORl
f5E+EL0ZVC1FLZfzqyAHPIbzBMtzlrojWiA/VnqB/BPF9+DhWid12j0bKwFP
xOsaacNJ98KTB+toSgcbaOSSwx8If7kvPXYxb9rgYs75mCH9LmGaxLTh+esS
Z1HpHXGM4gNGZbWLU8s982vuaEBJ+YgUFhEVLQa5MNiRngFy+ehs2YSTYzbZ
/WhYuFFe7eSFDb5r0Sz3pbtSC2Jvs3KQkSqejA6jKhVKoG9tuCuAsZYL1XYY
/Ab3lcDWZbXS7oG+oBQcTnymIzMcbk6f5zt2u0NraHCyQZ1toZurotGMqJCN
FH/foLEMPgQkw494+TFw7GCkpzOxonHPcsB6XyS4ehsZIHDZwGMgnTvoNYr9
Q+HaCLsPNHqC5tkJX/qAfT5YTFB2LGc9C7kNtM6rLeHu+xZWwMJE1w1BKj11
qY19pKHgEGcezOTWX5uLpvPHOJsWxm2cyA0gR7jvrW/CM4xyMnHC8uI0Ta8h
+1cYlu9S6aUQ0qLwuj1FSDQJDIzlz/Ls2U0cOeMzj9tJFLmFl/jT/qa1GWpO
IwT2cn/fBY1BPlHLrAforQBxkPPC3ZnyfTOA02xUCN+O0QDGqSgou6VIafWu
xWZbsoF5lSWgIM07vww5C7zh4/GYVqZSL0EDKW/5HFpgxBADotKA7ETlq/SV
bhk58JRCiIRfV/5mlznLFS0K08ISjsBOdrCmHkAWL+rGMegQSYcqqYq0+HVf
t3Lj6u5tMf3tHSfeIJZhKFCAdwBjAVmEAcUgFL/YrkvWYOcz7XamIMfxpg6P
U49hnKnp9RRTjakZuFt7RcNfk89GEW72iovTXPw4clNqBVZ5z/NRm2KbOZKF
S9dv1+g6F4lYzUeX+7isg5PGVEsb9JpZX+dOiC4bSyckTI7u0yCBgOq9Nsm4
ppt42cE11cUGDSFoI/WprcZ7Z62xG+Hz4rlYkWkamOk8TUR4aHyT8tO/GAe+
RX/AlXiRzDNRt0xMdm3w7Q8EF2msbdQ3tQevwOTJpNfJN6cFg6GAVOw3lgPo
mmF1wkY5TWXU/HO0yU96KFXaL4n0tHvHDBNo59PAB3S3CPBrbDRqA0pHY7Pr
lx5ULFv86M/zUFXNTDPv0u8t8YPD8+c7YzjDBWo+thYUdZ8vS5A7I39pTrXu
pcmesu7RG+7AsM/ujYCC9tJcCYxqNjdHEsBdrqQFa3y0Fv0dsAjDpxYwG82i
MZg/1dBFi8cwVbe5jZHmzJ7h8qTDRr/cMcTBtPuUmqmcP+gg39ksfZvxuzaU
7tcHZrkaLxTIBLEFKNxksMj4D3aVujeGDq6yQBEVJqckwN0OmmhNazoiP+5s
ADT5xskjante4NdCSVccRPeFmpWadyBHpLfKiyVI7B25R6G8PuumUMGRtLta
uj2tJ3VmNlqrmJ9M1pRmP7MiAiOgg/WC6G3QNd1FjA8a6DvXeWRgk5z6Bl9j
MSdjnu3W8jQ2omvdezwrB/mCrkUyVX72s2HZL8kLiwdflvtT5mbs9OlV3iF0
KjsYGYbrJUH09oohl8qdsizHJ4U/utaDo78EC+l0hl8HGccpj1KDqJaFGHVW
5gTIXA8ZIQdsuG2IDecMPxmgjcJROw6n4RfGfPevO+j/D4j5bA2XNUZWuVxk
IvPpZmesZxjuo1O4zGo0Bp+rGSgjHMs7fZYLzBWYkDwqps8nHiW1k5k6QkDu
qJwf/43BXgoXZdvuOiAdu8V2OtU4mKI+P2EmxyXB3dBhwSk6aklnldkxrbOx
2gt3gt6qpj/WBJE++qf6jSDbP+64lPzffe682+m1bB1/1D7Z1FcyLC3G14Af
lxA0tPgUM4+WuV0j64yginpNnqxyRt2zTkcAgNsfXmJopL8HJMgPJnGS4nqi
Em4a0PB2gySmVxHZ4tQOlp90qzu77CRqGZHK7X3BusPyeMXe13LQg1ZEe+3O
WNbnPE7uanSsY/SvoEYuKmxuczjlhig3nfkwE35HQw3uAsntcfkN83doev6a
iqJ04dt0DEIWEB8vW0Wts9ZUbUe6g+bRcCAT7Vo7B4Lct2ZSg1HzVzZDUDIA
pgxb4FlB+hRlVy9Htk2fDtJZ01ksG7lKibYPUiq/KJwpzsiSZc2wP9HJHURg
vBlFACqeOigRIPDPs2sWPU1rnldvCUSali5ehjHfTF+ZCrmXk5G0SYvu2fJi
sd5o4g97Sgo9+9eNP1lr8Ocn52FEaeBGxyhXGYH8l9cqmeBgPYq+oFZN1W/L
uSSOJ1An0lADer0RlZVljwS8A6oYzlGRrRXNKLAquC9Ap6vk9L7MC2M3Inax
/cvzCN734NFNG0M8EDiYZamYiG1OmWvgwLKE/8N9qHVG+PcoyhUJa4pIDMJn
Ctgg3L21t3+TXAiBIKe/PNYBE8agywaLLJfQiXZTFgqw530j52W6jaO/EpF0
njg9hzQCn5BGqTBX2IVk5PuRwj58QudA68FPF9KKn20ddr695elb7fB1J9sM
pfkpB6FYDtpM5FnMPn7xiXHuATcmYwk8CNzdg8eZlzrewnAwSlwLGsxFoiuH
HHky+v6bFK33KPza9Z10y9Lf/1boQPY2amXC3JBQvp/nybuN4ufOHb4m6MWb
AMV4oLt5oUukyUX3/iABBndHBjYMNi11ztXSZIB/znL3iPkm8RWxuLxZaJNh
Y5GjLrzwR3rBb3jBYSvH8UR7wZZxDPjjqdy+Nj84/Ttp9821FInIhpb8YtVv
EpNo1HxAIt7a5pWtjXker+P/mf/64eb3WikBNSOZCLAIshsjQqfeuhlBazxO
HVzsKQkNDfp7+ySY0ZIn+Qsr6ZjkCLGFslMpgMejHAHaE8WNoDztyAJkvA8P
zenfvLWqcrAZ6XmVcFOBK9LOFWid28NqQr5BhrYzOqofad8rGqLcO2fbo6IT
Fv8XFSQxFD77GrK4dk6Kc6TjP+tSVjacTY4clNmt3IdI2zSO5Cga7MW3cSoJ
5YA0NWbQP3THA4cvbtHiLGFtDiE/ZAPlK8ImYLHgXhwcr/MCa9+3xlXN5Zvv
j/+ac7t8ygmqwdAY7yAczOAiQw9mf62cVvQ9fN+VMvkanLq+GWRBYoD1HKHm
CrgLm+AT25Z4S8fCLZrPMpD0uKRGlU91yCD1qeorNzzl8wqkVvnD34U8g8Vd
yhkluCeiw2wkv27bSJx9j3ww1udRXU/aqy2tgRPVT+yAe3KN1DMZDDK5+Vgt
722TkLx+5ZnBB/IXnkkv2StdfYTCLCNxY/41n7kmwW59O76XESoleT4RTPbi
2Q37kVDrafzzDi7kMxDTtQ0TfQxX8y3S3mLK8+MvB6k2pTCnQSpwlJ0Qvjw1
Acotfpm2wQjI2s9Vv0QJdQYeR+awhEtrgE2D8p3EtGhvLM4kAKteU+BM25dK
YrnmyI62cjTAYejVGysw3Aeezt3LGW+nFW67jIuIX472vPDNQeoCMv8uVmnp
mthRmxZ166f46Qa76fY5ZGqL3Nr8W1hD+5odq73B0JqN8pUdMTMnqFtHRkHn
kxUanZKoxi0D+BBgjbGJayyNkh7lTJj2WNSZ5MqYhcITwPUHjwCosaJnpLnV
yeVf8hULNKFngFYmYdu4gEal049nN70S3dF7RykVwTTnPhs2SopZtkOP8Tnh
S8oIQAfBwXjS5BsVYQH2GNEYFv2xyUrasbbIEutvMp/sE87yapWSYcZ6BSnS
yQHNkx5gdMbkqsEDngXE/6b9P2k7n6hDqLJgRxfpNxzYc1QEcXg/vsV4nRZq
JBQsfUND2TvENp1VK9N9+FgNdjm6pgQ1CWEl/NrYyaUBliuOYoDQ8NGdpoRK
D/GA/9gmYJsdNhqb6qyqmM3/H0T3sLQYv+5u/ofoHFdAdOW//AoA7YO55CMP
y1NfnWQyPnzZSFcj6aV53jHnwG8dDgBq2/sWXNjbpvHsFBaGvPIXao+HnVKk
gaDIEgkOln7kJXsbR3t4Km4jr5JHAEIZOOuPN0ZxysZwSFbQUg+VHgOWZoL2
7Q2fE7shXJ38Ac0WuUJIMryPTviF3xEbPOMgDe7VBoYjQcNx+Im5z36ipj47
uAHOjm9KoCFvwkDlb0OOlQCTJE3zjw88Edh2wqtmnC3z47Fx2u3hLcMVQ8xv
st1qoQe6zgzqGaUyNlMOb1HMcu5GyjwSU4eiNzGbf6pwWLSaPptic/lpITCD
WuF+w8GTOOEn4BTYHqkgWv5om5vdUa0QvQ/9ZPr57B6Os2Q/tJnCsgZFLpet
Ky/GRrNecSlI8JxMw3Zl9ASHcL5Jba+VnKtMuKvYZGvFGFhifzFajpASC0cY
fCJr9u4q7P4Bj5H0FreA3IytWuSPRMFWNlOZU96J5Y/8FKMJc7BgKdwBSiny
71xcoSYiAFE1ziS1hDgRaHsZFdtTDhvroASkt1vetLc5MrAef+pRK//cQLPl
3IuJzBqd/u/phxFbvOJPRo55BTlY2WMeIT7G05lfjXL1JjfDqzxb+sbslDr7
+dHS7wWrlyLe5fgCZPNWtpPX6Pw4XBBqMQf+DWlIbXX8CwVFA8ght7Nizo/Z
ucSmC6vY5KnVBEvT2cPiawZMX1ZbM7+7a4e+tGwJfxDiBlNuUGWbIQpvcKoP
LXxffDZnXEcwBD9B74t0zNtm6Cb6k+iFBNE+LrZGpd7esCGcuV3/ov4odpUk
wREgIFvmX57fm5342yRboD1OzHsrfSJBYzhB33zXL1j5zg4nSREOrSYj+kS8
2rOdORePwLVGvI34YtUb9j6LWHKicEOCC7XQumGO7eMUNR/pFyEnSW1pWN/4
2EmpRMyVZH31QByzS52PhhWha4GDwWwfyhYtECxV/ofR7kcDuVPJHrZpu0xy
n3LL6OoJl1Ks3WO7skzPXzY8lIQf0nwc6x5fILmq4wuP/cNRFvjBEeaKFP3Z
lXffN3KViuEGPLClpf3Jy2mmMf3bYJy7mVezHfd3x1an5crlvI8EE7G0n96h
CtBxhOgmkl/KzaS+EmNRVrS8Vg25PMGxVU9k82sfSsaORo8UJr937o8hQtWy
+2V28R0AclOumYNyrd/aaxj448ejwuI0XAkExScATQgqwj3MFalyBq26FV60
nY7bM5WwnTwrI3qDHgRQAkzWh7NanqZRbPK3lUsnen0fQeD03ESGr7ylp7Z8
pqNAvCD/38kI4jIu5avM9VKoByoaVNpPNrSiqTpaLrmsTebfSbkullg+RlIm
KwboGKeP8Orfe9qSZZVa4amTcOksq6GkfZNnaJxZ9aVWiL3Pk6nSNmDgWWkv
HYS/EGk4UmRXDhUePYXBEhQSObvtsowxrC3pjDELo/gEWj156/Va0btmJBXf
hphLp6OnAKuIxSgQIT+mg4MxvOR/C23pbfgxvHp/DvPbq08hDWYOYIRtKwKE
lwXxSaVGIYeEC0ftr4aV66G/22SQ2chla4qGVvKkfNeqU7KVDClDVzLvWJPY
g2dZ57hGCdL5gtS4XiJs4dcUOSn+M1H73Shv3fZyCNEdo178SXHpFy9Gmoaq
C7+6rM6SJgljM4C9lE0GdqJUVvkQFfuyxywS7z8nqzRqlZniBvYn7EqgHnLo
cbOsw+qoLOF/x5aLjzAk0SCfvJhC5pE03spYbPsaHT3qcdbK3Q/yDAAZZTzm
DV0j/PaAUI5qu/cfi58W5zOK8Rip4PBhwYemCEQzNgm/1SVG5cBRNVMyx2Sk
iVUqCXh2eZ7SlDhFA+HW0m66KKPoFVm60qxln7ukyCnE2gtJBjxfctVLLVy1
SCHgMxg4sSGo5QolEe6apfOvKUpH/NLogU/f8RqsPv6G7udIqewdjqEOcajQ
QfZG1kiNOPPfCPUz/cxY+sW+pZdKzSt7q88ucU+aNEZCTm14VAfrPXnPToM1
jeFlqjjxd3DhtYA/jgcsalGrm5bt3OvYXHlOGrug8a6RZ3saX0MbzlGlmwMU
RGhyFk1CtwGCZr42xypgJRpwWH7i0/ZZfNih0w7sD8maf0vW9iEBHRStEmj7
VYwUlDohxvwOzqcjKH4CXQ3l/ll3/pqcU2mMVoUSzcrAZaB3sUh4Ma5DTlC+
FmEPI4nf8v1Sh3LTvQdzUkajY5raOB8ylquViCmVBLgPLKkzlq5o6JDVe9wc
QGcuxF5tHarD+FZ3rvUt74YXmFHdzBVAI8e76MZ6HPD1/L6DJMMiAmRjEOU1
7Inbh4IPmvgzA+mxC9RAS5e+zdD2GKH8vG4MeNO6/LjXEgYaFoDLIVnoJanN
qMHU1V0PerKZd7jUWa/5LWc8y/btEc3tr0tPEC3TT6x8cvTwQB9EcaaYhUwN
z5sdQA3mynw5fvoBXfEilvVN727O2XmjYWODVj0xosmT9rlfXWDYcMPxVXjt
EiZ9inqRV6H6OAmXP9lcLaLbvKtB6FlOIXGUwUEhMKR2A16BqBXn5x9pR8km
Iz64Ivi8qEkT8UboQwlZRZl2PN9RiOEFNtM/ecy3MiOM4qtb1Lb1Lahf6Rk7
q0ovsD33sfMWE4VraiUBA9gA/ugqIcowEPVNocilOuVQ0nCZW0X2DYDWzdKU
BMBzPIVGIkHgaOJxIDKheF3BpcJlnWAdCMK1kzfVibmP8JTlqYdezB7G1N5g
QRWj0CHSqe9dDaYCdJdjxmnWBlSo40vY5ISkEP/mxv5egybJH5z13zncZdRm
KJgWSggMejmttS3Z+lTSZnNqH1/9ojonTfBEs9PeGJK92g/v2PPb+ZEl3Rnq
BpUIVdGe3bGqnO783uWeLkOP+CpPbS44MjG3xuyzDSa8XTiREweHIu81Up3h
B0xLCeNF0AyNS6OygtGSwnneIgBf5lbulRgFW1DgZSPDamNthy8E/NWejoYJ
brTH5KJqlptmoX6Z6/CPG5URVffaj9I1GYLb2V4Zjb6BU3YVm8GJo0ZdSRCF
kPB3KGiInW2ADjjosSG7hSxSMk5NtCnYENBIpPe1+agkpMjwUPG0grB5QZtY
SIVUtX3Lkug79VFv8avRCrWZ4L+AK2jMEv/6YQdzG1lE1m1hTO38STYgdFeR
efPmFTlhSm35eIllP+LBhuBumFk8kKG0CDzqDkD43X3bzQ/BfJhBWbf58BUU
qG0vjc1y8II+8AzBJ4h+uQWFw0jIWPEUvlez26JHaAQKMGS0whflVH9fJ3hT
PnU8MtuIcRcqm9p8isUnWjjvAwZqIZGgD+bMWIdKems+puCCFuQpoAwU7Nn5
zXBU5bNlH4DCutzNQWq9/NGRy3D+2zLpqkIKBVDArS79L7pUULS3iv1fA/Cp
mlfwwzZteBHT3U6V8Yc7qRBaaRXF6ACtsPmoTKDsIkUrS8dPKBnE+YDiT5HD
M+yo5fZWnI0F579qX1Bs55Vc7dSHorXniL3QH9rEds0A4esgApFKwGOnzN83
ZINLjiaNGGrtROxUzXz1UnJEFN3qkWfa1+Yko1gFwmwgU5DOEDBqf7HhI8OV
yt1N3vGSmBUaWohQEHcK/aLQguRSSXf/2UDg0+7orZfbkx5mtwXSdJxgAJG9
dq/PSIhH+POo3EEAYR2a/1hK7GOS9LF43GfeN5ycaJnhwKxrTaNfgKDnryJn
ERWSmGQdAjlHYOB8Qp97H5YS2ADxig9vj6RpUKE3pjQsI4udH4/QNAz2oni7
Xxcjh3diQUS7j07E/yEHN1I+YBa7cVzKGOTYJGohgMbnBqJWzv5iySkSijqU
LvNkSxZS9ac/6sbml3dR/8LCX46auoZCoRU3iiF85XiO+XTcPtoj9/HJNkyH
a2B52a39bzW7avli56e8Av6agc+cCy2g9Egz5vabe/PjMPtb4pVCVEh6UEnr
tYKOBZS8B3GHNPUZ1oeCyZYCFnoVtTJD2DYyWRPRajBkLFBZAFn71quDQS/r
PkEwDfD9248Wv+iWSLiFZb6dc16whQ47JpRJVu8ITFCW5bx1KbT1/CVxHX7I
9YDtIsCeEnEKCLIao7SpYQoOjexrOipE1FYpFO7HpTFXEVygcNiGbUErdl75
JPtGd14Dg6WZoWvNXMLsdKPsb/O3HHsCSX2hTKyui1jEV/rj3d/Az6RFjKKZ
gcCKD4Cx9z+Yog0Ragh7eDE2KPeqvJVojHoIRj6AJRnRmS/M+NJLyO59BVaC
88hNI8YrLcr6IIZoBOIQ9CdJ3xPlXzXoVIHVnHYv+X9yBgrqTbNtIDX8SZ94
SrJi7oecu099O8BXrx2Wb4mcP6i4XStXBT3leCZUJOBWu6/l6PNnJNmTHy8J
GXNqhh/UXmNAr/faJKIS0UEhcSYnxJfm+9DW6/hCEQu4VJeA5Tt5rWrv3NIP
xTOTkIVCy9udykFh3y53wxmDsKJyWZKIwjrXqy/YkSh1yHmWBfyxP5TaVjEu
f1iMqx5+542EjAXDmLZRAi8TYXibyiJwxXtVSTR5SUBn+vn1YFDGeTKArR1Z
LIN0sZZdWUYQ8lqwteXCgvNp/FGu0F1svswdIoX36WCsdlQz5aBWqn9TqM8F
+X/5X4DODvcjnbNF2Kqrl3xrtb+9U3sRiMK0rUR6EeY2wNGFL6Ry6ELtvYpG
52q5Z8GJTcJx5kHezRHeJ8mghbcAoHpTHlsV3CNvDHXHG7C7fUt2RoTd/yTJ
uB869wX7Mn+17fiPyBIy4/OLdMCbMwGKF41fPIRuEUSRzLg1oNNlPEgazzbc
PYgZW2JDWDwpBsu/jVrjDSx31gWYTTJ7FXRtZ0mPeZTK/ZC/5TFR2nonjyH/
FUm5r88jf0F5jjq+pTQHIC3otcuC2xWGrX5FhI6YREf6NgZlRQg/UutXigNC
QZUQ3CYq0TLlnNQLcWYHWrd+l6jSyYxmSfgW06X+Q8RFUHYcuWO9S75K+mbf
TQicyioYT8LmyUiluQE7NoFM7stnoOydcyMcJ7QrTykLI2EoZ+zHpCsb0B4j
bN/T1NEdvG+tIB5OQsCF4HzIpWkbcPoZ268DOs2g0Hp5KJ33idSIAf9nCxdS
l15sB2iOZSJ0ft5Fi7ew4M1z8dpzpn7BHN+BjPtdD+dQpPGB9qvNbc/UZ8bV
stIGmLKnSUVWYg1hIehZD3gmE6Ty1qa41nF1aSPrnegfgHrwA+A6A+AN0S4X
JSomY7sgASdHangdrY5INgMeIDbQB9gCxr0duW2nh7i5d42V2P+15S7LGKGb
uRF06O8aeykgWfnrUl9VKqTwlrVLrWQ/+piaCLXk89nvYhbXhhvROna3YGLf
dVbRMdmOy8ojyGlxR4hCKm06UNrU/PX04W39JTWWfZfTy1MkiJKv4T5IkMzy
pAPC5GEFGqgUf4CDd8zhGAleK3fSt2nyoRSHT6AEzrBFziJ7S4piZCtbdh51
X4rrskJohTE1ip7fkmW4+Z+TQcpoQ8QjNDNWbU0QXSMDSH1OUJJB/UmKqlHh
J90n0YiRNorppZFQhe4wDmvLg0eyHUVf41ncgAGJtWGYg81H9FwFY4tU8n7l
IA+na/mSJfqdE9ZkqXnSAKqFR8g0+vvO8JKfpVjWroHXBEVgfPWVmWDU+Qc9
eO96hKe8NtaJZr30ZcOgHnojx+QeHWL2eSOWcQPdnSuwGDd4veWit9ZNMhx2
Uy8vgE7ZxE0gfwkDoxYiltXREVUgWoBTFJf9+FDVJPMebbS0XyvdYOiDuyh/
MGhXPdbdWhkoB049jTFMeO4VfzMt2ASgCHKlhNGNaIClmBs0lLf/KCIvFMAp
kJv0VGRtNzYkEICGzjymxXcCMShUO9oZeqffD5YfWgbXL/2SlstY7ONMwOh7
p86nJpSISQa57CnElfwRmvEjydcHTzr3kqtJBo8HpNH6VUykxberXOMdz4hW
uXadaL/4PrLxcd+hZNRSPytRnlXm/0jYTOIC5FB+Sjy8WbJMHjQtf9AW780H
jKRDi+xli3vT8ZmL9D1teeZxe94LcaMstsD+hA4dKKHY9Dw70rsIYNa8H+mb
nP3LCFMPz9MfB2BVnZ7lvmZLEtVDuzZrfIjJxO+DcnJVrwaQt3uHqvkFSn9g
mk1xuBPMuI1Gb48yVswntjwDYF/Z9abnmueBGwyhXIl0OFHWLzeoJa9xAv1r
umNkYXrBC0zv5lD6Hm1KBbRuO0WGAdC69lSOy1q7k9yjIHKeeTplZIk1FXwJ
71CgA/0cFSLV75iExDAQc1MDSwtH0Gs24G51WcUBWMPX2WSFHACVwGMuAgfz
84LsvMoOwLGRTJu9XvjhrbHdSYoEmpemFgWZgM+5XtyJRseg/MIG9VDBycWQ
G23vTZZ5fesBMp0cJ8l977+KqjTN/VtXScFTDcOqV8rNqt3EHVt8nMtLqNCr
jGIJqkdLVYmuI7SC/Zgk1ohjSXCxXBaJoadOdpAXAmEwWUE8Zl9NHni/M2F/
71YbCoX4lkz5rp/Wnt1t4bE53kawQkZ1U6DKQJs1l1o6vD99+gqyLeNMwq2b
dHXdAa3vUjriS0+1jQfqFiZdAbDjMRkX2+dY9JcIvjXP/WihzHIQfQocrG4j
4nBDUmPMlbOiX+bFoGzzxdu1rLCDtV5P7QbZywqpsK1rR4yBeuCroOIVBw++
s4sRwUnJnSVR9MmnUbqKNSjWqBxFm0+J/CkhfgYtz6SIVf/lIOpb1U8Kx8U8
Tp7E+yvNkjdPAfImvG1SV4O7x56fGMNau4oKtPzh1t1Ws4rHgN2jSTkyw2sU
wZ0PKb/joaLAhOc5zQgVXRIP60CYU07r3EFFMSgQv9bBS0s2koXEjoVLVlQ8
Aajpjfag0s1R0YPOz9M4pYKOdbIjJ25MNIJEP2OEcON4BAuNDVBwxeWJ8P+Y
GbakRcokMb71u3oJtw/KlpqqivC0+R3gn3aHzBbbXfXUOnZSvstob3qasUN0
yyl7+RX93I3+rcwngrBzkQgPXQBZtfWdT8srKjfyJf4qoRdifcwITx8sV+OL
LqFt86wjfsb+4xha/OVdzsSbhVDtwFKmJANmECotma/TMzG9Vzl0caNhlRh2
0XPh6mLmdzyIB0H7CoRI0dK66M+prg4u3SmyosTopWu+6XUWOIZv+iAX8am6
it9Cv7e/zoaKppa4EAqZ70lSzwoEbVqbLtXMIANuI5zFwRDui03ene5yChTj
fpZvDJQ8DDBx4YB9hLUfiai7E5lgbxRtB/u9hS4SelKcKAerlIjOsUp+zcp7
ujEikt2YKKxN+/OS5Mkxka4sTQyiIGk5gbqUQ+exmnmnzwyh3Fn4UucU4ucv
2bLz1sLsr/DuV+PRQvI6N6zBANCJshW5YwMq35VNwb//X9tjKKKaH/3UH9KD
VW17m0qyuFQgxWpsjXrqJPlJhQbOnZyimocGp9XisZM/vXJ+uL6vsLj1b9zl
JupSs51yZlmBmQwdXQrLC9bhcIyjgFWOOw711bVhgIqWtIiCj9dtqk2sCILz
tgXFgeh7lvHu/Z41VDjY3PsD+wfUdhkHwnHyK8L5/019C14EKdKY9FioQR0e
XqKVP5W4YD2BdbK/r1Xi+ciXH1r1TN7jZq0Xt2IGtr1arT+P5uxLatcMh5NB
ZzpIk/7IZkhmsgwy2aQm6TYiNMrxa4j93a7MhgZiLecGdXGxvWXWN0WEzSXy
J7HgEse81M+5KnOa0WYyZygXBJUDtFSe+ItufP0LhAW+oFIx2VMueaTLQRox
KrCQfTy3CLBXFY7/XR/fTWaw/gCoQeWYg/F027cLqTsFuq+kz7klnKZViuv8
URmIUBPHso16ZlYjbWipoTeaUMpMgTtP7huc58sgww9eMYmo3iUPTF428CC8
3sV9oOeTHMt96jrcO02+MXUOkPcH4LZXOgH1ShInC7XUzr2OE/Shcam1Gbib
DhGzE8/mOxrMMEASBpaeMlujUUTlErB6T4Aybb3ruq2ub0YpCwYURyTN6vHz
8vB/z742y/2tbDAox+pSlH3ghlwgZCss64DLl1h3coxqY3OX2+BNctCPkzmO
sUpHP0RWF5ewfxoJ8IKBrofI6F9e8AgHGllmZlsj4VH9bPezoIU+7xq6+E+I
StYB6aKtsl8APYXjWRQKkT5TzbrxQtANiqH2hPBFG35gd0IUv7ejYpTdl1Ly
0WMc63n4qKH0WQwE62+fXNnaV9cH1t1XXaliGt56HWn+XDBBMSzY0oO26DCT
eVC4xovmpMiJFj9l2NkYq2c1ocaCNylB1uonTGRA4MGhblVHg22HaguUcdFn
BypVgVuCjhnWJyVX51CJN5pnHhV9kcQjjLnpKk94PCSxwE8h0bEDI9ejUZoS
od11NfDJXr0rKj5zCGsHRWqBlzGVB+onZUwmp7CiLFwjAfqFMXQJY7BAF5hA
X4GzfO9XIOyDfMJmVa0HqyordXcCjRllspCSH6lvH2R0baWpZbFTYG71qzxo
W2JWVYCsNW6xG/V3tMDJEYFRVSkBHCreXNiPuUIj9s7bgUq0PtYFJYNxPceC
N1c8FrYVDLHTXjAkxqaejqtEvDBTwDvkrO2Da9U3UueHoruseJT4pvmZYN7A
7fqBFdbKlzeCB2/6xXwfyMMtuYNpWzgYPG8SKnXsrf6DSmYVGK8M2RtXiFfi
SFzVAvH0LYfuLucwb+1aGu0Bf2euyunMDwCPkA66LtuoXaOedRkJNWyajAro
88ycOuO14b0er1z1+N77iFsTQDX16dVMOW+o2EFtzJ7tcW194Z5/zrTI1ULX
bhgtuncipubjfugoR48d/HtayI/b1lZQk7KPKxhqFUHiyeVVhNw1UbAnVcEt
EzcqsffgDLfsKzS9KVoZ6gBuLEFvwEr45dYdIO1uXraZygHw6o778QAL/oBm
2sw+iol1XZmbh2zqE8G3171451DYrm42STEvj231LvPgNJptOYEBa6KeeOl+
Uy+aMDoi6sWIZLDqN2AzfIaPk3nxHW27A3ZXX11oryp7ZAPrBR7rPNmHTANy
WtqYBytsJb7+vd3tlLDis5A3MAcou3/TZfOjKk+0Snlos/OzFPlyTQz76oHA
wydWp+NyajsTa1WW3md0sIf0Bd9IWIPOSQ/kDRfhuS6ZnnfAltFo15QTmr+y
gGjuQIEps6dwzy3VxggOURT8WRI2mysqUbExJz6ieD+vOg+D3T2BiR/nSqhh
6F/eQsWpJI2ke3KskecT1FXaPCQWa3CchjcGWuHu0MnFX3rsdRlZF+foQnm4
6kRhT4Pzto+uPcH4UelfpGakZ/+383cliZ7eLkJyHVXQUK3dYHosG/TNgeId
EdDmIb+rIlDUNPh03hBfvC42SP73dd+AXHM2h/6rGFNlEU387ytbQBD03Hnl
XEghT5bv4PE2fZvHevTBwzkvJB4bKZHn+NmjV5Ns4HRegi/X0AnyB+uixBqA
a/2rnre33IAIiCbczmmbflqc5BHkLlIgdtgJIPauzU2hsNM7rgUo0wKM6l2z
QXTapw2eZykHDbV5BfkanBfpAqw/JOvjBRqC7MjGZaNZTRQkeEUog/hQxmk7
Gz0YoQ0AxWE9R6gmET1Ut+VoXs/f3sm3gOhstWGENNKrjNitnnjAFaZ9ALT/
/zGzV2Cka4g096hz/ENnk5v5ZT0sYYO4a28Uv2NxQ1SHsZG4krv2Cn/XdhqV
1k9ndxPWgdEr6QpvXBHdAezORKQOq7f5qSJFjdRNj14PBCMjvuYXgcy0C0pR
aNIpcT+K65kag7OJJGgfQRTIcgNbzQB9dBmzT8jRr5HjO9m7rBm7ijx79bZw
g07HhfoyiGd7nhNzhdBgI0BVj6BQHE/s1eCE4Hzk9enMgIZVtN+JBp7f5zb0
2ZBaN6UNSPIqUevP17iAYIDVrTWiPouXzRjfEj3PSrqAgNF5U6Mlpd4s685c
A8CTCrM9etVKjx7dDbwMjDg2syAylmGEnbrrLgKWdiXEe6rZifqi+NJDkiuz
cIl4QCmeW/2XctslpQS5ktQ570pB6criZoLA7hR5kcGlNLe6ZH/7gs3rTx62
Wb6Vx3bIKBbZMonTplMoFH8zI4BB/GZR2kZi5Xh4+YHhqfxu2zN/QZ5CP7tN
xoFWemZhdc1ukA9CyPbecW3NPqG+YRw03u+pgMoQGF4H/PFiLjERWdlig3sa
fjkPRTwiNefBxuFDwrymy7lC5WG7HncaOJiOaEvZE7IF9cbUMRRGN4Ft6EdI
woERH9zmQRu703OXeiptQjxbvFluZHCaDy+N8tOtZnvk+CvvufmZdy6R8PFG
7F4FGEt3NgBvKqg+9N7JF4+W6UI52PQD2+/bbjOsm4ybff9PcqEVx1+0/rOI
XqpROx+j9CesSvkw4zM8HroaUWu/X42PTRH/xcKw38XscMATOVO8KBHwm6q2
vJrQ6eJT+LRHtQuiLbQ+vNN+2eyiPXGHcJ39Bt34kCuzNc4uj2OuvyEJI4q5
km9i0bEem2VPUDVJfd/G4MBQvC9H0UJB8u4vbw/W9UeP0YpqTnPmlct7wNGq
HnMhp0y9rAX8iwChlkpcLuuYs1AwzYB6NGQgw+kigLjGE6kXV6UM07ULQDqe
e2mBU4c7gLwLZEPYF+YN3HMt4ATfdXlF3uArQsLcfu2xlaORQlIGjyRbc4QI
4kQQMumK10QnZUmTYeZX9yPYmkSxIVfK10VqUUVCVFT4fWdnmqdnCzLGLtsY
Cba9E8CvPopm7QlXdZthFXR6EMA21hMf7D6f86SSleirO1i8Jqn6WS2MM0kT
Whbgcb2d/NciuQtNXPJnJaGPs0bLutrnehsq379m1ZBnBBTrTGLNJlcV2ZnC
SuFqRfv9aQiUT2Fva2CDP9f6roqqEu0hsyBenDJXuuInkbUEOKih5rooyYMZ
/0VijUhAZhEo3w6QXxCFnoDU/HO2tB9POrmCWi/F3n90dx5jgKQB6ZHhkHyX
d3DItgUWWacVIPO2oDv0o0xga3V0bvpzhylnlqr5LnQguKKknAN+MHhHjj4U
xQyN9O1m3XQ3ANd0C5t9WLpGc2l8p1TxvybdIwHjgDNCN3dURZTV+tXGBHPx
1Dv0McoUaj2gXKm/LZzig6TqIpAauLwPP7pWgxhBZjUqAsZa20ThMX+ieBw8
Rs6udHiMQm7+8izyJWrgmQjDRgZwPs+L30LekuvWmiZNVLgLuRsRV9E8OS7k
Znly76tbGA62qqjllMdXe4q2s6x+XM2p99CiFwuVAapvP87XzMNz2E/yMJTm
0EqZFrEM48rC5ByQlJ72wwyatm1ApLS58Vk9toyXy5jwUoNdgtM2b8MZNPUV
5k2FoTqeZbSnT0fVgTRsCHbvzMikaLCLSMfxeHZQQTHwEV4YrXbLbVdzZDkr
352U/iNRqqwF3HjFyPxf/b91IP4oRSxmo/hxAMZgKMeUpLU6mOgbCwq/vb/D
eJH4QWKtSXcW1L30AriNz/wsrnGjOCbz2DAF0F51yxw0vd0vGX0iXQNt+KDL
JVO+Bob54BmsMsfwX5hADYqhKclUA7DmtYHmB/PKHh8h1AQat9oUxCqhspPr
BSLb9MKb/6QKrMRsYBxr7W3lld3030tXojXU2oqWvLiLFSLic4g88AlRPS6B
U4TK0JT7xGunK2MpqKcNRE9bx8+axxNW9ApycgE6CXUSZssr1UhqxXb6qdiK
5dDLTh/qUQCnrsG2swatqyJSsZ6ocFxobC3UXjm/2x51M560OLM+kim34lSt
ivwKGyyz8vrebiSufLH0OLz0QpA+1opInG/avxcQh1FBPCHfLnFRgcKxh+1+
kBJiu8pOfi/CNmAlfImAImxD7lnEtmfP8Ze7EoelDYc0UXVIQpD8akw1YEk9
tquutfXHFpT4GWNo/XXNirxiSV2+58hHi3CiA+MKJrir0ZJf2F4mH8jOx4Oc
NrMapAFeQYq7LAwbQXTDK+WQ3Fc0Hc1G9nNVIO2vQX3Q2KlEpX8x24hY68VI
nRZVKbAU6iKO7/vOqUbg1hl4PQ+w/gt5ti88SGjvbPO5uTJ0GV0Gm3OGRM77
X7EYixEfSQGAzegwGQBfgi3NqDO8bxrFohqtHrRtvanRXYD1BePDEh7nADEw
7qXYPRg1ovH18MEs/18bzjkxb6dCN1hxBMXo5VCuoGr3dzp6WRk/G/ihzwGA
XlpqjNIjuxTD/ywa0koX3Ilx439XsdnBoMiHMeC7VM/PTIbJPOB2lWwF1i4Z
O+TCNThnqQnMdHmaX+5AhLkbUhtDkODnbXc767ODGvq5YlD2dDTHnNTnDt5W
paZUMc0EOhHMYB+30vDFzg4YlBvCVVtRmmqogITGvZsQVvJEsH7H6EiIit6f
0pB2U2xn5k3lB/o9Cl8CpRhjmKTqUE9RCJuwku3N5cGuUuL29dsWgxRnB1i4
P/lMIXSZ+Et+WSbrb/oYMtzitmDJGDUhbWsT6KO/trzTu682IsUCUpUZvQOE
lWdFaVJmCEJWhOXfDz3akMSFJyckdtxqhzmO8EtrGIwGyqyz/A1kOv/muG1C
f2Ptdv61nnYQdUtvFo6lg0XvWvoVJnfWul947ArDLwTSkSTVCSrq3kJHt+zv
VmgnYIEKGj8MBGWetvhWwzwxnYW/n4f6K3i1N1fvrY5e6/4oNCzcuKJZ45lN
Va25uWov6mhxCNxvW8dK0gkLsQDeQ7EYKp+/9tjkx+ZEZTpCONwvbEMrPpSz
kEVesKHltI+u37hoW8dSciyy8+FJ9vFdNs91lpt9GXvOaEnHWHRN/eoH+GzP
8CnSW8YXjpUxOix5YaLoGfHESG/CI8czsp8KyHzPP7uhIXf3BRpe+nBx3Hz0
GbIz0viXJ5iH+TCFTnCijnwYGDRJ9o4YN4d1fJDb07o+hQwANfWgoIDYe7NR
4kN/DHagS8AzjvTprANIe6SWtjcOADl7xzZaSUc5/rTDNVLPBXGzNihfJvOF
HEE3Z72n++sCwVDO5gSM3US1ClCYVwD5N/G+A5Nor+8ySe0HFA2Pg3k2uJ2r
JpPp+hch1Gu2OB+mzvO7P+s2N/SPzsrq2EErLeig3xDTmunfWP+HbtlFZIfF
1/0jC0vIWhLsvJ7nwtffM+MYnHdZdty6ylwErkVarF3NLpdUpdSAastDcyZ0
REpZKN2B+nxMPJO1XVEkh8tDzUGgpHnTlKGdF5m7eeThE3KZPFMCECDXUd2L
3abkTzN4767Ug0QQa842qcaDq5D2wwR+dUQxt4D8SKb3uMTEzhPz1nDecx70
CbadTXa6tMjGJ+BudK+j4Xt5Dxw2zOHPh2FbQOzwoaD9Ieytzx8romSpf/4x
wd5pspH3PRF65xzI8e3o1BKHGot6sidSCcBJm7vhULaYTyCFd+wR8i3VzHhb
VvTVsjLBRsLX37jtCJ1QhXhcaHS0eHM9MxQG/lGzuAXWKcYchp6FkbDSNNt8
iEH5dGurlr1zwSA6solaaGw5ms3WATXAmZ29Su+s1/D5yJvQsQZUex9RmtKN
e+ByhSfy9IwHyCeP3F+OnCvVKei1Obrwf3x4/JGW+FKRamBt4ghS5gml8Kd3
JHxzJGkDWut2Ncklh2Nr2QG3EE5U+sjyVJVPYhrtijXnod0iwMz8h9tDCz3A
GTRTl6f+Lk0FvMDGIvrtzKNN5uBqL0yNE7M2oP3NtfilPlkoBJz1TR+euGM8
2cn3R4VDzmZ+YCdIYnVzDylYxJOOVu8j8MYP3Gqt1WYFfVkp1JOH8pIdLAgc
X1xgWJlIvN1WNrg6xswFpA8SFIWpddZpXrXLrHDYZap+bD3LK+4/tDA0lcmB
aIB8fMYFsy3Bf337rBp1FpgO9c+I5BdTrCgMu81pWsR9lTBA3dYr/GuB0c6O
j2O/7JFivSE7hheqkVAV6F2AhsLAA/dTLtpN70EzrWkwj8LJ+eDPi9FTvE94
+WXjfl/yC2xMGcoLSKF/ITnMaQeGdDys5UZ7CG1iLD/KO93zsvENpv/wEc7I
qgESmgjBP4ihvnPcEscqUP+auyMIDMSTPi70a6MCJFxrcOejruMti8KbYrLF
PZwy5VbmMWbv46Ra9W3CHmEB2vXwvP/cWGkvo0qniLh2QiEyDuWX8qtGsvur
WxAdzAvUa1Q0okImY3R8WIjqeTPT4e+K25sbLkKvah6KVwn91i1k2BYp8BHM
j2DU1HUqEd9ztdfbJVC17g7z2Ght2bSmXp4acyZM4hZpwtWngUqJzl7yuFcp
hHHJ31g5pni4iY7MK2BuprgYymJPR79oD1EJXIxUvKZTF57lBp2VrCsJOSyU
s5tFItyFhE7OD5ZM/IbIQJssq1U59ktJC06E558snc/gSbVAD+5laObfIL0c
JNPr+yHUMaG00be3Xd8FXgalt9KhCms+aftiUx+PpUo+B0xkoTKPQy/PW3Lw
nV+HlR9FGSQXvvpQr3n4Uq8E4R7rXcI8o7/5JwyASpdT6/qsGHVHMXvaBjsl
jpHvBNTvqAOGbPDavuv2sssz5rYqhzdWvDxC8Ov/TuM6WdtlANuq79WAHQcE
jwX4lK2aOs5nBG4Kx/ovBODNiCXbIH6NvDotv6J0wJyV9bIbUkPHCjFs4QWe
yeJ2Qhlojbs94MLIr++p15tse1tMZS9RpBJ2d/pEplgvZob4Gdg2tYl1/ITg
BKgEtAp8MN0IFh18qfamFovt2MkB4SgbcOfl96mXRNczl+P2FfLGrR2fgbEd
K01+dWLXm0VMqgxDcvuRWoPFbPTz0S9+kliNdIygSzEd+vjfsDNQ2ZkBudy9
LRLkfY/JmS+F/vEOFLlomC7W3rbyj/k2MChfB0Y6kRLw1BwWtXtCKlKVA7s6
BSkDouvKeQ6fcpQ+SiL6T0qzcJXc5eDbxBWGoXKVogQJbzYrl5T8cTalqDRU
xnyrRGYzwWOlWgyNy9f19vm1CoXDTO96/KSMXxwCcLA8V1p59VD0IRxXdUlS
3ekiZNUDOFbZVkAAOg/C0MITfcDcNAJMCR2Z3dve+j8f3Oaq4EITdyCYpARI
W0Nc/0kkE3BfqRHTxqXUOdqWZUjZ8SzfVTSCRvhw08yBor4/L3UNuh60oxy4
lPJ5lhdKp8hcPD1ent9U4cxKl+5FT7idvmdXJdDY1NZryM7m/ahB5Vg2Kv/P
VZyOnKS5vJn93uX/Zg5aT1zu8XdNJ5MxsOh/37/BYQEI/u0o1wof/L7eU4L2
vyitMIp4ZRp1ifg/SRYgn82vo2WEpcTGshHIE+oianYbuvJur2r2whsQCmjj
rDs81niDGSegt0ot9sl1zSOTQ33ejOw2OMgcnJJwKHZbESPPd4gbBg7HW2s5
9u8fqf7TXrp6B+owBim46py/qMuRy/d8hpCKzn/+EvuGY3uq7XLZ85Iy0UQd
YXk2+0D1BgOJ6je2bEeLB1muoyPNTmJMW/8cwPEoQdn95jqkuSBFTeeio96C
KA+UnGrITYPCPb8fsnyjkgdGeOVUs6f9Xn33xdnxCSPzY0DSY/xdFdIGC4em
SfWnd0DsrEhez8flSgcIsDF7npld6cUIaPyJcP1zKQGWQ4qhJ9yqJzjpaixS
NKy7JLVOZwbYH4744TqTk2T1uTl4m32MqjKxOxMWxaIFofr6vuZ9CjWrZXMM
h5XrGedMK3Ljmq1SmSxx9pwxXebwy1YziqpvHfS1Opj8o6TjoYygQ80CgR9A
AcJ8K1QTwh4jmkYvAHqU4t6nits0qpplNoeTBM3qDiN5V72eMvR70EwxyTc3
REBjPt3hCgKPmvAFa0HjuTr4N6pUpu9pRSir56M4ZPmiLMxRkhVBR3hCaekG
smiVbn20jigFN2U+2rImBxNIvMoSnaS/gWryUT8gOcw2YqlZhRTrG6alZh2O
n/CQ5kL56xGGDZDsHMm4yqczDZg0u4g1uZ7ICWYut6M9NeqeT64o3nNV6GsB
eLusB0QXPwEGksN0ecFv6llmJ5daIHHBJzFV6YLkjL9ykIGiS71GCcvw422z
3exRnjkhI7WxBuaoBe9YERSkJjYeeDyLzmyO9Ce+9pmul0zbIWZhDQrjjBL2
uSaw8lSXNOGJP7AwLypck28kNXMzzz4jnQqRl3+jWY28IPi+PRpHCoif2RTY
nw9dYJqFEgb6H3RLzdfepeRUDQt6C2038OwPCQEAeE9ZHDq59Q9OqRfjhIYJ
BEiYBwIfo1PcjXYmDtmBEENifFlQdxiqjf8nHus8TQNuR4ZRhVu8lsie+1nb
JvH8eYgmCJn6H0h342KwzcbmQQ5c3YyxSWV9KWw0Q0S6Xi7oENyl/V/F8QdN
bZcDTiTMLx/hNEpROOe+tkJy4gPRNXQGH05sEdNkVt1QatmsWQLwxmd/LlFT
xunGeD50wF7tAetv52nwQLD/U8QURuJ6K8H2AYpl6NR4jqW+NnZrErAh1M8x
HnVm5To3XugCBcZi2x5TeBc0Yx0hRFdTmUVUyBI1Nsny6U0uKWlzYIDs+reo
YHuYIh8wWaptJvyxyioSVD9nz2XvIcKFRyZXNFsYSQKJglVAbLBE5KKhm3SV
NM4Pk+njaUDUThfn+oHsETuOmhxdtCJ4+0wUU09sHLajORRXhRhH4zADtQSI
94rDLQFwODPrKAlY0RjhtgzNJYK1hqBwql8ELbYUrOntYvvd7GdJNA9u2pWN
hCaGTztm8duis2l+edrlMmJCm9Zy4eQLaFE+BwW52gW8ReBTnrJsBDZqL76A
jMdYtmaA642eXlZdT9J8xLAbh1S6DzmhOhTJyCFEW9B695IraIQRnp914rgk
aDg6aGkcKJJXHG0q1ds6hN+zvnd5PcxGfSmnEKKb15Fz5jpOEc8ztCcrSGOQ
kjXVkdK6/ZkzgtLdTCFxzQXt5gni8j+vwMEkiBqnuRIXYTkqKqt787p71oYK
Yyp835DaD2ZVjzdjDgv6/8aor1cDo7FA4HA2nchF/EuWUaneZ+pdGmBd1rnV
I5QaE4ugQw89d2N8bBF4QHrvl3XqiCH2+Y0D85hquyOEpREGBeFKdG/qATBb
MSxYRpWthZlcsMZpPja9DFMENMS+vuJaUle1byekkKC3+UMpOzUWC39NYwT6
Rapw1UnY4ivp2xWr8GeBhi4R7/5PEtxmZaxDkSi7xJD4IYwoVkzz01N6899X
fMqRUEH9hbqyeK8Rf0BDU/xDkOiMTIjQ1MbHKC15YW8VBlHsRTAJw8AamP0Y
MOUMQQ2hBiYlh67lBdFA6e+/8QFJy3Cd5rRmxgPR4+yX/A6DZm4scZaPgzNl
fQ77GOcJr9sx38dhTuz7CJgGVVhBqpen2dvs4cVPhuS3TM+DPlEwR16lxY7z
2mPqhkQmYN786jns01hRrp/7Mjlz9qGSI9h7J0k5PYct+2UGTYjPJaPuaAqN
KFzGc5fzxuINJUcZjmyYhyhraQit+mWNEaRN98gGL0w2Yd8JKvlJWStvwJo0
q+X//N7M8bpWyN0MphHGm15jGv39cJfXhlnXbjJqATFakSlBRLko48ePgkaG
KHoptgDT59G6irkCBjpC2fNz0blUKiF233xReZbpWJHukHZSo98oDQDWcd+G
jS11DgEtyoYwK1GELejPAzokuSZA8mx64WlzP6qdn8GIt7jx/akVhMwiu+ks
5cwgx9xpgRtPK1q9pyGtg3/HxAW7s85jlxEBHhJSChLRcbUuj6FXG083tOjl
Kb8DEdxdeAkYVSNbNDyCpJMULSeXb/JIBK0Wmp2zp2ykFyAy75xIzs04RkFS
qs5oAV06Q6y320jnyoywygqirk6LWyQmXg5oUldEIu6bQp3gPHPyzXEjHncK
rtW30HP1z/5pCED3S5/F+ZU0Xpklwve2qC8yFDnrcNoxbjtiMHB6oVtUzDYY
/9hlH2E9y2JK+ngtzPxYpPmIWIr+D7/NzV7o1hEB4dgc9l4zdKV3HyGUvdxs
K1xWCBKR8GciBYM0Dt+fdsczwFfubn6Zmj3UD2daUB127EHTQXcUYkfdvti1
Ku/EE7RF7JwHewitlfKAIqxG+wHK8b48CeJbMMAv/0hYSWMLa4muXBO/MTHU
b64iASRIzWUjM3N22KiWsYSzhHd+lBDO6w7azQXIhHDIiLOiDEvO0ezJFug+
Bei6YKQC9kkzCX+o59SqP/QttRaUMRAFKyg+L8KVZglKJ8ku+2S3RzT+e+/4
WHtNDyEAl1hw7rlyWB8SIJSAy2IgYjlQDcDEWlUT14pTEtv0GuODgwEHFo6W
TYHRP7VYmrm7dlXZCC1tmcdahfMMzpKVcpUPBbM5ru0hfWKTZJMFVscGB9KC
ycezHhvLhOHGrTAQRmNeyk/BLqZETbUHy71rutAtLJWov3Nz4RqtW/8j4pWx
K8BNGouFnDa9B4AF0K1VHXQ/fpUNxF5uruym8q+cA0+793oFlTflMrFXYboI
dx5mf+SA/hffRbEwilmsC7FgFv80HAO6EIaFnZdVgvcZP+H58J0KfPuTe7wo
tniMwuHgI3mnhcc6+BQhtYeB/AiNMfN1GnvgwOtE0Lt7/TC04AFzDbnrvGCp
R3FVD4D3j0H9SWMp1+4oreecgkaZXGWn9BPIQbXqIARjoN6qrCzRc8rWiRMD
lGqZVZHBtCyZxXAHFLl9IMDIi1utZ2ojZKzh5hQB4Q2nvddJO7WvKHSQvV0B
bHJk/wPz3IJPO9yoASAfEFoyfLMHdj8W+Hz8296BZHSN0e8mi8iQRO6nsOse
3irDxq+XhOiUhLVB0cdTyJlz6qKF0GM9mVDPlgiM/JHnh4kx8IMWqZT5cxif
NkmPcp68uPsQqEa/d2WRiDDNCAbC6hYuVbWx2cr/KiwLLX0E0cH0BeW+PbQ8
rROkYoUMOOyckHhTFuA50+lV7+fscq9Tv8HurOeznE7FZgkKwuMfdI+38AaW
FeTe4BBNXHeXF08pEEj+KCp8VAi50eyNrkCfwXzB0KCKG1jH6sD92qFZkFRw
VnGw/is4cpgR+1UElImi4wycszg9MAiTgp6outmc6tkGtVAxnXGmzIse9ybl
fKY49FNTj61WYHpbbrPBgblqscxiVMX5VJ3fMqWticx3YTERUPiiF+TeJrwo
ZXUHNqGh4pFYD/MMCezemYosJGe1FrbFk0I/KfO6z/WRCJjNEiHKQPFT+62L
TR695Ptx3KW22GthdXscAHLpuecAmbFeLTLnq2iucbV30/SIcPEQ61u+KYmQ
OcV1RTaAmYVLzucMOKOCdaQ79pwnRkBjuYtrTjfYR2MD3x+nIUI+Dq0wcZMJ
6kCuHLFirCBtlbl24fF8MFbJ2WRSNDhU2gpcz7etAuAbki+A7DAS7C3pvbjG
zYCtIY6ChiW80TbYv8Nbr8JpuclEK5xkDcHVg+4sctu9rXiuLog/rPZCdKdV
UHp48g4eWQtGNlgIUb0AT1A1IYEwDkzpkkVtm64AEo8NiAqXEJmMNn6yxR1S
3YSPtgX6RhaS0FDPWii5vj9pFSIWVH7MIVa+tpcZIWrxcD7KwNEvwLL63gWC
1FFO06w+aQzb0xi6VVMBGYbE/puQIeKTKEEgwHBD1MGcXL04R2+9LdlFiuof
O4XTHraQ3jZb07wACAiAc2tP4esQ5TnJglRLLRMVmuWK9OIAJE5G8zUGmLYD
jQdK3XRLdcJC+vb8jQyUdfXHf8j5ZFuvWQX7O70U1xFJ0A8Jr1/tVEVy4ELC
A5IvmSFFClljjRNCo3XE4AqMwLEJjFhfJfqmHzptYGaLweJn3DCDHpvrBrhm
Gwmtwpm7ljrYryW5jqCR1Wzga19u12W37a1JxpKrjaUY/7GgTFh92+SGsElo
NYPPf6Alyz35QiZang4qKVw7L0WohGP2KMrLrNeGdbFt+rZZcI23EEYQMSTa
tsSBxwHMafuIimyejd/afOtNdv5IaPpE7JJXMuZtHrRiRPjJTzTlUaKg7ews
/09obYzNs3/xOKSbgSUblLO924iRQzYnDNMF+x8QpOVf+SmvnM7bxeDra5Xf
012RtI4PE0eQMX903ILfsA9qzRMVN0mmaRGgJrEdZyfj/Ak12M2Oor52nMq1
8xfDe3rh7Lie7AEfUGoRjxVC1ciPPIrtTy0/G2GaLnTSaQU2DiG7DkjArMl5
bKK19SApVHbwDLfupGN+iEnMmoNVNFgPnCDdJ3Y3bG1+GlGWYdp+FafdBaYh
/oDJ4ikCHxita0kMTTpiOm2Nqp3qR78zrK7wkeUOjpmQ4/IhpC+FprOJki85
HuweRhbCP8zoYYWvWtJwqustS0IIpQBkAAZRxoxgoBy8lgXI4LjQrSKpWLVp
FkpDT++XLehpI5ICmb9Qe33XNYIIUBMxqqwi5EoDX0oGbic2m2GoPpzacYD0
0clL4lsLa1dWi6h4xk8dX4qCUKrLKtqKALW12HFCRWLq6n82TxlUu455E78g
cHxJjxR98CTbqn1rk0fIKEjvpwtwVv5+1WczCGWc7FhmCT3tW+JEBTqC7uLX
9F8Ooj+rNTbAuOidFRJmECgxWrk2GqmqojCnLcsYKHE2+vq2MNnq/4auqreD
qHMbmEfIeqS4sGn2hrUareaS44IKD5WekgUhUGelpf47hBQ9WSOD5swrOZIF
h3k45yewLF+JFFD4FcsOazUSHKDagv3RTilNud4D/cHQQEvSMwW8z8+nc/VV
tfWbnzYLtxlb+UsHisTtxon0gQCg6z5xoCG8pB8JWbV9/HOJjPl+5EoQ/Bgy
sbEoj2bSAjS3Od7vjLsRKeq2cIfMeBd+LyopevuaprtGO5ysimf1AeTqVhPw
6KpZTysu4h/q9VYZIaLO69Wa7PK9bI8dcTxUwovbC6yiJi8/VqD0l9t8UcO9
g9TZnE48lR9omcLv1K8P6yTNV3p+fO7n2RCXpUaqTH/Gtpzrz5GKspypKo9d
tpqQsc8JN+EwXljHjJc2LgJjpAA0zDsmeFKq6hG2ob3JavfDZy2HOeZSdTvE
9UEfrKhs6SirXK1UJRK3ekTWibGr5rsllKSqJx89RMHrKFaI5Nr4uzGV+14U
/VOLraa9PC94hKUjE7ZYZVKwDM50RQfWjG0jF7y62fIlqD05LxEDSMTrrvO8
v920XCAw6HkKOk9LrQK0ovob2B0VOV63CblUwJuH20ht/jceWRHvHJ5cEW5T
d6i8V4SUgE2g90/4dT9j0uhkv1FkjG9wYL4cN14KmBX7kHYBoX50lSF0Kko6
O1VWGKPU/49/uM4z7A7MAMbhOJPXVFbGcSZlLqEiAupyv0ZGp4UgkQiXcGEh
woM0XjjQvQX26WgPOzFbUdxLSvrH+MUT3x2/NYui7RhT+lbejapAPgZPNxXe
Sz3BrrAlhPxtMQHoJbbRgc3UjRt1t1qc61HUMeCakBA6pdivBstHhcLJ93nF
soeGt9HTkuIaEioPoY/8GCiBiUqLeNegxIJj456VQ5FmAArnnJT0+z61Nl5n
kCCBqQtuldegjeb9hGy+Gc3HaPR6cXZBad81sHG0X3VzlCY0t9cFR63u+/44
5b5pUOFWpaz69Tm93Ibyo+SLfNLJ4SJNLgjID9R4LFOiA1ZKwSUuD+sZlot2
TILfSbSaBJqEg4foQqPsvC/CsB0C0EycxGaKnQVcRgXuWw88ZoZ+K1xQZjR4
J47N4AFAvdsIds3HWjLeOmFcS3MRZ3DWsAKYm20skB7rgm2lhZSobVYBn6Us
QqU+FECOoI7HVrGO1V9HgJ6PovTpifamIFCf5oVuNRwpw2P3aM+Y0VBxZmmP
ZeZYe9D+IpGGAkggODRw2U1ji05NBtwpPYGmz6jZHqNw/hhU4bPYHMBUl+V6
tZfBFyWX/JOZlUBo7jlFwZ6sGcQVy794h+qb2dOKTFDkMzZdWXVmLPV/d3ed
SkDW7Y0iggn6mN8X3cn0S9cdsZs/G5vRYNHZXCY3giZSC8tOfMSW+j7v4I7k
Ij4icGOvbAhIf1J3bR3z6PpHF1JJuhHAtdvxN8buQXQU+pVDHwSb/PmsMnLS
YCWJU0asgQjgGNLORyAOUlr+ni/shAW+2ZMPuP+99GpXW3e8+90RBQaqeuhT
WKs89Tb3EC+PXru/5PxyihpI2dgseolR8h3IsfiRheNjGQn3vAC7FGKjwKPI
MOI52ZiARdbwXLhUHVh9S1X9V2EuGYT3LoiOdRwb3tsfag0cRW8bfeIRjOxm
sww8xHIPW6jy1c4bhJnl7PGSu1UbNM4/DRgfJRPDG2AUMep2IzZKj2ohJFp2
b93LvhtP7061OyUPsB55r2oBNdcWg+qv08f456XzNVUsiceLeqWuDEf+A7cV
cpFQFn5uKnkxXP9C3UAj01c2r4F0qkG5zkXkG1p3kODoOarF1MkjIPc8h3n5
LLLunU2Zlp4lwW8dYNijBb/0WXA3gvwv/QY1Bg2NpEhIG9Ho1HjDdCuRKsHM
eM+6CwKHq/JAXKbvM+sSRXHDyb3wdd2Rkiv/eGitBVLYc2ZXycDLgcz8TBRC
w8TNU/oR735edTMUn+ijOUaNodj+OsX4DdFTSIFaTNJRnGqj4DXDNvPbiRrB
TcH4q6OeG+nxXAQz1bIfBLIhY/8uuyPF6K0pu7C3rFLReue2fdGiMQyiD6OB
rEXjQ8jEVuNeSYjsOJDZAEw/fC3YBUsNSfckrNrh0UtF0anl4eLcFwVYBDlr
C7Y9GoKRH0GFeWUiV3z+8hpryRFrl7nAp9mVAUK0UIvP5skA0rxvyyYNM9qN
FMzX+xLoZUOuB+t0sZq262TrCQUK1mEiGgkiT30bSciFXEoEpE+wkM26GbID
AicP6YdqhMwfCFV1xx4b3ZPPdul312ClKd5025Q5znZnh9Y7fzH4N+Lmj5PY
eFj52VBh1IkfPOQxsj1iBm0qcF8o5GK9W4rPIwKZYC1kdaIRnPdpWA/KjRsl
YwQ7O+VQHzX05y8Sgmm74H4frUlsmBKXnDs58b3pRU7YCLAUhdCPMHzqaRKN
FfafhSmAYelsgW5L9AGEGavFnyYRBoalWMiXTMci3Zace7i/z+pNfieTYc+9
G7waoXYCmaJvMU/md+uOGa4yJs6mfM4G8R+u4doHQYE7kBDQAg+kUdg8IjVx
JcFXu2oK+TWay77OHm5la/CfaRMhDx+xOoFBxifpPHkSMmyYdJ0vq3dlbmVB
OuCjB3VsWqMGWTXtTmYZfgq4E37oBXlY+S8zmkK5ZZR5aAkQWPMoirnfZWlE
w+3eQaEAUJwn0yjy5OJ2ARelOAKNhEORpB3kYSBn8rn2/CM4VKHmfAy7RufC
fBwI48DEKMt3ATzvMy5o4000KQEaglQrzQtBdJ/hFbr8u17gJSDv/DdQdOcO
y6nPUHbP+E9C1vK4em8/kI7D+xR/9PiHbx9YGrTaQaJ4SBHsG1DsprU3CPhy
WBsmIKdtwWOT7bu6dZxcgV2awqzx8Dei4YKGcgdTG0U/IX/zLP9C2n3AHUDH
NGkInXgDlccn6a2AOnRFcifQ0c4c4AFJNyzhWbb51x7Cwgd9vTOh6Bk3cXJI
3xYhZHkR7MccUT5pEs8JuwhxrnvxoAzW0PtGmu6sMhhI0bB7frAsmOhaT2Af
ZBGG+V1WRWXuriaaaLbpP+Ooxcvh4XeDNLgX4QZJdwgb6QBqm/A58a2ZVYd9
AZUmgRtPu/AJqu15MOk+OTNppCT+3LR7KZR11eNP9JP3GP09gG2zaaH38kNe
D/nhigVaH1mliyPMOOBQ60CCvGYDlhpkjz82xk+E1QySLBH6S+v2FOCUktYV
Obuzjc1Ikvxw5oXmrNmXnCdIIqEZD2C7MVFVPlDNWIHTAdlvCHxVzB+5N6sR
ClXD3VphjdjDs8Xn9yirhEjugES2X2mq2t+LuHzdrxXycfpnSMZ91++yU706
Q2IaCJ4N4LclfYGvfBegFzSskDYMYUhtN2E0QlEOlQ7r821AZEK71x0I0dLj
H8lMe5a5bMCbRzEGD0thvL+HKLiTlhjiqLjUINElv9uF2j+UJnEr+nUENQLr
aWRyJYdPQW4hX5pDvFZ8U2qfQ6K2qmFkk4ymyI9TFZCtJKcT9Kay6sFOHEhh
PSzj2ai3RrqUZVxERPR1lCZvLcf9cH9QKWju3VOD4dnBdNjVasb0BcqBdQRS
6v36y675LtVm/hq5qzbRtGuiHgKJhCQok7qFaFG+xcPVrybrbEQT+SRN5Ni3
caDtZLPDbh2gy3RlCAgq56WXz5C7sy8GTDMOTIjVw/YRtzhTqD21HwW53RNw
Exlmh+dSzINT9y1QwR7Toe0U1GJqUGtIjTKeU+V6zP2W4nkLu3LSIiP3Dwfo
CMYdSbJbY9ZwdZvqJlOHCEYdVKDXaplPLJnXbZls7k8F1ttwkOg+fAoYGwwn
qDHYPCJcLJRJsInt1c1JfeXb0naVH1pbhwN1dlyID1pg/GVCyB9NY4D33pTY
AlXHEsU40vw386Tq+N2uiB6Yrx1Cy1dJC3nAs40h2H3CKbl+IaeAHJ07x6c6
/Pdp6TMGL6hLH5GgaPdt5KOJDza3DhwQoalE+m1gxwE6kyW6v2Qw92FlaBgc
kq1LUM8PKlSQeuFJM9DatRaISwzr4q2O69nd1W0CxVX7E87094SS39NZqHnd
GrQBjmVWxOlv+fXyPGFgsM9IAAEwUg9AGQtzvQ8TBukols5R68enzz9BeIDT
8mjKWxv702YQCHP9TNXQs7nA+WEfzbkQLKWjdxWRi365xTqZIxqi+fb0cmpl
fIoEB2Dw55adujNpmC4XnI+vvXALAY3awxO0tck0kc4fKuBjb9neoVCMMS3G
8B1IH+FrGq9ffD0CIq3niFWvpVkGpw4ndy1pV53j2BTsVvkXKaLTYAquOM5g
IHCqTBh9HRJi8jD4YSUl3Px4G+cvu6HQ3zgqf/6192QFqF9FZ9uV8mIC0nfj
q+TmK3Fyplmy4TfvZ4WPRqHd1dKlVlctUlc35n5oaqKreyWC2UHUFgcp65X0
ySZCgrn2au7r2DFnr8CrmwpJjhXOusTegGFkWqicy3IBP2ESU0L/knIEvJK1
YoJ9BFt+73BPVkSLimrLwpDWb0u5Eip5nd5f+eoocvYfHKgyI2sZJzn1NEQ3
cebQJ5LBe1t2q3VSZBmKHp3sku+JKLCOg+6mruqejMMufVbErGGrhvaQqUyo
FhQjAArhRv98PiFdjR/xcYtquQgkZMlcJVIPLWaIjaJpeworSsOFmADGypN0
dbhh4B4J5aKz88ViGnyZ+Mavxud4UMFJSj5XEZG4lrS4O7Uhiz54Q6WtHN2h
QUg1uhG/QzWKVaRXWVnptcpDwmWTlQB4Vfj1Nyh3uLWGWTPkTQxPyu9gyEC2
Xyw52UZLW2h6lbFRCNaIwFnjPd3IKPvmmIESHVTqPbZFHI/6jgi8wKx6p1Gq
gbN/IwSO9G/ajqHXw7vkp/vgCPhRMq2uP54WTqqWOmcavAlD3wCYdQqq3xXb
pVwQxCCtfJ9a/qGLrlaaQS8UN8PKdGyrOXWMJ06pYoE1PW/7YLpBbnf0tw4N
WDAah8Ot6pczd4r5osPVGxW52a04l32UVC61Ba6KWzuc9v96hP9Dvc71QTyq
/mIIvqun28Ponfn8wQ/HzF8PU5DrPXKsPDzCcK02cpRWKGmkW/LRZVYkr9jy
Vilan7STrRNyGkJXzXomYwr1mRzwSYagx+LiYTTeuZRcrivGZ+UOLcT9mEuA
QeDtgb7uuzHPM+7i+M6jjn/bU5nEgpMn/PEULgoYHkg1XDGfov4oiNC63F1h
sT0dltHZf3hFx232Ge3x8PJ4XBMbAUjsWMhln+KA7FlX1O946b2uWeqDPecH
9FyNYIlwWK/U4e+1sfWHujzTnY9wgYqIFh25eCGIOW1ZV8R+5WZmklnkg5FF
WfnS0n21EPuCUM+Yuj3asGWHFYI88Mcq6rx1qCdwUwuQ2ctGPHxl9l+Eslna
SvLDoIkfdR/PGGQfNFBWo15XxOqK/pKA77QHfvXFGSf+1k3f/lqmJimWN9pi
uS4QMPMfcwCosKTE29CVOA3cY/PGwQiG5qGY7wI/fikq753iMilQHRbKQKIo
FBuLTTvDye2Ysm16vYOMST3AzqrJkySXu1JwBswCazMedMjSERRkro8Ghi//
V2pQLRpuLapSMIWb9/+NLd2Ym64eKkszfCCRp/Tw81MfR1bkQZU7JaqNPPsD
GG1lxmeAXEIevtA7OHMdtEE+1PsyuTRALQCkL1MiM1mq/RPkmGhr1tjnxeec
hymP1E8eHjdXpZg0QK5BfqDAJg2s+SgRaVp/KrRqbmqKbUkzadYprwt3bMA4
B0z3WLc4vlWfzE2sz/D3t4mAutR0FYanIgJAayu4H0rN4HFkCrvvRXoUMpFR
lFrUppVaHsvuyh1qvum/BAU1VwnKA99bCQJcDUJ0Uu9AFkw7RX/LhmXDCzZe
74LzxqgtFwPiad7YvLMIT2dSXjSLYFBNLP8SdbbbsiF186CCEEFFkuxubp8n
DzN6suEU5B0RAVLrKvP/uFZ4bgqxTVQoIvAOU7UnfWvIV2vILF9RwBFEkNlU
SQzlXt1F7LndWacUQaCa7RZOssd3hKmP9m6qV5itBAcKjexmFady3VIvP3hI
Brk4a+fc8FxmYXMyLVehQiZTPmJhW3oKl7y6+U26ZPHOgYLxqTpRqZKaaDAy
PltdXpOTAAL8KSIMtgiD0AiCTmTklHKcEheuFz63/XvETgR15qq8jyTm4jxO
uQ9gQzDZo8xlTY+wjiCgjvBA7MGXYEAl2oZ0oCqRy/ro8jcXN9GMs/We7TfQ
5skjgh6060MjarzJ9iszJT6zV6mMvjKVR3At4l0vFCIx1YbRIwmLaFjpHGQu
R53a1rlhOF2Bbhv0o3eiNprUsItT2FeeLD5C5SVA827n2whs8VyPqftBgzZ1
elmTSFqnmyUefWcQ289XtLr1HuRn/aah8FFzuFKMZTUYoyE/h5yVkHOqm8r2
G18I3sB+JnL3SQnhfeCzDMGjkzgtaUy0oEgIwDNFqe4eJfZDq2+yZrD/+fAf
UQb7gaH0BcFMc8VrPFR5/n0piQmsq+llmIC0fS//QI+EhHDJ8bxFPE4taFFi
yObwdF0/3xOcmG4ajnXv8JhU7yMBhstqCQVgh8QqWyr25xUiJHzVyUtePRDU
+opV3y+nMiNpH6jZtOsY2c9eoVmvCpwrWM1zvSi7qyJ1dLOfFuEzlMHdsxwX
VY1rH6JfLVLuVHAmZAfgK/I2FYZhx60EVrIaHiniLQ9ag/txFiRGK3u0POZv
kCtkLj+wiEXA3fEWVvGHHo+FsX9QkMlUyq5sA5a88pisB6i4FzSdtXVTxuO4
sUHh5Pl7V0lhS/Kc92ogJXfUvW7AWYm+ql8Xt/5zSSQrFge5duBJzeve+3a9
/6Kic187kCw8XAZDqWzSuhxgDGCfy74JZeuueqBDnrc3O+kgMtfinefHKuoW
9lOeHLqZoEvYLRFee80tHGoEP6obCPkkLnJKa92bZFEX0kZrI4lKEjRIYtaa
PocbyOxsigCbNyj9B7phfDHOMuZPIafKgvhSDMl3myKq7tz7to5PjiXEoozY
ykjKbccAnlojejuCPhVk4xk06BVv69NDUfgw6U2pWCWuErveLRC0gSp3dlIH
KUnCmn0Vp5G4MF7I+IRnapXeODvXmzQ3vUXKGvkfVmA575C09dAG7NPGEvk5
rv0oZgTlm5SiJRPlUud6o04I7hqbpN1yLBsZC6wO9vtVUXOVyjCFSirRXGUj
7vVEJlXZXO5wb50dQYh8Q7CxbnafQogNNgZsGehtDJPuLnmWmwsqBU8yvJkL
MJ4AcWzIRCzZNFua2M0b2i7RyQZkFrNBebKcQAuAxo1GEmhnIbYueT9eFW2f
WaqIKnfLfIJYafQae6wB9C230ZaY+vIjMc4CA4B56Njy9adD+NJnEoK07hoz
tyN/a9Tm+Obmly64mIO/ywy270YKii2RpO1A5LuGxZEG0WZgALe3OCf6vvdH
WMV3iKOnDT7u7iq+8uPkYVKABIjh2HsidCd3PxXclAUEOeAlQWWSIoFmMj+W
T85iOR6v6IvosqxpxZD0gM8/2RxOU6vKHFfBaieoJ/RWg4yvIFu5DgDyyai7
BbxMT54hM2YdkJoSTu/HjoWcbLgJIcXdE4BX28SY2ryCxnl9WtzXmOgFJEn+
QDIMKMNwNj9Nw2sU1yzNaeAhxXJWwrPA7udwAQg/oc3tSJ9r0E/nqL5+z4wp
0wvsNXu24CfXlPa6SsQjqXx3j6pvJHqhIQ3bh4XUdAD7eKqc6r0Rk2f9QIbC
sDh5lz4aV6TsIVQhDuJGXZgqpPnFmp8ugBcXhXOJaEhXm8en3NdKwnjdwU25
/njAyaM3oiaYWE1tF26FBE6+Ek5aJRTeLKa41uBMDW/61BO6gRdshrakvWgt
CwobpWrRc+1NpXQKlQ9dnVnIG69wt3z7kraXSOBwVbNh6pEIbxkP5bU0/bk7
2m8OxLplUpxrUGi9SqSc6tuPO4Fv2leuPFx2PwBkkRSj0vKE6Z6I9iYqKuO4
nKhB2kpUqgxFOjmcYmhS07B4W4Knno1/YY6j7VQqs0+ws/GXolSfm8NgJGa/
uZ5ey38zc9/xXndm+w0bhwhdM2+RmoXFU8abKd6otV/FnpIHMokIH1rcVtIn
Vj1wkwzmUSLq24fRUvRQT3OpJBqMnKLj1VlFeLSTfOroTWiuMG1wfJg9eVoN
xmn5mD51b4sahgfYNK3CUawK3r+Mkm0f3eF4fU4qdIk6couvdhjj63sx8fmT
wyUSNm+Dodock1fuW8i7x1alJ7cOhswfWY8bDteyxFnjhv/XPPAIZZxZuHTv
ovRDssPenxDJf4ZDkoD5RnD2ti7+licKuYig63pxVrteGP1MqJK467DMzR8Z
3f/nt0OPTMWweB4gBjeSWPu7RQrkhXUzDN9Lt4Nnu2XeX0Y0jLlq2mFSDagQ
WjNAOxR/xdC9HIqmabweo5BBPHTycEvHymSuo2R0n9sZZYwN1+aBzudvuTyf
edaju30PDIjB5F9OljbAXScPkUotxRwk0Ot6qpoch7sqQfWp32cWaCE8pVJD
qrc/4LhCAuT44eQaMToDRHz3UTIjjEzoLOGVfkLE/V+z+A+u8Z9soM/eYZvb
hXi8v4odxN79LH4IsGVMiVJkvfvghwA0L4A/eN9R4CTXhU13wDhh1mvYyFbL
AEA5NzueJsBuThC2TSlovCe3PZas0mM31hHEjtHmCe3nK0nYk+C4jLExVrCS
Z2x0Q9ArrDOCI1q006st/14NyWRsLsZzVwq/cdM/1rThGnaR2hUb8+QnKyti
YOndLjDPwSHJlZX4moKg/5UH3ysOIMJnpZokwH/UldOIpJERTwltv4Kvw8TH
fvU6bgsiEyOG7hk1T9S00I1ZE00nASBHELAYAeiM2nplxmi/FZhpeTO/QWlg
tWm3ENycr8BFNVONyqbyz9XAHza2WgTZIpwjfDY40vKnxCXYiw/hK/cWqMa5
+Ik8VqhU/YZCCfhm1ecxhYh7dxDI8fM4JC8CVgHcLo4YOXtoEdffEUXrGRbu
IHToOyvA0sAR0oFGB4IIRrYPUvHViPxwpOMXXiwCXyrMbe9C+/cgB+IoyBZO
dqOucA2x5Ix025+9Qc8WamB5Ikq4ubuKb1qdA1zCXZtbgdKToUelT183c0QQ
L5x4Mej+PICLtUfM9k1N+AX4sMQJEnHLNba+tcphYGz6BsQlACh/l90VURSR
UxR8hRjfb9bVppleVMQR15PlWHk/1NmBgp62AywxrWs7Vd7+7ZJZf6QX6NfY
KasKp6hb+YRPxM+eOTZUOwNAh6S7KzkhnDHWVqA7tq78nN2t+0DXpDVRFZeU
xwC5hmC8wO9Wzr4ZRYG2bvE3LMXWqtiiBuzSDutciQOIJLtNHZlD5NxDXrJo
fEeVUc/8crzL4j4TchjFF/mAS4lu6HHiTc1dgnG0Yj6Ojk7hqpM/uGtOLnng
hHndWLz7N6i9uvfaD1bHmKgRAi88jQtfF9NgaTwN5bg73Z3HjFqpo5HKsIl3
07oIxwF+5AVweeIfghX5cbBbx+FKEODXPf7dm2z0Tq6RLEW3HmwrwxE49vme
opd07rwVo/MvOLulv/u8uwLLElVwQASGfzZahVLtlxfyTN/xnu28SCqiQbKh
YuG3YwoltoLTkv1IGSeaDb6RqQCJ26KHls9r8xxiUzTT5KBJxqG9jwTcUSwQ
fK7iSPsBZo/Etq6AkxfFERNT0FuGYXnfGM64pPq99Juwb4MRdE924BoQqmln
xXdfhfrva9tmLLD5r3oPSQBDctvHgXTZpntzuUb7XS03OKgZPgUc5ApbOj0j
eJJWdirMaf7qWwvRVsMp976sSK3tXFF6Qm8st+M9BIcwEnJxEDMDaI6cAkHr
l5SaGnkl+W0xljT5kD+U3LM16QzEw+Rz6HK2R5wcjt8rHIfcauDdmuZ2AaHc
hwrPT96U25egcenqUJpHjhHxyR2vu8JdL4dgxro8NqF443+GBtWW3mPATXf7
B96MNTDohLstlOgjmfG57kAXjL9cyTRq8l0Iy53u6XRxozIn0qoRY3qAnbZg
JO4qpMK0TP3u0ncD1BIxFtfJUoJ2xVV3K9c61SfrasMoo+C70Fga7/lRCb8V
+GbBUh9umUjJj12mbJDKghmN47hlMSybnli1XvaZURxKF8mt8HcEJ5RZRvgC
RnEP6IWduNXY0igCLy0o6CeZupOc5CZ1haYj/A14jy/a0jK/OOTIqAKntCMb
P8zTfJY4O2ivT8HV3kLTwk6gIzFOtS9y/0KtJeHTLBQxd3EgqLVv5gzWe4H4
uSFYo+FWOIM8weHsCLvE0e4FHrUrkD6MHTVpESmjWC8xvUp0mZQghsgHUIvf
8lRnyZ0f/X2J+Fsy5R8SRJFE6cZVdKV/AecUXmb/BNRhruqfMim7WIUrQISC
TvvNSfYsZQvYbt53Cf+NEVTkhdtfGAgpacWAhxjxKOUw/pwzQffsMW8bmT4u
v/gf1a3eAkSxoJFOdHmIezf4eFqhdkZPLbT7uvgTIBwcIz4qUJ7i0EWWv9uh
gKwQgy6O/DNbLU99CJDFQA2ANTEVaRyiRGqDpRU04PkfvdSY0TBq7wsEh39I
f3bLCgj/oNbVkWUCFEZcDp6Ovld1tiD2HWOOFLIlVfPT4c3PejHkvpjQQB7C
KtkmEjcMP4PooOI6jGst8NQU2T5ywWS9wtzG/1JApEWJUQkLF/d2mEuC2La2
/e/6qrVRa3SGbdx+A+Y+T3BHTTGC49fSDdXnQIh6NSG/UzOLmOsVwVYRgVxL
S2pFpSwAAeqq0AT1uEC6iwN0Q76wCtVpM7kTcd+jNT+FBUPF70vnbujo++0C
4TrZvNlURH3x8ku9ijzvjDtJ1lF+Mt0JST95DLz3dR6iOu4lirwzQIwfR/3J
6MMtcXqfQM/pSuTB7oj7zLEvttiywTS3Xvr3K2ykfeRj28Ama5sn/RNelnpe
Ub1QTO8C4oWU21P+plFt4myE/pAPTWTCG4aXdSWJXFayotmqx0D1tjLWKeuH
Y19WON1+acu9aAkug1Ec56+EJ5z/mnuQXqmsuCO+7JEY+KRK/qAuSCY9W2Gm
mrz77P46FGCcyAksWQkSThvre33xzEDaTybRlqiwtoywT9buNEmm8jTBkZ0x
Gf+4pfbLamN0R1mJvoVT13Liv31wmtCp1KrNg2Ug+dKCfmD1vggRhjvuSP7n
jXC5BVr/X5inJ7SeI1hh19/+apuC/oarqo16a/eNLuajsY3QTgLEBZN14IhD
fFmneuY5XczEUqA/9o6iE6RlzMLJVIjrCwJnTcG0UqjiIEXa/1JceLgDSgfc
6K9m9XQQb2p7AlYZVZM/EF8/3VW+abuEwppYhV8OxiAm7OCT1aQYRgSBjWqB
cavhvn16ElZfHCXGlZe7J7XvQk1CIh5PR/AScBHin8pXhB+2KXIleJbFQKyw
mB1HG5UAwJBz4EcdYc5wp5lYp1qPLJCOGFhQRgoow43qIOWwGv/rUfOLTrVx
5urINsKv9aphtfjm1t8wZ3zr1iYRpgjO6SDfMU6NCB2+k3e1Kt3kDBql2Fam
tXnr0NTNqhvIpnVn2tIhVDwWG8NsBYNKVF6f5KsCnZPHWyrxnifmou7goyRN
COBvQdn0gWWVSmHYXN/CcAxIwS49x3O8zuSsPNLJiri1PWtZSBlZsePiPu0Z
Bsb5aaeF6Ez+sK0Hp1uPjqEE1agKRFY3lCUl/Bgz6MROXOPqg+VlG2s4nIUk
M5gOX8Hw8MU3wlWCrhQ5ohLuNAq5aotxVTopc5PfoWflMOywlBgqNHEBB3lO
vit/JUrnnxn1Hi21qN0l5bon/sTq+MFuAeMprweHVktsYLQKvhtp5VuegNKO
V2twojUrUyWXx2dDD5P3OSlA+U3O4Ib728QXzv+svOKhTWnhGwkHCLE1WZ4X
skMxjiX4wdtaOCmqbK/uyq8SNAwQxYGvrbDqZu5cUl722SmYHjekkw1MPOzV
eI/Z2bixEO765QiHk6aZAEmvz9N6CkvmOF+jFgUWL3G+gQ0h8HBJYWiKQ8j6
hrzEdk0Xk1rnQika8uJai3Z+RuJ/4Dypg5E5ReR4VDkM9pSnOC7gDOz6IlFT
8uX39xeYKwPuKca4g0XertAv6L0gCsA51fHnZpm8EaIngUEXbQEC9EBX1R0R
IfAm478OGad08o+QxcWDziuBff9c39XWBqLfOtZMm39C1f9p/kwPr7NUN2aI
W5U6GIGAU6q00xD/2Z8NPn36sBEzKO513IwBumGYeqrK1j/UhKUBRFo6rY41
hc7cQr+MuhtmpcRQvYmcbBwUd7A0Sw0paMaZ++jyQCUGO6vXPalDbszj84RX
UHyJ7hBbwfLW1vS4AWnspsXvQ2stA6dwhLIjdY1ENvGtkKv6ahXZ1EEXF1Dx
czHrIOL9r66vOuAgNmtG/NfdLXUpVHEvf3k6fTGjRahFeO1hWxlPa+2R+z35
WudOrtTWQmqxA0P+ncPCqpMkWK3mDWjDQT6ocAB5tQQuTEu9B0cQQru7hApB
IYT6e2RqLHl06IIzG1sUhk+FGTRDGrM5RwHsszvjogm1oopCUet/RWzZwI3K
veWKz5qzeY6XaCX4I8aZbZTMTdvLhfDsNHzlEvFOHgsgfqfFr5YoxrS53FDQ
18jS9Wswu5jg4w0gGFwpfKZHY14RVail9pZP5v2ZyBfH+2OrSyMNGThEbGQ0
VQ9Pda2GImhEitHWq3pQervqHAi6nVTOIspgW+zIvQtjOTZzu2qFCw3A6WrN
LHhekLXuQZ+6omw6VnbwUlc1S0rNm5CrqFbV4r52ExmxQGrKxneI3j2IWZnT
ZejuR187He6R1fZXsMd9zWHCzX1lmsb+d3VQ/5SScR3ex8Zm/uYyebMiSw4o
ZXSryvteNgNNjxpVOkjR7F9ekFRjCzmBSC21eK6fXL/ddYQ6ljMFx7EQrutg
3nSA+l6zLQFECNONAaIxZKvHiKW4fjDaAqeO21MVxQgewCur3aCNTmhnwtlz
657rrLUVK/94Pz+KkGQbIugXJMGf/Eja4/43e+U3NJ3cm2kHKhFyu7X7KGny
6KxIKOjvD8dgQAyszj9e4gor+KP3MiEE2y1JpwuYJJiWzMYNK+fPME7YMsb1
Gs+u8/Fp659payndRm3EJgpWjBXT+zbcClzlxcGM2CPozM0o2xV+jdmDKoVL
4+UodwivpY6O6OBUp07EmyIVW5pF/WiyX7Xru7QMQc8eAdoGRPhrNkfh3m2M
ZV3PTiTLqNjfabzXSpqSDl675zsz7kT//Ct1kEvC0Gn13jD3XehP7EyZf55V
xaOzCsh1fscBoehw2C0goPF/lFTqz1xTjvmiBQ6B5T1QC0pTtR2w9wjVets2
kc+2Izk+Pp0Qs5wTtlASvGRJvbPeNOxwJWQ2gm2zvnUcFaTbLdpQF3ZFBqHy
4vGlQeOjwsaShKQAxCT1ydzsdm9nw63fXUexoZKRRntcTCV+JNSJ1zHXy18T
Wt0XtSRiz7knMY1aYlImTPvXxGF++ze8z/tnNob6ADd1vwp97W9upb88LlRF
FS2dhmhf+1OghhvVVCbtPAopK2LB9pNmD8thEz0GH620SnwJUhjhmCfoNQ1Q
Pw03u90O2JVveP/gtyiBNLE2nINGk309NKvnTxSethPb2dXGKQgi7e8X9dKl
128wKhEXtcHTbTCDl8UzAbWl+JdghsEEvIo2tnaMW/p9/nSGKxWwbWzmV57n
DL4fFn0Rr1bL+lU1/ExwOGAE8A0DB+mMa4EFaBRUAgTWbvSMUKtFuAccxq8x
glia5PeUIMblVI893ZqZvo6ZJBN3TzkzOvJAaHuOQEQBtsaOs+emoegEYMQs
/ALN24oGM91enEXDPQhV5/b4/RbHCk6yAF7hmtcixDt1AckABpVZ/0KDomlu
4mJyAFCwjv5m12H9OPJfK4MgIxpfFWkL4o2LY274+K/JBo0rvPDs7y/cICnT
oZ1EA56FodOs94qUc1R6CUb9U61Y+3TxG3KjeX38YPa8jPm6CS4rB4/HljcG
Uihbvk1geK5hEQmAsxxFgVxN8cwH1BzpJh7LUsmDpaxrx/sDc675Vu0fdPGC
FAPyWyKoHQjIfsVg8K8H5bseKlEsxADVbeyMn+yiGpftCdfRYHhuckWuD7ab
fGv6IC7tFXcT7hmpLs1IPs3O0CGPNGv/eOJG6KNeUaNin0VvJxspMGwQYwYY
kAnmMGRZVobOrXrLdWBCQvIA0bu5mWLzQsAsNhbCaa69M7NEqFsdSR1/5UP2
ZP6Zn4B1LxDMtLZENiXd8dg/J8Io7VzHa+ik5Krby1r/fPVoSd17BFUJUkrq
4/WtbwxVnRbReJwnQuWiFaHqqeZzO+9UIrBL1YLhfp6u9pjGAC9lY/w96reU
Xiney0aqNkuhwIgRrhxayS4JeQwpEzoBq75iSYO2u499TjZc7e5zOWUBj+Wr
kq2+GpolEy4TkSVLUVIC70UOKwUXhOC97aeba/8hXSV0HUpUTP9MHkPeuT9z
kwqBEpQIsCwcjtbthFjHj8EwYxYq57EOoH1BOmlG6MqI8bqc1CM24XLlliCQ
HUOxhgarAxuVLqfHYKwwcsbmDLp0I8tlkqalXtzQzmJXxrOx3Da42F5XJ1Qo
z5M5gDgDkwfcDAw5/8fNOFVBl+pEkmpxD9cRVzn0+UqfageskTg/ocrcy7ZZ
y7o+8bJmYbJsZdVKXs33ftgE+jEwfzGSdsMmKCtXnlYlsgZUtw4B1308zfBy
vSe2jDmAXGQdErnUakylwzjjmI2uzkz0Jim1xApNeaquFFJqfGZiVg1oWolB
JPaCAzQ1Omjm6mD1b/PzfW5x8VKfAzIVU0jhYu+EYeGtKvmBtYTHm6bjhjn1
EhS1A9/65fwZOmljN8hOP6t0FBqmQ+tKI9WCHHrMVHZtjLCk6jj+xzU0TiRn
K+Q9a5jIppGqoAUAtbKUz3WxRIItL/fkDUbbKHfIPM/Vw6372Wwamk/j3wbw
ruM+lMNeNZkb6UJaq6mhQbryR1E1nLPYfVDjoCz7QvqcnAD32rd6P3AfSpRT
/AluCuUGRgHdW53iVeFKmlWOTw01WDGib2N7zPu0cZwKu0B6CxZLVtpg8LJ7
exCqa73y5tsw6D9qDI/b1//3iqEMlRHAMuuuuAbjMYxsKQp3XsJAFatkzK97
Y45v9vm2FPuraPzlxGV3sjBpnc4LqB12P7qhbS8xyfSDfv5t+jyPUsrK6VER
K0tR7RXAel2Wydw2MWKLQzZsl7ji+VBDrJE8Wf1bDNm46ROMbCId3fw+flb5
1wV5ESjAd5OZ3z1wupNomFgTfHC/n2O3kMlWgd13CYj2LnY9rd3X47IYo7T1
C1G9xl/1LVVwNXjpDrsOBKiVsXuR2Oh2F3Deoh34PN3Tk5NSAl9HUonUqy5n
RsD5PkWw8XG0e7JMQVrDB567nsm73MVTTGca0kRw2srLBwf131/3ff3VZglV
2FqQ6MpmX1PsV7N7LlDliW57sYG/8PW7A1JVr8tehfa3r45EaG6nCahm2988
bRGJcpw+UcKmlQHlYmFxs0ZvOGz3/JegOSYdDVaSP8bu5KvCu7Whw0+GxbgO
3WJk6rc4c+ZbQdC3gS1gRxKp6haYGLZ3UhoOQ5hCVz+HrjXXsEPQsfGnebtm
HIKUCuhoPIAB7oHL654xWiWCdwpa7v+I93CYnhCLcqvdF9M10fwnhdUMWGWN
93y4Ch1LizBFryrxHbg6wfQ1RZL40HCbEKv2fxVqVW+F0Z0QR5jup1X79d6k
QmfVVRqto7qRKi3v6fL8RDgvseRUtyUFAdn/YTglZ2E9dYQzn2ROFLwH/cG2
q79Y3TSUDvp3wVJio9/JT9U9cYwYnvYq79h5QHLfunhrNtCyZKXNVOQ6iiw3
Ssy5YY9bVtO6KUfY3GKmBo4Puk7zSVFrhEQKW2tZ22B2y1XdhsGV48vP1b5i
BvLpn+t4KqQcXYoxFlNWq5CGJ8H8ZrpzLUNcxZ1alWbuda+C2pwZKwS7Rmti
MV8BySzmjI4o2AXzwaYWMEdEEdSm89Xjlyl5VLxOCdrsYPup44S0LTjg+o8S
Sma8RaDlD4fayai+n2bHJZ+cHr0zlyQ4pJOcjA1Ab68a/rrHrIsuj2F+C0gG
KHsRWtzJ2oI3hFDqU+gB+kO0GxeDhGHywfA4Nk4D02eQCmeL4tmF4Mdxhuhb
+9OY9KaMDwIG5jedRJynvNTeYlLZT8o1BeELehY5Y3GzQanhvDWkZ55UG8a5
XcpyxyZkXWY6HI88EY7ZDWqJiYLQCeylQ7XXG9lFbCGA65rsZG4qpplXGtxD
0xAaSaLSHTNyPaMd0iDerBQfWvQj3VMG14nY5VBvaNtcoR45AWY7443kpjPi
1NIp2EM7o5ovnFTAVhuZq6ZnuGWuXptPMb6y8M8KYbn9s/Ga1nSk9iTpTlyn
UDo0V4ytj65G1q/1w3qEppuOmdPasUy6fwfryYr/9R3E0ZP4t04cktf03R2W
JCrfX+nNv3nfm8Tqd+2Ifq9IJyvobx3Y/dh1ka71Uq1SFfnA3RqMaen3/WWy
lgJD9gZFr4r2kxGJ/Kkv7Vrk1q10pMy4e4P5KJa6/sZ3ELs7MYI9X6aSwusf
4dGaRtm2lE0Y0MJHvW3XYBuuNCWmkPQ2lz1CUFTLvHvPpxPH59hOdy1Mg0Px
rXJZhexR9WkZ3opiGDaKr+nOU8UjDOshaSRKx2jemfh161zwhGppG6N37fZx
ZNrBZ5n86cG6wivMBbgeEjFmPAHEJPxzZn3RS2RthhQo40cYIkYzwiWOmcWk
iHQfmXhMdjIIxkgZOS1OM/VTrHIVWjRg8sh4L3NfLIlLH0zPiG9jSs1PdXo1
oHTFM0dJs4l+uw+BG6M70C9ZUO3PJD2QVx7IyuIiqo0k4+4kpeLr4e3SLy9V
MyJafujv8SAObPVKJICHlxsVDFn1Ij5/2osWtUqhycmPre9n+OCxgNJLyqRu
NPwikjcu4B8cY0PYme62elx6XEGvYoLgXDCC6FYHDTeQzywhAV7ifWNIZkeG
SBh3v30NDf5L9K/4e49pExJ2zMPu8BU4aVzq7jyMlhdSuRN3EfUzyg7S33K5
P20TSK6VKH29ZWiHeAnJE/3B87HmxfaM+K90BpoPiU7r5OOLgHfxXnK5InhT
UEPAJBO0nQB3ryLoIP8RdrfkypffihNcdZMGsUacewVmCJybkkTim6EzyhK+
U7pC4ZGX/3+/FRUJkyNBOOvw2UA6WOepOiOVf6xKubWZnLkQsnGFFJilwXtu
NCswZ83PXPtXYVSxs90Iq84UDEMEgnxi5UPs6TlV2tn16enIfizB4ZLSFWp1
s4Chs0K5xn5d1bhVBKPqL1Hdjwj6nMDLhVeX/8EejxCo8t2K8cJM8p9Gr7Cm
lisPYvbGkJkxp2LNEBDMrlnCQNLn9DcrJ08wpNlfbKdP5mEQ3o3DR/QZnU8L
IL6z4ti7j+k8yTLY6PXPEejFXXfFNhJexmJvyF04jaencOt2Fz7Kba6ZlLmO
8QtmmjzgvfFs3jfYq0kjIFKoxLe1uc7StE0FPZPUFkIuB4Knvy8OFBpXCHII
7a9NkQEgY9zX3TrZIumibKNxwhb5B4N5juhkg1eoUeCWx9FuD+SXUHhK2oIX
mDOyPcSWm9iHcro0VqoODrilgR3KdyMZH1IbLI4JWgeH28Bwz5SZhKUU0aOS
xaqIvEQenchOOLCYsGisS3beZ7larKpaMy/Uf89WIla/RVMFBMTss1NOpAgN
Zo4QxWCOK87Cd2JhUwazQ5p04oqd8a1sipXxka3v2jmVn6FZXB9Xaoyg8Gnh
17GQjRPjDkbLWBmUU8P8CFqtECr3zhsRxSdmGzI/XnWzF+CHnhtF6DqOlXik
XkdBgItvupLwnJn3QN7wc7106iOja49z7GaTVwyS5dWoHx+gUXCXF/83VvYS
0iiFrscMQq7Cxn+tC0FuCZdoZ0RHwW9/uhnhWALpQ0PkuIq05dUu/829ZJcG
eL2TmvkvuQmTEPVSJ5puag4aN4CN/T6JuPWV8s0Dwepbbs0X/T0YzF7f+ofv
3GpWxAlwYeHaNLOgy9kHOa0tuktk2RcLfbKd9rmqNlJZdpG/tzX4aMD2crGo
T0XG9kxoqlzLmbIQXy5Qr4EXSSqpHnVmNyk/S+grLTgde5CjzQTxr+lCS/zX
g9gJmK9SjuGGIVlNir2rc20UI/EoO4MDbn82R/YrxYxSnWNjcGFgbT1/H9yu
NUgo8UjxPLAEzPwnKJuAB071BX+8zLJLSybR09QF0sjY77XZ6ChUnWL2R4Ss
aCXalHsF1+cmV18rbgShNAmS7tJNP8UD2LaLJ3GKOXFd5Oj0Ii049twC6SwN
9MQVJ/j0ROlf+a0f8/MaHDDjW4sEAWm38Fu2aHh56PnMBM/LNt9nCtmKxc5H
fFXjdrW4PbeBCo5R+sVTePGQd31wgkxiFoqw/dVEZu53mg0fPEY9wVeQ8Yo4
lkBN83v/q9lRZILNarNmo/24s6KmHoItdyNHdx3Wf40i6iNQttSExIEY1PtE
XT7DxX4hymLg+YeOdNQ9LMqCee7qnRqD4Jn3pofsVvKceRo+Gun9JQkAXbOO
7qYMTtxgsPLQfQxqixYk+zPPg4K+2fOjkc/fh02XSW6EFn+slxU18vmFyB2J
iOjraG8iDVvkFhSuNc5O8bJ9HDA6eOpEbD0h5ncCCPa9IePWkBuT+C0dWoaj
UR5nbfRE0w1S/z/luWbWGZtZp2YLmM04K0j4TSLmRtdtf6zuW1Z4QibxJxt4
DyhSE265lmCID9f0/4JnN6nNnB/jm2dhrQEhQPZ4PNs5ibohsGNmjrLN5PJJ
sVxdI4kmwcMXvyrTRh7tkGhiuItMJs2IdySQ+J+UHbxz0BPYUODXa+BpMuwe
O2uBl5z659hZiIRIFZuOACYlRwd/l/jkuFWjMNYGbNQ4b7eUTqAyhhNs/rs3
MdeAf3hiNibCjC50mXqOfk1GQZHIrFTcXxiUylNg2lsj++XYS0qx0gRGzrnN
It2it6gpL0BsUXv503jIxCNoNytBOT+kFrEf3DqRIT0GSXLuXsDE07xIKj1W
PQVBOBlYE5oLO4xl92MTMT2tHgH39MhYn1oRRNiZmuT4JQ8Hn4nO6aAL02/x
fONDmwkR5wtag1pHkQpZAUh+1yoP1RpT+Ho+s6hP0yU7dLmxABf4a8AMSC8N
gCsf53B8BuWcPG2zdB1hlpCPOCeNn9jXrF5kqrmNL6MHWSem3bij07BiKC1m
06SYRYx5qfUOwzFx6rEXnovm6PX+ui2HQldD1drPDYKOJlYRmHsz1LkndSMz
rPtuIvZbI4ovLHLOq4qQpWYCihzza9/0xLLlJwGGDMBYDby5NfiuhZO4fmlB
jmWiNY5xKK0+LZ0xDPpb8V/FdHLh4FJbTFonZqdN9dRF92z4/GbQYRVv7/cU
wkByxGiGeuVGbCxwMNjMZEvCQchV0hSpf7mvkiGQteq2xmWQXNOOe3D/obY7
dqvoUA7SDnK/NCAs2YC0y8z0EIS+aqyVBmGCMDTxwOehGKFEKwhqAoe/WHs/
JbSYoMXd2+UeRGCKGNjivvBdGZzfrXYsDUBKON7FTyD/MnMLI6ebiF+qvBCG
HO9BE2KLcrEsdL1R3nCoYJMCZD+VlxcEl/1asEBc5VtfQN0mjlD/fGW7Xnah
3Eugi3/EDgJhkoWpm4QsnlVTYw19OxJ2TZ03qamdOT8fIDQGdk41/8AF5y6I
Da/zoJzgk9MnhKCjGdt+rjpf9QyzEvRfOn7I6EqXtkcK6ocTKcGUCi9DzinE
QpWPyK6KR2opk0L+V5VmtR5nBtlEPBSlnmOwQVRlYLKHxXfMK++gSxYlII67
DoTW6wJWp6d/NdjCQoaI4zs76zFVB1stJ+eS8vSge9kJir/FLjkRLnetC8Px
f6ylL9V4e7jGcZ9IX3dVhSqqfYZ/d8wQ36qz7IgItCnp40devGd44VVG5b4g
ppB94Uzg0AFgaTtum4L3894VxWWlV34Ztk6oDi2QcAbbfecKCHZLJPJAa7Z7
Q928ug24tZhUQ+GpKzgc5NRjzlSYHItF5iyVQdTCTo1hcZ0l0+BiSrqDREmH
qVqcWdxMUfTCWLRnuNH56ct5Kf0tKMGJt9IuCTI4UdUeUH2pWUAeZWapT3sB
ZeuLRy9I3OIV+rYEftZh5Xb2wXSXgWPTL3w9hc2s+i5MJX705nkF7FGOEp3x
gK+0ajziixq1ITLsuIV4V7l30TI9nJ+agH9GX8tX3XjIgNl86sT6p0h1z+me
QnnTUUkH2pNfyXcCwKhvitpKDlhdt+bIkRceodP8q6qFwxI2ySuRJSbiMGz9
rbn9EtxCWU6FhR0vPjY0uQQlPfhrXdKaAdBF9lKmvhrptmyIsvecaK7V2Frj
U8TnfBqj/PL9dJDNbcjj8PY9RQSNKrukWKbv+fpcShr/Aari7LQHLE+oJZ66
RRArfyUgWNM5w4J57Fy5UM7rIp5+Nd920gvRx8Kt5ntua8FcsA5KEyjZrB+3
Z9BexSc7iBb7r4FUd9YezF+t+COxtnwhmi7eXQdTr/XLFVyjis5wt9c/kuuh
WFrU6PppCVPsFZCogrD34jtPvrVOLwDEY5foBwqP8veF2njJexeREiSfWHF5
dqX5WBQQC9VQczeOZZEiHMnsyCBunbW2EJkLhmKaaaYV0eWe+wEL+qq4SRWa
0k08OEN0se6AI5HVrI9CHKhirmoA63XC5Ds6joZDXveu7TyBCB2CGNwJqfaK
YBJYpkXLGzBephkjmbSiLbXRrrPT+UlbMO5yYQ0srQfBl1b0Emj6HkF+E1yc
nLwgipu8zDVGFdL2ht041qDoyCI6l2Hdd5RmEw8UI7XjnbqcUtzl7iPhrPN0
nVw+5UBQl04L0kAkCal7v0abr7veOnLApD9ktf3rO8Wo6GfnD7QGltEv3mTY
AHA+kKmK9EDe2DzH2/0e5w+3gGnYr/UsmHsLpI/f3VQ/atZYzXabNRYjr8BH
IeFmRnQNFQb/oSWWlLCS+8DhUozrMeEDeQP2EXWPjfDI/rwWiuBd+lZHfcHb
i1Zl3BMd95NEHLvOWAwDPtfGzSU9xcl+jAiB6TqkEy0XqoXKpNIZxuFBxQAW
RMqUkSv1uiudM1DNpXGo029NHdxw5eK1FFXgKC0Spj/4h8K12cL4dGvhqhsk
FD3IJ5OlvqbAgYHQqzMkIVog6ybmAOWCeA+g3SIpPE/3JfXLcKrt8jWlUBFe
8tv3KevkE5/6V1TunvnDPGWKsx0XtXZF6YYVXBf6X6KbkDgc022tnf34bflK
WZJRN5Tu9F4wet6n6k7ssGmB5fPq1hYh5yNldFtpGkIFt1dCqfVvPZSu/Fj1
A2kcISVz0Xz5y6fIvugbi1owy4F/Zmj7GkPf3FqZ4xwNeQ0kQpMFs3U25K4i
CegS4IAVx11SlxSSF0Y3N+//A/a1Hhr9PIv3exFsEnbdHzdQJz74gUParp6N
+QXjp2Kn9X8o/P1vASWmFoMyd1G5SVEaq3VKooFnWtO+dvTZWZv7//Su6eFa
nYwgxMLb+1u7iAIOXLMT9XK9zZLIQsbUf5okFLke/11tPD2mpmPABB9Ipssg
oSMGUgFxNnsQXCwEn/6eV/GN1YPzkajS/ikqpSWgZh95ht4Pf/uO/8M1AR5g
LMhSBXsvrDe/7SGnf3k1PQE4h8rfxV0s2mmxGuVTt0+KqTVIV2udidHMiJHB
Eh0Xa8gcQSb/HAm/mPGku8Bi83qDOR5DMkKbtxx1f63fzZJuB5eNAXirVEOQ
TX0qZdMvIqt0Ty+Edpd8OdgFkGKH4aZY29WWqDpRp8FII9LHgH4gwVgWHfHl
9AzPIZq1B4b0rZ6JBsgGi2ZY86M82S64TV0uKMw7Wp6XVkN/HLR+4t/ThaK7
gSc/KYcbGJAz06v2blIz0pRoahb36H9mO2qWPCbE7TJcb3rN15asIL4kiyUj
DfbMrYvYT0+BhPorAr7AqksV9mM5317VEi5KPB9Dn2OroGs+8D3yIOxGKRWf
0Mrq91hL3Q5THXECyUv+YFs3Pfw82ieNTnjHY+x2P1MsaP0Aj6WMt520jmif
zbBDIeBLwKwswyMJjDKqCTEJyVr/y3c5KRBw5sE4aLn8Q1o9rf8wv+1hjQTc
nDfSeIbra8KUpxkBSJqOqQHEFC9bOyHgp9jzu1WJxrzkZza2s2jWNHVwiUAE
sfgpXvE7VLOh5EKeNNpRGQ4/yttasM5gFM6BF3LuxlOZIuov/8lUdAm2vSNS
uekTLfyElwlcjmtLEA10akODbriN5pPsLTK75e39bC/5IqRw7e85dAOy1jB5
M6iMMBT2dxUmxtA5aPHVsNESQ2bhXLrbhQYF+53QTsStSgb+WMG70nGkrX7Z
o0p+1eHEf0TePP2b82INXgO+H1aEo6nc64Uchl3AQviiJZDCOx5Op8UO/05p
RoTSke5sx2Dj6NaJduG/mmjLYX2relHnYydJN9WvICBh952hpEVjhZCqvVdU
wTAJ3QqoO7jwaCPZnSRF6pdBpags80kATo4LChSobJ1sNjqw8k2cO9gfpAnV
j8ZUYAzUE9Iv/a77z1RIyccsT+TGO+UHC9sfaLFeEjKZbw5nw3+aOlsGoPmp
xUBgd5xD5pwCA2GEP9OKFFedyF459tbWo3evKTOCgzUbdoJlIdYybphMz/UB
OqEt5Y1A0KDlqjbBwlzlKejxPaXUIR8t+JX+SxBW0TmRE5lzQCnl8LHC32uO
FXk2yrmykd/kAJw2DjAwjBRIzU2D1sclPE/Smcvm5O0S8+Ts3gmxCvYeJQJC
/no0G3D7CN6MS6ocu/PnfrkIXNdYpUtykOklrhPGxOb4elKvqjgSOYvCWfop
uYlAXBePhqqcV7F/m/PkH2gHGcGVc7RRnbJ81ycGNM+2VjjKeB35numr5iJi
WhamwGYBdRl2bd/KV6WIKe82FTbUrkXmDm+OAPVc2fqEA/igCwdgusuHDaUN
JtcOY7Otc32e/+4ObWygo2g06u98DygrXAKxZ+xa3fX1cdBULHEYqnVoYJP8
bAEdDEG4paUs2mOdjtUtyzVjYEWM5g8ne0enmB7dNLg2evLeD9NSqj18rqqf
wzDluc0pZhrz7Ty646k7GkyoiQkrAEeDneDpg3LypXBIf4X1mCnOsjPTC8YB
+codGDYrAGYxB8Y9MVGzjWQdjFJasW7cV2Fc3sz3c2IHBFjuuC4EB0qe8xCb
vCiZDK13KoapZgZ4XIs4IxwO24ICkTiafdMRwgzlUzWUzlE4yFaDm8OXxPHw
oG3b2CHy6AkHOUsWY9liZ8hfAoMVyAS8PH/NrC/9+JzwwNmsdtISRrIX/wa8
iXspzoALFsSgOww1pQy1ScS6IZFu6lhSwES/ORD3tlhanxt+vZSxN9Zx7Do4
UdkeAX/KQ2kO3rO2MgTxPKhjo7EVRPrrSuBXbyt7Q9NKqjtR8CLSfSFiFEcR
wSPMEp/EkiVf2lREuIlIwB+RbLe6Gw6BvcOapga6MVazEMADq/zbx/L2aNYw
57CH

`pragma protect end_protected
