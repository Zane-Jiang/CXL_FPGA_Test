// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GYjtU6qDyyxgL6GBZ2qQsPgL/GTC+1Eg83UBQ9PDVnbBkYN1Hp0A3kq6G9Lt
CNKblgpC+rQd1rtNx9tSO4KM2Hf3C8QNo5HRkVsaQlMuWqcUNiujFt3ypdyp
4WigyUypTX47c4SD/igO9Rdu3SGn73T6acp32gDoDeLIOYckL+DKkYtb4cFg
TAVo+GEcrbF2z5cdHECR17KDKceLYABzMH73rkqVAyMIMk6hlq6cwFFj2LEQ
XD/+UyOlOCtEM/rI4s8Feyp12N3klVv9EC1lFOLMLiArDHyGaKUDTfUfCi9d
txkRmZ/F6YgxSNbYym0v0KlBuum+0bQajF2HS+KrJw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AVho1EOqdMYroxU96g+fHVjqfvd1XMuWjvTiHC/ZS+Ndvb9QGhdY2/2oGh5Z
19ZJU7EhTVxFpfy2+SnPHK1T8e1i3Q9dUky/mqOEX9dlQJnYq2Ji8vSiuPhA
odwwCfSIAuBPc7Z0JsSJvpFMOHNr95pa37EQr8Piij2NGg9AFAHpTNJBxjh0
86rktClX0fyrwTVNGdmvPw1yjHkAH/Jzx/f1UyjwstQMZ3nZTImt0BzMvtHR
EiS7MUD2YvYYglXoKi5wZy84uJiwze3t06vshkSwa1oOhRcJCYp+5wVgkHOW
4zYwtdNsU7jjcnPBCFCcRpYpn3d5Lh2BdBnnfuVgIA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZVp76w348sNqZzST54qzIX43A279LX1PWR2q5bFGKFK6Q8r3LOgYh7U4ZEx9
ezKfC2TeQz92JxtKL4tJZrt4wEN475aT1hSFUbwJwg5uiJfZ6FOgK0/tl4dm
RlFqmlfBQYmCx+EsB0LQ3pyMp+jXh0ncj28vBjl3rYHXsUMGBq4Ht3yUuuAQ
4cdgWf7tXpvGZBI0Hrr37RIj2Tm0+qJCd9us8fgM6Jrv5jwGs6v/DjycOwEX
FqFhR7wj8Jz+BLfEDPFCjwfAs4UUO1/6NIKQ02Ef5SWdaJBedkmtyj5qb3rl
3220fhe+9eryFd7ZfjXNP1utJwziMIbYGrcxksJ8Qw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KZ3tWsBaOrwcxG7MrISQkS6jnhnRhH0RyMMH11iDIW4NcvI2TNz7JQRWe/rV
1oDnib48RObGX41YABuNt1FtwGLvugCVsI4w4phZVhNlMk3gz/bpoyOdvUAC
rHZj97VbpVYh9wKl2shOeSGxt86rVu0GmkeyIUqtPHx+ZNMpkMo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oTmZe7pZsoKJslxKt+Jap0XSLWN4OlqO5EfZY2smYuZcwWJaYKlyx/dW1r+G
v1A65t6PsT0IKTU/q7pxFAHozYRlObs21v3TIp1sQqiHxoHfYr5t0usIH7HF
Cb+UBKEbJfQEXJILmctaWeZZhGPh8Ptv8hqd8WpMyv2t9CFcrVj+1kNo2fk4
N0qQG27jYaN8gB7DC23B0namaF92Tk71DdYWvuqs4DPCjCU1K6VRuZ2DVHBn
D0zdHwCnxfqoq8ySHmgiZkHgJ+rwnV2YRb/GpdbzwyO6xApflIKC/xb8qXDa
3YIXbvFsmYkmYxmtxDbllatzxWRF4PaAu3eOakV7h4PJv7epEu1UGau2/LBX
wjXdWzHt01MJBLwpiNsYWeuormn2kedZuT3TuP7nkMqnUDbf1Wuy/DCAjlak
mNLH+pEe6yg1ldQePSdhQleK4l8naDfBZYvZMIBZ/aZDfKaZARcwMWMa5pve
Roe594igJlHyhtYy2hHjF+j+ZPUUE4Q7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
u2JttTIEk4NP0Y+Faw1ZBL71w6dXRuMClXlqOnhRTWecO/HQDnLdGluUJHoL
hdVmKC6Wn+cUqkFLdviTJHery05yL/M00nOlrQ2dN6YpgmnmnDn7k4WyE640
94g1NnjHJQM5yEEZfmbFbKWPDCHclBFzOMzhVSIfRj36E44QLq4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n/SqAhxoG6cs93EVUittM9jYPI1gt4h6UVE0PG88gHEMVZpQa0mBwoh+f6Yg
4JA6zuEMEe8piRHhNNhzoIslTZlyauT6uYOlWffIFwdgGO2ILKhKYYpbD/Es
+WZ42OQIyC4CvtwSfwHLsh+YLJcI0lnWppmGj77KGHBscM9t+FU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 71360)
`pragma protect data_block
gAAMYdzyCCLVLBbzT4ehtAq2rivt66kjDGeZq4Tz4Ab/p7oS7Xd8GRHn4tmp
BrKbgpPspaGCz0iOwGV21KQZeuWWfVdJfHYD3+Ov4YGGG/Tb0cy6d3JwavGP
a7Qrc+YYr8hlzuAb7KAIPGAiSfIowzp8Js80SGtQysxiIyXo7ND8O4gZ9M8Z
FqeOB3qrXYRszClhE1aFJpRugtmAHTs68a+6rtbvWQ+twzx2j3DEcx/vFsXO
93Oh+RQMAQu7fdI84smju56DdX3+iTWZIzfJEmJMovhHQML1V8qSV7PDbBrg
XOvMcgYVku3e4/dn8RDU/9KSo2iHW92yQ186FjxxIx2hvqb32NY186Pw1trf
ipnh9ycemHiXSyYM5n7tgweNsmsmjC6L+/tLXZvONDITBitvTTuzWwSKa5Wp
a1dNX+xITIIkjgtJJxDOxzilKr6sS48Q3T5MLgcRxWEfKcCnQ+wfLw38KTa2
EZZby9E+hpL9YG6xEcI+ylXXdznHamLEWiovVVXTSwVh8Orw+fz40dSbt8P2
Ce6SdKtRPIXMSAH6CdeIa4wVdIDaIqU1wo7T9zTn2nwDkAp3IhaegAeZ7IlD
dejIG5mYsYjIPDlqSRJ+BlWu78WL/615g2ZAfNFodaGC07xbFsl3ipXn7C3u
0TlFn6YXKukZ7IbXZFMPcP/Gq8cDSrOzRelbqw7dRI1M5dIjnT6MGG+hl4Nu
igweHnYrv2eS6cqrw1Vi5IpDmjq+F1CBgpqyOb8egN8mTKMbr6Vd1cZjZCII
lN+rVIiedx9RRQulH66EB4Bd5K4d1ubxg9tHrhLlP7wnJEaIBayrphFexK/8
FtLBPFT/qeGXE5cZj90gUXTtU+lnCAl9qLW1m9lEJWBA1uZokFHK8ZkWUUZP
N9MXkraYY9PEllAEpF8S43AJKbeqS2CSPWkCuUsI42puKbZyriQHtKqwpLid
HmYeb41AmzS9yq8mIgFjSlv7obqTSYovbQY4BBIiJQFJCd50Gw9IudVGPPyT
IlOqK+N7y6F8GzoTtnz2Bym1/qMXGmyZkQuMiCGuSKXPdfJoz2/eg0vOGCDw
SxKNyNrdXyH0CkNSKh5klo4Kj4MctQPQJ+b/gvidj0e/OvE9EQs/xZWwifgJ
tUO3tYNqpucNnueeNDZbdQc3fkdOqdpcCjLvFCjOzA9b06KDOrkCorIE+HlJ
aqhAZKPUoli4koRdz0m8UEHY5HnFwDKL75kJPTtwFzXuH+SOHopgRWHhu+AX
Zd0bQ4twNpDpZW1+z6LUIzB1CLPHe8KVsoHGv8Far48wTSQZ2SoAVK13bucN
ihboHmqz5xzUPJBkYL+HnVwKbwDq7uGCTb1QqjhLuJIiLZJB7lGa+0Jv7LUl
d5vAvpzRrPSxubWHQh3hByQfEPE3eGS8wbG2AL74NKt4QGjAYf7dWeTp4p0W
IG84T9B+UQU+twXrcUqgIR+noDT07ARD1Emxnq3nsDk5pG70ZIVCuGFOFnb5
8xzgf6IWmnWL4vik4+bC/v5ACeDqzG2yFiVEA4KZRnJO/DjAQshJRIbvGNFN
H2VtJJs2EXWVOC3QBKGzzhbCmdq6toHN42MZcvtos4SU9ZTdVlUsY+pSKVXj
PCuJxpX+mh8E5V+V5UdJmYR66nZ96Puhdq+scPY815ozA67dooZJyinOhgkS
fGtPqm42yK2yhz9AR1TNVD5yQUN+ba04cx89O+YeRHcFroiigVLd6iSs4+Ey
p1KIFGaGc4tfa/JFLxRpdU43vfA5IUDugMacG5IcPul4HCxmN/o05amnijhO
ZGqQ9BhIQR2JsYHpkglPvPms2G9RP4rNNQRxEdw+9tKaLmsyEAgeu+MEDBGy
EgXR9fJk9sAmTeIZ6pZyIT1bxP9UYvhkpShRp3yrsRi1+2myV1h8EAsqTIkr
fkPjPGlNhgnTO+i/aMD0VeSpOGeZ6tC9Vr0pEMsnqrcT5iaOxYq3xmJQM0dk
1TsfY/zrG26PqaJiATGl2THVMdmzJ4seFkSzK/fblk88eSuTKBF10pIxr3lZ
b/S41si2WEcrNMI04zNcUCAbt8HV3XphJA+rj0IXgU5IrWwvzpPt1I9B+dzv
OZlN50bolhGxY6ABkUaV3tFn1G/Oc09Mtt8CsCpHF2Y36lpS0LTsy1+LP+cR
fqUNtBsHQdzDp85TL+9BMh0EBpLDJIkixyUfwFUd3ztywuGCmxMWJT58bJN8
bXxsk4UTpJqJI/jA7YYhBrPgRH54idCSmZwoJERoYLf75MB19G+b2zZMfiDD
9Xm0wOmYCiiBlGX3NTg7o514tKQ5QZCGqNLdT+QQLPnxbhpyxLqqySUQe5wY
DeaLYvZLf6oxwLby1W0konW961IZBiqmKMjuQwdnONk68uefH5PgenzkY+im
wu4tkiCYKdsUN8OVsYFNwP58PEAdEKToO/D16tWRa4cUtVD37LhaZjeCO/C7
Cbj614h6q3Hk+u8lOMsrtmzIoB7/b3NRq0vFh9jIGgtUTx7wmihdywcjooQN
BAA08KmXOOGldDZBVhHon68mRH5rQvgZsfTTvyjUpul3g77EmuYIGvqimzlD
/m3gdEJUlA88Tq/oYukk68hgnWb6E7QFKT5Qk2/DhE0J8NQCx9luU0Rn8fkU
efQrY1sZGGLhETyHNFpcE30BXCqFzMJIWAU3qtQj6Hr4M3Yl/bwFc4q3w6nO
cSBb41A9ALd/xFj+3VYYMqFbbRTTmp4FGtyC4oXU5EMXeV/A2o5n4KA8Eytb
n+yR/DVeQDFM6av1Wl+ASNw7ZbIN7qc2291xwXcvvOGS+Yjo6cdQAix8jeaH
CLJsFJVWNBgHVKwNCT5rWDPIoFBLMKLvrKz3M1qCsK7a+S/XqMN0Hg6IONK+
ire4clVXRtYib8zGzN1sSAuUyUUxXH+M9PPGyNTuKkih1G7P/RVbKnS4ah9d
lI3KFyEjQ7dUWXN+Es7Im63cy/gNOXeP/691cKmLqXbe7vNFOsOZusACG9Ph
jNZPAenvdX0PapkJQIj+eYOUcbChIXS7dmHcXiY3fyMzXvUyFarX9YHv2S/l
dVnZEiIa/hyzeQbkvuxFMvfc7gMxBhaTu3GF416TvKOzV3gfGg2VgWe60PSk
Nz5+hQBjhgHQS9GuZxE6p8Sr6Xm/8DTKoX72gsuTLmcnWhbdtU3rZ229YRbf
ZBZ7Bkk5PqENJ2j4L2QZ8mXSmN1ahxQUBtyX+KQ8zFch3DnIdsv/YvmPuKXn
lFtfIQtxCivnZiHWPxERaon1Xo/iaxDOIkSOFwzJdhua783jEKyqgwl23KcF
8GXSqqdBtctb9+ZL1BXl2mP7Zl3u0Tvkz1FJ0Fa43SpvSZXtr7pqPdBkZQpr
kPvJKgJYgCf4QemTFVjaVlQ0HHRDFmN1sT645vRYYpPKwhZIUCO7nNQ6NmfX
ftb3jGNVwFE5/35QSw/iWuyXFe0sRqXAHBbA1+jyUli2HeaBXe5j/PTJYG+9
b+KI3ZHROEAUv5DfOtzsWh9mw9GT/ATHALRW9yDyULPMUBcAkmBN6TI+0MKR
GRnZCKDxVwIgCsZv2dmmNDVI8PB9RCsylALlipBVKGTizEHl/5kc7Q1/H+AA
bXPkHHM8ev3cgHmWrdzGD+ifk3JSc0xuzgNVMZYjNp8YKQQZZGegaZwSwyqk
Iv2CFM/Hodzb221KEMrFI3GUzFztmyoG3P3IsJLbhluXMP3dbLoH7sqk09UH
CDVf/FNMh943kRSJMRdtGxZq4FxKggYMmd1Mb+sUxzdLXLeVUyaEQbWDpnMW
QF/+fsWkm/EuAI/1QOGNaVBrN4tvrXkipKIlDDtHCgNtMiUU5xKy+e7oG/3h
76LAHpzBA8cZhkgO6TLKyFP0DJQMdfcPdjsrcag9bZN0U6GMkWHil4iJAVL9
sB8qiSvdXRGB9S34zEyLloODxjqKrJwZL8PVOFP4JVN14ZjnZLTARFge16bv
bLP81tmYdf0rKkUhMDXqOgqLPvaeXrF8e9kf9cebxRCStasYo8QxO+aQ92aO
QZzA3GuVqbyLHDb7HUV0P9gMocbOCnPQmfHl4J/LR9DHxK8e2pI5TAUyl3YY
kb/imyY7M7KDfu1Arb85YgsXLB5nVtqproJ2NI0LuDxwrP21GcCUxGf0dkPE
dN4Z/Da4vHaeMDqbef1XyThO9hcRlpKk1dtXCeR+KTCaWsFf2PMibi1dM7zR
e/gZ99FrCZ5qZwSBDNUt2Ldwaut1a6EsaJ6ezvCLsQZC9wrpHPFey0Qw1JJe
jug+T3u7JwSV3VhedauBxcB5TnAghryicfT64VxoEdOLWQc47JhkkOgdwQkE
xKx2UrTcC9su5t0jGQxVBTI4cigdgufjAVkV1pUMVMu354mg4/qgGepIH81m
tikg5rtfS4q09e0tuOyRSUKrDOaF+HTVdAQVDwajLEJO9L1M/F0JMqu0zkuL
xpuI4sA4jTEhdL2meDquHS3wsHp+mSnepimjxhDjaCIuCYR0GJcF9fgTdUQZ
nsHPtauuo/tE7I2OxmJh3m+BCrLGd8JpvlA7bDRnpY1vi6FcH1z3Glq6h6Qg
p5iZpq+btcWxZR/IkiokwqDXmzNi0mZBQzybFVRYWFue3Av+ldnldCjKxscG
jrpdyW/hnlBENA5TIWFUoh1m6x9gPUpA9x0tKgj6aE/J/bvtUIBs4VWvlXfq
Wtr/QnX3b0Df+julPlyYk/cfK/mmPsk1/kEr8IQGQxfV/Zhl9jhS/axea6A4
4xYFAoB8SxGOrLKHpRJZOSBKYkJ9uElq/kh7ReFcrgrNZewzksI7KJOFh/NS
HvwVMXnv+CtFniKcxqwPshQQnKF4WCUfr4kwgV5Gr6QDtGyK+8yaZFNDCKwv
awxM6JMSqsc0RRU00RPjuAEfc+WpAiRCXkpj12+NitId9lpMDcNGsRKe0jV7
erxZGIsuGqk7+OrLKKyXx2ZRIrcu+4MOn7Ig/2eYF75OBRwaO9tFc6h/54iB
rZhvGTiNvLSD+LxtsaaUZKItK6KfT1ASP3ENvJQqkFQusmzUsvJuheZd9o01
OZLJkrdD/9MTZYkd8wFEe4t6jsYari7q3P/NHP1uUcH2988sI+ec58KA5n5/
VVhGytLS+O57V/UZAIGT6dJ834F5UMKaoWRLO9rpqVBaBBnl6q6HenJLorG4
GxMnfajmIrIUxmWIOqFnacELxcBdaiozD39wYGWSJPFPCTjMJpeTA/qJXvoJ
x767AcqZxtDnWATQZyCP1FT6ngQ4OSvAlnOZJvo2WMEBH/LRZzN3gimm9pJW
RWZEOE/1y7oThSmvM16CU2RKB2bsJe/XQGpi0dU52weQ3lcVjBBFtmseVSgQ
/yqbVsC06KeNffpBocPnOfsKzDjT+iW5ONnmE7oiX833VBaYdEkL4uQdLD9+
ArO5DvTzeZLYzcSyi9764l1dwwHd+vPRjdTvg6MJyKxfxbWPj25NKv6JEa7B
A2P6+mVkbRv2pr0uKtS2b7x1uXIwwaNoi+OBNtLgNdC1zNRr98KKTyEyc3Aj
gPWWqXweGhFMqQX0O2lfnL1QHP8XJWUlYZWC2CaKW2HE2hh0S4nFXRes0gTC
qkbhqEAxPCd/Y0c3q/PXiQUgc6HbHqzucpA+njue7r6ZzVikchhnQPNCRISq
ia824HW2fVXB/6UW9uA3Y/aktsnDtGrhV4VKnhH9QRGa2rLhjHioeDQ7lf5h
Xj6OQ/jQtHhFIH4Njzb98fyVEzQUNapQHDfsDZJ8tyuutzN0NwibT3EnOEAV
t/rjT9QGtrPXbZJfaSStaoyLUaNE1X2qw960ljyhoo7odNAxE1mo9SDnlIUJ
TVWC1RUDCXNbY83oCIIYAY8g++OvKx7Wr/Ga6VNzN2+3tFJEmpWkiyazinep
7eayqa2Kxkym/um9Ptz8feOA3v72lD0GYxIetFJk//1lzFcgNO73QjQaRNEc
7tjo6mIqtbtJx9qKftGEWqSpvRVEUPLyB9AczBOb+9mZeGD816pOw3pKvDcp
rMG5z9nJmN14d7VHK2PlCQEqbOSKIFvdWjXBVa5RAq+ekAobEYpOh6nDgwEe
+7SfzLfQWUrb4DsuqnweYdrsYHLi7afvvuBi3dtSRY5S0Jvi4PUyhOfJQkTg
DMUEPkkWjN7XY5VU7J7BMY9hPLeei6BYfgTt2LENN1itPxfHEscGSG9m/6wN
rzQfGiWSLV4EuZrwkRcgvA688ra7mdqVSK5ggRQ3seGuD8PUL+HEhfKEHUBj
xnbCvg3gs+8LvVH9tXkw0iBb6bNU57j+xxGbXd2bczSLowTwnCeUNEhCoYih
R3iExTNVypE27fW6iyCQwrUgC8Vo2X1cytUa9ak33GEMO3p64npmmY7u5pmT
QmbgB5m7RnS2u118Q86jdtFxrWcQr+lpC8BIjj+C6TkguykVcoUWbbH1NzlH
0cyAkYMrGvFrOuSN68hHE/NxK1x3dbIrAz8ysWJOiw/37TKHYv4yGCliTim9
F2ZoNXkbU4/Nz8qRjysQMvHmMq9LLVJ8qJaesDY8MtYscXwPwNoSIcf5ucvs
rwLWS9ihX1stLemh9ORzl/Ol2kpbzbh30j2ZQMadlSlFcGIVGJptBwvHkcRO
eSCpiqdwMZGWnti6Wvb5KMfJnIuW/8lHAGe1JzASC1AXxsPcW8mcOyuHhkUO
k21bxPspu5xes2EPjPZFUeDI97HGWNUWAphOpZaPFVi14lStvyUxE6F5U7th
Y0wi2KQUZkgfZLNPNk3th+LN0dy4VM99kZcugTFJ2ZVI0NPh6l9LM5mnn6IH
o10+6hoRO/VLWu3P/iEvfl59W38Jb3K/Cc1xUe+xh85sViHS+V8dmPJFx6qI
gm/vnCMwq7RaoC01wPQQLPpnUdlK5AbRyVnq4fQEVS6s3JqGGQQ3tIeSfy1B
s9BBatTUBVhr414WdoP3uWe+xBHNV43ZYvGdub49hcewHUTZB23dF85xWZIL
ahcUY8oyNOuGYTIY5pqrxZE9JtZU/ROQe2sNX58dL9BACuy8uPz0cnM3F4Jq
l3nOmgFBLBSAr4+yaVBqvKLenbzk4gyDhCcQRU5xgwcGyXi2W0VUmYicHmec
J5E9ghTv6K1iPrKMnuFRe4BWXrxW7wMJvFF7MI4l7PsdgKog9/X5DJdUN2/T
K4JcdepBT4yPRpGpOQ8Gl8lbckmFQxgtuaFpIkmL/ABl4cfaLCvqw9YXBFkF
xGbHIQEpBZgmFE0HObVCHj9OcRgYw8ugG+8jSU+dum35KR8RQM5C3taSh1bD
0snAG7BHxjL0iM5KO453WuEuY3wR8oo6HJiWn9k/PeTUDki3A/JDhJE8lXC3
0hxEdgtBI44yiqH/cXmOzZ3qnCMtl774CN6JkL3qBPCcweBSgATOB0p2q9mD
PEsYd3USuO07VAE+Ku6y/+CKssrbRCse5wxPyZIa6KrjtLiyCy+ZvrTfSoCs
LmzZethzI64/lfFcuDQYQubjP5+wXFePxfn4LPUj58Zx5E55v2Fpbfci3V0V
9FO/gz7gDh2VAt0LWtq0e3j18KjlVnJTwFsWOoPlntGLbEP4rux9ja58ubwG
0SMCvHupg/sKD+V5PwxBJlYD8rNJl1pWVLdijOFBzHmqGefXMKF78bLOPYwU
Go04BKp+/HFildGPX2w8c1hkB/KKfHY8IUQe/FQN4gvj/VtYo5i3AMEnHJ9d
IA8IqXqzpD/CK1Fx/TipjNxQNhbzmhnZgpX+vrn91ADDW9MEvOGyFkOey4ku
xf8vPzaweklgOzs4E5nY+6EzVbZKRFF5oa51KYFVHKNT+V7O4jQC0ZIQszoe
n1ZQ+pAyZwnsvSL25AIWQFmQHtqwHxTXT1KwjV9NqC5gx+tiAQzo6M7UmRkd
5oIFsM2+20NuhHoOAG4hQIFV16Ct77Ki5HyOEKyCHE+zNS2VY4FyUemM9rCl
JQebfB0vQv/YQ/vU9/eIwVlu/12SlXBUNlqahVAW7Pw9ZUF2CRww3YX0kLud
v518AokKJgtrIwtmtt2G12Ma+8C64nrk5ipDheJgZehFLOrA2JSaPA9lrtDa
6F95V79WKiSkSVJfYFVPJ6oPOP2B66G1gj003QJt2i/95PacYXP10Znrnsvr
OTW4rl7P4H9+UdcPNVY/9N56bP+G7mH/mEvh3a6f62BSKFS+MKdIlX6oS1O1
rlqrv4zlQFLkAbgstinoJ0Zv1SQi0OunlVwi3Aj/+d3abnwKUjpOYHHyDOuB
5qdeaDgV9bgywYQlz0Oor2FCd1giMZ0jaqjYcfeKmRApa97ho/ODUN4nS+nW
i/C99z7V/9lKxz34IF3EE7/c8t4Q5cs5lByDpdROhklZEe7ep/pbOweKkT2R
NJhCokSbXdwe2pQZd0/JYyP4zAliOhN+EV6l+tZV7wwhZpG6o+vF2XPfQJpC
XduyzdeCVrCu8PpeBabAHHSVFdbnSUnydOICf4eCMGoT95k5rlMKVeXT2iBP
XySMv0kHFHntTxQMvBlecfUn3cO+a0odFkVMWr/Ps+x5o69qF1axwSZXW4jx
Zmcozad9rAip1iVNTmj8aL+WY+It1KuCAnc4IR3jFkejap19MbnGYGviR95G
9WPWjCndBmwaCQ0fJUtC+amH3w7IToDSFhmA6wlplAKhVCNkf+aoMlIJO5N9
AODHevrVMhpIxgnDCyZWzq+88l2D7lRT3c2eB16jau2cQBg5A9OmEzgSWmqB
IX5oFVqxnN/GhktoOoT/65q+EXhvotEQp+iu61Hd92WylgOD24CX8dMgpXbI
ux3WDmr/y0PU6BDUdrt/fv+fbIRa8jtzEhaCqEA1027HfPdn3b6P0uJmnIIB
E6Ukw7Nq/qAvrf9V5fEHD65XdweJj0AyWIXn7m2rStozdwOJl0FY1oRygH+E
l5XthFdK9ObC1v3NUOjOrLAuiNZtoNhBSgepjxgPtgNokoznacBLh0b04Jte
GIoJwM2e85W2xn3XGv+PVmB9i5Zg3tvAzfQznU9vVVB6QhYpTDd8UdAX9eov
1I4KtSqFyijt+1guQcOLskuLPOQl1CQGXYRVwRZdQO/SsYVH4FKNGRqfuoDg
3sinOsYcc7vXTB1c6vvj7JZ5jqkHpABaXxMsZk9knyqZcETcXhuyFlIk+JW/
U9RivaOigOom2K3sy5i9WZZEzODeXur/jGm+pSmGuRMGP8tDse+/R8NpLcEr
+WXlDZtdAYahQKLBfmu3n3PEyfc1vkTpSYDNw8zVKed3ssFY1gZVI/bxXRFV
OgwZtzPv4nNhGeaGHev2BLYhhUsq3/6B8S5Z4vKUTn0Tc1GMXh6i1SyMnU/R
kwGicIDi3cpYlfCOxt/On02O/bmxI6KS9Z4HVPJZ1BqObLG/zKBvM2u+NBHy
k0azLmzsW6p3KhnNUMyC/4lHUR0azHozx6Nta6woTv7GN4ungU3xnsn9JQjt
aipPuD8CeNKVOELOnkKZC0+tbsZSi+m+zWobqS2QOZl5ZauIlSKW78pFJkLz
BEsULoq729ADkif0wusl2Y5bOrqubZh/hfLRTRuHVuMF7+NzSwREYBk/dIwQ
mgwF78qlDsLRLz9r/2WI3x+pekn0bDYPFg5aknpmpsE83nNe1fwXlhbrbGvc
0NIHL86eElvndqhsNWO+Q5rk8ewC4m2ib+3S6tQBYNlB62x4KzeZufY09V4V
aJycRutmi2PbXHF3Ad3IU7ij4fbo9mwOZCXFMFkJPhxMClpwG0zxwEdoyjuP
cAdnEzFr1cxB09XzYNu6jBZ8c0R4L6kGO4hu3zD5+TJGuqFHuws2+Oscwikc
1MyNjKIgNfglZe36tSJeGgw+T0i1VQWMsUcX5+AlC5Z6lMmaGydIBADBz/pA
wDf7M0sUy2ZwQZt7fmgZ353pkzMAZ8nKP6vy0/7c/ucEab9t4tiUF/UFLIiq
EhFhgIrKmYlKjTQT7zSH9Z6+yi30thrFkFa5ICH6BcexwvZr0bISwGsvCZpr
P5rl5FORpMLTUG6Js/1XpM2VM6K730s3LCMBvR9Hy9OwxUrhGsjb3j8AxAaS
weH8et0rgUqEYBn6OsioO6Hut2ViMGAR3zYHMDCMvVTQoJHmKeTzkrnv2GAs
A0p0BK7ip0rty7Z481CAtfafxlmu/rekMrpMqdBKVsNNpahRtnlaEqmZS5KE
Sho3Jcn6A30gwK2swQFUE3mVSDy87r1+ijPbBKH/o9gr8ZakcVvSxkdDtm75
Wff951muaBi54gPRa8ui31GlLCSQmjMWeuQHIJmKUM6otSI5sycJ8tgMr5HT
l/yAtImobFluLjwPTjIhdiF2N51TaXhOA9TAjc9E4LUvxnqCSAtak+hAupr2
n5/sAilpyMceS0e6JsAulQN83Qs+6OlICYY1eOI/PbClZMW/4aQHK8UH8kKK
BXBSwNDfC9vTtPg0aIymWD5v+HlBbyMgNIcTxOmcZ2qfSEnsprOkK04z6k02
wheM+kcuu7QDjyNRUQN6ZD5PHJAbGL7rfnNYqWGM4Jgt34xylP0becg4ZeMc
YMddij3yED71totDo+KOuXh4c+V0ykoSA9rYA4GO+1+q3PVjFh6vqRXmh2yu
WPI2yqpq8vb9eVZJLIaoUuXntiPHCdgCkWjmgE3729agwt1Xkag7JdCLgtim
xEBYbXGsN9ze3nhZy1Ni/pW2JkihVHQJT7tN94aTgsVoAULrY/4KryZlRxDa
gdGeOtXA3hoywKjqabCdNKM9XJYDbmnC4o+58YWDqQAnIYAqBqsc1/S0EDCX
Dy8IkL9oRM7BziE+oAgbyiMMnywe6AWeAFOKrdc/mEovhUnibKS5cz12CNGE
Gr0G1LdgU3PG+r7hDgICqVcYGZ/zGk5PwRzk70Cs2qSzDQKU0VoUIevqQ5rp
Fcz9EhTA+X7gmGROYBl5wDEOwuXuHer4KZcE31oyD9j6MRkbaoSzKcj1w/j0
ohbeVtmvjbc+N9Br02Ab964UWxuwrfuqbnrHgXXqLsBEac3VOqufyFMHoNIl
Lr33KwT2uVAvXHe7Q3/N3Pw0v/6Ip61m9An+13yeaaAsVm2t8s2FH52pD47w
LmnF7I/5opLHiDRWlzCnX57DpBX/YjnxBDnv+HZ5kQM/qL0b/W/sclar2xYx
7FVLP8wcKS74ur+UfHizz2MeSySyRlcmT8EwpttSYUzQKQLmae7bdVZNrYys
yQBW9WUhDiXXca/FrhdPaMf1dbwrVeb2G99A3QHOhsxoPAXJG7oBNpmpJoKb
yEUPApAt4so3ri5ngjM6qdfy7TCUdGqecc33ymrOSJKidTIfK0b9LphXHzcL
CF1Dy86umJR9nFhreZVjFwmTA6258jL+Y90NGYQT5PglZ/wssLUR0R9ggCoP
MwGUphrNMr0aBIbC7WsvlmkynH8W5SzvHrkUxr9LoJqUNBFBZLFM7Cl0ZQ7w
JEICRI70FeUSblj/RvE37IEN2jyWEBifUWIilNgZS2I8v15PrEuXgImlR2dl
U1nDrT9Lwu4rdoeLw2m77V7odyVDK7bqPvMriBIMeTQ+S1wUwSTkUV+PFWoq
vPc0bYDlh2K0I9Nkw1g7MyZHoqPghsRTkf1lhers2cdzmZOLIf8yxNl0q3/Y
rbuv6OEhNoSQWLXqjI9s0/X6zrIvahpFd5RSC8Xe9goi++ucKFYZbB9yI/z2
UVI5fdnpwcs3buBMNx/a14zOHcqPw4zjMmvmqW+VUz+NQYhyM4PurGWAMe9M
89wGwHUO1sgAxRpRA8Mth3nQFaJ35XJ3c7TayrU4mFx11whZUKEpCQiHLrQS
jQpl4UOlUosH7Em7i8rX/Kw5yqDMZjiQfHvYN3HyAdLn0cIJmn96B1YRGbMh
DqHyCJn3fhld2hvJ/xzRww2LDEPKltKlADb6QzwlfPmmVMeD3ArDzWYU7Xhj
7DH8DbRtMiuftNOs7iiDYreoOv4EnBE44GbTwLqHOAtzYQW4ts8s2sXV0vFR
t+oHXjD0LFAkltiVWEVPNs9GBWjwG9SqGLtwU+AoRaRCPlAF26srG+K+qhvJ
3iSEE1/X2kLvM2p7lpj5ysydl+JakvmmpC+iN4Zq4+z7daPxBcAKg2q1Z8gb
OxMoUqtp5a6lE7ztNTAqr7lf/5ibbu/p3w1u5aGcdtUDeCb94aeZdjtLM6ZW
8/2aM8ZuM/4CfNkVdTSxKj6BL7WTN42gLCjDQgQEkPaMov+YwTUkidqPzviO
xZrXd4X6qL6vvtKf4hdU3h5GBFJ9i3Uys7pQfDpCx9mleddYvghYZ7PJCAzC
X5t5lL1MdyzfXuuayy7/qWZFGJAOoOkBNTySjK37rRfEqEBo6v+OmvZLLjpq
UKrHXpsmrxMs5KOlma95fxJEVT9pDBnmWQUpXCQJovz0sqmYKW6e2GcaEiQw
jRGf5rhp4hNRxigA5Ou8xXoVKYVKe4SyJ0s4picKnWaay6r8IDoqCUgXx/EE
0WtdI7ySyul7Cg92I4FI7flw5eVDU51x10h6SMsgp4Yu4wajzReePFoarmLo
+bHZId9KD+o/6TlaV0RrpTZqlrNsK2Bm+Z6Vulg85Ja43jL/zl958WFcCaX8
Fo04PwFD7Zde8CSXT2RLg8XeY37ki8RLkgGdAet4QwDszvYkHElOHOn63XMZ
d+XcyUh41AiOGkoJ/itdlBjhw0ef0rlurRHQMlVtmqBLeRxW/c95sS1ORAFD
Xh+lRelmmJjoskY2l0wOS7EP4JEFsJh567rPB6jEPamfWe0veNJ55Rrw9eGs
FnvtbTyXpB73U5xmY9ggMIoHq7WpJUJdIiFnlW9UWBJ8BTqSwpddQ/Rb/7M6
9Yn4xI/lBmiQs/uxfr1kgFS4X75ASECzVYiwhWMzz4dO7vAv9gXQCZJafIsf
CpsIPTXts4m8M2xX1rfix3DhSI1C4ZpF3Z30+Z69JtVWqTH5v0k1c+Nc0Zmj
iYYTFxB1rDeEdRHe3+jD06VNRvd//3d6msTnwZVLgrnMCRZvtBhwEm+V0j1P
k0anMG5ef6/WP4082m85pg3SAvNRPjMQjBbFonoJagHJQ0F860Bc3az99PDm
0x29Ik2EgaFymVraZ861kuuwHSP48Fp7JzzOUHODGpQavrSBo5Jc64n1MQdl
H7M604/l2fY7hrbybNPmH7LOUTlj4JrBAj16cjvWytK4cLJ5EB5mmmT2FuwN
A5hqwp+LWk4z/124q7Pih2aAsM92IpGlEfM59Kl+0G6Vfy/ckyV6ygCr8+sV
P8/MnIwZN88XcI43ib+2IrXr+4mMGovl63epQKhXCIQWmYxyH3blgMOx0hTY
Ja4p1KscQ0UNlyoRCMxwVK2havp+huwIqPyjG9nCt8Qd5Xr7zprkB8CygKv7
eNwRSvTlXEscbQzcqpnbN9VBAezSXrTEl3G5BZZ/TN7PWPu6F0YklJS+53n9
Tadi5zJxFcWSiV+7KqTT0AEGUnqIbpQoZqd0BpCyWkvPVcNaHo14lTYB5pC/
qIo0iDn8EYpYbRR0nC6uGJSm1DXVjf8ydqraVBwUmqXBAWPROnrCcETGEMTD
6MJz0IqtWEq3R78b+6bw5R1U4tMpOAeUugRm9lFiO3D3jVIczhx8ny9xvNbZ
4r/f99958efs+9xnrf5+1QkjzGBm+ogc/mxPIDiW/3+qTgxby+Cv0v7bjCwu
knw8EA7qVXuV4Jy5dpuX43IVerL36jCvrFpb0XsIANHJI9CGYffkfm9gTLtY
9QEmhiupQRCZrzAhrsJZ8sY+zSsA9fC9eP7PLYZEAwSLIyw0TLvMA5L7EMFI
eWSyDfePmCgH/B/kOeA+qXxKCQ+3tQNZ+1rVZgXQSXGLRZplis/VAXAtNH+j
1m/Q0k+au0oCIx9M8DqZfJPGtSJk2dFgSbQxmERd/k2j+9g3d1G/6PmBp8hz
2yEPPnbs+0/djcN5ETegmtLnUZWN9G9+dWwnRYzIVvkeBe5iUUjwSAOUDuSo
kyWJs0Xt/gFiokqdOEJsZrAli6NKzi3PNvnY2e2gbgOXGKnN4dgTaKaVO80y
paROA4gEJP4eRsf/I01Ocv+ioYbrN25nTh8dNNo5lsgkFEk7h4tRti4I+2Jc
7jI5JDrfzs29ZLnOYXhXZvnOl7ICrNduYr/xgCKEJxTclPrn+i483G0QmbFS
HIy+jgwvwkAE4CZO3Ff5PKBG8K/Vm2xPiSoH9xc/Tv6jRmnC8Q4vq0Vkp0dV
s7CsWOlapldy2fozRrxnu8dnVPUMdbYJF72FwoRPcLGfpgaZia9O1MRp9WlJ
H6wtHU/pk267nQtFyCgfrwvixASFiDCm01nhb8DQVrVNWAxy/7OVvoUPQaWU
8MFe2zGZHVSlz1r9BXCJIVykMm1gddVMNcxp7xALjX0b47bVlXTzFK7h0w6L
IEdzD6yC8bkzQU8OBjevfXHJS27Q83qGToyzTIr0M3TlTSKASvFxujVUN+m/
RruJer71S13PfFGjY81XJU15yx/u6K/0NDnfFCqCuYfU7WWlet1wdm5Inx7u
b6mIXqz/c7ufvPmqowpOon9m3VJvFJ9RYFMf4kbO6v2XciFfalptarRKA78j
35mHD0rQMGoXLj1xjcdDoBhjmOlkGNZzRjbOYKdt4g+cuHZCte7ovEczR5vl
jA8bYjfq1BZCQIUhdGMibd3zQ/3eL57U277j6XRhXZxhBQGTXW1cMhPDwdgZ
vysI2aWJ1b1WVnNL0VnxcYmDFGpiqsmFbf/BrZlfGAu73jpGHF+sh1/hBZkA
f95vHpxNCsbJ6jb2KZIRg32P7GShbU8lQpePw7xd7g/BfVy1l715E6rBnzgA
OX7URQZLPVJ9tKjWG9BgaG4YNOursJhpPLObocWYGlU/G0BP9lsLfHHKc8Z5
rEA2BMfLr2bFKqItznX4E/Zl1ySt02caVTaUsw3AOhiheEocLq4ycl551Rpf
WPEFcjGqz38Hp7pEXxq++oMYWD5Qz0mnmHNoF1l48lzsQk5PtZ9IskR6iBTa
uU7JeIX/fI3UxGcug2b3bDUiPg48W88ZWakX+q0jSHthn5aUkQDn87MchZtK
hGnwPRx2gHl3mIF/joSTTbdc5R55UzMdfFyq60ti579eNx7Q2s5XP10Z1DH3
QVPhppvA81JRu2DEVqQMwB+Fx+IDVmrSPMrhrqjALNfxJKIEzXGxM0BwQ9O9
rCSrvnDOaQEpP9qw1Hoi789VFCS9bbgAzAX8TUBH8IoIZB4wu6CV84WhNPPt
QssuH9TZSBJ8MvGIt3I2FyDuaZIjFG8IHNQtHf+HcH91/sJJtQhiauioxqgd
S3Igg4CrIIDAdEaJusrFxf8hIs8AuZQ8PO1d9DIdMlxqBCt0AE5DiOD0i+6D
b4ZgTnhzyDCBFOAgIFZPeD4DbtUILFpeMUsROsrZhixJ9EpxvRn6dCHx0Iie
1xQpen/+Atv047jcoTkNhvdVMvQEEviCXRFsh7aFn0aSc18BxMyKfhkXoU+A
NEAD4tD780itKw6xDDQ9fG3EFijukMhjV1lzhM9WW2SvnEmaBoG+IAO0TidA
RN0QbXIn18QfjdOD20kcD5KyKTVf/nMmT0BVzv3xSnwtSUHRdMGFVbeYc/l8
mPdKB+mWDabZpnLps3iC1p3lc8ekw4z4uju57XBp31+vWwdrhavfVE2ae8qu
dv/+y3R7kXCayI3vvQ0P1THyYvFY2v18Gqlv8RAKzootlvUo3zJAGHonVVep
jLA29bv/sSgKixC1Ek30Uq3vIQiqBZr+3DLn4QymqKl2RcXAscXKmUvERYWN
Jr1NYD1Sl/Jt+35oMjNsuLffaYCIxrik8Spx/wiQPAkjz9Mjil1/Dvz5d3Ia
wiT3bzwc3jUZtR4KyPkPlJhsFPZRQPz+QyUvxUiGYUwqe/a0czRHG9FgFoSd
6Een5CktF5ZvNzheZTfvnl1TrprtESIEdPox0B+J9d9tSJfURAbd6i6P9Kr9
q/o+FEOF9Y78oFhDIzn6704XakNVghFGdkOFpfX2qJoii8asZtqSgeAEHybP
J+29YOG9GdNGEg+syg57ArMt1BvWeNu730OZKSEZOtkF7rulvWPdd+vuv1ML
X+DtCLiYpn9iXnD9jKqCnkUD3LPNScdjJ3XnvgzHfpbu2YCxA/0cxz2HwYhV
x//vd5aqsO27gSJdKpV1TsypmmtNnp3OO83MxvLAG8OF6WXiKoJv5ynREEyj
IbMYynGAsgZpfZLn78n9zQ3+/MlI2jyOMNERhz0D0kE25e7wN/u91P8raxsv
TskpQWBT4DwzGDkptdGG18TRL4Lp35ZgE/uELiwyy40xZJC2P0pXc2OdAbvl
HhLjutHwfX7EjoGTF4w1c9MESE9dT6W78xyY3UvtfGDpgofgAbpETbnsiaez
+6CjOKDt5onmkgGOlc8bFHVuI0q/NCAezZuuziosHrP0wIvec9VRDIrXtzQN
eH/S4z4GQnouu6OtaJ/trObLwGDnw7IL0vaTDeOO/BTMHw+fEEeGfNANLhnY
I4gZWEogWXxlHkp5VT39ruGPBCofQNR/4ha4aXbi1zbqvH4fbpmI0PGYhGwv
foFXOdsSxcAXCl3h3Vdajc4mKV1aHohOzwSmsThgpXZc8/ajkjyJJeR7mQgT
KE1tsFin8IcS+uNKa3o+M87ylo4vzXVNWbmIaBc5bzrgG/2cUN7v/IOh72Uk
FrfjbvRKPbUmBz9LmDp29zYvy3vE80BCfTTi50i2naJpIDIJkjuUnom/DZCf
RqPgeP1emoJPsWR5GFK/rEETg3kk5SbSz/rV2NgTD4Hj5WJqlEYvMemb8sRn
e57wC/UsS/NqLBVvtlSq0bSKhLgtee4WRlMW1sx4BJIwRISk0AJ7HWNKpDPe
+cby+8wVwcCzMOkskH7FMCGcInkxvoAl5Kr69caSiskIhCzt+2xCBB9ZKAEF
Aud1q/C3RS1zlPWP9SJDQ2sRFn8ihqY78ZC06828uBC3n4YVTcq9RqChbyDM
yMlmMIbqGgdMPvJUXyZl81YYxud1/SxOIwuEv5nAMYeiCi/w5wshMsbMbv+k
23ggohcmSYuHK2XufCXK2vks1AnIdhazbeG0yoPoNHVoubCsfGc3P1G2Dr2A
zEPCT4GE5U7o/w5oral491X372/Ju8Mcb2udVMzjH1d1/b7mqEMpxlWxc1Aq
NcUywdO5F+v5QCncHSvusHou9ua+H9TpLQgI1H4sGSZZAF1fe9x1+6d22T3l
/Z4jsvhcrAxsrzBeFLnd3sSF28OiwxrAqmg4/pkuNpv5PxztxRmb4j2cpgG0
fNGgyoOqMwxS4kuyBjFwdCHgSHA1y5WHmMWEM8fCh8UIhOkbvO/TFTopM0Ux
lvmypA2WtvttMkOCzq8whp3MTvujQzmf9uapt72E9J6Z2NJ1rLMT5OyyG+/f
u+lXjXuzxk108bQedFFIULr4L3ISQArkDQIH/8BosAxpb/R5RLmGQV45jODa
pNmcf0vxUJw7R6VoLhElMRq045dIsaME0TdPEGNwXLbRmqXzbeba04LXAyO4
VTssCDDL+yv6HrPO+HrRnvE8GKvkalQ0xew+ZUG7nUqHdM6ideFxoK9nKvXG
/T2n6v/75KYV95OTzL5sDHe8mOqshOJamiAbB+5VseCl12POXzpFj7/TZDjp
wzeba4hwyXNTU7+65/zPaG/wtH/FL2PjlWDW3ld7cnuwOuaITT8xSPkVCsRI
Kj0HQXSq+28mYb/9zXR3xxzmXBl3M0Fm84HpGCUcJAaDAYxc9BAZQ5NPUype
PWQ/ZBQ56MBom0h0NWxENWf9Nsb6U2sOpq9HKsvDVSfDfRMTq+7XHJPwNvjA
6Ex3VRdXPSTozVTbh7qJNv6pJ7C0wrw96c/5RBQUmV4cQPchj1vIcOI3WBEB
fdNpnMCl8rG0b0n8RVkxqyD8kjhHqDe7Gy+fhhJPzNjW5xQOqYsRq1tdnxPv
fqjrX8L63tpFpthDL1Jtj+f3B2isEhbRW/iSWNgh9elQSatPGxH05C8Y7rmV
x5lU0mvMTawKzF31E80w514DpzWPy7TNar5JdEpQ3ntXzAwSCXuTGZ5WU8lO
0/frg5YHmT4jw9HVaa3BOLJnwNS1rLxmZshe6OsrBHFuR2L7wyLKgESS/IJj
C0kAPEm8yLCZi+LV0FQY0PEdsUVo6O+5wg/QMkvtTm+tTZmLhdeXaDaA3BgZ
NQKQureKfOapMdzw/QrLNOgNR8JFrP01hRDK/B03poZ8bHCNyJF5b4eLwevO
dyynvkteGxZAwSkswttlqsdpHdskHyPq4vATD6GJob6rv+CPYnHc4HviEDtC
5LJNc7N2H9CeAE8hZcN6vXepuVI1F0cZ2leoOWgIdIGdWxargZN6T9J6F4OO
V8SiLL/40Fdn4zOn7DvnAsQX1bLnFGRjXREk5CpqsdIhL22qiA9kA3Wab6Ur
V3VA3chGbY9BlS5qmK6pTTpYpbkMk3tOxUsBL6KQWqPJ8EXFwQqNAZKasBoI
ckun5dO8gUosAPV54ayGkROiwKvtWf7x4MNrAdv/cV2/DNODyQTq5FzHik+k
Ry5dhxqgpdnR4WQubBSY8af9yRVLVO6/yHoQT3NSZ5SrM4n6KLz8sw/NafiU
WzIf+5zsORF3wD6s3gaHqgLiExUgrIF/fGPQ8+r5U31L5XMfUWjU3qnUbhq2
BqfRkA5rtTgIVSYIQi8LEEPdyYYzNzYfDvrrdu2mOZx3ga0Q6ztZujZjNMfC
HAPzilAHYO6gL64fl7jrk7hVWsV9B+GabcEH+rHOo+SK2QozZSAD5KMlEM5g
3JxyL9nS85AVmK9DuuAp8yGiGKR8YcrbdgQg6nYplMMssFuoBiOoRCXBgVRx
A6mDy63MaI/ZIc48yYFoO0bxXEx8qdqHodRRksCuIIZlsfrdqKg2EENg+xcI
c0hiGUbRZp/W6CBgIOROCG7V0Se3J9OnBQ7tZjR2cvqlgT7kRsygSfcGIE5z
YCzY+nnroqi4dBZe9u4vaQV949bg8B9J+bVKXgkSfHD+vJUa67KSCenp7NF7
+Ib5FSAUedoOt5DziKKPIIrcoSP+hZ1Dd13M1Kbllx8jI+mfOVOdoXKi509/
RwIUwKwNggP40E286bji7RF63mhkax/sKFddkzEkzLoZk8y/5GnfZ/L5Gt7L
dNuJHQLHaxslq3X65fT/f66EMSaW+4KNMzBh2LIB2jrYbpbcsG+Na6Sue1OC
s7emWwiTIyMoRb9C1zGt3r4zUPe1OIbrjLZI6NMm8MZLVyRi/OJtljvUebW6
7bz0L5Y4FhxuMZ2TLXcSCAR2PdaVkGp7vezKt1WKO09p3lLtROJt+ky5KSNu
3GmYvrF8egPM4B+ymXL8qLO+lr7zWdsmsxV8t4RpYnmtSvUZO9fQ9R+9gDuJ
Q3OtRPIWrXnGgpjT3OrzK31I8cxd5wzPRqgkjHa0A39/MGBI33+zGsCJ0l7b
ScbHLqr6em1mQfQuWTKiEHH9bnATEpj4wqOM9R4Sa0hxpLRMY1na7qkgf3YU
5xmhpKcivANK8A138v1RolTO9PiowiXiPT8/CwzqN8f8A1OfkdJH9ZYtE/QY
Slfl4l3U/k/rafrY/vO0s0ndvxd72aZ5RBt2YHW7su0E/2u/+eQd4WkE1Zp/
tazyjT10VoMiplmxTHPN7UGu4+aCgTJjulXjSrx4hMGe13rN/NKsohpcGkTP
d3IYwB2XWy9VbXgzI96waBcIoP8tbMKyaEhlwDiDD30pMzjtqZvIwmWU/qYA
e19FPd4KrkCjfkWZ7bUH9Lf7N4wSNbzfEol/NZD0B6O8O9QD1VxauaO6Xaz5
Sjjs5Ldm7xbRYJGaAnA94iFnoKYu4uhF1cIKm9/ufO/Ty3HB7DkaFXnDMwVr
3a8IGXl5OQp6nFZ0Xe61a74VBQOXQohT1C6GrcZ6XaxALdue2op35vM1RCfa
XA18Y8nGuY6mJ523Im7aq7KY5FSLdkLVxsJDw28f58GCqfGj8WVVtjduzTIL
71wtd6U+zIlxbyIOldnR/9KiCqW5XL81LXRF5ZrsWH+AigrV3MEc5sXHZgeq
gpnf2ztUK0ec3af7UF31PJRAOQ9S3jl/aGUZVACiVNnTBNSqUVAZsL+X0fhw
7wHD302Xdz+b1vLvS/I4EnuuSXeFvh7zjGt42+OLsoGVNNrPnuQCF7HvHz/O
IMHJfwAB6AyERV1EMPhXBa3BG94a16+KXbiN3vkvIehdDstm/8DAkAAc9FG4
GvEivcDqhMrdKXncOx/gfA3GbqP3JjOmY43mk2ig/On0FtZ4cd3gQmrOieGd
MzLOI7gnN7HGFMIINq6raPKTndKmgn23d1il5nR63vQ0Ws9AnDm2aHIuVphQ
ok4m2+gLtCRXvqQxsoJhtnxpDN+qrmyK6IGKrRAjr/X4x8TfAJva5bqLBvWM
QxXzXqEihC41BJPK9PUuJIsT8UvnbPWmaYAk3YRS+sNXc1Lb0b5DWUtWzh+7
iyVS6vZLNi17pojSHll98cOCPUL9RY8AcCwksOXls3HgwqKD5qqKMpgfV0D6
5GItwt1rkkeWEY5bQXj/Ew27KNnIFtIlNRYYNcc/8QCwEPShZ3Idt1v0WujE
RCQxWyr/2uA1L3+v4qEWkKQKOf5izRGN/CySqh45UK7bLX+cLOKaygybwqHi
1LrKT6xFO8POjj5yWGg0boSkzunIZFCOXTYGJn4it4DOYaeZBOGZPkXpa/GX
h7vHemMqJsNYg+dUex0UjtaPfVahPj4vx3dSQBZnWIeLD1NmRr0fEb5nv+Xb
7V0ahd2uoDaHNzYRi4F/ZP505uUXXIpTBn3R1tmCZYTMqprY6ktKQp8N51gn
JgRmX/Ydfw0VTBgn01NE+30J/+8VHLMVMwB603IiY/Wr8mySpfQEzr7nq+kO
x215DarKKoKSVjSmPJ70QyMLwpFvEuaqRbAc8xGvkT6KJXZtUddb4s1kC6X9
vioU9rqBw1S7Wj2NoyuMEAqFQzOadqeA1NQNuZiHdZAqr4tdCEibDE9nkaGv
Tgx1QL1SFYh9b0LlggnL3oxE1b6U/Jn0Vd0IozzEZI0YGzgVhPcn6GlNKzVe
S7hIV9GEpVvxQF4wDwtwjEMotE3CVWyqxjlD7xYphUQak4ukjruwjGCf4UBx
CQ0b+JVqwje0POOXgcMF618Qs3zK56DlVbQ/UPrQ+eOR7PvXIB/OFg5REPCz
NPLdAKzo6ox0WgqcgLTCz6C73ggQTg8xYMhCjEGIzKOBGIc3J2+zG44wrQDo
YXF3SFlJwop81H6Bv9lgfvntkuou6pdCTf2p/Ek5x549yvcHSwub6S7hcPni
d71SqgPpGErSgr9M3Na7piGjWblZnYSqi12DUd3d/nyBOythiJ1pckAaIiyS
nGMnfJqlBAM1XqM4N7AEb+5gu7XZVfsaj3cUD4FWyQ99/6MquuiUKjTI1CBg
D1SehRqhPyeplzUZO7IkcnEi8oETlao1UrAk6FZ8Sbmf1NG4Z3jdvIYExmv8
aRnMvWJSEIwSVv50urweGUTHu4IvgOYrW0Z/Zgk6aTre+H7h3CGGf5xgXs+Q
tLxGvXzAIJgKgeX3T0lHUDQgjOZ0cP4PqVYgYfq6nWIhbcX/o2k3lzkw8Y3n
bqD/mIDm+9bB9onMYX5qXTTCTjcSvOmlwpX0ah9RnmhRlOF8Zw6WO6MVdAfw
wv8w3huGKHKKRwKpkl51dYC0riy8pr1vUmXZOTIuJvZa3K4SnqaUjp9grWaO
cfWbvhv2IjF1c4GSbfJyhYU83agxvDgU7AxGGDjvYkuuA0/uz559cUdyjGb2
3Ff6COx3XP5/rKi3T0fGiDmSIQxkl8/cGGVo2bK/MFwY0Q+EeKrZjcKCn2Nf
m4emJErtDs3+hAM3KaSx4WuKqx24vfCD3J4X0k3bIhUhNT8Qvvg2nSLgrcj+
2Lx8DbYmlU0LI2TUTa5PtpVWB1KRfR0A8kDq+C1x0jq0MLIcWopyTr4Ksq6T
/qw0d1Q6M8eq7KP1fgDjZINXRbj9U2tJBi0nQvRLbJi5jjZ2PlhqpEHLoEsg
9p3Jr4bxdJKA5bIsYEqVMvNNJF7/7vptpjnPJ5tr+JfgkZSJiVGSxgC5ct/w
eLQXWhnTlxQ+Wc9d59sUX4TzBHPU8aneD5Bc0duH2EhBfgcM+uNzkwGwDj/F
1+iAdn5F62caaU7wFx+BKWKWlsoZKVzL3bEpT+d97k9muzxc9kTIb2lAs1pe
a6z8ohHL0qKAJ9iSYGo/ahrP2lMfy4hjXcRVTDbf7ReVfbIujpIbPxBkiHkV
hbG/sKInS3NMY4O1oPuHbsCcRaQietapdIh6zTye9fELma447YTFDqurF6B7
VAGOyVMQdWBY1uT3ZMixZTxEEJ5uZj4tcjgkOGcsdlbggwQkksK/GxnE6Zow
7ADTVRQABnyr7vO57Le7GykKOsyiTGqK0HVSTfgr3XowqgAPpqtmk6towpUm
VzqYB8IZdfVdbD+tzdvQPxA8boqnSl9hrdeeqjWcw6q+xaKUporSy1YoAkju
RWwrfvth5BTXneHcI+NkBpTEGbaQFa4nCKYAC2YpHR174dnD2DsEvo6/Ho96
MPne3pICL+HX33JAJDBMC+AkQ+upA2SUYPyWJZ7D3fmhJIXgUBct/ATwEUsx
HRTBa3c7Ae6i/WbF4Osea+5Xppkc1+btDTvm1mUBYCzsI2w/QfEF8S2tJAGS
/TGeM8+QOnSZovOLgCWGhtPrl13bYx0osiC1rLhfhD70fnMZtciaBtswMSO6
GPF64etimEj4V2P1wjksJvbcBEw8hOSmzKTBLeVATFmRNbNmdnIo6ACUBp5D
8/ek6gIG+/q9c/0E+UfeJy5V1vr8NjgGLKlioCmujbYylrZHNz0nAbca01D9
u7kfYU6xK5j/AYNAME8FQ/F3gM0zAhjGC8JZSKr8838DJIWmPCQn0uwt8ZDP
oiVO8LBbyDb9vNVBOKdNZG8ybX3pMdfrs3KAP7QWcbSxPPIAPHtYP2x/pU7z
hXMIBDCXAzBxcgoNokat819YiDBFRE2ip0HMYjTDq/9KoiNAKC6i5xN9HGZH
8+fGDl5j8LVqYMcgioCduW5KjjeCVgyUOEyn20gkmleEI/ZAUMGnlzcJvHTG
xi2LEvCFBsDGCeCBM9z4TA/oRto4D2PdC4rJxW9itMsRVviX7nR/NzQSzHro
jMjCmo7UYsb3SsT3m1LJ3PgW0ovd9eXnLKtPlYDwoNGEoA781HdLg4i81egg
tzaGnq6t6ZMR7v0PAAxSgKbi9MWOccqeDv2iG2u+TmwZvS3FHXXgfEd/ptCc
Jp0zQoCUSxkaHVAjfdSOr7jI8tqesTFY7U1BM2ACcuiYvqe0wGxaZYWD4L4W
PrUiLmFBCbV7nTNDdEpTzXC30uVSnDLk/tos2+Pzw+ZwqmyGKyy//dA4lgVv
qAz+xpv+o9TjoVVxKhS7pbFKKZ3We9MpByuyMn96lIrn2nV3BewBA+QAVY5q
PM3aUOW0pyxMCbLo11S8wl2du4Ev7V0LIj/cDYczGxgSRULPvCeW6ab0RbVr
LOg4nP7v58PBovm7+fhSc7CVM2KP4Gg/6Ob8nCkOVzBBeeXPL7nuxKzzvtWY
Su4MMRSmvkvb6rZlejnIlG2Y0KZlBurfPrDf6TYedQxqhwpBYHculQwZ7zmF
rHGuxkxpg1t9e4Hiqhc5hfrF5cLJrQd4wI5cUqmXge/M1vFcAKtriRk0Nb3c
o4EujYXdwuO/DS1fcLTfvkcF0TOZ2uCr6HXWgI8+KHYNBDgmpYz8ciqqI60A
/zGV3tR7OuSzKDy0cr1+SN4H+tdpAPIdb/5c1UdWn2r1QiWogsPfxJgkYtUg
eKOCHQ2nA+SPBUKpfvCnJBryz/xZU+9nadqgKVqy9JB0k9ST0jcXxKkl7rEU
RvyTzdRphEDb9cd5RrMFfvzoyWYvAIEIvuG6ZrMUEq7D592YFKfgLLJMLTB3
ygQTxo5Waro5SRjMxzVnj54SyMzeaaAs3jArYQMLhWnPIzZ5WlV5qFc9tkX4
GWiLzz50cAcfPsancUfHkenMMlXmFxWRBYi+w7sNYEcz/zuQD3YqRSVpPui1
xe4VCz9g2nlOF1vShqb1i/dEzm/JJJu6d+4YVss95mzQuDF4AJ6eeDUtFFXi
CrEesNUzpbuLh7gdIOC4xrHtbW38O0ixgCan9oEtMtXtn6wmhY9u9zq03G6S
3WRXvrf4SRmZqAGaMhJlPfwAuXOllPhU/US+l7s3tKlUrRgC1HloCQcbYCh0
5W6gecNtEKZBUJCJRgm/JHfct3OTLAoRaEoToXd782ZpQi/1cXmOP/rb8SNo
JtaXOrcmEg1mrdDovbalDaACHCYLs0yDfQIcgBnIPhiqKBZZfpcJNAKnOUkm
ut+0DdOzJoRvdKxx9xlsxd1SyyRJgpB5FQ5tgfuz2frT/g5V6OvvYdoG37e8
cfysbS01qqzsRWIbdKfSLzrgof8mpDluGJvMzjc7phVRnOZ+jMFsbALtoqfx
hrjtyw328krsJ0nSLi+LEP42viCFYDqS+pTCIAHUNBzd94XVcesXoO+dvCGn
izMUp0b2mOcacGc06+85k7e84+Wn61UDZY4cEWueGBOH9XLvLzEEtZKbQ8Ji
tpsjWAijYrNnywCRjpPxQDsXZdGyuMWhfG5f/PLcrBrxjtlD3V+vvHN/nzK1
dsF/guIKVc3XpmKpZ095S40pMuYxSFUUUYEXcHNgu+wckCanAggpIOGhh5N5
i+rNzaUMR6fZXmQBybVGkW04DPgVPd2PuzLKFtk+DIte14iNqHifN8yHie+G
10BbhFYk305MyBbL4m3XtOIEEiyy22hFJAUli3edjb7EsOawldOZ3/mfgrHV
SfucIumvUpYV6umo14hUsCNlQJ1PiWypc9D2Va5fqe59HqxwJwecinhZ9DSb
QUixqWD2T/1Y9sRwTZddVzUfq98gV0A7msg+uk3jeOlrgSDkGwcdCDOt80NR
WprZf//ZT7TGSyz3KFTQLdOM8KuyLSu+VWjjxBBt7JpuPB0gNw0rAxLaxnnv
fAIASsJNqbWYPtYV1xNh8m+3WjgHoccMj6pwnYRHVp488BHyfFsKJZOneF7K
oE9vINdm4txZj4jKPeEUF2A6Zze15ELWDzyVM1JQ6mXvwYP71+c77dH8GzNI
+wM8efPLezVXcSk1zqgCC9m7wGSTSXH+fglarzkOGYErG/eS+re1L/xxqdv6
T/Z/mfCwyzHa5UQIDXgb22/8unWsfKfrZczBQO9I6L6OFt/shBphDdiMpB7v
TQS2OB/n6xkcBZkIMmEtn5Pwd4G2SW0C5KYbJJOAgVptkdRtuyWllOKnDG5c
VhP57PlEUdbrU1HxRgTrq+2Zie1xch/0DLQeOlVmlsBTsz8SMmIw62Un5JWa
TN9TrInlP1XVIQ2CCCFb4vYU4DcJ+RMry/J8vQlRUUUzIEjX7gTf338vHTgX
wLf7Ae8duj9/WUFyEeI/IJI3kOcT0shkIMgOzRkpBAuSKgF/dBaM+wkV4tSS
pq0WH8s0GX3u+s2+37c43jcEvL0qZE4vKRLzQvJUF8Vc5n2Qz5B9V8m02Pdg
hUTa+eoDnOsm7CDk8IvdzLdo5RirZdw3Spb1QyeklT5FLTMVdolDfIvI/4Y7
RvGFbaXB8qosBejKb3GLDvtq2TGwc5yi2BBa8QDcff9fOuM/abcLsUST/NMB
lJBoukCBo9BzcvhdoeDVRyTDkg7bdG7iGQZZc0G7481iMkJjJuT4WuH1Fhi0
keKQC734SCnP/WgxWi1LPbdJOVkH/634y8QaCmSs1hL/LYp7OAm9ldjUI6PT
eIsElB85LHlZ34jeZMfgVQnel8XRY7ysk1FU98FiE8eJXN4oJcRorhAj1S8A
swhWJQ9H7XPSCN/AMbqhN7s8X5DkV4r0r9WbugVHG31Qc9csGq4+dshdUvpy
r/X+w2zSfTfRsC3tEpSn531JshOExlSFvO5lmjAsFjUqyzSsd2ErLZXHihPC
srxF+ezVu9sGYtbsrMRSgsZlX5W6JRjSl4KlkILZ7YPJxFG6GIavl/SUEIVq
4AAzAi2omhn0BrFre8bttUrgwrwGDQiCC6IoIK9+tUCwXJAjWsqHKf1tdUFM
cQufbc0bf/ZizeeKNGoLiy5BA3S9m2dBtkW4a16UK4LCyNxezzR+6HsYsA4X
OUGN46Y0cEamDdeFF4tM+QrZNKj/1PBcWrasiHJ75Xh2LZOSGwVDWcF7Ed4s
E3uHHuNZQnIhXOwSxW3SINcNgx8FitUbkDbG41PIIAjxmHseiMXot7+lYn1F
4bx1Nu/27cPkIM5Y33MOk3y17hFYhTgRom6uRNI9bLoQcEud+uyVXPpFtb+U
DGgDhKtP87N+3e0O/XvJVttVXlaTy7W54uZ1N3DkU3Dp2X1ZLkqEzzXSrMRy
1NM0rWcPnjcSPVCdMQJp9v17rkVuAx7+l1Fswg7pkJRUL3YLHMX7m1H5vIFa
jR36xKeNUNQVWcX1F8Vpi3Y6YadJffDnirR/aZ9a7DOavRE8MoLgIy7kBpFw
kNxFVc7aksAvCBBkLAP5kjjHc+ALNF/2Hv4bVeqJI7JKTopxZVy9wlphi+h2
8AmxOv5t3Qu0qOL1WNw+LnEQTmaUZ6tlcflfEJbtaUgRhoE4aiAjNjbcyH6x
1ZURVqvPAEPccWW2f+nTsd1FlFTPFy2rbNjMgU+nbMycZ86XEiTOSnxxlYLA
cjxPnv2FRSNZpgROp/bcMAt3p7qmZ86Msg1rvf8fym1q9ZPz1irtIcJyFxjK
NnX+WJYyc+avGRgeW6IrPpeR7YsfKLwYx0AWx5YT4xGboFUfT1QJAX/zfbZP
lYlqQ0uHFZUxlxxaLuQkAltE9WX8OK4yRfWnr72ok5+qxmQ+fEaxeAz43qLu
Uymksw4aQ8SJYLKNH5GHTcnCHhziqWM1liy6Fb94bjwrEkGIe7IWvJfU55Fh
5O+aEDt08wUoBUvdc0xfacAu4kPPj0jy8bn0OLIV5/LzU3Kx6LITOz6NtPSj
G/crI52ezRac2sl9FWrTQiL4dwlr8WrZGcJa5xS2uME/jNbUzFqL9Ac9b1X6
W90kUnW9bjHs7/iJ4N78841QFvPpmlhbJS7IdtbKQSpmbbXV88mrleoon83V
SixFmtjXcnHbp/L5EvezMTuq/95FafnUPUQ13hgTcJFXgZVpg0jrBBfIvX75
bqy+aCq4UFkZJSSuxFJK+AmR3dHKkpxUJUUpr8pIxYO2zxHjudiFqrjd10NG
ZkYHezXMR3IaL3rWGT8p5CRrBdheueO4SCznCjw0Y+I2Q5mzXPSxDa/VW28/
+WkuzUVhxj8YMZBqnaXv3WYjjjp43Tlw/7fUt5N1T6bzYw2/E0hAzqSTIr0/
iSgCZpH2bZhmKFvvTseUy0BZjidr6SoH4kcxVkU7FUzwK24tHAduXZrSulmH
BCua1BRJc8+myJt76eMw7QNNQzZQ5nCqe5brBLCdo8kQV3XhLoWdicJxSvrT
1G39QjVzNLVYZvkDu3WFW0JACIop/gc7BkEkwzVpRH09/z3+0RpvUzooPrN4
n4IZjMazuX/0S8m406el1cuEwV4phaTjTNIw8NZch0A+UTMEVRwiNnxR5pXN
aSQrsWmKUlzJ7PKNhOSFgsCowQgGN87Q3CBqUr4FfCLXjZ2g6PojcvobPlQR
fZvsr7GGFyRcaB8EGwatat15n9ATQLT9FDVIkiZe6hf3Yo6MplYUB4NQChMF
EV0kS+Elg7pVuFl00M5hINitZ0b3CJ+9E9945ZUzgEB7IWRWaLxDtAbiGBbm
4N8xk3oN1ajyP6xKvUvIenjjW7hLCFUtjm/FzNhajOfjgqpTl6Vu+cxBUxZG
w4ufglzJDNJkxfvlk5+t0//33SL3ASN6gECAjPg2+EMen992ff+E8zzkLgrH
wYPrTDFYo4Tjbx6RRg+L3f9Ulx2XyoQ/u2KpZCb25xZM8Pirc+RewdDuZTUO
nMemU94FPpo5wNgUJYGuUdAfE54FTriI7ZuI53ALpjUS3Ew8qsHF40rqA8i+
/IYKlpHfLQFRWXBFrxjDwbC3i3EhckR/2gnQ5HusQiw69RkQTzB/ONLRq3k6
oqHMpU+tyWudeTj8ZPXyuJJUQVp4A0HszHR85og4umIA11xlXdvXbWiCz3ZW
QuX81wFQ/hwBF6bEnGb8e5aLI1h/ND4qjm9A5RG41Mo+XN0k7ZY2R266M35Y
F0oRcWOcO/r1CQjeElkWJTRgn48Hkkd5SMrN5lPggOF1nLKcvB70TQ22OeWj
VKbH8GdnQBA1vXzJh+NPmPpqevoFpytTTRNORdvSMLu+1JJ3uZyUDdFCQE7t
x24eNXs7YasSliObwGcIhes8kiupYNikJDwClxJAT4M9hMhEouxE84aNGF4f
urMnjekNNOsdD147A7Qdq3yfyNsQAxEg8IHt7nrSNryUxmJbS4OGzqG19fN4
K7HS1Lil9cius95rTDX82P1ianWvS1i5wNjxvzkiZMIov5SmPZcPcXurd31y
9n/whTCYGov6h3aw8uw1uMbf0sNVNwyef4TmPqY+JV4rpNOx95PMy9tyep7R
8JLY7MzljfmZdMvm74hjvl5UlvOQEI17fPVBPxmuot541CaZD1WJ1pbxciZi
7FUrVBD+Y1hgY2tAiBiHAUQwrJN2Hn4uJ6o43fmEpDOdnLcAqQDKCaS7kWBA
jJed9eW/71pEn3n0tcig2sbjtKHn/BgKiBJzvRV1pKWZWgxTQsAnVWRF6Bip
AUOW1zMsBlb7WTM1hCqWz3hSPNCaW/E9BQsBeNjMg6pHv2QdOZfKWMCegNgk
q4mpzq79NiHxjpxxmyHJ8MTJW146dXdI4FELBbIfMnRW8yrwrwG2gO8KPCYk
aK3erCJTzmBfKUcgImIs08iaq/C5DIO5aYSFW6YqhSyHBCeb+evixf9AQfmw
DWYYsjmT/yYq/Eo6jC6khwq7js6teUbbkvmAAd2/itpuuZIEMi+fAvvci+dq
nrFQDGILt6Y2a1tr1naq+NSSwVVAzM/x8OE2tV2JR1irBZvmm2DzZQou4B0D
FdaBKhq0VTF8mLdUjr2aQci+ARoh4AE09pxrak1seQHVWRmp6wKfoEWAauws
VyC0HPG98stOknx/rudinAzmllqg5PzNmt1DNTAPs6zJT1ZE4e3EkSYSEjAt
c07et5yZ1Eo1tFLkv7uedCWkg0x3puAUwRV+Ho+Mh4+HhGYvI7qYCKgSsxHu
613xlhJdlAQ08N7P+NyWnxWoW2i0Wi8MESTeQQWYstDLGzPx66fRVyF5gDyn
6AMylj8WlFSAhpjT98CLtzO8VcqVNiYFF+VEbxy6ExMZ1v5D6hDDlsE/S9DZ
pM9c2stOQ64R5YybZvC5kS+0K5Xj4ZFy8KpVscSuuNdCjh8fnHsbctpt85vv
iJKWVjqaVPjMs9qRWAWLZnTyKF91iUXhS6jG/5T2vWWf/Fpa9DLFYzoFulwe
PMxNf27TezbuHnLjOKPpyK0SePbFoEMFKRCo54NsAmBYjmflEmA6UQe/sGrh
4v2f9B8jgP5aihOWfrcjBUX9lEbK5w7ycPd5KoZjoGDl80e98Z1t/Bje9b1y
luGoIfWbOQ/upqgduv6un1Z3nllbZ641aR3X6rocNYuOT4qOKH0/1CUqIOnK
rClNiFnLPaTXzc38O9HTrn89LPZM5fGSsFIQggyV4cZVQ68wh3U5fouwX0zf
BGUHBMPwSa5705y7oxXMq2OnaP/S2uz1HIacioY5LY8ScYSoHp7n+LjWDLa1
QbFxuVxpurhIXTo5GDLaXtMLyE91P+AMQylGcSpJIRiAOGy9WmyRX3vRpy4j
AG+oAF6NWl0axZW+2rxzUzIy3cfmKkXqV6LNHXTDX0opgCkxCZZE5frPjl83
cNqa9Wl9KFi5I4QeLFfiTXOnX0K9Sb/74hOXByOe49nAr50PigZ1t9AUCx+a
0HQYWHckroaW/RXPbW2f7HeOQT30+GlxkY38Q/ZQ/ESygy+cft0OOc6k/KKn
1yPjrtdbv1EqUIaupu8KWMeVoPufB+w8EpmyKrfChtTu5IFm+ajsMliwEI3R
EhdYwGVGRJN/Vo5QG2a6bLikTT5ikPPaG073Oi6sOXDWuuYg6xWfyPdhZ/45
38zEbw9krnT7sRVlE5nc8JU9mEB9VzbFUr7HuFpR4Jj6uo1GVIZ19Rl0mqLZ
uL7DlbCqqpQAYaofvCIlvUOe0x1PVlkHf9iXzI35CZh7uvOWBXuM+1h7u99+
SWyImGVEJsmuT9yp6/HFF8B8U105ZU9JKju9aEJTmW0qEoBtlF09bkaL9t81
1EF9++sR4TOBMCMZ2lK1I0+giyp6YXz7HFOq6nPLtWxrxDTTvtymMfhke/IA
7F7iuRPiZEyJEliwX/WVpIdXhYhMBTDdp2Af6JT7u4jZvwvNsOtsZoT7dmUS
dPxGTwTjhi1LSeeOgoXDPCBvEHrITLnhwVyR6P2+FCr9ySOb+qwhALrVmPPh
DDvDVqApDqRFe2KAhMp8yjOfyczxDSqCTUu98xBdCAxtBWoZSIBAky4Jmtsm
7nNQSDAaNXXaaU/jJFdLlw3PbiQcSVquNz7V+mwLJdAs9/coM+IPZVWxMszE
xib1N9BNsqbhyYi9xwKvPJ+Jx+lcpKu1ST9pI2PdIONyBxSESVoLNMN25uwo
vFFQgWFHFh022cEWQEXxiI0LdzTaipq0a86DAd6eCY8AOa+UdYC3S7FHWe0+
7k2pZ7ze55whVpkimzWFs2NglWkchiYDOZjLRu4MoMUwwKEvYOn4zSt0WCS7
9zC0w2H8jr5O7C2goIP0ofhYUBbgodp9rrhcIV3P55nwknZ6iPEQkpM3/qhd
3DaH2HY85L2pdSaMnRfrSEpye9dmEui3TgomPE8rOAxNeciMFIFiZQSSzJ72
qU7gX+fldUyYNJ6sqMqHutDPG0ViIUNh3kXyo7wr3LwFbnVG7IEheV4vdAnw
SE9XuGO8EbwDaj4wWAtcPQmhEMQkl410R2CIhCJeMCeoysk0V9/5g1a3gGnl
AdhBpUxV0PuBvHZtKxuthvu2iguNZGD0OXdGPWRebALIYpTJTWh2Xa8EMml5
zqm44i2VvGzw4tPsvGqB2RzrGzjQ+ZkZXaFOP9rjH4h0WY0OdSv6HKccdyCo
HNARhiMyxkneX4oSq33TA14rpVK5QhBumCdbV4gb09PXvgEX7Zw1PnGUjmx1
j3Qp09K4voq9/4pVvX3lSI7MwTxxHsGjgOEy5L6N9xJOAG1r309ZGZwvT22y
1NESkFGKQ36nACRLIHBqNUNo0j0aALyhSMNCrqZN5TD52HIeouLLnjPtgeLD
19Ez183fQ21a6oyZTTFouEJVRRAB4d3ioAXchlOIdt1JurFkov200/RGIAKK
GvwxGKS9U977wUvkOchRkUs9/LN38UWby+KT1wO74/qoXUBIJfHcfX6HGp9R
k5c4FJT/OZklYP5GTOEjRUPeAk33OQL98+rB0ef51NgfPDOSX9gigWzknp91
jekdhw5DRCFN0F1RSK96+ASPKQyrwtjlcKJC4sNFNaeZUAcvbAHTpqZabzmn
FpGgmb3PooDG2AONbnhL6TIBORBSjWO5UwHLObIjGFNlSLL8l8Hvbo+Mwbq+
VCJtqBf05eF/5KJHSzpudHy/hVIyxHYQHWOv/uky+IbOhAS/cYYQlfQH7aFh
l9fKqkhXf1OGJnlsoZwQ03T1faGWME7VRW4dMT8srv/oOJk2aldGKHoTB84J
yGjxWoQ7ThgQAN+RK/JS371ZGjXL4IRrU5cjBwBl2sCL2AROJbwB4tCkwIcr
VCx5FhgKWpOBWr0eHHUpkrQqoI3mmxp+L+uQLSyWrqQFawgqQ8OXxgAZjX7w
tFVKPTmy+6CUQMTawICWxG2L72XlotmHZvchf9djeSEB1+C7puigSPAnRgDU
NdlGGpPlpeJvVz5uDciKxT2SBPy/qmoEpKeX+HDwZkJix/G1KzZqeTVX5mSU
aMYEAwL2RmzCt3rq5Gu+TtK+u1sKNhkWbFnigeOCIwKwj2vNPV6NcfxN35SR
b7/9Jqv00653rdlMr0xukDRoIl9L92gW3T3K91PvdjNRbvX0rAi25sjEQQkt
pPAW/CtmhTe+X1HkN6gv6cvX5LA7OAFOmwkGVnNPwxLAIrDYZ+EEy0c1yHkm
n1wLygwpdV0bZehR5Iam2sY6vnt018yvm5tPT64eZBKMPOjC3MDXzGyAml8W
oUdGbvGpFJpbl8glBB4PRh4oczhgC4ya+ZqeuHb6BbKQ7dcyExutZpqi7Ytc
bZt5alM/PRepYR2P/WXq9fjHpju8dTjPcNn3Gob5r02pulcEDDClfQjL9/pt
DaCDml71H2iM2OPEzKNtqMmkck2EtU3vzeBsp3goEFL2qoT1sYjGmdTJ1Pr/
rMbM3zZ2q31+CgRvTT7nj1gASVS/D6kbAhji1faQg7qLDEtDTw7N7KBMlGWj
fWhD9CgXF9JJ3dQVQ/msW4nOQmIIEX2/VAiHdrlOJz974qJHg/Acd6TseVfO
yhkS3yjx+xFmNKg3/er87R9paD60a/a99/T+dAqM60f5uvyC/StHDLgT1qdH
/0i+LFkZThGIQRtq3meebtuUOHxuNxtsmh+EXdd9FbU3PSk2w7f5skWFnrUc
RUmfVlFGpyegd7wbFptI9TroAEHG1ELXbv+tMhqk8j4yh3+IMiw07H/sT2U1
k4Z438cgJd1RqCCk1YUsoIQgTRa8Fs46Pb+3mVuGl2RM88O0h7TXyde+ff48
owAcN7NEmU80MzmXe4FARivx1gczvIhl1IVmobO9B+fCUDRL/+sL/5XQAq1V
iaJ2eS99fLpCr3VyVaTB0ydfOxQ4DwdRcVsa15u5zj4bHuDzIaNW4xhGr71D
YLLpMQddTUYoVnXUtqmnjLFcumykctgQCBJbCRWsvK8R9uXZRRhiVBFa+acW
b4iyZ4vB+XALS7HMNGhKrc+T+Vtydnh2o8p/eQNXDyTnQNNeEIlBQBWWdqSQ
/SRu3cqlqAES+Uya9vji5BeqG7kxBRtrbYEQdD9IoOIJMvNtAjQO+8MM2dTI
/zg6WKQjc38m0fSZcUiXYCr78F80RQCnJ2jf+C7IXFxaLzY62v9xvCOcnlAE
XaMpMRfPQBmHZr1eIoUd0Mr2DQYJpbq1+35A8FpCc3ecI8moaVaKqvmUpKp9
6u3MiJCzWX919lFAL5FgFI1LWBabulj9THIu6tj3LItBuak7uc/62aCz/n1X
onoYBkThdJAQMbrDOmFrNgKmVwbTsdFnA5kBpyR9kReKBkCOISBGHzD5LTJK
PjHE43P3yn1JrBggbIl9LPgUPX0Z7aoaJ0KDZFaMmHinEIgRjKaqilHycNUb
KdXnmtD8VBitpMb3hwnbmf4reoFV5jnEfTkYFkyg5v08+OZJdatQ8pEZj4u4
sWgceq+cA4d89jfQPl5UZ4AfCMs29cpfhodQkVOqMFK2bxRExLMqd5rd0rVe
Sy/XzcvUcxhuCykLkAwShPfHqyJj9L8te36Y4qKKoS04LsL7pBWJYIpPfnR5
H2+l01FKIGmRPMxYUlLr+zVF6nGjpIvjGaqmqoqXfBiJByUkhbzVucO7oIKz
Sii3jsC0ZPu6CXs+/QRYA9Plhq7fP7aW2QVb5b5JFl1T58QBDvNys6pyHwHb
6ea8SUfehhJLwkL9WvnSMpfjyA3AyLvGyrPGqH8dV1wTlYzTkHwZV8OPeoSE
dVNzJAaXR6S8LkKe6DF9YXKIHhnGJYUHHHApeynqq19gur6jP0Cb8ppRSH/5
yQHBZvXlmgxzF4Z/eVAtgbH6yb2+Y8mRzns/aiCmmRQL0wkS75PrqLmGEAOA
z6WpXyIxZ4/Iorqt8UpkYmiTja7mHjoG34IAyEPj5JrklvhJ+r4q3u+Avw0Q
Pisn31tIONsfJsr/k/5FFQDu/zQPLQSKM54lD1BCc/1EU5Na9Oy7kEsX/Zpq
jnvOEpP1RmXG2BmbK39tlPLLOn6ypMP3w2DVv4GEoRufaOD74uGokj+6suZA
YwaTqFeyvssEo1FEF9baUQFf41sjBz8MK8oOP5cTFTQGgipbrq95qfbdCO9B
GhOFbaUtDpQHiZhYoGG4Ef8XlVd9ggVeAEDcqkV2dTQ02khVUbV2zyM5QttF
xIwn+uGclCPNsRf8JJIBFchNv64KJAM7U3Mxw8MfAlu+DAAacidpJfkPEHRC
Pt1wIbljyDpTNIKAAsWhIZC8K/hgFybPkwGXbxJ4H7qP9zr87LekaO1KbB+j
Q29uxUd5TEYpoAWF0iGkOCprdEbkyUuMvdNN55em9tSPiCJSziDnQsgBBYZ+
wB+WXhyeKiiYyVWfahps6ziEtPz7lg5Ah0IRvuYQT/ehTQv4QbuvXnLgv03p
6sfkStr7rDB2YDvKPv6jZPOaPEhYHCOZAMtU8qsyMB7S8wcq9wZ+XoSyzdui
vg61h2c0TJCiZGM9HqMtil0+UFXwwp59jWW/63aQEtWrxZbFCzVi8u3yKQCS
0h7xpdUJs9CJyXh/NabOMxVk1m2JnFxPfHkfpnAAgWhlOYX1LIw6lekWKtYo
d3UpWW59+Okm52doY72rDncn3EJil2d7V20JdKpkVSiWLA0NwUnAbXUUZ+VZ
57+If68aoDWBlYk1FfpSK4TjRoTRWIk3gz++4RoKoVevlASm2bVEfar5XZDn
ZZ3XFDshQykzFjCGI52DgwOmkXQYsqyF8Z2M7OaGlscgDgjgfQtqccATb8xU
B+l+PfWdHpLOCzbTEI97TxFqm3YXHsq+Ixyw3pLO0JZiNQuYKSID0KD0xduk
HXNDVSJz97F9+ObtQnvQpn0xVOaNGOKNUXSrJ95m3WcKIS7WxWHvLc+8jqpf
kY+sxLkVSWdoLEm7uo6qvsYt1Gq6APK5owhdudpgSD4x29ycB5jXUiot8D/Q
EHkiwlgSF9mH4ofiYQNPCRvQQzJABtMYZ1wlMoYoznE4nUynVPjGRK73AspX
6ad9aI06J7ZmLx3tKUwtKs04Eghem3ACbdYp1dhcmST71rXDAax0lNFTSfG5
Y+GY4sPiCVM9sFr2gSG1r+6UmP29Tg6JsIlB/3OaFaYCiPtuPDMY/ALKodsY
Ip2q5xQw+omo4F3Q9B/51MSotfsm+ycpq49ozhU92YLGNNzrol6W+sX8mGkw
SbKhN3zVnO4CRfQLFQtGbNBtDUoLtsqr+QBFdwmFhcYfyWYk656GdGfz+HUW
HtRTpnTs/kcUTDC+o+y0peST+V+jYXJi0ty0MzDcDJxGZX/GAI2wTiH5oXNM
tNjxkCOkLcYpJyuciPqwY/Boyf5R0ADErPFMUsxn01a0SZtMxQEHeIm5QJrf
fLFeno4JPmYa0vGk/v68uxl7IOE0/v0gnW70vRmh9VWrmIty5FehM3wU8LPC
VAiR7ipe51WF6KYdcDV5Z9tbWTC9nx5l4eP7aUC+lO+fyK4fcwNVQ+c/CZrI
mU0AcP7a61fS/olvit1MdJja94fa8fXiD0GvGqZ9ZNX0D04pY26RycsJnWr9
G8f8bL7Ip0qpGkQOI60PWjUsITOhlyhV96ZqjfWKEDVs6J8R3D+e6H9gLxLN
A6lg9Ha5+E4g1E6DjiIdUpQ45dehCoKyCV/8CExp/o1QnZlECj6tPc8l7YsJ
5Z9lYnrvstZBdtV69blq/xTDcoxzp0RA4JndCiilABJQW3/BPtO+D5XZ5Dio
oZwUYymCaWrOFy2nnGgCy5e3mwWB5b/88Eki32GsNff7Cx7PcSWFC+TD9KzF
YALbG+TW3SRKfH9vOW3TcoZyIcPQSIbPySOaYMS7q5C+pI7eNZFaDAf3A/o1
lsjc74spOjgVH+jLNNiwl1lz7a6BdC0HwVnzj1tZ+yQ0vZ1tlI+2A/AqFK6Q
suhxxVNZ+/p9vqQnQq0T6Skcxs3M+iR+Qq/dZvQmuIX3jobTLntAgw5SiU5K
LIv7pLazpekmnC+ld5uCUJqwC5i5cre8qmmGsYBWmBTygDQCkBWSlieGHpFG
yPrCBexDWNphFMl+yiZ8C9pa61VtxNWeSrySNC0fSD3IegJHmqHV5vb78Sy1
wpKKb0I6O//EF4aH0Q1KoqEolSM+lNkgwUoTdvT9WEoLst5haMEPUJ/FSjBh
z3EvcT4FWPzvlFyxSR0ac1bLGz6vV+XPNcjDXMvjwyPFYPSq+Q79BchvRTFK
5MvWkkvIg2I1g8nVTGh6e3ORrNL135KIz4E8XUVWjnqRelaDNl5alePN9kpF
UMS73nJcENG8tbTOzUE1wMsfow0woswVATDvoUTh6uN7H4D3KXsnCukb61gU
zJN70c38VsJSFaRCE/r9dPWh+T38HAc9tpmKPKMFrOHMe59APg6KDagjDS13
VUxAn1tPkuc5gjG4cVhtWGJc49DZQbNBzv11dYLHd3vjg0E37L+/P5AHQtr0
MxtcFm4kuz+H7+ra3i/AmS6yJDi8gsCtZ+oH208tHxwHikXX16G1cWYoStUB
R8iUV0GyqzhrRFXQJA9GT4wgzcrWRseryj2lqumc4gWcEquexCY2oS9x4yO3
jx2kQ+iAn46Ho1BZGUGMOo+lZRs6Qb+55ZHymAagM/qWywxjOmNYGJRoAyXw
XPfsfx6nttMFaWIzcRebHka0xSXUYtdAV07GTd6JfW3YQHivDihrctemIEAG
jq8x1qU7BzZu8ATjmyKd+MQx0nia/bxpRaG3eiXwhElKbg2XnB6NbbayH/IU
BuWFwgnpLlgt/bdsjB5MqCdzPRSNqdSiRVW+CoQQ9Rin1CpIZJ2mjkNO9Ob8
0yQq0aW6NHpQw19tCLYb6tsfecOqDbTh/JP0bipShRGPvUJSMlY9QDPCNizR
2Z14Fi4JsUBUhgWcAc1V6YfOPmj4wyGK8ujCY3MTifG3UKKIMRgslqnrjYSv
ojOi5RzVOckSCej4nLvmJDFw2ZEiRHCh3QdcHiHZj0EegtdDkixi7mRzSn0u
eEC3syq4yiVMMDT/xJR47YlJuAQnU6QWcnfs7/SF8uzmnSX0xHo52HTOTQHH
tRDVsHoI8uX6myuzPaJ15ec6s2DZeYdlP4amqFrgER6zs6q84LClVouRliIy
phy9ROOEK3nk1BwdJeCNsThe7eCTq+f4mstHL+NYevIwwfZQzrx2XXkp12p2
xM0ZHjdsaxKKIb3AUC80K6paqiOF9Y3L1/I2+AM2SwVTJFEcvCYirq4kCtm8
ZlFhvnumE4jUGvLFrvnBnNUGqEV6qn1naqHpuNGbBrbi78pgm2o6SLLgGrwC
yWZVm0nWs5yAMZ+IGcfSL/cmH0wPQ+ZsxXFBu9QSIgcyon/AIvwcAxtusRHj
SYhmeaFwiFf6g0l2QitAWZNqUrqw9Dpe+t93VRxc1IClNGeLNRruoCpay41h
jjpeHNodh00LJl5c1baCUi8RzYeXzxDlNJ343ZzuKkw90UtTxrhYMBBhbnEs
BJOI9JJ4ZKI2bG8XcI9J++874afG6O63FQSrkrz0ZvBjjBBvF0prwLLhzjn+
EBgqh9Mvk/HDlK55FTP1nk2QIhxch2FTI1djYQt27BGxB11hhbWD7sO0EoLz
YHgaAXG+W9AWuR6Lp7kW3y4rQXaOB1lcC6xtxlUveTsjdySI8tepwf05D5L+
+kiQDLYuTQSq3Gtn8ZLpsHqrMeXg7gpE2cD0K1zztvXUpp8sL2UtqAt1p81R
LwXX/bXMybBMAPyrPpaCZAdXunzZWdV9Enfj5z/V9JQrEEJpSJnMg+PiEHA0
pmwRe/Jr+kFgE02gdfkzJ1hJWRnMxOIWXqdACDXK0fqK0WKr/JTUoYMOCKv5
P8LK0yi2L751J5ZITXzP6QP7WFPvS2EmZbrP1Nv+44+05fAJu45LT+gotDQU
GFzDjLE3C/Dg/Rp1IJDcsijSDJ3nRBScov9qLbzsliknhwWfqVc0yDlpoNlr
sw9eQ+2/slHBnSEijVbsavPmnHVnVkjh5xWig571yFJSc0dMk0WutPug2WHT
XZ/isNn1Sp4wzy/7r7DgOyLOHx132IXtta11oAC/aBKUhiUthEB0NKZ9ksU2
tfhvjD148WDO76a2HgOKWUMCiMcaMuwj7lAZdxINZ0/VMMy6NtM5k8RZQCSY
I35Hpx3XQExO81hSM1zZ5UOQGV2UIlFrGOY4QTbqupcMj7x5K6AFtQtEVV86
qyMX2+bLFtxBlEY6YyjsD0KxrjJzDHBDNhe7XBFRxZonJ23pUZiLlTkVszwh
Ct+sUC6Z8xk/sUrjwx2JttXNXpC1SG9nJS+wbN8Hiy1iXuROlelHry2ap5sO
Xfe/vmzcD/m/f8u3gnaeXHcjsyz2LV1uTAAUMVbAAyo73Llt3ECPIEvweFPc
YM9Ydsiio10BhNihB1ITIUwCT4RZuk6k9hOesbdzlYooXCma1VvhDvl7yeMQ
Grc7RE+5uMxlkyJH8mNaq9DdUHgD6RrX+ds8I7ONIwOO3BxuN1M9WDux0YG/
qMoq/thJAPEWWPUQbZwpLIPwuWSWnPoQh9WrH3w6E2Z4vqB52lMi2eMlK05+
n+4uiw2yzz1jIgv/8eaZN+p0G4TlCKsfdxXogGgxibGUSyLH6+P20kNgIMiT
FIaSBaTXOU6xElYNt3PWLJcP7pXxvP0K5sERrUmGBWghS9d4Ncpzxhv6Y1RU
hWUo9dXWzScoNrI5X2bz/YUhYaLtr4Wvvp7a2xI4d/VA5TQzQ9XcAFmc6KIb
qtJtxkL1I9dxR0Gv/5leAiwvfXrRkEiOsVrVrBZ9fd2RDsLAEL9c9mVTK6Y+
64DmpXjqeNDEIEY0jF989hI5FL61PGEmoHoWokcbxXWH99RnOcilS2VKPGTW
ZCk9JTXqtcgmNEflz387madtibto7wdvyP3IHmKp2da8jaGY1anTtqvVXQ2d
PnbymQU6Iznf/tQxwUEuSMIRhQU3kuGcZUBrHDrhkMlcpKHU2zHJdX24ZpWj
OR+Q9yrG5STx6QBln+G9NGTyuVjLKCB9Efv2JhEGM3O2MqAodJWHL7kYX30+
fDGSE9Iv5QwG01U2Hk8+ukSJBZpDN1Z5Qz/pL6cAnBiGqeJZxWPqGKrw/1RB
25LmWEnZLCaacEY0vjPV8tBSJ1GLRH32xqpSrM/Ugzrfvfolg2UQFecHfeDz
1YDu2hTDlIUgA0k7lvSOGU72jHYtJkODKcmJ/wUIkkRKjvQ8aSJQ9ug16buf
GpFs+WYkP8W54RFhAgER8xVtiM9O3x/5ClF0dYvyd9FXzVPmaM3P74jLLKzy
vpDzQDLABe0ViVrZI3gYnt96S21d67s9v2LYY7HSNFqagOmbrnv6i6AEGWBt
IaX7gPkMTnpIRqxPG/Ty04zM1SP4iO1ne7IwJ7GEi4/KWAvv4fm2sTxFXmHY
56l/9TuOnV1H9mXR/iJ83Ft4Y/wXUJJWw8oZCe+DgPblEIoiQJ1WP7UEO9yK
QkBbVNSBQULABIh2lppZ+Abx1ZPMnfPv4ns5A1FLvUOvtiQ6JvT6jMKveM+6
ogrUQ2iAFIFBrnE2UHI52HZieggBDvE0skMn4ndY1t3MYaB/Rbw/ME/9GloL
CnlEEYa9I12KHxVW2t/Ed1aEmP7RGHw3MTzNvlD7ZsYO34GdP0ZDyhplg1MI
TowGC1YnDFg5Ew6/pL5szHO4sn7RuCoK4hK5eOpNjYp7kvUWKPE3udlnrO4Y
xuT6amDWEmjyuL9WeZr/b41Tz9UKr5BfwSixSNdGQ+xhcM6TG/J9ayCG8WSb
qM8KzxTzb4eApS6ijgD+Ou2CaEECquIIew4IkmR33L51Aaxi+q0h4duafsFt
VUiwo2OHhH0+AetJHDWP4qIrYAn9fm1igxgthzlxSt6qroPomGl8ZVJd0L12
SrKRHl30Hg3cs6o90qS6Pb0rewEyKumjJAKI8VR7UZELpEU8NzHZVJH6G/TX
U2U9ZwNuBrWQlLBkG7kJU4NLjHyJgyKS7z3sFF5h7rht2a2N47yHM9NrigHa
nxKpGfMRSpmDnpCLchOTK1nHN1UBqtqRlwUa7AbOj1IxBNOdzZshs/3AW5rX
LvGWcFdBKIKNMpQB0oMUbVu7AiEQFMmKMV45hs2C2sZWZDoj4Cm/f/IGaIkk
9OoJ/QVXVM58agiMYbEVsYhcN2mDLUyUML9M600Nt25sDuHwknwCPlspf5vA
HmkE56mJAfr3dMnobC4FT6li0zTBXQ2i4RPOQd4XXdswagJeyRig2CjRXy6o
YyPr2VaOmWJl78gAxozdHeZPlviYGQ6o2NF8XxVQKQSgBYWOZmNF8Aduouzy
gV0GO5xnk1E1gj4MU9AE1NIhufKcGQfmonIlCceFZ/6+guOHK5E+uPQHKvyS
wVsEUhRw0f/Us89cdU54vbOSHhMdh1Cxn5t6vY6RP6nM3x3xucV29TXZB2aI
U5XyLbEsGVmq/jdMli8wcTjUAXXFPJLlMD0kxN++7W6s8ZyXj2FZVn8XC+tw
NgalONc88pbXFUOZlQ+vP94yIRtQlQhy1qsaDPHrdiaTenpIQdEW9mLCnewD
r/K9Fk19QnKrM9UXQFHTbqK5eOSpOKBuIacLN0ziGX4echrn8LRcmBcDuC7f
qE/bgdcOGKtHgz9KsuL5SPbZoXOvT/pqYVGPWpO+RBx6LYHFFBuUjShXHF4P
kex0OwW0lTeYzew7miEEcOE40qfm6pm5KzRNNGBNZ2ergzMiTk1MynrIWXJt
ZIvYzzHFIOpZZI8oP1B/vwlLV1qaIQnhKcWjlTQOazfCJzY+VkaptuMSpTm8
0eqNcCrJfBL5il+fhqLLM5v75Rtzw9VrKRDz9lMG6Mou3SeC+a4eYHtbd5SJ
PPq+bvro7SarU3y3j9Aow+evgUk6XzoYCCfjKOPfFv62QhVg2L2OXt9cajit
ByndpEEgDf0JCsqdCwc3cAigWZmeADw/DFlCehMNAiqu7CeuiYDfuhGwS2tz
tzaXBxSbssDoQsQ4nxqS20t4HQobHW0tGfkpQYJ3GJBE0SldKf7o7/AJO8k6
zVhp2LPvGEysfv8HfkxpBj41ukLQkIIULXQJEksgDrY1cLZiI1u8bKWVpAAo
PbxkiIvfbAVUtpVJSXlLQ0pRfEKAMjnZK1/BkLMF5GXybcA/Nid2X5YElN2+
u7e29aQJWe8otpdXy7ESMKo1KA/yYxX6iOHY4QjrgzT9hqOmIHKEdKdyLfS3
8846P7wsXljQDBkzoSFK0iyUt2MgI2CE1hDTYtlqSHXa1R1IzFQsXF0q6DLo
hRDyi1jebyk9MSuU8UqbOKzEw1yWpebnJwLRVhhvHWCbtUCj5bVQqHWfQkBm
OWi6yUTtpUdp8bCic5qFfsBlN2tmy+/ySPtG8nFWxk4h4QeTJfK6sOq+8889
Zy4zhP3YEt9MK3wuEUdlzCIEFwUv95KuxZeNaSW5m2CC8Dlw0NYTzU6IgFmu
kpDX3ZR9YILX8oJoqj2TDiIW/Xv/eu8SpBVEscnSIdvwj4v2ZR48cMAO/voq
NNoI/VAaW7uXVBpkOhMf+9KXD8a4qQFy/hBQ8QqW5QmnNkR1yvnPZG6opM4Y
at60F/t4UTc/X9PFEHOQJZnbrugYr9ScuANFp5HPb/bfChwCpynyNPYUMTSJ
OAwEmFEwxD/+fEb7au2UdtATyI9jTFuHOdyG0Y/xH92wzBIuMhpApejc6Gkn
Kqfh0MdrbVcXFFjuCT9rMxccXGMjpmZT28nYA6xVb/z+IqfR9mAyiIY4YV8u
lz+mlK2rWDrgJszuZwwL7xVi+E6DdVIztIdaxDYR6keFCm4s3kJhdjSMuRBw
SN2FNLENs1dg/Wuued6/hAcZAz2DEFA4bIzqtjtkIl6ImwrOY5YQbPifE+8j
gGMs2fz9XZdn7vtwGUwsYU6x4xT3SkvDOE1cv4Xyi+P6BKtGqUJW4bf9puSo
MJKseX9KZ6Rlfd+Py5+5UfhJ8K9LsCN90ztI6CMLRO2yU6iuD1ma1uXPyoGT
q9fAHd4EKKVFWGtU6msKU9Yz2vZUWJ+Vo/yywQYywyDSYKHg0dlCXMaS6kGm
IIBa2x712YKYVQm9qJtzFuDRTyk4cAhEIMiUz4cqAaTXwcImBrhs3TE3D7Bk
Ea2Ywd4qwkYRjLrb/E9opQ8E9wGidMdX9pe8HSiLguVPKWKjpdvjYbReWXw6
CMRlu60RhtRR2zPgO7oPTM3BC4r/V9nbad4mHkg1ZZUq5KaGQWa7RYi7ENKc
ucolGu/U8E+Ld3NwO5AwlBr6i9QHw73uYxONbRNB/JxZuqW0FwH9lNXZHYxb
H0amgg3QphI+LqIAA9kFPcvd3Pcwod94N2JizarAsWlbPIEsV+Mw+x0Iqzc5
4+NKA8bOnVJ00Yz6MjRxIt0eyfT9LZb0lsU75mWAmp9gNdXJRHMuR1gD2z9X
n14ZgqEuGTZARU+5ScYF8KEE1d2DLX2DcTJzY+dnrm2y1mgNrX8K4HPbbEfB
xEsaOddecJfJ+U3wD90hqY2PbsUraNY1YeUT5pv0KNO84fjdaNjGI7iEmiIX
gjP9Mfq/xLAAg7qC/AJySvEIJ1/ip1NR+k7qsc2mD12ERx4/jJ4deHe2mauj
1YWgVBH6bUSB/goLINKVl+X1skIIw5bwd8Lsp1Bo6lfSeUbQhZR8gHrMva5l
VZh9QFALi6euxhTM6WmVdaUjzOhBBXkleor6WSKMCOpaAIHFo0eWisu7YFRZ
rEK9xxMsBvociCK9LykE6slfm/HKBDDFU1HjaYp3kyGdlRE3RrxeP1S8USkd
9hXgZ6G+q63XdHdgPgY6tcdJdPcudrpktnGwDdL6jyyYFAmPkjirssLoVzzS
T5S+Zm+exAW/4Vb+lqyyRLu1+Ica6MASRYffjg44n40wzQEksAbe4QcC3tBT
D5cWdbyhDiqpL1O9/jhFkWaqQy8SYWjvGPE5CYEW6u95+XYl9A2wWGnlSOHy
GdqcaUdFxw93oif77eHQMWuFpC3lWldlbaMYA2XE2a77wlJY+AEKIloldsP9
wMAREjuGk80G7B2MDyeQgZtf3GCXEMJcEW5UmFLIkrv7vvQNLW/Q3biKCVil
Q2l+t2DWHBfZsmhVJYg9zZrHTKVIrNIFYeSDOCyky5onlfSm3aORUqyHLeOo
HqMALl1b/zOCGTBVgaEV17BPfOQ0QGb4+RLLjpRiqpLoMZlif4j2zt8e81q1
H0oaCBBqYMw+XfZH2efV2QMuCzMFGTLPxKzwGSmpCsLo1s+AO5UDgfIvVg9q
dB8QYt05MiLWhPy0ex57IF/qUxKzfoTWrEl0zUXm1Zy2VeyP0O9m0dasB0Mf
FenmM18aYh14xtA8bNY9tx0nooPabHdpNV0FThmnNhxPDzjrOuJqyv5dq36H
QIdIyulG1E74uIDvhyDVi+KIVyngUQi+ojfc2h2R3mu+U855nMWqGhLL1pS8
Ad7jW4TTHYXpxlLyGBkq5pIeNNZYllb/eo4ZhakUeZ5imY1Ql9yExTO7o92m
bWFKPeFBPRfqyYoSKxdNZDmt9OyKWadPmtptUfkITYuIztQ0MvKGUOv+Gdok
LY7J2QMoNRCebfAaBFj76DoKsUmWFsN6V9Rmm32JZqB80cloBOW92ueTiJbv
F4R+yChkKc0ul2FmCOjSLcfu30eV8Osmqn54gEK1/c8Ylhimhy9hhlREq0QD
8rMYvMLMBIt3BnXGfOXyGdbDa2Adye1aDgGE9EgTdzIeMmM/kKNxvYlou6L5
bVQ45mCjC4cmnxGJ2F2eUV9D2AAFHbR82VJBeGgcmpTiUhoaU8c633A3pl9J
FNIRgUnE2RZErsF4bp08mKeDFnVAvGJM3b++pQYMIV1/4Bew2DRe+BLHAccD
y1f3cuRgXNj5gpRWajUDrCsyY3CGqVaK/OMF25/Mger1x2M96rdF0hdeFRMm
UxepG2lfvLj2hmiIfWAV94X2/U/uhmT4i0NxYoEF48Uz+KEIlH1drnnN/JKa
QLbhmIBgfj9UgdlGMoLQR2R9DEpvdRGpS6Vp+1A/WS/Ww7+c36tWIGJ7dzv9
kCsDTTq6+wsrDai3hH+rq3aFVvwDC1jeulep/Fu2d/HBM3wyabfkUcm8Dv8o
1fG9rpPkMpAgrvt8GsVGRU+BjQFYbMKjFfy1eyHa5k9ySGrqAd2wupcdTX0J
u/OjEOVZA6fKy3qZPh9G+VdgOoDtUw6U6CdZj6PDhc1hMK7Iv18fUVOWDaFk
V7ecTnI9NY1SFgy6g32Gwnbp+ageuFnHVsO53aP9gP47Guul4Fih+x0oATdd
s9FRum/WY1fYCAa3Yo8szrHGO7996qoapjNy/m9ZY9QJxbEnmS7JNf6caVhU
4NDKPqy3X9onJAUp1mMRcy3Vvx0WvmBGRRCmsjtgSa5BLYp1WgeCfNtDMQrA
Ehj5jTUE9ePClr8CKPw3fKvWKWBN8BNlLKIkiTBD5RXSC27ASOnZvtD//NKB
Yxm9BMOD2kZo/R5I1AaDpaz/RX/jJzZvkS3ODv8PEPqRQzgiLbg1LeXezh1u
ktdS9nQZHlvoPHk25Bcj8qmo7vilqmjz0Z5zAjA9+dspt0ZrSQ6rc6zeTpmg
C3eB52BULsdd8hOmRtHCBv18g33bbo7mfvMj0dGd/zEXC8qoi14dj161eSJS
pP4yVxODX12DcAVF5oK5e7t0JTr6ACEKCLVECDkl+CW5V+ARd85xEp8XHrPy
ysxena400Mz8tS2/vT1KzSqRXFy1rbVikBwCrxCV3uMcuiQbQbF/WGSe51KW
EHfTRn8/6qfp10E7EqDUXCCTSowQaMscsX8I1/FEnFIk5zc29qBcdfCKe7Ho
dcV00l4UUQyIjJouLx0nuX9l7Z3ewYVYzfLNMzmlb7h7144JjOMuaLabCuOK
FIzXjUSb7VUw5x9vrjBrKXZMjlm2F6ENKNERik32NeUTxbPr+hJWq+29xj+P
GV9SofbJIPkTaSaJ+A1DNVRh3ll99nOWY7wtfoj3yb1N1ChEJhk5jAWWP3zz
FGDwKEFOhcsaSRJACwo/OmPmNctsMww2yRUz+Z4xyh3jNmZR2TNFmr6nA/Zz
/2PymWGI5cxXB/pR1nnQQI2/ae0Pp7z9sdkwr1uyNhlc1RttBwJPkioWY0n5
46HLqoWd9lYhhPzxIHQsXzNZB3ahWdOr45cxXnSDff4ILPL+HVSfcjBYkhpV
GzK3aNlocvoKGjX5LxxgMTq30S2oWU12JXlmdyOrSdLr+T2fHnU6sHULNXyC
gKfEC96nX9SOoqNNaVz5JpdNQWQYsfLArjpKK3wqmQG8hl8gN9hacLJOcEOi
FaVH+Rl/lIHubwQaoi6pmzWJw33Cio1vcWxU9GQR1CFwrk3HFN7PL8RUIhC6
q2GgVYiyzxNBaOIP7TQMuCRMxE5+q6De4mCKyLWiTC18ecrjeh5L2g1VIC6t
zlc90A1HFEEK75wo0H/hDaPnRvqU7R02v3tkc+OVIkHHNWKbhaMvFuaxrDqw
WNEexnGdbABwhh6BH5FBMbpefcha8hb3qruAl3Z7LiDrNndiF+saJMpRLFHE
KzPp/yj9pShJvspUA29er7LvyD17+mTdRZGoTahTPGK1aMQx25/drW2TbfqQ
EBiV83RnwPMH/OOIL81PGZGrLdIesBzdH3eXlSG1jC1IvGNm7ZomnJQ6043R
QjB+HCFjkKr+Q+z9ivt478a7LpKO5wXhoCio6dPXhIp6/LJQDfDwlV1UZelb
dMGh71DvAtGWSjZ3Yv0xSN1IOM93ReYEucpJK25FdCe3fBNTjttV8gXsbgW7
9BIuXURWXM6TAg4MMWP0Z4oXvqEBVjpPEQjz6R9X2TAkutrUC2j5hzyNvsO1
yOjBfNnBuoI9z3qNu520aGdaWtELvy0OIXYsPCAdypX0vIcnaQtXjpXV5wmX
c5aenM3OY+BYu6UMmznIDTsBITQRxdD6BG5yVayhmKE/8fWv4zdZMAF81PAH
X8z6Jdqo8TOCVz4S7ewlADJ9Y9YMvbrvHxi/j3r1CReEcSij7glwBX3V+fE0
koFcbfAL7xlYHke8Wwl/52AEBDfdviQG03Z9Qpt0Wr9/Yz9DxOxegu5GjhbA
9LJDTs5ELkaTjWWo/+sYXIAg6iMdDdFLJJadkLQsALxHbwMZVC0yd+SRfSes
IwjORfkVOjlC3jOLsejyHonMUo4ZaShMLs+uGC6QU1RR3FV4RNaRSFoyhDh0
/t4iPLjj8x1vogPOqmaRUNXJW/JYm3c0tNj2vE5OyVTezBuGxn7E9sed85J7
wEw9qWbUqVBh3UIuqTstuw07D151ndwUGZBy09xhUMn+V3P8D6sTDsomkk0F
eJqAhAOVY7mC3p5cEM0MAhrSt0C0Vm08N162orKbM3n2wNw1q3NGDnrNat9X
iD2EIFELWzuUflo3sEYqpLgSnWbRhUSiyycwlQHmiU6Jjs1z93n4r7Re0iBz
7N5RRLomGEjGtCtmHQRFZLOXaFkWO2ecOG6P1cBF2tupJgaGMUu5AlaeHVsk
Ksi1jamtjTKilXYQngfGltcISaFEDiXOXzaNwmg2BNUWDuDkVuZsmf4aKzE9
k2ttG1xD9uNTxJ+9Hoimibc5xHLbs5jdYJFD7rP0FZa1u83T8xg5ePnjBzCj
bMdPdNWrWH/3MARtvTo1NUlnz69FBRF60ziS+cI4l0Tl6bHL1+nj3djg5+lG
JLGlCoKtfDEuReq/Z4jg7qPj5muIWK4V4MVf+sI4DFLwXdubl2O74Oh/48Mo
eAGuace3hzpuE/Nfv5ZhH/V7XpS1zQGr0av03JPlicz8gvQcbjDEwbq2ueZD
QRi3+kqIujy1LKLt5I1yAHmcqSKQRQLJLGttRaYrrNTzN4s1fzxO9Ye2h2da
OZcoS1F5b3UraZ4oJ0r77p9ttm5dWVqX+QW+jwu4mPNG1Sqn719xoVdP/a55
ALB+3kYvT30cS/P50axooU4jyEbgUDbAv0HE/JDVTlCk6gOTu1NN6kMun0DP
pjv1h9+7MqccUjrEY6tbgb2bkQOcX6FDILw+fa+Su7Aq+GIYYiPLbixlBX+i
VdRQqAOOAlKNl+/qbgYYXoH9yyzOhldNXHmNEEInKI03dOzRgB1aIVIOAKwf
/baA9cX1X+5ZaBwlJExen1Xz1iX/UyE3YR1yz2sMX35jg0q9rvd3EjVm2plX
zgaaS0IZlbXBTPMSSSV8GbGWa4yNTUS+P8YXGZJz6f2D5p+upf60ZKqFQa3N
tA9zTgPw24lvUSu+CK1iCZ2nmh77PO9xkmk4LukKyawYvKZQcp+sMI+ZjHzS
N6RE0hNO19Pk0t+t5Yl4aRkIPnXGmJf6fmnuH4IdtEGbv2fzPtfrBn4+RV+x
ynDm5P+m1yEoUMH0JP+UEjJZ80HKqH9uEkn3h5HfoOmtfi5/cvLLzq/kxMkl
/K3x4jb9NkB+snbk2a0zxdAbxaiTnn2cG/j0H7a6CzTHMIhsf4TNYWqOSP9h
/vxcCWjQ9lxFFQga+SClhvY34j5NCEgYBxK8BG1ggW8KMB0jrCTv+VMoRZki
ATnC4tP9CW4uyYWas8nBUnID/h6zPiyGQopveJjZGQcimT7CT2kOi7WOVF5t
vrsfxBgyflGS7I7qPWXI5qC+sQRW1VsvCprFgOgGFTBKItMDh4oDoDsWnz4N
gAsZPr0SEFHlDp8hu3uQvb0koJLzYBlYJCzgJ9PubtlAjVaIMM8ClFVI4i6l
994NIe8r8QANbhLbeZYLVe+URCR3qM503K5vHhJtALDVybciU5Q29QecRHSz
aYNyHaApz8TJ/xwM1Q+mXIvY2WNiEtmz0+gOIklQCANuFSAY4U913ta/amRC
t+4963h6wvjZg5FWOtLyj9jBafh5ttA7Z7oPjsXsPVdbQaqk+k+1eVBHr/TV
mwo7lNacWwrJ3bS30Q27ijNJ9Sel1cMktShzN+c5NNEhYEs5i5vZH3FV2aXQ
WJF6xaOhUCueAkD4E6fnY/BdbiMvLDzyJBjOgblVuFmtpWqquCvLuA//YZP8
LlMzFbaT46iGJI9MWvyhsnTzuqDYHVYH5MJ9xYtTwcAv/QNJYWkv/YJcHLyu
mxzcXGbvWRW7cwd27iNyFTnMpZWXivArVkjLJOzEJaUMrPbc88j2V0y5cnT1
yW1qIqysqdaGsTECLkob7UfWzdHzT5E/xYZ6lRlGi8/Lh5Yt4SA/WS+z6SLD
zvVMIH7NQkyCUjmSEF/yBuagzou4VXVaLQ1Zv71YNC0DV6KR5ocU3d8B8pcV
/fbWh+OPfHF7WE6rFWzb1V7HDfe8OygwwIk3o3KKIefMDYD1m6FFvgkIqrsa
NszSRxdUPK7pOasXqgQwhvzzS3w9IzF7C3+jOzrgY8OlCN7km51i3eMpIq/4
WLxrs8Ft80pYuzA7/Ra0lDrhQNcoYfyIf1GDp8CzWy9WPvPYg5urlxpnHyYf
4pb2iVfmSVbQXKemNrT8qx9nouot806DHrzZfQ0b61ShTlGqfsIGT2G/R9fk
0TY1/3q1nI1820O2WlboG81eFpjCAIJkYLPOFgKr1hVOihI0eX3wfkGuceut
5ew0mZN3jw7DXDM2COB6z572+jipInaRl3OcrcaVX/+vAhpbh9HuQO+p8atQ
mb3KcMpNfyDBNu3v9RtZk4WqQfrvfEXvRd5QzcuWxm0iOlUsdgI0FFzmQqpr
naHs3VUhE2ZrAuvb5jfDQJryF5LlrhJimScTA5ySmIj7Gu2CCY/DcWA14er7
l2yUiKvxD8v7BGYlXg9jrNkCXXZ68BBHS8Tcdtvdc4npEC3OUvRmXb+HSJhg
+bFMpjC0e2W9pYljpvu9DN0eR5+p+gxxeVCjtEcJn6y9l49mMYzVVeH95uSw
0AP6Q8MKFR4MK53mLF+0d8pbccpXQVGp8q8mWCHkbfx9YTjW1+37Q3qtXa7M
NH4LgfiS8gBLUVf1AeR2Y5517jKzBFpNdpdPHQO/whMTXAZmplt1OEL4/wOv
6MBNi1Ec7x09WQ1d2Gxn8tmhRRh3cBbjfpHxcxQRka10gDCL3HWLLqCP8lwn
eZd07qfG8gIJ9+wXUJguRooNdLliVsQgr3YpgGZaC2Vej05MwFOhaVtFvWLj
AmqGwPnAPOo06PsWP3b3T0KMzotgQnRc1X7YFAG/U6M3ckLHd9Ay8ylzsqc/
i1ZpguuqeD8XAay4h2FOm/SHPPpLtX3b8+sWaVRZZNlBkJNtGcKij17uPbI1
wRfzKTSQUtAVD1t9TkLuQ1l9BQaIJhehKy65CFcEcomnP5/rBIkRVKe5vcJ/
AGPT55BT36lIiSonr1pTo93GelvH923dNwjT/ReNH81WmSFj+Dm+xFiLhAdd
bbIrg9UFIA/iC5t2HQSS0l49J3Evk51btDMPpPDlyxMUzWpHBKPK4mMfPQS/
5MbWBSMDWa1quaAIMersMMWuvl/iBXGZdydw2m/PiB63hETHwu24PrJ6yXDO
1DpxaVvbHlWzvlBi0lBiUa3nEb+K07znC3oJj4s5gGcMfXrHseBrHM1KpxBN
ZNafvcBgHykFnSBaEQJf7j40rk/ItE/YxvJSv5m5rTw/K2iABT8JoFJzv9zV
68EuUYzz8tw2tKAycVeZC+LFuJMcpPLzBMASkYx6LgJ1oOqFgsjY4IbD1GZB
3BtgW+aRTkFsxcaie4y21dRd32gCqmU6aN7JWsHPW+jLWwAnjgbetuSsDMZL
olEs2q6ibpA09ciAV/Wwh6dATfaxTpZuAWIqSWhgaLYF696l8nIvMDogefub
1gPGeSYgv0PUhL6tjM+BxIf7vo4OzZlJTV4ZUnHHemE3R8fcT3r7KmC4PGij
p++nUg273t2RI002YkQKAuY+CwCQCsqC+/9Yk9b99T0bibv79fR+VURkb+Ni
9QcI7Sxjf/6J0s9VFV+qpXmW7eVH8Zz3Szc3grTCvTFndTjtKK3VRmD0zDzQ
dMQXN8GE+X4/rbAGPU7QlZw/fTVn2po3Z0rr/zPRHtgZaK28/GdH7kTWfOBP
L0nkinrVzqP9dV/LrVEUwdnACq+w7I17S8jFXWqC7XTuRlc4ni/RxjQgsxwp
mAOuJfBMethfU6BmfqECzyf5pSLczju5RHrlG+tizxZXinLuGPwI4te7KIQX
0naBEKOgWJzreo1ig/i+7CVsjnsqmrt2Z6YL7BTNTZP7fnfwcQ/DCBk/SdKI
9vDWyqVkh2GkD6uCJMMnA0bIuVNGvCjD7lLEgYXpVh4BEEoxnYvgvvfb4Cxc
3NT1i9WtsgcNrlpy4rOkm8v+GOGiS1+clMMnkxFjwrL7zX5uA+YDMw2qCZEb
VwpmZvKv+jp/pWUwkob7EMAsx9ogdYse20cDkEbtB0oH0oZ+flev4jHuKxyH
eCvmjDjR1nSjIxCQ07vV+EDu//JFuR4kdjbYcYR23mdiuUsbRui5ZOTbzB7X
3CcqJ43sIgonPOq274814DScLbarFOBKG9uTA+DHfSAxTDuG0BGM+FJd1Z1X
8VlPLi/3ffNQ4eF7pKw9QZvzyi70TG1+2I4eU3xem/+72S0r5cIWXQj/WN+d
5/kXnrojMBPSHbh4j95R2766C4ro+kEiC/r7BvaaFd15U06Ec4K9RTI6Ulcm
pgHuAyzJlbawgtbreW96OPJ0ZNH0l1M0uIp9YvcjGikcoRH6cjRtV3I44366
B4UpDp43upoyo8GRx5PF3GxZJuxmePq9zN+x+/PuTU1R8j14I5T9s0ECtTim
B7YeG1331LE6xH0ORUOkIRE7heumE0ZKG4wGANLBoeDH6H2+lrI6na78mQFF
6CrE+91rwPJBp1Oa7bqYrNmhD7LFcvvcoMG9ZLel0lVuqPiC9C8Hds/zS3wG
fgsiuQZ/1stjVQ4FNyKgV+r6lPc6/JVNpYN60WcW+fWa+gp4vanqUDQftD8L
9bkf5pZ80LcPN8iHeNnmHVd1ziSrvmSzNyHDn2OZYMmKyJ0zr8w14mCrnj3Y
y8mTwAhLbPQAsFGQ5M2zr++XIqamNiclWY9CbXUWIxAe5/Giq383j7Mvqjd5
tRHawcdujri5OqFAGOMwYMApOpl+pmcLI5r1liD1Uib+hIRUPxTNzGNciEac
KFsPOE7G2uQuLzqcEbo9QrLPqLQ2LqtN8G1aSwYmg6yMF7kNiLP5Ih3uxVlM
+JhMBDd5uzStg77QlmQ1PMNgf53+CuYvj2yW+b1nTLq7F9W8+VRU/WI8Lv9K
zo5I3YQpqrXmWxwysT7wLQPylxdc624icqJnbinbByeiYRy7WIiOsCbiSJrL
MkPH7WwK3HQ1UTLGJWNxMNnsJyJO3iSudWlpsRtLHMjha/5Vi3NZMF8nBnuX
jRn2rVwHUZr0VoPRPSBB+6VuekMvfPuf46ffhRgj+bsuI+fLp8KgaYPZmP1P
R1mhFlpeMp+DI0vxChekQREo+N2sjOZadHmpx7pVcUhIz9Gs2ynUCFwitPRG
508rdNrITvukvhtYkXFosDleswCvHlKo2Qz/Ri47Pu1jact5hJNAGjcwX6TW
hWdXy8Pu1fxf0lkzNM/xxaoUGVH957a1ccyvNRDyk9/7YtMbYW9jC7bfbhSR
brRH/3spmIJZf0XDvVF3ewryyNY90CRoKgDl0XAcndHT9oTrabWSTdg2BWhU
TRttxL5uvv+muO43P78LIVe9XCg2DqNooNGSlVhL/Wzu0wCaKdDBTv39n6Ze
B0nWVsBhQQ2ZLzROwFPYAONwJGF0RHfdaWRzF+63iZLkkl56SYMi55WJwCan
mkWdhTUImUykHat9OLm/58Nu24mNlitVXwSDiLGqWJSwi6Zip5libwwQK6oC
oCrvUcqaWPfnEEc/19vQvui/VFFycnhDJj7ckyzI/rOxhzX/8ubix2hCu8co
pe9K4pyBh6ysAdTM+y3yYXKGdd9ca8gCeC9bPi2HUkVZJv063WYmnV8en1zp
elpAwrj48M5Q2olDmv1pK2sxDBlDZoAg2PDimxfIJ0OVjfgrGYr/8+RWueja
rF3loQ/3waLagPdnmJ4iJ6K6Jk8+DhY9T/8z+X4a/HQJer+Y+xcXk91U5TXe
6MBMYlTQIZU5NID+2mxkplCLE+I+SNe0x0a/IrIy4hlV/qdCW0UPtHFcKu4L
Qqk6O2trs1um5yIbT0kLQ3LyhWUrBpjBjOkAsFX9Fa9hYPSOiXcmXr/JgMZ0
Oh+urk2D3G+f8Sks0mdlU+9HFHnfQKzhVg4j8JB3jUZCcvdZl0zzzU2kYbpr
15PVVFIlAxSGXzG1zzbv7JVXzZ6RjFLBucF5IkbwsLO2RsXqEmYQdpvk5a4f
GjLAa69UDRVYm36Gj3AxYFqx88poBtQz6l1WdVtfDe+quuCys8iv6Px2Lfeb
ffNtgMeLn5bYltxpzbrSxjwNZmSvVlgOIL+t49+QKSVLh5C66SGttI7N4vFY
kBGisq0d4aU4KGYmDJhh7s3WfT3T+zSzuTpEvydY9nDRQkg5szfVN+UQEWqG
VLDlyR5peMqaH0KkGTySb88j5cqzJ8jzQK0lUep57TGQfWyDGO5QMrEfvAMM
KHkTaKwqbIjOTj9h8hrWZ/kf4fcas1oSrdgqA7JN+7Um07s68qdY+baSL4eg
KOO4DlQ5QC1XFqKk6s0i+njHD5sTmrSyB4f7yQG5uyah2JsKjYvU6CVVGHbh
XqSXyej6+p4L6J7phgacHQihislprg+exz5jwQsiep4UGUX124tfssLBgIP2
mdvsRbAvBaNkRzB8l3plynSS20gS4H4LXzVjC1MTriXPCBAxPV9ERDZm7Ynl
ycGGNNYpPxVeH9kMBdTQy61VTFQaoUAEKHidjuXN9RUiMV1WiPN8PRRfUzxx
ACz+qTHWLwdPSyeJ4AS+Yq09NX0/UotXasnPA/vHyOhiVZrxCcrZOQ/EDbZd
KTeuWydntG9IOboG+QVm+g2+K/d0dXXE0qpgfoyKekXRRqn1zJb8H2vjxLS8
qj8b4V1Ojosmhohx0Pe6rf6M382GF9kdZrXp2u2VDEpDvWG/yrqhxhBDLeRg
D2IPz3eqG2bZTYJ7kk4aVis1DX2l30HlUNy9o6ObngPSjZ/jg7ytC+L4OBoc
/WwYqotgWc2t3I64g7sa4ZJBQxW3IExkcbh31yy5ZHHXqnBZcfNpFNxOy0fO
vBr7+8QsSPGXxexp8aV5kptenCAyxBZJGfQzS9CKIw1GTPqwupw50FOsnfWR
1VZrFrXCe/vYSbSlmz3eC+5idRWDJkOLAxtX1FxFUYY8gDJsMokzkd8UarFf
7YOVbjpi81mCdF0grVIxxMNZHmbtg4blUQDMAM668ItUS16rovzuzNi8+6cv
21brTcXWn3VOEVJkt8ygNMMxIx37782RTJ7iK9ycoEGUrwXy374J+FbHGZOg
PYfU36hcZ8kuw89dhKVxvpazEciyipO+g38HY2T3HnVOENwPrNWMnD6I901R
kin7KBbSifPnUTQTcH6hEdSgdASnIOhMitja4EzyAlFpa4m0Z4eDtBnFmakI
u5Jh4GBntqg05T0t9WFVFNmoB/JoqpvOPTkmhuVpLpDNahLv834IlGxQgBJZ
Ea0d3tPgyKm8FFj5sZs+XOdAaj94RWGnwSvUoFPatq6ICCyLI0N5JzH/gNML
1y7IWEIk1DgAUJRQ44LFUUSAB38nuW6EAL7yVKFppgffff+V5sRR0N4Vhl1x
orruxzFOwdRRegx+oCjgdL3DLo08D9M1lPpykMcYDEz1oLJT/9biHgU5WOV0
R47NSqjqUxghk34rVilPnK01sAI1VOs9h4gZ75pG0eEogjQSKStkA+ja5cVP
N2f4lc27jsWqNSxbSBfraIObCunBYrT4/NWlFvY7upjlfVYSs+RqODn8x/WY
kBg4wnSkAtsA7mjov+JqQYcfWOQJi6eTVTVP8PdLUyUVbN8qmawcCDwhCgxT
6wYRY1K/gpAz5+xa4yW3lT2GzlE64R2Ifhn5ZGF1msHXg8HmDV5oh/AK9N3e
oXitqfFJfFAdCGdfu1xuCcC/7R1DhSEmptJKrTo1Xxt2E6WiR4NFDA6KbwzJ
ZPYeCuTnD4F8IWQwG/Nd+BlvXY46m//thYKD1/J6UrbidMELWzgRTWDhDvML
i7s2vrR6pfnRvHu3zt3pBqmO3cyOYDfNk39Hx8X8BhTmpejb3MsAEBN01nXg
cBTT+hFBDaQGGa3Vwni1OewibsJkjMe1d3FDATS1DIKSABgYFAs6pfjV9dYs
INuGmVGtnG7YTF5ZxhccLJO2v5wxYK+yFEwegd7UvLzVzH4K3AWv0nC8c54b
vPMOb1yi52TCWaDCNzpBfbe/bnL45+0clOLK8CPZfEt2EavLlmm9cxVwV/uY
75tqSYCHzlD1lmcEE+An3S4y1oVCXilEz2ZAH7ebqRR5LCNoJN9lL4LGkmX3
XUNdiyXL4DkWc2JghPX2/AmEV3AMAfk1iLwTangxxQdJOUArPsYYtoFWHCVm
6enzQhTli6IlHxlL+W6EdCDOPGX0HDd/ZzPyzwio2C6+GznVgX96wHP42esn
3XDTlyAd8XGX9iIRl+guI+SJynNi26762ORqTBuJ6UTddZQNUJCdkTTea3D1
DCvjt671Oq6Loz3t5QUblhR19ISgoVQZLAwFM0LzMe8RlbP+FhI5NpYfxTR0
2Ftpm9jrzKxpQ0fLvlnlW8fAOt2IJuzdzfM4g1XKEdb78bI4gH2X6XYR76bt
L5QD6x2BzuIaAOw+iiXVNdirmqPEvW2HOEiGBsom+Ig9ErK/jNc7QLi8HEoE
Lz381VOIkuzYnJAWBI3IlXtvpMDsgf8RcDICSr76TDkvGfTUT5Fu/pxSE3nO
ED8cZmcI4f1xFOCwInVN2FF8eG+FVDHx8QCWgmtaiql/CuY02PsEGGy3qEuc
k7DR22oZL6zmcUWy1pRMkv4WFNrxRQ2eb9cUHn86mS/jlYEEJdGI9heGYnn9
/P2Rgiph6QULRpZ94Bg5wVJ38z0YAVii4znnvk4bSb76E8vmMCyn0kEPwyzN
jP6pawxNKFForLckwBFzKE7e7x5bZ4pkTJDHaxVVQM2S74r85rl3Rxf98UUQ
P3/YlAkNbokS/zvKsuoiuIPhFVWUTvQ8Nz4sBfXOGxDRFZqOy09YCEkhS3KX
xE0v6RJB5VRM+sUVWePWQ6OEBjiGEBGY1kLfGCxGag7LE1c2PJ5M9nvYe8rB
Fv8p/G6J770/fFsENn7PZy20a9UIv82RZKAFWhjMX8cU43FCzjbY1XrgYuUH
RBU89+RHZkWq2vMNnaHulRsLxcRCVgHOh0GQUd5inQLIfTglXHgaI1A4FMNR
5XtsiSpHnfVqkaC2f9GNO9q4z8w4pe4PlIX9l31/NSftquCaVhbQGbd3VEQ7
O1tDX2GzbdLdOddB4wUIBXsuGLKacO9SHq739ZOQ9Kct+OVzSo9AyS6gZqEx
LtD6iOSUMn5S1Iucx1zF1kHahFt/QWTQNaQ8lbLkvuo7m7qAthLAIfo4xZdy
M7k6by5LEBCANJqdGHd+qp5mfFPAuGnGYba4wnywSZTcyWTJcDREzeu4Y7Dg
ABKdGuNzGFEGvPuZnJZy5Kq9Gvx8kiUwJCHeKXIAbBCbr0hdvGg5AvIOa8o1
uN3r18IELqjzMKK4iDQmj+SvqYfIZH3HOcBuAH3GNwV6Ujs6m3EK3n0EdV3D
5o2aavSG3CKeAZ6I3QQU1wbkN7WDSYtZ9llE3UqBruKCwn5cFpaupA6XJj7L
S27JlvT95yX3sLw2KcYEf4JaDeOx9QscmcPu2fjvX0yAQczstlQGLnxok44r
gNHrkhQ1pB+f+VTtZzj1+bxNf0IZ+MetTjVXeNcTQzXYoE4ulaRihvL3LYU+
Ef4xVuM1X6USjZeOkAOgNQ2YzTc702vz3p12bn7QkAilwx9ZyXYLcDrQthV5
TBW8RGvGh3T28FvE045SyhJ2DTy/79HdwDenTSSQuQIxVqXGu5UTIPmLb40/
w117NMeSX/vm7DLjKiqylSpwqGxJ5ifbKBYK24J4pwTUb+LOvqr9lZF3eFbi
NIrOG2YTkVmINyovAizkXl52Ws6QGp/Z/G2JxgEI//SEMEOgCIX49uEp9HoY
SYGkj+Oa0/2Ve6AvS2JldFf/RY16GTSf1WANLQuwtwDKki6XT2MARdzYJKyh
Kn0loXD9RxDmcGGLO0VciWwsYey0T5vxtXh+5oBkHx5o0ISxbeul6CaZfeYk
EUrwp+0nLO6Eg2yRQn6skkSLTwiw82N7zgV9pAFLoGUVZkhO83VteNtpPDSH
kMKUYA4pqhI9wRJp/jdPVD+AuXvpYKYyh36vqs73nhKniyts29GfHAebexMH
T/tmQDyXGMuuORqkEcE8E1hP77lDiT3rwAMnx6pBuWLaR5HBf8DgLux6SA/U
dtjGHwCwH9Txwd59XLw4p4NW3v7VWAR2Jg2ohDtamgclKMqEmp9hKF/5gkGs
KZEd31sXByyjLzbirn7eyayZJlJh/VmGekkJSQHfnXDG3JvqhnqxbG35SNEF
FMzC/AP6urTuud0J7ErexHhOndLmKjULq3zhIzSKgzSR6j+vaXl5ERFySnx+
ZMcMpuYP9tfj2kTkBw2BCcbzQ38chT2uAVYrGwoj2hEdCuLkO19wqIVxo7X1
EWtdqohhU2D3izrL5FOBBzn9EhG1GvpOCdSAp4uXEKu9NNnaGndAFomcA50H
qMOXJgEMWql/urNvMu54hsef4awys8qPO9VB1YO2pj2VG1fdQAzaIeZrdC30
rTW8HFur4p/fXvlUFYiw89Qq393+86v9QQ1dIQzwd9zP4SmqhTqLTHAl9VLP
stC0LMuYUjk1xesCC9UEs1cEFsfNTZYU2xmK9yTJF/sU7OIdW5vYhHEMgVJL
xlzDhZ/IWEUpgoTwAAQkL2cwAdf3k7vZzBwarBlDcNMz0Klqd1+dTkdJk2H3
rKRrw1CRVD6Hg086HjttQwIvyVLOij6EtTwHkP03Yo4zOf0tVnlCtx+VkSqr
H9gBtQcWJPLOhjIGm/dwP8VP4Z4bxw7x7DRvZZvUvoXmOkQz6N95yxUxf3fO
7uf/Jim6ydtlpJUf7jUbLlfi0C0I9Q4ovpPi8v+xZ2Sehn+77VIG5pg6LUQL
kxT545vvNT7VB8WjqBnGUWRChZaGTcduCaxZw+rv1k7ApdPvcrlnlhmv+FYT
WcrByzQq7tAvaFuMHL4bh35j8yccXVWLq8JHb1CXo8o5FdLYM5n4nM1xqYyT
nK9dlVnUVC9inp+nNn58V81GMmLtFJQq5v50J8RhqogCfXEiAaSIzaZXH5Z9
glX0qSj0pqX2a8DznmeLBsPTSLYgJNPlWQiR6bXxOItDwviLt+cPm9+cn8Bw
Hb7oZ2QyZ8a0qT2XnOJF1dqHtJV7Pebkr4EoYFA2Brwz1n2Ep00aXt6u2VXv
ys1tKpJ8pnu603Z3SIeOegIiG7ymUB6jIb9MRlB9+h1bHtt5vz9Zd4LDjiB2
a1p2jIlYPxayvN9qoNe+QZfM7y2dOkxQpxPOaco+p+MZACIGfU7dTroaV5LC
uuRRNFjlsQUPFDtElynwa/O3jPbqIU+GjjIR81DFHCMMRyEcwoAVIBIyZ4V3
9gMM4RGQ3NmZFGKRwYvGT0WQV8UZi3EVbH2lVhwCAvWr6EhHynprWaqCtjg/
3UM4tRm06DctnASNyG2LbfdFx08fM9SS/nF9KIUraGaAsDElg4BY8+XJoBf1
Vb5YNHt3ygfwx3XHGXcOftiNEeGWvelX8tcvrAki7evqyNtc7PzCG25ozuaU
GE+OGjrS4BVNB5VW8TxxFmcoQlFF/gD/XqQWHsIxHtuL0tgGPNbY55Es0RRO
SbkwMSpxppbMu741UQyugaXK/tcPT7FwQyqeb/QKqPiAx4oIVOhgagAtiH50
ItM09SmvLqCukrQOQ+SNbZ4O0j/o30dkoqSzUdst9LgslM3SjnJn8mECOdZp
BncD7lkQWioU2SEU1QQ0JT6STGQgxqk4F742ZGXH6mwEjWYZi3ByEMc8u9Ld
2jjuw+qOyoNdprKWMJvnI9JhgbJ+SM+ocaKAJHT2xtnnTGDadabUOIXfE2m/
uq2aaAiM6DDNXQD8BsJKbYtIqd7ut/WYsRwNtQuRzMZBxjdk6oJN7Ze/tNA9
NO+4IKCh6k/fqW8JUz5ILcVVerFBn8fYZY9lDg3UBxp5Z+257SRwk1Hjia7S
qA5ccptQgwPRQTwNpiThaMFoXqYasSAj6sDls0POpmWJtodh1ucHoxM8ZpwP
Xeoj5mPL7DlhhTdQZlnjq2ehMKb3ws8ZreNliJV4c1H7iKjuFDKhpL3lyAOa
mkb1l1PAS4pVFgBqy80jO7ksW4fNCuF1+OWqhx9sJio1b/8nkKlbfx8mltvX
U78twtQLPvn34dCXTaLywVg4iqtYZaADyVt/cUExQ6XCluKfSdXYcCmwgqlo
+aawHHsiaDmgpjVf7Od6BQT3YKPg2sNSQYMBDfoKQL0SfHAmQ5LW5yPGnYUP
9HLZxqX7OzGtBeQcU3u8SD1iL3PT8BitzWxlb9aJRTaZezeU7Daj+1cm7mqP
EGWDkLotAT/6uQe70Kt/HVQodAGmdVzC7VvNrZ3zpj9BBUIUxXSUrGoQeKrt
EhqR11hBbQa/qnLxyw13y2A7Co6wiLQjKUFHlriIUnDgqlOaed/+X5+r/Xbx
TLRzXSXk+CRPcQ9sCqxmBhjdJXK66wovLaWIav+ckPmv4NiBVURn2p16AS2k
a571u342SOPlH/uU+dj5BgHpkxv31KdPpgYBZUDbwh3WwP0NaNkDt1884iSm
Ov4ltRstsKfgRu21f3qDCIgZR0J2tjvilCyKGJzL9xVgncVRAoJ3dLmZn1J0
9Vdfh45lF93NGRZi9ExeY242RqCjCi6hTFED0Gc/xtoWQcko4zBIViRAAZrj
Q9jWG9brDO0DaIkn2jwP0TA+M7UxTFds4UASHIaq+sU0Rn6+2nApvV1zcWlB
jQtPDfu3ZLd7iHaHCMRBgi2cSSycnUoYQGKSbGLPZ8bF2ygqxpjKHT42LWJW
rnhbb20Lv8w5YyzBqmytuBJHZPTw2OwxvDlGv4zRdR3l+4ECWwxF5hkAJSnD
0+QImqR9RwOH/iTAyA7/u8hNflYmDgZJnzcZzFFTWiSAzH7KLuc+kFpBB89f
VCItwPZ4vUpZc3vl5PC1qLdATfD5L7oxjAQj4E0Z61YYHRkDABKi39DYZLCX
KNsruZWnXsiU8/htwBl3BYr9QrwYttLZjJinCVKmNuyCXjwJcfo4KquYJcpg
GtN/UmY+VVw+08MQKESNHTGsSA/jws7WLzbfPWxWaLMBbycM2zcC5dXkmWuu
HCCd8Y8Bvr0YxiKyiAJXvhb8Q8h6l/DHtCuawRejcH+X4SgoCMdT6F6oYphx
eE3El5FPgXEMkW8CWfn4tCHBJQnQXVYfiTL5+7D93RByfVTdzI1/Os0zBCZm
Dp3FDFxR1o2bjX0y1YFJEFpfcgj9b3K29svdqUyagQp32092MYSXEHSKqcm3
Vb9tSzBUHFg3tXcWWmXP7THJrnkC8Jp5aCuItjevvkuzhrJW0LxSC+eim8CS
8kwRnGw+EWCYpdKq57bbW5OcNfaY216aH/8CCHETqf15GDv+obRdEQ8ZgPqe
4qOIq/WmHypA0gQqbMXWBpQ0HloEdfVu9PjfDhumqsAEA8+JNoDEXCmzL6LB
znRdAUWwX7eOerdpmeXEbhhIasOyUuHGHbFF7LrOlR3tNGiyN5tLn9bwiLfw
MxXKDodAPeLdFFffeZyBzmbw4N4yTGqkISq+qE003LnHtH1hdAOo9RIhyWEb
pPviwl+Rcb6avevofuUBVnZ19oD9EesWDyWs304DWTS6zV1PHhl1+Xkto+Au
x4273TX0iHOUcOMvM9WOFFAs5DgVR7q8HyHvBgrPbWLTPsrFhtKlzzTeJB2l
kN34qNF/w5Nd5lrP1E0cyfLwbZ145O9QZYVn+vtO9u5qNuUHoh2Jzw6e0/dJ
8CfCkDAmuSKrDzvQWHCXC3THcVMXWmm8tXDmjwG2xDciRvHt7q6l1XPwVZ70
beBjVi4gOUxcq1Fvq4febJ5AOw219yjRNNez6xbR10Trsd0qpx8cCcBsyVQJ
JBP45+ABv6UHsasUVkMcCMsDBth1oU0o5Gquk7VUBaWePFFqaBb10uLjbi9C
nrLgP1hG7AxhT3G1F4kEg0QS7SCfa1E9LlAkpMD+GgeL9OtrDRRga8OePPlR
pG5rvIM8maN7Xzhk7Fv4vs/mqexFkxHjvRjYi2cgWHDu0nHM8SgA3C5pxDtt
zdeo9/ZmbU3B4eJdaN3bX27u+RKIFF2tC1+/2D9/BkFv//Wolwi7LXMRkRcZ
/o3aEHXNWxxraF7pgJQCrhI9L+q2wD5JztWsCeWz1ry4Uk04i0BuK7G7oGxn
MslRnivWxNekSqcTDCTlXNGKXpcZPnU0WS+ihH3GCO17FGwRCYfp/ZRK5DmP
w0SfbTjVlrYdN53jDPiNztCL9kfCIkTmE4jzJxLhX4Hj9836IOHuxHBATR4T
uPJD6DUAZPFaE6kcr1nZYb91FPJITeE2XjpIZjvyd34hk63/M7oiOdA+2toh
bdm5VNAmLR1zQ+n7NnrP8fhllvKkrFH1alyTemUa7erAWAtA/kD/vaTzdesW
dUlVcmXnPu220v0bygPaLHyif90SPrTeUVkI1wGtt9wr9wXPAs6h86gr0Z3T
2UZ1QFG5tlWqnxSuOyLk1ZZWwZBM46GweF/thnLwN8MNQS5Cqr4/mGWOi0Or
iqPyXcq8QbYJnVQ7+rk2MQY+olnsBctdsKhesbIzi+47OLcggHq73ZWo1PF8
IqLZ9qwrf25r61XguCF8UpYIeTaA8Sz+yyNyzJKEEfL8CWtcx5RrYs8AJcs0
CKHmfljHrUifCxcXPW2pWiDMUdqq/cWyK1g5vQE1rlEVOkEudR8UnzVHJctA
L6mH8PuneC7Tg50abDVyyWJwpv1ZPj0MB2i2K+hNxVQfEngc4zoKIhClPyte
G1RTevfQwTaHm3Z9ZO99s3ah9u7rztW4PQ+Kk60B2Re1YWP+GH/46nHM0+/6
JaJ/HYUviXwXSewVWXlLXvHYWiHNRvJf+/rIVwh1psSXIDdKsdIMiS/v4uhy
D+Qo/VmnQAyP6Qr7tyNhU/QCghxD70c0UxH/EN8pd4QKVcHJF5np+k4xCcR0
YvV6mMsuTnMQr5kU4mpOUasJuXoGJ6bCT8Ow1RxZQzTYSr+xgepKr1uNEXyn
Gg8frUvgc1dis6alYW0D4p2qbXqW0BjnFGL+VqIZNEIOWoXZglX6r7Tw268+
4/VNjzkGiz8+KOCLT/KAmjAuy+a2J0gu/eMsPS+95j3TgGAOB5NfyLaUaeHu
S+6d22Bi7BgX+jrFBOEd8Q5yM4KBOtiuiLz7FFZpbZGmTemue4hy05y+ApJr
FcluFAf6PEeayysn79so6/3m4QNGy5Blaz+2T/U4kME/RzPaTjJ6lVik9I4t
bMHz7TNYlGD+SLBiys8hQcQIbpGYtQXYVzcEn6W3BJhKmRfTRyInlKzntJtt
UqyXJ8SmWURScFMffBfXIViU8PWJ9wMqSNrH7is/Oqg6auwEgb1LEyJSY6t9
FfupbhGtqrL9u1VztX/V4fADRSKpZzZ6FM/mh+AG0PuZKqY9hq2yXe2jCZny
d7y/lTKZ6dSDdWzCOZry7so9BK2fvqis8iAA6485R8dxepNWFcTRDOvyCJnk
oelXnXH3B0BAyFRV7b1X/OuFuYAOBWIC6XWwJuNFEa4mBGLRjlSpJxh+t/lD
Hsoy4oHei+NIcRzcXfK/8e3ASaZWOZNnLU1sB/nW0d5TxvqhooFDi8I16L/q
vzGNP4SKJWDnJAkE0lBUh+9Ri2ZtFuQImWa0SUF7UmMYfzPIGPViXowMqmCY
dKFRfV8jjsblynOSvT/488HTyVegHL04WaCFIBkNDr0K9u77f3ZlyiBuspRA
HcLzecvMOQlbCaWQBHnDkUpCnNgiSJ3pwg0kxOWcYCBLv25UF0L0Kuq1Id8i
wZZJ+ieXk9hji7sq0Rm/kLddgshwxQRTHwWs8yYbr2JsWk5SiWqsvT+cqO/r
6Ac7rLmfCcu+AJ2xaDVdElUkVlBYVNLa/LcFfy+lt7L2uiA0xhTiiu9VKvhh
DY3h0LBESEI/HnAB3OLb2g+vq3ycHnuLxyIr3GVNp5LarBbMruRVH14/JRfI
ID533Nm5c31xnF6AESDtg8qrutQ2LfvVBqtotRp0k4miG9TasJXQ9cV+FT4g
AzjlB7UW83jcbaFirErz/T2PGqJ9EYK7cBQF67Ekg1oTvrUIXfVMlah0HqVx
NozFNlC59foYIHUG4/3L3cjiePozN7moQoe8Pzk8Ui0KRH9W2YvUHUY1y+K7
XXLKk97xPy2eRsqnlmIrcBzfQaihK20BjrfzAcLkfs/jVWyPXdQGHNg6paEc
jh0CMUGbedLLyH5J4VE/Cgpt1sM9KlI1ZjvT2yTovPFtmUZN0xEf6jFSNzq0
HBUaiKQ+YTTsf9dFuKacGxcYBwD8sNOLAn+9BV6SzF6pc4cBDn1YgJ3/NDvp
vuH7YbTv5n0nsTjzm3Gf3eaLKgzbLcp7JwaYR5sLQXAauZvFxjnR3ZYxd0C6
QuasN/g644rtzWnisNOC+h0MFIBjr0u+F6dV+9qmYbTN4xaca3a6ba2oreSI
zp+fcZAdvg8stRsEMLoNW7FYMqpbdplJXBxBuemzJuElSSqS+t1JW4qWFpLq
TdhtTmo0pt0ItYWrZUMj3WuYLcQ7wIf4HJ98PAcMCX8ZHch9Cx2GX3S+27YV
jsgWdoMPwvoD9YTXw5h6Qo7AjawRiZ163+XkyIWg0mGKQzBk/uDS3bILZVYF
dc0XQZX+CG9KusG6EidqFFRBedzzonBjNdL6f9dnLWGzcoWl+camqervCoZL
3wah62KZ7DeeebaFXzu2iC7krpxCyBKGbbPiLJb84F7mZak+whAp7iXosdUP
oAMUoqcvs6gb2R3XtODnHqpATwVBe3ThQbnycQ9KnjUyNmaCR8tha0HqwEf2
VJz6rVvNMDgTiRlEONWMCN56McCkn1KBog8Mf3JuxiW5/ILUBuQWcguB71ca
vgSjCnz/jWHd598nw/3TQgTIt+2vjZstLAy1sxwiRsqXBVcgYLRS8nUsDL1n
lomhYSAh1OCCBw2pOKTkIIXH9uli/y7Ti9wC1dv02ygQ4R+PJr6NP3AKQv55
zdnBh8PAxB1jkjXWh2evG5JuQs9l1Y7Vi69FRhs+mFAGKg73HIU/+CfmvF1t
nIOGKAdBgWULcG63KeDUZqtPdprHr12I8Or7bNCJlAgYOHEVzMUG4rpAsGiJ
EEzCA5jWl8DrqG0zQIgTtuqjbl+fMEqO8SRvNE08dpOTXH3AGGPAsHFTLhKN
/neHPfJDLVovywTGUOayFMp0OVEnnJ3pW5rbZrMr7bQXpsQ/+uTsPLqdfCid
xZmwFxjRhchouG0n7KC4PdG7sXgUczuEa5zdbUEvlAxMa7U9STtkk0xccP4J
lrA8oIP5mjkoF0xm85ckZR2Rk0RpbNeAX75IxuVkDbtzz2elm4yP+99YVXu+
ez78KWWcyvGA1hz0BNpsNfwf/izG3FTziNlw9A7fNNskGAHt8dTlNP5SRTP/
h7TFnzWIGUaplcmqRsEGfKobKz60/wIyp/07BMfQqaQu0PHr8NalVcBilSb0
HxWbM+UxZifCkI3llWTdo8JXm9OCx/LjOmS4lCjmCXtCbTr1AGfGZy5GshVg
Dlsgg5GMBry593lpsP94IBCDcPAqUvgbSxDZEaaiyiGP28BxwjmrHZoqyPjO
0p+Fp/xB/0lDrIq3cfV2UZ1Xa/ZLUcINhZtIa+koLQJsP7Jj0fDcukYFd4Gw
uxFVPZHE2jyyDDQl/ke8YiVK1YgVvWqzkGF+7NFyz1+zNfNfI06SVBzBR6AS
2jGERWfadD0yvbLSzIIc3aaor8DrCzlVj3Pihw3iLlWhC+FvrlYAsRddUIgf
Lm/0zq0UVogiATlAk4Fqg4Y9PpzqdB0X/J0sgeB77DyihZ/3TiX7khut333M
CKp0cIaLjOrYwVp9UqogZfx/UtTRwbsdYd91t2FIOZH9wn0hPJC8VIXBJ/TA
RpOIYAoVWWOkpvFJHm1vIFe/Gjk5BBXMiYkXI4thpMWDQ2jz69+hqYdpitzz
suPsp5IGeEIO6Nh8VxahNECXi5SSXe//21KLZgr44mepImXn3OLjyxQdidjX
eoHBumjr+2PUMtEpZj+915sBdHT+SAhUHjm5u17nEQ7E1hLcz0K/Flv/zZEf
TPArosOGou1udfp7a28m3eoMH+3u08fR8ObjJuWH2GEjxDKvizSGgJcM4AhN
H5BZ/31eOtLA28Yecd+y3D9PQqPBgJzoar1Gw8Q56gA0uD+9m9s45D5OqxPx
IJhi6vg73aaDUtRxPiClaOeaQ0fsfocCZ64cF2T+58+sF0LnuhAzyPrlYBLn
d5MCLPQYXMN6BuSCgCedqdLvcEcxpPszy1d6ZFWQb0elYOZ+xcLI/cBO+u3s
FD7qsQ3iOhYYN+VXhnJFPsIUl7//FAqis029uDbT6ERLfvWJECp4MarDYc17
u6G5DHosCJtxMfYi6cJhMDY0rcnkaUL9f/eQkcfaW4whJJp7O8XbOLpDGagU
ckPa412Bc61Lq9dnM6MET4Do6+u/Qaw0ieLrnQr3/8zvpMMIsij5aRQjQmYx
mivtnSbtxgvKpZf8tJAl/5nvrtU8eRt9mLv+K/qPeyFot/d2XTvR2CeunL2/
LgavNEtwWiiepT373Llxe2sAP/xxK9LL00u6tStZvXoGE4lxDT8eWc9qv71R
K8PYnWE/2B1mdW5q8O8Z0Or6Ac8q4R4nkCf44TyBQDsYAPGuavI1nuYSodWq
aNroGyY7DOreRikhIQaam1mXVcXNLZDCQ8zHRjAbgK/YLBypv4xIIa376qHB
y2rpz65Cc1w8YZbw1sd/WZ1B+LU4MUYGHKDTxcnko2eP+Xg2J5HlhOFYTSAi
jwkzbwPZrmK5FEHBrSbHSves/2vbq8AE5PMN/7XfUO/KzR+5dqIsFXJMVdQd
+KXbJTebJR14IP2EcTela7TXAaYMVw1tKhzpQMcxjZ5lvuTSlJUXIkod4dka
TIoRY1DoryUmfdvvQNtSf4auqrEO2UgqsjivcQaN2ELyJ0rzty9V0UFROSIb
HrGcxxkIZI+cyHqKuWdHHae8HYQ4caOZ3v89iZATpsNHmRnDBMnLzWHzd4R7
Mgd1fojtz823DzoWVfM0KgnjNCRaP1mAmPH6f9DYQm4Pa4AM/xMo1xNkmdFr
JLJIC8XOgKMFEFkK8q/SFfdcxkO5tsejkQTV9PEeEnNQpzz8Ymy8zrqgwNo6
so7yBTST2U7j14FPXgjFMKAV3/cMMCzMAexbl8H7p/ZQ1dt4DtXjn+5kLuTl
HAkmrJFoGxp/D7FyKgXoaUdMb+1YqYzB6Zcu4krRlN2d2ouqmn1O8e+PmTuj
z6zZcmBQ2aoRJqQPQ4zGnS8CyI6pbtbIrFzOp59FC6PuSidR+RrD/Pcn71G/
9SlZ744HC9/7KVCZkZi9pdX1wnXHVFP+D++r0r6PQw8oD6VLkWb945oEzH9f
5eo9KuNbZU9G+B6PArjrFUDa3NWFrIgn1qRb1aNgHpac03tBW3HsRJ1Qy/qg
J9uiYLaNChjgkLNwnV1zXzFelvL17GE4xfssOIJQy/O/ctq3VGDniQU1IGmb
g34XOvUjyWclmDvjTEEPvzJX/G1JTZFxcdNwfednhKoeoMW/jW92SeIpYyKX
RraJgWbPtAhQSspslukZm/yBgE7xATe33GTRUSc6DvizzDZs2XWa6rk6EGYq
Ouq29j1Vee0Q5SvJ8Fkh9pZHto6lzPjHWxJFkGqbNjE5fN89J5+3lsXKuJKa
M5inqqORSIlS5Tc3tPanSDNMiE7Xcss+NCPLSAotnZwozT0yo2kr+M3Tw9aZ
uZj1qGuEIaYzyQUhSPpGCdN4Y4fBUb/nm8rQlW9cJMI/B5uso8EhuA1Yu5lK
Xem0pZV97P8SPbr8hOzIjv1Mrc03ns/galmflDMuHnTqDOlzOy6/Lc06tuJ9
YXuF2LeZO2kFCcpDGY18yX/7x3Bn0LHMxZuebINHjdtBCNGGv4FZQdFepzpw
l7UXCP3MjF1sHn7ePGXROXL/B/FdkIBCl1pIlGeBq63AQBFG1570u7kQPAH4
M6ssutx8hy09f6kFhE9U+OzxYvIhEV6wHhnLJHx8lZTkebmrFJiqpa50JptA
bxXPruM5V9MA4cfU+D6RTghaNzMXCpset9QzqPEQlJifPjTZZxs/nQt03LU5
DM+yRh/cQBb1PXbUyhl5IsmW/pxLWQYS+wP2wVD3DpGvxwWOLWquUb8Nld6o
LhTSo4y0IGPPAGVQCsDdkD4/jIPilBz2XTEppbYjtH8T8YbxSkO7QflKMui+
nrZ1XBIE9zqJetXWy2MdsMcao1+7iqmWGZ0r82Kpo+UxfvOJzlUZ0ceA/YwY
9mwXbB20JFiWfEsklN6+VwDo9xm3cw7oEE9XJMLwwte1DvpO9jrXo4Xg5ECy
SoG/DWX61OfHme3dgGVO9yQFZuAbVPYX3qcMVL8CrTMQk6qz32Igqk6RJblv
3CpFJX+v8+ql3SMxz9ny9JqZePNZXG8StW/wpVCJTg5Iw8mavEyhsSDLrDdf
0FN0sZhRAST06GjG+4FibCBCc00Ix+S5iVydJzXKKZs9ff+bxaTYzUda/nn+
u8ibEV8pokj18PLWhxCgliKKIkYaEOeva70MlmJgQfFEVgNrYVoLd/ZNWI2s
+q9zU80r8LTpIrxwV5xtCmmEJLp7rRf3srQBVMo+K54qln7a30JhwAp3Nky/
PZaSRTc8QEbfZNebsCsAv+AETA/bLTJnhGAAhfgdM4l0xoTM4JYbAcVbHAj/
WJyN4r87xdaELrka+GWFBcVGsJCQ2CgDfr4k/VsnUVvsBPX/tpXoEF0g4n7Y
kwYEPpMAfr8beGsbRMZ5FQ1ZrlNXE1mHPBXSbto2dEHnuSEsrWsXDfHumBbK
yJSZg6HOJPQqwWlzKgQkg4wItjWTBIzJG4mfRQoukYmmiMdIhPTG5RgIEBoH
OuZS9QpzV8m4yPPTthU+DTvFIjRD0pkQadTnnaOT913F+9BzZ04ky3+4F36i
qvRgLkUVWvN8f+AviM9Z1z5J9+YfVPa2U6BqebBIUa4HHs2VYCsIpNalSPo1
8ksVZf+JhH6m/7gRubPJ9mUACuuwrRU+pn4e60hkvVAt0Fyrom2pmlFkPzs4
zpbGBp0yfpSfsqFJyD6SC+r2bkP4UMkg7ELO6rrOJGWUj62aoMxNue9/u6Fw
sc7KB0GnfaCaUKDiWhqoliNuyFNebIB+bI9y+2+p2vPVSbEW2AOmW9AnKD8B
z5Mg+aNKhLT9L4Z0JIg4fve3oChTb47iHLNbC3TSug8iy7CzU4gps469egkO
n0pYGP/TvAMbSAuJzIXIIzvU6adSO8dOQ9NWDnNK+DnJ8Bs9ECXmnd+GnvMf
vqMjEadoPdofcHtIJLoi6cqXtGcEgr3YL/iHgXyLKj/6qYs/VWxAZUHoy+IZ
p1Pid85lSMy0SbXGH8sSFIE75a82vOrAri/sFlKu5KEhmbCnCHV77KvGAsRs
Dv84AEo6A8uWGmxltgLZnCPBlmfnWxyVPTGZsS6ip+MydyIeAGX5BljqPus9
lleHDyijEQPcJIr6xU+I+e2RNzJH+0pGgTBzeHcCw/IyidVjlqoWMIb9bL6U
KsevxdX3l7mRL5rzOfdTBk/9/HQk71jQqv5CDjmKmLM/MMJIEtRatM9nNzJk
uBMBzPEasQzzeC+dPIi/caKUWr6bBjopDZSr9mKc2G5uOOKyKdtbEk8hXdDC
Xmc4s14kBvz7dJdET7hCPOgEVAuOv/YSUuBvMuxMLYA4v7CY1cQCioqu4EM8
hzZKd7OcJDP6zDIzZi2VGgzvAl6VMbDmIbHXH+483hAS/TScKxIZDjVgXAiG
2N9fgv7A/D/FgtoP72Lkitk1aZSSlD3dp1ai2G1gxNagZJSicA8lLsm2ExtV
IILgxqajptGsCeWjRR8MZ37vZ/B3qOkpTljyXgd7YJScN2oQimafAx1XnFa9
hkyxnSZnicjSD0TqsqqR5mUJt6g859dsoBwiaP4SXMlfxkco7/7P9MfTAO0T
u+7yNm8T+N9UNo8RC2Is/zcRMnUwAcMslZeQSUwyFP0JSnQQDh7XBcbQcbL7
c7ML+pcoe9bSJct6JMLTbTJiW98Niqqj5XThOGa+In8ymdj0juz04n5zDK/a
RYs5F8PmEqOa2FA/VZKxXXVbVr4b7wIzeM5Eo8hXwTE/148aKLmj/LOb4Inj
fML1Aei56qPKGaMUTfX8g2vhtgYq3QMNkbC1KyNP/ayPgLA5gi06oJO9cs+z
Oq1UjAnWk7hIIn2pziFpAHOY94oGK0w7hAVkeYceTnuDuaxj87IW7ScwsyB0
zpnM1Yuu9aG+I3IbBL20uFJt6diabuKxKJONQu6zAc7owBXVdg2Rwikb2C06
GdAAjaglArLNs35G6mVUVsXyzmK9b+04YOoA02qInN20G9SvGNQeJvlxn0r6
AlWPkT9BYTMkWh1QKNgvrh4JxV6gpcRb7d85Z/Pnj+8obdm+l+LzeDAsRy6K
qV0WVeWCQath0cyZnhW4GO6JYlXBZW/B851CtDjsSHRg14JcUfqehzr5yIvA
bzdM7TWI+9zR8v6YOXI2Gh0bcJfBr3XBcX00LoM6c0mi/cR1g8ILehgBncLm
Qvy/DeCDJOxvsdYA2S1R2iq+Bza4wcdk56FQLETZM3tCERm8kJq5yJVfpi/r
2HpeDX65veEnUexDDs1MaC5eVvFTaEW3MYwmTEvmdU+Hn4lKzBP2H/i17hij
o3iHQd52pfzYS1tNzI/9oDvpwiPxaNq4Zg5q8iYRWpCFqm5/ofGkg2PK0XSG
RmpRAQDmuIFF2Jv071lzhFfbeNIAGf95rezEKLWQ6IgyqqEHzBmHBSCV55dL
0Y4N6aYgG75Pq2/lKxWUklLJdxQC4Ja3Dd0X33MhrpLh+0No6+1JwHzrHGwG
EZ8OdKdZXOezMySRZ/zjjMq0Mg5K1fXuCxujSBk3euqZcd0itOeDYff3SEue
sLDajv8FOA0O6ptxZp9DaBmYTXPKkOq3xEkw01FpP4Q0Hnnir/NLXnZcdzZB
ehVTBV8CpdD1TvJClvIoxQaywaSj8NL4EbVFyWfmqmPOlstWjkSaO7tP+BrQ
6hyiqcZh47zqvsdzMoNfrpFALl0jphQ/XXX3UfCAULNtgsPcu1i2AV/n+PVN
i7EVlUfbzKVfM/CDGO8qJlOpoKVoeCPm/Wm+0SGJraTvVrNziec07S3FIjji
chX7QpDgC175gEVL4hWLUu7chN89ewK6T9wzG3+K9rE9+hDNO4KrlAD2XJ9i
sSNHI9Ug3thwj9L8PMEcIxzYLndR4xyvt7PfIW1S3VyH9BY4j9VYTN4p2tZe
q5s3U/vtPmDDxOhLwNfi6AF/N3YgTJNq5j5Wz7cRoggyTrsBIj/GWAUKXaA1
PSRvxhU0/vlMG0t5sDniQfUHflZsZJireVYH18Iu1VtO4ZMcWY0kE0hyDgdT
nDnhRhC4G95lHOI4ZjBZMZbW1prh0NADVTh0UZr8v/il3XnZjE3WXrMgThtV
5PgbIOo29kRQbhG/1D4lWaUvf6jw8pZqB/Zq9gJNHQ8kDFWvuy8uVHjnk19n
xKnPpaLm8imlwW6eFRKM8DlhZP7yoSGTRHwX3KYSN38ldWhU4OmeBmBMKVfB
njgay+H2L4bTU47F+6ZFmEAUIzuZktI8fDtVdU5/d7qOxE6heRCc/oaK1KUj
rGDTEWxWcbhyTfjt3XxMOJyJycyJ1PjDkxrTvByN03lBrEoa+JBiR/L9VXQx
8KuMzFpQR3zjr18jh0dsQq6ImBEc1as7IgTjxO8y4lv9+/5rdufY09a+zfk6
9cpZD4qUM50T+likQ1i8rhcG/bgfgi59vo/jJTx52MfyFWx1h8r+p2PGJRyi
tgl3apk1cU1IVwYe2QwTixJwb2NIwXKaEjeZlkqnCJPWgYdbrADHgemF8ngk
b/9p9co1HdF4J4ToI50byP6FBrb9OIwzfQwXbKKiQTo+olewKl3GYJTR9L4p
H3WYNdD+WimulZXIdcGLq/XNcs2ZBjOJjlR+qH4KlVhkr0xUCET9wuU9oATs
iV2noY8WvP7dYnp6/P8XeLQoCfuXcoc9bMFQCWTRBRP7fi6Ldu7y5N6UxDEq
ovXYmvi6655nD04t67al4angUePYTHVXN4Y5DimhfnvTfKk9Kb/rXHQeH8mR
QCKzwrnzcaaXNkm9AvHKE2WB6tIijotd6yYw+iijeDYjAlbhHLp5JSNAsMeB
eaVT9OATPRv9CqLLfrGpPsdmS/gWV5BDQ4gNE3HhHy+5J7oAC5slARYCU+J/
HvJV99rSn2aTJiRyGoRIRtrwArynNwxLmmoumkWTLKmJ/9M4w+ItW1vaKaEo
FepLfFbknRSiVdrHGQKU9Akao9afaRIfk7vGBreXqdbQQhNSARSozASnnfFs
d6+Xnz5Csbw1x0rEOAgtNwI59Vjus0lqbZQBLU5C0iQqG4gZvEyEbVjn6lAV
/E4OwTqAgQjdi4+n7HTNpIZ0b6RF7vrgkiv8Qqcn7tYQhmIfV65J2lAvVqV7
nH9yQ5dWBzYv4G2rzrJGfVH83LC6dLPAMNAN/B0Owf+slstCeNLuDms4Rvqq
4KZBPpteOvGCtPhMueCG0naeXnnvbzQlfzC5DDEWp1cNVutMiQRxbrS4JRhv
PmeN2/qtpZ5WanAoNI5m0FqIIjF1hX3X3+WH4dyDv6F3ZUqaNF9oYGvnSGQi
c4CxAiiKSBis3q8kcwtc2T+mxFgQf0ciWVgKjwZ8+moQZkJgWSJoTFWI+639
zsuR8nYMhXvIF+9IgBmWRNcil0eCQ7ptu/WcCpykuneyFX7Oq/LeTPXwxchP
XUYVKMABf5BezycqWDSbmnp3aVdrKYEZfQFqzpd+BX8cnZ9Rly2ODPZDD4Tf
9hI/ncqqkqz9ejyxrxBC04Cc9iKHfz0KmvTbMCBFQFcysmNdJ8Gr3RJaQj9u
epXqXBmEkQxLAKCBWAEAdy3fvWCTLsaYhh5kuxcEnbfG4+K36eQ9yt4V/xd7
zczSx+D3CeMdVwjoJHX76UlxoGVDx9C1Qax6JJ/OYV0jPa+eg/flJUv6FfbN
ZSm25QDtv7Jor373/DmkADn18WnTQJwL2lamgCzM4Igyfl4Rw6OHLDDeXmU7
UuQWlecoXi315VuwayLpVJntA1Ty1IqWrHk+qTYBTmcbNrrvqq0fTGE7aOJb
EKRHNyTj0HeFUVq2dReLGWKilFfbvBf39pvnjeoR9D89WeZNvdKVjyCmdK+w
nHYGP3AuikfNws3q1bvCWt80KZw8ZylspB5onFoI7IggEXZLai1BcgihvzKH
ZqD72DzAcgNMAnLWl0GpDFqtX97ZDcUw+Ujn3et/WpWvyC3VmjqaTHigDA7V
KvRfjKhSZmQAGYnuufw3Wii0D6QKWBXbxn3uiFHHH/+pFmmEhGcoyp8A93O1
B0y5NuJmeAvlg89rhaU8kriXTFFzA2cJBtjo0SlAeCU2LuI8ot8pjnMAT+PA
8ZXIIXnUfpDO5ye9SHj940mYM4TNF4VLiXLjusfb7COehFzoRWM3TaicUk2l
zFWyRC4dEVEgqNOn2LRYzgQhNQA0IxAaBZK8uNfKZDgHbCbpLE+XBJmSknvl
lHda1S/eJbqVtWSvuFL5J9Oo+ualV0TEKWdrzUejECaRWsVYB/horXg5oldc
Z3TQltI61+dcIo8JCgg+wUdPxq29b/e9ixBFQkesiUmUZaR7d/3YDJ53Qcvz
qzdPC71qzo2UdbRvY7GmZlH6PXp664lwsRLu7QxHTQhKzPbyKDk8/QQXX+7a
DmE4tfGUoU5ccktwDVIdn+xS8FyOFMLvWa9xuJeXbGVG9vKvPUDRp997fZl/
4Xx6KGaUP/mTDxgi1pXH3EdtHfHjpZQhatZQuVzxnQyvanjC1sxI6BuK4PfM
mXSsOe6YcT4aN+cE/8MRjvcRka8n9/8MyIQO2DAG+5+ZTwSlCfnQaWlqkxzz
sDsALbnm0Ei6cD7aivtYlLBPIMhHzMQQeHvSnt2+Yx/QmbqqrJsDhfZVwYHF
OlNNW4z84ZBXFI535ebv4sfL1MnXcpw6voYUu9SwGN0w9fC31t8zj24SKT9q
h77cr36Hl8+NYvbcIX0sauDrPWkfngYdXAd9aPCZQF39pg+Wd+5g7OIsPZOa
1b7bpcK43UKxP4+wEtqBaMTvTWtvwHJRmWEUJ8dfKy4cPkki3+lNSDhjtkF3
UyJqj+KTZZEX7C/KRT0SrSG5cB9OaHJ4X3UYazcFM4m1qufuf/cFodhjeSDi
55HbGN3TDYJTeNbYIRjOLQEdlYl17BFNV7wVt4fcnVflHALjK37b7zcJjyPX
MdLMpEQOgQ+NRpSV9/bG4BrtR+H+dgKiGrucJmp58tc7q+Sn7PpPyMHiPRhS
rlHjmTcNXRnWGV7iUkrnBRXDLS6hk+g2I+Y1eXuBP3fI1D246k2Kj5bln4FK
N1FFzEJ2RCil3YKeY0wwr4sDU+ta+5uXvV+2/qoEITyL3BhdyG+8kWX/FMq1
zW0+gs3Jxn7YZER6cnp4DAMHBQSA7+g69igAU9InrYl9ygMXwjY2h5g9ky66
rBRvlXz/lMWhZSjeQvT+ArCMSU/PE+ZIYuAj/nctOBeaLfaeFL43RAylMHfH
EvIkesxlupRR5TQyk1fwI1dEF/6051Swld2kuHMeQmcJNpgU78RuK3R/yTf2
LMhUD7Kh32bIfBFPtxmrYT2WuZ4t4rYNpWaQbZfyOUiZpqN97wrEiKNuWxcU
HTpwO7Q33LHTNn4WmcU6AG8/hi17hnGY7ueWHaIRGa1hBAzTbzOJ/UTCX/g9
6CuAl3TVzrrULF20/RbawHeFcvIRWxtUbEjNWGzuZAwvw2viNS4kEJ9nND89
VnHQNQeTHR0z+YCpA8CaROn/6uO101bXke6F0LvWusFo0ESnv5Q5PDQok1cE
DCRNseqrv/Wvy6GbI1H8OajwV0CLAzPGFW6RLLcb3NbMi0HPjIAB8CAmG7iF
s6ZcjxOPPCtlAqOB3u55lbrY8zbKWvn/OVzYwAMBHafEPGDbp2nMdzlzDHAX
FZK9QoPMapMC6AGaqxNHGZfsThmsb9siabFMzisCoNGF794vY27ZxxlqpcDw
OF8USPsp9LnVbA6wPuj5b3lS43aU70q8gvmFWYI9dIS+EP/bYiCZ+4T8+GNY
7LUZGcEYs5v+2SD2jWv0QEjCd6IDtNSgEQXN8aF46+B0QYK0ziUMQ/33XAfn
ATZ9feU9PxeIh+LT+Ebc7NPG3yBLC+aC2ZFlY6+3dsaqD+CjdpQmGAyVR1yJ
1W0huwJfQwkJ6K5mBzbMkNEJ3UE7NV8OAr9NVeamhxU8SCbaRveqs+nvpwUf
P/jie34UdYectcfTeA7Oye8u+UKJee4aC8WOLtVtg6aRf6hGQkJuenpOFWeR
pAtsfUe3KXEyiL2NeGBLvbqCYQIhp/l8591EC0PRtj1+VCa4OZfhvWztD/lF
n4omL+2MYg5HQ58CqGyyIiQMLo72BdasTKBQQqqyo+KGBQOAQDbhblYe5/2F
qgTCvqaHNO78BtJgRvqBnx4+clMOY5HKfG/WFXgH9glsjyDfIbNUcdGErmht
xmhn9UYi2sGMVLXM0YRMQ4ghZnHbe47n7OXR1azFdNbzIBCEuF+S0diWPHI0
VM/PsgfM72Cc9q5p4tNYk1k0edvTo5QQuaCNzsKngEzTTl+Qkxks7DlFBEar
Hah0H77gLXAJKYbRLqTRtCvUiEmbNsx1ncuOfQ3B4yAZiPW5/Sfqj77QtO6c
fqfIpVBawFsNyEI/SJjMQksHdOwmLKM1jB2IROQpVFhoabxAUV/v1IuXtvp+
Q4uGdlbxk0+UhPRDP1lcauMGKojQNbueKtCbSorcELf9dhbl+SG3W01xblyB
3E40zzQgUhK2PlETG/Kvjp1WaomGCcEBbwGTzm2C8HSBZlWQd9oOanWz+uou
xNJ88lcJH0av06pj8e4WNDlzU39lnFrbWzqoT/8xz3AJjwck4dPuuG0xwqhN
BeQQHZSJbU3Oe9tXC3j6ycy0Y+PaeaGOwiFKD13nr/Y2jj86Z6jSfep3kTW2
Ui26aQB8rdQkyZ1ckLwF451Zfxfc+eT1jItwurkgCPu6NfDRvPCe8lZyiABt
o9CtKkVaVJblu7bCZMnTC3uhsQblDF7/fiI392tk0aW6OSs1bgXimoRs/EIq
fWCxGO2cJv8eEU8XaMmaCbogdDZOCnbn6IEPZ3KQxDnGrusoug7fZrGnSPvC
0jKxRW8DPZrrSkM32ECzpyPOlcq2ICGyzAniuL/ZbFTZmp8j3WnUTJv6OeEx
j2nyICJrulT+eLefvOG+wc3upU92uQQqTzrzaxODavaw/osQp4+Fc/kFvlDk
b81VKW6hNnZWZzASJjCg9GGkhQcuh2bdiekjDyirjDpOUZ06Z4zN9+jtJLZs
l5+Z9Q+GFpUap8nhARucg/P2uyFoTRfvmaxAAkwqHSOQb9aTHW7Srduqc6+5
jpVtYeVQvNoGvwc1ZFhSoavGwbMI1gqFSNbu2MdG9s3VSNa6BhQxPcjucp7w
sNd67oflyTzhNTb51TR23W0rNu/iNfCBXAwQHh/4J0vuPeoeVIyNz5+tvgCx
DkmbQUaV4JLin+9xLYpx70u1lt9ApUFsj99GqkWrWStL5LkGviOjG1QNMPvf
YJttopd8ktdTVxSPkQvc+iypt4wU4rmvrd11Ss2A5RqrnvxjuVqkkuSlpAGz
p3P5i/y4yg1X1P4Vps7pnzE8mZsI1B2SS967xOSFx3+dhOPvk10eMTS71wi0
26caTUr7GkGrObYR8IYF0rO+M1xzcrVAR92IbQLA/pTs8FRfYG88e50KtinF
7IE+HZBp/3ZKi7dVUNEBTEG/aAWnn4Ha0C68wTBESMAFL46emE9I1XrFbJxg
rSoTvGmzzXydxybqk6pG29IKymPfRS/kWqECcDdVFzXDUhlZVJP4XvsSRN7x
YI6Ie1c6eWOXNj/QmEoV9I/DDoXA3olpIV7RsTHwD/Wgml+FOfJj7s1M8iSd
YZg29ZodKLA5se4dTTwfJybSKSh722RN/w/VPdvpOW06nbFwkEQbtvKmZH0c
JAV3d3BBAuwlhoELsoDYoWR18K+ujeXvtusjSXUV8bWdGu54ce9Bc9GTrZVx
DeVmJcLPJCCt9deA9C6rEtQF/gXMo0FZZtNemOLQHm1PGIIBzLiYoobeoj5e
8HPkDTLFFSJvvCPCKUySHtNg39/vkFZ6Oidwv04f95kYmEjdrE00td63pa6G
eQUN2vvwEYRxT5OAA88umi7w4kXafeu+n/TDM6pNjda6bu7A6+PmenuG6Es7
YPFyU6xP3XN45FsHt6UE0S0P6WG266X4FuRdRdWcIVIDnYxTRqW23hdcDNDC
wItY3OKuNAF66A4rjAkojQp/WuVPGJkRQ7xwSOTLZFPxDbwPnpdpR003Gq9c
FHQ8KvCDC3Jjygd9Is4A8unBx/Jc+VtchwN2tY6S+/x90YZFliTKo0vBYaLX
qZNFrzSMMPiBs57Ge1hK1aAtMNMM3D2/hQuPFkKCBUY13dPYLgKf8hz4R+YZ
NKtU9HjS8mN9rXwnkjUeWXgqMPSRNHDXkzxIcmii2G8OSmyQ0t4l889TYtt4
kRHb6oqXazs+KWkIgudkTRQnCdfulGYqm0IB0KMtwNlm3BXkqUVE3lS1CGt+
MwurE4X/YombBKym9zy6Q3Bjme2QzOVFG7Tqavk6PD1Z2LrcxjqOZ+HcaoT6
hJAGqDXP3C5EncfrZ3AQBcty8bSBUwZZvn+D4De/bRabawaEV6wM/c0/Em+c
GbXApNWBozPe8Uolt4I5RbPzgKd7NJ/LzetPaxz3ZrUWXfS0re4q3FbiRE2y
cqy6JwvKsAhUxb83yWQtH3NNNYwFMT6Wll6m9k34KbrvtwdxiR/xKNYP2KCo
KuA2l1ZAiZA3U2nc4UO7LuygEeIMigDWLqQQHiKhCEqcdQ+8zwT8lVoO26Al
2EHsnxleX56yfM2geILZQrfXm/eS6NW6n0H6g2sT+SlzvzRyctd1c4X1iMAY
10iP9iF1pcmqcuIMu3S1rS/dvBFKX406+lRK0LjgbCeM/fMkPUWMYfbiByvh
H51ICbHjZFgWjEMeCQUBZayrnYKAkbu7hmgdED9DVPMVUSuOf7WlbJfDZ/pS
OBrDXQEeJ4X70VrD9znNFl/5xrutuAH6gsnOiom6heBt8BrW71X5wMw7KUi8
vJmVYGOp8GbThjgE9uvmX6VuXXou159K1lve7cBwwSxHN4ltLGXsdvTI5oub
R60gxd4RrqOpRMiLij0IqXLcJMz8uQ9Gr+jVOAufL3N1zOvaj2q7r+RqiLm4
sLd43VcydsRrzCME8R++ydvJwaX4/VQ+1mDyba3MmxA/AcVC+mzZrKoy49tP
sTg3JocBhB0MIahaGSDHP3VcDnPCebSukcbTJg7rljEZJlewo3CQv18MumH8
9dZGKtRJVHo9Lrg8aBdULriS52OThSdXr6Se8QPXdPuezqAB6DF/h0m15sQD
I190+G7588r38QeHQJO7jJ+8ggVOQCkAfOK1qJzSJw7i4GTsi2uwReUxU3zu
4NFM9Y+2YGv03DRHDkb6OS96pLXAheVDz7EJl9SBU1GCbG6i+IHUwICKTxpj
V6s3NRoNE8KpllQJISKtqcPoj91RI6luKrZFFyFT4e337pCt5JmFMkBlh2jN
FHmdQ366kagR/VRa7ohWmSriWwfepd2GQWpUeVDqikLVE+IVAmGBDIRdEyH7
VsAxB5PY2sDQeGYUFecdrEG3M8XWuukK7nrIUlOplh6xa8lwVRFUgBnBMVXg
oI2GDpmHfevZLK5nZezdIAAu8utUij8OXTKbsZoUYESevzJcpvPjbXjgzz0x
PiHkyUj8pGF5imeyVvSiEW5uo/u3e4P4K3r3ZDA/iiTxzOeGn3TVLTgEPntp
4tmOyL396U0IgqT1j0ZzUcBfIavzj8Kmr/ulONsdfyP3kXiEwMe4t5GNjsiP
VHra3lf9nHXNJFvkRlIWlRBkyFyTrE1ULxIXNtJ22ctlnNxnatt/Xu087Zh6
ubDGqAZ3JIUxtOUdOozMbOxGD1VQfrNciVcsgXSYzyXnY5LPDHG7Zt5v/X4f
q9xl6qchQhkvCnWVKIesniHkeYy+3uR2Ck+TKxXTRir9RFmJd3AlOMcT8yJC
7XgtFciWcofr8W/LQHi/BJWWfAxHU287WBCGZqmSpqAX2sPsKPRrxLWHKfx2
0dRLv9lXgwhIIBQUQoQ6Hqf9aYPP4OgEKdMy4+g6bsqiu5uV29Y9Gpyktivf
m3VCbwjy0ytaI7DcUN03/vpW/zXqS3JtrvADKHd2XkUEWNt+strIEqKePPo5
8LToewmoRpqF8eKYkOah2wRMBOPpohfIIr4HSzVGxNyRbmnxbnU+Dpd3Tbv8
9zbmZqCvRuzXjkj7d7pdl+A7rBkpttc+AuD/CJCRebB1LsGxkcDF98E4OXhS
xNqK9vCF/wS9G/2lGuWTT6d/gbgCWfkEjKCbOAqPzw18ip7JO0gNDWvMf7og
wz05g7atu80akOoZEIPAJNNjtWoviJbrW4tO/RaG5jbk+v2cUy2PCRD6YGuD
zm2Sa3c0/nZ2nqU56Mqp8dAOxHjwO08rtVMA8UzSa26HpvJwESJtSOtGfwr2
A55i/oBC9ZPtClSPqG9wfPDCYvrEXdX+Imy+yCPqcTbb1XK3mf8OTowDz++M
vRPyJ9OindV3HIEtYJYxCSgLf84U2wP1qhGj7bG5oz9g8FASBBc2gzqguuFK
Da5vXTdjpkvF/hVSeRSt721WAVipAIyNbI/16M4AvWu5eInYXK6/j/Ry4Dlh
URufzBkweD5nMzlkH3GMqViitx4+Z7wv7Vf/gDQOdKNBHJzOf27s71ixL0WK
Q30JULx91HcqfXcyx7PwqIIsVd7PJRYeh6MHxeMAmNFmdW9wRe4SSNskMRmL
nmw3/VCcVs1jD5d1vvE4NH3CI8RR9MPb82PGiOgzcM2s/TKTNDbhkSozetY1
AUOpph0Heuw1XXAvZckz2hD4FMuDyI4+h7aTZh+00ek5yCNM7Sn7lF5pqDR1
0gc0KOaaDJCUi2hOeDpqQmYTc0TFitVqQVKSW7IJGZjHAmK/3Wwi/ObP0CJ+
YgTZkkFz+beTFUp+hScYGKt4gsDjZvy4zzEZfnrfVoGhw+Us4ANkqAzHCXBl
x7tEjQcc8KW8O1xCiTXMFj4shXlqL6xL+yE07K0+hnYxXOvL3bTskOt+67Um
wy0NERbjJbwpLYqMOSN9vseI5zkTLXGqp2Dm0rYiBslwXj4V7p5uzkBV0Itd
YTUlCh1qQT/0W6g9BEgd+L8dPsEG+fZqnd99NfKhIUnIg0uLU+YL8PDnrk7a
XZAkMEq/ByRG83j7R926FLhbn5Gh6b6IlkJmAtEvklcVdMXkxjYCa+5HBqXi
jnHyZ9vFANbkN04KFgovCP4Wr679on5Vy7FiU21WdA+I2l3oGdC5bRPuvT7d
5HumcYziHn4tjjvpiG04P2zQ1ofAoMt8to4C0JqUNpeJ5ou1W4gX1lvg90Gx
tVgq0U0ck5TGHV0OG0juYZqZ2XyVlk3azbPJqNJrkMRVZgHcEDKcYF+yMRgv
GwN86xWmEtbp8GAvljfS2GxxYG3qwgZw1B5xF3vBuYzlQp1KUAMwjxwbCBmN
7lkvfSC2plILiQErPCXSyRw2h3oo5ftLoMxZ/12RLtyFRIHwktm4ka64c37n
/sd/+pRxvgUxpZ37t5+h6eyzKbpVYTkBhhHTHoCFGo37vcJ00teuVdGGMeu7
ruhRkEOwHCNNGhPBc64A5l8Y9qsYowGxFr+xrImj04ciz0qvtFuFolKi7X4Q
zdj0oz/lPBI+OpKm5ZO9Qm99xAR9vAMlG0AdQkkloOAjgVfHi6ANz4SUNWgS
6KTK4SVINxcYtTIEwu2839i84x1EZyJB17PIq8VQsshgQ6ASzSFUbFoeOtGU
Gv7bBxVI+DMrldD6WIH7CAfKFaqLI68WTqS4E6qgQW94jQVW2mJwp/9CUN9c
1YyUIU2lmzGv3xA+qUlkMBhNmZYQPL2CCvpreJ5E/1ZmF3Po9rK+svjqSUqG
B2251THgVRwWhyeheAPh+4Cpeo3/m4SElnBidq6HAkzxbO7tB+OpSIgOrHIp
2Dlqs8KhHZCMiLymbCW1RDKc3BWhI2uxXIKFefkoTyxJW6ceHIq8elgur38Q
HjRTdRZIhferN9lkvoRXqtUAs109cSjs7aFzjs4629alfvFwZduZPmIncsNn
zID6LjrFAcR0NJAAYM15OQ3TRw86hX5h1nkP60DMuHNdrM0fi86kce3Jri72
7Ovu9ZpNT/pozc3vs6ZGyBuD+xEwlf/jqnv/NppXAKorbGkI40V1/fYlmuLR
yh2Qn9FXxKTi7SAdoBI/1EfhLHAdQVnfdSTVvV6OgqlJlsKcf4W3fIb/NN7F
sYtZ3zPnys2VMLRtlOxjuEW5bO0280o/TfxoFLqCiTWsy29340vE5fWkR2wM
V7JdTf++VZTtdC3A9AmnCV9nr8mBEo2aGjXW7GDZ31psOV6MdwI4errvIdWH
rlqU1jGW6trqRC+xc4Eo/bDfZTaTho1jFFfqWU4EuJ3dzjnN4hhWaFz7pdQz
pXSDoPUVv+ve/Vn8zXHxToRwmslBRdNu3hKvPKdhfMng3Do2mDaRimJsC39A
9TBpdh1iPHZ25EHpju981wLymHfybB8LHHJIQDfxD2DzXNBSm9aGSeynDLA/
l2CcHcqD5nz/8zvgEwF+kjPSpv4Dv0mhgTYWoQwqha9l0u0V2fN+FjTMRdyr
8KtmtZ2NAu5+sFp8eJaVKDsoZd1NO8dO7ae/oISaTpI9RilNjOPV1lN/3hWy
R1HUsK1C/oXm99TeCREw2B8pI20OUpW8Q6oDC/3e6I0In9IRiOo4YFJCNChS
QjdOgQ7bbRuLopZNu8mrxeE4ATvDn9R0b8J+wT/ZvpnfupUcUMvxz4jN1Iff
gRnTnfc7/Eu11WXh+9T4prOrtW2aQuM6RTgRqdOwHNk8ymu1sx7p+VB9UTpf
Cg7kITWj7t+XBXo5w0TXgDLqC8pRgc8MlE8EsuOX5FjW7AWlSXcH5vwyc/L/
OlZRMOSPiYFbiW5Q9a2h3Ejvq9MtJZLT9/QevE84dxRkoAOhgUplNk4Gg3C5
QnkBAaqRPmOpJ21nrO2rD3sovtDTpDzwesJYMR0ybkhf8zaZcY3TtYnhFS2a
07S5NmXAIBWqV35VhVrAgLOT6OkLteHW875+AS6zPPEvjcvCOHZGrpLPIsqX
vEZ6DS+CUfni6qGHXJ7x1S1eT1Xbt4LbwzSyeqcfOaPF93YcAMZIhBoc2dSj
AWrbuLDdlS5GWJ9t/rERGWFRWTFQhNFpmbesw5097l1xDMa7C7kosMrmAb6w
5yhuofTuV4nBrOmfcax22Ww/rivW6+rN8uFxRTfynF+dnHOS+r3sDIhIpCEV
TULWLFUuW4Co6Vyx6JguCTqAOMwCwO3YbPZck/43TZL/yJCs/KOW+fcJL7s6
F4K6oyo3V7RhVFy+rYzTUgNkpTpJgfwQigsOFZCOdaStwKh993u6wsgiyrtB
Zlf2VZukVFe7e6kuprCh0hIbTkIGvb9R37PjBog8WbPH6ro515gX8OTNYy+g
13QF9ovvkp1Qg8GOevwbJcr9vgJy6nXxNBWJloo//pVS8Kn74nUcuyQsp0YF
DqN5VGrov5cnQhKItoguVvvuBiQ6ijN27QVTBZIB/RBp3RbxjFs7z7iLy/a7
7B4kmBYFUAXsZg4js5vi973rDfPjqigW4hWJm15dTPwERYn3v05Fg8nMzxMM
TpvjK5Lb9lrQTAElsueX00oLGGSjoyaeILuR4VVm7gHyv7bdtFI8ZiKivrfD
Y4rJquT50+PMvf+1kg11nsg0MkIuogwB0o4H8z/2JHZrTUpQkS+CbJhT9axk
ZMmLbrDDTGmtTwIuj+2wpZcKxefLBk0SfBG6VQFn6EUlcT4yzJ/DFq2AwhcR
9WyOlwhy4TuMSopnjfxD8fbe8xPWrWD40yN7oBAf3wi4zE98liQG9qoXA9Kq
Pe0qZYQw80fdFdWsUVDYQXY2e4v44fT/6l7v0oHG9nmYi2Kidqk9l+4T8Ydm
pK+F0Oa11wNYh80Z0vEPcuSgo1yLx5AbwMc6q0ihUnO/xRDsUudaf/dILCRp
BD0g+H8iyaBHxe2ng2mBwjh6/Z5kTokqRz7qVoJBezXXftMYo1TyXQvntUKc
qnasiXjT3CB2iwbFU3eRnboVoeggnZ7svN0cZZ9jdhZHwmTv5P9B3UfUDPH7
4fgErjondSJIxE2ezQnZecfAPMeB2XZ5w5g71cEFLkZyscO4vRi9By+Vy4mO
UrIBxAmO2Lc4mxVsMXNZUfa52GWBAa+rF+tEjriSi42VC7/wtFJ79F/HLUe0
u6QXp5azynaK+uvXHf3mrwT6dxZ+T0gVpq91uzsyGrizOOVPw/6lm3xIsOSz
e+vTHhkv2ggrblgPVpUtx3sAC/Gz8roPpnjXrF3at3YTYWO2bV8vjia0cSIr
nZ+Wq0gaVMEgcfb4YD2/B3DtjBPdyGxTk76V2hHl81X50eBlOsZe4LYWBxPC
cSoSb4P/LprzsEblQ64572rc+zLoSGir4oscDUgcY2kDWr6u8aIobKEVH3c1
ve9Hp/lLYhAUzqjm3Ug85mMxzbmPBJ6f7BFvJPfGaz+QaWnIwVgdPKih3J3B
3qP5oBDkBCjtE4LE8XR1Zuoiuxxd5AepGLiknwBmqwgeBu39FdaVQONdb3L9
RYTdPXjs+rU6uS9uE4R7jxqx+u1M0iigHM9wxpmrT19WhxkRklowrKfW83R1
pjHUu1QBDPHNSRK5h83O2YZsPd+vSYwCFlBNCTJo+BmMQbbgddhkmdqvBhly
XVpI8ii1U5ZdfjQQ4C6bguZJTjXQP1Vz78CvmTtZ9H9UfX8uS8k9DhP141KI
8zE1OUt1rY3dcwGMNrfqOycoAIDrK+enmOHpQLeFOyupmBD54PgmrF7vriOj
h4g2KZt1Y+umrcX2MSNVo7mkC1WpWu5NsE1iNNVh7MeBfGhltMr32qHCEOca
U+SCPqBCdXuS8Zma426pAGYJmYBfk4AFSqYhwGm0MsiIklXTO85S9d/zTHiN
rluO19ueHoAf427xqP+giX5YEuKCW6fPuCukhYlfqG7BagUnph9MArumM9gP
0m5yUG8aPqlhmCpmWhPt3mTpov9FtNlvzkZRDWx7TvCfEQmWzafKVWyaiHHQ
2AAO6OsTL43+pfc3jDN8SfwWgV6uwqkxv7enUM2drydfAR6ef58BK6VVwQlC
36eFnl4xxfQ/fowP0oyQITij1Tky5BaAtO5jyyYZ2n7xZRw6+DuH9GYv1TNn
qSOX8R++RtafOfVzsay/i6pU0FbSJSqrZCDgNhE73otZLqBzMrcbRQnep00d
7Qm0XKRziZ2evX650XezZsll/ReSjh4d8+DjfWgPg1TtRnCKoMckHEKIY1V+
CPYr3zaBqkQCqIA2iapEC0XgWQRqg6R5eROoarWxidnpRiklPtD6e7ZcFbHY
ewljKOx+ZjwbHmY3Zo9G1SKU0rXE7ePctWxTCQqy3uBv8rOwbHDJpb3WnTHd
ZnsJ7iFgCx3Bfwt36utg0ZvHOdVxD7eapjOmd1rQEBsY9yBDMWaviM7GkFcD
j4aPfzWvdLWXeJ+mKSS1uiec9MbkaMSJ9TBOvGZ/Rkb5cqYdVomkvzc5vHwr
zkEkQp3ZRLvjBYKOd7hOrikbp0FrrYn9pZxnreng+iHlqFhF/VW/43y5xmji
f/TN2znWPmGyz6uAYqPzwt/EDY53pvQ+u6sM0VSTOZguIxx8TxiC8rB01WQm
aqQkVD/iFNrb6iEvlraayzL4OGN9J+wubp5rR60I+GA3R52wGYr+boqzYBxX
+Q2u7FbuOeqlWLpP6nPcsVu1vAIWn6ZIkYYNms/7JN13RKb6mhFO1S6wf21M
yoVAzrTaPsmvdyjkfXWq3XVF//6l4W91dik7YmHOv10kMQZadXjiA9fBbh91
9qbrTF8vaYyHn8zaFDR54s4j7vHO1sV8YMpMLfqiflBQav5sIZcoFDCjxDh1
0yFJ5JS7fsnUtf01Gc2AkvftQDvxNGbRRmYPJMWOc7obmKwEeqebRYsN+7Uy
dJSsMkjcBMYtqEm73Gr7vWUEwANfsKb8aYHd+QDEvqADTjSdhW5IAnzvwyhi
sfQUXkd0IT8D0QarzBs5CPbx3+8Yk1yQ5vRmGWwkEqaQ9gXkwnLVh/q4/HLR
GedQx2z+rLYg2q3i0RyEssBtHRirdysgooidwvsTHMovOjWccY2bk7DJrZOm
ttQ81UU+5AAqnZBsVVqhLVkxa7tHvNd3abfrcOP+9jC4PXwq341bRnAS0F0h
Pe8fG7qVmf8jCTjlIia+PC8D5InUM09f/EJ5yIOPoWN9FQHHzaG96o3wbhtk
zVKSM8B1+EKco70EoPVpC9f+BvLC644bT1pqc23f8SOjGCrQKwH0EY/DRJ9A
VYwo8WaRSPGoKCeHVSGu2WRdkakpwNGBg6PHW2e6+LvoKI1M7fLSWmSYLgnB
4+VY24v8XLT0DfnTvGPTWPsbhVNmYfmsyQyorgQjP/lDAyHsa/HSyLzoK152
v6x/g/OhE803qyNDDC720+OPXJ/WatLKtEkYC6fANxgeuriqk0m9Qi4wsdz9
x8m+NYFdtrqNe8nmAAQuUzTmpMWIVEt7ZVlGhI+0ZMLGl1GChBIoPSGZBlZB
XesBvDA95REeNPxwyah+E6Nner8bv50rW7WKKKIV96/WfbHB2JRIYmI0qJAf
TJLt8taMFzDloNu/9Ab8XwS0UEvnCdEjtjnmv9VpHJlShzTz4rPzL7nRJRPX
KFFKA1nYpo84XiIzhr/oQNsN5mDlMnxaWlA9D/0a2D0JTO5ediGKSIseHTJy
wcnMbEhCXzVcBRAnKKu6XuFSm4J4AYM2PtpjzAc3ESqB31LQfozj7BexnKW/
DaQKYHPuq8CEfqT7Wz+sy2aPsSTGiIb8zYGyJR386HlMV6AzhGlIW+5okeIv
wzHblAi8M+T5w+t1/HRBCuSd5V8h9rBp6fTZpUhGSvuKyFz/Kj0/3E7sUwRJ
EPg19qQD1K9XLuE7Md9TCtEI0AjH/+7b5d075zxIIjzaaQENRt1NZkkHv0F+
GbJbX4TeA5JdCHED/+z8IDKFobCJQwzFC6yivpi7Z/aG1Xhrhs8iN/OvHO17
zNCNlTzmYxuhwmpdlc1vDPdxEbWwvfOLZn4xvEkrL/Od0MzTDAOyKNRX+GUH
5YZDRCMEPudyesOlPFusJajf3uPUJIIqv2soJ1hxiDhIh4kfpAkAUDwP60OS
uf2aDUcVOwLy+lbAfz6Em7MLUtfrWE6SCczJ4si/AQMldQmId/vG/GZHpWbE
PfvedMesYIZKMLZLx6hAt+loAni+znzv+fGVJZMp5St3WXUjyvQmCfuCYN9u
0PK4RQkz5D4LTKm4J1lIwOG6dQ1hft8Id1hkyQMvSX0mmCcciOyqjRDRpJtV
ULaPFgyIn5YcoHw3GS+lVBzetMrFLqdTC6GuEZB5mDso9lL5eMXzUWse8HjC
lLH9UDQP0XU4GNfw0Ezmy8viSsZPh57/GBVpQ6u48JESoQkDNlfc+uwbqOOD
+WnTQx9r679NDaryX2b+L7tRBKtSF84dtr0lwyfWCux6lwoSncEt3CXAohzN
yJZ6LjoSGbJtL9YAMEUDoJbME6u0uhCDg9ud64zt5x/lgFPycp/kiG9xgsqB
/j5qMuBGs+eH7bk+f5Xhk9TbnV3u4rfyt1z9M/ibdORsL4NwjkhumzYPDM2F
W8g2QTm1PeUHmuoTBJd+NVwATMEKRF+a6UKZN9oQCV1gbAsMot8UHOls8w7c
SzUJQhfYFdAe9Qmg4YhvvT6H8IZcWyHwz6Mqcx2xXVzSmqQSaHlR29UkqCS3
snjhnQnsUPCNzx/m5Ss9P2FY014TsYyAgeF4fJC9r55/WM73kK2Vy7gPVH3u
sIogZ2lX2eAbPxpV0Z7aFOOLBklYBjGY0a5Ii/+/tuBoYgDB82yfPBW3DfB4
WAMNlZqPryQLfOsgkbMCgqbYEcqDA7mAL18DcL1f5eDQcfTiU5gvOpHRbUeG
pLwy/jHXisp8hQ0H9QfLk0dqE1LS1ip1+XhmooRNt0lZmpUvifYSZtW4lBFF
cRE4LcarfWw1PjjKwYmH8G+9+GcnQVOR3gZdLO1v9K0AQ0BCFp/CNocjJdv8
bLOTunUZlnxCW0z6JS30zwhKIKtuEC4/o1RguXYLnlWWTWlSzwmEN4A5zGo8
JcFbNwLFr2DKcwgKuHbFXE7Fdn79cAqkHMF+lJXUnI44IADZO/royhLGrNBD
YOPNUmizXhzTUc4jto5omkTvIk4TwimE7Ntgr5BrEl0coy8xv+7MgSvWdd1I
c21tO0xlOixdk5TgCMe/oQARqixmtdGMbKOBzNQUjXyekpcoyhJj8rlLmxrg
Fs0fDJHiJK4wEq8K/Kqv90Cy4S++Gyo+0GKW9cEigQm1LrbzQT3VWM7spEVh
qrVq5ChiuaQ8J7+xtPTCb6DGKVpjfFMe2fxh2Kd6FI5Ie4jSuuhIdMBaI0ys
kBBbdvtw8wJgQ9jg3LCm5IGAWRaU463orG8Zh+N2vl+6R/co8aeZfWqk27mI
Ypj7/e1Qe/ay9OTzIyfinDIhaT4OrPxamm93WvfatI9UFrPdjzQaguAYPG9S
lSNmlm1YyrYbJNu/G3+0qVhRbqnx7LPeOnWi9IVsozbbCJhC39rA5iY+OFml
gfd4Lomg0FmZ6/3uex13aCVEc0GiUFzHEPhF0ETCW1DBTGwNoGBTU7uFBbcU
HmCO2q2wSfeMNbnocXKbMXL2J2h8dins+/Ve1zLIvLiwJwc9V7ytErh0Cs+P
6uZwQ6KUnhlLHU+ws40zwaqqglNPvyyy7PcXrZS4iJRJ9xFIq8aCWz28psVq
6ZKBdFuXntjFBjwLtptTxLtXWBZCV5CGJiZbF/gZ3dhf5X3eBIX3WexN1sou
ifZ9xjmt1DzwPDSc8KzR78DjGfD1wf3TCVbFatFkhq2G7YQQitCImRZbCrvg
Ec94I7er0GDxMhAvrhrgMil24iIZFUUrwS/kBDWdOgHaP3ekXrZGXEQk6+RP
NBIFlD3PfJST5kWW0rQLQJwvkOAt+6kcn3+XpYnOM9SHQKQwCj96PdrTzCNy
SGLrJZUDZjctW7a12wXWRMeWPyb6qSXR2Bqas9uz74c0gCLFP6HPkby10qCP
a5Td4saqElEDGANzYwqD4wrMp3iC1rCT+oP1DLcfaqFkiROLCjEWIugsQK3q
F5gXlP2BheLbvYAbi3AKck1UDdT32ZSYQoiYdIbbuEwef8+Wf+jnkh2X8InO
uX/YVBamhCa5su2o/ZK++Y3Mby2B3sElgaRE19+lFIBpuu7M2Mg0fxx4bjI7
XsWN7CdVRgnK5Xuno+FJTouseljIz50SKAmFjWSgXTgopZY9neaP3dA7f7ti
v5cMo41blgNm7Ns6als95FxcF44b/gXXU5EKahEN2HorIIm8RUiAKbCusF2i
q4ho7J8eke3/RVsqVb7yjTwPrewIoOP9hUqLycKveSfjUuUSR+25VsXeJXmL
cId2xJJ8key9kAyTpCPkgX8x3WJck9x2Y1ULZmB3tGNL0R7Sz39qf6SqcDYH
Ym7SfaMq6cQgX0GBONdyj2Eruc6wPuyKSc/WpVkryuZGxkg7ZB/LvVw5KHK2
gh/nr11ID5lvsczS9nRBlwjaNY0MgtCnKUZK1LiZzHtFVs/rk8fYXKE9SB0i
WB9M2KGixuVZa2hSb87GSTNh3ppaq8Muovv9UB53nrXZ2nC9MWdwF7RFYnIt
gqKGYdxmyHuB73iVEvlbl3ExGnpRVYwRQNuJ3sAppqU5amepBrD/efxftELU
MDhYKjZaYHWju4qVGOnKAFyiLq9SlbUkERNcp+8Mnf7M4bMkax9SZUeEUCka
b+wd5iRypG4DwNInRE8CIvU3LumURfo1iSEwIOb977g1d2MYNV4ofOnnpr0O
dqNdh4cuKyVR+zBb7eC6W+2Tev67aRCHQqSCnel6Gi10wJ1V0NN/zMShVOpp
9e2h4ewcWF+OZz0f2Yw+mUT9WevK4t4XKjykFTaaWCO0VWLfxyCq7R8oGMnC
3Gz5C08NIegho6Uz6h3srAati1DNKRjMTp7AC1czLuFh4YdKPBVCRJ3VdI1l
qkXSiq58G9jl582oi2Z1HNATvCQoUBsQmTtglJN6fAtr00IcI6cCEFgCwJpo
yQdu/jgB8s6qOn0DeBZ7xsm4teKaZRLUa5d+2ZTnA32f+3bTlZtgDREOcYTh
bdoLB+eGC40T6zYr1qoemlf5010Pq99xJGWG1djFRH+e8Kb+IsZmqilFmKQr
w8O6wV8/uF69I6gO7P2QYNPhgt87UGeZb14TXC4fSqabD20U4Xe6fAleULKI
p7mibiUZrMOjbJwEl7KxBkiEcAIMIfzMcIyKIwypa0my99kNHpbqsff7U8oj
t/TcoI16JUBWpy2rCd+o4c1EJf0FpJmkt8wIkrdIDS7+mb9Fr5BM31sD1RsY
o1RN3fN00WMd6gmPLnvVmmTmLisH0gfvEfWwbcjch8MR+5o4JuAPpNUr2I9B
4uKkli6/+6H3BP0oYpobf6uy+1czFWMPtCOiQfPV1O4fTGl7qpI5V0qUo8hu
M45mHxBVXM5iTuGrgWmi9WbYSJdP90AskY6P9zKuLxOWTpUnfb15sZBAUwYY
ZRB3YH6Y3wU5IT4Tfz6YzINwKStt/8XMKDCau4j6wpuHV33nYZ7bfTxmEjog
jsLXkYp05OC69sdtT2o9YI0zAHBTgw4WyJ2zJDrmcgrfNphJgAaLXjOfHlkc
X77/e53S0zDBQYFSCBLiDdBbpzcPAKb0FJpGRFR47kQEyEMZv8p1vPzNugwc
zcq7ZR+sSAOj2xzghSiwH1lXeEqmkZABlesDzFleGeKvQQLPfxRQ3RXFvPLO
WBOIlqt/zxxocUgSH2YyIqD8bl3NWW1XuOr74j4C/r4T3PC0CQiNTuoC43No
XzZBLcFA9M43wbrTbJQXquPu+12+t8gRe85Stu8f3S13w66Qbx2ec7AR/d0d
LYM9kbyurZipVfJANs/ahJZnDLevY8hW45umSOZ9CQcLD+nJ0w2EOs+PUGPR
RbLktNwIXNwANJfy6DAYDZWIJYS9M8/62KPfzMCaxei9j9h6BIBfjEvFqLZ1
IDXv12VU4f7bg8mgXVwtC0v32vbR/aRFawFigaKHrgpQqwIDuFR5Gkoi+SR4
WG1bAesn6cNJR2g7v65TP7lCVXgCIcpLws+yEtlhtnEokDKhuO5n2ChoS0CL
nywP9qnPyt452gHCV40iRz63nrSXBwOtKhdQ5wlMVjReaAJmB0lVZTWMSvSH
digOn4WsZ9VaQXvjpfAi160ykKkQYnXRNhOjNp6xgC482BKXorVJg3MSTHa7
7kLmfz2xpJ66Ww0P1CF50fmI75w1csMsJn+9Awbwvt4UY4FOUdZu+LBcWHYH
A2o2fcQrgm116AhTxwGyfrKT5YQyXwZYbMDrGWXm4G6pL/8gyP7mFwNsqLwW
wu80yZz2pAoOpZWshv0EuL0qjWCdH5PMlF2NxgmsLVPPXJ9hfMYvRVjIqfHn
9IacP6i41zFFuc8v3nk8y4IIjdlC4UbYC3pufhGNJolNEpSYGNqSZDchXkrZ
HpVBo4C0BEGlTRVknFJ1LXQK6GEFTznu+LVf1Adx11a7oM9+O9RBTjhL8ap7
v0isFbDdzNW4KnK0aT6LOIsrosySx7ayqUxi2g9VRnFmgKxodCtdYKmvcG5n
muU0N0JXT4n9RNDO6Y99BoJjZdvpS8Z+HP+RUlcZc8MMRti631ZaIVgcRBr4
jeZ3ByGQHRR6U1bfIVmO+Cnp/xed7VhwB0erX8XhRBAH5WW518Gaaawvx6W+
llfT7ktqwivm2/Z9ITRgEf8Zqg2CTnBdwxsL6uwaOD04i2U5wmX//P66uIul
uOuP+i49oHNQ3ZDmrmq4HhnQRyRvDamI0MeO341su6ozUfbW4hE9GhM9PHzO
FIMIOSB8oXSVmxdOHg3M6xUI5bJQS8QMktR+Eqo6s4h3iJOhLttoWT7WaTV9
4/QeReBzEKVvkHr7uaNJO+ZG8nDB9xi+qPjjE0ywlsWDgqd44ke5HheSwije
IGnamfvRMXY1Ct+AH9WBHqjNr6UjB61LZzeZpZ0qe/CiuUnzBZGhKWB6MXlH
FjIKNGgfT6KnWlyVBAGaacSDdTV3mNsEGmrCW432WVgClRk/3wk9iAVcITvk
UmLvWU+X6B41MDURxbFQCERh2JYwPELT+BaQejQNa+GPL8gE9qwSAP3dLj2x
biAEqYOtMjtfHv9clX8SyjE1oYWhoeShyf97Ol4E68iVkV1AaT6t2NOvQQpG
5B5f32TIhzgXvC+SwA2JBTMrNPo9mhHCrgrmpmDr9z5uN+16wo49sCWvFpls
GFM5w7MuIVhFvthig1skIo6/B1Tt3QWhg1XTDvmxOpCwICsTaYUHg/S7xN8a
qJUGV8kOuT10yrHCeFXITG3KNSEnD/8DMYptPUUSmo2Ia5mckkcuYzkwDSbf
XKFD3S9gSxg6cqHAnQDB8kyyCNe2bHYomgi6I9/Cru5By6LgwFdekEWxRx9d
XCDXzTsaz022InkgdAWdgjuq2YzxV8kLsTyYnTKdszJjsu9IdHVRlseXhyiw
qkP/O+CIqEbB+18GiCabfcbh569pHsHs5X3eorrxfJbZsx+LVmkZO3ELvg0D
31qG+RHNOesBxCS1e4TInBy/ywT5fZfJgCLTqqjGdjb86FbUv0gmOfVnQgww
sPuYAlMKiRp/JoWJsl+l8r0J1ieaCD6KVCinoAI1jXhwON7gSMWMpslQakt/
8wdRz8qhO9I48zEhXXTtIrf4V99LXR6BkZLTYKQJI/RLroTLwtra9Q0YrOzx
SJndHGpEZWnNPVeyZnwHn5vXJGs1LZ7t3L5Dlxq+w2zMUtYQhapx0sYXEXjq
QI6Z42Rk+k3nRTtPupJLwgQTJ1LdTTdRfpnnBdEeigbYB7DzAs4G6JowdIJZ
W/nwz2oNPiZtDm7cZL731S8zYa4rlkiN48m5UZlcw47U4wVptCeMsEX2/0cT
by8QgMI1v8TkfnCSovfn9P9K64qa6mYfgAbSSEIYsJIaCHxAHAWB7q2asdBU
R+ta3QSdJCmvad12UVZz+ii91piDYVLVw2qo9eFE7Xxn8eM/wxvL9WbMQG23
AMoOYIGU3QxfuUTAg7hRaDLdtNiaf0b10HJEoNVYpwzOnLBJph1AkcaHRIbC
L0BTalFAaxOSqWRU4qe8O29h6GbIgYOPvErTsCOkBuKD2ruD2D5lNdwnRlo1
V2fyYdvL9njyGL7UhUWBb4stQIJkTolf/RhKhEviguPY0iDbhFtV06FJZxbk
Joi8bBfpDFgZ9QUYmK4iXCGkfhcTw7DZBf+88LUgalIcB6FvWR3FnAJZLTLO
toG7YEevrgN2ZLrJF/Uo2e4DAHxxV0TG7wnsfb2ZJgs8fS4N3Pl2Sj/CaeJU
U0khe3SVX6vvSmdgdhCksy7wnvq9RKXTlt+zePqiVNJQtDY3eY3SwkOru6Gu
rYTfwNJPrUkoCEzOzuYJmGFG0nFy+bt6C39zWx111dePgHLBAsTkYf5x1qlC
RIrRF4n50B0p/BOUg/RxdsGtTMpuQxNPKTDUYPTAw4TcetmO3aPh5mVBhKu3
u82/kN2snApJwlX8BfI+xD//FMqDH2ret9a0/OmaocZj1dSBlP4VVCadFceg
/zHLb2j0YiP8o9lMOXK4TwMFiVeZizT97589adujUGDtSO8kaU5wVu3jei/C
3n48n8Ias9O7FO+h13UYI8kIDPly/5OaNJ9Gz/ybrjXkSeD2CwArmCZKkFPG
h9BEdzcH/5qf9oz22mZiAJuZFPIM/jX0tKooc9ZYB3j1CJbsLc6nCwwO9dX+
W4oI2H6RQc9YQb878Ci72NimwLXldOjExsOpt9PdDuK+JSDfBYgzR+4//7IV
W7lNk+IMNw4DVNGt/BDklzSP6z4zeMBmNS0uzX1nDuMeX3kH+p5P9sXhwfNJ
HVUtXDo+hHlsjbywKubJRgqIk8W564YL+cpfyKOmwp12FMEjMR9bX+ud9YUG
TRAzLFZSn5gHm1cV+WXOc+Aq9DwQ975xk5djTUvKBHVIoyTz0DUoAJf8vZO6
LbXe0ZDCAaBydYmPKvTk+fVo0YvR7NmW5yIS+sRGN2rGfbu6HMiZtmseriy6
WLwtGPXAu+0+B7tkgggfsidfhcRHfE0065ecOmOXUCH03OT7oLxaAzvi7UTg
ClwS4+MmgxdVowD0qAtkJ58wDAqtdDdDcTBGOywtGZi03Tx8ntmI1ZK90sS4
kX8ozInugN6j8CjIjGqYVWrKQaZKNEHPwhKLoXTI3AyJhaD+S61xoVitn4yW
fB+AA5kt0cJTaxgLjIy9UbcgKGgeaSeewDQ63OnS3nyzylf+I6g5XorhTrYw
sWfMagXAVwMwcPUAC1HEuo8DunabwMsDBOn0zSQwz2Blk9dGp6ykoZ0hJ30I
wCLvs4+y4nvbYkRX0K0RJuS9hUS81AKkN3knivIoUNg+LniehXpkszEpIOAm
XghIKJdtwesi5UJLfavrhbkKbMpqbb8rO7ACOPrRvW7aZ+6+5u8Rj3kZmvxo
68LTPlNovCOswVNOd6HhvcYuKib6pJm5OLV7osKLTMtAu7jDiGf79pdDrzKf
2OqTkxWIXYXmUKOVt07eJmFq57FTOWl6NTcwtWbxzyBH8JKePg33SFtlGFQM
ykavKfF4bJOohEg2J1Uz+2xwV1a0Zw79WOcgenaFn2T230pJ2ShUO7UDpxWu
dWpn4uGV4qLvzlag63+6pNB6Vd2X7GvXq9ZG+haI689hS/So41mPcKVuDx94
GqcRP5RPGupFp5jvwsbOCaNyp0092w+/v838xNEzSNyApydRCzwU3e/vXa8m
9lWS7ru5Mp6t/A2MD4ytfAN8PPhU3of20UjQpH9uFmI8pwVN+Z5FRw5ysHD6
05gP6leDitVzu4zKPd4lluBUfKguuEPZQsuCod4buSmz8wgOlnPogwh2Y1xX
bQn77sGU+5j7VHq4c1FWunZfMhKah/ZDMNs41pKujkNT2EmHp3LraU4sQR/B
G1xU5xBCoz1RMj6skKGdHVvo6qiajnAQaro2aGezPckfE9oVJ/sf8LlJpW3a
ldqDkP7n515A+runa3DVSCivRi2F6s/PlqH7ZHxKQHW1HKQBfss3VFyOsaF5
acVmc8walW/OqJjDrxHnQ/JF4pCt7rSHzyASWjDR0gKCllwRBImgIisFhrbZ
ZyQqcd5MG1whnERuL0PoZvDCPQiuOCIU8ZhD4W3pACmYD5Qe0Iply31+/NsT
8kgx1bcB6UxfMxlF6tFSerlmrQP2NbJlimQsYY+eapN87omkb9S4/3jQmCaf
eUWj7cMVa9DtXDbBzgtIKNk4Y+yNOYVEsB3JgbaP3tUBpQgIlWDk6vztKqWZ
idKBkZ8W6IfINzRpqooaFQN+diJkk1XIKoJWuHfTkBdEB7SrcoSQYpKx1Hyp
NXl3QMIvgK8bIejVSbU4ZM8ZqTBX2vzimNvg/J64wQu1Mt4mWoMKtTrA7U0/
B+ax6W3DNxDUTOcQO7L1ZZ9dOQk1elQKCfSyKFxtHY1zjtH9XcPEfcq0tFDS
xUWZFawluYvSwfg7pPZn/YXyjMd9n1W5DJZ8PQta54vL2MgiHE5pXbDKJJDD
8EjIv4HO5D3hd6EtivZD6vSqxY0fiAVATAMXWrNTlcHQoe0+0iNIUK/N9aX/
9iSXUCHTE+XjGZiABwhDGG4/pji7TR5TGud5CpS86y7g7l2HeY/HkkoD5WPo
+8N+jhDm4bTXc814rKJuBba5P/+qj8iZp5y9+aMX3uEaK7sTzfHGbAYMF5KU
XmeuFSeypMJ+3TxsDoVub1E7+kjOKQ4ks7cK0BsdSxVtY2cFK/ZqueoQdhSx
xA3wjm3LYwIPfPRb6vQIugk9OXeThWA66mcsf5D+qgq1DO+59upWsE7Q/HOv
qqhx0tJC7l1p4Y/Mivw/qM8rkg403Qru3S6h4bQrZl64H8M5bMYy3qJkNPHZ
PS1uLzA/3kjgIHyTl6xmbjibUl5XGIcGxoaHOApj3tSiHeCBnSUWkTghzzk2
EUGqM/ch7O0OAn6VTFHVAJ0jH8SZMDFPl8YAfdXTCnI8N7cesipEnSScFFMP
o5Lhq8u1WM5lJ3mtwn7Gvg/P7uxe35q2ocP/A+t7KqcefuiLmbg+TsyeXOV6
hy+xUBrIph46J6r7r7LWsLBCf+EE17nI6lXblbT2PfCX92hvYfRbvtGvs32U
Z2Uew1lpuEMe2GgDCAxm5TsrNzWsdQ2jevU/fMtyoQ3HpvMNHX3Lg6RaK1V9
VCmqGJ0OliVgDXBhXqq8A61jpOoUYkKmGc7LWsXybDFzKh3xiu9iOovshv/i
+Nx5j00bglG3Z6Gd/VLvX07tNa3HqEvqTjevdZx2Rs204xOv3Yn/t2PZjUJR
xrRL7g5n2JXpaF/sG7je6HEwa9mOWtHT8cZKTa6pgOmHT83sd0Srwnq3Hb1S
0OqCix1n6cM6R2Mvx/cIp4tuGeUd7ec0KwYMMAN9/hI+GxqmpF8UTTvV5iqO
kgW20e0k8RXXv1X96V7CDTFzbC6Ql9ho/bZPtx6e+J8fasdJqjh9FDlKsCdO
qohBT7ho3lxZThhGbQbDC9HjJU6oNQ+tw5KCaoXQGHUvmdvJgaQoDcuyukuD
cbZLEyZZKvqxaSt0Ou/g/rUNz18gOBBtSnCzxtw0mB0kPghsb2oKxNYuIdye
1vsXvsxr5LIDiLedCm2AuSTGpEuAOM/k0m0iiFKmN5Jzydt2uQyZH/1W3Cpv
OFra10+qsTypNG8NQmIvC4i2UrCRGQ+C9yE03GvXNzGiLi+wA6S9rVuMHmJ2
5b9Ji6Yrza8cl6xndV5KzKrywEWyAU6l+jQQVlv71UyfAtvjZrRKCSw5ZdMQ
hIBbwqIarlSVEqkT2iV98MZCZQL3NX8yoIIl+0mJ5fgZDSfNuBBuBtWF+I8Z
yBz72wz1cHbzuQXufqHZhX2IrsDg1EJ/JWuSo9XXUqGkPvdHjso4fQCZqKeU
KQXFbLm1/HkdaX78roLDjTOq3Z3YWXV/O5kkWnUjrQ+GDHOb8g/l29w17pGI
/yamWIYt4ZoO6B5TJrK7PIev5WQVlztUDNjX35UZjszeckvqZv5hZpztvOBo
p+/qjvvRBYIYrl4Xp89SDfTy8e92eT+dMkq407aG58Wc2/Xb0SaHDozIi0Qp
kfjbsGk2VZK1er7dEr/4wa0IUeseqhKYXE4oo6GAa7Igpxbeiu6eijdpYKYQ
6KLEHE53glVS1hdYjx5UIwWLzLSNiE6LS4XbOjsZl9qt+4Z9DvOIB6Cse6p1
2QyL+zazxtnCYS2TUIJi59YH9QmyijtxBCRnbQTfJBclZMr9MEMKW+/zo3uG
0xPUumRmH7vwBH66AUFxLtmTfPsDWehFDe/OFHVjRjfXvGJ5qFNTX0cveQCT
YaqnIuIkVPMVQHXtlcTuMoWtHPBMw0Yj7b+sKKCkklt+H9HRo+ssxKe/uz28
FctZEKEnY08Zn4PmxSyL+89UckokrefYGc0antYwgoMDwX4j6pRpV3J+YOZC
6JuwZeo5kT7uPmykuCkhCcv4VCN2V0vsGaEbcVk3gnJNQ9J2HSckmT6g5ymN
MU7xq2521cnL20n3pDT048rM22kT+p/aWXhdyuPVUbvz6m/gbdpavAXrISik
284blNkLlK4uBTIqsk+aAZTwZY4L/EdO82eHPBYA0IE3gj8ExD41qJLEgDm4
cbIPOT+1u/3BVMwVPnRuzDezERAiOc4qZZDb4s/pCj159baOPpqF5FUv24vs
UD9L85PyMvBcM9UPI44txqog85Boa16o/l9e7rNjpDWmS3tQPiz8kV6JalOY
wSQK3H3jsEvaztWrT6F7PJ4YPyhg1kHrvDNn7YHytwAm4cQ=

`pragma protect end_protected
