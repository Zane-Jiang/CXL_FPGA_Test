// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YplKS9ny4DVBPGxlbgCL2IaPmd8rp5JHapwzn5/3fw2r+286fD2efeSlsEF5
K5U58I/8IaUUYYmg1fSUcZ57LLCQLYpwMQ5MvxWC0T4nPO0SbnIMtWPfB2hz
23bpC11z0k7yt2+gm5i/W5sswlsiBgfvrM+Vw/9Ns5wejxUtd+IUZgjfcSZ8
9/ivMUPxEs1ncc8Ix8eutJBT8B/RrD5rkBMpkJErJP8vfBrJi3GwAP2Vfl7z
0a611CbXEajlsZQFXu4SB9zIyoVI31GxAPwNyULDeTlUo7o6VsLhvka7BxCH
+Gf5RLYLgqKWOErHWnbG06xukIg2tmHXpKMb2wnBeA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hHII7VM3RUu3HBD4JQabw/8Ebfo9Kj0NP0g/m+RYhropIQT83Vz0gxZkC6GS
4kgvV5n9AQVkXmnp7Njv2dpaJ1wHTOZpZ3i17rD6pn1tiWb8iBTiqtaVOD7b
yUwaabPckq1WGYs8t2Un1crWrx2xLF1IP9KUoKmsny/39Zw+tPEwRoH5PqRZ
fV8IrTz9gMuk3gZ9SkiJ3Fmhnd/hcLy8iLieSA2MKvJiXCxOwzfxG6WiNwsD
8L86QPJjjaVkqQLi8czrqPmVSjxxKf8TJQlR/p5V3DT3GsSt7lWYIUBxBBfp
ObRFqhVUPLvGgiU2yjqkKfd4FhAPQtJp2Sz4FsQB/A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hdzrdv3SMA/IMo3AZtiOJYSH+EPMDPHgxBQ7akc9FZYscMPktbEVGw6o3/pG
N0kfc4G6avHMREE7XmmveKR7o2dIvSEYW0XCbzyqbqLLkACc1/M0Xs0U9OAw
zEDpWYxiJB4vtq6xzgJi+xr/yAG5hTctsz/lBi380m5KO3lZuRdFXMaNBRci
p8Fy9IoTrzt2xMaN8TZzVdmGkjukxGMKSGrweCpRNR0/pEm9D8BXeficIp/W
pbx1uGOKDLT5qtjSZgrAeF/zxM9VDWMlHfQsOE71I0uHV7J38OWgAqfnO6EJ
B3nRh+9XooG8BEVe8z3+fklcQ8bf3Co+W5b10d18WQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hL5hh18JlXJ56ux03y0lg+gSiGE7UY9xq75i16hGS9O2IawEkItQzNpJ9S3i
xKglUHEOWGkZECniZu8+VUvIcyChrkL5N6PAQ8RRZdJpXMwCLO6ehALfaiUi
CLNx5bgPWnI6UhgqrDwK91hIHpY6rSutDscGHaSKMLycEGRWBFE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LYRjwR6MMDqzXGecS3gi4eplz17hBOqPOD94+4wrnBjOKpAtu2y0HYfsdIgm
1chBDC0uLfW1RX8GT9707w+M7Xlx+8PgxniC8PdADKK4hdY6nAWNXTxquDJP
kaCfcn13+vUf8DvkPR2TyMv6kCCRPZPweRT1HiCuiLplw08UZb0FOwi65Zjg
5/SXWsbuBVttGWEcY9NBtbMqANue18IJqw9NcVmsa4MAfNKBMq37Hp6JiCn9
gGH6y6LsWHDxyAMKzb4BgkqqzpN7R28BcJOS44azBFn4+qtAm+JdVBd8ThnA
c0XiCzAfYJ2DTAoAjf/6nRnnn7PYGTFZS3sy2kSohEaHR7JjLbydHSUsS11L
EaAneSCxHIlIM4LCdpdvaMb+P7rFexpDbYpJ8yS7BIw+rK/ZYEAayxbRdkjp
5yrnzzDDmJV5eBS026HzKGTP/s/7uI2jHk3XiCmJKRHI+GOUdZFAF0oAfEeq
WYK7RGYjppiMYqz/wz0UZE1/9E76cICv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
j9aGhNYDowffSqc1roKZaG/r54wWAhNmMLOVch5duVTD/FYm/F4l2x7CC8sX
snGfIjVIiWHfkF4Qgr28hXAwImYr/RvV2XQ6kvYo2w/lMmp9yOstbRbeEUA6
iUiJaYOkSw3RR/2JvpX0TAKs2cyZZhk8pUPoFZn23Y9jYdlsDu0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LSYUr0g2lECcjThpy/4Jd49wdw6qaDP8VpyGfdf/xttOxOLaUQh2S/XCHC8X
vYGpa9MzSjNetbnuwWfv6B/zL3BYM3+Y2Hvs07Z5A+U6QmwfWg4TWsfgl7fr
tkFrOF12dFmNJWKioNRIbswJ3bXaHF/gKq+e+LoE1HjNiOIqzIk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16864)
`pragma protect data_block
/9ofhZzF4tNgBAm9po04sAXslAN9XJYh0A37vDC2uL1uUI/JUmeuFWTWqc9n
qydZKeYQ9z2IidYYAByEJfqNyRqeb90eG9S4muwsnbtQqK3rQtU8DeZ5TlWU
7H4M9asPlWEXp5wt8upsmODQff7FpvlwiOa4QDcy9g5vyC+lj24my9cv0GDA
g8r63NhzO8lhYxgTawPiC5vt/8Icv4RsTUDSAJlkIy5MAUxMJxY8s8N4NG81
Z2h4vwX8k4eFw+NE1NEuZxV/4tsJLhVAC6FL5sCvezEQmFI5FsDgIv4fjeJU
l2wnAE82u38nJPvAX01PRuA1z4LYza/mmz2acj96COaJUXIuY/tWv3mdsm6v
63+O9qWMlWduR6HZhfUL5LQ7oGp2qNyO9PvnJ/xxdvUlWD3K2Yw6ewxfRW+y
9XYO/ed9F449Dwwzvbt+0zashKdq8jfamkYolsk1Wl/U4fUPaSHAalan6ae0
3ExSFagLZHgpbnRDxiYFjEbN0H500nL0vG3zElwf6WaIqY4bSDsh9AeNUYwQ
cva1cvlgk1kQdlJXWn7aEAchkBfX72mMZ8Jt11rT5GXCiNhWXtEb4ktAwy8j
TKr+XvxaFTokxUBhhPJ7gaLyRJNR58bcEwI18xLmh66mk97t2l35Qa7Daf4y
nQy7qEqX+XEX2lvK0Ig9oGAnsN+HFN49WRUx7vo3zzUTrFtTDas7CmXTd+Co
BkMhDfayqVquDRqkpJiws/Zl5glmF3w4YPVTWq5+v2Ex+yx9hVNfdOFIZ8GX
m5cUlri1a9Ynt5YYv47N4zfLt6BWPrt2YrKO/adKojPvlA7F10hoj9LC08cG
dYVZEWQodQOPaa2I26SjdXlHyXfKqLiZQXke0wJjNvIPJp5vJA7ifPhhNrjG
SnL0uAGeS+z0uHtNFm68su9Hlt25OmOEpU7y8JPHJ6Lid5xpWZWeROzCVJHr
cgSGdbXyDCPRgSi76iLqFpr2LD8uQ6jf0Xg3FrQ6VVBJqVMXoYGgsp6xZc1G
4xXMmjDH9VlrboSs5OI/ItazjUMBAhWUgxMH6uOFsCHkaheFt58mb3Zpr3li
ccc7UQFLuo5RUl4xuVEgiC471miqP/qGnS/MSBoJMPeHndc3WUotGmXA5PLA
MXeitU1NZNbbwJwjYzkQzd9lWRuRm4Rzjg2wjHgQVa1FwJg+SRdXREypmsLM
fP0qCNEOfh0K9Cc6MZNRbVteaHqPJmr4Qe3DyDJB2xLeOmjWm5jX5H17SggA
DbWlRYcI3blzu/YRcjYGWaEU6TuTmJ2dEuV9/rGFbUkzQ2tDSuN5bH8YVsaS
NYfW9xILN//ECrHaNo09syeeJktsWiNb+98h6+dEvHEk11yKd9O5FX9jup45
AVrz6+PFid6acIaAL0Gzy4Wwi1yJaH5/sTiNUjdn/IBGS2Uv9wFR5oQ6ZsJk
JF0QcsE5bAv9HntOU8mF+TOeibBvOl4mgdST+ozH5yE70JcO/q1we33/t6z5
izo+yA0WPiYCKsyhWSMZf6zS+pV2CzcljPSQEJ++/6XGhqHKEXIMs2l6y+HU
Ma6MbS04IocHKk2goukXFlv63Zsl440Ts8ZDR+WAsIg64Ki4FQafQbGFlmHf
JRvQEMCbMy68gU3RLGxyCjGjXafWzddbMlfjev9k6bV4cSf+YNTobh/sL2Yl
i8qbARrgjzOdKb//GMFmVlycGJpBhDzhqctd0cZlnsLytt3lYwohI1TaggTq
Ogcw1L8Yz4biKSGC5qUJ1riprfMtEXDQ37MyR0vtLViLks/AK1+oLY68lapJ
RuyfgRUiM6Tpylj6Q7GM9OhrN+vgFHFu9mnuvvIF2zGc7B4PpVoIflBPB80G
ZR5nK7mvNB4wRpDLYV3xQBMDxyi41XsR4H8pPK+OAAf+zrjvm6q34YjVjd3i
/c/k4h5N05KOZY9b+jg3ajLHQ2bQ2DJgJMtNQghuHBEqviRIUxy3PTwmddoO
6T4RGnXCiNeBEHmeuJf/yABRlVyK1bgCh5bh5l8PHQn7nf1VfDUSJiu6Z8aP
SHVibC1034jJtmMIsmapTv9+vw24wyABfdpQujYTRIQJ89jELVIRL+OnQf01
1ARM/h+W1TLvhOMfBdnCyVhw+J4204yak5DW9U1j629IoinqLJzurXwo415X
wimVFhT3w182Q7GgSCcuFHOjSXAyudDFj/aJsio2v8AzAvT2CCPjEujsEHk1
wL+eEpj6m3F57hNZgSVCCguKmCPS2p+6iOLGom63pwxoe8ln6/X8JKGY+MiT
Ywjo9YiD7mrA0Sa/3LU9P8nv6PYqbq1vRKn0YIyUCLVnjm+mmzMlToFQG/5V
o5cWqMTQIPmQQtubBDd1U/8mIdECwOM740t48onjd3lUonDqnWOOO+2Brv+P
QaNfVEECNCcvGmyTQSFOf3FSI4ueiHmSi8CQ1XDQJNAI5nnjVmwz4SvxpKn4
QcOTveetm3TSCF4mtao1L324RJnDVf2kCTPW7qZAp+JmguzIpX1Or9pjv/C5
2mu3UmRjV4unFCgvqpZHgVzLVDWfPXMR08zB60qagLt4pU0zzMKAQRGtgrmy
mBVcCV9OEGF/dMxyYEhi4dRZK23RWw7d1GwasOdOu75nVTysu4v+4rCwNYwf
xw38JZp3+zqx2KX6e7nVnAIaT9rZg5iZkyxrJkKqDrhiaDyvDdjXNyRjegaA
UDYbEtq2bkEBnF2qwuL+B9K65+McQuWkXYOwUvSaLpvccK4zjC/O/geG8Cdp
or/iZKttW+5fDRHuidup7Gn6h5n4S6nlwuDmS16It5raNRNBgyH33z/YchgT
j5tom3uwIlWqLJYu6CBbgmy+DEbF+uR+Tk5TBYHO4ysJqNgdm/cAedeNMZF8
RgOYgWolCrI6pFhY+W6rgodTJ7YoZ/22wPLW+1+pb9E6y75WCfiXZpwCq3qc
2eT0l3kbszR8v8vCSG1AzAwnDWgwh8gKVZY+5+okFcMVVHAHnUMamZQ1LP/U
gzC0MfHrtZ4YgGeq2hxBPWv/JUDAk4UzYta/2lZ5Y/V9Ztu2oc+7hvsoiM/y
Dr+C/OIFAO1MnPXUoPFUOvdxJtaUJ0sS/rO5yFTcQyr2zJAjQRdCRyN1tN1Z
SF4/E0SglazwaZCo+is4+fDxIyIvE+AnmnWMlwWc+5RIA+Cu36knmatEOhBx
4YBIwZNnOjiybELI/sm5ZVO4yIVsXwmJ+jd68SNWsBK/dQrOu2lLhXcjyloy
dUOyPPOFoF17XTAvEvq8LBV8vJCeorr+RpaAPkrKfTm7jmqncHyKFOxj6imu
rJw5JnxMJpKiN/RKpuyAtsAkG9m71q8LV/gQN2eyI8EaMgVHDHAZiPXxsku/
nxPgMJ49sBsi6xjmjXF9xnURyflerQSaiQl5WwByJ14PKEdBfGO7E4rv4IPP
vPaTmIO7Uo0k133XK6eaDTvbB2FwEDKXjhDueI+KpPEFxDaw2y9HC4HmHtpw
luldwDcTnvtB6k8aQeqvrqOPCjKrWUODgYbmBl0Wh3GYlnuLDWybYNBlLQgG
fm/101DUjhGRvnR+W7ACUfTZAEpL/42wg7uI51FiySkvMZ4I3HIWp094Dtca
Z7bu+iH/TAwHPz0lq/VwrqSzaTyniUzQFyE6BipRE2xDMePAS3TF4CHIN0Dy
nlC463cMPhJiPW/z2adzOFT42nszmlQl5In9uadPirA2HgC3kvJxBxV0IP+R
hlc12ZBotSqKmV4OOw0CCO0E05FhFW7weQFKuftj0gtT6SbvHyaEHYZc4pWF
++kGk5E/cDKZn4vRQ0LGgV4M6GraLvC6hk6ESYuMDXEWjXFnwKuHqOznpd9m
6KfjocXoQYJC5+XF3890rrKRoa9FlFAGgsISJQr3Kd0RkqEw2pkw6fHP1+6i
7yqdsvjyj+fRay7u2Rvh6lFa815kcTvAnQFUrfTRV4yP1VtYfRCl+ayiNP2B
1DjyoTP8kGFoORd3SikILlyu/HxxD1X6D1nlo93GiqMlMA01K/twAnP2dfex
hwQ2ESGeTZQKPcSCS18HgnLl3TenMsgUvdfK5AKx7c3uDxv0Ws6PYT3hW0ZR
NhYgqZhgyfz566XItDRZYYdO156KRbUiKTi4IYSljXJN+CPA06KOmmo05sye
PUipctftDWZbt+/q6j+NXv2lBJ54Tmnw8KYFNRMUKyiJR2zHzZBrBhoco2Vn
UmXJpH/6B+jCXFJEuQMHAfEta3NE4LbGUIy0BLxuwek3DRlyKjdfj9qzSDcw
Cr+pedupDg/YhPYXSrTgXfPb6wBaSBD3Eg1tPT53bg8mVMPIJtwTeLsNPQpY
mU0RX6lE98MYsixCfrHJEJA1gOocCnuY2/DWBGBcvzjsevNQMou3L3a1+75P
YMMz3EXAVebkjhhmNvffosafghyr1w8HQcqcNklrvyELvteBC8IKdAOmBQJV
T6r41vJ4M2NHp17Oi+lhtzwiIyDa9kvKk8D4Cp71KeTaFA19/IivlT7eq13c
sDwr4rRP3Fz6Uu6J2ZV36KXfiwPUcNiY38R21Hyc8KR42vU6JGe6M/daVr1/
FLVeKuOBSqQRf1aGphCQJ/1Wl75x+kDN9lEb0lYyvYcnolXF7FZ+aiVRvZ4o
yqm7V2t7kcWSnfnftR35ClwrdQp2zzzEhQvRpqdQHob4SHJDO5G8OWje/CYz
6ODrGr8J1CyDCOYDu8RBWZb4K3b1keMEVwGLoxQjwLUpsIcIWML9OcEfhDdA
OusfNSLHeq06ZrREFKpp+hFIf1cIpp1NfI8/czRndUgDJslxgbScn37Hi5BI
zBmAu/rj/0XE7ITVYHlDsJG1R3czK529wUzzmWkBYfIE3FkX/KleLqRrHHLQ
GrUdJMWt2cCRLhOrD3C5HTXZ8lm97qgIiML+ALGxi5J+zcGEkFV44xeINFzu
g9n8rMlHfIxkrpcbqAvW1wXO8f8VKvz0kIkDs0UHR3KUr6cGHNA3Q4NZkrt6
ahReCxKfIdgrXVIq8VBP7BB/Ddp7onPDDCEbmOxfw+NSjEj6jPH1aQzDWw8R
ZCqDQS0bxI2si4FCny7SDzDz0reNlNaBSeUCFUzbO67r6PahLAobI5XLOzOB
NYinviHCz1lJspcpk/ZcTwPes8VVSFsTdD/Z1aKQZHgwA6FiG03rl6IrEq1P
YuVxdVfbeztF1iUcP+cJFidWuFnEbrgTFojiJ3ua/rOyvc/FHSv5vpZyFes8
RvU5TdtbR5TxrcnLlofY6ZfYbiuzZs/gIzeJSWWW5O6yYje7VJ2U5fWS3isA
monEgk8S9Lnl0UN3GFN/flT8tKsJNKWonwSnOidWOBBxidICrAF1dwfb1nwu
mxLAPZEEEUrEZk2XGZBjoHeAokmaiKa7tiPNyot0t0gBP3Mg/Wl3LBGagblK
thHTU8Z7nRRmUuVNZITQeIzetXHStYT/5I69ZqWUtW9KZh6BBsFeZIZSA6Li
bE0nzz2rVaodenTG96/9WXLDAGEImQotsoUXjG5XTqTs+qcioU2qr0nNGtRe
HB1lfjofCwHq9kBkPpXdNTXrQcrbaAvl2oSCbOQmpcbWY5Rz8aFid+hvGYRv
pBFOEcFWdHXRd21y8gZJGJKQHof8vePIa9T3lyVktNk7aPVEy75M5rEAs9Ae
GferTifB3/aB+00AXLtAojPJ9sZda04T6gMl4683Ix5o6COnZay6SAcIFryp
LCBo5PscU7xGQvco0XQQPpHOAitcx+09jK28viwYL0ooszOXYMGVqWcVSCjZ
u/1YFtmLAT1iFFZOszGxGrBs7BChDAR3b2/LVPe+qJVyHFn3cLmBeMjd5Plz
GP5RPqejsBBMzj179ulTpQva3I9HWEV2Ylphs/+9gbWvv2NX5Nz/dW12EdNG
gTD4mWg0wskZKkzQHm434dtIWrascMEVEhzEXtNt9HsAKaPL+HvPySvR4mr1
YMs/e0oX59jdzM3QRrykEt3Yjp8AEqRBU5m3Lt6L7CMRAt0BlKrGQOE+xHAK
L4Lguxo3UyzvDGpTTNW+OxzmoWvRqdZnigsx42t5c1nFC30OeY0cDqHblPlf
tct6CGDEQyKWFuD3b+FBl+hX7Y1YJguYTxOjrz9Ms1pT2hiXoPCQRr4ObnQR
hSEI1ujY7xzxLklZYJKyjANg7QxMWDIM7smxtsAdGmuzBbPmevTNFMbjBzMv
D1kOOoSDuKN0ith33XCCJrWZy6EXfT6AFxgIMml3zBcb4RAZXuZ2msBh0ljs
yZbdowl1Yt3iY8G8h7E0oFbcFOpREkeKy+TAdAt1B5xy6Eb5iyF9lyK8lWyr
qF5b+C2NO5yTG6tJzP6V282eVxWk2rZs3BxC2lfVWULH275pdExTabNlPUig
EP2dd7zHwp6vfFUjzGN5j84nl56ULxnLqlFRhg/h4f31ksEFgFu+qwUyeuKa
m8U+Geeuk6FiBzlGPZH1wQbNmfMRuktrGMEeLw4G1MLOTxKfXPpnofGMiFM8
RdpcSv4iPYZuJsdyKS9O7CnOPlNGwNaiMqx/ajArY55O4jXJjgTGYbzNwNHA
jgA1V2mMbmcNKzqoahXputehwyxZ1qLNZglFslOXrvgq/TBK5d/41LUHUvgD
UrRqkcO1LKMdJBpZW8jb3X67blZNcW/qCaSrGoE4sYHRFBsbv7LWhpXyTEft
8/83gthVm1zcy+9YLmw9iED3JL0ZbY/B6JOE0d28d1sGTFSQksl9pIvaM52e
gbI6Ke3d2ffLRJKlfvQulxUccXw+IFfyUPJDgkULu0vVZGpqmgXs3sAq7Z3p
Q3jU9pfnA4NtWdZbJBJBrnwxhM4K8p/tlab1K7lqDydFReHhHxeR5PTLk1hJ
3Dioz7RUTaos/3Xk7xxTlKarLnLpX87Ehy4Tdmg0EMFN5b3F3tPFaB9s17F/
N5oaGWQIVBCegYfV7rADRHGY+hx23O+AvsZq34xWcMoQZ4yJBZH967fLKSbK
wGG4iitztoontYHRSNklJw20QMnEB3yspMD4sLxNxHV8UpLzvbBFRmGWskj7
sXWCVz0AdFqbaAVLY4bfz6NNxnY3WlUHm/ToNWZnkwWT3BVeC0r0EmtYhmw4
JfNWdh5WF3xjpBuw+Hq73u7vzkVZr+smZB8JxHdPChnuyznBsnWXsKtbDjVy
g/c3wTHESi2T4ZSkSfdPWxqRmXhWSB95FtRs84F4nZP86iFX9fDSftaBu1i3
K6P956pAdgBuvYuI6N5aXd3o/pwEPIfUZBlBw9AKzD18UnLK2kwRM++d3zZQ
EiVdzbtnofFp8yc1ZlLg11vfrHizIDSmVpNR6tvVdAvlvysTsImqkksixr6R
lZYC/ZuYlhsV/8lIypbNsZu2pAf7j9/Hfj/CiE9mBvRKx7Uzqv/RDkDvYFX+
igLnmew+Mi7+DnFRSDJaVtkH89PZEZmWD0CDDI51Qb3QIh+S794BGYnNAeD4
pGPBkgd1okWHQWt9pML863BqU0Dsd0X80jyWXqwETO27ntrbq7tWHk/jfFOZ
XIhnzWAJaqFMLTzuaOl7cTelS60CJorQnzs9JRr6kGFS86rvf3xqpvTXZ9ms
/9n1v/TiBgJ/GBpB/v068T+7l3p8BtZE/qXOzDw3E97TZRli7xpJnXOjavT6
Ha+qjD3mkq7V/ZB8iFiKbSOsiiVrb1Rc3jwf/VJiZsvnOx7b4+uZzAAhB54L
zkJ8kME0rCjv+wEm7VcJbOEQu9BL58/VwbhSm5VNIsav7KDA6o2EhuLqalNM
T+QWPWQFo2f0mB5rtphLVUquHNs89YBiixm8i4EU0tJ6rbZC+FWIUXJDmOVy
oiEVUErkeNbSR5B+aHCXbQmpYMD1YhcNzxNDAOF0w/JaUfYhFchVAOhhxEcT
Zzu5kW3vpnoqSUfgBna5dQ4BVJbdWCwm9VQe/T25ueUPhlY5ciAtIgLbJ+2h
F0dZypVKREQ1I8tXI7uHOnogPch9x6Pu3NNbSCLN6WtfmR3oaaOibgqQnS13
O3n0GiKVjbeP4GOxKmeXCDhWDhGiuluMZc0573fKip554bGWH1BfPRYCGXNK
GpzqWYYOgEZ3Sn2/7HXkCrBfso+KgzPaZEV08lopz10v68ms9o5O2DB42GQf
O1J+iNG8MXwrXd9s72NWXG+doa4aCsXoAqcaEv5thWI4we/Gysra9L+3xUXT
/qCXIWQtrq3KDxWPBxXrRrh9pzS/nGuS8MHodps+kZXJPvbV976sMDXj/UN8
Taiwh85HBWdgAzUf0CVjm22FyM1/MhcBSJCPvuwrOTkhYVRYu2n77Dd6jdCF
/PaKQQxPTy42uaB65dEMwLxnd4B9wieCyh2uqT2P8c3PGcfwpAA6opmq9tOM
hbI+EgM0iYZ4lTYESz8r4o52j/dDwBUK/os3eOBJEXupwRJEeh6CWc0k/Jq2
J1Uunp4iy/bXR8ffHWyZuPNcT3raZLB2muFlXNCxOPYukG7xFCqk4/HEHrVz
JAm3cfvEDgMwzgOTxOBhFR7P2ACCK+xOjWyuqGL9ey6oYAsA+q7dQ04vFZ2h
b4QzS6XBm8pShvP7NPfNon8j0qj7R+Mwpl0AoBxsUvtF5fiGJUTsHtQGJ5r7
AaHVjn5i2DJWIpcPpb2AFgWT4crLQ7ljuVeaXGiXNMf9zXKeRoLiS2/rxGfD
WjcomvD+/ToHA4KjP2iNVr77gg8Mlg+XFB6oyySPOhbssibfIUgbhEpvFHm/
+gPuq78cf8G/ZndX+eahK1dbJp8wzTuG7CC/xEYH5xW1YOShPbWw1dL6tmtV
aUMwDiw4cep0ZRtzK6pN4l+utY/J86JeE+i6OJV1mvGWxy80wIm/h1x/JFoq
1jC9T8xEh8I8owM5BtqBb4SLfC28FIUhWbvs4sj1uevcjRDq2Zv8mafo0tgv
QK4uxg6MQeZVvxa9NqUNq66R4sn8JkSXSAzMx9ZKfQDjC1Rdh3xeO8QF44OV
jBGsE465+FO9m1+7/raI45NnWK0EampOgQi53rvJDlFnREB1HmMdi74bd72/
6NCZojZGCP8ZkXWiirEEQa/HB2/xaGu8Di6FnCSoa3gqb64RnEFYqTQMkpLC
oeJ6TEIVoajclec5XcoBPMF3rveDEBy87K7H4p7DuP+P0jw84RrPnpzD6fre
YbbV9XzoAppvJup6Owxc+xsMRPv6+48VEWXx8XjsP2FvqOkHOsSGZslwjsdm
AKperV8pUyCXsO/NSwFZZKdzB1wSga3/VTHmDvFS+b5ZgiS7JpqD6m6vV34g
NCDF7ux+R1IJsAPdhLCFBzOzIm2qUMl7pviUChUAzCWTXAh4Nrh0ByDALmaI
IJya1iaEyjwbVoVsL0s9NePZ7zYhEhk1AEAxujV7gI4GqU2SSeMxbFEuua0/
oq1G/Y/97zjDnJMXkIU3G4oQM30Xn5TNyil2NJaLKSojG7hHkPZdX3nJoP/t
Fa7YarrdEqIJ5GVdkq9cH/kvQxuu27rV9H49NokkGXoZ0+agwItMXnFHRFcP
ApgBGDLvVmkASzS65fen+BH2TMPhOs+3m73Q+1uI4Q3hxpF4Zl9tenS/wQI+
JZK6KLOhW1B9EtbT4f/sDzw2DL+2duD2bb4nS/xUGTPrBldU5FVrukl84Hkz
a8LA48PARhJCfE2ZO/KkK1HmTkm5pToIq5HqV38a/dlqQTfW+NZkGvM6UTzT
7dctc1mZkM1i719HMZ6F7M0k3/RCqD3xtz4MOJLviqnCBvPvg+j0oYNkYDdh
eTkeUdRoCgaUoXNyC/exNzMLvL3FougQUQmGfktlDyP+/Buyn9bRCjh3A0ut
SdZaakvzdrqBzLHyawniqI0JCRdRaM/i3TgNj0MNjHde0T+Sy7GnVbERQGHz
KsUR8t2iBIrkNFHNeDUM1qmWfTj9W8swCOK09I7aIVMW/KL5uKHLsl03aJlE
fJFj14pMkpCddViQg7Bhi39m6oTgYNUt1GAT9P1o3MwGR/l4RY4l3cbmYG0c
hdacTFT0YCvm9TYrkC+lUnWYSEBqxtJnueJdU6jsXXvBwCizKUABr7rM2FIy
Gj106uGvdDN61ydPxAEcIlphNlSQrtJ3O00aNBugJbI5U5op5vEB6uHgwVc9
1e02S67Z7fwlI2GRMuNGCvna9R+3DRDYjkCwbcwTiw6bzHgjdhDRKXiEyMFW
/ZFg3w23BKg9fKexwCYiJJn7SPcQGnKA6rljB9621Xc2ZrUx2nZI5mDeUdA1
rzLE9j/AMKgPlGIUvASAUUdQu5tFUDJhdVzX7Y2volWmZCEsHvz8DDaJrBpG
FSQISol2klueKw1xD13E2FVcNwgidfN3yTxmR9M/TLQZ8u8NHMnJvyo3yhLd
a+S4mAlhDxwQ6fCpFpijkynrlRp2q6DIU0x5pCV3ZLzPt5e04sYp26C1iXxL
0nYgaaYF5szsXz7zMhUqXP8nEt6USg/69LJzc7gQ0mi++E5RevrPTsYFSB/B
lcfjVtLfSDIVWJLGkGFhaJiDxNjF6HFpQbZaRGiPsAtItT3Y9nJpx3uhlroj
qINewxDvDtmNl2L4nV80owjaIjZWs1lIRAPFkCM1brUwuLazEDgYHAr0IFjF
uhfFWHFpA9U+qlcXeBAGURteNETDBavQ/YHNQwyIEXebs9HeFm0cot5jMiFH
s4pWKEzqjEJeU8qBfAm5Xf1l70cVHWygXDbfgyd3/fnr7aUahFisf4X08FeV
dOeHZcUHhTYs3ucLKFladQntgNfS3amLuRT3gBmf8zILyOKM1PBNurAlTULX
Rxj4enCpGlmqz9hf/pRGoTOqBjkQ+v/vbQMOEWG2U3/lWSRldvmYADv+QNaa
Aq/teHygMkryT2OE/eMdlMB1OcCTvRvNiArV7dPB6l9/ugo1bNGsdMd4PJzE
bi7sIqUS26pWp9wTXTwvRuHTXcMH0oPRBVlqUd3Om3w7WTAz4helWF/zF0+L
dooSn9MEXFRqkglkvEKbDYnJv5SrwvINETAwaGTpG7vJk6YM7WnS7aCcJ+V+
Kwg+2dHcjg4O5yyneIHgrAFxltZfsK9RWnrBfnHgnLxItVag7xKkILvMWg2U
4TMRRd1BAQk45m0KTaiOws/y5l/OupKbZoc+xOlnhnq7LrmbrkKTvgULt+YZ
kP4VEgQZi4cTN51YBXCPm9rnIY1mp3TQAqZwGOU6Jaahz++PemFI3Wo9A2PN
no9j5j5N0PksTTKwCtcX2T4qw4Qh977aOXf4jis8E51sodXEMv7ZbLBGw441
mV/08R5kG5ome1heR2pcgofT18zz5p0hSiAIJXT6nOP9394JhjperdHiQOqT
V6JVlm4H4UtjKQNuC0aEpRdNl4Tj4PrJFWTkdwNYc3PDGlxTotBxtN+dR3aL
lQu9yW7pelO+UnRQmObFmjb2QhgFKCoR7zr+C/SGu4c1vlAHPxICphj2m6bX
+2YRLSVvG6csezoFj3KJfIov1LdOJyppdTUA6Dba3aN5mu/+EyJMp0mrzo1z
RRdujlDCy9tL6+GcJIomRqO3Z/CJO06K+D4i3PUFWiP8aq2QcPXCrODZoYOZ
L0oqpzbnzUTw5XYhIYC+r/Sv4KOdqrVco9LBNmqzzWN96eJksm4Wrc/9XjLs
leuk7jKm2qMz6rt/H6DFUSk9HE3wDGa9JWHxM9O3ZwVZ8xR30mEIzjXGpY7E
rs0vsvXAtbDv1AOIPu3AxseDEEH6ri48f1HW0Iub91Ueyp3qgKURFofWzDje
LfUKQ1gchjXnEgyYMbROYFt+aE9K2Ti7en2gZ0ixHUJ+ITvjdX1XteQ6ukAg
rDw1Vmya7hLarhAsMFSRYTPgHJLaGL54z9gJU83hq3kqLPgrPQCpNiwXSYtC
IabaKUb3uRwRz3SG0e5e7CIVrO/+FGxC4QGGEpanFdFdQJ4HI9wZaEutAQ6G
8uKH6vd4gm8/bO8G4v3SAhecjZV7T1ZEd3JZUsag6IugFnYyKVzqxK2loPzZ
iMzDLdL4Gf9FN+/hq/vXqwyD9ZI/MeP24/VHy5EXt/15owtnKGsvME7QlFmi
NjT6jYR7lGcDgNtdgba+5+QrZrt5RXQcyLLuB9URwLus7xudR+YxW4e9COPn
qBTt+8jfZNh5/HEnO+dDbBItvrfM2eblXSObfbI+uqGDp9XDEtYxPlx6vmPw
OJaE4a8eC+q5hxb1ruEzTiL+DE7qORPb+MUoJuzwVO7+XmXH4pt+9MqeaqtJ
bCBZYGqCFLDsWxjYVFdiHgfNJfFRGvwNiffSXCz14RFFQ5LsULvyLiqhoqfx
yo8S+oEP7bEbSzQXAss/qVagt59LsV/qrSll74xcSn2hycbyX9aa7WYHmt0y
1ERgieA6JwbQ7B8kmEnbRw81I3M1M3VSKWWl8+0AYbbmrJoMlnfsmhtToPlo
+rWYSXrI4UKWc8dRLRfC4B+Wbm+WBTB2UUhFwcFdPZ/AxDJFv+xasz+eJRbd
bge0wtzKr1i/mkANC5hxwbwyRWZzEQlahTMS/ba4dr3Sb9AKeylDmB9icutU
4tUvBc5vQuUgGQJwKn/jeOQo7wFg8TgcGN/cn/5Nnk5vXvb1GbDn4YKYs9xf
2DaWs05eWo1r60rJqcYj2orQ8n7I0cOOPX91tKPmSwD/kqvbewQpmzFGPy26
kQpV7138JZFwwXN6GPpuMrIqO2xjk+TWQVeQ4Gc29GDSA4Wo9X6Sq8WgRyUO
IknXVjGQyuKEjR4GaZawmnd+JDTosY8+cx2LA9bYAKU78khZHdhxBH5LPVwE
0ypANSi+6GlER0rbLYYnh+uqE62SEh/d/NzuvN3zeZ4nYXa5vFhmK1ipp3Up
17GA16AXNfPY2wGuhFixt7qRB17I5lwCPTdNwCOOdXvXGglSvkpwC1nrBkcS
j4ct0kJxhGNrGa2iSp/UUxjO/DKNyioPFHeDJRPaSMOt0GGqjgfJicwEOy5b
yXCfbRE/N8/EAcMxE8DE9LNBYsiCrtY3IytNGEEQDQMO2+2BJn8L0Qzvv5qy
CqZPLzU7bj8lUKLTSCERNJbe2WRFbA484Z9qsxDJwS1Qf/8MXfkSxaBUzg1n
lG4Kuu93SEE62/k7TIyTcdgg3fa5kTJeaVf7/Z54FbyQi1bhVccYYmR9UzTM
qG4JkJmtTJsBqxUU1aE11zAXIMfvJa2oXFcGs3yiG9xGmgqBxoS7Ivpm/w6f
etLn0WEjwa1SQgqZEeAWZfofXp+A5Dibiqs28PsJlSqAmn+LPSSO5LcrK7PC
ct91jQO/eHxkv71yzI0/FuPVenLScXi0XLh3s6sxaA7JqVt5p00D2E+wCoF3
kjwg3FIioYLJsZVEp3IBlXfpBfBDsBPBIMXFePOnKwJ+wcPUcdwBCO3LoKl/
saO7VwU24XM+gmUN/andRVqKxkrjl2CYjNNDGvGy1EIdAM6HL/DLP2S+E4cN
S/I6iqi6mWVJ5AMmR7R/K1uYMfhaX4Iq8gCEASsEtQTJYriZsUJY4zOy4ByY
3yhn90dMhNhWMLjWVJ+y2bYSD1Y8rMGpY2jAlRKpp+53+Tu4Mw3IhqQCGsTu
k/enhx0EZJ8vtbJort6aw1qYnewPg/Rem+4E1fA9RIeYc3sfLM/+CTCheG4K
yd1a4A+GeDCyf3JrezmfkVSqPk4/ERAb0omEiGtAJHKrbpuoes6Uytxow1Bw
xiziQDTgRFxY2Fdbij4vU4bfjcH3M66Elm0o5T9ASIoW5LkS1ddCd7tLYgBO
psUfL5EJRfRo4MWl+EEPcQYeFJPGBW5wojSWgZNXW5uemKPX2OVPfq6sQQi3
2cDa7VHo1PApuHE0XFWYn/z5qq8pGNx4n7KJYpvPme7FHkZZdGMoJWPUvErv
kgnWkI3pYSZ9a2gInfJrBFX/zJ17Bwj/wc+j1v4f/zuASGl/I1WJOiKzTMU7
qPbv9ZCq5bx2WBw8rxVCht6UGwL8ZSsdVUixEGMm2Zm+RiRLa3IfT6+53Ds7
asREgMtNLGI5iSbipABlkxNbKTmkAzFL1bJ5khL77lnOHFDIJXgxXrR0N/ts
2OBmXBSBe3bNlVTfIrj1n2j8JIER3oYF2+PdtxKHcM7aHqPwEEf7+k++m8ah
KCJk7qAn+ZbESgXMS8N91Sl04cSTCmLmke8c+iNqWiULWdRr9fIRToNXiBEk
Qdy+fvm6m9sBEhRlb+9GrGb04oECa9nB36WPX6oWenSjFJVg1/upWM5C6Zmt
a38iamJKbQzqlYXeLGwlKOSqiUiNvH5DOwY3UdZ+0lORbbGhph0u2khDIZlv
Zvpb2QwFUbJA6NLYMI90ziTM7f+lWgUfm4kjh0neivKhNLPOUyxmAg0Kfn9v
Yp+XLlcZb2AnMRz8P5CZhbKQ10kjo/FyURykYjuzgFnfALpJtq3fzgtE1lpW
5OyiZNYbkQ3OyRMMRBeNkTdLgf9ydbI5RP53mmhLQlMAB+bfEdHmaSkKKndZ
eztNWtvK5vIW9l14nu6iEvMtn5tH09FJ+6Hx6tJsP5CNX29baj5qERFZsvcl
35e2t2+ezMs54wglvMYwLatDN5EfN2pZLcpPantI3VMo+VBRCV9w6AYz13qf
sqNNmYATfOyUJGSFIt+0EtD0v6rH10ro/avFMz9/pTuk1LQZIRJ0UaorPbnr
7d4PTV/DK04Wra5Pi/dO4IKhU8ZItw3SO7Djclxat06aTJMw3XNRQtg4X2Id
BjY4XsMUbW/ylCpvYEGVTWUe8wDrI01P+L+nGazC25OchGc9H62o/7d2DTQB
AOQA3aZEE+rpGlFjtKMUymXIQLQM684M4/hb+tj3g0VovP1oEN01JQRZyUUK
otaAqZimmo2+OOZO4OCjdSbko8lschEGyOwqzzZOLmmFcdxFpD8deNoxaZR0
mtW1Sp1njrHNCa5OQ1QaC8hv/XJEHOAJ4Mqlu0tyRepLrQ0qi+f6WXu+L8xp
KwzfYBrRF9Ku1A4ZCMnJlVDq4iBNHIyiVnF+EAXOx5XKSrFuNiDbP6mcWEBR
x3Fqovr5Cy3JpZISpECAwxaY6X6TtSwdKVkNXdeh5gy3xUia2FRBglgZU6Qa
Uo7BMlPfCZa7Kz9V7FuY8qSL1rCy4qZbD9StrcFU9kl70qmO24cWtar8uPaU
u5QIXB3SbcbdlbHIyTY2KFmNhuRpKHwPA8jYcoRFz7bhBbHRLhDR9b1s1M+O
Z7Uz5QsLJkAXFxCFnpR4B/dvgLD7rjjxBv0bDIi5n+MKQh3ekJJKha7CbDIu
WazbnPwZwc3SfwLgyZz4P1roQD2JYmNJkxFJDdK37o9U9ghSeiEINUQIVFR/
BE5ROvccjEfmel+5Xn8Nr9hvLDUCKuhHTmNLTtMCOsX5rb7EX0Z/y21kEuEz
j3uwb15KrSUn0FEj7nl76AVfvd9B5VEkLxF3US0Qlj3rpEqI0+cgkN47go2w
9Rbj0Ahb5+iMBoqym+bZ76veyM2W3lBNbEIEoMgzNKNmU91aOwqF07adIk0x
by2sQksehtjXoYz4dxF0mAIalpYPArJhlzRhr5WWioeWfTpsaIFlss4xouKp
ftH4EcGXcVODDHD6oTKcSmngYZuTNJXR0hAtQS0YksdaRj7KDvf3XUsIOz4O
iH1CYtn9h6bQL8mN9HuhUbBZxA6ubx3bdBugNUpRO/TIgCBGxjx/RWHh5CdF
A5JzdgyMdNWBJMwK3IVXKcTos7oxGa7iE8VUHWHCY2G+j0bh8jjfDRe7UQIl
N/OiwWj29Sj/kcI5ztfQR70fGHkJdaI6D++ka2PYi+8IfjVkdIVmvlqW6jky
NNIHcJE61W9qAM/QfFsl+rcpQHgEuX/atspVM3rHyypmQvp+8RcgFXQaMsBu
q8HMrHimTYeZYx9xGbzR6fN6kwLoZ1W9FJRcqNu3QBrTDtb0dwC6lsi55Wfs
Bph+btBoSUBTZGBzWgrZj+9wFf9Z59EOeEGbszmU0BWWq7wyc9NBSypZvSwD
BvSkkWPME574M+Hmkhyhtudi+JkOchrsmCdvznfpEKRtLNjRhfUHOquAz+/m
Y7v9LPVeUGTRj3ACASZo4zY/TZ+u5tr6lpRFcKgORV9X+UZvf72WBVhIZiaq
AQnu+dEZNMvVPnZp086vEEha1gRDmc1Q2YBc9qaUdK36rGx8FJcpNP8jlH1/
4CRV9AkHHdcTbxCVFIy+xwTNgo3P61SPFpbtBoMx7veXropC6oYrJrhVfeG8
4ufCnJQKjkIqwzmR2AmZNi2dVnQvN+0KQFxDOZ+WnuQ5N8yxc8mBhZV5CS1E
6Gb+3c0LEMRUtV6rUwQz3LW83SG1AKYStZLs8DzzBFvLBOmKGBvRvHLJcLs+
PgMRDbTQfpbnFW3r1l3pt/YxlyWJIok4FPy5oGbletNNZI/tL2yHR0/RtKPW
SkdHjJTCsdrnIYgSWgCQm3K0eZLeP7Tlkrv58CbnUQvLBRVBEqlp4h6jvGLW
RM0EHWdJAKzPmsPxNlNY0NwBMPIW1qPGUiF8Y1bQEpnJ3m/KMONZbWEPx6Wx
M08duLP4yzJ3ITwI4grWoC0CsUtkWDHARlPfk6N3Awv/ZXUf7Uqvukv4tlfS
T7G0YASODOTDbz/N1e8orjdw+uj9dhclbTxqJ3+Qh8Z4ToGx8LUpyO4XAcL5
ZaxwZ+mBUaVDgr9RszDPwOnPQjs7s+8wETUTGOb5Rkoii+U7dJ/hdapGTozH
2iuDLBOuEcQXjsdivQPX1dEZ1Hz4QA3m1ybXRuxuEncwG+Tm6haxcIOgizPh
mvQBS6mPB9eKL8Ozat5hZl0sXPHwM9lKFUrCDwn2VKSeDv6Xc6/6Mue113av
Pb0mSS/GyR+BTMLOvsJg484wH0yqyObJRYwcGmBMX+gfQSTqd1TpgXXRq95T
ncTAi09ReZXGIT+m1LjytzDW8yE+j9EXyLIG/SNazrV1fjD6dr9Bgah+kono
CDGunrvlqDoCvbjdXJZMfKuNgqb0VG/FApahOewIjnzbY+Drrj6cn805ezjs
DerLglG9HirrEnIEHOrE6Gp0uiH3FaCnoEpGEHQqrW8TuayPFI+XUsolOFHk
MvCMELHUN3ABpxYTxHF2227Otrsy5ElV6LlhRWRZPEAysinQUj65BJs1zqRw
EtMDkBfBlKgIPj4jepLIG2qDh9cAYdTDqwLdUw96V3Owu9KrV0H4haByzAil
u3rKOz9Q4bJ3AhCsbR/h/IyWAg6gdNI9o2ZzPXhPDvTvd5Bioi36+Ib1Uo0Q
2IoMs0JIfC2CCBIaK17Tm9BzFizql3JKhYItdGlwfJrEVvZuqeGCsFexTz+L
oAG1G0K9SiTVYMTCe2PhgRIdx+MrkF1tMreHEW+ZZsH+Xi4LgmZHiQy+cFi6
t2IsjOWwwa9r67w9PxxFwcRgwmSHo72RKkV5kExn18Ke81kylC71N7Nh7KF1
3A/zUWgoECGeofFRziDca/Q4lBA/bsJvlHrEj2+FyNq7FhOKLvq7scYFhu1s
Alqd393WhLod7tBuvpKj6AnGdMbisLLi3LtCiytLWupif0d7RgmntEE3odTA
h4MKBQ7FVi4e9VeA3BmuPu7rpteir7NSqayNPeG3kCUfAXfyiwrQXReFfhI4
4iasakCUff5L1pTjqLIfAlQt7cUs+qCp+ke7rxQXS09onqP31iF2GVVrRhUh
9TY1xldPTvyIihPibWgEw8l9NLsGEEMUznhfunJR8/mhIOWYr4jjRhP2VjO6
IOrxTB4FS85fM+x065CmXL3yXyOlBUFz9KXH3930c72nB5ZuircF+WP6ujz4
EYH2Qk1f0qvQ2y74b3TKRwhAT3rKS4yZC9GCcn5at+zvtSL43bJL2wQllPSs
y6+E2FCn7YC5XdO02Me6tdDvva1CraYQUw5Y0K6Ca4CEYsbfJvKVLy0Mhe+o
40C6W0tSvvVY5WmZVe2/Wj0skwDNse3wYY1b7opl3009S8RbFqzWLHGS2dt8
b/9XQWEgCnyPJXAIWl6pOauuxNWffRlzoqNPzMer4DlCfuNe6PeTzHlJZ/BD
hC8U+lFqRu2gIgyPIJW56zpo7Jm21MJxcNwSLCedgy2p0cILt/sJ6Qdj6z11
ml7Z02+WBS+mJiYfX/SrnWa9JzZBr3iBf/FtDAXBiTilklLhOXZAciQLHfs2
/xJjGbVKBlQgseg4Xc8KqQbysaAk8vheLxMlU6czxC0Lh5FB6hZcn9i8Psop
SFQGnu4hP8c8b5gjYxok8eTNaqJq+0IkPqq4pp3FMguptLWY6w8fA6JkW0hX
AbtsSzR6ujXADB6U3ujSLlGKiMyXloOzVtwwPV0cMf+L0uDAkPHp1nWBv0TE
K5jqfy0SL3EXXLC+dzbP6izu4GyZicDhpL7KKBWwfpwhaoecJ3MAj4p6Mqjm
DPn1VYxC8WSksKVv02Qyie5hesm55yXzYMcV+vryh3E+DCqzIOO+XhHs/V/8
6aZhcOraAHSihvCgQNVHGhfzjvcpLDHCAipTmcTfIVwAA8FLfOJg0u169TL+
CTeLNqHZ2pWhwEsXivu+xh3YVia7C1wFgKszsk9XGA8GSJbX0SE2tMBHZZGr
gMgCCgeOGCoTPmCkZ+KxcghrvVWzpNrjbp0qXrbHtEu6jEBt0cQZJeVSbCQV
JIeIamPA+mCdbPFYlIp0JUGpvLR1VFpc9CTRLZPR4KxyzE4Tp1E86IaBNJlj
WR/I+IxaXwxEpiJGepoYtPn67SpPhNMaty/rI3r5kC0yFNgkokhi/WI7qO8V
jJ9TSWIRR4ZDTvF8HqGLmp2uIctHgO3MKW+WK3O+lL6Dz5vBSCDbMg6quMLk
LGIiFocadPxPYerLI9xiw1sS2QxxsAzZplGPy7faTFXpGMHZaA75YqI+9HoO
1jukWIdbN+0wVM8EOb0aOsLJukjcqsbYk1ZG6lLbgJ4dVVBiqTVRrNvJcjTI
8DoPlliavEjWWHGymFyQo8nDOV7ncXpv6+CnVEu0/vzUID6jaDOxaRGxd755
JBgMFFZeHDOKaXyxDiOYcja0awRMZ8EeHObnqz0/L6//wmApF8pRTEeQcYr7
w0NIuR9Xy5J1gdzabW2TCMf1OYBNP8u/ZFRVAv90h+jdAyIWl+UqXRVezAVH
DGImdrFLcHJJJ958/GDwmQgW+4k4oTlv4qc/55Sy/2dhKiJ9zVm8zqjWqRyr
82Dm6IIVP+rAGzDziteotHaGG2Z6HixrA7SkmDd2kuGP8V3e45JrP0hEagsp
GGrsXRxRDjMzZEUz5JdU6gf1SylnwEoBIMyc+dwxWtr+gy0mAxE5U3DzZn0S
Q4nWhUL4ZnbfgqNDI49A7CEEYqk/4CVER+Vk3tvoBSTzYCxGglimgftR35sY
OlusqpXtwgOqTDVIXPCzPYNVdpQ7Qy1tTONWvxVNHKnPkvmXm/9wUVct8hzE
2CX3fQAA+aIYaJNstTGyoE4aDffezS6f8YWdLozmCn530TD3JUnK9BkC2Hod
6X/p2IsHI8EeBZ9TSdQwiW6SS9Lp3hoDHbJ6HFvmNzoZ5IXGnTiuhB+416Nc
qP53H2EKcqYcEIdmpj78qj/2T1Eq+h4AuTanDV/6QJqaUjN5/q/e0kdLujoG
TtK1X1leS24NjNhyEK9MjJk3N3vhtbugPK5JewLY5bSrjnNk9RIbXYAYEG0l
pGYKSIqhsaSjZcFFGre2If5EhZosFmNV1SKrJbvHKmzvkz5Z0jxraXn1VE4o
wIZMKUCJqLiWhF7cSR4cUi2kiEhauUVtJTy/HPvnb1OSf9sMp58YWCKItk50
I63M6S8xruN33ZgwGzxWRzhTzgEGx0jMPUWAc4gg2ySCduSTW0UhFPKk0oCf
AZeaqECxGkqluB4ncrhhWFSrV9eCT1YqzKeuTPQzfF80iyxRTMDMdjJwLq1Y
1IvNrqTd18L6z4JBWTjpQVgr5epxtO+olGSyuQTWmjHyLFuS3lm8/AHTLhH2
/r/semdKK/DrgDJ+DALgb7P5gKLChNIcFYVTULJHe0gP+xohGLoUyZES3oCL
ZqESo8C++9pZVEnSFzJ9g2kbhfIpFapKC4bzluG03Ot0hJaATy8mealqcTNW
q+HJi/VAuXClhpxOW1ZVOQw4uK0M8yYcrOK6ecl00NkWcAET2gt+Wll5fmLi
p2sAHzHCvo6SRcVLfj9TxxUbjQZMEa3o1CaPMDFJXiVKBYr2kJa98OVCZA8Z
qGsJrAwXkf+AOY8VpHfZx+ZIUyE/DzJc56DNayRIlyIDlfcDsFMGb+q1bkre
xJWpyvrsCpGPmG/NbEtw4XYgrM5yJVZ4Ad8TnLPrFNtoXNpjLYU/xsJ6V8ng
J9Zf/57NEQyPzn3WsDwHRyeLj+qvcFccskFsfbOFiUf6y3AzjULJ5MaBKgyV
VUOc9Q8iTX1m+OuaPYwnN3f/9gZCJqw1rtoSo7ep4S6zEr9Vuhjd1F8oVt6a
mT393RJb4fwEJEYDmUf2f7qX82DDmQoj/3c2JHqGqhvgyq9xBQomzkrzFNcG
atQWivjV9DLtiwEUO/4ZjdkSBmJYQz8M13BCNVOqgkTj6gGbC19/Inwu39pq
/YdMFlyEv0Fj6vcEK3Ifoyk8KUF0UysPTsDahZ3BdXMwHtKXe1qVk4B0+O2n
Gy0C9VBhvOaysu7PX0AgBJAL+Vjq7vvBSgf+jLhRayQT6R3mEGEUvdcl0e/i
40Gq11I0dTmOY1TugPoERg/DlEdjuIoElasN800lr31T1zl1zDhuxIJbse9c
rcMUJxbkGQbbSBs0i2eZWIzghKTXuVJTKqGYWNU4Zm6FuH8HxC9G5EYi6yaC
Kb5Z3rXYZHuDlnxV1+dWSNZqoNm+HAU+QlCTkUdXNIXuQrkE7WCWD9rEg3U9
M8Tw1dMdotWMQYpgAk7eZQzmfe6nMQES0ZoJg03JBdMVD151R08mVXfeLe7+
BJ1sM0cNBNbCBbNDLTJyuyLY6Uwn6N5w8KaYvmTLTwSNTY2uJ+8D61UapmSR
UrXuai9Uaa9nRAvxj51Sb7WfjQwmeLQa8ljkZwa0NXvzG521b3UKC1wRuCHh
0e7I/vHQwP7RepNkt/JXWK4knY/F4rxItwKHGblK1in3DNMiK8gYvJKgfVL5
yEDmtbtSqScO8kNy8zYXkUwYox6+UNMPQPsU2zKGYY5bmtXwzEzsIOTjpihZ
CHByRNhwLKjbUbhOwY+Vc/+Q0Sbw8T+SLYj/+pDbzchcc37pWCknYCh0bi+s
OXByOYbXAcqi9Zyh5wxF0lqyKITdzWflGfGk1JrBvqmwb2BapXEkD3GR0ys8
08jBXn441T980zn7SV3LiP1EmAzVVUKj3K6U2hEhutOH1OQX4YB+pbOaC5VI
Mh0fIK7FpvOqqzXzx/ftQ/ZYvkWBdFEpYMZV8PAcy/Hugfc8K3HP0TBf0VaF
bH5QfGm2ZgomuqUsEdX0/cVXIsTr1lcL+C+XYyIGC2Fjnv7hGALBWwSjIVws
GB86Dk2Ne61iMBB1H0MdnLF5z0Sqeg1WWtA7dni4nFbUqk9tCvwHvJXJSG9u
EjerM3Infhr5KHdAGxbZLd7I3WLW1clavt5OX3LQxGMJU0JUUWfOAJnike8z
E8I1aq7E1263xq9KZMcWkdIvmzwyP8YPWlXmdETBQNGXhR+FBdFmQUE8RJJ2
5s5ZHzCcRXhfd10IabsGY67OvmSiwq9ciZpUJ6QKQg4R6sGWxEKz+NMkdCXZ
YyKBPKaA6FjzuSca4pQxm4vdW0EQXgj7g+97QIiFnii+gSbaH2MVvoz65yhR
jwE/juXnEs6M+FdwbVgp58Jy/CaKFGTgtciCtz077rOzHOOs11qisEk1YFPl
3F6gufirIxsfaydMzIC6nmCV2IaMU4X/dxYnxwUQr99ATKYlO9nNYCixZIJP
HO/W+sdLXwLXGReexQfsxPW/lhqYplgIkAUTzLWueawzbGvnCwwKaI4eME/h
GucY7vBc+cnP2bbyI81dQOibmmlx1uLHkoQtJv+VAYHE4Vwb+yopQcEVoolF
rhLYCHN4aLMtot62dUdn3O9snsgM+YwIryU95oSFjzzspotoYjr+jCpCbBZP
vBoGS6E9CAoffc3RG9ZMwBiAOLYEd43BKF5blEOCitue8F3Gu/POsQfV0Sdv
b5LvnIsbck0jXk/iTe5yihsxZ4NPQS5ySIbxmd3197wOcpCJUUzh39v82jmo
JyHXUYJFJNQzKEVsS4PXt8ga0qZnwH6c/+Q6rE7pz/RRGJ+DinJu5JLOujNb
Ju3SoDuyXta+rNUHvLk2FtavBypaPpQ0hdKNLheI+gAlUf3ZrBpw4emvkG28
59ENEkXrhQBnD2TdmfPWl23rnP6Fl3bGx5/g4p3zlQkUtwT6zgmrRJHHYeQL
zFxQZVCEgDNiNC9GKOxGzVRBQxnJ/+hsRcn+AFxnYms6WIvUoO63IScBnV4D
TPnkzuqMC9KBHbtanDvUZxxYgXR38CexpuzsCh+uVPW9mF5Xl0Ivrqbt8xen
148hFs9AjA8FfMN6U2dw94phyVZzeYZFemBvCfBE520PIVvRUWMVwYGaOT6F
7Hu56U02brjEJazRlYEFd4ikG0lJWacM4+veGGJjMqu9Mg==

`pragma protect end_protected
