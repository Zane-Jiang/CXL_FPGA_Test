// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
c3/dLVnFG5iJerVHQaKm5ClMixYgpQ6WkRoG+eHe/I+AC/NgnUUxm6Nhm2lRfABn
K30Y97Wva7ypSAC/VqhasK9mERM9SG8KaAAozIcDntl9R9K4AeNmAusoX6LRUaKz
K9dEHe6vqTzrcP7Sz2PswwrcTp30j+iqyVJQh1FFFSo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 71936 )
`pragma protect data_block
2opqDnbzwibdae1pkKFEZisqIWW20Iebf/9BxwiSku/TeKtSmSJPTnatv7qpkSBt
wicZbC2b1UG9W/41XKfOBUkqFW52xAdlQ9GLF/zLZEfmIvPHxAIHE2sLbtxI4Lq3
2SJdav3FZjc441XMFfqprlxV8a55jY9YDuihGaHrW5YsDGQucrnGfqHu9XjXNE7b
0SjjXWEPnSt2f7Qt1UkzQC84RNIV18zAexABUemEdyAyNVdxdx3VMssV3WqlUxZf
Zut0Z5rhFn/HBH0A21wmdMqQhCTLPsTcOPb4aFv21LsZOJp2p4x9sirtKPRbIcqq
T6NDwBdcRuzfUWkVhYUS5jEVRKjZb0Pc7af542CBDopEZ60Cj7AOCuXgtODqDCiK
fQIdxiBK2GzPC5QDkBK/VJkiOS8n3yvY+BLgG4hsDRzOo1sGWlDxO/MnK3DCRFR8
nI7VTWH9JiigImrhzILkn+bpHp6XLclYReKinrO9rXV4778XaDsaszBNzQlxa40O
dAmz34AUjZ9Lasor+o0Uq/YGmb5koUb+5GV1wiYcclGq7CUsFdmrrA22vK/jIA6l
dGAkXyWElnp9Rpv5fSd1WCA36w+XuzjMVM2nB1Lota26WhbRO3LuKci9KLrunnxU
Pwl0jZpgcJncEZVbwGMDMvyzvEvKvuu69TlERsNhnZIN3/m9CTBlMJczfsTf8kWe
tPzBw4nRDjgBHMQNJiVJO/ki02U1qKFQxU31NrtRkSsGz6joEo563hrbrWgocMQK
H5Vyek88vggrT96dZotwishowhSC3ecdjTRUVEw9AEqriugBYPyAc/s18aaPus9E
6CMXwNMsC4q1xanEFloOZnHKzBH7O5XfMQ8Xg5Cd1g5o3EfLrUPxjRZdUsAgQaqp
Bv+eBy+tu59bYq9hybuIE2JJn4RnyFpqQZQLCtKFqOYGOa8Knf9c+4bk0AuZgAVQ
m2bbZnwJhYguB1hYTknBEVVmXpiTAFxz1a9SO70lA1hUURKOjY9sry1oG3yl+RGB
c4eRHVDe69qCFw2XYZ7KHoTG7ZEInczMhuRiIomSLEKdhPZhnryCADhvRFqEVqQF
x+wWpymqTEzM6I4U58ybXvwX/tUxxLvERx2NyRV0KIsoZ8NVjj9WEeTe21jPj9p7
Qoeue30JEGE4R00h0IacHTW/Tu9RnlDUs0a8XQkp/Rc8gpUwlcSCv93uRXa2KBsc
iCfdIro5Dybp1SDRvK074MWLbTOLlsW/SwbJPHXUTTHK397+IH5P2I4nVlJe7ja4
cMGeklxSvWUF0390qQocS+q6CXTF/EiezPOVGG/JZ7wa8gqdrzLn9JuRPXkipCez
2w2khlVg57CZBlbgT86OFLrOiQnyJMOHzi5taHLrMyUMsn3TQWeuXSpH82+2lrDx
lVhe2Dfodc/3KJT3Mq4GGGVyOQGkJ1pTnldyBUb2rTmoWgpjCudA+zQZiagQSCVk
GjqBgMR0S6LBGq6Z04Twjsg31v0pRGpmOOJ5xbAgVFgeL/6rWX8m2rnSZCpS02pn
Px1jIo2fRHkSSAOMi1ELFGUc4GdAPeQDta/FKr5aOhNAKTBNPTfBqi7rNV6Tb7xB
WytDO+sdBcnnQ1x6p0C5IXNI1IzoQMqMW+stbC76KIBjSZNEa342nx2nniLd34pr
HUcDk0OzxgUZpH1a+NFOD0yLaw7SiLuOYrgNXvwYphmnDubUqmVD4MUlmGotYhVU
FqBy79hXjmbxNd2Ib6NOvOPktngccmZcPLxoS1yS5tQz/YSUVDzBoyHfP0bi0mpP
dwJFeyK1ZeAxArDnDpEk/V4UauNHhYzVW1lGEfPfY1I3ghDBpCCbFabtn7VF5i2m
4wsW7Fjvw7hqHtVVTIC64wH5LqYJeUW52IOQxcF1NNEsAG2E4PfC/lOhSjJ1lERM
iJ8XT14J4VRvqrvpp5T5JyPFHWRUv+uWoAHOwvwKA9U/S2rtQED4KjnMCuk2J4dI
MRfXHf4dX+ahsJtvu5aMik7wzyXtV4M+a8Z7KB+l77trcSi+jzdqqsUCmlHqHkgd
3ERoBt7fpGlvI+Lt8vucfN8PhwRXKv4vANzQ9pKZH7KsiwjrSitLioC58HTzi3AC
R9v6CSDucF0wpaSg0qsFzvCeKJnGZ5XxEOFK05v4qwr409+WTTp5/SmCl0i6CHRy
ZZREM6wZF/WVVbXTmPxaGhnN3Vf/Unv5SEwPeeaJXfigfDZY2wyp35Ty8rSWrBlI
JSh9BsWzWqnapPvfCLZU8lXCDqmHPyl0oJZAKTck5UJaLCsU//BhiIQEtfkOayyy
r80Ho8Hqh+Tv3ltGadQKCmKuW17dBaKI5BBxWJGIowcYn1+vcVYv6gT01m3QqTED
LSBoggHec7XDrAh7iOsJu26clGK5MVTjg0OH3pjYUDf2sTOTGHI7LKGf/8J6Mko5
lD/GdqipLCzV8GD0dHRmWX+5+HE8ri9cbWO+pJ1TXaaL5bHGTp7hR+IPTJYwPnJ0
Kb3gWJR4bYHlG4AMtZUG11ve29/iNDrUkiPYTA279GZVAMI/TLF2yvVHPTD4VXas
Nk5kxQyxqBEb3UTDZMawPYp/8jcAwGnvmJPDUWnYrprJp8awKwPtBIcaMZ2/fRg+
xAbtZdzapBxpwPu8UDaQumhsKJapyALza09c8s12E4gNWcTGKsWhbTk18d0jhwN4
B7Id76G9+o5+cP/B8bdPTsAwO9CaxtEIKvRsjbGvlww9TiUKnvdyhRnk+xt0BJRv
0M1fmHeqycK3wgjOLpeOY151rR+UnKdrL3mEtP+DA/tidlqZfF7D2g6FN7hIphGl
EzSuF4hX8AfVxMsGE7EqYps9KAUouwTDqAs9CiloJEUGCIaL1MSqV/agYf0IV9Hb
NWZ9WDGoV+ZezIBIPgQHAyAcp/QH9T0lKj/T5DWdxy4mGF4h+w5X6QHJhoYsW2eE
RWI+yd7DCzR8U2KzWNQU4XEwts5FEKghlAFC7w9iMBJXHUXKIz6mS2rr4v1H1FY7
+htgq/fAY6JJPBLLzoygxJsMCxiobS6fJ8yGSRIE1nQGpJnXcCp3TCvefnFly4gO
JtBslPMmBaO03Jmimy1YdHrL0JM9l2yE/BKhdd2Hhee8cMWhAX2rZGLA3jJgLCc2
BHR4sUmJSYi1d/u89/gZieC6XKVtd1D+8Hebr/mHCBs8DehPiYxAOsZR2C+UJ8Qc
evaVuniloJMDGXoucvlvLB3OD3Hrd3LbALdLi8I7cYDzqH3oithKGQkQ6GXkn+I3
/uSAUEvVuWRCBl8TCIRfFWxOJmuldnHwgznbQkdu57TD9ZCnSgf++NAZ1kX1i6aa
Ai00WK7QZD0qG784PKTqzrSe7TsYvOit88pw+bWdgOSg8dbs6VbCyZMr3+xCldtG
JMNtCn/FvUKdxTtMN+ZLqtfMEpGuNCdmdU1ljl9h2kxb1WVBVdpSCx+JmNLOJBfp
nBor+ZFak1gE1CMag1OK6fJZLrg49sBc7iyqK8d28a3Gg5EWppjbPMr5J+mlOvsa
u82ohvNSj98i0gut83RTn2rIvM3plrX0twgN1jkwD3osyaQM1woBAy/8o/4n3Ubh
ERm5oQHFIbCNcNHc4EQJBXVr+KxH4vEgE/AJHr9MARVaA1Tw6gpbiX7E6E0DLMg5
tENLYWKV+pUwD5b3hrvIR1nSius+DrgaOyj0jjUk76NS0b7kNb8bm1Z3pG4eHPT1
G+1c/M03VGAxdHWWbnziIpQ2IsrpcmLj0Y8QCeQN3si/jZNUwmemSxhAFCvpkRxR
rrw9XF8QobmnOX+o+4cCY7AOLDjkNZntp/yG1D0sHBGfqO6MkjBcntTmnm3EJD6j
U9hDaR7WSvuMrLdF8kgwEq8Z0BV3XuRTNjxskB35Bw1TEOatgohstvr7CdLAHDj1
LFC6KURVuQllXGV+uUgX78RaW51sVHNfoXhvpgFq+2LHopqGd4a+j7FdnGd9If/o
FRx/gs9O5STRDbB6vzWDJlPoEwQjwIhTmd8tzroufQqnaKXciqo3hFgystwUcQHf
nDeFdqxTjyi8LxFWD36jrDRBlyAqO4nlzVjkjF5+Om1MYf3RzOHJYPP3Vg0upWkC
KO4DFU0vZDszRtOah0hpMKPkfpCmR88LSgqiCEC7bBvE+zG5R5TvXVdwXtwzzgiZ
Y82Wssywerbp8N/mJIgHjwb5uoeqRiEAmbbkITh4xwLIfPhWcBmoqqhO4FfIj8va
i0zxnrodIvL3SI8+XLuIdyMzGyLVjnkxVPiYpRw/W9+cCMGO/DMaHdq1vAZa+FX5
waw05NGta/wCZA7ZlM4VDEQiDNAajuCkzLu6Crf51XfE/fjisOmkDBasa1Akjg1m
MspV3vsOwl6HxBv515gc6+egfsynR/xjVz8Mw/C633Gu5v3eXIBdk9acty4P8cI/
W15p4pMbW7h465omhb8VL01q+4jL8YEfvfhrW3vqS6mWh2EYansoLl0FZ/NJ1DyM
6E9XXLnAa8H1vXdTwh5WRIC3JghAgvcGghf6aq/DUcP8AmeNr5lBiUtauwpyOIJz
zkbOC6QtqJRTSFe3rr4tv2FWtZ6Ucgt7/9wIvrH+Xk8vTdbmHFhJcSfcGw3AkQYe
MLC6CxXbyedPZW3lia+eYfyA3+it3yAgo+Cv+gQyu7ptsYpDwzaBi1/t6fCGIzbN
YIDoU3JJnOKva9IJw1NiqnklGmHPiXJzoTRa6neVZf/2W+84cTQFZGBOXj3UL/WQ
cm/ECF527Fot/9DgQSe5fjhKMSjFAOdkxaU+5/GkW6f5TBFXqzJk/b4JaWOXXYyf
fzeHTyLR34cSD1H+zEnHtE9q4ISvavg45WtNjgMR7J/gog2HNdKrnk0kcSLctbKC
/yF2J889/KMCJiXlsoRGjTG18qUhvl68080f5JoH4+9hA6cU9i0VgXMgYUO/eHjc
417+kbH/6gOt8w2cp9Y+c9n0/xWGwn9I+4FduD0LD24DGZmBQoLZoQXvoP47cptY
2v6yhMLhhDUuzvvwidq56tpTLT8dnQ3Couo+m5x2VmkFm6b+01cD1fM7TExqP2sS
JsRQfJObUSd1tak8C1INjG2EqwR59qx2HZ3e1ggVN+LqNJGNXQ5hmpmC50ro7tFv
Z6zqsFfm41aZlM+FhGjm4kV4JwgjjQnm3Bw26hI98GLxEbaAw2XElWjMNWUD+rsv
/M2eJ23IC/pE/Ik+KzgtLjSYHdrC72yL3Kpr6ThlB8wxqLqpaGjqhnc7ysukQxN/
+pX1rJQ4a3h1efHZABsz5z9d4TYfyF34GqMYGWQ5YjhdvhumoHbTXOYq7i7qAsfR
GowGPRVQ2vK2jTb5J2M4PeryrQh+ojB0Q/n1eEHLCsD2WJKZP4KXzV5z4etgHv7s
JMzO0AJMJTnxtXMikbB346KYKMngUMMkPjZ6GA4fmRoe7PSt2Az+ixumE0gg/l0E
B3phREmEcmBbefuy1+vJmoaDA9ETsW0eHO4rulLTWDG3OhZDNqMdVNzme+BZUCuP
XZVsjeaMcZC08sxLyz3z4yxus5JO5XEj3wBCH53JZLtPenrcUi3/bbAq7F/K8a4R
+O+AzWgDi3FjUpFzA1oP5oX4b07ASoObYVMN03Er1clCoNsrg2i8PRrLTioe1BsR
2MsZ2zZdtDsM/6rK598l+KQTrT6J/JAYgFemZRr+xkS+UABtb+TY3X1q00ygw+Wr
u7DTR0hfgpbdPaph7El4yVI8oh1h50NsMwbqqvb8iJN8QNww4hMoUdakYl2Od0u4
MemwEVrykT4olTYDHHFC7P7ui5sqSofxhN6nS10edqN+6fzZ+53uyfR+9RCWFR3w
41jkwkloHvmeO0znHwSlOSXhjXcyzmrDB61bKKYmQLjur2TuUXO6FX/TKoHsLmrb
vFrayNKlA33O6WWT6OdyHy9w6kT8OWWcur7rcfGkJ/ig4qIqqiLJ+Fg8YaUqO7zF
WNvJE4pOXnfl/aSzpgOgUylQDAREYKRO28NPKq+YWbcuM3f04WqsBwKrzGWbS9sF
cASBLmCmM8iX/PjovyjixQ9GaDeY1Gu0jknXXiJOQB+FmEf63I3SakfHDYsObWDU
BYCV9z97TJGp+B0NLQQt8anDJUEI4g/frwDWgnRwJPAOIFgAqW5WKpyAGA2QyX3m
nOPZSfPIp75tDn4OKGEW1GHwzvDFiqVmHwE95BbIAv658SwH2wxmcYwy3wDBiHeS
H+J38YrIX/ClV/+yaXZOBa5gWQB1r7QkkW/VyMj/CKP2kFO8MLE4m9burn6Z1v1+
PZ2f18e8GhpGE4FdoyB/eNOcV9d5SWVMtsVMzXqIxJbzgrAdIS3ynH4Oj/ouh0Oj
QotHAZ8298ZL8CFCYwu92PC9AvyGB0lKho2PHszMqrWlzJr1EdeeGnNQg5A8mPnj
KpW5Khe+vulS3JyBlGDDWJJtLu4PAmVexJQWhrr6YgUWz+hXzy9C52aK1eu5J0qj
A33PeLF4HEoK8RGRfJRfHjWDNahfzTyzR6yffF4JZFJBfAGUe9nRCw50euzr/MFw
tQTKX+p97yeM0U/M2QjvY81fKoxcuScnQzg02RH93vJULa1UoNEhoM9Con0pu4jp
LlkqWEPA29NSuiF66fT2CKOu1hji9KPAnv+VTrSH+P7TLY7GiGFSRteTi+D7LOBE
cBIO/pykxhJ01zUGqqZHmpMmbxYkKzTy/piwFJBPlnnzFTmREb8Ld4+b2x5rLJHq
4Vuyj0ShP/P6wnRhDwuTsGNiGdhmHQhfqLPufiZfAMUwNHehgpkYUQclRjl9SXx8
SsSRkX/KbDsKlXaVHxUyWtid3rX/vLsN6ExusslMo8Hm1SnK2XzNi/8wqApRFUK9
GkIsc9J+7f7Pa6Vu9R3si33yTRiA1ceeEqMLjxENNsnrbbQ6B8M2RvD34BaD52uC
dG7b/dSDkuE3vSEQm1pEgib3vEE9ISvsjLEuQ82mj+ejhZbf0ULpbxOB/ZmVpbKE
Jz5DQE8DDuAEzpoA8Vzs9quvhRqONW2zEovBKhN7qqonMVXi0FTmkPwnsFLEmA9l
fyKKyG+MTEbyqOeifC3PyuDvag8saeDoGZPwp2w0bU1jTRAXVxAoE4TEY04I1RUx
hwIk5P8leeSQpNakw/xRtaM2FpWssqbiCE5Uqone2Eude9mgNsZxs/VkG0C1lSy0
WSTbVCbvbnZEZLA23ccMGq7My6vg1D+3MTBgbEeeZlNQd/i+nY7hGN/AnL4OROvU
gTsbKJFaJ/ZbHaUdsZpNXq4Cq9VLJVh6VP5Ce0jO6V1yjR36BCwDMJKvW6Ub7OsU
azdwk0f0sj/C3zv4L2cs8Jdy102zPdDNB5OcHF3LuueLr5k4iVfHbqUhb1LeHQRz
vW+caJk9ZGy7WJ7yhYCCJfrxo+1jIyYleOA2qkvBg8GPJwEOIHuV3J35/hYL7Xbp
nZfMdritww9/owQ7+M8J1Za10f6L7DSbdtxhvssfY2lCIDMwtmUb2BWWbN1dzF1m
D49IEnfVJ5tm6an0O4pvdOV1j+UWDQKdZjQ5/Ebv0Hpo8Uvovdruv8GyOMyk6nNu
PN7IUv7+q90XoGesIe1K/6B8vTEGt7yUWKYqU141Mw/zK0fGhk0HPu3R15uHDHJO
7hbMAnicPe5TXo/SRBG6Zycmlnqj1w1b5mYb/ANSjy7hzd3itueB7ydP+cV6YCv8
FwnhqGq8JYHCfuupewHyQ+T5jouWAZ1+kCGrnFQpptjI89PYZmzSL8JlPfnWu48K
XjaxIaPZ+5M39g4pywFCnGHJI7T5sfvQ3wSbRI+b+4tMMRmTTctlo1+cyrojldu9
NDWQXUUUIm2mKRLIxQUphOtXd8Ffc/N7VkO1lZ/A2KBXFutZxytkY9Vt8Y7tRs4a
yw4m8nLLozweuBoV6Le0P7vdZxuYpzmLVa4Aj2uRyzPokWx3UjnBeCMeO+ZeT+1r
SjjfM2aBMBdMzYNm3dIMPvbgV3rhjA5MOPtzc9dKl9P1vo8MEXd5uSB1iX/6/4DY
sIzZrKTOlMGtgraLsvWHsPdnHeWyVoTqN3woo9Fj29IL2VJuZJ6BkWApO2OOXk5I
fVQLvuoF58RMXSlwFl/zCVleOx6+V0kG1lDFYk7XeqbASaWj/VRGbGiXSFw8YVg9
otsIKidzi0t+EewmDz+i+60Hvta5ROfPq5tNHMs1tWdIWsH2Hns+k7IyrWA1mPtw
TbOHug1EHzMoshcM413y+YMChpWb2gWrIMn3gqiukVD8oJiWeUew1kfnyVEBsxFm
lCVDhEp2M9LKaeQEneTyE5PKHxWv5kANNsyfLpoE8Wj0MYUZHVZHuLVeFft5yAMk
6fMmg0WTJHrZCMBilEkYv+3oB8QABVsTJ9Zj1Z379ksLMX2Dxja11cByH9GHksWV
Wwj78gNNqdM3Y8jb/MbIu8SKnuskTw3kv5+cjjOLrvamnLJV7u+rJcrZra9ha1vI
PmBEKcR0YYAGQa89eZxWtEi8fyDQR7uKUrPlY8RD4ElEQapFcTpxT02rhqvBtGLI
+QsPBIlLDBJh52/sAEJjqCxjo+IEInhUV8/jSbrRkVd1Y4XpPL6IsKKZ7lx20n5/
Dmg9vb/3oAmOLVZ4ZAcqVgNwPG3sWxydR0ZZNVwQBQlQQKiDexoqzZhx+HbMeRyk
FUk5ybndPkfgH7M1b0EOjBc480XPcfm+EDf8sotO4IIhwuJWJKW6dhSneDNuJAiQ
cQyBHIwrfqol/QbcBpd2eICM9GVnk1tq69tiQM1cMOlEzSduN6DiIwfUPGQJ20xT
bLuY41E300bIRaOwHaXmAyA5B5M5luX5RDQdV/5jKtmZgUYSfbhbirQbMj5LKx+c
Yj1WGKT1uN0j0cHj1R9Zy82WdDxoH2YS8ksoShSzRdy0vtSHCvlv3gzkkDxB1AAr
CqVDopwNILUU4tcr9S62oOxFu8kG77gqAFFxFpdXljW21f4Nb/3y716lnLpGFKMx
K0rRNMrGiH7CeFU4q0ZRQu5wnpMGQ7HshbXFD54jld5UnN8U+NZKz5WBwilctkZh
LGbgK2HqiQoVSMRINH2OkPBPdlIRhweRWIcZdk5Ocxux1aXv8DYsx2VarMDHYQB1
lzIZqonFheOW4C55DxaWfwXnCZg4zBbHrQe2r87fCchzw2yosj3hEqhlM5OsnZUF
ISCBFOu/jr4de7zbJDZ8fZCROqjTg3P5RW38y5UJdqRM0E4Z2LlSM4Q8YMIvGJtF
uYUG5MgxhFH7F8FKsrGFRJPr1t8qsQHrwUtufvtls1hLZvwW4g2mK34XSzWBsesM
ivoiPSb3sVk0PKEQp7f1d8buRVuydqqJgXJCBtPZVZh/PGzVlXUidYaQW+7MLV0Q
mht8q+qjDn5NO0crc+u7ReTvRk/aecqiiw0xrNBhyrTfzphHbyrcwcF9FRNtXdqD
uQCvrtnaaDb81xDLADa8Vi0J34nnIRl8t+B0O+DIegErvpI0n+Jy5FnvaTws1XzA
gS/mJaucIaw3sED9gGOVh2IV2R+LATBKxHretPTaKHDj0c0nFFfCBJsszFQWnn//
EGtBBW6RJtGjcSQJ2LRG2udVcwY3I3DQlDCLrobujwdqHyXeDgRqiPJfG/Rz9aB0
qjUaNiBaslIqtlEVj5jY6B5IhZUiRusvK0h+GMrxNka+npF0lC0xmLPx/rELtgjl
OB0hEKH4oY0mN7EZm9/XZLuuA8FHZvXuc8k0nBhGi2fADUx3vQOlXL+gUO18uQiD
zQXclq6jY35CJQwkx+mu4VTVhTSobaj97FwAVAeO97qtem/tAewXGQr0vyhXzLmh
97PQrsh/Idu9Niki7/zP2DG2XV1u/TOXqAkz76wLjMACjVLJJ54xJEuQAOTvFpEv
z5pQvZDY5KCVpqTznXglfiwXsFaELOwi6+mkqLkOpE22qHYZPWDozToRV02vdOHY
wbDxZF3p6qqXT64mPJ4qFRxTnWOuTNMAFlb10WFtzP2e6CBmnFh8SOC0bhmG51sG
dg2xEK+gfdq8YqEb372S9sqjinBM2hY6KKk3WqOPeVPDddgc0blqXRinHJF7s35w
0h55jIYPDuiVO6VQ/HTA9lzYdAQZku0DT/XBkjXGztkm2gfgFDFaXMBpMGhexIts
R0PuDYyg5aOIUITx/ZpJgjYzpI9fMMZPkHzf+8x7w1SH1qiwA0mtjjEARlM/bZuz
BiG5Wpc79CTyeQS2TC6J/l0+4vwyRzaiGMW5tmIzAc8h/+mKXGjGsXx/SHPfCtg1
Vzc/1m2X4pK8nfmaCN6YEV+SEsP+TvEYO/cOrdjFrWjHra0DYVaOwbzaTEuwtzsu
aGWogRzbYeBDoBhmFqNGVkAGr3wq3sNGSk179tyAb/lD+S5Sm8oPu/eUT+fHPJz8
+hC1DhMycYM2iQoILDVfWK6M0GdlBcgB0giSq6l01Zl6DNurNVsnKC0yryNNVbSW
IqjUJCz5WyUwUr8IrltH+fUKsyx8RCHNWfNroEvR/3ovxoaq+aGckM+a5GeV+kQ6
qmIwhLwxXLSkft1/rLvSKQJe/FptwhEoLeTbkncmih9ECq69T6y7ItTQ4LMtRFdd
1f5ClWapvBiBwCpSFR9xxIBiN0tMfdCiYcxYTCpTV5GHBlxQvrCVzYwyUQZWcsLP
1ra5dCD7hLiJuKBAeZr/SKX6j1xJYru+MVcnhmIPC8y5FYGaqfXMwchWAPCH4jeq
H8x+UJZ0gn8GMX+Z925S15t3dhZ3vvOW4RmDBEqbt3MQRwN2g1ho37CusUD7RCF9
7vNGoztA49rfORpKBD+U/Dujs77D/j6BdGMu/ptSb4lcljRpf3sOVNOxtjG6LqDl
zAP5/oeBN7UyeNx73wQZIY6WBe1KVlEIBF3Pa8X3P8W4gbOIEw4N47E3LUBr1bhd
SPJTQlYP3izr5u9ro8X1mvFzS0Jrhm4yI1cFR/oBOeQCHZouieE+v8uVvTBkd/1D
MhyZ6SNESGa+FJ/AOZNLMFOHvZgvZjjfyAE2J6Ce7Wh8DnYNkYJP5frg6eT7yERY
Es2d18m5QS86DTz4kVTK5no8A33JMLIcUKPLd6b2xD/ppHk9abQVXVGrJLXNU2N8
4QH7MEqh2fVNgLD/5iEvnQCBJMq7kgEhcX91FdA0sun578Q0JXHFHrAHh+eBSbPz
BRaRg/im/HRSsbR2QrBx6L5h5Pgo3qdBzw5RIjXqaTDzme9b22BEWXLHlqOJ/g+8
jLx559eCaghJ9PA07QyPFDY+r3ReePolgF4WABuLMiDzmogGDC0UhsFca2fLxJR4
U8ZVOp1Lq7LI+JOuSGrW25FMZNwVK3lXL0zwKBsluotEepEZyJYt9qQEBWLhdTif
o82qrqxs0btId3uHWbWBv/FPPw7wWf26suqlAnVuSaTMwBjBsk5Y+Su8sgEnnmC3
+Ki16oT1d5NXyhl3UC5zblxQL1n2C8iaBqjM6xO3osaD8x816cgKbPy0RKFafK7D
vLR4MUxDDm0ch/FS39+QATKMLk97YTu4dThd442Fyeh990KkxyEGSGfy/l/P78AF
+QkJ4l9nYobNi02QfZqrvPkfWreIImpnlOKcPAg7UW9NUjgNlK+Caf+Gim/S2fyL
PEVYTU4foxU64R51kgGapDV/0og9Dx6bVtKcHfTDpXUU79Dir070TGlq2CnAnz24
us/87fCDeH9au1coV+Zi/maMYfDgH4PzVmKMzajoI2EBQmEvvQn9Jr6QK8lkM9co
9OhRZcZ/bjqkdKbZOr3JL/70Vw0EZwsEeZrHX5/yaTP3jazQhyzPBiG4nHJVihg2
h/6gbxuJBV6Q6afiOQPdvy4lBSCLs7c6I/8gDmbDClHwQr8CJWwgTAPcnkEf0ACG
GpWcc7FZyBSp2m8/xOXgkUqf7tnXb6xRRHLr5WyYWqyTFE3r5fNuxDaPNOfIxnkQ
cE7mPHmrNMZnTL87DQ4+Z7IrxWXWRiHPwaQJB1J5fmFHMFjtjlGXS6nYX4tjyJSm
RKRWxsOpMWrtIa5+W3K7nntjPcrdELmsQ6SWs+dk2CLi9we0o8SYqa+MUvmThgVB
ND4e7Kr8M235wH0Iy7Ke+9bbkaTAOqavYZdWiETAPujPOJP9YX3OXNxJAYCfzS6/
YPwbW/W/DlzPnC7LZ/C1A6WQOFRxvUb6y2gNtHBlIwGdjPX1MeTtNYc3CrfEyrFZ
qk0twlSHlUtsJcPErWCYU4WfljKBzFXw57wZxEa2hMKMyv9ec0GXZoEGzkOnM33j
1JADEUUbuvZKitJpc3lTao+Dg/GmcayZocJotUA+WNebFJ4rT3exNZf8sKsIdS7C
4b5oICAtY3Kgrcif2QM2bX9X8keof5j3Ph3vhg1eLvR+H4arFKRzDH2cHKZA5/rY
zk08PsRrMnoaiYHa4ojtZsz47sZFYCZzrXvQ60hl1BoWAMbEjQxSv+N8hO6lB68I
MJ8RVKhh3wn8A1lDZLy2MMwn7IHMoaxnICrNyPtHRyC+EitJEmhnTQAd3/EdzydL
q7gADgF5uV9wSX1O7O5a/dODqunLTM8RUb+Vh9diKBsYH9Li4dX+oDIqTGcOVEU0
SDbyZm59niAp+MsSk4Oq39yUK3TCOgFpu1aa47g8mjAmUjkUJHOeS9QxKkqb04oE
NQF45xhE7mMMpHphSkawoMfZDYxakiNdv4QdIegZ5K+QDziIp81zud9oyBSPZcTb
uvLNlfvjK5fk+76IP23vru60dHlFsu32uCvzTjDnQI4Ge/t8pkXG5FD4YoU6mg0c
OuJqaF6ubO/Tkcq7Go/UvoPKtNMnENSSvSyA4dEhBM1svJZsD5oAo6JLOkqYLNkV
PNJnDrFT+aDhLDnnxHfMQyeEs3Ig+qyTi2125NEObdTm/W/XjCdUkZrDlu0tVbCV
c+rbgOAL8l5Rs1bq9M7IhztftoRQyB15Ly0p/wfXVadwxw/0kKV86+FDsJVZJHbo
J5eaLZ0/Y5p4pjIDaJ8UaBeE8M3nV6cqlZ9qe4+JOukFOp/Uwqe91erb1qkCFZE/
MLTFd6WMoSGgz/itTWa0eUOOG5nm5V9Ska3AB+YUgkd3ZcAD6sIJCLUZizCZ8LKM
F5VnzOhdOKj7x8gWk7dKfm2Km45zduUk30sOc+KWfa8gYab7vEj9Sziq4NmxujwL
1Qql9U3kXKLqVWlY1SuZDuXmRsYLG3KewjMBC0baMS/U9gMPYKXz76dUtRnwGSW4
eHwzv+jC1ITU7uMKeZ4RLks0Eo3oypZL/dDx0NK3R+to2Eo8zlUSPjIpbgvosiXM
pN1N1ce+3U42FFSbQ5wCjLFWQb+0hdjEEHugEyNiP/x9G/CSDBSLl9v42olRar8R
Al4BufPUmEbVv65FEhHt1s5MhB3o7/su5hOfPJX1WxKbWlSg1QkvDDDdFxJ4yucz
CwMLmEkUHlogvJajSBgJYlqSDpbIun0ljhcF1Lvi6B/G/WVKkpiPY/Vj/Y0crFvY
/KqRKgTbqtry47cymC4jmXYBCeZ3Q8JmtCnW9w2LSoqSma7Anyyiv58RUuw1LAfn
xq165Qn66N/IeOl79Rmx1476Dvkf1MZZlohBxyjWSloRQjdtt9R+HzyMy1kFfpBO
7/OFPrZ9ePZAMgiQ9krBnOZgExsFtX/gLjBrfIe/OPPlMCgd5eO01dzmOhBAmGIA
lb0Zl3tVa0iflzd1mCFX1NKpHs/MZf1lPDdwWUaQLtV5MtrE8A3E/dAfx/6TY7dN
hFVdbi9iBSLOIYJmkP3WgDNHz84DPm/cA/7gtNG+bVzAEALs4ypbUi1IkVT7zB8r
yrhvVuhs4pCz0u0efq2C5+gV+cl+r9Gz09BFD8GNQXwmOGx2i4722/UnEXJMR2XO
9so6HZfAYPqQRus7WoSoK+r/GFNvnZc241DLmcahqedYQ52y1jAcpbASnLpm4Tn0
Wd61vcUB4ArgeBlh2BEL9TxtX8EAABrkj0yS0P6NMQpwoc2v0IXrFhzU3tdEW7M+
qeabwEAuBAxnVdnV8MpILnqwU4Gq/xmRcQ3mq1HlAOk+P4x6wM7X+MjgcxRkNBXC
C8JyoW2HXHEWrXEXX/hn1M5pGL7yH5wGJDw4uvKX51to9w2Rc1M5VyVDK0H1qRwI
WS1GIMzjcxrFpFZXwLriOw9fM3OMulepveLgfYghLiA0Q4UuyqgoX3ZBlu80XlQh
qsnn6dToNHJZm1JCn9mscJ9sYNkkWo8dP8l64VcnT6ywLCNK7x1l3VQRAkGR4oHC
hf1nm1fEV7PeH4KyXn21KeGySzJMaiukQwS1pBmiCZGW1bCFX6GwnQnFWEGeFSql
nhGi1hnkT2h9lg8hNqCXr8CQ17bnfA01n0XjMmDwiYlE9Fb2GzW06UCu9UnHpL9M
2ypKf2l2akCViRpQaP0CO6adRMWSwfdYiKcFTDD2YPrWeLn/JOGR3HmZ2gX4eIee
ZUgB+XWasp0kCznrbjP7DMQQgS8t0wkvXiBrjMQ2ks4ZwGE2DbSwLGq4SBhPRdzb
7mpxliHPnb85O+wIVH5gB6FqazaZz5kH16BKNHRq52o0uDrqNjvDY0uTxC6BRe2g
oWmnrnkyA+nrSDxuDEMppovtytjPGG4gkRAQJeQJEInV/CippaVL8m3kkOpQJlO+
kXCj1DSpChihEdCCdTdSc4BFhYLx18gHjW+XeoyjDyjSGqAdITm13nAPx2rXi8yt
Ac92d4FNsRNMuK59kp+UC1+Ru/cBkcHHDktx3waiS5Nu1/3q9A4npYaEM+cWZ9kH
HppUkQfltXjSsEvT6eXiZN21z2TcZyHsbMzcv6mq1EEe8oQUvNogyOkm/oFPo4Sn
S/GOe/hv/IMIZSxtuRi/WJtB0ORxTtlIl7N2SCtfEmZYGpRLRLaTchsdnNb3HVod
3BfxFqsKD2qAzHDWtHMuPLdi7AHMTAIC/++1d76xC+eml5pDpC7175uuKuk3Y9+n
/lzMqeu4jvretCngWgCoE6XF/NKU07WFkJq3FDpl9/G/TuvACAT3KAd7b7SUQ5to
ssYOzcWgTRs8NXjOYdwyIjOCTcq+GAvTYVxrch31yC/NA9VnyhmO/4YXT2NAIRWu
AJOj4RXxMYs8nyz0J3VC+l/9gz26Rkd1pRV+KFwMiP68DiakgEQoD/xBZxqzFjz/
4t6E+TwNaMhcD8c+VouI9nS8wwI1Qn38Lbu5vwHIXEsWuAuCBvw5BpCHoDy4ukag
ckgPYKzF5HdAvu1dFWroYQeypM2TCm+EUZVks1hOtekcjf/S96U8hsJp4aelhIUt
TK8iG30DXDgUgq4z8GUtv6DjgUXDlC2ZOFkuQyd3RdToQ1rAJKOUriCoj4j8V7nj
zlFdvVx175gQgezP7F0AhiYgkHp2MDkleKjd8cuqEs0rvXtpsMf++2ZQBphI256m
+eZ5Gp1tZuUkX0/odB4hGMkr1I70g7CrJzqzxkWHcaZySdw7381CbAbKq8gUt7jD
w4AiwkfLaTkV8TA98o/YvrwMsjLgPXxpViX+WEFwTbalDPz2N02CA0K25/+TY0ir
zobcDwdPnkJpEyz3V/S+nk8EcXTmi+MMWXj2SxWMfxfOdH9BmRnUnVxRBp43x73/
nYJ7A2vZb6/sB4Xz/397Tz0KN5N0/apXz5IyqaonyXADGac+kbUmdNotT3o5A6Bu
GyiSJqoJaHlljuJcB0EVI0tXIqJMnls+i5+iQlWwXctPbYnvlYfPE0AQbG34LmFn
eWksJ5MX7YN5/JB1OaTebDLcRWsmGUH0NA9gZG6r4OkViZIRy/wcDWl8J0MGcE49
S7pl9vFy+7YaV5MNvk6lZ4vkUjsbWmO7799Cv5AKPqYuZWZRPLJ+HI+1hcGUgL3x
UhZdBj1YjQIYAkJTrPXKNTSdaZ/ChlcKF8gMXY74JMy9tV6I+2ujLfp1JYDROHPY
4eCM7Ti/ldTpUzo7gudDmbDupy0ldAeXxkpOAFRD7zU8XNX8V4rkimGrlv8PjUNA
3v7XRsneYW6Rak1ohoJdtIGQUHtx5hBNbdm42BW5R0IpUuP6WBjW4rxFHs+/Fjwq
xpdJAtXEYoqPZTnfg4Mw84tjy8QQ1aq6v8Ftnkk11olrC/CmZGF6Iuc1gC+DLtbB
iEPRDl4vlJv0sJQJ7G+yLtwaosj89TrzbNYPt4jMFDbaelY39rOwq87XSj1XEy9a
ZCRUi7psI9Vq95CPN6yKX4Pz5eqBeHlAz9FP624FtSsZYszHB4S+NMPPEtZ4rN3l
lhGq76ayBx8AZ2B0TGP/DIZ1k7ZWFw9ZQLW+Wf1kX2GV7Twovctk1Q+LjiscG8xE
b+jzg9/XAm71Rnsi1/bRnDgA6mnRTSJDBpCk0v3tE+A9+lXeCcoq+STZCoRjMrH7
5Ey8/D24jX2QlSr7sS54Yd9ZpX8HVL/N9LImwKOGJdAkpq+mjK6OpOkDoqH8JnxJ
NEODtLk/Kgz6FLU3Lc1cNt+mX7AtAYGyysEm+ju2mbgsFhy22tOtCRlaGpRbUZu1
h61dWHO5kFEv7cIXPyZf9g15V2Sii2Kh6IxghkWIs8zz5CSsf+raJyj0//D207MD
izlt9gDcINtncStzGiyP5WUdut3Zpi8JLwM2+CR/u9JnD2eZkqjuViKlQ0pf0CDR
ck48uQuSP8E3SPGZFVonnnKOPTx++1J8C+p+Rb7BVLCHl9FwFZAuhQBv7LFMbPui
WOFgXhwsjKBDDc0nvPG486UVb5aHA00AiDqsfQJ+e3rmWjt7DMTfsK3d15EQxDB4
lkVS/vmfH/ay00xv+yvDurOr/xG70RA+xjaxviZYNohMjrl45mytPetahgmarRHZ
8RLE5zoAHpA7onpHO3I49pLl2Z4qWMzIQKOqDVSRsCJzQ+/aIJt0bEPtdowWM2rF
tikng1bHPUWtLtRAMReYjU3ejjyBT9fhR5RDiKfY1LU8Xek9aGk8z46gjd23T4Sw
LRWMb0s8F1amZyfsssdeopF87dz/zVGmazcVxX94zHl6H5sgVNHZ1e7/JZieZJjz
jcI8jQJNQNOMsKVGy61lMtp29526EX3GPfffj4ehcEQPb28o4ncTWMc1eD7JuE/F
DFyxMc+AcLH+MHq7OmjPQqsoaEfnfQ9nYbeLpNpBYg1PuU6d/YagmuA31yIwmis0
FiIS8Eu8k8yaZstxkPP5pwDxwmf7BpVn1F/0bsBZt250CCudPdCoz8lD0YJWoRwG
2xFiZwqTm6e3invi1r/KFy+jXKNxFBSV6UUdI685onZOWtgpzzHfcEeMrL9yIMdh
LQF6+TwC0kJxULX8gveqaxb700Sgfkksht8LuDxfQKnXjyzRELsWbvBeQCeDLzXv
V5ulPN4eh5RxTHNpgTRmRM3hJTynxdpvMBQN8xJ2petONYwq3gWInnIYSMPra9GR
19imE8DgGeVf31sO3u7c0a7YrIgAndrnwBYIK6cIUO+p/gAiSwzw8whTs4ZZvX8f
9Hu/sR6d3CZiKg/9UleUNf49Jh3tnr+C4NN8KaaoVEe/n77aNyj13e8zOSsPMyTW
z2BCqGqU65gjZBBzHaa9Q0m716ROVYR8Sc3qEWu/IacMotBC5gkU9oZ7W7q+59/8
OhMn9c9oT6Jm+oWSbelfqIiC1PSvBg7PnCrjUXikDs0UDPHjoC0nAjI4UGjYuhzX
yjGLyFSHuni/Yw19yvZ9/kftCzlgAHlaznmWlWL178RNugyTmkYeKTvnxcaeEb2O
wPDjLHlxQJXcRH95E/Z7mbP2ZQIpsN7+NmWa+3Ndpt9zPN5sJ7agGTz7/e38D8mw
lDUMliEyT7A7axyeG7nZ1y0bQIb23c/RkSmBmM2+o4Q+zYODJ1Nnn42ZcU6L8dh3
mzI3/zSNHwL7Kg2jAseqFPatBzYWzv0zQSzgmaf7+kltBZhPbavNOySkZZ/7MrL1
zZErDgQCGz9XHbOM7GV3j/E0/dwnifg3c9aCCWOUacK7fGspUAs9xMGdm6dN63Dy
V65m/wlTuhvpbrF7imI9w2YUAiH+4nw25HJa0DXySHD4rA7hnTNq1fc03VF8Z3f1
5FfJHYo5mzhfUyZ7PIKYRTm0QZh+tDYdfZ5ZCX8G5AMffYWgDkqU53qVvjA3kPvs
afjh8+NeXUfEiyGK8LSpcwcF2XmwZHHFozmIdlGfqSRolXSpZz70aOR+bQCyT3MJ
PPxt6Vl35bDPCc3IYN3JJCQAqWKS/Q30Foahn+L+jRS2Ph5t6+1SMOW1cPaFQn9t
17DVe7e1qTNGo1hCsyXb2HBfPUaA2pm2c9Gi5ewVYSn6QsNlTey25s7qsBT3wNlj
43XTecMnvMCTbZsyAL5dFZhNG3neHTFZ30thooiQ0gqjam533nNQfsScGJDouZyo
HkG2G8RvFAY4TdLCwPjNwgJJapzTZJNPCDwGTzSSEJQU8YhXWiiGSyrnhbduPeCZ
9saH/G5qh+76rXqVsF4EOOcyOOxzjnVKNf4wD/AK8+uyyW+gF5cluFkaobD3WWfx
ccUMVpxgCUhEigr9S60AZ0/UFexrblMX3LIDYsMSEYGw8ZmLoygO6lcPtalBctba
PiAlZ7q0nbO3ASF+aevnDEbdrIeu6DuY6f4OTmXSmhE+TyT7FqC7fiC2KDSuZNiT
DjltxAjaUOrZ0tDdHA8Ud+imic2R1vJY3ziii1aAdTd8hVitjfQEbMPSPjafi/BS
xNHwP22fndwbR7isdClX5PgiuIexdqxy+ya+XExuP/xXK/4EjDZuD50PBgsPZWI4
JV8HBUvQcaUkHZhFkC2wNx2jAZ2Ib8A0NLzqQRaXlms6a1/QSb+g7atSBDg3gkix
SW3gP46X10Jt0QanUwv84HaGb0h7HFdPTQqC+M8hEegN0QcAjrSHXaFi0mf5H5S8
gPPRrSP9zaIOO/K4PG6D6azuhE5p7hIQSKbIbcX7IvoHjvrMnoYfXbMEmJ8PS337
OSc9PIJvQ21oAsjXMecU5ArlcBPZ81zjFtWKlbwgOyUxFGepRQpOY0jOlOT1VHB9
r9IpOYswcaRzBq2898vCL/Xbp9GLV4ZEBkyvIiDpASYq8EEjmXuMfclu1eMHGOee
M3kteOiYpNnLb6rWRCFRyUL+pD+MqfTs34qjph+70hLws7lofv81tLUyVC6UDVpk
iClsLaINLpqTxn2Hki4vFBe3ks9yquwEgNSm9uTlyuf7gqPfG4WfrVA0UrHz2X4L
pV3CfzpW7aIpyAqtNShAC/iwAVAowdbBt6CdNykrKi3c7MxhbomZ0QPiWYzgzfwO
ekhpTB3q4zhjcXIhj7PqVElm91MMnw+u51eCP4KdkZmBbBH0tszxUQAFwtB7x+8z
M85PYBT9Mwoeythv3Qy9pwDg6WJ+yAPVqIYFRgnjJnWqSDiXjSJI9MlWEKR9MreU
5OGP9morIxzZPQv2MTqYc9ksxyECSop4DuEYaN5Mba3bqtKFWkepHVWwwVYHnqwm
4T/Y14HMQatMvq3pgE2QplKlkgPBQrW7RjM/5gh1uLLkNI1e7CYN0x4JiWqmeeYJ
JTxwfgV17UptjPuTBY1w7iaFJgWY6iyyBZLatf7OoZjX1VyPR9Mh/8wZwfXYQird
dhIH50gAEMlmw7rWdMS/c9aQsv1VacFjVaYu2DjVcyMR1DPR3MPvEEd6TcHIVZ3C
qxRhxd9EPtXxgd1VAv00dcNiiplmvLddx4UAWpogzdd8eNzQ4vpntK7GVfEJvXfU
aOtBd97hWltohJvOngJbBiIkz0nqGxtZOvw4YVm6NKF3kfo9NFEhGXZq/MpSEYOQ
t2ncPM86ICMU1LX0R9qVOTfKRNY+NyBiScqeuizd8fuk8Pm/mIOW8VUIV4LtOHeh
bHKHamTq7+G55bo7sJ3AhQu1+RSX/2q29Bvq3hqsCXnSsnUgQQDz83K5yUE8C0mX
jxg1m/Dk41x6ah/1W2HnCjERUiYMoxFHwF1t7PZ0XWZ5KgvHiJYHK3Hm5BEmnl6w
pDUQ1zH1b+LqDgk6Q9Tjm/c1bf91dPpmSbIbWl5yLhn+h2HAEBJWu2Fzd4u+XUbu
PuIQfiUuxGUtlg9jVVRb3zC+haRyc0vl8vDP8Bn9HDbbT6xmcFDVa9VRnLgp4deg
ZlHo7+PrPHoSojf7IXY843rAa1nsfkaM6wsotb3CRMXF/S7N+rfoSCFyLHxG41Cz
CmueyBd2ydP/+beJEehuZS3oZ+QZq/yLvGxjW67SHFbo+UvDDF5TKRPakn05lG3Z
7LJe9B8BY7Vot7Zq9RMzJUG8C8nXuYfer0ZF/NlCBWyQ8XKTiIc0Z0rrKDgOJXuW
H/coTlUPwlG4BAZ8ENwKdufpsLqGtMBVXeM6zE+ZVxokD9ADsVyHUMzhHW3tu3ww
+U6S0CmLH6b3VNo9JiXgZDm4xzN45dFnZ1sP+VeENb7hE8NsFhqgI708d4i6aNqX
9j9a6OMDj+j6vhDjjtXcOCMYKCTuAxlQe9sq9JBr0/ubsh4LXw3k34nYnqrqUbdu
72m2kvjIjWGICwpEMRgPL2m/3jV7gocWS2zXEcU8dl3FucH4oE20hRcbxIalUo34
Q1FJBu3uuS6+ax3KKSKPnGkp3ffna8Dn9gagjnEzi/yWRwBE7kPMS9LS7zGygYuw
ln/Bjy5OfgnQsZsHLRfdNpK9o4kxGeqwXIdaAvL8UiTYy4Rq3G4l0S9SnC4C4UtV
pUNp9Pweel/0lpuChunUkMXUne7CJatcEDgk4T1J6HJBw9GUWBMEMjAd20tYiWzc
rPb0ATWqUko6hxfjkfOyS6aJofGsAJhwxs7MU0lxFZJFiqVlCeNcKNJimObY0x/M
4a9z8a8pw4fra4nKMOt6nXOMxhF8OuhP7H+lTFmSlyqbmwEvysO3rK/6RrOfyG9y
STxH20kvcnPXXApTHXT1DAphtr/mN8j2WsZHqMACebbpo02fmzWuc+lrc2ukJgsV
BBa9oo/9hgB9lNHr6tFxcno2r713FaC+3LWPTi5TrWzTKKZ1Xp+CMP4xSCOAvfOi
4cR0tkkf7lS2ppoRfrP05eFU5Ovfh3CkORYmzupvWvdG3NdBrTQe+501ZLXHAng+
Xa67SWM3ZvsEViz5M6ArCkG3Ad53449QHV1A3cNw1CQQPhrH7TtDnCOOP+p7w29d
rD2pwK5dyg5IJKlvVD5qfPLiGlFN+7ka1NhKseNGuZ2AnVhZLuj0cvUGWwcMZ2je
NMggstamfSoWLf4gNc8cZQ687nUkMUfZXy0wl7FrUdHofMCxwksnrHwqJrHSQlK/
j5f67Cffpf0lMOlRhPPi08TBSb4ULxetJIp8s25c3N83Y6jIO/KjoqPz3Y0rnRJu
LUalFe26vk/cDHQbBBItB8uBgnHEiZXyThs6swzn90MI8wik+Zzre6Qoo9Xqw/oH
nmlJ1M6X3L1DrWFlhoP4AUulOhf6iQ5+1OhGjAH2GSzFXX+KTTPcIjncekO42fLz
vFmjtv00jaQd5PKFHggP4+HCh6uSPxnCB1SAccIvjUGERLYQGgvQfltYDhOqm90e
r/Mc0RzZ/kuYeeYdRj1vuVkfmit517ofZ0d4e5G9+rTRoerjjAtxku3Sb8M/dppD
PB8/jqSO+/kx/Gp4l73GIvdZ2EcJlMu961Qe5LWo9yErxhzbxyTcWtX5NnctHUa7
ai6Ekz6sdNp0vQ1zzUS4cCSoLv3ZeixcMlIhlFvFCZrkVbwY2pp0dtCGPsxWVoXr
EAGeSS9YlRZoQQVOsbVe9vw4CGjWAKPbYgJ72ioZcW9kWmJtSS0Lx51acAOeYObg
q6xCnKX11LtZA9h3FDrc1X9dSqfqnru/rKFhg6ic/meA95gnd1aGnnDsK4Tw4WK5
Xj7PtUa944B7cdKh1k82PpZ0upnUWhYaiEAaF1cdltY2kQPgYe4BDzIm+Co7RwZz
OKmd4n+O8tBul/AJ0vccJNuiUW9NIU2WZhCGIZomp67Hfr2yHP8k9eSOtX5AYwvM
V4mWOvWz10AtJrxwoRKBs0Q37NM3A9hGJZIJKGrCYimhGuecSqCRp0gD0C5mKThI
rS6jQLfTU37vk0BS1CGSt4KdLuKp9H7nJww83aC0rSexSynPl5thpT1IlPsn6Ldv
QwN6Q/VdwMI9fiUM/EbVmgrbfcd0NM8tIzryZ6k0i2rFCWcve2Ybedrfj3g8OPdb
Uo1f95rQCNrW2h52RrDxKAmrxq3DnSZloLN6CRVf0cUNO8hfEqBl7fkW3nwb4kDD
sHTz2EaIWH92I88h0Y4MDAGKz3vqu5YxiKeyfvc8RrTbxk7wNIO3SkUi2dYV5ujj
9nj2UWWoYgpQjbXAf9ugoe40WM7/Shai2lmlTdrnfA7ObswD64SZZYbYu2ftjoW2
/qADTm9Aq5Q84lKTc7KSNtSWKih9YAaHCNG6BMfg0yjvaM6/x91oa8z+hqTgB5pV
O5UAVA+cfkM5HHiC8qdslWIt+m/2DJ59Pldn2DL59lXyJYGS+K0uw+HDWokShsOF
WRDW9dHxbb7FcK8ic9Ks3QvS+qFIR4nvHE2zLAZQWU4YvADfQvqPMrUhY8OZjh9U
zMD/e++7ZuAz/8ptdIMc8EqhTIfiKQy+u+VOtyoaOKv3Wy1o7fIQEyCVolNPbQcA
qCLX0IltDnL6iKizPyb6iyGisZS3UtIU+DcUt452byRvGWrcKpCx4T5Zv3q0836o
7tl+wrHE2yBJ6L8fuTmqHa9y4RvO5xnvlDeEkHb+TkRvy1qXBBa9EuY2ZwkxJUV7
UtaS94z9XcgQIaY1O3BjwBS1sTqtKyXvT/JgoKUicZ6eTGCBkYyRIy8tZLBCOjz7
ihvzw3DAsxOvuabKG+NU99Sok87LBxk/IXKVHCG+mCGq34Gw5QV5URbUgKVAbxm4
bV3WE+DREKYVoIx8vwTsJrFLU+zYMGE9OLT36nM2TC0CgBHd+DbpvBiY0qkXQgHS
n6sGN0ZeN3JhFldEbp3rMmF/aaesWbTXckqPIvuwzs4RRf3vtt0XGUZ88cLmoixT
L2NJUl+X5whXpwNhL9vFi+blF9hdYU8XmsLow+GfPvKS+V0EyXHVipOGqM2fJoan
tys5BXbPfeuy2H59XFiosqhhu0adBr0FsHXxC+Uhl+wmFZBNGUw/Zj4M0xgF53Fn
3rFAA+05+FJydFMQeOt9RceWnPJBzxwK9gDjBgxln4NPbLF/0aMI+Ow+npTdVYVx
ssFFLItLDFeaFbNcQPTDK17RhaSqt+lzG6+mkUSz4cPflWwclpb/ah+5l+0BZX0e
8f54gDCOrcruS+tKp2dMW1mhC4QJiEoT9eWvGJzzy5l8ihAl1bWUyhlVegRrwbii
d42BhzipbAOpyGMr+XtrKRBk7eu6uIGGdNanti/YST1nQaQ4TOKbqp3QcCjw5S3j
KRQRHaS0urjDIZ/EI05BcSpTMBg3KJisrpNi1FzAyImYeLfYyMsQaEPWedmnVUgT
rGIwWGQLEEbvA/RdK25+3+3XpBgO2CFL8Z4XZZB1JE2eNKsOMH+BnDasy2JiYWoE
grQfPfcstkvzbfxyXIvG2khpViANFGDa9nb9suq2wUj4YVx5r5JivgsfsfhyrtIN
ZuDqzXdYjO5KG6H0Fb2HvEwxKtZxkxYcUhi22gJVm5lTCaQJ5GLgqcxuymFuWMLz
AyvKU8ueeWyAi4khCZeGlfDjYcpYbymroY26o7v16N5LDo8yA/exjT5NpKWdljT7
C3owlun4PFIn2B8n6D8Za5l1nux4hT5+rYl8Y+wipLRqoyFNaPIG3k759MfyMJc6
bK67DgFbmA9nJoVzYvFSiTa/u8H8laOy+++cMMdrZ6xAThJylHtjiSyVryKhzVQ7
zUqaZ2KlZz2m8DY4BqUA0vj2vOMsSCCaKlNbVywxRuve1vYBlDpN4+KIM61xQ6z6
A8WIhrEeVKqRuc2R750KHpl9ec06nfELlQyD8+Czq+we8v3qG3OD0SIr9Z16Ux8R
1O0VT82+YkpkeRUyFGW9ASPkJ4vAXXAmiFUW9hS4enRhkb6lwpL2ZGcYZBmyhIbR
dB/zuW2yc1ILaTNK7+lLArnpYDL3176rvVk/fMkYjr3w4GU7K2IZF11yWKts6lGd
dgQqquhk6JLgx2RJ+Y2+mpAMcJ5SLPaMNpDSe8a+XMMlUdANPhssUkp8lHSko0c+
l7RfyRXSH6TMQSXLJwuCkHSdJy8Cdu4I6Xc8jlMzdVrErnqa9BkHPsAb6ibLlVVI
Jeiq4tk0Ddo6jKC51q953IWgz8xn7KILaVUnkePms/Tra7eEXzFnPgfIH5OL24fq
qEcctEmNgBz/wa7ujaqgfvEFO+LjAnNQGzD/4QJIFWz+vYyJuJXHgHw1i5IeiiBZ
0EKZXF9zrs0f55fxl8Qj32KD0EJsajLSaThyzo1I73JiWOGiCrrwNw7NuezstuCE
xAwtGQ902W1KE8jeAfivjXEs92F2bTVSGu86oxkzBzDzvbuMwvx7bWwkw2IgTdqQ
0rPL4LXW5s23O3PTPqQmPlNCOwqltJT8D4ZkJPsnkSc7wZvbaGaYRzE+fN8RyedZ
uAOE86HPS86Vp1vMkQ45B0tj730/a79yN0A14utZsU90YfNxPSprEZWK1PACq7fm
oxHU2I4t+LElxEEA8E45OZKm51dREUTkBgcl72uzw9CfpG1SeYHX9/y8x/4hB0hA
fiGNw7aH9isyFK5EvtoHZ06QK/ymswRXufvD3NnzGRPBTV+CW3CfiQNoM6jEAwbB
c5TY2Bw2mo/fwC0/O5xeb2kZBUpTrmVrFM9v7BvHqBp4nfPhuQBUzNb07OVPFcYL
6vHyN6A34sQeKnddgBtVQQ1EqSlILku8OSwR3csE37RxSRHQK/S9nsmPqpjA3voN
dn6zEGBqXu2D/x/LLB/VYlKIVhbAWKT+4YhkJvSM+4kwKhz2g7SpMvb18bE1nWe5
0WYssMoh3Tj9vh9F4RTgzkz4SNeIJTeIXVpn8aKht7y0pH8bGzTJheZ9QJE5uiYi
RV6EQ4p5n3Msp+bq8ehbQwF6yR9oyJ/UiYGfD76/NK/zUQ7DTnJeO4W/pG9RBo3y
mORnSv8WDDoeif+haVydTneLjkZlzBn9ejCvT++VNqUDqKcFvB9shy8O4apGxLOP
EFpDTblIuYFiW5x8os22dF0VBHlkKSswicpzKnEbs6wd3tN7IES3B4gBHTvN3lIK
4fmZX8L7HzpVTU3s7r9sQ6gmfKw195+j6RmdjNaxhXLbYjSJXCzTp+qC+P1z1aV1
s4sfwBKtadl8IC+7PNdSo+K4WtInjED6n1S9UcAFz/wRwUlNL8CfU4sWgDUK875F
VEw0ANoaXjL/rEWGTepAt6qFDtvJufOr3kdWf/0uz7OGhON3eLE070+W1LhGdgsX
nKL9VX+zj7qBuPBw4Mxz6gcyRI/IEHI2mz5I6kdPak6RE+tcp6muPj5i0tmSSHl9
wSsGWg82/msFg13MYucll+iK+bz5d+OkVdjYfWikQFpPbmRP2KhSp0D+qCDewkrx
Q9b9flFM10GeZc0JmbU7fRIM6ZK1e4Uv/FU4kz+RbbFnK1T39X5ItKJt+orIt/Af
1D1mKCdAEb8N5yHrgTdm0qDRCXB1RgK8Ry31u59IsVo1zcw1TIXOjJsUnz0XF2yx
AqtQwdvuQqR8g12i4YRRruB+84SRXup3iycTmj9aHGNDvngJY4xrFXFLIVTfZFtu
SZ6rHYy3xrJXqVZjB5zxf0EiekJ1HOxDqAVP5f1ZTaF7762jy7qxpCouEXAR7PdM
YeD/5GW1FCOSHFRVeZhJsqNeSkLuBBSY72lH+4Goz5DvqmX68avx0BvCQn2KY00b
ISnqxYyjVEyT9zvH7qjXb2a4LjSAF2IT5gfGnheOIQdpA01KEeoTbkgS9iZ65ooj
L4vww5E2axWpQxjARYP7pZSpimqwtL2eFXwCIckx4T9imi5hSz2vvvvEtJiFXWs/
lL8S3QlAUMbqEYahH9oezT2n20vY1NI4qtHAL8bTWF8Xvtr1x7VepbN8k1K/Glp5
25Bj2Scx+G8sPuKSOPDOAXRLZyc5nJlIx2SM/59/WHMMtCat2upIXlV0VZqP9BMw
d+EtgQkzGE1FRt45+ruWa8dPH7TB/DjYUTtw+vOPLxaECC6EBzp0JA1sjiGpy9we
mR9H4DjtM5Er4BvT+QzehzQy/+7HoIT6Zc70+gX8CCOG8uNLN/4lIOkPPA5RzZXP
jJD8IEtWMPzIi9SHTrCPlNpgslNhpei9IQTsX1gwNaHkMWKrkUTEqF0iOoVLLoAh
4BSiayDVemy+hox3KoYFi2HjzNPoepW8oeMFTCL8bpaekr5Vg5c/21XsHckKcrz0
vApZjg4PBSCqNEseAk85AQ48MdjrbwanMM/8ACBJizG+cPbuhElg/sEy0i8xxH4w
jAntnFRvwCGAW2OMD4rqdYK7V19oE/npSuJM4ZeG4+94vFaIPiy/oW4mXc3jiAmm
N7nEZQ0lVaAfee3vrivtLCkWvEiB69j27cYjlPOOQ2hQH8HBoDMh4snKUt8hrWtr
ukTkJYbEFelyAQKZMKs+nqx+maC9HDgIeQFkyAbXSiXHRfKXdBNI+AOb15ds7HPO
gVtLvbm9KSltZtc8TvFfrztSBWwojkkd1OjCBcSeSNsJ6hHIWbacquYHaXZyP4VU
gWDNrO1ICsI/5DenJvz2+CyKjBPeLVVOXTmxrOI/bfhaZqrTjm7KJO/H2FwsrN/F
mtNkevb1A2d2xnqP1Ho/T2UFAEi598y2vVsTRXmhIDIJlu4k9GifcSGkdP7DlaGj
kzF2WfncH9AsDeSF54TREDRD1p+DlWLTA0ZMThoA3wuDLaxmme0kKgsZ97w9nVoh
w7hLrJkG32ljmaCIup93ZKZelyCvkm2hta7GuDyQIxgyd3k5DBWGzHEzCnhZHE2i
0HmdTxhdA4DU0AzR0ACCUsd9LQVVyhSwLEf+5HUd0NrF5xG3C+WQEZyPx8g501dj
n81vd9BaQ5OGWDMF56gJLOsp+cLIIFQxLUfm/pcyWVn1dmgShNXN/KZPeRfpXZAN
tTIvNVkpLvmOklqx2J2gPuYkQJikkIwTRXl/gRkVNLSsB0RH7NzPHuojOnT5KKE7
z1NXuHYxoT8fwgrqJ5uQMct1qJWs3Kp1hZFKALfzUKCvgRfajw+U7ITWF0FSXBsw
8NM3YlWuAFXzHR/IaDRv1NopYyydu3exSppkaaonXgbgkRu5aTN80ZFPWBJIg+EX
tYNMAuYxKfS8Nu79ygeGrGb2lPHEM57g2mYEyXDzvGqO8ktFhtIK9Am9qSE13uaU
ZVlX9w7AA3ZOCCVggYDxnTTg5V5tIt5kfncAV/Fr9Ei0JpryNCAT+CfUbri4/ek+
ynCye5JHNDImcCt474mLWqrKd/OY9NAD7BfMxs2n7l1kgUIffSFkjeCFtt6y7DvO
56EjPaL07MH6JqrjxjJMwPAIg6/LGcfuK7fi4/qSg5APdQpoXiSlpWv33F1TnKn5
ckjcy/X8gVWVu1F7mKe49IYqSQC7KEJt9wp9iGSQKSzppjjVkFlJv3ueDD7YOBdh
dNcc+eGSoThSF4ue+9PqGb3F1F1uxa6pZhRAhw5uHxWtercJEWAsRLQYX+zGdBpa
cA36ihGhgM1FXjzt2Hu6azF4Sr0ohEVoN0FVwFzfSDVpPmek+/lFMYbIZNE2PhEd
ibpLMHFHyABfLiV+vHZVUc95bHmsflFCPPMY4NYhA9FLdVqX7LIVjq/uCtYjpGBM
Wr/pfe+wCb3rY+U/BRCxN3o2NkhYPrREsYNMe9W6hi4QKLqYeh0g6yAwYaI8Di9f
6Qt3v1fJFEI80UvGu6nr9GjmFotX9KAWdK3pZ7KP/ZBvKeKAobObWJKpq/k/+tZU
0VpSKbG7Aeejnzcor0U5SJLe+ujvuAwIJccvvLfIKmQPM3yf6HhhQNi7zb1fxr+p
gd3gscX7CLV5CSwaAX1Oz1Bdvj9OxoGEMGntRYgQbxNOgmO8JKZolcGANy9CvSEn
aUKiXgHNCsWry8cERKpK3yfEJKO+FjddcrN4xhzMITpz8Ya2EzMFRNYRxY64vNxL
F+zTY57u6yUcouZW/BU76PTZvKSJZ645W/yTSSV0kQ5/n//k7h6TeuI+TQ1F4MzC
KhCHSqngM+xgVMWe0UjvSQTtW9F4sJV+NzMV+W0zaTgR+b9lBFZINurRmbBa9Ouh
ubUaTZ0zZamdTAkYhG1oiWLCSVvK9A8sAwGtLL2MHZl3G5iBSgvykg1SVK5VKdlJ
Oos4efAQr00I4bSXLZvgoXCtNiN7nGYse1FG9aGaZ1HYNg+JtcbPcpU6SJCwW+G5
Ai76MnurI9Ezq9KpzfUr4A4UwXu/1jjHPhM7i3cpnG7w3HNlyVCbeGc8aUOCLq0P
FrWb6dNMQ82FgULEMczcOipg0O6M8C+kMw2XpaqdHXg/EyH9rabg3WNXblHLQJhy
GX3UnT7zPld8kEre0ukbpsLwlClMwzyU3m4IGyQGDp2jK1iK04PUgHqXqDbrvoui
gFofMxOe7Kpi8MquEKlbi1vjw0uHQIiKQgHg4HKqVjfgsHkUWFUc855a8OesoA5B
ZMUkTP/rID2fqIBnRpjS9oY9LW2Ylud6GHSN3Vvh2CysveLBlqBJFBAqEcxhd75I
wF79FusxoPWEQmCAsWJ86CXv1/JA+ISqfI+OrEY8fZh9IKdMACM9UBcNlkKI3fqp
etT+jyPTzAWcMlhhxTVMMxN5YEfU7KKDOWYXR3bVQuymTT7BcQaqyufbhM9ebI6l
v1iiFQO/MT2WbUCoPuKmcvdBJZFccBXxhqzm6Q/B/8Ve5tk0J5dkdBZd+AajhmUA
o31O/WqPzjqUKxjIK5WOE4zXr/niLpZL6oKDdCnJkq7oB+sWq/IPv0mgxocMlFMa
m1cBtXJi87sefLiUd6AWc+tQdMzSOBzF9pGmT12pNDowXWS7msVJ7JbC8uxETK9h
G1u97iHBu5cmWm2HxgFzt4gpkUSk6e+fOay6cYzOLZSUjXL3jPdXdHw+BfCwD9k6
nxxpFbnPOWgglf7LzFMu00TaLPMhGbcdnjHTPS0jObmDXtj1Un/Ge3WPaX86MEEf
wXWx0lJq4igTGQATuXOUHneEswkAkjdEuYWUaDeedD8TRKJSJxXN66F+GyEaJa/r
KQBk0vKAMM7YWvjm38uCmIwumaY3eBCdQvYe4sYw+77V/tawt6Bo/h+8Vo7hbitn
zzlewZbcjEmv4Lb5SI74QW8rvSIFUgj6bYlvaEDM/CDDqzh1ND+fDJQbmr0AbIm2
4yM2T4qokJXaqWvIaXdTI8a7Ctrm8pNNVTwhg+cdjjpHJIHDSsYQUi7gPl+pAjGA
ljW60hpF05goq/MfJ4GySyreT9AxL5L1VdkYMJXwzBSEnZTP53VMP1ZPhBSEvKKP
yCG0h4ArVgy3iNcZAjcOdqvXNHVQvUlEI7qnFr2ec0UTzGtT8thLVvg+R03mBoPD
PicUJ6uQpWhe7QxFNizqrzggT9qV8cSNpYC8T00ob48iWdO+RlSuy80MOEE7gTMp
oiv/PFfe19RNsq+j41cmz1p2MmuKYf8Tgtom1l88FGOMLGZQKcsc6CcrB8UqCRed
xCdo7hupnCAyL7DwR8Eo/L3fbdiE6tO9XkZqbwuJ0xcY42XC0td8r9UJIQ2wkqhW
zK3Yl2wf77RCtN/TheQaoLsJF2LSWP8wE5BQkWInQYhomHS7MswCbGmagZn20gPh
QFxC146oVNQ+YZv0sPVBN72obYXDnnWwFJKku8WC9rlhik+D9+8y/F6KJtrKs41z
T+qOx79ko0pX1SML6DQXs8bfPzoSJkbc3IBo7zU9Ko9XJ0aGVeQtx0ZsvykFRHN5
2WGK9e2wmqaJ7XzZrTPZ0G/Y5/uU3QrJLRUuQMSABwrJDX8xRSjJJ+Cgzh4FxEB8
9TrzTRBlC5XZOj50YJvmKPBi1mT8fFhyIjGkB2TY+omHIS3uamb7McAxPR6aadR+
/cWWl9Loyc/rWn+am6gzDd7HcvGZEsPC3xENnkU/P2Rg2bTyRMNukKdHVVT9MaMb
z/ioqp0CBmjRlhr9YiNklaBAYp+cOBeY++8d2/prvuS7nnhZI8a3xJR9aTNfMXWV
ljJb/2X1kTGZHEGmnG/zkjNi9JNC5hNuPSxCzv3EUDjI9iQKp0VEuvj6hN1UZaXA
iU7gannckPunRddF+a9UBkIxhTrclTuGaoeZMwDmXxXBl0122pSFYL/iaDEodyOc
zKwknC4txgmT1M6AXN80KBmumJcng8Vq7/GtVjeRlOMFDA8mLDWdkbhLt7ijQVsG
aD3hFB9MuuyfM8Su9o1XpDN4AyZzOTbzNLcmARzm3F5p0Rdk1B5TWQ6GG7/WBto0
isLsZnoLvTY0oMUzM+HAOSRel5TUAIB4duwr7gRQIUbaaK8Nfi0KEQxnecItXjMX
hwsY1kQ7YVd1xFzmW/tsUFFntxhHIvh+hO+AmIS2tEBERrIFzl6KJ1V4SFVy+KPU
fiUBiMX9ErYbunnRvDy8ylYyUbrKLhGQSpKUblRERDxlQknEnXr8Uf2mG7jYNCrP
oqHyj4a5XZRAE5l0eqFnxEQObzMb2WZW3lPQe0d9X5mDfA80yhzRr9K3pd1OMhQc
WEuJ1ByWX98xCiBEjsFEgZj+6oW1jhyHLWRnpbxcN+tf9qt3rtgW94ALdiHyCTfL
grIQMXEYsQZPdpecsK/wKlcanR2OXAaPxWIML8TBuw2YlCANSLbImr4KGhta1K04
ssl/idz62SEHQc5OHFTHTeE8eT/kWDtgpoX0oKmH2BhSbAec4cv2XMoHoIYRzz3q
Gzqx/gS85GpBe9EOuRSy3umjO0kqHroerAEWr7Rhx3A9+ZNZ+n/Qlh9IAHnOyBkp
nQPwGMLKNRpPttnAblzdv36J1B8zt80tuDrVFiz8lDE44g7oDlzzTgWmtLeR+f3I
vUWrI0JdKzIuOn3nmDLDgH2Pz5pJnk4Z+TJA19eC6FhWBl4SzFIQz/zahWh5CViV
ia8WqwNI2tyAoEQqaCtijIW9uaucXVzuwLW39DgBm4m4TG5wKhvGEV+MvYWb63Qp
rG8czoqNNN58mtTkOb/TmKcnAAT03CH/+pBqOMF8VlqRcoULTW49oU9A4Vqg/nai
TXieWHIIBywc1tSMoF/MRnCB0RGVrkMDTSKUaFdsW+VoFsmUmLdwZ1kXhPfzKvOo
FTMhWfkRC3nCPcfDsDesQvYAtR/J+vUArGQjxkI1ezO/5eB7NwRzKW8Wcf7D4KLc
HpqHocfs7NwQsRib+Nek3moy8YY+xiH+BSr8vmXZDZ6a6t3NP6eScvomPYn1zQ5s
bhyVC+Xn1+lXkV/Sapbg25ApfJyJAxf+/uKoSBorNGkq9/BOZRzTGO9BeUB15GoY
nUrCpDdxBQ6A6Y7h/6IvY25Gva74b90xBUKX0HpGCdn+K6bombu4QceOnZ0h5EUA
L5TDJEF+sIha/H6ihf+yaLbNAsGu9/GK9FujUDqxrMUChSXhdNwy/eucl8a3dgiY
oPh3WxWTou+UBKtTqSSL6dVR8uzWvxBm9U3MC/p597LUjiJKK5MA6oSf8Ogrtenx
MCcb3sMgt9OwgdY6Sje/Bupf9/lOLoSWHudUxcCU26yO7Otw+N5hhs0DJN3znug8
TlEcbznxKd83kmFLHK0ZpwIfe4IKIoXc+aI8uMPTKJX2rV8ayoU/JuNQYd9Z99As
fEoIOfCA9uUdhRERQJYAlwYjSlgdHm/zEpdXHDqhoLs1UCPNxYnlHwVMNAXJbKCs
cNiZJTeLy7rdfcpgk57OTEzT/RDbtZoPndbchydYAiTXgh5mj/hCFcFvq4tbwEG2
LmNjgzzwXOZFXfMqwUODMSlwpQ7BDHFhzgQC7H6ixeFjF/4fiUoaYQDgUKBPRBqY
011ZiLJavF+KaH6ekdQxa3lGKeR8lmW7X9fLL0L9a4BCgYHWKFPcOPOXVVmvMAJI
irBgl5TPN5K8r3qn3tGDEbONNTVQTe7UUcxHXtxtI5JH8Sxy5bvHKdnEv+YCQK9l
YMhOnNxU+AZiBevyV89UYwkL5313eWjQ4vWZq4JbI8Kzk02RhoLAp4mXZhcGnd/2
vlmRDX0QSgP5u8dXBHxUblV4zx68QCshfGk48PgLYpIhW4fXP0XKy2y3sczsr2dO
VO+TH2lD2eRBxIq98UK8B3SxbSHqOa52MzaMGEMSjdNtf40RDX+ywBnpAtiZDbrq
OFw3crqeFjw4C7S8lMie3fyDbN29YFYikmzeDmJQnElJlObIO1xQkWQHrMII9DSq
v2Qu29amNiFIctCU+cRxyetGkI1fGBQv8tSVCsYQ185rNvez61SKY3Go9cIkxxTy
v96Lk40AH/59UVs2jDABfHV53tdxEklx9FzVLgUYgL+xU2f8Cg+njMvUxpzAa+xg
HQ536UwC6BG0bwCSEfZlW37pa/hwtE2vF+WYzXek2mDdafqNjEcpyw2tz2iNYi0s
w3K3nK6UWDVXnj8/zH+ta9q4iGzZlJ0pY2VhtqNs5S7WThSpFzkU6DzveCNMI8st
3/mgbzuvlwZihm5dgXKaAn3pfWMo8sQpOyOBPaKWAYY/1/tGocbDjzh0wUZCyciA
gaj4Hl0tA+J3rUdHYnMKohSPoTisKHVzIJMdkgP3GQ9endjqTVQ1rOY1c1N4PbLr
YDxoWLZOG8ffUeZIXmpvlb/DR64zS+ullTJ5gBH5lRPbp18yMD5b8SxEQys3DRI+
ha95VDyQrDkApDbXG783sErvmQPIfEHqIk0Jbl9XgT0m9ubEc7pG8+zaW25u7fzA
dz5wPYXH+/mlc72qHWb4vq3g7kwLqYbRjitQlKVkefliCMrPAx7drDx+oE0okPt6
BtouxHMO0PsN+OMbZ4hxy6/rFa7mc30ii8qd1sjtGKnAEJ+WLXW9jQyCCATg6ad6
SOm7dK1WTGcvZwjrCrT45i4sctv7wJwarSvB52vEcGDZqsthCW6atIiWLKXNIdXA
MIg/s7dz8hcklrFyp+6JmCkjsK78GutVUY7D/Id3O1zNBOtYqSx5YG2thluikgCo
7fcdX1oQW7UeClBnL5XJ2DuqRlK4wxl5nGgvW4qnGSP02yxVAz9/Pwy5KCRe1gSx
NbVQvfC4+zM2Z+yIwSEvdHly6zsvW3rptL+GsS5FTGo+bq1+BE/nr9DxwhWDdLqU
SoX4BCJc3H8TOkwu/tMcBPf7mqo88sn91bCbPwRfzRSoXmq8cZopH2ILCVyPm110
P/mWN4F+kYUwJEynzHFtS9krCqqW3UCN/rT+rz3vCxHL1JngnSHcS/7yAfqrFtGX
F+050Qhuq0CUUXmpyHO4Z4eCe52JDSL12BrxdKT35lHALzBey5tTgC79Kq0YgpYt
1pCw36+FAoJNznlQbUNBol0JJ+a/JrNm7pcPb4UsjmGg4BPfNoqjt2SthRcCbi7K
HK4qOfyYe+rbjZYEStSZhFw85FR6VxYB2HYuzbT4gg8C9myLWj+CxubdGvJlx/Bo
WFsmtxkcKBDjxjK7MbbrHp4BIN3Wqa7V2IblywZhNxk5T/6+Cr/Pw4yiTmwhOxeA
eLTDtIxzbV+4bUwdMVbmXs3p2brj1dlQ8NwnCsWx8grpYlu7uBiuzI9nmf21mIE2
T9/B9sia7yfGABZkokzOhn653cY5BuX8l2Lmbr/g87xbKqMGkvW1WHVciHc8lwI/
l5lsmhh3FVCOS3jBTe4GC9giIR9MOUjdk+5sOYpntxBao5bOdfxnyvQMm0a1CfSq
LKTdTg452GyVJ+hbvxY4VDEbCmIdH64oCiatjhGd/XB++J2KdYUbgJ1jzrqxbWi3
8nPJC/emPAqXjbxaqavU/Mbp6WwJPsmjSplsjHRhRj+hdQCnlY8BMw/0CYLbH8EC
T9HULJNZ7Kb9313rjHsH+DlfXccITz0rBucKuHjnjq12IVbmQNuNmFA7281mKEZY
pi4VXPhbL/n9eDArWt6TV2M18pTobC546nGReptZlEqcpYfOj/ln0v56H603NM8E
j/EMlSq9dAxnwl0h4oz7/6Kl4O7uCGDds5I6+FM5mLF1lmOFHv+aoLgfQopYS4y0
jNaUEH4Rgp2a+yWCq39oySmeepuGROcWfIYgTiADDBmNF4hw/4TaVT70AJgbl01q
XbY5W6OitrG37QI1BrZDGtkBzQTyAq6K7H2uX2IoTlA64q2pmipI374kaduDMLs2
yW1NZD1iTM2qe6LV4/aZGrBuumnV3FPDDcMlVP5LPJHJUbYFjajg1bU/NAniqiYf
GPE5NsjFlJ7y0VkW2Im5woCyxvjOUtFkwBMuJEA03zVuqfowr8IkwrHGzA3CG40f
MSJFg7mxLMarREcuoNWGdUnYvQJSkhN/RKRxlpeUeDkgNEmP3l51G918K8whKFtk
e0SJBZSMDAdy3XQQeJQQanvJhxC8tPNT+xuT1b3jP8AUfm/e0/WYkmmdWhNDyXUS
lB9l/g9CHQmklhMcQ780MQOOqtsuZg2HIyIDysZVB7DThZjRRRDvrVoecpJ+Ns7b
UXDCi9rL+R4FDwOXD2JA4K1mFyY36qeXahzR4H5RrNCzIz2d0/eBoJitZbTHD0o3
kgYPHB/xoUGL7Z2gGL/9JUyqWwlC+QM+R4qeJ0xroSIMNRjhcyOONsexSBglyAGF
mJYuu6q7sB5XGtniXzuFNeUfYEx7Nj5OL5GeevWsfjNupyXUtaRLxy3V/NjoLnaV
FKTcwzfmh1seWfLiTeT4nNGT/IOlVYFWcvxKRSFTb8bGu988e/gkAPwlyZ5AFd8O
jJJclpdjmcutgEuia8HHCV+KQFhhzf+u/X6P3sgy4x4avUS8BqCkBCY7L09XqueC
zJVVQMHjtnAhtl/3T+9SmGdl8qDvlaeLJxXr9BVTd8zINmD74RWFKhlKjfthduU5
NBS8VA4HZcCOntRFQ/DbABxf1WaJBadQKFUk1zdjc3mnb8oIb8Kc4/3QcbS1kzaX
qSGyfPK4v6CGOYuVBGDhfMWsoRemCdS/WLX7VUhZ3YuzXFskx06jDueCk+CfZL5s
Z3oP3m51BAaly9o7LxcEUjl3Dztaz/OA427gvbJ8ttlqIzuzOa1lISOn4ogC4yzV
zm4QnmrQJIRMtqdpq88w3SsZq6+2UAEbrDHLVIDoM1X9MsEdYXZ2kk/6CkHG+8+5
QxTesPQdyHcgbaMd+e6g8vsgvHgcVdmD0OALjuqkos6XgI4+KtVwfxqAyHkFTLzS
2/2pF9/NH4MsjqYyPDCPKcyC9ULcV13xOsxLJ6ieNOkyWI8UcHdXlNt7UgKnTqMl
OiHKHfC64QCknoom5qEYkcoqf5vsIBLiDeaC3FPPXU/VSxBt10bGUpUeYouzivF0
OnIKddX4BExCeI8918d2CbAlggvCk1+R1lic0xVviBOfT8qe9xjEMRO27R5eLR3a
rZ3QmVunVb2wypqAqJ0j4u91XYKNOYzCfSGPmTaggBYrdsOJAXK3EHGlnsILHaxN
0J7LRe+rbrehWvrGbFNrHdi/rA7erajGjE+ua4YPxfFTT8jnLrj6gecoSwYx2e8l
NX0qH9vCYpgvk+bLcOLlrOv5IL3YMAETEKaetknPs8sM6FQW974Zi5KawfJMkuEV
S2PnAj4BQEwQuuMFxkNnZ2FCGKH2PrysUYe5oXBF8mLs/qdVkOfxu03GIpCwxv5V
VM50yj63MUjoC+lHPFhIJeA4ZArcVJncgVDdoiK9oTXShpeIP2fmJN4xQHm+DGZL
NTFPv4lMAJElB0xxIqZI+9h8k32V6HXQ3M96iYGosAusfrB78ySyEcIieiOPI69W
4LduhYuXPx0ZKUv8ypnSQpRZz7oPBFbX5sFg+3Dc0aAp387W2KknFdxIBbFbWxz1
pPhrnANn4JwdE3vNFDnoh730m3oauhyCDFo7SjUlN8Xw0e1HOUBnT3/ue2Q7K8Dm
Zhjqrf/CwuXE7WGzJh406AkHcTpeyzpfVFWAbmOhtos5bQ1v8kZ+E93XxSYbRv4f
t6/EPhqkGrCUyYNkVSJfAUMIcPnENjqM1aV9vhp22mV5YTAhHkzl+B92UldTHOl9
HChcY3vHcLP+oowL+g62Ul5u0oqKUSr5Y+Tl94ZxoAbRL9xy5mqrwXywNj5cKSSl
BWtmURBIL7zbWcXIEP2Hn7cxDf+bp6r6pvlWhxOiC/MOLuxi+02iRtLNqkt25i+C
XXPS/sCDZ0M3EnDi/bioztVmea0aBSkxqSOwjTl54zw/hGf2RzFqaqINLf/EM8kM
o7GqiB0J/6Y+vw9PNWox+CwHEVXyyDht0yZeLRPCY6t081Urtuz47cv8hkjMyd3R
KTG4OCSxXUERxl5exnzn6aGZa1pGfBWQ5nPcUqwllX/RBa9wIOUS2KehL5gUp5EG
5AjVwWFxAkuvdSluG65Qxg9AJ4LjCKxngSGT3GeoT9WkAVSqczi2Ijf802uh3g4Q
nI5ehZmYShVtxxK7G1npfKBTJwXxtQuswnzQKZ9G0GUTVpSmhX+OVC7iW9zjTd5V
Bd/9vtNJunnVKQqndqUvVBoneHncykp1VMgwKWg7Q+TMkZxtBpOAgH2PJyXuokme
cpSn2yo3oSjSWq8hf3ljV2yzK6rq3IwX07vDTxS4WBBiO0EQcg98BZ7+0Tw8Wtc4
UyBzjiGLOfwzl30OdwdSXttQE9fl4HuImp6zV85ZsSl/JSnU8T887XmSI3tG2Ja+
dj7QxCnT3nqRVpdofsDNJVS1wsbJg0kLCpXRC5rlpQ+SYGCxJr31p4txKfMrprGm
4RKecTz/as75ROFtdNHufSGi54e4MnzITDWryX1SMNSQ0fepfl9yc2DNWUHbxBUi
nvYu+uRo+ygV3q4DnbJDd/83RI4ebHhzrhFmsM+DEORo0mZq3F3ClJGWlzgzjuxX
lP3yeP581frdP0ltUkyqGjndBRjvhvYSqXwtj9zTwteeKZ+bE6Enx/UbJ9JxI2IJ
ny4k6uHoaF7BRZta26y22wGmxqm3Q46Qjy2QOUhgPKvkPzUvwCtF0jiKm1xD5IRm
OHT3w71SW29CvC/1pIxfTOG8xWmoy1ozwH1Bg8Hjbu2y2vvE1XSj3jjKefds7KYq
5RyQuU6JGR5byPzmHs+jEX44tBYUO7dVcS3BkvMlh0lAZ2s5Bz2+gYXcMukm8QLf
RlJHQbsYG+BTLTry4mAV7nt68SBUFgFI3TCW3KixNBqw4zE/XjEquSlgzFmEr2EG
FJ2797GIzNiMnjSy93fQe2Io0b3p4L8CRxU1E19XZm7rCCKH7rgk9m4S2iLb+XJ/
akGUSHZHwk3XO7sJgwjKRU8fRpj3x8F8hDV/RD0bhlqslLGtKu1ysziilCjQrMZr
Gxtqt5fYpBRlYik54WXaN3Qw40ceaCp4uIUqQ5blgBjWVTUnBAQI5TFcRIKdBLD5
UryUhuG9RKjDOY4l6wh4uBY8ZEWWQFf0g3ci27YQAYAZYnM004xE7kE1y3RuuIVn
ql+IIeP2AqkIAss/aCXzAs7zkXlkatiQWEpvZWBVotjjeXAj/kj9EC0FywLynY3Y
gk+w9pG7HCIrXBMcT2yQ/JiUKD+19Vs1M9zfGmpFJdEOdDybVrSScFlPtez2Z3tR
YpC6Q1BIYkLwsobnZjH22D8l9vJTdKd96QR/FPwUp3oIFQUhwDC0QLxy9NMpe5IO
Yz/e6wkn0NqrVWPCGTSNPx6r2a9oSE65fXh3bbnCz+7iaeRGJ1k6w5FGIlli0EAN
9TlpyHZE2XcONqNniVjxYYgrap/3VnIV8BlUxM9fGO+ku1sMi+VdLooFQN42JzBg
0tl0wrJBcZjfM5EZef+koreQ9SPI3/sW+G5JvvgzB23BO+t1jzpTS8DflLv3ExpC
vKxqwlHI7DpjSntpPRMDoIrcjwwg32VqHilt8TrDGtnyPYxVgjBLCgGu/FecTbTs
fUiPWPtWkFlA4YWvf0aNspR+KjF1ZAsgOmnSYA9PXhesjDKL/A8XD4PmSnB07PlI
Dqd7LdVm6bGuTvr6ngsYNkNh3RtjzypMOvgUulghYd49Kd4S+yq7aO22GHzpzGyJ
ZWlez6HyNNEKJuYf3e6mZPvEFKH1XZdqaCFRMOjYGsCRNxSFpToRlrcrxmbBx1gF
+TWA7xFvaCbfgqLVEc8VrJAb+C1iHm/LLFxcrxRSctuZoCw1mP/8wwL+q0Z4C4/p
5j/lvdOhQYoY1mnKL2Z7ZilsnAVgry+YTB+VweXmlxRzaIwdnu597w5iPgv/jveA
G2uuq29+sXg2zcVOHAGNn2zmBFPqCQU5xSDv7hh//zhGjqgy9KGW0FIO/MShxYb8
03cbP2r1gOqB4IRd3LuHNlGDpoI0Hq8CJ4p6HcgUYvDTWTodGyBgfaET8Xt/0c67
9D88AeGtaE5jvSJ4UcYXbZHYDmkIY4P7K/Z29ED8owq099noQ+e9078VmV3v3ThV
GiLbSmE7HtsVO5E3VHWQjQn2KM+mezkrkJXI2euffMb/C2bLmASkl5CCz4q5n1ZW
vCAJL9jYpDsdpG2MboGlA814cQMXLgb7u7k8LakI/3PYiOuB/Z0TtP6IRcZA5Pwy
7DBgpP5wS22+2/NW0mmHtLLKFnJjMjUJB6/ZIN4dimspSJeGWsTkYl/BoPUjJvp5
q55pBsw9qp8dM5pEPxRfx1+0Lg243hLlYznuXMUeTMtMA6VpSjgfgIj0AdSU2vR5
RUDcFwPoie6U3GN2u+7e4sw4KnetmIzcgyblsyNmpsAD2xxq0YU7f4Py4mvHAe/5
aJwf2XewDnyn0gIvG74abYoadc3Jam1B8NB+4r4oJ9cAIdA01gVAKMZGF4UGVV5e
1M9L12VHqBpQC6fmY2KmgvzMMo+jdDmGqDu16MjtHYV15SKlisrA1kf2uRwJnVew
ia90nbWkmufoqj0we9uacDpPLPy2T83cL+d128XPQeqywP0nDcBQ13KvJXKa93T4
03KzksecJCao7DPKWA0q1kFi8vN7zpRbYst7oKhIV2D1LT6MBOIw27pNThnOmcY1
r3FCY2v9VB/k2LDfk5GzJz2QSBikwrj9oLcORiFhq14pkgh5AxcJb1oJyDRCi+px
bgdoxiPum3hGpmj9Voz6UoqX30DxhcZJl23eLEhFKm60n0Thak4rwU+8zFEhBFX5
3cPqo3hJAGUUtXtVccPaQ8Nu8y/Cxvz7dyteJ15YndfxOBsoiohs681CTyIcKc4U
VxQ4YUWo3UaBXe6Gqe+d0B9T3fM/+lWMxzswGIo70pj76uD8yQVQ3H1bj1+ST76D
462hHTMHoHTjiJSXlTQZIU6wDhe7FM/JyOxTw5MF/hY3NisvspSw+9+lCf+2BuYj
f6K7d5XHUgIpdsdnj9wR7tflWR5Ww/v2OXN3gpnjrO49SI3ULWu4UZx3TnngQgzE
r9zDd/jVa6eQixhl1FC2Pb8FEill2gB+/0eJqgblX2aSW+IASRIRa48FlVfNAci7
J8QBpDODpIXnRPJn68MRoIVRebSg5wVqodeZGPMpGDzLqMFkYnhPGK7GmvVzMMZN
jTdeKHS7oE+euLzuE1GcKYNI5FJN6Lgk9jBfmXfla/lXv/NJXnQqy0znp3H1xY0Q
1mP0ec1FJe+9/E15VJyEUlgqRbH8V4v3UuJu6x2+9cLWEjFEwVT7RdqfQhVwcUsc
qeieWu7e5EgVOrhwGh7f0s4wGwvDeFQsutav77jul2V+sjssdoE+JUC6s/PBMEv5
dcEYD+asVs7XaO1kFkCCwYzlzAbxwbutB28Q1KqFQOuOmjyGwrAEhBasuYi1pfK4
IqXlfBsNC9WKFFAUJokirz5yhEjleZFCUNruTKkpWHoxj1OsOqZFsmXHUknltPr2
QidgbnmzYtYwK8ypdNN/IkNvL2t11s7z9VKkDjXsimopcEUCig/t9nsbBURFZ0eE
iGPXKc2/+rv05M1uAhiYDCn6c+i+Uks7+no/VS6bLLTu7zTo/aNRMNF2A1llEBzg
K83Gl9lOz61QSb1eXX1Q1EqtxGB7j1CvdRxCXL+JWfYADrJnJ1OEaITgs0+waYxI
gkfEAmlv5n2A4tNPELSdSHvmWfW4x7te/+IoL9Q1qUJPa+zgyLRuhkTP777ciDxv
AlRLyI9psz+bkwknOAkxlRtySxuxsDcYLOruqrdiu4r5FFVQIWs8+xfpVsGlh6c3
EtDwZrbJ3nLvLWBJMUNjzSxtnSmGiB/ifGQU34zjxWNaUURJKE+TrOerhrdyk5xd
VxSPnwHhr30A0zwj8sbGuUtuxiHuBKtTVdhIkEpZ6YiytiZLI9E5E9M1R5jwTVxh
CXu6H1QY9gFQh/ywVvxSbDl0gbZlfbz2soSY5gVdLwBBnZ3UqQw7ix31l+Oqwr/N
NB9tJkehNC47zUUeUAUx51wT8OMA5bWzGuyzCayiIHj6+TUOl2IdIvp7PVgkEMB6
I74BNYBTIYQ7I3TKxl1ay7ScZK3ZO/4zMWQEQ3jeQSaj/miazVNYAHDqfHSICq1W
C2ObV/O5HBCj2HOozdVAC93N/AgUSetkduLapul4x82Ts4OFiqGP7lffqgv8qGZ8
MD3D144mkhJKrOAvUsr1qzp/E7e5EA75hIIXw4G5v0/FZALInMZuUi5cMGP+r8/2
ABPWaAfolKEWOxkT2Teb1MHxI+mhk2ySqLmkEXL2rwMbYQa6Y4GjtAdmh1ZHxQZ0
fEzdqtCovEFfgy5SZQ2bcQibpgdOA8+By+5gAfncdpiT9+jNHw4Tf/hkbg/J0azk
awxPg50oKFES4ezGzfp4Ih4go/NiLSVQaotVQutSEis2+szaJqusNN8+nleLBiH0
uZBfg4qGffz3AHEEg7KDdlQyeNqXm5ayAEGhNxsvlPenfYyNfR+puMtXyjjmzp4y
Jmv9eXipJcMFzieFSygG2OQGqjLxYkf2CCPkMo1TLUHMONPZSJ3CwoesUN8URLgW
jHdnenJ7TcKBDCvx5g1sfQMtp9JcNerOBrsfeu1ikqUKc0+i4j2WSby6Bu2xrC5x
jCK76rI95Y3MpB6kRAXPVj8J/LzJGogtJqJqqEoKFxXmkayKpLJQtuIsHTf9Xpwr
fYanCx23Bt8mD9RS/ah15Vv60lXtCbP5eEL2ySV4t7GyUbY4/ezycqa8E8PjYTd/
wb/EpeTN+LZoV3+mrRrAjs/6gM0x3mt/z5eRDbMKfiyftnlnDT27HlbeA19tdRGd
/SaY/2Bi+M7+1oat9uTz/O7Xl//tlUCdKZl8KAOp3Mxy+LxQi/oIVCkfsY1Lm5e6
tqH/PvLszmypte/8JAgmKu7h7uO/WSGIeFlyseJVwOWLsPJwBUsz08cxGenU7W0p
U28KtXSdy3mgygAqa1QoajNU+jk3FzbAGzXAtBPt2HRiaLn+dyKojrzXzJ2UM36Z
1FBDDeIWPcbyaAqpPeQXmbz/1E1pC72MVsXCmdO1TVKI5PXVsUbALaAZAULMy/ao
lBYkRXrEwpOrYniOd1Hx5N7Hj8LOt6TStQ7hwUWAs3DVTiRnrPIm0p5Os/6huF4K
dwMfEfHaalOXSPHTZpeb0uKCoqZZCkpe0gxobIErizwn+W2UbK9kI0ChRKiJhyMD
Ft6kx7/W0mS0kGtWzE+3WCYSMqnxv2LQZrSyYbfLUMYIcbBJ/KMMjvTDT1H9byQa
QH6ts4yAY0xPh8OLe+cXH/4+pZ4mnlWlfbwzlUNUCidu6DntVmjJRMKF7aG4OCUO
v1aJzDtAQxqVELusdb0aI/SIKhkZmpQXfkfTQNH5/2ZqSIEcM7wdiA/rEWoN4rGh
Pfo5bsraguiHK1o/OUt4POPd7SQKJScxcZsd8tOzbGCDRsH8OkO69Kzme+UyVq1M
TwcUFwuJ5W0EP+dmAUO3hBkzWz5+doAeUsMbvnxgZZ1+5d5n2PjcyacWm/DK60iK
e3elUUaC748ol2FsTL7s7+lR3kHGbk7vj4EG4TOlo4PGZmUUV8RE8wVPryFOxCCy
KeCLf82NfC/Koyhc2260mpi9YWG+qKSvgTMtox3NZc9O3Cauf8ogVHdQ4o9uJER9
N5jFxHu+d9QyltM72ihRhLfdn6fYxBsrzlSWWQ9uCJg0qsdWA23yGSgCg2gLyeAR
MI4cmhBgesSSBiLtq8nS3o4f7mE21skcDMIi43v1p5ABku/pnr1hfBp5RoW9MTyZ
prYslRHPfwHZ1kunrm2XHQWVGzFgdJI1cxsxcu5mOtSzlz+G+0jJiCpSRczAXz/0
pWsJwNdvB1X/IR6xTaC4OEOzuVIn221UoPwsUdhDPmFsLz+HK+2IJrprzs8GXWKR
k3LlVEoYv2dEAPWGgiEUf9Md9KNBhoWNMFt45jQPToGFhZRJXUdZz4RcmcS7BQHG
Qq/YilahYL3mhoTsI0HpX2BNVNP3vmh867bR9/T1uTNhKVfMb5dnGWMONWbPEXot
qfrfiKbxFU2+BN8bI3kh5pB0m8sIfWADPSNubR4jrrWYNpR31fkLutj+H195L8nr
pPWwgQaJdb/Ts32n4OtSuVHHR9bF2jyk8j9LVbVKuDeln+OUsMPLb9+FGNBP6KB8
5+VZsaiGVAFySVP98gWNatnUN359OUrFRDAw/WfQXLhG9sAOT0g4rVmsIcuTFI63
Tpax8VZXS9oX20z45wLuaRNqjoRQblfpHNdFgzjnewWr/KIbJSwWW0m8lz9gJU1z
kXiK1P0okCUoiNjLhYJWmlMwIxfXl8Gv8DSoyjZqBb5egClto4f/1wt++pCUwRvH
hbQPrZCQaXaUsd+u5WKtH6nysR33LJwkSBnUawnPHlgEUPGwQcYF3K//4aZSGjZ2
LvP/AD9Wmt5fdPzpoeYY0lr83wKG2CEXpoT+16ddBBha7BH23Sdk/nUGp2xofSGs
lLZoxTPkOQhlH2wAjvATLfYYYXAybqjJ6zK8cWjcXYig2zBL61dsBiii/lO7UEjl
GjUwj5du2LvF0qLYJ/pJ5MNCtebrBP9C0rizY9zVfH8sOR3RG7nyLjYg60vwfyoC
JEDprXTZAwn3i1tBerORmfawQz7UlbajphOgr2kDRe2OJpcUFqIxcAhZ8JHTo25u
It5fAnagUcn2jWJlTIIOtl3sMu9RhVD1CEsuX8xRCVnzC4ZE6dVJHgL7aHITaZx3
TYCr2w1o+AzFz40bOUQ2OwoS7M2xHLQYH641VbO+X/pL4NyRikX6wOrSzqV/On7v
weh8Y2YyGHzFoiEJFN8qVCvP9Rm2tocOiXNHrl/i9V40PhlwVubQyVmiq7zpRsIX
II2ArMqtyP1BGnQT8r8yO9GpNF+zX1xOW4K1zvY76nhMBt34fko7eTAz5F401zJv
BnSTG3fNsusBxNZpa0O25q7SZy7FFLUeqsLnJad4XfSsLzTW0+JnBBVk5U2bF3C5
hhZ4L8JSkmvRqveCXi3uE7OMaPb5w/dJykApp0k8Uea7mwxsDuIntVx/kLkCbWpE
ApH2/t91r3Vz4Grwpuvwh7tixCnN2F1Asfuay3jLW6SKBvERJMvvR3cBMirOcLBM
dsls6Jc4iCccetYOoLGPOHwLpku+CiFoMBRufYqh9vFVgqi4mIxsxgq620hUhTy/
rVNv4Ck5gUSWWVA1i2oN656lQH2PvXU00GMvkv/6Ds5z+RGgZI7e7kxpFopFAOEt
RBsaMOfPoHrGN5UOVrawuM79xIWShsiGrnOggLFEyLttZAN15k1AOXi3AlYuhgtW
n1q//qT7FJd3WafpVlory4fFOC+Oj1M4lSQHNADRc1Ih8ZaMEdIsECGMWoVDuEVy
1h4UFwvBUMNbCVIjRD8S/jtTGM0NgWUbhKiM+By3/wYUt3H2+hOWG/119prjn+hc
z8C8m7IuZivW6YWKNOfmD5CJMrWMB3wgxslc7AqKYNGoCTJMga9vy2y/2SNe//o6
38RIgBj8E7Alrw/Ox0AQA/GfF6WSQT4NgmftWkNjgLAOYOwLpdxlbv/Mti5xhwOn
gcaMVdvfPN6wkoYGTPTnUbMOn1LEr31oReSBSIWma7Csym4A3ZlZLPP5rn047IiA
77+8PrGXKT/55gqO+CdpDREu4Vmi4VpuaCasZjujDSaGPbHBTqIE0Kl0ywuUkyB0
q2lqyWtAfJGO3I1v56dhxFKSkmMCQ49c8AmS0/5u7VlmE05rF74LNDz4N8/zeG13
/Ijj7C4Ge1x22VTpmglGyYpVPvlBqpAh3yESAh9rx+kOmW3I7fyI3iAu4KEZhg4o
9QK91gFJDWdXQyIX52fXDG8QKxkC5+AupPvyhcw/u1tibbGtICfxxtv7ObB+rxx7
+L1RxltFJl8An0c2DTb/WNeAhh6yYD07XylLBBuo9kxHgfYvJl5DOxnEfkgVT37z
9P75HXUdjJIzC4E8ZxkmN+MPnJ1BE6EDi9ZV+lZi0a95sXyx0jiR1TwYK20ZSngU
pYmlT96jHm0AGRTT9bRzPenxGzXM5EoC2M62RjxqXmvBwBtcgYf9IkNIxz13zKu6
ZWEFaTHh+6SDbAJ+jUb79TH6Hc69fwmIGebhWxxpYsiQnIMcM+1fyp45UJiH6N2n
vDUvt2mJ16gW/f9ZIVnUK6xlUC9IEuct40YCW/d3FsUrx5V27JUgiooIqoqMj6LM
BRPjEk6Y6itS1pTJ4cmhTANFvqz9eKOUGPbv/8nmw9DdkJvvyc+M3kG5ym3nxq7O
5x/YOYmIj6ByHox9ulGD2PEAYixidSM7Lz6Tvvs95bcRRo+Tpsii8wpuwznNOrm0
3xZZ5byv4xF3DkrzGVyRMULODVonyvAl7XJayL/LN3F5iYzKMijIQwdqtffVmdou
237Wd8r/szQrl6fQ7znqkvwRRqIlI4qihSTtUaFuX2zvI0R+2AjF5lnSc1cGwnJN
Jq5AK87yTEMvwinr0T0NDw3y4SoYK7HnSGLuauVPWMIghvDx7h1cR5wPHPcBVfTP
ipGT5gBWnd4BbcciggKPMT6qtFMBI4hHAJgJjsbG2dCxg6fUNho9Ar2os2d5ZKM6
P7ZuD25dr1j3zbs0HcmeP5amQyoJYGYJz3G+Utl+wV7g+/9ZZe0SG2PW0dFFxQb3
wd9AiMdQKptfQcrdyHH/NBQZv3l+DQVv0BHdAKpXRW2JSh0Nw4v+FMHgxyOPxXYV
UkHr8cP0ksktkdDG3VKUn63CBu4f8aFLOBASeEYEX73/aWkHNMyHR7Qeo04hfFb/
Q4QGJtsnlHR0Z0qYz86ZcMFRbSskn9cBOc6IKte+r4sf1QqOYPiB42HF7j1sXdl2
rYksxD6PDoGfva+0BUQuz0jJ9XyctGnbYhc3u2rkboOBqyeq/VDY7MJZVPb9Btyy
BuDArdvOIZA7z7EwQK8sQ6Ibp5bWSZUs+eZoZ2ex+rxjjMjGYLKYBDvBP+s9DnK9
Xczg9jzKzYjhRaEHEKHNr0TMU8mFdNXjee8SKOESLXH6wnOKhsC5ADiDz/sTibKl
4UXRg3RsjNEXnXF7pGmmB7QGjKAqs32eLQsA3pUxiODffyXH3oR+esRp+EpTenM+
AN0MVVaN0blagnGJIaAzeXNAOoPEOk+UyLV9H6RQsF5aO5aEGF3WH0r5MG+5gsGP
v7FNTpDZUO0K6graS+zf/phcqLGRghuTi9BpsChBAP3DsTfdYZCEind56YlFOQm5
K49Ch0g0pKUm0wHzU/Kdy8tqBKmMLLxrVjc3YMJeFtQBDOeGnHY4HeX8zQCBAQ2Z
AiPUe98SQY1QCgJBhfIX5bIse2F4KTSXmG3SUCJU9d/DMc1YU4lDxmR35TnMMzOk
yB7ilsmAp+HRwiXe2A4oVwV4MDAnSv23k1oUGpCX5EM5xNR6oika4UAEy8/eDO8c
I8V5x4jHWbFtj5iU2srabuFdrkCeXFXYoaly3h9NGsjbDq2D7/nGFe9JopXxSQ7+
T8Cifk5moD4EHfH+z4t87K3hY/jO3bHbtlHcZLG9FkU83tkfYb8x9YZbz6vM1YJo
Qe8J42lven8ZxKIcvK2cDZF/14Evrpm8wPHISs98SsDJSgWiPTBuCVHRpoeEAphp
nl6u9M8K7q5xTxFNqcidD2NWs/NW1+tGIJJ7+P0XzuwotWWQn3wowz6RCiOITOe3
WvCIOzj2nPdYJ0DYkBFROomnQ43YoJNzPBT9Piq3TIVml/WmSh7mZK0yVf6ILavd
1bF2ZJj9bUy/SdZ5OPr/UCJh7Flan+yoPhWCUHf1UGD+xaPn+AhdvBV/0eKP9sXk
Q9WzFsIFv41freSMguKp3GaocRUoydFI9Dj8Hej3y89madj6YmEQvcJQE1I1h/mP
UJ8Bb3IOzSEy1ViHb2jIrOROCI35oO0iQaorrbpPj6NEtgiM0h8W1CUE+s27TSdi
/HcAmdojJ+U+8bp+bZhxyezVmrlytpfqwNDgymk1zSK5LSFaTZEkFVrviZHvugoA
0VKmDmyAZqoQhQV7dXDPWGNyU+schBfQ3STUmaemP7qULrdrmAqmn+RxaYzouirC
DG3uwpguqDDHedu5DbIHAYuSQRhNxFODw/gqlofgJazqPYqGkvnUeaX+iGbAzHNn
pDrqBjT/xPUmXZGlgAcasVp/Txlo4rLLYNCXwfKv0ipG9EQr9r6F6SzBqOqhy0qi
GKIGLWGjHgjND4rKkG/pBD9ohs25csQCC2Mk2hLb9il9X/xVfLKpx2eMVZ5/oMP4
B49SMUhq9p8CTvO3lHtvQ02FtD22fKY/hT9EUUc97EKzJboWuqnJB3SqIUT8oMZm
Qx4mrdIzP1jkdgdKrYzH5j+SIAdep92iMImDx55Rg2jTxeNzbPTdmzZnqjIiky5Y
ipHdgpt/1bzNzDucoxc+q2Q1HgyfkJmAwo9B+znfId+uPWxDzHmXdNGpNGOCs1E2
N3C+ZBHMndh41KGDtQyTRCd/nAuXkmF7hxfO97zFha+UybXzD3n+WEkHBPM08JS6
d3dcsVIqAyD/JiwygWDqhpg7xTqVnpFRCjQtL52NW1FjdFkRJx24Y7NMRmxjhHW3
AG2MJWiDImoN2jpqJYbfh3ULBN9kJRYqUmRrQFaPx+U5u4RB+Rt2wMLaqp5CUMrw
eFbGql1ObutRgvvvV5xubmDHNRC5XPxK3VLG/0zyySwRkjp46FL9v2gUHB/MjEFp
kfgtK83gDUQX4GFi3LYHP74Q2QFH6dI4czbVSClRao3Va5SVCXEwwtUMpRUVWK7t
Jcsl+bX0p6q6J/tLQC8lBKBQyld+iRPd2bm+WABwa1raUjLiwD3ZRnsdAj+kT3gA
IjNs+T1pdXqoNNjS/1pI6QeT+vWA26nSh++EkLR6SCPi4KpCp0s9ObrP473qi4Sr
ePb9BdygXkoFQfFhGSzxpV8OCUqOKMBGF7uPTkKSsUw/I2RhNdhFVd9C3/YyG3M9
tmaIjUAyef9zMDipY248yuHY2vHy1VZTDPlQuHn4kreia7XwbP8Zdjao8xGv4JGz
aKkxnB8Yun9wjYrWJiZgMIO22LTMg369csg+UgKQW3hcrOEvhChuxcq+tYkLLvn4
cKvb3mOhu98nIPj4bce11wo54kxaL65inlQPZKvQB1dv55dGMs3nBDjrrw7t9ji8
/9enQ6U+UoXZT6C6JU6ag6DsDfs08ZRRSK9mMp2h/RazXAc4HeySdzEspu7XIzek
g/IDkLGOur+6ga52/8Dy3Zu4DMid+/VTuDpuYxVxxA2eLWS4in1J+3kt8rH7fq7l
WeRBB+z82BIxdS5SZOPl/g/5yYLt8oyMf1vT/aF/rTYnI9qXPJyi10geH1arFaKG
I6c9no7Ly9GgdDcC1c8Jjgkg0fWUfhIK23fm11vCskaY2ufooE47Z5isKbdqc4Gm
AuLpIddkXz/ZIMYjpjLo6EVn6Dv7Ndgcje92aNnU5TGkLV8CH6y6f+dG8M7QFYeM
/HxH9Hcwfs09XJwZQi8RXIWmqxH8+SfgSWQEGp7YS3HxWCb9lLE/YeITT1gPrCs2
67qDGW9020pI6gfdeoXlzfbARCqoXvnUsq3W0w7ffWJvBt5VaoWppo9uRsM3HcEn
nurpF0rbX8uvIrU+5UnqP7XzPTS4oaHCc+tLbtI5UPTPjp7S3axKcyf+K94omM4W
kAZ291Fh37prPb6wUh6SBl3rHco1OLO8yJQLEH+owz/M8k2mII5RNn/OKAu1QlpP
n3aLAmEfsvg1Ek/8Mz1AKdsCEIpdoAdQmoWY4uIVja2UdktVPSTm5oqEw+0fvjuk
qlDqGFI7lKCSxAPderWjlWqvWJGrxVqy1+Jh2Q8MdEYoT9iLhd1dVkaLkSkU9qA3
OX1YsIXKlL4GlPRQaHTOPD8b+gMFBUf9f5OyydoRNWugen3P745iQV3I4qwmzG0y
0tOwUcgwFiJgb5tFtkYhAJQCceIrcSikI7H4+BJhAc91DxuYo+gN4usTERjX7K4c
Ez0zg7A40uqAB2xjllDFKe/4euPB/iD9/c64koeZKnzgA20IMlaIKCI9mKITB+FS
UMekVeEJvYjvd2BUoqag6X9d4t1Whm1iBS1f7idxxRKi/nDh67CyG51BihV5Tg3D
MvK8rnyGFyLeiiNMW5aWj6fvO32cnSy8Y2gAykeDidlLv/GQyOBREtT2vdn3SV1u
86rEGeMLsJFYPFjRjgsoqA+rdUHz09VaO1KOPQtnIHwQptSfN9XjUeFld8J0Bll/
O27+CgfoiLGgqB5k8vI3zVPXcPq5/1IHQxOZW8gusuaqGhNpCG8RI4LzidLTECqp
ZLwv7X/GGvRYbBCYgPW5uxoXFV89rgPsxaNNQ4NhAwtSlS4AI6voZyS6nfwFgooX
uICK0nQcgnTtcmEgdexTpBg43bkHlRk/FXEZJO348jp/6XXPCf5VOSat9EJG9vUp
q71ofwynIbIlqsWa1us0g5xvaC4DZUDHD0pepfUu7hxHft904MZPy7twdHpkIBB7
qgN5rYS2G4JGIGScBrRUogT3ijxdAhOw+7OL74G18OndPep2AAizmfbDn7VuFFY1
kxKh3G6qaTLRMnQIEZSSUJjnSYvjr2d3mcbKVqFVJL7klTTlcLvgWI+s/PWElh9D
cFDDgEFLGFVIfCPKGjeF8wtWFu3xB5GQV3Q0x+eUDXN3BtzgHv9bmiXZie3NJquH
qRtfp0/vZ7TfP3snQSEsZ+q6pL1XAfJsflnh16g6a8mw6gO4MpsxfwQYMK9GvTPm
insdqiDLGgakfyKXLZsBIRK2hnjw4rozg366OO6ZaYzNp+9KruemDPpDO/Ekw8G4
DjcqQpZPrNTFImYu8DXoWS0bNuOZtqTE/tN9hSgv2JR6HDyKTAczfZ58mgl17cLL
/js6AQ0s++vPZ23hz6YTN4WJhh+kCaT2xHcpHh0gHh8HtWNXfMLahoS24alHF8MR
Nc7oWvhN3VEZT8t44VgxgCrGwCQdK0y9zp1VW4rPyYFE0UfJ+O8Wc1PBKvIMUwKu
L2HoJCT2ldkm4xcAU8jPbXfhcbVKFYclPoe/4XFkYYym0WcKdQx87eu1EIIBUlEV
RsDmg5Xoi6/KIeAdYmhsOCatYYZbupdzFiEwllOCc8lOTf5GCH+KZBh+6rkI2IMP
k62IXC9pAt6JR7e4zRE063SKjGixIgAh6mXVzpmLALhR8KnBHYoSW1+pDeGjLbu1
BkfrPNpDp9wqY+KMjlT6CrQyU+mR1ckbW+k2cA5+j+Y+0uGlT5BHoibNk2LMJ45i
kgwFltVMEMEy++Gbew/oKi1UsavKrvVMkHTzynGZy1AE80oqq2O6meYRO3wl2QCp
vouVU4kSVf5IjrRVK/PB8obNmzZcCG9JZx/O1lrAbrmPVIuVThNQQr1yQlx5DLhW
pO/TZ/vQsLyRLYhAcvRj2ijx5f+/xuFspIAIYQx9zBa/kOH5SLtCaYwoMr6M1AbG
DPC7RspYrjRfnLR7l7Jyq/48cu250zLMJBMYM/06dkqBry6LG1MnEh6BieHrafFe
cP2X58GBE0Tt43TIL6DvdTP/GdM9ROV5zN8hMOYl88OzcGAyu8zLts+A29nOMCZ0
1b9tQ1QfS8PHX6pkvyx9tu313vOteaB6CNKNDFhqNilewgf9fiRfSt1D4qtIG/nY
Adi/7AKiQ2KKN1jgjgKfsStlwdhAwhFffZhyMPL35JmhZV7mnMNr1ksgYQKj6LBX
jNfGYRfbnp0FV9pHlQJj/iglcEtv2YUXZq4EI/uECXwfUCntNFmtFZRXLWH2MOQZ
av0ytRCV4jUn56RmHn89Pp/AyYTZC9/O1EI/ExrP6AIe9FPAVUmz1q1kIM7qsrdw
K1jTq7kne5b13nOyYS/y7iy7B79BO3IKSPRmVsJnRHRmTh1Jg2mBsRNC11yYeiJE
DCHyT07qgIfXhqFYFOlMPCuidtOyYqEH/+CxhRHSopG9KV09LmNsvGpyJbhjxfU2
dX/WHZptEXeUChDwFY6Hi7+6/4KXOLDvz2lsMbjgKwvCjpPvPCqhxakLcfVXTFn1
1OOEGByv4JVzPHfphs96L7IGBfi88bcROSJSdzqXgvx9K5EFgG5N5ki8L1MWlLCz
pBKk+3oUNMHMjBHz9dPB3/mW0Pmk/OnZWDavPw4deTbLtF9Q7bHEtzShOu8iVZ0T
Y7UnKT69v9DIhzVb6BCpOvDN2E2f6eMbdC3olMTVTBRHDnoNT2UkIrg/wZgCWeAb
t4WxXpOIcIswYh14JMncBav9puMv10DRZH1scmEt1iC5AtCd/4iutL0ujjxnhwJv
8y8DQrGIExWmguArlKmIBG6QX52VW+MZM+dMDcmRZsp+Ks+nBwf+q2XaM5GWGpKZ
dFoDbKdUF5e5IMK4qOUwT50YUs9nyiJM644lanoPuByRo+8VOD0TyG5KQo6ZvAPv
q1WkBrNtPoTiFD5E/uJs4gHfXJDc5VB7n0d76xLEtGFPbtiErLA9sf+FYTTEynsz
wcDqmUnnabxtCNxUcClIvIFbXzp/E505k9caMCSO/STfKJZJjzndAfqbcUuuMdQB
b0e4v2J/YEDKapm2cHyAz/JEOJHSyeRcfRut4ld7XNHa4Av4QW349aV2L2uMkIWH
qtv5LUY0ufnWsrqH29Q5aZsK6bmHp/a1JY8GquvAnPHZPkBHX2SGjwzzR2Ud6FAI
mJrgzqmxsReDxzXOnL4CXOVvxptVLzhin4hPWjV17G6XmAjFTKtzEsmf5PiiQvcv
EEmf4fdMGixZ/EKZ2kAO719FW/VduADKtfCgVPJwYVfZokbi18FaVEQkoEMB92Oi
iCt8YfKJviQHTHaBq4Kn7sdnSaYQKm5wYs+bu4w2xuowXmsNq+SutpqedUxlESMV
6uer6hRLo9wFoshYSOAs+6cXQo/jy5XH2Wkh/fSfyneMxzrHbeyvePe2EBBWFfY0
HDUf0eW0swvI7UB6v9bKZ4k4GK3zUflGjTniqFWer/hAoil838dqiBGMKn98DIG5
74rvaRgiMbt3+dj5UhTLHWV/48S7cOpL052glq7PGsPBNBKtfsa++OGdclg9M0so
WsYTgPmp9oHkOVSLwfBbw77wb5mSY9g7z+CX/nXZQSHnV5zQF73EeoQMfgpmuijO
7YvVLI6ydECjs/X+Bz5VGkREbOexdckK7YFvekpMd0uZ3ZZl4MS0R8ICTiyC7cfD
bFoXrEY8kqAPDa3HswnVJYQcFNHLT9oHDV7qjyb3NSGMLE1LWgjACMyV6vy3E2y+
kAy2fm3BSI/Wo5K1y5uKaNMVtAOklJxeL9jwLwPb8aPIwirZuWsqrWLRDG9Zi77g
gf0YY6FMEOOtcoSnQ2kUD0K0ut3PIRN/GZEsqQyXg0EBmtwkDSb2SFfw6ahseL8u
3BDU6ETnbNOJ7XL0xVRQOmAYC7DAaci3i42r2bqv0DBhO+U6Wb/vUk5bZ9vTN5tM
cbzLzhEsh/mNSCcQ9p4/d+QqwVEqEtJNT8F4pDTKYqI20fqsk5cP80ykjPxuhph0
LD/B4sDHXPiNd7sd6KQ4WqjOvqTqdecdPDG6rY1kFsJayKtvRMNrwiURfkUT1y9c
3Yv13GqTgQS8qGiDpzys34C4zg3ofVCy4SX+jLZZ12BOplwa6qZ/JL7ipPYXjcWs
s+Df/wgv8sw7naFe/mSXjRn8/Fcq4bj5UIhle/SGkEx++Y09Z1X3LIZjhMQC+Iqo
aRFxt4BpsFaXcm7lsPhQLAtObgAkPhCJgYR50BDnvGaRxAVUHjiC0CXnVxH/f09K
XNYhuDMHSVDKLkELN3K0ptxUqjTSlonbfoQdI+fKmOHUSTx4K0ZqjtQDQ6RITqdn
aRfVjvn1OdjR9pnoD1Fk37YOQ0yspWLmLU60w46liE1iMykUBx9LMGcFXl5KMnF+
g0Bi+F7jivxMonvWqs2bXm7IeyNmc/rUlrY8CYDbHmTTfHMNQJCFKauR3svt7jXN
orjIHXx/yb6IZ8hNGCxqBWxw68lqy0qP+7u8GYl+vWlVmpobEWqYHTeXZfnLTvyr
0tNrsnxHQXwuR+1fpE3ZwMGFJytsn60g5sjLizyJEitLRgk4Bf5RbqwwlTKwCarr
ooLgoxwYqwyZxOnAc0RtNH/sSf4uqtvfHaeK6S5Oi7z53OIxQvyjoEMAAsJD8kp0
Xl6UipNQCkespOGyNi2W21s61rDc1IZ2AI6o92sgdByoEIjnkkRQgyImX/eSA421
sdPRvEVPcUasSmusbXuQprmioQ0ucxOinfsZfTeLqSk+8K8sTTfPgmDZ+6F/z5q/
s6fyBYGu3zEeSVncMl/kSmPO86FzkLjHLS60lXchdHXYF4GOtmuqJCTK1Ei0Qzpo
VlD464M/QfU7up7fsnKf45FWVEf2WkQ4FTe9SjRM9HI6+YV58V/1IAsgI3Rl8mFN
jGX0W4ay1EvzhBqMK/S1auDPDArc3FRoM/PAU4+3Zt29F7YKGO3GT/oydk4J8uu0
KFZBLtDwB3/qqT8gc6h9cHyedWa/hXMc4sjGanN5fz1LY5c+tV1fTVV18LVPH9jM
KwsZyFOldfuvhXQq8BQd9UtlPUUlQfdLnD+PadUTfRohvBkiOHWTm1JyXTCFLj8e
Hu9AqEaOJCc8lkSwgkcYb0WUcdmP6lsczXiLS5uIAKviVI3+EoxyyLeoQvPF2dZa
0Pdb7o8KHcARi+mNB8EFGVBYKws+2U7ZfHsKu2oaAVxwQn0oHd0fLfoqPtuBazHM
Mwf9ml0Td1wOi1/TKhiCX5awVrxa/S3EES5xcqTSuB+Fie2o7XfX4ksh4Begj57B
jJyNsGKB6DM1xJIYhzUwfpoAa00h/8dSIZKPEPUBR6niEb/e3CP7tmWV7/PZ52x9
jC52QaxjWCNla6yoiOF9h9ox0a/Pjy0z6SoXmxzoZtP/NoGHCnx4RoTSk8f+cWVN
60k9DRICMFi8ETtf/ODZViJGpfbgIoOvtSXwDLzHRs+yERTO4Pj9GhJb3fnFdleM
WzvyzmUE/JeV0PWlf8fX49ItZiMO6DD/VXgJBPhvPaCB/CQA2m9orblnBXcrMnRE
DxJbOwMwsphjAWL/yS2ZGetIOcLk4SOVgHPExjVLTOj+OKDzRLZEV/e/T1hns9vK
dLYpRQEIaJZy5s+zIzhNVho+dswapvUozrjebcZdUbtBBkRe3M9hqKpoKs/WO50f
f8Kun8t4CngY70hNk5uHVY/W6M6HINliRrWzPOk/RbbWGh/ayz7KQVXmL2PKaBoW
K0u3s5EB9v6Gtc7+qeYViCD0mpVIRv2OQYmpIGuUuQ46JC6s5u92vxgRZMMcjTta
xSvJjbcqS4w5y9YMfc/1VCZLZAlG8dZHRnpWsTdKkkcan3iv3EQoZCBabNPM4ij5
6JsBTxSBOjcOFVKLZJ3mL7ONK3bjXpfDMv4uogYaoQalGh3b7DRyX9Kl3TSgLxiW
DATJ4jz69CWLWoT0O02YhNE6tMibJP2EioigP7tPNm/8KlidI68hqxv2eqR/B22s
F8UErHgsx3cbY9dDlx5OZanrsjmUPp2MLg1bp1N2WZewzfh0k1ZTWZHdnU7JGLF4
8maffu8K1f2OrVYhwzYhATIA3T2q/762NuQtgT+ZDTROhboZIWhDEJZmPM+qE2Y0
3fPLawxkQQU+JEU4M59MO8MKL4U0jB3AFnaTclrPTLF0cuYPWapa+daBu/PEgDf+
TtuKnK79p04gr8XzL6kS0z3dLGv6RzOvG6ac/pW7GPu9gIUnOauboPUXxvlCLE4Z
4PwoJP2EAdGYWAFLPH+V1tBAKNH+JQHoyg+pWnvGLmFeUc9h1P8EwW4RpYrco4df
q1/uOiQlnm+UXF7hLPgmMRnvXLPCyE9W2fnAI5GKdKf4tpXwvYOzuDNVQex8rwHh
na3RJXOoGY16X/uFyyuuUi+HX73n4P+5+yLAPTGrqLkYIJiWkseBjXXEJotw2LIz
lzuOwAnf6pZBSYUw8K1rWKWYwDNQxmlL4GyYX00H/89sFonOReqXB8jasCUxekc5
SBeZSqLQqBLJTZBxdGb4I4V2zyljSWNn+QGyB9mF4ZCBCMrPeBVrEg/8e2EyCfLO
aI5uJlneUH9fBOYpK+kFzd3btOfUvBl3nUl1Z23p307A1SCyl8mxnKjBZlBIMAwo
cxgPpyKpERxyDg/6uljyO6VbEI/RMv9UhGfCagTmsEFw589M8SUFMedrVRAglra2
BoxFYFOKY4sI9boIwZI+xPAUuxHvKenLMQcGeHJyNZ55E30mt44JxZrm0zEiQ4G5
oMf/db3XihpDVk4tMrBPWh49okTo14WNpLjBTDOCu0BD3cXHC4O7p/KaL5+qJ0S4
q4dr0Gt+F5cZK+64oaOr5t8ERtb7j0ifDjyffzzC4XxK3FyTrvZc3PPWCHWnU1UO
4AavmA19WPbO8hNa5eUKCxSb5rj7KnvyxRfwrVu/2KEne/gXnZ5mrZA76UMYO6Oi
2B2W0LUQtRymyap2B8wSlqPDV2AE3AC40wv5lddC11pM8Yd6JRzOKH9cnic7l7m5
+Oa1Pj7CzYZ2iUXjCegoYF+zgOvsU5LqbJBcNzo8nVrsff1BVU0zYeLZRMxLsk7R
58n7vwhKwC+KCTKW9WR6HJ8v/8tCDyOkG9gp2E2JlszS7tNPk2i0uB4kB1BhGtKT
GgH4fXW9GywpX+8w4yr/WSV+Etd9hENhFSlodvLeXcPvyCT3u5g8CXPgx1cEQiBt
DXCxU8cuiXqPFbOivBeqjVzBq1SHFreoWhu97uFXhU0CL8WDUH3xb/TXVjT0MZ1a
sRPMQ7SU4XPnSOCanGI+nKTiELb393X6InhXrkE4coVujLyFu9z/BVqd1czaEgQo
li/f23+obvaqnzPoFph8CX6lQBiSioiWb4tkuV+zt+/z2E28WG9iPdvsl4RU3uIE
E3rYdcB4W9GbQ1kkcOlx98s8c0ztmjz/rQKNocIQiJzwsmrbUG9B3sNqX/HQxqlE
2iYjDnSsIQ9gMhmEtbWPtfJOHRnCcWaM2r9ZfjP3oZgR6hC/RmEtDmLH7kNiYgEg
1W7Pnu8TBmJodL40ac508HVMrQqa02DQgLCbLrI0B6UC/z3+8TMOuuvH8XjWC2x1
dNnCaA/Ek3knWCk9mOsSYTWnlk8TZQKrAZD3+MuMJvfI+F5JBSaytMSVMUF6ZlC6
ZUoAF8lMzyCiF3j1UCpTGsKfK7ZAu19ksCfk6vEUuynwyVQks0vtalARHSUTvqA6
64ESFfxBYR5XDe2Cn/0EuGbLo4ejYQJ+i3P6+103SHGD0Hg/PVXohs1VPjLCPIpT
KZBSyYr8E8WpAJcvNwrnpAlQpfafYf8ts7wo8Z83h3VxPOkXJmBdON/M29GENpet
+5YkacJcyRfY5ipXginYo4AroAkzbVRhwltB9eWRlu8acMYE0Z27ye9D/xvMhxUS
ewXaXQr66lurNUWBBFpysTZrZA4ww707P0vFVwR94c67ItLcOpLDX/5bguVOb+lC
gQ3/3EAWa+sSwWYDDgzDlTPr5zp44O7MKmLKXCaI1uncg9CTs179amxbSnxcsQcu
ObFYMyzJ1dfcuT/PYhis3zuBPCDR3bg0ggx7G1Iq8ek7TLF9OH0AfWobNlQyIo3S
Kox5guES1/v+fMWpBRCn+klUV8/cDuPz8hykKBnW+d+fAW3Zf5Hy6qlcdZpoxSzU
7s7N/NA5uPPdaue0s/ub8CBcFC+UlKmXipUTf8oPRuWIL1iZ28/doAGAg6KFBIJ3
fNnXK3VBeuv7FzTFHnFWBHEs1RNEgIP57hBZV3Gd8Kqy09GyxX/TKHuo2ew3ztiP
/+a2by2+Vw+Lqxattmv7awDzrwPoWvgopWuEE4dED0NksLmoUow3tdZ2hjl+XohT
AV1KcOOGNQyHeaqFSkUE6IEmFkv2GB/320uuVv70u3fY9ZEVCDkikie8DOfBZX9S
LST/RJUj5SGoAVdweuD1aUW+vtOahzb6u70ImHrHc/nzeY+uDR4wrahAYhU3hJ8D
hLciJCJJ+AsRNRhKBIVZjeCPT6sWB2n2CE0mRbszhLHw2ZKUTPn5IbjW0tD5YT3+
yzpcrASe0438A1EICOh6Iw1y8k30QZhZ8Ghti9PBUGcVHk9Fr7mPodF5X52tnmT6
MlT+Lvlb6CH3IOxUfCtwDVlYxqiSRgkuGF1wfelEzvVtJgIvoRISY7DwYB5eCIf3
tR0B6eCE08OuQMba+ZmOBmFZCMPCUm1QLlKsIG7cGBLGgRHSPBn2PyLKZPe6AxPk
lCkmKDOMcD6GaiNH2XpKQ4zjAgYgYZs3GwPdoaEuTqntN27X4CtRa2mZ1ov84iOx
y/k8Fal/IUtXttoDPkG860+ud8NWHyGqAYob3sjUrq2gvYHnGEO4B6aDqErekHeZ
zjlx/66qGRPMnXd51t5v3ccSHU8TJqOATxuhCibwFn6hcnarEuL/KiSc6mMpoENn
dc1BjKruES0h6u08xbT9Wad37YhKJ8G7eosoBu+nizuRplypsYJWwqKMnLbfe4Rn
hvAYBaNY1MqKdpbVN4qCLDOxfODju51/z/riJ5AYTik332G90KsPWlolr9AjFGkQ
xasIdcW3Qf8rMWTBVV2oS3lDa8RtEk5AN7927gnEw4bL+y4I2j77JuW0Y7zIacJF
HTEcDs6vvIdZCqianJpsjJ/yeL0Un3ocH5bvf4C/KHc8XBpJq3O6ZlUFj+02EGxo
Eqel/bBfx+kVD+3PIDySgEeLg8ldytBC9zMxTZc5Z1Ul4LzzP1pWZL9vnxotgU9a
MUYGYp10dX7h4Sb3se42Z7r6UB7aY5thYoxsfqIVxZXETH3xeLVgV0rCvN3kTieF
nlaoev6DrQHCqDFJZghC6GLTe5iOcCTvNKvQSwuFrMlhONuLJLAodCcZPXhgRQPa
cQBU9PN4/rDG14sJ2GOfeDkGXuyEKd3dV6zStejv/4nHARkAp9xzZ54ARUD9T+wJ
JMr3kWGtcIdN+f7mMVMWmxTYKQBBGLKge80gJhgBoNm+zPg7eyOCTaGHWCbyBf88
EVJCGncSV777HmqohMlCWZTGEWmFchvCRF9ns77Hfabnb4OLpw6Ma9XnHzYl4AUy
pI7UZnWerceOky9UtMdSQ78ylPn977hpzygFWSDwjJhl5D1BNxd1xUvk/jsVFGS/
SntjDtxpRMV00acl5U7t7pZiCw0A12eU4PM2zBBan0YBHHh9DLNVws05RKqZbmG7
K//YXAf40J8fU4OkGLutt3QMsPyV+Tx2FKlKrUAWCrHNKAx4oJEiJaUa4OAnncE+
Z5DII7qESHGv6nuVDkEVFddhLCwPoJX1K8H9l+1c6zgqs3qtHy0rCQoDjKJCmzcF
PeyMh3EI1OXVFm0qcHrFc8Nki1tUdhHe7Zo4irond0fncfXEMUvXH7ccgZgLlfmv
pOONJjoR20BBDLMkx5M35+n8xh1wle5nC6fb3ERGyQa0sLdR3oi5z5APn3BCnNuo
1icqjzFBOfQE08KNY4Dh9GCg1U6Tvhzo67H0/tJDoio/gEvrtWZIM1Ac4/SUPc+H
mBqpjAgi8+twxl4bgErZDZPlfySnHnvFVS72hcBw711JZOWWGAWLtrr0XCswj9SX
tC5tcs4DqLvo5dVR4PjtA74DmcmAXK8WUOYW+KgjBbn1IyxlC2bB1E22bz/bKWUT
Wcz4v9HAfnR1r3/ulquy4piNLvMh6B92F9LR8fmK7yc2dq7jL2+vNWrYDFlSaZaR
NLi6HMP54A53JcEBRGjAPmfQk7Bs0uVCAu/sy7Xa+Ysk/cZHyFbOQLbieCkQLYnB
vo2ByjoXjy+TrFaJR+2VTRqqALiNTnG4UsElvrwfEgNc44WaBXCyG5moByzyBClH
+8LbmqTqmQa/HgGg65rVvxrDVhnnNTWznpO4xkPxZmIJG8d/3Q8ipnG+QSU4o8qS
RhXyJ+0dKH9Vr5hVLuOkOIeDO1x4qF22JRmLosZ2j004rt4OpsB3GEczcC6/pQlm
+Zw7ig6LnqI+qokgzFnmDCuYpL+RRMCO85h22bSbNNKFKP/vbH4NQegxf7i29mCi
YRXmW6J1bBgo7FirzobwFJ2ZAT1g33j6C+rhdlI3jXly9RWsQ5fYM/O/oKTd3tyc
qORiXZ+b5KtG43SQGB7jDJczLf7XSdp2qCSbbJuQGTOVqFSYx/MTIr7c2+9RZ5Ga
fw5juZOSDddS+7eqPlfB92j8ysV830HI+OuekMtDxpAU5HBuSDe4V4sp4lcV5ysf
5b43s/jfDNlUWH+4MqrQaJfRXnsWBl1nSswyuCxE/pZTG+N6AH2m02yUQZvzH0nb
ZgxpohG2aYSZI7DpauAJtZsk5PPtzIc2c9sj5IYBJG1uOyRXDrSRER9CktLQJGIW
xm2r2EmDjQvQceP7+enqVxSG1meR7sYP8Zzd3hduUYylsVQ/9KeWHQaTknEbkQzB
SORs1qB+e9a2HpwZi/+75gZJYa191viXd3S9kWayjOqe7hsFU103m3qMvcKqmdJh
HcVANHLJ8+C+Q5KsMtKoVvnWiSG6FAbq+TqgyW0jJkQYthODFURWbJmjxejab/1f
M6yD+T6sxnwdmlfam7Hi8l91ELOLXnEgOTI2/OeCbGeIJCZD3t3aALxh+6IpmkDf
WsxPWYgfbMGdeg2bH6SwNyMU8MQztCWnTVVUkX8JFxs3pZNCpYhVIrRnrZUaqXXH
SpTGKSSrcSiiC9F0Y2KqiTAy3ZgcOUQ5/AuoC4meN37gfZUYyZwsmkG8igtWOHOk
W9W5P1t80Uf9Z4utuQV97JJwPtYqwnribfa/72rnqrGgUp1pjrrCyyC30Cc/MUqQ
gLyX++dRQxBHCO7qAmdB0FJcbwMnl1aBtdT9kqEXqG8dPzfvcAuomDr1JMMLkoW+
nbseSQvRGLwuhmcIH3c2Om4glPAOlzt8UdPsDdDyBvG3C9gKPS8TmD4/os5+BUsi
As/JcJ3serM1tf/irZfiSJWtwVw6qjXxbxs5frwEVjaPw+rX7bjdN/tmI75X7XHc
+BA5Wc2bsi8yuYXUbPfn5HXuUOP/mwcsgXPGoaQme0m9tk6IBYl+G4VX1U88G0nb
nmJfEPFGYxvuCJZV2NTY+qkdEzp5DO2EEyDgCuaSvjXc8sKbTbhL2tJdKUhLCR05
wWtO1/HNJxr/ynr3Zm0Z4EPqhr6OtCJqImmpiM/2q/E1EGIVZMJb7mW10DMCKbLy
2ccx/ZF/27sZjbJpPmrFPFNMXojWbUdkwREhk5CdVrYFiNRMDPg/2zuZZcX3BXDQ
e6yjrK/mk4dZ1uXQ4CIcg63rI+2U2mnNn11ilqLvART2iBj7wzn23qCDioHoDuj8
Qklb8SBljdrh+oI9LlvDypt3KaWCZ4E11XIR7uC1uUM/Acor1Ayy0gAPmAe3QCzX
2pHVh/Fh4UiIaClXdFPJIJsV8jYSjdfoTPLRRxGJt7m/BY5gzmJOdsakWzkFt7Y6
TQq5PoIlke+kyW1ykZdkkAi/I06DxuAkM7nLtFOfrU6SkrYFBHfm895GbEgaQNUu
d/7Azo3IKbL5irC5w5yh3aOaitgrCUs9XgMNj74tHfsmrClZu4WBg+dsJLfoNdsS
AYHxtWe9jRLwsJJzzlTm1xWqzNxdHeokQvuE/XkW/RuzmOGH08i3bJYFNOvDD7B0
hCF7GjSW1kNe1zciN1aOcyL4z5J34lwrBGnMUMtn8EPQdIvtyqciNbB3obwt5vYQ
NJ1k35EMEaEL/wrwQqwvic+aoUYMvYMObOTLByw26lFGsoWE2gTLWv9Qf6H4+GK0
rNLKhdEWjiyetHXzXiCkvS1OTjaY4Bs6iKmilt3VFY6zKE2LbI7oaScIyGoBJCiA
yH8Swh5yjhpxyZ0QHptV+qh1Rcg/JYf7f+HfcfD/bA0snkysTzy7V1/YZQM0X42d
vN+E44UKHcDtQ/OLvYUdE5tSob/nBoyBRjqFyZ+uRXUuUfbLY4is8rUROielVN8M
FGSbR+V5yu3yEr+gkD5O48kQ3KNCRIvfPKbytdLNf0G6G2Dr+v+/C+T50UA3g3dB
uNyndqyMZ9fIBZK2WH8nfbnOrzjsd0O/HocmHrzdrawQ0dzWU9AVeWD82yAZHaqB
lmDXP7Rw8YbjBGXlDWQ3N93xnLCEeRo+gdcKzfjQgrJTWqMXxLawvxwyS9hUmVyF
bKwXqnZQHzYwMZZx1WpLDjlPa/wPRm/U1TZw4uQTmSuH8JvkH1NJKaXaq0ic5DwK
t7AAg5MxbSxSQsGel6EYoC/Xfp2JouW8Kmvsz2LBQm3Y5pxDD7Y44KNFR4XLi4aN
B/w1w8SnncqyTQOjWsd8efzYFl2+l3sKq9wmTalzx+L5rE/tzfNMJedpPweoQNqr
ZBesT/iYe+Icd6tlFa0Ohmlf1teyk4DzrPXwsHObg6v5w3OwnjB5V7sysutHmHf2
VJMyokzcy0Q0bC9XM78IPIJZoSeZwWhdHmMWZaywZ/9O2VgjFsUhNa0XyvxL9x1F
qC9qOTBReFcI7XlwsDsAqwjvEBaAzo7kCMRkLz9YXXm9j1MvIQPjiE/FMSB6TALw
3sdCWcjP8LgxP5JqD389NTNaTrFDCganeQbXE5xrqT8TzHZpEBvb5s2lXpUX8Lc+
oIP1z89eob8gu61byDGYmxNbp3T9CONgUpJyUXUSCIAYzsheiknSEWaK6uj/aQDq
jHlpa39nqt/9BYbhuhak2B7rLOrwW0lOgWIrLgSNPkZNnAMxujtxyoSBbCwgIUcU
Xh5hI08UCiLDShz4ETsrwi4jbENaroP8hmDkcgdnO1LclIyJsRzgfV4M8tWmU/Du
dcc1w/GW83UACl7zOYOYGo5WXiGyHVZGS43vNOZR5KL2w/ViECUjMp1CL8h9N1hW
LVG+NNDj4lI9ADAC1L2joZborhvLmWLhayH1fcwLMMRTmKEnYmWzkDz4qgQt4zfg
573POSOYUVEJitTQFXc3EnljMTung0GlZlMCChBsvndVqEpimTbnXDgvL0+oSIna
WO3JYJAg30Ra1DXTWeZAWVr+gCti/T8Yh3YOdpENpxcs+Eck/GxM4mSpy1t6Tpiz
Anx0mVh0qUPWmktHduZjQqkK0TIIiWH4lrDvPh41z5Iz/xpi7wCVEyPQYtUW55zf
ZHV8kkof4wf+pK+T/EB5gl4oEO5pYBWvpvI8QiHhy/T+EwmH+cwLFQDbgP1yXSXt
8X5fFzdg2fOnNQyK2CldeZY8TX95SkUhJm9UJf1mo+ayztk9pyScZbpFXRXDNroW
7Bi0ZYOj+ZSoUl4OTYwXwjvgL8uPWr7DHT07Pcn/+EfKNZhQS34R0eYTZPEEGCZy
AmlcI6g5TeN8FotUJmFXV8EC24CsZLqYn2rrsZHkIsFSQx9Gfi5YEXQO69cm8YDU
T4DNmf9R85cZVcmU97WiD5+ybCzBr3snNY2EpNKKdhQVgMmEy/FwIGMIz0gIRcQg
0QAG6rGiCU1RrYYrBroYYwdgyWIswJm4jFoXoE1bKR1jw6ayt+kTcqzyzjNh1kHG
EP8TVIIk17gPO6e+uAY8sDyYSUtlU+2H2oDOaTutvs4wGM2PHIIp+A+KUoZ6w9M8
Lnz/7Dmnh9EiBVKtIrReUndj2cHpMwBwVw5LWZrKcJ7gbUbjjKwS6ruYB80gew/d
Z0i1m3WR9XblhyWT0R7zl5Mi4wdvHMw+KgttfAcmgT1YJSOwfXAt7G+7L5c8q/oO
wEM3DCECJT/asR/eVEkzV+Nv02o32eDJ6nq/dk2pMQWv1v53Iq+lXWqoABAM2aJZ
/3h6S/2N9q0cKu+bzsuxedGYVLqh/UNz0wXj1oqNcPSw7GVnedov8Ptcfk/ci/uy
QgVYikfoZnpB/TOg6HBFfB/JjTKnhBURS+yzTheX7LfTCYAzSX87GCdARi1DI308
IQ6L+eTCnCyM3/PQ8VfGrgKEHNhX2QdwDb0wR1rWlY8MnX7SYysCM6gubcPNAwA6
gqiOkPAaxIYAScBhjegcV8dvupDgNhwOEPKQvUvjQbcGApTLiNnKJplHY7nJkcig
mCR1IN733+W/ROOQjWGJc0sUR5yjKmsckpmsvizjUZ5RtdS+4WtcVcNIc0DdIEe/
wR/79PgkZitds0b/or+v5c/RktTQKzo3lL5xORsUHhIA3v973UiabJZfHNSNkLG1
zlzUYfpALaw73w2rPqNFa+8ghxSjDH1l4qQxY75AkKZ9KDiwq40Rlser64BUpipC
HYUY9nhqsigSM0SIQnAQpAjxsAjhCUXfFtjsz80Q9R54FCqKQJRVoHVv6no4Jjwc
DX3GoAMNxdCWFwySeQdFNe7RRtTcuHdnh6pmcIZprEsNbT6Aug+/x6z4PW1IffVa
kjEfz/VUD2sHXRUD8mOkpCiz8nRhhunC5gsSSCFgmbPGtVM+jSQ8KOK1R0zIRLKe
JFVl/UPvs+RIcG1VRXJRYjGedm5rtj/sPp7JGSvAw68iXBdsxf3om6QDRqBlnSGz
EcU5zZd7bqVmQP7j6zP3uwilgBP1On2DUiYZ8ZD5pY7Df44mEzFjkanrJwQFCuWB
Sew3EJcAN37NxlYgnrmIQsKlICpM0z55jwsoR0nHY25hVYe1KAjt6e0O9gzhxFBh
ARagBtObtxhhttwBy/m+uM+XBseFcXK2sc62E0c8KSPN4o2FHWAwURxm/m6Azskr
WVDq6dwUDrcTjX8qX2/ITMo810wNFpUpWOw5Q7h2N/AbvCOS9aSwOdO5lqsLi7/C
+4Ymzsz3MntCiweSfgAknkhnAO8AIwPoR+QFSwJHU7sHP4a/atw/OVjMUiHawzao
MhANIekrQ+7gDRmShjlJbK/0ICD4kerQy/jpSwqwdVUC2NalzHgQCADoj0I3Whi9
NvUjw1nsyLQowZSZdIENI8G2cz/LlpzeFqhtDbit7NFg6i4X7V9PVPD2bHSdWftZ
qAUQ40gv9F1an9xGpYQTlBSwvCr9z7iyasSyCnIIZwihvt5I/f/G6Ksg5CBOojfu
0MNCQ5qf1erOjNePTmWx47yq+8WBP1E4MJCeh5ZCDsl+OQent0OUJPGmzoH6Uyvy
/WDckkH6MlBuookADl8qD5hSiE1YbqXiscCM1CcgRANjk7kEKuOizT0Whs9eEs+e
bsG03gyY4/5ltstrklL23xo1QDYMxdmPOKNMDnW0SiUbnpo/gZMZ0mM1WeHhdQ3m
CK+k0zdD16dFc1+McrxvwuGBtEiq88tMb8hpgtN7czzVDJDh1v4gMwtpsIDZkR3a
fyFbvywnErBNutNtmLQqPHg1827ekwRUbrM16gpgB1fFXruQLqoiERG+nUAS2aZm
h5V9Jdu6ZR/q6xkX/mOHeL/+LS21yOHKsvuFuMUz2UVehUumCOB15bm+PHUCmpis
falEhaRs8iO9jtpuiHdkgM+iN1NcNOD1qsw7545vdLDZcPaTrcnL8AUjZHpk+LSP
iuBHB14V4stVOgWqyKMbrgRKA5WU2Z5r+i4kcYAkkHqbSJYcfZrlmRt/GpRgwjoW
tMbF7u+9ZB5d7Bfyhw2AuD2tjxXT6wRiEk40dzfsFg/63gU2/BKZr6CRkgCFZw4K
ISeJrBUf1Ti5wi0EDMCME7KOz35qSKvPq+2KJyQbM3/o22MrWuRhEQJYiqSAAJvv
tJDaoddTqc6Z+Ff5dtI81oJzVLe2EFsN1H8yBRGxQfsbWtl5sEz8uI58w7aXms8g
0EgQnTGLHQfVn+KF38BD0tfntiNJPFPnBsk0DpV84wwCnkATb9nx3yZHBzzGLogq
sSmSzNvpwo9p+0ZY6EzSVbySpjG6QK7qSjasFDAXzmvZV+n5lLgXjSfjDxonoPnI
RjIBjdmCN6hjmRwf9HVgkYG8uEuY2XKNIy2s/7M2fRx2+FeewyrUZRs6RHX2qJae
KKsn0tUlzJ/nE2OVqhdLx64Mppo+/aW80PziEufQKJy1VCQ/cfpmD+JC6V7HgEaI
BbglibrC9X+4unAXOndvGdMdLJc+RaPLqkObEY55f1Q5IMPnK3IQKToipk9l/b4C
vM11JL6uJdlWh2CKSlR+loQGlC+oVDQy4RHl+75F+FPOoo8da2l/OQ/crUjRYWKL
fLVd/Uk4scN0v65rXPvkJnPwF/Ad37GAamU/Raw2Zfd1M5/v/A8CtqpLqVyE5Kz4
jWh8wJT3K54L/QJ67JON4IUDQ29gbqRdVeF3p3qYtzuqoepXcGHo5o0VQarR+GoB
KPXsb2ANM8fGO5JPzt2yNiLXkuRe1ExR4Cch+FsmKfbWUlr6KJ5ATl/XBV5q0pDi
B0i8DEkXUYEazYond8kcxwB1T7dRFlox2y3iZTOvFCHmrV1a/ecAYpc4eJ79ohtY
r2SyTCphvYnhspoIHRqmz49HGMunV3Ke3p/+Wb5Nk8Q1yl+o11EPpkdONYSYuvK+
S11Jv4IrbgNHfMTPDsApu406kv/PDFgwoU8Q88M8czT+b+kS6EWGguf0yCnv5so6
BIN/XkgWOD/DYVd7k+ZLPVksTpTqe/UbKJmAbQBQhqUm1aGf8tbqtvkDBpWau934
n792SBI/8bntd1gx0PD2OSijzRDum2Jw0+YKlu5/3nyt3srvI54QT5UFw4tB159W
IitJhqBlXKrGnO2oO3dFspeTSeF/TMlYI131TioAZwzKm4CiNQASzHOqbUeIFhBK
gG26IlWeLjdmoP+KAo7K563getY97qMK+I40DdGSt1rZ1RUuTGPMlPUoVeojOzOo
J1sxmGu0JeSxXKiZB5K0CbSQnikwTe9XPBQEcKUgFCEtNObNtzOWZiXINvTwG/Oy
PRbpX/apjF3bJAYg4PsJ4pCSwsZNUCwBR1J/BHeorVLr7SbaYvjv22XWZIZ45O0P
5wjp/GXBeSrXHoZk56Ce5Bv2XnvbMfpXDpzBa3iCGH6ouxNcd2YFYuNwIDyg7v6i
sGWQ3pCoQ3vv+7nwlbLk6dy3SxegunZm/PPYKuhcOEpGYhsXHA51cqNzL4hCXNU5
x3EW2moM7/w4Cgwqthm/BeD0G5Dd03+PC0Y8AET4HsbjznprrspTcOdtNMgbWGgn
nFk04AgXDm2WzWQNnC5mSf3aGuJybS9xqt89sF8UHelqCFDIbG3efMKwAkHRvQ0a
u814AmcmJ0gSCGhQnOg0tQ6CsoZ32RL2BHTKwomx1SMtM2+HiVRUpJ7RynPMZbWn
ulhzggDGzsARq4ui5oc3j20sE03MX44zFQQh45sZagoHAeHj5GG7iF0JXPsIKwm8
YP8XfszWaSO+7gLHi2SCu1fAPoMh0TZysk5bo4FRgrK4TQyKBdwnAr7Jb5a6WEgk
SgVjh+AYcwiZLu5gDk4qbuRh54EI+nwq13mr/U/PJLsnMqIXs3ljuHPacvzUMay3
0QJOfZe57SxHdL5rKyzb8swXvvQWuz3UESzt1d4B9Ec9sHCh3A48XlCUU83g4iUs
7clpdJ/F1mEI+fhLN7ee4tLVZAzi3ri4UNTUFh6uErIm0s8811iz+KHCQR84LcSG
wWFOkXByTxuJIq0K4C0XGL0YpBnxQ53IJznhkzw0C1gzCg6X1c0sOO/b2r0wzo43
EueBANUI+d0UNbFFA3lFJgVOMi6DYwZwcTRwmF0ktC+5foL4pVcZ6RdYpWIH464i
ymBks2aojekfmiU6V6KbuLL8tmGCKIhLWS/reg0sgiLySO7hxk6Gh5ZViZKnlU+e
jgwKgDFob8Giy3fw5eja/UDqf2yTARfrHji4iMPxX3csfp5ML/WqGE7b4QO7nSP3
4Niuztn9oqUy/N3cSezhTKfCg5ijT4SKW1YNrUCaTSbGp98VE9Iu8QRbtGp1dItf
mAVUiNL5qfakP8dnSbFX3FPTCtDvCkb98YNyfNWZDKWvwrRKLFPbLn3jN9O27wzp
JOFVBQKBc+Y1e/5euktKsQKEcePgEKPh0mSIf9qxn7pedKDTZROwrV1n0dh4u8/S
4JxifIttxcdSRqRvCB2pePuuuapDG0N16tFO4AP1t0oJrYCnqgpn4g8I5F+9IqBu
qdYEYtmyz+71q27nULs7tTanSQK6EQc9vwSrNO5XsiBfUHuiqs0OVj8BaLCoSQVJ
FEePo6cmaeNRVLaEjKAfNocpM8mJX7zPXi8G+1ukzRhU7PeeOdHPfH8lw/1c6Jdc
k6ABSgCkPm/7yzlcvgRLOzZmA5cRPqCXmpBfYO/0M0iog38gRHV6Txl6J9iFW1n3
m4B04G1cHop8rjg88kkPnK33jnDB//vT5lIm4np894NyD3sFJiCCy3Qgjzh0wm38
jGe2F4mS9TNliFP4jSh9w66gf10ayPM6AiN9LON6p6ecmVaWbhfY9t95jhSGvc3t
LHoQryefUxymPctseCjTh4Jg+N2RO+OEQjrk2g3JY5Xyq0bKtH1FSkfGAuH0rMaL
Zx9ymec4+lKFnTY1kdpsTep/A8/+1cYfnQ1rfudPktoViyNSiisba/PNS7Wy3iBL
aNURj0Pr+rMNlWo/LOdHVHMHD1/n2rR00E7mPgJkrc+C2vqll7tOGeyqYVBzYxnv
VK5GgYP2H0NaBk+cKcs+qLbf9Xdu6yE5ObDPKnPTzjfg1C8HM+R3TTKKCbrV7wwg
PdheFM4fsfz5SZM4kxaIr3mMHRhGAOELutYMYUs/RpgNlqIQTdV0iBOgWhVJGUV0
eWLf6pkuYFSa9fZJtiVKSjYuQAzEXh/b5C7ICnG5Qh4Aw418Py/hWfh8iZXJJ0cL
TYcXY9wMIoajacUNPPCZsSc5D+FWj7uUr7tN4rYEiMUmw1vkQDd4l216GlgLWAJF
2ym1nmlEX3Xb/n6PmUY1zXOBWnK5KR6+WJcfg40JdNbeOZHKfkXoWt4csnjPm2cN
/iONTGP7wxZcEvkj+xlW+GnMjnAHoOU4yY/1R9935H51KVkJTUG5C81W8sdPPZlF
rnHsXoQUVMUmJXSYefxM8/LIFCjLBwE5MGc6D8+jdh9DVidsSVYEdD/Fuw9Thtlg
yuUnRMezZjYAdiavRBktP2t+7UMhrj0xIsbqaqoMygRSQUiyhMy8+BTuV3D4k5pL
QZc8JICfnMsDGXGlF8LpBi5i30U2w5ihdnf165DJrAeTS57PVJgyxFjS05NGt/Sl
78i8nzqk0/Sj1hrCq3UTvO4mheqziynZrywWPQ2DZ9ALkU5IC8SuZoxYv/vFeyE9
NLohtr44+4LvSTAGJdbwyREMH+DXLI/HV9FzdfXZYzi2dB9Bxt3MOEyqNS1n80QD
HFS1MeuhOU6f6MokOVaKRPAmJlsYq+EN1FQihONKuOewd3UGVxZcWdKJRhEEcent
htdh61ypGMCQmkjc89FpLRveNQMwsbJs1PBTWEeDf5ofqMdyr+kS3uJtzymHr+OW
RAoQIRrt7ifuIicHD+h0JTLNHbbuyw0hgn697YYgltK73aD0ODq0cVYz9QYyChWa
VbLcj+uyj27A7Cqk4jdENTE3eTOs3cFR8VqVvPBsVaIDOPvkpTi9rjr+Rey+Dn3k
zzTrBO1KC4rtuwjZVHRbym9iMckDYSCiaHM5nurRIOhdHaEzcFoNo55ei0SnQCeh
SBPa1QlAdsC1e2Nd78ncLmVITmSswVSaMnlY4o9+jiujJxKWERMgRs44nZRYAynD
zfwueoMGAfWTsOp9Fy+T5Rlyu4yTmszn3KYBpQVIThCnE082Ct8BsE4MM/AksATk
RKrbVUXPHoYe1ftt56XFhL0Gi4Ve0BuOsyeeemolD7UcFkBkXfwIp76gTR3KNkEf
dws8vmCHWvVKuV4PRReCw3xMz+2SG+KrHz7QUPjXJgMoFhGo+sCSe2FR0iwk8/HF
YxWpN54mghe1BW4q8IRfqvvwFXYiRJ6FgajUl5z+Q/9T4VC+6MVP1ukOO+lQXmsn
6ubxzj7xdp2FGneruwFhVWN/9a3akbaiTzKk8OuhBhtJMQWQUm6QR6/rP834bn89
MFrynT2XMDvtmeFESy8yHJfSBEf3O0gIgunamCSsW//Q3/oakGaDLzxrH3flRlZT
WABSweVXK46qlZ9G+pWjcd9nQ2IHo1zO8QnzQerUMqBeyjtvQzAclh/nXRih6KZi
0IphUSanBlSCrT8f5xM+JBVdbpzXeKQ5B8Df2RDZz/rU986RsGcNVyBOge8JG1NY
bVde0j+C7s/UyR3fbGfKruUebPXymHWjYPwDBRXJikelJhNmyfYzacsLD3CgY3zK
unKM4iMnQkXkE4X/yih6iSy+awSb7egbZ8hB4WXfkEEo+VauyGwoFqjciwaWkECk
/yGxdgzpGuBJv3SEZRQIUgY5VNFh/vTpmlKclG3t7XTDDFDtGjgucGQaE4vrTvOC
XST6fSiQ7+9wqxZyEylmTZsMaiIiAE3ow0aRuLXSO9KbkcoLp4W1TKFYlIROoGga
TEVKaVhfxHmiZKChaXCC6+Pk6ZQU3sW0ML2sWz6uqIr63AMD7B+ilLvuHXpF6Biw
AV4dsR95OH7j3UjrbR2TXjdCV5izPDweN2cy4BNG0UZ2LxqE6349EGhMJ7wpkl4I
bH8kHW5aNm21BaFenD2M8xjIkhVk0g6In2V2Ig9FtHhR9mZwOpKhKaD274exGLUH
180ZT7+riz8dfMcKkmpQdZM621Co5GTczsMzfKg/WS6+zajbntvISA7EWS3X818A
Q21ObKeErCFgN26mcMYIEBGyFPUc73G+5dUIOaS0Q9d/H2D1Gq3HpObd/M+LPn4R
Hwj7g6SLWhBqA/2VE68Cc9C1OowxXa3WJaF9uwI8V9tDQeaitNtk9AD6Y9f9xVIl
K3usMCSJE1TLKs0nLKvJCFlxUXVsNJTCF0Dm2jxg5aLjqRYNg05oYPQ91HEj875F
Y4yPYm0FSGXI5Rgty9W7EdkXsBmOGeN7ug67ccO6i/cfS3ZmnaXkUVRuMEQy/BEA
C+GT2vuqQkyQPXHRMNbPpwtV3mwkoS+feMMx23tKZMTuGz6bBD6Lnfv+gOJOqg1k
+yESZdkrmEcrriVPpBAbyLcl51dShJQRgl9W8w2i699x5PMpK5OrA4hPy/U39gWj
3hjRwlUK6+r4tB0ljrzEyY+4LyPLI/a2upllntCyqwtOvPVtihzkBQi3mAfptePy
jzXXRV8IcmW0uxuAfDf1MUH1ZApBPHJCezB+pF/xjGMgtW51wlWfLcOpJHuX0+Op
ud0K4J3Ub5JLr/WLOoPW64P09ewjat8LYbJXXLCZGGQ08qRY+R/9UBPN8eBFP3tn
MOpNj/W/G9UL0N9aAL7pXCKaxX4dOyz6zfoZb7oyf+Se8HDlXrwH3y8bEapwmMXS
8CYMRlDwfIBz82XCf9wRa/7J8cokrS0gQQ9dFdFcWkiyJFUprVvi6gBqxkwPf/Pd
Iep5E8BmtRZXO40dwSOompnNxh7Kzn1hdI9P8ZF6VlOj/LJHPL8QZRseolROznn8
ruskMSnk6j2/2aiXLXmQbidjSWeciLfqtiA0QEKtZ400k2/kYG7damdjrn+4PGX9
oW/9Rz7TPKVeJLBHZuLWA5nFl4QK0y2n38BWQdMAKhI+f4lZEf2VAx8Ze5pUaMRs
0usid1V8PtIvYMHzW7V0j295OFRH2spKrxs7izNejSbhdVAsiLlkKZ2EDdLLTLMp
xgRO4mT7aL7wYCmUVCQtdutB/ysxyrrpx854xqQtfjfcyO9J21Mo15YvWXQqqm7D
DWoFy+8vz3h1pS5zjvzpfMaDsGw5sQ4crUF3sdosrrn88ziEHWibJlNcUZcfgjr4
epNxlHe8+JSo9l4W6VnwnkwaMHd0EqI8v9m7lQMPVTbzYQB/ZppK8OOLB9rkqBlR
eaQ2mFB6A/yZhEkH0bKbLcrMmFKQcEBn9qv1va+7Z2a8Cuho+s3oQglPlu5TfxTD
Mv8q6KQ3esmfO+ObBbWa+rz6dW8dSCIsn0dDYyX48hYz8tRNJnYeVm85PIuZ80fN
kOLAEB+cNTmKqHKaOZNUz6FtMiKpsAbXZMqRKkh8Hv3TJcRlBHJsDRy88zb5hPye
7MX00d48LWHivuIaMueDFKqUGh8cdgboxAK83+gfM38N9DUYUflKQwbEC2ZmH3Be
fGxdotqMSJUeoohHMHwhSuTs8ryMwm6MD5VUgBlYMz0HAkWknJCgGBG6XectNvKB
8Xn2rbStpsEs1z+OfW4bOr17FpFaA9jujbQE/evR4VPpfjZf5ZdHfV1XUQzDwXJS
EhXiUIdHNbNLHA/7XWVpBGhq/zCVfsnJodLys5nQMWcYFuz1x6K7ZWy2le5+RXSw
S/AiR/pCgSlXhysQMFxilfCDubHiwOlBIhsx5/axGU7QdHqP9xsHvO0CITOj0hd/
Qv/yeByeuaCbSUX2BsFBUi7dV/Awhu7rGjiMoIhLinRFF7Gt6yhTCyXLntsN/MTv
5cGnFqV0ehVJ4gbXJdZbmwTExkj/FCzjlNjzgycLIp0bbyH42xA/WGR3ZrYtLa3O
CN1zeFHDZK0i9IKezB1p7CUW81lgJwuqNYButlkxN6iLKJcIgJLG4kZCrjtqqjXC
+XsjFSCNBOSO3WJwCI60ILcxdTbQjNF+hViwE70SCtpx8tIDDY4zQYCRSfx2uCrW
nUr0+2Sb/2t1VI9+aEUvmDzlNruWZ45CDDX2ijGsuO+FqpYSpTguqxJ53aT4bzfd
2gV86uVGLnGG+q+MVQL9dxEOw2FawOeOk4aROMNShSvtuYdRzDggT3UWueHioHF6
76Y4xPJDqyW0u71ZNaaVla9JZWS4yrmj5UYBhKfzbV0Tn9noucRzjxorYMWQDLFT
1gYwyC2o9AbC1O1cAMNf46Iq9wUJr0wNC/wgFBu0UfuV93Fr5GjO3nIXTJemuRLa
eBRMP3ecRw9JCozw4zXkdUxHGQV7pjHgFPdM9SA7ie8QMoF7xnw324YLeSM8Lo8/
grEoIv7gEoqMwLuofj28Cgu8n5S0qHQbMD7+O0umeJJMryyMS9cpdlGGkEVv7ggP
E/Bbv1vO0PiskRgEpe2l+7FqLYhxopkBpHrgMLgHQBuYB7TL4F/nKbWC+B9edy4p
ALxXo9fEuF8lEd0EB8ldIwMYPOxTVQ11mFV7edBcHU5QVi4C7nQ0z5VTH03YKlyY
HYwy1fyNCJ1diR32aEvgi+/DKU2LSY4AmiAi+UZ1or96MsAnWVP7KgbY/aYWPGab
QRR+JfAZsjOWc5UTu1ezCpbowTebNscWm2o3FZSBy3VfogDPztYI/kVnlkfULZh7
kzjMxroBIG0GL4R4v6E37gFJqmP8HKBOY4DtkTxiKwkRxmmSE7K4CP9U0YQ+Hrx5
GSIR4YvIDeMAk7I9EE1F0WLRVVa1CVL1LLc52VXJRnKyW6KGpr6DJ8kXAthVbELr
d6YI4gLCiNJaoWQ1r0Ykhx3uQzFzER/X8jWltG42X9hAzjTjyytL6O1orv9F38+K
6UHYSUSD+g8OlL4V5MtZpPojG+KCK704ZDxabGqeLiv/eweWlYuu65lN3QOo81Li
yjlSHmqTcwKAH/X+Sk/t+crgYBUNZzqUhftcuB1cdlPWsGdiiXsIO1+gxbUC/L8z
4mR1X4F/VFGRii0KECsw0LIg4ku+PDdL4Gps0VjWpMFtVSw+IHEIZikUumsqD78h
WEFnmzSTI4TGGkw8885wfCR9SltJenWUouyG2S/J8O9cxzsYRKL0UR6FyWAWfNn7
JeXjnykQP8HLwbMyHsuFoc1oIJK5WVTMgGjpwaWR+3InvUZPCdecPPVs9NcXwoL9
+sIsvbu7Zt8DSXhRtlQTWWFBtpwgUzvp0LQsEiqIRyCG+gs9y+RaPYk7t+EmnFsR
NQRw/CTwMLPC3tYn81btO+x+4GaBbaPz43CQeTbxN0+Z4qSvc8CMxCrixCfTFYPo
oIFtUNOAHiNwwvNTY+4AzopSJq/Qks+ynLU7Cq4q8pyJFrFf40bEHCtzh6bhwOKH
t/PyPZNjXkpoy5pY6BEHcH7h2RtzYzVitsfwcbp2f54zeslDYcDB42XBo3BEq+3x
gm65T/F/lc0hbgahcx1crY0ljJWs2/59Q+aVsbZrpEYHIBhnWCiEPUMh3huMeHll
ttzLwIGeZGgz4DAr9PLvnVU2UYNLEK3AcFsvYn0kMJEs1k4djQ5QGpepn4NbwCT+
sgjAcNphtiECvPAK00N87fgvD7vnK3Uh8FgGMZbNswh0fTJoLKyakYpKSbXN8/rl
89XnSPEA7F3tSKHHbCft/Xr0yFriVji46K37ubVwVr5WGZuA6JNSsTjQWkB55oB/
2//JvAWgxlff/EeKabCLiEHzUys34L+DDXq32TqHuRnt4YK2wjH6AtKq5t8s2lz+
kizvhmFuKHPGk8ET3Jkdx/uCexR48aHvlidpwrVn5JAYKVVqezKaLKzk1BWG3h7A
4GJ5I+GTyLGIz2OyPVvFHI0w1oWPcbe50qukdxNClRubc6aijHF9uc172uhS45ua
USfS2Q01zn1ER7/xKipOcsO4SUkPMayu28+fHL0sbdLU4RVx6WIVCnS5ePfjutH/
r9Rd8vFIXyPTJxEziI897FNPOQe3nnsDGRelJmsAMR2+FmY52U6EuJYKM420JPzH
NHfvO4BtUYOHJCyWobmBp0fGy96V8rkZQuDDSldVqAw0ZDxS5hMtvqIDSHnDGK/h
ptpZaK2x+/0LzYDL7k0YxrZwY4ydRGqHq0iLA0CXiOmm1u1KOaGPA9DRB35nDvvP
QMLhqBd4jVbMW7D9iBGQ7duUnf9RPIfKbN4m/olRVN79z+QWbn98wUbUnGOvWL3D
iS/o3DJocyN4y5lhL5lmV02QTrJ146HfqWE7ccE48uY6hVGLDibWup67nTtpDbSd
DVYIcPsL8wZD8YVS+Z1S2scApcJ3X5HIm+r+nkeSrfRcZ0FhUqEVmN4k39D3O/O6
Jrbj/Ku3Znx/QembU+zwmU/f3XpaMx/8vu6uJDkrIcp1dSfXmWLXXayhqUWO1YPp
Uzj6FnYoRNU033+8zR4hNcG+rpbd9OwiLaN48Q/Pif91sbgPUBs++3I/h2lvsVrh
lef1d2zQ1l+11ML+tVcKa5PP2ZA/2TZiG7MHR7iRW0UKBFSjYohtNY3j8/0LaYMc
NOQH6ZGNsKN3pTinZye79m2IFh+BFEKbLJVZtrFEGsvES8apuFjoPj3kZcr4/Wwg
56/LDpz7/3lYJvYoKvdNzbRxsjJccO94V4l3Qy+rzbhh74xx4StSZ2uG+PsyEPoI
mvndIumkVAWRuy7YP5+tunaZIrtQBESauOJ3tx/1ShpiaugEkEdloX8F6q9j3esO
SddKMAJSnt06WtRhxkSScqwzyuZfmarxIGRxFpaNWpzUxN4OnsM/4uQlWI81z7P+
uC2DsAJXQz9U9HW2GheaqW4Sxv4EguD/aZF17krmaPI3j2mqJ/lElUeqSINV2KjG
0lKu9DQL3y+RCqTu04PAFJIRclBYQ5qapuvas4OXFTO0j6oEsD/hJKjJ5gpGrWDG
lQpDnyizyqE4GtJyTT9WcS/umljkNI6btvukQkX8d3/exURov+OJklL4kj0JE+gn
MI/QkUcEQs0l3lZ6naDAwYWa7subEfHDszVsy1GFr+W/SEV9oTYVYODkGe9NRmup
ZIKRTu5eWg2XecDMfswQqkiFCiO01eoo5uptSM82RlAsD8Eu0K4tJ2Hwlnz63DS6
fjWGNVW15F7TsFUCHnokc2SJ8+4/VNMyvk80dDSCsOU+M9S0iI+9hRscZuwH7oUX
E8sCh95P8o4PajGBojD6fvvB3IoyJ5RjSqdUZYvGTUBWZr2+16mBa9NS+V9bUGwL
+xqeodEuLF3YORpUeGUBj+sPE+3TUdBFXzyGkSOcpuaiAOg/7kuphQffmSygBivo
Ekn/0voZMit+y4tTbKwI/XLR48XPMrh5o65aqupA3zjvqBR+G5jNaBqtPzzslpRq
HtOLbXjwvkUaACNp2mMXX8lpqGRl/nnAsmwHDf7eXKn8zjz76AC/OtwJhtg64yVb
P+CawRb+gW9xMfgKoFGDK4DjhPpfWJMSd/lqNPfl0Rns+gzyvv/FL+rRAYk3Gerv
7aYAMq0pIqRFdT6t3E6B16QwUyNNEMjK2M/JrsVrcdUejRbTarE7xCVJZRIuGIjP
8OMZxxEc6Gqjl6V0mC4wo9dPXcxVDy4YSriCn/kFCva5sgD7ZgMo41kWyBmPNJuN
3Idp1nKijv3Xb8+LqKiHacaOulyCBHgu74DfGpgcsslrGoD054D1aYv2+6ohtjnl
U06dzF2apekgdJiinEXMrU0zcqdfrrTe2T3Ryaw+f9pvuZCE0QPfl8aqTVEH3cay
R9NT4oYsDE2Q8SOV5B/d42u9pwDymfK63sdoTf1Ychgb5GAoHeRu+SLvMBliePI8
oPMZdWwvYXqoNoOX5I590qC2i+4VqolLKsvpHF7VYnnPlWjR2oU4k1HQQaIpOpBA
llfB8+CPSixfBgXVQ9Db9YzxAofAFcXgnOvVtO7fCglSbXUT8vmpkWHP2IHSFULp
F+kvjqiqnyaDOQpcQFbrWxNmvOYHw91+j3oh7rt2JJNSsKP66Az7CtG2aZIGmALg
hbjB8c4D/bGT83WPBLN2i2qVWOK9ymYU5kAfhOQvNchLjIDLYORwjAdRsWbtLZcV
jXhFhfKT4qAUU7cQlze0qOz687QpraJFVzdj3VQQUnkb7+WgmHrtCtxUWiE47/wb
hfLA1tDSD/ZTZSZ+zJ+OAQhraHMS9zhZ74CLFfU6CMKHOmcDMU7xPlZrt/ganzIO
4rtya+SGD7SdwwtIYOxFAzFQxtzR+EIjpJ82qHcM/dZkcqhjGhIRxqOfrRtEqaBy
kI1/vO9KKLTcPJcP37Fe2YBB6aU306pYYENquF2nGfr0RTPVfvcpBCf9IeR3u6gi
zKMcb320Z9eon+akuWjecPSnT7Tt+bOnuo6AwX1GSzlmxkHAa+tfwGk3xKsjq//Q
3uOnTszYXfJ1VOGxQR+chB7AooEyFUDSSegRYyjjUhBdKYrFX3kz2lOxEg3JTpGL
GveMzGpQIkNq19PNYqKaoF08P+AL6Z/AjUq7jToPVoojJkBh0K9z5SnvzQVPhXOs
iTpCTZQVCmCBInt3Sy75aQOQCFl+vLKk9Gmrfw7HReZDNUQjFc4Wz/qNGDznDgJt
NS4CuRtPGUGW7ZdipSZkvUmnD0aC00P+SdpeiwmcqJsECvo3lyD3+fgSPz5JuTVq
9mDho3FU+4477oblbYI7XNvpjBL/hRstFRVO0ecb6QrtAaFYRi4edNxOJCn5Cj/C
av9CBHfEkvWqbZmshQN4Sbge0zqc097fW876XzuIVl5UbqQgcd2xDcaFMWzQeEor
l0yhzmZ2TBPmnMAoDeU+8WzcLJmIB01mBUKsmrOH0+1ePBsPrfcVZ/NR3YvXR+Be
kJMUwiy4q2+Dw+ura62gNjC4QWWca8lON+x/bpUIu1nF+4QSE0Hd3cjroP/KunHY
+HtbqZFdp5oJtnxe9TpdpHg11LuvUgAkAmpZB6gVszgWpY/LXmW3XjpmEMppMp66
en2bgZQiLRA8QKiJ0iRuHh0O7Tfvx4xwqmobtgB75i2in7sFCdHAl4OHqbCj3RIX
MSeiSlSc74G8bMtAafTmRJoJ0Uu2rd6pKlKT6O7brbN2ZQqbc0M2m1xPCBIlKz6j
bhsCrprsMuLaimCr0gCGk59kcBZplXOmtsFdzJbXY/jMarxG46grj+JoCjVB+TIt
WUP7YIcykzy9iGV0vpfB/Fos2jVZf1KZ+FndK7d7fP2FLQgJ1mayOsOSuJo0xLd1
IZKtouWZCBBz4SlNRjhIaSDoCuhu0SK93/BjzoJN107p/e3HEIOLJzbiQ+yL430j
x2D6hWKmWwLgqdmgF5cgFZ/elLCiEBblRYUkPaoVPAtj5BiEdXgzBr/yOVFVGnrT
Fz2s/lnm5ZhLkjyfLVfkTj/JJDe+I7wTDw/dXalNRWojGXoJ3P7G3uOeDkKRx6NI
BsFiXgWRqgvQHDkzzqSxpblQDG/GRtyu2oy6GpEodQZCz7ODWL3DNzgPBhWKdoOA
zsgo3OyYxAY8tgOloNMGMoIM7QjQQMj2fwMStxXrLjXMyVPVPiFguEY/diU9RYNO
dslQ7tYVQ3WAaeBO/0kH7PAWOwOTjL6KUbXJdrrZRerL/KhtmCAEmtrlmLZPpME2
qPz10hn8jWJwuSmN6k36J05IbV7zV9DdU/I1ViWPxRFjRxfZRHIZjsXlwOAzuyzq
qEzZStf+AEreCoIhjkwNoQk15ATCO4hpbbasfRHbqSfIsMEqgevOdaerM9R2CGeS
3i5sbt9ADXMjI1rqmrXsNXPgOnxsqIRefRc0J2uSiFkoS7jmnLWFlmvDhKymATrT
ksSLk0tnETe/HTIurbocLgxOD0wNDYoK4q2FuaWJNQkyMz3wxmoNLXvUlI0Y3IgU
3da60+etBzUFbxXt8qKNZXK210rUPWrLY4cqnz+1yBbp9YpIEMH8LmqVXVTyN0EU
D1pfgoEiWljXNU2VXMk/8u/GWw17EJkNfyV3ZPdTx6Lf3tVhfFrRsLiH+iDXCcIk
NuU09tosZHNub9vpaXh1lMzyJ083smlDVvqzLtneu0pP7gvLWvrXw+oEJILt18U2
amn0UGgqUS5cMMfnPhJIUxkCPFZ0SFXZdu50x2MoHphQEOttIQBHaYA8z59HxCWX
ICl6b/JruXezFk6SG2lATEZNUFLiw7ydArc3OFwlGOR4I6CEoACbWoHrQ/gU/Rhp
Ku2B3UqjQPxrY/hPw4nMPD7jSg/an6im6BZR1CBJ1s65dB7q+tF1xYKl6S5h9Gk4
Y41/S5/qc5Ke5pE8VXPKtp3eAuC9Fzu3k+oFmA4fle7QTZZ7uZry/uNS6mYapBu8
+qUH/rtDXET6GvKGB8nVJ2oelzE9A4sM2JAWRC5AlYPM6zhTSADSPx96r/BiDI1A
b1RzeoflA5miv9Y7B0enRuDSCTCMttV2YeUxJ574yAh3IEfDpbuoDcTyLAE9cWL0
fxDbRG3a2Ym7Dx2TfAI8UMq7QdGwFXb8gBiNZc2NEv8sA5zOy8ucbjBvj91Dr1So
eSch2ZqwMcfiUlW36aHzBjQ2aax4E0PfnO9akZVChLOtDWrhjyd5pXaxitsazhpb
1cnThgai/6YhoKYSl+hEQzAgT2aAhRkLmPPI98u2E5z4iOyaZDv2aMe2DdMZI49o
L0CFkGpdBbgFgMtgMFscw57V8/2D6rQEq17RJC7MGDBHnQhITeVQ2Jmcc6zpjVtg
0kVmfIeZpm8ffv/CiFcKDxeT9TgQFvnob5bdHwWNhTFuPOCKYPwp2O2jWx12yeu+
hD82pOyczDaZN/4IiGrb536RMCyIUSbKxOiWNWgYtIq+F6GuFSs80FmWENepTUYC
mCx25UQi/OrTnaUiEsN1uzoFDtRtH5hueNdJnHffJLoe7neCRkku9rD4XNug2KTu
Z+IXqi5efaIRcf6vuhOTKo+y2hL2uk/emkptzYqI3MsoWUPFdALgXP7pYLIueTWp
MbnIpHmoZcfesJVS/pqsSAHzg82exP1bIPFJ/hhX9iSVzE1yLIkV2QFx+EnInRxa
bVt+nlHzIUqdLKo3tQI8e6QwFphllWTleP4tetfl8JzvZs6YDQsSCzt8B0/stuND
pgcnU7itLXxEtQqwU66nbFaPLTuiuqH9OgN+QKLxs8rdQi9Ud4kGEkZZFdSvlO6b
mO93UmLYUI8TccFCLIlYdMJ35Y3ngBuV+ng5O0c91xDeOoLfs9XaUAU9eofJcDow
CuC6m7YrZmjsYPC99f7vffH7dfP4YoFGO6XmR9QGdssfLjqrDcr4G+0SidR3FJAn
J7xl8UGJll7Br26g6yz8+AU3hWP3lTD1R2HNYklyBsDlM94ZPtbsKzDBGSdwASlx
5lsYpn8iaWQ74VzdQ4Yvj0dUh9j/7HenQy+GEt98E2lmzVeiXXoCLnsF4f1lm6Rl
RLXcGwo0RM29JeJ7v7bRuERMA3rXWje6E3c9BKJQr/bUUoPXNFqKITlQKV9ggE75
Teo9PVkoX5CtRUM41QYFvARE8RJoGsMfTry9QtFPTeQUhWUTXeCr60dOVh9Rzrsy
yqJSzNz9jhpX/gck7HbRZPb1/vZBvLQBhJ+Yooaq9LWZbmquwu68JvDI2lMwy4Qn
Hm6j7ZT8PI3dJqt+/cx7nG0GlzOdN2UlQJ7m7GMco5KucD/wRP6OPGbfPdIZk2cx
PK8YCPFgHNdLx+8rfiyLECS9x8DuW4EiWCIZ7NPz1PP0tMpQVSq0jxy3PrduyMeS
6FoRDMvtXE/WW3W8/a675Ty824481mm3UR6LuEGZ/rwzsM6WcZJ4GXqbKabqUf6L
oas6daowf5QHoRa2TP/koc67aNcaEKPX7sb6R968s/41x4tVoA9wRRMU1cHSTdLJ
OCt0VXZpC9GelUJXu6M3WkjRjXHpKS7DCk02kkoXFvc/MkK8zpjSHbZkFa7f445/
d6wR6CMEJjlCid/C7+Hg/f6WljdhVWd13HDc+BI3gNKUgK/kPlZUtd+ymFtyxmp0
4W86S7mqYN9A//mheX5POBQkKmbuoo2IMXBjlG15oDAS6iIbGzv0OjRBnw85VtaI
NmH/+hDbnLvbewOactEkrd/FfRMhHrvmPsx0uU8WbMdJ8d9UDuGMSsXlGQz9xCWS
3Ts2SIb7rtg5RO+VFFWyPPVmz8rJRUwz3ahX3XnHeJm6dKpZllsgO77lIz3VY6A1
tupC6k0/zcNjfJv6Ie5gg/CsM9YIW7xM8qS0xHrmTLo9qRsBBdexCdMLX3g7j2Ns
pb4e4Sx1BeS6iwRBk9tM9gAETXvkdJpe9VNYYHfcclkMIF2VPX9TmLeilXJpk8nV
Qy1BbXGn7H4mN8b5O2YIwDQ81SD15oZ0CbyVc2b0zNG12G+6IqT8Wq85kyfDnzuN
CqRdq43xngQrIqUDLYP20GIX2j3quVdT8Uv+Quo0HNqnA1F9lbH6VmYULwzDK3Sd
6RiCbnfZxmMTSx9BfCA94jYPD/Tqs4GuZieE3XAkgCmkG4cZ9SNsDgUi3JQfS5/I
sDtQH5fCLa8jT/6ggOZlPVdsenc+L8ibR2gjAlQAE7R0nUExhGHM73pxWABa7C31
4P6WNrpnxslt4mndm5zAN5H5qmTJ1Wvm9azPydPaNu+F8TBfDEiCSu8zXLbFa1ry
3BkRp2ar9dyTTwwNDLtPZHSEEjVnPc0TCw3Se/rayzAYIE8cOPOXWKRCSQFT8744
Od2rmzqmNZ6teP7cjWjGMMImRMIiA2DUQ0R9uNZkn3BtIP+9Kmx1lVAnMrBiOqaC
7jvaoFqeXo8rg0LbmGsfA+TKKtk4UgTEMb3bC4u4ogI24GO0IHCqiw/raHu1ZYjy
gdBt1Jt265SR8eLwfsqEzJegCKs4QnxTUJ2mEXXUv+eMG6JwOpnNlScQE4wPUEg/
zUZUv/4XVPs37FIHqDRbDDq2KDjWUVHgwYTYwKmMu27eKW9dOcdvJPN2AFMEWGkb
PEnutAS+wLPpIWkyhF848zsm1ju8jajg3v/++x+/vfxzfOVIR83hnwRIunsHTB7I
NNDO7QdbxkOZb2JxsTaKBqiof79Dgpj72d6nxXZhKFwKBW8vBf2rY0aJmgsqMspM
4fcif8FqRnAlMfBjO7OJEGBxShaIz7lCmRtJIlgjMOn0erTXDlmFH+cmBe55AwHr
RCwHKsCm8LpMr84v2KaqaqB/4SYz+Rt2i5UIp5FhladD6Ch7+Z7l+NHr2ie0x77X
sqseriv9sLQc9W2VrJPRMo5rKyTcCZSUvoWdmMxfq0/wQj6aEbmzPDfdhq2PoFKU
3nv3yREazd/jRAuJYBBtk6R7tlr/pxPj2/lOJJ5nzi2Jch26xdlPpd+YWbu6A2Lg
7NfvSOYF5WDLH+yXkSKLCJG7GCRe9MUvDUuPbqsx2+OsLiishPDW8uBDABf7XlnZ
y1Br8toLthGfOGx0TnT/aKKCtesoMdbpTKROCIM0IB3cJpT7ZRhRNNdssdsyGPzl
iZCTlpyBMYVkVqftZN24ukKN1nuAerxD1BtRGxf9GPkEk0fnJ4kPOttgRz9WmUOY
3cX8sOn3mA1+4mJQXu2/ZZh+SncK20HMyFOWW9o6YnInnbtEol38YNdGNbZUoMX+
MO0PtjVpIod3tVzOkJW8RNApUWoljVTTsq9BRSKVB4PPZGdK4DVoRorByFMhrXGZ
zG49+a+ND1YEhH9VgLBpM1GKgmgPDpGy90vjyGuskmdIC1BtQ+vHRxkpM4xQIFdp
MiLRftAZlAFMZsHwPcflQusOrVPK06c8M/PyBrOPcIReuqUVW/6XwDkEyce2Dlxr
GSFMyqUEjkewamvILAAZmY92Cu+dcWcIeDckrNlH5ZMHB2ipXDXaj5+/QKFmfmeV
Xin1sqmXDf5w7u2r+9iO309qE6zZlGf+EVKGLF62zmkDAa2mYm/fnZaMu4kacrdd
a2BBYMefUcI49gScYIoxIN/lrJPUzKUW9vZ9eqYgsPwbzQHHqfxjrIa2YFYbkrW3
zKl3Pf/AGbVMf5q69+LCalcDUeXOp2nS3IZSnsyu00CKWZSK6UoNzRSdFQmY0Im7
lwJ0YemUMa/KT9pPnxdHGU8TBummxSNqnzBtTVULp9gLm4IW18ZRoDObngkqH/e4
TaKfZXZpwL2ysfVUMpO78rOOm479Uba/sqe0ExIKCbKx80n4Oc2sXUnReusXOYPz
dWgUbsFEXY/ImOSqSnImvBZ2K15ct8+2Bw3tsLWto9AuMvOIVYV9OCAmwZbs4lIU
DmeDCq2r343F8jsIafjzY3tM+LzNOh0KeEjuYUVEzF5Nev74snfSWGWYqrH2WO9n
wk69TWx9R95JDC4YynBDtELg+jQzFM+gLN3VonAfLRWtvsUlnfk4606zwe3guJrB
2Dfo7UHiHwIPd5lzT4my0ds6h+kSfbSTImZ5YNRo0AVkgqUt04bPu8IHcfOq1p+l
asXjnV4W+wwb9Y9e/zPUhs5xmiHDsOEcn2/ZI20TgPkWHUffN4PWmCBljWfA7RpJ
s15lp2OdMnycyCBInZEdqtFBpwa7nNI4F8v/HE9c1uPBW4kcjHVUM80y1uybJhsc
u54FWurcf7CzXl1Xv+BMSdllLXX3as9wfj1vspUAj9Kno0yq7ntqf1ZitqHCcC7x
cr6dN1mva8kJB+KXdi+is3wtHMjz46SDOIljkSljb49FNcfjOW/0+6m+2z8+SiaV
/XQZHIJohOl328oJkx9V1lZcSf4QoMbe7idw+aPgxQ4wrTyuR3zO5JyM+eDm0Xfm
RregP1kbBFIGkV/dnxX/v52guj2OSRKHju5e9+lu5dUJUHsj+c32k79EK26MWLq9
oC0auDTM9bODdXjlx71MYfl5J6xWFTpuaYM1/BYqQFTRMxVkGC3yxEW22mnOTZlf
qW0dR6LdDlZpjlY6L2y+O/jif0dlPbZLbypWYO4REuY22EllK3zLVQHRFTrqSTsw
2j5NVOGswo8NdJDqRYS/A6co3U/MwkOoZu4IxmeI+1waRn4j9FE/AYkZD1THrzw8
4DgJF7PqsRxZScOinHj4MIAwLUvoVsIFzWcxim3iPHatFRIkFK3CpbrrcoZuFJzm
Nx3HqLkE1RfBfAIhjf5hcLBpxcjnu380S61G1bORM7rK2R9V75EN5gd7/Je+6QfF
sI97XYrcZYqBCV0hKdY9VpkE7ohgAR0l150/ZEHgQMNDFBZfsVsvf8iI/1NSuhH7
e4z98LVZs7LqMM8R3tN6/vvAClq3lxN40hDgaRo+O+mIgm1ot9mRoex6qqcsPwKP
gWoNgDPhzNFhbYpBzCWYyTwpwCsDApCpJbEizPZWqeDqelYYXCPINCWt4nTPq+T8
6auUqFGkfXgIUMpO3SLTuKKS0+n8Q9AFjLpLEFZHsd+3x3UHwJewEm13WK/f9Jm+
SbKmU1jbPB6wVa1JcejaM8mUNrC++nkHQZiB/yoZFdNBg+iNZ+5L5YOKYol+DRf0
1bHVma4qgpVMhamyLmkGLQQH51NO8ViOmkO2VJLWumuJKwG2so5ji3ik1wvPvC65
Thk5oE1V6bQC8Bwqk45SVPvNlQg8NKpFFaZID4rCjStmFWxG2IMRVoknhcEq6S8E
xTOvkG3l3QwRV/ebHS7H/Kn6y6X3VlfnA55tdlt+6Xa3KUWaK5tzlJvPrYraHAUX
XQy/hDpE0m+EgMpXjwmc7y/it0m8DZIWh2W7gIiwTTslkBPUirnWFL2WnpcLkjEE
doNMLP5p/M5gGNisSgNLEMhC9SWQCR2Z5R8aA9Oc/hNaK9caBkqjoOhyf5GuOILI
aZYKH8bg2TLPd6oenyT1QJQ0yfKBSyBK+WTcsd6Nt4CUValQaz/jRx/bBtfNys01
PzvQ0P8XGOWeyOoRxLj2aiCZo4sSDk5mb9nqRZesY9CleU00PgHrym3SdrHHjqj4
W4Tc+Sft+FuuxU1JGHo/Zm+gT55Fjn28w/QXaRgmDWKQrizPwQcQ5RqiCVSLI4Y/
g3Q2/u9vBCJ1F+WD/rwCsbJ+fGkSASWguNokM9OM9os+nco9FtNTuWnmd7yUYV3I
nqEfcKSwJ1APKy2VdtnkqACKLgAOT6r+s7dM/8zAOWKEhv8QUBvNpjNXg4PdjtlY
gVKrzQqT8r9K6MR/Gms5tdJyNlXbb19sfykRSbnKf+RWx9WWp66UUgTWK6/D8/Ji
e+oHywacUzE6cWRdNFomrUKkpQgYnHTObY6ZhbMg0JDB2cskd2r2/K1hSI3c2Wzz
qpbkTauymLehaVtMIEVyT6z2yDrOc/Cz60z1tvjPNaXXj0epMDSMse5xRE0mfLkT
5MsuxtCKB+XxcyskNeMGZu4mTWymazhdclNcD4jNuH5lxh8EuUdJHKP+cmZQC8/Z
lg3Dy7uUzh1OPvsvtSoAEdBSCRZRFpdsAQL4IsK7Wp7sk8ZfujEpJHG08ghb1sbi
V5vCCPlyZXQV3M1AWAOIlz8JriJ7BxrBDjv0dwjemY50m+DN4zEC/38D4cDDNKVC
gs+MIu/bsb+6vI/rTvfuRsU/Ds4/g87VagA+PzOBzkNN9jhoqOj32xGqhcNcr6F4
iHPG+lZSWs9nP3oRKoQvIJkg5GJWSub2sTJ+Eq2pgVxJG9pLz1d4720uKtClYVQQ
ttzQjefcc9ZoO8Kurotk7xM9CUdUYRvDb0AWS19YYWipUq3cdk9XYDqy7GIVBPgr
iPsZfj9JlHrIdgIQxR22MGhoUVQLGA/Be4Sr8dy5O4gXsOoeUwirtg7Z8VuvX8SC
EA+GO3OfGpbA21UCncyLp0LbN2uIk69HWUq50X9dxha2asdYJkXVBOAbad9f/avU
zqpXcuiO8oXP16k1WTQgSm6MR7mRFyETt/gK7svX8nW6xvU1wG3pS0FsvkQyVo+3
emuEUQ4bRcfQVumL6MZj9de6qQAo3nZlzhRjbDXYJ0geZe9qH22fCDHSYpMTjjLm
DNSbY4I1JvKsuVfwPw0DN0oRPj8JVrTSNOXYyx1+t7FO8sdf/H/EC4h+R/HzzRyN
DYK5gmeNb1YPG8pZVwSv4lt7ZqbBTHqsQRKskjRaCBfS9y9bnMI2F3vnHqkVh4fJ
yxZ+C+QLSWNGxJ5o5F/CVs9huZ5fCRr6zCvKj7G3KGU0V5qbBgbKEGpKrGKYUfOZ
YVxh6BTPi8HEAEkXZrIkHRb2aCPe9ZuMQCNAz/b/Ocjnff/+3dQEvh55pI/XtfB8
C6ISmQAz5bQcIh/XBcvnjwi7TYEsFS0c585HUfZdY5ovNRNG+10TuNixUeBzDLpw
I+yPAFMpeZ61wpkuBwXUuRlM5yYQQz5r+3yyxdgnh+g3o+w7gMNKPJ5TQHZI0O13
vzsOJtwBDevdC98Wsdq5jCKRTeo3b61hreT1cQRnfoe/iYupx525PV/gcSoa5kTx
udTup49qErORgIbQf1npzO5ny/nDIrdSHh0n7dS4jRDe6ahb60ama8x+6Af8gEvZ
NZ8fpJofNtoXjDZtGtu75ODF0vnq90ene+HYQv6e6lPTXmTeLAp3YDYniNbqBvpf
hLSvGAErzpNKFeLRQKv9i8NVV9qrVVpG1VLVlc9rbd+875DZYxaNHsYvaE8oJWre
JuxKDjBwBYdvgrPyqxowyIsg5i8VGQkZJKxYTNk3qWnx6fvadZzy7IpklCmjTJlr
HEUJoC0QuVK6jddNDRbTFeYfIvJL+7BO/1VGwiQisH0YoWHL+l0xr3GddvFCLSgg
O+tCeINnk0zDtBvXQrwNVCtEZuR0JGexetAFnq7Fh4x6xQw7qpIP4EmFe1VMCeLx
iavQI6ezf/9bAbRlLwIcbnSZ/aKl37tqvuPP/cZqVneoYOvwFpDB6Gkusm45HZW8
4pe/3vwxgvmBuJmKulAk8rzDlk2yv12SPUof3BpUhvSn7+noRsV1dSZOExlgNMTC
yPB9OAEPTcSpyc6Qk6GpkAsGf79HLqbg4zl2ISQXSDRmKgCPIWeULxwGV6bPNIVr
N5XGvk2b3mT3mZI3b6NpnAgK7Ag2JeevNQt4C7Um8hMPvLnb8tMo3qH1euQnEVGt
Wu02JG3+0gm5yy1OroSiy8f6qAU6yo9GugSNY/1K6L4fAomw8zg7ul/I8ZNx5zk2
s/27KUhhZRMB+doj79rHLpi+z4ZZZCr8jpIL49+o/un1rTw8itfsAz+ZkSqQvP2N
JRFlmTWn6ex8VFO79wiye0VULcVSSPO+vP80VLRtqr20NDhLGJL+65J9wcAxzuyd
TBVonN/DQhZelEo1GnS0nU5WWlyPs46NiRMFEfegi+jUqookYazjXD/OtuYunFBT
HBvOftUl5HNnJ4HGnBg98P46w7+Y207Tj2i13fH8jWYogB3tqwpEj7YxKy5RPyFW
wAyZKaVVpI6MdoEi3sv7G5W/X1Wg97J2BbDydyKtkaS6l5OG8t0FXceWOHBOy9Gb
6hu99OInUoiI0tDzS5zh4TFy2Uzu7aWsIrNLCukFq4GJvjFdIPradDrW/qap2KqC
ZIEcXsAmnv580YFkk8CfQccHay0MyoZh8g85AxNQ2R+BIDkidIwO1bPmbPqXx2x6
saxa0a82Mg2YnFtga85mft1ACOMWzSwCqEcA4E3haJw8WASjo1VwnNB7c7vi/Chk
eL/PPHqYKdDLOKpJsHKz5O9W9TauLY+6yzEF53W03Pe4Jlke4Nv8sQMghqF18Df3
GDmaXzoWF+zCJ6vrlq8InEFb4otfxc7H02p7Yt06RNY5cJqmxLBdcsCMjdOqmCE2
tTUPolzLvqNsD+Z35Vc3EtJZiy6pQV2OXR9Y1AyBhpGJ2AYgb0gRtw2DUVOuKQxh
J+nnm0h1H+cmr3SanhEhe0qNDnJ4TGcxkvSu/1lVtGhERVo8TGr1Wm+Hw6q6LzX0
pyu4Wus6iQ6/cekuDG37+CZrC1vi9MwpvGuCu24JOQut5IOX1OvZYf8PDyFR8x4W
aIMFxm54g/xLLfTUx4eJk1btrMgsqa6NGzxFULfdOupDwshvmHVjbcOGTF3F886K
QQhyToVJp4SPUKztqdhU8RmldzX3+dj5f8PAXMcFIGNww8U/XdIHdE3Sib/XIQlE
YwEwPEhhBInCu+5yWRdwC+dxvjZKUPd43tI2U81DOSD47kiAvAmbvbbAD9NuDzlh
DUR+bshquJorFHCSyyKbvjMuZJallq6vINs6nd2KbePchqL2Y/K7IvBQKQnx7WC5
x0nEX9nxP3Hyp5mtyG3ivmqyL1/brq83YSTZMWuF28owtO27LK7vrre6+3/9g9BY
JHNY7jqobs22Cefmw+7YTjBItS55FVurWFdHL8eNgPnRhyVV31uu7nTOos5tzq4E
KpvK3lw2gcdDY7hjn3wwzf7MKzsDVmwU7HFO2kkV0o5M6QCo1jc5R8SBVVPSryCU
+xnjWS2c6pKr2PW1nbugfQjiXpmjD+szjdw2VmCeDnK61mXfsJPW6OCwPrITY3s9
FOYoXNp7AKBKKplj0KXIh+W8YjvGBMO4vCGH/Shh8wMZjGj+BZ0tEB439vR/M2gj
TflOFlAqkk0wnT6sfOdpacVG+lVTybkjImdJflz41GkKJNeG0nzXNEoKLslYxhZ+
PzelBNclF/UJ0O/0LWjWW2O8Uk3ivSJspVl3Fa0rolny1LmGxlGmmrvQovTGUJaF
5DQtqDrowIWVBw799K+7k14BmYGAq1XYhJwGEovGwPv6tS8EAPlNMESEwkibrbdn
bbjeMMs0DP6iGvh5tENnc+KSE5u3mxq288K2SmBYp62az4i4mKSwos4Qz2/rv2X8
joEog0leR4jj8k6YYq7eWYGr0nbbI8JO3Ply/hYUxdC5eQE7l8Aq4gIbUORwJCcT
TqjoO+4PKLOyttoPWb6R4H9n17Fkj2Ri0Ew56fJXBpw8z75InyvDtJXP0gsmNlmu
CiDVYHSHvzbiInlUbBPe4gPe91LfXlZgPd2VoQq10xUef12A01LKJaSgeGLJAPfP
FkKJel0TRmM6yVUypwaXOjFCxi7+LEs4/kXkEkrYH5GoyQn7b1+Kfvw9NheBpSuq
65fPkt4+1IpV3c9fp1P+su7Vz/4syye7qgXDKkqIir7dC1v+p71GAtbB+ww42MBt
0YqGlGhPawDRzxjDizyhh0rq9tFF9KuD+PmDt7aMyTnNZLK6rLUhNRc5bDRjKvp4
GmEq7XODDdfvAyPc4hreClLNCK5QmMxs85mWu9A3oxMxPIgMH0nEPCkL7bAaIuCo
9sXUjW/VNqH2rve7ykFjZJrXJmJiimfuz7cqCf4aMSwJcxgIqgdznsPNVvy2ib4n
JoXksq8PoVFuE8NWIHqnxlOXslyiL3c0cf3nAvUpl+4DfUKnJn/t4kEVCoJLowQf
RagM5v84CboMVeOPyCUOdh93aDHMJSa7GP2/R7qDZyUQPfqhPPG+o5+5ujm89nIA
oMHoih+AbL/egNTw4eUYu5UwBFENbZpa+CkTlGMfbu0OKui9b5iirFvh3ilsOwJI
mZrfGxMN7B1+TeXRN+J6CqTOmkA276CA8E1XNu103Ms/rWJPLxRChh9ZXJG44RS6
ryIQJnAvH0YM653adOFKNVeehrXzVte+55mbtDesvbalotS2mk8xua5VuyGiOSH7
YjIXqo6YV01SbGyLOoID2ktY+b/VrNm0oPRDYM9zyW2qqyt+8cXx55gAJzb8/jSe
SHaPJSW8385wrTXgNZLVgqjFf1Etk/Xe8SeZ4U+SpEfHlraTTi+6+cUZ5FoHyrJO
c7O3sFpp6+tFs6wIzEMoCticWhvDJwNskRdJYxSm+myOgtnn6zZISTVVkw9/9LqI
fKCVetzcv8FbMWQ2RnmpLcvV94ae07o8L9Q2PFOsWOLqye17YrNYhnmNfjEtQhZA
lzY3qDQmo3bGE+K7xLhQ4PmhOkuxXMK/bn6a0zme9gmWXa/+5AJyQoxDDjJQmSiy
Qt7Oe1FEUhChmQvxrRroGp9tvMEpgL3trd/rXYqjkxoJLCdTxTufb3++5X6sKoRq
XDjdzbbAbxWUTtN0Dg/7diSfhVtt4RIAcJR6mdVdDxnPx60RlaeMCUyjDf3s5q7T
hZsrWcBHdepazHP8++Epdo+18H1eJV4Un1K6Jrfxv3vCsK/9LFeqG3WRWKpPgte8
kkqcW6VQlECKrpXyB9vC6gmrPCUPX7uxc+ygstekS5BtSbyts2zfnVtCSo5sWeok
AintxTm1kV5quMKOml0XcPojDFa2bpiIYhNUzSPYK3OUGeZxzKpCxSHl8p9PXY8e
Snv01AKgmWOFUeBBw3Pkz2DqWNlTVgdv0TgLQQ2/dG6JBWxavz33pTLc+eAHhaFq
HeTpsAW2Lg0crbk8//wEHXjM/LRgqffM0T3cULY09rZCGbQRbeQZcT8wXnsiyh3Y
bprmdcGY3g4lcT1l68OYmFA41GPlF8xKLio9CW2IbumEu1sUFoIqaVY9d+rYauV/
+fx8LxsdP0Nx94Z0iHUx+IoA5TPspE2gVlgGmjf0+nbRSlUova01+//tRa4xAql+
rs/wfjOTRkNkKfsVpL4KnhvP28UP0amJFfn1twVg4cKe9V1jLwyNdL+QY3vyU9/+
PIKDmFh4sROzKkP7uoWwN7hlzrmfiuc4oGiuU2nmac8/pPQsWMp4wkDaCI6vZtOd
ftAaPon2L/o/NMdHtBQlMTVBeBcn+4FPTvsdCLqsFd+AhuBbqn3ZKaK3tT29otxv
+4WrAtkPEl2bjb9OHuB6SYEPA38WvjzrtYVbmyQc/Z9Fb+cQKiSfJhRgdSHh2zsa
A2BygbSVrX4hp94vZK48M+/ViEOf2J294+oda3CymMhTtU3Rw8XfJBGwJxVtVn74
74ohxFx5T2UPj9pSn0RizoGZRmXBABR7xRL+zlS7XqZEAa9Rqz2XsifPOoWvp5F+
GrY3Am4CZ/f4CwHpjDjb5L5YwLtrYXbezItbsvr0kFZT7lOBQCREC61QpoRelwfq
j59H3QXP9RvWuDF0EL3Jxx3IhJn7GpTJ2Hb37j6EgxC+ZR62hjVCJrErKre3VpuM
fowhZRZJVass/jB+9GZCDPE/+gMwO2sxkl4D7ZmeDHuuAs2nIVtXTA9CUvGil1lp
WUjtdcsIfAiD4hoSgd9XuynVYq3l2zsD5htEigEzchJvbvcoCCjQAtVfBW1U44sl
tnAfxnyhohzYuvX8Wzi4KPlfOQ/qBcV7dpyqnats11hF5LBIc4ExttM3L7IsAcXR
VZi3yCKvLoJqVSNPUZpPmeotgL8SJWq8huchRfxEzrZAWSIHnggftxQO9ZLtslsZ
TtcqMyQU3MBiV2spzy3ihxyKRy65aNLaSm2qJ8nY2A3AIhEW1p+wnE8Y1MlJD6Fk
FsF62VBApxFCG54ITj0UO2NZhLQhacRLX2ljdb7PqcuYuf3GyUkzckWgvQtQAT2/
Ew/AWXk+X9meJbxevZ7yL6mA76o2+NatO7pBYV9pUHhP1vuUu9MBLdRoUYdk4nv7
cBWySSy8coJj6Bi1RpgtEOW02vRg0xSeNIvXPGDflBkshbYEpbvCy3mxFvr6RPz/
g+DMpVgQ3nEUqD+xtVfoKqfrCstYiXqZDb+pNHv1nGypLZLPcURP4f/gb0GGfM5l
5YTbwuvorzZCPtPkXJSYSPWr36iKhH9ola0fjuGBwS5HSw4UDXz57VwZeQN9bx67
gWk6Us8gC4boEXq9GI+lIPZZ8NVVMDhTXrsrAkvFHdVWveBqH1L3cjxQOwpsxZuP
VVd3l/5P2ONv20n48KEuTZbGgVTmLWRfA4Ryg0CnzEq73Xl6TTpmUkwMrc0HCXRI
zqEQP48zkgbe0vKGGVMpfpebjiPGynDyc2f79YZlB0n967MDNe68/qdC8uJCfX6W
7es0c8Cz0PtbfKW1cRi5dYsE8qb3pC1NwhBEHjEiEI8YgNchz3hFgmQ/a60Kj6U6
9HAHT3MUykPrW6fEF5X58do3vf+1m4teRZEPHbuOJtONa2uU8XSquAkCSxoTOHj4
G9xjMWI3LsISJVr85TReHrheN4+QdxOU2jP2nieWFVlEfUZ3iRnuFO/6LafEYyzW
hfjou7S02UgTgAug+iHoJB7nM/mcVR+SqHmmJPsMo75+Dh6j/LplqX4kS/PwIKHX
+4WID8sFTDJ6Wm1w4pYTY+zvwHvOzPgQHcZPkUELhir+O72yYPeugPH7AFFGqXgV
ewha7TcU5664oR3fb+es4oJ4UOANqQs+j7BL35Fd/Ww/oypu8uyXpo5CvGHjuiOZ
79phLVKWD2qn0dV+P7HE3vp3o6zzDUYt6RWbCIO/4SbyWieDfmpgWSRvr9ctgPcK
wEnhWjNsKEnc3mHwSX8l6Npejjwh0BOBjmIa8JIuPqDxVwpfKnItsT+SA0wZCvbd
tiOhu9X/oyZM4Vw3VuML8SSrXh6+i07/Cyzl6YucRsGWPGGLxKEi6vuMOXSLEXxT
8AVPb2MkcR5PDJukztpNnDQSg7Kb1AH/wXcQJsLRF2dWQBd/upB4kLj1U1CKQCbV
oAxzHNRGobtvW3uX7sApY2MQlTF96HhRElSWqz+je3I9SFZV5c1VqzyjbBuGVT0T
O0ENg0djW3md/X/AoTMI8Bca6KIkybNL8lQe7sV1ucgN0vVuqJ0Nxo5K88v/zhxj
lN1LfHgM2hArEJjmgARX8v9Drg4f0mN/Wk7BZJ9hffrx5o45AZ+39WJ1D9vZ6npz
47T/vX7S8yDsG9exe2gmds7SHuVMKL1V/sfRGc6zhGZYS6S91cQPCSI6HI9GqhuT
jMIKoVJVOA7f04791V+1TWCBmZeqjhXe4XvsaFC/8repcBcbExBF3LRCTter7e/r
IZBNE2SOGxCjEUqi3AuiLySnTlmDzVezlS/XeEWyhaYAhZ/6hdd594upghSbImFr
XagsuT2zxaTRQWobW9UKlCnJAZu/tBRhC+Lymsrcaez06OnF7FSCZcgYAuPCdYQp
mNao+nPai4Du1GAf/L6zAeQyqM+0K3qHPD12OXMMQALo65vY2XhnHc1wGxIuyqav
Arc4/2RxDejYjMdtg9AjhnoWvgoLLKczLZoULTu9C0VGUgM5t3/VjOFleivJHsfC
vtyrah0ywyMbh9KKbwYDHmzU3mzcQJoC/Acgy2Xbgu3VgWpoXqyZAgzdLu5cSww7
1GJElIIK3IoM2m6CUOYiEyY+eSHPiVwOFiZJQGc7D/nB/N7v2Pa9GFS+HI/iMisJ
6OQvao9o5430JnqOAYri5+86hKJQlSsKQhBlYa2FyXNZiRTaW6I7BNjYynypTRzr
dFofUZqdIZ3nxF+u3UtGqbe0pxd0qv1o0vsMUfzEIkoIh1yOdwXndAfauX3fnb/o
sW6ic/qX/Mp+QjjOMN5Yp5jJOVCD8HIgWQVU/Bsxc3aFLLIn/uJawGEAdwCEQwua
B3n2PhGpWwdE3YD53F5CZv6hNNqvrDNNCELjr74df/TZxBH7+SfqjTuNtxd1xtZ8
RXKqSWMpfcpp7/WVFWxWPz6Yvm2KUK+ZINOOLFhmV5agbinCw79d/1ZAkBtp7vHh
D2Krg14EX2h+s6TCUr0fUsuWUTj0M+RlQBZFiBQf87tmcqIqPp2jAMiT3fLoyTIU
RglKIEt9Y725amyIgzcfP5e7TVETZfou6qlqFb5pebPMq8Ia/0rfjHeN2YV+biUw
ji9t5FhOeIfk2mcIYUdElqvKJS7jSS1uPmXj7UXa0wZa3YjepjNLGK91LE7KtQNF
2hkM30gJWfH1Fn+Cm5kYCv5DCbZwVgF1ESJ9CgIqxId4Yq4fTEptSldCQFWJRp8c
HS3OQ+vGy4jP1BblR9KUU0xjbmFtqx4mlIjbCPm4sTet+pXNBkWhdwv+pfW2/WbC
hLlTSDYQjexTpdfMBtn9cSxf5B8KYAoic4WZ0iZ94tCNEX4n+gJWxMQcV/5PVIPC
eztDVVEFNvpLyv1Vl6im4Z29nyNiiMFnT3RjQtLNovBl/Kg+/Hq2yZbEN4BzPYrT
91xEmR20yHQKuiN8AZqN5k2m21pzWe3mvtc5ox4e6RVhRVVMUqCGrOjmWmRm3aDY
oiqzIyza4u6ChQb1lCnx7ctm6hWK8AucvmenVSR2LgAu+q9Gqiwhh+vHJiV7dLag
1cnbttHFY81xQ2RGpOzRdQfWPbhIVWq1YHpQ4gP2hXOA61Int7lYaScrfwt9h1bL
jKwHfwfn90XBDmcNV5m6gX0C3IJG3Xf0Buw4BbLveDJjTXrHWfQjG/cnIjf3+Uy2
SwFSdfLpGNmW/y+XOtyU3TU8tJwJxIOOMtKAVPgVdNc9UQiWz08V7xksVytUEDQ/
kkCKTLhzz9Ibeh2RvT3fpUgjudHyQhZxEezV2Z4AHasby0KDc/35bzsJSD06CetE
aUgy5Hg/M8ytXayqLA+Chzpchd0TP5kyp9OQkPbYXLH0oKXPDqRVSdTLrIJHJaTK
ZjSRTErRnbtVSZZu6Se6WFZNNu+MQh/wViisXOIEg0v1l+izeLWzFEeJuoVPRuPD
hJODZzSZYnf8WjAGsxYJfZlS7VYFO/67rX1JxjgyTl0ibUffvant282yYq1YFbWF
FoObIxzFkoeKNCeYzv8t0gMSeMHsm9Q2/BjexudtXY7Ab4Q2YHQQztDOnDBHMw4M
84OdzxXVHwiVZasAdI7CyuGvuUqEgM6vpTxmUVGOaXZDJXzhFxav8Bw2s+x2hOAh
OzWUD7oiEh5aaSF2/e4qPeIfGw6YPnlxmF9h0sTZn+j/umpD1zlYE7cHI4gQx/xw
5PWhoJxcXEtZzlEUGtGiZ3zqo29JLxiO9C22Suuc5IHjXZwnHBZeuU7HYfiqiL/S
OP0pHqQvr/ITx9/18lcuGobXKtPfBu8hLFsUyEmXNu7O7BSJstcifoBZnpqmsxxa
EiZNf8+f7bydmk5VrfP/A2iV3DkJWq8BYf+jmuSWvtKIbwM+hjpT6IXq3050qC+n
BS9sIOZUbnDHgDeuaTYsIOpvfETjKEQn+WyZ3DtpWWOlQJEkrPKl7Ht60r5FRbJR
b4wUxjItFwlk8tO0CXIedWvxNuxC2+sk/JO+Z3yYmZLnDU8AP3BilpDIR3v+BWOd
PHfWdGfI2oEh+2NzolPSF5WrLdu+wqQaAf6s6bnhHb8p7HA53alxXH3fPfBO5VxX
AO6Vt5d7UIf/2IJQpinJHpaVQmGmfT3SYGOfMBxxY+1+mbwi8WrjY9mpNyCk3hot
EqlpF8BAnKi4us/dE58rTbERPbHBj7ujzANYRFky8LxjXH9o9D5BnVZtntYQSpcT
ioHPYxfzEOxwbAjUnorsxRhfmXm3mGIVXneScFjgbw8vaj+h2kAOz5zjzHMAHWDB
ZpKoInRN4kVOLCvPPJxAXXUR2gMr493xF99Btbq7dNwcT47+BdTPCJvLoMyCzyPk
mUyn44UXf1K3yFAu0uIAUDZb94yuwmpEylfbNfBkhiprwDLetxx0bTUhqk5tBVlA
ml38hE5IjmiQPBm1YcPtZIJUyyqYO2EFg+MZfZg9liFixBckWOGVDl0i5JtBR99h
I/HTW4v07MjYnJt+8XIRuT+Cd6zMxdoUy9Lvqx+gNxIJadmbvmloykxG5LDe3hDB
OGDbehQfVhi0nFkmihG3yuXnJaJVW6faWWfRpoXMuHA1WPBv+d6BXTO9dQOLkgxQ
TA6BiPEYEeh5RkRZO9RHwYedaDSE/Jx2J0e42ukOcad7N7fWXkj+lv649GD+VgSn
XgIAeorsOfPv9jWpXJF+5Lp1Jz/q9Wp19SmZRqO550E0XgphMPGuB5bXXgLzB0d/
WuRIUlgy4HznddAbfTCILWMnmL0TOLYY7Xc9MUC1bJ9m7OSSPBJMUFGDxUP5dnbQ
rMJd9I3Hyf1hYqU6PLowJBVMB3wVW70yq4wbLvKhdoEXKA52ztyPQ5awuAWpypXC
PKje4Lw0AxGqi3QadykUlumhm7efBQrhbPuGRNpnpy+dTTkpygl6VK40Ve9l0EE0
eDyWzmBZM/36OT50nr8HimwujcVRTxaus3C78NQ/vPDDJ+ZAigfyzGQWBSZzLQzk
cUuHOTMW5bUAftTl7kNBIvOdKqn0ZhTTKKSMvoCNYI4v+em5D5nPSOw+++0I3Acr
s35AAKqHDYKL/yOdThyIz7+gBM70xZroY0jtcDQKBcfPplfLtH1NTS4KOi/qPtzp
Rld1p4sgtZJafXtOGEYThgdYESbSK1VccZVFYHigiOiDeVzCJfM97FpsdQF4Y5Zz
ZT46fG2N7z67gKnU9yzx2x5ZifbUUuOowIJCgjLS2aFHx1Et5ldYeo0fmnUa2WWK
59P82KsQ7LE6GjftyU8sP6XaN0qdPIuYrKFfbTXp9nnVqFHuYWTgGSo2ed82cfZi
DTMQRY6BOar0MmDHMui5dWAh4TdPCemZ4jp4Fk+0y8DSTZJExQ+KD5eSvFMNj1wB
Lw0eTmX7x+OrEl4SBzezyhgTGZzRl5kGh65hRwAiTl5/DWIA/ySdqmTr7EejzesJ
ONbt4E1B5mZVSOhJlcU0fIcJoM0WvE+tFxP3BCql+5R+npehtJbDZoP2RTLfLfuW
U0qY1p+Z6sNVZ8//I7SJY17uL8lNx5YPgcJvbq2G1Qx50eIUHawUSpUeAE9MtXyc
ZHh+ZyAMfF4T1clZfU5HD9qVMgPpTUVXMUFZ3H4P9hqhgrw0aiH1v36C0DyJAtPl
H0ujGd2Q4B1y+m909ioQec4kx9KaPD3xPPgr8hO0cUHA+T3rvgyB0DA84Pi/kg6K
icNN7EYUfExXLNRiJiz9YJSLNHz1YmcTUZCew7TffUNRydVHESzbVa+rtCgXT+UQ
BQ/fiXk91iJcvQfw3VxdiPLZikhxvhanToNCPnwsuy+lPAeKdgNy45dln0o2J7pp
1h4ZSbtj52UB5CQT5nyyHY/r2GuqJ+y3/1o2VzCpw8HsqK8jwmoghM3F0QJAOfe5
Sk/udjExn5X54DjlcAdrKJI5plTitbCVKyo5Yk1fKgGoqInN74gnKi65mOb+yLBC
6qrd6ts/JqKe4tQEx3osE+gZnUmqgE7BfP1Ncy7F92j/K/lZPuYPUAxmdhpQebVn
5+gxzr2DYj66VQ7ppGZGVL+bDJiSZmpx3Vq5y9WAQpQSv55zDlcUhJqO/NjyqdpZ
XW2idU4ii9iA9LIuSx6bCQjB2Wluey7ZGpZJw3UAZH85hbLlea3ZzwOTcw7NDK9j
w+JohDJ5xEXgQIxB47+h2jmEnGCpp+7c7ivfE5TnSNfnJkNws4jjxWkFOLKf+h10
LRMBBXBt3AGc03ouBrJE8nC0B95DEV7IqJTFvLbH5mEWGoqoF8dfALSHzi+YbNfc
gEJORB2MDuhipKnFwKpWnQMhAnuP/SXED+dUYajw4w4Yfmo7rqD0Ap2rqyp5Q9i0
RZeIAynZxEqXWZeR1Ilf4x+OWqJBr5p84e6ugxptZbbOqROqj/8Hit0V6fvNXTru
PId+hPHBeb7qslXfGeviWz76z2Mj5iyf3bnzUt6sh+PIxl3IwW8CgItlnheBqL2/
RTI9rSJzWCbs5egJ9oQsn8jTra/oUUryd8BFcsSgoiKsNyYA5FkxR9MFnXuIVkVo
Rl7R+n5GrOvDHpW1Erfrv+/6wqZ1YxpdAQv2VCjfV9sTOJxxh+OF+zedJzU7U9lm
aGeYIAeY7UNcCFYDYqGnUw7RvSi39fEKtrDa1EVkMSwDjNUrJvvDi8yGXNFDH/Qw
veHA9+ryCb9FXEBMyjOSPovLqL90WcTa0r/L9xH4P+HepNpx40FX/A5qbz9Um0bp
oy2q784OSI9XunSWOr3UYazCGg0Hqs5PlsKeALJfZp3MkIrAQFJBABx7ek7HUkqA
MXYL7v/WOTWInjfmCAbZzzc+uuT0x1drgQ5iwQKfnSGxrt7g2oJxPCOa0ENIrYhT
U06b+9YrwYbxp4IQ3mgQwvDwAiE6YVLILbOkvPcwH68b7h6FfrJl4wjxepAmWE/O
YR1Bj5OkojaqaGpMxsgOHJOu/mc2HAfKzLUfspwJBJwwExIGBJq3u0cUfKUyPbQQ
vxefPbRWrGfjMFMtNGBLEDvT6W4HKs3cbT0WqIiwdLRGfixDkwUs990pkzVbjlez
FlfsTtKlzidvU1OUYit5wHV04P9C2qrBsvRaum945OHBQ82g+5JJ2c7HBWPkTe/W
lvweyFEdHEgu2Dg3dgw4TcSf8lQpsUh74n+1VPG9FMW9gwmUHY0mBL9WcgovTyk2
RJQlLSGTsTv8ugIYNEv02Uhe2hPIiXuJSd+dS6LWxME=

`pragma protect end_protected
