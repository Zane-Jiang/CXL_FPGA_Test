// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZIivsP6phbg4sE7veRawa11aBV16hM6wzJrzVhGds2qPVn6H4iZsw06nPeET
Un1TdOcDFCD3xOuWuxwbC5ZJMfxPiK3pZ43shB8mbJtVdn7WMyINus5ZhaZC
bLNFkuj0UmVganr17QfVGcKejyDKBn1/WH+Ys3jfdu09oaP9GIb3E7WHw7dT
SGYpZwVz1NDOi9aPruE7VSqp9oU3phxEEKoUPQIVwMZpbZlWpkc6UGiEg42b
pF0VOfdVYfkSpKozkfgWKwhgDwc2YodGQ6CoOg7o6gFXv07cZTNbfZdUDLSh
MssHOT8jjAQZhdoeKSR03HwudYuxe95eYTu32JNYDg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SRh5MmYJqPkkw26Y0HVyCiqxGbz0c2h5iQGJVx40zkk9CVexQsF8+m6yn2fN
Dw/iu4pnvAXV1GF/cIx4Vm+tvljGYjJ46zcxLfDa4rlcJo/H1jBVb5kumagX
RKFyf8TCiPE1HURsbLgyQq7YgUpTz/nIV4WkqprOI7sUhTbh6hfHo8R45TGs
G/VWMxxebELmJUjzXoYtGlZSN71X6jSp0LzW6hJ88p/WWdLCF1H36+AhQL8s
8URtwwhc6Vd4e7NGtWPX66fcj+rHFCrc87v3n73MoO7PieIOuhVSZHH21x+o
9an3mOZh6OI5WviWp4u5dyTsEB4lScW+Ds7Rf/SzmA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OoGPGIzXZtg4Lyhk83FCFvD7XHHPWja0fx0B+iBMCeuzz2rahmTGtGvHxRAQ
1YXdathPRCvMv95JOQWkE7nwZfP35k9Abm9D335RM1Iz5UR8m0JOstjxAD2n
KzHeJB7uVYIpFvRjiyy1baCiBKr1cb77j/b5OOe0wIYXEu4+4ZcNQ2I1Wamt
lSg0gTSqoUUPFKk7y9RFBh7FzEmL8FK28ROAPRvHf007eeaOBFwSYd0YP2hZ
FECbbdMf2SvMb9Khm0YGGqwSy4kwCiNvJGfl6S7IVVchBB89S1+0xEbqVdVa
UKVVlF1P1AoPN4DpETXmhWKyyfQAbcf+SmDPwb46kA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hErtGNMGzy/ssc28fVPQg6LViI43U6Ct1+qBoOL4ReoF6cZlJCcVkVcIlFe6
UlN5M9VoXJ398qg6BoIDjq9/0wTyCvnCXhxl0HgRvPo6CgoVbp40dnu+4mO3
KokBFbnpHTR59b8zwTll9tAUaoVcL1NSNUvHeAAuYA2Am20C1jA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jjL2m9iiZMwodCLa7Wg+zMwDZQv6xw3DCL/ZyepaMyIZY3RZcvDtvv/NB/K9
2j22g9yY6iQWl1JQi50xc8zZNFdsvw1al1tQ0dWAYnj4InDTMdGooxNV9bSO
Rn9xkl8IozHz20H9IUHmFliwf9jEe8gJK/6quG1SPLGW6B4yNi/QxjrTs053
mfcxkvUuSHUD+nIH+0FUweiesvm2vBQmn7JXxNWwUz1e3ZQrFxv+ARBkFDiL
sLKuOVc/XzNZNaIP4ZG3fNM2UtFisrdU78R2GJiFD9BSx0GpwzeHUOX8LUMN
dAbYsfAv66WSUvt8gMwdd5z/JyX8mb/j1eALMvm7QkDevciQ0j14xg4Ho9lY
HrH/rGfelQn0qpq2wmPoPhJGu57GDsUIX+oh8OANzmk3Yw16Kg4Gnt7hOO8P
cOEF45TyOs0sWAvr/MowkKldIZ7YzM2Wvc5N/NtGWWbdvyoy2XU0zzH/9u7m
blV631/PeuIXLRP2XXLhH1qbINNnpK8p


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Oh0QWofGTzTop92kVWN+cGp1eX715pS/+tDvlzgWIZeiEI9UXQjJc74i81cM
fWqlwdT0SVftXFY/E3uROuEggIlMS+Z73i0VXb4JjdNmtdDVzz7757BiQdNk
kkViso/inn1j3T8DYFSSJxQB8xHMi7mjGb/ii0F2Ugsvv5PiqB0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jkG72fW1DrB/vSJO8AJ5jKOmXNlwD3o6OywQb58s92gis52v4BiT78ZSkyC0
kHAxIwM4aXUXv60J97McVkDgInsGdF6NVvO4zyAA89qARUTkmT1vMyoKAN0k
Akw1zaeyKQxRon3RNxSMtzosDviKlshzqxOsWlst+fUPcgHnxiI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 22880)
`pragma protect data_block
dXv4RMXaK3K425nSQNPApXdO4W0CHUuB59CQlTxIW1rd557qrDX/6mZfSUTy
F4ckt+Ic2qJTBuG4GIdHy3wpBZFNXNPFmjuMricMxxZgkx8Ka6UGXfu/jt5t
dtu4NSfdb+gCJjd005EvDHmNUyLtcWOW7mmXyf8vSX25NdRQWYDIvEOzsyHA
wOHgM1fYQ64P4sfH9TBvlulIX5Vh3w7/24kkvmD0IS/xlaXRxc8/+7mF3hZf
v7gOUehBtNp9mqHyuih5PkfewhjPY6V1ajJJ39ARkUF+sfLHsYdjhf6fKhmH
C8t6WLRjutcTtm+POn2hLnasmBRGtkuhO9bRDov+locvKYUGn2c9V9XZrLL9
KALixc2vzYRslxQVjpBLyzkNPJ1FYr1EbtEBEqY44dVwPN5vSgylYxsdNaFu
evOlyJ3/CXgJdW6u6+gW7Mjdgt1vtSmlSftYgYIKqDUR/5bChWwG96Op5pdc
Hbn80SrMv08xOsJ7vnIKzRv6CHqnJgmRlv7nu1bUPhWGLdq1OQJFA2TTf2iF
c7md4Bx5LLV0CmXhzWrWHWzpXdQaZ8fOJ1ECHw+eYUDZqRJmC67v9QZkwpps
l+lF35bRLb7tOKiTl6yLI8XCQKNPlK5+WL9meFzS5Jdslqf27fXyC43/VmjA
F2NVpUINi/7gNEiNuGsNsAMzv6jBbP8MuwyjgM6ylsis+f73ZR7lFLJzAP0W
hcoAopu5wKqY+dZFdKfFqAMYoaRu18GGgYlUzUK1zsZjwfhqnRHhD2qMc1Mk
QmQxfafH+SRYRKWpDy0Y6/rMxmeeagHnGab7iVgTlUWGCZfu4CnySVCYQAei
764OCuySOHQ1jCEMUYbiXegD/J09HWI2CbKBcOkoB8vbinu/+n/inu7nGqUW
yUADKcd9PnMLuE29aDgzYdmAoBL10tCq4na/VSKrYJQA3/hPfJGKDJwQp8w9
G5BXQY5vnjSBZ6b5Lq+oM35oEQlGvD8ZMo9qQfBzTUPw6DYoJV+HVU1piT7J
UuI0hRPK6zuQ8RFeN4pC6nCzAdOPM1dqPivKQyiae83g7Pu1ZaBup/2QITt2
djM6fhVemi0em/ZbpgjO62qYabBMJyP5ObVuKmJNLUGNJBDhMIjOLQJaJCXs
VX8sdYDaQKBqSrFkxW8jLk0Kw3L4YDqORK3uzYAJmMrD2jsf68V2QMAs/kqs
luq5WHYLTUb6debdnE1NEYggWgbr9KxNUF08ec4rW46TWABz1sw/sqSZEpTw
rQPpTw6LpTBGo8mELkKyxzAGTzK5es2/gmMweF+dZHL5rQqTlp4sFqnxppdD
zAdK1Gm5+CbQhCjz/2LbiUKoUo6dYAjmcV2dRepiMBN7f0wdz54Y8hWVy3qC
76jYuIj0tzEXiIKSUm9sdzbd7t7h80EmP4BMlGSMSd/cC6LAMhXPDV5wQqoG
l0V16SZGVfjod3ADkIwwV+MPleBT9pg1eXesHhv2uoXo/S19YyZn+5AHrRyt
JM6rY6RVURmpTjOac90sNu+hSxlj78piU+ErIQ+rkZZ1VIF9IBVO7dSTNULh
ErYjrFKc0fNFEBJztf55dHpgCFTSYJmzoVciqQoEjwX/K5/9lW1tc+8DlEFV
Tzq2lhpDoJ1NdQkCfCqSkFdv2cc+px1fBImsHfh56ZZYPtH+SWkLknBb4Ke5
BSJw8SpjrVkSHgN4ZjLhyT+MK0h6qDOuxwWgPkhiwygwe2s6gRJweXo+ca6l
Qf6QKHHG3SdmHXpg+iGMkze8GEe5kPmywdNCjju718JG25ORdwTfa+nzdAjp
NYkVsc8B1IGBL7mNB0aB8/i1NIXhNt7VdpSHmoTBqwBvP6+xZLYAH3O6+PLy
lFbKl2d1lqHppScHxOZZI0rCRDAIXMBH8VUo2ZtOJMw72uk6jN5B48LcsBx+
I7bNY4u1PR9E7A3ZP9rLbfKE1cgnjuMRSF+SwAeNBRRZqvSLj2oyRkYgv82L
S04I3Ks5kkvsqmecvI9SjutCblVyUj71q2GVBJiHJhaZxyvsHStZgKjNO2sI
xV/uJhxTd6W2HkLiWm/+X6LWzJ6x/hetJAegPowU60ImUL8mWLOFr+qxtIPH
BmCO2RFwNcarByrWAjYV3r4g4yeC0e8FQl1qPRtpFvHsv48Wl8QbZA1EeEPs
6WwdP1InQlXVZSJUTzuYDXoa+g1rc8E2NeF1Uq8T4nT5R98ltX3+q5Er5o4q
pEnn2gN9sg8wSYDvh2Mxu5e43ou9ilth2TKmiKzRqNGITk30qFAP3HUcbqYA
2qlGNE09Ig4bow+sI8Ig88Wp44avcpcrEj5UY965N1mYOXU2wVTXee6UEJB9
AlrJZqmJHXPm0DBaaAbHBeOoyKFNSSXC72cB6IKdrGC7479NFK0lctINv2sr
3SE+SVmczakLpLiol++o4gRVC3nxHxbZMiXJqzqSQI2BDMuzwb4Vx7BpRUtz
47jfGhdMZWjrwsQW+xg01fUYAvFe69OFmYVK15k257Hh3T+T5G+O26G+is2Q
CmP1cE8o0NZa1rdX2sdY3Mlpo68v0w9oETxVnKfrJgbyfY6MBs2JwfaTpGaa
+2/VuGQ2ujo4n0ZdePmvnGgAAPXAkkY7dSBHK88be51p5IKEIILan3VvXFAI
aVKWQMZ9Gz9Tf8/BOL3ArfEffnuwiYMsXH5FVh4QTYDbZ9Nxqa5IuZAtKhk7
ULJd/6kePYwedWDl73hK/m2MIkvkHu5g5PAw832oX+YqtovCjV8jGw0Bmecw
SpGU/S70CpqUIhknSnOPMMwi8qEy0Mv68wpPtHpAmG1NH88B9ww1jx3vEfF0
W2nGi7H1cnQ3yvucF9rK0zAE9eNAQcEn/BBAbZtRb4VfHEQoFf/HBVhpHorT
eXsZI2OLFn2PeQLMnj2iw7mM5//GSnpdE8Z5S2NJjEon4no0pyTq6v30CaRC
maXoOv7UU/hwPbq5E4wsw5i/HmXaxZyJwiGBmNwdUz+5kYnKlV9oYY7U2uSV
64ss7Foy7ShNi4YHGtxyYbk9Rc3gpNkDj+cjvi2bP/uRzsAkW2BVlmFkc73g
xiCruyTqr7hBVBUslnlGb1nbNx55zTSkUvAwOneGXf+miHb6fR4Tb0wTNlln
WllVEne6NfLb0DtuVL2Y2e5XnEjjIjhAiZh7RvU/A4fIdQpp2+lNc93JHG4s
FEFGA7U3FsrqLTBvPdDn2xX+Z2+Ejs3NYCZofoqcsH/DMGW+l8XeydWhtnc3
x52bIKpsTpvM6dVUZ4WsTTBpGjbA/WzhCuY7DLVdICjoBCY5hvgsXC12yoMf
GQo9jr7bqdormJbTw7WFhCD5FBt9U/FXRn/f9g/vvgAZoB0ZlxfxdyTYEjvZ
b73T4i27Y01By8AmabjqHDMI1ZYdhKw6iSL6QRTurWzoWHlO3c97+bzYw1mc
Yri3JV8Es4/kBX3R/yRcYsg/y47bLTMljjr05+yTo8MuAR7FKl0XLhi3YYGc
VIPj06JcF+4zioGRBvy89anQKgsY3Yrv3ROlLp5vih3HZ9pLPW39P9t5vGbe
2bGklM8tHF7kswNUUtJdRzk0yofE03xvU60iLsefuiTexiBY9voIZ5XlcQEz
zLSwZTsF8FnmcDsydX8Exy74tUxJs1PQq+8ya7P0cGM+ZbEy7UN5LqEsGznw
Vjybv9hpdDJFH5jfMLjPRwI7gS2WEWZq9nXWPuu+2IBF7ctD4ds5v0XGo56L
My5SQKEZbxfNzBlk2jjLLu4u2CVVml3GBWaDw8JfGxX8QMNoxNsSN3mz1L/W
Alz/tbHjCCNFb+Ua2Dk/ccuuryQoLZZSMifd5YQGwZ7m9UdHUXkOQf2W/d2z
BgwZEKhubAtOo8eqj3PwQfGxzAmzu6DPk7qEM7XwxLrkSKT0yBhlgRW3WFnj
Nx7gew2P0545A5d5mHnoUmbhJ2oIrrOsIGGHtP0+GT6sw6wS8qFwiKEPau9O
1gYXZW8YV5WNUSAeRKSn1UHYWoY4vk25Iy0l8gpePHYWrNXHjXniEZdK5ocj
zN9rPocwBTkjxGS3BAKYozZ8pNmwX981hTU9YqHKCrVXk1uCJZNd/qxVgXNe
hGVMpB4SkSh3CtoESpQWvtPf9osCQKaXNywV/BEdd27BMEBamzOAxfIIOo6W
nHDeKaQLsQgqWLEFkLit9CooPdKN8ylaskO5VVpS6gYIiBevtRbzEEO/bVch
ZpFU2p6YrHKKjXVTQY20KWL7cOyYDTiTAe1QIZ31hmS26EXZOIDSMqhxt03f
atUPoO/ZNfeXswYOYxPL8zJdnLLBt8uKvK1oo4nLKmT+CTUW+fEZMFjoPB1k
sfuUs9CUdm/gz1xNJSxowruAJHQx4FvEHbvIoopi47Fr1qX9x3/h+rteGLOO
UR/dj7FD5N7+qwe4icT/1amqFry4x6MZsfaCQyr/601GXSmGsEfESVxV7fW6
YNyC+1SQKWTHSa53pj1zrCvlWkXEWp0ROvHaPx/oerc4GNN2WoiVbA+kotFC
8PN84czzZLAJasU9NBJdeY//Tmz1RBAkj4YM3Dpbo+e2dQwA/1QnueIcdFwE
K0fimbe3If6ydOWMwnORcKCmeRDJATzJKkwf795p0ncp5dxN93900ru3dNRW
L7G0miyuN8kb9VrEUoQeUqwfQoVdS9y9iJmeQYJkoMhl/QTQ6JF3EXlLQFum
iSmw3ZpcsTA0Kju3oPVqQpCKX4Bep5E6+VBv+CSoO+kFMsVRGr9pCUWlI6FB
n+JvoKibYXQndf/MDdR2GcC7MDn+QAhFBTAgo63pveIRZI6VzP+IOPxOaqZ9
JYMBJU5RxMvTkJEj+XoKRRL4v3PpLqgSL6XJudH5CC2v9TxcIHFg8yyJH2sd
2znuMBM8I34dWsLJXOEfCPVZrIY3n7vVVL5buzreHh+Tr2JCYHtmzvB6qj83
+bnpSv5DKJ+AsnjEI9nABh2cYW2fX6MRWdFKnkLsM+cy7NMpDMPTeWff4gN8
2ltpS57G6hzEWYX3T2sR2kwBLKpOtAeEepmyP2qaZDJe47HDUEmI909oFbug
zVxNkfQcDbH4A6nH+p9zpVphhSWoSUJE+L7InaIfID0uKcZXdOQ/PTcy10qK
3UdrYvXZaIvDiulj8iBcD9jxHo7NI+cnGUscAi53ESfuQZPeeZVHHomTWSZR
ITxWXUebTzeCa9CRdv2rmXWRyIPPSkoPkdrXCygGXbUnn2jrY+43r33O/uDC
k2xfIgXjvFE1rhyGqcw3HiiBzkDvJYTxK+YHl3JozKdGPOoDpZF4utjfztD/
l4KN6bjE/IAGccLXbntxTImfHYyC9QLBunhEyAmLMUuPZbshSZTLu4als4dV
haNr5pEWtmtRiiW7r8LCxQYwPH26Xp/XUeUkmN1KgtlWKy6aevms9bIxVYqF
Io9tbxlGGGF3RtenGHsdXywaQxlgyQcDBur+oLPyol875oKVAYRkYLSI7vtJ
iBCyD0RP0SGdRhkPrDyQl8uBeX+oOB4lJ2PMG8tfA65TqwLGJXos0mEdsAI+
NZzt9/zmqbv3Ds8A/pBlTnm4fqn7Ub22KqjqnfgRBjkjJP/oDuguSCTwzQfz
n8idmAwNhZu8+TmIbo7BSRgevzUQgVD8Ay22XBs5k84hCM6xT/oNorlrjT0D
F2jvnQz4w0FyP6NzPiTVHbu7eBHM7s91ePvCrlfn3QH47AMfTk3ScCf9RsZA
cjz/esKNa3ngJsgXHBnfVv31pWuptgvkt9uBGs0mn1/OXqX5O68CPne2wOkv
1KvaZ6Uad/DWL2UaFVzJwHITcIwFoijuqC22f9SJRqHmSHJUeFj+dSrBYKm4
FFYESwhzwCpm/R5Ukv/ALd2U1kbyP4MBNUv2XYxMP9AhrvoGZANUPRGthcRX
HjO/TwYAZz2iFIBr7q6PHI7qKWcCO5I+0/Hr7+Qqa1BogA60JT0l1FeIeRyS
caYA6/+3MxussDZmgMIE8jNb4qLCyc28UqqYtX4mlFbyxpgxLrynp87yu5Jo
VilsZLTSbnspVssNxklrcrG57SvNdV2uC/vvYlRSv5WSQ8zTCZt7Rcoo2a6T
JHF6vmMPsXn0VmutNtOR4Wg+csqXX3E94P3AsXt3yd4HVKfxs3UfKkvqvrux
c1qtKcIJKlZbRaSyR+EuB0z68q9PmFdC1XPA1QsHayxQzRauNqklxVV8NMVa
29U//kJZ3LSfpUf6TCD4POduswQf+tFm1GOoZvt9ZqKtkzbj2bmN5I6y19kJ
PPnKKXxSsrgmM4G6HnRD//BfyCYcsd6KlMjr+znNrXYogaSdva866AdpxQJB
+YVsz+vH3ORYa54hVgtjV5EC0paLMsqYsl0P46EFNAzcw/taenAYKQxQTe1V
1GXZYCpEx+Izgf4RnaxT8AGRIt5tHgjQSD1oyNL7lu1RvRg4GtdtaUGGYJ1j
L1hWkHKuPxK/OEKU4Y9xKyulNFGJwGAIUQ12vT+YRC/9r+DZh6THjQmvQeyS
NP8TZBxHBe2UIIL5zrmNHFqIbRi5ry/rBb5HQHTTib6d2BM3/QT+65N3S/vs
g2g9sXyJWnKQOMeY7y3gJ2uF8p9lKdqefJrTgPsyP2WfudRY+MkNEZw/l0vL
VLA4QPrhPGy7Uoy/AXfYW0FBDs4ZXAaIvAgGdoP7YuLOoV22aO6H47I+wHtm
YUY2b0ToU6EkuDqJOnjNalnQQeHtZh4quxVvg/Vh7OBBlUkoLEMxdaKLVDeG
5KbCEv3zfamYn2jmtXe4baEPMv2L0y2l2ZcXPMhCKWAa9B/mwgyDAUf3NC4o
yGBti2vZtbPB1MmJp2hCDYz1ZWH5GVG5AFTBmRyo67zYHoD89DRwtdXQXwQm
X/9tZL+FjjOzcwF+9nvwTKEWTp/8K8p1ocb1jQR1ncWnpidfbFvMuHCu5cZ3
VYK4M8zwBQ55iJ/QW1cPerNspycx2wM0RyV+7OO/et4YMffyqPTsSv+A9IXQ
b9tZiCD1KhM1zmi6i3Sl1IvezNIVoq0CpKU7JUtzVQZ4aVPYLXX18SL6LT0t
RUG02V7UboWDWG54waMkFlIg6O1F7SDVegGaxhH7rIz+n5ndveUHsBUjKa3o
pjXRrekqKP9iwe9EZAlWB/wgtpdFDCjuPODX/HCmSIIL5dqgTaa8VRFHCl5o
3Rq4gAj8DEsDqu3ygF8iwN9lMAk0ewfXradTFWadTh45gmk2lIuve4wbXAK9
jUaGWL4gtLnSB3/XrRezhaZgqWoGBo/5yqM0mEXO56D3Y1K84zfCxnTIqkUe
2ch13Xx5k5cVN5eVlF5nC8wtFoaGAttsNiF4PRFnmSfAxCKe0+IFSoLqWn+1
KiIEkryhf6zsHa6k6e7xUOsQtRM1mY+RgX+qrvvqiIobgxXoHgjTYgJDpI56
fiC99iugtg9w7x5hKABVXWetdId18QNqhGHgAoziiHGL+glmsOUQsRYALPw5
XbB90ivVQyxCGA5IhLQLyxov/yAt8teXMITqpSfI9yKO+qsWdQam11pGJfJc
pafTqho3VibwuH4flMSvuY3wiEZ27Yr08/ZEbxzBpFRlxJuBpFxFg8HjAuf5
60DbSVX3G0L4R4hC67q73LAxFJRRSr9oNLE0lpdIKsXp74d0pmi0oDp/yY96
6avkN026h+m3O+TiZJnGenDhu/9qWebWqm8ATo+C42lbjTSIZ51t1TG2gbz4
/kd8Hfx0ekr/4jgs80I3yFlvHdxd3rrQ5q1g/eW4Zhn1HXgamJEGtrYxXN8w
kJxgoOA0RNU7Fo12BRo6cCQ/JnKHRCL/yp7UV6Y23vXKCwIqLej+xhjMlvUD
bTbjlcP2I+UJ+JhhOK5qnXH8wGu3wrXXSivgQNMHsCLEZHrd8/8OfBZEPb7Y
CSuq3oxGcrTgykY4QPDd6ceoczgvk7I9V1LmQsXauvAQJ/D1NdXdlJGANt9i
wLHUmLs26DwqtgACGogb2547b2bZZilK1C49m1ywLga8L6PjjsHVl+hxoJRi
+zCDU5+wr/80VWrBSo9Ad/4OoZuvnnJDsmZv2IJx85pDHbTSCIQBsYbsMD5D
CABL3xwxCjgcU6GJJH4kBcDbGlw1N611b0GJeduR4OTXREG42uu2ZSZW10XR
SSCD51kmQMqh5bEz+RjR5L/m4RHcOk91TE3mwBYTzsAdt+A6WlFWFEWIyoVo
ATDfrS/ZcCiiZxMk1O3dZrZ0CXpF/cmiwrvb1nhS4DjXd1hWYZKWoRnaqvnI
33Tl2a2XjntqigOo10QIXC3GzDvsh8JYlH89CzTVa9GZC8dWUQ26pELfAJcr
ce0eH/lNdEg91YH5uIABbLng0MortfEiJx/mYzTgW6CY3VMAjwRaLyEtLHcM
YqMrqGb7hcMSgTgGnD2Hxb3h2QecGm/E1I6kSH54olZj2qvw5CGOPrQ8gARR
/ut9uvlJngG6Hz88u8qoTCigGev8GvwC1S2d1en5G22VNoDuaoBVaMZtURY8
pvLsyIuBbxI2x4qG6sd2nH9N/GkTaapTHWxBX6RcD1z2JMnN/H3ggEWJiEbF
kOlYXuctyYDGlYy29AWD2mmhRdF8gueAQdj7RtpCyz8EsYLbaLCiEAvvjm9/
9uMoPGuvAvB+Vcc+/v8ouqDRa8YBnjFPd0uUKYz+uZyEybGHSIDTBRvLc/6u
bCLk2mWPSLOz9Fjvul4mNU+HICOtgKFWBwDp5jInWEqBcpXYfGH8ZHrpJqgY
ZGUibJSpuqGg8Dpr1+PEla3TPMpfzmTv9nqJ1GuIqHW+nPA+JQT6HYEfXj6f
66cv3YzGGRN9QJ9AvtkWpiOxtJ5LzEaI0OYuzZp3yFSPHHuVH1nWNctXoAyQ
9pE912jVJVpjKusSvv8sxOBAl4V0Fcqzv9QgO2dCsH+jf+YkOkROjWsOtoyG
QiTy+ofvmiZxpdOhfkadDXcaZKMmZqWRAfbi3KCqgTx635Pmpj+0ZefxXA3W
hngSkKwHKjOyHfAfGLY/Y2DZUfQ5mglRpHTN30WxIyd42Bz/Luh7V5DNJK2p
QGOKWmTcXTN8y+LuGVieaaYfAVBtUoA180JvUb5iDUpMEhbayh8Zc2EFXTuO
PmHMR242aE/pBmATAsMYo+jWJM5JRpimo0Ier8AKg2WI8LBkYdbIkDhlr247
DAaNMkk5InIW7ZzoyBhSSA0XgvCA5G+bVDdkpkgdJCuVvaTJSewgZyk7jM1G
A/cjRN4PHx37df/JW1r8KvBAE6vrqcVAILPvQht2kp4rMMoUVQla224vxMEO
u+cLJtvoOnaW6wPZ2xEM8f2a9Im/cD2MUhnrQylXyEf6PhFtjIsVCNuMFydf
6/1rvLWMH5CSeC+GHMw66gk6AZYmFEd1G0qYarAqW7FymkmzjzXYs6tcbMWj
FLwR8HG2jE6dGLzqIgTJhH00jyoDsFQstGn8TFaq8OEzzknIqNgnbvizp6pb
tqNneI1Sm1X2dIIzcNzFwcjIKkbOaqL7cVXTXOf+i6/Uf0C3UpNhLzOP9eb3
+X3AUIGbUIDg6PwA1ri/w/zSMxyFoKOvf3WVJD+AdLpbs1lTyG9z5l7Yp3lV
uSmfv3pk8FiIt8cQSMnebQ2Q8YMG5nN/zgOJX5NbRoOaml9jj9UXUxsRFI33
KyFt/Bv18nibFGcvBansVq3njd54cOu/WW6CMqcNC/53FKL9bo+8vMGcDrE4
EQnVfZ6mt7rWpzeohCaRJNF6nm9FwG2/h8n3av6ksSjSmDkuagFe+lZx2w38
sDZ7gOQ9wY29q/hibvPEZEy7pAd+2RnEwV0t9+f1IVbP1sgiYNZkz5SKeo93
TRH/NTGt+pw/yHpFP82Hs9taY0bpzQ4PLzyoIOkX4VDrcySkBE/q5yW6hYhF
58Bz3m5mtpv09LLDia7UssL0oJqeaTPtiwzFPtMk9xbcRbERvwKtiKbnjWu8
zuhV+adQKgkdDcwWScSVF5afdic1WT/q0Grehro9WGc2iG889PZirjywMUrI
z4QfnpmjQUL6Y59Y7xug/mkhjx3zpAAXYmDN6GpTETCDcHtnjfA7/pVP0soH
Du7/Vcx3gGgl4zJyBQf45OpQKPvbDP4sXJUO9RqK1v7LwmzI6mPVPh/8OdA/
4Gjg5R+VmmyA5OEDTqnLYMYP5K5JmM+l8aFnU4OEh+ts0Wzpr4HoqsFFdViD
AL+DJ7lEIj8T6EPv4uyz15QamakS4EOn6ouVeKtyhNzEA2kmbcLVqkHhjdju
2qJUdYFWBLVv/T7nn7681sEhlUegvXDB2cjj6rotl0fspIPatdrAn2ZWeMs+
z/eIcMOa62Q5nnDzrC104snuOoTM3GBSgmaAtylBQgt5lvLlRNm503gCXXiU
tIHtvQ8AqxID0LZlMI1fONx8OkETGxITUlQ6BrHd4XCDHhGEoiW7oNuK7CzK
pmC6JWYqfdJCk+RTLmnjOtwX5cf7Mramh67m76Q0jfavJCUCRVQ2xWRiMu+2
WuirtkDqkQDvGVebb4G+UUqxdUjiKwV14109OZCicIwt8k3adJydlI9Hj+97
G7v/nAe3BvQhCbASIN9KNaOfFckx2OWHQ1OOUQ77whDW2MGHyZfSpx5t1zUu
aGqHZOhL0v+Y+gKEMzvcUnwL8oM/5NazWD7AdpqTNqqPTny4hQVjFSUVTZW/
zjobLc5sX24E6eJnK2IESn6KtMy44/yHlc5QLjemLLyyCsNYCeR80E1MsLDi
OnFLED/AhqjTE/ICDwDIp7Nt2n9Ud/0SosJX5bDNX1s2sFoQXYCsDm1HyUxF
qv1SB15dx6dNL9uHsi96KIX7kvG5s/5XzkEEEjaINdHmRtuT5A09vdAlPZa2
RWDZp7CuIM7Iyj5l6le1Vhr4pyK3Yft2hQBsvryb/2STZgy8Aps3IfA+6ElV
MnKwJYh6/ZW+/w+YpcLgMA6OX/TIoIl5mnCiNBStYDvPegBz3Q/avbd85cT1
Gm/vZhUAwGgevGcxCw1V3EscEGn1f1BfN0tupN0jwfNJpLKTogIUeSsV2oPO
qwEko7hM8VNYWtE5GPNV2DUmIoVegKdKewbARo5Z8vtKedw0Mmkys4M41MSL
Qqc5WrFgzLDWiMhSh0lmPFMeHRf+KNvgxPzzJY4OQwMgIKtXcMp3ddJYt65L
LOXXJpUIilhPLaT8tvz45ZsNa0kzj3Omie6Io+2QesrwLN4BA0lRrFMvRuZP
NX1SOx6Yro3kjvtFtX0brBMVrDJ3YifGx0L5veBxRusvbAOZoI+AdgQhWWg2
RMEVZ2Zk8/+oZnyjCjUVuw/CPRRE7vL4h+uNUB3dW19PnwcMN3SzzIT9u4y7
QzoG19fznDLhrEJPsUF7CUx/kCvxH89xu9P6ySaiAr62CZz7uUuiqhkFVjV8
RFEkPfO6xPQv6UKpT078VFEaip5zaTce1hqLOfegnrQLKA0IXQvCPtuIGGO1
RQs5WgEpoM83ERnmwEJsVXgVCbDPQ9QdZa6lymEfht9/c5WYzLbWrhWr+xnC
SRBQHUi7PkD0dh7IANEcctxfRV/AMpcv6q9quVulH5WN+/JlQ/fs53d7p5Lb
D1KYd4iNJqm9KrwFPwETDU/LxBGvcfcWYsN/HZAHtypG6KoQlt/O6uygUBr+
kiCaizMegrcW/AAybssz0BrZWsjVMqq5NVD/qpNCjLQBShD3nSLdKwj3Z86h
7BoX+4X/1MD6SO+mVjsmDlRWhJ8LZpbP5hexbYjweK/6U5mtEHuS4EJRZGs7
ZBi/8S0lF0oHN5OxSNGnp+btWCwikbpQryChMBoHohL7jnd/TrXmRYPlFWvh
VfrheBkaIoH8jmNsWkEuh1wf1kFQ4TtjI/Sf+VST58/MldxucVPNPUxWytfq
/QlU+8SeVwDRk/2iEgT8sVjaIE3aGIsqIyaViy1iWw2jmnTo6XvjblscJWV4
JDw6M3lykQ5DigbtcHPAtss2BAGotCVNAUoqCRVI4SpgiXmKcAZpLOSPMH7v
3gr/kRvcY/9K7wdF5usiJ98a1X38CTkW+oIuu6numEjeJY6aSbF3VhBHqX99
j9li6pxR9r65OT+ChpgcxWUiijyWTmYzoDKMiEhw3YKp1u0w9ezFie+GUI3j
iNROmznBu15VoX2Uv5B3RiJIaKMPmY9NACzdD4zdMr9E0oXZ9HYcKvahETmW
XS8ZwlFCbIe6/DlHmL4rBvZDuZIreJr6PjLwJgxgC7GTvdCUpOUTlVaPEuzu
Ou9nI+OupViYQRz6lo04EGXovyAVn+/o3RFZcYjTxzqocS4fCZj0NPyRD9pw
UcGbyCyj2uh1XMhjtaK0urcMw8MtNSi2os3paNvVKmrhu9kRj7d+oR37F3rt
1zARDdgz1GGRGfemACURtTj/k7OV8NB44EGDjcd+S30du0c5//p5oCpLGW+9
Gvnmo+/wj0gw7j7dIvaMn3NKR9SmaZnnmPV+UVfwoAKBZ+Y1t7aksyiB9qGO
wmwbyumLbo4C0aNFn+NSJZsJnYjpiakhmCZjtTJJfsUWcawc4BGjAfOFneU+
bITgcb4ZPLdhN6gRNR2ua+sVfm9yBW01xbW8L3V4alcoPchlmIzE87CHX2SG
tT1CMhC6aPPCIkUaw3B0rMvgQYUJf/nkEywus2oZHuBZ6RCfFlkQ7CRTgyop
fuLTXvbc2sKZbHWHnl7aHEmkgkzh6RD5gjuuwKsauz7QRSJCrFh/ACHDnT0N
DSfYVUGprWWP6GtwxYyI6vrSqkUbORXNaZoxe3hSXlzUE/2nPq07rNi/uXCU
/tsx42AQorrkpJcHZiWvMDkUZLSD2M8egRcPQi2OrO8Qtr4g5WxHicTzLvF1
vLeLgk1UXCEyT1sF2wKlE0SQ9jYvlNt5cdwrErPcD/ccHQkzUe8SqPaggmva
Py+6XsfMHnC1qNAHE5IzATwD35LFZiImn0x7L5GbOQ+N+Bhrse5WdvI+EywA
hGAeJ8ch/BIMf8MNqqtwGBvpHd7CPwYgz2UeIyCY/3ev/riCVPmJi/qVNJRA
qwnga3HcPmsz5BvWend3vY9nbZ3wAQqT2xPvxvxI8D0iqDNT7qxXkL44XZBh
SPdyG7DFGUcznsqb9IOP+/McCaGgugL+gh6VqWJ2Gajm4WcEcDlka5bJFz9U
VnnVTmYiAPuSTFt5VY7TNzTkXAMdorW5lvrID+St0+5D+/Cm3bTprvpH7MUD
qYo0ivdmhQVifp+Ffg/5iLqxkOzDmJFsYylVZHFN9ZBICLFm8u4w5Ydke50H
8Z6UI9D5rgSnS7CJycmQdUw2MtsBSJxUeJoiqW7vafK3h6PXzdF+VCfG1ggL
UVLEIuQK0+8WrarxFfo1fVtpXAfRSLh/tq3s8PExm4nbq5gT5YlvrG603MEq
LWB9djMN8uJC4ZuMlsB/YuHtCT8HoM8gdqyXzeG//afRQU41NNgvm/4eWfjl
vBj8Tg3QTdigzoYwUzLdwQWRx7t9UqbF18cYKP9fgiz3oZZYZaf0WkOByLpy
kRm9CdA4kOZzplewyWJQ7Wx3i1crxMQsvVb0sf7hs+PJQOfc0cBML/etk57D
xgzuUgCM56etzA9N+lCe7cctd+QCM3GvUxqM7q3e9KzbJ6wjMlaoXoTUhT5F
AYF9YQ/v1o5V48G4/pk/Y/2NzoxY8o8Z/rP1ndNS++IN9Eku7ssRa5X52TEl
6GD0TWw13/CNqinpah4H9UAgrGaqjOYgjZf1fldYSOyYYxqT5vxt+n8jdACq
Z93ALW/qkv2i55Vopefp5t3sCNFdTjMXXIvOjZovLUyK46mSyHy4K+G5tH9s
9EafyRE1xgz7ush9gVQ75vLHG0vKf3TIy4jeS+fgA54PJRhGgmSwfnBZExML
jYNjJTuzgp5qB/0HzP6RnDPpAMHjb/m26GFdKbpsqfIPRo7Z/l5fYtMFJr7q
cRO1E3taM5Md31Oi7rS36RJ3I5EwS9dlPFyiBoGnAsQ3e7UFLIgiNaMuMG+B
mVyhilqlj4kS7p+vvgkpM9up1lIaZmBvW9f0g7aci9PyVL35EIHlpmucd2DX
eNCVJbyvIsSl54g71XOGdHFeLL9KIwm8LmTlbUlUVKufDLTtMn9izNOwXyNT
dWFT3UFD3asi0dUmtaOCxmphtV1UCyX3+xY8Q+MEBAOcZl1SAmbMm7xqFlni
oGlDWhkXNzGcsoVU/+myFFRou1oKkkAIYmQwQ0nRsG53Q0+ZFFV8/G8SoZpu
nzkw7ouiZyy0J2Jdx4Y4+r/YZYAOihtNq+S6qIIVJbGcum6kHa0hrEc36p5l
PBazu0wmzbgg6hQs7SL9UQ5Z6QChqxQKvRrCCrw9xMFLVK6Y5dujdCAGahPg
aGgNAIryZQZ8F5hp2Ow4/4Y3GOLHp/ndFMmCZS0TKLv4gsozc7E/RzPFtI5i
uqJHDnksUV53j67rgWegEnr0eUtZdqXhBbGL6Y+3oCzpckmluEFCQoFaoqLX
b9D9k39WixrB6XtBpaiLY24iDhjcBPJ6LJYuvtAVfKsa97E2HDnGi4JNOAQQ
8+680LAop+b5g6EynBM7tsL5DwDuH0Pa9I+++qNW3dPPlQ3mzFiCyUTl0oq6
pkvHiPXkvQS507HIXQSWa/awivHqgYtonEA4rGRSVm8nJbD91T/4Lpw/2SGM
hevNUaL7BonsDsxQTB7T9xIAoXTEhUTqFEqa8z2m9vETTzaQOV9xHYs955Yg
yVB0bf/2NBCVAEnP/xw/3/Zu4iGkHfiqqvkgZUU/LsHemZtbYY3sSKJBr2M1
1d5i01vXRbKKD39C4qLohKUIapuZRHyUkE/ibrxTM6j98ENI39zF1l8OhKzp
F7L5LnPN+nZAzuSnGPztWFzLK+WhgzI0DtK7DeayftS2TooJZn/oNB/BqPO5
DF9rbVCE/VBOceJGPvHBzyCa3fxVcJ619/6A9X2ZEbNX6Pem6tGfxG20Oj2m
qkG1w1mpmabcD3RZ3cy1M/Yj4IRUDZmL/GP41dFbCQeXBrVu+73LyLB6GBXU
A50GCL3jdCVXFiijcSfeZbfo5AafSHx37y8h4c3lio3yECGc2aHxYV4aYkAH
NkHS7Rit2H8RxhFs7jCHQTQk0FAcnOCXFUVGgZ7ByRFwQk7C4harQIshwt7v
wSkviQWojYvraJEiNY/Se5xejV0ZOqjNoaMWfKu/99Zkpp3FST3Wtm9yhZnO
XExNWWJWtt/k1uQgUIZ8RgvSH5apM5jZnmSdPCBNXQMoDdAWXD2Jro1WbE11
fTEqokHjz2TdZVl25Oops6HLZfmsK1ftBmMHA6iXY46t28NHed2kQ2sdBhl3
1oxdIN1w9OK73NFGKM+iDMZxq5U7rc+JY5LPkhTfc/ZIKZjsVeZnS9EslcQ0
jLTb7NWxYwd4S6gW6qGru5bCFdy2Ea/UoWeLcFFDfrLCxrqSFqY8sacuiUcl
EyQEdr0FmEZJGFsUJzhYkqdPXYWIf757t05AMlgqnOidUjMAZ595bT8velLB
BYuvAtkRPMM7RBIQcGhd21nL8tmKPatrC+j6UZ7MhUA0xOO/kJyIl/mkdH3G
hxjmzMvPqTghcNV/z3/CzXfeYyjUd5Og46vIVeKNZSw/63cdr9auUjAwO/Zu
wMbA/Xspn9nIP+FPud3+NBpwwBCDXHMnWqBPll6JhkIxl5a0v1rgPUvaGibW
teA6TDxbnlj0D741G5Gupyf2w3R0dCQj8PNv6Su6b42+9PZz6bXp5wAWPaGU
bzGCeOnPF4z1nWpsL0UIC1iJfNLzTREU9hIsco5bUM/Im/CE/GeJvb36Q9Mp
7uvcFDk9+qV5SywMesJZCeF7OuQR5uHM0K0R8rUoNfaGoW0iD8gKDQXS9RkM
QA77AxaBvjAwbmXp/nGgssEsv9337FhvnmYYVPPXloqvhPFPO/HZ4FUDeriA
VV6f8wX//HU3Vo61dyMzEodKnw65xS0dyje3gjKpBDWjq9dk7/aiEhBiPhYN
cofYQirmTbE6kHd7wto4WaN0I1Q6j4lejDMzd/7nIdiis5mK1wXb/TusELT7
7uslfP4hPznfkaIMbmupTLHvU9n/Cz4MUOorp0D0EN2AX3lp+T+zvK0DScd2
B87ceMwX11NoOMNXIntd3kw5dNGh0Gw+PjxZAACFgtaKnN3rOoqc2WtPtQ6O
wnRVzJkNOPxlL94gxZCVh4CC4HjTpKbvYpsRcXvMxmwYNpZNEr13kbFZtQt1
buzwcFjCwIZ0tFV3BHTC99HEHmS86T9tL8RtZUAd0nhsXQqPfArNT7+FxgXo
H0PJLNcGZWCHMPncRNA9FcliKMVcjWF9kj+yyhz6pdiJ4A/MMXf8KOoMexpF
YWpXc9pR1dT5euO6bVdcu2FWC8mQNSz2+mF7fpkWNruxPcofFnWPZvmsSddR
CiL3l5TG45uxWxD49OwThsQyRlMKJB6f82M4xerjWFSORlw4WzlauVMI0Oen
adiZdvoL3/8JeUdl20IYxQkmJFooSZk5wfy0m/TOezxZ/yriBrITtKkSDpt1
awUPhWSFT+bFbDbYBwVFVnTRyn8XDMKemLTx1zPQm9NUH6vgYOXN3aIm5zpj
QQhHt0RCXRvPOJq01TdhtI8C3KCRBk6ZlWDIbltpsvxDjl7dQ8BjBUr03Xlx
UbEvoaCW3lMmEKQx86o53fsza/DcFSEgivMyueculB7T+k0NrlVXLng4nG9Z
2t+hCKshrRSqqaMEdoR5aQfpLeaiYOgNvvHa7kSPRYN6LELSriNFmMwgpSQh
GE8gzddXC9Zna1a/DSfhTyy/IYAv4/JusrQPsL3QSGyLt2gog2bC2QkuvA1P
v2J+0G8i4nMJz2X16uaEi2TYNmCUMC1nIpeVKm+/OFcKrdaoUXuukrEV3CxJ
Y9l30w9XNLYZmjbT2NUm/+s2DtzYpbGD9rzc5a+ehNZWZz2os/StRy1tqZqz
tvXEndejoKrKWOrI2ir6kRdT6U1LhS0jVt5JGNPY87iPUe4mR1NhvpxGVwJy
OH8kmoXzlYvX+OQ8r62MitEQfhbrQZdVgQMG0Y9a6rFelCXqkJ+GGvmB2sKb
KdJZ6g0fGBn6fo6CtJXySifCqlCEVQ66+y4sgNfa8++81yURDgWOoJ6XIcEP
8CI4tEXU/fyY9hMI84kn2JT1cCEgCvoYEZaXo1e0V2HsgmgNodcf+0dxQWyT
R4I2u8T4XUhcUUk4Ze1NxZ+//4EcYToAyJPcvWg+Sq1KxdlPZqZdDNEBh8Al
JqyRR8TJsXegMlz8s79+8OmJ/kExn/3GH5o7J81wiCkRhAmdcQeGm89ayYi2
BQM6VfRed4EDzmMb4VSEJfagan/eu6CjcRVFmz+ez1nPS1sZgFG+OIWok1lG
1kWz4t9m7kwx9yQjdO5zikrstBhypw78NbsfjbtUiffP8mOLFA37CBJjoMmc
dN5gTHNGWV5YKxYXCOsGrsQVsB4XsGqc8jLu0K8SsWPfmHtPql0q+/wY4/wS
x9nj+Rt1+09gSA+SR84K/Q3cFAp4J9F2CgTxq+AeCGzpqZDlGGKImXMhIZkr
OjiXJ4++0HsPIhOaHqvCPbBe+fy6rNJaJfy10ZO/VOa35PQkJHgPe0SM9rid
ljBlEYZZGU49bkg03Fbqone7D+cMjzV9Xl09ZA0I1ahZk6ZPD1FDW0MzNRGW
mgfm+eWjS6n4nQXYfICEJAnj8in1+FX5ogOmRbHgXTQHq9aWVFxuJxzRjxwI
Dr+XObsEYgzRNvjJFWDpbUm7cD0hTfCevp6kxDfZJKQj/K73PH2PQOdrcGpN
UTwdvHvZvFOo0EUmE58REficvedNkSDG0gonlXVMGCx4o/5FJJYZLAk0didM
u2swV03yZabnZqiGlCTAEYSwq2kAmclUr/Yju0VNwu4144pwhNKsuWNJS3vz
k0/lvX+N0nWGlfCeNAXqjmIt/JLskvlcbWZ2DXFFlMtc2ZHZVtsgMKF0P4My
sMEUaIqIvlp3T9DduCwirxOdr6XaZ1foNkRSEI4FslwhHe7rhDHqld8MQOT/
xyD6ylOMS5WRGEO5eDtrsAWvuNCCOepWRlbERTJkzqYIOjuYRQdI15mYaMdA
2WgplitGVNNopg4F04lPOKsc857LN9AWIORlOUhC3Sp1Ecf9oFWpvhVGk34Z
f0tPXZAeGn/TxtFrxYXL3bMPIQrIUcZpQxpB38TdqJ9EDGdQ4nYT3AMlI/CG
+P5DChX++425zTAarJW7+JhgFDprCNBoCJtH8qxcTojp9+lKVsZnvxDF4t8w
oiJCATA3XtKIBu1JK6qbx7Rf/MhVwrbUEUwkEnTptq5nKu/M7ezaZW2/PP4a
TjyI1Fa3KoLiLLcf7ojRZ2Obo4+U4GYe82Z6riykTb4LdIblAShcgPYPtI5+
T0e4/L+AqVxut9iRChuTeaJCO27wP4a68Fz6ScIlx9Rwu0w8KNuGGE3OR+BI
HehIlNHZ8TmEhdmT8+b0VJe+6HB4PquE0dfsVJF7/TyWzYxi90tn/bjMrU0q
kzjytmAamBPVt9hGAff0PggCfOWV0OO4+HYe2++fQSuzpJlMCpNpvuDTexp2
UObYzmoO0z/VW/1IWe4sm1Eh5O7DA75kZHOiEuaXggWH81OsjxGYDD+03k55
u6DK1HdS0jR+MxueXxjEIUvk9/PcwfNGAIHs+BUViS7tY9hg/AwZZA8mdBSL
W4uPIxGh4+FdlVFWn1MxJCGtONp5wA6w6AW/FUmvDXMWFezj2nCqt9z4d5aR
x/9eVYzOOV+urMwjEGRZPEDfkgLh0yy/Ebrfrk307is4FMtAconrTNJgLMm9
VAope7UbnULwdiPPKXe9Rn42s0CuBBZtgEFglvjTGiY9o2P0dH8qvRO7binS
YM2CpI7i6XroeDhyhA7U6PxFbx2OQjVgxh/ViUMYJ04RJ0ZaO6w8QVJc0Jet
hb42m58jz4cb0KaEvDex36ODEGV63ZP4FdIbYtwHnPkoREGhMejje/vGuha4
UVGOFTxy1/Td7iaGQDlA9UhiTst/9tsGmdItkfZJMUnlrMOzKq8ugFZfc9hc
l3DLYqzOH2s1JzMvVJugS0MSDzqzRojJMRAyhJZIEs/Xjtp7KTv7F1zQNs3G
AaPznx5LnayxDLiLCovOru4R5pq6yci1dR9B0ASFQMLz55nhSOx0rn1tW/Ug
+RmJMVJTTgAGF1AZ8RG8e09EpIhvgaVGZbo+kAJeTPPnvZq6Jtxft6ZeM+jT
nuFcFP1tofYeO2eEMT9V2fRPX3DhTf2+BNBKEFR5kQNvwLe6nM0dQ84Wc4Vb
NX6iO381y0Q0v210A37e9neGg3lh8Wqdsp0aIskPA5F9aV217A4Q5kIdpku5
6xA4ot1tdZsuCS6lpCGHdCj6gzvwyt8Q2uUJ4gnaPA8LDlAZS2ZO03C8MTy2
MJA4COhF8wOfrZyc7CWqXIrtNpaKaTaVuyBjpvb6AjsSE6cAM6HpkdLpmMbW
E5KH4ggbRa85JS6hmSeKgh3KIBT/te7U7UezLrLHNmwHONy/U7M+nkf+0jAs
zeWIWz/aDdgtJ0RN2jk0hVOZZSRQbPO6bFiQZdQKvPfaY8biKAQZLW7yodHm
YXqMYkXNZR+2amtFkDiA1jExXsigMkTFVVEzDVdHMla7mRFAXxp1fZmcS5VK
dtgY8FuOCKYXhh0vBJjjhpm8fJLiW26D+/adHOPKYdWf+edfFrkf1fl05e4n
oAgFwoO0DWbh9YGhTrvaeKanR5MVVkcYx9yzTqFifldV7+uQNiDiyrohtOoz
hPjDJ59Y32rfD6SXpmNQ7lT3Mue8XZZ7Ha5Za1gVfKNdvHiDXHWb6HMsIJ6k
5w9al1kSVaHqti5dUWVV3DruSjV/wR43NY12nTedzgVlT/nn8cZOJWTFfhyY
v3CgWW2RDs1t4ALugfOqcpAWzBVdjjsAOTJe0xdW3XGepto/aKWPzYa57XTu
wsdBzNR/BYtWK9OnG9AmmcJL++6nrIfA03VlwLTi665fLdLkIUzJDEeWvItf
INMPYs3Xx8Dfeki2v/xz7ogX1P8IdywdZoMunRAo6MLOTCHirsbcjjgZ09sv
Pb6rvtw+PZp6SDKj21MHApUT/nEBV9olBCPsaHpreXfQ8Y5WqvhenbnKN6zX
bdhG5pSVNJRKs7aRCQoG+DwnyWZBowJ3AX6iFg+zTEdhj1Q1u4jkGsM8WyYp
MtEfLtBYXGhtqApRPtl2bBl2hmSZdVH5Iu7GbTBeLpfgacWiHcEl0dTAyRXw
iGQed6oJlR3EAo/7WQXtOTvohNt/b+KpYewcvPDHd+lMD4G/u11ZTAwBChuJ
FGia2c7kSU6/7VrkouIe/TSY2JkpjC4Ya6Rga6gFzI/s7TWgLBD8SrL6dgco
CNqyGYLXNmK9bN012YhsubnIWH4yf0YGbYxYqAE//l+sqlCEsBJ9Biyd/UYN
NhypzkKZTSv4tXIcnxn+4X5IzCNUkWv8EsfR+REfAcfWt5OryAJlmJuZSlnD
wU2qwtjevmglL5JJw8U/lgt9gTs6qoWFaVcmnKGIkVu/K0+R6Rx5tw0eJcGv
BpNs2HnuyER44Y6hEftH4UWJZqChlJEOjODT533hHmRjrHRaLCFeUfYeuaC+
nN8CAXfE2a7kP5bOArAYNv4g4OsW0uCHMUVMgXp5e/G0TUgpFHxlU8ACxxfM
GJZ5TWa1UxFzOzgDQo2mSR5psrT7KPF8eqyRVzYomma5ZO4LQKebudWcOfFj
Oj73+Ub2jdGtwkcFtm1RdMwVMr3NT1bJzFdmgEHRinrZaOZZqTyu8nLFdKAe
xQJOTXZmN9imUANgl0URIyH8mKGdDsgUFpcZOfVvw4KeBVKYBi/h/qwb57xj
j4JbzFXAu2eaHwBkrsGHPG6OxJd9UcF+jkaMk01TionsBYiUF6Sy8DABZiGw
m13c3r1V84iYZkof2HqXrUHOkukFbdJVNxh7ChVSzdNMp2N2HEkK35OmsA8Y
Ez/OHFK7ahx77b5+K+eqf1+Yjyi0xoKFJSBZMwfru/0NKt/P/SOA4/bljJr8
7jGmkckgAx5zA9ydMZ8v1zocPXvDP57aswIXoMRuuzVfCbL8+19g/4M8DM/j
ZRFrnw+B3lfbjiFWYAcoyND+3ngeOh2XhSmkY68QorEuksKPwG9CQXyAIRg8
J6LfNCf9Io1TrGdo907bFtY3Lmb6275mo/gpG0z0BdhCG+HXqYfkQTf/KjBy
Tes0JS+3C/lXfzxevhovIGhjlgN27y4G786A9DSoI8t9CYh8BqvDYSY17ZVY
jx5gNIWTEZnNbpSUrlJFBxFrz47jnrRff+wGxrPERME8H+ZZx/2LlCF+bzk6
v3bnTEgJKZxfeXWYCN+TMY/Hn2HGpbBA63xDjC/afHwGUi98VPOAcEepbi7A
FGk7SjO4L/ALgilSGCnPdqdpV4RWZFbacTD+Vf/zZkVifrbnbr/n52oBZK2I
AEjurk98fSQQ8F4K40C8rN84BWOm/eqtNij21+igFODOipvLGEMAcPLl3Eqo
tEnIUfw89ct7Booq3NFWCNrnpCbuqbYONVmHcjtSqlItwBwi/QnfLmq/nIox
/t58gD5/mivzGgGIM+NG1AAV8rCk6zDapFluyVyIBTjzv/Ww70T3viTaZTyi
hKMnkxrFX6oArmqZQdir5aw+cPiu3A34/9Qlcqga3y2f1yR3wGa7WMZpNGYi
P7Ozr86IxTejN3IxRuw7KuW+OE73P9jnDHQ3JCKz8nxrMNT9IyjudmYK/eRT
DgnSaGLbTip+2qnkHhlm//05Bj20kyxC1E7tv0JFc5NuJt3eFsl8stX+vtgr
a3U+VFwdCjfygfbRah2nYt41L+tiE8l1V1ljh2RXYZ1tYgt7mDpO7Hmn4x6f
PqtvkEtbESKMc72N7vujovs629boqvmZhyIY9ksdBLvPcXmxFbIRolS2AFUe
UFwCbN/mV+NsLmVDSsj/bpCxhSDC1Mx80pYgye05ghaGqZGIkwLil6hHLPhd
FfaaQ0WVnVq202JlLoeAzj/diwHeUNda51UuLw4nxZp7WPJPOFaTmaX6VZSY
b/Xxn2QxtyzVwwyIwYM3mZ8VMYhjp0LkmzcGfsq9PTA69Sz9QL+pNFoEfsna
6cUjCBIPU6OHQgsCus4EyRRLvldogk2XhCpEbJBUHyv0GHBWNpGQ+4kmcxy9
QdBG8htp16VfYgWMLrlZoiuy0RL7eokSGzsFep7xqjfdUqiic3xLC86BwpsX
Xfu+soYdjZZyI3d4GCs1/Z6s26MZ+YR+Dx7uVekbBSkxMLo/nHc9BsY+PyDJ
p6YOQvfflWSm78PUFQGAs6W7r2hxBo29dyHSJporxVzQkWLrcKbW6WzW2Ltp
A8i25yToCM6PDzX72nnPtTcDLw+qxt8h/WvT2fpRMG23zxLJ+Z00REXu8dAW
FhK2cHGR5m++4sjH1ErK3lzajrKlautEDZbLO+H2kOofd7RqB5QpJ414YAdL
A6E13tTC9QkGqr4JGdIVOD/BozZfEJ03njhYVO8G5W2gaJ7V/4eEIAFZQZyh
cghkN1rnQTsbQQybN/uqGMJvzfyeQ+n9oHmZVf6uHMK9uGH/C43c+U2mhrYd
2gFBu1rkV7CNIY8dXwLLuo3cTC21m7+aBzW4gDUdAqW4c5q1yuk7ymMHA+Ou
hiClYZEfesrXwlUSJxDXX5n/5yrqScp05ZoKpnTzp0WsbHOwqeiO6OwYtT6C
FqrW+N2wNm8XFW/4P5AnquoTR9K9hhRiAN77Bpfo+oCe0wO8X1N8IPDg+ET/
PQb96mRLBy0t6uLh3e/VhBYHJlmWJWL0FY2tncn9HdSxv48/mkYEfR9Mc5de
c1GeL8FNLzc4Klrbfij/DCJ8AM5tgrNq06zUic5ynd//MqC7vQg2mE/bJt8S
irNqaV0/QD1vn2IG7vqdBdQu23wFE5TcAcxIXL3OY1ru+ytDZDMce70TKPnP
cKI6dA7TNAh8XbnA/CIAmjCzbv4GBTEmku19Vq8ysZa9Ty2W5zOWx4VB60IN
U0jDka75PKJv70xhH3kfr0u/fOCF0YYM4pA5xxtFXC7jPbLkDxajeIZ9bWz9
lg1rKDOH51lsHuLov1YuRdAMtbZ4nndgaNqeuFUpboJVUU1SsEkv1klRlPoX
+sJZFjUjKo7jBJVQselVYnjPIUjuEv3Fdejc/pury2pJiHkFwenPIRjk1omn
Ydbk0Zwev0/kfwSMd+H9xHshL45iA6W7hQUvQNslzbgEeL4p/nTKIVm8QWks
/Nf8E852oEIjt5OOgQa3t9uf+EdCkDBWTiY7rlUd3edXEf5r7IqkZ/ZdMoGQ
G1PlMDkoiHfGWbYfJAIFh7kNyl2nSoajj43FdJHb09+xzfXyhUx7Ar37LgLz
o2ZOULnfb1dSpgkLq0gVdNSZlepLYEHWPIfeMZVXi6DQy34mk1FyPX4vG7yg
PkYuAgwYLHyk+DVBFWyTAG3WhOQgmpuLKacMvxkAQgOoLZVkq7/17Y/gbtMX
dRTNKRUiZfJQqmYuraApQPoMeV6M6DEv1OxMqFyb7ibAKGP9Ct9P/Dbwh9rA
fc1Lkg7sxuuSRV4uHEmUMRJlS+GWAsB745RQKnmySYcjr8c+/LUtYlWuGucc
qEiBGNp7/oVpVl87Yl17hB8tLZGe817KDs4lKUXs7oE2TavArSOA1WTQJa70
E0PrPI1vI6VAJkV+hPlfFS4IuqjTAHq60BTRI2b0bNkMb1lslCmVTeVr2q0v
lS8JSt6x4rHjFQtnbV7wQaj8348cd7H2XJB63tzspdGsrhDYTgzKZx7mVRk1
k4W6kP9RabZnMVADgqfuXWxThix6PAbZ8ycv7bBdE3lWchBTN1/+yKUWaB5n
AxZwTwTF9SKlz+Vak+X+LcJYXz+WgLoU+/K+q70rcD03liD9LD9enPY5Wn+H
yNdt2psNi2kvedSh54Qd8r4PlJxZSDqmbIU7I1161VErcDVKn0ZahyG+LaNz
M/YtqVhb0rYMnv727pMUxwTCf/ZPtkEIlD55Ir4+7fcblCkRplCvJ08EK4v1
aGSgRzO1/QERtFCYgye5lwWp8TW4y3Wbc3JXnTsbPvMgrvqBYa5ilY28mu9J
i9yFm/aK1anD7iS4N/nJQymE3MlpOJ31CTsHt/1lNQ22RLM3Xk9Ith46vl6/
yhPK0mwHxdd00g+3Ol+ZRyV+SrntC85G/tezI2QFpCO75zgYyViFMWT+BB0n
GkM5qo5rkWiqf9CRohjsFiWvlbeIZjxy4bdbA/Ritaw6uGJNmr3c09YQy1sx
QlXPqjo4SCJXSOET429cG4yRuxWxT9Tl+Q8O/V6OHY/pEqeZzsIFKzxfwfGA
Q3sp169V9vQ+ZYikbg6nFOU2AqTH9U3vCJd+8bY+TlUN85uOmHPMRQCd5coC
u8ABleswx16SWPGcWAD6zaKh4a8nyfl2gdGVqhlZKZxnrk/RP5GUyu+P/t4t
bbwym3i+oCrqPkOUqku++WTv7xopfg0EbnjkWSysQY9Zes4QqNPcm7o/nUO6
E7YDChhD37V5mUVvmLpf+s1obDrE1B6CMNI6pcuptAzjWG4pxdMX2ezRJQb9
V2YS/9gBEXRG2Vms5dGmJtSXh5zwK4KxoAMitFPlXov4s7SEGSpf9Gvksn3I
TjkNrnL9zRwIDwunAsrsQPIxeFzJYIjwODh2Q4dxUoCmwRh41jvZEcGbB7YC
2kUu8KonGV3rHr0/haY0YGkpovkhlHrDCg3AcJx6tM10IiMsSvzpHaKI9To1
DEzRfGlBYDQnlMhQy5i4EqhKkenfNcitta0VQwR7tlbI/xUiiHKuvbYJsTQm
veGgQeQqYNcsmH2JnVUDXCAP52Sy8HGgK3TYf5DxKLZMuDIx4/eKP2KWg2De
naZEbBr/k+Ur+o+7BnAjeS/D8UPxFl4RerIfx1iUudIRfMSOVigFgyG5nurl
OyI4KGWtnjxIg2bDUpBg7ys+UdAu/eHpK3T6CQRd3/BM7YtiEq4sizLhhSGB
/9lU3eKq080BJGo3KkKYEWU+SeLttJoW/WNq4En5i0KOppxe5eeHAzQeh5Te
4+W1F3ORaOlzH4e4Iqfjf6MKosGXWAmKlvozDPSr6C236wrzULvaoIQb6nQe
Rx8Dm9yFxHKgJnguIQ2UTgaG4sXSUzbtcYVszubLu900wgJiZx8Z5DeMDTA5
eScY3aszj9FPlOVMXCS0fewls6HkMYbBY4xwiaWkMbJS4vZzVm7JVSPuWuUD
b8GeMQKS21HsrwXlJRbmCNHobILGP2Lb8QAw8x5nufxpuNvXvzr9+2SaosxL
LTLLJWKx72PhOE9w7HQdGqlO9ON2SgXpQSjDVHMf17Ei7Yfk5APfP/1C+UYC
mmCLnHPyOQ1D7mdoh++6RzbTJxMbyRo66ALCtfUo7NEJLt+jaf8On9mc9MK2
S2dExjVvhhyTC+Uv2UIW1PBCMoJwyaINRdB4hLCUg0v8d2XSGY4W+TRffBxW
aRyzSXC14mH5hjdgMx9pxDS2dY6tha2CJZcqQP7Q77Zb4pq4F18l4g8W8k1y
ZG51ntpksTbcxltpgw0+1bA3Ev6uueGsLK+ngr1+eHhsOJjAEvJl1f3K41T4
VNDWDZbEUBvPoA/h1QPJNLROI3XiE+FrFx3WinJZwb/GTLWgjBk4C7OvJnMv
eE+fZzr5GoZ9Df49PtKHBhYwmty94myIiNZAzPx3AKPozC5mdPl/PP1bnV9L
z4Yl+Euc6FT3Jspq3E2OjZuKVOiw+8lw4lenXM6FobamdkA7Iy58kJ5Su7At
QdbJ0DuwKN0DAh0V0x3MXlf4Qg2b/X9u/N98E9DUZiXiothW0Tx7vHMf3zo7
l+ZSz2/6yydlBqqydvese+9z59+5nBVk0ANawacSqTqUCYo50Qd7PJ1xjUHB
tot34FVEIHNSgAMTH7us0kQ4r13zk3XdJsmTY7rpw4o+p+nAamb4+23NSqr8
RYNOGCZZN6vx1qs2Igmr8+f13l8RfpQBgCzUj6agnxD2/z6TawqSKK+JzP6V
bACzS+4GQcQKQntWEzWx7F4e7LoJrOXDe2SprddyDnIbxZzCNFJ2fX+KAMz+
dVnb+uvmCw0iOuePzCf2Up/QZZRX5LM/p8Po80U1VvASC72loQjsIiCtiDQW
/l7N6UpakomQQLJRZ22YSw9z2Q0oe60C0tAfQ5GaRH2SoO25vIJZYNvM6FOt
ET7XYl0eqi9xYHj0gv1dM1kaU17Df5yfWyo3z1NEOGCyLd6LayxIcRA/P+pW
ybUWf/t5zOQlHCYh9bThK3aZ0YFvVvVtKQLWwblkNMrInwIDaD3KDIbSnVr5
FRuLC6GvTjKH317RgTON/wbqrj9bvRufrPcoyAQhvrE8Y3aniq/dW5zGrz9O
7C+2Z+UjUHsAxtYbP4BkvjtfkzgX3pnRhC/0I2Qr1E88mEgfuPvYSYqu3mha
WnsPOb0HEeLh8ZJkwmhB+P75rY4ZP44CZz13UhvvrQ798CDB7G9MIepchgW2
/M3APNMVOeXngsQ3M8onxsSPDtveuK+nLd7m1o6E4WxU0mFq7+UPujPcRnlM
hl0Qlw7cidGHD6suPOPrLoqQQDkQHpFtf+jFhX4JzFfpUjJ6Z20Z0hkSkvLC
wPejlRae5S2PgtNJYvnRQQQrR6ykFAc1cPCBbUPhTHF95CMVw0dv9A8lK/Z3
GDtlB+JT45Fp94xtMqmU8xMn9eIrpwtQ2VedDov/J7i9vSfAl84HSOF90D6l
oU+w4W2y58ILjn14qzFvn/SSiGPjsXFtSX8ZXiw6jhtsEOU/Sb+oPMqzo4nn
HeArsCDECqZUCESIRk2nxh8T+ALOEqD8oIA1B7MVF+uyYaldA+ecOstRtRO4
C7vabRbPfjV81dqxDgHZB8pkegUqj3OhrkYJvs7/GcmTB8WlBN+CmgEZQHcr
PLyWJtlVDMbesCsF+xXksr3+prvyOF2x10JksSwK9rErLmkX3USIMFIvUMVy
SQWBee+k3OUV6HoQeMbzdvaVp7AotfnUa5+PMz04f6a5v5lwTMf9vvajGWWG
o6Mu5k0m7i6aF66Gaf8Q6gknNAvLafvY+eufdBSenefY7BeZCTV+TNMETFn3
GomFPP9xyTucWDD57SazOMxluPBxDBK45+d7FqGlmFCchODtsTovd5k4BtsU
A3UNt789f7nVRluBL+HhidAoldOK3CFo+WycSM2aB01dbXMv7h75OGNqZ/3Z
Nt1NzGxYWTOqz5d0m+7Noxyik7KsUUOXbnWGHfmVvFbJ/aUVFeHpjZeCalzf
dxYGj1B6tXM7mikncbdEA2nPAsm1FAxKNLo5RsCq/U5pXAm0RLc2thyGxLN7
gymhCReRA4KzT/1b/4NvrrpqhpK+HcXxPS2q9i33SbiRV/VwUFlaWLp4f9XP
IZo3hI2svRdIEMkUTTjTvcvoss6aVQP3jK2u9CJBE47aDN8zfgevWNCQmG/k
YylbKPOPC3EX5JG0D41TYFNxeV0WU5fM3kja61KCCKV0w0P9Hbzi/eZSUx6N
hoyWbZvMDAR0LI6amxjmI6h9Ddio3jPzohOzDGLmiWpPft52EcDj1DRTCH1B
6kX+Ypo11Rhs/SVrELP0nNRGl182rsuOt+dHxMyi+c6ozJqPzrZN37q36HV2
9ie7/JFP8red7dkIc+yL6GWfrrRYlw5RyKu57Rchef1dXhVFlVM9bcO8zm4F
wa44M+kxn6kxwhUZSr0lZsrCe8TVaCD3ODNK+G444ZwFgYGhU/k6tWq1E+S3
Ly8IBSjWSQRJwo0a8/185tfOpY7poSWEaRblKP348gGZ/nrpnlEZSyVTt925
2AazCcyrdj2S4XT1IhqnhO4QMenP2FDj3tjbOtOEPoZveedKbyqQN/qs5XJM
CEzIXunMzt5Lfy7DRFHZu6by5kM4Fu++LzDV/HKSasynA9T8EP+c30OynV28
PZZmvUDsGx9A1r0Vkz05FQTeI9y1hn/sHrmOb0+2Y0i5syM3bxFTAE2AAbKs
91dkO29BNFoG2Nz5C47U7Rkmn4lgHIAyVd1PBSAopcEvNEHjhlD/6sd2QSeL
voPunRoxXqTzhj8xJ1HT+83h7bRwuA6hej2gRsKpAddqb5+/74T/klZg39Ei
djxW4xFwduofgZhlUPn3WbpxTsqucYcSXf1M3u9yWahfTyRrx8a/QDE88jhJ
+rUT82+epMJPc6+muwdpLeok1lISfEaMuwFXoDjF/I9Qg1hMwVP2hwFl31DF
eoEVSHtZrLmUlV5UEQwwIQn6t5tseyLg8X//El7Vd+ANhWDxosEU8QZULv2l
VK3aBDwg2drdRhquh5IlGLthoumgXrk7euaAQPpZxSueV5LpjnW1e33Wpxgz
46SFHGXitzbJwDkWo6cYj6OnbWEnkBnSM17DssvnWX1geG/lajTlA3b69+CO
s9Ax78WZhsldm4k9wzsSyfwd7QYDbToCWyt69QxRxXMLwPamoU95sdQV7wKs
bzdL6nfAQ7+aSMZZT9444DsGIhkgPwt+y4JC81NZDtj944g4N4l6Yj/EM7dj
/4C/6ZG7bp1+qu1Z8NUn5+soiSxLCdLtHZ7qEINFpvlV+rn39taNilA4dXhf
93vVKGqMg2+4wq0nx3z0dWLQvW1U78N7GXhK09CdWY5eD4tBo6gs5sDhls52
ZrkxO8+w1rQ4Nydz74HVncKgh9p0uOD6T/Ire7TTI42GX2Vup6Y7HEJsm5YR
0iiBGR2Wpq629vgbMfvcNESn2ldW6wP2tQnlekFEE1EnsAV7MdTonNMx2WDn
IetjCO2RNkmlK9InUSsUc1MYZI3Hvth4Kketgh2630CjVACo9lNDZeIIgFPj
Dflhn/Bc2BP6QbRETlzlb/LfX/4VHPxQYqn8vsx7OY1tOaGiZPQGy6sjtChO
P0yqn7Tm9tn0Yg/1bGKVtpmhM1h0m3MNlopU9CsuXzGFAeHsuRkUu60A51PD
nabWgkqn08ySqHWHllKw4HG+wr7DVV2z6L73dDnOWlOZeM4jXbPTbukLwsGa
fdljszoNJKOIEiFcId/MJj9s8bgGVgFtorgGt+zSraZXoE0pgvLa0bWiYXyA
aqtZJUuzhYxUWp2gkJ388EEYro/oitoINhnxSDBIEGHS4SltbCyeEJ2OAZC+
ivP/9WHuT9AwF/7Gk+JenO9lSdf5Knj+c2O9NsmuGdL0VKGfWvBZBdAivV2Q
IRdsnZ79PBI+rE3Vw3QYIxtYukN8Zo8nSJEyZb4PoaqU8qiAQgVG1zmDK7DF
6RuCYSxKqEJd6zD+C394w4mkJX7OpIOsZ4j5CcvutNKB0KBiPo/o7qBABYX7
ii4kdTLdr5rj8LLAsc+2ow8sASSCNItK85anGyV7C78Ym30ScRZGEf+mLEZ+
RuYomctelRYUioXuGvV/asdkDMfSLeiTxo0KZevnu7zhkQTgp/CaI9j+XF7V
kWOpEOtKU/r3sJXjacRfyRWfqq9pvb/jRLYTp5eDCUj7nSzK36gz5Wim6tKM
AlSBHl2k8nR+ebmgxTjSfA/mPFuyYQ4Lz3qG18gXLwrvD/qUKKvCT84A04+D
n2ViZsCvhfV9er2P8MNE39VqLvxok2wMhmAp20pmpC9kceFwmggtzRF4mnwQ
BZC0YpXMwh2uBRcs8L6l7+R6KfOc2Sobkvx4Ioz33kHaGfMhcTkXzgIxDvUY
P7g88AINA/APhgD1sOeSPlXOtHYHnxL8maQkBHFzouB778qE6DpmAKLBSSZU
hAk6kuzLwBIg0h5Rk7zS99v1SkWzo8cCoYhY3f1OJVtWrmChLQc/V8AvVaNA
+hgWPUXDNk49cJGYe1QLmBiuH0Cu/Gw5qBlsUbE4i7CO1I3WtApP+KDNIWOL
VNPIV3xC5FbAVmNdB59g69n1KsylWmSBpRr3t/IZNCWtBXYQUly1sWzOfuNV
kcsxSI0liN3qUeLP+c2jhYWSSd42VlihPA7HtRS3blbXt5x/eGBXwty68rDg
/MRdOqf3aAgIGT3z51joYSm1RAm+R98IGlb/0mkC1ZbcdPAKH457904BMJMy
i27VXQAeObktva7XXLAxSj8zt99TSzDqjTP85zgcrVaJsazGQca7mAGYaVAk
//nwsvHl3NYIlKh0VeZmMtVi0FCDeB0WG5HbSLLtvgYRD594qSgm8B/QqF5X
mGl+0PfbNDSUqruyGyDxznmw5DJSrDhAworuKizAJKOdZPZ75k9tc9px1lFJ
3F6WJlVHCK7KaCAHm8XFAyj5rsOoOXHtZO2Fv/VXOFfQZhQPZ9Ux/mUu/7S9
kb2YSHUOoXEVpA2Zja1hA0hXIO3JFSngjqWgjcvRVkj5mhw7cDEOQmeA4XoW
5SUD2BTt3MyY863hQixb+RQ3nB8BUjMk89HULPLT66bgbBQ+/bPaz2lF293u
WQOj2EmGjRYR6yc5XTaq8HKozRz+c7WL1KWG/0LDKlKY+lNxomAJyGwpLn5T
t7SRj01gZLQFXzV53Gsx9fqtJsOZbQqjKuXiy6/kYgbsOFWA7D1YbdvjXnir
DVilXSh/nXnQwXlwjOZhkNQqCxQ21K9SmbrwNSx0VAx0BaakvS1UHRRISWxM
VbWiS1mse8EG6/SYySpdr+9CYlQ=

`pragma protect end_protected
