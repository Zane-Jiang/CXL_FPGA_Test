// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0hOCuDuzuKiRlfwGt6M5WvbeO01oK7fs31kfVDzpZlo4iCYSrSDrXvL3xrx6
7MNMWDM0Xyce3ueMZqAixOjb1pdyVyu8ZpUpRGUms8i5DtYAjSh8gcE0XZvI
Snz5ZciZg2kv5Q1zIoNXEYlTJU5nqeDhdhgz/hUWQo/D+6nhMetVJHOC4UGz
G5qLUZ3DXfHJ9bxauQgd3yAjcq3XXjDaNGLKRfhgevJO/u05tzOkEf7iqpgN
Az9hUwpFMnzxqQMY41AJU2FKyj2lgUWDWPTpUDpLzv/jIyn/UXHTAZaVUJTy
7TGdJANdvhGMcQRmfkCOsQknAckH3TazcqYckDeNgw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GyFvga2W+j0twCzN9730GOfux2iXcLupQTGspRHjRvAN8DDmdy59nzbNNUWj
OT9+RuZ7oy+4Beo6zWVZkqx+DySIely24ieniazbVPoF3KoNObbumt+Th7cJ
wTpqJoGZareK7VV7mp0UyKsx5AD3TNV0GmEyGXO1rwFekoBJnUWxIns2y2/J
hmdI6oDdOhx9unc1FbM1H+Z8uezvCNF+Q1lxQk6EDK6VUinGpiVCGb3Gv/PQ
KjyXgaNn/TaH350MJQeS+82tLLwEG57gO3Ia41jC1q03mRGcT/UYuOKM3MOZ
6fW0qCAGDM5deWGnNv+w3qWG9dok7wutuuLtMAeBYw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BQQFBEhRcWTjbZ2xhp7Da6mMJY5T3UJtcaGNcca8oQZlc6RB1fJQ0sPuQE7j
qaDs6xi/KvNtXAlgnk12+GELms+3hTZU2uu0zYwbnhW/2UhgbCd14CQ5XoLj
mC5+rlV6cuQqqMFzWwkAjriNYwv1+9vRbGNGCmsLM1iOTPI//4/wUmrqkB5Z
x/01/jVGK63UsnH/xedkDDV14KmnlJCAFcX5dU1wKPz0MEJMwT/OSaQXaNKX
PYIUTPLBdHHnf5dgGO0IgbcB4GSavAEWdA+qVX0lHIFMnGS/KHL0ySgCVQxY
DBFtvotwq5tQabzp8MgcXfImGSGcewQImx9Vu0IgCg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MkRfY3omgXbS3+8u5+asFLaRiUScfJy2Fj7rPY15Mgfxc/Fm+uAjoPLjsqgL
DuJy4BYzJK6mwGdwPK6H54Y4H8UYjCcG6DCfl+noXs4LvUOkS3QHwV2TEu9s
SvJe61TyOe0jhlK+/6mU5amof7zlsBT0btnN1atFbE6q0nx0O1A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FHQNaM1DkOvBS72xYmWXcblSsJnHMrKK7pV54RZ9X/WicT9amCqLuNFUXZCK
oNL/AxEZKYdJKZ0rujjUDgTlOMtL9YgPly5hqeLWTS0n51c8LMggJiDZ6FxR
kecYKnNrtKpjd6g7BfXycyn/UnSkFBKsuRZwIvjrH345yxUGanODdgZOCdms
1CAt2mVHduLW6QQElTTyRxGRckRmrEZJegTi78JzXrsEBTOxBWotRWEFUXuu
JAkq1k/YasG4jp6F1dgF4suBw0RAI7ffmRSt90CEU1TqgONLMFBDIsO2t14K
YkpJqC8/5blXgJNrBMxRA+CFYzw629oD4IhuKrBDINB8PFmd3kH3KyW8Ih+S
dC5Dex3ZAt6HSbHxCcpHoftXrcO/Qr4ILB3O96wxG+l/o4DzYNLAPHCuJEe1
8a1fNHmssdEZ7NzpY911cTWz5fGLxOwWgTIj7LlduTIOXudNcM7Gs9Bc3VsA
OWfEoUDNug5e9F3EB7dSxIBsIJVaaDrL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
efyGR/r2dja9hTBiKsiSKQCEjZLrqlc4LAKGqrZCdnXoQb0WW6By5WOwHVJr
zC8gtHtx14Mcjev31WTEEJZIE3hprGFcAosGpWA3wOsfUpqKyLrs4KfqRbuy
KjdyEW4ifE/NbZOy+wILh4jxKMumIZqSKhXqUdRiBUqEgKG1hZQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eR2duLvE/KmAiZ2BDz8d64d3kBl7BLXVK5zxFLi43Jh9XnBhFwapAkvb37FB
wEmN++OqUGsksrpjGlk5WDQtBJMnjgKkSHV5oGAMln/uopYUkH66iOb+SfDT
LKkw2jYooLvUObZn7MXAAb1LNl4FcVlP3ftNe+0tfvbKQAE6AXw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 188432)
`pragma protect data_block
qAwSeFzG4t7IxiYoDt3GaHJHZFxYbwKXuKFPheLLjkQ5J3mQaA5vvaNBYDAI
4SFLYCpECA9PGUsC0nrCHfTVfNNxcnWo0F/p4mvaiC/vuezEZWxKeHdw42Xz
+xztNzSXygldfivMEjPsNSLYvKeyyQMdBHlZImSgk15V3ee0brTr7yUwakG6
9rqaJinI6IuPsRmEO8kucLENIDo6IE1OrSBdEPZFciWaA2IpkBjsybE+khi0
YVBm5SQJZxA+tVsR0QgaMe5qgVyUA2huzJNvhrjXPmqTR+1338ijnhc6U4dm
G8s/hhWcO2LGZ+UMpdxnk2fbq2622yFGtD3QDdmxGTrnj3CqPCwx19VXKPQl
1YrCtptX9a7QZiKuCF0OJi2FTeoFrgFi0TIvcYRT0+bvFwWnRWq4nbupSYA7
jKAwkaim3RtIe8qoHh8HLlA64o65MWlty3pOxHTY7PIF842X9bCueHOykaaV
PmyAwMVYQH6vcgFEKMdWqlN2ZVBia7jDsE7ck7zOyJhs1oCGiIjSXdiGHMjN
XueABcfkUAo0lzAFLfvUJjBFMuhg/BRb7J7E8fT1oSzKaus/uLQWrP9JmXzA
2DL/yoJin9ETbRiYd7n9X4PZyLVcJcOdeS+JEpz3b5ExeWKdNGMFAXTO+EBQ
SXMsA6oEoNJO14Sg8tOA3GB1ocSLV7NoBm2MXIFLPQ1hlKvZDiNJJjagsjjD
IfsxObZHA02oRd6lvgXuQ1Q/CGKcCNh6wund2x+FkH/siiMQhaLa/rbVSpCz
7DVshge4XG4w9Zm+3OzZJq+F9jC+0+Txj1rO4aUNFJfbw0cgC7W1r9tzDrif
I1ZVrKZRc9/WXC2DSnb8ySaajvJ91Ph/wWV0BcgW1mYIFb8c9QywWZCyFP+Y
W+3zp1LbkctmOyIU53jeBZnVe/1/f9ybtzTKnHCNd+xfkQw5ns9CYPs2rdKM
71V0Od1vyqt+bTRgBl3d1EcoT8pjW7pdrbuTBj14AabEEhqpvVctJXaJeJTp
fn2gn3J/NGXcDzpgBnIYTPYw3BEsmDyrglri0TZh0Zr965ujIifJDOvRxK/v
tC40uyMHaBRj2On7k6qSD/hU5MzIvz4OKYeaEvbrSUp2LQTdyyFkwKmqbWJ9
vx5MrJMGRyK7lE70kPZZcF1o9IJ2G9CB+VwqY9UojTO46zQFgocJeqdzN3m9
ybAZo2Zn6+fbTVsynzc9Aoivxhm/qnA1CgitR8KIxM6XXoDlC0/Q5+axJ6+b
g5mN41yLqwJy0XcWID6fQWUpg0T3O+XxIlvzAoAWcituojV4HPBG2sun219p
AG8VtDU6NhPb27U4eZTf6uIzpTcphdpSmIlwlhyGvOzBz6LgTi0xFijrSEqX
F94j1PQVOApwBK+xHtoSrovqsLgc5UTSaaMFqs/Bfm0aiuIvzFFCPn3/m4cQ
2l1tpspqoRk1VWlEN3/S1FmtbekyJoofzKaZXhtr5IlZjQXxvHSoPqnsT88/
Q0ueerQBIEecH13JdX8mrkGNh9G7GHqAAEAoHelYmVfFKjp3hnxr2drszAtd
r1CEoOdL5WGEEM6EOyiDmtay2+glM6S05b3N2Nso2yEbfTrCaoFod2roAX88
FcfnLY2GgQB3+rcbPAn57WXos4nyLTzqrR0IP0eTmJeYKvqv/3xqtrUrfQzG
UtGWJPkhdnVpSZJXj7E5cBvZDOwWR8esaJHKF6qGuhxOoWu81LFz7LnKrZgK
BxctN52Vyvx68GeV00+bphVpOYvugVkanCBmvoaAmNCKJd2/KNEJHVUIjJ3G
6zn8c/ovlrdCa7Orw3PV9kGbaButk/8bjIaanSOf75qBX0KOgXA+vAdJKRu8
wkACpC7NEfZihSV3aFrPHFj0Fztl9AC+tblRkHLGh/xYgb/G4tG+uvTLSoYb
ro9wYMHGRtoarLsDqspYzdbln8Vn65b3UEp7MItBmjiK/pwV4j/U04z+V+q4
ehBc2AA9woaSFbjPoEupY89k7Pfwo4uowMbizM247KlzUGK4PeqO3NGs2/n6
9op6W8vGqgf58jkVNAXcRKr7tfXnO4phiW6EF45EZqqYdl3Pbbi0Obh922o1
o9YLpXyTo6LQGF/uAuR58ZnTbQXHUP11uJCA1I7ICvodxQugrWjbcdq+ZubG
nRDzmFGVbsAQiDpNMvwQic5WROU9C91A8r6oIf6RvaP9T39GrJdE0/EXlkat
LCsUwUjEStLI7/vMIz7bLxJZnp2ROE6tYGH2zK6mngszjq04TjD0FhRxlDgv
7C9Ttxrhceifl9BV1UNXlHo3eAMtVsjmuAJKVWkI1rV3NZ1Xi9WnvHJpHluw
4pyhifoY38EqmevFcOfvkKFr/B6xZFzFWswnYdyW+yds/MeyYlaJoKJy9MK9
bxVIhUi6ktA7q7LtvXQJr1A6whLkVpPY4VbQcLt8QQLkKCwichnPRGS7dFD7
cdmT6jHO/oXcc/HuDgR6BCeXQSW5xYuIL4R8m2/rb+7QvZ7LCkI2JzbadAIN
aYxYGYgxJbOtpOnFGH09oGDPSIS6QQPQKqa7s9kKXcQaZDhYJfOn8BfY9WBl
1cERCINWL8qioBPTYh18KOocTzpF0o25yYQ8bZ4C9fyURw9KV0nGbn/VvXtn
vFwooPmI2ltYlDmO2Te9fH0k86Sypa5F3a2Sh0nX5f5tEqawNBn6x3h4S8E/
dKrRf0O2yFbozc3hSyHmFF/lIK5pYl2E/7XXATCXc0UILnxapM/SCbNQdiDr
sJu7MIay+dcXKUHJwN+J3eRWb2wRAA2O3vueU6qGpE44wpuxGPBOZ92IOHeB
/puz6t/oO8+pYAB+yhXefZmgUCJTuHgUfgXZY7yu+yjnQr5Y26oWMyjOYQL5
Tv5q41Nc3XWXDi2i10M1nYoTO1x1dieTQP9Jq6dkuDQWfuPl/LoSi+MO8j+O
tYxksvsNv3/ZCXvNRRNxUSJYA8zLz5pgA3Brd2LaO4mesS1sgQ41GGxD/7us
Urg5Mmr7vN8muEJDQsVQnFnMQjcszkubnmLqjDhzNnVapYKq/j9C4z/d5EEe
88np2LU37GDOHn6epeN4m0L/bMfM3KZdxV+j7D82jt+fm9L0J6SfUUw9Csj3
uZAMjsJhyw3hm7bX8kVnvdwdKcHiKtHdEjI533U/ID7decJR1DyxlLYldvNJ
Eb8vKKonG8IDEZVPNrtcVl7fTo7v2/otEEAzslHYK+njnxPW7mzvlcTIg6iY
DKaThy0ieJTswT0YkJz3c+Yy0zkLYKXVNpq1lvJlysEebVbPCp4v8pz0S9mI
NODxkFJ+H+FHnJeaZTcol7eZep5rM7Dw1SFogJem0GL7Fwz3KqEAFDyQuVeJ
F9CEkwYROHwH8OfeyrKvyAYCtIxP2ni9ynFzDi/Jt4/KHnRI3GcEugxAt6gr
wnCVXAok4d6+Qys9419eyZnTqdF6E+NsMBis2rw78jJ81OnnZ6GeYOwjkJWD
oXGm1D7aMGFm1Mvih4O5deuYvGzAOwfbsm/k6drdtI+8tVf7qs5SBrxGRWCJ
hHlaArMwnmsYNh6gDUVxb+/eNwEIMFklbY4/lLRxfKJhGdZi0EMvUN/Ik9HM
x/4rZv7EOiH4y9rcG/XT7kQXX2oeJICvuuX3UqbEzb7XYNNUMGX88mtb3FAz
8MjFyMSK7knct4ix0uKATzc7zFuxve9wdk8kkl0UbkvSa4JLkMhlc6XvHCfT
3apODVaOgYn/UWJ6ltGnTnTcw7bbp6ZfARo6FerK8bEVMJ4uxuQLKPuQWLq5
yPK7WbJKGj3Xx/FlXq0CSngZx7L1SC7HB3SrGH3bRzXFymI0awtaYL6HcdN5
uxnA8irfprUBiseaMaoawcWrorWewKZ4JZt5UWthzOCCtp/s5E7QFIXfuSeI
d15C4Oj34GEdGN9zRn1ymp2h/1xnsU2MC5+fpTFs0tPJm+UKofxkf/Mxrcfs
5R5Pm8FHe+9S/zkacj/m8CVoIjD1MhB1BNzZyoNxCznQ2S2SzgKNQE/ZnrUm
5MrfB4UdE7scgGRlon0ktmY7DQym7GDRGkqFlE700B/i5aQz8/OjS8kKlkEQ
q8IJ4yjgxkkFAl+wtVxAKKBE4GyBzKm7TkOTDEAZ9yBQ+60BeFy3YWZ2f7SY
5l+wo6ORiEirAEOPG1a3INyhu6vZleJoOs/HfRBChNfpvPd0lXrlix3rnZcU
NTFhUfk8AYhkFa7k2B9Y4kXetKrdNzdpEj88GseOhysXX3YDZaRfxMj+n+0o
5GuD0w3c1TKe9/j//epZjb5jLa5EjhSPv1v2icPiDETCwPEgwdY/YvVuEFCa
ogEVS93/OTxnBeUpCvY9GGgPNdTYuCIaPThmCEp7VXSwxD00cfBIxO8RoufV
z+T7ZNzUFz2ENhTX7MWBKdBRvargBTU/wd+dk7MKGAnToapVsQjZ7mgMFM2s
JReMToCxtnph5ghmsmxOLWJtObU0ZaUdJy6CX7jUxq7E1Ei1dhRlW9xqzMzN
Wprn0kkC54eggqjKpikWA64FjuVDCHlmmQLjsfT2qP87ehvOA31Xvc0Knsu5
qavF3TNK8ix/Ql7mLUWAckkzMV9NxDV8iWJtSNrJecUJkenvOgaWg93EB+vC
DG252vVoPzfeOZT564VQIrsrPNdTXQkz9YYas7W+lV+/5umbc5vf3/rlB5YG
UC7d7GayZbBVEWEgoTo/Ix8dvoev7+rY0uVN5Y6QI1Zgnksm9q2QprjTxTOG
blvX8aOloT+z6JhHPH2uOJ5eDUlYd9n/xNXgUX7qmATCQNKRiMrVlyUqhuTU
wU7weV0SL6sbC8MOfsrx+OMHwkgo/CYu1G8a33C5E2RpI8uTMflLEKeWfKvD
5BZA1Ejv37dFf8ANWClbtQRzNt6l9uEBvZxJuv26GAP/WVd1mkAThdomK0qI
SkpezqUJboNEQdCHp2g2MuYqJ/KIdgcc8jth0V58fDs6OGerSzcCD7zzIyHH
2fPbql1cAjTuEeM1dAgZQrPy6E1l8+Pd5Jj4HQ9vHzvs16o7y8kIvG+r4kga
i3gPtptKVsSpfRNdxyi8MImhjndTBG3eHXf+mjFpewsG/h6i5s3++VXe9Ggr
FLytemlgOiiZ9qEBH5gd8NcO5CedBA0x8jjxsypmCU1/xsKdZOU0nNU24VGC
mq5V3SnN6VGNiTA7QLAwCOZoSOiJLhsWbOhAzCcOsC3+Qb4NtriouaPp41f6
x5g8+Gc1QoCddKKz+/UxDORjCZiG10z8Id81ASQJ2q7WnjWW0pa4BsQeht+1
QoqjjB8Qnmz164LhLUh0kFBt/cFvOKyAL6Wc0m5d4crqTDGWs7b7sxpdkaMG
5h7apPDIX8lSKVDVaWCQCN37FxklofqDmwc5f1ronx4gFY1qu9zGBgW1NvBy
wmiy77b842f9J94DTrGDMDtfImM8NiMdQihq70PXjzqGphGNQ3v5X+kG+c5T
ZluA2/nR7nSZzjfUVciKvfiVD2gC4B70OnD5L5M7ChLw7FhBL2ofj9s3UQvP
PoPARJQNymTsLVzapojJLb29ghS6oxVyld5Bc5R1D9qZLBN+UROR8dO0QqxH
wFHgJ/WvXCng8nycU4avAi+SPsp7N2uYwDZqlypko9+eGT58mKn2lNiL65Gg
wdDUp16DErpENXxpQugC6zwLbtVkteqEDNLQ8pQS2125F/fHa3v0azLl7mTq
BJUd/EqI9AndvBVwUvsCZVLnKSepiEdOcry2L49Zzy61/eZT63x3wVqd56w6
VPejQPp18OvROMEMgHi+KyznZ/+v6sWA+dVBjWschcT1muJl7MnOFWRj/hOW
igkp7IIvqgo+n9lj4Tqy5S2jDnaDzu4rOSm0FP3++VfDNPnPxEIbjVw407Df
CxnhPX4XSXZu2mcxiKzyM2qS69Hv6NBlPf3GzdzfSpRV3Kd5yKujLk+Y1sVD
Q+bwxVxgKC4oLvULvxc6p3zpEWv9zG1XOpw9SPtibv5r0A14/7lKLvizoyQX
Jf5W5bi/lKeY5x8S/bR/Xk6wbe34Zhmw2UgDE7iGGwAue0Oc4eHR9ch7TOAq
KgolvKdIUa0hrbnaYCmYr2mMpy5n6N2uLXFc38nDDeyd61ZpnmvcLwzwfhCo
zRfVNgDfzHrDZ744gyFqxyG6vIEBnnigfyVPpVaiy6MMtkWYktzJmr/cuPtH
2uw4cIJdSpKvdiRcaHJh5j8EQYIwPIBbIbd6kKkBGmIr0LI2aY0wqCFWPmpl
3PiJhaLFYQwDpKirEckH0XJNQpmXX2+YIRvhKh4CJ008+frUrCdZEgjqKCB4
JL+H1MhLWgs9s08tXsvHHRVo1BjrMdrkIPsGF7xMfSw4atEm9BGWF8EO77dC
fV8tAW3yfein2W5eBKQ7S6z0ivuwt21kKKHygJ1aBzaTEEtNTpehQDsuD0I+
Ru+HwVOHHXGcB5eRaTbiV2NsdttEClqkv8m7OSWt3XXy81p6sCZq/gtO/xow
Dk1az88+dGwRZ0XMg2zWfqp5vnSTQykzOv4el4nWUR+1EPwLTF0KUWdNz8LK
Mae4hl/NEwMfoavOOm3KoivGfxEZBSkUrWIKK8Ikirz0pUOJqRm2NVQNdo4b
0vbz7+5UPSGHJa9qAiyhBHTR3NluJCS+OcDoqC5eAOSRfdyo5cqHoB0DQqdE
K6rbAfghdA0t6wcKSBDBvLHSyAZAkc+9kgXwZxN867ybesPQDJZpuSamDIb5
ifae4dJ6G4D4WxWlGyI/3AzDcHCwIP+zedQiJn+y0dYlYFZiT7T0yRM6z6tz
YOqcjcFd3799L/Cog5Sbj1UMIqbUmPg+2DdizDAivhDO4sqM7+nUEBHtF9l8
ji6eEnoR7o3qODrVH5l7f0rS0poGTAEFmKpCZsJeLefbVDTnmHbGo5CcRlRK
dzFJQfV7zoyJmpTycUF8SClPpDALdAKkGfx8B30meRkEf2Qa+L2cKyG+dj+M
zq5V4x4tMvBa3AA3AlX9SBnDIiSl/lpn1yNCgHCcJQ43U9ceuSOR1KP/xhmp
e8Cy+nuZggJP3K4xqmPtkR6Dlokv3LQ4au64JncM/KIFXhMxldh6NSX17GtZ
8ck6oeV4Y7cQXEj6QcX/vC3ykIC1+rveQBkiANQOoE/JZs03g9gXQjKy4WUs
siqJFFruk2npN0jvg4Kz8WgaZE18Lk6qpaN2fYG9Rt6P9mDgJxngYeeLDIAy
oIF6I83sb3+q2CZ8h+XgMuV4bPCJcXBB31nHN+9l/CJ5pjVSjrPYmCu6lh0u
0bkDml1NUMISk+9HH8HOQ/93IRe6h6yVskJmf51488Hnf0E/w4BVzLdIY2xa
Wy5J1lf2sfxakDbTuTGuFRfgK2zzxkpQ7PJHDTUsW5RbmScN2y/Petga1slc
42+iaPg68PtBj/IK8yyVx1CZ8GGHUR/d/JGyKc76bmafypnRJuLRf9xEecQh
A50UPEv2nBI22YdtP4ihD+nfyF+mHY6pt9X72IGHma2olbnwPQCpsYJ0AyuS
hiWiQnms+N7r7F1ccHdla/TXMVDTE6NWOMcAdELm6FjCzoCMyTZ1U6FlnUJQ
HP8EoO818OMQUi4d7Nnol00cPKKtLCI8zzGMYe39IA/9iGVxd60MUKMd9CHK
D8/jRkOMWV/YeI5W6QG2ktzel/Mn/46SSyy9vKLCnsLYlYLDgi+xrBhYaMoV
5qgV6xwa0QBCUD6CB85C7OV20HqfstjwZmiVo+9ayBTOIXEyHjfxZ0ff9lql
NIgqpnR+t4ydxQSjgHULJSQAqBjAu466qYP54qV8vdSoMmrKlcdPw2XqmBi7
mRs+BXYAJbeWycPpHJNTCVIZqUTJZfdcCKFAwFBLw4etwtKyguJC14wzKZjk
ax1U374DwXJN25Zwh//3WX+rXgViHMHyDNyMgDJjvCeyZfYRh/Css2W3P/8K
E9i4Dq/rKM+SAN4pYvjqyqOTKSmhy8JreEHAIQs6LUO+wWe53QkBCWRvPED/
NzGKPMEe9I8glklo/6HIx1Jm/+/sJxtdfoKb9JeyIDSV4dJP9mK5GkVS4F4G
dPWGQlmcpeZP0B+F52kULD+6SGQTpzIj52w8xg/+yh/9G+i3FEejLigye6aS
OUDkuD+ErHK2mh5A6wmNauXYGR1hCGSDf/QCkjVQGIvgbY8fo8RzW5WXMotR
hppcugMYvs1HNcd8v3W6eGHLVo7bsqR41UD2e1SW5Y+54lew+58LWTJ9fISo
OuTvkKlf6usnADnNQRH4FTk9Pl5Xc4NF/vWVdZmETYcAnUUXK6wgAD4Q3B7v
GzgNbK80qO9MTVp6QODqj60lyUxEji+mnhb2vYN8vp/AKeeuT8c4Dpn/eym/
ZOu24z1KEF8DU8ZmhJxIKGj7v/oN1irO6CThJBFO8PwNfcbnMZWB7e+fyXBs
o537jRpxAwr7H0Nf42frfO9vOFTrBACAEtiKowFpLTIKD2zjAe0YAAVsKYcU
FbJwP13fIK6gKzOb/RFV1Ra/6y+5Z5oDOg6Kt6oX29VrnE4CYl3LguBr5wEP
iSFP5pr8JIBvtij3uM5HbRZ/tdeEA5O/1rkWHehgkcdLcrK922+v8Ub/EIFg
ECXRBs6woW75yP9JS8XMMGjYOrEY4h4c0o15H9oJsR9DzZAeA10tsCneXl1M
VDYhooiV7xJPADlclt8S0j8GVwEG9p9ochy0krfQnnQ9r6+mbJd+oqGH6AnW
tuRx1toiBm0SzXqvG7CIcfA/qAWXIvW8xctMjauZAi2jAo+835UjFXoXskJx
R1WIiMcWfdadJbKB4GbgeHteGBP3UbtOJfD2KTDgm+1Qj6RGvrV9R38z2fO6
5d5hkRvEr90iCCXYvzEY+ZDGrAtVRt/7IiNnssKuwYbKcARddKLysVuyvlYi
WHcOaLiiZK8HXXMJGESzGhEFs2TAfO7aWLNlsIuBEVpKlsHSNPO0Wz0FLn9z
7h8qTcUdEs2e7wCezP8XIawwmoQYWugjYmkyw352HGnymEuNKDl2PdJnPYk/
IRFeFgiKjBbH/h90n/sd9QJp4qWfGU8b0M+u9S8L5vs66k7OyMVzRTYnGAiv
/sxGtMaUe842TjlIBWP9Pc6vSkMkM4A9lo3rzWX3tVYgCDjonJMOHDC/S55r
RQGcAe4RMViUSbnrqbDAMfyySOxgE1k+yNvzvISnW2xYqdk+eRwZKYIKcUBy
7fq5XBzxxf/hUNK/vPGDSdhFG6u8gGHbwP00SGxSoDcyPRop/8ginUKnp9JF
s+2AtGz1P+8N6jC+0WkBxPKY1SdVapia69jbP2lGApGg6GPY+7NFAATVR0qi
eTZOKqLA3fHb0FyGyP63Z15iNRqPtIzDTVto1fBrPrrXur80X561mMdaiBaP
QfUREnmIB2CZUxFyoT/P5yfAuP3z/6beBQd4LuYnbXlkgCSpNfU3ZQmoqwAg
6siSrpfG6W4kIzBFS35QhJeYVTC1tI8Kz+z4yWEBFxLy4dl55ogBkKSbyEMV
OxjmQ6YCHBLz4kN2TCxIlP/f09G4i0PtOUyJLNzImoCNMxoU0YeorZ908CqA
Dtt8k3L6q4Xx04JJ+MO3PkPMZniuUGeQHaV1rRjmuBOh6LY6SxFl0gVtjfFK
sAqrB++6kxfRngTI+0uOsRTYXjhNtzG+rdsJ0ESrKJudlxRzzX5Fnf89TZFt
5eZ1O30p8UTXB2JKPp5lYUvjbhwYMm1WnbpLPGzTVOWKGmUZOGaZ/xGhtedz
sV9YqH+btuLJrheXwxI+TiXBtlLtmVWJOdHqhafJ16im5SuCsHwMtbit5Rgk
uJQQib2OE0QU/b+l1lFb6vaBVtP+Nd9CkwmOqBMVDnmFYUVxGBXnNk8DSc6M
S0vazAse41xaSk27SUKWymg42ZcAqgoOYrL5IXrNC3+gAduibFKzCzu75sam
hI5wy6JVXzfHFoZpb3EcQok9gK0MHroCE8CeqV8A1uaPIbFixNKwgnkOwkzS
IHgtDHs+3BQ+uIY1nzICX3e+RtMplGeop28OIaqgBEKCbH9mpz2lRPNqmndC
kCAmJdz9JLYCINoTDkAXZWWXxcte+tq55Yiv+WULqVOi1J3/plPRKQsVpTmG
oHo8+fHkdVLpwWbhpokVJfvm5tPXqCpuv4EZ5jK4X/BwYuVw9EfELx1ypSew
J8GRvpZpV4euEp3FS1NveU4ibJA0DkQvuFogT7G+wgEF9kQuKwd41RT2DaIT
b+NKsizbyfzqbGUO1R79WfcXRftjOcigER1TL7ls75R9135vpqfgxolHkQJO
g3iRvGcbYFhrJr6wgbBDlxEpxf4lzMFxwrgki1/gl6zclcZIYvoA3qanYmbZ
SECAgnybRRK+u7Sjjoq29jQ/3wSdTUjyH6I01z04cVai3DMd7yIugLH+h9Uv
7MTgYIakWV2GlJpetpZfyUe4IMp5XeFJsWhvpCW0A5YDUcOJiaftpHTMMfxI
b4oUcVK9N0yKKdR+1rtZvzVdHNBKV/bvOmGIUsk0ucJc+jY9rEm1fD4zzOGE
hVdkjo9QKHvOxUVwn/ZvNrimCUlrrjSqwAAd3So4uNxnXav/3ehlbcRtbXwf
Vz+ePSVXIBQGGc5kN+WLWwLAw80Q7NtObFoq3uzRFP3ekw2e+xAwEg2bDMSq
cr5Hl/huK5xrfgkUMY1iJZ4Ig27vuwqHSEb2/ZPjA0UBS/yZ+cA+w+430Hkk
MwctkluIc7lM+KTNrkbPDFgnud7CcBMRtse6wvFf7hA+DdxR63nF7W6yh7F8
1XCnQ7cWbMWz4BpFzODN/r8HUGtC4JXIKckZdh2Qs4xc/2hHqtVmzEpehgia
Q0casobXWgUO/qJkmvb+WyEFE6DzLw93MzYxLB23oMmo4bxq85gZc5KqPbMY
/iEKz9T7fLjparuzGGgCUFj0t5XNaIpnGwAM9EmbX2UoNNXuTyz0Vg810x5f
ySjHvaquBE8YcrFaYCYLwSsg1pQ77IMz02TFQuxoGjGuOwUp+o8zr89vY9XT
l4Wo9PAKWH2fZHw3y1Sygmq3ZoDIZc82tq2dCmNUdC4t+j3ZjVi5MtQq9J0M
ktNnM8Ft7E2WvUr+k83or2rbIpRlygqmGJy+ltXJLkYAaYwx+4Gn9Os3yLmX
FTHw7OkI4+74AitgYtZkN0Az/5qRuY/IT2Yd7O8tDGqoYAedUfWi/vsQX+Bf
sW4m6mS/zTJijtRQ6AIqmHvlFRSz2ndPwJC9IFvYiLhmwR0S1pOCkIMyjT6w
Mmk6KY5PDbKHFSkgkhZ217MKluwJdrEO0MsAouEeTl4qdiOjekiDYyefyPAu
rVH7TY0iPdywLun/YE3jwTEc4UOVl28p8h2FoxBn0dbPd+LXkqN8PdCGu7gW
xob42++btBpptOZb3J/6zOMfUXmPqbzhpH69c6LuYMl3PoMO8GtOw8FpaF4u
Z+AYJxm2Sx8VXrOXmxwzGZ1lCefBVoT1m1R1JjHDUD7NRZ7B0ohXuq+jNj9Q
XJfpFrWMFY/GnE40LrGqDzZRDaZrRsEepf7yx3mR4FFE6FRRyN/FP3lM4ygL
GsYGMffRNa9Qe+1umVk2JtYCL+AfIzrf0RoLQMgq4JVRXypfX6/2dWJ0VLT2
RsgrjPwBr6eELiEh1RrHWlu2ukkUMXUbpfcpVWvzKTpDv9OjMOP68ZCxIUOb
DmToiLNT2545aJA8GIOcSyfGQbqFbzqAP34zuEEwf9/+JMwp8gRQEJRRdUjB
ommqP4m7A9ZmjZSy200kMfpQo29oJ/Yjm5zUtcGslPJ4i0Gv4LZScaEUyDVD
5blh8/PotO14FTbD7E7du6u+C4H9L0BIEj9jBp/jOhE+4ibu8GcJAerZ7c7o
1HkymAQU/+xMnr/1PCIVTgk6/c1Pw9u0lZ5y1qD+C3h5eveQvw00T47ZPnCg
hLs9jCXmjDJ8Xw1hWOUIPKEMHLPPeV0tfCAy8UbHSGNPgpmIHeFwVOeVWDX5
YZ4lkvPG5d873Mg4QltIlXB1teCfWMrq9wdz9w2FUltCBkMnIZMzgXoyuwFi
7p2TMrA3AerZHSZuIucQhoD2shdbhJbFCuCFQZ5j7BdDWCS/NDtntBii2jqs
o+/nt4DArN8yfF4RjfZxcEorMSZN7kexhp/7FOxGU66WRjsK8OQTNiJTIQXl
46ebiD0gk74crS/5eMhAdPPfTxOxMy5ARfgGjg9XPZtlsupZEDH+wdaJ/eKW
bUbVFZunzTcYV92MVqyHK3DhERUEXlNf/IOxh7/RIHre1XYe/zJCMIfNmnKy
nbEbzNR3fQJ/IZb9Ot9lWtMwzxBxPzwdyNF8oV8YW6xJy3ANmsOCBlJVhl91
vyoXuNu0M3/gOBBb7YH/5htmJynY+m4IJvubhsckruMsFmB5/EmHCD/pi+Rq
Qu2TDwVut9uA/9ujl5dEbEkRJVustHyXMGbLW9yuNEfAdu1LYoCZSVZQm2xW
+wPrf/warlxt0U56G4trd4vA6q2sEI5n4MemfScPIkaUl3iRemUAZSDhMLEJ
N9LOAWcA68rhlZ+o/CXreFke8+j8omCTaHtEd5wnBUL9fKaaGKIhrmqBbZ4D
GgRVPSGFuU5L71WIkbebNmx4fi3bsfUNiwtqU0UJ/fcLoQXjQxS2zpLt6/4l
a9+gLJTBwKQxwGEQeTi6FhvoUOtLxesGK3p1Sjv0xOMW83zOR0+O5BqkfxDC
R5xJweQzHam9Bca/QxKouORrKLXTsz+kHh19EWVxGFdh44k9Pyj5OuKXMLdr
0mlR9S5prhrYEcG82+XO27URyn6u9SSljWBjfbBt3BOBsznf4n26jz2eusC/
uiMgOyaGxxqfQQyBKSGzqsMpn5q9uNi8zvofW/T6G4cG+c1tAhvbQQ/9NcUy
mu3ewrF7hsi8CW0e2Sh23Qc5MzQC3IParYrOG6YC7CgLwAvYFfmNuz2FOJj9
zGCMMZ1ve5o9g1O8ysj6xaHAhExkJBJervjPCJ+6+fKQy2rct4WBtWo5NKI4
W+QYWyMMFvYqfmd97ppqUFnV5opW70AopxBkeu9Fv9Wt02f3IvJbP9Wdmvj5
vtcOSZm4OJ5aOJWvoO/N+RYKZiNCNhM6R3Z+hIgdPyTWkRiJYNi8fiot75ww
7xONk+y9z907jA+Ym4pxdDIobQO/S8QPcjF6PAFEXQqsr8kc+FDkZJMIFeSq
36yw0Vx8rRK6GmyrNPLRXPdgK0jdxOGIfGE2JhYXEQJ5sKT0ySbTWq7tqSsA
tn6+WrCqV86sAczq2b4PlmLLxTOWCkFtQaElipsoRCfrdycs8TU9d75Ab/Nv
1UUblm4TSLt8iJCFAiLPbBrcuqsH0QRG63oZ/WimYY93A/PdT8dfCr0gmrB9
1JYtU+pHRKd1PihBJtvEeOA4adqDqFWYOrMQCvfS+JpXKJX5ZVlS2HeMNc3+
z0TRAJcw1ACgLO65JEtwLkUBBm5V16K/uhkz78eFgXEu1HpyH0wuW/fZ7jOk
YjT19u0MPMeVvh2aUvURyGbxbpx330j2MahKKmI3KonsSY5RbOJ+6S/SJaO1
icLXH7eIYLUflpemqlQ08NBI6B4sLrwZA7eqh7iWqhC3WWggMiMAKnMe8orV
h+s5wWae4upOpk6TGHs+lhI7Ts6l0VHdMHL01SqnSaLNJFL43zTzusd8Q2bl
5r595kzBTEoF793OA6hgy4QVFF02yU5cYauMmgmaKqecfjKi4vOj4Yq19cbz
zY+2e/HxUT9vMcRiOtDoXmT+i7QgsujVHKW17iKt7eCa5tTapfSeIise1821
n/mQINqX71uG6tb+NjbXkFLlaKFQ8CE/+UP/XynA6jUuLsrEtdzapkOFeL/O
kHmWP76Nf/j2dPQ8akrnXorb0h/NKclgRY4xttxe5CXi0A63d2f5z9j9xwBC
UQpG/xXAVlj91CRWuuJIqR69RlzPbBKH+z/mlJdGbi/LrXzILoiUtXafi3cL
u/1pmbiFr+28q3HcExc0qoX+IYIe5GTguB+RO2A/May/hFaaRbjufMMKDdur
WTp3/ZN7pU+Lu/2Ev845AzWUxah21le2Qpx/jFEg53ZS9UKJwrA8rteGh4/Z
K/qn57iVn0b++RTjpJSw6uGADG8s8Pj82xFi/FJN8DxbPQaHSMPbn4jWGR5m
3HhiH6UfRCrIMxIjvxZk2J9yzd8BQ0P1BBxFonTaUI6lk796uyJGkWh1N7PN
Dah3pOQ9eh7C5cFSOERy2x7GpxsvR5bwIPRCsmUyck6zVB0c53wdgCQalSxQ
eD7Igom0qaqFu7TfH3A/Ui0IenzIMCneDosEdCVdQfxKAwiaZDK+2pNOFKDj
nr7rRWJrRTHsvHcTzqxh7JBjku2XiWh5fWot/NBgtO0fq0QWWzurA2xrCKm+
o0YiMkDV4vm0NueVJdl7xXqiT+gbKhXhh9NeZyfj8Cl//Ks49b3sWs5X5vgt
3x82bQMmVzxhBmJBLNkkNwdSUfo/h04aI3OClJ+JVCZ2RhiZ+oAmhkcM7b9s
8Saui6HeUL7HNk7c0l8I5e5sXnKRsrUMECW5hbDCzfxN7/kjhXAIdkMe4Ntv
7HQHITbZvKvoHJQ8C46zWVEMyznJVqlGwUJHY7hXsHEKeJ37hOYk3NQYihL8
xJqNW0+o0fio42whv0HqdcrwVrHm8f/ssdRD5bdxxz7dBKYcBC0fqoLVVYK9
BMoHzYyHlK5Ec4vCkNiuu/5EkG+FSIeyhJcZkn0d4WQ1zW5Btm4XBklhsBk1
zumDlqD2GjPB5o1Q95/DLas98xe2phrcfxcuEZ/waFCC7XqqHOlKo/JsbGxg
pCIQmK9h1m2ojkur5iU5Y13/3fZDsuW8nSieopVFEG/2FxB2NsD+ZYOFUZC5
iVGC4ee5ck2+inmiyU6Y68P3rvrnLB8ufD9k/elLRLJH0nfGmzhu9ImRZCyO
rSfJz4uCoxlfPiuwUcVaKUD2TZNETgLCo0Um+2KHujGrtXZMF+FVjPVu9nh5
AJLpU4O7hEZWH8mWPajRVYbAPRl6+A32tMDvDaL9p/47XW/48gGiUXs9Ez7v
wuDAFOqV1VeQd9B+Jj3cQL9frCfhUoDGPJnj43c2aPY4u6rwCXUCFkvtc+A/
UwW/8Q5FPaWdD6XdC2EvVZKQEkjP/kevFP5tx2RRWbMSsy8aED1tLR/hkZrV
0rvbl+sIgR8NOSjyT4jtbdgSti3WcNGhv5mt7SXoKkJ5Wyw6Ay9IHlwrire+
zUZ2f7jP+pkzeZq30+i8Ss9RYSoZZthmuWP4s32UFueLoF+bKI3EhVxflg7Q
W7qC++IJUo3cmCukkPuIAslSWGecE4MkbBfUF9O1nUX07OJTkOa5XhOXyKql
gzmr6hvIrL4S7lYYbR4Y2OXL8uACcvb0Ecpt9L9SD4h+goHHURoilYeDxyDD
hGwvALksX3S9UbDA4tQyqWaktjiFBWm6fpPX3P+bIHUYc+lEgGWLb+Kgf1A6
uo+ln2CcFiKp3VO3aNK4ZlqZacEaiLgPowBf9CWUIVKNTAvRFeA0/ltl9Ivr
Rx7jH4LoPoHKq+joQCjdQmGVmxr/y9hUOQtya/OQULoqJrC/HUIuZ0xUZ+7E
1jdpR1LUiNYDDi9BRWRyLFn2LUCOWu0Eo/cRI608o4ZvUgSHXs+CN29Fgrzg
jE+Wl6DJr2ONb8EDgyLszKR/LupShAkhAYwL9Y8r9CWUOL6i661W2AvoiRu+
uWPvW0ryMif6GmhitUNcx8KEJ13Mk1bvcRAThsD84oK+kWo+H0tF354SREW/
TnUGCqppikkyU3/0Z9/gWTrmDkOuDTAXEKxENgkWsVt6YaqVPa7OpZChUwbk
G6RJuwdqz9FxYh/8iWj8tDW3itwuXyUk4wdCj25yi3NCHQ8eOrhKWexrtwsx
UrBv9GSuMnc2IuCEGwdI93bt0WmgkAlPHQFTcAATIw5epRjCb9zs+He9XUJb
gw9Loy8Px+Wu0uFjBmxzhnKKHJLX1Sd4DUAB67qemavMTNV+iHbRcTxN6aZz
ecFRqRsvj/24aDpsQRgg/HaUxzIhApsydCd8E1eU4Y/LFAjLVxymPL6zYgQc
61QBZFZUP0+ehIKLPidsSw/j9TdptNPN4c4E/Om89Og++lP5PLuqj+7raDA0
K0Fu583eYySdrkv1nTUxeS3er4l7PSjG6kKAy4DyJ4Pj+po7Jxi6ssYL7w8H
ALs5g7hNlKDyynKeN6DNONpKmA2YgxM/QN/0poX8e4d3flU09WqSKVhGebsd
ZHCnRFy3V+JOZAScqqNk/6rZ74eEGWbRoY90q80BfQG6HDWFqFQOg+kmkI4w
Mg2V+7JE7KNvGJnvm9Ni7xhfYgMCxzf/ARnnU6DEMWwurMh9vw4cn7bxKwN7
DdS0+QVMXrzyI8XoSmnKoxO/RdYkKm6hqb+2MYdeHyfxB0zCb4Cup1WrQTll
/gWxa/WBjFVxosLSNshtkuJQUPm1TUyMdFIA1TgW37wPxS+VY+DDnGeg98Yz
UrOa79Nt74C3hsVTKnOCPJNEQCGWN1+ohfglph5H7+K1kVcsISl9JaSPfdD/
vhaNi8c3f4/1R0KjDlQMi5l74whKMi1/ExFQ6zIxCO4L14IoE5TtzCU9vzJf
05AnsYIQC4aH4pNG80SyxKTRhn78OLf062HcdnYYRamotvszXFgi6IZSFX96
tNt7CtMjcTaYKBzkouNNsRdvjgGtAIOTlYqCDjt8X14C0n5iuNriNmB1ws8T
YA88mO9za6fnRSTEZnwcImyUvZhF2/P5iCC2QMRsyQ4JoDT4XG2l8d12ZvGK
HulcZcqF/6HRG8whSvD7uW9Zfp4e/j8mfcJ+m66cPaQ+1gBOxflewZCMhTWD
Tu5yT45ZC1zCmRZlGa7yURnlxpee/NGXMC2Vel3Sc6YFjdV7RSL0aPox47fW
G0j6K6hUq8jqy/sVP/Vrm4tEXWIX8I0YNht7IzqlR5XV8jQd+wPwh5PNzRUl
R0cvf8l15ria+LSE++0ESiLBFHotJug9qhBwz9m8r8ScPKRnaniRL6BIdkFQ
DPBpuAAPGJaVBt5wNE5LnnUvbhRpGiG20Yg2QU6Ds2bQ+cnRafsKsS11leIo
PSYaHW0BwJweb/n+X6JCJUrbVydXPFcU8leDUqHYqTPHq+eFSNF/bnuISajl
AMocpmuuilQW+Ggel029j15LMwhCBGDHYZv6NtydzYfs895EJa0z9zitbU3z
a1DpKnREuBhcoYOweIXqsYYT0kjbiEWKvEAZtG5WrBFMxTflZd/bQOzfXsRo
VpMmqbv4wrcy981HyrcDsl+eCMVITeW9PGH8pV6zLDqTRzXLVV0utfICq7q0
evWRyzQXgw5hCP+9VEYB/QI0WTL4wqdgjlW3h9l7T0hwRocWvMCzfWLPzrrM
KG66Pg/cPLb7qx4yzBlmME44evjDs/IGgs63T9Et20Tz06nBPzXE1LIVlP/D
Yfa6ATZ0OJUEdOpvRxXji6w0bspDhXjbRQvLCF7WXGb3ejZtZbbs8XbtaMfd
w3B7J2iRCx0//kZlKpJmz2QorxOalDU8Jj3cRsmsuSqveGvdz/pL9iumJ5tf
WbO/5l1IiieLuXfoLraHysL54dWUW52jiiuh5yFUuEynjVecgNOJ6J/hHlKi
Bw0mclkxnMuvGpi4XxcdeIpbXCYyhW9l3G6iK0zQWPRFkTSRcxkV/QW/4xin
UUFzay82gJWAwgvMMghLaACn2fy8+PZh7vv8bYHteek7RQ717gZsEFyGo0Y4
G9m6sjd/u+nRysC58yWblmFoF59HlRlGJmJjg8EpINAyYQaQOcwitL9O7ZWm
H1VbhiboH5T28elDAGpGY8uKPw/8fnKW+aUu1mVlUJ2uYRbcjBWBelyvm7YL
z0y3OkEszduT6DiVKmhjA4cZdzuEJZqbIkFmY+9lK+P5peVCXhQo5IuuOrbn
e05Q1WwIIc6DCC3vu+koxNcfcnf23GtkbgNHpss4/putPhzT9vq4k97wzDtG
hbhJe0wM/RBM0h8x2+asHYpqOGsRJNwqcidJCLtI2+YzSzouxs+b3N0DBbhk
5Yf3ktsvTV8iIzsTbJrLrYhgBKlc6j+VHzz8msIBYRU1vuQDMSNXFzTdlu5I
aRbAqW8lc+LzwzFwJWDYaCMTMNU5imeeYOGglsOU+32VjaQDWXR9/66djnlI
eBiT3xEGNMFzPGPU1GkWdkIGHzEIbhvIu/aZT0fSrdy4D5CgLgPRvJu2Lqkw
gG/qpO1o3eBurRay/6SF66bGiTjzgB1LWk6GQUES5WgEelEgICzBSxg2FB/0
/kv/CkP33VMr5bN/YojvfwhYjtmyK3kvxLgP++IexPXRq2CUwHIIwWaeDGx9
8NU41ccNTvNK/YAPRFJKq9BVnfEiqjry2pvQglGHFLglFlhcvmazSc2XL5Tz
/lXb08Z07mUUmCAv6c9ULhtUqganCXqSyWzmFB6NUY0I82yQspzNC0iQniSX
mJ8hE313rBtHEbevc5pWQIIRxJqtleJYh9M1IGEg84q+OUUoluou7GNB7OeF
/zExXrv68GHvpD2YnjWNNzcTr2M1J1YY4aQid5KxWY0N/eA2IBlfxoIFcmZX
YfIau42eGto5EHYK0B+Tf/deuREw2i4ZGAkXWF3Tj9DXGjoDP852uGdLis+U
jW6+OKnhMwGxybfQ2KkloODZNvZCN6xXfyI7+HD+qDF2SPDO4bLMMfL/w1hs
irvADSQCkb1ZZ3eaaI05WHwfydDxK/9+p6/TvFbs0m5qExe1vxQZUK/jZViB
Cz0U/wDwyyd4UeYkTj5O3HCEpfOAOVucdMip24x4CxIzt16fR7wlDgXN2OFq
/nqDQJNnkdt11PehELNL7+bw5uD9Q065ody14yvE7pgMSHtVyTjv3KU49EaT
JJNBZyZrHJ7l7DC4qZuXFTtBjeylaqJm8Qew7wMB4g51l06OrOe+gby9b+ry
GiBgVOju14gHJeh2TSlaFsiWi6lhrmVziPNQehseqQK3jovZZRJtiATtCtgI
2I2N7lih6+1bGT1xASc7fVBNl1gb6x5BGor2ctPr1HAvu/jotOE/5YLFHhKY
vnTL4sPldkfSwKXHL5YWd5SfdCjvWbpzK/VDSQZKbx3bH8Mjji9RsNBPXdvM
mi9X8is8j02R7sNDT31FcABnYkygL+TKLuIysAdOuFn0QHtAMjzWdpBwyouN
0Y7uH92mherU992fvxrTMesJ/KO1s2gWnRx6l1E4rV2WubxKVsbW8t430Ktu
CbzXRGowvUAeW12atwNVYlEorB8sKkT2g8yAbjQ91DSMKDVnqLMvfnzNOlXM
nb3YjiQ4eTtx8CLN5ybjWYzQRRi0CERv+okTgYL/Tfgc+sFFLG1jf1uhlqAa
JdSIYRpdFh5JLrayjCzE6DjRpsGS5skhLGCrHVLST+0GfFUn37VFcvRDf3QH
7NMUg8pWnmx2xyw27hZM4UOtFDbSnMzhVYHirPnhsFrMSRdAyMCCkLZF7iPU
dkA3zD6IcWar9r972rsfOG+e1Kpfj5DhQ5zy5V4GbKuYP72KGid9fSk60p+N
2mSPEiOVx1zm6hx1zNCkRIc5gY/Ul0agbjXmNODv5CG+fMvCxk5daWgEd1sF
nD2akTQfKRhU2YzpIIn1NBqJ8ui78x5OoyPnCUlfVhp1udTRd4NDIdBOwMMI
bqW2NCygTVKzIPOKjSAY1BdSK3KpO0Lz1eLrZFBKMFD/kmhpYNkUBWj1BVOt
68obAB0HSpGQw/tnMXEFDvnR5vJh7cQNbeO6cvAmnV/rZwGBgPq/V7sJkF3V
8ytkYAHHDZVbTDVumb/IPc9KSYjwe/z2X9OpJXifYm2EjLHxps8g+xMLMJLx
om+YKJtDWXrHy7uzYhG7aAGxxtO716DXE+7kzgOWU/HlKJUUMZmmv9CxpYmE
WprhMf6MTGrsrjezGMQPmiYis3ldsgsHB5Ovg/A2Wc2w27UMGKNLFHQHehNP
ds51OqH9OfnNxLolNu6DZy+Ws1EGcMyGC3fBesJzpQlnYv1xfab0XJI9fcli
ICj3aIqaejaKiq9j1uYo9EqfsY5MgFlWAXOWpvmDXsj1dcE+n5/4jAeIp1oP
+ad4vbKLhmqpunUgNrc6yZAn9lM/rk6POtjFzGoxzKSyzDM4PUPq8/bvUKFq
5pA4eg6JKUUHGisSkGI6RCO81/H6XfWhnF18cAgamBxpZUt77hGIe45fXDYo
040JXuVg5XfrElzFRzefQauS6r3n2KIOA9QaJ9fTRY6Qf13z2WM/y0vgyRvK
lppQ2Nqi3gFUpztL2XBXYVXy3dqHmTWHJq21CHbCM2/Rkz9yDF+RsIlp3dbJ
FA2mTqdBZo5QjCA7Gqgo/DP29WON1+WXze6l5g5a4DHg0W+BeqChgV07Xzj3
Rcq/gSA7CxKJ2UFnLiGZSXtREv9o/2qp7SO6Sj/f46ZnxgS7bvef47n5Eeyq
1xe96BRCPoG5a8x2+8tBImxF2gwxBs6iO6s/9d7LoFnp1C3ROH6eto1CZif5
Vf9yYlEv9RPgfKSZH3DkpgjEOL7EaAAG0WU6rNhymrO7zsUsIp6zGbNF9N57
Il7+5bNENW2q0ltKGk9mcjZVsxjVqXPtV2mYhhp9ImCZhnGJqxvK+rSMlA5D
Ty/MsF+5HuvJD0028Goox6Xj5ECBvPRCkmhel864cE+99lMljGrG5+nZZGij
UL5a5o6wHv7FV8b3LulC8NmC+xcfFgUogw2xQcoNQyk0ZbC6E2SKTwCEHl9H
NjTOgVeEyND5HNjIjsvYODsUbni8sK6Ne65NjCxVwqjQj9VJiiGfggosxOUU
Xb76rqk/nhksgwGubtkCpsRvU9Vmdt+ZtUcm4I0SnLX270U0bjiZvIGJF6dW
8XFwUNn8aFiiiQNYNqXX6z3z30AXiq2vxCaTdoGRq8vwp/1LlW2wm9j0XXit
YzYPF5nrMFeVAkvyKYrMdt1Vp0J5n2w0RLQMVlqAhlBiFZo+/HgHNs0L1ESj
LCg1tw83lNZqFPbnW6QQ0vRlDcY9S2m8L/JYiycuI/vVwQ4eIDTSdKfySwJz
0r0C7JfDRf88d7EDa+ldQMW6HXtSwoejwEwbnCRTDQvF33lOxVIro7RYYoyH
anYAG4JZLXU6C4hsoPcJ1zcUVZ26cXXHViIpIBE5HwrOMKW9LoRTTbXuk3IK
KmgDNoTOHGvMkhJuqJ6VqbJTLRZCI86OYrXMT5JhYS8UJVJyIAXxJmAqY/jx
KXvp1MlKiLtlwTwFMrV/mHt4lqMcWIAr/ptmRkY+/yUy4JKrmleAeyDGRcKD
dx8BNV5WYx+791FCYBJf6Z8Ujwe+qS+tLR+B4ZX90alOO4J3Yh/fuL7fPFW5
cCEe6QL8AzcMUFxLljf9mmRi+/o+hFoV2L0Dm2EjNek2XGqAJozx2pcnDrR/
73da4ispS8dLvo3zGmOwyaBImtZHHDu5RhtQXX2dEWUB3F5ob9UwTfDcBt4k
ikZR2rEWMgVfgiKxobAP/R549iR2cJScvGOADflAr50s0+lyJbTavn5MqfOT
kPAF6zFytg4udnbt4diZ5HpgVDH/bAdVZ/8z5xyPp97zrUuMqZsC1mi8XzHw
bmNbUOohna9kVame53A3WDkSR1vnF0CM4tTdifzTPXyj8fJtGRcRsCvYTfVR
Rz0pD7IxOkUvjrAhS2DLtJmcR8rl/YLrOPRo8nDXr7Q5X1jNqsml4fzKAybg
dKmxshtoORtYdBbOPpKaPusXzrZnt5E6I6E3WSDQkQKjegZM2dWNp5ujmdz+
t04zLPpUG4qTY6yOQDJopdsm2gVZ9pKEpTT4V8ZZqh4SQ6QeMUeptQoJgSt4
Ze8Gvku2bHY6blrqvTSKQuEUBciyWe7+NpnPHoO0F317mAOf7kItbMNy9vww
NRNSlmMpOmexJ3hxyd3+3MQnz7TLB1S6iA/n8+iuTsCGzTJ8biCdq7fhI9za
1gQ/YDs8hZYGZqL5FwCWPnuuyas0LzSg4ZeDHI+bt6iprAiLv5gEjpv1LoFE
kB8ArW6DXOkQ1Sg431HAKuSnFANMT1Slo0jMOPnp6s/Bc+2T8rq0igEsZFHu
1T5cse4O17PQv6Mqpizzfiuy5TEWrUSWskar5hhlk34qfkhfH9O8R3/Pbsx0
iTyIg9Ars39rbPE40w4kPStQmptOmrlyCiQDbMTJrkYm4mDAKmAbgeZ6r69S
fVTI01ie+8CHGxLAVgtxJ9jhD1ktqiIefFu/nJXuCqV7PZKO9OpfIuaagQCe
IKbgmLAuX0d6qHTr3osgxkzRgYsNk4m7epI8rrLyGAAsw96j0dLtcfa+3lGb
b3iN2/veZtxAOHbgps1m7A5BpVbMU6qG32Bs/xfF9DF0CFjZslmg4L6HqhJE
apTtIJYp0Z8RNKqANv4IUNnrc7n6/M83yOrLan70jFkfgQBaabTl/YwQvufE
Qg+xp9Qlslz5J779GU1D4FTzT9K4+RWlusou1RvNYWNkVUlQIfhmE+s9IKeA
YDef+AeMqGwLnP6KBh4wLuIaOaXckVhzfmWjE2ysjCgba3nvXetPqknzxefT
9RGeSJcwxZdxHThWrjllvq5igaI84QDhEYnsISVOTKqi4jm1hbyCk0wuuFiT
9HPCb98rtrWGZhjo6NxLmqeBr28Py0QxGLBGbGQgc1HuKG0F0XlFTngCRz+f
2mP0JmvucsvbOahNODZb5kx86nmhKlMi4pDTnLNKx6p01QZuUFUSZlSTDGgb
8ILY+cdYl9tbmrgsrh1l3k7kSpXie+Yj6BiuIT+WwySr5mqTMe/6rCsP7NjR
wT+DR0t/bj69ONMEtJg7lNB1XgjQd/eMptR0OM5xrmL+BNCq102pcseAGYrp
t+gAKJms9LkM2G7m1j7SZ67e1bZX4GrDaiPOo8wS0rNxEAYxmBSTWG30zuho
d3rwCLIcvY9rT5sjM/d7nUqwjH5SlOGy13nU2MjSTMdMR0+Y5D837sCbpr4f
0/FjrUPGGKQgUapI7ZV38w9A9Z9Rc5qJ9RS4e5jQkMYcnCvdv3NH1D250dRw
uvxryvmRZ31huw4D1sVY5kI+10FkEGu0QszB5YqpMV9bBP6Zh3qODKwOQqhO
aArRJbAlDUAweSUJo3rIn2OdC+Ggk+3HHFsSJ9nX6gzrK4bkloPFyRSisleB
MPvkJXOzGipUG7X7pKDfCl+nq/kSPQns182Pl0glnztttf0RG9PxAyUmPuUv
ZyuV++qfUmDIti4NBNY5dLP2FRrgN+Bm7JAHwkPgOiYJYKNadvhYXc2OOQF1
YZmKd5tums1x709ai5VSbmYzFgmo3XlanoFeCb1uDM1pWRSTVrjusByEnlsi
tR6JU2yJOGwkdw2ioR5m0AgcQ1cZ2FHSZQw2RAYaoUoFmyT+KhpXBeJ5yiuc
Q/lVBha/ik2cGvD3fdA/MCyPO0EZl4SUAIf4HtkG/949ZIW3YHYn7Eqww9pE
RcGTOZvG/0zjvi6bqwEEVs3Uf03RwPc9H4f4BbC0aBgNzgcF8tG9mzDSO6F9
VCqBBi860aa1v4oxlw6Jc8XigmYyKAcAhAV8oZr4BHtO1FAQagt4sUMphiKT
rLlQXJEJX4R68U6Xl5hZ1ezrEXBtXKclAJeHE7473omzLWzc8O45h95QmLQ+
r0/QqGgvTTl5q19ShJY1muMmy4Ua0Pf+2w8y5cO4meFooLFO42zrvOzt59e9
FJNN/hOAKLXRWrmLarK8XRJNvKRxKYeU0S7eJKI5aK4z8efG5betsMVRNyGc
gEH2yg3l4HXBHnlty6LvH1P2h5aEXt5/y4Quf3Gg2clpIatCb93vFA0HQg70
e9Lf2SVfPNwke52M1G9nwmIBKIGrxlHzkqiGKiyDYQ5uQfe/vkY2efW2PeNr
M4tS91TEShCYfYmODWJOIad5Hx/eZR11VZleeTvmfChVvlSehrzkpTzvk1Fk
SfVcmUKawDVtZ/5Ysc8jfKjWQ25RY/7chjwgxEQ88+E9klZvjFX6rU/oc+nL
fcAIJF/Xn3lc0lxBWlCdTRcxu3MiH6o4JI3jejZEnlYcvvPaDOIHz1l6XYTl
ftmwDBbIk0hmSlH8PIIUd8tZDOeh8Z7vOhp3kLYUIff4D2VU1hpCL4KGj01V
Mpk899XPYkTbmdQ5LRu21e8tDtAl+YDySGvXZYKrIT+RAMQEulOF+uifd1iz
ReNCve0qdqVYwub2DcdPB3mPR7Wken5IO+LmK9XwxVpf9s3ckp1IJQIxhr1q
y3vq/42dl1x4I28uX2gbegNSgsytzybyA8zBSLwECl3REoVN+ZmT4F+u/weS
QchjJz47STEWTnjb2g7cfLxmUwoQcAa6BJNI620yyULoOBSykZPAIUiBwK4R
5WBMSA636AxsygLTMjQ9KU+DLtCZyaZ8TMo2o1bEbn4W9NiDkZKw43+YuPuQ
heKebKloEn6ZhlLZA5o9qG/Q4iVzdAvIjVAG57R38GmELTzfU9loCePOljZU
fdX0xGkdGHhyvfrgURX6LlKx+ZplqYhhw6b2BMNwYne7BpoCYOwYRayA0KEe
EzxRLgQg/YV94aumk1ltxNN2ru97MB5HB1Px8K3qISFxeKEy4DvULxFTaeWF
6ulx0uERyGdjekHbO/5I+hFAi0nhFd2BXBupPY9zhJcAqaX94Ozd570ofadb
niXyphSlbStPcktqyo03UoS3jS3iXLlKncT0wsrWNad4fePAWuy1Vh5saC9X
YEPmbWf+NfwhM4Ht8HG+s9pdhqfyMCMuXPhHke3s0uUEVpbMbfShqKD0U+Ll
HsVgnUGWB4E1kp3su/Tcz4n00bvNVqMKMx5hPoIK2dzeWEB16KoGSppszndd
HeXXnBXHx7uHrMZ49MyGdMOyQ2kpK/UcDbjqeNxMhH1Z/2yu+jgu0AMQfsrE
8HPq2s7zgQ9czWhRN85rFGz1MFwkwJs046g0QmZ/tsXdScue0laqPZFGpxZP
+WbIdSWV/xB538oQoktJxOsI9G3E6P8D9Fv2dGO1uhn8+bZXAbIL1D5DgCHR
XnBDFTdSq/GAjs2vq51YZVj9CnLY5loqCg3BTtDlTQV1PU3ltPVUqftiIA7t
WdLjaXuNxHqYm2HtQlLicjRcoin8FXmHyCUEx8RgJZrQZzfZOASPR68GUCqt
CKvpVE17tQ8RF+kTnfUoMMXbsjNHWw9eJigcbcK+j7j3zv+Je8Pwp+pS19sL
LyJX6K+crgrboXRvN7OY4AjhpAjnyVJd+D70rYgzmk8Y04T/dODQGF6cC5Nm
3YWlXEtQgxe4m7dZX+tkvaZBBA8Paatn+Z0mn0osQ3VNtTDeoaYStUGcgr5e
RVhG43D8iWhbzOigesqHovvirg711UQEWWj4iMAyi8mm9UrvS24F8ZHNUlZ4
5TYHmyBBQDXJiMy5L6lBUaD4O7gO4jbneccEvUmzlcy3/fhxyFOcub18KTit
ZTDQVtEgSz05dY5r5tzw7XnQt2PTY8m984g4JyBxEFI5iD0hNfWJMorKchrB
qMoRuOkISw+LDGul4pTe8LncGJP6n2a6Exv+p52wfmsX8osaLtjfIhfisYG7
aHfCqYztXh6ASqPPyrNnzADPSJ2Gl8VPKvbVXjU8aWFUz1wNAz6C7a55NAb2
AffCX5guGeAL80hF7VhlvA4u0ho5IeeVqQT3NXwCtlY3FemOnnQShypZ60U6
NhYWDM+umvrOtJQhOKlvO9WktdszHnQXMlpeP2OQ+NtfkKocb6PcqhjGofUy
PNqXHzrlHtHyeprT1dkRtP0xLLaxrQI/+alKuPqAZVKCocW5GEMZhVzh+3z0
ZF0IeuTImkyj4UYhrRTlOrlCU7jneaUXSFXmFJVz/rY2XRvwMhU+LrlPjKVJ
ifJTJ5z2aY67k6qXLSeqa6iEczngpoVQCk61iLGlU63kXKLfyZPJOFOPY9w2
26xdk87urL7/z2wnhvVbDIsrtFWHd1RX7prLDB9THZDQlmfwWVJi5QZ3ouJa
ukwbyH655GuqF84hZZwz0AV4uFdUkyB3hoU0DdmhunWWMv/+FF/6MDCq1g3j
pky85hYrBDR4+Unj+Zi3KO++yLMcDz/9pNVkF+lleYKPsIptMVLWTiZ5axPC
brC3wh0KvRw1inEu+iCo9NjJeY9H1mMWCPAcXmKsOzaijFhtdA5VuXcyMbL2
EGHXqK/VXsjTknkkp/TWBhTdRW2SuuUhLlZFNXpBnHuMAt3baK3C78OGsPXc
F3or/rQX+BU9cIxVhW7jOQgItQlYLw5B66R+ySWUxhdcyFFRf3tlDxZtjckB
y3nUvyYKUK5g5pTJebhYumsEnCgjJvNj5zeheIMv7IRuEXy1DNOe0ENwclnD
Z66WlkpEDn7atHM1Lr6ELsV6QwL+Zs8I9Ox8icS4ZkjpxMQ+yjHyH4BOogRk
IZQeEsMzcj6CNRf7xkqm9p6Ojn45O8cRblxj7bq7qyJdDI1IfnZCe/EVEIMI
g2CAtgTO91PbbBAWhsJVZuF8jPBLlou6Rc7Pc9ngTjc6FhB4/f49PH37E4tI
XTa2NPjeTxnWyizAKGFyX3Wb1KLvwoyXrNyTTuUesGjyThGEDzINSihmLjec
JvEMKtb+b9d+2o3C0hoCB5Q4gmdgCV2lvcISAuPLi2YA9YTEVxbNl6K/bwi0
/AGKa580itNqI4C2gyBHhqRrtZloaQImgtBPDPk4PNc7JMR5zsjyrSeRBeH1
5//M/JfJkgf3MrU3qAFXe1O1i0k9bM1nPXZduqS0aDPKcIgw4MXOXGV5AStV
1+pVqhQWBaBXsZVDvCqKk01wcysEOIRlobWKRD3BHynZ3jBw3nRmwywwzMhf
XBKIgsuiNnpHZLhuIXOckCSGghPtA2BpSBbwsFcuhoqJDtHeAbvks92hVc6f
U9QJ3NxH5IhibWICmZcHi7/Av3l1uRVtOpk8Nr/od6fjqRjvWwGdFpmFVnhr
JUWRpvtDdJr98DydhsIKc2f2tzs8hWl51ywWsX2MOEAm/7W99aanGt9+N5AQ
qaIwG2ZgIbPMTRAAUZhrBqeN84ni+3TANZsUDPnZLIEoOnhvH6UE5SfdAdn0
ikZMCpsZ773jUC2lY3AnXzSAhBUoWm2qrMOj4OB4z4YXaQ5dneKlAhNWX6Ch
j9xB0kYZV74asnU5V3czXnCw0ySMFKOejEEoMaPqXBknh0NcR5lMOWfHdajz
XfGCM6hY5I/Ksm+D++M1nYQVszHjW6sl8TCbb06ENkqxHjILqkZ+JwqBRAg8
YembAG88BA26UIOaWgbIyBdQ6zx4xq6jW+/99FyU5s9wPsR6fF+QnGKx7+I7
AG3QLJZaUqwan4ZklKaaVbwDwkjF66PD/GPTlTgXidlfLQSSXKRtmk5Z3Lhk
7Bu1fV+eatvNP38kQhFqGA1N0lIqwkHaDfnSLHq2yoojXrF7I5OUN4YJqkn0
sLrMjYAPF0HiUcpLdAnfFexhfexUMMppOOOBn5gNGHS5U1jSabWRH+P6PW7c
XyL7k729tQL/5kxAjCGjoceACH8qWZe7zg6AsWH0dZIfDcsB4Mh00PoxSvrf
4+If+1Od9diRIihJhrW5Jh5LLeOqMQzHwLfr7xJQoMZYHMK4BIY7fkg14mHY
+QGEw8cf7Td5/c/wsV00+OF+IqdRgMmpn7gi0vzUCJn/amwVizf1v+Hco0q7
j1A4wAf0/jXzgKmKMAYyS/W2tuCZ0ckvaO2XR2Sh4cauUgzzDpa1h52Hul05
x5+JGFF0lx4VNeFf9tFr8ao7QzpIG7WdFlBKCP2ffJuzGYt2BrvYxOFjIE7n
jRuUl6LFgba7b2/lrS1lB6QiLwVjN727kvaFK1cR1pB4EOOpg0IMvAGyawOR
/gNXg8rKBHhQC9kMe1wXcbBBfxV1rYM1sZvEpRvmMkg10treX50fNTM6yj1M
3U3zuW7suYYqoXzDrOZWlbSkwvH59OiC8p8XQX2cnkMvVhYeCJiQwl70kxJD
SLgcUSpLajSNjzqcomb/RXXaP/So3jLkUebrWs2JmA7ERsUEPsePS3TN4j/C
okk8LsaKMvJ4r3yXTbfRWummmp8fG5OknP7a9tXl7JLXZJjuzahE0Vsuwq0W
0hXJaA8qJgfOGIahClOEx4DL0AaCYeZUp8k2SWokQM0oMAPfhV3u+/RT8K1w
2188BcOYyH4vinc7rx8U4P/yw9ktEFf9SgCOWNbhGy0iS16CyPiytrkKd3HO
JnQM2Yi95U75wB1QKrZsE8PNKT8hwv0eMcEcN1VrAC/JLd3wkZwxKoVZcKKq
A1F/7ljkkUvkZFH6dtnhJ+Sp01AxPTVVaLqMWdRueUPWGwfgn8MeNBech4nH
Vle7DoZEVgmoJCv0sn2X1Z3oe/gbZQYW4RMczx2lN5tdCtASpA0+GvTXMRDb
QvAeas8zBxNcnK0aIYLatgqUiY3eM6IWnJr02DnVCRukQXgPHKre1leftovY
1kVNDFeVltRkGHekyCBvZGHVFpqnPcVPa0dixAaF8OsdYznGOb1chizZEKQK
kk2cDD8/O7mje2BDNehvv3amjeIemwAyQ/dG9Lz0ah8ZBMchHrqcsuLlYaJ2
ivO5M0lkKc3N98KE0X7bhTLyer5cWDbq609THUquEewC+OIPlQlk6Vy/Bl2e
TSwJRFDlNTyj85z5ppYZSs3bwIUdCtwGN1B8JnVYor/3GNeROSdt8RbbVfuj
4vp/xBjXdmbdMCw4k1J/c8xoXzIz4BAXLS0PGgv3Cgb/UGoIQdFQSYaDA7Xn
shQlOC9d0dP1bkTy8Z5tw9Lw8l/Nut8AJUT1exxg0mb9tZSYrVmFDu5rSYeE
7h3JGQq8fWSWKLnDUIBPvfgeQpXsnA1gQiqQ/j2HvnFDFGq7PyF/X+pM2I2K
aB9lJ9NsT7sXk5BnlbMhAfJlf+jvs+QjZ6FnbnU4pflbJxXzmOF0WE/0n1hq
utCVm0R5yGg0gTySsEhN94I3c8GwQ6jI5M39o13CVaRSIpU28+ydxKnxIqGe
9jZ8HoYvskoFBiiygayJoB6rbIJcXSzK5ceNf0BgEtUeiU1FjfxghyPXyLhW
rhJIabaH/PA3UsH4tBRXmxUNsju4XXIPY4i9l8slovA61JkZaPTuh1JqHXSb
gXfOTgzNAgs6rgYXhhcdk/EDIxTELqE08NVpPXwoDSemkZBOi6cSycQvy4mN
MrBAfLJq1snr6d5KGpeWXSsA8c6RmQX0/AiowD69SYoCWqMOGULl9tVwIfkc
L2BtiT+ZVICw6ow5JrrPF25d7Bpe0KUQCBHrhSFKaUymBz8RBngwYsf0lhpH
Qha5rc15ALe8fg2odhXFr+7HXag00luCq6jggWKOBX4ggK05gfp/5qURp1aj
9DJfgL5FYOTCyKwmz1gGzsskxfGr6jiyHFxj+UgMpXlZSqlyP4qUoznlVn+t
BfNdjhYBGy+d58oXDI4OlzXP6LCDke4JK0i/HEgM5w7Ih37FLQAHrxEFKu8V
H7Hm7c+tnfTxY3l9mHlLGLF36Fg4Tb1KyoA1HVUyeibGUvcsEJBJBVkVl00b
1PWW/K0sliQD8Za7VIEbwZJeupvxUU0+thZ2+mIJysGf6pcL+Qh56MLZMw4/
4vRR6mzkDHYYkJ5YVG3qhjnxgDCsPmdHJZEsJSPrWWaGHnGlusxAFsd3lXp0
bCPJAhRKyc4VeLXxMqsMgc8UC/JTKqNw3CmBbaew56BxG/g27jaL8v/cDHvb
EDvke3zCRJgjHMW8PFpLmqiQg8MZJ1LG5TsE/9RgkfoJ9SvOEU4CS0JFyArO
58nEW4jI0lB5ga7B+XJSNGbPCfc27YsLMIt1W8gk1GEtbfpeaAF1LGVfrthY
yE8CFlwVbCGSSqJl5nkJ96MqkiqfAda6j1wC2DmwleHLG/TWa/V/wAZn21DA
zgqYitpsyHHaVKrxUHhmtZz5SvpoT3oVBG3sUhG6MCGY8tbEgkGDrP8GehSD
WhEQvDTchV0EhT79mbrNP6zrii2yS6aaJfxWpCLN6F1rzRXCSyeriNhreAhE
9IVbLpCYpUWPwe/DIH1hM4lKmIcyGUupkLDmRoOXrOV394+yphGJrR8EyI8o
fLcdcF51HqY7x94WrllpCkUjTKf1+QAZus+rMzMVbSkif0rtYAR4qz/w7inH
owMFCfhL0wMY7OmXbhoNe7P2G9C2k1vYMAw0uSsChnABD0QKUWdClskMg/lX
XLBwtjfOT0skktviolV+/bwSLCBXeqOgy6lo87KEFQck1+nfPayUWXp9B/CM
yKccalapXoAop3mgPzDO77X9vysxR2N3+D57nn9EjwYe2hULNG+/i+gAIkXY
eBJRaQTP2xoyaFvaQsK0u88XwvCAOzFz+KbinUs3cUIb6rwy8a8monkWAGLe
qHvBQU9KNodTLSXxB+fciPKWTRkf9JfkSrk+e4HzioNEis9ZRqOaix4vPR8I
zeREHmp0hZpqTK0ypq1gc9PF71zL5iYpPZ2BTyvJO1968VBT6gvs9vf+Kdlr
cjkxNHUDbaaiNGLqvNEld+82RQNSIA9bH5mtkR/HK2tm2siQDRd3X7DVqnGp
GpYSmf7fMMtjhijjuAoAjq4bNybzGbpVlVTOw9zJhtB5BptYqCUkNbeGoLbx
UJzNnulhntx2ejMnPTsZ+eMhTegKXyFNA3TSGoufVrZg4eqcySqi/E2rWjCB
PIkuLIheguiWeSIXyEnuWh7BCO3JMjSIYUbJlmhfnxaibwFbnx34hQWg0Rbq
xf+N2AyMxPyy5mZmHJgvNnfAfRDzawHS1BAslHyxh2Fni+9vhMFyEWeHz8dH
zGO2CTDiQ/YeAYtCP3XeHLK6SyxuJYJPHdB3FlfNtr+8MkKuVsHFVRIsm0Sk
ZgqsGsO42GoHbJiq7VQUg/6201eVPw15hm0lb8s9KMN8pR09wCl5sHUb2YYJ
PgzvR/CPEEqu0M0rTzbqBinr4FlRTnadWYphgSV7Vx0YNN57gwaS1fPvuFZe
W5ucd3rcQqWHWC0i8fih/MEqGwW3lG2QzuWoV5NhpGpGVy1IZRp5MMCcXvLi
AkEB9izdYXmU29BV/Z8eNtyF1AUKYI0Vkr4v6RWshcEqio1b3tTjudn8Ekml
euxaNMYbodDbjtTgO0SV3cd4U6mYDDgZQNm928QhqU+4WMvdh0gHtqqyUtY5
dDPIB+SulgxZ4Hc4jA9eZf6LOMpPiChZJPsh3sbc41khdPVRFd3KcpYImzVC
iCVacSFQG1hffYI8k069AUEJgTw+5ZsEoDYZIwtbW5Jb4CgJ4EuWUxA+62Sn
snf38IeDe83oIQpyDBokSsepF/dEQ73K8LwsKEIeUyIDRH7rI36ydGQKUGue
Z/jRMpExY73lMiGNnxO2elboVJO2rqyX4OhLybF9JAACRFOPhKVBKum2/Siv
x42vST9NVeMPz92o3KjeIGCFf/tRX6m1yK3kTzHILFPb+Kawv2zP8ml2MSdF
j6GjnbNna6ZBNs2UJ3DpKQCzS7ZqfIfer82XaZqla5/t1yNwxDvlpNdCsA47
l/wlq+gLf3ZWDSCRcvw+NhKPWP0uqr4//imnFGaXsqUaiN09Cue4V0SMfJzt
3OktSdI7CZjmrIJT0PWxEzlWFiLzdFnMpQ5qLyLEt3Sy3NukesTjGEFby3ZB
oWkTWhgak93Y1j3SgghqJ4707O5I4ZUTE+6ea7OKrTE3kDiLo0j42flEk2sQ
LUZf23ISHF2vQveWpIBZ7ZABCWE5rR5cB3qGZZpHYknGMri8h9WNKFX5euco
JrPoqt8b9KvsOqdnPHLu+2i1ZIqZOZl2agkOyWrTO/vp4QeHftXgYy7eoIp+
inzO6d/3NdXN3NNWO+yAnnw71u4/uzW/bm339JxMCQQc0RGBZK2fVtuub19Q
WWofl4IZF3dMUSevSTTEuXEEKZQDNNZQiluw4MzfFww2Dza2/9+g7yIpW20S
RaRjMrkWoKfqtilQsYwUeJFAc8M+vIPEvR2MXC/qIp5i3DkrP283ARweA7ye
y004f0oO6HxOmI3SDHVNKyR8XD65EegGfjpYE7usl89drwLcxGK9F3Rf3uu5
HvH7SA4hV8A+jDJnjtcYUzOzTmRUqWmmE1q1evvKFeTcvvJpMAD1o3QWnmaL
5wKPG9sTAYCOmH6SNSucm7XDtuK0IB6HudNSKMO9sIyXxo9aOrsSSTuvro9H
n0Qxc4pwBngFXq+A/f22WC0PVvNICqVpsx+hqD0unpUbpKuWTkJAHbyLrirU
a8NnVJBbPtZxGTj6yCyrCX4YHgpaRPGEvRXKZ4gqGXsAPz0K2MTq01vO1S2t
v4YCosyRY4/ZEP63dEbHG0rUEZstjTbya5s4uurBMhZk9ch7Ya2btNTu1J9S
yiUl0MHH6pcdjyd57LtvXH+jiYnaDKKkYzlTU0RdT23hEeVhXHmDJuclFPa4
JJaVYCLZGsdfgO/JiLpyaTii1u7UAN7rsUhs2X9uSo9zIi9AQo71DCkEjomR
X8Gvq5DON2rw4CjYaeRdBa/SZvVLN19u10Fw+DiOe+nX/YMz18Qf4DSNhkdn
1hgc2Z21FcYTCuoYGJXOsvP+DZofxu2rtbALmQfWyMIWovS9f4BQCdg+iHlZ
ZkYrNsriwuWxwn1bdzaumlO+dRAQDGO3j9SQp5EBPv41h+a04unh4htgYpr7
+iUzy27VKoLpUP7zwulN2VkJ3hbCpaL7jQrPFjxYVX56PlG3b/QummJ5XCYd
ZqZPB1j19nrMWkl+1RQdm1ssS6n3rinHiekoj6PFq+M/H9frjOAD45YDgn3J
CRl1yC700EQq16o3oi4IUX3tvFH4xOA/UTmaIKdjmMAuxEHNVZJu8KkHL2Ea
2l8H0f1TC1/EKpLtHdaCePlWAhObRCZP+jBTUfGspOG/uG4bfa0GReFPkhyP
n8hQOlOmbjaF9k1tRVw0dTK2HC8lJsGr8V2UcxXdWaTTpXz7OjM1E+ixSM9N
hozZXZ27UsacjzZ/eKFNOPjcTh4o7pkwHvzjK6eiAQOmoAFqLRQusB4fIble
ozeG75/CKRufzFxPHOkQHrRP2bSFB0+iKtEmVR1O+EP0iXCVuVepnIQyNMeK
5brtKTuU3g3aGBdlgVrusPTziokb/Bg6LK+JGq+gq8P+0slWE1xDiVA6yrSC
uN/HLlMQEEIUI0PXbSdR/rSLyN1u/0VrWuqWn3wfiF084TQDjVJqWl7j8JgG
cnvippBUOrWwkQCkRwUlTtGFsTp52nLflgmr7MH80NuuYDErHDWup8xLoQuC
lXEEG7WELccg3Bwakx8GjYzYSLUxqMMfbWxmO35Qe9CI5T4E/E7lP2lEXa0N
FO3ZhIZTcE978eoALo85ji7l9aRQwRlHlM7WrqXDZSIG9LFSXZ0pdNzLXB8b
felVaps1XTrLuHxNQe7e43h3d0DuYI+bznzKCDQXrHarVCEShc3UUmWWGthJ
BAENSkbVDc8wwaBWr9hoqOQLqv+RFwfEUiBBjQJN6TLgUTPFm9Hau3m20/lB
FmPM4SgbjJidVEIEXH2YpUXmuvy3VdYIf6OQVC8EU1foG3ArCVHMWFNCRSY+
sGDVMMBd2WAc0ybSP825SmB+reV3W7cGh03mlA+3OFgGzESoqmEbt/UrLCXs
59smHLrUYz1UZDS4gTLkfVX9+OYHrxXedXOLZ4PaQKIZi4xMCxiqLwVEYH5g
Zjo7kZL8zD7py7I4KxO/KFTOFxWyv4zKRGCEuz2fFocQrCDEP+n0kB9Sa539
wFYQ5gtE/Oh8UDUeVaZ6Mw+j4JulqLZoGJID8NXV7GbPmIv6QJl/qnrEj4Cs
wmLBD2hUx3t+PN5DnEdkIfsOgw9OTV6CX6/B8XbgPlguIRi5wVBGd8ViSAAR
UFQktKhPQVR6FR5/np46yAO+ej4BSA9bM0pzC7MrvoajfsBAxDe6JBWu4HS4
gfiJPJnR06VXBWjeVVytBfMTfOZ0qwbJuUfVtJCPEfLZf8+WuyFpOJ/suDcT
0wOqO+qtedKTLo2QiGIvtkN8tiecDzuw6Wd9Y1YJK1bNlNPOsbX/CJ8NLVyD
wCPKBUBf+OpTjBrXSxVVRpfjssae4Vo4E09suTQ3nHtYj74xrL6h49K637r+
Ost3W36AGoEHYXII496pyxBWVeFZAu+CcI6GLJmtVY0Jz0fTM11ekI+I2NBS
IdLTUGJZNyYLYiCsqMlH4Z6rkxs0R7ZfwXTeE0gP1Jmfu0LmbhpeCXCo0VPG
U0n2su4Qu/tMLsPtp5PaMreTZYREDotOCGsKfqbjX9oN7n4tC1PuZGVI9lSf
mggGuP1GyHVdR0Yco2tfRGhcqufBp+qrxDKc8ZQ6zUiKCLlCFLfD1RA0udNs
os9zJn/GZf1P8qRh6rpsjXlKK2D5pGwbpytAHZMgmIMbmOQpYctz0HY7huD4
9/SsR6Vd0ZyG4BqZ/bq5QxhlJGjQOJ7BHvnd0Vfcxcip/wtJknU+QN6k2GWY
gfv4cz/3NuCHl5GApvJjzdjckmgm+0HXMvZaZb2GKilgtnlBc3de832Ec8BW
Pz4U+gYHOmUkIYugh3VJtbNC3jBC0jjO4zceTGQigRrJMwW8UTfqnDycNacz
Y42+GRbK3lBitcmmJ5U2QB4MfoqUvHJNQfLqUzqUCDAsz0nmyVwJ6ZARUU63
IyAGhGLoVsoh0IIFcPOqANp5Te7bqoX7VB7cvYns1W6sEUfgmEDHmIRdZeaN
50P8Kk841GU+fcsSV5Z9CjfKloDzEeqJaC9V+q9J7c9jLrIWKcPaFmOWsqVI
56zkvXieWtzKd7MbZnhsEzuSbA23bsgiwPA86Kta0c3+oJ57pLrprvZaUcHj
pI6sFXJdTqn+eKFRPsZ0tbznFLwerRCVgPrMqsOy8gs9/fDad6UfzVmuFu81
jYhCX0cf8DZ+yQe7UMdwulnQe0UZI96SKkrpkoGHT54SOBRFvfU3STn5nZoZ
adZJGn6eSMCKbQKAiOJIm9PWMFkukOY22waeWePq2ZKFxY2BAMaIUH5Pf+c0
kR7CL1ccmMr/g7XWDPjBTEd6Kmk1eUPacPpWIOnxfy9tiQN0JmejGZ5z/a3U
w9095snahHRl9e9KBVvD4aEHwN9KMwK31wh3T1j/oQjAKBvLtrejh+/HLUEG
aD+7M9fnli219BuL//XTc/Je9meSK5/Oqi7F4Fi8+x5wz02hnk0Mc+zUNUiX
a6+2sB/N57ATWarB/modCoOZNyjYe5pamMRJNtuI33Zp4TVVz7E+cs9+MB+I
w2RekVmrc9YF48OK5wxlrY378/uFn+8ypJeWWm7Aq58y6zzkX4vJs+ZLU0tw
rZull8RvT/xh+79cT0hVOYLXAQ15kfaQBetH8IhnF1My3MLhXT73FSj9UboS
yqvO/2rgg1ht01wSoW0929CS3+5zkByl1tC29lNvUb9KDt54TC5ubvI94Uwu
8KoDZwIgM0q5r257oDQDPBIhcqGmJ93a/eLGUpm0Kfu3oOJNF+hMyRXYLseB
/kqXtXFJNcdCbGd7mlv0XimV64hOOGO8VVfGWalkAMu/hVvjWNBEa5ehzni7
WuE0HEA+m5DPzeS0TPz/EmcvVRlq09GZLi95Z6E/iJa700uDlUFMdNtGNpMu
Pt5xcfXRy70HqmbNO05RWUfSBaLeky4Ea/WLge7DtMDAYMUBPfiUsIRjmZ+A
UlTNjjctP+ONpxQSVS0Mi+K/WH74vY3on5Pfg3vRKYnEAMbWjkYga0Tt49UL
rRDFwQ71vEXcfdOKM+AuDmBa/yClAEZ816sd18Qn0Mpl5tlEF+ysvQKrocIl
G/BdScUeTb/pN2MqN/XHiMqOdDPf4bX6nae0MfOlpm0gHNkhgs+Vk21xggVf
rc+eZUK2vXgBAz/HvyZ+q4apFIGHeMADp2NPNauzu5kl3YP/sTF8XoJ5K42M
xn7XjcQ27fq1nV+/3rKymwe5LgLo+1MJ2Aj/C68ce6o3RpOj2rueDY0kbghZ
cTWZ9fAnPrjpY1gax8hMgO908XGCoGv/RFeZxOTUs7rDUG2fG8a3KZKyPN0Y
bncCEM2c6+yQOcYjR4dQr8Q8vhHJd1HggvvINiayTcWU0cenaHcOTntuflB+
IgNxTbhhXXqm91zo7reMc52YwB1WQMtgQ3JvPtra+gBpRVu1KW9XHMNmX45v
ABidEfZeHXUh0lE5QMmfEtjt8/YANakNW3P4YA7pFc2HrS0EoJTyxwz+T7a1
LZNqk0Fv0W3cPT8bH0J6D4m5rl//tS752XwQ3sqNrhqt8XikpCV9nO2BgRww
aWKJHCSpoYT71TjoX+haW7soz6w6JZQ1/UY/YI2S1aHhwnycz2aMuzaV2EhC
aZT3uWZB5HSc+ZXyhgNAnXezI3Jx+q+Anc0QnZ2CRkX/BZe2cOVFSAJEb8WV
6iBDCNIEPkk8zmaJGGkfrScRGq0rzK6cTcOqHU6XxVKsWsE+ocmEaac6rRA4
q8zoYc9Q7P2iNrd5pLXBYUrNvT7OOjj6mscnJKAGxwaGU96RIM1kEJ74v/Pn
AbN/Ts07fMCGObpeEtKXrxzMmf9tCvMgXSiiWFpUAlz1TrN+OrN7ONoXynLJ
LKC1p6SbXyUtuTAQC3fcY1SnoYn0JJ5FpFxSRULURHSnjro6zr7jSF9CNpGO
kw4S9X+SeCJHbnrtuXDsOqOlB4iQjnskftON1HH0nuV59/kBgKuFjwvGXGmN
Dh+13PLNqKX7b7gDjhfBKPHKsxl2u3TyryvZ3puAdz2078d8avRGYeNAsI7q
Xy9vtWE9ahZZimgksC3CXM9Z2qWRHUZYoN9Q1qXmECakgDENQa0pgWIcA41X
L72vk/8ufBvgcdfC2qCqS9EfDB0IntJCsZAiM9hkRrmPzsxYDcodod0oi5Re
TSXJs+XZhZmUtcA8rxdD9h3Hp/EpRaUmGpmxOj7qWr1xcOZx++rFPpfUBGos
ufN8lDTU7TuYp+MPXfJpm+OK2l/KR2e38/NMw060HUY7wp7HPiFTDPyRFHHM
5aIr5v3O7tJWw4ABEQSI+VUjPfjjiy3GePjZm5tVxWuhq/NN9l7YNl6X49t8
Q3cZG0lOqB5XT60HA15q3gsQQmDPCp1ZYXETyd5n84kEtPxmYXiA0yOr3Hv5
Ez/c2ySdBDYJz5X7Fj582fS3ljQ/OzJFHAr6ckEGTBKXxa5Ilo9ZYvruJt50
rGMcjhzvnDTdvhRYSs/L6BjSEpB/Uby9jXVYMUa8K19adSOlOzvbbKbQVwgx
bw4zDnDx+Sye05K7CKYvODZGM7wqaVWeDBGzBhl4jueodf5ZoSt6NskxsM5H
N1y3efhv5nBoCTlgv8t/yVzzaAEx1BfmIU8P+OvvY1omr9FXVO88w0fsrlju
q+kNSmtjDrzCc6UX9Y/G5s50WFELwCqRtJedG0ID46tRzYdOLqGRouJsYkWk
HgdBWzeTSKqqwRihtLa86uZp3eZjsjZiWIaZd3JtFoenBh2POMnEQhCNf0nw
tL/WNJCnRPQVyyhAofRTZUv60RxsDDy5+chvpBsfGDmAVpKqgTd0loeWJ59Z
0bZ6J9fyOAS34Inkh4nym2Lr18emSlS/QeUKCRANmNHHpZjTznveZyTCcCHS
a9iqKf0BNn7dsMWv5YYVNULTRPFwrO+F8JsL6nvaYJPa/YKu+gSzGYHq4BFL
k1db//r3NtMpw92ykEhrM3FXXNCS0mSORxHZVhbjiiQYZR1FE5WCiPuSXNyq
DtXPav+b5ZQkylVixuDrb51WrnHkNjill9N8RfCmlkp2sIPWq0KTnTuQ/2ec
jEVFFKctOFQF/PBohtac9RPzW+NkK5bXjc8FI29ld52gWXSocqwVQv9KaYsf
5KSch1DYvXVvyRV+9oZnLbS8rnSkTaYfOkPceHJkUZPg/1wGz7HBr7bSmGTu
QBuixsM31ceNv84iiaJOvHYcKdSEKhh25BSM8oauGxilp/R/rR7gDmj3gSHt
ibJ9bG+VGo11miKPx+8RoTjsLRlxb4OE/KkUMVQKoLkENKqs2+PfjCGxYcBn
r2W5pa52ygmHDkFComsheEHu+jJWT0jpZLJTed6/NrIBLRGCXVNpYFs6FMKo
gwmaa4Jm6xpFAvXJr4CHjm8aIWH6z9+7Do4KmH3zN7X3pW030zWj/OqgsMZc
X734RJWIBJ2KcfDKsMBlw2FanRdx+tybeA96dwGrWcRCu2AGjEhIndXXNgla
9NntxJrveV89DEspYcRohqFOpOJwpP6nSiaL3sW7XZJEVUiPYgKvDjEjfiQh
Fk1tbTfuhlHn94J25dV49Pun0pBRDR97EAB4mqOvtaSlJ2sDHgs3w8CBTVGk
ot42XfGikUcw9u62EelXhy1thqrh0XGmmE+E1Ww7+h3pu+5TnHeCxHCRVP9l
7GmzecZkgE2RS3o9q9YobYU/0T1jojDcuE/gyPbfmhtIUg8ki9DJIM9nsK0G
hKb7fDpTLGde+IXh1WaG+eRhLUJxtpJkg2I9t29Uix7FFAtQbHh5SwigJrxH
1gMC0WJFKghmjrGGzlunej4EJh2z8lw+skRM3KhQdkJWG2pz95bbsWMuSNjT
QYe2OyVk4g4dgn4O5jsyUaAXx3PnGS4N7NUlBzQY0MYZr/ICMzCtDTO1Mw63
xC1LjYWhShfnaVs455OjpsyanR7fuAXFi+QmLpviZZnSnBKo0fHW2/jdCe7h
1ZMVma+RYG3jkYuAnu7ip3xuSSE8enLaHK1IJrTSLdnN185LP7nx8r4SDdm9
dyNVy8Hs3hTdSwz7SYqT7ZUeuedbgdBd2sX4tgW4KJsJ0BtZyW2Exbo5xAPw
hTpNutFNakR5dVIuw4aEAGUvMg4DhN1KYXq3dGSJGuCWMMsWvMAPC1o4Ex6F
bgWTB3yEU+in46ij+ZEees8P4ERkJl9lHULA4qsYZfyzVE5JtDaZT1swWXzm
9S4+uCSQHmDXNpHAcza16wSX+52nP5F3H+v1VaV/Z3u/wKlSHcFJU3EMe097
blpapOBiriHNpOlvw66+xJEirSWIFU5fpPLWde165A3/m6PA5o1WlXsac0Am
vAbS8MqakBtVQfsaVDev5NVEI+omTRBgfWlBOFjVXp0JP1fS8Y2HENTjlqbH
X0z6YxStltKFCGWtZPb4yzHY9diQSWuFPzoRj5odWcsVAj4W4qkwsALZSVCX
vWDAsTHRrODZMAkHw3uzAlkqzxUk5nPRnoDJSKUNn98G/3EA+o99FYLeaboa
muc7VCCTPIczdAdo1M9RRkBdazcJNCaFmLQ0zvq/IwFoKQm7KKuAEusxiItG
GGP6XZVomK1NCIFLs/l6JiI4Su5SDBbE0WE7e+IbzW4g8t6egfVWZpMbteon
B+jioH9Ld3ebX2BGmV8sEH49phXIT/AemtegYN9ox5uhrXTGPG1HNA/aoRWx
6oDiEXu/YPDfoJM9QqX7nqMh0ATbZfLKY36JGcIbCDRSLaJnjhGZS5CLiGu/
5BViV8AMy+2ldiO+Bg9uXa5AX1D5AYV9d18p619HHhnWAoD8Ch1wZ50UM01D
1okoQtsiB01Cfd2Mz10mjAx9I1VyvzqBzALb+J815iw1isPGzv40779up+p+
4rWovUK6GO/lvcTlPKaSWbToOJAspnapbaf7irxy22dNkFrU4dgas/kunkIF
7HvVrybMBq2MkCH+afuqtimbnZ4xaw88WwR9/zemnR47OZ17pcNdkh+62BOS
fSb7LpAfd4H/ulJ9r2VHlV/Owp5Tzip6RY9/VgC1Ct7ALgXEeMU66ZsheyYg
ItzeMkkYBEWjERiUX2IoGgrGTzK7lZw5XU5IoyxtcKy1XqiN1AYyTMoMORdm
BRj6WAuz5Pdmh6L435JaHYBLyfUHRu1Ep5naYE+gkow8Uv0d5IrDtjOB1PAZ
urumzBtdtcXpyO6AOjHv5rSFYxHGhf09jmMvu11vR0jRl4sNVpRl9N83HAzD
KbHLCYA5WA+F+lADksLAbiEYFwDHjMVB23jitvBF+RUd/Mx71cf71jzWskOc
FphHtr4atDQypjNkWLXWO2sq0XWbPymovKbVzkaNPizTH19nykfL2wBiq56S
mrj5NqpO103lGqKngtS7id9Vv+tQIakoyqFTAwMKaB4g9GMp9ZNkwjg+aRTw
nYlZ2EetZUg+k7XDUAhvkYIb9nvtnsoHtbEPiC+HoHDeoEJV8+zbfthm0GZt
Fgcx40Ev3eAIR7w4r1kJYtbphAYWEE8F8LvQzJT63W5rapEkmgyGIiKRs5P8
iwpTFUsw6RZ1GNNbzCHA/AhqtOawvaLusxIBc5c4O68uua2A8i9qA28U48LK
sFY2V4/LEc9xDIGLndArMQzLw7hfkXQIGASSqw5cgiPYlnF2Y/aVsVBvivrQ
o8OM9s+y0O8NJnTWHonYRRCj0i+gQd7GouAhNA9NKfL4BxGUEs6u87FNj6aP
safYiasuGEVV6RWUwi0IKCQaDMrNChLMrJ1wQf2sEGU6wXnK+MteWk1qlqiC
uXO0+/ksKzwawt/6ie9j5B4xgv6BAPIF09cnSxO3nlleLdUgdx/yYZxG0n+/
Oj7fN1JZUc6ZNNT9xzX3RDMy2Ym1zh44D//cduWtNc8lwIqmVx39CrZfAsl9
V+9H9NF2eDd78OQfR/OiJqVsl0E/7drCMzcKE9CL2+HlnGe89ixxbw7szo1s
tewKibH8hg/Ts+3isup397/86TK5WKAoxWwzGFp/SCnsUkEiVAHL/Y4spehr
5IVFwm1loYeOJ+/TQF5H+mJq+RjoBAy/vF5ebH4/Rmq5Zejo1FwDsEAcLnEA
jNJY9z0mu8sPHulTKhLM4DsF7XtbEiCz8vc2yJgLugT6HnWyJwR4eRzWnL7/
Nf5cOHlwuqswHqxn8AQ3jKuFyfLhOb2aXOuCxCu+HsuRkRNi9hVyM9h2qUMZ
JjA7DvuuzsXffmvS3VnWlEYsdi6lHHpKisBYkzUWT+rAh/Fx1Pn14lQD+/Ue
sOSNQ7R6OF9Qd6Z4R2aAB7GbFmJs8YIvrFmQSMXLg4yMeG8WsBBbVNso+zno
8sdqPhmfunKPhFMKtoBuPBbo2cTd8bkJJqs2yRLDl0NigS4CPsZUo2ppEByN
lJwvJ8iHEH3XuMUEWjl7NL8ofsMovXVVWy9EOEa7YKWRDRRTI5fHGeIQQJFD
ADVgsj8OALuwqBTGjv/xxUAEARirMQ6ZRrS4OBY8H+q10RmTZHDFOsDb6Z86
NVe+P1I6sZgGW9Ubie0VfeYSBIow1IoiUhjsJd3C5lIWutKLEXkfI2/2JgLN
E9Icv5VjgU64y3sS57NiTN6PH/zx46toA2NZmleIQ76PojukYH7bjLC+5r8G
1RdTP48zS+bRjAqMkMzVMAUBYqyGTobp3JYqF0+noGFF5LazWeuj2axWUX/K
+g9aLFK3nomALChHzI2AMXkUFUKCRiHJNJ2zcHpXBa3xR9KbCtFu6+zePsmL
AxhQrXOPpnSJkVFpxjlyiPBJVIWDfzXod2JcuF9EWkIXHpqiEJU0D7m9RRjB
DP9Ja8X+sOjIw38dOnHeDTVXXkUZsRIdnqWCcq6RUsX69MRbb//DfcyxAd5n
Bb6/djeJxRFg9E6dHUO0biqbtPYKdp0031/NeZf0ncSP8L4a1k6/mEe5FOXe
o7r2e1dMP+Pvdd1zfO4Ohb/tcK48ca4QfjCG3sGHo2tTRG/l3HiyIgIm5f+A
Otb20QSez6dZLKgSdO9sSpMWfai9NKy/+mxFdHDM82jK7ZZ4Dx8YYcHSCyyG
G4Xv6p3VrLpmeN8Ibjsax4kDoxcw49PPxrHVRFUsW+mryVFuSaUhhobc4jS9
JHvA+cwJlvRtZuUZPdAA46zrdmno6+TzGQJ2WpeckqxAG6iDxqv2fuDiPDbG
nO9zPOH9IGxdig+1V6D2Dq1oZka0+oLuO7CauDqucYsk5P3HlncTXxvOE3iq
D1kJVCzKCgv9Unfrjxs88Mct2Q0UJ9oncnNPt/xrRvKD79JxD7GcsyPG2PD2
omwzF8tfym8BAVYqanIQAZh1S97LNQBgguOer5z0icAE7YgHygaeZxumx0pe
FePX+PNvQF9qFpR/3o+wFqmaA2e/vSvJv9z3Bo6XMSMwkNMkaZpHCZySiAJ6
MLAF2Jab2X+uBwaeO2ADuPIuT7sFSkqY7OmiChoVJHo6u95PPJ+AQa3V//3Q
gSGl0keKyb/YsrKiBoRuNMrCZ3qtCY4bG66F29CmJ8jV+91CGHxSgOzomBRB
v9hVAK1+erAhmLjoEKvWGAOxNKa4UOPshVIgjpeVHvuNvfeTG75LZ6fpwW2U
72dbnSdiwfTYtT9cR6vgA3uF4YR1gG/qb+0afPQYHL4dl/0slBez9dK8YQmX
CYaBSReQjh+FgiBGEYwgZ8uc1zptHb8eO81XOKBynKfvBAQYVyVZgxRZtTjj
eRTCxJUs66A0CWVLl+jM4ZX+LD7T9g7HdhypubqUzb3cxD3vBBtRAMy8Vdn9
WhyM7B7j4JUhB0eh6wfEg63cT6NLaSAHFYAE1MUNvft4dYdtil9UrNUgH7+r
/zqIF3Jw7+H4egtoMwFILY0O8xjrnCtpaSBN1ZG/qMQEdE/Ftbf7C/qcLLXw
7jMGjopfjhX8QpNmDrPnSkFnILi5uUr2EZ7m5JVRsZ3N/QMHzH8+uG/aFfhp
C+eycI/QYsP6l5TMfROpQXqsXsjm0nhXwasGssIpL/awu/B+TtU9A6tcmkFd
FHwaucu2cc7qkYBfIazEsggdxFqPjJLUAfhEpG+rdTucpanke+tB6Vgq3Xgh
9+fQ7FPwOrQkw74dLKnLf6TNjyaqcrMFfTeyh3MyjW2Y0djpIGujDE7IA5uW
YI1IbWJwWSIJAck7rT0c1XnU1TnJDCez7vhCtNnyJkHoDGvuNiPMEdelH6ga
AviUlGYutxTBXtHjem1IeDoK8E70/D94xvv5J4Q+7dQh5BFd/u0SKNP0ipYT
YMStEDBH3UVtbQcR+aazThJNN01HHOfAfu8EtzkRZyGqOdZeaLLeDfNLZB7O
v6TKnp8A/19yKVns6GXR8m/kWY52fbAB1m4KbLo26pYfdi1aLRYNY6FBJOS/
VngiW9BLmkFjKGBT6VZ6oivRrosIs6MVJ0es22orFmn2q/If/sAka/aALeGf
E15vxfiT35gb3s1MScRtgcwwowxoEeJjWyHxZZedafOutqU9LvHGRiuZuWra
teqtSRZul9NAvFkkvpZE9IVeor42fmH5jApOy04/1joayW2bi683RWMkgTEF
qkNyhWysYysR2pUTQwUSZHNwNWlJFfgNJM1Sq4f85PtckpzOq0POSLLgQhDH
v7DfqoJDQSMO1do1wEj9zbYSovUrWNrul6Y1LVMeCzplcdaBLH+gn2Rggnpo
GdN+DxPk8rfOomr4F4+3ve0qUnlYcfMWlBBXi7LLBXd+tl5bKVldUf4CT+3r
r4rz6txy58KdUPRLFe4S47DKP9G4qsdVo3Zhm+utedyO4k9Z+Q39BqoHzr5a
WcGuMxAQE1MNQ08kL1ZGoe97M04yjqhn69pCP5xNhs64O1FPGfeCGiBqNVrV
d8pDkqAQ6ZeOCY2GCDIrHaRrkfF4OtwJ7tUvXbnZ10Vz+7q9/nZwcWJX0FBV
0K+cxkb66ftNbGKfkyfe5p/HS5dpl1VafTdwK/uooKf8Azj0UzAM0yTdlH8M
it4vPZEkZ1lwYtqhwC8Ndqb1hj+cQfLqPwQ+a/vSQIUPSrEQkNmuRWxCgV3K
qL1fY3ltXgQzFwUMQkuXLIomoIGZBkDuCk/6rQ74zKgmaNQjFbmJhTvFkaK8
EDrytPAQDr8IpUmi8UhwyBl3VGDgkXp/0/7y785B3nWWgkXDgCYQstBKI/qu
5Vq/3ydlZLfBiiHhPD90o1/fr/VoQT6BNkqI5POaEBlzgj85Hd71EodUXZMo
SaCgQzGyyzQWb/KiJVqALSPm18++NY9AA855oCN7eW7wt1QW/Z0uWVwAs0st
1oF5jNMHrxuePT3SrcHysVElGK3kqy44uHl9nT2zcj15xaExD5z4dbFNkEU+
Ps/xQ2etbyRFFiGkhUQ/XjpFwSjQSdQ4reIt3quWGXo7CeWjqdhtVi0ajxXy
J9bxqmFtl3HzRJ/0gjcqVaa4A1jxEErIagEN/3nnEJ4iOm71hjT2ljR9dFeN
vYzO6YtY2cNyomJOmrZbJ2Z1fvNYfrfol6qYqWqA8CgEsb8cGkseIGPnlwKH
zghmAU0aq3e22/OaamTl/2BRFTR7xP/agIPi/f7a61ubZJNjfDOxsgLq8Z4Y
EI3VNGc6vh7Sa3IMXTF9uFAgxB8yMHP0mSqVUimGWCZ8TyEr0jG4Peb1jS5O
PtyI0hOcwMaxoJbVlsCxYcTskF1YgtlCIzWWu6/MqRDp7kRuRz2HnKTvpIwH
fr5Afenv6bqmLxPhPQfMIae7o114MW9wOP1905O49x6voLSg5cy1eVvj+rfe
Kpk6oQJGxyfcAIfS4Y0LHugwTaH+A2c9r27SrfM+f1JEGQes6B+9jO8zoSCv
9zXTecHJC+nGPrNj3gFy6Q+wWEFYkmE2CQG1jHkRpFfbBNiKhML1LLwo2NNR
q5HsNFJzLG91boWo4A92siL7LfPfKb3lYPdt1vtOEKSR/wn85N4s3mJHW2Vt
/1tRsk8XTSbYbHNekvnv91kOLZIowc7s8vuem6mi93E5gpI6JztskzXOXu/O
0zE4vBnFKY/mCI0j5jfgc1BjMzdJOlA+XPqxnh2GbH/OEpUV94aNs/SLJrNu
G06YMLypRgn9XbAy2W9leFI1AgoZuDAzIm4osJ4bAKnMQ1pRUKDXR+9D/MBc
4iGUTPw5XVFRjqOtAk2fMN8De4Zd//G98RR1BT6Px/nsv1+mXC48YMjWmVMa
VC9j66NbEZkUqwJjjeM/BelSCBaJ0xOI82tgdfpmM5qMIIF/6cLQLSIMwAL4
Oc8lJ5c586XOlxUzM9oVSkxpNh1bGZAbGwPjgfkc7wZ30vy4fJdaZEDHyB5V
C01BYKpgKXCLdFYCKnHbSjdrqkCWlvwJPrVRZyRrvHUOx4h4Sg82icrCYK5p
OcO039E2dCiI/zJAOL1X+UYVd9Ex8NoBkvLXHQrC9Hhnv46h2SkRdjFMELMZ
rk2kABWsdNo13y4attF2S5G3atWn/Wz204TEj+JqKCcDvP+chf7RBtwpZrWT
2+E6DY5Ye8YbrI6bbekzzD2zk1BoC4OXUOeBp3sJAxf148ZU8akKGu+EU514
mccD+EWjh2MzWGxN4fWtnizJ9TDtmc+ya7ivB8QA5T2GN5UlUUtQ3J4nMJA2
+AKGENhm6nfz+ICnXDUYIOsHwpmbToEAkjeSXemNHpLXnbPZPeTcKvJXTc7O
WDEqWTUhgy2vIqqz4RnB5tzQZ2qq1gg3lS3PtuXUgXOkCMT7VmAI1wSVNDNj
/IlTbtV2+oFD1R3f2L7ZBmWxeM1+rG9U6JAMvsdaE38v7T+vDYN0/XZCUhmJ
mY/kiYSeducXWjYtVZgoC2ecO2uFehKKm7HbmKkdCE+gh5/t4lMM273QxFhx
Ae2v1CoryJreNirqCpJsrEf6qVLHwYerea49oj0NVMj3jEVu8MsTqOVFbutn
Gqupnvp2cenV6q4lecO6okT9NcPWtilAIKQ5goLZTGd0x0Ox8MZrxmVP/X63
zuJPaYpTebGYruhTz6Yn3FpvK6MjPZVlj/2iKRnDWk/caTNTUbk/caSP26rq
Nj5tYykUZvZHCoxFMKlm22CwLTZONsLU2IgOJeqFjwqYNfVDE0TVTC7rIBSV
XG8719Nu2wjiCHgEZ2CL9AyGKmEy3SZghFlnlNur2ufYEif3rM4lfQ+df46q
E8pDiZ5yYYLSl1+yFRfI+9o5DILF0aecOBcv1fo5tqT0oxxCMwo5XDwP67Nq
p9yAX0B7jpOiJdmzrJBb06F40R9iN1p1s9vg9SQ2n7IpdvkmI2yW2NtMtlRG
6aJUVqqkkpUUHUFutK55dAJ2ViYez0fDpRGUAHH0WpP7+uIZV3AmGlUURsd5
A2nq7w4DW4hRhw9bjEFhRDwzde7D1/ZhLVYP8TqiWbAHhrj80CNBEhiRoXvZ
UCzE0KVYkQv+9y5IawAnGMLfusnZnZ9dsNYyvq9c/ur0bwvVhRN6B2jTC5Eh
NK+DJMFcCswwcs92exbkhe+/tTgc3IV7zzcMkTFEKvf1imXpMu6CWe6wWgib
BUPbmV1VLBMbGyNNvyzclKanX+OjIqDOHM5daptFZbTeHhtAPgvFz6tp44zu
miy4+4AJ9rNkG1ABzoaBpK8OQPkOgbTdYyz7Ly2iOzs5zKCNwfCAo6f7R4Ya
QkbxXxP7JRb4ZM97pizgV7k2rY2xEoKFthVUavK0H+IwXLiUOdRQWf+ummdn
jR+sP1HIi0h0h9Sjvf5M4AEBvjmO0kcmzBtY5OIE1JLqLTbGthWkA7rLP3eH
coyv/k6ouJfW2sRzWSWXSVuacpePfHOeQZ2pG1aCRqix3PvKWIq0femi+8/B
OReB69IJKC4oYId+xY5g2pmjYgs6/Oq3VMWVLIkADAWHKeyF0uNsdI77a4Df
MzbahyHqYTb80oItpAvy5F+/zakwIvy9Yv3cvKka5LeSowKLfJ4cZLxUgaJh
DvbL/QX8lyjcLF2PNnOhB9ikS9nRRakiI39kilxzKscgbw8TajtqIpWLukGE
Ac7On/9J9RSAUuHaOVoySyi3VkUgxNjiwS+ihAr5r7my9UWZIxwISbA0omaO
33eKxMxQ1MJ/IWVOobJu4QOd4uStnxQzxliwAnMAezkNKHFq5R+3J9fZaY7W
iq5wD7yIGY0qVuLOsGpDJasvBjT1fvKMT8DlVTMPODIC+fe+cs6/kF5We+BT
JNXz4BhvxdLOJr/hF2RAuFQLN+p2KlJTGEjf7tUCcHEwgJnF1636Ui6OQPRX
dNSP0LIEHS2/Kc3EaUYbXdTNysjsT910FN9bG4KwuDXK81CXJbmqUnnL/S2g
kpTrNPV1l3BBKTAsmnOvKUvPf4JWrU5TYnWnWpBgISTtV7JN0rVz+tVF6Tf1
hxD8Cu5d+c5L7GeM+LfCuniqPiDGTdoGzl8408LsnrliszIEWPgEPsFtZ4R5
l2Pw95yBgQaBbGUG3kjhesYBlpQ0zbMWg7GvQAtuy/y7B62VnHDgi2On7Pkt
oZnmmSZvI0Hn9T5ofIxZwobC8WmwMUT6blMIyfjdvCMIZ3aaZeh8mEVCh2/d
v/JnRFpzLnsJkPxqY3BtBi8ngSrNVxtgXLv06VOo2va1Sv7C8whsJL7uPG/x
DhjXR0q/5iQqBkoK8DBbE3BM5SnUW8otFnR0rvbmbMP+bzRCtO3YNCPHwSRR
SkzRMydUtblLRZGsNhdIJBDOSfK1ruouBXjYpGTgeaqNUeVk6CRWq/5Vqmfp
u26vCGE0yLmEIvpBTxQHJermyHk1XQ+rkxPOnq6Z90uYy1/yxTpxLNPmoI0/
JGYsbLMhH8HHVk9t2BEIp7T009LXkn2wdPN2HIud+EPDjWhL3lwlK9mNdXNh
eT0leWfKolJ+UsNGfk8t6xTh0mn6Yo8dsd8gXufnEwJVDZxtEAHdnrvGcbDo
tYQY2uAehqtQiXYp2n8fxwa1rN4SUsdTKBZDxdrIQpdjkKgVGgi3RY249oTH
0xgTGuXCcbkmNTQfLgCx/IkEPspT7Sl1CRV15YzdfH4t/k46yO6njlWNY9U2
7edCMZC633B0hxE+WPlej86gcEMU4qK/OrcWw/RzDMUJgddFai/Hx2MTYCQL
9n8SfP4akxF8n78ehleaJ4KbsxdUWQCiS1MAdPWXEhFSzi7wvR6oYsGb02NB
My2GdW2CU6dlqO6NYyJ9jGQMIUUL08Wy9CjWnDvbCCV19JTqVd49ENMQDnco
RTUe6O8n47ZxvXXdBBNTf1vqqt6ojDG2v8IhAmFm2NW3wuSxqy85+DOaX2um
JjwEd0YlJHbq/UXjSB8aZTDWoT3Y44/Vln4jBfcfUu2+HRfg6ZFT5wxM0bAG
gA5ChHyVFmKV4ALSBIgzvyp111WgfSxnU3l/wpq16h6FF29mDvzikW8vDyih
1jbQc26oAEp1bWOYgnd236dFQETLY9iojL0j6Qla+Vh2XDRu3YHIfui8ZGuK
jBpGkP+bvUhr5BWRoFRP/Zsl6Xc+B873MZLF2P53anrxZ7KHa/tC0OLbsX6S
K6GXQiKaxWPqzmHp3U+Yn5Z1t6l4qLm6Cj5K/VFJkl4gq97Xrh5vP66rVov7
589EgzBwyeNHyR7SZgmr31bejx1aWSeeoJll6QpXrFHst5TIJyajXjL/Ki9V
8zTyUCqSg2NFgNfHvojSOIrjEPsaSPOnQduoizRqEbpqKdGdcOglCM7aOtYA
yOyyNmqxEJF2i6hMzAti6YN/+4WulUqB+sGRkIzXwUzAqL2p2qhzIws14Acf
5yZv0l3cXlWmZ+jfZI34GYjPzANaT7i3CHKi/w5Jatr8szbdeoIci8Ze9chH
+Y3B20glrV5s8VWqA6iBuDtxZtTDKErouHCoj+1aS/gOo3XvRgWClHHxMyCK
MkGe3ZQ1Bn8ou5Gn/nNhkwekVEH5DzDYaE56QrKex2OAo8KbkdHIvAtoX63w
X02J0fV5xSUCSnXe4ai5rv5Gn8Hk6Rw6bmuNE3iVCLD4ac0BQNvgSg/0qCVZ
e70rpB4C67uyjpOm4WILkFfsKe+IRvT1oRScf1HFh6ZVYIUfu+ZKoheMw0os
lU+OaYWsyUFYkPjWIDfpe03ODedkGdjAUMJPNt3AbGjheXbC9ISBch1+SPOP
a8XVjkTJbfNyflvJo9780g5nDzJy+VElpLvpOnU90KVKVgoNSC2YNPs+HIQ0
93tofyAu5nGiLHybD6eDy3W2tvOeVgTgM+40Le2u6XPKU4h5ChPqmlp6sH19
BVNTODUbeUcvig5eXSbb9vB11pTDEXuNihrC2ndJrJMx0sQY4KyxRFM4srOZ
ow2ZrtLGK2i9wYGM/ajiwsmRCWiqBkTcrDw93IuyiEAi9uTO0qmnpDNeDCOs
gjit6tp3DxY43wmpadm32ESP+Ph1DRAlfAlEYhnJzBOfaOi8nB0AmtJX/7Qx
ABeTEoLFgA7dtDc0kKzaKgUJUpoabtmhprEuqqmqYLxmwmBgadpZ7GXftqDl
ouqprEdyKGYDS8w2icCCFT8O6mu0EdshpeAWlB9qiDHPVWhhSvdPOddvY3+U
qNGNYMkMljqdAFvnMu6J05RxZzNZuRk5nIkHsZmo4mhfkVF8dfqM9Z52oMat
BRnytn13pOdjmyu49DQ1ASV2f0DfgakcOq9GXdIIE0Mz7mfZtjKp9R60B1bg
+vxEincodqpIV90sIRwy0Ak4r3aoZK/H8oCYVj+iF+jYc03kDGzS4h424Pxe
orebDiZJ/ta7AGt5uqiNRMYUSzHjtu53AdWSzleVNGbQoCi8HVlAH+VrDzgy
K9a2/6f3v9e1SqZ4q4ViAFzG186oiqPMaH/dwpk/tCL/x+XiK07/K1jm8MY2
PfvY56v3IlT6mq3Hk3ZiewF94mvsr/IN65k1lUEFLxu59Rcizdtpuh4S2Id7
ooZNh/gGAF9V2vuDKmhUj+6zu/NxXuCZQGeCmZ3q9l8c2q+88KGOLB8bd4S4
A3YBANrJtGvuSSLN3WTO46PwU8IupO1vk1h8oIlV8FA1Ty+8aBli2ixUloV6
yTMIFuaZ2j8HH32amrlJA6xuARYytuPXLxaPMvmUMezKQcMM8up1xJdctmjG
Tu9Gg460z36peaiJNVbOxc0ZgS/XvQ4ZFaYw7A8haJxzVS3K9BZdiYh3w2et
mrX3gA/QIT4d262j6YZ8pO94a2gIbw7IUvWROgr1prMFmK7Tr6SPcyfWHmEL
AId9JSSGO1N4a8lrd7fb3j9bD5aYwUvHmWK3tzGBan7MT5p9WP7ix69o1Aix
pmIvwJ71RduJ8RHLyhb303Q7CbgX6Ie7Ojj2KzWHGJV62Qg1R3OtROeHjt/x
RswGKAoog4OJBIENr6SmjNCLKQs2sSZJcTLCMtyUjLDdluVZqfBAMvMRfFJ/
1M5trVLu0gZW2dieJlSFSlmpHhM17afhVkC+xIPbCAy6NvjRxWrKNgGEcni3
Hd9uXburbXs31u5nFLczmJQ9+acRE0kjZgzc6fedinZ9mMeQQ8p7qRFZRBwR
OvLW4I0Jhbu8DcTP7Y+wrpr29b8NPn3y5hxA5RZILRfabCD7c1NIVNKlb/vl
LXna+6lVO61Z17EzXcWlXF2b2dBWtwF8BknYy0DHZ4XL757NknO6npfiDAD1
xWjHKS1KG1QvrtYRiP5YwJwfuKe/cDa99uuocOvCyJykydnpeOyeBGIIxE81
X9AmA9CRBGW4vVCkelXqWQBOldzODz0aRIWq4ShLlVpBwndwFIS9OGxDiz1w
aR2LOslhNkvWxiyBf0OjEXEzgqxggh5/Anlha6hBZn/4wX7F39RRegzFwREs
W5nJ57gKvnx8Xg/AAXgntsKFlKft5qWFgpog4tynP1XGQisyNFwtdJ9PmmU2
4445IDSJo5F9rdIQohMGeTPSnYctqKG/OKpJfl2JZL8IgWR93s9BUd9jTOFQ
OicLW7bEkWTb7RLyHM33G4lwMQYfxSuZigm71Z288J0B+SL9C2y3jIbqYn0l
DaUHpj8AZ/AwpLQ3BWH2WxGPGCJrMdBdnd6UwLYdFPYD/RX9sE2SJvezNU4V
ACChbkhU0CGCQtirtN/UHHioGcUieHviq2P6ruleGTfERqu9UtNGvcm8ZZzs
db8vrAXM9fnAo7Inf2mR/wQfl4YbdNv/EXZrnXji8MAB1MvZXVHAwQQTaK7q
ykzmSrzqS8u3nkkinZW5Ha5GgU2x88lJcn63GSp3hUVOmDTbV55+Pb9ckAdH
vqcHjoAlozdeXKCHtaa2WT0Q6C4LxYPC+q0G/Egbs+KwUSWmkW/3dtBOI99B
vG1XzUkgwRRBgKV+vtOCb1g5L33hldDbpi+sd/q3WL1J9F/kW/r8w9qWYYIR
XB24Qqw8Up/zZtd36NHTFg2tVdMyqUXjUrylXU9rdpxWt1melWe/BIzPYEdv
PKiHDqV4nc6SW+U2RYJ691PljlGAW6EAn1h23TeyWu6dak97y9zI38O/9l07
AvRaRGRO0feX5/7zN6+Bbax4rknstMmhiokiZJ4r7XRioGi4XGbiTXJNhJYh
j5lgOSMTGAUSyOoGbKHHCQKh6ksPJK8YEQSav1ujm6gC6wAoAfH73GwjE2oQ
TspI9b3zzq+IxM4+ULGHMOYMqsw2bMfyFcIxuU9xhLdnzi5i2J+YNUrhdpWL
HBHCh1nRhC2ZPWp/J/rduNNxfVlGbpvglPD5r6kZvvNzV4xgqPFnI6IVMdCm
zNknJxVV5QkSPFt+9uKn3amlqkszv2ZGQkI75Iltbl+0ZTZDUcnJFVDJXiGH
ayyC1Y+ivdHZ0i9GsA7j0LGiGpDqAyTDxhfpj5Hy7MuWrtivO2SAdZlODf/V
e1TL25tzkYL27zWI+KgKGIyu8U2f7nYeFJT1EodX6xyj5t8XYgBh0OeIb71Q
DNI2vywcM54xivi8Rfv9j6h/YwD2ymeJf58VEIQM0lu23mncfNGWssO26Qha
DY6Txa5eJXTTMyfNA0X3Opx0fjXGok5y3XZUX6PT0B7V6KJGXBkEk2viBXit
GisyEVVOXYS5zwysU7rf9R0xB+Jay7etAM+pw0VB8uczoNi7x0o2SBF0YEII
mKwa50hwOlqOEofXbyDNTQM8a6/Xkf1dy4u/QhBWUJ+0i3Kgr4HF1KjfSaTs
MWHcjHvmL8WoAWpmb56hyL1jQkKbb0Ku3RjnoqlCcwHv8UC51Y86SqTQ+j96
t66vRnkfSwCKb5ArvLdKuEo8T+rnlfQNG8/majpY1lR4YPLu8rDe6O4/Jy/F
d4BICn2/gQ7sHSEsJNaQWK53AGRv0z3qk7XQigcBYKBdfF4xZ84BC0uinHDJ
6zrOmqphGG6w4GSVwIKXjvgZ6eefJvfKDLxwu5svImZvjjIu4t3q1ql1/S8K
xmzPmBh9uukIMRR2UbGP9MdgN67qH+M8AJdgf/7VPMaI4dDpp1WF0KK0TnlC
V6mjT/L5sBiJ+Lcrw9Kf0Gqst9TmGAmttI57sdPwP1aV/j5i+/j0ZB7MrkgQ
UVI6cvwqvqBNRmJGcffkc8j32zf7ww7Jr/Sw0R6iLDD1XMW0B+sKWW809hPq
0/S3GtAVepmJo/KLfQjGpDxfWou9dcax5YSQwQ9bdYxlv6jv8UAvpjRAUUIo
7uJ/l3C5baQ3nHRiZMfst41ql1u8Wr4X9e0yyAAkjxyHO8rFK3O5BT1m/2uY
rM2Je7Oatxhriq1hEFYhhVE6kUnENIX4GloVUR4r3IR9uO+LokAqoymudWZP
4dWwoZahWt50lPtlYM/17orHoVQWggzKUfxi5kfn2QhfpJbvHbczEXIWW7xE
SlB3XG/uHCtbYrQSn88Xhx/11lSuDmCj7H1kmYbJQGDTcyILf1LyW9J0/L2w
ie1XpMIL+TwhceeElW2ZLc2IvQkkIRwqzcbDFMNp3y9fcfvK99uk74a+h2+E
yCAPY611pR8423ajndVsa0Hy5/Da+baQZfK9H8Li807UviXo1/XvXAfCn1KS
FRdUjzXABf1wq+v/w34B7ce4pBuQ1mn/mCt26dKQ6upl0WMW9zXoDbqxs5tP
P01gO8z0V1FLnD0t8YHN95MpfWS321WYG/u5iU/WqmItO+PHCS0JR3656bnD
V0dSm+gnXBUhaCSS3IkgHirkQbCseSYnZokIAIj2WWjT48VwpmOAs4e/lhd/
NZe5lHeAzdpSv65em0cy25lrCVnEqmbd6LpLOMETS0U/dzUrojsl8ScpSgFZ
+Zdw2RnYN28H6gtUv/BsRjwBGW5M2prR4N1pouXhQcFa8wRmm9cKR2r2xgTu
ax2G3AlkDMFFpkBuZ83wOcpRToY/0hPeitbp16q3c/tqskbl8zCnUJsObMLS
vlh2Q3Zxn1ImEN9t3LkM1NeCQL0MGnC/SbYhS+NCsBrhYx1QNnks4wzbJIxg
VQIX7SOR624j7aa5Nm7W6f5JF63/8isjRl0idiOO7HAwaLrTVeNgEVTiHbOq
7VdMP+lV5thbSGZNuKkg4fb9kVcSf4dVbhvTYkfjOcyh6jGD658fcK2RqwO/
+iw7Ql6rR9PrJwl2cYwR6iHN3sqRrDVt/z13K+EuaZOd9QH+3cLyJdSzb6v7
QGx+qVHqXrMIjIsbBb4q3q1+nS8EJsT/Xgxc6hqej90iP0kjRBmGdMLlrZtn
ScmZBx5l/FJEFECVu4sJOb5Fmg6wjGctJ2gcU2b22tfONT8XHJGdGQGNVujF
KNzPjNbo8Sqcxkml7WX77x3rX9mZF7wtZicFFAnBJU10AxrZgMtham3JopIA
OXmIYPUoopzQlHskZ5Bu4sc1yGTOZjI3OQS/Q0KE4wv8FT7jPul88oEJBsIR
xf1jt9OQsMflgHkgN832RRFjVuJJhAd68aivJHZaMiQFI58OptPhnwAALptK
leeQbGd0zoYDjTVSyC9X48ADyUDa1Fb39VFM8Ek8LKaXHk9tAs8pxklY7RmG
zkIwX+gZUtN5wxkBDb2FizGwnaAJ/Ql8XGwKeig3OS53pVKP1wTEdXwevngf
0Nr9RG2/YYhn+i1FJnIvBDMt0R2tjJSx1dGe7eq3ASkCxzKkLTtRXVBnLevU
qALFVKrmmnU6iwxLAaSaKraNU6PNKEegcrz94uy4NNAXHAonjFYgAKkPt3Lh
DUQJRlLHS3NNz+u3/X86JeYoLsyFKZFe4Rox4CrI9tl6peXcq4aRbNCfTgcd
UBQuRoArMzlGA5h+PBPNeqMWqzjE8EE3F0voQTTC5gCk3T27aaAiL7E/qhAw
Hx+uznpqig1kZynMMdAOdq9Iu3169INfzbBZMt4bSwDWTy9g+xWVxdPdv5cC
FZJgR5N0XOKHZFJLIu8vCUtZFU0ifxNmgPzesfYH1veH/w8dPwAv/f5ItTRK
vMrQ8lOUE3KNbZxNSOrLAxuIAvxK2abzStRkd3U1C6ub/XD3Ex0tCO++ZQNT
IsEOOj4aB4hjFFAZod4UASD8KRFf4k+Oj2GcC8WUflvXx55fMTQ91V5SCOFp
eEguvFRbH4wCOYirIcZSmyfYmBTwl7/bgj4IWfNSezcXMSL+xZCUuQgL6rwk
eDAB7KSyfyCHHnkpu7NzS/6KaFCtdd2Xd8wq4yIV3VzUY9VpIhHedOeAQrzb
KUU6maJTq4i2wzGjSHSWuzZETBSlMgnk96Cz8I3BBiv610UNkCGEEJpMk5rz
wXBTaORqCpCO/JW9jKHHSKYdDuhUoUD7CZlKtojbMm7jQy9zQ7tYmdXXoA/V
KFVx/kGPbZy4hnsiprJ+atuGSAwVTLVFv9HCcQI4Dw8hjU3nrLfhIXDf32Ow
M70Qd4t6ja6XpkrU/xEbTSC6Csj4x7H9XMGpMc3NEHm6UmWI37mkiskbubqh
jSdidAxPOu2DJqk8CxNhTrjUFTF4z0wklhGox+uX6wOl+tRQZZGGNb67XtME
niT40SCyq3VvDQZ8b3wsxauE7usYqik/t4SA99UL2yzs9eL2pVQUW0Adh0sr
b/9cI4d3YjuJi748K9ZM/LXHQLlVvEa5oc79rMvPaVU6SJz/Nniic/FD4vZv
s8gCF438w9I4ZJ0G9a/SzB85EJmV7+CFv9m6lI2Y+1qAjPET0raPQs+aVZOZ
MjwRl/y2nX1NOu1GeQMCNNViE836NSEgWMC6nm8uMc882KvMnzhjCDNuRIVk
O/vCH/8pNKsU0pY1MnanI258eIIn5jqb90FImvLPmLDe0E6jo6tE5JGZ+bss
lWhboExgaFhfP74FzEqcdqcXdYWzirJgim1wytlC6lSNnqLZWRm0AiMbyj2b
B0srdlXLt1csj+TRktSkM3t6gKRxmzxYjpHJGHVne2RbL2DtXY/Q4tlMBEHo
9IioZtogRTOThCuwNXV8AO41t7JEeF7XXACUSQR1u4310XF03vAzF+Nn0xnx
j/LIOcvrRW/cRSaUiw0CzLmOlluNIe15El0CAURdbPXTKo6aefP9vpbU7Dfa
adv4u/Ogr+wIHglsDp/j1INoS2uQ/FFYFVhjkjts+qyDBQWS1AZEC4JYE+y6
XY3pLFNiWAlVJvGpdJ1/MZFPj6t0H7LvHuB3EaU1WUMGx/xjQDAd4esN+G3B
iL5o4vTdrujVnP/acN/k6FZXD2iFzmiA68WDUlkHtzwFv1SIQvF6jBpG1ymx
KUL+Cx4Q8gG17lchM66jyFeVygCwD4/1JFsKNUI3EfPprToyI36F8wv1BD1b
rd14g/HGPSj2KVHEBCNpUeEm0DHgCBFcX/lOhe8GX6IUDBqSFKNwolhmUQTh
INundEFKlMEdFCmPQ+447lRYq0WHIVlqnQ5YQPwOrA76FBxbdfdou+NMwv7P
YB1qA1GEiaDMqiCdAqkjroyKnM6cljkSsY0/Cn28f9WS6xBlc14Vei08QIcE
4LhNlqoEdq/mTfdcBbsSJRDyheTU0UNvo/DebApi2MBe8bzkFd1wlawtss1M
cq718UIx18RusqaKh9V21oVPF0Nvqi15bENMoQUfJqlfYdUpzaJ85umQv4d+
IM/QJro1qzv8p1sOY42EoltwkHPjTBgBd1vMQg11fGckyzQ3xte10jI+g1zz
SuSkmAT16LTh0gKsVUrD06C5wY/jbu8ujous3afRR7B4TaL9Q72haF6+jmR8
ZT6Gq9amzkSJnhEVKsdQZ0vLmu1VzeqfGucyXpjPJijq9NOsv8UQcUNPA1EH
j70S9hriPTunV6QNJ/CRiXg2LD8rsxhqRweBDmLm+3+/5GrO67SRdmrpI6jA
hACm1q0TYVJ/1q4XQty3tW6SanL+3KvPWRWXzxVs/IYNAufr8uqA/1LBUZ4O
DYBATs5pvd2FvcGJXVcHGzQQDWdpV+Ze9FfcdfFd42srZ+KbhnI942Q11jRn
y07DELzwV26qCVrjA/G4OGNv60jbQPGl/HC0KKU+Co536ydHwK5+3kP7e0Sp
Cjk4SX0ADPZBnkPVkLbN8LeapzLoYThG0OYM2RW0vc5qtm8kexbDBEmsPMEY
caqg7eqeEETOIdCLTcatFD8NIawrt/W2YfIBjJ69nfN3mMcar5dx9DjxL9dd
DmsKNiOff30anqU6NNF44RrFgxoc5iMsy3lqkFeubGhmwddIJ5GLnStLQIXX
5mvUQdPQpXmj5UO6vewcuRqKni/SLr2rDb+1kQsdSoElHh2Lq2wgWr3BGGb3
GdFc6GGvCONpCgwFdTzedQiOP0bi4HF7g1ypWsUAfmVdRvXet196U2xwWeJ3
imA1dpZQDaK/nkb4XZfYfIX8dZk9OSLFiD0fp/ptPy6QWagWZ5k42fgZri2q
8GykFHdTEr6ZAApSSg1uzr7EY0hwM8ktc52ZN8MbVc9o2db/ze6DOIjkmtxc
mHn4imfLMt/C7HO2/eHG42P0sQYL88r5eVb5szpCbmfrrNtznQMvePT1oZ51
D9tzgtLhDScQBL9xwygI92vZiUdgAfkrNUVFvGoMA61qs1Icd8UP/EOJXAJG
Ipuz7exJJAxpQSWGUX2ZWxnLMFMcTQrPWqDfPEGIBEHlm2QGxvr2q70P53M2
8PhjO+6bGYec9J1zVi3TYdwmAnEzDkwCMbXPCTU7xQ6JVv3GipPCr9k0fUIM
WdYEl/y8l0PXVIIN3xBpI5uXzl4CHKGshTs7+lAdnx1lh9S5e1HTg+ie8Ksd
8XWEPupGJ3qwdXM+MRZuv9ukQqINpm6ICbiNm/5LY5RAXErTnyAb9FwSRwcC
O8JR7aCW6/ZDw+ceZth6vTDRnAyzLF+4TOAYZlsy8BTXIdgNhwaT0ATn2EgD
YZJ6zZPPCgQFoGJliCyE2c2+shEAditWs/NHDKZbmX18HYTkkUP0aeFxozuW
/X+WbbWx0ECs1FwqlW7W00fpBNnlYMHZCW12wzhktz/R9OQqnxWFHsYq/53r
yjW3QuiTeI3X56bmoKraO8214zSfaedwx+ixM4oL1jVcm8nEz4Dbn8orP6SV
YfjA5vmLvW0rtJw/JAuOXZdCsxcTUQAwjkZjdDeI+09RmjxfHPbQ3494Ngkp
f82nA+/o1FqYVoeKI5FN3Ifz8mUs44ZrTo7aEhZLMcYIavq7yYiFFbSpv+d0
9PFntl6WJOkhOhCI9uObK3Lh6EMpg+w5eiFptxeGBiX1XAbv6vQHWLdMCCIh
QG+7Im46ogtAuZxkvboXq4iX2QFvwzAPPXNVAig4nXhwY0UDis4fbuPThQ4X
MIo5KW3kkBFprD4SGlGlyPQ/5GsNgsQQ6yA6L49ory1hsdHsaBDvDpzD1RSV
DJEoEWAajkejcJLCpIj0WdTGjR6danGTSKLLiNhiKKKe0a+yuecV0lETkhGd
E9lx9DXvno1OE7i2MhyodyfpNxOTT5h+wHn0oB9u+LXCJ3OptfaEVpyP202E
0Um+9RJWFJYRvd4yUl7KNGDNNpsf8ckpo8mZNG4nNyyOZh6vVpbY4u+LWD2O
WHtLIKtCqQ3zoXB6WEilgcxpr8D4P1MQsXPye5qWsL8C2u3zvIYb/n2dDEvt
kqnsy+LTwQdLLxHH4Uubddu08xgZXx0HCpP85hbPvEv+wyT9AbYNU7G2o4pk
3NKa/lgedqD1lhn7dBYR10Pzgm1HKVZaXiVifYIdPtsMXwlZJPzUJnWcGuUP
oNNWIOSrKfyCvbEauwJJrvbADJl7Ti/KUvyb1uPrNjeXzmcBzL0zcx7hkbb8
0bhYDTxN1v7x7ICFxpCkTHwFZPgegK31rFjWOXtY5aqQED6sJ8p1w26RmxrD
npuE2pbRQ+OOtBmDQYhno2365QiVrMO/SGUn6oaoUgn7sD+6YV251zYrjXf7
+ou6HQCh24m2OQnNiiIeF4wjopqbxxE1s0d+3pJY+OKbfLAPS67lnJtqjAF5
nPrK2Kkv8RdR+5pc7qzRp4WA4jucp8mK7FyKA6KKFC7nPPFwhbJR00GoPZyF
xzqiBjC/ya3ndeuV/E4MmxQ/QCylZDyLkt60Wy5P5e0KScUKAGWZulwhh9mn
7bgR9gIk+hejxshFnMiPkCNuq35B4UQB8DT8E3C09cWyRZJwFGlL96JK+6fp
jg4LHGJQDFJla6wUZ32+DRaHMforBwG9DKYuXDHBstI7nLp7BYFHMnKMrm6z
cGa+wMJHxrRqN+XXw2NhGKWnxJdBBQb1icRgoHediL56MSQ/NTm2Ts+KlJyo
Z4Y6khnR3sZnmaLejO/c+1NqlvWkIw2Sk6OnGvDdOhLDXH9Z5KF/MIRdSI7N
cWU0XriF50w7dgaaAC1c6RDrJw7+ijusiaRLzLXWzTZ0q3LARDbwLSVSX3G0
lJaXR2n9FhXqAqfshvZbfW1T74m8uDlcPMZHmWhRaonUDQ9bR+MSMBWqD1sU
75uTiP8XMFe4oijZP1F+ZZH/nG8decbDaObpbQd8NMk4XNsRs9aZKZ0wr3V6
3HLU66Jnw1Q9bHcjfasUbfa6AbY5ILjBKGt0HSRt9wcF7r0CpG6bGUp+O5Mz
JJbp3hh2/enubGR2ZyEpk90kyb4x+vdAr6Z8D0MJIIyU0W+sdCGzi4JBJ5R4
AsDXZHn4I8Ex3r0HI6YZAAupxtnYOk0iCsX14v+vyZy1w48njSUfg2wafmYr
I/rNSHNn/A1gawStR9opJVwFxGB0E3J2TC1Hn6137/5HCcglc8eTRofTg6J3
fW43wE/gGTC3/B4FscPtlyJs2DKOmkU4jtDMS1p2Iw+3P7AEG/3WVxKtDlS8
OFjArHmFUhychaSzvcC1da8Jn9M2IwDPrl8KGV3Ven295XCF8txpxA5MU/rj
munPYI6RzZHpK3KK0XXFAyRpMMmNFHZURiblm1li+XUM8kn/5AUVkhrLbkyz
z+IzPAWgtNdfNGWxy7XjKc3hcHazPup70bc3EDvFAIk4ffPoS1pYrJ1xrkxv
xbEiLO1GVs+QKxXuYF4KfTcRIQNnhdybjS1rms/Iz6SDQGLlk07YyvxM6XuN
5kzNzAJqlBz5y9ueC2cnRA5DSdIW8G5ge1hqtpRP/al3a0ERT2xMf0iVfOVm
TQDlHu7zn3ZEBgEOcWFIFPGBbkhGsNz60BYddJuYC2/4bd6y42HEqMFDp1+L
EkPSYKZfW/tC1blX3L0r7aLIEmq+r05FQtM7qHZBlyIHbNwERIlQoAlasRnz
Y0DGlj5LGWc9Bv1DcEZFK6Kr/bp3SeeR7JZiO9H2T8UnX5OwC3aj+zzpZC81
hV1dee4XKmxDrkUH92dMCnUnyzLjs7Zi7z5inOehKnZPDQae6RORLR6Dl/Y+
PbKToOUgcV4EoXMoRTK0Ag89nuVNWdzjgnz5KcTf3grob6s3P+1MDbJDJHhJ
zcs0473VCnsAAnTTXsb0O2RFf+ShmiUTVk1J0rUzZkx/bkIEtP3udF4qka06
gTDLXvJ2aRCBH79WkuG2WJ08pUTVskrzjR8zRMd5U10xbYdGTY6BO4KozYyQ
ohH9uessj3MVpIaT4pFXFqQyQemDVMvJvjZhirvJlQQm1hMaJ9iZOdK3IaMd
VTQuIq80lpoWQpuPw8XmBF3MNHrG5laaz4FNXN8XdpV1pFBKZQqcTScPt9jN
WfmCiRM5me010Ukq9TZFn1q6hWlabv1022SIwnzQkjTDOsY2jO/E/g8mZRsX
gt/aetf0a3iWp33Q16zVTsmyweJvueLPgLfF41019OKa5bCnpUbVlazSKst1
bkU2BQb2Yh+Cd6/nN1vMtiJM6IEX4wY/md/WH8eYjA0VKnlKmjBejOgG6UB7
LIIxNlH72pHOMIG4r13cC50r5GpcB6kVF09PreXj6do9caBLPzPf9H6I/UGw
fbu7cOl3ciFJKR5HYE551nUTjruMwUGUL0hcldPjP/w8RcCANVVAB2kpGASH
wTR8tRWvJ2NsTi1ZEE3BQaL8Y3JCZ9X3QSSxdomLM8IahaRk2fKIS8YngfJm
URqDkKa5azBTdffirshxJFLfyj00SabM0Lguzi6Wkq8KXORX/dW34YLvi6nj
xT9Z/bYGMAMp5ppZlURj4zVoRSmVtqaQAb1bN3bwkb3iWcU2A7z7mHTct4sN
vDXFBAfBwPnHQs56De7tJGRFdaqRWNMK/T7PGm27VebYSDyp/w8uGxZ18ruv
Z+rCl4g+62+hoXMfFjKG+zj4+/z791WYwrHDVbopfmWR+tgZJXhvyirMYchM
tU6Y0CrOnZPrGvgSVtFcx08jWT3tzY6Iz6Et0gvgJBsre5XDHwsO6ZVrfwRz
gqv+ujY+2paiBtlNl2KpA3IlWb8i5/uPmNB8OinYU/Nt60mmk2mSkOhyUs3N
CDQmMx0ZAj6XWE2CKZ8IgdXld4869Hhneq7BhyaVXtXUj1vlBXd4cknoEZUy
I9GY8ZZXoUKaYziLsUwFzOABXZwYSR0N+H7Ur9PaCsmWCk+EawaIq34Cg1H6
b9XM3QKotaBBHLI/GcjhMizJLy0xyhUKiJP0DAuyo90TH5ziL1ly5I8HVLMK
HPpzoDI0BiOjo4e7je5Tg0Ofj8gnaE7G/wuHqB+nHhoFd5GnjsnuwbNSkS8/
TFgzKBLHXuZlyDaTZ/FM8SaBfcmystPINw1yaOB2952PYgM+3kRVYcq/hYGh
RU5SU5RUdyREVPyh4SuF42F5OliiZR38gHN/nIFWCrmWQBHJNZLpfTUtoD1S
YRqshagbGNCEJURCCH5EK/6nZ12OGu7UkBhNe6bvUUbxoPyTx63CQhdiG61w
Db1Ne66y4uxl28BBLMqcZd7Faqpx/UB9P3hIEPaaZK+HcSquIj46x8F3Gpbu
27VmnEt8XVdxx3VGqwv7b/K04hAcWYx6Hx2UNSUhpXFmMO4PxR+eW+uKxlcQ
4MCWb4oUmYOOevueUaXuXJwvCiLZndDEgoLYYTp5lfnG6yhRsqeneWW6UdAK
+Gqz/r4WX6o8RJXZ7B12+vpvpVG/Q+f2FgYm8IawHvWSoB/ZvVhuPG/KBdER
7Vjqib3zEvYhqfX65TG1x4w4N3TqAw2b8xS5WTNtda9z0xqGBrMltkc99vD6
nL+sm2N97ssStIuHUkSorwJ2DHOuzvNruRB0djqxzHSA4Vxysj9smFy/Yfq4
m+NM+fsbtp/9xElUN+EaYgl2KTa5NCsLJ6RrSgaviaGkL6sEOxvYbBzu2Tj0
fy6IdvXthP3y4SSjpbU6hX8IoHDREoRzSnu+O9GnKD72K7gRed/xP8jOa4oA
+pE3UfxKHhC8JZSOZzfz+vUiIeAu9gRBFVFdQA3WJgtkTbPSXQBxRjLyhFGs
XVMHcDZkjMqvKheX8FVKHbXvEtWD+qAbLHwidZpH7hBYMoj5Apko0zawihfw
fmgPSRjf8P/yGMj//5CyPG9jMcRZmO/Dky7NcMH32JKKO9+c5JazhHwBrnPh
sss8cgYXehMmTWpyCpuZbN2i2qYz8tx5CF7OqSECAWdsb6tnpLcwnhuvXrnm
+yIqz4gcaH31exda1GG2M9dk6uva14cF3J6F02cXBJSo75XnAMhefGqjmFQv
qgZ6qpevgDUlCfdjmgQhoT6WHk+b1D0QL6E67yTnhkl7TdcOqC+wZDAbF06a
UlQXlUVQ0HXSSW3Szkf6xcBTvjxph9MAoTzj0T4Ut1TcL3vsO6ezcTa8qdHR
XnzlKhW+rdaDDaTlZK19iOZJWaVcCzArTI60VOVi1lkXfqe60YA6EDrcC6Tl
pdKQq1fP/+PVroS7meIXtv5gWNIOjcg8LyYYvtXgLv7nqp69Q8VmkTmCNUxb
HUeAYYRqupCtP+HEw/EBqhCCAFuwa2PS6LE2ZcHuEcx+Z4prszESODa6uX6Q
OwyrEjxAAH+6afkAw1a7Bh9QAkOKHlk4nOSTmspXLpyjKsTzU4YLLXbdPUBE
2VrAS6WXNullHJXFDbD8DrZYK3gnPtDi5e2KPVfcZfib3Ahma3lJbMcXXVo1
t5CNoj2hinPfuvd/F6hBfmkC8xNDfxn9vtQqziYg55sJz06RscoFMhm5MHX+
h0Vm6rsQtHdvgpwBsmeN6EUpFs75gWMKO53b08zAYk6j6FDBZ7a2nxlSIbEB
6RJ7Pl80VYatV4g19XqmTPLzYMUqaiAKj+4o9NvvvOQGkw9v9HP8P6fXUVVf
65DT4rsK7qiQzp9Hm7BqibRaOSSnuQfe2QpKEme0dh0AHsRW7NAixhY7gIev
qet7mT+N3A4bct/XdCaIPntpKJb/CWJjIx8XIqL03uXSFDsAYxWcwXWmWpvt
4mDjmTugs0asvPX5GwY7eEyLxkBVwE/aB1RcQ7jc5Uska/h8+TdZ5hrcftsP
KT410C/ArD15D+jVKFIVIAGQe6bvQKfzv+6vWzTpUCnxgrhmz3Cb0B6F5SgI
FqGZnDXuND54JBF3QIcHrPME09JDT4/oWlVVHEO/bymbdndY9UBcELRDua/d
qR3wODyMjTCmC++Z+47DeAI4j5KpJBFREz73mC43iRuc9ERpQu39cY99IHiA
8womYzT73gEMsIxRVGpx2byyHK3YzJ8BZ1DxTkd39RO6nZA0MhR6rfaq2+u6
/CfeVfPZ0DjhYYNWgR8q6lql3aP5VCUnPf3wS2niPdmeRt+GBmTrV7gGYJ9k
eHShJUXg8FZ1CrJpP7lnBq7168nBRm891aqoxpZ3yngWKkLriAohRQI7PQjo
uic1yY6oPIn3n7q8C26Dc/OaLownmcN21M/4sxSdvLRkB2On3Nsm/GFzIIZZ
yi7nFMn+uOLrkJkdFZvSbA+DE6ccs+UqaRVjWARUahl5JBU1K/DZklYAiaoG
k3z4mAT/kIAE8h7NzR98vawfv7xzaHxefG1/LTxl+0POUTVIxlYFeVkN7IVi
hZwfC3ShqCxXhHONtZ4hkLvSN+EJOMgLB59Fe9hf1kzFHwmoie8mLPJR1cMe
9GgTd79I/7a643OGnuRkInwHkP8GPEh98XetoYEQJY0o4J3L6S6kanaCzgXf
J2JYSQPIKhgHf1NKpnIcYKIDQUfSx/ZYvNhW/vg5VTsTmbMPQd8GK/lAl5pD
0y46JvOxpxMBzpwguMFSo9I8xKIrpwIan/R7eQJcOc5a1xn+x99hqxEJq9r6
0+lQlOui9/yVwCHSm0lFGx4J/LmsRTP0RP577iy3t1qUgZGfMxgdumpogafg
yt0lUMx6k/obUBbkALxUyYpAfOUUTr3baMOUZd0LM6y7JsQZTMOqpXwSZrGR
Q3KDagXHK6Lq4TOKKgOTwyRYDTcVlcFG13G6mBCX8USkT3UYjLeEc+SXHUhi
mgSvacg1CgQLtdC/WLLPrKfQq2jFw8UuZ8JhFNLI3I6BuqOgXD/aviJ/a7FH
Q41qdqN3Unh+Yp6njHDE+92tKZ86Xlkgfe8fNi4VPdBMO3cgvkRV+s09cokM
6oSQhBtFYJ/xoWDR85NZ1TUSrF+YUDcQFrtdKkiyUifEfl8cB9iRoni5ziTB
Te2+OmqW0UogMC9v8fq7J/Cmq3EyXL7GCOGpFEyFFx7zW11e9beRscCjBqdg
0NOZ+CVBm72xvh6uubqnd4hv6335pIIqmkKumKV0zUdVzyvQHkFEy5oUTQZZ
kmXvcc2Q34202Cp8fPma8UWpHMHnr6RAoQ4jayVV/4GLjbRrv4A1VKQBsqtB
rKDu6umDl+As/2DtYSg51sKmmRThlIRy9oW+ecDBCJKZlYCzpB8B73CZ/jQd
krf9axn+/UJ76nCKNec4qlyOdHSeCzDTYsBUc7HHhdmS/QU3iLcT2scwzkP8
5vFI4TrGQfI+zaHlCGRmLx3GHzVd1D+EMh+0D5F2zwu74fODmRlbUpcJmOVr
dicsWIcwPDuOlLSyFsPI+Lx5c14xh+YyA79V0/iCuQqkca7HZ1FQaaR2tA9l
ylLUqoAbQIm3M3dEW+yzNqsm16OGxdmueC/ADaopf6otUa14PI+f8oyQZOMI
aN67jYsNeYmiyipvGh9XSg5A7VT1ZrCbyvzdaGTlHbDQSmRpxdNyCTTz8LNY
cGxl6o/oTYzVwtyDRRShKMXm7AUcrEyHFExbUmi3SXNRu6DK6b8vr/f6Eshz
6raPTlpj1jxN4wBraP3hzWbt3zti1z7AH17Xsbx3xxhGtkr+TmVPerRGBJ9C
DK9TgRKD6I6fcgq4WvtF2NGOELLW+M1poTNi70MgNVt+d5BfLf7I13pV/zob
tvL3lgPElZSRnvL9XVHBBERzD1oKSsWE6lpkC529WDtwQeBXhmTmoPv0Uesl
PJ8nlqttGPOUNT5lv4Rpbi1M1El2qLQuU/vn+F3gG/PTd83gnxJJuUrlWXp4
vhVgVpZewwv7qTOSXF+Uspt5HKVbCPtwxPakrvQ1mwdKlf7DovlzNWayTw+G
OJ9SU3IwKzcvjweIGZq+juekUeaH9i0zdRSYuwyycZNC3pCkkIYfOwpFN091
ttOO5T6hu+EiJOmCvoEtbsL0+Arz1VL/SKeu7NV6IJc00D1sgXglhlOCUS1c
j+MGZksBgt/TtQwQU8RKZ0DgsRBpcSmjB41RUJN/pqMhvoZjuwfwyYTgPZoA
flwvxQWwPA/k2rjG/RTQlHWMaZqRjGSBy+CbDHXUnDSh8DH1MSQEmbx4rWGN
Ly2h+PX5GJ62KfTSuAS/Oq8r8Lh38Sukc5sevozMQDDbTeVX4FZMAT3bc7GG
LZk7Jasul8piyODlhZQSjU5ZRwUYvrukDdF+SoK0McWlFGW8JfGrZGO76L09
ru1fUBDBp5xmSFCM6aJiHulYdYD5To/jqCk/jO3nJ52mOm9DDHIy7STvU/U6
WVVrFWe5q6gcxghQ+2ADERK0ET+mKRl+A08ej8EhKh1q1HXepx40Emac4T/M
4Gwtnvv1UEbIhCNozXl23QRm5Gt4+h4gC5eMdsABovA0kIOZz0rPnc/aZ8a9
6P+FaBX/Xrt/YXq/JyYdGOsOHcprJ7phcLJ2aYh/pEE+hmfQl37EKpHs5HGN
wkW0zrWZljolui08fuKc4GVJo8z/bauD5RY/7ljkA9i2o8yZys1nJcA96WLl
PVVb327AJSlIdL/xlHmA2zeDe5X24hr7LH4kLdkVRkPTn1+KfD6ksYxVf+G/
+g46jGObxDq/GTJh8nNIpAyIhFmv/NsgRFHxv2knAZm8TbnihY5c1zjBZ5Jo
JYcT+jBrTMkLbWMXui0Cbnk9MHYCN/nNW7+5ZgnRP+eFX4O3DueBQEHva83W
1fJlrehAcZgaJzORSz5yW0eDTgAHRmpNC0Pby3ajIXjPs+UxG3tO6NVik+//
lw5FU0ubHtBOxm3xy6juTv5pHR8Sz2eTvlfm2dRt1xYpX6wzMeyb2icRUREs
HI7wzB1D0PxBiYYKaC3p8sRfKygpwXwNmn2Vc7J2Jwx/cR9wcKjCJlnOm1Gd
ZJqBXd1k4TgFLQ4QNHN53zsupgrnBWw0wMtyyfc8eSKUkxMgmJDxzOsbxPZZ
ZI9miGRck0xVEQvewik7LAS+yi5XrS1nmtMtEHtvpyCiYCMvbd4vUfDwdlOy
3lfWSUb1G2TcJmKf5svqg289tQ4GAOoHzC1nIjtwDMwYsnIZ8YrCH/pgj+pY
rWOa5jfitr14+nJFTLxzBh2C21mJXt0uhH9S+tDdAwp0C3U+bf9jGYohwgTs
YpwZwbD+GI7xZsQZVNL0/9gLvyNdtlRM895YoqEWo/xx+qu+Kg68IA3bHrK4
zloVKaYOSBVnvPaho3OwM8uRtlAKmeHo+4OcOQqXS/QN8DWlaRdzCGvpRDQp
0teXwj8Dzr3b6PwYspKCiqHReQl/JvnuxQ5/nBFTla2DIv0HelbS6D6NhKVh
7U5RPsHRIMUZIoP/rH40P+k9bdYvvuJ+KysND/KfSft4aeaGSNsKuPUKHVnE
PRDIlUwJR6OXTafMKDHkPFSLXAV0vqJ/ZznHAVoH4VpzENqLv9JkJkm6/6oA
6OyA6GyDTPR8oyS0rVNhehQk9EqFat6kb17GgelFfQdFmq+yZWky42tpHbuO
vi/d4bUJSLIwNnFEXaQcy6ufsl2yMvv/g40H0K2NHiTBrtYhBvS0X4kcY8dg
3YkF8xHpBlvCQtcaFmoQyauqFnrWVH9p5J8Q85HHrnYqIYPMQphGn8pHYTqT
PvajL4pd9OJV5RRWdM7bIQe9YYw7GvTtjstELNqq7SV7DtRdO0uKvpl2h274
hBix1gnjGqTUICGPUjvA7d9d8t6J6xyjqwim7IXwC219sxqwp2vBuDDJIcL+
QHrHJv8R1oaIDuk1FGcLxikYkg3w+TCUPYnSYNCqcLIb26FN6hiWy6wIGqu5
Um1TAQ+yMFiynE1H3O3uRr63Pv2oLNj5Kf5PLhKHcwQlHozKHhjr84mzoA5W
xu4g8MLouhbT5g3AfNA7PkOAOGbWplIKzt6phMj/5DkKqNjx3L3yztc/aIcg
vKXRTiqvgex1jfJdDgUeIwAR+EZ+BpyHEVpfNdXdlmMIHj6ecpYcBgPMe6Y4
LLfXrReR6PMdPR92EodRn6WSIKtMEnTjTkaZXxGF0g3QniGFjiYTnBasjbUx
+8DxMdQmGEbTbLR8Xk2Zms0L0on8hUSoFR5NRhXhXKaKaYEwqYBFTRlBsveI
DzC2HwAmDAZLuS08ym31fP8g8xsUlpo3Gho1O0HtDsCf9An4NdKh3w20FLt2
XfZVCtYgb2esUosG16AUtAEzEY8Fbfag9QQGQ9D6l4vtHskGOAPJqFU+a/7I
uLg9uPnsQy2o4ZUbCCdXOqW0qgDgmboVh80tQ7FV1zZnUVhu+hVDWCb9MmVp
iem5jhtlNWm81G5rRqr8m4JCF0sKs7VLKAAThGq5r8nJmZBYJc78/x6hA4Xz
Ojvj34kC6aqhSxd+fUZ+R4dvmLkw9uZFcCUHPZvWIUmguU0l63Djb6JhOdfd
X4TxKs9lGPnluk9/yh3deAnbS5RvB2X3x0RysBpXFxRQhLfSqyffeEwT+kRp
pDJHlfiOAkfkqU92cJ9uBnLjmhQAXTBEyWg+LR8zAqIvmYMwmqH1JeGQbnMK
61zAfUkLa+4B1fQDxioR0b1Y/pduWmQ+HVvIcPIt59dpgGdAbFLcYGSIQWZ/
FxPNKCKrKLcZHeiJxRkeGXeKhqVAwIZcA3VcvonO4JnG3M2C321yAftjM+4y
dNoxQnFv+tITNXesTCEQxPXJZyCnjR6AkCI4xCoQen9RNQdmiYB07wgjBvm3
7Y3lcwpXS/wvOSQa98vnnv7sC/uRYWByuHnbX380ypZIs6ONiDGjFOHIYiXF
bbvpLG6imoEoB6BSIYX3NfGTCHlsqn4hUDASuzbBuNYnDsvxPgVCfHfjD418
TQVPAF3z3aKBW7EvmFje/O/QR+hJFrsxKc/loW2Dg6TpBb75A3wH0EzcAF+p
X/89g5OSuJTaYHEBYEICjOWdDa+duiZXapH9SHqStjNzmqCt64xaJF4e0MaB
oJPjcRD6uqz+bH2oOUHFD3w/J49SAQNk8pQeyoh7hsSS9Ee9fEQoTeXKwfrf
dNHS37KunJTiJGGuB4LLpUJs7BiHhmngdnFRXquDMD0Mp5WXXaUOeI9lVOgy
NYOJMHXL08/QiBx6dWYiF3Jt8/2vk6YkBojRle6JuNK2WsUA9Zg44BNfDgze
GNFo20HpBxf9PCTK1FoqB2Yt65XPLFlt+9V3MT1tzXNunNSlxK76pEWf6j/+
JXnfCN9Aifqoq0V3x6vZdcKtuF1N19HH5WJGi4ZGorfP96H43StauPyPoLL8
GsNdR7DqvpGfYrUWK05roYWp6L2MBQ7xM54ukgw1Dle6iO9/7WD4VOzEHETu
E3nuCDjcmPKGynflomGexQsXsrSvvRYf4DyjvVnPbIugVeXBz/+ZVPrJ2K0x
IOVWc+mmy5fZjHNN7xBdgXzS5dDril0pA1SZCfxiU27PToA7sNBMXlz5F4xw
mFtuPRtHA1aeOqNnyuTH1PRFXfVMnUgtHswzlfMe4Tqc8M72RuR8avryJRGn
+DU4yxbi2hENQo2sL58OxFhj/s5m0YOJ/xuuOCkCazC1eR0XFFD5ekj9ROJW
fY/M+5RP+HFScpZ2IZc2bo022QLZ/H4eFZHGm3ULP4FOhGibyNOojf7Nwbv6
S+qaf4SdPJ08PB6O3Gt2wmoYIAffwFW7kNZLV0w9n+69kbMKGHdoOqki3bnK
Iqdkj98kVh0fUR6QamRZSJ9EqorRNjWPDzAW6KrvmJNxBl9NTc4LY6W9GOVT
nRVKsO2/9ZtK+z0cdiFkYKSqYUhFDxbbkeYpuSu0szrZNUiVYCdgxCkH8z+4
uF/Sup+4eyHby5tFqgBXpReX5JxiI/RlVG23o3rG7VNuXJb26ehu9fMwwCRS
yrwjZa+8qDCFZHiqcghStXSo/1gVP2G9cV2bhlKRA29N4TOR3A1NqX3a9FxD
JUbfv/e4s7fxS09U8tAkZr9mlGUI/w64PGh1XqV0t4MGuZvE5uNeTiMN1vHl
PxaCJwktjxaRlQtr+vG2lJSjZJk5uuUvHF2C14lqA7FrFGkjOrtEGQfFLTJS
777gXTMZTXIDpOGRdTWtxwshOXC5fh0847DKJ/NJ6JBCGJnWS7V/kJDfjUDE
8xhwM6AVSTJdVadtTfILffvyYVGtnA//SvPNYnmunZEFuAm03VWh7j1RsEdv
Eh8zgj3Lc1vWlMwPksaaK1TuujiLv8IlCN8nL86k6jP2yYKFNKvkSdU6wiKm
hXQLN+u8+aZt/DG5EYk0tMiRWphwM9+keNs+v2a2WIBpmIkfi/IYZ0UI3tRB
Iay82BZMjzLkjeBuhQ+NZVZ4Ivc4zr14MqainVVXMt7AiGA/Dn3NMIYiawyQ
tBmDrMe+MKMXrGQttcxJDOaSV3knPs2qGsw9vgS+5e+OCYcuBaUdBe8U/Fof
P/J3677CBbmuRBfhM1QKBUn9YSQhtxyGC/6Waox5e0rFHvCB7lg9sHLtBOXl
0XZBpsRTzsPjy9uxz2oRe7RlwwkoojXYAaqqgMFUdQ6PhQzungzk/TuWYzya
GLSmXNVAJz1Ge5BrAKxGS7Bhd/Zr4UBo5qmYMnajI+sCkurLF0oj7KpkIibl
eT34DGy9jxi/Kuja3O0WY+egO6QrbKsTdE3xQvKgSOrInvnw6uu+R5P+DbGx
zuFP8eZOMIy7gioOwQlOQQCDGdSM+NUwa/JE1KoTdwkdEPobIz92xbOMsto3
XAPRaJy59kBoqZ2hLQz4t6X4RmQAp5HLpLILzPQKojVtdy74VeNj5h/y0xTr
Gj6WZgQb9BeEbwJPcPRT8fXMATKgtbGrUecr+2onoKfZ2JiPwpLpKfyteIZ/
xaiAGaLUE/HQ/R15iWzeFQ92djHWKk7d9XOgo1ZT3Vw2wJB6cswPZN2XqFB5
Gxurt+zghvVWdiH08690rUQLmpWyWw5Gn8RgCF43lZoa6Yo1HhnTELQRt0R5
p252rOwGQqUONwxWRYrUK8QTnEQL3j/HmpXuJyN9OEOg5z31hDFTGtBcRIzK
eh/lVWtVsPjqNpRiWRz/yFBM4MqWjJYawox/Xz9ulnRDNX/+clkMvHvo/MLf
8U5KrpTN5B3uctCVgMrYhRJtDSbJCHSqOL4ZwwBKENhMyyU02vQUb4MhA756
mFGFdj8kj5QPqF8GbHfDArqY0VKZikRKv+EAd9mwSt4H+/ZcfCEWWwTDX1Ue
97VzPZIwdxWK0tyzHIn/Oq/t96giClC0RebnwgbubRu6uy/OSyiDvRTefh9D
hdAMYmazBGhbGKJWW0+t3rsScUe/4SimvtywO0pWIk/mZpnLvS54FVgcOVCT
lZQtln4alkY1CSoysDaFV2luzsV7YR5FXfUSowGVwxy80jsmnjijug5dKFrk
LFXavJt6oY2b/2/gzmOhop6UXvrQya6rDYqQlpy3iB/XwZ+XkYBzGBziX09R
lF0w/6Oz7iq7BcB3eWAljta4UD+CSjHgJHgIjZl/CBKuf1vpKF4PotHZv/8K
TJPvG7sZ2qtlAKwHwexhHh8iSsUW/rC3ZqlX5b2ezyzMliFFG2ve0jlDB3B/
dE4dtn7+IbHVr3HZHt5r4jsYEpkmqC5ka7uQBUspjocUZyJUjE7hAqlZJykC
jn8bj3IG9QVegTTu/+qztOLzSgiGHefQCXcnDwQrKv0AOExeRHLGYQrv0HNv
EBfEh7u2oFZROKkON4Eb5EMtaFCE0iRqu+KNK0+op8rVqNTnaf0+JRFeWaXK
WnO+LecOGHF1lExrtMgh9eDAQzb6KR3SHBFx3VvWIyZocGeBln1EF9wibf+J
TzgUnAA2x2Pq4gk7Pm5boNTsrbReRsUFI1IxNOPOQNg1B7u4QABqDWSzXF2q
CefRjvtS/fWET2U0Wi4ItBD7v/MR/PC4aFC7C84yZ+vJGNIiA3tSdKUJFON4
MqTFepRaefzsWnnwzys3CpZ/fhvpGGybG/SP2H0Ow7oicrLy4CJ8nLmSy9sa
0v9MyefZVQegftEVE50lKq9zpcdTl2sgkdQG8S7EKrnHEIH0UvVDyr9kXa7U
Hjr0EBwwuharXSFQvKouiL1CRBEh6atE/fsIRda8TFzHsF3/vMrNtY49qhzb
BMRCSR7oeXfEVO3NvUe7lZil/NSM4IDy+qUAmd/QCzFkeBSWvCWIFe+mhdXQ
zsLwqKaZUA+qmLXdFEhe8+Byb/w17G9DxuSvRXJbIUhAedgZQFgEPjwIs5kH
j8RaK7lkNYu+XXorULxYlOwwY+XeWKTcW748kTBQN9Kx70Bx/HeKiXHmrbet
E4lhPFyC7rDfjXhYoXImH2vBbU0ZSYm3zmd55JmtX08bEX/2dh71OAmGTPDX
GAalY8oD5hTIE9d93Jt0FquIou9jl1Ozd8qqVG5Z0W99MDE4/rPj8ODW4/XT
OoFxuqgtKQHPfYRp2NcZieOYLoBRZIf7767DU+KT/r7HY/Lt9uKrVqGJQdLv
yspht+exz56pgjZeJA6a8TEHYaNUyc1xojzbiyK2cTH74PlkcI4YOhjxP3Hg
MZAG/pxrpK/7pNtsmGeV3t7zCwgNo+OhHr7c2iJdi6GUM7ayOvsyGHRJNNI0
ZrLCtARJNjrnH1GPF9tl/8mHli7yXx/ATyXfwAz4F7MTIi66vVOw6TeHxNQg
mZBmwuldl40W0tGYzv2E893GhTAEgRQ8ydBBTZjVcwUNOCd5Etd+75OEePv7
wPGMqDggn+dG3DV4LgJhSJMC+hQQ72kC5tMEo+5o2xofT0Tv6kF+ciaQNA/R
uP2rfgsN0LO6zDnLUPUeLcalSucPHhMCvkFGRp6cZPXAjJAAYzZQ2aUoiNg3
5TNq3F7ZCBWTWhu55DuUqVMJ0iGU3blJ/LPQQ/AKBs0atBBg1OGrIJkbHxWo
U6rVfD2cLonYW8HoC5GK3PRkKWdksjX43rML3GU/8gZGjieUNMoTKcRnzNwo
daLy4/KCTwzBp2sVTRwfLgB+KLzVeley28rSOrHgGSERHk65iAZCG49bmOMP
MsgKyLu/iN6M/LA2FF4afhUhZV0NuHpTr3j8jCZX++neXd+U413xaZijyK/Y
yPmpc1eLVED7lG8cIhUKzdQ8AKSr+cCxp2UsoVQKj9zrrOq2rxOfRluvwPdP
AhebR7X5+QmWCLLXDz/4RvKVMY3y/3LMtGevEFh42M+o4Ay2TM31rKE/Voqa
M3AWh89isxFmNlTLy7PClj3fhmEtnLXj6mT5PHUZS6U4umc9k49soV88xNGx
uP5m/i7215PfcW/QFg9ZaKgiIC9PsaH9EogLMMt8/9NtYXyZbQ2XP8LKyhyc
361X6Nw2NZ4xUMQlIfNvLDH4FlG8wnnE6A6WIS324dQyq3hX/wBOw3o8fv0J
SrNngHBGsAgyMFpLXThrZPyWmWOCswow9HXXsWWROeZuQn6qPedPqqC4mkUN
1uBRIuKLEMMBnVORi0HzzCcRXyCvBZF5BtrlARvaY2ACt826WWuC9H+kOpuZ
PaYDPjdWOBU2lUEM0B3Zb1y4PJhXjn08slVRg69Q0IrNeUHW3Oyq+mqzwj4e
FpxspQecUHCet0n05+u0qYiTLbPt7KDORetiWL5pi0f6ltZAPKAwjHmR2uyZ
Lor+R2a3SGRmCsedfN5XvGRsFpMSigHOkeSuenINx9FrZKzDiHsf8QRVsZDS
S3ginisXYVSvH6GUY8JqLODveZhyXRv0efYbXUOzscLhjC4pBhhWmoBOEpJP
5FnZmFhgb8tVWgyv33bZy6zcU1nv8Ops8vCqTwAn2P7TIAziH0IIoMXnyBsS
OFNXWWVl1SvoAvB0T4G/UdeWdaB0ReYRKhiFVVkTARfxr5Ma2RvxF0KXICgl
TtWlnC7z/OAiDOOUhoeRkK+gskp5LeRrFehq2d8z6REr+U/jWObW34XdV7u6
YgNKGqyXVMT+pN6C7uO9h5erprtx5y5LI47ZUvdk9zWIJKUy31VGH0R2eZz6
UuNmSJThlU6cBCEf9rhQQx6g7AbycWmqDZYBvmf2j4XtI4SyrggL93eGLlto
Yuz/usrRMhF0G+mT0mbdqzHichhPu/pxNBHvSGffsCCFsON0FYUCirwdajYX
HFMtjsZJuZf56pLGGUNaz6B082OsVLuB0CVGu+rVqQDgdz4vU0/EYm3lG69Z
MKwWUrj7wr9ns7KFYKx3iu0WYujipbKvBpqcxdoOZCDGEstiR4kLB/k55olI
CAl8Wkhv3McwOEf+CvW4KCoo85EFQbcgjH16iURPUKTnYqqCTCXgWHcaN5HB
8Jx8a1lG3Ocgh5pvyR6ilrHC0QzC7oFfcS2hD5F8ilixhGivsyHSQ+1341ID
LrBMOiO0c7vjd1xOojOJnWRiUrHOzHLqpPyHF9SwyGOJUxZHHS58lN5f91sz
F9YFFG0d6Ig5A4Gr6VQb1BK9he5wg4oFXFUeYIPj3z8vfYRATZHB4tyJdyDp
13igv232+ckPVVplTWuVCdNiu7WggsTqtHnGZPIRxtmih2eDSW+294btNTkq
oGV4VWUW1epYKoPDus1e9RdY5Ul5ltd0+ZrPaaN7g8wQJ+wPcVWbrMwnI8RJ
Ww/sbCQH2siEF4d3YjeUbmxadJi5GcYeVqFsau8gN6i7A1wk2ert3VrWVhz8
RudYDz+cveyq3SC9EZTyNhxwRXkB6ijOkdrgCivZpRO5W3hkTbTtrnmjqOax
PaXHelTN0PsGtfR7BGRIg/d2zbARhUQPmBqoUjZmx7PSEzjJmd16iHL1khKu
3HDJ//vx+jKnbLC8iPhRX3ch4Ihvgnm3gFRuX+wJpZNxesWV4WxzS1N8aff1
eDJFPUzlKucID/M2kAZ+GHBMxogt1+XXqLDbN8OS5kaN2ijVgQfWdWXoNGpR
9eu3XmcmzY8jHv6H3A51DjF5qXIgIZg9YDJZmDPMx7X60n+ydk3DglNa1Q+I
0CjUnlJycE0pDWTYkEiHqWlD8TT+QZAFgdqQUV+qvCJYazzLcFZGP45kBcNr
NNSef2ta4hJuBVE4jmSms/WP86KM6YTAOQJ15jjST8jOLGegiE0XNCX9D0K7
5EtdmIezO90TeLut1agcnukSil8si8mNvzJD85bBIwuB1I5fmVU59ZMsKC0K
o9ey65DeRjAfOKUoEWifNP1DQCrj9zolG6k8HPOMRGciJsOugizG42zygHCC
HksdqG/f1jgUghiuN06Uw/qbOslHyAkWxGUKB4kY/boFAVaGY3wnC761dc2v
0hHqs7bDLGvjo6iBXqiNBDbcdBt10qJ8BTYGvCS4RBS64jYSLJLAwIm1o1f8
e4YjRUBKF8Qa56Erx2xLBbUYo+jC7A2ZrgYHXX5u1AIwP/40Gx+ZnGKnQpcZ
b84FfOI/xcjoF91iYQv+0OPzdfFDyCgRT8VeC3CBstlmB5QmK2cwMO4Whvmo
xwsGv+AqETSyOO1PnRmIRgEsoIknWCUz9ZQZRjAcYYqcIms4uEUVvYrTYy53
lY/mh3QBLcLieRlz+pEAvcvl/RFARNNJopxQ/EQkLR0UFt5fgFpB1Nk8cklg
m054IBFuvu0uoimPZAOoGEPKLGKO6YKZcSnCImkLfyk/LizkNrlyzRPDTQap
o9dkWmMoPdLwUVx7cl1SqELLbhayWzoL52zKtquQxyDpKXU8qbEE+FbAfBNg
paWYGkSM52Zw4sUp2LHati0iWTpkOVppokQSdR0Ws+AQcXNr6mAtYCSJ9SAH
hFi8cUzK9nXziZrFYHb4tneqjw2CHsBPgr2Y2YeZEfpHuzp30bxPhelGsVgt
TH9mkmtufXSEcRypZqHCkrlnu43WffDxgfhlVQkQ5oHDNFN/vQggfZip3AbE
KQt0gI+pTEN38eMGmOR9VOs0ap9TeLQnhQrgbNY1R1jj1NzTH0mbTSJyl3hi
460raABlOQOVN8hzvOxnlUkjLtJANS+gVWSVj8smT9bQ90KuAAVLdpQFcDzh
p9rsJajoDm90fGOHwV6oLcDq0UOk2u5i7OutbBZwYe5Lwdt5haJ5d4lrxH2U
AGD6mjr1GRVljWYh9HHxZ9dwtLzuYo8DxIpFOSL+gXGPPXkfKubH7BN+8RLZ
N9ySnreo3QIclXiQ3ZC5b0M0rOVNIWeV5jM/l4T/lTIY6IBXsr+qUTo9Up+K
qesXDaSJm9kmYIpCu55eD0jsvnc1gpwA81oCUepFLSKOsbbeCcZbUPnif/BZ
LTYdjmbiw6ZtdWc4FjgbaVOz2LXinDY7jF3WvZs0g4qLmJV/wi4AahmaPiL1
18YOY5a0vIpjftqefRxRZJ50WxJ433KNYFoNwpFTPbvzchbFRKVyq2mqh9k1
KrEj6c76noRJGbPcEIbDcWdVVjyE3IdWdTNP3MtgR3qd/TCABK1swIt755fY
O2I42wxZsTlJf0sllOqkzekRUmb7tB7lpwp8Rr6YVh/A4lG2nNMrUoT0s2yT
GAH9qvLeOg6qZToDiMilDJk0ODCofCySVCObyJ0sf0sBPxKCFC6X2ldSlKNY
o5mzsjw+ntDHJTdPuqtDFn6YOMf+EnhoOR2ni9l1qTogBOlX3TwxvGXkVJqV
+sIG0DLDbwk1YcSNnPRqBXpcIs3iLN0AnvSMngpijn7hSjqStpynWpRH0nev
HmixGMuqbGHe42i1gyO2B8reP6ImOGB2RHgOcQGofiGeYXsyGOsTsAJM7VZ3
ZzzvM3mKZNYn7gbfdhhvmHqUhHOmL23TqnzbbrF+nIzFO5N1MugKUrhauz1J
C/sXOpAdBcAT/GYagLa84zhS3SFl7XTHJhrG3CPJ/7COfahzxtFrObgcWl38
jPWovOMPM96XXu+7U16BBtv56lNMZkF/QLLDp72gXcV0bHS8Atd5QDlkYXRq
TzIfwNuhJv0SDDUAJE5KgQs54dNA1sW69HS7CU8d/vqSE9fkCTF4D69UhEBD
8SOolqBpVoQNVqQ0pDANrFKcvlli97+4ng6Lcl2jgC0UQW+kYm5Ng8VI0Oo/
zi2Vfh3+iEliO2qV71mKGMT8x6hvPxJ/YI5xTZkysB5oHArMRATUNVe71ftp
2O50Ib8I4ZLz09VXujSnW3zOmio/K4JaQBulmjL8sK1irNydl1u25q++T0wq
2nNyr2vQDC9dr2gg1E77oVEBVD6ejqQ/anwesWiowLOqXovlp90NWHjO777T
xqSZg1Kcdf9MiaxchAZ8Crv0KPVEotpEomJgxarIybV7ALwJrs7gfWKAIM0w
3Iubx3H7vkaQweDSA29SLUqpUkEtK5ZyRgZJOGAtmBFY4rqbOHo3HEX2yeJ1
h3HwLPfZKjugd6caby4rrVI52oru0yZk6rcrJc5a6kACGaK+pzy5p12KnR81
z3s+YlkCnrfghaJ/fJXH5BYBabDurIE6+5XnDLd70Lwi/9IQYxy7+ZFUTTD0
9oC965Oh4vJAMR46DHQvCOvx7Z5fOeUnmKxWNSroNcYzgF+7SdOxdj7ADo0r
KRZt0EKyRPSzRHL/JAOG8Hil+vNg50BC7x+7kpCopHA4X4zbCzsyCLt+iXsm
YazLezgSdxqkaisy6n3r5S9B9SkAAXQRSYL+IpX5F/7j1LXyaLAot0MfrxKX
4FJmLbqIbdmmbr5HA02ODMx7dECRIYz517gGPMLrbUHgL0P1SQBOR+1IrWzz
gv0dLp1H8qKYUwcmjlFOlpH4PhueYso9XfCaVBLIUXPeny49yD/K81kHFwmI
3vd7QKYZGS45NsGz5PrgtIRZ+yNDRuBuClAGOoX1s4zNMMYavlLmtt/xf6Q/
MfccbdWvCd/a/TGGI/y3sY6hHD7cweG+MSD7s4MC/dfoILxtHjcEMcaKhK+/
DDb8MvbNLktSXznMDM0LLe+rmlCHMo5hTjI7bM0TwiN33ENxoP2SaebVta4F
Gol0WYW40XM7tCycKe61fHm6anZoRP+4Juu3GdxckcZqPE0jpsswqwxrkXPB
Nrv7PjcqU46UsTusDHUaHBOZYdYJcOrf5933o1pTgBRgLoEsm9WU5bHFlJFu
HKvtOG4GhvFjoNuLHtgeuBSePZBYL0BRmELgEGOya4dib3VmfF0f24CHZm2p
wNcRIN3WvmHQWS294icWMDKLXK0I05R2nkhy15928iPvWTWGVYEYCuyUy3f8
UfFQL2LUPux1uiQFRyt7oUbCBhLMJd/BKvFIddL6iN8BX4oVeWcK3ZLnY5WI
vsApEyfRBOAIqWi8H754ceY2knxUzsC0PTdudqX/ffmaDbpgqHJBF+aOHLV+
LSI+ak2fayquvl7MCl2OUvtyCIuHlfRQu8amulJ8mnQa4gbKmp5QtXGkBi+n
z17QmkTelmT1ocvCPNOtB4KpYvwElXS4i+1/H1dqM9aZt1nIll5K7xBaW9FP
g9MiPlonbetH9Rna4wRdF1IqfPymMJwHfsJzHjite1GQRu7mxt8+b1+jx7/M
/uKDRBmtiILvEanh/yP7SawNNZryNEwfG5vm4PNwnK6M3UAaHNUFYhvFaYrx
IIIRIVmKlFdB3J++ME3xecBRB/t32PQUrB5qAS/SB16qeAwLN1p/0rxSchGD
xoAxLOdA3HmY8Qdu8ys5wKZIpFvu4NNn5FAW1OKzfVraPtltDo4dZ5fexolL
36p4GreWQSQuQpnHRFLW/IElRZQ1rzplpnwUD84008uSCEMItFewyUMkgdkn
pJVC6H03/GKYRVdY30qlsA0kufYRR/WqSNgJ/igFYKpd24dTS/2LbG1vZQYP
Nm29aMD9+DfT92DJ7lIMh2daFiei/ZxsaR5iLth8iBAdzLn/3OQecVjq0pHz
6q5tRchHRtulnLn/yZFdcCj3V7d5uA9dlVItTVgMfmvfvig3cfswGlRU5c5j
W/JbZzXF5Q6T0Oe9FWouG9J3S67WGw1P8nnclfxvnsau17EfZp/UQyNuIr0E
ccPF1fQvmSjBBNsn9oZUofME90eeSxeFx6Dwm1f3A7QWwfhrJ4zWNNLxd+Gp
p5fgAfJInh4pw1Sim6mgC3vT38XhmaRVzrWMnNqDWpTFts5nwSzEr0XnXb6S
UlMFwuBXdMzJlZ0EIkCd0ft8DWVOM173e6FQilXorvU50UU7JwjDu2aGEs/p
sIyk9ISRyGUZtSo0z3vK1yFbdChnSSW945cW2VtLHZoTRqW8b5PhZhsC/SfS
kgLxg9tnuU/huxgaW1kjvnQpixGNhK5YKIt9SQ/+TMiGhSm80jvs6DZGmG/K
JMGrf9eWsExLdpOqE9rDyDIyrzsdWwgByh7g8X3RKg0fGQCQ2YinidgE/uRn
ZbyfUztHn+nICasmWRoaDifBAHoRIr2XSh2MDioPyJs2WAoFfp7+i2Hb9JZK
G/VVvhxxGCnicvsg1LvwKGxo/BFGKG6evBmdsQYxAwBYHd1CSW5fiM3VKhwz
oCWs9zhalKovu+pCibS8GY/Iw5p5X5+ZJPVwb1nd6YS/RKzuXeK6l5J7numF
XDplnyVRDQPbX9JO6s+8c/qOtVG7IEtf/1LIYEDT775CxMoUQLVRnQUiv+3y
u7xy909g4bVHn/0Pec9KvKttcAUG0ZZNpOlXagZ7tawpjkRGC5Le1E30DXMA
OLbHE4UWmXSiM7sJIxLXgfCEcnQ7N3L65G97jtyJZ64fw+WyaQ3ntyZpX/l7
7bj0PNvyRQKpiH4tQsq9Gbs/6Ygq6eXu2cfr2JpWdsEjyTp+p7QBpPEqOzMR
Ho97WrafLNdF+hJ7VD3HEs8ZwL7tTqH/DuyK4akIWgAG0KxcNniN5mLk7yH7
5xDF4eQ0sYWvjrgCG267f0kqByGfVXff14A7lM7ryV0vH+ChWlYJUniExbLr
tH9TaDDdUk0E3jVJZH1LIHtQuS/IOk4G2GrcUm5j8XIV9N48JEL/mpIT/ha3
5Y9U3gwnkeO8X3vFCUkhgDTZDnF3jFYMo/HeKJA1h6KcO8gMmqnb18yK5rYI
+BU7QZK2GKGO5HFBvo7X5mH5EmPi/+7juYVkEW79Um2mG3m3dSEYsniazYFp
5rpo5QRMVOpHk7Z3GaVEZTSNIvVgsztOhf47qpyaJoWkHqnTj3WhFSrbcfW4
qJkB56mYZJmbwKt1dDL+xRJLhSQCvgRA6ifMUEzYRTyNfG36FhbcwXHdjnkU
CDjjWtSJZJKmrI9AUfn3VVZBaGxWpBdR/WNWxc0Va+cpa3DgwJFNnOCJu8lK
QHGG06KaTaEq9aXUxqHmv6G+ZmW57jJTFeXCcKGMYoL/Csu5ExNI4egjlWBy
cc/piwMniiJzKolc+9IOzMofYqHFE7E/um8efB10zA3BNIKEk3Aeo3ul5eU2
3g++dACzpf33o90ml0SwJ+/NT025ckl6CxjKTfveT6Ulu+eQ/QdRxdI9QW2p
2RF8DPz/xMjT3r7xGeazihLbLwnZhF9vVa06+BAa6weQyIyWkBOfySiMXVM4
uPGeuiOdra51ZmNva4YqDolBjLz45ZQWh2YXobrFfrvJ6iY58IyJwbgq777J
llGE5bCIxW6t03Lk1C+w/kvkAR/GA18zAb79JXVw0P/yHi0a3mEiY1Zmjg3D
tcNU349S6ow6psp1yTACcu5XhPTGm6Vej83e6Jq5FSMYkkPgDDt4C/7ARakl
uCuT2u9c137okXoDr3ZFNlv7YvSoyabUX4sthzCu1IIaQRRvjYOBFLJNWTJY
D7PURxtYIxFE4dU4nx3EWjlU4GjA7Mdw+2auqYQAM8Gwy3NlgNq6FJvC/IdB
aVR8o9kRunZ4CBu9Db8HSJW2qxhuvgFC+KJvUaWXZx1s4Pjs+sgNP24/wauH
ZT0pEFW5q0behrBTYFkqsKi7X+iv6LIyXunt5w9MFIbWZbHo0xxsklMRlLNj
NW2EY015Q4T3B3HsO0sBT9CNfeVTSpnx/oEEf9tqcTkrF+MELX8IjIHVRpwn
WJVZGJUIg1FGezrhott+tU8+P5PMA07LmWgIPWmeKKa+LLe9OBXj0lbYdIUt
86kgRK/JlsijRsG5NYZDmIBudIbm3//O55gj1addUqAENpr0hRV3dRvqnMHh
eF2T1JBrxoLTopjS16W/7O9vmRky1Qn12AWUHNgb9g3B02m0o+g10ZHspTSS
NMK7V2XrWQ94+TN/L50PGgZyJI0cneNl/+bBO7LqIz6ihZIgI2ojh7vP2pFB
NJ+LvQFqZbI0pRzaSAq/nfPHllH7Qo45q4jEB4jyUTFw7+TW21PcYCG8r390
Wbj0GQi/JR2CNzJbr36TGemtehve3ulaZ6Ww0CoJoapg+fjod0dsEzJgN053
6ykS39cGJ2I6+I9oyLLLDTdK+6NJ3dqLwj4kLx0GET7XpW9dCxGj9yuadSDl
5ALks67kGKlNb5tGGQxi29SG7PTgvzEcPX4awj1U4OwQY01awqHxggtR72eP
C8FBdeu0dMTu9HACsRfsyz9bedp/ftEUzmMSLhRnjRe3FmuAb/bcm9T1Afdo
HplgXrPwQ9Ni9ez1cDSrIyvPRNAY+QyHCGuxAb1SaK8vmYJ+68IQeSklCGFi
s2PvBYUOY0ZiiOneqgTiGpqP2BPXjntoks46TL/rZVSt5JNKrg/hGcVegY58
Y+70zz/X5qLkDavQRFCetiQjFM60UAW9LaND8tK9beqPUMK9XNjHgcxVbnbP
4TwvGhN4xPsNVcSYhRKfgTW+MT5g6zRTRFu0cIySttmQ1q3lZFF9qMya8Kul
+LAnBtnHBkoFhS5+FpkGggoo41CtYy4ObQB2ounxQx6mcz7qE1ObIknvPAC8
fme+3qdYsEVVT/58nGhgvzfWg+RHtmt7+t6vYDB6Wlw6AQbvuQBUqjqtSGZ8
d6SzwT5y9cc1InNquwkGRZSezgzqjzVw6RqAg3U/nhffMf7BsK3jWV2v277w
3asjfTmDBzWY0NclPwsrQ6VHeatejn31mUAbDz+uSXoyT1u/8INLFAraAK97
fTnXkLBC99XM5yopRMHUcGwI0npR8budiVuSK86mLBCKheddN1JeAt8e295t
JNyoj7E1krJOnq2XBrED3xH67pwSXc+qmvThSyTIDnzEDT0cJ9DGqH/S/z0h
N5453zlm43Uplpm/P/ufdk03PqAHFl5YGoqRw186EEnlu5kPRSobl3U9ofUk
wt1SQl1mAZDaohVWY2uoWXx71K/RajFPB0KYtC3tAuuZGD77ZI/aGd6v0NjN
d4p2ycdxRFIzld0mZ5Mvuher3z6SwZRiplUnlqBE1/yGjpgGGBulIMUL+LQx
SF5kolSbtAqcH96ehLwuyGhSKgoGtMH3SATbjMIQy3IMI56Bzg7IEUcVYFC9
JLqQsovQxaCJAbtjENaCt+0XY6G+8VRQer8x3iz/xdhlwsm1hMTx4EI7H19D
cbw5W3meGR3S/Knz1aYD0d8HTbvpjBHql6yZy3he+uo4sD/QlWBl4YoC1ANd
D00jaRQYchY5Lb8tiA5fW5gbj490vr718WLJdQJua9SCaGNblyJBBaTsf2LH
0LCfWyU2YYSWfbgAkiMQ5vHYDkOpwiCOP8+gZW2by0/1DFB2eUyeuHdMd69g
zNeLRV5q7e0+7e2NBpo2okU5zH6if/ZtzuN1kqZpeMlampxeyzunr83Q1pPX
90t3XWBVj0lVWJC9Ia/RrRWe+lHXaMFTFsZvTElBaPoxBD4zxJhEac6iMFKE
CgYAGXknRdn94123HQc3cnQ8i8iCw4zsoqvHTuwrv6LN3CSWZq+noj4i0eJh
rCv88RIvIrFX5Erbm1hPqCfzPiMprZ2+gX4jxIj8zS08XCITzqzwRfM8AwaU
ESCIsUA8RYb4dXTOGtwBTU4iU7aGaU7wuOJBLLGkNBIc7U+DIkdmTDRULeGp
mnvhLYymNnZPA2tPwAYN6xoivHDHr0PqIT9YiPIWvGWUQv5ezVDNy47kgU8f
xqc+7LniZaDdUHkBaljPateP0Zmh6xh6p+htiW7J3yCgqMH9JafYz2xhTq7d
vi2NTIzK6+UasHesxzTlWWaKjXgox9uz3RzGvsoBfnhPAnT7rrKya0hmSnf5
1CxZpPUwQkJxtEv1OGsGxPZS+/YCvHGgs9kmDwgdv1YbWH2rxoA0ag0vFEku
Bo27eeFbuF4gHJlcmXaxRfLWQn23a8Uz1Jx9eqBNhcGVPjUIDT53oj7BN4Jh
iJLdKQE7/n1eEuM6Z7j97G6Hx6+Th58erewcfd1LYoPa3L6Tvy7BYduGdaG7
ABk5akUOXW7lIh1yJn5oYfB5el5XQgztnfbjmpUPL7avwYB75v3bBOq+Uvyl
AiNkb5e5IF/1pbWsMgp1aLSbrWVGW9CNvyeQa0HINlcripLi8yn0QXjTtxRK
BnPYyrZJcEO+ecbaZ1CFlp5U+e3f3y8k01xrpY6eNCwg0xt2uaUdvesJBkxP
ZDi/2L5NpUkC34/0L10y1GTUHeMDkAp6eUiJzeQ5686uL3LR56bG1MPhIyIv
gJQMdZsvyTWVSQQTF71tYSK8cHYvQPgYUfnJBCSDK+IHA4D0U0FWVVrBD30q
VMsu0w1WE8SZ5PgaGY+F2zx8Nzs6ePzYwbSAgLNvB6OkkaTitpGsqjoivt0i
GtHG1kdOAp9o3fR1UGw4DrkC2kRK9pge0v1CnXl9ALaOT/Wpxs0RBTMCUCi6
1BTlZQcxo/3+yuCWaw0S8oWyS3VC4+DmMX26beOpJuaRcnojEiRXc/0Mfd4T
+rkwlWGhJm5rjfYdJtQhs+rWJRSPFr7Yie4nLknpuB6C5wF73xAEVwu2Bt7Y
2S1DPFkoKwCkbhCj56brksedxE+cdce7QML9vXING+Usc2mUPlgaXBjlZFG+
5CbX1CG4ObicS/9FdBZ+XR6UWrZ4EeYfULqa9Xj+l0//C/4yHD9w4TIMblcV
j/ofwHSsbjvJ8cJXu4oGN52MC7vstG2zUyFJCs/8XNDFW/7vP/6MJNCxXZ3O
OlsyNHv7EHHHCmxv4yKZlbY6I9thDnSv0WUExXgcRGDMABHsFaEV50QSsnZ7
ogFrRnwOYSGUO8sjWoKlGY8/za6wO2Bw4QQjH6rPuqmfrf3epCt7B6Gu2zsA
d/I2RJHZcLPtCd/Hw7duw5aSgtPsXArDaZasHgaavLXziQzS4jJbHeUGyuNl
NBBxyOl1NdhI78QSV9/DeQEQDt9ZFY7D2TjN3ac/u8NtIkVTmBJ4RvWrb+iu
pETlGsjRLtPpYwCzIAe4HHpwc971lC6CQ6jqV6P//crHHE9loeBZyEqxgWJb
nq6QiKFIWejJTpDjFXwmeaQ7E5IQr3O5Lj8ZqKA7JRN4OUbczj6Lf2Y1U0+k
nhaWNsJb4GlqP953tfTixcilpUyrO1r0ty0WH4c65k3lP0ByF4yYAI3t8BSZ
JGf6nftrU73l85CoFjexklR+rUSeHmIUUW0rgqhg2NgT8VY3U8bNCzrTnp7Z
HzlvKiaf6gdaq9wW7IYxgAAZqSMeDoTyyAQthwhDd1m6TD+GYqiWK9pRsehz
y5OnZs0ecLPh7+akukrdKPdujkvwDtLtIldmenCKKfjL1XSovY5cq3diSXWi
nskv8YD8yLCKUQNTUTPNcLLefwlkofCxJqDE3ooIrLpZ1osY0K0WwSxiV5qa
eGkeUtCtbv+nitCA/rfAbBtRCD3SKFRY/nM+B7fMmk4/MW8eYyNuAq0IrWPB
PCgGCK+v9PCSGQ10hevXKcB3ytf8mKgBysYg6V0nOhLolY7KEhRl97fW3aTt
lVr+PTey1MkV4SZMmFe0uDS/jt9betcdDsXwM5cmyPaqE2pRTeyXoxK97MK8
TW/0RcRtUHxwq9qzb96yhwDvG4jq0F1A1Cyq7XMvD6p2p259HDLisc9Oxbc3
cUWw+oFxnwjKlPZb5KuEicYbwris5/D6tse1NdNbFQEMqvh+bM8YDiETTb4/
qLMjPgKuRBEQHldpgWfjmsxnOjFU6Sux/8suvFhxZ92yiXEbcKdBdWZ/Bckr
HU9J1/bGSjI7EMijcygQLoxUo+gb73mFqA3y+8aE3nYn7Ywgd/9KFCDzZ9oI
+0AhwyQxqy6BCRmonNvb5ZpBQyiWP/oeYotRkqymNZaBtZxHnR00oKailmAb
aOr9iKl/c6dKi/4Zf+Q9/QzEUY1EY9Q3O45TEH9PkrHuRRQ/Awuh/pwiKrNX
gfQAF2oamEbSvjN5Mifw+2DcBKrG8Oz5TeBArdxi1skosxq/9NRdTBqzV5iO
3PU2VvubId0H9nk7BBzCIIkoLCwevrTq4pVrK78kLKRyCgnkxNi+2FPLaDX0
XiiAY5/pUglRLvhi66b0EkkJH9g0Iv+ts9BhyVQjU/xKRCtdHWpVukCPCCNb
6hnJVQewMvS7/Nqq6+PZ/+GCPVShtNkTgh5wDzcJVhA46nLtthXMfhljMlJk
gE9WuSjZ2id9OkdHkiR9atix2xTVIxuzCJdPKPRApn2c2yhKVcixOcb9HjWY
NwH70TUSk8Rixw2LSHMfL1Y2DAGgzAqM+cwHwuwhfortYkorHeYpZXslaVA8
CVJpdgAxRwKxaIiEvNkw2rmin5l/jJv3Fmic+1aYLoX3Xx08sV3Ai3nIJcy7
S5zEvk+kTuRsGO27GUH/BIzqYQkxlrieFFOA5dzH3WX39EvM8wOlZ7w79XmH
BUewMFvmblLVebW1J0fAkxcMtKljJUB1rllWT9OlaLr4/UfbWwkEkJGC9vt4
QdNsHAWuWbPaUwuLuNrBaPfgEiiFMQmQDa5PYgB7uFSrCSftAawDpnYdW5VS
EjJs1+Vd8fStibdUp84bzL0ZkHHOWKX8hNGzsAJqZN03gxenEB/HxVmN6eGl
qEgBjFOYQFpIuLhEuVPCjFvCOKpRzUDKv9ejJG9aEgMRGzAdVCwAJM5f62NU
gXKrwMj0jEznjaiIMh9bCI816KCamclwhxeu5+TdnNzt4/w1cCwt7N453cQi
BJyvbioyUbGofz9VzEVv+l5S7B/Y3OBQuupoOfR4b+IRMb/dLi2XG1GrBDuL
LLDqlM8LgAEtsp6spbS8KHB7J6Yt1xvURFVKjb7MaOGkBgwK3tEH0YW1/dvX
LbfX0CL0R/DFaI9+bT1TyW8hj/vUwZsq2K246yPHBD/JprJholLaSzQ3AoF2
aV5RrnlOS/ZnEDf38I9HPTzqh5mgkVhD3ema3XLlESsdwqiDBFh+2XTVfkWH
aONRhKJbmVnzgTet6/wTaqej8ouasmNu3DyXta7GzPiDj3ilh9N6hJiJ3nZJ
2wM1wMz8bE1G6hjr8HE9tBZZn02zKJeuKaeZG97+8RDWTYkp6YOnGT7K5u1Z
PfWC6WP5ehMjFmXxZCiA71FpHV4doYKVYohkz4WRjBPzP00E3/1cuGzsGgml
nYYxOQrb/pdXkmpU5cu4Kvj24ckKBWMfZ9zmmyVf7TQGM0Zzym93ZRYf0gz6
KxJuN7mROI106OWJcOxruxkGs/j6PoZljveh5WwDyj6ruXcEyJm6wWmgSZSe
OyhXqeb6mqY32zophGbETH98gKpjzDMGkQfvsm0/a9NO8znAbX5Lxb/Vlc6Q
3ZoQCmDKB4dpIM1dJbCYIIN0o9c5vs8Xv5WbJ4bkgxYzViWpuJcHNqq+lshS
tUkGJz+nOSAF4t592G25Qyvuc14rjQ0mpYTvKV8vtfFcIcft0aOy45F9ZEyM
unIJ7LYffgLTWsplgpahTgZCZPiQyvpx2qqLEPPbp1NDmsmhGyfQ8SgWe7Qz
MRpq5Fu1bsZ2JYv9cdtYKjhMxJkFhZKZE3vhPiNCLjX5bSzMJHOuMDRhmd8o
7PgVvFMmpD7s6YR3CwjS+87Mbf/T7WsW4AybqicTj574M80yiSH87zuCHrPg
0s0kGeH6TQBRPMt/KSwGgVaMW3MMu9ZE/lXHq0vliT8hjmMHFbXW3Dx6vy39
0ToAqa7aEUqsJfALXO/QMvHJKmLTnE7rcd4+1leOwfLKHgYpbUqTvAsahVLj
Bph6w+elrsLCtk/0ZJDf/0sQEjdV7H8Z9aDgkQ/UAGr6V7hiH/bM6GbHkjHE
n4GVFDXhLMkCJv5Ao23nP1OVNjaDc6JGkmw+83pkTTzXiB39Qs2Im6OXQXZU
eZDMS7+vgeNObdOeH3EeE85ZY8od662sAvme30uK6abzDJdEKQbbDv6dNoTu
zmb1khf6mQN3EMxFJf6sSRUhABItZ+KYM+7QB0Af8BzQg3ad11u5FMkUetzl
LeV5SojfvL2yfpbfmF1BmVgVp0drcFTLqjwh9c14fyp0TmwPPZxfH0aFHP/e
L9bnqxGIVKr1wurXCcWQAB3LVRpbtZJtOxesn0N+rzzsUV4z3KoPNG6gFj1F
jruBNXU5Vx+Q9ygkG42SYc/9TsTFlR/jzQyvb+zHlESurfBBmSPzedor14AE
gJBiR6KR8M1g39zA5RORt0ErtgPsoPDSQoUWeB/f8ATkF7MBwgeNq2E7gIil
ckhGM2xzB1czcNnpzBc6fmdTEUAFZLZOp7tGx8zpKmLG6vqUVtE93weyJ4MF
+cw1FHVyWvtwwfTd7g4UdqrquvaqOz7T12G0cZkeqe46m85RVFEWSUR8HvET
WsteWZ6oPla/PWjkB/Rttnu+3+J+85L6w1aysSvk4MlB4kpeEOf9YTg6d61k
FRZpuYSoC00Y70od3xjaXL4CgIH5I2lAoGA/EDpYKsuyD/76Y69bPU68xkEC
d8UiOMKr98Fuu6Ho2hkOlGvalOFU20Kkf7Lw4eDMvZ86zBymQA1BYSRHePz0
cVb+/YaxX18nTWoAPP3Kb9/JZxxFBSQ0nDU1PLYmJhFjeY+wuRumD552HNsT
wiyqbgTpuf1qFwA2Qfzehzleyf4iJqPgchImGGVuiIxYD/2S97OzRaDuNKlj
LyfDyRwAKnwoITIZ9bnuFzlYkajPSQB8MhvGBsToY5Vmxa1UDKlDRG/e3Yso
FoOMN68kbmbZqtcyfl7xxRsgJA0TORIexBHoaCKtsF2AnDsG+EGaGp7KDB35
HjU8egWLjD+pCRS6af/01qcPa50d8LDo6X0tS9CzqswQcoFE9j8h/pJPq60S
q5Q7bJuvhh7X9UN9BCDNhLQhuNOsyxxM+QNdVoy0VR1QcFRh13S08klEUCjd
LGTzeniEXD7iqsDHduL02f/Yr99XLxtCPXNvVEE9Cdi8GgJseH3u02cTpvR8
Taa4IRvO+PLn4f50zP+5gfR5pbV4l+Xdi7o7QjH3QZCBi/AcVYfqKHzHyHcg
2ROUkJGqM1Rt5xcC/z/XiSOOhXuE8sNCVVH9FcnhLQ08JjBvVIuwjsvoCHIj
BS+QWsFFF611d3hD4Eo8IdaZE0mYuDBzZ1KQW5ywcN7JF973ZuyXavnubi7h
gTUToyoHbDsVas3AXGsrhhCCOhWYpT0KFJw4cCaV5o1WZAZDmUB+CEr8FiDr
Nb9kvH7KGhdO16WnZdS7979VqSzUmGuspWVmdEyVvnKvKfzq2ZX0ICD34gbL
NV11EXtdyBQQd/Gk2BWRocnvbdF0JytIEjfhwK3ZhjqpqkpNmA+YV02SFbLf
GU5LtvqIenirkX8aJvdDIu+sSQ6PVVBKcOkxRUaYL74Juh9paMkxR5XHzpr2
oZQ+k7JYoVXPT9H6sHrqxlEnmRrtppxs1IGHwvN/6o2PvDDeswJkbzeiE3My
NYxggo5nWdSrlXB0AZWelnVcune9+37IOb10rnKGksnD0VIcqAX9NVAOnImD
iw4VPX7qsjVN+a5MlLg87QmeLQoc8wCk8UWO42udhgdYTbgtTQb94TfpR02g
3eSQAY+BUMjzEPdK0y5pUD498B8Ch9+erqaIhPpICfyd9PQyCOrjrrUE0N+9
uZXdBy6OtP6hv7QTO1hDH8xss+08L1Tcu3/en/shB6QK8yu3jY6zOBEPoiAI
y6yyqGgMzKKgxUlXh4dRcjbXealDFkjI9cb+g+ZRfvE8wi1mXwjntMfzKcBs
Fak+iBdiHCGMy4GvhkmbPHWDK+i74jkLBuFer/SkCPGLmeppWmQkAUfVV3K+
oYA1oYhACls4yCw6sd5jxp+5JJpsWgB7GX4diYuL22gvHiuGiSL3UtDp+fBp
/G9R7yc5GvOmgCV3c2lhFYzrHq8oPpzC+tBYTnptgR9KHMO4tn6RikTnXSO2
o1tm/cCGeoCPZVpwMqiYQtuLH/5S8Pw0iiCs6q0hPf4uARygD40FTeWF6Aon
5JSHKvBaFGvMtiyP28CMskx2y7+OFMhuDhNoiJjHhOlDJddJq5ixuUWqFg1b
NrAkRK3Q853EkhCNfFwZ3c+iO/46VlObCAA4D60wA8NVeHRww8VLCVdgfnT8
pSo4+wF/3ltD4KX2yCJFx1EThmdzgg4LYlHsDjncF+/hfAuejp4fCBGUfQgv
4eXfknvCQH74ECREbm0lHYjddGDfBAeNBkpLpQ+SgafaFF9VAlScjNnfmQ+q
y8/WJtwz4NiCEOYRHdeomD0FXxuEInfxWL/qP++U9UCQYKTodgxkzpcudC7p
91H/7C8naqGYr2+V+TXaYqYfAyymplCVARH5z9KEZwtewxEmqvBFD+jKH6Zq
wlQg6rULsglUqX/5pLPsQ0vRIt36373Ue2d7bMKC+s+W7K0Mlx+lyPURcDMN
fp0dVaDCVC3oNpogVEZE3ZWLzO73h6I0bRQwBzKg4URm+UyMBXubN/KpyFUx
bNs/CbB3hOYTv4aPLGWd+ZnqDZNNP88nsriGpNiq26yN/HorL7vsk7Mj6GcI
qBinKlV7W2ITvCBsL8XzhYjgddyivcIuKWDPAuQSx1tR1WCnKlj7x2OaPwGf
lGvlxzyMxOOUlTuddlpChxRIiK4TFP4CziFgXwbaEk34HG8Uo68Vzr2ptBqq
TnY8UlR2dZtDMa5b59ReYCbUv7FyTWAnJTJRDPm90G3hoWRZy74SZJlOHaBz
Duo2AlABcoVYMQgw79NxWSbyyCeCsELHdQzBBprpRgTOTFuiC2RY9pScjN3T
RUrCBSpWYcfBeM8LKvXHdHpjH5RY59gphhHkb2ezsLGGN2tms/I1ZFE1hOnR
sqr+9b9gRpSQRpIliVSW1d85t75orz6OWHDCDnnu5CaBYDrq1s3adm6SIwnG
Sjw1IzNsG3mONe4AfOLr0EF50jbHSsKtoSMHxroB79+lG9X9JjstQ5XEPNn6
CFiQOfjUAc8gDUJ/hxs9lil8EzMe78iNoOMYZVgfI0s+vk94OmtYllqPCVWb
taoiYraGfAWeR5IKA38voHQP+b3q881WAKks/0vXVgvcJiq6ZEOLcldZ7wTZ
0UQoH215FRnZgej9PBGhHwZe4TJUHB506BMWqYkgpkdKqxTbViWk5R0vP99J
fgimko9As1Kgf2jS17Pc09yCJH2J9L7dbKgI1EY+si5uUZt8SaK18BJd9CFQ
KYd7U19ULNIU8EcDNlFLbxRUsIKEP1ePVfNJMUolcVkzGsa8zR6kRMW1Ue59
FNsUO+wsTtkxv8smhdbFd4X0enMLNtP22aCeRtGWuW+F1kD1fQ1OZPjNUVd7
qceC59X8De/4E4syMHDIxs8x1GEPueinl56Q1ZAVUAWLf8KrVwHudHlMR1AL
CDEZsUsSwzvv20yDJhj+b3hiMqOaRV17UGWAT3X6srsTP4Snv7bYxW0zficn
gvDB5pie/uhPztLexUrnR+p7UuTo75USr3c/GPhZUdZ2vvq/J85qyPax7Cls
3DQwAxT713pl8fnR2Np2A+SutXRc+hdQrlkQtIG3/inZD3wDUQH+9iwh1361
CtDtzQqndTBvSX3Ig4YAYSxvSJW5Auh2XQ0AoKl8FrvJBGUQJnqAUFVxoYAU
zU7ZYnVQxDY0yTbjS4Fp6NwxyfI/UIrl4jbWZANNcs4PAhyuOib0JVMU4Fqz
rZ9hH+xFA0d0fl/nuXx0XweW/ShEoi3GMQPsXLJnYzeEI2ARV9pZ02e3t+JW
gYtaEadwRQgOqHDfT4h6KysaMglFnMMfh7ScRUZeu47CzBrY5TBjgzP/+kcl
WpOv3x/K/mPNboawLagngiWKaQ3kKAk/0c5zSUTcXt2FGb93NbbQgf/U8utI
XKIU8JawdkO9PFngK/Js7/VPghZy4EF5cjGKL014SFVhD+guzX8+9PVRe0Vv
eT4YgYFMnwEhE4yU+6CcSCJ8/Zbdw3BJ6MosAc8PxXidkp72bJw+6Of5/kI2
ZtzFKhc9+iY51aCXKBaDwByxyo1v2eDoiNvnGq1CztOrkEpMBuIQtyvk6VFK
nq/q5pKxvZO2ut7wv9TNeQYgakqNYFFicwieXP8rifxIJHl1nGivxAVFEYZ4
zGGib7fTN7xErTBeVG4HMnfrLJMl8Ag3rnGX8/jkd68ZtTN5uHue59nfCbrd
cmCR8kxE3G8qWdWVMX+nuuSpi/mx0l9ukvnogSy9bArErtbTqNojztioXLtC
yNVFSO3ksY2dJsBTjLn4BRZD8jzx8BFLC2DVKo5FpS8HMC/qwSZEnCFwIehz
+pgskXX0rPEWtfPRea1lANdh2Nj5H/R/KOMXT7P6X3O8kFk/8x5UKwfA7bQo
TavpWXvXWYgNdpWL9+Su6IsT2hvgBqbwn3Yf+NW9O62MKvqjPrF4yy05u558
xhxjHp5ML6VeX5sS+QwMee6ylf69jujlLWJPPI723FsjuWxzd7yH9uu7YCY5
aulkfpwuwS+Uc4pzuqg9aT8Cn0RyLk1+57IcOK+gEEn6fBdBG/sMithnop5Q
lFdC8v/Z1tNH368ZqQYfBWZNBvtvAvOi+S1cZqvPAsTgBqGm/GIM1bZ1gcbC
ktuJ6NQuUH4TD8eFz623hAyRLyOriZXaIgHfqvVAMHvZqIZ/x5U8aLtUzmNT
ASNtGtg9/KRuL6mYyML0pbkRy9WJlPPjh2YuDRtR1/TmGUAPBZqQsFyM3PWp
WdzKV6B7PuOVOhLBb3PnZbbcbvxW4glZAeNf1GkKRov1u4mIryqQSHXAAhZO
aZG4fYPAeI9xb3Mj1PmrwDlNU4GlIDOuGJGfUwcG46MrJWfKHf9VXRywJnal
w1OIMMsgDZoylyo0rLYQo+y4COWGW3o+4tBacS6BxPiCIIu/ShwNvuyASOWA
7DOTyPFwubfpCiAIeEJQT/ywQaxwKIYUkutijTxe5diED0XEFtWH56pLim60
DKLbjKnyjcOUAEAZcyZ76ROzzNqeF5ClKbAOf71GGNyZZeQgIhQgakZboPM+
wtrMBY+wShrbOKU7fO298V3+N57dpGoy/ppCio0N44UkDZfVa6UiZf4Rouoq
nDMn2CEj35FWAR85TJRdCC3IQGCiyMbbmabVSFTqd9oA/U29gR8YyH9ZJTp1
5ooRUEilce7+0yKO3kH6Z4RXorlWUCUINHOPzGKgv8f3M81DaOSheKL1C4fn
r+8c65k40qUjyfIvRc3oGHK5GYHZbHo8jHz525V3JvJK9Edt5y89aVYWluTj
qUd8VqtAdF6KMNfvhKLLXLCSfLhRCHINJpR6BSl4HabWQoIhXxk1bx24wCPP
ZzaYSpqtpx0O4xXwu+XHkzZ2i+NbZG5YmSopF7JZwoqfDNMuclwOLBtHJAWt
2X2nADRJqtud0lInu/zSIL/b6XufFEaTvfjdtVR8t9GkhWpOEcwHgM2Oo3LH
dU7c4F4HqiVvG1nqhRBORznc7WMtWBJL4u4OoGo6CWNcaKyPvd8HAiPyyr81
tyXYWhxswmojJnv0Fn3Z7fwKA3CTTF9F+KLNCjyonojVcpLZjnf9+gxWIHYi
5DwGwk5YeapzvoklDIehTKpgl7JraoPAOKz/gJ7wQZO3hb0vFoIVsoNbYMA6
QA17en7FM8729htz32c2347fkmd7Ly7w6eQek1M9v9N0wBkvjsH4snAoD/h1
/Qx9XYmP6Dt3xxlXIAw0M30oNHgw6upo8ayJMdlSHCgbyF5oQbbro8r6aUeR
Z47rmbQReJAdbxZ3vSkW7NGbPEQoNog0HgRM7n4fU/N7UOpi0wLk7WHOjssE
F1blRpypLMy+48YDwoJ/WLDPN4FC56MOgNxIE+gcoH9kDKPhy7bnGDiMoQ1N
8F5aSke9yu34KAQ2NYBFSyp66E/KHsBXaDTKksradkJdPXEzWQKjImkCnGXc
LcCrlMbRES3lzLGu4LEpV3kb8rmDWJHJfWEW88X69O8aKGZO0BBPQ2ZCu3MW
EbNtlaZROUI5uKFJKjorGfxX+DtZdLwRqNvfQWgmDgmA4Uq4qUhQgi5jLA6S
cnp7JZg+xwKumPP+/d0skAYd50bTtWDMRLK7ul1yRB9MAJ3tkWkhY5BMPkVQ
DyPs9NFiKnWnlih+k6PY/wJEEi0HqLZKCsPVMeGSVF/eQ6W6826ELiCwLLtB
sBFaOc1g/BC5IycCNfT3xpgjMEkpgnOEcDjUgximJH/ZJMuarW+uW4Oe0TgF
Kk91XAzHUIrNH+5mE0gFufolshPABKAxT7Wd/sSVHVdmbJLpxxC/OmjyViu1
dUC7eQ/WM/7YEm6yMISTGtV9yMDwWfAyFrfhSbFF+UiIhVYIhBGGRm0k90wE
gwOq4aHBwB2EZuyhBIbuliutCYFf0bcBbfVz9JsE+aEdVBq9Vii9BR4upOGX
7MynFY5gGHDujYqaNn9ADyzBleMcffuuY92EjMfS/VfPS+6JnC6iF8a5pQFo
2CedX9Bism+xufPWqLH248O4O83MdkU2rnIHxr1Eo67KsPwpYayIJEgY9nN/
sRWVNqQJ/GOK+Ju5whCwrBeCVXWJcnFPYkOhBPb5IZyf+ChuKWEaeFETz4Ht
r6OLa+as7TL6Nh3c4kYLDCYBt8s9g/fW1Y/S31zNUu0Lodrwlj0BiZEcfL3/
rtMbd4WA/6IxxF1NgT5rC8fLDX/QXIbT2+mlHZ9sw4knTO9VzaNuAUDc4iY6
54Vzy1Y4qJP8K9PXv1Qnca96rRsqUhm+Rpl8jHmgSDt0JqUD/xqNFolx7ULp
lvBCPs2RFzSAwmFHCC1fgcpwtBiJrXFX2kMiXXBFVOz6Lqo1XYNfRsVcZGe3
Ud+MY2dRhX1upzLr9Jfi8xkQJnpaChYK6fSMtK7oqe9Q0wqPnv2rGFwrNcPT
ZpF2eKm/D8ql9nf6SJbh0NOGGWXKQ/Th0cesk64PyeBxW4X8dVyAFp9yG7mt
ZF7VYwGpXeAoUDOpEGuebZJGZJOGzBGs+nfE04GPMx9mWdRHagA9mno8QAx/
kEYKBElhNVPpINuEQFON0x0ffpSknA4x+8oIJ7QcxdrVnS+npIvi4WC2lnY9
2bWPdGUrScIGcJIEnE4vximzcz2SAXudrtTBf4g01kijMFG4UMv4y1L/w09F
ox6I5jtTec2LRDxJKGX5KSmmgN/dIeWDwYSNuVvu1C1ac5ACJEsmQS0opCoL
7aeSTEJD+aeK6FGKPKIlrCOMGSpXEe789vZ7CEOOnkwVs8xjebOfDSm6UNdW
uBuhF73yEBJffFSWnacPY3CDKw8N77BFOh/xx2hxIF9dQxBo8wL/hbINRRFt
p1KndyfSm+sF9EMYq7Jb+b2nJ/iLU1FAgJCK7B3jrfopLtHZRYv7qMpqSU+s
y8O983lQBXD5JqcWSdmwufrVclCDIPpByKep16UTtG/h4ZItT1Q1RNAwMFsi
Z0fPGOcDEUh16E+0v5JClHclE4UVfcgTJo7qdMWVUR0aiK24XnHk6cRXncr3
9TqAxtOiO275wLfL0ZyxePzX3ESqiLzgugFFaliHhwIEzn3XGJYFLLKAlRGS
7VlIl2TtW3Ke9/xvHOcV+S9oDS6jdEPW/zH5QHaJdb17+k4WJJDig8lZTTSV
QGCANoJVQe2UbRjg0/WYhWEV0psvj+9NO0CkH9haF2QaU6fwifbK61XwYHo4
ZDBTYIesgjmN0Mif2X3+Kf6qb8D4qZtRBZuDpS7Jccpkp/zkfE92w2m9/LvN
nNHgfDfBkR5eJnO5xh/U4vLdSr690p31OhzgcamtEb3vGKZSVD60GHrL+Vm1
TiaVxYZ3MZy1j4PGuIUKyG9MvtXnxB98n84mAtLgbBHJPNgZMFwseYAAJUBR
SvRGUo5nvr4vV/71IL/mWgf8AwWDHSe54MECSazgZq/0Qx6UqxBHnLuCeAhC
ejQ+1xgsfKdVlbDHNIvGYpBOrQO2yujVsxzz/CxhGMrR1tFZP8LdLm4mkNFm
bVbALxQ7FHBarqynwSYbCN4M7GE5UjZVaBGxUrtCxCLLiF5bH7c97Tc5TNUq
7/Cojdpx4Dicej2VgxJF0wO5HtrIqs9myPcb5+8sZY0NdoldnWtkNnvcKGXW
hGLZRoKd3jxN9Tr8bgolk2yL6uHwlOrGdGBjaPm+etGJKSzARFnKK+OoZcam
wnMlOmSf64AkCU9uA/ZwY3hFdBBqYUp+BfwinSLMxYw42T4GgFIYF7YzANEE
zgHrvvDiiIMff1fkphS67ALsBpNejKUf3OF20+WUbriTmHnH1/60CTSGbF00
pKOkFYON8ReH7in0NAL/GuALZAO+G5rkKciSBwlieWkBkI6A6I1ns/4xWpck
MKcEkcEpa41cx0Lxaz9j9xHY7eU/GHbOInz1P9ydnEYy0ezJnhbEWOebfiv/
KKmr74YKBU87zsNU0ej0XUi1QheGyLNtMpWs8KIfJu/lklAKXMiyPQp336pm
CgLuNX/PXhDETPwHQl5c/rXy3MwnnXM+VofR6dXnz2DUbwlCOw+pg2yYVRMY
rqWGjGadoT7ODmAov8w5qbdNabD7TDexbk7Sak6MNbX/AdEREpGE5cLU/DVn
53QhrM3WeFB70Ug4NeCK1k8dtzGv121jF8jllkBzV+Ypo6jTKv5kCQKv7kPu
FAON/HzdS+MCFm6xMVrjcrCXqvjEIqt0iEBNpWqfM/+Yx+PbUGZDlGPH4Sm6
OdfnpPGB3SGRfs6dYS0GcvUs8DbjR21YaT+HGPzvkhj59Q5Wi2iHsdKLDjyf
+Pquwc1KgMVnbG1P99nzLvRDQTs5B6ScIcytS8IK1tLQXCuIb4BU5viv8Tif
fQDBGUKZ1fTc2dU+CceXjkGaT/kW5Pdpew6z3PV7JxI7LtmX1BKQrC9kB4WB
Gy7jiUeFlC+i6mSG+7RLxewp7yP2oHSAu196FbAayuRHpak/RRTf1USfMGSo
Yz3QsbtNrIKtbKXHrQt+sigjJZFckizJdP4jX/Gs/2N66cNx45ltmZQ9Uu18
/ukXxOCbSugOS0u5GpsxeGMJ4qPrLwmTGtSCxiIc2tzaXI6G74ezz6iHSYIS
4SF0LXd/pOA2sLvasgNNe5dbpJAKdfAUNS7qO0laa7wjCNb8Xnh8kUKf/Io5
HQMQWERxg9Fv9FxizFtcCJ+HWCxoP5qsY9iwvbMYMr1ZQDu+zdTCPju67uuL
7CkXWFXoC5F3qE6+9PUHSndWmStKZbqweAkEWVcfOT5b3fbV+TdyAZHymeuY
KrEOcthcHQz4urqZHzXU2wbeOO2as7i+a9xb6mlMFV2JiNlWnQPejfIMaabZ
p4egbCWzhj/l4LuTK54o/JSjci690ZfOHjNlTTLcqvUDJqHjTFdiQTtqO97Q
BT95XrraHpNwQVVAkdtYZCrrt3Xm0PZRyoNXwsxWOTXOVkRelCEf3OyFJG9L
70K5VpZXGSuP7fG9m2qzXOPSc6gr+5psitIofViBPAdHu6oi+T0KzR9egIEg
pYN4DToOdSFhtYYhSrcLic/UUJb82rDMEq2Id6mxJRD9LyaNWdEgiZS61VfU
ebGIGt3MykCDeNjOGrGMsy5s4H6t7ePRX5iLo9iLKNM9yDB59v8wDowtHNC+
KKylbEbiC0E1hlgvXrDVKOMq4QUF478pvCLIfYqb6Iu/0/b9SxnL2ngxfDq6
EOz8TLMvacq6Rmo8xoZdZCseR5rkt6MdyOSmSGaj1Yj/yxDnN4TEtV/SQ/uD
c1O6vF7t1x9kVkfkQMiZXYKDGXdj9IEtaB+oGVNX2ELqCW1OBF+nAKV1P0SU
sM5BoStzehH+t+8yNjGHf+xLm+xilfbA8MOH/lBpsUimIOIyF384i3OKX9ct
7RQ+8uN+PKLYcp0vB36RmeTIFxGuZ4Qu+vrObUQoT4NdACCZ+4EL1OI7NgNz
g0l0AVOphME2xQyHL9ianwPbOEz9GYcJ42crIN1kpSuBaMuHRhQv59mqeuKO
S3uZKjavndlNcuwD/NkBZ5khFH3RQp+zZNVL/S1VLdG8EMSgyottCbCZY+B6
Uzeq8SZmZ/xusM7d5lDneNfPhMYy4nd1dbLxnOi3nXFwjd0t+c5YK7iKLmmF
w4q50xC9kfkuSLyUt2+KVNULVMfx6+jipurOXyN+ZQPBbqNuSFHhtDVnM0tk
9EHP2wErnfLksGJY73qQv3aIo9fWbxRUh98g3X7G2XrBj+1BskivATdcbO9c
hPSKS/DkvQ+Sy8x6YN/bL9xt9X+aYj2gQroBBiTf5SKx3BrIjeol/SM/q+qz
h5c+RXX8WHt3sk2nKPXvKG23ZkFmGrv7C6NQsOi4q1m8leoyH8G2+fqNV14m
jgrUkm6FRysLg5/bYlgfQ5ErxnoR/qPgGA/OB5lz9wKMZHJKVtGi/hNR/eB7
3vsrU8ze+TQTF1NH0jONPlmTUoFMOSd5p6FsvElJPWnhQx/LAAe9tL3oNelu
2vxZiqRBr5NlvZuK7vmUe7iZ3v6R2pL8twm6pnVE0l3afalCyuLboDxDc+hl
28yZ+Fs0pY9KNGbebFDRgHErqOQ0VyP92quoqIqdpPLrojPVRgxUNawtKd/s
ZQ64QnVKjkIp4lnokxnFmTSDEHSfVENVtHt/C8cGpBa/Qum1X0lLrHN5+9jo
AaZHsval0L+V4wg8ufzGp03/7griSfkcx8v6ols0BzsYZKwpNk2vgSNPF4Jz
Q17W5GaePC4V/LddrTlR7rpRrqSW7onACxg5FNqCy6hh4hv2uSsKeb5zmhQT
ohBmsFW0/roZd1/yX6I9jx09FEDqzi8gQYNybQBmbugcy0GXTBWhjESj392y
4f8WtwWEIQAqoQJMyvxkmJXjS7KI3UFneYdv3Bnp8JLXZdVq2kty46mvn+tu
K5nObZy/8VVdoXQUeGmsDIia5SjVZ3tp/12b6vcwTZQcuAuYXaukGBsQCwne
4bDlfajKK/balklGRUDRCwMHerjWzN9ZpqPAZaGXqw8BjzDgCKox4eQ4vEjp
2dje80CfUfAcbPtvvDrCrHMPtzE+RBKrkEK947yqREQBudgNmLwyyUUx/1iJ
ZHIdmUJKXY2YLA42dbjqHEIXPOg/BBrYxZh8/eL9JkmJKGxh2Uz2SXNdoeEK
v5D+m/r1bT/EIRiaK4JSDdznyDjvduTY5k3U2BRxHHlGGawlcXfNu7Ze1nEu
mJVePLM78rxCLxUspJ5QyB2ZNrwUfQw/Acm+v6StJUw1zAYmXEcb2UMGws1G
WAGO9R9UC2TwoK9DZmBdXw5aze3kV4G9otqawjUlh016WaEFsA6mNbM6/qGz
R0P6WuUrLtQlevFpJX7UfdrhwL9DgQsMSmqTR3xXcjDk27Zn5/+RS7UbYUFr
5EbjBweAgA/vU/Wbdao6pB6Mbo0Y+/555Pogj44h4605rDkUscaUh/R8pEZA
acdXnIFm5Y94W9k1uUnz+rYr6MRDqbSoStpQHB0nUJ6lUHYGkhu/EFySuL/n
mNci3XN8FZRVNVVfL1XNZIH5JGhSgdbOa/OIjrqGODU4E6iPGsl53R+h03XO
SIan8vacC+YOUM2yUBXJ4gFjvsLI09rseVR5529qSoWd1eNK1mT7fSCORu1J
2DXDvMhlTGKFY/OEbFz3JCyIP7SUFDWJQH0634XYBFuRkB94mXeQSr4m1P4U
W6dYJ7/tjmDV0vaH1l7bPu2xZ++H+T1BQntzsrePCkDwfvbJSxEafehCmr0T
w+VjY4ZHt2UVkivIe/TbE2GuWgHL6C4ydd3rmd0EylzD7NxRYTlT83GRAsHV
KZ4B49+ngejH0+gZjNvSnEsCd8w3GJk1fiuB5SKFNcNB6E6JUN3jPLPbRb1P
BCXTHl4tOz1VBKKSA+lExPMJCAteaF2ymXZ2rU4pyFm4+KexqgIlrGhj6KR0
05AjrB0tjO7BnFP5YmRhhJydL14aCJpjGBwt7o/TgvaD0b3iaZ6vpkSHQg+P
y+RRoarDBL4yslkGjvwFtTBEFHqZPLU4tO4f9nMoAFoCefYZ96elkZYBUPgN
6QxzC4X9cIN/gaIKU6sHuPT+ivQA81IxmUFYtHL+1zDj2qZjk3DV0+CgUQb9
sk+LeirR4L9Bm3dbrA/wl0Wh6UOotP0TWMrWzyElG7CF0lFcKwFNw409Faeh
5CwKQTUQG6AEw/MPfwpGPNQsOH4Psl88jPoy6hjCTZ8lDDpeNo9yYFfH757p
fkkU6/6FoJ420oKqAY00m0iaoQccQUfS0B1SqzbZ+FQFUFp3yXfTwtij/vUG
AEv2tN/4w3p7YjsPO1m6792msPCwiASJ1SxJ1SrzdMVHw9fPyI4RU7/CiPzA
DQdEaPsc1lIHkr6aD/qwfgY4ArFwvqgkAnu2NNuCajsIzYBkyvxZJxd7CxlV
rHF3yDXxbH81h+JiQBtPA4YoIWSQokugTHJnXSHaZrSK9rHXCJ7/nQ7pCqV8
xSELwcFIC7+9paScx6X9kPMOvff+0cNygVwgqtrQJeK7/xF1FYF3H/byIryb
1I1n7mllBs3DYT9jFHLrPufX9BpO8B0CS6voPJvEFvjCWflNhWLpDMXHeAPD
LTGZnX7+1bh9A3pNPxPWwvlR1iYlDzgY7nWLE2z1Qj6Vq8ivug/Jx/as1yNF
GllZkYO0FLPuwWtTdOdLa+jTlhbvqWkCgLYKcwB5ChY1D8jq2/wWcgMFAqJX
7CriZducZTw6dGr6AGvTo6Zerg6+60p+VcijvSUyqBCqiaMU8EpVcPhRu+WE
Jip38z5DQ/oUQ487xFeMDT8jSwmLkv8pjonB0QQig914v9bnFX4IH0V+v8xt
kExC+U2V8E5kfWRxFVw/rjZdG3BSoifm1JZzbcjxIU4pRqsKyAMXV5ycRI7q
bhLF1W/4GUwaq+pfcR1Avq0S5B2GpUb68Pv2SFg29HhjU2L1kclKXnKuOJy7
9J7jUcaJbfMkboWztsR+0BH/kflLCvFRjvi+aZPf3go+PFEG7a9oJZICwY2f
V1bloR6PGmJ66ziVNDOHLlHUnU1804O3wbSAIew48iUrEB9SSThL4h2VqERb
6fks6GbJ5Rp0J/XoqGwNwJ3wXjeo5xrN2ZGyTPcmXA/8iVCe4LaFtyTArHI/
f1skEsN04uCABY4hkyXO3T2nOYYTEJ9QJMFrhN0P2hshVukXXlMUs/3toQ+n
JxCoezKtLYxhXSClvfqINCsBpxAvm4Gi4qOUxcfyvleB1Kpt5oW7fEcwTK2w
XemG32qc4Mpw9XVyRCoXh7m7hn4NMXfuJ1/tfilClagttb2b/yJS0mkE9aaO
JFoZOfQaCZpgCe1Kjp3FfTEo3596tpVo12vLB0z5dwYieWTLA8fRWGOkUzEa
n2wbUY/K6nJn0ZneexEZgDcsaDfYPsh9uICC8FpHUUmQCj1vi4JLHdkChnLf
Q2QuoMtAKLpmaGU0BkzZ5kB4CMOfoIoQfXWj0UR/hl8tgoUhq0/4TyWjJMh/
48uzaqUIJnjMp6eUU1duLetwKOLOmoizgeoLvnV6ZW6Rhg4aFhwGRBNB7Rf8
ugB+rpziVtJ1Nw3FuQi3NpZRpM22BSa8rUPyFVJztmGGu/MT3dXzXNhFEzo5
m+X6BPB9eXW/ocBxN68eH6YwTfsqRFSBmofM8OodQPOM+0cItyUv1vw/pn4e
S+Dkw+zghGpVVlHeznfBrycB+BaL/+bCmBlLMGxq7c5lE5vatTAIAzn39xY9
5N+2n6l17hxztnYGckAVP/fHQTf0VpafvtX0uYwG3ZtqzBliBJsJdBhJYKRb
jLWRHMVotyerMvnyz5/aBIY6FBj6cImybQvZEd8pGu1sIemihJqdvz8fJgE9
0qArlzYCqbOGdQJ17i8oGfH5fJXqyHm93Op5cQNtWtcXYyoEBx0bcA7G8JDX
2JpqQuItui4hbRWZyksWEjmgvJ4aZTyX09yIE4ZBRpOn3iVLGDqZCW5bI+10
2u5fo1egT3NkfJIgxE+wze946Mj/oVPEr+bIvAGp1++qQmIrBBtcB4zIecr8
ur2J1fAF+6Xeqmu2sOD7rIUTVAgCfBe15mQFe1Usf7u7Lhp8t8o32JuVe5zS
Bv3008k3iZEUkRYtwTXrciRpHhXznDJazGh/tPE9NGb2Tgk57FX1J0udO6St
2Gqfcr/8kflIbhSdGot7UFnme4VznF62rx8hM/U9Lc69nJI94d7UM6mHiznn
F1rK4/iYcHUQIVZxbVUjlZQH3E2II+fgfwlpXDb7MvDzXeOPvHMyia4DWXhu
dOaldSE+fVp6ln6uhHfOg7b2NQFtPow90fjXdXyK/1gCzb3Bon5uiD31x7PU
FgcMvX9iZe5fY7QPiMW/UTTnPCAVBZw05HBwOVLov26GbQUb4J9Bzkzaj+iT
aiS8YVzY0vCMwHyi7+Sgqe/85Pkyr2VBDr8KeckKGoyJZKlLB6XalB0bXkn0
DIY29QapwhyW4zFVdA9VchiFts+3ljjSk7F3Z+9SDrf+pRpgOlA0vV4YdgZs
k9qddUNE1/7TaYrMXPXHKlZP4cTseia5lGTeghFEbdLayg80sLhgIZMYbG4H
+UIFSxT+SIryliXhla47LcZoAurZya1zQVcOHkSGCV+EV1DlkVjCjLjv9Q+L
DY3S74/X0qmviRDXamlk4lc2RHajzREZ2uoL3E3rWx7kwx5Z4Mlp48j0xlvh
7O021pZ51i40WL9x/Jxvuy5vRvuR8BZ5pdcKz3SH57OfPv8eJYT9EcCMIsET
op2ZqNSkPG4b4a03VS6HNeYONvTS/Ppspo7IPCe/iH7URrDqLKL0hFB6f2WV
7e2pjDFRjYhJTy+cVkykVm+zuKbDRgccfaInsLOz6UsYMBZqSoZSK3NP8Mxq
iAaqhxR60Ly2VqOJURA0ifklfmWF/vfIPYji1CJlFziVp5wcu9xYwnO0hDi4
o+Ozcs48ADiXJb/lKWVL81ots7/quq0Xcr7VFM4XnOTalalDlpkrGvnQnyro
vJTeE0c0sXmZQSmL8AG3/6AWkNJJ+l0H8xkcTk/H8NEbrfb62TFADcaYWRir
fjatQ5njQxIjYmOljV2OkkH+/etXx5CwAB3Cq+GZ3WU+xavVDMfz3yruTy49
QnnVPvVdamJeHep1w3e+c6PTlUEcD4s5d/q1kqQSehA4nG+EFP8XrVPzYdrE
YAqMqAO9TXgUcj6RRx1+u0lsh+ODjBUBkfLHNekJyMRfF60VlSMxoZcesZkz
qAITjsUJO70w95rqWHc6ipb68QZk2ZIAq2hBio1ksriVXKku8m9Z5r8fEWJz
ZNIpG4D74v4fbt9iRrkEcPKoPSXdd1WY1AviCzTxcZ3GEIuCD07aUB6/TBLW
PWJXzykYlS8Aa2MYau4xqCyZiELrk+JbPf/rygYlgw0T0d+uAKDcdM0vMnTk
OaPKTkPM8Z6uD6jjWzcH50JS1w54HlkKBmkAvccZ9eoZ+so8ht51YRw97HXQ
xums1SMbcmRDUa/C41z3YgjQnE9Xk3qwvXw2KOzqZKtlhj3EZKEk0fMWx2XF
LKm57anSzmZY+/NSd3jEWoWOTh28ch6v0z3AZyVigPVbcCdA6h6BTO1+CS2V
z/M2mgVe1xLlfIMRmZuWkE9By6UZr1slIzPzihTYCfcQhFS42bKfUQ+VeVy9
9Z/RSERunvblvJj0qlYPlQT3wyuMv8qlqKSGPshhKInyrw59Cn2NrEpioJH0
Fg9ScFPQbGgT6DCKW/X8eujXc0fdHWxfmBS1YBvHsAGtlpzL36mOz/KYwEzl
Af6PuDt0LJsztXQsQfDHXDoW5CoqENQoVeRt97cH5QsaDpeOq3arOYoJjRdJ
VW3Tf5K4IGQIiA3Jco2qSJKkT8QPfQniLBzRGvmHr8rM5xsywDvaeM+PVpfo
DzGXtHdjW3yQ5tS+V/JTh7S8g1I0lbI+VJbEXe6wXRC5Du5vLmpnb6UGN0f7
YtePb164aXDxkouXyWVceYclfoWwLyHTjJn76tgtZdLDGAMpwJrbpzgDjV0X
gj8ywREc2jKdAXdx7IrNJgdVQzSiP/ukQwhKi1CQK2s4kHwWL1dfjbmYA/Rx
NJd0I2m46UAvyjK2oqMYEV6+ay9xnk24eUiN9ZAEAdk85wQp2Nb7uyKrpsnr
7st5FopXjyFZp7dL9zPP8HKQ8O8c0Us1XShfgS05EpfetO2w89ZIRND9yJJq
uoFWD7eNcVvfza94+JsP3k6t3gZCsO6jij6wv8n8LVi0Fjd7C3LpoTggKbqB
Kh8T+UZuQoAdOq9xR7B0Wwk7yZhObwu0TrR6zN3tmSWNWHBPxXAk3XF9ScVV
17TW4Er+FrF321MBb9LNua/OmM3vuFUoT1voahNSiiPfC/GDtBEQROGVkm5d
3MDj2fpA9UnaDnXwv/X6Pg5aiSQ6f2YAT0vxmMlxrrze1UTNQ4VdXLOIZTbP
I5M7g/+P//x3FV11XKRwavDbJTyijtDwWTzuEgjbXD0ubvPEc+lzBV73hy4b
rzTfebWKhlTlEM7qyKDEmdIVrr/CnWKP60LKsHFa8ZvcPwHyZgamWrJejfCG
NT90UnA+Nbx83fk1NjWP7kkDHQYYhKu3PWXTUi1ptBNUPLjHl7uDXkQHb6j6
/N9p3dphcLnxZfu9NU7MTqoI6w0cnTU0SWYBQRplhi86smvTSuQ8AcKZN7Vj
3KEMF8aU5bFPa7UXR7DFsdKzGodnMzNtpnhRoBb/nJgWVlTjT/xynOWjaSzp
wz2WvOrPDVWvhgHJSJbxCeSfJdgAMbm8boGkV+Zm1nbcNoKR8oswiw8LiHe4
1hKttiPQS4RyhJXxMQlt99ZibEXbfx19gosJ7G06sB1loiRLBR4UCFGi9lF3
gtyCkw6V+x12LU7tJzV4fcqkjTwXoIp0Y5dYd9HNtKUgsFsZejM4mzoCMbf7
Fpuuf9flJNOjZWPMd1vZoSldKErXK63IRo0ZhFUTirhub2SFLECD1wSOEiTj
6hXLgzTJ92P0Rd6WjpX7zzthpsI1KzkJqOF7ACTBkbJbLW8Re67BYdqMfLVB
dyx4BfP1iGQl8RCYBh+el0boDc6xJuansDfnEM11iBC8aTRujwcG9bClq8ty
6ZD7gRmpLVq/iuXvm+HYoERXTJljYgpl0gHtowxC+dDrWp4Y4QSJ8Pdxn3UM
sTG02Qhad1q7AGoqLKavxYPNfZ2k9iWRHMBjLYeFCY+qcYtb2Umua4SuMtgU
ABnGYNZfCHl5PrgTB9we5W/ggtJgniDBe66hAwL6kKuzre4UP1JZZ3jVZ/ie
7k3rArMIWhu8znnJL4yqnviJa003qk/FCnRw9Bh6nS8ltF/MgZnkl2sWhMb5
EoDqKpVcuV/mEzq8pVrwfKI7j5cP4ZPMYBBdC+VdjHi/EvNQtt9+cn337WrK
BIzgrW8atQ9Vt104K8qGmV8IoF3INJfMJoTtyau0oyx46exH0ZMfN2D+jZY+
Gc1FyPU4kKNELSM/F8qDrfToDLEfJRoZeMzCkJ6sm9//bfmutJWSOl8PKdWH
j9XbeU/FrLCshoF059rQx+DxWu1GWhvgtJ9yk6w0Xn+iidsZWRB8lsmfZF/K
oEM8pEGP5v79lAO0Gog7a5wFs3Ep4MiSPUu80UlHsA4W2ifygu19/0AdcE9i
ix+soGJt01DNCOdyFVkNwJhlLNiQ7RLvyKL8Psr+wNv5jW2ROfkc6iAhlWG8
r1KNH3QoD7nbTg/g/HXYIySoiQBKzpVe44UeVytn04klqTpZWHFhGgVlwt2p
IuUuuemDm8gSf9meiVaNo7t6pjP2uBoBbyviMTzi6MRzNqj2xog6eJiMoqAa
V3QM0A2XHJP7xW2df5z+J6DY6yQNyGEjMii2k1aBk3TQsaBjNpvFc3r6Jpkm
IJJGEezk6dAJRcOjo3d4Rmq5uzmFtzSBbsRs2EMA2BZheigJWW6ZEByTeujg
dhCrkDXlNiv7gmkFI9rfPDjoJtYame2O0OsNMx0/YS1d+vzF+5FlvgYGgEwU
N9U0Q2gmJik5ssGqkiivCMe0+PTS+uDPeC5mYGPR1A+36gSB1ZoxCJjMQHCC
ZmbCp2anmvj0N2nTuxyi1V55OhWaAadc4qPjU+pMr5lGMgjNhDjh+MTYvoPi
ILtmClQdVQ5P1MfsVqxgjtbKhm55Cq5vFQD7aBatc9eGthfwyqyc2zW45Jo1
oWRvFFkkKn8vq7FqQckUkAYiDTqq41vhooGj1iZyZCAiz4x21yr8t2QvlGcy
qliQMaKwntQ9lhBuyFhG0/fxOYKL/JkrwSQMzxskH6kymzHg6oFbca+iEygd
ylbQ/EGkClNP3TYuhzAz+tgvJDZBBSD9tC5mgxfPYs3EXlNpRJ5akkzt/19Q
FTytSPQHXyHPM2c2yMYK2kKCazTPWYOuqiwo8nBU9TV/grxMFfoxvirdSy08
j4/kDpESpWWU9yYianCLbW9hJ55Xc6aWGTNgc9Fqq5MQGKv3FY8qhoCNB7Uy
f1P1QmqIenjRvXhoFuJvstEQQHDwJPPPopb1ZEJNaKwpignnSLYCHLQkpomV
xgZEXTKzfEQ57fcZ+OHweW8iqbbRa9QHzT3I1yFzFYxbbBq9yFeyuths5Ow8
8ssq9lgNpeyatGPbSf8Zt5hrS5HiVkWFPAbPffvIo0zwBqdx+H4F+5pNVdFN
ViDqfpkFE5Dfb5IkmD0aEDtiT8tFha9kZugNkqLOpPBpmxs7j/+50z/Yd3+O
YpZIdhKtPzzdcXdls443QOBgFJrlBMMmY6MaqVmDN3ZYeDNcsX3c4MWLcHzS
1iEjbKqo0A0swLacY/BH6wcRUEwrUonDqX+/eEK6MJM96NnOSgwUBgdekSND
EOTo6sdE3EhkOFCLNBU3EIIrQL5JTGlEr44qRjZMV67re5NW7ZA8+uXow/r3
v4pfWg/P+8wJ3qTSfqY+VgfazQhh5gUr+eyNgnh3rGshw+4/n6NWSedKBW3a
1Kw0vUUHN/R1wyqfYhMB9apKtIKO3VqwN0p3QbGvx9asyMw22bp+b9I0rFgq
pnsZHvcn+aP1G98AcjFCDqefN8EjcHqLV34FmPogmZi+U15ZcYCkReqCR8Vp
HjfPveUvwlBMDdIdmwEAkh3QBArPqDlNODOYB8FXyG+Nrlgc1iNhy0Unz2Cu
GRpbzIA467+lTrPyS95CoHYyBM2CkQ14iI/lUq3lIn24qWveyEld84+aBUWV
/kppQNCOGuN3hTtnaNC2hUK+e3WYUPoYzo+D2HRnxCLSVq8gsl3tWG85Xbir
a7ka7Mi03kWwbJ8aE4PuCd37uLAZ+RiZLpD7TjV417gT3DKRlrZo3rThFZIa
HLpGb5XvuRYxJPC1t0mdb0rSrjR+am4LZCV2yZ6REUPQ6NPRj6LPl/xf9TLu
dTBiXbftTA5Pd3fSf3hG9fT8Pd81lXIcCK9cRZ6C/aLZiVi2u6/o+lJcbwQT
FRLCy6lYiaRjme6rRE2jJLxe3mJfbE1hdHgWHvfV9/7oNhJuq2LD8KuRmyLr
tFNys3ot+inj2HKFSSrt3mh5RLu8vGBl5Mk3yRuGkyaenJr0YEL1D87XToE4
+nxbnWLLUG/HK4QkWpdbFOfwTdG74KL21CnS54S1EoBPvGMkZT1t4kulpUGs
bZUxCxALo2lnJjgl96AfCtFE9GaJ2V+9njuanX3p2cNb0HvqBo3cNMHt9DFH
BpFc7mg5LVmeDTRSx1YZKzHLE66z1Q7+5XybYKtfVR8HEjgoP8nYjsNzz44w
NLuGlp+1Pkra9DxPUknwQOm/YnONFl/WvWRZHbK7mHYOHqMXizpn8Pk3keRR
AawEDRYu3hMdij/57HoWRBvk2z3lYGPJS34GbfSCQqdBvh2WHpDUdWWX/fPy
IwEmusyErv6ul6/f//v0OvYg03oLKMGndLeFw/j5VMmv+T8jr09o9MXhPhXA
/UkT8mqt/RcVso77W12rXcBKf9940TolKT9XLn7lLKCBSjFE1UQv9+QXkmnO
1Mp+mbG3UwFsxv560Y7VheHNGcqplhPB9FSWUIp41/n6fNsku+tbEuLHzQ0I
KVGi8WefctIZTI4i7OCItTHDUUHNAnqhvEKG6eYYD/XbEysF6JvthLm3hhy+
4CO9HmEKm+btzMQwb34Us1BkNk1P+NHpGOkfyueCOeRp+Q1h93VnFNcMDkXE
7ODVKKT3S9knF+Mth4e+lcms7fgVQ8nlwRAFN0vHBi90RyYuKfD0m4HOvnjf
ILEOC2qajrAjLq0RNaKG8ngLJNiRv9F7pVHHh5/tn/CzMBYfm+V9PUExNxNI
INKpzkYUwC0M3M4isuC6DviU9l2Zj+YesXd6D2ZtI8SiITsTXRA1LCfa2JAg
4LrqzyFwpT7JrrFQCm9eZFvr6dcY/osuCu8dt+rDW/uQC/ukaEAJRK9hxISl
vUzm8Rn5z7i0zA5v5AZKsFvBnH1Ut16Oii/BUUmG5LNHgxXkYZd8YX0cGrRG
YabzSElsRDs3UrJf98WaINx8cdCOMVIAnMqqD4PXUv1OBfZcHK2nRDi4VF8R
uBAAY5W7Tu5LvB6+2J4XAhb4g/ccBtkgvIcOzVCGNW7zAbIqzqKYeQXPXdKG
5yunnFt7pi4qUB/grGu+rPZZfSxkFynF1iPDyqMOmn1zBuvtpaTSduMKMSFA
xBtE3NHraIn/3FcerdQ+i7tpPmFbeGldb0Do7cxGGjw7m1L4+1u/yDM5t645
ehZflBvOnZdqZjRz4bWuItr8uQKgVAXZYOOxFwsDZgLBuctFMsDJkgi3xaq7
XugfRecCgahylkx2lEhRAQxW2ExyoWSMqStIjE3iYpuEtUQNaUsowHVNxeAY
CuAH3Rm0YoCc7ap3RFdrOzkocEd0uoRV6rqP8oSzB6sqMRLs28iFdN+ma7eU
VVvFefArR6uhMJF0SyME3l2xU8xC0LztgQqNqQl65u4QaqDpSeiTX9bsoruG
ntj/RGNZop4/2ji4QOW8vbA+ygUvpkpKx2uOXMSX/L2UjEz2pOc6uEqisBBF
GPIe2NZC4CneKEULzS4StBUgR/1UB1NLsSfUU3POcE6CStVYtZkmZHVzHRIk
Jp2u9uDw2DT9CzcYkLf+Rcsd8AzWX3eyfym4XE8Fv8856nbEuikE+Wn3bZV6
mRFVkNc23VDwXtXDsGlvIx6AtSCY1LBJmUOW2UjblE2XoXrPj5t+BroVFc/g
s8Sl1xcoZHTRep6guRHwbA2LCCQ8QL5eewxtPz7j/EPE1UHK2QXyDD9F4el0
Vz1XxvWqNu4VTByl31vQqqP1qmATmAzBcx52R7imzC3nI56gecrJlizo4vT8
PfBrtVUyXYSzRv9GUo6cNUi+3DQU2f0Zeu+X7xVzAhP2oKP7PQO5AZ/DI3kH
vIOpcNlXU16ngE6oR6zkXG+rnh4QM7kG37WWANGhy7srBblYOvMLOcfCif/x
zOx7ddybSpcBGEQjycutsHJrS+aQE3y4Qz15eeJzYZxM6bWINbxU1MS814MK
ptD6v2TKKuLypLjss4FXCKx+671aIqzEB/vWgJscTrUKcyhjoA1oaPzSHeCy
/4DCOXeu+90ZPSfSVtMK/UFTzStwIkpflZ7Zg5gUqo+jrrGFaNsJ5KSkERU4
BvddAwNGYNdBHbBucm2iYC0OkjsN5U5RpFdWJ72K7Ew4WnHPNnkVePgzkz7I
WRD0uEhdet2d8YUDKAUt7PklNixTbEpTt5gQCCg8pw9Pjnj3fSO6Bv7zfmOC
4PmlXCKMMMYqlQMRzoxB9lpXr/GIXHdnaR0h5FgeFrqcH48ax8lF3tRrApO9
tWnEvyiyijCUg6XBUGdNacXCrIyIHnh38c8fK2bWJB2kVRizdUIzes2JWBgd
/u8670LlSHkArSmdbyRgA7wz3uTpPsyRx9t3HpxlJ+SNoz0TnUcNl4Fr7Oef
Hyv1I3LHkQDsTPq3j1R3nVRf9UCaKe4F66sggGAxlpi/4kWcdjsaIdFKWeAq
pPpr83J3LxsqMF5KS3kjFwyXxNOMYR6sM49K/E6MlUw1Hb0z/omq+iWIfvaC
wNBg4BgygXRrqLWvIhMZLNl2DnlArn5gYiLFpjLOLdBTTGpEgQcr2u3EhZYB
BQUjGdEkTkaVX2/3soU7Gw71gtEB7sZ++XM4KsryQN5MYbARhvm9wYLMK/oS
IfAhL10I+YzgBYhdkAEblzQS2vkRlJfTcDOpW2gkQIOd8BA4Bfj9e0FBRA63
IDLE65mVuc31KPqa51dtCwVMvaq3s+h91VGvlQAp4pntCH9CyVCPsbN/hKfV
TZY5Ek58VeAn7VVDwqHW0pVbSdvHL7kJJCPAG9s8W5ERNZUvuogqNwyIPyuP
mMUgvNNuqpSUuc35Ll6KjtGmSnel8K7JfWd0ud/RNV4Zp0gRVDiVdfZTPRZa
qzj659XTECiuVl2B8VdiFkgIDc9ogoTGZeq2xUSkvAmVLbaNZ3PZzyxV1Gx9
adHhvHGdV30rhNXG7t+6fUjMvkYCez4kpD8fPEWSbS4esXakzf7CCMc0H9GC
XM94mldPg804CU0XiP87G6/2HwUpt1mrEIPjGcPAX6IQrvHlD8yIpx1IMmR9
ag1Ds+zdWlMWPGAveHwxXIHiBN+r8PnjrOPYjgRRELxrK1Ix58Io4c0HA4Qu
AlKUssvfsyO94EQtRHzykQenxLU8gN8FjcE5j26cam8Pih8WwNyMsYrfElY4
/9/hZNbQbD7B/2df6ATux/Va/8IfnF3jSVgGboeEuQuMx2grjaguj86Pw5Qs
RDkiLrvdei4IFeZ7udB9dJ0aFelwqJcQlVqzgzQ2SP2jl+DcL81VYYKfjswV
JK+AqnNFxz04h2HmuZuyBCK9h/ETKVEIWjpoH/vvAw6m0sO/eAGzpMObwxeV
/mkfSEcsDF/Cro82ddqaoIOb3GMDxaG6QKEWEEFNGA+IKVvhnk/A2bWb+rUT
kWGYQv0ZFiV8raRlvjBFBY2RJcye/DHme09/6SaWsS3Is0fyGjrCbuWYcOVH
bMi/H5GtJypKjF9OC14uZyLvWC8uua7dkVHzbjEnsvkLV22hBxhUR8W/5nd8
QfCE0blvvjO58zXAoxoP6oZhR7yp4iceBVeDABH74xSk/a4TTvtWA/ZJHgk4
1Wg54N7TSlymsZrA2bAVVMu6peboHQ25XNCvxZ4JVWfvE5Qd2A9I2G++A/Ry
lWDKrdEb/lfjSBv5d7Cij2ASXvy7Ji8ryEjGm+SA2tdghUurQx5pfnIFBEjr
MsAFl5PqlZH7+JVcDGv4JbUOi4OJD4HDBfzux7yu06SFkr5go9pg70RYoXg7
xsEhmeKR1yu2/fuY7E9UJXE5nsxX1mdy2QkpOY/x7WXrFOwhPnr3DjgW3YOq
mELoTbBLeTOlh4cTouUEyqaOT1AHIaQj0tM4iJqR5HdnMny2LhVJJfLyKmxV
vPFnkV7r+vdMLhr9upHTyZ0kCzMLN7nPQZKIEdcvS/OYvZK3bFwFOuJa90b/
Z2PnyjMyVblaz9gx+3VRn5UFcZLZZ0RH/BZ5oYEnye0OLZ6y0Tde97Gt2GIY
anVQgm5vCNpe4Y2FOZqUly3LQW5irBQ9uAQSmh2P9ZVjivCX2fJNgl65dw1c
gVlQEG+Q4LQNg/ctHeAtK3Uvtg2QBv7SnP5j2kUlEvFyw+3bN7sn7I6FffPV
Ovj8wyUr6RrnHcViqczmb/8ghu2DQHsRwA8afkqBBPzSkLKfHpI4MWWz7zIr
bXRCvyfEu4reoW25x1k/hdpfzM6YxPExbnRCNFg4mYrY9/JJrY6jVErZjDWG
t3/w1gR8K3YAZolcnah77XLrErd4H5TraxUUzZY2CjTGGb8H8vtT7kRPO6gT
xUJAQW+dgT26a6swtEEbMKFz/wsgMznq3q/ehU2gYMN24q+ItcKL549h4Rwn
MEANepLABFb84w4ToJnXZXz2QbXffabn3Er6MKWfumID5eIR+QjzsDP/9x7t
+wp8CbMjcr9t1Tc1UU7eBOpaZLJsQA4zo/u90m1z8aiABetqve+J8pMxYygB
uM1fmrK6f4nO+oP910eZK16V7g2AJq4feEmWWbBrV4ErzZrRdnjv9bBo6inU
qCFDM46+6NFKK25wMMbkL3PoxgqmsdUBVGquR0vKsjvVU+648M2yYhYQ32tC
FlBeFyaRfMHq2PAOPqF8IclFbm1FDcXfUJLBv8jOsS7UxZgZcwM08S/gLg1n
v6VZ/ipUUufz83m37p5AxtUPEPBf8VnuS2DLb2adQazOv/52ff9fnNm1+yHi
FrZ8miXwQFhXbckQHvv5vXb9Z6SeXPheGJ7h1735v0IVG9lakTo53bUQcxey
HTdqV0QlSxlx/rCACmBmkK6v0lLrZipijFQ0F+/5Zs4YvN6TIDpxhOPo1INL
EWrD9IRjIyFmEovCtiQyRgCBTZHBDW6KVTCoDmSr/B6c4b5sC6DLyuNjF1K3
iEY9ImBqobOFEpEZck7/wPdiTYFABhOLoVYohtXQXMHceLl8sq1N9gg/LigS
OIxFduH9Mseed6/qEHq6olY/KmwTbzmKHUQgA2aJoapNxbRaU4zAGEAOXTtK
YsUXoIK9kbVpLtZxiXogu1GqZvlC9watW9Z0Ma5ihtdGzCeVuMxNa7k5DOO0
1jyTHXgWjss6hE1JgorWEK8SyVXMwqid1sZS9LoF74nMn+y9EOrqzOfsivSi
ZJ+IYTQtx342s4DUKT5hRNXfjdAJ6WuJ5gHcniBNsvSlh9VSquyFbON4aZBD
7reBsnjdL8L5P3Ks6+jTv7zjU3aeNTF9cJhfQPkrWl9MJ85xKTWzH+Pd200G
NlrrlTCf5EU4CYCD27K84U8LirMLOBbjzM53ApmSzRRX98Hw6g7tWtki9lBV
1eyAz7lW/y4Ou8YodPJkE3mzm+m0HXU3bhfjlm64EP2DsghPxW3dKNtTf96t
b5wfrTvH50xzSqfcVXVNCo20vtd9odmdtsaV9RGdCr+eT1kqiBOYOUIOOYxr
qDDnj4sXaw/RzPwg9YnyAnkvlLc3mmTiiXcm5/qaVczPtFUyYf7BehidkZFW
K9gVr+ZgdyXE2raiTpmYWLHhqKr76iaau/tpfZw0byWDQdAmPqvZMxXLB9T9
0H7krkKyesp95HclcvhINzRkqs1odNzDjax56GudIMA+YRkAb0Zm26v4xUVU
b1w4pK/AugpsXV3kDwHOVa5XnVA1DJEzq914rr/1usUJtDeDCi7G3KtZO0+e
bEZeMCfNTStH62TW8LVOiMfSkUiLYit8TmnRwlRUvuavk0cjv3JQuBdb457K
cKSagI3nvPrcGrOoHMYu4GW8EyEQWC8o0P/nRf3BAjT3UTyBGFpK/2dxYS2/
EgO+ILZCu8wa3lLYtQfzurruCTKCcXHpS3d6GbG557HsZQNoDi/bliNd9b5y
dDbIQ3gEv/V4bB+RqZiaEzZLV/f8RiQ8XLlaYzq0fAjMuiNqh9nA+azx1bR/
yE7MI61O9y2uEqMMwFl5hrIpSjVEPtNf9TnX5woWqY3cIt2Twp5L08PNmHM1
uTkJs2bKSo1UbrMsyp9zU5j6aZRdYTdN51V1Meu/px4ZkD3Uj4C/UttaU5ym
497cTXK7vA2fTCNvEVPqO3cYpe0O3xV2IRGBih/B0JXH9KbbYlFyUnJVTMzM
7cps8SZB6GmaUGnScKpjbcXWqt3M5hWAXt8vV/ylxdcSqasY3CVZbgEkv9af
jXbKXhjky9X/AZeUBWeZokgTzAj7VaCs8m52Bx5d6sN/R4FgjJTBNPczOgYO
WsllkgLwovkS6qGXMd81s1OvNSI/TsOMKKLpCambcqWwJFHX3vz8KCmMAQ9W
mS17krdTABkE5X776IoKzztFAOyOUPnCoWDBD9ABHStOvcdGaVzLPcobZ6B9
DW6Hl5I41u2CjlmI3+dDBzt9xSY242g97yL6tundXEGlJqBYHK61UOrk/Vg7
c8J+tAZ8E3yr8wXu/g2SbxHT3Jo5uvmidPZDdcmHsDKBgr6+JMIDUkRVHM3w
JKEVoADmwjLQWKYU8IrqprAQV8WiyERMOt6aJajJApmNsxyGcvQb5SJJAvYD
rrDBedWqtWdCByxsUB5+cf8jPcPk+0TDm2keYVG0Vn1EuEdtmt7vqzYyRY42
UeII+mSnks/TJfBXHQgmBxEkuQV++lyUONFBeJm+iRbLOi4fHWVU3GSpicwo
uMhCAHos2HbB+89daAVGsE3j9VAoiXbNmTTLJ3ZUsCRtWbtlz6KiFhGUhGBr
E/R4WexwAayIaG2dEt496eDlOhpge4rym7ZjowlXwHT9WXKwPL4QLevH/BJd
AVtNFnKgbNMdi2FgP/U2bUZlw/qpFpKeenNHC6BFvKX9DmFmnbEv4Qsi7WpN
BDp8oJYFnH9/bpOxlLd/505AcZDRPugHSCUVmzDl7U8yfchxsPVTEsesMCDI
3jTMcsvz3BgVINe/Vx5TlCWX6KtgoPbsTJwFAAU6jQ316FzKiKXDJ67tCTZ+
KuK2ZY2Lw2BWCtpa8HHR5dBXrgc6km1C4aXCYlRxf/0IxjKbbDjdj286wHaO
y6EX6rwhFcug15bC3oIthu+/x+5jSnVvpCurwf48a64Ae5kYzUThplSJcjtj
rS6sLatcpjse06acxVWIfPElknokRpJcwP+FVklXDZNDMkeiOSGFwzt0DG+9
b4EY8bh5qDHWmZ30v3OQ75JhcONucc0Wgv/V3zKiQvEexW4gQik6PRnsxgvU
WfPVTqhgaIud73Ffxy5J5zTaX1jHmAfC6m8TAU+ZMI/cNvKD9giutLcXkybK
XoiTJuDl2HDvDBOBaiC97xZ4Z/SOSQ94wBx/6iO/10MhrxPTAPcnTlNYb4gM
fKbgFD1wHWmaXkCtNoEOKvuo6yIY6++zmEkIewjOtuTOqIs1Os3OGRMHKJXc
R9ItJIoOgKplauPRMmKyYajJbFl3OEjSU2JetKaI5ruC2nKH+HJktZQ8KI37
WjitiGDd2HrBV3RddE3PSHgpfIYCNPxlrRZ0LR16hCm+u8NDiZtVQ+/2qLmY
Y43eFcqz+M9F8BImkZ/LztDyLroCn/gIJL/vwsksjtGhd3E/RbmbX8I7UBdo
pJ436vYlstz3eq2esNHqEZmfXXBtKg8fZ/l0LOhZSaPd23TTo5WWY/EY2S54
hEgAm6+qgOhRpycwubCCUflB2KigE/WQp1Mxdrg4mdb02KIXcvZMKfmRGBvK
FaJJhNBnpZrxSCxGu6yzIzeu1vOS2Cho5v4ZuKFfDpTiyoUHCamRMkEh3fhP
atPOkY64KANDzT4Z0N9KZqibrHnte5P0yewq2seWMcnBqTd23U4QXAe8z9we
q4gP5sJ9l1mTi+q5iyHz2PSBcWZb+542PuZoOkwWiUbMC88+o4Z+k5ttsb5a
K++dcY5VRlNqzBsnuKqAZd8iHQygkQq/pqXmMzLncKakFKh6YKD0mgiaM5Ji
yasWfuPmcR0uvkC01d1X1oSKpC0ChVLfi2J+21Rubub0O8CfeBskJxh3bK5m
XKzbc3aI5FbunAdmpvvhGPO71InOsyShCTAVdl+rWdNZrwZnBqsU4hf4yfWg
esC1Cv+HtPdDzYqurZEw+EMIgzjBqlSq6pZCr2rvFB2LRDx8NVnRHW5ZGcPo
Q/cNZkMQPL6F2+OLkJfddnqXXVNFOnwfs6x7mdhaeCJSKE0Hc9knHaqxieYI
sHz8gGfLCt7PzmusUIz+jfshjeJGEAaAqf71xy1SNNCHIMjOeQTYjqUinidz
IHTiGGFLdbHdPmQHJ29JXcKfzELNXyhLdDa0NqhIXIXUJzi/2PNXKbzX1N3s
YA5nQISpMpe0nMcvzEnADSIcdimmvxPNIfFGHcBf8s6yAuVraSWp5sSy6Z8x
uJXGVA4jqZu3eo4WayBpdtdEnMATQJbQj6HKoAr67Poxo3no54rX7UBXk1H6
z8mGTpnHKT9CWJt8U5a8tRCmqn6Spu0BrjMV/M+6RrPcE5y+zjkuxy+yLfB/
MEj+2SWBN6mTo4lWCzQv/moN4MW2j+9r1M3gYDPYdSrGyfDPDW30hbQMri9k
+r0UkKnmccw/4CRE8kvma9x8Y31gW3i0XYXKmSKQ5oT3omMEOt00rypjnShQ
e6FxyzxZA3YW+WDJRrEuH9aAQ61hHMbtprPAtc4PL+f2FAv2x3DdzlWd3MVi
tKYP2ryWPRuEWSE/c+nJXmAtK2se3tpE075tm7PQSo4ah/QpH1+kfrIUkb38
7NBAk8UysmQpBnaATMRSLT8dJunyDR/Zhd1rToyocNsy2bUcRljYmPmqXztk
lCGDgaqGdQXvfTdj921WEP3PZ3tzlmMgY/0fHheSvsnNYyJrnlCWmfmoDQlz
ePWNjBZYwCgUIvioPONuRxFrBX0kBFHEU+DdxFpiFx9kuvljEXIHyNIJlOhB
MqaDShUzgrDBmt9wiTLYXfIZ2UFVqKR6jfntD3bze6FFyEjqKW2IaibadxOQ
6YXvEUY5t+1AOUw9WMH5ZaV/wC1TazjHY8FhFLdmJraQthrcbZ0mIjVg619R
c3ECKTsVZkqDkNegOjUnGJQAjs+KAuZtQg/fUEZduTuxOUii9IBeuZIEnmf0
WFv6YjMsB45+6W5wIvluxGKrSJTsKUvOwhs1xsepiT+/7CTMqrc2DelcmZzW
PLwmvRKnFKxUoKwUaIvr6DDrdXSTDqe4VYhu9Tv1FXX8yqD19fmyKyhSQtsF
DEOoJJDl1sucptvTxqTd866OmQDVBTISWUzGeyktBznISzZsBiEu/bgiJdz2
s/6nINOZy2mWPZxpjIBsC6jlwXsFK4yBk8lnzZaIFxewC1PspsymHNbK+8Mj
hyn3nYC7/M3leZfbkfqb/L435+LHoKrL4x390Q6sttBhDkKpRJxz8CsLESXm
tdGrfyglAeNlKggBfqemzwgUtlF/lYB7vxENXKfPdv1x48Vxp0o268sleIrN
PZGpWj/hws1W/KV31HZ3IOwxL6FYbQBsYehfsXcWNCLQgfSTTDGGcZfkhU3H
r36eSgu9HxAXkD3vJ79zswPCE8TRBWQBQOMkcqVrPL8FTKSrz3InJFuR5DI4
sZ717/XlXjAI73BY7abFD/92/Twjso600anUruknb+Kn2JJvvDaETtoakUKY
nHqvhX5mis+4w6nPqrCCG2YNWPI/U2NxZD8nVbaIUUlXJBREjmadvGTLw2s6
kfa/H4YPkZFL+/QGaaBwkqmoa3aPBkRYFFGd7qWYbI0pzf7nkjZhCZn3GxkZ
aRivm+kz0YjMtffeOakXIYV5LfhcrwiD+nkjQRXXN4DOwNZPJs1lw3TQQiGr
/gkV6MuOtyNerAWF7rZgcOWwi66jVk4TSP8GiOPSmKjdz7Rnw+p20YcvAkhG
Xe5Wj8H/lgqqnCiPGTAuvEPmIEf2R40WbM5P9OLuVwpHTl/ClqnjsWoXUXSg
PKBhvkVMmN4KHqW4w8EdPe0gHo9NUkJcLKtVmgUs/f4AbixYfmkWGwomiW7s
KPCmNA2WnEwX9g8n1J78UcjMRLA45H7jW3WPjsuGg7DrFprrgAhhFAbusvrK
bz5cx6XSX3tIr1p3mpSYsNl1zcVIpC40FttoNB5g0KcW4T0VIxC9CdDHaUew
lh8MiYkjUCYF5Fva5pxSdYpqFLiW/eIpWsNNQYd0cgwBreyBNaKJ6GgUc1LY
LoVNYAp5KIuj+e6u1ISzMEBEPtlEd4VSKG4rPf88ycqHpkyFkN+cSoDfYjXu
s+ULjImkxoGjHgVL16pKFWdH86TDhfO/WGVZ+opBNuSq2A9OOur6HPWvGvOM
Jx25DRacxRr2YStDX1n7IxWzZm7NoecFlIxNgfrgeRrdRZxsjkCBcmW8nYiE
MU1+MfBOo6hwNOGWDWtdHRDH5t0gzEoTDGrY+RCMdiORI9gcmOPOuhXK4PGd
GjDiplL82eaMdS5cCrj15AQNqS0DLjnA3yD3spmvE9pKgqvg+PciiBDcDu5Q
nW4ksY96SuPSO7ul96GoA9lKQwjhaEAC7BbHcuL6+Mq9F17QIbU2dTCOc3qG
YGMwyGevmWA4uUf/JYKSCEqCtiZHUscpQ5krObEG0npb7tqpkZ7C1jAIMSrI
CDdkGkZLWfwCpuRYXtaKKOWS2RNIvBP/7umBhIaY4lSWknFgB3ALjGlcP4AV
1jBUopi5t16Rp5FAbvm6jId2lsBD0F60T+q9MCO2WomqW47LVAhfawlJnp+8
6PWufcKD0W/sdRqX1Wx/tVzmJ/R6oz9FrH1avFJvKlXrOE8B/xj3JHkS4G8F
MGisRuu/JwXrDhuIHZDhzfJJzkRI8YaeQ+ghqswP77heaQhcmJWQAJ5KM9zF
LHHhUQ21MTnd/GXzqE2Dmgrpj5dFBrQhMXPqaRodE6wVlOKvQ1bswEh8scUD
49bl/j1kElojH1uNmV+q5PrztJZqEqfEvHcbIP0ljaadwQhRbUGK7UBo4cjL
k6MdDDKwyNXg5g/tb6wm40BOIa4omiYXU1s+Oi9fnLsNlG+uxoc2zy4C9J3V
AG0nEXkhgJEIJ9dOdF08gfzSrf6AyIfc7VnUHay0NToxTJ0jaiboeYiGUWuN
g7ugpg0WKPdzvXx2yWOXQTB/IxqA6S9yJK7or4zca3Xnn4Be5p912k8FcrgY
q1Jfu3+CylOWPFHUeHWA2RFpsxe4BnVduXYFuMDj6Pk3WpAODEV+p7dU45Xk
kkVhas5h8uV4xTd9COP3V3lNqX5U56Qm9FsWc7fyGdzBhVLQ/lthd2Merlpx
z8RDvuTmqb56bYaREtd9DVCb8IZMvcs5+xQ07daQ4hMTmPvhqH3XCOliDUuD
JHa6tJmv7qpxFl35SpBvIemEwDJfa8ly/VljpI1/bAmv0Bm40wfcTIDrgLI7
3KQ9JqZb4aA6MBp36tWvYPz4ixBnj82g7L8FbJMndanCddsl7Gu33cNDk8qx
03Jh2Piszj2dIBuNdqSD00z2DVTLrWE9XygdLc48cROtes6jYn6H1iXYNGD9
VhwhLhrvML6u8vvO1tKzx0r5K5zdDoVLaGcPSfNI02HmoDNvXQCAn6e7b4cW
mZ4mcVaRA6vUUL4PbUM40nYqNvoAPqH+mSG6270zoaGFbGt71/RsGkJor3In
UYFrA5BonhN135IaYdxuNGzt2mZsFxK2kWjG2ZLsGG47s7M6BWY2GajLSSjq
e5YCuxSVMcYyst9I7a37cKB+Zqa/kVMtokLb9Sg/ju/4rLtVidumkSp68Ee9
m7ALKcyX7ll+W46UY+njHBDejjRedvOP7Tv3Az/Q3BlNY161Jacrlhwke8WA
iNPYZX88Ksh0XnZRPSDalodUcHBU4XcdASJmK94pchnZcGIuA/BSv+iUynfP
zyVFMBpXt4pU7OPmcMOdsYU5x0zPvwsgn6wcLsbHuwqzUfEIgz0dMLc0HzSD
/NY+aUL1AGahS85xYHlF9cWxB2ShfIQD4Tz6PcsNyVF84kjEnXcg9lf3Bkzh
HulNdSuLEhoYPv1J9+PlAKf4Yk2znp+Yz6ItKfmtnmPjfPPdQcVHCXdPJMTj
64odkelPzQOHc/7cyrhp/DzpGct9rsyRVMOBGRtKPp9CQBYt07avMCRCBOXr
kEaaDKOPQLYN+hIbUzB7j6ntaNVjogpNXXvyeCneZfAxiCHHJKIAyIdqOcT3
yK7FvP0fJbSuxGkfqm2LqUg/t8BfGQSMZMrIzq8OU1ZY+Z4dd1RxCzqZzflC
YzPQXCdWxQrFOGUqznXDXLGXCEIBAG4rP8gn5BhN7Ykso4n0suE4FWjWoysk
iwtrJGWAZgj9VVTZ7DtaSVzdGpmGKprFaayJ5eoveAr4p7sy4ZbXq+KtBwCf
zz2/NzL+oyX18bCXzgS3dKz81KoC91KL6OxOEjWLnKGCdvFvWm+9dOd+0M2Q
IU3hEzqV9e8WRUvxIYivTf1XRvIANV+VI0wcxdQetrExL7AEwd6+FI+LxE0G
M5Kit3jy/9HgYCbsEUq8T6oD9ZrUvfo7PAyH4XmG5jpdY03mT5u+vveGEalO
2XBfern2J4Eo4Ir5uHS6VAwplOkv7OAS37Qs3bLzfcw9Nh8qFqkXINcTkWIT
mlHeIfiKF9OWQ265LdezoK2l2TqaM6kBfZsOxYIME+PLSWVO9ru1iG/kOhZS
DDnwsAYsiJIX0EtNCLhxtE4luUkDzzHMNCXb4sPZ30IvYvX1mBJf5lGY+HW6
XTqJChBOsfb7nnZTjbhCa+vqutANG3M7q94DAlYz62tcA/0AoJfNoJnsFcHj
d34Zn7r8Y/8oKa2Aj6GN8Ob4+KEMcrvCKcHf4ENy8+m/WRXBNZ6H40ZYhnCl
Xj50c+FEPArLyRRk5l09V0bxjXTHQC6txJpkkQGF/HDD2eGqOts0Np3fwMIL
sErZqYxqZBu8W186hWDLJExfV4B34kVZc8MjvCdIetAu+G7b3tNvi3tCI020
U1iU5uIWtasgcywRRk5rDkdG4l9gt7Uk16h2gDglYBaTE/ZX3nlCm+UvfHpa
x6JxDp6Rz2RecD7xEs8Wq1icJMMY1EYp6vFMqtrGyEUk0nnQTWUXzrDShtkM
0lH+OQPYiCE81YFH1xG3nUe8cLymnJOCzeZJHGFKvAN52D6d1zsnfr0rWTYD
2VbRZjAS0444/wF2I3RnhlCqE7K/jKkhk6BcBt9K/sT6TNcYDxuWxXdhmPYs
LVormeVVu80fPEc6j/Nl2Ry+a5oxRqLrcMdciwdqg2kNNpIlJ7mgHEDElQgv
V2yjwoePwzsZ3Q6MdYh4gLcaxkIvftGX2mSV1JvgJCgzh8IJBAxf0/YgTJ0M
hNiZDziXOeGzw/JMYOh5r039uUm3BWASmCDDqpe4DZpLMyK419dH8mMACcKu
xYCfKTwHFMZ2+eosEnY/9ebDsp2Cqc8sIaDsqAWK9wAquYcTdIVSqjAMSa/H
3bAkQWcDqw+rbkBePKaUyBi14XFkUBcAAdJC8x+PJB2eCFlllY4Btgi5pUBl
OHZaVNZJLhvLi3eQXueuVZ7Mpy3ZWM7e/x3ah5MW0d7kccNptxVJ830dxspU
fYeO+eLiZXhnuicTni+0mbwVTprle292uq7StvgU8Vx2QiXE4snLvFbuhqkn
xcZO5hCYn4HWQSTC913lDlnCNBm+vIF3tAVvyQOoTzxrkC2itJHGaB/a1P7b
UzHG9nfYUwJf1cWzSK+evUBt4Fw4ixFnr+3xTMQi8YpT4ZWArjBhadz38GhI
reeT4FPZ1R/OQaXsjXGtIHwa87xnb9HL0pBTHzJ29BjIUMYaGMAu+9ODir7H
jvEi2EUvJIjA3DAH6OsXY7MsimRNBUaKCvADXbNNSJs5N5zHkmfoL++9UlkU
tQtG1t4XsxtPfv052M2S6+c8a5HmyTuewlHh4fwBqWVSg0jDgCBCi+3gzZhy
a98LKe5JDA9hzBVVOHYb9ncCSPJcqtFRCoQXuDrHmAsa2ghGx++ugliOaEko
YNHfehSTbvA3/tNkC4XzHMevcGYrKgjsIo3JkdfLLoVGhB0LV2W6zFSD/Y5C
Xr3DcRy4r17YNQfs3i6cMEkhFyxsYVhVNv4LRj9Yvn97n9gfxCExMdZ0AyiI
INTgOuDu+FtPLrzmRTAqF7v+kM0UBTZTX+OVLuksYcxefS1GhuPgkmrKM/DT
YG63oW732vYpxoSKKaYO9Ne8+RYh2qzt/cSELzRHqp+973TisBuh1fY+Xpax
RfBjBpw31WSB2IZSMMi2zgeWRaoM1gscju0qOfYkUeOJUbWptwkT8abwNvHv
yVd5TfEQHeJMl0wNF1z7P/gDEFWYog3bCbJKRtpyw/98Bfqyie2orBhqoQpW
ZZPkN2y90CvZcMu+sHGATxZ4e6OJ4mVJulYdQEbk86h4nNjgDorqvsdWE+2A
R5rrpSJ/b10mgRVPnuNwOqKIb+3pyG/4ilFlOLZUMoR0c84IxLI6bxeBuzFg
kDr6mPJ83lf1OQWoNrwGrxMHwKx1gYNOC97EUp/47ERVg32W8yz8AQeNrmJ5
bDmfsqil8uBlLWzcZssmR9mZGjfJctQF+LrqcwiaH+hn5Uv4XOXdGSuzRSGq
MZnYIS2rB/zK69fFtfEkdKn99FHV4UKSQQhe30kLvk9/GtyS4DhwF+rOtopO
nlfkw92VEYIEROHwFMc/KyP7H6w819uNeKLDj9cITVbM+vSFlT6LWI2uUNtW
wNIgoCN7/XTh0Ej+mTxAGmtIzP0jA7vxw+wb0PuiWAuf9WiasMmrKvbA+vLv
nGff5FXfVYpEWyo4XcUHqxGAM/EgM8SoZcGrkDI6NH/ZEk48TYDzK6+oAdqC
1hxounPIN0hchbGzySr6Xzr582oKt303cWTPlSmNr9Qydn5zcuh541bbsq5C
Hxk068tiUpsFDv/zrXIvNoz/egmC02jvps3lTWfB3Kl92TScBiuMUojqJ+c1
GqTn/92Pku/HF9QeAqFenLLJKioIL6geGX/8FvoOGIkSMGCcrQWF8heRBA/W
ZomCL9gsOEoVt/TupKuVWPJxDd6kMy0zTKYnRCfmVXDxnNyXW8MIeog5aFv5
Mfhc3lrefrqmcsY/GI+dVi3ph+gYz1+ekMbhsFzOrKjeF5jeeQS53ZSyyCDT
ZY5H28ILProomAmA0e4KzGwq83labCIhtntpk1pgaBcUhabQ8cJImfmddAzp
hT468XhFovo8CxYZ8blB5gqFp/YgLAuedsW/ECMWp3YsYcVwMdG3xjsjoGks
5/Mvvvv8H/dOvDnqyqMVGcHlH1KNF0s/dA9lmXtFVtze/VDZJto8LM70MGho
dsoyhjZRbuD3CxeGNJd0KyAF+ufp724T0xp1gBEQ4CYqHwOM5mP9JrolGeHy
BIRvD1YtzDoGGbvTNxMNZ6rcLf4BpJXskZ8GeyVHjGKCoGPW7JO90xsVfQwS
KG0DDwvPlEcfgIiGAiqJAW45CfWcmfPtiHEeyY+gQvLzQV7yIstWim85Am2j
cqJolklp/ZuJNmpVpnlN2lz/y9eBd1FXE0/5napgFQ6FpyMI4rdWNx9XBo69
bFyFQFUcLsIuKMCtm4H9SVNzAEEDokUDbsTP1DL+QFipVkZbM/+StnE1A9UN
QHoGrYaHApBBf44WOGAuaN8r6TJhvNxRfhxLpocaaStnH9aZYmWTVX+Ar5fl
4WIEtwAzwq92XZe3QMkCzOrSOsOeG3kdAeYtTV5fFxTcRMFT3HAUAqPoZGMC
BlYesweoXRMTtzcbmYyX7kRmlnCSjHpdx9SvNTMFkVjJrc+nqui6eA9Awce9
hKYOp2n0cHWCFceR8PyyVBYnOMbn0pM5I2YiXjvOpN0t/adZ2Wv1En+8uRQQ
U+5yw3wWR8/Xi23YF2qeCWymZZoeHEOrx1ZM2vYgpyxU7lPDYyaSeINI/v80
N4VVuxmQ3RQ3taACK4oV8e+vkLjyB8+pOJ8g5CCWqO/PBtWnRWDl6GzPFiKK
cZx9bUm7lJ5yr/vJNJthB5h1OkeKVHl+ETQ19P2cW1grGsMEQ5EF7001YfCZ
dGGFs4UKWsWtQpKTNvzzvpUnhZ7HO7yWKez2y2ChEMWkRSjENLPHWNewDdCf
IhHBACnfE3mwwGoggr/0SKx+UPi3gEqT9/C43qnPfsiUppJX0OzjQP7VrtW7
WFpUq93Z7XQaPP1nzy5vwQOifC2X2xVL68BYjq376fC2u1z3boEYbepD218o
qrP9eeWihHdB7p7+kanCPqoo0USTzcwjwx1SopziMnW3mgJi3fIZBVxkYpsO
urHlS3OVS7x8kF1FrNf4IMmA6PTtUlXf++KIsJq6i8yycNGvxbldP04XpoDr
tbBNWk9e7J0k4wJSB6dPvti9z1lQYfepXZjbFJE+qw6Snv4tFFIflc9aWWoF
YI6Z05srn6Ff+ORDcmz1qrzKsTCwltsdO3IVSuHaKUZdfwBXrIAGWf1b+6nt
wiSt7q2u9Ijj+7TRrY3zzQKmGENlreyEXT76d7nYnyD5gXwbwrk4siP5QTpH
oTwvbWJL3tn9UDTMl/BsHgVef7WY2UCMCvhLJwPZF24KfaIXxsbesXtoqksq
Mqwe8c9aOfUCYQtcPjucie/NQVvlWOuWRTns6wH3kiRZ5Opkf5WhVM94+c4/
FjW71fR26xZBWrm/p5mf7lvHLyGLnL/rEE81Tas2nTe7150VI/ajKnhg4ybG
wYf+lXFqRyIlLlHVvOgPLv/N2g4QqUIHPEodSuWu2sd9P4Bq2R3k1OkpzB/E
siZo+Ia3wddPxX2raNoHZQq87l+/vFVU3Uo2QHRAgianQSlC343v4edhyBwr
hsha099vONPP/LB7a8tIgohbgBhi/M4XyW6KO5PY3GbOubIj3X4cTG9Qor9a
JlygfUCPDBHbugAiFPBuW8t2MXwfglfPk1cvS7TZFUw9cG5Ir1MJNB+txwjT
iqAFJ0YRZQ/que0f9upsBs/d+2oYqx6uaWOxyV62R1v7spx/jYl0NxAPFYDw
nPZjL4ioJewZl4amgMf0mVHy2nn5icGe44hzGAKQ87xWFBudgN+jiOZa1U/D
HVRVP2143fYplZPeZBIUa8IrFqfrRwwLfx0riYlMnHi+gUSUO93hFDp7HvzE
qzCoWuP6CVWdrOsT9oOVOFcTdUF7AyvxnXEtOjFcyOVbgiG82wcKphj+gRCs
r1ZI7fJyfRuRFExM8Em3rx9k1BsRr7BtooGJbWvcTJ/spubk5tAsl8fxl2CQ
mjSgcY4uq5j3jn+qhc/y0HKcX2sE9gA9zc0dMmlMqzsmHOiFv5MZRsEBawh2
ncYDHk0ez1yZsxNP53XA27dONOvTq+wa9IzPd3Hm1nesn4QCgjodraG6dEZJ
3DKJ0Xc9SQu2MeOGx8P9PIZF/QULopWYURtfQi27OH3ezw6KxYueM39ec0fe
AI/rSFYm9nnzy+vvQVIUMJMZWzebT95C8mbJf+gxx/sWfq67DuMcT2YbYhGH
Wa/NE9OupcP/Cf30KZDmQKxE8qQWmqTRvygNmHZL3QeqyNAbeWpzXxJaXZeW
yvstvB15NjejzqQXx1F/aKBbWDgOE/U1hLLedrN28aC4ygZRyp2YBmCtd3rq
G/I8nqxUuLTQR/gHMCj9T1vc6HkX306FD+6Y46YqqQrc+fQPKtmRD9UJ+z1x
z3Tk8jvEOSCOtDuy3eYUGNNFdCFQgDXMTwBqwvJyXHE2ba+EqsTXR2YZD2ng
E175W69MRvNLcInX2v+7WzKxUUjcBEkHR86f0Gb7480fpm29vOU8mOlpOci0
fDU+UbVfcALUqX7Ljaick/vEKlJmYbu88EUD7RsErkl00pcpmp3cgF7Lrdxr
OhO1RSDoVQcV+2u/GM0KtuBBn9AboCLWCQSeWyA8FyuVHsLrqdc9acEZt7Pu
pftn/0F/i3T4WtvDBrknV+H4FZWte5NzFjmTt/jfRJKZTPTtCmBXz+d3MfLt
NJJ5VOEyfNnDecGHp8WNUas6icIbwuuxjpLh0miMJAIvrwCeSt7y79UXe6Yr
4NCDUtwhi5i4ZSxU/zcEzuM6TpIMetmsLmRLsSBMtOP9CZrJmyQ2RPLWsmtf
wsAd57vuzXP48CcJ/q50SwS/xVVdrCQKFcl2uwY5Q1UwJ7n9dIfkczgXgctc
JyDipyUJhgYVVj5CFQyrRK1/ZrpFDwj0KPsXyzTE2Afcm/cX5ZHO28R2I7ct
UZlQdVPFo1o5icxEWqMsTUmNraKE2RCXD4S1dkl2gFoiPe3C6O0/4pOeuCvi
quCCad3CDue5kq5Z/zPJKpW+90ReMOXL5HfNOvu1K90zak3CVnQU5HsPlwOr
CXApqD5SUsZYHMOVJuoi1Qv4kwQT/ESiTGLd5/96dxXuHTKHsXsLmOMKlBGB
ZUk9NBmp2vFOFdIrsRpoZefBOqj5jViz7fumY36G7G8mOAsdumpkC0WAGvAs
Qw6rBURT9cIRkcnFIdM81ZjpOmFVsfx1EOE3WfZvFHAI01TMKPDy7EPRVHQ1
EscSp3vSlT0BMMSrbIyz8c14GjYwU1RwolpLFxY+Z05B2ZN4hKrT1PqQH4WJ
jFP/I9iaK7DZipcZ7MYzKwRVcArwnf3sZqmGwi2OGiMT+VayWMBkAcEo3Dt8
01Y42LsWgl0DBdURFJmyMEj6juKUSw7r55PNd44NIKz6EHjop/6k4LTX7VC5
wzq5sqnps5l6Fhgkpo6zZWyZ2ExzHhRjeUdtyzjqDgP5qHyNBXm3YSsu5tFI
/FxrY8a38fEq/AwXBZNTAcRFtZ9G0jUyE5K85h/E3DnIMTy4yRTJ7N1+mzVS
QuO1hyieGt46WfL1AGZP48xpc2rWQYErpEae0mll3/KLeWAq20iUJ+4rwnOn
oCRnS/DIzCPlUU+D4HAz+XyCCxDozvkqua5xdH+IstPAmTqKcvnPbEFcOOEC
vK9KAYiL5Qwke6abHnDPydswvAwAlodD3daOXlo6/4v5y7eGdJYFR9MGzhHc
487qtMsTa1xWJua2V5i6oK/aQyCA4Ts/6R9Uv3WpyicaN4ei9F9Vrv9F8UxE
xia8NclP7btB0L4c1k7rxVnJpUdcjUH88Ak6gO9arrv2gn178zU0ZlWF0gZS
XNCjus4B1NWKAbM85PzBs3wwH/+rVV8mUXjty4uttPOiBIEPlKHuRPui9ndR
77tx9N7ZfmhboREXgCUZwvE4QWjgoehQ2TIcwXb1lKdKMHD6uFnSrvDpZGZA
DOBwG4jToU3ASYLohTt2c5m1mPYC75L3jnfxH11TNxc4ZDB8mww0AeazvB9E
iAaFOOoDUKcr6Ob4p4PsIJVpic6YG2EEvnQNojbcQtfFtnnOJi/rcbxnXVbA
oYKOu0j+UZGJnaOVCmnTcrnyPHy+40OcrlwYNxDPTM9I3yXjHVQC1YIAKtGg
4FF3pgkD+508yZMhhoLnCgakF+K73ZomqF6jMqii/8yAmsX2huvgQfhUVRzF
9aiNqMbUbdgR111a4ZiVRVSZBxpHJXXr2fkAasEmS7EEkCGr1Lcn5kD9qCsu
4X3MQUhX9PIpCjWZV8Td7lRbecwnET5+WYLBVQcM2H6lqeOCfRVD6Pv/4H5t
wdaHu6DkCI1Nhfx2qGoDRnGMwD5+LjksoNERhwdSQ8q7jVaR8h4oFCt6lBhx
DaW89QG6HlAauTDLSoB3itZgyeuCQT/fMK6Q6GwEsthaAIg3Lsis/2WJMZ/K
XhbmRRXlYaj2ePTqriHAUaoPAJKniJStVwQ7khc7MIxZuLe/joY1Na4fD0C/
g7NodxYH36otrWih2j2lEHo4cEzWAnicpUn/4uBwqic2Ym53EvOI3+vOOO8q
wWP7//ot/HusVBiw08b5Xxyw7qDFr0dOe8L3cU7THsTxc7xUbCbiQCOBk4H3
JA9yrxL7fG0MEO+1J4NRYsjMaWSx2hGLyDlxLtYZ0wAFmJDE0f0zUwhgYaJM
S8tZfzVgr9TeaSH+Mzzvq/8jPfMaFQh9DbcD0ffkIloXNrHeHYSrF7Kh0ZU5
8TzmSwFNdyFlkYN3MrMbpFnlFZ5my9d0hSjojkWwsQRlllHvrnE/CXn3OH4x
Xps/wzv87KMxAxZ7Ap8LWrq7lEHmaFDaLiwQ0JGzmiyJPtzSj5bAUhTYXdpg
h/LyoZNldcEoYFjJJib4ndCbVLz2TFBRGdk/RINrrCn8k36LYlDD9y5CWLZb
xGKfqiu1kpUMWSZuCnhpNupny60htH4Hmwnj2ygHAQqw9qlzdYhkpZTw3mxp
e1Q7aixDEo2x+BaHLAmsFIlNNaf62P3t+51LEQfp7G8OBcJ4A75BtdS2DthX
zLu9tYFPN1aeDpDqMFgXhTz6WWRrzplNb3QRcCno2/O9V+B78/8wTo2Xd6Fd
iLCrmeQG8ABGIGReUCKwgRJ96r11eKQ2/xbzmf8RqO2Spo/v1hFETtf3yNzo
MM5L26zQUOHzRukijZhy44FtxvECKiCqnWcRIm9TVKHKbdk7LvPFcBdG52n7
kLGOC/kLUXOGJdAY/BzkPO6Vs6c4T5tjt69yMC1aSfykr0L0MspMTeWeMMeb
9U1yMF7nXatXXr9EuVTNPvTHVJ+i1w985rKnLdxq4ubHZitziRfqf1FMY09k
wxbureqq5dmWTrumuX9Fki+4SoaOPJ455RwP2id1akWlcg7OL8DcPymfCTZ0
HV3SO4Ar0NXkU5bAdaMWAGhHqyI9YdJkjAeO4OfudhQlm8bFORylhNx1vDgx
/B3Lsoe+xiKFOfX0u9IjvLJxLUAolsf5yVAxHs9K9X1BVskITd4p1rGM2DNS
j1iOloEdOnoeqJzw+g2RPlOuvjckeL1PPua3nArxxMb9kWwncqS6sMF61a5w
HN1FITYnval2uabQJ82/RTQ4QNMGIy1PPV7NBeYb5YtejPtY+lBvKClXlY7i
bAUVMuv47e4Ka+X68+y0m8zTUwBDPr5jDS3txs5MittaVLOjWXtE4JXFgnoF
tRrWemstOBDhcc++PeBArwnfmBg6CjwUq2XcyNj7ubm78Hx/Po3EPehp/w4i
9Q/3kEYtphJPsU/YpG4XRTVsnR5wN/rNgHiUgXQeGa6Ij0yGlVX4va/kEADZ
+ZUXQrofEhuYPuqdpQiu7Ylx2vCeO0940evL7r+OIfR0x9RVTyEiEZuWtdun
sGFW7cPCp6O1wISU25dZT8ORPYWkO7mtr9mfbueoK6oUXMVNYpKWycJdSFFI
3OIwpkypNgfu8SR5oVhVhRj0th/9PCwBZAeWLaP0WwHBI6p0wJX+oH99SJEp
VvZJ5B/Mde8v+h2TW+BeYKMpdFXpKFuI82kHVwbyj4TUaZYaZHx6l45iTF78
SdCOa/ZnwfauH6CkgBwkaHVy9nnDfupPgy+TxSGyvxyS3+N/jnFPnf/Q3l1W
vmNQ+LbkYTlrkaCnAUZUDCnSXL6dOLDHP75PO5deBMXNL6otnesd09uomQR+
OoGarZVFIHV4X8m14YBy5JM5+6UaLlEFI8mrWOEmmFmP9wWNwsDaZx9MjQVB
idgHS8CMZ8T0cyLY5RuGejlnbQD3MTVqstvAdxIujumMJ9fWo9VowA2wJ0Sn
a0r8ufK2agM/W9iRZLonnC2Eu3d7BB2MrztnGdQ4uW7IGXpUAlqFdFbZGZa3
/CFk4PnCUKL5KD4nVOJeBgCF2gaIDEADb5keyg1uN8IPP64thLtx5fSZrxXI
d+sCQkNJv5fhNY/wfME4ZuIgTqiSxNdZw4yz3NP1Jl12QQ6+Yl5akqxJyeVA
2UyYVeVVYtbBXpgYYOe+7efRg5TecQHBIlf0aFpu66+6JNKBN8SwIYc437SE
GB0WPP6tKzeWDlZ78MaFnLRrQxTcj7GQ5jNjaXwmNlB5DCKW8jkw8p1CC/Xs
4sPYckQhbWoGrRRPg+G0CRHy9BZqzdey3c4BzFUgW43Eh18ky89VS2tNdQk4
GbF516I7QHacCJzp8rlSkunFPXOxnhkq8FO1LP30qDpqUG7Wl0XC9ZfffHXl
P1ME4v4f/jx9aVSf4EBDeIOsb1FO18LVexfMVSYIF/ZibSMS08KQrQvvW4v2
HDI3mGY6yJMvcQNRNw2hfwBs1ck1hkdX9AKL8NA3KJNAjpeX8lmo265PdciE
c+DFZfUx7DiLiN5UKAAauPLAmpW+lxEW5C3aOjh/dhACIr2cW/aHBsG7X/a2
OODSUIh7UyDOWdTsWVvQl30FEMNY3b0HTy4ybapMDCssPQ9VZ+spr1Z2GkdZ
8lNcofl6Bxvxq3GSM/1lmVv7OctHW1+oMJa5DjX/B8dXW7iegCbGR9UMw/5m
yltSsavpcqA9Ul86V7X0BIFinho3aoX8UoDpx6IaL3vAvpkaPce27ms5FkBn
mEZQW5YZ0OlJp0HpJkkfoocAXaqsOFC1cNew//iMciFa4sJtUBHIuiL1eUfM
VxDiuRHIUmW3cPkTDCr6DG46Lq6li50JReAQnXfYCdafjY9r3LyaaX3AZ0cT
SkUGxu9BOcsJdAJLv3sYkR6HZsmsIOMT/WDui/UM5HHK6jKAYOjt5kk1rRxU
2Smwr1j7BBinrPt9Ne2rl+Dxq9fFaYFvBaRVR+ntxXuL0YnGRmQApSRmgZE2
94tFU5oAE1+cGUcI//hb+0lgSXQXlVv9Iy1fiznUqhqq6WUEMMgIlDhSxdcu
SZfhajXsUsBtzTct7Gg32WeBnq5IlETeFpEvQYEcIY1TL+lmsGwkHLKa4QXI
9ag0Q5RWdsOHHfLZqjrE4pe7WPGGTNW9g3mPeYtTCQ90Kk4ZL8CbyLhAeaJo
OYFKR9fJKF69KU+uNPt7M4TH9gNjyEma3RGr0sxwputZ19qCiu57FVrr8iUJ
Ph/4kTpfmIOuFfXPQJEJ6uFZtwhru118INWJQYU6or2eAwj1OpKaWDdpli81
k7AYbifppRC0qCo1b/M2JfOX6v7M4YqxAV2OvQAOKNbUWKKdu2k7BBdR86ir
ZgHnmTXdjNyQ2baw61KMw1RWtpZSZjbLc/I+kINgyZD9heirr3IZgb54Ni9z
i7ss4Lh3x2oSfQKAEhHIiabnqpYvY4IG+sxJx45Di4JuOABkH0hMx5e820+B
r2+wIjgf0+GwUh/QOziI0vIyxEIz+IwzCj6NrnO3oePGY7EPnt1gfju0/3wG
PxatKef92NgoZjePFPWLJOue2GqkttcsEusWtXvnH7gHYjEVBjnlM63+7fP9
NTUhIOV7Pv/KnBTLexv0xOHe5QUCt1PzL0ZC9eAzWwvJhDp3ida7byXyJf9H
wgJ/2h4xr/6oe2CR9V6BoXaipTUmc1gOxbLq5vHZGwr0BFZv+LjUaR1jRUlg
MOCGzn+GWTiL2wZNicigmnS5ADJ40uQQgb8BMcni+H2i0pL7a7GUdYiHHM82
M3U2gBeCRe7hCkgQz7LnUzccMClag/kFd5ZGtOZu4N6qYHPAjMXSnf3gwfKP
KxyyduX5tXkTYvu6UowAoSzpwI8IfH8qzVf101/E4+ARhiR99RZn2oySu6RM
GpM2pvpBcjWM5QOsPve0Q7dpqfRHj0ddZa/PGQfRPmsoGYd46PyK1nUedN6X
CbMYSNQ8CE2Exlzr3LLaEkC87gy69dFfFy0AKpNsLpDxpF5ajIK2MV0pbih1
Lhk67Aha8/ZjJE7lPUqFrp6z5KXCaasrN/L6KyKA37VuZwFIsYtpcP7KoihV
8cRcPD5lhmQCGuoKVxmxQzBy/t3mbTT649mOLQb8w1cVczeaEvGojsX/InKH
g4IuxPGcIFjsL2fEj0QCUqJos+GghJ15IH8dpJQkFvJfD0NNSOwVfgY3yeKu
aevF0ZnY++t3MvL1++mzmoKN4RgQLrRuhkOrEWJQqGeCbjy4Thrq3TzBkkZo
atYpLayb/kZ8SkXSzUcZcAgIBiPFlbqF4BmpvC4TaYPrRx1PMCKXEZdkgI/3
ygs+EMUHXhtSiBGk5fIoO6MAbJGjwXWj4qrYndfgPrJq6WkIok0lWX70eOm5
Xf+KpY06RtL6C7x/hKgqAoB4aUOb6MNFApbEYBce04C1UbYWQRuI1vyNJkeH
uQvjeDRyaODuah4YtLylvKVbMyjtSmsh2Ftg92ZSyQvOEEjOSp5lyFz8wl0n
soWm6kc7fr9dK91QaYMjCzUqorqW/48WFuuHfXDwYI7F6Gxe4uLRbunCYBFr
55oFfcllSZ0Ci+smcNfSJj9WH+S8AucG4TS44NzH99Jck343yKaNozSIpDRA
LeYdiIp4uHWIFmF5J1Ur0YO9nBA7DxdUcQ4mUoIlWi//3pLlW0egJFEdzWPe
eMUz95WZlg9u+v7TcSKJva5/xoBv7t+YNpKg2wr21x5E8BcsCHTvBvKVEeAL
XSP+XZsc+HyEMK9aoJsAM6t93zO9SNn5qolEatGyy4zfCOkfqgV60oTHJXXh
SWXwX2OxOagGN5gNU0wc75Fk+L1BGxciVEX8vQy1VOWiv/snk1sN6h0U3AFn
pfMDvY5bOmZ3N/0Yn0PaF8Gbcd4wcONCc6z/xVy8Jjp2L4NIvsyCnU5MUpng
sQV3FOcA15Q0RbWiefGGAi1fHtqvCAL28zHsYRoUbHlHs8ZTMcnP3KpUTdFT
6shwDDwXhpMHT/ueIqhbcHUQuVxCLXM+/z2UXeinyYeasVzREIvBDkF5qUG2
jH/+ee23SnCaCRG8pLeEEbKg2Ozu/QSscCz8D3+AbPGJwwb20n1wTzvwbu78
Y1pgFw/97Cnzfe7vh+yp4HpnjtvAyYVqEKN7rsBS7M1AdkM226BLjjstk0wc
GzoTh1QZaNFHlapMSqB1IVMrIt7JoS4h+8M4sfRUrgmkKLJmgNAO1GFDPxVB
vzkQGX8WZbQ5gQ7g3U5JaI54nV2RIfc7roU++J/wSfKeBy/2uFek3/0Cg3NO
KsaFPqPlMV7EsQX6F3tnLNWw1ZLMU1DPe+7aKuHoB12jelZd+D6j7Dh4aMsh
CfywTNOwAQl2uaHYCal9AuU0jK1vQrjhpG4wPz2HhToyQwe1vqs37c92JtgD
/8xRlOIIFcKiy1P9lzxxQVzxELqEJE2ckfWAtP9YJnLpSc2WSzloOezLB5gx
oYkbtnh8GgVlvQbwy6xqw9dJOSPfI5vo3f4CyfLjYmKicdvH0QYrBlnUVzEh
rO1dHmUxHaeWPWtPe1kYACZusVng+73e0UHYXK39oW7Scz0h1xFQGcosBbDw
9DK1OAOuNbkOULdUZ0EtUBly+8jMT4RWi5agzPsIxR53rGXLRqauvBY6FrLV
fXx4XjgwxXYQ9S0hyYNwk0N3LZV7+P+fAfqA/UqaXRhv5G2HSHetIjxZa14a
/mcYEh/Z5ZOBbQUZjBGL6iiI4L4gxvZlT6XbVtxuYQkGC4b7gnLKDg6TrvNq
LqP0Or7ws9c/xjtoRdFm2TLIXDWQFsGkgY8A36lIO2UeG7XGq5LTXhQpsRIV
qRTYBJPypyeyR7O5QiH5MbEtsecQNHB3fksYvxeKfnktlUBVTp0MCTnmTgP0
oEOpCQp+ll8x9lF7x4Nwb+hHrqRzFCPuQzz3HN+38Q6PJGYsuKB7vejOwfIT
LjkaxzuYu+BWufMy6zfNpVxqLNnp9hOIMi8f22fPH2g9NFhGSyMvjoQePJR0
4M4SUwe686Ngf+dKm2ph1HcYeukpsjATKWoFWx136QjXVgUBUiSHCw5eV+N/
NF9soUx3vZXkYbYPVuKS7rrar0s+28wdGoVQtYrt3cqYaElYBcAUlk7DN6Sb
Xm2Rn0jkY+AmIWA0cU/6szg0HvyNMyAgb7Q4pkV1w1Vm0t7Ii6YJWG+8HWin
e4mCl2LRxEZyP14FNPq6jWhAuBbj0pEOH0CqmFYgD9IhvNiLs/nQdqqxC71B
8agvrj6G/oaZZ7I1qvYAKQhJ2sDT9cUyb6fDhACJmXEXsvH5N6FlPeE99Bhb
fY7yntq7tH2oPSIymFjheJqXiuO12kqf7+lFmZXwftlJjAfMVCUNbujwPQ4n
ZVZ5SAVLD8n8lWNO9OZHR5lDYvxlyDiQmcLGTaljw0RZe4MLEaKhcwRrL8cY
ZZSbJooLb1l9gpgKFWhSP+jx3VOYCLFZGTAbFXct99ksSCvUYKwUq5fzXVhA
evCJ5lTHzfQn5VRu2dp5Q/5MQts+AbH44Vu1pYHE3gdhriR47nfvnIhBOnZ1
ccDACI5E0GuAODKzgaQwP5h/T6RWfVzKtRFvZ6mFVx7sKjD2gXXAMqMpXeWh
7WFehaZ7EtAZ4vl6pIiu8rLuNM6yHeGqnV5OEn4o29p3w23e+dyCv9Gptd8U
5CnG1xQOwZE2kuRneb4Ss9+3r0z3BAZa2sUNICpwaGIPn/iCytkVNmexY6kk
yuRhbyAzrDfj5b0FVVqYRhQI9J0XJhc54oPcTDiGAGcK1iKEo8ejZYWOYvhZ
wwU9DXOs5kiaLHPjDq9ypy2+cViuhKHffq26+6ctYAlLXuOegvD49G/CbD8s
dpHRr6c/+TWheRY3sYl/L8I96B1Nk/OPXd2m7PTNdcZO4X67swAlT2Q7mmBF
GuxqAw3EwhnaUcnUsdLlxwdRSQKvIT/TpA9doKolTpi3RZFyrlmcliU+WnR5
91haoWHAtpmnRQrnmLCnkNYG2aVGL8CGXLCeN8daK6f0RhdVCduzKrYYhWAs
t0Zv250jpFJMAPnRNvpjZegLXqynqJZpSvEok3FyeX54cY7nw5gjo7hi74Ox
7Zx2LSc0+hzWd+6McSFTOu047HWku0iwtvJzLzSQji5FKXX1gSJUNQzUeX0c
9mOu52nn4RtfqIqXd4fOvf2Uwgz389ObLACTxvluxq6jpGG3t/kFOaLP/qhS
mBK9L28LwLuAPIypINg5QF+8wJvziOC+vD9h1d/s9aQStMDVw4evbiQ19VGR
XlJ+TRMkeviCWHTgaxmrLbyFItWaxeYXC8we2LxD59PCD1iSm0/2NJNhDsvh
VT8H0YTknNI8Gwb1tbSPtqcaF05CHRTvgxFS7EQ67EOl324cbwNelMxQFi9w
OysK74R3C2jPqdFLuBeeYjqCUWYKD0sHdYuYJbVYWv2exNydPJwEknGVVVdo
lYShTDFsMOUweyeh5dGkltE9ub1uZmUvqpIJdSntXsbLlr4mRJ3/+tSNY8Yh
rI6+W688QD4nLkmky4GjtYmODBbM8TKlmUovkkRvVceIi2P3zoR2GZIENZzb
mNtdUng4t9rG1KifLqTAEhYHmEUhGT+uDS4+Qa8OI8Udw7dF/ypd0p79OKTW
aK2Drszh/r6GUAGvzdrO4D/rtdr/kIRoPyiX5D0e9MZJ5iy/+hpIHDrl0tpd
hpAV9t348Hpshfc51B1zk3PbmYutu3NHZa1yRbcplNOP0NZNWYqyWEUEb4r9
Y3ptPxBCsLV2C6jJAKGpCsUHWk+mN6MLbJ94VxrqrdFOWKrHJbGfF/3C2g3l
WCuHYd9+e6x/0JTljK8itHYJ6r/aEbdttPR6osNNVKRGuHfF917eAWD0/0bC
GiOIXOO3F0sROLbn+3eXWeZDvsFYoXhOlEijEc8xSarHlYm7ireTeOoLvv6S
RNY1T0QQxEamwokosMnsY2KE54nPibV5V67z//eRj49W9OuUNAp0dUkLZCfY
xb3Vk9EtYdyZpDPt4ACrf5Zb/WF3gGIOTio9yjdAGXtp01rqr1FjUOJX5h2l
Pnqno6yz5/PLNH3Ry2rRvVnipXGVpy5QojcgxcGCB0kLjztPmw7cbSZ4yNo7
bTQ0DaCWuzJJdAnjZOxGzLbK7fSHdPmBY+/oaNl4ac4bLucjOjKfn8hCDdrS
PuYxUynJZPBMWKfMPTXu5YOK4lT4mWJHyAesUMDhBKoZMTwuyCmObud1OMQd
Sh/bK6PIv6z6leGhSwzrG4F8GiPtLv3GbpH5glC+UnzSq8A0X/81PilOosuj
Q7ZAv1TvejFpWBtdz6I/RTD4AY1ljeoK1tfCh2ChYFV7tWeFoeGsl8yrMxOZ
1eyBKXQ+7ECNbXtsvU24HEmqHadiqyRmU3O2yIFzZ4Zk64pTkJfNR/m04FBM
1iX+sQPxphRA7L6pjFsgvsRFmoyKaDEqWUfS6yIjQca/RPLeQtJ2MsiyJRBW
kCgSt2soRNfWdfag+LpswKZOu8Th4pcKaIgwR/hqM0nqnlK6kMBF3vMe/UA9
FDRZPpGEhHbZgA6Umj7ENvuMJH3d93dmoc6rnRyVhRbQs5HrGLXL7pkSSqyz
p12XEah3+7PnwKnjAX1F9T4X0yKSBhbXxKmPKYLqPs/Z1M9wISXjzzpReDNx
9JJCq4R4gDl5dmUCWL5pl7FNdYqTIPsLaZbK65Y54LHP+Tvhx3FxHqhQksl+
6l79auxabl+4PddH6NKtPC4xnLis1QpteL0yGIPTeGv8hsn647BD67TjZN4n
FfMeg3HUD9ArQUBzKWc8hCkU9O3IOwisZK8onpQKh/lTOCk6pENLsWpSQu7G
dqlu1wP59M1XAarz9bQaB2cD9y3283rzxEY+S2qBbJ0GH1zRfbtHpu/JvsKw
prQPo1u6aiu89pUfKOg4hxvsdQcfwJwPVuV7IQm8bWznPLCEKkFEN/tzPAE+
WZPnikA14y0wBU3IhktKcylhSeZCDOo88CXAoIfvjhmKpmXtyj+cbLIruWjv
5g3qOyoOQw02aKP1zFmXv9V8IPjUKOeqwHSEXuN0gXEQYF+QD2Tr5h8vzFU2
DlEc4B+dXYpNQifmJDmY13OqUZMMCTSe0gIGFMLJ57kICyVvpk68vpmXEhXj
b7Avk/AkAbHMSfDgTSE4ctP+iVou2Ncrwhu36ua8pLBTnwkX00rFcC4OMVlx
plLTq11e5uFHw78PcYMCTbrkP5ZzqaUsxovESAdtCwKmi/kQ+RBr1SIlI2wq
oMKkUwvsOTU9maNHB5VuDMsT/IZtgIM902YZwAOE8WxGOAiZ2VUT296GKgCX
0vZw8DBmDglmSIMAZ5nqRqT33QiGWxlDm4p3QReux8Im1vquxEGpHWrK9KW+
DJxDy9ZmzVn+tNUM5e1CfXcVJ4FcABahw57wAaRE8zjciKUKSbGXr4GgjX2O
dKpV0N0PaS2tljP6anXxvJIlMooQ5YMYBPYYeAw9lledyGBjNFL1tyQDKgjf
0XwiIxpHtU/IMGeiFZ1X+KVdMdEaKkDo/B36BbISwWmgv8tz4K5BMZnEYTa+
S6Ux7mDPhfUaJTsjp+Bi/LKyZNXO83vXyRpUtsD1HEYI0eXS3HuYMMK2tOhT
lXCaVgJXAq1yD9y2Tgz1B8uj8NszdGwgE0zogN5WKrFbFOkEAxYT7/1r7dPg
S0NESSQLwWGjeZkdiQHJvVBIwPbmthldZLFhUCGFGC5vMkvOahocDU6cWfIK
KmQNA9uyRWxzdufhLRGKJAQO2UmRloF8cKIHhCK6t61E4HPv6kLZ07CcVkvb
BYtbXLP0gYi7M6JeWhiweoN5fHhRHzH1WyCFCUVxcBwjpP6wRzTwt9MKpdKC
0vSLEt2d9goiFceFZTzXcVlgym3MtoPDByUGS6EDNPXu3xzLM2H2n26rxQCj
uqjXlNFuGJ/dJRnGXM62fjYId+56r4ZHnL5mwgVX52MvRMp503YAkdMRf/eR
kD0Q70W8kmXHDRM/P8+91+gJSHiaszaHqSW34LzduQ7kP9ASnseS+ELMxHys
IYAYM3RW39p+R/D9z2wTugS8Iepids+0pvIrMyfbpJgcxogQKMqhJ7ONN3yh
NW8CBAL/Bi8xYmgTa2Fbc2Ry3QiBjzBNV2jBncV/sTbfW5xyiLYEvlCUy3hI
Ea2K5RuiZnjW8+LWBVktGISjaxJmfXXcvDA9xSJ1Fqw1hsanW2IJAYriqfDy
pY6cePbVOoGhonKDeW87JpBl5yljq6pl4/qQG6hk1IN61cWzK/FEaJRjO/cP
zYKImO8GCnuXFGRjiGW/lACUubd9wxATWPTTfcYbWubUgbq7fZwmkeeW+qNy
33q5yCb6tqZBkmBrbKNIsj9g91FCxfIErrP3lnKs3fVckK2R99oYj0MG0UUd
t/XMbPh+t/so5bTJjRchu6IozOYICA/jOlvbQc2NtTAJc4Mou98mz1bjzNwh
L462nByNj5y68OcTuUhIAmgxSOz0Yap7PLP6r+yTT1CdNKx5lssdx/khmCai
Y8Og3kT8CQsC0J1A7loJR7NWe8wEkS6b1gbkRhlttJDQZxCa5FHUqN8N2mlG
8+2BKrEXqcdEbzSxjaRyhJ6G5td4ef5jpklL13WTFbgkVWUPhdVvv68t+dky
HUGnTgS+hfzlIbuLXrXWcvqQgCy2flVYYC9nqgfjahLejLVtb9nXOPGQyIRK
kdloKsQBrmMv/ZZuFCfrN+4/lvCXCMohDfEYCwfk3IMb3AX/JVz+dgLQFOSJ
1B33c2V4ogB4qfsYOP7We/SO7uKvHBKg8k9O6SHVGtXVvyDiBAO2aZdx5EdL
2R2RoouIMPIZWUDFIArpB4VNtqpbOJaI+j8GMxavVblKRjdMZubQQ3JyQoG9
qCJc3Eam53AmHlJ0J2zb66eHkerz7E3TbUUOYqE4S9/bwZUZl6Q7+lPDGuD4
YQOJIo6TR0t/550Szovwqgx0EqSHHZKrni6UIm23qhNB49L/A3Hc7BSnXw7i
rXHSxGpAOWxEKukFeIIjPSTv5yZ0rZdXLQbHVys8jhuyM07dyLRnC/2+SwMR
K3tcPUkSbHkqtveDh/SukBEBtd24mKG1Z02r1O/Godlbgfv3sQ/0umOUa2ew
hVwtU1dqGxrnljeOrh7p5LyNsVmTM+cKf059vJmvioQ5gZZEW3STDT+Fv7vr
+0aCx48omiHI4C1kDQkoWdUWgYiAgnT7WQunrp8w1IFV0oQEnVaSkg93JxoJ
PwA0BD9shR3LlE6kx+COpp8sjt01xLE1a6ukyUHrWouGZ+zIfLpZo+a5q0xq
ZhyLBc/8lyUq2jhon1gZvL4qetZp/JdKsUZW+i4G7OfkbAtgpqvONhLPQ3aL
A73rI5uxJ7472WioEdqAxlc4c0okHcWJ7L2DwHJecJeuDlhxycMo5lDDU2Y0
XVZE+ZAN+SyihEv2XBVVj4WGuqEcPTYk71IWd9rAekjPjZ30IjsuzQpuTtj0
W3yYOKY2OKQQNzHewXiA2VsDD+Hg0IMehbwcrtSmIAiield4RVKtJsu445Cv
GzsxV94JcVGWmN3Q0jTCUa6HpkO0u8FkYNeekCB6i1q8jbmsOMhwVJUVaZXQ
bO9LzRz5VouWJI8QSMhl883EdfSS7u7fGMe8+lbPXQPTOaAIhDKz8THnkEac
QP22PPleNK1ZtrfP7abxjtKUASEjba8JG0PheaRqbzNlpRRI9c530PaupETp
bI79EsGY1rzfa6xsOA3X77rMdFz2y6Jhyv3qw0n24NG/MUGmY/KLmnVOKHWE
ipr4dordN/f4eot5iLZYNFS5avMQVjFo2WHvKhoQ0/Kfny8+XES3YBwwV2TF
gQ2JUx/hjyOBzhxtaOn+zj4gV7y6saIT9jypS7mgdVfS1uqCw8F2FdtG7g25
G3Xch3vBPa8BF6FbWfr6xF4/vcRDFsc5p4Fn4ShQ/MyCkOxrToycs1I027cu
/gFkdZjl+PlWXVXYuNsu1oF5G1jzAjsvSfuDrfA1euYGnpmGtTu/jY/F9ggu
4a3ESf3WSgwGklpNrMvj9zUpt/IcFVvHlDTCZZSt2ckZKirSDbX8+WtGoh3r
d/xpA/B0tS7hFTuRM0ukt+5WQHsqv/dSuTZnlcYQ2IHkCTOeQYpVo+OgEgfr
QCbYuC481JykQ1hyAO3RlHO5mvrm4yi8JhKIiHkOXZJfTJiYUw1jteDWKkhc
iLEEGlPqiNOlLdYj2dAN6WIZQP5wFW2fM9Wd3w3/krcJ93NlU9YxYRxc9xHy
HF1qyuCnjlIhjJm07EpDOH6HMhmQn/XGysjfVW0HGJqRQHfMpc7aa3T/rS/w
JXQlWvXm06RHwscECD3kuwnU7aVxTjvGO0Kd2qVUWLMwBpqPp7SaTQ7dci/o
UgSqwhHf417v5Wxopfmgc0OgtiyRtdO8hFx8LXzhdOojtxE3x4z63HYUwCD5
5Bj3TjBmz7YezNHmdeIGp3EfegPdzlQMsguuSwbhd/6H6gOhfXZDcvqG4+Nj
t1ObmDGFHiVOWsW8wRVh1mVC3HklU0g1x0OxYoRgx1CjkTxWlby4ZaJuR2pb
8Q5cAa45MCRXIkKFTJ7GbBuuhlfpLRQQ/jXg6Y1PW5COJIQCPH8Ees0J45hO
gvr/ZkZy1zUhcpsypDD9VsK9qI2glvViQ5iGa2Gxzqx/spuoz8OD/YmsBSF3
PdgzAXfPOUhqTprxoG8Y6cDk/GYU/z43dh1xeDcviq1er2SBchoDEQU0FTZe
mlmUjcWRSiYWXBgCzk6R7nwCQKYQplMUZJ02uD07hziTHmim9mTtf/LPRTNF
Danh/RlIbHGPxKr/IPZ4Cv3Rbo88kGsROEsV5JQKLfaPCuc8CgnuiDihmVtJ
KddiUMoZhe0xfsp/bhUAFox4ThfI6eOT8FMMQJKRwhDYHb2acXksr5pMvory
9Z3Le/EKdS/HxtdW9os2H/ciDZxhtzQ34O0gwmasIZz3DEj9CZyJSw/AdN7A
tdnfCb4w3FQYeW/a/OWWDXgPy3XGvQ6Xzw0U79qVUWBc/4BmJi88Zy3PAJ4Q
VkTCJQbjzAUoHD6z2MrAslh4z4hGOPWIoPkkUaGg3SwI03Vv58ngq/1a4kyt
xBsXJTpXSJ1KUxXmOYwWinXwhvPikctqh6+1LaEwAxnhbFz/7qpfAKOhp9Dp
5uwGJXK67PIuzEuHeWoZ1DFPxLr2Ipd52YJZkZvoVszyZzknkscbFn9HU0Nd
o9pWRGp3qIeGZXoLdLQoRbxs4RQVD73l5ybi8H3wsDbGSFEMi8lzzlvHEo3b
P9qUWNYI/ae0g+pqmYCfUnrcQ5u3j6BVYJ+vFC6GcRpH7ro5sRfp516irrVt
5jiISf2GeRQFmcf06PMnsEBpkkiP8nWIXZaPvwf0EL82jj5XCazabYsj2wcP
jxRq4BH2dLdV6+bb5Dqvw0MVeI58qz2J1/8MvRFaE2ohkjUoV2NDhHfEWROl
yFhqE8t7lL0VrynIC532tqgkMncUuzc6LBhwlnFSw0M6EJ3NWW/jT1PJj1dR
0pTFUmpSLQ/BvgTZBW2ypmHx3W7qhqRuMZ7QZt/YpbfzJaw1lktR8JYv+77z
pgiiu/5Fj7EauAP4yy1wWABVA4Op4jackIv1EBvQ1hDJDKE+UKyeTNF8TPTk
gGvYm6uT4h8zsTd5poj/vZjg421LVB1UlhiT4KmYlpx4jNHFhgkVR9+mwtlo
Inc7V40+Le5g6JEH711X/L+gRdVjNTDKOwv2VKp7vPV5xN2sBcojG8EumdwL
oU0UzpYq7KmOrVsk0AH7FHIssg8Oqth5EeqUzTQBDwP8s/4uHTEgqFY+Hgg/
XIQdwryqOQPmQlepCKkcsK5DUjb3j8oZsx4G1dSHcReytmZyYF9l1cb12bmE
ofG6o5Ojn7EoGHImO8j1kh4wqfPo8aDW9qtkHLFzLUdRiQgpWQRXu4lbeCvx
xvTy7OAdw0n8uaz7x6a+p10LqQ2Y3pbnxisLvOsS85yb6FZBeW7/Sfs+/iTB
ZAwHSH9CSjhhV+yf8R/ef+aKNNbhzsu7A7IXbWLXVV9NOyhROTLhWe+CR6WK
xRGNcRXDpbfxofmIQ8CSmJKR2xKH4A87f4KRZNC/YslO1cT5YLW7H41tf5Rs
MKYpFWbT6porbNn8YGFrT/em1dfnND6ARo8YB7hWQ8jWpHXRf+xouA6f8ysG
7YZyO3Lr5bTVY2nrH+2jrbDMiB+ee4enO1J5A/QMqWrsL6gziJPmHG5dktmV
uni5mWJAFfXKC1ABCL0IMCEVe+prl6uMrebg8E6SWud5Emg2wPFlYa/5MQoU
CM6sunIVmVs3cUPxow8fBEQwrNuyAdqBVpzKAU0dSXEig/CLaUhAGO5Mnc9H
zsvufq1R8UzSCWAo/2xZMIId53jMvIX7VWDAHQo39AGDV4I3y48lhC/WDCyM
1EkhWxhaxf0uzvhFm/quiVUvx5/EQZ/N361ugMcdr6off10pRAFvaM+EhmoU
Pk5g4ei3JKeuA3vKC9XOAj/mtYCEBZmD0Xg8kViM/y20nMl8ywd9YQWt5+Dd
MdbA48Dji6tahz6KJPNVemf13JPRJUnPYg2iNUMtrkrzFmw6jVgWF5IY4pSU
aDXlBdfoC/x+kwSBpeAhPkCcIdeSTHU17oEs92rpFDsTYkas2mhas6gklm98
2lFLtwXCLns8KzdsSDgHCchD5XYtxdrRmGjnegNMyd5bd9WeOlBff9CTdaUj
5dE6FZF36Aw3KB0qyWmAdUlAjIykXcw26bazpasFT8PcMFZ1mD+c5o8E7xAR
TWEmrWp7Pad4kFy1mttLGjvkR0QW/L+m5riC1EaHpHMDsAY/Wd4PegoJ7aRp
HhN/3KInlLepEnQktoAmI9Kab7rznLCXI/zu8PM9UKKIWm0oJDCp4trSH3lG
kzg6ZnbJcJTk5IaVfHkUFOsXOLZ4T75vvYieaDorftTLhAy+ZMqCwnH8UmVQ
vCIrB4n3nr8jl21y9ykSUQ0nOmnfpyXwU+OHHtpBMfxixYWhi7KNkaDEATqJ
dgdKLU4OkQgWCKHGWwJrv2Uk1m3ADD3Tr3SKWXYzDtfPBARXdNea4WAMuOlZ
tZZzvws7jRd0mMmqMeIg4GJqFrwE9IZvIO9yYS0bCzdHgh/0njYB5E7cOHQa
WcOgPZlywJ64pz9DziHU3nmY+X3XVD+yZ73PRpQWvJgtilvXjmKJ9Z1aiS32
QIuIbRwytRXsKISOKajePJfQFKXqKqS6pVpBl/RnlDnh5KftVcntdHLOUvhR
iS8WFkgrJMBC3UnvkL4C40RxTPTyP37m90/zGNT68itJmESwoY/OkQ2r1xxB
DCeJ9VW5svDCdpUVcDZjvAee7hkRUa5bra4feoQ3HDne2RMxleYXVSgjPkGr
pAP6+qARowBO61bCvDTng0ZZdQeewwtv5ivnN1tsloH4mtnNFJOrOqHWmObG
Y2IpCbHyCCryvtd8gnUj2/qTPAHFLIHw7N89Ur/fQd0CSM7zFX4k5KWfawz8
nw2uUKpgYvKZrEOrICqYwRyQnti4u15SOVelBlAYDUJoClK8AckbZmj68t1O
qQSsvh8TJPQfWuXFF5+b/7Xbr51iUgt1njpewJL1FfK2APLA2h9MX5r8cKyt
1Cf7mxia80HClv/f/VbmnLbVVW8O37PfEhBdEGZu6o8CbFtFD3mvZn0EmxP8
tu7meOFbGYj0X+0NoAsrw0UQcuxsO16b7wMlS1wSXx2FR7/fhiTLa4/EkeIK
d7ZKoNc7YB+APvZh9kQ+UzcP8LEZfbtDoomj2k02kAMvFpFcAImbMWEpjG7F
9dogn+N0GVVgPnQ2fdz9k9QyFNdZvp3aRHOmu6Kke8UUzhX9kUvse8z3UoRz
/rPB8d0bwA6Uf3FousmwMSWKRSAiSCpnZsmymiS61A5q490Wi0FXVkGFvEcx
CJJscOkj24bcZwtpBqLtRWZGgbGeblhSZLb1bb9E9APIxwoQ2Vns6odXxCmM
9sNyUEOOu0W1u9Yxjl/IaUcxCgfsHeXTpMNDafOrhgIMjTXEIbS0CzAxHePn
oAy0l730B9FmSkk3lR4Uy/JgN7Ykso21FjHpMFXvqoS36cP9o5QhOWOzYZN0
QK3Va8nGPgbAeQPD1ITLKpFmknfw8Alm+/3i9HEaMSVJVhPQsYVDMOdpRnFe
my0wLZ1V5LAr4FzXcCBWvpe0pgI5/eGm2CTYPA+TD0WMA1tAdehjKnBLHJE6
YlOycCGcFlhqpGMTE+ZEQt+EEyMkWecp85YY3xunfuvhXB6/MY7qSPtjvn+U
8v7Y5utMSKH+oultkSGumhNmWfQrer5nWBw5wDWN961MEqAQPWFDFbONVlK/
bSE6QrnnxHiY1KbUYStVfLUiqDPwSDdrIdi8S2jsSJt6fcFzS3oubeNJYnkX
/yeKvSa8kj1p8m0ueymd+0wcSlqkf4MNX5V5wSGtaZKJA0inQShC405SQZMb
KBDdpNZi816Y+rmXNhYKan0qRGu1KBBrqSAMsy69Pr0RnRUmlEheTUM0kzTq
noEkRScToPlSuo2sXvLEys2glXaM0TtTxzFFNrMQ85gtFI8mxbxmvTCIbKcE
LWLuitNF9aIDOifc5wyZl9UpQ1FFee6vQq5fRc4fMaLsPea7lRq048vUaR97
7U5RKFGYVVK8AqLjVMQp2VbaTwbv548a0Ajo3BXiixdguoFKd0NbAn67/M8G
QWzStUuga8FDCE/YWi4nF8uTbo7BmRXdbfFdjH4NnjihCED7CzI+mrEpYmPe
ZY3pz3zYxl3YzBRz0gKlVHjcGsS/CMdDpl+FD+C7mM+TRx+Bu3jPd66lA8x2
50/L25sPM49iwQ8HpiG377u8I0sfuGdZD+5pBAzrc8cPK1NJFEoTJBa33WoM
3NQMXgLCVmDTXbxC4Gnv/zZ05F1ojwjtolel4ysaTYIrIxRnwoUAoPFAbg0o
x6md+9m1CFwfjfFEzKlpUUYfGRe/qCUOguHKqzDIG2gsRr8d5t9JywQgedvK
/1aKj23Vse8p78CqTcBz8x6EraldF+lnmrmQYevY1xHLKNMKtPKwHNIoA0Fc
3T7sTv1o9h7R981Dbllk9YyudSLEfxov/emaTGgLnYFiekCkzlfp8tJUsG/Q
PXi2OeJfQ8DJifXoJBJMy/r56Ul1nUfl1ZRIHAFc0pTeQI/dZEGOXDv6slXD
uxs8r5nbeZz3ak6ShHyw/t/QvtxcKqKIyfnGg0+50fWQ0ITO67zue1Egw1kX
OuN0g597c3ZV3wQ7C3pSkBlvdNPy9b9y0kXH5++hnQsKcfX+YZAD4/oCoE1n
5Om8FsBiXojH0+98HGu0flEamnxcqHYAx/QBSlvfaIDD0/us01dLhedZ2LX0
PvZRdZOMN0vV23pTFyKX+lUU16D1r5Z44KgnZRx9rSR27bjppkpyrZQnyK8h
zIMtnQhcdlc7f8/W35+gtT4iL9XObEe0Y5/zTi67PWmUQAXIwW9kOy4u5FXj
QcskpbOiFNsk/Mr+nJA6xcLk34B3tH17qoJ8P1OmQ9KvNg7kPQ5crMQR4Xdn
vhtXOn0EL7wwxl9XGvkvRh8eF8AcXAOY/jscoTUcQR/2zHDCm58EosnxGcfe
6fuho887wrxTcw9uK37mCaJ7RuxHraXwlCuJKj3YHtwqf+Pcsx0EpN+MUF/P
FErN296dapXBkyIbAZdUf9DrgaH0f2kXO20aqGs1GLaqruA0vXbDQbZRSaoK
WKznBT8C7zgY0EgLXVjsrfKf/4++iiWgFg3rXHyeqeyG3Kyt6A9o9qR/rbTx
WwCBMRH5uqFDkUCxe3WLl6hjEjcrqLSoTo2Cndmnn1v0esetXLdp2aRNphJk
prBkLr7QwBzqMPokHvpAyiJPJbMxAYm4iV3SEKOHktWVeU/Vh6NUdfYkRU+3
nnKU0as/QIItHWyteUqhuS9ni2k5Sw4Rwi8alJk3XrKv+MzYGI7r7tB7I+kX
9x0RSaRempIuXMY9EHc7+ALCRZaE+6dyztjmKE7UUBDJBi20xErfUzoF0kAR
cklDpU7e/2So839fiamNreCmMd7bVOW6EHDosXOoljliu/pBfjjGl6S383sw
2+OE2pnG3gpcTqSKldw4mToZo1IeNkDxS7qOpaAmfqokqZ5BEzsk2Idg2pMi
mQKbbpHVDL1qaN6hX/l7P48a15VgD3dNC31jvoEaf65wSeSRksSWiWxu8RDg
TS/ZhI8nYOZkL0Rm8Q5FfuI3AHZfvffFfruDPJuzb2e/dBt0TUsIJfXYwqnB
Or6fEDT7nh0K0DEZM+TtYHqdfaO+hE7BGQZ8sntCUvqvNZp8ptXV9xOEpRZ4
Eo8Vp72s4NDjfVVS+bRhhJMVb17lFzEw7yRDdM0QCNItO9aFxSnUCSge9TyL
0185s0BKE9mwMS4ACr/fA/0mU8GNj/qd6GiPmaqq31iKYhv42GV7D7Rjm7Xa
LKqqG5IbB7fkCr/2Y0Im3m1EPqRVNtyFtJACsRsEdeRyzSPsh8exDl5c+0D1
DNiB9ge8P4ku9Vl2btfhX1NToSySpRIlBIT3WcMVgGkMFUeWjwv30EoDPUTn
dTSDRiszuUzdguaJj5NDzPSkBmzgudJdk1brlnXb3zSaE1IsQZbRksqwhguQ
WZN40qlDR6FyHyjWh9zaSg8USHvF8BuRHJ+ZWJhbZ0DvibMxCP+CAwZErKqa
NzO8Zdl9ZSKxCx6Nii04dAsasFhoITPVFCdzxgmmCSaPaM+tZjypWngGGC2a
1eO0nZm5o8tgLCbUKB9hdajIiitOdXOkXfsJJY+I3xk5C2ETnrbnqMD1TULK
2qnCVMfcyMrP5JZ4UMaqsZugbREAF0ntnSOMzcoJfRIdo5tiLvY0fM/Tzp+H
nkiM82jEEuq50luTslBYdeMFL5PYxAZ5OscIwuTntyUgzue2qaqMLsTC41c9
2hJyI/Gsr/Fc5rkWAsIxusoFgsUFnXTDs4N1LbgKafrwCBSXgkdVpH2M3gQx
XnfzhCyHFhRN9vRKZXqa3QzSHHYmIpz52BSxTbiIK8ARke9Gpm0Xca0OqKJF
ktST/0CRn6EEAvU1B6SLy/95ciGtshxPN7jOn2Ck6g2YvlGFAm0OjxAs2mgr
3G4BzZuztMjHIDFOelWfj37OSec1eXAp3UUicJUyUiRC5rkoxtWKSN2Youyl
HtfqTq67lTMTEWvPdZLj7dHmMmtieEcEwWu6mGdQtSCfvcL1HsotLOy6ympE
nhRSsmDJnNhTc2+ATXv5DZb1+HBJtSVXnl0HTanzFs+eNHk90b0CvKLRENu1
+NN6kb1/zNk3Qh2y9n1DqT8ZG8VnqkCzkQK09tImK8Px87c8sXWtiPRvihLJ
dOsZodm4DdjHA9xLbaCNB8ti+yG79LP88JXxI6LkSyjlZ4Hm22EvPXqWvw/y
6M6tDkXPVrPKurycu3/5wA9z3WAflhhLlzn1+jzTYKQdWuzfLOdAstL7Rwdu
NARSwRZT4cnidXiDnXB5+Ve3BdgB32/xqf2tdY5+63hdRMqEbWarapwGdn2U
ZPp3nGnXT+mkrCTHGngEfspafFonip4HEkKxCh+ch2KYiGJVpMyQDK1/QSbV
DvD4E/gFOdjUUUF+ocfWFrZBMBDszV/7p1wQVskk/nu3IwG+OBjiISjq2+aR
2yS/AsS9OfDM1K2QTRPE3D222/3m52eGnO74WcSTibSAxmWaZ8hbKcOye3LO
KnXc2xQ7wK1UAnyfgR8v3nkYDX9/eFr7QBbG6F4MVZHsVz4ylHFar6LQqlgu
7kLVJzti+QtclHfPUOWl7E1PMHPa/1VpcPljuzTMUQZuEa6PX7gwkkZXmkFp
eU/s6rKgVW4PTY7l9BEuj14ikkXEL5v0c113oHBWwo6SioROrrGSJlqjy0xo
UEeXmb5BIph3RLf8Br3yRBnY4LjaXyEVNzKVlL6zXXU30mKlKaKF7xaC8Ep0
OzPAq4WQrjDfDVy5Pc63mualwS80wmio2EOh+A4lOP+Z0O4bSHr8izmWAyOP
X5yvsA7bvwRKlJohUlSoJRq4AXoKFDVxblaGJ9lSoXMNw5lNtDzr3ECaMPYr
lBbUZ+3VJX5LfawIuuwOtLlNrxprJ18Mcnamc9AyZJtmV6TARJA9Aosue+qS
hCxOH7hJxoh4nltT+voYwCEN/BycBJCnoSvrUhjgh0cY/nEjxnV4ZmtkPAOo
SU5QrWr0vHv4qh9KvvY2SqSVwjq5DEf2VYnAy6qHZaOifGZaYlHZs5gC4Y+S
/EnMKswey4g1YVp55GdBR5tISlPY0hHNnH3sGlPLJgNa2+l+2kaCGZPM2yue
kOl5l6SGMae1semeNTsL3gHDsGuBRhxhNmjWt5X1myDXgiXkVQQ2ma1V4pEZ
8gKEMVJ6ibRW9b0XHMce8pJIAQoXInUbQ5FnJOtc4XbakjV1ohsvyg2fFfom
wQaj8xLm2Dyz5AW6EuQ0YBAyt4q3AV4VI5y5FpzezWWyWwS6M8Sn2nNgUXAu
9dfpW3sfp/hR8mErYz21oSH39Leqf75+MKMmD/gAS5yTaeObd6MW7Q3WBPx5
8n6kKPj5GL/0QufH5DAoGnCP/APkZ5BTs4N6KjjURcd3oSxRr+YHsoaikHeu
lh76ae9q9ybhaY7J8npqHBiUjm7MvET3I0Cq89RpmC2A046EQ2B74d/EMulw
b/PJhblAsA2IerWZE0J8keLFwS9RPX7HYRYZMStszp/Fx14qsQKqbaVWhAxK
rXK4rhVZMSB+R/278ePVjMJWYpJ5KlJ+trw1Lbx1dXEsFhvm91+alcLrlrwO
vqCEYqeU9hLwQbMw6Gts7SOBgz7UU2FH1T1iaO2cbWCDU1TU7C7wUYJVcuR4
XH9kx8rqQqSweCk06+MYIvyJxtR6m90hFIf9rX6LYXFz2/C+ax6C48HXmQJU
K4R89dGI96Hn2Fr4fHVwLL+u0tHvCjml+P3tkF5fB1knUV7tAtJW1tGbYrvG
9lvh6Nbz2sD8hYjjAMVatbLad/3LF3vSlozTbA1P/fVzgXx77xVG3YrSZC6I
Qv/ncC6h+b3AzhuzXHvv85JUEJkzZnw5s98VbqpV6GXU/VmUp62L13nWL6gZ
7orawYmjRbg95b8cWqbc0GeNBfJQGy4in3UIqMOE5qlQPijccoh98dIxYcs3
DrvVIoLDRZx4hbusdrrEGvEXnoFbuUkXO7OKF1CSgV3BWGdHsykjddjtU6Zj
JmoWpyEdDkbymzcDuCdRpknZ8NSwIPX0JqqWYqM0SzyNDDiTPdbCPCOTHgBO
XIvp59IQLB1qs5ORoHSnkIz01CbCmNfY7dAMks74Pr005crf9EYsAsRnlgAH
TcYv6g2b+LWnZeCJEKddokKL8R/GD8AWShO0dyYhSLLxuKoOmNqDw1N+62CO
lLsoOgVW2OpkXUc08mGGK07X6xXVuEwS7kogrXgnLCmj/LWadHU4Ay+IH/Xg
J/fKK6Dh57oW3iKAWW0XKtFQ8G8OxhjCvBgRCQnZYBb3GU0L32yMgpXOFUag
2gbxJ4BTssHmZwusEy1yK8wHDeU/AVTKD3ZDVpPEgRFiooW8huhv6wvbqmPI
WKAJovALvJnztVFoT8tF5jks597HtGyj0fihE2m3IuEU4LfZAYCMqAuSxRCK
PS7B0jmrEyqTPXGzuDxk++Nz84EARf3Ol7LKdTPOg2Q5dcm0ab7a67c/QdZN
/FJMMEPXk5+APSLVyNhcu0MDrINxL9/TptlLYeItcGAe6KLhtsyTou9NOb7i
A4FBw8z++LeIsaYZkeS/as8fVONgTW9hZdFGgy7Y1PvvwhgvbHDQ8+lG/4SR
vNW8IgnTJP11SKiA7kFwGbnZ9t3B5At99EpsheXDAI/iMtoPPt8YBKgJmcWp
ny3o85qRqGmgZqo/W+8HZACcIRh0wCVgMF/rfI9BPTdVc0CmC522Xi3lIFv9
RVp1q3Zr6BWKjW0izshDlDH468Hptzwto3Z1dHoKRJweq8uDEAa2HlbE961V
sU1WgbzULISuXMyskRg7tOk4X6M0CV6b3aYy24FsxV4HoQDxD2J6tccREBBA
q2Tk1pMgPzKJqJ6eUAGnobl4hvVVwjf9ZXE3bQ7el0Kcl8PgkvSAJfHu+gOu
O10t7y2Z9lgZrcOg5qxRJJ3RbGjZ33CN7GjrLYVZQhu8ChpDtal2wjzAbgR3
Lokr+nY4ZqAT1xoAfK4044oeCNhR8QAqqYlmYKoSmxKC3zl//sV/G16+eamv
JJwUPOY5wEGuM8ob+jfpCL5JWqJMXdbSieugSgp6N398KorM5SjNJgtU11E7
j2KUIFW+v5izbfg25syeXRBM0QGLi5aJuwWFJrmDtMf9N3IJHuea3Ao9pTZl
MxycxJPxP2A26DN/DraFeo53gs35GrJV/H+jEA1WEFfvLcVVByuDRJApZh8F
Ha82YL/WTAocW1HkJfVkFk2ov9LND4C59/5xzBBEwU+MpsEGdsx21hlqgYli
JpgL1H2Q7YhwjaYvf+wiq4x1qSzbXAbAkt1c5uDSJxK709cSHGIKC0rwlTbu
1l0m7tJ5sEjmUfIxHS2l4aiT2hJgv0kj9PhWOXUo/yhGG+SIW3TgXy6HAcN5
58eSfK6J01CFCdXjjji06K8/cR85L9mZEWvCv4QaZsdq21Q/XEG66qPDbsKz
zn8GzpxUDB9jAPrJkoMeAimW31+5lhAMHhn4cMKSsLQRxwwuZ9ixc7jiSwC+
aNlWwE6DRqnu9caTtSqS+fwUcHrjiSEH9wjCWVHx0IMMPrtvSdceJD/UEDhs
4HBfDNiLK8qtx8RAscwUad3107GOsNizi8xkByigLyO7e9txCdzZNXcuRRjE
yTfOwQW0Dj3a3yZOI2LFCwl57Gm6CK8VUHPWmTWxZQjcRIfIW82EsrbytLRU
YUVQowheYLflhT9R+e8xw0wJtUikx+eaUrxxlYYe7eIdPXBWA4AOO9kQlCfJ
Pgau0R/cI6KjZSpO17U4gEoKpV67lQV2hE1UZOi70FVqflVsP22h6MEka8Pz
mMmsCAG67MhWTXfykn67V2hSYSOS3x6m4c6cezDq/GhDmZnjwLg829fnoL1B
65IW3WMjCNCGpmlzLQC+bgwF/lD414hbUpeZ/SOLwdw4D7Rqd+w6ZnwJ6lBa
5S2ltGBVPrlII/EGaVw+JfAIp8JJeZ7CcNfPknkshaRkvDAi1tarn0KAYNXZ
8WI/f9RhXcdp9OMCR2Mx3tE0IuwGn7ldGht51QNnW5gndNIOFGKSmC9f+Wz4
CAKzqvQWrfqSuAPQz+Nx+kFk1jENUgsZv9PO6fmVh1qaQearC0vZqlvULjtP
Kt8TZn19hFFRSUqSW6B696v3PTQyFKlmKdQp0wGkTSVILolo96TUCM7/MRkE
J2CesndjLYA6wodQtsgmR6sNNn4Rf8oPVby7zwHFaondTJ69nHwzI8JOC1o5
8A7xLpIK9x9cm0vQwjfhtzF0LiRhVEGgfnWU/oVjce2TeUBu0SeE9CD5A9Pt
qtz2MyloBye8hnoa6iD+DII5JpocE5NRrDgKe0z93Fo894Q/wrNgRF5VEqxT
av2kHvvflBAwRIfQknAuvRIkLziNCmDkP2eyg1XSMZQv3aJr5zI4fSscoPjh
LhYfyubyIeIgLcI659kWRaqBBi6tu7UdH79hiDjldaG6C6nbqT5ryNhjekId
2LrKu0Pz3OZMZDaoeW5GgDHuZ11uACc5nOMw0Pkp00hTuODeRIVF+onOhA3t
5lvnfc13F4g9FyUkNXWnGiKC/kKdofA5jv+6cdAHBeFrANGC5r+mZM5ROEKw
5FkXgvdWF+zlpfEpsSUmanbYkokAVJcjF7/iEf+VFSWNFaPxIYaWyHwuvb/S
z3iZVoHSqx1MePrnjOliu7mqhFBIoudQ5uxvcyXtid3WGVeujKXnQ+bBwQjt
bypvxHfUuz4iHh//YKvS6I9X3cC9njGwZZbzBERXcshzKXHrDXIePP5EHCnO
Yo5x6m2UGyW9oS2T6ZYnjrJduRj13WFmyx/NrIR3iDt2F9USZKAffK0N7ujN
9R/yUIlJHDTl60lLmXpGPQEBJfewM3xVZoQNb3lQStdE2xfFiWJ7xT6DQC05
sqS/yf6fm1KINFQMyF3DOgIVMzAAQvyPR/tTbYOw68dlDbClNcjr8kRAbaow
pi+jSGss2wh//NLPX7RWw0LgvpkyxuThMmuOKgSiytkcLV7iJGGEz9uR1jw6
ummi0HabOT60VsWLN9hToPUL2R7Vu9w+ctJb6a4Mt9OGLjRSbs0lF9H3Bex2
rSS0+SMf8sT1u05Sc0rAsDPagJZz1dIt+yHI+fIo7y5OZp2bRdARSZ140xNJ
aunfToWyGDwfSmpNoz4cHnUZwxa0rYtlrpykfGdWUfGb87Wj5D1HbF844idb
f2nsRSa8f/gOZUb2ZEmibUgeRUqMG4AVd2gmHf8dY0mXycagjWQPbkgOtR/c
/x1eOGqEs2YKHsPnYztXWz0kZ/EE3YxNdaCA34zZNj0uHrDtarbS1ibc+YyJ
ZKfUW4ScRj6PcSKQ6zy5NNZqSmzDZhHZ9udwAwaI8U6iF2DQFvgqgUZAQVY0
mFZcqH/ulbqR4Kp+QR6sBBbXyoHHH5/gurHfzOU3+bMsfBbwV9Vzm6oKWtEf
/hckijvpFFUDVzTOtAHvaEQ5C4QbKJ+yvhaVpf7BJwgqsGuG7w7cE/8NYkao
gZviuFd47EjGLiZkCULAKLs37hN5aGZ8ohMeOwN2qtLWCxsk+HeyqPJ+8UM2
b4guh9/alaE4AbTp9x+sTGOdc5zpEvijAj0oiQRhU5TZ1c+jX43K6Q3EtNWp
upBIgH1m1Rd8tCSwfK03P3nZnjkPV2Q5QrpM6eDq95Wf6Vq67M8qiGWBxHNM
XwAIDJ2/3OZ/8WUyV25RBt9O07OaMfi9XtbOdGp+ngc7eOVEi2uQ60kUaJ6L
rX/hP4zPY3IZZewcRtsO7/zpdEDJxEKR0X1i+J/F68tRGzF8Cv0syPj7Y5jP
BQynGjRxzqJYF+dH3Q5wleXoyeM63yJ7/O6rLC1PDdHwx24S8bPemYyh/s1j
7W6KC4rTNIpouPSweFbN5npF53NAdbMJzXxxBiW4JVr8pvMJvL2HucUv7Qtl
45J/ojhtPgR5p6rQuOrcunXRZzHBbHlM9yUzRlMQz+kAV65n2CilJLYVckY4
TWZVfERHv42OcS8zmWGkfOOlELRp2/uZjKiphgi3Lp61gNaBR9Sk+UaH/rG9
5hZ0IRMsUHloKu04lBO4RHKpM0+MGiiLsRXGfo8lAHhBSFPhZvPJ9DAppsij
x7m3T1ftp4vx47qEEvmj6YdMHm87ScD1wjJkoVuHkkqLs/fvMeI2LqPNnzGm
vnwo4e1fik1oXFh8LRckvbDmHiHmihXByikrgrNN3/LM7GnP6j4/pgMNiNih
jbnJIktcGBkl+Kg+dgeNOZkXx4qELRyvmLE49u/tqht8BDTHdhggJsvbSdeC
cmpZFtmTMSE7EKu8v0mJ8Er4Gs/oeX06F/0FLaCjJUlCuTKaf3kfij25A4CV
W0NZcBs1XxlRdvSge11vLFssR4sByEPtlX2kMno0Q3B87WOgvgOlvgmQxShu
Wgrv9a3qiIkt7piPBEhED75fxqQDPSgUpM0RuYo+h/r6o8anfZ5AEOHz45HA
W9TuPLjJB5TmRYeFvNW/ZBRtn5N+GdeWmahnH9JADBP6rfcRXDTGfGPnZ2br
p4CYqfppBOfn5UOG+hxfYpysE2fD1ofC1pZThg9Gzo0/C8oUnNrXqA8vC1Up
L3c40VQkpcpQdlBsRMD8z8bS4vQIEv9/0ex9WcIsedqVCwUUvvp/iwTgHmPX
JMWIIxwx3zqReAr0Xwx0Jaf1Qs35kfdd4ED2HYtg/Mo4sDG4O5v/9jGfArjq
tLnqebc+FXY/mUd6lTe8xrVkRQB9rKOxZj/WcRvlhU8NKPZLov4iwk0qxMub
Tr8fadNJq8z9RTEeXQsy5lnAuGBhYzXba+VnIZERORXmVRYqcjHx+egE28BK
zLPRHUDw8gSgOPFvNnwECXdSbyWSQ0k1+/Bf9h1tYSC6fsHIytxcWCJSLOVv
HUIAZZNTDFHpkZ91xx2F/YG+158aa0DENpR+622yahDGdAJ5Z4Lw0bpPkpNG
neRxInysRVmqCM+99sSWXY5ImkVNS+gpprT5kPgPUP+OH0D3x9BsZEnsY0tn
MeEyAIPqf7dDwQqECW0DqGyXGBFQTZ6xp6o4kHdHwHaX3/RHR0TYCDnedY2e
A5NqsHfYjhnjGxHMIARcSZD8K74PVNk82deKEPIvlDPnoDGP5E/NltsS2hoH
fXb0DEpi3cZuD7vdYP2lZNdpHORVW78+QmkFJnSZjz5oe4pckBqSE0oesvpc
CCCeeIqSV1Pt4dqB75vIGdpFfldynHvU9yh7Zc568gdlQOYKsa6q8diJELdr
Z4gURWQdloENHf07h7Se4LiLxKg0WLlg/1GrK5fh7FUt13L6QRdxJf4fJc5I
9Ra0SGwjDoXjwFGSHohcZ9vKVYa1sK8fL8OZJDRDmoI3UtLEKG9lF2kIK8X5
aK5UeOOuCiGUHrYSz91ZugpPkAPATGVDiH5NocSEd8RxYYWlNtqtQ4MyiUMH
+cLeyNBp1N4QqEP7Pdw9hQlTIGiKxPfZLJXoWqta4idj6HZYFw1hXJMLNhbW
UM1Ct8kozN6KBn2wwkZDBe1fdtsaOy7l5873AGd2hly7zY5r1cF1kRu6BkDp
T/1CHmFb04KlaPyuUaBUf4InxrJN6spDw4kwS3EHIyd+D+esAXElX6n7JFw/
mj9TDDl1nSBx+oa9pA3tJ0tRDW8h1rgAQwKQaoB9kStBPF27PgF9tKJwzIv2
F2jnQvYhOfzojr5csWCURbwTGArmjyoCAzGRH70Aj92JoEulfyUI8F9C9rJs
ZNUEfapfHFo3/Gr2ZRk69VU69n5WGpOqWjwx1LlEC/zpS5OL0cZHyC/9fyrO
+rcb27dkYu2x40jcgNty4DY2CVjD0i/TDxrWPiRkDHtdm7iuJateE4uZxUvT
m2OJzlgfWQEzpS7ipRThmWpVlYuKBKAYACCYlQ711tM9e2NDaEyp667Ma0H0
AiLwYRIPwIRL6lutz+bcE4ggDuXvzqkyRovZu49ljXYB8i3OSYTDpMUDBMex
Ko1zXiu5qRowUBbfn/eMFYARkZMmhhpV5oZXs7VtIw44i/nc7TWsfkxI4+2k
v7sTBW3koY4u3qwlwQ2fco6Zy1AKbIJZVSDk/KL+eQ2H0mtdw21cghuIzr47
v4ee51UsyRjhybcl/LWPofjBLzjjkA2vqn1RFrJfxzBfGxgFZudrorto4DV2
DvOpBxt89+iFsvEO9oWzcr9LqbegPyy3b0LC0V4vs/52fG1DcxkV9nmioXw3
lOY1SYzbhBvIPXXhUAvSoYccrQMZz2LMdIwx2k13+s41cAq+LwKfMdmKxgds
a2SQYbTTH9TlluBT6yOfslGVOg+x88hns0lUWwaOWuPzPL2WDlV75EpGLyON
hL3sPdl0fmHN9zAnmh/9uiPKigSqxwtKCaGye7SavlgA5Pk5EV4xPmfLc3Hf
179j2XH/r0/TLlnMxd+i64wcd3Ar1RpCslRbOwhySFLT9RGC9wzbupjZ12wp
JCbRi5S9hhUzigqe/iKlT98Cv5IPXdZDHe59ci26zGFqvqY0GEScsvcnY5A6
pC2FudDGNzEuspwpPuHl/gqYQwscY9m+i46iW/locQh69WqIfccK62obe3A1
8TesCotj+lb4RaFTNKnnExqeQwSPD2GDchyjGxEa5nfSOknEmkdX8B8XCgor
O40JOuAf/PB7TeyTS3zE9KzfoMf0pT4PpT9A4Igg3SmbeKPjsruVUbzLdarN
NajvkgYKbJOTaHgwrKFz4RMu64sgeq31N+T10GRj9V47OyC+hanQsluBJUV9
uDQ2Wf78YNyoQh4vbLWff7hb6OqOMMGMQlGd/ecfSC8e/rBLJfzWWRb/LAbt
Bc2VnZS9QJJSB+pyk3n5ZYsExjxd9sChdHaFy6h8xPMFyJ3JdTFfYQs3C5hX
7FQFgjLIPE8ABavLk2OR+C1HACCXXBxhthjt16HBsULEWBgLaAmAt82EP1ew
rbdk0NJK4D3lx/FfeBx39vyHDFoEc9uN3Yag2z12+Y/sMn3kJcCqTMmd+v3q
zAKYav2fcSQXQqJWs1Zuzh6//wTseCISr1vv5cSOVhLIVWphFEgVUhhfL3b8
+pD505NRqYsU1BcxJOPiR1JT/xRmzvTJgyWGTemcXovRrIxA6fN+bIPc7mbF
KO3bKpcHgkVOES5ZDtccq6+dpvqLhhk97D9m7rKTyXZ2dRQRnMUzOGG1WFQk
/lbWWtYQX1xc+HG7B5PvKMxFVTUTWIUf68evOaZ/ig6lfJ/hCjlU2QeeG5MS
nkn/Pm2TL+sqx6SQ7U+OZUcYupXEiCWraqIIiqwKvXYS0drsF6FnROy4JVQl
EYIG5VVZMTyTHc9VBKe3LKioXyXDzmj8L1ZahzuvAbPg8hD4x6pj7dWQvC4R
UQZGDneWqt6TExnBINfJlc1Y5tWg6NCJdM5xQzinNBOZovsg1ejnBz3ip0Wt
JlRw+YYEbQhhTWUeJSHxIKZUQEQeMeGUC05Zzt74iWg8kf2DEJmVp2vvkqWa
u0YsbciuWZk5WIsQtXKauj/Oll8RBsLjyEloE+zo9fUs9j+a9DKUaEcIrFey
itIJivFdNCPdgb+J8cziMhjT0KQMngKNi4TZB7AzpTCGewCZTGmb3yzl90X0
xYhe98pFOq4k45S72rtJ0pnt8PnJWWm84YXcX2QB+6ByIwgUoiQLLTnYBgd8
o4kq7sQfjCzvGb0nv1ljvRIh9qBBKs6bPIm8q51cVssnlBOXafOoK/4IFVBZ
O63pLae3Z2f9gOa/ysdZ0ZUvS0PSvU165ToXymZfR/NRNIW7tTU71j+Nyc6e
NPCAv+9OCEKBlbK79cdgxpIFIhjuf2ddQo/aQDEAalSVzDtvaeu+UdRCGMkY
4GXToG4PJ7PnYZPEzNEhuB+kg9mfWJDzu65XnJkz5ryC6r1fgq3+pZ3fbuaK
wZvcHxd6zTu8fDaINsPksAI/h7ZrVxvuH7837gYgqjffFJ6kH3IZq2mHqLXE
hYXL8dl+KIbZeJeF6rnPfC5byq5NDgI9pS1LY2flQlOHJJbLTiELp/T0Vch1
jc5JMuSuVJOAjb9olV0KNngQ42DrtB82pg/PMZQ8+wYkzX232yORrurkL7Bh
pxLVA155A9U4vvKLyCApX8G4Fn5sD7C+7DmHcg8aIx38oiIKS+0gWBtZ2qFe
/aLEBFcB54NjTdsewMt5w29wxEmn47QcylZsfaS+xyg4WAnrbCbl+LIkaAUz
CdS7eARCDTaViEx505FAeMWTGsrk2xBgihPyirj851B3XPs8JagOtCIh0GDL
kl4lq1gZdUoC4wQmPkLN8OwAslBNfTSagzgGNx8Uj5d7CnT9FVB6KHFJ3ftL
/hSTX8hl1kCOota3sJg8NxbBC7NiColonOqjQ4h9admgaQTEEyWi3RltMymO
+V7pH+7Cnj5972vGc/yxLvw0Uo9jsF+gZdcc9ZYmpwMFWR8qYssT51aq7Bpl
h31bP+N2ta3ycSJ6jAm5v+kScqt3nRNJfupsRIpr8f0usGpFsPWT4XxO3ECJ
QNuaOArIpkvlC7vGZCIDsJH7cNEoqrtA6+bi7QbNxjR+C8kyKReAIL72Dw7P
B7yxIbD/HJ5idF+DlTm1zuy737njwHgRJPh3b6svQ5Dico+56HpSHS2Q9DGH
Ce4BpVGs0k0/79skLMUtDrHGHdjNvsFsVA8VwmSsoL3vACXXVYRbsXIn/CuR
w+DqQKA/nvmIc1lMAZzPChn500noVFqAnOlwrQVULU8fP0AWPQo41Y0IviRF
tme/gEIZHmiD0DPPFS1iwOxj1jJR+r6fVodBSDH73s2NZl4hN+ip+BmZYoOf
qRElGH4h3aMIGg7/pcQFM0fAJh98PvYnv5UESg+B4kjR4E8JQppb88ZCdruJ
R7us1+qUUGHlCB00W9dfiI4IHVDwRwD2ybC6xtldFPWl07r7t3MEubICc731
GdySRdjeIhM5hKUGX3eugp70QKZs8yMCJHFldSlbxawWa/1zK4B0Ss5nl/8/
XRXulqCSJ0mDkDoYAKo1vyW6cQ4i8VS4O8CkJMwQgykMuZJRF3WIM2o1B4Ja
ocSRXo3F5of22KPAe9f5xeen3Lfyn7m/+64ErVnAMp1Low84Xov6DUkcDVws
hzGaFSNzYBpnDfwEWshPTt1TEMIm5DWpoff3r5Gf32lNo9EG69WXEAKBvwI4
wXyt71yOWXoP+F5mXstyZjBTnHZmDG04j+xmqkuUHy/WC9K6h4j6faaE64q4
Yq54EI9LB6YG9KqAngiEUOoeH1t7OP0qkttdCnOs7H9mGJRABAxfZRI2WrFx
mo7IkYRQdShCQAvTDpeYSnM6HNaiCo+PMs44J4iQ2f6C7nxGP5T+t+dUlOT2
HIJmGp6fJKhJUEk0loRd+zqZ40hM1gvdBOrB4xnoI9O26Ga96l0WT6srF3J4
rgHlfahK7n59ZnYOMD4O2/jYmxds77UaYz6oLr8twtBCEooIunUl+1Eph9YE
5C6rEku4S8Wm3tkOTI1a2UTeexDfG5NIa3GgDwm/M8Lr9ZG0xqggmDHAxMwK
VMC+Hv7WoyzjlXHgs/TUoz/gISYAKRWhNG3HH+zYDa4/29d109/KsV9FPwpc
d3FO/P+N19gZhEus3DtYubRUGKChHmnM7oqvpk9My3xnBpgoQchdU0Yztk/5
wOSYo366UrjIYSimJjnioeXKAms/NF57zfVcz6IiMFnYjJqtrb68q9T3/ghT
uiVYfXjyOG0zl/k8M9M6aR9wBk1yWMJnsRU/cRbdfClaFWMNxVrA9OKypawf
npWdF+uPKX/LbrWdWvrUExuEpUFM49tzclIC8UjpyvXN+/0YHcVAxkfTVvPa
0lJSu0ZMhx0bsMAjF1Y39jiqV80Kek5vxukaL0/cDt1sHl3MvzfpzaTgAeLn
uXtNEDk5kQTeqWKhJ+0MuxMe9XGQLgX005REGPWyxHBP83iAXu+407/4dZjP
qGy/Ul0V+hpkG5uVpqRf4pOaZUXtFb0iOG/6RMlkWz+toHSjlb5vhQnBp0uC
gYXirhyOoMNMz5AU2rHXivXzS3dYH0DJo1ikVZh4OOmyU4YFDbVyoRzTctCO
XHJA9sbtVePo/9bPq9sv/WoNK349nWoAr2NUkNuV36TgzmyMsSzmUmFqjiA2
juV2M53GaKbqDIDbbialgIdj5GC1rSVBMQNC/cAs14shL5dYnpzdj6XHolA1
vd30Q4kj2/HUuz0Tdby7Oarupmp0TO/9tXf2UAFj6TZpAi8P7qip1qKGf4fE
82DC1J4xtfhEwx89NnAZTmv+RAlT5+uBJceV1q4cPheCmMa9cRT8MMUaNhwk
XlzvVjsQ2z4nbnJiX4KVxU6JEpijDLYtAu1rlJWHOXj+1owCZybDNrPoFLoo
ngWxTp8SoDb+Y0bQ+/9h0bdWS716R9d5o70dxsjmZeq86zWtowzfU0nEYuOv
5T97KhRpz8VhLWOGLFRximwnOn2ooz8BCE/gF+UrSNa5oq+ZSODtr5BEWSe5
uezuXAvzGAp5WJgs9YMAJ+KbkuqiYSiEdKcM3UsP/8uUoshUde/puGLHMJ6h
/YA7eptLxW4g3rztKSxGiq1wqsw4mMCnhDHB1wsHxzDKZfxN4G5P+REHqRq3
dK2DFY3txup5TrLXjyPS3hBdoUGgG4XnSK7v+0dxy8/67bYP7jlihwPvMmLn
tmxFrWWOF90rwToOtgDU0Z97obtygklxcrfbExcCOjSs6lH/HxfmeVgEEaOp
pbyyIj3lnk9CQj+WG+mRb0ZCnyATCLBvOC/TL4GMjvnxCQ9ikQwr625sqwLm
Ee2DDUEMPQlxa13ydVUg/m300U97h9UXE2a1NZfIu+DO9VNprJtC2p9uZwMt
nF/cBsZq7e2tN3RrA7tpOnCcNOChJ7TnnwXGSZtYb++Go6fB3pqOfs4LmqgD
5nAdaYzqfYwTVywXGcF26xByOy/iAnVB9gTQW77utIRWR7ggs+Gk/9V81bYF
D9KrmzCpf7gsEvj5460WoM3jD61u/ekDzCS06Re4TzwULJyGVefwVi2wySyF
SrglRMBfJVDQCdbN5n2CUKlReqMltUPJ4futIeyWXRlMhLz5Pl+xD3Pu/m+t
kNLUYyJQvAgdAwx9Ak767Pv5Rfcv0RlIuDlkOeXU+loY6K4ZQaTx1IK5C26S
drMothf/SS7wbkas569+H4oVFNUXN/VZE4RHeq1venbpOvUaJsdY2TScvjbP
ZbX4xM6jKU/xowRnv7QZCRMSplj9CiLIJsxl2A3P6B/xGPF3dqsHgwvEqaql
gia1c2Lj0xufCcNHk40v76vWFwtMAqjWK1JQ+R1PwR3usKvuW5I3AauW2WLC
/8Hobr3QzSKyna4Yz5FdHbnaFrgquRc73mOrfDxrHJN6T0RRTvzyAbtwJgvU
EU7Ain/Nwu+ViAHaYNOuX1WIYnQS5bdh9GLEPMprrxz1ksIeOWU3q2LdRbdF
7H8M+oTQAkjhM9kt8QTVNSQjPSFK5QQNo3n/qir6qqeL1Hi/MHxXjl8/Zbgt
cgxo/Q2ZR+bBt5lkO1wP/fSssT5mkZFlaBNDOfZqwW/qPj6XOHocnIJ213KI
eGHhezvVJWcaU94lOZHw03fcBJpnqk59dRT4y6LN61H3JOaEmOgIAnovxWC4
H5aqO+KBAy4GyJjvHZpih504hZjDcB+krNwJ+vDbGQltGfJBB115iKl4bQ2p
j8F9pQPdxXN4ilDH1gHmcSvm027cwXLHAXDfVCuI/k6Jxt704tc0IaHiDM4a
cdz5D3rz4OsEftWu+5p8y628K7ATt4Lwk220X2VKKXL4yP+8iGWWobCjT+24
3WH+9+8DNMm8gq0t/FHaDxj3WCRNHQNBJO5RW6moqDi1j5+snE6vqBtk+Zii
fhn/vVkIk5GUsysIj2rW/RyFLI3EONGssZ+6glX75Y340s0VjBrOF2SXhQbt
zeoTcVneFMXFawoZkK6GHhNCX+nNwGITGAnI/8mK3D+P2KE2MA/ngBft6xYe
nmxeAzFKJLfYvQmIoUw/TjSJfkxPiFZ44X5KM4U0eUQteSfyQfIVlG6vGsCS
uSovQd7Jm+fxPZ2S+UGdDivJJsi9LEtopHJnm0icRWW4Qp8YcgWNKt8N7O0v
Hs8epXt2yVz+Fa2HDQ2ZcaOZFmK2nG1meZCE5pW+r/GMSm/GnMl95j250C1l
FyRAAHMHbgdSqfZ6nDSyS+4bjdT1vsSuOj/RaRH7qT4AMBRmX13Z9sW/9Goq
zV65zJa65O6miDI4JUbSWrnWYEZ0dILbzLEHVcIViMT/R0kqm9qnzQFUkJor
T2KZY5UN8gECRUIXAm+RhAcUt9Bk2bZIR1yYDSTcoIRs7rPKpkKVuoU3j0yj
Jo25VW12jSbarRnlPv81CMYEKiGRrLR9p825sgqbIXKKbenFl/Y0cn7FdyZr
DNBb3mS0JB3K1tFAY57O/ZHmDIn8xSDyqCU8IVbxrF9haM6xvFVoVIdsHr6y
QnQlwLCBFMAYmar1MsuvJwWLN0O0qr4VvnP+IQPORwm35sgLPUUYU8Nxq7cg
ftKSt7eSWW51zRm+gwnXxYaxIBNOW0Yv8V64sW4mZL7B6wIPEcP8gJJrD3/9
qdzWo8ZJY9opcgt/PO03izGM36HhKj6PHPg11pOmPQYaFfAupkNPrmBvM+8y
yBUOhknwFo846Zi1W1hNNVpiyEQOPKSD9lpi90OhvuTGnaaPtrTJbSgr29jM
lLRL96cC9+COoFIqlIl4aY+mV0GTsW1KTZLJX1QcCksw2hixd+tMLb8myGJL
zbkKil03zwFGFQbCazxbeQJrPwFq7lKPm+47+WULhDJATDVCGDnIzGzpNikd
g5Ytl5uLiDBS8WjLluQm89iNBbUVPHBpdcURob07GZehDAVPaUx2nA8dri2L
znNQRA/LgtAHE6x+44yrIueVNLn7VvjuyFs1lgTzLYIzYqsT81h+hQRuIAKh
jKimJv+J/4LDQRqOlhwLi/QVYZ2Hy5FKh+Yn5I4XWppdqIL1/+jWZHEJ6UHV
ZHGNSlgFCVaWdPHvnuZnCGYThqbUCP5x8J20okbTQXw6fRLQLU8SPuAqc6gz
ZINFOjtVPyyudPVZ/DdpdIUbEvHy7qXKauEyuyf+KSf0T7IwWJX+KMjJ6h/p
EKQrUvzDJ0A8I4mFZ/BajnvYvGOgWZVcWUAvGizn1y3P6NA/7pfsYgNpJvOX
gOA6Nlnsos+hHsF3/xNGMTj8N2AIw7lfy5K7HE1YdWJoSQnTYHof5cgsJuQd
FVDobHBnxeCS8Dt8LVuQAT+HYtu4aX77ahgyiDzgD3k3seVfINFwS8tTS/gc
J2iGStPUpbcOiy9qlY32+TEg0mIWMq8lFN5zMYzZeSgi8mFSW4idbyAIji1x
Vn8izgt27Kel/cEKBMPKYuUNOtarIvytuhmFGo2noJjTgn2jV/lCl0K+LpEM
P001GEfMBH2l1BFJyHOFEAB9oJfWbjN9DbzIGpw1x3tYV0nsuMCk80v/AZBa
DW+Ehasn/r0uB9RwfqHFTne57Z9r882DLMSJ0xsoBXyfDjUu9MVgEhlRnUO5
ybLKdZ8UxrGpxUWCkaofsbR6Sxs4rK2HDJkt0wFva+k5n1LlkKtdHm+J3qzy
i0Mb50yfBY60dus/MX7VN+1/3YNC4FskPrUkeYOcHf7PbpDBvbC575Q6rree
XcHEPiacmFFYKGeD7WtfQjqS5Qpmj2ElVECe+KxPkD81dpm9xAfOc2m5K5Y9
y/N/ocBqClYzF1wnaSMRtixyXLD8XQ2lw79cpFmp4BEAtR5JL/hSRQStaFzZ
j2zkRAArUB3hsFTJVJgr1fdB1dHDaW8TwFkqFCkisSJ5KHkFw4Z/5j4ox2/x
wdNaw3Uj7b927gJsy4VDNcKLpfcMd8OIgyPFTH1cY6fud2hY4s4hpxtglBjI
Gn9+7Zehjvz6ahuh2cqQ1T/7/QO9HUveY2mHYnE3XeOnzThGWBac5hzgkv9K
43RqvUrA/hABAvDtQ1gLhz0mYqf7/ex+1CCAofudWu53NyYI1njpFUjYZS5H
R57/Ibb8WEpyfVYR8WsWh20VwnTSqxST0qLAwDClOV9/UF4n1ZAcvaQvKDWv
6I9k7Gj/kEuAjYd4lRxkG1Emqq6MuS3InPa8srmjFSzLp7d2NCQL9bX7tCi/
/5msyV1iGQid5cKJRLkl0vMr62vLhVXJgHzY9Rk0d0iNrRX4n9ddbHVcRmMC
PJSa1Urru0n+8p4IHHctojgJu/MSLTOBVQ8SHNdfZNhRV02YBz9ZpjRifBdI
P3+c+OUmhHRpMjC6IR8mP4gPEhcmXjFds7gwUEWIxYcGTkoa288vRADwrtHX
fyq16bR3HXhkCCu1CLaALp6e//ied5QMq+UpNCH20mxtXBE6LklYcaDNNUzJ
w17x5Zf7nejEGzxKknVTsWMMYdpc/lfuT4V23mVCVXxeukZLwXytOFI1TUqn
4/DYVUt9uuNfyStEap2y4B1BL5zjUz1he1FFNR+7yPrNA834ILPVRaRIq5oR
4DMrwW3xyQflbGaXRaPh60oKPr/8uUc6vrTai4LG8YJ3B5YUApHwdyJBhn4v
2d9rGPCXOGoiZ2Ra2/wRWimxjNMAnG9yxgfJB2/rBHh7ltRUogKniMJkfd9w
wtai3aG4LKBUkzN5WNfhWSdA7dafAylkEeOI/sS3YGhW5QDwC9siOSD/Zu6Z
/4uu4yrergtz85TQ1JMZgJ8VA6x/deo+hFAkavHcwQebPzX33sZGLVUgm0Si
zIERQxrq7l3ONqbM7yDn+dNFiknxUgHh6Qu5rIB7ehfXaws9W0fAAxAcO4G9
IxQz+v2ldW7rEZkiZnZkHSIoZQGhd9gqjjGGzbwNL3QHBw5Xf9ES31QaHTkb
MyAbDMyLIiRcN+Krn4I0d7kgsHaIFQ6EQicKGOh9iFsRKFW9gXUWQa7neW7l
xNq0NKg4Gv6TTOl1/ob2S51YbNye41oafD0lh0IsGUz2Ava1cUNO3cpIALCt
3HGHhmetmrVHnO1t9sgTvZUQQDidD+tRzQgRJWL4sqrCT+zIAkXVUQbhQLEG
q0GS/Sab2FfHW2XOdKXJ8tbnzHzg2QiqpVfqJygfUmCBBp+5oJEtSe+QialC
XRNxS6Vd/Oz2KeR5lOVk3Y13zRNYbunun6Kp8lh7u89P6VpkEDRd27/Yt57d
KQOa+8CismjPMF1ajUfxd/EKbJZH3vXxGeDVniqxSLzmibcAZ0+bUj5IIf46
BfN5IJ7NamLF9GVMhVoBLg5IwSkW8DaoNv+NPd+jS0cuqgo95Zb+1TmnPmRr
YTNXyHvv15a2rxzpgPYBoKSR+/dleNDiafI955tu1jkPOGYQaTASLw63fRp9
StqB98g4G0S4+bkmXzEkSgu8sbBZ5DDxKNqLt8AvetiloFGgZKPOfCyWcAOI
PmEZIyep+8CJdtzjmUxVCuGzMQvj8HltKC7+1c9Tk2YZSXyQnG4elnFW5tIs
lRvVeB6sZ6/ayjud3DNqwYGCMCricFOjhAfOhIf7VVk43TUOzzEX4b73esaz
J5pR2JlMcKExEgmIOqfWrrMeL3vLLOkn6cTP1m7RhSp+n4IikYFFA+hohKAb
o5Xstdpp3VyVRdNAh7wIm2Uo//HGCRp4yzs1vstrJcUzjiNV1s6+lAdaq86r
aXswmtyrR7oiMAR0WPe3GyUvoHyJ6VdMUUwnH6NDY+ryp94enE92GKjS8VQh
VYlqE71oMRp2Z82rXiCs/Gn762ymgl4YOseo+TN9JuvjXzE2djIzgTkxaJVJ
dN/YF8BmKsoX5V54ZvRwQE/QiRlk/J3Oasr5tLSepot3yqM2KpemIHApiiOq
2RpJQkQEqAq9dX/rWvE3cydwwCyJqqpuPqr2yXIS84NEs/jWaGgAYSg0529M
BDIBKNhLRp8f0Ylhm7Y+HSs5Kbggv0MSB0T2ygQKvbT6iMwT/P4ipORviVI0
XPbHEY555TfgN4d09e0Kn1VKCuYzSOiLAVAvSEOGFp/os/x4eJPtGxX7SKPj
4S95SNt+oQsZdYpbF8UlE+0BWxAbOa5X1EZcxyYOnVAuxK+whYJFbsSyk/WK
03rHyh4AycYQfLh1QO0PrlsiTCsylYiuOq/ndrckt1iBzQWPMVA9iW073Cq/
ksz7UypUt5XvDCEi+mohKBheK19DNlSaoPdFTsFTmr4SIrs2XwBPRsW2pPDC
BBCawR3T8/Yp8IYzZZ+vHLamun6dLchEst9bFO72eb98vdWBAHb4PBA4Wfeo
guJUElU9AoN5gxx5w2kjBy43w1LFJfGNVanAQi+Rfd/x3fSpJNB8ZsXQyg39
VD8OrRbM2sQIr2yq7nb9Ux84ow8hSBqndRtws4df4xVQjIflzFYBhPl0vhTI
5OaXS7+Bl5zbRkb8sJzTfMP5JFANRvETLd3ZBl+ErmbfkyvHC9XoBHnrsiI8
83ri8491Ku1ulmsnwC3rgdNdKWB5Z6+WD99bESBvkC3EUdT7bTtMzMnpRVcC
6+jpI5mXFg1QdDPIhyb1/9+6iceUk8AJAV06mbviCkXrApm3Bu6DQP2SwtSd
yhyuR0oQ6DPo5QfedgP6eSChTzX4Ug4peNQPwP3a18TagAPnu72GSi7XXCcX
S1q1zbvXoGOxHAyGutaUTagoXC/0pVMlb/O9+U8cfT3ICQy+xTpTF7aAKG/4
NDgz9yfKWzn0LW+n4o6uv0XbbhiotJcxkaUOnHpb8WAiQPNEUMVXstnmEE6y
ah7Sp+tvXzdW8/Vjy57eIHjcVRT2brQC2eNcGf8pNVkvnQoDalheXJwPshzU
sS48Yvra8GrjotsVp40ho8WCW9V002i5A9vTZokh1RtRCf+gTGLq7ZAOckVZ
YB+Sfn3p+msebR0/kxWxdzgKfYvIheoX9yhhU+hw/TCI+FAvtpNxKS5v9ZJQ
cliuREmBEcoxSB4v9FyuFnMt4s0FDTLhttgqDnnZapMwkJ8cnhzznRIVL1ia
s1108ZOiHuCZ/YkEVJXNkPuJj5lTTOG8NiebZFZYmi0803+C7glZqeFVW16Z
yIDkk8F01mz4FBbnzN/Tfyd56+eNBh7I3shkfwqNC9r8g4jJA8gP7AnEj/yQ
B6AAO152BG3Q2EF+TXJ0vTvzGytv62EvnfoHTgUkOrrl0bEgJ6AIhjl83ZOt
QgCJMJ4BPxg6goRY+ytOaU+racgYM+TFZZhnyl88rVtksFpF44yf8wtL7FJ8
HC6FM1gqaMwZrsJp/9o6McUPJ2yhRQq4zlVj3EpChMgz4Mo9J3GPgZZyJAsh
BSJASB0aPPoaSOb1Yl1tkldWqulld7tsMVClvQJqaSYF+PMDZYRGHAVvfJ3k
yVdinKpVpgKc+XIyaRgu9cbtQG5v+hnKXpO+mgoysRCYXhz/IIY0oDjZHXcF
/8TXi8c2sdMPeQCJpo6d13zQ1j8zMzov++z9Z6/I/9cfUMxKVCm/qpvP3FG3
78H/lEopmk9H02hr/6B3ErWL+02Q876MU0LPwalX+GwupEMeyhzerXqCTVnp
wYgVpkJbQz/ELchCdFXuc2r0VnuFEC0zy1Y7sacbv9c649M+hHRk1Ft0NMG6
ipRsACczYv74QBBidwCwM8g9jyBewrjf1+7fxfY2f6fQ2ZlQspt9NVgEOoI6
v2Kn3wd0sk5IKVOlzsOBerTk88BduGGkU9q4rEW+X6xR5FCRDRBD38YjIsiJ
Eh1boAqd/n02ZvZYf9+90NIXhj63lHrhfbc7YsfYOHG6HvRZ0yqiMiQ5U2KA
rFUZHGBkPZjrMwjGDqW7mPmHXqMpCUr9Jxd6PAj9GhLTZUP7RJOkB9ukzp/E
a1n4LO90jyYxBvr6sfaDUzs+zjcn1Hd2m1xjGOEwknj7Uaz6uBYi2/nvPbVb
hTbUZU+nCzeqsKm+ECje9H0kcdTLHHUSpiYHHKx/PP8O9CDdE50KwHK6m8vx
hzYgE+V7PpPpWzxkDtwThFpDKhtgE/c0laqDWSY2cO8FWbZ8s0lPVo5JBZEk
unCWL8u9h5jfeXIiZa5F/oycXweAFvmXGsH/W3zfcddZtXd8uVcQxY47e67u
1znrUeFH9agArL3RIop+GJ+pLGq9/NtM3cmVzv8J7A58cm1Zov54BbMlgGB8
pLNBezqYHcZvX6xrvaNa05ZTCf4U9J233/9noN0/qGvdLDtywannlqUSGH7k
oAXxoYvXRzp7kz38SdfAawXZ1RWBAGNPzUN/JAD6XR4fDgK3p8pbaDX/3sCO
NoJgqYm5BOVRpmcsHEynG4Wod0J/qqWkHYyHDcV3Hq/Bxkm/fFB8qJX1NPgq
c3R07HSePyCiVepMnWu24EWf36/85OaCyP8GoGRVnxIdJgfIXs9pSp6CDI77
Qd9pjcLIXe7x6RZfTW4PF7ydN93y4ojPQiB+RW3duhnoV+6LSpil8RksZXVQ
Q1W4gakfGGgUc2HyIDnG8qnaiN+mKhgRfr17hTlqs4J9sSErY+SSIvuCwOMW
7YxTBZvb9ey4VHKCwKmqcUE3uU4186owe48mGKkjbup6x8ibviU7yFzzXXH5
IyabIcLWN+UBUTgpbdoLjGZKELNmFfySGxUStE9cwOxjhyc7urJc1WdEMTjB
/Ly1mYa4NhFNbADOxQN/D39CgLFpTt31e4mR3x2aD8AsPzFDyemPC2Nl8EMB
y/Ex+mlnVnmzSpMk/FX+PQS6NNoX7yOn3sVcuCz4JTauwh2Zk1lZEtbXDnH5
o0x+kukVts2dfSwUGG83Xi8uiYmDIhXeJ5nJPn+olR8EuDiQ9DkalzUWJyGF
If/h4l2JyEfuwf6rcVhrempJHCllr8huNNBm2/EaqVt6LkkbuXoWKCCr8G17
+buA+jrp4SW67oMhiLM4sJ16XQlsKonc5IcDljZv1VLnVHy1PTG5yYJ0i4jQ
ppE5/CYuM74Z2WbSfXmCtU9pHaiFYSGcGtJRv42bDxchxCwF8TKNnWl9wRsz
8gju7ohY9K68/PF9b4el6tFsJtpyLP6AEdEi91Ky0X9SeHABDjI4YYru20Fp
7UidKxf8Hu4bU3z0LogGVzregW5J9E2lkGWOQAmaorPRMxG68gFgh6yLf9BJ
WRm4aOnXlsd2PnvwQDpjrdf6EglpztE7WJh3uzk2Hf+tcLGWyFaqMXp8h2rw
zIim9ORk9p5JCakdnWx0fUuyr1lcAuetZ27x7S1sYAZpfYED3VeMZ6qzeGzp
agLOPEeV2gJWB6EpZikEMV3RYvNqdqUMmldn95jZcNsazems6p1kTdtD7Lw/
hc/RgK1txWj9krRT7ErZFe/vZhnnOcUVq6DBw19BjCEdm9fB2+Ch5XBVa8X0
/PRo2SlAI6NfU67VMFXcoy7rncg1rz52gHpD6FLpx/tEDY1lBpZ7eSJIY90P
RZPweoNbNQqddQWhURW1WuziZOnvqWhx/2REOCrSRQdJ5uZ5GXkyToxyPzXt
hwm0NDTvXsMKOiGunVR+CNnK7hq++110s5X6U9X7pwCF8i2Qg9CGaFnnFaG0
Zc/How8nNVGfnxO+XKUYMAhc4N6lpkAQMROBkJNJWBnVmFIDDoqR2k6k+wOo
BG4fGSUUYOtIi1hefaSdtrqxBF5FFvlpQTfnH39FdResFsfNxM/cto6pjKQl
d451Nw+jp87EV+lZU9NVH4y1MY8EKaIvZSIR6yYjMn357pPGODYMvvrFMXO3
6KAOg6s2gRhauit7vH9W62EEJ5kosEHWW2dW6cL0WrT/1GYgcRv3lpug/PWK
K2xEq+PeDahvHx+Xl9Ot0V3hhGey9NzXYz8SndfdWjUnA7oTyvfA9kLNdzfD
N/YM4Yp0iJnvJwd+gvDBm6V2LzZuKI95F74eNrMJ3fa5UAAhH8raqJ1rSitZ
r6a//iKpdN5nugqrjF1QyzlkcvEZRJlcbeIHo7iu3sJ5375h0N6x12oQI8Id
kSToRMYOdmlCp8NnBYam7PDznqUJXoH9s+E1bLcfd7TKuPz5RnfQ3IW5Dr68
bYRlhNQyfMTvBt6jnbfWYBwe2TwbTBcF3AQARKCVI9qzMu0ZJqSqdFqC3PJ2
tLj1C4vjrA+OEEmyK/r+lw+QTAZ8jklAcB1TFJwxMr9vH6SkT2gRUvVCydmn
/7YxQ+jB8p7Lixkvls0OE+DnlTkZGC3BBBPOZAsGBywkjMX+KYYGbuWrdPX2
gFodIpuB7/VnDMO1h/SqugBV2YdOOxtUeq+cSCVntrdHydD6rMsYtXODN/NB
Yb4cQHWLsBRpT/z4c6fotqJUKZMqeH4mHcRY++4CDUfJkiJY2svBzUcbFmId
39K1KrNBFnn5hLpMT3djqOlqQWAbq8zJHOVFDeHmIkEIqwRoNkY3jdDqHAyr
YZHp8vqr6n6sow7kxBi/a/B+BTxdtTFZZ0l52Q9Pt8oVNzE0GEigCiHnlYJg
bLhrP3uXlwV4+5tZGBqnol6NS+h7TAkdg35KV2J/PhNRJQmkb38/mzLTz8Xo
FHx7ZB8Bjxz9rIjVNkwPxEtWn6LlEmh1lATSkKYYyNqM9mK46gML0VFqwzmF
GAibNS8N9gEqBCeYuFbVSiCR9+S+KPUQ0uPrc0+C+oyN/V/C0SOOI9qapwy8
19pbM+sNWYTSLMycB/CKSAPmM+cSZnzSUPaOu+j5EfDE/Hic+SEk61rBw5oB
ep1M5JnMQMWeZaFwEt8AwZp0JsqfqpmUlXpMprX9/Tmkt01jKnuUrnYEzX5t
vKaJjCgYBSsmgAX+KQcq54w/1TPWgz9eFqx4lXd3wvH08uuKADHKe+Rq9Vd+
HPFjIxPc5yg1oH79P6TG5ph89vWDeFnClNYbyuqhgBWNjviGaJf7gOjb1UOF
nxOcV3Q6qRGyI0xQCsBvgehf4tUH986A72C8amQtPi99pWOg3HsUg4d6jVJl
H0mdOoTq6WdTR6xVo5fJB5QEzvVta6u2IW5SWlWAHib29bTSLUSTbO9HfnYZ
IKneBzzPt4nf3As3Le6Q/e1UoDgJnfn3fJRPY308eHMOOfyX2PtLipLLeer3
aBOFGCZA+M87yvpiiRF2kbuS13T4OunqLABw1ENid6aj9jkZuTrPr+8BR3wN
E/mpDe9GoNLZ9CnnErP25kwCzj+6/7hk4OwAeBM6/flXWK9kewkGfJ6gsLdm
VF1FgCm6qmFiTccCQCGdk3nkaT5ERCjpcENgx9RG/8scEsdoVkIO1rxHEDB3
wo+Y2IA2VK4bh2qlXWHSC2lc8xlV1eIAq2jsdyKiG96cPGWxOOP7YyUXQJ1t
lntDny3yHM+LU2KIVfP7bZJtoX0/2DxkeaD6DfV5uF8N6AUYQdRjzwcrx0Ok
bnDsoxPAqdPAM9ahvNtklIPmCTJx0dw/cvMX1uOJaLHAUb5GFYF2rYND96cj
yU6jQAGUMrihYu+9PO0IefZGI4/EQNCZ02NrZO0AsfJmKvPUk19sYODg6Q1m
4eFFNyokXgDyEppgbhyhdRdIp4ABRN0fLNfavufexWfyDvasDSQYWdJWI8Zv
8UQGyC35KPIGMc8/eSFZUs8lGY9oOiAqNkgrdXZZJC+AcvG4YRQqirFMqFE1
o9PQulU+y5FSTtqLKxtbkw+HFSnwctwfv7ipPYp1cNBW3GJuf2cI360Dj66Q
a2KwTp7aUFB5smEfica7gwohYXGB0f+H1hyAbsMMu+P39KfKBbY1By81MwoR
0/77aaCfxZ0+sRynVt2mWIWUsnyrd4NarjwVimvHv27srtg2t4BfIn24zqES
BszFAcBU1USorg2+1e9WEEb+bO0uNGSiA21qZv3JxxIFG/ugYPRA1WPmdyN/
XI2iQIbjh0PW5b5npbaYgV0a7RqTgLcmrtIraD6oon0ZWr/qrtPr1cKWnD2y
pagueAiBJZTfH1pQ/8JBa4ZYGGyxlpUGyNoAgtblIn7Gq9SaotZLvH3WzdUu
w3tCzcqDaAo17Tl/GdZiO+a9IgyEBxgR9K3200ZJCcTpbS3Y570CeGOQoBBH
VtKeYsODldyOt15Bh9FFd7uBRG79vOPfiK8dGOfvW4toe7uXUBlBeHo8803s
WC+z554DTZN3jS2XGLf+gmoajm+9YVZhL2r4JPAuMOm3OXyHedF42jKRO8Cl
dgCgsbQ5VG6m+Hb6wi3R4bHvSlPxMRVT9mXXvkFZkqLz7/R3S50IqKqM7fHR
DMylirrmeJj9+Y3TwB7irVWjpcPBdSH43RzYkZVKiEcZ9eCUKghj9f5Ko2aP
8GR1lI/B0MfRzp0SUZIhWVSjIo94wPiL5HfH2XoZYOwtJLD5rsyXWNGb7zl2
ICS9M7qiAGgLAK61ZRARAedU57r0Ih5qYhuKJ7EKIrUyYWu+F8yw9Opgg+9G
yvsYDel/UVkgG2Q7/I7f1gHfxvrrW81J0uEW+TS33abVIQg2gltwpzgkmRYn
UtYohuZV4KBIIJJtZoIVw8jVlowzH+Iqb2fKm6OBDDEQywsxyZT5Mt0u37Re
6OJKmVWdioU0L0JOTVY3+ajZyAVb829XOaJXx3JqFD7rQPG7fQWj2o2/SToh
gwn/sf1FOxFV6NH0CMp0EU6V9SiTYg7l8fBVIpgZH6l7DkTFyipnkz3JKzkn
MjdCB7Z4xbn6qyoSVrfIokC18S61Z9k9Tv51FPuS1xhcBD45YgJzD1XeVoc/
TajZvLHUIWNjzek2bI3LWjo6joKUKECyFx+83kFh+7TjrpDMXbnRkDsgjjcq
sPj+O4i5yh2Zryw0eK3oCdNd1Ca2yDBJ9iW/hW56yt495Ng7KW2viZluuiDd
9RygdcNkJbHC6Qg+hXD5Yrw8mJo60uXUmG9PwJ74OtR7S7yN94lgeFiKf+ad
oM3YVxRArKo2LyChndCBPw/cPo5RSHOJK9mFiTalt26xUxeazjKlxFAw4YfE
mTGq9NpO5g20Ry7vj4fCQn72YLAiaPsvFX6XhSbgbuNAyaF/vzqymSeeZeMm
Pj0M5XD9JBcTx6WlNBKYItoi3btnIGFwoowbkFuWLEZsSJ+kJ2kOHUTMYAqp
LmqmxtkOTbQaHe0e/EgslGjrPbdWcoC0i7Hp/Uckfd2G40s12bI7x7h714cS
ROeUWSF1KVwUZYRt0XP9ovE9z6iMDxZ+6ssoscz9YX+DyCX5e4mKyiPNu+i7
ZGJzVfqMh+BAHkb5pvhIA3dr14j/mNFa7/3YJOTrvyMbx42p2ZdyTDmasF5q
FyDPm6XFsfLU1aNzmribWfgFSI1EZYVlHd8VG4fDGeNEchBMdedq2EUf/WtX
nLutUB6I/bjV7GYLQBlHc2DJk5+YvMYSD5/7Yya3FjFpMXu7qn8W5fZvLtSr
bbRysa+PP1WFiv/qTNJWJKYu7RRC0L/4krqloxTQJ36ici04RvU/ZWFKQQlV
yKnikPOR4IyfaSF3OXBTxbRqDjKsEcctTwaoW2MlP1dKkmEF82NxJGKUMELE
6ZIuFngh4odmV2zG2Kmtmj2VLozWdbkaXkCjIUJmkhkN15ETljytsyWw9B8m
YKgdz74d/yqjQIeHzwmjccMnpeAEtNmnjeVZ/HJiULih8rBzkPIItJmTTCNh
u5CXjiwgTFOoEv0eZ7ZyKifGY8dpwbERYNE5pjzcx6IHNIy8nnBtQlej7NgG
ZCQyQPyPotNPKzovX2v17FvZuX1m08Fm7HjgvMzuRjQPdz8JEfDo31Lgxjtx
PfOY92QFMBngCShHJ1em0dfNtlM0tBO08M414EBPip9otFHzTV0bjFe/RC+0
UdUFKr7cHla/+sWc2yHiKVsUfbkFX/h+qHhcgSilTvFra79G5ajm7ELceF7U
oSTLxEUrZGofLmfsipG+3AJxtu5qxjSCdj429QxsErn8Mzborpi3hm5ebVyC
tLvHQshfvk/kIJhsrOqxKpQX64KvpqOlW3FaxD5aNUAyGg0FlVlewEDaA0wz
97QUpF7sohWDI2c1pVWf4+6TSuT3SgkTCxkh7csrrFkdnrhzdOX3MzSLRXds
L7nL2Kk4GQT4zapLqTxI9/5db9gTprles6C/ATp1EJ/xhrxICR6HlbORaWK3
4T52itzdvt93H7Z46YH0uFEerr6A/yNqygIcqrQJ9AuONdrpha2seYbKcpqL
qg07cCOgfl/aF+oG5Zjx5NfAkTk1cqWq2LKBTd7s97Lr6yIub4yYe/vmnMBi
jcRCq3LU/H2/4yHmP4MJHKNdJGP+nhwI2EUdd6nfl+ZsmPjL+v/1jy1To4id
c91wiEMjptH8eVcoYXKEjHWIfhPS40ZeJgCbADWgFHBGBXLusDRUbNlyvObD
UeGecDg/wiOtjVXRSWt6w+dF+Th8gJqo6gQ0URtDAnNJbMQ2XLImV9dRCiaR
T45F6jV9ATj77tMR4i2Eb9CaBcbnFG29Qj9eprNf+El3ryL5cxphI/gCxTU/
+GVZFU8pal7eZCYCVum7gtQfxMxUIcEYJ3aY2cttNPCFUP0jKLdQG8WcBKdb
HXmOs2iYUIBt7uiZaPilqOn9u2Wtd0a31iRoF0fqRa9MWuzKKRn3pQ27JAYC
W6ES7+0ookjiMqa2rSVRh8N6OEqfy+nFveTjzhOi08cFaCwsn9sVdQp+pFDH
XJQ4mE6MY8DU2M9/Hd1XC4bCyztNNW0dMiZc8Ov0OY3724cqnZS0VaX9uNNB
/+fu/humt5OJUPtdv8qLe0k/EmpytfBvnm/X+WjTPVvIzsjCs0Zm3at25gJi
WIvU2f46bdGCm0tfk7lUBeISkRw8tU133aqIKdrNpZYZZX4c+55FcrMPn6jQ
vaa0fR7oA1QInQvtNUobUfN+RB4y3DExLjNhzWTO4f4TU582Ochppt35Z52c
4bwaU+Il0KeL3I3sS/327M59Yv91sr4AsBCIFwG3fDbW9nMtWTxDogmcbfQW
vz9CQg8WLD7CB9zA8BJg3HB/HQYooKbh3SptU/TcyJb2LzWgBkMhaOVDHYqK
6h5muAmcomlCxn2c1VzuM2F984RaQWEzCgw9omX105glsZQB4j1puwg2zNmk
7iUJI1fLX5Smrw0t6sgKL+V+MiNWeyfwcD0CiUMrV6Xt44JttA7Fh0PnthlX
hbN2vHo4b1C5yTtOYPr4Vt7c+jJZbssdHdN/F/4PMv8S1gkKZLSuoPA243Xq
/VNo/Oixd/48MQhoPe+j23eQwpwtwKd+BseZ6a6h5Z6klayx0tKOIMqbBgBP
4ho2grZDL9ee6yW0BsBa2NEBgAhdA5oGIAIBp26jcXz648kQZhQLDbg5bDvV
95XplT9pw15IkJiRAlvfxxlOIXtv+PEBa51aUqmTtydmvpl3T5eQOiPtVrbb
csmu+n6/WGaAV3ZSAawPyF11POT8/1WtNCp0ZCsW0gOgN9i/adDpD6MNi8Jb
1HDPwVW0OeL787S/xc18apWxqVsnLhLwTJftjfKikEhBqHqeTnDThX2NZIkM
nDUWlIEgy7v6U/bD2S4qNBqUynYaXZCWeJHvuujAxFmhB1uYOQrXHL7sMUQh
Sk49JFcD3TY7haUctjbkyRPr+TCtOH82I05W5mNczUAt93Gp6M7U0HKPPm4K
tr85Mz9VP9j8pBkwDDgSSLUy3Nm1RZhvbMY2PnjlFTzEqlBWC+5j3wFGSXgK
AOg+hVv7bkW5BtsVYqbfeoNlXpB5omIApHzHuKpgTJ5VQ2m+1rn8Vzrwj9IU
La7wCoueuo4UTSjyK8HS2f1hgu9eapAfyu9DcFpPgVriiFvAGrZiHICVnzPv
pn0wFKym+Bx3IZwQ6x6HdXxRNHox1Ff68F0ULJQs3b9bGElrZNwsof9riG2C
HvI7U/K6MEkGxzBbVhxesx3OY/dUX2XGaHrEF8iNU38mYu3G17DexktD5LCF
37LsuuWsBvSN+yTyd3bNwIoZsPMn26eJ9QhglkGep64gd+iRnJdwoqpX3/v/
HuLpBjQf/OC8cZ2J46CTx6ln6ezJD8UOc+ky/ZRfuOxjBAbFPXYuVvWiaEAk
u0tj3MTuZHeXJnyYN1uNBTKtYUOE7FHkscfyHtDgIuHnlxmC+1TuV1acZg9Y
2yNm+HdNbfiAPSyWGY9XgbvI2iA88EUwwX1SWaho8rYNKbkN9cAGgDETozbw
OgMYuPoWIS2TOYwqlnzIzW664JUhbqq+TlWQ0N4wgaLc+KWY6agbzI9UCaXB
2AyztiJlH6A8rjCInieU5cR6+kYOJpg4XMd1Zx0kex2rIgw24GVq/25HQsd+
WRpCKwPqbVYpbaDiEDK44gIwtCFM6MozePYSvKp4gGCSMa8pi0uApFW9HkaB
Z7JWU8v6EmTtV1pJEsGUlXd51FKZEfaI3mgnPbW+DMhf1gUQ3We4V7kMqMPw
2V5sCagR2zSm34ZqC5mbA2rflyoqyk2lM9mJjUQ+ZGfC8KXh1mcngPiyW6tj
O5SISz9yvx6jBrOwR5u2BVqwtoTRji3Nk7LIoAM/QQjM2g3fmAjBZvAEnSpz
M/t1b7xJNmAgC3slAs+4C9fFgXVfduR4P0SKchS46QOhzc3MfyUZnfV4zPe6
tSzmQh8/adaeZKHUxTaK8qGG9YPxRltNvU9fKtjbebAKwao0VAlX8n2SV+Bv
Y+9H9pclb7Zy8I7UEMXgCjc8ZthcVkyMCVBsLli+8TyZTXJ09x7nGhWBgmMc
jSbjOYrQnmoKF3CtpnpHlfV7X9r41FuyjZULELfsXkx3Ig0fhZJN0/iwBMCZ
s/DEUs3voLPBpBVEwc1SO/I8TB14c5qMB/SyW9FGfYZGAuHuOyozWb9QjHsZ
U2PGjEAhoUmrOD8X5mQMmiej/NMPougcy88u09yFo90Pq8+EDp6uQrCg5V+E
cweefdDs3I3/t0MjhlMCBQqbV3+FEU/ujzH4kwl7A7gvpmDWlny1LMa1wJhb
IU19Ox8ny5z0MS30GwkhVtTVJpDcIcjRtZeXtoJTyhkxPdREQtltSqL/zrun
SgZUAA/T4dAZ5rLgbX0+VwgJSOWjUMV8gxAID4su9DiWZxht6o2mtwDVrjMb
s648nvOoI6q+04hO+2bHaa9Pz2ULcnZfwDlabo3HI8959r1NqCE94WgZEBFi
v6F0+uBsJEK9O2+bCVCJIA/Pg7t5ux9hsqEhH0GVoztOxsRp2iZ+qpaXVcFm
Wf6DoV9sB8aeUl7+Vee9cQKr5itVYyce/xKpHRarrZgNlLqnF3IeYVstFt6R
5Ul7qQ0o1QW2xOENEHRNTOM6CZ1xnBUasjRLgQ8LCOXrAONpcdGOTUJOW19e
IGdsM6N55k1pXjgb9d+9pvQDlWhEhRVwUnaBrNxG0N+7YAvlV/OqtHuaoXQG
HU1k6vDUmMtAzOVhyQndi9up/JlGgHAwB2OKLC7ny6kBI3xGMJvywJYFwF6y
FR3XoxIPWWM3grN+tVApUodObQ0x34ZnpRtxGZFP2kbRaQ3oKvMnj3sld0/i
OK5mgrEgrXBtzEuqN66M7V7E1zSqYBAfLoJ2qz4p7CAgmFepkicD7OR76kAA
KDl48E4bGdov5NDcKB5U2tsAM/KGuIoX4TvRjw43SdJQHoURd7eUHO4+DVjA
s1cTOWU7hjZXq+WLGC3ZA51+xTB5zLYUUteeV3qYAi5hKZwEeYJWGsYi438e
VmcW5HOLdEpOerD39Upy8LiCZwp973HSZVGI3cTz8DLpwBTNJsBqCfJXVFdK
QRUcZrRV3rP7hlgI1sJxjAzrRD5v8KecB8Yr9tj/gvXPIoET0KuPZeoncjqj
rKFH6Tkjer3wSGbzevMmyazJFob3gN7XsOoyeK3fr+FhEHQZzTWDfHLqcLWV
MbsNmdZOcHVII+vxrxcrOznrsw7+Z+o1OPsFKx1nEMFI67oib53XZwIJp9qM
JyRLi79YkOm1ZbCdGHBrZ7KKOLy+d4QfZ9rH9d+W0pi1x7HC0kmHCdT7ftf3
yd1Ze5lbdynWtxUIG4MEdrpehb000shDK/83Eu9LNPQNEVvXL1SLrVVHIU5x
Bka0JM0VFrt3S4MVO54N7KV7o88QbBpMII6M0ysfcagKj5lEABLOmMsNpngv
sLN30QDbSeMc4yEWD4R7AGX03c1hiqTP+sIWV6SNAFy1BE1bK2yvgPLh6Ey2
VzhS8Ea2Cc3GSVqIuLhpy1mgdnSxFfqARkP1Vu0q1gae+OpbpvGNO3eS4e/Q
ClFp7amnWS+x6/pYlyJO1wOdcpavphFPmxHz+Ytuai5EReJ4txJP8wjP/MG2
9NL4LyqDYlJEdadSuJGwgMdI+nDesGwQhpYkRdPNaBej7ZM6rzzh+gyLecFs
Fzdnm/NUnzcLgaQ8/blSHbrqNnMujxblqOhM2yFi16dvGTT3ZUzrynFzQSE1
jOds2hhNwOS1Tb5QaAGKZv5PvZfmfY3elMf3mOO8z1NZmOGsfW3Xy3aXhdio
4ifMNpWPXemCUA5srA/q8J20vBQcck3XhTxvf4S3ooiDagj+Hb+7luvaARqh
EIwABkuzh4/ku5QzOPhxR3d/eeCxd3R8z6GtRm4AUpLHGRXX0NmFG/Zvgly6
bYnqWf/qb0whCkQLykZhyJksKItVVd/LdiRGVQf4OEvt/azhoiiPUmStogxI
o9OKZiFxzKWXo4VPeOUNO/BkDjcPNmQKNKtUAsQrFUIMD4Cv93Uk6oUof18V
TMXLYETwJvWVzyPbAo1yZKH5QncoxQy124zkf+AkGYynftPoqF8OWObbdqFr
v4zd6phTGtKBO9JoJ/SXmgi6bdsMOb2wes+jcyJccASbU05+2md1A9ApOUH+
jeD77QjQ03lMGd68k+Ci/U+MYisLaFuBxvKsXRiofGoHgL6hQC0bsoFR5/yi
Y6KAve0R8ohzcFE5b5BeG3YyTesztVy6AgChKIkbRSClQBS0diW/9ehhIXXI
5BYsotPYsYsE8MoowX8Na10U/S6Itcd99Sgvp+8kCjYT2KzgzxLvPY76Swe2
PqKJJySmB7/3MfwvVYAvnhfcZZ9UlI2XjvXvWYjS4y9iHG/NJBUQ/RZb717R
/2ry4Sb3APROfQt/uV1W4Hhd50jJrtNO7dggi8f+tzj3H4l7jFQsNbn9EFiG
LKwEviH7m6iC670/K13Dn9TOq/PK0J3OeAxHAC0GXjUKlBpwlwu6zYxzkrKY
Q8ZTLYcyjdRLS4YqLRpwaPpWQ3ZD64Bqp5LsM05PfkU3FN+0LMrsqbp4oQno
0YKtHUIwvYj2q3bjyKAFrA0Pn61zh4+DfnJDmhZn1dzAFxPnNd4ow6pDWA60
U2BfZFHoWD/j5o1yKtKFb/FfFoGrZWNHezYKie3F6+ocl3TBYyJdE0GnSsXj
DlZSL2e+vbM1Cap4G9cLEPW4pQ1GbaXRpf4BcsXgEC97o0mN2DeaAj6r5nvW
9GvTlqx6d5qhB/0mhkMy7Ld4uKh64V4gFEWnEu+673BbJ0/8a7zF3wmJmK6Y
HT4WG4NnK6vIIaqIOBSQAVrHodrc1iWHtwdOmIr8Olp808+lbJ3EcL1EDvya
Mpthcz7ieIkuarTd05VWwIv9fxfl5JH7EkgxEMfCNu3XgEv85GuS+7s2hWWg
rjkCj9fPyarDr2juSb+8wjg1clM4Oi9XubqHGXL7gosiNsjIiNcrCCY8e56x
fH0hkQQTFZA+y4l3IbYYSjjx8CsAUxiX3TJ3tdXXdKUa5Cj4QUi3UcxO2Vcv
dd4c9qxUzjFjoYiD3Ra+RfU+fnkMRwtvfnFzOt0uRmR1XrmNGNAouFNcqYXj
tZdn5C8bC/rCDScLQnLjqhjFHvLdKjrJ8j/USrmhr2w4WNs9c9J0IyvDFeMW
0vs8sL05EZHpgAeoyXzl6Wo+aS+DcyJiTA3Vct5VNDl2N3CFYH/+YKc6zERM
PU5WTOr1tyxwrfqmhNXWYEAHWWJXRKvfTlZV2vMTa4LZUMX5doGxPzyl9Ju9
HwOG79jcK/3xZA/n9KYKJ5PRMP3Ryi6ox4nl/Qud59EzGFsvzRLFeEHAll3u
ZYieoMV3QoRC7wDe8+B/A1xcA/NMIwJjmbaYjK0KhK3iGYcg6Fh9xHyWNO7C
NK8pnHTilj8EBDoDron9xhC0CDge3LwOjqU6R8k3GMhdrlHD8DpKzqOaaudV
8yr6zy9TTJoEtT6LIeSRBHEE5yrrYO8Vef3RBD/VTQwA+8WMblRjpPH2nANO
YLrkrgxPs00Gq3w8vdAsGRc2ZyPCquwRskBTXsUqHebGgiJL/N3h3NCRB2m2
chYljB15qN+RIRNpC4lQ6zTueDEYZDr2eI5AVSsd1YKCm55XlizAU6q2+e/J
aJR5NFAiSz0FxLBzlmJfLvBwNVu1kjO66bg1bS6UuEmA/nNrlA1GJI+dxgkn
RgrOfIfsfLtk5T4fYiH7SEEKsKw56adeFe4ZXP7/f7/onX6BCoYemfySXyOT
XKxDb9GJPADs5y1rCUNZj6U84W+QpZyEb+vb3rHvGZ6N9r8VvCxxaPsd2T6p
qbb0dqSnWVR5+Jr9rtCg5vy3YzgSUMBZywKP2/yR4753vEN3dhbGV1u0TbfS
fyqvKA9wrcVV8zTAPcDpNqTKbC20svCycalKt5ZOLeDiAfl9LvUQ7crr+xKr
s9AvrbTaTGbp8+uZ6Od6tuXT1eKoO/PcBvvOuMbJVRz3hAn3F99LfgzqlSJF
jzi/wAMZbV2wj7JH3szKO7ENBNWRfQ3XxAkeRLu53vnpikHnb1SffQii8ohT
hDBI7imKwsGR60q8Q6pGSbxbto4pEt3a24Pv8sV/LVd22CybUnXG0GJmkHGO
FEutmZcejLl9/TM0KCqjRaHR7RJjCakm4M9BiojOR3MTY2Y/iSNIIlP2LxYt
bLInn++EVcuRMiKUN8HQMcykV9NjsdOxlQzfIq5jf/Lpbj054Pj+NmoIMm5s
tRTTpHwwNKfVjB/CoJgUzkDuZcdJ5jhX4K/j3CVhhUBhh0fbTGhSvJqcqPnv
po9zrhgImB/JEpVXQU/sZM845aV5KW6/IkHt+DP9fC2OhVPrvnQsOh/NwzCZ
hkugm/CYgkYN6L1Azjpdkid1KCQPvg0dxFuG+82851M57uwmOgYuxqq8Oibz
dpFUHhXiJv0pHK8kn3wduMAK/9LFG3pewEqfKCwIv7mCc+d0OFF3vV9Sfecx
jAJsXiCgxmPCbgXANtnye3MxBfSG+cUt//IyTgfMVyoFihAq3VVb2xcpcF1x
RD4j7RXIN8SayeMRJ5py7RfYirtDHxlElaNJlaIalDrE0fRy2Y73x9pI0bod
6bPJspnQqx2DYM5mmYHEVlkFFuqr2DIE8kcTzi9FdNVf/H9rqOiLsGT7hgPs
XuZj0L3i9hM2VCdgjOld06qRdQCHpTmZ19o/mDXGucOhqr01l1pXSpyop7Dt
9q/OzMZ+3I4riySMpf++OlRNNJO9g14blPEy/L+xR4KIFXhCB9GuZD4ry0gb
EI5fHwsvfukW+H1or5AIObsghnLPthOZvJuiNQCQYrXj1TJ0E8BQpvCHO1+i
LBsSbu10bnrfmxxmZfkVcQtujr9EVpJ8r933UWkWAFW/4/FipGDl27rkvLJo
p49gz4FP4UtDQcwMCDyBCoyZm3ipQQz+MX9elgrUa1c7rC+mLbcUyOnKYiNU
c2+nQa+FldPhBUU4PJ0NhDzYv6QSw7eo8isNujPLZ0q/JtMrP6Bvwzd9tHg+
ZplwJ+10rcyymS/GWcXX0ndGideZCue4khSibR9Mif7XiITsavESL4twa5at
uKHx6udQt5WSVz6ZBOEkUE0ZQ0K5ezqVs40s9QpSg4qcOkZU+0pCU/G9+btS
IA6OON+LLKbUWL45OOv4+kIZ4Q9jdkoA0I5ymndLBknrxucpGCyFsT3pSRQg
t4pTD/pJB8o7Bnt841eZ1k0PxvcrtXhbgSEaJ5etgFYftICwpCQEJvj4LaUA
HihipbAdDkkeJ5bWjFh379gq3IAUH4+lxxCllS91Cqf8Fk55IwzEFt7Z5eQz
n3THMjTtBXuCCRZS+jx7bplqbq9sIX805OMNnduL1rpkfcvcqA81zy12ibQy
Y6bIPViEpbRbj1jOtc6mT9wMjSi/cejA0mUWJP8fIlUkXXk746xtQ0JikTh9
WgaAPCjwJjP0AxRqR0xGSDAEJSRBJdN1gy+80lj5u9oJzy0CqhlY7BAavlb7
Pt36ASIZaI6YKxrDz8DX8Xd/jgQsDyBYvQ0NCxd40QiH1SsN8eEvgzmGooBc
uIu0WoQ4wfEB342OaIPmwKtf5FYJqAmBVmZ5XDCbiRvFTvUgmI7oEMyB2jkC
DOKzN38dsAofB7HUvhY+AGAiTFEzKxYEbxF7vVpuBddSFlTtn7Zhdi/nTmoU
5tpwmvihPGOmsW26MVIm249nFl5P74wJyw/IPRxUly4Mnk17TxIj5pA6U8OW
qKi0soJigpEHu1Ovo/rH/TJtwgczM3KlaytWSQPEETG8pEPOnNWSQu0S/+Km
JFMS9rFHrg4/xEe8uF3gu8+qxyrCfYVPtpBO5y4l0/IkpFRfjF3yCvlJaN90
vqjpJI/Vcv9W7aPAhlOAYZak6rtTLBReuf8njLKax3UPfYKH3IWKMe0wmENu
UBl/NXEKqWsyD7Vc0FX3uNovTQzsOYoxAY9jeq8PYbnoSYMV6IxD9+YzJZKv
x8JltzjtnKfloslXw3vlgwoiT0ThdAG0JJU7OlWieVPgVEELk0/xJ09XMnm5
2prEcUkHuunhKVYduD7FXzWyT5r70z3/H3zPsQwPQpPb/0+7wldNdQSoX/i5
1FJXHBwPv4AO4A2Mjs7h4se6cPpoO+pDBOMk83CoLCA+xeVtmQgc0lSfgLkB
0wThTLpb4x3Mp66Y+oTz7Tji4XcqDKLoZPUTkGzViP3hiT2yqKbkKf2g6PhR
p1ls+X9Aitn99cs47TaaRa8javJW+4C6CNHOdviizrMkKiwjk7JHCdpmOhHv
j1fSAdxl/xErSRAn+PQRhS5lzl5c2gMvdfcAxpF3CtCq68YoXJseONUwNaBT
xTdiHG5CRYvjTu+HSEduAuetLnd/g8oa8K9z3ag89Z4GXB445LB4N4Ty3fRK
DKlG134Xj969N+y65bgU2c5NuIOO0RYFAreambwZo8/7Zu0Lq6lyiC9fFsfJ
N33WugZgL2VXKPa9Z0pzamp9UZfnOeIs5xhi5qGNxWbB7E0ycqrhV4i2urYm
I6sREYKIbbMMRSTz9OqkrKOnsbkq+/kOwX67ssap1CbzlFENKnbWDzq1mLq7
t8kZfDoRkuDTx46X8MG2aotv1Lr2y6zxaV8JYCQQoquwdULYBIh3yp8ia53H
qvzNdq4xSMIEihuSb3EykToc+syS9bckR/f50tmayHN4U+874m5Gmy59Xd4o
B1KTl2kTDBA6M1RlKoxDVJMn+F551RTQ7oHPcbk46eHSyWc4gvxdUg6TIvJn
hnlSDH6dpo+j1XUuiJ373iRHTqatEk26cXYFCLFvyLwbSH8Do/nDqTKk853l
4s9GBu6352TJFP5BnLy7H2wDCtQNN2nrImYtfLAETa/6H9JETNSWXFTpSjFF
RKu21MjIK4y1y0NW7Un68BGVP6wp6RW/PmlxtMLxC0NNrmrNrvxXerVtZ82H
Nh9DiZ9ZgFqnBBmTvu+mpmWmLSzBLlE728auBKqsaHstvjsgxVhSAvgfiV2K
ozaQ3tUjZm4Qq6/olzXS440A4M47nOnx5xfhoghdxS6O7c3nW1YmVI0p9n5q
TFShkalgggwD1I/N6MQQrwidQBM9KS64axbBfQAoGFYTjJuG6Fx4zSKl6T7R
3VYzhm6Ezn+FZOL7I5KBnjG8OkCLcJW3bRukHIWcuD2pFfg9O8A83RAq8Zmd
A3y6Cjfyqwk9M2Zm+Kb9Vhwa1r9Z8PZcPzHUpvEA3cFFsErgzarp6jvaQv7e
eRl3wclfysnJCoH4NtAn26np0k2eMGLCdffTwwW+hjTZdvALst4y3C4Yq5/j
0LNJwgK2yFwFtPnan9VoQ2cOetdxFxSwIzD4sdDUIcg4ajpQLNNmpQJTrq63
i5M+PFJ6Z9cln2zQ/T+Qayy6O8leJH4zBZHZ4sn1AgeNBdFLiOs3fU/FH9Mp
ycxRt/w9pTvQcPbJgXmNxJBwFVjZr1Tku2PtbckmAUd2OFWJ+HJI1zL5BajD
qo2USJ/D+AQllMfQUdhthEnkf4dwkbiD1wNVevsaXrob+XoqwOqyhXOgBjhG
N8QhZHO7WzvPNG4/tgDAJ6L6DuV8Tps6gaUnmho0lDMMnUI8HupPXdPBEwsG
WWZSsyqfBCr6g+C/uoyBIzTverCzzzQCARotsBMApzG9BwJOnuf9So725/Mj
jV8P9ZhjwZvIXfCyd81P40APOXFEgWyB0HGE9V/uQfz5lczw6ynwX/5eMBJJ
bVXvQibsGdEy3vvj3LTii+NmLycc/u1xHzgEonGP7qBDTDOkegANDuVvKmnm
DkV7A/QZ6rCamNHDpA/e6UJJu0vORmRl8S7Mp0s2eIOXCydbFmABGY/oA12v
xpaNLcVTpXym0Ywgzho3VG6uEOgX2zH/uBuIqQl49zPz6h4ZBdQQgiPdKbjj
su7jX5nT7X9o0j+3q79K/ccK+QHNblp0kaHDTN4+OAhSvG+JaR1E2XDn/LyH
K8mFRsJIn7rfMSw+/fZZ5QnXaDHVmNDIRunaqqVMALwrwVQKu0IZ/oB/upcX
AaCl9/qh0A3FpU+BKjZA+7m1aZrqCzd6v4Rz78JOgDH4g8E0yGvl92wssPr1
RxKC4G6iNDCp2RtTcUfcwdtP0FMajdEnPELH5mp2pRYWmauchnZi7wxCW3kn
QcvnduZiSdhP7lqDB91f/wPhScytFEXjb6rsT1ij70FAw2nzrVFnX3yUiMOW
6Qq2oA5vIBk4o03RDdFhZFC08+eWGu7Glay6FFJWvEMxBmdD5r5zwjDEjGCI
UuZ22Lc8m8n+B6lXM3CYHDPzfRuRXDFGSt3KF9FmEFrjnkQFShY44GheURuv
eO/z0Ioy1Tl+h5DHLdFZ65Z8FJXR21cYanTy7Cf2FmeXI127dtvqn8ec2Oqj
y9XMS2X1aDMz8Ce60I8uk1j5CSa7X+3OuATDXH3r72sPXkOLezcNM6Nn33VY
/ObMmMvjVxDANnZAbCtzqunGbE2vyWU5b7AmbuJgURNZTLxJVgIXpHRNPxeC
KJpzcJufVFV45ilnvJF5iq8ND+QWTUkj/I6zICiGDdD26Dzx4NNZ9jUlsZv2
8AP5QNEeqDr9RFERtCLRiS2BRTMWrRNUNuxy7JmZiyZUPxDpUQqPAfuVkUGD
xcl43LjfduUyBkIk4W65DUSafxInvctB3+/lz3RQLIyqlVvv1VYTjaXWkNoM
U8/FUdyrKfaHhCkdnUAOIECNGkijsLqiQNYlQkFan/prvAwwY4qv4HunC5I/
PVcQ7szsU60Kk7OgwJEOnEaRts3o+VUgukfpApOlmLmhNFhWx3cCCZmIorPl
/QrcHxOj9zyskO8rL6O7GQ12EX4vG55UGbAHLpoGmOuIWEHiqXl0fePViHEj
xxy64iBDybVxcCMDRVmx2wWgpOfRAV2sDJe49me5kwf1WYZrA2awPNSjr0zk
Mt2hoD5akGnlhn/MmgKjlVZhocOG8bDl1bE2cY4L2pKght95oRTa1AmzAx6H
3bh9i8kC0AY3UL0xUwKmBHUfLzrk2CwVnlw2jrsU5s/0c4bUPG4FSPOK5mKb
higauTL+445nXUFiO9YF2FQ46N7pL6iA5OugsUWLY/O6KPsz0c4HqUzWOJUc
D2sJ9D389w/qKQ7cLohuzBp430fEewhJ2zSCrqI5X0mVmco5TnC4YD4BpPs0
qDfdwN7rBi/TPjw32IXgNWl14T6ZLNnc48cW5Sdl1HWaAeNF4LYjk6+AiT6V
9yuoLyCO9wiFfdiFlLsouSm5leBAazSUHvkfZGqot2nXAwsnBsEv/sELwSYP
MNBZ+66aCmo7VjiZ49Ho6TPPsIXbpzmCoabQuPrtz8DHJ35gZ601gFczgyiU
MbeIXwAdnT0mte1Lt7EL03JtxoIM9DZ6aksamm6ytciIu3N6UJ0pYQadIknb
qdahoWuayO+VAkbJfXCVVPAFluGVCV1TxixXmthfozXN8QP/TthMJnOJi6gI
c7C5cbVjjVkeMiznDLWnNzVZTRXz+OBTNUyoPmwQMmfA7jbWXiZxcSzrv5pB
nb8wFNJh1MJwgIMt8kIJwZ0/tly9yOilOIAnrEYGDzbYkg6AVYMqDtCyXZWU
TrwG4VfCN1wWflVd0+rBEUSyLydAXmYD6KktKjsQQ0qAQhjlGBaDfYPUIIvx
vgtGf8v0tB4DnTiW4FQdgpKu+JgdBea/Kn4q4Iyn9l+EfrWy9PsvScHBfs7n
Ff8jX6CN0qkwBfmh8ML17PadgYFOiSLbvYzmJ0HAzzngGOFPO9GPsHCJdQWV
8vT7N6FpS8Nch74BR/OoNURJ1dRJbjQcyVPih743/0/7wXrzB6sCHxLTIcFi
OCHQ8Hnr37RIOYlp1TP7dTF9Ya3l78qR7Ifu1mNIstfDU/TWphDWkop7Pc0x
Grc6Iyy3Nna9hicM3uZym1QUZuMXo/TRFdNXywMuiHL2/t3pCWB6mleq/iMj
fjzskwp8/g5KpyUc/bBZqb3NBbMryXHJqAWjpgSrVUQvB5ITzwTl4OLCv1hD
gjLuR99ZI0oMlE7YCWtdLy/ITzX0RnwI+XKRHel7iz5CwSwb9D2HrF0xJnlU
cIek/SQ+P11MryxUvHmB0k3f0OOhgRxlX+RfBN2et82KeaY7KdKV4IbAzC/c
s6w3A6ZjTVTZlTpPO1S6l7QlwwBwk2hP64WKJlhaQ8D9Jpd7fgQRXsLwaIg+
aenArfvfV+VF1F12e2uIWxk61LnrhGiS6AFT/AEBQ5Jy2+z9fYgdzRgFUHzp
rt/lWL4zPzStZQRHQ/iauiKgSSYKQ2xlAB0eZGMctiZYERSZV16qJgd+rkIl
nm5CKnpcR0209mOTPlWSn/9lho07h3PXSPmzr1dI5lwpInDMg6YPIJpOJNNQ
qSyiJJsDGNtuqLyObu0z9iBNOwUZRotl/pQ4IfK5asaTkt3dCrxKUyg7eh1B
hIyT+07a/H0h57KGXdZ+sNHD8eQNhC69jjAwQNEs49j18HDe268PkQU1qLP7
EDEHj0Kjhh5MdZ4rYYZjv7ZC1W+XaPFBZcM8NSU9XGtbxslt2AHgn+IFpL53
s+WZlRNCuwGdDS37MCbULOm13CIjQazFNRuuR9dgOEgsomwUcq5oAXyXumwa
Jn5vRzbNc3RkcX5M9xIxz0EiCI0vxrJx3PmVGWyfs/MuS0k1DixcS5qS17wP
rZwBx+s3FtaLDNRn8Yck5mS1pvNkCrh1lhG8FZMfbwsFuyXUuLbE0iLq//Y7
eXJ0axoRdehqhv92j9NjjEV3GB7iT8SMmuXI3T2KBxAm9akfPcY4DgxZPs9o
HYwmZ8ak0wL4ccxarUQZWLYpr/Mb8P+Ez1DHAhk+zltVBco1LMse8LMY2gw/
+mTGO8bYGMgXZfEnIVBrbbAYmYuHVTSOJx13dq6wIpMkAzEDUOETqoBsxiFT
tVh196d6kEecJ6rkWlvJJqdbKKbahctGqFX7981K8DOXqm0EvPQNOPuKPuoV
hddjM6/01oncUZTdefqEfR2rNuz1aAvrYoHGL5QV02CI1FrzTBeEb3RPhNHM
X2ewDqd2BtbV/iQdaFeL2UBS68QzTgoISitOHmhaf7eS+pFwtNfPkZEaSSQk
ReHxnXPFy1HjT85LFIGi3tvVhwbuJ9lxWrn/5fWUF2XFA8izp0xUL2LtYHw+
PTVdPrVP0mI7TwGhNIBrlGM6ELJrThw3C8fgt/aCFgt5xDuLlRrX3CWoVj15
fIbnfHnBkP4dRuWeQNqAKtNhbbCgM6cMxXTQ+1r2u/wHjDzJOvjGobBAVbXy
nzoCprK7xfyCOA+mWbCHfEBRVOcxoHetqw7pIUBPPpJ/v12Whf/ATak8ypEM
qSuF/hbXn0SdoxdDkplZUajzWc0XSlGiXeBosYlx+sqcULqg7NfZ7+1b7Pz2
/UCVePxmb8FbUwsUsyaaQPhhnZqnCe59S3eraVaA99387GCVVCiutnDJutoV
ba9S475IKnQERDrT66wjaoGqMAa3HRA/FZ7JKyElPczzqkvajD8/d1aS3lKR
7BwAyKZB7IOX7bED9lWDEX4SnIrG8qwF2Bpv82rUA8+ZTbfXqng1WkBVEnxb
Co1Crm7dK/mTX3RtlnDhrZ76SU1ucUvagHeyQHh/7TvMqkM4FSDAtaAO4omj
L0UIeGL+MY4niyd0PABXk/VKeyZxfCgFA6nCQvER68TnhmrFmm1IxP14xaTI
kji+ynf8KJljCXQILbuc09afPBMQZTlEJx/R3VeddxOoqkB5zL6jBTkrVZPI
teA8Ge6rBixe8fuAhLIyxGZAci80EmhaJ+6JluyGxyM6xCDbr5oj25fNfF5a
Cn4t7sIZ80vvlk5QqQrSqCbCVUe5qIpJZQntAxkKXFyhpqveGM7ORNO6lFGY
Aye8VQSO9gvG1UsqvJAcI0sIJEGJcNcm5aPqtZng6m8RJ3C+Rw57OQUCfqD2
41YiXSD5K3F6I3XK6lVqJtDBzpi17xiZya9IiX5FKe01yXosJYfOmVs7spPU
kjZz5LcFnOTdbcUhOvmmH8FR21GU+5gpzoxA7DSsT6H1DfUv4DAmUwnWAJ2y
qhfDJStUJf1XReQn7gSKRJdNzaev0j3D3asr2PO/dTIzY2v+bJ6SLltKLayI
9I2shwemlv8UdbAvzD+Vv4UgVIISftZ/7/wHb2sN0NbGplSuEojR68dJ1qjg
jzaTVm8JoVkcDBxcz7TKYTSozJuL9x/qSdByIOpYCy+PmXpcVsoOR1RM3bs3
gy/3+rgtH0G5EzvaF8g9/7iYkKHlSmsnZFvhWiY9yaEn9b7fVBgAsfSyRtBE
ldG1OX96Tgdi+r8bsF5zfe5NsbOsKEixX5tQqXOMkZsknbKEi71RfllA1wl2
JtreHViAufpUs+8JCDzBxr6zOSOg9OECtOztXeTtJUcG6uaj6V8Dr/weWVHf
+/qMEmi4XtlZGfsQPRUpA05ZGRZyrYit+KFi6pszE++/1EzIOGpFU+wRoCmK
OJ4Gbocuu8nBaffYuvSFFXMVsHuWnwWaAg1TsSsqhUZoaTnEe6h0LDM/sE/N
eqUf9q9D6eAdg9/T1S+SDpDSUXm6z6ElTeGpR0KjY9z242YQK8XHAssAIlNS
42kFFu0xTjIyEYqQKqGBbW6qdBpHfgY0nPgt/NNpmD+a0mKh9c+b2zj0EU9y
Na0Bo7WELDJFqL+Rq+RVRw3IJr9kPQeX/TNg38+LLLAPlFpX6a0N2PKmLDf2
2FxYIGKDaAmoja2FkGKkHrzn6B4L2MVHIZBdW86uNwcqMOZEQAwWfKUhYNFf
ahCLl6ji+U7BkKCpB8Vtj5gEIwZunqZuV3X8/XIEI2oMXGkN/gCPlSOeSRpp
NcaXNJsMsUccM5mPPZyZErRKn5qXGUTefzhRqo2VAfqQftXqNMQJffU5o55U
sLHeEDmbI3Lx6cG35jIegNwSkNK0XqgDQBtVsGkMdWckcni5LBoCmWKG2DtC
Ta6Fvw8bEq9qMiOPOINpJgfjUKud5CiMQYJPCgjRpo39xLDcrdMbXKKLTtZd
LtMr2+FargEVGcwNuH/nqcT+8Dpx6wFoEKH5Zn5Bg5MZHTN+B3YlzP4xttMY
/8SBAMAYiL3UTEeFCaVhlexsfnrOYuVmQtSgcCCXbq70bkXCjOMcXKVJzoNc
KWRto5p97wSdBzQc+SENI6J6xGGhltmxox7lwvNeIHYXih/y3mNrcGM1i40o
rI+flhTZighqGOAHgJ2oYH9S7pEXjQfwuHZw4hKvRgIBc+mToHP1gaTQSpHx
lkGK3DcWYMgRPqOK2XgmhST/tBgX/zQWwXFIAfTrn+XnV1DlhKeTIrT1Bum3
04/X0+MAk7j6f/u8fQISmE8nBcfx1BoJIE/68A56pZgpk1cx8XXWoz2o93T3
lQ/qLKtt2bb4gbJBcgECC+TlNGdTMBOzByQGw4C3eYb3OHmBCbSD7CyK0Fju
zzmDx+G6oZ+wlB8OU1IaEH7QMy3/lDvkAZuQTMdCTnVN49YBu8CY7zIOsxxM
rKKkEcpULTyo2Azjwsl5SgeffvngZvJiqQ9hDd51OUrmFcVFuUI/VFaEACs/
PPoYLJTbLc4JB47M2NT1D2/x5VkMEZoXTwGVi6WNJXqSnbR8JPg3L7e1YqNr
PTMrqZB9zkjFLDfWR+086JoXvbIh8CdyyZo0y06MIrrbbAZX+a4a6opzC23p
ZoUZ/QpdqH1kuFs92k5xmkb0MNoiBHKhnOBt7Wa/qkt99cI/EkpiUWBj6nwg
VdhWMADVuSEEjP+GOmYDhlLmuPpVYqSmbzOsK2KgdgM/MgsTiMOojyNPibBn
9u8Sk2vv8E1AlKqhKSZzB2i/S0e70XhTGiJMDgKUZydooN6py6Wepa4YRXoD
PTlBu7+YSpngxXn0isX+XLtGJj2IhLQtuz+IUtKQ1L4dqXZ1EgIfuZsPGeee
gYNDoue5K7kjcuDjzKgzA0GtUvlATmEbKTyFcgL1/eZtnWC+DJYyyvrlX44a
yE6LNNyi2utuhMng1BXuLmO3IVTKHJ/A4FYs4eATUfaTNTBe/KnCu3i1raGR
WqpllWJuogXTkKLneGW6An7Vnd9r8EBjO7kQrPkvVn0Ae5wZezNw2G3OY9IB
hBZCUt5gK8xNYoRXGoNM2JjE2aesIMJ379oS4R/4Un6IV1ezjwczoAth9duZ
r6t3FUkqx7TjJcnuuPouxTDUZ2OlZQBHL+a0Wle7Br/hicEpYyBD5wMA3dCf
FtGFht3D+S2s3RLQheQ879CJvJFcFsjqdMeaZKHUnb1kW1zjZmuE4Eg46TGe
l5MZPAg2JWb2ZO5fYPPW83bCb7Jz4kmBekQQawUvZQi/rKOlkC/mKwLAUH3T
1VypBNnSRC0pF4vqBF5ELdxrOHDicWeFNWC/GC7veEsuujssHhJJdKxQipIg
WyCpkahtILOhsLmRv+Hd+S8Q9uBrtpvX9qsheoQDELvJK5WR9ItHlTTuevtn
0YymUuXfud4adUAKKPrK/iC52PfhXdHhX7SDAIoSWXK4iV0wGQjFy5f3Z099
1/02qJCuMM5304s414kEntRfCLhZ/+gEj7mWa6CkpBMBCFQZx6EolA9AI77g
uTnjE9ozf7/lg/Gs/yVTDzMb1hNr/n2TMYfvwFdSlTv05l28yQlUsl/MQ0ua
K80cjxr7DbDHpbM9QWEyDSrt8PpqJbTje8N8YnywcV12Nehu0zkG3Zsx8VEg
EcXrNR9arXByMzldj19+WgHTkbcUhjQm54M+8Px5/l0bDmmJbbKK5IvrNqXX
keZd99txfwqq0xYK2PdOS5ejzLOesF5zqCxYHbVgZ1Gz5nYOwQNfCHmb065V
2RzYbaapOJIaUJK5/Wa5tyo9h+S/Ykdy6usvkFH5wDJ0ZLIwxl1cX3uS5kaX
E5NYhe4M/oiO0sFMQ3G5ItkQNr1zTHtKCBA5rZD/fLreWFORO6qxFfhrJ9Wi
sgFTo7H+jsMTBE1Gh4a571at3JydpO7ZGwxV4/jhewXW97O+Qj+fepsjLxSk
ymvRV7nGYHlAE8qnxWmFWoeYoQmbWQW7KUzm+0r8nc2YQWq9Z8ia1bAizMQP
cdsAFETOYupTfi81jHI0TZzj8fA005G68o1lMjXHdKbhKyyHC5x5+Lyp8jEi
m5ccWOGzmMMg6Aenx1mkukzgRdl/H+WKtQ0HaS/rBkmAniNPTIQtBj0lQn8B
JEZ9TSU1kiJFCet+p9Qs8pFwYuoraltBmNYFZhx/0ejQPgGEqlxcZIfiCLrs
BN+PfwJSKcsD1hAoFyOGdLNaMoZAAcxzi9cyqwKotW5li6X8KXrg4jTFt8Qk
ZGFvof3sSfIqUF2SP23gmrIuTRHzRc4pwTDWpdSOXjeWo+XjTVoa92LI2Gtv
uoXNDNdehaiflJ+8Bc91j+g3LbK0jl+E0SRU6gDZX0v8MI6QtSH8OJDHqFZN
gFrW26W3LP1HC8oPqYMINv3CpOJPPlnJiCofB91uBSrlMry42RXs9tEAYnEY
a451HPB/vlPOtBuUmN3eEsXy1Op2et5xemo+6Kga1pek0EzmJZ3Tjg+qrPEp
IxX4vIQD9sxWodaGZtf6cRRaGs9i3upjEn5pN5krFdYI25cEtd/ofrseZqw2
vONuk+4wFltJNiFCTkvsF9Mz9QVJale2wv8X/G2vu6hsApplPMx3p4jYFuht
0mLHWa3noyuCIwd5HexP/XPHEsivMupnee6McYVx0WgjFCvAz1Bvyc3s+rbi
Wm8iwv/Kg86DbR+ogItUdqVuX+SkCkX3xgXtsoYk8pji9AFpgJbGHtAlZgD2
qdRoomUPFo1F8lKfGyZzgEYOKq7Bvof11ZVHG5PIoIUcpHtFJFN7UNkEA+2L
mVq1BLpjS4fG6P+67OShXpcBnXeenogH7b8h6vUCeCfUapmsS6VMj4VdpakW
xEWcKYNnIwnjvM1O51Z3JZrUILXmo5yt76OlQsZGDt+5yOhZQATU4dACYQhK
xEsruwpVBiiSmKHnLBUA2flYwG7acZmrAGhkpm/6BuJ/qGO7PMbyCBv0o1T1
HK7hiKHzj8k6cg4Si66NxhanwaZ4RaIo/vbwp9KDswRXb1p7BX6DEVKsYLsH
g/EZGr36EgsPt9bamUT6pzgUcD7DRMkzNisveYt+jkFIBIUs1aBdgk8AkvAO
RQ/vvD1gU0du5GWDqTOpxw8PJXMzXMHBoTH7oI6G4QTxt/44rcCTPl7Vnn3d
aFcqzuq9iZAaQwx3QEY8GyDE/LrLCWZMUJKikkAMMVprV8Z5SzPArdUstTg4
C3+VWwfAW6aYRsmjIyOfD2J3alop5RkPom+hlBTZ8YIr3vLBcu98xpLuxBu3
kJjAw4ZHk5LOkiQdAqQqrnZR4YexYpdRs0/s195+tuaxHK7AWA0FoZfW4qJM
RKDKUoQj7SFwH9Va76CMjJK5QQp5mCgI0Ha5/S/PTgwWYZhsKn99e1+d1V+s
GhCNmSY43eODB6wH4EY1T1NAUbLI3wVTaZ+lHaqH8xO7+ItAA4dGi/nyLZv0
R6ZV9CUvfawOfFf6wkMZG9hhXAtfaOC+arbxV03ixWA+e/r5nftk3zFwG11i
3wDLq4pp8HCZJ/wgCjfZDZSGPPScKxsOpJlPcLWZwsKan8XM5Ri2J2gsHGtZ
phZkUaLm5GlcjTOCuPk2y+7lWQ452j6U8Af9Z7RtgeJT05I6QK+jasBXNt+e
/zd0EU5aFy9oQW5w8KpIOL88/FWnYR17HQccCunC0+ZjdbUG+5yUhLkL1/Go
3nf5K63QZUbhcKA8tJiEGtpfB2qI/FQ/N85Ejphgjo9EBiCBKYS0MqNczHyW
gMQwm6Sc2XD2yMs7+0QG6+HIAKZfYuUK1METat+xKD5ZWTAaUVA/mdigvjYo
/pVYFOfj5HuL0bNJff5zPKv6l77bceAtZngIFOFWpbakfqYb9b1s9NpmYrtC
m1gjK/pH4aimDKCNlA1dzmFX4avXc2wzhI7hepDoQV6LFc2d7PRdHD06devE
m3liNfo/wwRoPg7HopX/yfaPEkC6X8/l2hhf8aB+dPkYvjbnX3X7OPk5m2NF
EDuMyUfYPTBH8vsBh8almVDFFFtAutipa2utI2iJQd1cJF+LPHDcahVl+VvG
0r4TO6q8egfLCfqyQTqk90eriY5+Lf7hph1aFbTV1NFoIWLrslyi9fvp7H0R
Bu/TE5/AZGjz86MZyAl+j0cAlt4Sg1P1wBofUvI1QfRBQB6koP3ryHYkkyGm
FwybdQmEobBqgH76wG4tB+30Qq4PpJVPXIFlWg+CST2EDHTAzpmuQAsKemTh
TRzADCrCH/4+ROerclT/9KOdH/cDlRR69XdyOqi2f5alp1AildInrgG1cKhE
1dTXHDKRpLFo1g1z8vh6TqajKHFrc0PCfK1jW/TgKaBzdzk5Av1KUpayIJef
c1nCC9fxq8pcEPUQT9B0wnGyUS7xe6mzC/u3UppksSP1Vxk7zJA0emV1XqHg
cMHnPQ4yiqohYoHjQ17yMUzJuRazrjCbUeReaoLA680txWlz7t6CTQAztwr2
RzvQ0OV2soboeDSqVRHGlj1OXoySwBJEJ72JUrXxtQApDC5UTP75hGTTVgIn
ZUVQsFrCyt9QDZ4JZXHJ2f1fgR/QJkG1UnvVc769S7XSo01dX7/C7xxFhaab
WRdJ3Mm3mRFf27hpWJsDyIXs3SwyjKEIA7Wdswy/uHyJuIfItfqaJv2z/71J
Sypo0SM8bKphu/hUMA/LddOt5Mpgwn1P1n9yReNu7pMat2bOnlFIZdZUu20p
jKljT9/XXvkl6fAnKjUiRCuUzvslWeB3RUoSo1yycAYQYHR0R0iBN205m3NS
o1JVT/oNUP9QmJ067bbHnv7SKKA4V0dMYYtoygnTxUIYkp1LeA/vG2hVH+ZI
ZzzNmCW9MM+3wilub/WIBECMIsJ2ELIMayTDnM8fTMOySXxYd9NxV9b/G4UC
K4oiUKBQwmWt/taSbL4SbEgarIiuDbGwEelFsTMSxSMH2Jtczxs4f3poD767
3mbqUU2xIaUyEV+s+C8Lf6QDQVyF9rOgLUlYMwWq1HOzaclUd0zv62RUF6SE
j4ACUDZHT/HvrjZch2HuFfIt1EGbHwRTK88LC49LyUhvTZOwu7wTa5Ge7RLO
ICwyke9mt6TUgbly+unrF+XxU5K6qH9EoYyVlUNzZ4V9FNNcPTZlzqhnHNIG
PPHieBpCgacnIwtdGWlwqiDiDdrjjpA4/TCU18RnK993IG7YIy/O1JoWKUsr
Tue9uyFpIosmQYy4vJyKWU1uaXR4/LlT1rtcO61yYHW+QMWF/rtMvF39hASS
2KsiIUCLxLz/erp0da2mKPQPh5etU/Z3C7cV1dExnxtJLngG7T1Yv0qiQ/QP
Bz5I898EjG47yy1/UMmqWxer796MaRt2U0XHiwijCENyEuORUJMt0yWVxCQY
g8R7cb29/4AwHecHWHdw0OpZ62tkKUQVmjzlfb/llA+OlKg4Qe6sjnz0MDvs
fzEyzYIJ9kRr6zA6Kd+TJjWcEw9WKbWtrz+oHtNkkh/6M0NvZqw9ZmQXPJOX
GPH/ic7/JQHV2ZfZCHd+/cgU4RsDFL1T0zbfXrb/a71zzjFdG1JiSa4WvV+x
XRyM7Km/xmCcm4G+nVuxqif68JYrxbNpnoRrA2Y4D40FoefTenLeyZc7KH9B
U5S5wUZIUxKYvIK8eAhWzr5/jXfL213NNKspkOWSa/0kv2ZtuPEf3GirqrYC
jlDd4MmQweNYihy2wcL3n1BZnU2PY/VRAIZozpVEtYbZG2cBz6+yCW1BHOqH
sKlEvru1YWsJWR2imG/czIFkM70IxTxZWZgDmwBKrhr0NmTEY9mNKGrNMHVm
PKJ+s6VybwLveMf69EyCRZRu0qDtvP7yXeWwLDATfJcm+AeYMHq5dKuNR2u+
X/DgP7oKP1tMti6T2eG+lxKMfNYRHJziMExcnRtdrnddtmagEZWCbtaFtaRC
mVVt5yjl+jC8IRCPtmo+YRbmUd9owli7/bS1o5CEmhLMSo1BidHt+u2M392R
NwtOxHZODuOT8dK3W7iSWCG0sBo1Wy+6KPTcR1DAbetg205+2Tkj63VFH1qC
49ByXXOK1VJG0C1t6I++vvcwUrZ1uzUq5vB5NcFTJ7YYLolLkHuMJ1yUL8TH
cv4jz488xxVC2kZgkxH1nEtmP3yFZ4ZjTyiE5Hjr082YwqeHyqOBUBOOPtaj
48dOUxDCQKPJoWTTS4uiCkJk0pu/BOy5qtlGPvR57Er6c4/7Wgf1r6yo+5pv
GuH8e92QBgWOGC+FXK+lQ/8xPPDlPG+9mkZhMYI57U2ZwdlFxOQB6IdzNVq/
5r3IBIiHSn2+WJJpkMVjY0D+NDC+mvqT8Om3IHgmnVwvMf336wP3W9AUBdHi
IcqXp+3krruiW8dJfTcL0O1jein74am7xRsGWux4Rdavv2HyIy/bvfmssNJX
sLYUY+rwd/AGtbTiA/0wOcLMY5uJfIYD7Uw4ZM78M6GOLbN/R5ZDTz89uRYP
IUrmxdDN/iykJIzlsdCNEX7WnC6IWlFVbMBkYLN+GrP2wR/TpdiwaUoBJ4MS
Q0tQIt6x1uyLUrGFp01szlmuN+vs3DOMYblweeg3l9wE8mVS5xw+A3eIVuZR
uCEHanJ1jg6NOEeEvQXmuVlODbpdz8OFSwt065jFcu6WUv763TAQTL9j76pQ
q9wtmuxQWAJ9p5KNqfAqINRUWMwAoEMyld7ZZhwaTdIEJb/2kIZCnopml0it
hBPXsL1PMxC4a5sJEyEv0NXLLXFWx6xakUv9Lms4Sk4LkCDlByoOkfdHhhNu
QPLjyMDDmgPljmDpq3BTlk8HDZ5/R1QcEGvVQbH5FolWQjNfyK9epznfPo0C
qttOXu9dV27DFc77/xs5fMP/ji+LAyM29h0yizvjkBSxVJruRHsJkQnXCix+
YkYkLsbf+XoR5fKPpB29dLgp0TKfvq8VFlarYmtKzdgSZAI+/nczsUCZexZI
WLibXhwp9dxiVh6NxD2nfNjDU3Y8sX0qEJ8gZOKHFtJQi3SQUyEpWEbonAIU
Z9Zfd4SPs12PThaI6EDVlCu7MiATm8RWMSZwPFvNwlArG2/hsmLCQNfAY5Ps
VfWnbGzd0hnZQLy8U2F086/itzafTST+KRY7jI7CueRWfabutXeZaN26u3D6
nlOeBv4Whe6syfTZbzTQ5RhO+WQ/YYvZWh8L73Cv0EQXBW0Ta9snO4kGGzZW
sIcA6d97j9Sh8eBwKem+BIiOptMZeN9myDiivE6SKLpB/mncX/ktPe99uiTR
DxydKLQX30UjpXiVPRHETp1b9KnDH9H/p21K5hge06hqMMu+09aMq5gaqf61
lXhYoRpN37jF8rJLefKnVBYJzBYVNHsgTilKNIyohmimiP3Dr/vjD7cSzj5j
+WiEaVfDbLMl0CRj/sfQLyTFV/9SVEzduT9JXIaPOGCjE8E5hBf2SLE893S8
MSj1qsd8CY2Q32SJgqyxCty7fqFId74zMrtYXHghKamNA3w74ZlREnK9hEtz
eiDWdufj1cScJ1mDyfWYIaqg/7b66nJOTx35MFNooov4YBgN9VQYP9UrPUfX
8rHnwP/hOwysMYqiiHi1gVq06bCLRenOO2d6ctAe5F8GRNR+MckOoN6bGAG2
GFn9SftWJi/i/MYc7jdY2qsj5BOTI2W+dOvRBZ9eTqyFWM51hs3dC9UlLqJs
IArawqhCIK4nOW6SAzju0LueGG9FIZs3W8Z1/+Eyr5yRFOGM9xTtjBbNKGQv
YaxfyoPaJdK3v5hkeoUDgEU7Y19lXbo24c4dwbb0oVCzSZzLt+LBy6t3RFNH
o0FPcmBwnWWGBDlHD9F7amz2bHdo4DlNIaZJ7W7sBGOzDLCPKe+411ef19ni
1Y3rEfvWQk1g0L1e2TF7jowOieRzz8Inb4tkWJHXCC4E3Ods/xsT+kjGTaL6
4kZFddUm+D9tTy8YqyVWngVEkFd7Cj/gUz1g9VzZj9HytZ7jzJ5UyBn6arcB
Cj/PmmMXyPq7IFtIEaxmTh4moovzG0AyH9TFikTB4lMF0PRy/SN87VxPWZ8c
Hczrwu70rUtRITLHOsQ/xYnKB+YAP6+uIFDpkVHPesg614nwMKAnZYLbn5So
RlQlv/MiVWhnuQKSr9hTUCJXmD16AjClQ5i8+bPPg/ykpOtZl371PghXpD1G
MMHx64kyImWCk0SxN4bhqX5QNyMdW82DhcovyCLUczG7tzveiJggBDMIQz0u
4fuLaTB/GRw3m0fSsOeU5Q/1ymZjq6qduSgxp8HaO2Ud63nLylQ/wT0pEX9o
9cPdqQ/OfiJ0Fw4X3Tbcs7GzcPATr7Cm+BxsxdX00lI6SLP8CE9ZFUITCwiv
DrTS+8X490wD/PAM5b54MPYU5h0MsX6FVFR/uFqMHBvPyG4t4Sui54RY8c5X
R0eqCd8i+S7g6dYosDKvJ8u+BHQQRsrH7Ok+TWSeX9jE4Ko3BKkiFJRv4GKi
rmhozPntUpvAOEniagfjucQk6j6t+xwRp689gdE5WQ7xkJVVAVWovuLtlMRV
vftPl4ei1AqhWtqdW4+J3T+jwrn7BRf1C1ryouFhcUcHbptrdHFTx0sBa/k7
Q5VsFjKv9Kp7gtxzJYTAN6cJEYqyxm+AeZ77cNJLbsaBio0Vf3UIzap/63pV
4WHV+qWh06UF4tu3G87ihIflCtv1/VCJTwf4lnqD3pbbvHnxibXFNdmXB/mV
H9lPCtkP2COZPvhjIZQHY0uAPBNoDIB6t8pT8QZk3A5q0FrYQhXGQhbymSEu
YbKaViLn6OdwU8EPR3qGhZevTKX9TEHOq/cAiw9G2G8gsKtX3hVmU/KFG/Uz
EiQGL3lC08yXnRb+72Bj5Ahpj1LPzcC2CEmncKZswylOiuUKU2bRjwg5T08j
vL+VXqx5FiWjIoP9eLBCSa+JdyyyT2kyuBdURI6W11HoGRN8ffnIrGVZSajQ
/cm9QhxcDx7XT7n5POeqJu9B/EP/hkkciHF5mTR981HXE7gzJdcvKEsyXrNb
udQ8g4MdPRjatXuNdZiqwraG/sKlEPGuoZQ6mZt8iJvXX/EYHkPrESyeUwis
M6TBF/9k+8+6hwMIdOyfrdvBILOmtMuRwAMCi0zZmkhZcWzQ6KzTL5BWszWQ
x/uroQILUL35w++RsVB+nfupCIzQf1dU7K3nD6dyHpvti6hwSXZucfcMPtGd
0fZDoKCyTFEC/YY2+YeuhuzKvUH2rI9i6n0+75WzcJqDpJbSHJdDvFyt4MaN
aYtzZxSwWCHyDW8KDmapHQRNZsmxxkkpBKYsjD58nZQ6gOOVzxuEOyXdNsSC
T7ym3zrCeMSNd2LLAIGWg0/PyhZnPMiZ4zgpEKD4fKe5FRZAcW2QG1p6lWRk
SQwkFr8hNcR2CFqJhvzRwmcup8m/nGs/VAFPM8lDWuC4BtCqKk1wwOb308cX
bxiyGT88grb6KzUV6gMyPH0uuPyO/kUUC8yTT469CAmqE7rUEXah4teh3SG6
/KWKy320prcEqCnmit7O+xukaXHtlFmUaQb0Fu8troL51dipz00AdGmrwC9X
wzK2IuFJXyZb9Lw78S7P1+a+7EUFCjQvhxEZJwSRztCPK7TqJIR2jaCArV45
qI2pp6KHKy+TOwro8+uoydJDkQyjC/RGGnKYZMW8L7DJKQ1Nz1eSIrau39WN
rqhkebaHzg6vGrfht4rTHlbV3XA0bSmaIOi7TnJWKmDzqlgK5mdZaHSPRciX
cY6XkC+0pZlGl34Ng3kOZHk2DNW6gFDdkTw5gYfDu+6EPmxpyxZiMykjdkeO
+zIK94x4Mm+YFTI21LlmmE8jj4F3lcoYv4YD64nmNizwEPmic7/hKi3qKBbp
ewJFs3zqgZdzHFiGYU2/8R51Vi/svOQSm50T2mTGdn2DyXtNBgX7ixpeFEzV
LFv3GvgC8+1UOYbJfFFwhvHw2zsdsRaymTZ7ICmTzsq7rwZA1I4mRXAZ8riC
TBhgyWFyMCs5veJrvZhbRQUdQWCtitAngxvKRhgLGu9JB2D86Ovp2V3E31/8
N5Y22FYLVyhWms48l0qgdAO3vVyCqKpnYK86wYsMnGx4jT7+TNln/3NxbLb1
kfpvhFDb+91/vRWQ+YPwfGlUIaqhNGiyzQ/lZh6yHKnkNXsD9TXeN6ZL0NHg
d92zi3kPbc+G8G/SrfFw69wRtPu6nMKO1DnEB1Wm7ELCX5vVZWcTbb5Gsm3f
ltXF5AWRWEjEcucrIigg65QBklGfkEchtLOFNa0hDZMhn7V6X/NM1tCpAauo
3PwZy0uSAgNZ04wbHvx3ILXvIjOAnZ352WbRfcbCq/Tt1lBAdlCZZ4kpOawj
fG0lUkGUmZHkJT8rfUqee2WFfcF26B3kagUlmZwNts/e7DWtfbmCqyCNTi3n
OFyn09ar1DtfOw9vOVeR0yVvAJLbwt4Sirc0XYlO9MnzViHpQGFh+271kF16
9JL3RobVkiVfxuWOXAkTTI5sYajhPz4ST/fo2B6DkWWrywApSVJzc0e9MkA7
4EN5k5LEgU/4JljFFRYoXnIXC++ruO0iVth05vgZMVSyOx2HcRKhBgHWrjUC
nSlbslpydROmxgdzUKJHQmZdFwSh4VwohucVF9solfyl7RVgSyDDFirjZkbc
o2YpCSq9QpIRfswY6mB8TpJVvmtEbY5tC2F7ZMCc9D5Z4rjIy9hK1CzmCzvF
zN0fbRvA5T0xPay0yMwYfhagT8cQXJDLChtkd8/FOIHbiqkcaDEpSrkef3h5
nCjV8Q3Xq4pj9ESoxUAOnSRBXsn02AL1dLVxX/fDRraKNxWsgsMoPMnHjF7H
sdEPeEmCbvq093aZGN2gxb+rUcHf9f8ajahJmORl1Urag8R0TrGEIdirDy6U
ovpZyAXWcoWdPtxENyMWIG4ZBQbqW1AAiOPrvOUQhgVI/5F46QY1AS6ZwMCd
C07q0Oh8LJkhB3iCXLEUYaaOurrp3MpzhfSkDzz2VhZ43x+3U2z2K/WiX0sA
rDQGZW8AgxwLXHQ2jGXUAcUZECuVvPwM3175evRPmYzI7Cro1Ga/fuzz3Yty
8uMHrS3OLBHw6oqebR4XKrz0XgrbLoOssEkpM011EnFx2UKJcTXvSfm+rOr7
uLG/Pr9Ci3HATzA/UXOqA/gnwgf8L6nf4etqY3JSq+wWk8oKVKWuKOvIyHq6
x3IZ7UdqS21kvZPJONASaf+cbG9BHhUYEWc4FNS2kUf7OfiRb7QjHpkFc0O6
fHhgla93hyUlZOXy4/G+j+N2/R7N02ivsg4v/Oz0aQNmzuqoMklVJTK19XTp
Ewq/oUGK+vH6nRK0TPIcU3xq3uJMtIWjo/ap5mJftLDdL/myID80buAPCKXY
JCPLOAtb5co3npdczKe8Gv/WVibS5vdTG7SxJJtG4ChpN2IMrJl/3re1018s
V5PSiLWh3FkNGMGsCqn6M2k+rDvUj8doDfH005sTjWmfulokinm+2OKZzigL
h3xj0lRbHISn62cd17oHVD5UgSVzl+Osb3Vbwyo5KdLHMILNWyCtQLOdpF7q
LDhT0MqTr+Vs4D8awcA8c7OxN0ySjYQEhxYlT3nYRBILDBQPcvKD8YuqWSkI
XlQW1jfrxnE2IGJWlUr3rlOBnD3NcxmM7Ku/bxoVu8WJmz+9oul9Djc0NHtV
VctjmVbOEQ+pPhspZ/rlI/NHeZsfeYeE0L+SxQ7ZzbUOM/SnxIZwgdjjgXAC
W28AKMJNxXLj1tOhrpV8z/yAmq47Zk7f7VnsBH47OJa8SzrqgGTSQMiV6iIx
DXZLP95DVOAVruvrPDXv39vb3S10x9ziH4k6c5zFLCYd1fOf/veLoya9Rz8w
W/VlM/R4K4UuGrChVcIaGbLCPUwbVEN82Z9AkBpSklchXpi0K/24w4Vuo20a
EpFnqDjZs55A2TL2vOhu0cKKXtReeriOu2wbfuAxhX7QilkC7skX1YBE+6A0
BL/N+V2OcpR96Fal3Xn+4lZUBrtDRK+ob0B4zDFgbjPcuuz8zimACrqaqfof
llttL/mrybQjSLfdN7M03ctADc+Qwr7hA6UaESm4SfjEF1P829z3kDCQX8il
dFqCbKP1c1btZH2OMJZm3jFu3ux7suO6kxel4n0G1CgMCfTzfHXe+VYTyQEF
TCxnFVEmLCRTn9mgl+TuUtX7OVG3Q59s/h/TmBh+8j1WfjEEq4JRazUKuDPs
KvsqnwYmGZU1Fn9deXJDWGnIGFzCb80oepv1SQIM3ywqReSjxYls8HkpN4Rh
nRLb25APuvntST4s4eQW86ai1d2wdndTAY5wa50yLwSj+SffFDrptqu1FrY1
I8Is0IVLeNxl31fZ8hj4FEEG9tXMJF9rzWI477R+SEaqfBuTl3ub/q8/MHML
9OY/Zu2zNSzzxuS6A/S1DNH5iOkpSTXOPs/5FY7MmEbJo6/TpkzzK5OGpzZ9
QyKMKShIycBHVbwQJQgTnCc2s2Kf9DIlLShmekFp7YQpTCvTeLFkNsmx5UPc
1cAA7f+zJ7MiB2ghinvmwwiRcadzSDD1ktfgPZ1n6AiVvPAq9WFRgU7tO7r1
fgjL6/wV18v0nZJTfisLWAV5ENemvrEHv4Es5aVgSHKpGWvKNuld/eN71ES7
JswTpiVxEjZqsSINPI26UPKLKld6nID7ReofgT6/z5IwmQ6+EpVfq2cn5Ybf
n7UEBBvHMuFsaxdtji+uPzk7jvbUV3x0yXRvC99tVyL7LtNlmTR1jVNY0abh
CRUx1s09Vj7q7Hin0mAfBCVUm72bIlMuqFg33v/i3s7/36e9Tn8d2Ci2bbeE
PabVjFDsoE9FpGF40pbjObigBblG6UHrquU3T1Z3qJ5Uh3eiUGsAE4nwTtC6
p5mpAw/S6fPeP2w660s2jww47Ntk6as7mbMS6ixkcKmPjkoS6LYo3zaGVNn5
cJha1yfO/ihcG61j+xe4f0dIdpjuSFrNDcRlLSyPcuZu21GPmJsa7OP6X1fM
ivwc3Y9q8ySgI7MQrG5tAVstlGLUw4+I/IqZMiCY4UA27PuFiTz5DaurBjiD
iTC4kNqaKrna9tdMuKCTJUrozbSmKRPNIPaMzpIVrOf/FZkvcHheVjAsttGY
4F4CMR+tkOVFzLSwE7JAHVn7aQs2wRWPwpkcpRvehljNuJlOMpsbhn4ytSRd
Wr499XuCKrLrVFq8Rs6EsQBjUnunhaSoR/Is2lG70rTp7SOkpPGKPQfvns+S
6KtPbP1EriKCu7wXvWFhtCw3aiNIVdLVuQUCUPusNaEEKtuJf2IKgRN9Oa0W
5DnV6ps4l9G5TkFgAvyd2ZRxTWwGntIK3O02dpiPzFkTKXHaJR2v4q/yHdtm
E1TbLmWwgMzMpLz0O/HRdj5zVlau/x8a1t+F5jDNWnckbQgODHc22LmD12Rd
1ojiMdowLMVyHHeHv6YN4C9HT7DCEdGyMWU3VoZyAWREuQDLTpxRVZdu9kbi
Xc7jEJJ6KhfSIiEd6ZqAecg2notHt0/nwcKUIOJRdLYNEnqKFn+kY8BR4MVp
tAvMHrSOlYDQzT4Xkwfy/bk/eyxSXw8ekzZaJ0pKlAU2L2OReL9K5h12jaeA
eNo0mVMm9WwFVy6L+Lg5+B4kWXDtaQHyy8MKyzfKZcXOQZzFBOWSbtQTPdsy
/Qiz5jO//HvNFfKkvJHrSuVTJE6wX11r+9KsVqyOzaECaK+L310yA3SMNX1m
ngtuDFQJ0Z3HoEIET1Y01LnL7Y+AvgH9cAM666NMTLxJyS1DeFk1+7FY9SAp
xYgzIYsJWdL7nmEe38jAydmlSaPAOfVV/yyXw25fh0UvlmVCvUgXeZDTtBAS
1kPlXrht0UOqafv5MMlLhF7fPLhAb0B4MO77CQ8ssYiS9IrY7qLNFFRIAcJT
1q//UlPjpZ1OcXMaMv7LIjy9IeZ2i3zjRaDZElnSmO5/hSaSrrYsN1C1Sz/P
jQMySLAunPZnQBL0xgN17atkT0hZw9QmZA7K6ZW/EsjsOUfRjt7WZ8A6Kx2t
LsKCyeE2wNXOftyZPs6UxOV4plQnf2OYgs74W9GodnjNWcdGwP+5dNvcn44h
ra6kI0njNV+fveCuy2ZWCdwkC3haax3cARiT2+YWCs7bLx+5TWK3369GIpmN
NfCkY9kV45fXA+z+uiCk6nBFPr78kZ7Gjz0vaIBmrelH/7W73auQ2wcNm7o8
b5ROEw4xAv2XB4B62GwLUz43rD8imFFgLhq+74ox6bRUF4CmhokI7z/qxBiu
Urosvdsl9/uOJKa+nqfDMzPO72t/0xFRGlMdjA13xJlEW08tOgUheEkAD6NQ
0ymGEDCtJzMti3GhEbjEsxYkdYlf9ss39DG7jYsN/CmIN+AwGs7fb19cPngp
iq0xuuM76U1ksLGSe+uzFCswgmtKCLObT6QvLQZJiKnWQa24A7N08Gh+Yh6y
BwGWxOXcSrKoV7BI/pVtoux+cjuGRBfxkgX8kdrg3s3geQFSBXGLv/CWGE5E
e2XkOLT0h2XxdQ3jb/wEKbsciVMut+CBR7kRli0uZh+DluGKW7ilRst+m5K3
ZxPoFNhrNMD8dRQoKmbcs+Vc3EXIhOBeRWJ756QPqriusS1UXf55lKy4UHOy
I78hfUGW65W+zdcr6JP1qYUMbVbr5hFbOUbCWHmTFIvi8fc9/W0RPwBXRQ/N
EShgkKDn7YikznzkvAm5LohIvV80vTxKWdV7/oXwkADsmDK24W+VyD3+LNZp
izv+1nsFCOZS8gV2xQEQGRScVZGiOF9/eH32sdcnj+4oSPH/vwACw464g619
l9qCVa/mJJ28g08pQ8iYBUBHRPbNkpLx+H1K8vXvoW7Khun36ImQ3fbGHcW1
B0xwhFTtGmvUQsjof2mxnROZ7a1Nz7V+Yhtyda4VF7SrsxRYaIOgK5R1KWEj
brTcNJx27bCK/uqKiuoz2gmO5ECRJKfzxygEFUUopIalchr2dwPTX4C+leqI
9lUlBsQDEH+yN/UNfN+BY59kPJQmaJ/ooCRsZXBx+VLU6szQhGlN79hQDywW
/gq9/y8y76YqOI1kv4Yrzxz3mGKKW6QUqfoV751ThnmMrma7bHsMQk2qsq2b
aAkEbobYJr35P3/NlxHSuHr/w7aykYDzuopzsJ/dDTr+LwK6/IViBqkZ9Fc3
XCrKhss48vLBnGDh8AvrfkxtoNEBwX/Csh+1jzRhnbhQ5Jp4QhwOxXHnotKN
CLIki3MaWQ4HH057KLUZlRj9GuChYMjZbRaKIFKYi5Hpbx18uht5RLucpetq
OYQQrMafVFEcFXnPgm/+1pAvqMnjC5todBiRHODpk0XmMbQasF+03vWNoFWE
0RSmKenh1Py/UjN7fBqgglS7+DJJ/6BVdU/z7mUuF94zBhtC7FwcWcyEwmV3
5uxaMIseZSuo4Iy6qHpRRxBKqnQVRtROWGNpKFlN3gCdaNMA5Uf5egkyETyi
KKhfpMLixj/dmGb5Xx5Dxc56RTSncx7OgG8jz32kIYHA9cQzVkqJ18oAdCm3
KvD7HdnFzJMr+sH+AtSFqQxu5vYDWat74Zys9eCagcWFGObJR3WAJWFSGAzl
Ra9kQLjYopqihg+xAngtg9oZu6cyDhYmGEWiBvCYdagfrMOwnGZNnKEZdnaL
ApmVbyNyU6muJuCYUfU1bKtOP1I2lVRZTE3VoiNyaI5kZKKLk2sGcoWqPb4z
IgDf4952kIyPNiHlDHzI7qeYBLdhncBapx3TE7lekejTB776G7U6PQ8V+rAq
8JWfnk4h449DwD8IkCzwyFJ+vfrXw6YCoVG3mt4J3HvxHPzfVV5R/3qjlAI5
gh7B4IgNtjxEIR8TDE5dHDJjtYTkC+dGFwOUT4nwczjYPGh17eyKBqk6nRWV
vHQtBorWTXt+3Pg3Frn2BPVkERgceC0VxNv3KtySJr0jmiXaGpOqANvDFYp+
odCSt5F5kna2DMbKzJfcHqNrRjKiKO/4fppxPZWWhbbQeHBzs2OkQkkN5E51
mlT6q7xmF1FALcnkvmvIKrIMuub5Weg4y8vOiCZSN7ZhpgANHf3qrOJjkrN/
frUy6SpjKwwFUGGOh5u2RK/9ieQLLBSn+CUAil5IJziJXrl9Tda9ShVqHFdJ
TN74Taas8jkZRNrQqaoqzgjQUAitO9x9i9YWn/3+CfTZodAt54tZHGtlEmbE
c6RueP/38B9jcJI6f2hQMBMNOD9V5mSz9u1nUmWJiVhnkF2c+NoL9IEYfq+Z
tSjo7UurdKTpfcTNBYBVSdWzX0QPJuDKxn0cSzsvR0U5c0iHTbOyKUmLdSx4
aF3Xh5uDBQlkXqKPjjSRjenm3i0aQwb9zu51GQI1KXeuWzLZRIwj9zJEtpMa
2M9ArzG1NXwjJAXwH5dwM3TQyn9zvVYlT5IvpOCo9oEycYu38ekhsle20N+e
wLac5J8ownl1usm3f8/XMSndFseiCuXxOq9T/jWD419WyixazDTpiPBgMk7p
ASqIFIUXgMtWtvY90gLSEMI8TpFf5JxGxWn9RmKou6mtd0PyGxK4gUmX1Y4/
dakzbIplc13L6uiH2PlkeL0KWJJ4zALtctE2qhfTHlOWdoYVbJ8hbJFpeD1c
LUGofVgtvZ5KC57NxCFauSKeaSTAXPBuMnGHwAOpoHaPC8eaksGRkawEov4e
v9Y32EtSgzmWoJTaoaKEJeydUYNQrW9RsjkPO6n/loDhKfE8xjRcbH8Q9E8K
wZZDpAXiukzxjwXXdclYLHUVl9l/bOGMd9E3tQsMdLyQxEI7xsnssMfQ0QNv
wIPnIhJp30UxqB5ChRxkGlfbLHljrRTXwt15O6u11gZ7euv85P8bzFsIGhlr
ZggYYG5LMcT+gAMofljDwWz2H1j0vPtfKdbys+Rh+XcFmNSvInbstMTxA463
PX5K0Uq5nZDkBINiq88/hOzDl9zRLNN3RIBPaAl1M/Ez62ULzQ7DgjoVIF36
/aDysX32aXosycuZQdUKuxyDATwMD07U4pJdLgLO/qGkNFfDUtP9PvD4Zx73
DjXRYDHM5ezQh0GVTsz8qn/3bEU5KqRIC992BQZBuae47CzXxnGUMa7OCKjh
Wu9N3WYRxrxG6poVzbQR5PUED6jCt0XXlOat8xSB76AfjVSmCUHds1lSbC0g
IccI4TqLivNaOUlqbDqRgNABPFnLfDMH/kDTyZ6WsTA6qJe/pR0Ffg++bGp2
9W+AwZBz0CbWdnYVOh92vRc1V9dkqyQgfg4RzvjSRKKt1QU57Yw7YVEmYihx
kPqJNrTrBD6Gbp413rDYfWstrHNF2eza6UTHbZerh0j+LV7lqWeiZtc94Otq
12CoCI+BDdEGpKe989IUC2KFiF9wLBZ8j2CwjpEG4f7gah/bjP0+LECxfzEB
TZCNr6z301kIchYm0qZypYTJQsvvVYgz3rBmk9zJ31FaeRt07cABJdiWnyWv
1F+V7GN1mo0l/avsM82qIkuLtjR0fUc9M4OUdJeqC72+3GGfiYvHGjELpTYA
r4Rc0x/k8SmoUwytNl+zczwNvxCA0BbJvwgZlCx0Qw4dnzxAaQQNseK/NG8G
PyjeXmkMRDI1u2X1f1ABY3jxlEfCreZgPuTykoJfLLtlV8q2kVdqDWdbveBl
01HN6A2+vKXrt+ipiSsEaIPp+w3jBhhaTrTZVJosZ/kAtihFTs2vTkIyfaz6
yWGo9QoLwtq4NKpXJBwuXwqPPsBnCjz5e9otJmKglITiCtMAkWdzhW7p6DNm
RgYb3w256rDcv99hOtOm0dhBpeBlyj5NoOhWRMT5t8Z9KMrfkhngVqnlul/s
2PJJy9Q+Mcxm77W7Zjy9/xPazzKgix7V+sj2lJ3B0lHNVETu8mQUZTFtjMEa
0tpYwvi3tEsrxvJl93c+jfNC/GcawgfURfFaBt/HIiRKyhT7/CKBcLc1RQlr
74zjJ3vyK4NLwMTlPg8s3IE/wkOKokFH9jJGP51XjOrlNTGEIqKk6/TJaZOi
caS5H+fDk4GvF6PJWCHnxTvpsWYg6y6lvWYiY2lwHxUQoWQxm7puhoW7NVhG
i/ynN0qyOEQ8ZDd20B5Yn4Q4tJofkxM4oAcEZFGqcl0zTkDvTvy1/58u86rn
Ci4GHiEnqD/VbMGAOCqyjdCOB5mdZQ6zmPmtiaZ44ZcF0M7X02uNEOPh010u
1fo8DQWp9hXbInl2yqZbC54UrzG1ZRTZx9K9q3qxDCTw7sTXpgYYjcWvp0EV
apK9kzJjJffp7BIqGq8dlQjMqmDVNTST6ZSqwzz86yoedhKrMld5lXM9p4kD
m2u6+W46vKF/77JQviws6a4HLn11hQmvI+1stQ77wEXDKutI+60AWxFAfTwe
RQ8RKn9kDES1y9KtmaXi0jKQD3T0CJ/zz5+gZACFvw4GoyvU3m3q2Kr7qsmM
J1sol5+0jbZ3SqUp7lCJuK62fO6MhyaRaYbXeyejIMF9wnxvG3lDOuxX7l/W
XG2uI3jb2/2qxgWHlWblj+B5r6CFg0Qlbcoulppc8g1UynfEZdLlxzdkQaE2
14350yfenybJ0ONdRAo3LPW6iTjfgaLI9GnoRdmwfUne2bXZcaewmXuy/Z3P
5inynBR+dUXwwXPUJplIz+/7lx5/qvFGYJ0ZjL+kZZV6fP9gE0uG/iQdEEdb
OQyaPfGHk9DgpoOVoNEl1BW+nrDHNznaXwOCLEWXrrh9VpwKYgzdflsbD/o7
+3YxkIDan+2aUoy+ar7RMOx6YyvCRtaA/OLR323QUNUlFuQjJrsKA4Wdmafw
M57zTopztxbdkCodrUEEETI4ApXkgVworTGrZlfrxxVkxlbjN/Lofapau/nA
g43wp0VSICJjGB3a4hrPqbog6PH6r45I+vPpV19J6+vWpyh+XZjkKhFRRKtH
4v7j7CSK0PCeQ0vhuTs+ALsDLSlbVtrUYxHLGVv5Gqgl6vTPSK3GCDYfF59i
vX20DaPB04dE6rOyQjhDPeMC2Jvk5GTTImKVASgGkQ0f1WS6Moa4NfGpWb3p
PL+AeW+IBqMw6jBMgvD2+NVeTn2EpWENcHS788JGfJO7hvZxoPDW5YwQnmAG
KVPbQG44kiT4kz43qxu+YcyieghTLMbxLsowyp+Usa8Sd3GQP/a3ibNbWEJL
n1p528XCnPLlcAYJbEnZ9j9LO8hEXUvYOFGyAVLiwJi8g8p7LPsAIzcVmJv3
2zo1vremBcqGn3CU/LPqtB1BFcRwu8h9dDz4mIlIqSJh3fIGgizb79A5Z2Sy
w2Z+jQ8Uz0FC5WXXV/dQvlyZ0xTFGnZYK/t40OkrfGIPexIh49u9MWXny1Zy
Mubbw/E9fc2gQUCX5hd1lXN0Uu6SF7xy2Kb8/w0jY9EY+CFqmHoRbEFtQsmE
8kF2BfVoOJe0ml+4bUGTZTNCH2nrAxlEmHsdSoy+8y1opke5fvwcQp/NgMCj
SeivBtGBJz2MatuvulFxQsEw8etZz3gqcTe3pyZtEJxx0Gh38GbKgteE6/Dn
b3nSeEhSM+np0FEfQA2j/P2fChoEZqB/5f354Qu97Vzx2TUqg7VFJ2VFUykE
dblGtGEe7IpyfOMLFl5bKrQ1JZUI/9D4/lUgAC2mfE0Xsj+7hFjYZ06Ce3o2
BYim8S2DzdaOEOxUgmItwyeKyU9vjz4AsK1D9zpOlAB0EJPW7wyWvArXk/iH
dGS6kgtEI4WnXllvrKd/PMUuu2o2BTewAhDj+eeY8vZy8UBORwG3TLZdfnxC
NTEKaTO8XXqCDdu0Y87ALvyq5jheRiSOGsireQ+WvClnw5S3BcweRNLS5kjC
K8A+kQzAfxiT3f97NOajghwAINuxmGft6MUWogs5Yao7DW9wR0uX2GT/5TfO
GsieZouEyzbeoUUfdzti9JW7lta/HnNehgYXBIQfLG5T5kEkjN5gLsSIaZ95
FLXPrsB65EWCEMlMN/L1HNz+65QoAYp9VpuycsVi58HLBjAKbf1nr8aCyoJV
IHXVIX9PBPY5SJLxITHAMr5rZ7yai+m5HCil0mLHYrvN7/Of7FjfuqmOcOQ9
R/+tmuvNPTzu/FEE6ZcbzT4FXtu8is3IR4yM3NpWn6R7OurHxcSsedU0UqGC
MFJRUSopGh8I+Hu4+cUYV6ou3+Z9n5hbokXDVOgqq2flq0K5RoqGNJGaMbPU
OaAcAxl0zr71lc0ZFvunWyuSz/hpNeQ5VdXfmHBRSSCoGfJXQSmsvQU+l7Rf
L5EOhK8abcnGbNYRTk5FA6fJHfJJTB/rp1zim6CgXqcE0PHFVMCX7f2RheLM
8k9igNbJU+dXvyyIR1iA1P0hE9xuibIQ4bly4D85oxUB338Fh97AYk4HTN1C
cIiI8s/+CyNNe/kSIzeNBfwuYaWS5cwfEtt7cb8WOZ38PIYteq8tLu+kEYJi
Fwve7Esgo+4PO6SxZ5js3CnwOJrV/rmbTjFj4hDt/E8WvU6x+1A0GBBKCTJR
CSr0m7hRPh7r02lGPdUd5WS7dFR/OqGiOFkXIDM62gDll5Cz8fugLndAG4Zx
oyGCgjEKFltRpXKM+5lRDwYKBI7lpHtVCbijtvYVmAMEagCcf/aNqHKKpcO1
mcYLwgP0HGNoFPFOS1n3XSkgxc0anZl44CKjBQ4JFCC8nHJkLMyJbZ456frG
9hP9DRmXNCsaDTzZoSTkdPlF0fEzhBA7WCqd/cb4gQTCC0RDbCNYkeH2f1tP
vL5kGHfm+0+OxBL26AS1wskP7EVZPkBAdF3sksD2mDSFzYRiDxtwTG+aq0vB
yFHUaYRsC8mXoOmyOkhcFsVQa/kG2wm8OjMSREvgk9LIK1PkAHTCA4S8/q6o
Dsm8BBIe3VpIXt1n6cqzHc0Uc2uO6T8B01tyK0AsYFbJVVb+y6ffYUsgIrZ3
de4p1KxcRDJ0Sfo342vrAwTEcyGua4qpjf++WYZnOyU4L5xuAffbsor0wGzy
GK4QxkdYELUJdZvGCBo6V7H+b5cRHLyyXv2F0fh5ttNhfhUsXyEPVsPoAE6P
idoB/dJcUIeVdapi9zeGa+JU8Yk35dztQ2FHyavFbofNawMGgShbISh+ovSm
qeoHf+n6vSeWHhnccsE+cSFx2Zcgdeem3kDlk9f2UI8mx8TgRNgFBIcsFOhQ
6FY9lGUyH2NPvOM+l3thx4sKcQa7+RUeHkIgaRYQCd/8LnwkWtfOsdnDzbiG
WJEOf7h5C8u7LBM7ev9LCLdVWxhBLcGyoBLhsJCNUaFHm4lozz5NglJOF1Db
dK/RfJr/NAOdOcaBXzDQLqMd0hPFY2OVMXgPmVb5/DY2+wWZkFpEvqnROG4i
U/zZpm3Ezk/LGBLvkYevdj7TCl2yUkNSiz7tL7xlH/6OBoE1YbOrQvaOzFXK
EnJcPOs8bd2LnTaHKe+9RrSa9U4IHUOTqnxZjHWouoQBE6CdN8UvUwn4DGrc
epotbHE1d5EK9fqT7pzEgQ9INsm3G8WfaDBfkh2VcJhp9/Z6ZBvf0Pvvpxkw
epeyLbyWVPaohl9kBUj+Z8XLs9THnFyoYGPV/Tqdh78rPCsvVvj9LfiuajvA
CRwFOx+logrZtGopQOh5mhI/6duaNPKVzeS30MvTM7WYlL3z4E4JaGm3ZzGG
O1tG+Mn8rgDoC3VnJzwUs6AXIzbv2yi+4im/03kRjuZofBnmGpvPxzOvNxrD
blfLc1a/N5IAsBtifHGJA9VwXOvNWE3iSkHYnOqhCAQpe4U6GV74o5cJ4R9D
It9njsO4Y0IUBrfBiQfZ9TriKW6fwKIDOp80tayxbaOC9rgr0rwvC/fhQRxX
qWJqQhz7oEnEjop0ZUZQMo8qwz1PLX4RoVI+LN+4989m2BK3JnaWiUDpxXSH
KfG4tP/HKRDptKXYyikUp26sPkAnx33k0XR2kIFVigyMlVmnMpZLkj+UsGKy
PB4yZ5A6VpEM2ShCA3ZKSyt+vV7hLe/PMhI866ZEEODRIO5JZuUf6rYFo21k
XeeFhHh4pNiL7VYNoi07xrvvPeysoXIOk31FxwCKI0Pd/xhjMNlo6gPqgG5m
cmia7u6071eq+a55DBnLqhHhbf+bFFsOmSknkSv8scR1XVz5d0DDj96Jvu+T
YXTed29aJ/4y7UQLk0z1Zu6383Bfr6YD+fft0R5cnynn/yRvF9GbV5EPq45R
amDYOpchnhOgkOoHCdVuywIdFgEIC7dsthbxq2i5u96LqTk3yqafYqzv2oW7
bmknhML8Mr/Mx32GzHSLNESO70MpkLJfYO/naGYr2T5TawPCt9OXViS6lkB6
33ZW6Uh5wjE5Sv8bynreNSkg8IYOD11EceD7CW+/e6LtDKE3DPpU8hyjMpu1
Y7HGJexhgzyrngC81Zp5wlAFWQL8/F73qAZw8ZZrxEPmAubNOPGsSBAhNLUt
gmC+Z4xdW0d9iARGmy5uY0erFz1v72r5gLu2Od3vCLGxLuohxbrFnwUDL5EK
Synkf7MSrwmR3Zk7tWCQfAvNR8LN9JQ6+a8CWXIXNJLI4rek+Pt/iMIPQZcA
Z5S5Tv49VUXf6495RLaFTvjcNz6g+g8CTvBZTRiXZoyM9WR85XXnIprEltHw
bpMXaehUIFJP7Eyv9To9XT66M/oISA44HA0tuDhO+abYaXvgfxgN+0SMTqTc
VflhroEiRbIhG68QQUOVwp8+il4s92rpVJcGDIxfNtNEtUcpEF2c6ePWehSS
/xUe0FOXU1Hz5TCu9YS4poRsuFYGVGfr9EEcOiK8qxCaBgQKK1lqmvy1YO52
QIMcSBir2khlWvA87Pjk74O+9oYyvz274fttB5rT5DvienNJzxifX55UTnXh
FfdWUv7GXwuauwGX40gA2ilf7ZMlKayQSPft5Y5x1J1ZbVBm/u1OvmYD+mZd
k/hKGpSmzL4B0RbtCclId+rQ6tSko9EaodPWok3WMvENqrsGRBAK9jjcPHr1
K1cGlhbZwwapeUmIJpDWwejNnz4glG85yXf9bfTCLIyv8RIKigiJ9ypZoPmg
hzEotYLje5uYJGBrEyUwDqNzzY6AIvH7ykoIbuhIZSMBNXoPtdvAgTqUDkkm
WiE9P5kpQFIuflbtVuKKzYIW2z8L6YCM3XChbeaTheUn2CLd0JIEW5W5Td8c
BSplLNuNw2zbjZiX2ldmcdX+C+Os758XJza5OJjXRPYxPgPBbk6mWqgBWMEx
2NCxkkehRV7c0e9FT7AjBp9HzKWV+NlQ5iD5xQl+T4/hTtkwZPDiaO8FH3Ht
PgEzTS0so4i9oBXeGHg6tPfJ+wM9vDC3WL8kne72UFC8cGR9Y92xGMZQ1Cs7
SLaMmV4myCcBPKYSb44yKfuj6BEjkx3ABAw/sYbDpbMCsvSsGC3suU4GDJUo
kxaGfXTnR0hJ2ln8+ggdjetdt5QG6QSPRgpFtUn7bLoZkO7mIyNhoXECDkes
7uRTniabDE4I+MBU7yN9AGHikU7njes22TObwVm6xgLFzcLvYWtR8tYfj9aN
aFptpFlv3tRfT1+P3H+8wrthlZnlJJKroqbpEFf11bO8tEcI1XXLBoKboIAi
IVVgGGYn49rXrYMExCLDqM+8eImpYMJD9bKMCnI8GejYiilA5wPfqPFHznaA
mOuPtEBctMOWAufjsAXj64seZPxueol1PrClh/jR6Oz1g02Z64AFMf7rN3UW
D9KT5BTreJZziUUu32a7FjnjNeIXwwKenWKdIniQ/z8/4Jo0VxLFTWMPa382
FjNSjau6cM8tR+XudmavT/hpcZH4tK0jLlqysQsEVJjq5nqIsngMqSzeZfK1
K+BwDYc5HeE6aYeUobntif5djYQ/pejlVTMRJ4BHFTjHG8kqpQ2V8Ph6iTFh
kI/QvoH0OlRt76y8sdJy88kThGm7/IcdnPINZwAlRdHUxCPrKuAjK6a3EMBg
lDLX6pHB141OtbA4BqofgIqeiYPOrBrUeLSnHVXWWVteyubPDRLRSlvIMfWN
kp9JzPkKLdvVjf6FMYJypEzIbfr8v0AhU16nfrMs1S7Pc6b2ypJz33N9A0Sl
6Anw4YlRWMdSRLt/xQTtPXZo5BUbuYW4Q+1QtEwIC9FkygpFpNipVCfY63FW
t/f2a5sVkdYll2TB/CNcsq2mWyNVtR+XrIF4am7yibWQ541TtTmPbc/4mp0X
xTyBBiAIipcxXe7DqeDs2LkaO2bPHATTsBQqlHovEXNLiBLau7Tvkv7xfWpl
0t9CoiM7VP9Zxwyg/KQItzK70VGyVNfqj9EkFAiqzHGdrpMmOgJhBsy1yCyr
xt6CVdFcgKWagbn9uEHUYHbFfGEyhpMmhyi96zE0IrV15/8G1PHXKrTN5Kpe
oCwY29nrSUdcyglzwbT+wa465/GeD4TghCXlrkUDfIMkay4k32m2LWR7k8Xf
MKNsLMX1meLpdpM2n/PUa7UTr8T2OvW7JbgaBvjrSRwP996KV11MrquvacJO
cUCWPZNbpWAxveFjN0VpXGxZyGaKRueMyADTOFHVXoVTD5Eu4+6M7QsOc5PI
xVcJyDmq4tIq8ylhTFKAmALHLoA5c3eFzfRFnqHbnyMKKp6EUPnQ1ho9AyUV
nA6/wuT0QpWqcCHgxvGo7cHxhnu10Amq+wk3vE4nQfS+PgKgTMg01dxlK0wc
e84Ed3cN0GD793e2FvrZL1RllVzv8Xkf4aq1oyHBZcULiABT3X+7LnWegX14
sRDo3upFU3cfnnUgzH1HXWPOeFunWIoGI8wsA5qDnbc7a+NeETzqWS/eyp5H
Kihh2sEbqAuV8x4/IPTpiK9fmpCmVR1FygCrlTU4HIZICc9li/sJV2wi1PP3
EwL82bZRv2o1/kMidYMoWXr4lUUq+X6leZR9kGTJ14ae/MzCba0se4bHmGKn
aPB3r/2n+vwoPx6YAVnpzFll2Xs6MfZNNpq5pNTV4vN3oOR8zngu4ikHTAFw
JJN40nJKdV102gvUf+zwL8jAvGN476iR7FG4hPSbPBBAoD244v88ymz9FaJg
6irwgTtUhUJkZQGEQCRjfsLQst3vRIruhXHzbMpIkabW5bTJYmiPZ3iGdSR8
zO94q3p5IZ312uXrpjXvRxMuCDV1Q2eRrskflnci/EqAbg8whQVwNhlh/Pr3
P5NCgo2uiXXV88wxjKVuXyzUox8U05JKH4YCTgVkT9yCiMVCA2nF/QHOOl4o
Z2/pSpUCAIKUBIrdHFboiPIbrs3iwOsc2sTGcXTv+clPXEJhYRffg0QvUrsr
KZDxg+b6I/MeqxU39zmlCbzZlRl6UXKsmgerqZjkUbXWqlK4hUriRqWTpvH7
FDMZlJAZwvo1mgy2eeuVJuNaHaG6b1pmYfr240/aGtB/X/jkA5uH1VPBtCv7
VlOn8E6HKNWCw8nKMAyYsE3jMblnX+WW+JHcKa5a2aVsMEFL+8Z+aLM4X5Ca
vQqJmEfomVBWD0YvL6EBn1yemyLFEDYbg3h4lUqw4PMf2uLq9k4V7IfA1nq1
S9PYG8kDcCUuaZZIVULsr7Az2qZoaQI8VaCSwdOCZjNF0pMy56Yl265Iny9m
d+3e7P0B1NvjlQYOJ7lfhIuC+zdwyzK6bzC3igfSsy6zRTWMXCUfdKfirraA
ItWKQlcNLEGSHkru0u7VANhPxbF8xah+7iUwQAU3zeysGh3dNYFtiFAGV4Sw
eIy32pCb4BzClVOYKG5pazD6qTaFyfOSmIiHZIhUwRUZh3/W6He2OygoJ8Ix
c1UlqAfLUcYc42BWAg5V8fKMdkgyUnX9Su4Kq5IFu7rapTjBTmX2lJgXftBB
E/ZGzOPej67ZuR51ZMQqMJiipYj0JWgzad/R0Li4uf/3Mvykmtm+RwqS1yjM
xdqcTZWnTnGcSCRvCKn6B8NbaGqCZYQQartiE9UvpLVjkQ7DDq/823lKDFAM
qq0uCmpyOfkvZ57T90sVUDFJjqaOFLYPca9A+lfgLaKdeFcKMbHdPGQCKMIb
LX8I4WoCEImg1p7R4sdejG870OhGVcVVttkfHhMvkljqRekK3fK0p8bQ1FRv
jUH8cafzhFBruiHbTiyMALNuvvdUFRBSmvxlp9t238XheUtLfwRXaZTv05RD
BK6KqodIJ/yQSciPmFHp7OYWClLhA+X6Y9E/QNpUt/+ycHJPZflEYo3r6oen
CtFEfd6OGzDP5imWHB2P1ZhJ2cACJOQXudw4OTIOJ9QAOd8WoxajWNjkuHRJ
azVNrFS6ACTWONT72v+uhkX05GCCET5AZ8Rlmyf+6vexo595ZQIt3+DAAwJ9
TEyp0+Sye0LerBOGk4kZetVT6uywTpdbZ8FbCxQ5m9oKepwxCY/LiqzZXqPT
k0KHKIn6bOXqFjHCRZ+vDuYu5j5w66gkeEEFoRdhg8sTLjVimsGuemow5sng
t68yWxzUT7kzLbuyB1uX8iBj301GCvTaUZTEJ6CTFt3Bvz9GofBmmRidm91P
dZ0YJ2Le0erifucErW1MelbwRBlGOpOz3HZHYUnS4shFXekbxhugmksc5j5O
EORXxsUxCGsFRsDTuGd8s9rpW0NV9GedKVq6NDGxavDrg8oODWakDeImrXSY
xcx3YAZ3sxPqWzgia9CnV4uYpwsTaWVYHvl+QMC8Qer8UjTwkeiyqJGIHABK
j6DZYF/NiYKB5aHLk92+PdaQa23HSdVJIcav0NeymdIJCLwFy8I8OUAgMJEa
N3xDzkrIN8JLyDTSzq2eaOfT6XgEZ3zE2hNnQWlt8bFYZfGwkMdTpx9/BYhh
I/3HuE7ixpGAFDjDQIitygx4YLh81hXZwdJBYNoApMK7vLi56U/wh64xNyAc
2QkPgSYeT97X85WujbCz0Emd29c2F+WwoDaY1rxZYN0QOGKlnbfNzAorMZBg
zgntdcNblh9KMbfYIabcnaZ0ugAPh3cfOwhgBNy2RxgiCcrAdy2fYFVVZHeh
/5NagEhAql5Bqy+B6lPoBUBRI4WDSIouCFsx6WqdqzBXdWc2QYaukMUib9dJ
+dV0rH8CnqoXE/WoMuSTkQlHUEanbTCclCjifY51qPaIcwes0MC1dLPAvba6
11sF2EBiWcim95tsOqaFU1B3S7URy7Q3uwSKkN9KMKRB9iDcHdAewJiJoDUb
9e5Bfs+3DbYAUUEh5YFlNk2KVLQqRbDD5/7C43TNu28Vtx7fHn86ORPQKbiS
Covbf5xUFn2LVFQyRE/zbR+Vjctinu3VFooifoJ/T7Tv5L53wJewcHa0IRVB
GRW7anzGFv0XMl+a29lBLBZkZUPjlnoo8t9u57n+Q2fGFleXScIPZUyBAqzM
ISvziPdFT7jZq00GsijjPmpBiQoCSJbAtPJVHVLwzYoEEtsHO+CXSRwcTCs3
t6PmTNWHyVMRVjyVlQVnwYI6ndFvzW534yfpKXG9ulyTDG3GxHhdOalq52Pt
khKMeyyo6X36UGYceWtlMmDhe/twbUwJvbxfZb86JDnVn3hsGfynehNFmxOg
VZJAC7BK7cngEA5DWOLvBDCYiAysVXtGu7wvqqG9TxLqZ2cwyxtt9KD26GVK
j9qy49WB7nW4cWJ2tUfEqmUNN2USB6MS9KnV8RFwxlfFmDnMJl+JAsrHy1+8
mkM1HlWT0vYmZnNZL6x60f0Ky632DMo/yrB8A3Knr49jF9DxvrkLJrgrDtex
qH6VI/ExVd0BxzG059xYR7u6zMUbfUGaOgwZs9B/0yo1F08ddJuQ1nwLNTxA
ab7UpUUwtTO6aZpjVClCkyZ7yj2engioUD7zaw4C5KUgZqWYoXAMn0ZCey5G
qT8mhet5m8u9kClsvFXCkjW3T1X2FhRThR+vFOTOz+t/wsOP8hWtTB5Y7ZGY
bMfvmVpkzbu5M7UztJx9EYJQprZ53lD9k0rtSpKssOTQ9tPhFDM9BSgiJa7G
WmCfTxde+FEZP1j/OFbvS20xCQk5iEzY06cBeAzZCq0QF/FK9qdKHO3NniPr
57CEcSDoS7E98tNo5fDoIvs1WyInvCoDlAYBHXVPGx/bFrrm6YWsRHyDPahJ
Ns/0nskwR4r/qNf8x975cdQiiuBsRfkpl9qm/BFZyEyNM3h0OZECHrfgC4Jw
T3+oFeGu6TrGgr8tnNcfLJHmHzXMVKwZbbNaVTAah2xZLkdE0AG5/XT5s89N
tzJ2i0pIazz6rsfACXljeQA1y0J4PEDd4Z+egm69PMGmmDtI6g7X4mnF/MC0
hZoO9blI79EHWeCw4tL4pBH+MFL1IUZcrUvBqZAh+00e2iuYL8lRDu4WLVg/
1top7cF0ElPIklnlGSyUqFEbDQmcAaSKKb3YgbkFOvEp5ML7/bG+3BdO9Bz1
HIKsRmvaDA1qTnudt1RIW60C+cNpfuiFCsn0mA8RPrVa+zUhNLOymLunFD/U
sInSSF1d6inc2V6TUlgQThWjjIU/OlWL3RLTrdD7yPMBQjpsKwWDno2RNhcG
x+NHWxu9cC0hZYXg6oTjZJuFFPhR08e/vVjBDzXmkyWaTlR6GLe0MfVvhALO
7IJ5/b1sy8SLN4bW/qKRItgxZ1FLgY6NNB7N506eNo+2o0pE6dNUzlEVfr3T
eHStwPKwSa9cUlgigOPZSZ9IUnyVqu7q3sGOiGVUo2Kq3BxU42xYVmeWBNNU
HgtpClJjxXoO2VsSwULvA6C5fSOfGI1WpPJun3tDofIAHI/xrlwLJuz0lsAh
nV79yKyOLMHfIB/591PzTfChYSdeJmYw1f2uO4JGB41QE2IM/AdbRJKaGKfF
xmwXyfBl6VDh5e8NQ7qZ6/6QkOKb8BvsoiEccQJO8XvuZibMKXJYfs0az3YC
U62CHkaCQ9p/TwMkv4opRWHAgHjB6agFTT1uMZBPlczJIfgBvg8l3y+PY3Xe
eTKuRTWZI+IsiiKhCOJm6RnP7NSDi/ZHuuLhlNWKil9CypUti2fN66XKqhfY
nRrDipBIqXvai8VGAsKVxJ8TVjV0bzA6daZGy7AFQx2RuJ56YoXUZd1rj9/1
tePnl/BkK3kQ23bAQS0Nj0A1cX5uSSqohrHZwdG+66OAmRwlCu69bdq/vMdu
u7sGC2T/W/V+eEbVY9Cmqz5iT4Fq5hW8dLAZqEccgJgK9LIdA9N4053NmIla
Ol+NdOviJQHJvMfGaf9mxfzwtkMVxzuxHzPyyuTbIRBlyyPwETzWDcPmb5ty
EmkTfjlzKtkQkK7/tn92Q1wkbfPsh8eDEnEM/4wLS3mgNqBPEtf73TkEZMAE
q3zU58YFe099N9zmUZ7NmtRYURy6ejadfc7q/PsRRkrt5jN5B+6hjCECiczu
mxBBYOrQP4wYvZQDqASC2Zh20zBtlP8yBudtxQjQA9lsWG/gL2s3lHui2AyJ
ePwo8yq+Y27inpXxfOEgKSaxbZMcHXmURPtyD3vvp7GLY40nMnZegTCpRIok
15BYX8qdab9OYiwiQy83W2rQuOVYalf/0s9YXsYJ7kUnsGYluNYyeqOBJhsX
YkGPcpmO77MKPV8Uvdj7QwdFy/LAe3tk82DJpvJj4Q4o6YF744BkviSe0mv4
1qPS4v6ukeiemc51Yd77asi3XNLSrKGuG2D3HfbYhTBi3lcNw6rP4zEFZNmN
/zUPCQIkxS52ZJbNmN/bU4yHKakqDLSa2FiTI/BSCTJcvXuWnmyNUjxtqT3u
TqcZDlmdgWC/E0mmVNZGGf5Ey+4D2CtVH0ZogF5jLADTTpUDqSCQTxh1fz2v
rwF7FuBU2CsplCGxi1GdWBnKYv4ODW53t5DCJRUrQJodtSlTwR9YvcwANxwT
GW0Omh6KZuXOsFkfncXtJ+qjNc9vLjJjAVkazxypfDK71QK6xu4MhV/syc82
IQvRqxxNFlrmHC5yXlizCEIgy8vqiklG5b+PwK6WFqB3kgIG4XzGza/FCJBl
dEP8WXd34j+yTi20zFDOIq2vlHPB8iEMm7XIV48SAWORFKfxwWHtElwxB5h7
J8NfuOXpzOQ8dYC0vZzr3Nv625ebokX+E/VCN4u7/H8DPWJHI9q+NCRiNQoS
ap6HawhINC8cec00xqXTMQOMlecrfbknxsQ6E45YkBOY70MpAe25Rogti1i1
d/+XtqHHo6XDypv+uJ4aFEbv+Hcs8xsNDgIT8MfNe3Xj33qVtSa4VJfkdNW1
BiMxw1fW/B3n1+Ho6MJvINXmfHveL18elv9sPbIunCdrefHNCmMzq9MbvyJ5
SUfv5N4eIUYiYTzJXieWucrT7uQCuPUpkxi5sOFur0BoufPh+ELDCytNVoxR
UhBWJF+rCNSYieg2MUewfci4xYXMAfbm+1+Xp8GAdCCY78HWiRzVBHGm4Rny
I2j7ByhvZW2jQxwSPR/Lrvxscb6ngoccey5WLl0YRe4wGIp0fVrhCCr+NNQ+
Tg+jxz5mOYVkLh1qnXwqrxR18e1yOgu9s4+8yYaj0U57iZfsjYsKXt5S4lC8
swHmLXE4qujseRBdZtg3sEMRR0mAhiu3s087nnLBInNHrGrNKHVHWcRvNneA
JlBiLMOXGx7QCI7pcaTflxBFXJpt6S0KDMJyN25hfBaZYlgRJWL6LLUr7C/w
trSgnyf7NDyrhG6SgiMwQZxRpmtjJdspstGGmgbkt0SPtid9NBdBTwxdSF4t
/kWrE8Ncxk+GqvcQWcNTzZoCjKwdUu0ut+bGELBeN1h5X3VrEV0VgsfQnCU+
dwBWRf6mW1c2XK/ksusTD3XqQQoVCMGrm8gDd6sqLX3vmRVrJTkIyijIRXFj
Cd1rzfcHoh5A0BQgoNfJtKYc4QBAFr9P678X1hQpEhsLcPqY2sN+VjSW2u1c
VhQcgzi0QXPgJaKBAXrNsPobvMl2ExC2ygjtjaeLh4GcV+zKHwA84AYTojhQ
p/uQLjtdSs1dBz55bH9Yayc9GA5MQziVV0/PVH7sRlWXixZ3HLMo2qwPB/B1
wWejpHaJbC/oBAs6BGXwSAnHiYUVq0Eww0aj5L2cRVlMOlUaKMQPYlB2c5Wk
Au0O3/Fxk4/dxn9ZRA4CSAv1G9BA5Me2iLCFsUA8Uj9RWDuSq0BZ7c1YhKX4
jVq+Bei8yTUk7yy4GxCf8tZOIUkhMEIaESd/ZhsUBjvj9SuxsocxmbEImSZz
3dYsPHj4LsBoeF876LvKSKnwggvtM/JByyEA+kvM+RsY1K4n5JrHdTNaX8HN
32u+kaGEyCugaWoYCiZ1SQ/2h8OueQRhW7S1qcFinJlEe2SEvxwAGNmSXnfV
D1DSQExAfobAOF1bEAWJsjoo8vAQbFZjs6TsWfqpOCtXyYFVEzrByiirKlUN
6CpoT5PUUOMidSvOSibc615twaNkoY2WUu+P+OWANchq1NjR5tcal4iOf9vP
kDKBqyp1LBW2d4d5bW2oTJ/ov1cF55aFLnfjK0LEQ+WAyyGFbfXReKgpz6zZ
PKmP8inyuTwJ/cdUzFypX9LK4YJ/5cgwsjx50DhngcnpcaY8tDXie0F45t9q
8IogXXaKUn4KihjsOqVSzrvLzFcOEHJzQEo4C/pEedimg3CB/iPzguiqcWqE
0OQjYRS05h6PfttxsSWPPyUXZFs7f0Mkfm0fzn9Y+CyBqPwaY76uE2Ut14H/
mlmtFR4Daon76v1OkHZRjWXaQeAU4WKqf9FpJJpsfEg9/+QveintyskAP4T4
MEQHAb5foGWPNUmQW1jH7SRZWggfO0OvPqaMxEPVbGXb4dlO5s+dV9Mcalry
pmHIUwDW0fj0EdVo9fEKbKzNmydLJNfz9OCBWTlwSP4frUScHrdPCN5jzHmc
xdZGc9rfdgiT+ln87Wg0A83cKWX3jzAZ2hzbVsWxCmV/IbgHcT8a5qhdIILz
XazRtnlz0j9b3Qe2fonDeq740kPY7+Vy28WeRPoYPKlEWcqtnuKTzWtM8SPS
rOzxJcfFaZOhr88PeUjZ6t8U1K2h8mM75P/8BaeojMuexgnDeBLHLOmppuNi
ZzBqk+e5AGqNRa3FwJ9eiylbw7thVMZ7Lxh4K2BWrsd1OnOyDZa143k7Wk34
JaFoD9ZniDjiiloO8fpkh+49EAsAcfOPWNrleN47xYxChqMH+srKhVi/3fYL
jxAyppsa5i5I/rrZtPQ/rUt9+8uO0HiUtMewIPT8BR8VeeCjdqkLTIxcGM/b
vhoAl5eeUfeMZHjxEf0bpatJnEV2AO6VbVfakrTB+TIonI4q3iJFRXKDfa39
jilWiPsaxzRpvT+GI2XuDQ/DtrUVPFZ0ZJ+ZZ2k91h/ebX8bNZXMsKlEQukb
s06eB1kA5jEOc8H8dG5QrftKnIhA+qJW5Zt8iOKeI8a+hG43bC5dMr/qomLZ
XCLNV0IJl8pccoShIR+NJu21sdAApEPSkcUfhIPY/NOGGhyUDhHXVBl8OBKS
QVbpWRxxdf/5eSdcXi7pa2x20/JmC/QNMNIPj8ET1jYrB/+K+UMMMlqqE2oT
R/S85vzatrM5FAg1inCnkrhJnhIrzlVV4TVca7JO55mAPOGv+EkYzT+faIG9
osx0t6Uk+74B/BfE4RkUasctK481h5UFSu5aUErwLXDCscorqBdEvPu0kpU1
+8iW3TQyTa+TQ9quGwD72js0/2pAhpZkwBUDDo7Cy1WKeX/rhx6UznS06T+/
wdeCNfT9Vv8cQW6EaEFdzwcqevWut4/lD+nGCKOt//sVyYJlvjpyTATB6cAC
NHiHtZz6XHskFJCQMK+dJl3gxu91ciG6gdIuyoV21D+2TCQJjJ1ZpaXItf5o
FKiA27LyyAjf7wyTzKddpYD/ZJEDO+t0++XmErQbx6J8ejbkMmQBUuTZoL3r
HGbevxIuiNQO7jPpgJqAyYhQLg9jz7ENPjDvNPt+p35rG9HkgVRMRTmvpwS8
s6Dw2yTSx1L3GHokEkWoOVB83BHnMxYzOUSnyhZGeehrKWP8I5MzwLnSZBKt
muzN+S+8EX4lUHmD5zgB1Oja5EIIL1aULYakr7y3oDw1x+wrtcrzqWLEK/A3
KlZQrawGLWs9yaNw+OUBFOfVMUzsTbQgfIfMyrhlzy+JSVwPWUW2XNtFydsZ
EC0+vjfvywdBmL1uyDhALr1zgwu5H+XMRTy9CuUYNE3cUCQEkUYDdMw7NDiv
Nxwv02626b1AZnsVCxFdWvdpcZVx2uyMk/8fqv/RBlRPY/Np/KF+2Jp0r3Re
3kdVPiErbUYHO8lihzgcjgLiJkSaCd7Us5xfCxKG+c6z8j6xRBK28ZtvHh1g
RPyQwYuH5GvZxizFrmTTmIWg+Zu8CdNfj2UvryWyDIgPh9aIgnmaP8XS6Tnc
dVo38SjQdOchljZLnsCNQZ61bO59Q2keOaSE9yYDRy8cXievsK8T/806pObo
MJ0B1k6QKhUl9vt6gEdFTQz6s64tVpEsBWL7KTXi5HEJY0FC6Nibm5ezdqvd
T1drjQ9B461KoHEzX1Om71ElunnmtSi/ZniP/yH7A3h1DoqcLMoEjxRKeC+P
p41su9js3Rl1O0QSgQPTt+QMtuJs2VQuuv0YrqgPNFDMgzHqccXc7dhpMhC+
EQ17Ai09szAELwzUjM/gGCcEHeghpUUaXlIJfotWjRiyNKn8W2EEcjLAlVwS
U53wTeGj8+tuUj/2smSHDAPjVIIZBvinlnBQiReA0GpsKFH0iEa0sIwofdSi
o3c0WMsct2Ziqv5Ej3CiRanBw05mJo0Z0ae/a5NJg7HzRNMEgBH01iIahMwI
QtTVaoIr0400hWN82Y2yls5Kb3OD/DouoSmuPAJqygT9kK5O25e3qjkzEWFj
Td5NrX/SzFyZgO4Ht+nxPK2hRZwJIqLKNIzfxf1kJTvfDvRzpfYNyfjpBBBz
2YFXu1Ysxgvt3FDzn3WIgnnyZB/XvCFesNzQHaMwp06UUZIuWjxbHMT8yrbT
/U4yQTUwo5bdcVcHHJkSgR8RkMbee4SmRb0kw+NhOMMs456ygaqlt4wuW4Q6
BCchT7eYgD9goxtUlYRHrtFvIy1vQeizLj+zoMXsOfGyN74CE61Da3s86CS5
GN268o356H3Fy9u4fWhC1kCtzH7tYNMfX5AzoyikNgsKj7Acpfr2gkybh5dh
fyNFvlL/Iza1UhOjwt9kijbPH/E0VerTR+DFPYYgTheJ7C4d4+gx/sPlflIR
jGN78oX6e3x912KUJBWvN5i7uZq21bzOdUHTpMMLlKIv98UEmwLIqU+ztgFl
PR2Uryep/xNvhgY96xCLbOrw/P1tgIikJBOLQ/5PglxEpVyXIOdYvFjRsXPB
MKBzpkuOpGLjCe+kD50V0EepQb78eYNSNWdlY0cHKSZQgoykgRxjHkLx4jgA
czQLWeU9zQZKD4txpyhd4Wx9OKb+UmBjuN8P7dPWPMFLVuAFsxis4YSlBr64
wXcWNwMZGQySF8hwmWh+wPasRKCAeXAjCo52btMeUr9f+WOUFOboNJKOsfLI
2Bym9s7vY0Cgu1TUip/Kr7F5xq9Aih4oeyLphuwfuYfvq5YSVtd//td5iNRB
lNn1scF/ZLa7CzFY/ds+KEOPVnp08+RvL+ulpJD9Z37eVQ5uYfMHJl91N8ic
4BxKP5Xv/9rqvXIIwFugsWYhQKdFEm9CkgRF1ftNkmKg4dcFzM00zGNmDA84
vyKMmvB/1nFu1AjZ45DOEJlNnvwfIfKeJe6Fd5ap0Ev+RkFFQEBpt/YOQHG9
KBDZu5dV8TqhupbmQ/45ajBbIlaijGMzhIgXGGN9GldyNN6jsNBtO4x27XNh
RyLc0SBn3e6TThEUKsXuJ+jX5iffBJXEs+SDIhsd4bbexqHYLo9Ap8E7jEVV
bmNdgI+AaT9nNX+lmueszJXF2A6HpK8TeFEhyUQPqwgE7kpNKsA4SdXSOLgD
iq+M/D6zCCaqN8NIfoS0spVX9AekoDCXsWNI7uEKlhsXjcyoF/ANtmznufB6
wOZE27VHsB3urqPsuwiQvfPwmGf0JSFC1vLzrz9etAb9ne01QuGN2T2opzQk
FvLUJlVYuDp82p/oLM6Vy/joyTnOLEhnMuGMKdwx29YeXCHRpZZFVZk0Pyal
YsP4lIT2SiNZqbe6UTn+YVMULpSM14gcKRZztstW8hdF26oHmrh+eUppD1/L
U/vH92JwNUKqPFEV/r6xF9SrD/J2OH6Q1K2JePx6X9DSGlJACcNjO7zE7lBa
ak6GfKI26cQt//m1lqtnqYM0H3oVDtzDm0TIdeYE6aiVPbgOT7oo3FfTn1Vx
lGMnYfBxMGdWv/SUoQy+IEJGuQ0sexonZmiobH8x7z99EuRPcSoV8aGSuPLe
6+HcAKoGD1KQnLr8wC+sdaxMu3FrYuqmWFWxOwLPz//HNh6mxVZ1c/VuoSVb
gB1UpqEdv5zY9bFqAV4tRUeUDb3bXPIvxGzViO494ZV2UoOxpKJGDlkOr5Pu
RSiLp2BtB1D+t1rmU54ZwAfBGykFYQuATfav/aPLg5eDWYG+majE6L31PQk6
0Ow7HQVbWHruJ2sdmLMJpf12RDxl5U80vZk5bQWs1upKmMCwK8+pKL8x3A+J
PggcKlNYbECWdxEOIrv27R4fIFGkKdml4EIu1PN5pj+2+8t3VP54MzdgLQ2l
IRREl2iRM6XW7kPuyg+0RZ2XxLjwCazSv+xT9fQZXBGWp1cYglHV+KHR5bzS
2sXMw8cN4XK64MJFMvqMDEAVoA1hryv5II5EI6w9gASi2Gtd+XRUfplgvbMn
mwSkQeMTaPlQRHkATQwZ/jUKkw4idYRpyMmDj7/THeAP/152rJSj2eOrxGhh
JC/qR1F6kuvMd+Lo4+rYORhSKcbcFA/e+oYt73v2ug0ulV/B3mnURtmvJ0GN
z2BVlRrRr4/SHY4nDz21Px0RbCHd6VazlqRgsdXllAcu8o1n6caSBDwrsaL0
g6UZT+iKbL2AKjV9VsFi4t6QrkhNFZOLvDYLA5mRbjgiTZOYZL0ZvmGmCvU1
f9S/eS6kMsvv4k4zWSyedC2pWyL6IJrEttX0Dcgz+xbE4RvpqQsXFRxKkqws
t64ghFJS4GSxTq13UXav0oAMD14zqWW2x1pDOpMY4o0P4TnEjJdT6mGnaq7y
LZqOLWncBi/kXlDJsvyv0h2EsOvIfIKdadbmMPcBxnpL1qdyA02wM+ABSuu9
lcZ75GzRyuwCYOU9FhXPLBYOUFgvhqVXznjwQheqGc3Sm77zlBQEyrrQarhu
PdT9m/On3itHJfcovOwn/x6AI44eHtKoRGLJDWAncDM4qAbwkNPtgJzas5Tz
nYOgyBdUf7whmWMHG5D4k5uuwJSL3D0yvoGkRf2f9tmTew8HcdF8aeYK+E0D
K/AcWYzeeqW8csqsV5EfYFtqdF1UyipXAYBHEcwEFsP7Owa9PrrfiUOy8H4p
xK+51okv2p2Jv+OUCwY+mAY/JcGcRxa/3C1/43gbk7NdXRdQSVGlZssv1r7C
4cuAeAWI+K5lGa2YdphecdEibBviL994cKnBG1zCZHTAPLeNxuY6Vjh7VrIP
nIMd+KfohBoTgke5WHnFs9Hiqc9GoOyZ8F9bcbfMdyXvk7q9EFYhZ0IDwdf9
4a8sEP+hph7vfLebCWUNrVvHG0LO2FP/Wk9Dpbz7L6oJY0oCuX0ijoyrjkvF
AhSlvuVO8KqXdPBXclG2U77Mg2RoPOp1lENQyANI5KzRCgvnI65av1sPOePX
BPmVn0hYKX2CII9bsQGg4SOcZL1dZer8BEw4N3f4WN27IkSMAKHL7NWPGcVX
R1e1COMUTpHsATb2l+vx3KG/EzHzurSaLZp9zHAjHtGwWVOSFk8gjJkJsLKk
8IGOyttpQT+scEGt67rXxmKwy54P+x87g8T4D3w7QIeBn8UBbpskod1q+OtK
IQ/PiL+JzWXTdOxVn8zDGEH8wFtxB0Rhmic6UDT/9a92rdqEhIB+Wbd5zze+
wSOJG6Ym9vuXL11b4U6ESm6MpcDAVuDectbDIMemCg3o4vbwlLwNOaE7fCjT
EZnWK4ogLS1++kqyF0LN3y/yZYIFzKlgYTyORQtiRAMo0ODScHW0sVH+DXdC
yQBmXaI6/Ti8aawX0JUp8+pZBS7gpeewCaqo9yQPmX4scXW64QDD6gqHwneu
Gl6EL9fj9Cwl3DmT71ewfD5x2ChcHdIRqzuSAz+tW4ZcMyEIlHtK6AOUc8t3
dj2+yYT420A069HULBLWlKdCaTJlRUJmQplsjojYvdBVdCVoy73zGpw/1FZH
F30vd357i9fLPxBGfS6RS56ZYGPBpgIAcMdEKZb3HHOUTNAvcPmYhOeKI1mJ
6WvyKUrhBGFL7uf3it/P/x6B2cxEnZ1Rqo8k5uDFH+BEfneyJtXFuuww5qbN
sIfZpr/sxl6P/PybDFJyy1Rcf5Ws9BTmoUj4IrR5sIqKEJ/b7Nwqhe0ymd0Y
mbyvIfp6VQWQ8EU2rsY5mh74haCW2vG+Fpd4pSybFrhHM0CXVUAYIw8NvRFX
0Bjml2d79FnsBG1X7WWtcNKRjpt4Rjiihdv1fyxpMTWHwLOT2+8t38z5H2tn
DKCVltQ2skTmZY6pfQV/HMgjNHMpcxSjXil/A1wQxV5wWTGdlfB/sp6RYDob
gMhRqV0bRmVVipledRC987CRZxbhu8gJbJQUjKUwweq5D136HbPUTVVdeIT6
7c9/qeOs2toEMB3pwooL2gMbCpcYicSqP/ino0lIeNwgWb1g1TYMYteuVCXM
u/QR56scUuxaUNGI79nzT8vQ02mWUCUhv3wcaptBb3l2Gk6UQxQzsuXmjLcM
47piARJd+dJWdP/izRfMMmDsRvOxcBYeId4u56gf8kKy9/NQoaXAJ8RRZ8hA
VHT5guUbR+rUs0Lesdbe0YIW0YdYiB78cuNhtH+Dbz7y56c8CMWfzPp3cXdX
js0yDUJeDcbntpnodjgBIM0mo2mDBmiiOeCIcKabvNBTPNLxmUXNZafhs5OE
9qbFWfcCI+aLv2WZJXMiikPnsrXCyga7pq25XOAT/raVFQDGT+Rgyk9RViLJ
rZL9jQXtuykZUQHKSLNdl27jTer6kCc6NXIzCARWEZvoOXmlaQoqzMP8IIvW
IqtM+LzVVgmNwMPxYg5+BIkUlPeqQNgUFH0AJYUg7OzIqak6+Y9AVyv+Ltui
240npx60+cadoHV2pbqcAF59DzgTG+Gz/LjYEuv2JG1nb6fiL4RC7fc+e9Cw
cLD5li6PDqsMrc2PuKsJL0g4BZG0KRkeo2ZKMX5h4DWIvnu7H53zb3Bermyl
dCi+ed7cEU9orGk38jDtRDSvu/is2GJ9IUxfbXg1SG+e4eoBOMXHjRuOhMhj
jEeV//XjpA1xRK1gCTd6Gge1xoP8VDX/5vslV+WWSARQK/zyzcKsgHYSyAGl
pO2bDjTqLsYXOJIZCqftzcPHG3l0O+apdQ3etl+3fIyy8haeFVvCEeaAXwlk
JW/YDVj5g2BTmNGnF+cIl8+hqEG592OHd+pIzM1uWUcdrQCVap84X968Sqku
mVTZSEKqPS/1aq9tv9FOzUvZQhnNmYcBRkOtI3715RSyEiJlheORPav5hjyg
I96UVlzhQ9Q0dfaEKcW8NOenrE5Cab3/1pnW1Wvcrm81PVxvuTlUBWvLjhMh
Dzj5CsGCYmOXwDciYggfwi8o0Xie7TvOi1cgnXsQN7oiF5FW7hgVi/3zIzju
CMl2yrUyhsSr9ZBDNp2qb+ONY9ZKBamoT+Qe2NLbHDraUkFk9D9SQ0Ya/DFX
FbfReUOU+yCUVTnY5ro9q1/64hch/cbflTFeeDv13VCMiOOJHyLK5K+NAspe
mDSb3WlpTHmIHGR0Chh3Dzeopg07aKOWVqreBgAEFmFxrxqLZ4IcthOZjGS8
UuhhLQtcWP/bDf/9unAiXxP97xevGhhunY8Z2kT15oHUIvP6cFV10Hm9rAvq
ZlydFuaSmkhOAWvbME8i3T1mHCULRR00AhzD4N+9ORI5z5KPrf4apSPYWaev
Jq76Vgs7CLhoK0ynwvcCMUO5uvhUk8c+SnsMWfnmLhd+nFwLAqDJoG9D5Yyz
87q+Iy6/I7EPXYzaQ/ndJRt1Fxr/MHYmv6qH7qEbbYk1vMO7vFr8t+8MHXTs
yFcXNomEvxkOuUrMH6Do4EbIWLCzspFqB7K8d0BEDi5KhjUYcceda7K2quax
Ihuj6ejnLwNWTAlHZ6z+DFnFURCigEz6mDcndpOx+3AKV33w3h+w6Dod54rr
5WELP5EZRWOFZA3mZgjMazBDiiKc7MhJLyUCrls5S7N+S0q+QkHhPVaAq/Q7
8KbKMKvO+cvyx4Fdg8t3H7Kcudha0aOqR0vR8xGRz/dG2Dv0K4dTi1DjiUsi
colRvgEmCkmI7LNW91ciLFsMPpaMeSSIU6TGBIpPTHvQRXXNRVv6Z00mzPnW
DwgqhmxRzij9WnfqmL4O+aMdYu2iDWG3W8gvTZB3hoojQV3NOpYxoPc1nKM3
WCyeiF6yxFBv7G0OyU/xy91gqlbPUNmgToVtFb9OgDGJowg6JmGWNFzQKoZT
hIjfshRGIZNWmcyUNrxh2zkrbsOcAHx5bzdiQkptVAioZpjAmvYTyDlXXWuY
ajKqIxZEnZT8SBP1fxOSytwrJCra7Pay8NGi22IzpUIP/ESup08gfO7QjTIH
mT5zGWN4/Dz2NHqcM3bJ3n6n9ItaTVpk+MqTbqKAGfGM2T9CNtgff4krqHsR
nJHx18KStSnzbGt0fA9r+w5Sylt3LL2reoSemz43SadN9GTES0iJoSS4Ogao
boihbPO/YQMkaVOdVSinodAkGLyQILkmfLNr1OPkvRU84tUE7hyzFSdQ5u+3
j+ftLsBLiuhBBwtxEW5Ng1t2zj1Em3D0pv1+q+diw8rHizqKJ4nyuOhimqRg
BYhzuvJ40satPZnQ6CJyP/+lVdSP/e0UpmQhf93Uj29muC/qfiB+WKDDi5he
q4xs6Lc7icip+q0QgMcMroCtn87vN0ZRP8l8ALYgIrLyaSGtsIcaP/Neg8nX
eVu2jMkdKTyj1lJCq0J8FgZhI5p6WZp6F6pEOwHLP3sMOKP62vm1p2vS7wyK
II8s9bTnR/VE1zfJvr8GHKKYAN/1uuZuhDssTNV7U+3jD7BqbGY4dQGm3tYv
Ym5d2E8vZrLaMb7CdcCBFfUUZ3lB0aja2MH2H6L1D2ZWVTQQOxghWPykwNtr
40bNi0salIQlsvVhSX0Uejk+uVt9ffw7yYDwmMxK3s1dnt+6N0GpMGXWYMK8
f1QZ3sI1sYTiWJjETMT6hCTMzQCJN+abM6SH25aV+YyyY2BPZmzg6CpifCK1
/boYFgD6pEalW+1R7JN7TvWG+PVdXR8k4+G0aD5yykIBJa7Spppjf7hsSq5O
4Kkxe5J4sZlN3KG+MqRVC3Jfd4+4WgNuC1h29iBwb1a/+lNBRYsILGIc9Y5t
hdMI3VxA+2vGxQnxmBBaXNaEaCoCajhOVaitWo2CaqjZWRbQ0N+p3Uw2INBa
HZan8B52RVO9aoD7VNGe6AW/ahi1zgQo8lVUvjq4UXeEufazNNmXZ5YaAGJX
43cm+Ju2lSvxS9aKo0VxX6lda8TKspvp9DRtzbUA35GwRdfPtf2qckO3+4r+
IGvVuZTwOSsdlJevMUL9eyzfaUIKSdNHRBS+GHH4MJFnvvvvZZ5xGd4hfOxJ
oAWJ8TJW1eu5gMz+BlSVaFTodVjSoY0EFOWS2E2wskRr9CcrdGagaZd42UiC
QZ1c+Ftg7LoDpDWkOdX7mw9lqhUZmAmMhQgPuwuozfG3FNKIbk1KqFDVFUfD
XdpaT3jaxE0J0sE+QZSi2Lb9FxsZtsLf4SqjgGx0W27JCV7CdMa5rGvZt3Pr
XqBMsiVctBWwnAcx5xp9eDaj0u483OoJRFT3GB3Z0oN3Oj6RAc2OzAnW1hJj
89Y/4LHayGIC0Kg3S7x/gP7N86fSnxylg1SaML/FRU+D7CZD6NdNiYw+NnzT
lQd7Ww56cIrbMvRQa631b8u4gO8b8T+xrlpp1USWpkvkCDC+MfvLrgajUUro
DhL0eqtbzGWbjDEf8R754X6whhkuwGf9nx3N9wzP3HPs0f15I/wiDEpvG/kR
aMLx8oi2JlHcxAvNSYOgDzrHH0tUpg9t2wCtcOH/MX3DeWwswodHYwATUsz2
V/i5W2fnFoIKA4mU6/I3hyIy8TCH65NiwmAU7ajonIzupjjeIxZ9l61fo1xQ
p9GVvQfe1GgE5T3ih/OAsmxby166+Gp1ZjHIKcEr179jzfyoWSy0UmP9ebDZ
U6raWuro9U7cH77yLnEUVWP7q8zIBZYjnG22xnENvq6dpYKF+nDokyKnKcvD
8NDVaVic50hlIRU7pE29BgJb+lBkGWI4HZHcPpd5nPio01YTXin+pjvds2Jx
+tPzrLNC2tEBoRM5JUadPyWj67WDJTncctHQ6QjaCtj7Ea+O7lOJQI7Lbcuw
X6xqjCLjfl6Grq/PFqe2XNCISDudpKbAo+Snv8wIxzCXg68lspyfPzDz8A91
Gw+bM0O3m/WB+L7wldmkDH1nWQnE5/PqJbmspBccW+q5A7LZ4hqLLmEnO1WZ
LpGbFeUndYRIGkNRXpPoGVKNgUonXrKLJSCbyuzTWOu/LVagNf66Nzu7Pwgu
63G65EX0GLdj5OsPjOkMcOsrKP7mgtPZnQHZRRExQIshHpfe765EuGnT58BG
JcES43KFQ5ulqHULLTGk+0Lo+z1epAn282ydv3rNL/FQQEPwkEJsGzC0OGRi
boZ6t2m7sgzJhVvi1ycOhDVW1kehSBe118hOsQQpCP3rvR7T9+4Bb31XgBHx
wvUHKd2/ROp7pB9n0EeuyCIvbla26fVMz27wQkX2H3KnATumLOrJmqXrfKBT
B6Eqfuk4AzF+enCT1nt/5t0YOQ7lMGEDsVpypOvBR2gMUp5+WjKRJZjEat6D
3pwmRoGXWzKGmEYc7i6qzg4uu05OkXymCgKN7r/txBa0IowbOu+esZCl0hNX
GuKlMBd/QLd1OQ7ojUTVNV5UeZ24Fc55PYcluA1jg7cCbIPNjlK8Twvli2n3
DAFMa4XM+vtWdobUyDrJp8wMcfey9BA9YHMTcGiY8vodurQIFP0ANRTkx/wZ
Ua1YpQ+bW0Lany/E+Nw/wN60cd4hnkhB7JRtuPsa82BwIDJyiEbNoBg1VB83
Cqv315I+4VEomDplvznmLLbA6YZtgNhmO+pU1BvbPOvVR1GL2bgYSUbP56Ca
cmRtj+mBlWP5uWljQU22JPOwGaf0Wf9lJxQ5Pdli1Us1jArWoeWHqw/mjqO5
7p7oj337LOBXDf3P2Bgekk6HcpyKAKkN7SVkSM/BOloc1iUOK/Jm+PU4m8hC
ArloqCYJ3U176GauZUjvoXuMywZyocry+qLfxFTO3/MeneCIqUEto2Nk+48z
ReXByQT/nK4rnBvnzYCLr8A3q6QvzkmOrZyzpVCWpf4k+Y4LDj6yTUySxIa3
iDdWe3UQ6F0w7Qy9hTevAy6fVzaWN0hONNTxwvTOXSmwG6ww/u+G8T1+g8I5
ip/YlTAYkds/4lJ2eH6n/yyXo8QM1Shxk6pFkTsxm9CVVYjG4hxE7UN7kTBg
qfqUf2qkGKx+yPDaBkXCWcnVRuIQtw0+CfgGfMbTZ8DPhgthXy1fyBFehwuy
VRmRlCwyZKdvjE1W0+5dP/yKJJ03jEO4J50odMDq0ynEiUkHI5jnmRDLMhIM
xlDcovWgzct1lJ6coZB2ijrlcf/8EZF7EWpgD9erLgKDojkntj+B1/6o2IPK
QY2XEbjmCNFARxEDtUBrmDLtSuee0cfMz+hx+rmGU8xX1W8AFPCvX7r73qA7
6tJeuuRgtA1woCt2+p622THZGP63/7p6LtwebBC3A8GbyY69qS4IGTmUnI63
/2xRB8j1JfNIBzsPIWgE+rKtIg3qaCK5OA3RYmj03Gv/N9ilt0glXckcRMQG
LIrNRGXu4NJ6X+2JBG9a9U4EHswiQeCm/JKgkYAefShWP6go7xhHUXswKMsO
bNU2h9q/S0hcfu6mgxW+HCWKIhGGwFDAr3SfXfrI6N5YFTGTPTOPlkiWZ07C
Gpz3ecHj0RJZMOZQj+rB0zcXiGVRgYwI31fQE58NLBKI3MyX5G8R+n9sv3rJ
S6ZHqCLHBlG6DZZ+vZ/yDAYode+cO+we8W/QINMgYXCAIqpGQv1F2/8LF5k9
huxmQz5a2J9Uawz7dNyPccO2d79/JQXseph7isKQiwfeVSUNbbvRy/ahklB6
/9zphfZsug4Hexc4x2k3llrqDwfSLAS5DyU5Zp8zC5a3TAEKqt8VhSB37k6F
7h3B2p7JmWEwYcOFjgKB4+PHOs9xoqEbD4F0wC8pHBeU7jw/5T0HHaQjyNZK
jLl1cXVhysLmRF9Bu2dW7mkn/Ypbcum++a/Ne9wbq0ojZqhD9ZYEY/xUvTKc
AojytkZjQicP53Rp1yTbGdksSF5lxkOi4MkJI7qlHl1GU4+XqIjn67b1y7du
HbwTOIbILcKMPXmN15HcdgKEEhOcELeTK+cDmXj/87WA9uaGqH32ymJZcerm
RTCVb/FTz4WRIjgclyHwDKbbRNuiHy6IADOFhjC4OAA/A+KBT+dlHRPb7P+x
VyeImDW3T/isJEWoZFTXVlqyIFhTJgvu7TdiTMUFxcUMDje59bRco7mCwzF4
DZ31B/7Mhpdo0SGmv0vUq2CxbadPXzNHpQaOjmZ6F9IxsYBMVYZsjYDWdZ8o
QqwqfbqrPhcITCSfUiuiEEFJU3kXN3NcLMi9fqhe/n4Xtru2p2ufd+IlDL7g
xMyezfrN3wPwOsZNARgjqvyrvr8AectEjftFdWPAKT9LMTStZ7Sm2EPNx//o
XovVKb+IA6Hv3DsfhR2++6FDTRmSI2ECd5D2rPuMgDIc/g97RDwWfb7KkoFy
mc2ggNTovYQ4qq7KoR8InPdKGBub1R1v6aZqb3X3ail/3q403eBat3CC/YvQ
bGdvPFKOMY1/zxuYo1p1ttlJexEUK5LE/ljQf49eBzRhx4u9qdei57S3n7Uy
Qa/InBJdU2VcnJptSwb4sNIzZcEGXQ9VtlwWembNbpCOy0+L52f0cWkgx8om
QL+o6oCxVYvO6ch8PM9JtMRPpOIO9riHHkC+KCES8JpGxON22DPlmJvUxVMU
L6a9C/Ei4aI6DCm8HYkSx65mV73Pr61h8JuyCTT7ribhxR23OeA31fx7xBNL
C16RRZmiasZH9c476ei+EBi6qwyViH2EfRcUkkDiEIFtyvI2sOxbEibA82Va
4c6SsuXmuHusdzrGJG6MrsjOMbL+noSAjUelgWEHyXwOJQLi4yYn6BTrG57F
x2xLUFtnMpjVhJJY7Xt1WOjHqDKA9xMV7XHeZ2OIAanwVpOFji6YhQnDcaBi
43zz4VdwBoq6XcyScNAEJ0XpIeRRQvtB9cMr/HDHHAX+p0BBuufDimLfFLnf
X7spt4afuZTPrk6r2y9eMCIdNQbbvEnNxCqpZ4vPZtjAmDFcezFv565uAASU
Eb6VxQQj8rC1Au651qbhJZgBfuvoIaEErVLPO8Oig9VSHvQP86ZL4FmJaclJ
miy1E4GCFI4k48/Goa6RP7X3XJf1tSZP3lrUDXSbKz2xE/fQwiHmxaCvImzI
60/1ABZ5qmlqdLVtancbnfwl1Tx9HvfQ82gztktFRCreZQdLa/67Q570sRnR
VOHXdAAGJuNM1DRn2g7wnxEg+FwvOeO82nM819V8YlqZ8ezLvpkhxN3EuB2+
iQFtAHXNPssGKi9ze4lMsycQysey8p2fW/ShSCw0/vvuWh45j9gmvuaVGPjW
vN8vcMPL4xrJFYTXMycaNGY7XzpTm8zqC0/3WdYtAhJECWMt1egZYojJ4PwO
88N5wqmmLs0HoqgUog/e2sjm+eCDL2MERK7mCBVAXrnSeFz29FJvq91hSvRO
5h9vBPVAny3RBRRwgUetzprQD5S/tac7r38M3Y505zp5LlR7T/uzDKoi1Bdq
hx6yXlicqJelSyDqEhcjgdC8hrg9tOqJO+uz5vhpLr60mzYiWou/v/QtmpFx
z/7Y/WGXvGY27Cv933HGwSmpXKrZc0ucOfl+TJef3jnxmfkKA7NRNzcPmDcf
UCEBeAqntzkeN+MsYiw7BDowocuIcR9C9+bm3zWd+jFmqfNOEo/dwoXajiz7
QRiesp9QROrRD9nLkK3SQR1fWNIKvRhxxRx01NTC4AUv4IkycfPDN1tpdg9u
H52VCf3nu8DhP+5zb4lACIRglsmvJmKm61ocOz578zRTEtN+rxth3qQpQCEU
2vQPg/lvCDjBnXU/Co+2D4gX8MyVryhtbJNzD9k8olx6Q6BapQo1+jtgF+Ub
QrY+FOXUkfFQBV/kuAXpyo7Q0KlRyQpy54CLPq69MjrmTVHQPmQ7B1VMEokd
iXCd1mf+putbwwPlkKmEfPk2vnJQRueVVeHoMcBiZnCvSPLYbG/WeuMyNHgq
naUk/TbH6Vv6j8vXLELoRvjky6JVGx0f8DMrpjxDYaB33msCiKJwOAGldtEA
9uqNq7d2rBtejrJgHA3sawQ7eZW6w1XVT3yTyqxIH/riBOvvgIQRJHIK/x+I
ImNo6TWrXjhHB/XbXBNN0w0OCBcAEYLhWdYEYJ2A/z1vV+8lZfrc0RND6sKd
LiiWtFlfBqUI08a4mKpb3b+yt6cENrISn0l/hXsm2B9/NCsxz8E7Hi5s4i9m
7hfitXQl9MFiMTFdDJctDE7Kp5PGT1pcLmCIx6XkG/YykMzdfk8uxyK2OVlI
4tYzxzqRBm1vt7Gg4W2gvnxXyTQ1TeU3Q0Jn6EfQmgQqT3SZbw/GMO3QPYaQ
oCLmRC+s6Yj9WdGO5zuG9W7sT0+VPxx5NNE4GMgMdFu5AyRVhjT2mI83HdGF
Werg5fRxhZICd06vKxKHtR8uwvfH0WxQGH6SosDhFOPmMazGPD4YZc940zJ3
5dI1V8qet41u0fG1+fUbfLWT2ToRTGcJDl7LoiJa4VFc4JhS2FhZwzHv5699
KEqMk35sdVQRSBLXsYD47S4T8DybH9gUU+bwk87UGXGkVigjE/yna71mCGw9
Jiv1eefo3t68KtH/d5rH4qGhXAZLn/wWsFoWuPKEvqiZA78O2n+77a6ndNMN
CTG5Nib9gF73ktbhNUHRuqc0lTX7ZKUiYtphcEhQut2wMQ9RXb18BUW9Nx6E
ev2LtuAwNi69de3+nCk/IPeE8208fk1sKIMm4rY0P5UY3xFgiZRsGPZJTP68
X4HSZKVSo+mW7O5/OrWxmJX3WFg9+5pamqw0y+y+6Hu+fWb2GaHZPu0RFScq
UR0S22yNyGk94xNAmIYHEIo/igYROKuLV6WZVX0r7YJuHkgGJj8zE7s9AvPP
RhRE7ZgniE9WklSZRweEhFxBGLBB0I17RXw70OJG3D+UHyTzynQ3dj45xjvD
tD1soI2vQlB4Lk78/Ncul/LPzQ5uDkyETqgwpPQKFeTJzLSA36mCQunIf8fT
arKMli+OxAgHYv3D1WiLilXwVT8A4n0+ShSo7nAPxivt8qZA9ckAJ7a1G4Cx
BMUVYQ8IMdMgH0qsePp/1XGE8OEbzTTbkOYcFGbzaphxAXrIuhUt1/a3hf9H
XQlf1Z9MWmTN9TaWI7AWu4i8nOn5eiirV6M2q3c6qOSCXutpBBgtXBWRdFWF
/qbVY+peeekESC71YpeN/EkE8tKiQzxVxVntbpuqE/uh5lZzZMZh5am3Y9R0
lJDd/wt0CmW5J7HtZVv/xR5mlj2ngz+xD3DTua7AYR9OoIuS+35dcjvDLX0i
Njw3YqMCIU6e3ABuLyTYqbAVp6PKB2/JN9b2rC+1cDQSOS8YVNYWuICzECwj
ES7w0bAdxZg7EvuhlHxfNQD8Yg3Tnfzn0iumBixVU2QbpqEeVIVpiJ0rMQln
Y0ZpzukHpfnIWlUXDe6hxCR7srGR8qBe5GW2m6Wy9UXR2z6gxOWEY3XL7zqs
qw7QzpEPwxTX/7/WC/CXc2pU0CkNKaTks9F4wyJjPu5sLBVjZCUYGk4P+Ogj
bWV0yPIhLYYEu+pgr76IBP/XfeyiZD+xEAWeJ2FqkFGkrckM4eVo5d0l5wQr
Br+8MXpvihCIWgN9qGnr+aS83z7HoZs/DL7eqeVIeLpit4wQKVM7Bfr5wx7Q
1KksJtxBgBLwtoANPTEeoQTOxwgrhj2mBM12iuCsZwxl78lpm+U9sS8Rg/nj
JUhdy2F8TmVh/ooEVEMNYa6rAh5r0Rp1p0OOsHHlAqrec+0YNRkS7L93SlcT
u5MSj649Zq35ZUD9IHZedmJO0qrsxCeWW8Hj5a+toNGHoLOi4sT5mspu4niI
yitGtWyONAhwKUwNHeWPo464JGBBBBU6eB2AbhIRrOmKxhPSKrdQWOX7zL8t
lC7E9jOnaUjO2fIKLRmdygi4+fyTeaCA1yWtVqqNqiASm6BoN/Nr8NMtudTx
pDB7XG2V9RzlULYBtEy0V3fnqmlfeSmmazhTRza5PqBhgyE1V1YlrTLw5Tqa
gsKyYEv8MAakgHtRGs1QLBo0i82BaUIrRF/anemWXe6JukCSxyQlpj0MEPjq
Iq35P3OlPRrUaOx04LNczldtZHHXTVOiI+K/fTVTBR+ryh2A6QBCycxJzS+S
T8m0sIVByqoahi1yNVsO1+jaAv+kv7amvfzEFuawzvN1DRylhhh57sLTCjeN
c1iO2nzfxwZPiFnq86gMR/CDQWua64Cw3PSQjHlxMoKLnWqzK4GydlIn8FgP
66F7y2bo2UBuN0Lp2Hoy/teqEqaTHfo2Q96+jX+GCvduRukj2msM+K1xgzKL
iNHAIWQAvfSQYG/0FZ3cAdww9ozDi1HTLHFMd57RxfMeVHShCgkmKhqH8sCf
BtJmKSLOwJ/7w0ujLGIvYo7sRBWdI12VFoGaAPacsvB3XMdbNzNY0mXjBGge
xIper+Mv3F0/NfUBnbEjGtF4V/94VHXIZ9rFd4BZt05TTp9U2pcGlRPkHl0F
MfN3OqFG3PhrkQqgGBEPmN9MJhsgqAoiw0xgYbTk1q0aGf6sii8L/gNVvC8j
SnTu9+1NTNy8R/sM980nX8aT2/+MgiylFVITJ5Z8tGoOBxbSivOE3xFQFmPl
ToJ2rHiFMbACjdrrBYjuv1RhcDUPni+5+5EOUVrScKzRGkOShjkFnf9y1e/3
/VJwJy56FXKAm3dB28SQLhEYcjxeYtUwViR/XVMo51CUAs4ztYOdZW8rfYD5
rybhlheutkSHj+ZA1CrpX0wdQPmCt2F8cnaqqdSgmsNWpUZ52z3ZuTt9iCBz
+Jg7bR8nH3bcvtfqeKnI0SVZA0HlKy/Z/8c6ToRTRO1QKwrYx2ignviWvGXq
8a5z48ZfQXcO21chil7DHb+ZqQoZNVH4opMgbVEj64EqQSRUTuesfcB8t/an
1C/GSHyO5rmLTvW0WlvXYXgc4kbuuaGx1EwUj12gQSSvVaTWQAmZuo3uqy85
d2HIyEquK0YNbRtsPBCINaYIj1g+J0tFsWKU6wqQgYmLxswZIuaQgyd6KNOe
qF/bH2mWbL3IG2hGEFvmZ6mXJs9QQR2plEAWFtk7SuU1oT/Q90DeXm9pJzxa
NOaO33zgmS6SKgAY4vnbVDt7/WBXJQtZKwI9ObT6TgtZ3tRKm+t4AsxFTRhg
ftTmDB+5RE0XYlTF00IutZgPP5hLYH5ryYuvTLNSBV5PqIb15iDAsQJwZa88
0fWagTQCLsH0HtCv1ZZKEv98AwINrTd4yVbkrExixz7cPxlc6Aksx7v4ejZL
gza3dubPhSWZueu6UYLMrl89OZLqH92aPNIWubQNh5pGSuiJ9Zp3J32xFKLK
rTwoi9RCcimMnJENrYDWf+YnZpqq5AVJciaDB2hjNynVulRGezZ1eBzCvr5+
uK45Ai6zTjah7pSIYqvdpAf/LEZuGkmxqyyQBtcoEM05cg/zpJ1NY7S3N2Vm
qzBQDaTjpGQZ7myyolqdc1W+9lreBd+wOxTZxs6Ih8QI+Z3KX0l4zxFYbgUF
BZ2mC2vSLM43nyiWuJWy0Tu5kf/dn2769vHcXSpY76ebKyjRJPFLF7T6dDjo
Tub0/rQLzhjtyPcxZV8nQH5OT6kN4zKmr4ZkPAp6zfX/+Q4n15CwrQlKxkSF
kinR7VfptjUk63AQsePcfv8zqzKwf1nQe6ot0LAmHqvnWKIrey5O2SlEyuhb
Q7n/vw9EL5iu59i6TQcwf5B+9q3mbrH++4JhbKKJ9xQaDZEDjN2vRcKfeEMh
aA/WYbwt/GwwBxj0hppSG4d3ymfHFE/7DaPJzh+rFdVZ2krMsdFliKjvChW6
q+r7eU7z9DZ+pml6I8/QwZrKv+O7hGWUUgFzUP7Er+023Rxj3igQrvsQ1et/
Diaz9k8SbIhrlSzfLh0xMouQL2EriEyYuxmp2eUeQSk5Nw7S97qvuOP+9gyF
JEYp0WfLKdKdX6kafcKEMZRSvGTim76dvg5KyiCXrRgA9DZc2FET5h0m79tg
g4aYpxmN7nAjOE8WvuCTuTpOlBNY5UIoEwOxeQWGaYfh9yiCKFJEqru8LW0I
RhxCT7bzCF8dHEHUPSYWbtOK8lPBAs4O+Lg7VW3JGLQJPEccB4GfriI0gCFG
tIBDnC3yqy+JGMLiP7fDooHBh/yqCUJoZPUcjTm0nuRhgPAwyTCap894469t
fKsXNRYrEpN1XTGDdBzDjEaotFdsMYfKp5lSz6TmFF9ZjW4vw/mY2Yf/OoZx
yMj3BzSN0wNNavqbkdX50kYZ2ZrletoumZBf5MLzm7ZhCFV8zyxB+57aeA8D
wSg415Efw99SeT7iPcJUncJn2Sew9/ZPvWr/9TTtcg/E/l8ZIkhcHu1z6t0n
xgzVHfPfrknJoqDt0X53WX8DYU9Q7uYilAGDa63+d8/E9WqlR0u0ocM7+n4s
GFCzCjVgOzIckW/Ydh9EmKZ1BLqPUqCq9izVNkl3qc3ULVwxAmRraT1p7t7x
l9U8otR4rD36mDwTHhgHKK3WDgWqbOxVHiW6IlSuIfeYeQEtIBi7amskF3Zd
jgPRF7DGXgruC37FjQ/Af376OOQ/+gfmK1zR7GYJCWyQxu9xH0pKBmBB8JHy
rg/OWLSmXqjfKaF6eUQYXbON3O690mO0DYS+6K0uipwUPvNuSSJKAbahRUgf
L78ETZJFymZvIgJ82+x1KPyOSk2Ed/LXJAt69l+iNMLsYX9+6T/KQtTyCGP8
jlgLrNmhbHAsKDJ9rSrg8TUuynMAW6VZJRTW6jwbNYKQK85GkUq/kkqN3qnv
/WCKQmRnFU11j3M/BqkzSJwXKsztVBbf5hN8xrFRSaayRBrC06DWopf/0MNp
HH9yIS8MG1axIK0T620by8sQy2+iYXiXM7R7tJZbyWtnHzHWs5Rk7gZcbTDG
kNISJRQCWf3eplrU2+ZnDx9yz5YomN8bO2kzcqtLccLSTjfNEpNINNSHhvNs
4eIP7dkQHOi55ozCBbjskdog1n7emtS6MoqUcKdPQJs/x5yc/i0eFigX/ous
s0pfZJKx9uwdgZQI+uzFqXNgwGm77pwGjqWJY5Ia36mk6UCzbxQw2vXB9wct
DXfcBytiPrj9th5iJzHuqJzuKrbGcla1Prp63uymKB+7LoD9WYjinPBKPAep
xzjpqAaothNepa6EYP/bZn4AY2XiERK7EK+Xw216046fbbqFZHpBzSC9e37u
7eJfWur3xLinUz6Hx75T0ktgRs/794i6WokkquLMJiIDpo4iwxw0yiidfx6a
3EBuj4VTy/y/SIlFf2gm8MF4bgTb3jhWkE7HQaK08zBWjtSpoDpV8hkNpxvQ
xdeFZexQ0wASwZv7enVXkt+1FZWqSNc0i1WOISWFqDorkcI6dUH+O9ir7MYv
iV/A44AcZIL2OyEeUq3K9vUrS3nwparXbk2NnuPQQPiNkoA2s/8mukgYRo+3
ks46V142lJiLkqH3C6a6CclYDns6qdTC4SzLCjLSQhMOHAw1Q4GmmQOo8+Gs
1vyR6xGLi3h6yyeIZZcXUb7Ka+0+ahDsIYjP3SQS2CH4rp28ZVsrbqrRFj2G
DnpbPZ4/geDq35KLDmIB1Dw4PfFmEoY4ipbuGBqM3e9IXcsQux4GBuO2dcky
2OmLggnu7LmIO7xhfDSH9HcBmv3XVP2UVQyUY25Qx5mSOkY1JcEDvE+DWQFW
o9zCES9cPO4xEDdfsPAupzX/7447ItA7VnEW2BbFqc9MXXgUgR1o2eK1s0cf
hlSM+uEjvViCzOLB0+NQ1LPdixRRFuIHHTNOcMZRilBAamdFr0ViytDEahRt
kC7HRkSrT5pFiJYSX1BIDrSicgSZ1h/szxjowQZP5QbslJ+vPO+olxmzw9AG
q9eCIHIXOxL2IVLLxtXQtgwnCObnGdrmTMHfR2BhEBpR2sub57iDtYnyQmCu
/MDrfN8mD2SfnBfgrfmtyCqqRR2iQBglYZ+pYwoPzyplkfYHnjXTY7TNbjOP
X7KLjItX6hyYRUfiO/kJH7LxObYWqLKSQ+8fKbowwJYfJO2qxgu2BzZAJ6C4
UHX/bbz6+h7ZqsnmT1m7UrxrwTJDycf65ysZPPv0uWqSKBCZoJkTOGVnQodK
egVPtShZ+EoZCcWpmRx7LpubG+3DgXmlzORsYNKuXhNwkFblfgsAjck+eOFo
u3JaX11wlCNpyVSfIvKckm7HLMQgft2likXl3Dh/zFJKQm3LVq2okDj0fMJG
+IYSCxTjYYUmuFdRKgAfMLH3wEnY2a8lk3LLU7JZtJTaR+iX3gHh9WZNaWrn
VvMer5aMuOkAuNZp2XNI8QZdrlslbMUG+mN7F6nQOilhtEsA9EzrxJZ4gzz7
6x7z1KGFuaVdp5zFLr/JAWBiMWRiofYJS+nDk5bwQgJNsC3Aw2HY5wopphKX
Sbcz64f1JdEl4N8OYNpQnsXCJklEo4YCqfwoO8VLwGH+hoO6McQMQQQ7E8eA
QDmngtliP5k5JSDxMUD5KWCur5PgjwVUD62sGkjKQcmoKS55cfIDJtpC6NJX
EMUBF/VyajeZ1JORq8r47EtsntC0PqNlk39zfXv2a/mBnSjswc3f9KMEELkP
58prUpkimNywK5xtdAMnO9Rhd2KeK//dNl43RXin1GDQyubh96PJQoe6bfr9
vxLUZNgwllkHIp7leH/6ucz/WaJhk+irlL6wGy3xRuMQohvDoOonjoRI1NbQ
nCuIrMFIdiWjnbrP3AR91diQKRN86SwKxQJJsKFd0DlFf0Q2Jws6sWnmgt65
kyp/COqlgzmGbuDWrSnDuRxTkSMwTHJz77ZOX5iUAYwzelvjcaEYYE/V4nJJ
HwiGuEmV6e+PXjpvkUd0VYJi/teBsbcCPLQZBJERxI4JQTTNkbf1psGad+eJ
2yJfMCJu0n2HmmPJ6dBMd0ufYVJShQBAjy2B6bHregRXWaDvEGNRrXRldKga
TO7EtXdFvfIP+YtNSRMLjUXSV05fcrFlx3RXHacLJ8Dlug7zRl/8FTXPj1yA
6k9F+UShciL39Wc4mT4l0ucLnGWV7cL8iI7J5cHqWaQWVQ/651QDjWge84w2
pkoZC2OlrpNVshwEN1UVPf2fF3nKhuRQUO+o5PHjdiBZmbeun4l+dgWD46pN
Jlq8aSTmHxiS2ExJDt10jFs9tbBpoozRMkD8TtCFdrFYwjXrPIEnPfTZp7FM
K5PvbX47FCJNEgDD5OAAUuHTaN33eaEkd2DFjUUl55/CpMI5mfYzxJkVS47s
vB+R7h7I08wWERYQoOnQwKHOYYPlDXY+OGKCw0qHvvXqy90ZujrrqFHzx55U
ZaaZmEbi4AXZ5VbNM410h9P/JOP8q59JKC27EYmCA4RR74nf5dD2l9Yi29FS
q/zqEDCiWrfyqkhiH1XHXuzliCOTnOi1vv6byqX6UTvfr4wc7VHxQO6hXoDP
WrcZ00CRAzoDfb1kPvrggtTjVl5NZT2xE/vV2hG0KDLU08pVnF3WUkXzWs5T
qOKHrtXaVDT7lmvB7p5moj1iuk7MhuIWi0O2H3ItppAUPUiRHjPegcgd+s+Z
1gCELZ0z1qJv3Rbs9ALrhbeVIw1q4z2tB5lcl1NVDqRHgHWMeOV+iZL2dMMU
ealv6t7ZhsDjMKj8Vy87m4Wf96pJsNWqXGrEt2a5VM1SEM7vva7UODKoZF93
2k/ZlCvgBJQdCDBwm3uiCDzYr4cXPPL04TxdyBk7JbGyHrUfX3YKz6BDC6+f
2+Sg5nYRAoQJMrmQRLn0+MP+vEgPE2LdopGnVf3YRepuhJDz2W2x7d4hTmf5
FUzL/zygVDHCeNleBH50CkRv05mAe7CXkTBC88bYagbKsQs2PhkJBHCl7Q63
p5EGpH6wvR6lwXuL2PCYmjderGMo3qjaBuM9tQNexpY7nEmt+rNBy0t6e3+m
ZbNQg+kQi0d8ah5S3fKAwaygqtnrsvG6gypxPK1BTMAt3DMeVi8eRkDrMJQo
8gEXyIVCc9RcVH/Wt3XVBzR6307EiYmvXghAOFio0o9GuKy8GjPxxOE9VbGz
6hA/p++bbTh6ADi2ue5l1I9HuNEUj5s3gMOC2rbzGaY3PlmTMbFA0C5sVnq/
S3TtNMm8jTQCCFJXrFlLnbsLcS+gRD+eCciVzvjn17UdiQ7Z2s2hJU5RXj3A
ryV69/ntsklox+OSMC5JWP2Hcmyj5xna2Srh7+CfhTcwWIw8Nnm7l43m0Sjh
02LMricotssG7jmoZ4H/JJzxV297Fsfd7y92DOpNPSVgAMv7wWQtKIksYLdm
BE+VZ1g95JhZY2n0ceF9/qL9zf645O+ikdpQNu7Eomrx30CflOvZA6pUwmi3
YybzbtI/P3FF77QFcmIgVqVdBGUjBlqfWK5b5SjKFJsctrGWhJoxQPbfHv3y
1OIgXI26mkO9Hs481TKHjQAd4NjghF804RxHbupDAPGIxvyKQwAlUKFVb3ZH
xVUMKrJHi0aesDUAEN/pv9fUHmpwELm4HwHmG4Qgq2LM9RVMW6vjaVifS7j3
hAxcQ4OTiSP94QLQfQe8Wm2m3G3t10sPOUptZZ6K14ve+9smwI2MB4wNh7Ua
PNTRCQ9hp9FyUWrkEZK+tF7tI1YByGwSURpn/h9HLGkzBBS3FXXLWoyI8Vqm
hx7WxLDZq3Sfn2xYrx1Q0jsCB4XwOH5iTvAXLgU/k9Fi5mcNVkgyLZynrUul
yW63FBVVNAfjcDIlVcRErZl8aXFvytdyucn6ywagJT19K7JC+yyXO34gNYjT
uKiBKKJJw/jiiVKpUiQ6GUbxEj8NvdDoR+1hSUEnsEL8Z7ea1yGgw9pW1nkZ
hDTDLpgRvF+gBLLjRYxQw760mdRY6a/q+ZmjQKt6IxzOBEtyinAjp40cTIzw
LIz017TQmEJ04o0VXUPU8BPzEEmtS8lvX9lEtCVExY43SzOOpP3JI4VJmPfj
BsQy58GujhmMGVAA7emlMfLsa8lIbcWzHqgTsyptKlqNXsd9xzn7ndNuqGv6
pim+DeVA6rfulOoPLlqijKd334umm1EXNQM+wgFR+pkN+0cnyxNvzK72uT7L
Kp7unjhNVS47B3YUpR1Rxpqn9TidftQF35l+PepJ4kjqYP+PxnpZXXPaZDRI
5HQobiOa22ONccVMk4aH9K2ppWlfG5zarZ7uhyJ+9bpZx30hMzcHgXWITgZl
tBl1nM2t728WmV5JDRxjdFpZcq9xqESyNrcQMH3qH2UrGd4ArFk6bccHp1z9
62+0AUAouXjz1dJreF7owJBuENu9Whp1v3H7NrG+RWOg23vvj7MNIFtzxAqI
PUtU41PYr5VGQyTsiNZBQMM5QWIy4HXqXrNjSw+08g5OoYs/97SsNB54LKtE
jCTsJjxSVHYhNdNNMwC/DJNUaE4WR9cltKENAPZquuEZ0OGa6uyS6o7UqpED
rrNbbNubtS0Tbou5uVud16gaO9oMFWtYuPexq3qIUzbnftSZZvMZKgZtOnx0
SYEjRI/9kD9WIiZyZHeh02QTPIYOLrzFgz53fjb44fr3Q7SHj5SHV15RDhvn
L5tuGPaAVrDEgLCXd2JcGCVdNd46ma3bdbUduxrXcRQccV1Zv1SnXwdkxMX4
yfFlGRwNmNNqn0s6pjPAzzLoaNlbhY7uchEh4jHRDkFl3QnujAcKGVI8JXNn
slZTBXGTGVvIvTrfBvLOiC0prkDVpnxmzRnTQHYFmdQS7XL7eTDO9XdEWQHZ
YnJNlO/dT52/Gq4smdEAeQRopLm4GF7rWAYcFHyYc75qIj7lA3fU6xcECS+p
jmKrvj36gdNlFa9BPfFqJzbUa4Py0Slbk6F4DT3YN+SfR/SxTRN2nPt2VB1g
EEQpqQh7xxdSTAWb2t28ukF2s9ZjgpNPwnd/AzPoOpg/B+gG5JxRSiSvdHcY
uLAS1OmEyuODYdSxWvxgpEj2luEJf4O/hqjQQDIFIzJjuwxbQuzgjCwePXgk
VIZ1579b+dzbQjLujehN9RK0+/o3sKRMCh6lZWo8Tu7T4Euv84VZeZSLVJY/
RE1XZnkRiqz044ahFp3Vi/EqUocsr716Wzk6oYvisRvLVk71rz/qiat0ORpU
yvPXMfsAr0QCHxQl+Y4DKJgPS278N9bGoBDWAUZKSdfH7FfJxYdGmgGzNc2D
xOo2OXIbxp6yuaESEFWxZp1LZsopk0jc/Ygnvh4d20rqhTSGkT03N7ncfjuy
W7/iWfEaN7CMzn97aUL5C93dEYYPN5EpbQ+URhfJcu+w/MECauF8xvj/txTh
z8mtMJVTLZMalBYukzFhFlf+ue7X6M2mjNjQlipzVXHi0MkTqmGfAf6/yTpE
ZL4LqLA1Bzpv6HyVGfIyo3jdzgXRYbOMAoc3fvVtmChcjlTC4PIlRtUcqhPE
IkXG9RuIyfikhFPXVe7roeNFHdg9tcbOK7hWynHyMAI1NYSb+NaOscA1X1YR
OijP4iUXDpkXG8PjTwLetXo011BG7KWUlaBCytBXpPvv8+imhP6kueacq+mu
X+Wmioo/Cr6GReVzMjEStliC+uLTp8h2O5qOXokNU/R4PY1y5CDLukx1zsG/
9L2HmUYYGL+mCL8AeouHmJcob4FYlCFbVWUKcCTi4nWe9sW5auRit7I2fk4v
azUgkLyY8/dq0p/VeNdhnFf2IvJkzA88MRY18z3AuZkDPXPp0sKBqT0WdHrs
2bqgfusV+hxM/x1xnl8FfMlpxMpapvGn/nqE0xQ4uMwlQcqmmceaFTv2Ozwi
t3iZQ0xecFWxjwVauwK3Lo/rr6ZMZlhlZ8AMTgZzUWhl4NPrVLb0NecHduJe
iQSe90VaSQ4FNzCjITMJsJOhHJg8FhSy6iyQowKcyOmyLiUTPFrm/BMHzLqb
H3ZoUBmfk740NkjTrSv75Sab1Gam5dUE+aCccnTijsmkKAesEpaDfUY7YUPz
LYmspfvwzoMSLg1arppsOWCwpuHLueJ7/VBQprZ47E9cdHZHTynd9stT/YvL
rxFotO7z9hqdUkGTrK/s6DzRh1YRxav5f0S3Okuezn6VjkTt4HN4FROjMmRJ
mvJs/tmO0I+S2gpMkBL1S8ZIfTyFIe6axKkHw/hFZdN/27XW4AEHt0wr1wN4
0op/2L4md4fBdL1B4AkqXF/C2FUkCfqLAL+5KTyfx0GrsTLYNH/y1R0d6gbX
JnbPVPjTdsUUoGKXJEEk3Eno7C0j+41LSkjHwTGas/jrzpN3VJhvfWMebION
j325Dg/vR6nGHRhTjYstYEC6lReBH4Oi+nO9urNctmKFJvS6UWfIvTpOtNZK
WavJJzKXPqT94Df9qIHtgz9Bv6n/pBnYTECRXdEyN8+BzDW+0CsOOpkTTHCh
ujonnGHUaYtpIjvVuRzcFGYNKXpF55Zx9Yq3uYZV8VlZGSom/7C6raltg7lR
O7XqLfmqKNcFdSWaYi59VB1Aad18CrknQfejCyKg/dSquRmO50Uqg3e2ajBy
WqWxEmLJ6E700An+N58g1ALsHIsDdOalGC6pooGuO85uMlPnpeqqsNSvIEvL
5RlDuZGF6AqxSlpaIXh6L+CYlajdXLybdDpoeVcL9jjgG0pfLLvMacPxGnAZ
LL+y/Sdt3xRDO0g6ZovO/4QM9lbcdMax2659+l3ZSqC9hkR8wwHy6A/k4H/Q
PMS29xi+AjY+tXc6fSI/5RXcU0lNidiNR3qatfqvcypN7mipIia7RJr2Saqt
xMESkt7mad+G+m+swTxWPl1Gcdvx3J07Q4GBtkwPA2FYPvX8Tr0okeKT6j7z
Gmgp+re2+xr6AI67TgwPeO+RCq3PkKaKh8/42U9bTYW9jNcgkqSL+m+e95tQ
yzVnEwGyt8CPQokSED5GVowKJzWXwsMg0iFrpdEUcv2eCywp6Uk39cEoJ8Qz
njmALOZK0o5WlX8xyGtOa7zNW+JVQjtyszPy8wSJe6mXMhw9UxhbZAvdQwIA
yknrgErl012H0Aa3ammxt2JuKub+VuWAZb2mHoASQsVZX+xDGlITimlsukkA
Ptbb7aB/Fs097Iw5APx0+9w9YGiXdnMGb9AkJmyl/MSIHktrQ/n/RV3QgFlX
OtbJKJUB5/pihwWONxWabrBXTf5DIoXq9BgnGDrc//C+cILGXZOQDnU9bZiE
bjVBQ6xkiq84vMlE/dgn8eQDFFOsJWkHSsz1hPJY1filiUDCme+VRLVMYhRM
U6YplvMiM/TSAj7ZDRrkFq3gDgpq6jEvY5WrPz49yQ5hjtSKXY9dti05ydJ2
wDMLMJQEl+o1Yq9Wnn2K671/JndrQIRq4WU9Rq9UJoqUrrne7xDRZLNEp0yS
sdqutU3YgedKdPg/mc4I/VZf/3Anl0dPW1lrVze2tdeZGEy8W7X8is6zqoHM
w6/iINe9k9POYNIjKUCRll49nMS25UJGjLonDq/dipoc8PYYKy19CQsK1hnv
cpzR1IkbA3k7XITILp0UB84ejdbZ2LcOMuyNuHkqHkuPP4cHYXrbiaNH/4Wi
YBbQPlp88NJepenPmGKaebXplF+pdgFakLZdsmvuhalVQUKnZ9qWeUIfPkw/
PbgNU3TZvOUkoLLDrrgNo9B8t/ojv108tT22iABPN1z8cX1dFzDAD9kaaKIh
1+Bgn4fmFXRNNxazdnYJX1kqlgyCgjywhYaz5gxFfWZUl39PLO7fgPYAj+vA
Q22adj6JUSK8bZEbNL90CW8dyvoc8i2iq0EAk+iS/LMMGbtaps12kTawQlxs
G2fReyt2qr3bAsXjz5gCewl94UmBzdtregV7p4CMMLlf5upQ+NeBsk09bpW/
VMFBuubBJctXeDscxW0VE82d8k5igNs7Soo1NP6uG7OUAFPufVALWCAXjzqM
4rOkVNS2vcUsWrkFBEovDo/eBNvbJ/TrznYgHeRV8NudVKIzh71W53F5ol22
Mno6iErM0aaZlHRsFe4SBFdP0vPzo9iYWLn8Ze0XSATtLKkgmL49T7USTG9c
hryWTbqiboCtWMwTrFiPNptZYEdVSwb9TU1RGi+Xknu2WwvfR5YkKzM6oPMO
KeBX5OksBKZCDa8p+4cwP8wA4E5AXyyz9uUt6ExAPWbyzEMusosdqJswFP3e
i3klRF1NVbu5Pon3BhMB/TEd8uUeWHUlM+Lrdzgis0WJM8borD77YOS8EUrh
czOIQojulff9EgNIQmlrD0UvZEAkeRhUQVPcjPO33jnpGmEy+SYjKt0Casfu
IRewEeiMxc/PU+Hj4jl8fe4/32LTiWh1bN6hL/soGConydxfvYY+WmWWFXXT
Ml6S67eLZiyOAdMr5hj8aNREbzWU97A72wiCepzmDrvHN1AkfCTrnSXPPIeS
HIrLbM//WhZdwJcPfpfdmNUuO8DE/G2+K834vR0l7I4GW/pUTpm4dZXYbBMg
nZYw48K3FzKTNMUB1SeLAYt9pngYIh/iN6t99epxvaCRcZoT0Yuh/BAjppuq
E9cFT8Mzllf/jqnANmexHwxkaKndCYGDrAHf4K13enZKcuqUC+WXwDcOfOXg
34Yysx0Qof7k4b26hy5p5F9mTUFfpR9FZDPT6fgaukNlwWEg3OPb3q7yY9vR
HGI9DK3e1gkfFcp4xon4OoA6TP8N68csxsmxeLGTHjjPbhaqiLyzk5l0pMus
EDsNlSDiq962bi1ZYs2MGHNscpZT13wci2MV6x7z2N2DrCps6TlmtAZPEFFV
nviEWa3mRBTG5bcZ3RbiBWMkOu6MbP4sNi6kc05AuB59ltzCgDZTv7t9wvxF
5J0tV8SfUH/sIPvS5L/ASc3oJbBlfOXeKq6weFvYoHtv7yIKfx0dVN6QlK2h
lP0yEo0Ghpz0A32/VDOR4hzOQZr1RwZD5zq9VcAf+uXTxxJ8VhL4tpBRLtlZ
fix/xQSLmUuwvPEwGFuw7atd1kfIIIOmd93Ve7JEwg2rEQWNcf7jWNartztY
1uOpIOT+zuoTgRLsevkodO3DaielS3bjZIeNAMo40TBFphOGlFF1uHE1tvbt
AMrvNECBtPKd7sTi8b/yX1EZJ1xtz72rzJITWh7MKF1iCDYs17RFUkn+Sln0
Xfs2ogaYLl1m8fcLiSvgUhtVcDAjFmCRHwFVGc+A5oqi10aBgie0/ghBtTel
F01j4IbGR8a00+JocFj09MFdB65MFh+NRbymD1zSkK59q0IhGR0ceRrh3WrL
B5Yap0WZVvV+95BUnCDV5eZ0NX/YFaPU9TQojNgMdsSdxg12Fucs8M5NW/T7
wDps8fSsfF02CdvvZ7+Yv88cC5RdcNx4JQDhcIJyjZ5s/vQHWUY5W1XYLVhk
PUn8wv1QcjjFPXQWs7qXfJF9qmhk1LnAWZsAnURbKgZTPdz1UPCG0CaJqPc6
WtzUjrkQguB2BKXxXF2b/0F41eMyn61kVQk5vPCjjtctXPU9a/6Yz4gIjvWG
QQYzGuW2UoaG9bPikEI6sOYVGOj2BB675f5pwq5suLgS2nEanjK6xtLCdHqX
44sHb6q7n2nmm0Kp3Pa3Jsy7HjZ86NSj3oHqcmYbt3dre9t/DYadxHgOIdJI
+OndwIKw7zxdVR9UcKgqwCUJnZB+YSTRUR8vP9U/y8WUybZtZGdT2tAOW5t1
PLW+XbJWuZz2uctFvDGOSMwp9GXwchEUGmwId+txdA2F93s9zg4DM8BwEmoW
aNZMAgu4cow7m7dJ6529PkqaEE0n0t+nsX9S//viNAyo/mf3b9pNIZszsQ8L
RVrCNmM84gLEdWYzHVw0UX1jEytfgoBezRc4t104V2LP05kguJ6hSN1zj0U+
zT1TNhAnpvCzOAEQs50Mh+Zd8/J7kgEF+AdMYzHUlB1U3yHCLiJGSMwOcjf9
XO0BAjKXVwS74jL1wfY8ZvCG7jA3DPNcGZ0NM4GyUP6qakAZ/fKBLR5HU4Kh
ctNBOs+bQtUhxPtXYgwEHQf5DmK8S+d60TcbmCDvRgbPVX7BdZn6YHSLoWN6
nEjMJ5m6CufpKZ6C2rQJKLkuOSCf35h3acXGCgjDQGiOIfM2JhpBXfyv9Wj3
VUvKf8U8xBQetpWRjVMbMnFtlx3NLG5jZ6G05F9qOdcWF0pAfnRJU34wL6E/
8EMpdWwf39L56x7ZCJQLovbZxll3gPeZMsLkQAwakIugFUZIn9c6JKTJAlTu
itq49mR8ifiOSrIq3gRCEOF9+5FZdQm/aTnYINXUVf0owMS1B1MWEnuvemI+
WtxHaWhrLlocQ1lKDbq8QyOFxXZm301ty55FHzcVPYYWshbrnMkhmvCszoNO
6MJZDBu5vHiOoY1ituzuFcTAxhR5A/ErxHTgcDeYU5ESwtOzQCuGy9RVpKJL
hkJFgBqjS1JboEanNBnwDewIgd9z5fyF5n3fV50HhyL9cBd2I43yYr2lbNBu
DAMIywr6FcnIRb5Gn7322FQ4uOdt6/MBLnifNZg6tV74et8cETMA/ZJZ7gzo
2NThyBkE7wUNZpMGD9dkKHI7g9QHGCE75f5+YkBNv3z4xSt7SwqxOAD10M6B
VDPrsNRAMBXkIp9wlgiDpySg3aQQ08gelnQnFO7SA6BVMWwrASZsoRX+xo17
hAb5hAU68ms+QCe5vjJr8bEp6eh6fzsapLxVcQs+vGYPbO+LiT+exFI1Ols8
VxPP1cSjH4wjGCdWJmARJsybwVEgfaOmWVqjRaqopZ+hciXe6rNm0hyyzO7d
/27JNq3IasC2csnUZY2m9B4mD6m8zwBDjmGAMh6hdxviDlyMzYcKmVygSBnu
gCClId4aByfziZqr8n4jJMnZKH7paEiEk4osL4KK2MVJFS49CjUJYCqG+3o0
mzQl8qkYAfJsxj/9YEgmXjTg8z1Wo39MsmSlockzvxwJMCgiamoqKoOugNCr
/X6puMOgx8Vxb93Lm/A8/m2U/SAhKSEn1x3Czga6kesaAWMUo8KbDbvwhoTy
dglF8LAxOV8ZeO8so/Azca8N4J/xlyRrXZIRrufv/jy0J3Ifosd/SNTPlKKI
71r8Olydr2dl/eYLuTSDM3svpjE/ondeV9A+zS7YkFxHHC+E3WoSto/0vcRs
vxT8j7KWVmL2+Icl2auv9nhV8JUxr0zECQWiYD6IXpZ6zNeiMfJ+3i3Mazw/
mZE+MRzS0izz0Ylj92C4CM16ZZqIlqKW4Hns88LG9ghQq3s9u6hGU7iNt4TN
IU21Qn04bUCR2hmPNnTO3ePzkL4oPQyrc5dwlThnMC5hMTk2Vw1m9xMD3uuq
LckFzOpTcvingHwTX0R5VSw6QmKkjYoiZf6IZWTeL/QrB6n/V8n6pJJfT+E6
Sqpt7XoV2TXxf2fJLI0qV8qCcZ5cTu1wvoWOlbCqhVIcyP9kvyKE1PSJiweo
lLhnTUdC77YQHVpYD/SaazV9o/Gzcdh7Immct57CdGn30p0S/UB89cqVsWNr
zKgQ1LfEW3mHCPpoFCTyMV20cDPE+OcOFxQBT9KJ/Iu4JJgvzE/ujNvK3+gl
XvnY0TmW4q7Wj+zedQFmd5l6QrHDcQcgFkBkHWttLzF5aoGYnXExsZ06DxNM
SMl36+HFez1bN+BAfia2n3msnSL6m5TnHVQFuwZyd7fm2Ud4M1ULx+Rvmthd
QboUII4/7Ab6qJ2C14xzA3EItcV5uukzVnR44qB/L6JTKzZCZHO06pWmu/NF
yxWMcbILr1BVSzAshdw7NB8KxCnLT5CZry5vmqRh1SLCj2yO5ozl8wNCIrT5
rQEN0XCgj/KOT1wmWIF9EIISLVU4PWmV1FRRq4V6h6U97CwK55bRKTLcaba/
Pm+0N5xy58BCs6C3MOs2OpX+ZUQJY9Mv0zpGeootFabkCUmG3THWCvpNZnOn
soN3uNXcMm0wpCzSLDeKcASj9ZNIgKjiY0klM/RILl0xHyf+G10lw6lIR650
jubJbZWcpMJn221zX3J/dU6E6DgpIG6YIa6yLiMOOyix/AzEqn8Osx4dhTyT
l+u1pJwdGoNS6D1bU1mcP0beUC6hRVgGAkgeLDnDMfIC0eTKcK6lA6d7J8ZM
A9hgIt14LnPEEyFTaRJEQIpab2RIS0JXtAqGghfweIvUDeFSprWDcg1X8Isg
BryaukFDe/Rx64v44qEZRz0mZX3uXMGCt/fkH6xIuKUPCU8h5PGGKGKTtpSO
GGzTXajIMo4mf5fq9Oa1QKlt1qlTz+4Dnz6D4IyscDTn2oG4uLDEjFBYRzTb
dwKAE3Sh7vVTvmtjVktY6iGawSLdtT37vGl6Voe5v9f/u46Kg1fVCty8SYmQ
nHxfxkekh3ceKq6SKbN6TRAtUPeAodzjUJTr2PdW7ItY6ylTwB2CxzQMSgbV
iRUGRrudBBvO3NOCFl+F1QQTQgszEqsUZOA5mRb5RKmyROQ1nYxFOjoNR7Uu
4BO+dcgBU+RCWFBKGWVIe26QwLJaxBjLMZi62TwfvAPQnAbIW17XnXbIkjZ3
fdIoHE+V9JqmEKS+X2PoQZBnT7sfG1Ay/4M5wkjtSAfYckrIja6BOMmVq0Ny
m73GMzwydgl0lQy/k0B3F+nUdCuAFGsz0z2MGH5bk+XqxlOnk2MkZAXZH+tW
TjWO4iSnnhRG6UuXm6AIkihaevBgn9J8faQiGdBjtz9ZcJ9QUpqKN4K+7xVJ
U41bfUQxxR3VjMkWh4Z+LJ/WZIZaRhP4Sg659NyvnSeQVO0ZIm5loNfJBAlb
kCOS92HLDb7MZqteQxGnuudV9P1gqgRHaQ2enIaBv0E22ee3qJpT1Newurk6
zU/OhiypDr8H0Y10AFE8Woonn1IFCsht5uv12mlSxZq1wLhRbx2ToTRekJHk
pokWF/3pd8LtGrLeP81ZmUt+UNErzd/267ADkuRYYlcLAxQVk1SEBt2uA0dJ
vYkVwtE0xOORGOlzjIQkP3YLO1JltnhEVO7ZzCfXwOFVWwLIHkLfJEvBDhno
SkQw7HebrZiza8xY2S551niKWmmbHMCwjjhOUqLSMMDf+M9eg1mm7Cy39rqD
rqKfeh+5HNIKMRASSHIA0VW4QUd5z9wONdMQyQLJBYzmhjGieFlsvuRfSsZm
ceXIrzquD+s49qDYzBNmegLq220NaVKk0kqkq1cTFKtUYUbQqnweIepP3WgO
xkz5fZ8nVkKvL2vJhpIejImn6Rl7izCGNWz+RmLh+kFhRK97wqabugtyKuIt
u507VVrqR+J4tiwm/ZySD2KMme0NzDOGvCuqyVEtV4u6fHxhHwG9KK/Kabgc
hzlR3XPK7018kNgJZ4mqPeEAn/X8WHXpW/Q0ymwjrVDjoOxAJDVCL3wf6heg
vgI3BAumSzJoREwVda4Aysa4SGZTCnh25iVvGQpShHBJXFQXQ+9f8/kyB/9o
TPf6aVHfWo2229bI1jRGuks+aSkTJFTkC+4IRDaa8+P5QYJpe7zOlJ57sRq5
wWwF2i73PpCph3OwEu0Zpd8v2Ib02onZOZfmtS2L89ftOmVHSvzy5zzEBiye
iYqVdoLUqCLdkYzLZmvtk6WqQK9ISF6idRqyHx9gS7W1oU/GVUXz0LxEr1vb
v85ZUkx47kvDJFgcfebT5mblJMRnddva+DanafjMiZpzk+dAfUdWEUePKyCu
zodcFiE2j2pFyfZTcFu0GVAU54TPWE4y/jlHvaW5fBHPIEqq5X34Itcol2jM
PbHyY80csL1z0ilQYcSWU++elB61U/ZfdhjLYVC35/dT5S8GZFYE1zZEsSaF
9xJ8VzubKkNUlhktuCTtTUV1WIroJZjenaaiR0JYWrWK32EIUW3yZ/5yaFBL
tiCRVAY9rSTTs7sAqUKLWVgquZfR+bzHFcCYBM9oZQZLIHPuV+uRFHAd72zA
z4yx/Gu9+9GE8zZDNFmJ9/BHbU+44IVj7pCBt25Iq342ILAycTnV7AKtczUJ
zbjMtUptJtln0z3k9S/cHbYwGPCN54z7nFikZoyRrezh56CeYIwbTy87q1DQ
hvtcJr3G05+BaZywCs4CiQfM5HdopBjy2dtsH7VJN4QCxldeSH+gXMoUezdO
nMXondfb/eITyXIqBrP5mGqpSNvYh7MJAw/yfxOg8E9MIfxVIjKCRiuijvBT
yo7bsWcqkfXjbn3uWjNtYYiUSBZ/8r4Q7qtebk75ymoNXmg1jQdgqIFgUsA4
11V9hUfm5f9LicXvnFEmOsagj7izO1FQJHJ+KoyC1kGBB2//1ubiR53d4BmX
4Qk9URClq5rcTk4iThpf4r7/U/I36ZzWWrzJxAMSvOS3CdJc0mc6i+YuGJ8n
6KDIrqCjMAC7sGWsYx2EDIlbih4a5WwAHcvo3Q6U2XuJ2Uq8cLMUQSUqyDvx
Ww4uRi3CmS6eTdBmrdwLHEs/E4FZzlElJA5OhMOyvHxz+8doMrlJLw1AVMT/
m8EC1V0ORJq4oxNiYnmYGhsAgIfDSJwhmkumxyy6EtNaHBP5aBfhPcKrenJC
0nZEs8Xl+2DEuTIJZhHAy1BSY1BcJ2Ah/an6uVKkW4MPmir31C/07bvSgm5o
xUazQFNXAbVdD0NxAr7otCzeM7Wi1qoJf5/qMxMMcnYziYGaiNBRyiY34RiE
ft2WUUy3+bGtGYxYhm6ggHp5gVwNroe+DFje1YWKSTbtU6j3KdDgKz2Dmd7j
r4YDCQ1rg7Dgp6oy/oE8L5tctAY6xra9DvIAwCXkiCFaIS8XT+K2Ol6WL789
LADsIybsltk8n8OzCrTxfxj1qJ7mMiutsYOb0QIV5snEU5k0M2hU8qBuEgEt
gykRwG7xuG+9YMqX7JuYu4IOkWzw4fO711TdJ8F7jWtUDYkjem9j69TW73KW
Ncs4dqC8p4NZ6wVy79D2iHZFyq+ufkIpPNLyR68WZdg5+iseq2yC4bpLw2Qh
Xi9DD53OMZ6PMGRIuK2WPBtW1cd12IAu+z//nXldlAMayt3ic6UUGzSoAnbu
8qd1lWaeS5EOVlxkDTS20R9BJpsS2xZH/Ah9QwISo4gjQ1YVfR5T6mIfDjn2
Zp7QyMs/ZFqbudVux5dn50shcbnXIKvPoenUhC+Mr2Zz0t2natuoymokvzZQ
qUVPirDn/YeRWM7K/gdXRCqhRBigyoRsCLACNhjR6kn554QkvC7p8TtY3Cgz
XAJ80n5asyjSgPjXMo4hZuzHZa6PhBFD9Nr5F7oNYRCyk5vyjhpPLso0+yTe
MItS7agJSeIV8XGdRA7VYa3SvLKaslXPne6o9/syFPXuaMO+PRBNLTJaxmWL
jEAVT+aaQd0Z1Ay73BEI0D7LvQYUXvuZ3eeYOgCSdwpvLZveia3aKVMzeA8k
yGRmMSjlGcOA4Dphq5uLei/AS00TLNlCPDzwLb7nCpvENmnLXbaPva7n5a91
O22ZlhNfhIzAwm1KvONFUQO5RtXRPDqzcRo+S8nX2b6wZvghqUlbcd/l4QGV
qNCa8Use7LCuZeRgO18gGn8Brtlt5/UNW3rWSNeeaa89cBb396dA2LDqhBJ+
VSLOClhNCzrh2BCaKJjZOHMBEw/H7EoqPa4V+ZU6wzWZm95cG/gmX1IxHf8W
lkHM4pi2fiyRhP8frrBLe+U3aEA2Nm+zLXw32gXrxDlsT2CgfhXEP/guri18
8nkdwFzQ3v93USI9v5n/lNhC/ekxkT9vddqMcfK5+Vkey35ZDg2aCo0chYIK
G8pPJuAe4de8YjaUxKBfqqmW9rp9eHnWtPszxSEJgkwuL6FA8QHsUFy1q4Qp
b+YRvoqYE247XN2IJsX7HWag2WqO2jTkbZ71Dj+/D8jZ+3tSiKLOPiOSHKiW
pYiAwcQOoREj7s1cLwzmiq/ELsPeqldEiNNyL9ds8McBdcZWS6sXwJk4RELI
udlY8brJWrPkoIXoRC+4dfVZfGmc1YY22m78bgVD34WFYqb0bNWC6Zudr0Xw
2Gto0l2sKeC6XqNwH6vICmEIebUC72Qyshd5YI4R7q6sV81CqbzDjDN5waBu
2yL0L5c0ymbFK4ZASZdMooI8mwi0PvI6H8nYlcMumAI2N5lntF7uPC5tmJtc
WV2xLOxWFbx666jEcWpY2jBCb2u2/Spu30RKL8oiqDyiMJVZlVvf6/EVx8BG
ymgKJvRvjjBSOTwg3Bd9tKg=

`pragma protect end_protected
