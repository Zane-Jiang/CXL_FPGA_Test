// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HyMLkDq6P7BKGuzfFbQztuedFPHX/SVCi2TatT3CXHJBJOXnv3SkfEUJ7544
8ACTpcgmzEbHEQKWE0i2GaykDUoHfYKjbla4zReqjj/ccIDhzDAAEfceRo48
jpIqwura8O5qJG+2ud3/vZKWslk6kCAL+YZGBl9X1r+z5ljvxkFkWAtgQxhA
Dr3rXtm5MsyIFoMaaRCzDcj8LtenLRDuBB2ILxIyPuGh1Mmf7oLwKjXTZWKj
ygH/P8E0RM2WDVpPdKCziyCPLytKN87EnCzPY2+z9TLFPo2twlSjRfU5Ba0L
fWUUXXhAxDhUwQxI//CqRy4dXaH01SMGH4ARegbwwA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V57M3N8N9yYQgRKxO0mTcTtqTkwN2RnKdjeorr5YvlYK9a/0WEI5H/hmtcJB
DV0bnPZkSVxqfsqfIBvXrNKhl/VNg/LgoA7iBlKIAHRWDPDrPvZwiTv1vgGo
khVl8P5d4nmfquFb5+hqqHt2aPfdRElZ0JVtnA/ho2yE0EIdPEH3n5AvWpWB
WKZesGUIvn/YXtz4inPbupCaFJqmP5cTlznH6qvBRGojsi55mZORVYgtAtO8
ui32GggJcnRdGGRre5mP+P0tXU2uu2e/UFJslJ50HEfrGObnbOCVgCrEscuJ
wY6AH+1zFLsfGYoT8D4ukvifoP9329YgiEVIlv3VtQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qBogkHNe3HQRbMNUf9zCVXPLw/k1YSzhmFMyPJUduYijqnddgpeL1b2yTRW8
YdwGhALKzOYcKHSNqyuyPboEpcNWIn+kPe7X3jXKa99SVOmmmP9BPrH70xWq
pKtYXW4m9lHjDO7c8m0FEsfBZ0fu68kJfvcHlQJaqogjLw9JZ/OnfCJ+Nym7
TP0YUb/EmPZqgeZBU4qG8yo3mEV1gd412Iyqa67c2Vle2ZnlKv6Cn2neKDDZ
KdJikihiz9+wtUbvJ0wnuqxoO9wHYhiB9tpuMO/RySgKqjUYiWRLJMqK3fH8
22K9HI5DNwiL6UQ18Af+h1mY0/52PVpXoc6EvRLTOA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
C51fE7gZwwbNh6jht4xkBvVUjUFHBiCFLVRTnGG9ojOf9mrkOUdy3uJBDV96
eoqgCaO0vjih6rCRkhRhzmzvfB94qdezFQsKzKYqGOxuuvkIn/izAK54KIBO
40bvDzebMEh/urZ/Opf+GouWVt+IVw+eh0jNyBty4DQ+BQ/2ohE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Dsaev0gDRdItd6/cD0FiKJP1Db5Aujw8YhI6OduKgV1+sTWXqyvxjxSZ/1W6
SY4VmtQc7Z7mZMuYsbHJehoZsNOZV3ZLexqVIeQn6OkuqS1ezU/zmy6E0k6G
w3G/n7cJr5vBgJ+p2WRKhyxOPKUEFHMKzkXwyppK3I5suiSr8zZGQHLmZmKP
MsS0ZD8jTtw6pbQa5ER/GkULa55JjKzwO+8F4IiAQAGHNTjC9e1S/RIsRLVR
z+NCXShteQYvw+wZF8QQKeFKtUEmSoEw/KNW9dHZhyKxs6O0PHo6pikBzhl2
SNHNaeEfCsqbwj2ipfgzYTNK9f1pEh4lQAtCJuLGasVWeo69NOK2XWY5EF+0
Uz6BD4e+1fhbolozxqCIinS1p98PSbkHci6cGKOkEYFt3J1CbU6KOU4fVU/6
c81Rqexn12OQbukkg+JAAGDrl9eFGV7YekAnq2ZkAA7TC6lUEBFzI/6NZnLB
WSYNwHnpYB3AAb7DKgkLYr4yLFWB2k7L


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TM5MLGbqKWquMSGaZQ1yjpsg4c2fPahkpY+Tvmr76O+lvssnUdyUCDPDFkhe
56x75O3PR87i0kBXnma7fWto2jmrqzD9oripOX1x7d46P1DycxyJ49CJMVXs
QJd3wgx6asNdYwc09dYpkyICXCocAcpcHe0RKdcicQrQlPCXAPU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FMmGYgcnDto73iV/vxMayiTE72dDeWAVdYpd7ACcNWfsTQQJu0cyfZxgSzJC
Ee6CCUkceeR5cKYRf7gNvxf1T4uvpLitbCjd+XCLiPLeS7/ZaxH0o7h/EvU/
j0g79UsTixqiPZ4RCq6+9UicSTLcBazRymqnIJVO52X0ZnJEmbU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3344)
`pragma protect data_block
/+fu8lLP4SBxb+BgNnx0KrWuTSepAZAYp70g+3/bGvvMMvcQgIypS2SGoBIp
z+kvvivZR7G/z/ZL+4tYgG2wf7nt5JoynLZZgFUfR6ZKMenh705W66DFMqE2
fhEyOnRKYGCurKf/punWi5Thw/ZI9g0x0hwo+anG6PRD4sblgvdDHPje9Lw4
X1a10rw/3Gs99Sqhs3B+Vz+FKlh6THR36IMR6USZ45VL/ipzg8t/GpOb58Xv
+CPlpXIm2QKy4sG23wjWGVGxwMe2dkrZ54s67N8s6S0WejZ/wZraN9PNpC+6
iomyE8uip1OKjB+bSfSXNDTuEa2Z/zHKtMufz/w5bfQ8gOHnP4uKQPGn/s8/
MwjFDPfdFwSNgfkza+Tl4VZA6UAcBPWIr6UmHJOZRBNjwI1aBaq7PX1/Haox
0RsQBzQ0Bwx/NPfQftTmwY7UN/PZSgoqnS6lZE5HW1EeDch2QjkScZWEzGtM
hyvsbSgmmMDwHScGxkNQhS7CVkCXIo49/HwPszYZhhMeE6PczV7kh4pFZu/B
nHFN7c+XdcShKZAjdhUYc8Se8QCu9EAlvlCqX9l6FDfJO0tDjoPzr8zue6pH
ASTRSpZ+0t87rak0oci5duicoSfMnU3H+2gsmL1wdBpxWaZjC/xsi2o1Cgpx
mGOL5lUGhecWFz3edYUCbjKV/ThaUlp5CP1dZpUHRa906WBupXYQK+DlfdqM
wqEcQ8ZgKwTDg6M8Pu/0d7LdKSkubCHPcI4K0KAUaCsLfDwQtjIIy6slOS3E
lUfkziNytUE+Y2SwtPWdqyfmE4HPqnTePeHJ1ign5t6OVzFSaJVsK0QTA+I6
yZKTw79r+ADITxgJ1jWLbAiY6iF9+zQtkOmMDVuKZtrxy+f3p61Wbhuv+CgE
1dhnG+sk0CyllLjGHhvN4vWLj/ctXhzrLorgvSFp0ioevL8lbhR+UoeOGbyG
Rj91Go1ifQtzy0N3gddxXxHX41GoGQz2R2b3THukJ6Hc3jXZmNTLaKsAxxkd
otEVLSWr9Hr84hJ8iq6EkKnNNPH1mxBnoNqdD/ZubPY/4Xph55O4QlPIV4Qm
wvBSK0jb0aFpZMKgNxy6KxJUkNZh86nHml77fE4KtwWqFfYBYlECpi9cuXI0
g+hw81lLFPWY/dzPdMlBpbGBFIiLSFPN23BIjtgMeKOOWrZvoj7ODZ3KQKJa
GQ2aclQ1uRg0rFckJVTqsPUuG18m0gbTb0yEVOV2vWGPfBD01KhE3cIMgwU/
i7T6vajoodW23P05aZZLPwKatvgZQd56ueDm3Zfv2okes64ZQRr+JNzb9/Uo
b84pIyDb7LAMiHkx5MK0CoPxclF0fz258WVy/XEPvK1Mu0fMSQEditwP49mq
QQEPms9o599ZpzcS1dKtEOGZxCo5gQPN04N2ZW64M8S4WQx5bHGmcjX8HjjU
oER0c8PiZxLvZ//8Bh7izDtZYXCXslAGAFxuoe1tJnQFLCpgt3R6OzBusVp+
2rXkIw05E1hgWt1TsJDaFTtJhpTFBGRmRxeAOglLcKqbHcnADxy0xy486t1D
li89VmAv20LowCs2heaHgv8DkIg4eE4TLKDkqCyAeXRW1sZkPtJ8rxCmgb3G
CHS/kIvux9o7JEX5X5gbRayx4Yu8rJ5jXIVRhL2B0h0ihddPuPj+Y+O8N/rl
s6+UWbvrg7wYLPQS774Hnk2WkhYk+XwB5wAtzzr9T9o15JgJ0ILtC8Xlc2h+
IT5VDWRmhdqXq71ALcySgzlGY30nGvSuobWjH7IOb4SbInPMPYsNODlJ3d4M
AhPXTXJKolBGgbbXSdR6tVtEOB7TgZ/WVA2wSFlZLcRLwAcYuvQdWf8l5Lvr
HXhrHW6BWcKJWs36sRT5p5AcTrMfl2x5As4BqZipx+kihGKxblOY24YrPRkS
C8GE4UTCk2oavwL6C2DHWWdbkKRgV05VdoCLs0t3OpaSfGbyqfJeA7cGbDEV
5+GzSH9LlYAV6xPPzV7gDZFdHOnWXuaW+aqdh4oQ8/ywB4zT2HvtuhiMAHRl
dHVYypwCPy4md4EdSr5TG8t6MY8GS7g2ErZQauQ9NKnzRWjcTORS3gxtv6DS
xlcv8IcxCYOGyzLdGu3wpSJLKfSggG11WJ1SqUnSqfdyn+ZqvejIFpNr/7Vz
E/UzDAqF5WIY5mHf2JXDHDjMBo0ewQs32Lr0XHxFyzyXB7cq6rvF1FcGGPgt
m03fDqiNHm4nBXYA0SRrUS0kgG1cfI8oekNjKeMXk5/d8V24fV24mNXnPzT7
vzJ79R2ffg88i/D2IHJaiwxkryUcOIip+PK6B5cIFnGu0LcBnjZHVv1XQ1sl
j+Qvb/DUM3MG3hCQltqvqFlQ6JcML9FswIDPKxJkSZORaRLq4b4kHlXzBfpe
jylJdG8+euGm/bFwDlNQiV6FWOKJD4OObTSyuV1nNVjcN405O/vlwftxXhqF
frNIvpxIIgPeBHidleawXVND07t7bncRtQYINtDN2PKy2k/ScMAYu/INmXr2
gwBs97p75s3gF5VZLKVVgPJ1KBb9SaSVYGDvpihBOSVSUwZ7rMyNEcZFTYLB
xILkJjAUlGjjN69bNR1NrW6NHcC5KzQyPX38TsEDVN5u4GfEf6hOy4LGYNKK
mmek4Y38IDUwVxLbg8IdxH3sit9/2Hdk7ha1vMPveMbJhxx/jrqPz4F7vslG
ohqP/L4Oj6088/YvM5JBZGEgQe7yro48S+Z4PlTQTVRCsqFzygXwR+q1zBYI
6wuenECiIxZHsl6DH7icm5OG9StEL0Uoj6H3uQUFRi+Lk0icw01bBhDHzpDx
+j1nUF2q7NJ6aDO2wAXQ4FKieuALF7hKtugdB23b7t4rLm4HjvLlUt2Y2MWf
dBU+NoudIorYPbRCHzoxea1y2EP5gskR8pC9L1dGJlM8ZnX7Q+hMqALlJ2fE
tktBGy/VlpgsaWummFLuhjameuTLRjpbkLlYUnbhOjDwGHfOzQY/AZTb7lUi
JKa6Fr7a6be/+oYgoNoVAxFT48slyyLp8hoHAPBykEXhCgnh+cPL88WSBEBl
3bF2eqvCJHu1ozukjQJFdJ6s0O8wNeBPzDA6/jUp5/5ZsRIfYaDsCDPQUYqM
bAyOSw4qsZUwMr5WVYc9xR7uvkDpzcJTFzS0e6MJHy/uOTJeAbq/WUFN7TWv
z1mXlWb48xbPff7CufTpDcRCdv1QZwdX6NJ5Ej989vwXfUzua5w3egWpfA44
9xOmugd2NzgD8TxQMcqMEnbbM9vv49ZeQfJfGF3j1UCY7+h94UoJ4q4OsFRK
iIIzQZFTk1fziD/OKG9iuL+hufdvKgrUWZ6EDii+MCd+psCHPwKDL801nULL
TgC0LcTsEWBz8U02FbyyI0GP4rStfXMOO3BE/AhYWzEDU2/XyLkAz+aDO8xA
D+dyeTFsgDZ3G03YmCF5t9wiZrDa94pMrxU/JuMNzliqVJekiGn/UZr0eu37
EPpgsRNWkzsi4BhPyZ1A01Uha018IFKEMZl+agILEbnt0e5aVPlVKM/k379+
VmCIdB/ronms5q/vutMzpEUQzJPIrwjS259m75iPZVcG6chXgfqqTE6283JO
ra2uQvh1d9qnz1AYriJ7Zf8JH5oDX0yMQTid/du3421UQqNWl0/UT9ErUZm8
5s7rWjsYScsWKlpSD3KLKJtajeTMef2qOL0l8fVUNMdCaSjEh4XBeh1vJsAS
cp0NCf0CqZIKskqbLyIpOc7BpfX3iHV8aw5Qj0fHfjspAWMVsGx33xz0URD1
5yjE//dXrVNAeoUvJV/Io5J91Y8Eqg9Ji5X2rPlz7Cju2AC/u8qOjFfojdpZ
VteQXuogrzLKW718dIb2NjcXk6RkK5vpLdmHBu0TGed10Za049Bu9g2LJmwR
SDySOmIIRR63cKuvD9ywIB/2XTOOWpeAu+FMefYXahjOJ2ce1uIgRfPggf1V
7E/5PvJO/HOfwoYavQzoK/ZHxAz8i0kmPwvk7zAg1zbxH/3rQJw32bBx+xta
ewY8tmgSfPqges/6KqWYeEyB2OfD2wMY96K1gXnBMyQF4I5inbfQYGGRTLaN
b/l/NuKzsOGlJFzvPgxurirgyLW2+EAS+IHWQlgk10QV1SibYfAOvdDNvLSH
hJO3P6Ch9jgf4LlJCrb+T06FuxqV3Z/U87+BKHhZjtidS0DKZ0GhjTTN018B
hPnizGFx/A5MIwltXw4+ZVFmj2pYCtuNt+a0VFSvLuZc7mKy5OQ4avHlpbd/
9Fg4fSQy8JsSTnyL0ORKyZyssXa4naf82g5Dsk0r/TrYXSATajaxzfKeSaUA
UUzTIzTgzFzQ4Cn62T5/ZAv9bIObuRNRKnQbAYs28nopmftaPH2bDvTlEbp5
gNn8CpfCQb7Zx5YEpbkqmb2tIWWdBok/SiwDGvjKoZb2kQl0ClrClTZdstji
KWHxf/ZQ7olJD3ofsDk=

`pragma protect end_protected
