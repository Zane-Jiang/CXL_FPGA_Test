// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VO3IQN0nK/kCmZ40NPWpdZylsCUa5BPbyqby40QtOfYAH1uZxNKlLsnoPqzs
Z/03TIL6fP4JUwlj7ToBofXd/3gd327poB5ogx7G7q1PkfDbUOxa2YQGVbHy
fwo9bh/km5EdMsNHaHE9YUBD1efLiSYXvSVnvfcUFzJax0JnIPkPnNd5UYVD
hp4RmgEt1VMmrNHCeZp+pUWJNQ0d4yStPjE42fAUGgeoDgsQ1ZqQfLThVZ4d
c1XHIadhwrNsrOzaXNmj1A9bXCzZQwqRe1P5LYIAPXernVHhYQir9XrA8eOS
mB/ITbo1JIqxTB+2xzB9XrrX8bobeUEDk+uGv+5uxQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ykh2H3ULVZqv/vyIUrS+IeXXWtcNTuKFysjuHZ4acswDaQGrmFu3NgBoP3kg
wwvvMygGh1Tlm3K1EyQ9cV3Vt2OcgTbEXrqJrGquAeCztpoJK+kF/aDrl2NK
EymeBmVqlCf9Iw6XnjHVYmdZaIWNio+Ya3w3Z09NKL5CM2EIyDLVKng9g+5I
rnxdCrJuc+ItfwVg47TxwacRDOL9fWR4txkj2gy8VxvqYtB5cgf6MT2MO75G
S1QG2/6fDpLcNoHKtWiQtT6qUfnKP2YisHQWoFWCZcSAATlZOXfrVtgPhBe2
4eP1e/n1JMYftsSbluL8oHxtL5WCGnLiI5GuRWVatg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bPRxgXjUpyFth+37tgDZKPmcW5ViuwdGgzqjfqXm3lWRszaKw70r9tNSsTdB
MqBz6ExFYnukSsSQ6Anh5Ty9E8FYNGf+yhNYqgvnkCGWU9zc0NRPCDaiDex2
RqaQKsu69DFRKJ/jqCwXqat8QpibHhSYHRh/NvsuKKVhPM91ockbGQbhvPi1
302VRQ+d31VolNXbFtSB1K6mbEUTx0SaJpzT/kKNj+3Xd+pYwzZir6B5OzXG
VeexQxr5eVOPu7gPQYxQCuTl0TvxxNWceuERhQSSak5Nbjkl3Zn1mvXAYPeD
7tb7tcsMe9X47757FsykvykCXPlBXvG1LQNKBe5Udg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ltb52kk9t3Ve/LTvhEFoi0L7Q4Z/zwkizsESWhKQt7fhW4hgsxPdBLDnXW9i
fCF5rmTYWYatlMZvG2vIitd04Tkh8HmXcwV86ACVJMN5hURAVwBh2Y+yEkOF
MH5d7KttfX3nLCQ9It6YsKp4A9MKgyy6O0Ebk6IKp96dPQ3/+xA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
iyPfni7V66UAboPdp7hIYQymVxom0aVEL+mKSIa+TXGhq2mwiAUpYSqN+gpp
R9Dra5vazckYtj6DAiJWBiOnaPxaOiJxdgI265S2WNxoJSmRof/0J3iWSDC0
RvDAIsydpyHlcLRSUb+GeMlnJF+VlIu9/0QBlLPijR8Xo3ivvBBMvIyXE8Fh
Ob91X8Hh+SwOKsEBb9CM06bk6A78ZRIzwtb71xMt5e594El00oW1xAYEaxop
oHG3si8Yj57cnI11Svz6RlWJvttS7Wb0TEBWzDD58S5C7IQEVlw2KrF3dOIn
25DVSbJZVaOos+h8dnoC7dfaeTRG7v+bEyVB3fnfnQnf/JL+ryeioTfs/EBW
D4TVpy48iMojCkHbh9pifXKt0BCtK2wNMhUr5FaT+CM+JnHY2Is0qWZsmnSl
IVbWV+zv1j/bbPj9KdrG+ZinNoedoYKAFOBKnDvUzNdS8xpekjw/9xJzKAd7
DpiiswWfngltjC0LdtH22kkPkWzLRaPn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fd/QhbZhF8JiKgpZ35Cbz9pZrhQZ0/RixnhXji9ArwUBrfP9K7c0qRSFsQzL
7e5jg4acwTC5Sjs1QBseLf7gZ9OTXFs5FEd9O5ycD24OF9f6VcHwEKHshlLM
F1P6vxsJQM74QMtPCLnjc6+oA7X61O0SHkPTx7gsC/Ih2un4A8g=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZeYc15dMhVEeoDo1e/eIa4P/+HE7sKlNowgkiEXrQTyIfL5GDA9qgbL69QCE
n2MN3OL12yuB2nKES4FWI3bm8bXERPzdQT0JF+ZDRm61u37xpBl0zF/35eXr
AqtCesNGmGJXVWWKkb28qDGO/41LZhUT5Mjw6nshC3rC3uQy4Gs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 84400)
`pragma protect data_block
hU3pWGxvjsyTKbqyREZHa38g7ScqG0lNXEJcjZBZTVr8GP5QyvE1P5ROKGbK
Zl9nCJcQKSKOhrBn/9MQwHdqoLi4DjqS33JPvAwDu3/dRr6VsJgU7b3ciypW
vU8S4PDg56hPD3YXcBmKKlugci62NE+TjIh5L7WJs7GUQWDKlCItu5nfHB4K
m8+vUbHkF1aJ9NG4PBJfFYy/+q7HSpgfOTa4nbcmzzepuGb8jZDkhkLmi+g+
rXrPqvUijThLvHGTCOpPdMKPbpFDakeFe4PQ+S47AzgXqo4RdMYP1yaoWoKT
uavd1OCLaGRUuG+oO9Gn34tb67rkKaHRC1k6Ah40cu6syouXdEfOPPzn0B8V
66wHbbVl+pGl2hgHpTQLIRqwpusgLt9PEsHijuKhs7nC5A8gQhL7YWnUDsk6
CaA/GT9x5ldymVanKfu4yHjHksPvvep5GUunqpjgSJDxA8OPtBx//K0M/nww
tWdeDfH7r66T/SLi2vX0tTj/GW5NGfotutpp0VGu1donS5MWRhGVG5Nd+B++
3CRlQuz/IdY8r2+MfhNYWuHwBEIBNiVMkoRnbVXiWzlXomzmTk33jDi2+Kqv
soO+sFn39nUQliReVsryDsO5QEtErVF1tLFdmQa3nyHD5BYkWVSsxmf9t+BZ
3Ld78Q491gWU3emWRTIm/3cl/f74d7qq27ZNISN2W/unhEIDWJCs3Rykgcur
kYEGfN+w1qR0FAUP/zi79vvjfq79CuVY59GAwPFDwrsTIkF6LGpXSr3NCNeJ
/XczNomrC5+2/7F9RsQOOmXbbFGPn9oLaBL6STcBzzngpTGeLKK1r4ZOm7Ax
p5HhVY/+4ZVHDCOq1bibzKdGb/uYZavb+rsETq5GD6WeFC3SUKyauXSGIZ+B
yFA/Q5ALHU30K7CDeYhWzTo6PgdorJirNW0qo1nNmKzhXk4nUI4IOrZMWVOH
FOgOL71zOLs9vMGOQ4/ehELAgg+KeG8dzsjlnInb77O5dwsZ0I62pjjuMLzM
KpxtbuoivlCmkwfYKE3RVxg1yzDQMj4GNws15fn8QjfrGdQk2AuDChaO+t8J
n0Gar+T1dJ3KH0sSJ5ypyEXAAIyaPDmeDwP0JZcoSmoL++DS/3yIFQmMTnI/
BX/qR1yYcCQYQZ0mO61j48vGOMqZ6dUylRY5TJG5q1KSBJDyPH9U/B2lkA+n
g34Ptav0Daqe3oXAalTZUw0ms/eJbFZeQgjx21ufonRn9hYbbL8Fo+CK/FlX
c01H+XuJ7hXF5tDo97NAoV+EQeLtOiNFTbmKvoSLHBcaSOuGzZ0sVRKbO6N2
915xcJG15OKZTL8DRJKAr4YqChcc29LrdFxZ5j7FqTaGDHfbriuQn8bvFcuH
BO4BSqiuRjP0hJVmAhXMa6RkYFQNmcuGCR2SBvNZPOSgiXcEILhx3Bf2/Qdh
NcT41MMX2lV8ypc8O9DRp+1MHrStOHvfBo7cEhAIPcp3GJwxPy12dItqWmSM
uvN+JaVjP1t2OTnvfNvfnwT2lkkGnpGlFZKEcSxAXIb8g3XbqFxb/6SVJxmD
wdINfe4L28n34TJ2d7xuNa+gJbpvgsUwLOMFXd7k91yW+So9SfSbrmLim9Nv
QtoZ6UKd+6P8l7OTYMmH4aMbvonPXhS3DGlF6q1+m0OBIA+9oMuliqCGw/dZ
7gWweyDN13VFl2bGyNwzso85aEmlMGXVg0KtE1IHNzuL/LanWqBIk2SMvGhj
nYEWvtqDDBqhe/q0UItz/6XO+FOzNnBTb/xkkigeI7REb2Ams/Q44j3+Hmal
FC73nAZva5jKHZEv3ZZ7UYRoyIQFXBry5/yRs/V+CqEmKifQmllZH1fDQ8gj
cb+dcncaMHZkumKQBfcbwCzJImP5V7E/R1ykTe7O4U+nV+zH0r9VWuJ/yXSn
MqwiZBqbr1jyT6kU/X4knfSsL3YfEFOJDI0RM4uAE9/K2AJetDULLByJa1hf
apzoAKrC1kfvMu+dg8MS285Qyhjga95L3fNx+26G0nw5567hhgk0OgXp3a50
iJkrv2/ynu2crQP/mJ4O7IY1zHrjLg3xTaIK2mZ81VfjEWkSHq+Mq65nsqj8
zCImglCxsmZdWPTmcmvhdT4pQNaQMJXmOf+cfCBiHDSvuwqlFSuaxywPaou8
25CPIvrPcWIbk7vNqashuFfRILqfrZ/T5B67GG9tnf8CXz4NirDjEbNAqOTh
5wxaaL++IPRdSUh0k/Uf1OVuaXXZFXfadpszq3QM57sQUhxIl8TQ1JUMsJzV
Ntr8VFaM9xMMagc60a8Tyrx+mzRx6f83nlY/oEqCzfI9npt9+CQxbPOlYHA4
SpSDWv4/ammeIgXsQ0uwmMS0+bg6AEei9t5A383cP+2YMxq/nLapytIvM+/R
f9HA6UqonI9vV4VoET2UStLA+fMVKEsodbHAwGEuj1ZSNbVLWIhKXcCvpiOE
nd7J19k5YWJStdYE8GD/RE6dUhqV6dgvKdPP1Xk/bEpAIT3qqfb9pTcEXVGM
zdJpmisk0lSfP0ZqxK46gwmB0/WeTPPCseNDS+ynwSlO00oEfanhj8p3L2Rv
BBdxhY90vizKFtLeMFwH8fs60dIhWs3kDk2qDHMizYCx2vzhM+xhFkZIMhxO
9n+FuOzVj8qID9Pr+MJ3CDunynbrfgZJWaWVvxzmt78tlJLhy+UD7oCpzhOZ
38kqQiH3K+tiUxSnnevdipWUgSOsWtCuzy6QDYy/OoW2q5yskjok+dGqx+vd
R1iIHbCNEIS1wIu6EAVfWK0XMfY1wRTTSuAudGJpdMPZpxkpMRE+hU28wHEU
0sJsjtS96/RYnAEsVrgj+55QPifg63q78eliAaQQzSfFEaHI/u6cbRtJPZHI
vXgT5JDbvIGZL7+WYE3LQUhZhoFngH1xc7te9Oefwgv6zV6R2DRd8ScIwXrm
srXABjvgoAvEtt4vmmUFeoJ3QlAd+Abobor7LBBYTxAJfDZRwInTRuMdJKtO
uJNa/WUB+0UfwqaBHiFzE/yirkNw3nBRsrTdcXe5qYQPv2/iHhdqvUvlYre1
VsYlExJYqJca3UQ39cVgYQVDBcaGHE+9kPfqRFp0JNy4YLqEuosJJWJe6150
TAPKCcREGrUm2fN3z7wZJsSW2REMWfYFF43rV+RmosUWFFArZlbgfCisFboq
DaH3vEMu+VlG6xpC2ljVKOj41WGjUovJs+FYzipMDdXCKYOeKKBg6WDl0cEZ
49Bd1tUjN/r+xP8XZJB0lXw6pXhj99U5MCviZI1XL3HxnaXm5oq7VeWw6nwX
y9GH5cAjxcgRbtBJ756nTw5HNngztZdesfX2CeggJzpytB+WSJhZT8po97cF
hX8vhee4fy74my8wVyw1OGCJizLsl3ppaazd9HAYQR3/4MTPPhj62wpF82fa
DuC7zKRQXpxV3jV5tyMzgG0GDsI5gkYvrEUO9VhvjHEP/12HVl2Y6ofbm8Le
g3g8C3x1aZ1q4lQeJ9mBkj0Z5lWD1w5Zlpaq5u8MZokvjerUFZ8p1roJQ5RQ
uYDX02s9apaPAYJa44r4thL8wtz9VkGeyqtHKRt9SPyB7tEiYtJEJanfz5mm
8w+mQgAQcc2HGqUxe5pfecP2XbyJCJHwVlZNxDLx18E9B/0D0inpyi7evqOC
mJWDXNj0LRmHmxpseQOiMQImi1aqkNwj1WWraIPxUdxSOpjfN48sL+YadkI3
id7YChsbn+Sk4IKtgva/L6m8wemGSbgXxmEGN8L+Hzd5JiXECMjZIrzQlzXX
wy1XWCQd6DqZn9TtRRjKDFobyWweoCa04c8TuPx2KiNiAcgTXapajpjw0YPi
e4uEl50A6DsudHAxiwSEQ813cCSDJ66ZOqELAaaL+euDkPvBLeRCEuLWPhnR
/pXk9Zo7qo31BFgzZSONPPH8J9pnIQ+3sLJTCDHn4sqNtW//lF7ZUslzD7I3
ti8yRbDOeo8SpKwxdcKrxy9lfu1SWMctxLnTxISrNvwZ62v+qtYsnQFh9X5W
90Wtlt+vjVogrB4DjHVlIvAYZJ7pZy7gQiij0Fe8C08sFzxClG/gfEDr88B4
iKHfIIdpEl1j1vLpdSJiErYUQyYyUq5Ie9x1rXlii+7aJJEI8CBqpDwPN0Dm
/eXHP9cdPZrN4bdB60mA3mXEslF7seBcX9jj3fZJus9a25SAcZPCkqwAcrCq
c/R8seO4tCs0I/e1SSH+MXuRllsorAhibc3Ko6mfT4g907P4oLiWISxSbuQy
ruDKpJ3RpYJJDAge+oQGzuLxzt2y6XUk6MyGOITbRdLEtj0ZO3OHcyOZSsKt
2ESaDZZomfFqoLvLr8u3cBULnllGiJSZd/0ze+vxZzCbS2pqh09xhFDwpFc+
KGB88R9iU1IAysMHrnKjEwMUPBfx4s4LqiXTIarExWHl3bNNQ/GNDKazBJ37
blytYtntyvBylcq1CQLdqb1tI3F5wBOwJuJ+0HGvul9/ETdUhyiKfB3uZzSH
+VklI6virsIbMlETTFnQEoZ8f9HTfGBI1dLt0eQ1N1iDy2I0QCUqTMyEKiGb
TpDkFajtDObmwPTUhmTxuj9uUUoKQo4njmakQG+pJIT5CtppSpoe+vPYTLyf
B3TvyWgcU3hH/JE6z3YzoghwOlOWxoWG59ClWaSgN7l2qnGbtGpth9t6j24C
JNhwsOUqmmPsc+JO5BIHOyZ06nnlKtd8cTItJ0enly6Oxb4u+Rhvq1JvikQD
kUEmgqEkZOeNTBAFvdWKTCvJXCy4tE3Yrb0mtm66yeQSWKcQABsqgnpC4Dmr
DYQDtcxfNpTZTpmb5I4Qyvs/0iUfvCLri7LUZMwoUbURg1FIvh90rYCIpoEr
d02GtGpbUh/m6mRzJEZNqN9JcFtSmi9DnXV9nFKqP54QGs1kX8JRXta2XERO
uEzFCf5zEpiVliaLJLgKUbOwd25yYS2ukOc/TBfTmHV/9n7OQUr65ulvonzW
gvNZg7EXcxblygWVS+qvqazykzEa8Uu/uVX/JG0oqhUags+pSDWjJZVAaEFD
HABU7mn+csYlAhtuRLr4UXFOPWiUIuRpircTid5B6E9kYiKw+IOegH0SYp+P
/mJbsVcjDUhXULnazRe4G0oYWgTCjzWR0+GWKVOywc8tRYTSiTA2RAa6bZy+
AmOVHlhlCCseqkCGP7hH/Qq3zEwbagbI4C45iE1Bcj6Ugui/AbcJIZx4EzPK
rSYvN6oTaBOYvbhfnP70I1Wd1eks3UNTQNxaEb70e7y1Cd1sgjQ3mCWludq7
m5up1+DkpQRT0J7UooLMjXoafkHn8WWJNRTRuKhn/l0vA7HA4slXnDGUn/Hz
didr3u170WCIzTVMUG2eLonwq2ov7xWHP3VgZTPfRj3mY2/PHoiNGgJbI4UD
UVi1+0FWj7jr9si9P2OlICQI8lYxfUNZAp/IeuU2g4XYJPTW395uj6zaXsyh
Hm5BGmEnMSd+/9EF0m6f+1E4AVkgHmMj7AaX0fOlN/Ig+Zws8xC1K7mTuO4P
DP/XwLg9IXiNMElRzkjaXDxAhSZFI6t7EHtR6u4EbK6CQxCfy4q/Jpbfds5t
5Emxud7uNiI6QLX1TnXFpQ9K0YH2ReVXpHx5FCPi58Nh7n9hDV0wxllUPgwZ
nCR9gRiQsHbQVZziZ1ud7jtFyHm50HO/mmnKIX22XztkskPn9i4Lvi/yKGxm
z8woefvLqg1WU/VyAgPsrdREnlHorGusgD07XTglJzIYxnIHrZIWNg1zdcg5
VWZNBheO9aMCOKTTjWJUA7i/j6egXCMl4y5KH9TpH2m4GLJvyrr8TmTPoHwF
UeTCnpi9RQsDYxhbrJKXmD0SowCL7eVN55hgtG9dh8NAm3Kg/FRZ/LeTMD0V
QkGLFp2POvbLLYmUantR04jgr5FCS7X3oyCNNXWEOnTXbvc8/K3crvW9d6AZ
bTu+708PYtxtbCcvQ2uoyiPKYLs2+GaqaZ7MH3j4jS8cwKdkt+wDg6kFXv6s
C3KNfWsiHmmZ//rdtA8JO8uTdKsIfvb0a7n6zQhFKN3hEPJlpVsRFghFtopY
XBurIV9SVPu9MOhKFoJqr3aJ5XbRxG2Zp3VF0RJOmzwgL4daCfXXCB1NW7iN
BGXMqZ/rF3uFFSLn9+Lh1iwGAkiYoXYVB5Ptiv2B4nykkH/Ml1lFKbtm0OyZ
ReuVkgukoSrYs5gbxSSUhfjis0K+cgYYYmuOiUH3NilTZbw7umlQSxclE/5/
nywcDXohHQN0ngMgP8ml8pvK7mbWiwchyT6UA6WFcxVxNiWXgy1JMJspoJvB
28lCKFYRXu4FwlcDSdX9slml+qeMcfTIGAVB+KeqJtYpz/08zxw67LwmNX9G
zlVGdC5rZ9/rWoz1xKmrGJNrdcsMjzr9226GlyG1hLGj3jvtTkN2omeq6sMP
f8yAsZDkGxHW1m0aatubXAN9ceyq6cH9J6Bpo5GLMSZ8ZPikO8bE5Dtf8ZE1
VcHpdf50RjWLu8LbbBn47ACCYN4tiHPJ1rVQrZoPt8Rd7Q7L9B0UDtPRlzT0
3jPfU1ZyNN+kI5p/kqkACUPuPH2AxkfY8thF6QklIQxIIIC0rwk/uOHH7h6O
p60/qjuCJC91GDy5a/ggaPfGKP8Kg+1te9u2mP6GSalmvPkAP1a6NozWNBzk
CrHSYvx0372e0F6u6BOtH1KihcgrBveE2OqZTnbQwdR/OhpNkIheHvomqAnH
JupTrKeSCEA3jI17dHscNNRRRzyDYvZjPdkYRQJHQ09VTJo3+zfCSHPY2tOe
LFvG2oH71cnElPQhLeTFVjoKOaNJnUKv1QNyI8fuP4cRvHCs1dWZtbaRdc8V
8ds+6/jst24zFmxriHN8+k/O+mMT87ZhmxWb+FGfsGiLBQSfvZpvc+xGcx4q
tkllMVwWVj3pzaiW+R+EnxzcTZPJae36Ll5o+ogcOSaB8N8woymadGR5CEF4
8Ui8k4QMUauqWg2wC8CoggtKpRUfLj+3QlT8rF74onysUYpukxGHpJCDZkfS
gNF4A5f63/MxzNMOb/mCN4WQSk1+FaQtShxESQpcW0k4wpWtTfiVSkotXua3
B2beOMf9BXR0BNrclwW0JbEPp6wNO/agrruFLteK8vYS4Yt82iJ95tH2BPta
nhVmrvw2QTruUXFj/9CcnSagtQFecXvDHFcS1Vp1xVbvft6K/WjXkGf86eJd
MK1jKo7clknkIYqEOh3ivkmZF9pkQf/0KEFT7eTwxopfnTYwj60GwLf1TUqp
U4tIFRFuk8kRvJ5Vd+V/xdUZTlJGdN5/l3JxnHfeGwW6phQ61iv/7hgS/R7H
3EErrttzRHd9tZgfDt1CY3zCjrr1rJvExBt5JrzsE7EYCD6aXrlYxKkGjHrJ
PmSM0N5amM1yiLXQr0mxMfY81Lup7zzcez6kKUQmVUIXVp+5L8lAdRCn/rNi
9BdEdIfSJlp1NK1B9KldiIHwWODfWN4CwnGpbKzo47bz8+cn7NlDNYx2CgiH
aNqnqkmseovKo20tetrhcKfuBDkighNjKRMOs0MAtlQduqqhKUBOKJk67hJL
TT3NwQRkCeFzhSlrUmgy4eyHOUB+XTObQDwHXauGwo3my/xhpNMw8lv1dIRM
VUWCddhYzdNf0NtiiMFHk7U4hdDUqcmLr54E+0DWErJOQc0sa6e4OM1ef8pj
TYhP5PkRjmPqqVWcnwSYECdTjCCc2vowji8fyK8P///PyZhdquPYNtWqEbCs
dkWdqffb25r9Qnuv0VZQ/ud+c4KIfMJSU6l8FtT//iNJDtLdav6771XpvxQ0
bNArzUma9nwv+2YRsoJdS+tExhcshLr2lH9B/nx3UzzwSMrK6Fz+jk+uCGIi
dVNt7PRZJodkIaWzjEGo/P1kPI4BVu89PMrB6Fo6TJPyN6kQQpH7i7V0qjgg
TM3W2KMz+4yQQCUcHQ/OpM15+vrJMCy/6OmDBypJrBOyBPYBQlZLtxBTfks3
luPItsOHGISfj+tZYxlrwooP0TZekmap1j5kUlNzubWS6LJyyhL62b2O3642
ORIDqkZIdrR77DOVrTIeJm8VHhibZrJcSmFTIZi46dH9Rtt9R2hT3dLdgh1B
9/p4AcQ3rpNKg471rcco5rtRivm/CFvld57n4OaAtUFm1Pwe6qa5svgVsjiv
8yxjutYx75JUnCmk2U67eOB36Wt59fB4mteBoGLn6yHY/YtGS1GjJQFTv3Oq
MWzk1wqZBwAwzl7UgEpgl7yABZb2uF1yuJaAK1hd4pWPKmsUwdaDRodUhyjX
dv2Hgfn+VO5cD3i6BMCGTNkQhrSSHNnCvuznKZ9mHq/qpmKEsbNSxj7MFFhf
svLrcQ3JRcy99Me3odFLni5dHyyYv863JOhQWsCkhNG8Djxm7GVvvF8LsukI
3s1OrOzKVERwgAHeyl7Yffb3VgNDFlrGxOmBXywXySs0gXrZ3llMggfrKz/X
mOPKyMr2lft871VNiDdhsh//Oj4Gmgv9yX7uipoR17wOQ4iQwN4JPWrK8jOU
SuILBahP/LBS78kZuI0Y6ahvMaRzjBv1qSS6qbnogl/yrRRXRInNySxbROL0
q40gBrfh+2GeCx57/UA6Q5YJHo1iI38JCPyGqLHCiiCrKOMjGqxLX8prYGAD
mTOLhEIM5uSfAUWlfd/ALQIRw9NObP/ydHH3a4mIR6Yfw+2/AKGKN8fyZZ+9
qhWdzqquQV3bUPtnV+R7U394Z56RLtsDf8ZsZnskqijWLV0G1aOWvIGnM66e
s2OYAraEdK2fKXV6/oAipjYn8DFJvj9BQZCn/JOzRPeQxkI/xKFodbwibh/8
R0QEFtd1THxRnjALGX7P1KDrCN+LztSlT99Niay5V3b/EiB9D9VL4QZ4uhSq
RUS53vtcc0uRLF0PhHxYFz+WjSeLd+bAhPmzXtdZTfkWey3mRIriX20VsWNu
5ND24+j8+SCP4lIvO4eNrK8Pyezv1zEedbbFG8H8MIyBquimBSoLQ45wUgJY
lRz/pxw9aC9sLDW7FJt3NIFEGf/Hm5BF4jrsckeREpJw1lOG5mBAPphKnQIe
HYaPrkp7gjBB5fE3Tozwgzx5p5DpXxo6SR7yYM49zChbK81XApK1kR5ly2P5
H6sRzcz1tNdHB5m21y6+BfZxo7DbDrDrTiHaoL7yoUs6d8ax7W2mqqPQsFwD
N9SX9H5UCCZJ0pREWD5dyFQp3BOs5sryUT5uB38AmL2cLyw55zDGAYXHVgnR
2kQKjGw0LuCB/5Barkgr1Bl0fD9TNnKsCQyh5qX7+o4myFH6hk1HwwTC380I
W4NwI+FyCenIx2ozcKmLAWIxzXeVpxGeqf34lhZhu7meujZV0iY0Wd9rapUL
ccPNgbdXJDq4U+Ye47pa3yr84Nj/MGK+HCs6vVOwEt3V7Z9r4AdMLiODuWDL
y113uf3wABqIedkxhKeH66vu5rHLqpf9AGQTjlKsV+zuIzQPlBaH3KNnN8j/
+Tx5UE1C0JOMzD5X5PYgY+AInmLANSzR8mY5+Gcsg9V9ULypclUiLnKrStm6
NZ7kxodzqtd/DGpndlISyO+U9KX7Co6VUReO2ZJ+piw3GsljmHM8Crzdk55N
fr0LuSdUPwsU/kl3RlgW9QYLLmSr2qhLDUt1qVELxfKPeOOX6or52XeDCOv0
rXStqAwWIPfvdtZRQFV3EPG3ITsyi2b6r9TegzlfUJxCfDhGAS8Sg+8VKqrI
BBmFHfPJrZw/nLbgXgoggynU4poOnrPunIynU0HzBISqz9mRc0lE4xPe753T
WiaQsFLHTPFvJwI7LYW9YDnEmRyUA77mS7yf0s9m4JerXhTT4NCjfDsCacRj
Y3fEKU4fkYvGts4mUN/hjT/OeoAjqmmfW2vW/y0PvVdeovufpqRFBeqihBtR
nweBMgeg/y6eI9EDxCmAr09n/EbAvMdYVsJ1ms4PX6N+h+C8wDtOzY3SZQ5d
2vPRMEgEHwS2R2neNmLG7gqMv070ibputsCVgeOLWsvo8/P2qdsuRqTMrQYq
/WS6zN6F/XwtCYoXZ6uJOb4+uTccBkZi1v8xgldmLw3GayjWNCq6ODkIuAT0
qk8eyvvsMQN9SXJ6aUL7oPzab1HfstZHPEaMNiF6RaC2xfuYGCz0J3ksZzn2
F2XkO2AmVCf8QEFy44bzHrPDlFBy2p4zROxH//AUCeMDdComlxir7s6HdaQf
kd0vHH6H3mZe/DL+gkfYL1nRVnQp1pBAssmvHndDbmQXLQ2Rybg5GezxeHeq
xIgrzBWaUqLMufjkAEaSOkHjuVkcSQCeiezGH+daapO4b7CGd+46Rgs9PkqJ
f8xH6m3RzouYzLlnK2VwCcgrF07ZnXgol9/OChOdYFzuz32c+n/wAo6Rpoui
OAGZLwJWvOEhOmmCrofLaXKJjjNd9nUjWV8VueASRrOwJXufZ/tgFK7V3tFX
wywNd6mPONlYuH+cOBXB52JNCSmyVKf9O76vwgovGOux1DFDYGvpkVRJbJYu
CgBNDSNpgFri7edgtS0I69JKRrtP/3wojyyajeHB0U2sxrVQQ+Oag6Y1e98j
0S/CNIxazLfO9hByxkE28MdIp+FPXEmay5GxjWj8OWwL1aabvqRirimcA/bN
p86Kg4v8bNrvUSWphnDg/u4r8fzxZiCpHzlnQ5cEzxeDgusZxDlj4zEDnfFW
doWqAPCNCmN2euqbIoUR6xmaKr/v0+Qyhvd+cJb0Ewi4+ON/Vjv4QY7Lw4j3
eGiHHD3bfQGpGh/d5QSB4pS3a6445UMF06jFrhKFT6CWi/Xq13gTweXZ5mVE
m0IwmCXCo2Xkl3y0NLbc/al89YPnNujsWopdCWFXsnJBcTrQxIAmWeh3ajZq
CkebQakw+WHoPvFTiue43rJY6LWFRz7txAT3zf6NuUhHRSz3uX+7oohwMLyr
RQSuM679obTs6j56H8Re8ISJbKKwhrQMHJm2xOskfR86/7eeyj2kc3BsLHg9
y6CY83JA6feONPH+gB0MMpphb9wy9CKq1i938VQA+2l3jIloGn7eLB8noDRN
Al/k5gYg3bLRBgAmvFKroyRfYVKmJNAW2Hgx2eeChwjdQvkCzG7AQurW5InZ
RfD2qeEM9hqlJG55avlp52PYGwrjMp2mIO0KrG/eTOYkw5N+3wpQ7XwLufHh
5ZLEhZ9Rh5BJIXmoIkJ7Hn1/xJnXYfSnRnPwfQE39IdI5PBHQ0iBlJ85vP5l
MgEKo4T6QXNdDHti17ltUfs69uwT9b4AmRvqU30AcGnZCiDZqjQ+lslf2PVY
qvsXfuBW9S3Vva0zhjea29qThB14Jj70zm+yUMOo9Lx2yuKz4nAtC/b/gSYo
PnXpOLhKXRV7YKxNk707UXBdRRZ5HqFTOYL5mlf5V+L6HwonV0x8lnixyBcH
hhTYVX0nhbHRi8ptbamEaS+OSfRNTM4P3DSUlgvWSc+IKsLHbAn4+QK+ynu8
deQ90sCqbuKWYRoGht3yDhPlxAN/TBB0e9gdw0/CN4sNdZhU8aZE6NKRq/ZU
zhOkkupBTvqIsPe+kr0ySlDEngxMgc9KBPX90ifGvWjSPEyj04wpTpJu9bwH
q1UWPYmcvsVGNDLsqX0p6ZkeHwqfW0pHYs+qh3Cgf1iRvb+67R8bHUSFPP+s
xdAiGtk/reabmySl5tdND3tXjLr93bFv8vBGVMBR9LDOP4HOzUWpko+tvsFJ
dqO44OhpvQArGdsrOQiq/c0yzQBdzip194otLTdmQfuHWaFM1kPmEFlP7doq
BkcoYE33k13t8MacBDREhuMAw963bT4h0KmnXjGWTP6qbXLVZdQzVqT8RxRJ
1zAA3xVM37ohNEoiGjuKbFlpRQknv1idWWSY2TGNEN47Ga2XgfdVGUI5NfW+
crFXFfr4f1zHSmu4v0WuhZQI3jkYWdU0JPnCbJpGwuz2rM0cQzCYdPwNfDnv
tT6twIYv3F50+YbVNF5pcJhl/K0PiGL/PnHqg+UShIgxFc7WIrMUFrPTezv0
I1bew9I55Ls+VGYaS830nBkuNNpPIjjLvNBlCy8nYIf7HIhy1PzEmPICpCt+
SxMr2gpW45MnCkDjkq4/fkO17I/TuKSlUzmKIjNPRtyRjVm/84gYzZGb9xiR
CZjvRqkwrh8+Sbft7JayaspISMnjSgbAhwXvHrHGj8WD6Db9aJA7ZuNG1mmV
VsR3RpWvyGPfJCMOIVli6BcarDbO+ZQwtxBJYS2jyijLqJueK+agEi658HUC
vUW8hdUNuauPTONXDNFUO5lUYKvOtg0UAIm+2p7eeqihtS2Lrv2lUhqrvtHo
QWB4drBWfyNMnNQKaDLAWh+XCs7S+sA51pH/48BhdIiDWMDfNBrmwC3gWKi+
80Sog/XMokMakTuvd6/O+FW/eDP5meFJqcf3uhzn1V3kgh7dwnYgyjd6wGIV
snVvVcpl7KU+/jST6rFZ7T1BzoI4arJAyCmVykMLj2U97G0q76zoYFAC+Tyc
KiMOm/WUmsO9WsGgeaxkyqi1KjcGzroEN63DGxSTha4dtD0t5ckFePzpMV1M
t/e7tQAwKpEY8GKhlJl8RqAOX9VrHjX3RKfPEiNGAF5Lo662T+d847fkEpnM
kxexorfS+FLu/vQyMOJjHpcst+tOvFLKMfs7F0cn4KknY3D3q9gr58JZm9G7
Z5lNX9C8Q4DTaHXzZY8q7V0laHGiJZWqImPweFajqKQn/uD4PayeibskNNBf
dqmTu59FGceYHhHhcDk5iExdP8AUc8QKMfVE4HmuzzvL7CTWfWUg9xHY6wwh
92PNPDKYcddCiUJfrqi+G4msSzQLOyQdXGt0PM6jwabe5TjINBQbByKR48Ce
78MNarxiWff761k7j7uGYdhJMMnptCOqcnSns4qOUM8nk2p4qkn0HEv3dfsf
ZSVg9GUVIJi5v/A+TAesXFyORlQ++yaDUrygOT7dXi4hZOS5CPd0LU2yZ7PS
qJdDZoRhMIcm1Hv20r9fMEdpAEkUirQU41zhJbmSTDVehIQUSO/8RloXw62d
sFmJ5QuiIYezCWZxj0E/ahdQ/3qsfGEcDfg3wcNuQZz4oI/3/YYkjC+mffiQ
y+BlqcSsIhMmd7Pi4vpdMPJFwvgt2BEqDHUsEtUwscZVtVDfNY84OEG4YAFE
B2fmgOtjn3oKbd2lck3+zpWkQjk6u4HFvAFEC2qZyyRug9qFB3JnzGv4711w
Cfi2i1NJ0fpEaqBFNq9lM5Qj/k4x/y/KzKFaxHONNe1fe6xMq4NL1fcLJWEX
sH5D80Rw+tZixJ15oa/3DuJ/OKP9DIPI3N6wYKnmUf9Dt1raihFpcoEjAR47
rBN2YvGqZIPks5ziJQ9jNAN2aK0Kl2KkbH8Nh7pdzf5AOJIntBAtK57pv/er
FVyOyd5nPPQVxo4oaPLuTsBIxc5bewHfiJUQ9VX40csZ+QFac7pKZJf6dbrK
75LdoK3zgEs0i+RIK0VP401IjDkWdq6tolkEgcx1a3LfgfDmvy345qN1IEfa
1m23DyDNsVahh/mOubRt8HzXSQ+oGkq2Y78QLmsxkiB0CF5wx3NgFzR1/7Or
WTow687trGwHXKXNAco4zcD6OjElNnZv+XRaCmXJDLZA4BOupDQmdI7mR6iY
GG8xWHUbEqaC6519HfhV2jrgBKkQ4WbfpckZnzxbXdWFtJ2llN3L1LxXU3Qv
6NnDiByPUAJg7LMhsL/lnzLfQHV4JMho3ln/X0EO4/Ce5qgM0jhzEpU9K7oY
sOcLayi+ovzyT1OnJshP2rpF39D5CgTxgFItUTqlPMWLhHy1G+48CLjnon33
kc53mv8OhArDHCDsIKozalhKW3F8swfcWI1DtSFqsXEsH+CxgB15u9Lp5UER
4U5o35ALUxVKMtQko4txOG5Q+qVEWRy3JHkRt8pYvwR0LhOcuV/SY4n1eH3m
ksroYi9fqDuQnz9uKwqJteaO6VhR37Ef+OZe4vHKDWxT0qS33LSd9o0ok0si
zz1NmyxfXVMtmg4Yup7isOHG4u9yVxlDKSGdJdmJgVfAdaTbcoLvUVo+eaae
Pq6uttjmhtVMefrEVYTSldqPWbS3Bt+X8h89bkAyzt0liwcaSoRF+orVhbWx
WQwrJQi7pyEiQRT+NStkoCHzSqWoQ+VIbNRVl3CdbstwUKy3Gk5wLGbaE1Ov
zXOftPGR5bwtPcVF2NQJ/3kyusVCDnjTfgmYob8GjwALy3ndctuvercJKmpd
KqKGRctN6mPlFrDyFiSBY03LlBw/wYlNlh9eYOR3ibOD3CyvKyZVMm1ZgEy2
Frb3vGQf9ggZRruLGV97DPavgmMEMHjpgiwMkJH57lLEB5zw8SgVA2Chye2f
cem8gXRw+ESM9gqNKWJmy5lq/upKgvFN8p1IXwX8Vj3vhSr1ih1CgYh1mi5U
LHfHSAqKauCo9vthX92QYrn2w0iT5QkfZrr5V+Q4+qab3blVGXAVCLXWdCQC
OrTJSWRx5Y6gS1wsjQKtJ5gSA7nhJ2QXEPIPA3qXiTh7ceiQyJ3MIr1rTV4d
7Tu6uxHTJeON4y1/XM/W+1YBuyFZavY2aqWVvifOtGQs/laH+G2dURiKJbEY
9kY+EeFRwiuxQALD7rCB4lNUcpa3XRlrKKeBYUg17VCB5Pq5WF/2wSQNaDkC
iT2grEcRnuymBi5U+8YSduKYg6HZuXrCmeVsvUCb+xksGLuQdGJxqctC46v4
2EZBqdsKJ3JykqRNfdOrLF9ajkGij+xmgLhq8H0fq1JF9EpS8Mk+4cOiCD5H
0bnr4pq6CqR7hFoEgVG0PNXRBBbWtcuWcl5t2cETzf9kfmPNF4kbNai/M8tb
tWxSFZXKoXdE0FEJlmY7sT4Ijk3mi1CeDYZtZLDhMfWZpRRqmapzWLEqkN+m
BJB2Zr+dfFbTzwnqma0QjDz00HPNThkBC+ds6KBnJZex7sbfla1j1lGz7M5r
fBI8ZMgAlXuXIcl1jSDUaJzUYPhKbkXm+kuwGukjPllfqHYNHWp9+GAei1Fh
QR9MJYGtdN9rcpVEJefMQ38nZdXck6zUn5rjZ34J89dy+FdJQYpAj90RxGmE
j51A71kQBSD7vPHwMArLysoD1lZLEgHE/SXjO4AvxVkabQTSW4pgnWvrbGSi
TrHL8/WQ3xTF3WjmvlEG8f4c39/XEydqbgRHX4pepN6YbZ8OQrCINhAIHtpm
aurvIZ+MEPWks00bVPPDevyT3DVqaUaAmvNQBH7umRiPSQ4IkK0s2UnerxNj
F0/xJBBBp2wzYyDPYOXDDMQqZrRSv6Ff9I7hemsxg+pmaklmwuPQOZkU5oVI
71jaQft+Icm0VJld4upaxhgLU2CbdG288jcda+Sb7Wiwj7ImumN0dNMKw0fe
NFY5vMAyQRbc2uErVLk51M2q0AvlFXJ53M/g9b6Jm+3se88FQrhOK4pdhJC7
lqjKKEJdWn7doMmq1Gsw4pgFcmh/1K8VWeBkH4RXOQOyNcwcKUCXEpiGS2u/
J5LL2XJn/7Ld3+vU3+0QwxIP8OJiKFyajbTU7vDoVaGlw3H+yfRt2p9CaEYl
Iuwug20JYbPIxCubAvWvgOs4CuBnGwuQUtgxB2z2J4GGA6DO/0UyhoVgcbcc
CVuLJCN3NuANQfACu+einmu3EXZf59vSRUxO9FaBJPsQuHM70VEm5aF8G5Bi
nCfbxjokb/giZpBAIwsmPv+N0hz++eQhc4fRn2OpIznx1ysUBngUdgc/2TDm
tN5yXkTDjPw99hB4JlPGFDrMvByEuuCxtj8APyf1CCLDmrk/IEqC7aBe1H7t
fi2IrTKsFVhhprSuiubYIb/PPnu0IERA2FLYCAhIoSFrc1+wqwKeZmCCs+Lt
mCOFD7VXN8oWeUMSxj9ss45/V7sMCn7W1uCI0/gCKyjB2U7j5lAn4yIoPJbB
8MxoUKv7d3FyTUJ+mENC9wkz4G4cNS1pKUyLtk8Q1/PDGTmBkXk17fQWTuEV
SoDCPhScvtZSe/5W2GBWJxk8xibZxRLELebfJ/J29baX2rHFZ7dka5A3kMXJ
HZHpY4hKMYecAtaZT+38Qy6w7YJbdKRl0JUyrHUhQvL+qW8XKLlvpI8uarRo
LBGxGP4jFxna3zcO2TbpJBDMPJZBIYIvysKzHpa1MIqeQ18jjHAPBccrckcw
fqNjXtnMXUtU132cjbIW6hSjR/S1Ma1VGcCRhSw+P/+LzhAAp87kvy2xpId3
UYCGzsTIzvbPg5L4bMP20V4m48jY6Lv5QS2n2e0c6KMmZ1Bn4hwMgmlwO2pg
oMgcS7DjLQ4f0sL32utTnvn71hBWj2wufuYWBHfeAi5ATWa5UrYxy9qt1aQE
AyEqL1QOxH9wwoPoJkyo8bxljUEyRzljiD4RgSW+slrhMI8GlCD+P3yvujEV
OHN91VBWp54acY+DfTqqdv3Hk0Aniu9vtXHud8hRveIArbTHgE+ba1USui4+
FvW12nT1yYW8XgcAAZCn79wnp3Rwb6Ncgkr4c3SpCPjbI9RgWvIu0iY/jjTc
BaC2fKwcrYtZtWIZZqdwD/vU6eotAtsNYMJjQZDenwGQ4l33vsRbueVfKgKq
5FAf+SCXo8R6ONVZ9XQEtRVKSgPhaubED7+LZU07D9PTdEdNcize5/9I0ZNV
altHlPjvk7wnnMZoJDfnx57A21RfC9lzZsDjAkQpWO3GIN98fNPGpChuPabM
yMmraABYBd88UOTL05CrIJFWMj2+3gUMkFnvc+Y83cYPgM9vY6sVoz1AYlGq
Rg9XeCgFHEdNV5gCmrvJowtgL6gHqE567ODMJG8V0x7mB/Zy4SOXAWk7aQpc
1ABmlI9W9r8Yv7DBNshoNQ0z2kz6D0iJwdTyl8rLusYb/9B+2e/5bnNx/etb
LbMEZ5w7gffGzDi2nK3YwXZBB9AYmh20NUxvq+JmM8bOHsW9jxcRxTN0SW6v
13P2ebhTYChKH4WKCyOO+zkcP3p4RfLtOSL7K+9JIgF86XxgZ9flacPEsm1d
QfXi2dYGi5ivwF4lCSt5hSyw8NE/N5qWliYQv8KFEWkc2WYCFvVwJ0K0KGG8
1UIL5+WpM1Q3q6PgTpS65cied27TSctqpu+bTGMI3psQ2uKpNDl/7lFfOkHS
KOmVtsGAyIHvL0VhcULGkBKWcFmpCZz2lTH6zHgvr3f4MeHJmUWsSQPRCcBu
UGVtRw9XA9EAxXTvcerorL4OZAN0HNrLzrlUgnEry9tpr2zzBuZwUBnT/7IE
Py8J+0/vJ3P8Ott01qpTOHZPAYL4n2653byhmJ8F7PTMI+DBcMl9nq4Rx/+p
O0u/DV/AAfNyZDa/LqBQKp97I0Wu8Ceub0ik241u7YIdTIH5chvO8Lx4HJrV
gdCkuGcOdH5o4DivG03KV+qZXmYtobD7ObsEiCLir2V0w/Ns1Gd7k5+lf2t3
s2q3sCRsyfgievxKON5xZG2Mkgc7ksgbNuEMlXRSJSB9b0MxM54KJpIBee6u
sf1dwkkYX1DBclzfG4sU7uPxMxxT6NWPOp0XJgICUltewuydW3a20XhsE3C6
HVgg4eJ0mly9rU82yr4RJvtpuotLrokndcVDvos68pgAZ8yRifk5bKaui5XX
Gtxs/xr9cbyxglDj8x2eX3Tc+iBOtAiLjMy+10Hf19r/XAD0C3l3Rz2AMmAp
WEtfSNTiKb4XIvlGHktfrfTL8lpHua6v1s6/eS7HJ4nCBw6rFUtygGFEFoUU
MB2sFlrvng8lIlH9WU5JFs55UwC05nvzBEnNFC1CvoE+nG1PVbjucqnRWMQ2
37JMHpqF/dhCJ24JS3jdPu7MMQI9vnL7yNOFmoyECPIQkdDKKlIkfjXYMs4A
NYlKD0cQz/qRn3NArP5L4bU3TDsN+yy64SLFkFgR/k86rVY8drJCzfgaiGY3
nHpbizbZ3+rmXgF+BcTbRJKgILTgFTjVOTUfX+P0uW/+LE6jpWT8XkUhjmeO
k3Dhv5qtDNeRqJADuSwdonbP3X9iw/gNP01cYGtkZDfHl0tA3aog2+1fxU/w
f3LHqoHnIgaY/wAicPv3H8X+giX3vr8FJvAM7/4mbK0MEzU1vhOVVY1390RT
1Cknp8hbdnCpho2kyjfOJiT6MPVX/Vd/7wN8Zvuk2mS4sAgjckxBBQpEZaU/
ET95TohC7MRkhFQHPBc97TFpB4wkt0uoDA0j14evGXMV9R2T9Z5ltnDprV23
sMBbjxN66tHmXzb3du5RwKyfLG8YQmxSZHQTI5JkOM1e05jFS5oARRbyXiEL
MRkDG/mglfyKuvy3oQw9z9t6/FLBTXXltYA/BYjxrZ5e4nfb1wfP86CrQrxb
iVSZ10BGuiUttgDQb70ESPzf93KkE8A2U0WH3oLmojru9vLwupYWFPbJPzkS
sZ3wiFtKzDv8a2MMjUxJi8vZAxDcjyNGBNy1lKzQWzZxRuwKklZDRqaWB+OQ
l9BNQ2l1UsGbYQZY3DFr4NTI/PBI4NusldU3qv03PCEuMTlsoN7lwybAGhAi
wpqAIoLd2Quek0AqXjY//gdPzC8BFpy0B2UoQUTK5MLH58VACF8ExHv/Q3RT
jD/tPAFJV9o3XWJmjPEmuoYv5itGSYmWA9tXNHKqJiYFdN9OmfHoJs61rLGF
JnLam6iSo0E6rNFtXhBGiJmGdny5qVejQs/rhhys3Kkx5NBtWhfAjHsn1qWK
4XGAPkwvr4IJ0Nsy8W/9rNIVTY7RwW3gFU3bpOKW8FAj/0hdY3ZTU79KWnhB
x82QImF9LKYJjXfFm0K5jyznx+VaQGQAKC5t+l7tB5G5VX/gs+Aay9p9ScRQ
CZaa81GzbMzjQy5K0PT5ixe4V+lzqNii48Cw1fmNJSrohndrCJ+kRT6uiaqd
f9wwsip5KjQ9fpj+HqC5JYDMqiazX5ZHBql5iqi5XfnZYbfdGx7Usbda+1Yl
66G1jIQCwffDIrtUtyQT4PcBy2tMRy4kfp+SdwiJboA5v0hzLlXRUCc5gO47
kUot0dZzeOW9A6QqlBb+63U7huoKz8LHMKZBxCuZwtryaxQhUAYcRP33oxiP
N419kQbtQv1hEB9hn3uRuFJOH0l0xSCY0Cl1xuKMfxcpGaPOc5YMgnh0rRnw
CJcSUyqBzazP0J5r0QWadELhkVFStcBf9xcaMQExiZ1XdOf1RncuLHpTp53G
pqFX1a/DwG0sqyTSOVvVg2vXniRrplsm8Fvkkx5DTZNKbNxvQASQOUOIEZia
h39RYMRA9d+2yZjZhzLX0La3ZMl/spz8ZK0/07qfnCaOoBcxVZ/qPPUKGIa7
RBNnZRe0ftfyL1fd8rCRU8RdTQwwdoRTqv6Ag3PO0Oguyt2bSIUc2/wHGYUi
kOV4GBLWkbUpGEg4Bb0Lg8E0YU/tnR1h51ol9TGo+d5yssVmReKX4yBID/59
tsUaD9eSyaYLL3apo3OrBS/LY6YsCibNu/SLIwqPbYmog8tFFMVnvMwu09Kv
v0Aul+9h6QDSjO2d7a2AZW9Qds6c5DMZJApgkINS/uDftuBtGotrX1I6dWYr
hB4sqZ/ItBV5z1JS3KfPSvYIwGR9pj2m88RN1uCBEWdh9YQVLdIQdWPZfHwp
4KtbE4/zHwwNdZiN9m9RmQdktkzV1NfzUsoZ8lIn8guvLbr95jJyJEnNwJ+r
DlxeH5f2eJH34UXAHryUdfF4LCM6fvPT3poFvsdLd59yj6r4ThNHtpLyDhqf
q824Jzr3jUsqKzxqDdf1ZArqZmPNNNDcCmM5rznpJWL1D4pVQF+GHf/qIRqI
cl/KFmkjq2uVxiw80yCe7mMuC4+INYmkUl1MtfzRdzXMcnxlwpSXnkRTPnve
AdcdRsLRh3zoJjK8w669JUbzOk2oxQB7xyYMW7JCfTcvz4pm9tC6dYPseF47
3OEUTolxJlj9/zQbJtGhjkyxTLDfCnJxOlidf5wQ3zuGG7F1tsl8yfnQQjBx
Y1yTk2sZwuQWniA+owdvxZTCf+vJBVIzQ3XfPMcFPZZ2LxB6FnD0jP0IELcn
vsOjL/6pJ4RX307astbN5xGMJXG+JCJB2JrjfwShM7Vif68pxe93sUlLoUNd
4QqKDc+mw87rLXXORTRc9l2vjdOFt91BguyQFcK3bPeW7G7uWInWFlP/gVhz
FcirJUnE9TRhh3J4357KoC9ZFKVX7CEEbGuT+8/PVo7KgvVza48j+HtZtoxS
MRoNJ+lufezj+TrOPeQekZYPTCVhzthM7u3eN5ihnCQMdBkqg3lGNUSBCwP9
V/hD0AXXnz84z7ZmsZLMaTenuxoXFp+VlkrLu8QI51V4Ro6WcpF3qVQLITkq
V+wElTQhZ8OjBePB++4u5QxostOpIFWh5IsB82eRJUjTk23vZg4jmV4gRHHH
u1/sdw4t1aU9kIX4+1++n8rUu22ZH/BMjjrgLKEFPlPZV/P2ZK1SPx/qAtLs
NGhCz1PAvJEptuzdGLQNpZhAx6z9Ym7l2VuxWenSqBHImhSbDUsI5sX0Ipej
6izH22HSDv5Bw8F4Uq9pvDQieUFa4WhXsn/CNGI/oePdA0iROehnpWIlLUaA
t92nqqKYC8H56WAm1Q4qMZrebYyJSQ/0bj+G0gzmEbYmxx0QrkBqRGYR3Es4
JRha2yla3VdSicp6ROf4SckeqCDM45mp4d/gAyVM+xajOriB64M1qvhupeB0
UTInX2B+yHB/jKkomE+YE3IbtIdzAjer7WSBOXKc7jTqg6yIR5JJA1tJRr04
5ehwI0Wi/K9ABgTKSczzm5usF+oXvCZROlkBr+dpRkH8LNXbEAMdDsnhbvI0
6NEK4IsodrQCgQRMfydihVXJOiZ7Q4bkpMZhdd3SpNDaOsJtrMg6QjxCU02/
JM2kZGmSBZs5i3nAeBZuG59FZZJ9UMLB6b1OyHWGSFyw/8c5WpdxlWwBRr9+
wHOtvtfJygptuG1N9KEcU6Iki/cT1eEGDoyqb1ZvwG6sEk1dD9hK7rQInFUC
eYe5eLDCQ+wMheJCAlotlXvkUw3kKMZe5B9fhaiKlqZJYpyKXtsx9iqh2rCN
u3M8gmwIo6LnSvMgbFxeEi106axkZLaRYRLRaSO4nOCJO817SDoHdIdLReow
umb4474zQmrorVNKrEaocF4M45BxUuPmEgmq8AuQzVhUlg0ioxdF0cXYGa+p
BM+Vd7nu/9dG/SWUEg16gFzYPRwvUf0XOZcFoeu6SqitBFU/Ol+ThS03n294
fgqBaRYDAciniCgu3KiY3hKP8FejY+4nBF9Q0gMZbEMZB3o0SxS8MsMevzcW
nA1fHgP6Cq2jzjx0jhMVH9E36ZoOxQB33povEfjuJcCu7n03rzY2lHnOm9L3
S2cJcAA9d+fR1kbotKf6uKmt8qnLjpowajZjKKVhVPZOUS2gEAZu+/XBDAta
9hQ9zO2mUWaOo1iuinjpDxTGYA+5Fxb7NGbvZF/sg80bHrc9eksCDGQcNIjO
hIIxFsY051qKGdXHRH96WfTdV/2ca453NcLd/1UKxDyAOm/tm9uOiqnpI49F
ePLxNhHVnK4NmHieDoPKdGGHVk/6cpNfJtZMMhnbiru1bs/YzyJ/uaXGtdZw
LRlso4nMJ4dIAg4cWNyG5rgIobSpzHwodTD/bjNNnKNBhtPT7d5FdOMtewYB
5WkGc3Owk3GBVjRn8Cjcb0AnolgQ/aki73KOE5+C6UNOr0VvoR1jpge5ntr2
42Dpgv9FW4tNfsFWDWMmLQMpXqS8qU2rcDjJLGk7++wJ/4c4NGRd2skqnlzt
HEE3VJxT+7Qy59De2lsc3m0sm25AwfNIAGIFZSBIu90eV9R8Rh6cF16EoFei
y3RRxTfozOqkPYk4i9I1wffTpiqYf5Bj52daxZU73EfBLU+lpozqZ8VeH1sT
dxO722lq3UK6fVx/O+WqvXJwmvA5wO4LT1L8TwSwwdrzNGjerPZ7IZsVR6yK
32987djDt2U8+KlPcKyGKfcFBeldEvGm/FlI0T+2wuvdf3lFVM4IvaBo/JUs
BnZghZyNkqDmmG3yiaU8hlhnO1cBNO6tjR57yf2uOxDay8gJplxYsAu5YBAg
FoB7GcuMYFZVfFsWqytYFQFBy/cuivgQnmIBh9bcZjhlukW5rYuJP+cAvBrg
K8dgCM/ieANuS9l+D8E++UnLi2MBM21d1aHCCE4FmORI6UY1KAA0DcZtLFwa
xQxx6WJqQujx9mQkBJfdFITHoPX5x3ywIn64OmJgzq18q1ImkkhplkRlLiyA
3kIoP0TCfyw0IIqBZlnweItJoZADqgWAkXKirWG1DdU9gRHRkQ/ySFgQ+rIe
reMNBEaSiqn6NHpavlhyL7obWgNhp8+inPkYfpTnvoN9iWel/2YZU6KrLbNU
Xu3lsFBzfVtVzni0FflhImExWH0fPg08AsqlqbGZcihDmkwurAu1GT2Vvjbx
r1biYVLqlX0C6YrXxUNhDnkjtpujLK0CdRTcAzKKcJ9qnSg/axXDCD2WCm6b
ST6+yPweW90v8aJiqY7Roe667i1W5pHEXAo7Uhix00LgI4FwpDU3tNpx0Ewj
FyGH5jRLpOCwnXSHN/YHCWAW8wImdIE44ZKdwvuFepiYvuWkb57+SZClndxC
H7DrPhW9stTbPGlHyu8CBbK9ZEzD3VvhfEpKV9YlA0hXnpui8VsPx3fCwTiY
tFUQ2U3uTj/DLlPMg3IFr3MAdM+xh8Lus19K2XgphuyBh996U07y7Pqb0zxG
6mgUQXn2w9tIY42tNd8QU5zT5hYR7PEUkIrZxBSTsxANHEvTF3TpxlGBgeZx
G+QHv0ahhEDx6HOcISdPNbTH4uorEPBTexR4uF2zgicT1aV7sWCQ741yCz8i
IuuV86106AcSn5wL5AJJBBIMOEmlUrs51e4wmMxIVFir8GZjR/3xdxkdkE9K
vWFAs+4kEZdWr77G9kXNTR0BRIfgP2wzVG19KB40VU7B1gwWiMBC+ndFFUfp
pp143Zz5BcRnw6IT64XvC47TsJc4SZcwTzMJ4OxYhFiYpdHv7hreDEVTS2vh
Op1k6ZmMan8rIBmg1mAVOoJvCI1GEcD9y10ZGIOA2bVi+O2ZsL/uOfbA0U3n
VWEb9bxc+zznL/sC/iKtWQ7TLw4WGqwGimPNM0+tjKVZ9ymo12s2ZzfCMqj5
bsKWSGjIDpQ1xEPbxxzEzXhsEEt6rBxvalJQFiTY8Z+NdDNIYQyZquGeK8gs
cSSWh4pmRGcIyGBziWvNKcwnQ3nBngzOVtHLVyPgEEd/rtE3DJ08Mu0LVN9V
tfJGpP9ChIiAyz8nyU7XmOLMJ0R70uP13ccvHHlxpIBPD0DwcELhPCNlB0C1
nZ7hs2y+dpHLPg/2gh97RBtrNocqy5zzPSmaG0Pu/fDkCBOvgdZ5oQSz7+40
GW52mun54i8q8UUD6dT+kY+zlsGKl903QsC8G1cKrCzJ7CEjM90QB6cP90Kp
bIZSlAongHE43WLTYH1MigC7xGQnxEhgNztKQDbRuJ0HblfUxLpyaO7r6kCw
dABc0KhLAKrCMNnga1Btl8m9TTt8XnE8wByWEtOEyOhby5XiJKR+GkLayiN2
Nyv79817i6sNwEYqxuGmuv4FQjl2BAsQBL461Hqt1VFMYtyQA4C/E32kk2t5
YHLY6bD9UlFcX1vCbQE3Jr4t6BiAA/rsblEwl3gV6dlDcJKFyH5ifB4l7S+3
6t6EhRO5eiy7DjoF4dI/EaZ4mAXafjMz3RZfNMoMI7WsgeXxypjn5A4kaCMH
rHtQu6nK2Wa2g9sDpPUjafi3Y6trXKcjxjH6J9PTNoVa6fEA9zJW1H6UIM0q
LKuiXaqZaWsfO1RE8g8TnGRRxuHmaOuKtWYIQhQuhztpuA2h3nWFPFnv/vOJ
ZQcblLNb0lXkCyhT1bJXacEOd+tOz+5tR/ZnL6eZuecaoQFUasFi4PwuXm4Y
ueLCh4hPLnDrP8wfWtV+c36HzDOx/P8U6r75r2RuNV20HOc4EkOH/J9p+ui9
K+OQCzd5/8hXfdA8ylgekNLrXv7vTOWWi2j8t6d3OKNrg3yKfY3BDqf93o1S
ljEaUn9sGPkl5qrw3uwk3mDpQDltPCyO3eYvQZdpgxNHG2gs58+iHiZp+9qC
QQLKEzziA3E+zFnGHM3OjyOBB+OkNt50iriwTXc/rFec+Phf7dVkKQ1M6IqX
qPFksiFoJ7Jix342efRhpdhY3/dYfjnFHoFsfYFgzXTk+R1fh1cLbM8Q0yYt
Tezike21xHXmcx4h8FcxAjoQ4xhLdukIqR/qt8N5BiRk6Z5JtFg06k3v3kpn
kWrnxgD9Ky/1UG17GIcOnuh5tQYU964K3CCOF8Hr6u9M/FnA+XEQL2sc9d9W
lRHR82Mqw3222Psa4nKOCHM/f4gY/4Tm/usDLw7PzNO7/0NtVJiSkoOi6v19
QOc5BpuCvb8d0dkmuj9DeFYSi8LE2ivDnDMIiVKDzXOKluVJTqZmpm159Z92
u1jzDAKAZzlZ9nEoYETQPuAPzJPGhquxlKm701SBATq0e8attZUXihxga3Bn
bXy2pLrB6CaAz9hE8DsMlZcD5ft0r6zFlb5y1LmP3o/M0EZ/Xi0pK3WloEvn
3p01o/QFRDiL+mFXd7OYvbbGCabZ4zBaRRcbmOWc22SA+FZVN32TvY6zaQdC
2LYVAeFosiuFkpFz1l0GNiv1HU/1m1HciZMBlKnM2YQCuQVbgZbwJOVlh02a
PAb6ushxJP87Hm46jpoXuWR0hDchMwqmzrlWb5U1MbRsnm+imcUlvPX0W1fR
EL7OBbBE/cIG7ZD9m5wO8IESkznyHnSnH+vkkip4KVJWU2Dl/Eeqi6AL4poM
HrAU1c6S6BIBS/7wFZwXOAuPupvaGfEQxq/HXLhufDVDEyrlBFamOkyGWJPp
AM8lzZZW9+6ma7WLSHwhlBWZdqn/npCWI395uTjkR9MC1Gx2L4erK57nx6wN
iHESU9COr2+993ZsN2mnz63uZpubKtJV1UjjKB8U7eQLQQI4STst6tt3ya9C
aYANTFpX30vEKtEIgI946x4biELgcuj5HLnGgkuW3MrEOa0BibIKnLhQvThK
MQTd+bGgVzm3Vk+ZUmZhlyAMro3ELBu7r6JZRtV3svotzgdDsDReSuC68DFg
3m1tP6pgj1nLdQkoE6jHDuRtOAzk89QRUyYVXxJAqqOXVyWLarUYgbNqjFaF
a30iWz09HiSomVtu1ptBhq5ZZK1t14oJ6l3D4er1ibZ+UK03QteLEM7lWH9M
yOHnfz5a/os7ZJ+fMd6iPS/q/kVVX2u6A2Ikym/joi/8ir5Nk/e8MCQjY/u7
iCbblqYOkSZRqspFrphrtnoo57rjgkUpe5nyGHnW16P+WFya+8GBPVZW6Mo0
w7coY2O6qN5l/eYTXfVTmFnHHqQAqo+5bQTKbQhvU63eoW9MlKQpYj/E5qM+
Qh63ZSkzAZD691BdWRO8w8ci5rEQVBM44VOTToABr5XHGXsnjMEr7QaCFWVL
SgQYwVQ3ZL/Eq5rHpvHd36dYptDWMwADQ4YxMUBZKiZWEwdXEzFkg1jYErfG
gIemhFTyQt/0JxYZv2wy+8MkOJkgGlhkAwJLK8BkxlNfnMPZKpUaH6J/GX+Y
vktO8DyHTVRhsvuBrgqIIRHIk++Zp7vA2cfrKdziZhB7aislmX57pATBQHpl
yxbJQ/q4Wk1+i/hr2T2f0Jh0yHFlFDqz8oJ4dwfm+ns9ZvGDc0su3f6uFTus
ouxOVXt7pxkiDg7W2mBcd+FoYWUuiz/pT/iN7Xg0TEvtsC/hEieiv8y0b1N9
riOVMXYG5IZPeSgTZi3WxvuJvyiPyRW7MTMg3kIhyFV3lrpRu53vYQmziDjl
QKYHw8TjaLfKGpgBC2Qbc/A+FxUo9mY9+DGA6xPT83mvbCMy6llOYKb/QDpC
MS31RmWe0cgzSplH20lOJahOfUTlLfvJURDGHweSWcy4fpDvKXWApGJaNwQX
ay/Ulwn+Ho75VO+EjnGS8yKm9vUFO0K4NaVnyCnUro3/v69Mrnd1POpNojgA
QZ9NTuRl1bvAiFmxFEtTZiWzqGMYDEoIj1UZgiItAhtRJ8VVLGzhvIxPoL7x
t+4Bt0bGj4IdCKetkcaT7E70S2pp4NYwqJmpPasQsLsjt7TTioeeWc+axu4S
GW/MRzfFGnn+iWg+O4p3NN/TBRFlrIDYAmMaO0TI/PY9uB0ytSfyowG4P4Fs
1kyFmBud2iI3mks3swbX8ft11yXiCwLrqeE/UU+cxb2MZoJcZOz5lf08Kwf7
Tunnpy+5vmLPNOrdi8Nnfw+X58JQOx4dOeKHQCofrpFlWyFtfmWYW4eTg3JV
TVRrjc8SdP0Gdyuhr9EWtGlrusAXLoDxUE2aYb54pB60v9z2BTM8nysgnOz0
Fj7d97OZF/vYVn5I7xyZhpj+FivrYCgh/XQMuiwQgvWgEdDCIsm061P3HBsH
8vbQflVeH/TV3CJ2iYdo1YUATu8m1aSCCDMxf6CMy4DRUrA2xFC+AQ8f1j1+
k8CqP2MsohLuepff7mEyyd/HL26Ie5TJodu1V3qwU4nDQMXI9kZeUNFaSW+1
2pUuukv+W5CofnZPCiRmoL6zmey5Um2ty/+x0c8jfC5pywYHzguVWkWowwIt
JCwwb1Ot7eFk9qztPSIHSPDacKHjR0jhFPbNU40HvruHE+QBCQUGUDyrioiG
GcrxXQHMCOf/6MXRahjEpSD4rpeZQoVLnXcozFrVA6QhpWfcyDTLbWYdXUHH
ptg5J7bXoQCrb3UBjcQwkN+VJao9gaI8LxNpBue8hvxctFIXGqsVJg1NNQCJ
KRDMEYop5f7L9L7FATMakQ6KQWCLZglxdfMDMlmA7FVj+9yAy8khg83m/tq3
ApoAT6NK21G59oh/WXOxVekutwLr+FYElV77DtEBGbBpjYD+if8h9L165LbK
0NWU8/D/sV9SQ/pSaURjhtgvCDGqw4s1zN53gwWX6zbujTdoTd3JqWchkngJ
4HuZb7yoeblptPtHj4ocd+LF7p1VVum1zRNjDTNPk67oNluomALr4HnZFYiJ
BOYq1X/5pAf8zo9HU2w5BpQQ1eXS3EYSoXpJWJ6yrluoYWux2CGRjYmDxeB3
mWzyWYa2YR4JYEFmBIhDlEEqA4N3/5mfOq0MUQG3McQK7/bU9dB6r07Pq0FT
/KNiUuVoXwkXlfKpDxRmI/7mKPLy7/Dz8zwAQ4Lk2AJfWxs6JZ67P0VVqhKB
GytPMQwmXJI0JmTc5I0crSoYg2V5PFztkV+KGoZbyIhvgobBrNKXGcLX+g9w
DBq6GdjsHMMtsJhjB70tSkHCyK9OptNsdni9MPT9vHyngAQQmnvjUWJnsLpV
oyRB95pUciT+9m+JSQIEu4YFGKQ47SvLe2ZfJUrOv2rIPlQcy9iBuBNSPEXv
fN4fpC3Mwq3AVE6vabygmMjiQAoK08dJ4R4iK4JmGBFUmzpf+Ob63kuDurJK
DHOf61TlMsNVHFlhA6h9Ue7Tu0ZzjaC7TQ9aG1nigMdXBvPxHKgPU4jF1MTc
ekeNERjfkIOpdja4cg/oXYs8kMxfYnxhWQVvU8WgKBnxs060Ndi3nBwlAoTK
ioLdbTF+d2OAWq3ynwAYmctwgYOhDRzWq85LKfH33nvEIcRIBASGlDHt/V4S
ZYuvrY8WlawTBy4l/d/Y/fVDGq9rBsb+wJjy3vnln5ma6RH1Tw2EjPmW6150
4rR1RJbj0Nr2+StKyFcv2N7g1fkwOQR0z6h0to/4XjgXSV/zLsK8Q7ZLa+Nn
uz2fqnB7GZ7W4PoETyT46VQgFmDDiKyBf2p778YKXd0kAVS2bGrFnR0qNux/
6tPYX8n0FDOW0OnE69BO2jhgLTJeKGxt9h1KQWBvgkUPPZZRzRsbjZwoLPfQ
p9mtquqfY1gzm6/LhVWE8E71hx5Q6BEOMBaTP1FwM/8XcLsIG6FlL99iq6UH
aNjr6iuFjQWK7xoWQQ/9Kimg+PCTgP0pXNybbsG9F2WBYc+kGNPcjgd6TWDD
DxJjxSgzj/Ib6IKRIrP4LQT9Fz3mF/pETPhDCA7LWwFy9egdqJHUTAcvPljx
0820p5RWmvgxZpdEj7Ot/CH1wrqFU8MdHoK8w3djgAxeD64K7bKFsd/d/6gx
lu7IzYRQ21RQpAT9zaRedy7h4LAkmqoaEeT6YoHczKw9tFGdGUrKtSPOabtg
GpW/XPdvMeH3jU2Y9jvpE8lYWDZSHIYJRFKDm6XSSdGcg6zQQS9aMAGVXT/L
GFUZ+wb/ac9MXXwo0Zz53hhClC1E8nqoh2fqln7GPkpIb/LZNOZaGlWpeEdT
6euboE1ObtF9sDd1qMiy5gvBccy05HnzkCE9ejnxVtA7THPAOM145JVFiLnd
sb3EIp0gjAFNLa1oqgGaphFSvCqknuemVWR0yoaHkvDQb9ykjOzUzN22UA+z
hskVt23OEyaPPilhDOU/94dTf8CXjHXmHFidJ622Il+xoJbSxCAQk/PVruuR
+/YdcuWDZ1LziKUAaJgsT/8TUxfUK97WI+p9fjHlmCJULj1DEXYPD0F9YyWb
TktzBD1LU2zUDw+INHIAU8JeK0jZA6gnMBz82TW/AsOCHbcu9speJCivskhQ
TmiYnophT76ULsf0MIjl6ixXRh0pyg0fzU/1iCuy5R7nVkFw1XsWI4KDHmcq
yexyJ0DEoajR39p0zQD5jHJMAw3MxJxsXI3IBBFL7YpCxeFs8VEHB9NtxLzK
lWrUlSo2JxDDGqFSA1b1oF3pmd6tbvCkgf2nUwEqAK2q1wry0Y1MVd4JGbmr
gjaumheNaBpchusLsvn6qJaS1a3OQtFA1qxXgl1AAEHiuCUE1U0HwlAnorRR
TJ4nmVGuGB/bGpEyZnJRfUtqpPOVUwQw9reI4A76OGMMKBGvlB2Q9LvcJOdj
/i4oeSdiKaiXdBCjl8zL14UgyJmAP+YyRa+d7IrmN2qct5rztlfvk71l9k+2
rvGySUWFFdgllObPkoKtMr1B+HJxqmCjhkRurCA1zcpFBtlz+JWrvL9+cyQs
zu60eFn9t9BL/H904Fyie3F/t3l4GNxBp4GGnWHEErP+T2pAGh1F3rQFrUOf
b+Bswojs9Jz/df7FhPNa0hvquJi5ajwaFjsla6U4K1J4AHl7zdLXH9tU253X
PNqSNSqqmiXhUM7ita2AG2ZmJvQlWa5sZhPjQNnW0xvGTwtMHi1lRvvVCndh
QiaoZwqBwBd++pkKEcE9BLCGwO9I40OJ6yJJStCrNobaJkgt3OJrqi9Hpi9z
xJiKahgaenfLkdhV/MePNF52hQqBCneeYe9T5C6E3irbOXo/bAdYkr2mC8Ou
5cMPDQiiwOPej9Kr/cgdZKG7KNbeLvqRxw61ZWoHGpds+NYcjFZRQJx6+xfK
eEH+dWpX6Tu+yBGHaQg5n+7tktJqZO0+SDP2GnnQOquYjnAGATjemeLnPQsS
SMywVYPvzv1tgRpc2S+km7bbHynq/bsHgmvfjjHiEAKrZBi/LkCEUUMyl12r
7Zg2urys6H+c/EwCn93C1F6FlTRggxhHOkRLxRyxef/Tq3VNgk4rbq7i4oIQ
HVh9hVAevKL2KR6833xYjeGLK9LtbiPczkxbL0sq26jRLnPlp/eC63ECuUXD
8Yhfq7Hh7BJUaGL+8gqSLt1yG4D9QsRIU1+rVjMRpguz1BFtFzKrIITXJheY
sbNHViORgXcL4AWIhSYjf2P9yCtYDp/g15+Ivy/fxmahr3Gfi3xwmns+79TI
UdPOCnYoC4/ClsbTmNNYkEtXSHjJGqpjRKtHYD3E/UtU8R437+HIJ7VgA3K5
CXSOePMOq3SNUXWQpTK2Wcs5CLZktnQSozGZz9PfJWrmMyOIM57+ikUl+106
j3UD07pKs1alEdJATUKK4OI8K8g+DAZU7S3PpwLGIuJgaotNzxqClgzG99Ie
jdF2WDHXaI6t7ScWYt1t9XNocxbmE2e3wlE+PzqY7OvK4b/Fu+AsLexJ0XiB
QeGJw5reL40mCd5YPvZP5ICNxJWz6mxg44XJ1nqYyCh5dpr99HX2eqRR+Z2z
b+A7JnGoAIeW30bK0DPpIcg/cH8oTvAmsv4bb21AsrXg0dLhv/GvNAwTp/4S
DH+x/ANLCyiryYc80a/MvF4zHDGHdkdK+ur5mF424IJgm59HBjJ1KnI7Kqea
xtP2e5OPFquaHFFuiw3yDZ2LIGu/xBcWHRJw6nQw2GawHAxAuNBim+ne2MeX
y+r66DSAb8/cfFNnHefAoCNsuhFZiIXauH6fZMXqBGWjwmnpCTG5zDP6KFD7
y4T3iAKoTTFm5dtPTRtzVce8KQoHWIZXn/efZVZwSdeLg/9mOoGFkw2tyezL
LqFSwDiFEtAbOP0FGJxzPg9HhxtNImJpF9Do+t4VeR8ssrnm2Am3FZmGa/cm
5rYYrCldiQUNlVOsalkGZRS0XIaW5McFLH1rGr0iphLkad0XrDAn8iJLg+aG
gyS9iBITDR5AYIzRtSmaXnmz1AwNktSfviP58G0mdc8BupVYyCW8EM2RqkEo
tptCIEXcMHUb53YmOJfGauRgOk2Lgi1MpkmKXPkdorzagG7EecvzbHi4dJzg
ANtzUyWhFNuo0AbHOBuHtj1apB6AExk+7rIxjF0Ng+0QLHBB/EgWz0xw1Drr
xYQwFuoLRO9JBZjm/NJy19vw68aRaBh3G5OtYWEvSTQ3b/frtuhofMP2fImg
1NJ9bcjvCfIJ69feUuVKdCDFFGo9arfD6yHWo+W/H0Gavn4giCGKqfgO0ASY
2PjaUJzAHlMqlNnRNLqsP5ES2YkdjrQm5O4mNrn8JPTS49WzN364cSMnc2kj
UG4rxQjjSkNVogBLQ8ZexXFIOPqNn8JNd8+GB+1ir95uzyEfzTsrjRTb7KJ+
9fY5GXcdf1paZiV4Qzwq9INlcoXVVtHj83Tw+GTQfOz/I+A2vRSD7Ck7SeWn
URyug7AwXs6qysBXG8pGnbSDqQkLIO0qyqhO24HbxnvrWuZSpg4PHoF8OsPH
LgvXNM+wibYYL0NPSJCt0/UivJz4DmapwRHBWKH9Rvo/EIuM40lWCsjC3JLU
Ff8uwyc3IwOYZgHSSBhgL+v7Hq7SYQAxK1DJRYEyecpKR82aOcy+zyLbXy7o
TPJe/bviPTM7nzKK0p0nGU/GrqbheZwpZcveo7tTRRkUouUvh7+gYfArs2Hc
1BQQp0T9K7jJ8yS5Y2QxlUKB3QNLP90T2rXOCxnbTaGKvZWB5zbJBQT/Nu5e
qvXgbcGSbOxEUH7uKB8WEU29beyM+Am97gmbnYeIaL0P8RLmjgAK/34N15MA
9hlS1zgVOkI1qhdOHsZ0rOF+wBRoNGqP12yTsStGKPTN12tlEBEbOTE6pOb2
SVheAKa3bnN7z8PYmvDfElTUQ0Sg4ScCMloxt871MbtXGI/M5xLLcaBmz6Km
B9C5GiyzxJSgbZWHekagnQO4V5UJGlXrewI/Lre0Vlr8pIW+rURc8nRcXfd5
/YHx++jT3eeHUZ3zJ/UEP2RKNnFaXsFpQC7qOkjMF4iYhMJzi9mTgsHiJBqr
EzhKmFrgtLSQg0iip1+B9wt5Gc9o1T4hywAaPDJRglrrbE/ibRc0mU8LY1/d
UAfKwoRhxurv2Xv9tsejCBc45hnHtWk/xTtetn+B76wjgi5gpKmB7RkPfLqc
T3Pq/kDcW05zH2FXhUiB0x8IEaIt43Svu19Xz9gzKs/6Hweq2rlG4lLBncHd
k8vJQnThb5BMxyehryzJNLPdpi1aP7prQ3p8SxihJzFIygYevcmhjo8mOtw2
Jcl3NwpyqeFNQV1DI90XCU/HTMp4HzHjKsHk8OyYK1w4w4rKnumIIe/ea8TN
QrVFqXgnGq/dkIg2ik68eiBoY7QrPUnwNwQuDK23JdAyDEC+2deDJZtTWHsL
onGneE8+sfCx7qFxdhFyHoinPW91PbhkVf1fX145dkzEk0XQgJo1WSY9HOqb
B4FwaNfbJftOYKOBANrB9h8ZS+qaPbwCv4MvJ7Okhu+CaU+mhxHDrwxV/bQj
FlPcTWBSUUcQ0qFOvaujPYUq3It9iUohWiB+qqqwVib1FubAXp9oi7eEhYur
Zl35h7FtBpqOj3zGhkAacrUSI6Racf1oP+eyvbfVz6YwoFKfIpMVsaMJHHsg
so1vHAXhCD2akGhfGG047rMzz/TmbHAbGgrivn45YROQpze8p0X4gbq7CHOw
q+cWg6JXltDkYVuhiUp/XfQEHzkydk84kL9rogHUVQf6QK17I625dIeWVQgP
5/XFSJySY/CzzULz3vj3QsjRHiXOEFvbsLGofeZLk78+l07tqh4eSCNvRlpR
a9dPWH2Ulrs0miIKGK0IjJ2f5MTF3uQ+i2XX4UlnAY5Ht37UA4L8+iRQ3S56
jTw4A8IQsW52jvwIqODP3UxjIENhoHpX05XnTFqcvGG9bJWQL8pMFNeKmxZR
NjrFd6QpsI/+rZznh+DhPxjUk6OzZw6l8sN80lUa3OUlOGsu0TF9JrN64awC
L2/TdEc6hKm7qdzAnb/oKKhsdnYWj8MlGSXmVDrs0WNY/wu0HBrgQ0lrv7Ft
w9NFnrRQJTDOb4q95YA9HeIk16QPVOiz/omsTSchcsb97KILyqLScv+PlZ7C
f5cuO8H1EDhz/x4j30bD4tbQ/j++Jki4JzdQ6Gxkc78G5NQ1hmKVnpLRxoE3
T9G1wvqQ40dmlwYdvjJA7kEQbHT1V5Ftr9DSLccvYBs7til0OZLBg2Nq5Z6x
qCTV9cM437ENVwDNLSMMtA5mmetwMt1iYTplDO81R+dLgpxlL4Shf6pXeyT5
Rsa3qBub7kIddCddHKbLQOXnVR9uybi4BArNquBC0GPczFvWvDxKpmFhjnS6
gdyWq9g9U0xUWqTmASK4Nb0ub3yemISKwz+TM9OE2eVrZrbisEAAKKPRsGkx
6lkwyB+/h9JXWyw4GQ4eSflVY5gfOkn4r30j/RNuyPaDfq7aFlEATy0JD/Am
KQcS8fD4lTqQo7+gDhI4XsGy9093L1oDWzoGT0lhoAu5hJK5wgfDJFq9prso
GfauyZFSTaWcIdFYVmIww08BzGXg08A4tPOeXkTLP0wmlGj0P5kQ6/rj2bJL
8Yarcv2w3/J2bnJz2P9iTjfAorZG3sBktEAMnfvHDDID6OHGf3+eB6v0GfLU
sTuNjT1D5TsjcfXUrjGKilbDgICKFp2Wwq7Q0nnCabnDXZuWie+7ARQHSVa4
9RdMLkajUhicg5bPTwdmW3a8SETghP/rI+gnFTMetWJo1uPZUD8lrBx7bdxc
t1UUWvXPGHJG4dfGkmfEPPaS4ns4QORzrZIOuVva//xlhTbF8RonU6MQZyzc
ANIozN7nQMSnzML0RD2SISFonw+osAJSRUDv94ylkmXKDuv2w7NPOPA8dLOi
odu/MpbduMY9YirZNBxm5V2U5rIfxan4WF25kmSmXXT+2Y/trMG/Rpb0hG4w
e+Lii6ncEzr/CsIZjtgoheNlnrHFbfWUCZGVC1VA3k1DEY/nH2ddzlZ78JTs
YDbQLsMUsWegLXqtCrpcPRI1ZWC5aCWUp/h8sHfu6SudwV81OzyxGDzHEYrz
axxdqPtiwCcAO/Y/MKMlLQkgWRyF3rdqaUTqCXngejJFc4PzLPDxT2oTC7pf
/+9ayIr8DzSSS1pvF2y4m6EAWb0xNOb7hde6zhEIvrcqLLJXqk50lo+CBaWJ
tMEQWZlYOFh8o4DT+wEkrW5kgI3UmI50nprTlh6FKO847soi+x8ocnBAGD26
2KmS8WEUXvgdxx0eI+HFky/nUkg3sW8v9vjvryzfAvuQwZrtWDKt4IU1I7ab
HftKfjpSNsxNHIlxbR08fjUzPEhAwV4IUpNLBVMLNAgEr2GgfItIUHhrCuj3
AzIk/6446pRex8m/tPE8a7cJzpop3ryBChVheSuUZ3FhHqvRXJHHGISeHXvj
5nvNYwHdqYJ6Fi+x0U4uYS31qH7Yq3A/1ixXKVjduS3auqb8wllzVm4+fRrq
nmQxMUNKQr85MJTjDH9NwIZ8YFbnpE24erE5HlNKg2b81PGyaIGrGJEKKVpW
K3+t6aVgzd0EpjZRCVB7jYjNXVqH0YfapXPI+h3B3gd4XKAQcbe2UWAtTyNu
05pPFOHBTznUjHYAdyyYsvXCrlPi+yVvz3dhJSfyPTqX8adFentEcZlCudPj
6w5AV10T5RiALrhuG5Uz8vmj1jPhOgIQD52cr+aSCrm3W8jAUZtqO5pxMa9T
5hfzl+ecpfay+y3k69493RPQp89TW9uV+0tvVAaEzV7YKqdK9MJ60UqHCEz9
RyOOqsJ6pyhzm4RjfanLQz01J9QngfskdzKb5cEK2RqT/dpVVyVlxUL0ci5B
p2Nk+BePWr7nbkFDKN+BcTQi33Wd2/fMCDu1pPAPDJ03Xdld2+dIvA3WrxnO
HqiKTey+himzxK6SM0nWHrYklM2AQg1p0yyOY50EjqgEca5EUVcCg7CTYoym
ji5Icz0pIhMB+dkcOO7bm5cirL1tWJ8Xl4Y+nY7I7jbEEgBoedP+OmbjSpqF
takFUeubASqeAR79MS+qiLtngy/wGg6Weg02pWPENWP8pZw4u5L++uWX8oR+
5QIDsXG4gpXCStKJerO7TUj2PMTq1EDNDQZC6nwUz1qYeYxfTAW5N0huWIoe
4pf/6QhXCI8qSD/k7WJWBT7z8yWn/misVMe4BsIhwYy+f0jYBt64xvbj8Oi0
DERi7uoQtDDsUoeoBhuxoQEC8KpnIy7IferR7njZeAdWbWFpNCR2/nGnp83s
46DmvwZyQI+GnvQZvkDOL4TUXwmkSeuimcn7KN8YBmslt+rJLixGNQ/+lY0r
/NoEB9IlRg+QnksmISoTU2ZXrq11xtPwhal6pqcWlTPJAnw7L+oiCt4hC3VK
GQ0/bIokkyou3zrzbeV23Fxre2JfttffFLCOgWj8DbtiFWngc0868Rj8aqkt
BleqS19vk0sz4KS2CbSK4iTr6QTHhI1NF/d1e9GdlUeRO3Xy5XLFIvfLJPKN
ExJosgOHoR8sD8F2VKpaUbuocJSMgiCPAUugTdJkmiLCVeIpgurYjfoJCnkB
EarE/WymkbGnH3iEWXKljYIOcLETunIggVzOdUabf9WKe2xCoxpjkBHxPPo+
6D70u9yMrjw8LFWPsYOTbQaTQ/UnND7XHH9WQZPVwQhKkRjVG1Ei3OhSnDQB
OGoTXOMZFyk/Yw0gNoKI7g6nk736RgMqAXNAtapDtssVmGeRzUGfevMk0+n0
OOig/v8gjEORfFBY1X6up3c/sH6Y32r25Lw87I+Pz7VccFq+POEfjX72gpgo
wS4vWbUulhocsiUwCY2vV5UjAfbvlb6VwuG5KneqeoafMniuE5w3c8fut/zH
qa2qvlQKEekSNeVEYLzwJ6P0onKNmDsv7vxsrM33F+umUzEmKdLFCTxMvLh+
7hiRuAnbPYTnq34b7/EMStddBP5CzTMDcBV1EIOe0rwCXFLPG32Yv5v/keWq
D5W6KqHAKwWAOMBLaDZP4xKsJzqMkQhwAE3frsauG3NZWQsnZPbZJIigiME5
zQW3uC9pfHWmuEgXq7NLukGAl9Hw1V/EbT2WkT2wuwRTU9DMKrbY5U9F7RZv
ZtAE6qAXBN3AtmAWt85o4j6mw+dfmq3axXCRA0OvrF6oegCZlXfuycnkJkJS
cBauBnUu3CVu6lCe2ZgiOGi9Wvky4xmY5jejs9oCEemImYcF7P3vx3h9fz1z
cWeqaRHkDxAHbp5zmMaWrpLu4dTzX9QbPXzpggFuqQVUTJ4ALHo8H2SfMaHq
DAyki2JgewtEJfWlc6Az4eAvYLi70MmF8epxisIVasdJDo1L6LZ8rNotvtOx
jpDIovffGJaGmzhcLN5nBDjTXTktbWdXsEHlvoHFMdh8AzS5ESw+R4CQTFuT
yv48N2Et5izZD0XNAWUugm+vtjamSGWI8Ccz3M4+nLoLdN3oLP3URwS4XsKq
HPEVVPTlXTtiPOQjI2t2m9Bh/1LecWXIjeHDuJfqkZkGGr0ItcdxmqJxIAZZ
2fCOFIiQBpU8pQpjz0MTd9D9AygfKb5AN1ZJXol9H3S+HQOrHKmUnIJDFBKF
SdIfZIfQ/ca20Z2W+uyQFhnEhwN3+8IAL/pWWS5++mn+Rk9tlu7Z2k3R/MKQ
tqaG+aufWJAipR9SpbpU/g7z0xd27EVbqgX4Fnac07Ia0hjLNff/qEOsY+gU
/lbKBMncjJ+IQAKI6CuIB2W7SxDGBMujm0c3pkbNsDU525c5OQFJ/Kb/uVc2
8qvrr0YgHFSdUeelS9KJOdRfpaov2RqXJWUbcxKIrt+gM/bn45TlpT/10bog
aLt+bnQ/6vx0f40dgpxDVYRK+iUXcFxKfC8q800f1vHsNFrMX7oIlr7TU3ZJ
3Yy81pvh2XOQHDp6zPImjMJ9Qqu5Q3VNACmP+YUlGrAqJgYCe3lP0BkEsPO3
RdgwTPGp225waEwV9aliEKfNSa0IGC/2rNFohCfP7mv+T0Htx2WlT9fzolFg
0O2QtAUWGHzRBtfaP9LVJ6lvSOOSHtWOHWfjeJ1L2NU6Z/H5/LNVhVJQsubG
lwcxXQ0sqjVA59FQTdK11vd/mDRHTucNA2aGGO9J+4jeVAY5omobUtQz5+ce
zEFh4sDLRFGYwtk/XJPFlErEWw00CZ5QRuJ9OdTzstUhmHG1hzO+YKX9nd+O
fIiGq5ZP4S/E3zkspQh7de0MJVIY00uMK2Tb3vvJD6FmyqEKvEjR5DtZaqXF
YAHdCRJ7FJFH1DbWr6fXF1mJYf5RA8j7FcP4OnAPyshVndsXYVVUh+eDVYm7
1ZL8aFnG7obzO/N6nV3IM5N4TohBbqquEzBc/sfzbTe7GYW5RbywfZINzPcF
xZ5KNAaX88BgDpX/BxTgYHM6bT7iG94QqLxT/IH9v35eD025GG26RHSdcsU7
IXaXYSOFAbvB9f7ULgknba2Jo0FpbKH0fwX1tc3HVZCsqo1oiCjH2nzCBwYC
J7dMmzJbxjatsHUYV4Nox35LN+93uPh+nvsjUBf0wDbSrNxnbpI8mJAkt6vk
6AsgkZKaqywvKEP68oAsLh/cMJrCek0zRV+phouqpvrPQS5LYETh0eyzoQtX
KnOLtYpNgA56llwgWKAhPP0LkHO1ak6RmRsWpiYtLj+kfYlRJ2XKFD1pKtE7
etxio5J/42pHrxdRQpeiJEkLWkkwTqYQ6avlT4A+WMnKUrvkYYSVrrRa0Z6b
2R5ZQ5BUoEZX91fvwbk6QEz1HGl1hkmwE+3II2RbPkhd39b+ndRDP/qilPWJ
F7eOzHepuwQgyWLEBqrckiwTT15UIQ4vfFrBEPJrBUxEqiu5fHbHEfU9yG6A
QOEtFqmu8XkcdPpsRK5ad9GaOQJdoaB4agCB7uVTTgCBCBatjzFSJZHBcui+
/SItWgc9znAvodzbRDd4NgeiW/JhmhfVZH8i6jq31kJy2QP+mx53hPDbxRbi
GI0TeOFzTtlUz5NGB9RYJ+RQfjGPVbeFCFv77WiCN5QGSwrcNS8S+vxcmpxy
eRtLV4jIeQPR07nB/YG2sXP6i01rFm8zcoHztcZssJovk8XrTQCkyk3VCyg0
X9RLkY8zAt1lQoqGRdkgh+ioxxUrgRqdGCX24h9xcAfWd5fA6RArMMC3T8C6
+s5/hJIX9XbxL6+lJUiS/44/oB4oQ/6wNfZzrvR0BRt2QvJ8yRmypeHYqnr/
a/YWqsX3MZFsKvVbNzFroV+9wmH5TnoOPXXDxfK39rIwvDe3ZZHt2DiTwYZX
hkuEMCDHJIz2Hx0Qcwe/Wo3vFGaqzV/g/k4x3ATelU0IjT/fcqgd5H+sd8hs
hljxmPr7DbP3X9FMLd/JYq1T54hFUiDAqvf9nTqMk3C65AyaSZirSC3+wA4x
pJ3zkc2vXYGEMQvjmZ5mlE0g3mTTcQ7Gc9o9urrT7uFFXeFEwYC4QiGZx6hV
FELArldZl2LiD7ZX0jDgf6AvWOYSdIF2wpCbKkdPzEsyBo73w/PPsXLwyskb
ioUd2HuhxY0eFtDu7oNuKupDTDYF9zFzbxGPKl4pkdY5yyWJ6tu407m/uvag
XURAIIkAs2EDl+Gp7tDet5hKrNx5yxausvl/Wq7AUYGam3/kJ0YLVgC4khE3
chxutLgFH+eQG6sxKyd8ZgjKjPnXkKTZ0NLV4NIuq/OJjtwSv74B2k78FqDU
FvXmzTzw4L0AZRyn9+7hZkZSunxGs2Py5nWT6yJvGB2U2dJJtEsmepMN0Zh8
quUY0aNs4c83ENHylHhw457bLTH9sActyaZ5MA0By7Xo0pIgaVMSmn18X85c
XCzHVLvwI3VziORnO71oQZF8DX6jdQ4ip0pbKvECt/FdJG1fyu1R6zk2o1Qj
CNmUDCaUGjlkj0Wm3cOy32BLIxJxUzy+AW6utq1zC0+C1uUHC8h4S7ZLGxTq
DxCvGoVbzdunsA5/l/xNMbSmYcAgDQeVA1MM87WrY8dQLLRIg/2/1u3awv7/
A/VGjHfjCxzl+eVOHogLtem8mjeSAJIMh2TdIlzs6Mex09Tw40eQxXmwFoLN
Ksd8eBqJ829xI3/wQpzM3+TmlbhQR4elYoB2nmP1DWEsrAjMNn2h+YLWOb3P
BZw/e0EXkMR50o3zXLWGxcu5FciXXBLBOj1cszf8ZEsa+IX8TyBBvXdICXnd
t0cZSh429wPoCKAu2GHoFWGFActMX92tsqZ+KVJArLq/wJ2oYwz8uCgm5s9o
9+xZxL9tHDd233XYp0WlBWkI/BXLlEeuxPCvxpU9LUHeTLC8aC5p28bllyOM
+7jb8OC3+KAQDj+q4tZRO3DEOBIkd2H/5TMiHFNBfhbNjvi+HSNFZFHf6Uh5
X2vf7EMX0qL9Y8blTMAafzidlEsBGYRLtUltBgUqrfbLNRHHLFkUHBCgMH1j
UcSnsndHu7sTsIsuv8hKnzaG5m/wJNC62/t7fu/pguv0kOTBsMKALfwPLVdF
0iE8gGQgvbaq2QynmnCawi7ZNWO7gzGcleM6i02VwPGioF7wQ6J3em7oMIHy
DlnVozHnd2JWKYXe8bsdsuGvcwVXfRQavv3adCc8JR7U2wIvpel3A9BEMj9M
RageWCBJFrJTY36vjbmwaCKcma24HQc2N318z8c7lcUZ2mN08YfyfdNMW9Kw
/sTef7b5o1Ja9TPZeqmdA3PpKkR8QrCjdjT0Vs4ZgqAGxH3dbWp0SAxpEGca
vQFhzF3AsQzh07YUDcGyKrsWDQpGUoa4EQJt4gs5+li8kVTdY/DYypjZxHOA
QykoSiibedeeI1M9vX/UZyjUb1T1YUIiScNNn8m794uaQ83sWSUPX4ys79rB
NsLEOh1RwtWTFiFco89ofOTnd7htTPnxhJe0DTTeLwk7XaF3Vc8QKCu/p/Cc
kfPiwYcuYJ4lUx5oQZZpWQLp0bHQt3cguFCDp3HHGdk3wKJPKJvxGQy1O79q
H9m/xAXCv8Vd2n3ZlOf0EBeNWpkdBJIDcWCo+bjeJpbJfOFYIUVf4GA2swyK
IqXPzqdTvQxfRrE3LI1X7pu090mUMN18jtwd8Qv0+R3JdKokESCgpUQlVg4z
ZxxkaXnb6ycvhC3BV26pzr3UpEsrdJQaU9jgOtHlcKqdLNE9htqn55npDsud
YxZg4Z+t1lxzJYUNQWWUahN2FRU8TNP6RTy0EDkYMa8qMeTDiWDN1/2EAgB+
gZTWlxqsLJA78lIjnFm8toipEo1zjtPWk1W7yllNH/+b2O3wtHEMh9x221Ph
07NX7jreqn6zv86bxOUY1cCPu+k/Vn6UT6Vxo80CZbRB+8tkSHlNnNOScw3l
pWN6YcgXFBJsi0+wIeF0veYX77B5BiqID3Xuok3pfJacRN0Sw1yFHQDLdDur
UGi81b2S07z6x+5M1iCR/VOxsrw8Wms+qkn1iRmiTupUffWxk6v9ctw2q9eX
LLiue2EhxBZgF5+IwR/uahEGc/ejhO5NCGDCCyz4qVONW1T6ncme3j1tuKxs
mFKxzgyP8Vko3ltR5cuulDwOVNNU2O5a+dQxJ+joLWQ0JjW37Ztjvdpsb0fC
0brusSRiHyjJDClNFF5f/fKfsOmnOCAk0xeAW+dbG5faSEOC4zwPEUdzuVfc
w8SHL/P10yJ3Ksq3ah5U1qFE9vhBC2bOf++wwUQKDfarJ++8yNyrftgM/4sa
3EkRz5k9GIPzlNUpANxjSptN/ao7bFtOh54TUf+8WeCkBmYzlSu5CQedykZv
Lc5KIhDJeuwHdhgUvPmXF0dqk0BKirz9rmTK4Swan76p2Jucsjg1itu4wMKj
LiHBULamCKc8cvhFroOgr82/dEO82fufNyqELg2tUaWyJDprf6cwT24mkV6b
lxOXx9QBF54hZlRmZe2jrDMMrM6MXuNn3lR7mrZp7+6Q58x+Hzse6fHRoG0W
HVrrTVu4QFgqjQvZPD1xMeE0snLIXvQ31Dh71ZUgPkQjPhNRxpEImJ//o6i/
xUKevo2DTqsTaGwCUc/pAcy7m7LgoaCzTb08bnIywlAVB4yRnsLVFK4KjaTe
KABizkdgX/+ydA3bBUlTuryIVDDkNTh63x+OpOhIHIS7Du5TZ9WtXzMbiRIx
Ka90eh0wUbbCFW88zjcTI24zYLzwiNFgQmOMhXToN2YSa+oq8h7ewacWCSen
DiKquFiCW1YUF4paso9rc3Dj9c70gTaeb17OcCNNXdDGb5lc6jlvT6+xfBHs
zfZCKzl6Qyx1CgRrLKXTPc0QIccCMsXTDjmAbZvDO/mTvV6ttozCJG/1SZDp
fUwHUqIwVug9FKFC2QHcGy0ZV2u3q4NDvn/FCb5BvBqZeBZDIsbaPTZjDNOB
VpSPzPi8ZSLdVBl/kqO1nD2ERyd/I4S2T9J243mItqWNw9u8xyzb+Bv0Kvef
qAoCcj4ucorSt/ZIfEHnoQiZr39Jt3CXqrN2CGxO/ur5ubmOxrYzGcw4NpcN
1ZWegzqVrUdNkVp2CqWUwqlivk6HNZvf+jjPXLYprgecX4WK08iwmnpoeKM2
ulhAKx/4n4aYa0MteMcCJHz5EngqjItIW56IcYOJc02PFXXl+s5Afofw9qt7
mIRi/I2Kov7yNKOXKRnwIqA6ntFh+P1YCq58L5QcyLZePe18O5vfGS24lFg6
irO1aeegliD2y8n9nx1NRix+F8DXd7GI5CGajl1HWqW5+E8wsN1yvoZHrZ5T
8KJjK7MZDWbXkZipqFL/25fE4z6UGxQA1EUpR8pNqoYJdR0rF7JlDm7ID4OR
cJ5k9nzN7/WSe5o0vgYv3EIsLzmqwUr0VeO5Kurcj8L99ju3v1yuei48zg8G
Rc8vqdOGlgZ3FLKawssJGy1uXvUbgACubjuuXgBWS/P9cITKWEfB8gJQgvMj
HVQCqOuDNvrenO/Z9laKUGLYIXHaEQmy5sPtewN/JLMIQiaEIrOq3Zp81tpp
SQOLHQwzMXNqrls/uNEWiFtsapttCG4p2aIdLdNSDTJAxASojtswCSLIBDJX
tUC7H1zOEJF9caLyKiL/+UkXDk35bovsorMf8q0edRa8IS7uoNCX/rQdDsbc
PN/7ogr1jpbUY8LuwiXYZnjFDaKgaw/GSKXclmfU/2FVpJ4KfonZxS3hrLlz
U1vYxyy9m4z0pD7icmNArQ2CkleEG3auba6IeE9V/Oa+6FcYfAaYRyoPlapo
6Sxpkvhz8MJeZRNfT7Z+rSmAlJnVdG52exjBQMPHaW6peJCvv6jVW0uJQUSk
/VU+mJOH9cOZlu9cK1HjRwikCgXGI3xm3Ba1E8h/O50WXSNebwoEYtJOim0r
3e1UKYXvbDqZdyENsII/5VDBAqJYYY4A97srRz5N24R0RUCIL+my0GPDOL5S
5Y+Q+uzOBh6RwmmzResXrm5mn07CU0oUE42Ca17+xoLaCGz9k2AwCKD3Nj5H
ElwbQfHRZWRdwnlh8UACDoDBygGF/f2yn9iFLogVz2zbD5CHB5vC0/zzE55H
75sPaGHm+f/8hmQNBCbZ1fIQEVWpKgxjkPemgNhE0OYBE7fbVYuoDUyV8Kzg
E3/lG83azgUh0slO5yIIRXGg6XICQFhggMJqP5Gu/VG0HITp8qn20NeoBbre
X1e35Pxkq0KnnIkYWm8nN2zQMeeyQOKParAkO6OuKEpGFGQB4povwb875pso
UZS6FQs/xHn5UbfUquEeo8C08Sm1IsY9sjjZEFGXNJ/Qag4u+PMxmvt9KCgT
PMt9pZfFEaxtVJNYit6+kRED03d6hi7SYoMc5v4jWIQ8Dage1KB4ekHZjA42
xXpO/UV/uLqNaHiPrw42aon3TCcdRCQd+ToOBoWXk7Exolg2Ym9HowmiyzuB
GMBSxA2Ow3L90RMmtbrKDG1pKL/TCY8WkpB2q5KD/P5DnHthw5xFfw7EJR9Q
wKSPFmClET1g8fLbWrHygRrUVqfEhpSk7lwB8hvDqCerMO1cQJgT4Ql6x5CU
g4x/Gga9Y2IETz+I5u4p6eBom961/uRYHlaFjnH2JaX4Gy2wmkFLe7K9PvYw
O5KqtzQhJ6xkNhO3mGB3nE5bUYgIAasbH0KPHOBhxOgg7zT3e1p2CGh87L02
K7R0tz5PPsxqqvMTmAB95OvNTvA//WJbc3uEbM6ML29RhwwtBR3E5AGX7gpW
ZFr+fUTzd8qYDF3Mb2yGizaolnZ0TjyOnlIJL+MqJq0uRICwUgoqYc2bbJL3
EnoilDvB9LDm88tApsU8x5ovntSPuM3lMAO5a6ydh7vx5VNRcMzEIA7LuvI3
+JTpcNyDBsYT0CgvZiTMn7EaNNj4D1/OWLsLazeBPR9A3p81ciI/nh1ZJqIH
oiAwr2tABvxq6GDoYbE57jbS1elQ9fJG+MZZ5CFwOtGcwkzgOUYbIunIdg15
UqpyXsley8Dx7X/Jgm4zsBf56ZbmWSEEAp6qF889l5Hznc1hb5Txoj68t4jj
/FVpi8d/gDcEynOyKiqfstXLAF7n/7muw/5Ilwih0pm2RaIv2g63KPq/CLLm
NHCiDuHNMRe7LcndWGkyds8zGCU+tDDTY0c8g4ixGuUFUWlAJhk+PT8Xj7BT
9oM+zREjiDbHCQ12hiLc2jOmado7cd6+8X0VJmw7Cz3uwXgldPIbKtbi42hn
cyINrs1eIfA34tH3E6E814jKQ18zfAllXLa9FaImRjKMm5qZb1N2mkLG6+F2
6sOmA0M9m500h+N5b2Awf6XnDBiag5wSLUzBHxmrvCqMJI494HPLuX1G81+F
EsD9NpNJr3PGw9ubiyfRbIVkAGBjzuyuvP+Q4+rJ7AU439mnhd98/+XGsGp4
Fz5BCOKJoR3Y1XhA1YrAW1t9Be1ISQ7yGTathkVcTbehuyDnQK2RU7aUGy52
3m/gxgZX0W03hM63z7cMLHeeG+UPUtyP+gltcUC/PzOhyxul73m2lvnOATcl
7axNShK3XTsL1UDN49mVZQcc1alLrUG4Vf3HVszb6U3E0kyUz03iIlBoHifY
NhKR6B5Kl1Pq4NoE9SHmbn3loTEQ3t3Gh6I2BhZIMV3R6C5eVXg8Vd9FK2kL
WBWkfbr/oZZlP+r32PYTx6wcE78gRm1v1fMaTdUSe880QfcI7m+GAcle5LgB
swLmIb6cRu7E34zc9VP1Pfu4NoWZd6hugIiet1vZijrLvsNnS1V7V/HIleCa
RZ3xe0shDS+WEuUsoJkMMo8kKuHNjyNeRuR7rNUhHwX+1BmbTSYwYbWEdfSH
Ayi9T3V982SdvZ1Vs/WvHrOjnqXmRsA7ATuq+mZfxc+9ksOl0e5gYOKFpPwR
vtK/bRO+lfxrUfdQ4r02zI14AybggWYULyZsqBHUADLHFe0aONvUeAiDHYyM
CN6/qLiEJIsNe/w1IRbBuxZS6FDhMq1jrwvMrkaekTxzaaCx5m97ToxBa/PN
SpG3tABPi0PQBV05X1r/KHfloziFOTHGqOnLpwywLbrMDu2o5AzJ0bqVjL0d
wYqG+BF+sBSLdz/bIRBi581DL6Rz1fKFuo0Lk1y7AcL4vD7y0rW6mwDLIsn6
p+xNJ15//th1z2dtNXavrigCRAA1mV5D6MmQo7VUEfH/bccsZ7AoQKcrpTkh
S1l9a3LUjcK2Ay6qGGUR2kn/tTzVK1kXOWA2TkbgH9rLlYaCm9oJlxh1L6ii
/QQviDGNDDTb6Zefgfjil9vLhdqwPveEjJCDIkpSHdZtsYFpLnC1NlMAZYCj
E17fgFU+Pq9RhpyIseB+UsR1+EYJoBbjRYbvux6qWIIb8K9drySe4L3k1uyv
wV3ujFPmdDAJG4olsQuRp2PapoRRBla8/gNvdmEVbDeBHvKLnoG5WM3CYUGV
QRZ3hBMZVaTYOEH5zVhL0wgXpG/OxoKNTCstWsBWF5CNElgn6ImzotiiUrxO
b1EEkz3q69yvWoKmApCINOMH41OD9SlToMt2dnAwMe8BzaTYKTpvo2ZwzkX6
eIaYBAjoCG+UzEocypwJwk/Dx2hWSis9iHGwFhVslKVNffuobk77mGwa1mwf
LeTOUcpuJvgl9wiNwxzSNB6BTyXNXVah8+Fy6tZABlsZqbK5j1R6jtOaTY07
mLnwebx3StEEAIgDEg09nnTY/gKYmoLBY49YSolW+c9QN5KHA82kyz4JTtjZ
rE3/wzUVLrCHgjZp816ouj2tNFRZ5AfcMwvgzHjZ02+mm2qmi0XaQUjBzrK7
ttYp8v0QzaT0bkQc8W4f7R1/9CZ9WtUseve6lQgG3A1yepcFgjYYQuuVFoU6
gCmAO3kYxwrMBGdJsLNH2T5k+4DMpmeqTzOd+LlyDwiH+GYs8JxL/QFARad/
9ugk9BjiN/bAHSFYXC6+sqg/csOFHi6bwkwOoO2p27ocwWHYeVoH17FeoikU
JgDUJUnKXGOwOSNDj3megb3tWanfQsXvz2IRBmD5uMf9BLwwwhoiIDsWpCsP
xZo0Rz5W3y7ihBK9TZgaEQrSfXEPpmdoUBDImxWCnSJmfTrsBH8hsMVBd6Il
UfkPXZ2ZPiA0D9HnChLiCRakITV8QzBbLkiFGB3lHMGa9xD4mGBGDdghQW6f
6/P++FwjaX/5LW+7Gkvw1Odozg5sKEM8J3f4fSHqQMlDCX7cT8FMBB2ZJOxp
gR2Kf0irnUVLt1FmhU9P0h6V60+engW5SOswbRn2VMaJfC4EwQSK1aP+d4mK
YT0zAel1uGCD4xiXYVEKHqx4Ww9Bcy/+iLiXNL/dWmqTVA6xrnKKdSGi36ff
8hLKayjy3BV84iA/f8C57KOFRMsk6c6YlJQ5PpKRmbA7yxIHDjkrRtln3jHH
xUehnT8mHip8IKSrEGLVfkVGWIcBgq6W9hHnvTq73qtnFE8MxcEFPkXtIN7D
H1Rl6b+QlRCoEr274Fcxzpjf88AxM1OhA3/bmbqm56U2sRVxCEJ9xMFV7JRT
UwcVnHztbvWb9oUlz4La3jrL4CLbZXYTGBFguJ4nyoRFJjkWjRQWV1AHwzEB
bqqk0SmfsfG/MTcFNIEllB6SU30chCgDnll1YmyQ8AO5WxXLCZRqigy828kD
vXuUaOJWBqw9QtN1VHbU7t6dlAUszTpANTee+xF9NsZdopS/XDFnfZQCZM7j
+gieFPb7CSbQN8CaWlUuquCjzfH8bVT3tgQVaqDkmBhMqfZK5r3ht5WjjdeT
0EwTIEmofavbXvvwjcS9CIcz6RtkiRWWawqO2x0GJhBeTg/E2+YsTBOLebhO
xoZQN4INw1Q/VhYVXtZOinbcb7pIWnmhhxVc08nUMX8iQA363oQtFzGlBQZu
LWG2WMWyT93N6JLLSsTrZJwmJLuBNPDg2RxIKb0kwMwsCI+pbMGkw3YM9xIR
8wT3eOHsJDoNcrKOCl9js89lDRQsK9QLtnukdzrUQUwWKSHYDv3DHPcEeKh2
vbZhEyZyO7KV6GOSaxhDAoKU7p+j9KvjWPJraBVSGKB4rbZupCYDpt6hBc8G
sNU7gbhSxTJ4d9rhyi+XytVEV8dfn7KwV7Jii60uUqqvkkmYYLMwRLab7Yq+
HcM6MCS2zWlne27sxoijSdHQqmVXdbDHah1aCVSXUbMqZmS8Qfz9LJR84X/4
3uCnQQdoObwFaTvEP0GVFcB1sJEk5vF3mh05bY/sXdNpr5e9QZ9cVbqESBTu
drlaqXSuFjxi8b/G/rUHvQB27Zv3/OVWcxQmEL9BDynVJ9sMLIi3JPaSesHD
p7Uwptt5EFtXfN4UHQpViQN5CszapDDMTFbWi+q3YRWa5pj3vtVUQ2HQTC78
nHnzaxn7qfFiXlBhe4i6/9lawlUolbp7DlxibYL6hcEa98qN+SjKBjBA5PY7
TRGL+g/jt+O76cglGcgO/29YtOrWMtMVt10DZGS3ycYRCVGct/8TS/qCXTEB
CoOU8PSZbzg1giFLEBX8zaGCemXlrMmM2RoJbpYE4S15aOLLkC4WMWTqMvoe
FXjR3WO4hilXxJfKRqPsUAlxzpUTLKsl7TckVo4rD0hLZK323z2Q1nqq72xd
664f5BkHBAOyyFRX095oNf1azRHA4BT7yiACc25n1L860vCf+DdLJonL15FL
UecpUApVPtXlJRGOQw1gQG1puz2r4Ejnxv3R9p/2N5GWgpCnpN7nAZenBlQn
BvseGR8nIRmTc5GES3d/XW2zvvGTrHf9CeHpKhnlCA1osGyHHQ0FfSKPXcdW
Ynb2/HnqzIPGeD8h9WXfXLlTjY8CmGIdyWt/lxDGaB/v+buZFvdAFL9Iwegk
W9EDI/UXj2AcFjwn6ibPWH8s7LCwZeqXFEmBgB1Pvep1TpsuajmLyuY9NjRj
SafwG/X2gA5SgWAEPJNIjVyHbs1J+vS71fAIfDcLdwldthWq6u8P8VZ21wsc
gGHogz3+5FBdPt7XlR2CPv0S5faNuwFpB0e8BqljdwpSpUGL8RMCuzVHeIIh
zD13W/84qStCxYb2L//q6snKzMvlEaumUlUKGuOXU117fDTIcMA25M1CKsfW
592QDWLbN0omlzHV/nrmSVd+1EHXZ8s8PxMrlisjyrZ8a0fsKSTX40wNk/lZ
rspOEWuNZevJlG1xPodirLmjy1z10YML5OhBn+gjo32rK7bHEKPnIYaFwT3c
04QLc3KfoPj6JHhvK1eqzO7La7s7ql9Ux0xoFw64dQyNWT5t7QVGavIvCjAZ
oSLqZ/sfv24TLWK7g24Gm8CvvcptJJs2gJii4q5k/GHgScubh+E4as7gy+At
nnk9texTbYEXapQmGvTSNV6eBcqQErY/qEtUMpg4pQeLys66fi9SoEuQXlPb
6Ga9FDm7HLhuZv1SI7GJyKdcWYeZj7SaZr1+NASs6Gbg9pptMNL+oFMPJqsz
kQzD1hsOUHCM0UZpvmiKg43PbPh5PlQrAO1nygPjo0PDln8B9ZYw1GWfOPvy
SNDQDDsUSz7QxS2zgxDQdLsVJUAKHeBqAfjh5leSkZxH3DxAaI24b/UwVPkI
ok3M7yDp6CWrS6YmEEqMxnUDDaRUdLVR5I/K3G6uVCk9MFW3GMLtDU+htMdU
FnWgloCO/wABx8+LUkEgiS5AfSpLeqzvqq2i/E02SD3wZTbFTqs4aVr7LvC+
VASVRBSxtJjRA7JrhYpNa7kQDyP4rDx8nzbKMoxx8oRZkTNOEDqD63B+IeSR
FrIUzHdDbSaCbsZWI1aHiScCoCQwrHjQeYwKEsSPaos4J4/PD3Wqa9PrkK71
Sti+ebXt9cyXXjkqG17W1+hSegpo8k1A/G1S1cDUO3K8SdsJBHlQOtIkXUml
zPTd8pd3ZUJqaZdWelDEqnati2bcXwhjDU1aJluNkOm8EcR7wNTN9kGBpBKT
CKhKYWD3RoORHK8Qcyf4K7AzXfIEYUfEzy5WrKd65LUUL8zRBxSSSEZRHZdP
Tj7HRtWaOSR83Czj64/Ouhk5sIW2mWSGGmddPU3iOHXF1fHG9ElwLWKk1Xte
0FE+BvPbH4luTtbzhwNmIuB7izqb0DPEO6Ac+DxkaQKwOw8rpSMv1Hl9J0XY
iCJwUBP8iAsGhKgZmqtzC4WBDrPqFiAHPlCCxLJZHPwqY2k7zF/LuZr8yFdv
mgk3xQNf3SLa0vGjoIRR6uXgnopJX/h4G66RCxsPf0Zx3OD01Cv+eelYriRt
kPYoE/ntvrQX3IvZRcDvHRjIEfTFGwtF5s0OcyMMDPez06n9k3rQrqC2L9jX
vRusS47MyNH3IZdnxBTi1BXGyhopO5muHfMXwJ8tzUeZIOtKt7Yk4lBOvF2k
bHX+RYEaKOFoyC6HcgaFBcyCcbq9vEx0KAlpQ088SfiZTlDZjmuuTZlTD6wf
58qalx33e1RSfgdPBF8YgqdOb2J0cSthyrH1ObOdb5d585nM808YnURbX909
RXqKkOGkdsnzAJGklwefW6vDZfMhmaUelnXjWfgSPoh5QQbuG7DTmuR6Qx0e
L8P1DoVlVoJKO4cfKMIB/+34Ag/OG+PQppxdPVh+Aa3+ty8pOngwM/Tpo8iv
xZ9y/1m8C2+uAd6NUWSQmrIYftYFzPy8eX9D6e4mANRCendP44E0LM1HVmHa
4NCHShxjD1Bi3qVAx3/rkDMiSdCUdDU1VR1WBVnM4whNPA+2ItSw/dfO0AOD
UOH/J/+hebrACZjbyh8clhDEPf96cs9Twko8C8A2ipyP2nBlHGfAyK0aTt6Q
U+qHCMmjQJs6khNtWelZKovXckC8ygil+3fZq3vMtOosTCfcEmPBnVlb6/VK
cDcm4TXbAbPPWrINCpkBlQyewhnXqi4GpEUUXtfgDvQxkJwamRLNW6ZNNo77
BDLTUBmSZbF59klwF/kmqQSWh1cPWqU/9DgXPmpFhFdjcX58Qbj9ach2cPxX
VEp6GFggUA5e/sc0fVLhJB0TUZEShnabKWQl36LRYwtd4D0WIeNM28mOqOSZ
yZDZIEk82dSoV6qXhnTEB6uGo4NhLxQup9jME1SYF4HWh4wi1UvIkjE6r8qn
oG0HLnKyaIMCRkbcedzpLGSuvsAtt509YbRlRCOycA/cIZ0jt5AEXNqEQkrz
2rKafmo/Ko6EKaEFoI752IvwVkV4RRzwhUYPtjOD0cGlIsB5WygjogJ/T4Al
H31/VEDJfVRJ3AypdBlRxqTxsC2YoDVqhavyG2X9jyp7ASmAWP7xydsjiDAD
1Bd4BJuDahP66U0q1f0AhydRoKPDUFNuCesqO0EYFLfgvMF0XxjXkxTOmAye
uhJpqVKymd6hgP+sHP+09xzMdq1RUlQEkil3ZGcB4TEJOItXhtpltfn+sS5/
XkSJv8vZc8cXSfs0JfQcXo8kE8ikR4y9FpkVWTS9SKX1JuTP9vYsbZ8p45DA
tbzkl6rgJaoYRqjTGsj6r8dWwBR8jjy8Jkt2dBwGxJ6NFeQKYgL9cq8IhjII
pGPEt0lavbDEY1QvCfVlXZVKmochA12nzobyYjQcdbxYEU9VBYaYeZM/2lHA
b8zKJnnHhnV0pa0/lh5sjFP37g1O2SLsPGGYqMAO+qHEDmFFAIG/WQHabpON
hVBLRx5WHtkQauu1rw1qB9NCQN4G2tQQIE4OhgCLjj7fAXUeclE9YGvO2FXR
xSITdwCLyIeTkZt8tUV4nhMBd0HFwc3Magt6GfxBfmGq1yJ/3mIcAZ5gvoNu
RhCTrYAivn7YNHJO0WTyOhA06aIdAO8fv5Ok4o4IzOrElVv3aOkIQkV1mi/q
YcUE30nULXqXgn94+GkK+UAzUNexBbxOMUQEFHp2SD1uHHZ2qriMUTQwCH1V
6sx33esaZ8CN6RUkokZ/i1kuwXWnpDcE/uTl0adqReRCADJw7J3Wn2cOw9OZ
xEZBYqI7TnM/OCZ51p9ms9BRHIsEqdeBlBGu+t+mj95//DSReYSI+PcSWCWK
L5lcafnlzdafU8JXVLgjKRBPAxziPkpP7/FnUKddHR0ieWSPde0sgNgjfVBO
ci51g1WK1G7YKrMAm1WQnJg0y5AIjB4P9xMgQEvOKea8tpq6YSYh7vqkdqRM
V9FkYp6BHRf0MNFt6uFe7npnzm70UyQ+974KvYbSvm9TAWcSee2TFbfuPO8D
6pCD8j65DGf32rHF4CmKWjWFZZzriykMFA0KSvQ2wn6wQSwij1bBQmnq2iGf
WcPTqebcYCvlUFKbGQytWTPSI9ej/l0mom2JXDpMoSxrotQD5UKL5v69lUfY
/e++7PtojWdi6UJjIQE14kshSG/I+cLGnVNNpSQlXbv/Y1UwW/C6V1Dbqr9K
B03p01HkHxBV0vAy/IeqrBPJcOOAGhz0s/RImBjjy0dV+d2BwSR4bwMFI1Z3
x2/QsHrULNKVTlmY7fjx17DLfdXTs1oHnlcxj7TCWITI3M6ptdQyuSGcmFML
1dFvCAEXYhpgzFfodoSaZbN9XBa7TNUdNnrIRt/wJRFgOKVvHO6aAjwZNiwb
jpwQwCy9pZWOFutPlc6aUBYHMNHOAUmy4MYU53xA5Wxz+tA7BBrwZjp44KTm
30LTiqXewUK0Qpr7LxdSkPl373bqRY5hG4aQEsQ1LamPoKsYtrrC+I4v1vlo
vOqovpkNMsiM6PCIUFw9AnmoO/fl6dbp6TjtPldBEJm9V1FdCMvHYiq5Tjc9
l9U5PgTc80EavTGjMKyn/7fTjUw9kcG9WvrWGiO4lyJGJqk0ezZNKH/btwnv
FG3jK/L95lGF91vUkki78jkfaPo5pK00AdsuOi4XAGYpIdhEMfl8y+KcmNST
kZGFRrJ7/zqsqsYVfaCjqK2l7hre5jHgfvRwOlu+teMvJX7lRKXMoccdpJO3
rS/leGMeEod4nxoImMzm7I8SKT9WUsIk9D7hgCTVw9Y56llo4wqXR9swG8pF
Q0TZcguTVuaeoqvSyqDW+h4LPjZtQiaNoCymSj1t6lKxCD2x/C29aexn3fLm
ZUXsO8f0Ke6dqgSHFByV1BRg+MyN5dK9VVET5GuK9SdvBQWu3GruIrFcX5H0
zSFvoVzvxIKNlYLE0ktB+dXxcr/+yme5j+ktMmogMYYbsaYuweIxyJp9HnpD
9E0dj+HoGtt7+HJN6Yp/4Tk9Bmw8UAMuL+2PUTLEX++6zU1YnqPOEBSq7wrk
oc5oaNjDWmRoenHViMmWsSJR1bCLvYmKBAq614gg33GMfyj8Ya8XjRdawa97
TNUoJIOFdyfO7DIf2NIzcsa/w4ieZ7gxtv8PpdNavNOPW5824pzV/pIMf438
Zpri+7KMpf/TyPJwp5rhWUWfPZcQftlLaFBYL+h8pXQH0rmZd7jyqi6hUred
17r7r9BnOTWABA0TOUvP3TADHGQ2P9BlKwnePknNYrQrJnKcMpdL6vmpabIB
z7oliXf24R7GrAEN8B2+Mni6GYM5DHMN2gAuKAvz9mzWBsjGkBdBLvcK5iQj
YnGGF2mZevek+HkkZGzIqMjW/Ntg7GMR9NhpEKxm/oXWmJq6pBhXxWmO82tu
N160nze5U0G3u5S9IO51gD/AZCVSS4fM0Xc2Mh8cQqQ15wY4qfaeeYKk/Lxo
GLbkwqEYszkI+LRhPHnzBKdqJ7PrmojteGR89SM4XwtYVXka17CymljXmz93
I6skWxBVOU8xZLCqp+9pkyVSN5q0lIjZEs/bCkX+5FHx/5PgxRFXJG6B+MwH
fPUGbzDNiIatJFWy/iH1g4eUIUw9HSGOf4hflWNG2LGVuU5nynNJJ/rSehEs
4bT44m3XoK6VSVTMtL9Odk0Gi7nN4fJQm8MPx2kiTj4SpP/WLaZJtqG70Jrr
Tz/WZth6e9BEN/cK4PnS2Qud6Penz0GcE+bVjj2gqrz/JzFfrJy7xd2W0GJ4
urJUdjXc85HsnD0SpQyKPgt9zDSutVJNU6umV3n1ppUgeDm9+lfJM1rm7AXS
0XmPUkR2D4xW0Ij/TEauGg3uZiaDTG4dpzg8g9vmDj0qQ4i7n/Pz+6LFK9h0
bXa+kFJcMbzDX0MkR09I9H5HDYgms9w6qmb5dPtk6zVXZpBmkhw7yh1CPWBV
bxJk9tylPfWU3Amw+71KfcSsS99Nx2cPqfBTCFPNkiKx9y70WiosZkXeUkM3
VzwIpnLiJQrRBAVn7F8UZqvXefFS3fYhq828zk1tFs+oQyPRtfZQuI4RmWTo
3ZU6cK2oh2U0J1hq2OxulQk7X22MluFeBGXSPrf7McwSaBsKr0JR8KUQMqf4
mtujUIryKWxCY/5D+upxhzJGrUSpZxxVV98Z52H52Tju1T3w634sD5OPMw6I
ZE7OLPF2SjalwGWdn2QsEUS+PjXHgK49IOf9wFjJDgyTbAhdC4DyZ4MbZyQn
M1XdSwtm8a05n5MvuYCKKAhwHPs/VSa9L7d0mqDitngNt9QSwrjMd5O+mMIW
dQ0hSybnPwf6O2B68QfVVKzweMtJa7Pd4GGEUOT4eSrpLK4/i0caSYZOMDMd
vh8XhvUDfobqr1cd2mYkJb7pqArL8SP3S8qC8tMz/7ByasdJ+HNHA4FUa1Tx
aGPdQujJtmvREYfR5ZLpqXs4m9qXqea4Y4h77G/s/EZUe4Tjrf8MHXWztq+U
UBxxXJM46uzFVTZTaiU1nuxVQd0SRrzfyF3MVj+AcVchCkO5hkuw16a4Sj8x
5qCMvqUOzGy4eyNpNTDpxRXEQ1eqC6lGwY32BeUI2zoIm8fZQpZLpdwufleZ
Gjxj5PDFpg6uPskOOhPGFUHoMzX9Vo+Xm0wlWtE9lnBD6F4GwRIeayz7GRCB
maYVhglZhsjitpi8YYGqwaREt5CNfFwhpZEcO1qoejqQqwOoFXMn6/ArWShJ
pbTd0i2ufXrfdkNS033U+MB2wX2hEAKCh/MlkIT63Q3c2BxDJnmyKx8t7LD3
qbeshL8vKavo14zcA9MplIqDp4AN/k/45/U36xOrQmtP/EgD98RF0NhXJOX1
5P8KqFZKr7+6l45lq+r65JqYkrHBIdfjcBFrQZPg0W1yCHby9cM7RfXKCbf9
/f5FRKbTBXeNvYvAPEVZubW/uqrhfEU2583VvEs3CHkD2EInygzIT697yQ+r
7mqzf1a1b3iSwNRWmkUXLHoET53t73hyTN4iqGV47eI7CofiZxuAWt1LlivH
iETtpgEvw8QpOIsEhIqow2IdNJTIEfBMToOYn568kGinkS2lPweZyeBARB8B
GLFN/jZGqjiaoiPr2SnCUiytEaaBD9mlER/irpMbx6l+x+YV0JiLIPy/BWpm
RHRVF9pzaLv3SnPdbOnkak32KZ/GBnfV7qws60KxL8C6CP1H4FN/2LOlr0kx
Ff/BckmrQAku8sVPH3qbAGRNQ+4vKRPsZ9ZAbgksjwA7laCD1ZmJz9XulZWl
YZzu/1DslBaqI1G5ddO9yqwSqY8MjnaPR2d+liuN4TeMG3YOm5z1CVL2zqoa
ys5Cs/L8dJD+NQr7ThzeJBwBMMuzgg3QesBBEjb62WAdF75eeMiXDKvGVW/B
M2vuIshQWQAzRastCC81OWazlRo0sBD4ZY1bWGiUMfOWJi7gR4LToZPt531Z
cmoUYyOMMBJ4xJhYRPWL7U18keuhe5T6FYE7q5BhoQHpYpqa3tMuKU4kgn0k
Gniw+K/FOCbnfsZQBJzEGQB4BIfHlP8YIH8g2PbRQQs7BXqXTpRDuMyDScxM
auX4cd66WjSXviqUgq8axCHtX3CiKvSVMBaMtO/Tm+l5qT1jCBDu9QVaSF4K
omFYY0NGkTpJ453bZUDIpqwlfjmveyx7R2O0oS9geJmwk18e2p19yHCqXndq
gDCQPhrT6N5ldoejUKdHdJGflrcEhgRKhUiCwsYhZzT99w42IptLLmf1TM0L
NkPKmNxf+B+fWhRydvqQnRI0XylW0SQYpElCrgOwTT/nlDD848nKgKRLKB3G
IVC27q+cXwDhJnxbp2U8pmrlcqGjRAuqtZfWRFbtBqt+vUw+zuVt8645uuI9
2m3D2bl7oaGFz0tUGNJK1iY91dEbkN2/4uc+dvWE6QzrZ0+JY9OYvb9k3iPM
zjWQ0h48PyGq+eA0OFISVhVvPXIyz88vZ5n5dVT4VDZ4n1jD9U45+PYgkJz+
CrPslADlD0g0q7zlhP178NHeJtcEmBG5D8mjDNHo0+yzHNW+QOW17gvrWxlx
m7Ss5Em12TasFkQYdKETeSEmsrQxHhKl0FW4F9/BaJy2+aIX34jE7gLOYk4y
E0P8uBP5J6ur4XCdwwaedJgZBGjalgS6VaYKmYUjXyKEF+qHsqw92olJhczy
rMcvBTb6xVThlbybZ4lX2reSuAfiaVa+c3bSdoWV7N0wu0hD5eIbdxSFl1bX
yGcroAe9O5Lqo39QEpTF2Cw+42eLEV/xw66HelLbea40g9Q8nhNWUM2lshLl
5JnnyAOOsLjzpPudYfb81vy6b8RD36qgEVULzyF+80cFFVEwL0RWqfjYas4+
y4X87y3F4vehXXHnetVZJj8bd9JEaBbuR/1v/J+ZmjtnyhTdqvX0riZL/pG0
NSwR5sRdqhZVM3/vDv55mmmnD6Ejqb/WtGyyON449ra9S9He+hpInmLpSaVE
P5YGAsBmK5boE64bO8u7iFU2qnP9vtpV9OtycR9rwmVOZE4kSN7Qq0o99PG9
VY610UtjUcX1Smx+LD+w1tP5VTxajj/2hxwT0nl4g5CZAUsthoGZseAgk0d+
dT5AXmJu65DHy5yMFnsErGfYAS27zJ3cr2HtjLAzbvtQqTC2ozs/EeqfeqJu
YMm6+PfC90mM/PikmS2rCX9lGnVGpGf+UTZU0+ApHmqt8CpCobQXtyKpGlMT
Ain90ULlhMXDO91t0d5nX9HX8mlVMZAvxHKTZJPpDHFgFAsBCY7NcPco1+ER
3bedmYssU88JZJwrHoUq+Xr0goAZB8r18WLJ6PI98SQNI+dTUEjUv/vKaze7
kK7Bl8c2JQoprau3BZZLQJr4PY30+kT5gDGErJAYg6JT9FZJ6TKeBH14oxCw
uHBuHpPo1cucxlMrsksqJDd+ggM9An6tlkN8ykaPTiABUUoVGNrU/nYl82CT
jf/Yx4h5R8Ba2TgPIGyThcxpapIFszaegOV0/nVzFdkcL+m6OKwiRJC+ZBQ1
ZVZMMsoP1G908c4uFXBkutozpc8PzeAv5SyowdGhgwUljLuJN7q2GSH+Jcih
lDn37YUODrs3qeSEIyjaSxNx9etUjIpgVYrbba/VvNn6w+Q4ggP4iwL7eB7F
kDF+ERS8QGsn05k67Qmf9yjOpU8G0TxZDSC3ChXdtd/t+mS79TC4IeXNKYye
ceBVpvpTqcSvYogf3PdBPrfi1HTKk2sBwqdtZcZS+znWu01gz2292V1kXGXn
kkSsI5FP2vHnLwNV6Dsef7S7WoBqwfVm3Jmje9ps7SiVlJCFl+WVic1KT1/T
kAFWPRXEC5Q/QF3Mk00etGMgLwWgB4EzX7yjI+vM5czpJo3rMKjyde74my/0
yn+4yxWgH08yhrjOQ/KbRdYUHSRH9nWJRf0Ig7QER4/53OQa7EU9ZXtuEPvI
DD+4t3NCYH+0njUOPd8ydniryUrvz7dcAQD16dgKOboUgsYUdv/o33hZgAr2
ARc3ZJPETAPcdBeAGAGf9A2kQOc9erOi2zFoxTGRHIAt8BTTPkeuX1e0lJuj
PHRPKTgyyrrUqTloJPdnSQt/5hlpRMnZXLvhwGKYJiPi4YGFniPlxV1jBUnp
ig59CG054VYWDidnlo4g7MwF+p7OzrXp/6Cj4J8Mxr86e83WAy1a9jrXJaMg
h5X9gUjMlNriEzl26i0QcQXY5AcAaG0qwkOCpyX/8UqT5bX866zrFT45huS8
Jc95DAZgTl4BpK8k5uF+jTvr6WV9u1Fpibv3g89xU+QwFle/yvOnf/CArkE1
1+xcdEnpeeD9eozE2XdSyrjt6wcGO23IruzM1FyXXcNe8mVD/F3VkI46aK+1
VmUXBfiIr6Mrbs3hpvRdlOrRTr+GQZM067bM8Dh7OpK5ianN+OtnX+77VFsl
BVCCY+0FhOY9gbDpUdHUYFuOhJffXv+Qdq9JN5O5JlbsgIXL1YJl7hODpEOp
PyabqgwvKFakzyVPAlsne9E5v67tUeyA7tfiQ0XLMO4r69g2vRcBwpTlyjVX
4rff8/CCNAxY+EhnmWYDnX0LNlezLmbSvSGjuHFbINSDIGY7A/nCyylZF8me
EBNYe8Tt/eyIO54eFg60ZgjtGIpe3ZAlueEOzjjtYKkorIARpyQ4ytcCbtPt
XQmaV5hfLvyok5uh8hMzPuy8vZNCpjooSkZl/GKH9H1Hnev6PjfdFZYKBsSW
p8bpzK+tnzfXxe/52XWMXszDDEuv4/BriM0Eq+RYZ/TkC8KeeV63zd0wtL7+
EYrlRbGKD6jaBZ76ZuYHSn9ACqHbAifOtyx62QkTacJgqogKMAfjkJvArwjm
prXLdss2Rbjr2i3f0gEx96D4KVAj7922W+xrvGonWkXOpiKs0NRgu20EBWI0
+2T3RSJ52UHAdN7byp32v1KCJpCoWibbIBtD6Rn65oDaq9NDmuUS87SUwa7u
hbMP2aJNhCogrYI50LMtuiUeszz8z5gof29ZsVORkrl6WEbhzQCSUsIRfLHE
1RCyCNlBDmmcG8Ih4pDt2Zz5uOnetptu5Nlp8ddJlIwMzLeAApB1ZYtJKgGE
+f1x9Tz12IjTvg31Qzxh+/yGDFTcz0cON2yhCDYgz07fA7U2lLAHGX28w4wz
1Sv+Dmrzf6Wi9TG5zVQS/oTzugrrt9LEZ6NvA7CiCfqNDeR8upCP5aa16f+/
//oR5F8eE1/OJeQ/TRYW/h1OQB6QgELmRUSwcpNqJHHmtXH2X+A4RFAUcX2p
ydFGuBC/SYWbm8naocwi7AYhlPU9Xzyo4hdmNGLP+3trJcwiwp3Uhv7h8Sjn
2iRUkx3hvG5zfcKvhmoLi+uKgShMPcayDxEyuy8jSudnNRGvAvKEI48qIRYt
JFqBCXM+k1Z2z3i2z+bFzne4pqx3ONzSVrBZDAV2R/0H43yEzmWGaj1uBQQv
2f68F873hqjLATWDM5KMyWRaUSBPb6OKKR/5xAO5CwqutnBsdkMFcjsBb3Bc
QO41IeDwxAyZSkBqHny4mcXJHWD6IMWh9TKYRukBtWXsQAiJWeQsxXYoc8zt
LJ4gG5VmU/zyHc8XCbKTzvJBhfRaksjW5NkLY0JvyE68QK0eV+kBqM6/1Oq8
kC0PxoIZyhitW1l4CMfD78vSNYAQij8uz4ovPZ8SPPfGahttmmSLGX+oHdjc
3i0Ed/GH9HydF76iVsxWkSxRTBbKZzctFotJfy9EAfMYXb1Dq/iOtqEtvp1V
F13k9EKoMxJPxUNTnQNm4O6udSr+CQZj7dVTOjavlrFWFFCuFZiVpnRVNXK7
X/o5m70r9i5ZaZYoOOpsNDDGwf24ltJuWmBqzDiwZvUU41Z3bTBTaiAejGvM
wvsWuJtIpudfLAANPPJdqcBIyU9rHCzlBxGwwkuLPDwJQIwHhOfzS4738ER5
0BxXdAF6iP0qmu5DNfptl01nOgp8e/ZOHL4YbAAQQL1sM9v+fNZVQygLcMW+
dTuS7YTR4oopXtSElHMqoyx+uDLiWD5DcnybtsB9ofBSpfLBL07WzRRIkpnX
G5tXHrxwABIfL6LbZmVjuAvjAEP2pdg66MOWPQGzLAMvAYmMJ1MLhHPLkuii
ba3C0oph7E7OiIBc733gFj2gCLnsZdhjS3wR8lOcY3FBW+PAmBPgomZNaJCs
o+ECzlX7Cs0u2EQvtO/1qU4RllmqOCdx58p4795J7YzBHWzJxynfs3BRXRyQ
0jyGyRJQ8isBIoDTe/pPPWXmmwmZN20w7vjIVgS/M/BwW7OuXm+R+Ii8l2ML
U7+rXuaKEkVFl56pEWfwJlvu2/c9FLwBQKWPkpdBd9AD9E1ntkLJfeEveawG
MoObyLoEfMnJwR+TJynke3Ppe95GPUCYGAw19ND7a+cMl7+QP3m+5Tly4T1z
MrH2cho7IfHQsthw9k5JzpgM0+t0Be4DwH8Uxqg+wezCl8Z3t/t0ujWB+Svg
p0VH5DeunGB78hx3Cf5xHjmKNglbAoFxxvhZETx1fBQr7mJ11JmWpHCd+bGG
W6Afs81RjwH4wl3jOpr9zeSbzCgYzAconQPXUg0XfkiGjjNos0pWRV3kKWy2
ma/nUoBQzW4VrlbJJzPKZYvE5rurBv3ssCZyvnlY7LrNxUeOGwVvmhaifjnX
CrA2kMA7MxFyIXy1FjmS8F4zjAl62MRl7LWEa7RfkNgOgeK0/sWWJ1s5Xwi0
T+eGULNkpgXBxSGRfM2c2MKydSaopKpAZaIvpJojk9foHsZcBm8k6ntrqhVV
VD0xP1+JoE+m0PurfxyEpsmzHINhSmHyVEUcpMj4d9yNGzQIi0vq5fgNEAnT
FFbRWwmm+0EnXgaMdpfxDuIxkzH0kJ2iwoUlxyR/tbD9YO3QLQnwNdULoWWH
pj2uI238zO7FTiqhN/pQ7pYB44NVjBbd7hHkoeRWkNNWl4D1TjC02u+1podH
uE5S5atEgaQx8BmeFrDIHitrQS7oFEKUmsX0V99lMOFJzQElosdzcitDAc3v
AfLMNUA5xWazfopl0FisBzv2PNKrYPqNW4deXvnbBTcXuahujpaR26Lqi/Lp
jCYHyuKPR4BKcGU6vT68N91nE/dmK9EJlxVcNVEhTTnsnWvR6j9RncaxCKeo
EJIOEfGRTVey/LnqC9Q060Y3rd9oT0nbI4jif0TrfUAAfNma4sS/dEyg7Ney
r9JKx5kgRri0PxAcWGccSggVMLM0K3JdUjiC7tkSK/upFzZrDT2VdIeTcTY9
APiH4/p8dzPC8lu+HEt4aABQAF+R5iYgSGbNhI4zLnZ9hNe7sgXkQig1nSUp
3Dg6vJ3U0HHARE8eYQKxuGJjgJK3uk22gsheq7ijum866P2r8+gVKOqVcXSd
mJ7CGvJA3uB+8Voh84pkGbAfkJ0wBVgKWedD1cd55Z4U6ox9m6N/chPXbi7X
d/n6b2DK0dsSTvNVdPK5zadHQjcndqATAw4bO6awJX6/FHu3JD4qh5tLC1DD
/5A/bC44cMCbwWsOPMR0qupkHzt0pQshXaVEbmyJL0DUN0x9nAs+z2ylZD+d
s0UjF0vF40x7ROeoSl+UJogC1L//gt0UyrNFj0IrrRH9XWzRg+ZRkNg6CmL9
eUM6BJd38Pf2UcP8VkY1zI8mApI2VZCRCLucyYWq6MQR+mVk+ukNVlADx1NT
6QYaTQJ3nqs0Ikdpr0sXV+tEbZce9wQXkouLHjaj2rrVKXh1jY5IKwos5dOy
wn7/JKHcUVIAhFtMflrgcV7+KDEtEcnHGYMOqrfK89FA0LQHilk8I1ivDmiC
ebEt7bZXyCKmRyCsEmXLB999igvCooHh12WqRBysrLAuQmTO0HhPgC9Of38p
rt4aalPqPkteSajR62VDWT/0ZOluXHcaYZ+Ld5TttskIzgMk0ZGfswQQSNI7
jJOw6grhZTKTza+NOtopUDSdpXFMD9xk+H4J4eZ9dyno8Tb8JtQOI/3Ti3k5
NGVuaHRVhICh+LQm1BGLja7IjhyaT6mdR7Euver7ns/lo/WBKIy8wT6sjvN1
7qe51to5OplCBf3uOrzusqIq+sfI8NRuQ83lqRtruM5LmY4MAMVVVanKtq7L
M0in3I2JOIdWpLFqmfjlCQJmuHNzK1n+N3WxFDwsMncbi/c7NA+1kymsy3wZ
0Z+SGd3bGA+oduhmi7lHCZ6k+Y81vHJf7oFNROyLqvFYS9GPJ2rga63/+lOa
lAfvSBH2PEa46J225s9RKQI9dKp/hJUKgi8Dii5i1Ov/9RzFFXP9+2fK07eH
DMYwxIPZU2PZA1g9oVFHcGjBFUCoW2rrCPsssNWCKxzBjX/+bdE8dA943vqm
7DfQCQ3bCIl2rfK1mQq33SpnnR9shhhQ21iNDX97PLZh02L8i9nv67xD/ksC
U3oHtqfpWC2HyU9HcgqIoHQRW88G/EMBXu9YDxz1bdSSesQ+bYM4RzQ2o4gC
kbl2+nXQptf1nSV0DZr9HGogbBDriQ9TX6ZGOGClBF6MCmL8rx3mfTQJLMXk
4FJmVKIhU4huAjGqJujyXfUNRvtnnVmRGu6h6M9LTfh6Qrgu73ynEjQy0G1q
AyKPZPdUeiCNF+TUTihFjq5sAtp3/AbHqHKWI4RdFB0eomx0DnVqgFJCo3Bg
9SvdqTqYqpRA0PpNeQ7IepsmKHn/PcZn0vFwbjpwBl0XkGJ6karLUCzZYBHN
EBKItzPSy91Y5mmCq4WUFHw0HMsomNeZoQ8+tmNtL5W334jJWLACT1VkklUh
m5BpOImq35qDFbZQ2O+4Y6CLB4DcEjU2pzkcOFP3y87zgo3Irf13VRlMWzoc
x97fEv0Enl7hX10FzvhKTKRe2l5wfahNSfGV4MOBQriBQ82+63ErbIrWPpOB
VdZpm1a3W3TWh0xC7O9uhQWvubLNWgGxXw3GvNjqhvYxpwP7zVXc5suMD/dr
hgW0c06LAldY6xbUahfERlhj4mgBBd+qlmBFT+V6jjjyIzr7rW5KSK9owWAT
9dWKe3tJbZ1BkLI8u2O8ihw+tWyNL44KVEheWAZtO6ZXwavaPBAm+eAzKLUK
qq5CDAcvCvnyi1r1ZUIwORQXWqXa6mKxyeBHZBMer8AweSLZZRlZNRrNJNc7
ZMfgj0jLx29jxcc0TG7RfLmvCMtwq1wWh5da1gMxr2Uy8J/39gY+S0OzZG8B
m9C6RfZf9+o9ENI8KqytcZOAYmDM4sW0oztFZ2Q5Q9NOODCNVvJRchOmfbR/
rHYsb9O0znNjK0BBQmVjaFgV6D+ubIrHJRXTkJqj1GEtoxN0+IpOjD3EwB32
QQI1pWztfL6zoMNJk7Zlu2H1zfrHO2bUDm3y8KZVA9Hk81U6kONHYHDiouSH
vZC97/DwkxQTJ0PmgrAjU19a6Xh+iwO6nAsi5mGt2T/Z2pce9abCgk1P1ZAs
z9EHCrbg+Gyh/+zsyRIJ8zBNdjvMV1TfJRzGCGNqnUyVNPUKeJNrl5in7qzD
QO17ZkTCBXrynOrCQ+LRSQNQM6J5vFSRjKhnbaQ7fuTL1zCjO9DxBOoDcRXO
CR7XeuXqwAsc3H1oF/6+fafNKH+ltPLxESwm/X96/fuRh5+mYTpn1GZO0lyg
BdEucD+lOFUY0pIJoU6mELPIGPXqcb9iZqTcDMbbmuZ6JtZbmfNoFRVxNGwW
eDHNWFqrKVMnf6J+W+asLWBwgmFXX9SxSf8S167AzAA2yBbQbzvDdqu/95Cf
E2jRwO+I5KQLC6CcBOPgTAQxyDfVg7SUr4BN8sTYRgBswgloEAZ4ILhawJtn
3Q71jssDHmpI+lBoknDqtw1AfJFTzJpFm++73DzkVj7O2rqp/4ePs6k4VnRr
r3iJkVlRN7lEMg2gHNJKNZlQKAqR1nptPc5WV34+cGQocL2SEn1k6ulae4y4
3WuihlgJF9M9qs8QJqtjYsjyIc4+tB/MQNtG1I1IyN3vIQ1/bUqKf5h5yTc+
X2GlFE5El360qI4vOTtkcpCqTDNHLNobwf1Kz0L+0ixN/YJxxe/tmzmukb3Z
yDYmJ1XNnjy07M8XyVQgwGXHC4DChJaJ0OlgfiP6pKRALkpzDla3tFNcBB3m
sFmRrYNGY/210wJSAh0qEXygmIgXjqPi2uxxa5fV0A4m8D8cY+wKwcGYQEgV
Stuxq2B5N+kkS7hsErSazxfTd8nQa4us8CVs/DgOdU3hiCyaLCkBhXwMT2gQ
9AwF7yJq8HpM+nbDh9N/N/VHX6BrfmXnLE1cbSDHfXirNy6y4jZBDNzI3Xtb
VtLheDHjGxC/TRv4Kgc2X1PJWu7lcAtB4i8OGgVsHRhvnFzLyL/pCPPPNfJf
VEufKxAeYPZljDOWl1T1ycoyAmnR6Yaud61SMywg5pzDNfoiiAYkE6WB1C0c
PLN+Bu3b14paLNwQCLaFwM6r/2/ZKLYGB3ERrPSkh3K+9JAAnaPPxLXcXE+X
UmEea4np/JMVG/na+YOJ7VhXz6Fn9nircb3YaMAhOL+IqufluOeYHjeQMd+L
Bh4p86inu8zhLpzD3dxqSRaaCd1Jh1kLk78uap/J1SMKdfK8FTS2CJmksXnb
Ouctdk+/F7j05QsGhNC1B1rJKGqaj0L5uyQWuM5CYBWI3A9zthYYx3oK9Ihq
ECbImh8+Dcht3MsUS7GLSKDl+SSgmRKjDVTnTNU8pcS07UyXyVoCFWJg/LB7
8weOIv9Dl+Uiqg1zoNWMrLwBl/iRxb/AYVow0lUxZkndrGhfy2MbHdB2OtsY
nLktPHb7WGLm2dtCxTP9clZS7yJTI8B+ekoRt7sGg8J6IgvoBu8Hbmefh0zD
4shl0Q4GudymXN33+kQ9GFP1fblQvshx0FRMX5NxfWtb0oVPmc+aja4w6jbg
6OGFve96gYB5+w4/pa8A2gIepCQgxWFhQzjI5B18lMC3LLDCVzipCLbKNBWI
xNPpdsAN8UCmg5mAUm2xBY5PTst23iUr1g8R1WWb6rlUR/cRN4F63nOAWKDA
0M9H6VIQb4ymtUx2kC1VRVMKpVMRflWMmgS7VjkRdK+G/g6Oe56nCIr6/wTB
JXZE4RT7Ftkpp08QLDZ+9ZZWGH7zulUFZvxxNde6Iv9g6ZXRXHpwEwTuKrQb
sRSf+nmkncONMTBipt8iWrHsG1fQNs07rfmUMbXCIo175ruQoygSMaTt7mZ2
NpH3aZPYa12wSbEzk8chpJ5rbDYmeiQUhgy+q/mVIkh1obfUvR90kRbr69aN
N67P7cIruQhpH7YAN5CWyZUy0sdr7tuljASQ8D5xFgLskXqU3Fw9h2Ye8Mfv
bYsKEh9IItl8OkrwX/KnQDc5XruTsIxGokExZL+RrNMtxVbwc1pEAPalVrc6
phJuDvPMHCgvcXwRGkPX4BPbc0cgMP2q19jndEWeZED6POhfSuf7bosGheQw
SucGGl2VbsD0ppYRbgz0OflJFtauyK7ytDbxr9EIZ7VaXhtraE6gFv8QSZUI
0958KnXLHq7X+Gr1aklS8+ZCdKQXQ87ndtnhoJgcAD15iFS7+vtV7sWYEps8
jtpZZKtWAuwpN/jd3QuvbwtFg/fbX9SLoLbYmePXnTgq+dA/VDvEpPsxm8rX
amnXARtkBrZTEAJ8xpQNxk8fqsP/nc05EZajza/gLM+tdSztmH9fnmPOAmbs
Kb+e4Zr/YE1AVFyEP7DyPlcL8B8QgPmRczUFY7MnczuQzC/cqK1i7sor9wwX
yIEAzui/3g0MDLtCfWANWq9pXUMOD8ndX8xqy2xE3QDViHjcFiSXv83VHrDo
tcKWAe1pFbJxuzcE1dO6iKI+bR4c1OG5WLYIFG3Df40kraOkVwaZv7Qdif0V
M6Lb2V1cu7pqYvlT5XxTdufjb429tnM7MnjEaPp7sALDVBZ9yYNeztd5Ke9x
oCQIg0gti3QbNoYHvhGE7tBWX1+d8weLl5Swf+UcL81YCuvMtaVd2lymPa8l
lZ3LgL9vE0fiTOPMKGayq/+nOY6SM4JhS4LgMk49Y7F6YUV/LhnlqYjTF0Qf
SNPUEWXDruZVT58WlcFizMWCcSF8WvqgGHYNmzS+9uk5wGJ2LL5qkbYHRjqA
dmR5N+5JFJtAgbs+moba2cNE/leVrw+NfaQ7kBFqp0kiR+0RsO686Ai+Myff
uytspdX50doZOMkzq/Zsy+vciiqDSwnsSUjVkTMAQpr3eF2po/0vm12aYsVv
ur36OIGHN6KnRzBwQaRbnEvoFgtgsGAJF5zHu7z4Gk08Ix6AWrHvMmcOW0Me
DcBebOXtpUT/UDroYh5dp7XY4x1suDnJev7/J32W8l7VYs4ILmX6Pm3rUOUy
8+XB6bIB/sUGaoiVP7jXjIZwJGwSbhci2kKhZRT/0bwVFP5xnmYQ3HtsNFhp
JIfBx5j97/Fu/8g2x/fSPvLh6pf2d8vJbdGqhuOwvAkow2GrOE3v7U9rzQiF
K94oDvseynPf/3RtwQEGKrQm6gQbt+ZqreR4FBdIMAjKk0qoArQ5N3jH24e4
NgCMcjimNZAk5jcZTzBe0Tf/iYtZ16R1xUc7y7+e9a4qzHT8l3EK3ZjbAHr/
icKPNwpD1QjsRUIoP19YZzCQA6cceVipuYIPw4eDTVl5QOOrZkeLBb/5id5R
QHV15WQoF3XT8Ag3oOkw1zqnMpfvX0LjbkqCuruyBTwCnX1vTjXhHMDbELk+
NeEcbLPQTjH4HyPOnmhCH53+zwSG98fGVuFxJcP67S2DEKe7WyoZEVtGx7AU
ehyMWM4RnluEdhOo1Q+54SA+YwRcf91+ifJeaY3q+9KQ93HClC8x4VCF9VVk
dfoykzT8rMhp5wk5TwphtjzCLMe14kTLGMZt1JKMY7vzoQlgFwpFRBdcvl3r
OYa15MWV+7i1DJ9K5/6NAPvAHgCYjCy/SHtzsIMBnRtYPFPAjAWXpvsF6veS
WntN/dn87yEMZJKnXqd5AIs8THcJ2zL+DFAk1qECpkqLGMS4K3vEyhKW0xvI
FeQy8faEbedvmiFZPANozew0J/R1NvmGp5Vox53NnvEFQm3WmZKGLofFET25
LnJ2ZN+2vnpBtggM/j4AiVU6zwk3bWrov2uZviDhBKvXEYOG8DnuvwW6hZjM
upKX5MiDAysNEYdrhIqnIIGelntQJuR+tY2CG3qFquylIqkDDePydgZzNbHg
1z6t1dCeV/QQ3q3z6HkGQFo4onysDPNLBeUjf5/z8CBdMOdMfQalC1FZsLb+
32uwb2QCNjAUuTaaj+gg7QnA9do/H/sZRoIMys+JDGga72sx6upzSbFrHqx7
BPVHBPG46j2A2LN3aI0/0384rGRwv1gjWfRZp273odSaM+U7iGVV14yAZ+fr
YiT7v8RlurLuZN9OKpFlvyM35BlpnYO6IN4wR1DjS+J2FTTDrssRyK6cGsq0
q/gelRzuYmI5Eu7siHl0SgbKCixe+pfUbzBpyvpwaRoLunrfzo2POX0gk155
25O6llJntILWws8V0UIlSIcpkgsMBR0bvz3sZcNGPwod4w0fs1JCbjjVzbQB
askUhmNaAsfayza/PPmdK33UpaIfLuGK9/1p2q2c3VfUpU9rImbGOgoW6CeU
c9V0Hnl1iPqnzt7Ke7pshiZ2mNBZH60DQfZotCRE3s2VmeNP6D83mfxmmuNg
ijavM4zcYeOk8UGXcSLuH2zYnWvxSuyedZr8vX0TlsVy+h8fGXzd6FdBlq9N
7l1IM+YikwAnWlbsMRt58Ws5su62EePfMppfc4s24zH7DGxvunetNqs/oCE6
pOyTuB1mFZdULuPaeuSNlWPUPOduafFcFiwOMkvSbQo63Cb3lffSB3qq8nKS
Y05NnMZWwJzits1SMKcJFrQ+eF1hA8B4AylL/DSgPLHcvu35M7RQ1xmNVOey
d7azS8lEMdOMDQ6G+qEkt7YUUEeqMnwLvmp3zboRNzUV5ZKL1QHjTbsXZaTp
1aHtmri9C33bF698uGU3efXvTXPKWKnHaQjS+iub428j2iIGiKt9jaGKaJDx
KPrtAOOdUkkh3TB6DCBZV3zBXx+cecb4ACe+POX/hsk2TN1QUCeBQqhAvnWL
gTc1UNaNc1o1yZmgP3Nz3kLwFQwH5e9rDqVSuvsD/36XocEOD0Kh13RYdOIJ
1GirD4jG1ugCYdseOIOSnQL3rZoqDEleRUAlql2sJPdrhe1vRebzH5kJ6NUk
DLemg3pJbc505NPAiso40wYWLardqnJ5ms+wnRns/e+fs+bRzDQg+mo7ErxD
n3ou5GEYItZ6YTlH70fuUeSEeaMWptafWVO+riPjoguv1INvaf2hwNhU4rVy
HST0hpvLDWixrClKL91F1yVIvdCO/V6u3hlxPUg3zu3Ti5ikHN1hH32O/rtL
7OjCY7DkqXMA6dlG6EmDc3Gaqx6MIL0eIhs6cYDSw0vpmy7DlY+lgsZojDDE
K201N5o5tM2JUj8J/2kvGuSwyn8Sy/XtKLMF6gONRdKqJIxSgDp0lQlLtUAj
PgvTzA3JEjTKFUr5hI/DznX+/yhdsmYi27hTExvlcP4C4x5OLPlzgVKjYb8p
wfFEIjLFv/+bMdBnlWTmCGcoJvYrYlgF11fc/vvtiL0ojZMKw8VrIpyfYWrE
bGDKmrjvz8lBrhCqKzkM97AJjlzonWq+o3ttgQnW0/ZZS7Axwbt/PG63uHvN
rOYOskluivRx2TQCIXw3PuPIJx3tOOHy09Vv4mq3bZxlw/Xy4Hovn1gPeCMF
u5CQTiIB/GBFXghblUhoNdMl/1hIHu89WsN2Brt0UzNYaNbfNAHRiQ8Ssm6C
d5DkLGdnIwXsn/aOHqK1zP5KJ2lmvDnKlYnMfkXnIVb96lnvER8YZpZdW6QI
rAR9ZP295iD1tI6sNNH4IHloCvDZl/d7ZFDAjmVgizEhZs+F4VmkWS1IHwi/
oIBeytCpxqHBWtQmq+EJWoj4Uaw6QTlh0RaDdISKFAKgKZ8YHoQglca2rThk
QDdqU3sWR2n9vI0Yu9iW2lCkDuf5s1n2nV9TKpCKIcOmL3U3W4DtP2d0VEQz
PwjQm1K9M+WYV6NekWW8QXQkEy27EP4EBotRdpbXUM+mkUYk35oZqenUzw9Q
wEu5IF8IAFyw83q6VriBucYLjgiOk8pgD6xK4+QBXRcQR0EnvLBmddvVyu2U
3xyTflsUytr2nNb+SxJo1we7jLmfSoBEBUsSSitgovTy/wfCQQYf8mbDDSql
58pZcVII/5MYhF90TegCGfzF0k4Uy/JSNm8uuB0IZk0GJaXhEmx5QFF/Y3OD
gjd9afiwRpHkb4amieZTiPUDyt7Gm6VLqQAtkesJHCldDA7yUu+m1S0YHoAd
AY1hwpkUp/G3ZsK2am9lDHbYeMwUBRL/hlVRRYBZdUOnJaNZ0+8s8qkhagFP
VJOokdL50LlyWSGuObbhyKB3KG9Gtyg7XgWFRIeZA1oy3khRbnhNi9G7JMTm
HIpdb9ZGvWhGfWVzikNfjNyfFhqmzaVGVBopsRJV3qupAVLz98C61Lo5UQVv
zWGLCk/0qxudh7zUy/m1dh6f09QhHUHyOPIuX6xYrWnQ1Og1maSxfvhil+GV
lx1XrT/8L+14uN5jJ5E/C9Dw+A+qXwriaHytpNe3UQyE1uK9jxTyfP/9EY0O
3eBmEfC2LlGfP83PHfNovD+d6HzuMaOz/6xBxwbOFpL0v4wkgkVX0cDOWo5V
7bMDwQCKsQCUmeDNEDhW9f5QQduh+kCOD71bG0EspeWx97Jgt0YDSWQjk5EJ
W5h7F46ZLf4YNnlxhlh31CGFEcuCImgqWkaSpZnq1YAvGJTGGaIIA2OcB0vg
59wu5vF8hTkhUmINDXfmS3c508JcW+G0TJF2U3wdR0YDJ5E/FyloaFcU+RZI
8+TBo9RKV5PrlbAYTMLBM8uKB5FA8iiwHhCpsTjwqRAfWIX1G0v+uH49CfGF
rB/E1/dJ5yF17DB2Tll9tRlr27jrnmGFAl63Hh5qtOlTR7ziZy2aTdcBHbpB
DdPIGYDt1Km7I6NNaImgyh/68TaYzNIaRGs1hXxD2QBcG9cFvBid7heKeaTM
bHus+q8LD9unxE/8/TIhznE8bK7ps2LWsjpByyHfFwxbFmzPJTygaEgf2zCb
EzCZGQzNTOQiRFdF+924h8LhMDxpNz0AI8MTqjbXBkqB8HY+x756cC+aKI+g
7qBHhc5Sa8wQrSwoTO2jDeBDebi+If3or0YZV+JV6Lap38W/3FTtfmZscTiN
lWh42LE2LOeqHm+uk7yMkq+GN9/vdVhjzqBJdebb7tR6Xj6CD/Rfn9AlCfaI
voopoW3ND0YyNH79bPPrzhBgxtF+p11qoVnjy/YejDlwtTKn2Jfyn8fc5geS
XDaO+ai1/JVTcYmqRBwKgwJRmXc1kHG6gAqp+HW4lrAeQ3WieO6BOBA8QENF
1M9DkWTX4k3c1d8tkaH7DMe1qbn9nwaKzVs+xLiE/+E1O7rg93DZbumopHL7
JJji2jr41MvINxFVxPXE9MRDeEkD6UJLmubHvIYOqBUwAYCI7XOsU4J3+ICr
I9+njMwPP+iT9FDtBlTTmMFSXhDt3zmYX2hCy1E6s/MVBvKDjwCucvCpPP/p
SXBtKDTeJVg0+yw/BrOHXZa22kOTjuIg2aYYGjecqaVXHje4i8YqnVy0Ydr5
lZDa28JqviKCldfiUOf6IZtBtG1xTpfn6Hguzh01Cm9yGSxaJbEGW2gZ+aJA
xc9q7sjdaJfeU5gW+ucnRYajdDI9RgObgGrhZusQloFYuwb1Wk+riAyIXwe8
0XF5Ay+KzdsbNiSc/YcK6UWO4WDIlHeO/q7BaMRj+C+2Mfa2nhTTfGvyhMEW
+jshxi9JceJXoOFkN9e49+XWh8niBVbarSWEeSUlfjH3J//om20GFtrxswur
NvoZ2a7YCTxBup2qcoHusBU1Acc2kPowT1m6p5nMpFlcptU21p7QH28Hq4Ij
38uqvr0/YxZdhoNgjnxKVQttDdTlGpnNbZgan2O9hgfcy17UQcIlqNbve0Yl
nlBQ9glDfgSB4Okx+GGIPiFKZ/hrcsqz1XUKa2STgeuCBAOObQFRZ/87diA3
ZVk33gcW0Dxj+PHiTR//4wDOReOwNdE3J79b3gllLT2dG26uVCoHCoX8+9e7
e2XRze3g9g6le1oYH1zcXlv9jTnbiR2fObXBzeATQGKVCwzC2OP4z4w41LIn
3Vdfz2T432N54q1Rfe+U1xlpgjJOrRmXRzhc1kG/QEiw0le2hmGlnYrCIGaR
sYjjdrsOlGd9pajIyWY77KhjN5h8Y3yfdopXTBpuWmQFZqi7vmPN05v/Kfj5
ddoZ9+hL1bq8ngcL32pYhv9FcdSBMWJUiQ51/CeT+MHdeK9ZIGNoCa0eaLJe
Urok5jbsboBT7FHgU2X3IYV7zFJeZIVkTekfio0fK2JeP0xm/u+ZVHI61ZOF
8f/nxe6IxwmiyfR7khswgoYqGq8aAYGas7NsZ1lm24rmFOYCs5beK6X3Yyib
kOyn9J+k2O6y+g3v5dt3HC5a9RNgj9oBZbhJy/Q/AAy+hywFRyZl2LSZs2mE
z1hL6XPIiIYrbt+oQWloYt5oHA2L1Gx1sqY9GPJArnqRKRPEoz7DwY8UVHqL
HNdXZQHavaEAEzX8zpPehhu4PFOiUiNwwrIYwf0fr1BtlsaG74+UPrLb+2Cn
IJpjj1UzwNG5qd8DgE+HwRLpi1lgOiT11V+XJ/TjbcEIoAco5SRH6FWZ6+qL
IJV4Jc/IBOH3Dk6Fflz3SDTdBUZt+nAzmEQVSKShB/Z9+p690cI/cTt6mil4
losn8W6+Dei734XiZ5EvNHWbcgOtTyUF4RYLFXyQOGukrxmMTEn33OshMGR5
njLyMds8dRMB9liDQUoM4lyqk42f4PupSjNfXnq678MIWXOgEnFhh5Hgeqej
/Q1ZEfWbiyorQb1M1ghoPDGcaLlzUdyzArBsJ6LyEb2jIvsEogyXIJ12/+7V
LSg9N62xva2LEizhYYN/6LkPssB9NWrOgnf2OxGIH3a69IMiEAV3OzO0gKOb
YuxgAh7ftAgFF4ZaZMKivvIJG2vQ9aB8OJ0SCkSUB4P3YtFkDFi/gn/6bOFo
XGzjUBFFNn9l/JqSiUZRWDHbXmPIqyvaSfya/WtLE5qElgMa+CzCq9WcIZ+P
tQna/vJz+rMAt4arglENg1YfK/foyqay6DdMHbLk4vkvzquiNDQ7kcmpq6N2
f/qWCvbesvNJG2cLPHsbL4OI/+ELM7u4s0MJy6GM55S5qevxfoLO0cECNsec
EPNjuElseCHDTHw7y5RIRu5oO8md49GW8zyb8yB3qL64DAyFrCiIFiqXcTt6
teZLd8wH79dUci6LXaQKjTaP1EuQCsYAInkWV4X6TZAJpVGoVQvJ+hsI4j5+
S9C1Xv9Q7r3v6+e/oMsDCLlpJZyK2/UcgxTuLI03gWDKuwJq10E0668+0IO4
SiG/wf4Bkw89c41vctYgUyNQoMSdZ+w+ZglzZvb3eweVCbasHnSxvTuShdTp
ufT2HORPFX4hZqrX2s8/uVCeWpkXFmsgQCz9RscbJY0ZYQiLFawPhk5T0xOo
CQPgTKIGLqf9mChWH9pInhUqrZTYfIH6GqMWAfJjctXgCqOtvhV48ZHf0JqW
YM4JADYkg7FDTmIM8oocoOdaDgwF0lHRm4biVRgrfxgLLE6SmIdh5EX3g3PY
Ax1DeRYDBIDA3EwxSxf7Ad1hEXWWehNFjQFY/COib0wZcKyDlON7pmYoXVVC
Mi3MziYCUAFTKhSYeTf10rFRo+KfNWdh0sw+neavoN/LkimAYTogX7ZHXKNt
oqtWOETxwKhQnyLBwm2dKkjTqKxMZaM/Fs7rKtgIcAG5yu79v4NbZcJ9Md2f
u46Ywd+Zh3X06wLFc5SbBj8bCLCocNVmjjtK/8FiVEFYQt0KHR5AugjjzQP7
kDEmHa8Tz4pTHrlEdzsyDopHtlaowSoRKoUo96uCc24aq05P0oCqGdxj2dd/
z9a/+/qltEDdxZKLLEaBmRyFwNrMDz3XPSQu8G/LPWr89GIWOJlmdJH4aCH0
bgBu29JE4zJZAzQn2jX3G1cixY1FNfu8xgJpZGVB5tJ7vcr3mwiikQqWqQ3L
e9oRoFdjHURhn5pRA3pFuWbg6mDhugrfP/l5H3FBhHmollAlsHQyAEsW02UH
auG9D0lovPh5T6Aw2dob/uvULZJYY7O7WA3HNWIGB7XjeUL4alFZ1n7azKPi
TYGJ39fPrGEQFf9QbMxbQtg3Lm2GT4bZo7HR+ATSdwNbYkGfwJI9LgW8kw/A
xQg0ENB5mN3ytCMbLnBixuZnExeW99dyivelzVPTo25cPsomOwRALXouRRvT
bD7EnoHoFk2WLS4qhJRbcxToElTKhAIxdSCpMSgFgmhiMgM/CNT/H52S3OGP
zMVeaC9n9NgOQepNELNxtmw/CF1x0+253dlIU/sMCUeBkpEFJI0EbYKe8u6S
T45sOyG9KW7BcmS1V3Ro6mW9SfWLWM7+xAiGKX09lEyypFn6FSdiEyRBxk28
kzewmxjcTbXklKMuTdQXlGuR8hiotUBLWNh7YJ9u71kdPCCwXRA8bq8PQWol
HGLGLGWt2Ykm4vfuS6hRn588szl0lp6I52YMI/38RALVK+lR1jY94R7c94gR
XZNN5p8J8XJZwa4e3HmYCXcC23b+mVyGIhNDodJ/D7UstmPQyoa4ouYRjyhI
mZ9xT3d4lJNNu+nXVm2x+6JZLTK9xGGfZD0Fl81WZlsGP1PeB7LFettNLyyw
I/rb+SrBe5LJUlZ7xrrAG4RywCBmZcj4eFgAsdo5Dq4DIk24w/r8J+3+oMdC
pRrphp0dNuknt5i0GzrlKBUPBW9+0SdFeBSGioiZ2CvceqGy/CR4/SHSYZdJ
J7qd5vwn0fqXiBU1Vj7AzfQ+7f0KafrO/GGbt3sOdmYgttsh5BZUK08WTIQC
AfTHeo8b0Boiv8fc8PNCzao0U8OJWUbmOCMHNNqeZEkUG3K8qNrWWoILsdBU
xH6O1BTQ6vMg3rd7hq2qZxqwZ34Y3oYXFjpjMciMwhewvNYHzl+KGXcLkQmb
vVHwQk52NhQZUtv4lKpk3Zc0JGEmiGgWDDU9TN368OfxmTkeZMg/s6UykZFA
kbsgpY1kuhvCnYziq9b6aVVqHH74ZyqIEcg6LfdaEzY4JQZiL0t3x7FHNgXo
3wIDjT3DWDxQyOTHudKfY0mAClF6s5hu7k7XwjrWHF6B9dsBkIVLqSnp9JSi
UyhB30KwXsN0l0AZ/A1qwXVpvqG1zXz9T3j/zQ9biI3vsJMdWQpFPJNR8kG5
kKAVNwWYQ4Nic8f3CvM/1urvGb6f/VsHobDspsrFphRY7Rhfj7D0q3SGWWY9
mw1o+Vh2BvV5TsO+evO6fh8bOpNlhZbwRGNQfK2w0srKlpSnwgAmT7bnS60r
xwXMJEuIvjk/9Vu1JIPdp1RJZhZo2UG52oQQJItd2E8u5tduxL8Ws9UX0JQ2
bA1zR2xzNrmvhuSW+FWTQAprsSi1zETdDFHkqC96qOY+EQCBUgVD/n7+KVnO
x+ya2GZiSXiYyg54KNPmLqyPGItWRjHyoA+zUE0bPxOS7u6NckXmQFIt+Tub
fM2jBSRbXJNvnB372f42bGyocTmb1zAvKLEswxs+qugu0SPvbC3zgbYqf5Nk
lEwjIwqj32dnaF/LbIz7LK9p/DHJ01EiBgwfUtQK08EEK6rPqzhyX7RsUbCH
Zxm9aIGI7gp1YyKYCpgyMW6aD+l9fDGfpi7wTW+c/JebQ9eUr+S9NTOK2zrW
pzjVDFZLLuPRnPixFVu0eO2k0TT7MJUpPeRTPsJPtE5HB5jtRZHtjd2pJ9W/
ITtGgoVJqDbYjcQsvN+1WFJC/anuT60Q2+MIe8oEXb6iDXoOB4DtHGQ7hry9
rqEtWf6q+917bHx2hYpTlgO9l7srESAjZF2snOErIj3+OjZbHiqRTMVruwmN
Vnb8b1K+lisi6+Nuwjw3YTxGSf1I69JFKGv8pJRBGs3k3Laeg0v4vRX2EL0u
wtzXyRO9LgxEfYijFxNLqAegc0l5iVPliW2PkPmHaen32DtjUdjPoMm139CI
H6TPkg7Wkn6jUNX6wUWMw2ZYsUw4yw8p4I7DHYpcoTVwTQ9eSVdlP6b5swNe
HozJG7gqGf83ZDGDE5R8+Jq/DPYhKH/9niKZIDk+hxnFqs+sXZqdBoeq6Fev
37QZt0Nolra4mGf3EWH8lpIyLIh/6TkbTz1aUWAlf0DYj1PP8PTzAnJiIplI
IAggyRQWqvGdEgsX39KiVhLf69zx0V+J03WTtE/YJRWY/TU94wbLH+uHXt4e
4c8Ona2WWYKx402LItWCCtj51wOxDilTmrvULMdqz65PiXhImMLHEDzY60ho
soL9Dof7Re6b3OkmZmBt25Qj17Q8vj37xi6bcSALhv+cAdo0iTJUnBna6jHI
sbrKcp2pLIlgPBZYmv+u9Nt80gQH6iSTJQgYjOx0R0TAN/rYR/GPyFrv/u1L
YORNyPGpPwR+OXvLhTQ7Bn+g+lcB+P09xnu8NW+ndAZHshfDDY9gKAcdO+6f
geBA5xLFvAC29W1aSkDxo88VkERhryVJKg71rjUbrO3uROjh+MNtUHFlTWDW
xoaIotCzJMNqzcY6y5QNnTtzmwiddZC8/oFyLkglhisDxKfj7onuO4oxAiwC
Tt3dhheTaCnbfUuuBjpYa6qY+8F583yPAePJq/AoNhpzyEyIWCOxuuPMtaSd
A7ZcuKn78G63dGGWY2JRGCpBWz44CSn5YWfrfuYCRA92c9i6H2E5GfqObfqy
IcS3wOxK+eIalUl/kanuoaCWT3O0l4R/L9tD5H2DeIq2W2OfihNL8KDCXtqZ
4iZp/7VzPOD01Xu9cwyA1drP7wiufXPgz2gH6+KufjQKCnlHX3ApneroqNuK
gKwD2QbdRqudffTJbmQVox2a+H9kUqsyivZpE1+M9gwpKylwP5p2nl3d3aky
3SGB4Kj23UwfC35V+ZGKiYzPmnGWDT1KrQUWUluR6M73c+5rnUoWJU1vt5gQ
ahz4DB4cK83oq5cndpj5oIJSEMR8b6kJ9+YTrcas2sgmtM6Xo+kgUsExUHvn
pJopGKSjcunklnFlW7NMbiRbleUmbcLynTYrD0AnT9Qu9i8G1/umPbrz6Gae
8M0x1zm/hq64mjS+hwin3WzGGifM6nOQU5UvdqtmgO8jeUz2VJR1rJnJn6UR
GajXSdegqmBTFblI22JxGlEwcuR/9SbHfuMN6dKXdcN/nrakFhty++R2zu1B
2MpNUIND8e6dIczqt4SOYUtyVR/0JBLRjWnuYZ6Rc5tR2Lnd620zNh0Ie8DQ
s6AIY0XwH7Drs6EpoQgnsA7NSV25XaEyGXkjlfHEeqEUazZllIeumE/zPV3D
ZG9HvoDvm9Z+DKHOm1gnWINanBr24SMBCwfeNXGVyrn6hT3hiElIRnAxvGMa
Y/hDcUzQdlpaZNKuyWgJ4m34skxZIuvpNfnr5ViYJs7z0ONzRfZ9QEOO3L9o
hN59U0eJD160bn0oASB3okUKgJ+jtN4pqUBSBfV/04NaV4hv1FQjcs2dSrqg
ogsY4sVibbecAEhqZtlH/XaJYhJ71iN8ihhvsoRf6am5fb1JM/tED7VuegjH
nSDgEfyO1cGC4X59uMXv7ofp8SQfU+KTBE1l2RCF4asD3RHslNi/uFEddxWh
MPdPRuqlWcmIOVyjSvj6vtsFYByJkTDeM522H41HZxZ+CO8XJ1giDckU/FuF
IpXPnffQ5ky6M2QluJ1cB3HNYLBc5Wa1PgNOYZM0OT6aDt0vVDt/Fo76Mg6p
EhfMbtes3igW1iW21qLybuclAVKYawX5+ZvGl5Nip2w4JE0VXpmsDqIQKlUl
4t324p9MQkBwIFENcQbka3ZSPCiEigrZpNGV4qWijLhnS6jya1ADBHoU2oHL
ADa9gj1dpciPiksm1eHGQef6ESgcquFLQiiH/gi4mHqBZae9/uOcs5m6EN0R
MzE71zqV1zN1Y6AXWkyAcLKviyDKM3aryE6JSaI6EoRljCG8Xt6IYIq1hk75
+xreHt61Q8QZ1s3g7+EtVZVKes5tTqyIuJ8I2V/Ly1JJdvI+hR6K+e79oqeI
HW+sAz8m8elOERkhnX8BVXOKOVHtyL1Xj40SkBuHCO5jsxKqFT6nabWjC23c
3OfFTLulKUn11g+HaqvtSLsJah1VSAuYy3MtCHMh9WGMx/fyoR+vPrdErbDx
ElEc8axvs2+xjnYfsru7exuAb4ePdNagPSxskOvhM7dukeDtvZtYcCR+aNWY
X0XK8WngDtA9rlJQmTxzyofvV7dR7FmSYSJrWFAbNQ75bbA52wPAlasWSvMR
3UanJiGm1C80E7yYnHlJuwltVO0QpX2cncIXCaYx8GDvGZCiGZbDULL5Njs5
1JLc2xOhnNwBhVdT+RABP5bJJa88r/2y4ffgRyUOuMbEywBjg7ALZqzL4Ghq
8lFDVbSImyavIwsJzfW+aCJ1JJGj84ZA52BU+ZE0ovRHxfYYA5d5BEL4n0F4
+sTMkP4bsm4SLZNRIDEmXf9B0Wr77JR2yLXBPBcQnUGijcKea8gvuGQoaM+i
n23kqhZx4atdSqv7IBKnYC9g/2804EMf05wfx/3XpReUEYHuCafTPLKDem4M
DB4zylqLiipOVEf2SzfWk751WpGJEioCde30DDMsX61YwSVTdVmAl31w9CuZ
cYaKoc0myfzpVS/jmX/Ha6zVEvuI6f1KoKU2D6qJ3XIagaXL0lXke13UbUZ7
7xPtegXhobRDvpM0JDfrbMt4X0dMnH/gamdz+3wLPOz22HZa82p0s2rDkIHP
teANZEBDcWQ+bNZ61ehlvO4J+XcYeXlmqdTxcLg1u1grgkZtx9mZaSdMalsW
b/zMLgwgzdxWHbNN33NJkhpQpMq1XT4+i7u5X2YsmTcfaXQh/RTz39/cfjq1
/WuWaTKF1VRp9SPe1YvhpNs1xpyFVqu0Plu0wXSaEX3H/+9JK7KfFir19TXR
g7as2o8vOO5qIeknnvqrD2ROq1wrjtizohhTZoeo9RtueFEXR33Z3kRR/Fa6
J3GLPOLlb1stXsdSNfxqq/uHYKxYAYfosh+n6A/nJDnwVSMmL6tTleT0M6bO
EsRl92GMoilnSnNXovw7Hrmi3VAtiiHX9vPyK/XAfmc1LnjFWrz1wuV13jie
SNb/BMYq4WgbMTS3TOLhlfhh/X6so3CQ/bqn+ZTgYwCiwywRLDGWm9K3LGpp
Ho7K6WKyXY/P3SomGo/0r8IbR7VdGVE0D7O0u/yEiegkby0mHXuwD1V0hV5g
V2iCKlAhxqBJs5Ld8uWQ+qeOKsqfgaBUtIKTvtD9rOZBrN+W0j9TCrrb7Kcm
RAdNDIHwP/eU72aANAHp0SRDxc6OoT0vosz7otUwVQvVJcYrU7LaQ/WjmG3x
8votE5a9qzDmUNkYz8ofH8OlwjxMX3rSrCIjdnUOFLkgo6gMgZTd5oEmxF02
48A6fiH8lpBK9fXmizd/JQXW5O7FQdFTk47AgEgqPC0jfQb7T2TeCc8ivWr3
v2h5ffbAHWwvVF1mrcdCFlcFvrSiuIsCIb8DMmb6nE54nufcpBDIZ5LiLr4Z
5vdNfCCQ6uAfnH1fZ+6xWTUtFm7qFzXYmczSU4+6Sozfiuyv1iLDZZ03saSF
JWnx0xwGKuKTNm0j0wwf5pCqMxhKZOspyDNSCX6kLm45E4bJCq/wpZazXoBC
d60aGGjxFO/KHlgXNV2UtCjPKJSz+9JfX9pDl037q5mmbLjiIZ/tIUT1COJS
pmIl4V69mwMJ72/k4tqeJYdeWYzhTStbgJP2Vrk4sqCadfwsrip/japRgJyt
kKFwbc7IQ9tApAUX8MJOzO7/fPdYIFDpJ2JskkDYDDzGCPZTOZoR0kQVXozL
BsdXKQDlPxx7Bm20dmMcB8u0l32tGu003VGLR610RkODz/sSE/gf/rLFgwYW
hkbRbBY6mfzyKoENSV0VEJe1pxCJz7VMq2OtyCrH2wEsOXWcAxacDem7J/Og
8cL8EYsCxYVRFUltP/ixuRiPuf0ArIxyZkfgUOrYnbCaEF/7TNHo72OIuMfD
x7+OhTp/+CddsGvKqgQLrC77HERiqYvmxmkio1DiOg+Po8NHk3yZd+Ey78Lv
+lU/sBHgIV7USAzK6oR8ocM1rxlhwDZQbupjphsjfy6ZfwfNU+c0v9u/D08N
Uo/LqiFszF8BLDcFdVToIkGzT+9Yuk/NCZmnl6te0KlqhjOps1bNdNGi39mD
3pWd8kc2qQKk4bOk6xFvWMXUuE07K2IXXxB524SNlBE57CnvTnn5ye3x9Th3
ZBwuGAAgFswSVFJvcS1peQkb3gCNDjpf3MRvTrLIcATcmJG2fBoTwe+G8USy
0+MqvVyRjqM8NGCaTbYitNK/oDfsGY1TNLx6pszF05RTOEXezA3Bi+sSU6ND
sUtF5IF6tgo5vOMde/1t+MdPWw0FYN2pd3d0x2ao0OXtSfEKH+Mv6Gm6oCYM
F4GGHMwyE8/IMGO+aCUHzc4jUNwbqhZPgFzcIelLZ9ggfdwMS8bBUQkkSXyN
ie4ZzxoLm6LGMAy7lRZ1k42pdrQZAAQMzj+DaeSY02S2lcxDeuqi1/bNQ6QX
ghNRv2987ayS5+LVROS7+yCoAc1twS7wY6LsHuzD1CrgHbhGQyCAryFNB4+a
BZKqCYYbox9B3aBGYLRtv+uC67fnGOfbZkptL0CS8/YyawFgOi3C3BVrSW3k
WBrUPeZi3UEuhkNE2MJukxK2WyGz8K/tPwUDr9z7PoWZuvVUyh+dZpakIRBO
1Nn+MfITp33X0sfrMEq66CBiT3xg1zgx5wlGFsAtFJV9JDchpo/l6jQ5PNfj
MNrLKrHKYE7/nNi7q/Lz07xWerl2HU/h5xLSUMAWkFoD9CcjDxkqhuHIFTUQ
efY0Xgwl3M6XzCh7MJQqM5hTY83dj1BF9zR2Num3yAO/BOaa3JQze7nYQqhq
Qy1y4VW9Bucr7e5S8k1sYCF3Gb5IKJ+kw7suqaGeqbVCU8PN3M0wEVSN2tA4
ALWgRtU/gWecubcQ0jm+RvKRSAFOQ8fkj8tv7tl+hUTYfrvpmyz5KKvXfQcM
hLt2kUOR2tNPZlmd1i+OAmVmbvshHxzix7MpONzGV8qiMBog4wohj0prNkAD
h71sjkOSLKyEBHA50k/sf59oUzOn3qCxKBCCaIjV7t1jxCsDocY6AH/Rux3C
1symgGc4aCR1Lxw4qK+EAlZiIuAzDKwLyQzTXokUUBRyHNAoHcjDRcu0Itm9
U7J+qzt27cAFFUJpV5XwMqpT4iPJgrGqeHf/lRMx9zDxOg/RpTrpHUynDJv5
7ygng0z8/wv501ltWZucp9TgBzt9gA7rfCv3VIGH4vWfD256SRF+trTAqFYM
4iGFRG0uN1aSA/rniFJ5CLjTfO+1wjfM6Yg+pBUUs1gXZF0ZblcZ2oVGu8YS
gOfQ9RhF6k+koNrolwRaBUzAKJfePVR2x1c1uErAcqVf/uhaIDmMiBM12r8I
hoUk+VjmC6+gA2iqTDJ0K2PY/491sA+xYyYg9o5SpIKMCOx44RWO2keC3wbs
xjYcL/vKzW2BAbgLdUza3JWoVWrNA5YqaLKMRQpU79TIp9xpDHU7j3ph9Jv7
NocOP1/Jas3xiBWbh5yjNSZY6UFDIK3jKube8jb11/6/b9VDYQSWPltuIVSR
hMc1/QNkY0EiFAGnyv7C/8OSm6K8DbtfsCSB/xHwYS30tOMwMMs0FWRRyaWq
9AkcAwRd9gCFK3IdNswFLlFk4lS14+L3xjRKWjQRkAMPX0YlFyCdrjk3raZX
6IrMOSpEi4Qg89320byrjjXL9odz+DNyoC5pfCrftUdV7I9qOTefbXbGyUhO
RKp8hrp/c5AEgCjqkszovFS3puoNYAyS0imMfQPry7ORWOeJYCIc+kCeSnjg
xv/QLAx9OSu7dxXLeF7jq/LBMzqLxIe3gMnKWSjiMrHDFPan01980bWbW8P9
YgAraLsAsaEWkROzkRGG4Te9HMwJw2+c0wFW0FyUotlqvHSuW5Hs/g8+toZ2
GgwF5k+IzLE73TSJ+hOjb0zDUxKl9bIWJekjiwqk2N/JfmoDOcazdOH2OCZA
aYEw5nZQkhE8jRT4l/WzdqYjHlakHq80Wzm3i14zDe4vMdNYU0JMVaPvYcGF
tcS+UtnAxUspx2aqMkYFl4u7y1W97zWbnw3AgZ8bFviA43kMWB43QnL1QNLr
F1hrWrYkZgaiaIZNYs+WlfH4j3hHm9p6/pI3WQA2ktZW7UnMidjAkvJk54qL
X0zDVuD1IlShcIqD4MBCmLQZPl4azVyMYVL+lBwyaMQdcEfo3CC1S6xxYmmy
yYU25tqokOVZaSOYE2K1aXcsfIVgKmyFBoufzUbm+k9DkDMkvVsS0sOMRsiM
FgcjT6PxJhDlXJeZhjvYWmy89X0xPNHui8qpiz5/ykDOMvVbiCxKiIxHnPXz
dK8uqeUAvUfPXVMURFitI784kBRPPrTMMucPY9SKNjNgPdRHbXA3Hfxjdeq2
DzMnNvTxyO99xt7NYJ2eIuklZqsLj2s/EcYp5QXFKRfNZ5op3slgJDFcLWJh
tuViGgy2UvaqNwSmHhIMSyhF/dqD1t+g4BuoMZ/3dPs/iwS9b5MxgZgW6adx
UrwUNxt07NBUrheb7vvJXqz9FiCebrl0BIQSkzQQGKRsTeaE3UO7Un8z0mGd
3kHBoUbyI2lQB2Whm73bjUyTJ7oLcDNkRjhV0kCJ8dxbfvqsXgZDM40hUTAx
+0bm0gBAlNd09cBQKgB2DhA4BUC5aF6ecQTQeTMDJDfhWDAPlbVJ7+55kQUF
A8NxBJWIUoIF4zztcuPvKRfuXuQM+eD6hruRMtMcDpFnXMnUBAWpDa/+PPhA
EBpjVM50tKapvodvKGcpJyzFu3/27qKKvUMuRCc71wJAImrBJnx58eZCTjP6
/UDf4zBxwOy+KoocbXKk8m6JRjr8+tCae2HvYhycQIP03LQ7VnTlW+1VzOPU
Q4whkhbuJxDMofRwxwmPom2oJIoxdWSdPbMOe0K9XnpWnkwsOLnm71qXExs3
nXzpkxlWMkcRNrWJwQ0DJQVZPL3kqD4sO0m1lOLDQIyh5bEguVtn8ZWMOUdY
YzWHit4g0o0h91TeDYgfP3b1b/PBi2ZmowOh1HSWqfeyXQHDQ0RHn+uF1GSc
AxIqcl2jdVLCHIt5YMzWP+Q8wbVp5hEw8f9bbksgEEm3FfUz/Gn2E60CLvPl
/uTW+LQhv6Jt9ZphZ8SXF7cpqf/E+6HVN54mtQd9pnvZ1tYqdPacbJXlNswk
SEX1Ii54PG+T9bJnKWwtuL24FBtECx3ER+4AxIN99h2KW21Gu2Q/+Mh6f9Io
/5ztD0b3HtbwicY4sy5nTTQcg5TrkknsB54/BoONcKUGq4FVvQqfhp5jbZcn
MIdUwuphjSv2Zif/H4OGrbEl5gRpBSKwCoocEV4tklBVQ28ib44zvYG2/fqo
edOa6v8u73CWebDqlTldUBbrNC9yjldU6pEwdskCjy9AgkD98Hfu55hyZXk1
vkbGQwyKXbIXJzXeC/6TQGH3adtXbU/YkLnjd3H3l4N5njp7ATZgXYeg7cz9
bji1tCxiCtkSKcuiex1MOpkEK+EVZJ3g+nWMXT3HmjoNwgt4Tonzz/Hy41UP
lhW23XE6QLhXzvwHbLWE0CSlBOPQF2xDhfauvTw2QIh3FXfchSi5GY/pOMMS
3jghQKmQfLMUXTKm1tAGkr/B2WrNTdgwvyz/RWus+xzVY8/2HLf47BEeU/2t
8fDzj/BYdJWgm/sBquehC9eXUqE/eg+I6EmM80sqfsQE2s113xQmsbj2Td++
FAd0Mmm/H0Gnlqe3oS145HzJGQ526hjhQ++v9ckNXXXXJW0vsOUguifvLnhd
7AEDALkRgZLvrLoHdpqMXClzlXeGAjVFokAM3B1Z50Fn+jLt/mcntExY2f7R
16JZ8VKGIMeUJvlJcfIUHyYas0h80N3pzwlmu+oCkMAx4KxsssoGidzs1k/8
F2Yjr5HiGtifrvd8QmyYOLjxviGjsApQULFxduAi79bQPuvS4KUu4bOs6I66
6HnheWaA9qwJFi4N2lhda4/ervFf9Pdp3RypGSbJ6ZyMHfEDb5Q3OPXz3yfq
2fL1L3AeoLAbRm6V16qg7nGdkqv7637PklquieaAyqu5O8WwazuVyvFI/yI3
FjGxxzJV4IS/CWsb9UWIl1saKU8imC/BzA1f06Kr4h2pqEZY4DtB6AGGme8Y
EuszNOo+UwUpYeWrjfYNb6iJWXjDaEhUlGKfkqaUpXufPP5t8G3cvKE7KHX7
/APbk66ATK/BPwpm50CCyEZGcrE/LWGLbHcgi/q2TlNIRa6SOXO5VkL6hI2k
tchnNBuuw7VcQunD0UgAZ++sdID/koUOVis3dXCBs0919XITkw4G4ex27Iou
maR3tFwo/ZXqiSdaAihLFSAobPRKdeL/qxxqCZ04Qw7mQjAu2hrtEQ1X5lyA
pATM5OdrGVbEmRbtNOcp8V2RTmItsR/E9nJk0xkxCO1YiqaGXHkmbkXeFrqw
wbRgk9IT+WW9BNVNzD9gv9VBT/WA1Nbmoz+TrA6grbe6wtAeBV+nVwP65B0A
I7hU2d0/3H7xlOrN3TupuvBwODXb+PEMUpVQayjLKk8PG33V9zcV6rFJ8kNu
xy3gu2WKz1XmSdxUwbj5c/89VEYfB7VEOH8OEg04CTTqqJ3Cd70fbdXA0rFH
j3yDUne+bGCoQYJy5JABIZEZKDPpV45Voe69BBIeAg2ad2Vw74DDsvSiqWFS
1OicxwsFDR0B7m3TACz814zWY1r7mC1L29tlQVLbbOZ3TuvCZTdpWbz0gEcC
kTQsleuklAhhPVrM2HDgpDj8IaIevFj1i7TVM1ANgJMEtd247Q5xzPUBpnwW
ZxXnVftTl9knuwzVM8zQgxflmiAVvgIV7DiBWVeM4DUOUHTzhtm/+BcYG+uS
f4HsbmLDqaDJRtVRO0VZCHhiciHA3YJCVc+1zswP4m5AHUkXR4sxNrieXFgC
Drv0fAJOobtxV3dM1v5NiQNvm2bLhE5TCy7CwVQrozqvzrQioYGUPnTnvZfq
L74OJmoiyqES5dDf29apPfEA1XAPkOKgOui/tEn0qrR0QJW0PI7ZLmgg2g66
ImlGz9UgFJqjm0OPAgIMwNlkELcUdt4vKi68hg6Bc3y/6hkWsu65osLfTWb6
95dBmSReGSaNymIujPuOEzE9sREmqzx7VB9BS2q9LwjAnrzuIBwZcRJPGYWN
gn9QducAfRV8+8a+zPqRIPO7+rZ/pbfF2DpyCK6LEO3PBeYQ5380zqC+fpEB
OmDUwePqAz4CIoXV+CJJhqYEOk9DzeElQ0o0fIwJB7pshhUeg7YPYDHakzZU
CA882ZyZNH32E59+11V+HAO6faM0lar7lqFYq/4vee1AtYGJL0jMsoc2CZo/
Jb++D47t1aJF3Uxw36JWKcb7kAcHoKOszjYH+oc181uCB4GdFlX4YeQTTFJv
6qVHN8rRJivogrcmb/3Uwt7+ufTISYGeQ+oyt5zewT3bdG+BMxCzKDTEqu/7
m9GtKuK7MG9fUbYvX1pt1Fx4xAsib+e1taRdj/SK6r5R7dz+jSwD0N8LT8ES
4LXZJXzRkoe9t3z4RlbT9QxY9BsN063deFf6A1XkPIuR8SkBtHPkWKwAccuB
2TlylveXPD6YzsX6HYj4KOhTvJoEoMNTkXAR1alNvh4bGjx9/ig3IFeGDNT8
Mer99xedGuPn45lwcKVsPQ59JSbiq6XxnqwIwgibAB7y6XheAG6q5CwmrEuM
dZ6NatCHnrs14mIjUG+W7dv4eLqQu2gf7E5w1eZRmswoMcb6xFNSxGfi8cG1
1ecAo1XllNJIGxmp+hBjiFZoybiVI4z6vAO4CC/2Or7g85eq7GvCk0fxwRyS
8x+j4wg8Mdp7dsC3veiFtvK9eFGtW2j3g8Z/wFNpH+p1qWXTe+OaMv2HheZU
Goe25oVImaInKJRVcjMZiWMjn3O4QR9OU22Gq9HjrzL8kJ2whcoF2VOkW7rZ
vJTfLHbGrrDPj7EnxWXDlP20fVO/JVYGRnnBXsMGpaKmfBrInjZbZV3N92kn
8J4WXjH1ZOTngP/IaqiqcTje0SvN1USiRxvWaNcJKR3ydsIBCoc0HMDj37Zt
x/sOMXexW0O21EPFexpw1Hq6MRtPSy+GjbYmgUf4YaeFGfUUL/lzmoZVNr3R
FqtQZxGRc2LPJUe3Tn8YQ2C03J74WRhzO+KiIjc30JLH3uqdTORDvMNZN1KA
dvMlGoAx+3DN6qt01pMsoJztJmXh5nlIXcrw9SMcgXOugYB27OwhVFddKjN2
44V3TxJbE5SDFhO7zr8NOoyiP/by4zXO6rct8AR5y/W0DxxnQ19yu09SHTQH
hzuLAxuRNzFa3E6o1qnBowXay6Fm93N7PkiA0oLqi2Vfdds62+RZxD53Ax4G
HhQrGM3L6VpumuWt36Og3GAsTfBdbyFZFxMsAQssmHFIz4EdxOOhQF4E6ulJ
Yx5VZtyyi+YehYSZaqUmMVn+eDJH9lIQ1pVcojfDnO8K8XG/qbMK7cTNtjXq
CemuJ1pbrxQrNTEY8wTWqTYwZU0kWHiZv6i5DLCymeYrnRkT3AmWsQhq0FJK
dGka8wEciIHNGELpBFNzeT1PpnEtlDGKTsUqlwU1bolVXrOw+ODFM/Vd6fqa
pEdNVSeViKrhKFLY93KjDEXWqtwaFzQdcnd++713YcDIAPnW6ffXamjTQUkQ
aG0u8cm02KB231QbZah32G19fyW4u+xnSp8De1ofoPa87GV4LohUOMRR/8zk
hu/iz0qAFnFUnoqHBij4Gml8LFAuwgsfQyB2lBtUVfQQx3hW6QjW1TVqcA+t
suq5uidb+bpshSQ2GOmIEbOQLSi5iUJFvKKeoo6e+fvf0IX5TKTKTmOfHaSJ
xZCxDCKb9AAIAYSV0z291g8mY7aHcB5GOkdnpD+H3yJjolFtaAXJmIPB9OJd
WZi9TmlPfVw4vnrI9DzJnzZKOJSQRb261w9CLM0CL9/Q/3972NUztxE58kkB
lGQh8RNDS4MS2OND/MgA6Dr/ImxYtTzmjUVtZoParHeH4WBbBaW1jx/Yg0A+
tl+P+LOTx9jDQq2qQDeaYxmksSMh1fHiPpsYdIc7hq13ek5v7wjbmst/gLL3
7i36MIr5klXnMH2XD5z12p92eplTP7vUz9fwg4cwsRgWotv7YYkhxKCh5uRr
qH6M15XrqtMjyYYgtnoatV3Cdc3diXl6Dfqw4rS1YMvlX2lh7vcsYxF4xsar
z2fD+zBSQJl9dosh8DkhAB+NOpDpypgf3m2pEZX8Vb9CX1yRLASv3BVthcRT
XrM0t55FIz/r0xCix3tU+OqU7oecNhtkfcxNrry0JIOH8gaoQR3CPPF8PdO1
WHDeiZXmb+pPypJF6sr4Yo7UPPjzfV9O59iNbfD2IIT7HUK3QNH41PaJrR4E
VmoRHl6BuhweVJLNMZ1LSeoktFnLEmk33Ejoxka1oKyI718ISngKyeLljPKx
3bg0EogBNaRZh0VS2OYSnk5rZz1f7YGI9IRp3W45XKoeYATq3OKJFkOodwko
QEFG1IIkleCaMRZOQPLcFz4OXf4/32rdIECp4WQTKx4uUyLMAfdGX2jgxJHN
r8h3XwuDfSjE6CPy80xvyvjPxHMQfblhBbk9Qh//FS30NFcS73BfyJBrzF5p
JbGS7w8hG2IaDho1iT5GoJhBAZFEXpBJbCKr4/zflFzfvQaiZW3hZNAEtaI/
d9GYQe7Dbs5LKJ2EvIoi99/ys8qGmInzdKfku1rPkc9Yh2beLT2854UvaLn+
zusfEfzLyIctYZYSzslYDhG8ZqcmaYFaJ0M7URbi+96QXiNctkziF4e3L19W
rz0dh2ncwV6aIt40cR4s1hMUeKfQ86TO6TifevZXJeVuIxAqYYDpHRJ00qs+
I/liKKUf+u0ScZ0fJi5OZPd8RnHFIGbIie9wJ1B7x0NwVGwEBgub6OXtL2V/
87IQ8KiUG1zqDWl85Yps2zwMv6fOoa9NgVmaB76gc6jliVFIhhLkJG/xg7Q2
YXQdiuJnp+Dlf+ZAxqoI4ZV7uMCXTNP1Y5Eco5UFXFy72w/+cD+jWTt8fk0b
uOjio1Fj7C6zNwX/AtvIsh0IOIKGEKOFZxvxMo8SENAai0ABE+eBjrPWpqs8
km4jzJRodcpIdIiAZ/TFHmn6QrWjkIMwYaDAiz0Gr5CUhfk4/zX1bmUljZfG
fB40j+femDX1BMtsjJvBUotLdpNhYqzyGWt6ogNMOPN5VhKYBIiD122mMuXo
54BJZOKmS4UEtytnFdhd2oJ55SmXTCiUdC5/S/+wCOK/s0jyMvO6qvVrrJzi
/+iwWk+/Sw3OguavM82padJYKzx1a2mA2dMz2/j2nc/b6U4wH8r5rWryPBUz
2UhBJmL0HTm+VJR6GWuGbb8+PSAcd+HFZiOo/jAsJC2k9ia0dYBG2tpe9cNL
yycVce52SM1cRLSh9b5ehbqp7sJOZ07XF/sNIyZX8hL84OJXGIqKyptDh9FR
+Rt2D13gJNnWc5diL56yImMWHkgL9vDUyANNgP0Lob8P7A+R7LhcOpXhscet
730CUveKsgwr+OkMp9ZPETdox25Ekqvo+6VvsYn2Qfkvtiqu9fMz3bs7Si5U
4qsJvEQ5sOu+1gYGTpGamuiXq8T9mituDeBzUByIowpaOMIBGDBzSmfTMC/0
4rtOzQf0WZzI4iG3il69Yk24y6tEo+YwjiKh1ILUxPCvPRO8AV8P4swtb+MM
jS5/NMRVPg+dQyt8ZK+aVKquxumopOqRJuJuDbql9eDdfi7haPEiWTWLmcDk
AcvdcWhwkkXJWl46LonGHPYMKulv+wT7AE3jahnz17xUSaW4OIMsSfo0zWlZ
WELCcG+6Gnu24B7R0XL/G0PvQnnqTpDlnhW4wpQsP6ECFLQiuOXXtyUNnicv
SL+5mPMQdQVIjc8Xfu1N8o2wI8QfDFv0vRhex8Bo8IxGDLJ58N9XVD6k9iyD
j1dNGwIBCOpJ9Jzaqd3UaCcNHJbpI/3ZMzwVBi8GPzO0asbKQ0V1W91dWbnO
L1x1mKg6vckBzCKfhWy/Ufu0Bdj3QHMg9vsAGb5l0xo4cV0yokhLyTJzl9RW
jHkv79/IiG/zVjS7fHXTwrbn2mcTTXUncOV2vZt/Z4fHn9Fq7s/aZ1ihB3Ri
ujUIVLZA8MJQHlF1CHE/2YWdgyU8V7wKJW1mZ7xCCdo5QXEbdkZewqz77/yc
JIjN3VviRz39RP0bmkVJD8TmCbGGvEt/Glf0aWV7B2PPg4YaPlm+0sn3BIS9
X/1XZ1uJt0QTizTk4EyL1y8MrYs/z8d5eU2MVVMgawONpeliPCkQntR6Wor9
xBj7AytX3/rDsRBPM6cSOVAGRtWXgpB4Xwv9Dy8Vd9ktCnlscyiX2NPM6vIT
0frWJDWgGxbaBMIFusdRL/hDubCgQTxu11c31hCvxG9VycEFvxaNthY+Hhbz
25qS6lSD9REO5VnzOyu4Tqr3thoDs82L95l1FMAaJ+q5ByuoenhU4LvJoIia
rvRl6juk4ZiYlwagMAJpIlIz+o00I7lEDJhJ26jTOTuIC707d+N7b8eIMMch
ITovQJ5KEePeYOVMpaOqe+EfjoZWpIvlNfmokcBS73yx+daGLv+5mif2Ol/U
N0Bp8yMxhlH+JMRw55JhiTKiCElqQfoNLQrvzSjIIJLxED1RZhjGdnIXgd1h
hhICubqQmbJ87VREnAyQpKakRDrvpwcwPhMXXsWbvM7ajDD2rxa9CbVM+r6C
CN9Nb8ahv4ZSIBHi0Rp445GEOVpJ+kM/fTze/SXg6dZJctsZ6S4RDKbe6pzj
fGRAO8i4ffdFEbCtJZ1IRR88qJjwaaEAzSmsFt9jfJTyOAtgPuxf/TQx8DvV
kYZby3DMxCmAI8hI+fxSK5wWNnWH9bp/rjIvggKvnog1g7KktHHsP9lIi4ZK
3qUXCsdMHSI+jGauWK3/kO8ehyXcIHQTLUertEaBTm5VxJm24CeJDekJnUoj
fzY//jUxBtk3kMlGyBQlaff5wWJk6CKfb3mXaqYTavQv0Rct/iWsbQF4m7uF
ByXd5nyBw8QNOQqfhSd4jbCkUBHsm/WwlXM0VkF6nuyBx0ITAeBWZXjPFWvx
eFL7xsy/NEYHihtUtmDi69Fk7MXy+UjVD+a82kTbGx7It9+SFS7M0Lj17vUT
36R/mt3Y1apGWjAPivFZodGPk4kUdv2oRNUjtAVyfBwD7/Z95c9hKOmWzXJz
WH24oznyrvslItny3gbnWyg5nbBf+1WCNMLD2HbmN6Jkt+IlXtowO68kBFx/
7t1DFzWhtKCZGKR7DRnkm6hZmYWjMYVPLrsVD3QSDJvedtxyCoSzV2MxFLp+
d3y5m/aN+WZZ7Cdyb3wDFlHuYT0s/v+lzD3BhZDjt70ZjIpJhDkiOCf9IMCX
kyHFmj6fnJIpTMKt1VQNjRWN3YyQrFPH68Hyc8pZ2LldIA4KMfGsSBXrcYKc
f09iU1DzUmDga0fS8AM2w97wul8V67p0MIHqF09CJQOsZterFOd9RbeHIpxG
vZWj257MI2abAgr5Q1MCBY13HrTNvj58pfJK1xOpuzmoD1Nxgsf3HNHhtql4
paXskMDhrtopIl0aBmGTWmQVjX5EDRoSd6NCZcbAMxDeI15sO0+H+aL929IM
Wtc7AND2r5qpPJsjOW4tuVsq9voVUUCdLSiVCE7ILy7CXcbjugwpxtWfUMFb
mwnFON2PQ+G1PIFigz3tVWUYgbrQZCm1C7CgMJhQbSq3DzIVfdSMhchSJczK
SvFFBNlV9cND3M4cZFsELW8cZy5DR4c6RdWShXRsbn6GTkeY3l1o55pz4zrQ
7w0hiSqB+jp6F6Hmi4Gu5b/ABxkZ/Q68dzp+7rR5/2yhB9IoIzPlXWifuv4j
5pE8vUUZbrb5I20BEJptupdarKvzkiWLbzyFLXaFC9AOSAXitD/kbzGxB67u
Gku1aHvl/lFyQ0SBN5csXWlsTZXAQ3zQnCMCtkGgUZfrBC1K8awHcaeAQMX+
FSr/uI08WPayohUOnpOMCV7Q6WB4PqIrDEFcQTO/wBKRo6O0v+UOHvgHhYd/
MbPWEP9JmY9hbVD9IFv5FRj590eO3U/m+diBTLPvf8WQhQqUWATa0Yf3/2I9
1vcTfjffwXQMaZpNSklIAyn4CoqflU2xAU1K3drLAYNYQYJj3nY7DnCaXrQH
hhlGuCnum0wRW8CwKJ9vk5c/6wtML7+wa36AKl9c8sj294YvasrhEph5RtY8
LtALRFumjG259TmqB9tYRyVmWFT4BebepYPGT7MQoPJiLW0WetnE6fmqgKk0
4FmXHZDH5CHdEEMwzhjspAqYdCCSR/rKofveau5GtTw3iFgjIMP+3rOez5yU
P4+cdSIvZVcIv1VMlUnobdt1RB/a1vVQrnjRxRldeUlfKU28N/v8bWN5n9eU
6dJ2/cTRlEjlkDLYZaKi1nBgioWMKIEhoLrOUOqqGgIhrpMUjPY+7DEBhheO
OnAXKIxoPO4FaeLhA6zk4zUDR3KsXywLhmzMg0TMO8LGWVDlknsCeWd/4iGp
S/47NQ30LJcB9iA6BLyPhsQ+21w7AomUXvtwNjYHjKu2YhMMKBgZBa4rLJ7v
RvhWnmWaSXMO2n7520OkmjFA3JQd0clomttcEHtaOy0zu0vPM2LwLqm47rH1
8uREViHDK+rYcEWgy+r3dKAjCDDW8ZqKGfElhd/QMscSxsQgNOFl695Zi78P
ifLcHJSdHlcZNknviANM0cAwyT1xfyUNtiuRi8NcRKkHb7y9Dj18p+Ccx5z5
iPYTSm8MF4e5aEwX2f2jiwAri/uoY3joc96G1hMZyMHRGZ1a3XDfCVJEe977
9zUbQ2DPIt35yUltCAr2/Kx+uxpuOBNm14wmomcne36XgCFhVSlrvjAf4GvL
aVq27CZVim7Z9X4F6QX2xsj64sqq13ZhtMKylB7vCHmMmN/Xj/OQriT6jOGH
H809EO7KGHFOIXjtEEIJD0w2tujk/hg5B3tTULkz6t+sIpSmclHCM7Nxs874
FUADzazMs0HsefOVfzbrN556ut6Y9KeWjJBpxyY8dcznP5Owtk210SVyJiTX
e3q3C2aaEaMCQXZwcO3JJQl9wAOiUXkU0+IhA4resj3iMyfdvaSNtUzCmFTu
qEa3v8Rqe5RVflm+bKZn9Wc6YfPvBbQ3RGV1072Icq1+6rpQFjvLlbdv1NO8
RXG7VGpSwfg38VkA36vzmJ0klkaOepORsiwEQ9KJRpseuxWrbSRDxy8239jO
EL54GOStRUOiUJKCJpifkYq03l+UL08pnzaYz9e9W3kwHdnTz+FtwZ9Ib2qU
mofAnCeR5u194EOmUfHh7QiRMurbbn+l6qguNL4boEDVQBfgk0tMdGSJA3cp
E3Pda1QxVl7XHxW1uVni2EbTOLWKcVwmGwTfWNuC/+TEiiL/6Z641s9ejNyH
pXIw8RHC9sVVZxyeVaSm3dU1jSYctHcRkVl904MZHnSF3h1u4miQ4zmkHLDB
wy6HmoXe7pHt1nJ99TrHBisA7VNtntSMFGBQLsjxi8jZJVD4TXMt8F83AvKF
uaH909CMJbIJEB7eCEqp1wrUvm5zAoFhQk/SB6crGHOYGxUzIqqDs7PItA1n
F9lzGVJGLO61vTwFi8KgvXm6XNqfppaQJBNv1APmEZXBR+R/lLK+46vZPx7w
zilf6Qr9VVFGdtL3vqVkwg9x0+kLqPmtdwwnoZuP55rCIp3CSI8H2AWYUJAZ
GfHWgaURjdb4iImYhhJIOnmuh5oFZ5N+A8vrwPzGFS7/KQctYYn9O4DSuBhj
7t6CBp0UwOHB4VaCXWsiaqhqXg8Hv7McsnI0xcn15V1AH2av0r83M9roZCMZ
oUuACGF83Amdb49h0DhIoLRhvoDjlYSmTO1PPdk5dQBNb/saMnifNO0ZtqyA
Loa8qrhEl2jTnrKG7B6M4v1aexIy1NmiZrRuNGsvsJDlYBclZjgCJEyUndDQ
zT5qtTaGP1U9IWF/VLm+0EalJ/z7dFLnIgLIzi6QT8Fjv0p+TtqUlp4aPAGu
BQTWIe9yZnVIP2skGJADzDCYUu3X6pKZxv2AeDrYfQI1835cwtREyJienTPM
vgUGLhRfyQVoM0gnHcAH1zYi8vdey8Hf6/m+MJXT7YiQM5CGNeyIiqYOyUYd
4U/97H2cKOkhMBaOdfQTfE1ZjbJdEtQO9QpPWNEWMxRY5eyKiPuL7aH7EjNP
we9Dl4qrDYhAzodChmnoUsKvXK+2tGZViMz1rC9ccvLn43J68SjwGwZljEZC
2dFwtHVOGQAuvrSXq9f+T9Ay57VbUmH+0rM0voLwX5jGJ1/01fv2W6CyjeT+
dXPBv90mtQex56qtoZyutc+QlHZ1itzbEWkq9YjuASkjjvJoJTuEzxdVcwmG
FamZ1/v2yskY7TqSagF9PMTnZO5/kNflRKQsIUz9OIYr+LsoIn8b7hQm7Scp
7B3u8slmxKnr6wJTqvGEXlEWE0/6rH0CtUu5m/CpetluAB8D5iF74GuVTPCB
qYNyaBFnz2Ghk0LsGAkAVGMBkM1jnjzvZX7pXRABcEnrdJaJ8p7YnqYTRdry
FuI0rt5Javx5AoQUL3tIvWEHB5gLqmpudGrvTXatDrjNz1TtGr2zEDqY/DgG
2MD9zAdfEh1dSsL20cf6qPhdNfybhbn5FDSvYFtCidzGdzH3PX5esB/hjuUN
iJsYwt9ayqYAIzJBHp18W571y+IRSnX5n16fJE5Zw5hBVP3k3C9Wl2tHJ09W
u/nV6irLAkJ1IBbJhAi5iQKMGxqWKhstfVshvvdKRz+//gN3sTkPoXQF+Qkg
JX7zYuoIIvrjlAkbVo4qFQDfJvvi+/8P59h9+QPX/EBBYkwQQYehRh+7Nrit
yzPQC7TDZ4hPFU4Dr11y4zzOTwWnGPTd6AcaYiBk4puwTzBtoCShdAwnc2o/
E/MDW5s8SBeYu1uVDSIRvZbnZWl7KlB0DeVtqUA8T6slYX2dcrUoskPbcFaW
6Uu/VXpZgbzQH2XSmZ8CCqxfccKcQ0TltQcvDA2dPnvBstqx0krb4lEjiQ7Z
zx7MAfW71T0wMt5Zx/XCYOzjkL2EcUUs/LF+UepGKlKe879fvN0seAWW2Tio
nqidLs4oJh+eiCYylIvZ3tmbVhmTzw0Yl30RX/1FU7W7LZvDyR1Rgdxfn8J/
ZKKe89c2lLd3ZR2A4PjbsglZiYWPsCT4IGSFvDEZ0/bFwZb3g+Ys/BEV8Wnl
2+056PKw4xdL/GuVYozyKmiNy+d6UidpViF7MYkYQXZb49bUSwwAH9BjjxUC
P7OW56YShP1wocFc8N7niWJzC300apjAkjlHFRE5FWjp41TStfoHey9Sz0Vr
+48nDIsz41Y0K5aCSEDBNEkGRmKj+97E+gQ2t4LfWqFHsTlFK6RyvpJFxsTJ
J9uZ5ePs9ynfhLanSyECMHoMbtAejmJWAggOSWFaHPEu0zB/AyuuPd8NIgnh
TQrd7sAVbQm00Pk3AdZQyZQjrnQfOJFC9SCP1cVmetkLTfXrbAFoDLPqPo+b
Wafk0UdhEDLfPlkH77Cxe/CmspZPH0rMEhhhWafzfSm7lpD9rT/fy3ZHGpcj
WVsooa/iOcjsy/e4aWP2EB+NZFRAzn8hq48YUVZBPwiEe7z14hnms2II+U8R
eLKLjm/xE/oaltIx2xu6TgtVVKj/iD1ecwV+rnqzs6wxLW9iHMJU1kEzvC6G
ySYNU74+S7N2xdCoVligo13y27dcJ94firfc8RJ8wYEsRNAodnZse+gmTSH4
rNyLOvubcc8eGyVMpmiGeGwInV+vaj8emFLuoUIHZC39VKf2lOQLTLgUIHZx
6opNjvOjUmxF5HuAk+1PsRzC5h+TuNdBBxYjDo8iwIWGUJBMvnkGEqRwP5i4
3GddNE9lVnxB6vW6InmOCcdhyBNe2xW4W4vdtHeHswrqzlFfsyiN5H1kSey5
3KVW1ZXNiVOpmq9Fs4zoBjd7dPPlpasWWsi9op3YFsxtGZtXukoIN1Y7E5q2
K/QhmboaR5NClHRYuNR4yaBp7bDoSYbAgpXjbuKb5hBoQOEsoXABn990XfwP
Od9NuWNLWhENTeGPFBIK2/mHtE2VLI+Xpxcx02Btyq+JQxGA7XJ55Dxk6N8A
WFxOLkDpUa94H5F/1lixe+eqGsg2Nrzw16s4uGXIcs2LSAGr2Ls41oQQwNsL
C40GmgW3o1WdkE1tXuwJYnCTSVMH2YSDIgJ56qbm2S8vNUJUb6EzrCjKiVhY
UoDkLI46CM25OFwJqijOrYIPgdLAd0szrEQNrVHm1CpKdd6JBLqDX4OpTsuo
iEOaaMTRfmajd8lGtVdkBCAO5stlCQZ6OAJ5Ywx9X7jMPpN93QWULl8zy+E1
3Uy2bEVwNBa2KY4/++GikMU2VX/2JUfigsndQV2Fw96JW2pMpvjrd1jbChj+
8prCL7rp2eH7Vurstek/n7gQ2CmjBGQBcE1NMXi2TKXHGoyeq419TIvkROV+
puUinPEklOYU6cFblCNSsU7kvKy8bAsq6U1LjFV72xVahMBFg9zOwaS9082A
AXF9MjaY1pLmYVAHoGu88EgFRFN22YK/V2A8lI4L9TBJW/lOsI/EcicFYAoV
Yb0ScAjb3/8aFdeNhpfGIyXx2eNo62KQ2/mWAD9yKonRs+Fg8Q8El3hD7CyL
T1/Plae0KCohrQZnPRhoBikzb2wbRzdF+QqBHhfa/2/nQpzXgTK7lAjORINn
BlRpkhJNh7kmNrY6PD8i5MYjfAz7T04gb9piWQFyNI6vtu6C6jI3YxpOV42M
S3YsqiKuJxhGxp9eiOlFFPmzpWY8N2I9N+VEGmD5V2xbWiAtd8wf0pNJTMSg
nKmiYzevUC4ObmUwUjvAfMn4XyXCzhdhGG4Niy9CIFkLPdLtPU5HmoCbaZj4
+KPhERczoDZABdCHoBI13LMrMF+/0O3qpWA981YXjWT+HpjIuuIrdHVo8z7D
fxx06bBr5FakkVIjKCBNk8WFkeUq2jxfmIjGnm4UrTr5XEU2mQw7I74nAKfy
E25pLUgH7Ge+cYUEaVpua/zeSMM5iexRGUKmArUi23x5Hf34TDB8UYHmTfm7
zAuVRr25k/hAZbq9W9k2hZgRP6DW9toLIdZUehs3iRRGaR+zI4cn2fZp+Kl8
zubm3CBItZcVIr4dl+FIKOzLvjOfn5ScvKWzw4Pk7jiUM7Ke/PKxUfHT7/yq
1K8KXu7Q4P6jKR6LWb1gunG5TSbioR/htDQo4PsHScjgcPKeACA1bL9q4AQk
Zw605/SaRh10xHk+HPBRzZzfAkeOSIjit1UEZrbs0sniTiK1ZdVocxXbJqc0
78buAhBIl/X7n2YN58TBw7j2+PoNpuW3NJGh7skT/pPIPJjXAGIMYa7IhNbK
cmJ49CwA6y0+f7gq4NsIEQuRwMd1pQLu8ieV7gdpZSVre6Krl5kVkGbArrfx
7kVfyNSfUi4+Lmwo2Rrm42pOfUmsDypDaAImGfuBB0yulXC2CjRwLvZiyRFX
pQV5rvrF6Re6ZmOvZUR3gZUtbsqeSuiT3d+LalSaK58tFzffJPARgXY5zpNg
M2VYCTi8GziQKXQzp1JE+DZQsk6yh1wlUqbKJcCd8dZZ4C1cjHrqNRm3y4Ba
PDqw2gQY39NU1koyotAJGlN58TPqRNw3tTN7/2mlVtKATmo2uLp+ahy0OTqc
nBQbsRf3CNmoK4DkJGrWJhakkuFU0lwjdAC1uJsCd0Z5EErRPuxkRhinrWhI
2UTLISlKfuwqGWweglKRrkMXTAA7LeyDJfuxibi8aY9jOjFOuDa9CI17vgRc
a3Zp3pfMGLA9hl44AaE+vclzdMcdqHplM6CcX1DSnkzWoTWtrGz7/UtKLBC4
yW35YEgrMrUBtx5NHgNRe2JDgNmj62I/QaAxAxonYncalsQsKPpyjRktvTwH
9LzG7ibqmwm1KK2hgpu+tmVxP3TvoFMhU/N1igkAs9vRD4dpPBD0vqGWJ66l
YUA14X6+VuLfh44+DUj8waWjaPfYblRvaF76hPugs/s6IRP8d0nPO4Xp1tsL
LGQgyNkpNrGpWrQ0WB0YPOWvee0lP4JcONKv1fNApZYpdMolO8rFawSu7ojx
ng4pCmTQkf6BjhMThHWSPYJVIBkC+eQKDSLCv2kbBSWmFvRFLfHGq2I3Zgcz
ud+Us68OigLlfsYRXcYUM/zjSYeZQ2UPXYe8GR4rbVogJw25G1NnTL+v4j1v
NpUsicbsAom67Jaiuq17G3jXlxOlM9mslSFrbS8sjBXx0P8DLy7iuUFChpuv
pfaewsUCXvzQ6Y+7BoLDbijx+h0aCxjj8eA7TjbO124mu7UVV5tdQr1ia74I
I+J18jI4qRlS1/jixXqdZL080KcWJujLtdonTfc0M5iOWmrifd2D8K9Wte8q
GBENAUaU8Ir6vquEcixBCkPcuWzNtAU2IJc8epiNZx+Yyi4rAd9LsDqo7jm1
85NS5qjYlTh0K1nPgfC6SpkNuUH82eok/ogbh0izQnvCMCpYc8wKnFul2XJN
rf8vBolYqGX3NydLArYCJ2YZAXkv2squ+t5pmabk4KjMubgOzsc7JSttzofP
3MbEKNFR6DnDaJFSZalAqNHkp/RhkHPTusUlMlnpMtSfYi+qbyizzDgOZwfv
LSkahvzu7Fsq/2d8AX6RYi7dRS1oKLtEfU16EndW7bcQVqlfV+H4fCoPlLGh
DSe+07Dw5rWLY3AoPl60GWJk6UMG8eTbjHSLIrHsfjjw+8iZ8z0GLHjV2ll3
w6XzUcVoY9HMPfonRf0fVs1hwYijsayp2Cql10GC3dwSCuOQhvtaOmN4aZ/J
4HWh0bjQ6gno0NI0FrkCvoclW2zc7uEa3Gi1+CXfARtV2WUu7/RS5wy05dI/
HkiRq1CqhuMr8oCuRf9axFw86meKmTV47bHv+60bHZAIMUlAzu/erF7LYFzW
T6XlmQumDrAIhm5Kj3R4fGQkJVtwz7I+ZkkErb/E/4tUmUJ7sNttosirM6fn
VdHN6X1GiJMTwDqJxVyHykDRheZFuq5ZnmSr5RgdrUz/Nnd+Oh4kGweEn48z
r0wU8lEZMYtA/ZbjivYj9KUGItVHSRTFWvVKOk73XmxB9DXwxp/SI2V+SPNe
PV4cFDTa0FvJDxDg0p5GnA6H7lFZXNmzTmY9XBWMNdtOPVJFp+aCz5tFBXvL
wcWF5TVHtS7rSo30aveef/U/hHP7WGYCQYUfhL+dw36NHxGs9oLShmsB2Wvg
s/GjHGT/M3RdFD0GX4LcDZSyZk6u0RSQDCU6pkyveLXpdF/CQed+8O9HTpkQ
/W75hs0XxdYQzTXsfldeB/B/1TJUoF3pY73S5TspsoH7nwbIsXnby9Xr/zEb
EzA9EB3kHtfrO3NMQC1lLpe8I9uJRKiyMSyKdlC681e55uJ5kIiJdJ/g2EkK
rWJshr0eXTZtD7hZQb3ZeZC8gl27n2tjx2dh4SZmQ+pKMTIZXb+GrqJLNKtU
P75Q6ZlShor8hOalhb2nSr1WcLBXtp4Vm5CiJJNOnrCzJh/zkknARyM0nh67
QSGkRK/UdKRZz96d+M96lM1r+5aMgl8MqyuLZwnmssbVSa2i76/cdOC5JkVj
YR5yKWXu9HJk4bQW5s3KTZIOACifbW4lDRm8P3h/ib0Uq3trqJ7QT5LIJwUj
RH8aoGnAmFblH0WdimXYeznWyarcA6/EV4VwqqlVLEyOY+C0af4h05Et12ZR
GAzVPQM8rz9BQfvd2Tkvyb0J+/u2GvJfrDjRcQnaLvNrpIqhEY00SMiAl4Md
CihFlKqg/iFfkG5ar60Q58fARuUpcPkE1FhskMQ5ZaSf9STe1ZvyK/B6clWN
IOrIGe8NTgJtonU7HveAXWjShZ9njSb0gIDi1x5Rf73KibsZUzH6qvopbnG6
qAmDRPc9gJzktje0Jd5MXitD7Qi8s/by+mYf7+Xy8yEQUBgroBlENdkcwZ5B
senL58RZ6c+8ohup/UQQjvJykLbNa+PIML/k/bABRergo4cIMXqLiskleONe
PAiUWvcLlyqzaTHFWkcQD1uTOP6O+gvZShxzIutPOXX3Z1iulJH0Hc01bytK
zdnZxAFe1uemav6gMfcbeuqFRnpbcMkOuZBezjCuq9D58ni8hQLhF5cxw29U
tsEmBb/wwRfk/lDy20uexi1S6rmBV05okt0WCgbv0BiPp053TtfQbC97Tnjl
OIHvUvcBAtYE6qK7JMGouBPnT7yg8xlQNaRvbTEOEzOanm3IZx9UmORAniMz
F4b3xAi5f2jSSW2g3Oi5zYR6mG5Xs+6KzCJU1afwWG1FICCEW6Ypk3++aFi8
nfF3p3O4lexi2dN3o3TGx1/1Q5K4MK52bbdfQw1WgUlV44+dh4Y81qkV0hkR
7IdG8IJrtwEKj49cemEENljZZWvZd6HErC0vmKT+jTymqcvfAJwhd4dN1jiL
eyxaANWd6lJzDcugw6+A4krLlongvi90LHumcMPMULcM9Nfv8DVmGgwpOS0H
K0jmOI6Dy6fOyYqODfSiwq/T7L5qo5UBAIcngTEvAmJDcA2lU+8uC6X6V0q9
zIrawT/oUxqsMhM59WEOUVBUmGqqSoZYsr+nd57s7qTvtpyZ3WNV0Fr36vCq
ZNDAvlBT4J1n5VgogDHJ/XaIdW7GnHqeUmA/5BqKGeCmKaGzVm5Vdo5S4iPr
aj0gHTqkzXRq/HUbjxrZsya78WyKtprxtbYsnf2KJQtqLHed7vpJUSu14sHL
j7BtBfoPdDgMnT57pZoGlxnkX11jPPKyZG/8Y5scmre6v1ki2Mm18woH6lJH
rBbAUg09aUoKmyc3wsQy7KNGWCnIkhBP7GXG28xWeNlrvLlyr704vun4M3OY
CXECeaCVcPcDerz6JQQ2SZmsVH0DI1bTAfHJr06yXp/0lGlCZsSqudqKCXFv
RwyiNPJCYY8vvjj4BeomSrXkm24FukdK8LyxcRlWKcLdejkNlZDklevScEji
felXMZgptfEjxtZ4ICAE3zXIys7s8fI9HvKdF6tu3UpDpMP0Tm29jiQaqZVj
bekVjcgXnR4GTU1RmHCjTHsQqSBGanc8btozSrAxzoIk7C0jRK37iunkRRAt
xamXxHPIHi6K3kW82tS8daUbHIsamruukx5tvoaHnhWS4RDZvSej8G5I7kwH
fHOHld76MwzF2unWqlcJHmOGUVSZg7lCjTEx37M+XkPV2hN0Roko5b0PkOJq
Ns5f44ncB2sK3DihSNK+2N9jnl5j5Mn7LTTegLZVJfB++v94Hld+suhl7XEq
s6Am7uqM3PdwKuKGvCZbpg75kLghbGZL+5NvpHGiXYAo/vLjQ9kFNrI4avky
KNJqvmMCvLp41ahPJKabVq05Kqn9K63w7FLPdDQfVYEJmxNVjYFXD12l8LdO
EliUVwl1Su++mbEh2fxrUCRTd5YC9kAifTY+HKB2Yp8VuLBa4sYNFF9xH2t4
2vomz4nLUukx5Vm3lgvXCcYBpmKCsU6RRcDLlnMpFsNplPFAPtb1fr6Ogzys
H6geVvmgQ7ZA1hCL0bKztihljy+DAl+bXC8s2X9qtPx2hmaAIz0g7RKyXjyf
OUfPGzYNK1muMoje19MJaknYzQhszG+UCDHrfgEtC0sednMhkcOmfadoDobb
mOE3+dKV6lSrS0JoCvDrDVEpPCKZVUiR1BB01d0wTTdnl620CLGMTQTF96KC
/YlVOxMXXij7FNEKXHsisF8iogc0/D9LAcimpovIrKVuWdFeTetWgs04pOzx
OgCcTVnQUHmv/uRPb6AdnayQlJnq5+qzhCbsi3EB60vTlfNxKitnWwK5QJyB
VlaQIeFrAUP3wIQAYTteoAb+7wIkMgLrXzLzQ1AiSwy3UeWPLtlgpu88I4yz
6/KngSDyvzkZQwA5U0A2dsaXeI+cly9VIPq0liEXl44HkSPtgllcqd0aU3nC
ZAZkva4YCyj/r+EVtZErBxnoKu1tNvX2TWXI3W1WWDukukKeuldyf3O8ILTH
05xDAVIS/wqk+8XuJ8x0mn2Me/lKvnM50WHIoXjO7Xm3XQEoE1+uthrDIgbN
yaIUT4BZD4LVvRAuOTzst/+F615OPCScPU2Tj0Knqv+/hb2NjtbbVIPLGWGs
p7GR88pdIwOQ9f6sp6o6hw4wdHgyl669+qKF2IRhYZShy6PyPaU8cEWTM39f
4rbEsYZ/9yo/23Cb66aBcbo2EwmZnk3cwWREDKek35/OAZCm1kAZv+fm+dcv
za0EiR/tPSxP3MNVNSM9+SzRTzc4Op9r95nlpWvOSPZdrTxPV1wXdB3Z4asf
SJzPbv7YLacLOIh1gFK4HyrC7TbEBGkCatQm9k2BjtpqzlYkawCkMyj7hcIq
S5e6wVAgx//7haoPJRoy7ewBYGi52DeQbtXKcAwE0LdGA4HJvG97FuQDOJPo
XNcd/wfbpDHdZhkxv4Bn7Q38T067PU0TBoViEhDM0gB1409XaaiBE6Ihy2IO
mBTLIhzX8j76I9/YaXqzeqcfNQiGl3uammwMiu5kGY0GGUnUj8Cjz/QBl+Ci
bMUHeDdvlXOH0u6njRgS0aEY90Ojx+2YPXws2/n/qVLnqPXRo7Se19NDNCdi
7wx00ZIarH5WScEyUoVe4HdOmxHwFjjFwUXJqv//zQYu7AMlx3yGccA2foun
nELIJJSHyGJW5AFoSziEPKjyHERJeu/TaAbNkpluqIJB/S1gZqo4R/lFLkku
K6isb1dZG2oIz8bJUtZFjoPYXxtTqyKMCYTfEm963fNXwjy9+zgQSiDI5E4m
ptYGYXP4bPYV6+fy+F/RRmyjHQsvt6C2nrm8UyVEUxYTbvyvAJO+yqepGH5n
Pihl/Q4J7QHos0qlTlWiVBOhJE/+W8zZz/69maB5j3c7kHRn9PMR1H//q2qD
CvH/a447y5Fp3Yw2G3E8IECYqND+iweoq7BX0nCckfAqh+0EImpADTVT65/h
ZG4uwO2LwWe+6QWu7R6UkT6cJUnZL4W+0t1IdDql/wMDIEtDRLGy21aWnVcd
6Vp0t4s2OXNKnIHfIfLNzb7nFim6k83FkYFa61jO2bM0W/+i4mbo9jl3ujrN
H5JbACxhXYHZcj9ohDml5Kcg33sfKi8wEF8u3SCOO2NDA912Ce7mQSWUFaAv
ih8BwyWNiZOb9AQRT110n2MIK2l2I0OcjKlfHKxQYt0RluYdOEuReSrEAUt1
85WW+tCzxC1iQ3l6zT82oYeyg3dM3fMCUIFr9Lj7/rxQBy5K9hF3gN6ltJAY
jqAc24V8PdcVZEWoneqQeySRh9PfioQMAnolsjwKTvaAaAkUHhTc/9kCesR3
X7NyiTe+wW528ZW7IXIlpyo3HMizLNMpt3LWh3wHAN9r97F4Ugoubz2c7L2h
KW9uQsnNk+wZv+RTApXUsa6jYYS/xeJidiLs17bgvoIdI6MN1f/ypA386kiz
xdZed3saJIFqXBCbvJM39eceeTESpu460BlG5qFfbAjwzyg9dbV1Nqe29Bbn
iVAfzpz3LkXYYf11GQM4LlJBsG/flJ+HJonnxmfOdRMyF4w2SuNUG6SlYW8K
V9nQ15nxPygLpodaaSiM86wNSp2E1HqOB6590nXQDsdWkid0Kybg9W+Pu3CZ
i4Z0rSXXVUvipmiEFhamq4XmKv/dKN+wEnzQ2kkiDU4wx8yzAP8XD3NnFNC5
igk79XI1pJuStsCqZ6K8veqHyJMWJ9xdT2COLA+EMYsw9zbUSMVSQ2L4bfMm
m8Z40eqENP8k5stAblPBbb+rJqAF3MDSy8SHpYy3EC8lAb0tKQi/MXO0zY+0
xd6FrodcS3Q8+9gTOkbqdNvszlfz+jSrbgAafrxaLlO/IiSsa31l6Lljhv5S
PzJwxCOMS90IWWI8vZiukFJpjmOuy9kZP8g4SHutPBzfkPId0vg+l1nKt/fr
ITlbVH9c8WQD0/Ssd+Dk4h0AfA5ChHtCXQWnLtFcSqKW3/o5122v5o8x4CoA
vqQbOZXV9FiKx9PWZjVC1iCwsU9cItLeRXxMZQvwsa+KTTLzJWdGo5eqxnRI
+a2q1RnHG2NGCcLq6vBEBQvrY0quh/OtFDtXhxUWY7Z/RwxzXLgNBztDXvr+
GfuQdXVBpZsIA8mx8a2uQmH6OgiK/898fXDgJ6ay7WeYusQdRAWqo4cx+XLw
gUfvTwkPHsHUqJg83E1F1wfIS2/foluLUgbClBzhES5/r4av7SRqXnDzpBdU
FGAyvjKWpR3MoZwm5JsVAlahIGyufM0G5UH/w6tGXbb1bAmQKLwxbJ5wL9sr
R5SGzX5Qe/poKNSNLcwZeNYWA8G3qh3D6VLCAgfGfmkequg/ANpGHqiGrQSM
p5JqywBTXXZ1uSU3v2rIv7mT379mQGW/Wb8QeWVKpuia7qQQAOqANj9ipmlu
RVAoL9jEe7JXfLpstLOX/HZO/q1S02SLAx1PjdBOQWR1/B9bzykQ/puitZEq
0nTj9P+krT70AdA5glL0vibD/Q18HIYGvMW42NMNV2kjrboU3nNTCdsoyCNt
aSJ1cVEZWH7O+cv4WznIzIbO8hbUaFz6B/w/xX1KUF4TVg5zfJPvAsmFok1o
7VMuJIRqTsSJHYcK5nZ0evIz7fNJ5T5gHYV0gXA89SRsz6tAyh5sKFXLkKgv
n7QTTgsfaauov5xlMZiydgbwnBu9rVwtSbkN9ni3MDP/h0j0XZNDMkrqfAjB
ZX/6fol9dDjUqX4EqSzMfoRMG6qxBnsAseio5ry0+t++fqpqksz2edlNfeCT
rCylYiugdZZoUOV/XQ8DYMHgc8oaw1LtWw0JGWT2iIJGl0UFsxyXk/z2NBgv
gRGpMz9/VtEWnRSausuFSdPH90QUQx48nsDuCLOdj+GH91GXmynANTFKAqKZ
tB9ehJMhv8JLxkKefbDDc5LdYcrJZ8rrUfjCFT83Bjaz7xzBzFSnKi54aYfU
BOZ3e8zvkxG7RZ3gXdimu5FJ3+EwJ3UbCoMSQTQWe9iUp6tQP8yG8uIBdwpb
X0DdjD09V8q+pn8wWBRhiihDI8Jb2XBFbGFFkq8qvlXf0e2E/Wm25MvOWCA7
LeUu8X5WwhyFPkMO7Elhms7ofMb/6za0ooDHDlVyAJDUPtBAJINPmc3TQqjh
33hpllDHKAh6xS8ObFNywW+wGwvqosLWQR5uqW02TvYqkkCzP1DJfqawS41K
2avUFJytUDX4vxahcZlZnUupL1eu5zih/XgZLlGjcEoLRuqj/KaOfQxBoazc
tYVvs77/WYKKWD6YNEQE1LmQIbyxNDvtMULZX5BmpjtG2kKvvDguzJTH5G4T
3BhWdO2QeXydKdP3n6LBMRVqE0n+U5HmVEiHKC2YzLrZ0LKv85tRbd3zFT8K
ybyFsKjdoLO/MXrtlSXFF0oLKXJIZNzfyL3H6IVG/cswJg/APCUs0UNdD0ms
kD34Tk7KWz65kAVWtJIfukb34KFBue5PCIzlPYPV/tHScUEJnPhy8IL2gbte
465nfUujTBYvW2UtE9PvXISgZN3DHe92MOsvuQSk2KznWsjUsZ7Fe3iTSEuZ
kJy+5slg4aZDJnAKJ9HapExmmAuimecEFpaeuS+pgMwc/PAxKzXdcOpt2nrK
74/iHZDadQoQKPaW64flJ+JnG3mst+cjM9FSVTbZhsN+R4wkhbEVy197Q/+5
8VMlB9vI6QTfo9IjrdfJuWi7Rwb1GAnWgHRebPMTfvhYe5jk6rkzEBRtxbC2
e9dgJYN1vkZmUHIZP2lC1LKFcZCcquiBnKRsO9Eim1TMySdEF7iYTsEqiYLr
D+Wk4dOftVWwQVpB6RTDkk/JKJ6vqlp53dRyCm2SKPmV4uwn0ifWtVZIpiOp
Ee2qWx0z+jRMeY75uTb3XP2Y/OKUqLKyMWM5eh+P+98ME9dNJSSaIUaHdb0K
0ap41/R8KN3Rxlu6YOJmGB3LFNInBcRBnzCdOTfVr6anT6SecImxvMmzvMgk
0SFYagSOK7DltL/qiO09+jrGdTKxRPrKgpf06bIzsOvF/ZafZFnW9Qk6URp0
f1RBe1A1QRkkDttFYWZfzClvG4lxcjuglNbw4Acj/T4/DUFDmY40XACMfWy2
T5c905LsvInd0l7Q1nfOFvqs36B8D8b7W9JO2BPp4HdM4cq/H3ECkkuq+PsP
UvLFrEjuy8Dzlyb5ppbHnClkClWCrjRKoxvG4+da4+RgTmj57nWgid2phAxk
mdqQMU6ZELdIgBX3k8Tse9j8us0NqTunObbmEdX4ulv0wNlZOBkldccD1L+Y
g0MY+cfsvGWhLGzXmMAc0W3/HhCOPUfxPX7aONWrq7R0Qm403GPdNIxuZ6Ce
EwIfz0s3ruxr0sHU21hii/lhvug81rNGtjc4tedsB82sAlTdAFp6UeIuHmby
FdCPQYiuXFYP3xAfdq27AczsQUVZOP+DYRqFwuKJH8l0TVGVBG8eEvFwD4gD
oWOw4Uyc3bgTvA8h3bYp0CaotF1qKHrut7tD9yxPPcJJFQf1n24R+AmIqte3
0+0AqJdh2IuG840C62dXvGScS4gLpQa8Vf0uN3s3GBWYRd3Nj/0qR6eDykeu
y1auvkGl1NlbwtcRhdK3ypyP9asGn176oH7CE73YXyGSdg1qc4g02uAc8OCZ
10llL1zb9A41geJEkF5On8Buten9jReZgtS/oHNHrf3F8PyqLK1PAE0nKSJ5
4Zx/IEO8zKyiVhJ6KNKUyRjptmHH+YzX3E5APQHHtrObuhAd0VXIsl6mUfrc
4VhCyhW/MRcyCdlY5cNPpAGDNKAv4mwv+qBSJqoOz35ZxXmkzxtXloLd1RTt
f+Fu+0I9Q7+YiD9E4RJqXbjxBWNueOD5dKq3vroryYogMpHbbeXrhu8UwJPx
UrsoXzi8dIte0ekPElIMGHSFGI8mzoGyy4CxCAotIeWecH+y+taxZASxnP3P
SnL/ZvIHWWCtFj4isAoMxqhADJJgLKg53UyI0ug6q/UmRnp7iVHv74Dk+II1
PqXa86fenyPeC6H3RhRy0oi2x1x/IuRRDPL3AobEuxI8XRO01xgpFmllN7Vl
8oZsrBbrEAA4pnrwbnNUI+GG3ALfozGJUUQd8HTrYsm4Az+qWw0KgyY4/Ixt
wvaoRx9D73Vop2/06Vh26fn+6zShN/jexhgldZOZAVtjzl182edQgmtXTuMq
OkEIPhLPHzqsrAX1+EcDleuJqf0TgM6Giz1PHhd/abensDkUoYn30b6P83tK
+g9TXrDTbkDibH+moJYM/Kj+yRz7nnEXhS8zFLRBreLKkd4X6EFq/NicHG4P
MmQmBvGqcfbpFt1Q6LLOU+v15i2YOeDynm7iNhSv7TL0YUBXzZ7qXhw0w4mH
FlS/zaECDuhHxrO/EIz63dmsk6aNTXPj+7McecD24uJrZ8EMEjpRvTWK1Wwu
yp+SrKTZgLcpy7oco9f6AziyKm6BlfJoqD0AhQ5CZkfgezMOr/4sXtloONdA
gDYouX7T5MAAJVLFZ6+hLw+3kI3Te1J+O7DOtAr7Mi8x4BFCM09aebsgd+OL
fuhVFIKBKMwYhiugyFCZpu0cqrGC0P2Y3cOwrbW9EzDYEaZfuTp+ylWsZCHn
q1m2/SYxKTGVPP5wxQ7DLqk9kFIzHYZtNw9XrGbFhka5QYZlPjp4lJ2ECpIW
dJdRQUuDnyGugL3gjFaoJpOSwVj+RqsGdNh8R2dpgcqB8wAcZzeEwj1wq7U+
3A/0oX1mNHKDetp9IDgj9tBm5FeYrjhjz0thfY1rlUxMUJgNk+V24wU6KSBZ
rbXlduI7PDtrjcWujQ3deC26PcovKRC2cnEtSuQ5dKgiayJb0HkOmW12wY4g
cwyxQxz3wYEdH3rUpMFCXCAZpm3i/cx4G2FXCGtDg6P2hCy/ZGWnTCPcLezX
Exi6ED1XqzOwMiiE6K52wUkragacD2BarXEz9n+IyUKfdrliec8PHTD/Tp0j
2oPBO3ROVoNdp8C7jZYKf2cQ/vCc3FcuuDbUahLyGB0mL+o6S3WhGTYMKHNF
2FpRisRHO6LrIQ/ZBmU972DT7ld5etzJWHz1Ncj5d+C/FpcQ6oTbYbCQBYj6
SNm3piVWa72F218vV4GvlIWRilKy+lyAvJzqSVF+9huF/nprCz0Oqd8cDG2D
Xu7IglWE3R6WXQNXIOa/OUrgmCPo8NKJ4RaniBBMMq/nTHp2TMC8JbBrmCWX
b5GNrL/RXqwSJVMSNQ03WmKivceAIYS6XM24w/8TzOGMwvEumMqn7feiaTgw
JZ1P8v2GfXgq8c50sLE3o8Sy3jHqFQeyVUzytM24bpSqoQUECp17rNO1ckPS
ghhOUMu2DRmjrvHMadDyfeQ6pZQrb5dnJ5y6G8+kk4i/IvlBdkiCIGYzvld9
QHLhDLWi/PN4HES+lYAGAVB6gsItp1t8gM+EdjFeQL7Rm8bN2UNXnLAmegBV
DcV8ltj1M0XLZobLBncEJzw7cegFtNdE7fPoYS6B4YcUO3+eRRnPbyO7QnIo
Xh/5HipRM2FoKUxyMltjmiqNfQpxZ2gDXSFlt1UfzczwjaNfLDMMYbPO4BD0
VuPeo3A02aAxaPCtEOTOd/Jle5brdjMjQBLkaY8x57UXBYNTo0byVjepjFo2
svGD/F88EFip8wwG4HpiiKOjyz8fpmtpyGE390rMCdGquQEGOPXtrYH93MR/
ep0pCKuqhvsQzv3TB0KxMya61imbg6Q05abTZIj3w2LamZhsQiyKwAMgeUcb
7pjOBe4Lzveeni9MaeIBakvrblXRVuMOayzwGwZztq4Tt57oBUGp6iZNaPZX
5deEhKsqi2KTF1EtyPg/tbXeXzFBYMPwSLQpI/uA89Zl7UUqVeKtSldCy4tK
24l3LIg8QaSUT0p2Dmdcx7efLPNG9ivFSdAt8rdBEUAmG0kRMyNwyWsa6GuE
KuT3EdxCfvftGxzH2+w7TEMF3iExHmngoHP6OTGjdiq7Jwb/my3zbKtIlxAp
xjdaruhwV5gb9+4QbYdFziqUf7gJ4f4fvQNDRyqFnG3FFbTwZNmjaYs9cubd
C9o38QZSXRva1ribh24M7DHw3qB8r7LX5ulNbuM0Qv75Z6y1H5ELlducu3fL
DiFnHIGB96BhIEj34pPOcE4lnAuXB3O+3aL2/3dFyF3AWHA2WTOZc1PFJzwR
HsmxlR8yBbj6bTkb1FQFTfFaY1aNB2kJyBogePEcV2vLHmysBt8aAv4LeSEQ
cT7I5mlzU8YCBdo1DsVUqbaBYV8H1x9pCDFHCfE3RxdQO8NEbn0sazX8sf6N
e0RccRL6WZ6giFY9GkH9IKr/gRXTfr7GQlbn8pI1wLdsffer56sAJwigbstY
txC58MLQY882DHHcyM9z+OGUpK0PKFdTB1opdBj4/Sx6Px8aq69LD7sEGF4l
+2A4MMUj9AOlY4UW1CdBznsVMDXGuZfsu7MB5eOW0vOBQdoPddcW5JWEKZ93
RIgtSD+vS+mQ8rREtbuo17aMlcOxn41ASd5UrEdoZWiz1kVl74V2VRDk9SO0
fDi0AuuyrxwOx9dgxq0YMo5J0XnH3noi+QbfmaNIcrt1V0kEHCs5FEyZbznL
w8dAibdaX9UZCR0CbNkfLQVCnQTJISTllUZ+tzxdRwzSOOowNJR3ovqfN9AK
qeNVgsA87KraL5YR0yG8AbIARrMqvRhw2rPrzRbKB9sbv5wSRkBlx08DTQVn
VK+r+oFPNcgIYxapN55udnEt9nrtNDNqbcsRAOp6n2bcBiWMHRYkhIr6nlu+
/cW4sVzpzubJMbIjBt6txOFzcQnJJTYS5JtUGUf/Eqo8gEO+0TVwZWsf4L+1
InsaSNHuUTLT7svANUrde7oNIAAYam7a425EQLDU26mHPHyXLZ+EJ3G2U4eq
TqMDQFHRbC2uq6qp4qNVyjZfXjiATE3iVZ3yLTtpcDu260Oxj8wMGIKs+cbX
VJ1QTd5PPjEKoFTU5SNISseJJfOWg71zqoYen1CniYxgeQUVU0SHrVDyNPqW
NVxlzu71hb3iD7OMxiJHmhhMWdNnGh+wmakW/y0axVKxj9kqnOxsILLHGLQ/
96kFA1qbcmvenrpD60eix51FjNEzCDidUpbHP24o1/9uo7cU1/R5EDhqlaKk
OuCE/jCayx9WLlHGtX2ms9y/yOq/QEeV/7g2Ddvkt13WgDmR77B7on1jsYV2
iCD9pdQ3aMCxdxC5BifbnmpZeAngBs4GMW14EtqwM1tVBxhiwRb/kpc0N0xD
ezHcPJpv4jLpiykAEKlvYiLpgEtit/Dxg6z9kHpNjgQicruMnPKRwr4dOu4c
aI+2LTYbzhIGLEVEh4CzzBStELR64Zx75aIgxbrqlJLskC+YmLe3KYF71xWl
01FV6Djdkm4mbAJZc13sIXaohlTQWgc+hW2soHa3XoHKScOa4CP7wuX7Qumm
lFqIxaRSAtIYVkwmgx4VtBtlvVFmwWs6L1o3H8XFatQS3Yl5200It5Vaz3zO
GWQeP502xcFQXyrWpMbsfI1/2Kosm3HhzBP0QyvYEIxbx5kkNzM7qn2nw7Xk
5/2fPvPBRIYvKHq3HKGEh0XFgLJ5yLXGMFTTRZEfg7SJuIFjKenZgQPuBM2X
zL9BfJfV2DU+eHCBhnKKHQDz2fnedNQRTenbBcAisRIebkXPciTDtOzuCtIK
Yzdyeghrh/wJm4RX3XTM94Dbcy6PULPrkqz9Bcg+YjzNMA5w/xGslGnvJnxK
EZ2oKQmiAdcON6XgRND+CDHJmE5ds12oCHgyw5vHMJTcpCElrYTlhcytBIMC
zAYRPn2pTfwqGrAKQpJJyjC9Iamn9ljEN7ftToIsN+3dZecme6QoaXkZufSL
tOWH6dTMUjlkSrsq1LFKH10KbIGXnQ/Ov4Mx02k/VQkceEy7yQ9bEbJYQoDf
XqmtoraO6wQdJdyo+1Puq9Y9XiZu5SN0p6/9HJgYXycC7xAw8eqMOK82UK37
waJUPBYQZsHcydckdeOHrCJT3+DSYLB4DBVJZ8Pzc0SPHWGHwmhSSNJ5EsYy
EsdZM3ZYuFAADV77yEqRxpxSFVxuNxSWWClkLMu8FY2cAnbC954E0bOFZSDk
qOySwC5mwLFXyCnWlN0NMCp6t+Jx+dHljZq/EAVvmmG7y1hTs9W60qPESgbz
GOSJrnRzwXUhfueaR3HPhamJmIA1BQ83xGXWXZUhu+2qzrhas9edSeRnx2La
5SC4FKfSKPKOK8hYDCiAfzT+xllD/9jINvSrs9h4v8+DUHHpf1s65XxBWxi9
rWpQWUR+oTCtQtoR4ZBFK3iHd/Hwk0gZKjS9AxLsp93hWkcCUwc9CxXwFwfA
4jKl7J8OtFiNWVnwh7cdCFMci7+83xeu+MqiinZYY2ZFwjgRk2uuNJ21gHZ/
/XnWChNNbhljgORqlTHPsicZTvsKfFyIZfWdEPwhI5I2RR5bIs6U2b3+PYpg
pMApLfxdA2ToSXTCGkrLQX77ZQ9E8+kr3CmYK4Hjl6RwgUEMdYfNVRdOlaGV
sFXo/CmeSOsBDeAfcAuiHeAvM4K78gDtZmYG2VsFdbYQhM6wm/3LpIbYgTQn
eMqgEQRD6YFfEznuHEkvC8KDTvPlndcqkm411qzWdxn81drpJ28vbQSMxqWp
0rAOtrT2CWYMS5x/ltjncrZKPh8PlQxRmZbpfRWeQOFxzvSB5oGSDqX3UYDb
JFhYVgxXm1nSnX9WKv6CVF+gA8SD1UUix+l079Te512zAr4JXwemMpP5uL9G
TDQ3hM9O7xZkT7WnlSKhf3K/BQZese3Yq0/AiDH9dBa0Ge+sw9LaL37l+fuR
oeAEYBnmu/qQ5VYWiQel9JzTdcq/0VRLjRcUGlKLXy6uh8DycHM1kD2DqCqi
ZcyrEptYpFoszQIQukgFOaKqTRfwztawX41Q61C2JJ86CBRtO0NYerNaiu2M
/RFvZvLNy9xRldwmk3QI1sYsZnds/YnyNnXFhaImuKoEevNm+Shg1JoRfnvW
Ch8PHRTwKPMPImHbWHEAXQNvRdv+m4a+8hM4PBoCRMtP3uGopFN314MF2EBG
4uhkLW03KewMbDEx5UwjHQlCpD0wm5fXqcNdbFQCu/YlowbFADk6WNY7Os3U
gWicjOOsIp5syhtm63SdMQ4CWTh/56H4w0zDtNhzx/G6F+u7xS8acjUOaW7W
nGQGxg5VfDY3uOYG0bXwbTVNoOA6Qrfcu6acmhfxPNbBj7WxT68j9q1Vlc2Q
DqiDNS7kZZr+xcPkDmXtZGa7BSdj25YIiVLuAPgLOTHoC4oeVO2kanZDK3OG
vzHTBEf+zZa2Z4RNeUxV2RXrZhXJjDt3ytbp4hsc5UBSA181sJMcUnKAslke
74SMvmQybbCFPl0cUw7sKa+0xdrceRe+xZ6+NF3YECWnp0nGGNn+CMPieAoz
KwSZJ4BRxONm/Xrhphv2Mv22hnSah+zeMiDQySxaHGh+rfyoLL0cS19ndeC7
zw7xYA0BNg60nygN1p+bg6kRnEGbDLHdpD+04W/30M80xh6r2E3zAxGtqlft
oXxz+J+JHx/RyCdwETKGsd4COE8eoLtu5i+CzGoVvpLAWk2AkqyyaHkTzQma
O9tmGIfpD8wJnlsko9oVTbjiw8D6hFIQ/4bwfMnPYh2NeiCA29vXeLs5E6qf
0fqFCarp4AeegAvc6Bsn7iiL7/QXaJfvYcUihdtj21YJsT7YCxYZ3KmX8it+
boFGrI+GtNg/PXPXQobf47VC3uuEUgUQ9Q1S+onkzAF0wHJfmSk8GHiOI8Fp
9KKOjGgEaSZQ59TkHeJHqRI6tgYAhjxtFyzIjDLqYhR2m3kF8l1DeDYCxet/
sypJJ2egc5cb9ZnUdfupb0dWqnCqC2YzQsLIEKVbX36XDGxuXbbVbb6c661M
AtOqrNNh/84zjB+uAe53td1pQGZlPkTU2lYbtkBQC5BbJTEupRexmfekLSY4
ZhgKHVZ1nKfIVThXXPMvOAAJaQ8IE9VspLq5BRPW46QmvlUzly775hkUY/bt
p/4fDuU1G4IfHjNQYKgfTueEVjt+1YRkoqGD8SegLd1Pp7hRXzKVlFYjo4aN
c/j6js0KJx6uuKAtgSNcgpQuK6T+TehMv1+ASKndjJXogpkRy1ptRFvi6Sc8
hbazKXM9SZmU6xDw4C/BBT73od4enZ7EUDhu9tjWr8EBpSx17jKJthn8TvTQ
QWHM6pB579aThhTCtKKG9g5bcW5INBqHvRDSfaO8cl31ksf/7+OGy30huGUf
7fommSmVm+PPlvz5vF7u0xkEQU3IfOBw+BAGic32VeKcaCvWNlRjwmwT2SN2
P3z58V7/qpxMd6ybQ1pNhiyAziGK++oLmUWpakn8lO8m1FDfQ/x/nBlb64ll
vLiNetANBoZ05KBaaqoRPu0wn8oOFcw9OSL1p2Ef1vHJGVojBgS7+hTMM1Em
rYTEyKAd1FSIXIOOkDzDuFSqQGQDTYDokI1l/eDXShlKV3v6nwa6T4JeDKJ1
JCjLSOaP+jfG04ALnD4lWBmdkWr76gFurUukmNVNnjJX5l12fLux1UbeNe01
8DYjHNzWTIJsNiIawPZk+C97gjzyiGwdo31ijQPf6a15Nty1lJpB+NV1yKRN
cCu3hmg6w12Teyef+T+Bi5DrsJsHyNXmR7Wz0ZcfByHcaVbWbvtFSrBWDnLy
0vrSsJGhQO9cIp9St7W7qRg6OqAV684VSGOhI4QtcWmUmpsXR2rfmSH0Nwf7
58qTwtfg/E9zO5Geoark16g0ck/vzwJYF322MsM0hjya9uhfRdvLin8QoSVj
dL07i6ty+JcxS6PvnlNK6Afo+0Vztl0DoRICSOQ+eACnyT+tEOhsMwZLXQIf
eLC3agHsKbeF5Q40O+gB3AiIfD/+DajW20pPM+EA+Sr4CrI9jxZPqVhm513O
0oQQQ3PZjBG7UzPbKXQIklaEiYVQFvuuVk4aYRmGJRby4JgwdwKHWoT4AWvD
zWFHUsf59OEWmQMZUw2ws1S+duXQWc0vf8sQhuSXIYFdbBSYMzHjcjkM1/zX
k554VnqK18XI7Llho46EHHidYBO0epmZ+cH0jnDgI7r3f6VRreflHomdjKCD
LNzYkQGjYVq8Ru9n+7vYqzwSrUQg123JW+1UFvFyeGyz+qRDrJUdwvCCGBwC
gfiP6d15olAY5sp4RH1RJAdeMV4AwgKBKyLeaag9KwUbgjJJJL8W3XFBJUXs
AO3hdOUZf8eJFesYH+cPFgTjMI5NyAozmgSFOGEAAnuLO21fIA6AFX97CVN+
+4bsbbO4D/q4fz9qyo775Wy3lVGzKQVUDUzh9T8qKyMfLjfJHja3wuxMJ4pU
DcwzVEpdFhpgb0PkKEO+UpVDWM1RZJotL522bS5Es8wzS3FqJn7NT5iuFvJC
UVnc5PFWK/qxlH7fRut6fvCBLDJk0ZC6Jj8sxzjf7VdBGZWBLtMW/Lulj4j+
f1ocm0kQ8Y1DR883Qwo41UGl9+a5YaYLckwyLETahYtJRsAt8MSa5nc+ubO8
nOSWjpVY2k9jWfp6M12vRzWuddfDfTE7lfrkRA7Rh/fSAFDYA35EYZPP2Mvi
I7TVfIhsD9IdO8zu69B9rzFCa6aPfAM2LBXP2IBtlEHrLN5N3yrWG9FledFu
3kmvtps72X7r+HgTvwlHBQ5owmZI41/mrYI47PEIBEIjbYr9wF4sKogCs0nl
TqsyCCjTffUgrNBjes2iAoG/cp2OUYTdJ58mLQXcKA0Hwb5jEcv7MReYLWkC
GHDmsOCqXtZ5OaURYAaIdWCCBMJLqq8bwTM2368/J4PMLT1Qfzg6dio8UwmX
zWLc7HLF7oNSi/e4GJl71+80mZRCBey1naGtt34FIDd2OeDPebsZbeLbtkti
zPJK1bM8xHPuC13VpzS9YEwNZ1QB5EbD3KjWWMmMFYOE7x2bwXUAS96VtWJM
e6Vbx1B1YMV1/zgaoFS65TV0q5967EpcLQuf8b9CW2UbLHZjpPIHl7+JF8nM
xv9x2abxRt+Xg5MwdfFCQkmlSjFUyTgk2oqkEW4TYUya3fGURfIQCCIQ5Z6w
ldtliKc9DUHlESxnB33jrnGLMeGEVdADZDWfoev80L3OcDqxKBUM57rqXASh
ahLtMmWr9x4zFhl8QVNe98mCwWl6JZWxYAAiM5RPWmzbnX4dmvoQeT5r+t4N
3SsvR4GxZq/2aBzRdYPwWZ8pPrCdarhN0H/nmWbYGG9mxc7c9hBB6DNWdJL8
KEr5tlIbnmRKfNDNW4okauCnWAVk32D5DdVhlZcs8bxM9e00SogTEIO+KMDf
y4lKnNWhftAdNqEkjhBUVSK7Su4aFkOWOKWw4F7aROxi+lLMljRnliCt3CYn
72HicXYp0qj3oOuOsZZCTeSGP2Q/rXMLQJzwH5Au9TVQDtuldAa/KMSrMpwi
Zcl2iShNVAiIflf1Nzq1a0xCpQIKhlz5r4DO13BY3TXgETjz82HRzH1qsl48
7VVwD2zF+y2QCfSVGIZMliUD5fjKOd+tAwIxtnJB28hFQVx9OoBQTSaR3xe3
uvcK9m/tZB7h6C3vleaTYshesCO5YYLsfdrUFMFVLf9Ou6cexLjy8Z1s1rKZ
8TLSXTyoHmDYqcb3P9MzcawkqyNXrHERCU0FXgnpCHBMf3X940n/qct6i1JA
7UTsRI3DOVsGGb2vyZeM5/afI31/6yM3vE/IramJc8VIx016k5103tvNK60d
xrUZgOPuMLUI1BVr6YONj5cwH0j0J/l/FbMrqV/KjF7nzIQPfiElBHlcgErm
h27jA550XZd57wdglPS3KX2H/UbjfSLN+mCzVJXURyAyYKYXDQzZ8bM0BcUi
fRl/S5vmffqyeKNgttzNEtGQ0xOxkVSHgECYibOIESNaVZ7Km5LHfCFx3uas
Nmuj6O7ineUmkDmnFgOKiB/TaDYZwi5joUdKy5WH3fz5hGpIWO9bMRRKxeu8
a/CsG+jlKRsw2Z23uq3+GUUGUtbUezhUzMTuHGnluh5zUlTn0LaPzOMvNf75
YedP/Z8pXpuymBn+qMBIvf6c2RdADSXlB7tljuWDxcUvX1ldX/V9IDBf8dXA
cifjYsUc0sACA+XYcyIkg7xNXsx1ylywAm8O0z62ZH0eTkBE6y61AQ6w4MI1
2kkVAlkeLFgN/TrUyVBENu3Ti74uUPIgzf35gSkdhLRy/XbJsc2/P+BGHjUE
o4bVruEPoR+KbKCg7tXW0nwI03kp70SdhN9YlSglHP0jAeDU8kTgouFgBB97
L9pU9B4m8P9danxlS3OLMHq16Rp9ciQKZA9A7IHdn9iyp8THcQbDupEQSMXp
ZiqRPLF6bX/M1zVJRIweWetrtQKn/+/W6XbaaO417OqLVeXX0bR68RymXPp9
WbVXwKX8kw9FdMWmwZ4MoMbkdd9yektm7gbVGwcP5MbrNl5+RCa+WEI8ifL+
aRsc1u+YJGrL6UMlU4g46rKIe3M3zILzmV2hX2j5fnazxvDEpU5ZPVljfaPT
XWb8/j8RD/E03TthoE49aiEsu7w1Q59FEo67hZBfHuzQ8mggP1UYv2KiW2Pp
el7xqo6AcKG0daZun1zFQlY/1mBOm6HIP80YB7FiVIbK5nAz0+TEjH0AVF+4
WTtK69bKxbP7oAlb5NrhV2ye+pctK15COQUMsk2cvmOoH/iEVMwuT+fFpbjt
DBFw3sosAxAOpSBJAf/Vu8NTWfB8yg4LHJFuBNVH0NAtixCDciH4Jznjkhln
m+XVMN2PEFEufwABCC4QAhmKZeQ8ChdYaQgcKk4sa6Wn1NznsDDfebCW/LYu
gwlBhFgQ8JTA8StQiiHu2Ve5jQQxp27vggFnmDACo+xDQSD01b6cCFQv/Rvn
LrCCo420zPn1FHNIeqW4omTCboI30w6i7/FlY8Sy+8W770JTf4YCDZrAJfuh
AfbQyIrjoidWVPk7xthjwL1d9T+KdJ2CC81GU3s4CfxjuzFQ5pZHOVM7PHnI
zJuKI8tcYZ/s4xUX5BJw0jhAmqR6qgQf6g==

`pragma protect end_protected
