`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
pVGgweMpXf0Bw6XvigD+ZW0fz0EbigbQZyCHsuO2LFpS2sUKdzl+FGM1Vz/eXGWL
Z+lSpbqPvB+UkLbkzmTHDTvCl01DHVHcuB4BwC7fidjLZ2LxwoQjdMIx6OsamNO/
fknM72WLoREjIeFQ+iG9bKgeGCLjnEfuDWaHltR057M=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8544), data_block
DeH0lDgNjPqaRiJ6vtXmNlGhPpihUOMB/Ds8uPms5M0B6Vn7cK9LQGcFcO2TVxfe
m+iki0iCioRvhXqB6N0z+YNMIIl04TLfp2VXKqkGrfaeFamKgaNFMdXQhpQqDJ0l
AqQUu9E3zohDuvjXHEHAfM47nZq7YpZTgltsMsUdxfxHGtvT/0Br97XQbdWuFpck
nnyNkiS2qd5xXcm3I8nbDTpgbC8idQblc3QFjJLX+ztnH23YVGazILmdmnCP0p1r
R2J7zIPqahDyjqglQLiLhtm4tRJ5Ddc+ZWzquzw7YQLg0CdmIU8EpF0Dqy1KtZx1
hkD6GB0MxMHMwnXlTm16XkxJnLNHtEDeVUHsjBNlTNfs28XPdOW/IvpMJduUD3QH
MW0m4ChoLzNmDUamn7vwxDpSGATmr448MTVUA51CV40wxfEtXaD5DwG1jYB+yOby
S/LrewNEw6BJpDpSOpOO5PJZnURWAPMawnQbXG2Qf5WZ3kSTrufBGGnU4cIL4wKd
CA6Rq0FzHIAEQAnLzyk78ZM0yNYVLicgTGG+VkL255i2d1Hf6i1UO9KC1+Xg6vsv
l17JmYVpQsTLxYqezXKJhZJ3mMG8SekCAEsW8DBF6WuYa/vQUEjX02cYitRnyUMF
6cs7YzOnPkKFTfJl0xSyDoERRqTbgW6MsCjM6llI9w6fZ8NpUiDRMivqgVLIzM9p
C8PE032cFjtwkQWRGtj2OB33iIQaZ+8U3tzq1MlDLCLe9eokVBSFX+sHoDSQd7Sn
mY2kg70SS2hbeXiT1AcBWYhsrkxWZH1Gds/gcAjYxLxRFiwEKV5aIBEGUEASckaq
VvekHifvIIazzFuYW8atbWY36Bl30HhsKaxVewSDzdVv1aIc1MW+s1cf2zcUheKl
bCGtDFH2vGAIbtOyVwX4Fu3KK8hnio5af6BOn4DaOB/Kjm/lyO5Ku2Gpjh1Apcve
UzjaaBdOnkRw7Fg2y+Xrxzie7b2jqCB79P3xxfPmCGGDyWVvMuRJ78sYCG8AELr5
PlKB08nMj+X36tAxOFHVuTwuwFqkWXs3tJT5aluOvDNiIWLddiilaZNcpOdB1TMz
3TLID6aWUQun4v+ZF4dFmplx6HEJ6ffoSDxZ788kLfLhuevT9JE6XUIo+vu+X7bC
1Ur0I7JI3FQrn0M9+GGxkLryrUrqjpeBeh5He1iUI8axNXsEzGyG1exG+bgRNUjx
S7yftLWVG0TQQf0avy+wMXYQc5t9IKH6ckvci+GwxJX9psYVOMCieidXx8V/s4Kf
yJmuZyMp/6ivxRIspb5NUxwlyJ+eQutbtT75aFXkBOZLw389MYuvFafloIfJ0ILg
cxh+lgjuqniSqbN76FIp7z4/A1in0qc5aZNqhnpqDOKd0qh3YvUcf3qtz0lx+wh4
K9YwmeSLKLK250wKJcVpvzIP7mulF9Ta5oVikIUzG5+KBEbFBKQ3Lrq5JPUARu6Y
epNQX88qsyMl1idWKplI3RMnj//j7f5zhQuzxyBfYMp6qLcsMuvkV6hwzofqBBjY
3XqxzehxjnZ6GKwabWDBy/dtD987gqJVkfj5JT99CtjnxZD512c+3kgPYVQPnWnt
bRnpJXN28cb0B3r7XAQht3QfHaKyI2lQTo+9fCBrFVUhsquJ9H0k8oPB8wnSdlOC
ihXiVLg0NqBouTjRSc6SNRekGS7eZW5lTdbgTLeENxZTWPProjGhNLAlxrz2Kg/p
h8K4hyFChcaFDZRtfqy8Gnq/8tmi6SWAfYcrQn5Nu9+vm3W6f6bRNzN/VJbGpxTp
UGd2jzVftqtxody6IwY0FLoyYwN3xcvkxS+vaofzMRTjvUlTWKSDdeDaD1eNh0/d
bkUKXnD52sN052k8nqUE5TYY+aOIYIXm1XguT0DgY0RxJFCBCdh/VMkl+3qqqfp/
lBR9qzyAr8P04yaCjRqUhgyQi0cRgCoJRIGPT4dzlnANFqc5Fx20w/M+z+W6NR4p
0Cx2IkF3d32K3N2SMAY7ZCakxjzKq/Sg7GekEd6tmKAcTubh94cJHn5mkj6KidUK
2Zx45i4GIyuUkKboKe8DqEY+spVg8J4O1we+DBn1cohqU2k7iW5kw4qABVS/5Dsx
AYqlGJKFcUOEZ5Y1cse5qv7kU9oKKC1vn2/EqEEbUtu1wi6kVmiR6D8YSEFqA13B
G8hbjKxhPr2YukXKe9vxV6htwB34YOg5MJYueRDu17fnFJ3f6jS2Aatpakj9p7Q3
NODNtnIy60BRKUOsOnEVWtPDxflvYQkx8lhFrneepVVaaeT1IoLtVCy47xE7GC6X
RBzLeNPkmq+4DrGu+NmGBemsWUjniI8fQnzGYhhEobN8z60u0oiYvz0fdPuXJnI0
3RL9d9KSYHfXF2O+HEAP4ZNreUR3AgtazaWrO4Rq7MhOPY7JyQUgD8YwEJ74zjCB
t5YhLbI6UiQLgqTgZHi+xT74VEuM7kLFQhD6BpVF/GwGnKhmU7H5XDHHx/sxg2BW
h2cTCoCxAwAV7cFwWI1rQ9r9InjdSUpLbQKmjw2BKigVrBirDMyc7TQJhvEjbKXi
gMyBXeeYt9v6fJ3/AParU0SxvXvYQYljQGDeooEIJOnBaYRwPWO+7UTDPlJ1gxxn
6XlnIKLeVOPnm43LWZ4MxWd4ZMNRbsQIwFvpzWlwMHmMOTAwD89SEjhGZsjE43fO
7x+LvBe2Fq1eDdr4P9ytfrlXLMNWR9rF04bnk5jHCwjy20efg8NiUQg9Wu3AKooD
bURAhDP90+vRyL+pMs8BQl96ubsuwehJtR8XIlvLmfIS271K8hFupUngBDg59Zaj
D+y27lGN//XLWLrcQrfKe0s0Egd7c2dB48xl4+RhzkVKf4TC7fIDeTc0Tq7RKT/T
3sTvftNQDXOE7gb5w4SIwiov/opMlNP7IZrqXcyq/ScB1hIhbqr5gbO1YG0M3m+U
8TalcnCSeV1JpE3hPkH/+Ksj0aTTioHfXeqb2ikHqmCPAN2hyuBP/NSSj9ryIhYz
/3lZXsRZ5hg6AMcDzL8CKRcaLJG7dnArPa6+/XxrloJgh5EtDmVXAtKR4XblXygD
t1ahfOJgv+Q7FmJi+6y/RK8lYooEJFeMbpTbbGrruurKpw+m2IOH5cQDtPLrcEqw
2Zwb9o3Xn/hW4JcmGvT4dVh3FUro1ZRDv15tLdHtWqkUZ54E6lChzcUWuk4eXfob
Hw76yb0x0RLscdgLXs7YCcuciOq8b4nKJBu3Ha6CqynTZDR52BtYN6WpN9CN9bgU
CbiGqY/q611NgIVJkW5TyDgByJ32HsanExHee6NEgOY8HtCcIWltKdtVTuMZq6Ej
zkN4DtvN9hlLSz5VdUMzTsyw7XVdUo67uiqmpJD8HJz28Yt9vD23SZZMoeObGx3a
3DG5p3xQ4Ovqa11V+blaoQt7JWEDQgUK+aPeS++wzOdWAFHlUkwbB/AGODv+64lJ
fVBKoZuP/ADo0XC07CMR+ko8pmRD+pOUBN3qPQy0VI+bedKdLX1WrdjiO7Qn4OL1
FFZ73MTKV4OcNB6a9Ci097roDbAwPyNIVrNRvoEshN6aW/VLnLTi0SPxiQkrr5Ni
yqMkYG393ciXWT6WgZQ+xqWENmBZ1TKTGp5oy/j9fYlunO7kC0J62cEc84rnavke
QmSN5JSBL7iCb1b/hMbLP63gwaRFYEq+qQVmAcosXSBTS9AWJJrHg/7ivQhFYu++
gq4qu8LPV/WDVYlzGIbsxQvP5Kc/NNKhic5xD+4p/8sCIDM/Gc7Jsctxz/TCDRQQ
Ut4B6JcjZzSGXPoQpeit3WI7du80pZjQmB4pB4FQZgikaAVHIp1IFxTW4JxoX/EH
qjABIWMROlHa+N8W3MSBNuUOWWhn1VSZQfcR+Yn+NtvC8A+dpyz+x/lOyQd7g8+Q
M9pDA+W04cR1egprZHdGx6o1amW/GcdTFRVE8Xt9+2uSzjORVEq1iPohgaLmZkMu
AJhgeDTDkUIDs6veTG1w+ne7lA4CgTMpATNb9aRjmgF/KZ6cnwK4gFP5rKv29GX1
RKT5xZlV6G+0KZDg05U1h9av0VpK180KE5n1RX0wWEDsm6HjsT3p2wok2cV57MKb
VCZyT+Ns5gbzXtQK11c7PdcR6ObyA0qJw9B+iIZLntgEHHDDnDyn3hAtc4XxnSuS
IHWsytt6Owb2UrR2sKjYUh8C0eCiDRIojGUm6VrLeqv4kJXAHdkwMRx68JoEJG/r
MeoSEEgqz+1e0sYSO0vtRHeJ0FPbVaPzVyUNZlLp3ivbC8KEOjPYDRm2a+wU6+Xw
tsuganjsLDcmmSJCBLT3C6SaVUfwgwGDmLC7pBvQbn0q+vF7VcFwdlMT/ag/ypNc
KqPN80meLPXZozpEu9aPAUAmaRW2uftqucmrpbsj7cZTLe+Qpl8RcxEtdAMz1l4w
PVTZq9FQ3IinN1Aa7mbG4KLEUfnT5dnSNUcOZDQ8BRU8hCbM3WjxlNZi4CTErred
AwrikfuYihV1n7lJiA5yqUJAHZMswkHVYIgGSpisPOWXVd/5dELXg+E8hG4n6LBf
vBFVZrh1G5PlnNmaYyQACItZrqDGruENZWnsQrHUZTIfaKHLWAm8mZ8wLtdD5TgS
VeLwXDOYwKlKOv8TZrD10PdpczxbD0L3c0K6stWNg0EgdHCO3ob3WwajsG6pl8oR
8f1FLpgB5PADpQa3Z/bM8bP+gwOrIx6CGmppeHAmzVPGCvYd9JUxucA2NND9SC8y
Tq24cmvTdoSUbPOk2Ek5mlXHItGLiBd3sc0WZGtfIfCncmcgozAkivWtyWxeoDZR
+NJetyZqngJtU+HfFM6XJ6gy0ohmkezMQcQ4PigwjCxCclqTeVsGeSECmIU3+h8f
K2XSJxiAbK7FEqNNrWJigUrmVg7IoMrSjY5BHDmJjIcM5bLm5tNHcUqsQhNJvePL
1L9S7kO8AOWDEJrLybev2JOZkLZZoNpfIPtTycj8Bd5YMTp17h8ZUIwzMkStSIXN
HIl9SJ9jjHkSNILOsG1ohMfGV1rrx1cMbvZBwb2wtGZ33IlDPJzcR6F9JtV3WNkc
ysAYLRtaYTzPzZtIbr60/JdxHXKcOtBhheBbctB7HrstBcqCTpR1InibCeMdeqkb
myNwco1aw5CtW1timZdmzD0CouCtvfgpGZBqskFLAjoCPLnznSQ/Y0nwAgj/DABA
49Rmshf05m0PVXtVK7Y/nmlQZbEpCt+Ffqwj/w61pyHibsNKQrxtvFLM2dwAqvnH
n5VaPgG0jHQH3OE5mSt56hQwvEnSNEDaumcmxHvBzC73ZfDULoTpjSZwHLvwwi02
95cSjDC+s6XADRry2kEs/5Y3DLfL1s/1M1TlQTsQPYFgZ0MpxaKvyJSTEG2iEk1i
Ho43t95JC4LXeBnqzf9HvS9DaGz4b3X0Z3kQ3yyikKd9BzDQBbmEC1T7q6mwQRN2
o93ux/xZ3hPvukW1Npsn+0QnBCyjU/bAOZbgmfJddww/u/OlhytXwwTv8GKss80S
fPyRxpgs+KDkHgXubS5Rn7701WXFPrHYDTvgthDCRf/4zuWEmFVFQ7VN8vBZ1W4J
my4IcfC78B0oK8pUvgBAOclSXCPKHspFjBGMcHbA4VKTyIbVWT3c0yJiHGC5ep2I
qLSvXj2npT9hNT6eSfRIrxQBFO/eO7OC9CKpML6E73PiP3eXJd0b90+cxUgndTDS
vucezr57e2UZcP8nryDIhu/bSo3jJaSGjAqZ2i36ZbPkOYUv9u5C4i4hmNTidc2J
Nf2Cb8xyw7BpyWseF9NXR3YTb1IJc2EtuckgNUJeU56ue8/1VxaK0muIIeOdoOel
bcA52dXnU4joviB8q5iw9BbMZ/SXY/fXPAdI4HiWXaoHjDESHeB3h9MmQFlu2QeS
mAP1l8QoPUfwqNerhf+DNCOGu9VvtNTKn0pJtAwjEEBZemBsYbn0gPKQsq58DNwg
tDUtvifkoyUOfQqstN50J0aR+B5hESZQCtuRyZVTEwrzOxNyhbH1wkhwD1lecdkY
vzpKvzfYvecXiXTg7JhJcsZYthGnj7y0CkN7g6uEDr5gS2d5w6GDEopQHDEv00/W
Urm/MNzEbbR8IXt3lp4Pq/U3OW5EkF81QzNGmtah0eCXBv2YCEexkRN7RKFayg5e
wDr3GQyAaJJSM7cFVx9qNFu4CRRCROg8mHLW/ZcUOAmBZ3WiAUZCF8L4rbKR5Qyr
gasi3SKGErixs5kXBXoxWl9Nm+MzFHTyhYFDkUhkAaBZukbxSgzAAIz3VR6kZ/El
SMJoHW4WRPWeNci2y+8v7lqYW3MvfiXlVJz2kvQyxoWwCsi3BAlLNbhl3iMyBH2W
nbjpHjDadnTnH01QtwX0h4Rjr/zAut8BdvJiwVayXSsqoOxUhop0Fqhn64PFsIkE
Mib9Z97QS0DKLtLaPKvnwGekJKcWcphsCOIT4Lb4CWGAdnR7Oh+2FG8fgsxqC1Tq
UBmsXY4McfXW/TGunnHiHxyxw2JSzYd3biyCWzB7kgl94EnIF7YR5472VT4nyjZt
XL+GdE1omkxZxFJs6mk0gK9O7AcPBrel1k9E6l3IjchMk0WNvkRpxiHidiZEGMCJ
kvHj3WFQ5l/SIFz0HpitAXFocPOAYbsHKH97i2w6FKRyMN4B8cz5uVzaFVR9R+PV
qREGL/vRWhTG4cs0BUWA5f/evEt3r4g/nQCCQptYFuRUWSz5hLR0SyeAWdKAyhXu
Ui73VTO2UKaW7HtBGBL5OJBtXpY/XMhKvuq7X4w9sAbOTiYxWekdf5wxOILJCy8L
Bmo867YFm6btsiLv28Q6OFwvjU8iFIck+S09bCLXxXMlcOc7xjziVze94NP9c4GP
LN2eAnFvI4JvAlN0VXqHHmRdqyR+rbb8DxKW4kjW/OfmN4bCIEU9IkOEdFD2OMcv
/mh42nDrTMZ8faZaY2iieGxYx005LxVv8hSMMhv56RmlVYs7mRBzlAE9fX+nEwRz
TL1jyK+bMGfynmKo4uXU7TStm6zwnShKV0E9dn/Jt5O9gcr9sg+i3AoMlmAdYv/y
H4TEvRxJCvlHnXIHWtqd2/C8G3mJ9JwC5rJe2nMFbY3n7YhQ8kQzlPUA4QDaoPMi
qfxlf4c0Vk8rs/5C8+8bwQUErIcW4Qusbq9ZfI+hb9Ae88x2dEJyfFkkfVak4if6
iF969bncH7iAsKYyYGaaKqMZBZJZspkh0tBFKnrvuxsE/s+TI/qaJjELt7LX4jXl
LzqsFyiXhU28jdKMRGIHhBqsiGZxch1wdMwT3UwQMz2kywqZSg6N8GeIrdMZzuDh
ovNEghW7so/SH3xbUikHCoS8mbhfh0h+JFFKgtZWMsT6fft9OcQPPr5piHW6Ao5o
6ex5QiRhbKh1xrRtYd/VsuMVGOvp6/QTOV56YouJuwBMcltp6153tOOvxA4lVBEX
+/yGIORGgU9QG8V37ZmExkwqrwXhuwHBUEu+/Qmh3+JAARZKPkc62EPsQvaB0A7T
BrdCDf4WMAiYk94jinV3cd1cQG6w014G5EZ+wzAgyt8vOEilcSgmrTsub3gNJvGZ
IsO8jzFTZ4U1MhGATy2256yvS3cys/7GKC8g0IpNhzbs+Zc3YbEiZqGz9asKblGk
MRwxbAWd4ecxVnr4rxADnTwYmsTgtbld/N7QFssDXuMqAOUoi/w4zztwAx89NwQM
lX3gOCYsAGfFUJwLUzG0b9r6cstmvwbut1hnzxWBrgTmOBdbm/ZJASBaZGM3CJKH
Oynv3/LrcUBXwbwCpzJqZtXwhdDp0Xjt7uimM9e46g+iDJ714Aul01o8pguK6KUH
LbNVpJolQIeiIxNcJGIy9VZkLOdO870x2K3+gDFF9KJYm1z7MIMPrMXMm9WSfKgJ
xRbYcA0kxIXYLfz5MoCvpoTsf/shVrEdK1I6/WxFYOdcb5O1EcqjfFXRJmIvwEIp
pyndHqKi7foJO9nir4kwNDWV10WHT2wgMcVuPI9ogSkRPZqWvb6MPRWsJy9KkiTY
X6A3BZmUSXr55AKs2LO/0Hr9+U2sYJEzRlgxSmg4bv6J1rsSZ5gOzm3N9UoV05bk
8cigjwPzlBAKtQMMUwM67smaPD+Ac/bJn8194YLn7Kq9rqjsuwlR7j1k0+vWvYjP
EdMkRn3U3pJ0tfXQioxZzGKjhlgMAHOFy2fv7iGE/zo4kNTFCWbPdvQVbJ4eo4VV
13mfV6tXZrm/c1DaORycJd1H868vu31WZvUT1J8fkPT7VASywoHy8ga/Z/HH9tmy
bpFRINkRZQf1bl//qXrHt1axcPyZAFcioqZiKRI6hNJ3Hf0X/2dxaXV6RniwFNjT
qr0k9ZXIIEJ9bzAyKss7rI73Bjl4G7QsasyX7q33Dea+kzNfcSuhfstCbvPyg1Sa
49rvMyIjFnNPFxYoFmRAE8sZk3eou2cdujkqnVo8V5vrsrEaXhGrlEBDcRHC9KGd
nJ0IhkVu9HCkMC8MtDwvmI1GTp6bc9X4psJemvLFikpajL9/hf0/5Nyxl3J1jC/j
ncXNsHjFzMQZnuQHlxWmrjeZeV1XZ0zP8lYJdw3A9swk6sUwwdsgk3086KlrjriB
U5VdjVjvArjHA8qWG3af6UrFI27YzPBPlFPcDrex6k8c/TboR+h6mcWuNSXJeex3
KpGJKtBvuk3myo4o9e1reMeWDGW12NHfvW5FfbiOVk5+RzhhryZtKf+ce4Lvt9tr
6OZCYPh+JcmF6DnlXH0nlbx539gb3gAhlkp2ZNNMCDXH1SVyFeqNs3MF5gl4V/mI
4OqCAadOBxZqNTZJS9k+nLuQubuq83u0L3fMiRFAwmU+QY9ySOXAJ/J+ju/uD0AM
oNadVvDZcGslkMRnfYGMbjCvSoo6/XLXRkhNs0OLJn101FiVGI7973nrYn+wJxVn
MaZICCExuiCkX/4yCOTZ0MRafDCCsYnLY/ijq78rE3nvZEQ3JsRgCnmy8DiFHbNi
j/IJE73zGb9+CuYySCKYZPHcMusRqI4g70SNDhN84h/7opNPqxg8hOQftb5C3g/S
az9gmOqt620AOlX7YBBYHLgu6ICre38BkgV2rDxYzt0LqmJPIwKmkfxvqbmxSUKG
5irGcoR1ROL+Yf9d5fj8eRmEiYYk8zdl1T2q2iA9aYcEH3HyjUnxnh8v9+cfeiYR
RRwWp+4XUw1tpjHuQlBdq0i0mfDl9etvqEpz3B7MFPNwmhYT/d4aHRSxI2eos3Os
MLMDw1a8Wvub0Lhhd1xyPK6vky0Lp+ZIyT/AjHZpRpcnvmfos6eTltfKAiqv6sFN
bcbe0t5MqGPP9Zjll6X9q/2PacW5cj62w90ntn1hJ27KjXOCK81rLCo9O9Ttg9gJ
TsBGCDrJ0K4VDENQoN0KVcZfDld1+4V+BB0FAxyqsXy3vrOQp68znNmu27nv1fTz
ZF0tWgoFOaaQj6lWcQlJ/JzFiHi90NA6IVP/k7qt7Zlq8niaoAFmpYhnq9eEhWTm
hqCfG2AijVqqEZik1HcJTbMRTKbCIPTnWClzQjyCcJn8vkvUfZyH7PEs3tFJ+CVn
NcW5uiczhUvewtbcuBBAFH9pz7fPsmzDfKIEazjIx0g9fr7yszckgHpRwGInwnZV
jlBiZ2fa3ncfRCu66bZRyYtFOL0SBZytzTdYpAmd49aSQ3aOvQP3MYtzsm0c148Y
DK17MxPkFdMiscqrZ6tT5IDrtEa2ttTPe+qYDU/zekUrixRUoksfGkeZsqEFvvTH
WuhPnsp1uXYlz7tDMFnX2ogZk0bBDuQodAJ+VDQWsV7wPbXSyOGzZLXgPj+yglZD
qyzbRTI4OBX365dY5O5wq/6PfnP8HB5ReoklTR1xAgJ/aVeP+yKAOKVDOGrC6d82
qEng8L5t1fA2tnJHd5zdMyNYu6pgRPtCnGwbYAg760bNTsBQXBRJop9cELXU2MEj
TiAgKGeB2B+hVo/Bk1jkgtZ9WAAdUJQsDtkWYTnuTt4ec8kLdRu56tHFixxH53UZ
6DUwfPpC0+Si7pCjiXrjyw/UoVxm+xgmDSDWFCFquyuqCdLiH8dGr5qB0pRSyc8L
ErQXmoC3CarMVs6mSabJdEffumuGiTVdCeeLx2ISn9Gg0LYyNaaGyyqeyASr8G9y
ATP6GG33OqfjSaO8ZMPlONnJHj5sCbthkaOZgdHpOn4AetlKY38QfaBfy10ii/bm
n4GahFztm6BUY8IF55X7JafLhqjfVxiJSQMkWmXZWki/6NVcpdyg4QlJ5y1Vtpzz
B4yorNa3OTU1S3845NLMB3ita+CxAL6Yud8npTPyiMApdNxX/f4O3C1er7Kwaozp
AfUiVa2QBKAIzQnNedFWguvFFQ3r3w9OJXbTj9i1/S/3Bw4wb1Oe+3fo+q7gjDMy
B7ejzbefyMVYt2KpH5MdlkoUbLGrzPTcg8uKFbkLT1RqnvUZb57cN29g8Ob5rbMb
oGuyxPNtNOqPrxyhXfQqS2fmogw7HPkoVNonqiyNTlFEnsKpkSZESkRCeYot6UBE
IXkh7AFo38DrARG9cTt2XasNwa2OIjP3IfDEEuOthitUyYrOP1p66AWlVoQHBj05
m2dws1Rd9wevYH8aNeKrTncHsCc1Vr/l3+Th30Qas+6ZwS6xERJXwpmvIfd26ibE
DCdcxBhQlq9VV1foRNKTIkzIFv/DpKacIER0gi/T6Ux8ma2W+CiCVXy6IGSKU5CC
JRfteYFqACVotRPAJTNps3N7zIpAlfsGdiMdmD9oZ4J1UJ2N2VBavW5YYs/UTJBC
BbAKAYfPK50srzdsthHyJDHUUVyPjsJJRZgCqSYKvolFGoWmBOhzpDR/6Jj0Fu+B
TE7zsjUq4ORz9goeKSvna5aVxxzfDX49rNIIu39nRNIn0BhC2BH6ieWvb7UtMGja
QQlJ72ttUlDIpbpomSM6jJKW5aR8yZChnynokc/UjlhUfHv+F3mGo1oK9Han3ksi
9a0WksEv6jWQYkl+6tbSrC18GcB7TF51QoZCKBitsX+ej/WogJbs45/qjROnL1tu
dnlQP5Agzijaew+4DzyC3577cF02XYW03OaLCj7m8eZ0kiukx6/ohcESy8Jf3uz4
4FGXvrwilrt2zkCvPeVSDGrlT1rFmIa/HhKXP8MqHZRA6R1+Nr7OTpvCjCkTL3vX
zg7M/3wv7vA786KZThVAD+wiTPU7QwjAYNDhl+jA3doVVurN8N+HOVhBHNPtrp9C
UMKEWVA0MQE6hgz5BUzEGA/3gRH+xp/gmjS2nbdVtavSPAhwHipdNGbWDDtzY71u
X0U1k9yMQEHUJw6U2jib2DJsx7GbuNi7P319OT1ffET476hX9FPEqEs53TFKmEsF
AQCUveCj6p1dMYXG8ZRxJUM7RKofAQnYerPYB3QRBmh93+yOddJJdcTvcVkLTAxr
`pragma protect end_protected
