// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
T7fVtZmA1bi5btLVVBkrVj68RZbaZbDo9X+aiB3RwXnSWcKHeYZ29MUMFYf7t8Gp
CcFauzgbZ1FF4sTqu+DEO/ncmm72vh92sBPErsmjMUmPrFp7P1u82rePzqcEfK9r
Yz9AX0yzn5LXYcdzfW4UAedcqzqZVDR6MJ8ujBEaCOo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1012928 )
`pragma protect data_block
9GasDXIx9w3ejmDtTZJVqLdfypechDJPIhi5zAeuAKtvcu3a3HGLLEEw53N9WTLv
WtB7ZKzcAzX7aNCD5Q8+MqFE+iSleqW+2wvsBRFJOISHmgvvzBrGVBPpD8X+EiM9
mLjCDdrPdm/a8IWozFu+LdYLAbTe3e0ctnPebZD65wQj3BcazooYVWkqODK8i25c
j4OXcJyGFUEEU++viq96sKHTiXl9eN7bRuoK9zJJgFaKtKxZd18TfZV2bStkdcVx
7yYrP90BhtzsgMLdOU1u2/5rRimX5VxgtQKpdbiH8k3VGIm2YYBmJKl3tKaUUThJ
nkXTHP4k8v5eGzumbX8gCOUw2C+ODLSTEFyG0JUKxekm9NoxnUD+r95M924gW/8M
B4lHJWS470jjKCI/5TukV0hFhC6be2pLUEdlaldRM60Q335Lcs18xQRv7DmvJJx8
2NkvPff8IC4HvgftVvOa3smpnNQ+LOx21YMaYOzr44jrXdvHWS1gvrfUt7Jbcc5i
XVazE+sUQN1eBbGna6Z/NRYWnxepC5ez0DqBEE3lFivhXYFWV9bhMzul0KZb5nkb
Wkfrvnnz19UvYJxq6SVV4GyhkXLaWOljLrOzIiWkTjcelkDX2Ln3bnp4irr5TBcL
eXaKOjlT1sO7Qwf9IedhrcD4rlA6PhE0169pz+pe9lHnFeMOQXTzAOOajoBg8I/Q
DeoqDGYPOg0NuFHOwsU+nLMS0IFocajqJYJcCRWsQrbe08G1u9PJ+cxEQfbU9tC4
7G/sjB3RCKfAwWpparGWexb/b9O67OBROrv0syB9WxGfhRWdhNHa3pvCOWgzQJQN
OEp3J+urYdETLd6SMvr8qxN+EqX8yZ3QKT9BwkFjM7eBwXH/nmm654iK2JF6i+A0
5niug5FmNGtvRLZOzFuwZjgPnUVM+bRnZFvnkAsF0JE9YsSqWQ3s5h7tWTu/+1TU
AGzPaFaZZJeW/cQAGNQE4ye4GelL4MtDy+o4WPzQLRSvSQel8b+XEbzTwT/7GVTP
A5pJQoQ0N6EFDzjudb4VIS3ANb+31J1iJhc57WwZ529+n0vjzcIvGkdAnAawdn/K
LGlKPGlgD4y1Apki3ASpjd+tvatEnRdKWEW95/ldJQZladtc7J/DC7ztTKywxv9l
hRhEXlW/nGW3wTgTNeC/7JtCoNA33CNQxetSc7aNwbxhyW1XWvgQ8DKJvi7YJFBd
o/+a5xMM66btcVj79eA7cmQ7aPDFA9Q2upyIH51iltWNpF1vJ+nxM0icGzUNhRy0
rMl0z9o/6iO5dwfG5+wisHqeisQjyXIcMFvyhI6GbE36qzq/lyAzF+jISCWgi80V
9KGnK+xehQTKVhJm9TvGZuS0XblDYP+EfT3wSLhvFURf5mStbhM3ys5FVeo3UiIo
XFxPvI1nOddg8G90DxXJgsl2vgYUUnvT5x58nQgdvg4Tt08SIlIcGehemxjobpNL
nGzrDvvrGvbzRkA0ezDU58hSbG4m1Az0E4oxkffAnBn8uxD3l1nmPoui6S3e40H/
IKVI6gEedxO8mbcfNBpO1XbXw4pOiUG980tTDKQJI8SmM8VwmqnM5leVSVVpnV+c
whbarkyqWfAdwa0Fo27mWRneGzVKjd30u8Cffjy3alsuPRv9AvMqPwtYnUNWjXAO
jnmqk7KMBaLFqBlVWrRtGYnFSqQ6CxXjUW72JIS9o85cgoy8aSViqEta3GQFI6ls
vYnLF8+pSeJMsvmTloOaeR82CjnTRILya4ubZhTOFRBbobIuJ3R+3FF2LywR3Yvs
CXTslfISJ2e/EHVCuNErr2GdgD6+Z46OieaLLIpxFHnbCLIIEuzbahkW/sfqpzdH
4FyXXGM/oblFvgtGxR6lyX7L5vLATj6jpNmO4ZCbJCVpjWPPkT70TqY0LCheiz3l
q42RlMipNTBj6NDfnAKHCh7zd++t9GN3QHRUNNg8v9ib9B6UevTSkJMsGBDbJIrb
OI4IcLenc36BQhpJYGbCHujiwqhbgciPXKqzD8r46kC+z7DRb9VyLdbA9ffLjLde
A1Dh7D+eKALQJ86Mkh5mNi+z7JF95WqA9/Nyi0Ztfn6Y6fSVTJyUxKRuX3WXDdFv
yvwfKv+0G/5ybxZ60zPYK7L3QdeM28DwblW9Bnp5z5F5/CxPEtZ1jLfKeJCR3z1o
AnoJoIpCzlPMLF0b6k33tOQxs5TELFF6bXXVbYSggrjnzC9/wPY4Brxt36oK3496
kwlZcItLgXkzL/FcvJ+8FjBCC0i2uymvABy7ZIy0PD4/VcVwv/YCuRL5QqxjIvSV
LeYD8M5ZHMzyCFjVcjCrGtby4DD0qHHjQ/WKPj/xBetppfhWutQxFpiDtO+9nHhT
qiRPXE4EORLlNAM3KI4yAk3rpvQzTvlVrg9lddgxTLz1q0zKw5G/ubK7zEcjbEJR
MZrxPpBBak7iALywwRUpJmaksJ0PeyoqQbXeuOkLIhQLr89iU0xNouhviVbgkfae
xHM2Wo7N3KcSp6IseCHBDZ0t74lf04OkovWYQk66sNiQvbsyGgNjRu+B37qwLSX2
6y1KYW5vE+9ggo6aO2/xIdQY2wFDi7zVDHU4bvD09GpgbrsOwf8Qhev5udmvBr8x
ojNRiFAKuepvkJqrcNXZiQ+tdgBh4fuOLQuKNqDdEKWAxrKifRrM4LzQmRzZYiMM
5vag416w4r8FIk69879qMDxJa7rRHyDIJvtslKRYf5qz6YoR25qqeYn6th9TYUDI
v1/Kku7ST+o2r5Dsy/+HbFv/Y/FUcz4U3eK2z9yu1R8E4iKLrLPE/fgoBrY4KSGe
tcNWy43D3CNegnGAyjzSiyhur4XPx8kkugEiBCoi9ejReDnEMDgJLHsuyR/bUWTi
w/kch1lV6AxHDsAMzyNJN2fr5orqM2Hiz9oZBRvlNJbk+gPlhd2S5GwFsWftrdJ+
/4Kn7k/qVnJiyZurlBdBKb+A7z2vwqOV17+wv2Ny0PZiIaEEbToHcRtgypVAd18p
S+nq0u4/DTd5kfP0XqdHqcJPWObgSa7Ku0e7E7l/Co/1s+PQNFrlbQ2Qgm84j9md
ccBCwKSP/XYj+Ec/WGvgpul/iXJCNRB1711hfr4Hm7HueEPGNh3yA+TZ70Oas2a9
1va8vTQ937A5bzhnMtjYE00YoXt5ccceX5qzg383jWjFW30LuQQQf1jT8X8pGgtr
MzalmU1wiGdTvlc1Pyee+jmjAcgzBesgOBfxOjHa7NntRMIi/towgf7to2tX85yH
H3kdn59gyeBEok+DfTeErz15LkAi2sP9j1HVzdWrMpZz/NrGL4R1VKxu4B9fBzI7
Qn7CSCob3g4rlaRG6HZzGzFeghYwVnQIEFYIH1pMf89X3wf2rbJwVwo4XS+UPif9
ijCBTojkXHsR4TrGcDcIFVPK0U1+g6/l03ogAgWqXzpAogKsfN6CaymtBgIvdzq1
8SbzXMjZzxz3Vw2si/PLl63FNzT/6Tr4d9iXk8RRGycqF2VhbNCkDe+z2nxbr4+L
MUU18TQmENrQB0cVlDvxzq5YzMq8iAiqB8gUn0R6r+qR4yafLE8XPQQCNXMFzU3t
M9Epa/PWULvuGizyCC1gUnBNB+UVGl8adRPFaFnVXusWxhgxZ4rhKw+Lud2snuHf
yxW9Ex+meuznBzLHHu3mEmWjNf/bCAV3ZrGphNCNmNDCSVI70nxE4HvgxfewdDyZ
kiql3tCatD7iX5gRv9XGiS8MsCiP9QFAzbKMIRWaajSxXHAQF/38ndOOmCmhkYNJ
n1y1ARsi3qQWNmpMGwd7xt7xAwX3srhjfxr1cZcCtJmpWb0ihyQEIZaNQLTAaGzS
sFW1x1OHKGfBuWmCDcHfT7jYOY9/ttFu7bGOEIn9EGRv7+1z7ZIkW4T1FcnZ8bDg
Z7vUz+gzMmCybEJx3ZJZq1MRjmXJ4vw/2tUTr5WKfNJqFL4DZqnkZP0vWe/Ex/4x
odKLVPFBivTrnOrv6JujSswq0fi/3yEmoEMLz7h10bgWxD3DMVDmgdn7U0+2HKbO
Xo4JgeRScSreBDn/k3xZyNQ6ydO22PWXXq/YJUdEkf3/gGmL64HKh2RmekniR1ao
Onin/3SO8XVwWbDIy8m8Z3fp6goTJPQD7uOjzX/GW5HNv+3eT0QnFaKPt3xJ7io8
ZVRJMB0Zue5YRD0ZX68tyDaj1VlM6IKDNlLQqVcHSZwEtGSofbBYUEYMruSe9eNc
t4penc7HD5L7XhHGMJsUEdf25u1dCL7JVECdKL/JsWcxT34lNbaI9bk6KcqlNUxR
kx6q7tFiVuIsPi78yekAc0mZk9vjMW7jimJyGdvNiFRuCAZJZXYO6x62iY8RP0qD
XXFwqKZTD9rjAVRy9zQV2fer00aWRcc7X+5Mx71ofUkcLdhrGraPqb9R741YYHld
zsRMmJIVDPkzyK+LKgz2sE3wqf8uKIfLfGAPJa4pGoLChUaargTeEy7JTNKUVqCD
ysKs3O9rR/M4xXPgSmJd0xqz9GF38781gRVA+ARCtD8pZWzi8kt9PaReJuV+taXu
QF2Bnee175O5tUARV7ayXxYT5neArrLezZyBa3g0ZNVDuUykTGIlwhtql4ZPXIfg
lEraIYzjUvvNv1dg3tSRGeggzy8q7MbKXfy5NoRdZAP9XzQrnQnO/yccvz45HuOh
sy8bzHAA7Ci+NdCRrGa+H9gB8CavA85cQiQjxRwobsFk589VhR0J3KHCfIQ41hpC
idDKHd5rbpx9A2HL98JQhNLTZ2T6y9JJBFqve4WgPxsBw3X+UwWd+AKsSG+DDBy5
+l3P0vWxcdiV63dxCe9MLL09jRG2kDok7hs0K5Nu+CiLl5CVUpFicbZcnkyhEmL0
d3knEnheRQI09jmZ4TbBA983uSNsML7frW+gLkGmtas2aSlzuv9fShThXWktva7U
neejvsp4OFiugjfJ2PkAA9MNsEF1iVx3lTBdZB5nLqpqM1IsGIiMmTLttbtzBA3q
TI7dzXwJnyOS2pcIpYI6Kub3/Y+P+5JnlPyFK1B0sknAC75igHnnwWHxki+213cR
StC1x1LavzFdjO7aXVecmWLqtLs1GrcvwUaWD83FzJIrZeWFpMz8hyFteAuLTJaR
ERMJHyjCoBFrHVgre/BuyZ/4iEhsUclyHnEi4fo6PIE7Y1NiNdme7N9ETklVuTA0
j8DJcLbn3Qrwtxok1Lj5G7Bq2ztUXDN0xAPyqogbQ7ohzoKDDEwOUYN17b6eV+rj
HTZZ3o/iabs15h1CmtOWa8yA3WSnMsqXNnvISYiVhjylqfd19ejWUh8sHUTfu9s0
AZOPLeQDMdChREmy/VxPuD545dQmppIXKtpYWEFAfvIQkaemGHfyngOM88h+qdLF
us2VX4ps6jEEPN+HBUAVeg9LfWdGckLnUwjpMdqvd5fVHPaMDW9wRWhNzqssIQ7x
xdsUwQYCWIudYr4p/imZ3YVGItzTVPUktLw1DkK8hfhsfqXCXk+ThAunD4LCE+na
9izpZeTE6HfjUwsDYhOb7jtjxD66GY5WlUF+7rGyGa/QWIbrt2q8mNeSE3/p0Uuw
JxClj/Ohr37K11Ug8ppnQT3/cNz3dr0m5tWMyUbptIjHjLZd0nxTX7fpiezoBTYm
iEjJqjio4qQwWUoZXeRwOlrU5pflJ5EOmGoVDgxlRt0gbKVqQNZDxTHyU7JJBQ5Z
ZmOwzpEPUpGtTEnEPUHGMj4rIUAKdP/INtDNzuY2VKuP3niRJRza/n1il4HQYKPz
3B9w5iV5M30dLGXjekNzveaUm+4SdhImg7WL+u71dm3/94rI46l60ACRSGp414nm
aQ3cahF5T1fGkDbGJRCrSMW/DVYbsrFiYtuKjLid5RFMAXFpt2q1feOVtgv1ZEBK
/aXqSPiY+UvByj3Knlb/nU09M2Ilj868cFwsQiUGKfocO+O7VHAK87FOKjr59kgj
wVeZRQgj7k4+gUu3v28fvJ9UROODvO2s1QaUsz/G39uJgH9inBwCSFuPCiJ5/JHD
5SPWykJo/7QTVdwVDySeRZDau/EfQ7z1GIGjSeoQC/SFp739CdcKxryIdN6dwG/M
N4xBz9cffuVk+o6ia9kjxAE17jayl477om4EQBt75eXBEcxOtS3LlSJyK9CNL1Or
G1AXVncwp1Tm06SHnQcTelGezxzfPBWCC7JkUd/Rg7TM5O9woB/qEJZf1ADwzXQv
JV5+/tX49ejNc4PW8tckP608jx6tbWkpUXLI16qEUSLustDQRq2BhalqT62XFZax
xnNM+gZnhq1IX1Jwkca69KnJUYdcJ3FKG782ojFe6YW6gURNIfmz0kUKhFofOPrW
ElNiqJJbW9P/Nk1u7h/8D3Ghfgjx0LY3wmIvkxxdqeqHNI2jOR5n9vFusGuMlLWJ
Qo9coOa4VCjqwb1aXzSrZG1eQAFhbozNwSsesQLh1UoxOJLW6cLDyLrfcyIH99xx
K5qOFnrUZiooPz54h7wsL5uJsiRgq6tkE6B4yyxy8B+ItkKlK1qJ51UXSfnxblZc
Yma0AdijIEGm1J6+7ibQD8EJGd11eHuqKes7osaQgsVgE8qkZe4ML4/Ut5qbZFhh
rOnb118oPKQdx70BRJYsOMT55ivQJ1qZHRPCvrtrvyIHohnOAX7oWTLRspTFjSj6
BgSuRW/8rIyhFX4jg6ki+qQXls64f6AqjG/xRgThijEOQebUfa8YNEp0Ga7E/Ntg
hUertVC5yJnxJukAKdH8aG2z3Lw+TAi4VdEBR9KMcVQmFgNxfLXVQJSyMGCyz+Vj
xHikhFRMkH+I5OSyr91BaqZaw0KAZmNZmAZZrewbKX37uBtKgviKhtJDhhr2LE3y
KinnUoSREJ3n/DV6f3/4i8fq3GHxbNIAswo7EQK0kpPJqtRX3sRgQF09yE1tLQKz
y1rspOMrZtJnyUmXI7DqPhBusdU3tGuQUemjpMb+36tkhtinHnsvQswSZ9U8EEfW
7LlnUKP8V8wuWJ4OBYGeO59dMS4DejmpqLjgdfrIBP2alT/Fufh8z3JYzfnca/vm
JjpWYndX1EZsBZAJ4FYT2TykUNCmPPJ7wwdRY842BCP0172ebcQaEHRJUC2OFBpQ
fYBnRHKgVSt9749hMgBPrku03wFH9LqAhmTIKUVO/0lhtJg7OSU1dVmhKT3wE2Os
up2hHcJvcX5oTTXXz1tDxbSV81SKZgDvgWFGGhawrU3iPWnnUWre/hfADlOwD9d+
BZWaO0fsU8B2d6rZIFTD5oqfw8toa9G3DuaZk4vhnMLLwTacf1NPoayD3/32QOSQ
x5P7XPW32FTe+ZRdgyfeYhQuI0FFc/JRKqMc+NUWMQkcs3Ei+0CDtlfLNt8CnUiK
zz9gTmENjaQklkO0hdPDzG7LAFj54g0vWOktmvu7CcgkXmGHEca/FINeaMWepdMm
XMluzdkMVsRkTZ6k4RKTKZuPDh+GaXEsIzHvLWAwn2y60ERjaj/MvA7om0YZfpwP
1AEcJ/EV/VprsofbGW3xeiG+10zO9L4hi9EucNdYK4/G9BDRp1xZp4enB2p9EG0p
e5eBql0/BhQQ8kza7S68+Z6G2q5Mqo/uPF93T3f670xJW2sj8M+HResmATMbMBPT
dwT6+8+igViD/u+5LsFCbZiPUnDUvXNvvGcC6Kag7nI2uJv9hkOiwGKEdMWnpYs0
CqDlsKaSOQWvc/mresvqNu6QBtZ0pp9dwO1m/laQiOThFvtMLtHF4flMSF2p3e9q
mQ/ewexE3T7evmyPIQgNV/eq/KFk8Cgt1oQJBY4q/KcGco0PYQAAdjpnENGKhfN2
/m2CL6w0rEMLm1g5YZmLR4DjlRNEVGKw1KHVxRKzAA0u5YKu0pdlDvKvd58RFLkv
OYI1haPPhpi7HtEGeRPb+Z2Ui8jwiCTHAlAgm2tbvCxLTP/LT8Xklfcpb/6YpOmh
B+pDeCK5UMKZKIBexhIfFeAhvmmXac5e7YegFCDcQibTCgCcg6zXFF3grGntBzlk
pTHi9CDG1jqu1/8l+ht9UgdEUJou8s5tPkN6Nl5jIEMkK3HjOQdgzW33eqAhrZJ9
WqEU0sbJ/k6CdQeA00S985TQE7YFHDFK8EWiP2g4EwOKMlne6JMo07/nXgA9z6fB
JwdLevopw5k6YQh+6sU2fBpZwo40DmsZXr2E6S/LyOo0O8UTM61A3hZuWc6HtJtV
6YQF+cLu0oPWDZjQTr+84n2UUfyKDqktII1GV2mgllLcTz/DvQMnjKsNFrczbhgs
+uQd+u3aeX6kl2MZpIXAdvoFkEtuOIYfjH3J6cVV8KJk8n7I3Dq/neQCuwx05CFr
1bD6W4wJWSXI3YEDxGlkuAxijq0tiojxAn3u32cY45yb0rdei4mK/b6D94xkexmu
cHIMI/ishrPl+towORQaWaziLCUR9jymnZl/G6f4CuT4zgNB29gKphuJlUg/5oPR
5q70LBJlTiFh6chPMmF18dKIWZ1ru1PBQpGlzAk5S/7LHZ9H78LkkfFdLApKjQJ/
sTVfOcQxr8K23EYrfBadZaQmw6cgEaqgm9vCZWzMdMDRPMUAohhZMIeIMn7HpaxR
LgQU2hao8ahnJF0snEC4wI3Oy301/8lJjqxgh45DvmB/imcDM66dekK/nkBee/xf
/VDCLmySpbZ8UNdxLppcXevsIcGY5ZQhdOEFOFaegjl3zNKhXDMg9+bZSwhjRkZ0
s0x9REn0x7zEGpVA7t7D6HbGEgfrOVbganOc7OMvLjD/dtjOLm7yxkiTsxtkhVyO
/jZXHglJR2yaPqDpvjXyUR5L2+OKEjitjq+bW6DWWkP3BPYl0MqHBrTM7/F/7hmP
ZTFPSGvEy6ADPKOTzLnIN6N/jpga9+ndhjgUuLS/31fFYF80qmkEbQ1Ud0eDgPc1
CMFh+fYSaCwieQuqxF5MQvmf7AsaPK5A3147vAdduTmbrEc1U9f1mZaLWyLXpUDB
j8JkTMN+A4kiwiIWdk77JPSK+vDV4cB6QZ/9cW/8PMHTUXdI2c6i3LG60tKui+B8
+bMXop97lLxt/p749X6NvOUp+jA1EJ3qHrYbAbo3tqSJiPPQhdiGBQPiSJRcjdDe
xPF6GXxSs/fxIJmPmyeN1bQ4PXrCCO7fleUfsQOApHUXV9IYXpwsBs02HdSeWTx4
D591m9AXbr+tHtqFWkqQYvAjY8D5uLYbVOcw1+lVqrFtSSnIStCK+BcWvOVtKf8R
dbUH5QaQUHsHDSLx5lg/Scng4lruUkJm9z4sEMA893Ub2JNKoCEwbok/T+9t1PK+
r6abBC7xUC1WLvSWvCA4rhHbBBkRlvzqAF1ABJtmtQSpw6BlF6NA7FGcYwv1N+Zr
ofxWLqJtMEb3bB+oWUz7kNSx+WrjOALGy6SmEz1xM7tHZCpODn+vZQZLANoJDerI
JbEVE7SXloks2W4mU3CSYXDsPAykE1mVwqJuaoxa0O3vQYfB/Ege9b1ATEGQMxwy
cIGSZieaC3SdjJsXut0KU07BWfGQgvltSAKp3SbztyHKfYKE4M22tEueZBqg1M4f
m+IzWEDNGn6Nqiv2JhecsxOf+b1ZBO8CWuDcB0uczEpx0lfK3C1NzfYPGnF/Dspf
7D+TZlQF9otbR0CHJTl4+NnrKluYojUolqX2csy0g+fQLsMmvKZU+o31E8kHeb/5
CQmOTYtuGrN3vB8OJo5z4C18BAGmmMeFznOA2Txf7Kt6xTeL0U4NZK88TW6H5cdP
Ju43rekzTnFtRnzoy2pShiguNzDSpMvVcCpFbjv9tJhk5uxmJ6errqKRqrVmXmkk
6h5uxatXsN0JkakUFTz0DKn1o64sNcNEcN3roRmxxIEkzmGq2191oM2odWU26r5P
dsfRPrSZfnkkmb9/SEBOqWLk7F5qmTqmdfJTNU9dao0C0IvJAoKCUjhp/Q9INP+j
tTJIyCiazcseOD/WpAvztr7tGteunyGSaiCglg6KfrQQCWuwpxCSZDDn8sXsxOY3
KPcenF5wII65/QxLEHT7TxSvunbM76TSdOQ9nogvmR6BMnQU75SI57AN5VfV2LmE
4/Sz5k6PCsEr+66fWq5gtoPZAbUlv+KoobeOVpn+TjRc5aDvmhJos41UXz/CeVGG
ZDonI0qkpcGUecAR1uXiOF56gJqHggwA/xmNGz5Ga4fdX9TkLG4sp/ANlHT+/W0P
OJSlPybmok5A968UGgrR5wW76RTnJJFumS254XqyPyzwmYSEus4c5ki9bTZ/VqgU
hhuboU8WvKweCDvRdMD7tMgPH9woausiIwoHakHwLx2xho0rYsB1GkMib+5ND7gN
hs/VE8EclUsUie/h1gOG1LK+btpvDS6VFYQZt6a02jo9IyhnGRHHqZGL/ouHETdu
NeyGYVe/uJQNbHI6Zs7+FxC7Chgyc69nCJgSmhQkkLmPuoqYzs407KXwxnBEzjKm
NnoXsu8nK9tQzZ8Kl3uzfnW8LWK0b/8oi2aaK6wPvDZ30iDQ+8yNXaBHlWqNxNNe
IaowIfffkHzjQaYSK4G7Um2Wdf85gfx50FswngFzJd9xaP3cIH5Eme3LOZO5/glZ
xKhchJiyh55UAe4uOUpwTi43e+aBHIVhxvmdLh8fTywjb8QVVUX3IXrvDMVYylOG
1nRsB9mLmJ7AeaUMsSdK5AY2r0KORGphGwlDbJ4b2WuSsv63JcqvDOkHVmwaMyLJ
pDSMqkNNiYm1Lqit0C73jBLlP3T+6woXSUktPWd8MuJhciR7Nk6o+3mOmXSPTxWL
8qUwSfZOy4reFyV0TACGXyDf4/K7W9uJI5RI28UvTreh+glNQuVj9UL2PCWuJ0QT
jb8xC5wsN2lrpg8BIQnLBJTfrlWk210ileXwA2vP03XVKrOLDaHhKbG/jN4zWy1J
PKYUASOPKV1fNSw0kRjYbWSNG3UpU2pe/dQrRE0/8nZwk2nVnb3LjbwbbdWbW8s8
76fs44merHEB8ch8WJmSoa4E5y1Kg8OOmT46Vh8wbWI05vx3yu/rpxi/IKy/MiIS
Xs6ZpvcClTHYlhlOTxUTL5oxuTH5agZsvs0NwSx86I/VIoxg0i23/sHpirBL6uZs
vEvSA5EbS2yFDVGXjidErYsZ0U0xW1LX+aQu+eSLhfIQSmeUwtK8HYI4cy/FY0ce
YoJIBllLk75CtURk/7VwOuDpq0YXYCBb2Z/ctxTfdR8OnhEy3ji8sTL4JWShqM5I
Sa4hRl4VjKjIvdGUrg/IwiYHpR1K4KcS0P1MmMWotKMOzhq6SjRyLJ5t8okHmKIl
HGnEVxWXwK1ZTQxpYVBVk8QaVyHwV6yMAgeY0psWYtzieEfEatRwdGg0UdZapp6D
jwfw55KwpgMawgR+ADDAiszrklHyUqf5IjcsxNHQ46ibDzJswpxVBMkY76c285fQ
CHCndFrjFT0sleROzA9e+cygGcaUMiMjr8qbXJOa3nZo6oSdWECua38n00eLRXdF
7DLAzMKcO9PsWGE3Da9YyVqmUWTEAF8G8s/8WacV0jtFHCisflnl9Ta5DrldQ95x
FV5U6xz/SFHfojYPF5Antgp3kUhD0sVbMtFf6b8wo99kKPQTzGF+5Vi/t+nynnL2
Gq1qY8iofNTsWc1lQ4Vp/gqK32b+Lg6I18uH913Qb23FHqHGj1XYZv/nAI8vmJYv
51hn0m2IR/Dc+5ZYNrcxHwsbouSXtZGmVH8oox02bvHduFc1ary0IG0KUeWH3cOT
28lrK3/hG7GJ9coa+gLZtTJZfIRNniyhQwuIXL1CvImfyU0f9xP9jYhPmsX499tG
82A4HDoxSlG0hMbXbP6KXeIGt9mLZZoRiOU+8+EzFabAHJFhuqMUQH+g51/JnXnG
VNvZP/scivxpUEQgVK2qrtI/U4h1pMdb6XQ2ZVT2AMS+85opUXGOfnU24qLM3OQy
4dsoJqVfaoqXOM6B6TdjP4EOFeZ4qoGamLlO77XoNS58fpmU8XtRDgdjk/9HZcOY
9uoyCMDp2tNzcvhVPzf598PM+96jwnLPOCC/Ip1IpYQeaKQIwRbdPT6PSFWjh9Lw
VBdpfc5P+UmjfPUexd5BgX2ce0AU6YkMJ9HTvnel5xbRPpFcFVwWGdGH+LIMkc7x
m933EM8F/3WZYXuKb1wVA5usGW1epuGv59PKOz95X3vTuvnhfyx7m1Rjnc5u7SPg
vYZozfKmdv5bvMB88RtuGFh3LhZcfH5MX7jTuo8CFDxx6OCD3hDs8Ud61rm09pA3
qvQNX5C+ztOTJ+AuKJFJ21JLVMkm1E7rSWNhsLubjJ4d8gnfy63p453EdD2XJv4I
l26iaxeZXO1CJXMPc+TMj8zpWYQ/KDLIM4DJ3bkNQHJONBOv2xxxFSvvJ0YusUez
7pf5AWE4MHPB5z9FJQwjQPudTIrqpAxJ62MzClcmFmfusZIlNDUTg1BI6E4E4VXr
+ERUSJXkaY2bkDfxv0p0evAhSL7/zYcAjoR585djQyHVJqc3YQyby7zpjRNtJfoW
lBW4HZzq4aSI3x0KnVvtOtHnzu7nnYvdRe6iU/bGO90frTfJbu1ZjN+B4I2KpSnC
Y7vl9KFNNZNa+fDazKThYXlcTtS9g2geMGHlWed/v+kdz/S7L9GiKN2F1Kwg7z5q
v1qttei5VG9KayXnR9QkDOB8fxwuvw60V0UIjDYo4B30yTelNFeyTKMlMzKEy86X
rqzPRNw5zQmhwTKIWOpxCSkbrc/2iU+wQfh2dS3VKzIAqRmdWn2R5xkh4X+jFpQc
LtVqBAeIObpW4FgfU48sh4nMn7KS46NptiHFYxwqj9kckRZvwvZrjvb1MgUwCYI9
dc9GZsnhHJ/XDtHnzQw7N/4Lqs+TevIJ2XvQHG0eDKRMOLge4Tt4XkAm+2j5r8S5
stayVCulDewXWMll1AB7UstHu/bcMi/0d+WbL5N2/0uuE5k8Kl/LNLeUzG1vFKUo
ZqL/6IyLj2IljOwGYwtgyhJzVzf2bb+ru4PVHIV19V0nyEX3zDKf2ywjdiWtdyMx
hPCrweSR+ErIg1CK7WlUo5BA00T3W9LUZBtrtRbuDRsz2BdOsUskdvSkSqF3kL0d
zRai2iiuES32Ypb6FIzsHAJyXBmcXbYeN5nD2XQjjmIUhMQm7QLGOA7l1TxrusmE
faGN7aTXCIkGsE0XGxSEqeWMOLcXNAxsHM787DZD5gmP46VN5o3vvijCqGV8y0RP
s01enOQ7CVgPa/p9D5jFJqLC0IudKYmo9lB4AtqxM2UP2RrI6fbAgullKJB0oide
qfiDSQ0fXVqmqvdyUIYPuE6Tr5gtgpeM8CHh8Mca0WjG3lcxw0MwKeVh9yNsT77E
XzfkzRmlZ95X8y/QV/3vxf4MSw4OgkIp1lrY+Eysw//AEsBAV2gJ+WzSX0ntCacm
fICkp1a9Vnmq9RSBypqSTnzsMRLavsWV/Mx3YgwYvcs2aHKL8hyuuAfwnhFsn7+0
oyrGAg+uXps8yjsj/C/lFPr1ong9m4muN0IWEAEdbIT+3hRuyM9xSYTAeZMTLDys
2tmaLsqKF9zZf9AIUQaV9sq0MZAGdpX+8mDXSb5y3i4H25m+/kSPw20vY2IMmM5p
Q7pxEwXYeEMba2q5SXll96o9FagxFAwFcG9Ftwywp1tPrJGyTTX1ctBZg/KVoXOQ
prcG08ihEPlBQDGv2S4aGA1Nk6jhzja2WaYwvc2yI8JDaHotz0O1X/HgH2O62kjQ
zSJAWk8VJNKzsso4uyTtt1tIXzTw8iq6CVuKxice7IiCD5vtSzjfZ/rbxnuLNDCV
g6znFHH3L1kpgDdztQ3RvZeZSvjtCyjoWU5PoUFyAXVtjMRSiNJ8PKqEgZPXlDU+
4la7Pt92hq9wF96Qu2hZVfqYQ5DZ+dfnHIPzuYTeAe06iJFmlXbgPRndrJsbG15H
VoOdm4aWhEQZes5/tDCqSZsTDyjTMnutECgoRamPQNgm4nnkxtEMxqHvnGjIlhy+
R8Tdm/NIbPUzVPRMmt478FOINT9qucoJfZ3c5PyJRGZrxoktYVvo1ArRClgo+epB
aWoyfeZYiB/sEoJmt0ODjxwKYl16XFeOUQWzP1s1p7XAdcUgqF1zXw38wfheDi7D
3j7kK+tVgeFxrh9NQ53QbZnl1ZY8FtTAT9KaU0iOz/RHGgt7TsQTb1492fT28JMM
Q/lZBqyDI1hcDqMJ4WfDXTEpRoU0ifOtECDb2zFx0BskeQh5kKKMNClOG/CLpQPO
VoZ/gTBDZwRGMC8eE4LsLJsrO7P4EI5BzPc8PCK+XRORkUekwufB+KBjngMwZ+3S
JdggpcFHKoCi54Udph3oTHisi1XXVq40R/HvCEKMXwG+8zuYrDDnTJhEoENyvQho
1/Lxy5GoHyjvFlJw4fEXcB0IbbWkHn1IFt4UxvxHr1NHSOVmQr+1KPZ2beefoXvf
D91GXdNrl80GqVIRXPvsVMI905doQp1+4bL0Z7YG++uPy4P3msugTa1f0oYED+4W
UIyoltMFdz2aqyKSs2jhQbcRwOx6aOnyfBQWZkUGlLx/ccPPu2r25+1jlhcUkASG
Rp5R5FwOK5bIKr/1zoWQz361WHI72Aez79dH1PHg++ftEBuH/46CpIa8WvO4Cn8t
nkOIzVohPb7Uw85tDr5EAQAgkt78Z4eXLl9bei4E4tjE85kcx6L859VRj8BRojZv
IBGJVchGXlit7ll91qRWG5uzttsWXY0Gjwozm0CyH3YqlsU4mjHx6nrgh0O6iFoK
m8PgZeT74rm4/9KqgucEDgLNJHJUJQOnL7EdlCEGB8PiPK4PohGk6a3XOi4eIsNA
pzbL3kIVXFzwFTlczmOc2SYZIJZt6npUXpT0lHnat8T3xlzCg6uuvtBtkB8P5T9O
Y/ko8FWrs1vyGNYNcXekza19vvhheDH+j5VNVuWKrrs06qZUm6TDogamPMvOu2NU
ZQyQYutfk79p4mqf9/CxPcQUXs2f848SqCQXyiZxLoNhe0kc3xt1ji4Kb92N2nIq
x6w8zYDPjutw9mt3nNR9r3doQ9sSGkVMI2h+/U1FwNWDFd/r39mLOizRE9dYii6e
64dtToyRWhLb2HyreTQrHKVB9t8grLq2obm7FV/JXn7lhCV7+S06a0axijPAnrC9
OM5w5m0y8Q9h6KdphxqWdttlVJm6TgybRM+PZmc0UKX39E4FMYUIJWIVfw88Nhgp
WmRYKWXqvCxmkcKRgMobwja3xgnCsob5hHP9YjvtusFlC/VhgTTbZ/mURDpXcUf8
zpULYihga4tv45UBTwjyx5kVIgOUufbTaGqzGZCKlyj0JvMYkyw228Yr15pRvulk
nubU313wM6BaNNiOy5sMt1jwy3YOwmgPhTtRJ0zFRgm4TSIdJzZoblN/WeNJB23l
mlO1bRnHNcAULQZFrENgPzu+d0NlczYTUZ0HVjQgDWFCn5Cg08sP8UIGZnMrTZ5U
/BrfkIoc8FTcLJtZv8ODzKros0txsXVRtrtoVNwenu9PpBkIIjulSNwfnWPDkWrn
CWweMfFclV4038YSdzuoPmsEAyNmrdwjKnIeJ5NkMBIkNDOXdv3IDtbidlq7JZxt
0of3l0SEA8bTl/blpphxC+pmpydf+oMgtdDw/b8SKHswZeLu+PbxpKGYDIFCHtiK
2hZRHocVD6ezZzzXqcxdMhhdmt635W/PCeQGgCKrWBfgb0MkO1QzAuBxh4nwfJLj
WjjAGqno01BfgfTtaVZ1cyh+DIMZzmJZnkWZRZAeA9PRO/jf/jGxRo4IZSDEeqJl
w6OE5BVzrZ79mvUFmuWnmlQrysGS+gC1H+hr6Skd2EQvSXG5FHusrQ50EpOclGSp
oxpnd57foCInWzJbeXOdlyuGdzCEIbIh7M4n94cuuZrgwuUbvMMX2R9+hjmPzgI2
xq/gtpqHCMNhejzxbMLVy5pHiZa9sicTKKmTOUhGshY+8NDrXtBSAtxjgtzA72yP
B8R+5c4mbvftDK/mDz6Ne3mSidnf7HAVmv0WDbMbcZ1nlBqsGm0SgHsipexLtqB9
Viv9flGKATGUNXsp6EYNUOE82i0S6wWD+v2EqBw26wwfLa+wGRvOJIGg+K4JAt04
XWzIq2jzobS8h0o5k/YYjBeFk8MhH3vZ2vmaJ1oBIMnnJ32CwOyU+HT2NtuiA74O
UxYUW/G7MmkigfB7ld8HRYqxjs4Wj5hOXdpbXWgiq3ketN48PkHaVNdMPrVScHtJ
epUVivQeZQunZCcMkfVY5wj8A7+kcCa309paFrlw4y4XsaTvEXk8bcDIjtVFD4Y3
MA/RpTfDCMRaYGwZNHj8MZNk8fa8AkyvSqyylrt586krxdELUE4AOqgyiFCmLzI9
h1vbVNgAaWt1lnWVeF2Gb4dR4Krb9D0Xfd46ef07Dlfd3WJibZVen9eiW3W8o1gk
LZr56fQlR++kbaXlc+Z8IteWMsM5uG7ffjmLBcpOizhRlHLm/tKZIr85EyJ2I821
20hBiQzjeFZMc76XbsUL8mrTRyh8fK3zZmDWY9k+SO07qPk7rqgzdLj/3rcNevdI
vQ5E2xwTS0ADcz1D6y6T81HwWBClp8sXAck/LERNy7FGGbbqgFAIP9cEvrhEW1gG
2Pq4wau98PCFMnqFDY84rLF4wgWVSHimPs0CKwG704GUMK5y+qJDmSQr9YKbzpG5
5VkEAqEtpHfDAlYhfdN6ZttK/jZRoc/ejzLIO7lLz9Y4DQOTzE94nNgmzZ1twX4c
e/wnVMfAGZyOspour39QJsy/8AByn+2s3JXtrYZjMsHjvFJZd2YGxihOxug+n9J9
ejVKGDFe6hCGxOBW2nh3FaOLNKbxaNLdzgeQSY+nJg+Psavo1fESZlYAXgFS/GSv
HFDYIWZQtOa2O0ybN8v9pgItlybIIo7px1sci6od0yRxqV23e+aazYnsEVgUnx+p
l/UhgMTyeKP893Yum/sH7qATCQAacVmyBLUbwELHM+zOwNw49LCoXrxZlh251rBl
2brywPSoliBfeq7qBHpFylWJ0xFbs/uF9lq7FlLho0ZVaJy5p8TAhhxVLRmTpHJW
ZHsqLdj4q/EfAFWri4bzQ02364iJYEmlmfTirTzcqynK+ZpIYxbVpb2Nsc09FK/B
s4GcgpLN5X1RgsYtnNd2TOyFXLJj/uy8pi9V71MlhacAfjtAqlG4SG7MRVoAEmJa
McmNftRvGwxS4LHi5lZZ/izycnpzJL8hBpK8DSmibwhoK7NOvefo8HA/RPWHBMKr
MtlRfdv/nAAZSlB/aTRspG4IWRkqo6MEtDaQIvwLxid9HW+wUBdY2I63RDXbM6js
jQAg/J4vMrhiCSgQ92vMTEkg2qJqMTS/73TgcKFJie0Oxd15UGaXbsxGBQbIHDee
7TNP8Es1OhQcLCgclr8Dimi0gXOe+4X62RT+t4pLo7uUVhLwO5chM79XpLqN/Oth
46iToq4ffSTy1mBidcBQPaH6oFJ/IRb8u7xtF86fe/lJ937fSFZuznr8Dk3lyc6g
mSKBzcqeLRNGNiESFKZVBmzPz//zOJhESldSbb0wwbdrINrrdJVpyFU82fmZS/Ge
wirITxT5Autb+F3730TA5UfkMU6gyGrvciPh3SvvDIJlXxMKWTB1kKPjvobPp3TM
aU8QohdmIxPVtKuX4ifT65ig95J1rA23PN1Ytg1aNYzbxYcAR8ab8c99zKWjod7L
B6O7TcgZOaA4VMiWiMpeIGf38M7NCY0xspXkAglj6B0bVaM6dsSs8SAVhCnvSNGv
RYG0F97KIJ7tofTIPj8Yz7cW9uuKMS8fO4zXdyYUbxcMqmhpM+X8H6RBU5+Xb/hn
2rhCJDQEIP7bU1QsN1bhy/JzTzfMpPf0RIun33P6IsRAV/iUtqtO/IyfmDQ6KDmu
rNu4AeY7FKe+3hc1aUaOLiAOs3tuIimeSaKQOyKpK59vGOjU4qfGd5K6Gd6U1tyV
y3dGTnHq6FCVqfNKTGemZ91xa8VpxZ0Ra/HdJ9I0Z6pUEPpFxRwhaMMkQUBRbDsp
eGqun8SYOUbgMEp5eYyanuUI86qp0PpIyx3XWYOqUwPDhata+610Idtlw3pE7G2V
NgJxnjPGE/F5jI5ayJCa4VttX+wCJjeq22C/AQoA9vpuobbbxGPVNdL5gPdcUiVD
zYQtc0YHUEFtCzNwNoZJfwHkc+JZyfvnZjyg+dDHipW5jAkSZUt7K8aaR0wd0UYf
xR8JAiNKdoEaYbAGsnXWiLIf5Q5SBdrr+Nos1cxU513hbRT8w/DLyBzdqZCzW/RW
39memIgqfM6mNh/jtK1CKYmMZcCfkve5yisTX+x63PNASf+Bb9MdI6ARtYBZirZL
oKLouaKvFYQXcL8nKQXNYgjXZz3l9K4Gq9A2hHUWj9R9iQwQykgVB/NSxBJwcio8
M1z2lx5v6SYcpGB6eKL9q3Sp8GR5kKQq1Oanor2MgZoURKvgjNyYg6YH/o6B6FXq
tcinp5t2Yae48qDlU5Sr8GJmEy+MhKefZnUpW2Byh1Sq0k9kArK9501OQMhw7htU
u1ijZPeyjfUPOhvp4wrugGW73l1ngIWvxGIyoQuPpw9HLBWJWlJ9A0AxYsbX+hAz
6r0/x1ZsCmiNGIiwrskLMH1xP6G/6rzX8kcm8UkoojBv1Dfrd3akzRKc/iClqWqK
B90/6OmYO8RdCb6eRuurNcDX7JwkxgwihOndXmQR3xJqdjwg43K5aOnkIdvPe0mL
MOj3gGE7+c1AEVcvg3lZEuhiuUDZ3lh/n1Xo0iUVlxx4DbTf8SiHay+xTVW59CvW
DuqdrcOsxEfdC8x64h/kiBMPFghbsf7D/uohc562fAnCPlStHe2Z1CZ9WHSV/e4p
+65p8YIDSguKGcRc4naNmaiAkGbS+q2Xipl9hETr00MoJGNTxIhHomZnOmMIUE2Q
sDYIG4djCosTiAqfEcK1vTCSn9tmzj62Z8av4YqUbu3tbK+lnFW5ZcBxn0vAO6cd
gduPHOkapbPWWLMScTZ2SpIsLWnDMYyeQMmT9YE21nbs6rY4kvMTHOciRm2z2DkK
0F/usw/WFMEE+m5sFdopz4SJZoJQ2BV8IDSU5BdEtnuBoWWAKxrBgOQ1C5MRyajV
qGIe3x+9julcIfUrlVBmLGl0hq5cavssfvpikCNmdodrT0LLj3h7u5lWnj0ShwiC
9f0+7KeUBUrJZvt0rn6xg/K+mUR8Aupxm0E+ZjHNk1fd0c4wUfhb8RA3zVwlMqJk
meiiAhborgHlKc8OQo/OGq25C11vdde+odcg5wGmnUcP2sONs3GN9baPHOmro4a+
LNb9rnT577xPFd9oaPE+wvBsiUEgfpIHmMIPGn50K/dHmF9MBsnu1l/YBx71w1mQ
9QIncg/lllw1+c8+pAgYRPWXpDqDvGUWRl6dslI3icarAP93vdyIWCrTyCgOVYgG
B0Na6Tkib+UKrqbs0A7qXxFZK0HfgjS55qNYveQ9s9zjORny+d4Yl2qJkDn9fXuK
NPe4qsY59i9Vt+e+M4slpl8WpdmqAQsZwvlN59o4ZCE1MsbrnDf2QUfhgFGu+636
qb69HPIsLZ1N5uu/vPqbudKn+7vHOjoa3jByWwBAhzUQXmW2V6dhCAQsTGPz9rgE
F12l/73cu95UjAwFE7DAiSL66UlE2olDlCy3Z7Wuzxi4+SV+WYPnBEoRoQZlz/6P
847mn/kXBzpWv1XMjYvF9C8muTZ0pEa/zeKPaiZwUL2HiM4gvtRzfSc9PKsdSf0K
CVVXDZINANPBH2h4AfAyRxto23yDpKS+GiiGy+W408trBSPFgx2ZLlfuvzgHhPjS
89zNO/74TTHRtc7PCid8V9tn7E3Z160dEVoLnQNFD5YiZcEjH/IAdzBfpJoUzs/5
vzOdKLykIsq4y40Mm+tuoE4CVaYVznEmvyWv/6vbOcDDxBh0Q/2yeu7UfxKT4UBq
eRON6E52WlGSl1TCzQ/8v4y2+8JsC2lm0ZlfzsWPmwCVDJxbTwynOULdFp08v2o1
icobrW6/gJIE1mtd1dfes8eSq4lwfrTUCo59GXbyjjNdTWyAKvFsHxifuaJ2gUbe
B39Qiq/esFvJsu9pIuq0N3VvI8Ziv5ALj+d5bYV8GGOZeBnKNYhnMSy3QQ8kKHOw
FdAlqerBlNPyvIqfdvx+NzgI0OXhgjaKpdszmTpc+V6V8W5h++6j/LlAIvrbZGWX
Zdjd6TTSeJv/WzhPlydc7suMxjW7d6fLEI6SQmHswNbyz8LBi/Tka9SOmRrV0jEz
f9cvtDyXlcfxasUtkr5F6VXiSd9PC/g1eWZdorLe3NFgGVGj46zcErWm4wgxa9N6
rHl3Cl4yV6Cu6YvziSsuT5Qv60UavtGIHxrcDWxd9z5WlvRg0AT5qgtBFxzmHkv3
NBozw/UEMxaJS70nxl5cR0TW4uoLEfE2sXzILZmyPu7Hu+xlUosLbB9G0p5t3QmY
k+62RYmpuWpILgR5ypUkYJJQeMoDCcx7f9j8389nK6FtLB/t+Ktgr6FeW9q3wqQI
RWWHNu2TNnxCs43WpsN/f+KH44fHYuPOIbk1awJEtL6i288j5Z1F4J2JheBqF+Iv
tHgkMdEpXx92cE9koCstcRQXuqdmEp7CgJ7zZlhRxkTxw8IjDto25xAHywlWwcXp
ECj0FJ2AUJ5fh0oPmSPJSxsX/SIGV5gylebBnhXweF+cfd2scZk8EnCZaevyIx5e
00oLAOz5queIq68DDydPr9CUOt+isAdgpCjj+sGzv8dqKKxWBh+SO7+uj+VJheMY
wGQhhMEoxHViHjY7oLKJKW65kQVAT76+yg+2sjfTUpqHOuR1Ifgr8lmxMIpBmVhG
QI/vgspvQ3MZZyGquTgu2ZZ7+Y7s0DEAfyig++VE8tpnySRATOiiooPcO/N7eBjw
tHXmbASsU8cdAjnyTiPhMCCKH0X/H+whCwB86VSDu4nYojwaCf98qlT0TP6bDdJz
c/CwA+K1gASyfSdU3iYH6DO1JQfh9MvDQKqPSWBIjr+rRgLPF8LgwvZUsDVhckEW
NEZKbIrNPJJaZzeh7ZxaqTSv1B3TlS1lUh6Ays/6VZVT+Eznk65eUCl/5s29/P7E
qOrQqWyP8gEv5LSV+ORhT87ZpltszjDZ+0BwKa52rC6MZmF/wCzbqLS/3FwgLgBx
lffwXC8U48L5z/K5c/zS6LxvxcwzpQHFtPt+c/xsdnB07xh8BXIwQMAxJfR6OJ3g
cAL8lfIn19Ik2qP3cW+F2Mv4xDCETTX22Ir09Rl7xPAl1rougyKXmz4eX7VGEfLJ
3ZqYgpfP5zWP8xPsrf1q5jn8qskHH+JUrxFYRBk9MQ+OXUu4WQWKchQlYesITVK6
VkStGzyVKH7H6AzHDKuhmUF8aPoLZHvEB7UbK9ok6BTh028iiihQaaOv9GOUr+3Y
ORjzc43G9TMqe5NfGedP3SNfEXsLLKjlGouVWLMQpnoe/2dsBI/SnhHJoKGS+3fH
zxm/HMqBejlCF9x4a4e4/rWfqM+alrPQ0dsWEHvzW6w5PQWro4w+nmB/2SfLULej
vJhD2fgUQq1KacuztOBFC2YkYwg8d0jOE3p1nKNKz8eJfkfbWaaLSAGZHyT1NNEi
OdHq9z/X1SLYsV5qnuOj2XAGRauZZZ/LY42V0QqxN11I/kXx8s8JMUpjgp1pKIXu
OAfzAg7dLO7gVdaBF0LnImlQ0phgyq9wzaFDIv8CnUwTFxrS+EZHANvyMBjhibIv
GVSoaemJ0bMaIiw2BsszH6j+Wwv+pN62T3q6vMUWWalIc5XkoWdVTArG7IAzgCaY
Sw35SVjMqKNpCRLbY8a8ewVyW/qNkLKQbs3CB9WDpwzZ4ajkCUBdxXZqpjlIaGXJ
Kqre4LqmcONbWhIkvj0VefewQBvRbYzVRMhxjXmNCbbMN4H5FbFSiPDqI8qMMAct
k+z7Vs8LOQe0MBoFCzsoAcA5xd1pIqDzXrNSquIpBrkNd4zZURbYPeW7WTmY3bOG
y0WWVExCW5C3QcPxpnn5MO296chAzjBgo3OQ64rci5G+ZbThlfOBNEaBIqQvaUcy
v+lq5Mrt8bQYqa0SHhU8tqZ+6GVX7GINythTQhtvGQ1uLbtj68jbAhO4OhtveWfw
sG2CapCryX50p98D/LG1cuWKz1BXh+fYQZ/dGNs0QQl6yoBm5Fb25iDwMzDj6RL3
8gD08RNszFWByZEo7Ja78E5YlgfnWKyuLLbg593aBGSUCNUYh7hcEtx8XMQjCPbV
d6VTDy1vVeHqeQZiHqKHYntsvdE2LhZyl50rLk91Nr/TZWoA5+augTq07G4qCgNb
tHpDucJF+LaMmYw5FqLoFBZC/1w7bYlZMMKAJMyN2r4wa69isE+c6lNavvjbpNWB
x5vHSawMgTLNYtxOXU9otmh1RqTbuRW8nha8vCrfrxnA2C1LkXu1nUFh4etmASJW
e3uFsa0fXo1/Vc7Le/zBTBAg6Su6aF++WfAmqO+WcXZztcVTEqO3oiLH5KDv3bQp
S3+FE9z39WYDbApcJdD0qe68z6mxffOKubd7S+s2phb0FaQelZ9I3yoLDP0qZK3m
43rL1iO4vED3PxZe5Vnc01WLvX4ycR62w387p39bWgdFv2bBSTEqid/alqksyqY/
XV+65JQIBeCWbEPka0iKyVECTqr8BBFsWIzoKW9du6vi15pGsy+QcV2Ru7OQa5E9
ahdeP75dDuWRKoWMcaa2kiScflLp1+wHsHYQEkr8bHOoWSTaVWYGpjOtqv4Iv5te
WyZXk6WKQ1XAcDmk40boTeBeQC+IWaseabGTA14NWAYoBiTAzcnU3GK7N/qJFgzP
T7iZeCJ+zbawmkCqHD23T8t2Qce1xPqJM+mPae6WyVmtoXI14ZkoL3tJWJT/k6p8
ElqL36jLGcq9q2lmfWcMWqajCs02mQtBF9SxOMo3pZPiUoUyEzpKhnlA/eeR8eJ4
9HCSioRW/mC2s7U1HsJWOaQB9LFKuHM3O4ym4qhIUEgr1Ivm0sXGdOLEL/LbbK4H
dyQkUMW3+TIZQOtYBXLmMLV/V1zmSbSRhk2Hj+Lb6cCeuyQi4URGLZ1sTNpZKdwJ
IcMyzgZ+2Zhi1pS3IvthU+zEmmrRbpbcJqouRETq8yQjFBgTrE1FR0ZoFWTJ1J4p
GphuDIktshqTxuY8pf3ykvCAk9wiOOJdW1zYL6Ai5GulUbyaeBi8pl4d0xH2zBdx
qma0KyyTYsNSiYWi7OhmgD0lTQKwO7EhW2h0mWuQaBlrunGgtmlmM1noqlWWthqv
eBQ4YmDWmEzpWd5r0+oBRcKyUNLyHlG2cuHrb5tUsXBvbvVY0OQ+jVCnsUQKgC29
3n4qwD5Ksog4/1soY+xq98CMHwEsSDWprzZeHXiqaFYk58Ch3jRP4Jn5fxrQvGPb
9DNvZnK+nZsvB7hEAxyNxqwM6O/4I/IhEHT/vqUCHApSC7fLKCfggw0lHxoQ+TQ+
LtBSUciGAyDIu+DX8kFiZmP6dwniAnZLJi09sD6qAFAIOLQcsq3vT78OBgZfD7dn
Fptx9plolqAnbH9g8pAJxAp7E0cMSy3kSQiF8z/GuS3w78W4KTJulf+nBOTrh+eL
vHBAASUyAC2EoYH1zdipeZlRuDG5zXw+y0FH3MY0TOG1hjprmUTMaeAv4MMxf76R
V7ddXB7CRPzidVFduiWgtl5tO3ZO/eMZRraKuNdpmbUZca1Uzt3SIjD2+MILNZdY
O1Wr3LejTSWgF4Gwg7YdAUUCYBmBh5lVpZJAg6AYv98kbyJymKNQBkeN9TqAqOYt
dzlKo+C2F0+ldOyDfHvFTcXTVnfEnW6tBOKIByyjotiYkTtBmG0V99fIWCiwUzXN
frEBKhD6ZVJkpu19Qa7naYeqp8JKjU5DbxwkLL1sFlP0ZjHkOTMvuG/CLDSEuNRC
z6GBKvz4BHg/enRLYq0BcHmFnNeqwlPNHngIPqthA8zVpy5N8Pd7qQ6FY8BSA3vr
I/+FKXqB2IJP3dtTx6tTFBpcoI3Tw8iaMhZtqK0GL68357RmrTZCfB8FGI8eCDQ1
kpUWAQ9Pb+Z2TWGqNeEcpHiC4uNWoThl+sTNDAw3q4ZZ2JvG4g4EFvB42FCWYMx2
IXQ4/VpGXgifOsp6pLrxje88F5Iyb7O4td8haHNzhl3TDdq3TWkJiRcO+FJP8yjB
ohmymzAkj/R0PYoeLl0hxcZSez4m/1n4URKYs6jf+sOfc8Wh8p7IZ+RAMS0x+cmv
0/Uq1Ba3oTTKRfTzl9pRix1Qd95hTs5zJSn4cniUg/qVXorGI5nwlJ5+yu9I250Q
N3sMEIwk+1aeB//ickvCvgHXCs7qfiqrFdxO8RQCR98Lsc57l1wf9v+sBdMhB8++
j2ImYVEyOpuByL76pH+msKNQJGzKAvxXXsz4SsnP41LQ7Ad8lT1LPkrCyPmMlX+E
uFytst1Jl1mOmSjv8rWUL2e5vtKDXzQsqQEmm+8VcranDU73mXhi8Cyi7+a05vUA
ELFbLPzKEXwXuVyHA3CHljSu/Pt0vbAxpZPElV/Kg6byyJmJJtOzYSHJH5eTOC7e
ii+DvAKTh3GSn66C/x0jJeH1WGhrRp8M2WkBvxYCBmTY+0RWWy/uLK83v2CP348/
Z108myRyTqGmI03xAZaddGG0KUPmCpPeRCITnoR9YxGPMcIMObE631F9ooIvxjiS
XUIkciK1K7HiMRkNvcLqYiYxICvUNATkQ0GiVTlr1ypGbLPZ/DHzP9Vatm3KIirS
oCHZ2EJcUZiKWssbLrdXb635Msg1l29fZPx2jPYE9aZSt1gtPaFAsP0Z8y6InGdL
KzZ7iec+u9mCfVVds2+t64cnWSlde1OhCIbVbwNMhfIRXrORrE5+R140IKWqUcCl
ccTnvboSGQ6c24q7mbG+On/wqLEuZfecRzdKKLVgq7bsGZEMDPbh5aC7I03r3sJM
UTsANjTjMKsV6x6DKvd/Gupzq/LgQUR7u1JSsE97BHCeUORBFMPtCPP6g1+pReLh
GNq0ZfqnZI1Q6XjYgxU5X3IBHcsYE1QRVHgzYefXcYPBF0W+PJujHdnPDUZr7l42
3LReTvTaJvzi+OE8pCXU8X3wySeBA7KKQ/cBQsi2h0n3pUDrrsVUye9hWpdTrZZA
hPvhtvqxRT1f7YzXb25VeFXXUITFFQIbQNx4L3bs6Dgd/gGvacuwgV2gI973v4IW
4jsL9aW+F7F/dqqZlbqwlF91rDP+9alY2xhKidXS30g8tWeNB7I+gzl9NgWBoM/+
9Ld4HkUpbdIktj2R+xHp2IlJpMmlbCCAdAiLGJBZ9yDLcHQrxCalSrUOZwtArdui
W57Uf/yBaBw8qPB6tAeTIkE9cfWmWOuAP1Br2oOZY6Pq4Y8WiDHwlS7kMSenhBtZ
/BZ4OfNDQJQ8hPBFf0f1G/Ftma+YQmSf1BdeEOZz5mWKGcw7aaqQmyxCnPmRr2lX
m11AbKZodElGdafn9BHQEVQ0Nfc0JzxBreCNFUCFr7H+CBXahnNLW9ZNg+IW0JA1
wZPnBSHc4p2Cwwhb5/EvW+NrPZwqp8+TQc6XQtDALapPAU1+gCEOyCSr2q51mhnz
wGYWhQOfAaGhM4Ct2vB1Kh8zAEZw0r5Flze4i4YplvoM9PHzDVk2mXUUCCqOD2+C
Za1GZAKvvXG8ImNNYnZGHBOnohoZAq3b/9ysJ4zr5kp2H6bCGPNf9RjGhV2nwv2/
dDDXZ+FTHWFb/FPbL2r+MX32z7MS5QZBMP8qNmCC/KJz0b6pS32wrLKeX87BK7lM
SSfZX4nf/rph1vPXyOxW7cy898bZg9d+PW9UaCNnwAuASFIO55h9eLLeeQYwZfwL
w23MqsFKh4HBO2dnVKu/k/Ho3+Wk/9kdA3tKhHWnbQmmiRVx1pQUczj4Y+AYf9Dv
ZY7to4jU6cf4jDMk4heePNpp7dOygDNh27dLGXgoMKK+eHvZu3YizrlMxC82uYUJ
wbt6LhRUG4NxCl+pCkDkXyBGXW/1omTOsY91qave3SAvt1WChM3yzbUmEjondgso
QoR6GJsnW8wsMYyeoa3zO4nI0jFuHFysrl6b4aXzZ06vKOy13naCWt3T/+B8xfer
PpI23P70ymoppRrrdU2dVyBtaAvyizGl1nptDpl2Ky67CB6GcwiLSPKSPk/DDPko
OeiQgrEPSUMv30D/KtZW1dYVuSvMENCG851VBZz44M8a+6sWrAdZ4+9Hv4iimjwj
XhzOfFYEtu+RTZ9hOEZg18HNCdIxEfbaVDlSQZhhGBjoTXElNkPpalHYkh4ZD8UC
Z6DCBrqaR6XKug2WaV+yBtZSRJdefRf5UQ+zSpjIR+REv5M6FezU2BN+Yxc/rg0c
Z9cAj0ur4Re0vcV6GxnFsmJQ2SW0eH/oolE1lbWgrK+OT2jsDWJ27BhJRTY9mSk7
qk5PI172ZjVFsjJNIxn/i+JXxxlBU4jzVnNY8opaFbYbrohW0ZCbRE6JhuiEtOqJ
lKZ25b3ZYMI65RPPAWOp4vQyA54XMgw2Z8gfiORwry0H4lYuE/pD2/9hiSdOJHLR
4oLD3gEwcWDEpLSQnKnvqY3GFguoMcRzigAJNg/HW636iELv6vEjMqeXlHOUbaaV
WJTCxybQ/gjD0Ti9FFxc5915sEwMDTTBmYNM3NuUK0eRCY6W3rmaiBetPc/+Sx/h
poCyhK4ZLqaXLhhT5Rph/8/CiNhRiMxjU2hqpTHRO4eL6GNxzyRt7zs7++2dnEOO
GWdel73u1EYs1HTD9bzerjdzY4//FdhHE8UrNhFq3uvHHK3WKmBEiP5EL9pCdGwq
vF+EfA6P6C4ScwvHk1I13vTldpvCYT24SI/zlfp40NBoXJ+xaBYAV3UX+qXXpjnh
6kUqOxkMw1LKl0qll6mghTJDxeDKBBZwv6xwL3cRqucnJE2/JNzpdGkrrwU6cjmD
CEnUkCWFvDCxhbhnQGYiCInzpZCSGUtyF0cdqecpOQPR0DqJs9EASX5kJdVZ7BcP
ebFdkH+wGrOHRaov1wObHtZltXcaAQenE+zEvGwnqk5k3rlNalAi7mIKg6K1xCde
L24+ad3B0eFUlJtNsKqLCuoEgEGtgyoI1GCp62NERf0bYdcsUsKg5lvMrlHOxGLL
TqsMRycWXGBfqL94qxEdG9pupC8peLw51KMea6aggOZBqkQHHItc1ZF9asuloKV9
2cb6yzAeLteI5L3SAt29GZGojHKjqVZQRtatC5SG+Dk2H78Iyx+60eIPqGvrYcuA
sPT6C7ix1KsizrVzuOUEBHe+UftUfK7mWxejiy8Vq1CJz8ZmHQ9uBxZk815QJGkU
NmDjhLrQqmEANuSZ+8s9L3n5sBKRaoVe9ZMCgYwKtW6xM7lmrcw/aESJnpud1wWZ
1t+MnDQUpBoXIi7OXyxkHVKD9iA+a/byTFx1fOnWg12bSw/28MDDMbKWDoXS2IhI
Cfi7sJLvkqyCN/EURjWUM7g/zCF6fAawVyEkQYH15I+knt/yH9s+nzA/SsfHCRIP
/nA8vS9heiDHOoAYQha3NgBlqEWOFHjm6Q8tRB0du475ef2SMcT8JMLi6Q8ZhL/6
RAGHEHRw8aRT9iNHArraNH9f6YFLZ87urRbVpy//heBueD3aDIDruQu0adF5oKvt
R5l2RgU0XQkpqkficLt+5dBPrv3jKL7ZGcU8oO6fXU7dsLO9V8AIbns2+KDjbRb2
+ismcuvrg7EWwH/EoARhT+VP0PcrEZ/wx0ggw14EbI4rMGtkjRLAdLUrPkvIIf3u
1OGxTX/hz2TzEwTMPalDNHN3oPpa5Yx6GpBjemuFYXyjYr8OJlkZgg+vf4nw8I0E
G+3T0NsJyqgrzGBATYq4YHa75z5hZVARbZIZ/EcYxc8f4R56kqOB9H/Dm7Okj9Pg
onYx2Cl5w3DEE1Y7Kib4vsaEH5fCkZBgVn5uO61ow3sO72xm7kjckniDQkaOOYLo
8Wt8X9LAK37Y/bw5yjZfkjLFJd8y0ytZgYf6ZJoSIeZKCkTMrP7Jv65k6R5RKK9a
Zlzj5GK7OM5tibp8QH2ii0X2D6h9IXF/kXZBqIWJNxzlCJMZLZCyaCaAIolyqiCa
PikUYNnDOnxkDlyF5Mw46RQW7gWzyI/aki04823XAdTBR9Bpa8J0RZj/pCLU/z11
nVxj1qxG3++JvheQzmwesJ+5yCD2G2IisL8+Ku7GfS2BjWOtQ9QXBktwSkIr9tIy
/bJ/QWuFR5JBCDcA7V3OYG99d3xQ+9bYNeCKop0SoHJ/ZUwtg5KRNy6A1aqYT8EJ
ftYx/EjLKcxL7uKYTqDutC6KQOFWxl7Yda49UU4ijH3bfuUwKS2Xbe4c6/HMHJiu
dw0BbvY/3/vG0cAKBNWvKhzz5D+/dXcQT0sB1JkmUKP9KI0x2UdXFyDHOcSXxji2
+ZRpTsrQ7cVEHyfHKGOvqwOFuI8vA4RpffkVSErbnPd/PV99fIzOVgqpJJm3IYUh
t7jBKxxuhLGouaX027UmzdsZyK5r9qaOxidrVnoWvppr4XTjS0cTYwhanKw3GZdK
Oe10NkyTft/fH/YifQvnsjIreWUaVPK0xF7e+IC5Fsch8dH6rL+Wq24FeYfieZtp
RO8mmKPaO9xx/I5dU2x5+eA3C2J9wVB5lNs2C+IV+WHack4iyaZrLANAjko2chmF
zsQiKdezAD10L1gtCNlTw0UkXi9FtmpaXZVKiIGnTTZzdncsjllYxZcpz7zwYjX7
sLho305G1h4iT2s7n7INZr+U8HxnLFgCK8FFiWbqu2b/XEKWu1Y+dxjAyQnJj0CJ
UZmJwatulZ3ldrT7ldd1sYjXQRuklJ9kKOUOw25LteDRWr4A+YBAkgqwlH5p/Hv9
Yz+rvlMMDnvsV+H0nivgUfW+7KPxemvQO+0ZiHK++iHLV8YM+qQ2xgDGfHDbiss8
PC5wzPZjPyICttSKXiDXi7h0OLhObW9JMYsZCEoFyxTF6gyaQtJF6caHA6K5VJLQ
um7YFc0XYSR7w8rLhlSsKOoS5+X22JAuo9Xcp7O0Lx9hdPRsS8N3mPVEgOTTAwza
SRSfLbyGeq3ra726DGqLyWs5KgRG99hUZVtYk7Tp4AxxIGxf1+KQUtEPeBQsVeFd
OJi6+Z1al9z2d7nIbjfVB2pulOf9G6IOZFDI0SSEy1K3xnUCo3WBG3Y/SBJ/RQ41
zKPfVe4blEwEPX3+sJghTBw/vkAp3QuFWGIg+B4PnVY/UDXbcaA3A4R4eX1EU1i5
0oUp30Clcg6PYQmO7iwSYb+HvlOhjOcXcd1anOe3Z4Hi5BRsVLjQURYcPyeFsSqt
AtJU+9tnjcyV5JEnWao21gRKZEZD8EzYTLVB1vg5YJivFlOgwPFGz/uDuokiMNym
cgxqPi8zfQUAYl5ZZi2AaGXT/HbzNUw4zQZVWjmkbCBI8oJlAbfj5EZsR9UIAZMh
Eeh1+4MVKZ7/UZ1UkRZP1vt6zNbsm+zwGAejySOTdbqCIYSNkkKFYJ67Ie8V+Ssq
K1l6m4RWduWWUySZe7Lg3PkNUKqTz1q1cMmbhdlA6l7KUXk4XHPbe3b93hXReC6s
IE/nd9EqfNJ13hoTHTXD5mu8qQ9V5sk0cqYVAdw7GP7Q6mKgFiDKOEOC7L8JCWDv
HqsPmhYlic1rs9N+j9SbL/2JiDVhfii2DqxlNLknoAmaQrNERbP8nqi7f/xRCyrW
xWzaWFdzuQ5HfLJqa5anXXTbaY+R5QAAUAhgbLdDUVNfU1pl7n1sRxAi+zrISazl
YK8nFZrj0msteQzL1dJL1OYXhFLDhAsMZ+LjDatCLEXfu2an435HoCpXLcuYNyRC
5yUkU5g+nKFjNTd095q1gAM/Om/ZCIf+LGP6Lx27nygJHacpB7qd8yPGu/XihvEv
qoM7BwooF6daWe5ssd8rQvUHz2KoR4bDuMi2w1JCO6hGLE6M+1qvKdq1fULbI9+9
Z2NpmxeYswdhI0a2Y8Ho9wjWtDVx8YY/EBzEcqeJqCCCZmLjTHrvqVZA+w1OTKxf
qAdLjSJvp0CmdgbF0hL3fmx1Qu7LEgkgKZ53JRbtvrcaCE+Nsq8bS5fO5j7M1VSn
9a1XaqLzt0LFHf0X16fXxUQl8r3SqKBSADtRlbKZKaViVG4n50JMl++VDRwPVS7t
CdBeQk+7VmQzuI1ZuukRprU2ozGFm5OarKncnGLNdl7Nr0G7mESwoaiMXF5Z4nz0
gGrxGvW3gymbKsCdnaRm2dGSq0Csf0PzS21bVRGhAK3pqpmvKrCIwTMHG+YxIATw
lGX/r6r6wHRdGS2iZugsUEOIpavaKEhvocbF4tO0H7KBflmMQ//FX7WlMGAWpMk6
u5quEiZ3862Bw8GBH19bI6tirJnUBrqG4if5d7nrnoBPipyPU8W+XpP8vNmjOglU
Zlo6OKrmKmNFoxTUYenYiziI5+yM6NrqGfikPWsvsezcyw0F/07Eutv0oF2gl6WP
JyO0iPFmWRP7zmxeyEjDrzC55Z0xUNhFUd/nXY01B1YOVi5c6AGSGFS2T5Ml+UOm
UT/QytdcgHRUUoPnW8MOvg4ZvXUXs9eMiyHvk7Cs3PzXblzVAOD/R7s7eXqdvg8f
ieLTJi4QA4qkMsILxsPme3wFKjs3gN1I5NttrowTjp7KJPSCMWEnCTJiuuaFaEwf
OGUugF6VRt2nVlNNRgVzKiQy4xCuApmSaKLnE6yxOZt63lU+9Ao5FM7L97llY7Zh
b9JDKSfKqcx6zYUunXjw6FfVbbIWFx0QI5HdHcuQ70BLUty/fsFTmhLPuuOLyjXh
EhQAsfz0LOQjLHGDv4arHKolW/s6kYq388Hr3FfSXEWtHhghv4rUu0IjiaTEjLCX
rM8bGTZlc0DOzFRVHvc/KDXoRoAGWNW2mSolTj+ksU/bEslHLWE+vi1Uzqk/FlBh
PaBu7WWTZsJCM6vo8TXlSeA77SGXjdrCcS4ovtqT11KlXQmMNO5sS3h/23zWmKjo
hWHO5m6/AvuKHcxHpbHkvRuT6wB79PnicoSzConJGmbRn57F7lDskFyfJXDwitNf
R7ewCw6MlzGQGonf263583eMzlZ2OjUTcIlEHp+iEHbE/ukG8ZzoNqP6t1bpDwNb
D2GC1P3ceuqzFG1j9h9WTWs/MLoxrAkQlIyboPAudzQfFk5HdwVBofnuXATAbsZB
xI1LRUNjJVpPhFgxDFZ8gpGLUb8ay18qtWHUFNJOYd3S6MOu2rh38KJu0gD3gPMU
g9XWITYkdZ+B1uNJZXrFmKpVpyvN+D6Fv3L+EpUODEdudaEylcP9Hmr2QWNw/+VN
JFPvu1O/JsYg3oVoGU1/tT4OsefT8Vq7FpA23ZorlEqMhbMBS7y1fx+hkm+O4yYg
M0A/Y8EgloK08HOBnN7rNHTxSp2ZqkP55AtCPKOs0r54XeZwv3dmiMr24f8R53kr
38cG90ee5xt85yIkaPjB/k1wHzfQKDb5wAf/LinCbG0q7ddQEzqlkKpKkfizhzqL
RfJ+f8wfEilmHRgnQzV6x6Qo7JkJx1c0Di6R15ug2C7mhUzkZDTzLz1BU6lirdWy
sJTgZfiCsI4xSQWT/M4r3i+bCCRpzmhetqAV7KzPSUw5rQuajaVv89dmSLSdt0Ym
pdzAtfULmq1vP+DcV++/SGTBBvDc1A7xvIkPYxXKeswayFgDx9NI1wbT6mShwy/j
tV+x+gL5+TW5hQx8oRGJM5fzF0FtRTSrCuupBFL5EGoYwY7CsLm52YAWJi+wBSpa
z8bUYAptle6bbA6eSRPtwDzVul5t2SnpRDIjMBpLVbkRIWZzfDAmCk7EBGKZfH5C
gbo33UJq0000OxWkgz+OUEQSfIYL6/Uia/iQEkBrVXiWnBn6l5mwTxLgCZ7aSXSt
Ei66nCopQ4k3LLFa6I79lEa8wSCIzf8rVOphPLRQdHtZAxiei1YkKvhXqbElrEkv
ryqeuFL0jSLP5+UQmz/gnMRItBhruo+2vZrqEp9sgdURhnOUwmVqEQys1G1yQHnc
WLy4U34hWlOGyw8eTtkG0PlB0NACaLb4rEnaJ66bX4XJ7vKucK/uMQM3r+jEO+NG
WG81gRmJAY6HhupE4haTPy7RgY8SOyFgfVkLqMZBO8uXeI0/HpfRvTWVLJGKboGS
iVm3d0m8KCyZvlZ1gBizcLDvkWQMPIboSHyJ0RpBawYu9yNX5gzJYkOtSwA7uP7B
5gnVzIRlr1jJDpCkwMutX4+O/7qY0jxkWjNCICBEuYWEgz0rl7EnDV+6Wyo1Fp6z
0zl9cWN0r//cOaW2cFFaG00EsgXVQ62fDwcWaZ952Sv4UrWehGG/L9Gkf1HZkVXD
BAQxFkC67vNAv9SmqR0dAwZYDgqKscBimxBVQ4c+B3Lkv+e6OgkSWiUCksTpwkFP
yGd9umiQp9Ksha/fL7pmyFld2hQGBCQgsG/7WgZpZ4GCfzXsUJHXI1gtuIKNtDWw
yYTUlRx2xrLadAN10bGeSFOayjueKaW42cjWBM0P/l2MV6aff2yBQn7IoQfmThsY
afPhjcj0fseiuPqpBu8MSlrAH4ffi7h+CmasVWCqB9MknS+eHipEexF79tDNROR8
Iueeo0Jz27Ex4/PpqFDd0A3TumC85jTtEDhxUPj3S0dfNeDOpIqn90zZYIQ8yjHK
2c61jIF23+WxBQSPPZX7PZyQn08hTE8mtSR1GuNltTS6CsTYPlfKBoLtbD/y1wOL
4HKy5eJpaP+QkglurxDVMe+czLIz6ob7282EzMKGYyc+IOeWWQx/9AG4ph0bChcn
aqKaNYl9KOYl/x8trKJTGWMtx0OOIurO2MZwWgAYbQDsHu3akzRxOjxBXHGHsiBq
ab0clkhPpcN3U87V/eIv1ADTQnUT4vLGiTQR6foFIpA5tfnvmNO4Hf0KFOakKchh
2+dTTKezk/3I+G0Yyl/3GfoLmQIbidDEXORGlLnGYE20NDKbvBr1i1QQEpTQBwKr
KarbRlCgdTI8bgzQz0py67nRos1kuhnLAdSa99I99Dm6rooeQHCZT1vWV+CWO1Rd
GBT+tvakwRDttMxDvCh6Z9rM3bzjmhbSkeN9qAHUEklFW3rh3w2/POkVmlSYF0Bg
WGhF+zWPhrHvQp/khK19YLUYcRyTqIsGBSS3FqiU8DrMqm2SVe+69jYBuHaOli9v
SJ/b4wBfLT1XN4yiH7udisIhK3Ab7Nxe5dWpjD/uO7QKtJq8CPS1o+VYFFW7+kev
RTGvZw2WRns+c34sBEN8aBk0d57bxL+fTus4byxdmPiOy2inHVHED71+imXbhEhN
idSobI0nmAQz6kNJ6/byxpBmTX10OKYk4HwW+Bo4Tp00fVjGNjGWOzWfurDu1RUl
wCO7yVCKLDrUJ+tNHLc9JvLKBMJENR0S3xeHQAyx2rrTWQDmYSEt+qjSZEX8K05f
m2AqhaBw0ol7AqqFmx7R3+vRbq40PJGKk/aDYA2Mr5TO1izM5vlwn5cV0iV+PgW7
e4hMBE9dRwD9wBwI3MQtFTzbXNJxoyl0vOoHBmBzE1QVnIL61Wl67jEI1nuCIVc7
G8mEqcZmhfugLtIuWm7ddWURNO3X9c1FkU2o8CEQF+s60XpuxZ91t2sVN63P3cDR
y4/G3lGRjLJmVBEKu4s621MtFCELM0rnEzXr2LOOJ7y8DrT05b6HaWKJ7SIMgvgy
cx6WUHLy/pcLxx45qRG2b+2N5X/qK6YtXG6a4QZyWpWiceJqOZ8y9G6osjp+XLjq
2+KuIkd4eJdZ+svo4fz8WdlzEmwFRA5giJjubp1+R7Qz6k8u7+D3EZykKj15GrLO
2CwWeF28kPGDRjw/dFyBpMmeNrNpLSdeMB3U6Gs4gbdDaK7bIY64z4Q79xK4PmYq
gjxWxALLfX+UE+A/n31xcg4jdd7fKNCfTThzYixDFn90y0ZdSH1P2kMBLvtt5IhA
/ceRCuSVdMNQDBg8aJfnnJAN7b673n5vCCbfMbSHpYUNAE/mAyxiSDI+ow0LhEYB
lZxwBwoqiNBjGClhlu09TP9gI8q4sZdCHForyVgaBTKkjwvatqoI+4P606b4dPxC
Ma+pTAkf7huSsuWqYqtwS8CSKL9suSi/m5aGLol/JjIY/AZUf8aUtpwyFginswhB
vKsQiJi7kRNwNcRUWhh6eFt3QNMY4vieRuYs4gcb59p/xhFBuGPOjVTzfujogdsY
9HlY2+AbHhwERspky6fxmRudwdPdLxA0fn/uLWWTnOUNIGToaGvJeRK6VMUb0rAt
Tr/KlWPiZM3DbE1MIQ46zlimpwNjUKpXChnRGvOEeUzzD6iTS7t2W9VpP6upegSU
8PVaqf3sKRwofbldiGMOy/nae3mQ5mY1HZA1Kkh4ONyqX8EtvYq4dHwhIHD9ta0e
MQ2eZYYGvMw4f/lORd8dSOM/WTYtV5G8+Y0vgu4xP9r28/8ekum8de60qZ0r6QFe
pvwbasTgeW81c4/iPEOBqj9OzU1e+nZYTY5sIxNSCZibyMncgl3r2bhiDiDTAlrZ
B1Ft5QI8DtxRO7mcsX2fVebVHjwVuNzVH+guvujY909zXo8a1EvYHnRas62/wCqV
HI5/ItL2LK0WMWGlBbVERkH5eIzcSCEC0mI3yUAY4Y4MzqbgWnBxJvnnHmuIY+5Z
wvl/ka/LtJ9qiDunUDHiSOUkujgZsppaMex3tDzGCVY9wqxWxyDDKoYr+JKFB0ut
obCmaIoW506efB6PCLVXEiKKsCIqsZlqRoSPM7ZaJPhhD/olADnq8OOlk3GVMHyC
FnHoOwpYipoZMkW8v3qEQcdN6cO89OOS1/UunouRyIXST9GoShSc++cG3ujjoqFB
gb+g3YmDD8i9k4ObCxULHgRrQ8LnkSKgn4XOHsbVNpih90DwSrICMysybWjrA+bi
nXIQSRT2bvjZu00fQZH4rBtB6T2n9N4eXyD3xIsCIp+9+9uNKD6CFJero2VwhCtc
KbJmvY44N4EMfAwKLRb1ICHdDjIEVH5JCgIzJYVEjDCLxbXR55MlNVcCJan/PLnQ
cC6eqzDZL93NJzb5rSchrcJvqB1e9EVuM783O7nWo2Qa5rtxhFX6kb0rgz+M/uGP
vouk/uPTfR1F3xC1xS25gYjH0dBfFtE2zrkPqClcPPNrUfN74eUxxeHtG8d+Y3gP
tciDcge9lKsWAw/VMoAOtmZbugUrqOYwBCy1gRIFWeapOrtzrw+tzKr7QnG6+2/k
tXX0lMK01a6k67RNh05CBN21G9GVLqF6lXJHf38g3G7sKDqdVuemB5nEa9FdTo62
8F64HPxXCO5mE0sP94wPG0bwIEpdHlig9+YbLAFnjmkYf8RvnkhTbh/6CIiBZuw/
hTsL2NUGMZ/o7bVYjoUMA8odQTfWfpy1PQVUdcTYI5bzcbS7no6CGLd70sY/sHCQ
ZeSM69DBbUtsVV0Zmdz34ouacUj7UT5aAQPTk4UGQL0+OG02hIEj1VC9XOPafzB7
QgM0ERfXPnUfU+emMHWIS08d24Ldjgovj64vt44H1qGJOtcwtnNpH3e6AWNv2x9g
BLbkggVBKqKDFAjpgXP/v5EIlli+Qrbh1uArApPJtWz3HlipWavcKX2IY+l8MPwU
PsaI634+5cvW/ufv+uE+9fXG24EoCA1/MnQwv35ZmxAN7Gh9tCroRh6H06Nc+tEt
N3dGE8rsC1TfobZIh5wjTsRP6YjFV0Yij5JDpMW3R8WdD0pt8QHmA3WflYV23dKy
ZG6mjtxna3kFqYPaVClE0Mu/016rehDE2siD6vV9i5JBRsQFjNho2ouXANE831Tj
xc3RjP00URE4M0eUfuVjUMEm/uPogWVjoqJ7R8DIJgrX88L6UP88jOanuACko0Mt
tklm0ZcNjZHYqHAzubbKFnT4n4FX9iY2FgkbmrAxpSJCXEZQDICkBYib+u9sbgE8
8m8HJ+ywPAxb6HWdXi2DTOFvspA2b5vuyXoKPAgYy6D8zscn1FFFGZaWMgXwBGD2
R64aAsQFfPqlniw1lf/3XIghn8zFdl9JhKn361zOhyy/9Qc1uOPuHcaoBYq2Ho65
2thp/r8OwriUX0L/Bk1Mw9C7iNKx9rF+i6/ze57+CbMtHqBLHHwzBdYLCN6Ov17c
rm5IhXaxPJnlg67BJX/AUDGVXPJA+ZwfX0Q+X9NIlMWfdbQilj5wqRz8PlR4pC+7
gGGoBHPwK7TrnzyHwcAzSCzcIBhUbM6uC4H5FP6iUfNLuH/FwMI7IwqkeWjQ6XCh
Q9jQDY+TciFBK42ETrx5pR+lrEzBKTDjFWwjiiX0duDVO5awHEIJMWgCwbV2niug
cr8mRiCVhJWiL8BCrjZyuxFSrP2ylUx+jtBXvP8w7opEDE8Nh2FeoBQgLITJN8Hv
yFcSRaqOsVrav03bqayceb5O+Y6VgxY58LxtwR+1n4uFwrOCFxuDWSud8HYb0+dl
I6PDRQYI7CytyD0rqfrSJsYHTkjiH7oGpzQSL8aWKIrfRXiavKM76ALHLu2TY2q6
UZe8bRZ5kZjL/Phspj2VZciKNR1J1VO9Y14VuCsfVOElUNWi1Tzm3so+Yr1zkpNQ
oeeRJKhdjw+ievVh+OsEM4iMl9xWIXW+nGwulIZ51if/5674nYPYHV6IOX92EJVr
IeiWDFPxLPZhzjPAqhnV+IP8u9NjxZh9nShcOCHx1bdeNNyC4Pv0PCkyRSy3oqqu
2DBK/PpfJEt3fYJgcldj/ONysiK5J1o5l9/Vcy06dkZOFmO8zA5AUy8ML89kqH4q
l1fNv5ny7T2fERs7iMCNUoP+OcflEfSKBbQ3xZRcv0mdYYk++csK2hZCyAZPktrp
Km7JR02RztfB76E0k8EbN3M7Ig5o22VvIgm/8RuNZkYO2cIMaPbSbj3u95C9BVFW
tyqE6zRg81PJTn5DKhn7qM22SynFbfLq9XHMlQ+e3auzZk1UAIGsOQ6pd97olDEW
lFc8nJ1oI2gsfo3wiftrohfBPNCJ8amQhf6fuGZNgKltgdRwiGRRJZbaSZvPFs6X
FqLiVE+f7YZ4ezWmUrm1cMSLIC1lkS6YaOlilQCuhJLNq3Sk7b6jqfrfOt7aYNia
HPc3urcmQAoxsuLJmIHZJc/98Too+hbL1dZLR8jGnmcdUeZI5P0vEWem1PFcRhG+
LvPvuhRXwSppzMllah/g7QRHmJIN7mddKJ8Xv647gURIqeroEh0JsA/yh/MwtxWu
LK7T/xR2DvVB7Ory7Rx7DXepv1I5NexxDGuig8piBW0b7xHxhKyFpkEzg8tQLFx3
/Y2fOXFC7wgo0KuSmPw0c+RxkL+7Gjtv3ZAHpkyxbxIhOMQWowlKI1XramfVyDo5
QFyr/X8ghI/womgU8FbASEJ3s8VimeDTk7f/EP9TsFzpeYQId3WFf834rMdjeIJV
UjY1WNvJO4/sBWWiUf0+AOvnqVHLvpnXZV4/D8CcWspShoR9rIB+34z6InlWnPCU
D9FicQrMJjafGgPV415Trd5fwvf+N9gqBjzmry7xkgmbCeTs9Ff5NHi6wo23bKrZ
r4wkdqwqTYRgLgnstuNSRtbO8smUG27/1sN1HMz2+LPCFOP48MzPh5IPrrn2WSJ0
wtTVyvT/FPATSPEtAeFvKtSWhzM9+Vlew85HURvbHQhA73bHnlLgBtsQGsPmg3tP
qhW4xcFM2JDzc9aOjXGr9pb2NWVgE9a7kVbW+hn7rY6kKVuZYAwKDWBsAJsGUbQ5
EkVlAq6Q/iUHXHI7ZHtXC6HovQYCxuIhMjoLC0CY4HDTEbAcj2201nFWoy+UCi1Z
UiKqElet/XuKA8rFJmm3YuPkmfqf9FlJYI2xl4fF/KJiWbXIiHRkNoEUxvmDDEEL
zVuKKo8Lfrbrwy8z1+dirFSBlDj0SHCNe1vS4xmxWQFJqp3mLoT5lr+6kSjYmYpo
xIrZfXBFeFwgI6F/9Ise+az91++aCGY14HFJkCErhItB7Kq2baaG0PjSQN0KLJwX
2zjhoWyvwXZNHEl/Gu2xsT5vwn02JcCtfG3WVGjZAmC1KXqXAU1D7GXupAs0JaNf
tCgYlF7mVQ8nUuCKf581CremvyoN5QMri+TF3nUJT+JxztyRJHiL2NO7jrqteWl4
V+yyJs1Lab03oEAr9kFBobX6+vTMIYDc0I4B957wW5l/0bLOJtxS6xqZRb5+mZSa
OZ2lWcI2N6liINGNQsoEucFENR8BuB4EsxoV1XHEkQduEvEC421iPveBEf49SPo2
ES892dlPVjJ1Y7kkeFYddu2fxd9ajJaEBS/RmYhUZtyKrxqknBfaJYfCKq+Xswdi
nEIEYIoi7DeuGL+4+bW/3fJ2cG2r20GJR5tfi/9SjFUFKPRciISItNAK1hJjrRZV
bfO9DaDvs5rsvNjV3J5nRXOCsh+oQjx2ggWrN7rMmnKR5qxqMeSljuaLUax74E6T
LlITzhEIUKN8invq++xMyUj1+R0KoJfVWWQiVb8bR4dc+QB/4PKOYIFueTeXsU5G
wHG5h8emQNlZJ5KwVrLClqcJLzL4vXll4jwCeydmP/P7ZuH1II4utfrN69gaoTY1
hbgVXqC5ngVRwxIXZ6uSTEJRs0ZwR4SGmeYVeAWKm3uzNgs5F2zsWjJ+00rbCGa8
02KGYUzpuGaIymn+p0Nd/js2NC40t1wYr/wU5cdAHN5z0wtTQir22JezjtDw8D2e
USa9EmK+6S+uU3d2OLdG7QP+hXotdSmavMdj8gJL6xbfOWbDeTxPdcO3Ij+3cAQw
P+Gj6fsKY8l2yWbMQNo/kiUK4anUN/ZvxfXUkrjFduSHGmaAIJ9UrIrXaaRoohdH
gIBQ+/5gzZ+Ub+DvOXJ6p8qUVu33KpUge38paBiOUY4mEChCYgCz5eqcW0A9hZ+p
QGC7FjIMg/c8xLIPCH3g0kMvt18D1pa+0UMGod9bG0y7HAxDMC+GRl7WPLv3ymRd
VVVU+dwt9tBe5D7eOnGCPVSeI7iPFGiCnN5kKw0lldwqD4qDgOWuyhkLJLyOZFpR
xKSW/yq/fuP9+7eSOUpqxKCGaCLCfuFpFwGZUJIoTcjyr65/+qaW6JINFzUS7cBO
KEYzr7xtB1pmzTHNQTbWMf50ppq+SYcpEsfFOCXw5lWfH1GuSxsXbU3y0ydyEZy5
y2V/82qFd5yvn3k05HczEiIKhw7xYoBC4lxRLWVEkRoiEqT6sZAvFB+sgNxANrx0
2LDfkRKMzpxdoFOj6Z7JkNmTaLroMNJrYKxkVjL9Eh+eFcoFuFUt7TUEgeI+Evqr
KHHPnGc2az7kUKQV0kWdUq8/tGbuvQkz/9GS7wcHUMICzLWoz6fUD4C0Awo391Pb
n3pdabjDK9E6cXY6Nh5h8b5aG+If4xvE2ZgdxApJRFiGqKERzJUGsF1bUjy1VDK2
1Mas4pMOyPUbU7mZa9hjc3Dv3ClycZ62cCwT1/Vmk5FZoeWOs8/NdukdB58fDc3f
+ohf4h4/1Da4x8p0zr1HWPg3PlvUxlduYzV4zhMcWgsue2HZcZBpqntFj0J9sFYg
brt4rNZzRWUB2XhFEeW8WIdLwHINExBOhINTGw8FuMWkuYc4xhak0m+SVQOie59n
/awz9ALEOxs0Ywi4ckzkEx9IHeAH7CMQOLOOgp/eEZGYJDjvGXXY6xxvLZ+VTI7b
fr3Bhh0i0D+tJaGdGPrUSdQC/qCgpX8R5bxbBaUexYayxrjTZ+X9PiVwitwfMNB9
X4qJ5HcJI3iDTAlyus+U0WWS4aEf8ojO9ilmyrgUeSoGQocBWTX/ix+NLEc8KEHf
WvtV4jZ+YFf5SgBgCdlmFIYBfOxpn3v1oEIBfS2+gZAVCF5DkmHhIu4xKkCYeUd7
YtDXZiUTuUZx+2KGOy5oZrMEbjKoh/A5P+TEvpezPy+QJMeD7IZR61YOwNNjy7Lj
zufSYAIav/qiM4yf0PaqROxuUW6ZRW6Gsx3FS8HEtk19kIWQg8jsV3oTKW2IzeNU
ZGg015y5KZcz1SJDOGEMnYks6Ld1cC3RewJfKSiPx1TRLXLBIs71COp81N4OZc03
lSwPphPZlPK5QI2rVG7v/XC6dCQp04AsfFxTBo4e5+ZVuWVMyl9/xLAXv+ShJ8Z7
Hmlw3UcyVmZkKYOVhHH7aPoSpy1SefmID2OxZuqJ0RNM2cEoqvxYEDhYrlNmfLCc
7YyS0t50YJeQ6oSEzVv2u1I1FF4dtWaUx2YCW7mR8+5TjJqy+h/amsyoldeAbS/S
Q0BNtOKCiExIAvr3om2NJTWMgmizB4z9h3aWWnoLrPOq66UFreUA7wI0SGvLg4ND
v4Ljhmn7XlM37son2nG5uJiQrdWRI/CJV9e19wTrPsTwhXWdiqD+JYVAQGisCRxA
lbNfIQDF+SDCz1T3h+mUoIiGIhu5d1J6G3wPPfA8ow2NqD7JLYba2iVHdPWSBxZP
i0MSCf1duAI1YhyEzs3JptKnelvuZM2GVprfM9bWSZb+s3ZBORasBociL/yjPcgq
hqiHolF1rr2hGdopAjeyROUWSQZjAW2GmfReJ+rIgZ8RZA+QuubpIRiCaMiyRufW
vg89g3PZtIJIjXwHtJvy277rMu/NXIvmGCHYMGFYS47mQfLwu8eIRqZ2nu9YSrgD
489El9wiMPqZ1nKwdEMfdcjsQc+5Wj5C9Ix6ylrhn1FG3fi1JeFgWaJRlS8dauYn
0hUugj7nppFVZZuYbTETUeE65A0uogSX+KNen76pZhSnQbTYBuP/KWZrCu5DWYMM
m7if0ES+h0z/Qa6a7QamrtmgycAVPOpPrxWAXgX5TrReIgpT9CggN/XNPvTq1P/n
+Gm+Xms7QwjFRZ1e1vOe1koAqFCIvEGvDzfDCcz3ZWJ6Zzjp8R6XI+CsaPysJd9u
ZF1jhyqJljr4tT7OtJn6LX2Klvhvsr/vhkniqvHHnL1YRqIVgt+TdOixWb6EX+gA
Yu9F5c4mu35rXjor8AHGm+5aoU3WIKlH7bDfQoNb+HHsABg69hUabrFonal/1+PG
4ugR2OSMmxYyfRw9m3fFYiQtSxOQfUKISk7XuaX0y1OkK5vwl45EJTSj62KazNN0
d5yDZxUKz466ykvbMgR3bv2/O/w5ePpXmY3wa2IFjG0BmeAL1NYqecw+hz4MEAKU
v7qJ/qFNWcwbslZhVoZKEO7CEPz+q30sbQKJTk3wZFQIkmrtmvLRXudfcReRhM50
mrcEhu1F0OQzX9Sy7JPCDHWXUIkkMJyMvZ0L2s3IrHHzzGiZKOuOVI7RtG4rEAjw
PdriLEC1je0bESkBfQuHlhFwgiVc/IokBMMEcOFcrzNKhxQDB5GeJV24grNYz26k
mXXwnnoU/rTzWVzYqrcm8QWMPhYa7Bm8TLyPX2VASXbjcEqtHDxD5nwlssFCN+7n
TqWoDP7vYEUwfk03skNY7Qr0I/tSSwvEZmJFJFTcXSU4ePZ45Vi7IS5Cz6wwFzX5
1JwGulQ/+rI8+I5gI/SrdmPwA591GMIXKoapASz/fb3HqpCHHT4koYa7Bnj2HTHU
1novRw8UkhyH8I5n479feS9kAotxp1o7oWLp7tOxr9MkBwcMi/tstlU7PVcNf89T
2x+/l0dSklOzuXW7bZIbBXxyESDzjuunJG8cJV7+Qrmk4vYCNylbxQt3G8P2sVks
aSagezSIALjPqFBDC8AzNBzUA6f1X5UUoaXEWBYlUMoFJXb5jhBcVhbJy517x5iX
M2wAK5j51YxrLYqkHVrYSqyncXyEsmGMMm/asUH2LBVN4rdNCzGpnPYp2nb5o/Rg
INGKRYTmUJzd5oUnBq5zwY/EIUd0jMM4bLq65SUUfJ5Hs4HdET10aokyetQPByuc
I/JwnlUNbeMBJ0P9IE+T8sHYtfLXX6HEfkzrLoWhKZDo9iYW4lCQC0gwxq9r2KFO
CcOZkx5PezknJIpszkuqQp5hCAh3VcVp1knnHxqjSwNxtoASuU0MLg0OVf1v5N6J
7/RxL8UcHT4vwrLiYaBWMmiHSb841vExnuQhDwKXCDy5FaQWZ+uiBM2EIMZZ1Pws
1IoVjUAMncdR72Gby9qN6G67X8JvOq10KZOkylnjy1rzHvscPDAMscgdF/wUNU/G
31jILa0ywBeCHaY8zfIKHC+I/upQgLouq+evRpkIRj1apzFNzuzjgWwdmwSCX2R3
G6pPqoyg9f5Nl1vmCpfEMrIiy4FbLTAeuHtm73+VjJXLn33cjExsIZEYuQTMsXcd
kDTt/EHw420TPsnakMto6deuhYem5u60YooRFECWpruoIb+ChAKWzNlKL3xwh7SN
Bi4FR3R6KfHKNjX7KyI0bXxLxm7JVccmq+gTeA7TyDZHTm1zj7WdJ5NlPasZebq0
rsWBG7MB1u2+g32UVSZ6tdU/4WRaxLLeqJNSoR8LowmbGldGM0rZkDq+YM0A2qIb
u+vsItT/PCiNPEO2GZiDCAN5ecOUfGrxg/vLDi+0AVKfN/4TR+QrOma6/LpfgCqU
RkcF4Ny+Vi/feyOE1pzTISpiooB74iHyjlA7JOcuRx++nWN3w+O6tyxqKyRnczOk
f48cCO+LfRjqnUSk0bWpFsPugD2gKGEk8eQYK83+nzesP1zwF1KsMXv5+sXxwoGe
hslkf/M5q8X9DJBMETqAhGUk81mJGzwYGMps1dSpbGVoZDj2TCwFEd51qQ8BvcD2
8V6lCJV76zhpJVgygVj3ntxTI0y0shoNv5O53mno7ctYOiEbJzgt0A71SPKaNmcO
A+OKHdVM27jBVlSyrUzUOLi2IC5t2hSusRiHN7kqDRJi/nb7I1YTPSpA2WTAvyOy
Zr+c34rr0k+V96opE3eV1ELh+EvXu3eZW5jYXd/Z+0gJxv1vYtlwZAYlBOof9rbo
No8VbfGmYEEajT98iw2Re7Ve4q7Mtt0tBXUMK/bGnmPCD+6bj1Eq0CCit71z8o1G
0qCqGkuRwNrxasber6ujHb8lfdWGhZ6vj4ojfCdFMz3+Ii87SrST4C2KHdTr1t1R
vs7jhoq5Vxx5lmm0lvUdLzyz4yjpJuqmvd1YRayLGIImqUYWTI8c3s9Nbx/HTAMx
Q0bn5RAgIgbYLHVkESzWH6IcUv1U1gDjMqmjLNV4m9WF1wviIsXH3zcNegDyQ+Rw
wiwnob77blQla9gajyzVgtKjAgAopLoHFqM6rCxVJv+JNlBB/lt/znP0mS/BYPuZ
5Ir47xDfXJLdJOmjXa16VeH4tPCdJd9iVDty2Y5h94m/FOCnX1mpMO4dyRt9C+CV
OEuFMvvf9LS4PwZMpSw1xmu8R/QvticYm206KSsperAxZSwtjraU4vwoqPKrA7Wh
RbqwHYYhKHZrmFVc9dgFA0/fCbbsFmhx/oQ9zqq87PufpOa/hTZityBXt1aXZHCH
dtar8o2nWKDzCi8AHIzbHWlISPw3IphWQAQbP88j3e/0HAmQ1Ipy1yDcB4ZWoTNu
t1cSQg1Oj5/BXs+6e4YfG0DxpaV5DBShXm3tcG9v3RFSJJfNKWbujx7QBpckydO0
sPZFCV/itig+4hUph+PaVRjGObVgIx3472d1azVc6f+EpxmHUG2Cpy73YFvR6JR3
pCXd3jcoQ8E/utXJ8rpXSifvzVzQ+sMdQAqCHClyajvK5KW/87tSBcajrNpbh+vt
7q8732qh/XkouUoutCc+F0fjuwsFJKYXQ36J66cJmwovwl3hN2MntnbW6Jfe2X1Z
hKlgh7uydAX+qcJAF7hhnNYdufdSiog/CPyQhf0ly0rgi44iZRN1Ze3fFMko6JpR
+oB5Rd/5gEZevHLXqH885FgTSdKW3ubLgUg4Z4jS44DmtZ1hIFrcQxTir1nwKMCI
13VXIjdToxTwOtlNu0e688Mwe5ey85NAvRpyKvRjAuBAx7YD9eKcd2gae1cjNPgY
PUrbBVwFx7Hz/tjytAjYm03ZAjfayno5chbGrwUgz8pdJDCjZPOJ79N2AFz2tORt
0n03hIMrRVuyeytQ09eisEkYAhR8RKq5259eQEUWbP6I+5RRuAxYE3IBIm/gDqZX
L2s8XJFXzWS0yBRDnSYJkmzyvfowS5oa3QgNLl+b2NGeGXactOfVzD+PH+uFeud9
SpBTjyrv85PbdSkkbtPKHweUVMxBUi8SVlksQvt9UEMZ5yOphik0RfpAn5WL5kkK
IHkWHkOJnkVfXrOx13kChK+e+2iXaJ36ogOCnmS30blCEbuP4+Rkm2OZhrPQcrri
IUVkmQrafcuFhpuvu7g+q6yZCMbF//o2RTECJ+EsYYRVhDVD0Fph+CKcEBqJ1JqJ
Tcy2qUPe513ir9eHrQL87fh3ClIANEvbMpkRY29osUsfSEIK9SO3pPwf59Q31EcJ
rg34IWGj6wXG7vpAnIb11nbBJNWUZKmcWime5QKGjA17MDRTSrUvonDYo44nbAp/
RmQCdkQDq5NmzbBfflQ+y/WDRlN15e3o7F9KavZ3oL+dy14YOUioYjuFSPea81Tk
xss5BdFO48pAC8ipsxu1iG+290JFXKDuGQYBbaGQRlIZpSwOnP9ghN56bNUtrDsx
0ICZAoHgFuq7sGUyDubiidqyCk53CyGfAlD4XhfCNZIyBKYcx82UpyMHY2l1w/qQ
FMD+XDKTCnU6uBnnXpOP3b5GI9QPVorOerYCb36NtgQaLROw/kzGpS+qGkfI320g
WHzgZLE24mXBUOtb2wBLqjdRK2v/ponk9qWwoilsN+CQF7+v80P/mnFOK78UcLZJ
7zcfBTAAdWR2Chcz7DaNeNY5xHr7u8lOWiX3CMu4PP5M09f1f0dEfMb2/1LbgrWe
wx7GFT14iwo9mwQblEk5lCeGOknZDTT6lWG3SAeRJfqvBHG5IaDglPu+kwGbUfpF
ukKstsPnJkWqAF37D+jTlwrhWmVumq/GeKphpauPbjPIeGnZVaWJnCnANA0kKCnh
rSubXkalIcuubn6IL71ozUqNprZBmRZn8LGpJTrV+FekbOPXOYNQ6jFV1Ua2F2RL
EZieJ9ty+GaCvZaYe75VExeIoRAEyfXAprPjeooI+TaFk7RChzPJsWxy7+s+tTZn
8yMI9MhtAhiG1j+3R6shJPO2tatqq9vUTvdg5pWtvylfn5r9bepTibs1bV/o3wTI
DzyYLlbg+NU8v1TTnE0U6cJkb2/7UpT2ZEptYdkCjwRmB2ebuwWrg/wIfBIEVpu8
iF8HwBT8cxJkZqy9L0Y2YzMjgduoILe0NcW5SdzXxgO68xHCYyFR47CsPmxgGJ6P
9UJuk8g0POrX6m4N6viXPgiosmHV3rLWIJSe4Ia9yWh/JvT+4fqS6qFZEfplHI2x
TzJ8jbe3tRfoE7qEGO2sT97qU7PsRsUGws3vvz7aRaRpEJP6xkkOsCadkNbAa9cX
l08Jo/LdY9BzN/lVBoYRD/2KHgPGyApjo5ubjVAkUTRTipk5Jz9WpFMyKOPCRhYc
vxK44o43s5oHo/ZZB9gBze1TiNqjuZPEQZ0gBbLJkxGCAHiyf/SBVFenLcxUV9GB
qgUYxhJmDFWe1ATnDO3f+WdcgTljqOJ00uA8jAc6PQuECXArfdoRejZ4QtEkJG+q
jxm2GpdbXPuaWMq+pZZPm3g+x6723q4Fk8IrjLQ7kFf2KjXJiLBMLcryh/zmOxdQ
jSzMyPrG3nD5EkjzN/AAYvARIxvvjMT3/ekJBFgMifE/dkNfy2s6Md4IQ3N7vVr5
bvjleWK+gEjEKfL3rQ75BGcz42giBYFBB/4rIh81Wvk2W1sneS1LcWvalkLGhM1p
bZRMOaV09DVV3ljdaszNy/tX/r8KqVITJ6urpX/FZ0PNJPiQzrtAkqZkV1bBiOOd
if1lNkOZnxhmdnsW1CtX854i0FQLqkO7VszkGG5Hqu1msB/xcliM2nOembaFV7K1
ryIZqxn1cqKypn0EpLKJ9sTKRsAgFUVE4AM+1u12jpRFK8wC7n3Wl6VGUjZWLzGw
LaTNI05sHSqb2qIl2HS2PfjSwQUndfOVB6kj0sN0SVhEFoUSaVjLm1WWa9VYskeo
kmUBD3kdCUA2L/wpXKg6qvYM52cCykS/gON+P7KnJoHwR+VYcnG1caW0mhsqGAPz
ZVl7WTnu0kY1Ea1zMR4vrZMrV/EJnLPdyEZI3PLs8l9Agh0iz5h7iQWclvm3YdKa
+KZbLKcq6iCz0iMmBeqE4/syhYn6NrW+A9Ky/sO0evA0Bv5mse5HwpVLKNpMGLFx
wpibBIqAZeJJLahZzPiVXMW8QWoyOPRXofsWDhbk+YbGSVhtsPe8huiDCVJXahCR
uVktSzgkZIpnHgqVV26LP65jrCf/RGsdMHDrCOs2MRAF0D+4w9iqZ3ayunoHvP2e
qFM4MWtv8pPBdGm2hVrx5V7M7xgyRZigBc69sXzPPQafk42PbUc0IBrwQv5Poos2
EUxvfFHtKT7OfXzxDrc9faukn+BBR+M1c0ixBstDE2oAzY9YDKcp5+f6+IrhPFVx
tK9cLRLjMt7DwzSPwCWglJnrqACqF8dkwGlUh/B23ZrFE3aCYYMMkwF6CIrc9AlO
BC/RRjLGljGR9Q0+w+dQPjYN6RMv29xKJnnyHKh/oEiur6iM326blCtJZsV/EkRy
YAdVKNx8mMy9piNhLstGFI2YxukjzF5VUZSLVIpxwjk+dZRU0HyXq5aWkku+2VpY
X7gM/qqX4RVVakWzOnV3+5DakGU1GgcojwRFBqZtI5TKc1/KD4hgrnCAw6SAhSYl
+Qla3AP+6iZHmmFJu+0G5H7EU1cQGYFYOAD41d3QrYX5oZIaaapiiPGyUwkNfXaP
IRx7h6pPXKkBOyiM1zQIWDCvnopRb9WQorVvb18Hofr5ZXBVUqzW/+JYV1QLg+Ns
ancIoBpTN3MkbSvX/Hy+rR3X6gayOUqwl3nlYkIGE+S/gqoLetkXqqka7BQJ+ugY
YcL4P6/So0iSeARlWrtxxEiu4XhWJgy58j8t3PBQyfgF6ilh2VG2bh4BhXpSl9z8
LAcbUIEBbMm8+Ur6tbDKvgLXrqz9OchByKL2o6BUfGH9McqRZ6vvYQojYbjbl1Xt
DISlFRGpZy5hSlaG+nDGM1vLFOmoRdV48k56kV1fERWHJoLnP1LX9bi4SZ/PWLdF
o+UjBJ7zgzSj1ZD/mibE9bXEO14e8dLfyS6SDqGyt5/RpWnWduJ5oFvSimyVijAo
oHY860R9tIEcrPTsbAfIGegnCo3i7iMIYY/q9oPxoLovPG+voOx0qdjqmY+lLLpo
p/HbKO0N9RtbdKRkqgqBjn4IvdpPGzrAb60FbYja8N3eV9AFL0DGMalGiicVg2Jk
iBVNJh4CC0Z8RaeRe0aUlA0CYoobyGQ9ZA1N8fomnBVV1YCudrexiDGEgQe/tRZR
hKXWd47MMJeONbcTXkQ4eqOSjme8UDG2hmfBHHX/UcfbSr8Bm7N5YYblBisufmed
6s8Mm0r6PiWDz82YrLXZ4ZD8Oeo/QV2Vghp3w0uUCULVlUlrti2QHMa8y86ouUUc
bRhImU/2CjAAe1/KkZtYuWAsFcjvqqq+LFOBl/oB52n/EBdUKQPlIInhcjOROhUp
5fJgAGS78PDzQTHWO3/voNN3e7uPRfoTjBlQVcF83WT4GMmwRUPGsIIEM9M8gxDJ
HEb2wgEaNnNkWtK2Qbhf/h36axzDc9ipxTSRNP+6kxRmC4+rHd2jlHt8zafLDPgV
AAB1xKy9Si/AgJX99jT6IE2RnrMbW4krxFr8/7RXrV0pDqLa+POBU3S5JZ043Bu9
u2kIqXao7XcMbfBK0cSFZHrtVc8gWwUcudQMXoYTMgMUKmqQT+SMCh21EFXF6JuS
yDS34ybFNEOasa3oi7AesjAv1wy0zAqUDtiQM5ojlZ7zXBkDTrkSRfrTyvvnC4qE
R5+Rr5xAFZN7qAlbiYyWe61YzDg8UvNeQ5g7CvReiescZ4T1/YzctwbhAVclcDwd
XIkN20C99k9R+k5vk2lRIpDnq9zjlqPSQ7HdcwC2TTt/5lh9B8WZ1WKllG3jxuSl
sDi2D+zAx7v314I9mI7CEUtCD0hmA4LfYsiShKgX1CRVPFuafnTaGGDtMPRv6Q67
i4t/oT8do54CixRjqxgjhctd+vraCyeAjthF/yl+/01v8fyxoLk2pIQjqcmG3uSa
/hWgdF1HEZfy9oBmh2HTAtM1JmCP1TB2zlOX9gHh8O1Z8QH8RPJzQDswsRHdevG5
GdZjXkLdNI2eDCSqS6OGErXMOJ2bdzQpkhn2WEyJcDUvuqjvRKcHE85ED1JHIU8H
UlpiPrdsd0OHTM981njO0cWwpgju6G0tDahSnZTrgZEyWd6yO87FwuU8Xnq/o7SL
cE4RnagggLf/fT4Qmo2doU4IJL9RzoJwSyWHGOPcdeQbbgMlujxehkDYSx6MJo5s
8fWS116L9Px4azKCgfsrBzszBS+i38qeqY+gXUTXWwC9+uBtRG+dTzbCK2ekCq71
P/pqvavh+d6AwVJose18XwoUScCiq1xmesizVJrbhgqHzWZ7qZIAPXSKriP7GwRh
hbJ6pySF47JitnbWcIi3tz4LTfKfzKS0IiuLyDTwMUePpsNkfxzzndqe7FQGxiYR
lJ9o68lGv3Yu3pZoi6zwgnDjanR/OmLIc8rCYUg8eBVautu6auWNvRpz1hjqZHPb
KBldc7IT7NHKDBHPfWYy91hqFmdkVn6U1dwKNg/kGu3hKXlh36AotJKtx1Y9QulM
dbjVpM558wbOyRXVqEhJxvo4rNFDPUESlID761zKnan5qLyJe4EY7dxbyBih/QRi
roiF1V2KQZJBFywFnP6rTPl+8+M2MY+Y59UE8bA31/7Pkcmx4NZU8pJMGNwI5hhi
vW1wg7La5Uv+ioR40UM05FOABsUWif1fnMYvHOMUyuxXf1NDWIeVRlqX2iPF1nnx
BwRP5A9RmoBFpBX/tWBIvvka5JvDkv4A4fFTOVAKBteZ005IpwZBZZ9QQ93R2tP2
9oEomGcZvko4ZHF6RFIq8xyjvB0zcxWJbdr81H4yVIqdHcyC6tjV7yJpIEFart0U
YRf7O6tlhv3tqA9MYHnhsYS8XH5/jEBc4QLev1aR3LfXd9AEBMHrBghD90LC5wNb
JUVgUMmex9Pgh440OcRjhDsw+KC5xs2APBU1pxHjEZ67lS0fIbwbIFdjOtnHccQR
v+DWNWDbUb1IhU/sdqO7K0J/Hif3olHIWEb+9Qt7JXdiW6eu4iwrBZtQYS4DjaeW
tk5J8RoJT3KcKMbJ+lnoYx9k8sT7C/r7fwN4C28oWR28Km1bhpPLp72giez5nPs7
BjSh6oo2brgIzFS1uLt7EdaJTcw6so0/So1tUnqOp/7lvnC6Ilsv1xDyCuqf+Hf6
LsmhCk00ZjTHgkLj+c3S9CE6Ib3xfLbw4Bgy/5tvNvi5egm5yrIKoMFNPtxjAb+d
DaSOQ6lCm7r5kx8weDFS8EOMfp3mJTfCVdRo76phCVK93zMltGyqxskWUcpmh4xx
Zo/fjtUUsEbP1w2zLZ0qlDL4sIqVOQi9ikZoYh2tufeqSzMzlcskfs4UvwLEEsyu
BkyVYwm1wD77chFlsAhwVmA0ND352dRkmc1pdGBn6rrTBlbmnkVuGwDaqPg6AOrK
JuQBnifYGlO+xRJAucksQeXdkP61Qv2OMFcSjSFbIFdA1dF42AUeCJRtnKbssoV6
/94+kD9yqZce5svkDFWDMPTw07DTCc9H/S7VCVazPWLIFvEafEzn4lTVQr/0uxKc
AyNotCo1etgc+0wEFqUX1M2Dn6kzIlH6EenzcAH167NKonl9BKR2CmVafFKljTfV
UrZrTgr34rbXwZzjKYe20WPI1q5EanNJJ1pbn36dbwbNvIjn65JzlvdXVxHPwF8e
deJMWjwHyPey1IYlPNN8foVYaD/+uOAjT3sI605MyPuY3JB+0zHVlgGu057OIUM4
c5farpoVaMolORGmx57bwfQITQS0+OarjjB1MtahxWzd9GzIckrC2mf8qH0G2uNh
wzrhx6kxcQwnvTD+LIfdfj8zlIxiF6i7N3O9puQ2bgvwKtZHX+PVlXGXDkj2SKZY
SUjtsEsTKvsJjUnydMYh4ofnvUCE+UuXX9NtFhhP0aLBfJQVkiQlroAiIEJ0kyor
ULZsDB07hwIJc+HR7YUtlgmQStjLdf0gsccgcyq5aTedFQU4bOUR39Q89XjK7ToZ
cuHH0FNxCGF0XxcSCrBu8n30yUBzIAH+7gJxHCMJ1R2uOG+8a89bAGx22mK28mIF
nmxL11U+VhawTo6aVE+YtVXqpPVXvrqCYXHpp7DWOFLFKywf48H1YcMCQVvfKQ6b
StJkgjHmxokauurIhPpG0IgoMgKoXSnqM9+WM6U1bkziD8OhJibegO6bZFaOVddH
N79k+bqlC4JWvOONtjVdRcG2ZMJKHXoLvnsqHaGEeDjis2g4TZUWo5mVpgQJkV/k
lSiGaLH2koz9Lxi0mfshAinMpSGbdJGRYb7Bes2KWvgY2a+u3XZQ50BXEVD/63q0
BxPgxvePaIelcQOmjTg/nmrew/r0UfaB45ddW5HS3eOz/7Sm7AwYoK2ap96Vu1e2
P5P0zBeJeyxd110fTye8aQqi5w7hkffWHj/W+gjm4sVIZ9wHWjvVgki2FiX+d0Tu
GCV7ZLjaS1oDK+V9G9Zg+O2odQeyR9XnUzibj8DaWV9KKqjp42lRqcjSpysuCDvO
rmgKRKiRa+iR9PELcDlcxc3092uqQqXfFZDQEPWJz9jD/nxXNlCSf/i/MfltcQIw
9qfpvKwqsibfUOi51muJVnDaORN2ZAKal1S/tb2LdTtLu2SQVWxfyQ+3wnSheP2I
T3af7x8cXnE6YCeq0Fb1l2oJ/sjUg66JiDeKRcH9dxw4J5SuvdEkKzt7NVyYgXc4
3QsyIS594xCfOwJaGyCHsLYvzooGo7qujZvLt6smInDA/yGxk5oe6pJ4LbEJUiaY
l2Wv5acXsMVbVrcDzRy7oqawq1VGFoS13PCGsA/479NM54bJPgYfk4qS+h5/xWYn
D66PuNHMGlXhvmPOY2igfZz5wEgLeEV2Wodh4ZIQaCzEHuH5j6ccCK31tCX+l20n
rOmgJFH/sgZASonKBUSL+7CTWpbeEuAjFToZpxIrkqmG8RYrVA19JmGTnof2yFaG
TJngJuPEGA43Qn0P3uIEYsS/FGwdVNHveL4rdTguEkVQOYthXmqKzVbaXkXxCnr6
t6wdnbRO06Jwe1wsdNurPKLvKTne0J89eiMkVCJM3YzIF62NUVoBNdgQ8Dcj3+xX
d++moZEWTsDt/14qbDReqgNepmDQpa6cL01e07uyqDDynYs6GrJ0jeeg8vRv2ryb
h9ExEMv+LCI8+qFr2Pa1sEuF+JkII07+wqkajkjRX3hAPkOuaVy3DOBb7cu5EC34
ac5IKUBptOwlQKjURv4SGHWNvcnth6U0revjCYwDyX74+sJzFzFt38C4uaqSW2eD
hcFHMcjxaHETXZ2PfjYby06hJRtof07J4ll0vMg27I48cZrkJ0+HvBk/MGDQL6/v
Jj+/vvUQV6YwQDxNhQVgT91n5krN01TalHcluWVyCrU1+uhCkr7Qkfk78220rlql
D0UopSQ2Nou0zPT5VZkukh9lUI3nIhAuUawQ4lAdC9hS0oDXtk2iRXBaB7/EKUZ2
VkxATeNJxz9DDlq0KS+SnDmradBJF4lw9V+/dTris1HYSyqw1M8Uv4VDiO2fgs4v
xPr7zT9uDvNLFLQ04mTArlOXtbD0ZcUsZj0OJ60GerEERtvHxRpM6Ar5ARGAeoVY
U5ROzm8r+EIhxNDxPvpfqvSzVHA23x0npCKIuCDgeg3MgCUxlVIWoq55o2vvpbs6
9sRbUP81o3YjEYQO6p7DVe7feYk+uD4rCc4328jExqWEv0FBZ6wPXJIpgN1kUcRN
3rpQR89IY7mCMut5G5tRNU2BVjk8fC5Fs7L/CwZfY7AbHIAYd0gCojKgxY+M9POY
BsSdyFdgFpzzoK9APOvvbziKI0AuGoc5A2gfan7T3+XqmSryn23iQobpO9dgNNVm
9OVZgcXa1vmAX957t+51c9X3wMFCHgVkl9ZFEcP/hyAgDsWrfUDQiKyKooMxk0nS
1LGpdXevkol+bLA6xK4PlMqKgcDlTvrZ/m8+3D1vMmw3ZU84HBQn6S6n4B38QZ5E
s8gpgILYjybttThFHfdMyhrZyoGxKua6omo2w3jZXMcFk3FdAdhEK22sUlQnjzEy
M7LEAqN2NMa1tWmitVh+V/DdIlvhHqWmmyDZDYnQtKMYrx02OBnR1jdr7+mTLP5j
UXXksMuBuifpMsH4OQvVEFR2Bt/L0EwJ7EjGyFr/XFy24lmUKHDzFivZeXxxHW8g
HnYxHe0ZfLDoeKqF52kMx3a+6yBwt8iw5ltTkOeLDACyVlx0UnhDL+0KLJPZvhuu
lOdFN6KYdu1Nd3NynoJvMfyZ91ZhaST3coQUcoaDEf11CxToD4qXQRRNG5i3ERCm
iaMEliigkVwCiVArz/fClazRd+SYZfifyAVUfdyexLunMjwp1w596PFLX5fJ61my
3prz6+w9TVpR9J/9ytRLUZUEw8U0ADGQRIcgbTOcD8E/l63jvJsohjPAV2GkbSuO
gJrVCCIMWLgqiS5Lxh/lC8rgIv5HyaonlFYgJMbZug8j1VVF9TQUe0RLI64m05WB
wHQtnUNOmSvP/6mF1KJVtJWWlngnNGyLEHhqDT7AmSNIYyP4p71zbIasxvveparI
wzbMtxtTeg3EyllbfOaiFr1E0Pg74UKReO+qcKz5eSUGY5tyjhAxnSv8UmxtDul3
A2IRU+4puA/Q+LcTHqFIvr1KGRZkVNKAEQdmJdspONf3rQ5Qkvpi1M4c8NbOp1zc
HSMcFGogSPY/1X5MO5GYY5eehK7cEkr0CDNJNcM8pb5eEfFaaQrI3l1R6hZEcht0
msQ4G3iVvJZ8a015luq74hPuHeoX+HZO33y1j924z54ZMn8z4Phu3e5R9MGBhUf+
BtysMouRDlexDDpvhBhpAYvZVWu50VZY/hbZnqynYxCuAwXxqUfsEAk/JgVBqP9n
U6Fc7tw2H90KSIDF6Dk0QXDi4zq9yMuWBA1Etk3I6apAGrsYGErAZOzlS84U7lyQ
2dj9hv0RS/1/gK/dW3C5ipGrdrxCv3qmSn8iOG13SAxgNyENeHKEnfZm02bdSplD
9gSiSZ3HFzShIqlaujCga8T+yUc36PW4FNkc56IMHPnS+7g2AnEE0Ztmuj5TuRMb
ftg+yJtAV/9vQYfVIUinNl8yqyXQEkTowHViHbvvhxKa5orC3ErjpTDZMT9mHchS
McnXu0il7GsvL/vf+xBpzfb/n780gWaTGTTDXjUxPD3uuERDL2TeRQqPANSCBjyy
QHUEWDxJUBibE70teXmJX2+E9oGQlcMqjE53ynrjM0l9AbGu3zmOYvUS6ZpMd0Uo
7EK4Dy+vT92bcR+YiI1/UfsiVQelEG0LeDSQaEovFshkpJD0WCP7fNtE9U3z1Sv+
GXebBL+X7YUUYp9IL8qsjXVl6dfthcXTDk9/ekzbhhuiHaID6sq2n3Y38fIyGurv
6SdW980lFT4hxCVU1MGBbS2t6dslXvi50o/9Z8ZVbQr14O8BSh9MIarX7iTpn7zL
lM9scv6+OY+IWUkQE/fiT/2VfKvMhzsB+bkWmf285/j/BfMemF9b3H7vKNw41iNk
zfbPve0SKlWpqthUjdmZI8s5J4UL+demwsoMXf+7a0wq0+pRU8hUAICPHG78p9RI
lDaUN97nBdkL0KwyQiabJ5IkENwlLvlM2EU1APgxCFmS+Lxc0+2u6+ROdrIBJLea
vJWeEMUBIUF+MSCz+2Twv5lfPtwd4tRRFAxjES+1Dyafg4akFN8zw/9XPOXV1KRM
8nh4YbsVXEfuSJ/cJt5hCn7dqms0tjejLBNLOU50q+jOa2JozjvGa/DVZuasvn4y
XopY/UAi9MU6mM4HHQifSkCaOzSBygo2Hm5xQLL5Pjrp+KH1FEG7ppWNjumIEpv8
tmFm68gVWbeQclBevoIt9F/bRbG7sA9Xmt9XBZeBATrDFdBv1XRFzUQ+PkJLBwzc
GyPG/YVxYb1o3L4M9umj/AxqjkwUgcfFyrCMNFGkMXSgdvfFOcGjWzoRjHqw3off
3z7yHSd7MylWsZs/VFSZZ3cd0XorockzIfozxSqQ7IvJeSeIaf4r+J2aniHPoSrz
nbfTJpLqp6RElPLlZqIuutRydO+8wp2WV3u3XarEjlv4yT6ffngTFeougjQhp05m
wjkA08MUWC4bE2M6urMLJu0uoRDDai5M3JOoE40BFIxUIWLwAn6XiDZZuX+7pa1v
lMb6kjyaIuzNsHYzP35r4ztp9l2DqHnc9WmAcaGUOmh7B9ZUfHaH9zNW0oY8w/52
DRBD6oYITPja597ECcMAU2MAHnndJdnKApImYQULBpUKwxBEksyM7yUrlWJJxKQv
LyR8+5PxQyyhI+EXR377SH7sU2FRK460twsTcsqW4NORHhAOEC8dUzb3BXLefDPS
jMdiuPVe7hnSh6uLYicDMr6ed7yQrQ+t0joBqV+HTuJMxoHSyMGgQ2Ww5rxoah1d
SWKrjgXPsx5WL3SJTEqtBTouzK5zZpH0LfWJFysNyBRNYJK8AlsWQvUR6FOdU3ec
cysdca8SZYH+ROCPvRmBZdNCNLoDlTBXThXqpUeVJOq0L2C2TbjUrXupMHNxhrI1
T7SyhPlR28L7NtWcXZMw8Y4l6LkGpiD9y80Kgbl427MzI213z5bC4Pdyq14vTlvb
gfaWynwu1HbozhrsEWrVKISxm3rjroTqpXjlUh+XE2BHWGqjh+s0XB01LJ8lW8Xc
wXMUs8MHPaqxreEnxOwlgbA3RLvsi67HdjtitVOcPuLo1ESbeu/KFZ2Rby2cVFsJ
oC2ALkQNAm38cQO51C5lLqp+XNh1ewo0Hl4TQ+3fU+J2/67feifV2YxnLfJevr2J
k88PI++gjh2P0tJWjpuh2acbB3HfIwu3al/eG2TQnWH8hDFFCv9sU9xwJV1augSn
NtroGLQO+lxPjmzSTs6KnJ4W+bv46NLNBRn5sfTLkTE0s8/dnZ+iGz0aI0hiRS86
rk5EYYCt47I3857bIERfrrcnXGGCG9diIHGsQwlDZcq8XdvdTUQSn9H9XdEaFrCE
+aBd4vlJtuDe0IIEY0G7gSRwqLKTb22Ne1hp4qTaKFVuC2AojLaO7KkdoRfLJECL
Elo5WKZ0xhcRjgf3vyQA3ASp0sb1XD1sQPvSgOonZ2Qo+5eHMW5Hz94vTkkwzvmI
NzqowcFYKvc9XXJHJCJIqpPFhClR14hoayy67Y5aSBfDn8PsjVho74AMTJsNb6nG
+OVgTbgosCIB+408gQ2L3M+U19EBkPE39CZ31OmcqYTcz4Jlq+zoblp/a8+2bRho
we/Di2shB40Nsxd5BlemY1rSk0JbprOCCf/9Ee85K/Zk0lf6u8VuCY91u8bgGt9/
LuDQovyZRo+qjI4H0irkGNCe8xOdiytuiKmFedqeM09ROs6oj9wsyEscKI3/aCw9
vxKfj11LUMnxn+xE4QApAX43wC8OM4/Dmhy4M00EJjeChack5mukZ92H8tEPT8Pa
1Z7PPx5UQa4nZGxHHLpeLbro3hWXRLi//nRZg52q/EF7oW3HX2RDGnOsu2vmN9Wm
IY5hAJ09SvM0qoky+UkSIGxyG6IOaIhcuih0DLpx5FSFie7J06zZSPvBJ5IsPewt
dGMdhZJ85++51RDe4mKBJsJGUJ2uUkTFUcjDoaMWU9lrQmEX4o+iKI1bnIFOBCGn
PUvrivz2XK0HdZheXiDa4Kcr4ucLxor5l1tMlVzvn4KoJSTwzPQaoAt6bizlryHD
bRaUDKasVqORKyhK/6pywLNf1BJT2z8LxbgFSs6O+bibMwW6lA0tMOUG6XRmBgTZ
M956+EOHQQ8T6phCEDgheOFWy2fGK/e0l6NCVn+JC9/w1LfkJhAvSBMCloSy6KWD
94n9eB8OZAQhhhou+GCmpHzFH0j+/P8qncbR7JSxjpC9oBR6+9cmytUBbcg1qS/e
AHtu81o1UtCxPqCaONtgSalBdHtQhQG+eeviAItLVw+Ejxrl3KxV0zR1DRYVQOWD
lgl3Y3MyZuZmJVE7VADb1cFS+W9K1X7fA9pkktwfYGDV6jV/CZP87mXKuvcPvwk0
ZeLBouUUXSAJVyyzToDWu4mfDnY1bkY7PIdHCHzz8JbVILJMKwXM60PMpNtZaL4u
LJbGkRKv45MRa3MMG6vKl6x5LVB8G94Je9Us/bF8t2L7u2RI86KI1bIAGwyQzIxe
4VhiAE1sLKihowPnxHcy755N6O8Dt0WKBEj81DgdG231NwRvloH/f8fKCFsgVEF4
SosQZd/44zEuldC3J1W4YmVWc0uy74xv659B+ZB3saMsZTyLVhuIboEIjo8YiKg7
xhLRAZDb8me7hx+mDrKDPpnpN48WDfbqsrXMF+gjXPjHwuaBhOYUWUq4s2vLZ/mA
t1u0RGeXNYJ/9DRIV+Qnu2nN4vXyHgXuoUgS0q+69Y9uZbSfps96Ja3jL8iga4hp
9aycL9GzkqKFvnjkPnKh6d27jEwzHFZBh0hENe6TdUIdQGLCksdoXCCPBtmljqnq
r9dfuVwFrYwCDtfwB14u/9O+b5Qxeof+HtG4aZQ7cfTThrRHQBI9AJtLoPgiiEVA
Lwt8RaaJYb0NSzcI4FlNSkZPvnq/yKT/sF6VUKaMGCLu0vcioy8RgheSJzTXZGoB
hT0WPBXKJd2nvZoLWf3ARcgr/KtLaHcI5RGsHCssta0r9Jzpyet9eIls+sNwq/sL
3w1fgFXU5ZSWWmGcen6FYm2kDUACpzdQ4zZKC6WGThqE9b4WsmPUxMkJ/I7grlYL
AaH5+SSD+r+91qiVlII6iy6KBUcCmwz9MqNFGYhhnV2V5u7ahTl4SfIHrDCtg1Uz
tV5KDvkrHdNVqFyJdIXzLEueCEn+RNuMSewJ6y4/AH/pwrl8KYrNhBOkdBeiuvKA
4izESUe0tJuOTKCFgJt7SbsCGvhAt7pCcjVuy79tukwNL+OXHIT1v1wpHKFAPhi3
TkaLJIxx0Oa8W3Gst1HcXYxJpKRMjH47lQKAmnozflTzRArzEJMCArr0Atw4sMof
Ykbxpq+tH6rbaZGj4rL8ZuGEInpGgpXgf95e7Mj6yshA19ZiGNFDbo/pfA5eixXo
Q28n2tPM/+rdqUjtpsDzu2avh1aZtBuElmZyWYHGTa5vnxF19LOgt9SXQ4KFyM+t
iLxQg5veofG9B0JNjITUgqtgJSHJOBq7qpytCbA4pS6NF4sduVj3oLZ+TJzDWkJ/
O+I3CkXqz3kV0yDGqE2lfec51Ora/NccDoZ3BUsi7pOYpYsl2rwTUXaM1oguMxg7
liZWRZhrmMn1UWNgBr4wMSBrY4B6pw5nicVFwtyVn4565uKpU3wZhcvpyuJsmhof
xR1VlrIshMTaH1uf/GxUrFcyK6cUp5SqU0hK3Am6cAzMbY+wy2UApnKsEQO7Vq+k
AQUqQZILhIcO9RzC4FgZMbLrEKOj8Q2ySgtFNiY/7hYDyFoYa8eHd+MYY3tc6hgP
eg7C9fKyd0REgv0NslouBaFrKmK4l56g8IGimdXHcfPDvLuSs7FIv/piCJl4lOi3
81qxoHlnGRnQ/w5qXJJbpqTzCG6l7dUSSmakk543U+JC8bLdrgBTAwBsD0Cb8Nza
GiMPRp5eIMLBo1m5zTQKLRS9MqWafHoM/wDxXRGdn7BPOJQ6d0D7Pz5YuciXPbdU
6ommdsCbWqTLQ1ezqDxL6gZLs3nMHpuJKwOG33ERL5fdXjiWjcPefaZxqTn01iQe
n9NCB+kqYZf04pCX2mGIZPuvz0ujIkW4vy1JMqcMrhMxGoDj6I0unEiAo6W/Na2g
X44RQ5uzeTH0ilix6zYXvEEAbU7XOtsELb9RoxHpRXdTkT70GEibRJQ0F0p67SSx
17cu636fPEfF1sWUFr48Nd8qrNAxIteRrj7MQpllmDW2yO0QU2rsj763wP0he45a
k8sDrIDjQwxgGkXpcYUdErYf297I7F0Saz3aNBSwwBuMPpPOza1K+Fssavwe34qB
udjdeoN2elpkrmte1g9YHUbE83M7Vb9ZcB8tmQXEP0dxxsepmiQWU3qshcfZj/Wv
/G6bUZzp4S63OeAJ3Djx4PjXfXiiuEOgC/UlA+gDqtzBibmssrnNnX9bE3/vJcXT
B5VQQpCfhRF2eeOpzuQgn/SGuMyLE39x4SNLaYmXoy8hQdOLihF0pNr+shRbcdQS
MwHXZ/42zzong7HYr3bEWuiIiTP/iCDQipfeFePaObsPzXSlXnoFb8tTxvWQ1uM0
gDk8lkTamgcS9ZNS2aUM64SDPDOMjZeD9iLLph8hx+2Xa382Q/0EP41rXFKc6oh/
n1THRbXa5mOHgKyND5blVZCtIFiadQ0SPg/1ih+d2XC4H6HnXZvmb6JYC6mS3Jme
DWUO+3vmSJXPT6T6HdliN2GJ2kIJHnOSurrRMvsYnmrIB0LneYmaRuOcAcSHy9D9
qh34LY2lEOdU2aBt9s0molamshjdTpTGMmNDSBMdIMWkzW5RWUh9a3dBt0cSiatG
vBL57EUlzEYzyBShKvmgl2rRKKXN2++P6vG1VO5I5KmlZWuaBXzgjilsqGv3Ba5W
WqlhjLxEHyisVr96ybkD5jeEC1TbbH5jcB1rNG4umoQnFdIK90enUGFu1S5B7BC5
ZCwkW3sG5cjl0PxmCt6WjGY2027RPVCTacGEf8oo7kTOlRQ2cM6dRIxe1hv/LojK
p9FeBj2aDDsNtBmqhwkfYjBlccM/QNEToNwdwHP1voUsmfhJSirSIwMNdIg8XKco
aOyvjmoXzHzApiEzxp5ycz17YnRjbbKAhLbWE1dID3cFZBvbb6JfpgoDyAGY9iys
T07xkSojms86brvFBaXRfwqvJfQZOtm7q3YLlht9/auujVxojnLXgnIkao7b+CB5
G9cmLhbtuInf5Oank0sgARhXgHEaaVFww9FnGP11zNbUEB6+dhBtwIdyQ48/6fie
bcInkpFcstfKoPVWIm5MlsIU/y4qheJkxJbM8B3jWw8W5+7YYeB6F9lLCUomB0jq
VgF52Iu5kZ+VzglwnAz2ZIZzJL+kzmC3Q0uaXpDtAHeOa9541SmyQa1uPFYOJEnz
Juhfg2y+Dp+T4DooxZBLusHkkFBDeEQBkpiRuYCFcOrYBhsvnn2GoaFS0xEJVrK9
cQ3Mijb07ZnSQc0+cjBv/Gvp1rv2hhPL/njgTGa/5MeCdwwJQReuYYPQMVV2gwP2
gWk2yPWg75LdnMjH5NUxo6+r+fySuqGfwp/T23/IdGxtHMeEoPrr+0wf8EoaJrI4
gOWJ/SIePinBS8cbmzZ5NDP3uCPAyEEFMjpbHdD7p7W2vljwJFKdU5Zmf2OJPvgV
N0agN1B1NBdVDkwrAW9v3IMsaMGN3oqhgPL0MVoB3FOg38OtZuy1UvFHW/P9Y9eD
ygiyBktv3Z56iQhfaqZamouKNpIckKR7yZgijWwg0CFvvEiOPxLkhXwu4oB8ZRe/
P6eeeL5kp5fugUbgV0jQ4bDK9mGzXIAx9clNMb8mtClfTQqF6u+Dc2aHOvvQDAxH
f86zCpEZwPpXAqaitmMVGbIlsemYwHRzWgKrO8XmHI+VzTadgi9cNfMHHkbuGzTb
pzdRzzTqtZHQ5nqQawvFy7R83lSxrxYSPc6eS5oP5sc5KGdVt+w8veo6uvXysoOY
FSnh9svQRlmUCk4tjVx9zQQG/TuDxQjHOD9kecV+FnsVlUFGxTc1eonFaZYvkeZz
4i3TQgkgd767AqKPP5jZfAS2OHVc62asINEpXFeL7nAk/iWMJW/vDCd8OvBMKTPu
VrflRgxery0AvG41KMFC85sjprCF0GLt+wUqhQ69iqgPWFh/YyfcnQHNc3I7h7QR
1M0NuZU4v603nn0hGUmWyfxPtmx8TQnVbc0lxJE+82VR7W90BMdQO/RorHs2qzWW
IL+RhilVU/WFJcxWd8wdvwGgtvrOuvgW8jJDZQPGXLcwahWTuPRdoUtbEjGP/y77
tT+gtp+k7KuAImkUKGhC8IHgJ30nRECuC26W8LoSMlT4SH7B8+vrbri0Y904ydav
TfQ/9Nt169cCFnIkmwTNM/+U7I4UwRkNkKD0JZ2hQIuRKyYmIMeeXbJ451Aqz/E5
JnlLYjf0tWKh6D+JgVhSUZSsGk7aNfKNNXKjZ+nleHvOWv2t+3+pXHeH0RKWBECM
nU4pNqvXWir6L2kcWvXuLVQXHllkv2JLvx60b0QF7s56m99eqKVPZmUnXVeQ00hS
LJTRRmGy845f9RFYr0VtfXXwedXW/MmRFz5p23lW0rWGIDRlIdlcXzR+f0YD/yrK
7ZlGX09wMRXWz6/tRzsg6WuXkx9214C1m3fPe7i9ZD91MjxRGOmqy3/mmf9rymFH
B4j1E2cy96x7kD+uqlkoW3mc0A3T7I9H25wqFV0SnxZYPYVWEBFi5ncHCGwunMuF
awTXZnvAeIkiOnZsftaY0Fn9o0PPKEZSBRORz3B/WDpqVJ5QPFE2vhKDA2TnjItS
biYkxt8ENrUAP8OYdx+BOl5WCIKnF9zexEd8ZT05XVGnsE6/S2/leZrHLo3AXG6u
Yr+7OJN2ulR4q/KfvofCRthmS3gOTQdPX1gAYNHXowtvs/oCoNmc1TFLVOj43efS
DX46u8ib5oc+Tw9XCrtbWht9JhlzN0oBKkeMBAv0WaRboMqZulDY0awSSREReweE
AlPCLUj+j5z31LkXqcp/V7GZ4bGVoTVmJHaO+NY7nD2lzB1kCzd8ASNjm3/BOomz
KyrsSygN5SvB4sR/kTlqdVVyrc0vgSpuC7c2g6lNfFqC1eueBb9tB58jetnE6P6b
G72gtjv1aRu4sPsVTHEL1tVJ41eKMRdvySZK7DnEiPoXrKf/OFEJwKhov+8w4WHZ
mLWSLB45TBzb8zkmxMjYckr6ix6L0CUYreIoRm/O+Q5Oek9LtSwLovYAHwJKdgLm
/CAs/XpUmK9wbR9L0X5hIv6FOO8zX2chAiVidJ9V9UmPr8e3DgbBXM/ndPO1mTXo
FR1SV6+6ZK81t6CSMtYlPQmZxA3NJEgyk0Wv+TgYCHojEh9JkBOFOQp7ZiBVd66f
fRvZndIUrlRts4j2luZQ5E3+zzE4qbEYiDE101IR0Yj+c5THBP3ls++2Z/gSkwLh
D0V+L9nCjtqmZcSa68MUsw+pQKcVgyaFnQKpye7TdFcnPBrw2OycMb6v2cY90A4z
Ve9gx5Pgpk0bIlwnERAh/2B126I6tEUPZnGBdx+S5dYkGVp+RuODrC+OH+boXBy2
EPBsd0RHtva16WsA38zKzJJl6aOpnZMIKoTndSqs5+DpCMDGreflBqpMAmRyA5GP
UOGsNlbdRZK/TMH9lC8EAg5xV4v/g8TNrD3QhO5RJRqKcWjEwM8rRoG6MzBWoG2H
ni+5KUFJBGqA+1qszfwRI4nuROBagp3XfVKtrgn3KYYyVGYqYpSBn1TBQiM3W1xL
sYAy1geHinKoiLaepEmaI1FHsKWu0vKT9NJtfop/g5ZwhTlQuoRMHGx1z+Olguli
f+bdwcTdgbvyDUiyaVJ592KMKu/VhbWWwTyvhYVQwLGQ68Lqs6sHvwGuEQmP1TnB
33WTpj25hhG7+0NCbz8l8xRPOY732uvM++rk7Z5xd71AmLNPvhOHbXxwQKLfNAtY
9v2TREnIFuGjMXHlVmEb7+i2QjsKzgIFK+2Gk0BDEF0Qnna8+BWBdbj7/UV2y3qJ
XyfETXp6MmxidsXhSS68CSEw01i6FecvfE+6wci7aBeIXj+Y6B/qlBsffZFcGwls
b7EI7z0cJiBYnY3H4DWckSfxzIOvBNY/mnuy6D1XmTFxeyjwWfL87CGZP3gBWKI7
9tz/T04JxJ+a8/tCF8SE3BYYsqEJdtYFiR/Bj10aC//13CkOqHkSWIRkCfLJ9dHG
rlP5vTG//tAM8LxqmgWiqkHvIx2s4i+MBU44LM8ehrYQeqnn/pzVQAPzipOoDT1P
5O7DeAl6Y1IPKQKeoRsw7MHq9jVUW7WuR9egIxEf9Rtf3gnHpdOCNN1X7dS9sdOP
iC70DaxdIaNfr9nx50zetOb0yk/qjV0ce/LbxlUC3eGsbqv2x5Ny9Qk17WevJ85u
TMADgGUHKKTF6U0WLzLfB3jssp5JawUY3J6LY6Y8/3QXju3FMVuGT0RZzLkRZ0iX
OgIxZvLRD5mSbMzycwhIm5+hS7KiGS4wNxsKcQET5VRssfvSbJl4bLnZTTMYlERY
tRP6DNl+8A9kZrtc9sf7f3xKcb1F9Vyaef+4Vq5wNBlMyNVGDJd+wnnaoPUs56n4
M6op6IXAToFAG3gBVameelwuekt1jlzeTjn4goJ0gRCmqRATM7Eyc5RjoisP7RUx
yK2HlR+6ywZxTWHfjr6KK4gFt1U8XPZ7jckDnDPmvt/zMYTvt4poUcIBlBm1sIaE
Klhr3FpnWpwTAfOrNf92HZnqzL06tgaaqIvPCvR8x2CK+iZGiCNSf4JeImO1iRoW
Ce1Q4B+274eA7yEYzo8tJpfIE/ldHuofxYBXboN790qfMLHq6alNvoyFLqu1ZEBc
nXacZl3Om//qdkcvjTb78+MfpVKM50WxysFkZ9lpJEnF9uWvKSmbOYsPi3lHbTMt
37UhaLVZjShkOnEzPqwajMbfhcYLIp8CgiY4b829DTeNAmg3ALm5VvAwBFZtnV9u
0Hm49+dvmOj+pE2eu4XmSC7DBNUP5FJBihp6C15CzLeNULyBIDj2DkSt/PdpsdE5
qfzfOS4RpRl/vVGT2jobQKI8hPan0WP87AbrGmvHa6jafhAMyvGwjECzK+90xXBu
Co8BcLOXxVBU0xzcUvT7D6ovp04ypp/17JHZd7DDKdrM8WddiZapsJjNKIL5tMAn
PcCGeClPeFMhZULz3+lNmPlcO49x0GxPDBvLFdsk5mrn9oYw3MEcMwn4Y1t0es3+
pBWs7IG+eo69MBRC+83kbbOZ67TrkkfmNMCCtDUnWJ0GM9dBHifLLyvITC6X54e+
YoxPls2G33OWqnBvf96t38I3A1BReHlCXjexPpEvxSojxuFNoQx1F/Nkvx9WFKZJ
qT83J/VPL2UlYZoRrdjwqyO0sK6WAGklxxZ+UqassGy/o/NO6PCE3HxZjkZMLKW4
snGexUqJahWewxzKb3H2f95l1ZABdyZDBi0C5T4dYCVFNl0ZKiQr2jA9dqQnd46G
SUkvhmlYoUECSlXvQ4330a+DeuFWqtRBWAjDXwirAsBpcZAweWQMjoS9f95i1bSn
wW2O+2BMZdGt5v7Ch9PVU7k3RSLq+09rAFJqCRaS3qU8wk0lCt4QXkm3/ekGb4kU
eg/xihJGL+1jzH0cOjN/A0Q0iYORfqsCYCXTFWzBUEDZtCFja+S53yb+8ZhkisGV
xob2mtLwcV+xeIDhgaLz05pEB9gfclgnDHEq4wFSueM/BN8Oc74CBfc7XNvl4dtP
L0O0G9IYUaP1ha21cSdUW62Frbl/uteuKLuL3BcYzleNtRgBLHdPYJPoUNUGxXL1
hqvh8+fz0c1vCNgo1qSnvzIAGuhz2UkDPxNQRRhTv/VZt3Le+5DQyRw6m2ri4oxD
MQ5l/bPeKJa4XqLDfX5/BoxTFhtpRCEqa+tN5qX41avl/SYh+eWjkSdkafG75Cq8
zdIjVzqLgqwJskang3ZO5FW8m2FTRg9epb93NOJrmhQMAat2opweSPEa23w6FPtu
36lpxXh6M+DX/gYJ6QGHDK9zx7rZEniyS3eNexA1NWHNEf2SXEyDKxVhI6zYOieU
WJgjca1WdwtpTWuMN1hSdhlg9ZXr1RtRhy5D3PsGbne9AVGzgGtmf/7ftrbvTZdG
bdrqvKdespCRDOSUWqL7N8cZiqbOpmM7bSqNxdFm9YbD04TRMtqbCyBWB/lbDTqv
rqlZMdU1+9ZXznnWZm4KxC3yOjiL68VWVDh+QIg73/3Js/CA1EvXgi/is9sCAhY5
+XYUDaw4NodBRWFNCI0Jo+x7WjcKyv/HqphHElL2xm/LiVCoxFeqhsWvtHa4/Llq
JzUzrp4AjBsTBL6AGODHTwum/YMC/Hcie+YcM3TjxrBYSa8eWsDGnf2DlfOXECvI
i9ZbLhZdaTMsk8tU4rw5O8J1D1Jw7LVtFISXCpKmdcU36569ZXCzwQorIfrwfEhN
G+zuXbhfDTYj9X1Pq6uUkl0SRMgk+kGPHAAfELdWGoPUWUVJ84Y3PPDHBX+V21mq
aQkLAtpUscFCgxmOW//YuCIk83CDcq+NQTbqejzrC2r3y5g5dqZbcQUVImJIICQb
4Uzr8NBZJVZanFUKA3AmUAPSksecD3Au6q3qrTDYGF5lpEj2TyPqsgqywDvWMaf3
CX7jKb7C7QiFZmSNWaTb7AUvg38NVaHtSPl7+dwNzunwpg7UiqxqhgjV3MqR7xyF
cHzJM04AfHIT0cqoq3PbaZ1j7yKcbGxb7eXfZTOs/QRpz9Hy4nDihldYZleU5bvM
cKQKIRrNN/8q7of57G7/C2zAE50o0dH1V8tDLlSBl1spBf9NIZYsIOqKXUTGqvWj
etIjlwmg6RhPLh42Bdn2gjAqxfqDT5abNSVdKLUNqnCuCtUn0s38qFb8s2atqiB5
ogEEmC0Rc2U1Vd7KUSy47EslDAPXVavimgFSqs79A5tBd1zThDJj1Ky0YLlBq7hu
R1Jf8MJs3kY/Qt5DD8Xf4lfYBVXAxVE4BY8SV8eIbfcfhbBCv6mJ5BSp8vKXL8Ei
fZ8znVHWYLZgs250nDFJHXNkUKkL5HBALn6XHM2Ik0tSDo9yBYA9NWXbEp49Aj7+
t3sNICMpp8YFiAHuk5w7olSO3oVcGVfphLQPtDE7aIiu9Z5rgV8Obz002IR/Rt5W
kyPJK5nB10S/ujQPCgArLcsMhrb+dBsgIQ7qQ9FSD3YR/nqPGllYDU6yMnZMDxRy
X6DlnMEQH1oYsgiUZr33l89/MVcPAxSizWMj7XYu15ebpODiUbxTvY4jqRAr5QQT
BCcUJA/BWnt+iqdSrHIGAqW7hCYxHosgJIMJ8XBY6Xf2VR9iHMepQ3WiONDy5CVn
OVxgxXFmSfDdqpYN7HRai/B4W3lvagcjfRqTPOQExiAvrfzWKfhV/DOWfwACxMdA
7vYBkqmHfvTGnQ01LRwNtYDC01toTGMvDb1QC4713h5U/wzfd1O8JMkM5T1h4y/X
lg1gXB3//ITeb1P2A62MM9i0SKVwhd+vmVhCT2De7lzvTAcNNniDBErNJ7pkHqKp
DB417K89//hctyAJlFuN6r5i7unHHiUJs2i84aIe5rQtTdgwJG7hAW+XXyXwIj9G
0eyGD08GsDq+Kb/1+BRi9l6GCgYEwSDuQhhttL1E85cj5JtIM1gnXnn1YRgmFrha
xN0TXCxsDFZP21EhKViRQUMwvxCVZ6SquUKwaJyDRAAdOIcc2SE5qWoCOo5/AgHT
cCuqBPfKlTG/RMDV3im/7esc9ZX4ZxXqrYdvy7FLVxGcYHpPRSfLTdbhABb3mDDH
C11qE3HdF3JxZdsU6jbWR6oleIR3e1bpXRTOFlE1P3Otpdk/RyldcLW+E1A4u2bv
iZpmcb2f3zMds2QlGSl9YQpIw+qQkXFWNNNJPvj6jMKjte8LC4ZZGL01hh4w+ag2
UfbXf5eO/6Ftr9UT00bwauJbNNsBrUDozrPzovOpQPOH1kA5hV1RSIJf3frug8VE
a+uFFfPwmkqct7yqgzH3toUDGmELTKx+UKhKzc1XdhhJHE67K7MlNCEXT0X+vPVb
6eHLhXZfdqscqcv1HCpPT8YEES+R/bq6MJNrbo4oDti/RM0kEfCNR5UqiZgcJivH
gMOdJAu+f3pEO8NfctwJ4KFJkMS0PhG8bHTM6OzUue0zv4hqMONwOoIsBbcTjkqq
xRX57o4fRAzZMb0GBOTOHWEwHaTAkrzwZB51oY+L8wYreR1NlE8e6tFHXGwi/LZ6
DzI4xCJbsNVGnMqPGjCLJPeuCtkh1WuvCOav81MHxshspg/ph1Wr4Wkayf1Vg79x
SamUZpRcfCn0wH0G6IbS5sBTIeuMmfNCZ8Wks+SapL1GW0eLK0l06+OU0FIZ4YhT
IyYPrek0thPCYdK3E+mx8JWGLvRlm4bWSxAHE2WtYV03hHUURRPVn1sqjD47U5Cg
UcJ9RaK+O5SJY+CO6jgSJHbLB8gVayLf3YM9un/PlW0frS2qq42HhOCc54L7PLbA
l+qwiASKKUXFuz+nriPh/vSFs9gZjh+ufaogBr1RoI1cxOEixYbllP9YnLF3kJf7
gQPusvCLeqEIEmDL/wKn2TN6U2rO3XX7ElzKAoZfuk+sTM8vQsVESSmRXNw0TyzK
XtDI428PCUuwJR0p4p00FwIqkACa1k/LeDzxqLQVT0Fs4V1kT1kCUei3pjBguv74
IJwAYTh63dtFp3Y7nH0hplFQUIP/btkPLucuuPJrdxxoD0ie59ly0GlE0tghvLIA
Hybwwxk08JaDhHpmZwRhhCMJGOZdIU/ulgZgCtwPvRyMljGvggFgBnxiRLb/7C+b
7Zwwls1br8yAsTx1Gpfqp9aFujgnS7oJOjz4YMfyZUrThwehz2wKgQ12EmYRuZ/Z
Pd/0Vzs99u/pUfBaNqvIMFR/mduq+WhwdtnLatdFfHKDS1TfNXnhIEEvCAzwEE7a
shBSI5LldOQ4QXrMfyNKu6f2C2qH0bnmS07AQKdgnWQ3myuy6oxB3lJhLJndMlyW
rSGGk7/RdNqA5cE8MrUGLWFHXXvdTJrhlc4OmXeo99QRUEfYLp/OSsvgCDFwsP/S
VPMhQZ4TUVm9M2SqpdFWayWJnb3oQVs/vrBTu/wQj7ThlcUEnSAbXsPeGj1rORuM
EqZdRWNHeNLvs7o1LxYCTSX7gjpmB5G4hRAtfDGw1VoP8k85XoHZSGyN1wxIYdhE
No2L9FhdlhIdrk6RDQxEEBosbpYdKSvo6+8NVjESFvQ135R2nXO7dZuyplpb31ai
b3IMpYGfJMkPcjsfYfR8TeOL6QdN/3HYrUlDWJDCcGqv9ML8sLJlsHK7iCKJkvn6
6+//PwbIOsANvKafaloo2IUTsE+oZxIhZrLXBzUvASANdhRDmJHoVVEwOhzK+pvN
7dpY4HRr9L1RvBdbaEu4DFVUcZnOG4cVxR3Cq8FptsWrZMd8QR2OsSHOxwBrUUVa
RPRg/CkmfTGp+3c2UzoXewOJIculD/3qIc3p3YRe0iCQ6PpWMcGHzWx1uvwx4iIT
uc7uDf9ywhYUrceisSxgfmCBUsKudVRhfMSm+buLCQtbTMpzthO7QItcZ5nWEZyZ
1CEENQbyE2znorvsAI9ZVYrUwE83y51HTsn533bOaYSfxi31np/QNsWywAuGSK/A
6LbbS2/8C0IlfZMVt3MtNodzFR1ywwM9z6Mtsin3DwDVOeOrEXfh+MeRlM3d/jI+
IvK0fXNKNdQgzc60aEG8SpVT4yWJSd/193K6VEMRkzB6kKcebymOjoyhC+5vTtwM
jTD7V7N3m7PWstpKBQ8SkJXrQ6JxV0wxGZfW+2JfyjYPamc1VlUFpxZyTj86zjG0
9pg9jMLdL5JxhGRcYNT13i+riz0vtsFHMg4xSwtPni14mVVJ3tnwNQ6CdJLWG/nz
2h/zlnUbu+JNHA4AhVez0VVZXSYgdDjsGl6dubEKAxsTeX7oUO74JW5VEU4fq745
Lrl+XgU8cNux7Uxf4pG2RiMSuJsc6dzhktJQrFHjn+CSC8YHTqtL5So51SFS3OAt
vcWHHG8ZONjneOkpnbiwRg28rLkJMhk8C3F8UJgtDfrMzgxsgkVPIdruqGDDY38D
KVf9ZOoDx9bdJKqLQdFKB5Hplhs4lhISmxZbS0q4v9A8bDpj6bbgzjb1zflHP/8u
9GrzSDK+EBjnvNKdY7RaIGLgVaKIHVTi/OkKeg2Cp4yOGttz7ghdET08njxQbRjE
7W+m72PExaTVpfL/ZWMmB59dOhiIwwTLC0M+r56TE2FAMRD6Movhnmp6hl8ydhAv
Kuyt3/ZguvrA3ihkL3TeLSMS9gbNOG+MOKSTGnxnOW91U0YT9u5REnU5s4BKHMsX
j96ECpAQ/5yo0a6aR4xTSJMDughbqNN9KeQ+ilYY23GsH5BBDkP9DOoPl2EgYszZ
kykZ9AZXY8MwK643IV9mGqAS8HzBWjhVgJP1BKH8in0bpFJ1fei4UcVsi4QoKgj9
0IMkLw4ZOJANYauWtqnDdu3hsFeC/+VbGH3RdWBtPWHC5vYfCru83mdPGAYoFLtd
mzQ6w4o/Hee0Q00iolPZiqO/Z6K29XTKg1LVOA8we2xwNLzu3iyXr/HKkkeMv60E
3wCaLymyD/qDA8iHa+ExummLa0OClQbi1yFeDSl/R5pNec5fEb81GtREikFk5O7w
PYYMsBeSoXhXJzrh64Wcm17s+gMf0eAFURDoRQpk0b9u2s5cZaAokmlP3CxecFlx
5J1o5TL46RazWajpTt58PcTCU2NUrHRZuVt0CpI9LrwrMx1N0qGZpa2hd/ey76Jv
nuhU3uQIcMZnasEKzqusSmHBxIio0UDq76dsWkkO2YfWsz+S2KLq8eWpv2QdzfoE
X6FUo65bhRCl+SfzO3h3jpcyuC4JVH8ExKrDpvluEANHEZ/T1uE7RovOWOxPFceM
JEluw4IZLFWJeqFpYFuKX1umtfQhPeoUXxWmS1kW585urYspSfwg6X0Wj9azVJqe
ttvhBb+LbowsJscoILlIiPhq7CoARFvhS1+ktwmK2/u3VH5agCp9Z5AqTxdWgncj
R/e247SO8DN+qzkdn27XtT+lN2hhxcCmKe2u8TZr1CCtQ06YY3cYN9ZP7xFaLxqX
Vqc50oYTDgFr/qAkMIqz1paXBSQ6PskvSecoEFLugNdBecMF47oESyOWSWExSPBk
1rOIbBt6shs7u8Ier57F2QZf1N15D63KFfe/SMGd61hCuiNoaFkgCY9IoZr27Mny
/LRGxEOEpaHHZqBQLOKrm2b4/OIXAu1FdcJddu+5fCQST8vEMySUNYeEjHtHkwtw
xjTblqKR1sgopBSoBzzkneBAMzfiiTn+LzaDRh5wMAA54j6fTKwvS+vDde2tnDLm
v9ivKUZ7MfivGgQL0An77d0LS2w4E9apmfJmIQLP4M/nvEp+tR0OITdlyLrMzoJt
Q1aiLYMlYIQLxgA3/Ahluk/5k+PwNbOPRdHrI3Jd0N8u4P0XkSNiddVrG9zdyUzn
+bk6GppK4b1eGZ1r71fzqYWpQKc5iMauoq54KENJkZyvReHefS8dQo1Hp+Qs3yHA
r8Bp+owt/cBgssnTFnKHPcUn7iuCCl+MaXRhffLsD1sQGlGjiD2j5rBiCpijwk9i
I4UF9EvgZtpq3hvcF/+Ok8YRyEZQznaMVMPlc9F8u4s+NkLFg/8Gf5kdm+gNhaHQ
1Nu9rohZACaWuvcGlail2/Tg1mkEx58xzDX3vLluymtAdGRNE/FwdkV0KuviA1xi
PyYh/h7xbCTBF0qeYXyep/P7NJN5XQJaxFy9TKyHgUbOBpguk5dENSxgc6PzPAeV
q0qT3FE+6ySNQjmaHmkWdaAMW99uUN4jGSzzfFXoec5Y9VeM8nH5loc+IJXVCTIq
MAn5X/m0gq8b3hNpm8QY1nLYjYkBbGciTpq41VHp8wnHScMH3Jc1IDrbtzcYiI84
29YT/xeCTzJ3jdiufkut0kJQhVtKjF98nwsrzwuS5s1YGR7H5HPALGfjUswLmG4T
S11UtsFf0ypR/SKxSzdC2wuw2W9R+4EJ8STTVA8wDtnpsEGrby6FtjjHQPO/DgkC
7igwnYrbzEbgWrmggUYJd4/yyHAaEll+Jo9zNYvnmwJkCbcw0uOQWRd28hIGIPBK
zrlE+3KADdrzuVC60g4xbQrWjy+nGralnrb/uTiCk9d8X4RULbNwIwemI0dfNEx9
UEaRi59myGpI8sibZbH6r25XI63SLYInzqBkUfSB1fFjjwtIWg/BWy25sPoJm+c3
vcNmjmybX5+lkAJBXFsUFq3fbM29CZ3qiLm00v/JJaA5hkDDFME/D4W5lOF7skkQ
Hql5PMVsC3GynQY4GpXQRwhxLk8q+f3MqhFFKBcSH4m/u8mDorC/HFaujdI/wpI+
eZtMmszGUfnXnf+dbytQUie9afWrCV5nJyuYYrmlefKbo9G4/iKbEnf0NJPt55D2
nghO9uRP5gycBAeZtqvfbDx7YW3QESnzVvSODJDn1dBSt8l1XGrVpPL/wvGO4Ekb
T6jTQTNDZnJ/qkc1PWVHaQyWDMiQR8sMvHx+N30Tfo+dxx5VYCzR9ojq/mEsWxUi
Zc4q6om9vn0GIhGGjI0+/PuMUOER5ZvpwYKqEl73HiRVCZMJ4NnWQ/X9b1mHdd1I
Xk6GYcvclyPcaTospYIWI1Mt+e4O4kIvSvNJA0Oc9jsMqMDwIL+ZWgR6PTI95XjA
uVexI3OSjkUX4rcUPBXdqT6QjVHQVOLlCm85+vaWih9b8H7DpqgKPFtV0ovCBp4L
hoKikslKFiO5CO1MnpN6jB9/rlTs3MpGdGEW34irdOYCKmVLy2z7GhNZ+a2tNqXq
N4KHuZ7eTmiZ6vJWQEoWIhJZHYbDNLJHz66Ftu+mCMR3WQUaWs4Q0eWmLwCl+sT6
/FIhzJby7kDK090hPJmY4gqKZZxCfqERKX21MnmsymRyCL2WtjOjUJgDxFdCWL8U
u8qMDaiGMQrp0v8+FZ/8Z4vDQ6ii0RKFl30mpi+hXb6H0oVkXzX+MKUszhlJwlgK
RSU9kFST/e7IX0s1TJQO9lQ5UWlaHpop7k9+93HbLLpX5FCICPhzNNgiUlp5PVq4
9sb+eGzCti4lL4fVTGKsCPz6vBtqNXDYPupH70mETOi27dhK6rC3E10SgTOqQsLz
By2DqPnLbw6nG/YAyRXyGyMAhtB3b4Yn/Ip55qDpDe56SdrY7qEOZs0fo3H6ATsm
sbPVMbwtq9yObitMqbQiWEmXj6xkPFyqHdXnMBxzl2OfZswZM3Z1UsldOrVWqemc
gDYp2dm6D4XqAiiIKyf/1f3153peFiWEHutoakVMMlSrPU70bVU9aml2uHrigBm9
pE3SLRJiTWYa91dqpnjsGj02tCqnyH34jV6Fcqts5V80jHTFZkcJx6/2RgrQjxaE
cSkdyZqSn63ZKH5wBSny1b8B2pPfeWh5i589pGdg383uyQPdGBoZOz8U56rsbIdA
llXvYOyRNR4/8W6OTfRMmDszGaySGF5jaaQeZR6cwPzZV2joQkrvME0pE0MUgqCs
+gRMERiTCoOaNAVPu+jNoxK2cgjZhu1pR+P2WI743cPfQ0EI58ltPnxA5KTcAimO
Ca961wHqUhR3bY4b0pstjhPGNJVOUQfGoPg6yb/Pl/h/UVnBQj7uGeMFfoFf2OqQ
j31uaqX59JthbkdOAcwt8TBlh1rZYl61T9UyeoY/RrZFEVEcXniVUKp6p7dd1ksO
ynz61EBPABNGqEiW5tT8dkVX1vrKVidiEbAYwUFWw0KijVkOY7weg8Zr1VS4p0Wd
jLfw2BglxM5LEqJhOKcTDHSSM1nnLnIH4wKV3Ur+vr8JmHRwAKXwmWXeUrcgPMKb
injoitFU4kjxSea7y3FQDtVy0U8L3nwb+C5V3FhTShhTRMPFwsOt1zaXJVYdf1xa
IaiPMwxiDyaBNXuA8Xu4pfFrQSGZkMzCSb7Wf2tsMCKgLc3bmhxXpG0YSymd27QF
sdGd4UW42/4uuQNMlmuJpsZa81YCqyq2dMzod+whuP5CQBUhlTFiyliBCqXOYaqf
lpJ3Df4DaOTemUJW0BG7X7ajG4PNxTVvalIdBHaMGBfZAz9mpPd9mVKsgNhTGWZk
T67Wy5TwT4GyNNOi0huQt0A+t6C5hVTz0zFjB6m8ATNFEWCpeHHR2F7urOXGmTZG
KadP2XSpCx/bxpmQ4KqP7TJ3l1j2eGyLJmrs5y309C/Ea9bXI8dkpmRCZoeTMyf2
J0vs2B4kY/20BceIq0lkHjBvUX3Hvc/JbeBgiDvlkjfetR+H7SQlKR40CPjkbMcY
+kokJjf8fDLGGPNWqszLd312iaA1+W67R6h8ZynY/zUg9au/Y8UZEfGAFMM2YTCo
NdGcgj9RlAdmqNTDX9izw7U47gfgK/qTkHbXiRzMzJ8RcazLc3UTFxLln2/TyvA+
2hya5klNrM24PBRSY99qWysIcKJ232vn9MJIruC9RTbG4J6zrw/vQQ9m9KVgMiuM
i17BOeJXAbtlGHi0fIqjcOodi+g8NFCSoRTy4+JBfBCof2lbyXUwmLm0ljy1GBp1
pWSRrlo3Phrbl6nWb4wnjZL1jXJ9KpgEyTS+9QzNJMhYeN7jC7H9FsDJlFVFKjIY
+jDqwHb5egUgTr/mjcWf2Nfqr6rSOETRx/C5k/KmVRp4cTair8RYVpcmw/4uoiTE
PO2khbGflhjC8MwmuC7zTb1fXeTwb/z6mqVvys5gpDm91bGpt/ujP8AorjiA2ufl
Fc2zb8YSJa9jXBb1jnIntKzq7NpHMO4OyITHncuiMPnjJbyPuk7eY7mv2pCOzXJN
ylScsExysQSZXl5ShllbcTqzwhnXJbrzrA0ArzX50OeFP5RSiYYBLcA6NQzE0z2W
2nIa+fSLKY0NcGYx5ggZHPO+48genSiEwQFVhRRGNf2y5+71vqiPHspjc26Lb/Iv
AGlSbgW43urHKj5pm7QW4BrodL7mm2R+PjeU0hlwqvW19bRlcAc4Qn6ySpdiPous
2tP8peFdBHyxSLvvTbbo6JulAkeHkP/fiSd8kpgTruHTLTr8xnsXbPM03x2XkdE1
mJ4abN5wKUoCHkzX9HWad0mai83Lbr9P9UhmVrItmwBApit0gNjK21ANVHwAIwCQ
j3sMkeCkpTVaChu+nXhPJ57GfRAKx3i0WEBPuYwOG2YmYxh2EV1dPr0Mc5wrQAj0
WmkFf9IN7TbVZ1X+TwYKmJyYYjx5aYF0/nV5o2MxstYn8zfUOXZIgxNmc5q9pADb
3JzN0EX9MPXkLADD2fPq1B+OLXcIgnRFDarrsd8Kx6A8dyLVJ+qtRLThc8g7apco
6wfPGhjCyzLYeKEQmmgupY6gCxy8/GQ5LxyVW9tqjUZJiOTkEIWtbhkubloKnY8O
8UH26WYO9AKczXyeDO979NIL8usqzN98hrK/rvFnygtDGvxpovq7wa23wceOAj5l
Lxa9TbS/Uu9K6yFKjrCsyMbckhYLs9J2ITswRDwN14Aiak69LhmP9E9VxOW2EpCw
vFXfS8zC05xuFzO5pTXGxU5AdWTZU0jRcaYyLiUkCif6LWUauq1jOCt4WEg7dBw2
xtVQmp66HDWXawH/z0kcDVw2OVUpWFz+lC6tupFOD0Q7yRKYRhA+YQYRULSuMdOY
85KvMoQaneWnBGQ7RFLWfrXwr1G41nauHrKtqyMYCMG53c13WDq/wZLcBQylRgF1
Wp5VM8SRVHGpvMYYugJEAy+J7FXgVrnqpEE6C0CP+KwXuy8w+Qf9ZkXzmG39/2Gf
KGmzJRvYrIVT3XnmfoEvSb3YN5tB9G42XBeujdPXsg3WinIyEi+GMZu6ejl2Hvtf
c7XRVgTXVF0NuE3OixcfD4U7QYIPWXmbrF1L7ZlfeRuSx0BcjnLE9dx8umOrsSNC
RBWPVstOVqEp3iLr8EJooUnD1EeHgwsSNh7vITttow+o2Atr9N+IOhrX7YRfSAK9
sSw2rQvBeE9Hj5OJ9YNEKsCD7dseAyV0/yXqDH3ZtH0mFw59Nnh0T2+IybGeh6do
yUgDzRq4x0UrC7o2QF85Z0OlU4sujDhpkYLvyrPuPXA4A5GH2AzkmpfATbKwH8FA
bWOJEQPPRKYi+fUiRzhUgGG680XmBCzv/wAtrksFGR1ZBprDA9y+skDN8d37kaGm
P/yzJDIhGDC9jOelOfSaemP2yqbBUR0A2YCoycF9OQZ0Jay9YM/TPAhaqiMGZXOa
RA2/p1YodC/BaxOs32oWiO2YZo+75ahm7AGDAPxB2w+8REAB32FF3/GRAclf6LeS
gp8jsOEpPzML19NRlFUoJUQv4OC+5H+hpW4ffbv0RxYsJzNKhA3CjPuAN/3zTajb
UbdFeVieEugO4JIUwlq9Mmvyckp5N09doIP5uQm5sx2WU+uo/WKgYQ5CBRpBBGWg
x3Z/CYv4Lkrx6kKuswlblcMFXLhihwSN9DnZITDgOp2prfD5m8/uZDq4Dh4H2ptJ
pdI9RuEDkYXE5jzRYG/urNTTUfFYsxtIqZvf8+spYZ3s3pqJYzYsuwxR9klvIkEO
G4QdMnVYeKkJ3aa+hbWG+2pDI/rGznc7qJPDR2ZQpT13Q12gI0jmja8vwGJEJGbz
WswUzvxXBShhCrXjMC8UA+Gsqz4Hr8cjJERQwUYQ3PtOjv066gDyEHfrv7aIH+hQ
kP6/+f1PxP8OZ4w2NfEMMJMMU0ixJfuZGmvGRCNgotOIdmJOg1VEqmzbX6fJwJtB
LqJp2pcVUqSfyOxOAlw9jshmHs/KmCGKDMkhTAr2yN+qDCMSWroXOWtuP4IbZ1bj
qWL05ML/NyFsLEpJfLpCqQZ1xNaiUXsyDwfW81nYuK5EcWxQ31Xy5YnUYhjwlXE9
AVY62bqbAcb7Ko6CEYqUEJaG5gQ2ccLJuTBiKGpQeIrNQQZthM42B1KULNNS9lM0
LY0UKGN+mLSZfu3gpxpGQ4ly2OVABta7bMzppsZeB+/w6/lIt70cNSdlc/6ttDGK
ko7eOjR6DAsJsIrL8Jn4mMew/XBB4NGf+4hN5dgmomQKt2ozeVJIG8M6NvgDPv1I
E+L9SUWeoyDNsnADGvgT8RjGulsT0INtIbjZvc7gUi8PrfvJRX5uAA54sbOxo4xA
6hIQ2dZGeqx5BP96E4hkb53x6PWgHPkmb8kNh46z+tAGGIvpBh275CJxV3tlYZMQ
V4M/wXJ/FYnUF6/LqjmOh3l/tJu58anHBtduP69FGDyVm29v+yKq37rRvNHmVL2z
nQgbUjYYEY5cVV2EGDQ0gfdK2s2E3D+rPTEsW8mF6o7K6tIkkJG55NylEmkWRC3c
GWPMOWNq0rwfQD+SGNUjyN0ZXJsOmks/8YiHQs1Spz6NYBYlATU4Lposa7+wEaU6
nqkMkqaaQsP9PGjfSg/PNEMVsV6Mi5GYaGxPwQUIBifxtVMF+gVa3DgfAucLd6qb
sUxYZVFZr+ivoWEpcXVMe3b16aJ87PQCpIo762CgQx/tEpkElBRJXjF21oYqjcSC
bNWRT/L/Ko01Dq2ZRl4dAS0Px3b+HnQK7ynWc5AY5g/YbKV0CEfne1I/F4dr2Esq
sTSymGztesUmxDhfeiSak7e10HYrujI4Z03wk421q1gF5cWzjRGkEhsLKJbguEmr
m+kqQQNdn+WQtnUb7ki6t/u1kl6uMYnXnSEgEvJEFvZuyH01qvlLsE2JLHwpqX/0
0hWytIyqO2kahr+9QAdXiQht4e13RxVtfJgyZEyXW0EdfSPj3/NFAzTHCJeKj2gB
2rRyw8ZkwFlmYCOhcNfyLbTlEoYFMr4NW1D7EzlHgej5xUIHvhobF9rbIrCToj1D
FNGjVQa78DUFkZvKrXogFJqSHzNzH8Q0WcQ+yRj1hBPixhxCvNMxK03FolXznyk2
MvUsizgj5B9YqW4Lpf98nc6OET4Y/Ez081V9QX2pPzuS9iUJFudGE5J7yzWPt0FT
gYC9oap4I/ac8nU74j3PbAZlC13p2EUjNIG4zvqiqLQlcln7p0jGY2BHr5OYoDN9
pua867qDmqsc+nBk5fCRCKgNsQErEeMh3StUFKKxoAUV7SZ5T9Nk2T5PqnAnwU+B
QUpZj70H+eXhbbqcjGz5xBYh9anMUPRzmUDNi+TzefqSqeAgf61VhtagmuUUqufi
MxrqWAKrbL95u4O925M7AO6ijhw02PmHVLtLWMZbd000Ao92SlyuAu4mmzld9Qm7
MmaoB4849FvhVwxCqlRWDLgmB8KCdBBIuNhoziPehiHiFvO/IHmi4U0tw0rfl1pp
s8lqmLmjSQ1XKhNNvl2s2QLzIdbhh4jJGmSmqJOPqT8p9MqdnDdF0HeJZW02YZhZ
dU49R1Gcelbt1yes1ss1ncGIDmKwFA3hMpIlDeTceAUIHvpGxg55DyIkWSVEINo0
A1s+pau8lpxgiMnnYZJb1XmHd/Wqemlyot9cIQY3p0ez+yXAzW6Q63yBelfkFBkK
u2wCvw89McWFdVyZLlPSOA6S4iNdhKNLJkGlwjpJ/lu0pJcNEL5RUEn32icUPaWV
EPHI1dBt0Nbc6AF8/MTE6aszMa0RpmF9x1LD6GukjZsDlJwu+Gi52T3io4RtWKBn
JK1J/myWxh5voY+rMIB0hpQzQ24TT5fuOILn2UAV2zLePrFrQ4JPcyhM54k2RmMI
IOcq/+ynKi4Qv4NA1mbGlKZwKSmH8Fiup9s0xbeEU843Opm/6IvDtsXLg9aUDAHR
k5BUYBtXhUN97w0U7LrkgsVIwNmQryJH6TQJDKtq3GbtGtMrivVchLm5RAtunwJF
fK+FgaIgVyAi/IrWgLWimRgdMny8uMOMJdPQtOpz8OLnffHb1j3/DqPI/Bq0y+R0
rMiKBYmCgaSlJ91eGHwCN9nLLKr9qDDqO1K1UxZwmyMWeF6wIAQaPdR7NA00KgNV
eHGgZ26YgtRulLg6LEmna/Yfb3BAV4aSea1Kxi5c2rP7SlOROjlcG9RFsGnv530P
sszEOZ4apazpcSPcWx3VSQdpmsr+up1vUhi2D+SGLxRUd4GgmxSsJHVtd2PvbVDU
4KRdjGDX513/vo+KsYdUWRcTBD5h/WoHuiIHnet1Jb5bnmzcWsfc7E6QNRzWuEOA
E1N1lF6PyTNfrcMxGgYspkOXNq5g6gojRODY0QTWeI+5lPjjVC1m0m/idlsaJ3oo
8gYG+Zmu5gLIgy/PrYpVXKU4VkzNCgTwhrXYAaa8T1T+b3JmxMvOrZU3OZFfg6WC
DLtd/GuyC0EQRSv9o0TqXhAz8Juy6tVP79dA2CHlixJAxTR4qHoEfs5RyxxB1ISb
LXYlGt1pdCCuJJEVb3UvzCVPx6NDFHN0rPtPAEry/Xi3jfwe5GmsZjmuIBtyq6AT
zHswuZKpLdPa9f9Fwu3AtSZx4PEXP0v/8pWPcmO2q0HI7zI/W/h4rmgHHs4ZlZRh
+GTZjficEckxQTFhH/0tb9ZdguckcW1EJJKiWN11Y2s6NBNvnVkhJb3pmOaiGWsf
Beqh97EoLAb/mZlnSiFh7yPa0Yy1nCCcZxzdRW9OeSrKRhljQ7e0YffQWrhqwYLN
zRrajUldj8kwC0wFpqjtslo0CpxNGwTVzQ7SVgMWPfiVlsfGgoZkZv+LtV3BnoPh
z1uW8Zjt42iCMxgCnmziJz+fxZlc3vunkm92AnSOzj1fXArv/2ip9kk0UrMGFTrU
o0fOFogpRIQOKoD/67IgEv3q6Ywh73o7Xn9WVzXqdHCNKG26fhP7c3cpOvXuclru
Kjcfn7odV8b+ADXwnolrtnzcvIiy0SH91qMsTWZZ0PsPyKY22+idpbr/3j+JwJNR
l0xzJUUxsBiCDQzs4xMfa9nZ+QDzl/QJXV9ulg54k11I2KIKQAx3snfss2A01um1
yKNpVF4oBfCJRgwy0f0VAJ9MN5Rr/M8wdD9J3Mgr/g0dB3YyhyMNbQY8m2Vsbyg2
/Kww4yaefKrA0b8jISw3mx7yfhGnMYCe21KNKV6vPZijsk0BwsDdAu1K/lWKPURn
3ZQ2JKo9a0/TB+qIQJFgro9yhNWkQVU9qmcJNFki2mcKA0M94i8ckYY6r72RBaJS
rQ2DV1h1L30IuhqfkNgihT/cTuBqg8mw/e3EhpYhHL9cAKtWlqzyh0/fhK6FdyqI
MVTjZ+FWrLrN3S5IaUnz5kIMp++nToP7qPt5fOCLdzj9qGRxHvoYU0ZC1nDF0HS7
lwah70aui0WOEPrMDjNbKklQaiSn0p0VlSJeqNxdHa+EpTqhCj6RKUgwWv2NHa4U
yFY7aJhd/w8lznszhICanTz208AfsQP9dSN7D9FwgfwwA7mIgXbG347AvKS5U8KU
ZProAaWEiW2VqDb1RFx8CE14aQICDQV6897/rtBhv+JVlYHPrJqwmRmgH/5Mvnui
mlhdx4MzFswLX1XNa+KUWIVMALuLHhmmNLrElxHSu/gsstRc22MdqiyjgqV5VP60
Q4AQJOL8RqyhFYnN8zOKrZQ6wFrWhGd8PTJUXDtoTjxXsaBOA2T6FwAC7I5pbKOW
iLxI+9rCNuc8jRG7btHUDy12cZSgZcaFr9QIAt+4vpdlxIlDmlmPOByR5ROfRk+e
yOccwt7AUj1rl6UqaNv3hS5R8NJdvTHTknXxxlbLDucdbZocbVASCmk4DzuVKA2k
7EN9tshV/3R+U5mub4A8Ggk7Ecj0rYNogN+ya4PObf+nciLvY2DgMbSRXCsUFyHW
qEA5hefqvPu75Za1JDzmv9RThYxWOESPoF6MiCS+ulMwLE9LWCSGTREZ61KiakQ6
8odIrbi4bHU0TTFxB1IBOncTWboGKB8eVa3qHkzCw0fbwW+wLFuOZ+YH9tjonPXl
vacsj32bIc44L9j0egJxXugNsx0FnJf1/ndgGUyiGBN/tgnk2ql8oLAxfLgpYXLI
aHeotFpYtgdKtWjS4WM8RZSkftP5iHlHNGi9hoqC7FCmgHUXyJYTp17SfLSc8V+6
X+PGRnrG5eZVE6bt/83VrR9aUQPcu6UyjdMgWr1CCBGSzIR82jiTGUHBUk/Nm+w0
pptc5H99NvNKHPCVMB+X9hHZoE24B8T3aIy9bdFw5zNAb8eJJl+1/lV83a0WBqFD
L8wwtID0ndshVcs5yCWaRRIbV72bosozXlkJdHQUGLFnaTwPqpQOGVenOe70djd1
3cf2raRbhTTmw6xHzaUuQ1w+6Gjl9ugLT6Yv8NwXTRdlzY9/+304lXcT9G035Jqs
yWArkCLfyh+6jIDl3kqViPT4038DKflqcOLvHENpf4d2Pyz53aMWUsjbMZR6Po6l
F+KFwXpLk2gleP62aYuUdAhXEkc2j2+r79IW/TExxCnxGCLSNWwfHncuXmcBSBPA
O79DUMLDSOFRBivqYqPgHrW/MXtNhYhQ/pJS101YV4GQEMv8mDsb9ToOa5ZLqEzz
iTBeiqnHvGHcOzm6RgnCQGn4Jr8nzGyzmk9tLjW16dYj3uhtIzc9HaCXN5pv9c3d
1CA0ViSVVKPuHiXPJJqgPiy5Q1UZ5OSSE62xm5AWsZdmBXCown7gvY0LUVC09p6i
fKfJWjAFLGtdPpCNFL8/wuPqAvrzT/S7XGr60WxGRfiUVyLhNwzbTX6Slc55BMsC
txca9j5LnNzg60NDp3XahHyrAxYhRi1LlTRW4vaQf8+O63sZuDWQ01z6J7iPHy9D
ZHJBgvpOl/Lepogs16LKSYPQz+gMBGGTPgepURnlFe0jUcFWSpmEnOidn6mfz4hD
XbL4zWF6xn/NoLvUlJEFr5xPMBQlaqBh5+VR5tAA7WKSJ0qGKNLukhCF0KnRcC55
NKiHyI3Kyw59d1rZDZa5EP/m9HR7plIIW+ZlmUcTUG5yFqwj9/gqnYWRgErA61tP
ol720N3T0XrU3yMRwT5ionGdK0BgP5j9k7LWOaNEBoDzrwJovG2+G50r0XaoX4x5
iU9M052n6lCILKnyaZcAWuQ3Fdod5RrQ8f8K14JLrfu+vyKOzOaJ0IVHOqsfYZF3
tTHIMUidaA1gLloRyUx7o1msWi/6akcfDYWMRw7TcvplEPm9Nv9nQ22WQ4rI+pl3
L+Sb+88gJGdNiZHhlHsOMIE+sWeyrqMqGgpFXVJwOyXw6fWPpGsO8oTONMu4E/Nh
z6jcjCoxnXneZMj73MJuKAtz4aDjYAmOBKmV4zodoAx6kqXmBDh9Joq7Rp89Muvt
SdS1B5OLDFXEtSswCxdpaAnYuYxMokDrWIMUxmUCcpK+K91P7cZOqbT/+T+LY8LX
MT8wiaSNXXQy+02g3f3cZJM7z28anLmG4bFcePAajFGVvhN/2aYKkOy1pfdl98RO
WJL+jWvXNSGt8/6ZCRKhF494p897SrbjmWjrt8w1F4LgbU32tnUNOCdGxa+shR7Q
27HDnTOh/IGwi4zJZBObIH8J46DWb7GpPe2SQOK5H6HEwjYl57dy03FiWWLHx7Ey
eMLT+euyUALiYNPWec/IPcnUUtDs9NXWJ1875Hf0wcKXe12R1Z0zxT7jLpWTEjB4
2yEDQ01E9EozXchDonrgGrmtijHUOikr9x5QAfG/OjMtdkRwV7CwfU2lnXG1MyWj
WGOrx2rrxb1XmJXalXUh6WMTnFZHm/t3PlPBYd4Yfttci8ev1MoEASsw5Rgr4nTp
9YECgEO3THbjnH5n3/lsvqzRoS6ZA7VZ9/e7VYgQ8j6EYI/6i50gWBs/DmK5K3X+
aphsDbBM+ERZFnsHslnSkkrOEXzYw7hcAnnsTGOBjrgzYj9R31+q2jw/pFxlYCxD
O/s0ehGNLrJSYUAR5otIp461CwSq7uY52BTG2BXVBt8EGFY2giXM2Ora+0lvr5gj
wteKpgGicpnE4hIZXqPbQMbioyCvxWw3b7OtV2jvnnCo7FRO8VYo+UCtfWTrxiwP
EjsKYXF4uFGqphlHkrzuuA+G/eBxmj5t63M2nbWKYUGleR7vani7G/Pj5lr2zmIm
hfkWLXZChaoIGckcAUxwi81jDpUSQLbtSPRcHPc/lgt27xzGGt7M4x8eYRtWCQOL
g0WcjVvY+FVapUCjtgh/Eqe0yX/ahFBZM9z70Wtnc505X4mr1/O3ykz8LDKaFr9g
+9nVQZD03mmnLhqy4Iggd73uvbPZxJP9VCYtK+bDgJ91oiPm3NSqbcSN1M4FsdkU
tFDEoxGkNcbajifOBnqnYq+W9k5W3EjiXqBrMPamDlzyW/xnTvIzVIANx0pBnmk5
9hB5cC6/2+lYztJJD78lUsJGvDc5kgWYhOfvXV3d81sBjdak2HnJarVxl/lytX2u
MsVY6exgI1YfxM88DGLSJQIqomZAsSsEKSKLyCf1noY1YlDrBE63xfym+VnrEHfQ
VC3/6SIiWKnos1lz1M/10RpjFGpsaWlJuf58eIE5OyJpkQZ/n3nhRJZPtcWXrWhx
qGdmFeav/csHFWTo5+ELaBWw1PYEfstekslQJI0vl+zotPhZ4ehYjPj2VeUDDQf0
HDqEdHdeFLg9TGhjaB5iXLDO27IUPUufbL1th1/4/dhK5dArVBJvuDHkTkM2JDPH
s0ZYy4El5mlSKC4ecn89i9m9X6eX+TOqnck934q6+bsUffvuutvhyPfnHx/p9pv+
JbcExsokotYmQq3WTZenOeTmbqNJha//ooZPxvu0NgsuAlmLRbVjFF1mnjZ+dlZI
PEV6nmxCD0WbHYespQf2x1il9KMuW+HWO0s095SO4e4iWXYi8crX/1imyCfoMw8Q
jYngRzBsOZjGL1lju0lVsV0E2o6uvf0KVMS5w7riWb+kAwlOkcwW1/gDdN4W+xDj
2yCFMkirsnbWUk45bs92UM5jGCmVV2Hfmk+UMMFE9nZnp7EK3rzTpju7yBQ304YM
8RcmB2FVVspeiDzQY9K7AsUBD509D7PT6FS85dvRQZJBWtzgHDB/fBQmTFVpXYTD
GASKTFC2U/GoqxBXMVF1t4OQ3bTPvhSHjWf1qBgBOboKlW+8vT2civ7ajTOZ39Wa
Do8Mx2XeeUDf6ycqtXCI8t2+9MQLfcmIr1CqWUWAWj3gztAPlq+c1RxCOzfpU0I0
l8vqliZTdbNTA3ke70hmFAyKG9NqN4gDcr3jLE5nolITNLWdn1zihmmUQOUkDxR0
p7Rt/sZUjNcuv+q0qA3s26FNhbzXxO+UdxKNXidv1g+f5M/BN7H9VGJSrID4+xsJ
ZK8hsl62w9/nZ+Oiuq2dw3pdptHst5zNlxCaKTwHEG79ajZ2F5y5vcoe5xBOnc3W
XEa4EaRpoTCGksC9ivqJKuZLiFZtH34/OZaHUKxT5S27Wyp0qOhlwDUFeibamxn8
vnB/ljC3B5Ucb0G0eQwe10M0Ms+2ufJuvQivD15/sdqfjFn2kIqhgDyNvGWbnPjX
QE9ZL4/ANKNKtFm9gdsSZjN7mygELJcHANSXNOHUx3Xp7ZTbHRRtImP4gLD8Pmym
rr2xnFpbiuOeJjm/tjOO8cwmND06OFIoOWwV7x9kiy7UKnTB95F2/Re4C+okwhzM
Fe3IAvamNyrUC9D5aEKnQqqo6xVABo9XVrXuisKO6IuHj0FR1YSv/Y0vReo7GoDR
Rj1izlBU/6zLGvmRnD1TOtgVYC5SnNFS2CKjXRFg5NTDAufxu423D3X9Z2qgYpce
J7udpG0NIWXKRUh3jkHO4Ts5XvbO0Hfbziy1MyB8Yu7TM0u8eArn8AEeqxAbL6i8
JV9jyWkpX+G1XRMulhTwiXZLXbu4XwgJrXZzmd7e+1mYC57ZHTVTLUaQN/k17EfO
7pcGFvlGFXiP+SKMwWsK8r7gOf+sVYaSYkYk+naa6mAi1jmffJejWSwlU0X1jp/m
nPQPf/4auDelLJ9YbvCM0Yorbp1CuMZMSwbhqSTIMjnINx/hTZJ6DTbfPBiEu3R5
moPcvvWN69jEMaDGYpb45IwF78d0XvpCq7WiTxwesgT06FgRJgw5DIUoAun4Io8y
MBH5SFXu/aD5kTK1wXRqwnKyivJDN7xZSy7qtVqByWrk/f8hZf3j/WCzItvpkeQd
HoZh3spu7aQG8j+JfALDA79gpzyGk+EBZ0S9yE688wifELEBJm9pdhi+rPqKczSC
xNP5SKLtK4Y4S1nz9oVR1QoWGgSQEF/rms+zJEqqEVySQ9W+fbQdGhq9vb+nRmc3
jbWEgAypHRzGkm8TSyPT4YeCs0V6mxxbSeLbj2+nRT1AbTA1WXq01LlW8IrwaKHq
TWf/iVd6vo90KqSvALs+8csP4QaxwY7tUK4qjLGE4y0r6nDoX0UG9SCC1GgMLaR2
eWabs0V/jFzpSbLRL6PxU/PmIGNf3LAhnB9jck5oCBVQTX1kL/SDIfGxhesqDoSc
ZWFXwXO2w1241rjdmG2NfFk/5L1UWTll+2TwIZCL4R4QEiBq37D9K+/9BzTFwj2/
dOTpi8fPvVF76DeKr7qbcC/EiIrHyF/2GUuTKIlf2sw3XYSmVuydYhMbGjYr9ilv
cc54hRya1N8L+nHdkCFG/smd7R7/yhSuh0FB4dOEQ9g+SoRSiwBdFe8SQa2xRCal
aZToALpt8yjAef9ZaxYlXtUxyiznYvnOAhSkBXXj++95LBThaq2rGEvXT6H/q1nX
4CNIMslSfCj1fUiuVBUwz1csUhbEO/HQ39XB0oN6LHl7+5o8xGMN4lCXb92GdMty
MgqcEbwsI2EsoS3kf+mXDAQUHLN5rINeD2jm4N+bjAOQIJydNxtnjD+sTprQIoxQ
0+LioLvxyrWU9ZI09W9ebFNy2Gid5RYngkl9865mjqUA0XX581ISyhTGsWPxXt28
Ux7+N5Y/H0vRdpOjFroc2SP1ImCL/k9IjrfhSq+1+6SlDIJ6+SyGcI/PFTiQYatY
Ts5M3Mq5SVCilrXy2lxHjRa1T1AOsvQo/VoWsRf8kHr4e8JbS7XfrpEzZxw8T+Nd
JyML2gyUr6iylo8szDY4PJpmIdRF7AFR+rvt1Y3uu9KtbRTx6wGBL+fjxo37FIyU
XZvhxXkD1t29qBlvuvjyVlCgXQb/GD8baIy+sNAiAauzYi/zTHzCNZGWRPGBndUe
r5wkhAMkOVxKBO2PnaXw/z6JHc9IJb9tvqoo6MIjfTt51EzHLiy/V/SG61LuCSup
HwGrYsgKrynCCl0tsaqs81bhHeuPuFAUWNVfcxIxavEKIh4tcJCjlFKykJVaa6gn
ksiz2xJ0slEyjYBkYrmxYrgSjaEUQaBusMD5uzKXdX36cOvJ1cLYg2rbiTob+WkG
oAXMTQtQ0ykpTY3UE/INPrHo6Q756IScEm4AGpu2WA5SIawdQrh9DOGI3a/P6CE5
uAeKKL9nyFAYt9GBUdSUHGlpDdz/BEptcKe5ZG3XuvYU3JtODoHVQwF0QSTyk3Ou
KMSUzGOX0WRxmfwRDoit+A3sIrrIsmQE0xGptvm0pO6I8cX4mRmWWLkv7vkOglKQ
7PVRkmHsGOZMWq8fzhiUbcscjYI05PdNfD8Lbri+ebY3u6vHmcYIBAAk4zBVRk0f
BmgXSngXfLqK/krSExmcn4V/HF4jfnAVj5BeI17RhMNZxXp0kqkSVl/S73BoVTgy
bBSPoBwmUpHAfvWLXEUCCJ6GTa1rtBOUS9KIZJMD63UE1Y0sJR1k/RPmztuifR/k
QKWiPV0XD5QDxmw6oXgn7h9MmCPLnWL30KFuEoEyRjtYD6CmfRPeCQtCxfC48qym
x/HfDeF31ZApt9m9unDx8P48QQg60Qw42xWabuiXAj4OAOFB6SHi4AMhth5WcAtF
pDwaIXhVW6NdSK9EGDfVjvcWXWE66vLLQZEu8ka8l9sBK5Duu7RxIRfFuWKJUnfg
XZcxu9jB37P+YbVgvRlfVraiPxSM8Ck+A+OqX6xT6xHpjcxq+xdbZtEELGu0JTEs
sRJs4k28TpWJv0CdJNjNplEQ9NERn1FLLZxevBsFXHYi5eMumZDfvlAWFAwPp1Ru
/nYhSU9Bqy67NDbzIwbQg4vWwpvJjxYh1JA4s+XTb/I+GnnRN1iGmqk2iahnK8ue
W8xifGPUsex1NKWedJT5e3azhsgKE7vPYmfyV6boaeUpsu4mDIRXQfmNLGhuJCj1
Yjf2y7dlqDdfLnGTKMpUQlbG6BlysD8pEMSt2eRwE6MgNRpa+Slo4Q28/nQIKHQh
JZ0Uy9J1vj9XZQTHfDio7IkRUe2Bxi2mbNmu0vr8o6SFHAgeBmMxhG1OIRpAf0/G
EfY6LN/oQkROX43W3A8i6BURPQOIS2q2s6I5YaS5uCQmuzi1rfYaJLfoBrrVC4cb
nmXXuhGT5uSkc0gJZhdITATJwbyKaftXuxC+lO4WtdBX6wIURnS77jt+K+KOwt7j
5tkEHZMj1KdyykQgqYRiyaqqZOEW2w4/oRy76IuNoCPWDLx1rdNuCsfNOV2KHXcD
d5gAba7UV12KVj7plK+ioFuquLy1pp/a+unMah37qohYMCva4tpMr3FiS2lnVBNX
tsqGzmrBJfjxD0jN7QNU8/ZSKxN47H4h6VFoGeDidetVXOsTODEcZSlvVis7TET3
WWFPAlL4cYThSP7jzURZcyEYIL/pFdRoAhTyMh4pwmhxkVyOEZw1FnxUYjtxmvmk
RfXJHwuX7jrhYo/YIUwXkp+/PjAPRMe378/NndF5RKBZSg1NM0bUxKUwji0FnGaF
/z4E3I7BnswymJuc4zjtGh4kUmE4gqIrg/Bi+VA0udtP1EdYstpD4dCcNIHcAVZQ
MYMf5qKNkz7ugdaYR3SpJESSw/OSmiZa0OwNzTF2aLFNy/wFCt69ecdiJDIC64nJ
046ph/o4WY9VsNcRgvIYP7AOcc73gVGpozxpWBmuQZkp5sKv4QLpc/IVTSlACWYP
qTUX/JMBiK+q3vqCedvDW6iYRv3bVbr3gh+8oYbqfmpA2R4QMUbknv0Lb4YIJrhD
lLfmJSVaypF5Uro0IETrrAop9RgXxIbq16Pg1HZtfFeL5Y3p3vB3k71MvoA+BjRj
f7wgk2xGB6qi2GEOiSFVS1WvYJ4pceyz6avBH8VzoPM7QoHtZt/51aP2nX62s6KP
zqL8lSjSV64T4DBtYPZEWdC77Dck8Ybmbk/giIvrxq4R2tic2lonSq0TJiiJy0r3
cPni+nrSY5XTir1oO1XNToCgZ2SnYL/L0HV/vYHIcGDHPzRLXE+w78b48QIzOB0q
V8NCrsyXTg64z2q5DSS4vSyvh0YPtC1u7MYgQjnOlhbqLxzAuo2ij+MjiEuRUe81
eaR2i5qBjbw2GlJ+SBY5zcutX56gOI2HZTraD2phtv710EO8ndnMROOWXGRbXDkc
MqE8Vv3m26Z+sW290K1/2C5X/jr2TqkmQFrHofCXXReyb7WFLkAViRX6uDJcxlny
WCrtv/bJDvrlVTBCYQZhLqFtT7VCXuqcM9ALIQoUIOl/qR+whz4dPaC0LNkyEl20
K160Q7NXx2mE8WtjooUVWk/whnvSkYuS60gq/eU4GDGJeCdHdHF/BNB0L7uzTrdE
tt4TW5CkjO0lCZWUQaD9fvtrc6Kgf1lak8Dzd2Iesp03g1/y0ggJQFvsAYpSN5bk
GdqujOZfuyVlMpmzcXcTSNRLNz7wurTvX3bXkdJtpYKPTxpmLk9Ak84AY+1HtRmO
2aVhmUqfoLSoE1JcUHkViZP9PMbe3DeUMoJ5N7wTK29E6Uju8MPdwhxS0r3u/ifv
9b4mQmyqaLTxA8Jdctyc11I7wPl4ji5feTjuRvxWUwH254JDccoAJJGHAjRIQsd9
Wztw7Rhj0hHRDFcxboPcIIGc9DUxi3MtzT2jSmewORF2101zBeIhawYal5FlY83r
JHq8txIQUm2hl23YlItL7BGLEcCcZPKPnjJyQZ+EY+9pa2afvKlykjIHbnJfk7wr
bjO00o5whDKT/RmMKxvpAcsbHsPV6hOefYNvZbE2Jk6GOePYeqPj6XhYA394sZ7U
GdEupwZNQS3wM9Of+Yqfs7XiQ60G+F8KtlaiEk3TEiAEyAGFfkHGItYiS0sPbTnl
WFe+jRaOKcxcvQ0Y0bNzaVXSQSnwTswcqhmTOCKC7H1B4ip4fQgOjNipPRQiPsSq
lootoQo4/AXy6DhUGeoi+aY3VzqMRfRqoAYSgCjZRhnQwgd+eXpY1zPWd0m968Tc
QPIEpvD75Ylg1mfHXGypRy+zvfGCPiT2dBTOpoHe2sqdR8L3R+70cw/WbPJSeC+k
p8Ydj7LbNGL+Jd4pO5059XwLskHzMfX7U84v1Z9FYue5ZWkVlsEs94umkm0xDYm7
Nermo4n4W+b48WDXQC/4w5L6oJZHv4e6n2EnOY/K5/PN0tCdRx8GYr8WphaT3qNp
lw3iX+nQmiPTOVYMpbrunGDqrwD5gi7F1Hz/xYEN6Vhdd7yTpD/JmMFv5vgs3var
b9y7qjAilOC+GcCnfXs8F9JTF1Us/A2roBMzmRkCc0KY1s5IeUioBiJPg8JN0Fla
SI3X5ud6VfNJtIEV4ZJT3jQW+PoPL8O8oXXZOp1fGhWq//PVSuIG3jC4UKp2emZC
F+4uZBgbaXi9giSA/M5KYOZ/6tXS6qr12JHEgAoW5w9VW6BnklIEe3gWJRJkNN1y
KLHL3mM5T73GQOOpxEApwoL+9YbVuBOuHwDphPIKzxFIDHyycml09GcXtiaQGuEw
VObckdz108kg1Crmdc0/+SGQ901RFFby/W90wKgBVhRLivxie8Cc+wo6u1KC99Uc
/eRmgVcn2+9KeE7SBpsk8UtTKx3yOq7uLdgKF7Sstxk6NsqPuD1tqQL9EWR6ERBQ
3OayyIYrC1TMQ/flfrHILAiwKJAZpUL599ymCDWI6vlhImuyCgQVNrlKXVgtG+1u
9O/7fNMawYXpw79jc1UVCOIB6A/lTL0R2L0n9Pk1JJNa+pjSqrdGIlYZNaiePjgy
sc4BkNHxQoYHWhrM8di9aUKdnCZ2YewnRZepbTxU7LcJ757sG2sH/B9mfq7SIJX7
+znJ3OT/8KGxx2gi7o+wthYvbVosHfWUj2N1abLIbbItoqOoikyTAicCjkPsL2YK
fhF7v2khk+pqWZ4AixtOTI+1/dRYK2IodK29nuztAflzddlPe87ojJOX1Gq9OeiL
ISqWd2YWHfb7LkmfiNRUtXMet4iGoPuYIsFRVMV9UZhKseLdqLpVKWahwFISJxuG
yX/W2V6p0NH1+qmedmZtl9xhsGCSMeWd2QILUbq3qn+YIfbhZCDRPlnUA+wOEccj
F7cdaB3m8tFBrXT29iCeING6Ya0n9TGnICsVNjhwwSy/gsrWiiHn4yias3BANpe7
s8rVjsMjO3IMIejtsEwKfheY3nCcUBTIXhoU3vQkhAt+hnSTQEndVsOjjLsPt6p0
dvflELUrD0VmdQnPbtkDec711znYfsNtelx3CCTxogk5k/tJwzotuukir+P8Frf1
KQiJkHsCxHyGiK0NxGxMnmUeyDFJYT9fBex505lEZsjnsgN/h3VmGb9A0+5QeBCq
229ZXpys2cu2mqludw3U69Qox8jPbBxmlLLbdg5UdfQ782fpjLnmnT5CY7q4H3k+
aaXYuVlPTOS0R8U1QBAVzfBmAdKx3V7koXKBbuwzTlH6ix8hDDN9z10l3/O08vZ1
jD6fCEY8p0RDbObRq76TcicJKZyxS6TBrBeq05rrJGfRmbfSLPARvnHtIliHNn5y
EFq/PCDyq4GA2arXzsJJR7jenctyNPBef75lYC4Gaui8OxphlxbE7azinALDe/Gf
KGWhuaYzcfQGVOl0XV5YHnfJ+OM4h29aB1jXWJTdKXQoRAmbAge1NPSPGUfqG3De
MaABCFn14RNB5RizhCu1Jor6XBKbxM7R8Pider3PHVQajLK6SEzAxuK3n7BvNdl8
HjwOO0pQf5hlQ488VdHojdbXZFP1tBxnEEVGoxtwZOF8yof8zHRfSgGWxOLQzq2Z
DuiR0eFYOM0geMsPrh5MIJ1JjpFeBOdoKbprvp70ptURfmZhnM+sBpjjEvIhis8W
40BslKiDfO2OEhYpk62aZ2yJWd3YHQ7IGY51y+ljIe7ML0dCg5lVvS6TPuRjIE4C
XPOq3Bs+8J33KtfsftqpyyduKZFjGN348R7jNgWb+G3KbvZvbbfEQTELvnF3+7Zz
JZLHrn9nSc40F0QwwrnXVvINaMAunstcI6f1OdNE84I23FuCY3WUAIj95/zGsv+F
Lb2gqPtuiFaLoFTlSv6hyh6EXjNNUCCD/9ze7CTDmHrbXnrI+/8+5SIBF/77eQzS
JEA/S+blmwKxTvU45WG0PFR1VsGjxX7OgogxFwumPjoz+7WEc6dIo8NGC2gdKlu7
PsI+mXeq4fllPPgLcZ5qtPuw2B8X+akvjNr4JC9Lhsa5c/oq/gNRBDb63G7l3QB7
egGfszxDEuJ0BHiPKnb5r7L+l7rXQLIBFpegFpAnT4NTf+XDQCiDLxiZd4GSYLKJ
7t6rR0CiVz6NptRzLIccS240jOfHogwSmeAqVb4k1m/1oGrRbPZ9DhT0ZYu/GKUk
tGxb8flkLjKew1BWD16LLijm1m7Y6HVm6S9Tdwu9FSMAVU4p5mgVg1miZhGzmjYb
KpLM7vkdTcBsLQimo9l9Mkp7wdTqcnkxXam0GbFGxVznNtJqnv68slvtSYBQykIj
9Otuvb8VTppmL5QmwWXhDQrSlwj1CqOtdjc2f+4wQq3/WOj/zk2dl5ZmD5LmkV0m
0gx20n0mdfz2RFALAq5AgtN95tlAVwwGbRUPbXzSKGdXWCuj+4105LpqNoGyx8Uk
0mdADFp9dCEHM3xggVmZRCK5qZKMKp7qGu/tNsxaoSBkQEEUkM1tqO/Rz1kWOZhN
wzut2oQbqfpPfTTtE7b1M7neFPuv3LL3J20ioTypBGPyLNiwGjawYeOAEmRlbmLj
msIQYZsTzz1reHkQQh8X0lIuUoG00niUrJGSgB2uYnqgVkvUhKv1fIWi8TIVW7Eu
rlX/Zbv1EwYFxw4SXE3XpCPRKsigcH8Od1fWtWwLQOcstzmMkFfZx4yw8LgPlnsj
mHfZbRKX8CVgLu+sUSBiIkgHDbOXbqRNDuNs+CEK7+lr8n1nmxPHq+qLVCHkdGBB
o40lZxB+2uSSxc2h/Jmu45eLHRwrdwXyqtnKlU9o25D/HPnN+U3eHAyhuJS9FnhR
Dtw4aPdl4wJYNhqTRJCxkYzJrgtUhqT7CYFQmvf/00hB1PMmnWhnphsBfDyxAEiY
nNtmef01j0xsZ8cLe+KDhsh2v8IO8yp9fPelwzW8Z6y766SYF1vRhCZyTBS526Gg
h1pJSbTaTN88MUmzbWEb7OaaiHxvTA9NsdAmjDmv8kkHxeaZiKaVBmkozvqGOJzC
AdSwesk7jsk40gZ6vfNKBtfJBhLehnwrRZ82+EDl09zvuusgCLi+q4mjSnRWxqRQ
hU16r5XXqsoPJULxhSV9MABS6c1SaK4iKRPaaKpCtp5wWwKnwiyaX6XECTliGUKR
9K3b0+KwO+1qgxLyTD6Yhs1cSLwBdp5m6E4fp1p8gpOZ8RXmljfYRY92j9XlQQMF
UHmRHVQUQ7PUQ9niiY+KHc4BGa8a7PkSuA8Jggie+3KKFLaDA6PQN8BdbbYjmUNz
f+PBrvlm1i0rMqG8SqYUrEpi+Nb8Qw/NzkzjZNCY2MjIOZni4002PaG1GalMu1YT
dtEcr8EkTmxT3+iIBzEdtcZh1KZpa4/wJlHM7alVFG48Qg2hI3YFTxWc0rM1WeX+
ghEGP2ibSREjK0SklKbVt1SjUEZEn8m9Qw5XZeWQ64CHfeKIMnravO7qzDiVStog
49b6xVEyQi+8cCL5e8vWOTHhyPwjCfqfxzvp/MfuoLUldeNNocUn8AStVS5zPeKX
m0+13oa0GW+phP5wXSM/6dafpcd0OcqY3hu0Nu/dmBrL0cLT3iKzb4JYsUlK5d57
KrE9BsHiDEnPYYa6iYJ0JM+g/iTBlPZWWI7DNVMrOoAS3Tw8oezHY7lvt9peE+CP
5Yg2HTNvHLlYDOZ+OH6g430wZ+cWbdxdiYNM3uKdSOYU5oqBOc6qrQ4lDoL2REkU
LIFg59rHyQhq9ZPrz+2VDf6cS5i8vT+PsWyEjbM+EshOFmW9DV8UpEz5c04+yZVj
sYyceL4KaMhVQgnGpMd0jJxicBQ6Xp5LIU34huB3gpjuh1ZsiBQJWqJnbwvue7rB
mxg+R8eqca43GU69KVjpxJteMAzsaDwIifrwx+JzEf/7PlV0u6wD9ojqNQ/Egkeu
w+kstgwyifGXjOXSku+uF7a1plFFry86RcVWabRNlEzI+La0kW+AkqDGj6cV2gDM
vLUZ8hpJp1WrYJfiiEjmZmpLsGVPpzwvTsCzxatDIv/HZxOPGWyR3jtBXpM6qp+H
LfFg6DkkbLBTpBsdkn8nIrM6NW02RFxfmMOdirVmUoGzzPGVzc6JLYCq9vIPKPWp
n8TYOn7vE5q2Rm3Cu1onbt/WPlTBVR9bjWO/9/JaJDXsN91jepp3y24EkYOF7HzK
Usjczj5jsSSg+NAds/gnj0RTQbmwPwJiV19kPGmjaQpb+gafxory6hvvLdq4KP9h
ySNUq8hpXpJBvcW8A4jOcbtQ+N3U63A6VTelz4u4cOO0os1OOISnLU5HGinp3fl8
/KX05gCyvN86PXICJSKKYNY0lz6Xn182a+4r+r/e6NuBK4Z/y5tXnBCOYoOUh8qB
DZTHGcY8QOMFahHpWba74/b6QgASJQAxXR1PUwTdy0g5+ca5UZImGhJ2OXX8AoH0
we4Mk2kmgVfYpfFsHfBhi3eMYdyOr2pdLexbxmy+i7fesR8j+mA3Y/F/iqZOgZQB
yq+LSrijG4qxny2+8LW2nm/vi18Seq8cY+zpXq2E7H0xXcMQ59lYFizi5p/wul8D
Q91/ViyGRjU0kxHKOS7mTe9VpvAhG+p9DC5QtPEwY0+UeW0DvdtOEGdIW/5OpM6e
f5TQtjE1mUdg9OtuHFQ7KNyf+eF4piakOr+6SQGzK0AtjkkgBz4DdHcnhB5cN90m
TR8Kaj0dg7clNCQrvSiRMQvrvegLnh5FYCZLUFe2MGbwIro9oSdwXIdT6aVD1/i4
tegQ5rB3H0qLmwbU/u4h6MrmoZvtB+0BTIgsBN7gGoCi4Q+28iu7mOj9r35yP1+k
9laeSjmfvdVAXLHt81HF6kU3VUF83MpotKbsJgGtzXQABUsqLH2Nkj+oBspRBSLC
zRlsJzgVw9a2+rZtctG/Au/KjRVI1DxFmSV2Y8Oh6cgmtI+0NUVwGv6eYmznvseO
qqYV13yY72EGMGABvOrpU02J4TiMLBRrE2Ur7I18YG1i+PGw+oc92LhUtBQSHN4w
tOdlS217EmawQm6s1bNBgpbj7AqAU8L8xrxb7eALMmenvOxF5NR9MkXkFI7Aiyvu
YdtVwFa0BQXkOx5PLRUXh06d+NhRQ8f4eCbqKGNp9SxIgXY2PSXRamt7PQHCmEVM
6gUox7OG2xpbMi+ojIffnnX0bqBFyj403G7W5NgX4tE00getYgfZBFIZwo6hbPC6
iv1bzdtMNkOqzFQw9Alvs3MjDow6dCeFjXj+RnG4PzhCXicKa7XV3H56E60dI+NH
1uXtIy7WYf3wtoWj7a8yV2obJaooIB0prjM95kjp7DF8RpkjObGQ5aYO5X+1aqKK
lCtVtLEhWFZJnsOLMQa4eFzJlIuX70GOUN3+Vcw3FpicUVyKOdu5mto9tgngSGV+
brby1nmgf+QtnZJn9OAqIM84oXSPHDJnqRs+Am/IiZy4LhI1vsk+YQsA7sNIg0Hb
3JhXzBAIgKqahFIOkiK5WNigPhDpXB0ua19EJ3q17Gx/HBubet230XpGK1NQsV9F
ZdChYGYHgSwQ2vFnqk+BkoSjn0gZ8L6WYtTINuERJTZilY21k4tKbnzD2cFrOWg0
lfiFYpygsSaTcIN9OIuv0DfT/jdow3vewri2HAOK9gEAJ3HDkAN4KY/PJaLMeVVB
y1Bjqn765yTXV6svmvgHllBA0JktOsj439a2mE39asmq6LJEXfZ+Ia3vcbczfCYt
nlf3U2DgkC4OZ2+KDRrBMKeGZdJv7RJcmI8K2LlnJuLnVXCtksRJXJZ8DS6Z2i7y
VeNkbcttFJUaUgNmWCD9AnFQl+t6+BZmQ+zeAg3UUwnb+YEukcn5u2yEgXUskUw7
C2ieySXjYyFkSoLfi2ye0fAf35658fZouF2+0Cb+sq/2m5aYGMvq1wwgk1Cqv2vc
TMW6ZvWfleYiapOQuk4DzzMlQVgnFKB2l6qPvIrh14uNE/LHgJfWJs45tMtHv/VU
uB+pYKwqbvbd1Li8q9QmZTuPMREFGkq6xztz7QGrAGD13x5VQN4Sh9HYXrIj8mGW
QtWzzh6I1yAz2fKE6Jw7hr3Qg1/Ut8VXq6kWEJgziKMlC9Gc3ZG6+r6E8zr8Vtu6
iFc9HmpgghdQtWEJjTkjgqid6aUhgMQuCIQwpbCfUtXTSSJ02bhbJC/S3nT5cc+f
MJE7uPQ91QtYTp6/aWAtBlrECdYzfKR/iE1+oGh5Dwl1O2KRsRRJf/m05zLPpfco
Ka7Pg5S1afO/RCgA+ADPQnsQNvKFesM6QrydJuxrpun8XmyXqdtyRhRXN7X6Jvna
EKn54Q+K0PDHjfyYaSq6Iv6hb1pXg9bsuq4d9B3OriJ1Nw6u5nz93lWe/sDAEPza
GXDwaxlQNgYlCJhHAT61q5Nh1bSUCip2zE+T42U1gZZ7+Bpqr8YT2tC8Dfj59XHZ
V2J2zHjeH1ZI9LvGY1J81dBE6FCwpaSTu5R0lMwSqt/2NI5v/olXmx9s+8EugnuQ
htk654MCc7Mf5quB3cKx24hv3uPpp1T2+EhEKu7qsa0VwXBIPypWi8uEf3o8FVt6
DSseHAbB5cvwr7cJsK5t5tL5B75NL1kXNlhEX6rcq4P1Llsrb1JLiM+pkg3KhP7i
uxWJBtFl1rIb9Q0ygQqfK2Dwd1bCcMswSlDE8ARH9ufVQ9z52sjZk/b0/B+Ickn2
EamnZwFVOPn7ixixNJyIE6JiLbvtO4QLJ/2tgcfTPe2M5DcplPtuMnQ5xjERL8f3
2REymnY3frvIGkABU4DWiOg/8/NddhBihGAZtImnzV/v5cJdmp24aCOnI0KZP9LR
crXoIciHnNdWtXUJNiqAwsTuOyvn5I4ZLtCa63unk3YJOqtmzDyKrVBB4OIzreDw
oZbiMksdZr2AlOIge46Y1aehs3C1wtWxK2sZ2+b0PZJH7VfHghTx9yWOt7pOTkV+
IplhWyBNj8eJES4TIpUe6vQcpZ/CB+2p6Dnp7iAxjHiLq9r1+KYnoW41lDRAhDOQ
x3HUcK+qZTbJoAdBBqaKAQwR5Ahz+oqPzhMg1/0sNcbQTXT6MyThywGJZANIGgjJ
RHzB4W6VE0uSJ5osyhDDyC1umTzAtoETpZOx+Qa+canP3R3qRfHYEMfI1lviBope
dSP653QSM+Tbo+2FGf75WoxKe9GFJaXQ8pnDuSrrbYkME/mBW66jwzXY5eyhufit
99UzMrER6i3N6+9beDnc731+Q7jfSCMXNAiWCFEmNvZAMlYxbb3Srzo6F7B5YR5Y
+6oD6yJhBnJryuNSPfi2Y0+qJo+rAmaf8nxvcndNOhoC714mhkhGrI8HOeEl3Dow
KDEp2pNbQw91zsYUu9GJz7qcYjf9YdWx61r5S8KTVXHWPr9OzfMMgdDzNNuRqk3s
2abvVJdYjT5Px4vXA2TFMjC0UUyYHmT9IuVJw3P2c2EBQhQkkz5tPtiwECuXMB0P
5ELBjBxgmdVdXAi3tjIzXue6cXvRKg8jT1kWa48witInQ3h3JaMzuyRP1scXaPii
GtlzMK9eAa7+kQ5dHWbE/ibFnZboc9AuUTZxL56iAYFSxmj56YY1TFa5glz73gqg
t1O8DnbR5Q2UO2lI2UMAYFGnu2scmHXd6tPJi3U+tVa0OM07oo0d9YtGRbW6UHVy
WbOgQnWc1L/Fuk0OhEhX3r5gSnmjfbnGiS6wh5aqKx69bx3JoV7uZfzUyQ7I6wsw
oT6I6HlNZxpWMHLrhYzsCQ3ivDA2ZlDis854zWyPmrEDtcANfiyXT4RwhmWIDrsb
uMnestB5uvrCyNKyws5vfR0Xxb5WF6WQFrAtPGCg0h5DbeAlVgUuNlD9FKLQau04
lnUPBPbcf84h0nNOB/ZQ6U+P/1bqssH6Aj8qmK3mHa7xTWkHA9RTzEPnQB5PVvQK
3kBH0N2cz4mRKGXSvC7Ip+5f8bcf1PSzxT0JUPOKA5ykLH+4FXMC7fdlWZ95T9ei
Qyxut0SuEn22EMzY7ijyQ22fN4eTWCYnaWRZL9wPq8RZ1CMs8LsaZO+gtvx0q864
F7Vj3m+Dgu8FBhopn+XJdTcwTGLbuszoUZ3bLaX77XrEAPaVlX+/d92jHWHW+c/o
FCFflOz8QWFa7QYxb6D7a7VoVfA3XZNbS1jFEUQkpoliorOHjayh3FpRn8ddxIbq
htbtYvWRW1IfuQvheDyTqbwHjlRDbtEd0g4ljkRrYqLR2GwhgJREQAGnnLTOe9ey
lOCLGpk1HzRDEKJxfbK3v6JHKSxEAexwFk9aYuU7zJ5sTDkipT9h6atfzrKBij5P
7n1NO0yS8WfeYFlUy9ErCDDGrMwWxY9N2E++Lbvwc1HJwr+ZYRbt9dhvwJcTtzII
5gwOTa1AzIxH/oGHv7YwjthUvphAo9RaWooxZty+Tk+YFH0B4yZmPjqwv3WrtCxe
TE4oNVNRWg3wsOXZMXm+SA+4KW2hh2MTBFiCxfsvqCIFR1Xioxqkr6X8DiOBwD7v
pq2sH9GbpIdbSiLLao9jJzphyYFmcquXcEFiHxd2BRDLUBufLovv6j7fvmIS84PZ
BtZivP32V4WNVGsuLQ6H3oEXkFKs7P3jJuQGGZfsrrVk71qWO7pSLOpl7qDPqFx1
dFHdPtGo8JcfENMW/dbWJEhY5xFLE4KNnB8M5lBjyo/rf4xIZYcK/xqCl92HrLBC
gwNDuAYJ4rvfqaFhekSPYRUYuEhxb9EUJ0+Pb2WSHZtx4iKcPagaRaucp4sh/Xne
N5GRRrzbLHPLPmimxw1aTSITeg36V0oCXHt0eMkONaXlbOJoxXeXyiyOYz2otmqh
Zs8Ke+HCR1MyPUHsJZ2Xw9S8AIJDC09H5p48iuS8QO86BOdtGv/EJQzzcwA9vF/F
r6/7vdHyYJ5ux7zYxJembCcA2bVz6Gt3Gyt4q8mwDUVmwZm7SGasjVZozNJ2w3Sp
0ejVfQGhftoD+Croz10WcEhZstrBfUA2i9X9WrVcU/c2m1Aic0V/A3SaevJf/1Xc
pw/ZqyEZWEExtWrw/LzW/B2BP4iIpvZYDXNCt8uS25vCqK1eZWU0PdP/spj+QOat
9dOFV9nc84inLLVQXZmZ+UvXSODyWuujDUnKgiQQbgCy2chUce/CO3/A43ztZa2n
ClWYGOMPeJEj9RwutxuMU3RQTQmKJH+aGx+uq3oSybM+9ZIUz6v/I9SimVxeWJFH
K20EQvntu5tcSfQIlX85snq/3m+2+BLQwwcAmFPzKQHlHf7yswiiwY8Wqc03mUcZ
StJSGznuHLWiSWqVJfNUL6HLkEzHEuIw+PwhhrlpqG+1i//q5Rr6ZHNjc0uKyxzg
X1CHj9S7s7vB0S5zEBjOTW5/OQOXvEqpkwdPb7jgGWvpMv5JlO0LXeLknFDClIuM
ahD7Sv4dce24vz7hMgyoJrXeAFPik/Az0qejzOMMQtAA2F49GvteDAIkPY0r4LT2
I0BO+lecdMRKS0WFxgofb96TKg7Gkcmgavtf+fPiyYc5fj13HqRB0AT1u4lhob1M
nhLMyU+gLlhHlYKYbrPewBDzJYq6BsKnkPT/jrqSZTo/Q+pI4YBICfB+OXJjmZm7
nevQWm0ijow1JAjJtAm3Jt3e3Rr5WbCQ5Tqv9uW1iJaBMo/s+KXV02iz07v6JrVD
9P8vwpLceMQOwPNiyDkBxqVdeuzp6HeNXSgWActiotGQjyU1a2SkVNhqjuQRqbYX
NGINXEb+H+Op/ydJ+TiuMM94MsyFhGmaHJyBHpeRS39pLClxOfT6FX8L5cLkdAjy
dMe/Fz/2+xeo9ViGOajQ0p9hwm1+v8rzkFCYNc+8L1kHo4JvZW37qWeK8d+pb9M+
+bbfi8yjVOrB/wkfIOiRPq21scxs/o3lMD+mEF1tOtfMQucibYTNEbfa9c8LQSG1
7BU87GPdyUO7yCf9j9dMCo3E2HbiYgnC9cPS1cpMI6A0Dj+ph8S0u9LfKXWajZD7
dmNSBCZDpefgKcd7ksqUoNtbE3ty5L7P1p96MwgcFkV6g1rSM0yhGpJqdw/rigvA
OmAUGHCHlt2mZ73sY583W6otNGUy3R8foENEopy4cg9zDMPYdwyvfcGcHNUp9XWr
9j+FiJ8YUZep1rF/HPTzTHb3f3orRxdt0rnUTTpfgzuSn6GCGxworL7RZ+jJ8P8O
TedXmOg/SkTw+r5HKAncHH+sP/iVOKNMUvTZgn6p8u85LO2NuVOChS197xpLP+BK
IHDVNJwcnUFk20VjUspUlLC5c4ezK5thcQY6e83XgnSGnUGTTqXV/Ak7Iq4Nume+
CPvRK0mZPH9B+6jKR6wG/WaGjwz0ZTKBXOxaqHlCRPGeNTqczOjmZocl7szpGcdD
0+88kheA5m33F4ECXDauWkuWNscoITnBIxLG+HOi0ORp2qPVELrtnikThVr8AcsR
YayD3XrbjW+Ud0KSdustOdo8kc5bj6ONXmx0p9SafN/jmwyIREJ0w8odGNiKWzvn
Sqo1wrjwx+ysl5WJLmtYgnVT1LulawTVj9xOb1Biw5Y6uCkOj9MFqDIATp+7hDPt
NhthEwQUKlM4kZ19+dh4cPyx/mRwjsCsKi8XmreXxsStavlegNhKSpyEuNxxjz16
wRmVyDJx+itoKjy/N5sMOiDYTKeLpas52iSpaTWWhbs3jUNa+ywYJd6l82BHwZbG
/B2J2mNbxfzD9KVGmtcU2FT02vCnM6T0U3Ph5PNfrs1AGQPdIWbnjarCY839KR0m
60UTYC6zeALlzfXq+/DW9f/ttHXyZkTfZSDkw3OwP95j7kHbRZfnsighMlKiKAXC
ILL8bfWaAu6HoetqP6nH4uGuY/GP//mjJZ7E3jy7Om4XnrES2g4qXBgCzHXJoQa3
f336D1bMDpIVMhllKeilBdRlcrW17wiY8yBKoZ46X3L3y6ITdpaYHeJ3eKEwEn7X
EvW001u9OUrlY0FMRdv7XCO5V2GqNFPbeHj6Xf+q52KV3lmbWk8nk/7N1CIhfl40
pYnAmuo3XIFi7bvX8eCf6+ENnt/QMIf+N9V+0dC+zH1OEok1PvzuElhzWGQI4ORL
SifjzCae7nVcQLdSLjtV9BDYuhRdCuS5X4FXzD/NMLLJ7NaLryXCmbFdl1R1/L6l
7sWvcqxI2kHR4pktQiB4hG1ZHShQ+zl8w2c57HEyiGsy6cSAyTSNDpqeBva1pNX5
pxk0TMuAHg7ZC57lGazem6aKBnlhw/IhQ5/PI4JPohh6fW31pTkOMBeaY2zI2mz9
UPOmyxQUerrQF+hj0aVD+K2mUu+91mHBXAC1rg9ZT0Kk9HO3ULuJEkDb8eoYfQb2
jMpKmUc2yi22mATsQJNusR9MIVPjFIQeeduSKZgkev8o2G7umcffCvNyhkxyL/bG
M1T67jXtvWm2fxyT+JgROT7i4yBOmjF52fkdrVgSl9VALLoipXGTdD+WYKmIOLpB
5k30iNEjHh3gnD2y+6pDbhAg/nGBiN7Uh+wqEAJJpFhn0Hq0VwVBBK67FGWz9o8Y
WRcvxWONfjlJEE8atwqHXMpTHDoGc6gBexE8SCxfh2x3A9gdi3eBBhPPEqIMFB9p
ZejEKj+k5ssX9TVHGC630v3xkNbyHJigoQJU/no916bjclk6s8l1fIk0W2QfLLYZ
J+nL2vW7potRtOljDjr+mOy9SbKsHrrBiFi3tCZSg8VbiveZqkHRBAhYQZgga3Zv
6+/FqeIPPlj1CqV6oZ4j9isK7mdXzSkneXM3zQmG6noIJWC9N3tP/qPxQZhic3eA
XxKEXaV9H5Dk4KhlA0Se8sAYl3ODixkSKjBA8cFtdb2Zrrk/x31m9xMv0w8hQrvB
akJmuj/eSP9C4gZ1fUWAgO+fs0WiGecFg06qOvhHHEwxgj9Q9O/jx8hb4d2nk2w3
1UK2F4Bl48ztrdwbi0G/zzfkalPaHETcMX+THL9pJunEbM4XPmKDBKPI3c+s1L9a
qt3H9rfbC99sBxNcqG8MUJ73EM+3Z217a/ww7YgCZi5fZlxW/2veRWZUDA0dSSLq
mEHFLX8RKOo38GtokrR8sinQyKmSTZLaBQuKUscwvXW/4rDYUR/Lp3B15XxP75nN
opfSN06kJOPJhR/+DRaIOhCYmNDz5U/JFsTMSZeI4o69ib0uXm8K9+ydRRkKR6oQ
Ih3aAxm36VXQbab0sI7pfzMWJRTZokCwcfgf0qk829CBzI532KHj/AeuWpFnK9aZ
HYTVkcIE8YxlgSFcdcikNTrVvryAhu0taCcvA/snSXvkeFviNUpRy4YznjSwcBT8
tkU88rBgcbyxBfPHubsI/vbiqywnegVTLTm3KizTfUqE76uNrDJdNYiPdfczAPEO
VKn2bwdb4L+WrJP7B0KGwAE0PCXa4PvK+LXurkD237rvgg6wtKcxQIiSBwGcPHbd
ZwCF5Ehrg/JrXp9Cz7vXJ4NaO3eLfdnARhmAH2ASyy0H/6Ng/U2kR2PDVlnwKMoP
2YWT2o8L8P85rooJOF0D9g1g8bZs0mWld1uRLeknWiWp10F18113RP2bK+roqXV+
eS9qxs5kjsemrYq/xlLa4mDReWU+H2EYP2TPs/QoqD2ajxHTetvytE54wtuds4aC
sUakH1KVg3hHjcxmWtuI5bFRv2gTQXBxdMJfSv2oHIp6FEyGO+wmZbcDpJVEVWFB
BAyedFG1GxTafuX3+0txnI8zQvrxWQbQh/HxbMHUXzpAc6Aa7btpheuIhZr2IdyJ
KTas/y8t+J1Ieuh8JwN+tnzytBw6HF1mmwOpXl196JmR+Hl1bXG2A+fHZjwCAvKH
IMs/t/aEzAVwfzR6xkVlhchgVyqX8XQAapbp6TvkuwR2TDFqaPVjFDv/vZM9FOlD
fTtB3uwBgLDeKv7lIL2qejlhdoKWLc/U/Pu+t7si4jJgfNkP6TwzJCFvFXIE/JBQ
5w1CJKAPz97gz1XR4FjknvdzelPKJGvhoRehAJ0XKL/3iO+oS8diN2caS22qzQGy
bWKGuLr4AkLG2QIG9Nd7WtRQ9v6Nq1KlX06DveD4v0bds9RGX9HJglWmVspEnIsu
WYbBfDcjuA0Xvk75WigwRjh5/WYbUkHQ9nJepse5vou2X9LRFOODLM0SfPBd0vXt
qiXA0ZhIHmt0JTQkVvEfwOaVJF2PyCEhd+QzHrT1gO0WMY8TN3Kp54D0rBnyAhI8
7glSwcV8+G977NqxuCeK/1MPknZZO5ghLbnblfEcwCIeHpnh6l6kybPPm11yrYns
R7LTtv2Fi3WRHwjx4RwG3iq5S8G08cNFJlcc4hG5dGy2JS+0txtqiY3ocahFa8Fa
+xODzHquaAm44nTqoxicLz15XSZYEqf/XjtQhKGfVwL4rg102QF5BoRUQ+0tuQOi
QNwS9jK1UJAA11p0D3NJVMbbCMvinGLcpAGzqLm8DFZbtv/dYH+CiMCiJ+BA6KOh
n/TuONMfsBAOBlaErmYTQgcc6KUFn6SRBTBib9EZuBuMvo/YELOYy1GafT+zDgsJ
R6d0txcj5ODoY5BgrWb1/vGa2BG85i2QH700AueLVEcX/uOlvicjKNTkUs8Um4u3
XAe2YpmhZ5M1SdzTp16xg3GGQp+xRpq5jCcIZHBgdw35o7E4pSGSEERoXCpCwTxc
NKfZuLHMBySZdS7vr6daZUUC722avnbuOcHayPhBcDayWu5nzWhung4rSS9z4NmC
ljsDn2VxhybshxQC8BaglRaaqEHLJxiq9a1KqIMhJtr92BZe4Dwqa0Hl8a8BDESJ
/tiPs6aWPZrRziJGyM4+9GjOiVA4emj21Wn3TJyN2VSU4MePsmV4oROfsZn6mO24
dDKbPfZtG1OWaLe47BxupUpRXNmPdWBDI3PTZwhGw5yjxyOnOWFZZPoQxFD3zRVn
vph7Qt8RKqBKmtzaSYsCK60bhLuyvUwCEcswncSWC89hLq7GYnsjbvkX3rHH20Zh
AbtXIjHZf9Qb5uLxrUv3IqzNjhd4jLy0UOsiRkiwCm2i4EKHj+iLJ1L6KJPk5U2f
hoAQcq6JRVVh1lmZKwDcrC7X3UBH181i1IA2sy9HxHYhkVCKRxUxrQpLd1iiN/2l
uhNylxTUHZh4XxAU23gaYASaGFm+906ZAWqwLffU6EXmO/CZ4hFs0yuEf8QwHilf
7Q2XQfmTvaSgqrVhqTkb2M/DcIgkDVjITqwbSzHclRWKwN18iGJn+49CA0XWplMb
KVG5FGL+jFurCUuWbkf6MBFEsw09tEW4xambzbujfDJtnQeS1UYx5NIf+8O2zqC0
neoW2zeaRvPjGxUU6a5z+2VGeP2plIEwoJ3/ydsC8b847EYO9mT6HbDr5oPwJT0U
qsMvuIA2iuJU6a0qvQ37ZVVJQXEmfLmlDiLwE/IfZYr6W/TTNt7OhzIwidqV0iA4
FZP//hSkKUrlmaQexxVHokZlXGKzUepr/Sps2DtsE0Y1WMntOt+oW8//MSp2VYGq
OsbPUpO9mWCr9vkHzbcsrECGtwkagz/Y0RmPwQH+pJwPAUzkYK1xYS0TbQHcb1sb
B2BscBbFvqH55uaeXFZJzbIQTnvpGttHVWLsLEiXTXDmTU5AemAvO9IlCpa+nfuj
MyhEoaKezK2cHPq3/b/EPFxsbgV79CXgwBMX4VNwfSYue+L9ZN3dNvOq21+JiQ44
7QPL6dywXti15vrmO71KGC9mtNxOqVJGcHHubfqCqHxJOcxYfgllHe6gfvRpV5YT
4PXJYrXXln4G/mY5gJ6dUwFkC73HTXSdoCjDl0T1ktAXngg+owJUrFJb12SZXEdv
eOoU/0nw6fsikkd2qp0TmiTel2zNwqs3YxGDdXPxLa/DOP6dT0hyKrgt4tvnwZEA
EYNur3aYwpO54TL/2ahakX13btDQpbeyNz0mnCOp7hFuaaHVc68ELmKHDWknECM3
g1qyUK3s1cD7Iev0gA4qZH01qsegmgougwIMRuFbOYs02VNT5kaW2VTeIjb6+Y6Y
vbJlVgpKr0lfnxFXNmynpnzabHgqx5oO7cbx52tAkG/oGW0amwNQJGD/+LOJqpxg
PQM8kgPtKiedwSD4UL2J3gRhIPCfkVUFpL8tz50K8OPT1m35ReP9hyfOsksSLLPH
cky8pw3o4D4iZOj9cPKS+AksSHgtjnjPHkClPVz1kQ077feUd24c1m/dqjJlChUE
GRpRd5upKPTnqKdAmsephJS97GF+LBjxYIf5FZyQkDRcP/SIw0NzlZTWN1rr0MYv
/V9YJAhM6SZbYCkTDKPyTXtFjZIws6uS1odZNnAQc4UD2ISV+NIUVNWLbskuSEGM
82v3w9+VWw3I3ud5tDDt2mhQ5DwXE9OvqjDWDsTI0x9DSqUDhJNIez+JDZ4lO3Jn
wsQ9MFUJwG0ulyyNlhBE/YUSFY6z8MBH5BxCe5lNzx9LrL818IHzZfmTH0mli/0y
mGdhTMG5A+xinCJiJ9Xt3xOliGxtKOYYKM6wKlkv+HvvluJJMGH8XXkAV5Cte/xY
edUmBloDxq/md6CFqEXuahiirsIFmrd6xG2xuP08dJ8XKkQKGPcIz3Sa9IFUEPrW
dVm10VaBKZlCXbKSh+7SLhKma8KWRexTctN0jb6ESnDK+O454ioEwDNHb2FL1Urj
3qpDSXYIyRdDSmlPqX1CoDTFt3S3avG1FvVzqJaxoKDL4nPyjBTw4OcNEfJsRPO5
CYb2qR9uFlNUvH9/99UWx/MGUHAMnlaNux+/IjNwcgJP+IijgNycxrajMXtSOW/S
FExX2GIIaYjehreunGQyVAvnRItBVbTqsRbO4e2QyBX8AmWxn0u/ljnjx52Ivaj/
3WM0IaCCAJaf8MwqKihmCnPd3RJ37aWKP15ap69T7DXXfsYn5+2qHPvrlE0cpYiP
D6QJfsedWFEPbkO56yQIz9xtvXn3zyHXyb6DleFLmCULVvbojABcNlD2IGobI6Fr
xlRKch8xYgFeeAsjV9HJuRQbYTJUFpZ0i47MALwLodyN01Q8V/sHOyOd+0Eg/vn6
LaYfjx6yqLgHgGiOGkcC5zbox8flPPRyOk5RYJLSxbPiTnx+P1HmFOIx2O+GkMjB
EGRSNQbKpIXHWF/QEYPaTR2kva2BuvVNjEOdKPTKlrmmIQgOhkjJsa5DKGt9OLIG
tzdAhwpsr7c0jes9+6+bG3c41tph4z6V6mjpWnPbpuYLULTwxaK7FP7JO9uW6sPr
kcbNK17yKqKLtVapso+lXI60iW5Ubmy08dNzfKkyOViPDZT0fw+L5u5LY86DByvP
Vua7wsUO1/afeJ3HFaoUN51YfujRnlkRlUebBPUEMe0M+Yw2Z7AwCy2wQURGOw7p
aOCAFKIFFMS8ZwnJBvlTlgqF1GwYrwmm+JoRVlTn57McX2MqKrYfqqrCzFKIj+1J
lhRLkNTO9nyUfovblMpOMqoKDF00MnVIXu5g7GjZN2y7Q2SR4xIneV1te/GZAKgR
Yt4dB4pEe/m8hUXdZmbm/7j2eNDOKa8vJCUqN7rmyEc7PLiBUPK3l7qcZOl09qK4
XNSl+EZU/wD8vejNPEEVRzm1Xxte97xM4hgRyut8K+kIzKWZPWRWMPHYVZU9/NN0
e1r0JeROKuWTW/tqYCfhADHrlnaEr6Z+NuSMHZd5Yq227Dd+nHLYDPZN87GgMXWR
bYyXUkcTrCgO70gF/MBXIth09SlOUWsswXS2giKsXLhMM+Vaz0q8z4h1L5+SA8zR
D1oZH0Ah6jrLOymM2hSgg9Z2cMVv6iz0Epj16B2SjiW3sS23JJzv1XNOtZtNN+np
JUFCxOTSRCoQjXZzubNuGPWYjGzisK047cr17/Qq5T2+K3Xe7ZHK9on12YOYwab0
8NuxL4d5g0c4nW4GVYt2KP6Yr2LH94bbVFsRTXbbp6empDoXoN78a0sPQZaA682A
Zy7XznfeNG7Fh+uR8YDVX3yKA7shtZKv3mL8eX7mVojygH/S2l7MMClBRTuT9wh4
HOtUm8zqcspBCv9p2CXOFK4r16ppElIhPa1oBeY/dwh5AC4WEbESsBmKSKJlqP5B
dI0oJzkdATLaNetSYZqeRmRHk7jfBXug8S13PmJ51LtMymWsA816uDen9N3Nabzk
R2G+ubynNoTe+/u6RHE37ePNaOXSd5lFJZai0g2vmoB1EO0sqW5FVqbhvG0mYy1X
pO8YOUZeT/yN4MVz1U2YHoeLMGshS1ruZp+0qvGh8FSzBXg47dnAnA3I7D2j3Kyt
tMgV5fLGjcPiHXiCw5ZQb4cAYsgj/wLRTZDzM5sVrXylI9jHKStw3Dbl1eIauYgk
KXuXt1CT04Av/HMUIIFXy2uN2inJ+vwyknYIW78NgvJN+Qy8b4uL61eoAzi6MmKE
T5qTHNnKFBsy4LPeyHkcffio1KNpdxB0Gts5e8oJszBRdEj8l0nmjVMqvpSmbL6p
q/HbwbGgZA8gTN3Q+lyRtsQsJ2VRd2neYgrRa8aO94LFuafXy/v4v7btom8LHnL+
OOM8VH3dmITtDYhdX9LTY6o0IqiFil4K++VL3TGlBHlI/QG/WlSjrRLMNjGjeCVk
UhRlAOyDSyYuycMAP+dF+sE/L7xVlCrOhiZfKi5xQiayhmYL7xvfQP9j+8+FiI8H
Op8zPE4mH61s/BanodynWL6v8yz79n76g+DEFQkEWpqQ0yDvSiUzQklCpOlWU1Yp
1Odc8T16xtL1+6iQe+xAEZ/nfmCMspAM/eVroPRtG0sFVou7LUuiEYjyvFWGZ5FP
A5wKCP83ZkEraghKnW9OLTH24Gq5hFxbEANkfmEIHPQcAOoxpfwMYR3alltJgoG9
96Cn+psl8rYm6RIm8QzqFqs5jpiVxU4mowZm3cm6qoCzcuuNi+NfUvKPUuo1TEa+
CTKyaS+GA1lXtxepDCSzbuLUDsjv8XlikC5RvtDkzqX2R03Fw7OwmxDZFQAA3oku
6O957iAt61wTHs+3EiiIWAkk2fURGv8L85xiYqyfyDv8CLnqOevrLY/NFFfwLil1
pzjA2SjWtxw3pXpCPDEqkZ8TsiB8b+H7+gs5f0Gp92Yrzvw/1PybB3eyuv2IOkSM
FNQ0hR48BZmmIADhjDqX+78VaRplmRCxdk3PDuiImp3TUBB6diKNEedrKCXE8Gnu
0Cz0IgIWUgSMqo8u1OSo0Z+rUaQx4pcMoLlL9JHYftyMcvRiEQfo3ncn+sb2kae4
Ylkbi7BD7xRBTtsfwCqXmTWxGfA0ULBLR2Qve3UWpdY3Vy6aSSwPTHGoVRtR+RWB
L3Mn9G1+YGV9ju2v0THLy4kahXxTiEsx3q3glDyn1t0i7Q+q11YanMw07ZiySfOd
rGTcAdSWbDI7Gsw0sqpWtyUhp6VglL0ryuTj41364/5972la/YoIH+D2nXANVBrD
VmTCIS1PjZkv2iEpnaGe85qhrCk/OTW83V17Izfn3lEcuLrI63mYYBF7DoxzQnKo
XkDv72AR0P83e4HXMXGGVtgaqU9ua5fNDMFPhFoFGPSfdy9asd+gFnh1gLDkffxw
Ei1K7PLFxykkcKp/NH7xMQp8eDVEr1BeZuNR5UECbvA+7OscUnCykBQhIjUTFlWt
dAi40+Ynvnk4zbIqKn3/eQBPYeVwwhPZ/RU/Kh/3PpdisQpIoQ5NKnge/Qe2c0op
8vamheVd5NabMWBrKA4am8Dpa/jgLomzQrsp+9qF4r/yzZgAfYukjpAwt3+5U39s
BslcOzRzGeZVHjgff2eaV8QZ3xkb13TJWyR2JMXbO25xfN7aB+DTlnRAF0yDOyqN
jIFr+4EQ6T15pJtE04mrZoJ+Uh9FzlK7ZR5T+2BCNR9cdeEJQIl6edmGaJKGPxEA
jIuLgZVNvFJUNfCLmQcDYWZhs49N+3APC67ghEMiWslk6Hco4zEHomljtuhvmPMp
2bL1JIRT5QvSFvM736U+iDD+X3Z/PynZ8CFy/cbC2HieiGQg03RX+lrjrYGINfZJ
0DVc7C2DbAxlGnthrs9IThlwezau4ASiM+l6iB2zLNMHD0AKjiKCtCKPAhoX7cE/
dMT1G1ZiQP3AV6HEV5ldE3sInh0v+LWUkJLujGtJedLMdRBysuUEse/0qleunPEz
GrDAyLJavSemN5ibZ/9Z8TdriTb+JtSKP0bi1fQ/b2rATwbKx1YSOT9zvHUd+30Q
tBjIFFL9eC/GL8UCjJdjoTeU9trgYlx/DjhvRedOqt3to8YmoiM1wQxtlsu75l03
z1ciFojbayAO3uDy2qo79sTXp3Nb9ijV5YsR5Q7xFkpUh8uumzxJJ5SX6VEVsJdo
DvtIAQjgZb15VckjuznNJOVM0eBZ7TcVmyMYWLbXIJRhQXhFBXAW+gfDOv/gIxhz
4wLwp0n0PJwfdinG0qkFPMeSld+DbHv4wO/Qea6NNFEk5uNWhqpb9yvKzGzpE7SX
M6k9PkDEzYLCDgW1l0quVYjl5Kj9zVnla/ZfwhGDx0WGjpFsomVaeDg5h7jlkk0A
NOm2CJT/13I3ywMZVwDjjoCuumhsv03uCSVrU0j+vyvA4MlrsMfzxHqAA3OKXCqE
YAFsovTDSm1Q0u+nDR8Gbp37p7xsUOeBmjcBzIAfs/g69Vido1hIQhfxHMoZTEkB
HI8b3UdZg55T/1hpDMnyCUXuQrMcwxvoiSgha4t4KzYBnsULOF7hT7NUg11TW1GK
CMmQOkeuBdR2eR49iovtkV0edO5OZiQWyZ4HEVwBmsxZYuK1B8rSEPPvd7annkjy
2Od5XAxza4KBAUqJ3LgG7lKrdmFfelAF2DhlAZcjMQZqLH9OLTA33Ux5h1BGf0lg
joNolbHO0pj03CDAWWC+xHBzYgu95xKYj31F1O9C/M5y8hsrRyz8fIiI5bIPARqv
yel0YUoGmqkTzLv/8O9hjvWHxyRiy36WUN0UOhl41RZl4eXLZEHhRqTCdPOavBlm
RKRjetbD3N3OOvp99jH9YPxLEFPQory8t8zAiksmf3/KeLe3LTrY2/aETycVnsFi
lVDFnVcmj6nR7ushkwobbN+aEo5/WKM2RQ4KpwzD/UjvdZkyWAL57iORMq5EcAnm
JFmk5nXAsELLR8ZkRvtzTY4c5vLWPeYAo7ONbHazWBto8HQIQ8/uLOHmenPAE5a+
6QjuahMZ4i5/AkOpitB9AQmmkvB3UNcfP3a9p39JhD2sDfscgGvmg8kybB9pg+h7
27W99Mo+7HjV3+wfpEq5Y3zK8yPNrLjOu08yP1MTJE2AinWo6ng20sc2FNKCqHMh
/hVD+4ckpb+ff54ZQz2lhaf39IyrXehzcLm15IpY1CIZbr5WGHMmhM+0EhHtVH5H
YX+KgmU2WOHk855CnFLRgSm/eNw7Bt65SrX0l4OZ59yZUHdf5B9WrH9uk6YbIlNE
rH8WNPPUjQUJGQ1F19bSd30bMMwQfMpqo/YugZJKh6py8VdzdIEdpmCt2rL8f+qW
PwGfDwrVXicY7aX4lLhfLq7wiMnDN+P1fJXrHlP8bq0RfH68NTpdljxAHSgeuz7u
l/Pss8mtH90sKZQq0JDR9poGZOUeU6bQyOQAH+zA4ZMs8nkKN6n/1/PYZSpCIp/i
8Txf3yC8wXCVfKCx+nTe3Whfzr5CyoZdlK4ou0+cR1WDUl3Cd1sOflhXkXs2wFgf
MbJN2zqLGkAPhIrFOfUgQIlqkgo+2jTKPm7nQAMshSYmcj745UtDLLF4HnrtgK21
EaxEifjox2zbc7HnJ2e4xJqJknTGdAbCouDmLiTIZ1jWBpCR3LHzf8+W366co36r
6lHaBSMEpQ45JWFqOXV2sAx+ngY/7B8cfYVc3wgunnoJwJASW9LPcm2ZmzO3Vh15
6BMRNSZVlqOvld4rNDKU14r/qW5tKumTAKF0yGQDO+2S109lf4gGwxO9ZlFfGrmV
Jc6yAPxPqVGs8rOPVSC5BoiEAX0LdxOnrlRroNmU1Yh0Bg3bHNEkPoLLiaqr3QJP
hw7ZDRk/+JGZl/YKmx3e5X0I11Am3YadnJTTEgrRPdEyw9w1lJZGnEb2WYLquJKn
Ajv2q7OJDcKebEPgP7IEKikKWW0biXxQ0RyNFLTXSzOnSGsD5dmhRoHwniQ+Bhzf
+RJLSe8LpPLVQAk1v7GfiG89mDoZgCX8bafdV+S37RSxWF3znDAPpRwV0cpLTLhG
eWVo+JC//3iJ4XITyjJG+3w15FOmRRMbaqtEJBUftSU5BMiirVAS9zwQyr9HZTDg
Ff8WiajZpJvziyVYPiVotJBXhNBrn1E6ZSwBVHwqVzYXvGlzRnrFYfQDfkc6w+IM
biUi2D9SlDp1OYXhta2YnshSVkUcn0NYbisYtDXUHj1smEfoqoXqCHaAlzGCLnno
ZG+BG99F4VcbCchlsIRhHgyhNx+R4qT9WOXlP0MGva4gJ4Nf4sDQ1xNB/J/llm2g
8/+VdvwPgwEfNEJylJGIVma0qA+/B1dJEZqUA39MoQbVuyDXZFDpJvUIYiHVtEpW
1rMjdslGv3teJCYKolRgPi8ez7MHbDiwOatDDrXRT0MbHoRBNUUuNeOBOJbFQcKj
b4TXEdx0cSJK2fMFMxc0JyNSaNxQb8fP7n3l531NaalCbvxP9mXlpVcpMQxZsKfE
qGbZTM3NpBbctS9I0D0pnksUFFzvW31i6FBOJsr25ihOBDOIF7dFOU9xMkBI/8qh
q62d2JSTZ/bfIXbkNDcwswosSN8ex29dybshpm7mMuugDa0z7SvF1eXgtVsELIwS
nO4SKuhterIygM2kctt7SAPaS2Y59xXzvHQF6o/PJQhpAT2h4bWJb+Ttw6/SA+Hg
ZKohoz+KO15ruDabdDWYU3MsVh+wyBPS+Q9csRfkBC/ZvRPQqnCVPqq5LAv/ET4H
sCVl/HtwuwIaXbgBUrBkrsGAapnD9Fqy7mZe0PdxagLT57bT3Q7K29EkTDaClenu
L3UgCgbXODdBG1govOMJ/3lpe5aT7PQvFA/2YEkoI7c2OaTUgrujnyR7sAI60HAG
AS2E54ZTec8SjVrf+sqS2L8FcysGz+FOd1q1IZ+kJLYJtokVcBeGbVLmbRMly9UH
SLRymPxEv65WcUl1zeQjc+ihOr7EiG4SRoDBksUeTAoqA/kyHpjjol4xrJC8ER3w
qIYiCULzAZA7R+9CWv33xi9Tll7i8qu1pstR8+lUoNhoUw7AYwKlMkNWJmctT3m2
n/plMjSdN3i6raBYTC06cARxtRoM+3Itm1XjAiEEVKfXbPuZxSOQ45B2eh/SDRBx
P/YSq3UL07+T7VoBbLixbjej5oTD8WN2qGPhjkqXEX0WEkWi5LksptqqDLKcmkPr
S12qsqW1sMkcWU+kCNzQGPKL6bcKqFqerXMQL1MCTvubteCa4FqjB04B5vj8d40T
RsbX2uZq4miLHpgg0zmBgTHhKAVqwb9d2kZd4K3X8DlSB2UOeu0rT4GxsuiKo5Zv
KKCRDFmUhSHQlPsGm1K/MYYrFTqCq9pz/PZxN1vnas/aNawLb2xkzMKwNcAACKoY
Y7P5KLcLqQSTzaYDiGRyqd8qgsgQLHKWHOHMdXV5vMTYCYf/8C97wTugiRe9YBOK
CZZRVyWu3iMVBmbPtxtgJggs+fPrj8xiYCVbNBuyOzr/68MLe118wFancAoYfDia
/r14V9vPg6vR0Ulb3gkaBI6SaedFd3pr1elBJnUEqfQgahdTFP7ej9ue9ysGzrNA
yuESpJna4jLQcIHpVTx9kP4lzK6AVvb/r/G/sx09pV3jnp3lk5Q19ilOCLcMNnHm
uZTcg7qnB6h8fTcVHHknlX64ntSGSRJZ5J+5Qf3FJjtDW0WyrSWtGXn+g/cvK3Xe
xb0wN/tkYqxHKZDFgmgN+4qq2mY0HYi2opS0gRulDnionzYJVP1DvDTCelACL6aX
+oxQSD5zyfe30+KfSeAUMeQarrpoDxQK51qm6YtN5I3ivEUp3KKTdQY9rB0DU4is
cUTCzrd/FVcu3WFSUhBcuBCQoAAOk5bpKB9O5V/qw/nbc4wh86QuNM5puQhCNudc
MLAttB1Hr0ms+DkOF40qJEBu4wMEnghKPxAtucwukGHHoJMNxJ5bd63MZmIkz1uu
rr/ML5wrvmitp51cWY8toynVV2H7iNtrW25AeX8eoawa8u85vyIpOe3ifGozbjnK
XJkn1m4y+jFz1VcQEp9to1Bapt4ziT/XC6bImd5Xcf8sp/LMv7OhZLobZppG/8ya
Ox8FHEEhbkt2939BjYubJEqzBqbsYjHfWakMoG6xqxHFM60yZUOGUwrrNwlXyaZy
Qg93NQOWL4kv7SQizZ4H/9BQzdueGDGBSYYlz0amjPqGOQbqFxbn1jDeCXlPIXkq
jtEQOVv3fAiCLdzSbWbCQKMMj2BzTXzyCdei/UXeRJfBdt9XJJ7xVP1i4UQdPBH0
kuEv5GKgcgg9pu1pYYrZH1aK7lTUBLSFxPEGMJNY1VePn9REGj4p+VsY0ionSoxz
+epTw1kpkdqUmDhHc2Zpv3QnerFrYqOXUK7Om3BbOwYX1ykiT5N/Dfk9tLtZzh4K
MF8f6dBXBHGvvj7lGB2vqkxSAwUydF9bNuDXwAzUeVdlo38xa8coldQGzB60Iokn
5O9dKeERVzsYzrW+WiQ3a2imZUwAIcDoKbhg258Qf0p7jNGJUUHX4j22PvFOhyN6
S1Tm3CkCyJ9BTBcWowBRqIk8oT5ypoMk02cZ6fgCWnNadUhyyLSHr6uPIs4kwt0t
7MXx+MCbo6Q2h8i+/XjN1YDv46Q3Ob5mRlQHikLof58ZenBMwbsjVkLozF7a9Hxs
PX3bK3TXX+NyZFFOQG8sBoJSChmtzYW5c83b+nrfbXuw8ublsRlBHrbgRo/nCEA1
MvkLLYvIhVz9Q2LfD5Qo0On4Ux8Os1yP58o3WzpjmV9Nz9ajIJxf5IgQkftODlWE
V6UgFBLE8i19mhUmiNVuoYx1ksxoIbPhzWZm7ngc8jwQKyViU+ztflpwo/hgI/pt
+qdeyWovISZ0ksCZyN0s3FBfLG/YuspJz3Dt+QtjIA8oGlxNeIEl2ln/uLRGRFzY
DQcrKPbPUwUWd1LygQa7xq2DO7WUneE1N3LR5H111v8leZJiOpm/oPqYVzcq9Uye
1HLXCzFDoi1bvVshQXxBc7mctYoILvO5CIiO3lbeM8IlF4orAqdHvUPbelab39Yn
cOe0hmHY8O3hCqm8XXpKRDeL/EWLm1qEqH6qmiJRtDNzy1drTOFSdIyew7iRcFyc
qK7AEG88fsoC3PefDQjqha6b2m331ylBxZkePgp4AkUvG/QLSNncSGmCYfikP5lw
Zfk57qK4f3frR7DMxSn3bgyWt1dDgU/ATsiFJrh3k/CTJb9oFb+Ywc5g4aysyM22
/gI4oNwALNnzmGwiq4o4J7K04pv5XoJXtdobUkQYKubV9QX29OCQUZvvcQTdqF2H
1ypbw2d5Dl+EheWmYG2cz6wwQwh4wiUVmeQ1pTKdSY47FEjqL3FyCDZtBZcbfPeA
P5ALzR+2/Ldt/qiq0mTneJCXPOrtuov2J7dDH4fzu9G+/0dKOpF21rJvhqzwGNjX
hDhtbVtlPUKwyDCpHArxEk8c/hKnVNyFCmeaxVSJM9QXH1xCDOaBRhD/SW4Pulf2
ze2Zk4ahf1nYzIUsJ9lG3s7wLopGHTi2A1H52iDzmdxcx14wWKAWa7n20FY9Huqu
9H6QTv/n/VQxOEY0TQctuKGJ3d26W/qzqJanGT0xExf8AumHZdKtnUJjRHKBidjj
pvsxw4lK0QrkmGaVy3WHoHhmvQbhgLQELCin63IqY7o77HMVP6F2DF8Vlo/erPXe
XuKI2pCZwOfatXydz42hhxTn8P2E/+nKjCU/utSmshuJoPWKmq5JIF0MJtEKKVKl
SlrZiWn/4nYUIkiMn9lUYAHq6B2SApqC4F4uLJ7rcAkxijFY2K430DXpbwIT+cnw
AIcRXppZmWrrNR7B/hB2cKiMSJgDB4t4bCJtfgivCnnCeGx2jxsLfjXR7oO9E8YU
8qKpMhaAUWtucgIU8h1S1dSSJmdlufjoNks3VD43FpYb9FuvXZq+vn7KnKWjqQS/
NsQP2UtUW657Ty4gZsOB8i0Hz17ENPJhn4DKjNaXe9iUhPHhgG2q16i5/UaulMQt
iDXpfoVwBaIyo+VyhlCKlcEX+FIOAwkIWgsGurTKj5V9ugK2xq1Z6gUmBtafOXIi
rmsqxpXIpB7uMV/wUvJzpwPrJTLjSSs+xoR+5zXsyZCYvC5oarYjdewi+wM8hPu8
Vys/2eHjVVV4T6S8UlxKbGanpCVpdCzvD/sk4jOe0T/13d9FTSVd97P31LOPLwtX
u/kjAMlhCUKnlZFlh5LdluKiy9WUgBFHrC/jKzvSjcgyPNWJXTSRtvjsG7lI8USB
3qW1dSUtFIxqlhPzvdGOwdC65SqHafm60uPcZLTZbyE9hlk/W4hMRJmk727hkOBc
//h9DxRG3WIJZ0WV2r3xoZkdfy4N0/U2+s2Q7h/LE6B3/kR+0vzuExchOW2e9Y6r
dhxPQkHH2jzSZJHZTmdHIzzfW4ZOKWGqsq3kFOMT6wjSU5uYi1+4kK0r2DIEkyTz
ODFLfDe36fKmNaIjhw3aSvfJm2OtI3cYGQfMxWaVhbgKlAValhuDR62irML0ORt6
tou5r2lQ8zhjzlyqfZFI3FvTVjPFZ/NAxe7o+nr5EZnW0W4NxyiANBCHF+Pp4C57
mAMKufr8zCjA6ZbjKhukkQ5HiWYZyZo+uxT11FlqdVHjLaqbgjtF8gKOk31+NogE
bwWlLw8fkDJy2C8+ZzxE5KZ7qiLKmaoS8Bjf9xnz0m3PL7R6JeTEB2W7CabfCU8l
xqnNhuId4aBOHdk89sJzhcCbdPFZtFxboZlcY2s4N2LjFruBSXOOPm1MVD+mEu3O
w6z9RUmqlDjEN5EpwTZaspaLpbxAVcOg8uSdW0a0hkw22Q9SO8LkQ8BeK+qsYQz6
m7/V8G+hkLqsXvngNrGUSVAv1dF4B0qIw0EWJ1OvIgzrWiT2ZpceQlhu77HW0SgG
jFrl6eR/F78G8+fTn4X6HRYvVq8TF9zlLEJmWuEhYw9lx6GHPtWEdUGdHvN7kTRi
U4SNMbZFaVKvTKLtGHCfMULBDUJNsE/WekJiOzcphtL2PSjBPdBmdV3MBIX0n5Wg
gsVRAeUscTaE7+yB7EmzDHPc9bg8ru/IGyxCRgDL2S9+WxyRtep+zkCivFXspzRB
fk1u3gN9TbmfqfUwD1c67fwphjbEDbNHRysJ2p2BjK2+7XwH+7poYfoVhdYSPJ0o
w5nRSQyfLP1KkIvbFD+mz9aOQHv7HpCmNfe67IeDwl3EoGzIFoFbCZfUYIToB4jK
GnZD/uH3SWZZkvrkqM7EWNAjnjYTlAiVOygcWutU2yfTfNwiGvfMxp0exZwZF1ta
Xow82owZFNEBjrsvMEd+1ZselVfrNPyoMSKIgXw8Cn2JKtyepF2pAtHJZfP7JzeY
RJcd3KQ3HgEMfLgaRw5SU1H6q+ZyIkMe2Py3OEA+Dv4TggT0D26YjLSp9aO96pTy
Dwww2/jWqmRdreyqif257hyYkYaMEfxFjZVIu0TDJesdm2TWAN5PiJu6Ipn9s41Q
FQwyfCiCTVdqc5oyRMrPYWojovQtBM8uUdWGyzCpjQ/odRc8By43yhb//Ki8nS1j
zdqSKHxhVjCzxNxqtRPTMIPxP527yreZiJW2UwlDVXtgpOHi6QufLlg7bQfouhov
uQgqntJH1KKhEe5QoPm5SLRKjQLQd73mpUXJ6lCDLoPisKZMR4lavBKZ7m5mARhs
nqHatfoOWvivZ7mZZVLuUrLW9U8RFtImZMXSsTo8TnreqMrINAkLrrjfB070zVqF
eapq4p9ULLepoQALu1FE08ynKYPtOz4WTGDBkbE55dtEuqPVvU23malLgz35gnW5
KFszS2YHrJaZQS8GBbwFraVmld0+Bw+q7OrDB5niQ5GU2tExj5t5yYt8kB3oIFn0
s8jfNop2wUcA38u5L3YzNPPg1TTCHB0FpDNNo476KeD9QDo8FCZCgOyiNiS5wKQP
wIjS7X7im8q2t68g/o9mOrB/Bd0OZ3SaEXybGKRY/M8d3dSeLKecawwcWM67O+72
a7vVVaW3QR/O0yPc7azNQt7mYtOX6V2UDtygFmxmzJXgEc9yL1VQrrFnLQSYIDwb
1xnWVsl3wP7S67ewNNtmCky1lvCIclJ+d0tBAqgj0gfFFd5JHOdo/uAZJbCBJ9+g
YxJkBUlPuOePT+muiOsncfOqwy5aM5Ed3QNHZR2Woq4yudn2CyDUbfASu0rSO4Vq
lK8DpDb4Oy1ab0OvupheWODxgmzJZr840OQ7poh3+xhLwC12PZ06QRMyuoTrShn9
QaAPrsY8uCPOBuIW4CIpVqIAU4+GdiIuACYLp97KcwJ9AfgvinvCZAEOTAjg6D40
EOjHw3GX8fDFpEIwYBAdaFOC+HYNn0vupRfjSWw1qVpwN2mETBmRh6JmCaWQ2YwR
Vp0AAZ8m23BVFzlnckdzk7e14YXQLlJhqq7w8HYWSWZG46d2QWI+qlKAwYuewfaC
b2jUG34QDMvsfoj20OCzvDyT8WkrdoaDPZDdoXRCIuB6S4R6Q6c17KIOLKev8E0B
lIW9hmEaG3bAhs80ZPKF71BkUQtq79FgUvkzXBVyjazyKI4bUHWn0AqFBA9+L06+
B8YW/bqE654TQR2kKyXaONCr66qQqwEZ7EU/1FTU3mhB5YcJb/rlRV3YOJubNPie
GGdrnQWLJK+KJgTFncWobSPMXls17GsUu97MqMhFfL8FbILMuZ+H23DO9697Scgk
ChfqbBhHU8fUJB7W0x+wHbxfCeJC6Itwc5hnfInpnQVDfD/3O5rTZ5CuCfsDT5qd
azxju7yXl9rYkKuUx4eK7hOR4/bVw84V7DkXTbVybD/wXt13Yj41kJe3juq3dpcH
MhKgAlx37qHmDJXTupCEXlAerDk4Xzh1Rl0jcHDaSLKLR1oBok7X/SCTmKQeEYsJ
fg5fpLwp1VjyonMB1Y5YZyplArTAe358dIb9MxcbkQ6eDvyBoFD2yIEvt1aGv/x2
7urccElt6veeEh1ADhVJMpwlXnEiZdHG/9sBOk/0PtEci/M59ysqdnvliXJEPs/I
ZkiOiueNE9cDhIx/0f9ftpudBKQG9r0ua6vbukN4tfXmdU5tz40sctTGQqh6vrN8
i+mmD3ZYLl/FxvMGa/GJWH6lFTG3DXQAK7fsUTUx2KRKlqNSFQGfkC2wv2zsbkHZ
HnOFNXDywZgcHI6s++DA458NrRwI0pE3zAG3QBNhugXKcoNBMEXi8cg8Mrh10FMA
KPf4i5h9XzJsnS//C12SAtm3I8MdhM+gwZhJhXVTSwYo/WX06oZBIlNnPVlsoCE9
PfWJdI4CT1HGtchb78yeC7byMJKpEVqR/q72e1e8Dgfu9LsWq3WSMPTM4GRfGUZS
VcReErJOkPY9SrkcI+gn6OZ7Hg5JhAmDROoAkx06Q2+oeetUU3PxqfU52MYwFLvf
p5CITnuyNBlCN6Pj8szvLikIzDXPeliK8WHq1LusvnziEGpapHuWdB0o/0m5NVVr
EhJDgksYmizQhsz9dflt5Zst5Qf+Ngq+bGyPmidSy/KLJT/WbDMKiFUF3369QWGl
nv4TugwHY8PVPjBSKBGRGlMFaXi5YtGrSfE/7K9Ck9YjCmBUvOOoM3SPi11yW6Ic
4jjEIvIh4skPZoEZGOeu2hN+rk8QnwNtzoneZhXYowaYlzjAAF3I0GMiHdXM4n7R
OOfN3icRKrJqq0ttNiBrryVIitRLPxzzyYsXY9c/Kex0c8/GRP0frbqvo4rFDtNO
zy+UpjrbEgwvKraXufiFP5LPovdjx300YY94mhOsOGkMAWXQkR2DQ0c6nVHItZ0b
67CBoItS47gnmC41EnXSOjyjUwfLnkMzEh19aMyKMSZhK1g7N+DQQnoHosW8Ft5O
NqwH8dwapHl/t1tKuwpEC/gZypfdPsCSZGLQe8vH4gTM+QNPyYQQNqt8bkATwtDM
2Xd1jlgpfX0EcQe3Q4F0Nny5BtrApd6B4Du909Iuvyy2wDNwxLxDIioTOvfA0U+C
UMbJcuPX+xrTYKwNI9ixXS/V85iloqjWlu3pX9gSdY4R1W6H8jWBhZiH7pJxY10t
qi/rmfQSli1uSayLmWWXGpzISkkz7KNgr96J7ROiCu8u0EQv4Xsck+FxdjtRS07G
zqRKxOj13bEU5ZBqMShrQRQ8uWD2QSeVLde9pX6Cuxl2oJL3u9sMyihMI/uhCiA6
j84EG55eDW6vj3ujGNeOTFIlhVIRLLgrNrAh9cLEKY0iQdoc4JkHB8I53Gev98XO
gWs6kyJO0NTW96eZKOSTyeSYJTEFuQsYuynZqLiZqdRQWFDUTGlXTxQS0/TlrEDV
zHUAeUHwsDLLo1YfAYvBCIc2V5GSA3m9+s7O7CGoT6roNfIZNd7Qw+DgoTw8YJmz
NUav24eSfplaIA9hOxw4F76bhJ0aA2yyNwJGgtcBeG7swtY1muVGg6t2LtQCzKd2
jprkj8t28Ce5A7ZAMpFKROYfRruk9nlpwsNUQbVkvafe9OD/01HPDqA6fcFrZT/H
YhG0jSm4l2RASZAi+Bp/sDKd0ySmDwCFlie4PMsU9H6rrsIa/M01KcYmIcm2tLFt
bUlCDSEzIrJA9idtkrsdHe7W6y7FyXF32n/ViL3Xyp7fB/IpwGKX0ozvqOlQSaRK
izq8yLQOqH6O4Lm466380kPqyHAoLGG/Hn3qemlwiLyiernPmqoYVdIAcvquLBIH
ewOsQwDBAASKpz4p5mL5BB1JR4r+d17jK5ulPGoEj6z8NMIIbpG+zgNkks4vtCS/
IAeLV7Boqq1pRwarjCCdaHkmeuL20Pa09gtuBzBN38p5JjEM5hnOgBY9i25Ws/z/
swi/a3VUyt3xNuuGrgfo5bq/MgV+0bSgHrRBtY8P5YH/mjlEWuoXkZaR6S4aoTU9
mbbFanvotWrOZQYslN9RubPT55NpaJaJEt1+FjXRyr10IClT7Ke9kUMSt3ZoKrTv
t0hrriOJw6h/Ob5+suJhA9N/uERPZf+K7+0pwN8E8VJkZSc6uyRMCXmnfrBwBBYj
VwMdPeBVwLEjhI5bLd9pXfs38lMFCSWe3qSYG2AycRHgtnueLVyG8WamsKTWRHQv
N1Slnd66kLcPS1XEey/wTpix5SR3+Jrq/DeiY0ADjL+RmUt0CUQ0XqG2e9EEh9GY
ffTEIwNwYdwv0DMMFcd8wpBgM+Olr0C61EqZlQvP4T+xeBx+zaRmcc13PNteVCeu
/CuXUsb5eECtluKqsW4brWhDqmc6H4Y1/IGyYOVQyiksqU3Cv4wPdjfTiKf0JeBv
xq0NLZlk7dnvDLFzYY5ilVqKDASeQ5CZ+roR6vSU5sim6qKUf4+HEQIDGg8kVsjY
ciAoGzHNiBA6/fxcvFHSL+kE+iytfEKTw3EJGM8KMbVcU8L5Z/hmCQRdF2HG4DKr
5vhajuFmUgor6es8Z+4En3DGSiYeVQi0+VV1qAtsV+5cIrBlOwAz+Vy40lQEDdcu
sHfrrA1BNcOuaVPLQd9SXfQ8bKE0sMNDoPi8tXqQyx4By/4VT3bSenrwoonuuwTe
AzrrgCMp3Ko9bk711CaQmuLgW/Y6dPO2J1l1Hc3kGwBbvHjAHWSKxWs1fHDfA4/V
dYJWhslzxkA0lhgNBbLf83pDdeN47aXTl2q7rjKEqYYWxtLTcXJzDuLEwIofDCyW
FHuhgfBs1tQvZBcFLIXKEVgV6ZcZ5fyRn65Je0tdM9E96uOy1nIkWdYtAJhrkbWS
49t02JU1+hv9hQmuri7FMGbnxZfPB5bVoCGjoa5kmZP1ylBi4sX3uK1+rB8BR7eD
4X+mwXPZPm4tX+esoqzvlKd8VJmbLBRGRcFdJHRnnwVdFUxUte+zK1dsdkttKEVb
/T27aCQnmSEjNrQXLNivUJCwu4q/y4yyJObfuX1IgtSstgN4rDr5zjb1okWSUpBv
oAO19RCZfSePaK0wN+PdC8F9sFXiQZDr6qFq9UDPILD/qTgTi09hQBjRKLxS4fQT
Ek7LcNQAi/TrUYNSQR0VSMNMio6uNELhCY1+Xl1Bw1i1xwh7Jt1bWFZS9IYhgoDv
kZu23QqVePlOBdU282omv7WgFQkYNLQiCGKbYZgND2kQw6y2hy8R/qiezMUTosOg
7tM1YJTqZkYYuhg5dcYUmN4UnRYdo73VSX91QBV2u5c/YBvc7SkeJoKhSUxJxZFh
rmVJZn+K1JqHotEjG0hm+zEzxw5X60JV1l1kCNoJtSyGIoL4Fbf2516CdGQCK+SR
MwJBnB3w6z+qKnjVJSnWhOqIcTPpufFetxnbzkU1FeL21OBqQ+DZwrkTKwJ6Ic5x
Nhx10mKvVWAwWvsaNfOEfA9JgjuNeZ94X7+Ap8YhYMEWPmoAHRiFbx0Kbt8UUtCU
jnXkHN+6qfqPbPfi8XPe1hfCjMcozAkHEELnQUCHpTkLgdY8nXoj1ZoTErl3zVqm
irJ7BF+dwUooH/dPEuQS3DlhFYm8am0BX9uMjBwIGAc6EyEd5msbF9D1ogcMmJs/
IRtKZZmC3ZcobucqW/sIPZmVNk07Mbz077sEQxf54ik7qB/76eT6rT+iPVE9YrDm
BLgSsnKFRjvx6Z99QJ3W5QxvK0WK6Xt2q9EFpmyvOqX3mhTnrK7km7eQU0BcJb6C
7bp0BsghvyyTITB4sx7NJCaWYAS4DGjncdZB+YR0UB5nkePP8YrriATOkWBHP1Jn
9ix7pDKUOVvC7uDHJqI5FOjGOFrEeCW6IJNXxfHnwObNMhxS1KYaAf4skRvL1f8Y
Ysti6lbhZ+YawMJ4K5OU4MTHS4pJwYsd4zXbk6yex4+4VDszPpP+RLR+ubYJNyXx
vV+ekH4+Y/N1QP3I9brq3BlQBIotrwkyRebQ/P+PzbcO6l9gbiKwOEb2oe7fv207
gzaOYklb4L7d08UCOWwHvakjNPHmCQPRmkqA+8VSi8n0FmixNIjddFlmOToJY8H0
4k/rTZxTzx5pAXMkKlOUlOSJgMEI8X0e1xf1aHAJ1U17UWJX4TLZXhYhKNF2UxbG
jve/WkkHuk+5k3U9uycl4czLFJKHAhT+XM2/LmonRfL2YJQW3bKvwF7s5BQL7cM+
hB5D+kfcMGQcJaRTJ7if/b8PcIX2geYWgejHWE/uxVKs1Cy0f7edr/e2aTw/WVx1
k0D1d0pedZCFCXNtNVzAT9NftBhRhBfIOaGTudXwDwzttIN1BZafaZldM7ORQG6K
jviNW4Qt0Ei8TXGUGpwMed48UFqJnrMgopCCJNbrl9wmn3Dh0LpHnMb+S0qFj7Hg
v8KZExIoKN7DAOfViKeWygU8iVnfF5X54SVrEOu0odKDDJlLE+ULlT0El5C55ljH
mk20TgPeN5rDzt7gHvCL5KlUTTk8A1ZSkq6MKI4TjIxW2kkyjV0etPwyeUSPrTOx
8x6KHH/a4i8bgrjWCj067DcLFmT2mHDbLG0N0Xu8tHxLBpJRJzFPXwOw7pEveF8d
xhPoMNKhjTtht9zVbjWG5gqWLjBvN0NjJKoPUsW3Uj0NtnLtaziwl93UGY/nKa5s
5TT7xZuzkSas94JRf3T1ni84feo1yImuGTYuB3cXXVGEoz19rNsiEvVdsTXLviyQ
xHucVQWam3x5jV/19NjWO3mWJz0DS5Iw07YT387NxZQJP/B5K6H5c5lriHHIFnrC
crqtsNm0ytb7Dmymk3cWFMP8nNKVTOe0Kr/YHTI1q/McCGNypiAGrZbDjX+8GU69
lfUL1tn0oLWLsdqUiSGxPqPmi0N3W5v06e481wcMVivENEtaQCtasekgav8YfBHQ
RohHFyFyPZIbsc8TAWPGs4CklXQBeYOz69geRjb0YMKnZrqYnZQy5SgLU3nONgv9
LWJhydtUqYqRcMwrg/X4ef70duXYcAwAAfCh2n1XgYcnXABNN4QH267v12YbvxAs
WzyjaXPRi9YcYX+rNOjJxYEPsHLe/APzGBVXIYYmChGk/zcnQ8m5Hx8/TQ8WCOZN
kEnlm0u+HHwcgDnMib8hv8tAHxPVz8lJ8cUlwp8pgx+ns/knjUu0JleY7XYDm+XD
OClCUJJK94u1KR9a3v8rLr4ScxKwWTrN1kSLj2v4Jtf7+6V4WWhUbZdHw6dj8tgN
73GqKmKBlGO+smexKLa7n7mvrjcjE19Xgcj9l/UIk2v3CY3IcnQkIo2qjC+O+5Wi
iPZJWld+clFpGJDwdJ1EfSPkbyh1NdDUs7utNGTPNfzO8fpZPuMkD0xPU94ly+zu
xGEsCKw6ylY5pT57eXV3M5tSnOXIUpM1ClephrTevOW2oLBYtY6T3nUSMH20U7pl
wPSF5kHYhceh44alX6IN4kPT3DQliPpVe84nZvYjAmppeMlxa0uFP0FKHB0HPh7p
uYFgUKfwk6vIrCTwqzLrXEPL2BIEUPEckoK0Z7mS9WaiEC0fUnBARczzW88SI9Pj
czQwf/ujYn+OoUyJVWGKmFFz1jPllb4NHQArHZSOMu5B2BtDh55azRKlCwlBKlnn
a8VXB/0wGmIsVenvOcSxB71jGpcXbsq9Ee03QzmpHXP5jz56tNJJNP7MUlkHiWaA
brsRfQoNAaEdcQzL7Jkrr5qjKjp68x9g6mpui65xE5BpWBugj7D28j7jBwoeCAV1
XbdkzbprdOtGkUkBPvgqYcMEEN7D4cuwFvvoeLaJ9UwsggWKV7HPogB2nvLK87mN
8YJAosuQl1Q0eOFvL6RyKHrwwPjjKo7nXnZneSB2M4H2WZH/7uppw+iGIyDdO4sL
fUoY3Y+k9qEKMwSLfal9jouzSpD95om+qGJ+FCqEELCrYYL4Jjxvig26qzcsDi7o
WclY4idwxfL7foyQo92mEndy/2+ex/PkU1mGlJMtv8uMl1kWblIYxls81tSWtXhU
suf95jijUrDtxtSZdfmfIpmCt7jziaqQUFzOVRarN3zyxd3BJdcE+dr2W11rxupa
wJ5SZGE/KpybbcmGnGAK6oIDCXdYfnePjXLlRMwKa4cHlh0vG4lwZWcMsjuyCXS/
+rd7+FOcE6WNqQNHxdTQVEFoz9qf3Z4H66BrkPM6DZRZRFlRybssJqO3BQjn/kXw
FNFAUNYGdiT5l4MoP4P88YS1/+0Oa0Kb6z1D7Y4bXElH7PZepC52XCmjqZSzOQQt
E4xrLvmKr7J5EVmeYbUfims8UvXY712w9srDmaBz4BHTAEyzluIbNiTpylv2bGQ9
M0AAGhTvPlS9XCOja8bIZR1PvAcgE/i+z6lAFKN2CJuyDmSWDYfNsWBIh7h8oaXC
wETGqSp7C95s26TdxsipMnSzaQdNnWvua5romwQURyZFqb3bTfQrgdUdiFj/VQMx
5H+kGewe/GAkT7Ry85r01kTdupp97gLzFFyfYvUMsKXVeQFkWDaXSNEg9B+Yu/mG
/98KJassQNrfD+WJ9FJIk7FcsnNEfZ/3XuChGNdH+ntGbub+9z1p+jZN+6ftJWV1
yt87MUsO5h3xTp/0tlDxBIIR0TrfoYnl4e6Ai8tXMpby63pzRp/RooldiHGaQVzs
O/qb6PfmlE30o417hUIz8NEpwVNfddwFb0RCTxT3erbpsGIMRylH6lRA6Cz68l7+
uzfmLfzfGco74oxKFpai6IdWmW/lhRaAIquMOic3qP+mdFPF6HWVXqlvlsHp95uf
yzVV7RKVhaezioXluHikxWCK5RNaAagN3+lupuHZqhvWU0bajkD4KBFZS/AysxCZ
Rubih5jYri6WAZj9CChLgAUKF9Uh55Jm5u85B+49UcSN9Vk2QU3A58nqfneG7ZsE
jJcIIXrHoSgVcnCHV1D+A6vxOHccaKzhpoZ7sEeCBAM1FZmf9OiusCQBuBpzhPWT
dFDHxutyDZVQL2/xu7na5GpEWXFfwvXjGdb7oWrHN+XG1t+PQlrPC26lFFRtgFY+
JORPN+7O0mHeP+b5NUOMwJunwHtf54eQQ5cCKkT4s1839atPA3RqpSZzMh9p68yY
oS46fP6O+8FGtE1LJDLgMnAbNrt+7lMKxbxSoz2poPcKH6x01wqTCb7YV1s1S2ZF
U4RHftJ8BWSIMLVwijv1sM+VQLoWVO4O3hTZ0/+M4Md5zwxjoB1AGvuJxdpMf7XV
QWr79WAWtuOkXCPEI7n6Ht3geAbughKpIxFYlf99L2SZBp/meMqEulWih/DJv/ca
nOMin17u2WVSHnWU+xhLzzzvLVD95q+wkXZA4NhyEQGMM3WfS57p5RzPIIB6j8qo
+m8oE0sPmiVvrhMBaK0pvDKuStWCVOuep+Nu5kLcE0wKj0iJhDLCTOAHdJ/pzMeK
Y1TJTkvXcxZ1UvRmr9ATDUbMOSU9fThSWSG+t639m+Xr39eW0svpqR59JApudzbh
L7zSuh7w0ER6eiNjbXhRYwkuWgKfTU62PywBWt2MJEysTHoEJdHCtevQJHaCj2zg
fudqh0Ynuy/tz8bxsrQzssmcx0OxgDyNAzA4IhY//5SjLoqBbhqW9NsTDuAQ35Xv
NcScYnBHKVO/r3hpqsQF2U6I+NQbp1ZHLW0mBKk8XHOKRKQWrU3XodOIJAcv33Ff
Jo1bEUify6YB9c28IadF1cE1lh4v2M/jERCSI+XpPufbZp6BgMw29L22LCdyMCc1
UCXIlh9QBjb5mHwkLCfG9HI7Bhv1Z9c3LQ7Q9THDAjFexdeXb/wAW4U30P0MGVW3
EMm9UB/fZZBBgxEsby9hQzC8z8CTfnFYHnptFSpsbWvy0UskNguhJoepEwF0XUKA
ppCYqkdY4y98PkKJbqX7EP9Y7qDL4pnUPtR06GsASlrygSQzoIjNKsBtyJu9J6eu
lBUXuK7lkhNKl9eYU3eS3V2sh0iB413HW7htm9mZmC6q4zwesmWfueJkv2kJ45nN
70NWuGFyXXDZSn26y5IpUdShI0++u/zvezffQP7ChXgfGlM25vEAZHUUSqIDv84M
PXi0xYtgDEOLHbE+dPin0XolcnGMhlvd/mS3QXeSWdel1cpnpfpWztx3hPfqkgUK
vQ9lLbT9zRTS5shF+ktPwoiZ8QpXjLSYU9NDW4XQBj8D30Ic/iOmpAkAEOazvnuI
lQlEMBCwfEKF5VFYnEus9hC/mHP06YRNWOXjGyGm7dLYXQpyW7G6PGFYMtLlZYcU
gkELKWGdBI1SGTn/4v5TadZoOHNdQiIrPBFKJuaaKzdJdbp+Yam1JbykYyuzYYPu
zs99/GBlqY8MNtuDLy/G0mQtP7lngzQNtpvGurODVKiyKHx9gnHDz59Rw8ALARFV
/W65mTNmKSTLdGfahVdIHFry4J9wms2PmL1FxqyEUNrIH39JkzEOVSzwUwsq12p5
mE9EDs4ww/I+pYagcnVFbUtcukIk+wQeY0osoON7Ze+wDapbKaSbNXwvvVhHfxYv
mpvfGt64PdBpEtTuHK4LYAA1dYHy1GV2a0aBXtt6xRqF6JD05BCZW1fy7Kn9TgXB
LiBACGHuNhPVU7Zx5kqTqCzZGrBKwvhZjAYA0b/H5aQyqJzBNMp9zkuQ0h9yRvwo
1wp05LOO6LTwu9z6o8Hwoy/Cb9UwKZtDqMzSu5wlsIXODR1pf/+JfHZ97Ifw+Hyz
V0s9eQC3WwTRdbZaNWh7RIG5O1A7sbwAmcKj8TFKpIysSczVfIsOCyD0wXkLfN1l
y1hCSyxHeawhgI+YulcWbz9v0/a/QN+n/DaM1ya+B2iKtbNk4mDX0eVr/ZUuz/B8
HtmOmQhV5Y7JpHD+e1vXfWVlzOckLChtkrtgF5OABNun3z8fj0DUSHXXpk4A5UnS
M1gsjwWH1fiK2M8Kuep4Oj4NMp+WU4StnKSbTssfgtQRaAZ9skmwIISR1q3hr6/O
MT4PU6HwBChmuH9hxM745f0Ye6vXgMqNypLoXyBOuaZA037B8BYSQfl/3yquqEc/
MwAnl1nkBo7X+zFaVdhh6YnIWF+d8e7oF2dM9+edCdlECB8suSamYKpiLQ9hC5YZ
7wrBNm6qqNQhmhC9ygiCkWrDU1GK6x8Ez0G4GIl8hpefF0xKaUEZWUWz5BANkruE
on4Sd13GIgMHXB6oEMWMak+R4uOv7jo+P8MnraVw/IUw6d1U5hvxMgmOm8i74nE+
e2H+45tSaXQksePr9aWAUaWSubGJpnvZFnVAd/WpxlVLw5s2sG4LDCFXbOwpqZhJ
rywD1ru8gSqiUIScmXeKjpk2hQau4nt02eZGwxsVtep2Sf4Ii+Hl/jhcVl9ZAfgc
j/v+v1ksIas8Tx0TCdt65v8O+84sRboZ1OU1z6KW5d3jJG+J3iQ2kF13x/kmGi9g
xWSLAD9TXPx+9AnawnHH98Ok1czoG9abSxwJhXBIbAXjxvnuPnDRkhS+oaxROpp0
CDYkjhQA+q0OKhWAwHX7yV4wOroP1nTWKHujz0eF13SI56qsZ18oS6xBvhkpZsWP
hn6hNo9UjoulQyjg+W1unXndclFgzEEc+Yg62jaOVlOclTrkKAnVeodkY5wQX4rx
5TkFxT+xBzFKcGC3HpRNSlxFwYf+f2EwDBVui+aJ2yiGWcSBcL9gjNyf/ikqBOxD
TQMci52ISFRZ3M5evgpt261bSiaxdquZ6yKYS/HrwNGCv8b+Ku3U6k6x7kOq7fjV
9IMm9QgK/bwoBDYR8Rp/MfwIncOiugcYv0CqPCgbXc9d+pIk+/24NPEN6NvCBum/
VIb56iZ0od+Bl3WTndQxFfTaWJDx0ED9LsLJLACsft7kR6rNUPoaHlrMqITvB9Lz
82oUjWSiAxozF0HzPwS3f9DwfSh/oS9jbnuIowtNnMQYYj/VjhoL098LzFnNHWQA
2FYJYlVIN+rdu+OJiwjjMm8a8IQHVE9wDoTCS/eR3TDxdMA2Es/Q6ZmbvnfXQuZs
Zesh+WYgua/evinkWn08jkGQAF9nA/VIYFQpQBUcQbdohQOjSuorbHRKd1U40a+/
xY9C5eAO5Bg+XOGRB3d09zPVMwGBMmvsdX1j3gDuOGfvRWVe7tRET98GExINR1Bv
JOp2d3rmxt83SxqPIBfMbPyZMJd82xEiEEIhUaqIwDznyvChMzs777Szhu2Vn7d4
8ZAWYC/8wyP7rZZ219qEZmyBW1+f36MQaqQthRZ8qK/YIbLZ+Vk9358VBNGAYxza
i0/Metu7efPuwzPiMZzH0UmWc5zbw0yyOm9QzkF1j+ZdfA06nj1rEt8gZzeZ1cX9
4pu5qX7qFPo7K6OcGZXViHl1yduRgnWB7G0+Gxc53hSbG9OS2ZFn4fhax8zyu2Tj
Mz7V8/upQOElF0T6oODokSp/ZQXGqcKUFwMDGs8v/QcL4ZNhpn4WxBZCgNPGpm3H
J/ASiX7cF22EHnq5OjN1hx0bF7qPN/5/rD0RI1a897JcFtVo8tttlrVS9+0V7M1j
s3ZKVzNJXtBtFUtPsUx9uBemkWfDyJ++dhiQ4ZrSWCb+hFyZzgbnJiD2mlHoEt81
LWJGM452z7XzxLcdByXrDiuAppOsIMHAy0m5FBW9LvdxRVN8GRRNroNQt8Ne8WMf
MIIxOPQtlfJP+J5aOb0wQQpKPPAiSuunECqx1b9OWomW2mAqXN9rF9XF3cjI0Pjj
dlPc4NXSIpiQ5fsLjkrRF0CBFX6qJsQrQCpW1QfyDX08SWU0rQBhnmU4QlYvJkV/
DJIX3i9R9N7gsMS+qPfI2mI4W9ohpl1yErLF4lt9PJw/uszUVvfMQ8Bdb3XI3/Z/
sq+8s44xX/DpS2oLpbv8AJr08mkrKIkO2FO0K0HNvQE4AzN7IMgs8RfOSJIa2RDT
i1Vy1IN5v8xssgNOiFySDLUCcqXDYyavEvmGPUgBsMWUJsckzJdaulIOTy/Xtl+2
IVsNoRRNDl0Mhf1uG/XVdLiCsgqcr+Ka2gloB20DKglSa4A3C/YCc5Or2fpdBFKr
K2Dw/aBoxNP5rqajJaATexGtLLZkdMjsQWYx3pSxT0R7HQKdxSM5HBldxehAbHGB
cq6Xfrb8GFZWyr12vpJbvmmwfbXzV/tVKK/V07bUSZfdzhMHDS9gS2dtr2nz0yVZ
Kc0NJRnQUrCsRSW+DvHiHPTSVW7hC5oeFwgSa9dqL2y3wXlY2OBdOyaUpyhRM+gT
jhDA6SzZF6zX04KeI+WuaI0dZZSvBdXhyQbgcHgtcyUEcXtbDsQ+udHq5GcSrJlB
irv+WI1fii54CmQkVfk3BxuNemTd3JNyTX5Qd9i2GhCrxCFX9oXnNbTiGqPvsh82
I8VlLh+nUGIdevBuRvfLHQX7kB058gJGpmSiTtdOLghwFqxNHD57cbdcm8LeoJWz
eHRPTsvMdDQNRYGe8QeMUufKKjd944zikh3Ijltbel8STv6qTbTcaqBDZpDeWBVA
sGI7sLcnwnH9tzlIBG6vhSPdz16bW7iH6U2nR/nTbOdREdkFvM0Ef2Vq8wljpuk7
hVsiWZIc3OriWx5ROw0+Uq6GHiRid+LMsIx73BGOOuYZGDOGtslWHjNoKFdNUzJt
BCMFzp4gPaReMiH0k3IIY/SfXoBRcDWiwYQOgcBqd0ZD3DVsSxC3WDo8GGJ9ZFsu
ZETMVOYYGEXt6gIVonNxiRqYIA/iUO3J40zvrVpna75TBdpf92mmh93QxILtAfet
s45hlAhCoZd687noDF4A/HnZgkFsCU66UrW4E1NGesMpu9jcLIXMa4/sz5jkmuUd
io2t86p+mIa8FYYPZgStbRUvq95wknQolF7JNBnBcwq0P6pBVLMBGrxCqPLzt302
2xUofEK1h3GEhx3D6Sm/F7vo4sjtGF/a4H9rTBr4U5o12N+RvzRy7Ko+XcCHL6Fh
EGGWQux7V/XhEpjxAOsgGoVpOeXDq7p6KqG13AbTNhDeOXgPmz3Xmp258cQZqDQZ
onz8JpGBT/7T/S/exKxKbfeM6z7a2P0rD6PD82T3LMQNbBKZKzkyYy1M8YxIvDM+
s5i2s3pLAId+NyF/nT/U+BMsro1adr1QF2gT2sYsHOzJ1dEtU78rbpdkWF/xSQkT
GcUeSw6PUQEBDcR17KpRBf+VV37SanTvWX+gNJ7HNZdALeLwwDWyfDX2SHghna66
xPOotyhe4KxErEcEELt5yPNxQEAvpYLbH4DxexALNvWv0mrvKgUV/0wleR7RVbOo
VzwauK0m7hAW58pTsZeiKnDx+7hUiKCzYD0xfVmfRZhVPsT/LVZhsNNndGia/rGQ
x0Cuu+grrkUGJi03zam9U2NU0evvcj5KJldhm/13T7EqPRbYxx2Z4Tkpl0N14gDv
4Rvv7rvlxwQ0A32S4LKZQYo8U4Y0Hk+Y87qrF7ToEpeRa3kbkixomEHg3quSO5Pq
RHB+6Y0bK2LIrtkZV/B1HBQ7EKb4jfek+aP+b9rKWgiGFJShBV85x6YA1pPcXVUU
IE6yCcCwxOoH3asnMe46WjR4uTGp8pOqCWpSktiHaxjhp118lINmx0OZPRxirIO5
kejY8UIghW3+S93sHqAF1zibWni5VNYggs1Y/nJvLsSrXlOM5hsS4p8AiQFC9CuD
ZtfU6J8ieNQRhVY6m2g13aNfeCGyrRqKWhogrTcbY0P2gbF5pYsYqlpCIOpsSmwF
6K7xn+1HHooD3JQVRs5VehzFRm4cRmcaSzNI4gOx4O/t8PS9YXiYxjWsnQCRfZZ9
3Qv+AfYJqGlgspqAnHeQgSSdcitlFBwBVbynhaqMgxW1r7DvGmAjAPcB4D8IDbsg
lorgRHxv/adlN5SuMsvfUdfem5HnA/0cZ3chivl87m2u1rdlLAOroN+fxySyBwvB
xxcBh9kdQzdruLk7ESpwd3eV1FbUD9CBScdFPsnku4KHecNNEoktqI901dBqZZQU
z4PFCXQJOFZ95AkcsC33wiHOjaGJybNQiH6pplB2ZysGn6yI49eUjZfExsWOlTFe
rcc4CixIPsEW72ND8Ps/+aCop2CQnZL4PtwcrnjpmCp3/d7nIv1WF5mBi1fQbUph
Puw0Jq6KEdZvjrA7Sf7rcgB+pICeSRMFJ32q26TQeXmjV2KzOgGfR2rIxQaExhDI
stSVCTMCnvGWyxAQ9d/Q03PYuex53M2APiTM1yseDPDK9ZrvWRDK73aG81oZzB20
KOVjoG0Ylm8CbxO+C3u6GAvXC/5gGn0Ahfg1owhUlY0C3RztE1cxaZoV8vpBIj5z
ZwcI0RgaSHYfFNklJpm0C3ZxPWT26n0P3y9IvQs4cX9Jag9CHluE4Ui6szn7b0A1
LNyD82anl2JeDflLX2NWBfbpI15n+bgSAUuXx0XRCgInqbTMhxUS+9YGfKzVnsTQ
aBuDLNKpusB2MMtDl4d/cbYtnktJPx0oO2EBtYYDLcEnGmE2aq6eHE4+AGpqp9P1
09yPi1M9+kcCZsWfe8AW5BAewLkgJ3NOG9XhZKB4e70YQXffqyWn0jGrrviZV5Z4
AFaXrT8hjGj3Iqu4MLEVPvHYdEgohZ7CtgmXA0Fed47O6q1bzh75K7dxj24dPAsg
cg26eClA46Z7YTQm/LZbk2WQgKw0HZ2tWnBq+xafn44MX/VRQq1kRzHDTP+gKDI2
X+oShykjXeJwDMRZXtKPG+PPv/Tr46mmltbQZbnbSF2GrPeD+AQIbU5bfPydXMSY
aHTUkpKuQe3ThZ21jpOo4nRQdMnNc48JflpbV5yTByuF3lMxpUuB28YcEkqBxpev
weoVP/one0MGgxemNpxUqBqzPAzjcqUpqC0P+LyPjQZN9KNmYsjF+EB6Y0F+hjpF
ddUZCaz7/5CRzvNf39AfjTOlxArzljYy1sbplf9bIV2dxJVWEZADoElzt+jh3prv
xgL4fzsw+oaceTbhXwEXG0c4Yonzx5+XakoFCwK7mLgQE5hyXS85Zfs7a5k+ouE6
vE58X/3A7DBRQ67EK6S2rsqBJEk6GZE9bNyCeyFFCBpx/K+DjDFg3U44HoY/oyZa
5UtVkHeIzUEgHlPm3/KCUVyZTWfCBBV9wJqORxq7ZTT7TN+etsyPsmC3KjtV2/Bh
5/Jw8VcPj6VQnZ5pHyZizSo6U3R6FJLYvcW9QzwR8i8ufAqGvr0335lqvVFbTS+A
zvs41YsEYIv64P0nqgiY/I7BgtkRqYfvEPir2r3Kj6RdK4TT1p3gWFO2yxrXo0S6
rrKLicNtth+OYlqBRprBqN9U/4r1Phiw9sh8tS62GURisAGCVmQyxDWF+xbkzUaY
bw+F6sXS1aFgv+9JMSwJFugPmS8ZsUxXAef16jHPsr9r/o+JnCUO7PileKEt4+mc
EPQqXXUxVlCT5OkQ/LDGOzuAuxr3UUbmgR4GxXVbAsbFFfWzTDbRs5Ozu33p8FPx
SZYRLZAlH4F7gQfxhHCkiAZOsS3yAznZD6KP/kDTDmH9p9LLAwsTBYoFQqIBzsz1
cwm+NMsFNaToO3vnFB7DxPhpI8rrwvBsIxlQTISJsfXqi3XrKHLxezKw+5u5er2p
b7xVhyA3K1tcsz4rhCM7DOf51vAxr9vWnULkcwGb5lhchGSr/PucZm02O1861oMv
62kXg27pgiaALxBdlz3wgOipmh9yCXp+wfd/k99/ST1W1GyWrephPnE+zsownpIL
4rD7VJSxr98AUUQVxU3TPOLkAqZBINmvRvt4W1Ca2ALzRThRgluxg/HK/ik0/ndw
T3dQBHIBFUQl4Ao0vOoyS/5U7asz2lLiN7Xo1igLcVQ/R1dl0SrJyswejuSIKnzi
igSm78ktFpCFIPCI/XMR9p/mVv9lY81sygOUP/41SGso3ZXi7HJZMN2LXE97ZZXX
8lc4f3xEVD8C+HZYGxfrXOfgwWkNe3qcii4e0C/JqiB38WqJvMfmPZbwMa80t5ic
c9Qmr6fR6zAcN/TUu+Dg0y1z7iF4U5eTZ1X87h6yanTJNTdRgFL49ZUoSauqZ8FN
0dK3J220RK+LTxngNV766eP6o02JfhM93AiPzAqlYStvvStCzeZxlpCOGd+fzTfR
j2z7uBof61sLDE0j4VuKTjAgKNoi+HXFf452094CPY4URDU3Ks5Rjz4IUbEQmtZz
3KyqOV6KF8dqs9arH7J0UNfMpK27SF4z302p/xTCVb6ihDg7zLo7Wxq8F6YRPE2I
8wv63MmVBi+U9ESK/4xVefUtaMvgifmhOFaI+YhAxvxO/D+jMSNBYrOVTQz4w8tS
aS/rW6EH/Rdu+VHR4Gh5MiPs3qRC7R/dpQDbLFZu1HMY0kDzJqTgnYR+kle8hwmV
J0sqqbGBGdpFsyT48OH7HSwA/PJ35yKjrgT99BwJyAnYB2iTcdxEegIB2L4fzS/5
Cso7CEfhc0GLX9K7yyuLjhED1+I54thmWRFpICaUR6+zDKfeSFmJ2jQT9ga++rfQ
74bbXOm1RVo42Q6ICis9iVItwzHCAXqWJ0GymW96P+fnWU3bVsgt5lDaxdNI8zZn
5OguVjchD4jfULjTR1t3mt3vLV6YLyoxdrVA4nSySz2X3f/W/BjALxGRDKNUoihI
0t/3RR9y4yZD7hCsztl/1JNWRF3IVxJi1GJoHw8vW3G3ZFqeJ9rt+o/lCsaRi9Mb
TTYkHsPJj0ZsgRSCyDGtp2lIsvu42g2MXhAo4goe8O7LfWNA3NkYfVrtXr9fZxvR
upsrAvsrKDRxKf1FtnGK6sKJpd4NDKqOWNVdDnUxCfYa7Rpgh+dS1eLUw2JinHEq
kXwB+Jm9dnnlNlVJZYKUSRcmKqlw+sq9COoHlO/DSf7yWOiakPbPbe1pZt9XCdZC
/r1NAgEW1o4o87NymN4c9xislynJkZqai3lsAi8pObHoMgocQO6qGGx+wequWL4t
JGdwCZ7hY5+oM9rKTczWECVw97owsu9rzD0wqy819XnpXaRoqfj/6VI//A2cM0Is
1R2tlQ33nOQelX8uWBfJI5eHE2wTGnsjekjvxrD8nI7abnj8BVsl7qL7mxcRaeTc
SEPDUi6HDJawbDugG/dGwcOI6ZCoXxo/pP/JnAGmaQaaOAR/dHf75gb6JK4A9Y78
IIi7o3/NGEsUyk5N/oqDUG0Kq3J2kVeMtIvjfBJqnWHxLN8830kOT/WZpsgwQ2bm
bdwkqVHBYUN/YIFthVUM/LCA4oPSfDRoU0BuF6QN+brzWI6NKvfKaByNq7gOWc5J
5gI0dIpZ2UuL+5OgXF4zed8CcwY49vQXNKg/IIAR0wMmnDo8xmoX7BcnJWMJtBrv
go5cyQCFchNfsZ8Ugkuh7AwgQltKXGjFYeBaGM99VMgTKpBpFloAO8rG29Flipth
qucFHirCIDYAIS2BQi/5spnPqwYAWuBo/9f2LFRx0QDcAub9LoYxyU1/DcUDgdNP
w4pN9ZBKLaKYgs64N4E8D9zOrmcXTxPCukXywABvUSHsLehnIGrEbhB1ud4jgVV1
/+ga970wCoscVB0jjhV4IX50QLvyZFXJPG7HiawoTX+cg3T56ApwXJUAiAnbU36d
g1K7nHdS2qeCPVtMwN1cNu/r5HNJlELcYW2ve7x4IzgOuBTboefeT95mQ6vAKGR2
HBNPPNwuhPEPR1cFbLnDVfv74doWtCby8Wdi0idNuWFsLrsxtWIZ3IHlZTzEzruX
tEbAr3K1VJWP2RstED/iESv5cJ70CnKQqzscYMfvSbF4N4AJFkQPlvnQ3bQa/3cH
+tzAQlvs7mh/CuRkT4vzMysH5izaEWhJobKo9q3bdTSWACsCeZqCHAqywQBzKJ8F
64fCMKDKjFqXrxQRBjnwK985IvAQanzlq/b27s5uEmwUEO4GtF/2dIPxsiF8673V
6Fiq8q/MP15kf4orgZzdkl3os61B6pG+7KcXtK44+icnHJxVvdqSm1CEUa3yTsXC
h0HAbgD3KZ7/IWor+VmAGB0aYQd3Th8U6rz22iucsOIshBv5e3U6OdpAw1bGWuZ5
JMkWXw16GwalrkmpYKdfKhAKZaNXKKKB3V1OOZspDVPXNK6KgDZni9eNuzTn16pP
+vZhD9qDT11xwPCaFHwsU5pjzng+BKzy4l5+DmP7BfTxWdw24b6SK+V8qZbqpwt9
2STYHc66CxEUy/YHQJ+qmELI1QVu6O8kJwAGuMP0YB473Q0B5XUOIGiY55EG6WPi
cPd1UuAUcnWv6rkPsnnTAze1T4vxvmd4bAaTIWozQB1u/MhM7TY3fP5lzzRjzWLA
I5OWATUzbgtC9LZtv2re2HShqKeFSZeMU9GFR4LDcMl/imhGpDl7DMhakbSbm6eI
9W+tZYaboCK75WTQm3e/9DpSNkS/3iL7Am1LI/xevsD+ZNjzorXjyid44IbVVGON
igDCDSW2DM3Oeq6itG1UQKpT9IMbnSbdYvNpWSItcryXetWBwkQYpaFBb3DM9uXS
ThZZbBQjo/gbrSWTCXKBXtSRV2mq2kZgaYuKrhlXtem7A9UZeKKE+bdL9clUPj0w
5tCQjts1EdkHsar7zXk2eBeZMxKFtsmJQN1Nr2av3H5p9y1m/gyOlmw7OwxNOC+x
h/auX8WqyNy49punxWmFOLGn/5IgcwwSW029fLsHHVXl3X0ATZFIMt1f9Fj9BAlJ
xFuz0mIW/p7xuav+MyR+a7Me1+x6lZ1l98Ta7ldTwxfQ8vGvFWkMnyucWKa466V9
Bl0xPN0S/0GjejAltwJqKr/NTMN03NSMJtlLSznlR7iDqIM0/HOxppF+LVnSblNM
SvLgNDSqZ+tj0cP/NUwMXftLrwspfkDKbn+yCE2YKwkyZ2I0DgvmF7Z67HVZWKZV
FCUQvtRuyo9429f60xATqXhg6Fad8jLb6vfAWAznakDzu7siWJsMrJDJ4rUeY5xM
OeEa/Q8kFHEM8G4MUMkNM2eGquJ3jMOjXVzmg0ZpqGDlnlZFzaLDmeHM6aDkWZoC
ECq/rpAEwVl93eSWI4Fl58fBgMtcq5LQrtyoj65E57mJZRuWDoh1rWPIpO7jfNbp
KbrkOctETwos8Uh+cOuV3PB3kHBvftAn9Q9eBmyMsd5hZw9YZOvWOwSRd3kcxMMh
sv5EtD27VHlPzDDNG+3X74fy9gWs4iYPLQ6v0Rc+CzZVrS40jgI8zT4GxXeQJr/G
u0b2lB4N1EmzDHa/asLmsgFeoJjWDWbSAmYm5AWdPizZigWXpnRt92RKV8BDQsTX
5tkltnuwZV2k7Toifreb0DoNAUM9WtE1dDYIDtcrW1u0jT9VV8ByayTFd6y6o3gy
2O4QBgfxj4cI+A6jjCdQHbtu/qXg9Cau9A+FHWne696RzyHqi7tHiTnLSOrRmITG
jzTlVgdNxMauHqMIgjaUfDj+0MoSRDEUB0NElkm9B5AZqwyBsfK88oEoF4Y83TCy
RkfytpfaOqnr0ktLa3FubEiUVNWoFC4/z3PZL+ngDFIZrHl1QAN8hXwW4z1JZ7q/
swNKfzReihsLuJClrNpipCZN/srVk+hfFGvrsiIgbQdv0YUNNvY+37jKPRF0DX0H
fq/mwi05pulVrr1nayafMkRVLwtKyCGirCunJtE4+IPmDLU5iuQmDPDbfattHHR8
/5HwMqpXWxWOxnlz9LUy0UL0QZJlA10CK+/0FjV3nQFGuwUU1sPNmOA4i0a1qMmb
c75dYOuJdrtmPS/CO7hSyUgb8eihYmuAYOvteUtfADUc4MpDcqV5fzpGMD9pxWQK
vrOQEg+hzxXDFSpYfDrSWRfHYda7+DNFGoCCHbUNupr2OjCAjPwK5TnDJaQXC98G
DkMArIooI9Nu6XKotP3ciE7bOgXrULnGdtJH3ZqWPgd3Pql5wnIjdPR45lqVuPKH
y7JuM4fOGqG9/+3UK2NW4dGeKyVNu2Rm+LCTMFUGTQmod0H6plIz0+m4mBg8DrnC
2ouLchv9WoiPHrphoV1PUWNDJeDlhGV6kc9gOOnngymjP5XDiSRNXjwx6UecW+Ix
5a3ueL1lMCYBIAFmoBUre+BSZ1IjJu9UQkWtHmrr22QuvIdyYNo1wzCG5MI5e4BW
JK4M1E/Ehm0M2dQKY5tR4AXnifPpVcM8XYAypkuSKRQDH1Gq7/bZQ5TgMf9+S+kE
UNC/w3RJ0NJNtSUqWCZtaeEVD03n1fK9v4g+B4Og+A6l9gQkOx3qiBfxkKVQtYmw
A3hj8wq9quTv4PGARWrQnSjsqPLY7AZn90Xl0P77nizkN1KBGBkvojiKtOemsVC4
9B0KyqxNgrn6ADy9aRufdD2AP1dhFQi2OJJ4a5eixLkDUIKtA7x28IYwsmFTULW8
cY1ncNctOnZPkObAih0pt4YUvVK2jjSZhww2c7A//mzTBKJqLYbXcgHDgPb+rwDa
XaK9COU5XCBkuAJZ20lJhyDcBeNpbRHC8uozO6g9ugEQkOyexiMEH6dL8T0HWb83
9CbkoS3VzmlwdjVBfXIJYqve/MiHSBUNasWQQ7tFkAQiiYafEYcs43JgEX7fO3Vi
GtR/tUMzCdOtWpLLro3oTlgrnHsjQZQdC56pmtoKv7BnI3Rdxa4tOIRxcMvxRmRT
MC1QNoN0Z67c+przDrnjAuCfO62PcZ9P7a1RG71hXyl7ISVXErHmhvNDIlmOvW2s
VU0O9jwJkOFTxrj7PJD5im1Q4EIFJn0kwCXC8sfqurN9hAQXxNyUiqKoozVgJXGz
SV6Nja0CwHO8JUB7OpxhHbaRVOMRu5NKOSN2eT7k/QWCQVTc5/Q/Hqhklwq4067c
ibc4vzCC5I7+TvvPgazBBesG6kNWWn4UU/wG8WkEUnFR+8c7xe3AOSoFeFcNIXH6
LMxj48T8dwo67RMM4XMj0B19Jl9y6XvgPhehSjy4cSHBD0JGe0fg+/TcDnATX7Dr
Q+05QNQUuwq1vlPzATThqH/lxcadbt+dAtsIY9WfLT1taRiMxKlyGsEvtxY7XsSM
yCZXoUUk/lSOZgZOk109tP6tFX3TH+BrM3E9VZq+EWQKNe7eCvHKqLw6FobQjeg7
kU08rpbVApd0wD1YtHMlDFIizJ98ulorM3SRbDe+ub9yXb5kl6rksXFLYXudGgpB
s0kOSbAkOCSRvsI7b4QN9eCgmHwkADyEwSdAQcqEGT4IHonpdqhB7CoQhG0X6Bt6
g3LdNn5qcTTlC/cqZy/i5H+PMZPAqravJBdpiXx4maMGj+BxmDi2TwZinCG+4nNE
FO3UywTJ+uiYjBbtkghJpDvBNTrpCjJNBejUQSbfmMFGORw4vUmfaj9cQa6JI9Rl
WStSc7yyOwFI9INI5br6i4XU6LGKEW1QYuW1iNt9AG4JOQUrI2F6ocR4Ein/oJmY
KsMrQUdZbfV0XCWAg18tlaSexSBaLsjj6pvakI5IDjU+EP0n2sKnCKGXib0I80hl
z90HJ5EJXi2rqzJ8skwUZJlo9SyduJHs3a1m89Jn1preT+wfl5ldjVCUkfKdKQOX
B6dod7TSe377x+jrGWuOTxK385p32KH1F47pVjiO8Sc8s4k1Ht2AqyU7Eks8HFUR
PZDh1MWmUwbgQevIYIzQ0vlItjGRyiqxdNK/003+34LtYm49Za2D+HcDNsm/sziu
yxuberUOpMqE+jT18f1t+O/DmWMNR3Bx1Rj8t4mSx64CTpHA4uetA+7GhPugl/8j
kswg5veXAsqk4a8pnlAu6OfIuUkG/yCtg3ztQaYZvNxTWE2nu6gBSPQ8BYrYNEFS
STtKV2bHhaxhmFlVj0eY0ruF9r48bTvcyKnadjCQTW9ikbiKKXKYmfO8Z3UzcmBu
299Yt4uP6l1w8D3HPfIU7bQJaaZKahdadLQa0uW4V+52w9OBcTaae5SwGKlaaWy/
tbmNCVLvQ3KagTNKuBc3Zjz0F/BRKVx+lDDwO43sSlY8WhaKVzIqtnE6jBcOSL1R
qls6NCAo9MMC9JOVmYjLPBloIbfqSkd0DYKzMDXJolo+YCzfdv1yS3y088M+iFO1
Objjuj4yjSRYW4PqVq0hmaRtdLREj5mab+hwm5Dirred4X4r0rTTv8ijr2oX7AqW
Ha/5ksGr7erL8jpIL0u7GF1nEsse5f7q8rf7qEYyCElp8Jbjlf3pCo/+z5EczHDh
OKdOR5jHCNFQ2BMYbkWrVzcOQyMjHk1RJlzsN5yihuavpwL5F8TH9zSe/feoTOxP
ZvEM3m/1/ZMWaONtw/nR+otVHAHoZ9HCykdCKBsyv7sA/6sfn4JomphjWNt82arN
DY8a5TCTPPGNSDioNogs19d3mcewzZpqNG0nKi0vDJ47tj9b3QLN4/LLZBZtoNty
hzlOTssDRTeOlnQVck9/Rm1G0KICXk5JMY6ZwQqgfHGkpS7s7A34qSvRoRtkAf+5
bHGSrRqh4V3p2/5F26ZSrD4TMABomABFR4NFDtTAT8KE+ZOqWZhFH43H8s6bkwrc
dMECfdb6klWeR/6ofgBYFYP2/X0IMSk6DvSo4rA8sD4+seWgpifq4+NYdAWGnTIZ
7ZwZJrygWTeYXt7CfdPBzsbzR+lJwMCHpVx15jJDSXPi8g2jq41TDiBn+e+S+dp8
cy/9NmRpQugWdnDrbLjnBg/Gjn31w+8PQmT+FWr4ubEvOheuXxzhRzrAl1ae8AwV
nyGeVu8EXPy33cZ+lu4DsU75MSqmGoux5u9oxldyyvaeYfqXzyNhuaMeAlygNZ9E
C8wU8j4JVb5EeuiQIknVYqyZuEw61bDeMvBVw6Ac0dt5jZkWv9ctfufwEyVD35Tq
FF+3E+KYvblrG8Oijf79MfcBBMoIx2N6HYxfdp4PaEjDDmWYVTvzsq0WfjAW+ZlH
PH81F/nEkGfz/PfKZThjeuULAkmLrVOH5PiW2Z2BT+xDzHg5jnc8JbbTcaLwDlNl
FFCEbnlVgNpcmGJObti4x6lSi9ofIVppEDcD6LEMev0j94bubQgb/Ai6IeceTLjV
M9IH//4nUZB4aw85KaEPh+CO3ikkdVzqfptsyUIv2oeKLN56nK0zHFIa4hkC0o25
vXe3J9icT0cUIqVmRRsrp9mUGWimRJC8XmYd4uEjbvi0RHzQ71X7AXhqato6vLaA
RrS1TRZIuAMRd+EDWAod5lU8mHm7kkHskGgVyNfBPdPOvuIIUWUG7/ZC8EtSGIg3
lKPGXUJK3/YLqAK/Hc6OuxkeHe+MMKTMnLbLeLdc26lE5wlK1/j50WVqsRReqo+C
Gm42jAIEOf0Tt7GM0/7pE17NZfETcLDkCrvY52rQcjq7vNLxjklLoxeIR5CH4+Xo
Uo0gYseutKdutSafcJfpBTD9KQeh3PRwVcPx2huc92VYVHt1SbOeeOOZQLBR/RyS
xsq9uT9nSdNz2HFK7fdDUEcTElTNXh3/MKioGx/H57ezSAwewz8BsFcwS2n4vfMw
6yo767oRftBRjkGnKpQPBBOOlO2HzYrbqr93buveEOWkuUPr1rGAEcAdGFMDN44/
bQbia6ctWCB2UjWyypF3Db/RQpON5LgLtRp6rIWWCOqLrAb3lA92xOkSWNfi5JKx
vka9esQM/kAUx6GR+/dGYQxixvFn8dxiepJtwhSwVHi30gHqsKRcwxUuWDxgjrdI
NCPV5GnpQDjHjAWfF3SaWfxBDYs1SkJFI/Tp8N7dX9TBPNvzIgKbArqK6FwqC3qW
0fzUPZDl7qL5gobkE4diF/y3JaZQOYbZZaBxqsG+s1Q6mUf7eyJrUIe2VcwDzDUR
KzJM4N9u6RJjtN5r0YLmYbxjtqGNRIiw1dPl+fWAruK6COCo1Qqiu6qQjQ+eJfdg
tB+x3Jl1FfaS6GlDZ+aM2N3Q58Ljtn/alx3un7/VSSWX9EvP18C685OEbDHstYlS
TcFBokL7QNBLHENjQFbSTkfOb5F18ubBx+tfpXpb7LXFC9lUnXZg38wTRnpEYval
41dopR1OqqT1pLwLDMnu5gb8uq6KyXE68xSxQEHQDIjovdNyWzgTyeRO9o5jgiBy
h0C3+KWEpPhSEDvpgx1rUO1pgC5oZR2NB1CXALppLUqeTsF8YIvFXjAH42ke705E
E7WlJFRxPISrhyx8dziuMFJxzdxuQHMa8VdZhwxO8XLrbjI2+e2G7Ny1/6WnphMd
16tffjptNSn84y0I2yTRnHz3iT59erXKSiL+U9LBUi+flEIcjRcgcrprNLU/i89Z
bnylJmS0p5bMfTTF4Y+P8C80R+dNV2KJ9b3ToiBYfBQ5EmwAFGlgx3mVHbkbIquk
W57X6MWNBn2WrOPFbq3Srr4Znvcm+TsQxkfuiIwu05eBNDIZCZm6E0BiAp/Q0iup
7qsTpNE01syhRn17SZZ+DBlEOlVr6lf6Knv6vzaYOJPfbBGOn+Zaq3sJr+kmuMiH
EYnFUcifjHy/2GBGYPaZrJsI6sdqKh57nWfExodUhdYKwKE34ZquqmXLzBUg6Rth
g9Tw3/EzFbuisYeYL04hZEZvsNvgLRY36RiNsRsyylnDOQZ0lTfCQb3CeX+7wBQy
/aSotHoSfyIvSCKvP8O6eU3pS5iI26HveDpchjImds7HP9oqR5VB7yV7PbNxZool
Du1WwFCHCgyHWN2MZLDfv8Jl/XnNHKgj2bP5/2QpIoa4zAbICAk3k9J35Tk0fj3l
L5SHjBuiEMuKajUAc23YGtIyxYDmkPfJ+ysQZWe+I0+xSg3DIhZ4wn1hCT/rDAg3
Wcxmh8vmBzO9pNAnS3iiHPJVwq98q0c+fI4bBkolDNF83QRrwHYFu3zq43If32+H
KNYxh5J1wdQ9cXdrr7LOX5qbS9dP9Zjb1iabTJ+HiuvIeGIb8N3/AGb0WgnNYrdN
DYrJJz7w2uMQqL7Ff3APoeC9sMqAVg8RxEowqbhCwTMX2st2nAA/kRb9MArCXNoz
qoJFXFIDAz4OCy3+MRvfZf9/4gJO2EaOubf1/g+EfTxPFKXWLQ4K8UZIZ2WEvS8M
OW5R3sFCLXd3JqJxr6FCXSzIflPD9Kof+MDq7mk036DMp2XBr3jbtHEUJpYPEfIs
KeFSH5VnvK9dLoKpA7oKMMvkyNap+q+c0oj1FTSpsrOIK6PcOQvBKAofnap99qCq
522N7v/Yl5hlYRcSevA2PL/eIqX5byPf/CjxmYDEbVtfhKWdo2wCwVuiFoH0To32
I7XH8xjY+X8bxKZ5YUktnWlbDPfXJCaitMjV9TMFP0e0rOsUov3sJbcKtmTOZjGB
PRzfm5qvxyCDdF9Ok4JGQ67lD+u2Bfpijy/7p+wtzbdOccMKFXbWZVmGVYwZ3um8
45YAELEkYq0+D3NN4hJFDWdpfKZ9PEU6o6AvkprzTwGiUVcftMc7B8rHUL6bqtJT
y7BevmqvjIeES9ccjPoUDAabBWQxh7QTnEcrEPAT0BkEz3oH7yXycbrGrlacJSon
Ch4xgF6R3Bvffp0uHjv+qi87w6kWTwMhj+etF3pRwARERIsOrMdgi7lowyEqLg3n
4SCfqQWilb0d1lN4La1PWadkRkCwOX/QNUomioTymzxTQ7gMMPI6q5ADWdKc4sgo
SygcCpYZfoRGpS0WEWiR+BnKHU5pPMCaFxSkuMO/MrzRWQ70z9nPmK/yGPYIprMd
+xhpOBqYdSRom94UC9e0ayJqVEaVZd4v4hzIdnj/z1CqwIvQuxzp/ot0dT7TUx/h
eASEwZADde5GM09K2mz7EkEY6qvUm2w3tgNviVwyZEFi/OiwvySbAR44jkGbbb52
9QRLuBAPKrteGLZFBDKLVm3fFoUpnotYiHCSRQRGlzohf41jp9cdPLydsNrAVX/q
9VqhnPBtZMmmVEyrU3P0TkXA81Sl2IHZFg/zK63wRGx5qdb1tIOejPeKjb9FzxsZ
rtRVIcM9IxSgdXyP5fxu2zZ720P66bBK3EaVkA4xMfDywtckGjhGA6CCMiHz/kmP
yv/5nxQE9/KZkYjAG2wJFFeo9S4e8gCcQrcc/ll/Fp4K2GNHjwRfJeSk7xq9c1ia
dJQZIeb8htkFrXlEojqVjzfUMLUY+I4dcKSYgoHe91aV+4zZgR8vu2WaqVrD5zJ6
+0cLrlKbMo8xPtqnF1NLX76odswIPQVynfWmSfYRZqx4CHwgLxD8jwbxVWDdmVyD
yzr6s01FeebhZtvWLmn8MQc9ZYNHtEY84OCXHgWH2WaGjVTNMHv8QzKIFKUkJBxQ
mnnq/X8VyC/U3nIOqGuv49ZM0Jg6h1QVBGO4k1Qnp8UenV2u69bP0YftofnsPC9E
mvpkr6IeDMINzkNxN2k0DwYebPVjN/Labx1avhfJvfR+mTrH76BxjG/ErUp5YGLF
lvHk6v8OM6SI8pmyXAl5L4xIvc2t8aN1k9wtAVjqIO1EifiAn4wUUy99Yqw3rTj8
fZ/TCWlKXz2f6qXgRVXX7F54pgbeqr8hmdi5IFTaXmPxalGS3sycvt2Dmz9gQzlx
Vl+WBEVbEU7AXXKPhYUhOHmaQDU5V6AF6MQRE6g0ODZHL/S4QJr6Piq3DqjevHjw
RwYcjkLW3IHLyjdID4/ys2WPTFdw60IuT8d3hvqFXlMKNIx3vCUMcRnj6cZoExlG
Bs4Hnaw19zD7j0XDE78FOTGXK8SFn5FQtj8x1d/MxorMmCx++8KVD0KzwkMm+Rcq
vFnfQNLAYxzyIervdlKxzYNrzFYKaXhH/Txv295uxpgDdTffedELdFexbiud2bY+
CrJIwzfdnmO4oDqCJIezElR7BAV+YnTh5GI5ti8NjJEhV1LdgYtPAXXOl+WpAQtm
aEEd98y9VVWr9XuD4x6qXElvlYiix+sklWGoOMd1pMEr5q0bsR5YeXQATmHJ7HY0
4opPe4rG+qAvyBzxSv5X6dMA7YRaWvxCCdqrIxO7BRlZUTFhNCiAcR3KoOPBCDHN
jchP54pdgdIY9UfkNlyQwTropn/3j66vumadCFsPvwJW8hIWmaPSsM4aEfjW/NGK
mmRrLS47hThrmymFAFC6pgxQMkySsA9Ov2IAlWc/nzs+XwWadwqbBc23bJzPxiO3
BnY4zcg4Ma4Q8hEINx0VY/4eTR8lQlHq7r0ZwOVbxbzgnzbAjFcLq+wwH8l4XdsI
G3BEx0eGkSXoRn6Su4pqjs0qDugCERce8KmQMlY1+fYtD8tSgjPOztgHztUckdAy
Nmfuc7tyDfkPpPXNzADR5+LWDVoLGNTWsg5MERiSiCAQ07rFB1mzsBwERiS9bZbZ
4kGYunyEWYowgm9lHkiyE/1uBmEgtiWoZgUrt/1DbvQpZ+HxKTQOhhRjzw24j0Gc
xAHlkX88KBgh72AXktKYLiaYpFysMutpLiES456JXWjhjO8cdQ1Abb5kEJGzKrC4
1lDzq03u7sJBFdCq6kAK2SARF3w3zn82WLfXcpuT3shWyu6hm5spcmHYRKgTnS4X
iUZKAXSOccOh0mbrLOX9nMFweBOpGzmR+hddabUPE8AamudDuG4zj3NRj/PsdQe/
aajHPIJs1IpRFqyb/jyFTpCu2eSBboTtJwA+K22KW7pXV4Id6afqAOlsKWtjQto5
rlhuVmCaEfnEzVhrdRSWmIlAQxuLaxmV8sf96+G/SfL1d7OfEGdBCsTC7O4DlYaL
05TvBvz/DGZQV82JcATvB54q6HLhBEuOWoB3LIaqivCAJsg5hCNHMnP8vMvd2LY0
8sOd7FMxFtIe5CfntORXo2BC16MOs1Bdp9tLrZdQxC4OvnbhodD7FmzHMTtiP89e
FN2xHjXoIPac/Ahxc6cDCFWC6pNNux7VLHDYHdahHmRD3T+BC7iqw1dScKHmThZ/
pozfDjyR+0ufQstc1lkt04BYfJOw1Km5EuehxdrZ1lupKkfcZYX0gaDs8Gbmnc2z
3R3jGQkZ5nanvZX0l34iCpjOsLdRN0D9XbDxyltYOf/BYtM5bYlbB3WbO6nHY/Ce
kP3OOtqK5LVdgqdM51IYnKDz+4aDhfV0miGatAvWkimvcXdduk7V7Bexi0PFadXs
yzXd3qtmrjQCJUN682MBFvVkNsULMmyiGuKzgaASZx+2V8cMdVyx9yNj3nfQHUyH
vnXhEx+cmOOMOzTesRozoaOga/HDY/090m+jMqrLDmQiAMYpt51huu3bv5oCAbeq
EspPEFnmMUIHMrQhHeB0FpJ/q+hhymTSUoXNl60CEmMgfOpWlitRmScZoUJ/IFOO
Ci+R8pi64/dSP4VsT0atFVd45HwQE7XQ+aNj1xzleMkCaYdOW4jm4cAHnjXFPlQ0
JLCIEg0MB2W3YATd41FCzL3daHUnMlktreYL3OfPSc3S4pkML/s2Qe4NnZyDgCN3
WepS1JDPfhkwdAQMoJvI+4Ki3noi9hIuPfGjGMoZ9vn2nmK8738lSEndkcMWJYXo
84kl31pg/mAr8Y9/IbcvqN+OMGJWz+Cu5Bp7egmzQHsJq9xLe5RX9iFgtggdlV/H
3ztGRawhvAqgcOi8uQ9Q8AxsMMhtUuG5SyigTWommcrqGJZ9WpjGQJ7BNKEdFzuJ
LxlcYEOR5Iy+NBqP8FVOcpNw6/szkAZQDh2yeJCLKM+BsZXFOuLlU3ghhoZqNmAI
T0WnQ6qMpfDb6+VbrdODMp3WSUwsmek/N43fDpBmdiOG1KDLOj5eHqc3WYirC7oU
g93GbHuIF/ZgAmqCMg/B+IqrRZ/dwLxLRsHkiHgfZpKI9LY9F0ygnfdGGg3vkBMN
qEcjz/KzfTq6ZETKfset5MtfS5iT6sQKB7uJJpwwlGOnXqaUQLZMCO+zm3rvEYpM
E0i+USVfbhJSUyktMWKhsmcJqTL33hmrg7Tor/qFbfggZKvrztnGOZARYAr1R8+7
C8YktT49yGNbuVNgm3GCAXyVvD0vKxZnVblNx74vE4EBzRzuozjFOpjoNUupcBQh
9k6nkfo9xNw3ZuPGucuivL9tK9Op471q9d3PAwD/z6869fOxHlhTaEIb3koui/Qs
TmAB2YugT9+AojovP0YLKXMz81vGlbKxSHeoriLqtOoG2ZlWVQkET2pwG0aM+I+O
DTNtjYrI2N8em41byAs4ZokSB3TcWuyUNIV1iRWQmyXwMcxuw3QOgjR96znoN/hf
BXNwNzZ0ENWeO2QsM75O2hjzBhzc1bsE+vu1jRqnqqXWenqVjXC0e2ucDr02kmas
8tjUcHBywZkNPxaDwtJroBc4Ndst0MQeXbBjxERuy5+lmcd3us1qEp6tXFPdBrOA
6L5ODDQEB6EVESm22CDXQBUaWli7uhfd/oMA6bO5lGa3+eZf/p990TQeeTEvmOMS
aTJ6/7IYJq9tBkIfLDiINH/TPGzuOwChsvxBHYBqJWGtL81hEfCIGL8PMishVyIo
Zc0BVRuy8YOqjX90ySwy6FIHKtSipZrt1SKh2cvNCwiKG4Zj3n7LlGuRhWyhBYkq
0oa861AN8D3v4QNwbo4PXPclrYHvlEr03a3LcKIYCZFr4zsjNkEHFYemi41gpzW2
1Nlzye5UujMDKcybBP7FHw7It5nl2sD2mFWm/Gm59qpczFrbg2zmUwdFHFQ92bTt
ezxGMCnhmjbDu2fCykg92L7SpZ0+KkfrwOgLtb568MbpxhpcisR4aR6nEUSxDPyJ
AtQMFP7Wp2MMAN7NjRITiM6QmSwd/yv7ADglPsyxok1fXp9fhtGoCsq+a5K66M2f
CQbHpu4cFcURX/yWl/XOI8wEzhg+DCmK/Q6wTnIuXRTqt2VfWSK6be/iwr9u/CCN
eDGrs1Qu01hcqiDVsmoaPvNOfZ36IeJad6P8cN+K6L6eBgzBuBrxZWItNJeCMWre
Bb7IzJplSoO6cNPWotx8LXibcA9MEmIsu47XqvTuyIQCLX8v0avXah8IkZEyicR3
cl0ixN0tuAfHC904MpNHbyYXXo2051SNwHXrkhM0Y/Sci/gr5//76Zv+aeVPx6nR
bF40CcMsFLTrIoAywMdtFagAVHkGuXxEVNHC0sj6A5CftF0tSOfKL3Kp0kpB1gRk
3IiGO1rX9YlDzeo8Yk1qKiPP9RdHY8GE7NpQ8esHKTI9vlpzQFmEW/9u1jc/woRR
4/xKx7oN63mK7h1+6+8rsGP7N8uB+Yry/sa4wATRNmq9STuoMZPwIFj3JMrjtCs6
x0oLe4RsvtB2sMxJKcAoXeT/EX3NBwVBtwGgJnCBzIgDaW5jbcWPriyjvgaTVnmW
8kVkUjASSOkZxKmfKe36EGLkXzm52FSC3eBvGCb9y+qUj0U1rFawgYLdUkUQMwxF
imfrk9gDdTl0j8Kk7+rW7h2H8k5otFclkHLde7/jTjWN6M4vbhoD2xUUPG5I8K+G
v3KiE6EAjOgWvUaBCJl1EB/kM1szbJaWS9bDU9Saa0zbjcB7yVC0B5ngiJWJkDrr
a1UI7ofB1Aqvq7ICGtqGGT4TfPEgVHfRneutzK/rbPaFy93vbCYtp7HoLaqTqDkY
6YAyh+3n0gj3vRSzZYnxSLipWK1r4vIOW1XgirlN7ulM0v+jBSlXt1npEx+cfALy
Twyc2yL9a7gcpr363u/MJTS9jCZZ+EAe7cR3fyXjVuB7BOwKZ2NuECASt6jGDs2R
340n61CKzhBhklxa7J8GtD3agsF3rk/bVzDQC+VC43uwE3edHjO+KRy+2BOYQZL7
CwTMy2TW14h+R2rxs/kpv1p5tiRB94qmSQwg9xgiWmesiB3VwfE697ASmzxebC3L
9pvDRIOrMaCfOTfBCywEuQ9c3wTSHePnzoLzmnlEDc07GtKs9CrYT4tVg/Ljzixr
1/TiR0XGiKqWxqErsx/vbFh4R4jklqh9pKnRmDuGuft3tcTJUQZhI+y6wSjs3PF9
iIu7lXbGgyYmuxw0bQ0Rllh/UV4iuDvtgQO8QJFmu6XaOc6jc73hy/Cc9nDgqO2W
gJuW7YZ2KWsOlr2pVe/cVwnFJJym0yql/rFCUyB/UFBx/oRRfeh2lHCILL0k1gtJ
Caf4aMMqO32sj1PZZMSgjcp24wRA0F8qjCcl9iEbHtMA+2uY9C4yEV8MEcNhvOez
BAVW6rCIWhk5eGvgadEL5+OsRc7RpcpoDI327SnDIsM/llV9p44QOjKZMHYGBKtf
om79heU3AkaKn0AyfGcJJEoMv37zdycTuA/q9pHRyATa7wi+rdvPMiIFKnmoMlfF
NSRcH5UHvijvHtHDhnFtRxJ9gUY8MbcL2ct/BZHePmWEwKykkl3VItvv4/5ftM/R
YyaN/x3yS7SbcHyuSs6BelcJ2Q8/dEBztczjjWM9Kerb8OLiyvWyNPEr1Nq0jOLq
EkqFjq8iPkPQxPn/JHs8Q9bNOh3fhevQHUNNsPjBxsqsLAJI/zdm3JYljsl/yyNJ
lBksRO6qozQPw9p9GxK5bXw6fuaVBwEK5GnaJUbtFffifRpkgTnqjYlf2t7h9ivZ
TCox/RiZ3FICRZNCmrWboYfmu/LlIfKRRXG7BMeZKlx0j62QRXgR9vu+yP8CXO0B
SqVEFncbkoQsBHhqCW63NTs8gak8MOA7NWqTRV+YvItBw4EajbhPAEBXr41lgckF
8/ShZXX4ou4poEzn84gCMlo++NpIOEhWwoJnzy5lnRmP202W2yI9rHNUdXUihy75
G4G+//YG5VGjf1yxrahYhuE2YBXREroX85FPIN7ttB1Fh/3ePclkCZv82jYw7gt7
4PUTbkMrwEqaLq7EJzUAosteSPxxfWyjikCMe7gRQTiyC3CvOuuoNB53OBDH5Yol
5tzJPCm245W4Bk4O/IpZ89B8LUvi4FIIsGw5vlpT1GVuwkQuhVf6oA9QSf03h2o0
rkN+WbHL2NBODJSizIJmkan7lW6auOoIksEj7cPJaFjiNo+KCkcbXiDmnVosmlDw
bunxlRqcwsSl2PMO9B7xFSBzHTCF6DM/qGGg+kkbFdkJAdy5H+/lbtILwzimLbs2
PUMkKra5y5lTXHzwymEGPJFrk2kZbKoer9/UJT4bJUjs9THxujW52csv00rnJ9YK
KOb+jCEy2Vb/uqcKnYznddrjtFy1RsOO2AIwzp7Bq1Ow6bthJurKrWDwSbWoFjiU
Iu6FVvbgBNnPqfh0bbAqu1wM660m8hhjrF2NHWNM+m7rU0g6YuylaL8FJsZ8WgHx
+wZOTJvIWJ2mioe1aPvTu0u5EhBE038fTK1vniuqyU+vjzBqkBuCZeku4ZIdxVYE
KTJfjYXmuTHeQ5G7M6K+11NQ4aRIfoVu26n7balv5NO6w2gFjhkx5NKZBuKCl2U5
ac0hRDRNUY/pGJBmRGD6+/wH3CE/8THYd19d39xGseGnuG2Npzl1qFpcutUfeYAU
0VA3ePkdben9yNAW2C3Rt7dugwlQ7dg+iv1IU+fAlA49lsX0tKfjgaegmnaknqp1
zpuX5K/rzrI1DkY9JgQzOxAqDtD6ZM786nijP/sbzZNlWKB1yvCANC3ShiXfVNA3
NzZYoAYPbB39lf0F99indlLwIRiLbjlFJEVtF4pEWqC0Y89M49nBeegphqsUiLGh
VzjrAQ+LTMdSmZh/wp21r5Cy1DLIBOn7Ucv53A0LCAJpAZuv3QwnE/GCdNemksyD
jQD+xjRDALeWzs0D2ZP+JEvD2K/vgB5rWVm9DdF+tqWZhpopi4PSTKZWwliWWztj
bMZIPO2jB1cTKaW2OzPQOzcLeCnP74cWJVHIIr6UzHR3DyfDFc/ks/PZqEAQLuqI
z5BW+I2ZJby1OQ9sw1u4KAsuDCB3AkM2OBJI1Cf6Zuj3WRP3wVeyzwES4NrcQKpY
4joeVG3No7JOTgJOyvZX9FRWvTBATsoaQDxXJqWxT5E+y1SVKTQ2fQvrCPazeyPI
i1vjhbd+sXOlxGOd7Fn+M8guCAOTsToPAwE6GlGSQvwvm7Hfka4QFrJwfqcQENrR
2bkiORl81QKOEBSNJl0tODL0+K0UetZ+au/7JtkQ+SWF3jV8IrH3YX+pQE3ePliH
oEcZm60Cu+922/1TOzLCTsVc+jPjMys5YpRBD7zY4+bLNW6NmFLIODaYXp9Z+gth
vB+nrsEs6GB0xQTpQzGhg3REsFBFGB9DVLtEOsTlD/ajPlCmRkK1BQtiYTNwzKra
kjW/PTcocLseMjrY14Q6UNi7W+5OI+5TgG/57pbyH3CaBA3MzbXfqPjU5l7VsEjX
gTQxrjOkguJSGGrzjcVzqwNQJXp0UkbVMGMbsxKgEGswyOyI98ywOKtGmSUoOKir
7vfHsVzv2zjf1my/DnwwW0W0JoAptQYF5vBZ5TVdv4/GUP4pNdkvHYY3hdj2sdg4
XBRJspNGS4M6waLNhj7ZiZkLBAfaRtCDvYP730uwVYOqyM9WiYFIuHYAwVRbPxfa
Kr0gBR0YOrpz7itAVMyyoYGfBO5Jtteua0VaPObqr9OBGTEr2o0IKXn0jQ+jAKdF
u9I+C0BIAuEj++JiZFu2j/c0Hnz2Pc9LdfJkBQ/Q9UcvmtKVJGanvFhJCzYGO6oF
iVLD1Kp1UcEeeFFD0BQWIL8g8UjBSCe7WnQHs+pKh5B2aVnTqvHm69xT4nntbdXJ
qJb8pG9sqo2uO+zYd+xbT3IWzbKQxpe4Mi7qDJuFzvrd3qssGZV4xSHshgRTfgKW
Y7A3U7iWiuRmApO1l9sOzoCCq2ceGjVM5NUMBw0FDByIC4yG5Zwx41/BLUAHLm2V
8Br+D8x1+QhrBH1If4GQ2LuegN/mG/s+waSLb865S6WW44nDTTVOtvW2vNndin/P
nNEXCNhElsPu2wA39YS6QvP11OkjZvdFv61wopPUkaGFhYV1+cMs0qAk4Chp8uSa
t1nLZt8ClibbIcUN65eYdKGDGKtaRZKSIn0VWbts+9xkoy+eEdT38k+FvYJAz50k
1eFnvkJuhYFwHrpCSC7GUTluhZRl5xvTGMR5BBo98xTq3TNmy8XXcmIFRQpA5WKE
8bS+AkzQfJ/6EfOJP1m6hKXW9btGqwtOttIfbav7NTgcxI5cesVNA8WpfCK72fp8
MgPTlg6Y5rRs4fcCzZkM+A3YT8DrMRjbST8c4/rXfQ6I2NFjy72IoXkbI3I1xsBv
jgumkn/AWBvxIf+QF0TAXZe2t4vyRecig7/TnK2T0TZx5eK2Dv7rYRh87l3O49Gv
FN4ac3DT+YdfIn7o39dD/UJplFkajkXmDAwxAtt8VngVFuud0qflbe29nu+u8N7z
3Ov1/vzYkVxG7B5xoFGViaxTwX5/I5ZwukEdxAaMUew0gR/e53c7N/WR0gr9CZdx
CsiiedUUTIBAmSGp31Nvxa6cuPEp/N+Ppf+sAqqh7Rr0wd21EsbPCExvTyXm8Kr7
NSbsHm8kwRfceU/ZTOLR7QW/5xdQ5nMYONtlhi6bwLwsRDk+cHcZDUtAC9aURlYo
9Cc9bVv7yT2Xu9zd+dPAXTVMYQtWDM6fK4IlWo1rM7lyrz3N/+xVl/MTjfs3L5LE
8uVYeG6w4mWKIm4a5xbR41yjw+aRfMZMdKXkNw199w6KAoRK2GC4JIfypkjBMTYl
Qt2Q4knjUm34ThKpMP/P4HNtIptkezpBgU9Bw57pH0IblPDkgcTpQOpvyqPPSwN8
fxohfmbUN2usSKhJZfF+Zi9W+thKQ5op0FESW9l7my9f+5QbnvrslFPh/pt3eXAh
OPQl/bh3AtJYWMay5uVD3qt+I3n6Fl/ghU1+UI03m4c7SyDacUvSfzSQHDXT1XMg
sSgw2Hk0tBmBTYy7ODLwYBZ79yIppgAP/likL3k+p64zbo6vCNoLyYhE9pr7/xDs
3dZhgxTl6Z+09JeY9OXDEKQIMMSvufJWEihCkntoYPaXaSljUrC8/QVW3nWpI2lp
lub3QArMaM/Km3u4bO00sIesdrh55WEI2jAnCmGXDzlHegr7rx9ywJWbODfKFryo
OTS/hKjS/+H6NJoQzU83ah/QOk2ANjMDxcsm/ddepJ7nS7Nffe+mSd+GvPtVEf/7
Q9CwzE5V+C3ZrM78otLpihApyQVqywT3mW2m96qWC7rL5FZeIijdJ4/KmX+w2rQx
hcZT087+XGOPZkuAk0QDMDLTbVlC2h8FoZNf0HFYdrjtB9ZWNLe9xJ+aISjd10xE
HJ5SZtU8kj8IO/Cl2BsVf43HXkxaEknC3V8hXjumKRTwcMB3b10rO4ewho1SRKjW
XwuH9I5TU3KWtQ28UitJvUltXcYH4xV3v2yDNZ4czzVwykomALI44RKjarmluVNT
a8+cPRi+FqM8T0P4yar0U/x0vV6zRd90GugjNDT9tCKNet6gwzGzGNHWrWNTGfK7
j/+eO8+Ojrox4wj0iDlsmXCBpdkh3KnQKhdGGz9gCKHNtBmkMOnIU7R3vb51/GM5
Fxt78jfLHV+3pYFC9zHrD0vBUEhAalcHSDfADhQ+XA4ozqrlZlCsxQVGE4GbtROW
o6acdyuldhkdnVyRwgYjtGgTtuj51q4jDXOVCzfTnc+gbpdNerOvZ0PutwiQzDxy
Re01WqKUxnCu2VcgKmkLB+qxnPgyTASUqYP7HWz6uNSNrmYz59xmltJ9/a9Zy41f
XRNodAMgUc1hiewU2Sutq3/dYzc8oSWBxVa10YNlDBCbn49vLz7fDBiIECYxBrph
IgXVcNn61xq0peabh4pCqMZ3Jz2MJ949/3vSxSB4An7w5Lwx9pKHgT8PmgIDhggZ
Qizk50KyCz64F8WFJnv0XjiB0/hr6YPNMGnflUhxlSU2fyRrSoSsQYH0Mz6CudUK
bW4dxZ/+TSOsCAQ9+dHGi9FaKpI/Q3yiYcbUdXwK5TIadZhp5EtIcBTIUx9ytghz
5PuM9U++6uivOJqTn8RDUXzLSIHkIjWiXAjuRu7ymLl37I0EE/dESSV3SoHNdwAg
5RRmFEzDTqfvWWn4lN7emGA4yGH9PGh2W0b5evn9et9LiyK4GXSPGhRRtAVVNsec
F4kVjbN51HTsExZZ5QIKmnTvTxupWNnIN0C54BbsGouFG/mKk10xucf5i6AfocYb
BfoZsQQp/azSho2ft7ClW6k+3ad5EvwzEdWg68qVVZ/kJAwJvyWCfITn7upNRY/X
GNv9p4AbDqSX8tzMt1EmRb/vySUs2EvBH+NkjPIDgkol+8/ZTMXmOjCYe/FyXVit
YMLwFUr+Og+TnZJ53ABiEyvmCtybwG+jakyPTJCxQyWPdmVVgvtqHENe7Q/5F8aG
3bfsVZMFyTK4+OvIDyrXWSwQiUgI6YsukgMwwT0jP2JH/7sPlPgrcd9lklzFUKX9
TtaN56bfi3MI/ONLONW98FAYJJAUxmS7oeyPgpraUt6cNYAyXJ7iKGSrpi2zQ4X4
1QeLTLWmTvCvvvM2G55iOpk5C2V3XgMetZgVGsx0h2ra01J4PDnZJmEsMtM8747F
PjlLTq+CQ+/MoXjx7XARCZ4jFNktoIhAdspfdUqOmW2AU77KMqG8ZVQAmBbAhuVW
TvItrPNiB0ZiMCi5fGILm3lG2dcWK0xFiitqCE/5lVWaue/21BEdvyvz0RCxuFZ6
4UOH6QeRLC4UbHAMf5DHLsfoLKCkZU/2iUfO20ckUSeLMw/4DVFNwSImYY1yHbd8
Iev6xwa6jLN+T8U1yeR550DGxNL6531SKghE/e3GVhT6jNsvU1V/EWOA3PK+sN/O
JIlYMR3UKBe2Lhkd3pGXr/S43BF2xLBedgEEKvJI1rgWeVq9iLdDqChBPu0xU3mm
1pvzizj9NFD51+hIlMOwu72+6z0HkKRPN2wGjxqrAp5Fu5FtbbjW4in0ug9XgJOH
qocPOrXxUmyWgBKLr/D9FRfJSvJB+OW6EKkhpg6OMWdEsgXP6RdxYhXcPezptdHj
9IrFWNWlIvp6LEUjfSLgy4QcZE0VqSO3PfxB8KJAnTxF5SMsptUFQVouDx3RKDJC
sMrJdERhS8M92qE+7Oo9zyAcg4FoTI4BisMMRdo2fn03z/bsOVWPNzqEyi+dK6n/
2vMRmAGeB5XqexHIGknQK3EVdzMQVfJBk+srw5D0LKVgYrM2VYueCIw1tIf5sUG6
0vjeSbqUmu6wjZi0WNRaGOZF4ZgRvmZ8oOYa+xhFaW+5xFSvs1JyXqJKuzX3Qahp
LW3r95Mc/BFrung7hkoiqy/xS8aRLSAT+oiX9rYbhlAe5gYFi+2N0ftqZi2kW3LO
15CvYmy7EGDAIIl2kb4gH+8F50lxvapliV/hLqxtC5uRThIO6hlpk2EzXP0FC3pG
fwUtwto4XEamn6TszV0rVxJ2WoDgW6QUzvEBUUjFB2tAmIqWCIe5zvzevbw/2YPf
07FWvEMm9xtJuRbeF+5PclTNJCjdh5qgz26k2loJSpe2O9FRVIWuWHEPHmIuhY27
bEbQ37eJFdaGbZaXCc26IL9OEAydXMLEFLNh6I5PYtZNxz+7m5QXXdQIld0Bo6li
aRt8CAyJzCfoS0U63q34857rDjctY5lCwAta8cdQ+dS6kw2r8MsGs966kXuw4s7D
z+fJaswvbRwNEpBZa2ozpFWK5IxOVqi6pdJT4ZkylHCStVtCdgVREVLcZUvc7HDD
DgwaQ3GHThMYALW0pz2LDoZwJ76mdMNLVOpJ2QFsCJ8wcyBj9ncVBgGqWul8oz+B
2lYSmR2kxxVHp0k99z5F3nt8qWw6FDTRvG7hyitfWFXGdwTRL8pwwJt/yGwDHA4e
3UGYWZsbxPwWfH0JSMV6ndGegaNg671zwyGpkl4yfYnMekpBs9gqrIL+tFkEB073
cYJn/3atR9htKG9roLlBaJau19doQ6S/ENWhUfZFLAUPL1ojibRH/c7TMMLDqThX
msrj5n8jGZgzTKGRBCozfuSsxMqaGomeK7P13ConS4Jo4XBzAno6cZCOo427FoMP
lHjpK/SZHRhBibwLX493wGzyJD8jwFhbgAl7vnGc+cfnO/OWMmPuQfi7jy7nrdRo
qhsgehkprDnTqE+62AKbEFcF7m9J4MrErubl1VG+hA7aAu+diAaBwtMbi0Drq/7g
9UexqZxV1t+T3LnpJTdf2xGIfAEc/OpL1y79Ic4m1QtApxGDkY1855ChjAZ/DXUy
NEKemt1P4PeLCLGiFxDaiC2t0tg25jPoqCdq//Nb1OO4idVJFCbMMG+SdCJyEs4O
CE/LsG1vKlpIxMVM5RZqtLno09SN8+EBZo/Jm7T763SG9FgIFbKsLKF/jZv9QCst
XkFEPYfaYzG4f9c1jL43aFJqiwENCt7olkePsx23pqwr0FcdUs14i1JbeAEfvdSL
jIIZ296D7HzZJzPgcpQLRTP2PG8rOLPDHWlg4wXVR4jozKcfdX5sEDjhX1VEDuLs
c1sqi4Jf18RnWgRs2++fszrd3hapi3wl+nbiIpPedE9AaQNQZlDNGvtKIXaFCAMN
PK1q6by6ab5QhWuZ3K2QZkinx8fBBZvJRnEtFnCxKWePSINDxn3cnSxEveB2olZ7
YC6CLD/G3cOXEQ0vFN0kMHCtbXlsr7I8+WW03qb2guWuVWIwo9DwrUZMhk91Hpeq
esRI/wDYcsDi/opJA3bmneUIEg5NIXvNO/CqRu7OceKbiXirjbRxNBLMWYdC3wzu
gDsTBD4Jhp/NNJQquSmbzhUZtw3PZj2c8F1G+GRwM/u8eml0tMiTIp5y3Bjtvtyu
l8lvdInXYvw51cGKSGt4sQU9noa8sd3B6q0PtmyY0Xys9ciCd1Mg51ChFoPyITDr
3gIajDsxQcczbEN2e6R1eITxxX6Kj61/SV6vJR9eQNiJ3l00OR9FMvL0AwtRvmHP
kt0AZ9OF9/dWuua4amOVrxihtUqTQ7VYlO4/ihHsH66yHdUTkfL3Uq5L4SdOe8yO
MPxEex2xcz6UoN6zgE0279BEzPPwnxbjrYv5tW7uDU2bjMEn5/bEOrXBdvEvHBvL
o/PmuJFqI4FuJSASXxcuOyUnWfqcy+wFbNh4Ln/YWLTy41qroC7jea3aSGW/XIzX
ob/ihgSe2pwUwBhYbEhD+7M1wzDoTAGLtZ/+39cRy0abJsEXj3Mq6npLtJbnW4mw
LhuUG8kFy3/QKhjaKd29WTIrpq+0oalJSkhsiyLYpjjNHuK3MnkZPNf+F2oWe1q7
0DlfUxKufSIhtUW1h1jbmMZnK/B+Agi091uPnChSiM5MAoLEHSDMFKJbGnhYZj2e
oWIxagWMAfIFwTsq6vtuKZuG5WP/cltB/eCAf33p8BdX3GZKlkGorGubjlur8/OO
gCodLYSLr/E9HHUc2zKKzQeqgMAJ7PgFOhMXc+860aOUtwB0sUtVjzh78zBSoNVQ
LuobJam6SxJgSl2tF4Qi4DdHKVCtI8VZxld0vju1bTBhrmDigTdF9ovxh2DG4YKC
n2Fwht2E3tu53wA/c7gnAQJNnxFdFeCBpt9TnHeuinnJkHvACz2agO/nV2Or1008
oWbSFX3POVdxVDGcR6nb2IDA8Ywj0FpA4xfrX36fZPFZAdih30R1Do/PkuPv9xOR
4jBGdNkiVlr+hYzNp6qoukeOhzmW9hHIGkkrP2Hl1W1R6ry/wK5vGrNnRbvwhjD9
LgJSAAurNlVV/TXtxqIhlCrjxkUOfnoMehVbS3bXZjkDX/LZ3nkdlYka8fLQPn8R
QXec4TXx3K4YRfe4LkPmnIzEIzezPcJ+8XGrleCxQyf+XFjWHaswBbIex5QQDfns
dyZHZBJS601Zmf/ikGdLsKkbT1fCwyLE+fSRQWSPh2WJjKS+Jw0CKIGyjGTHRs4l
kz43Z8l8jQC59xzfOnX3hhyplA8YwsszFF/S5g7/GdDr0yyXEzlKQ7IAKoCaNm/R
PAZf26gJjTheVMrLvgDLxb6okzGyo9GAO43CPR8V7ckiog1Y2ZCWKh21Lu5bz9Zw
lqY6q3w1GsKB80l3rUioEJA3e1YMkg9Xn/G8HDn6aI1G0m8qe+taWiL9YKke+1HK
9MoikV+VaElgTzOF4tzGpFMe/P2r1I+vlh8LPxZLtE+KDU2YkhCdfYJtO3/ESTr9
SVaX8LHYJuUQAE10XFOZIIO8waY9Va3+hgOq9pw21noV2LipGWpLCWRlWF9KufOB
5eoy2ijo+1DjVZOAYcF+aqQ1D3aLSYLXekqtE0V7xumWg2lxjGpSpMp6ejBffRCl
JvIKUs7p/+jpH+uv12/gb2GO+1uAwYFNvmGoDNZbtLlZQaMEmo+hdzOUbIyEAbmR
gZreOORsjr+PXFTKlsZ8qnaqia+R3ZAb+SLetbRO+2/4oZxHx+TSVxZmsITEsUoa
IqMScp7fkKhR/D65ahoRPTAafIKMnwtVYuPb9NMyvgbhRsRZ6Mq+mBImyw5YxSk/
PkeFY9EjU5V2uUbg2NtYev6FXsXlRNYQouzbkx6yV86SQpXJVe3IzlPI5PqnDpDi
EDqPyzM5Wr1kZFhaJxF8lbt0UpqPW6xE9GwqVq5fCoTCHX7UZseA9BI5efxrJmnI
3SbMNvrOZKslb54V16PQvQmlgkPG90NR2jFAWkQPL3dukitwzWdDXD5DTd8WQ/EC
46h9SbZ7eDq/J6Pwck8bM/R7QEfVSlGsKmQDwyl8FkTPEoWgH0Y2QuhyzJCCJdZb
a6T2LF2JjgMyHxHi+pgXV3qevnn8IXIi1Cxl6J7ztPWvdFgrRk22oQdb9nAkKxbH
1GmmEHkXolHFckw1WOh1zAJ5R5fxXx2cRWynbmwMhyD52n4typOo3lb2Wo6g3A3V
izOCi55lotKG/6fjqvQatANCvO9kbEbDWpZTKOifQY2I8I5wWx8+X+rzp6E7gNpj
3VP60bCMsUhMs5ONqY1X3RGkZQNaA66wz+aNY8O3DKDggscUdmLZbY41WbX6/XYl
cXTZwn1sL0sLs/iQNsq9EUDx5oCX4hyQQERSLxdK0p1v3dWcy0mSLrCfxSWJQx82
+aqMInEdw9gB8OGw43dvzegbOoWnFOtYsjEtaWLvBxASuSlbwxKj5nYy2GWkNB8p
Fbb5d0GR5JjGJDnVFX+2X+SmwCYcI7Dk1fdwym0PucfQmagIx2nU3iwXEeScdRlZ
CMaYKCmRHbaGm0rqp9Wvi5YWsr8NhEIUZH2eYcJgqTd+/G5VTNAl1ZLCBsH+zUcN
PNe0QWBelg7rQxdu4v0OPHINAphj6yocEZAPr5S2ncpBddZ3bHizAgz06PPO1Bi9
M6b6CWnkgwKN+RvnipNaxt4piuHPPA8nFCpVRMCBev0E9mqOpfFQnnhoMnKhacPr
TD0CS0YBI3AXiUJsEGr8i+l5lOZGR/2yJUNFEiPvR1KcwZKoArV5XJe7t0SKaAX3
yXInBUglF93w/1vCNifeNgNbSeuh+XWsv2ZbPv2wUX9USFwEFdjNBhbUUWfMtuRb
vjG+m69acEA25kY1nmvsg4pu/jRQ3j2CUAVFFHsFg+k1Pf7eVgtFNQ/s6IILbE/J
lV7So5/MEwhWaGjQwCxbqWQD4Pf3yEqFhWryOlI5Epitj/AauUT9Yc5ReKpX1R3D
UCiMrlCvSrUb/ixHbvMrpmEtryvWXk+mthaUy8KI90WGwXerz4auRPZoG0ZmsCE6
5i4q5p4bLRFsGsiZdP9Zzt7LltOlnkurP4i74KP5tGHfushKtXoBvL5U/9Y61ius
abwkeiIVz9xrftf0NbMJvoE1YEFOcM76QZBVqs3N9btwLhw75MfHSR/LUm9pvO9y
2F2V5h22bEeKj15GO+/H3Pih4iP70wGPNugcnn+OOBS6cW8VCeoIkoqN6QIoVvGO
3YMX66evsePs8shHYFZtf2eV9dgG4GwS0V1hecfnyZKRGU7P5c978T0y84bJmYQL
8Mq2tf89c6vN8Kbq6lS6GRiEZnAQ4uMU5+VFbPGloeKMspRXnbBLwwvkotsFxLfS
073S5FjKENmqXC4fo5LZYtHn9fSejAmMcJv62OlT8bm4gwUm80LUnBRq3deFBEgn
MWkpZTBKxyUhxu3QG61VCveLIARr4OmCmNbwNF9rRKlRXln6Vd4BlmzZo0F1Chfp
7FhXZO6kKwuL4ovlCinHDI0gQ7UfgydRcY7HyH+zZrYa89neseZukz05/3g5Ht2B
wFxmmBeG8/vhufykuBAnD3LMq0j5kaBdW+6Hgi1BrUTBIcMBdldiB9I/d6yNiUIe
Vc/zBhBPGqTh1A0lSgXlvVEpCZn5HKTHylSOJ+OVyJJ8Kn8+Gib6Qz5ykV3AcLpJ
zVpZXY6iPfn6Nd6jmH5n/0XdqQh7p+FHVxuST4XSgEAejO3SdHgKN1/KCQ9c9acu
qxZr46gJQikg7aE4H2bUeQw+17KlrRJmkI7V2yDZPY3pimqGNHnXP+1Mpcfw5dzv
c4eWIdj4dgsXWEAyyMTAJ20n0FBQWcWhV4HJjMLUWSkHqX1+qqL7nQyjosq0P7AD
mSmklXL6tjP7DjoUDZ38gWnwpf2V28LB87nd9YuYiF4suFTeZ9WfJi66vJehJuiX
nqdF7/yD4Z7ybTnJCnleyXSucwFUM3Z6pVD5tak0lZyzuKywqJquRsbdUoVN8OvT
Uu9uUnjgdY4uTOzekHTxPXHtT/qmsKvejyJdOE/hxYT9Ds5ij4skME9W5tVh9pMd
QsA4LYx5lrEU8bpgSELrxaw/oRNYu51tRyOjXFFiT4aLYDxu9j1Y/2TONaGUjkEP
TGf115hfYC3gdZrDMfXgIZkzMrKa8B7e5F9dupZlO531Zmv7c6RQc5nUKm+M+4RZ
7BfJu12DsvgVVbRq7XYwBz1h2AAUv2wuPw0LEQT+ro1Qcf5xzmPEY2yRpO309XFL
BKA+BhR0ABJBhBeWjjkHdhODmT/2zftmvGCPVkEjN3XGcpCOb/pROBFut/+452Jo
v5hqfwzMU3VlKQ8cS3PJ0oSEOPA8dO1E1Az/DzoFN2uS+ZochLftikP7/npa731U
MTBXfVRkmNQ3o/CtQDYQyB7vVuS47Tbc4WUqymZ/HF2PGNwrBLtuYaaFdDXx+qM4
Cnmcl6a7qfi5gchX99BhdU7/W2DsHrRUkgSr48+BiDqp9FHOEK3/4UDkaOFqVySx
6RawiemQoybsYOlQ8Mw8BT8EjHX/bFP2GIqcFjIj5CQylVhcb3HMFqf4w6JpwiCO
Uzw58w0svh1vmRF4GWYU4ItlatIC+RVKPZKc0cORm0V2+3tjA5oe+Lq/TYd8R4Z+
PG/HqITn0fZdMMoWr+D/hVNNZHBsKAnLicjsS8eX/MDq5W9N05vi7y1EE13bA2ug
LIeSVMKJWlp3TgjV4lcbDhu10hIB19SbqAqSO2SgHXaF2mU4I/cl4fiRSKZD0ZgT
ilUvQkGsC3HS+urMdKWTKF8+Lfo6cZHW6h8Bo4klCd+zsce9IZAWI0YyNhIvHw2e
ug4zmDXXVw56kiElSvlJFbAbqaeAev3nkXAjC7hGeA+CO0NmDk9x0IOIj/wVRddp
7xOBwcIObCuTrUaQsdNRgZDlH1tkJSV3QUnGAyyVuk7feNUV0FBq7aFket5FBedz
t3W3JC7PXWnS51ybmdPn6352mKAReF2Ff8GlnOiYRcasxBKNNtu5MGCDrp8zcspZ
FFmKpLyXIUmIfK0wjHRmynC7oW5H6Y3uj1zrWtLMkEKOtP3lHgnPHT73tzD6dH6v
hJ2LqIwdYFJyUeMlSjX5CGcrK7AECySU7RinaIW6GUbhPfq1Vb0/02MYEM9ro1oB
3lqUN9JckvmU155l8dcK2MaFmCV2wPc2g8g4d/lqPkNbByh3KnlUP/gcC0f0kR3b
4in6aFYLwie69JUhlp9yDBOaKoXIZ35IJhDY2GTFJQQDxZ20Uub+lj+cRvJS+UR2
BwyapK1oNTmZUllmQhDCyPhqAP18xFI1HP+Hc+Cx440YM2bufUgWKzXA3XkLPyQp
w2a/zqwG9Vi6glrb0OAJhY7mEMuthnF82wRGbwnegYNG9MfTZ/cr4Je3zv4atEGY
WlaXvtdFQ7uVm3kDOPItW+fIN6kPDaW11eDEiZiJstkNFHYGakM4MGOtx5BzyJcf
My6UdFMvU3vS/+8iPs6P7PrK3x12crQNjINvIuWg4yGB1iLB0Iwz81pLROyaJC1o
Ih5LdhgNOyZvS7OXwLc+RuaZX+JG1L/mg5FUJnw7NoAth03ZmbF/IyKOVM+3NEJT
Xv1YUkQ0Rq73St4fzYbI4WRKzJEh+W4oImTsNeNK/XEVTvb9f30PT0WmApz1KNbi
V9v7Q0V53+nfndTEmjlYXVlBb7w5cAnAyOA6H38sKKKeSvQc/Rgyl4QBtqaCfENH
wLoi6+6ErhenvZkqVkgHKQucvpWA2eqYTgkGNzN1aTt8rYfn2hjbTqW+kEdxDlUw
uNPLTDqHXcGu2rrwdEoHUiwwFU/nRYXWRhBZZZN81yqyJE/bzD+7wxNnGJPT8qge
R9HyHtgCLoPSHDFAxWNFnE6+gSbPM9V6ENlANgSuB1MV8FJb/inbJO7+gS3t0e9f
thwMwgCyW4kGffmgOED4PhQ/TQcUV9mZd1RHuOry6w4f9LeWVbq3WaDptf2oUal0
47Ugrxjq4550fj1wTCGQunPutOjCayZyNPaDP6Lh6YPiGKdRg+AFwxmzCGUd5Ajz
0wt8KGAZncLxF7uAhdSTx+cFI4hKzWrpEyTaCkiqV66so4rvhWFJOC8d/A+svsw4
/C15U8y6WmRTVfoGbqEwu6fN8VhGfqW0a7Xg3KgZeO0EGAz9LMOzahQcAv6Ce4Iy
xvmcmlr+h2y24AnGH8ERxYeB1F8oy1ldFy8Os0btI9QkYmVlYyxuapW+DojKSfX5
09tYaAwzV+ntYA4Igcb08qd1JxOLmPObsrKpLGCr9JlKu58wbp5JBYcQATiyC44j
gIZFtB5F0Fh/Pvo+9cEo98tMLL5gX1w8R4NiseeJxrCvlj/M/rp9Lb+N6bWzQVEx
NdmHeobf+ywF2jIB2Wfm1ZjV7z7LEuTx4oeKUlF9QsZxtOWQCyBzqRwNU3f/y2X7
mhlxCKuKRYh1d4kq3+Efj7AZZx8qeqyb2a3szNhi2oGQYjUHVqBSNTZhcJqIyECV
WWBRKuTXmeyyL4jMvncSC1wl70SeZIeoatsl3vPRD9AxlShCA15/IRzwIV00Mpjr
sSCwYCRXe7Q6uACrsAfkLnEdFCcTl0md2ruIUjgvlSgfX1Gqi/N/Sd4w3ebFhG9J
5GhU5cZ2i7eBKGo4o/ZIjTfCVKedy36ltKmXojKcXnlcm9qBTd3XWESTvBVV+mhU
qFRPPLtjAUMzLi85rJxK9vrc93OJc7pp0aJuLVq0VclUbNsgtYqx/5htXE5yLDBo
A3xgF/rB0rBl75bqzrSzQLDwNMr0vQdBHogdXvNkkDLW9Lh13mFuA3BpnVZvFL78
WRNuyhN7JlGLY75DhMBB+dcY6sP6xnjcXZq5PCQfPn2IpNr+LjcIJCMDe+rxswmO
+OV+8lbl5qWL4kWye2LDqjqriyElGSvJ3TVzr6dYfhAxr6C5GbWjM6Pkgv0vCfQV
371G7aIOaFdQ0VkwYB15qL8jDQdrDirjB+Hr13U4+8RLI8Ar9Si5nrSwvKlOyzFm
umGQdmnSGpGCsr3TwgVOJeQHJF6aBUqBZ6MeswXdysYrRgQEWr4k1qsRbXGhaw59
iXlZ7o5w7KpYDCBolENXM//e1wFykxC96gwtLsPplb0yfNKwL6bblvbuJ32lmxuw
1jmWnWbIY1Q85uylA2lhJ6/l7nNI+u31CDSgF+Uljj/ImGxYHoRDsVBbJSqUsz7q
dH6WYlkOkijD+vnqg7prntTT4wlZYFTo9FX2GnFSaObrBIp0PtNRhjaExU7URwYs
/MSYN5ShJlzRi63oZemql6IC+lJFkwLSdvO4u40hxI1izDsFjVrh8v682WtER3+A
ynw14O3JtmJLAe+Gl8KmsoY2yc0t5cK+nPM3rpanC7+5TmtYXmYdDVz3HU2KLZJU
dn577pQ9PIIaVyNGO3ixeJHJX9F9WqBsky1v30kE2t89+IOI9cEjF7FDajXJ6nRz
qTsC8BDe0BF5M8BgILYo5tJBvmdMsteN3E85HnjhHBPxjUqROMTPCwxDHez3vX+l
GKV8GGH0noyBUXnQauLSCcT6MuTbEA2ysE9OxWpb0sp1/IBbhtLMbsOKCP7nuXbG
/my4qkZrfVIYX1kUcvPHPvvLNE4FFc2iVw1gXp/g/GE9/nL3EHO7bhMMahQ1mTYA
amEzld3xuVlWD5Jag3TyOohco3DiRKOGM4KkM5g0n219loWZ76uioDSZSROWuSli
TqJf3zYMtUppTYhDamYwKwllwKw1N+xA3pJWoTbphOKQog4tpoKGueRuUIOvQgJr
prVKN/lXcDbDyUSD3ROtFbucYcUYMpfsrpT9axpz8eQqTm7sOcXl6hCb7HC/MqLS
/Gdd98NBo+RWCo59fJN4uAYg9MbWkiWEyxJEx+nb/+/0l9O3UbuV6E5qZrZfCX2O
sDt35laD1CpnZdpMEcsElZXg8C4eQ9Y+dSr0Z3Mpidjx+e/DXecNmpupof4iAPdl
yiDrKTamr9FQlBV38a8W72diSQJYQwO9LcYwJLzOqkBkYwixhHufGA6QZb93LuQA
CFJ3pm6lfi7qskAX39ZqfoZCH7ampaPGl+1UdQ0VWk7w9rf2rTAFEDvrM5U8Ua6a
/YDUwkJyYHdcT7uDYg2WoOTtBVI3SS+/za+AbZx6t54a7zsDhPngzGnW4cx20CAg
nnJ+/63yH3+MXBkWtpmfOmJjMS0Iqi817kfq0BCEJPORlUu3D2EL5i4r9P+KhH2X
MpqYL6roq6+DG5rnbkK0S9brol7vyov04hUlIk3KVlFRBE05kavCm2VlL4KL1b8C
PI8/Q6vq5n9ANLiixtbRmlSt0zxRe6acsJoesQJ5gTDYLb7GE0ZNMVFcxymdCcwf
QVP1p4ikN+R1a4yuTmt2mQEjQx18je28vjaDQJhwu0p6TvTro/8985hMb8qWR1U1
+zoM0CHuzU4dnC7dA73Cshhk95XPJWG5tHUbuoWNfpQPAWu3KcOLmz17k7GbpVDl
ve+M/d9/F8lYQ+HfzJmV3qQkh6ujeifjeptCxxOIHpNplEWF54IJwp/h9kyowL1b
65iGuodLPh2ZX0RNXHxG2lpBJ4UCPlcsKMNwwqhS51Kh61DyjnqA/eoPG++aweeD
CGb6SrIelJVMtoqezhUF2ZnhFUeaRMa5WYM9WdIzybwyNCOTGjb4sFEfOByKtN1b
mpR+ZB+SHV01qzDZ6X1NtGL6pP654wLGhtXiqiG7H9CawmCsd6f2lG21FnC6LaWA
trCedFdckR3cHOTUkh27SyVQk5yh5s9xuWL/U0L0wEvRJi7VksnbT/9biPi0s4iS
qI/nYoRffKUB9XO2G6V8o1kIEBnRxOiIK3mXesuiNXvsRkWHMmSujcl54BSusUTc
OorRg+WhFZAyIugAGc0nVIk+o/BxSdrlOTfvFMNk24K+mDZuhrf6fU/UPNA5j8qQ
KLbO5KRtzGp7uLH6IHNzaWLT8gdIMz8KN6XsW9h1dAg5vwkXzcpBpzS/vyylD2JZ
8utzf/yun3d5xzos2MHgDDi0xREX0AGwgWWgo0yilEfa4dlYpBBNZm90hBDpFJQ/
BBPFm9r3IMra+lFuTaQ5p7l8M1pOHuQPktTZyE3WtCIIHGNwsMIJ4XByOZBqVrhq
knw3JY3gcgff0mEITzDlxafePpPQf59oxxlWKaFVfbvLu5EucIsmwXpAuSpm4aJ/
ICq9gJ1OeZWq/fzGba9aNjEQAGhnyMomPY6ih5whxXThDG0ygdS5nhV/yDoAJbKk
Z6Udsvak6DRgLKmAE6/Na5EJu6sDW+C1oCWGtf5LDr/ve7plMaTf8CHlpaFttzpO
KNn1m+Xk3P1b3iwMypKA93722DQuJDWo6ZG0Q1FqiFfofHnL5s3w2DPX+k7FpLt4
d7SyLHCuvrLVQj2YPWf+1B5tkknsjRpzUEmGayiMH7Qr935CH3k1No8YR1kr5gj1
LE34akeIoqTS8ptWuZ9IDmHXjcayqUH3YUvI3e2gAL6gPNDD42exd+KizAHBcFbd
MVqGS6JRsSrvYPdHhD7SxbMsi7Uj45n25EUBqf8RvGzdEm3xJCVuQQeyV5vNm5Pt
3E+TP4z6SrE6+WUQBBigfFFEqbFhs7ehIFXC76Pq3z3b/7GZMaDH1r018BbAAS2I
L0YmR6ffXYeWZFCF48vxG3mhgQKE4iwn3Sy2QlEHpNymKKEtb/LfsHEARRuq/KmT
a448Lhl1lNCNcTgJQZpTi1Bx+etcYbgoIdxmNy0QBD0DyOyB7svAVXBpk39zHrvA
u+Rz3ZJmd7lqSn+3ut0wmSjYQJdOu3wWFAIuGODba+KhtM1IzpSivh2iwRFWlDCk
iOhMaUhr07XAaykUGpSPa9OA6ZuE45q3EQEFE0JHcZhmC9YEkqd8rhfSSSrjLc+6
5XJ6uylqryEPNnzte5Jkkx/6HmyM8ePbHMuyD6vIaIBEPdTDx37VnkhpFzbUSP6y
1E+MCbnhWW+Aq4kXgh6z7mvDmhmn8t6JgyFMlELShJpL8ACVGEeVraEHHQ4RUBGe
XGbIech307Ne78+2SkBhF2LDUOaPDRgvj37PP1ef300fOqCbvkVN0gaJADtgZR5t
Xza4EFtCU5ODNUrbHJyGyVGjaIo1DkwDYq+a4OOWsoGLEf+sYjcxuQDgObbb8D7h
8NYRUjxYHbjm+9xgrzUp7vekVPBh4hGuazKQWA/ME88qfj1Moe/rJeMOx/KXt4X6
W1oY1HMqZ43gxNJndheQJSMi5iiARlgPtJZrUEXVpoZj4lurXKc9OLzc1vPrd/Cd
cJE6WGSi5dMSs6D8feMny4e1UvysDt0r6+2kBwVvE5dnhmXT0HwB/7G5H0XSMS65
dvsXM2KlTaGcuvZdVXqjNl3Bjm/yyC1y/YaM7cgxW8d6RC6Y7bMzgac7+gE0JZaD
RqXR0VuhFpLIWX/4VQtHKzuuR8BC3paMjf/TfJT3DKwPXkks31xx1ZndDc5ApU7m
KNhjPU+x7TS1gB5XFHY3Tvv1MCKRO9RRuY5JQhwEmC0SDkqweXFe+3xCJ0Uo7AgP
G/k9R5XOO2TVI+lEdZl12xHE8pXLn1jcljZH+PoYuctKEbW6gxzEPbjSZ5H2T4BX
bHwC1DCwZXwfoMMJ0pnP5Lu5GjLFeXGVJaCoYBAhSWr64MIDL0xG3Yd8gAOn/3nW
7iUbKXAND/H7pOwBoaaFQglOknct/5dReNUj8DNvTdteUNZvaBrJGVQxqainHsw0
6YOJGMROV7TdE8G7oqTUOIgWR3Z6Nfn2KXnMUSwiYJ68nQWuCiLJsXxqPe6Or2ow
Mkpe1XWBTJW+6XYs2w8r6T3oInLEydH4e49bUdXFX3zVkDWA8UsYMRdFRM/9iPS3
4RKFFj0gCY4wkXJbYwgNy8tbZUSovtMiCxzfjO2MbqrqpfO5pu9mtzcIteMmUzTY
7LaNZpez5ZF8p6ANmYWbe8PF8uCfGGy4nUDI3x0ZYZjLRtzu1IMHDKoWb+GeVXx5
03M2mjKHaTdxJhPgGj4EfUObcsvUrR2S9mW63HfF+m9GB8QcC5zv1TLbI4VcOTrO
8b+F57bn8V3zJYPHku+gvAOXAN9mogU/WynxU6lBBYDz9LqfdYqL/vztHeDcdfAd
sX078+9BWgkPQ7hNsMQ3YmrvPnjXwP59wezaExUK3h61UNDA0ThkEC1XNnNjcgjW
KWKgG+SRlDzBLq6ZnbeGvbiU8V0xF3dzmXdYroKwHxDXCoJXAtjc12Eb1XdDscEc
PK57KaRzN2GjxuroxGDvI+ddkhmQRcu89RRtruQAwAo1M6/WHjx+mYswqRJkOyXl
F6AGzPT6hrABHpcJyG5tLaC5Rc7Os1yf4B0nRHd+O0Pxecm+mojpws8Dt4JW5HdJ
osMAZBMi9STAb4lpyWLAqoXQjhtiGFcWojGqjHzGuE9s0JFzmlxJgaDaGUKh2sz/
cw5pBjl4IMc5LCPmQ6tt0qyia8lXbT4mkTI9BBrhaUN3eDlevb8V0j8wLJLLKFaU
wcjlLr5GDHC5HBGlA3Q1T3E3URrizud6DyggQfz3Fyl/qUv2pr2SBL3UHiL3zgFp
0s8/RRpbD4/CTiT9mvrnFfm9HrPt1Mgpndc9am05YQak6YJwNH1Hp9Fu5feDEtU2
mddJ+bgXJdU8XQWsY/LWosozol3KmQ4b3dcGe1K3S4fzOjxWu/XhOVCgRPTxO6Fm
quM2uzGYsqFXvvonBsbuyGciPrPQE8X8+X9Lx9Moyq4VzcNs9l/d6yA0md+q/gij
6JyHw+LAHhv9W/5hcB3oDB1ANp30ZLotB+wTmD+2ubiwuI5hEM4w5kndpBHEoexG
6YjP6SsFHbvqC5mFgTPh7zDMORTFukeQOjie6uP2f9d5MvIpajwh/chge6cSo3QJ
JsT/R8sZfUNdLAsbDRXiHKkH6/51AZ1wUswRvNTaArx+cJjKm5jdxOT5i57RhQCF
ZfGUAR3/ABSdGtsCfW+DhscDDEw07biee2MfVRCsGGCGnTw3zad+75iFkXwqSFo1
/7AmQhiVMdiYIrsd7a/Gqx/YEigA/FCdAG14mdyxTXGp3QdqgTGK8ugTgH0EktNg
glpYhHNDjZVH35NPnobEWd7WC4PQSKGNhZnqkcDVse+50IKxH5phvCzfpaYQggmk
2+4LLGei4FOX3203wvHBJQQVT0qajuQLChzIvIEPbgm3g/E+3VRDlNmabI90rmCo
JAjx3yFhlv4CfO4xelewOCFwya11FR58CxpBRtzd+qpMv/ebZaYVUmDN+P+Bwpsu
GyDuiY0M3heDA4sCKvQDaATiAeVB4LZyubo1VQBHhU6YDi6A11ZYjAXduXxwNnsg
+ymkJ/PHqKHvZNErgUFEduFIuA9OWECp7udclp0JOb0tR4YB15WybcZ9JCjnMrA1
HLCJ1YK5cj6n/g+aGB8GHAAg03gbQZc9BYy8pHTB1eqRQE3BOGMg0DR3CbOKxE1d
tTvTQSuKbHfOtdNNIGN5EajWqwjPscrwZfRuOMXv4Ai2OwCCNqOb6fFbszpaQT88
xhn0uAhIdZd9LodD9Mp/homCYbR6wkiD8qYAzjq8LK65fC5NSyw3HvLnEVKJpndQ
ABS0paN885HtaWvTgwrPOHNXKBfmmzhy6PPa8nBJV3KFi+dBZqGBlL1QBtKKfgkR
YG+jTkVSPY4Z+ERPjzigKzu8s999VJWpSxYEPazpBPp2LP0dd3tFbkoakWrUYp/P
TqmhjwW5yK90Ga1uvHWp39E3cswCEtqLswVO/aA2XMOM2+jITSzQBxiRnuR+Vbiy
WGMZcuHRpl5AahW1xJcbrGJhwmFp4M2cDMXds5myD9ASHBqqFvnXxaBePFo01eRX
0o93ick+vwXg/Jc+CKQQihGVoWs/+lPCyc4gjF/WH2gHq7F0fiWDPclHnNV2050n
2dec3gy36T9QG4TFkc+xoYZaaXQeJ5EtIcw2Fr8GNtxtjwaWCJhdD6f7BEHJ2nId
xi7s3vZ30H0ov8w93EzDi+rKtqRoQ2ekWRG5BlhUGkpGMdTBV8x+gn03yHeFwNUc
2rIrMUxNvc56zI20n4jI8lVsHD5L9N1q0QsbD6roIZpfl6rnFpkhW5aZZyD3sPQz
c67WEWx2f32BVVXuZK++IG9jsxIvN7RkeS0p0H4CuN+Oy3IBcbpLOhdLoYOQdoXP
f7ziXei42hDUw52h1zLutHHwWGhCvEhtGP3MimTLnJOLLhD3vBBHvh4UI0dxqGjY
SgjEwh869cS3PMWimzWFlnpMAnG9PdSg5OsuaP6jJqobWaSh2fAQPeChKTdfG/IM
ljQzGuHLrx9K6GZDpOJRYbt5tGCTP15d7RNFXLO0cf7OZkscQajmebnfT7FyONV6
S+181WRUO3+JdI3hRzaT6/IZ7NJ5BUjtBqP6Bbic4ubznyUnBHfl/WiNCTwyiT4V
3zk8wzS9Zcri0SRvmnODwVXh3hy6xLLlBdVQ2tThY7cRWtN7ggt+sKb0vIb7NNsR
OyUJHI4xEuB6PZLCl1FWhjERuCKcI+X8Z3+lz3NI3pXcrWdiY9gxrKVLG5q6F9/l
aHelfsAASQwOPoJ2IP3Ty2ofqi9+MVfZ3eb+ckMLOiyVPv1aNzjdw/vZ5riS5C2v
ewhrvdXGw25U5LIL2ouZmxBiNa5/JN1WZYgz7N7fGJaGG+TTP4Qgao/bedT1WR6q
6lZQNwGRi48CGdl46DZAjARaFEOauopoDsf1Mwm8ATSfOYdBTHYwZ84Ba8cxdREZ
5XqKGICVvi1sUF4q0xT+Ouh8yRlYdrMxAicEZK7XBaVPLWUp5opEgZLPn28zbNDo
2qubCHBHtR8klFvhA3Q/GCEa5Ir+0NGRcimOo++vP9mvZ9ZkHxNZ/7+CTvCbI2cd
0yh7coTUfmaA0CqUsOqgl4fw/gpru5Qgpl8s6lNlJg1TyC/tUmSSAgNcn3zut/WE
8hwE3mvnjrshj+uM5O3qenLQulFNLW+Hq+uXrE3DPYWU/JWxotJSIK57yUmM0gj3
kmQA7Aa/nTwp2BAeE81bBgqNp0P/XCwfres+xOI7mbJ0QpJkC4I46rxQowvqgvc6
hk3bI6Y9YJFOBFz5EoX2hdSqNGZxGuu/ZmxDaCEp/Q4Ei8ppFUD8/1KvRHWNjDvD
rbQG4JsQspPHJVeQlu9J0XLH+vU+hYz5dDxf037RQ5REdtFEPPbp8n2Y03T/NUec
jEe/hhwJj6VT2wIdUjtIi7v9n7wh25qoH3SGr4o57Q5rarOGy0q5kLR6iDPojN6g
ulDo/LHh1TAQlQC1o0mF9BqxUN1x/TUz0Cpbdzlrj4nanhycsT7QXCzigCky3+YA
GRtBEweFP0daBvset5USG4CGqBt2SuvlFggjzC2re9Ymg+N7HActwznJPSXeP5GD
x0V/XwKTO4V6/mXWCWSMdf/fvOfjiuJo8Ai3cLCH6HjbLhEaNw8Pl1G2VfsFz9Ri
sU5O0pNxAoEhTADqCTfWNiJ5rSn5b9Dg84ZyR6K6/jsGH9u8YsFfBZh96SJ00vQw
rd5LiumB3akTe8r+F/eTcG7XcVPms2VkC3IwMNWzvmqPA/vnAtmHoqNP1oUCGAsq
mJY0t9tsiOI3/itnCaLMoTaj6UydRj9bYdqDG9/V1fp5nDpq4Fxhg6Xm5OedMcvR
i2aA4ZpeYftYM3rmy1FeXnq/6QcZ8f63G8vZKqTOJPpK9WbDR2X4+Uj9edP+2FQi
SGFWti6MiYwLSORbtPQ/SEZDt1kQfKPA6VCPwVRzB2ibyv9i7j4RoVJoevn3YyfB
0I5vYFKDf5cIASIauuoHyyjkYBD4LL/HkUGUHpTyNEsFWLZJByXgbf6MLZNrUSrK
t5yRrbntaGFtdmUU/XXwPq2bMc16q+asNtJAABo2qFthvy8CVlC0nzmtl63yDgSF
eDbKW4+E+5un3omfZhh9VzDnD6DYwqXDZrUcjgGW0nDtpf+o1AqjbOHAJblrcuuM
bAkVyD9Kag91D9hpncN3wMxuhdBd9K9Se1QvPuvvHrMGznbHtXgN6c8iuL6MkK5E
pBrxkKTQ9VIcU+1cfYCm/6PqYaXy03xpbIBNipdeMNWetjsFHV7tvUjand26EnmP
9s6FTP5GW75cdoM7WuSyqVeipKgQIlGXD4WpA5dQ1vHXR+OKHY4NGBJofIduR9q0
j4ZneL7oKst8qHoh+Zgh5qDjp/7oaNphcEreOwloxqWJyOId3XRZYWzu+Wq24CKZ
41CAo5e/20cvv8uIYpdaWJk4+Sa0qfaU76u0exjb5pR64hN4iEotGSlFKjp+/tUO
zse0qi8Ucox1SM+6u38rCaAZQ1MqqCtMO3CooTPBCxMQDewRWy0rOZGwy2KB2AjH
Z4d3iw/xJV7eVMUrhIXrxvZw5kDUbGfLk+QWE+I7FfvAR/xTqAfFzA5ww1uIzy54
Xr2NwClACuBUvmMDgSFdT0tyb1PYsbGUO62AQLSSLGvkR9Ld95dyV+jKRs1flt4R
1b6VrDt/MhKf2Q+dQ2noT/gBv/xg0F+OsrUcfR1DsCiTWnNdj4bP2oBWHc+wjXff
lddstVFNB6/rp7HnMgFaqrET10R0Xs4u4RGC4DiNjw7G7NQN8o37dtVXLPDpdcHA
ABP88BV3OHBTwecTC/dC2eYRmjTD7sC74eynSP/wJG/j98WfZvq8fHYFIsYM9Yt5
jFmSex/DH4QnYIzL2vNJhY2Xd7/pXx3B1vAFV6Dm2c/Oq9VRht1D2acoVW4exrMK
gKOHb0RjF1Pl9eQsc/EdsQR9fpqZ/P4YB4/qJcqh7Z5WjG3YvodgeGEky3giDSfC
vcmZyDgDAYjLsi2BlE3BMrvj0O/jHVCAPQFFmOcleSx+p/YvMctpt33R3vHPFIN3
LQP1+R4hWfSVvYJ3jmIR/ANKRhkgTeyWcZITBpffUmd/YmhuOk5g4mDjszOKRPnX
oTNny5mbDWKsFT5jjMfNKc9IZX55cNOp2yZDL4CiRGbL6qvKId+6QvJS47e9Vogc
rdkdkGQkbBTlCQozGRKJCj/vk9gXmOf2IYoY3hUiSITfMZewj13Yxk6UGqViG3oy
ihpVt1XadK6xWBWiJWgU+shGkLTqD3eIwmAIfVFlw0FEGxGg9AdbkoGvGanpsWpU
80D+cs/ofEolkIiifxFSbqzB0ZUS11SSFrJ37hr48F3x0ezGejfCkFgSzwvdBswj
LtFHscrkjdBViz31JpCsa7YFwaQPcqI7gvUs+nRx+FjCTpdCuQQ2ddgQaR44ZvIZ
u/cTuSUFnNQt+UA5ojfRog93wVn/4U9Xtdm/x6I9GvnO51KnnA1aDJan9WCFQ9m2
qm+6VerpJfGLOCCaB+8T/2mzkl85X27/NcGbkoH+UqbMgJN7yLgZ+s1OTywbHT2x
9NQkHRPxK57mr17gVIxWf7OsTP8qNKsJgKXGRZbQPPG8hQnzHyqhbXFb7KxqrJOY
Y3j0/NWOP0M5719otisY5TH8M9oAOyP8okB87Q67bDQV+02GsAFDSq8TIxJv2vPG
ixfjUKFQJ9ejyofGPH13ghCzubETmaycH12TPzZyT8IbE14tKzdgPTCBr70l0nvA
ocFvlo1qXWgmHPbumBg4ZBkHXWuFuBHetMDEEHqVZKcplIfmrgs+49YnHP4eHZzW
E2fZRC4ZWpckatDJ42jrHVtQW77AO6dFHWqpwlfkq8zDxAx0fvte36QDByjbXbpV
WU4UdiVJwzth+/FkUNFT+50dfgNtauWFCI3+sEjxTRa68/yZ0z5+i+6FOe9nP+cL
tOOcHTrp84sY0gO7cEHhqVM2CoqIqAkqgzWsB9Ce6g2XbdNiB2IzKdgp6QALgr07
P4NMAC0B5Z6Lpv1twyt5wqLJNMugRURVI1GOKkFtgEIeVbpPZfXfqVXmr1YjrEj9
d2q9WelQ1ar/WUKtGHWbMmwl72sZDXq8noaDwweq2Mp5N6ocsb1np3Fr/hTYGCRN
XJD69nYIcCcwLhi8HdLkkjEFvNxrzQMQ/tmZYQ5l7AJp5TfmbLFMlRh/33jQlJiT
apgKYIEPzQ7MsxjrpxlfiV/uQ/Xfd/ARWNNen7szX/VHcDUcDUNVcaDL0D+xBM2T
y8nY7jCxfHLkP7AmXTYiEob8/3OTTpXfi++82uHKyLvA0CPp0HknbyvXOCQsbMJw
akkkR8ZaB2VG9EuwRAUbYR7k/cQXFHeVktg65gUK4Lpe9OSmjf4bpvZ+RHI91s0g
i9F8H4vCIVVkEjWERhQvUzRBy8aH3m3mKw36eGuiSxYO5HC+IsR1/9Yraeek0Y/2
I2YfSr8lpcwVrxDLhOvnowaL+61xY6uud7cB7EuSmI6t3VAtQlR1ihh6EUsWDpN+
GP+GkNRxDcgst3BSklTNH+AS6PCOG3JmbMlyE9B3l987ukH/GvEpCKp7019UCdFJ
8zH5aNVqsHrg4TQ6+GL3l/gMcAaWtdGNAzmTj+lmgChJEtb5M4yDi+WJyKQJN0K1
AcyWrH4sqDpbeBVD5UY/xZkjs6q9P463KX3GbqZtM0wpIcSS4j97F7p7gB9eQyWu
iZWhEv3X+ejzzclPPyUyTWpSeSG5e7kLP6BsPp7MQ5c4nVs+9lFU8CBwtLfegq1P
I8wnp6it7PpCYn1hQAZfg7Z083TcUR0PucZRXF0PKHiUeuu5cpoq6KPCRRT6UtwM
WyTCf+czXqaSOZL9pk2v2xohDmTxQ3Gvgi4z1k2rDa6C5qpdPQnG5UYnPsa5wLAh
r64kJOEEih0stbTDDXelWOtU6s+h2DqQ2S02NSCa3poE/Fbdya9bA18QKkIvsJQ1
wdYtcuF+FmwtQfMQYJCYKhBF6L8nyRf/XEdy2j13CipwPWuMWz6eHFnRx6glJAad
JQI09CUUeAbVM+jSOZnFiHGTBAxJFS/sA+wZYkXntSpRwNPcfDBitsH9jNJmisvG
fx7ioebo8hb8ewRwQ9IbmQtaWEL+xQoQBaVVg+uHuUT59qJwvONTHw+vBwAb5lvr
r4zEKnorC1dUEy8k51Dx5en0InVaw/8S2EbS/h+93Z2XYvQWWYJUYgII/JRIUkk1
cRmdv/MMFur5SgtZS+bZ0K4BjZDJWWKuqjy8Gk2qeWpiRVZolYUkITbO7KabUXdl
Ud9JPdMSHGBm+3h3N3E0Z8aLo1pKUKEJOCc0nv401bH/ZleIVCPdgVcU8I6miVAp
k+tlwxYJUSEqUa1MweM0gJoTjOfc85qGsf76F8cXDiXZOCspJwsZ+TX0Qo6eWT0k
umXrP3BSUNmVBXCRt6wYjhdc+DdEpQFavlNPf4XYHUDCpksyAyedar36zLcocSfN
MLgAOTbaPc662zNqjuZq0jWVWM3U/sPxZibtKoUWoWMg23ABOeeVd32XCfOmBaiy
5JxTwkXMqvXst2X2fnL0J8SLTElm8kFzNlV9oeHRrp5fAXqiNO+Ia7qu7lXKVy6X
StxD1rc7ylk/xv03EjZ9vkcIBS703daxfhcZ+7ND05vpX5fkXkM3arFY9ZQ5S/P9
rIC5bO/kVNMLAolG9EVCgWyz5KQJsLcJj2XWCE8lW0TdP7oR4/8xSrWZ4A8lEa7s
Ut/Ht4SfuZF4uWgSkbYlD2zeY++B7YUOWnRE7/XY+2Yky5LvAd9YQ0Ir29IdEPB1
6Dz7XqX5BlsTQw+GwYrVpfDthywmpfSoh2z8uQPyZpaME0fNVwWYueR5ywOiAOJa
fbslNm+92KroAfH3LawLNk8V67SqTWTRa4mqVOpPBMw1Ge1d333WEHWNUOwQKJYE
hpFffGOROZL5rXyiSHKR1WJnl7zBvZdzbdU8thT8TGS+YTARPDnjQhh8rSOsVErl
cii8wBtnGkpZaFAkOMPcZg2d0/LTYs0BbnSW4cGPq4TB+xIXwfcNEIHYSI3rGj6W
KyER/vmseXJzMd0eG1aiT94/mPWF3wtkPru2nYZOQIgBaYue9XsDDszTSTRNWVQy
yGgTQrMpVxsLdbHB1PElFTgc5H+jNm5QJyMCkFRV6ba4LNeddt0qgAQlK52pJjIk
gCQjy+f/1mhOi/GwP0OH50l0ZKR1cHuHlXZia+0w+0B6SDqqr6MXym4PvT5AnKgq
7auB9/rMU5mvPnkCrnlCXVnl/IDuudxwuo3oTOuuHCM1kfAEqJdOEohGLCBYxmtX
a9vbPcrksXoMU1+CL5t+BixJTF1n1sxby87iYiNIxpBGfEDqtfhxNa9U+PpZXmMm
Et9UJkm06dlg2o8CWPvOisaFzWeCp0HsDqzXNDL3/TboYiPoG1ZABThplUlldWBK
rK1t0zbhtEYgKivBZge/b/FBt1AxGxvNxaA++UpoMUUuTjAFkLFOZ2nSqaPjaJfu
MelaDuU3i/tLBfLlDSzpqVfAYH9Gq20xc5JaSmMRqrjo70Ilc8xBfd67AcOYO4wm
RkmA1btlL4j3M4ZxU9nknwAnEoq6TjS+10WZvScSB6CHQf9t0/VMmPMty94My3St
XpGHyCx532gFBHKp4jqGOkWlw0r4i3LF/vS0WudtBl2JddBDoN8Q60HlUd1CXrdO
qXZ05AGCDaimXr8U+rSxvTVrugBfYH/6dsfgHKtxaijVMXbVVP/hWOqXHXEEkIXI
QXkMHVUDmNRxiNyHWFgG/v5F6shQUxPBid6DI12Fp/vT/2YffhiEM2JBEeMMEjpN
nSJWC8OfEbpd5Y2bOmBGw7TKXXdRSKu+k65+oyQZQAcEoJD4canrmjNhnjkPqDYo
hensq2NUEKnPZivL9VjYD9CYIehEXCdtH7x3UFMKqBJcjcnfVD/N1ygR2TiPZ7Qp
gPdNumVSRNtVH9hpRUbvex+m/+tqXaBcvaMxEOYcl8EFcn74WnGslpaE5G/dy907
mdvloRn6eZAiEZpRuDS8LPfRj9oTi1l0kmRXtsoS/cvAayAURH+XeE1NWBd9PyYz
n+kvm+yAahyi8doRVDFuU/rY9m3CDzZ+mh99NmK2kXQuaaCMI/QBk/TAiEvknRU8
oWukk/mNiEzM3BRjJPm97esfm4DFrIxNvTJCjap6f9fOneDvQD4XKWf3XWxhB2OJ
3lwAkr/DCGB+uhwbK+vSaFQo+e/MYuSvcZM/oJnpfxch23pFNwobmYPnk+yFJNVS
c+IPoGVRxhm6wVhRdrzsKIu0UUSPOTCou5QEpTu3gRJm2n3658GL9hddepNLOBw+
e/CQTSbwrhCIarfezgcB8oRMdZX4zdXWpuHTj7DQ5KrbLPOQ+gmHj7b56tSj/q+5
HEURRY4fOTeTdqaajJ6HRag2/Nh+SSG534fwei4ChV72GuYYONU9PoHxWnVq5L3I
jDnpf2oMetuT1B+lTXIAYgoNF8CGwqwAtJRQaWRp754jp80etWUe3vjSf/0Ihu+s
DEh38cDsBBhAqathyfSN2IHIUeyGXALV0hvLW2dEXy7P1rxboWgCbM0T2oknD3fC
c9jZhUQbYFsCYWgGaZ37I/DQMqDczhMa0NsOa/JdE1MasEPcJE/Y2xYkTIBXbhuV
wQQX00ilC2xB9PdK6SPsN59Iz4qIkMK0LvGr7mz1Ke88BNZy4JKGryu/qasBkAAX
xZJbwYJN1mvQde4Zj+L7Od+0dRs1XA+6YDbQUUBMtkY0YNiMGHYugjA57zlpXoTa
QUMULiuRmf+QWlosyDmwsA5i7+rNb113P2WCbcX+QNjpMvy2pXRKE39qwalzs+Pd
+J27+XuC8sd84qKDYxDdi2Mi+0YkeQN0Q1e92eTAjIU1Xcow9bxzsXAb1jEv/Wo1
U50yoFSW/kfCnK+uXQR9yboJEzG0CcaCA0Q/6srNCUDU8H0N+o3n2dKxiQp7D2DH
W0z1GWwbZc0Xi00VIXD0UKZeJGFFCLd3Ke8aNu1QMmM9bSlKKpSRZw2WANCyzxP7
iENuGsYjV30DQDRinBip1gtzRYc+jmjXJ6uLSQLEV83D5OhjBJjUy8uDgKDRwfwW
zKNCHh3eWseB8BH/1U5zkA47itE8zULJzvYuXPgzwI/wbaDjp9wIChC+w8U8AAsI
/J3lTHv26okTCafxXksfVCuaWB5b9hmOEe609j88SyzgQPxzdUiJHi33AjOOzB6I
BUBLzceupEgknRdN93f7Cd8DEShcCrrvv5v28MS+A6+8HzbyECmnJjDexOduv3OH
QzxtewNSwG90HOFvLLlLf7/+Kw7AckVIjmq/Mdvgp47MDdI9Lh1RfCXJ6UdUfB9J
ghsQqqGu19GBA+P60MvevRZkc5qTDSgQcgIDqJsrNii/D6jVrYO9oI/8dyh9MC+T
Tqq0k4ZfqkvCjEHPTpq92VPW9UcSKhP1eI2oRWyydR4ST2kJQ7NPUPBc7eZLnI0m
kqn7fqEnklEBcb6KIVkBvci537ItkO87zlxJ6oOspRlZ04z03usJYKc6aa4bMbXh
IJ8AlaBThzoKOdMbfTOAjztsMFFV8NR3vpmTUyAxSubaBX8lE5UlDOIwLDMHODBy
kkusER+WztF3g2M2KuMDAaKAsczawUAGMl1Z5PgseoGwvU05/qx3I6UTCPNq9QXU
xrFaNessdJuLX2WYmsd8vbZh+Uqiu6YXmlVDbYXrZUbq6C7wXdvbRnNAn8byw0JF
8TCGZTim9o2TcWvCvQ9G9qVTjoRSNpm5Bb9RBfhuQTvswXSHANg+DpIVveXS58DN
Eqbw98YHOFGnvRlWhjvL2hBtMX66f5DGv5jMke5rikWVwaJoEvlLLUTPEssJw9ji
19JWGFzdDGRycuwfdANn6ZYjRtg+SZadqaEv66970Y/oAhTR7x4HhdrUzowQvYgw
VlpLhgFDeyeehPL3VZPeCukpJsh2gZ6Z5AF3QNwnhWf7hozC4hKp8Kk5nrKG5z8G
2m1kS7s/PvOCB4/VAcNnLdJdeJGjHiHC4vomiSyFLMIreH/dHGM8qWDTpE8NJHT2
whb5TKpZ/aXrqFs+qFd+SkW71/J7uK+bodZ/myd/jmaRyP1GZEVb4Eyp1jqdczdi
WtjLT/hYeeWOdLUIk/dODbtFh1eajX8KR7I0BTrLPsuAIjwS8wSDXUqjaaz1/GMX
euroneYVzbFnaKNS2IB2w2QC78l8GqZhD5UVzCxj0ZABymaL8nHCZvsgHI8GyRhV
7ytawHYuX8eFsJf+zgwmESRjQFHjy4RLtwADOOhjSR+Cy6EBwL8vTuzmLvuqy3NB
4jkHPLaEW0Sp7I9GDC+lrrlqIjpyvo2dEuLY55wAjLAy52g8nfvwZ2hoX6YFuGub
Dse7pyJ2/a5kuSXwgvXSwbBXpGhdx2ax9Yug1LtN3PJM44mCwGCf3UgYvtVuNu2Y
02+pTelASOQ5+xQoi4G5RH++M9iYJ5u4Ec1sR4mZhUy+opYAW2qtBwdy6h1uoZkN
nYiXAcOumy7kdFMOuuEjsnd0IowsSM26j6mHuunPaH9TDyhtcpsjXo8/1scltd3K
IAE4CmsNtqnvoNR6PU1DE9lVqTS9RBHpi0L5YIqz3xzS8L74J2zWcd95nLMlu52M
L4ucjQhYFE+S+vJZuhQCXqA9ApWTvoy88B8vcM8JIuHmXrFL0/632BoHWhq7t6w1
/4aIxbBfmDVMq94Farj0nzjce4vx+xgrRPcBc3vgNoQbxDy68+Rqf9JnNATaAJSN
rCeOS0/bOcFlAq470sNhxMTEGBqLyURsH4HDxuKkajKVYPaHZtR9aogGZCtQmvwJ
cd2g9hwSvydc0bs+AhygP7+2KN51wbTT5RpDy4kSTcqtmAfzE1ZzPpiaiKEu43QU
Dg/CZmXoJzO60turGRLJ4TkdOA6YdToPnt/aJdP50+4AV2UwgKDjOL75UDg+/E9W
xBVrRemcg3wlsotbFkj8oUiutpAJC5yNzLGr3wiM0sIDzw7LVIEKfRFKQf878ulH
/u3wm0gOP5DgNnjh3Qn/9YoeHOnoxk68+GW5SZIpAgfyBtlU+hwM9q9Wykpg2ENe
GlVMsqzFIbQPA4qWtOQUOPQd7oUWA7mUfBKS9hRIsb2LXonZIxZREudW+0CmLkWD
9yEkubx+2po/QyJLTTXZvqa9UUGy5uklthCwrJ28Oswfi/Hw/WwThrLvH3IPByhs
5TCKMrUJvA3ZhgvyY6yUbSyPTb9ABqrk3e7mrtT3YG+tmtZYru6HNTGiZbV/qwyo
Eu6ybU6+i9Ppgqm/pC37jVPr1cufHbmPEYBovL6jHCRvg1ZgY3DGg/DJWkdIZJ0/
k66s5HM0s2gRaYu8g8Df0n/syNxuexFWseRkpcdT5DLZ2Fy/XjzO/ko94qOFdItP
8lGJqhDQ0pANHog7sos8NeQuC4cyNEO26ZG0mAmQIXjioHhJfkD+5ZgqngkxpWKF
g03uVoNGT+jaxXiBMlcDr3f1eMgFyWuz+Bg67P9AC8kaKbnP5kckWNC2NsN678f+
CyvVr93FKdD9zKbDXaqf6lUNAFLwqtdhQMaWnNTQbpmJBesTXnt5zN2E8P/XWVDx
k5ruBJPOPM4yS8i4EGB91CMj6SM9EwnpTAUx1rJMum8+/iwzTA1740X3p5asq6nH
nVf3AHLrC5opml/aNBiuDs3Juf8Jxd3HKlQQKzk8VJb0ZzDwLKj5fHjbM5edFE0N
/Np0pwUJBC9hJwi3D7uwYmhOi2vU08ruVHKO5Xqy0tGXGpSOJtJwaqa2pD7P7LIp
daQdDsZee7TcfnLGxiVjjIyClVnNi54Z7AwoMjLX9R1w8w31i97W+ILCXE+kvlpg
iWqbXH28fxc7J5WscVftMSMEJMId1Y5gzE67+V3cRiUwEPYYRdIPzvmVjZ5GSrLy
DWmiEIv2yZRPus7nXF93u/eFbMADaniUR5+naF12NjEu10CGm88zJSGg3zw/Vn6B
X3KpZleqGuTad2NRTTgV/n8B8K5C2rIa6lgwRkfT/7JCS8uswETg69btIRQFZWoM
GLtp5nHDEGQFspdsiIUcrO+MDW0UaAlFgKsbFmK0TZtSy1+0SrRcy+K+Bt443Pcr
SM5Xg066X5wTntfXa5U+DQ9fKzlguoDreM4tuISO/w2118OkIColn63RCMl2R4wx
YA2E6kfdEEstkBk85m9H47ihdzsK2W9Axuh13TDqrDwGLdCpDArMqaXLUAnwYNUk
q2cQtyN4AIC6+LB7mStpXQPStSSHNdHR/eXRwqbin5uufbOKGj6f1OJpa9+x3ZFS
LO7pHtopUZzZngJf4r/ChUeAvVND/V4YKJ91/lFOclo/SkSaxlrTe+lIa9uhehqV
PcxLJC/1bdV+VDP6CV11YCxVXI9ECnOr/rM/IMxZGmOXQUTGp8wLErEqh3EVbK3y
zrdaq8BFErgK+5Pam0GXw/dmtV+7Lk4KrJRa9jn0h95iLDfdIKaGtCRqfRqyNNzK
QTWwLnaAbNZm7nIkaK+LcugBAxqY9OShQMMw/dwqjpYLPtuyAzjw7tfrSKDPKJmZ
l13yrokkmgvnNX5cIeObRLnMsZXB9UCymll37t66SKasOQCCXXoRbGAa8HGuLPB5
41wb2JqBjM9YGQZVts94QDvxbXuzGS96ZFYvWXNtAGWgJZ0ozyrwUUIZf3EhbRdf
GbDehO21JvzYbkIPW/OSSsuldLlTf9T2nizuWBwk3si5hwmFGSIp/cOaOAR9q2ro
mhpCDZHQdrGCJzBz+U9CkmE8pvWgMEnw/W8zG0Amqb0e/SQjNvzmm4tUA2Pi21Wl
cCmZkE98HNSjQ+k53lLV6CjBu+YS2SjGGX0NnFplLoSoN1Kv7SSHo8gQT9zaUtb0
dkGo6R5dGRMSG+Onl7/xEoZNdPs834njvkCJhQ7dgoYz0/wFYFkt74KtfEaVBOP3
Px9+IK88sDvSiFqVTYD/wzjW6oQbHKvqkoAtTJppIkp0ISxqbmZd07FatAJ1duyr
nWGq03Ye/9aZHCMXHoSDcJ4PnPFXf9+JaEvE7qOr5ppKDetXnEI+4AgOZM2h7GfW
zNUzgJko3RHnUpJLGyf4pdUa9umMit0qZeH5AWTM3jndlYX290vGh11Fy9oZABsK
30xTUvb/sDa8Q6avOe3cxDStiqQG7wnMfBztfpguQnLFv49ucueuZKR9hJZyAXhW
raPM6utAnObYja3bawx7sCxjOBKrDlGuTawx3Hscr8ujKeO2RAwmwLdVOS0AkB+I
yVfE/FX4n35SiW7BWYWJTGtB/AoUracDqeNTHk5bKvW51Oqlv6RG9k1zk6E3+1YN
UazbISZ9pIS5RzzLWhPGrnpfUulrR6z9hXt+4Q904E0+MwUQ5Fn2RDhXyPlkDe5k
+jR1T9hMOsZ45/77ry8hEKZqM0cOWIWOa6Mlzui2noi1aRtXS8xOzgiwwqCkZo6V
ZKOrDATA3SkY68OHsJRkhbYDOFQy1gJ4v0xbBiVQqsd9OU2I2y/R1GjZjFCpgYR8
fC26EqDUsJFc+66xWgMoFb1kivCT3DJcQuF4HnzK/wOjn/a9V/1FSdWuylFhlpd2
rE+sntEMrnHBNpelKXCgnlAytMs8Ae3EGtMxeBl82Ok9SooNf1HyZ8Flvr6ZXBEJ
vSRrxVw5HrjYw3UgSrUhN7/dID2tQvJxcsuJJK/+KLIkxwCp8Wf/N69NjqEa/TmR
0QNZbW27grXptx+WPeNvocKtwmIHCvhkxyJSeh8mrs99MPEJA9mrdez5TLrOvXXW
4549dYCE4y7k9jK7okpY0xTz7qtUapsRUIF6x5Ea4UcJxMnzn9jVNaD+/Z90sCf/
njayMUpd/COxxCW0KbQSCMcOswLHzcd0HRIrFgWzidOFzJ3pDqWvIh6IukR53vP7
xxPXGmuNh/ffdxMSBM3Ec83nVHC/KzkaF6hyypaJ4dDvOHjsyvTq0qB3UnsVbv93
cuGVF2gt3el2Dto2jtvSnmOV6PWjXx8EKjyOz4FBbWeBdDxz0zl8qCZ0ePtEhudS
8p3O3EyzQoP9Tz0bXK6RluBvkvh8T65KBSYyhNuJg7IMPO4BGVfoC+y6vGnGOlKh
9RtlV0ARCvYfBEbE/1VuD9SzOuDt/bKlG/mG46uncy594FJRDW0bHUPcIhwhGqzd
2eO2JPvI5yEKEsMLsyj7MLCWe8yLedHwH7vPc4cgYMAz2+xsd1ZRPYqBEiJu/n8D
EtN+Jn7/qkrzfHG9SRY5OWqtmdrPEnFeQDvd4HDEfMmOeRIE/TjGZZ9QV7oybqht
sjfkkxWBaRiZSjCRdhIWTfi2QjLJzpLHbI0n8uWH+/VPghu7tKnD6hdMjk88w9B3
bCQTSDwWBl14gc9bVpR0+/aoIzFUh0PcvGaB7XAei1DrSnyUBvwfa40jMEtnTg9K
z+qJGSLI4gHF4P3b/Ca/f2mS21qKBy3razrreiJHBYiL5evJdQxdsJGVVN59aFgH
lmvZsyncVWZ50abMuG82PyH8bAdygc6sp1E7/iHjwIEbmIMGi/YvxKkn8eictjrw
PQHXm5CAwi19BQf1z6cFaUnywlpMD1b/DU6HZAkksCYQ+oTPmhwe2EdJJvJrc2Zo
K/EQmxsdrqbAMEqLijhgjyslKTkFuXDjcz4a1DfxRcEiM2t80gDvXHQEqiH524Wp
FyzWcie3Xl9bYlQLROM1lrA2IaadaWqVnZzyBCsqhSktMiM+cAvL1sxCKF7W9eV0
3xz83EXDOW8uNMg7BpI1WMBBBBpkUhCkRYx8I3dBGpZy9sVqzLCIQllbh7VW43c5
724JfUwtKOON59AlS62YnzFNOPKtRCnsuyIZOIR4TDi46ONXbT53lwGbGKywGUhY
ECuauiZccD6BfAHYoJaZyVYHmJhbBJBdmZtg9fc/+qTtzIRlLND/Vk7T3252o2Iz
n+lyoqXdTlwO44v6lcVsrs/7dyMUbQLfYEkbKnsSpsXaguPj//78v9lajleBte1Q
yFr8+/+OgedJasBHbb5UDWp42x9XuPssnrVtbdyOzCMI8fejEb6gNj3F4yJ/wNPL
y4bAN93FiGI6TKj7KnkAi1B4RpdoBni9S1AmNF5l3Ywj6RgRharPkjMUPPAIFjg5
x/nyTO3/6JDos597vZFR48LKlsiuALgws/PRrvoIsZDocjwQQ8mX+IhC9c4fnQwm
0lszkhHuejHnWTFR4ioHImjIKRVgWaWEnOMwdVsXyHXaFuaQug8RP2Z4AUfBv/KS
iZgQqx2Qss5FfjkKH7HJsymn+JX8Tx+BTjQp4R+8QTPojMeeaN15Si1JZi+rKAsC
RwEBtgJysrBBMFmVJvUU8Do+J4snL/ZVfqfP11RfoCSEKm6PM1wka4IfSQrBPPLj
17bOLhhiZEDN12mQg53m3+LiQzNrorqadBPaKxGC+S7wXyrL8xIkQKykt19UIoyu
CL2e6NXcPOKoIpqLeD2H0gzC3Ig5ft9ektjaTqFsOr+M1UxGXWrhU4jmvZlVP1RN
y97ao9HekWwdM5bOXYh1YLOITv9ev0B2FLDi6c1aulq4VAMkq2s7os0v6tbU05l4
9aE9FItAWxYswiieqft9DjEqcnVh2YeiJ/gvT1JDuQJnq9ZZzZrQM6fScUHAV7dg
fKWIeoUoNSngbTmBo4PAqLVOdZX+L3TBZ95r0dJ0V4EcSst+XW0SobWbLQ1o5pUv
K28OksKPZKsQtygfh+8X5NhA9dgc8a3VHBVVIFEtm+5raonmRtPt0nYtLgsOGSj9
Nvhs37Uyz+KO18gNglb6FTJMMGSJ1M5hZMM+JIt7BJXZSBvVFmOjgSe43KJWHtPv
yfcJCdKAE5oehY2mK3997cf//FNZJJxFQ4nzXmHfVldtVO7p7ArlVCby7i92SY9K
3C6YCO/i3cKE+rsfCy52CsGVYZjPBUHKlMUZ3wGdVAfRR4+YKnwMkH6fYIdWRzov
ThVTBGol0DIhsaEYvVTtA5HZXErQJZ5lOPtIlIuMW8RbQqelDs0yk7emIAiPvAdY
u150L9+oAA3b3F/vK+Ybx6FNuMSyqaHPUk/iT4HdQH2+srQot+cEchr3vd0LIump
V1tmOjJ+hAbtWuVREMxNOfy6yUcYWpsKJ1Ff6R363iCOyrjj5gFSwlfj+eZIec9M
iNAxvCb1W0UFg/QF92wl+SxATGZ14wR+B2N0g0sXL2Tlv3/bFQpOB31ZdGtqaqri
iKY6zhp1wYyAsDV2qg9R0GZMvplXXf3zHV2f6muYFvilEesFdjUK8xzShqkBoQmF
AVJTZcWLFS9tftkq0G49JiV3sfg1kEAD4IwKOZJ3L2wT8H5QsY/odYbjk9Chit7U
dewR4JioWBYE6Syujy2ARwQGuLlPx19fEdkZU7nYAo2mJ0g/XI0mFAFGNmSBmtpD
Ff/olhDrUex8GNGX+98rIWdstXWUkwYkD2nyy0ecsVRnEKA6a5QalilPJ+yvLvA2
SawWz+5cN2f8J2ufCuWD42Gv+FnipxM9PBleBF/ioiEy+HoByisxoZ49ktHH1rOA
+5bzOOc9nn2NKLrUeuJ0bbOrdiLPIQsIpE2+bmQvudkg+Cr0aKB+FgbhV1q9VcrS
5+r8Z1Xl73rB5G5nLUitZYiVI1xp4DA7voKgPlCD5XcfTQ+vFkqFyKiP6DHkC7CJ
UBd8PcjpXwkWIDwsLtojcRuM0rAmdZrBvGaFspOWR5xOsrh336tNri5rqUZv8iP0
fSacxjxcK93+Lf8TJUFel7ZeeCMWWy4dQkiAuGrCcyxk1D22HttgzeEfsF9+41j+
htQtbwGvcMipbzSAxLVMnPlk5xHXnn/H5+aRAHLfKzieGWRWd43WNI6NAUHwJkB6
5hmrwo/Cr5GyprXUI+DjRX0PlQfnb3S/GmGLBc0QmDm8DJl3RBthTq4YXRHG+cge
ixSnv8dlLoCY87rHa9MkVUz/jffGKAkHRociPiNMyRm2R4iKwwWq2Iv8Gdwmal4v
wcVFz7kVQyw8BdZatsYVrSaqtnPhnDZaRA3BFM6tSFHDr6Y30ROed//wDda6Hohu
EnCmMnxi4IMJPBZhOtOYsdt4H4D71i0Qt5HyFiFvxkqHsUVgioEcU0GVyBV2keZL
PimGg15gsHcmR5rImOt0b3UUncxhhR3uT6BAEkwUejwopFryVYQJLNtxcYtzxtEL
DTQxbk8fRMp3yo47ygXV3Sri0KDQSrMD2AM1YKaVQMQa2m40d9mxwtTEvZ4+4dmw
ISfxsWsNY6HKK8S1FUpA31eNFyyonEATMPDlD+tMl9igOjg+ohNKDEjGt3hwciXs
BHfPukDgMIHqL8AhVmk/p7LuB+EvMeYa80YhdSACqsFvWV9P0vbC/57jgp/PCRfx
8c/HU06fO8npVnMslF0BqTF3RzKmLVQd9W3c5xQbMiUQ5AE54S6cryQZweCAFXab
33P9D8pzrf/+h85JurTQvDDDAHwpzAzNEob4Re6nGAVb0m2M9FU04D2RlFXprTJZ
PmKi402Fop3LrHkklt/6YxCKRwucf++hrNbL8ZJ2rI1uyq6Pqglxah+Z7tlnjBPG
C5gWhJyAlBEJHAWLG0AMa05foaWAnAFvfKpYFebOBp6Ib+3zlHLLXmJ9SC0AjH0V
1zY97P8iO8B5yLCMc94SlcJPZjlFQc10fUbmfEfdiAR1d4cjotYAjMauVEFacOFw
3UixJDtiFVqG40zHVjhhRaajLo3r/+G52Rdj/QkukDTBxQN2jWQShkxxMdKSlsgj
JP7JlPkFLawzzXtQ6KB3AvpfdJlaU8ldqLHvKT1Czu3/g9cIMwbDQSyHSa8DT/Rl
qhT0GFFeNGe7N9WDXgyEeweckC8q1/C7BMhguvL9odZSS+kg6AXcPB8iHfvzVJIx
iTSd+yahWDAe3U9znhU4mFRVRRTZ3m2AVVz1ryokUiwdmwY8d+MXP7awctyj2s+H
PxgT69XoHT8WaTvRDfJw0uo+dQozLhvro01OtY08p53FOxhvuupD8uAXpoplMhYn
INKDy3nKiST6ZXdvJJjmYBuoLyCdG7m2JWZfO51E1Y1MVHOMwlu52wVVBT5e0la/
0TUGcZLNoe6DRifhsvYyWNvpqeOblIiY9i2DNKJpO+5NjbB3Se0ie6xebdThCrMG
qpfUySoQ8PMczecrsFZRqgDXV60IhjbPAJfswD1RCjkR3k8NTTZhA+5rJSVUMKEo
Mr1nqwSxoKry2ND3VpoqgEv3RKf5WiPWP+7H07ITm92u3oU8r9Ze10xQgrrvohUs
+84RgGhdsM6fvvEBOdLrUg4FSuIqzPVMjGFhI/D5YusfN1EJAA9rAYNcJLD+XA9Y
PRF4TLotri5zLyxBiptAgFHNOyW1Wn9J40bbk6mB6aDk0JrZshDKvKksD6vuKaK0
h8CA1smnS0bLHX6hPjLrXEV3eUk/ApXOrUU92Rog6vkkGbygWXzfgxCNBf2pK4qF
3cYQpzgK8zwAlQsSnebsYEiO0W8jrqxavC4+JhMOhVcKUGXesEF0v9+zVxnRXV88
RRNfjoDOCs8T43dtmtnQK+3qELclKtMbiLKDdCOK1aq6qcL52u5v4SyTfj4UQneK
x2eoMdKTHZ12kwRKDG4RcG6VXIk1M475xAbiOrPIBatWGdd4j1RXOaJIFeMSzdXC
DtR7+C8TirIfnx1Ry2GrL6BO09fUVJ5OkmAEt2OZn5pKpss3w4ZE7TfGSMsyG7+C
Q5UzRz3KSSzmb7DWTZWFvJvnS8ryuilpzeN6R3Tz53Ltvqau21DvOxionuit1WXx
VKQR8WX5xb8u5vxzXJ8L8qu2q2GP7C+SH+NBCqz+5LCo6QlHSEItdNLajRpuEHim
AXv5VjxMdNCX/VG5JwayZKRF2JRiBF/C5fSqmzd0ytiJpl4gsiKULrSoFAJwD86N
HVH5TOHd6jewi4QyJPy3pQdIGO3DeDlj6Z2DGGtlZEPzON5dvmSUkIq95FKAn+GN
7SmI86x4yRqQ8u9UNKqU1ZHZi8W7O62ZEhK6JfROSdKjvOULu3BIxRoLsXMUOWa6
uZ9PMA6WC4DDHoW64+Ge3HJhHNAM8UjuY8uABsnXObBGAQnyDk9oab/hb3eZ2e0C
R6EbCTmfntXNujNGMj9JPEVIoK0xuzVEk7bzkOR8kA2YnrrAWPt1RErezd+yz5HP
8fpRgCvhWGJOKgNIIM6YZzDi/UceNAVUWR/SxIJu+F14f/p/uOM3h11POC2JWZlY
sgbrJRysCZ2Cu2SeT8h4JvXNCQSbDcvESFq+G/5TNFtLusTLR8DTq5rDIWItN4Fy
0Ei7Wl9McoUJDHM9rctYJAkxcK7H12/2xnkdEkg2m+tl1n1JU0zOQmNU2EhPmWCP
61fPUi2hkvYwgVEeKPVhpnAZDo0tcZ5mO6vBOT/iYnycc/YYc/nE275sO56mKzOU
tsC3hqEbTWj0oQ0JObXS48twmdTHXzfP/Q7RyQfgaYhIcguyr6eKrBCJt79istBs
2yMg3oSY4Q7//RSpMjYqiCnMKeLLTcL7sgsVpug/Wm7Nee6D7xm5QTn4XXRlmcEr
Ez3XLXQuhCoOp8u12N2c2s2mkqsyznYiYPjLpZAo7VtyXyVzHFlrYQ/WJ3uPukG8
6Ep9/hlrLyOhLFXQNG8eyI3RDOqB5veckwcrei7mj/1n3AOPehm2pXrncRtWOZLz
FljEkUBwRr4vz3Gor2gQz2c9PMMZ9ptBWRmQ8M3MnSiE8TLZH2cCDlNIhBC6JYBf
nd/SHBAK96g62Z0l4QRUQyK4PNph4r9PH70SrFT3bW6PQ1NL0sN9fgfA3Gzb67OX
Sj9i89kqsMlbDCRPBN19/bF+5lipJGT2zYqwrtS99CI757cEB1+49JvATxX+pUrn
BNNgoOR79/rvpra2ZrMVT5SyQXvvaFBFfhWYkPTODYlVTgJ7YBdURLj7lRPja6vf
KgFc75bveH9Jk7nCqBR+Uf3k6S48BpFHY+HQlzM5woGXgCZQBgeHeXxnAnqEa1w2
Yzq/GbQ6PnexsagdlH2KMLDmwkWnIcuuTJZxmYWVRJZJcQg7MhiszQhdn+abmt+l
oVTQ+qytJx1sUZwhTQVvunxRtXbk506ANJCsIesIKBzUjVaonZvv9KWOVdTU/26D
HDUvqoqVqiO/iEPoImibL7oRGUbBqp1vEeF5DdjYVcI1JWz+uwILpLf/jIhkm/yl
QDMB8TRVDERCGSqhit3H0Sry6DrE+dngudfrCtwFj2DfsqNusQe6QGp0nY5w0OwB
DUMmpb+tiEExo5SdY9v4AfWIREeDMkqcvHA94e0jk09LlgQRhXiKsYCVvLe6SuTT
1DQ9eOn2HgjVlhG5Cf2cFvs3AngblPsRaVn6L0SHQlddrwSHnyAeLXwFCastRNG8
CwJzSmDPO5oPHRoORSqa4XgtYPItv1GstyvQW2Ya4VTO0qVnOkMpNwh3bHk5gb1C
clsbVmik7V6b7sfY5FdIbF7WS8N2UvVKG5xOhctxBWJu2ClmhJSepG+d0JlE9eqc
8LaHtwf7lv+wlHjMCrRhuwFtoaL0Q3pAW/W+f6DfEpr+smDbGgIs3xOaEx2lJin+
bbj3v+PFfMlYTjcCvcRj2XKsM6Yv6WPZRJpMMHppaIITbt8GSQ0ULaCL864KVx3A
mX8oMzkxOJAmtIcwvpfY/LZixOSBX2cmhJxCTHejmaM0lijRT4gJZQASJw39h7Xs
AyeSqWYQaGnrQjbdKGpMHuM9IRn1vZzdrgwP5bolw2hgdkeP6HKll5sO+SidxZkq
e5IDDeK8M+gjV3RtbKWmzW24ojkw3wjVrBYBjcBDUqIL50zWx2vAGhKkRGsOpLyW
D9U9YSYSrldLNRvrSqWBrmqKLc+D2rl5a8yTWkTNBtYOyff1ImrShiCvEhk8IVsH
dw/o1OJTRkfkhW52diq7UgNxfXb42lRpCd64BtO4HDeMSnaUtl/JCuHOd5X8nYYs
j/W2Dx2SCpE+vIShRMTjy3g6yzybZHU8ldVK360fsYWAkIo+AD2ZnGUMX55gavOV
cfTB/lDZNCD5DTrsYQj0n8ZDvI1tmf2sKyGpIeUzH78/8dZVxHL86U+KwbI61Xfq
s8M6JDtfKlXEvAdNc0aPkT4omMhI7epKewejYmyd/AaP7vIauml/aCC8Z6XfkCEA
jldxPNcrjfkm+iD6akm7NhyMz1djYzGgpJaqAIOOPlDykd9PhfAiPhaREiEIAMZL
fLaj2ZC8qfUn9Ah72wIA3q2mWbMsoJELoMgd9fwFnwYvHXdFngJbofnMesRZFzvI
zDChBTVG/iHaPF8f9KJGci5azYisKCZTDFa2XNy9LdYbhSJDiJWg29zd3F/QK6qg
UbR0AwHOpyiyNfPjx2mR94NwLRK8bxm2uVudH5YSksQLdH9knggTjv60R2VeG6Mi
qVX1v6uHAtzmwcCTH7m3DP3mFaTp7hJBWbpQ5xjp6ITHUrtICdGUJ06JsOvG2WGq
1XQIF3juU1b5Mh/suwkFRewesVGoWm36hYsXbrXIjzOTl96wu4kYYk89q2uzTLe7
a7kt6g0aLWPChXcSUnP5WLlztugMc3e+0oy4ToXuhcEu7GhscKYMFRkWKDZxFJeR
gx/D9OvJquGm2AfB/NvA03G0wrrLQNuQfRfBsoskzkFyzbw1QZtPkHsYgl875ywj
TtWNLGPUhzrWIYGxHKeZyfWJYLm3A2CnvzkOv4AmBDXAwXpu+gIUaAc1ZUo4ZXsf
s/KqKBWcOCDlP6b6TNU3ULBDftuMRAEhjMVACD7BGqGcX8mFRzImLN2c+0oI4oJc
kMYioW6MbZCGfJy/QRs3Xe8x2v/0sHCaOa02MCMnAVTTFOuo02TfQPArNDHjgb/8
C17SJgqHTjYyYO+bmPt3TFB15so5C9EeTnJerhTh3BFatamTf5Pdveq9S2syw//4
IEKK6lS+MLJe4VpqK9NgLI9wwCpwgH68enBHDcHRLOlxgfcMGiiP+XOuwC+7JM2N
QOI+TtW8hlH9fkOUIBCMEbtcTHycgv5xOOKxH9bsPc+TTHBVVHXCfCfciNDy7bsz
NnH3zGDY1xGiw4rCvsjeqZFKdVMM3XqtpcGMmxQK7sk0O0s6SB6vlp7H3ShNZRif
pmQFGOf4AYq3OpG3mh4dKJJq8Vm0WCU2g7sZhoe84DzXJh5oevb/iduddx9pq/ym
25vfPIFGoFyDYCVDZHY3wy0URuja+rh/ENws2RYOjtaj9Oczs/C6Eq1qAcHjeZ3O
7QGeQCBXURXAzTMS52LE6Lz5HYBYg8npVVH262/7qLj5yfrPPunCdyBDKQNa5PXU
9P+L2v8kCzB6WYOAwWKTCHC//hYcp3+4uPvO0AkdhAA6xZ9pQl1by3rSRqfDeg39
vH8+eL6Aq4WLlUuU48tY1vyDbJg8ScWT4oycy8KaAWSHlZ04WDHuguglnbW+jQoB
aaEJoj20Tmg23u4W9xM0jGMtKR507aKxmfZyo8WCkrJqxPhOt5WcMLGX1zV/ySk4
ldriyvxqkGjxstQJqHgfr6DcRemegJHMr1pw+Yv4b7QQh4a+dvNK3ja9e32PbbKE
uGBb8xzQKjWZwWLdiQXe2M149kpFvOH5311FwBk1O9iIlG2vhrikSjwYe57quZVe
sGPaGDWvRDieyOAB089cRctFFk5JgcbeIAb2NAyu7lWlL7Hm/nAy2Gs/6MvVtPkS
ELmodyt+BK5oAArPOb14vk3n//ViUsADwT7rQV3BDeaHDPKLOhXpcy5kiYZ2Kuj+
1xJ6g8+WuOKw0fGCNgpHMPBCcCuR8e25GIUl5yNtG8jz4JXB9zGjatOIjhc8qeuP
9OP8wC/u6qWqTRqbCb+xLHmQPP5qG6/ALzQtMzITm8dd+LGBU8mdxpLwy3cHM+Zt
mM6xN92iUHG2U6/wqvXL82q7bemv9mCCiDf+Jj41I7fljI3XTJBDg5Y19s6sClH4
EyvR/by+2icOLYJ+oczS79pBg1qpTeR6MXbMxP435UmTzHK4Bot/U8VwshgRkQ9O
GyLiRXyRVXrkMYoq9BAIp/lPdaFElS2+uuGzGjE8zFCDDPfk87NmxJzA5ZefHFc9
Brx2QFj+jFFqx8FtMMOLX8HejIf28oXOyLNpeDM3jFzDEhfL5LDtDdiw2vPx7CSW
YJIch+IOYYHWSOM0H85W8XcbJhlo5JEMUbSakxO8ex/1e4qumgn/Emq1x9uoHWF/
/a7vIuxJnCLXrPmt2+qBjYtmZiW7pkuMXdHnydVOqLx3UzFd5M1ZN2NKs5NewWxx
WDMmOkkoHaVjNln8lXjqiw2aVJ/j+NE20D9c6XhfRdNkT6yBVrg9qVdFsSBPtVEy
ro/FtVYVUH9TUQfYlVvKYxdXQKsKCON88xg/T6z12aWlTEAMWmsDLXCqVkVyBGyt
5/tbeVbcoHEFQSYQ1AwNt73qYac6+2iZYOqTV8xHk8YcXDlrEJviOwdlkZawhzqx
m0WNK9zCfi9zM1YlK4PrB1M8tIaiJiYo/mOU9NLKPYmmuncqmLMqdv+VNbRNFOzC
EP7rD57KF5WOhdwy16mQySSCckrRtksoEbtjVVwHL7/WanVpFKcO/v+cg79Q2hUJ
y6O1NhHOZsJX7shvv9oZJmGDk/1aPs2gFO/D2Gh2Oxi5g8A5aYOKpxBGrckNcQXM
rOScSVX7jXDTJsrKnQCUPEq/JGxVU3hAHU6NY+oFDQ8jcke9nTJ/y+r6+sYXXgnz
B4lzuvOxoCKC+1a6E2cUlimoma224zK9w3fnHCGcK809dFzWxPbfV45DvROO4CTW
FNCNa+AGtIVWQu3ewsrsFldxGcKloPzq2piY+AFNWoOe0SCfIinfD4cscpoPdYtR
L02fVTI/WmJADTa8Lt0FRtbBQan8gIDoeCdzT/UiuAZU72ec6Xc9ya4jopfqNgIC
bZHZSqqxVSmTIfpk9Ws8Z2gXPu2FUd7u9GzAGnRwgA5wS3ZyYslnFlbrNtGzq1Xc
YmNpIk3jR3itVhJFkm3B4mQH5psPveW4Bvd93/vbkoflRxd9GqmtwmhCxWeAUNEW
ppdhokMHuXg89IHkCcrt2bqafa97kpRIQxc37CE3NOY2+sLmQb0aXW1VLz/nr9Go
r4n0gh5oVFr/oyTsqAdsjaDkvcy27XWuAg20MOIETQISA7E36SXRIt7qc+kmTVrv
4qnWTOQ2w/lsgAtW1ZaBaaJI6uVCywUmV2+OVoXvotrgJHZK2PgFHGRV6x9hkwIa
1RjC7IkYV7VOpZyuLcPU6ynEd+IrxvJ3TLPMiy3S8FCZlJvnY2gkSXe0EM8aY7Lu
R+IyuKVtS41La6kOCD6yJCrR3m+vPgHHlzDpewXJWYmC9NikKU3/F2m5joaY8YMu
j7GxDdyBL3iqeCPkClCkesAlp3I/6VK1WlyZ6z3/xpphbbNhPwQcc9Mk29rclV7E
bLcMpXynncTtvUHJUMf4SqQpluzSNoKurVTnzmvYZKjyZ88Qvi2WyNNYnearG1dr
OHd51JXQAuiiJh3OcQl8rYTdQXnNpttHvZJm96mEp6XSpKPDZ6BgH0E2YWHlCk8e
ibGZvPHwbsHfB/4oVnsX1FFTk417i4M5h243PKlD8D0uPoyfffoPYfcArDIkXLEF
mqnRocEVgr/rReXeAreSxfdn2cSNzYt5VmVGERvocObPQED5kXiGWHN9G+vGpaFe
/4Z6gcUe72uJgYlsrXYnneRFbsC/W+vgvXe5Tz/DHcdtYbi5aoj39Oh42RDalNqG
hkgNXKlloszG7hdE6EgbxOSlff0lkxuX1rHjKGzFgSi75HwodyCudbENbja9QObU
0YBuOT7O55UiAKHglgxg6jLd+5dSHLlZceVYHZEaJ0vIbWEqUaqmllTL3bjW26JH
/kWj3T1Xco0JGjY7HnnI3ccce1HC6/SLDzoVbIq0z54ielvlOQNmr7ybBivh13CU
8sJkPve8HztpZSn/jJnRa466I37mMy6HyooRsGkpjwL+AVS9KvQrhvcvi1RiYBpl
kFUy5IiKJaygdgUgaMnoKIXJgy4tRgg6QSuzdWLp6s4gAll7Irm8Du64KFn5yiJV
z/hcM9gDOCiSCEsajQk1nqIvTeVdMM0SqAthtGQRTGJ0gxiH3hNC2f5QtMxYQLpi
nL8vZjvTDxAq9ip2cictikikskc9n8cUPuD98iRTlcE+OxDeKoZ/q2filpLNJfhK
olY0b4crJmDE7MVrJplPizPZhL8pBXmBL/UPWun9JsIC+iyDBYZdxtZyt3TZwutR
TdxnmTv4p/CGEAhWQbIo1As1+31v7SZDPPd01rxpmQ2QrJNZGK8WMMbmzaa+3KAc
Mkd65EvtXNW361w5BTX/v3pTnFsZ+FpTBkNWEMDjmGNHJdfRjI07hv30F6Wak3lc
MZAKKtt8hT79rRNAMbY+WsxOmY8BWkNwVjorja8Efd9jX6Ji68g4Ry9p8wKOT7uq
wlRMaFuPmrEgx5YDBYIlAi1AGLET3Dhg2rEllwmCB9S7u6lSPiNBFuMN8mC8TbJ0
wMC2qmTPJhj4rQZYlFwCDtEoju/O2lXHzLjpWgm/HA4/sBTD6StS0ynJaHSPGcAG
OE1EIzbmQt+KUPyCQz4fGA66VvIrGvYcL+6vyqU+BRXHyYNgetHn8EAKDcsFjjWE
wmvc09msgTgGtJg2+eWJxtoB5UkCx6TuMNFcthpFWLDbOcbBfVt9MtClO72kz7fT
AFi1KpUGDL5Ws3Vg2vtEQ+pbR+ac2ZDM3DPLj16WFEXjD+ZqVHchgXRx9mwGrfWn
RsdFqHa6Ka5YLqqUoVlolETSdKFRA1gIQtBdWqidqYpLbEAdbTo+Hz7I6gjrmjML
LkMPHyKGbHHzE/AGbjgVttu4t+XGAJiVK79KF31Lt+jEumhktV1dt44yCb9jCb67
5bjZ2mnavskAdkSJoyVkTFX6/pi+Fy1UDTLcwZ8jN1OOEF0jf0OtWJsE5e3JDOtP
zCGxrmrCq5Jt0Y5AuVrmVUBfwC8nm0/Y9ldhi5hrQF/RNIXYrWkWcKznsm4JEcfa
s3pfi2kP6t0uzTV9sPDfhnjetvp9r1vjJnAxj8D/Bp9C++rrEF6NNwd9rkBtbMm0
aMHoCn2ApIZSUAEHt3EiqA3XrSVqmEupWAcfxNEV37iBhJX5npZwk7HTbqUoEmun
NXsDm+N4TAwPmilwDO/noxZnV8tFwLQKpKapzsZIUSTbDfJAW+GVC2STc4UWtp5b
iau3MYcQvq7Z5a9JhaUwB5PgSm7kewquGBi5OG3XsoKHMtSN0Tje8jDRt50tza/v
UStvlPmLL52QoGM5c///YICxgXfYIfU3gO8gpJCEq1Q1sTcCYZiI/nSAZfC16bn9
sI6Fny+lwdDOSOqVlCkPsqrvWJEmPwPjY+lx1YTHwqL7LzMugtUMcP24Tlvld4Nc
hFS+gaYqKiSfwarG5ZmVCOOF6VFmjioB6IfOt6/OxYquwpInD12dGx9QFgVXIk9P
rzudb7XitJ7KCnbyQiyELJ8X8+yP7qWB90tEioetUNxsctCdJ+Zam3w+ufejF3Dq
wdqOuP2PFVlnpXZlIpqr1BeH2xikKOHuvLFUGeUi5s5nPoQkajAYhb1VLr43ZU4R
R3apCyD74z/BZgZgooN1TFamlq3axpAdnuWpum83JzwWLty1rtecwJjTTsMYaG7/
AtgT7QDRJzq36N97G8r0TgTDC9jGl4F8kqtlEn1IsvlNbJ3S3SnUEXHHR17QF/Ob
Qk1l34KRyWuIWeHN4LD7jaqftZpK6SF0sPMHXXYQNnX5ZgkUSxSk7Iqm9y3yfWau
XzxMfEcpybWPkMix5d6HKZKkXNDtSkLVKjeb7U6boQeGmEMvryrXDihXAOQrJrtq
1a7HNQJfVpyQPULhEv3vCxNAOBHgPYSskx1XP61S6cCkqgNHYigKvcNoKmtnQyOD
YAZ/i6IeqgHGBqyIlR9EKdfZ0BEz1TGHKMN6mW2hQDL7GUAVhY4fO4vC7z9zlMxJ
P4Gdmk8+OYWv5UJstYFwnsMZmjpv4QKdKi5zk1tNKcNBZWKt0ftOLlGQ+ysBViJU
9sBjQlAER/J9nNIuqXXF6AYVU9k6nOq2/BjSZtFtwaoOkYN6k88xChYj87Kcol/u
vvlBLHn3SD9y8B5Awpxz3M0t09owkl3EhYeRRFOIDeo/kNkCFeR1qUkKUgG1fKbc
tRRSMYbkcPHCFkx+h64RcHf2zkde54eCbZIjcBJ0b7Aa7prNowd1EbNSPW716utv
Ard7g5sdXfABDWHdO8JV84FqNko3Lp2kylLSxOdS7NKW9tsSi+qI7dC9UhcXMXMf
iu4oeI/joz5bgnW4vZ1hnFo04n8/nGcxVMt+IisJgYtfQmyEyeUgXhP1bLjuUlP3
IYWD0OyD07NAd4uZSzjc+xgZqPe2jL92xzPGXe7+gIwNWLEB3d2GyVQhOocvREHX
vr5K7nB6ASbIZvFynE4YNUucU3n7UrguRWDd9xYSgPsY0tmG9WuO26Jv9k4p433f
5AjXJtlEyR+R1BLqvOSFZekLMSmc+pMNOwrjzti78eWal8sP6FAaaDEMCfpYnlVA
vNcHG3nvtQSGOmY31DDu76HZIP/6WHXNtt0TJGDhXtXC+YcsiMJ/8ELZFdiwborP
pY/EwbPIeH2DgUoOJTGMhuTclsnEoVkucSsUDCQ90rORTHUtoktmRXFt9//sk9wB
ut568Kw2xygWxLiI1jW6lhsAtRzfz3NjMdhRz2kOtdLaybWaPNGjcbvEx7HZLBJa
aTJ4bzYOZeRGoadexF4IpQiufbx0mXSl8pobrqRC4u0L9ePbwe+5q3Qo3EYS4DdH
EQMpzJrR2TXic5FJlVI5B/wuIYDZhDDAduVjxIzxc9ubpgUUhFJRJ9qoM1ZkFFK1
GO9zGt3Dk446Gxf3H2ToWAmQDGB4bgIoM1rpj3l1xUCb+KZsX96N3Ph3HzGRSsLe
FFLSlX50x3/anbACqHxCXJSwgVhfxBxfQ9LzDDFXf7dXF8WKWyMZxuCw+qIZv71z
1EoQ2mtfHdWPgZIrEbgZ3vJWe9IfwgoJhL/EnzEzQnJLcwXACHegJe7hCvbyPAVJ
m/0zA4ayqG9acDq93i6f13fA0C3JpvsfdhDMkT0CKq47XNZ+ehOHXGKY7+UYPbx1
vzoRwFfT7WytfangMN8Dx39xSCLaJIv0Is3iPD0a1wcV9QQ9E0nWQ8GxUosA3zeM
SbPe8rJULv+cRmzqYNGzdlMPv4Em8NL24Qth2tuIRdZJ+x2OgxGSk1RQ1Dg/CS4a
loV1Au7PvNWg+/AaiyZtoTtfh39RvNpVESD+za4PqX2rJ2G2IOgYjqBKXOLXA2G7
/SZYjF4i6NNAy/P8pX4dEpgwd8vSGVrPjVUprOfdYLnA+y2JrsvHywRnpn2CRQDW
MHxuUtY0J7vsgbN2pFadozOnDMiLG99S4dEYjhwCSPhCJhkfCclBaKRZC6CoCcXY
8yp1RKBSd7TGvwl8GTo2XkGIhcsrvksHPl3nJRLGT0DViADbgduIBQR5BNsJ3+s8
bENsTRaeu90ARZnSz5AdkmRwTOYngn5vlcs7RScKPUVfyNxyIDJZ8tNLXMQRao2X
kXtbq9ZMWFtVnFMzQcZt+GHO0AcxkYq5GxYty9UcfZ6+vPusW/cV819QWTaA16NZ
79qJsQbzvT03DH92lurKroP6Nk8UJQJZthljz64XxHTonJgpSN+2fivsEhQm7X27
axTxAoQfwyV4m3POofS7RSWHP/pQrgunW+mC/mMun1v1JzlD+npGi+cjks2d/Iz4
t0Ye3B7tbn9Awp/FJyqyGIr+8K6iaCj8tqRoZnuwWwjwJIMf6j+7tfM/t459CplA
X8Ao3gh9AD1HnB9Nh4QjvO0cckV0b4+zLjwgGxbqqXcC9spp1ebCVwRdZsiBzBRm
jjFq1DAjzUdeGy0ZzjZjomqS5c/4RXRPE07wvXhc/iXEDu7m95ThGwia+8t8bLnr
vwEZX8XHWen16+sQuVlMZjjuLKAFqYs1gjaOm/A7UubF65U+61AScCd4lq5flgHs
H//DILjfQ+TmiMIKXddldamXRsb1G//LMx/lnyGnZLlz6NjNLcvn69XBEeb2NKPS
ENOvRThPeIY9a9b9paopwwU+LbvSn2643J9HbS6VzaFNH2dRikgbjIYyjlbxjchv
ki4C27Do2dKVlWHzWXjYYdjoQ//q2H3nUvT9Ax+MycVSz/KoL5fzXFxEacr0QPiE
FaQ2ENoykllOufkYJBfOwB+lanR3Wzqt7ES3+6DjpRk6xZ9sgTf4wC0vWmxbsKFt
Be95nMNP8DRe/70/EZNf7rartpq0jMBnNwgPwowSQEkchv8k0xJWM/Bx6j01fptM
Mlt02mr5r6Dh/UKN2ufZxZfpRFocG1zd7Q+PQc2CMt4OnJXgwPGna+nCfdqRzlOZ
u143ZSuU9extpoRram7FZ7wFErzrN9U3RPhg9C3LigIW5b5e4MquNZT8vYbfYF8g
AUoj3VRbUVNAFJ9MAOUKxogeNSSkptREB44z8nfpf9rlbTTx29uw0/ctXoUcwP+2
/mZwM/iIP6FcmYiBPPoMWryivmF9Eg1ZIQ8XOWIwb8y0TwsNIX8yt8xyO7ZhkoC5
AO/eEGN6nsmRvKlZ4UN/ZPxZa3WQNFLD0jM4or9llbCiEn4MWBDZq1+eZzBWd5Sl
SJ+PR+dkG5LkXISYqe8fEo7N5FmLvfTeFjGo4yxCJtsoZM1lWuAwHL0wCryovprB
0A4EAlYdtuWfYB5eiPGPS3ES8BaHzq2VfKXVpH+H/+kiLk48tLzMaA0tcrUTaqP4
gBjj/kpiYGjcklbw2VyFs9365ryTe/gQXjy77yaw1J9Mn/Og6cuf7aYUsM/EYlnG
GgSUJh7mdf4y9VtvEJFJW3dcoGbasCailYiQtT7XVmdLLl0qiskDNBkt1Sx1AGMn
3WHE95HscCPvNxp7dim98tRGroAR1UTCGeJqamEG0ERtnecyhx0BjHVNID7tfI2q
oKaNGKMFo8i87zwdZ1rHzgenSdEnhANDRVQNhk4ab0tyRpWWbtMUtus5mz/yCcIe
4TcJLc00fr2NOLeV+xJigmAwsjHa+gNmc/HbIRxS+5IrcxuArr0keWvjOg7D4QgO
bW1t4T3G9Qga6Rzq7za0z3PGe5f4RvI7DZEVjSFtLS8ZkUo/Q6ka4hT/cgZOdscF
pvE7cggChZMHzXoGxNkCl8Rdlp1auq3m0S2xZ4K/5rWDsVEqA4dcBVMtQ6EL8B/J
wkWIsR/xQeOEi3OOUTc6ieCTF1X3KJ4m2JulhD+JaUmbDcyfDmyy/dBlS9zvt+WB
k1n3T1cXRZuwfgq3M5VNunWlNg84xKmlO/IAAtxZwLehgcIk/26AmISQSmbcUAyu
bcPpoLlzxgKBC4z120vdl0+jMpTT79UVRYH09n9QRPppVVLfzBzfKSe/ATKXDvos
RhS0jM9AdMFIQP5DyYFrE6a8y5eZOHp7lv5eAaHz2EeZMnGJlcKfkghqrA3Spu3k
f5XEUK8NTcNxnkD+0f0selHW79Z3Yaqg7WB3BALO/BMXU6M6fLuiinMq1UlX2BzR
IJPCrMGQkwb55iSB2IAHxyLwiyB3yQEgA7jxy5UG9Cgq/LE3AApriEQDhetyG4v/
EkOmS0AzwMwKw+jvDwky/Neg6a8q/EA7anlvGvvWFWfUMvq2z/NZMhJIRrjGfHKP
mUqz8leQ6F0HzukWboi9hHr3La4qWrlxOvYQwaYonG2jGF8aJAGdlpGIVs1ABa1J
AQvrqgSJg5yhTyH3o1gwFWWtAsn70sA3nmtON639Z0Fvvet0RPtACUjnMYfjL2do
g394D+25aQF+ShrwozQGKj95UKoTbf7F9FKLGT4RlnF7SiRPUtM7ZMTEmb+/W/3F
wrsBEuq2HmYUu3QH7maEZ+OnMGedItzKh/c3HnGplJVcjzB+9QbzGFHmXbgTTDnW
gsl1zwkNHWPRtHFYRp7eMKr9tnJcEiGRbAYmuPNNpFkfgEP39TdY2/yRaREhXhsH
T20lVGEmr2pN78m0ybcE0brFl1H/yKWCrrqOYhMCY3lgh1C6jYGnpSGFHSdzJBgc
m6zZI5Z3c6KvlwKl51tNKOqILnsPI+lWy+0t2D2GYKjgFWgf5C/rafV6MaZJZRmR
fJI9NsLi4rHd9/P/E6xo+4lh+zsO838+wiuB30N6wnOSdNWLFGv6i6Zefu++o7MO
EXADWms55E4ANXifAm1GBJhGzxllIlTOcLYAv0Xm4hNAegVbZWkYl0ipnFRkwrXb
Uc2bAXXMSL/6eaWdT0FITk0nD9HK344La8HTlz0TyXtNGSdTN++RXedGJJtSDZW9
usH9viA1lqQshD4N4DMgWeT5V+QJrvbsbstOyL7SuKtsG76Sa1Wn91QseScparkE
/M4S9n0WD7ZQYUZNnFeuGcSRjCqe2C3FMuHIJhLROdjc5M14nTRF8SrgPpajo7dS
64tXE1zPhRgJRJeRjrc3novAB6prDQWVZzHpODkRxom2QQjrzBoO2vLFFEb8bPCj
QCzha+CP00sRlKo7f/9lE6pibqb//dLcBWpcCfgpEc2Vi/RLLe6pbcyv4HMoT7bZ
5rxUNYEeOFoTU937bDe6JRwar1qO9GhAQn+iLCNTkaThmBNBcEta9hUgc3kH9ogJ
cD5sFtvObxkS6i4OroRiX2KKr5E1ZfRP4IxP7ujztpJOPOgbFYhTUfezKr2JZvjk
QdYJT39hdaUTz9NZPHtPNM4i6zU2pmgUIJqxISxQKKZAsReMMp1AItioPlXZKnAS
oYpzctjnkbG4xbVNVkIdpQywf4eo+xgc8Wnjhw+jePemGgrvUjNmZ0hX/tZUsC/w
xNSCN4q0zGLZ3WlO4+M0fUFy3b9gqPnJFZSmIrPungcSAGIf8wI71VIoQRn+dn0h
YpH1QLutvmpsuuNofV63qhUt7p2L5yRwRtTLPieK+PKhs1BDedtDrNraT1OtYcSl
JZNrFirz17TzegKyzPs9o+2M3SJO9J5idqzqSFo9aVSrul4eR4PT++I1UWC/X6X1
erpwZkLLTaGiPT0+3LdMp0G2bti3548Bht3FBrWagj49XruE8suIvqNVIjW0wtz4
+vrY+h7xqu7sHxaRc0SxYj5GI9ZiR8ZCV9GsnijKzEzsrucUzd7vtXYrqm0Gytu3
r8FTbkADWXmbLgP1S2iCh1PRg0LtnzGntVXTkfxsZzmFgbHypWoSJqak9a0hcXbU
RQ7TBSvZ3IHGxSZPR4JrMLGsItlkEeSNqkA0Y4+EbSzb81c9e1yKqD6S32yomfT9
lWRmKy7A/qZzZrNsbqfzEhejv7WEj+SYTiXqiGqBuH4MHovJXZcd9E4Kb9fZmeXU
y/f8ZoMqIXzIQsOzoXatRu6nU+3QwWGqsIBteKUVmWcBra/KQD5serNipay8lb55
3keSdMcft6nGdZ3yBSAhYvJUMG+DeW1PyvS88ridmQX6G6uUrVzAat2cV3L6Hwqe
mZU1P5tFSaGdJCFmZCF9k+ceZqQj3sfhjJeyDQ9VTlyPvJnmb4IY0PsAR7fHb9BZ
6Dywdw0wxMlKC41yvCBEejbk2AyZapCzNNciSugZdFvoGXB3XmYrLSwqtjEvqW9n
qMPXvLwbb3p5GyOlP10j9ZTaNsvMen4s4xHgvO+oV+c55lgv3PCRCMBbyrpQpRyB
+A6EsLvSyu7wQsMCcSAmUHWrJEvOtZ0KNP4ayi9Dgwz/1cNAR0xxDwW4M31/Mo+e
/BfxUDSZzLKoXbzLxfU0h0OREQs60I/3cKN1abWyKxLGmnal5zWpK56zngsJ8i1h
38poSyIr2eqiS3dYVKGuuQ6M8a/BzanTjjqJQ++c8xskxRVWcST+NMcGaa2DRVV+
KSOJw99M/aMvdAPnYzJ+gAtTf0zD2666hx2hbjGSxDvOilenBxmmWyE8+XgIo9qP
NMtyW8aui4HaF30gUX6BuupAQDeMAs21HUitEWfG7/PoL2jfKfPAAV+LuoUTLS9q
P73RPhesv8ypOlJbPapy6Wel5fqI+LKeR4ih8A5gq3XfsC3nAUIdq5RJFXZ60j3w
IQudEyk6IAB8XYFL9MSsw+f2xiAJ6Yq2xWCAoajS+SUhpXtIMiVr7XpHOFu1qzV8
+9KpXonrFQqNO4k376yQgrWnBu2PWqHDXIR3ILO8sOVRsROnn5IUmyJwZSBJT+b+
HYU9/gwJV1AejX3TlSRoCuziQuWlauXS41Em0yQljAkLynoQAw4XAIMh5J/81NRZ
jelPUusPWv3PJOZYNVy8X/eqNVX1BQcgfbPQ+P6GajasGdlgEfp9yhaUT5GZmXP5
JRV9Vj3uZYbEOFwCPKY6pxOwcSQGqfIkIk5w16q9k/3VGLpPD21hUskOXRzuPM9d
QyG0oXqQVmPm0BDbJwZN3Ivc0FJmm15xAbiVDgLPrzxYpamxlej4LemH7iOPXB3J
90EWIe96tOW3NOmBhIu0DY3wxMy2aIerjeOuGgFrXsTNOsklINdRrfwM0Or1M4Me
rmlJANgAAsMQknMZ0sQ7bUQanRR2voLgWCQKzMkpY2EUNHPdDKPIaA4SLPh1Wscy
qFhS8RVl/QiwL8XMfY6ZheOlLAPWmOURwFtjHwTvRxXvjYpdy1VEvGWfYbsPbQur
FLnWz25mGqJsANZQ2ouCuZdD1ZezRse8HpkAta7CfARZgvoSiGAFtqtLbRKv10Ss
Ntu1WUOhKI0/irOII2O57Zj91bAXT2Ho5PM5h2WWxnd3JOLagjIgBcLt6R1dVUto
td+ZYkbYORulSFFLMejO7ooTfeaRMjqeVbToHXTIsgrzxvjP1mZc3HErgw7cWyCf
RzrWlEAIj4BLX1rchIw+bDlx5ukkRqClzhbNrBuypTwCnYeTJMX+aHPCL9hgRcSg
zNxwXQxcvR/5BPHGXWQa05QdTNX33LewpiAOPOgYd3baekuDpIRH6kSA52tU+p3T
kCp36n9ZlyXnbpxgnyD6qxKwCu8dJkZ9vzFkXkNZ78vBiOVxMT3mcXfa/EzZeKy7
qEnyPVpxzCXrPtwR0b3+Q2SyenMIy80c5m64bywOeW2aACaKjeFJlX6JZsznKT/8
yk+JhSuw2Gz6P0WKCgYgLD5cBYfDuXfMaY/j+vF4zt2I1SShL1Q72L4tk0gpIJp0
b8KjkG7pZZYn6Xxb8PQ5CkjZy4SCAYNJUqM5eWCj7FpF+nt8qkncOXENBqWiPK5S
SgulPc8ekxYKUc8DKsbeYAhPc+4veZ6kU/LUlGzBWgKgYkGK1FgCJ+KuFUsNIrpC
sgpaseiQSUmw6JtoplNrd3ca4NM8E0JQMFF1KTrBrGn/+woha1pmFUKtKDhb1FMc
6KuTy9is/wFe5JN/55gXfVKOpfYnDM/f7k9Sh+LxbH/UN/PcgB8YT43pJXXdSsGC
TxRm/mKXZjdksl6ITgG+N7XGzDjH+nSGYTq5HdxgnolTBU97rkDJqvHItA/tyQ0z
UWMXfUjIAF+hkznnzH/BRUunLuh3S4wLGe0lkwKJ/6wKDcJ78JpIb0ym/OkifUyv
6L5giG2LCDJslk98EmtHZO9KdjjbfivntqmAb3JfHZtQa+riwUzceu1mpflJrfDI
G6dO/kDovtFiNeeu+GwrgvBHYwBMQ8zLveej0RxpJhsvEtDj53u4oL/rO5Z1MIsK
Wj7OWsgU2dFVdSWnj9RZpULUyOEyPCCJun/aMvHTSQBaLfxy5F0wWgAxGNmrNsZ6
RxmrGvxeSlldVYTcX9aaSJluiH2lVAFAYG4pg2HuHKKYsh0IOv8qNjf4gs3sOHBd
T/rGXGtf0Ec9daol1Abj9g8Mzq0asUbd8kgDyR7tXUP5CberEuU4T951vl+iEQFW
j0VnmpNQEGP+/JKjjKfatfmDDuvZ9VnV56F+58f2V0Ds5urWsoAA6qLBMcGnG4oO
WYgim0o5DTVpXt+bvjY6/uUEcHtiVQZbDZ3Eu99/8LLMZ1SZVUTAaqHn5qWedOUQ
CWauIiU+C7QyhEh/PO1cd3nQPh97pK3PCKDs6aLVzz8+VinFWcg0lgp6g6DC59WH
pfkuD40MsXK8IirGDOd/oCMlEiATYeOq5s0Y8xr1aR3a6IFLVKB855xxpoH2T+As
4eBNnCyYRi0mLhORwIK4uOIPRhdhrEWR/BIRMsha9G5vmGyX4G/9znhXLrNErg7k
9x3seR4czlRPOJD1zdaoLY1ZZD/oebBv9/5p1IfXEzxceO4poIHh6YYNX09S21VZ
i7Sh+nOPWz4A7EF/kqTc6rfRYOJBb/ELWZHiqJgKVJlnleGNZ4daMv4cleJPQQBO
NEu6W/7/BIqFqGo/cKHAYWvuuJUcnhH3AveXiisPl7M/arX1BMnyuh5qV9PYh31d
1Nwscc9/GaqVCcwsom2GYgv1QF6NQ9qyz2EkJRIzjx1qqsQ1KHwPID71JlGN4k/V
KTEzvsoU1A2CwmYtQxX0aVNFMbuG85Ep/C8YYNbFhdqEcwOMgwHsc4kNRm2BxBEe
4GMnsa8XoRsDE8ostLx6Vs4gxaxSjw0c5Jhc/S598XtWn9XQz6NVWym8GCXLkuhk
XW/tWRB/W0ux2GCxHZGUwOB5n4nQeiaU40VcHKzrrSZ2iQg0llSBfcdHTEt9Lg4/
SFOLh1SMWP9UIYYQbRKTxlrOjXGsE1BM3+Hq0S8dcr59nA0x0bV5JNLrSEvVyO7M
DdZDMoD4Iz3WwojGYqCyGzCzC2LQub31OtnIVo2r+K4sI/cIwYQD0pxulJ4xES4K
uC7S4UnxJ2Au1tw2BU3LcSn41HfquoRqHXRZAx/OK9/4JqjKTcfxnE2wrX+gOPGM
tuKV1JuIjoEVodBCbj6Y2B4syPTdnvYMIie2M+wslMdFMpjDt0vMLIIzKPfoYi61
WYaCO9i5Uun7e3+q6WUEsuC/U3Q329+rwecoKHb8KaSdtCYsurRL6fbxO7kT21z7
cGNkkg//MfO17tAKgqfVHct3hbU9qk4qh1qDCHdMyzkHXgGChw+IXyhnUzqz3xxN
rZMG1hobBcfpQebGTU79oCEaEfMJkqHpqxTjtYaBcghuSKcMF5Lpp5sk0aDCPCBy
cbHg9ePdPUQbRkJj3JxRYLujpIDG9d0aqDoeWx1Zdu2PjyLNYGAzS8HcVXDjOlZa
TFc+z+7ZWMrxbozEVbOrNNAoWSSMrKjwDnxiLEP9+10EfWfcANimIElGF/v5JgT/
pp1+wWE836ejd6OvPk3aQ7zIMXAVvh7CsaSRXxVOutGm0BYbyaZ6sJZJ3u69m4rl
Hh6aS+rRJ6qdI/IbudKBW8AnUqWQCZXTj/53/l+HvSkgFoGRMcR+m7DgdzbApiBT
1oVIAW9HYDvjgfz94JvFazDuBi42cuzpOaB+nZwotf74z8b46j+qy9pq+Zli6jek
61ZfAlHLIbavZUvCUS9mEJytg7JG8l8+oOAseQnla2ZOcFziRYkyqurmUib9e2P8
tWCjM+oF0fjHminar1NZtyOV60lHTzv9g4vmM53V1pLrWOxhEuuP/7GZSbvnJaqq
+MUdxR4PZyHNpJezHsegwKMWGpcGWskVafY1h6VUPgmvUMdsms0Z3CFZf7e8Q0Ww
Mg7lnHrW+5GOQAdYoFt6gpe8kp8eGZeOYiqBvO3lm5/UQ7u1WRMI84We+O0NBNaP
xQKaOfeumGwdhrHEeYwkQDvpNCRulKY367LIYfrlgoFmImi/iI62OGRxIFmLyCZm
1MTACBQ2ACj1QxcVO0lie21FogddM/8SZQf5LpKhWkgfv/MWJMH/pDoQLeUx2ZZ+
emk65p+mU3fdaTOgQE5n5kXWR1O/KoiWoA7nCzTrSGLEkvFpDDyY/NGlg8jqRoyb
ww3HOmp5MSn9JmJ0S1VGzj+c2t6uqcAjDJ5oxukGxCo2Og1KKh0hH3VVSB1h1xmy
JG89vvy8N0OM8pT+pnGDugtjlHEyRKs4W8AwFUPPGpqxgqtI4qBwJdl05AF6nsnY
ugY+cngLNiQiwlbicRMbDDMsmJKpg6uAvJ/9azGv8i4P/oxPWnhVQUl+9DoUCc6/
DNx3ne1vJQ+zcWUxmW8Ybb7Xg/1mBYG1BEKIcQzoDfiow3cKNS7KOpn9wqxBed57
9EPIOdab/9vdaNqfzedTU6IIxIv1imuHhjgt2f4pnkk9l2FqTiVN/4dUMTLsd3N6
EEjAGdRvS9sTXeAIIx3ZcNWPqX/cmj1qFmJXZIH8uQE06ILiZ08cUIbGnweXkcEU
KU42bugBXAxpG95rFEimpUeXbTGcK39wjXRypK4xBqjfyuWT4JL/Qu4TGV+ELj8r
ov9bAfiaVNgfmqNZkeefsp2NXEFlwlrUzOpwCwWWd9OwRu5UEf11c9uqMmbbYUJv
q+9TrarYN7q34KWZsHTRBjQa0EztJTRThCViU/ARD0xZdUHGwn2/fmTu1TVninUe
n0L8GLRNF7lFxczgBUqbYTAw0toaH2jn7vm7NnvSBeXnk+fn9acTF0y40C/23UJG
ka1IEq0Lo6b0gMbRivZmKZsm9sc5iceuVfbzSI5lub1/xYFZImzO95GFzI33CN6L
icuvKSzUf+n9eTbAY5QR/u8A4bSWA3U5VokF8c4n6/k4bB89KeUi4dWW85Fq9kEu
2Ed2b33oyPZx5lV0HupWfHG1yHuUOxBlrmR+yhKmHkoM3K+AoDhxz3YNyApLPSZY
jIUiOk1k1bMMW0E82ntllth4ZXhu3sbMs2q3ydEGRDAbVJZ9gwsjhJIu+7NDZsV9
wH8AvdtZFo7401XnjtkCvQHYebnHrhpw9s7DhMqjm7nnpBbeompQCsTyGRFAwqzC
HCbBaePCuucxVl9b8VPNmwaViJRaHc/MXOxPNEXRipBoWhwre5CeKkPPbOTbzqxT
gZX1xqls7tAjVUge4nYOqGwVSKZaDF+xtTZwfgkaaRwyJhHEHULhquSt06k07Tsz
8MasCjQwFctPIk/tltgPd7CDh+f/nQwsZDiODZiwkiZlzupc/vb3nAlKL7a4DhZW
vhvcuAs4mrFhicNAVf6KWUvzMGjb8n1rLeVNv8+zRF71WG9NAl22Fi++yaD1+HeT
HQBFN6giG6S179gQhnZBuLgSEjc3pgJ5qDUMfDKFq1m37Y1zcgJHz82r5zlUQfIq
umletVOtintlkHqpHYcKmhhpErMr1m4sRJnRktcDHoX7etpHWtzD+lSDfHg2mrlf
l8yu58wqkGmko9/WHuqZKrir8+t+4ntR5Ye8tplZ5Uy6STUNxz+VuepwAASjkKxk
fU9gbhWwvZ2Q9DXAEhj1F6Pet3WGW0dI49an6FYRy/HduIVzTJBckFJ7W61snGKf
tsmpWCFpr4u6wCJ0WMMKVf1ckBAq32xqQpsPIiduKSPZqqHsWgKYRNIKNmTeYAW1
sALpfSOU2AtiezPIIzLDSZj4FpqCEVnm/5ZAE8pkkSGR2EHrfgwAjc2xCgT+vqEQ
LDcGqwpTnL3K7XuWAm3Ic2EAnUNuwtzXbb6xRS0PubdD4ddgZANGi9p4JH6hmz4Y
GJu5cAYRKrNPDfPMHaCbZh7k3JDl9NQMmk/8EdaiNnot3n5qo+VPzF9o8asNMB9r
OmALz9L6x4hDMRHhskrJgc2e31Vd1Z5KPIVbFM+wIFEltT3dblneTvDFFZx7Rv1j
4wYFNWT7qM5bVp9Qw6uB0L6CkFQv16DXbEB8pP+Y24VsxSZiBCDlN77xx0UNhBtW
TvakZds7fvKyKJhnI6Hsxi+8hIzUXFZTu1ucn2BuRngU2Mv2zR2bxKRwgfoIvv2D
92D6W7YTSojJXL/mlBP6ChmHFJ3tjbpiqkAAeVYGpJGTGVJq//j90pXTCVzwrUMu
cpq5nBinOZ+mOeYOrjNS+HbdE05PGRPrfIeON5wnT/0O+JWXZKjywVOiJBEBrKgn
npAV2r1UwUl2ig2EFaK1Pgv2n56cQLuYkj3ZMlJOmjYf0kvEMgZRGQNtvz34Y2uG
vn39CEc8ARx7pznKMeCWxV/gSH2PGojwajSs5anuZLnGqle6Y/Zr1aCbyfp31Vhy
4Eyri7UAz1tTYlUNEyfeqa78HERRVyVeYZYIu63K3se8XQln5MXuE40vToUEnMKy
OUAxUMtrzzplUt1mbgtyCwBIdHdsb6ed5vIpEvv4QPDV6SFpX5TL2acMnC7Wi9Rc
7TThv2EFwutLEYaQBojHY0i+5edEUz3kj1HDd2z5axyZlDEBS3unfC+NZ5GWTD73
p0K6ASwgX/lO0T/4t0ajECbrrIhrRfLcJspizng48xbVCyjQCWYIrVjX2/0xAHWn
83N8eGwz0EQFY4uWuX7cF2MsEej5PCd55Y7TGp/xVzKGvJJPFXbQeoPksrI9Myg0
eWdDdz89U/bUI1/faYPVGrIdH4fKeBLhu3KU+PsIPeZf2oanU0P726vqUPvoTxNa
kN5aBMt9jAIbpy5FMm5RxCx/NRez+OovXUhEFXvpb4t6BPHGRerN4nq6J0p75o4G
eJBwLBrZSjgX3apd+3eoR52rnG1lUbnovvjQD7Q1N8nYnrBuyFhNwsgpbfJx2NRs
FRVLtbeNcnZLVTiBnyMjITJSocPVB+twLXq/5gWE4hINM9GTyw5Fc2yrtu29D+kj
ekrrcTTF+dYLJAgZrd71fjjO+gFMBHWreIvneZHaStYNzvyvY3tqgPLDkCmjM5M3
uQhBKFdryXWwDpvL9gbGDtne/XemHL/jUcrdyIr9nfclL6aI+V6gubfGHpQT14kf
dmlLt2/Zhs0xgsK46R9Z0Sle6kczPIDb6wwmKsk7YT2YxlrAbK7j2d8VPvnzz6YZ
W2Ztq2ZFHwkgHhLk0u6kUffI+r7MbIrwmrznrW6NtF24JzW0lRRjqFp8NG29ZGFx
karEg0vtmZtzMFSj+1n6EDvAj+j/j4QOBorSOO4VtZZwSz3LHOihdNlMa3KMswfW
53GDmQlpXec87ywTrEfuEPz9ycYNtu5Gm4Y/RgFGh0jh3+jsJG/l4GaQdbbnLZ8C
y4yFuVIcoH6of7UOHoz91Pzy3tizBh/hk3K8P6D3Xvq6itBkEXnz8E/F1fOI53PY
aMmmNLCuYw6+9so+WLS80QrGGUYpBNjp4kftLw5n6uN0/ZYqlEjX4P6PNQl1ebuh
L03n+T/BCGUvVopyRgJAcqQt6qXdbRhtFaIt97IaBBscYoRqjPeCIqZPWwZj+bH9
0Qt4ViKkzx2Q9IScEci343mGzvXdQ/A42UNaKWVvJ96hfh1Fy0iWMqqmIKam/yNp
/rLNI0N3Jx3lCc+eDXAd1247OzyQJFmfQ1S8lORA6LrGkmL5iCynOWx988QEqSEC
rlVNNw7XUFpQVbZhfnpk+drh2Di1yJwVJbFULAfjwnzW8cR0AX3fTLsRvWcnbeAe
JaGkrNRcMozY9BiwKFg3/KC5NCaWbN1wBAbDTjaQK/BjW8KcF9/PjkBYGZ1xcrH5
ooBIPO2wr2eJn7OKu5y+5pbMI+SzNeaKMKB4JQak/daLTgFrEOGY9wwFHgrFVm7q
NGx+y9aHw5fD6mkkodgFcC1gzz8Q21oxrbn2dcUk8BxBp9lm2Nn12SHLdUHuzhvd
9ceEZtpymGVxkALgN5x+m0p3QokZrgrtzZxnefJCkU5+tsPYL5ZRGJH+ZozyrFy3
tiSuZb3zrhemAc/mh3o+z60oSayVWVM+NOTYw4qxoGTUYILl3/vfn3SWF6i1EEMI
ad5kfM+NK6/fxAHnbv0Z3lkyG1EN9qQp0i7sWIJDA77il7U5sY1PFp596GvLDmy5
8ezLBrXep2mUHi4Hd6voP6Rb0mKO0gTI+fQmP5TpDuFUuydy4x0g0VFiIMzhbedf
snQMsDcXwHhfX0/KbF98jxj79YrTy6kkWTcMOrKMxRwtdYIXr5fQinUT+/SMKj6i
nu/pENN5Oj0pdVBPs6oaNuffcCcOFvQeyrI+3FDNNiHLaycfpErWZY/t/SWZxyuE
QKRF2O3+yanCP2KcEp3U3PC1h/NmxPR75tZ+CZxjWVrRVk5a2cKIeMqChtN4aoXw
psJOi8Fhmrr+885w4ZvVkhrYnXCsul0niAyYvXQ09tLfvY/1WJ3DunPPeYj0SPL4
i7fLm5PcmHIe+gYWN+dSo2VaAy9PuSamtBRhUzNqs2mCOcVfyvczvp677+vmJ+DC
3q0Ki1/Wy3lN0Xq+f7H4j59yJpSD30f+4CaxKS/k2jE4CgJu6Xb5yOpMsikZd26v
H/tAANH6hJPsXGi1S+xL1bHiJ00kmfhLWpgirgOJtUX7URgQCZLp9gLXMr/w0SaD
/YKZkvfpZJJ/zD0zMSYnui/0ImyrXHfewm2WwCTmVx4ULZQBloT/i07V4+bsF2aH
VrVKDWr2T2aylst4htRSN5745RbBkc5TmM+lVa8WxUMKYsOxIkNI5XXemwBMcyru
tuBmPuYSRsciv68c++wcKVnjvOZu433zxM2EWH8NL0GB1NP0m45YIsEm2xiti3ew
kycwAyxAfi871vYSSB93e1u2vAZdXL0JNR4JDrWfSj05azlFxT/Z4ERaVDO1j2eD
0bIR4yQPq+Z6s5z+Hr/dVsbXdjD/qwe7311HNR3n9YUV6NGtASqbUrnMgh7lQmRX
9pJjfeVYGYVPpAkVBwpFpui8FsULRCILrTiqPQglUtKTxGyaelLb0MlRb7/j2Nut
e7EhACSJD+uQFa0GWcoZVUf9NVv8p+6XP+fg1SZ2z5cCN5jYns+T4Dl5qeTr8Qxy
zP/irxkiOOPhn+5SY5XxEka40d2rB/wTPn27oK1O3BsqzFUgiZ08lKw3xyYzxUw2
XLODUDAK3ovKl7H8YH42H9MT98srSGwzYMj95CzAxZluhDIC0yt4Y+HoteQ4jitf
aS0ngDb9o1fNx3sWCoC9RIN8LWJrEjgddtV/KSR9VzPlO6wtLSYnHr/nxDo3z01o
8q2DPfKyS495bDZyEbaz8JNSeCjZcW3DX55heNGHtIjkKsenBrhJzXcIAeWjiRbD
RrCgtsC5MdwUpbNiUm+3rk5nTN/x22DDzwFTCeDTtI4EgewCpkPc1+rGqxI40zkz
tuAgSD2NHGcTrqV3+8me4TeZFzluEz+h6TaZpHGx3lp7arJXKM9nKCxcXSh1ITYS
Bu+a1bkvfsvwer+RYjIhxvCP97xcQYnK/MCai9IxRYqLNHuf08sseWvMtWQiwSCs
fIA/zSkYfsyxezT9jsyFpNULTKWodBgNFEfwMZ70q6x1PPieS1Wdt+HbFc9ta8CB
puaXYoakU0xeg2GVCG4qmD1mIkfm8nvaxVaf5Sy2qnlO1Qm/1i8EVETAmdiD3kem
xp9b0C+apb7g0mj/8th8y2OoJ8GvQvRgkYoJBunw5p0C1ZSWIFebqOQfAantDhvN
J7R72NoiPEp9So0MN2tSkk+j9LPIPkIJ1tLgY8GZCDC7zGiEOuOkUz/R7L5D05FO
bYxgyFvWi1p+h0L2MFLh1mWMqefex9LLIrRi2hJ900vCMd1Aj5n2N6vC/EKC4t0j
1PQ9mCe/IH68l39hv+eBzLcb2+BiC2AZ5ZqonJ5ULVONMoPRgNgqUrVcBYLsmLDV
Qf3yOKaMkNdWJrdt03QQ7ACYe80CBfQ4xn7V/m9opHKmnrk/AZq1EomCxTQjJkVi
/YogIXIdn9WhN846n7sEgClZ7SJr4MQTuldVBg0Z0uSduirwyGmfM8xDCS7Et1kW
06/n42nrunXxxNMSV79vWxOYpkLHRtme35hvGyxNYCEb92FHb7ks0DKYvVwZ9mAV
6owQfINVPuY9TSlESjfgKwNYhxQ8ZSKlPJ1o2PqASkA9mFk2G7R1ITd6OJoHI8p1
Ap7iL+bpP0Zmj51yqi4T/aKA/4n6WI6r0BwmTpbXOxRrzd5JNPBYVaslKQp6TiL4
9PuNqe/uys9YyzabNjecGsvo93Es20JwGCBacnOZewyhzEmi8SFmRv7PcwfZykTq
wUFFmgq5rHNwi7ZLM16TMlFqicXiZXZDjpONj1pTXCYSpZtJZwuTCkgqL7mHKQW/
CBqVExfljk00qRt9xxs9AZ9e4z8oTdMUuXIblck4RDSt1LD8yOE4cC6ArJD8HbVl
R23HPdwuv9MVPt6LioNCgmbDAgolLrFTUEflcb+WzZx4MLy3X4PWS+yyPt4qxbGi
nez3GgaphHrwJQRV4Wdqa+EARmrASheRyf96e81mY6IsowQL3IfyVeO1NA6EEqjJ
17RIqS6lYbmlYvHczltDrKVJ/B5ClOqApSC6HGJmrAOUZoYjMujo0EwZiMFWFgON
xKjlpV3wk8sMEs8oPHMKNHoXEzSkepxpgsoHvBrIJCmIKFlUBsEOYgDL+D1cY9nt
Y8ruwJ3YIaNf8ytKuHYLD5KIEBXg3RYw6+rw1oy4F1vnwEiaGkgorKXno4Ea89E9
xlitI8ccD6P2bcRktITH3xSg+ScFblVJKxACFbrqkDMNhZ3wQLupiv+Wx5nxmkvw
/dP9RNKgkh4i6Rw+8qb6JT3XCV1f0djDzwdc1wlGH1NWU7pY1o6JnKVPXQcznKZj
5+ezrVqqDGncsSwT9tcDK/H/RSYeJvb+iawmiXjYZZi9OHqbRAYHbGAJqBdMBzIl
9MJ68igX4gmWK2IhWq0SWSJ8lNs4sBhfzTBz3doI3DBRvVvAH8Uv3Aq1OrGy8pA7
VLlxr2vI1dnNetIeCJ+MTgfsNQ+kqwG91fX0RvsyYxg10U/2n7+Qd/oAPpavR73U
BVkBKlijUD8VI9nvW0KOnrJh1p+9UXev3blH55WNKjNKB4cXeZRObI9Rptny8mv6
+giTc1pQu7Nknknb6I/ST2KbqxkbnDsBsfk7p0RR7CZbhUwlMu6ha5aEGlxxcKNU
ZG9c3VWEVILxwjaw7mbJuBFblQDI0usguErx9eUjxRVbQexvdVhZMxSjI5AP0fA/
PFSzDb7i5GAcoipXXFgWdpFq/ZI/vVrq4jTIpgNeUZZH5R/LthbOk+qE+wY5WK5t
pVccyTjD+fEvklagw7S1X+csen0Cr9FDiUwsWs0JKgZz9tJbLGLaVrlb9T8euWgz
GFmMKk/QGZuFvC3CEqDXHoaGchzax8QL39+UCtY8+mwTAsCa7LF4to/lk+R2qmPq
a3dinTCRsG6LV7taESF+3hgE4o4la302iWEmbJP5Abc1S4cOzK/e68Lr8M9x/l2c
Oprnulmf3LvrOTBpfiw6SUDyeWDZGj75uTDpZtiQwW85lEGmrmIIIVKiCncQcmzy
tTPeku7MhoQ1Kx6kOT5RNvmEUE0JhRFC5kSssZns7Whg9FjMEfztSrrzDqB6gwSH
thnDKQyNleSUoL0XS0VjxncV0q8Ayfu5gJRMtNSeleZDkI9W5DAH/QwgqbWbAl2k
HsUcf473dMjvm62Y2+85Dap+RAMpiXpzdreKda9dLdiDqrguQZsxo7y1+Wac8nmV
eHgYcC4Q2WCb0mFb/nFPl3Rb54faT/MHq3xD5k+BNoZedSId0BxTBCTbaw4ziLjX
xhHz/qJ6qZulxToygvIBO5l4hmja2IWel7bl1RNH6j8wWeXhvAlHDo70XIipwPvB
iInHfprWUbz3MGVs1C933Q7P71FQ9XZITlACS28Q/Hk8gMX6wYMXN18pdu5zgRTX
SgnNiFl3/hxwxjgYySGVecmoNDooC8qIARFA3DfT88h82Eb+mWJ4m0/kqdHz+gH5
Ue6iSrSm0eS2lRdtR1QFTUy/dWPIWikaGQO1fAV+kIMSfBVEdMkWyLnvWE0K/iMv
Os9dgSfQuL9+BDY/22yH26W3HzmtTYkl4DzFX1Uit6maCZU6SOo8e9dD+2h/+1Wk
XsQBfZ4yFE1xAAVWIe3/iND5Y8mFCFvZifgPqN0OeTHW+uVDAebRfDQz7IxbddlK
Cyq5HKBwwaTJhnYxNdP3A4TwYoWd3+KCwfChd6ew6Mdxaq1GQisYenHxhorp0bq+
0RfVWlVcsmnulcPEybTlwUx5gs5RI31QiR5IowFHZgp8gSxnl4+BcHyHI+ukh6ly
Ms/rNja1BSHRioBI6HBfDHojB8aciiy+I0Uva4T7X26V/pwuRIfj09rRDc/bH73Q
yjCsTWTOfwMdhnpBIAq38QBvLUhQ2WufaEXSKwktIqpcVExfne956I9W4UlIHbYT
tgh4dFZy2BmTqPfR5ntgWbgiug/1QRvKqahDmdI3+zrGmu4FBZSL1KGdUbZTefO1
nzKouqTCQqMcTqVD4iizVkr90Ci8/8Qrk/BHSZx6l1lhzm8ONJCFZMSPf4eU1Feo
yUg2gv0WUpA33y90dwYRz4r16PepH9qA0db3Kh5NyFC6sMLfmLT6MQM9rNAe0yFs
rtBkXyeaish3gx1u3SFRD2tu0gCF6sLsm5E7V1euY3AhcHBqf9qfV4bznKlhqFlS
akyfExfzoJh13YO31sZ4gJLNicXH13prxEs2lkyHELZya2Jb5iU8WI7+DEav0Nor
Rc0SfgunidlKyRvxILJs1C0p2TqGmXRJx1aikKpBOXSMGfX6Yru6FrhwKROhP5TH
RLBBgwJ7Q3cueM99LDFxuJ+f9DPbqzR0OGTJyD1sKwdN53t7beR71dmj2XxRWPZt
hHmHTGIEtoTKx2aqtzW7rZphvvicyl4NKPGjGyWTiH2a/kozy5PIV5EYMazR+31H
s7aazbCNAHfZBgrR34bDiAWgzuVEWupD32M6IvVNIveKFSevC/EOwnKpGOl4ETLd
oDi4s10CG4OMcm7ahjBIfaKQgugXTnKe2q8Bom8fB4MC/2rA5Poui6pLVEs7AY5L
5EB4tQ17PONNRQAJzPailBqkOZGbrVNYt/TTEt41dnk8Hwt+PLHiyLnu6zuLrTJl
VMzxaJbFMrpJnK1JDoRduXmdOUeVGKphzzWgnVqPIigYXndYeXS2XkZB80wx2wdK
eyYu7PYrYefIuZmuvN8tmBdOHvymgTnGTFcxqhkhfuHe9EEoGm2IlXHPnLWJZ28N
8Sp9+jNxfkA9MyNIHdHoD5+BtrZES/GNT325S9hVbbnMxlT1hJWWou8a/CJv8nJj
HVkMPBxmsiNTzFCe+yfGmbmv32PMEGpsfszoutERVyoo+nvuP0PF+KQEc9Ryrxiy
KXltfQpWnsDTTGnI6K7YckxYxleHboJV10+7EedpalFWsP4VQHCEVQGoa3scKv00
Nc9YytBptAdN2lW8WaqEbr+eWhmBhW5t1I3wA0ZZur46jck/KrxF0mgQrVhqwWAP
46yqbT175fRQPyN57oQh0bMxbmbE7Y4xlZ66F5ORhdkrhye1n2/qqqSN8Lhg44A5
8Ur4CWi8dzgGBp24+sh9R00pX9pww6ACkrwsElOT6G/CiNUchAWtMrMU0TgeCYo5
A0FttcFtLRofYkNjWqwnfWR3cvRqUPzQNOLYKDq1BI8Jvme3Y7E2/Y6S97e9JSNF
gH0PvbBj3+fPV8jeCLUWNhJTB854wtNiqfBtq/nbgMEQjF9DIwM2ZR9PkdCAZT/Z
13GuhhI8gPICdW1vd9SEwz4S+0Eh5EMYvkYRzUkxY4XQ/whADHxlgWZI3yd+6+yU
zVcZBXD/2fFD5o9zfq8c310/ekvatof5WCUZ/SiikN7/GiEpDCDb+kHAL+ns7ykv
ngsxsrypn/CjoDFxTseDvvEej31nzyjG6OoZyt3Zs1X5STlYeRenmYbn5miPNvme
U5r2wCc0CnvjS5KSzlPZjgYoPNTQSd27n9KudaNzWSALmakNpW8+SmDLKuewNEyy
pf6Wo0kilJeYleI1AoemtNiNFD5qw5wD39OSlrCfiJj0aFy5QylDcoBZY83RnvmY
fT4YHVs7ZrWr15Vf255P02Jn8UPlqHt7oDoH+I5FnFfw1n2x7+nc1KzcwMWchJWJ
7T03fS1Fz2XlCQl9G70kBCwa8bcYCJ2yucutyrWAZm9uGo4b+Jibb10rL5Sfjk1Z
o1JzOrLiPSICJyRdpDHq7Zzvg1P5ydkal00uZyAUKRp3aE9hpVyFMMkrDhVlZHBN
yED4gQGeWoNP4wPceFGHcN1rTy7d08yJGJAdB3EmACeqZFK1GjTZaJZrCBwM6AI5
p7ph+UWRgeoOR/mZvNa7rryTz62l8pUiZ6aX8I5nU3AyWT07icz1CuD1qgMs3rq3
YIXwZI7k4GeCGt72ZI9kL7D9TUgVHWLvNTDlqPSvb9+rqF5YA0IB9pT1ck8JRFGB
sAp5ojrcDD0FL1XzZXP8otn0GVVZ2pbcOc+ip6RcsHYOPl1gvVKq5RRupxzt1TDa
xCddrInh4WrTA6i1OlvnqItx31LIwhIHbEp7UvOJIB0x4YDoHNHGW6FDaYkA+qUI
Go/Pk6TwF/eCfCUvD2nuCR5Gv2cBJTV/G7CySIfGu6/fGTmiEhjKvXANDva7wQMV
g8aZs9hl182J2pMPcU2bhHhntChm53qNMU8xKhMMx5Wvky/hIvdJD776lOd/GrEe
zX24ZYh5vFR3QKJRbgKlIxL9OyYfuDbKyptHfYeLHODxqaMWWhouKkxkXKdRKD6T
tokxSdfCFF0hehj3BPK2PprvMH96pcdBMPZyUTyUD1iG3604mMYICpHNheQ2tV1d
kdQe0VjzkQIWDtyIidCYLxMmUnk6PF0P8dZkTJsePowjEzEK8bGLzTQEtHmeqOol
8TjUACSTyGjDv962HiccWXuh+1xOrZWMBVDLWYVQdLq5YWTbGvF5Cs1RdcRv+InC
yQPWMey9hJ0trPF7vTYmMjiSx3HgBrVa8YfKVbrKqQXh2dRkoW8029uJAxOTRz+7
M5wyzheYk7jMIPKkbMs3SWsmrn5lQBCvCWYkxXDcrlSSXBWOEYGGoCn6ck8SVq3D
fBrCj+b2OVXgvzWND/Acn2tIXcyjnwcOTrN2QPn1HUY1NaXGFVGpSwngfIcbaw6Q
/cLsJt6IPfO8RQ0w+jExO6j2dfliHbSxsAz/KagI1DYVBacdeA5oeiUja1cws2kC
iDJ45hQzJovl54Le/dqosPyQuSxJOVNUjmvTBbnEEELgxy7pTrL/wMVCg1QzTmAQ
nQfuKiahhKi7mn+HavB+C7X8Yp0tXuvJ9IeQq8MIcKxa3Q9sM7cVVvDXoIP7v5lJ
5od2P1tj4oGi+NH1c7Tvd1KoYMWZfFkg5i/aIYenAEFtajGJ57eVnnjTFwhLzr+P
5JOHxC89GVwGqQl2uUOkaa3WRbu9Ihs3oroWbCfoRBDLyfggqMbOfmMeSGMmpBj2
ph2y1BfRu8H9VD3sJNsgSAYUBn+nGFEONpy4ZHlK7k/GDloZaKyFeku827nlInGg
3Mgju5x3fVdZ05jlNwp5YJPGGPxmMvwvDz+6Hg17tam2BpyBzIGTU1NntVacfNCD
X1R5sUV5H0XrhGTYJPtiUR062JfdoywUCi+gGeKHiTpih0v1iVMrXIO1oa8zcf2S
PTIbdzBVP+RgMqBm67ueMuqQzJQJ1ZVHO6IKvyj22RFmiUssgZbbY6jvwdTLjNk1
2ZkwhyNvhKojGigkTSKNFk66baY+d6eFsFpZ/v8dRtn86KUxl5ZDqqomBtXI9Yhx
aUv/46NoapBbuDANFROaanT05pV3YCQjBfd6XoPPH8wtqdunsB7YDCBSmTBeDunl
RE34AvDyU6zxFmSwScH4G010EkYxvSSHPWTjPo38P6wXU7+xw7KAJDbhQYzb+qr3
+j59yMCD8OZOzoguBVa/ME8UiuBBf+EiQo14ECYHVJih/m0c8HeESzSHMyv+4mLG
Bqj+CdySAPJjQUEiT3AF9420od15p0+bG3oSjFclRu9GXkdQOp/70i1hzqeO3bqK
QUuru1nUItFFLw5wiXqXKNoV/5D9yiXvcS9uw2kcmnpM1OSW4RKiNVBhlIcbVGIB
OifemhScD8eThO6WX/3CNN5Yv5byDYWqsICtjOAml3YRTVOyaa5HqY5Y3Cf7tKVS
6QYNKzZefTVz1Usc8F12vhIgsqygAjDxKNi1vaydRRfhL8+IkeAPFoQgkz6Ff1AV
S0x0KfFGiWCmTamALW7uGb9l8IbLEzAGwmMkyq8AFucJqV9Q61w5zFBEvZBBEgGJ
r7RNvmCsS7AOAjlxOnc8EIh2+h12onAgkeL3T8xh/bp4qNUUGcXZ67aIsOn0LkmA
5i3F36OQIIRmbGUNDjviYIiD39Y5JrtM9z5PSKCRaEGMKIvDPezwxqGANERIrh7w
Z6MoMXjl01ntz1AfP/Kk/qTOWwqmD+Bal5Mc400/Wr2YxJFvNc13/h7FOFf6NnNo
ZXAK9PHEqkENMjcGW9axhyWGBZKV+IqfxePs8/RNHcTKzBR4oJ6A84v1h8VEOojK
2d5DOFs3ntGu0Mbx6B4p02HxRT8NCAw7SKWocIXAb0n7730oiABAlkmpf5v5J5tx
Co3GbEFMjTz9FaHLesPtdTtwuZ+d+dTa0dsEg3F9ytI/+GZl2e3vO7mK+CNFGWbU
z0gNRGzcNuZx/IzhRKdEso692D9K3jAoKeFXwEuSP2u/NxXLrCxq5sUvzcfDwn7e
fiZn8FqfbOEC6gHr1Rh9hv8U8cjY9XZ7nuyUwVOxSf0yeWR/rxjhg6WkSJV5TIrv
BEeq74DmUUmFXwPwuUtnNBsx606j1UnOb1jyH7LCibyVnBNHhojP/1fwRBpDaGNq
B9wL559+po6FpWNkyn0WUcvKqYpooOPreA7YOgMXDreWWavKrjjsrNQUTgagh81a
hVvBrIjrItLZTo00x0KesZLGLG8XdnwX73RsTxpjlqEYJZNEH89xRVrMdkKXZsFf
oPb29ly+7bDkrgI+FNz01HOwRdWb38W38lV0aAYxutxsZmxalMGEerl8nNLQqZ6h
ynL5TQ3LOowmk4oasq/cRRnvPZt+vnvA53L/Gu3vwg7YG8CQSUf5uFsszUMSQHnv
exu4IRHKzHlNgBXL8YnV38eWlInsUlGbwmbFq2fMLMyTINFOwT00omg+CDYsWgtA
l3eQrb5D4ox8TZHrXWpRz5pCdCnv2sGf/MMOiaiaYizHhQK94kH1yqaWTQd+O7Ls
NfL353WoMekktNKy+bf86fIzJzvLoSjFTot4r8S265Nv+u+fjB75X6M1apF9i2E9
dqCdz6SDooDHvLihFVaya9f4JuZ8VUWUBAu5kBw91Xjrf3NsM84jYrjwueYQOAE+
35dWVcGjQJXKPjcoWU2jKjl6dploslOxHUnOs8nWLBIVWXiMfZYMWNdsHLwSpCDs
YwWpvmzu4KjKm6ESRZ3l96phVH+qELtuHrjPhGQosarRS7hX6a6thT/gkTegADSX
osP9YukBUfF2wIuthEF/sFa3ttAJRJ/33NXb2BQ42Nf1TGfqKamEUMO47CafBRH9
sao4Q/AWrcm5vaK9qh9LK3TwmA7pVcLLFyDnRNhmiIwR+aA8D5CwvoHVWNXYeN+A
8QItpOe4Qjs9GiHHMJcTPi+2VWaZPrp/8b2XY3k5fjs6x37UroFYjflxtHRtREZ1
ahDdSuiYl9TlgkiVLNtGz9t0w0iTwJAize4x10aRaHkqaAKK0l7AijTIcA+Y/ldB
rUZ8Q8aTrr0O3SboVbBptruw2Mx3LcMsejTzo8nvcmOEsDIG4ZynhTvPs1ucTNfB
rlPImc92zqN8VQ0oIV/fntZdbWTvw7Kr1H6s8uGDv/U/0UFKlhB2d9tSdjW884An
IjvTppnFaDPEX4x19gvNEFlj3oZ4yyn9VlV50HeGp74wFfeQtFt8KYZCH3WvaCQR
Qvv+n0uhOHSEgFKMJQs9dcFft0+3UXbd0MM2+fyPs17kSyoDzXf9nhk7+4ef+aXx
h6WOIF1cnfiCJ0yciW539yu3IagYpguSV4xiB08D3icPtF7KOQzdrgXW6KMuIKoR
lDYo9DEN+k5YBnKiaUdxL6p8s6ykwuEfBvV/FYOA10Zwux1w217UNjerQX08WKue
JPwcRMU0rS7jf5mkvJdlnsoLi0pebEyMOA3eHjoPU4j0+zxuVpMeWo0SjMVY/jpI
0XhfEh6FT6OFbX//+8Bxx6ACkxMQyhGpqglgRSM6pmA1E+r08ztb5jb2SgyleRg6
q/RPulj3sJ5Pm88FJal2EY8QZBENqTCCbWyOHVtcR3owI7i3OtOTdaS50192nmGm
MtBKkBUDWRpJxvLLDRMRVeaIeYSqTZOvxQuTUYZZmCtqiaXHlD2r0LgLuYAWdi1l
bE1hO3BS/B45si0C638OTAl5zPqEMfkbs3Gx+NPTmXajKxAOv9PwKjFcxRDeW63l
kYKdPpI+VkxgZbJnGYNTa5pEmJUXT+7AC4Ke7X2l4Ix0XwmaP6V5YDeDGPmkOc6f
jLFem3YZdkWfzbEZurHslUlVamyI3F1Mg4vZRHjJbek8XyFhgLU7QR98YAcHic/x
yDv9D6wfpCPQNPa+3LkmOT8Ji1OclaZbYw6F4VGgnpfvXIOgsrwUUwiyseW3RIfN
7HOiZ6izQ6Ad5J/DBm3zQq4FukFioepviD12eWYudn23+Si8Txpt+N1PPm8nL6Ew
Vvj+Baq+mjdhDyET1r25TX0VIEfsdzhIlM1VBaSOmKrObH3byfPhCIfX2vgLEiyj
rTBTqhnNysMMgkB4o/dTUrPSL5fPiT5w9Bdz/RKpm4uCiFdLJiLDt8QWqlpqwaaJ
148CRaw7cbA8mVb8zUjouDEbQR5vAqofZBjwVUWBfKa0wuh88jkiAzBSaqRwxlRf
jxUci25KGql9R4jgLxFL3V0M/PPoJTC6T1/AH7O3PCY2MeaxF3UnMmlg954+kQP9
BJ1J0+i+jFt5UgotFdIhsb4tJ03vp9Ge4SFMkmfmi2IBngSW9jjPU2wFwaCWxU4L
kkYCfhX6M5Hu8Psk6EcZOCc9zw+W7vD1uar1R9Xlm+LzLGmV3PP9DxeyJBrLcB7o
Cph96cFEuGpg2J+2DATe86Slrv5c2pItqC4+UKVLsECNlYJf4zXAcCTIIB2n7MgC
jW6PzCUkmH/hYQYbPj4ptzkFVJ36uyWAD5JGpBpoaWRO1rKL1BO9w71YAShEYnXr
sdUZevbfkh+o/3WCOSiMNvCJwk9I5VZLlJZ+rxQuIgEg95FDGOnnhYzxUtKqtaaY
dbqM4OiQPHWAQK4722eTptXzh8AdQG3xwHhvKzhO3WDBGpSvkqtbkhmTGtE49RIw
8GLEqCqgksyGBhYHIrFkQA7867mb1jtgCNrh9TXjK7xUyTT+/Iw3ocBleCiNCUFU
VlyjZr6c5bbamzR7NvAdbIdkLDW7V+6Nwn8Vw6iQ7hq7SVM5j21vNM8UHLQtxm92
sNzGQHR+o3I1sL7G+PhpRCsZJtXPNGSSUvOFp0Hf4XhLnqTV977MzC58MZtwH2P0
ojDxfrGPn+i9s84NCnLh2aO68IRgMT8LyLT6ckBtr0GxbPB+tzKcmqQ0uBUgBKLr
RIREs/94qe4LJGBy/E0FwI3qFNIzMvocCMk+laFFuu+9/ifqmRksYCmzvXn0wM8F
meBWSwfIj1r8w0hOuynreLapxmtvkm9D52z5GBe91SE4t3yIB4rKuYL3X5TNmtHl
dQpWhFiNM6f0PB5h9rf9tKLDhFmOExVctXZR6b9uOs1j6SFrXJdMg3laTBR7mQSJ
uuS/Mw0B1FB7b1CGgXe67McUieN7PR7/PeGo55fUnXv4kJslRvEIP8GX2cvIlSiv
P4E9m6LYeRz6tSpMrA7EQZtU4gNDHnK+NTmMs217ssILnbvAsWYoObrdhvW38zrW
Bx+z5EwyTGGA4DjxzCtrNmkc4WnzerXhawdpYY7/igjWJuTvAz908SmroFzAmTRw
F0jOOS6Nkia04/PVfyT2jRT5PGBtKGoeVCgdSLXLdheLS+7b9jVXfXxxpzMbfyEa
XCjr0/GlqiwBWuAum+8U5J2J5QOvp8O81F6E25bE9sQy59+cHKULmhOSZAEYWggI
GxhfWK87CyzdB78IJN/O4UOdfjNSuJYNG8tkbLSeHS6NcgBZSD3+EwEIN2pIuzie
mG7RuFnM/dS3nnjqyXike978t+hQ/eOtDv8Z0O9Xp6+FUW5qrAGIag9tZ0k3rJkt
D54XWEe3mWKvtFiAtXgzDs3kWYYkwDf2WEtySHS2W1okJlVe+U8DSm5pxtk1Chc4
F7Z0f7PotQiakxEA0C/vHBAPdCQJPgJu59UkeV+qUkyB/80jPpWa/ApytlhpZkTf
U2lDT6Sfe4PnGF1Kwlnflnq/yqs0J+AV135Lv3IwHrCOdh1PKN5SQCzEqisLsNWd
0fVcE/A+2zDCN8gh4R3O4cmvC2rllRjjD+TEbVNfHUwPigSLoNJLRo7/hNaxH+Wc
QtiuW8NIzaaZgmeeYG7s4nygf5hie4+XdyjaZasXSrR/pVB77k8ZGw9cizuRaG9o
k2u6Fa1DizsmJqBC9o/ZUFGGMjMN3zpnMIWamdEfueAscndwRoUst2vMa9NihrJX
OIzch70dtUVOJB6+dNxYR0CYQG+BhJWrT4E2V70lRDnfFpbcbZm6mjgEtZWc2xRC
I5Gz8W/3G6D5Oq2QIBYosvWyFksAbbDLVvfgN5HVonFmFIVWMxw4iltKw2aqWNZa
v/Xxi00ieaKdSQrssLCqCnqWlkMSDp2Sh7vH7fmX2kzaSj2mvlvVXFTXK3Oot0E7
JfUdz+BIXck6u2RK783msBoxYfc5rC/XGTxpsi6KAzURAg//Ff54pTXdXWTBzZRY
pPQSvUMGxZivYXZ5g3ZQ0CnNcRg/9bFDipWKwNpbk9F8v4HENWMKqhmsqIFxIOmj
FgL48yPlyfRtlBa32RX2ytzvFr++fcc2OI5Objcc4sA1IKG/GYKDAkp1/zwbrqvn
Mvdp4gPi+x0c5GgI++v6MN1eVIVPpRgnHBp8swaAQ1iO8Ckw80redBbW6s2gDK91
d2TeMskyL2YF4mw+MZuKwayt5MHo8ukhHna3rEiBmo8NxeELShDBF9+aO0bvU897
ZpbaoCyFttlb+F+iqKUahBAct51RcXqw3BRpaxCdFFKiOJlF6hQvCI23RVfohJJQ
pRSweMkgVAwy4gEYVExSmYmB/GJIeqWEovH8WfAvU/Q0OQRqx+Ze8nuzptsPnc9d
d9bTkbuJLYffkvh3c+7xyzVTEW6WBXfztUUwEGxEeuexKuohTI7ACopBFXCVpuj8
nQBVbIJwkPhtJOopnZS3Cpb/7CxhiODXngCy3lSLHpGS1oEF+9mHjCPB10E/60qS
XhfPYaViwjKIj3/LxfMlx/oxcNr3uOYqMmnvzhF3COh2aYTz7UcoHfX+8uM/LiXE
fDcWKM1f5N6+GToyDJWkx2oQOWf16tp3m1/s75MXL1VdQeeE5GXSsDYYO3A807jP
JlRgVPkWeNZq3RSkrRGoqHWBjy0zbH54vA4HncrQhIKUkTsyMpuW6oKHD1kjOz/2
EqhK0AM2SGU2d3kgJWEmLrFnXasZr4/SXm4TnZynIh6R7QJwvXe8WNq/I/k9CyNV
//YcdCkmHSmhB9dgSiICc3XEpyxgbXRrubLt2wNg1kZ71avg0glCS/BejocaN+D4
HmgngxT9YXoF4LC2vcdzBpBRbagClwN9eyaXSV93d1t3m4le0w2SZaSOMu2qGoCS
fWH24dsGEEJi9IPPQ2nYVwCug1IviLCSGnDGdMDkIC51YTaPx/aBVZ2VXW8dduwH
WodGZ2MT5yPVK5vPunsR8Ay6FtmCSpLBm9JKEqpI3PQozC2WtXOCtO3eKtSFPS16
ba9pLT+VvsFZ5RPiR7BMseCV2A41YIS7gmksu4ElWnMr2foC5PPoGAzUwPaE99wc
Pfro6/LFByJGwmB03+R8FRzclMl5/5IdCaIp8AiNd1DiC8TCCdQ8C8ML8K8w4Skg
HAJO/I8QSG5MpRkvwMHJQmKpmvTEpAmNLr+JcTCF0TPIo4QnCtXlvu4ED7OW94O6
ibX2gMmuDSyHJlZpxwUvqT0F67R+CS1JvZpGrbMrGzHA13B06KUFkxC02kzV2/ct
Y8UjFfD43+GqFXdIQi1Oc6pluLm0fcWYpwak/x+KbSNNPOj4MgYuNqz2m5elU4hg
GlXqF0xLZA0aIl/kve3+cdJiFyzex/ww8atkOptEZmSKrNnbFhNqqX3Ydhr3RSCB
RDXl6tBSAe70GjKNqRk0z3iVmZ8nuM0fV2iDR8eHAY5MZl/VGEhO7zE2qotfAmBq
2zmY3oHOAl6Lu4jrR2QNCBqKED+M5t++55reN0A3WHbTuE4vR7VhGFxXe6dU9s0/
YEuq6uS6D8t2DfQWU2q7PlGsccMOPVTLolMyShR50Ya+4/KpyAYPRtOfPl2CC2m6
2J7yJSj1csmR/813e72S88VUyX+W8A/d2QohHWnDeZ2qIHX5dvyiHORwRgsMFC75
obz6TjdRFUvzYURgknqn511malLTxISmrtz2Am2muosSOoPMKk6qJNEqdflSJEUk
ZVK5mS8CgQjYfy/a2uiR3ke0kDJZkp6MnMZ3UapFHpKJU47Wp0DI/mA9Vh0p5elK
zO+9uSQR06Mh5hkxUlN3cJ9uFd8D5ef3eyMPy62cnUuu0Gv+PupEkl1PkSRPke+X
6lvkAm8+1ZwuYxX/YLvJCcMcpmqCTPbrS0KA3lEG+Te/Xw9tpjDOn0eOfzmny0h/
Sw9RvPEFj3sjJ+MxDPdnmm2/JlBFsPC1p+O5qvITtFuyRS+du+wS4ntXF1HjIIvf
HI2a8DCPm2p5oZbICYqi5skz/h61XKpB+R6zR+6LbXBWKdL9DuhLOXpp62OoOPIn
pug6BFLKdoIf22AqfyBOMqV9I2847Mi9xs7rYQMxRGGWHusfQhWEv46PVX8wfikb
/VLR1rJ+wQtGdxL6KiqOXJqZhF8iIGhI/qeGjwVR8bFhrYM4oWjgUIN2rbloUHww
2rqzAq6M0/zDuOQviiBx77jpUAFCdNZ1QCP7U+ShYlhVDaUiM264yPDGbPUjNtSN
EqkIb6sxt6oezxuF5dcbx2EnbFj1qskqJJExxZPnSZ4IrT2dxrkfwqQ+glEuIYW+
kOExu0Mf2axImc6guvhD/LLsdWOwZSrnMMdslSEkm/rrKTFnJWcdsxyLsMVUlpy5
m7Hc+QC7LFR46iJcyGer2oltojOFVjRsroRs1UKYuei/N4chkaGBWPR1cZvbeyi9
X2LaJpoC0liA3S3245i8owJVjj3BZ894/HuUm4SX8+WA/UScn2aYAr74ZCYrdHmC
wJ22Ik0PRMqO3itSeoomZ33jIbyKTmVU4FqNwAmjEkrE3BL22Llvv/oaYVOQmwBU
pdgrIxr0L7coLJocl7nx8nAlJ3XsFcLqXoYIMe8aQToKxqqQMO7K8K1NcNt36KZG
AuVibjeMtaFnyg0yZaiU5V9t7WZlIRrr0lwNjNAFTorLnp17O/rSOwOsDIg3kXPp
QsVpzgdl008s6+raqafYiMt/dtLv0dLJb3xwLa4/Jd+45fvYU8FRkIP2RnlHGFm9
tdA0YcmDlipDCawyJvAJrqhVm65Re2/ud7AQURFo98Eiji/c7aW1/5EaukvYhKIH
OP2vRDXXecVCLR7+OlSCZIR0PjGlkA7WlcQdGFFlx4Q5O7ltA7+H64MBnOB5qi6k
Fj5U+bdRA5p8SRKHQCEjXFjHXHi9OVrJTgVkc1fLUVnOp9PN0PkuTfX4OkJwNeXk
BpTmbD+9eEmVPd+iVFYdufNHXEhYrqMUxAUtW9iL6KI6SxgGKFHPznIjqANBy1Zj
Sho9Y/PhfkoDCGoEGlU2LM8fA5AmguBm+YI1W2DmRBM0rujT1AYIPUDikTEaU/MU
XnMHaQxshF2l4s8bH6mv4FRQl17UX7BiJh3U3EiD5C2rHmBmdrZ5VYzr1wpVWk23
Vqp077gtT8cgCYoVg+/xvi8lzhDtDVwof0iwVvnrji61xKhfc/C+3aE9AR6KLiSZ
/uU4YjpQo270oRgDgHWFR6zEICkYHBSK/zGTz7HR3ZrYy1EP1W3XrXzmSmuLhTZB
HwT8u62azToEoBBZofuFtCM6A27gkQ0+7+lPgc761K+ocxRzSXL1O0VGf0HBVpKu
K82cJdr7kWD78mUKZENuAhH1KcCYYupSe4Jhohe61AIqXs7cRz0YFwDxVJS32seK
qLJKb5Uwsx6928Rv2Sj8rN5Qihp9dp7H0Ygk+3Ff9wSB/HC30Qv1YqPp4YzDBO8o
Fxf8LZRD+hho7g7kr8uvIH11VfBVN5qK2Pxzb1FZmhtQe+EHBJWT+/xNEX3VVNb2
fG410nlyqFVDGxsLQ45emXUN/6R9Cpn7YdSPC9jfCTGJu/fBexJ9FwT4m5QTsJyv
GG3JQL/fMxWvcBNdKUQh0e/FRctVZjbFVe+36+bbQysZOCFp+79eXL9ihMSUA6e0
rxTduiMpzaGGuewfQz8JgOVzN32S5rIgOLX8tF4WzGs0zSr3orV+NVnX07uNdNce
hthH2ijJGZgGXHXtcNVy7rmT3OEIrffKHu+heLpV+JlkwR+pZgvQIFCKTKtsQ/ma
F3OeuTJjrvF+1X3lK9T+gU2lUjd/+EBHqtkZzAtpnj9/MFJEaYBZ3X0DAn7JP9q9
jcdtCqu8+HeugiAtdnHBsV5c0glSe3i0OHbuwtjnN8GedUM5FqGOl3XnJrJpLV5A
iseBlT+V75pEB9Uqd69n3T9STou6ykMBj/vdP1rAeJJ/qirMefLFhkkx/uXjeC8f
EWdnryd5RabsHkXzSv4h7xd6RwvOu/DeuKOXhKgnQeSQuw+lbdcy5qnDGEL8UHpt
02OYiz0TzFj8mMTU610+nmlszSegumGtHuS1W1Ae4zxBIfuHgPQ3A0/eD1NvYkc3
4/NjxnkglSSMNudvMXV3egCnxk64IBDVMFmreri1SdDrC4Ntdrv52U0gj4ha0dna
9m0QjbMLufRyGBQRP3KHbx3kqqF6vl+6t/9DN4ITjxgo2tKLvJlWfAu7bQiM+EOo
aj8zgeFQliV4bD9x4yjkzLPR39hlvklvVxQGFFpFsISf6VtsEBzv5iPe4NuOqJHf
FAY3BVCdibORvNkke/dlv2zSm6X8K9GpTqXJDnptfk2VkI3RRQtfC7fowZkVfO8m
gu7nB45SFHPU14DehAhGuYYy1YYDhEqwjAo/HsnCSuJ6PEAvv5NDbJEIvlFaLqxo
D7VPmrEiTioAbgXdEIGjn+nGH+G0fYQ75u6nBCnT9wywP2Bu3mLSPXXDBLTeBzNY
mtapfmF4+6QrfRlhoBaES0clN72VP7Rt1Bgek54qdM5Vg5HcSOwxrMsxvfzig9IV
+2Ml1CPRklT1JcNilPhqjWaYc/Ej6hLmwhF7Q2OmqPk/Dwm+eJty/qnRHnLM+rjX
mCg4cWl5nNHv18ntchBNOiBA+s8FPpjy5jJ690XKla60vyt/DseAbQ6JQOLwEAB/
9u++UH3AGYCd+4eJ/1tt7wIJEO2TYmrMrIavHNmA5o6cLADLIXjEF3KB+IlCl+8G
tQqBS63YTlw+BExVLDr4P8IwhU6oaljKJkcEXzpcLa3rXTrfH2/YiRCJaKkJki1R
ulhEHwDJGyl6Q1IoTJiTO/kDc6pqZLtUTHvrmzVlDK8q60jeTnZ9cv2JlyqVrTXr
FlZE5hcf7BaoGbbfcKtc2QJnduBu6CnrS9JYdwL6ChZVN+KxJ4/T+gmzmPAiu7CR
h0HdTJFkqkT2CEEo9XYI2NSnP8Vo+drHaBeKQ1RyJsCMxvONelHijCCvUoPWLutK
DpQG72MvjWb/rg4BeWru2HpPtRWdyuSgKQOmYlH4VPR4jdL5GoOB9gad9x+abXcU
zXDZ1VgLOT7523GM5DVqrv1B3nyF4U98OgEH4KJiILkN9rwILw/Lu5Lu8yWH8Oxq
wFmgsOoYIsOXKhOIkB3Q31JOsyrG7zOFq3BotelYQkPQtMZ/EwYcJt/2i9FYUhbP
YXEAGb9wnrs+/bjOTngvwIU3dxfOIaLyddvMPfPL7w5rC21CmkCfhzIhKqEJiwI9
uCyijO0BdmoNSePhApuMu4nXKstmnMtFfPFKx1li7k/+Gvc4sFayvKW2MIXPY+YQ
E0jzAab35w+TYgcsKltVOpDoAAJKK1oc9Vk0h19AwrZKV+2VE7frpK7DXWC/GGen
ShTQ/r685pxcHrqQSi0WvnXXkitmvdNl/X1R/lTQe3iUtmX2awlUXQc5ZBgSgFD1
KR6sCAGwWtuYDxVi7mC+8VjcrT+efjzNtv13+33/Buqo9kIwnusLTMK/2ZhX7Aig
ybEF7EYN7jbXZA1rlaMFLu1r08pVJ/KUSshepK7bg/FkcubC4Ekz3RbX3/NkaEZu
f9V0NRbsWGm9KgE3qM1D8hwJVWr//DSRLD6X8RTKQF5jfyNjFHSrwWhSncOjWiKx
h4BBRmjyyTvIBRlkl9J05eaeWiINT2fRVJV0+i93gYC7KZy55eq/b/g05bjdK4WY
dgYmro+Zz8DPgq4c9u9V6CJvqsBQX2jTCovdYAV4Z9q0DvnvTRahmaNSUIzuozpt
sOO1/TEcXuHXNMpQd6RNrOEr/CBsInRi493gd7K+e7ddy+Gcjn/UNfkZkOPvlibT
h63t7THPcWYvUOwKqt2p2Jv4tuSrTbfAR9gfV3EiwfZvGcnGUS6NiqKI4Hx7bYFt
EPiesvMYlNYjk/zzM5/khxoIgggczwMxd4QDKG8m8zr0P7pGNNnwJ6Gyecw/IUM8
wvf6to72dpFmKxKQRqv1GU1J8S6LS1Xq1v9KA3une1Rf9GzWzIUqi92BK7jtMaNa
FreJdow7vPMDPuTinfW/ZvS7fCc0uDiPg3N1vnS6cS6oiWF7SBuTawI2w0bN3mVU
OWEH1JjiJ/uPHVHu2cEjtAw0HHPC9tkUXlMehEcO02gQK+caqLh1RsMoXGByC4Jo
yVLeV7bTe98nhjR7kIUQrw1jiWquODmJ980VRkjj2kRE2L4x5ASNqNO6EIJsXtvv
vvmZn6HCqX2EacfxbKfRUwRNBQ1BjXJYisRZlZ1hpsS/bIIJLEBSDEJ6mbJ3P4N1
AWn22pLMWa76n1BeRO9rN1X0BPWTkrFc+REeb6aPriEHhFc6XrzpzgqXkFTZgRQi
y5cSE41e4WI6f/pr+tPBK66Sn/il0Oeo5gSZCtATpRF9v2jJtzZQRDaih9RmNtE2
tN1fTXBwf2td0I+Pvt9CJv6kjSdA8hjNg7CulRxQipKD97dkqqADlxWId9Mj+Nwf
GCJBCnE5F7O3maC9DxDuub7HD3glyrl45+dnLYCC+wpZTR1NxKJGwwoeIkUWAVwy
Bbwn4GsiNS9mxiIP+NPrGSlU9xP/ycTRkOIh4X4I1D9cVe8p11AGkV4viy31HxFp
sqJmel9yTc5M2vv7zbcv8XlWyAeioFkKWuV575t+6OvJDknWv3gHQBusqH+06rdq
2ysFccmSOwIy4Jc3/4kj/QFB5fKIL3129PrXuKGSvvOHzTuqcFj/9m394XqRvCaN
gXDGilJR1dhyZQDeo1kOoPvQAiVsfzZha/InFMskLuTg56R8tBBefsndWI1axKvP
6AuPG90a+dfn7KdUs5JD5C3atX+yVGKvlonJGsXJyJuJsatcbBBmPsOyObJA337k
14EFSAgiE/wpeUH4vk/1jazq3HOWUpiNsHbEdQW5FRp7zqZtMBu7oYl1FofBN2Jm
QsjA2/0UPUyYzbMlD4W5lVAUzjsUyTW8n3uUSmrzkFDkH9oMwAcy24e5xAWCGWoc
qXygZrxjJWgbHGMoz5/RM2wou/o1NOtYO4ypV/xqidJOLu+qnERMLO/2sFPRsr+Z
1FHCQOKmti9/oRRzMzuDSjZuz6BujaKHLiqTzUzVotc1o6V7S4eAdONOJzyvhtiw
z+dW7GQsg6qB1zx702atagD2nLOQXuf5HL857HL0jpq1FVFtafreVtHGcDY3nZws
b/X9c5tT2WPLtci9d1nXwXwC/ruuH20xBN9ZDUbWnlci+p+CRyJjZSgVHPgpzlrD
X1/QmI2W/Qyw0W3O4dDcXxe2SeBIkDgQ5BMCIMj/lpA5n+z86z+hQ6LjDaR9IA7S
7Lj1onlhpMIE8kSPwF7DskOdSMMLRFVPhWC66TZ7lWnI8EVsfrz6TZ5ghlzPi7DE
wfD/BhlfVXFN+loVRVZ+F7KVJifejO7fBKod7fFsW/JWLkaarInTT5bhCdhYZQxF
H6GnRKu80vx/0uJ6pwKrsGPG6LBg10ibBAT2ftfmGVhuYXBcusyWRi5iMmUrURas
L2xtkUVWjULNB4I7llcPQONG2K9thzqCjEqSIEj2B1z355PL6U+kaqIcHS4QXaFm
FWwFRxOWLAXg7tdpIgtvoRbRQM/IzAwaBNigq7t3KmYIUCWK3jmm88QMdwb+uq+X
JEtZ82yw5K8EUruRk05UsuW/9jbwBHgdXhHdIAiciuQQnhkHZwsHygHqmX5PlRHG
3iVEwnNjyndmPKTn14vg5bz64tWeQBasn+e0AvVlx9aT//TysK+r5EJNELULNpPm
J+06EWFK7Us/7rAC9e7YI5VaX+x+fyXHwh8WnjWWRajaRVAUZwE2PjdRMdvu0+nn
851uaeNTDEPLMvMn9hD7/5drkbi5Mf/XHh7lfJVOpCQVGoazP4p534CynGx2+nSa
cMXXINbWpN54+puNnd0XOFZoQskg52fZ+pK8i4y7y3TRS3wLj1OKbptF1ex5mfdd
6PhQJkaiApXsWz1gz+zxtsHzwAWSQE9GhkIIdUwn4lK+JeaZ5SnAYGkPIGf4bYtE
iTNeh16eas5ejQpJbU12FkBGz8F9eed8mr6EDjEg7LoWHFtQtqUwUKtnfPP26xX/
jumsznAECBuBzrywEcnYDEa9k54UZoQvj2p9zbGaS2vvQXbrDcrJ2V6AdGx1oPn/
S+IdV5C7zjP7AnWf4XfuRtTFBJ+2Wxe8uzN/5rG9jtygNnKQy03kYMWOUHfsBF+C
Vyc8FDrzaRDULMeOrGK8xwKEkfsfCSsMCTOEBXeHRhXGrx9mASl9UGoq7qCPnq2m
RDsMB9yGgM7KPvb+6CyW9fuuPeMmi1FQQJS26Ckvm6ZjVhZ5yKi7no0QS9b+DIWe
YXpKdiIfOJ/gFd5Zc2xkhmVpP6iy9+6kfzaOZ3pb0tt0MTSppZEhoh1t1vr/Bllj
2pRHHWJn6rkkslRv2Sk730iGC4lQaIGz9UeON8Mscy2LC6Awg3lz0qhjG26Pn32E
HNFEQKMWqRFBmaTi1bV2KcEeV2frhRLo6QC6WK6T/yYzOFkTrompHoHcOnv6sBSf
ebCJnApaf8fPQj3TDN6Zd4qLNgpTbLlHNjvGZKQnxTXEmvMO7LIdJarwqH2ztrIK
qabFAB0iaT8okM8SkZC6FbcrdTiPgfXDGzLrvQEyGPwmQEeNKIBpYtdwD8KBW6ZE
KTuLkFYDKfw0W0tCSI+1RmXywPNvrBabjGLKDNoKiX1hkxLA8yjYhfWk/PtutMcO
db5xEq1vnanoPok88oariPgvuq9C8cUNHxWUlLlVusROuovoHPaqqSUh0sWwHKbn
ueXRaJBKKsxx4Wqlt0a9abgMsfL64qYJ/KS1QztO8JISRz3gsacNeavovBr36mGo
74Iew2AF+j4Qt882HcTuLqI35nkqXitI7EBB+xjvKhidFl8edcp0Bsl1THABIQ0i
XuqPbxflCz7UDPS5fPI96VFy6m3p6M2+B32GjpYRx1APF+YiKLcPkUJloI8MSwYI
I3WCjxtUR3QVxXNK7YXVFH0YBfyyQUoWW2o36EFC2XmqGp2y+eIGbTPg9XigZP3v
r1bYtDqVs4PPLZyuYRKx+RzOmvJ2n7A6NINUgNBhMIrzditZ11hjVWZukueZ06FK
e+jqCHSbvc+4/G73VYJL+jhXDlq3cI1RsGtYJ1faHSQGPOxfzhxeUIwL5Ot1A/1n
GwO+lelTCSZSfwQvIjCzT/rGORzDX3c3WGaao/6rNqP9/7rFsYdUVOBilEEOAKfL
vGanbZYNfzFlP7ghrY4W2+t2b/Mffr/vnux8g2ioH3jG8duYfyt6a+ecPx9wSpbO
SdWLB1kNDJOKuy6V22tNucChM2PqZW5BJh67NjrhgE34XoPAjArxAKb5DvsZ5Zsa
2wwLtzaa2hDiN9ykjOLMGnRVrMO7gmmjs1tRyIyjPMVfQ7x/apZX9ZTAl1JOKFm9
jMWNMWlJ4jYkHzKQdG+Cg1zAVrOC6KckkxohPyZ2kAxB9N1l2l4yRZxX92HUdylM
RuDzMNLvkyR65DGy3l9nH3qtiJ4bsaldm4ph99feD25t+ktllgUqrgtn/TMRIRcY
3LjFaotS2k74BDlAovR/ehbZV1YnPcr/1W3sk7iIvRQCJNVuWFMFow+BWamLmV+c
J1zGxK85Zpktc/4HaAIgI5fk6cMiIi5aALJ3euhOXVt59XKGgxM8/wbBwWvVWW6R
OJaafLCLJVHFGq+JDPJq6veciD0XD4m7/Phi/g6vTwhNzHkX8qNuwp+hB9qQGab6
CuOrWNHOHVf4h+YQzHGJumzbZzDBUToT+7lkvvrSnLhCVs58tgnle7KL6VDqzPNq
d8jqEUerFiM9ZX+HVNJRdw1R6OS74wdLGY7RGzNe+Jk2NLMyiKa90aWXU++4Js4C
lLuHWS6L8kYin+p0HaUAZLFnHTDwH/JUde8OUnSLqzU7UGNBGfeBMBJ27ZctwdcZ
6IviV8jNk+Cjdd6rLsRsi0QVf7a6YP+W6pJpkAg9+rJsfZunIiBLVfn7XxV6xbYF
RIrpjX/XjMZfVTS8rMToai4aDIMKg0HXlrF3Ln/sstcxWnDvvRJzgyaGy6A5OZS3
TNO4YYFPWoJ30GQ+6K2S2rsUux1GncnjWPvJbNjoRHajyTPYseJCRLOzqLOPh+xj
kpkFll5/JkNlW+Pi4+zfwKovwYVrDb3UVw8QbIjXDgtvJZ2+bPCc9+H5JlKiml2B
F7WF5hxHHpJxUFV/ZJbrj3SEFD2qHeBYq9R/NUi5rQGe6Qw0lu7jn7aHU5JdkFqY
KOr8aMt/gTYY0vAfgGhHuV75L+A8ip/+iSApTsu/9FU23i0c+hywXH/n8UkoNa+1
vPU8JXESGSguCxD9KvS9c4wOEg0fo/zMCzyg94sV5es4oUfRPCtrCBb0CDOHGQX7
19dt4UHpPKG7dFjDRai6K1T+yOHTiYcH8YdBJet6EhXDPXp8hnmPMILxzvFdDmTk
baVc6fosn3iJOTdwt2hqxyfnJMW+XhGrLK1N2yV7B1el3aaYftk6TGFPRajcertK
Hmv+s5B5Zy9c1NZ8KaCsOZ+rcw4nQ675SgsoBh9MEcA9T4UwHaipLJesPFRoGkb0
ssjCqmptB4cqaDEP1EPl8VKGhQsf4fhpKylURTrooapK1uy7COoL/O2K234uGNfm
us17Mxqf+PRkd7Rw5adPxrh6ecVt6fimmKa8ZvgKpQBxfV5QKjx9+YsH3Bhi31qx
EXJildXODj9BVAoUErIb9n2DixthFPHPGA4xPUTYG8kyyFHd18s7Aniuq/8ARBe0
0fuIbWz12HgI/v9ESlVgm4i4OQKMxWuOXHbbfAtzJ5TZlPS36XwUFvzWp3HU109x
ihaK66VSJ+r4EFdWGdACn8qxv7ZskLbanNfkA4vUJ1evtFRg9sg1itY+El/ZJWpb
+XvpP5PpNTvW2d3MkRmFrFEYRZcp+B+DNoHHpW8XrP5UIKxEyd7/ZBpW/zUVspL1
l1/bDt7Oj/rMmPPEQ1BAoJ5PeL0hJAAMYq0XUnHdUJiaNjWD6/HaKZ0xdb4vaGJ3
X5SqPyqGoLllU2YKPy+ozLbZomGjtmZqm0p/mSvsTde7FYh+fbVoZKDyukSbuEnS
LPZzEnbhUsmE4KoKOi+JgjBRPGiaXhCV4I7WrpsTLt/vyx+AopDZr+hW7zWdwIkL
62I3NIN7DSpxvqM9mQZjibUfLJ59voVPVH2/MuWiD4x9MeFHnSkxuNu6d8eSfiFJ
QKol0gOrdUUYoQGUM6dUyBMXQEAAuHXLKeafvA+akDanwaQjFW9T891OFV7UKgrS
pAz21yw5BFb8yYGjnMmZKWyNdqNhLIgZBg1bsqEz9ml6jLpPrpJcExbozvRI12HX
592GApcjP5zfY8hbQMHUeZ6snR4kwEgFWebuyW9WufVARMXdJKKRZymI4CurtAIs
sPN7NHqqs9OjDAptXW2nYTgi/43AAzDtylD+oY35gd9DPdeYmdaDaqAZDMAVGfcd
of4L8MCi2qYDBcblo1KI6T8jgcp9U6qBz9yd3yYGiKphTTCstw/3voHeXumgE47u
XhvAmfSD2KJMfq+lOxF4oiSKvydSFNFUj2rLzQxpACBmiskdSzY5ZIeWEG/xsaEH
wCYsB+KfV+mtjhWSiBHesquITa46zw8AIufVpjqKpUBhC2jk04WsC8spw9TBasjO
ks82iRlfHeJTpRuftYn6woB99jmbQGnu5ASt7leRDTbi52uYQRfEmkBBmScJWi57
SDSuLq4YNVuc5eWzRcBqx/sE28cHpq6KWvtL4vgGxbOOsF2DM+KTmqAFiIKH0IV0
fSEm7xt0zo1LfFakzQqAYCgQ1p7tEldZrlWVTzEi+onnsUokdpjaeyBsVpJ2VDns
MXhv9pNC16KRIu/zkS4tiuYN78m3MwAIF0hnlQQZ9F2uyvLjk0mTKza62pdMc726
JVQNSJXaeVhhCrpPRN1/mc7AvexBng6AtAcFei/SIwEXzZZf5kDk+AdKS6SZLwMI
zkT8MfDWFkGvm/wjDq8jBwWWdU9rkGCfqt12JMxo550kpB3Idgnx36TX+uWhTUDv
g/ZNshPt4lg5fR3cS2MITDQDZcx1efc/V69ZElsOXM5m4kQYESDyR61nV9yIpx3t
o5Vvi2o2ntgo/fdwKPPDKzjhcgVOlFxxTjfwvY5Pr5qHDLrSOcX/r6LMo2bVwSU+
0UuOYgh6byHtv9ZHGqXKFnCTqNqLFAjykIMd9gcZpweItDS/69ZSVhn8NDBZq22W
erCzM19w5p2rm7a1SIv/dg2nbuKW1+bbchEHEtPFBwUQ+OFRUSSG4k8Kmf559maq
EKBSfYd+e1m8WCK9zsu+NCavGiguGXmwiASeGtthuDMmQTjBRycSmlweiUocuVeI
tjE6bGooJUAsH+RHwu0AO/buH9Rs2QGvxpZIewdl/wWDnjvlNzRtp8DbMhGu1STp
j3Hjv1w7OxA5apNG+f9mjNveEkdxXDYLi57hgK5/LQGzpgN+y7Bm+T6yoiFFjX0g
X5DuPg1W0ZWiV0Os4xQOqIYsPJrmnD6pVIYIuX8u/7SMiGBd0nURdeGOCUPXu++p
ER4B6YVM1+wJAGEPRlueVZL/fgIJAOuXCKyLNATfGtal37fmrRRjfdrRY+/XneWQ
94PqehTrolFw8P2snpfqcDuCCHg7OrVgQQzoTMk6W8vSuWZb5juJnQqwmMOt4q3b
cQSlUT94dmiGkdIeGZo5/PVBa3mc+KE9WVXMyiLoqVTetj3KH+e/ByYhbLDmhE3R
XOuUYX8t3f7LOdlNSyI13yCeNLkub1oPkiN8QeMT6Yjb+NQ7AFsCdbiDxX/qXVDz
dj/oZThgO1KoZidmHYwrMiJQY/uFL0UhI3UE+Z7jg54clYdjK1BO5KWlDUTZOblV
wPooA0fBa1uIu6OYKlS7CWgHV525gg1gYu8I+TcA3QOKYLO3gkXY2tIvDd1Sw1tj
kSi5hhuljS0/KoWVm9bUjii7OweCm+mWaFePMLFC5cFRXiGZTX5MqG3s3t+oan3t
n5GZot/gDkvSXfKPIF2oFnbXmSFJbjSoBS/mZGZHUESgsZxvKJD1o7VbR1ikbdpZ
ZQrA3Q7mNE/wonIllxrb3zH0wj21L4+eQ63O0MumlovKcjup3cgUZ00CepT2c5Q+
wbLrdxiDKA/Xemfo1OWvSsPG1K7aneeqs0kegEp8YfFH1CbtfOgGTxEs/dnb7TrK
qtkLyZObK4z/6WVY5g7bO0zC2x4+563MQE/FGGT4qBiKDzKuz6UHj+tLN4oXXUWA
xj6IIsv73TkUkDdrvFVMyus59AhwD+rs+Q1qjhvjGiztEsLjhbkE91QfEguhv1Qw
fD7z4qUCgv2Z6JG0U+GHv2ZZYejcwKy+auTiaAnVO0miKXviGqbMO2P/8Z5u+fnQ
WvIGgdX9H/8ap7fRpLmgBBzLKzkZssY9z9vvRcxFcP6z7a6SpJXVsB1KLu4lfzP3
Y+G+2hzZBGXdxjL9qXyyptVrv09FJwVh7WzhjWaKcRosze/YTiCkld49cz8CrGl1
etOJaUPjKz9N7iWJLKIa6shGDjMPCQ93VMOyLQyMpnhOe8yUpcwX5wRYF8Qszl6y
Bjm/27wSJwT+K90/Dk/GJZoru2BlKwzCsPXicTr9mcNSkuS2gZmTjotjz6euJ6R4
xpG2A6SDbueqbFNziNyECr2neMfjSGlGwLTA4iO73vp94U0IpOiuvH9bcarxivJP
BFEYn5HMDiui33gFoPu26/KkjAQxisYEYga7LLRNdlymsMtL4uqTXOyCn8yHmb0V
J5adr2Z08jHjhTMgAy6f3wg/s9p7WXF2MtJxQU2vkjMJbksEjRD1TNI8pP1C6jKN
1MFX821M6lYLLlJ/qoppK5WcNIDBjEirDej6Oe/NAxk6qLz4KyKoZ5TbvanRFjHq
B2ol11v6KRVt6JgbtzEQcIBDBVPOTwrzQTtbjDB6LmBAzXLvd10ICe4FqLgJmyZz
2moxcSZngNzBzYnEYdE7KntRHqeZD5hLRJNkO4meRhfbP1yj3s/TYXZRo31U0GMN
Yhfy9Fq7r+t+b2PEsC3Yzc7DUFCQjJOX9wEYtf2dyeUOqOFHn0qm3g7AvceZzXL2
8lrt9pqarjIR2IX7wiZr5QdUiZlBnbTHtORqYLoSE70Ns0/1u2jkZrBFfqtVBXwf
Q/5WBDT/UdvGisQ1u0LeiVzZ45iUFRRetZSr5zeL5eOCjQV9ZcDEZQTjVTUve9ui
DLnnU/9gGkVvoyoGtxdAlIPDWrIByfgcrw37rMfvLzP6EZwFa+AeugjNVaTNdvl8
5Xl8d/Y+vneZGZnI6ToN1eDzJzMl9tCTqu5kvcT+BExjs1kgrA7jjYZvwunilYlU
ebK+iQnrR4SxS90DH0y8EZxf0i79tgjXj9uewXCSpTxm1eLr3np2IBPXCdJ2mBx0
7ORApYCtTrkarZbRwR66m3iFb92UHhiE8tp1+HO533Pj4N2pIYA5lVJt2MwBLx2X
jqC2RK5bQDlvYo1ofxSO+VTzjMWSoHUI9VdvfyoZ6aVgudwM66CBpL05PC0Q62Nq
EnaSwwjZNr19Xc59TY6uOZHEqo9dFSoF7+pDHAO12FVoZkJWoNGtObFBCc9bPbRL
XgOHjmqwXuXFRkN9YWe1+8avlUlJ3rl3NOGi0rYVSAIlTCHsI4sFDHHIeSy1fJXb
oWQg5nrSRVSc/AZj9aae2CI9onBi9Xspp9rJ1JW+b0pw0EHEpT9ODxLgPScn+/zM
ZLUS+3O7Si8VtIGnSy7uZuCUTSa5erA11Ctvbf/9iy4ef2D8lh5ycOK8fd02UN8p
fFHZBp+NLyn732MOoN5bMUM9rec6StzOfr0krbuQtk8e9vEak8FtHAE8bmh9jq8N
0sSMNVcUlzb0LicSWrufXmcwRCB+LVlXvwkGutmLw5StCDPzWdT77xUK1lL8lWP2
IsKY2PteSTvADBMaRTSOq/HnX5KrBLFeATfbsJxypglNbIz7qowvAhW466+h7D4g
inle8qIUe2iCyLD6Kpj2S+kZITLxaFRpZ26TKBON2m5ml7u2k7+gHfAvQ4fXPG8B
uzQdeLmbi8MNU/T5LEG86lEfCWtZor8wdKDLzXMngIYk9b6VfXR7kkqh7Kf+SZog
UaQyrZ4rrVI+QMXyvmW1Sy1qhtHFOm5W4XfJOBBTpk91+R5upN1KBuk0FXN+q2qJ
S8BdHuujRd58S6RBz+QDtBc0xdojrWqQhf3W/8S5fGz770/eHEmfW1O4QRhfidse
AtWFSrPI4mf8bsvJ6SgTNXB5HxZEZm6yXhkYLBiyQ5Qj/dTnD5COii6uuO4PVM2B
Se/TyPMYaxtrsD02mBWVTz+yI++XH2kOCKvKGZqUxJTaBEQAoIbingI3za7j/cES
bIgp8v7wD3rZ/82xeCXMjHiUtl3E7YFhEziD5naOnDA+PdaJH2XAzs1QpUA5iqXo
kiyhdFfnEpwfzm9yuAiEcKve6v/meoNpb4rGoBJQ7/ugNHGaskinjTFACCdqCRZm
EAf7ODOFNztutE3l9KFUBIC0frRJSQh1Q1K4GyuBYFCimEjZsqTzzj7eRkW0oMN8
9CtvQTtNgcKYHI90/NzYa8ItxK4QiiwpdvQoMNvFxafWwuqofjgBmouo7zKbIjEF
ArfZTeDimm2YSwHlpNTgrK+Gq4YVnxb7UsX2U/7onJBmGwbk2cUziZT6FyzUisoh
zWdNShR7yHawo+35FuTaEYah0BfYyaduRnhELHBpor8JtloBwH3fWQfYgiKBStLp
1ZspysA/I210ADhrya+9pRfstX2hEz3VrLLkLhEFekpE9EuIKUBn4aNxQIPXqhuw
v8FT+Eh2GkUrDZ9kqJMxvPWHebzO+IiOftjh1X2ucQGpSEONHjt/Fx126Cp5zIPR
8+tyImKkJaPmPLvV/Rsc9Xa6T0U6IacfK8RsTguqdL9F+sqfaCq5sokD0TOYHBzB
GnucqcDPEYO88MgamzeGbsuQO9JqDWevsU3E7CfCe+uvtkbMlcGuJvzj4QgkLjK2
hj3UyIUzowFaPpOIUh7ZvaYwV3GVZRsO9kJTRQHyRi9tl6DLsZBONX3gLXxZDzB8
Z0V3LXSt0Yr2itETPnv2f9q6cdGqP4rMAD+r0XNRbWxyuaIgmwyZTxfcvu93BKTC
6tAXMRlySVYUgaO5lIyBUSC7Zn0oK1SqUnQRetfDodpFzsJWbySIyLDrgG8n2Uuc
8FtpmisvxsqpBd1k7LomyNyq/rgSTpZVkk71AmDNl5+awkmMCxPAf1C+Ms7U+Hd/
qdlbdRBivhCyN3w25VS7o4QHYGYZvPvjvs1/7Q6bJ9NTzf2TZToKwuJsNAuDnr71
KrxG3yOFXJYZyPNrMDgeo3Z+1epEqf/Z8qHM48bZqgkY7s64Bu7DrsO0Vxkpa3gC
LuVgQVDr4Ngf6sfBGgw26ZpAybSRY13R2V/W//mJXtfM1iPtwMST32Ixp6WbSDXl
jI/PZjm7W/SW3/YMcMTFyLvx9j3ob5kn5csi6VGgRahMNKvZKllg9G40mQULqQj/
pVf7itXiInjEztIkBtarpV0gZsSoR/V08qxaV7mvJcXSmwZhmzQ/IFUxqTVT/++X
MIw6I/L1EED8uNFruvb9Po4+mKXavJxqyVg5gsrsFAmvzllYS0vbTB7Y2fTiurZ3
wEYcoHWfqQsffFhtyTvHVWlSBBSPc2py4W0xltfa6ZNpfEOOTGZNtMpX76y7LYpy
tv7/ZN8cdf0/MjTI4RDgRzTo4l+k3k9/k9jyeaixj4H7ucDt2GeMgu3qYyhdZSHS
+FahT7kbExO0CySGM5X/wjjSfLSdh91uaK2wRf3bVllnc05aQX7YXEW0q/KsK0Hy
fz2EiG+GiYRAQcfwOB/WxuJNR35LFuSYPB+w+nuCew/9OwbanP9MQmzNq5bgz+pD
U7ov8IWyATTTeAoAjEVESkF1uhQmFh9+fThCKvnym5NwtUJxMgklBulRiwcjCd5x
olXKpyS6e4fm7Mq/+T8IIRiEEQU7yETnYGapcoottSliGyVE3sYAUG3JxRSHV1tR
X9odvZ815EDNMxGv+9yY47fdIxTmovOxwJY+S4ULIJHAycCxmCAH0WNHGZRtvW7h
8rib+WqBDlH0l4jEuWZYuyMlprchMe3JAxVqZDAEZlsBUqgB0rKE7nEM6epY4Etm
TwnVjd0WAzrS4yL+1wE0W0ovtJy0lRPBQxMiw2iZJ3Ll4LHqt3KOPGLZ9/8uxZ8h
ldpDn4kUaCpoFvYpRVjQQboCWhIEuVZ3VO9CbJfh6c0hwrjYGgOetPg2IVzkeRvS
F3AO94SP8q626czTTcOLgOJJ3oEaNXiWGiEZMgG5QLfMgoFaRMaj6mGrrroKsoas
YLN0BteVoRzN3TrYYAVpUwK98TBUsq5b/RunKbxsncNkIlcBEhAVl4Fi7RSusQds
KBESReD6KCB6xcV6YNinYlg4VynhSF59F4fuDgjnLmPnAtrGjueqIe2oqjIw2IYz
x88PS8aH3P2RdBWPj+N6uc+SE9GrrYoo9tWQ4UYBJSgEx6jKj/QKxRk5u5ZNJkMZ
IxjoDTjNQZHh85rzhYoCiJW4Hy82mQYTcCdLXn2oXArSbXyBloL0om1AQi14fnVx
DbW2ZGfX58xTBwQSJQilbnTdlhVIaOLPRYjN+3JKDudUopGwWoJhwHjs9h+nJFhm
sp6ccCT/ysxWU5N3qkzd1rwwnZqlirM7BtFPDMhOYox+ZSHpJUp3kAXvoCCT9W1S
mxZSx2YVs3mxbMjfAxwxhpYM3WXHHlWGDam6qKkL3wUDOZWgNf2iaviJDXDEuTwK
JFGFsQs6owKXe369UdqckO8iM9jbBWyFX8aHsA3o2AgP1DNdT4ZM0ltxUp0s5ZOM
r3RYlF01t1OxRQUaPjTA5IyIGfWPytJ4AseUAZMwaL7RdAhpsgBkR60djX1yh840
At52eAlpnI7RWwi+2bS0Vg9JIgQmbLRJpkFet7OPXvCMRn1HA/ab3Q3TNRIOfHV/
triiCFUbVzcrAG86Cg9JHPGt3ToMlBsDglsDxBNl+ETC58qdSL7MtjLQIRK45gwu
JX2VclshNJd9QzW2hYuASahqL2vn2uje3+1mAg79ZYzkziokP1Bb/0UuYmeOjX4O
4akKcfZUgeLdYVUdq8it/Sr49X7n9NmzD04Tit/Q1OErmck10KsZ5TUTKw63jR2c
0rpEB599kRWyCOXgNKgfxZqArOVQ9GVjkN9PUSQzA1m9TWHWp6v7mxPNbBA2wIdW
aPHbp+zcCCNN4tPMD9ySp3Se3qBCIARPMRLh42yLRqfNICwMZWZsG42eOgCujP12
URxU1D3a+vqmPMFgE58F4xNcBSsXKRCLDMzuG9Ki2TY6sYWWwcG4+R5l7n1ybdIp
klYBhWqwWkzhWxzub9FRIa5nLLWsN3xnb76DHNA3tR4tIldvRgzQbZVtx2/5jaV2
jrD2b2a1NPElnZwrsSWL8JE8ooeeUcnDW01BPfH8ce9w1qsvYB0YldfqrYjQylyT
rveoVZAMzchat+FnsFQIVwg1EAopH+Yx72PzWEMKa57BXVustASVqJ2hSuFrZNUa
cPB1ey18y4sMztX5MNRj7ZGTa3MB6iqmjefr5BjuBXaRr/3fI7xnLvDEiPRSKEZB
j4D4cIrujU4RbLeT0esjC2l3/o6NtkM+IgszSRlMwqCvsxKvOV79tWCw8bv5nf/R
zoJQDPrk8LK7qRNz7uuOl60nKH9uvjdVV3kWWaGpshpjQSz15J1dyetJ2F2kOygv
NoMpzMdop1SsUEJT2IQ1zeqDZtvFktBuNtJBbEXt2kQoD8eRuKgXAZDQd+b5N209
H88QvxV3kdGI+neQwIGf51/asIYfN1c2znhK7Dc4B6bCqjZeJbnxedboFlzwf9rX
JCF4DTJrVEYJR2JlCqAFQdLOy9v1b3qiqmEHGhQWbH+WU43ZaNMU80uoxtCTGKHn
xIqi0xUslmvOML4LIxWE28ZqiG+a80ujPFKJ7sP+K5xgE3A2S1DaRYU2W1p9Fhqd
Tf08i+Hhr5+k1MFGXjRJwrQITgXqJHk2EASDvXhSAl+6z2x7IcrFVFryuACVPXkq
ihxKrjsLQgV+HXRbU/xXpK+NcE68TwFVwS+mbMsq6Vuq9fB6QPx4y9ZcbquXbmWJ
Qn9fo0FGkMO1QQDv/uEdLfApqUrLSTuggDYVqeIOsNt4DhVgZmf2e88jDeXm0/+o
vd+wBds3GZqcyD9QJDAdOwxFAJ/poAhMwNGdRfl8gXBzEBI1z3sPTYarVUTm5eGo
iNtg4dJXYOlPRVWYHOHwvbJkgECj7VlzIcTeYfoQVZj8WEOHgI0LQOZTOazH6n+w
oWun/HnvLcXmu0wZOrvkJzZkPUd6GuX4RnTL/0Z37qi5UcjHLoReILRaawZ+GTcj
D3n3zyXr36dR27UrqUHghq8MiGv/2mvzniOX/pVUF9vYEG0J+LyY+VV73kvr6wVd
TNvd9s3Pt09hLE+1kkIeKaZern2JKlPYF8Li/VD1cfFmeGGtZ6OncxUmm7SHfUu7
2goMeeI3gtraSA0ORszT8XgFKLlnzhpQ8SlQBuH8sixIZcKF5e+QSp6bZxWRCNIG
+MDx2A1z7RZYrgGaZc5sNWq701b57m0CL+If713BnUzag8v7wTsWmBcc8XwwVzJP
myNkG1uRQCe88R5zRWdHXXtfSiSwMxuabufjqUn7A63TwtgC3tepWkQu4bYXnSBt
4nKrjnOFP8nOcM2+qTdlKhgsglCU6kBLL+yzWDV8TJroBwFl5SA1IRLxFH+lDR63
oAjepZgf5grapjYBaWjrul1KDkG+mE73OuenyoFRcoDFIAfE+VpDEyi3S0eAz5C8
bNU/sxYRzWI2D1pWTVVTbZNkAse318H7R66sKG7pCc5/YFVqcwgDAEqf/EHWLBNi
WoUmkI0/Ta24h9N3ZSd9XYQ6feEmgCutnT10ixHOiT8mwLpdFt4MGSS5s5Cs4GYi
m5UEvUOVr+s28rh8kZ13JRiEZU7H3930BjpEyU2NJD23+pqTnYE+uI1tvOxrZfgo
eRzYs0Z+YkPyasz+YRe9BRw4zRvH8Kd4+6BqDufh1FmUM4wpx8xAslplvgixo6pw
WSq5/c6Wt0a6zI/4p6Uh8+SEIZOtVYunLFx5AswxPHLFE5B4EVtdjy2EzyFt/X3N
mt9KUKraVTaVRgPrOnRVWUOmoxzlxCxn4UrFNsRzLUIMHYgwUuiUCRCmKiZ9Whuf
cMmMNFuqjyrtvPPMYUdSw7oTulNdnjwuxPaA0jSopBe//8JQ24dyVJkxxKRMp7bE
S8fUzYuSh0pFHqIo94HUivBaMixnCmkdfXSRM6MuBEBHnU0WuSvPsc9sciuS0Bn5
rUAuoZcvyA5FfiKj7G/4QZcqQAduxr0ilVU5aLV9ckhXDuAFLm1awDxD9zYyUlOj
8AYIZx0tcysn1aP628oJE6IUP0N0vmozT+TJq0svdVe8a9ve0QnZ089UEObdqDgQ
v1ymp0jwQx5GSWxvx9ux+G08S11FRxM9EfoH0wR2lp2oyJ5AEBCN2MPQIJnY0054
Aa8TDI58QtKOj7pqiZCNtmaRgymdKggZIrpx1GFCbLrGo2hEqRhWPczq2/WVC+y0
bmM1zvZUryHGHZROE4xL40h6+xQZ0ZcE50mj80Rio9k52ATr+IEpCrTajJcH0qGy
NjJbT+VC19GpohhAVaODd1vHbJucn4xj9JpIdfjoGqYWj23iL761cgR1XwHaSkNq
AuI5FZxEY6STKD1L7XpRIcqStkZoxkQRohZBd5tjMt+hhcgTYxIJqpQWShF/21/q
ouiDT8ytbFZlgeVRm3nvucb1SuK819HnDAon6QgBC+VXKdTZV+50ow8BFKwpE6xj
smQ+ss4/Bwir1viJeOpDZC7b16DIbtos2S/BFPIizB28OIu99phpHkV6L9t7GW40
1TM4CRB+L4Amib5FDh2ztcJO9Uw2BJpdLTBHFfrySG6A+QUq1QED/nwHGE7u1Uc9
l9lak+zpU+PySUJ0Xtwf5tCfMt5WUkEIYg7DTcXiZ1/aZcwPhyjiW0UoB+0kNOCv
UO5LUwUrD8krnLNszxGjrPlgm/RBnHyzFxjQreS9Y956OJMmGZVvGCv07Md6rjeZ
CmrYSGLWVvlsZgvZxJQtrl7KxOBtG4eAqsP1E6I1ft3MSNh0/x477wxGO7BX1DeP
EQIXJiLf5KRsezvT24YwaC/XN7hlVmi5SpvO1BXDXyHgvv11U6irmT6sg4tqXOQd
rupUCICkIzD681kuoZLCgjq7PNoQe0azOXePwNCbSusaD6t9HdOl0hAnfcA5c3hJ
AyBOQxci/qkxsoLHS2/XJPbHLtjmQ8kOJRVFxQlpnEYxaaWc4rH1hYkWSiTJj3Ej
LkTFdWzk+jC0qOCNCQFZA6FJildp+Te63amurNZ5WracMhRfltGhN0eJAxS4tLAF
kV2MWj8wQ9IzxnwpH8KJw/37I9+V1DMlp6Wn6cbDsjKXw0hpOp8pTd1U8uhjm3UR
Z4IhNysWHip2nc4nopDwCG72rAvbeZCfZUud+iNj1b6LpiMd2MAMNJwuZYaKn6fq
c3fLuZigVWbAwKYM2vQ1B66z/8qg3aKmAd7ZKeewstas9/pWhaM5Rs8U356EUxn8
NzNcPjrvuKmEZ3IWWyPLdABcsvItTWJvALeDlu9EVDgqswqMSrXrqDkmL2RouOuO
gqm/Yu+6Wnwd+KYReLoCSZ2sOpzuqlkZA4k/N4yM51KQMLuhPw+LeZ1QCmnF/0uC
HDl/FXzf75ouRSfVjGpBtmo+48bCKe+Q1RtuUVbgiUfyML4nunsvFd/ZGrOg60m5
LidE10yXgNU3HhvHK6ZyLOvRhWpui8/J3zSw+tFw8V8DrycgiDsU00qYeFKYR/7C
yQZMLHsq9lUKMeA+sLJr5mzbfZetB8qtuvTV/oQ88Y3rMeFjMViLYUhviUTQdJO+
BEvLiiQFsuKFdMnIUJtQyDkiNSUJQ+/u6ZvDzfQJosnpYpwQLq/a2JZXE1jU5apA
Xhe0VS/Nw3cydg7aL7UomQ2mKgzPdHFvZk5y18YL8h3oFfP2t0s+1qk26HVT7eZ2
H1m16bCqiOZEECIthq390KQsz27G6So1X/cZg4ISE8Y8PIrVlY2lx+dLVy4WHG7c
WsCtvirs3P0YfZXtrstRObb50JjLzHKmOwe2LAClIImk6/2SA5kSvREIxqxyeTef
lLi7bV6qEkSZLEvBAX/oecmAo2GY/wfv69t2h68MCMNrLf/kJeUL2G5gTgXNtXFL
pjVV5gWV2bwGP3kApk7YFwD6SkDRals1zyFHaDP/sRx+QpZgsA5tdr3B051K0SV4
rpqP4JlonkAseX4uMPMiIBFi7KuknDRFdw4nhy7AWHchNuxG843TxmikEQH7X8Ah
46KI0yO48lYc7rryzaWXzG63jQZBcbciyW2bTX3Og5sPhuLokH4vJjVo1l9A9tGx
Z3hHo7Y9NnilYVxwGdYG/vAUNCMZDrqRbgdYuHHK+6lgmjxCIqpeNVfiwX4MLUF+
42dCiohGl6TjAq6Bx5Fyjbs6YLrKBWd1MVrE6zIeOA2U+SZliZI9R/Zuqr2j2m0m
xylice+ACrMpGf0npJTvdkFXshJ3qKqrcdX0zkeU1mvKwHGrUUmn6rt5lmJ3RkrJ
Mvc0Qv/hqYtSeHZ/4/3kEJ4eakt9oHwhwBvitZYmRRrkgREL0hFT8eESps4/w3AE
xCe2oF0FrIpZRNM+j9Cv5+l2VpzfyTZG7ULieLd7nRc/8vE96Duebd+Yj9qJBbml
14/Rn+EwriWCjELffvhhqH+JgPlQNRKkTjQPHXafsc5mpIbJCOvMvJ8pWT+WB3yy
76N0Bx0/I4PZqLIFwXdvRcwAGi3jnBqjJiU7F1fUAmam5XEL2DPbyIIhoBTFqGrd
m6iRuiHY1+PB8FAyTGU2TCzsV6XYHgX4zTux6U2NChMXSnW25J9zMMw5Y2uaXQ7Z
wN+DBnFThCFi/4bXuKkjJInP+/AU8371l3QAWdhd7DO6EsmhUSUQO65rmsHGPBz5
+csXnU9mIkFtb+UB//bA/QtD7/PIocrTZKk7qWFX0mQL9Bk41gZaWAQWIMguEmS8
AXHdizpNROxWeWJOz+g+JnCxTY0k/0vOVmbWnq0FUdq/ltqVLLJ/368WZKnDwZ7U
dh/KA/xEK93LO2yvQXN6J3VZ1JgFhFCfPN6DNX52cEkMednpN70yptmHYfLaE3RB
0W1wi+2AJNpkM/CZfLJ4yrXC8Q4fN8IifKVLc3gS2seuoZDfYYZnwogF794SaZXI
YMkOorFhbJufBaE4NYe0AGIIRW6uwBN64k3vmhy4waLX4pXvPyJAuoyVHv1PMKhZ
Mi+c240Za9CkxOybwdLNGb3OTf+McmfsaFOs/5VOlvcnMxWGtZiukyaxSKOeFvLp
KugfWwMKNUjlk2/heUlxRg5aB/iVqrlMy6BskiJHHMqCyCAuDb8Z7Q04SyvCUcr8
oNideQW23ShvuUGEiyBM8an+PrHkOEMMHs1ewVj5dvlF4ZhrXnG3J00gTY47A5Mq
ScjoRHsDR3AopSia4E8bQlnvnDeC1ziZHqjAx33TohHcnV+bMV68vNdb9bXy9KjN
Vmld+gsm6Csxk9K8EPWq3Hi863g+eQWCyk4tOF6WgiIArmdJkLNKDJ/attf0kPHR
QjfCFH6t4I0BLRaeifERjZwzBHkMjYjx3mVxa/2afRnqXG46qYpON3//txDfYnFO
0/EDX4t2gytRUHbsL0nL6do4wecpiPTA3/nLh4CczNCK+/OUhLC+VJwte3vSkm2+
j4H226JG6yKCF/EdHnSx/MqQ7d56xNvTcoE6uG6FQRW2ae7MexuSyigX+wQ5Wl29
EUCSGVUsMhdrXkJgTwJ1il0CuORS/Qe7fNKa04DxgrYOE/lcsW8HcZo6W2MdNpqK
zJzZP/SR3j9PbrerdPAcuYXQmxEr4wfn4gnaFZhc9DwiBmjvdq0F57bIpBylj4gQ
ilMWkaA2Z6d8uUF4iu2oD43wyy40z+uP8JgmpGZqAjyc4P5ao2QZK7S1+I4ycGYP
VDnzm2R1bVRkzVszkllN+bKoSE6Y+NfN07oLmorT1qid8Usk3W+Xftoo4pR6vtND
MQ56pVxS6eV9yQ8kuGdNMUotkJ5x57z9yqdG7sw0j3WiV3bttzpij+kr7Bgl1T6r
QhcfRUC88pH8drgnHXUhlUcRRGT1Wl0f/kjlog/rck0Ewtjt9eqZQxDnGQaSHmh9
/RIU2Xj9j4MPWPRzPlRQeYJhGSsLcixVfH2pJdttUbUZbWEer+OmYTDOx01dlLPk
1dSXn9h63BeEwSmyxDzU+vkNyqLzLWnrSWO/kQEViThXmVm7pHf1O88iGlrOHA1r
EXgRjV2JfHG+G6JrL8BGghfjX4pgeLxjO3LGTfDLbt48XGVwA7c+yrU+ZyVUjZNH
SEDXrSjVL20efm4Op8n6N0p64mE3FtGuRRvCduBtPiAavWnVe1clrCxVpDageozR
Ru+Gp7TXayWGUNjxWwD2fdbV3NkoH5W9xHMMYmym6vQODpnk9INz5UUN5RDFcrY5
6WTMn3+Qx9vG6adSar5cRz/JA/0lntJUrEtTVHVDlYG4gQzN8oUSO77R+tYTVwWc
P9Qr5BIida3DqLmwDcgt578pEKhakwjtY+5zCMOal1SdbgE03fqp08RvKmg6pY+M
FsbGNQJbBZzdIpCP1ilWjec9dj9d2hIgFEDIzWLhsk53vvKJq19+Q3cycQVcGlH8
73TZ20WACiIsJfzxVdNNctkb2zSleLOkHJZMWZC5AOVv0qMJzERVvvfZq591jtiG
+cAAsDKCJWBq4g2NYevt/jfLpYanpUtd0Udf5Vbr1Qc5Dnrynm6sCD9xunFM29Pf
/WeS19KQwocgFdE8B+A2hQp9MX3uBl79iMnF2k9RwYlSOLAoGt5cAo4gHr3Ha9/S
pO0HBAP/d3x4g+P3+tmq2CMkVwaqDtCI4FY0cDHobCJpfX+YZKzdb/i60FW3Oy21
GAe61XgP8IeQVrCKP9NMMZupXeb+2lcn9FIsvT8gmDn6jQ5pIllqhfrI+cz01mmY
yZqoeo37mN58uOZ7IYPvVuumrgb3F0UCXtUKTD3/9h2w3MSOE2CYLN3kD61MDMKE
+ntY0xX8B/ANj8LYQeAafHafEAzpoSL4La/G/hKMKEbZAVvSfHaxdkCErYjiJ5sE
8CsAjh1kafrmA/a4CZgJeV1dM/ZgivA76snnTib7NpcmzUvUlXcSHd9EpL5uLJb3
yn9kgn0yUIOYW84vHErMt3NGSW4cOBUHT8U/s+fCkwyiiKzwjA8x8o7HDRWHQYbz
XK/BVccfMCY8qdPkrBkaR9vYTDDBuOJXbFBYvNbYZk3a3oWoqEOZhZMvgdjwllyE
UDNsG3mIjg8Zx2PSCpmStyP3LHMNSDXiYBB+oVnSVgVhuaMHfdcNps3l0j0e8Hc4
tC2VsLPy3OZ23crkGknLoC1w01u1NZ3HC+BJmG+D+sxIUzSvcHmR/1ishCJW3k+J
R5n2TS18UCO7whOFD+S2VsS8Mpn46iLMYNZ5mZcZfUI/QtnqvX3hZxnHYmwMinpW
1ShpMZeFSmsrM6bsHd679EMPGto7w2dLiDD/4YD0f1Ih9vC9lf12LzJgF1VI7xSO
UOws2wTZK/FS1jZ8AK6FEBqFK5e5TL28O/7C8SjRmYR4G9Rp2VDZZyUBdrlsGC9T
A8l70pStatZQ9mjvcdoRYCEynt8vIrpBkEIhQxq+ihd4nBqx5dvyoMno0qR64t3V
QyPBpPgGVCNCa4CJO4wdyAPeoPSXUpJ1s3zTPlc1q7EgD7Sbu4uHlI+cpocvfxVG
IRjFnrejfhzmfBwzSffW1yX78rxhoL5yKAJRmFeVL7/OmMMztey2zarAZbm4O6fr
wZ9doHuk+5zS//x7WafoEt7lzftk/3REmHyAUmwxKosX7k2wE43uQvDkxHGB33A7
ZOKP3XxDXuuLyXR5aim3kBsUK4lf4KTPvEXU7iZ2FyB1EhYLUSnUXp++14PPTCwW
yTXx1dG8nrLYu7x7Z8gGBE2QPCB/lYn41ZKIGiuDAxEvh44/RwW++ALaLgmMQ6rJ
0LITV7NegUw41O7Xt4QfcepJPRsH87Vm6XeQxmHc9w4sPsHmj6lKC74lOuB3clTY
FThfLhATvfmiWwdy2Bh7NowqTFVf/U5gaaJgwGnLCKdgQ7XjqdwTVgAh2XiLt5bU
3LTc2Zz7GzYHF2A1Oj9GgFS6QJzVo/4DZf3nWFLQAC2PviKyT2qvM+ftMYsHAtRX
DAclJfcTM0Yw3a1pI8oA+Lsiqe8LtiaO0fvnjFSoFLwKejX4rg5xgUHxmeZIIoVu
J8+haMY2VjSMWnIlNFhiXOOsKW5FE0BpwsJEj1OJwrxGIBY6E43dX6ZSLYvrSq4o
uF+kdwUpSVdJ8A6Ihb7NTaFdTUWgVBTG562MdcsuVgoeY5TxIoSk1KqZJzaUCKKK
IOSOWYkgYcl2BctJ8kqtAbimeaC56hZAlr1Lm1qWYoAFBtScjfnRX9AVV/l47FF7
Ep5vKWzZMh4M+HaVWQHguG3UqG+zHWaqrx9WY2nM4lRR2jiAclzkcFxNbn3T4gCv
46zMYcMvzJhtr6lFugBi+3kDhBIY4ZYCDilQMjCxWAbqBlGt+BtUkcFQuDYyHvjK
2xq3W5x+eH3vVfMMLde3aSSbcj8NECOUWJ6Dj2y7oSiqdMvivFPHbJSANFowxWxo
ANgrt5dS0mhHL14wVtT4r+Mkb34S1nC42lKG7PH2l40FvObQd54Ep3HtUfhhJfn8
EmdOGgHMJ53xQlC6V5/qEGMvDpt3diXXdSTPMFbHjyQpDA5D9ycwPURJ6HLxdAhk
K+afzFL56A3BGkY++6pQBxJ9XsngJFwXgGpKWfI0bZjlSZqPO9vWT2z5TEf2/fuw
1HN1QwwmB2qrO3ml8tnXCmU1KtqjVlJgM7e8JdF9pGas/R39vBJ5uP/VBGwRKUea
eCvT8N44ulPsE7h8kQOPfrrlepql4Q5rAn7B3UHVr07NtrHCSXVyQoPq6RAmAddZ
sLKBUiemNsnDp+01a+w8owIPF3rdymke1/iRlNd6IHGsqZw1grg2xAedRI+aoaZ2
Q07dtGezxEkWyCcREGDzhNu14n5g+ioZFzphDcBunoxe+eYlfaA93r7Gp7JXiDsO
zZrs8EKOUe9XsPsysQjCZrSwk/CH+XPYKWQx5mHW4V+5Y+Ax7ZLHQtzUajHwDa3x
fpb7irYppoFhTV43p9AuVRuDTBP2buaKi79h5mmxHbd8BxzC5Hi9oQoub/ZqLvTz
Wah6Mlq06bDhg7ZD2NCVMxZMhkgOD5THZSTcVmFYZbJGqUAYum6wefP57OZbrvRY
HzWx332E8ny3L6eijL3jPy3WJDkcNXiA5JSIT3J0XR3Dtg6VoCltsxRKu+5ufIIK
3T7yH9UN6cE+Is4GgrDUe6RK7cWELT7Lulq65x7Uw9Iik9z57iNooMEz3z6FLGoJ
6LebANg2s413Qwaz2uf7MbJKGrcnUQGlwmdi/jEy2Na6Ye7+EDi58T+VCTzU0414
zdoPliTtyy+1Ob/lWgKd54rrJ3fke8awqhZBZhwWRa3LdDaf3sbRXqmrYaLjUyEA
O+Vc1gBLXrpcW9+mlFBLVu6hPA0R+pyTffMJJEpqTz8aNx3ivng4DWam58hR+tYa
cw0l/rFGIoUX72Riu/A680SK8rvC9UrAhEyN62aLYMOYa/S89qfTcfZKop6fGg+R
FolsCmeECvftlH/TeHBzawAGDJiQLadRKNZqzKBvsRtP6y+zhaqR4GT6Tyz1eA3C
zEBTUXhR/HOPfZTitpPl/yM+yFyqZNJ3iVqq8zs2AeiS5vEhp6ZmZ51eKUahaR1X
PQ8bSs/tRANfkH5QLFHKjvqjt24pK8r6xNQM2LNfV+SSsQCP94dgfQzJH1YMrD09
BcgMkpT/L/Eqmp3nfMBouuGcttfIm3yqq3H6hsCzqIpISIIz6qN5i0Bv0r7VnpqO
tzTlDN1lzOenxwX2JRGXoO8zDMo4IGvf8sQQgtuazOvjm3cpUeFXppvluUuTn4xO
9RI0gJugNCTiOZLhzLNtQipoLJa1vuT1gxGiF3AFWVZU7DM2RFgDxYWtCg3IW7QK
ek4YYfec56xXKZu5VU0Zu4NHoF4fMnYPvVb0NNiinaVYq1cy13HaCQycliFZbkzo
S5SWIre23dpvW1HTm6Y2X+9RKli1whV1yk6bR2ChvJoBW9iZ+OLYMBeA8PGQDkap
rn70oAX2rCEt7zqAorYTf8YHTXcrhAmz3r27Ovi8KT8RFRVw3NMRjB6Ak8GZX5Sp
/qUVwZ/c/oxEyKKHEK2cpHqSJygXZ9YYnxdRwf7ERYASWnof2qJc4xsYLKmOUX1p
O3vkeQLR3lHl9rbueG3MUc7LBDcfjz6erxaRN/onaduueGalJE7986xgfPPo6iTi
TG+pk/XazY8OfcPlzznJD09RCxwzJXYDdxOo/AQvNOGRdV6ulPxczvzLZobZUUkv
xzd2PHtbkAlxcjwlbtT+DFvIMobwkpUdlqphkFp5Sa7PV5jmIk7L7VPsbqTcda0L
KStLlYwKrMqt9TOcDLilvfwPDYEFKeVmRSyLTMz5n9hhtoguAh5PI3uLQ2FqV21C
cORD7RVEEAyPN39jgSB4+7d1dag2aixSlK3UTqMF73thcl1HFE4Q+GhFPmrVNLSf
GtPQdwqlQjl1dlSWsCDEO3m92kV28gzsKiTeOFbE+1frnVaZEWQFuaFF0MznJAWY
0i9xvGSqg5GqmstQiAD/DpLcZm7Pb4oStHpxL9bSbVP5lLgmS/FjgHWW2b/I70JY
9A6Op+MR6JDsbsgbOVYg5OknDEUVRQ6M3zBQFNI7smc8V/9ozG4uApupU3Pxqyzb
tZwN6EPdzrsBsXCEJMKxQKlUwwnOB9muZQhfsJRZCHHXrtB6/8l8NK1kPJ9aGd/l
ghyueaFtff2d8gWbv74QAHULytPngDlvXWvRgz/1DWw+RKqW11n6zTP0JPOOaz/K
SIID/pMHAyeQpeaCqMPpOsF3LilQ28kejRLUlrTfMULJqAV38gW73Pr/kAnsHPbQ
Ct8AZvVIoZ3f6fENczgFHdtId/lhdKVz5R6r9j+3KM/QEtKpYf9YcBTl6VdDmz8M
0/4J4FyKibZEfj3dUmXV9UI142oZlvLRxU+Pr3K8JIV6iTxinHTpx9aWMpm9QN+v
BsVd2AsS/mXQnmhlCm6RDVAytqN+qrpLt5s2AZE5buxxYF5/sTC2KlUyxiwRv0O9
0fC3NNxV2Eg7e96D2dl4J0ItGCwb3AkeIshPgS+W3N13c9Xl2jnhV+PvRB612R8B
9wGOtcOLZmed5lQ7LwRM5upandG3/rTh9OsEzss2Gc1x1NOigbsQSxOzGymSHp+t
3Xu2x2/N3RuOqMwR3gNM1IRFOD7W3koRDyYzvW4sx0Vi+tQjia4XqEKcVW47RjLA
ZER0qqU58wx6uzMQDKHufbyMDYUUKk6dwHKM6Cm0II7y2pPwL1DQ4Zm4tQj0PGPm
h9F1RHCi1UROmROM0XvoLj64V2umXoCdNvMBFPvWMRoH/8vrh3xHEXqDUzGKvOmq
kkYJtY3LO6b5xtFY9E7oK8l6bcgkHUV7I3sqgWAunfh11q2Yglpz3wMz7mrnN3+t
9PQu+AYJh0/iKY1WfHiH8wfJtr3+7qIxF3NLmV62CsUYTQc2bxaaXj7zZ0HHDJpE
4S6fyURVByKgk/KuTtdmq6Fn1Se4AhEqEbUnXX3kb6Lssp/Z1Pj4ehOKdcMBuLSc
EPHaHCtDNpMfScXLz475Neil1wPO0vN4e3Y1f6P3BmfBkWCsWHqMFTm7JXCnGmrG
GMmGziK0E7p3nq9N/wPAUFPRtWtnt9Idno6k8xV4RjwPZbYG1/2vimtegTvwXk0C
oMALgqaLlz4jtyR0rtxkbH2+6Fp5UcudKIb3V0MMUNxAYJlLBYF+fw+3Q/kcA7gW
Zkzr1v197sbFr8Qru6oqGVXvIQtYef3xc+mt4oiqwepDAHqIZJuPpe7+oervyg+C
mFVpOlCwEsUvu00Eoi0UC4zItpyzMFMRuGS3acI/g+OBTpQbYXdfkVgJEiudg/gV
YSbI9XyyMwON7v8JODzS3jLJuSV9xk3DBuHGRLvKY/OEJvLdgZAlYuDVBYmtqnJ4
Q9KUdstUlGwUUemhzlGB0W/2jVhTQwLWb1dNwO6ZiKwVbiVXeB7D2L25PXXltOkB
nGJA4/5ssmd0EoUAJxU/jYI8wIiI0gPhI2aYALcW5i7ysc0C1teAT0q04eAkVQNg
MpmD+H7CuNoC5KlI2wd7GBabDIdiqi+ZECNKFRNUS9ObpysG/JwW90BVS6qiCHE1
t6wIkZ/0FGnZvuPWdwSUQIyllXuYVW8whexEMELiG8WorHQqYD0CQ7b4PfEruzq6
XyAvzv68T0fAytqs5ut5R7cWyC/t+r4nceb3Gfdny3A1hylKstSR51jUo8sLdF5y
aYbtyNW1riyl+tISTVMUnL9IJkqLIpT70YTJm1AfNlD+fOiYX5gW1v+PPj86y+S9
Ig7MMK7e8PzOKUxkbtX6Is8xqjFcg+AMEcLeBpiUXZ0QvpNsDMNMXVyqywmUF6tS
/2oCqhR41lJEiBVYFqmGGFHoNwrJQcadNmFYmsTftvb0oLCWphByllQbd0ifE70Q
EPmcoFapFmco7DkmYOtS6R0062M8s++S6USPcDNgtNDMfaepbFhmGvUTXeZdwH3r
1ZdxcElMeyvUWizAxiv5Wi5gjulRLWK7r3w+MP6IfqECGEncgMdjxiEBE8ElX4fb
dWtuXPwrKKEOxaX5mndvRn2qU5JM2oTZX8XV5VUYKb6kgcKW2B41RAeIgw4x2i2F
ACcbRZ8Jkou6DfCqaNLMgk00PhFLAXz6g3rOX3RwnMbmzYZD+GpsC5f+UsiAs6ZQ
fIoufr5HsTAndcVMEYDI+t9wTH/K3nlkahHMuXx/WnuY/PJzntRXXM0jgMZkq6zK
/O4Nj1tzl5Wq0zcJyKJNkPYQuxfWjdxT8Ke6RsBgowkE3zzliR65eHN8afklRuUl
NFORRfZlicJTzJ5FbVh2zKRTPVRWO6zh1xPjynFqhcwc4iBELbcqvgm06eJFD5Bh
tYtSE1DVBTwKhyvbs48aTNbsVLXFHuloLU8O0GAbgvDmrjHFm6aTT3OkE7g+PLjl
uznwAQpsfqy9Ryi68r8tnGT9w4NjSWfhzvlIqwQsA9tmXmhlUlqZUHyScpVeCr37
j7jT7DqUokM54pa/oYE/dsR0E2Dh4Xp8Shcg8tFxK46Wb0e9CDzVOtIH7g3ok8Qr
Ld/BbCR8rM7zwte8M/bVtmkoCbgIgo3FDY9k22UI98AIi8sDspCa81V240DS7LxZ
7IhqI1oJKgQJCH/H9ZEfKP2culmRVsVWiUo6za5pPLr9L9JUFUSN/CT1D6PdNVEX
rAQ5iPA5/nQ0cR090HEEmDnLfIX11sF6JWDgb+aqqHU9gQfcJ8kumuE0zYbTMjBB
O9BXEVHYLUTVmU+jfgnIdTPi86elPm9GGrMQFasI4ezQUbrBj6LRPax0nuPaFyHY
3tnuA/+q29fAb92tnta5g6DYvfPQgpXNbA0HumcgZ19PcKaV4/0QnODgquyq0w6Y
tIwEFwCF3fOlPea2uql3mrtcrsT+pD0BF2Xu7MCOoJaGD+ItWyDwP9H/JfbpcF9a
KfbKAbDGcKjWzS5RNPR7jUFfsIEe1c63gS/IcLjMuEqKVBdwj8QUuPSrRvLvfi1P
3vCBiZ5cQ4lZtNKMeQBKKzv65wIpraTJUjF/p/qSHhAiRQY871VYv6F6V2empGqx
9b1LkRbCzbcWiQVl/xsPurDxxC6zrYnd3v+24M85cuSztXJrrieK3F5lCrHWoUtH
S6pNYowUDe2itAC8Bf6yBy1/VgSZD3tNFzB8dVQ6e24eKFSA5c++W1x8/NydQC/X
bjhl03XOqbKoPPrhBcWZB9zt880izaZOx9ZF8yTizjb47VwOTnOKCWpTZqxW8+NV
NR2+e77mwZNnfvJdptCNOdbDl2smFJiFsqmvlcZBQwrvrDHkNro2HRp8GJLkh+iK
d7gFdfrMrms15BUUzj3UDPGyEsI2u4h6zrOUAuGE9TkPCHTwO5oYKHUn7aZEsH4m
IWil1WFVGV/bl7w/KFRyUDzTvkpQ/lZ8LnKjDMdGf4GJn8iI9OaJE5IZitOb63/2
XyXlkvpK659CAsaplFZjq9Ai+Cfnri0ze995HjHec1L6LF3PAGbk0zaUELRRFPZf
hpPuvcDgQrGRLhL6HCY+tBr8lHnwANeNWVKQMPaOzlGG8AvznI81RYXeL8Su3kT2
dkLUV2yrVYEfWpEGRWI0c3bYufSVAaVvAAFkRW8TriDNRH/QwAm9rTgOC8ppCSsL
P/hBSFMuCwTdNhLdBK6Oke6A0rmGg8nkoNzgoqiNjiZAUrxx4eyR6jy9y3OiBUR1
DsPoUAWovHJpWsdjyNJlyNQKEV9IgsbWw0QJar5nuCvXwf6zAzL8yKP2sd1c75DO
0Eieeh/vGsDeFKghLUWprS02wdIW33+Z97ellhr8VWM6voCOQhYG2o9rj65QOXs/
vevh/BHqDpdZWYyMKzj9cAqfl+4QTUCKu2+JlnlIiJMJaV1H0hZ364gmGgyvLMpx
IRfXnE/X3s54slIGXgNvs/0CHfz7IAuoofB3Wrau1i8Ax7ug7uyJBmStMFYD51KT
Ipyl4ETEpGAQTNPnJq+sHPcCGjlf4oc26LNoopgo5sU30uAky11iZNqiAQ8JIO5c
5d5JvM8EW6ldK7htg+rcKmrgRpl+Nr4paYK9eu55KI/16Nd9R61Jo3E7Rf4eW1Xw
pSponJlpvqbEgYzNfvpsgZXsN6UmuAeTNpuSHvRn7wi6Jr23wbXGulF0psIe8KvD
BsLUGj+upzhMZRwSqkmHNEJfi5q2oyF27mtp7OLJNyPSCcb78Kd6SlJ+LpchH93h
nkXpbQKVUMdVuaa0ga6VBPrAlA3eJMmMONqp2P2YOQq4xFFAdMADBmHdMF9X0a8Y
Uumpeao7kcBM/kUzF6VihApgtgHhubLMquuwft+RXaCkpOz4jtbXS3NTTtD+roFQ
iGk8AjN5E1913V6A3hd+CBrSsgiHUFpkhuXPi5U+WfWbGsl61Vdkmqm102pkt1Or
lrQ1Lo5KFduyZaAsGdQRHIEn/6c5/mBJXjSOvslP031mg9MQKAJxkgt8U35PPlDX
4a6+ksPJTJih4SN6N7sdJqqv5dYNah/vsgJqCWOPiuAHc2BFZx7k5P8tk9OLKPnY
/DCHjVYY1CTg1ausM2RF2rc5t3YiwNx6oYkXz9k/u44NUpTH0Zer462dWSIZiaZe
zbKoLPxDPn6/5X2CATLD2x80u2ME8AqqzWAwFqYivXqj5yGtYbe+/jwMdrf4BA2N
efLdydQWC9N1K2Bp2tBUaeiR9dmtDw4uJfNhvWKXqOf8AGabHvRPMRLvK+lyg3ON
5fwRTRmSxoUf4XyFopCqwZssRyi7vl1zgVxzMR4viy+ysSof7I7ny/RJkVOcLnDJ
dX+v+Bb9LcYtwkYJ4eM0ovXYICWVVemb2acOoxdZqTtZCsUb000txAnAqIMuHSX4
HBMWHfHk23MHL2h4vI9dh/lLu7J8Ul0cvqbWYo6IYahp79/QQL0IHVygRutDtGJQ
L8Rnd83GIoalV6lpJStOBYHEolm3SlmuWBragISDHuIMsaEmSgN/fqlvcnuvKGG9
cTMocSsCwdXS5gpIyo4kEpPpmQlrkJMnEd9EAWrtHxmbWjiNsjJdJVl9X+ZNVDRk
XluhyUJEUaN5P9/PCo8mbycM0qYV7/JB4XxJ3ex4N9SmtrrHLn0d7Dt4Mll5Or6J
KBqhceGXet5zwVlZtFjH2O7xj26zM211gY0QPvrQ0r/4ly9J0ueoDPol7oIEZYlv
PgTgxyu6sGBs2yT1coWHWMEJrs1yrjQ9w4yUc+/fbdVSIjGSWMcHqVOc35d2ojI3
Nn/99/NqlsVrAmv8HVxrarCd9QkF/mnvhf6xfdXM/oOgJ0qmfmYqkJGPwOaQbPDD
PIDtRx3YvyiKRvBwwQwfocG/YPfBSQsc9OXRw344R24GAzwHVtNh0fRrDZW6+u2Y
RxtR3mrzr5FYE8Lb23RI0sfC2usw7HnoB46w9zJp8Sxc3dvA3gZipUQUEUdQ8hBM
OBgcSgFOjkFPAXFFtjMpJIOZHmZLGsWPpRreg/rU7OjJJt7HZaF6n2Sa8zgzxT4e
LSWOzkpSiRmNmfIP8wYJDUKlmq5ssdKArJvF3wwFWWcgR6jTo45W3/End4Zo/y4j
vqfVkAG3WNamj34EqkKkqvqVrZmIOvpHow28HfuSq1zQmUY/QYv0q51WG0fDFCiY
1rRLJKemaDjbj1Woq7UcRKg4i06qJ+H4SyJn2XWUx8Nxmg3MvypJ7gaiH4mwxPAJ
7WV3tpJCwCPpxp3fvu52ZAzQti+jahS6gKi2W6DLoJE6e1bY0NSFlPCy2BrO6z7/
0wRolFr+5COe++h+KrL8sTkXZ8fEH7XqXWrK+pOOXv6TPNRbLlHapyXBZ7XeL6Mc
QYoBcSd7jHX7PjudQ6Bmfe9gcDj/ZZoPrjOLwnnxyLBIXNpmCBC1wJZ/H53ACHdK
xRCLjKNDaVy5NOXy56uHtSsZUpHrjRiqUdo0qEZbrJkbJK0Phs3lPjcTC96l1f/p
haATaZ6zfUFUb1TweFIYP36BT6u7o5hhSJFpiLIlAbOFG2s3xZCVP1CNLHQDxTVy
Y3li/yOOPNAbcPe9Mp/2whLbqGThf/1MWeGoKlwUK6C4gThCqHX/+/HevMN+uamr
TsvWa9vebgvpgkkjIyd0Bgr8UFqN2nanwZLCVXc2kV/W2J4eB0pZD3X9CtyjPKgp
MMsydruTUuT0xtpo2ILqP4TmJNBSJUjNJu+agL9Qk5OcvJzsoFGe10yMow9wbLic
8Fy2/UtFb9DMiexsNH+H5mTM5agmPMSvr+n2zXkd7EVoVVw25n7cbzPjvk1Briio
lJyHPge6fVuBg9QaTBHBtCqpZ+LdNXDX5iN+xxD91rpgv8mJq3n63GNj1zMKTqtQ
vJOVdF+jCAvjhG2zR7yj4TNF8MxgKn+0j6LG5ipJGPigYWOT51VbK3xSFPdNa8gD
/IlqQ5CY8/hsaukiRZL0Ozhuz/dGBH51HGQj1Y1drOzM29ucV+uQdqS7Z9liDpCX
Rx6t+PR31Fg6v3gltYeVm3iTfgx25JnjBuBAVTU19Q5RJ1NTSBX09y66DGibNI9P
qiO/+tMgFqEw8hjqmQOGxCmila9c9+3M8R159svGTiNvyeV76X4mFvtTl8WYEZZU
qrUTXNvU7z2Nu4qT/Mtr9bqsKrCHaxslEJzXaKD284CyDiB4NCBrBvUNK+AHAXNa
mNc5yG3Of9dfCLR2B/YNsQBCw1pkgk3/hSOOAZunY9LLYUbDDWelL632/DSQnPZc
XR8Ixbq2qMUsnrBHX/mp61p4KQNsBX2x59fU8XV+wFkKnu9FJWh8ty/ln3Qb5xVb
pwPLxqOVOnwa0lTeQtHfdK6C2P6nfglaanrbOQDoIfxlm3kZQKav6LlCqXC7dCXc
rN5i0/i88YruaRjW8JRVtKGJAMf7Z19nNKUYNgORVxlvNsPIzgRoLOTKUWKqKiIs
JiZd0wOXaWHrRrtjxDy5Yzmhgpbkn/abKIxc97k8FfOuWXReM3UuF608+U9pComD
UI0CPgpibpxp2eLSiYB/PyS/5Ept7WiUc7lsDfnKpx5aDbtIfUaF45nTnSNBJMhf
0zhP3c4FesSPnn5HXSFqGTFCxON3Mv9mu+UzTizBe2OQ3GfQbSERsaUX30Z2/Jvd
Y/Ee0RaoGUL6XvJ1IH6FFAuyk72tHWZRrmGVOY0fQc9r1iZCm9R/5JripCnjbF/p
1ORzgObPcYU40CPhkTaO4G1BKA1iApL+SYKG+W9xLEX3v4NplCQU6rTnUelbbwGs
RJwWV7XtAQCuAIbmK+vAuRIUAiUPjh25OrFyTsR1r7nqNs59+L6VWVRu9YG9tpMh
zpAfTvxNTSLpLyduLzikrM/NwSvll0Avh0gIBD6h06bkA1/2tlnTINqaGH67q+yR
4HWNdKfeNjWBQ+SVgaNwlgAnHJXrdX8S4ejBpYYvjeRBTTq3FPC914bV1KKnwRn8
rANJ45ot7dYaG7pNe1zU6orMe5K7i58mNe5S1fbIWbOob28ovtn13f7+r8lbJZ+V
FsGtWMFwXy8yJdpI96L7x6vCeo+7m2QuJoQnEUp5EB2Y7DFjApiTVllBXGQQ5QTX
u6T9kaDwcUYaNtGVODnPDFtOjiw2bZfDX+/dQDci8jZb6DzLYoZFi7iach9tlHxW
+h+mW+RjBOHRWPI5Fw9HRjPhbk9kL+aXYFRhNlknLCNeQZUpzQKZQcxL0y0Js+V1
ca1nPo7mfeT2z0ZiJ0D9Hu2kgxnWHxoF5Izd5TSTIfGlkRK6CYwjvEMbX0989kru
z0oHy4q34gJ9cJKzVQaO7MFpt5bjZVHdBQKYUuozZ9/ZxTrSGGHNwMZZOqDfa1g5
s6dqcWF0LaqJydDaHtAlT8xI+1ZOJGov2zhwodl0ah0rTaHEAK+sV7b42Ht2Qv82
a/kCWHMcDC+9PK5RWIl5HsdB/Ijss3aZXnq/Y7o3Sw4wJLYnwx+Lk+EbUZjIUcA6
aX/CpJPBMkUV/slRCaQjmaJGyh/0DQn2BFjK92bmZ1nvqYYcUUcPnLYiwPTm47Jy
/kbZ/a+HXJJc32yUlJE0nKnLNA9gQ5HwI9+WAq6AKsVjWZi9wb0RygydyD9WWafP
2rihrHBUXSbkx2E/roKrEL4mZOvYPFuyZqA5KZauLdBTGxauibf1EovjMMOEKAHC
mzrP8DJUhauwx2MTGhCTbF87IjpssS/BaiIXnh/J59Hsgp/LrYqZMv18i3jO6zz9
6G4XwGibFZ+uTxmb8yUwGTXiCGkwpZ6vs/q6yvwIxHh0FcZGPoEEai0x85Ua33PD
f8VNPHz8aIl/ktKKvcwTm5Xh9mRF8l867clrFPSW/Q1e+hlGKnRFQFbKGImZ/I/8
lMRJgnRF4LxSfqDk2ITvR8yb3U4uPR55IV1K80DhPIYB+tTFfBuf/FlEmohnihUF
uqc93+M+ZxqAJgy3/y3Hbojur6AZn3PhYYT5SXa2JMJwlhQLnwd0c7GoEjcNNc+W
DU8DYC5lfP51CFhZ6aMMCjDOo4Ai/wvuXxp+gQ3KMKOPXDjWTTfawv1kvznYmRHY
T2tmQHWbQpsftiKzHd8lOUfGvvVCCPxkhPZZLRB4dNfvOZL4ofiwyxN7PEnn6s+i
TbsFo+bNkr9nqii9AZVoPS5acWc2P8CHzN2ZBVAp+NxUg4mP0wUzxeIfxs8oDBhy
2Ml4Hi6OdIBvkp3e291JBgCTBzNUXFr11dYdH7aamyJzZgWrHKnBuNqHGUexsai/
t0jcp0GwmJKj40zKMGSc0C1mgvv+ZvUI9TLwFIsTk06cv1GfAk0NtvaMKBdZIzjo
m8Tke4syu9dsKq5kDotMBGjHL2RJdSmDxfNBswAO5wXv9HODtrSyY84KYNFwz0iQ
5LIwHszAmv6kNRRaaq45+xRLfsHhmzIL9Mn/j5EoyDjuCtZUiBp8lr0SYD4B9rBK
96xmwE5Oui8MX1pgdoNDP+d/ZcIUCjjf8ucaGu+sjNjEw/VanK7zmPumINIGe/Lc
TbUhd1YUoMdcUrzLDT7KOGn8yBr6/WG8qhg/OcdvTEjN6jHRWv5UVtBlybzu+DF4
pVk+/D8d1TIJmQXdKFvYH1xqdmau17PxDgHoMXDO5Q8De0u3SLnuLcavU8ERY/Rl
WN/XtvvUEpZUHiKhhNM1BauMDcewh4K89OoKbwIhviyewxfjR0v6YlSvkAQek3t4
48IIw+NGMLka/yZAS31aUP1JCYx9vXGUt997ezzCqdfujmlXC9utI9RjL1T5V2gU
LstN0SYcAVmrZqL/Q8gJX+sHcVLkBrw5PBtZLOTI81rPLsURZoxHhHWvL1CmoN6P
a9MIm8tRXdxJnwEk6NX7xmXCwpxFzf3Djy48VUQackaUw1baVgPwdPATNUoaiUc4
lNBBNtfp3UchDzLpPUGAZvEnl9YADPIp3QiaBkf4IxThQuEEqdyYmC+BORxMX60w
s3vplrzenWuSaycSLoE3YV2EUYc6oHPHBvtB9AUn1rc/4zu5a80io1lM6ZPFT4tg
hAoVsKe7ml0UWjAfr/LGMIEFmnKfsPFCg0bbq8bCAUFkfsZdEvj5epIhll+sMrqi
pOnmj6+hjR1cRPFeZmPWWng3eBrQnFHVst0Py0aGpYMT0i6X54a0kYysUdWPBcSw
sA3BC0JoomRtRKvBB7JaJFREGvuBS3xb0n//GW3GGLGspPVlg1dTFuevNd97Qwnc
aHtM3ZC/XNPA0yWclVk5IpjVGk1dJA3HX3YsyDPTc4eq2vmvjDbektC3ookeCoHb
fi6526GfwyywKc/BCyYXQ4M5kQaOu7GqARnfjK01xU5UflJZTd8RlEYc2KfgDVBJ
z7t8aOkIs2D5Ifn+Rau1sCOzfmEDZVX/RvbL+zQIro9rYuIkfmAIEGeOlPBJpFst
1M6JlKXXl+XCmOel7GaZhzNaI/cbFM6B/2g34Y3YeHljdnmmIuhy9wxnVWZ4Yu1I
nj8G/WpZtybkDTYiNQLC5WeCQWDJkWYUrcpQTVMBrLy1kf9N/z3DXxTtTZ91mZeZ
SqHxT548fhI/2z+1zvBtNhvRuZy+b2FSxxJgDjUr8aQ0U3o5Cy2rqLUifY48UQn5
u47hClrP+uh3mDHrBWjV+YlB9NQe8qS9GY9v6mVeFeJySAO6gDDzxnggEYMbnNFi
rd9jTfBX5yRXFsHTx4BkzGEXGW8W/zbbQ/DUldrjMtLxyuC9sw3EgasCbAfdofqT
MNHi3lMb49bSnyOXT+EBXCapgvufSn7ROn5ZkdaHjL48IiLz/msOxw+CZw1qcq31
+BAOeF37DBa0x4zpnnxGHCxuYmnjvzy919TIQ3ZxyM/4xG40qHjpqVXY+cFGXJnz
yUyQPplI3RqY/zziaugoq4tWgFCrRnPePe9TCmhFyIZe7JGhIuYUI2N3uFfMgDsF
pVnk+pOovra56x9MSw+59wrhjk7ESForNbjUlFXPSZEfVChn+88CfedZTfFdTz8f
R8XoK/TBzIl3OkJbz36ggUOrzRVO1JXp2UiBdDP+nCRTAAMgBgyo9zI5PdkquJld
RsTbi5ZRS2mH3HT6gK+uMok1bd8hJW7V0yjwFK6mOszpBt3C9d12gQQ7kBj+Zvnn
t8Qxm/TUn9HOyKa7wl/Zxm2yggsj3VXaEryAIAIa9761NCFDbrT5ZIyxVveHZf35
0nZylTuwbRCV9CjWsZr90f2daVVcjyh71BKVSFcJPy3gPedtkhr8exhTk9I0JYo/
QFNaVYEBEjT4W+ulRqR+AD5VhglLyWvMjTLoD/mrkvUYlwcH4z8nmngvXgEPqKND
I/WbubZjZ2FFb8I+zojH+KF7nfqvMUkemtf+Pxj5Y4qqS1ZI+0UmD+kUMw+PI7CH
w0VrwBHVqT/Op4O20PVV+qO/EMnTbsnAD3XPJhOY9NjCfxFsppTNAoIfvScR08Q/
7907l9CUhiBQ/V4yiB0G0RYxRibJgkt1lgINMrZwjrXH2bs1rTvRFnKl6kRMKbc7
0zLoy84Ac2jdF/Ap7R/aHG1cyBpPyVYnUZKjk17WjV+RHns+3rHDDU2Zvhhhr/qQ
sgErzhlXa2H9QPMQJnwLJk/bfQPFV4NbS69TCGvPnEy8ck0A4R5rs1vvxHr4N3GB
RVQkVFAVnv4vLN/0Ho3rIbJf73USHQ/Z1X5nTdQk0Q6XWDjvCbeUDA1P6bcdhnne
eqX3GUmqJ5NHQ7Luz+QIKrotG75jl2ydH00ZZOJxEAn57sHNb/x1CP5OqCdRTrNe
558a1IY2ckooU5xbOxRWHUB+iHgNfBvHzuinWH9sQqtKK58pUgtKHLpvKKBuIA1I
XuBumGGeBdkGBgbNACylj5uaGVW5eClKqcylDARI9vWz8liyU2KM7TIKR5LdshZ4
xiC8AqpBoGP4OM6jkOl9/Zise8lCDojg5qW6jS6OYLXbJCoYgdWiJNZWjzF1N+/N
mJvnc14Kc/SJLKZ0+PQM4VXKfCA4C7zmFFbiNWgqmQ6vpBY26mjWyOQ9vg/zFGTR
9A7sAypgGQ/vMSDS+pUtEE2nhLEplrews8f/Y0OXP9hpSD5vtUbw8eVLeY7WiT07
wiNUvFDiK7lEWBAl5dGBTr8kToBHrkp10XhKie7uV22mJccaJfVrJw3jHPteXZDE
LMMrzj6GEJv7n8Plttxz599JHnqPufI6RjkEKKoCD0Sa67e2+tiAIogPicNlTa6Z
R3P+wdvsBDKHjfYsjuEBjLKNa8DK/sS0FOul+8TW/NaJjCrWqQW5FwAdqa3jubOO
vJJGgSz567kO3WE8hn2ETyb/6Hr1pK8xqHAtVFODq4cLcdmu73jk93gVRgxjGHOG
fgHZvVXO7lslB7mabRSAONkALlUJjS0Dk/YBla2E0zu65tZ70q4/t+vJdp12vRDv
+gW1EIUUG2I8kNA42Kt5x33M/pIolDF0ihMx5zG4A5XzeSecNMv2snuvwoqyHz7y
QXm3AIOd7SXagAp0D+e8Iq6NvovQTUfdh6Ie9x9Wo9TS9ARPRcTwH/xIfb93bLpQ
nYQS04bp/EMoQVVqjp88BB4O5+ESemDqnmzCNH6YXl6jIMmL8k228mllkUXV+ebg
c+XlrS0w+OOoDM/GWk7XHr+XVy8ILSxpBgMOMn0CjYLb08bFTiXIp/VsWWcjsT2q
HNbMK+F9W7noFNoPkHTUlM5INbZq6PFXDXIx9B+rigzbdamqhkM6ddbEu2kkmia9
9mKgO7RoGgi5JWQJjfzjyj74neSmZ+iCIRbv+aNcZqIufHv59dbLS3R4MRgYTmY4
JGpAXKr2bth1wcxTATmcEuUwD56k76NBPKDX68yVEZhbjrfJWGuO+z9YH8hXLVrj
zdyyPHfL/sEr24emdelMbBkmsR4/ouf4hiCQFBUwNu0zoM8W8YMGTK8YmFC3RQAu
76SJnaxFlX72Z6UM24UkolKGef9PHjVVmPAwKkGVa+gUgumWTqjJeTHiiRwTdsbe
KJB7ktx5ydNCyrgYFbNrKtdJ9ZTF/lVb2CJoLkoYLB05nQtJNstTXYn+XbxNY1oO
PishgYxkZjXO2mXcSajwDGzBqcAb1/sdFOs6z7iKR+qbfjX3K5kyUodFXA0O58MT
yFOLeKQGXxSmSjiU+dVmZqzX0SY0tkK6ugnvUVy5KXK/mAIyEOqi5KxoLYYCY2m9
dvrmLGENxDBqdTGD65ouD4s8B9gVt3es0YnBQecE78Bxjxi+lKMWrMs2jECsAGij
f5Uhd529gfD4arHvl7T97Y2cSGccosWrjStOigcHSTakeLiq1U5u5OJ2dYjDTZT5
VQVHNfomWTsNorWTNEno6115Ucv78oGPAfUkK5j2wgHok+HnX1UFfIqM1ydM3esr
m2oq9fiF/WExObjfUl9wdCRBTlQqktHJXn6Cd1BQjOPqRxn0JSGdbmVoJMqEv/ZF
uvaPkvgbsnbgdb+DFS3mUdB/rGsQTarEcYkqIvLrfFESuw8ho1qZe9OvQRu+1/nC
HGsTOy2bf8hSY0+tZ31+Oai3ejeBwgbGCyiJOEyR6AcToXiiAYwOnFqRpf8XsYAq
4+7bIjv59J7cJw2DFzBNbVA63dow61LSOTiQ/Mhdgzlc7bl/OXfU17duLDe5gwLK
cqKLwWOQmcT+2jIPLx/NeGt6f40w+PNlc0NQItNV3rwDVwF8c8THOeGwjqAsNqKS
AfCjxp7X7LfpevhmhbJv6cJyuLKjoDI2cX9X84TPLhQASOCYcXTWjO9obIqH/lVm
JgN9Lw8i35p1d+FayHoP2TNp0OXqQUn/wIHM9fGZAWT6L0MP29rsBEMAFHaV4kkh
AJH/haYNxLn5cQN8RtxjPj18m6oECp9jjyK7hyCfWzTdDi3jNtM/WxQtHackqDB7
ZvQ/+v0UNgYSK9dnpz7iqJJzmLSkwgIRkNiAvvRIU/uMCdjXvZT4fXSBIol5zGgs
jtHhOy9bMHzWKoIbtVRFDAvSK8wvv1Lj0en0oJ1Xc9mNZcuo9Dn9jeK4W1BDM5cd
PY3dixr4YjtEu0lDeUwxq72R/kp1skUB7TgXhP0tvOU9dyAnRo06NwK/zEbE7T8f
oWDshmLM/ipqshXxDwZNojCrecNdcOot9a8W5yrtM9hMsH66xhhG46NkQRXCy/F/
AQQc8DyrW3f9jAQbfI8BTOgiyO+yRxrqrOMtKWiI8+7ErCccYlA66O5QF+4NzdHE
yr/5Q3k3/44hysPId3+4fCkfyaqGiNtiXM74uE2evfmHCj0A+NqXRJfTpPBcOO3Y
e0oC44qSZigXaq5M81qfgLGOfX+a/Wb7QzezQU2vArxDLQvko0UW9rb8QeLNFfLh
VN8tdqKJByrZY8IjjzF3bwwM+f86Ea04cDlU3CnuJ12H8UfTBrvaG96dnQlhc5i5
08zZnXfIwPsGogaJTLemsocZ8yEd6ebcBjQHFH6NzeTdFOkq6VFyAsmCZnLHdOO1
NOMbstKjoMqO2+Dnk0w/i3tH332ZLhK2J29/RnSMRqlATHI1ErIMcm8Gntrx6xAP
y9HZPxueWmFdkEzbfJrcG4LF9I0mAfs8IHCBHZ/vsWMQmCTIHODy5+oGTBIjTlTC
v9/xvklkF2GlUP1tbTQbUGjWNzx6OSro5YibyP3+L4WqaX8/7ZXRjrqHyT2C4Q98
WmmW7JC0vmTazpk6e/4WlOil0kOoupPyOYDVTaKfBQFdZaStHOtDUp94i7pO9Nyy
3SQlp+LoFKjiGX3xZEBpNiSQzMdrhMdWslID9aCbiKPJ/FxPlNVCMBygVXQIMA4z
Ez39YZNyr93ZBZ1mrq7HjJ2PJGtFVk8VAoPG6hXYF0SY3ilTX9md3x9tbGk9nlfQ
vPmU29byNMo3SYcD546riBsWjOPxli3mHaEbD/wToj3WlXzJw0+vhTdKTQ9acDgO
aHw95znsY6db2AXWIqM87K14DuokZFPRiizHC8PvMG/S1f6KINKt6QqyvouzKHS+
hXt+ZqSCUFnYhY0PWoujNfn3pX7D0pAQ7NBFNEj3TgeEMObjt69FeXFKk4wus9kU
P7WQ4rCtJx/1m6zpMdATnWse0PdpFx9vajnx4mJdbDAl5KAPM6GAMq/3QtjJOZaK
4NkR4rfnB2HuE1dgnQKV7UwzwFFG80uRKc3sTzuPqxNj7rQbAgsDpwcV1bHHi/58
XS9CY4HgFiJDkztFHYskk7IH5u0AFwUz1zoNVoirtjy21v0vhlEv6UczfFKGEE1A
aISt45cuOhuxsvPRh0BtdYYcHwQc7WqXdM2IcaL4WswkhdUI2C61ze7rpMhKRMov
SCf5LHQHkvVC6LEDQQZwetcln9cvaE6TbjlF5yYwUE/aUl38PYf4eqrbhGfr0fXu
iIc8W6nKWUhn/tl2o3Vwr0HnQIpMCWUMlpUQa/3AYbfGJ8tMLN1X56V/5pxSYgfR
ghBxknIS5OPryMOltXNQK7yDBc8x/sU9qH/5tsl6qliZYO0v6WO0OfvfeIPqq60T
DUe8mj3LhIvO66v6WkNFQV+VlnChiXZHn/JVF36YiOBB/dgUkIjOFQ2jmCfrPxpC
UibX4iDSTJjiLB9W26oBOW0v/jQmiJjhyx8RKy1ynEeA7rdi96hEqXqvpXs4n25W
97FayZQyXKGPfPkO5CRgx5xRyDXjjIIRYFOMtcdVdtRYajvBwZKy74I2t5banTSs
kOP2Xa3pGSHAHqvuOsa0Nvrz5V63cTELLJfTpwuyeKPsofsYFc4kVW04MoGm9gVG
MYKnTyKzK/ssRHOM/7wtqqNe5mldF0IB/imzCxhKU/B/Wr7b4ZPf/O3+fnvZW77+
2udcnfyPjxT4xn8E7MTeg6ZkxN890vJI2OgYSmmIvuhTSEOCWP8hJ3E3SiZQp19P
ioz5dywfaTKzmDvU8fk9QHug896zvcdJe6hpo+Ibz80Ve6Dv15bGWV0Sw6rRrURy
SqNdD01chPX/W98mweV0FomyI57mOgcfL0WMa53ml1whLHlJupt9XiQAezV2j2jb
8LFVzrjh3PDSFbQD0BM3JYUVR7hCnD8agIJK9d/IrZmDX17g4Q30skUgfCiP52rv
Etim4Ah54ZnF4Vh1ykRG3M5rbwuTBxVkEffDaEFo7vQz4y5QAOzfsNbp2AnGWrBi
FjIlbfJAOGLd82YlDNrSdmnGT9M8q29JP8v0YCiX6gVS2m4VAe6aqh/YfouaCY2r
rI7i5EUMPYzHoasRE92RFH2/snvuou8WL2I/afPEl1CZiLHk+fa7TFgRKvbW6TmU
ZYcxXi5yv338gy+W89OaSFsqvdTN5ZnahITctSNKVIvj9tpBKnjbfhm6WTjN437U
yFx9bnJCJ8kcfkTSuMEqqW5ZlV3da1vz7MHEJPLOcd6IX9BV8W7vyCwxzNSSBZ4h
Cq+/LjpC6vLboZYHd8QVixLOEAuVEYCgPWvErkEY/WpHFGJosmL5BEPfzyw3OqHt
Te78J5aVVY/fQF66gE52PpZOrgSvn17inOU63aOdZ/pRbnZPseZLXXrhJYglO2dx
drrGvd2TcpGmGXARTNxypGQ+2VGYV5HxAy7CxdBnnaB244DUYauc+kI5b/RoUKVj
REQU1Wx43tW/ewcKaKRWMaDNd5ttF0AoS72u4erRXwLgixOKwZPaUmhsDUW27AfM
j+aiypxxurbjbuAniVjAAzi6Rzd7pWjTK8rC0UgUSWGBl5zYnBRZicEXc1MQcw6X
ybh6IvEdPeEGdrWFz20xeBWZLGNr2+bAJeUB/7k3eb96VCG0HrkfnMjRNn7vLCyy
EOjkJBQsWT5CQOlTeUfWt+Od4wcbxCs3uJBMe8NlqycxF/bGGIjrolkr2ZYT40WS
vdt4AtIrVeJQtyeVlVQdoVF2L75P1rXZEb4adl+I9XZb3ojEB4Q/mma3LP0VVAP5
od0vU8JE+C4eKDUU7BhrRYChuibvEZvjX9c1wm6ftHGBv32f/rILsJvGa/RYYnfl
FIlwsqkV4gWgpJRGAUNL+j7+nOIKcRexIsBniJnCh+KA7FIZU9ICK7kS3q+HOD9Y
LuM4kNyoS3aJ6NbI4OzG5eAXXlYIr4oV0Tchsziiqdq4dDvqHJDoetbrn0mzkMjr
O7SNeSiotWDlh75ItWIsBHctNan1zHmtBY8wV26UwRxwr84nDflV4V2MzFzkCV4h
NgOFyYmBwTrbuAyHPF2AZLQxD/dwbiWj28GRg3xNNuyDGLQXtlWpYQ3eywsyWXU/
m59d28kqVSGdn4iW+RKlVtWPgECiECCOtS1S5JQTnUnREWorvg6Gvw0x0OGjQTj2
gIfCvU9PFQ0c04/m4sPSt2WmiYjeyNPVHdPfZMAK0cQuBb6ZMXtAfa8/xx/biLzp
h8pLKGaQh0msumX3A65PgLWZlAASdAT8kBwSpZ3Z2DeYhK8VGvL+enQIZAdbtDwF
T0THJlzuWCCL7+kjgB315B9A9XUhJrc58Us4cMIlmRucyNv1HqPg6xmuMyw7fJu/
hYlB+BnaEnGKJG3v8eQ/eA/u4LuiIl4OmNXCTFXQsIcLvLUMG7yqB9SWYIfbCwkP
jb+Gkze+htzwd8+AtwNy01uRwMYPNi955fQz3pbofTAIpmd9I8ZdyakdNDtCjmeU
49WUjLX2hEilKuMQudJ5cR3kh6qdpDGPgL/ogavNTLiBPwfxLSjSl8EWsAPOjMqE
XWuJzir6fviNiVsS6D1+z/P/AgXmJ6pceSBIPqm+aMePWJ5hCvtviK5Ue5Mwm84R
sS6ifWoH92fWjjaGOjguIQri0FdCpPv6r51y/XcQOG2Gz0Me/XN8wa0zTALp7Elf
d7iep2Hv8ZwprSCeq7kDeuemSVPxtFwL+sMDDRr36LHRpLKNEVWG4wCHp3rm//Iq
X9MyShXR6mT3TXQLGotIlYUCJtV6IGIQtBFUVW6vNk3Zq//qI1EWUE9u1FFRIuIz
WahIK2Pgpb/3seM6jWxfN7DhZj+i1EcY3NzkfOAjV89VcWvgE18yg4az4paQ1tsg
voMzVcyp1CDdilAyTgVKnL0LJbS5Pgp5inJyk9dYCramsn33G+Eof+OJtPaxfGAM
cNabl59TvC5M2gLDLyXwfp1XTonK5d3vPya0mgz2FKlPTUg9/Bys29ARMi6eRM1K
PaYynSrTenGpBQJJigP2f2hMSBdB6Dt8X1pocPMYSdaG/DEcyLLFZ2pPhBnzjs4w
JOAY+jMrs32S0wlyeHyzxPvdxkSVCH573Wen6NinfDp1W20zC1jJopmGNMdk3AVH
azQE7whlGoIJVFCoBjbK5+aElxAf4bfw1AOPBABTp2RrHKyop+igHpGnZm8S+hUV
/peiWrnaSLE9rxsT3tAxJzZ8RiLpRPRklZFi75493u1TJkDOLHMBT2i2EjyPS1jV
d5A+VUmi+l3MenmeM9CkkNvr2z3Izp9u56E7qdWbzSyfwlajitgxLgxmy5iN2/Si
em2sXlOGW8JimjeJh3ifNGYf7xqy/+3Vu1srZwMPTnnBQzdBy4rAQaIPeSFCAKBa
lXdc/dMbrDUlf7rE+DZNfx9d+pxJyCTbT1Hl/KJEQIROgASq+z9+c8TqDzJquy7J
7cbNlxr2iy9r5+3byEC7AEEcmic3LC0LW0jbq6cd+PnlYWb0DT9+zS315EGTyAzs
NAEcVqoexmUaRCZTmIkZfLAQFwNvooyMMFCwV7M0DwFC7SWaMi+QCoU0fgPPBixk
dDzd8hi9Gjgyx2rszlayhBHZD3aWEkLEyDdzG2DzgOnA88x75UjJNRPcMD2Z9Jkl
oy5r0kcVCy53gKNamdmlvnGfUwGNjvlroxr7u33gpSbpjU2xEV/Iwktw028sGN83
Dx6gflyEdRvBEtABJF3rzs4ezGoM9XjgcC26YEyXxQfQGFJZZwGKGuYytcIu8Mwb
6zKHYysNjtfZeBiWUKQW0iUNcN6FZMBUl9ZPG0jZ+dtO6LYiZKg+5uW2G4paPeTF
QD1tWDNcbS2qSzUmyxuTmMJjxiGkSCXyoJ+cTVtJfQ5WmgZfuasz90jPlcPQIsA3
lpNrUJmfryA6ZEpbjvYw5aGWhfvsRrlMLCp3sfcn93ccSsSrzkJ2CVtPChoZGCxl
bZQYAsRWyeNjav0d2TSTZTWbHfxcpFI80yRKEG/TOKvFdtmPmeVMK8O8OzqGeewt
9s8nOMZAkj1DWzEo32L1gFAWVVPhnvb5DSZYLO9fxhlGsypM0072ZMwQQTPg17AC
yVikJ5g+j59kZVdTmmW5SQMbUEknrAGf3wrq9KgTs727uI8NtmoQsfxgvFGG1C/R
bLEEhQPrXbjuTM9l13YSPcHPg+t0ovuVVVuDdeRvHxGtb3s2KRW7Y6uY5671+bGc
5uUmCwFVxCH4AIg/DcmmU11ddOIP7axnL0ytCwXKWb55ETAVkk/uFnL0rM5J6hlR
gsF1ArtQsOJONXudnFqK2OBUaN8w3j+hvX2ggEnfkfRImh00im7bCrp7/xwTnWZ+
QSuceTUFR5atbLy9W+24MkTSB7wZSWq24HwnO7ZG7GCCq1kU8/Oki3kM7RON2XJh
VALxb/zxuT0x3+iFC+tnXRoHrK4OvpCaFxjSIqMEWDEvmksvoiu1gSCk+rwCYvCq
rB7veFjCZBA8DXIefWv4QaFxGy5Zjzvi5mIf7sukJdxTdIa64QPvqHyA9LKB5YF0
yuRbMQiIKgxDQFidouRKEFDQxK/b2tzuMK27VUdihRNQ6qeSzRTPJCXST+NV0oru
TzPJrg2ZtE/tImzlRPDaCy+O4/WICkxtKXjvYlw6nifdY3dwWDOEVV/sglnmNm3H
eOTcHn/aJXAcZBnC9Z+86uPaXO4M74QwVS6V2IFVsBWTrJODnd6kPOQ6pndECMD0
nSQ34GnrdEisYZwB5ruz8FeEPMTHfi56VCz2Dw+3B5/NOIGPySGolKKM49wiXQGl
P/AhqAMZt1/u8LTMQY9gulAoVW0Al5fDxq7Vb+R2BZUZHPSA/rz50Cjj1d4AWZki
Itosv+3HVZWCCS4ImPk6QOAKOVzXMW50U9FS5pxUlcDoiw4KGWqtOg3zLxQQ1jNh
moneMW83jXIodfnj8mAM7s4FIx3QpNpUybkxonjGmTyDRNAIzt95DxwSMp0SD56M
z2SGf59Q5PAxxnqoeWMne9XAPay3m4WxTjqPJkNQVEMepzvwQFmlETssGBSzu4ld
XDyDb8n4eEpwi3w8bQIuL0ZvIxZnnRUPY4YryH5Hpi+633fNKZVU5QiexT8FLLnt
UU8aa8yWWXnsNpqZoaa9vSUEXHSdSj3IPSD0CzOpUc+SuQ6fMzHW/yegDL5W8lTx
+qqdVpSJBHqMD9Kvl1CXeAp7ddTpgUb/vjPXPzzbwjFQX3+tcBc9re84dTgmBEfY
E7EKLtdbYm5IUfx4kdx29uve9oemMownS+4ukTUIwy345MNMWFIKfwd+GVU9qXoY
+EKp25qduMb5bR69u19A4XveGbmvlM58vp3fM0tRaFiAQ31o/r1lRSTLuR8V++Xd
bogXTsOZKqLtuDFulQfs8cxWnkJsYHtLoXJ5HH8GOBQR8CilJWXwyT5QlNHFS1W/
Wq4meUcKS5O2Aifap/Gx/aTRr+Y/RTgy4eYENsCHvg3n3ZAe+sraaUxZDk7Gd1Xn
gyo8BGoklMBEgrrZEGiVO9szZOeK9WAWLYaAC8CvdwjmSQZdOWOyRm9eFGSoB/Ds
8d8fBcop6lTdF4FSNTkuXzwu18xRPWZt6gtEyIjcI9np07x0mIR2eLj0rnGiZNE+
3ACdwnLotZ7C6jdd2eqqbXDdmjU/Jh6YxSqwkp7xLs+Ez3E/d2G4WgSAB/tOU/nk
mS0AGjP9soh2nihpjrK4sjSnWrAIAiw6TtF0xNtcmmvzCBVIwskSpuZQ4yBOsSGb
Iirl8MrBN/d5xQwMeo4rlxdtwcyDtfXu27VoijdpcF/d8sndajUQTrQ+dDDoEM3P
G4bW9hie9ujBNA7I2JMSC9tm7UUTKjRcZ3RTv6COAHOjJecAfMcLEesOm/q3iDQG
GG7w8tqUVVlC8B+YOrrdo0mBzvHqf00guMyWap+yT+hD+yUeVoerMlmpS82+yJp7
9S5J0IUlf/LW7gMU+mlPrK5YFF6pufYJeTJiwTmhzcVG9xXK4CxegF8We9lwDtFK
vqi/mim+vzQpmXCdl9+4Owf8fN/EsRNTuFFgJWeKb9CAYCGeZBrcubl8m/QCrCMb
QNHm/GufmEeNl9/ujA3RZNbHXZt70rkAntCgHzL3ezAPUieQd41ht+lYztqJdKzK
92rnreFwOkh80uAXxp9/wgwHwOILYEtY2loIGx7sk8iC3kik8NmjDMlM5q+y0T2T
SzDN6hBKvqiGJls5HTDlUVJV5Kup9IgFr/F63f7gOudUixZbmIdco7BNfWVRqzzA
l4blKRyyfhXNlFv9Q8QFjrciD1KL5iSFcInHa2QEY4FbADScIkVoLqxK3pR3px36
BPM0Z/jRbacbbRCJ+kdO2lRS4oMeF1ivXlTUTNWsK1f5vRAmCy40pe9HzT9W7A0J
7HwSgwggBpAbRr73rf2tU1j5BICb7aFNqDlxnWrrOrHCHrjM0V16/7G947OaxOrd
SDD3S/myIUta9lP6szeVwtI43Olf47wfzD8KTzBoIgybkooCyfLs2W2wr9wXsUr7
kE/vF6Z8giL1ezqxUnOb3ic7XCllTEbrspFeNIaVIxWCt875jMS4mR44hE1efeIo
uOkdjr1J54Oqu7JJPmCL+TPn+VcxdGffnP5xpUAI8WBLmUUReECBZ8jTs+dfleg3
0BuZHA5W16Jsw7+V/YDoM0Ltj0T0y0MiDf/4nEcU2NuO3EO8+fZlID9zbbpaD2s2
bl/D02sBTt/8wJeh6uQP2DXycB4CxbsNrKPb1mxq9RGoKpxSTXG1Oz2k3YYlyAVP
xm2+FQnHRVmJJ2VFOPLEQ3uEYbpDuPD3aMdbrKfMlhcCvhoQU7YRT+z3D/0JOwRo
vnOs2WlAs4ZyoBY5rAQO3w6Jb77fLUqAkxj3q0YOS1q7yROXLfuOFO1arSOKLSqA
R0OYZCAzdPL9XTTaWKT4F+gad6r39/WvhAw7HXcRKbPzpXkSMMlqyGHATUWLA8qS
ok6tlc+vOAeQj0r6f5gYE+swOi/XHwqxrOEtRGQMQEVxKYI2MOLL9n3kkLT6pbWv
9aXXHebs5qkKGPRief+QF1COLZz6CWoUAosQa8l7bAkjtO+z/iR1+bz9uuQWGrQb
hu2AMelSa8hk6DYlB1em0Ln2UdzYyLXP6cbyV9j+jIm0s4F/Zp/4kP/OHW5eyUuz
vrCvGmGTNsAEOs13KuZkef8dyHd3ZDX5//+HIY9JDoOz/zqKxHw8kLvP36UwO0tV
JIuFvkg5J9kx5TJ9BHS4nv0IQFzFRZmFtMDYP1XlQMkhFJ2NgqyA6MuEHRNBnL9q
HU6q2JyUuxD9jo7AGWc4G8Z3UVrEmy1cqk5ll1yEYLyAYBcHMzlfTXe7zsFDBXv5
pnNQXJeEK4UrHQ++VKg7zD6KOigbLgt7okulb7ZdIec7W73lo43URMw203xWhrxr
THHmf953JcsZEnWNUdoy2t8oZvcd63+ToQ0N+hGtqSw2/uEFBOwGV5T1ROx26Dxh
bLvrvqHX69Neg0ufZYWyC+iij/n3iKovjV1KVD2yCck+n+AQOkG8l5Uh0+vTE6qJ
H6zl3JTmti0c7FAyZoOpdWiHoJAKDuuvVLSeYbKvXKqRMZ2bLz6vGC+YHR9G71bP
4RUl2V8UmmE2OjznqJehblY4DYN26bO2+pLeqMXD5YnOzt2EWW0uWsm5S9QtlHes
IUbQDOggNpkUSOkVrZq7XGyy2jR5bErgP0xgEELIfS0hjKfdP2c20SphaoWtk98N
3jq9AQoFaN7oC5p/J0ecBIO89xBE9gukb46md3e9kErX6vUbLbsrLrl0b/DLKagl
5H+H69gPQNctE8YDJ8M9eVlrmvcZybtXvUqgMBJ0BwRwUyQqXXqbzWYaVXRNXdA+
CiXX4aKbNoMwFhBUIbxeLfVxq+joLgMKdQMyIR+qvTuK4OpCY+AUdKxzE75zMGdm
E+GZ7mZcQuTGLRnriMdool5RKEAOg7RKbejnBiKCaiiG4r6FK4ytstvIA80087Qy
earhPhcE/t88zr3uzaEunbiYRb3fzRh0Cn7adr6Jdm/3Z5mcwYC4rfExBwwGWDeO
gWtrxt1mMWmqzaoZx+WDpMzadAL3yrB+lwL0cQgRo7QwEnlFlBvuuyPEuuovdiJh
1S9r44pnZUxLBygemDb7S7AIoqWF1Mz5p8FBhw9nZ0vLofo3OoiI7Wmo4/CeMEXn
UJE/K4w7pffnutRQ+4glJKs0KbCv88gW/ssBOMy8SRJQ/uU4K0QJceXQWz50YVe8
uj88SaWBf3Uq6fuB5AVUZfgsIC680VOZjqiMQwUKWUsPY457ipgHgzjeaMJzgE9x
tchsbeI3NqQUSFkIlJWFzj++EhrW3aB9JMV6aLkxObPclXjGualyW9X9bYpklpYO
341JueQPCo08CtvgAZljdoZm4jj83RPltRTp7ImXHEfEW8M9K1WZMeiBK9ocj/Jh
j15l0FYcQD4GkkC762s0SMlU2MRYOrObrbtCiMJqsQv1ZJ9IQPqf4cmBvpmcEE8p
21XW034MPMVhV+Z1ik/n1xusEtzPmn87q1YJ1M8j5B69OWwdI0THAmoPgc3nJX2t
j69sFaikHS+prAidxwUTZ82SqVPptkr6cBVvI6HD5NShw4PS0MqFaS7P02VASkXT
jXCL6fVS9YDtxYn3GpmdST5YQnTgzdLEvZDyOpjb85J90G5ltXzGuigdY76ejAdE
v8ctTyN+WxUMRRhwxIjjnd72Q0RtyBiBiRw/ISUSGYdVYT8A+dV9bnS+CKj6BRSP
KVu4x37muM7r5ZvFGZGE242isqrp/uHo2ZjPF2dxycn6vpiR7KkmZPyUcsxUbxyx
NVuOriLkQZ5MRJNxZ1QBXEz8+VhYvKM6kfKzhOLQanZjmeITPxSkiJeCbGELfXmD
Q7DdkzWnQGTAhQykibzPwcgp4ARRnmvnia07u7UWl3tAwY7d3c2bK0dts+0rOSDf
KDz7DE0ycyJwckO9snD8sESd9zHR6vZ2Z1Kti8mLBhapxm/2MKn958aOA7jvWa/8
0xIobszS5dQheLO6ynVhPmIRb9kZU2VWT8iJRUPnhHLTqFqDu5NZoV5fgT+jDkWe
zHlCrjGcMI0WVj+ECq9i8YmG/WWDdhn/MaLmW5dBq0e7JVi653LCGmxnQQUd2iU4
EnLk6FvnSXjWKZ/pVLJ6Ctv2IHk4qqayag2y9yhZFoBfM3R+s0lv4iZePVHmbdxO
COy2ZgOiWOiGwVerdJSB7+pOdScTyiXkkSPh536Hj1BsMSngXDPC87AnhxXhf28o
biWn7Y3iiidZCqdIuUkndkAbwLzqpOgfnGRHeY0a78JEhR+LTBHIXwIbNdYVicE9
97Pv9L3G2rsenb/QRG1nA7DBqOkG+K0WSjmOKUFbHyNytipq5KibW2llY0ooIhh8
Z2WPPXvoImjFI0tcOJtDFEzHRhV33l6w8RE1UwQX5hWFxSPWibsnDqlRH5jGvch4
7u+oEi7j/GHtEEutVYosKlnQC+s+fA81aCvgkMcB2+OOXGzRnfg6VgEBtqJEK50V
rpLQUigsbb38Oz9gqKfkwbGcSWpTFInmfCBalWVEJwBpHGxgTzk2KyWBIdbZ0gU5
Lvh9J7JI9EXB8KW4ct53AmpR4BYjhFSzwW1wYGQRw0fPVO6bL+dG83ngPNNGcvz+
xS4kWWZ8TYniDHLtbSaAxASlNxyOFLSICOHnlff7hyhIi5udmFaWiHZRRF8zBgmA
ABlO3daYFbORP8WrQNpebCIbHKkiY9W8vJ4hWn/j35dpEVdnCM6mSmcQafsdLLdQ
gXWZ6KIhYJSZukZ0JtEmjxF0mwdkMXdh1RtV8uC3rGKxxchzcPTo7RSnhWm1NQdI
/yjO37tEEm/o//NY8HzH80rUovG3iPZWrcZo0ZmRrIfCcMOV7Z4EnXIjXLD8bNeZ
1nCnGsRHZ2qSEXrzhkeeUT+OjHaXlc/9IvbXrW7PB+8npIsUuQEZdV61YzlN2vBv
udD7e78Tk3hu/f7J3MkkH0H3zrDSY50adWydSxhhIT3CcPf1nxrgtQ2l7D+52WdJ
zOc5l56Hy55zX/X61nHi8INDFgFMFlbhrJScbMRctKWmaLG01fuQCtd3tIDjP/Wk
UdIPFXNqoznQ7tlSa9Wsgy0Y7WEM/07g1k4V8gUiRH6ZDz0ilMqv698+xeNDX6uA
WCZnHp4jjSVmZcCRilyV/funmhteZlLP5FYDnn5tTKH586pAa3Miqn/G711jBH5s
7HvZ9/UK0/FHSN+6OYwbqGy3rGT1yLi+t5qSgq9pQ+HmCQRItPA8kdZal6QpYp3y
FjKrzw16Mx4+LAT2iNFcCYspVRWCmS0s89lNuP97kghPq4DmFugF6HeDhbn1ptLu
M7gBmtCm1+LH7g5bP3Y77eQCGrOA0W5plZQedWcsMVQtilNkSUa8Rn2ODVMTl9ZU
/k9thuagSSzcbilUzRL3W0ACXknMx6YVXnscgVmNEPHCkXmfb14Pg0wOjQhrPjkU
ELuOI40k/B9K2B2iKKoMxDqnXcfx8dcJ1me9oDi0xQdJM3NgNMsmMhyqgRyHgQ8M
msHBYpaNMUHAE2VEilIYRVUjiedx4BBEzb2vPc4l8404+XdOQO46MWH6i5ETv0Ze
B8Vo9OTvz0LLk3ZrJYwmeyKGpBvWQYci8k1ugJwOf+QmjzVdbu8/ID6+UCX+Wa9K
cLkXg8CrnKp4FEWsdLwr//+5w1Qvr7jdHwOqmdMmxVS/k1DFcP+yIBcGOLpwT82L
KQe/WlWXWO+LKHMsUGjyDPfTCETqvyW5aMxbcmDbe6Wn2wn8fE+I4Hni1u/QTEc1
MsF05pdpW9wuDIW2s9EIHmVrr4ToLUqTJl+L0mpNCaG6k7jGwXqgjadomY9mvYG3
MLRxPEtGQ1Neqb1rQwzwKt6//Ik6npaSLRmbvRyeCzdh1meUZ1CWG6/978urCkWX
pScRcTxdoLgwdijf8M6l+6MYr5OCXrnaBmNB/j677UpnZrU6JDRcikhjiBgW2Oco
XFXMRiteHP99tz7dyI9O0U7vDyyA4HRPp70D8zSTF0wTSCVI4t1UKw7PxNMkmqYP
fBUQ/5WTOrcn1M+hvdq1IDjhwUDyytBVjZXZVjzcBSz9Fg+KecphMBDCWtOvfaR6
+BQv2BULtXxFYkRMU+sL4N1c54OIiK2YXl5KY1pGIWULR6fNw8SUy0G1QLuBc+QC
Nk7s0fDQ8Y3PiRa1/skONmlmRHdshdvB/xaDxRKcgoHu8J2UX5bQSS8m4MZq8FJ2
HFbRY9K/I8nXQawLXaJ6irOjDzVQj0qq1NG2+F7dldETzsgXjoOhQxkc1RHkR63O
g7NriaojZvzdzKxg3AjPwdszpHqh4RY0DJfI31CSd1dGaw2RituuNSG73DYk3IaF
IeGtXucnjuXc28Z/xV8QyRBw+UsSkFIVJu6RpRSaeV0EQq/KGaSeBDFxWKM06CHE
CAh36SriifDhO/7jWv1XlJCB20Dui52E9cu4snj5WdHP7w1oLRFcFvXmqXqMYyX5
H3RRp2pQ52JOxys4Mufnpz65QYKiQXG7H/EIAzM8U5GhAZBWbN6a0oZBI4H+HJud
vRO1MdnZAjvvcrWICykr6mw+Je5ZDT3UKoJnyNsYYU/S9TRUKjvGQ6QBZjHne3yN
/8D2cm/xhdIO/5hkjbG0ZAS8q2Oy+EG/PVUgE3umzZD99PJCFX1KNF7z9XyjxAgn
E59GfDWRqEL+dhZg/XftG3DEgKaV0jn5SwqdvFmMwJ6Ou/DTq1GtNIjLnfTpUf1G
vcXrxQ1MUYhmxkghdNhCsaEHnFs4d6+0CeaP2wfnKq3UL9jAYAYmXSw9tebUiIGA
uwjb4OxIXAp5uJKLmDDhQNGf2tivi0TvI2k2Z4z86AYAdu/3v+a7C0H0lY4Q8W2+
SqcosOw68dKeN6hle9Fg1M/qSlT9C5dWclF5hqGGkcaVzHGePPxRcDnYeRXSQgZa
z0d++1JzUOAD+xfiYI1ixKM2Hhib1Fm8+xS/Fpq/vtbFQKG4Lta1fz2zlhVoJDJ7
CQOgx+cJ6KDVsxPicQPwi2d5cA2e5K699YBG+EBdsJUyQPhQpku5kSt7SaXD7PhY
zZmW361m/i4IVcQQXAligiJ0nY0F3keBzwl5Vl9NxS8xFzoA177KFL+0w79uFsse
XAYV8qCcr/1eef1GvXHMi5ylGQ9voZnZTdiQGh4JcsEJGLRobxRiPGy9ZpXc73Ag
hBXihVcelKDI/aVzA6ZLanbQvQx5A9B+zG3Q+Ivn6M+PovUHRVsV2DGW06sOWsNL
pCenUL3aOtclibG0B+j2xMfGYJB9bIiiGjY8rKUUqQrfN8UJL7Gc4qZbEU7Z3MfW
WSlLOBU5Ii0pUA+n44d7/lmR4jbVRMM4UzGJDbP3CMCBV47sTp82Gdre6nsVnn6X
PJ9r30R58Ly2gc7ZlBCiGhn/01OJ+dcAm3dRwGG0RgYOSIWoorg/fZMSZsRb4+GU
EecneAUze6dkBSieYrfpxGfeqMr2Z9bt0726SxRAOik8e13cgqI5WjyFcmFTxNGu
UsGAh1K6Wl55WHCuNdHeTLr7o+H5VMj+4t5PSTygYZEu9Cred8p9l4ieeE+ivR7c
/JB+ctFj35gZeLznF0sZD7FtbqX24tiwgunDcVE6ip0EmQiZgZNALtm0vbB83mDp
vyD2jTZDiM8a9bsSUOPcj1MqfmP7k77hsTM9rvWhwUj9IKGKfXdES//in36ZGlUp
4OwQTwbPO84pWWho/RtitGozSZ+wxi5zXRw2G2o9OE9C6AWmw5MK2PURtKZHLZJG
PwHpIHryJiGJxK+u9G0QU53j4rnOPgAyw/pr6fOTEB2xPfBKPJnb4A/++fQR1hf0
umMvXjOfkIffMFI0yVDOJ8IpywiMMmEmuRFDc11Ckq3uLKVHE1lNBRJKXK1eCpAK
37FI+E3ObjtzchMZn9se/44wFIwIqszPlqPuKUZKeZNpSBMT5z0ABjA3l/4BW4Xx
wm1Hz9JbUpuhZJQWJ+BG0BExUqqq4MUV5WR2U/VSJ6HLuMkzN1bkYFdRQufPWnI1
rEqaUaCbUGcK3fC2tpKIaYw9M8dSi1CjZsTApVLWiI0S6u2hjGn6pDv1pyo/HJEK
hPfMGtiGjbgpSOBHcI0PDyGWe5VekElz8XdHekW/a86pVnfXIItDcxo+9pHrF/o5
ZKkmp192T4rA3AmPOuLZPtGZAyq/EUkprtpSn9H+STKKYucxF+pqKTGQy0KvdvZ1
chfO0d424n/Z3ceNzgxKCU9oyuik+xQIwVA+e2b0XBGgbcQkJmYf6etiEn+UbBsn
Nx1h+2h91NF7u/URxE822ltV+t5BT5KhySE7KNVs8QPUEdPfs89myQdVSCg0UXD5
RsbqqeBm+7FcMVYrq9MsiST7gbbFNaNMxJfZDaJ8jupUYakPKhCqw83aPsbiUVJg
mxzfp8T5n85F8B0cFAgICGSdaTfSZSlz56KFBUBGWTRAQHeK0DqGcrI9vmFkVZ9d
V5tFNjVySiu9pbYNTLTVOvyX0YgO17P8RRtPpWphKUCthmv8T5k++xSpETUFzcP+
nKZC5rom6/F36oQpRnftfxRNtJ2inXU4ZlfzofvxmlPyAoiIsw37hAwqZDmHFLOD
/Acmh1NSQi+b67ystoGV3kmvoZfuJg6msMRxwn0iPpbQ9n8XmCd2ZIoqr2h/JVbk
dV/wkb8Sk5RliWaajsmhRYwYxcpr6pY+wCsbgea5fmWtR4UxPrKr5uwTf80rvdqX
N2TJiO3C/Nz6241VohBzDExS6V9jZqHuQgrbNJS6Hr4wEQIHDDRTIKw6DNzuoANX
Ro7E6su4pBv/GIN78q51nHn6fEQK+4qGHAiMvknXhPCUyjKDuhEfIxjrbf9i+gwG
MFZoyMH1g1oaMCzZNUTHEIw95ycSr8WiDiHDNH60+r2C1LjerQNS+FL1/Ol4TMUh
lkPW7IoZ8621C9lVLhz7YFpbpvIRr0yyWWpvEgQs0wFJvuviTUvKf0DIrQUt7Ufw
wrYfxgCo38qW2ZsSoJbtBXVfgtvntOS87Xja8Jdv2T9sfZHQSBqdGvO4dTWCyo9U
J7llUIQM8o1Kq1442OuLchzenWRosWEOoszm9WouPQbvXt5u94lSZuy/sKXxTaAh
Xa22hoir4FBS5mDUihUjos2v7M5yuNT2hXHjCxRhCCFuTsxvGkEufvgiopNVIuSk
66HnGUXGQd+bF43BYDv3tefKQ43kNrNTY5rspnQHPdPbd+QCW8k8jZFC3zIuWoJk
DJQY50Po4uzHcoyx82l9QC63LaMWjU0+RSttCcJYUh9227F5wjkE0wagI7yBKBSQ
B2iJ5y7ZM9kALC8JI9bL5ozlC0k1xVvOPgMetMsbApRce5A36qnPFfUDVv6/bfbp
YHW2P/Dxgi0dmKUUFQKt2Iw0msjVz4eaXCkqmq/4MCD84smYc1VSXBdvUKhJyqph
67hFgZDHrCBpjsunz8WxqFU1KNMJhktDWKqyBdDhJx+s6vIS1oMOXpmC2YJXrO/n
fcIl9zT++0+zodm1gvAyPJD20B7JeQ6sCtO20I2f1nDtrY9r3L4K8WzG9mklSdeI
XxILuB1ecZUUEZHAvAOzUaJtF1uxY+wTHTXzFSuejU09xpK111iR14l2eKB2+9RH
4HKmi/tjNOp9BCv6k/29s44WW06a/WcKNY0OPRdUQ59fN5S9GEOEB7C9y4maIbSw
aoxeSATv2lwIMokfytjAQfA2OIA8fdKaJkdy7EZJ4WiULg7zRkYitvv/rtxgAZxk
QdyzmbvhVfDVuhLPDuQEwvmSzM94ZMXYNAmgq5OPFu0u+y3yubf4U0eGHZLImbuC
QmJDl4/j0ryxgwBNtFqL8jXByqRMkwHciXzZf5A3t+pszAOTbVI9A1a51qtOYtTS
bBA1iBFbKmTLP6nl3tCYqQC34VP9nVvZo7kyf8+zNjvq5QbvYs75VOpTAtePjjHe
K9+Zlht3Myy0NEEZnGQ5Mc1YZExla+nKpb+8ZfnHSmv2zGdleIBSqYdj7pMd8Ig5
nS1A3CWE0/78mRscC9rPbF0PZmC+Mdfrqrwac5bScgRjZWbYWEDsBNOVx//LCBs4
0p/1pNXujkcg0l+IBGUJzB41k8M4MyNyN5sr47o4pRl1poj5QW2YGpNQOOsTiutS
PlCJOiz5cktHM7ORCG+LNtJxs8lMExu/mnOCYjDFvpcpJ3HYcrpI91h9a2mozj4O
Z6SMfin0upwCKIHoRS1ceJISdh2cimEXgnoEbzD9P20aFvOAoRue6SodFsdcoA0v
QEhiPBQZM9HcneMm3PdH7O/jB0/PPafq1qZxzvlFYG74x5MCr6H9Rzp2Ok1sptwD
t5YADHyWfAyoC+IMqmlK73eodrmyNZbxHWVwX/ZWgxsyVIjqLtbo82yh1FjZE1DY
Qn7QRjHTDsiFyixggXvYmnHMXRHLjiPsgqyOXoo6J0SywRodSFTZo54264N8LBiN
DPNucUQO+XH8HrkUSXYAA6Tnpu1j8GqY4fW4jRKDP6k7YUqdujeYvWt8A8A1vlc8
Ai5tYPRIRAppPM9ea7HFcObvKgpaCz1pZ5c/zxP9fH4MxmwTX/yj0mGeeGthNdPg
/Im/70a5mzIELLDkTkU59eA5fwDCH8xFMXt8V/UXT6eB80xFK0E4hqLGtn5hIKkR
un38L0TuctLxewAXd0Nz8fdhihiG1/MwIUfjwLcD85CfVanb+6ZF5fv+PKr/TZnv
/NmRBdlxTpezXlVawsP6IdIeAJTzbWOz3GY2FFZCMzNH7pPCxm0ODb23Pkux1SBA
q4IaRfCliofgCK9Pwdyx3vty/hJx7m/w7+O9G65VxQfweRP+a591c4Cpx+27Ztx9
HOpBPdrvCQoS6SdEPBiIia4WagqYKeTpWw8ICcz20ocAuwtCxF8PuKaW6SgqRypK
vOspwHf5lgaukPGbnuE+7IogP1d2X6tVinT0o2vDLgBX7UkilI5zs8r+9bLdQSal
KWmVqcHR/xVrOd5SvzVx64y9JRZbQMz1wfD4La2jwS8QYVCh2+mDlgOEY8KGBTF9
D2vo7QLJnpT+y2Icc6KmjiRN5ezehOBVcnDXh43x0zfGp/sV9cksDtNa03gAdxeP
9WANQ0QKUMjzUAM9LemrXpi0vfHlcMni9XMgyHvxMi4b7TRZiuI7RfUZBL4vt8TO
yyUXn+fvKfckGQ2dLymQkjS8WuYeQaKdtOqNtmL9vDpZDtMYgTmq4Yc0T6lBHOUP
BnnI0aA9qafobQ3ho0J4DLTqJTAvlz5vDqUao7Y81njhqfg4bWayld/L/IIh7qkw
Kju9qmpsZBY9S5Mw5QwruhFeSSUDlob/+gT28Ovt3Ed7Thjt1Et6Otw+GAyBTjUh
zzhlk9dpbrnZU2CN3CdSTaGw/B2lc2sRJYcFDAN9aORv+8nNXc9NY6y0wKhlCVsc
bPrCiJffBX1VMNy+/AbCZPVSXHl/PoR8ua8uixbGW17kN73j3jh7n+TUG00tdYo4
e1Yd4cTKEUDFZ6fWN7TumWjd2hCImCzOaa2e1SG48PH18bnV5gbHuyTem//+pGG6
GjdUKzKWUvZL5oQ/8CHi4j/FG7pSt5g+L3uB6YmUIEmarys1rh7j4Z+nacK3MxHJ
QWLW0J4eOFiNeKeR4xX5Vd+VWYUb4OPVC4I+GuqcHPrvf8JzfcUfWXY+/RaD35e3
n4m3+wOWL/5jyZKeuj4zUyaa1yiwXWta3a5hdYcEi/UXxafU3JklFe4t5gPD1ETP
QjdNqzaOhIvJXOJbAovtgyJun62XdkGYfFbHXXhQkkWpmfKZejJ6Gic+2TXozoWR
lTSHQdY6QeuVgssYmrCZE0CucQ65rXdpkXb9V/Tyg9MSbrPW3kUS5CoSJnNAFSjU
QjjYqeHHsftOdeiTeQmMbhNwr1S6J4tdSd094KVhyAtUUyfu5SVBuGumpOay/2/u
nJi4QJphDzTSQdqOlZ++7TLhyqt4visWvidQ2braY324qsWK8fSG1Yi5XoNddrRm
GHMlJgeoUPYzz6GttCgwHwUD6emKrzw3+orE+g3dTzjrFkiU3r84wApglkWGcrpD
DwSFgzD0nSzUEtQyJqAwLceHFaOi4KbM6+jJZI61CBP9x2y4Q6NIdtaNazTSJCfC
Wsj/lE/xH2CG7XiXfiJq+NrZSazyRADTb8niPMY6AyLATfuZrWITXLEYkmPjNeWX
dao5yA6uf/NQVZ0jvnEsHxQHozdaFWKZW1hA0vLOC6wW1x1ShJjOlxwm4K1lKVgg
RRe+MVuRP1OcW6AkFoG4qcAexOgY5lXC3e0eUZFz4Ru+6/FKhPvN2iA/i0SVmKCy
5Na7lX2O9/AmF4DjPrn9lmXPLnE1PHJuqhAj8Mx0x2/XzP5TI9l53Z5dYDM+1bKg
0SB9tStPp3v3dju0S1cjZgAVhIa78SfsSRB5GaKH8SR/KNgMgkefWKVD79YlHcku
5+C3KGwhLqO/PABzUURTC+YNEMXuL8A0RARpmPVCqGEwM0Q8ujZtCHh8G80sle8s
R3Qf2sMYXgJ9oBjhCgInte8M1h1NzeACkuf83ZcPCKkE0n99CJy7jvZ0LoSdop33
oHtBpq9P+XB/9+jWKuQYRfMsgynaX58I6T0ye4QPkOZGfw4weAEqE0/+MAmZJZUQ
6ZsAo3NMU3BRttH1o8wDUmY6GglVRrA23wbCx3UKOrjB8WWIiAs9oU5Rg/OB+IRh
nHowzqQNOLIpyCkguvHUrNS2A9aZbSc21P/B7ExLTBIAMOvG2C7Uv5PAPCUAcEeN
ckvotJ0dEpJDLC+kP16RbU0zE8zOO/ToGYptthq01IhTKqqxGFLjzCHRZzyj+51l
3I71PDd8OiFlQr/6cW33/SiKLhvQPvMH3KJuYbkvUnNXjDhyhn4YWShTWFucM9w9
8/mlH9ua4kdVTIvlZEBgF5riBE/KnNUwhTGTp+weHS5oL2nQBhTDylR3+LgRiu3T
8JNSsSFmhvBIyppAbbwbPwi7q2IxnETjCsvVbVZQeNj7DZQFnrbF5zYpyH9HkX5X
b1uvWbTeegrYQmLQw8vHpT1c0wBIfzQfV/qkOYTtyTagXgy1u6BoRz1t/Qt5Byw2
QDk+KzsKKq6jSDSooPEeLqGDhS5f8YInB2p/2muA2BT2KOgdyQB98pQD/jyOZQ0b
enlSUNhtaOhga5rW4pvq1Ca+ishwGewI0WtFlrwbFiMkESA8CbK9/YiuWJjE1Trf
U/Jm1+RMUqy8XjTWzUxRuS7LUNB6lW2UwLOCWU071e8Qu360cdqxDa0x6WhXe59s
874IMMKlINlDESlCGMm0E+HSL/Xjq7IcX+IEMjvZxJB1ke+Nhny5IkumZrdxxXOp
rD65S+gg04YcrfzydmRLvYx2RkaVL6a0baBtDbhz8CWmA1/WOMUdKBcw6LOoiMgy
OlYb3dQkIbpAW3OZZO74VmxnS1eAa1D3SWH/xeNUR0owRLJgv047jrW636wAT19Z
CVnOPudkQ80L1vBKYSjPTfQyfKl/LzfNJuRHjdioiVo7yuNMk5OWtqhfl39M7ce6
Yvvo+q3XFnbI3t3v9ajbD4U3GuPhJ/sF/6LJqBiQr+CvmGiVuhtvO7Yv35rscrQf
yFagbwB5HqXMA/iKSAhVII31Zclsrrr+8Fvs6UGb+8wpMlmXMr2ac0UJ0v0I0TEP
HapPgxgKvxiIPgRrnncYzwPkLR2sA6aQtXux+fODODMOaEYC4QL89Xh8PZRvOtEf
S/zmWXc9J1+ksv+Tu0qcn23iD2NMhdusr2DlehSl1EtfHak8CadRfAQnoIyRrWC2
wQJwAeNgwhQs4HtoDdl24Q04AZH3ZvZDgJgeDmLuAX78GU0pTOYB+fgtHFCmEWra
uK4RqpCzfCz0R8tsWLN90HSibjv5E7Dru5whNP0kaW++dX92lsuyDXRCrAT/SKTs
z4KA2pgPeDpKc3Khi4RGuuuX4VWNopS3pWDBDvrduspJIO2f0qOEJFX+66jtIhBw
XOSHWWj+pcvE2gVKUpvHpJugftH3ikBE33lnQFO+zaPspGwV9O3F/72j2vepavin
46of9CMxdjsRTIGTvgQXXHAMZcWcUIis2bqA7lMDTdbIrjmLUczbTmR4ONKbtPJZ
o0CkaJJg/9+D/SoQClrGx4q6eAJKpC1l3Es0xYeh6v0zLMHNJZSwbxarO3463Reg
5Wg6yFVPoqD5Ti++fiaAN6LbTr/lTFNO524G0al4VnJ5TrM+k6GxgfnuTVIlqxnY
tP4tx7JJGTKtR3/UnD+Ya96vYSscMeh3GN/fes55uiir08csbqFnYki/JlC/fgkZ
qvYYvpcYgGRQ9N5BYT+0m69SYoTXaU7GN7yMsw8fYVu8SIfvT1UCeBu9YMbS2QWp
GAreuSrR9ltvnwr7kI5usDJa9XP12b50HV9WDzTIoyjbMKAIawSBZZST5UOCtd5F
8RmB5MhnHH4PiIQrQZ6jxlix7xFPtjYhDxM5jOIFQ+CKKcMw6YOuj/Lb38yOc6GZ
MgddafuP2I5U3TxEaulKQzZ4K/JqYhKZBbHP6Y2jYU940ePhgcpBy0werbqjwr2M
Vsmpmi0ZNkjxc6ubZjBB4K2Im53fhT7jJUOIUpKGlQvw3xrGz4dHEs2i2TG+1rjO
ntPuxWaO0WLD1PLFgd5tkBopoKZGTkERSze0FEEFtCiYtLOyKbvzqIFN6SXalp4c
3v2ayV4v+oH5D8WGvkHIgNJWh++PY41HrbtiL+JJ6JCxr3d4x2zQq+yDuG1kqWdV
AmI0KmLM1fJ7pF9yxBsmFkpYefmGUCNr2FHb/VPHtmHlK1BstLCEDzWAUhhacQzs
HYcRlZ+uz/6jdMVkxyqBY3kpEFVQJl8qYCF1+0ZW8ommShTlS5s6DRImtB3ZXphI
xJBhorZyZK0ZKtWbBpux5mc8jhG0WQIunzDjIY8XmmKeReQA+hpeF6tVf7AufeKO
R8cfu2MHXSXMoqI6sht8GnxVVgnzbOxCHXxNw32OWFieWxn/r/EsxY/JcibslNgG
c7aBnd3Fb61gkFe1r8M2/jDmNbAQaXcIGeEDo5of2u701A2sRIBTxqe29ru1FSDO
IpbOtvayWXr6KYW0sJEV/P9xiX/TVQWKNX1a9azdaE5rHgncwpD+vgnhpVHMsSFI
XbbmfM3Ave91G3tDLgXUQIV4DEJTTB9iwfdMMGXONvrSXmfGSvMdl/h3bA+eOU5O
CxX82VrTsszeOVkr9ZFe/lhSFvWW7Fmm0L29JFCGl6bG/upyn9C+gKaz/7Y3EjTo
bL4JCRQGbDz7EXVsskU1X6ACY26fqIrcQYxu0hQQLt/jNvZXIc1co3DWFvbGJJeR
A9qQXA4lKkvLDcVVe+40JWr7oWWwW5NOG0+Nt50moVp8B9cenwjEDJfdZnPUcd5h
BBzxzTA9cj1X3mkwIyb5dJ7wwummbfdCv7OemY9WmmPBYiMXKQbxx8rkNfpEJKCj
2COBmocpH/TReQpxaNWNLm/zBdFtRnJf/Lxrjmm5HSkHfY51DtkUhS5PlDquv4yM
u0TWnkSXj0HtRrMth5n9d0t8HsZoggQtN+lpyhsf15XKLxpBrY221ThGlQonYGve
fPV/wAQ16sdF1inWyXSXqpRup3sARgK9FLpj4UowIJzFvcyYm/g2jM7Elw+IrGP8
xryJLecXqe4QRSYOfO1E8P6XuYylvm/tmLbmvqmf+cCXxoTbvwVJPhP6J9sdkPBx
b0ciO9NN1i0BhJSOgEqDKKmSFaXEGs6LnEAtizAEUzlL56MCFMHZtxN/DaG6nBbl
AeME+42uaqbv+xfiFwozeb5yCzrSFJAm7xzQSBl8rk6sOj6QYiSrhD20kl01s/jT
mSnJgKZCF2x/+f7hg53nSvRuTsu1OPleNTFHWG0B3g5fj7Omhmc6G3mkAt26bUaV
owpquzjZkv4968cQp7hSsBGJ7W9BjXr/KGtQIxqAiPijJlT8FZE2IzqhHIDQC7cR
Zz/nYPL9f2HbQFBWtAb6xKEA+hf8A5bjyhYkQHPaR7IsErdyJv0VIyXERxUPCTk+
9Py1z7SywxFX4xV8qr62WWPGIyV3k/YQuCkyX/uH0zaxr3lf2TFIfy91v0Q2EEXs
7x0QPxPUIOiymZGmQE1gBLgVDTfdRSjXJ372yTRMqEuIIC5Ofk0F/5tNoWCg3JUi
RRy/K3p95hu2wbrfP68FSP7cIgRNHfDLC/c6qvdiPtU0dSakABqPy01IyuBf1Vsn
0OaM4Dv28m8I96rOeOKZzkvAPkt15cb5JlvG1tVpga1x5hHTPjfv/hsMth6wgeZh
vuh9Cq/sfKkS9BLbCxiEIVT715sGceBZ5YGTl/UvS5u71mpiOUWokOEdW1FGyhnw
s0EaA3aBcj+hruc85XBKKbCNi9xUMOy00zvFjo+LwxvhmJ5DNMezzcKHta3eKYfQ
QA7EjmoWBF/PHJ2qN4mp2eQb82b8p5S3WrQLuZxZ4BSwqcXn5tbMGSm9cqfXmAaY
ZT5chcqdZy2mZ1RZ+t19MVcJZbxHoI80s4qC0jEmlJJiQC/2N+kBa5ivQ/ddnpbI
BhotmQ9naOOoJa7s0o8nKSy45EU6AdahQsA62CxSwXH5scCmhPh2ek7h6vl0nWvg
X1P2aY3qBy49RjNY35H+jV6X7ISXg6okvS6o7HroKtXT4cjTU9GNHlvqenUp7na+
vfY4SimX7ix3H/3p7Zsr/CELvzfbxw9vvWjMcNWfgBsEZqYFW/pFhbislYnYqATf
BEQiCT0APP2GlM6y3RIVYJ2VLpUFmN7B8HgSn/Ii0Oj6ORRODuWnbiH0/MqJ9GhD
3AVtROX1LJSsUy7jnExyKRBSZkPdtLsRk7nQr12r9zyguxjoM5nj5Sfi5fWG/3wu
c6loI5Od3r0x34QGHL2jaFHZX2EJ5kGbaMfqN2hLNq3NRnd0zfrjoNikR/nGDctr
OUjb8Wt5PJX/UUEHYYYwwmW0wefthyK9E54hPSVkcyW9eruIRqw6QVsxjaO544+3
tbX8aLq/hJARQ6vHUQhTwc2KpeY1K4Wvdzqt6sr4f9w3fpGisqqOSZNIeWRPoBsD
zOG9IZ3SgTE8tEN2ZaKg0Bjri/VFagylYZ9mTwo+0FlDTQ3Fhr1UbFWNqMbwo1o/
seMeIysBU0lLKhMLicGFxAWfB9XKJjzrigYcDOVIC5y8AEA9iDgK33ewR26PNW0F
uyjI5xX/wFVvWJj/Phv7IBggtqymd1rYMYSTYCTE40eHRRy9uZUtJlqmDZzCzp1S
7vKrd3l3cwMZpr6ktkxBzE0JrxLOHW9JwIOLMu3nzUs/FoU3IAlhiM+1nW+rcR8K
KL0zmVS8q2GAXo3/MG7p7N9P0OtiXqUZ0x/J2Qle3Na/kx9gaDy1xxgZVc+Gb4D9
FiOFH6vk3jB4OJmosJh4u6RVEn2BIAUw5bsI1/qok9MUNbE6ww4r+eUHm/TcIuDf
77yAkBIhkXV5D99/5QBq6BKM/dSMNRSW+Ma+2SG3ngRO7AWPX7nqjKyCH9qGbooY
Aa97qgRxjgKEibeS5t67BpTz2GoDBsA/mT/uBxrZbP8vdatRYiFkuB9nWr9IYdJX
iS1nryVDi5mjUY5KjIoRZZ77ujzWDMPO3Per7M3hG9o/YMC7wGK+JgKMYQmKs7lH
DkMHdS4NLTlDQpcpzite9h2SDfsyP7Xqs5wDArjaxxnbkq0GmUtXV0fV+e4LhV7M
K7dqfuMiVnEEk1n1Jzv49qqRKOKMWq0TsC2owH0Si0W7E7DRsEOsrmIXw4+Zfsas
EztciVBSfT6d7fQ550QZcLuiqzpjPpa8qR7KTGPKTUaQP8XsVVvqKe0+PBO2ce0e
AStyehOS0/NQpYObPbuQj1RmB35e4bCyxZANNDmv0UciSzo0PeLpL/i7vY+dMCFt
+0brOt/mZiGQJSkP0+uV/cnXtL+z4ei0tze9Tr4vlOBsDG1zC5cO5pRjOXHeONot
RXThwa/g4TnBlbWoJSngaZvrb0f4Dxhty8grNvLvVBot0tTXxZPVo2nAwdaL395/
Dm/6/bu4juoKVzHMOBSuD8jbZyexoZnl6qmxaAuekSkxqmuG62MzxEUOZZBzZJji
hk57SDzzs2xM7qoqOGzXtNGEGVp5//GAgwKPdsDrVjBBMqWwUIKQYnpUKMr0zsuy
ExhXoH/K7nHIXRTXv8CamhKKwc6/Cyq2VW/dIs+n5JH6sg9ZSuV+9OMNgADYyB5g
0KVv1fGNgfuXmsyMqAtLdun+mgcFi3cUgckwxpxrvwWBlsSaMxX4xXSylBQbK5yY
smdrDds6ICaa7+nCFCY26AyRxsCGs7sUWXOlpxuXyLgT/GSgsME9b7psSPExvpjG
RiZLV2cJXSiKRWy1/t4fg00SFvhl/5NRZk6y6cJR+SQnO6PkoQQUjaMnplRXLnUn
Gnl3uya0z4S9bTZVxcpVCiuzn5pxME3KUuvKvWzPFozDB5/o5UahAn4BUR+ZTzRE
GtkjgaLS3sQB7BI5pZbhCPShtYSq5ufLxfTlNaHR8bFeDv9X/LRt2PqSr/iWBdp4
Ii7c/Iq+QSNXdV9oL0vE52Tc8vGyPl2UoDIH1OAR655Soq49Jp1SRNfh5w6JmZQh
PPeJPUF19D1RBdisgT390S6AlgWgJCybHnRLxH/C4i+bHGppucHs1A2HCN2whBXk
TLA7p9IEZVfSfGidPE772VNf7okYcY3ExH85y7A+Mw+hqsMN6iNd0UrrLMtguWwM
IcEEI85AF236JsIaVkIKpDU1mc+bL8rnNzHm13JnwSunSZK53UMU1p4Viy7vcUGW
gILwMla5ZJuqt4n4MqDugLPfiYARrZy2xsTHxRGGrO+s5U/kB4o51R+5rzh2TSkl
+lc3HvwOWj76WiwL6LJ/E5Br+tWHmBUO3vq+p+Jecqw16C80XlqWnPorMnid0ul6
0HCi7r/tfITZ5ZdCZG/2P9LB5BRoCOAYEBqEexSb2rERVJW4eWrPhLK++73ZgAm9
JrUrLgnFu4gJpI9FXkjJzp8xoeQ5A30UZBXens0BJD8NLzh9qhVGp4N+wfOsXYAb
SEWeSAnqfNs55emLgD0FvFufMnN3Xylr65XgPg76VtdJjedKLc3dHEfh/+MwaAFm
zSo4Pt9H02gvR+jhVNwNEYelgb7xi96QJwP/H3vA51UOFLmG1LebHkhoK5IjAxEo
vSCI0JETN64o0JuyfG6TwRM32TBkcQmDfjZisA1ri8KEgC4dxBGhsM3m0yn9iIZc
HfZC3EFs1IMp25LosVQDgYWN4NsUQJRuIvtNNMrfXUfKBk79cX45Wx4g4l5WU3RQ
ZIvw8sILrOEw8xUyBACa8qVekJFOwcLtDh+rU8q0pcZHyuIkEcPuTbYg0uQCgKFv
J8dLAX7iCYApGUKp/AHgs1t6jTrf0dkfAESvMQJels82++wtMBJ/0R8GdCdMlE+i
vyV08wxys/1zWt1O4WVCckN/oMQcbS9RfuH860kETHpVbJPnJR3QKF+o5syxA3pH
dCmdveSztm4IyBUrXDQH5k+LWu/SKkz+j3wM6p4M7zscQ7AbvFtJ+UEWWuXPcXMC
+/NkTjpQmxYqNSyQWF4Q3QPh8hGk7f9MQojj5mdxuRl28Xo0S1592DE6KVSOMQUF
bmjZQ5tT5hoRKBvWUJw+lbE3EBhBW9UPnKEy1qWRgCEKvM3Uq1Kxmq5KPrUfGTSr
9e4x83nRmLttZKzgYx3SKbEISFZBe2E64JuGTAYsiOR1wUEWsFCk3e4Re9ix0MMJ
uoNcDvzMqhDZGpgFFLaI65dV1whGjSi0LX+5rRc76wOEdVYWMs4q+q9aBCdhrlNR
sLXH+lc873nDkLUDvtmSIssfzqCdeLl9WMSLb90uR27ZTKTGAiO6nDbUEwuWP9jj
M2XknYkpCI4Kywj82VGUTuSdk7TQXOjRQyned/dnELp2ESOol6REL3TH6dj7JYyT
lzWknhkQXmBAJQdRtYbqOIUB243Qh/eTHHArW1CZj50ffw+uDhOcmN/KvfHd1BmO
J0t8gxmv7lerftHXsUOG/PZvlKghCRNSU/A2A+AUa6jtiTuBw3mMtspIYpDkCIRh
ABJHxBcWIBk2fS05AEVIUzKFFNHnS1wtOiOekJYajH1NhM0RnXPcYWDpdWRK2kri
huJx6d5+vCl5wDpcwKJNLRYUHvXeEhIoCMUBj2qv7c0KdqdH6+PMTt3PF0UV/nNk
bZ0XksJijqf+jLwNhxdiqfaxdqaxMRPdPw1CuXmTdxRPCrQzQC5LdH1sRrUkKdCk
yeakt0JvyM7EAWF39PvP1EPRLkbBhoRCMVCHNbY79L9oo7BV92EdpPPFGa8Qy+WB
thXUjuf1WYkrPLq1IemHWWnNREDxpNcAfXGkQXbcIAnAkKnDuCDS9gKHNGIQnTtY
t/MIYjUU46VLeGGfWYcd19AnO0iEzOy9HcMieyHf9z1SyhN1AkLdnt9I5fwo3846
d/LPs5L/Z2r6GlhJYEP/optRQQv+v2Dqai7tqIxP08hb1zFuQm2gocAUR8T2Gzww
NLMu8Fs918Zo25wi3SnDOGh6tMebGe7sjaPj7+l4oOXQu175Z05BT0CmnaE3noBz
mU2SgxH4ibqYlqzkmIc7v77oGR4x/0wJXD7Fjh2JUjv8lahRMBbvWqrS9QKzgC7c
2z5luUdcFymnNs9+xLoOtT7BY0vQ6PEaACppUEdLXGd6MBqwKrTJ7iVfQI/PX8kD
3CyBYEPTS1Qr4hKyUsw1IKxB3ead9Uew0/dmpdg5ymT+9aXfJ6JdpuE2nYkbp1QV
oyWHU/A+8AhCr/OXZW/8n3Ezr6e0+2UzD9rld3+5dfvWoF21iansoFsVB6H5xnAV
0s37nF2V2dgESlsKzR7ushRNGgeDQwn/jH+acA2YY7zkVngMPH7f5q4uUSkNW+Uf
LW0ywQfh1hemzf3qJ7fR8L3hnX6jdlO1IQ+Xs+l6M30ux6uL+MHMVVCLzVnrxEvV
bSMK++2cPsOrq4O5zRlgFkJiyAJWkglAmnsBj9D0wMEt37dotfKU3H2Nt02lxv5+
Y1KwILVVFFoEPa1M4ZFBj2yMxGtsQpyYzhopKJWg3onlwvw5P8AFrQAlaC6fw0j+
uDDoU4YOyY1FR/fZsC9rjvwKaiPtkueQV/LPEoKJrTYB8e6gNmU/Rpj3lxEVxM2m
em/VPqLY6tV+4qEa5mlPDfAQcAc5rvV9a9MbCWO3VVkPQPCdQX5GZK7lU2z0xY4U
yC2aLVAXJua2T3Tf3u4xsLhuwi+bXdCr6MxtNrBqPgWr00pK8ouqcAkSUkM+u0RX
34DO3qPHhSUnMaEVlQtccL8MDHg/du4/GqJdJtDXUWsEDh1gKvVLOdv8qYtWWqVt
4SbT0R6VTmZADPfQTS/grgexby9NlU1Cbz3qYmy7b0E4x/bmu7Lb6uVlaYfSSkD2
wWnNqo3RPmUejG2PNs2hS0DIn31mnBhT9wyOIj/1D8ZVLFb7O/fdzFX98Pm0+Hgd
J1793T5xOBVfFn5uyOBKAmqiSkWyX8fpPxXosROrIoWDigsDHE7T1YTTmHO5Bd4U
FMh9sQDWGAqPSNjaKGqhH3BZNByMdV6WgUXTKmYYx0HTLlp6JNsgWOXktASb6FXo
HFKEqJi0SSYy7RGKwY8zW169+f95qs4MiGtbxIdhjIyUb1jTWcdl8Qtd3LNR5Dkd
Cacnnf4NsOS1BCKyxPrcOqN7x3qmn69PnB9nE1iOxcmHCNZ+0FZ6QNKrxyKl36kH
7NjATEBtI9BBK6ZlXYKfUfhAOPkBNugmvJbD/RDYS43EhE28w9deLkPQCbTvteUv
zbdZEWWBukFqJWB1/uJRryMNOkbU6rwEy/E/2YNp5T4lD9zXY0Fi22arq/Uk+aTo
f0WBgnTSWzEJ/2HFgT42gMuiO2csfXPexW0MmZr+KzGBssPVDiBKmjLruPDjxR3g
cSkmpogEJTAwIXmavi7oXxRspx9zXmb7GsChfx1WyHjD63q/0uzGXMw8eOsksvrU
EQQ5jgD3jXlLZmg444aQtRAIl9+Fbk/jqazoIWY5aAX9z33FaAxcyX3tGkBUpcwJ
f0/U8YiIIZxTJTsquuiBJWxEhKSARXfIoPlPYq43dRs3ceQCKGJJhwYx3RyDdIG9
WN+LfAvrL6IMgDSgbGJ2wyPhF5Hy6Ka/xyKh/pXIwisf4hm3XU8OvPZrzqBWa4Pk
ysC4hnKIOkP6G4ZCVJ/YKFjL4H8AGS9pJM6ZpuJpPFTvJ/Tknuhd44m4fH6qIwqS
AF/Y/DQ3odPusxkVimxHHcCMD5376D7awUhjD0QK/frzrK/EEi4/oUuQcdvJrjAa
JiAAiwFAEHuaytSVkWJRxyETW91IKXYmqWzVv7Und8DoxtGZHhXPnvdZSdyqVWdQ
90lQQYV67IaYwtjUf32inFnJ3PvH6Y1NiD7z1xsvez4HjR/IAWm4o/v4LjrsolcA
QYPALO5HxDe4xuWr1ptwE1fA+3QcEb8VJdIZWA1MCR8n37WgCcljSktEdYudGbog
d4i2TU7VPZK3a7rvTsG/IZzCg+33HAhoCrNCU1PKH+VDLVGdoZv5KAIddR3zJREr
2aP2Xq+Iau7O2uk2YmDSpoCOSbJVHvgqxAqjx3HCP/Ca0C8rBTzw44np9kuj0i1S
pl4armv4xN3yBNkPU8n4MuE4W9z6PvntqP+v3EMoTbOfHKP7PeOLfV8mAYBlv5HU
8H7Pdm9laa8ewRMOtJUEUE7eKkY8KN9eTytjrkrB9mmu2GoRVvZmfTsUpsHREIAi
CLJ+RkqmgYxh5Tsiub8xP8p9oKFIEXu61NR4jF+GD5OSYFHwhUYnueDUeuwESVM+
+OW1bG/nPWkS61BPm/KvcOiklYS7YPBYeG5/28mlAFQhK6TL3jvbLCbnfKqsAReB
kfDzfVaZBROhrH9Etq9m0W0bouR/y/6etfzKCR72AmSk3J0uQC9yuKeezwpXTvVM
4WGAPL0/s8iWVpdY4XbaTekJGnavUEO8x/D8wDLrX1nzxLmGlC+S0v5iFlUULRDq
DjW2PL5J5fP1vekVkgUxI3nMtN/W/goxvff0ysy6i4VUD/RfyR8eYcSRxa/m4DrH
C+xUNsVQisMtxKDjBox1U/OZM04IQfzK+CL2cgxGK0kgY6hqdG25tWhzXieXlUQ/
76yEskA51YMYZ8ovZ4i6ZijSz1qWrtfs3xEvlnoXhUjRedmJrtdEc6kXd/l/pE9P
VLbnpoEYSgM7eOOosO6znntW9VimW3zC8HbAwTq9LFYtl717BU3ScPA3Xz63cXSu
rz/OGv56hYO2aucxQkp1c3S/MVUSHvW/xrsgfJX76Y/i2WhE3BL2AXV8rooI2If0
Ax1G0GfAyzM7UI80h3scJqhg3PSNX9rFnt/K8eHGP/DQQ0+kOsDAdw1kHFi/d9cW
9og/tGKip1g0NLX6QO+Uftkywr8OsJGqQzn4vyg7mDjYpi4tqZ6smJkUaloKp/7f
hnbwq2go8KWy5I/PX7DFi2g4XPiqnU2QVaoFgxGEkuYH2GFZcDnHl+aVduwi7YRt
qTRESGE8HyU4QpPtade0yn2KEgR5gFoZ32caG8lKhdAGsy+/S87QLOhZ2mh3RI+F
vOPy1rlJhzkkfm0/ofkXD0k7hungj79Kozj5hMa3oEgGXNPgNu0vRKw6+rBwRl6C
h1ic0ZBZz3jw0dbrno7EWkD8OH/a/n+SxGBHum8BzHLGRRSdfUDUpcrmvNex4S6n
yKYeNklzHl01hdvGAj3PYrmOTwmkcd/hvR3B37Y6xwfleKnJYEsF1tXI0mgnNQdg
5OAbWImxnftgQReaC7q/XRIUFQBKgH654fCejeXJtcSZEAgUVXqc9CNeGNnfzNd+
zKgSc8zUNjqG9zN7/1wqVzshKGsmFrSOmF01wCooah4r2FzQSHBvwGPTZ3E/CHLe
FTo4eQ1XlfDEYlhGkpPFNJpedNxV3hK8PaV+B1KafV7lAmxx9iP9oREm0V7yrjdD
H4D+xjLSaZsASElAXnzAA6WYHqmpMU9JtGS30F4CCqofkvd6Oun7ZHucwrrjgxRp
R+3JCoBMkGp/qZBgIdne3M5G8mTlpl5Eat/3LSBw5twOE+MR1Txh4YR/F+PLPShq
J/pICKiJ3z2EpHGBRlMrx0a2RuE3MTnJYkK50HY/NIh4KrZAcT9zdI7BZkAhPTkd
h6KYhYdywWJU5JQ8WZxZo9lcYDKhiRBXVbv+oFgJcp6pU4UENysNAmzbw49HgnTK
jpJrgrJd6VVemD2sfzmXad8CxO+KHzEl0Se2L9CxwQP0dMqHCIKieyukcoIB7AVu
vY6s8E84Vqn1cjd2y9PKbHHLHygkqYDIgRY2hfMwSAr38m8xAoWWDwjGylI5INoy
1SPn6DgsDUepc6/o+9NuYNyKlBjz+yoxoGAMaSNzWx9wSw5xDeuIbvy1MrAKmpe6
mDRS1psDCNu6p0k9DcgFPOOGpICziVJALv0pDoro87c68RBtbgqIRnK3VQyo4VLF
7KwCL8Np0G9ib7bqaaekf68SIAot2pCX5mq9w2GmjYxJ9XZ+xbzuscD2p26vmYRj
l+jJVL8niJERUKM5sWq3Z3Oe4JFMoS5KyymnEB4ZGEtuWGJBci8QM8cD8aiESoTP
J66rsODi2PdxWRNfQJ6RJkYMEtkQSuze0l7V5oqmo+AW6TP35Xo98kpnb20k+yvk
ErhK3gItjo02re5F7I5FJGrAitmNJohIqNn9ZfSf84bP/nTvaIdSWqpCBsuVIS8T
41zHByUSvMMfMtxax7+GC8X8SEJqJ6vienwYXDmc3Cc76pRuHBmoj2qUNvUzRZGZ
KqF87DYv9oP4GaOjOcVv6pWMDvX4fozWhO6WiFeVHB/lr5H8AstfHo/7eU1DoFa0
oSNe6kzhXcos+JqRqYcJeeFUfbQhCPsQko6Ii1Dz15R87jpl85Q1NvVLyK2a1t2n
jaUKsylkRwQnCnVf8WN0WkKbwu8CY7J0k1ktP+iaFtizNl+9bn10t9ylyGN3s2k6
hlvrWRUXecfOGaPB6VafhYpsidjwTGmxAy5yDNQOZ/2xWiPOpR7Egbz2USB+3WFh
9wydvfi31z1o23LW2fYR+J1V4UV7xUwMHpVhdCgoU02OwQnIZvSlEcaOkVYhYza8
K8IXbD5Mb4bUNy8yR9w1p+rL7Gz16wPGerj6VzrUSp1iWh73W53nURDFKw5W8gep
LWd/Nbyaru5kq8TWM7l58OqkNakLO1egDgVLm0tv05yv6ZBvLKX+qzV90UdvcELe
aK5BFx5pdWGYUuMouKxbcfn+hmV6nPNtOz7PIF638r4V/toqQSlAtWTrHEIMn4Jz
BHES49tl+ip9IhYoKx2tEU/cOrgauDXwOSluBU/GL2BEaVXiEoy/lgxp9GPmfhu8
TzSgVUsBc4Hkc7MIg7Fugbp0VOCQ3GuQeT9BMeCqmtJXORZvO7062tL9pgqAJaEo
q1FbQOykjep0H5At73X5Vcvb64iye347URSOSc2kgJd2o7jpf4EhimgQI0+Bhp5p
L7L4lk7byHNY5/VMAKQF0bwXeI7WqtBXzPVns80H4ua1A2Yb1x6RnW6oVjotzeL/
2SR/wULqecKtnBPtljs/M1kfxSA7YdZkbgEvE7MtwUvc0ymSO1K0DSf7Aqaavxt1
vUBQdQPQeIxiNFkSEcdHM5ITuwHvtGNg9eDBCQaNFgrA0Hlhvg7CYkxzdGg8HL27
czcXe7ll1KK93riGFz3nhMANwVd3P71D+Y5mUrMzhQeJXxIZJz6vhEwlu0q4TY1G
KEAWq+FNisn3IgkNtdKE6qFpUNj31TkUTWOu++WAk18IgmHVIlOOhXSj8FE0ch3G
a6LEwPIlkTPEYHTzJCnxndgrbPcDZgUlmeCxDl6wKpbZedqAQj+zcfqd2kVszMdz
zHYPCm8k3VE/B3cOFUaCRAKgS7sdSRXru+jM5EHd2r7P9zpTJnvi/ECyWd9z7w2Z
mDqyifpQrcYUIOxFPHsxuojyvWmpXL0RcYdBVpQjbAynMHSHHJvazIF0U8S2qo0S
YF6xJwbMBkspdvLGZ+qsDH+JJ5ZUEok2qDx6COSFKkEkV099ssg07hIMM9WLf/BT
aZaQdcxJf1gdGQPWsH16b7+XJKFGdlEZsxr+ob1RWBPqAe7DMky+702YpJTuslfj
8AP99l3ls3NShplNy5x7L9aXux7Zkryy+GVSF5PLU1cudTeRwztRcLwFF+H/g6/A
mvOwXIiC+byzVfndlZCvnXnwsQE5MVlQv/lW47TF+b/gKsyLj9w6UquC4LxqKax4
lFERdpuPUbTJQiNECpTBisT9MxduKxpMntOSyTi+YoVHfKkjyn0y18n/kYUDqXci
xfCqAhoDBZBcEbZpb9ArGmn870CQCu0RDQARZurfTu0k3OiMfkbqK52O/9nLHFxX
LVOatzgS5J1wOkuLcx3nX+DSbRCKkdiBQ+q0jT7PmFsqpfPgBlXGgFQGk/eKA8CQ
uq7wcZySUi82eZMhwTJqsi2wWGDP3rW2W9tedrbtLupREm/7pNPkQkfG0I8hrCih
vM5DujdMTkS4FhLroETM06sA9Ize18EP70/ubbMbAvWNMcmw6pdPNjv4tQe9oIhV
QELZd/itWJbL9Br3AFF8ErDBeNs+ardpWBfhCSUpJguW8PJrOYuKfVnXou9OsgBo
zmWVY/jfQ89/ycgg3dAX95OnZX6VdJuv68PoH2YVvW6qa6T+VbYierYeNCvOsJ0g
SUEpok9vQI2RiEfIvUXzaOl+eyKpzwc/qiYi72tLYDaxthexPyuII9mNgd8OA+fT
YXH5ghY5+hTvYAD/pm57r0iY+P/BKln7H6sNZF99BSRd3wIXwa3Kwi77XkpauhFq
+PjDBFkm9YszFaVkpxERoptTCd7UkZzYYZyvbNRclem9x9I1nl8ZB1Mre2zhZcVr
S7PEKsgmUF7EFrqC2gnn/iL/9x1OGXC5djY3I5n7FpI+gzZTco3kSjtvNl7Vh8yy
DZ/FYGpRWXNPI55/grSe2A6zbnQpAZC/x9bqNnN3rC+IMRKSgAmklxut2dzk9vVM
AdLMIAFGu/EY/OcynvDVBG7KQmExxGzz19NzDT3BQFgOr/sFUr4b+ekGaIxZn/N0
8r/b66bhxOdMegg5wqLGyhpPynbap3N347be39B8tN/wIGNdZmjpgzTcneXXKNdM
KCQfY2GeGUsnRIC5soxtAw/TY8RcOF87E8StAfU/uEAKC8zU128TsECs16Hvyz10
2ncxxQFfIrp1oerVjGEcZtFvuNJXNWejS0+Hy7P+HecTxioFYYjpPR4w1QRrr64W
Y6reiKlBxeZnyYIaKHmk/NimuW/wK3VIq/SGNOwXUHrGxA5Ygub6gZZ2gtTrY1yk
nAxkZr/Wt06PTk6Ug/0nn2K5IEwnt7CXfeeTfo5cEF6ZU4h6vScV/5uFtdw0U3yJ
G3+9b2QNchSZ5QhJswgXzmKjgLfbY1vyVCIWu6jd6lnjEfiXKW+JIKcUqDMP7DEj
19YGHO41jasgUAmL1EO1behCQAMbxef/fJnyOlpSqYXU7gT6GH5dwZijVAGSqMQX
VHSEyfJM9/3AIhRYWns8mbk/m9eBLCHaLcjmLnb4hyh6IWfdZKtl0S9WzlO6aizC
MEe3s3B/WR7ItimRmI5Li+ZcFFhbtl16mPMhw1vrb1zTd6E55RLswN4JYDeBqMks
500TJZRGme1/plLG+VOFs8NP3YklRNTsyPhJ9shJNkj2tpF/iSyAL9H2oUzN/QPV
ilrhy0hsRenbxxwkJ/QNCH1d7QN8sCdbzOSaAX/ytyAyNLt0Uz75j3QXtoymfwwE
3UdqDI0slW7N4KeNnQm0lqBpG3d3kS2bNvhSHaCumOmFisUX2fpsEf+3Dph14I06
TgCVplOn7RVlS7PvBaUnJei5P8FFeuaq3KjLGMNT43H0GuasLUmhWBI5zb02YMh6
HG6EuUyWTF/zrbIuhg6OhCVdIbszgXO1dSKa1ExKDhpvpjXoxTDFpQr75OdX/hLD
xHAIdXkGkZ1Mr5v4aCP7qp1AjG2rDv6qURAmikEl8aviZ6N5ZQK9w/q4c6CnNAA+
dPiIvMKXIpwkZ3uuhlJu1LSfBWcv3JuRj9zFcR9Ffs7aPs2WqD8gSnyFYjgJQShs
95aaYlzp9Di3F/XtTHK4+sBh530XG3QY91QYuRUbQk4S9Fnd+9Z/OPrLfNkVPnxK
KVWtqJ737m36nNZH2SG04grje7+rzOClSq/U9wxdYIlahARxmSX6tbD0yE/dM3iR
+OIB/qikoMLw+oTGp/AnOabvKriC1FgC7Q4HmZ6JWG9UqM1CjdixgL7UVdkSFaST
jSbrbgKGfa7hsxLeizrZlOZP99LMZKknSR5rf4EcNugx6XL6LFa3pTPalw78Zyh2
+nGTwY/KKEAOyzdJO+ZMs2FzAvBUU0bzCpon7eq+H7ZM5b8Nd9y+GlE0PGAEMO8y
Y34NYWBjz8/Z+Dc8UTK9GRgT/67NEtjjt+vRhszdVnon1G+2eu3t0K83dMfffUKL
/ZmvEhapkwrW2/GlyJME5VScxtcNSLJb/VgWILJMZeF6qGqoh6KvspQvxcVNZLSh
XIayUw43zFUQSTsuvgOcEgBuuUMZjhV5b+bOM50ZTjnP+4U0dsRXSEGt/hoQrwlP
lMaKeyEUlOzWy3waXCtPPIPob9KRU0Xcn7pmz7AJl8K/Xl6X6IDA/4TgjfVjV85N
AVLFA7p3OdIRV6aF9REORcR+Q3pYcuYvC0DYpXOZIgVl6a5diCICB/OWd/i22ZQ8
FZNGaP5FanhfBbXmxdb5n2R9TeqG9RDjMQh0cv/mHP0k0aQFIlHk1Ihz8OcycjXa
riyxh3hhXyF4CrEYHQobMm1S5z6JI59OnytvUQcXOO2W9U5pTy8uKHSiCQ1Tn/f8
heUBwCgMjIhXa7BLuPGqm+Kgt4BaWLM83/aHITzD+zC3iudUX02kw41fMuwlP6OR
FX7phRz8EKZY3hVr30vi0A2FAsezTZFTrLL+NY/bUKau2scJpzOf2GdyjfUPqgur
GS2usr67PGpsHUzwjWpjrflz0grEnbXUFfCfJE1ad1FGnW3MUNRrFVJIjJKV8cHv
oSBrUd6pBQq7Bn+7dpAKGXhD7Pk3Ns2TPET3bU6Mm+/8znL1Qm6ebh4hgBiuAyAG
wQYHsLJ+b99FLRZeO7+wglgKAgpNc/XFpfcHPtsrIyu4GlC4MRhZMMVATg1v2jrl
PXFqufMJJxOtiKQ4kxuCb1PuX325YlEiGj+TFZpFX+jlUjZZKKS4oa1IkLkZuoY6
/SQK/jTT8HRwiaiUGCkYpwpLFYyQ35xC8LV4IwFW1WM1ik/YplJbvCjJMGs+Oo8k
0g/TzS41dwGzvaJcYXH+uarg1ebxvtX24jvDHBLlFPEaAGClIgfVcz7iF7ZgzOD9
RyylA6hw63T3XAOYSo7h8GvGyQfVM+GZ2SFcbyI88eYPD16wdnV2gmGIoSRwoOdw
btG5UOh/wsny3H8zpjyCZtiil/FP//4a4jJLf8+GvnaTYOZLlNwaPDomTA70T9P3
ufockxIqNn4cX8G17tVACyA15lIQDX2y/WHZEYO0V3Ex4DA1o2VPMWVy/nQACRvm
KiOnZS6Lz/ru4xIzSkpGN3/imvasQRjPQfbCxyfk92jaell+SNl78vp25Cdryq8t
W1Kd6TVM7eSIbJBecxXFgV05QpisPx4MjlaPX8I50WNX1E4sb4RevNO0qucuqb6v
4M4tcfdU4274cKFEuBq+LxnmQobxWA5+DvnVBI80iwGh2Qxosn0wfW3BMM+ak28U
mnKmBxdhCsu14CGfEnsLtWYNckCcdK2JEFBr995oSlg1sZw5n3sCB30oqMC4jrLw
9O7x5BldIPNHyyOJiyvYlrD6RzSlmG7GHyqBUlqirb0MCk2va1uTB3BjfAFwOrYQ
eweAfiJsI98RV/8EaaD6bpgmU4X4TQRZGcqhqj5XZj34ahXwLwn8C/HhUvq03MgR
weh554bmGh0cjZJEfHMtzEfuVvYMLI9mU0v6v4reWGcf28kuMXKmUb5ORjzL69OF
3xT+7SxKNihY1yp5m+TjK+C9B8g8g5W9bRFxZOuxU0X8vv+/Y78/vLQ4xwayd8SB
ZK2kSefKp4ID6TcL9CuZsF5TUSuMc0kGjK5y3P5eqGT0eJ9zHBg20kg6V792AKpB
MCQzJRPbCNm3k192sadxH4Tkb/xwXg08yMKUMaeFEad5WonTmBB/3LVnqbXu/YyQ
OXqRS8RybCEHwVJDyd9Bs3HHNPC3b6ObFW0JQwiILeFmIDjomtH8GkjSNdGngb+o
4M8gOEWyVcFls+tTLjPsnORFh0vlsgC1Kqv3euPoA8h7XiAwdUwdMwg7/yBnmFFs
lPfZqFHvJ/wz7gS1thZLubrbspIfAPauKUIKPp+rUhop4zdTtsHogTk3nFT8FvZY
d8JI2ACgcjdlbjfFJXLd6+HrIcuVxDLPFueQfi4nMJFp1I57E5mCtHDl37RumhZa
O2uRQX1PyMupwBYcT7dpCd+k/cMuY+5hHMZCBc/VMukVA1zTcWFMzkAkzupiEM9K
Tcfy7DWN4DH6lxdtcvkU9M2Wcnuw44GJYTve7SqUmbwSbEbrvl8CEpzrLwjeBbcJ
1RJ4THkXwPoZZwZMo2pCZ5mQAszd74N+aEqctZcJzJEQDvwsmRj3NKXueBTryye5
jPeZI8wnXZGi0VN/1AFu1E6JodcrRClBAJlUbB0OuYzIA+ChiU+YBdbJ2BZd4FWp
FOL3YUQjQWyZDSuwy+qDYqDJ7jNmr3wPN5/j1KOKOx4b+In7i4w9j4jVJWCg1Y0M
qYe39VQ4nQgPT0TEx1U6qTlDythoNbucMOEO4zGGQYVRbceuLFTgCQGL36ZUhS7A
vv7fL4O7ZYz3r+4TliWaoHWbG1B32omkNiqVHpXWj4BZHYH17ocPRFDaTw+2uTaI
yYCYGVpVCvuaIq1Jj5eZmXwAiDu66+EEieZ0Na8wLH0j4dT0kJXbw37uAI20vh38
lo4aRyUommUGk1VtCmNBucgZAS2pGw+5CLcXJAInqyEYrOQEgTWKomvWUnhPG4Ha
pRHoa4L/Hh3pNV+wO3HjHe6pVHJHkvTgyN05PmnDIoT88uxH8bSPh/Oo31wR+pqg
o2DpZIsju7+NPhDbiHAW496ZQsDBGlu2dBLKJ72sWZHjxbETpdNNxLp2Et6SkurX
YKBRvP+0AbQ0Y35MMzCVzhV8WpbP8BEiEo1RDu3vlTQtKgyUOGXLPkAtpj25m5Ui
5TMdhrOfmxyEI5uUJq6V97S9Ot1xkaOHsKnrFm1pPbBvTi2YLCdDgh+3EkAdOiMd
Qa+2nwBXBBXrO8KskaCuypSnNh3VIYhb8wTg6DMU7mZEzoWOctnzT9kNzUReN6++
P2m1EfDDq0HQNWqloDFFgjZiNrEh3iNrRoMrO/1Qc6MS/ZZMUh49owQlNsRJV1WF
zv4A+UrlOrqnktIxIqwRRYO/tu3up0T183c/WMd1wPACAyhHoMHYZEAHf5qlIhUN
HkR1WdM9y6H9790s60QyM7TG+zTSvNgAT+079FifYuIYp8SFe+XlzmQjzE7wQjIi
m7iIL+7yGPg7SH5ICCEabDqHWV2fWpkmvThC+yax/tjaCrrPy8xFYUosuSRzL/hR
AgUPkUb108A9jnaoKuRIHR4DrsGuBHlLxsmpnvjyYjOGTWQp7Z9q6XEryPCUODOv
bOO2DosWpGpoOBumz6M42MRHS3n72jGjnb9qp65WZB4/CbQCwGy/kbI493isMAgg
gATM48XEL2loaq2eVgPTfIr/c8+DwxnK0cAGeiqzCtFyjTkwj/Pq+RKN7yq9WjC7
/69R6FhweHfsREp3xpJJUA9EE+h2tXJlIt26R4ZCk/eQSa1m9jidXLygSnnBZUKV
hE3Jkjz4H8Ww+GRH79wklRF/c4+X2KoDyBo3+4IHp7dbXpkUrji832pFTJ2DkoDk
UoDpbToT7nFA+9Fc+W74CKbuohmY3R6GSNKFR1bs1ePisK3iqMlYAFbqfUH+/yAA
VhyJgVg6FRdPz9NwqTlFkEOr5t2u4PsorZPJdEshZWBjpFmxD+ZrTqLNcXPYqplf
YAseFEiC/L0mCkmVLdzFSxwGJoALtFuMElMgUDgMEoM3gFx5yFBtcdIjhJ2urh69
QooI0Lah1DC65tT7qnZzTPNwVz7r86yi+JbOxwpgMlj0R0yZqk0DS0CGA1dSWb9Z
f8vY4QYNlXcqjqxhgLpBzQj0Skl9FisCgan5xulIEsLHWoE3T+DfO2SoRwrxCQKn
Cc/lXr/YvoeIeHaRMpFhfCpIPT+ORyUgSQ1FfmY8ZmF0InbmKseXE4+rXIRMzjne
y6vNn1QCFLexoXoXk3j49YMenppqsi1J3Sc7gdEONE56253FYaiafI2Gw8f6eWnv
rZL+ku0G46F2kHEIFH1YGM3J5bnTTTxnm70qVSzY/GnqSkGP2kcfw3g9CsU73Qc/
PgWtnQEqQwVwPXwZ1yR2vYosmhu3UWsYjHqxJQA9D9zwOsBr9LiV+rG4ySVkT0gr
U55gf1rOfnBtoOLsMXtZ9UvpWRHLrrW0rWhUezDNKCHxHlLterXEM8218r6CDWUF
EQufbR/fLUW+5Yq71RWpGelCf/Y3FO78Q47PPICjXarBOvAbW3Df9Psd7XLgOOn4
yRc71lN2XZUSoYH1t2biFNE55HyiKdry3/JtvkBUDNvIqUyPiJ8Hhq/bAoZ9Alvj
XyclOWHQrIrrj+pDfemZ1mTBjaauMBa7tBD6YZDU/JUfmBmMirocAEGo7pX2eQy6
wYhjx2Vdoyut8VzdvQBLM+IuGuu0u2HHG0Lnyid3XFeRP80bv2ch45hI0XLjIf80
M7LZnjb0ci5sYKNnKQAnBpNUACtxRzUEeuIH5nDxIT9VZRc+cZtN0FOdLfANUw1E
BXL4XYQSZWtFJkuHUPrBC02ij6OZi4ili3XLejq7j3ea0moPZA8c4DXspoB742+s
9lpILRbAXkqj3UrHnVfcTMYmvIVneq3nguEwhp4R7tq+l04GQsbdeq5Hdblproca
6uPlMb8LqcGkj8ftHjxv1tvdrz2lw3y8+lYlnjhMLgJA8D218lBibM2sE7XohsCT
hXGhlUxjj1HccTQ2wjJxZw130KkZU8ZYZ56f/nvlG6wyB0+R7oULIWBb5AuGxEyp
W6XqB1alTLc8EbnpyrajwYhcSW9cTZMjjQkWx03O8YY3KwrsHKAO5mxpxLDum02R
DAf/VqnBUUGR2RQ91xcBxESbpv9gOxazMeY9pm3ncTluLlfBEqZ6GlVlxDV9Jkua
2E8X5LOETexjmUQG2R7AvfDu3f4yFoMQ101s2FTW59VXLIUwDlYBQ9npyhCZEOUZ
tkuhBtpSKzi43qYpBSbP9AhZghNxHmgIp3n4ZwmoM6aQLL9R8y4dc9ferlCB6I+T
DdfzC+dLrrfhSeL1KzLkJI51+vMl/DFLoHjHIU4uND/7+YP/4ohGDnEZrm+SPQcI
Sb9QgHdcEdOrSKzRdPnHPKVrxxlxwGMegRD/JxWm/rnqKGRM37XicNNyAzjqUw0Q
pPiFEIAOy+T/QVZT6pb7mKnsMmfinS53eO0w0RohEpdf2HW9vRNGsQm10wS5rYup
2EDseiCWcrN7S4a4qf8KtJURVvx1GCDp4ICN/qXFa44gMRD34oUdSSZJDfosxXuK
941acFDwXjXVGiABpW0XjDO71KM5lNWBRr7KtJ+3FTqndB0ByWGVzPgLCKaGDI33
+ztECFOQqjXIYNpXLwRDpAmH1+XUMNN2HjaMa1BuMfWUVYA/33tdCOLxzuNF5qs/
gz/mdKlnl2UeErtz5qg82XBL2Ymo3sOciikHax7dVGoDM93cPYaMlZt9mXLMGalq
4gYsBLr3CkQsEimfNbjGavV3BOnn0TpV4sF8eUH+IA4o6im/p00Mo6tKZdmhVdkf
rFtnjCgObtQzmHsBzc74Dc1RE+uZRqvskF3rsoOM34Z+F9K5TzXZRmbFXFusZ435
y173mfeKWo7wB8HhN9IfqEs3RoxWfDxnD+30rRUiUZRRahp3/2i2iJrxEsRt2j1Z
iCM69c+n/bNbeYktgX/Q7vmKVgZ/EzbN+lumWe5uVsS9hukdXI9vppuhJcIQECky
J8zIPCIHKysXrtx6XeCgi36Asa5Wma9q25zolMrKBDNc3Yb2WQFwzz+fv4mzpBul
p5SmJZczVshL1jT35DK9CUZaczVt6iURaeZXfhTkKZbCRgtt/gChqCmQDd3Fliap
4eJ3mE49qqeJz2YmDpYPDooe1grbIn6ygT+spfEAJOdMV2aHQh5WBgP4ullPO/+i
85IEfrIqLsYmmyRh/SnQ2vFV3mbzER3255nm0yPYp2Mi+m9vtougEoBlXN3NbgEz
glrV4DqvOEYkldXoUBHJzqQ7TWQnsd8btaW0fx9k1WOKtbv4Is8Q6qVC3pnRiRWU
J20fpBUpkV3NjP6sacRZBN6Ntm5v71yQCS7opiGsX6MfrgLGmBRZVzIUS+TVBKii
wON66wImrviY8t6wQAbdmjk3e3nZrXVJB2AEqvxzat89L/VXG6DGOBKAjQFJ1bNB
f00rWujVNwBbubFz55gdj1GQR51HqAY2prumKAs3P2nNYBK87YKk/QiunueQ+FCX
7vtMrEDwj+ffNrwrbDLBSvzyYFcJIyGoBSEzq8RzBKuQm0udvsT35XPw/FpgRd4d
NnrUWidgQ1f1bRg6BfTyGRQWsxtPOUUBwlpJalhTDOOfIKCc562pp6FdZTsAyH42
n+o4Q2iqKxhSrraqA8hW+nl+0mkgQfnfPGVLpp7Sr/rLXhI9cxZCZuW8t/aJR/0r
nOVUW5LK5B96KsTqZN2xHo6i/jKTVhCaxMAc8jqX3ij1+0zefmIlgxlLUe/UptqB
u6eDHFjF1DHC/JGi+qPKnhyirxCmNUlY0mHcuuOK1oNNtuYrmOOz7BjvZZ/R/1KL
p2LxO34LB3V4lgwgJ+HbDCIyvyYlXKP+9CRhIIAJRK+5RZ4sr0o9G+B4cIPQ/zdq
ZMF3KtL6AbmxdftY4SCr2O/wALxr3v43MiuxqDJx8lbBNiY6/F13gEaHTkmD0BON
0e4VAttkvqFqd6RWooESFilkwXB9WMt6N33Yq+4vNZc6ukcxgt2rSDr8FBF5jwjy
CCSP6xzV8uUiqxmMXmViSRZZ2SXDnx73Dq/wZnWi0U8/HHQxBZIb+mpKuXucSnZ6
79wG951Ddq1l9qrKi1wZ1aUfCPjh6uD8+4D3AlvvFnQtd4fJ0Zr4qhyee32JhDlR
CphOAy814BlsrXuygXjLcPQtfX9kv0aOcC1/KzD7bwAaRcc4E2R3FqFvbFfqhlON
qC/WJNof1Eq6Oz9C2+L3MXMfDACPffCY0GbZFrbiodUfUEIDIZf5PsGpwcSpCb8x
MctoifW98YUeBZQUCsyVsxeCcUXnYaV6mlWi9oLb/Slkgz66Knla49gv74WX4sog
O6YgbmJhNnBxW2rPu9AmRrhUy2o407T5ug5IsifHI6r9buOhlMj9k2uF5EyGxB7W
GdoT/Czm6oBHjY5K5JBLQ1f3qy81lu5PM3TRHoDRJEM3N9F9FwzFNCW0h2ec2rnt
k2M5pF5tSMKT5AA0H8J2BIpP0Jghwitm27694sbnG90lKuH7DQYqyRfUym5jyC+H
pXRKxSyMY5v6qgPYjfeyaQdVnh0WK0KWKT/PopnzUAPM2aQrZOnwzIPbkuEsRY/k
NpTeBtnIYVAVkqFAE06ZILKLfA233szfzsJql2kE/7/MQSze4mO0TCwFdbmgTlyG
Up5JcxmxeW2bkPbaZBJxjN4jZejouB5MIMNynrCIM8Zt0A7AuYQDIxu6DFOmXvyb
RmPlMHn1dwi7I0DtoAjJ/JkQnssiscaW6WHWKhrqQqTPvZPk73ooQ/haei0Ag8uS
RUiwQHQrgOW1VBGEEDuO8KP15te/o/bk37nqUf3dBru4HJe2WPBgLU1sfNyylPX4
iKucOzOVxQYrCWPuOhG+loGXbRRIP5973h/8bEvG/qVSFnZxSmnIrnu6nr4JLbhm
jIk5Vkq5RFjFqNGHFk2lAoymNl7cavpYNTCshGGMJWswEhtVEcqx+K5cesDH5uAz
dWN/qTSv8J/llVRed80kSgQzj5E2oSlqVE3hLmNdQsCyazOg/GHe5aMuQq0umYFp
7hVGFlyE0ujW/K7Y+VfHEFTnnZ/mobJ9XOY/5OhgKgcOEM5XnXqO+MJYGQPrq0Mx
T2rqrqKhOSAW969jKnXMkUtU3vvett9JsAXhA3plFjKHTuSz9EPLaRF9z8+fit43
o4NAMZMyB50l5lTxCCnvPGdkyNjeu3ZrMo64oLl9LWKS50DAviDLPfu4EoP0a+gO
rQELLPB1h7Ner3tvL+M+pREnYHmmr5OapxDnjWws/TfLkBUSwVRhe1Cq6DXiFMI9
l8WtB79NvdRiKuVLM6DG7tZ82R/5QLJSAKj2SXL0s/MhkzZTz5JVFCapz3LKuA+I
4wUE77bO8qZdmNvBEJuXkCURmhRbGrHX/wRZEkp9gS/7IyejEdRjdcLV9fIUg04v
fWYCzHeal5iksb2bwb5ZhvaTX/7BRJ+8QrEsnUxkoOhq7IpWvrZWTJYVO8iZsC/a
nNehbYcHm4RRxFOqiDY8F5ILWdJwYpX8taljIgWkXuH2X8pAPwVPTmm/sW51OOs4
hQP0hVE4T0Z6l4SJCYw5saeSRayeVmFQzOpYwpzeI/mTyhBz8MVEHbAn8ZwZpDrr
caqwq6t57pUVzmyeP/Yoxxs6VljcjaFNVM99/aL+q/MaVPOsVK1U10t3lXwBJeD9
aFh/opjScYQzyRfHlwDCFMgVEKCSWtnSBugb4UjcswQ3nAVPaRuwBVodRRZt+7PP
Lm8ye8lMN5y3mRtlrXC4Z3nDYSdToQFxImNeCiQuM2Oa4S9iHK08rtRBaD9yGavZ
YJiKlBl5wsDm5fkAo0HxgBnLV1y2rypRm1hFKtdzCUbjfTW5+7W2vAAaXYq6yaQs
eGOgAQ3GFPNmzCsQTkjkYfSwJCHfnPbbmPZ1r2906wvagE6UPzHssDkkbtMndfKY
xiNO1NpxoVh3Jkib1Fngp/jc8Q5R8WDn8HVL0/uUsUpXMFOSBKoy0NvastAdWKwF
rGWTdk1vSvabgl9Y2uTDnQykqv/5cFYWXUBi1um/8G/+I3iZwYVZjDd1syvKcclo
qziNiDSw+18dYuOwd1jpvJjJIH3Dew5MnQVN6Ag8BT0I6KMg5Mt06C2SnKdiKbyK
AGmOGh+epxNRaaiIGuD/lv5/8u0oEyVM/6jlB/AM3gjTXg/0hFw5tgaToxtGq/q2
YtthMySPvLipXdmdF3PAxQr4Orsmg8Bi6cV3JScNApnu+Yy9KWiZz5QLTOmgxfoU
XlJjJFlHn+sBMBZpodWaN2uKECL0kSzW2fWltfsBBcymOE0R1Pu5MOLnda/SkoIn
uc085ZsNtqAvtks5SfMWsICjKsuQ/yblU/9QlgjBpESt+/g6FgDplbAF8WAiSjKp
tZ/4PtzDFj47hGyNocv2HmfOPRZZMbnejpaV4/ItVkYzXHqkZDsfnq5qzOuAnsvs
ei6uvlDHfLqdoJvYWMPeBdxYHB2y26paDdR13nvGHVayQ0/IeSAxe4z8rSB+Astb
j7RJ4jV33WNQAdi5OKhIBxCp4XxWzju4A1u+fh6v415w0FlIRRn2dDs4i64aoIoA
r/iTAl+UEw29z5ldNPMIidBiAVwObeqi5mWZdLObdj+A+6K46IpI3wELafeFjzfh
tCe1OvC86tSnxG1gAZTyHV8bkrKSUEzO7gep8tv9LJsQXAcyn29cv3bKoaoNeHN3
jBS+7szm6qR1cdEz4ttRDjpZdxvD73BEmzHFMqTUcL4pWMaHBz4iDVP+TB2VP+nY
3YcS1A7Tch1l0Pfm9Oe7R+7YxaGNtvhHUAyNMu+3/pQJY7IPS69rE/aZ7giVQXa6
3p9AAd7dx4CW8MXQp6wIFF2qUrrPtegk4+QDXSlXYafe/M/Vs9kdxNsF5kIiMywd
QXulm5z694Iw7VpA92XsNT0kop7AnOmt+wL4ysFWI6OB1bYm6Epd+zd/9KFz11Wy
m4b8TiK0xnH5u4dQiP4tXEJk20H/7hNmwtuuswoc6fZmn9VSu2P/FuBbo4amfhIx
GLPcOqlN2xY6nB1R6Y6Ph3UfHHCb5VFbgdhGWc2TjAkVqhDPxU7mDlQQxm/e1C7f
aRUloWLf7FXUDKyeT1+Z/4g/JgcZsBrEN/PEnjfB6NUvJeHBo50CY6Qk9uA4vPMx
wLrNUTxe1JJ0imdkc8kYWgB+DugJOINj00I0vDxdSpI9YrjuwIevulTaR7PFMLj4
Q+XLYx3lzbIHtWHrric+WeG98HEEqpijHjZ3zTEyFfE4LdJQtL3PCS8vS0T3v1eJ
CFDQZkBnZRv157j8ETnOH1nTa0ZilscAsUS/hTH663TyVqnX+c0N04zNlyRM+FpY
BG6Y6mRL8pCqQ0ScDIVl/SCzNz3aZhQEX+OE4pCIemdUa5SPxhrMk1Ot1jQsYkoA
TrnTzjLxnoj2iEsC4PTuylz86mbwkhGbxjOyhzJd1UwWk3lbqqrcYflOQwSfn08H
1Jcw31ENwKqtGZ4uBMuhGhBMv8p/csE493ck9MaMXfxW9iG1XB+pAz4DP18l4OrM
hHWYIV5cnOShBlODJEhPwHgw4g8KK0+cFZjx8NnA5OcchHz0ieOrEu0utMnKdwAJ
QZH6M1DKA3Ois8TV/QuYkF0qfyUMOoYNNpSpJ+2x3yn6z9unAyuOWLtoTBPc5Dvw
4jbzU/HP7Hrx2JtdsfMBD1bNEwTvW+bMsAwcU+0ygy23GPDzzhU2+N1bja7cUGHg
9mCnfHg9V42EWHr7U/Cnu3B0TKh4kt5yUbMduEEMCQb9e9ZTRcKmjQAxTQel9kha
sjfoLA1ZtLqK6rHsAkfEbqRo6ICRWTYj6AUdmy1p/guVb6LoY58cmAiyteAJ3Ees
exs+94j9DygrWXIpn6tRPXYoaC5pmY721wq9Uht80QjIKofNhnReTc//3MTlb/ms
aZhR434sCSxOzVXiZAR4JI0duBzse5xvg5qzskL8kPNJ1kSuRnoZ6NP9F1ZPrASh
ykPhfEWb+YtxJdupEQfAyLAlY9rmonIG8D3Xvi29jvvV0Pe74yw4u43biWg4UKu2
YxC3aSZZR4TLyOPlLjSFDrGj00NWORWr287pG6uEpqs495Ps14DnBuiamoP4kVzv
JpMFaknAy/uSizDNlrBDbqTRmO37bG0ct9JLb/A5e8TCKRcQVYtCtDs/0pXiS5Y1
CCyL9nJ4Dn9SudZ5qYkxK3EQqaGepJ4P0rtQK0MyLYeUgdWe6pXMht++wLJ9x7ju
3+CQizF95QnIVj0VEjGQp0nZ6hz/y5FpRSF7mk3Kv3MLeuBkaEj5ukwieQfta6uU
0X/tdhLcyrQ/l+aK20QPHi4/6Gp47rAY1HO5rzmti8GChg4Eiv0fbFXbsNQ21xZO
z651bi96TFklnAQ+9/vV+skpRWChZfet2u8m+qyaPmRaXrJC7Gn9WcoNvmsKgos3
NUYrsNrQU7TKPkANrPGPo6ofw4X/GKEPgtmOEAilMD7qWje5eOtuMij/s3kXLJAz
yof2txzu7fUlPk2WXlcL6WCNyHXQDteQ+jJWoBqJTC7sOagzlcdiHsfKpZf3pLHN
w3PxzuIBrXhmINMlQEXhGBzK6CsUwF4Q30NZM94o76lXlIhBLC5eAjpCDom/1jbG
7KuqhJzj/oi9MJwXLlENHYJiPvikoBit+62aO4ASCee+D7Pr4yZh1f9ho8vbvHyi
/r1cMqXniYhdYM/DOyuzTSCHNtC1tbQcswPBtDIxtFv+IEPjGABx5qFu1Jq1rF5K
Bk51DZHoHGVo+lbmmmCaqYYdyS6DQt0UgX5IP7CqgY1dVT0i9WKgyqHkNdKAqBT9
SvHb+yKvKMUf/sW3kNy8adbMwBAjkpTsB2qDETi8scutsW4M+0B8EqxwckBTLu9v
CLG1Qr/FX9ss32H3wDyf1nU7GgklpYwdDf/R0OjOEAWSD+TpU27VYtDgvbcTRf6K
GmwUIJ0SAbxNpXyLnUysLL3AByCJQdyaLsy7nWAjolIjYmg7o3yf5X7SJy0n7Jvq
3/rFCDhenoajqIql75kSLJgb5tLovBd/pbxpU7kl79axiHv2RN8m2CKaE8QUNcPv
iah6Vy/BO8+MAT99tqiIMR68H7xpoH4dkFkoG2TGWLnLXoNR8wQaXEOM5CpQt+Qe
JpCC3+IjL9JQYTPa1Xa/rgEQgkHse1qHJmAa2PMDPc5FjQsgCe8Kw5AfaPYQ+1uH
Uf2EWRFyPcIHwwpC7z3XMU5omLxsF7uJela6TM74i86KsGlGiuyYl3wvC7MTK/z6
QfXsh4lJm1HoXuojctrfdaOsQInPYwzbD7Il2eUMf1okRT7tykhv37FQF4l1BPF1
LF6wrreSKQDMP4dP7QER0lVPJGQYO4gjqo4Sep2RWyRus/sJ5JUlDj51ISPv9Sfc
HBM/ndmOFJjMAxrzcgrUGHYT8ofmSq8k8M7AfRRGvSDHEgrxZ/8Zr9f6pEmxP/SZ
sJ6buCZK/8nAqzHAl7OYxk4ZKOWOyhRb5UgZcGn+jLQ5NALtnNQ1Q2UwygVv0qY4
U8OaRxjP8xczaPkGuDVNgKdNeCflrmr978KUS0TPs5kEGu0pD0zoPZY0n1Wmlvsq
nZTJ11s2k2enA8p5PFhypGVPt+I3VCXfe3qptSSrgIZ4FV2IRifdebRDnczg8shY
tok+kf7YOjMkY+9H9K8it1SuqVW4JNh0dnMkMnk/EEoek0ouPxuowjOj2eC6oAr2
wyUQGyKQ4nFjx/JDLxSyVGx+NzZwwwOJJqvAsPgaQ0k33TYfq3V27xbekIibQIsj
xMl8Qnem+gZDq/RCiJ0LxYRBUsB3jfxvhoo7oM87CLLOYbsSKbpujQfQwt3i6ugq
K+jQpZLhWw40Mz0nWHCGjl2AJveNXtMvbOhVWF1F+kgrfMwSJohoLCn8iy5Km2q4
BCQxilP9uoUbhVLAPcqWPA7cwHZOmYyJHLJeQTHCxeUds+3uMHbPuflRJtzg3sK/
OOH+uESK6Y3zz3qXbhRV02AGEkaEYvzkCcPHv0xPpCC9OWAQJfLrzELz9sJR0p/g
AqDqaB/cfT25ex+9ZetKiiisxwkSyjjLgK90rH9QbjgQblEB02CC1E5qn0ZJ9dNG
Ufx5VD3GsRw+GqCBXrVCJEBjIASULbXTqwrn3szI/ieLVXhDq70aJCtCS3tnnDgP
drg4EefjfYoNXgkCk33gbdfPA+KAj3nwjAErjiymr0NjQcNB7mQ4ocq7g1BTk/uE
625nDn877bG2yIjtww/XSjsShy9BVyqymbM7RVQSaqkNseu49G1dklqPyo/jbd8S
t+KePWEcD4O0Edb1Ip5plm9hoOaX4QcI2NMk2jQgZme69PMcCY9YAOelSq8Swpb8
08cYNT6aIas//Md8vojCZNFMrvc4ZT9DDQougAY2T+zugcfwAfF6iTtnswxeXfCy
COhwfGXV2fAoKypJz5N/BJgCBU9T5CSpPU/TjMFcLRlWI8eeusU3XDEGBjzEfGNS
OwAxk1FFGjlTIJ7xuDDZm27UeX0pcsQ235UlIvSZlASVB8nXlCZOXahftOvKQ99V
qSkzEHX9YRLhxg9y/uzXb6VIi9gjDLNMqOzJekheMMPJLU7wKXNDdNRUee6k+1+g
FQS8d+dZaByY16Fe4aQkgkU+J0ALYvSxQmpsGLWrgCxnFRA/ObPLpWKqu9pnv4/3
jkl0t65YEr7ZO+Gpo2hN2xJUabNMFQl4u382a3Ij/zr7yjWZ7p8Cxj/9cr2E6uTp
33RNxy2fjbbMQ0vGKqaF377N7A9C1UKOrTaOc6cRKBVSghoftS2CBVDwY0/lnzkX
QNyUO5zEz3Vz03rvt1LR7MkXmdyTd5T0dPgZoRJ4FSpGwmQYEMpBVrGH2mTMXbcZ
yWDxYW+JVxvLo0+tnZGB1hiwN6ttWLcV8JPSRCpBeovvyKrCVDK4ziLJXbLo2ahx
CzQiKeMkUl7YUmUky9aqM9Sc5eOidlnR2e5OFfbuHzpdM4QK5/JYBXw9FmzavBw0
IrMaGT/CbGzxEQffpUnAfC4saTg6wtBjwrijB8WFzPvso8nmKLjpZX+x4T2Vz/jZ
8sTd4eXrahiknMyVDeUEjoRUxY9BDzwgELmcvvi6cUc3bw5uwWpH5yTbrkhr14xh
Vu972xYwKCecaRKQrDwl5AdRECS8lsPQHbI9J9nF/TZNxFeEe8CJyNqm8iKPAgrM
ihxChELVbB9MmyDRfqhR7V78j40zzIr8gSQhba9OV1rupw+KPWsVfcw8kdyT0pi7
iNDvBYHmx2sNkfsiI/wXnAn6OvO2cg9owVb2IoPyH6DEv5bs6zIdp+Av0tQ80Ejw
TU7ApDYQFaai4HYM9hsW0wRUkJ/m4OSBnAswBLYGv//sfokxhqOc/SiteosmFfBC
mjdUJoZnOaP+S2FN7HQoghm83g3rgTUuzpRhVQe6tWuq10RCj0go0qNuPxB+XuIx
yiLVI0R1PM0BFhGX6yn/V6rT9bD8QYXRYKvxFnG6sMNnOiRASxVuFr8LNxwmz6lZ
5puBVMw0br+rsNpUfDqx5tSfMg6isfRJCEDC6JmA9n+JQQtdbZ02WNWEieItxJNX
oHXBMcKuNideY9yFntGS9qSOTq9B4HPuFr/fxhzWwvi2WRaLDZZutN/N3bbRNBdK
LTsNgik/Fx+Qhm2N6VOrD+0DJZmz3q7zycOBhWjYEWjtYUN9bW7CdTV43tz2//CN
7Kyr+/H9xwWCEuzPXbZL0Zt0GussNL5B63hedRPloRyhIUk18gtNeO9jA0pOELBM
aBht+SyzveUlW+h5zjneBp3e2VFW/Lh/a985us+ukTZaLsW22FGJ+7aPYl9UsqJm
OX5DRvIhmQVEpN6MWrBtZdpHBevmaiOKgyFMw9LNkXim8k9lK0iwUntdo6+e9oKd
4WbnAGcOpkJfnfVbNosbBVsG3tIdnUdxGaFcLCBI9iXcG/4W8H+4hGS7DoaWUO5R
3cCxaxPGB4mxeRNxliimLNfSSdJLk9HwWK859pA6Gp1L74vGDRF6QnA1rMRlR4Rj
dlj6hM1shOJkPWUM9jM3L7MIfV1cJYOx/P2CNZTpJ/xY0YZGvQQLP74dPtKMFiZq
p0N8qPFYDil4TJOa8jk/B82MoubSaCqFxZ3Rf9ip6y1iCMKg4vFZJyYYVJ+KMjai
F9jE1koqgkXbv8xEVoPdGWa0jB/8OTPHUd5i86xZAmqRbyN+40WXsLaHtJ6qkYjL
TdXXGVpQxBMfDJxOK+3DHT2MmJflqYurzK0gVN5iGHvj/N1Ylc8PnjxqxS4MlPIi
a0lXznNSuYZmTTqr80EK/FCSet6tOrg8J1UbRHkz6mS9sKQOR8A+Quj26UrmWWgE
Hp9ZoGPq1q+yU+oSnNpUJXubRpl49OFnOraBjI2FIbss1xqqlKG7CKRajk0dSlHr
eIOlefQZr3iV/CCjPAa40KQ7AZmPly+x/pNWbHkxJE1AHyEHi7PkuvF9F9OP8DJo
saKFOZ6Ofq2Dqk2DR3RglpulITFQUAvrcvBjNSKkubij5LxxlJpagwzdUc1L8CJH
Rz/5i8s4PXIqt95PJ7IPN6esVZjamDCGN8HKkiEUCVPDBb3xPylYFq7RX05BIwUI
7O1QKBykaxfw4ipqozb1+bQRxY1ydjQ/Zc+XveUgu0vY+meP5bnPDylCx7n+Y/+0
01T4KE2zFBUmM85eBhVikOtyVzPI6Dq4TwTdOWu4sr7delbJroLO2BPPzAt/ryXi
9z1YyS/w1HEsYS98KLXD5qEbYDJHPjliP+/GxoqI19kvsJ+pGfVReffNB2mtbXtZ
rAkW7FrUGF54yVhLUhleUeDAMXkQ+wpZWSZULmSnZH4XFcMbxsIMf59T0+Lmy41u
7IDrenmYJjpZCqnuKqlu/bfgbHgdH9jUbD8LfGffgOLyXavk/blxRm7Kl3xXNqRO
Efyd9VXlKzT+PMNpkSTo/pxWcpEOd34mG+twfvAHbrdsIQxED1HRXkrcTQ4d7bc1
ukwx4b9S4TtSJh7tpGaZnJIZQ0lQZOBkAR0uGf57tc7BxmQuZMh3C2TpI9cXrT5z
daS4xxkAAC5NtWEKb+TCzIuysQD67q3a2GurPM9lNb9VTS3q42Gvh9WzRJsebZEo
iP43blJCnMXD7ZyPUmWYXwFnEmdsmxXri1p4VvLCb7Chn1DQZ1UJW/o02V0oiOrT
WDVgYKPO7STbpOS79mtHU7dkb5TbSb1xPKI82XdUnEzvVR+dJqeS0xcoKG8w6Njy
4jRGYLyMN8FLnRcOuH4hWtadpvXEvZ0XQzan81AwrhItNMun9Xh0r9p4LsWJvDCo
gJJqh0EXmfI9yVSI1LtyHsj2PKlxsnx0zaHwfnN2iLrN0Bg0ognUosSen0Bm8sa3
kwkIuyNzG7ISUPwOpPuGpU3kJ7JtI0Ybezi8e0M+Ejur1jE9LijTZj8BJ69W9lyw
QH2RB7PrUSoO0InLa2Gxx6K3/4jG0yVEpKzaIjH27RRTuZ+GvE5ZXnl9w8e1XJrI
EReb8cdJtBM9+lLl3vm4hJmIol7G7t/fepgCBoEmkXwYV1eVJTKIlU6fBBXoLwRv
zdqZ/whbuTcCh+miKCsPzJ+deGveYJFCCEu2214u36GFKr1yr4HDQ9CygFm5eHP/
HUl8AYFdCF7BQxi0bq6OLXN0DxP2VB04OTD+rlsLxV8r83kCI2BotyUc9q+/rQ/K
UMDGXjJCPPR6AqvV6Z2OJiyVJMWujfTnCPbgMDgii7sTvVWFufEra/t4KMjVQ6y2
yj/cOHeXvlySWDCrhQJDRg1QbOMISv8yQf7lIGhHuDzoHIzOnzRnMoi3yR10710K
DkNAwD3NzwfEhxZlw0Lhp207nQ9OiZF2b0Z1KrbDiKBp6mv/hE2XGKTkFpV2dSeH
VW8GUnAU1QfgRVbitQgm7pFK0w3prN3JM7FOo7ebgTC4787DghYZK0uzHPH8uHnZ
o0x23CGXk8bHFPbR3B9zsx3LPlikKy7ZJDRj5UrXKLNFCRyw229Rb4dyryPYweLu
Jlv97m6Rx4AWkAvYtL9Paa80DCwMVvmumEfxKoufoE8J0BJPLw/MyYkNuc2rACO2
Uh64q9GRu89+ho5q9/PFDpEdU+d9jzSSlnR5Y5BUNmwExXfGeK+DZnCsbgKObnb9
Hfmy8WcExmyxjGZDq8hFiAGmoBWLL0wMr3JcAcEUx8VABGHg+OxWDmD4W9J31yfH
6m8uxHcUxBwSbYE4cobXapvyNNb7v6mbn1Gp/lrICNGQb45jeLcJOYd128k3b1Wj
ty5rWxPExsTvYUOv0DVUzrBkY9kmb/nAmtzRwS79fzkPNM2V702DN7RZgRJ5oqIS
Yw/aJHS3EHuBZwYDKxubRvBYvZLxd9ESVmyA8i5r0w+77cfX027kIGIjU8hptFAf
/pjWv4mVnneth5Zk6e+o+bUf0v5ADJWssaJfk47VpWwVWDGB+CkE15qz2tm7k0pJ
E2r2zWyR6DuDg3sr6vDeh0rhtpUZS8FNQF4Jfd8ufl8OisWL1kzkchciDZZtZZ4D
MvUGg+wHl0eE4/oXcJ2YpR7cVcPLNPnzoGFPdfBhtuyZ5fmnerjW/Iye3RUU8K5k
ydyhQGUtj8IRpXlZtYS4/RaagUd+Mrt5EdmUBuPRKWSJIzaMxyvTbCjHz1fb8K4m
x15PA7RnxnxYo3BAs7Z/EfNJNOEe+HL8XxitmJb7i7I5zAdG0H0jzMcD6C/BMq/j
cqBGlcjgV2NKwI0mc8SoMUHPfbqfzBPzD4SUOhgKOaz3ckubyuHdDM2RhtwJJtxn
sv/PwVECFsrp6CK3my9i6zL+08JS0XXTic39mtd0SGu0j3W6Fvf55Gy7+zyPXy9k
m9ZmZL9jLURAwj0FTPmFrau4f/lutpa02BAHzuEEtWrS75hshp93ttHPMG/QZ7+Q
kiGrQ01jI1dvKy3e4IfXKerNzvu5QoqGmY58R/AP6umJC9Wz+0P6JMffDQU10P8X
Xv7cZu9uzFIuOCueT+2zTdidfJh8EWkj0rRiBBu4WkQdzuPlOAqKO6hm6ych/mq0
2yWO+k0vUQOZnNwcROf/msEOMQM/0uy/9UgB0NnxqC8lzni1suaCmyqITGp/KWGy
Nr6sHcv5HvMrM3p9GKQyXLdPGXUB+r9M4Kiy2hBx2yUozQjYPJzVTD/xOVsNPJuT
uh49BumGXO6+ey6rgWyl4YrmaqHT7QEXB1edvtbctE3dzl0RCusjhrN+jQbSTpTQ
+SNPZZQljSqfYM1xmZaNHfJU/huUg0UojXHdxb6FRM5nPUjnXrjFGSPTgj2SDNcg
098FFWN4jwObdoTyRbi/+jDZAH/RAvFZz3MByoupIFhn/DcP2EDzUeCCjHW+JB+2
AaU9Yc1GPf0lcK6uOUY8iSccXy/voOx2uUxa4oHevI80x2eInTLP5Rc3eO+FrfK1
DYwav+S3MQF/7Tc9UCRQAiIjY0JMmQBfg+j0ImaoOyiZR4HOizyhw8GuE2SgGNEH
jC79aFXIcopcXpBOaDXVOpWIV6yXn1mNMbj2qP1nnyB/EAHChRCn3gWU05RABSKB
+5AOD7OGTXTBF5VgmKI/1X2HgB0yrceXIPn6R/TkWrGUFLSpThsz84Dbyla6BBeE
3A5PcpFr6HLgbgbTgO3OGgIBLWqqK+kCE79kO2s79ZTq/+dNjPvtjDzmkss/VqSQ
XWtclsSss608r3n+5F6gTExRDaxQcbas5osmcGvg4tXr4fKbo5WC4NMMU07MzqMM
WnF0j7nFhmKc9FwHprHZmhpspAWMpjO/fsAFsgc7mcmqoB5MpWXRh4+h9z0BQ2NH
rTvqxSP/tXIeS/8IN5D9SO0XQgE68UtahUVW+MU0OhuuZxa7nbtd/0Nod30ijiO3
8NsIIBqdMSE7g4W9e1pn454vNM3qzHfREl9iSeLiKLDv3KP8EFNPXtLLk2MYiPkm
/CWyWCNl05Nev+41tCWvteAO9hC1tqejzGA7Wo3fxz5681pcn35a0F2PB4jBdJV/
oeDsVy1Wfrlk8NnCUPizw5HDXfL2E/yVJj33SjvzE5F77RDbdkCtxZHqGsd8/MaS
M9GC8GhfP8iLHaa4djnMSlhrN3TrL4IyiRVowQRThY66tCQDlg62ffOTJK5Vy6/1
YTrQG1tTZnk5IvZwrcgXY6ZFGoySV6zqpsoYJttPTvE0VkUk3WUkZHYz8mVfEEZ7
wAqOSPRrSF8tHzgvfy/377ryZCn+OiZ5LeQiPmFs4KiJlHzJMOhHdX+NppsIFzEL
fqK3Mu08Dc02A3GBTtCCdqXHfK38R1HosPTaVEN+Htw3D0zbR4+KWphy040TxliE
GTCjh5jDKKs9YSb2kEnPNVR6WAK6wZuDzmL6gDSx950C/xcKTMgrVaen2QJ63P84
rrNpgHm489N0hmFPWAqobWcIuxKXpd8580hNlIrZ/HspcyyorXWvLlok2e9kICy5
BRCHWg47mOozWuM+XVaqSc2BuKnIByxKurLZJ4J/6wxkuMiClxv59WOpyiU4Ggzy
vinj3CD9n1w3I5npH2XY/WIUB4+Nw3RqgNWOxx7vfLi6ratooEqnvamUGGx0rKKe
gWzJn/WEy5otEMl9rzMqNmZFkaQJ0LnuXGtE/OVup6oErPwVNXy8iZTqtoXEKCS+
45EmXNxwPTtBzf58qYHubJqXXPiNsW+k7FaUMRRlQs2RD3v9hUimolHLD3VHNWzH
ydBk8iHYIfomYACDi+dUNpQAtzJx/KWpeYde19nSR/eXEm0rO6xM4YcF1LWyVrPL
m7JcEQSJKSyGHbDyxaOXqXkebTEslWTFDttDPWrsQeLtHXjVaUiAvr2YAenRg/O1
1TuZ4sMdaWYQhg3bk7x1xDT6/rc7vRtVnNG5nvXxyHmGkmrfeYEk6SvNzxW9hFrh
9M9TogUwphcogsI+6CYU8sd61qei/Zj5PXOrjKC5suPMKCmI4anUMHrAsRn1Ipsv
Y3j5OZ2esp7jXPKiTS66DtZZbX0hZfctzaetDfPHxv2qcj5LHSwYvj3HfPXmPvch
np+NOz2ivAr0vQq6SpAIVi/SX+uxeFWekuGoo8Vyxfc408J4kwpvmaXC72aSNW7j
9gyqePaV7P1ylk9IB+R+9yfTjtv184AX3VsV61v9+bJmF0U3g8kH4m8iyV11L4f8
ev1kIZRSUcpmLLhHL86l2/ktw45S+/2fxjOQB2wr6i4GDzzLixj1b7BGJ5yegHfN
XmU3DyWkX+LORBIVBXPST8G7XhWR+Za0AaLpTJRwEuOs4MTtkTkpmDN/2A2/bALd
nY7CJdx4Xzs2W4Ga7V2lgksP56n1UbXf2qxRXqO4Bu3m7eLtUignky2TWUs19Gr+
8cGTB9w09TYORS3uWYql1DzlC+8LC5ptt9+K+wMzGbR0Xvd4ZqUR7TdjeRR+Wje4
V/9aRJ7oh6tQkcwT0FOaH3hO5/M4uPGS/tMySjFWM9nHmoU00Sfbm7Cr6bax8b06
sb2cMYEnfNzFQPaiA6Lhl6vDT/EnyAKchNjmUua/MPnrFGG6r0qrkOB9lEIa+sVO
pc7trU5kE4jMMxGkrjvmD54krjzsp0ztrzii/7XLZPaeLplIv040UaN1xHGGQbpx
gt/1+37SzqCW6lDpFyU8UdBEQr1Y0e147Msd/sW9IOAy+jr1mR3qbSOioQ73JblE
Br7uUy/S/1rrAmqRPPYwt+dayNbpIpqiPhKhWyP30dpECC/u7cwSwz7xKKM1XOBq
YYc8COhXXEMAzWe7uUkF/YA/HINKdiNsgSpruiDANKtscvsFE+szL2WXyXy3jpZP
BqPqpIL9WLpDyw1ogEBJeRPu+jp/TK23Zta54PXmS4f7peJN6m6oEjJGEI3Pel7b
sGrud0RVbFZbWqb76J0u0ZcnXhLsL5MMwkIX5iT0wZgYvyb9Sw1ui4RtWuLn+ml+
3D6GwjhnE7cXunF3sI718MbkUKk2VvTiozf8YudzwbCRn3uzvKJoT5S3oOt4hTvM
Eeod5RDXckBqLP+bAyOlr6O/va+ZgMIh9yFj2BwrI0+zM5Xxq94IQtu/a7r4lFEn
lGA+Z0Ij/mLFiiuOFyq6NGe6QckOtr6WnbqoleXIcK+1YWM8FGiyZuhkk4RhQMof
dlOe3fmbAfCzIR226P+knKdHZji7RBzN89r0GPGKh2rAZk+Jh5wpBsMiNrlcnR8G
CU4r4LYOoaBsEXLwt64uq8AcengQtyuk98Vk9NilgR8xgSlN1gGZHfIa8GPfWTQd
4is7ptJRmcGbRLx2ImfJXuzBu5YVDkqxyynSslFt/sZRnpvT+5bV4USvTO6bPdDE
k+VYwDLOtCm3y9Ip42xdsCPfMH4SHeS9WXjmZpKG4W/e8b5FngX00j3VCj77PCNs
N00Nxgiw7PmE/Cj11X7e/YWtKcSPeCQ/R29SKj7aVBAb/TmtAYsOFNMWoXT2D9LN
iIEfUvoH9WiEP9TyLatUF4N6Dzk5k/Lef5JzfzHbTny7k+aOLf1BICadI9wJMkde
w8L26hlhvGuVNTIFeJE6ZyTBVc2fbZy3JyTXUdJZN63g14/5LNFxkIRRXINEydY9
H6OBh7apRzKRbMd0P1mQr3CR773RA+aZKhRmyiGQwlhLPAVczlNu+2/Z5GFswuSy
vp/q6uqrK4XABDt38FA4LGwStRDYBgcQgxCEfqRs5OnA06gn9cfPeqXxdMC9kJMY
FL95xNhkJJ2rHfkSk2WK5Ta4M+nevThpF/4HlTM9qEwOOWRAjN8PhsAME0ZraXn8
mD0a0OTrWOsqxlUN3ZBsKpComRky4pxCesX8+OV+M1Vx00SMlbk04TBk17m04yum
ZKYjq9TTLUPoMl3cy6JLUNS+XY7AnZgTMPyU6yX+QuA2Tmb/4SMxwnTFOTSDG1m2
QIcjAZPMumsqpDWrLiQRw30hYiKlpUa2ro5Qv8alUJwRMC2HfGIckOX5o7sX9dfE
a7UhWgx6PW9+5Y6mpRzOI8uezzdUFP8zAxVugBQKX2MhBr3YFuJFj6ox1/bJoFTk
XeALPg9MLdK9e6v8ouqnXyOzevgo+DQbw37WjSy4Bz/P7+RwkVapw/1t0HT+rDSa
1t5UwK1n2Pe8F1w3RT1Ws8WzRmbCFxg4qYtHMhiBiA1x/ANMrJm6HBaSWoaLMvz1
gRrpQcmEcNtgF76Uld0VwOwHB5SX9Xm6020RLpp/Qu3DrUk1vNhwR0ktx7ss2Prg
bTD+COWR+O9D2YRrcwihX1ww0OjnWdnjPJ8huCpmIjsiJnQKJ7B2SWEcLN7+AHwK
G3Q+1OketfVKOYuil06dxIVxXkoJwwvDyh/fCfVUnnMggo7Xpgbco11zzln4oVv/
Q9TdlOGlIqgi1SxMOUK+uVHga29eiJty+My84KW5FSxduVIA8/YUh6YvNOW5hP/h
SkSwOygQ+ouJyIrIIute3D/4XdBGTaJmxhq/zJSctF24Nb+HWWjMl+SsKWLXNPXm
5s3DXNslhvhX4G7fks+qFpx+ZpbeGy8iM7eMVKb3SBWHV2z1dLsns/J0UAnzdBeO
g+zPUmfgDE7eMdKnyp+zwYFJSseLwbJspMPj80dn7eAjnURMUeqQkgShPFUSAD+i
bMM7yzmhVp86p3ufTDoksVDxAHKBv7giudFS++KjxrblxuPzT0pOrCe8re1avsmn
Gk6ZDR2aCOS++MZVPj3uQag75KJuf1TRB45AnMYjSEy8oaHubuj9imyl5G0CqhU1
5heU2qcqJ7Pe558ogHCc4bBwhA5jb0Or8q7+E3PUzE6qM6QVcTdh7ryIpYhchB1g
PYv8K9pFz2r6H/Hazd455xpNkOtChzaePGqUCNehrZCNRZY98Uz6T/7mV2R1Ae3K
+GvbfxQYjpayOqOw70ej5GCVkn8Ao4Q5Sj2V7N2TQYLIWmR+iQeluGfS69UaalbL
eco0AVIoE61NZ3y7tlj6J9X1nhPQoejG4vv3BeCdgsda+2HeQvzO+NvV2+MmLJRK
N5/r66dgE3yhD3g/0D9ckCnXwrdFPs/GY1DiulZ2UHJpGodhNa/1oOsuuOI4heL6
C07A90VhD1yhJBJymXJzkiu43BsTP/gm1eNxBpgFgc5BG0IKY0UpeMj0ETgjncNL
qolu7LDw+kMtp6OjNuXQ2RPYE4lLdjGZHcZ91qJSMNuu52MiFmWJ0mEbj6lBIv7T
2CbGMTdRzyf7ebzJ8o8JqZa3ikzfJu8LKnOkZkNYGY5PrNt+3jS4VgDIvI8aiuBP
imUZORJI6wRWyM6EcPbs/naQFAJCZtvGPCqn4l3cH5ZcmXtrSELe79Qd3VAdPyrE
YDWuZ8fQh0CVeKMCnAZjA3GzzsfxZqGUpYqmORi8XPSQwXYKVsj7OkYIUq1yV1Td
zI+uGRyBwYdSfot9/ypczIAEwo00HRru3DSxX4KGHklGF5IjxYgeBrz+gMsYYbiL
kSlkD+grBAQNHgPsPqagKlPXPiud+lYwYcEJyOM2ZQpXsxCYSzHuvNnjLfzsrO4Q
Qi2/rtdfkJFe6fQ1lBfitgd2y8ZqbDyEuYCCMj9AZdSpqZfKovIZkTNoSIiTQIl8
fbgR45nu9N0zekqDfhKLdo54ww02fQ/aloqWVTwjmY1hEqeju3JMuXtYZbAC5qn4
LQpwtnCwIoMkOPHh9wge2ZjUb3tg2H7yhrufa3085MVugIC+QEWCJW29KbVNpX3a
k7FlaZzoBIJd4DNKghyc7BrWwvDA4xLMoh06Johlg7Hk2PEv8HcqBdJWUwpyEF7W
dNBj6H9avNqaC8M/a0ZcSVy71NUCXwy8FM6CJLDQCZOMZEX6fwUMD4hJ3vApV/8L
VLC2Fl37WiQc/Q9d8AhapaFoyuAL86TPtfOOQqQ7NBi9giTSF04e1r57PZb7PNhN
uY/6xk3FsqUlD0EhSPNVYu0UwAzvPch1aKEPRzZY+gBSagykyJSK1F1+GiyvhnSs
1jmJsZDnmgG6x9IU1fNkFr02VH7GN1bkBt15Flu0pK57ycR8BrpsQvy0VcvpTcYc
642vXmrowRnnNDxSZC4+jI7XbYX0WEHwPNKIM7xtsx/1AWJ8aTAr5TEaKua5sb2U
bnLPxQaFBPi+YqOQ9xaWNb9+X2qumoEsUVdJvpftqPgsLzzdp4OUFIZ176/qga66
QMlzr7tU6piSPtRrzI0QN49EuY+S5CTLq9/woFFW+HO4PwxVBnr3BFXxVdZoAxrj
B3bmIGdLfSzrTmNEI8rlN2B9YYCEvip7v3OkOIBnmDVfp/K7CsrqhNQhrsWFamUh
1zi3NMI+OGHd87o9U8zw4Ei8Fb6+O2HkM7gzAjFcH8sn3q9L/83UqWqBrP75RF2b
HJf18wXTvYpfPWFxe0bGT0xPoMpppidL/9reoxN98Q858oqolrC6mp/rhoYtf5fT
oGOFBRlXjUausE1FGWfwytXgiGFgpaKOjIeT2MgsG80KsPprZawtpiDnxNPp+RND
xRJEjix/QC8spdsWxZ6XW4RMluW0wKC1vdpJsuTjmanaRL0PcflL93uDFdU14Xe3
LDyiBx4K04I7ipRv4xAL+9pxbrxBvZSTjTWmhLu4KRkWB/m52q5Bd0nbx4Ve7Fnc
4GEti8vrRDXCXJWY0fLehPrPUgKBRN1Q2puNDHd9AW9CAYjU3EYvaHf0d+J5ILVW
UfS7+Ty/XibCGmfShYZydMWS+6N8O2C0DPtbvRtZN+ACsoI3//vX0FUMTm3x0kBH
LZEVwlKKfHKqdgLXE2tN7rnR5Mn4ZDG6XncFFeTNd0G99ui2ZxOi0avphLhZUQe7
WB4Dk9AR/s/hWY5emJ8QPGAzzLOsM8D8wBDzwfEIvjrTvB/5hED6UkU957k1sCfC
7aGeYhw8c3iuOgayUToZY4Z09WRPeQFTiVkf5bFabxkbb/QWxkInqejGpDzASfzz
p9a2alPc2kfmC3Ss0aioXCx9MiuwPNRdeKr8HlmeCWsXJHI+beZ6JVh6Hc8mXBla
v/vH+mSjO2mHfcjRsenyf43wWKvRdmjg64exijW2nQ+KaW9b5JflrbrI3nnHCcRR
VcILXzikIf+gNTeVCfsXoMbmAuD07h8TcVJMvIHnYzkdXX1BmazyzsQltLMV7orF
urwStY35UlW4fcO/A4709bf9eyX4TpX06lBgm2COvr2oCn0zIjjfLxZI31uu4Dak
onrPoZnccdalBKdhCLXBW9ZVBhhAnaLkY1YnZku1G0C6BZuw5fc9Pd/aws2ZmH8M
u7/7/P6JYXczdzNLUXsJDi2/2vzXxBVWdDKJaicDodoppwhrxNz3bI+fVk03SGZo
jTkpznFQMM2qr98k3dtHgUR38AipwCCwbNv3sWNUMwsmKhPKAG4B+0RpC/j1mN1P
zAQg7dFxDcc5aM+4Tla7ddT6exmv1UWm9p/vMCzKRNDOtwakv2Otdt7StNRtSNZV
LVKeUKeBKqgkdcR9oTLoB/pInj3Vke9c31ez9tkht4BcqinVsJW8fDF9x3yKnrlO
3VEEtly+ZiZibp9qHI1MbiPNcJAgGfmHL2mac2fGx3trBD/Rv+/yJM/0+b3vOyKt
8Tp2II8nT3RI/K0qKCCrMlg81ciwsFQXsnzrKXuilNfTKwjPBWO/kWnoI/RQfu+U
znLHyVNsyvsUgMEg5nHgMVpKFvZbF55JvEjO9DJX3KdvusK/6zDPn0eGFyK327iB
4ZhjbvuTcj9VZ6hHUU2iKrQ54scwAP9iKv8wID0FhZk5SaaHRkkjE3kQzVWxTmPD
5HL1vQ3JuXTgub7MUoJg70bENdgVPVpwT1rwJJlcn23GRTKvns73uUWNdF5bukbA
ujaT4g/pnusoVCTi++c2O4pF446NLyBYPlzguAbj4u35HZbWKzTBXNPqbWQ+cjDS
eoGm899/DBimvQdAR8HURp2A5UZkvWiMPda7e3H/+GuiuFvQ3D6ldmc1m12592WJ
OHnq7CE9JWJpigzLTxKyegF0Pft+h9FFyEYdhiTIybEHHAishcwcsXYFW4CMX74K
LRRlhEx/rmbkr4809kn4a0yS6tdhOmxeFV4LH5+TH2L8Pb0adEOxy3DYdpuB7m2X
KPiIcRKTDxT/lsWVagz+QaC01FE8MaCayZErtnnO72+sRKqvpvv9cbag+XQvuxRG
kfv8CYBcNgNoWmxWUKxmsylr7ulnS9jR5cfypSHJ/TZRXDi1Gw9JvwimcBhzlYJw
eK1GMLfKuxBh95hO+ZrCorvw36/hO5iX5giW6VCowYJTd/j9x+xVEoSSKFz8r0MS
OihYd5M8IUSosMRYan0pokSdQXFv8aR+FAXcalfkibBnvPUmPTL7KVw82Za5Nv+I
xDFnq8uL6mpS4lqG6hX0TneHLfzS3M7bRPOpvqgELES0bqEn9XVcRCCIDdp6ATvg
lDchAHWtIHkPXQAVeBCEV4susvSprs0tvQwdhdYJQ4fuuOvCvw4JuhD9BrgIU4jf
LnkdRfHAcWKWgLvg3srMNDOJ/GJqqXuamOpD6Snwd00QmtZFp0IgKr5Bovk49y0c
nFtdTUF4llS0FRKf/Mzc3xEOUxEWE08P3oirCg0aOKnWXVeP3e2WOv+Ni3M1ACcK
BFLludhP/BgdbT2Kyo51DXZAPTvnz1e81dJOnHZM+xFaPJoL+XbJZ986IsWar00x
8dYqpw2L6FUB8wa9zPq2oUuLQdZXPAreioez1ehbuxndaKFHHkSfzdcKmRZs3yQ4
C+l3Etifhkw8cxEdHjBoDTVwEu1gd+aGM4JmeCQgOTatj/YV3rJR/M8kVduubAqN
9vo6YTd8C/CloGIN/S2CSDgbWQ0enypTd5Zg2cOhHGfDki65UAs9yeBnLlgswWM0
QiendaaGs6TVg/HBbP2PA0oUjuNxOh9wwsk/NzYX63tMXo7HKs6AKyqem+jLaE7U
iFHqtQ2aQ3bW85xBeXlq6LeYV8NGzZn15U62YUx/DaxtOriC8aPE2Nb3BeWsV0U9
YwmWerXO+TOVExOwX8I9Im9slid1Az1cgcV7t8UT33MrrmVgAf8RNCqFsWruVXWD
/YyS4t6h5B31YXHSsAoU49M5iwz4naF6JIUMzbzuwZPC6ds8E3zYnoQ/FYogpHqC
mb2C5pNmackMqa6RfFO/jNW2oPX8cIICzwM3s6JCt8I/8NpCsulwB9JwUxfsfDrZ
61QWft3usggJNxpFLLEpTr4EfBLrG9jhDCFk2sxoM5LZsANaE+RODFizhkT+NtzQ
DhWdtNmY/QmDzcK16lgCc9zzgFOTSLm/EAZm5lnhVcA2/ezqzm6R5Ny7cLTzcmB7
Fsr8JsCBQ21QnDr3NQxZr05OiIDVav9Jj4pNW8UW0533tsXYEBEBZi/lLue7ULig
oLPk0LeYbrKyDUpe8UmJtpkLLAJuP7M4e8bg98HMjoHCC8U0Kx7139oje64p9Ko0
Fnlztg7ZK0mP+AiY661ERMpkYLoorygNIGbtizhk5jO6MRlbSizTd0V8AKTnv/a1
KjkMkb/iIY/A2/NmOjHiC4UihhzAGnwSOrpVim10EgziqinIiVH8+Nko6ifBn5K3
aDENhgq1Rq2KJg4ni6A1VVxcU5CZVsAnt7f0s3XonqLExJNoXQe63kuCS3zFb3ub
dc7kzx1Rs3z4Q8rylSeCkEtd3sXI3bbLKS1RY5T+H+vECdSI3V6HjVpuB1wmw2e1
oTk4Wkz5ibEu4pT5/aZvKIvIszLTfPlNhHNGdRIuFHitKPMZOvDH4xSM5hA3LNo6
TwR9l6BefU6roytSXqxkAteVyaWDwSQirytfF/0lfCpHjMuqpwanS034ouCd2HZ/
gY+aIDvzrcKT00mnyj7iRK98PrXgoVYVyxlLC+XwUSNPWJ2nwr2aEvqHHB8obF3l
m2eY0d0PlPkLD4AETyEB5wMM7M6dx8ai3jNOJ0pH8PDOV+5k7JkE480KYAEgS6C5
8X01QcuLdATHg9agCSeVHx5uOAIiOWviQJC3PSAtfSqzvcq+0ZAzkAe4OCrU07UT
yHaIR+VzcmTd6OY7PYgN1UGGNSMHu0aBi8IV3BH0vwTN2XC/Nfe6ZW12x6Rq2A3g
6mpUma9R7fW7zL85nuH6hUA2Uuq85P/p5BphYENUTRo82eps1zp7EsLsnEzAWtj1
OMObMR/aOlVbUL2FBpJdMlev1R3j+cB+MfSDW8SNYLqs76M7NKkGFiXhh1LcptJV
AWbvxTGfWvlf36l8rQ5MM+aYV+NeZgdrbaaCb6H/AwI3NokX7WmFCJHpzRVudl60
dl/xfEGzFgKkgoLne3XugnMOJVxz0/Mb/tLbAJ2UMzomOg28yctebUXuwDafKkzd
1MuFfD1RZ6YqxE3jVL2+RqGG5FSiLSQSTWHMhcjZmK+b9hPkl6y5JW3kv4u9cK/9
t2VQY1oQBHhRQsU39Gg5XSsiZkTTF72RzXXQYicHQF1E0gUwNlQ4SCRDVJ7r6szn
EnAPe3E08MhzkcjWzoe6Qe3igBfc1WJltzNW3Puqvb+bOxs5NCNawto0vtNuI0d4
Yi58P73ns4Z7F7PGzKNs2rC71EbqxWYqq9+/7UoNDJIOTuzwL119cPLxR4+3tf4V
iWzZDmSDK4QQu/K4s/sSFiKSn5IzOW5wTTru5npMvDikDMNo5nLxT4B4UqXZuFda
KKIjfu8s5Rz0zGaajzzbCYct/B6vCv3tQbwyOl47MJpdjRhHHw/dp8LqDBEkW88h
A2/enpnQvFOrmIqz1Pj/wx+MzTM5nBGm61ksqSVSWrkBzGUj8zyIFf39J4HY0s1M
mjFvnkVWL+2zMQzttyRpdoolwVdNoNVinRKJX+8tWAq3FHYdkDFVbCIXKBu0yC97
gSyC67/7sjqmFzGKILOV3RH5B0N5UTUdIYIRo/CEAu8HAQDrjXFSfTrjNrn9+/XU
GJyIpPvZmFEX2I1ZNxklIOT5eHl8YK7NMIkntdMVoAkelvMU/MX7vS/vjkZK4vyn
ze8+/5+qpCu1FGxgT/GzqduUyHCR5NMOCYQ2eEOOntGobyBWBy2RxFnHWEY0E7n0
hYRpn0DVxdzje4StHfSFoWJNhVQ0a5F7ptp5bkF+zqGIFlPVM0O9D5ZvNuNItCdM
JdH/+XPSxRVKJlrNzdeQ+4/8YLuG6ggOffvwG3wN1+vAznx9LU05y9SPWN3uSh2D
trPhfxtTKgEG1ZPJMBwcoriT0jKuj9DAK8aFTW3yx9S+1SKHwyW3COGt8CJVbR6U
DGLOvBaGGlxkb7H2A4+DQ8EZIRLEU5vxGdXQxpTm7kqyGMSWEF3ttt8B8RyP9Ff5
q/d13uZRSriUOb+pGTu6sqRfZip5yGSs3CSom9ZPmsRS19IVzYpMzbyueWPYglku
Gce1+3e/wW8uKPp2C6lMtJx9p3qffhQtyqzTGF/PlYT8SnG9jN6uFT6vU4thRCM1
ZSfFmp/d0LGvnYeNeVcNTEHGIzLBJpjhm72TbiA3gRcgSB0jSxOEScVEC7fVp0wA
FBRMvcJkGG9SGnekARytswwrEMPg8BUm78fM9Rj4EYAzNHz+yvcdlZwGUJIAJ6BU
DXAszqi+riPg+YJFqsA2Grahg+P4xpR9pKwwaUP+I/6ule0bu3W7L8nJ5livcrPw
oSKbtDSVCLa9jGMekX6ecYu9QI6yICOq1/Eq4qbRAINKrZCx9Xs46hBk59O7Owo7
zgNOdq4gWNJkLjQSR4t+NmxQ7k+jZBygsdH+Cd3pay12SttX5/JX42ydtDPvvpjx
N5r1kJmMdMQTfoNtZ4I1NpLpOVRToTFcQGwLvmAudlQ/AE0VvRMED1bXiilBA2tV
yx/3rclSOlN6/xv0u1wF7uE1Hz2CLtNIuV7xF9DHPrV8OBd9dnT0vg3fGBcZTI82
fqv8qx0ZgPTiegHnLwJ5agCadRwchC/cwbzBzZhJxfQHuMbdnFif0cIvhXVGdZ+d
HT0OUnBG7N935zKCxChcHV+7TgGkV7WMrgdCaA1wliWcLCjcTZIo7tJSrFgKZpwq
1qhQTRKUgb5R0lKIuB1yUHjsDl0xCaViwtVhVBNhsyHs7wkUGJoG6Ice0OaTvBuV
5pQgbGx0XPyZ+pPbTAZIOAhDmFBYa7ZqvlAh0GPknMrqSzL18MbkO5sYu3u4KxOM
mHxVaNFH/U+DrReQGjBCgQv8XL/4hjFh+XDNApgXxfUtudCsDwZCo+WOq9Ym/ZD+
0KjuNGB46XvzDEN3UwkG0J0ZHbwIae4npkK27OiRwBzDlPV/pcweKsTjIiPvrjOt
UIfh0ePE+XnP3SytiMUzCveKnSMRGlAw7+IvP44vuUHTicC6oG/jUaW83BwbKa1V
WB28mgsr8hP9hKmqQgsSLa3Q6aOBLMWnSUg3moROJeMmRmedd3mCRCj0p/LHPPVy
E8qFd+p2L97h/7+6QxntDnhXL5qgpyWG3EDm58ynM3lqhI6i/gB1XarG03+GhtX6
n2AxJYoP8j8hI88r9WDSZkA2vRHvzNtWiOeV0ytsSr+F3/0osgAzgjcA0BAPz9iE
6Pfp4OA/hjNJGVfRqM7R0QNo0XV6ArjGQ6XSApfPqTFMqqc/8HSpbj1GOlM+R1wE
1/MajgUL4hh/W+pxPU5CTN3aF1F21fAnYyJCq1QsCrfDRdprR6t36kHSiVkZKQhp
Kv9cn82IhAdEQ0Lj5Sl85dYyYLkCci16L2qixa/ewxELZxi6n1jLVCcoMRI9ie+n
DP+x4L5SHr7aIhjk3sVTB7TCxDkWQ+H8lljR7LEeCGi+6ZgKAo91eLA06nYP6IPw
/YDs6q1py0fTxr3tp1W4tnTSsHQ2XzowAu/iftM2GRQT67RL55CadzhD3JENvwix
EQZ6Wbw4HbJrQ5jAT3w9lmP3vnERiA5i63DeixiRJjlxSVn/sDi776BZzXw5k310
qqgKsT/mCsSKOPaAt19gqZ038rrgMDksy+hUAncK0OHqrtebKwZWbj1Hh1yEh6aC
q3oncwTq80BxYqNfxPaflw++W08KEj9fmOlXXtRsGjDZmV6sHifvmCABfOqaojZj
cY+f3aqDkeNvezggW1u/LLenPlP6SGuurNMQT+UvLx5Yx4iznX1EDjwdGzFP/EQu
3qlOT8ts52ydOXDfBIAHjvlqN1g7i0v1FxLtyxHpwh+l7LVmMYKN26uF8V/w6j+c
4sYZIP4itF+9m5YN1cDCxEzVawog8e+zInDcLJQYifF3vo2xPIqnRZbAgqB0wibH
LApMb7A2dAinqkb2bfVPizlSUebw78fbFjdejIJkeYKTfxYqaRyxahaOSeQ2Z2cc
ejS5odtbczrOR9URVwsFSmzarR/p8Qibffpb012FuWnQUxlgvMugMVjMdfMrQzqd
COf3kRym46tOpy+VDKQocY1O3TJx7EHEHMBv8St4nyRSUNB1CwWCAAZeCLo9Y5oN
YZLj2AThv2kPSOzjHea+iDLifE+MtxeZOPa4MGolCxTWbh1vwlUxxHC2eVfhgMzT
6+BGLiMqsyDm6vS0ZfM0MSIVdhXSmG/YcuL6T1sEZ9pPY1W6w5oZBcPhzCIB/oZd
ee8Oh59NgUHnstrpjL4ElZBp3Fu4R9C1R9nMZdxtuZo+bwYR7KoABFlHzBoBqolb
PiX3fr/+VFIie+BWJFHkpZ+H1gXrMWbGk/jN69vbBl+EOj5t564ZD8Vh4YzVE3jB
uTubXJMhpJ8EsSbRIohIu3IwU39+UTjBy5Mvzy/t017Ob4zOBUtMe55Z4APv043G
bT1tdEBdC62BSKZBSL41hmx885m8R41srlRYR7rE5ZiWoPDB14z13y/HXYbSXxHp
o5gnCRDUQhrMTX44zzZFDwYfAadPvwilVjCM1SdmxzgbCbLbKZJD9g26U0zdpG2+
5JymZlzyIbiVjkmYrNPWx+QcX+mR/RWRRe3oIGyHHdUX6L5xaHhBybgkhWrvN8Zz
65YiMoIvNbVKzeZSmGjhbvgkoNGAdqZFUM22+Y2o+icuELZH1hcPqkLUdprT8504
7sczdhU83aJvu2n/4JLgOBZ6d8ORKZHEgdQNVrFG/a1XmUnIiFNZovSWrzXzqOhy
GpJsCsUo7gz1M+psRY4Xd0E0vCRDWWqc+hlY5Luhyd3cNaQSwZVm/t4iZYeOfnNb
80cbUBpPbb7YX5GjQyfm7xi2h3+XIr8T0UPvxeJm917socoFRrspAaBZCCXQ+W3R
ZDKPwglwEMuigzvr6a/GEtHMWM7NCz58jG4nfFVvJYvJH610IoqLtEXzAMA9LifV
NZYcDM3hssZbjmG/wgwo9rb2+JlyukjomQa5+kKXcCDTJC4Bkx5xVSxk+pJqJojV
9RoERhxJgnsg8gCUNxFYjsEJ0vlavzy+2Kp0Pot2n5fuJjwNkY6NnkVRxja8yXAb
aqBkSyYkkAIzXvqXaWkrBeXNLyOwphFZSlBBh0BTWITQRF4js4TIgqM1gp8lc33N
fdgnIj4ma0zqgVc3p5VcasKeR0lclXRhKZ3oZAA/i3lCaXKSrJo5NcU9BlFKj6n2
zR0hxrTBpKYeIoW7rVZzcdkVom+nv2O4hJ7PXAVWgdhE0aL77m9RgGToJRBO7wGA
Vp1IallPI0XHUzGiEYsMyerbxhvuEk1Bg+lOD3A/SUTobciEQMb9lCLL3KeMvQZ5
lVsoas4S4zM6ZhuwKjcf+nBJb4oseuLB45YOqNBCEUUKghOnhsm/wy/Em59L0Jlm
IOE++gHdZ2ZkFjJbU3e3u2Q/lBO3P2E3mhzFZ2fqq06d7yAd4fICWhiWwDa7dSML
5mEjqChhFmaztpA6BJgZVs+RXfB+K2A8CFreFIU8b1b+SRTvl6NQPPZlE65Hp7wT
OkUkdy+10N8iE7IYoGOaedYwowsVAt5DHjvvr+FLWI6MzcMtZ352wOstMCR5kx+7
/mcFaiS0zLaz8jU4CogVJZ2wU41ZhN/yWqsfbGL7iOtZ/YLuGMCFjiTMmtgD++Yw
VHgK2TvmhTPlrElyo2CZPISSyHEPwbiYTTwhw/mDbUGr4vEefFuwQm7niw4owz/5
qq4VmrBh61f7Ecjr7HIAeeQVLwDXWruvd/PTzt+nzWziIP3k+A7Diwk/OKEs/ZK4
Vk2ayF31OBZh3rT+5xQTd0x5QG63oHIb8oKJOjNNwDNuegDd/fEFbUu5l8++6WZO
1aI7QnSaL8GTJ417L+MikWsZNEa/WJ0Xp4/5xvDIUEd0Fa2zutZ03rRziNILBGoy
b+BWLbZonGQwa2cYze29TEFKxXZ1N9RuQji0o2DoDlzJ+h4kN0aA6x2C6O9ZK5DO
xRj8leIwkfvPzrM5v2JwBJkyjGtUK9obw4s/LgAWZBEGBL4qu3BdL2wJ54ctLJqo
0OzZgLdMK1MSaEIVvEYLVA8XG7I6EfdrheGeVE0Oa7uNKk+KfQPRVNdxFwAXr6po
QITSp7ah3PNWIfeyXqEPNnMl3mEqkDu1nHxSURHKGl8aRKFaMNqkxcTQy3DHNCVM
VP2sKqcVIkROKXX2BhuOHJ81Y+JroEqnWhvca8nRJV8q7LdCo+W9ccWJgJwXmzNq
AvQgLXDF3Pcl97Ltvv8K5vXsCr8C9PvNta3YzN1bN2kk6pgoCR6VtOPJozjIVm7B
2dBTLC8lVyXviySojDHQru2salp/9oLw1buvJILVhiC3EnZGIX16BiHaXTsDYsJL
gBqXhbdiN0lBMNfBtepwNzuhh/SY7TodUlxpXN5/Y7a4uMnwp40nX0kR3m5wC2F7
FmeFUXZSlkLqlwmChshZLn0fbf8HXa+0QXsf+oVvzCQ3i1jJjy9UhC4jz+MVkqF4
s//tFq+B+AyW4Cyudzvg2V7arog16BONkZByILv9Bnj4tZQllIXx1LkiNaSlHqq3
pi7VVRM5FETVXUYsGtK7kfx+gAodZKiKFlcdAvAmiH6rcjULHf56b1y6j2Z3rdIx
qzAjQV/Rjt82JCmXxCMpkz7HlpVJY9M5MVXdQgCZUVirYYKIWRz2rsq5dFUAtmCV
eSfBL+aAFWqAayRBztyHCXBMYdWGeeQDfFGJlpIa8u+d1HQ9nDxVMPfvzQSoiZps
SSqC2hgnxjpoayoSfCnVN5LCjbrtlxyzNATUPqXgyxFjh/xNivPiW2mmPDvJAIfn
qgRnb+DOkRahblQPZrRtTytvvOST+z1nKhpsSoSAMPgCHIO0ll+/2yXgV8lnVJQH
eAYnZ3y+ArqxFiiVuRwGgDeiTWferCawpDCAKFefKsK36BNvaMhoNbwo79bYdnFF
SK7cKuj6gzqYO7UtKoSinu56OZNctfPYq6HzfYuJqBIpAYm7WALg1lPRn8/xBsKD
u1iysITiy83bTzKzwB14WuenMAeBiDC9Q/jY5wQyYPRBMfQr6rrEfT7836n4En3Q
rKcPJ/WCYWVHMWyi61Q5UR9zi3YgduZU7yt61V+cBLaI97Zp/7nDCdJ86gss7Efg
Hfa5j9Y5OEJkYK8nih3Kc6/8xBo6+qgIjUmwQAC3WbkAQ0lWk/xOdMAG3F/nVy6f
jBgrk48Y+ODEsDJpMsGu+c9T8C0UNW+12ScmRfzFS1I1EociQ+ARxAuP+j3gi8Pi
5JkO4L5EG6LVfUw+V4S2mZKcAlgjEUbGXeiDrwnDatlFTs4aJjczSfhFi0zHXiDw
MwL2ZFKNg4ERDdTMnZMRR1dtZTE7n12sIn3NarcxH+qUBmuAmZza4P7Y+rS0ilxC
qSqfG7RE+S8uQTANyZJQITWGPf/O4QBvWjJm2PtqoDinlPYrSvQ8IphK2stLmmD7
nW575rL7Xa4bFEcqVYI590ivVfX3rXjRlINXzGOCuKy9v/P9qi91dmbxSJzySV05
Vt6vkm6cgQCrYCs9JgD/Z2gaB9GqbUixuUVpXc6EUsnmcOjrSLTQmyJfJPQzUa6f
c8KrGBKuftwTa1r3h922y4NBkn8R2BwoZ9pBoIM66Qe4SqVqtyJ0tvdOQECLlov1
Qna1DJTHqTfrdqHOuyHVIFmgpUNhWNI888eEG/pakM54d+3Lt3AMc8191oqFDFRp
944ia342gzKdV7ut4+qOGfdXfdBVYE/GZAFdxmzv8Et3r++PGYJofaXXmIMLq/jf
sVS/IPY8RKujl17lkMV38dZJFoclRFBEM4Sp/fOP+X59qDbeSu7bz5RxeZFRsGP3
wjrwUBaITonPBdx+hrWhVU0J1qfdZTk7uASR3oh5TFoo4EG+DqUQAzW2l2Dy/WnY
2yPgW7oATq+ZGZmUl8Grq+bj7rY+KS7PIw5z3f/vtQ+jMjmxcJXKufDJNDrnBFzD
1+ly5+Hsr/Cf1izHNU9RS6aXuqghkPHa4qay2dlYEZJgTNZ19idyI6xG814LqiFr
OX4GfPPzD6ZzQYJRnvAp9BsSkThy3O/4f6OPqkXQO5QCNIcSj1Yz5Q4WGfB8oO/I
Kw24ghXdgBgWQahyYeqLV1FbjqkB6hLpqcIOrimRR2AWUOWaF/A/gfJh/h7kLVF8
0A36inhXNq82hetwyam/L9e565X8jlEC8oKnTltHc4UyxfsuiN3b1sqt1EO48mzM
DOr1SMkzLvVrXM+ihc70+GhPtT5Le9ZKimGs5cZ2yJfmL/d+5+qYSQL4wpBe6dda
SjalMBLsoB8afOogaxkpDt+7C2CYfLnEgiWwr2C8k0Y8BvsQCrgS2sWUoO5QqOX2
jy5wpBDA7wvNxthqeVh2DpLdNx2qm/uJKrcRqcbWamPKYQGDzOS4sqYvepud8Kak
q4jk1eGElKQ9wEhtYAVAaaXNGciV8YTLBcrs11ZHXP8CiJli86uupF9KpFgmOaQh
A4TVHnXuOOPnEmNk+fG7UR3x2zXI1JAP8Jo2BzlPyc2wty8JluToSt4Omr0H69UO
I3RvZBZ/jZaumDvbX4e2PhNOqif6KzywKYmTZXpYi9WWRylkFpF2LqzJQWN9gz1n
Ty0wna0HprE0c+oopFkIUgIO2pQvlIMBICwiC3vWj9EXTY4cc6fnvZCVE9lmL8Al
XfJUyuwALLXZ0DiYLGbW8rKNygTI42CEhfgzwDDYcAeVcr1pAZvUyRHjDy1S25qS
Miqj8B4LHiZgiZoMPHwaZNHSReU+t/M5DwWYrkrFvYMKpL0N4+enloHEbA2reu7x
pxvOzYHoDDEfsgczGC/2CquCJt7AcRqQrbg2rrt6Ae9/rGTr9a04CI+YXHR5b5Tf
ecDEWp41y9Ag8eWeIhQUHj++nwvab66lEjST0yZymdDVw8SMUiq0VuxxvFpBNB0N
s14F5kMIdYKY9DBHlxLEIKI0T+qUwshQfJohUx1//1YzMeM12dQ7Cr4FXaHo11pO
kWCeet8ziERiKcK9EPOZRdqIqodlPp+5s+9SvGtwtW/oBJP28r4QlE7HlGwXT1ml
/nElIFAHXY3VXFcWOnRCREGp9z1S10iTaH0yYkM8NOWK5gs9zTPTnaS0HnokGNmZ
qv/ZXfGwVTxcz0XXyw17r11gLyBWwn4NHg7S2DqjGmPcsQ0YZgn+gOamMrDwJ5TD
8G48BkjyOiUseFB9cMGFMCjkjBu4MBjq4bfFMmmpH5KjIA3ePreabgHgxGKL9L0N
jiqMKIvtFMOf6bUl9JWOTPvVS11efTPPR+8K+oRUXSnOj0HH8RMPcYpc/D+Gf1fA
9ulJR1wUz6k/ZUUmyarci9p9VeXdSAg/yTgIdUyN91M7xgg5OLm5HFX6xJKHTNsh
Rs1/7AHA9h/QDsCCQQymmz2FLLtA7nRqoy1XS5ETa2d+DVS/8cxR/BCGKNMwKpSy
Wwd6rINbPjozGBpVzHZSIM9s1QIlZOueVMM8DE4dxiMm/TkDEBMni1KC+py4555W
5BJIkigm1OoOzxU4GNqzJcowSGKnALo/fgG9C9kJOh+pr7szf0c5V7CZV3JP8CX7
uXwQvlGNll9eyNIDuyC1+cOQ9OmrwgSNrmXpD+FU3uLtr3jHGn9ecO6juqVmPSpK
HOBIWxd1pSjt6uRS6za70Qi5Fk61rmY6fZ9H5csk4F/E4ijwn3uzicpGc1TVA1Ag
nmu5IE7SmvEeqk45K0QY1PyWOkYV9Kaif/39pChORjCLoR2Bew8VFcbMMtAZbyx6
dzJZ5jIal1YWiZLTXmH7o0hOSQu3amD+pGXe7pF/Kj5usAFrota5om4DNeF6jVmk
nPdXLhNdDGQcv+xLwdG/frx4qeJui9rgRATSceB2CM3hBfuKW2HLYLPBVmltoiA8
lHmqFv4wL3nPHm79BZ0joeSKKjwN6eIlW4YCDfE2lHigsY1SnBb+TtmzNMenS4c2
uTSmXvG8H4UxsmhxoS54lICtD+qgzrfOEInjM4Lsy4R/4a6eC1WSUF4RrkDCkHX9
jOMmH6GdNhtIaH+84KVv4+w1t+E3ZzuhbDuw1JeYPMayvPyLdr2+MaX/1qnCR0eM
fjcz4dnGpVIxqhNK4Pp0yWHZFSQInMm7jUQ7q2kMO8MO2J22Vr6lodklc9Fj9zg7
fxpa68XVfgM7OqTY1OuEgCXUP8yvh+AEcdikWj1QcW8AfNfBjVr9iGaAH6SPDXqk
gJFrw8Mp/oOKaiXQZmSeFnf+UkQfxq+H5KoACnjMQ+R7ZmMFE2rdFK0wKPVE9owB
OJFlBw/yGg/AvO37BmQ9WCyyiUkU7xCfakz1HKVbheWxd5IWzVyUHQ4UYjR5YxPZ
fT9AbEi+OYVAWAsQFoXFkolfmKGACWMVy8Uv37hNCkmKT/hDI1/SfkO0w68OJRy9
bYnnkCDBiezVPgOoUUZPM9ERr3lutdAVO2rS43tV4ZjpOhT//7lhkIkoo1suSMkp
mkJnHQSWNTnAyfp2fdxKD9Uzf8IgYpjOeZRqvzwnUu82r/z8eRLUTEJy3APoaEPp
s6QOjWdaMZgrwES6FCpHDb9YMNG6ZOwpivWRvgJi/1Gp6sadF+QBTBQNgiKikZYb
judAnJZm5gF1rSsjyxy7sHFZw+uVx2Ma7UK1G8Rw4Hil1+8VykU+rFsd4cfllFf/
95L91eNQk4nnq61qhzlf38HqpdBdKaAjwTgAir+0eJPnJqVzJDc32kKxN3K5KCLn
NayPVbSW1dh/pYVyg4KTjIkA2f+o34FDRXmSCF197EXRyH3WyT6HdFVKFZ3C8RuT
PT3J8kqWT0NiGlkPVjVqE9ePs5xcpmRtp97VNipf3O+6YzBT0ClGGGr/ZjNrnfmd
9ohQTC6GckoL5apQu9IBp/hTF2i8/4Fvb9Iq52S8KQWxSFCXFJ9Hv2Uh8O1qYPWF
kNz3wHHgVeUTBVpDokqGzNSIY2rltgGWKywEw4hEP3B62Aab20KLJlKHGtVGThOR
lH3nnwZ4y1CCY4E+R6A7F0SvduuLbk1VvWnisfSWnBkBazxmncbtA1pr5w6l/8le
2s6Dw/HRT/jqzxbfRxWLO/4d03+aSMlE6n64AE1u5sY6BCvk90BOitVTXkNtAwih
2no8TQv3FBFywYUZaQ+uauehFMmupkXTcmfzDUcPPzW4/HYcL2hjTb1T3t6avVQ+
qs4Xe0IznWxVrZfXJZ9LnDywPWRUUw33vIIst5rnmp1q+unSl77ntPDSRoy3ga1i
Cc4VoFogS8vEQoqIhFpP6EB+LbBVdPmNm/pvZUzkKSyWWnVbQSGL5M6J3kTB6EE9
wgOYP4I+o2l2zk7BoiJ+mdskA5P0PKAHR9z7w7YG8g4OzMk0argHOhR5keUj4WKh
8KDi4D2JRhgcfmOhedJI989L3Csyv5XqzUeyvZvAX9L+fFwNmDm2Bgt7ez1UHzPT
n1NBcbDmywC7VnEwk7eEXqpjJyYaVkcGFSyrOjQJk/f62YvWCMFalRbUcAz8PT6J
ZCXHJK47dAQ5oaHcUDF9Lcx5ZxwijupXjETp3NEsEs1BRCLwV2IY5Z9XrY0854pk
i8WVaBphsLLWDILeFklOWoDLDlCVKzEIdmHVWtFGSzLe1RxjmE36tCzL50QMiKOC
c25K68IEiOCAnUhk2ZXI2oMwEmCdT/81yiiAxUvyG3tXo30DGuv8aWMEbY6kl6ey
wSTjtD3bfZGqdN2H0cjnG3NRKVwr50IVIIMOk20b09at5Gm1mcORXO3YdTo4Ujiu
WDp1XNfkCI4bTwVqKZGje4xImE5+7sRLoLt6Owo6fq+iF7v9ZdjROhQfv+y/msKy
c6p+Kkl3wKmbZ2vszteVLTUf5kUhb5l9xNpTIAu+nZHaRoHBmjmMIjqG+ao8Fqdd
Ev/+Dh+LJTGrKf8hQ7175m422g6CExn13C+xG72f4uNjEDjtJf3aIT7KQKjyqVrD
+Huad+c0m77OTFDnGXXEzUizSe4UXpNgZrBOdRgEsMVcPTmKUdNX+Qdc8LFXjVi/
i4MmInLElVfxrVhfYBH4ICR3mKvOhZyP+IR5w44WlQCarMpEEm+GOv2dPKNMByvF
q2SDQi1JGh/z5nGEtueaBNOnKsq0grFzGP77FCs9JZRF+QcEpG9YxmGDcWBllVZK
ZfAtYNx4iQNjjUNtAceYEk7lZH7dyoX5QQrp2LfcTUftK/o2gXR1i6gpjJcyQZIb
43bCvkPAwSWcouLRrLKBRJnA2FhuBr3TfJCp/C80GxssVVS8MtN5JR1aEcScClnR
XefQIxsfcBU6nD0R8swuad76l7uVvPajRUJa7eiC/clWiimtbqwqIUZ8doWCtp+T
X1uxR1rd2HSVbcNVPVxR8ASaQNHVpgLE7Q0o4n86cnASK2ZxuGnllsslWhXsvJAQ
u2afdEhV26W2Teg9r0cJYQLVPURfQlDGGNMbyyA+KI09A4+tcCd4Phm0njL33eTK
vIvaM/kxEkDtFPHl80TMd4i8oBNriZsvJjWxbIFvs+xgnyrNThsp8VbJ9MjvkGef
LcYEXr2iABWkebiAFqtom3r3Hv1nlZejqAN+8GozMfZdzYh6Yxq7HUYtmpoGOyO8
6fJZNFRanIt1ARK1kNrl4GZ7KEy+Rf8n0in7c5L/lBmK8X95m8RM+NKmAI79fHDM
UapbQZBLNR+y9Cpe7EOYGC1LB9xZw3L7egC4AsJjp2916fkp7VVUscu9ZLtlIYkt
/AalsA9kMCp9nt6tvLh8XA963o8dOBK7tA5rOLP+j0rtqU/euMzN3JtSVk31D9CD
SlhE0cyxxnMKXS71+FH2fPgg6YFTFJLM/n1Pig3fa+At0ZtF+FPshRoF8CCdmwEj
M0QD1VR0uSi9mf5F+fZbAu1rx31z+OFEwWskQ7rI71MOeIOMc1g/472fvBnTupdC
ux+P8MgV5tiQJdZzgRUMhsaOlzSqFM6wc9+Wr0Dh0B7RqXGGOZf8AglSQDoX35qG
zRO9/0Cc20bux/uRyzQ86XSFZJ0a4rPt3GNtcdEArMDMncuVMjvR/yIttvthDS/u
OAT7h3cFYqMcAOl15OhLP0ZTohdSNIebucFdQjyBy7827baUrYQFvUlZJqPKspm6
oavozFMDFStShtFLLpGkNxfrLoP0dEvb0abskhsNbVD1PVnkZ3q1t+0QH9laJsUR
6jzQsQhxbETD8A2RGqwXFWvlTGh+3ONUoBh9HukDnMsz24z3ME4UI2PVnO7AIV0K
fcGxPNBxncvGFz0PMwyIcYAVfvkoDakMZeKf1+SXY0X710AIpg28v7o9SNSxJf2t
b7VrLuVadutscQMDsFKHbDUx/eL3AQIJuDOoox97zS17RWtAlHTRMpmjP6Ia0nJ4
/v2nEgyPJr1mmCFiag0HPz+Bxb79TiCS3NoQCN3qxGaDYshw9WCsTEfsu3l4u2QE
PJeIjAb/sCWp0QWe2AUF2XtLssYqyqVe50clR02EQL+uYxWxrJupUAwXySIOsW++
XCJehy+mU/h1rllP1kCzT/H7DJ1h3B6dLNicmPSYSz3/5W+7K+b73fg+5QR8nsM0
+45xW2MuHJEtFNo3qWGs6W0IWDJjbpwGm/3jos9y8p0WRCQUnpFM+lJxNJODe45V
KIhjJyPCTSeC6HJW1vfLhBuWIPn9kllK1JUxk59RLoR4B8OicYdmoI9BHIkV1Fmg
vxpJT0fpSDqkBgDaQacDIXCHfbvgkMT0nPao6ESDBFpt/zQDJexoatj46pyZL81M
91KnW8px6gyjlqJCpK1uC9vWRebRAQbEw4/wc8XzZO5ziPWh6+Xqk6MdjJCfCEzs
us3peS9UmK93IVLMIbS7BR2Y+jvdKqRnqF6f/Z7gOef0JILPmmX2wC7H6JmQQ+U5
VUACEMH1Qp1Y/Iwe+EMSoHgur7LH4YcJHb5ZSPesPFEvYfveyuNR+Bli20WRJi1v
3v3j4iTCLQL9s2O7f9dtFVxUMUQRKl/ixRYKEIGkoOypsdM1uSyhEJjGJ4b8R8Lm
enA5Jue76i800u36DO5iK4dRFvPQCLFGStQDRNj+ceiZnlabPRa9kyccOT3ixl8A
Zsu5/roPQ8Ojr5ufN4FClJQoad16y9aJdcMjd40n3JvxQNcaKcAw9MqAKZsiJkKj
L+68xc5ZI9zGiVYH+DPPYN1rWM6MdrvEXEePdgecNSD+zPpN2Dbfneu9q/9wj2kB
JWiT4WYhyoZRGFrPOEPCB99dizaApHQ0zQb/rBE+cMWLzd1dcbKN5wi/VCsBB6e7
72KLpvWlU+D7+fnlddga1Fe4Rymhk05UimEk7H3e8QtWIe9AGFDUGbd6Lslukw7J
VUb6MK0dPcsTosSBHZnqrm8Quix+TvtGcQ6cT5rMCR+L8HkVhkxnhQTXCAw9GC1+
Ra38XlBXn26kmBABmIDvGxDcYE5LlmkydIlhCOTdzCnPajkEYheFoH1tHQBzMHWR
qsq1BNQjv1FKTg2l0+shKlo+iO8+sd20Dt9E0Q9m6k2MQniDY9NT3+X6OfQ7ANyE
N4nVTs7kiQll7bbnHXK+Jf9cMwaPRp79+2bKppR1lPjdIS5ObLS+r38PlchUmjWV
oXlcDAVu5suELhWa+nYeiyvVSwEJHNEFPq5h+SA4i3s48o7KUjWRpNLN0a86umy8
5+aB/4PRvv4vpW1lk2P3YpTAjgKtESYFwte1doqaEvF/jmB95jVoU/Ta6a+VT8Ee
5srZXRniQ3Mt8vwhLzVZxAkbKTo0PZrqZma2WS448n/eH0FqtxWctX8hTCXNhsPH
JS3jOI44u08cVtok9homscXMRy3KEYWv86HhCIxVuHko89yKwxkpqSCjrYucijxZ
5sjT+XoTDrjMmGZbcoDqofhcjtQrVxI4b8lPSFU1w1TL5gZeYow55HJxAuRCoJ52
qXlAK6T03M1TJJOI9LBaahQYWma/qqsgjvqkJDlA6IKYbYazpskmwSEb/c8AU1UP
awL8WaCFSdQsCOJKDPitLHXSsTNP4FQCIkZIV2gBeB5BEfKLorRDJyvvDqxkLcYI
F1lodTI03skR0enYrBpnh+lwbzzgJbwTRpdm7Nt43Tk6hzMLGpZNx7wkUevHqICl
CWsEBkncREQKb8a8Zx4H9iuZFP1auWUNirdkcQfJzK0eWoJXfbYPazPiwAwlWA44
wlTCpJl3ep9lhzlkBfvFdW9Ej2wM5mtHc+QaCuVieNuGxkYMBEq+4AhQGQ+KQqAH
9yqK/PGf+jxlOes1veGPG8Sp1LfEnFlAYl0hmVEkdfOjl0BUmtjtSNDfxt67AAKR
ne4+mDsJnztVUV5fP61biKOuC7AyZ84irp8xqVAEEciusmOpsT7bcjddD51fS2oO
6ppIpspYAZOGhtdL+hjmkH6ZjXGeGZUP8i5WJcD3sZY7geVS1NYg/ooJ3BpD1mLO
GdaBf2Ugf9imZdEPCinuIXOrgLEuRljG1p9UUNQKDm268POaBqk+n4YIrvQItpoe
ShtPA0S+BgZz70lJnnpGzJPAOoGvRlfytxYF+SNeWO/jwdqYvCn0p8OQR4rQiw34
OIZtJxF8dhfXvB4H4c9NrYront5l/1e5KDmxDonrotcqNLNap+euXZP7UxLizK7E
AnbGrnIKNyI8kr9N/tH5Z2EfI4Q7BNGcNNdl9oMTh4mjgOmZPTHSTLENvJyCoxMt
/+iVGFbSNS5+iPBcfF+LG/Li+wkt+YRoF4pwUB33nEPowHLFsOO+/bWllfkM0OS5
vFzzu6QbH+wwHq15w6REypFwksFlbwleAGbw1TB6nstN8Jr7AE28reRDQ+AW/bni
vPbJefmiejRzozNbwl9W8AkXWLSBE3d3Q6GCeS120NkH1juaF1pRFxsjhL0pmFIW
SKbGo0wwar6YaZJ0DZaqxdRg+TNpnh2eZ49ShDPyxFAUYB+qycLXO6r2RCdaa+JT
wAZsRRAdS9v0vT07clK+Y+1Q1brzPCEAmc85ipHnp5Mgo77BtH+vZI2XqW2BkcOy
TBfYuntcGvBAHYXszkgOqjK0FN+hexAeXZonGPtU6cDk7BgIaaafpC7RdH1KJlSe
NbT+vWaC7ohePXWT+y0tC7LaWzjv6sygA92ZRnthILylurNHibWRyzlIrxbZHUkt
fqgjax+NIwEefzu+7dvQJ5PU+Pl23ctuEiLoOZEvnxTOA9gjSPCIJP1zzc4JE+0W
wVmGrCIiYZa+tSkgsRiY9qyO7/7gKBtl3OLLAZu7fQXduUYFEX+czitQpM2O9Dyp
9nmEBmrOIK8vMCSbRrA+pNPQVk1id+xB+69+ueyOWHejB3A7KgH07FpGuf9YYjZb
0Mk/O9Y2jjikfWhXQh8zGpdhGnRZiSQdUiAXODBbHygtgt8UNJbKPBx1sc7DuSx5
CmzGfiUCKJbJyFROhKjufNkWq+klSth/XrmIRvuk1f2GfE5S93Kq84MHeLc7C1Fz
UNiNokfajSrPhtKSLe2V6SOr6yCA+XfUMrIkVxfb0c260sGcfQ6xBYpYz5Z4BcBC
kNdeX3e+S4tnCrByZ3V+9I0W1wLgdUFb41524+X0XMX6+S7mpTzk4vbryH+mJ3ie
z7gsfE+5LKq8CNtbRqIAaqEj5KLYzQ6eWRiVyBSvRWBORu2jOxCZNiIgvB/2KscX
WiKzemgSDjHGUQojGkC9JdKMap0MyQIlKnCKIBtfYm8lYeMzSEGjiAEPrREE14Cg
Py/Ymcs+poS46uCwVyltpM7WgcEFvTOwuvjNSGJawVMXmodGrji+k02u5oAbBvud
usL540KJDcV10c/T7J4YPXRSawHXQMjfiOO/+FTLn/b8tJRYYEAD+fgv5lHfhtQ0
KRGpegSi0JWzBMTnbe+mpWd4oqAdVRM/O+B2177Sxh96oYHCTlpEdxzm3/rfUyB8
MBLYOQMT9K1HRYBquWV9XbkoW0psf7yhRDYj+WeRrRbEekfm9UbKJI4GWnAHRaPb
qCbgPw7hLNnEFfO2Hsmeg7nQIacXzTvp/UaaEJ7PT6oHNW7FO0ww3rdKFN/5o8DI
nKB7BsxtpAulzsqtxDjO12EFC6Ei86uZmVu+rcNSlxKm5OPXQHqatMEZg+ZLmAth
SCTSfMDTN4ZlPcQV6+5rHKt3iUxlXIW8+xg9MYSgRW36yOmDAVbN2InUybC6RRqB
LabDmxI8WfXX6eeoRQOKdU/OMlgvj1E/2Bv9pMCtfJDttwo+CyEt9g7e4beVEmqM
1zijZ36CpfJQKKV0w3XktnpE2xwmDEQ3nQm3vd4az2xhryfsoXqJ/Ya4CoZIYOlJ
ErslXishPwGnIbIJlVw0F1TIWKHGIfxq3vj+OdQGlTlVSdIMp3yw7mKdkPTOfFea
mvu8PxTXABFJp92e8wgkcw3g4KhJIZ2teoAJ4tYSjTtNNcKbysIZRyGKJkphtcUE
mLEElMscV7d7ll1zMiTVmkstWUDBKU0708IhrauB4tbhVpOM4MBX6iZKoBINVfhZ
fb+9aRX8Zoiv91PFhpaQ85nSEYbAPoNj3QyrEayQ5oqucelgS01/laB8+0eJEpx9
pLhf620+om5quG8VOCv3SpZVcTSGk9mjX5LU6zUc9NByrQyHinx1Twku5U5HE7kp
VtrCfoITrYka/W2T6261WbMb1lp+nWSDqRxzRTlIyruuUX/o8lSykqwgfvqMiHRM
FNS///XFQElkthBWPvYWGcjTszN/To2W9D4KruQAZsX+ZHU2m85N5zKglfyuHpZX
h3vOPFSoz6xnwp13swL0NrAlgqpavNlleIx3GkTDRrHjHjcjpm7YBMxzzeIox2U2
TMjLBmdJw1LpqOXyOU3MCDU66QJqilnYoz2s5sfiwycrX49uIKRg5yqeSnkAGH5/
U9CtCppEZRSlUewUh2CKUHUVbyStRamSlI1g8zOqyRLTjr2fns3IbVmQzVVLaKYx
GCym3SJuMUlel/vQO5vkaDcYdVD48MhPllzn6ZXnsY32vr+VJAr6Lb+oinLZh/vb
fD9jmsY30Q7U4AYlWo4MkWldM77ZzgpTGBc3bIQ7ahCvS+xYqyKTSFTqEhxHqjuP
naiFFWUPJnbRs2XW8ZDuFw4TA/MsSwQfzmCPWEQqTzyB8dOM6hFDepikB1AFgLO2
7I4VLep7mKDrODk7xPQUEXUcNvHn+v31L5VUPn6rA9f8lYj8a8aG8lvO4MbHgE2Z
VSwDqMrKgt5iUCmFzI/ADXDCSWsxMASdoRRMWa4kz089WTo+aEZpsjUzxrPRrhaY
NhRuALh96Xd/IZJCnG732PLGcO/i91g+D+gEsBUIvh138D7YNEy8215MVuaooejG
NsrDXAOzlJl079McM78fbqUoDLGgWUKvZw5FkeXuAabJBdPh2Y2fwNrtdtirfZCt
eqcuYx3STtUQHIvFTL4DQKWH/yUMo4bi0/3JmbS1HQksoQ87ad+8UFfN0MkLumnY
1cLANLbaDPSXHLXRAtxTOYhVs9fhrLZDmlWAmAg5MWUImxkT+TOvJ64OG5vj1vIZ
azw5GX3qCjo+ZpWt48GEA6F9F33+08v9B2PbNaZd5JtmwsAGpJ4hAociwT6KQIOm
82jvOScR/ORPt5Ok6iIhX7WAJPP9wAuJO8wxQCejko/W50mY2dhklqFWASHogiWa
5WOqYmNKizbnMYNUOCvd0M/uh1IsaOSwQmxiPNWXnAmlLA32zgFNRFFi5WJby7iw
26Fn6KFHsdeb8Vu1gXHr0I4E+J12kqEOH9j7CFidlQIZla4abrjj3WJVqNPOoc2l
RrHwmg2UjPepp/DAogn+Sg+iBfQMQnBP9vHfozaWH0gIO2YypvWFuL3fuLE/TItq
fln878KzslA2RTaAEUwE5F75v7Is6uD6nvQ5U6Ynu1/Opej4JgJ3qzysg2aNKVJ5
avnVixQafTMjxf25GUlaXEiqxFagGnWfrdKIW8iSqFqV2WF/ayotymdHJ2nYAzDz
4l34Nx6bVBNTH/Oohy6W84Q2K9JJR68l9ivIlySQ/ZpipX6Oskthjy7W0UB0O/Mn
+/zsexfDtPhAcmUpZbYwp8ltrlostQWiTm+SniJvWVld5zacAbRX2qUaLauWTjny
Yvz63fyreCn1TzoViF/VXbFjjw38e4I3l2Rw9IJOioHRD1MX9dTGHWhKw1/YdQ3h
CHr84l4v70pBKtmNZvhhfsBN69YPJ8+JG9iM4LLt89+eP4YYKFkMrD6HHWw4TrMS
z2FVfS3jtvMuMgLi10itBDT1bKwEvOc6c04FCryb8/jCfgErGhFpaKkKsqrwQr1V
QTqw7DD4tS2/0oC9ooWg/zmXrOksb434gF+cOu9y6SE/uKE5Fm3/hh/0VR5JD/Id
jIUuGScD55dO086w3VDIlLHYj0dudXXbP9wYNsDG5+j7YD6FvZpFevqX5EgKzgOs
8tJxgNO2mj5HZ59jGp//ah1o9Oobo7UVfBXT/Qh8PgDmOZl5QlgZfepfjqcytDjb
oGgQWGz2ZDRubQuWpnpPlrWUWfS2H1Y7D/Xkhd73dvrnFQfDBH0UGWPbqz7T3OpJ
skRrMNt1lKjXxiuPlS+4p0RoxYHJ4z7+xFmR183UVVrB+WoG5IWrYk5VKzuiI0/8
EiMhgwEEYmVil6JGset4JjME1kkTw/vgM744CHglYeuir7Y3326vTfxuO6Vmqq9k
P3lE762mMHtfrM3Thxgj7fVMh+LUR1mJhvPw5CNqPwWWayUBNzIeZrZNbJ0hFCsp
hRVPxePMk3H29Ur+iB4d9zw9EFhfhaa1n6JfeoAStV7KRnHvMKDyvmD2p1ZZALrp
EP3qBZjIOAcHu2+iTk4E0LCwKjbnHhLUAiHReQ2qCA0aAyWzkrwRY6HGHG8iaWPR
3q+bSY4hisw/09akfX/mMLvLLEk4IOz54rHrW+cMND1rNl/2rJv0AxKIuVDjuyBb
HQ/H2k2UTPZTMQyaku4jMkpvvBH6zEmU+KW5IbRFgQ3Ux4xrxrhzRLnl9xkuQzeJ
QNM9qKqN98le6sDBas6OPrV7lmhi/z89dveoHs8qum+CN5iM6VC9i6YbhnlgKffg
JNveum0uAKqyqN3kgvxkHjav/OUxE2gvd8EJBi3EzJCMyH8CHbL5U1RvKzjyF5z1
3uVFfKpqW91HAycDel20zpKwqYDKBAeSWyz/x6yUVCpY+xb3HXXOg4ImxLy0EKfG
SoCfTcSR/t5tG0W3tEylz9Fnw9+5p6aBzszm52bhCbiPhF+GsrYVtMSZvCbKlUqI
Nre9MXmiLZyKHH+ZmplDx/8TwzTjrC3Dlpby6pDlM3rXJ6n620hwy88lRiYzW27W
7G5IXSpezCaAJBrhgZq8YqDCmGSAivcEcao8EnNjjbAecS5oXLZfNpGjmIrcgdqv
aXHfOr+yUkprZj+bAYWOFYgoRyY40Dbyixc8LkbNrDktqsbbn0sR7UhUac6DVMwi
zj48vq1ep49bXFk2gDCWmzRIlAkhn6lNvJiGIu5vjleqn3RpC8OXFwf1Wq1p2b45
q/oT6f2wk1zoCF29PXxAELqwziMDN3X42xXVknu6QCYWKq2Uyi2hxxSDhW16Rx49
yNB9ngeHEIL7kkpWL3vuiQZ8uiiALpIkXtZDqNbUPnrz6E8k54TE81DHcxgYJaCI
DKcsjd5N8Lxg2UDJKOv6C4XDu9OTseJzyXiTcLSdARkzrNmVipHXvV/GkPIq87y3
GOAUBjEyT55v49a+PFFC5uw9GW1299CfN8Xksv0fJXn4fqrXX23OYo9VaaUeWtyI
l56cEmSXeIaJ5u4y2HQBdCjUwAR9zJyhwkUjZz84Hueg8N6AqVF6uqvHfC0h0R1O
sPm8fhJa5XUyci74SWcJskyLoYe6RRuTXEHNrrMhy3optnksTCLjCS6axbymh3ZF
Bfq+7iv4IECdWErs0rqlwFMCRsf0Yna7IgVrJwK0G8TnJfDxMMybJXi1ZjNkfWYU
Qmvh/Q1A572nYZtjrl8ASm5JW0GL2BY2i3eWBMbJGzE4EXmRPh8gxRQV/e7EYxw/
j1iWML/LBbicXCmYYL+Isxry/CTiJO20vyAGjlGXqQOiWHFBwNyiFTrMtA4uSMNK
4v34nUfBmgsAeSumT+ZegX5fvF4rFgEqSNiZpvyUjCqY1il77fKDCwSpVsH/EewK
2UXPGivTud56BUl9dMa+8VHc6HtBC1cQGiGGcqGDgnLKpc1GuxlXQbCoX1S9ICli
LxnW2mnjTxHryGSivFISTlfoOQDCKyKcRfM7qBHSX8525+zou/uawzAzkCUXIF4u
D5BfGxT/uaVoef4Pltc9tLIlxf4WMwO6q6gqlNjm6xAsYMeSmGOzDl3YqgggdR7v
fnce4HFHwrVgozf79iz6hxX4cHvNQGUOAX+91XaaIM9IwXlUy0oZUjS9Kf4saq19
iwSap9ZCqS5EjPhSr2IJVTPSdiMxMFOCt2uK/LwWcnsx1ptLPSYE9fqklW0oNHHB
vhYzzoE+07fm2e3A/zbOGolgzm2xgnrIqcp3iBbm4Bjzxsj9GBkn4Tk8TTdSo9Sy
4PZsVGO6gKVROvS3rFOKvEwZUVCG+IwL2w1Ps4YvqKlOczi4Yg9oHpZrRS+jjJut
ajSNkB26hmDW5osk/6PSDaT6OnGOxw4RFBRfbPhS9sNEGuS1mkBA7K3RMMrbuf1I
ziQwXdILrdtY1uhl8EEpz9se5d8cRLedscGTwfY+D6vrAZPFmfQKwiIWAQK99t5Q
kRikhz6zgMzyzy+A9QEUcOPY/eU4V1399CTw267DgrtehW6PQgeBmFvvRRt/Nmig
b4Kg9j5q4ECI8XMyzWnYfSpRpRra3pLeYo8MCcB+gRZC5IbC7Idk+TV9O9VLkqmr
dC6UPWGM+5UEGTfQOStWreoMU3INfRz8Tbhbimn+hcqEPA/g6IlmRFt6IUeJYSO0
Z+zIy87rjB4qvcwTtcsaJJFh1IaUYxwfzDSzPfAGb6IAOCIuPJZ3lP9pUBHVErKL
LbAe7XNzYcal0+y+U8QxOcL0J0V5s0aSsOk7W0SZjmF0Z0CIaoRbyqQGDE2FZIsg
Q17del9/JrEbRT10s6lmQaiwa/v2NJ9Ow1YmJ4YSWgGmDGPFwKntQLZZIFljZtUO
ptB6RrXdkxseTmP+nBy/b1aTG07LCx0F1C6LKQweTDImTq99fymlO3rZ0M4ksCPV
EpXpYkZJUBWGQv5bWcKeT1mP2LzGy5A6Kkgvp+sdCy/XEjzQlgn2WHoXeaKHbxh4
GbXsmDpajdFarQxXiI46W4e8nNXU9jrh92jnhxaPOd5daCVPKnEoy/pIbdSQN68M
87RyRkk89iDuRBLolcF0zZRHqYl8zbUUCRrliAj9ZfqsFyxikmJWZRfO7VqZ7+3k
+noLDnELX0TuVMIe8SCfIQEHQLLYWe8hsx+t+hMEpoSGOpBwYZMia7SI0e9NxdX6
qJJuS3Vb2sT1/jvnRTkz2DWpljY55V54HNoLiIjtlnTNwkbRoPeB1SRdr+UyKNHL
TlLmWTvf6X9yjAEw8oXOWuTQLUFjwAoL3Y7GuPZ2cPFI+1Py+NKe2Wr9PsiqL/dY
0lv0w15h+VR5S4AnJB7TaOgYhrFa2MWXJ2nQbDzvLYz6vLBwC8C4eGSuNpqHl+c4
8up8xR9b6v/6T80YWuHrnmrP6PKEC+w2w2hUmCs/GAMFiiyx37DLm2K2qmnPtJWa
T0dCOs6hrNWJISJDtbDqh/gjJ7RJjWB4OcVE7vE5TnTO7YmFw3sWooMzGcAdXXiK
ZvpSVdHmdVYThaJN1XY8ESYYCPsL3wNN0+ezeqgcBV7a6/VuS3hdc49Ram7QNP+k
aPyIYyZ8BCnFDV2lyreHPAD7i6asdb/wGk3HqMBpnjzSWDLyG6d+b5SWDjHQb/LB
qYi5cpCqMsyGBj2ROKc+Js0V/nWAUI9WlH1qFJNPACpJbaNFclIq0a7dS+/SF/Fh
yz93pv3gLGnfxkEhhRCDJOiIfOgH5u9yrjUwKkEahPl0+lM9+Fzdsri0qXZMroLe
O8avZ/zz2QcDqBEZh7DV6WcTNfdU6VvR7UMz/HdAYE7h4I6rqtGa+LB+tuND2fUr
PD2mOJw2lb+P00toZW9H98WtGHHp5Vi5iWVkjhUGShWKBgpmVDggfkBOOpTctpB4
F/rO+EODCWeUGQfLEPfBBvIsUCg/9ZNGqzb4ffGpa7/NYvJUg+Nnwc7iaxu4E8W/
szzsGC/AFME7tRN9E52QwRlX3d2Ge4aQSirXQ6qgUakqHNGX5Wtn8xVRksvENZXf
RjUGWcWIMtCsvxNLdorCl3WRjf5jVu67ux7kSFIhxx7Oy+L81fyp9NdLqnyiyz4t
nqCzB/XlkD+6vNpjqWbhmTv6vQo5W1Nf9EGtcvfvec0mzmTD7m2J+zUPOnpfps0G
u5W5ZdfjwXsBjG4cbx7pbtW9qyjMjvqcHCLCReTK8T07u8ByCzVH/pntkYbTnNUB
1khaqdWQobqBI+6n8ltj7M+bbUjYV1ffdH3BFQKnwREi4PUacZvm1SkyWGgqlxDF
2oxt4xg08U0HGbjAf88j0Ld/pCQc0sLqNBCDq6LipOeLAdoBXFbbbcvvhLdb6qtX
Es7YjJ49XVuwZYj9j3BKIvG7nIboIi7p9u7f+Kbd9oBNa30yQAZGbstUGWCpZzzr
qq0cPtB7UW8A8ZF7o5oVOZ6MoWoDOYwsjpyjlRRr6eSo2FpQBywDng0GdjaWuFiL
JxiaEJTksfryh0OKnTJ0Vu4mfyxt1YurQwW3F6zyJazTfckTq9txRqCJSYQtV9CO
HgGmR/mrMMJhuAVof5No/6CDsztqxaCiI5iORatitb74uuJ/EHFDUq1RzuXGk6OU
T2EtwmFty9Y47fkjhXrsft4lMC8VKOu5dLrJSzh7L2DodGWFY3hMjGQDr3M9WK/y
a195YEqk11llFZb6N5eUYWLrJPgH5fDChKSYOGSWar58fkayjX3nBIHekflXKyVg
JsqY9u1igXc1OeGDV+9qjvtwLcvMbkMy9RDs1FKQ64AD1uZ1A4jBr+3xJ08efuou
YTnYnVmqUgATsEWXvoE24ceiADu1jVOExmXE0WXdkla703iSqb4FPdYNX44/s9HR
pDCIP+BO2xFr1zbhxQLe2tfffiGWTgCyJVmWeFRhnBXAO3pV+ZDaekj2ZdSkjCIX
qh+BxjRbm8U1dHEbdGQRAXwkZl3aBd/G52cY/oQomxJK7x4d7B0c+3K2//CpvBgk
Oimmj9ncrGHZk1vemoo/xHjO2kzMN8vQwBxy+PxGi4j8xZZngDWyD5nerTewLBiU
+Sw9SxShnd116mUnMI1aVp+Ma0R+e3WxQfM3fDK1Bwdfh3hxOAkSI7QTh30vRYO+
BDljTIESb2rCTZ/l1mqxXsf3YYRxVwq3qtTdAtZL7e2XCnPiO1tXcuGXyUqJAG8f
Y6E1Cl9Z0NsE95yyV8HVUH8toA1wkJffj9++9UghOlnlD50//UYPRHU+otNUXM+r
LXUdBQxwNlNW3BLUjiSI/x9WvsOXE25XENDX68JNb3WIxChRu7ZUPGSoJ3NTox6G
ldajVrNh2CXXgDvbSwpLA3BwHkwiL3yqDZcPHHjk/k5Edj6d3TP81WKb9WnVTpin
8k7eOPC5YNAzcrKjFhmB3SehLgCivy9VKy4EalRC95U7hegkGCitPqfAWfqZ8oIS
tThhkmAsOG7JBqUIuZ//z+q8RdpIss4HuDHpNm7NM2df/Z46MslGK+YpwyW4+Mxv
Y/a6qprwbnWAUJVPa31xC6Stsh7iGte14alb4UCO1LffSegQrWq+ZbBg/bZ78fhh
jr0iTWrJ2iUvGcbjpj4llx7RaWIgJZ/G3BHUE6SgjnAiNfHFBFfLwBM637YL3Byk
i2NiILKXQahv2zNPoLh6x1vM8G+Tm8zEGsLuCzJuPYFOyJ68rJgYrdypbKUBb1bB
ZaMjimJZwNwWhnJkJceVov+B4yzLfoMEDZWH6xI7T1qm1fmWf6zg9Tv3qmsryf64
IZ1ZrwE52FKw6MAkyNpQBbcvbt/HCVhOQPBTN/tgedJpeteaGvdSqrsLEmPLsaG7
Cg7V6ZWRzlEFERXwKdJTReTEnF+ISy4W+u+XCH8Gvukc82LVfH8agH8GGKF2Icx7
RAgjLdyWx2wNBty+wfZtN6zFQCqoX6VviwlFke1iXRbQIbzr6+BFZkq6xDYVdpm0
4NHbDtJjbnJCjzbNQ6HtCdmzyzrW1mY/VAHwnCISSBhKXkoPeqx66lWzlS6HnmlV
KibZlxq4U9fYEKP8Fu00ESndsnFkqJB6CrmVcPIBnwRjLF8L+nM72023K23EQbnV
kN2LCstFiBUDtdJx2b/hBfTAawwbneMaXppfW3/IONcbspCF6xvEiKtx00IgMuqG
d5QQxjeU5onJt6UNfKZO8YD2Y8VbnXV9S8UR4oo8sbID5mXeQ66a5JcWMhHv3UoE
hhuxlXOkT3a3DW3gZ6RcCqFs8YxMu4ndc8x8FsS6KMCrPsjJxRmdedWj75YW+5JS
tzf6J4xJONEfcdpLtScGNCSc7tb4CXjwfUbEkIyepRp5K10HpJ6KE2vpv1W7SaQT
FeO3F8W6mn3BwXCc4xVjPgVl9cMVyj+jzZbuT/GSCTFqL65Tuei8E187d5ru2ZBE
t0/uU8pUQAgbOUYc1+gLp4lu4/Z6xZe7A70j6XDYkxAUrIsMENgdG3FJMnDYn7RG
i2DClglN08qm5ERGdmY5U/2kRdB4DciX64SfNSB4z2XV64CUvvo9jqfoswu0gtDh
a/KYmdv7DoOTN56B6D+ZBBKTFmyz5Mnbagi1/7oCFoTuxpkWzYuo0Wu9916H+lDQ
yiRHc0cgCL0EJ4rfRgweTVI1tj/n9Y5Bx5CQQdJw5uIaWiYdDcEsL510NTTm+xf8
E+TB5Fln1ZRYjA5IUCRBhvi1lXpSeka7yxdWLcD1kXIbJoAJqrFaXfhuGYZTjIKG
bCDnfzMjMNbi8t4bctaBRUQsBejTc/mKm2olp5zT1FyvFO3SeD0RpCS+xH21qXQS
d9h6lUaLxK+C3D3QgjniRxanbxV7pYheUEAZd3Ww7dtxDlaft0zx1p0K5q49XdZW
vXO3VKY2uydkwPdxU4m1sKYwX7SRaOAJJotiLLieQGXBJVg+GmhGsrPdzwUxkdR5
R/mhB8L705EqrC1hbsa8Fikxe1wIesC8SPRc9ZWBwZGK7wj/1qQxDK4+mQSE/Sem
co4gjjqjd/gr4NSQgPdwJEl+ew+KL5dEsmxdyKxpXLXoMy20lvUAxl1O7nicwg0G
Y+YMyD5zS0jFOjvKgpUUxepEFUt6Yw1OvxisAYJBvnHs7YwMGNO7q0hMCfANcUWV
WkfD/rqZKRX5+Kz2E0whdtaJ2gxbmSjNPVWJFMfwh5dDTmFqdsKpaQ14FDRKtOb2
do75fDqLQjSV2Ql3lVK9rEnR0Dl/oWQZoWt6pwqkUAXHiLbbV4fS5mg9q6pm9vWr
xtoHqoYXfrKBT5aMZEzyXC3TCyjmHSdJ+1R8ArxbiwtYv7FUjYYt/V5Yu+Uqpe2R
w6Zq3dxmtoAJxYPxyquQMOsSR+Hz/1ToHs+sGdeaOGB7b0gO5/P46BJatyhyJKcE
/1B+gtflsOXEPkUG7CVrLrMgLD94vo7CIF2u2FqpNxc/522eelZn92iTnEUwk/Af
+KNyqyntYGMna1le3eCrAbGvzgeOGMrYySSlK7eGdaqqq7W319hnJmi++OSVFhlk
KhH+JC291y9L0H9PdqBF5HTX3ZGGmriftidQtjA7p15QZI3xGW9r/Y7OMkzcWZ7u
Uf6iUkjjUcTpclhz5+QnDQ+2vLA7OAB1nTMoPuk+FGKBCIS2YS1RF1pSaUcNfdaF
253xqEuUn1EGKq59Tb6Ig+vJ52Q1DJ3oYJx9OaAMfVzgYUd7yYy5jwYEDwBiyRtX
9rBRlYUAVP0+fRhE37FDme4WTmw3kXUH7OklgA8AhF2C1y+Tz4RKWQpNOcgBDCfO
20Zs/jSeS2u3hS0JS+cQaIbSd+cMGgu4X6BkNWpEKY/wk1AVcmPM17FbJCPqT1dT
zWEYeELt9nfK7K4GORglo3ne9ntQn3fUlnGIvK1GyEBwx0skoWfsusrYmqirPBC9
knbVlMxINavVkSNelK+vjWCsAKMbNw/RLQw3iQJHXjMt8wCprBv3iRzqX2Ww3KQm
Q7ClDMe4VLEeD86dM3tXX40N/ptolCJEqyRfEQGGrX3NMFt4LaOe+2In5VsQvKsS
x/J9tZITssStM62vNkUALB3hC3eD7j1NheLrEPc+6DAFC+cNzNzoJQR+K/4K771j
jv2otdB3RrJeKq7JVgyIvZE7KkGGrpfL7Hbv+JtingKizFVNuPkLe9h2Vf2JoFhm
5qh5AgD35NhLySiISvAWzDYJ6bIxH173iJML5uwAmQQQ738C59aW02kFh0RqgJwD
1GuUoYnjw2zEnPqcwvI7kw9gr5G0h3bCZw64IlMWEA1h+EQaRJ2s0CatA03SAo3h
QGCqtqO8finhy5WDI9OPs460Kd2GHF4/R2d/Sw6E4op00kyShQV0A4y2WbXk+4Y6
AUp/S40PU/fGFRgyj4EMgwiODOQJewrwnnch+8Wdg2Hcxn27Qpc+mhZjli+eoi+2
Xc5sDpDr0q0DoUZ/ci9LLbP441XVCbOPmEsNZKh8QYNQ1RKg++v8cvsc6sbpBPz2
jTK2OQuUJxUUqGMd3v8Chvc3wuqiqfvL68utad50zY1ZclpdVX+79i0+Ci38aif3
avBIzAdoB8VhCw5zOimDVHHjVjSDpkW3OSqLefRc38gfkQVYsYy9wDfpATuDt+oi
S27JVQf6Tt6gPCMI4pjVX5xW9NkO9OEWhi8y17afG6u75nYRitKfpO5UGDJMa5Pf
ofe/NqkJe/q1zC5bxAOFWN4CQ1wbYEbKZj5hPN3tB1Iq+/VvPLh4zn0pOLdggife
sv5lvPSzvz4EDMy2ILzsbPAJUVZlJXjeXvmznXfd+1/C6Vp2fxLcMMVUNy8gpwFf
MEbtjlgVHlTdCCfNY7zMNFcauivh04/WcfYLNfa14w+9ffnfgS+Nkdx01i43xTCm
kfTm4L1Mc3vFq7IyxQfOfaEY3OjHzVULeF4te7VQwyuppN5KezB0H38SxmNgBXjo
ku7s/LgM4kEsvOPkR1e+n4I9C0Oiwd7x9nDw7CWuH9+LG+uLg6h9gnjw6QfHLZW1
GUOGDQfF/3W0EBnQ1q+rywLYRUkMtnmazFi0BqLIdNfEd4k/pbXFp8NnMOQRQj6b
CayHbdHo5G6a/XScosH2WDlb4/+LubyP19S+YWtiQP0AAR7qcFqQoWYOyEzgcztx
jtlNX3YE0qP4ycf0vYMi8+7NVFEtv5cvO4cMy5Xxtc4ZNioLbkaT1Gl58brnMXmt
pJtlMWi2Hnxa0gmf/iF9C+ekSK9AZB+CDg5VqlRSZ4LUGL1hYMKJvWZe6MKIngTl
RkYIVIq4r9ihUfY7afIS9YW5g6iZ0sRCzO7wJb/4qRKdI5km/w5bmUKPyY/7YGCh
tnuv7sqVUEQS6K6U/jHKdMEdbTEY/1Y54xQAK137HjXUIbI1DaBxiCqgUzlvSQad
bXut1LAx2Jg8uPINALA3LWajAS7vViR9CYhGV/Q0GbqCDMlvVj5mIGI5u8JoFsRi
D5QBAb8dnVEoF9hdz9Yyayl7OOzZyP4ZxqSCMsmHrDSq0R6fIs6LHtp3kHcYTbmx
CjTtiB6pAcuxjF/ctfpl+O67VWgEnt//cUYJL3BT2qaCuea4tQfIqGNZ5CC1FW77
vkYB20S2eiUJnk3ksJnlvRQyOnG5hR1cVl+9FZbZnCV08OOwzaz395JjpehlsKgw
7q7tbbB6spV8Sjqo6kXj5zO2jrnDtG7MP/BR6Fmld086iniWnwPi2drZyWZsas6l
BviO5cNJHaUhqtEG0fUQV+VrrDhK3Fwf128xfXHSf7sDA4HMpK8LVHNcniJcZrHZ
rIfE5UqaKuVDHxob7rW1cddBcRcq3OEXIFOiFIadkeEflkifkJ2avhQ9gsfpyquO
C/+g0x+Ss3XMVjRclgPUDvXpBl6kMtSalDh3eTMAm1wIwt6bGKKcGdI7xM4J/vER
ZZgRqlwKyegOlTVCXebWsJ0EfTZK4kIuvn25T1j086AVYothoVapGQdQHRvFSGs/
KFfv3kenhc9FJJE0SBTZG1oUrFzdB1KmRQQAwZH8Vry4TkyQ9YPgzQrij+kdXiN+
mWRuTeBfEr0/yU2OlHMXjQm9nj0IvvhUh/XvA7kBc2q9ivkT+3Lu/QDHo5PJi96a
/nwoXPIXHz/8p2rI1deL6X6gsYDJL3W90QINdkPGMA323YoQd91VffuMG4e7YtUM
vGrfWGdJ9BlL1We1bSn2vI+HGGhpVPMEA22s+QlblkZ4TAhfD9WlKjB3HVave9lj
eXLLw2zl+KIEk736B70B8g9UK15PkV9JvruiHnvglwkP8qDERKnyIh6bX9sQ2Gw4
weMbF3F96gD15UjxObMGKxqnbhk/D5eUFtW2LitBd+47n+7jueWKp/ABfwZ7Q7op
D3+oZfoJoV6xjWH3g90Iyol+Amx12piuvnKuAXSQoRHJ+mkdpBFaFCMn9bHan68Q
O1aKfrSerbcWkKZYxZKtBD9uwqWf38EYufVQPS/b3mmBUrVkAfxZguJb/0x7KelV
XmXJ4TbsjhN0QP/am0c41xiFRtqLfnIRuFMdK5CD86DGrdpaeCSVy6nABfiixsPX
sduJSD2PU0B5qBWkEgxZVC81WuiMaN2Vw7K+OnooNP2ECttgkIkaBaFb/4dMIR2g
0H7MVqpgQOQukcUydGz7Im+ROkaa7LbT8EaDaQg9aE4BY8CLN173KZfA2D/AUA0U
yzK5tbOabU9bydy0dKxYK3+kAwxRX3GKF9FJYtgPZPGmyNjs2kF6YSn4QxUXSbBw
B9WbKy1cB4w2TbV3k873vgu2sacutd/XwfTpmJ5/5nxYNtp4jRgqteneXczAnJ8g
H0RSp0mmdGYJoPmi6VS1zSFX7+ONUk1OEhYllcEZzdewE5j2oyOgatn6l4m8B64p
u1w72aGovQesFgjQPqP5/4OXhgQ6pReRc6w2MgONEFwcsbi480qnp/h23NDmigHP
EVu/8hLUkNrDN4oa2YGIqKOq19zOBZwIjv/ebSjeIAi2mgtmY58Q9GaFQCPnpotS
Qy7J6r43Y/FHo6lqs0riqbhLg0O/r0H7o86Qw4TUt4GhyPusH05WeZNf3cokd1u8
Db7pVZGaqRQlMklip5mmYD+vNEQnngozdIAbiSTkBEMn6dWdAyV/b6bCD2M5UWeb
Yhcd6H5f8eufvaIOkyHGz6vi5MIG7LbSlkQnQuySQInhusfJrWwikjl4IKyrdZdV
FMeOdxKPEcUUiqcDKpqM02e1/Eps6bAjop/+QgrQ+qOj5njsSI6iiTzj7mCDveOj
y6uf6mg0+kZ10HrrdIErl3QBZ+uX5upcw17Y77m4rHFgzGo5LZKubsijZH3H9Fop
4ZQ/fHerkVr9F81AepksDjdddL7KDjFnPfY1tq4519kLSG0qDFvwFFJSbSNaIeA7
pPC3qD3LKZ1tTBGdNVtZ2Bd0dc39QRTpxAykEpNAJAfIovx0BF4RHkXgctx9SPaG
DHGMDXuPqAvNf2KZgPoK4i++V/FRpADD4RfBy0EWPZaoPoYGrdhcERWnBp3/Rtcx
jevRvwjnD/FYOWEHXAcPQ8svNbhKIhxXdKYmH8MkSJztP45dAuvfppqu16lstHrP
hjTClm5AfzHtCM1YgvEK0Q9xuDwfPpegcCJw78iVHXout45SoXnnXpec2Sc6Ipls
x0Dm04dNJW7qfKehDzhuqbWPr0PR6oUoYFkHj1B3YTDHoclTOttL8Xqcz6uO25PJ
mNUOB8V1/FSsilEqMqVRhCQU3g6BLS4OMseeOlUHKFLp4O24pVJhZJVYOSnfgPC2
5sYZPnv4DgwPqJIDtaC4w+1ZbiBQnzROMBDUy+7FxI00TPllmBx5339fW+ryBreo
xW+RXdWuttjGh++XHxbL2rwPtjkBezAOoAdYrVQAZvAyyfgSivSlhicr0JFLvHXP
ckkq4vnmt5vBhl3oL1PXxRlVPysE5seOADcYlPCimpGeXP9XsFfq+V9TDQBBO10j
AXsYAvBYRAqJU3YAI0xRPZyWe+KiMPw4KHb7BJ2v5yNVhFfZBFNx+WeZps5M6a6a
5FdgBnQM7IUERNRDds1zo5x/PEUpuJjYAQRoJzHbRiKSTScAQXNCSTr7L9T3gdZS
p3yLMc4ib00tuqx7YU3Nb7TzklLUcD3wFSUO+sZzcaoeAm0m1xoVp8gw4WuKjFWw
uNYeQW9a1vSJhG2yr6EvfM3G3jWfSxtRptdHVyFUz4tPnEzHqJ873VU55lcp3mAX
urn4uD3HPm/1QHMw4676e+0Vr2UHjNSZXQSmJ4yJ0HLO9ruk1JW7UvSjXHELlA9p
pKxPn4+w/4+cqvpbNvtZGMlqKwAVVBtcXB/Y8lWjODa1uIoP/75cvhaUpWRbRnJG
By6XPIxvYmB+DzCYgDucscyit/8fyDgwFMMBUV+dqCPNqq58P1kmKuu9uETK4iJT
cIelXXfBhe1Ps+hX8/W7XG0bjbSPkYbTBvR4/017Ek4SraDpVm2jV/SCQaFPYgHd
k7bxTkGp5DzVqD3ULJt4xoChIaFCNhGoTdkhDG/S+FA49V8SlqKb5th8nDgaEWqo
lQvfRhhRolZY2GnB4on7U/SMHzDVw2TNb5Fmpw+g+76hol3XJarrxAkSV1UnZUTi
yGCZj8lIGK5+WIzUcW+ZoTtw8P4WN0ICVi12Tim9abJ46NNl3o2xPvimFuDqGyVh
d9RvtkWKQ4AyuP4Br0kFfdrXm4xSBox57b0aYWtw5iMtlX7JRLTY1j+8q4o4zilg
zw1f2w1P80gDEJc07oQj8EfbNmb2lNnIHW7HrJ9a1rIbzBVmfEs3IF1zG4IxXbBi
/x+DO4dVrNkQUkh36f0NlNtlzaLjD7gV/RjJVyagqITiclYOddjWoZXHqjD+gzeZ
5mxotdE8RhEGbqrOt2Rk/9NU8nYXB1P/DFP57YyKJgM02EhFowzJmFwjZ2jOJL5K
pjf3PQvWGKNlk2L1HHLjqLSeIr9i55J9vfxUg/QzjM9WJ1dUR7r/YTz7dvyLpOHC
/maDTQh9MQ4QOntf9RIML1zuUWAEyuaY3t3ftRKQTz/9R+B44ni6o1OhjmqS1AA+
AvzSm/TAfkFQZsPG0LME5YiGb9tN2BB91pntVF+PcYmpoGMAN+2TjPcBptPT+gFq
9zOKuyHwv1JdPgbZcAQ3S2JqkGjyi9nrT/ZsUY4th/viQKyzhrXG8yYZgF4Nk/TB
IP2cd6iyrGHTCabzR58BCwy0W+84PcrQtd/05NLnMYahH7UQtTGb0f3mm8+Kb0Rn
35n1MHr0i1gwU+yTCUFKar3A0dWXRPtCJQaxA/i8gp28HSV+X1m1zSH4WWj2+aLm
NbV51qVlphzWsxJKYWxmxZ5uPqjq+b5Py3zxyAZN4h7HMbTE71E4Yk8jBz4kJRjZ
pAC0IDFPiFGmLSkl4dqC/LTEXbc6O8d+9bYpyHNVEC1Tx48OQpwL4oPeVscdifUL
exiLzlayDy4GUELD0fB4I5InCev/zVKzPCj1uxcDeurY1poEPUejgu36I6NtEFBk
jronNrP+6mBAr8rzwC2hh0eU1kYNnd5gYgkfRdBKrGWUT4etiiZYEOM65TdmF1nH
s45JhLp/vPPjYUFJDhO769l2tjaA8WAWH/LwLOc1M/fVgsLQMbMuY8RMs8j306nU
iIm3ENby7ezFHSCpjzDMsG8Hx9RpZYvhzBshROyT8c1xAzJAjFMNrP4i5gSGTW/L
LHB/0T5wCGJ+uvAmkGUV1WO5cYt0RbIoGxbNUGloT1/qGTGKJkDU6qTUnJLSs+yp
b1N3BFtf86ZX9kSTPa73KcMtzlijah5/bQVbrPLCA+479fFWoS2CudNCky513+vl
tuGDCpWfDbNGjxeozOzU33sUBRTJAnd2jFool4sC76jJnG3o1fe2vHOvJ+a9cEgR
nSTMHICfCbCb3kftN4JRvL7Z6fyDS3v1Dyh3BPNwTd2WCmTpYDjsjfowfGzjjJPR
nBma9jPY3hYvgVjXBSlEjKkZ7P3a+BhBac8ERxMFBNbhlAg3c8N9Gj6FyAic+9/Q
JPcXBgwCHq/PcEpFkOArRI9/jfEw/KynQpoa/CwMq3YCvtD2AUgNefE3HBIcXqQG
6nAI3A9K/gL6g9C2Dn7RvL8KrSNqYIM9/sauPTGGs7mMTibnjVnHGb3KDuD7picT
8Eu7EqEfN7eTQtWomWkITjU5ipV6o63SYO3ZHHe6JPL19pcac+kell9i5OQsjrUS
gC81efYjOmBXNpYmkTUGZEDxzT+SFOS6N9m5mEr3kbG7oMrHIw9vvTpB95nmpTLq
dqeu3cmgkpkITopiKmUqBlettv+XgZDycRvXGpFpNwQinyNKRVArR/0OhVXYbDm7
IxXiGxrnY05gQFCnZLH9PR/+y0jGaCQfMinBK9C1Ck3qjgXW4VMc8OQDTuOCg57T
P6nnoBbDQVG02UebBjJ49YkpetD9VyWOAHyItRkSyj2fJXU6vaO1qpWRzXSyIKNg
0xTIuga1+B0cA6OfVgaJ4ODa/CrRF4kx3TmT7DQYLMN+Ci4g2uFBMmsbXjaUl39c
vGhfszWQLMT79rOShm+S+J50xv+ZuYWVIh/TPx9OSfCamexc0Ub9/QGdSWz2gYqg
ymcN99JSGrKBsm0zswsKuUz7wxiyvcO6ov7c87iuS2OvHOolgsJSixegxd9BB+Ne
sjgP9AYXFafVMurVU26BD9SqgG8UdSlpCa6ZUv8YNwC5S3bxuifvBe+PyBIe6r1S
axTUkBR9Q9D3LRzuVOSxo/ukZjTHdQfv+NmsWizCf9t7zi9odeQF0RFE/dp9xpmh
tZN7g4jHTU/xpYMzD1RLhfYmO8x9xEcItFDMqOe06EQRE9D++vE0zFkt/cUKZI/A
rEHHkJig8vAzNNJENGBXd0Oer95iD709nz0H5HysNauajUD2V+MnwOHtsXbLzUdy
RMcwkEAZBE0c8FtovTj6CGQWulgY66ZLC78rJHW2hscEoCVxunefF9nZrhJeCplL
H++pUklRC6WGb0KQfjMEuDz0nZyLm4Ds1QY5UeFh0j4PfMQA4Eneu4a7lbZLPdWJ
OKNAFsMN08KDIORpEW9LSv3yw2F6WyGcT+kJtWDH78GqBnnw0nlsiiyr5sMTs+h6
Ufw3RqiFyGPxTdR/5USG/y3Db7Mygr3BhAtaLMPM9rzZeu0p29eBv64JWnu2TkRU
i2A+0LzU/ynkvuld0d0TSIAHYKaXri0Csb/jvPtLlWdrRdyOd6gEZ1Abi1mJwqNR
znVfTdjC3C0Xe1N1o0yPWT/bE0v4rlnVfEkAklqXMSU2YHTaND5E2QBsKmKxspQq
WChWDoUPuZddG8lDjJQCkXKIuDSGr52LiASNw8POT4Z4OP9Xtv1cJgdHWZo4C3YR
8Xt84xRBk7sWm/15sU32eaHyhGA4iSK+R7aClL6wL94iZhB1fGutCVSRl3AbGuau
69zJpTzR3RTcfnCwB0hqKIV+U9CQ3KY337yIiRZEjnvutaaaSUhiIhu8GlhT7F1C
Sh+Ax10OX6QdYDYDuzcQ+3fPlSZHDVBIyQSslnpqEuOXgbKz7Fsyh9zz5VU+Uz5z
blUoslVwfgOY9fZSHKh2oVeL4l0XLhyZkBL/5Rs2UACJoDDdKqqiLuLZiFwE/NhG
ytUQlBOE2LK0fIdPx+pOzrMRL+t6uqBwmAaXky7A+4A/Eh+BTNEQ7yqaVj++A5tq
MPmUE5qw7F431FspGuCk+mCF9TzrzKt0mO3D2nHs0LqvufRRWPB7iOJsYtEoOad1
v+BHD0fybBDfnumuBbpuCsMIS9Y+rd/JCt95S0Qss4374PYn3MepsUykWbUNO2yz
9D3TdgfkQY3BMzlAZsOagAuyCyE4wBqqv0ctlittIx5a7i8uBrc8RLcCyvTsRYvf
1lYIQzDqis2iTLGJ6irJrKo5/wfAZ9TDdXlqG68LzGIhmsF7yy8FJeLVdipwulvR
eao7be8z0gIKvUPHDKYJJaXpH/6fwqUzScEcay84LsD2IiRbmrumubOnToHiUYGI
Kygbf1UwrtKvIImH2uLm8fDhBsEYs1SyWTo9aUSXDKajYaparthRGop2L77Gqcg1
pALRki3nAtp0p61CfIWr540tuGRXUPNVq7Tp7e4PAEh8EfpRQvx0fhZN4EH2BBuP
kBO184RLTh0cJGOSkJ2nSyxRNlqEgGD4WHhIINb2dJ4otQrmlHgUS6mZ75yXgPJT
+dW9SozlNCP94vsmnmQp5UI8slPL+xnKkejifB0+arxZczWRfkzkpulg+cHimcqh
VEZnQGtsq9sR2TxeCBvB2SDNvKLFwu/PjzYe3pVSWo8Db9kEFLdoudfSDGRHYQMP
ic90eEq+WbjS/aHM5FODuLlbdr+zUtnIX82huXSrTD7u1iXX+BvZpndd/TFNIao1
oBoOuTh+nC3WCjBKSdh9UArnm5YHLPR3cXgJHHT5Fgy5J41IkzNyZ2C7xG/subkZ
WKN2WYEcbwmmsgYFXJHo/0D3xQb/6+d1aQusQBLRVJzRnocMyoqwyzMeSY8/qYZr
7EWW/smVil/hSKT2Wa+Xf/DpPKdqBfbOp7QQuUDUD0Cj2++jF8dI1guSv3yhbCPJ
LxCT0adNDUTGMAxIJDWYjwPeL7MDdNZbAGE3rmFEXRfeOyxmoyTYiN5rxVihauN5
d+I2nXfPG1lUmfJwfV54JvqLNRIomwaAz+w3EMFaayjQejy4oM65eW6C5LXI8SMW
1bQEgYNvXB1oNLDusmtYK/ndkvu/n4ZlY8s2HabA+I2pgF4q4dKTgX/+3ozfji5r
k+wVKMU5lzbbk8DLZWUKGVnXAlhDeI6TWjoT9hnPDxHR86IAn/6OcmSgcy1FlXgw
wPTXRNnzUNCkJqczM2YtdFd/aMKEc/s+flYPsbdglH6AMABMKZLbnNb828MGZSkO
2SPKmusXmUhiH6yF5lxhE2l5QWmU4vRNQWMzb3vWt7NzynwXqEYz3bvS5Dg4qTD1
Gou+f3zAS0cG5HO31yLj/tkkyy/ySOfyjiN0mRat5JJpzWghWLTFRsDtsrybWT7K
JzgeEJTfEkoOXK00oicISCKQFp0hfYr71Y3tj3W7DdLlYE5r40b+Hh1r+9dKQvs4
jze6vooVNoEvObtV4CvliF+w03ZMC1BsETWDxLVWjc4Yu2wEasQE+/dKqyFKNKCZ
hkrn1WXIV2w2OUVBh+XSpruVAEq+I5M9vKuLURAmTZ/tXYsUsf5ltCYBCrDAxYwB
FYFocO9Rj/YuWlYmEtVskX7QFhCvC9YeMoaGUeGzU43BrC1wxuZF+F4jmILY4Cen
lHSHgRkAU3ezZhaGCqMKH4QW5o2tC4Tb4EFjgZP2dy0nzgGrsFzWixKfDoZm9oB3
qlKSyVr5AQJAGmQgkD6FRvBX2auoKjtbDxhksKZLK4JGwM0qvmTaAvb7s1sHRR5M
XSoq6VMEDuFbHsxEr+gAhqUfX4s+3kWYzn6LxkYHlz8Ew/8dD6pdsHvHaiuPK16Y
NL6RJ7Ec6b+SK5pb2M3RPAM0ZVSs7HqjbuoX2bbJkOR/IlO/L37abfTueA3GZFDn
MKbUuO7LlXsVuAk9POOz0i7chTykPUdJKBG+hM996MEYkWRuppEFB7rt8GsvOXbh
yiwMi9ywXIBJYXm7Xq2aHybKFGWzpqrsyM34GXbUZe5gUNwpbV+0baPi7CxbBjHF
Kb489dFcdqABaZHcFwISEj48Zu8hw83nLS2HmDNuY8Mamm35oaIVxuk836tFasb7
IcjPsY1F7NDienK5sTrqIv60S6P4xrVzMeJC0DM4bu2n6fygf6lJzo0ckGhlCh3T
rNbxO82T/zB9YEwxpDQ7uMtIvJkoagnkwh+2EmMyvJjj8BhV1zjQtEZ+w4Tu0rSU
BteF0iuvBGXHy4C3RgH7+dJ0JiTMT5cKkpMbmoLKN5vATM9jBh5gf7AkY8mKAl38
Q1+ppKl1qbcYjRDNw6od1FyDREkcmsvKPPQKwoyV7qAs21/l8m0oBbFHlFlBDF5t
6M61Ag9zcVuf7QZkPWAL6F8UlfImuOTmKbJNlGJ9kbq0l6TglMXX2kRJJ5EFr8lf
fyNhjlrCg8Vm9C5EjrovO0h4yyGNNeslyl+bde+YL64paLuQPjkjrgNjBZsMYIwK
8uKkrXu0breOej5iImA5WPojMzluQPte0FjdFBOjxk9LYIm1JVhzTm8oxNNdKp0O
PFvBHem6iDCHRRLjlX61I2Wz3XCYoFZiIBtN+h0DmEM5wYl61zFXnA6cTxxT0c0Q
uhVQ9jQNUG8nYRoMHdZ8GHtq63eLInnDdf3orY0bCnnyDEIvACglh6POC3x9B7fk
eUzKwXxbh/yfWUQ/pWETaDtfQD500ypw9BsrjDX+CNtn5hr/1o97UnSgCkEagOOS
HOgjV58w4/eJzDljFOoC65rCl6VJgBM3EkefXhLxGmLZPBtkoZ57atkh6LibjRdo
8aBBNpTlHQDX8tSSQidFtijh5CtqDdPHr+vrO2v32AgnXrsbyqi1nzm9ErJ0e1H3
Ns2lSnyWQVGc+i0cxnv0/70osVNxnXHkPgOrWXEaBtOBQMU9dHFy9UUBIlb/QPbM
emVLOV9Xu20Qy9Gsk+hXooUlpMcUvH+zaXitRsp1HQFo9qrc34gPq2G7iAkN4FAY
U7om5YJQPu8pAILxBV03wQ0qrgw0NUYnYgCp8lYX56OP0bR/noUUhAKYO6ZPjMzr
krOx7SzlQQOCNIftdX9tCQtXcpXKMFifTtOZaXUxqaQGbDO+6K+sfk6kUzcaXKb6
BJzI4tMbHQMEHAiqZmqpKf+lf5/jSWzVlWgGumgB8VXdItybE7aERBuDb355pjqA
rkc/orrhTNo2joL/MzSrnkSQqhO06LvQNTpy1kGPBFLeMj1YdW1vHvG+3ixVn/Cq
hRUBXKrguYPwGMQpre+WFqRURqpbyTi6AeK2FT4g32K4BPtsSGSXNZc+7M85qLXg
PYSqCUnvRC9msadPEMLkaxPuAnDNxKLOkU5cGYMWipmu//tbI/vihxcidejsin5w
OoN/JJxedFRz/8n8FF3LrxM/m6s5DJhxj8tMTC9aAupAqEA+NHXZHzzQHuRVzhO7
3iwv52di7LSWm8zMjpOy3A/za3gz5rmT+38XCbQT6zMgqIh9fOv8Nis33Il2qxD9
4fiO8Sv8lmDBR3cIbOF7vFPK0cfg9iZZkBrVL0JuLWTr9usvG3ONX7/VwquieQdA
FvV9dqov0j9H8KWS6ijsrRQqYp6mCAmjKksOx3w+3tdvFX85mEjCP0h7wN+RwK7L
Nd+2CiX09tS3pio4zUEBFcTPtZ4krdgh4Z0XBDu1tYsEdFohnEo3fdp+bwRpzrec
gp5IKajFS+H4K+ZPt5RzHhwuXKvaThfJlLxr9Y5G6mHMSA4S6YabceB5IVToNVf4
yFFnCFeuDmNxZaMwxht+zdq2DCOv+opscVnTPZU45pju4pq5rGxbBKR4T6sWNete
7gESFgIeiVbS8Fu+cD5uazBF8ASWzT8asgiuKP9Qs/fvaMhZWgqNV5GOg7mbZjBX
aJw78lcoewoRtaon+D4SEPOuCcFKuYFCetOLjNWAtJp7rbceGEb9up8JWyVa2nYV
fRxNtbZ5YO3f2sC1kz8/c7x867CN7+K93b0alf1p5fF0nKDQH1bLtEM0zafBjaWu
43b4a0XQZbawSJkBp34IvfW1y6FtLnfrf+BlTeyObaLvR7jQdvmLNnlnywhQoWHI
/deISkBkoUZYtj40q33HCn3H+SaJfO7aUEaFgHAwcJW7gEvPCZ657hoJSEOwKWLa
JOZASyLilqvMnLjHNCavhxlHMGURClH4Y1qp0OaCJTGJNl22/E5uSoIe9N1VGAjn
ioMKMPTU9xP+p8g3JGqFhmE7YFlbTDVFXaXeFerqJAjJ7WMnaaV52DiFcNaBePxg
lKg+uco6a9mP0dSAdA7xChtQhMnzhkFLvrCu9FLHregbqQFY3FUIZOxlDNCWK2vk
mbTKbuOBeSZ8/aUB/V8Z0laPhVfkaQlNOMXt5WnSmNLsrj+ZKLiDpFvPgyNB3P+W
LHYBzp6sgLfQ3vZuOPijwlGxwHz+1bRM4dPq17J4Re1BLLNVErXzow+UHLynLg7A
HJbuw2S2AmMuwYd9QXThQ6zZqATarn73CmGfI43+5knC0hpYDWfxoj/EpI+vxXsG
GmLn6hDYmJcfcMGH9Iv4zOblARCsQNflm4ITrKVwwBteT6HaVk14omCB2r/LW4Ai
lPsymPlbSO+tmxRgt4jHCh1bpWg5sHyo/jGnzHq+xDMTzPnbURV2KbDD7WkQTOVn
xsrx1gwuKMW12xxYxrvOyszRLWA5UmjqdYiL4MkU130OR7FMQsem0/rw+GFpTigK
0mdYenO9DlRe3si8pRssedwBvTDxJukJLwahyJVYVduHzd4CvleFGbrkY7yD3rm6
hrA/cym2/Aui0ZpSfLhz+jKlFVN9vDfAMOACSWQ/97BbwvEz+EDT4EL8lrPWxSxB
u9d2LqngnpyNRBmOF2R7nQLnjaXsmsfkOGqg2i8ztzCUJDQPMgP1oLN5rNaBtn5V
ujWBGzAwmOzQROzwlD4BPxJQPNjpvjlLRW11O74WbUw21qSTBelR0BkvrEkGoNDo
3ZJ3d8gdDN2kRW8BTtFBftRHhna58bUE2N/1u9UCrTj7r5ghQjgVkIV2NXUAIzL2
NhPBnlWmPwizLa00g5ab2g3jTT59dZdI3TeNtymA+FiV12UEaItgBQHvrL9VHE1V
8Snhwt5eg5VATOq3TKhKtH0MrLCyXLkP7jET5bDgptkHUTBnwGoqkSPVaSFNpnG1
4dCEUPOktxzvneICvM+SFBEcAOSKl7X894s1UNvayYf9QC3Q8SXd9f7IBIgC6hMx
VkHZZjijpGdAPs1Mzhs9ajemiqKXiJWnvnGpnhejA4fVq4GsxI6H2cNoOynTS9/t
9ZguA6MuXfsrY3yBKaVryiVjSEUnAA7olieg9Vh3kp8sMHkwXN+kRus/B0qGmllA
CMr6iIa4nhBkhabpAjgwwFh6B0QYd+nIAVjZE7DsFHy256Ydm4dKC9sATzpteEBz
hD3TNj7Kh4Gk7Tw892+A8Le57BntYQL3FK6Ug1EMosdBh/1x4yRARJBvvYDy1NXl
tR+tHPK0qtnTvE7liz2/iChb7qj1GiChqT5/zdnAOJaOS/81kLMu48L26MWxCeMG
F5Wl/a+cTWzTgQzCz9RcVMAH8j54/a2V7uTg5duAu4bT6D8p3wqIONbQT7U0Imak
5rmnXngf1sQF6nu2TqhpmiWLnFCccH0S7NEh4+UEYBWyDQfIxj48ogWuDKNKkBYt
cQqilhGPxD1vaGNH4FSTSe3FME8EvRAAL6WTJKWuK7YSPhjfvsQ7M57MaVOWTyAw
++607hov/xxo9OnkDXphkPoQK7e5npUpMnP3Y7JfnD/z7UmEZ6KGVHk4hc2GD0wH
NBNd1Tldvx1y0Vd3+4JfOkvu1/fn1XdK5D9iBhONP9UUEW0XyxvoQ6YHgtTeA56t
GMqoVRS+jjHxUkqCESc9ichaLMTurm9UYqK0hUD6irxIFBBBRDy925HLOgLEhmYb
zmMXgh110uvYV/tc4ZPFuAHZ56U2YPXUxcQc08UvReQFA6HtkeL8ntwEzd9/Xq6K
4YFZdqiWKbipGp81Y4t0HpCxcTlFE/7DpRKT8yK/31H6kEtuHbndR6DsBSk8rMI7
Sf9oHz8kadSP4+cOkjgfnFKmE9n7I1jHpLeR+GAv3FERDnfYlS0CDKM6Wce/rvQD
Xjst+ADwvD4v8AStIPdAonsJRkiGeFcXtkYgrOY2pGfz5eZLXDOnMcN1KVVAnlyP
209mj+FRAbK+Mu/S6vtaHL0ZMqxib0XadGIvCjhupjJEGiOPb4WhaXSXvyj55gEl
5wLdXslRL83CFuLyH2N2A8IgGeViMY6QjbPSBKTlyYKC9xYHSBkTeEsbiME6NFTE
/j0KL0D12tRTTFkzcecbWdXFoj1uQPHzu98JY+x2nkmIapOhrTa+omqUB1YDgjSF
7AamOKlsporh0M9onSdm4762Iadwj2xDBjxiYwdBVztKZdqZw06xj1l1T0BwcqGc
Jh45fFCo/osjDNSRtWmRfyoK9gsfDVVBXERqHcP9TyhtErmSPL85P9gZffTSjT5P
zOjF9/OIikOjP47lK+Np2id3qKVQeJigWkLnuCM5nBwMFqeD64CQXP336rCztlEE
C/TEIaKv6wTb+L5qCR41xJkYardVGaAsPwRAKfubb5V/f1uOYguof1/P2f8HW/aC
3Qtg299npsKrFZPu/rhfSkzSqACbY4jjJy0Jzec51zmA96LrTP7yrHZKkarw41Dm
8DtV3xHbRHDFH68ejnQBxWdYiAqo1x/mYa9OE6G0O2z4IkP+y2kTTYddorfGdPGM
JVRuIcqc4XpfuijX1LMhNhnOCmXPEkKBytMdJqdqO1881PIDb4vG7ZZR75EH2O2d
X5p2wmcXQepPAiKTd9iHuY2pAexP9/ngRyw1Rxnu4TZM802fTDJs6xtgQ4L566N7
ng2yXVQAEz+/5jJiTavioGYqGlbfbDIJzblH6b0TDj7twcdo+jLn874zpsqDWwoz
0qCCVJeBoJkPU9x7K7gmxHLg5GBuZloHq3lQByw7JusP7e3DpnLiFfWWNXCnCAAe
VElTqTFEZryBpVFSVC1q6R0Xrzoel5qE/JeJw5Ra8gOYZldd7pqnqnU7jM84XAok
JOfnkl8iI/anEquyeKGjbDEJJOeugUEZIYM/h4uel1OAW+1HEAsP5n7zmSNzamZs
6igwCROZoJqEr9msAfRUSXvEs+2Q56H6RASP843k+ypyYM8PkeyI65pFYooqXgzc
9VVNQFRLsDaAQ6cEvr6oAOqQaXIKB5UQim/BhSV7jfCOH4mlJiIwTE5FaXAuhcD1
VPfJPezemKaPNC8uNG0svToxYIB2K47bPD03fl/n7w9qGcMV6s/L9ncnMszE0y1o
af58coiRozuF+vjo2GAyuq2VUubs6SOlmVzDfz5Hz/8ulx75GaBY9v0+P/pOF0G6
ARIp+7brRjZ3dhzWiiqjOLxaUZToY8iw1qLTpbaFooAEYVRNvRNVXS7tsoMfn0Qj
fj131BghZjUp3f/BoJgZSERRLXaBHmhN0VaNvOsdJKhNQKGgUbzaF5ZdThzdskPO
jFs7703yTKoLzKOqMrMlYhbt4I8E7vWUNHtBkXyCWLv1tv3QqILRBnw3XHw2och1
39TdEXXM1q+HZz8MGn9QE75qIIhD7VEAE5Flid0msbiL293gGv58fdofU5KtO90q
TIiSGsbSRcqqy6hwpn1RdLUnKxwPUYtRNtq0hyRMKS/PJ87acRmF1CNciBlRYliZ
Sqt6JsESYYNg+lA/n9qCh0N5QUuSHga8r8COA71DOPox1qjMdb6oJEDSRwRMy3Ym
e0cVwx7tfCMsfHkDvz3r1uxgYc7KrLHfROPRDDOPdPBYkZ3eVTpoFmmCCPlwGOYC
B8NWkg4UYqYUZcV+O8wbGNiJ1Cof8S2UMjEjTFnCTDED1dn7ZOundVb3HJPhwEbp
Bem2IqkTh9VsmNWkUKibfufEu91A8HRKRaxtwQe9ElXWu8kgUWSip1+URmRE3Ro0
Buu022rfGiNcd5pgm24BYZ/WDS9cKZGw/aRIhij9VPp7wlVTke0Z0mgJ1g/RntnA
KsjJVvEyRWsyopRSL4d1rklCgJPrBmmfjRqYaP3X3oSYNkFa+hzxrb7FRhi5u53a
7bChuoPwtW3VXA2PfwfHkFfeACHZOy8+8lCsJl9GRBeXA0avha1+p13Rt/QqaFwe
ZshShgxV6zZNMeIRqV+1otUHXY/AgBn9qFoD/fpeCFqhBjd/3wSUra6p36OAU7w0
ZCBM+IKwFlvGtXMvhCE6XZukjeLYkvt+nm0qaXe9sGF/QiRgeJon3ZauzQvuLS2B
5SYlkF1vWetIOJ6Zm9BrXFsTCKm690phCb/pC1okTAWdXo5JE5bn5Vus9oZyl0dE
cFBU+b0ija/zcNwk3G7n7Y8IZuO6hP893aZvIBy7RvdhSdgkAWADqcRAR9ZOYF9p
g2nXU2Y1Drox0o5F6f8QomLLkB6qXDaxlOaJZcvWFAyt4sWd3rFF0NPYrEVdqEDF
xJuolkyjowsNA5fd9hk1s0haa5XQJGShTjog81RhnkUqj+uCWgYzpiWyexCuyuGc
e2BBC6aJbzdLjVwL7yRD1E3BxjuotpyFHBNnkooVedmu62MNcf6gsQTSnSIZZsXT
5Fgqi4KuRcx+089whdrf1ms6CJVy1iQq0o9JZ9fYJn+Es1mJIUbcPA+C7gigA3rs
FEtxgUQeOhB5RUc2PVvhqgmAdjdAS+7EQHKFYTsqRqcxic5qwh9qvCZ1Wa+ZuVTj
wSedao3PHMPDKa7lGG70qKQ4qObwjkFN8tWDBHnU2IbBbLf8VxG2s+G0oKGUFDLG
rngwWhqnDiYpey/Oh2Ndrgy3HpYggsfDCu718nUc9pYmJkMyVf/P/QmkPSmw4g4V
0s+r+TY0jWszNorBT06ukEUBxBTrCmPuupi+7+Joy1DjNPNQhw57fEofYVx082+s
DdrgR71e5UHAkZZIMl2ZSLX7uTJvDcCpgQerJyMBwtgxCZHbo+AwVpR0Oj0fZaGq
tP2vPSZK2wmJ9DWI7jtpki/Xw47tbIVqKXKjHV1ntow40Quk2ZZ+N7lwsEGX4UKL
S/TYjrYryA/yK65UqR72PKtB2zENmQUIINb4Xhw3Gk2mzC5kApcMCslO9CCAZ0ic
frAPtkvwonunobJfmW+A3kC7xE6QaHsGpVidGpDEs7kvX3kIWcRVV2c+hAOrqiet
4vVKODuNcI2QEd7SFiRFJ5hdClmi6uOjTznV1mL5r8uc5hF3PVxnJIrktp1iQ0QA
klW23SaoteftBMnT65LBDk32dZJVUSpbZ8qDridEHhwxNo59lQNeUU4/bgvw+LZT
JUFCXpWYZLQ+ycyTGbJf6DvWFB3Gw28TX2o5KGMaT/6jEA8bm1eT6hZ1Wh1X5YUf
i43zJzxI31bp2eJ2T7yGpzg0VRKa5nq75ckSRspQa4mhtQWlftPiKl5xpHkQE8WO
DuqwMWr17CEIc5NBxqkUFuC9qlhiZphKjlzhmlxULcjraKa0a95hWN6NTyQngC+S
pq92hSqGht2ZanYrpa4k3J6kUg+rVjYPXEE842D5ipIEq9u7Mqg/M7rcagIui+WU
dnTgEtDYOMaZR++MRWYg15Vq4b7CsQLtkrBwS4Pk03PRgE3wN2ddoZ5JqiaT9UkB
tjWAUEgcEdwkEBRPFZu/XEzZFxPHbMZyDHsUQUSGzSL+iStoIN/vHsQ168oHTs3p
C+Ig2OQnyMpNIbK9dz/dSX/bJ5f+i2XaXX93Z3EMIAlDxyPrVXJ+/JY8cZ+p8bQo
SX7KhrGZ+/4rOZeTCaP0LHYzO0dXY0/DTEV1nfYhtVZP2v5BqkNehFfdEzKyIUrq
OZT4FqCfOiZk4bd7d3toliZjN4ihmzv+WeLONJOi0slBV1fRskwdVqw6IkxC/trB
7To2UhRMH4r18sCECJcoChBKf5/eJOTMIg8oBSHSz0Hxtk924CUlgo4cCD+CmobO
tilM9wsDKM+tA3PvtWHOgbXBvAfdVksp/IEU16hbL+N7gON9qw08pxYgnaN4KCUP
qjFheZtBHfMam9NcDywSxM3/YIOrPonTEjSjwfh9cyp0AcPbxJN7QzRdXZcO6vtX
DwE9iklCk0CaLn8cSb1fFIPyE4iNDSIiTP+KmBwlq5s0F3xX18QlT5ds9D/Abgsz
2hXk0c1dsV1aIriTV202nWQ/z1IAsh88qRJuD11lf6eNAwjshO61q8XOIaZNe2IY
iLwwxddYExRbqPCKKSzhVmhh1v3O4xH2vYdPZtPFJbvg3IuxBtLDIikvM+IVYR6h
zi2iOILEjmkCQTUdKNwBLT7++RiA7l4MR8qhWKNZ0wBZUwp687hHkKAK/Fqg4/5Q
b4QZYCgkQ2DPZuwTK35jWW/+tQILWt02dkpHnCjNNhnYMqAvWR+8julSd51dqzJS
lajkHSZ2L8pm9bg1zaa0rg6CSykha2YJcPKcD3OMeWGY3DqgA8qA32xeTj/fCetd
ghfq4sXXOdIyl27L5px/AJnlqu6xptpjQe8nE42v1gIwaXJuc/YiIBZejzeAau07
pnE0xryqQ1OucNSXQMOb2uTgjhQrlLSNFfsZNbgmuhFXvAU2L/rWGGJNfjFqQpjD
LqsAb+FCYqvN/3wNvg6pgMktsMsU5IdaZw/6CbB6SX1eKjUz6hLO+Mie1UJNx4/r
IOsWz6WeoJnjGnO1xWzSJgMhDoYy1/VAGF81ugpb1fY5BKEwk5e70M40y6aymAZ8
tyRYtKhUt/Q64GglURSi0ruF4BgANNcd+r1BE80gulTYR9QlWTlthqNDl4I3sYb8
MIFwmA9tRxbt7+x5xfxcvWfa46AGdlHa1y8qt0q3hvCj1jD65WctMOS4vrrVe7xA
h8Ln0apuKVSXeS1UbbtyWcL619zTjQ7V2ez1GsW+6xV4P81mQ6eTBJAvDsdLBr8h
svYSFLddsVTkQ2Cbl3PXDG0Ct1wXkqI4dd+IiSDRFzZA871VNQlvdQL53WprYIT9
EdtvGD6Gsf2v968WhNPm4lO7CQUUZD7Z1SWSt+fdtaf2NTFdrt0okGSlWUpz/YKo
bX7/uQtrl8h5tPDsQyl+F5ZRysCFf2DSWw3eWX6qHFCwOMn6fYNQbo7kJhzhjBZO
WM3E9kFtgJRKyw7SaPe3dcF7ejLQLStubkU5EcTyF+ZodgeUf1Qj6tS4wLFFaA8k
Fme3cAqJkxEc4HpPZwsw/pS7gYp3QtKUY1JZA4RB0kulyRV4UQ9xmI4iqJ/KVxJE
S+L8x0CoXZuFQttI84dpgKQC8rkBOnJcqtr7PcVcdOLXtiNAI0E0LSR5crb0E3bS
ewwEHHNJlhJnoilWwBV3JEyumy1yxdaUUxEgwmu0lmJLlt9u/E9fwHHl022mF3TM
wMRGfzN9JmeJvnGa1cS76KkK+6G8tpnVEZIEQBQUZNA0+dK2X78WpdX/cFMQnfP9
xAZ9vkIl9JhS0+RNCxnxgyfNhZ49pt7acfwPM/oiGg44Pne7wSm1u3Bk0B/F8XHo
NN5++8ZoDMhRIa7B+JjOW7VGKhizIYsW4tksi9947YPLRW8+tUncB0neR7Y2jyii
LmNF2/UrrBb87fdJyxbZdZrLHO7Ufbzyk8CJ1jLBROqjjkwLgoGa0ge1hlIG25WZ
s2mA74VgcqIkRtFe7hNjCgRNSFJdCATI8A4JjcVmlXViIkvM19+I2toqMSJijaxt
boYYw3I9fa0elExmngZ6QVwDA2eglPFp0bFkZ766/BJQtNM+L7Deih3gchGH3aAe
9j8Y01tpSy4DSGRAKd68rpnyAqL+iMQLsPSfh7pj/dDhLFYbQELbGJKrsLj7dn7z
fPBdjrkcopoZTEpylurG9l3OkJB/22C+RP73lQVykraP1kyqT41JBS2wxLUb2BRC
S/oC95mGLxgN2y0tyZxMPUaB2LM9xBL7ZQxMTZ4u6XsNZXy/5LNGSHyQa3VC8uwY
Kw/blfYD4yhC/QViGjlbG60TbzSwGvpnVgDHQ0/2fkguHXQ2wE7OJyjQ2M+sQE4S
qXsI+1utpzqqKPu45nq7HJr7WnuQYOEhegj9lZ9zJEwfTmU7suYG0m1/oBjayO4Y
I30MnQ/soJtEQWiPFFkJjtV7eZfJwl9XqgwozUQtFngK11ZIjkfpl+U20fG5lx1+
HmuVhag80hbMscIzjCf/8t4tCT+YiPlieWWqRfF1qFtusxOCw3LI+UCaeeMnlJth
OrzcXHULnUS7PAzvDMqc33LtZsANS3klmKt3x9zzWwxfp8JDPsq6aPe6HGc4r0/F
FyOTs6lyhauC3jX/P63BgmriXJKXPhf4Hv2smN8YYuEkAQFZlsVS37XJEJVdj1Fw
r+8HRrd8qut3vkcLbit9R20ouubo1/RUL7GHKuIiJucaGmAu9QJAItaZ39ldulPc
XlhiHLlg6tmS+T7FHIYQyXL64T/0AY+sEzoGRlfRMMcZCyLzhoHjzjdPMH8t2wju
zyjpbY70HJygCdXt0OS3/RRjzs1zeDZTeNjI/q/nwOBMvRb/nBX4m4tG5iBOwY4Y
rijLg4FHgJ2pH3r04xxyZ/v4r8m50vniI2P9HWLwWPSlwAF9/5S2xiNBgSJbWhLv
OKQwEiCYo9bLU7cSDBoz3roidiMRgwnV4xYSmS/5xXsWkXrzvAG5nQTVHcqvZ6nq
9bdKhsDuZv1Rl+aIulUXBVlm/J5iSYJ3LhFZqLjv4D6nVsAm4dq1QVfMeSpdYnX3
+7VX9MOzE3HMGWVqr4FNO8gX7ECRkKNgrdjV9AuUnve3AtGaVk1DxgAYvKcCuJf6
klViv6Ux233BLMZpO9DFfSg5wVx3aOVVbdDyWKHMHugvKIdzdspVPlhn9cnbOW+H
wdE/vyzK3kKMWA9FWBWfA2oPQICPwNh982VqmkpORzuScdYg9PiVsLwdxvZkkowJ
bp6SA3rFL9SHl0QVIvdVfDQUOpapMu6eaVrrZHfxEIm7MneaUhJWL5mrvJkQSf3l
TDkChNzSAA8UYVKXMYRe4qkFJPInFpdx+2BMW+OhE++MCET+ctQBNceWO8pqAfsg
94Jvkg9jK/53kMOb5rYdXxayE3ns9pE3YZsfLJpDKuRK3HoQWXeUNREjbkiFeLKu
P0HoJ+bsgfpyb7Aaq7W7qpMEs7imLRZILYJpZbc/jLJlI618yxzg0UQRTNQ2CY2Z
At3MpZxPJOvQ7bFZ3pnx9s8jeopgwbw/YKZ/dHrK070ayalSx2Sm7GaBBO8umqVK
nzLu8ypKAxfd/ZN7kKUSIBmGLfy1LiYcugLtkTxn+8RyP+cH/2ltm1nNdjnIFhRN
7d7IiqNLx3ZsmEXi+nwpT0ajXdXFpnVstT1WkqcA8CW2cLcGCE0gezcbUSorDRir
zJankggqdyyseX306hgo7P70aUcdHpQvd0CrKvbbLRwNFJDrLZdl1qcTde5dFBrt
Y3qTwHZNf0Xz+k9KdEh2BMglYPLN3+7w18qqJBaAvDFTGOwV1MjRQxucfV9oLeWf
lTVIuy9YQuArIbyxOPrkwKUBwhTWbzmCQ5yIiFGQzD995eUGTQ9rdGGj0FgvHmmB
6+aZfZtmq/4lDN6qD7wo8ZUC0CqBYokDRLP9Txlid53xpqbkEKocXQH1gpDNbFku
evgif/RTv1NdtCXL6mpd+SO1T+ObkUesQuNb6b/Gkfs1sdfCyZL/B+ytl8muRV7k
ld9Fpa94edoeS9zHMzEt7flJfUvjfao3G+y/Lc4Cns0aySMCMk4OjYTWLY32fAow
j9GDK/A8D0uA5VBFXiw++VHSXmCQoi3CGbkQ6l6h4VPXkEWxzaP204aVXRu0768s
7Tk8LqLuAnQFC0tekDvN+MawGtQBtJgNrp5PpTYuJ6fvAApIZjyzpDdvfrCnyeZi
kvhvp9UGx0gV1bFij5dI59OjHvqb8OURaI9MXiz1YKoVFfQvtRB/FysIQnJq0csz
nXb9vdIN7uQwGsT41xIJoO4ly9FqfZ6BettYCiGZPPWRSOyjhHF/SKsSmV3/eBMr
WxGPT382k+hehNUQa3WxeSb7l8XwJ3KFA0jSv2Qt3I9A8vXCC32uAz16ADcudEF4
Bz49k0mdtiXKu8bGIVLOdJF0ynOgdGfb6lYlqbq6LcbGODxb9nXn+Cnk3CGc8hPd
KeblKUcqBsJyUwjzhoD40neoxByMC/M/CTvlA6ivWLildpceRpsXgsfrAO+AtXqU
WO5r6elIPM6zQA0/32B8dAcurr4LTdThV7UORzvFeflSIvexKYdjUY7oFxs53Etc
i+NQVoFsPiDoZTGwjRH5wGKXqu7tw37aENvy8OoGzL1DgJxlzr6/g0BjYKVHGMHH
6dEMuUBpsTe10aQ/asJxxRxTD+6kKxsEA4WrbW8kSMpqmI/727t3yakpY+LjNskj
/KvAqerYeK1VDkom0jFVS0uzsvOrCfoGlO2z+Dj6E5ZHjuwIpb4r1gMoib22nAZA
eguVthFzWJ4jcvK6Auttz96OctbZ4ZWdgQEfOUFU6+Jt5Bjll4QpRRjObx+c3OMb
htLj6Ldn22tfkyviv4kN3Hnjj+204i5+o/VIp1YXI/aWVjGZm13VH4kyPGqxNUNj
vnJR4lKuj5dmMgKASK60k2nCOBcvzvnFBZHauBRgU9rL3TJtfUVGSB8yXwuZ3Ywd
WRIxuuPFt7EdQ/zgR36UTjpNV73fEpGMrjgNjsSy2n22Tov0WZGs87vgYu/tkEuU
ChtCRgc13efJUEGPXdBPuZf8GQej/NOcH8UL0qB8WOyqyyUFp2WsdxDIjlqtLj1J
uLCV6iYnLJw2NIaaxuuRJdpxCGQhFYiQuLFCxelyPM3TuioCqxu+xBj6zJQeEL2j
AjuTUtKNvvqfRXJIhH9mQnUfGWmOCtyU0v2EJO5s1ApHf1ujRtPsMO+iIunB0UR+
25GzAsoRrVmvsqRA0xrIgUUyCbfh8zWzNjoE8R0eEglxDrUJOU3KAxC0bhLc59MP
AQXtOrPTY8swlPyRDFU6oifcw+7c8xaQSO0req2iIin+maqQckx+c6+Qf7XbOsV6
sNsKTUaa/RDRcJ/X6h/506T4LoGoc+GqZqeox8aeowwYbHmZtOUggGs2PDuwOiMu
nKS/W3zF0/d0fE0mO0le/FzPiR2Ma/J4xfUbARG2xrj32OXZdez95wNY9IkkMvHx
gzjj3T3j0TlAuqZ2NfRmb0IDxPCWhEmcEaeaNxeVr5IvRWlTQYEzM8jtXGy4oJRe
QUkwvcb4NmLI7T5Da/uXxcOMWpCe65qJj9AEgkIyon5NHUlUdk2gBGXRMEQtkfgx
ins3fzxJmn3B4AyVkuoVmNR1Mah/Dipe3hjYVJQ30+EeEDK65h2v1rAvYw/mybOM
t0uhjYauxK+S3ie/g6Y8n/r7COaDK7tOCus9k75d43+VA3p7SnZSuREeoU9BCUlq
1vVdJ/DVHn2k0ISNgX58Le2HdbMFtjapdp7K9tp1fmbtikS2EDSSnORHxBw49140
EYb+k8YKHXLYA7VfuswVQ+HcgMY1j3t0j2e0Qw0c4vnGhsakdgWzyDDOMdeuvU3u
kJG8ZS1jdD1Untqa7Xwoz+3K/FAfuZOsLeJZcQiciHptw5BddJhaY6S9mw25BNWT
oJ02AIcOkpP+o9OjkKwDm9cqqxc7Hf61TUzJ1a0eSOKL7Fc541SEQKBVQUXYfQ2k
XEHlGTfciLYNm9JS3NecWkKw3tuXm2APtdUfXOko0PkP/fcpcOTIKuW/pbRHMXqR
jP+fubdsV+Y6m9RnhcAbul6dt0XdVM06yqy+Fg1VdlNlSaECvr0jVeI5vN1mjc1J
65ogO4lAsMhvcm8OPhqa3glUinGw7/vhXoFjzrDe6pwGQ2Jnjt6HxaYIZXNJbl74
0hYwxNgb+1+ecgUlx41iMd8WIPhovhuc+Ng3YOK4nMKdQavrS9tDKgHuoCRMbEUO
dz/WsGx83FHbV6hr5j0U1yDEwJsv+0tOd9//rNsOV1B48UjpKxuy/8AU+2pn7aXt
aUIudAiOTR+jB8IPyHx8aZlTCY5zE5jak+m2HUUh2LM4lWW+iyLm3L0vIZu0xnPQ
ByY5Z3nU1RmU4GGdFlpLWLZsZi9CL2BzO9Uuo3N0ybkrbAIMzzhopl2AZc4yrRfF
WceDVQaPJzuNqFxmJ+UOFkGASwxJiUQv/3OMa6ZtjuewNNcQx9HOwGoGuj3zYxQ4
r1Q2KRXLvMN7prtx2fE5Hamma2QJOzPYjn6FQ8T824LMR4KiKn1wwhieeuGkJRIv
0XnkfutuSNw/jtFxCJyaylvmkvXi87hWvg9GJ9KVfbT81wBa4KwiFImT/2AZYdMf
7/Q8WRaMIPXu2grnJvP4Wvbze9eY0UGoGkIaz2APFM0Pb6RGgzChQziZzv9nkXBY
EUwEGepO5zcDCphr8+cRMHzas3jd9F/ja+06GXA04jZvIUcGjhWCSEiN9zI6BBxM
15J36aj0z4SezO6851qm+lU6r/jsFyGzZRKrA1KeU30OzpxkSCNAX2S67oQaWT2G
7WYbhGZHmvhNfz4wXE6WPNIgM8rZQupJ+ZS4jp8+Qk4O3MBqYCIJ8y8rXlLMaMHF
wysIv43rX/dqB6riH+O4z6eEvGFKwjRzis+9XOG+Enb+YVSPApJZuROiJMKBzmjA
567YyaS4Rx/GkY7kgafeWXnuFBpJzHUV3e1IBB+7sLgFxGbEYcqUFMJ3eCGc/R2O
LravpacSVR5KPdUH/SHZYJf3l67jAMVhJEUe5tzrFC07EbbvYWxCTgnRCdHpAxpd
ZVgsk7ExBajBltV/JB00la8KxeWSUPceEVQ62QS3pJ5+Lq/Vp18FakihO4XuR3F/
E1k8h147xh0pImBVYCK1UHyhQ1Pnwpz994amw5U7bD8EBYNy4C+HeA3mIBXhwLlb
iEZzDTjJB8QEC9D70cETOTz7zyFXF093/yEoT8tuV0+umZcInDboUsQ+vDpkZ7p8
1ZuAwlzKv0dqm7jGaxzu7HwpveyIusA5w06sy11fMstZzrXuxWTLYS5rwzEBT4z3
Kb7vlBN99vNL/5/fEMckVAUnUrdhvAfHTcP7hKtxF0v34A4kqyvOtRw6zUfDB0Dj
ZH+j+s4tcJ1nnpsrYuJcQ6b7bOt5GcK2ZjdeASI3PuXwzs49rAH2sne0Hc2r9q0D
15r2NR0RYWIfr8An/0w5qguZH5/aeoSNq+4cd3SYDvHGNGwFhWGURKWaiH/BMWVE
lMOBk/hBUwEZTA4J4oS0vUn6oh5h2DJuHpVsIq7b319Hf1s4T8oHIpXQ9Hqt1c1H
ff21WdbFcvOpy/CCegma+b6hnzoTDLBrSURlQGiXk858F3ppsjAtJax3IzNVoVtk
FAC77ntWJdPG7rOrOJvkmS6Eoa9duptNxG614ntTAbONnMypqH+HI/8aGwvk4HDc
WNxObHZpgDEwlO52DhYGNlBEK/KO9PNBURzx5zyXYnMsUM801Kue2U8BA2tBw11U
FXkz0uUCHws0KQWCLZg0+wXULhGSWD7N5U985wZOloY338VLoGYYE+WtlXn1vZ9C
8YG5uPoFueej06s5Jyu4jEoYYYHFMOsL0xSCyOQpbsnNaFfZhhIVTRXr6ov75zk6
yypbb/C8uvOSlfSpdfgmRzfTAQJGLq4LmF9tnStXMy9hwQ9pCgvd9CopHTbaE1/g
wFXemzgr68GVY+n4SLYaHC1uIeObZ8CBf3pwgnQUDcolZJ1PCBfstEELtyVLTK2+
X+2WUcrA+qj1O2AGR9DTFCHvBjnpodn5iiY5l6cCgS0U/Q0/veAPN3U/E1DPbdOL
G7PB5BcJ2MGnDSLxM2BaEIziwdsdHLUWqLLOkyiTONZPxiULvjlNVsIdzC6WyIGN
feKxR3G+DqkgE1OqIQxBddXZS5beh8s7WtvK02Sc0O5h/QqLm7eZaP3GH2UNAdaq
lvGMwJafTWqRrUicmowixJejSdxE0hhJzudULBfhxfAdyfA8ltt3hYTjEChFpdGI
DldoR4sSgxg6H68TxjT/FIzddip4SkI89OkVuvk06qZ5NfrWKbjJHBQr0Li4BSK4
JTbxNgGAyEndSweh0BKayZjXgrjMzOEfiGCdGuCvaMt+1bl7fJnvtT1vn/hgITEu
vLg0P1fIt0iIsaYuyUCb+emD2ipy5SjSCI/qh6ZF1EWW7q2EKsyr83lVlzKYkutr
ZmXLtyL5WcnExMD76qZAKJmPVRuNRliKn31X1/sIIOzJF4FQnfHRFmrf/BScwDrX
4g6SBGIrCKwG1Joqp8vNcdp8KkUEAqn/CBaDDzEf/cq8luhVbKTXLCGfYiwvNSqg
+ebHUoV6CUlT+Km6g4FSAUtM7z+2U/CBWLuY/YBoQcXfnb/azancadrFD+MPaZiC
/S+8Bl0sBHRn9Tgo+b99jqq+2ITB6GsK5BxbBF6QU/RpwdT8kEejxz0r46CPI9ST
czznaZ1L27KPLBOW4BNevVCmtIBpQMdzrchdEMXqICqQbcpb3Wl9HXVfExlnufs0
KAEkL5ywpcZxGigd7ecY1fKx1CEHzuPS/y6HU3Ovc7zuT+AxD+gkGNoUiqE6dqL+
U5cpVSWdvP//icQbiBZMclay9dOQnuP8vvaKt8PrKD0OpO3TfmkG+2JBZ8Gre9H6
gto1NdutJzwYlUWE6uEDKKc4g0OM3a9K8+bKx1vlRmdkIl99qMJlUaTnfNbdET7z
NiWB43FqGEjF8o+8aicX+BEI8oZX9Z4grjh8rQd/SZLK5zqPUAGg0Zj9PP5i6JKk
1OjQuZk8yH+TrdvmwRwUHBbv6Uj3brXTc5a9jrAwXk1P+k6ACPKAeml7HpbAHf9Y
mWzr10jFk6Iw1xJkalkWah67CU+rP763m7/AELFb+xwBOTWrODbbwDF7H6zM4Siw
KxfGbaGzcnCYcfAJFlS1Bc//5uv8OnbbNyoSDVzuF/syvu1VfntTf2NEwzG2fIbi
8gE66BILw3MBvpOPnOh8NztA4WmBKjq8P8hyTf5vzOtFXv2HuzqKbZyIbVrcg3z7
YCj3f2akSmCpauO5l+Qkvur9AXoCtTaeZ8fafZXDZLvhTNb5rqmXuiNwzPWpGtpN
ydvJEQtDKpttr33ZsM9amhZ8DnTTdSZLNgBnpG/sNJkbgmJX1eYnM7TPRGBYpEDG
CTSmYZuyX8vSetNq8O7MJKG/bkE22VYRkO1tt4nKbBwKYARcNykVzixK4dWOPiHT
GIMLjU88yOPaGVKRDSICU+huNArhVwslRXGH8/SpjI+sPMNT8tuC4nkmqHbXgAYL
IE4wcsPseLix0Y1Zl2LDSKEkp7/Axt5ZtlhUnWz10T8doT3BxYZ97jpE20OREd9t
jR0rwN+79ltzQO33hLiCcMptiL+b99wRtxWOj7wOdKXqDXHwx3pSz+sM6LwAsDpv
USKW1Wjd6PczckAEQVzz5aRgVNO2PX7WcGh6QJiAqAN0s+ND+GR7qTluE+WNy2sL
EvQKLPBYhhJDCZIEC/4Uxt3+vVUCd8NXXU3+B+1bifblzTlDFTvIOFoCnfdA28Z4
QODF7EqPeiep5vEjXy4EhtfG5Wq5/X+GSWpCJeprG9/VEg3QdRd2tiKgvgjcmzLC
MGYhmE42gasTPclxEdgTN5E3wyCrEDGpmcBNGMeIoiXZXlMrG4OSS+50R03HcG68
47pf6bP17MntvwCF5kTEwT62qYBo9oeD75VXL+NqtXB4SDRI2QHzPjA2f9MZDlAr
eymkSeL92e0Nm0oG4wBTtyMzu2jONCR2A5WWSlBhpmj3dUjgoFTgzrmGyBMlQFvY
D/1Dmefs5aeW2xW27B3m6Y7qEcmB9cQnqF5zWdfiH7aFLF6CzjpoWPcK4yUF8mmv
h66SaBnTufmvqm1U+VgMvweddnsloZfArAk2yvEKC5ijqQQCLFafI4QUFH+IPLAL
o6ai39EoQa550JeNhNC/Ypv9HRgkpT62Z907qUGXG08mrwB4Mp5/AWCWRmBaVZBB
f+cRi25UzOu2xa0cJE07dZGozgs/UzFWGPvxx+K+SCihxWLY4dvAY5VE7VI8VlCO
ndYrvxIsaVa0x304Ck7VQtsemtP+45zPYT9ngv0fqvm+4oSa+aAPUCAzykC0vNFY
KOUGjgambFLWh2GTmZ7FaUhdNnuGNEKwio/HpjgaQYH5x9lgqMbShdNQdli3VGGf
r/f1admuwmwZLH7GpvDJsPJQJjcxyJKVPs/ZACOxDC418gWjDHTh68vzb67/ouPi
+XUEXnE2PWXoNOsdmnwmFs3gIRq1gzeww9idDHAQgT4UyTMvBGt4ayteaGnvT1eW
yEwKW2+1NNRhqDZ7y3LQydsuxTFcs609VLlULTeLFaHGXoIiV1zoJJuh0LpdEbG5
+RtTqxOKKJ9plfQQm40aqsvQNRsg2dS3oxYiOlbgl88+/Jk4Qul9qyzORlbaNV9+
gNVAij6ig+E3ZlKH3gkos3EKIwE4maNt8kTD4wNUBO5qhQmD87SQ8mdcxzIii26m
rsKZxJhHzfybF6uovk+RW2dqSIE+d66pQiLNhcoa+4js0Ij8KUjH80JQCPjV+kqJ
BvHsc+asxlHSoacRMphuqIaLbZ2cDWjwiMyxIZOfYF1JLpHVFbqbANnuIfxevKps
6De9ePavh+WpmOvRnoNGcOYG+/nObWB3VawiiirLC7ERZean1pUTzghCaM1mnUb7
Gh5M16JV1LlYCB8S29unz1rPYhacN0xOdGjaxDulAbkLgxD7nI587jOugImQFoY5
vUHWWLzjlxSndPvliuiYp9WQ0O/w9JgFllESjqMLpmlhURUjmMuKiEl+MiHLRKwA
444EFPAjgcb1g3I0ARqKfYygfsrh/uKeNnWK6fPfMrzgt7kUX6YdqGIf0ONXcf/M
q3yfY/Dp7uREJxF9c93q0qlAcHvKWpTa5sIvTGcBCvRY3jKupFVt9kS1OXEi3gvz
rPR7ojUZ1GPtOltgF5LpRx1paCWBKT1RSJxE6xMNZKxTgL5tLpvxvG7rpMuc1WIH
H+iByD3icVrGQqF0q9eVcqooupsDEaSozc9WAsOADAVgk2VGP8WxAr47ibBNKgJG
ONpRbq3f0ddBQInFaz43KjJeIxK0xnfmE+koETWSZe1XPKPDzgjL4MpMuxaiwH4c
dmx+qN8n1YTBiQPKoQUW66SQWX1zUuvzLynKpR1UxJr69wKrlyMMbV3BR6fJ1Vq/
XQQvd2fiXOQkrE0AFl1DM4LEalADWKiYQBcLdRdt8iAG95IfakJV/wWE+OxxBrzC
x3dHY/QMKVcG1qNKcih1S+qAxoOuBSiIH2Yp1lOzIXt0NMPthwkE47OJgdYxhFAS
HBAISP6ekszJnCJtX5zesSA/xMO54y3Zs5SmYh58+C+42nB/jwN5wXaxHQVAHIIa
oWZe3d3GcRIudQqMvXnqwaZ6VCZ0s3+2GzTiKdsp1z92hgxYFS5ykiFv8jLVykD7
59Yvd+KYtS3Q8Gp0g6Hj6n3ucCilepq0u7HzVmrQz7zduRWMBdLIdgjOIJCCyz3j
PaqV2xJJnHfpXGWv70evn/JKDtAnqBgOvatZ1/gSsdI8Wt9eWbpkZ8/rZ2VNiura
xcEYP2eHGpoTREK6OYgZkHplPSxHmrYUIKJGhvKzvIOxdmDNGUQ/hCoJyY412TTB
ojjI20IaWPEkHjInUgOWb1es8RCrjgThJjWv2DtYqZNGrLNTcXJmWKsXkq/B3y/U
8F2hs6j2k5aIVAQcj56lfLnLIYTkv+0znoW8rcRWcLFrQNZTdgLpUoJLWAc0IK5C
l/QCOCsrlC71rvmBmn6IXng2pq7vAYhLSqb37joPgSrTUTMNSjN8bkwEqOrAFrkZ
YKHSYlWetzG1xLXm88F/gVN4jjTnOqUlHjzHP09qqM0gOtjQ6nvY3FJ8LF5a6eW1
sGXCUTeICj6dMlk0bNGtRQLWF9N6tB16RAg2IgKZ5luDIU5yTV94KPxKTxhR6RoS
EcAW9YC9dgx5QqRU3FZfVyx759KlWeOtuhiFTNGy0k0lRtQh0OYFnCuAxU0rhcjN
oDTYr5lhMt+0etWi497I3gXgUq/imbxTDygMfmMnbjydZPseZ6W6uAcXr/WYQkm8
lfW/odGs66aoij6drpdfDxCIj/aXpm7ZvQFvuXuhb7+9CUiDUQ5liUvBuP7pQSKL
aTuyQ4QAdeHaEx7qH5TEhjqKtggKEUnzsh00tIJcdXNvDGd2mACRfLOzOMDJgqkt
7xgKmKuZqfSZwBlQrTlCegjh2ZWFDGDgZU6+htJNfUC92Q/c9jFXaqe67X5jtw3f
NjvsSJZKoKw8xfyBm6RKPLhsvp4kYGSTMpZ3uqatB3CBxDnxxZMf8IPvY08KWYY+
A7c5McKDNUMNY5EkxiX6ApCebtwYjb/dzs+ER1q2mBybqTv/Z365TlQ9W+xaJq1x
mu0pcUEeuXUr/6ZkrVVz2jlHby7PYK9P0Jdr5h/6tcuH0wF4mG0nBDKhPw48+dQR
I6UWVa6wKBvxtep2GnVgEmFLX7cdQt/cPDXTpb6EQhzCNDYT0XFWU7dvtiVbnNNl
++xZi86HHcFa26HHL8rvGUPQfdNqnNe/8rWe18yIlI6RBsBq11duKO+1/H2SazRN
2FhjUULWBfzbw+to1sfwAPKedlFZxB5XRGG5FAGKAGAYvOiDXVunzX46u0PdCgwv
LipKp2aHrmHJZrjxtjWDSYA2GOjAmnF0+/aOdzaCcr12KMgWRaGUVnXQ9qComsfh
XtwZjB4l+67kcD7hOik9k+3OzkbL+59gq8SKrnQJWzV39u7d5nO4Sy+T3taJYFoJ
1WkE59KTsk2o7J/VOY3u0/fgHKw0zkYlEo5t20juKgyJMJK/M9T4Xo2DujjP8+Jw
Rm2BPTqpC2t0gNjTedbDBsK1WaLqMbAdPJYDd3DmZ8XTqRVPsug0sNS/J4vLLTNa
iwm6aDM0iPSbcn3MlvSetKSJSOtxYBPSytybJQM7LeFUNYCFKAj/wjCvxOpFGaD8
ch+xd69o5FiR3mD11Avt5o5WrVy5RVL+Ri7RVz8/ZTmRzBc0aXN/BiIcz8e81tzr
OnQg2wnxjWVa4B/LJv9dgMj952AeWlDpDILHl4CYGova81bCIqmBr1njKjI5BGiJ
zQs/8oHGYpNWHL2dMvHsprBgpvUtgH53+keS5SRaM8QjYVQ7TRvmKWdhZA04c+vO
JWqdKwwbjft6msn4u9dAaaBTupbJ8ShKzKbEoMbPwznGoyIbZNrO9/oE+cvGnCj9
WQG4cFvoET022Qf8f1Qx+9RtNWX8LhDluC4CBfu2ZfiEcy8UkzrQvSudUw047xGI
FCtmJ/CHg+ges8l9eXGkxloe484eP47dJ31ucNtIibQ4NTvvC5YvFshhu7ijLMPW
WHzphQGMxDmxKq3U30R/AJf1Nt3OMH0Z3e0gYAe8H5HEjVCkVtyf5E3v3VWHlRkc
cW1gRxfH20S8vxpbwj8ETPbw1qGHvRQ+r8/aZiEy87WlPaMDX4h2R8Bw3v7bMPIz
Mj0/bG43IriofQJZnpgxyLFKba4M+9ssqWLX3PO9EqbTzzqmfvA9yucGf0+cD8nU
aR1RAgHgW3XmgRq77vI0/o8GvqJqtcSP7YT2fdRlziPuJNqKe6MKH5FWVTxgwhBc
Ht5w7XHcSv5657stJZ9gl8vTKAkh6sAqcvTm2ldg1pkR1joB1X9xj/nhDWte7+85
yIus+pgzNIC0HZ1ajMqV9sHEEjPfxdwawPGKH+bW56iIikrnsxG/CqrKWZ8n6A6Z
KObhOG3r2VwekAdQwosxvSjP9nymiR1YhlLcbt5tH7QhYbpOAqGuW3etdFrQexUF
Xbx5+mXmUraAfo8QWfceaw/CaJTHxrFB7iBi9yBYqwFgC1YM2sYVd0U3v/BnFTn5
MsJY/+MWJ1SRWl50YeXewNzuoYKQwh2jrIFXf42zFvJF3aXf4INavmh6D0hJZwO5
gTJQZHAGPl3KlUXELMhf+TyhKlMdBeb/mocUWGc50Utogyrcrjow7nS4gRsJyJST
l9AyeGt/mn4UV9sgLfhM9ZUuFhDqbUdQWDu+4P+5l/KNs1rgJ0gx02gMBQNprA9I
jffe4VYKhlcXs1PXr6QEsBiTfU7uynBKw4IbNCE78h574mHuLpYsmYhW8kGGROKu
Qsqe01PrOd/x3NLMKAB6FZzby1GwYzsTgR+ztiBSF7W5WYf1BjiQQSC66Auux7F8
kz6fBa2jY/0o05J6O9F7XkwmhNrWL2I1wgQ3dMWksuW9mF3fsMhqvJGJHEPpYhRu
xPFciGo8NpgfVVIAqeqsRPaSDAU8md/QXFpTWxrM+xxvtiy0iYxJN2wE/pVeY1Ng
Qz42/T7OAKVOmOexHY1//SZd78QA3m8Em20+QSQRj55qYMWldBja2nSKuUeC2vht
LFWuNUVHnzWlk6w+xqvav0uLfYXLNEmbIr0Wyd50EJbUdEW6HacAe8zrsvqfxWGa
aDqvIaK99H5ShGaZqGQ8N+kaFG2ftjz09dLNcRDrefFBaUwMQYO3+x/OgH5iBUXj
vuy8iG31DalVRfcvJRaKbQZwEz5/uAWbzyPvMdpFyq17SZZOJ4XJoo04M5gRG5Ni
u86P+G5xhVeJqzEkJUNMcmS+GOJAH7r12bdFNnFuDGQt2Jns3Rpl0BK+Nz+ybeCd
AeXCLe80r43+lwqWWHR5mleShpv7dSkpxdMtQGMnj+XE4spzqLqK9PeuGmrA1Dv8
wTEqPMWPDtH2++VNEm2AExntz8vRHsyzOjUNpzHvh3I+R4AKIa47NV558ovCJBJs
ctHUTAH7/2nsNLBxxeSeDExr6zByLh9n6YsLqh6gOdBw/0uamefGoyVDRDAc+NW7
oBMPbfhr86CTcXbAuHHu9DD0wTRzUTwMxduIR2cJ+pbkhKFTUwbJ0iaMbycKH8vd
3kSPXFQwsCKS/fEvYWw1CWGqWkVBVmwzi0IySmoy+uFUC/7Ar7eEPfau3v2MOMVi
PikdztwgmJENorcgiotYoPCuwaY+0g4Stm92WjuCNCI9oflMobr5mUz0eGS2mH5I
1KQqPCdVkGBY0XmTrSLOSlXPp2qKa1nr/WelNi9AvMvV9ZmI0c/cZD+gCyoCvjLj
g0sKKc8vIa+1hBrGCpCnWi+9+Azrot4OCJ8dceJuCAfwuVqPbbCor36icnSionTb
qdWed+R/KH/jhqs0ReavmAIMnxwBBSJnBs4DrkFg3MnTPjKAhEryM8bNZHlYej2E
c3biALLz4OOu+WFbFznayKprEdjktCbJPTEPSMuQS182YnbSz2i2BJa2Epl6XM2E
PyPQWBZwHbxxjfKKygddR7/zLva3C/PLDj8++JXXWlV6SxK5TLwyAwlmgG3cx8ar
JA0b3QiiIrBBhj9kuR5ackWA0uiPLbXU6M44ilv5c2fvGccT7qmOeC5e95d6M+tl
JzBkZDe092FJUSteUJstxLk3WL0uJwy9cOH0tiyayUVRL5coL71safRLC/VFdGrl
aQJ8ZXr7IMDsSCG0XVy1eJsD1GNYim7FXWFW6RcY4shNdBAcVhcFMAgurQhj0ea2
TlmchKtANEhpPTXBZ3yomKwg7DU7zu0NJCpphTZuZI2fc4yuJ3WksbBZjtGbVutd
DxugLGHFi5+mbJaWTuqNdjKnE/lbfXt30UnMez1py+F7wB+nnJPorYfA7MY7AU8d
6iqlRuQw/2+/wqpU0YfxQnMAzEDdXSssqjl7JdeNqnYtGfJFuzmvxzJzG/KE5prm
hiDr6OFKQnNW2snmf4JT/6etGEFnl1EFgwI0mEtN3rSbj+z/QhX5J0g4ICq+ZVd1
aWvmzHiA0VNUTFnhHq3W43XRlXnhJ5LmoRjbKgMEwNoIGpTrL07wzD9Zn6ynpbeB
Kr2tmB8x3T+LhFs/G78UiU11Bnwzcu1PMoD7rELgzPAsRkIjkB7eb2/aSGzkZGhh
LmheyS29wgwbujkyPrwEHUljgZMNwZSKNsywPiGBOyZD1Q4y0X1efWSl+pDzMsvX
mva7X7b0BE5z12IgPReUx5Vm0zmkyM7dO81/ZnMumbyvQMf4xXSiWLDFl3EfiM2B
reX4yYTVvTGwIXlcPbhv9fHNl8I5Ao4NRck7jzd6LuBb4U4hO3/d51gXI0GX7FcN
FuC5eaHKxVHiCDlmrG5IK5BaQQ6M6QwzALiwopUCvzc73ah0bcAxGcAzTRnFgTP2
yNulLAWCw6i+Q5dQCGQTgOAY01Gz2A6Ou9WKJ+d3d/tvh27jMMtmpgASLaJ8fyMo
T9ONu/ofW9XFl8mV+Op8Qzkvh3fTW9trBJyecw3qPEAk4p8PQwwtwycNFGhc+0bt
208DLL1eoQ4zuy8u7DyQoDbTuhXassN5D/3XjAMIsCcCAlEKq/O1xPlaRtC3gdNZ
Fv+QbaPHL2uoZ2lLt4YjBKxKh6MUEo69yc+7GOn3htFJuPn6XeC5vqSHDtHQPCEI
fpN6KDS4U3VjKL1j7otO1g4VKzvdrUexjHu1efTzyQBMMg8q2vzRxlJ0ULJPTahf
up4jn6ukDoljrHHZmmJ5vwxG8pELiiaZcXhdFMFQtrXjQVEB58F0D+sA0VYfGMvF
a5UjuxIcLHEBjmgh2Pep2lktxawVYZE0doObtpBM4LMyB1gg/e8QXnGF68NdISKU
LcoF/3Vy1j84TA+Zw8cC11JmIxZbzR5knhIoruDia3hOVKkOUscOl07qgyqUgPrb
P62DTK7khaWIh/B+i+njDoku9puIlHyF6eM/y6TcL10xpRhPQpPCb6wVsO1B7klC
C6Go9m4Tdre96Mb5NixR/n+b3dS0HWnizjYK8pRJxVcNTP4MtsC542+2yk8gtAE3
TKy6iJ4eEytRyZovvWI/3q3m4t19R7jT8bC10jW+kfXD7kV35bT5doJsfT5gbMJF
SlLqaabpMzAYQfvOw74Udtc6cgcDI95x5zunxk3ujiR8wPk7pl6Uw+9f/qjvMmnT
T4GHCWQSdhMCrhKv9DU20EXqeUax8228XJyIdX1ozCZUM9BZlBiwD2QkO9nIhHx6
8LK5LjB5T8tfClZPFnHMITf4IVrnKj0KmnBmU0/pjEiDkn8JuTEjUv694tMowtKT
NGyomLVpfKr+HVt4jkbPR1BStJn8MHDG3lSp4c2PjTBPZ9m02vlSCyPPPFKHeLSK
SCYC9HS0jkQKPsrw4YFVMtlxBhncYtMwNAbjfy4V+lyuh+kAUvoMmcfyeuqEGqKQ
g0wx9OsWav704GGaa+tWTjt0XO6Tj/x2LzkhsLkyiqgUlCfFZmhOkQDjRK8xZIFK
WIhmRktEcvuqZ1LXzUG3n6AsRVg0PJ1pt6ffifYs+x7/8WQbQltcr1KU+VgxzK9d
IaONVWR1C6xrd3kgP66P4zJCulV8xqLkbUNXLJIOlprqwNiLPHXeVnivKR7ZhPLY
U2rt/bRzgN2piwi5mz02rVYQfj1VdQ1dYhOyj5Yce4ZP1W/3GxkZXUBSolMxC9CO
1cP9/60oIL9qrMdabRu3rU/na1jNeiRlvifssk0HPcB9NBcj19cUYxfzs1gZEAIv
sQPNzk3Li/cop2RsCRwxmImKt4B4in7en81VdEV93oGQDcHjw8M4kAijVJc8QwdK
WdBDcbZLNIYErFzKQ9L2hKvurWi8HgA83f+buFNTwvaRU8UR9swnX0gIVHHw+sFp
zIf4fIXchWLfHI1fyrbTxlacNMscY6t9mK33OS0hHMtdi4mra4bgBUezpSOw54ty
xxtsAGi6sh+9EUk66/VU0/UAe3fYcUdczrluMBgZvKl92cu9gnBQypRweszxur5F
G8KC3Y9XW2IhCr1PKXMJxNn5RR/0hMSdY0f9FM1LT2AL+LIMIV83AzColJdqs7wZ
qGCkHKQ/M8uMx02zy7NZi5s3UsernXqPJQHzhB/6lRfSg6LZJvpyOzIaAtQa91Vn
qcPn6i5pKEjRRACtlibqPGmONZRuKyEzLOD2F6J6Dd3wJMp+WD9XphYit2S3txUH
LVvsossfHN8fGNlUfrJ1fx4MZ5cPR1sHDXp4agQg29+PNG8/N1lAh2/cBwhnC1zK
w1Ronw1VBWAenhvwwr30TH61PRLnb6lWVNSd2MLPoz6ZNMDphlIDAe/P+vYH9WtM
+zIL4QktsGNaQleRWUYC5UIA4x6yCk+O1Xkv3wjT2UKzhTH3/St8YTbIslsSnhlr
saWUX9GzdnLX5gq6Pi6lWm2IAJgWlO7fA7VttBXr74V3/bZPOTSfsYCqWaI4eWcj
x2mQtx/mNm2fZ6DXySBQoIPlNlp5r5ofNlBts308nJUBaZiq3KcCMgIcpqrC1sDJ
DI8iuJOiIcS1WjpZp7SGvfgXIuIvcqcamTXDEF2OjY08gS+NDMqLSKd5VWsEy862
LXLOMYGgy+1dsnTovgpxnPWj6kCGS+YQcvASvxHrZF6jtqV0fgNYLBvJ7i7BJ3CC
fSv0Da0SdBJ8oYmygk+whHUdRaQBaTF8TQJ7m7YL+qs9iUwPWxKdQF4knFb0AlMg
eF2CCbaS8fJdkvkt7rCjShIvy8A8wXKuYdckuuXg6wxLNJ6So2OF0JjIKA158DTm
A2vxWjA+u3fEqHwNeSCKVYPBXC0BnL/7H82zthxwSjS3tPD9sUvGLbOhyc1wl7Py
jZjs9yYjDi+iCIS8OQ+9c7PmnsojHlCxofyLxbT/E1M9BdS5/rs11l/Fe7me0J/l
vS3qmKOIFOVKwSeMjahuTbOM6zyDo8mv7iXZNwWq+Ycy/aRwzZ1DJ75lmVkrSqak
bNKbAvGq9gw1DyC9ttr7zF2A2tMyymbQHfqpnJzbAHDxg+xyvqMK5b/LlfMYvx8T
WE4VpdOy/7zBUGeU3Ht/t5R4SUyO83PkovhcU2tTzsS97liAXGGCc3XD0M6RPdf/
FrwQrSvYGiCs7+F+Wn9N2AkC9YoNiv3aPBMlXxiIwESID2FJk4d8cektqOd0ZviQ
b/lrz3rgi6Ko0ktSMOEwh0tzIktIIizF0y/dxl7bIJBX89icRHiAb7Imioa74zOW
FUUz5bZINKBvY/GUXytUSj0/Y5lJUGXQWGEMXhvSXT6AW7uaam6LF+ON5FfOoWGt
5vbVMdrZ6CaOgEn4MW6DsVpcEtOearVpA8wUGxHCB/EdUNCA6WF/jIWpXA+WtqWJ
XGWBUlO+BHUIEF88bsP2vu8DdGYfM+7NFNCZWHydceGi9Dghq12hivP0hYMmU3f3
3IBqazKCmbTguGy4hTPrHCtL1U+N5XdzO1h30OSTpaiMGpJlPfSHSXImn2a9tYx0
vGR0DTNcKz9mqCkhGtV9IyMmL2wUTKlxN832Xq/TAP5Nqivjxj3reD9y6lmf/e8p
c8pTWDQWkNf/kia+5/vvjWBzHY9/nXe7vDWwH+Br+WepuECJC5cHiP7oHx5XjM/q
itMBeRBxwkA6126pJ+QzWmVmNC8ibg8Yp0O2P1JGIYtJFodphusJo99wkI539w8L
gnluydH882ZsbJsKYs2ukFn9A5315amoYmlfT71iox/qKcrKeMdKhveXekpa++fF
2fx1XRC8LbeROuHQgAzFm4luVYEp4+doSLq7KR9Qcfzmc3RqkuIqKDxlhReBb6Sf
RRXi3e68NSSIyJryzYEIF7qx/rSZS7CPzKKuA3pqEv5R8/UdTgNxOlQpNJ78rJAJ
b3DwWBPtbG+UH1wk0zugJtZfW1pRNicmJNNRXhoXECEZGVL/mSdfY8tMeleXshCf
40MPtnp6uLlCHcJNhvktwK3wDRjf4Ry3nENsLNnPnvPG9N8UM/qNeOuBuNqvTLq3
hfN6jmRoSrrj9Gh9NhIqkYXk8hf9ywEhoFtcQxuHU+OFBmpJ+AVwdC20z3VEYwzK
Ar0yZ+KUpsEg58A4tkKlnv6X35Ad3lwTBG+l9UKkQQQ39+RmTF+thF4krSE/AwNq
T1yjtBhGB7y/yEBXRrdLafJ/pqxFQOxKTaVxk0BPB13vHahh1MpyQmipQX1orpb5
/wQnAHkt33cNNJ2MeXXDh9O9em9SHse4DNNG4en/+sOIXu1HKmLzj+TnCYIxalG1
/bb3FmPNFR2bT9FmhUB4kGLs+YSrNQ2tRQ9kOaWKCnk86y3hC2Sc7eQs6RcKlQzS
XRzRq5aZE1tcQ8eUNiIYGw6Evkg6XNOPa+VPvVG3lFO4pIFL+Xcd3X6W/oAYKkJf
fXkQCGdqi5I0YxPpeniZKdZ4Qp5qW/3mT7CHNeyP0g+8gtg5kfLCkMarOhtJEGT2
O6xrGRbXt8oRT3FZbb9f5t5QenOFUuAVdtmgOS/3qZiAGx44wF15vSxNA+4KI7Yd
jzIR8VTG3G9sHZtBk10Uq8SI8z1nD7FTPtk0OeAK18RCx75yMHb3Fjk+UB8e/05W
Bz8EFHTgil2VnmyR9dP7loBc425V0d63uXbRQgDjxLVgbA5EGo43tLd4j13wHr2B
CqplVDaAhu3l6HNYZTfCGOrb1pr6ELDUKnfr2AEY10Q/FpIHRTY5nfaCa8r3w44S
geILYD1SmWNqzA9J2rU772vvf/oFGcmnDB1KQLo/aFPdRYqz7x6vRBdl1gGWm0T9
H4a5tbwo4SUAtfUQ0JCT6yweyecdhoSqvjyTobcEBknq0syXXVVKCovOX6rdcIId
D6T81kzAvUWaamJv7TVLji06qZBXQaW9g18usUi2Fwg3iIeyn173f8cQu+4Q/Fny
8M+wMFzizK+ji+t/88pucOJVWbj8ZditAiUbZGrrwbHakaIQeTE0To+AsPUYlL3m
ZfT1ihAIaO9iBupX1kiavy760IY7hRSR21/0jDR2FnPq4TVQEf1XyVRPEoVzBMUA
RHL+87KlQdIti5J5Oxh6uLp8mtT7PwRtbE2Q4v31IDb2llQhooZS+kywr1k6WoKf
CpG3FO/SddumD4bLxkNWtaprTmy/7Qpkb6IAin9i/xEkK4t6kzYEMqgXFE0tLFEN
aJO4WSHUMmQk/XtwHAX5yNZBqNN8p7E4khJ7vPejd294UH0c36OEuNM5v2KEyfFw
Jdi/6hWZdpC93PUqeFTY5M6AP2Mn8eKWawqoTkvOqh1/C8ZNgVRI7D6cx8Dfi2tu
JbuOLpgBdnp40fK0GsnszYSIZqNtH7Z6Ol/Ty/9UU2XqjcS+XrOujesRtdPay43P
rnlMSEeAvBWJA4nAebESmeo9ro2Gx5B89+72OUTJB6InQIUO/vOAffbreV/7v46s
nHZZ3sDlaxH3wL9CkEVl/ZlndWIS4lDv1PGdLttoNSO1Kp9Vbts7nD+DgPY9lpO4
LJ/c7dtX7uaksyxjDPcw2Hb575yOdZZ+VhZLAAuZaXF8T5l47YOf7lyEjdMxjkGO
127uiZ/o+m1qafKIIhKNrUziRKgfuzUajByeNlxXQ6eaB7nbNfY+AM5uFwus+LFm
8raYcSe93FNihzMg7buLM/P6LqT0fk0ZhvF63IQ/Ify8FK2vwh7GIPdBs2N7AzK6
EVA1LN8A9NPkUgHs9IXJA6A0C7xS5kRpUrOfo7AG0p1gptL0zdRLbMxBci8kYJt7
PShfjkVI2o0+4B3JABEQX6fWPCu3twPJLhVkaeXhfTW+Qv6FEEMorh6teKwV9Xjb
/8v+m9GRMYACvHbQUPYibQkf+cpQ/cIbtHtDbQfZQPJn/+QE4JjV5aDFlI2joc21
lKrteZoMGO1fBdSI7AVsT9rYZ7Y21oNHGcqWPJ2Zp0rmvaNW2GSnO6AA2aiBrZAF
klserYsaTEk29zGwGoSiPzSgqOfkpzn/Ym3Iw2dszayw0BczWadbg+CkIRsjZZY3
G+0QaMW/HQ2g5xv3tRHXa0LS9YT1vuYQBixyeLoZ2qbecESbXHsCkMdoRG5GE2Rn
1wQssYQgmWa4eDi/8rRqWBLK+1wdMKEAYbIF0iWusI4LY49SJZO3L/WIH5jDgsqS
59UpzrON/JQs2Tr1lRX6QYveAwrOMdKaUAOmqQ6wUJ6LYFtH5RUl9re9Ru1Y6d/M
2DR1oQRRV1xHHbDKkHr7yDWXXFyX4v5WkuFzktB0Saok2vWGEAwwiShVzL4rhRVy
HyBA9KymsSM6dBxKjY/3j8++/bNkH73u/yWIUc7WJXSgYl+8XdyhialLa6UQQKJ4
j3N7RIkGj4hEMu+E11Ks69yz67JvDYfLuZiAgUViJ5Adzh8+4U131tWJRITqxCOQ
i6/WcUz6Bb5Q4CxOcmR1+oe46mc4XJwMNU1aIhtLWqFWDQUFyBLjLd8eJnYnD72t
/7CTsRM9RjOAiRLrwqWDar7gjkACkVPh4DCGFsrPlqvUEvffSyt3NTLT0eZ8Eh7U
XS2/gZ08QrcsAuWXw3RxuinbJTi5DtOKVFq6AlTB5nl0VNc5XPj/OPfwTsk0otv1
NwCWy16ndk6qnTsT+433XSANc5MVxMu0o9OvjJbSwRt9T/OYDuL22GTWeo6RNoyR
1SBVBqnHdUrkjWWye37HbEhQ5I5/eGL76KNLJ4U/Q+ZfvRrwgHDob6bhgbvJZRM7
IDB1xUWiX+7RyP+3WcNQugZzjF2Hs2qr1h0yTkQM3RdoCkONlxmlBSdfr2qMUp8O
fJ2OeWETDP6NCJTdVeAOJ46OSdvO7c0gGrgBg2qvQesi943gsvNdrawEhbxFgBAf
ym1cC9zRSArlcO+zE+i39rH+MEpdQFSwHcdpFvKD/LB4FVfNRQLLQg1tEQJvNp2i
Lt1gzquTvtU0tXZgmrWlZLMy988DYF87gmKOlH7vHDs/CQQAczPFHbpRCzJwT7HG
/DuTv/AwvDw45qRlCbg/7x9XIChzfIIcVjh2b/odwqFE1UBMWfSCCDh5hM75lRC5
VPXw8F4zRvC6zwdRdOyyDzy9ErH05iziS9sx3UH9b2ClDwv9NACNEmXcYxCb1iKc
EINfs5McGqXtYQCMKBY7FIbT1xoIj0YWkx9l0Vx2g0XHsBtA0+xGwDNPDIBd3eGk
hw9PnP7qlkZ1o0KWH5z/RworbKeSWShkDyYMwmVVDN2RrcATJMq2BXtBTTJ4TFPD
EoB5w69QXzIzXiMPuTbjd7OVSuuwNz/aLtBqNUukbgRLMjEgtglXP1CqZuUH60rK
Zxt+gZOXbkIVO/9fPaU9yt1o0kV+yZnPc0OLeuBSnfT75mZMXNudf2CQ91krjHL8
rzBYeTpkB+tTzU4Vggo27wSs3EEqe2BO5eJOZ6VCWLvAmbTorOhx6MuwdjnY472I
sPtMKX1aB340zWTI5oWP0yy9BTBI+mv7E6cMyIGum/O8/dnu2X7PP8IZp8ZEYzdA
r3MbiNjhJjv5L6BXV5fOTnBfxNkvKqLIt5iTJjzqAbrtJV5skxDe053k04qJYzjd
i4uOLDZeFuu+EpUidiI6iiZUP5X5zfg3tPEumbbwjlJi4p+YCeE8Y2zqCrDRlE/C
/ZlWJwNn+mE1eNHrg2tscIe+Xo6DSUqjbQ84/gfQxysM8YTWuB2Vc9Jvim+PnF86
ezPaBu7npO2e8dc7/Ax9A+wiL0ggnX+SEicpVuoTRrScj/HG7G7xYjprC3+btRc2
Futm2mCFh8YXtKua7VIsFEarKjhIEeS8tvaTr3Dk66x3Wp586hfOeD+f6NkoehRm
VqVSiFLNyui3AdEMAYDhzqAFOjSU8YaQB//JH8wzUXL9VRDLJFoRdkQt0Gmuv+yh
wYD0NZOFKKVJKGvO8V8JrfMRRj0s9qvreaY7qBlgIcifxgGkmAja/9p6XRFiJamf
hrZPr8wfs2Ad0nd9kG5wjw9zYTBEdNsV01UlB+z328OIfLdX6G/mCIW6Mwo1zhW3
JxonefTLlu34oKRaIxqMly0WKoji7Y+ua1gyWE4hR+g6IUsNdDOPJaxVAJjoC23r
5uy3+cluM5tBvTS5F6B22zkURS2MS1i0Z3lro8bcK1PhwltO5MIGcBd92ut4Is9e
rZ07amaV0JkGnq2UlasHnfZLDv1JYtmD1SIGHX4WUvKkvusXMXEzHVjp6VXhhBnj
2We/dnaW29irE6cr6yqCrJq3M47rQzff7gAsHueWjanh8gTomwTTXg4s8/zpp0pP
vVWGZr0AO9yoFRDzhO3GgD4DcsID2H/m5H+UsoqHJj+4cCRXFp5wzK0I7Le4D13n
2hXURUU1J89sfX/vQ/yFY3toSE3N9PKanh9ajNJFDa2Ybw4WWiFap383JlE9rjFh
+p/E8AYbJ4vPzyS5IFwmwxC2DGAcVXG0Rm2h9mFlzLYt2+yc7vMNcCVyhJDT6qeS
aPjoAmKYJbeba211a2UYq5dODXHK8DGSBOQOGxYZ6tyMGQKeyr7WHa1ooVT1Doy0
hBXSpTk/8jhtrEQTqkS4h6GBeMsMwNedArwca34nHkg8l2OrvD7a9S9yhcZq8LgU
FylRnjU6k5/++Oj097Qi5s7K81inkJZeqKyHu81FaOiRLTe9djUIjKdv76/ov4tA
lMLUfiPhetvEwDE1Kpl5zEmzIDVn4uV16GM1jrc4Nc2tgPl896gSLRsTuX2kPa2x
gvgAiqUoa1Ha82M5fQQfRYI+sTfVTg9PwT7/yIYdL1sol/h+PI/xDkfcxUxgE8BM
0T8FeUweHzLu3/pL6m6yaIpmo8hZK84ddiNjezKVPY9LpURL9ok8poYiLRGtUGUb
e+IxNWlIsRuqUdGDsbEaC0TbZYWWRmwyfR0MwqjDYPnYglNWmxSD2SXLjn/Zatgc
sp+w32f/t07cUlmOiC/qfM7GCBM3WcDl9cUJc2TaV1ImzRmeoNuH1swiUY+Z/KUq
NJbBtH/teg2pT2z0tn3w5/NGXZUQ2zmUZyDhv/kKssn4XEjUrirvwIsUHbcc6Yj3
eBnRh81hlUaGaYXOcA+I2wHlN0NB/bc1TuyLL3Ko35MGH/2UomGg7bCqbkU2eQ8F
BNOBB3QT+FJu6+CIIPThmkP+AKu5B8Y4uaQu5pf9Npf6+r9QsGBSIcDj/xKq0x9e
NBe2lBWYGqJP3BkldIp3n014SakkntmJporXdcXLVzIhjRX8OZv/HSIYBZP2iIev
Klfmuv9i4gUyNDmSWXMWi4L4lTIYzpLSGGcwUlgN/Hsysd8dbQsT0me68uXqfD5k
gNdlP43dfxpqhOAKhT9q/ERW3sj8Oo/0SKqTWjKu7V7Yct5kXAUD2a3+XpWwNQJv
ys8B2mvOGO/vQB6GD1VhcGAVHKMoL6sapvwvTxrLjiVVx5dSsWXgMh/WHZzT/emA
jzZnyiZYirDsl+RNI3L09bSfjefoujYkj3FkaCCtH042sWZYm9tL5qM+oOU+RRXk
sRhHAoq7BWW0rilKOhG2kC0Hd5fRROI3zDmU9LCUQrlzAjkCoNwILfBPGis6BZI7
lsxWjYvyAXvvAdd952kjG2vMmCg5tTqIwHcYrs8D+ZfDGO7+5x0u165280cnPU8G
NAfeD3ElDNRXKQ9Rw6lJrDZXQVma4bstiRic7FPvtX0ARvR2zFjABIZL41/bgHTh
qzr6Fv3pJCmMYGbyjUswpiF7WBLOZt3REBD60U5w1X7tbJVahc15yjoTi4T928Gh
XsiJy2n8yF53gRwT5GvVpFaUWRxIR4UQRNjDrG5mGdx2OsibS5EKn+03/ROgFoEO
HkDkALSVHYiop6dyLODBZincb03MvaAgRrR/SSyq6wtwa5bJX6+W6w2eDEGuGll0
XdUKhbMc0N6mS+Zi6Jzdx6u3PrPCm8aiQvzxNzQjKtnk9uKB62KrYsr3K9PnmX01
BPGjL9W2tWWLJjj/DkhL2M4vKDY2t6xTO8YI1S63dVcBHaFEmtE29+GsG8dP03pk
XtAAjisvQhIjys46IPN5tIR96Jf+3eheqk7w3N5BL9QXF19dEcP/eOUtMPn+I1ma
9z5HDMUtQAuRFxQs9LHsWPxF4FOcYXAdEi/Z9HrsUKqH6SuiPhGze9TBSrqPPhrb
VAUnTlNgMjB0Rdh7A5i4fQkKMDvsyHNjYglHYUXP5qt9lnrsHrw9gyw/C+sgapSL
WUr3u/tg2fL6h1mkB1EkZIEhvDm0RZXy1ii6WR7s+5PQgmqyOOZdbw4BD20RCYY1
L7mxctAdYDzd0eEzxkuTJ/TI7ZkfPkeHLwd4G9pM8XnonS8C9WDYQHXP9hMke6Nk
bdbOuq9BnS0sID6Sj44w2ZPikrJK/DOM88tj3eOyhU9G4UFUTcd7pYz3FdiOXYr8
GcxB0Bz2QSdtykcjWs9DKJZwN+s6tI/F1lAsRBBpWOrnM5X4G4nohZ3dEoXx1OBr
Wvflh8vkGCJevyl74DhZm/y9Myn8lh2pvwzlnEnQ9H1IG1IvICzF5/IQJ/fohNor
3nfyArVukFVZQdss5tDJmc17EBBIojKWX5Pns0vExzmuh3EKbG6sJVvX1sHF3SP4
7lXEYi7KoAZcBBqV7cFCuLBivAzyy/TYuCI+j3qm5x4OZyvYJS8DSV/d+aUGtKJS
+0npZjYdEEyY3zMBfdRRYcHHWTTVfbI8Rfje6cCsQl+NebITMiUNQ/PxWXPZcrmP
FCutarRGjeaTZOwvyv0BnJ8h4B4ZM3ulmjhGDJTebmuZWDEwwhoLKVGz3AB2Os+T
CqvhMspOk4HxOnslhYcUxcTAUZvH6Ne+PEs0C+Cdnvp1EKNWPxBSITMDxX3Vel6F
gC4FuQLUoy3ajZH9V+1HIUx1TQipCXt4qT5Lgzh/2cKdubSABi9eYTvZbi4psJ8k
vYn0e1EXhvrYIgBGtJvWgHnNdrJ28n2qJACUm8FnfQEYfeQjczNp26MSYu1gaWW3
yZ/Q9Hhidy4GVZhdl9Cc0LoFTOjtIEbm/MckHrVRRdfZVtkQrhkOQcX5qqbxUC4y
Du3UQjZGrsL4ucRnr165o2XeDzHq9lDLXrpLUUF/8cbB/F4e85RTP01dn3j/Hg9K
cZjA5UK/ixFvxiUTmD6L538slxjVKc2jp2CMG//o6l4q05ZLq9YAUEIwwvwLduGO
XQpNtYe3HLcei7iuCxCqp5QaJ4S6LvuJH3IOTTLsOTx3ROJokUN5BoiMHF7LQW+Q
5/aorSs7pVv1uLNSW5qfkKjnPwFZlALfbz0P+HtQtO8xbA4SRCQna2OoFyIHRli+
DhQ0JtptAN2811ixyX2MQBQkdciIifrTM4kZAXtIG5jNh64gPsOUnELBiFQI4jFt
sJTEQIO719zP3EZdyS/SKGJ/xp+FDf3eVRf9ii5mf/bhy8aMgM2R3fUh7YVGdIqW
tM9MQZlw6R3ZnAsMaGqyjGtIWI5eTYseNWx4q13HAv1EDZgA0jxEVdf8YYQ8MWuI
pbld7UtcETrjR51WSluMN3GWSjjvu/S4806uOZDnxyG8SsSQdN3OgmeBEIjk5Jh4
dNvNy2hFxzLpLaXy3AFxAUGzDdI+3pyP5EoEqGpAl9b8u1jnNSt7b9ggcDB7ijbA
jF7E9snXziv35rnyVrC9Ws1LBdQm/Xg3GtGj/WkL7PxCN+27rrCy9Sfn0RRfF98R
w8byOxZ6/VcWxXe0xdo9m2ZLA/vOXKmu9j8gaKlQW/RYdGkaWFjOwUyfu6PfpkZw
C0hlRUnibkNOHtW5QS2geHSvQFFxZpK0u/GVWDHTV6wlYoVigIznXShBEfFhibVC
nf55YF72Zw1hKWRMFZIfpU9RlhHRFF1kapMg9B9voV567Wj8rduHmA/KcgVKAwGO
rpYFmM+aqC2c0OOfJGgPLKY6jNVI/mHPHv5MvQt2Q8v4S39dXL3NvWHYYGhCoHsd
qiPWOJe8gxnHEpJ4Cm2hpONU2MLIGeDmENvunmuIaL9zQwsT1ZxaXSEsxIWwhn8v
08hPoQblNEQcA5aAsSWTEBtQWLXmIJsqS9ZIN8glqn/bdruGDKqHltZlu3gLShrk
TVrpOdldoKMMNZjV9p+7Xr5gYgtge9jg1V0S64s34jzV8eotC3wcelNPTB2J5818
/gMmJVrA2J5V1mUD/kfWb/8r4aNi8SQhfzEASvMDDQXBOm8DXn4CwOn2184Ti+7z
yfFLP6rr3ugsxOJthMIKssfz7UbIbeYYQrEHlZcCXsbhuZVLDU/bGQ0L9N80wwsQ
NiXfYb9iGFOrUvFxXrj7oSrqjCjlmVhl5387mcw8Bvoic+Z+N7RyanCXtQR0+iNr
oHDWRuTePY/a7Tr1Dt2u88XiScGAk6CZZXoR/nqXfXmqcH+aKl/fnYTxAIcqrN7H
lIKSi8qqrLA3eRvNQAgciB4cLrRpQZ3Si/s3ihk2Y9WipfyQiI/bDZd2F0g3bbCf
OcB25RZkei72ANX7myPg5Q9xFMXPvLbade9ZA+VOJfykr7uLzsPenNq3/geHWTDk
j8rTd8HgmHZ/GeczeMqGJhD+jniupfBCx5Op/NdHRBaU6yOEGmaMt785TwUJjzqd
eKKbmX35NbFk1TEFtF97Zo5r/l2oKd748g5mUoGukAf7P+35QTPKOWiORT5tUPKk
U8uaIC2PkLY9eFkjhp0zvVeY1Sy5k8fgRGFJ0XlLMQ3xYwqJpCvBpfXMMC58EcJh
cVpsO+xju+ansy5UslcqEu8BdfgWLkHMxIUf7BbcqKovVchsxWhssjyEjPoo2GjR
W4QKcJStELCYOtCDCAspILoysArqYPwedUrJEgN60XyoUcpNO7iBk1MUgtN6uMhx
PxEnAt7G1K9zgcw2Wo1B16fYWJj98mrrRov3Kkcm5RIkDASJP52PDKUHErq3neYj
GxwPxh7ibg5uTf3HMhhHjnqKQ/gbGm9YRU650zP/JNjhO+HmGTSlqyWt4L9yK0Gn
FRMC/8JFgQqhGmyvsVi+0hoAeCs8OiEu8MCxPu3dfZs7IFk94OU7W0AiZSF5Z88Y
+O+W6zH6hCpwc5ytSjVsRaWpI0qKJ+6Ax8KI5W72u7EOtlQxJb0fiPNcP1Bgj7UW
WO3Xo721BFb7AdLvdKbO+TLl6yJ0Ut9Ngc4PI9PwPlOJKVH1CgJ1HOeCBWSME3u1
9T238lye6ROmcqay82ev1OZDlGMoKNgSMrSajACmtIVxB1UMzdVsNaDu6RaLQYZ5
PC/l6FTms3tDANkweiyivQ0Pjjf98xWeYyBf0d3I6NZ/1YG4c0mCcDWfEmyD6rbx
byLnJo2jyqNsaued6/CS3DcRtxx7UNCsApLZZ5ev27eT2SUjm967ua8E9k/NpW2/
syt3tX6naii9BqaAbK1FpksVyMteXUFq+CoKQmcQKK5P60Mtuf2AzPlec2eoJjda
ZQHP/7hOuGLsuqcuGwGLXhiFrFqFyaxBeIkM4RkAOLZz8L5GuZqLR8X7ZhNt2frx
VUCJhn8Er3f4SelCk5zONm7AK7dJEjTHyYhuKMaShgX+gwI/soUZmSrrcPt5LYKB
dG/rmg5XwSSi98haNUrKP/k8N92jcdX1uJyqE197RkMO+GqiWUHavyfqvn4WZ7lK
gqA4sjCTEbQrCDDXyqO3ZeWcynbHiVAcG8zorUSI5ccx9pEHlxa0CpDLUGBY0apV
jM4zfceCGf9cwyPDQusqM/IyOM7jMAD+01Tsh8MmiDkh7eYSu7QRF6f/Yqc5Apwx
nABlNF1RuXiDcUvtusXbVnHOtbVBHtl2KIYxTGekoSqaW7A3RasmS1zri8bZPk+g
s2r6fauIpnwm6knGgbzdItZwPALGzUditzj8AdNnb+NTqe8jC+KsdroJYGKcX2T9
kksG0vlYtszYRj6eYI4ms4SCeHc+1imnOLsi0Uc0MSvNhhVhHtEf0vUySjQ31jOM
64AKXnF8Q1VMf7i2vkn4gIO2dum/ld8cEVtDPOdbpnlGt/2yfkMP7maIdF+xyTJz
8T5RDLhVA8Wo10iZhLAU6HRZymGDO39dP6AZiKzjgJ1/FXc6NM1x2td2K1+rFLAQ
Xp69YGw7k5gQCPGqwTtY6tkmQH4vM53ZevA1lB4gjnjjf8NhViyfS6kDJtLhPU6G
iKE/YeySnHg2NFrqlmvKOs92+AcXfmAttaz2TyhCm+atvGgiSZMC21dT2qQGOfnc
V/wQLfu8KDVlBYaW6xPM0SMeJvbI69+0hyYdkj6kXrxXg6hnRyUXLMveMbMfBfAM
QM+lTynbgDRNF46L82Rd1owZQONVbKCrKCog2h+l6O3QBaVIWHY49yHLuIE8KI9b
McVoCYQpJnb9wp+81iLnG3O4cQ2zHHgLlNDrOQ1G7+vSMjNEsk/2+XuSVu4Xv/0j
w2nkd5A9y4KUPEcsnmBXPZUg7jlEn1x0ViF+jPXfYQg+DfolmQPslei3DYFA5tc4
3GVxI6qMLBqyxiU3QlvQYA56Qds0+wbxM19F16PgQG58WKl+5sn1jLTdvpSBFucW
KYRWBRcGvJfdozuRoRRlpOZ54ZcZqWSxT0zLlIeL/6q1YjHRWbDKShTq4k4rLGMm
tqCThCvQD7sZQVsAIR0w5a8qM97aRU032QmGPG4RtPCz1RwPMBG6a8eKUvmguG84
t93UZQd+CwxNbDEeiN0OZxyE/lQRgyJu/5YF6w+WPzDqnn7SO4JjbooH/kMGEg8r
V7FjAOLF1yzHFgR37x2bSdkyVZp9eBGVqXjrgDYLxMS5zu0PpRxb9M7f5/EUgqZR
iQPMzdjzYKEuekEt6wy7ERpUxzuHdUE6QtsoMcIOaebTVM3IJpeZMjX8jFryPhY9
POjPkP7j3gbrdBhytCE9+Qb0fISnkhmKTjW9fwJlnt4A0LvqBjLjDSVuaz7bVaRa
Vu5U8pUy0PjrK+qeGXSGru17R9+X5m+AQSP02S4nRzLAhRS7O90JsjLSyrDxTSCv
gKKXu/P4fIf96W7nEw8V3DMuwyTRZmZejfW0FeiNYblDZ9q0xJRI92VgK1wE6hxV
mkW/fSN1K5hKon8VmhBcPjTj6vG7RPmBakv/JYx8zTJc/1zhR7PAzLBfikD92jJu
Qr9S6gx2m+s7qsl9/LvliD+2FLiijH0WQniVpiFJSRTEJmKqkTDN2xU7QGF76bsy
zzRWjFD+/1SqA7IfXGIuzDKGEOBGo9KqpeEUuH/Tnm9FIQQulhI2HHC/z9k3LmDL
tbn34WGrb1CJICFpQbmf+AOU43X+d7/BGFLJURHpmTKqvDKamkY1tX2mtYdJCtgQ
9qDxiEAV83X+4fXLPWnBho/3uDIVXJjt84fkDCiR+dnL/9Jct3MP/lLlzOd1T0kU
Rz7NmoEx8QL2UU4exPgZg8gI6hoaAQ+045pqHXJYZ4GWUsNMLKbXM4LXFiiAU7uW
ZJRTgbSPhV1HT7EUQr7YoufXYpj0vlGYLM93jm7UTehkbo89RtcsICGVmXA5rcZv
pxu8sGPwRHlxvAE9Ldk/PgEDawmhUsVyDyxXklgH+VzsmB7emkMB4AK2zqe8YyP3
hGG7vd1D1HHCYH/mACt4wIeOVs0Xwgj8EA0SY74zsnfahQk8anYrm75wYsB/FWzD
UB9TA+CzYE1hKg/AxyW+/Nkfkj7Y1E0LSYoGQQhbU+JGYIJO8wZBeogaJw0lsuEd
s5SQFsb0aawYWrZBGdTh8vkfQwEJAyDnWbMQ8Ox2iXA5Bpo7HIHHkFbHhHybGiwA
y8BmQ470UJC401YvgZZPdSkw3wgNQJ/YSuSvKfmghHdsx97WvRFXUtilYb/mUe40
sGhcJGMwwCeUTmm7PtSmBD9cQirNPwkgpaP7rr8U8sCDjS6hptbQx6ikb8w4BLIc
ALJBx98Z4ztRNncBYauwj7WfuPhCX0US/C7dgd4mFXCDLADQCTNvj7sZCPkudW3D
x9TsVuN2c67XTucbc7+lGRBMzwcpAdcHRhYJfqVKZ2w4EretAWdLndyS9gh7jxLn
DuoFnJGSZmR0Cn6NDQoycDeVHYERHzPSiTeVFr0VEffRzFhpKHOjhGsedJfhZySa
VSPWA8RorypFQ+qHvdjVxtAOb6989qQORvNJRLyVjiMTW5ZvBONVZx7uUS75UGdN
ISWZ8JSPP5D22Gb8sUQ+/xOQNUWroIn8agjj3ZbWCUwqqonSmQ4/uauMsfh2336o
1d/qhI5iruhluHFyrMxkDIwUl4qd5/BBUlSQowql9TX8s3wbnNBhCjMJgWAUxw1R
hZr63zWhe0zmsZzOmx0/zBRy49q6rioCxwa6i/gbjB7qYRdzOOjfsKbazcuV2vpd
nZYccBCNbRhwtAbf/mOvdIcNYjyTtc4HGT+bs3X6+S5bRwMFMcuY4x2wwpZw5wYD
XhAIQIavOc2JSEVHNsiN8e82iEYUAr/tonJ2fd7Nf8LZHjDf5dVql3jUL/tduinX
Wp0zrc7auert4xktSRxtsjSz8rY3iN465dwJT+LCGQcAHN0qJmpcYZwP/ohU42Ee
hKB+SUNz2uyJrvSWF/NllNNqYRXCMHGM1BkpCqr8eVw8BgNM1UzHP6H1VDoJZv/n
CfktPlOH6DK26zkWhJi39jhmFha/Dqq5ZYnzHhFNtWhEct4NnVJMJdX0F0hezMoT
VicDLp2URQVy2QWyJKpCCKQDWKy220rl6TRHjv6QEehAU8a4zaU3keZpzfcoUqvB
JxZ42/qhPYE1IXJja7CFkWz7o4CRfJxUT6GkiIPNEtWGak56+A5isFqS8n+75K5z
6iEyzDUzxKRuIInoy1Srb9++q8bzYFcKU8z1GKq57mRZpIfaslEx5rrqBfyHkbYb
1qG33D/QGtNz4rKMhqgYBONmHn92Yq/lHbbdPTQeZUM8iAhC49Oqq6DC++AiDOIB
j2VRr8I4D6JiAUeZj0T6QcuZmfx79QNXqOT6GFbcxVw1t0v3IzpIakRpxR1/yUz4
dIkZ/P+dnyzm9dlWTMgC2pXWtqI2AriEibScmq8TvLe8l3nCkxECjKvbjoe9Tziw
x0E2M/6iHLoYNiCFZqkk8qBqa8fn7xZJJ+y4R5+HiDE2TP2R+13z0f32eIml1bIy
L7DO78nlEgO5fnZmrpsIx7nuUEQkSDLEaCf6D13DeUywz81xMyrge4OAzZbi8bGF
3bA/RRY13H1djj+jZShB7E59bg0Sz1+z61VtzPfvDNWGZ9T0i3GqjHqW6X/33Zik
opKoGOtgFgVp/dmjUnv+0Xr7YiGbKvTQffM0XYXOSdIZ4O0CwKFeSOFCYvBsek63
8qTWuoGN3rpTeAXEPk1jcTvlb3bLxOIn0bECz8ZVKjOd0hIUbYPMaNCt2M0xF2QY
LUHJJp99JOTkVRgrSkce2hcm8HXWTMYukrqpE7KCdidwtJgl3H78zVG5bgAPU+AA
yYQQLsko1X6NF8JW/GqOrRVHftTX6UyFnXBRXDFcgwyzuvvFM4dtlWc8PtAQUuvP
Ul6xTemvEV9HixwaVjGZAB3e4lYsrYNj8EBUrH7rHjV0iphZjSfkzPVj1P5JviW1
7ZcNNkEy4kGdIbhFMvXGVk0xbznilDYOLYLs7J/xKFmkSCtOz3O+0wnJTnPc0Prt
pTxWfxgNkqf2QC2zZMLuO6huw7MiT1X0UURhqEhXxseS4chroBbwmjjXh4II8YjV
nCAqcU6z/e6vwF6PUB8HS+w6p0yOHFy2txzvR7l2as3QDmfM1JhxBrWZKYJzzz27
u3uDu4gDBfKm5F2mNWqkSy/tq873JEHTznnoHJ4UaVx/VOnaxCAsgv4HUVRRELFG
oO3gGkBsYOLQ88r9Y6YO7TJnJpVU9HytEc/bQVrFOAw7u5goIwQYXg+CFnAlglWH
7Mg54bPLDiKL92kzXQ8WHPxT6/1/ZOTa7ciX5NXMSziQ9a/GXQn1lDDsGN8yzAIb
QeazT07eNOu14AkfxPlObp6CJE8ethAdBcWX+BjlENQw4tknyVJD6t32Z78z20Zz
++WwLX+47Rmdnumwd3NEp9AqJ00wVGUt+F/3p90NcN94P/t9o8PssGlBuK9ZQChs
LP75X0PQNDHL1sDFOEMU7nw4uB0L/Dgtx21yEwlfRAJVyJ55amLfc/1lmc9CEUXK
PAoztjBzffdpr8bFusy9C+bTylrzOGYZTGmC7E7cwzppZJ5fnggj8BqRmoDAKBNE
OMuCrugkMHx7cxn4dzEByzdSmPF1CfNnwRZ+3QG0yL4V8+zxz9OEp9d/blUzN+te
NmvDP7zIrRz4dpFmZeUXIuM+cZuivypNbqetAmpMxANoe9vx8bzsjKhIlOqXd127
azVYECC40Z6DTGmt2AuvtRdMV6VVteHhTcNN5kNAzb+6jFrJF4IK7QSFMSrf/VNn
63mIFZQ0SeAFwMcP+Hb2U966ABvfTdv6k8ivpOygxQynhCz72d9VaYJNbWv7gGSr
e9yiJ65s0T/vjKfj8jWyKKuIYt7Zk29QTFkw5zuIAMuiASBP5v5K7k3/5rLmsmok
g5SFN0SBF+pplDphrkCk4UI0H/NFWfsRwLjTMeSHlEsaig88EaxP4JnQwo71vBim
UXYnSFvhJEdVYlExiEQCiQSIm5WAUJH3CKz4FhOi1V2+/KI5JtI4N3qXi1kVb8P7
mFGelmucxAkA9FiftPkdJ9ykcLzL7LPHYbuLTp1o4o6deQ2UDC1xGoPliSPUlEsp
oglNrUB9qSzKVOR/NltSdWd+HMa0tf9KC11W5XnVD2X9+egtlk+DrrLQgl/3gyrn
bIAoP/J+U7w7vSFjQxO02tFiw4iJkFkzf4RfbteUZ/2/PFZzvlKazow0DvMeMNYu
Qqp3mnH/VZ1vpCk8ucrmOMZzZ+x/IKaaTZMzNssArJOSAt/rfD4fmj367dbeVi1j
cK4Wpt+T1PlT6K8iW9cgxgnuJqJKQUnHNxblO7PIY2clqjMPDnjLVWI5hg1+wPH3
WTUC1P6wFFmiiOTK9t7Hd2FPTQymhqf4M2T7K0B2rVmZRkzoTq+eF0HKk6/enCma
n35DTyM9xCYfP9BpluIdIQN6s+/R7nHvyK8ZRPx4raFpzNf1qP+pYCcwEBeSmo9U
50tgKiyQFI7en+spTk3P53TRhiw6IYzIUhZ0tdNZAIsW2iqRZXkg92znJraxaYqa
23if+n6dIk5cyfBQNZmv73iRwscFwZTYWq4LJOFqTfUe5i6CGh8PaXS/remmMzzN
0uNw4qIjIwBggOQ7j/EoKubeKeKjgCO0vTkTQeBe+llw44IOywCVCZKtum3qxF0H
UGQq9BsB7wwqUqzCtUsUMI2FD106/uqvn7su5Y/MKhGL00iM9sZg5dD8w05U6PgC
eo6jF5oWuOlFdaRCkP+YsPurOBO7276LFIH67nrp2jAwr8e1/KWSsOJSIs050oE3
+Bz4GDhyKiP5f7MEW38DrF2TV7bOgftxB4yxKlhcpcEilXcw/ypORdXiu1mLoytg
FXY3a8t4O4v2FfckqQcjONgU0ccYlO7K9gpCAgNarKT6blhWbVJmerl3MiUhJlaA
NBFB4kON58sR1IpuayoXdD24g7kEqonaTuCEp7AnMqoQ0PGkJtNKSBOFudLuPB5z
+WNucZulhTXp1UZ8KVU/8XhzzetnwAOsG1G3Z807s1xZ6OR936wmGZBU1vOvorBE
N7XwvQDMFIgN0jSPdqr4cMxCtVhDQV8lOwhAkfsLWXnE9ka6ix6p0xEjyAZnPaSV
8/QYw4lypLQjs2CZCb3bfFVeeBUlCwO4GDzoMqAQseS9RBex4rVlCV0hMv46e+IE
lZ6jIaNZLiKBpJhxI8sR3eXjS5w0IB+2c0A336jMrB4FsrWBEdAjPDQH/qdf8QfH
+ZIU/5TUcgrW5jisfDm2YQH0Un9eaUxqkp5JMgtJWgFw2csfpGj1HtayeXONcfQa
0fiMwQIoxmAMTSau/wLgjBSNshn7fcBrh6L9K55LAe5iPDV4HJxyK/gWrfs37lZ7
RoNTQeXztFuFHLr3E67+gmVcB2wcqe4RxHPTlKT/iMdFEWlJ0BiSZMwLTnsdL8Td
iUFw2rOaw6Syrfj0zukNwrmoWV7TFL7xvIxvUb8dz/lBszfrTFHC6Bhw1CccPjid
bLnAaQiSJrVa7yzKoNcn7A7JatK3cAFthcRL8I4zcwiGCf17jb2hUmt5SfZ+NX3L
lOGPZCtoqTwP3a4/iUw8cegsakNw3HXgZM4sEUH5x2S9PqDwk9+IjntAg9VeuprW
filPFBsxrzlgtuNtWI7E5Wog02LV0rrhjXFrf9KtU/O5T1MH3OxhMPpdTgCcZz8s
hsh8UeRZt3zNvDaX3LKnTFpDFHNhnBkTtv1HKgs7EU8Blr5soJ83ScgST+QVkCXs
bJw8B4OLwPr5Nx8vjhXymtn/7MyliSMUOGpBv/PnWAaPZ4lv2bSiQ5OtNM44xg4N
2gHSt/nZ7lfACse/QDNbCbB69BJOMb9wsOhBDmCV+j/S8DhDIKK4avcTymXmxb1k
pHRBR7E3xek/xZtviBrbCXQn20PGp/1FczAt6hn/JXFl86cshnD8SqwVVTL5gkPT
AKk5zeRTzekW4oEn5cfxcsrssggREYta6IfvDAOz2Sue/ymY1zrwXBHmN2K2q3ns
BnPh9jk4ZubU5lJyBoxqob26QttGasuiE94/7BnOdrMTRiOtFyWpblXwBajK1e46
nD4whxz4fkwMtneIHd7TFACFyAq2ldYmPLsbIta4xgDxvAlIXRbMCO5tzi48jqVU
GQjXgnUeZaQeB8HbFKS9ZveH3YogzKRH/d5/AOIYmTn56fmBgL70ISLGQcnKffyM
P+0sYISlPodFuzifG/qIio4qD95sLAtJV5PJ9qqDraji9GV9KoyokpgDO2O3Yd5n
BKdCDBaI7Nh43wwS8lPO74JrCVGGyL2xVJZY/hUKRhMgbpwqohJ5CwBF5eiJsLRE
oNr88OpbzzNvlgZBnke4oKJxahuTHqjWZyQyRVkJJ6qJ7URdSU/bkD+uRu02RbRP
Jq+DL0M0Ug5qYOQLyogXNNt21Fg1tn8F2Oz7LDZohjTVlYgGEvm8F9F9XSLkQ36C
aZfZEO1PUoogve5IbjXM/fImr03m0lpG3vz9nUfU5vqLwYOj0DvFnWYyhv0WydhH
LFeAqFYby23CJ5pCaNcay09ZjayTx3nvgZ3BiqHNeRdr9EYTV3/jTJ5TujDGWODt
mqM1hbZkzckFM00I7oYXJqM7g2bGRq/8B9JsxoxO8vcW4+ai5bbv2rgVWK9n2lCy
HMdkL3yGZVxxej98zCnlOszj0LjlnrmMM15klfzudm6MsO5CX0WoTiR4pM/N2McA
vBIKu3MLKE8ii2qmOXiTGtp2XDA9ogMAf7PjHgWsmLj/7GvbiFqMDrHcWiE41uIE
FEashoJ1E/PQwyHNRVPiCApHZbUG+ZNpEuAEf2m1AfBKNWMx2/uD5i0bN5hPha4J
r3E9/MB102o7mZlS0yDnhO/XlV42VTAVw69qap8z+CZ631+51ttP9dGf2k6Bf0/m
kfol+DH9w5/UbvACz3Rjf7ubJvTsAF2QfEuz1Gb5q/AI2uHnfmEIU6AtkWKeYZVi
TO5shHMsd6Z2T9D2y2+ajJ9j8piRUy6SmmfMJX7+4DPlo4HDZ7klvYHjAcub9WK0
gpo5F43IZPP4CN/e+SUkJF2mTBtPBv+D/ANa3z2gW8wU1qtEYWOWRrsrg/VeL/r5
LSfiByZrIq/URBf1bOVCTYQle+vfesgoNoDJNp+qecRQ8EJa9cnI/29cQG6L9RFH
vXzV0A+9N5SSMWI/yMQZ9eyRGAOHyutyYyXXFLAWgdEGNwFcwPV0c7gGZ0m0mXYD
C6fMa68wFEqUQ2rtpOb4MVUx+/dolyUKJezumehpkjmuVPM8gWFVo0WhC/LCqPej
hckEg1z8xixowVbKXB1YhR4I/drsOMdjpm7TT2Hj2HKrc41pZnJ2pZl5/6Ep3hov
GCVYjp1eFIJ7hliNPQPZ5nR6/pcqBktWU0ay9AdbZKlCqHunbUR9y3jpUFIey06H
Jm8w7w5Ma2glbJP+Dkgpe671H07wDHpFCbFCt7SspokTR1UAXjla/Pcz85WJdwUK
UVx5MO5BGjbqr0h5ZJ6Oe11yKdTz0AwTx8lw1wBmDBdM/Mdab3Pz9yWKEuxiN2U9
xERVSHYyF5LptUYl+jwHbTo8h7VxTP90l2pyoiLUec08OGzXVgCqr3NESAxDSbIJ
PYa6CDWiXPJX8mzgf1N++YkUR5P7ZWWTgSZXAMThzv3VvP6DdIm6uDoJlLxY1dUm
m5DqlPLZm0oCc9RsLNrg6XQJKjtjc2cfVCNs/o8YPDRDxKZP+jK2qp/6Rxtlf83S
2zOpVAwK6BDy4CdZ5x164TCIWptPX/oXFqJUjBlqMeSLGMbw6X5pfMBrzS863N8G
G9F5RKSLDjRwGsGuTnqorvA4iRAWfv87MvmD9jGoBjzv5oWMWxELfMfpnNnA5Xli
cW7FvCkeDEh11Xd04fqqXwKLonUFEM25gsSTqu7VaH8rcQjl8S9u1HFLjaNFUecP
wqQMadXmURRfwdS18cwwvq13Cs6mlsTD9m+LeRz8BWudIPfu5J75UlDAxRyhH4vv
YKpvYxd7Ft8j0gf4/hAgTPriqzA8BqFzwFiGoFfhQFbhBePe4gEQbu65AsOKUtl2
Zb2Y8jWKm4MjW5/Igczz2XwaID9ZZ6Plexht2cozs/KHbyzVYHzOFFhhaGZipuqj
TqcYVHGtOlo8xwnjj71jg2DVceGPGyV9Mafy9DjPVyGK3kcYqHgzmRO2T8AlpFgG
DnEIMX0vpU8rHtNfyXHhH+T8KjMvbpwQ7mZKpgyxpBox+Sys8/aQkuYuQE7dp53Q
+Kgyq5NiEXzK4+6IRtOu55Znz1Raai6hRU6/xb0Q2wqu7wgOSu8OfsQM9lgVgSnF
Ck0/yt7T06e+ucz27EKBl2/RERTO6MmmMLOn4jv7lQRcInMH1DRCwP+V/3uD5yVX
+8vLA1vL7Z1Xym1Ei/odLqYqOsuO/fVIjbBEwk3qpQUonAdbPBR6PlTDTTfQ4TVB
seqeJC0NtL27/aR025NmCnrYf03K0sWm8F7uPVrcy/BOfE//r3oyZNUmpp5VhJ5h
7zX1G78i2Eo3neGnUB4ARtVDvouYdsWUq64mZ3M2AiCwrTzLdU/Z7Xig8yoTTbtg
TmIsugVvxHY/BSuf6TMKhJhdcbtdPkGKG5Ok7UbkGV0yF+M3nqNzpXRuZtLBx0Hw
+CdT0fNJPcKCB5SEckmtvJkuMt6U4ucUD6k7TNlOX8uBCBnvQDhlZKc+DjRanKsy
cPXzZtFElssj3h0sAzo1Y5JBQjKYZe48m/Hy+mmGP/KWeLYVjcebEYgQb+oh0KIh
jmN8NaoPXUoYVzsz3Ub01SLVkAbadS9HAmh41qWcomNDpeCc1exesuMYe8q9CGTF
kZxW7GIulfMn8Ielzo4nZGktP3Nof00j3dvadGFjee+PbyTBvMtu/kuY5saoIWNh
Pmuwug7ldtprf1cKELWR9O4jAgbRwdX76zYJNjVtu+BLiBCQLsGLKRGxqhYUCcuH
xKuTZ/m9Hcbw53O1yZGtFqKhaVyCmi9oCa0ErZ7giaSySlTGqeQ+N5aMgteNNBN4
H5GwgXZPb/C8GUu5ti2km+kvssITKzKg2zsJcIna+yrydnyNdmPfjP8N2OdZq/MR
gVuCXcelHhSwFsVe9sBPkrmrLZW9EyxeBR5aiDi5OHKPL8FSiUUbU5K1qCrbOu5M
8QWkTPdF0C3NfiwC3zN4kDVJ5KdK9m2KNfqJ7h99LrGSOk/YO9kPfAypTYf3NqfO
Ez7rNFhOnFEQOPVfz2rdKCBLLjhIBTSIECEksx+heyHJaAG7DFzBC2kLSBegZMO+
5gF8yrk6oubYA1Ku1zgyoa8ZPqp+6aPrgidhK+dkSIo4+TkY9ijzmmqLytSQO/wy
7/8TINgnZ/Z/RvxrY/xUNttLEo2YWM5GSg9VMKqctpAa2uramoflj3T2i89Jslk1
tFFQOZ1z8aWocceAIp5+hswqO5uJ+CEARBm6jzGB8RSFy4+Vu1nhljSsOiGmSRVR
jmjDNXam7whYm8MtD4BFIweJGRGorEIoO9cPOnX/YuMx8tmlqD2kIybwPwRMuEXA
yVBj5J/d0ODOD0STSmpWdFN7uNPzKSsQYLLY5x2ZV8SqFs/EVWfOPCN6VpRKpvQS
EZOkfyzPUhJ12lmBw7VnwDaxAmvn2VMZokHrNNnohFHpvMTMVSW2Ii+uxNTEwDY4
/LzhnbfMZ+50ElMMO6QOz/ANohDnwVS3pLdGume3f/xkH0gUQ34MT0QRIIgu0RRm
CO7BuJEvILp/XWEd2xkSDRKUM1fyjIWCqVlZlI4y6eAEvLDo0BljA2VY38cKdvqE
V8/MxZTwzyex+fHHkYSE9RdeS+LM31WcV82r1WCAtpYrjqE5wYmanZDscCdXDqOj
aq1frtYwmNK079+CJUGCjx6Ur8aK7RGg5VT/40hoGlCLlRuJ1eDFktAVxJ2e6bjk
jjxu7ok9FSlaWDeyf7k1uUpIisSqp4Ig64VjLFtTIeF2z7tepDFBWkHcbNHcyf9w
UzI5G6IbEIGfMBU0GqUAoY4iobf7t0PTAu00m+z2mA7oaccVfXzHxN7AqiOW56XB
rCcb66AIcPRFzm3Du4Hr/boDN17OKTgOua6OAxs/S16ZdgFJgw4CAyQPy9UmFYUe
Lu+Gb+DlCgzvQqKoIATfRK5G+o85lcig2C349eNapQjoJutwEemqpcIjAzYDF78i
GE94Ttf2RxBSJcdSi8e1tz+pyn9wN+JubcvYx4Eq/Dy5mjh1OW1O5ZLSAwoqsqgr
1dwEnziy9ak1L7SFwT+85HXXt1iOCwy6igD7FasFxW+MKMJjE41g8GXEKwZ8VguY
5rBNpg+NcyPs3efqv6jo0WLAQAAu+GpUvXN/DNwmD/I5N5iC/i3k/ndVKsfUMTme
uryWQiKRTiBpcOxrCkzX9relFsj2NL5ryXaUTTp5lTxvasG4ADtu9dk4/uMdkBC9
AC6/OVmsgJ+GZnSioIFkVf7yInq7PWY23snpBTduYcNInHwaPcR1Lull8O0f3F8A
g4vo+2K+E0nyt5skuMXsLiSthRp9blDKlTJYWH6S2+p5k7T+kMRENsMCDCjJjlyp
VunHDMLqOMEOBh8dUFXBWXhvWhlW/r/ncoHD1zXpHBkOgY3vMDa9NIfbGsT4j7Pd
1HH82qC1VoPVz56PA6GzMaMbsAPeZ1ZhbcgI/0POGCQ+hA0iRVLbXMpcvzeWDmtY
AKoLUPRokbmraTbtV1MFeCXZPa2o9YG45hxee3scrdkcvTLIRwzglwJJHGnmkxs3
BL1ojydTsrl2gXgH5gQ4YmwFN+H7NvOjY9TSHqYdnUnA9DrjshGJdLcBInKezuiO
mBa7xGjE/eRYwlp3Zft069mC94KPI06hBhj/7U2t2WPbUchweJLCoepKf6RJiMFK
Kg+7H3tWU5eC+UoToCykucGwmu8mT64OmCYcGE5H5Ect0v8uhEtzaxYg96qZBFY8
UwOxWOd4tF7ewrMdeRHW1LenXEkv7CuiFhS7XGPSBHy7oTDB1ZtWlzMjJkgWP5uF
RqDaoFsRy8LqS84SdZX7AhjCQYuh4DqYv1C51eKotecBiei42afFm7LldAk3bQ4/
gwZNVmUiufn5OqTh2IQTXxKW6f941VT4AZmpV3EaWSh+EMRId1GGo764OIyqzrxv
lLlzRjgw26ah99dCrqVG4SWgiBpucuz+CLUOZEwXZ2X6yffhQYt0BIuZt7h1K/St
ZNRPZRGvnkxGmDYiSbL3SVwl2UPKNZ+wtAIPxg70divvnPJkgB/IC099tXNyC6Ap
3svJ1aatYi30Zk4LqwgdCycDAY71v68ZbfqyncQWFooa6RBQZ6+t97A8WSpxPYGW
pFefSqyAsSpVr44XojMxkccfPhJRgYdeVzxlBOyjS+BoStCXMW6qwptCLVUMd5F3
EJyQP3MgbrBqEMlJrk8kLaIIxH9DUjhN+ARcYzWxqok+dI6q7D0or6Es66PwvHUc
+5VcEHcuv377wi3XU9lcTF4zHecN8HronfurOmxxOP6IwiNzsP9YeYBj7Gam86Xn
L+a/LI1gyFIqcGHZSbZwYrzDTMOXv+A+afkC5Uu8zaRqzKMC3+SSHOk3LvMTwrew
t8tse4lLdIgH1aCwK0/DPMUYVTTqZuJJpOd3zNARW+2RRgEQP0WnvjIwR9kLVRm3
W+PfcRJt227n3TpwuHXF++AoO7PK05uSX6LN+HmAGCVKgJJsrzdDP4sC5wYVE/Ct
HDj5Xy2wp09y5ffFIyIasVZNMVrQwahf5cxvNQUM7L6abhdnbjUNaJVpXb3K7X3D
6IiHEI/qI8Ayv7dsmBighadNRa4Dq7oUtGlLIWOdGL5gPrnyiOiFtluFmN0seonX
Hl2BNDKDxodzPFtDDZMFiIMFfMQiCvoixFSTxTNsht5Y0mUVr96HzVwv/xlhp3vL
iKDFrsIL0LJS9Q0zEk+kGfigpr836iv+Wx+WvmgqzAndsbZ6CyztVsffFm78h39d
P5LSSmozlRR9meXaKSkhFtXPgKTvMK6pW0YpJuo9uIlQ10YHdzQdUSjXDfxjYBci
V6YCMyXb1vwidYoUWTfGx7J3/hYMW3YfQ3WSTLtIw4AXKb4lRsMS3y/Gc3nmQgkx
lP5E2ynL69mDKHj1+GCUBQ/UAF5vL/wv8cqGD8iilz5sanu6cKOew55+wmNhUNXG
+oRDOV+VPbZRBUbq5ou3/UFOTL8KqGKOdOa345E+oo/qC3WvD7mohCxbhqLFl/z/
9SbcmcWiKyMphGYM0I5pjb8IFE09s4TNllt0ovyaBbUQM2uvdMniVnvcqOoxYmVz
0LZafE3wQMG5wQL8jnxggFd8ajF+ojTBc0Ae3vAipL8ncqbRhqtVRkzvM7Juawk6
B8vHGEnorxFloWr4f5OBXGHwvgxVOZufcfEXoki10hLPdKOxj2yIJ+6R6fVJM3JZ
5+TWZoAN0QcFYWWCFQ1FDdv+DvEC6qwxqgQTNF+SudzLq4nC++F+lCPumKtXsUGA
DGWJQVTKLKtd5UeytRlIkKcYQzkaqlUxQxpxWBaxj+zth+Nn1M4/ZqFqXF5VBBjH
Q5pGU9/G2fcXV4dALSX9c4U2SBDcgaMOLs51t9Jp5P8rra1VFhrxToQms/py2IIn
o9QyBnB10JeKA5zRu4kovy8EZieVhmuKyPmH2mmMOugxmu7w0dqQdTHgEssjv3GX
owUjvRrfIU4bGKmcHHvZc338ibq86XmLbZUkdRlpy0yslSfkMzZiInAWyqhL+HD1
rObopFRG5tshdfyK8cO4lxHoftws97+XbqJvcaJ/rJ7NKsjMytl5ia+N2kXQvdAC
j0bbJV/oOc9T+F/TyZrmspAkfQ8nC8v4h2juUC4CfQrmMFM8w94b8jY2+TVtGySG
BZtlRn2qeSHPf8C6Mj3AUna80xSxQgqkzH+urFlSa1i7nRFQDYLEe4xzzXE2XY5c
h2kGL5LXifAr9tI/8kdO8L9XQsJMnjHf4Ni+b7DCSbKDzgptpdtbPK9BD9j+ojU7
8lj9vH7aAt6lbsCrkDiliu/LBE4zl9NA5cZggV+n4If0g1GsXep17eXOkv6hSpo5
Tu9STAgkarZVqPoV6CQGnzMPKOHaQuKx1t1fR6cFrwiHYorXlSynjDcZPWz07vyb
lUBe0N3FB7I6+/fT8OPknlblB/khh4X3sUW6FrIVdaOLJWNixu75no66MHxCa8hs
VTsFIo59AbYOyoVX0rfT42NoP0fnIIuP4peikMOYU8wMM8NPlggF+OZsDHv4NBue
2rWEHSO6C1bXDzJRfZaKswcL9yWJI3aw8JHuC6/1EPXSEa11trtBfS0VJ+0fI6T2
2FFySVjE2zwWPP5JxQfRQWvgB7ZKewJdpVSvH31OJcF/Oz4+KpQTvlyupCvoB9Id
S7nWLDXqyqIfPix7JB/BwTPAq8Es+0veTp60oo1eZI1egtwsgx+7zNQisGOi+Zkh
zhfEOM+yE6T/QOlIm6AudPVunHgFpHqAoToO112RaW5BvNJ3EI0PSpN4NIo7DVxi
9wdcurE2n9x7Wyh9WMfDfiRZ+H1UUD8RZMuOLx48/yvrdEl4vqITNbTVl+R9A6iT
6JfaNLhvPP5eGMYLb5LsmdWmemtQBxYcqmws3omGDIkxkuvFMuOPiu9+C+hhvgOK
wnDI8mdr5SKjUAioRtt1+c0QmIi+r/v3t8tcekEXdaX/0F1dlP8VIQwLF22sgjLq
J6YlBa4ghNNWXPeU5QOcjfkmefqa7u+qZbUqRjYyRQzrDHV547dd20F8ctkSdn5a
nWdCPfMtpJn029kzUUE9jqIEFb2KUEhcACviSnG+Q569g5IVy1GhBEbw2RvbGWDy
4wDv4KY33JYidfhMHnPvvpNb7q4M8d+MIIWdsJwORcSwkmZ9DDqcSra18n6qZoyQ
ULl9DtsmH+YdoyTy9GapDbDFlknkk0ZcJy3L+ZCkG64sLyqX5U5FzaRgO6eFYdOc
IqQbj11EpRG+A48hD36OLktqyDOVxw9E7Pw21wIhfUnF1zC+PQU5jE7f4OiLhzR+
6n0mbH97onSpdiNFtAowaSLRVVPcAztjdXPixD02xAqm5go+FsrvYptMtTdnArcW
UglcrHO8AR2jNOgORAfYDjVJ9Higd43T53h9SioB5BbL0bHo8fPFO/dkhtzuV4y4
V8NmioRAZPoA9Svc5jkKaTevVxWylqnneYsIYc5aCOC0CtnGZa4up8IcWY1q4wZf
ehNrvtag9ReQJ09uAvuYjlS2BhY+Ho9N9qRbrJtVemfoUNO7TKK/9fH5ZrBEnR9L
y6wdQ4vHZWcRgI+wgJ91Vu4NjNgff0vyCuUnx6nNsbhRTkyVfd9sdLcWUdclkpkY
ZZdksJBU+fcu7hgg0eUNmh8s6vVM2XRlISuTKKOqWRkOSlU9IcJrCsQDy04rLDPc
llFW3qaDpqlyERNJJrAmbKI6aG4nzEghdst0DhSo9J27EnjMCQjV+zGK+dq9PLXE
B1EgOQt9pBC4rdusB3Ona4ohaD+oFZryV1LyyRx7SyUqfdoaly02fwRq6MNAFqI7
T6frayyWmZcKrb+x9S7Mq8hIySpKKawul2sh1nP/4VTKyW/5LU6UhG/Hbsz606bm
Ro3sj0MNxg5zti4Szt1a/tq69z8hgg0/ewyFlz51ObBcuiSwrh17fYZOe+c3vOSL
k2dsTtraTSKvCi1x8lMTS19I9XV0q8LLeMOFltKbPc1zpfqWLW6oXcJBRomVrk88
3LKenvtUyKYfBceRZNvRbJ7XYMex5Cp5ENCnrMIPdFutKva2Dwo+PVhzVdebgHex
rhCWJm8Ev4TrAS0QPg7NzwWzb1rKITYcbeXwpGnD3JlTTCXX2TxPKw82/sfNBZP+
PzJ4eDeOyLKsaz/WxWl8rjKh2/n3e/OUu67nymUF/lMbD+0YxUAmr9GO1+g0aDi8
1pnt/iVnLoJX4nOfH1GS+h7dWje8E20GPLZXGYgv60bmrTRk8PV4hZXLTbqWL7lQ
1oxELRDOP1abhT2nUOlyVH9U5+JeYHYdjRjxE5lPlYjp50aF1SNlbE8QlObAIDHh
i3CO7i2ZxyBkYadljUN58R1eUj6kEF9ndyi0qQ+r+S/JFEUPOkefJND4yL1j/u5+
9zBkPwC+6y18u4P7pks5HpbLcbvDr8rgeg6trzMgBJjVx8hBXdAQ6/afn1bc6zbg
H2n4dookyw1hFMjhZphLEJALaYFw35k/xnZnETPgnuMVNV4UA3/1VKwLflj4UjGF
9j1U9tv7f/1Z81QCE4sA3OC1X1FuK9+ST6uAHTlcHIY1OzDVnAuvpiWLqlIsd/xt
chYmWY3J5O3lBiSXwk/7X3SYzY4x7KrnAAPohCD6TgMzp1nRKtpGoQRxwAs9xWDg
C/WtRhcSqHhe0o74BZd22mWIIPa3xsYv3nCDH6NVrix+86Sc194yFiECGL+PbsJ5
HlWwloCl13iCm1+aavYWxfaIZVz3LS690QMwXY6apfWxcQhNj9rXvbo+vpJ8RWJP
rfYTWuZ4KeLCbKWFo0NdSpfIEfbyzGH+3J3ZjdkeWPt7bfERQGmM/XuPEKOsyvka
b8idl6JhzAIoUGLEVg7iErxDjFl1L4OZkUvpYs/wEC9q7HpvaO8wp262dj6af/Ir
OA8NOvgLv/kV1W8a1zN/rBAGWBf55QCorbrcQA/W/dBac135RLZvoWNpevx+mKF0
VQHvljlQkx9/nqavd5z9fuLjqdvqKoH4c6Y1RAgWsnlO5YicSjeGr6Mt/CNPH/0I
JwLjpxxpoQ4ucptEZIqTcEtbdIYWiLqqsZJ0Zq/1w4z8xKZNiOSxC6BAONz7wzo5
45o+hFUHlbSRh3ZDhi7rCTVy2DtzH8UAcHTqE3IQq2mNrjOiMJSpG91c+xkeH7Um
JyzUUrwko06/AycoX1KLzLmjOl+2zZtjMEsgvBSDCAO99ejgEeW/6QUtW/xXoj4G
LKOCF1/8eq82xBN79V1EI8LkiOSMe+De14zdmt0LXR3ZBwZHA6O2INcMvSIgO2Xx
C/3WqrZPIjB52R9a4PFZK8WJ6R3yuDlY2D7snS/ob/PWxQuURQH+xeK0+B6ljCYr
xPbqN3Kiu2K84Pz+Er7ySECcxwaXZnid0LBszoe84s50RvovtJByPtO1oOvWxVV/
VsH82pZ1peaMp1TAfDm4L5EOAn6AtMwIyUNB1P2mBSIPekTIuESayqk777zABwnZ
bOf08/jFLcBou/4rjaxkDoywlVcDgT7IAGJurPUiOoGliPa0+qlho1b6aW3knqQV
u3TC8kHNdiZbbJ0aRqgvjsfoChENZLAeOYPNrURIaXng+shUCj6deq/d55djCS6e
99cvxVkgn0KLWa43sHsvVGBVNtzRk6NeZe7NcME1+Z2yCxPYmPUg6ozNfzAprXmE
faO4CMsU+Gb3XoHi0rmKIqsrjjmdjRZkhBjOPnn/a1nwQ9zPyIgpY9QRNiJFoI1c
NtViqRwoOgRbKs/JA2f9i8eVF8hSoic0EItklMk63CxDUPmxKOQzAM/aUwndUzqB
ZkoUZOBPP6pQ8l58os//Va0OdZPW6xRm0cQwvtAmQROhHg5+qdS/5JCRktJJ1DdT
8HZ4mv0Q7ysxtzz5myw0gvRS4nVmFdqJQtPyFw4vwL6nowsbdkY5TChYnwJG5LJq
tSDt+kUNX+UjLd80ktBR1kqPBhPbM+vBLjk2Rv4NLR6SruOZ0kq5+ZQo+MPKGbt+
XYC1niH3jlGGcjUma1ezVmeCudjSTLLcWFORI9V7Yn+0IMIBrLxPRnNwIjdCS1Rj
Yii3nullnhEjNuH8jmhu/0CQ5AEBxspYj/nEj+Pty/n1LSNJG7YqkIX4fH7MlvCI
lfnP4ceAOq76VRJo45qdD2Eme0EUxSNJYHcoGay+tUbjv+274ftotPzY0F8yqGu8
klwyiRDx98ps0/vMqEITkAwqyKvlyQZezshBCVbsras1arbdyNMFY27gLX3n+xlv
Dfdhag3nssyV0KyEoCryCs6iULLmd5TX0VbdKpkIfIxYLMx/dPAyST51OMKmJb4y
TKZDpesjEB52AE+obBvpOMejVMNwM1E/BVW90ZtCqaHvY82D+j7jVkdp857GEzCb
iaNZPMYKyQaJ70N21w2aMvCi7uvhBLyqTziT1iDXsk4qq8LpRw7neRMUxGPH/xUK
SKA3saRuhGCND+AQWqh6S6ieTwIZdDuqVb6mpxgvgb1zShbpesRQxtDti9aXVhRf
gfCoPkiAvu5ptFJ2R4S8LkTdRVJidSfPlKSF832+TaV891uLPTF/ih8pYV5RUXdM
1kxE4W0cWegj5GDYXZMB4poC5/clDTeHfY6XTjd2Y1dfuLDbrHACG4zdQ1+CPEg7
s83DNBCNfcEW7b2icDy9BbV15h+mgFpx3LyQ4ijr0Kgl4tFnXEiQOO27X5C4jOh7
ClV76Qq9Uj1x+sw1ImHs4mWAfkuCoJ4GyPke+i2Y6I0yjA3bUgnQkSMoraTuRDJw
udG8mcvrgrRN6Wx1nfxYAeSXuv2nLnTkcRU/zuzsvam9I94hHcZQca09BUxum3tA
4WpyObXR+rnh1JEMwVRgV+OKrDN2b7pGuHlkloWUjD/uw9AGB5SVHeyzbsvKh/Vf
T85EeIrXsw7k8q1NgvnLVb9Gtz9hJhCQpHdTIa8ssnRYS0Ic2vRKk4hK7TScae9J
j133nM8b8lRc1VxDhbLXk8KdFhH9Ux523oCdI79RDX9OLNt8NQPMJSNmh5oUI3nl
7JaGx9OrfIWv8ve4MtLZG4JrrEH17CF+ratUYxLavk5WE3KsZas+dHaNIdTYd2Kt
s5Uj1YTS6wxt8L5meDypjoLXdBI4rzjUMArGRS1M8zBmCbzKfwU8kICaq4DvlkJH
wsg1Yh05IYpo5Aw1UafnGSfbUD4hseUImDq1pIxGM0i3p4D4xz7GxViXlosMLpXS
KjrAMQvxRH4bglEB5TyCkPOsDVxjMP9bObFzquYxWyu85xsHzivViq3XuUrL8jhe
n0QElugDhISolZlEZTi/X2dYCvBsogi1yt7zUGquxFLjTNKXfcmfCZ0MT7vAbEGY
OtdlKyrIfsGVnHduWBZhDOLmL/8ShBy5N/KT75ABirRFpoG1ryWWqLnsugLfV2cV
S0PuzYBnbEO7E23Xc3LS6FwpO0ZNcpBZUxJYX0/LQyG2yb7R5E3I+T05GKrXu5Qm
wpQaFGMaFA9vg2fFvjc4hkINv3vIRJYxR7r0xnFvCSuteSyIJzl9jPEf2gSt65IH
HapuZIozYKeSCnb5lD+1iFfxj+vwJkMAEGNtinjf16TIKxToVXYnRderCilmQbT5
qT7q2NWu1lRYQfGr5UuNWGE5bjXciCJZY1mcxhAm+3/U8Cz7qsEO7+Go95OsXM7E
Yx+w3q4+DOrUhlANVugc/cL0oqhhFJivjDYqGe2IE7hmqC7bzPlx+f3cwtBa+GnQ
BNW9Tnky9f1936zv3O6hL11T7j3dDq8cicPZePObJZn3+z2vYr/IXwHB2D2hCazS
k/bfpmuylT3FcoqCyXkwGoPJeVlL3YbkMaHL3Lgs5THr8ZppNLBQVR8oxZ0R7RHb
KBMK7g3O1dFmraXhfnnVO5RShBAYLU8Cbgq/MqPQJlMAyNrDvmEo1bBz70qGP1jR
rZjzCje3Mav+yb5ggLYEvPbmKUGeDlka7A7jb5JhaNNnJHWfnyBjQh+JHXNQ0cX4
xwo+dIz2C+kcIZtxUZsqso2XyGG37aboehzvqAiv6ILOq38X36hmzgBo2vgi62iY
n1nS+emqsCWXuzsGE3Svklyu5uvzhRO+uzMI9ObbMrvQEVE3ew/1WTyohUslFXFV
N05xIWcOilj0rP0mLKjePNqsT9lEyRqPMyRq1tQcAlAtTVHEi+gG/BbFLRocZYLK
ZTT0tPEQ0vk4exJxqOMn2QEOPa/EGYAvB7hRUGncU2Ad+1Yu7u8Tu0RYO5MjSqF9
3XMq4dJ8sh822WZJgtQqfAPEd1ybSVc3BG1CW0KtVqhmuvO08PXFl7aBuw3SNA/f
/3ajutXzbHZ7EvvMF3VpQLkGe1PMu7sZIrmLrqKNDvUIAbnNBE9nTicZTnZcOQVd
bBA0b+rjz76MjzNppkdrc2QV+BZEwAQO6a+O/OTmGDd9pnDnxkeieys8w1zrCcYn
AmAUzU4EPjq480aGt4xoftUM5FqW7XZQkZ3Sn4PTyG1ynd4FF8sA7VpBlA9ydUFF
sqc1DNXUYgODl4/Z8x9Sv9PqNw/IdOl9DelsHQ9k73S/Dz6ho+WqWdov8XQ9HB88
CgkfVzkgSOMsSF++ITo0MFB5BT5LxAOtPyXD7o3Cluh8j5FoUelY+Y8A43yO40y5
SOc995C+4iEIe8UtlkRRrS+IN6eNPlu30F8dty1sPbFpQ5VsN6iJWXZ17GQANVc3
UVtJExksQow+VNHUkOJ7W221aFcys5qRCUxfgvRsLOOWRswnZSu9/NZnRUz00c2C
K2Flb9WLreLGoNBHKLTA1XUbNngPr3/oOSO1/tY8vqoZeZQf5DyYvlAZ5zwiaEEF
LYmETni2Md0Vr/sn6zTQ4Wime/VrvNz4PV5SCcIr0kLXIhBZLFdEWSEbu0DIFp9A
yU8KkLiEQOD37vXRfmm+B3ZF0zbHgIe0a0xtsl/tleXtPcZLs3q2W6IeSiMmCtnc
8V1SzEdBm8Vk1wBMlElu9RaT1U43SrTIJzBPEEKLRB2cqlDd7efDSli7nMC/XcP7
7U25NDob8/wcx7fThm5HeY7yhR2+2D9eUiW+BjrfuKaeq3PMckEfOOAEYBt8jB6N
khS+lRphlvaGuI2AefalasRVUFe0zsuVIvhNWvFEpradgsNUvBiXp3l63dAV2K9E
AQx7ALZxIgFgSidQoBrORgpDtPyhcK7kvloNM5PPQ7y64IsL+iJAbxR2cS3P0ck6
fi+USKMCsLIpW8DFqs7akQd90/PtBOJ4MmFlsS13EXgaSgvtpVSVhwKHvn5CJVGm
2LEV2oJZILjbOOB7gvjwL703AsblNFGFngjwUrXAN9s7B7RqQMQcZNvM7EzhgVdV
39wjTaAgqtBgeIh90KKGz3lDNf6Lcf8pACQ7SFInR6BURea8AZrRDq6sIXyu+bZh
ITfhKX7xYtxBpg3jRfzZ6ocT5ufq0BbdbQ6daq/aYLj361rp1WbKBBoYIIVsKGS7
m0Cz6IuoSL0odw1F/PzA6vAnuraDM9tz+kNpk8akhozoL/SetlUlEQLBxBhgS7cu
gc7ohRrWK7eZiM2vUSUIfE6qVBuLLTo2PYA1quybQfWEyDjri2PzXy5JixG/gelA
S6N6lU3LTl1SCgGqUkKIrQ094aty7xITXRNiVYYkVrEYSny9zWD8q7nqeVtOjeUZ
3oZerty1wYx8DGII2XgWRUZCIYyv5mrZyZjVE6n0MV+C5z2K6eJVvWDChcGC31kW
ELuxOZcW4RUf5RZ5luOv1qTBbja1IAcyNGt3FUoyh7sEFL0Vf4V9p02FRT8Rb4ym
IHDg80lkR8/bwC+1Zt7MH7vO0Fy+vE12erUW8IluHXTzCAdZxU4PCSWlLQLTdLxL
27dOS2XUpyRMSgZov+RHnddV45JCOTsncx1n87VXSlIQLjSeVDiGX52lID9CqE7b
we6W4U0w9c0iA3y+IUspnRwvK5tZ/ZjM4f97UjlqBGUhWxys7Uz8xH3SN0Rx4xag
0qEdvOcr8c0+dfXQNofle4TVa5wERRnYpiz1vSwojTZHOUuRjAA59igGGQBaLPBw
Yg8fr/shOxSM2nyk07Lyp+i5grBU3bqefBqnZBGYW0E1VnZMeC7jP0Z9QPX8zfWt
XYTp8DinEiODvOx41hFS1Z8bHvuYHUwbs1prG7Nyr4qqkSbry4ZDEGr1PGKknLA5
DHTw59pQtHuxTIFfzHdLx06ZcRP+DhxAfgMlhxwOym/UDlxvVfUngcdoRs8FnDYx
jLSA1qGs39jbM8e4lIUmfSDg3x+PqZL5N7wVePoV9tihrL6HKLkdVrfGj4VQi9jM
kzsZZF+1vWUqBw+EY2zlt3dXdv85dOEWQIwu7hwFPEOPuMkTJvb524GP0SPKegzH
40Yv4sW/lLeREMuuIlp6PSSoUiBKYr75i/P7B4M9d7CRur3gL6jx0ogw/Km8TS37
XDU8zTaU820hL+G5jsUPYx3pRFIUKJCM7kFongO9Cn82WdcOdUs96h/kQ1sDw605
/5gDZxD7t2eMgHz9MdBp4zI3gWCC7EuoO0MkHGhuSI/pU90HjDQcFpBb1Z1rSLgN
nIfwgwfmkdkJ+4z423yHH8dpxbO5+NoF/AXQvoV2cxFDBsOJQLp7jMNwZAZOvMHs
cParkoTroSZgGNoEdj6hX0c495kiH1qU+wXCrYvynLb+UkBcAC9ST+U1IyARNZ+v
G23P7sgsfD2B+LGliGIWKnM2wvGSqTio3rqPXegO3eJQ+LmmMc1lMnYuywXXV3yn
bNBMk38mQwjaaztolcp72NnpUcrdYdr3+7IHFfk/Q2q7LsQ+cueb6dTOICdNeQJp
QAswqkcNzrPVKsCJHCprw5cNnNZqFxur6zdNWjfnIuq+N8LOayVE0tO7dleyQ+f8
OYpeMr+Qqc7ypBdnLvvhRPpFMMiF11jdysTYXRgaVGPOgPZQdViie1f1jhxCfd9d
M//dbd46j4Gjv1OIfz8o5DJR+ovW5GdEE0IphVCkxDh0UXSr8QcJocUqRfitOU+K
QITg64lF4/tQsDiG/WEWSCIcbrjKZNnbYdAkBEZ43rrC+s6rX7cXE8QSMy4bUuO7
UBwgEOheaqw6LI+x1R3MCC313Juc87I00LkPBoyvnxveaWUgG+FPgP5Ttck2Fqe2
8+9qsq8CVrLDTb22mn1JQH2yE177WufjkK6tLDW9n+ZipQ7yF5JnuKMCUk3ldY9G
l0fnNVZq8ZNyPnUf5biCO6akMPpYbtpNPvX8SUCvKhSwE539rR7SJ4syBpsamvAt
x5TKobWIQO90F6IGzckXuFVgEgUFPgHmIZZimeifW+XNoH2oh/4eB6HrCHDqchTK
PDndkNFLhK7p3/xdNRGsckvedu0np3FaByBIhc8E3c6NGdd79zGAh8YwjRaDVotb
5jbbKBipp2d7aQk1M1LtowyUyd3+tNEM4vyCnIL6KcJZgkVU4z6vg6tKySwZosSJ
6LwrZAnr3eKx/UImZgXeuMwvWREIm+2wIGrpY1DDY+BXhoVMgdqfgnkJSiCGYy/N
+ApZZ1GTSqBDYXMCPzC1qZBKMzRhHmNjEAbtrA0BITC8Wwgxlez6JdtyPQIfniNR
Urd3BVnqkZGupATiJfSmWWP971VYyUzQwQeh/1QYU/27jBLM81e3ld7nvCXe7D/o
KPSMjh3OZzAnzVAzF7qLJ3HXQ9AOW6Dj81N+VgMbMn5pI6VkXqnIR89Dj99zF8xW
lvd0VLGeHo7w06yLp9J1q5idhiVd1swL5X/SUB8f9QAPXFhD8WXmjawmSkzttk7V
/eTmAg1hZ1oddCWhkxY7SuPCM/VnqBTho4trKNdJSJ+2G0IMMzRjYTB8Gtua3ypv
EMtI+9LwxWseNXAO6mcYoUb5jdMI/Nf4ll4FNz9J0V9VF8w1NOxcKzprMbIglYoL
xfgnKC21QYp6JIu/mU7JZVDAQ+K5+CwJ/sLQ0KH0/NE3Se35pPpq8vxhbLYm07Xz
B5nei7reDT9lUszfl3sIuvjuZP3lFYAccq/ytWWGnOm6K18jqpbUUYRQrhY09LVc
oriDTSold2C6p+r9+jT9aVqUg9KB7aHXM6GfDLD+UoEDdlE/d6t+eTZLR+gf471T
axRgE/JZL4AAbyOZQdoHFTaPIdLKI90EFagE3eNPSIRohfiJiRw5M934KjT0Lmyj
lRwNaclDRCpNkmwIOXHTwjnayUf03uvAVdAc4nNzBFzOkSwYis37EFY70KoZ3LFr
VukK71FgYdAPyz5cYgd1VSB0v47bwc5RS6f9QeHH0D50LwCGDOi+234/IhD/34e5
NZ/WjX6DLpBX9eTp/mpratezFM10t/swUrdMnPqxDJdadtERVz+2lkJuW5/XOCVx
qu7r0iePKDSKP86SEFT2Ig6+MwnhCn3Opd1qwrozKNRJGhMZOgLLQOIRvOY+kRS6
h3FiFRr8OpYQialbCrFpS7v2NFwRgeaNkpcqDwZ7GnCBEXvED8O8PqwaAF8JVsNo
8wwXe92HCNKkKVhhZkxPhTLRiVrNh8zjpjl0W7ZxKLe30BMjQ2a7ZL/nUJO7vaSu
FqBbT5jRSOkYYrAmZ4Ut9GT+lq5xt/U4smmrR1pVv1Lw2Wpgr++/Ecpy4wA/RTDL
Z7CFDis6HbN6vktZ7PZB+ebDKjuK9zmdzZVfoKUmoIdXicd7kq+1+bIuRPlG2YHO
FU7joH6dPgLcBEJJ1bHS3pSuekCrDrMRqqmm+1fRw7BSK4JIKfotrN5Oa/6GKOod
xUfPT7Un4m9tybYq6do9KiE8aMIDIGb1FfvuFf8kxyWMsIEyLcoktsolGaI7NxHT
tql3SDEYiIJjg9aL1N7BwSHCHGf6n4bNHpBYme2WUF8oQctRWLehzasgC9V6PD0m
GNgTt74xUrVPUWaDacfIr4FAGERTArVh2iFr9oe4y8/UC7wb2iLfNIXvaLpVttKH
tk2cl1K/GXY+zCk+swGS3Xu01e1eFOwIqjfmdoCLatCOmcpj4Z/N2K9p2a5FQ1O5
Lg/tG2fmePRZmBcstZp6gOz0tpmGLc5FFGzwg4HJcdURFnpyshydS4NdA+I1/eBi
RGrprYh5BIej8HeOoZc0B8K34IE3aqidNcPdOb73csd37R3ySvlYCz2XmKZfrPfw
peMYkH9JM/8b8l21OHVcByrwt4UeuHHU1sDcDSXj1Nlmpe9fpT6uzQWicrw4I0vo
sYu9V5Cm3ieX0lyoS0Ui+fQ6aEAph4UgABOfIwDpTZzy3lRseAqRgYvZo46z0vGv
Q2xhsFFO8XTgg3JK6n5b6IkRwgKwgTx22Y073SI6unTge+xzFH00KiqtGqG2gdgR
7IEAp6E2PymdkiRbVyZkgfwDZGfnydrLPoRhC20TzMCwB7WcBdTA8psYDPgbkODE
FjbbpVlkRWqxeAVkBcnE5xlDp2nJKa54Xnyl2NeWY8F1H2RcR+3xVOq9oozA51wi
Pfkilqkug9ziT4yNUoS+/avfrm/QjqNYfGnJfv8mXQYGYcM4WJbvebvzoSZ568C6
nlRG3E0Tqpkflx4WKYN8+3CDPUYHImRwvJ+LO+YnVKxc591waumL1vkGBBF/IFp4
00FMGB+4G8jQdEUbQ93gUbJqGzwg1Fefv9kwM4Icj0Ta3B0qLamfgDBRUfS8s+gb
jupe5RxWgattOhvvdDZRHLeK94WYpGltJkK4EG4I3RWv8FmZn+xxW4AH3W8A+RbV
n/vyqbug//iJxSemWdpFrI+LFE/WKmhqwGW9GZ6mkoUYQL/MZSTVhFRFZj+W5ORN
baF7cLatHfIEGwyFfHLcQcu4dwJ59UwY9Hmb1+O8B+FLc7dblMz8++En/a8Yj5iY
zOiHoAfRLvK+XejLKdyrTCobiV1D9RuNMfE/RjpEwLy/vvr06CPM56jhjnHhdQNn
YMQ18kqCqcVzjTxDsCzQEpK4JOOuzUPPR1JSlCyDHlcnTdAT7nBfclb+68ja0otK
zCjvy2rHyx4f1o+HM3gIyrHAF9evliZ6x8tlUrjqfpSwxzqFzVC0UOlLWfKOFRaY
IrGWEG49l964FFceVDBI4f+u+A44DzO3dNtjQq4Utppf+/F38teIGzkxKTB/USs5
wRJnSXPpUsYXIi+lJkDk2gDknJTpdRV2oyRsLPzl+TG0jmvN198Rfv5ZQ4tQ2r/k
BPq0/OkqM/KFcnInkDVwP3+aw4x62G7fRp5BPAfgQ1P07gVpdwc5PkMt0xTS6lz9
IzWgzVfPuGHyVa/POWx65fihzi4f3IpKlOddkOEKcQE4ujy39fkRNswowdhFc5EV
+HYrMEF17TrQOyBBpGFj+HftaNpbNgN31DmPqQjsxDgYayCYoju06lN4zl7ks6OQ
9gUC8nhsnhVGzp6v1fPCd3g1/d30iT9V4lZFDqkgbmKi/wDTJW35lS+LdTuKryns
f25d1pI16EcS55bH0xVmBNe6qFthBFtp9sap01UvL2m/03P3xYJG0kpAIGOdgxxl
1nFh5Hag64IImbW8nGEs0qcHoXAsvNqE/zSY8TaKJOnqYnhq+wkh/aO59DLIfYVD
lM1OxyTjT8z/RbL+yO3Fx63zFPWZ1AQPR5SjxeSTi1v9ygDP3n9CogIQBPw6p+Q5
KuOTR124ODldJknV75o6slISNQJhlfxsX49j9yx5V51E4ZCFNsb6mfcwdHFQdR2c
AZRGW5zQiuOqjshhaIpvNpE4zYw0oQsKhEL4d4e2gvN32DvlcTdg5QFJ8fkr/LMx
2xRyAyNkuaDUNl4VBg8Iy6VvhDPp5P83xbImqN55rAXMDnHigMQ5W6RZwgs5zjlu
PbzGp18d/tJApbv0Vp0pvlFIa/F1yLZV4T8iGGjgSfab/guLNFdVqTcxzsJ4vYxR
HW1Zi/3i7l+kHBpE9Mq5cSObxbwBa3N3QLu9CrUqT1PsxefkhMg2ZpeiRZzDDxS+
xT1V9gf7QiA0PXnizL3QQmaKVmvtRIp5bXTunUGQ75ADJT1W6cV3Z8F7V2CS1pu8
IKJNyKAmJSreCqL0UitfWV13Qa7+OxjAk73fnvvz8K8+nVmQ2JHI3Qjja0Fp8RL0
dJAJp9CW6Sxn497X2CRMqGy6FJvytytz16ASu6gn6SXy1nossSAWSyiU57ARz4FE
7ISD0XOvXg1SGejoPP8D9d36eGVQcsM+cZcniopP1roSU2T+DWg9bO4L2DdrezG6
UdITFv+lCGs+zrNuNRXHvm/2BoMkVQrODzPmrbIUYwBfre7RIqYk32CLWcNDw93J
7stQXrPp5c+40uQ93bmuMfK7pGOFTDJCiuNYhwYAjrzXC1ilRWsDWKYl58OPPr1/
knbhdufxzaIADwpGQe4NveLeFzO7Otd1dbkA3zefdZxIoTQ+cwI5i/sx64O83fgE
zoPO3WGe9ooTfino8rIuLS4/xhjtu6W2QONfL0DwUnX9IvyRIfloi1G1xt8zExRN
EG5KL5ThSCkx2JPgDIJHGDz06rlU4/pMXqIqHe6JBzf4gFMx8mc5wXVSZpK23Ak2
n2TRQ3VT1zJLsAHbdB/nwhAJ+8cRdBRBDAFnemT6jKTHpzWmnf0eurwSqcI24yhL
KVCqRGxxuGk5/AMM7poW7Jquu8vZMc/BxFq1/DuS3lTHq+DkMu819fU0M9rxEmJ4
CLoydxSbPZ4zhietp24BFD0o//69QQD/I5dTUnT7uQbeLZ1Mes9dn/YdSSjk237u
hmNNKJkDq42nzm9nR5cXSx3rd57HG9DSS4NcGBvh9FaTtlQh8rWCrT/qXGg+Sz3v
ewsKy+vrJjZsLYPsbMgXdkAu4wsPHaGj+7L0axDKE/zXFxn77O5UpzEyEE+PA+jA
dIxEi8NfJTHXqaI0n1+3O7rp/Gp2cdh9MCovZFdC54XJh808P4005+hUqP2+vSbJ
GAHYMwc+AnGr/cesYfCIc0OFXSWrTYN9o8KBsufx0PlRfknNVM7sM/k5Nzivxm4W
WAQlPO91au4J98AxPv4A92MEOIxbkVs7k7QzQ48vwr0iC50YNC9WRs6ZRrwXnJBd
Xfm5S0fa/jvIa7DnVzVINr5p30b/T1KgeLSMm1DSqGZVR/es653GEzGmuHUAi3G3
uLxELbb6wKOF2DUPa1bhWnLkkLtCKxNtN0OjTA2pHVGXUObOE7sDdR6w72NKBMpU
cukZCaplRfrvsOuwpYYBWlncp9BGaK6fqqzhG+6IcVVrVl9HzxnKlFuSJhK1cwXe
rcPXXM/bkGzselb2tHvKHYur5Q28lrjN2C8O1XQiJmKcZjyB6t3ZhSfnUCHdw8N/
c+MU4azNDsuss+SYY3WjPA26JmMW8C7AG5RnBQmSOeRQzGeKkAERvCKORShoIQXX
ar4Cw7fOwM81B68iN8yzr9vq852LEii4iVNbsp0R4KWEF4SJfxexOMVFfYr7JfyA
MwlJzF/FiItK5ObeUfxhxwXsgI3Rn6ucqd9SU0VQD8tyltM1FR04KAPzf+IsDXd7
fQhjh4l6YN+7XbnFr4Db9jRR2DXtDERRBJIO9A4Iqg8fwKRvNfIlNnGAAGLnRS6w
tDQ5cxErX5+tEYm7iZQJfaV+4gmYW32e6KOcl68HOoxz0UfoNr5muSjaRNvSqIRr
ryyIFeJmYl0KlBOY73zqmnDKmG8UgINJf5KOo7cpGjXVaFV8kzskBDfLV4ya8G2W
A/aZ7ip2BOUJh+Q7D/tx+lmJT4tqPK4XfS8fzFh9tTkBt2plAL6CwNQhQgdVayBx
SbkK7gX7boUYmZeE5RIagShq2m9KTd2zV6MPnh3pVdNbTPeqT8ZvsE4o4OVxODD2
8dKlpX20Yry10dExD6bXbbxjFnbF0vejkKmlv+zxTv9+hmPshJYUr+lilkNuY82O
mdo8T6WaKt3DF+4nlQ45TuEFeLUdvNa0cgvFZcCWkDIhCtKZPkgV2wCnOfZbYO20
VHISzeHABfm58X3zlvjrABOJnVeZxtHk7mL9NQjBd6QoeWR5mqEu8GfUjtxgdWLJ
beyJS8+GJw3K4AYIDgY2DfIzlYdtRjrA7QYpyS1KYoMUAh5W9fR9HobPc1sTItVi
guGnctITVUrbEZNh7rrZLjH1j0/eFHqhP36VjQsg5zxucY7dpduxDFl+lnqks6tF
AooMyPL/wE1iWJA0HUSpAUfbAPWyjjn7pR+ooSx+6Lxs0a9FmzVuI0sjxgqBieDu
DYmcv4gAbVBJ/UGd+0MsZ6ti5O2CdwfvG4/d8gpQ/9q29Dd+s+dGpIsleWAe1vr7
8maOV82ixVkNS9ykbo0p4IIY3YaWSGX1tEUmCBY8rNFki+OO68sNJfIX51cATHWa
eYh6M9BA95P1S2q8urzMJMBgfXsSYtBH/DlTvAApQD4X5Fa6/j84OL0vcmivzhQb
DLgtmiNUBHqiRZFORPWAK7aJdffmnm+QZERhSgWE8T+5vH5WXqOuaRp5MeMtyg+x
rEdb+pllLgOs3Of7OnyOqAx6JA20SgUd4YMH6/WjeclLRwVc3tJTfadpqOVOnqWv
NEkDyEfec9h0LEuCPnfzcglvq05R5PDQKA+qXjd+umI0B0JHKkFCHqbBog/Q9kbF
a4V0nVQ55ds9hDD6U4JxDBLppgcI4qprrvXjmhm+mMFzUUnZuO+D/wnw2LbYQSXM
eRSh2yeGlPwf374fvrW1sptrUNmsuugo0p4RFgRzB5KUihqlsbjZVst2WIj8m6cb
CoSTcBgmJiqVNH4WQI2UAPhRmUqEQ7gOx2JOBj89aWTtKQqkH8CW3aipwjwduExP
F+lgqgwvXHe6Lt6nV9yYp02BiD8o1j+ufi+WtiZPk8rDYAm5K4nL9l2QLRFoW1j1
QkBZkdHqyVu5jKbsE1dGG7zKEYtPu7juu3Vs+9VLCPaNhqpf4kEVB1LaXyQqU90j
wcDRicY1tOtEyRqm+ZWw8J5JmO56app7x+fWkB0Dn0pcAHdD5RwmSf7KXjO7XQLx
xmdNuNkPa4bLMVNdZFjbtD+kqj3ZJqfk+ve0wWUzDTcNgbD/CuV955SFqptKyF63
tGzwypySvwYzkXYnb4shcQEk1OzNb9dTjyMyKu8Ng0ykPk/qSwcjJ7Y2xVHr0tke
WgCyKXNGV8pkzlpr2dz2JeJQlOdiSyO5cGQZJgzZya/Mxc3JR5uLgMjVP1+Lk8WV
XoR+e8aEIaBR0Fw4acxHo0j39TuwAbwljUAzdSzE+1C82La2rLhhHvrrJ2LqvkXb
c4v+xV7R7WigJ1/58Dgmqpd6PNRFTkZNDLgdu+7OThTBBC62xvyk37RrtgYpNu31
Lz1q8EUhLJ2tlrh9T31o23gPot9yJDnCcYPLKDIhic4q/Owxixfg+iaaws6NZaTt
gPVy50CDhwwbsYHvJ4mdNtJHUeLy4jVWf9bz6SxUZdygEv7W06Di7tvk+ZAqciJ9
H6cbmcOh+UTgA1cXtVpgWygeOeGbi97XO8DAwtEU+2nU95jNrGhvxt9ZeW/e5is2
FUvucQukAsZUhp4I3UkeSL98UNKTbivCb3VnXCHWdTA4FzZDA25DXKHtOybUToOj
GSO9KvJuFdq/pTtFkN/yTkrmYBvTlYxkpD+MMPSW1CKYMdVfKAWaEhPzDaDY7Upw
BqJebwVYp/0ZCL5cvpPIXdldQ+KiX5DbYndfCIah+T+5ArXQWUPNKjeLi0xIQ9dO
yJIAA3viiTxRIAtgMM7yd42+CkBo6Lh2DS88YHAxyiuRzseWExmbkVOYMykDDjqj
fFVnaAlz53Y7CnVSgF99/VZZFuVymC4dtGVPUpx2nSb54ZtYQpngruUubIfpD2E6
o3sDwBxH/bGEyADwchpanJJpLdlJGz7ChOmk0pGDzK7Z4RuQlEo4va/XL2b1y6Oj
/QmRP7x+TrDVSuDOjevipGacBMvJk64TqQitEd9WjQZ3vfd0WjR+8ElMvaNWvZec
BOTH6cvoG7ruiwKWm1aJl+hvCkaKrvx8purjiOxyhWMARwFXy27AU0lkQcaa/485
TGHOY0mYY+4NjWGzl8gk4rUpybwOIlIlAs1Bd9q0isbwXD/wVzL2qvXV64V4ptfo
eFSF73wUs1ItjgbHyT9fT8uD4zvEaRyfmBKXSbeXQ9uG6K+ikTcqDjSqCp6PenGd
HoB0lb46yQRBgn/Pqprp9TCQsElRBHlOpJg1IK4WW7uewl4uO/bUzemy/xBuZar7
x+ZT2rJtyhWtP9QmG7zSIjVtOC/wQTdlRNla3dVdQj8EStMogGc9AfFcdLieQ4We
t+6b03cD9ene6yq3zP0pW5rhrg7URFr+iZtxjBIhqv0uBxwNQ82bWrXOqMCPB0S7
hG3iwnKFAstUbumZmdzz3iQco2E6PNRGpybgsHsqpnr7f0CwtW6TTgMOcQZ+5lsR
8bnWnVWMvpB4YS0Tfz9RoddaIF/o3B444yrUY1SYjxP0zUs+aetFtZo92cnXUoBM
I7rvJ8M5yEDOzxd3yHSQKaGuZCToZkcvxlBY+GJZNuJ0PZyhjRFbFYMTOaQ+DJW2
ICSbC+lW/6XPlnz2U8KPR8tb4G4DOgbHDFZoWO+DMLq5HRgbPJV66uiT2Wp41FW/
FYigdLEQN1RpkpzKw7Zm8YA66MdjWtuvG2IbtscnCgWyE+MI6vLctzZYOMn9TaIJ
ZngLEUYX/RaxFnkfInuqiNGc9D49YvPrQGQAXv1mYptEDl/V8G8dGYz6aUE9fQ2N
RnGlUdlPaeVQALsB6FbkGK9cZMogcoopwbysScdXs1LUwD18LAEnJR3dLKo5Fz/x
GmwDSVvgRX1BJuS2r7Jucq7fGgpMmI00YNJKP9JexVR6x9Na0oc101WLsvpBjLj6
XAp02sCbDaowjPGshVHaf6Bf+H+cV9FkzRdouuLuMyeYR1e5XbhF8aGeD3bAn5SY
UaiqQhBFfmK0iy+NT7fFBnYA9YV8EDSQUTRlQqknLQLXwN+wKuswwxlTcTB6XnaR
ncubgAhPYnNxoSHsZaXdDrFRbH/FXgfvrrHvDF1xaQG9umjUqI9ie40bkeOFxtFh
DnP0Eg0pcdnGao4VU93hZ+tF7TCwMvNlRJ06PMZM758q3VFNyg7PGB/MytpKjK2N
aKZJ2H+J+qV1sSZ8fOorZX7sUZzRgByJ0olr2BD7o/XFW2TENxIG+4rS6EsTsz6F
CJy/Rdy0uQk/PgCyM701oPag10x4vPdkQ98XPRUbF6subqssg1qKFrbx+uZNtbdN
mAvGKKiY1/cR3tF/CS0snPuAv2jNPexHyQS+3gbIFESk7Qz/DZusRcYrtFA9Bby5
tLLCG+8axW1xfGzMledfRtn7euSr/5SHn0Ykko8aFy5YAUlGflrYUKDtJPNXUE0m
K1dkSBm1U5YM9oENmkClrQIiuJabdloW2MCeipPKbP3aVzYPubjYxTXiziOuPBue
R5G4HTKuHSHZjSP5aDe34K/A1v6Hc4aZKRvPGkGpmdk+H+2BTS96Xkccy4Ue2fqL
T7UgKP52keSM0MDMS+E22RLHvadxto41XbahRbHPM8MxsbZceOaAyUjYHOaiR+Jd
oA85FKUI1U1JLds11ipyZxPbniwApY4c1/13UUcdhCFFmHGlLNZdn13YE+z0h1Xy
SOoOzniJhAm5cw6UdRGAtgzh6PcMq2juI83YZdyGmALjdkRwRcnlYnmAX/Em2XwD
C1l8bYMdFx3iZh4IE5PEBs03xkL5Ma+ygsDuWbm4Lx7Bs40qE2RCHosPS+RVXAHf
J2yCLf8+Tvfq2zJz2zMgkpAVBZFi+bH4WUYBbstuWUTqqlA5fzGP30NIVEom9Ekg
zWcAXHc+BmkkSY50erP/oqV+F3YzEsbIu310MDUg2iZLUf/7794hkagj3WvzQmkh
uGiVeGfFmXvILZJMM6vj/yD9LVomhKnbfWtgIQ2dJgGMMSy2SwzTAQrwhn1szPpH
ihjXWPB5DHAPZRy7jj23ppTFiFnMMnobwK2L9Lh/ji/UI13eacxgsp6LDl6MVdXO
fGl5ibWcV0BS1/re5W/zOUt8VBx1t3e/0TQ8AqYpwsFkO20S4sy9yY68VX2/9CYm
jgOb784Cun4FZh7/C78m0sTTQ+k2CYFpkGYzdKO7AE8/MB7NcTO+EQoXrsR7Ekpz
GdZMQEMv+hlsA6uoWYhXnjjMH257BZsUXZc/wfL1ujJiionLe/ofdg2rmapxGflR
2qdMIcKdj7i5tl/Yp1sIC262+MCGyaXO0k14gzO0UtVsSyUKxA5CLTAX8VHrWz3S
CKJfz+MuKV1H66oFzp4wwd4V/SX5pPooxNjhjR2iH1IHIqc8mTTgCWw0guBUuXG8
2LDqX8FHiyPWjHwQLDftD+PQ3DGQl4aOR7VZY66B2UnL0VMbLCxW0koHlkSKSyhE
6J33Wm9RqcXVCp+KJ6AE1l0XyjZEo147o2miGbeG70gSONPNy6p/JFBCgoW8nqFD
AaCMiuzDz1mGCxsvh1qaIqdu5FP7UgKoWKKbCRr5Pr+MUl85UNHvop5KUpzWpYZx
ENtjDKXQegUFKg9jr5lS2wA3MVKeCENMZzhJcD9AfxCks32FGIxSmuxyg00JgNZg
3ceoJGhxsZtYNSNFTxNMxKB0LYSMCjKM0UeGdz9SBbn2ODVdnOXu0NiLuJFclgbK
gdvGgd/sfqw/+ZA9hMaS72SQMhYoQzkBKevTIyD16Ebi5kPagOJE2c/a+GAJPS7L
YE2OvzVKGIeKY1hJmBGZH+XOmbWczGpU08Fsv48AG6DTH9myJDt3GAoT6WjdqFAq
I9+THAfOJc+QTsN53E+p0jQta6tHnkyZ4fJVqXqesQtDCzeuZ1LiZm0Vp94pRa9m
Yc+J5WZGrpOKCSWHy3xJXI3Pkjq+DtoXCfmuvde4kKR4uPdT5C8Q2mDRuziHCCBg
2WaE4lqKm9heENkTL7PjB/YRbc+CEwk2/p0bCP10UYbTVi6hhuS/BVo6nbCS457Y
RhpxPLGr6b9nIQqouSFKA77fAK/OTTBYcj0IyFuxz+i/fnLu/i4xWl8XbFgn3v+L
VtJWgwnWUUTh/yVqI4hYUwm0W6Cvg4MzVFzKPywNpomCwUGwzpLVaxiIT8yJ4JKW
oiFP0yzyhoF2UbtNza1KFZKLLouNIjqvG01u+E67wLbMIo9IUAh+1BioDCh89GFH
oV3tDFwHO6+8QIdkJdfKTUDSiBHrNbHSwStizjnU4PzU2ZXDfrHhVOe8c1zm3DMc
tVzLyNnMVk2bvs3jfyqJq871xF8tov9qO6eJ300emn+wdVpfK+J0Srhh9D49XQif
Sfu72ZP0cMAF+lC6YQts6jmxfzrwpdroaGndw5nIrOd0AFO5WNLGWHsQRtesDZP4
Clol61e5naHNtxH8mbwzXipk1hh4OQjikKK005Wqet6C1Zk5bf28Z6/pGzrbZJas
QfFUWc1iWKWW1sI2OS1/OMZpWWk8cE88YbXHdetaDTYPPc6/jPnB09R1WvxKag2V
eF6RCSlWhNsXZOGVn5qh7lWKwAq9GAa5d1yxAH4e0DBguZTA8fffGNWUSQ6w610a
h5JpOdh3Pvt6RnTcW3afIwIzfFOVYwewR6x+4pjSeAgWa2Lt5AC+wfyd1p1NL+To
NppgrRIX+e1r0kwya6a3al0z3BDmW/qjoLhBxtZOukF8Hl6GVB16RhKSgheUwz2V
Oa+xv3G+qErQvyX/BEKCXYUOlNFzeUBBlNQWLQqAkzvL0GMcgUeMdcBteAyoAbc5
0tf6w9Htme57oITaI+/uJGq5qIfu2gQSRyyk/cAodvxZN/K424BYOVkpHXo7/Y6p
J1pkXoqEdOjLHgD52Uaj3suiMqzOB5AWVKxTLOWBmaMHxX0be5bpvX48At2EJTGW
QrlEpz4VUKRt+cYVULanvbfbSiunRe0ETC9auDm8gs2oYem5u4XXWlWbs86/S4ch
BFEqqYA5OIG0pHY5lurBQOVZqht0PH7OKPt9dMd1lYSc0KmRghGqxUdZY2O8rPh9
EWthSCLZR1dicLUwTR81zOfbdlZksPOsXtYZpCwJOmc3XY3YjUjt5vRlAqBLjYYg
rJtZuR9TRGtJX0sYEL4EofGmvyYOu8cNDhSDhjoE2GE3FIWCy5rVlsuZaW24FalN
O3RX7UOsv5KMyjLWmZUpcgoeCwRNeA0FY054dM1lyUrXd+vyyF7/hxnY7U9LitP6
fPCpPY8ftAoWP91rdYw36/bB1bW3vvnxi89bCLeWtvb9gLJ6aPX2Ao5lSjRS5Y1O
768Sw/NP0O1303Rvm2Fhz/mBTyzRuF4wqzj1y5IrjxyKzcUUCmpVXcezXlonZm0O
A9+3S/bEcTzxzmzFwh9RkAbkakmKr53cC1Ty4co9WMc4LIjqmEe0iC8G1QIG4BZy
T35ponY8Hvf7kAxS8UsTJ+l0VBustlPpUCMzdoBF0yhwBaeIWrbRAFZzw/sHktyr
ldWfiwmng70awpgjFJJBLtiO1Az10apRpbXwAPM0PKaOXD4zu1Vbqh1B1k0ldTJD
V1he3BzV46yWD9O7iSGoINYjrk5zaKAyxk9xkLJAxygMSPqGsWqX6w/jNBQBPA34
7WVATBt4gL2IBCfo5/s26+O8er6fR+ApGay3ek70o7jxjDf2EOhqnF74hfkRNIm5
kjNe3GfC5bRzm5kd27sfFKWQs71VOcMgP1U9/xFKffrto0TrVMHjz9I68PQWYqZB
ddQKg+bxXEKS60lPCIPkYtRaU6qCWxp6lSRoKN1Y9w0XMBr7BIjuNgir+H9j0snC
+/lhm0kroU19h8FdQ5GvhvB1Fil2aKGmoRGrHmc/C1eJGio437loIkcdHnNQR/c6
gDabT7yB2r91gCBeyHK1N7/LGFmejiGGfCNfWvNTw/eEnJOx7kIn9caK0cepeRAR
gAnon6uV4OAFYRPNKjBNe7Ij0ikVyukFK+WV7lDOfJaEPAcZc3FUZM9h83fzZfe1
5qUAcArnQ9YFL846W9NV6aZvVpk3q9CXdsCSo7nI+qEz8k+iFEBNj3RAnR04bdxh
pa7cEeKoRPC+GuVtOODbbDdLswLZoJowaG2hPWWwDLXCQc2nwMF5BcKp2wDT+UjA
2bsydl6BJPgb2B2IbcU7YpzTHj4NO9SWc/0rYx0UBz3q+rpq3n3FgYpp5QZf7Niu
lzHLAEL7k/YMe7fUnUHbYSujUF5kqZD80RHa22TejE4yB1568szQUWKvoyg8t8HU
9bQIBHIO8eD4dQPnF0eHBhX3FTv10R1/Z7z1PKAPWRX73JqyEhX59CC0mjr2gyTs
EEoEX63mO20KuzreEPOVdW82yINRA7KRzGl+jaTCh/URpbXq/yTItGEfdKcC40v4
f3UIfXZRvYBXoTO/fOWuLGUImIu6mW9HOlLMOhaMO6bL8XLhVMOZZ+v7ox2TnvHu
FkAhWQYGEjyQYi3zn6rHcNvwFxsOhtWuN8RXU+7ePx3+DgkK6ZYBtpdhWCA63cDI
bVtll+TbR2nQWgt9VOtch0h8F5ZDyacMBFtmYvEMvTyR5lH9JAp/xRw2hD4c9p1z
HFAd4E6FIs6xkHMFuo9auswaLhHHhpFnsJltdyTHmScIFn2nfM6y3iTRQcea00Zn
JbjTgFMuQcp2UsMpZEWZetSta2lQRsge74eY+ym+oT0Fw4sNQ9dGKdpu0Xem289/
uOD3GEP04t8J/V7GN7/lic5YMQABggp6BO3wpBaVUqngPtOD011coWP+/zqu/Wd0
HwTNk7mF+vhAPFzpmZw9QbFZdMGuISIdfOSShTt/BCfL+sXRlRtqBSZA3FYb42/j
uyZiRpTJZ5oI7KwPcvevSMODT1jrur2p7vmZrEcGdjJW/1KB1xCW7Yl+ZsfKiNMG
FFyeOEb+gIyHmt2bUhx33/kikSHghWp4no1c9i1dONj9VOF7gp5Zf7i2gvCwZ0DU
QscU2CvQaQLQHC3PTP8VRcCK8r/qN52TPGFeEg/HBthi+kBHFwMdm7jv+8tqXVx/
1ZAS48D2uoTJfkMMI4SdL6sW+YzuVVrF5+aYdUr3P4ktlkMu3Smo+dHj9Q58TkTb
Msnna0HJqfagqkKPAtt21idee5i8y/1HlNmyE8jT+LaHPy6i9zOI374LCtsNLmvS
5zb+agt8Npy8ybllq4BCof1wyJVEQZ2HS6oTSNreVaNPdLOgkb9gyXXCl/DcVgef
biOvN8OHkVGSBk6duE7ggHEcfbB6Mz45W7+yLaf0MHK8mqZRY0cf9/p9eINMehhO
jHGKCb34A1OR1TcSyTGd5R0NOm9wiNCAaN2iZSIsBXOi+Qk21jFVACoyNpB5T34W
P1lAErZCe72N6tM35bLsdapKjhTGNMXFWmsn/KyAaKLvNeFQNwz/Mezoa+6yt2F+
vBmoLwd4EZ4mZQbGxTeCuXg0fGt6PtBD+MPEsD+uZ0ZeGH+1rq/3LexfYWwYf4Ez
K6eXCL6X+7oF6VBt+gQWXN1PWzmQauJXT9T12KR5TIBSZj8K2W8jwePPvmxp+Iea
SlwtNDo2Alw6Gfn9pC/i+DLbaEV0dqwhS0RVO9+fZAUvmdhMwuX/t2IMKQVg/IVB
LFeuQ1S/9J3hocVTVCvxM14GGWyrWHsHH/Uci0pa4LXGqlfsv0WRkurmATYtEMIV
Yl4LTwpmw2dTIgtyxB04vFlaq8ZNyiFTPDZOA/3xtpQuIc5GHmXqvu1+St9lQuwi
pwjJfTtCcYUsaFgRF+XuIxr/8xrZ2HOEp3xFPyu7Fo0PjkcO9/P7LNkK3G0CymNw
OBRN0raK0Dz5JX7IZjEfRsEPoYfWURUT77AZxVGZX5l3FBSMw1BI7W4Y6SaADJeL
pkMwBReJKmu+wvTbGbr7e91VobjAm+F820eEfxVXKNBljXX74OSW829nVjWvoLIY
s0eSY0Nl8FrF3U4vw6mzco/JpCWxDKXioDfPQlG8tR6miSB1e5GzUJgxcLPhK0WA
IneYQ5eUDXPkgtfwC1GEyzcGuMuu8scIa+mBuYVHGe8v4XN7x/XHCB6F18P/gIp6
dveUaCZZqE3Y5F1FiMd2OHYLw1QM83ZI7vrt1fBg3Oo72gtj6uBcRb7SbghOm5bL
4AYJUS8FY2XeoqfE5Bod+T+1DoCtCKuCLQEI1fQWjYMbE2s4IcylYHz+PR5p5oU+
aqXSruPKrfsIkxSKYJdngvAH4mPH+CGT8z/Cv31kCtLJ6dDL5D86txLCXimfMTsf
jHP9B7zbfqHtUhq8AYa59QPVLWxdvuPqBFPKAL3O3ZRjr5qT8xF8uRfOWJvD3D7Q
7+PnNZVv0XjtnZyFmCLIuaPQmu+6SDblwSUxWvMPgsLvwX2g0KguZKNddWCKR4Co
vAjAebuT5zSqPWyE1Vs/158WA14xTJbN67lQkkqpocKdOTSB/ePWHos4pxuFTD3Z
LkbR9IELVrl+2yv9/ZveRl85jTeKFUu2o3I8P9S3TD8yYF1e+9Bw4vBRHiFTgmuo
cxwUVmF+BYCu6z04GtreiAc6gDfqLDGdQf8OTwskEWsWmCea383pHh0KogCVPlHP
7TOMmZKkR58cQmOV30GmD2wwopPPiSvywNJJLEDPwfC8rQ8PlMclwVGpR+iE1jwZ
2rorwBD+VCyyV2EYXEPItIAyFAlgiuLsR/HRZys1XaOcHn+boza58VpVB9ilQz0m
Jzi2fMaPkDJ76gsgmnk2zXh10kVsCeyDW05w1sv2G1cyuQ3xfEm78+y1QnxxKFI+
EEnlNrTXWlNMSfvscGgiY2aVlP1PZzraXc5dohwLn2IYaDL8/inE5EAlUDZ0yy9A
EtykPnY1Ie5k3tLPGplc93BPRAuqkRE0GmFhlRFOCSQCxFMFN2OcRDAIS8j3IGGr
bByPQo/1lPvV9K4orbWz0usWTxw7N0cyqHJdjJ8I6SVRNrM5X+72BNHOkpEAI/Tk
ZxjMeouAYvhPB1NZYJEJ6M9Oe6KmNlzOMW8gcPJ0Hj0wFeqlYCXNhroISUbGtmsb
rp8iM3A7uR0R8fub72k6B/WzmHWuLOuE4x2zWLFuSsDKMvwYRF52hsTD4gXd4tUn
iTQOjiEqT1EJOe/kkjC4Xpf6C9WRFUOS7x9P3iOljsrw2XNFKBv/ptJC+97w7sUR
gMsWWB9w7smDGWV3zvs4dkLVPzuNB8/14agOyZVwd+T7cAAs0H2Hjh2TwM8jfhQd
u0/T71N0Wk1rYydMrcVLX4El4doQumWhtiAnwcjELUIZbtvl0//IHbotH4o9aFrU
DGjYXOSvjzwWn+0dIBk0wOB2+qYxFqEzYaeNVpuX5OvqhPzJ29e4iRYYxFMVphQ7
flxtmgS5T4IpD5IKgHSm7H85ax/0CBVCPdjOf+romMRFAuF1jMQdyLfBSlfYx+yQ
c3BggL44rJpzOs12VAhSPH0Q6WrZSgAcCRdss6nyI6CjgGaO5xFHzXpRs/Mxzf2o
hx+aiZd77nAwJiJ6HyKMMBN11JlCv9UEiI/3n4l6lYk14xTjneJPkrHom63v3Hsc
cijnkMjWYkAzYVUPC1uSyGkE58jF9FZHsMDy3qW6wdsdWfhVIjIAxb7SbGE2Ex0y
vu3gFImZakNhfNTHSSbp4mkqE6O6Yla2SvP7sN2EFpzn9OYSBfRkwrXLBrqAyXOA
udhRMkVJJrQJs56OVtCW7BrEAvoDeRCICmyIox6lpmlCn6h5J1mFS7x7vPozKyKn
77TchN9RAGpiay1+ZQJgwtLLEsZ3z8Ijf3Az6HCvR4PelktDWZbhA6HBk5y+nhLn
Ua+ZkUqT/nvztFKGd30knSYn2gLnVLHfp/qozweokg+gorT61R20tJX8F8g3mK5u
LLgapQRszWgj7LLEZHF2eME1TPGHjs9VjeLQn3ZQpWRW8vlWDjT/wGE2+1T2Dbnx
5FpUcaq9Qj+ebbEXgAIlISA+4Ew2ZJmB0S3GbQvFYt15JmbQAQZkmjUgUnRIohPW
wjjcQ97qKAJ66DQ+Eq6JyLuCKaYhUPZonX01qDNkLyn1lbyFHD03IrmNv8GwezRB
JNl5zzhZdEd5fUF4D9M3PzrygvqI+EtOL91Mz/hZr8aL/Qe3d4aXt84bK0AAwacq
Od6cluuirJoMuLP2Tz/3dh0JJSvBls3Zuc39aFjTMnCD3yzhAcCN+8Y5lQ7NA7cs
qL/wrK0/WgCQE3VxHFjuekbuqoKxJqJmIR4w9COl1g9mDsU8eEINRjQv7zyKjFLk
08qUbN8RRjVReuF1MrHGYgoUJgsOuZ7vNO2hFM5UOTkvvN/tq6jxX36zjHdOI+Ih
qpnlNtZGtwed6Ht+6YDBKHBhE9KxvfCLxSPTkM0FNFkEQGKLemVqipeNzhJLQjwP
Gqo4ZgQYtfRuxd/PpVsEnvIlSqpyr62Vph1W1XslMmdtvQfmPauf5wdtmimF4aHA
9NqNuE3L7XPiAl83M1++6FUiG0jgOoOcI5LfvhPDa0X89T9dxT1vlVzCVNlh2M3a
YP7CgmO6mzd0TT1pHj57WS53F+rMSlyN2dlBgnB46ZbzzYoWjYAWCYzQj+zFKz8g
h4H+JunS6ZcINqQ7Hpxb/MGpsi0Pro5G+UiHS7RVMrsE/CfryKvCwz4IFQY/e67F
wtl8YysEnP04YDQMdcfNQ1bJhRjrT8mwyAdOQDS4HdXYTJZmuu70zEhP82juDd+c
UqnW7Mry4FwEK5nCRrAI/UcDw2g9L1hSQZ8Bvfkeyz3mg+wdVETyxU/DpJUxPabX
Oebf7zIcAFIgdDZWYCc8WmuFsb/fY7ftfMlciD0z5bslZVYJvi9OUyZFwsCWO95G
XRVfbrUPDvizUvHX0rAXXgQfPtXKw+CpsU2iCgGiMn/LAskMMNJCWOKUxT5hJLh7
M1okWeoPnht2iaB6YUTXfdB4CbRJjA70iSPvI88J9V5EtVNKUabNmXKxOynhM7vG
w1ItInffaApTaNQX4LfdY3LxHOayNRQ7PjlM4eJyZGueB4BngV4vzLuiJTfGnLuW
GrWauxBgaCNJRdiiP6rv7vrwZQJcGfWGbIMYmqSwGn1fVwdkcu7x/GdWk296eLpd
AmE+4eovLmDooMgrFRtcJOtSUqYxVtFEZ8KPwQbw1LScMUKQuwD2A9uhbGdQnNN1
TPYQzPlDOBGtXM02cGPKqWs8KTHWmTW7vl+4xwp3d3GaWKBBxT8GLMaNEASbp9Mw
QPJwpyVHJb3soVHumW8K6D5TyhmNRL+2FF50zG1V4MJ6HGpKfq0438J58cpC6zFl
F02IuPD50rpVZc9Zh04TffNleKCcgbVc71WGFurJJy7leV2UtxFYhHRIQMqJC+Kv
prfdB3/+TQ0MapOqWByhL2pIwOXs6XX4B2A8xBv0mITusesVxtfEbsG9xo4Iko9q
p/SOqkQWcOU/RkkdjQGUJqsgLvK6ZaOI+AkY5yzrjPJe9u8MGpTA7aDko/I4ctq3
qeXac58C+sfY4MA+N6dx991EStLqy1qGToNnkv8yRCnwkmfYbYPjZX0rEy+nyEq+
990NWb8FaAzXiyjFJZ9r2a2Uuhns92iQVDPc+uFdKLoU3RKx/OjXg3lu2jf/66KX
HiIytp7zTu0yDXct233AIO+OPmIo3qwpOn9Wf2HZpXcVLGJ3zMe/zezLAbhkd9D4
9QvWF/sxCfBw3SY3LT7Et993O19bZOnXycKQrdOQjO33sioLdHEg12vuWQ0oGBTB
ORXm+dELuZyq+ACXjdUjTiLDRAtZ7UdSkAzXAPdrJvUpVAE3/Oiko6DO9UOi4SiT
KViYlgaerWZMjhd3HmgsSbRxxbSUVrCu2jktej8/DDTnEOa7ICqWUWRfgwsHOpQw
soOiVq2NeD0HC31EEiAsq4ByvRSt6EpuMmfseegqxCF8Q3dBK4BpoO7DrTbt9Wub
7UBlHExAaw7BoC+svxpmTa6MqhmNz6wlu9WEyphc91PGNJwPA0ehtY0XA0lGPf1v
SiYMulUpYiv/JK6fFOrHr8kahqLe3/34YeF00jTPNPa7pPkopELu0CFPiKzLwPnW
/Chu+V711TZbA61C56AzMW/fQpG5rHblxyDvb2roBbE0dgdMIumx3jxRbNECDnsV
ckJJ6N7D1KVCgDR9p36xY80yqtjXPQKc9olLvrSGofKpukaG08AM+eYKdeXZF6bM
KX63umAi5iLxjOEPQVmUFo0c7yRKRpYKwqcj+51+VLWeVSNHY5TVqBRwh5EG/RET
lgCjb5zUs/zpnuKUkRyXab4e5GPGrUsi1JZP+ImK5HEIEyqYjGxHubDivMWvoXBX
luJBqka8uxMTEao3meWemoj+vReDoeHFh73vvh+Gf6U83npY66UOr3M0GOs82aki
wBYakH8obCzoLY9uj5ty/TVmWlPxVlqBzxxRYUVhsVRvmeepA3GRDLa7xRe2mOJj
POT9TwB63/GA1yQTfPZl59eH8R0BWWCYAkpATXIQwTNo3XpkU6HzzrQ+A+ex9d5R
PUVgmGYAyeOmQEMkt1A0SK+Nz751PuisC++itzgT5eCjdg6rxqn0ANzl82PSSb4F
1DSkHTfRDDTeUtW4HevUvLdHc8/VjAINfdPAaZmsCt1nBXhCoPfb3X5KzYDXOilL
iwRe11I32Ni1S98Wby5BhM/bFfXDEGV02NdG6z41R0fRFpsfgPPwF/Wx9Y5/K6mT
HO01vfBmxWGW0HcvQD/Tu0mSbyN4Y+yl3eIulXcLZgBWOZlKjrSmXIuPab4GbnL8
nl4YVYSOzgGmTfUUQyjvZ1Xho7ekJ3JYaBgFHY9UjT1xtXClC81KhDqod3UMfsFx
M+pAEDUNHitb4/2yGo0hGKAHXHys2C7hqrx+Ct6HLfTAJhGHcmV5+JVo084ubT9j
roGuDWX9wZ/ahpD87OKtxPc8exA0vDpOW/rR1PXWYkOdCcl7c7KazIG/mlgCPQdV
OMjIsGp4Ieqf6boRIOAmcAnzD7aOoksHHNmlEzzkzDv7Gms0heB39bl/u71DRXSS
SmzjC/vxnxRZxNN0OWhiCfEvBeCYJVd8rRrL4KK8GjPktk8AXs5cnuKO1ih6rT5X
+jbmfY4iEp2cTephvKwtCD+eKeRyTxuMy3qmZ7FXHctnw2er40UHbavePeSmP7uq
TOpNifuIcGpRQdNabJUFG4JJg6I+lvE0ItzGAWAQUopl5wO2KNjqVvsjP7WFL+T9
Mtk+HVVTLxrBkFOlLPxpUgJLROOUnJFKzSU0N3RNGkJmzGD/N4nhDdC821fssOIK
V0GsHrjanGQf7QaSTLrFMCf5E6Cvl20ale93FxRi26SNMyGL2U56LArGny9BG/PM
5mG3R/xjG6CY1v//QzqqNbM31Sv92zYHLcCGMqjlyTVPtboGYLNoarQrR6JIetVP
VyJTtYRW6FSRefGlMI++CeVi3uw+6+ihPZxyA12A9mKolP1p7u4SLCG8MMKt6Et1
XNq48poj/FTHkFc3wUSk/QfmsThDD5bt5CqjHIOo4wTPOxYLD57rS2OZI3oy6/zb
oyk6kqGhzVT3QiA8cDPvpNmcceT+OZu8ZkTUIZ4oyh6Ik27hy3MhVGkrxg+PMO8u
cG8F3Drcd9YKoyxYd5+dy///4Ii2BkNK3Vw/Hw834J57P6kRGSPpa6S5U+mq6N6h
EjolbIAvPDQoRQmBkq54kjBtLMLABhDV4U2L68zdkr84TccysClIrwXyTM8dQz5S
EpEgHlDxoGzpMbKj+ZfOEMghza/Qj+mY4Nk1X0DAUMmyZBHBQIZPR9WhrGRH5X1C
gwQBLg/NBSe6KsYJth2ZM7ZURjZE/zDScBJ11iCwBEptoXc2q7KL0ewz3zd1FWR/
qOyx2sQuep50VacwMa6MIKnA3HTR82hSfs8mC7QuNl+pP8u9IuDk0tZ1uJMCysRS
VwCpSpxTi5O6NDqJJUP00WqGKGfbB1XMv3/WzlTDRZ9aairAl9+UAy41UeI7bfup
PrKrDXmHBk0nFrJGK+6LUX2TweC7q88jw4SXUnZRd302gbNEyzGEqPtPemZK+YrF
zuCHtV+mzIK8Mgx46LDV6L3YHIsozvq8AzRUVKIhUhDQhDG+mF1ybwc80kuR249b
vXnOV4Qh9UVOE10aNmfr71D8gokNYfWzB6rfq1Yz3rrhOMtOKgJj5DfU5soaP6i6
Qc+tKABKA4piAuYckmIfyC169CVE1rTWVtOnP1l57Z63U0de6gB4P7qIpsGdc7Go
aErHZ06H4reHS+yLPC8RLPJfQZQbAN7BIcgXdrAvnQCTNRVVW2kldz7IFFo/4ciH
6UHBR4AOPmVIRq7nLeoCLF85lBuePmhYSpDc0Qqegv+h+0KBA6NJWsiXnT/cca95
OM4cH0wQg/PhwCwlIpReRJOh4be5kelP7M3s1/Hapbz0M++Xb5++zp6vOV3lvc0O
jSYmW0j4f9vPNZL6L+ZRe7MOatXxLs7rhXQCrLNtsoa+GUPD+e8uu9AI43HOGhKi
Lu1TTUgemRkhwpTRCClMDipDzplkI8wOJJ/gjw0bOqnlURJpM/z1egz/L6qhwGVn
FTU57xRxHSEjC4g/JODkHEr9ziEFTmu9G0o0Y9AC5rnFi0M6YF/6SQR7KXR98Gek
6RCRPjMZ35zOLhIqRDTNeLY0AEkZgfu1leopbInzLXFFy/vvGTNrXw6Wopa2bRjH
m/Mv2mL/bvtg6p1USVn8NXEtmJGqe/8INvRFVKiCoPntVb/iYqAdrW8sWTPsAVa4
T/fHXbGPMV3yKzHC48rErZf43HsRbYbPy42QNAteQ2wXKDT4Y02aJqw7pRin2wnd
FbVGb+EBffhOtRHNIt+uQMo3yGJ9XGv5DRH1Ub0/pjvLTVJcUEY88XuNUVhqIh/W
c0BZC1L2wa9OAKgCz5hJeX8c6o9JPAxgg3MmkKnIKvNdRUwMPFs3VTV/i3qDmJlA
cmsvpvXStBkocBYxRqIm2rs0f/Eo3O7wQnRYgrRY/F7SGFQbu7eGIr3q8rGi2Noe
yMMM19LF1q2Z7E6VxTv2+h4cofvuEFIxpoWu3I2dAMF4kNQyYNj5Bc6JlZAPy9XS
iGjLfO5RgdrTcC/5N5I5v3+wtzLzIltGZ6T+yMlbxq8NLwsGub1M2M2x3+W6OKj0
8w3XmFz86cXMOhdXxmJ9IMi41rhmZEKhFkEaxIRgu8C6NSkpVU6YJcS/UmEzimnc
ZHOs20LX/XTPdrYO4j/yICzdGPoalO+OccprTLkDERd3ohOS6xn/FVkdAMejBnl/
TTtqRKAHZeEVS/t5Q3WUFgWJVbf6S8wqCKT+F1XDcnIEInDx0A8QYugxT/LToGJL
VRvw7J6tyJOLDruytouhQWE9YLPCbBUflN3XjN/RCKo+mWAoOvYnCNMUdiRNs8c5
hf5f0K/QoQPmf4JWS9FGLxFjSwUHAs02ywJVINps4qSvLTJQK0j04NU6R9XW+gno
6G2aU4HrYmSIZA1IdFZzoQb50b1wAgybaDQ6/hFHxYp4Y+3iH957TJZrv2qn6oV7
5+KQWnZ2Jiaob09q3MGpOcxt2ppIBB6PDHuKjdYxwK4DdHTSrFGsYNfuhJaMIHKs
SkzWAvpw4Q1fTQKkvyXgZHFrXO2Z0g5sQj2HuSjpfehWQnyD257RHGVyXO0rvY1J
jlHIpDVOlYYFtZt0ceISo8BpukYp3YXcb0rcqOWPspjM8VMNJVrm22N23fYk1gop
9oES+zwVwGgu8AallNI0J7DIgd5ie3A95SgIbT8xFeF/3hlib7NfSIe0PzxwFal4
yyCTCXrJXRG4XpPyttPaU+uTXVmO9+rhf7p26Ub/R5xPJpHuDf+UJ0tNOv+DfEcS
92nTh3L7Af8XMzSvZEqyMUcr2w3eJrJwnb+eh/FMyajbmptuQhyfrdQB+AUeVcB5
1/7BTq2woUEZgtOzPEKG1JSXOa5UkqE27stqm12fSLMvsxPvCraUoXUlY5wqcT5O
OxKxhEJZ876mGV61AQ6wQp7ivli68aFoq9Cjb0riQZSHscLYxQCJF6Pems+nWMhm
+jCDIakOjrKjwt99zzxsCyoivCx78JdW8GM0Qc5/5qS0XcbJuQiIgnLDoiIx1gPy
l2S9x3RrBF5gIBfZ19upx2668NL4rQadv2n62kyFbK2Z70E9doifSlf8H1Bzelun
5MKIqCUCbTSOCgPnexXy1H9Fd0ytStFTzhSWykM6mBN2dxyCO8JLYBhcqYRjN7ak
2xWKaJNCGQ4L0AVgQQ88vTfkygu6Z6KlRbx6Y8bjsI8BnOgkoCBYiqHf4itKYxzL
EvrlmaTsXwAb5wYWQFdl7Ah0KnC9oP2xqAYw2+EBoqGOMm23DBYGLbJuBpQQQ+EW
71GJoZoCcLZT76HHyC4xWOc2rQw/rpXOa3IpEDkkdlyT6gbEaLPgtjxZWb+cPWOk
gJnsrFKqMKAlGSzQ/cwZ+W/t7pXBrHtmKBn7C5TQzMzbk03u12WmFLrKr+bpRv5T
FeTGUh5haGHuBtV1yco1qtda29DVPt2Idh6VXib4TL0TLs8BEQjXpQjUd9xsHN13
MSWDW3Agw7WW0lF6v2pwmhvon0YtXahEy7tYSEtCxFEEQKqWF7Wjc5G/QCaE2NiB
fyPegQkSt16Bm8o2VigSlI404pcny7Ob5AjT5d6Tt81sRLujUE0dcta+ViT2FYZG
FWDSpGdqPp19alua16sp+0Bc2Cw+h+ECjxVGvxIKT046vB2uuBo3bDweea/hx+D4
ErWqPR75smz5+GeiuEyqw45q5XrHcuFfYIEX1X8wvcQwyHV5yqvtZhRCV7C99ZOh
w/VaMyi7l4gLE+ITsf61QpQ5JsEfKIsYA1hzG0k94mTzwBDG9qXMBQ0kq8+xFDPQ
vY6VZZAS/8J8ONFoKfVBfCPwjID6t9rGhJe4dir125u6o/MeLM73rv/BzxgaZVCm
mBpp5lx28EuTxopI8wAWBvnFSAMhA5h/0IBAp2/nsAV6BJTwybL7e2OMlzHzFWso
JqolmPILpbv+xvr2SjVFE+FCha0QyvcLYtJ5R/oItxUXyq8DuBVBZBZq9VPtrIfo
QikbIHlMpQMkSzslrcEHLzzPNjSN4YrvH70IOEmWJ1SP5U4iCuNex33+/H12sgcz
6tnOXHlgY/ZOD9EpuWcierfkwQWyP3ReDX+kIsOTNhjFXDoVJ0Rji1hjOo5oE5y5
M+HOFMz5Dt8iu1vmPdMSJs/LcoMM/vrMkD3WNHFnZpSksX2Q8C97d/tnd9nz4Osu
FW+kVw9pm/EjkU6k3SGi8S1hJNf+9T7XMzUam9TUyrCbuYPumgBCBbA0U846vnf5
sI4WK90B3dHD0LynjbV0Q8DpgqAJtASmftrxILq8m6VmPfUqp9H+KQTNJ/wWcJ5I
8GfgDDQSGpeNN2pDXY1awGUIJVKl8AKPkM+HcjClkPWh5BSKU99Ad6EjDlvqN6FL
cqVwY6e9HPbkFqMz31EOUlWhaD1V7/02NbFYrrgcAmeJO1Xzaovt5OoL+0Ev+EX6
tdQT7Q8I2cZK62ZBaMkUCumB1Fyx7n8Mp2XAwsq4Fidj3DR5vGjj+i4YBWsrIoae
vezg3RbOWbPMBbn6szunksEf6f+F+wHnJM5FrDF6ZHc7owrCCHlYcnRS3rvHxbUY
lsbZidYybjOve13AekJwS/rsvW58mi977ajmu8lyNjUUfiX1Sw30Hbq9Ir0TDHqG
SY6+fnOATljdj6pmX6FRx6tMIbS4GAghe2zTK+qgZxYZFWOfXyoiL1ODIWkEQTG5
Zk6W2+Bs1H40XIt1yonbjWCrztt6GN8IrpZ+mynSaysXt01IFZH1uzhXIefCIMjs
ngXwqIJ7xYPeCsC1HotLZlniufzVhPTNAvgSFvkPeyGmRZer+TC2BXnSyHKURieU
eeujsL5ueBdFGUliD9dpqlTIGfj2eVLoR0ifyMCW2dQlk4GnkrlOF+ZRU6OT9q7b
9/EqcVKHE5e97KdwSCSEjGQxJRDHn99b04WTJsJqGAojtRxBPsHBysXBC1QSTN8K
DhD03+6nL/x1yti6Yt6aWrGMd4J5hIeBPG3j9oFqGC32DoTr4tbMVnyudjMu77og
Nx+TqakamYMTc8l/F+zPLw0p8Zkv6fzynlIX6daTD2I8eDZJtLnF/TuHv4pmT3uz
iL+ryRb0yHAErC4/1jaHfqJFlb6RMGeJX2sN3B2f/Y4M/lO66K/lmm1ygT5rNhsc
Snbv0FP73bff2//suP4gG6Hx6cEqTXXVVAqPZOIQ4AXrqPs/KyoE1cspKYYMpwGR
NcVHfP9YVE3imPXABOpFvD5VHXVM9r841iKzyGngDggyooumpN/p2CdpDPG2hA4s
OhEsjSPUXGHItZ/FtEiSRUG8bJhLxo6EHG0KK+7GKDFRjjdcUjLsl6HMBegR5Gno
2ow0Rzhfpy9rMmKXBTWylVYBDNEpHM8k9kfNOL9RREsttmEx1fVuf/XV0DfBZSqJ
0G92UyVVn7GaFFDP4eb0uMrqS33HEtZvch7KZFz3iN4yUXpAYmHFnfvgvnMwCgrh
9oQaxoeK7SfKFjNXiNI70UDJUlidXlarmFqgzFrZ5LecV36Q438OSXqfT2omwM6L
VTmGfQmEnpu7zoo4L3CVcTXzXe23o94jRE8AxHJUUfMtUKUS/vaA9UN3o8YFqQIC
coXWC94WfEEbfN6qJcXaeQ+dCHTONp9hdoVTBLU2OA5hBzitfgwF7zsD+iPmYaV3
aRGbcRRGmJL8DrGkMaU2eYlIebTrqxmsLM8kh92rzfXWyjXKHAkEIvt4j5Y3jat1
bK0KbZTBHzyFfB76b+tmTHZXTj1aw6q4k/6+Zdd+9Z/2s+5Srfv8IYkmzNXSXw+q
o2wI9f8fSjnu+2v+IFKHWsAYCY79f2cXQV9Fuu25wq+yvoVlvw+DwCTPpd2BeGHh
nHpWKNhgRyhyg8HAijQcCuSwNPRnn86vO0Lmpyxf5ITWNIhJ7Kt8poLo1hPTdYFb
VlukyhT1EvJMpWrbmIpB86QD+zFqsFLApZhSifDI1WXaEnexcTA0N/iWSxqxWwiP
IpIwtbF9UmWpWVE/qEIzJ5K7aAwl/I1YdKNO1aMXAD7L6fc+ZzYitcOqxyC1l4eh
I5sbZTW1bpnKMT0ifmuTPDGHBrrNWq7qieAq099IDx2I1JrEoH8p+axl+Pa6DoFW
D35Rfn0nuLQ3pwm8V+tVM7cCaxahsuca09OH5IL9jD/9mzzCWdFbTvOOljzPRZTH
skkzpESv3fkGbIxqAsKFi4jqFsyX3key2LHk6H+OPOB0Oe7Yd1UXlJ4ibnWpQV54
TP0tgxKLf/B7SSowVaC86QakjGKhlWUN05f7nUtrDC+hTMevAqF4VCz/eU/QPhre
IM6V47+k+LxTjx17esobcV8Jefozay9qfs5FZ8g0IHW4FDFiO2kYi4Y/8glTkorA
xR4hSmGWyFoCoxbQ5uADc0Uyb/t9KZ/1MxUXA+I/OkSUbf+6A2FAImEv45yFaM4K
JLOoKYh4qvuCrsBeSpjHKd9sxpKZku6bBT2bCHHM7/y76CiTPE7q/6qgWlneODrI
Y7wGeiJelVWSYyBVBDZUCzOK2Qp6N95DoLq7ldX19frmDCdDpQkHdJL/5Qg2b7vZ
8su+yU6DHbT6+Dxl8d1urv4Gk9gFSTeSWR5IIGO1G/sr1ycXkBCyhU7JTZ1zevDT
CcIMUDaFkDhqu0TwQLymZjNzJmBM1C4IaIDQJx2yD6pHY+q0sYNEQ4pzdqxU8Poz
SwtVn4D3sCgeIcLudb4DaUN9fR/ouTxVdSy4LuRRjUzuKrGaF1jiZlGOWbPzQLJc
Q6SGnqz9riUsllX0jGUuaFy+vNBmbNG9kYkm0vZwYr+ja7eJ0wEx4lvOL9rgjBPk
OY+wXh51CTetXDq/He0RlUaeESHqwFj/IGbv+rWFSkG7/YnQyEycJ1/JQIow89PP
sDACHSaxJ4PPYQrQY4eKN+gUUTKjbIldHe3uj1tElN9oA6RFiIv/gr2CXrAz9bae
DjQHMeBOPMdIG4EE+Fujqzyf05WqL2/lyvePL7JU0yAawCHqY5aALdUniq8Q7rvU
HD0bcI7kMW9svdF78HZqq30dpTk/XwSggyiAMu/vkNxQchP15PAGtHqa54394fTg
nOC7j8CauZV5LDUCkEzt8FmJywGxMiMnzOgFbNSLxmh6q66zZvembaRH5c2E9H8Y
QhCt2iGtOQ4GKxBhdSCPSRDuFhy835IpKNXEMJkgBBGymoqtWdmE+q+QY9GfGbe9
UqHHx67uk/VFPGK2T/ogN+6JDSqnE8VvMZbpg+WqrYUPhc6BVfmC/06uSmjMdBJN
hX9YaLQBhHQeM+mWxCtp/0HVRHPQ+7x8XmuYvxxv30YS0928h+U8pWSVmQBKaYy6
nLwzc9O9bhFNUtcyHsT/XYw8OtVF2JYEz51K9Nwz82uxHC4eoEzQCXZQ6720GHWV
ExDy8H51Nyp5E0edZ0BSoPWxxaeDkOS1h7x4BYP4Cn7MVbAIm83VFu6xLBSr4Lz6
WAEGwAVSf3P/R5OSsbagZek9GOXtmU44R2Pj4oSNsc+CyyhzyK64/lwmL5/tld+d
PUWl1OGH4MQ6K1rz8nHyd0f+jmkFnVnMW8WTz9Tn8Bin/v5ZRVQ9FCHaAAtYBLL3
n9QFZ91l4pGd7eLmnAPWRSwimyPty3HLGBYYWWs9eOM37dYtTO7W88P+mbSwLnqM
YcnEKiqWoyFM3u4D6U/O8dQqoFJV1przdyMOBQRLY/HBUxVkQz1lpYG/CrxXKHj1
TlaQd1MtH+PQxxKo+NMsN1B07H4/IwIcwaebL83yZ862YyuBG6eXRjInO5v8pnec
kG9DMxnrVtMSWt44UukZZsUCvxOi/ia75OFFpHG5BmCeXSZspDJ6/DDGdCvieRDk
rGeWl3QGsg+EKwKsv0Jeon/vbdzZxkCP1cNjI6uAd21RDbP6187kidCoV8NagcQ3
Xg2LwoK7uteAd3EOeVYGpqIWZc21tqo0Euk+W9VLw0/ViCqfl3l8ef6nSFfo/E4W
IDbbmmS8wHsdGkZ/6NRTLhox1xa7xWSx0NDzjXle257uraA+fsMgsVORCr6+bLru
hVFjZk38iB/dGTWf1wjW8N9VkUVxOTNPHU8QnpC1CShnTTc1gNvTpq6KjNuhaJYQ
ji/71kRFCMoQ/+Dbp46y2Y4skFLxWKxUQWQejzJYP9mLC5waSuFhMCFln7Xa+nZc
u/067OKA6kzCGbbkZuqopE/TbfT8Xz4Zr2lj1OIyXyowEV/BaQkzXlbKHRrQU1FU
QjuLA5LQo55OI34WhuRJ2qP3Q/ApWwwvwbMPxB6iOs0OxTcKjheJpBnK4xufHZYn
8DmUJqb6TgFPxbMHqlDtusudRLHEyv7U2gaxtwiV8XL2SJRwlWh9Ibngov36JLGd
wwM9/SymAgdlJMlQbQIevpc86LzcgDpD11BLwPOVc0cyKIWbvsYvWD2MDf10zgQ3
+YKAuQdO1KlAWf0+7z5lL4c6WSGaOYmD+GAq06E+kaBDfRDofWD9ZMyueNNyaE3h
jqzNGcZitfsOUDAg527HakCq2b2ayfHW+E7xXA+N4Qr29Gb23ryRdevNwFw4+Ldf
ipNR9i2/gRg96IiOFYpVG4VSFMowKiNWHoUx5uPiWqkT/pmaz4hdv3VcJs2V6qvI
PEpaiCGyTCXj06dGhDDaefissKJ7XMnt3HqmdnmUl1/ajH6QFJyilXBXECl6t5x8
5/8dpnFSNArQS6GoBw2sKimO8Sgxeq77eqYAA6qVBbIi889RKwbzytY+qtfLuweC
Kcojq2pgrjKh+Exb8xRCA6myapB3VnHj9CB+M+1JyJlFk7WG2CwBWXZCqtUw9XUS
bfghHsi6007PHqU6zOFq/Lq75pDpXZK81LhP8beEu2KJHyGoLkzU3K6je1TjcsWM
oZSKnlgNbkIAFVC/YcWwWC8Kcs61B/BaehybcF7Ga3B8QLMK4/5kmiSIYimaitps
j71OiBJENZYkEcPzXCgsrLfRVR0rDaM9W4AU96J0OoRixSQanvkDr7sTHdMmSdEd
POaXoZiw4aILAKvDV89OeRxeArsErwX02j5upB+Jmv2JqBMMcB+2TUAZ1KYHBnxB
74PtvAao4u5B9NfT0KO6dPcKoc/iYnKvbe1MIeZzEiiLSEd1oUPt93wXAI53HVGP
jD1M9qHJ+N7Sumj0EAiZk940Rp3GhdtIGjt82pzoUI4ACwyXsXnU5DgIYbjqyP3/
60STmS78rm0uZD3CpZgFYJ3rS/Ngi6Us3OmDAmd7ikPgQLtDInkXWyIpnjuREpM6
kFFfVbFEYh5u2wcTzumiSiriaYGyj84oewdz5uzvkF7T0Fwr/3XtCOgjI/cbIDOY
6LJmo+NONP3IFfvN/T+hXX/y5sp85p217Dci/eAsK2lMndZJT4bAEd0XqyqZ4Rdk
ca9A89eqj7FkuxrPu95mjJtwhDBqxgekwUF9bnW3K4uCJz7pOYJrihbiwuzNkwdz
nEEaaIkG7HQyql/TJ79HLkH7spF6bldK3vZVMWbaF0YXS0qgFXqnFPnhB7OnbDWs
Cak6CVmmo9WhPMVsY8Jzyw2vjdaj+ycQ9u/D0QHZsdAKw81BYQPlGFcBZgrIW+m7
DGchLKjDkdi5Qg+ZOy+MIsLfBfvizN3jSHm9HD1SLsCoPVFDFzB2ik73pl43ii8R
xg3fK+trAcZCrRSfRQQETVTAkJ5HqJ6l7QYnT9ByG0bdhAl8Rk8sZYvzBMmv+O8w
CkkSw52OEjHafIPN7L2PIgXrkQdc3yIive/DCIhRkbRUI+rxc1APICgRzJXb7bKe
NiPgVZ5/UA2sXZAR8qc4z76ELiRmEUlI0ym33u3M7bVno3D64d1WsczWXX5I0n4Q
SrWizGIlapm011fmCUe7FpdnjT0EjB8iD8dCFQ4Ppa98aDtF5AztkbIinrA/BHst
pw9HbnbXgUwk9Jkv3hHUOKfGHIGFcjzxnDMILR8VMTf9g8lZBA8v1QLhSgWKWKeh
lPIuWvgpLA/oFFOw7HAATxKSp8CKL5FgsYZE+AKlywtv7PNYZidrsVNGKO8y2SvC
7RLVEjjTP3WfvVgczkUlvXmSCkna9oHkGPTWlgcyT+A3M+NTDH6iN8zJ52bAZ4iT
0V53BD2SjATwiCiQWypQyAbcjsIk6+lsUEgwKZbYMYndz7AXxRqqT+Zfbz+5wQLD
HS0pv0UQ3OnJUjEm+mLaXHSTHQRTbm1S/WYUFDFQkV5IKO1pzx/n6sx/ADehtY1g
vFhRsvRmygYH/I1d8eFbsOtXkNkaXL8y7P2aw0ggHy0ZSXXaVzZFKmCEMARRzLDe
16j0u5UQW/eT2yqNByEUXOLLqFbEN/QhVS05smyBc7suq4HlKf3YnryAtwtQD0Dn
Q+8Az3u/pBiNXbkl35DK7sQvp921/5Q5ZEZ79pbk8nFEMyDSX+h/HzDmdS55y5AT
RCtB6nsSzO1vBivoGnT1rDh4qePyeewhIOORNXzWgS/PliXe3C8Guoyv2VkPqxlp
bFsgaHv752XuiIuJ5g0b47mDfXws1YhIPYjRNTx4EBc4tagdSq2UqvG/DuZfbzJd
uF/ZSuC+A8MMk2p/uL1DdSL+c3lVQ5BBv0iKuIimRqQU38TBP+C84f2se0WEntbF
m/XVsHbropAiyYnc12qsPTXTWxI/U5LZlrutHkTtYutqp139pEXHhahTPqtar/qv
ebNpuPJYbNGbvBS/M5NHtt8gQ+cyeEfZ0R4V4B3Ht1KyaKOlqZanaaUq7jBcb/QK
LZgvBK0svcUtjYjrcir8qaTPcu7xBjNptNVM5dNHzpQ2oM1KeO6eCNj4xnW/sDE9
BmxyUGhHEUS4Da4HpiPWTn3dqKTMyU4Mh759sNQp9DqkC1VRpromEdxpk/9olapR
M7P+p1X7EJkTxpZly3s396qeaFaWCJsCvl8CrQJ5e0SiC+H6HyhPhq9ce9WkMQ3d
eVJzT0mWerI5GUckpe0PGP2bhVmgJF7RJ8vX3DB2fAGi2AAsGa5b0h0HBs4SEWto
jYuJrzLHSLZBGm//yBRSZt2m2EOceloBZzP9otbTnR9sh8EkuINQFiR/Rr0jNkWx
mi25QJdUHbbD0cU5I2Iv6v4A/CjlZb0i+A9EiZAsYxXO8V3K3MZy4rjpv8aXnhry
LjMatE+DRKa1VwkpZFve13l6WBLfnCmjwD+YxQ0fz9ZdAnj5ACpH43uvbK9xTJUY
fuKzeVL+Y3r2VTzpwfnqE/yIfC3wM0gGJzE6Y6FDWTRws1E/2Q5+tm3TZ15g75Mj
01LixjxPHrP7/di+4Q9SkiDrbRWVynfQudp6qfedDdBgl6Uu+wOVCNFMaDh7KffZ
4dqjg4xZ+x+99mmLDnUoQvmrJpj0Sz2iZrMPoUoP31Iyh55v6vXONVRJD3sYGtQW
jCrEu/TYsAqiFmRxxwW/jAxOm7q62ZGSi7jZcY41ELD90QpkYm0MKy+7gg7Lvpwb
hseuMcDzVEbTNLp/68Ru5kE7gxBR10fG/5SlSOEOSZgCGs2969lfIIJPtaFyJAR4
ivZ8GG+UScygnwxVcfi4cNyeKYTGmsx/F6zi5yw0Yg0oyzNhzIvCo0zlfhlmhswG
ij8iW4jbw3AuVLoOUO+i3vaQM7OFRwWO34150JVLxK+AgQy5sn1/g140uauwuR+O
VpRez0uzy3ErhTggcuXm32Sq0/vgBUP6lULfQFBE+N0y1KSrowkjlhCZsnQAUKU9
Qmguq3GCFogegBCHPqa824eDD//609no4XF8tAgOmpVxDL7DzZaHbqL6GrkD0Ywm
OwOJ2tNiI1YN977CU7/enII9u6v+XESuBSeCEM5/0awLQr036dLJ5Z0MSSNFi1F9
dqs/JsL1a+cbyltJmbCKxz96nyi9hWArJvqvFBj+5XfwoU35ibqEU2x7jQYIW0mo
x4P8ggyrHbXZy6ZLZwhyc3PPsBPgx+Vyn1Fr3HfkbSH9t6BdEFVrB3coW3I+ZUzu
L2N5M8HWsevoca77rpflfvz7zlAfWCuLAPJkQhaRfTV9mMDL248WS7MwsBJGSGPp
eI0U7WAlVyTThL6Zr14geWbubOOaxQ+st6S8a4sL5RVIo0J9BHWPkmvM6Kz64TeD
WmSLL4z6nWb9N8jwR4GDdpVNqaK4a49X1HuEh2pqz3n2SSzKVZkbZ/XgfuWg6K1u
/AudzT0ZtAeRkBKsPLgfNdFiZID3KeCMiubfBrt79Zgn2fiXHwyb0dADWSNosQh9
ZgCejGBqYU/4V4MoV8Qr3kxRnl+3XFwdf+XmxyCjeNqfBKsOosykM2U/+ehIIpO7
3o1iASe6OthbHhU7V7De/Nc+/UTHBcgBV4rAPG7Oorm/OcFiFdSq5VoLdASI3OGm
s4/NMRvD/M9kmEoESd1qmLrRqVVUMIxNs3cYkZDU8Rpf+VXfOoZ1QY/e8u3VuGEn
m+c54bvGze6mZdjQWQnxfI+Ki3Lstu0HEeII+zHI5pX/SkLXmNPWIH3BzP/vnETE
9akngG9E6nfsDwBQce7zjWNp6f/d7Q6z7On1gPGjAICh4a/LFcXLZP06M5oSY2u9
ZoNnhrSWe82juUvQ1n2lrO8VlvBlyK31HXZ72gjjNYrFtsS8cUq8MOSNOu4euohZ
QjrtWnUqw+66fE4OiPgZB0dm7JysS7DA4hOKt14FDjEEUYesV0qbigGJlm3r0L00
AW7z1UIPBa4W3b4/cxyvomRg8cKWPM9gGFL7r5/XOHvMcP109j1KXztXA//lkXCQ
N8HmF06g7L+XAwIeJ5smUzYcrPT6NSOzEfwUH+MuSrceiABV7i3rmeZ1AC7nPEQr
oqaV5m0BkBtnnEz2huD7nhJmeNVVDbxDMf7WHzU4xDUuw/DCVsin3yEDXnPDK+VC
4F6RE9x4H4nNVTnI8SKvqT3z4sEssMzQ4SK9w6/6xgGx0Htq8TVbfnckmz8Y6fcF
zV5+hjYoDCwoxj29PZxtZ4uiXQAO6SrY6kA7hHOfGBFduesXFLPFXwQx2fAocioR
NyC9+Z+QY5zYK3XtwMP3L8O0b6DknfbpI1c+sL2pu16eVwPkoI8rgwGTovGAFJzU
wWJEJBtaYrX3GOGyAvyjeEbUHq2/bPad0wRSOR4eqXXT5k+MX//3rWv3A85jTbcp
G+JsE+IAkqOJbZmtzjPMwfGty5k8byS6pA4eq+VrJY2qvGeay29TF8pXo/mUJYAv
bHguhDOWZD5jOlUmNQDkaee1rTRMVfKa6gOElQJ2zFS57Cod/CGZt/VLJsWdMHtz
7W8iTcdjnirqOObOKGlUSFIrgZraN8IJ2TV+G2moUucgxSnorAnMU2qF0qces+M7
rG2wxbNHPv9DhCHcpfbaes3tOXptRheR7FVFkGS07QRnPEuFUfuMqhmqI+aE08GP
w4FjppdY3XEDlJ8mp1xTcihrltv3JH8E46PTpqykvB7D7ED2zCQ3hJYWRuoii6CV
9g9zt1rHEMajb1tGXZaOlDm2Syt9p+x5xGQlOTsGYCZKmk5TuaXEDFMNdRL83WrG
26cCilIdkx1H03K4g2UQ51JtxYhVSddTK6dqKtexCr4Qth2RTaYkiO8UnhCUxjRQ
S/A1EhX3QXpF1CCBjRhLJuw8DUZnvozD2IIQArOSogM6JKF24Os/tOBtOWs3TiYQ
LST6/XBqUrsH8oy1B95ZGama5arOVYU8XdJfRetXo7SwJwmLEKIdlppUIhmDwGg4
zH33ItFNpf/9OrOei9vzk1AArrKZEfuVepk4Oi2Bv44W8WxQXaRSaIuJ+W4KIInh
NKpI5oAfyTtPwbEszlPpE7abPSUGM7k9DixvL04wfRlS7eBbTun6XVSRzzlk79PH
9Rniz8xqSrVYRrOH7kC6pbxzGJtetxBwdopIukk9AVQ3BFWQv4HzwPpQ4WwDJ1AD
BUfimxi6f6+gZggUbc9fPtAK9/lISK5l4xg9Hkdx4pY9bJ8Ag9Dr4/j6nUZLl0tW
z69ynmgoDF4Py4EeKRwQo/TzGlR6X9udQFCEr1mY92NAf+S7PSjQ32Ysa7OuyJaK
Cq7WRfGVpxJ1dnq/fD30Gnizkru2+fOmUhgLM6KQOEVoqu+J/47A7A41JQTFhNuJ
YAGyqNoKKkf/QM5KkwQWEKJ5/2fKI3fzJ3f0X7NCL74hMOHPlgob8YTT1A9DxIpg
VPovQAbx+vfPzCn9J+VCiFnVvHAH9klyEhKdpuuzh3CYq3pYhhtuBCOSaQ5Owz63
md4hAUw12WsNBQgdfNyEGNKCE22WFYv60F1ttanRpIc7SgVuB90Yg1mEt+NwIUM9
bcwlr1+YX6w25sHWsz5gQPivL+SFhGGeckeXeQPXYmiztVZPLyoJzeuha4g2ipv6
VK/QJ430dpsOVjNiXKyW9T4ehD2hRL95DXU65YBSdz+nDGEbm5YRR0tzVv5x4e89
1H1WTzzoG/aIUFxz885ZAGlK20yoD9t0zQQZIBsDZm/RNUZL3xLyxTN/78Z4S3hP
idwsa5tTrSpn61IcP/zJtDLtrSkxEAjDVcMzak4bia5mHoaD3KlmRVoS9v4sgAHJ
zopZLGYXiodd6IpK85+53N1h6eFZ6WYZyM0Knt7cq0p1hsqe5f9TNjK/WoiKpW9a
lBCGX08q1KJ1baLZ3lsQPfgoq5JK3IYOko4lGszMqiwlhOZTnyACxof2rBVqbIwZ
t1ZfR+QwGV2VIpNQsQZdV0+PNVax6ZKrhTb0e8nhyoKRcUehPeE0Y6iQu+pnMX41
eEn/OD3gOwNaE853fva7P2vZTldkJdzeXlOVluaEFrit4igEZ2dgcZPx9cbJ+Fvd
5+DwW5T0TdwDkJDCooWdycu4U+yZ2+XclkdiQpZiVJYgvetP+R1XhHgcT4ztHJqo
Vs5T6/tRMX9puRf/w8r72y9fem4epNKDR2P5mNPAXEuik0Hyf0J6OaZUqlbLloSP
c8DSJ5YKH2xQlpLmA8Sh4MACTaUc42/mkJNkxtseMFlpLaLkJCVf6FkZWf7MvAxG
/pcy3doG6htvmFxHrpGLXFbut/iT7aF4p4Dm97JPxC2q9YXGHb+Rd5JBN2N5qsFV
ERWScCjBmB0hQsCLpaq56ncX6i8pNkuFUoRwE8nmvEx1en1ooQKOtm2EJryEoAc+
xu17YZ9h0sL8VvyKcohONRGyxnLv1lL92TtkrgIoFmRkoRdSdEj6TMI1U8kc6wi2
fSO5qCliG522yUMI3lPEVNhWx5uS2My59ipC1QJzxN01FOMMsCD3XE+pCxWfQ+7B
H8NYXBHcHADcq2i1xZbAiar+CFQnuWPrLdatTWnvk2iqKOt2RoEHkVMqEfWuURZN
P4q/ZbkC5fPnLz3RttSmgH/zVSUr3A4p4007C17R4FmPooow1aePlhuuW5CFzRJG
ALICYFF+eHuK93APTrQas0oCXpZtA8qLDnA95YYK2xLSwu2aUq4puQw31mgn7nhI
GsC4BIph/k2e/Wvjr/q6IxVnv/JG7T7xVItNLJlPJsXs6bQMMPzjIoUUTE8vvqOf
T8TCUYwXIdxL13lkR2OhaYkUgRETpqK1mZRMz3iFDioAdNn6seYG3v4qyl4oXhlW
Ggk4bxSB5c03oJvy8tqe2aSbkBVS4hdHJ1A70Op537BkqJ1UBXM+cNtyfUtyDGz9
tIo4esdCV5zo0yuJJfJ29URzupnOm1yCQBr5Tz1O38Q2k/hPHJH5ow1fMAxuHtY6
oYTCnw2hkRsQVm0yhrklwcAxl+e0JATr80DaG64cfjHtuSIzHOV+vFwDWlc4/dmS
Kqfy5Ww/a1eCXWMt+7Cw6kDCWKY3MFV78b+YwM7n5xmQOTJLzyzTPPkUin/oryLt
me5aaOWfpLKh+jdiGd8/0dx7P1d2ctIF7KnFGY7bkBqSe3fC6lho76x11gwS6kYR
gpvVPQ0dAGqw+fWJhfEGpmJSiU+GpbnR6kUR880r76z+jmIZ89v5jjkmhW75EXeI
FMVgLaLvCidZy7IFfnmQTMWBhAd4kUg/7I+taZyjnCpz0/P0mj8fNc2PWJbSGlfH
rkrFuHe/wspZVayXhuRg1jum/LDy6ym7gBnV5XW4Q192YgKEv1QJ+giBjW+qO4sB
J1w5LtmlwVzDb0Y7hYA7RxBfRis4VoI+HtZB5gFjL2QW6ocWoTCHYmgnx0KlUEpg
vybvuygFRU3Ycg5EuAyRLqwtQJmLOxP1ssHcUe+YlyjjVrXx+WHW+vTic2HZCkWa
QCRIzMej27hr/NbCl10aXsbT7c20ty73UxbnUgXBhGjG+fi08+fDLtLr4GNVn7mJ
vjR84vE3EM40dWWVD+D48wUO1jyyRK62v5QjL4NNrGBx4YajVQOg9QczTdmajn71
daNtzk0T5sOCiQmZEpgjZZRhg87nYWLHuQ8Id3QADty3WfuRcmZmp/h3xV71SP7d
HjDwC2PXGhs/X2Ay2nG/V2v4w3W5njBXEpnE6+C4SWwhAV/zQxD66dobgKJZlx4O
6AEVtbxDwQLl20Uvqn5KQw22/mzvlIS3XMdY7fIXQqMzTfBTiPqyZjrPuJenaX3i
HALJFpbxIaNGBLYF+xZRN6V+FJh2SPjnM8PR4qPMDBvEmQuPbI50UegZiBmQYYMp
3JEu66w9LstbuFFzifH2XuUFrziysdpVek7l4SPqDb8ePSU0/qoom4z7FJrFG+XN
FDJCPeHPjq4iiriGKJl0oxAMyCWSO9jsUtv7Vfyz0D4xmd4QuvLJnaZwm17ahROT
hROpSCeyc38h92iwg2Af9YUsPx99tbZl9hyOEMoELuAsKD/JzCNptI9RpRd4leqw
3fSVL2TmCWAS8DIELJgMEC1Pf0QAySGssfFufIG/bAyL3QB/wDi6x2wScyQxSHFw
zVbh+41yfi3xLtTaSNrBrIaCAAW2ut8/lJdpwU4TaIGbScnzrhEEFfuellItDM2x
H0DurwC8KIfPmFsFu28OqvUYaeCSm/K9Gw+7wDTO0JD7fhVnjp0pj/+YbBwpopG6
cXW1SVSvEdV7TGDsh2xB4Aw+Vx030lG/qgThuDS0y8J+IwQSHwi6qO/EAvvIe64F
CcdxBf3wyP58L+Wc6tzk2ExyBAZeZNxRjhu4MVsJ6CzsiOd5Ilc5O4G23YN0lq9e
Si1r5xLZakUkTWOITW6OKXVsGrswzHHySNNTksS2R5c0mXWUY5B7CBdrSSXehlz7
dKaq6Ozv/CnE9LilVk3WWGkFe07eGkzcQbkjVJzCp+W2PvE2/iNI13Ws8Z2gR+/e
NL4kIiFqFqxISviTcc2qExs4GbTHu8ZEE3pJRJxweqgb2I4f21O9vy9m+GcO+9mT
wIaL1i8Jv7J8T6/gnjUpzZ0Yk7+l/X4DGrqyNLKc2wSjQVd8TF2NkRAyjsB4njX3
LXGfFrvw/cXeHPTPabpoL9xNhe8FeQbrMh1XQ9EtKrnaRG33oYCm0OjH810fgVAM
Pq2uGcwO78ESh4++y7uE9HF3DSUxtV4laz0XjvbkELHaunN1wBD+JJygVrKpoOZY
1zu/ZGUfWU/VFvewlfJQ0CyFW4x9HBZ/jhgC66r3UX7FrapDxcnjFWYCEwiYCyPo
9rFAAA1fVUaIYI+s8bN93fbi6EEcqE0Zz+4gObvdkHTxULmLerLeiIL/T2Wu/nh0
8wslYXTxOAt8e8aLuB1Pd1QLTWZIku9RXsiayL3OCF9P5yu4GRBYI3G7olh5ZMye
FmtQMMBcz+V1z9cWCApPjKo3feLgUG04ovn1N0X6tpP7DNs5+BvpunEN564cp457
Ur3MVX4l8FdQm3e9ejTZN6nonNKnEuHGIGG6Vy3YNHx3MNkxOmggRIkWyCcC0x9f
Ti96pnA6fpahzU4YPWrerAM4MlvgCBqFSwcv/9qJMQHprvmAzdr/ggnJUqXDXhkJ
5NrWAPYYpkhgCfrXU7ki1iVbJJWREN6zr41mZteanFiVyc37MapriYJpQRWzFIJV
8l13bqOxexQXhPA5nZ7WWi/cYRs4OUK6vrpjzgvxQbPjuMdi57GZYuRJLwPBUkJE
dBvmLagJkkNNjXtdB7DCv9rRwMRBgsniB/FbcKDEARmaG/1P6+5MCcMH0YbpJiFW
7I703ZhUUKODbGV9GPAGcWEy26ykWoYIubyG81Ak3UU5gkqljsN1qou70cluD95G
frR3SfVBmf324nOC+E+Spgwj6MlBY8xEfTtBqlGVuNvyzkrGhRuvXl7UTnh4JvOw
+QRYxzH4Im3b+lgng1nY7wg1osrTz057v2LsW0Li/6SZI+0SpDRJBlfkmCdSni9Z
5X/Djcesd6tklh5P0gM95YRtqPC39rhV2mEQ84+Wdye0sja777+OTjAwlrj03JTV
0ltQnRAdovcRvYwDyZLaLtjlx6tML34qtmqxpD8O/mDriW6DBctGzYrQ9/HyJnHH
axcJQ3gDcqBjq61gbIyhIU0mGM0TqBj2ssSXu6hfH7pRNQEOEfJmVHUkYrJ5Eq9l
Z/QvnHHQQ7G9lVZQD2AzaWnPTpy/ElXEXLJr7LqS13ucvx+kIzXPothh1dSoGkol
nFxybcROd5A+s/yynFVbKzAgK/8QbHqlLoXm64vMbVt43KwLdyDF79Hht2cQmFBk
rvdbPmvnivt8f5Y3pFCxhU4IeMoYeyPyi4r94GkQcmLVD7nW/I1FOA3aeKwAI6W6
/qns89KGPsXsis09+65vJT1rcBrZR1BExFcT6gCH4R0Pmc69dS9gwZz8cW32G0hY
7Yr1/P9qN1pNpJkXlOxiKL8klhY136m14iiX0z/oKtZL/rh5Cx3IjDSZEq3VfJr3
EosW1qBRYag4RtE3+Dl0hon4duT44vq4hkfkX6EfUx/IARCIRJKtxamiagrvNqVE
IpMn5/fr5o0ctrLkwpx3ijBeX/uNFMWCeChs6uZy406hLNbtmro4SWEZ9LwPMGDn
PlVKzZzfgyMunyR0ux9hy/4WLCUaG08/MwVG3xRWsr0SpVbC87aEBOsJ9RIdT5Ev
qHw7Es7nTZxBfVF5ufN2tmUtfHD9NjnheXaKPsucTBC1bweqvi0ZwO0jLjJecDIo
a8WwcfVMYppoeLK4rvcdzajSu9YdE9s0stcY+LBWXqI4eEl5a+fVm/sQoIvGH9gq
nbm/Z3DhpC/0rNrZ+GrRVAvw+KQrVYugt1G/7/tB2is+ro/3v+/nKL2adM0iGSAs
raI99kiesU4S3E9S3rG3NJ4QROOIa7lk8SQ4wvyoLvxbYtVX9+b6Al5UhjaMmUwd
AdCu5rVL42KvbGR+ZO6sCA1Pm0oNxt/8OD6EqOViklvTJlxaQeE1FPY1lTmxEmuP
AvUBsBqV4TG8CV7jVq17tZ8exJfXf9AeY8jO+c4l0yia4tUkJVyqnZULLJzydAqf
1McodrDKDfveVHqFtJ01dclzkqnSrXWHG8Jqwvoxex+oKi9GC2j/uxQZ6E9WqkfJ
8SXaR+nOL5FYD5KzBegvEHuBtxFXlxZWYwxLGxGmcQF+ojp04iGZEP03+rwJ2QkN
nBZUhC1OSCt/uVtoKtgCNSSvJ9E1Wl0ZYW6VHonLTWBd3+8wyMXx1UaQOX5URZXV
+FBILkLudOPtuoni80U48O0TJYDSUwzrDkDdcQdjdeBGa68QoKz2VUcxQYooLl0m
LeB8EqhZaibE3d8iAZjbd6+hZ705eQ2DI3urMnx3PsLJ/wnJZMoHSVPHdB3GMjro
wOdwRTumclLB/+AF5XI/OOZUt7PBCUHIVD08WAI/FcqJCYcpIusDp4ifi1YLvGx4
rHLdnwr2miBG1nKJhpg6xPxpSN+9KC1uitky+qKsfDB8IRHuqGDcUcRdL5KLYIP8
+4+DfKxN67E4cghPvaCVNKXpUCgql7LSm5haSC5S17a296cUFvI9bYsIHdQDe17A
QlKurC0tYhbIqjhHY0EH796o0/eNR1Rug9IdA/ZbCwKfhbDm0zA8SOowxkP23z9u
8hx7AFyD7OCuima64CftNwOs3STK8ilvNet5DfH5bW7PMcFtyn+G8JvhSOF5Axj3
aas6XyONZx87ZCtvH9rPCOMKHvSZ93gy4w0fyz1ycbWGPWt+DizT9T5e/+l36iT7
6VwH5NQfbli6NVpvy+753BiRqdV81bewxOojPaBMTgdR0Z5eo+NzI/1YdBitFVrt
phb1FpZwVAiEDHTC7JkgxNeXTVzJNzAX33i7lLtCz6zY2WeBmJuECi3eJQikROop
ESavbEmNOwU+mUCJwIYVu5KkG5bpPVNJH89hV1Wm61stg/2Btj3N7Oj1wmZ/9sXo
AImhMVeppu5gR0oL6zt8o9Gh3znqzuuw42ERrEhFJtijNzJK18fEhZ26hwSWm6ua
gZcXjiXHeSrhiqFJ8outgmYm0R3Kwsf1ooAiCbaxJe6V0Jj+JYp0gxStaqwN6PFt
c1MGTQ0QGJakr9YZ4xdgm6QFqOgOLn5JX7bEDemG6ySGBHr1a3j63/HfzDwHU55d
RAlu5Es9MdVRqnu3W2GwoNPuwuE/ZixKUms9U60t8Uk8/kdnYtiDr2qyosNAX5Mv
PHrQ/c/+ZD1nqPrDSomn/b3ThBhyDYlkKd+B6gA2csqvz95FWFm+0OR8FgWhgfLI
3yESgfOAgq742bV8d4tsCpLLf6RUV3j0yXlOW6qmrFmTFkPOra+lpy5QlkNBtys7
3xWxEmHkVYqr59mfgaE1lxq7kQuxwlTfWm6bDnLWmZKRIEVQEl/7A9teQGo3YIUA
b1I4Fg+MLs8cLXhCzEHP1ylLXNW+dE5sjjxsB5yXqvyOcuE0DQGtEEtz+q0MN4nS
lz0+edqqIgSm0Gt5LAZ5QDO760XqP9vZn+rZoCxCEqZtWTNdn6hYSEsuo0LzsOQZ
6Chqcfw00YvkGz+WQeC9Z1JXfWWL+WaYN0oYnlbdVR4zjWx8xBB0+0BULAZ9eFm0
Pg42Bgjb1NGZT2qsYfAYNo4QnjwiX/US5lXLxawVV6SEKHjFKBSXYlXUAVmdTCxS
jMs17PD339wYmjFeXDmuDEQPl05E/PK3Dblz5tE1FlZL+0P6hWQ31/DpKaCfU6pX
+nbCP+yLUz7MseD3jHRJ+oPpHIzeTkiDzgpmnLjvjL1XfsE4ZsOBW4WA6gv+sAhd
cYS1lvktPShqoqt+9RytfnvNRYuP7r57d164W6qZDQ3+GFhcpRLvwWLcTa2G0anL
e8R4N9pAfKdRRgTCnp2X3iCLmoLitAOV2t0VnXcKRbZAKW9eFBQRgv0eejqHvzYV
XW4O6MT5VD/5X6mQPmKR+M2YpqTKxdwxRAK5DkVxoUX8lt4DOT8HEJZKTZf0Z78w
FQmLdKJkLAtmjrDgrCAXhj+jDWsVi8gM2f0HIB2Naj5hcvgKQkVU64GIeOiRB+H3
u/3D53miPH4d0YU0Wgggy9TGoqYd7usguIiShrvv1aNUDTXzHLaVWqOFd7ydovGu
VEDRCzbF7IsPRkvLaTNP3f3jZlLfNWNiSLQbCb+kbFXWgfwCOy/Vt35BnpEhYsAi
gE5hxJAwODh3lTetsL89/3kNdX+x3fJJWwdqNpZiNo+sJtt6zdGIsOPgMeCJ3Wsg
lBhXVWVd9ZI5SKfejS3Nxbsm24XNgNA+7+nQXGYRw+IE5daNf3dDaSpRowsyapBD
xNd6FGlfh5+x7DIKJOCS78hK1eQ+izk7sNl1LnA8Dc6oRTuX0U8+x+zdVzjP5dVl
YBBhuz4AMrgiECkxJTHg85rZvk34vn/neNqfMeoi/5uyux6ev0y1m9EpAFnI8plg
THm/u9FrKA5My3xBCfeOLC+FDAis5Lj6YNUhrjTgvstUkqxpyIlQQCtYOdm+ErTY
Mbn5cBhunE7HHOpXgWs6aqaeRK21K8zPaAFJil6gBluc1XyvOaoqEa9Kq3w8Dr4h
9wy7kWyMls6tc2PtIL4SxJp8yPUadno0R46wPvXGXZNkqxQm29x+YfhVG5t7GmD7
C8tIox8bq27bek20aI65plH/eEQuNbT7lgbF9hjdOVejvZW1WK8aZok6dwvGyKpf
bUqvMdPmoRCQvQl8K6QyfKeZGpBo4NNZ5w36cAgcHopC9a6bnlaXqknQ1ycPa66U
hc60A1D7/nowWhpwBWxz87sU0Kvgt/kw922AcwYpBVipVV5uitqNfwDOlJv/78SD
EV78nIBqgcK111oC7vHg/x0smlQUH6FQbvCrFoHK7bZ594EWz85iTmh1iTvSsnjW
Dc+ap7lHMK052Y1RjlGFIpnApfGpPDw3JaXfgxnRNDWaENhzE7MjkqxDY1NpAkO6
7RKf08EAR9+CDI4rGCZYn19RJ+w78Kl764lbvdF66AQSXvEW8IYQwEzf74uWMm9q
aZtKyOTzsQ2qgzDUhYkbn0BgOsiPRrLTpCifr8egBtEsF8FcMey0Mw0iZQ+QKaFx
zyWZm+evi2f0OgT8twS5U5qpraeQamx7GpKHcDoeZlEuU5HT710uqryhJm6tJujQ
sFCHMlYw2qh7WJ2H+sgDU4i8shgBWXwZg/ib+Xv8zcL3ceIdOuD6bsXIH3MQuUCJ
JLGtV/7HtmKrrHqP3ezXRytSLI+tnJlS9xGAPr/+mLKq2TXpkLNABbPoSZWEqo2x
HxD1v5yvmWI5TZWrgKPMOg9w7BuwYSxUSKODtddpZHFxqAla/SQJJl+GubbzXCGr
zbBOyvef6pVzfuksBShAHvMzsnEZ68++qo8WUSKvyA7svleTDKf9GBFEQuMvQU5D
XQfme2K7WeUG+wokG5PtGPJy2r+L6nnn8pUe3JM1tRAdl4Nwrm1Eh0UtPQdozGB8
BcLTSS16OA72bkwHPZaCdtx0fGjYDpV/ERqZrwnLPhOVgtDQQazs4BSOEVtYzCV1
sjYVlER0IU6cmjFv1Qk8rzS/9gRtoFCcCI8+yldvWsr1BBlOjz9frPtdJeLVGUJm
6xc+U7IfMtqhE8EKjeD03Ka4mAXIpMQL7zPNUvWfug1C+I4hgmNDPN/1LLB1zT6t
QF/ta8W8GSyBvugX50h2SqR8kCGUsjY1Lz6MJIdsGHfE8FfqKCZDLU4XXD8ch5Jk
pL8ZUi2Rr6hcGF9j+6/hrnvWAOO9m6Tma7dVJWdMcGsnQBTKEG6vYab5FCpJAej5
B34I/ry7tteVzfagB9Q7pkzyrBMgK7+Yvg6KegkE/FA50OvQIeUIiliBBP2vkUHm
O3zl97vK2uc8h4YiL9TWEoh/ZeFvpuH6k3DgK9LQeftk8E4hU5eUXkFkIZPYVhfj
xktLOUsWiaJ5uzM32wzuijl66OBIGjDwSY1AnBiqZnsBNH8QJcvaz+pSOqE9Lutp
RZLcFLbNcgiKBdK0q/Mih8ws4nwidYe5pFY4Dn+evYKNuDCn7dA+tw0wCJOOxO8H
UH16W3O2/c7XpLijdycs+Oe3wJVAExkNFf9nToOktPJb2OtUj/IyB0sznbTO/qPp
3Avsp2dCewUbk1iIbu7UFnSc3Xcq+nJkm1cuc443wQb0+n0Y0cL/5tG1WRUI3yyM
sVxkvXYTfSzYcPzVDJ7Ly4FmJHudPPQsYVW5Ngoh+Eue85syG8NLOoT9L5gi8A2F
wbXRBnARuMpjZFPZfxVwBwWpwQBJ+NYv85sf4VO4PfEmpMZh5UzAkSvY9NY/gu9u
9p7vfcCf4j+rY0zLVhHpQcl6+bYPaae203p1MfnbCUhDwL/V4DnspSrmiwkEgZiN
EztJl3vvi5ox7T9PeXOB8jY/hHXN6/t4+i8TiH1EGjxTGETR57q9UQsHcHC1pCeW
taktV6IflkofOKww+dY6WntbFZ60ZnuvUpM39uC5pwBiSNRop8X9LKuMJ41WOqxc
Q3Zz54DDzT3MDC1k8ZHvin4R3HISFw1t4GHQCD50AqiVgjmPZzb+DKo0Sod1Nz1T
ULxIwgaUZ1F2GceLBvT9vVfzq0jGL3ix2vJNBE5ow0FN/kJURzQTxUr6gOARq3JX
7IKbjw8uzWkO1F8lOhjzvWhO7B1Ah2cqDdD5BfKBdOmvuHQgNbBh6wR24DoqBFRV
+C9FNYXWJOtrbDXbhWuLNi1XtdMViGk2DPyPmGzYG4UwnQI15LU/1bCkJxQzxM5r
T/4bPoLqwcRQRwFNIhRCJMP/aHpsjHjeLqHDMvosnum+IVHJ3w4TKqYTonlK7nnd
JHeOKYyHnRbdQbwwxcSVarLxqvIbkPT4BooG3IFE88oYqTwASp2N3LFAVHcpePVM
ojmEHhatk0+YAGcOAmIqHvj615CfvbJ5e5iDSlI0su+YKd7SEZSo0LqTwPENRG9n
Hwju1/xAzx/O8sMjiohf1A6hgxycs575mmSOgc83JNMdk4nOS+Kn9N0lARQQTob7
aCZsr1FSU0y8nIcxGI1RK6LyA/UhAYpQplzOc1oqOkH2bFPg1uTS6GqC7JLT8hxR
ii7pdEX+c16WADp9fvTee3lxw3dbrAmY1xc0PfianT2slyO90/godaA8EehL3WpM
qNLMgeTgikbYT5PbbkFJcIuIGjGWw0NcX97O2Z7jdeXwbAiFU3lpGSz7za2YCZ9J
KX8f+K+T7C9cVPKjIWwwp1I34B69yhneCHFg7uCW91p6v/fikyVsId0qQVqvIs9e
yCwK760NmB6Bt++VxfBospH5c3dPVzuMMJiBRdWq+0ZwEn5ZBp04AFT5pnvNLZ06
BX6Pex/3CSvYigXCGzH6YV7gc7S5IjjFAjqCNsTt954yPncvgeGkYROXSgTtEyxu
qlIwtGKuttCv7bgnGm80D//v68LHjmtA7KyGX5mc8r8AwHpj6FvvSzZure6tmUaB
iEfem5pqmlK9zHyjsT8yzgR04nrF9HJ34hpNdPZXyZ8Y6sqkcHEZULfpYscFpF20
u0S5MpwlSi3/Z4whgT1huUypgHK1SD1fjj6nuhVB/0QWo/k0qC70OqoMicd3+CmE
Q49qeapVxp5aOshGLSab0Nm5dE2TrOqlvD/jYcjBVbgYSOT+fW14KMmdeK23+9oW
7TvN1h7PF5LpUZ7UhFVXSQsM3lUGWFvIHtprTd+3io0R0SPlPaeQgM541a79InuO
6PJeSFL1NXd1gKrwDX48b3T/5UhZ7i9tCqjEaaDLhJtU7Ek25JoHdqTHtlLnBg9z
l6NIxd+8EmRZAAALS4lu1e+zrLrCExWWE0cf/fiArlOVOp0pj6mBYKR0DtCwGvQi
W/yqua2xJCffm+N8e3UTj8FLMs1SKO7kzwuBz/Gd4v+PMiEzjcHDlSDGWtw59F+Y
18NP0ZCG/wVc6R5vs3YKEqa4SFxrJQK/v6Kc0ahKaVfP7+Uktp+t3E+BrGZZEa8M
rn6ljn9T/NU40deX3aGPjCP5eS4b+0BpY7CcMkteBvgAsOEZOC2ZqNcGAh27LUsR
ejZZW6Ir50OpW6IqZ5HFEIRJUgwrjsDJAeSkqtTxGly5zLkU3UOcKeXpHPqCdxnf
ym3v8OZI6dWiwfiiBlIgu2q+w2KOvDgBmwJ0lSDf3bY6GXUtpVybFLC/GrRT/q4M
KlNkKdwKvQBFwOyipV7Yv/p1cirA6xnC5eWli3rKzfuDD8IwmLGsEWGMsfOY4qwW
LdgojpzZbZLjRYrrjjGSax8s3QKiwwwaJpM26qqOH0Ret58iKRtwCmsm5cOiNSvy
XvPjeJpl9/o01rctPteCD4d+ZzbxFk0nhU6o7I9baRbsm71O8wY9mlQi6FFehkui
q6rJxVpFg8mUmwc+RYoJml6+2sEqsX+Sr8AxtAWj0DcJCGfLSsnTpCyHWRrFG7b4
xml2WE0/iSLhO3Ik2oYLFeIIagJWbAuOmIUAnB00hvMM56WK4Gp0s1BIsczSVsYq
Wh2A+xPnRhUVCcWwKlBC0glUN+/I48NdZfVncJPq9Ka68CmPIWgBBFIda3wAMSG7
EmUkoRP7ONXkuWE7CL5pA2av2d4NoHPE2IlCSfo5Is1itJAByPr+hPQSS1+Ex0vL
0Kc2MYRjDC4ld+LAyR4ybngy0rDQkbNla/IxQoZcwJ7mCG/O74uzXQU7Aj8UMPDI
CIYlw+mjwX4U9OZl4vzqSOWthPAYS85ttzqmlVnFAgUQwgarEmdWs61XkNhs3vYB
8ysuD/lZXpQnzaLrP1R8bx3m1J00SvKlGGcJLbH5IoIR6DX6JDkPsFZ+okwSC3OV
dn2KqbYEEAUR7uBD3y3TV1QTjhXdPS3oaI6f9fW9U4QQ7rAsKce5kOJaIh8OTrcq
f/8xYEh6oFoBOaoWCIgJNPvf12UzOyvukfyU5kj7OafmCI17l6U0u+4tsggb5i2B
Q9JXtX9DPJ+cJsdX4kzgAx/s0D8LJ1/hy2yb3kFoONn8YGcTpzeVlBLA3PYrB1W6
25APmMlO4ORuM+HYmh0PN0C8r2rt5Hf5M8kZUoSC1JbcEHjx+BF9vZbS/DtgAELx
ZLdTuH0cjQjvpsud8W4wDq2dSG9Lq1BptqjDWnuv3dLUyF1myGph8T8mpny+kaJO
X9+1XYfCHXE4JuTWxU0vZDp/QhPYTIyRuOoiVj2IS/B6ujMNnAc8G6GxXLDJc/C3
hjIEzexfL723Anr07/vbdixEgY/KjvAvKireCC5+WflZNjIe8tDJT1uXPlRu8PYH
lBxMWIwTDr401H8w4phfAwRYHaE18ath0FW1DjaMNhyvb8r7fP9COE0VgMDAD0l4
dsROhhWffTkpf9XX4lDyBL0Cu+P0QhW3cMKZPMinCS2JW3AK8crE9JZ7X/FsmHiO
844A2giy6s++PGrjpMuxDk2kJRYXAHZVwPaGdxu4L+wPvwn1JU7ductNpTW9ciHH
SVqU3bx4CXfbkvWLccVg1prn4O5v4OBqDe0c0ujisCWD1ivNQmQfRFvF0rGcfWi6
0g+dlDTovufEbT9J+offm0XXLPPjgcrY98RZ9NxizWTRF4J5Jh0BAkiAzcZyzB/H
ki9hk242e8WKlGP7TSXiyVxLpjKKuZYmDR9OawaIR8qKOpg82SPsp5VUDUQJ/PIu
u0PJEJllYyZaZ9N75Q4tCTxLmJc6SXtErduYAU8H6McWZihTkWCzjDZJwo/tBwYv
mxc5pcx6Tv0mCjJ3PnYht0nZsnC+V4LwYhLB633sLUljxVZHKvf4zAaT6/4pdO44
fDq9vNJzYIJaOLq4bT4VZuSamThXmwTXJ+AmSyycFQm5rjkKy6wv4NACIqulB744
peo8Bhuurc7vfKikmvFdu5XEZeFLsBC0EgP9U9o0y991tIhMqoWZWQDZG68EyEo8
98/vX1ROC7+S/hYbFw6X356mZEVGAdxzs2Ecpt+0NTC18xn+kWlRG+gR4lSFm07v
7IFYq+uhaokbMMgx16C9I+bs1HVJFi89fK0nejekc9KKI5sH5UzDYwoN0Vh6uRe4
+G1clLMvYx35tUVhM4h0ilMgsc+QwqhMO6yzlsdF7bjApgwHT4xwSv6I6WsS/jGM
wLApjLtTpr6ZzB3ZjabPgNfWHbtFsjuMUHPHaOGF7ocOU84KRHQ0RNRPJGzX9FG7
aoXUUPnpRnKrKcX8tWFB2UyXVebajt4sFFh86X3o+R4gCj71Vm9SxJDyQQ/hZomF
a8LQemizfDhejUgwc6JyHuqBojCS8cbuyCVwYYNI4PKPauPjFAMqppTH5h9g/Hrk
Z1OacOkdbjIP6YwrXx2jmnafVOY+1yWQ2UEsp+zOz3Wqq+lxl0qps66yEhyQXIWo
AQocheqLrDh176ToxWeqfh1W2A1x9cHDNm3gEPdh/2DlVa2IuIcJE9ATrOuMgGWC
1uFD0ZW+zROEn6woNAzLTnYe8nUMLICvYKsPuK0ycT/2UBXWZvJAGiV+/028mf3y
ngslaPj2OrULthQgrj1SL0YiAIle77ctuQTy+Q8w9ucuNMToOlNLDIe4+eZt0r3L
T6PTQu5aw0eyBqPNji+pLqsMxgUr+Xkj+dNPbx6vpYmcIBG80h9HISzCOVC4WWFp
l2Ax3Qs7TVzmJrfjeMmv7Ph8T1FGdX/4Nqm6Ll7azb/YPwah+eSPUWjyJ4/q4AqK
ZQx5jVHxNHI58BBE32NKEMssGZ2UR/GB1OYgWU5sBevJVM0TvixxZ3iqr1nMNpUi
9jdkTUH0klp4YXGk0f9sc51YQP8tvNKSTjC3rB0cABSa0gFQdIwEvExuC1ORM54e
S8xKTfcw64vuE87nRi0v3+in9YZ76vzDyyE8ve0bIwDgxjmP+vyxfKuca7ZlRgKd
UF6kLCbtmdLeYqVwSSyDtV+iGL7K4IbfkD4hbHoCbFmUbiogpMoTAl2JE6SADc4h
DkbH2HWQ6vErr3L3dhNKHhVR+zfgsPo7mJaWFjqalHySJLgm7enTFEeiflp++tCt
rNAD6qLhoiaOw+v8uOc2LNGdu7AmA8hkEJxEZgoeVGp4Jrpwo9D/m/oMEfstj1Of
ozqoQwc3qNOl+hkATFEWah/G0fpX9JIaem2NeoSU/iEWku7BHmjGNugMRBkI4Z4i
BheHEv1fO3SmtR2dmVy5V/2T9ZKRrIVxb7prSEP66mIs18dD/YmHayX4R/itNesj
5SD7seyQTjqwKcraG4hlbFif4+gD8aUNQhjS3fi4uEqFoxwiDQsZ0QUwWzuDttoY
4Nk0j5tnm46o8BMQaH0+x9Jg6NBpWn+L4Ppa2XJXG4or5RHuOZxwnzzK6vMR0gLg
IehIMx/Q2UleLavl1E6HGz7cqbNDIK4KxZ9tIILcrkjZ2JwlWbm+zGznrjQvIQjL
fkZ0VD9BAx58Oui6ZB/3ILAL2OBkHfurVeGiH80m9T4YaG0zUHEaKH6loLNDJVxg
cgwjgKK39qCGq94V2ZTkTnAcmj7Ka8YvfnN6IVELX5hIz9QLKqYScAVtuSideRvo
nMaKtF8xo4dytdIFxJNcdGVp9SpqvSVUBFGymFUGo56RiaLw1NQP0N8UjynCzsm+
P2g7FuBb+Y7FfqTqxXZPvdUWDPTKd74uxIHK0MFLGPCmsGirh0wKekcgjcluvJem
OQfA4+KDbjtD66sBeLARr+HWmfIonYu1EecFyja8xW/V7Cj/XdJVzANXy1JdFgCH
HTKgvQcsPtnSs3stT+52FX+LC66/Bi8ES44G4qaw1njwseVb4MWfzoCYx+5sI8ox
aU4OIUpN6pJqPyEMNQH4Z0l/UierhEtCFmmULHPfPZienA3tUXPNxjQSjnYQOgLe
XnFBC33/h5cLKlffoW+mb1xs9z7rCC2EigKfKdbNMHdQJiQSSFvU+GsWmrgnv/wZ
BPOUxEiSXQjjshrdZvjBAjGid7AaQQEkrWhJNdG1fxQhLmvb7gZvOGbrOrFZbk+r
xqlXxZZJJuGASGx9ptSg2IO0wrH9FujRk+J1xlLxTDj9Dqz1IFlVkvEUX/ip6F1k
RGY08k7ftA/rRiNrfn31t17vxCR6LHX8WjmFOb1ySSz5DcdNOiMjI1C1ZxhNmZH7
GOt5b+cMYeUtN5aE/BpV4FoIzf1Y4o6kZwPKuFYTegj29nWe4RNBH5JlCDR+t2MW
cKa31QfUmNRwcj1/B1ANDbQ6jHA8gtnDoKoQHNriUUpBEB13TtCO4av/y1rmaKN4
9oNOvCYlz5KwwRQooQ27b4UzJjAOQ22V9uFlKQFkcSs8c+vUERCM5tr4XdZL6vTs
KX5Ur1H/qeoJ7/7uToulJyJ9H/vL6u5pp1QDlhGKcp20EGSPkr6smHHBk0PxHJt8
SerNGEAnWI1yMktopZKFImuZb8PFrtHvZ+3emSZMSEqHPqxlDnEzMplPPK3mPPcQ
rmtm9TFtaEKHXCq9IXhSvLKA9W1VrKeN5kpNaRAZGPSmUo1d/tzwDunBSODYefFB
BS8ufMI60cyNflpTVLNj14ONTxkAxl0D3V8ck8LO2gi8YNcx83zjCXVPc9gN1/T1
VwhHXPGjDUku2QPqRKeWzQb9zon6SY5nEueSCNOjcW2lSY7n6GUe7jIYbFgcHQ2f
SW9hMlqKzJE0YAHrbKA0Ufyrm06baiKrmyfA+k+PMV72IimnBgBp+i5CXmBa8CpE
dX/ae98ueGb7QSdj8q8ZcaK5s2ELfQk2PXRqCO97oZbMu5325ELnr7zmN/LhwYSG
2gGkUU7WIxzK3uGgmRlHgpKAmaFH8e4Yuzj0xtlrBYOR3nhL719KNU4w1kN25AVu
yE//f7Ss2zm5Va8692WdwLtgndNq42ikJF8WCyDN6Ss/4xVLRqICCOL7BibBiZl7
s/qq/WgxUhYwlKYfaZ2oxqRfDWGhfdxCJxcwyGyS04c7P/zalJo39kT90KfVKRhF
dn+fASD6JRUP4PDrQf1PjrCys5drUXrXlaE38p1zPIi0iJJN09OXeoMP93ctlj7m
+ej7km26VM6A7DrzShW5oNzaGK+SmLKVlkcEdHRQqxSOHdubzYAXyCeABOqWoqAy
VPaHPtswbRPV8mqgBtVG+q/rRuZmofDOrE7ikTKGNljDrKN7IqTaCWMZLo97AM/8
+5vTaTC6jfJ3DoTspVCMw7Sk/0msfQZ11hGfzux+ZdBEBq1nzofpzPDPLgRGcbv4
aoRSkIYp/72GzvJUhdJKSqqRmkI1aBLDFdIaCVifs6WxUy2xkq6qakzKWtJiJbVS
8es8AyPbcPYMx+pGKphSFCvNg2sjpub0T2tNoO2YjI5J6T2ogXZktRDU+loL2AHd
8RcW9rR6b02C9f5oM7TgusCFAp5g1e/wqIAnLQlWEFy9sbkuPHrj42KTp16ZsbA/
vabPW1ALySDldAC+h3870XNm6GOH8rAa93VLG4WhJHilWAGvIwT33ajLiIcKWhJ9
so9lP/jIv/xgx5KKYs2hyhZ8aHqUCUEgOTnrS8s/LAqDrgm2TZZdzyB5/y3DQRP7
RSJqEgfUwqXkHiulex5asd1WahoGW6BGMbf5yabDHpmuQZvKxhJJr8QsxD8QXzuO
DQ8X5vNr5/IDO8drMHDa6qdQbhB5YjTwCBGePj/6wYW+m5rfx3SA3N2Er69AIUt9
X2g5vG5ZmVOOSX29jCzIE6M//oFfspCJpFY0+gY7SZB5+L4POX7LI1TI8b1CkGAG
vgHeAe/ATAV1upiQVidGYyy/oJy/OHsN0W6HE2P6WY5BDXxnVb6dwZiPL48M5tat
1cig3zR/q7G7NTkuBRNC1XnmDUD72WqhnovR29d+y2hhWTtwgET/fzVe6Y/QNKV8
JHjQ7uvLCNENJlAj7IahoGLBww7vglqTyWjU5FFiaFRFf8Ij+CTYjEDwxzzuffrv
NSJLp++DUh+jMxybkbqb+7SdgJamg/Dp+GCOaLFUVkcFMSLzPasPFvyLw2jCwPB1
k9XbvP1cd3buGjRLq4xaD8gzJw473G/vH+0gQOEarluVD+AkkadyMtff2da5NhjF
7Fo29MtPH4mFNRUCFL3+sXSnCl6LbuQPKHJMgZP2XUNd/yG70mtnATeOS4zI+rnG
01z+hK0cSRyeCEMds6+g4in5/ldkoWnnjTnQyckCv6SUkKvz46+qa1o/Swrk73B0
ZxF95ca5TYEZnNR9461Te7NOOywsAh27KRRHK13+nufsHO0Ns2IuHWJsDKnClQnC
CudH6EuZEkhLbuScx9Njgc15ArZppV29JaGw8qzQUZAMiIktMSSauZXSZqS23sIg
GpGRZFAvx9RwZRp9Cvw2zAeq5Pf+wkiIu9xFaORRrhSU14wUCy/CDYmVaSxoWmyv
vJzfrJkYWGhSj3RwU/SBKNuwG/aQmdNA8zO9VWLdCF49KfgyKCC+AVs2Jbug5hwm
Om3siM/gI5FwzIpZCuoXc6Ne8wZqumNmQ3TN3oKzl+tu3uUuGqAFVcI1FUPH+iUF
DpV2FGnft3j0bkdwS0F3oCJ1BeqtOVbVPPA6uj3vZoL3UyDUaGNLq3SlzQpWituj
UgnSaiTU3/OfYvzFDhuT/5SPVWrCUQFCB2xG9cNz/69v0/KURqKhKSvj6oKHpwAz
qPtfJ1UJAgytJGl7KIEMrwR8X+jq5o7tWw3DUEN9lY3SrC7zxbHUt8rYnyGpMvwT
TVWo0IXrNt2N0B0waLuKKyYj/WqK24jlJp1Rus1qG6fhzfzG9tEcBgH6cLiq+FK+
7BtYDGKfFa/yIWLUntF61JsUt6jYMLIhxsehGchXIUO71HZQE5BXdOttgGvJfkb4
Hh4/N9+NRAlRxk10oAXsLEfEK0JNO0fsDQgcOa+JH9S0XjUBAYof7XkiSeS9c6Ph
t2cFSOyrms05+856/5hXzbludI/BpvmfqijIaQ35IChksG3CgFYeAEK00C8zk5Zf
NuUHJcAFUCHMnTlq2HyL3SXh8PcaBA/q9hcspSnL3ej65NKj01tHYDst3fekD18Y
dKeCmfaUl8yURt7p2TxijPyn+7UDq4VueDJUw1v1RGDxwE6KCgnMCqQN+grVWw9J
ZvGfXW6VelULt/tsra4a17zDp7niFTNUPT0p5wDrO/qQx1GZOhXctCrMFDcZqDsN
BAgAH1bmctxkYQlHPBDt7EkRuj1/I0jNPMt+0yMznwjvwsImKiPK+vhielLmK4Rd
hCbgSLPA1NFq61r7a2gf85+a/QG0QgQ+TDIXDPfv/8IlyDMqmfRzkHwwPgZsc72h
EJL6HrHdF0EkXIIitdaqEFMkS41BbluB4Attx3WUE/33nFSwmHVhEcZUTlYcnTbz
7a4NiskGfKdRzmP9EbJIeTrB4LbPiBhiqHb5IiRpO6qspZM9akmdPWogxwjSNgYv
MzOTzFl/in/WtjusfgnptAGB4wWhUbESSYPSKdq9KUJvMuESI8Fko5TqOjeyovcl
0o7rcCu0bRjjn6h12B4WQd9r+gxmBVBlDVRUMf52lx2inKYTZYJFMKy4zy7UFPr+
VQJEPX6b2pWEn7hO1eRH5M8+zTecfFEcwp36l09RwVN88pgNp2X5Xz/1ZtNuCeCF
L4dHKWQG9UzpSSN4yWivWEeKTpiBT5ESvA6sAhhxZVKP30H/HUW2bsRl1NyJ0aPz
uzbYmEcWNldQ3IWRPMmtSWvgEcgPCNsQfJEAK5UKZmh9aD2tHpi6vh3SVs9jEGV1
PwLUYH175yBkGjWYbqJnHEALZCub4h+g7XpcsD41iIL3En6oGEIJrhbWB8BCXRo/
3erUx9xDMyRi5XhMxxvc43uBP1edhQkn0pUnRpF+Ql6jdkqibpp2m25EymNhKb78
REXw7QEF0EVNx1GHauQmnS5JP55LcJUCDrgMlaUDAg2xK2xyHWgDBIYJ0ejQ3tHG
LS/HArE5k6PvYfAGV/vLuseZyEZ9JIVg5/0QfN/MP6A3G0Fu/cAQZV2ROv+wses1
eVUsw/q+cM+jnktirZNYlsmdDz6x2FkmjgLXwxTP7x/YMylxnz1M4T3upYUoGEQn
gTUR5bSktOMu+IoEJHIUZVWKLwrYXwwFiT4D/T+PwWHfGqZWgIivWx2u3cWQLQK7
YFTpRCApOn5m4urFdDWI0vawB2M1cBVB0SitDKtdMZwIJH1NRoaAWpBiLuM6Si5p
KB8tMVYn0CAvPlD32bCzhuGJ2W0g3kDwNS8w3kQ8H98G079ajR3vMuCwvbM5KnZJ
rD+Ob/+N8/qxcVUrDLw4DAr9S0KIt/pBA2uXXeZoxE8yiT0lBFYgTIEHvPXj5vwk
Apqm7BVtYskP77klicknZi3GnoFiW/n8zeSNtlSlstzeJ3xrneKm6D6oxC66RCoD
DNyJX/j7D+RGWsaSiAF7JuL0Z+TtGUQFzQNY823PA2X+jMXlxGrOI4n1cTLXkra9
UWRcG7dDk1Z1PyY6/qQgckFT5h3QiHQJSk3t+QCRVFHOKwd/QfbnaqDn4DD94e+u
WNMXFJWQN/2Zda9siBI3CgL8UIGlV4XnxaCTOtZLL8tPTzjHg38D3u+FJaD5sqTi
Gvrj48OHaik6tGYK7BCJ41SG99d7jCsxtu8d/Y6Q2dwFC7dZr05r3A8DkT6XpGXe
9Vy/i0EE3WNqgofu4k87aePNbZuhaMt5WCq+eHhtaclJo/5vdYFNI9zagXhciN6i
102YIrSCK7JMkyYKAsqAS40TYdbEOFIcHC1hG4s5vXxQM0eSwVz78gwS5KvYOxqG
YByrTQW8T8NDcXQ/03oglVe9jNw5SHh1J/amJtb/Y8qoiHh23OywJHAeenHvzSkZ
TYQoH4Z9xMdGpZpZVK9Dwxt4n1f0BAluqEU+YCxteLPKP2REY/r6WyK2fa9W+oJy
ua4I6nMF7TY/dp1jeM5WaX+hXaQpoRAbtMAkpe1OIET7RPnVJDdPT+EPbtZx/4da
2LEfT/6H/evcneXp1jsBTngO8kIf3Mgbv6QWiKCFoesKJOP7kPn5+EgGdmqoyVZL
J5tviWe+4cgHwN384p2y/xCE3QkEdzYgehPX7T02Rqq5kTzg0Zh2BJDiMO9B4Asu
A0jWSCScVRjvXWN8sJU2ddKvqu2ylb8GO0+HqjjwgRg7PvUtuxhWTIQDW7PgnvL9
Xr0RQZRJxfQxMKWXAEG+iEylgak5x+uSCDr+iQ/s884/FHjJ+tBlV6X6Z9ft3xra
R2bMM3ZZt6qzeldQnbcNQEuKIcna8gR4iZTIhlFObkfFniMPQBNoV/vRBQRaRvHT
gadsAblNc7436szTZbgO4hqaNM00MIIHKcGYQTJgO4YzOzfnI4b2B0p2tsXBONs0
+bUW6u9LC1YhzLccW/G85U3d8x4Ed8BM0R2mogUtlJOuXCqYJp+4FERbqx+9LGeQ
0GyXthH0HwX7Hz2hvDB0XNNscFVTpq1yL6CBhIaz2QvK+RG6i/cdv7ifhXj1xt+e
/qM7nO69XBqyrwOprcPpT0zlFrEV8vVbKjq4YuYTPPdFlw3aqdxcGWlNnTOCFEGs
nizjMvbf5PrZ9ZCbquOhKyfY84nGKlfrxtYi9tpvmJWTAKo3fOC5EuiWvHi6DSZ1
Y+A6u/BCI9SUqJNvNe3wNCeCorUKSbm8mKamdd3d1ThBM6tHqV4Z5uOfOpWAv9w2
eePbjLne6ZEPzIYDtnQLgxyGttj758DQchUyHni6397lC6vBc13LiYDfO5mI/2wC
PS5GnzbpenBkIQj7kAz95SwImk4v1I5opO8eq5A1MC7JIBPC35JEPwKpd6ztJ741
0LW6riO+SNONBSck946Aucov4BNvYkBNkPbMSx5vFAmM3H24Rpu1JwVq0gwwNvst
6ovH8eMDo0fZmIXoiT8BLoEkON0Vofj8EGoTu8CoORtkFhWUT7tJCrzl5uiwOLnh
NmNIlyrJtDV0CLNKke2NDzBl/T+O1EIOFRsqdZ5FqpmaR3UbxNymG9OiJ4i0jkZ+
Kj9F/RjmWN2/ML5RBbEUE0vQ0f6BgSApg2lRC+wtdVhW58TpwjBn1FmkKBolCMm6
ieRzo4QTDhuCmT4sbbc0cQIli1HptzdEQTRIBv2XWnaFIJwl3ElQQB4gbT8++Uvv
Q0LMVZAv/zw2aMyZMujvDwQZSAJAPn5nwh5x4U1a1UKlc7unBFEjuPpCyTFwMVwk
UOCXRMe1Sv5MkSY+ww5xHSzz/7qe8b5SLjfOlyNbvdz/ZecAh/iZ4MizL/vCMx/+
qKHORRzPyfrG3hggfHziSuPtAzYjfz9/4/rrBHeF6a5SA6ewLqPnGzOQlr505175
BRbB5WzH1gGos3IDifynjmVEe1Vi/HPL3urUXqh0Ju8rBY3q/DsCgpslS0ZNp9fO
RocJkBf9QeUVQzNAtbX8Tq5EYO4C3dEMLSBlQwQjUaSnX17JGrFEL8bcaTU4uOZM
eY5Za/7wePfFv7mFlIaw3Fi1+RaLk2FGmJooNBV5u5s6MVKIRmJ0Kypyr3A3Ra0d
lVXhLNSk9yITDilcTneQGraxNwSuFgWztDdAvDoRtS3gSUzGEpQOKNqIUtIBt4YE
RzPo2LuvsDr2+TajpYUEqd1XyohXZWtdQkybsXncNnfBFaWGQPtNnn8YP30vgqwF
vzSCh/H1t5W53CsjoHvezeWfDKp66KwB0sz9ZLHc5kz+Z8Sd/FIoL2kC+lj+bNq7
qYfyzrZ49f5qzFq4itRYbZXZkNd6wCrHmghTKbEpdu0h+Ifz2jVKNxNPlU15XdDc
PIcJ/ZTnru7tp5KkBN0mRb4+o0Nvm/Xit+UuuzsCzVAB6qPmSnfPqWfRm84zwk4b
lT3SIvwm7shRycN2sPNmcNqKmCWh+zm3cl7G0L/3esysuk++Bk8mjc2bPQUIC6Nr
lLCS/2cje4e+0XW5Pq8xs+EQ9Z7cpDq01ckxdA0eNcDUnE5cgMRgQhAU3L7S6b/s
Os/1Y4UJy3LA5gZUubQGnsFJyNp1c5ce/dI4RDxhQtojPNUpk4Dvpi86bP8bhRoH
MTmzMGn4zWceaCp55kJl2t7iUIJbdYSuEkRKmKm+/NYXwiLrV1dpvNebuX3qWdSc
nhYWd504yZsxp67wKQJI6p1H/IB8AUfhUUBrliXcHj56NSSP2yntm1ogcKpyWTQC
Q9eTpbqqCWtxMPvhXyfh2oKgMa0cyu6EoeEkzXtN3tbiX4tSivhTdCT2Dl5jr1W7
Js9gDH22IRHOQrI1Mr/kehFiGz5TJrOrf6KB9nCNBgyskwzeRrH608dzf7//N8jR
4dqn6AcKObavMdstR4M3SC1FbZqphqBkLSYWzL43G+cddx0LNOJNeQKa6C6fZwk5
MdqANgVt1TBbjIlPY6uKQ6bW3l0ZZr3on+9gwI5+KDmWHH/4EDVRB19vvFaKdEiu
ItA1A4WwX1h0PxFskimWfx6tIMi1cOx/yRwIArgSujIO1/2f63WudQi8h3Plz/rM
MuZEhfz0KIP3d+YIlfpMZUWHqMr1kfedQLG3XfA8PmybxD75+AER8BpGSPX+ephZ
Bq3iy4auQvTjXW3R9ID/gxx7veT/j8q9XFg7v25LDHdr8kiTK2HWcR2dpfwcrIeM
nbWV9pZarvmRC6vkhtqIoHxquBtHI7GfWpmb+Jo5LQgcWIvvwjOuCTUtMNluiBYM
usKWmTyEbMapfdYrBVUO2mkjIIRi5MRypwvV86J3NgAmC7Il0tRqJQSF2IwyZ8z7
1DGxBp26RMKyMzBKA8K7YeqrpAAy5skjUVTTJ11hf07rK/HdzXS+qIkcK+jTLrFD
aPROTj6nrnj9Vw0Qkfr778klbrJ9Q2A9TmdCMXAiIz0AGhfnTPidHLfzmLX+RI6M
mR4Ir5inDGM63UTUZRutxWftaZaxmkIzQwALSmN5LpJPVwe5OGn8loeI0n0EdzcH
oqsZVdELHba0W0H7lyhGr8ZpwKcoAQcsBR48ydZCDGtmhIgRXeEThA+TyIvWS/Py
GNoCLb64nFWNlAStOczoyR7uHFwFa7UHQL9CSQvJa4nc8DWNIylkAm7Mo1OPePzl
TuMW99Av5NdQQjT5qKivjwX3quBEteHCgI2cA4owVWBJb68Y0rduFskDWjl1odde
aad+TYThkrnGD60kCpH2fyge5qRc80UuVgWnFqIg/ELZp8XwoGwDk1H7f2/YPuuz
vBjrvDJbOBrcPGfKR4l2ZNK42FU1IQLwxwwuvvEywUCtFMvA/5Je3s8rZ0SGAfIA
adqVwkCW1u8iwZh+RcOjAvbXn9mmH5bX0gBBO9y6M6xE5BAkW3e9X1CwlKk/d7J6
mSILm++EEiUF7PhhFH8LEu5j4oGAzVSxIfRIclw9qLY5+LpIr1s+nmByZhZYbft8
cewPXrrKcucJ02H5TfWrE1o78xMk+Iblphiva0ct5YiP7SLtcHxSseeOetFQoyBX
XZ4VKU9RW6KqDeCRdW/huB97vip5PWL2Fw9IoIl6/1tIHOLLREmWHsMnQHUeqko/
wuto786N6t72jRGVIrfyspRyd8X0T1qpwpd8wFnP5vtdgxnUbPeM7Am1/ODS/N7q
aRynm2tEIVe+xVPqOc+Hph7J7i/m2RO+sSloW01+OaOQN5odXpfC0RfrBupC9c/t
QqUI4CMrnv2xs4m8o3gNQUlmPaCeHc9DXjrEWNDmxoDjtNzduPOXSLVVt2mW/ctm
fYXbBelmDk/s8P/L+Ji/aXthauIXBcQBFk0n4/5PGcdlhUvgmk+uuFTTC4CpdZGV
01x2J9P8IHPpev0ikQjNspAH3y/nX71px4Tn4DcKxEQDIfoAc654McDDHi5sg9oT
5L95z+sBWzdJpqb/1xzvMlFhN4N6ugKKohqDgNCYj+TqoH3wkw6eqFW5PFobZs10
cAL3R9W1emPX0VV/TKBvvbxXO/4ulPMGxn+MB8AtGGVVgSrX6rOy76ET9p2RUIhI
IyITU4dIkjcRNjwfBCxMGNmF59UsnVyROtRqITIrT1YHxCZf9IFt0rdovVIr4Jsw
aFdLZTxHXThmProG29KBmyHiy2fIJo6ixMDjaYJa4G2drXMbCf+d7L4BMEoabIz5
j0bZGWV40nguLNLruYTAJUfkLmUa92qQSiacNtL5YyiM6AU7MegvYZiZiWHOmSSy
YtMbGZX6xt8F8rNOoH0yJk9fupqLp2IjzI/uS/OuXvdQMxe+AGFVYo6Z1wPr5A0+
eGf8f7/rXZLVIHhm/sHvRlk/tURmcOHFUEcR8Hf49mk8FDg02wIHAXipSQ/0g1PP
lOsoQbr4q65lwuhtrqEvb2/5FP5EomWlUjaFG4Xd/qFttyfIoj1Lk4fBj6pldDv1
fH5Qi7XFjoXUCtVeEQ6G7hst6WNhiKBtEYSTZYppoYA8ihlJj9a/rr3LrzFg5WDk
QqbFn7+7457YvZAy9gPeTBSsv1WCgzLTCTGGzie/AKjwPx62qYqGOx3BrSB0Fpre
dFT5ggE8qbZk8bUcda17j6pDCeJXVyz0CGjI/s+suVQHYAPO7FT875vGVDImUxEB
3A6oSN4zFjMBbmN7NkyNE6/0n1pJzZ12h+XNmRakNO0HJ20Rafim49TybbOKhoVU
PDixvIELtbKMycERGu/u/3ncXDPJbnoJVa8MqDhz96lf3i2itqZVbAdc2wePXXO+
1gXSh8A5lsr/f8QE+RkcDPhLEvmTRpij0HnruTKWGmJhcYztlwJoRCiyNMRi3cgx
5V3hyt/VSARiH36otv2LqPmlJTH+cImCHYOSfWdtjzUPPin0h2Hg0QzLp7lr2SgZ
HK5a0xa65Pv51clbzC7z9jEKIlu+N4aTdBQXcBNnpoBZV/dtbcsF82OPbI3/IoOd
JcbaIGUDWmjlcijpOqLkRsaMRmUM7Y3++JxH2WHTEaVaAcuLgHNoNhuV8p8C3RqP
nyeZjfnkkZoKTmlUC+k/DMPGq/QlO67E7fcmZxAsSe8T7UnBVKn6Eu3VsR2hmN3i
VoJnBSSujzfHQbOH5OJV/srsMeweGljZ/A/2ftc0ndArWDUmoSiD1cYPiP82iF+S
D2gAVi6rdexyyqBRTEeSMb4JvPIsZoF4ASO1Bx9rIIQBuuS4C9gqbPfSMBcf18wK
+5Ut0vll7sBij797Rhf6iZ+A2cT7y5M3iyHH/iFvKF/3fmJgxioqJYofQhrp0lcl
PTvFt+8EDea/J1DzyLKhxsLQcjvA5t58oBvYOuqanYkQD9It+31glYl2sKRy9jbz
BIP51pGVU9YWs6v3H0WXt4sYeg2hvSBMuM2mesfMbACDqlQUwh8yG5+vhDpx75K8
gBh071vGPCFCILQZhuRNvpOgnqImQa3wogZC+V6QiiJerCHl4kXMj7P/bJZbvY6X
2dWzsGu9UxDtC2vvVaRL4x4+KC/5M+vPgjIm8OeNZ4qD0ie9d++9TTEV3y9Je5br
WDPhCjeMQ0jDmbl+1JcyiDNtltss6IHJsiNPdgQGH3Z9sPvKLKkmAcmVfXYVfWny
BoPEa5o/Lwpeh+34XRBC07AcqmXLdsLiV0l0/K8/0aoyOg8hS1CbGNpKXq55guBN
vyyYNK8U+MsVobRH+kuf0kD/NikPtqJUyY5LiG2MjJ2ABL2HxE+YFHRpUiYcQwIn
IbR6qTWsL/CABpPiLpD3tXswQIYCGg4qIHU9AcTdUyCx5Wbhu9tt5e5kl/OOfrZH
XQZi+33P7OtIh1BA9eH5PxbKeQSHTE3hoo+isBLnoH0aksIGkOTmer6daNsDZUOK
RgLoprXM9xxgM1Elc1dj4+UNAAbjv7lI7Py2STUUPxsJ2PFmZ3YUnEJlNk+RrxmZ
JscFFF5E53EjYVYTJ5/IJU+WwkIk8SX+1jW0mxfX1VUfCwse7GmHqy+GUqmZ/+ZX
V63NYsHw/3KFUGN95ZmJ8ebjTDfhKkNBd5/SaPBo4StJvnOVHdXngUKlgeS7DcWT
PgpUYnv2qcj8cv515qJbjdmZMn4Z3Xg2vi1U+btap6zn80U03RUK+OyEXXPzJjor
tujFaHbidBwId51eSat6xEcCHggB4u2HFyZb/og/PyLxO0RF1BLG35ZJAhlFKFvh
X22utPAsL9Td2s0Sxh+Esf19Ko9kEITNGiwHN/kE+tO76CDQ1GhFphqUbhzVhki+
t0lJRAQwcRowJ7yf5rDBCo8cEVH2EykXlKsmAQMEK9bh35yKrtfYqn88b+/5ytju
Y1tmyILDi+UGkFy2I3jcmJdf/qPTXSITdKnSkX1Jcok3p+48MDzj7vIdWs2m96ra
YWw2HrksQRVR2pqmMsCURCZQi8NHiS4OFHrcKiy526NSGDgUxO+JnbbdxCeA6RgC
9PiWq8XCHufhHpdA5qW3DXb8cN+hXgUK4eOi9uDuWK17l7gXpofkre7+/kSFf/KH
muWB0w9UMH5Zwc/6lqAMBT9w0RHbZO4P+8LRmOpiaPpaWHY1EpzPEMtbDezKucr3
V8RyMWIUL9QJm8Jg25v/yGr3uObwDaGhMSGW1sNFGBZu6rsCTjjpTdnSWTya2WpU
ABic1cvaF4kR4fMsu9X+2ZdBWWdCliiOkgp+GytF33oupApKFClwj9CvZZ6I+AmO
Avc4WCoyOsZGJkFAAbu6yR3g1my0GmdSoAuuXMiZujQVgMUvzUAQSE5cPXIRvAde
Hr2mPBUPCHwCSy8HBj/kKqz4YoREb/W/TNB+OJa3EWtpFFCI8pMdVIiLTznEYUMI
qseia36Zijox58YfWtu67YWcYENegXHzEa32MKaxXjB4+txGN4vuJbcVnN+olOVe
XIUci4zq1o4lLw2IS3Z/Mq97sOx1XeXLgYmfP78br4f1Jjn7oEeGE38QY0kHdVRs
fz1Z9KlEY4xRN1azPP+rHmjgUsNV69gWmfignoixN4Berzz6c0ZoxWq/WgisvV7u
Jl7ocDwg22M/RndwX7S9xJOE2yn1maPUSIsmBKD//B95J1+A/OsFeGPmk9ouDJCI
+nPWUxvftYjnns5WIzTg7BXIa9PQk0JSDE+pXHFC01Z7hiH6ekMyJo4fpF+uYpLJ
F3qdDGj3J1i4wLTRAuw6cGGwpJJ4GD0RKj7BSQMB+pc9CXCs31rBJTmN+1TMoI3M
c7epsWp6w/nKvXFgoTu9uJvstE8Ou5ml1XF88al2kA7rGPtdN6SblQM8L1pfs090
U3I2ffBGepdRWhBnK1qPbxIyMdG7TEsXVrR10W5+oP78CfwW7GRuvGCHRDERPPmW
hPu0aSWVKB4n2z18o6HHn7MYxf15C9icf1FSFl3ZrWvSkfRFT3ZxdoxHEDrr95X2
N0Tz+o0GQt7EINDEiYMk9M0kIOjktN+CcFu3FIjhiompbUtJM+CumZK1PgkKf5Pc
Uz+pYKtTs1RyhnevI3Vmz6lWpxPhUDLiq+A8uapJlTdS2iJFPNdWNty08JJEiOQ1
+gnHe96XtHg7L1Ybdm3K3xr3v3zJP6wS7e96DY+0ZVU0Umsbg03g4TWN6vbHOvBY
O4oPNPZMde5CMH4oSGSrwtQwHSTtNyvHiM6ASe4Kxvmean0sUJwo/g8a2NB8Edod
mnWRxnRJdHxGTopDAyF4hO16gpKHY5e7CUt1nt8hMWxIl2VQ53dMmpiq4fZHBH4R
KSxlXG5otX26+puFlou9+PGLZVNzhcZWUA/JIB9dmRG4tnsNRc6+p8W1yRJutzVh
Uq/poFxOWpmG6Ox/f5pTHzn7qNBKAZ4YxQR4NUtc7U5IjhK7bGmBW+qY4knn9JDu
9n5sY9klwur5ggIyk6RZaVFY07Os766sbGEhzyb0TaNCvlPJuyp2MDZlZJhUaiht
T84H72IUfXpD1JHSlH+wZIqyAtmf8+MfVfvGWgdT8tbgJeBLBZNT6Uj7wE3qUMgc
IrpTluKHvagPGhVms5xicHE5z0XXRB/RWeyOUX+xwzr9gVZvpzF6YxMUk3HOmtzY
r6aNL8ClrGzXNLMz0bHgCsJzC5291Y0P+AsLNRIbGDUYbUQ7fB9Xj49uFQtQUoFz
KLGiXRKhgwWQM4HRphHmKgHrXAa06AgQMe+rLKslzpaNGHAvL0/bansyNuQ+yTNr
nEOTYN7ZLgTwSK+AwJ0NLRfVSOkS6VGu0JkQ21uV8bEQcSHVqD34x7CgLRAAfucn
j3pxyHT8POD8TbBh2fj2ZZDAxucEyaSMZP+6+KwgTWOWYgSkYkWyBYM8JP5k4hre
RmWFIRdsTOWPBQKzWoxdonmoa89Qr0S0p2iftOZ+V8kfWCOZle5oWEKg0qvP8r9O
n/AOSq1XUe6oK4to4pRUVDz17cVtIm5pbPUWF/X8P15M+1bpNHUsEOOkq/qJdpCm
fl5lEbXL0iKIuFLyXYiBDHyGnisDr7s4w1T/P9wIXouFc/I6t1LHxFla/5lxA0B0
nkPX2a82AjhdJEQcmJP+AIhnwzm+8Fmd7gLsefyIV5ddm7cY+M+WfUBrcJWZBgkB
QggqtouCFAexblUSUbLzxL9pryeBQFBdwYApMlyp86bna8KAvcLlR/gmOOKN3ZHu
16v7VsgDOvB0MUhcY+mZ2Y4ibmwMtGdf4DsK+wYcPDa7+vetKZeMMx0b3zm/Wnty
FjHGx9nPyjghYgYHeRjmpFnwA3XsxqTlLUUHJw8+RlTC2KwHZw0BSqLbjddpHg40
j8ZyTNfClBovL86wYaMGTN2gpN6Xya6KYtnjb2rgrAt626vzP3P9JYs6YRwvW/yh
Qgzeb7GaNqpS4KfXRO75Fc/r6bTDwEYNzy22m/TJBKzbtGgCZYTtBdqoIqBd79Kw
5tMHnQ+3Xgn4GPNo+fccjOBkAcY8SzOtjdaOyZAn4OOuxHglPrWUrKq/ufouoDLR
4aITxfQy8CvMePs8hyHuNYPc6es9azqQFcEo7keBIv1sKen0ESDmIcx+d+mB928I
qbMzE0rk3NmaTOPvEebmc1y+bB1x+i7yiaCqSDnpVxoqC1W8gu09wTjsBBtIN7U9
saVpe+CB1PjsuCnHW9/3olbiNAPCBmhrwIPK14Yct4eMycy7BdCuUikA+GZEb0AA
EVQ/4U6KrLs0M3irpI3B60TDvolpx6Gv1eQSbYPD/QD+Y3QuMwyXfJNK+Qc7/sDd
nhNK2h+dtqQ0mwiIr0fYrXUQmjWsdNBD4qeTxKuOPhKbhJQvjr793eWEzx2ZGo/l
GZZNE0ueeHth9G+I6GXl8iNleNt4PfHlLmJn/SnK4daiR6eD+NZJYjrJ7XAShrwg
nFt1LO6l1DOcSLHdXfDCzRF4aerl5L2Mm7uYfccOSNjDqeZJ5nfCfDxfdP2Euhhk
UzW/OaNCgYjkfj0IVuWa7bmmu6eGywlgkqvTNHH0BVJHItNtw9X/bkVOsfNFm4Zo
nWA1/HO9HRzB+C78d4nUG+X6uQduamSgrIfy9Nb8Z0jsquMW5+yZcAr/wjml3+pZ
dHV48Rn7m9z3IRAiCHnOzFHiZPA1ABFTJg6bN8QD/xNKhxGgOo1CImb5kSzbtYDQ
j6E9fSg1JEYEEX8Irn2oQgJFFG3kUs+z42byeLZmv33rpCIVqc1CRVaM2RQ7qoQL
L3aoZzjbqBwBTkcYdS5ZQIXj2FwK9GZT3r9mnGa5J5pLUGgTvZ0Sc5AX42MfHQGr
z+Y47NQ/v+fgtkStIV4IVV7QfSM1FRU80Z5fIvoy0fmkY3Jrw3W/YUyT+XKBbN9E
tWUWLDpCRsr0cEWTaVA5UdvXm6QsRkynhTL+3Bk8i/W/npcYLKzHErRokS1FHfF5
l4SRnIaMWgDcT1dIPy7MkvcFYMk98scxLxSd6dULElX6ng+di+LU+eQemv3xfxCE
Bp2Nyr9069kESac/VNHWMEtKqLtFQKtlxtHJc5CUf7qGgDEByd2+YnoeyO1lGfjZ
Jc6ePHPh4hcQqv8ydotqizc0IlbxMddNQcyaFFt0CdR95nHhmtd5cJm+dVx8ACk1
xj9JIRcNjDvbCVQ3FePY2vnOYeV98TVPeFVmkSJgQ4spy1GPZ2Z1sz2dhDxbQG8N
BT0cpYAYjJPY6x0TVBNuv6Z2r5QR4LIfbZrU7zNRDjpmuk0nkg5C/Hlz1Sx8lORc
eFE2Z48VuMCRF0DyAOshMiPjHfP3hZNkaenIXe3cKJxq7Sy1T+kDltGSXM4T5Pn1
DAU0obEjXhin+HV7tYAnqIQzEXq2KC4J1+vr85LlbHprFct+UYILzkm+5GZIv77M
+88Y1d1cwEX12kFhj1KfOa8IWKvqplT9HgfMPmXM7FG0ubf1tGC0axfHtmQ5Nnky
33FsVuav+pQZbVw1rdicsJx1PP3hmI4XNNgDqC470f8DRmbqQJtfYwFVWOGuVROf
rD7u1K9EnP4T5613lQdXPCyGr1pb0ktGfujz9+URj8RQOVrkAZHcrP9YvhErqK0e
ikfyjXjJnWwife5g/NLg0GanZHbt9/g5ocap9Ji4ZUli258nqxUhw2wjKJ5Gaq21
T+9V2dbcmhUmf6fL5ymssdIfg0HWqogTfk3KY0rSNEdL5/mzvoBMoG7KoO5Ryzat
LsRgztmuPhJqKEEba6GDziGbKvQo4ezyzNxxW6XVZrnDJXOMXDg2SGBmrVn0IOL8
9eZZxv/Tls9cvIoo9QzkRs7zGYpfdqoeUu36w1UH8WP2/7PNKzVQfEsuR0XhFW4m
HddTeoy6qACDqnN+t+3v6jVMR9hTon3RJ+q+5R/qP4MJry6S8mDiKH9E4pcwiqjs
w6zC2rDJDcR86WVb9gKZrxljdgrMP2uP6QQGUodqLvVS0wwkTosbnvw4ssOvmsx5
ZlxWS178xYfw8mm0bhef4famzRdnzoOb075T3niXhaZpyixTWlZCno8SCRvlPFaR
3EOtDJursELb9TE4ENSKIubCdQxdrtaOp0+BqW7uFwmVDt7R/lfsRkYz4pdj2dBP
lnGugZqWJTHnMlTwKUGgN9b9QCwLqeIS5DYNVDw/IXkr41qcVKJgt0U/87Hdf6gL
850+Vcu6oR0k6b6grhu6GXPIfjj1C3BmguqJFmBA2ez2rSsn9lhDEx/Zz+b5vbm5
K+USrq8XInKQ7LZndVLeNYIEtAKRfR/3HoF22y5G6VhVLz1z/Q5IL/ElbWLLLzGZ
wcC8uZSSIGM7xfTw6M0TEGYTzVhCDIqLWs/9vgJbgRpmYymbKDyV7/4I/ogyRFF8
jLDTbt5JN3jt1U+L3+EznrnRLxSISt/LXPh5bmL90k2QzJSLneHowR8UoIF1xoZ2
oeimBDVEPqxyxGtG1sikWMBvGYkRPv13O45J/GH0rlQfoZMR1WX3OM/ujvxNIoyx
5xs0myBn1S2VJStHhrMuR4r8zhP9iR4FbPyO7Xsr46GFan4uQyA3U/77U2wK/VmS
GBEr8sx2BMhPZ8YRp0A/fHBVXBwYOxi9AMRW7rCCj48IL/7OPEvIBhJWB2yGTIQf
r5VTiK4Fou8eG9uDZLAm7RYC/6d9mzMAc4+ojUjOZFxvEnwpqmLuDZd3fR1ZBDfh
EKF/ml2YfMukLBYdlT0mOYYPy7LvOWn7lX+2F/voKovsG+arFyNhCh9wwrRwTAnV
kReB2T/5Xu/H/zw2cWfN72GYkzYBdqtCOx4mS3nSITlWD1fbtyy2AKnO3CwhB+hM
+fZxC3TbT1S6QinJxqxOGsOjMUmPFR610ijAgbVx3xb7jnkAcEvmgss4g1xana4S
mO1fxK/eelPOFjqK/j6xZ90bLsDmiTR8ZZnp9b3dFIqoScK+YibxViEVyc2KylBp
WCjFnm3B5R17a7NQR3ftbh24TRPmhrndl8oLa+ZmsYZpP5BmAo1QNnoCUlU0Dn2r
RoMH7IbqEogH35yf6VN5ti5RQI9CRhKoyGpg42/4LAFe3nHoZuTJX8XEg/yjly2O
5yh5LL0Nst3XcjxxG6ZtpfwYzyG6tF0B5+D4gWyTelhHKTauYnfQ6tx9gzX4Rujn
pUgxZc28H8iCrA+R2mqyIAKe3UI9A7Bx3TPW4awzDsxmwJyW1LTrPJFFNsEPh64x
qE2UlKi0ck/5uluASQbGw9CbDBgKDv/xWXxA2WujKtmkiITRrZjCQElsryb3eMH+
LgaM/gr9z6vvJ90UvXKlsCp3nzmrBiUtxw9v47RYoEN2xi1Ujhz5fuE4UJBuHslw
FMZBMewwa1Acw8spogRFmwbMPEb3F5Tbl634S6YRc/kH3QrJZK/dZ2VVNkBr6DTn
wVf88yR68efGOXlQ3ojg+Zsw9bAHFNqxsSv+PVp1IV0l79x4h9JS1hCFltRdW2cl
ukD3X8y1eEphKusB7td/pKZXsZpittMzTcoTthF3foufgwlGsWk1nEmguaC3KwwS
2jFivBek98+Kuv+z1qzpiJfCmvzCKpKnjzdle+lGXadQZz8P+7uaLqxM2aVuD6EC
sxDvekGtbJ7h72ngrTVX49IZEXSsYeRfXkO7aEYncFOmZbod9MC8ETV9rIocokKF
saqrjL8rBhIGkNM2GEoqAhSBOLWmrIESMOr1laxILFVMCOOLM8G9r/zILiK981Ga
QgiWbbyPkbZDPAvxOAYbiK4m0Bc3zCypPbRBMTmzEh9GmtoKh/S30pHA7fl4qi2V
uJiC6X9qpljpKnHO1qTN9/OVsUTD7krfdmmJEgtuOBrRYVu/43BDS+NDNuMb3jgk
5eNKAUEavQDZdFD9lEUkpu36IEsycRisXD6p+TIJX6NN8fW3p7miFDwLcq2wPDK0
BK+RtnFluMYiJKMQ53heJOZKn/azOkaRz1ukHs2MudOybELLUCh0Ka5dwaHP4Er0
4xY6kfcvvB+JW3JYYjpS9jdnAypz8DCbSswsISj+4ivzUcqOINYYLFSFi7WGSjxA
LulAlta4dsz2l5VVN81ghfH65Wl1UZO3ubfKj9mocS4oQuKlhkepcuP6+pXabVNi
vf3+1Ol1lmnYGjoQHr06l749NPtZpNgGFJJAjzttwWPXXtl+znroqNo93RLZHFe6
5m2ROw9C6LmwN/uNBRrBLJffqZ4ue2guo7GDIlGubInK8ademDE9MfxxXfZIfbHC
9ho4iA0gv9xuXHIwlvY8OI3/77opeutLPAM0C872Vwju/IGUTrSy13rnpxnsm238
BCHGXdgc5O1K3EGuApNEN77oMs5C8IO+0PNxeVzUsSX1H2hMRnW3ueY1O3lzwgTc
UOmPBulWMaNwClM9QA8QshNl2bdII66Pihj7xhSrgTQtkkaXVhBwA4VaKl+/+Zd5
c3p/wAyqrXOPpiCIeRpTOt+PhOL3wzVlDQjRuOsq92fsqTOvFoHwOmBZq2wzlF58
M+TD+1wQaFEy8pAOISuTqnV5CI/Nu8NCXlq79wbGUf/c1gtZ0ZhWCfbT+oEp6kfO
rwI+DVIdaYMBuuE+LuAwJp/LYp4IsTnzfurcdfohByr8Tv/UT2RgAPXj0/bXi9zC
K2+YnTY8mfaGrNhHGBoaWLMsIMeY7sWSuFUPYfn9dTy52jdj/h2/oUOffagyfsJi
pmWq95Py+Fs/oG8/Vfl6fUgP07dy5ce9KfvhwVnLzAx4hJER/YqoXSFZnAGShvAG
NLQ6hz4Kl3lrvxmfZrhFXjLFtnGNRo76x93mTsHgN5JWSa7ebBpM2GWL0zzGFY9b
J5uIieBvEzuEdoTRkcmxHVSlUAvRmINoF88bjip0WH0ArvgHxmkeQPVW+TwWMIFA
QKU/SIHGGJxfIsuo4K8ssj193aEw9MJ51+Dmnt7pmrllNpQa0aq2h+QYrRw7n891
0a1BN+673aEFRiHz8cKd1FJznWu4rBw/dDAhyE8BVROD+wm0TXZRH9gLweP+fb49
Fmp3dLUkpe0vFqOyDyWcK0QqzNdMr/jnQzIEmqKPIizQSaGLbsuEAn1nBtS3NmHl
i8Z9rOpWC1kT5Ud+i2lkJRvN4KmTwZ7WrUZIDmFY3e2Uo7wzAp9tscq3pU/mf1mz
vFSP5cecgCNq6fvnFke4h3/FKDhgOuXTpA2qUQ79Y5doIzUQ2reHFDONFhiZxdUx
s7e2KCnPeq7uu8KrfeYGFkAe9DKBiHa16ibz7MMec97xyp72O0yq9e2LxJx0Ybrk
Ob5krOCAGtERnmw5mmg+3PdOggTifggmFiwqdINNTn7X5QLgkFD9kgCRBtJjGmDp
RfJ9qFms0jd41QwEfa8FAj1tXKPxBTIdw9LEEr2UpfI6oCi9/mx2ggpP/UdA6geW
0xB7CFb4BT4JrHy2ohOKC9y7m+QTphSyZwLyyYtyGIuK9Kwdxbd4+oonRO9CqZbl
L/iuFacX8M7UoQ6Yu96Dcgn8TgDwyYDPdtV7shqZG5+b3YEbw4rrfOg6HV8sof2L
Giwzy/TiFxl+jjUBevINbk2fHqEO2hcNBaImy0lZB0LhB04FcoyCfEpCbC178AeE
uFfWrpqT5Z18CckAYos6JkgSObeyoqcrYPNAfdSrLr4Cgz8I7JOoaLaUu2IvZaaS
FRmo1/kJ6Ds8VU/EJfbYvXh7yz/TGasbCxFXgQfFxt4PDR68l84I/i6C7n1HQ6RL
5gJtgmV2DYJY7Ki0yAUHOK7K3Mp8lm9DfdZOmZpBBmPFt/Xd28yaX4o2zEbGU8K/
fVv1qhVvKrACRztbKJuqdkM0ZRJn0KIrmx/SoZTKfnIjaxxkdL4exR8UIbJ/BFgD
oZx9b1PilVXeixd1qwRkmNQFoLm4gVuGGgkzKmsWxPlknTAdxfa8dLbFKcwBRVrh
0KtPZe1LafaK458sJ1mz5BCA/Uhj/E9VJFzQjdNqXNiNJr1O73+wxfmMdhO2xG/u
qc7v/HdqYpEnCjP9UlOL4TAPne65WEBHCniRm+ONQH7XNZyGXFCMQ680w82FlDW2
/3B6Ttqb5jMbCIQNHlf32q8BRG/SEXtnA8VU7/UbP3+tDRWPFLLIwWYF3nTkGT2R
fBn7Bw2UlEidCa2AOsgek9td60526hLlZGdO0WAeiR6hOr25orQEUbKEozRFmXR2
OYuqOThBqynC4aGYIvmXE32n6ftIQWfm49BJvLOghy32On9LVnWt6MDXwAwzF40O
fMcJR6nftnCRT1paut/1uMkIWZAN9Ad0R3+C+PoSWsKpp6FK/NfDJAgJ65pzr2Gl
5S1f68IUAZIduDhThrIXpFiiQ3+KijP/u2t0fmTvUe15owHWWLwU2kBYOgOfQ1aF
+EeuuD4FaTV/JJlWSII+i0IN63N2qNQimXI/K+Tb4lR2t0Kkcb7BGUZbvgChh181
rkezayQnNKOD3WwnBZEI+ocnBZ8MTJooJeic/qtto9Y49H/IIWdF+nzeaizEzFmw
CvPrFxb6hQTs9x8Ktq/QtXAg3o9m7P12sbT2cgj3YUe5KfQVgiJp4V41hZSzymNk
CXLg5EbZNMKBndknciYUy3FdKGnluc+EKTIaIkc2hPXYiwGuH60h4ObaNSVbwl7L
K/dx8nQdVWgIU3mNjx9MLQ/M2OpfLBIXAUYkjw7RHLuh8spBhvbd06cOmI6HBlyE
lDKvjIL6ux4Xqa/KwKRoHnWb3bVwcaLJgr/KNVOPIxM/flPvu9HOmdIQB+Z77JNB
FeLB3yfnpLeS1j1+O/+778Dm2hbxJZzFmhkxBM6BNO4gwLGaqtIl4kD5nAAz7glr
wOTRs1RI+EnKeldN6vOuFPAmRvl1DZr3r9KKOPkutbZgruNjhngCfL1DPknwZZsZ
yxrUl7JntFeWXHuQfgZKw/mfqzo7ijE7ZbIspIfMflebzE/IIWxT2okN5duUACna
xTXt5urdsEvTetsBhAlQeGV7kXsu+nNpstxP9/dC57SgLS60txPfFwBx91ObUspb
9zsfQ4hzSgcfiTCTLrO7BkEcLDWJzlNR0gWUDUBj2pYN4E53egZvvz25Zbw4k9wW
HvpCstpNHu2SEVLBtf5uznWnc/BhMV68i5OZtGwrRcLjS4CEyQaiEtpb1IIQR5BF
HXjRCm8f85gOAFtMkQLLazyLuPH0h3iIf/wncRIwq3MsbnFKLvDwhvNdVTbSkqVf
GlNl1Cd8sbZrmjvfpMO8vzylRlakHbds6FQIiCoAkWw4q6UrBIbiZJo3SHvaFvfI
GTtsBH9UdkxT/YlQ69QFbzqxa8yRVKvFA/85uLanXOuZi7+XhEz8MjTACQNC54ED
Coja3zpa5ctuDp/1Zthdy4eUHti3XxYwWrh+orHVOIRixAKWlASki/omkMPwvI++
+o5nXm35yXH2DoLjypvoMbb+qH/uCXo8VOnYFVFBrZtf/DWf0Mi7HMN0szyPqSHR
YYgZKatILRZn1eb1+eWQ32sjOfzIU9eJ/3hXk9YQiCSjJpQY+EDzn7ZPM3QjpAYg
ML0sVeMF5jPd1beB9vF7j1au+RAgEuUeTL95p9nDtWC5YZNlO5l8Gj8yqtVc1kjP
kGp7/X2nhlxbAtAKPfGOiQa5vgc2zbKKuGqQILXdvc4p9Rifz/FRrnhpHSJtQ1Os
GlGnH2f+PjeHvFkqJuN5w7W18hgELTEtCRAtQqLGqzsjycY9nbG+7uEPByMld6Fq
cxZMfcQfZGeC8UZX1DH5GOhoEphRywOJrh53suD4X7Vqp51ZqdeCpyEbnAVXcDKl
jDMDk8uJci9UQ/GAmo3Xqdj0UBSCinZvKZf4inUaYR4Xbt3XLeMWPGF6mVFuS1X1
wCuhxZXAfi+EUME6N4Ju7D/WMPzseXcKypKtWrzNOwaOQLv1zAVV89+x5A4SEwBu
YDAakfWmTf5t+bWI868QZ5syPtgkpLX440EyyHtOE2Pkp/OEK1z7Srl2ghfYMHpu
I3mT/jNEiABzR6WuHgYzygrc7soI8cOK3obozLbBXGuBE1WNbefAcb10e3X0/WKR
gXkxPPuyyWcIB/MEh4dPZx5GZbexb0wXALQe8kO4FxDzHlhjNOyVriChvqylQvqD
mrymw/pX67hXj6fDu4NUWUElisTF0+K5yGo/6YZS1Il4BPrYtNJfhHa71EEfFsdY
Je/rKI7FoJrXcCsU8+0IyyYHseNX13mPjx1+OjxubGhiYynrWTs6CFTRUw/nWbcd
pieCXO+e6Xzp0ps9TrrYIsAIlTYsI0Opz75voxvXOVhms85qVdPgobOPJSqq4Ehk
s2EC9uPj57TQi4gaLxUBLHlvL+wxrYPqZIlia5E+LZHYmp9GWi7eUL/ijUan9hYp
PUXxdNP3+oSiu4dpa9XWZDelzw91c5LxQmdSgvZV5Klz4nHK2EVjiQ2mUW4GM6gn
8OXw7FNRHQU2oaHfnwwYgFAWYruS22sZJukl2imSo/9s0jchWySuvkOHZqzm03aY
39oq9V7Co6mO+RAh430XXBx7BfBxPvPgP26CEbtNMcJUFRYuUmWf26A796KF5UdZ
hWWzSfd+tomKzSSJF1B7CopHuGXzm6FIAtGjnMc60B5sq+QpAaddLEniR+5esHEx
1ep8N+nMLPeNM99lxEL31JP8tUX9yg0OptWzjNNk4vOptagNj76tqYNVrgXJOmxh
17gW210l1IR30yx3GHOGyFbtfGAXrOxxJtpshwuUfjsUCn1+ckKPnnyiVYfc7Cee
yEDD2MT53o1wsEhMBIsEszNlLz1S1XcckWo8KhOkjRIb/ZYG8/k9uHf67XXeMQDU
a0qTEMo7GBziOSoTJfLacHDCJDwUkLkIz4r7eE5sMVwWzXrNuA7fkDorATBRBXFL
vizuu9XNY5tfPacN2J7k6dDQS46JWMoZDfHnntZ4GaPcBevZwW6nqXFVKuhQXN2D
mvTPFsm9tGzG2wjTiUwQdzEIfrm+dt7YXwJ1pQsqWNRqsSpZWGLfkbQWcs0XwDJs
0qAErg86HRHo/BaAVMG+EN8qx9VZh7Qy4C5AhzskP49M/pGckkMWFQmyp5KApYSt
jwwqtLlT96ilszXzt91NXGYWHzuSFaE1Sp6zv/Q515YhE0g1lE3sy9q/Q4Fl9EfC
pfZjDJE0XetsAWltUt3JyWDd1K1fIC2xyfCprYEnFNKp15JdiVFUw9UfCfMZ3FoM
kSB40sgJURyIT/wxfzl+sA+SSafTt/OYmfZxsYoB/DRFswr4rTAmDCfnu/W/PKp5
b1DXPIW2rDJXmtsxVyEL+KIHohUDXSLwCKlBr6F5HsSArSj0QI62Ce41KlPI+B/1
Eu3ObBXbBrmgECYYj76Qja5S7BSQSh2UBLSW82dbraUMUhwfsefTipCmjTbkaXQy
XrteIBBrJz9AaQwCKbOmeHBGvnV56EEKgCGioc5/Fma+RfBHP90P90+L8BiD90Gf
W8rz0DgpZacPTUsYQHX+r3l+IA7WxStDKvGuBEfUYknJMPVTKp6YaVCTkHwh9WG2
91bhlVyX/A/bpInx0OTf/QEPqDk5fDCV3NCZgPcHVEC1l5FWKYzDw3C5/HGefrdi
f4FbXg3I6Oz+uc+WjlY1forbWv+qK2KWBx1gTvRt1RD3dqVWvvddhi7llTLxuRPG
N1KK3CfCxIbKPSpZXkSfn8XOzZonBLpAZ05x7SBcqL5ejyXqFOISENBx/739boNC
48Wz699EvWmGefKmA0DMQ6Tt1jtZwvxngAIgNgadOzI98SDj6jaPfqaqXojkR+2k
ivzwY4wz7O7qjJ6KTPMA04RtrmfNK9vl9uugh8W8TVTqL6MPWweXyIEs2lq/xULP
A80rTSH+5SN24go9alG1h6y+BYh1rRTDEmufcAIWWLdq6fBDEo61ASozrpfPOweQ
VleIebcxwTkX/phxi3c5CzQE8gJ1J5Eknjocg/2O/rLqYunE2hda+9xdiz8s+qpp
ekBgqZKU+T3ZLqCebu3S7JuL0Ii8QuNX5S5GV6x6a00mCNqwEX+9FM7B0WyqtCuA
SjwoNHX3bOPag+65ct+DSxmuS+zGJMtTDToL0dSWimdiwGZEv8F0xkP1PKw/DC20
eB71LG5knkR91vUJSp6iCGU0CwJLjYFVZPiveULe87ucBX8ZMw7FYL9c76U9PlVd
xiq6pEv+UE9h30NtuhZc506HK336C2HkG1rv1bAMCCO0jPMuS26nX0WRlISiO3fE
LJWrYyNAj3KBikzSrb+JA9DcdcSjt6Nh+ii2o3ws7iPJbI47sTBJigcUy9+8B9/C
YRobBhLj2GBzokd4He5jfrIzB88xLJsaWFU22og/t1bh99jfJzCmM/PRIsvF0HwN
wz6FhWVX0YDVxL6AWoc0yNAEOTsCXL6YHzaRYA68QsHNWDFxXYGrtljjm+QMZQa4
ZCrsAZMYiRADwrpXLXDIsQkhYR5mSPi1usVUpujTbhuy4VFumkil57hPksrxgce2
TBwl7ebZrAq3lqb0H3ddwb5v2j4UUPA2ordt0OtREq61ph/cw/Oq1E37XxsNQFYC
IVqlAEtbVJKKNOKdFcQq4nANOeS5ky3wECxJBOdFHhbrOrN76Bxesiy/rncD/DuB
VrOt1xYC8cEV67VjBq0GUctqtyWuZ8y6AkQGDfcMsild3ci4xxafjbuyzzKJNBwD
br0hPHf/HE6q1zY/q+6OtrgYSQvQRD3LwWnhjnrMbthsdbALU9w1WERyhApsjx1s
NNVIJ23tD+cj0rE19QHxBdC30Ljn1odZkPcVPQyuM4KTFS089l6loZicRjDG03DL
EpD7DkIwQ99ELCWGoQw4OotBXdib1NMohr5u9NrHAVfzFt8djjOWhDf7KTkLOHYo
6YvRHWiT7Y3hIrLDI9frCKjJKUlsgwtCuWM69/svUokMSqR6hy65AujfzO9kdMLh
PXr8oFJKIlHiA2PDDcLkeQS82/+kTb054/7+Vr320neGH+6GiCRrUcbMuD45to1k
m8tr1Vemd6Y0SLioeIKrUF/eVQXv/MpaK6dQYa62jUMgsNannsPCHZHcLHX8xA9d
AVg7msXc2YgEq/JrbWKwbpNEzLEoNBl5x54gOA+C9A7wHM2qdET1K6/cNMOfVl04
Vu46NOw7QxysKFg27X/T5LVpJynCoEAaXtEn95pOi6V+4C5UfoU2HqBYkD0rAWXS
Jb/sD6JDl8OMz3bnIoEo5tDYlQHWJsPW4neXmfpjrhaIrYlBi5r8c2PT9VKWhSr3
z9pcc8KLER581WxOVE6zXuPSKyLb/0u8HcdBtNmaREWXcQn9gZQarHg6NOvQ77EL
+thxiKB5aW7X1krp2nzlNWi0l10ySUcS8Wth5R4tPm76yiyF1pOWLM8qIfEeP16+
t3amn4bdqO2XyIcIzjpDdR4ajH/6y387etRlLAbgKhtF5Hr/IyMQUsNsARF5IIIy
aDTPL4Hsic0J9l3b/cNiDWdV5wCbu+uO8fAk11HOBRCdMQDIHos8GYhj4PydW4bN
+BOUlAr4BwirGbiLy3pY5SBXyY+MG2hMSRXxowqdzmeqXZ1OaU9+/Ysuxjq6orUM
p4dYd7pXVZDzmsOz8hUHbHmcYk+KHv6baHYWUFIVoK1BOMUhmE3+GlF0Rk9iaDM8
x25nR7PZjsiPKP8+HMpM4SXLS8mBLGOjKCaxvYrUJcCY/gYjbQffUA+/A+l8wtca
mBOAIMmC919eMFCSyctzXrY2Y39N5UfgUqOW1iaq7UopnxI/HwksFtH66rqbpQT9
P33JQKKiig5KH783dQyL9/VKJO1/Eazqj/ht64HzSHs0biVWiUAZNmzr9qhGynAP
XAPale6z7E8lJnJAPh+S9AWoBCkO2X8ExorrsCiRrk3Q6PK1SClPcYhHiuXBlS/t
E6hGc2mkZ8tLk0o9AtPkEx73QP2/H4oXFglVpTN3HrkYgh1KUTcFU6LVIqLHmR2r
Nupp8bDBY4bkeyZoAMjuHQf6nhpS4oUEhMJ70Ly8FYcgLNqr9BUY3EHogR2MjK8L
06W/LTHlUnn3NEsk4miaP1lW5H2E/dJjjrjJWItPAAk1ocfzDBlHBHhIy+XI+aE2
Movf496ZlnjgeXEUxJPPM2QhfEwSj68TXPR1FcFvc32kBeG9yuN+jykZJInb7Evg
SbXxkUZKkLmX9CWUh0/mux1biHO5jmcyWVho+liTcC4ZNd/nboaw+AU0n4kvI0vg
gIhaEdH92rePAana3wPZFpqbaRkJShnHQgCt7LvFthSixMCspUxNLt7o9CQoIiOy
PnnDb+JRJcKIwPsPMQUpDpnw4OSpkITcsUQ0pvvWdJdjStOYURIBzd77ioVbw6bR
7EX6ugYkKCyTFS4oMq215NCG418N5KQHAyURvxE+J8sUgjXXy0mUxobt7jJTEHjt
L9dptdkzE1U8IHSIhYphEDdWUGoDXdMqnK+54CVacX3vgK2QRmAgFqggkGz0BUsO
cU3nSpfhq+6MQREcyF/m0BcGClfC5NE1s8dbMEOfeC6QtJL2SKNOax0iLOSgzEgy
di6yC6t49h8Hg0hiUpkhImCZLLWaJwFIUyUQEz0oX96DRnH0mYMJjwRhJ4ZddbRa
glDdc9MVxDkU7Ke/H7k7gicT5xg86oMmPog3G7DxHDI0xqZdTZb2KpTb+3AX5CO7
2py1+26AXBIQas7vBGlUBMikcHEa1RrDdSoKztonrQdLXtvXVKC+mXjrDETlP/YH
rS7ORTG0Vsl68AuVKg/omGRbYk9gnCUMbOz0Koi8kO44jwTI+DdXbfDJSUZ2+Rif
B6NlHqf3x2iDcL7RfAQLwQfWZq67zHE4sR/BZLZkxtK+hvlEbDC5aasBN1xZbi7m
qpgWsMWaWAMbT+WMJ+tLho+/eWtQLGFbwBBk8s9x2uJp65tmiEDvrHwylVaMQXfH
FBimkfYRrh9nMA+18FfhjxGplwfz+7878kXNcmBhDSpRfGDEb4G8ngoVivAaNdKN
F7BJpHU9aSVqqv3nhpGeX8+gpmfq8DyirodKXSWaQ3wWieYiwcj7UElf/pQt7Ptp
H2NDAzf62Se+N2u5DrrAkqera+13filzjupzJgKx7ETtnPVfCpUoL8vgOuSOP1q9
lyisj2OYpwxwN6XqryO5xVoVWBGR/RjebGnqxiYfQ6TjvYYqZaQH4iYLLdHNuf6E
uRB9UdBYeC6twJ0IPWYoK+E8+5QpadMx/CIlLdHNdrSkWoVDMJyRwFIZjCJcyFpE
qaO05TTQ19fd8LRsARLQ3yV1/CzvofpVot9oBU/qf35+kjIpgbadS/F6Iysp5bCv
wgaMuTV2tYclNP8Q/dajS6BqmSlWY1Gbo4jv47LiHEh5rvl0v64EK6+fYyCdC/Jz
nQ+NQSTespqzU/mD4buoOjkh8UZLSbCgr6DgY1mcKCNSnsxjvnGSGVxPjtKrKW9s
LVAZ30pRTSzdvF4h3xQmVvZN0haSOMlUFFQqrb/lsSJ9iIuUGnZNeP8HDnaoGx3/
opN7mN9SBZDoBcbXGxDyoT8CvxWMtcfJbR4J1zi4O79oIp0nt14pz/3pueR8u5wu
QNCfSishmct312Dmf9AqyJU561AOAOSBJ63Vzd3URTwih7GCUgFRHp9xJ3nQeGHZ
V42XMG4BSz0wVx6sz95X6gskuqWm4W/w4t8sbld+PCUciAwpV5g2PnOTbi+3PYuR
mbt5UuKcu9Rr7n6CHKSClOPJRngDVFpzEIA0UyKQKGIHrA4TiLVVVk1qOHjedbz6
YbNhWSfz6tuay9xDRoqEfFPqheQrZiTkx8vtNGGT7BN6yQLG2tor4kERCJ2oAyl4
WG3YrWX0Y5Z1zEOo8WiCV/PtwCKorj6wTxDKLlrYl4+JgLaWFZHkPcJVUJ36C1NF
2KHJuCvTv4ScbdpB/nan7duNEsWaToKcUMun5CluGrmW8GGkqXGWpmH3fZ51rwhD
ZVZ/77fRiTge2SS9YPSUAeNwoxhKNZOhIqaFQEX14tMITSf5SvY+xzB9MTlMYCg1
sf+HmGkhOnKpbq5NfS/lqo68CtJKUevNtxfxtMaQgEGwhdIzWepteM7yFK2HqZkv
po/ceLUDb2uNct0n4EmL/1MeK7Q1ipn8//i9Z8DJpHRahFAoDsdPz6tTYWueoa1x
QBNnAPYCGVKrRMRwRnZKIMqZ5JDjnkcRduItP1EOMglZBjNYJGvj1Mux4r/YoYj7
GwuDBLzF3pNBS2l0l4MpMe4RYhwNFmx/OajF6KbLVcH3F6iTUAGj/fLGdxPBj1q/
G0GA9A/YsaA9q3wSRsOzX1lcv4Glf99wF96fhxoPIFXfuEMrgqxAKArnu7zNjwNE
UZNfgXAy8i/m6fwH5iHIat+geuNPajwFQZ1QTmVL8AGm9H6HYpdnH4XWuBDL7rvP
nLfVQY9jPXP5pbLrqQLave5f5VZkGmznZbqbh3t/qrRummi2uxEvVpkV1fOZ6PtH
kz+6OtLKXWJmd7R9dIrrh+WNgkrPykyu5QtTZQ8jXXuAooJjxA+ic6CnuXnxLAlN
EQcuclaqO4eYU53Zic8kfpHmcmc8T9tqKe1EWg70Bu4tzLSJcopzOHc0TL0mhxxZ
C4xKqbG2rTmZUkYr0EVaKH+TfwUs+V79Pgb+UC+MR8VZEQCZnEbeRR5gTVK4KrvO
+jvdEIDrI6QCq05nuiI5xOm/AVbvjDcbeVG6h9QVVBFNMLhyiiRa4L8T6GNqUZXG
0ukVVqTj2Bgl/PmS9zQO5bWqsjSf+QLCPLv+ahv7xbwIRQp2/kjHaF11QLNquNG1
yLmbOkDSHR+VCZLzLeTuO2XNAZcGUOyFvixHobpD2wsjU+TQxij5Rti0DEaqq199
RB5AjGbAozbFTkqSV1vHFifJeceysv9wJjbG2PIS1OZkV3tiz0MPE0mx0CLryvYN
o0jvPKYxV0/U9iS21coIMxdzZZ3d4lv7ARb614u0cx3OOycZAB/U02cHkyG1/Mso
0Gr9qnBO5TzG/LDc54OG05Zi4c3aipZXXv8rg/NLoax+HJkz/t5r2hyGtuIUBbks
hwdTl5qjM5Y/s2JSZQwPQ3oci4bWvx5J0kdx2soXTLDc6mqSMGZJhh8XOjeHIErg
HI/+w659Lrz6UnWMJf+8iea9DeAZBWyZU9XtNhG9NuEjifvrRsJf2UOUiMHyYJkN
uisMbVCqhRqfW91EDkXfJYxy1vfsm5p1BzD7Q8rZUdmZz91oNl6tVbca7lzHyyB+
ZZUVGX01Rfy/D3Gtk/HQqmo7QcTwRVLoNoKGFtIL4a7bwBhiYfJZeAMGruoFVy1I
tfJtLQ6rsqWN+BbTuXb/LuNQhpViOnVREl3Ej5vvHkUHzzzyUT+K9L9rchFDJNlO
EZwCKRvwGbVe0bgM5iiTFiPYrPauRH1r55bDCZQS5T635Ptf5K41oNT7NzpYJtZr
PRdLudMN+7GObAQ6zUCjUpCKo3BRBMR9qCtTO+aizez7LBnDock/vkEAhn27xeJG
8RdYKsYOksok5BhzK8X+QYWlxTgZ250B1TbFlj0QYsHHwWMwNWXIHnBA5xMdorpJ
vdhh9aOKWWtXbBr+Ui3QBzUGIB5Bb1eF9yl9vxzzhAcJ3n8N40hXlK6aLLb1B7xd
EXvCv7Tlu02LnGEetew63LuzvcwdKfTtPXXg6sNgGX3pRv2JKQgLlmY2cUfWf32E
oMrBep4mL+83UI7lB/HiFXaOmjuX8CFYRnpwEPosAPKKKDp8FE3Zr2kMUtwDWn0V
OnswfUkuLj2FPQ/NpyuQtG+lcOetdJNHMQrtArop/WQqfkx/LbpojANiX+GpEhWz
xhrBaz3ExSffqyiO7JMpVZ9jg+/Emiag4g4tmrZPzI7lqTrbmAEPHf6+nWCNeTWb
X338K29eI82evs1KXINJRFsOwmnBMitXUh20Kn7++qAwFCt9K0SV7yADG9sS7ty3
UtOUdupzRor+mJZoM4O9e6zr8r1WBUYD3OyxD/PhUhRdlXjeg/Qfl6E5ubRGtQPF
eT9hGeXMHAbnuEO5dA09ZXvI34GTtkYMK8vWrdTGceOR3+qRrKPTn0u1ASPsT/ou
80GvTCOFoNbu2+TFkZkqeDUGXCYxKd3VQQnXU41d3u7/KvxROfPWDMCcKxsDZkXD
8aaiKdlobBAgm2Pq5KNA/7aqQ5D42oC7usd34itb8R5hmNkZzVn1m2GIRLvpRkyL
abnK6sCPlC/MAw5gIIW7h6Va1vD3m2CYm6+6BUC5zKeqALjYbWzYU9IdeCU5LQSb
UXteihUD7yHT/3veTvp79Xsr0HX3OBs9+t97BpQbW86JFmjhXN7jFuw1EGnWQgqT
2+fv0Bjp6EkfvjrVy9IhNYaSKaIfyPlR8+/hpE8CS/I+LGXD2TMFkvXWGWLAY4eV
nHHrrCWVrJXbXaHLLhDLYljIK4RXDVmfDABcImqij6ZCprgoTnjFm6aMhACWQtiK
f0b+ISx3Slwfdz1oPsO32dozX/m7T2aSAiZ11uHjoR1nGvwg3KB4zAUuKr5gLCtt
eTxnx19iBF16Yulf+EKi601AVtl9fwjreSMeSeNKtxrVF41t6G1Y+N7YuKAdJb9y
ycZWNqTzZHDsTnAHAEE7lIgOtN1TFzqEcFtXEmx43sVXawbe0muNdJMIIqaMydyA
WdL0+nW9++si2YPj9ZwQVqGJfY+7zv5rwF8NqbfLgbJzbZ6qKLyomRlm1dP6nf5h
IdOgHy+T6EHsjSSUO3xyDhWqgDUBDlLK58tz0YL2O/zQHa0TheqRrUXn/bJajyz7
VtOVP+NQgES7JcRrgrC0Utmas/9gF9omsd9ux4Zz0Za0LTbIekMu1UOBWGUmxXsM
VqPf3IEPgwpdgI2QXQABtrhBgNR8Fq8qQArmhDtLuQOlHpTnEwtOKzr6Wg/lKX+p
pu1I9SLj6P2RihN7fn67p9G4AiDCP4i6DOLvdku1xx9o40gElROskgDBQsLUEINE
wQhdwqA8zjnbe7Sp2qwE/0Emc8/ze6LlZvMZNESEVkt/MJ98vY2MzEovQgsU12Jc
45jLC2gxzbtx/lQDvY1jl4nXYOqqXDSU78pnb2Q/PMKjeRZstbTcx1XqruZe0E8m
WETk8Gwqg/CcJg1QNLezADvfsFgd8XMRwhOXWMd9rtvjAaskilG89qx9tvMh6XXG
UqWjUSkh/W9jiPLGHZ15MjT6yKUTWLX/gF24bn2FSgA03Dfwa9ADA4EYfuSEl0EW
jk1ZqTHUpMbfr8qloGvEYhc/gtZGcijvZQseriwqhJPy/2CDC6rcQ72EbVyB9QZT
7EgRpe+qHcymU/wkjzVYO/+pM4wRkKqFrVyhwj4tXt8QfVUgBCLKU2qHZ/qdj047
JxMOWWUllFX0YJKLzxHBxXf5PiYCokcPeLapYcOYjaG8Y//q4AbqjLzsKHd+tfzK
HQIaeof/o60DC2Pq6m98wbdhpxbwuaqShrulAuwcxjARVHv5kOTTYAn1Dexc7e98
/ZRO5gIG2+duHyQFT9f7YI9nYk1Vk7FKoHVvAZ1jczFrgj4pJuJgkx1GjJbDt5Q/
W8DmFC29zxn0K+AfI2wUeD2KMEbwrnLmjANDXICAsVOcos52ykvg9C6bhTD4UtLv
M17u6rimS51W9h/8iX8u7MJBlpZAbC2NLgxIkCyzDSTtbwqSLUhGjwReUS3+ri+3
v738vHLZg2nj98QDAZ+zhU/4wzthRzPRgSuSSADshYJKSoRB4DAdQbD0gRkgShVT
l2kYkfk5zIdhmpZ91eLDr2AMyHczW0UVmiIFqupqwFRe+kWHJo5lqn0Z53CwIj87
IciJZRWCEPn9v3rLOchaII/nicHK5Nbbb3HsiFRBBEGRD4WCxdHg45LQATY5jODw
aUltE7w39fjUa28JDtCrKcK/R8hw2M1XD54BO7ukU1ySyu1WnycmyXRSdT9rUMdv
C1Wlq7s0xn8DDdQ7MIPUhXiMQZm5OuTcVJ76CYqhVPkHT2kZthAJm2W4+9jeU8iV
opqcVLmzG1MLiMon3V9bLLE/mnBCB1uq3kpNVKFnh1Om1mPyTYOQfoU8k3JKujgE
XGzR7tzQqn4zPeHD03HN0PBVy7RxX0y9HO2GbNstxvSmzkcZoHIQ3Wwb/1cgOSnG
VVyEW0B5d6QT2p/jmIUXBzK4vkOL3Tqpmb+SUPwwym6taIpKpolM7YVpWGj5Q1il
nJMCm4laHEs6f2VgjiGbjc47s0uLEnEhVyVRCycdLgZbofs7owakWefslbn/a9PW
U3yNPMaW1oZT/q0yZNgvHJ4J0u3w+bfUTuRSRy6fw/IG8ZUJ4wKMtEHrLIvyZmo0
gsSF6thUEmh7LARYpeaICcVHCTzXEKXzbxLXWP08Tbelh09HrUfOaTo1s7rDDBaZ
gEBgPKTcWq8exYqglmnFVaoAhrdBrZrO83fQDBRwSRMnkDhwXmfc85TMw4tS26We
lyaalm/ErnRLli5JlkrzE2mDSTdpqphef5M2BFqnR6Vv168/Q+IWL4TVacAm1lpF
LCPKvJxeUnqiSWnM5Rup7hs2ajIUh0CdjNp2DtW4oX2SZ3lKHapIJNJV3yXhl6Dt
E+82k/V4xC1gehmptxh4uYsfvXEr+4oc6A6KB5S46unXha1/aGui6dlCeh3pVJiW
M5Gf/arSo1egdx4p/OqzpJGevYnD29CFn127emFRCthdWAcscqcsOYyStzeTfD3b
y8tkquBrPRDNwU/Flq49DjHiv8iOaEcHlz4MSceBnA745WmhfRFao4kZP6dBx1Q3
+U5hX5kA3FycueqBehvRUJsGgOYoaXVjQKa3TR1+IFOgKNjzFFFr2pRei0KmVRFx
JZnShckHhy6IAm9SjKRJtH6B3Yl7Bcdnq/Kj3pH/zgKNApXYY70g6nsGmZPkrGhs
IbkteGcjGYx8pgMlPuitZFdhuNgly6oIWpjtJ6+ge/WnyVhfqtND9MfPFtm5nG8L
VbaV2dOyDdai3q7tIa7ohRDZWiCoHUxlRbE+eB+thvNRj5sbm8L7GZniFBiCKX3W
jhgH64kQOze+aJFcApVqgJF8nv0F/ucsBQe0tWwOLwHh3O2CJRD3gMdMj3Ll31qR
uFDgcwly5VAj8GSaAt4Lz6GaUmPMDj3JAoZ2BRsYU6PBjAjq5SG66WxuYghOyz7V
Q/t5WA8IWTa0VkIDXj1Zl9wRsR3ltrgaCilUMLjhOCsKdtg0EIklaGJOVUlkcIl3
Pgdhk9133WlnfqNU+N5nc4OzLpvbI9cF501J+h07Gt8sDV2W9b5Gb7JwvFK751J5
0qZKcusmBN8emq7FuJqAJHYugIYxQUx/c9zHKoQ76+aFHs8uK5csFK0SoGgkCagc
ig2N6HUbWa4T9dZxmjvj+KCb3pqwbskQbMkA3cONFPSprw1GG1kvIJ0JJVsM/XA3
Cd5yOxCdJku21cQpc8kWr1JrWUNtblY8dRTPgurzG0gyjPLoPxMhgGrEZaL9A63u
O0fbnzHyKDabLW5Fw1X8uDVgisVtlrh0/nMdZ3ZBUL5/LcQPJZOfbmedWlRviIbX
jZl3VGBN2zbHWOUTr9vy0y4yC+RyxwIWDmURkCEQV8XZKcWyl9gObHgbnHQgAikB
cB3uvyVWCxOAAhKO3M61e2/0drZAV7IlIeB72PcttLWOSvuIUROsSbpXD2m12v/S
iHx9kd2AUEXPEerCV8/FHxdXiNp9CiPRjfiQnC2UXP4SYlpQZ2g5odraCyzMTqfp
afSHo7FjOrEUaKyRTaAh8/0/i+d0PkjdFe4nyfYTHVlq7DFzWqehirewKmxNYeDC
ylT5/lLET5ohTYjS0EUe9rr1v2p+BgNjSBp5wgtL3l98G/hq2gKGnhYGRo+0gl0v
0nL/RuFnzH5AHKX9ldnunfsyxnAWH9FItTKNHkx+VOPiWehVXfDUe4J0vC+7Y2ld
k0ETnzzESSBoB67bfeDZbzRtgSfLhu32cKXe12QKapzbrdJkmh0pXCIzjCSXbZ6t
8Qt/sFQW5ACjBy88YkDvIDQLgkJjPQur34AWNV7FN36ghcK2S5atSFtM7M0x31Ea
hZQYgk+SUAmrOFIZclC+vsrtTUf+oKjl/ewCzIDMGDsW2Cqi9Sq/kpOxbxrVWqZ7
OsgAN6Vj+4QTUaohJ3WussEITpC3y01FNYQIRRY605FTxRMInSmTxkFBXWX+FEt2
JC5RLTPVMxFq7kDfBTLOj5NMYnOXqlY2L2vjpqS4mp+geyE06ziZpQPin++7u+j1
34tndZfn3QgI114t/WbpbwiPQXFctf0pc2mo98YUKcblrYjX7H7NhAFXNAE6Cc++
8jYiqUwjVo6Hn53s7UH/zGQRon7BBILcqJ0mtw6gBauYcP1Z4eixO5M1gt9jOlh1
Do5I8637gBBCqtkjGeBoxlqjyny6STtBo6nIP68tOM2xZ6NeOETKw/i22oqAbv6C
n56rypmy7r0JmgFfSY7Z9ktMwAzJskfN3xT1uO1iQVdA5GfPBDH91tWH5Aw+RtWo
h77pWEKeQivyyymq0BdwmejdqtraKc8okRPY4uKr2WJTHgiXESfvFqup6mx5DDeV
PJnrRQ2E+xDyPAp+tJcD8eLroVhWYNEojiCMoQU66zs/HMIjz9LIyky9e1/lyTHL
0KfUK8EZdKwGQ5Bb25uBWHrPkc7P8FByGZTwLOjAvz5VoBwLQNugoUSyDrKcf1Rx
tvCe6+8YQqym3yZbHxI2bpkO0RvQHmlvfhr5j1U6tTk4kxhp1QZyspsQaD/xZXK6
4H6RhtCKDP7fPZpoxYSaD+M4CyKXRUF4f7NVz6cQnlLpm1tWd9fV28wKhlkGlr3Y
N2DVVZ5i0HCdFyzOCBWNS22Wf20SFn9g6wYo454MuJ78BRmU9mR95FtX1CDoPbHr
VFO4qHmGEKnsI5tC/LbYDwiZs4Xtt2whpbNgkdu0SXOGZUz4/7/IY6lZJ3p0T8/k
UoRdFaCKmMEezdlqWsY3FwDZaFcjeP3xBT6w6dsnF3UDMIb3fBsGT1XC6GXhAB/i
WzDZye+E364FV7FfF4EwKdqQr21AK+Cr3MklbLX+Ee/M0whICLPKSOhWNQ1NakVb
Y3r+abx6Mfwzqo+KhW/8aP7nF9TQg2uVPNvTi9ZmgKb5vnirsgAutYr/2MyvLHx0
hc4qW2qWGoTUBbrenhVoJXwxsYsARYk9O6JQFp2zllMysRwd2v5UCSpRCsjVq+06
p9Ozdhqm7txK0oUFVLtN6aQYOz+wjNqsY9NiuLrvrHBxb28uvR81ga9LOV2rkpfY
vYOOsshmxUKDjlbbsmSpYNxFYSM4ietYD9mOqlKHaM1XWdDThdztUVjxzPqPEyJM
Zqo5RnRJ6tfqedVAUZDbJ4nF33F0Qjon125Ix+ZDMKjnl1YT44f9H5x2dTrokKEt
QiAjNjwD8vJmyo91ikrF3hutMv2MsJcHk9T0wMBiNsi2k97AURiIelba+qrS5H0A
57LmF/ASWW2j01qCoaPJeQsMFCZ3Lf0/dN4tRlsTwQAKnseI2eyp6jIamvCgr3JG
Q5anyjRW4eQJvRCDzxoISwjxEa1euteW0CLTAn7uZcoBPhdEZScWgJFwCEUfs8pm
zEFqRy+bRL1WLTnKa2Khw8nHgsh6/UJgeWdQ7CUGp6p5+Ob3vNs2JVcFAWblaT7Z
g/87Hk1+zItJdF+Gu9S4M+vB2EovPkVsEw8JyWES7aAxa04t3ac3TxZSMT1nMTq+
ftAbyipml644L+IsGu4kLNp0/52P8RzVSDHCZVNYIIBCV4z9E5teHmWRfaLjhQWG
04rRIyj7MLFHMlyC9ghPWgImI+0Z3hrQmvtdvfRgy94syYlv/UZuu3YrGvnnF0PA
KI/C+1I9lHQsJamMXCJ9NfkeCpVs5iK0Snxg3/JsZoTQ4KhF+1tSrjIXHWw4NUjc
uDgVNiDLkty9jYBhTvS7AEaG49IgqO/dVGupneiI8iKuTZwOUNR+3/kiNefgvIyk
jl6n0wPOqvoslLZOmjn5yuT5Vtnph2YFkPhx2L8LXfd3SL3I3jXBN33W5R8kJ0Xc
e6VIOjgI7hwhnbANEYuu9X7ze3lHPO4+gjYYvOIvw2H8Ksgzb+q8W9PT/Y5CbvhW
D9QFysA/m/mKb3O521yjQ82oJVsVDOixe5XWWodBD2eY5W6FLfwP/TajpUgJDvEb
Ut86ca3mcaKhs3EpSihRoKgY9xUDUGvOq7aHAF2J1XX0Mzg606q0lM6Dv+8ZJNHL
WDLkUESNc48+VoIpNIxjE3eDXikRBoh5Dq6v+l0kjhaFv1TvmL5skPOAz/4X+H33
JlQesVBnegV54DpMn6KxBN7agQD8PhiqAICPmpLUmJQuIGiMrPr6Mi25bnVPiae9
LQ1RZ8noSy+vgGWKKHVmM6wde3yzMqQAVm2UQHIZkywheNNNzI3weyb80GQe11rc
7m3qVK1//T6WJY6vLnWk6WpWXglK1nD9U2WBXpN18qjA47i40IQ4XLK+iPkrHG6p
e5SZFROCvKef+IDGXg/4cZWPIYjtMtembL9MCEC2+fPvghHsqhBwfwEDooMVcAQV
+XIkqhgI3Y2YJs5z2cM26Pjl/Skwpm+DSBwAKRBqwfmXOGOP6YRpzHvan/qf25kg
GEBCKzucl6/vn4+d42daGvrXkot3G68bj5j3zfMnIfJAIdm1RSFx3iNHkPKQ57d0
OrEQYCebiF5OSS3kJ+9xuPn8E8FLhdFeZ+LimHY5wYsIgfd/FgLAwOxW91xzq40J
h0X4I4BK9mraAVokDZo9J3rrSAhUpji37lvHIHjgfic8ybMLideni8jj28VgzuIF
QtzjBdfQIfWku7k0lxVYKeYwVDE8aI6AX+JZTiG41HOd2woL+qCdtmY5Ol9a/CTH
hfHW5lRTOkjzGAHFrv7Ho/3ymg2MysSOGgxZO/2JOdWHNtzoyfumMepWXiHZc1iN
sMjVEOexZUCkJNnaZmRLeZG15VfPTYgigJZ4EiRcAUKtrSAqS6hqbEYh59PbTJSW
yLmrHjuhTmO14Fsj88oBevXa5ylgdX6pY9ZMSUP6MfXCfu/Tl7VEdDJpHGfqMvnz
/I9PoL6rigYs8Y3I4/G54tKnTkyK7Jt4/zmtWSXQv8rViBbL2W/d+/sfTYdqzJYo
iGJGR9p+SdZCtjd72XWAdcX0emP0BLnZlfpxDcRRqbxF+9xsoW5wHGuWVRM/F6yi
8zH3IIYT8RuR/hbdK+fyFnOnF5jZdJ/izrn1IiB/48+sx1rWZYd4HyTr+Vy81Ymw
Qy5VAKKc8iGJVMr8ZwiyZ2CCOaxIze52tVHY1wuawVjTtS0CMFj/bbYhdrFQ3qzC
uL2OMOrkaA3yvIy/VMzROQUOttQgxOicTc9jjVVoWSd18CTM0KEYeNyqZUySXBea
46CyjP6w0FIn2+zuSVq0u4SwKonl3p5EWuhzUiuBMwSpFC9xunAL6bymgRDzWI8v
wrvWglcsHjGHq7k4gi1J4Oe1ZUw3rLP/JBQ0t2knNr+XWnfehTbYVoGNNo+lGoiY
WnVsJc7Uh2vG5gFeuqMe81SfOHf9jB8E4TRV78xezf4m5/yVtTfzdAtT9KRP0rsc
G7ZJchg1KAkS/YZK0Bc14CeC+7dRGRRxcSt80pAcn9sgvyv26N4FfaAV2Lc7XxXA
LIH2l01ky2dOSA7nXUfBENb1Y0CN3yDVTN0VgWaxDbxDtrzakCTWMbye8PtBAAzg
+twfx/ffO1Qk6ouIOmJTLVrc3HcW9n3obRvpBUSP0eaaOUxlQJnLPBliILqANJpD
kZPyYXEK5X4IfrNtXQAzI33V6oh6ppQnd9Ah+2NWsUcAte3KH13TBcYscDm8qYqy
br9GFY88X+CoFC36ljw8MODwutCkRpDNactqgaFba+4flKSEGKvcgwfaBQ4hfYn4
/hNCGZoFiPFhDCWgUTD5oMxKy/dU7r85zOOg37ZN2oudXxtZRW/upTmev0g55wQb
+tisUSFBVitYfIXkd8hSm6uJy+HsmHPY92PGpWqRoj1jZf6x2ZuisuTSw/+7nBag
whAZnG49susTpMgEWavdg/roleIL8jqjcY39TC3HW9XGK9qnfYKo8G/Asj6/c079
WClY4tEG5oygljKTqD0O9erOq5YQEfFsEJ2SIitDFAOY1tGos4S1Y6C10Dqot9Fu
78wUdUQPkuB9FgfmUtfMiCMgMX0P0ItCJLeKUF8oh3QRSgvl6kLWqChVlHLlNBgI
LTVcqqqDAQVb+f2jzjMcLM6PHIl1yVH6H/igI4o1GkFeFhFKe5H3gUrGbcj31X3K
P3DmsX/iYq69DTmFiWPZwoo2QpCOxyFjsEiLHgvO1lOcXooPrMSTKoLCFAe3upQs
P4UQJzXQDd3RKcIjdEyYUr84qiX1P2oFhfBRB3AekeOw2H1I85vV6Rms8uBeMiTU
bPcpbM9qaVMDgznZmNb84dG3vshTichoRb08AtCDGP54g4I4BWICCXNevUBlM0lb
g+rXEIpM0LXp45+H942kGwPdxTVdOb0yK7Kc3uzm1YbUioEOPxU6dwHr/x9dbHTt
qe4MG+8xq+jz1d+3/fQkmyC+6TCymhuyAW6Zk9+ZdyFhRXw9KMQVRSiR9Qjf5Ykp
jSBI67ggghbyRLktX6tbhSTbwdApfZekTTqIG+Nt6F1H99UlEehCaJOQAyJb0HKt
m+6xno8+tBWFiQqg5fc00xaYc50ylZEY9z7TfdVvF/xM3RuvT5Ei1cTpoJrYfXm3
azPmSAu/XvjWPjB5PJUvj3z6F/g/gCxS5JwfQvSazQrXBdiDRRaeeIoa5Ym1F67e
VXowT9gscnNZj9r3jGko6mNysc6p0Ofb+8WMZDNImmU/ZaGgOqb4Z1ap4kZf4zE6
V7hz30hZ1wTck6KjOzWMZ2+qriUiS1fagG/QJxYJQUC7AVuzAYT67az07xJt9auY
XGcoI7SNH5/YopgrlSa8FcgSRridm3VPAW5YJD2W5JZdWHgiXl9PAO8pMwB7UBgJ
xp2bzBm4chyStSsohVf7oTdZmeXaTfWHBmhEaBihY30OQm0v3n221z60xa03ud6Q
VcemcYEOGkzGsJ7hZJiZF2xhn3XFfHC6MUkzNblVgsayE8YchDsSuPu6iA13tP6w
7Qwoz52cMYUQN1d07nY9uy27nVKFRkf5p9KM+KU8Mp46ku1RgVq96p5X5UYJaH8f
zDGBi5KRnwjidHulps2NaB1DNyMtYTlKx+Y3zEwbzWrxBbHNlqg+/lTiD0nb3OMO
WoTW9g07BfFxuc/MF/YTKx6rFoV9U9BKVAEXYdA0J1lnAtufaVPpwihq8F3s7d9v
jdXKjcNtgeUsofj62RFgY6VNDio/Br8szqwHxT2ichl3I0kTu19g6P9Hfj54sK1S
uJr9ciR9kI4kSzK6K6vviENgiI1BFpE8i7dfl0kIZHYc75p5NDQ2JRQNoYWR8iU2
JuXKPnda4ooyMOp2cmaBJ/uxoJnFN6lbKNyYccw8b7PNUyufDKelZ2mZG8PStA7z
PCGf01RPTqqj2FSn0OUNrc4KBOUvOXM1WBg/8Q0BQ1PbdriIp0J+K/az2fM04EGQ
IokyAF0yvYdDK2HStv+fq66GmlEbbqWFJrjqKD7wpQikqGv0S+Ow2McE6V2STzeE
ptOl8iGWTMG91vNkPMA39xHmccALtlZvNuRJIPHtd0sv83dEwO74evPZ8StyISmf
SfjdrWKnphINhsfj2d80wWAP+yqBa9nQ1zYZ7OrLeC9IMqriMj6Msp1vt+9RYRgW
Sbc+wkgpHUBnpAb+v+2paLnswMzTyxmLGJm1uYMmgCV+4kh1gMn/AqGC4CVVqdPy
TLpD47Q9RruMbuS3MBUxmw+ft+WZKgWrKIwKhAnLw/wPYD5J2Ut1qHjWr4DOS5cq
nCo9mfq5jgB+rkn12wRmLQcjO/rLenp9/wBAyEtQcgOdlbIkgBezPAXzb4JMyqFF
JJc0TFZsg1fCX2LBoGsGiZVcNyQIqXqJIbHDFZgtw/oyoWSj1Z8r8YdBSLx8/sf9
zvNi7sNHxEC9hENDMB9ReXfXDic7qQCVsJLLUdCqaALjnGgfjwWf5VQ90JOMxn9u
SyyYZCXHshFYDNYUwgihIt9Mx7CG5PLiHL8JZVCivLBB3Ktnu7ypvoi4bY6m3cxS
0A5g4CFim6BI4zZcgRnWCFec/DycP4a62xHDMc9YTnfE48jiQNn67YbXtt0tP/FU
2aIeVKuIc0EHd/imJ0iRca8oJ6p81Tv+1p4yYicAuWPogdBvaGCLXXYYWdD/APWL
vBa7SfprumyFVqemtTPP5L3xT4ATHEknxgtHXAF8xpv/c2P0VSoLrubVcRu3JhNK
bwqpo5+c/7oHfTu85XV0eH2vD8B62AeaB6FKjrr8OcqCcA1VtMif/c4zPZyDTnxp
uKaGCp0u5Tlv13E8FBxzJz7OJfmgZIh8i5/Z+p0HZVkCeS7e1gpPtTL72t+9Sb4H
2po+PhRdhgiqL1Aur+8QxkkZ8PYXF1DoDWB+bXRFQvtBA86SEJvjW3bEWhoGPBU6
/mq2Ao4J66d6KcgpXl0aZqWeeBMA1h9dZ9v9vc6OzvCwKbkWrqAHcJ/nkDpPoFKU
ldRzJxGlZ9IZzGhVgirFIo1ViUT9E7JBQwYrCGYV5n9Mqa/uL5DUJ1eDuPxGNone
dEDv75NUsgCwgnFzJ+6k8x5vQ8ptnNthBEKvFb9aj41L+hbuJgSegs98B3b/muFr
Zb9STZgE14RIC/rk6YYgEvccCD4h3+9RaJQuZjdeJWZcY5ZMJzF1PX6oQMrIa1zg
Vi2EVbAr9/ShBFwsuyEBcFhxvPOGF62N09iFAJFAToNBhG0F9N14RrtEhzUIy2PE
xNyeofUpUQgylETX2e21Dc7bTVUbNIQS9iaZ/c+c1Hd/r847Q5ilV40+qlBRyXVU
Jy5ns4outQ+b4I6URmGrRu4BcicjVHofEHCdI91woeF+6brAmVfKFUMu+dY04fmg
IyhL+oMiRN9cB/cb6FzJ5D/W6JP5AhK7TXuoBy3NTF5qWUvU8iekWxv/LbbG1edt
cyDsitNMYCMVG3n2CppaTNBp0N6T4vjErehGy1qKqbj0EYW/yg9f0IdAp8zHxCAa
YrF3hr75vZUgjwvJs8Z9c7mEBKu9oieYd9ufvYjeyiY9BmG+bEJWFck8S83gOsZr
AnrHoDH+vZ1A5c+txGbpNVEXzP++3yGSaHLN6mAeNu+sB9AT8E0KeVGWOr+OmlFj
dbuJwyE0Kal5YCdAjrya0AQwLXWo5NUxBi5QgfCprnCos3XmhLD7TZXTucmNIEda
EeB5Me+EjZ5E0Id2pMvPUT83uDWRRJzmPeQGH2+1JzGjhOpd93xuuinaOW2ChYF2
kqs0SMABVkzxQUNQpcVYHN99sOinz2jLwpGkHmXIYVvRbpsFYSy718+oOx4sAJu3
37+H9CL9j/dAOQJGiXQRfR77sNk5VqiPsDJs6QFvm04RqJ86qlmw/ZCLoaOvUrFk
vY9VRNUi9KqCgyTmNM4o5QWlH9tB3XAtmUpdPk3Mn3YJ1oNDpRvx2H8bDpv9PTW4
5mSGnpWkEiNVDMFCkPEpZK/UCR1v9KGo8KC90MRjbsfO+5ml5lzYj8k8GI0YLPGh
IRppN2TzVZef/NljWLvjQgQDo2HN0H40B6Z3JWvQSEnYD7aTlprcaOKqjbeE5feP
MgdeqruZYnSeFd3VeJ+X4wU19YFW3e8oxs7gkFr4zTjO3gWPEgmkZYkID9bmh+le
M4bAXwuvVZAs5zb7CpOBs8HqBXKM0dc1bBHbr7yN2KXUC2A9uPFvHnDztqbA7mIR
0BOQYM6rz47lE/Y+fBXsegTd39mOffXvgr4Rtpsne95yAbHEbm+52XFo/PXcSQwG
PAykT40Npg2wZubHjgdeLDWedoKneER1O1p4AGzybQQNHM2nxRRAaR6pyVkz6hKQ
yEclkdihLUXZVA2ycOpRjUZRPaJYbS8zb4MQ+zbSd5QzwON7mO8r7q70aVnrwtFT
U8Qy8tva9zp5QrMmgs8NfAzARk/BCkTUO+Atfdw5xiwv/8TvRPw6v1IvQRXbrkzV
/ZyGKoAMUlGOnzRXvw/BNAdfjrSH6ydXAcXKuzX9zws5XzIv7qvBaeCN1EzNUR5d
6/dg+uYga1hT/yrZiAvh6TVY0YrEJWnVFBLZmrOJ1kwbUYE9gEYTDCn2WiTYWKhf
FLd5bkkICDB5YTt78a/SEV/WZA/fr+aoYmQ8F5wtmm1R0Y+ZHG8+SL0lIxDwiCIA
g8ijeXGlkyR+VjbbWPEaiK6IiCNyeSCGZtDUaghao3qxfiwGoiJH/zNiJJaBy9fT
S6poEbg1Yzeo+UJ8F+fifc7pgN2H0FGgPqMqdycfd0aPuml3pr+PfWdLFNpFp7hF
LmUHOTZVx8hZ/lN4GvPv0Ez47rdIau85NztBRchDABfPpOio/OjKs98T8T6Uk/RT
+n+v+Zpy26pO8C/kFpyajDMeS+YIbLd8k3CBuzA9zdGqPl1ZD/KwbanmpVvonTJD
J2QJ2J6fzXeHcv05Hu1lynaLlnBhdmH9xFesDrnvfzOPZC+CWUwlMp9n2gzipRpB
TjiKrhx3SjP7TAQYAkp82kQCuURe0lMsYKweMsLjj50SdZrO34kDTRxYN+5TKQye
MacDq/6AaeInbBrQPyCt4TD20vmAn9VQg11RXcK3cSNCKNKD341+Tkejykofp/FD
1DCDL3af5UPu0fkNy/X6g1Xv2F3gUl0SEQ99BUET25bYHmaj/Qwa3F/goXPxOS09
qsWGtBkB4q7EcN/a8axtj0apzt9fGd8mQ3l/1DRfavgq/ax34dyoE6ZYNo1JRVbD
RODsam+y39kSWAV+wV7gQ8VL7HIGCs/Z7KKqOv4DtA5/CaG7YjIyEfoiXH2ebjnm
eqV2PjL3BlsFrNUtlH341wYTSE9b5MhouPR017V4koc4atTkISeCCtJGj8IQqttC
+da9kspJtgjIiSvuht3OiZ4qiHw4YWLNH9dc1qo0Y5UyCDKUQeNfqsSk5vDsuXpj
ntbyaArlke2vmwAQwRvUBkl6GrhDiVrXccyUR/OfHDR+KleKo4gSMQt3InLsCrlt
xT8Y2dbhowXYTeKdX/ZIYw29bJG+IsygXoYQGC78vnzEqFQM756igIN/JDCDGLlt
qTiFa3ZQTkf5ujh7ouXZpaU2JP8+TGQINsAiOqOR1p1TamxlXNFPtMYIzGfSg6Dy
LPxeiqWUN036ANWg7GCGb1+UyVK8/5JqlO8j3XKTKo+89yBxw63L6Yp1P7vdItc8
w6KvUqy9aqVGt2T7vMcXgG2AiXuyi8QpftK1hD4pA661HW3JJcdcHOwi+Cuwxtf7
9+eqWCEcSC2aOGkyETgcMnGgiALDZIg4gM7wRKs3DDP0vSS1wCvDs2ZQZRLnwvSq
uHUObdMYMH+EswmKUNbUmm8gDzmmVE/TkNY+MXg1ubrHHHvyYtOjgyruU7DhGIfS
L/0lBwQgLnLv71d/k4XnGpuhfCFG8RYbDsipCVf+f4w590S7nfr/0KoWbTX/x+iR
+hZaF4EsGbxCcNqQnyLDYlkhR0AiaiseRlxCsd/uYp7tPSi8VMzBs+L/jGq85Jll
6Rggw+Dd/pdZm6pJJtqn9F9B64pU/mmfrkxXtDJ/U1bcT6abZJEUBWhh1k/mjf8n
G9aRKRItuvXxWOZQSdb6XCBkEbIfaRVXXM8SCGiJgo/Vq2qkmOudsNBIc2OP8Jit
R6loNlEu4Uakd8KVeJraLBB5mZ1qHYROlFG+u8cb/OBriXFtHqgYvv/eUL4R2Trt
NAynkW7teC239u3JQXoasvcm584moyqfYxT9/BlKyUF2bH+ovNHlg7CQzU1Kh0Mo
PK5Ap01VW8WoRXCf9ghbWPm9Xr3TapJasR3Q25MMbncmHHdBuL/B/bgGHmh5jDaK
STEclBQ5Ic/vN/eJ6j64vlj1HK0S8+iGR7LXm6KNA5X41vgbSh7tvzk7DBdIOAfv
wEyQIx/dXY13hpnrjcj3cuNp/IyJjolZoNDIMtKWbvvvrm/SRc7ctFvO8PH/41ul
rj1xgdMhgQDBmIGxYAyYT6L47AsdHZJXGPyW8DuWtSjH5Bgu9jeKfUCo4y/CDLy2
f34D83sz0BcfZUdtHnOboqOLVdyC9rPXqWNiw8qe+kawGhDyQ42cq/6GdLDW1lG9
CulV1gRTjvATiEvTzW7gKLZob5SzuJ/QnFzpiyI0H7hG+3V/g/gOMGuuFfy6B1e3
F+xi848/D9EP3fklnk1O1zvmj2yhe7p+CyKzBtCN04i0eE3erS4ODMZT7MBGeHU4
KQwYUJqnGl3fCWN/wB387cjzxkkY8DswALTJpTw4ETHVRMeI0Htm3pnP/J3S+swR
Gv4z3wF3RUYt7suwNij4tTDLBkIUlx/mnbVZxFDmT+plIZZDJr9hioDpHwsaU+re
qHtsNvhwJNpSNgGfX3h/3FXd3W5BFcOpb/yJkdYc8OymuS+EBFIqNOmS+uiU5cXi
YZ+LEdaR/flqJmsNOCE63AYA5foq1OT8SUh2GbUcZGwGrGK85NKf/ptSPoMGL41S
9AjvaApE4D1cSImB387Vd9jZl1BmSLjBhpp8caJKlalQc6s5+Xoqwe8yvkKdj3CM
TGNPu8ucFfpSitLPThLx9ykQMMolSnyjAyBEEwGlfmN5lzEzA+Ena/1/4xE7XEmG
T6YdLyQ4MMwY7a6+Obc/EGcrVSZwdDpkGkPxEv7l8RE1DRlfrwBIlIZf7x7T9qCx
p/V9Pi8No8OH1/wS9hESJIZMp3lZfAqIIs5jYFoN4wdUSZWHHuUak1UtYA7P0Bs7
Jo+vQfDoTxlTdnAT7plzt0zbEKZCmui/WzFbQDcx6K2ZW1goG7kOcfiTi/WwEwr3
3XXXd3vn1AfDl3wqE/TW7UbbGMWstO0O19OI7rhX4brLMalVOWxoLk9fsVWSRBOr
Jtz5XIy+WmHq6aQIlEuGniKCY0XfRBq/Vhuv6rb078uFlBfOYJ7otmWS+48BMzqT
CHm/8RGTZw/qx9jhxPq5X6Jzx6bx+VrQybK1wiYHxSG9ea6mxrRkCnTtGiaDgl3f
ouI1qfaMg5CdNRcylWOhx7ssCa1DpbKoYfo2HN2DjLP7V5OIXidTFEVj2We4+ttW
O3WkEbAU6t7MQW3x5Ybl51K0cp8uBhcfLKWyKb5ahL/Oz/xC8n631n2kJ85yZSf3
/M+4lenQgOCaaZPGW3ycJX501TZRQ0g6ipbdm91NRN5pMhTgnQyQHMTEqBi5TV+i
KPbgBairpsjtP7ZKfuY+8SRSEUsrpxPzTpMfGgEeBw0vxGh7q41AnoNiPaNrUBgt
QcP/H6SzpbURGSsOgDjfHHvnnuGPHybi4BqBszha0FJcAX9AK8xtiTn2XqoaoUGJ
Oav7+HtOEpBZv/f9Ui/n0ax8XzkSSNRPRh5zPjC5lNGQhuGqNLgS+9qg9WTwYMn6
epmRgumD79dOAHI/nP/q4Gzec9WLpns35sAk7CPmhPG9LbMxqn3g1fgORqoZTp3V
9HN6i/p68oWBXEn9XRg8NBOe2mE8s3rF1qY9Y0YV63tLLF+lSZfZk0ojTUXOOnVt
5Ya04v77a9Vzh8vyNexaYWHyA5q5LwadSnO34kn0tN1d6x6S7Zd9GGA7QZhg1UKR
XQrN28jxGSe8WvyqRTHxof9Ij9CKYujlijeiS/W48bCivBUGdBjfLOnECyHkPFwI
FY7pGvl4Ypen4vQ1UAcpixi6DYywPkCtrw350mIeWiR+n+kHI1oELc7XpSf3wZS0
Ny/MEQcu04KrQgBDfNTq8KxY5l1PK++tE16QKB0DF/pxOGIzCjWYWH/owFRaKIUf
S0fFQ9NHQ2n7ty8KvQhX3VDpFPY+NiN7gXdonjmfanEStbvrsjw08FqqG/ZHfd0o
feiDtCzVy/m5Oam3GDC0KBvvWQ1xXSh0+WCZFESvR2RkUbbPuEdkPzUrzt4XQBqm
bklsizPbArsWXHX2pHuSy95nUpA2zitkdC+HpHcsu/iKVvA/nBAK/qNmgrLjKmdk
evSc5rhQpGspiUorvFdsej4YAlvdQrZL4eZmdRBwfACEDZqeomt65E3VRg75wkgu
ypgxJSH9ztqZY8k2teU3S4KuYT8YQSGGwYIFnllNIuFJ+EFDFp+sZ0FI5M6YSTDu
OxHazDF2mUl76EnNOBPztqEviu1PT6PYD6nbxaN+kxe+gSzrO+PuFOoUeO0oqaJ8
cXG5/ZclcSNMlMaQulPjwnKm6UG6BH3TG26UzWYUyvxFXjeeNuqJousBA/9pJEFs
pZUNIU7+URR8rc1aCCy2zdNrR7/xkr2thxptmOOq+eLc47pRvN5nOY/vD635P2sS
UP1qqPeiKyCDAXkqqmwI0WfgdVAAPkQ7sST5YfoGwjoTzMxaKtPuVdkXwbWMKV6X
70ipGy+Fydt8bHoI53exLyN4h2hgr9mdifSbeNJAQD8lWl1PVt/kOzV/JHJQsuAX
2PfwOPF4AuhUNK/Tqx2MBW7tnB+nZz0Dg0wVLajvgtmfgGOhTH8wBi5M/zSih1Jr
MBnPfIDxoWBeVhiBEZ5lGBA2EmPQau5MjSiOCFxceb6F/6cYXIzNxW/wZXAmXrwl
4Z+G+XsM5KNvGG99zP5KxxnOyl5zLBoNH3ML+vCY/CR42GH36mfwyD79+oUO8Ba9
yM6aPj1PcT5/vMpRWqCGWedXeS/mQ6hg/w6O6CG2uc6Ix/eYeTvhIRnq6mzMBz7L
fauLHx7VTPd73aEH202OwpBnzRf15iXPvG5nYjUdrk+227cd2QG2BB5biIqmCSRy
29X4lP1ClyNRLmA2lP4TBiH95n53m74UsArD+KjdFH2gnRai8k4OfjYaxUb5t8Na
Y9KjW2mk8MFuLUN+MeKW8HjGvDvtjMtEhlBK9bt78lIjRf/heHOICThlyk6MPpNe
Z2mOhNxmiYwsm/BPLrDdjxtuTBRTid9AJG4n1DMDR/HemIZFwvehB21w+S9kuGcZ
MwEK/iEXQB0z0Flak+LLvtJGSTmkDPR5nyOkugWxY71CwEtn/y9UmQyVQXIQl18x
mXNTUwXkcvaR/xxrTEQrCiDziMijzb8kNsrCq+aSCrS7FfozjpLznc/n97vHoXjx
wyYFbC/Nap6mMFunUUxhzRqpoCIdzu2YZpczEbAKHqYqtOcW2HwCzYCwG0aNEmOM
SbIOf5cxXUIAK9neec37iZEZb0Y8OD9E0+E6MzIwTfkoDKpDQ9EjJh8QlFOjmFJK
2A32vdCVoDtsw+QL+QJZjkXCK8gDkxyQeT4n2DzrJt7X/QpMlekYn+ii2jmESotj
n1xRL0yqginFOspTzPiu2+7c4LMbGzH78o63csShZ6L3Nu9A8Q3jyWo2JV6vi/ER
9K0gJVk9NTQTnMi3CF7VwHyLLmmsXU5krBjddnBPYLG9hhMtQXdV6gGLg9JhOfsq
4KrH6PBbEtMKTBeUpQQyagegUvMRHjVvjBOMqRZ17FiCd5V0oeJBtaXlFjWMPGgk
hzFjLrNfI6L8uuRe43CrPA0b1YCUjF923bMUzlroVz+AsEYckXUVEr/kP8GsybhI
wK/vmYCevYgDO4dYzIdJ1DKVAlO8ajcqsCs+utzwQUFyXnUJ/3kliyiPCF9Bzrbp
eLEqtZPyhmOd3QoS4lTJBWOdPMLRO/4JRf45zuyJvyvHnohmWKi2fW+k8niYWY10
YQTmsW98iyeMo4mw98/YQlDqshqyzgj+XOBtHOjxwzsAuRH4qPVALRaVp8R7LhTl
LLEF//aHKz7ra7+faM7pLON2ExAhYF0u54Q82Im6Mb1gwkaHrZzGH4AztMesX5qt
CQf1/V+/YAYrn28ZEao1mKQqJW41Ix/1pKc0viQe6zuQ4sciPDdSGmTtqdxFGGIF
RLWDwVRy55dWd9EaHz0sHCmOFyBqoqAe1PmZqSujKIMOf49HXNW+IQW0UHoS1cky
Tbnh6kKT+v40PsGwIXMv04bXgCXW5Q6welzh02EMZTV/0uHdF3q4smjo3ogYX4n3
TyM+fdshB4iPDVFXzBaiZeX3hp8IsTliKgGp69Fp5L+KC+GfhfysnXjoOHEOaMsZ
IqJicy9E+cHDMYquYHBEiWHYP2pRv7aW0lPGcGBDCKuDEWPSbjCwcZ4rh33w4S71
WR+tjYKneM4Gx4Su2h9ZVaJ7SjSv7ENQDd+ARlWaFUzvhdxsRlbNwQzgUWZmiWS/
JI7g3FskhhUUGJRg+hmlRTDPMtJnewqqgoUHluWeEF6MDu47nzZnD9vJwfszewJN
owgQegLuLAMvFCQ8cErrzCGa/H/ZtrxqPLOef1mu8acpHuEf6GNcZA8DIOsaEQ1B
c/zP5oxL2oVTg/+quMpVT7LYS76Ddrwh/uVawiTHYRVFvoHrZhzrQH8rj7aPyQen
BqeEUUy69C5wK0eJHadk84iOFJG9ebIo6HJIAxCuEIXWNM003QW/ggtApYln/Mo4
1KhSJkpdnhhu9z9sDbfLxJpCElNx+GhCBR7IJdJM5Rq7eL2pQxCd6+lXPwep+Q0C
D23neeNvGUrNmPFylpBor9L9pWYZ7d5vRZwo0VUVEN5MS1fWjVEAMc4Kk5HHfUsH
AJ46bYISvkP1CyTWIw1XWXjv5OfHxxwE+0EdF/a5uFi0+XNtls7voazC+OuIaLJI
IOQ/nPArFVfp+RiBipBdVRTxRZI5jVicIcCDxyg6qMhT2OcTl/aJu1+6E23nMS4J
sAf4fjIj67FBTvPxvZFWAfl4rqv4492bJ24LzTPpi2+8gZakacto7XaYGD/03nSw
wclH9nEVeG6NBTO5tzmRH8LnuZmpPoXCJjGyJ/seC4aMBrczJiBbo9Q/o3wPuBZe
l88MuZgMX24fsET8PQiulbl4LL0h5J6zVwbkp1xtRb+r4uxeKikkbuL+a+vSz7/u
wdAdFq1RZ3yYGVHG52S+uTWTXn0AIsKT4qjDV1AHiTEVY5niUL+jdUh4veoVC/iE
3uu0ut5xfFnn/RJXaPK6z4Mk+2RpLoNso90zxBTXTmuTbDS7i4iqmudcWpGE7Mxe
wNlWdzGKWrq57zCoh99epsG5E8Qa7vYJK6GwBHJ4Q7AAMMaSqitfMBgxlv79ZoG9
9beknAlNeZCos3YjBz+IFQjXH7XtAKPkKPQ9/Z2fcQ0l3F0fQVvptR7cDbc6Y8MP
+oRUoMW5j2btEAXguGlfDdwO07fobrWcOUvjsID4H64j68JC7iVLgKnYmbuId1PE
q3PHv2B9GI1ALEu8mOymsbm/WvyGkbnVhIe/mZJ4SAy2m2JHiqTv/Hm7MLzrddL6
QZd1XywBMepz6lzvh75y4XJVUIjDaoGbv5ovrWtlRhlaRk58qmLvW26jwCAG8eaQ
cdp/Cyzwj2xi8v8/P8dXRps9TEOxgw5l2TYLmWHvHNgIUUVNO6YPK03UaKGLxBzK
HOWuaTG60/wGKsLEuRXN5jLP8f0ZpWuvK1lyU710yPlYbZ33VxC9qklWjt8nLsva
tRlVssr+Ae6s5lFbcT4clPMRhrxEwAHcl3tZQfLXXEGyriT6xz7rd+Jtkep0Oz4n
Lk6HewNCAH9y2DvtLb4VLcgGW0WSnspiSSBrX4MaEPMbq74Aja5fKGwSLyQ57ZhR
+AWQ3crQXuwwjAA7rCHxZt2mAtD4/YK/8bdqi+1wgplxtPkwFkxgybYQJfZOlqJT
YaJhEjGU4cxIMbH2I7FfqmfNHNn5GYFLE5eS0kD1HaD1ppl/dKqFTw0iJxKqn7fy
LtXU99ukR8K4UBGRQyGasKMCnKsCAdqoJIHiOtiLTC3Y9gZp/3MBOk9x7hvg/dMo
CbWUFto7itinRo2GLfKEXfByQx9j6LFgBG1gJC7fWbNE2s4ODswgztV3sSh4fp7U
DEUpLQMMpP65nwmYLvfqVEwtinF0zD2WdAATh2QfZKWXOUeBu10ePXycyFhr8YCT
CXe2+jj6NjKiIWM0g6UPfFDqQBrDBBUtRRJJdgGbetY0LyKBFykXMUGSIbe9uQbx
y/OGigrORic5/WCaa7eDLDlqNRBP/+V4QGPcM0x1lDT9RF7EC97wikTjuYJVxuAy
sFUQ7iTCPBeliVfhEXqZ4JcZpJcpZwH7Sz4DdWKOj+5AkkayEDDrNn6UBjZQxLiA
EXyuQSJaMjCSAKjhAJViDy3DbRmmayloZkY6my63upv0GudxQxhDF/vs7phcDqEG
DvgGkZ+vRr0DZCVXupj9Yw1fOlpbk38AMjQKG4m75A0mt3nrO+/lHp3BSsnS/n+c
yDqRhNcw++jjJvEAV0NjA/rvVf+NVXMPbj3E7fDhc/96J9cSCCZj8fkosgh96Hod
rJSdC4fB3NIOvUG1kmr0q3tXrM2dgEyOfIxiuCI5rOXQYIR4BsnX5oASP1eaEorG
Am49GGA1tdCsLSkn3zvmTFcBMkECTlPWDJZRQdWANx0Fx0HH9BMPaJTMLda3j8c6
xeXq/6R7iG4gx+n0YCO1GXRaepOr8j9ZJfFrOInKEkxcajAne8OBcyhBOOTlHYhW
mD0a/J+GSJyaImn7cRbclZbTHw7mGGTUnZdz+Z/K1SnVgKGftfU7y/jogpy840gP
niI7i+dB8mzqK/SjgF1ftVC9wJnCpUNUWJD3DJWy9tcodW3NUx+G1fSfBLEcufgV
+1aR8qJipUwc1jG6pGLZV+fX1SfKLXQSEIpFcCVEFt7hDvs4yjr692Sh3WbqmJry
C9OvKMgE6KIC93xYMcaqFLZsY5lSqTPUAR4uuS8hiUFadvcTejHfevzSpByufXe+
ktvnRthzfbFXqZ6LIm3ApXhIOZCS6vfEKWOusneAd//G+AnCLuilblAZ+ps8Hs3i
HdiMALIlytG6HPDOsL/p6PiMbPQzZHulmW0JPjAQR9dDNwzUVGXr1grq8uYKLNds
35RjgTQQmp5WBSU9VTV61W3BLUDwJE1LrAWE6YgHDeWOcv0zE5nI54FdqVawM29+
+WdaBmzMjkptmx96hx2kGf7FH6aBA23yqvv95QZLdkH4uwEXjq+ppADzlTyrDMxN
N/mnossoVKs4XIj7zh9MYnlmu77fkjebXiyHKnqUgQRtul6xqx7EXQyImao8wxro
UPfYqEyKtC207SEpBkczM1JRRGuCwC9h5CrNiqJrjgwaDhwGlvd3EGgE2C3t5rV+
21Q6G93HvzG81inR8vbGmlf9e36z9+SrqmHWnwGJM2Xe9WIr5fKctA3p0/t8xTDB
U5ZLCnXPpitXddu/QDBBCDEe5rdbe9+Q85gOptIN4uPLvzMxdQmxHk3M5VzbT+3J
Hbaha6KU4QmVE7+lNYLKBnXD2FJ4NgWvZ1pkQiF7Y2cs9a1Je7DcvXJ0UzNn+Mm0
T/AGuIUdjyMc2geigi9stB41FUazmiSxEtlcdn2WLia88/4+Pofv9uzBsXzNyK5U
2b6/nLR2UIMylxLpi5pLGenvxh0whjVUKuRu+u3m62LjzhsnywSq75XEztVHRL8c
ANR2favS+rEMqMNl4VSDXcY4LZ36u1sZjHmQrNgjSkqnid2gDbQx2SIpa+MQutT/
Mw0dexsAK151cl3UIVRASHzrFMoNIGLLIh96cA/kSdcgtKInmYD2B8TEI7NMWDI6
xfnpf/wtrEPnmmGVRalvfFXj73r9nf05844fT8/zhdibr84EztXMNXAu41HWNRRC
lHOcsoJliNBOqwhQe5jnlQkVxL99PdETPQjHX+o6MiWhhKkQGAc1ENf46ioYeqxj
USj/1jbsDCvP6Q0bNJFIEkP6cQqxxeReo3P61W+bVXGa4nMHdi3hzQjukCCQ+1Nk
5E2SvlTGJfnDyEGUwb438mC3Mkuw9QwU+UNlrNzdb2X0K2bGFz6l8ke/DXKflPs1
Y2BO9uAhk3gfDGwbvKxsqaXvYhwDj39XhEfiAjXAqDpcFHv2o7F4R1QK81nNIEFe
G3jwh4jRkxc0pG/cLtQLvq8ZNSQVpab6uM+yhwkm2IS/DDN/7lydU31dYNQyx5eI
2eokizfEwY+vkO4nWR2YMSSOKz873zhU+Ja5YRr0cTE3KjZClbJL9F+JvTHZAdde
vFQ2ti23zOd013kP10+3zG0PeuRuzkEF3c+xEeEKlQG5y+HasW5ohIBA/3TrD4gg
sZxdx6JF5Oc9lT9HU0UbCGhoESl4P1JrEf5lcWN/YFFagcyiP5nHZtVXJOl7P+KN
d4W2px+CfwFoBJmVbsNiZFsFvSaZouxaAXy09PwNcTU4LrQYgxrJEqERGPQ9KYuJ
ffY/micwdrMusdnYvRXRwOYbiRDMWvM6PBAIW0vtEB+i0tWbFph1n+jaeeS2T4c7
2lkk8Pfck7SSQGDV3VSKHstalW7V63tvKqjMvMpHl87EdyGQiOPdezHlmyrfujf8
4Hq8ZhK/aUCjibDP+557/AwI6yRzVTEuE/usD4YpvzD03ZcNDb9IagFK3y0N+42m
ZV7VCvFvuAKShvCHjZmWbgs9uJ6mIYDbT1pSwhZBMnbS6XFuZKsC/+cfrwMK68Ue
rgECFbMVvZcvR/Jb46c2+yoESWIYDjXOW3iO+megn4g2ugqP7pqHSOu4Z46Fwwv7
KcphFbzyQkz/CktIUtcNIywWMbeC4ZvzVUvdbMi8pGnBcCyKw9u6gLGrKLU3WirN
6HI29VDHvNyMLjzgfueYWFIvwIV5PPp/cWni+u7BfCDDWKUqgKN1aCrAbkDYKSL+
Dy513SHUtmM/iZoHIEsd6iFUSD1JPOZ0GeS+sJCaGIdbqv/J5FwpDC94Kd+4MLxG
mdtIYViD0Fkz3E/bXxxM+mndLs7eTprKdr69RKu0MKYScFbHlCUiOoU/ucucX7px
KlCDoE4DlfT4XlUI05Cvc3cRVM4l5B3Hkzdsz+f2bzBemMLhV+6LZAzqRw8RBPYO
3zUnl13JQjSvzOs4XqLAwPZsJNnxlRb6CtBiWqRFes4a188Bwi1MA8DEpVaaQQSG
YGw/maim9JMhNVky1AcWIqxN4NGuCPYDPJNN/qw7xHEztBZZRW0b15wMQuJsaq1n
fgOUzjzvDEidkkvdH/EjWZBd2VaDanwwkCw79j1NRFQBxE8sl2OBrWz/fB5VltxI
Tg+EwgsRDu/BGoAO+lzEN3+seQDEt7SJhqVMb+U1LeOW9b7x7FiVN2/mkcbrTioe
/61BEf+GwgGz1TFH5Ome/h8IoCsWi8+MLS3HOidKQ3oGcN+9hMSfgayaV0aGcSx3
nlTuuEyWHMOyqmEXpzmKTJlVvxhmqmcfML1s2QWwo6POXHmqEWHf4fen9PEehB5r
i43jy79Mt9gV2fxhB0twl4yYDZo69QegC8veFGr7XwOxMOxL3rmwcfO5VC4/gqhl
u5UZ191WxEwjlZOSmkT8AY5MppbVvPcxDAALFL3s5UghZ4Iidvmqp/pVqh4M/BY4
K9snlXuYpB6xf5NbPu/DYjlJ4hPISxGZxWCjckozhe/CAhpU5msEeQjg/UknAeeg
pbXRGhur+/dG2H2HdfDM+OOGT0h/P49RNVeXKmR9+E80VRglJOgNNMxfF2A15ziw
hCS9oYLAsu2AAmZe/O1EpGZeHuE7iPpZI9XnszfxR185qlq+iniKvp51K04AGPKQ
lkfjb4bwyS8VoF+Rf5whx5ZVIAHGU7WI8CDn7YlB4WhIH0SCiWEPAzTg5RezuEHr
cYfmlaESBphpiJ8PSVmm7hYNz4L7I3WwTifFIwFhULsNiKHcdgGz5Vf4ci1BcKlb
Um/kn8374oXF/4LJU97qL5Uo2CiU6rf7hmoRqn1OXIZEtbZR4O4GD0X+IqFxfDMZ
aOZWXq9Xjs42F474R/E/FRL3uZTGL52FF8BeGeXW8FJbDS1BGtLQhHkku3ylxpmq
amDChYjSjF9MlJBN9I4qWvz6SvfEVui43vMG9YgcvwdvvOgJXAe00IkN9AmRZxIM
teU03QSa1Rce9l4MfuS/AvDoq7whnaGJNmQlWZYO4I/Vqbq810xjD0KrBzWuY7RJ
X0ExAdkaeHFfLrG1cB07OjtUm8F0bP6jCRDYiRPfuyi48P5qpfXdII1sKuzPKssk
R7h+nmNwHLHAuc3p11kA6Ny6xizMCpvWmOW1uYzqgPRjGc5nmz2mJZj8wHwYPg5f
n3sK+K6vghJxyw9VS3JWNYF0CR9t6VsDQskSiWS3DdJoSTxJoK7bVAspE2EnGKR9
mQuNOEiK4drLWXGY6Jx5EvCvNOsRZS9SR2/twm6jwIPEU/R72BQsKlfZJEi6J5a9
CU5E0w+Uim6JO6LPOaJnMzEAwEdvGqAUtuQeT9uHXId8rGxTojEZM6v3JQd935aE
Y6d67AmJA+Ti+8U0Temx0ffPzzNc3i6FTAU2bLyoBGkQKc7mDoxWrwZZ+WtDYP06
WkzSczPUsNRrCD391QfzYGer5Y/tb8d76fRTgRprHmmAxEO//uh48l2tzV4HILzV
6weQfckFv+QoLbb9PVr5dd8EFgvtINlQ32abZ6gU/7Rq+y0tUc7Z1YJRYkUihkBm
pmzpC3nE0ZihfBnSJ087X9UfGvKLfj878ODnjoEQ2MvbmxReadlxLHtUuGtXxquk
qWr770RHbNJ8giHhiScd8IMSCP4wbrEeEfwRVCI3gdDGtUbmutZZhhbPQfZqUu02
ndsATzsJY+byUynLplJf3KouTR8y1SzwCRk1daI9yf4xDsOvtZD486nAQg5Murgm
vl5F+voOcDs0DNDKj7AAW5CQul+lI2QYk+3yogz+lBhb9WyrD3lDO7v1agGotPb6
R2LZw7FWRrG1XbzdPBKCHPhUN+LG2oyC0O0cVT1X4rzOY7seXUtplb7Go/zDCJbE
prdKdFy8DXhSLpLj/endF0HBZZlyBUaFq53nYhU5ZCYIHgGJU06YYJCCd8mQfICl
r91LjVYl5Q+wHIZE31xfmdgu59QoJPb0T98mt688mJGII9yqdkTD15zvlwwa1R3V
ZYAHhLM7COKCVVThnO6xppw1DqhOtF9HR4EDQlikSGoRvw3tEop9s9lGI1+UwotW
m9Jn1kJd2kfh9NCzR0OzJy4ysk0sFMXGo/CLc0oPl4QkVe06AsGe3mCYu8katCPg
CMNx6G58F/IDj1nsKyGdm9g/d3MiASi3ebUGlOPPLrlzl/cQ1YFIRVPgQZ76KJFr
jeOoOLpLBlHz/YiupMev9dg+6uAxpnObwpAN/d0/ULrvCwE/0yhpb6/5laUT/ktn
HyNWSM+tcMJERaoj0wCh6D47Flo2KPedYnBbsLrWiBpTcQTiE0S/wGSF8lwJIKoL
UOfnzzeNUvu8qroDv/NcZpivJFl+xZVw+yYbNjxcV/bAV5JlgJSRpEaXKKaTKLwW
XQbK31Ow+2xylE1uzYchwGDNYfxHHTCHMlUP55yCfWnzFqb8nw72BG6sFIEkBmMc
DyZA0c/LYiku3jNfPIqehblZ2CYUOccgJErOkdEouVWI0Md6/QyzhwQqe9zyBr4R
nmio3uSNIg4oJDJyvVWbjwvZf9fpkru8rU+T0GEXoBk2pJEZdFSEDAy9FQH5qdn/
NfgoEadt30b50+m4M99YDajxjqAKcQJqHTJ7QpD2qoJ22fwwwdJRl1wKKzQxFGuc
TvbooPONf25NTPto4OmFWpt7k2iEJT9Ph/Afmg2XXZytXDdrq9dI+5Y6+mOhYE23
vcxc2rst3nFNPNZh6HcoNK9WES9/zVjTVpZPls+2ZO+HpL1Qm/ooGbv0mZ2TSBcg
xzRzAFsH0uOUr5+Qd7dOwS61+POo628iZRkRP3dkdkqYc0xJa4MAvC7dp0DIdMEP
u9IYw1OT7TTDcuwvJi+cRNWRLq2kfL4ENfeGnQTxYUBn6BGLJ8OOmBEV4lFu3kIS
xaTHLV9/9uv9Rvokei9nH7D+ZZJTPraR4jArNsuhABjtZTIoBCnYfprfE6qD8q8V
buCpaDBSzvkoVBDJvZTuCGTtBjT7PhI0MTmq7rKmmtd3ORnjqYh1lx8I04+wLMzw
H+Q54Q4iaxds4fSvcsVDwBgeZhXCDLLXc83vsk7F3RnGCy2OciLnEZo/yp0nqOgx
T9h/NnXw08F4ELEYt/bF55l0T6+b3CBx8wVEhceGkIdoxbT1dZxiaAc8JIimVK9v
+PK0FEIcRMOOvwUevhRggzjb9l+n5HOJOiXeErPcyva8orgWwgGjnQa0Vwz61Q61
tLg58J+V7rhl24wZBWds7bh0jv2ocVJ7TZYkLnE1KAKSwy+rb8cJltkj7JCi15ba
hckKd+wHyGaVSfp7pkuLOBpMg5yCjjJK7tn+sgfOu941BbKUvdwiZBCQJsiUM7p6
Fgnu0YaY8LxBC3O9nUamnDVGbkfPF+H+5dMAJNCet+Hj2iQq86Is68A11+prT4My
aIkm/n/SohV+P2uWdtyeMOZcOGLauVgwn6w6amElGNfdpsX5T/ECbT0HktFSK4BQ
mE/JR6dtTMLAr26f+wiTGFkxHoYl9MtLf4VhIx9nAK7kdRHfou05W2C4kuYZ4xFR
dmFIj2uIhGzpN3uldgPeeBKFKhvO05Wr4IsOz/rS4293RZHdW2Qlt7GiZlij5LLw
UShKyoXz7P+zYNEiSnmS3LE7QuCkGrOFhmgitoNyl7UQm3sHd+5Y6NN7bkzwOibS
toUND8yK1R+IkBLVvje9Gb0s3/uOuZ3YLU6XjqCS2GyIvGNbywQdGKfDxikolaAF
DB5WZBUgkaFp5ybKe+I0UDGu3WM3YIKI29sloY3Ey0f/4dlrt1ERr2lVH8kyyTwC
mtalUeFwCI6H/uXL4kI4M8n2is7f7P/wQQdPlHjwiLwiFh03Zx2XQpiHiVqXddh+
9nIlUMLGVbJiqNZ0OI+A1eHmi0q8gnac9HT4IDuJczkPHeNxuXrdvTouLTci3wDA
q9m/vdBv9/7+RMj+DGemiuOmd4tsrf1UCfLxKCAm69vyyIFl1gIW4/MLcfTpI+3z
Je6rzp89b6OTn2xcAI1Gt0VHGXsHG0Rhd4w2PLeDbm+ipvjouQvAtS2mCSgIwljx
6dNRWx9A9ByBtSw8rZ59YH29T8RUj+TQWWEoRQlKwKos5T4HBPsl7X23UpEvqsnT
KnzWbs74WKxu0+Q/UFE8RLX2fkinygwEtffHPxOt1ZCJWxMCbTbUae3NKqcGVb5I
UGaOTILZFV6QxIHvIL1G2R38u1sMqwzMxW+EidIh9sK+E+UuR9LBvthtUQkdHnOR
M5BjbUVZvj0hI8EMdp9lrhcOu7QNN84FTpYGwFy6B5sJC/i/lqm4RT5ZjdcTxjzc
CW9hFPsHtEQyNZqthY3vqUD4aWzVMWF27gi4gdv8LWVg0MUeX9xNRpwFx5NqTtRy
7EGPqW2hQc1ZHTwG9CmWfMaa8xHfBylBtwAw60QUZn/IHVLG6HokcT3EBJodGQQe
3m29dtRFQ520bwfeACoQr2Edp1V5AXuLBUCx1zmPnfjrE4L5bnrz/B4MzQBQDSEy
I0+3U79PuJGNwYhV5TPNjBorNesul4D0Kbgl8o8NbEdikcBY84NQVE1VwWfyZ+pe
rA/WlABbCTjNjbvv6G4X+PgUIeOBeenrEMkQFqgPgazp5o4vwVZD/R4QO+WwLVYY
htKwvhgZZPDiRpn8XWLAUpRljGc7gHriIZtvuEKU05PHUUZgEQpGWiVmqDrCD4W0
66n7U3Jowh5mDBK/kQPzOE5PW4rO7l3eD+/Nz6GJfF7NevwuEnpYBVXDmFCjWzrQ
CRzoIiTe4CbOc6cMqzogYuaUbNo18uq7MeMIHFIx86d8GzgEXbXgarglG7j2+mLG
H1b7relxMO2khI0gOAKUdUEYVNskNvy4TxKYX8b4/wEsXDINyRwWtWiUlwNVdqIx
+d0DWoIp6n5zGIrkONcrcmVx/2tGX6O5wiNeFNGyL7RXRQ3cA5OAZqNCqXf5Xo/k
ggyw3xvmx+vGFUFK2w3lFZDLwtXlgyXYuKiCrD5hnt2qwUXX2WURZdBg0DQOgezm
toqQSWIE/aE2Xiuu6ThCpdkcfjPBRcIshHtqpFoI4cmAu2awHFeLfEAVOhnBzoDp
cw4sUAclQSZTf3KjfSqys/jPQ/IN14QFGwUqMxaFcTRa1XYts2EAQ0ZhmiJbK9C/
YUb4bECVJiQ+kNb9YenoJRhztV7iWQkz7nt+C9xVGJ+Pj+nA+vx28zwoJVXjFtDd
Sg1DD7dlWH1M1RiK0XIADmBYK9oPoUsim5qvRD1ZWHyXLeTX8kTo/a9snVtZWOag
qqblzyxPzMc7a/2Gehm7J4fGr7cazXWUNZ+oSowj1+XVwhVSGiGPKe4U9xKaFcTY
JN409NJG1yx9lRhknV7qRf+poRM2qUnAv5qw6xhaMt+QrYyGD4hVewN3LzDdPHI/
kALK0ltV1WZNDuMIJHfBqFIOIf0e+8eR9hcBwbYqoBHe5UrBH58RWX90JC6Q4ABq
38Y3dAdMFx6Lz573ujYviTActx7ND4fnG5dsoKxIpGp8s0zr0mFeyt19eeBcOGS5
wg5CfNzYwtkl8VwYXy7xBsx3W+hlQaWN1+31xp6KDHSzJxIoUaLZjXgD5uO92+X1
wi7XjmmqmuOocdhz0+yndgaD4RonOUgRwlF9Du+OblLR5joiKedRPlROtr6hoi9k
hTUaf/3KSjKfbjpbBudSeauEf+l0ZoYenQqf80lFu0kl6Vv/oZjjulGx28aAFVex
JhxQ1HqiFNwlPd9/01dI0ycZdWJZ7w8AK6VNHhXjjP5sjlGjeP0fdmI8gFApDI41
HXwvRm6D5oz4QQkcHa6qs80qMfvdCb6qHIoUOsf/qGL/ZApObrL5BCUG8kISUZO7
i88umwudbKqAwx1hgDKUS3C0rB9QpJJOiWnwQ9WOBgyZsF/MHe42/VJeLd7aV+Ob
QFnnX7iVpBn2JOvGgC1c3KjiRqZ2D7wJRu+ijL3fUrqXcyq6aV3Lymkjo+HzairO
Vjf3Rio3tl30tB6fgN18RCLGIiQiMjn90MT06hONuNggHOztFzeZBLHiidM7Z4/r
S+I+GQ93hR4rJlkQOt03BBpx1TaW1p6VtcLH7ZIKKBHCERlGYhDUg6GYUpVfYmi8
EaURQGYiaxOU8V8k16sCO100z0+bWhBdxz0FSRTx5JQ3r5I8ZNetTmwhyyJqaVfB
Ddgn7uFFxYSyd1iR3Jj9kn98N3xJvm7obwgwinCrF5On4ZJgvB3h6wNWRmol0CbP
aoElftyRYjkU0VeI0WNwQPHdVCjwl9YXNfotdG6gdsy0fDZpJStvaV2lXnRe29Ap
KeqhfMeQGsHhhqD99swFI96DR5tBkQcOToIsK07VJLDmpOPz2OhuR06aSBXlRMd8
C231cYmblQHf4ULpNDCIYMcuttOeCYlAgC2cnl2+T+MAFzzQ0v8wiqcX7bvuiovv
rpdprjO6gwE6V9yjVFSeKfHPXHrAN2Odhod89i4v+PReaZI377U9YBuDvsi5wJPk
IeT2M3xRENCenNNBc9sq1yuD63ujvoc/P6oHgI5F96dd/bFSmdmKBZ0MyZ508Mov
Lj1sIFB17H/1QSOGoG+rm+IsBQET+wuis1rNHcOGiVndSpYFbMlOwYPARZQ85/k3
esllv/W/OAU3sDVcOd8uGd3FCqDeX4BiLDCERcUmUddIyJE/xfvQCvYblAs5wwKI
sMgrR9AdrPiBwCm7sujDlmAxKxsTtingK2k5GMsRwHQOdX43bTvY1VMMb9DkeynP
VHaUxqLMgYnfYIEi85GthMelh0fkgqd6kdbK/yB2rStR6PJQwv/5np5J9DcFmcXC
m7lzZRFskcHEhkNGRLlk8A7j18Z78+6wNS15hO8zeAB0ojIm6k6+Hs6Dbk1u/o/s
WZe2UP/msXdhiDdBoFU0n9IKj2Y/4QgkaRPj4cjPkgn4tetc6/MjCC/fVDNfVXfh
BXgxDkgyoqA7u9gcVqRVKk7qsgePPEaNXVtE6ikiPuA56inXtuY7CEj/2nWuNH49
c3ZvG6THYGZmcR7m4aGb2WkXDaHYafLvGsX7jYxo6PNWLmTr7tl6+mqPxFQ+b3xx
E8PPmGHH18E6+04/0t9lvmEgleAgjEJuLFBIs3CzwkO+HTXLDSJL7XO1odp3Dvhu
i5qChEYPFUXCyxVd49S8aJI4N/u/zama4vsECEHEWKgV5sMvDssbn9E4AkR7Z2ev
be4d5Krw1zQe4WlXrUppqzH9k/PY6lFlkes/jBjYYfccpvFZGAJ/r9HQzIICjeoS
jw3qcAgdJgBHyJhXRM967JenbOQl7PumRH/0me5I3MyygXKXdIhruqr5V1eEeWk7
a7oGPcW76jkeDoNGpd48PJ8GB0ZQVU/Xb588kYqb1Dd+ab8qKI34d45O3CSo0TSM
aq3wSQvWLt08HxYT1/gcTQCyuQqaJzxuPt8rtvqzQ5yneRNGU7HKTWbFv2awDVHG
mR5F+uMhZj3YelmbUNM4joGhrDOvrXrIli/7PiRppKzjGUByx8TDOIJMeK3ZFTfx
MEMrWRmHwoOoYIhEfdVI2Pi1sRqe8XOWeZIRXdV/iyi3EtgtwrigP1Ch/PUaa2Cx
9PJHaiTNU/fRjuqfU6gUM1vLNUNAhDcBu1C8g/LiST/d9BO4pG2s0miEYBKoWdMq
nPCHppLntwj9kS0GGCGRIod1Bdi5UPflIHfIL/zDPh7P7oTwOwzTv0LgJygzHdSf
D8Y9QAOOtQHtsK4avB6R67Ms+oeINnxf+Z078XKGzGuwdSzGtH8tIzXFZ7rSctvy
OQDPPtnptcLiYoA930X2aI/MswyH8RhdcnZO+fe3EIlruG9lFeOXhdgAwzYChZTl
fVWoGgkPz7h33WtlN0tfwO/ZKYq2TPCAA3td1xjuYySrlUfh1wj4J3PBmSK+r2I6
rxloyehMvaWJ21Aa2Vi+8zmU3nZu3cP2IMXIquQ6puSglVIhSIe7mzRlP9HPaHel
2iduuRH4IlHNrSOB7L9yg5USJUtuxTGpEYOHxY0NBSdEHqH2MBUAnWQnK8FipkhU
qDK2lA1MAYHj5AEjHLEfWnBAuhE91n2y9hHtmxnDDjvqf7dZuprP3GQBbKftoBOf
VX4QJJI1fV+ICw+wgpVQHG5k5LVOlYV/p7cP9Blp2R/qlBCMBHfJnxDZczUHH/OH
ZH0Zf/Rf4nzsoPC4GPrRrkGhiMQ9ZoIher8s07Gd8hNF0qSiNn19R5Brez1VNnhO
sZpPsTi/D3LFrKMUQboxZbT0spgZQBSMgkpa0dM4O2GfaHE70ERp93umbXU4TZ2G
Q29tzF6WGyXSF6RA6yAuK+m66BFy+vGEkt1ajQkF/HYVpmdmktCXMBl0JVSL9X+7
tz8ckdxB40n+Yk+NRUPBe0RHxK9fLTK90b9wQ0BMwo/pL8IDMwhhtHIisTrbkZFs
1n1yctZKMhhxwY3pnIn9OvCo12pcz4a5Pzgt43cCEXBT+EvhXhb7gAYbcgyqJR/X
jt9v1NwJYVsK5m6PxGpmbypHy86JddJ/dPyOSoZQF6ZRg7/DwVgxKrTU2+jgmT+f
mwejYIPrs6zlOowSvRo3iGbhsUpbnwsRlVXrvfNxhjZEN+a36DcAQ9Ae6k/wN//b
hMOMb6rmNLg0iTCk67c0tPI90GweezNOwpmCMtGNCPehCgz1GqUY7YSJQEYqV7HV
G4wqPxoudN2Im1gJic6GUeN7MjhWQSbYMq66jHqg4/m4ZUevRep0LkQ+m8NlpaXw
xumuBP2mc2GuMjtMHVCQKvtJwKOU8ty3Fo3I2tPLeeJxKKMy3SV3TfR4t4a9PTsV
TywQpfu3MZMm9Ur3qLa3/8UFWxM1Pw6hh0EdhKCQFCiwzb1Y01WDDdbukVud3vt4
l0NbRQSG8RqjSweOK5QEMgsT1ApeqpsRJdxSUYeb2XLlDekl588zY8sYovMC66A1
Mjdsmy2mwvMsxaV2Vj22quq6zf+ydYx/ttv3SXwHaShk3YkgT12RABxseJ/pSXB/
CGSY6apbD2APxXsaxWX5ye7LKjqZHvG9ff65L/5VYcuTtmVueGJ+2XUMlypfhaPk
euL57JXMjV0kzmUytEEtz6AAXw3yC78iF9I8tRJL78ylrR6H+o54N3PkwDD7Uyuc
krgbRxasCQ3Td+dFmSO1N+ASewB1QGM33hc847AAVb/cQwbHVkO6iMEEB2BFl5GK
yQM6jv9e6rs8qTqzGxQuKjEFLtIhwARJViK/ePBSUOEUr3YkrW+VngxR+uO901t8
yQm2achodOe8CVoCwKPhDpE3MvFyVfHU6RWIQqzZQy3oUazlLpBjT70Pgf77p9OM
4BmU3poG920IFsP7F17eLhd0hNcJCrTkSwqY75krBy6eoUOE0BMAaej7NVkLTLxO
Zb7p6PC/hDHzDn5IcJYov1/RsI4GsLtFr0aXYoMNLf5Bt16PDZ/D4tH1b8DXQ1p+
UXSDNxEV2LIqalfrecjjGYVPEGtujtFlZ+PkTt8anZnlsajWnedPwZRWiJrNs45a
KEYQ/1ihe6Ip2rXVux3tQupHnYugpj8GmVbOh0byBGC5RrX3C6YpsmnxokqK9e0i
d3vh9te4112OAZwulJPIYT15Xl6AeKLqwJE/PhB5vHtEoEt3acMRA9caFAepIfpW
5ucHCVYbpAh6GBTWHNoze43oIlNlKa7ByI1ntbbCaylWAWyEs+iIi7yW6U4zyAkM
ZA5t05LvESZ/vxvKu23lNSK2rWsE0WnL5PI9PtgENedOYpVCBInDvSAj+6XB/GNq
4Wp/aS9Gx4DaTUSwrVNgZ2/6w6TIdHjtxxDlzQNvf9U+j65Cyunei3Q3iM7mcr55
ZDNG6gV8c143IEeSCkQfMTgG2yEeDN0vB21pq2bEGL4w0mE8VvlchigJEcOY8IRN
k4AzoJltda/HKQxXVTqE3hG8VD3LWjFaDT9fffby1h9ztmNP8ntd2zOd+R662UL6
fG4lBo0rfBYIQe1FqLJU8IABhNfr9CQ7+mET6llrXf5To4n/RR0gvogfUhebwbIs
/C9ukg8E6FIq7gTVRp8Hc7ivR6o6Pjk/RDYLBMGKXfGs2oCayG4qYsek5zq6+pDu
iIFk2LC1LgiBD7JmxR8SyPwjSQCLuYzxkozqc+LWkuR55V5kfFb0PafR3wmucOOE
0UwQGfr1tMWOlSH81y66iNykPMI5aYfvT3UvOHfe9nb+QNoHDWSlZ4zH76N3EewS
vxgPN7PMFwD4bSeWqt1YzDPFo7GbuoPlpasfwESxiKWZ/wrq6rY5Kta/T+YLlz/L
3eH9NLCc2eVU+85LgOYgoEA2nzXVtZSY81yKcI6+xfHfHO4VPvSG14fdHHPeg+ZQ
MGlDQF/7fR85V0YcM3AIbsv1FKnh/6/fykQgHaKQl2J8Ba6AyVVQjZ3SHLL/NIXk
SH/94nhbLbCjWEVX45+cKs6Nj2MxONwRrltqntGWmZ89LSqk582AmVH9El6xwthj
BzRIz81KCBDIfNA11x9lzIGFFXMxKAJoQTRjmgkViTYfABYlrXZ5jQwQFBer7ScO
rQVtKGeOlDUSGoMgK0xNJ30WM3dhiyo8WDdsCWV8fUDIs6xtj0nTbrV1OTt/nhnP
egCldlNdYYqx7Bt5RTvLXdeNQQBSGlNvPSJnWtPc5Tn/GNcAMNqZzKth3YnJ2DeL
ifRm0UYzqPWO2Kgiy62aNSU4BrIK7a9Yd9AziYxvVqTi4IxnKA1amH8B8wPhauHj
IYQ0qQwVx/t5f0b8qZ/2s3m9fqwNOTmbqLdJFf4GHUINgcxmXUoi539lIqNtyzvw
p7/Pcy6aF1tmoAH7zAVDtuEY4WzNZ/ghlynqFTSz3vgXjz+p6XTWan0g/NVJrOt/
p9iYO3S47qN92usOMo4R60gFju+auNSRrdUcpTZL97fw6SzFjsot8cENI9WZWv79
adIzGXwer5UmoO97IS0I18pC1MaXvCQH4x/o/Chch1XjayjgKrMyI05E6voWLG4r
1xcWu9lhmWgWW/0BA1qqHT6wPGumNjq4zk/IRb4AVMr0vX9CGMGyqTYNkVBkJxSB
wdCQ94NiKAjQHNXTdMPX70HtuZtk8J8AHzAz91J+rY9qQIvlBL0YaaC+ZYCKZrVN
yra/cy17RtJcQYzTgHZgUyZ4zl2zmAo2+TjLlu8pxmx2/tO8cEOrFO2LJ3rUxqra
DqntnBRZ39Sr/VxPnN2Jlp8wNYpBQAFrlNVyXM0cmBokI7j7JkIYgKIlD2rRWPdk
AgkUzCvtyIPDXor8Hm4Iapnghl4H3fV73mxvXKhk9GUpzcHw/deZbKgMv1RRl4wX
Nfwj+rZr4fNEbo2yGQCDS/1zQbL3MgruBpJZSRrmp0oCQJXdTqNRGjVN2W+BkL5f
7lRoip4O70hLW006vMbBqOoQcYi4BaDqAy88uMTJ95EYEOm+qBNDdTmNL+9sMq+v
gXdgE7nMkfjgZAgdIzW/P9xsUoUDSr76bOb8zftzqrzB/9KXWU9eCz6RU6BNXbuN
QWPOUG8aR1tLqzG7ukJtJPoiRiAWu9qrj2Cw9NFFYJKofMqHaLsh8twqXXQQHw6v
smqKO9frg9izGDJcKxvl64BoVUrMKxaekqZ/KFryxScR43c9SF7Uexs2vCXIoAzp
9A+Crc9Gni+xXS23FsxiWyaDPzk2Irx8BskLwiHMSzwEYKkD8m/G7KE3BfH8uVt7
WKxLYNBhfexRGnj6e+EqAn5K2Tl9XptkXnt9Y9eXo4CWxhJ+zPQJmrqcAweHlW1Z
uVKvoIsTm4cQI9arHhPLEMPd6DwoC67HYQcMdofgtGN+Li+hDyYTECDVfUbrebRM
3/qHEhq7wcjWoGCeEe4StqoaEPkrZMiTbZf5UZrkHeqihX4Sla8vzQZNeqyqe9y1
tXwQjRrhb/AsUwyE24JuGyPtg5QTNu9cz2OWmmkKZ045h/VeoMS+BBZvGC5GRVMD
xWkanoRZsT0R+yn6zgno4ZRh26lTMu7hB/5yOh/MMxs04wd0BeyFb+fh+tR6m1b7
mdSd98ZarNBhlZZI5oVtb1adCbzxv24aodre5z1NJCepA+S2k2daamy0vIsrJf1l
h8GjvqOwSFbS0GiX294hk7H7UrkLN4RCSpU/TP2hBZ1w1ALyQRXmHDoMbfBoTmSX
bt1wvjD5h8LEHBbSN9lgwQUhspYatMYJhEAP+2NrXF2yoQgINc/1czXJHTQq+lUD
xd1Sv92mWGmBapgtDWZT41pE39ZQKG2Qe9XGcpINq55xdGivonaq1mtcHLgtVmSq
O5Ej5PkLCriN3PJieBtAdcSwt1NhJbjVoECvOqLauygZCkMWoscvxPS+K0AuBNj7
bItMcAZGIUEbc1haFoAiK97RwELU8UNq34dS7bJey6SUMvPuGG0OaFJUrpWqZXDZ
AUaRwEtNYNpYe67uWaxyYFdClh+bNe1UTNCd4khCfhPyy86Pr6FSFdSQdNR5YvX7
s/DBi3EBPvA6QBFefgMlrpL8FvGznW1qgwaYEhBCi37OyIidiITuY7Lu3UFlSFS1
yTUNAGEHjn79gu2xYvvWmdi3qrgKzvsM8buf6k2cBPM2wpcNQ3vwpfQYlsi1PSPX
+Uqf7BvTpxrDAVpeMn+RTXq8XVmdy8Micb4hgk8t0mEXN1FD0ZoxVHn4XR67dtjq
CdzLDnVZchE/WYRFKeG+uazBA4NIcC/wSespFqImzkv2PATJ6i1VbCr79DG5j9J9
5cQ7cBjjTIXGpJOijW/S205mrNkpyFoxBlP/E/QieEwtJOHyuK7VxsXLg/J7TiUv
Bpncx3lebYSqF2oVPApvNJYDHv5KUHNM1OI9LMFBoTqeEEUTxHTtWKwUy9FWR09/
gMxuJh5P2Q4b1rEHAqUY5MzHEoRp39rnPm17SbeXOBTR8j7enuWZjPD258ulqtyQ
pVbHXIm2q7uGE0GRXSmwBJOLPJiU7mCCqcwAJPeHcNtGGQeVefZaHaxyNEjpCdU5
92hFbWpo/cYSxZBbZrQxzsDODSus97Nf5a43tciPyTmm1gwAhdREZNwHY/sVDLOF
Yv46WfAYSJoWQTLDFyIR8A6j8gcIJ+EIjdM0QJkF2pL3/cboQLWkboDUT8t1aiNk
CfKQdEbWdRQOwiPaXkw4PInEhbZWuzxu+zgNsNcPrvE9rGzUmeH+S3TVJpxr1PvI
ltSevOzWF17AKPI0cy2qaorNezjXr+qUkf0LySGPK3IhyIBz0aCZes2md42IJLdx
dzrrgEuql+Ud7atGoVRXATA+z/ReO0zADSWzvQ1KBudnNvNA2t9XoiUhq3fXe91c
kzYRKra4q0v/obMczyox8U2D2KKQsHuxywPfVIA+ZRGeuC+xtaHPPL9zmNLKX3v7
lXScdovOZaxXsGbldieCVwFS74DB48EFITh2jVZilVnqtsTDmsIWNEDu5jew69Zd
kuEH2L6EHmyELL2I9luGJsol8K446lfvSeB8DYL8/C1ouK1bPHu3ooI04154DCQ1
rj1gvTiTKb4/lwOqoDGWoZaqVRPazLcDawhKh5Zge2g/FWzIhUhFGkiQAF98S3gy
RbyzynKI+vNFEuprLK1w9RguwSfhfR+8pZrsv6GZJLtRPQqkQwkvHym+yxC+vhAq
ufVPIWc/c8Iu4B5/g411hvmcYbXFC+509weF9HuIcSa5UVUYkjG4HsdWW6ujAUlN
jQZdRoVf5+F8iCUo9+DvNxQGFw1z0XsoTD4nIjKrl3vkgPjDoA7RbbR0kVTC2vVS
7pnhzVUZ87Av8tfVgmnAtXC32rIQ2Uv7ssTto3tvSOPLh5w9rNT1GqhPP/ASzZ8H
z/U5QnH0GHc0Vv9DuHPdoI5E+PjekN23lR4NfoCOTzl4kh73hoCEfCiwJJ9BMDL5
1InmQJvRbj9tMTYlSKYBLvdx+eNBfzVdP2LDs0vtxiJRn5GoVuLDyDMu5X9lqoq+
kCrOUpkuF3AusANUhTjq20LO+qs7XXt+07SnN2uw5YDLC+sQxvaL770eS0w8d5XM
5calvJ1n0I+zOHGWb+JTwmUpW51EriZXVmiWXtILTz+uTVokCQFa9c7VSZgaCY31
KcRInu3U4sKvlRJpDpo3Ihb/1SINOhpyax4mqMeqZh2byrmy7z6kJ+NE6BPIaM88
clb0k9r3Q7LcNlExwFuEs5WksGaSVx2gTb95leiM0kSc0oITX2eb1i7yEPAtHd6M
y+0p2LXrtl16RaVB77gTBfoFfcTMFJgupyy8pj9pFw0Ix9yj1i1LC/SRWFe0WPDU
I4HxbIyweI7aPsgvviD3pakRyudXnBVylMbNoVxCSmwJVW4NgjndMZ2SASl/Efes
y9+WV34VgyP6DzYlIIPB9Csf6rjVlJEM2I4QvgHI7CFNf3b37vzCksWQqcOoNNY7
4CkvA2SoSDk5DsDNfpbYZGZKbU6YV8FzX7gUohQOCeDgOlmaLFtvUtGhfTZ4GsVN
RNvmEOY/MM2tWAlPISWCgXvlIiiCRlTOOl0hgFdzT0vPa/xj35lDhSGGtKEUppe8
cLN5q/hAVrqNi9KBobuSpY/uC76w5y1xe/ttoXbj62NcdC43R0B8Bfmur8Zr9iwL
8LjfU9kPsXqAsWx9G88RVamQltgnb4Nxz2QtqlEHD2LX98BpfMFGGAwSizh1YTxv
EEWwm+VwfaW754cc9F0ABxaU84wuzeMRWeC+BfnTjZy3OgksdALHoqCgjeeE3JRq
ui/HrZAaZbp3yXvRwjcGNnHnp80/PcUA8eBBV/tmHDiwYQyImRXY8cGXVnYQIGwO
SeJRhnmjeQFqr231Wb33DMnuLhZgAL0J2M+ZVL8vMi6KsN9r+pfdTmjDgAC8ZKse
HPLsnlwAu+kr9NX1IY9Oc6gxcL5PmG2YO1Ojrxsh/26QYPMr9CAPW6AbLvLWLI2Y
IUFK5bUy7gnjIf9W3MiTRYBwd5RcG0Hk1NzEGd4Hb+FHaK96f1PAhJMvLZThlP5k
piqnpze/Gcks7LfYGDkLKjkwUzDfifpLi9hiMnoHpxrz3AX83bDEQBpabyP/2j8B
ADNQ9uo6cinA42rpOZvLFJkvCYbNVshuZp7tRO6JjikYeYumalBNe6opivJqJUJu
/EF2FRXQXRIscYRIy0Jg1oh0++xMg7zfhsXaMiMRd2R89nDWWzEF6G3b5AVcrMZP
LfpFwf1zRfLqWUcqqXS+L43AdDXG5YnF/BpKgGjNRvPK/wotZHAnF/z6Rl5Dlndc
kdSVAzrklmBGYx9axgcaHT02MmmhAyO1aQKIFL8xBc6s6jRnAtsj857ZwznW18u2
uZyZB+YHEcVAuF5hn5Q9EC4ZtKytuYOoOpHZXrN+o+UhBuvl87W0abhy26phj7Vh
cUrxh2MPKOM3AvUpTyrJnIqLhpBgdcSMO14f+zoPS+vhCcc/l8SWd/dw3fBRVrPD
rbQHeZ9IoV2rpFT9FaIbk+pi/yHOX7pw3eDiv91yU5D23hwt3uqiC/waS/mJEjbE
1d5sJuLJ10lsQlKMFZbytUg4OCMiJsO9tqLyYxYOwmTiriwO1cteRhQBYw5hr0Sz
iqydkIs6nvHV9rL4yEfYJXhHFjjTt0596vi9O9XPBvWHb8XrA5LInmGomMRk6G6R
DBiCA1elVPH0pwXtBKOuHfpRTyN7hLp9+rdSy4dDSdhseD+/oWM0dXHpy/QNj+cZ
zKYqhqYNnsdq/Yw/ALRuC0SZ3dhawWdP3w2GCi+YVBisdIoBMeFbiHvukNibLmfD
MgdG0sIb8j48nOOgdIlZpHS1cWSeOUx8+efNxu3bPliW4nMVkG91NUdmMn86tDno
GdRKNXBJqYFKG4NgfKXlO3I8PsjnC3jdTSOUbOhotdg8o2sx+adhu+kqA7ITuyDy
hOioEzaFHV2Mw7KODuj8qomAbAZVeGwcxyCKnZkKDi2GtdFDPQvJRa4Yb2i9u+7j
ornf+Xth9H+YoeeJbqtXYMhMq9jHTaO4VHg8gfAHxVX49eZbb1AmcdygG34OFubr
yjFGyUnavLa60ti7M54Y/mVc2RI4Ta4RvljpwDRHSbgGAC4F9lQFWahLEv9i0bSJ
eBWpPBscnb1dJvMZA2dwnHhj3lA75kpgLO46IPI8QP3beMuxR6zEGHfwHqhThnUA
k/RkdtvbLG4uvjo9gIBZRbXo40+cbY2ddOptToTGFiOAbrVfMc7CdOSAvUVgGevD
L0OHyqon8SnZnCCv53MIS5VBkG8Redvzu27d0VinxhmnUb5IMUO7adPD5TonLVsS
xUW/Jt7hwhb1jvXFamZvOYkeZEh82Dkq0mKSFbyZfmmafIVX5HhFQW8/o1KCcU4G
VEtBqy6C8g8GwUOUDZBP1HxZoA+IfN7/o5UjpUvVyJBiSoaEo7Wxs1iMAMiPHJCe
ox3yKLF78LUjTK7BvbHjn1X0/br1lwzclXytDYpM1itdBV0g2rf+zsMyx4jaWPRm
2kR4QwRSB2zGdEhWrRzfQRBwoHfWTcwE1wrlgUbJOHL+4vJbiokvvQOlsqJbPatD
K3RdabvCV+sgmFXol/iIIF5U5NStbzA+Rbgu5P5Q5bD7pYluBlGWj5Ck4TQVsK3X
bVCkGR6mC/BbpTpNVQJTQAFRZSBxvUQ6SAwzERL3/qbmqmBHoMU+oPg4ddDZwjci
TUvDp64FkX58CQW0ZZl5Vmfaxn4c8YBi2Z2lWC3KtIxLlOh1/tEAWOWWAh2irfky
MfeunZwIE1X/CtgkblhA6XCHeSF7JzUEIPNc/T2rXL2ZgA0pQPcNg86Ikv37/9KG
4HDigJfnA1Qg2/4EVqXFcEszoCj1oUR5R0CKwgWnYVwbKigvnay5jv1wvSVUcjx6
HpfspT5ZfSd/G2mNVPc5vRoFoDTWQBJ1FrzvFuWDUtmrr60SByPJBMwtA6ncXnkN
59ocXsFdOwi4oKeOVxtWTYJTT1DxdTTRdw10Yr2iHpznrXuxAGDTDPpCgzltzz6d
TbgWlkji4mY8zqTo3VsFwJwTJNlgrdH2FHlvxeF4g51rFqa8R8UPZESUAScHA0gA
wWOU79iIC6z5zojMmajuQNMI8TAMLauWV/wWPxdatwoLfCU4CN/mei4n00XaVEFi
8P+Vsus8A5xsza2TsQSafFEXusbDZkqr+JqmLJsA63GN17+MaDFhav40I9+ruGA1
N1ZO4GVEQhdOKvAllOUsTSCVwUTtEbPS/5gJR35mnXGSW//z6YLgws/K7FNqFo0L
NFjYFdo3Nj8ByM/eU0ps49hzOM+ZoFur9QUWTxoL4sk54yB7opF/G0BMNg441ihG
psaOlL+blZFb4/Y8n01H0SMCv06WQ+xtRGqsazBqbs6/uwZveVrZo2rl38pFLIOx
ppepzHFszN/1CZnfSd6wTXvHqbzyqwaAq6gAix2se4ymokfLr+xt8Ansf4ft9QkZ
kw8OU+mqA1p8YHo76ioLVnkTNrhUYiaC0g6ybazPMmkXyIb4ZEqmaSccRWbr0T+I
C/jjhPu7xUIbRBJ4IolR8cTUbu4v4A5najpFVZR9hPJzFaxBmuzkdcHb8E9zAEAs
BV5j3d4NfHcq4raoUD/hlOvsdNuYohtdL5DQTPSNOU/f/B/wzhC7kzJ0NcncKXEH
KTfNueMYbMVn9qoovCGuW1cwcOgdS9Erac4NAWjmh8sJOGLXuDEwLFe5KvpgOCTD
8FUGn8x7ITIzIMguzKkqN4UDrpC70sduhLIle1HP7hBPmU/uKHFKpvYmBDLb9ysB
epT9+OxINpzesnMJsVBnNlJS1UYbzAPlIPNWs/TrUFd9tx2n5GgStt3g03U/murU
WYKEx5Hy3sppmDQjRrnY3s5RgoW1iotxfBqKb9NtuXe08uRyHTHS6OhTTUV/8zIg
OV2kiz/LSdjgUO3J3/y0vJ4z0d6rwOYC4+SbhfpqQT4Ep1tl3TVV5P0BkFR6WxHU
fh/027RZQ/B37hWzLMhCud7V36YpzlqRCCQ+iPSxv7vPKpM/NR23X+32BAKarUQH
e+Nwpop87G84fpOe5s0lGALkOFtxbE8NReUgidjcqcbKXXkckaxxEgUlIHb+T1Am
EHu1vdXGVNdLFsqZnHxUidwJAROLG9Rk/DeWmk//9CBjXBkl6w0eAI4CR5oqyahv
Jrv+krokd1mqk9rR6YjfmywdMdkrq6Lmn+TsrPOzyIYp4OGs6geiEttBb46tuPKJ
3BtYpvHtrylgUyhI1bDRW+hRgh3PyoaVLdNYU7qwU0n90SIsxhUiFcJA8JavprJ7
KQy5tcNI/Vbe+UcIJczFYzwcM5iwkUdGRUbiEPvR5Hoe5PLtO5ce/3/mdDVoNtte
8BQPyRlA5Vl0WXAKpaMOeypR1oyMl2fzSLsxFlP0Bm4l41TGXDYucGSBh6XmdVHu
/5SQYHepWMCOkBQTjaTFTq5SwzvNKGBdkvaEEojwUa19pAMompP0bkOxDogGrvPc
n6i+s/pSYZwq2vPU5OcKEaGJjWpAXqLxyzJ4ov3hfFTNThka7srMKFt385JMJ7ca
SxGv+EBLciL5c78INEy+6OWcg4nv23Z/u3EuQRK4/Sam/IXyzCZi2G0eQ3Hw20pj
Evzfh6eV8KqZfxm7YQVR6gDiqkkHpizglrMIbciwkb8ioOqmJtlVKoRkQ0ywOiPf
hn3hMEj4z8tfsvNXEZAPt+JvSprN7YiaNUbJWsF8u7TEgcHDrdElXXiXNbq9cYLz
LomC822Id1cgGOpLLsTTf3tgfIFMwcgNo8K+lYEn4hEvGe4Vl1Ht3Nvr/+q9BJeS
nemFKqxs0Xiok1PdNmkE0oaZd6C4IIyWBSnYdVEuzb2KF9u3u8W9eQtTrqdbu3mp
GjNB3OZ5A9FpPlP8R0u0AV6ZFQQWbtaB7FgAr2O+lHO3Fb8LwxlBAuwc3wNlD+eO
ucwT2grrcmdVYeAz2YXCnQIqPMLbv9uXWZhB+8MHABdr8mCCtbr3vPAOz5uWrr+e
9WCSZiV4dAeZEe/Unt2dhVDKZhiUF9ZGRBTsOrFPTVqxZWzqS6zBVU1+8bfwn126
sPst4gAhLTedp4Oks68/H0N+j38qIEIc6wGEYigYjaR5HAvbFJDXhdYAN0W94RD2
A7kDfScQJXcCKXwL0dg2IFvUPXPhAxlt9NxTOY0b3kg/JTQnnk3az1twOLxbJM+z
epkmRv3Z2E5/pTuHecACd+gYT4tTB35aish0XbTAQuSI7J2h39Tdtv4cCYd6X9Zs
Y+nDudjLYAB0pZjlKeAATErHQale6ZiT74JjygHVpphxfomnSTXaultdNxwkL/GL
vUKdAXQTWucCszhC0y4I3FVAtUhZ2X9VgNVC8z3OqwmGU2aSN/eHA3QxGRxNizsT
0PyzuT/BGvr3MqJ4585eFOChFV6bsE2uVBDMSu4XdeaD1IV6Q2k5xbyHCu53HAbf
64sYH0Al2goxrVt36cOZsHn4y9fHKOQFbg/s6WRXtyOp8y1Y1+hYSk2M4L4y51d5
YQUHB7K9NFnov+5mfV7fNC9ENLDhygTNvsVNOppP+cpBKMm3aNrxfQrrZwLDR67w
RMhJgef0+RdpPd9m6c3ChYtsg2yEVMOvwS4XSr8VEr7CUV+ckH5PN6+WPpP2iUnI
7BQ1GlSDGzQW631WVkJai2SGZJfRmHn1LkDgvtiTTsPuXgJpZAdb8+9OTJ+cdNe8
twlKb47AubRMNFSTEfagIZEFifCukI4scooZRt/FGehG4WaeGJvKgEHgyqj2b5sM
E5+HOVlydYYkhnpQTdSOwcdtjOwyHRTT1yufbn9Lk2Ne2SeYpkIzYO+i5EXGlEEt
K6iVX3EYRcJ0jv7vIyGQjgJfR4x1VzqqAh/sNmy/1QPNyDEaNEOts6at/6KcfQK1
GjwbiMvGufSpxLQBX0EQE+acIgGAd1SNNho0+fhvavxBi7yZVpUOeN1Iuv6QdWvM
TqXrGDaiQ/n2zuBt7rjssKe8ONhZFOB9xfFNFhwIbApzOkLGI4T4gOXleuERzmJd
iFORjqt+87xtVqCivo8LXfQy45lUmvCiw4U9hVRo7fsc5oDNeMJGf8o2WhL/TjrP
NyDTHF8QAZu6DgBGVzs+9Mz1Yu+QqCayT2zVn8nTWICqj8e8zmfjmvhHOQ9qzL+6
kWLb3Er4vhtHnSFQ/S79/FE/qLcdWST6wBHrkQxkWsqNBqvexmhAIOiCOi86dqaw
Wn9WqGPqQ2m6RhCV58JM7baXzr6AoNgRGBR6viH7vkIniNxf0S6caX2Fjypcbe4v
92/J1aMFyrRQwcp+wk+6JHALjWAlqTkhak7wo5zrUn20zUgEBAuAH33gCSDd7aZo
wqivxtTl/7+DfpyQeLLz4YRqh2mEHqXuB/U3V18ycbFsjzNoMt2uPtfIMIPt9j5Q
kjaEbxXmo7vJqHO3fW7ehl6sOrMFY0PseP9HKT08oaHxBqOqaDeqUNSC33ly1PQC
5CZqJj/Cz9Ts6y/TailaCdTQmZ9G7p0vqpQw57xXfzcIUPtV30jxJHbxBtPzObAW
VtiS+XGhrKPvzBL4kCjkofzNq6nw94VhB6a3EjXiu/5ySlOWprq8RO//BwNgnJv9
ncaGBQXfUHS6sklPi2AQ9rCqOGJHozShyUol+9sK/22s2RXN9m5H0eGOeeTzTstF
rx4jVj8h4Z8/diBu9bfuEFoJ1V7oRb+mBLlcVfqHO6l8yAC7pe65EQuhVVqzp/+f
I2K6Wq2ExNPFmZ/380fedcjIOKdxWZ881rh9ceEghZr1Xi7Epcy6LZt1lLyEROyn
csNGLCiXa+jZcLdrcO2kBBqVd3SmR9slIIdpZ/1V+rD3CG/uGFxqjnKPaeWzqPG0
0JYrgtJsHbeMpyFnDKWVNgMMLQZf6MdadjlEoZjRa3C0+y+gJ+sADPYiMOnphX88
DrsgzFG36QNMeePl0KlGVaarjiJZ4eWpch4bejfRVMpN/McVzgJM4pacyYQwGMK8
umWWMoDcxTsXoN3xFFKlNxffQ42i5+5de7T/EwukMcY8+jNQMzSS3GS6E1KZbMQo
A8OWb4/Wk5xeKQwQxBvVBy6zQi39T9LSB0XCyoRudCp205afhdc/2y43fJ0Th0A7
H8sxykY82eVGmQ7M9lRxJzdrHPPyNlUYGk6lWykg3CckjOMkGvFtMPk2bqgFLrR8
mVQnxmqrrdx0F33a3V5seEm3fYgQ0Fv5IDS+Zs4bjqLhUGurG6qJew61LbbRFqCq
G1ZCIHK1t98dVeqVkW38zk1FHkwHQrHo6wjwguKnGcShk52QoknHpDV3PoB/ZFiz
GnLbTc6VgYKH84AlnYFAp7hbXC1hzj3IYkYSSXbtTehCxOXsH9SK+1+LlLCjuc7z
I9ZwQ2/zOCMGCCvLAuxVK9fyPq5s60zAZ83JDK4y1tS4YAFxX3Z8Btqet7g5cCCG
a8EAKJxS8lrA1qHl1vpgbwdAZFYAQyxYa6dPW6Wn0k12Cu2JSAiGnd9qiWec3SMo
TrOmiwuOP8+0N2qv2kJDn7mteObRxM14W3Zul/PjrMju7CLuntQFfra7UHcM21rH
HWMsEXi23PO8fClOTpxZurNvJ1bmiZuALrv99ed9xtKdFKICxGvaNP4ZC+bsXz6L
Y/0KWmEuYrBQF/NDPRZ64uQg/EJf2LAfwP3YEFWzvjvTAWTbpmpQm2MLUfZ23B/L
QEloZjvweBm1+OwHUehqf90iOuQjbktBIo2ipc9cwcvnQdewn3NgO3h2RpyQ9W9R
K5C4sTR+ceowwIDelzAGM8amqOBLzhFOjB8mmYEcUVQshla6sK0OjtLq1fS9QAz6
SH9doDpTClc2hj3c/FySiHJl26MvWV8NtOvIWsSNIVoxoge5GWuK8OOACucLmiYs
HsTRZY+apcYyChI4TfPcb5HL438b7dl4SyzfchJx9kL4QO5ghMQCeYEbhDZI1Z3f
0Fyk8WpJiZd6nMIWAEZHNamxut6fbDBlXCJ9/P6HReaVxDBK0Ojst0CxsXBAReoP
VW3uHNZV6/zDG/rhqRPsRw3++s+dqReY8izu4sbOr5sCqCfsNGQWTHItZe9I0/Sr
5kyMbHkSR26XpIDh8S7UkE16k/I0v+zqAQSLNw/LtYVyB1BoOulk7kS8rAXEpYkI
j+1ALPCrfRlzCN2fiXhO4+q1Et4EH72VS6sy0/jBHeC2nPtgQiwiOA91lhXDTWey
DFGJEMqB5DW6W2/MBVzATyB1RF27XASmlg7hHrkc0Q976uqRfP/7fwm0pR38qNN2
s8jM8C2nzQm0c51yTi2Lm5ktgLPH2Gn1ghV676AeyG5XUQ93WDhiI+x43xHSsbyK
XtgzLslSPNIqY+UgHWoUUXVyvp+thMQbZVx8QC9Nap3MfSeGX7QozU/DcHdFjcev
rZ4ZMsjMg1Ibeb7ugSrY9ApYT90I3+t6GB/lO9GYF6LwNW5yBSjATJMUzTunTh7U
m1SjLD0hWj9gxGiQ2mJkNElRK26JDX2KH53XZ4tbG2eAd0ekxFbSPNNVoCQ1+hws
IBuFeBaJwyQUZs/7yoh8MkwZjDD13FI2/1XdsEQxBykS7frf2KuqYJXeuCLMleKL
FvMXEYU+oMxDrzYUZk2aMxwn1m+uqtZXEiIGkN4qhH1C6+owsP+KE2v3T0CNhG9F
trTM5nvJAl7F2OKCBj075VF7Bb5Jc5iGYpFJciv+ZlvV5SMwOzJEOnouptCKDL1d
ZuNw/DQEE3wGX9bRpMe+gdPNjC8Rxco/zQQO1AiziGzSu41WKd9Tz83YtN7vd+dX
+nGoExpsJ49Zx8NdEqLPyBPn796e05ktJAgEx3/y5EiIb+BEsagNtDQDLuB5Ut89
pDKZ/daWdlwyWHLutdF0dkuhg9B8KIbLEn0M9/4fMISKFXkrPOs2cLgl7ThCh0FK
VLa5JKxT0Sf94trTNX38H1b8vvY1uXwxdZbmY0oC4totzFsh1KWs2XFykWvaRhjn
uTr8Xur4jd5cnKSZ1Wa62M4ikSlztE9wkyzrrYnk2eQrVuxKCwxfVa60NV4mdVYj
PIOyokbxRfJroNLpjrf22GFcfAzz5wlf58sXtiNqn+IRGf4ED5pshFpgItY3HkpV
nX6ySmNJTLLSYhtaJGaXXZ4FXPjLjhfPotu0FwaruValUxEzXJWuCSeEYT+689Be
gq1SUvmQqD+vXCWJdIJGkKWL4OcvAs2Iock5dub7ylLGproql7iNwFRMISVOIzek
KZ7KLRZSzOn8HZucTEqiy2LmfTdB8ZhN76efY/wRX1wfGzVsFoTMo4AILgQHjnIG
naK5rMJzY0o36hXCy9D3D8CXpThwtsfD/pQwhGv/2O05+Y7neDpBfjiOc1ConaHm
/nujmN4JZcgQVLaE3oNGmzWLAevDQUaRRFvkJlzXWHwyFDbPFOVdmfinaXu+gvDz
S/J3zl6B4Vl4g08AJNUa87ycmyD87+ABcERpr5T6BGwb6MS603nyXtRm1TL6v915
o/LWEuF2uQ7eSMZxnaBfgNFL3aawAQwJn9CQUVTq4yEVSvkoZBDfbhvy0Dz8TvUC
y5/4gs77AThoxYY1DJa8SJxYYiN497fkXNVEoqYeczAO/o3ESG4Wx16QLXtUHpz1
84jHdlFtK94n0LmLLZUzTzr6uqV9gXiKUWAfX0uP4wP8SiT2iz4K4ReVoQ18l2P5
xLj4RFJdxOwxjg5oxkno9EstAMBNLHb7ppGmZvvXT7CKaipt76NyUmOVwrnNTEuG
oXFURgrMMxMxQDet3xBMFcyWtm/uuSBP6zynMIwO6HT6lm3Q4F3I0BWXEUHa//NM
JXhTYZ1tOBpgw0uLdY1KAsQvcAfeySrgZ+Lfqs3idzZtjAQ6lBVP0TGHe7DotfyO
VUnXg7nK0Ns2EZTXKV5Ysa62/0H0tdoSjMc4SrDf6iu8gGnrqTAVIow9+v2PPrIR
+z3PEuTE2+2iVw/0tBYY5q34ZuK3ABaXJdgSeF9/oQvReYEjQNvu91aHfat7JTX8
Cofj6ngkB051m/fuzNvXk0WS7YQIKMr/Z9ugw9KM2BQdrXvU+64HZA4LgbPmjuCB
UNysiuQN5mExKC9f2kbc5G1dyqKXfdGlB3CMhEc8Dlch6sFKugnPF8IgqR/Mc4j7
1wkLqJ90By5AvkC4rKt2rHw/sG8a0PRhKCMGG0xjic5/wqVkQCVWQ8N+NHQjlUGB
CDJfpnmhAQC5RgndlWRMJI3ht6Wh69ELoXwAl7NMjcL5/s0L0L2AcqjWjxKqsjVC
NGeBTkE05mQqRpUEOKxxWA4DKdHh2aWPPbwe9UFEqRrAvjt7gK/axMJKTq7z/h1A
+plee3I+HmYHexPMvzQVP3nBt91LrXlvOH955LLimo6491Ro6kCW/Gmks9Bt/76I
iluVPDx0xdzWwRpkuFDLIXYKjE1b0uwbiXx47e8egCgwRLXDHI06O0DjMXQUGAQ5
k1v8peVOtpmq7vo7xLcc5/BNxOQYl4x89zfiYFYgJ3E0lU12x8uFc9MCvh+5k9cl
UCj3DP3eOC025dQY4TYu096L6d810t3EVq4TOxEJCpCTLSGJOU3JNzmvnYgmC3p3
kMCXKwWqugUzc3ef/z3mTRs9PoriTjkhGueZDsrICJqwt5mMnyy6cQzhROnn5Rbl
GdWeCGaV7I3EJFs9LeO2oYPZLyvRvGsImUzamhUbn88uGptxy5/SpCx7QX8fe/am
QHFuvAeM8F07CrUEjNAak35J4vBsunGmTOOTCeFCTwWtEuH3La5eE92VzBPThK3w
qaJUvT/0VORXmYZ6bQFQdGofGqSLmQCd7qDNaA1ZSkPtTpzq4nS/wSCw/W8JDicM
/v2tTsfGLWML2gk2JJ1qcFMQvrcYVysMFgdnD1wtaUlc8hZaY40MtpS9m8+ulH/k
JxSFueDAesITtsVrH3hVsLjRyUoarVXuDg7aTldz2M6FQj5LnzxvbplE0610t8nR
YRQQAouq51ZH/nhESGWBYdvM6de5vFSzDZE+3WqNXm897joKOgqJJ4GWJNLMti3M
x9nA8X6NEpcG/BaUPZDrYp87PJxJGbqVpSOvA73XRZKqjjJGE1xzWeoA6jwsLULZ
yB/wzZCMokB4onh7y9pCcGLNd/mnKvV3xwGDS+HFNR6mIbHterbqz5K0eKIa1ShH
uGzpquTQdP7VqFHdgTV2QEnYuTmJr+BzEonANcGAPqgdBeMF/ZgaF+tzkmExQUst
C9Dns6Etr6bF+h8dzavX8EUNpMXzDtZcjtXD4NDqiNO016UWHyVTEw0zrT1fwU2R
D0nOeRYtqHoeT89ZWVwcj6r67CBDKaUb4s9JMkpS4R6/G7CA47Wdi9xLwlRi8IlB
QRNXOy6uDWn+1AgxEaZjOKL0Sc0DccZKD/BfMwYIRd3TFIC0p3/m8RCeJ0zmSXF/
lgPKN/aibX38JXYJu9qnvCpU7ek3XlPKJ9f/oF1iTfVz8ABRf3ArADGogD+foDAw
ZbY7hP5TB8LJ4ADiq+iQVdwsSKX4kPmnb11HLZyE+tQR/8oriJKGQBy34k5jnnOI
Na3C84/jEvtCBPrGjh/KPfEXAGZjnfKWBdN5rHwNmivBbKIP9X839BXzjA9IU7Rn
jrmlnlnfQ3B7BgYjHJdICR2adzt9aSZdj9rGo7Qg+7bxVYQ8J/aCMFMUe1G+LRm5
OuYoHfFHVxgttqT/+mEqWHuUyVi/zuJTiFrwrp9SLRqe/owRWDVqdEyeVNnxkbNZ
s2nMis3128TkLAON2/rwYGsW1+DlAceYXJkstJ4i6vlDEy5TMqw8QwatgeS02pDz
cisINLWI+nN/059C3IVPRW/Z91kjp4y2d8Hq3BGsE07kjVmnzFC8wvxa6MtaYfpP
4P2UbubeCXupcY59uuV7TxWtIaUVY2qspFnhsBp/jHyKqBAkSPxLc0gUXU0qrnO3
f6nBLXCM9nvxCxKqWHmlyMiU4/hfNSqNg6Z3b1A0VFCfThX8vSt83RllWXnPZH2/
EfqqotpEwkKqLrG9XtYRfZmSRdBxzEjm5wr0K+yzvtXJh4J4G81luenwTEMNGYBC
C0kOa2YorrzA942bVHO8JF+hWN88fP7T3GfYBgsfIA2xazKlPPbnzXdxo3StG7he
La1YlSg172Gz4xlbgXb6PmmdmGaEtrmYxPgC4Tho/zONc6zu07mT2vhfjT3lVxxk
34AcmYLJ5XaU1PW2PammkaI8bZXbRY4rtVWa9FG6pVnIqyyF9UqSnB4Ra3LZdt5t
qX7IaVRgq7UNbjxCVFDxJR6Z2r/B6MyEbDQODBDwiRVN6ZVc5LV9dMItfJIbSTbF
fUayuKx/ksAMB/qWN2xwohhP8ESFz2cplfCuGRXyKLnJ6gKgo6rvh2qUO3dmIq/N
fLpiyWioGfzisPUUpyidrzgJU9CopfExjOebTjJAEOFqDdbiUeLKOoZiNiHEx9GR
rKH9eNX0rDUeqg+5rU0G6w9Inw/MMaoz1tZYctzw3DAUi8fciTxYoKfSLIM+xyuf
ftDiiDijxlUv+AQeLXoC//Tf70FPYU2EhJ/MeJCLY5SksYyie/Eoouw2teYkn0+1
5wssELx/Kg+te+njn58a1JgkqUshexxEPifEL9jswiVbxow7a/TbSR2LKYMMVpKe
rDnAYra5pe964jmALHMBUSO6ZEabRgnV+N64DnsVAbIkyGTU4KzyWgmBIzeBMopA
vvb0An8s0jQLbbhCZNhlw5uU16oYL46AwJhrPbc55cPZz3IflxQXorL5vNQ6rNzf
pG+tKtYKer4EeNGQCuVhLG0PJ3l4vjxthxJNSKJV9pTcNAsvELh6y5/zAM6+Mmdb
dBX/8pfYQxUfKNMDZ/cFylJV7wfJaIi7KK8BRDH1LAtzU9EzYLyaye3whXELc6nq
B+yfCThlQH7dRbdVsYKxx6HKgcm0rwqUPD+G7SEmTNak4UBt+95HjbQVOGHz9jJ0
UjdD0/G1JUfKKEp5d5ASXJkb969QrBXsnT4LWgOg5AofziniPfLHCPTfEFHpwZkM
TuK5PStYzpLKdHkOOw7VcQScrEuzgTxfafy3EK0r1ahR+gvB/OnaQFx1aa15diV5
yoFrxumTgSsaMnKQ4o3kmJEac2ok9G1jUsCMcEK4RXT5PM+c30oVyo8kLk4DBM9z
WgfanUH16k4HhZkokqcKJG4wP878KSgMGnz6BNO3Q/1mMfXHp95QqZqZ0XogbFLw
YHEeeazj2X1aBajYz48+XHByIwdVZgocRNyeaPYUlFcO9MVY/GH3PIpfZ/cEgVf/
9UZ5mlO4ySYnVH1kNhwxD02UAn9Qv/0YXAYRuQQ0XOn7v0eQsQ5oVwK+PbkUXCMZ
HB1qmIqx5KHAePLEMlKrQcppV/tXz368UcadBuptYyYfGf98bd+3pKkL14lHjgOW
dO4fMisjhHps5mib0yjlnYX/XKTv0RKRljr/E/M8m8obMt+Pxdp4dZVoS5sPSoBD
qghFbGjDrF7SEptSWnuaPQwS2Mwx4qQo9IGtJJ40/n614ftPa6HNlAbRTIDAmMzp
6KJkbAA36oOINid45MtlxISWGuMwfhhujmsBy4XYB6PMNYGOi9cRz7tqpfm0W0qx
EdUZ9Diju2dFK2iE+hVBCteX/u8sKdIZqHcS8cr48HnzszETtHia5Zvl55H7U8BC
AjQBO3r3jLpSNaElSkrPNHLNRRvxmbom2alR59y8a+Hu8Avb47FHiD99f2LFtzXn
b/LNFcAMGD4Db4COZsRkTphNjXzSLY7fvwciJWKEoD8I9CSkwXcf8IIbdvTkHpuZ
3Qggh0Ss3TXIK6LkNtKE5ipPiiNtpUDpnfAebPM2V7hY2inc2pP1JpjgiwD0aFRT
KeLBisBIsjXsMfmjYqb8c1wArUthYk/GyYtRBZoFILlWu7hpfVaapqgKtn8jcGid
J2zE+z1j59SHfszc6uJhMqTXSjZateyqZLH0nlXzeF7yBvWDB8hrj1mV6njcv3fp
0CoboU94fzP6Tkb0ofGbTrDw8FeGrVvZVLDUCSVWer1/WQn1qvSqAG4obLstfc5L
/vh/wCgw229sivdNL24TMzmkkrSExBirIdOKGFbHBXQR2rSdT+0v8xY5BReFu1et
ZhmclHNxdCZ+4sjbfDNjkcy55g7PT40i2tafVCc4cTNXPE8W0ELlv/FDMWkrlXzI
2Vlod2MWmHlotfopohLyAJecgusSmxK/Nxa3bQMHPHIqTUX6A8PHRw2L+31oq5Jo
csTyjwG5g2oCIwkr5I9CUnHEsk6Ze15Ox8XcjyGBTP8YhTKrtv/p+cmSsZSgspVQ
C1lIT+JXfP/8RJMX0fX20dXYHKm0qVxD37me7XY/tFe0UasmuRpn6VVPmEbghbhQ
YkUb2ib0Fha5Yr0XIAMJHxiZyeqpeD1tC9eonpROv7uDsedb3kl3hCRF9fC59m2J
uQRuSYshoCoZ3qj7gc20PuZGWtRfgvh1SoqndvmIfom/uKSiu3J1vpWNXtp8lUw1
/bOpCljOzMT7oLTmNP+XdYdYcZpG56uvi+auxQ9dyHE4UZKurKsUYYenO4HI2W7c
tOBKG0R9VH18ol8h0JEcVbrl5YtI9ivUUJpllx9M+lLwcV4HGVlNYenEJ/KKF7cK
IwYQUu1vuY46FzOMGuN8iXQta8AaeO7WfI2T9/tZt0gcIxxrA7TAhkUMydLAJU/h
3CIVg/MbghsIPRIjBvh8tzIJS2lhj/WKDUpDYPXQowKqYVSTAGZul9AXfNInBGGr
Y0eNwkQxT4Ey2HJtCgk0XsW6s6h0Mg1wA4aaziiX8X4XHuNOhe0zJklfgDxhHG67
5BPvbUCKqX0TEh/wrZzxmsKvwE79HFEVnwZ3RKJlVJ8sc9WwFtI3Y4Lfn+NKKBKT
sZLs6Co/fwUeXCyinOVhTRBVFIkySUKfbD1M3EcqqXdrtu86vgO1nG5E4qWT69r3
xJrW3/bkG7kU8raXamQs5s9ft3ewD0JM26j36t0M51tE3J4Zpxf+ftvqioqmdlmq
XHn0cQbL9FFjOGi8w7qkzmy3cq45PfC3XdWJNrteQA9g9G8cSxk3tpOqr3+UzipB
AaBbIU1/NfT3VD/Ag/OkbrUSGNxrcOMwd32mHwsejX/1I6Fy5i4BxtjQi8O5RUz1
viwD+rKspGRiUSDKHhn988mVbCVBEu+QoRYrutFt00XJ1SBc1P0j0b2LpFvPgWtK
ySJ5CGspDrC7O7ycplo6VRA8wEkRvaCnKnWJAK0AlbneIa/mbFWi03/+NTeH+hhs
qpvk0VagP+90ruZmaSutGfr8xLhsQZEVO/JA7FZuiW4vE8j53EYhUrxiO0wbAP/i
XnFyanVU+HU3KLHpZgufhoJ5nk0FBHI0cYv6Dz5C7MscHovSQ3Q50aIbyfzW3DHy
ens94euRyXLlhF4VnOCQ0PdNjMUofsTOKRSyxwEV4KrS/h7zrNxFFgTBNGfWtLJp
Ag1cQs83zQKMIl9vQuCgge4MZEjeyYPmlMuxr+G+5Bx6xdanNbDQrZNC5qoB8uRT
hmd2UKSHDPN3T6ASDa4EkNc7tkgNuz4zebaBzqN8x/TTyl/DWnEvTUVYuteP0MIA
Em27sUYCQ+HY4IQCM+YzGqA9jKG7PtxU0799NOMihLTxha3aY45Ks9nVSnURbeTi
rDnqI/aay6b9Kcq/4cc1wgk0Dk/tC1NIBFuCS2AnNn+G/AQj+fF81yCdzerYClrL
Mek5oStNXAye4pevfXYcjqAx0QC9XFrwJDqmrW2yDbXpxIy9oQu0CRccoxk+ry8Q
Z2lZ/kGkLPzHdAhyCfKUlm25ZnA+45aOHt1BMjxGSrNbBEnIFOVY1288R825VjJg
FaZL8khqips5vh/np0YU7jk5gqWo8olQ8mytripNSOaB7mNmFqazkW14aI7G8URC
aEgEm2UHKp0kdHxYRQiTOhLmk91Y5K9MBKE9vkCpF53KCr3dKSoLotJSH9bd17e0
TBbNJ6jWy2bxHhliEG2F+4ZxjWM4jLhAaHMSBm5tk2lF9dnhmf8/QpP9vVimCX65
M29o3NuB7Cd7Dwlz0C9qk8Pdyf9MKfVCX+wvKCC2FP3kj9RG5Z/7EDtrnyX10g6X
9fIi056SieGiFPuW9wl+FdGIVz3Wf3p7FzoBa4CBxXHWxBiIE1DPR5mAf+PxJdfb
C6GkwgAagJTgXttosJvxyuLKozPGHw54k8FiGvuPEcGMR/8mPA2fmTTbzzPHiC6H
YbWJ940fpAm6o4wNs3IvDyDHx8MTINVTiZOEr3tguSqnVD92yGeYI5OMSt0uCriU
+2rt8HGRAuRUpYW2qbBiJymfg7QTD6NzcT419eSvLi0adjszuJbJc82FL1C/qJKL
ITMGq5sV3BWtknUseCPCACsRMMijPGy3zgWXrHTHb4432vBlF6EYCpZEybKI0snQ
sdNHNY5KdmW7oI8XGGvj/S7xf1raYUWRG7YR7cYmfaY5AtWjSn2njYdv/IuFxTYK
DkhPavQSvenJLhTe5wSjrLXKJD3i3R9faMU4114GA9UyVjjI9sapYn8t6GyG9vUO
exzY+QJD1i86BEDZ7xDU6BoryVPnMspLhtNU1cCpugD8XfvfmfSucqG79AAVT10e
LkAEb0hUbMa7Mmwe5aKuqH4sDgpY+VKquRrNuq7j1XBPDuy/tfAq47yT3VXj3iRw
hh9p5EpYATV5KiRil784RioKdgT/n5Bx9uMGvTieEp34EgfvuLogNnOCeQmBXhfX
hqalOHksrUoLaM56Alrz7P97+9aPXzlCj376fM4tHqpfgMMkvjj6SNVPGWMNYg4r
AkAsoffwB7gvvWY056pH1mD5bhpdIaBT9Bl20XkwqfBy8BIsOvxHlbrub/rD/neF
ZqTXt31IgkA6s3oR+vyKFurVUvMQC0Kd+S1UUYVMfc/sbc53GXCNyRLNuW8TeorA
lKa34BQPe5TOga+HEJGhJc/oRPBimcR+gyuoQltKGzUeSLfy3G+IEMBfpNyB/264
gRZoDHL6z8zFOq6zr+UjATEv/rCtgz06KKjh3v1CNHA2yshnP+MLtmduJBbnio7f
Bo7a2uPjLFn3/TbipQeJnU02hYSOhIrJBVmhf1N0FWhhUGlcpAEltq+UEN33NJys
cnwB9R3p9PTjiddSalJlRw3GTVjIbBvSxZjDgb26esEqAqsiEQ0N3c92wcbTQ3Zp
cBEUjDESeTuow6iF48H9543R5BvFv3rsVFrqpYdywYjsh/lNeE/eK1K2Fz4U65Zi
qq/pj3sXc5SD/l16E6Cd51482uaMYDH0U3mY4RByGWboZK6xinwthGlzmj9WfVqx
lZ0yiPgufV1Fd6NRGWHv1c6XWGt0t1gZGJf+KjAIfO+K56E8TXsO3mW5nCY9Xu9F
ruYmDCu0wtEs3TH9vUKh2V6SOkcTodLw8kBYisNTArUnkTxilNiHGoyYFu7u/4lA
+xzivfYjh7EmYOL9N1CUJYkt6vKvysiY9D0gbNQo45Y9FRuZtb1DGTAt0UYSv1rQ
sfsAz3v51jTzxH8qGDX7wXNOVvOn8rNuhJAODQ5CzhVmNRiJvCrpKjddt+9Z25YK
BZHbG1/MMGI5ZMti8hlHKDW6bPOTKELc+SzpXle/ftIgLitnXqnmUSbQYJIbyfGE
QTbHyXhEGWEx73DR484+30OejtmTnwk/8zt+5RYhrFx5Z08FH37xRheP8gbTeQZ8
8dwBNeXZ6G7bQEZ90eHXMZoLBmo7ETsFqLLcHnYuqLVhY7WVETHGcthZ+dW0mQFA
5O1SokUpW0LKlJPALoFtkreVd5JhADJN1tH8803zcZnuoKd8QkkhQ7BXI5GiLiK3
qxYS/pajbd/pU2QtovqYbjGLUGjoOkZODcAfRuwlyCQrwsa4J7wOT8s3kBa25LGp
1oTi1/Mw9lVa69bcB3AWL6Lycn1u6w8JTZ0wCL1pBDLLcCun4Ju0ImjAR/fVB36P
52KpcKm6EiYrFjLYBENH+ESG6WuKWYYpZnEVw072GLysh0T1Xh82Sqe3m/TWPE3f
wmZ1PsKK69Vt3mObYJhvpmiQYDbI73aNtpN7YabWSegAwADJ9wjbhf1XUcWRN/DN
8ge7QcHSqiDlWUN4CJmqSlBx30yGXiBMcLYYFD3+xA+QL5rACipYqxk+rZxDKmjs
T8ACu+VdrSr5S6N381RBJOHSIn90HkLrC0SU07Jot2IyPZe8fiThghjvzFQ3xhGa
X60jOMKzaAz4GVRZFjhSeARIuLYJzoETYc+FLs0UOVRmzC+XwL4R+hmaUH+c/JO4
bzu4VGGfPEPFKElF5qpFPEicH8l2whApuxNSoXCrfeaQu3eK+4hSE4fPuSrtkhzx
0QRTBz0OCf03d029YJULNdFQ8D3zys4bN+nPIX5WXioeAPLaTclOdChY9mqq2Ili
T/hNbLv90e5D9CoejzmBAQ8Ftmo+wrspv7vtCpikDgNW5XNASvd7ZnjVVfyH4sO8
+fWv/E5ECy39gN7b+CQOggkzYGlpK3yxrByTAKArQe47vET/Qm+5JgCJnZb7Exv8
F9nLdlEzxZ05O4MZjAjjCriSnVHhnkUMxbD99ZCpRMkcw3a/gdnib2oGotQrkYkx
UU1GEv12MAS6pZB7w6sEKRy2fVZDkR9JiMEiEloMIuA/vtj7XI+x18T+GTqHhB4x
K7ja6pCl+A/MCu922+53vrdAonBsU0Mv98a4PyAjLAPnWzmBw4yx0SnJIHlF8iRJ
XiMHqSzxZf8qORWQTee6Oj3aMajiCQoKV/JnbLs0r01DFPSDifilIbEpXYqLcRe4
XfPEn9m8+xiOIDfV+ImCzC8pR5iXNixZ51ZfKqFUYcD+X/SlQEM3lsoH7t1XWo0R
fY/A0GM1KetcmQNCNtBPle3fMvKqcspz0oJHgcFumedp2/THNfbxCmQs7AI4dRnR
vrqH8cwoM56+PlFE3vUJLR4iG8+jMnjHQZsKULCiIJjp0eC6vdwevQVizGDf3XTC
gq6wOoLlm9Z5zp7rf3GTIQDPtlVU7VczQJ5Um93fJGZIGYt4GUyEDp2FM8Ctq+sI
3LR3NPgKL/ryhj3xrQDeAOvo9qFEUYD6RlXtzu93UJr+RNC1qOsQ4NFlLODuQCkJ
mum9Ifjnvrcgx9NJ7BbksbOwJmDDCC8DWfXjqSUfXm7loaNIUV+RRiZKFWmgVf7c
NAefv744rERDJ5GNciB45kCN7ZKRVWb5pGOR/GQiMAhbZnPP6TwruSZFZ/twOygo
UY4gl611u1Af4HaFX3lk5T6Rc8wP7RIC1rRMvEojmtNvZHt242vRvqwPsq2sixbA
scAjJitGt7upGL7SC3Ygp8ncC6PZIdBmmKI/NK0MDw32GiJ/sRQBrIEK3fgvMEa+
/dl3eRbjK4sV04GJIyZqIsCRNLPw8dcwFeiz4Crxz3S15A1CkDt3iSB4Y2HS6gTC
z2pHzF2yOFy44X8WYjECe1avcB9xQNXLoyrxPpixDytsOgI31jr5JuZZzMuVyzMK
zOJXmC/2JKD0YrHO8Y4iAWm0iHGlAEn2VppS+yvT1xfIul1wC30xsiRJSaYbTA+/
2DBgkxuV3s138o4riCCtR5cgTcW2Hj6xnPnTxNOnIyd4rZ4Gmvnmg2rzQmUgEhsp
6n6w9Bpxx/rX8KqudwCNPIEg/fSUulLaqhQtUcE60aKR2qLda5kOsSsWhGVoOYZG
/Pknsu4NmMQNXFprLOEzLB65rjFmDg2OAjE8Fr0F9qTtVEbJ7grg377pCE14pe6b
a70DXS7YVcUuG4Ss/KQ0ZWx3kI8gOI/huVLw5PSlACKHFzlvHGuJQF2sXjorN0EV
jNfh++Wkv8oTJMNnAhrAnpGGCJpl7sKmRZ1kQ261fXh6fuyZJ9ox1lvgmHF/tYM/
RdWvkg7PLP/vqkI8dTnNJq7pL3GRPqsUCA7kO7qzvvHexVaX9EqsRgPJUmtOa5Bf
tUVXJflrv5ujQr8MpkFGIxxnmp9QquHBD6xhL8fUczwKb/Mo/zfgrx95Z7I6dQSJ
AMosX3CbXRnaAbEZLeqofZZb9itfx32sFG/hGiiGPQ7cQRHSc/bGCUeU1XxSlmPJ
0rq0yWB0klpktkLGtXolHKrrwQ0HzIOZqJRWnsicPBRuFSdJ1m/SJqjWA9KNGk95
KNWQ/jQGvvss0u0tq7ThfYO6qiuSUthwXVtSeUy16za0FA2vJVbcMPmUvDNe6Acq
xGlTNpgHqUTHnOpfoi70IdNg0pysAyn+MIYfIuYIZVN6C+XViUVCJaQVx6AE0uzw
W0HESo15IXSqhgfqTJriin2ezsKhtJA0P5s8cebibCrIvtwiv6AgOX18hJ3LG/jb
dzyss4wt6qsq9eNL6aFxaX1Attl3GpluirIf2TcaYOam/qr00y0sIoKfY4POf8gx
TWKV2EJymu58+u2LLlOohbZ5vW461YXPsk/oIivR7mipSeVQqdSTvjX8xsd2yGRz
BkTlu0wJkMfmSvW0s9/9nJ+O0tp2kETPphV015gGeUW2evuFRYpW9yh4b8xM1q11
ujv03Y5L5fwRsXWf5x5/YHo8MRQKO5n7+tGVAJJmt4jnzjavb4klKyQIuigW/6xG
f9VhXQc7LHejvvQm54ESjNLIMMj/FmQ6Eng9ut4KADo9s+sDj73Web9UIXAMa5HX
OPQwj3CRTtPvwhjbo9e1KfPIR32OL0S3/cFyclcVX4y5ttxljqlKoNPOhI/t+SRd
AEibtjR76Y0lnpHnwTqEW0XrPFYz35c9si9w2WAOri5z0iHJLcmialrlYP5/yGUp
n4aQIWjkE18y21U4q+JVJxRxIHqm/O1z1K3/u9tZtMBTY1cR1F1XytvscOKfKWDf
vcGg9INvxYHz/LHFB3g7mRBgHezCcFlyVI1sF3r7E/+06ORVEf4yx4+diF5sMTjK
7uzvSRMWRjnEPd8sD28Y5ZnMz4Rpw2PwowMUqDmZzvNYyYxlPVRfmT4/5kG50wW0
MxkaGOux+a599dShnRGhv0X+ZSFYdMxZwXvaKngDOdaimhtxx/c7J0O4QUheEQat
w2PD1efkeFt01+yjoAxucsv/jndKqREsWgNBCtHbT/k1+ISlsQfb6NzS1263MISx
fXFUCUm/PFSJ9iDPlGOLtwtaE22SvcTaeLtGc8cTMsSCcn8JPGaTeB1htpxJf7zG
KUBY0tXEvqMa76mdtl/z1V4zE13/QhsqolNUBQUXEw9TkPz4xF2+P6DbFZoc0SUS
99Xm+TZlp9bmFybEwRaCyJjSHzBia2OUmfudujNL3kvfjCBnabDVnmrIlDnHY0SD
xr2QpQWO0jMVWdTZAeJUMuUWW8xmBnTwhVaW8B7MxYonVhnQFpNAgcPtekQsNeDU
pyCsFfPc7PFq/muMvQjSL0ruJUFbOV8IhoQJDNJFTrl9Jq+s/zb9IzyAZAzWJYn0
i642I3RCDy1Qf/JXEgPp6aN7Sv6+fBmLlKYXv32R2DLhJPS01U7W4C4AcfaSTakD
hS/DRH7hlnG1C52F4q8S29ENqFB2p864VOQAGT3tpocZwwlQ/eH3B6k5xTCWFFdh
2ol+tRAMaUqXN2ojalx+zo7Z24h/zV+XRZD0wqeKNERoW7CVHafdqETNYlj6KY4M
VNNntAigi0IcOtgkja6yYKI41CPWvvIZLS3e4wEHBsTKu1AjWDVRJmDI4D4GRB+6
heqiCG4E0YJ9vVPoKmtDAjJC5cV4mbmv1XRLHFaLn2SOSmzSlcfBzMNY4eiArw+G
ouYxuO857vBmgshU9RkEljRvLhZlbxV5H2iIFyylHoQC3DpwmAilej162QjKf8yw
Dc4GFWA0za0pxf3kaMS+s6EVHAI9zPXL9JKhD8dCVSZ8PAef2to3knRW0YMfGw/X
Advoj4nfRwZPgVhJ5Llxn3MwVlFKW+AaiXu42Vf9GKF3GP2solqdjRQiOZjSnf3a
e43bTGt4Rlgh9opQ5CB6kpiKPFObl/zKZEopbGU+cFQrXI9kLOprFqv1qwOlWKdL
fi8KgGtehb0whWXVyCC5Veg/oHinFv/uVj7N4RZsbI+thf1ptaGNI+B1fdmr4XRw
ktjLVOX4ZP60ViJBbK9WQDdV6gV7+MTTdakszx1QOOFwXID9cw7bJwNHqyYQ6hmP
Hq8ORTqlvlLy8mjq3fIgm5rtE5Eq6+oVIANMLxr99/p1KMLZT1Gi3YmJkkCu9EvV
OJAwpjAA448s8Lh7DCWwXpy6N7IWh+H40OQvZhh5FomTWcKZL2Ht50Xm2GOES4GA
6EI2UGwJ4c/ndLNTVmHKGhUJsmdVact7JVburPz79k7ne4iKnRq2LBpFlkHpxDHU
47qCBhWvtP8ZjGCQmDI+DlbUdpdGGH4EKsNovn4ljZwpZWLhQOUR4MSKv8NeUp0u
1WM3sUxSDHGbcjaNVw7d8dSSrVWNIgFkbekKojoaMBt48qYNU3LsLI44fTLC8e1B
frXEGZn1uNRDkXIYfbcVk5fjOZIWO1H+I8EUqIb7/7kBSy7d601WxtLQnAjrFzG6
REqDRxbRF9ILeiXx9i0pE9wyJyw55H3EW1SaXPXEHmfYQSXVNYnwHBRWFOh2lduk
/ui++5GIkOkjUi6pem/Wf/6F3c23/5KHheD/ey1nvrzZVaEgnfpHz/IF2CaJRvaR
F5L4pb4EcoLosr4fKn4CQyN93ogrJAHCGE7DCCdPBEALTuTT9rTiC5HEecir+Z3R
U4lMhcXOaJMG3X5rtpWBPUq9Houp5B8nlNzg/aWD4xE+wjNjFZ14D9oMYUG17Qbi
7OTJCt1TgoEdCmtPVHqaON3pihfynCmpfIRRWEsV1v/895IpSR4xEuHcR6Cl3016
PHRGNFWgp3wLAiNIVpZIvA5UjvOdLNfhL7qf7UaHaCUeQCIhgC1GkCPac0+q70QS
+48wdRmU+XlKhe6qax6nkPqQMcGYujGpdA9JesYshpYGZv/rZzYBvdlu8uWRWeJp
tGJ1NhWwgaSNbOQzaHqSuoZlqNtgRJpK7C9NyMaFile4REY+S1BBi5BEOeOwuSB0
OwzZn9aPPDHx2CGPNH7ESONKc6d5LjoYV8+UfVzlkvYUUdv+4ptXpceoLvyMV3dC
GQiOAtrFU7QeKYjGHqZ5kgWaUsJ2oNRMk94lww3yWb+zSjp9D1YItwUyIxaVDxSH
XCVgG4C334rdkY2iTI7DnA8wn8ctqDjDbO/9L3Q7U5hDUqgsrptOC85cD+fHbR9a
CZEhwRNnS9l1lJUj41r/sYbTEb1+5kUA6vlzYR/zlTQPhtIcHYHzwAuZs74Q1U5G
tilhPY7WWM+tgj3zfl65rN3hxUChXm9hf2byumzJA9qLo5PXRPkwxA+QERJiXVJZ
g4hnvhR7xXBzVTTZc+7adoQC0h7pCGBF2cCjv1sOUjH67Z6MEjl4Khlw0e2O0Lmn
YuRgESa94DmU4hzidZ5E0GkEZ/p8LbtWCPz/17vq9RaH9ajQ+AZBay009lJ+ftyb
A84UBuJv+9vHOEVB/OBmGULfXWc3w8dDzHETCnuluTWqK3K4WSxmbz54x8sT/EM7
JT+pfi+5CcmZ/4oK6nupjgL2REs97sVdpZa6hfyaXGKSWOoxOBRGbE5+4tUk7Qbh
dqIPUCE8Vclf7SKFOfBL/Fe0hnHgzYfHDMuGNo0uEVe+bgLjmr2i7aBGQE26XUbI
dWQ14RYHi2WB1zp0PQnqhKXCCXF3af3QqlETy0d6j33ACI1Da8AxJ+RBrJ4J2wSh
uLp/epcBMEtpHX6OgbMe/SSnxmf19H1djnaek4Wq2hLhSP1ihPXxVeCQWJCM/N0F
Bm3xZQdxpcKqPtD42ntApEenXxGLPfEawudjCab3TZVzDOz+wkrT1lg6LYw7mp2w
2C14O77IDNY0h0wJga+XsQTTBIHJWipYsoFKn+y7E7pASsfAzY9aFvbmyRTagXNE
WIqe3eE2UIex0sRL4+rdHH/+TwyJ/UcRFaPTvOURZ4Vam1QeqpubYFhVXSXGz+Z/
DefOZAIv4CLsGrd/t1Za5dx+EMf9SExr7hJY1xyZ2yHglXaKG4o03MIYgPw8fXJe
dJyw+GOeqqdOU1YwrhypfHLu1FbS6w73o1hMXYeL2JVIvFe027GelutFrj0xfsi2
ao+MGouQQ9vul+GDak33qsR4UG15G0XyKVzorOelgqmTFQ1vBkEsBZ0B1EjmFt5Y
k1VJsSY1EcdU6kgY2qhkRr4HBqacWq921I+mS2AtHlSxvdFH3yL18Mgeg3nREPRa
eMP4nv4U58vA9TwXha24AoVrSg2Vwlooiis2z6LDfwEN9nd/ZE1JA55hE4u5JJlc
K7unygIKr+I9x9W1Md08RzvGwbqe9JTvd1TOSSD60gFkX8Z4KTY/dOXvAy44ydgV
XRP2B9cZw/0vCzvP1VIf0UXd2t2Td7RIloOyis1XHE12KFEcTdMZrVpUi/eHjhPO
nXdqPZHDnU+bvu329I8/aEPKDhWc94Xplm5eerDXLIMz1VLjNxjhRBFz+rUZJtwu
JVCwRqu3SyTYQrJE+I5upbWYvUbIfGnVoWmUqtckAYuEGqkJoikpjvbMKpLsG5R9
K3MD4/zEQiYOLnWZdVktQcq2+ZEzFj7mOWmCcU2K0/6lWRXxDebylfhpXOItOafy
Ransj3mr3tacKI9PCZ93fyWqxFFRXhCaSrBRzWrbHue/ufvo5YNydD/bWawStT82
/qZ0UEHwp2Z0lFciqsduwr24JopKsYOPIW9/rItz/Ny30CH0iL/55X3C++b37ZEf
pkpgiUgjQQnYJ316xKIXYMzQeWsMPvij4GqosNo3G3ddrVtlLRk65u7f9rU1F+0B
bQHaZ0SQthtyD8uifH35DxjaFOEj8EcVpymdtusIF3QNy9hUhN6Ore4AYVlwrIGf
OQ67viwixvoi4TO67z1CXmP4bymclyzsjXznHpxo60Vil8jZ2wXzRcTurQ2Bktfy
6viRNLATUio3FogWCSe5wfCvPZGwj7MDUYtMXd4mszBsjCPGv/N/eWgpJRMpK6OJ
6jrHcxGHVC/VEl/EUqyJjpRF+LkuBmUr4/XoLshINMzrW4y6i5W3tGjGjYxySPoA
0frspu64c2eplFmUAURJwb4nDVibEqjwqf2iVgui8de5Cew6RGUxKnuMVPRxY0oq
8On2TjD1E924L6u7lgod1UeTWCc0Pr5tGcLqIDBklww+z7xGP7+ByKyn5xXXzEvU
xk8ZjecuC18H7DybOnkfykEQSxugXgMM3DtE+a/Mn4U3acmpG8IujFRC0KxT1xyf
Rc7pKstDywLS8KEmUZlGVsmOL+3abBJnwK71onATpj4li6yBVXxI5ieun6XIEGuE
bLnJ+Y/5/wV2hq1ftDENvaXwZJTykbkelEg+Cy4g9YjHBJdl2/w7VwQUpfTioP8H
Zp+Jwg+N9i3xHZP62robqD1P3Elu9hbsAkdtooVR1RmBDMnuJXqni/IAsgKTRDWE
kYoScY62dwSeMqXcEkm6uJo8EvkluH9SKga91P3xHnSBiwWnZrWxGrlrzZtdkx2J
6mGR5dWTnmy81YW83w01MCecjoyVUWK4v7yedRD3dE9d70zGT7UOURkBvChzrjnC
Fl8VWw+5Eg0hezWWPmg45luClt57xssGGXGdrxiX/YOiuglKhe107Y05ieGtqRSG
iFKxs0DKs2aBKdCKKnmvwovuvQ6Oe3QiEUjLE3TeGN9dXD+1HH6l9B2jOewE2vpk
y9374+5cUElDs4Ph633sc3LdGkI3LAkg7lfiStsyuol7iG7/UAtTqeGv0Zft/F6F
K5KX86VvDJNuLBZlGKb8dpTf8ccDjf8niu19MSL0xPvmjc+lzMpr78C8JBnb1ggv
ICIwowpDcj3r696XVsORAYIQ84KV8nIO+yp3NGCGBT2AIyNSYzN62U/VLN5Dcc4l
2y+exdHy0gCnO3UqHReAbdPCXf9qlh3LWGhlXEY4uD/sdOgKXRxIteIXbhDHFjU9
ydlB8R16kRvtPRHfe6DGlgbpy/YuDkWiVkWC0PcuFjxcn7TSelOc9FxUtk+Xg2y1
1B9nn7W3h+kZlgyDKqk0W25ozV1WtAMtyH2StMa38X+UUXlxhQcai9ha0/Iqnqak
XCv/3mNc9Y2nOKfJF4mNl4rn4DxL0b9YZJo1f57OP0uvoK5tcOSDkA6P6gu22W1a
UmW/lcxVBS887yqbnB2JKEvb5G3Jdjam2t/Tbnw2SI/TS/ISNGbmW6DhXCoGTga9
ElFquScu57OyVGy50bMwEwzlJu2KZ6IvSx5PJwN7czubsaPlFEUvdT7Hua/KETfk
WpXWeX+bn7m9YBGDT6QLl/LJ/BkGVDnfvMJFtbmb6N4+j8F3k14KmqZ3RI2fb2tx
/Io8wVgllAsOBHpJqApJl1ctuq56MoYd7ZAUV2l1udAu4qkq8FNViSbL8Uj93uQZ
K8kjNIf3bJflePbm/XbCzlwtFj8DLPGSS1Gypjg1xvIs3aWs1+Y//wh0AsXKUDSU
5jacFboS0dSSup6im18cJCg6aTYT2fnSUzISheqD2z93MT8rUmu4DAsLh4tRvOO9
8tdkkkhsKqltq3SrepSJfLkw/7+6mQ/Xnkw9034Sh9u0hoMOUg1dZCe8EjsCp3P0
/MGMpnXlrRrIui3S9LhWGNbrJqfkIyYtv+QtAMsnGcZbVPvcTLDd735dr98XOX8b
c8poc6HRrXbFoSbeCW6kOKJzRIVQbVgw68aYcSt+aeiEo//Nx49L9Qzxu5TymaRD
Kw05Zw79WbccoaBnuerNBNpZuCS5rVGkH8O0a+CqCOEyu8hhLN0sRPP9PwUB2AZf
1e/droAjy7AUcKBw2KTqgTCpHtIuGRwUSLIL4D87EWhMaGtU97jgne1hIc1QjSAf
gHqrd099NTDDOTfbjCE5+e+YCsO/GDLhtL4pB5SaRzP1Rk/ZsGwqSa8x19RqPbop
JPArSH+p5h2e4pWckQteE0u/+voHerzeJHxCM4HQEyvUmpJq8Pc0M7GqdoaGXQcL
QJ28/VcG3IJ3/Ply8P8wYyHKl+hfNKjz9z9ihkhkdj1Yozq8X7aN8TVxdifvNkab
8hmfN2i6rT95nWAyWE8oAXx1kuVTn9Gvr17hhNi85+uk+VrtRh8xrU93xIv2mCqq
T1lYQvN0iMzRenPrbM7aSWXWEEHepSC+ifwiy+KAt8INE6wiQBnUSqjeoqqiZEOp
pxrNPh1svIexv9usRINAVd76heEMtxCTt83B/ciwcpNAbTGru2NLMWW1L0jrW72F
ngMUsjstIB2PiahI5Vk9MjJJ8AT05otmN1JyC4Ky1NAZDmIlxw5i1EFAw8T+1J9l
9NG2bY5m+Lw9WIj7Zexs0TsdtSEyrh2CACNWXb+LrP7ESvdfeQSPPpNj+tl1mgCE
0oeVHYg1J07knH1GJuZc2IkmtpEO2dAvUIhm4AY/3248BD934G0GOttxwpyq06Yw
oiAMaBTi8TnoqwMANP1h3dFDpQmdpRwtKYb2KiQoDHpIJ4qfNi1bQ5j+udGdphnX
4iR2kNgwLXbFMktjK+r9LpZ75sl/0ywPe2mhhZgzHd7yp7WRbEM9l1NSWRRGT/vG
1LMOjM3BUi5nz0TNK3Jn3Kh0iLOVEKZJDU2litJY5iC2HLc3f2Poc2wbd+sXTEmm
owfgvC0Qp3x3i7rmX2wYRuqAwL186e4sQePYv/RbODfTp7IA2jAKNl60ILrPg2bo
csC5liVerKEunhuKIj6hvM6tcz+fucYdl3UTY0wi9X7teDhGaf9OrZU+xie2JiO7
IVTFAMer46wCYRR0fiuvBX1YRoO7RgJvHn1y9gSKUtfrlFGpm4vhbh+bnT7Fxpes
SeI1WxPj5V9ysIdiz8dpKhQa5aqBGIN62mNRQKTW4zN5qIF5a7tfBKDduVFAcd6e
0JqQPEOYpLY7iV6/dsG8orhhicu2hVxrm+01NqxDolyrAkRhLHMPYd4GHZhpj+hU
coeGCKAM4M9jo6wceBKwGx9/+/QF3GDN+p+6EJXb/lcBo/jQvu8/82TA3TR3msEm
Kt75i3vInP3sDjU+xWFW9c2gzdqBe61AH916uXV5Ftx/SNdBfjN5aRjlQvEPalUv
LIFn+A7gRMMEaPwybDsYLDNTXnyukCyIRNdroXCFnZELX42a+vasVbZC/fL1cRSv
HHUmygvcZl+FMPfMLqYIXgmN3cpiImNJHbXuiwgqGyyAZ1scNMDTsuFi9Pk6op2E
QUbsqJTErGK7KKYeNUQ0X7oG9wLFKgIRvlJeI2wiN2oifj2ArL2Du2CU9SuEl2dy
mFsSWJxVahBv3n8DRykbHU6Db77bfREfcV02TPWiDmaZ3Q3MmZ2LICTov+5Nm4HI
AdNjgq9IHNYJdCD8+TY41MvV28eHpiUJ0JsZMGf6HSkl3y3YUu6HJCR+BjaUADSf
AYAa6rE/WIDRMAsVyTYaFZACidY5RD/9pAYwkT0n27NesegZMxbnLvLY1IFWVax4
5mrwNC7NJ8vvC8feR27VTlusq7nW9+av5iSJ3PhlX3MJBtlFwn3mGkR7LYJcuEYU
z3uVOtMntWqHkljizjUxtSXg1o9A7LxQDvfW2W/v8emCHfcbqpu8aCcmLselDbiI
ccOqgQ9OqCp03hVls3v6jK+1zIyG3cxVD4Kunc9D2bpil8F3E49ta9ktCYdGEAXw
gd6boSvThczlBgp7Ghvf2IU2icr1PJyL8GOt/RYd7hI+ceMI/rYLxmtfNUT00nmO
fgkExsnIMM4MDZasNFjRzXfjoTkxqml81GedUVSm0CfQ1RjcgYwhElWYOLqJMJgg
hRrLup3JpWrJcOe274NVNrwaGp6O0x6A3eIWNlhA4Re8NnwEcO1BZK/g05CJiDFz
w94ftfpjm+PjOAo/lp8+syf06/Nj4FZfXsXILhZ7DgFn39Lacimf/NRdM+9fkFH+
qd4gig91yLX8v0zMTox5OPSoeOWmag6Euy1QcbfjivJRZkVUxd0nppfvuTKlCGFu
XMBDet+AMKR3MRhmx2rIepS9Dq0TxB0vfcVnXsmVjNpMDm8s6DyRfjt2dHpWPo1j
r6uTBnA6apolBVezz3uXCg7qFU9HyP6uRD7VScEWWRKL41fL2NOqEgzaVfDVXInF
OkB5XNbKjz51iFPT8N2MJtgty9Qqq2l7q4Ilz9PKivDO2mU5eyO+LPRFr+epYmyy
qp57lTmwWVNgSaCLd+Kf2DkOfUrcZaSjKDRVkYLVeOMH1ZNH9HSjsbSxWkIqIyzp
mqIrluZuubRaCZlILz6RURllZDEKPNbVTeTxtGWDRc2XSXdVh1F5TRE9EKxIH4QO
R/psmBmR1WWhwCl7AFsFR/bX8qIB54/WeRm9nkWIy73hXG3b1P7U01kQy6gG5r6S
cCjWmCI3wRvIiyzOwMpQTXFJZYgh1voUDxIu6xn8iXHMDOgeRBBhJ9BXizafrn/b
wXMEATJtmsw5yexIyX8oF8x/BsSo9J4QJepdJwTrfkqhG0JJh3myl4iT+IT+P6hP
ER+XxO3xEkFJr7/WKQBAcRGUy4sTHz5j8v1SaBsiFTfrX575lHYsQySla5CxSHQ7
edGKVm5Df7jgt4lumO50hrLTSC+ay+rzyFsKssZwoPoucp4igKczxe7EtWLmPBdV
bvfCH/2R3Q2wyuurVBcMoHT/sMGJyc/jUQsqVg9nD6u4jcSmcJB2k8jntIuUXVI1
IGJzneCht9NFzIJ7nDCTI5qJAZ9jYKAnAJvh8i4fWMINxooGjTodHdBbTH+sm74d
Q5YfBZhoK8BuqOTCBCh3Mua3QGmuIyajPVmhJnmNtJnzutvs3wufW3Gv9FXhxtnI
Pgk5m3IS3vWZzfT8+he6GjoJk2uxKmPj1TRjbXzHbfy93Hzy+87wPgnUywNWLPWb
783dOpj4hGnP93Q9eEp+DuuxMuc4trHw+HJF04R3/f+0YkiCZN3VGrnqgjqQM2i1
k06b1t9pvseA7ezFh4DGYQO4jqxnjw5Lz3AUo99Y2FdTuxiuN5zIWTk6dYKvH/Dy
T/MhjCtDud5K/YF9fyDKaohAoQF/dylKIOOTIMpdOX0y5BeSr9MTvw2kMgs+Us+G
+RsI5HKpfDPzhW70zBzSq3UbcHZDlMN7jS0vB6MvNS6PUDccsCZHg3zQdjZVA4R5
dm+UDpZp3AJ8tpffTLkfqVeaIrPHMdx5YUVeTl3c+ujryR57goO5HTb4LQ8XGCOl
CeY4jmaJPEwobug8B6rPe+s37DyFXhOJjVM6ClB1YJWxGwQ2U/0WX9BB7zDPz8Ad
fP4sp5NMWuGHBCtQQAtBSJO8fTjM3cuTKgHv9r3V6FNT0vA7jAwXWCL5GUgCcfkG
OEtVlj0y+6QCKgOZwxeQ22270oD2J3zHtRJVWTgF2P7f4Ua9GMevIoGTzw2dhMAx
Nbmjpl1N6gwwZiBL4E5b8xpJgedJHcPcDyhMzhhHiS9D93378iGacBvB/W9FaTOI
jxhpmEXm0AgBCH2ONV+dGrW+YO/i5fMQxQJnsY4f0N0fFdMY97hHbOwqDzLlCfG3
gjPnXieb5CfVH2f59N71GGV1jdYxiF6f4uHFheYsiruQP9nqs3g9/dZPk8zf6Lh6
f9fXwSP+FFHHoC3x4yWcNQwZ6Cr/+ZyGrCkLSEaro0QOlcru3Mv8q4zgdCLnGdga
UVgnX4N26LY5H7lP6SlXYhIOel4i3OKoilHPwU2Mfs95xapsFHqzL1JlaxYD9wG1
QPgB7VMAhhmvafeAyzMpRki4KaNM4g6KMebMbU96CQMn+zbhgCX6OiGPQqlPtSbX
65WIqN76gdcoAblqZ+GvTdX5XF7wdX6zSf+wtdYrqpS6666HvmcYnY6VsVFpR93X
aR8VFbeqv3c7BfIn2lzELFH8BvPON+5bKXsq0c66AWsS8DTnEEx2eiPHFzoUiY/u
4tf31eEVVmzupCWeNbQE43m5ax2vQKhNj2NZRFdmNTNovIdlhRvxY5ceovFqXGIh
iZuvm0nLFNh1TLbASPjtRhHguxQh7kQzmVgJLfxpyYmx1tC1C93oow98cE/yDh7p
owCfqu5mEO430vGi//YdSMcNIlz+6JPhR707T7041uovvCq1rHcYOY7SLN4xTHiB
of53Hxx/sIr8g7qyCFIRiQDtmuIQHO72X5FP2R3jxRiG/N2I3MvSqeqxrLhSKG6M
ILmCfDI0AX9tb5B54EdxpOlBB5n/HFu6XJMrDgFawSQYojoNrAwt9MC/U6C+oc4b
Ch5gi3s0PrLK/8P0V0nrMQSbGIACKnlfD3YkdE0O7Kkhu3SU4ePeZ6ls1S/BozSq
NkvOgiBkgx7PTzxRyUNkfb9Q53GBn2/fCS71EmMYSVEDlZ0f66Tt2fGpbxHUrc6B
R/oowEb+9hU5x5OcjESIr7EmHYvdI+7G3jSNgu90QmfFqZ0KTsGAUt3mNvuo88Sp
jISDSfyRDUru3vYQpnwrLBmmh/SQ/PFf9M+t99wm6h/9Q+43gtrhf5X3J+7rCasB
h0HoUjQj99B45GNbPmpeh/BhCZQeVCvnhaIxvA5C41vjlioxVlJU3TicizqJJnz6
fCoCxu4Xr6Xtk/9dYx6RWz9wNO77iCCdyv53T0qCXMgqp/DeGwYsk9Rbk255ajRn
0HdxBqp7DmduBg+kl54nr6zJbTIW9RDqcMwNDx6XIagfYTUmdlKkq4buriwLo7kW
qWJZEeM7Xn5LfzsdoB5XrqnBvy2yw/TXAC3bN5ej+Mb/m3dNPKZS3lHtJ+kCdtpC
oHI39IpfoIFlUD9Orv4pcK8MO3ZmlyByMeQ0Z6B0KGy3429UpbwYceIRwiaxzk4w
Vx1TrkqL0/xTFQBmAw0Ac8Gq6Gqikv6T9YiWSmXZHL82rRrxp8IcSUdy14LrDYEm
Dc6sFvvemJn60lH0euzbL23s/AMo0UEUDtnmwyHW5gPg3rNmJ32x2mXpVOemBOC+
o78otZLJqncsvyLNSl8D6aWOP2dd7+N8DlwL3GbyC8Z9qOrGDQwL10ux208Gnm5A
n/OvdW279MQuYTke5Fa7mw2ccB+UFa2E9VGe5/+D9vCL4TTVYhbE/V5s4Jp/CbO1
hP5s/55OIY1Kx66ELuKLC4TCWyvgInxo1lnqOyvL3tzt0WWgr90TCD1QBDpomH1i
7EJ59rgK7HJSso9Wqhi+kqZxm+Fg2b8Hc4dKASTCHCU0Rz0spiXpnoO5F6j4Z+NQ
Y9OEPEubNsz9bvHdQzVskTldVFPy/5VIHnWYwowvUuMMXZizcHbwuMTLe1U/KcPi
N1xEiHFDTL5lTGky5EYetP6grdIefqFbDLDxU4FwcHMtzANi8PK0x2c+wF05nun8
ARh49/1lbC6YL5ZVHRIGnnpvFYGU8hoN27xyBdJnixK7AjgP6CCZs/9KZSF+1CBL
YfqfefphpYNNrbWqx8K/c4wWGGJHOSWI/GEdiIr2FP7Dah7waMlJ4LHqn1I2vBxb
rXU0d3ko5OVEKleJBZiehQVWGEN3MoQ+fQ2V18ZYaT3ccmz61h54AJ6n+Nqg5quL
KOXHZGX+N9AIBgreLojPGAFXUQLDH7LCO8qs08nLG+ndfPBTCzJydC4xbYVvmiqd
O480nRy2j/yW+ki4h2nSdRuH4BM2K0wKDi/VaX/+ZomrZUwaYwrmARE0tnxFjoD7
pToTyzUzv+FcoL+D5RwCtMP0GeZUNp1VzP6LgG3n8HBZWHpdSoH/gwuh/Em7AdJo
RO/8mYF5vPc3ANeviLIIoAY+619Ww8/Q9esNrryxuVeagixauqvZ3GrnmqZWfPFb
4tmAWz9aiGCPEJ/RrbSRX4AWtHpYECPHhuFuPjZFI8s3lp9duZjmKRPI8pwPJc5N
KR81asQmoNsV43Sl5XVzwJ7grgujVKc0CShulsGjLlwBD41M78woCxEPAWNMHRwq
wtzKhzt2jsUeLhSyYMkrlGBqlWnq76o7aTFAyvOk4IaoQK8Kqe/6fGbr2mBKHHyE
4X4bwGCOaG5WICCSyO+zxpeqcTzUzQGNEyZZSP2gx5LnOfoElFL3PGmR60xeqoel
zvoYtZuPb6GOO1bnIIFCzFRH3WkV0thE+xJq5XmF38tLidORDDWQ2s0ZtK+UHcsX
HoQD8BjitERocZMErb1xOluAbc5IWRfQ0ZR7zPJ8usSWZ4ts0zcP3rl0FzfjdvMt
rgd/zXK324PhA1IZUOwSF2EX+jc+ZbNeU8AMORtDzHEf/EbLH3+pQ1jmQMP2sQiw
c3NcJMDHn0pdhd6xxG1FFgf2vlCWaE7V7CrXx5aKivZmFlftxqPcpU9ImzMfj1OY
kqiz0sPgchuiYdyKN/wt5dbZhiQzfXpdsAYiyUJIB58brgccQYlGOguop/ppSqzl
TOUreOC+yFKvxxIyNGaroskEf52bmMpafBlsLvEHF0I6XW3z+2TClFtAlFnGJ1wP
HggyzqC7qT3Sr4Vn2XcsZcmbwUO8nUViSm8hk5Z94T2OVunsCijVGcmFKMW7m9TB
vz3anoFEvIWSjXU6mFhVkCIYYq1QEO+w3wgjBNfsraVdIWuvCkPQ0+sFSTDKYG7t
bmRG2EMFyiv4SXsIyz3j+6S3hKvQ+VbkTMZF5StVtobTZaGaZ97q5pLcgeY+h8id
FyVXG9lrATTWejgV0DTJZo5jnCQCw4/30pziiV9W3NwLf7kCtP+xlNVAJBhQgaMz
HxFm/pcwFx3c1M5D6oX6BXzKLItf58BJqn+xvW45Vt9MfvYEUsfpkgkYBzeVs5cE
48x22orbCMENFYqnUulgbQ2kvwKcy0EBrdLpH4ES0duiNQYZ48MjTFEav57CiwYw
Wqu6n998bzEcT72PBJ+SNsSUk4Hc1Z6foBujiaMZaXaLENtrhs54zQTy/fWK4mql
cRo2lV7KFQZA1Fy+6cdil/4tjpDM+7Wq+u8C0xia2C1G/Rh7uRDELkxvEiSR4Ucm
kkyFIdWvpUquCHb7akpjX3GaPBBo+LtY8BCF+H92CqX/WEvFPg+tPUASb8hQg3WJ
GiGBY+FVqP8fiia/NN1jVny3qPDY37MXRXR8X0zpWciarV9+QRPQfJ08xUnBSfjz
Rh9lUj9N9xqM5ioa7HIMngjd47uUrH8YCySJ/GYTvcEJO7ELNIsgpDG8gPifFufo
KzTdpdr0ydAh1vkOBVv3RTi2y8nXgx4Sw5LjbNd2OAtxj3oIuLyZobQoO4ZiJX24
N9sEW0KHEleoxx+JtyHl3ebZdRI3OikikkWtJiUr5WZSOmi6v6Y7zApoXZ7T443H
EXbdC8gjoFp3fmQOlO27ZlBM+Jnl6cRdGTZJNctuW1+wcGZthP/HhY6hZgnLkQxK
6krkD6cDFfCKPdx42yPGXs9ZPQ1zXtUOHaDvj9o2gtHtTLeRqjyJ7/7cO26yygNC
qkIpTQieomxtBNgayy4tmNh1hsk+O05nrh47kT7vcO0G1SX8Fn4qb/Y3L8IXEwVP
2IWAieH9RN7x62C07u+fEea4YjEXxwPM3mWexl4LS9jYwB/Mi5yR/SRKxtDyBTcm
UIP2mU6N4gz5J6VkI5ZrzvM1HFTaLgw5Dfa8e+UpY0p//rbC7N1S5ZZxnPmMQnsq
9w21orsgI61WZn1eRl6f9NP9EzpsMnCze/lj8rIVAry7HvRp5guUAprEf2N88mMl
nhggjnGdGXUvtAiM1RNWY1nFQMV1/YX/1xEKbWu0BsGlwDKLKzJP33q7a55rOyr6
zwSjMfYT3QHpzHip4yjLpw94LANfiElNLzrNbe2TKdSzTO2iym1RjA/bCUI6qULQ
eoycPYucd6MHKcAeAkBTuNtnFeT7lrxDRFeh2lh1uShQNL501jjEOmtVSVnFVETY
eZ3xo0xxbp3QC+kpVKbrQJsy7vP/1WOybj8Kz9yWpaLwF8e/wtBPId/PIT58KyDI
VF+w8c69+t1rvx8LgHlTIJJyNIByj5pzvose24Y5o0uzq9VqMFcCz0OkdEu7Hmzh
seZQvfdWQeydui0OxFuUHnITnqAhZC5pyqhU6PgQbN8OBB/IC4cSa1hTnqwUbhdr
SAMDr8H1LmT33HyOQjkZF6ujP6leIiiibBJCbUr/zWYmXN97mDKGbZKYo45mwQmk
V9K5t9SFA6aJ0yEGrOT3PIcn0b4BfKqynGOCWji7EeI15KINdvcWwhyLRag/Z5t/
4YzuGpMeeugEuhO/AywxnlA2GfAB4uExFSc7dT2bb3piPxrsvFh/Qiq+iuMVW7Es
57/g1/JHgbvs+D0kiyVdJQ/ETfgOkNQCyOPEl5nrCcyB+2uAEXeOqK797VzKWiEG
nAmKJVLxgsr6C3NxjOV5/OyMm+gFsBvzXmxph2RNyoD/NNrDUmQ8XWk4Ci6wo4aU
gfuzQNDfzq3xRQY9y3U6SKmu3SgAQlTm9UXSKsL2BOpnhbOHh0xX/pSOJCX8nRHe
EBUuEelHU7zxijKs22EdlEkQI7hCIvq6zhMlhA9254sTs7vPOmbxaa7Qj73iPtNY
Cl5DXQho1+1zkrpLBECi5gCDnkMGiNIeiM37IQlb7nuevqi37ARFKuRftGgaCwcw
aCdHZGxc9bD9EZ6oY+jeFqGdmNClN54Xu/PAoNKYT8HVY6ftPCbxAWG4+y0220CP
/LrRQbhAlYxv9rILTaKRrjj5bv/qcOkzZzfISyWs0CqplWNgsPmwvy2n3oOy5WFY
6mm1deSsfzmgoi9Jb9zLxf/Vj1hhD5gXJ7zhwTSreONb77rlyRtTP9P9nHiGQ/gH
6M5MwfI9QAmwK0q8JMS7JfD03IvgSDZQikasIWLNcKhDlpbK3BnDhpKEZMEU2si2
3BCHRUy4mMNIX5iBs4hqm41Rtv/iD63HgAs5DA/GacRVFCpBSBEu11afqb6rBh1U
KOJDdjeBqu5hs6V30GkUZdYUw07emZUnKL81flWsn2vSehXeW7Hvoi2OoEZm645I
B/liuk1rMODWhhq1hBt06aXc9tTO1V04xoCotT6JLaupo+gOWmkpKNx3KAFISYXl
8Mqy3mpecODPR1EtRKMXQcXObrK24SvklhgPm1cSMzC/7g96gM2eyYUUT9U1POtM
vKxNb6Ci4bMvtay2VAMAF4tpCNv3/ZAV+fzUi5gi4MnG1pWl4Q3FrjjTh11hfUWd
v2vqrASjPd7NyKmbH8Y9tCwFtQ1/O3q2OZYW91UTprJbcyR1FCq30y7gTVzSXJ9w
gKFOkuV6PJQQkg55ttc2CmxkME2aaiGvN2Lbkfn2W+sFiSaX7sRQ4qNJqPAx79dR
yhVHMA4aV1XbI+23TrUBUtSIMKT98g0az8o7fz9rJ+ilDYrtys05TFiuKxRKs+Bm
z0SRoJSKSypgkpTf9bDJ396K3vzSowXO2c0TA+Jx6iArArNAwAhqNZp8E42jd7Dg
1oWcqgX1GIw+ucOtB3iODsY4ffnUo+8GwtyVtl2AnVdNa8XmGZKcwPpxw2cxH1Kz
CyhigFmDp5M3H3O2XJpJcXYLIOu2p547ZgqAJI1SIzx+LcSKW18CFmCzc+2G7OLW
U4PvOjYsG7OLZXZ9Nkfk7nWenpoPkHiH4CETrmFzDyYVwK3oXnheym9Yhd80MhNc
t/mJP+EV85rLnZmPi5q0cTfFS5i4z/SXiNj47thZNFgnb/fYJANW3ITOm9hyCaUm
IOIiKysJx7vQ9MF1Eyg7VLOrlKxJjD/iOPAyizjxPCrrw37GXBCgm8TwREmXXId5
XUJj51kiT8YHbijlnFaQ7MPR6stRa561FNLSwWZMyVmdfFE5o1zrG+h9UmuGKN7M
X1Fm9dD8YtwwhkcKpQS+UJBny4bsJwlIDIpXRYYq3iqAHbjUHIVut61yeYNwTQTq
LcGl6VhY1V6SAcsSTt1mLHmeWObbFMZqVceYf7NkGVMXOtYYciGSkPafNaGZPAua
7VS2ITgDohZJa/v+tOOrVM3gDZDh4t9KrlpAsEbnCE9NTk+Pp5V+RO8LCjZwq6rR
E8zv4EGGehMJfRo0rFPMYOvJHGL+7oo6Y/SlyZRKTMiMWezcFpEck0M8LV48Momr
3nEQ6VdBKCZw0gAv7zClUlg41WMJIpMwNslFZIPodkJ2KpidLcnSj625bhlyvD9o
YL7mi/EiloZQqLI+IY27b53JLK6l1D0mutOk66MLNnshbwBchsJS/xtDr6jBX7cF
aBRgPf5d3nabPIGHDkmArZvVHwRfLbqLcOx0W8UKzo8/7v8NJsNMKNMtGH6w8fOe
+7PIK6y7mEL4QE6drmpsrHqn1Y7C20stGvmzWBIgSmKcNaspy4b4mONmPjhPoXHS
qZu+VQVqs9M9waM9MEGGWULDoyxKKgVDrtmU/jYqfiWB0n/2sBo9QhZ9ojEhC8iD
9UfyoC8sTXmMAe9ygTCLTS3katxV7pFTWAN5/621C2RhacPe0S6cqrvVv+VC+J7F
PUSP+cr0ATmPM7bPIbJ8uMekjfdyVXs48ROE38w/cLlJpjFq1MFEX72etNKwrT63
7pxvlQncUyY0hGT7XDM0bqAd8GW0hQXDuaGcPdx/ti1OOgazECSlJ+caUDs03vib
idA9Uvx8VK4fbj86cE2Lwk8BDCXrkhBwJ35aE96n6A+/K4nz7sem4Aupt/198ks4
X0RV6vSoyAN9ijTZJXpK3LWCL4qbgdbYl43FDUnyT6JjoygJ4Ovw9spqqC1DJiCS
jHaYvq3qCVmq+6NLapUsgpgGHkS0BEXBUz18u4avr2BeUGRbS7uXBL02WFWQckdI
aIXuqsrIGMmYwXEDQLMjJeF4p4G2QhghH+kAw1M0+eiSKQUJovHKHgzlMC9RADba
ulYBXqMUBNNWsx0WUGTVVpKSaPZAU1BVMsPYJHF0l7ry1fm0s/4hQ5IkF8M1AjhG
8a54O5kipWHijRSTfB8VIcuweUQza6q6rru9m66KPbJPqi1Wbn+vtjizfTjwiq13
kp5w1E1IDrA+2pbqZmSlJ8McMBeqVgMR82axQBxm3j+reKdQ4x/mVYIb4Kf+gqHw
1kTDh0yaqUn5R3/kjqyGWparxtmgS5quJVzYkbO7h7nuGsZ+x53t4gVtTepYREHL
6jdswzM+PnJMYQvGxXvruMTKSnJbaKDZe2lfwxmddzaRBscRMIPujjmOQkznlTZB
PbSrHP63SAvLsYnxNm8b1mbYloeAO1JkC8GgqvW7ta9PX5pEmuSH4rM7AQr/di2Z
X0E8gl8zvHEgKsT26gD9Rt+Y8xFV2X91bTAnFS0Mz+4c8B+U0Z6VS77017jx3Nny
XIzbpO1zZtt1cTqKa+Vp0lmrpZy1anPVPZfqsNaEeruiXQpEdsgSDl3RxvR9lzz6
HOOojLUWo6Swc8wLuA1hPhOFwHQKGj8HHS0XE/K0hfbVT6Am++bYG1jHl2EqaY0j
S8+qkeBYR/rNdtr6bncoGMVMwWMU3FSzpLFxYIurD3qgbA8Yt7lXmyzmGjNXq4Qy
3K9jAiL8V4JG6W9WxaXh6X+6SBK4P/6VN1Zr0pgdgSGMFJBRKBDD9pwWa+ByZ+a1
ej1hZWj/YGsvBs4cMLZI+HjbkYBYu0WfBgXztGOEiCXe3gtuvkXCwOVl3KapR8BO
u8BcBRl4tipBtW2aNzDozCMyZdxHiXXHbSLhyr3nLiYBbrCh2NOiLEM5E7FTbTRt
BrHJEpwuhFgHjVH8CkzmbbIRKlDiB5SUlPTfwgJIGn+djhctfDobiAOsHaLJAG4l
W2L6luOwjOPj4+m0StBDb4nC6YWJZC/t1fTQw7MPTFGqXNsw9kukgACYshpLengD
RHIGMQ8LOfuhIdjCbirIOHZSX7uSH+TeokfLiKAJFCqXarfV6Q9RLG6NbBlXOkbH
hKmS0udLcQflWXhXOafUQIOIT9alMXIGkokQulSFsiJ6gWdaAIVWDg1Ara9CtmHo
HULeep9zlPGIYxlE0uw5J4+NkURw+YLyZRkNc+JSwOMULKaSIQTGOXa9YM1T8Lhs
knCGW6WhAIoRaAmxs4OHkKsezCDYcu9YBsu9UAFU+7GLsYBNprS4LJy70H31SUj8
57szCB0jLmkrF3jL/KPX1wFM3mx9TLKo2GKgZWERJifjqkIxuaLlup1Un54S4pAg
tAyeJtaCdGZGiYzDJj6niEoFAHZL0M6aE9tK3ab0aDtR3VOCuDZ2cKgAavkr3yS/
KbIdg10SVjcPt9mvb5Omn4J4lte42pDyGLAUBUGFabGmD7LZYolq7mt/uVzCPS43
3Qp8h2/PgDi5cTLxN7aclCGymSwGaAZre3G0Ym8Spd/wgLnP2SFaqR6xzRMGlhwl
O5KtDKo2RbcQ3ULjq4nbnG/95a5f+XyyCeszFIxiyRS8Y9QXHLNmqGCf2wVtnmTi
HZyDsFNZPGMc6ybhXcB5FvEOEUKY8m1HpyZtYPtvvUqyB6zgxIJKpDKqkoNkgjoK
ycoPlvacwXLJIIRI95+Mzchk4bht1nU+4ndGLtyj9DTg7wSeuF4r6+v7u8IVjXl4
N20zwJzqPSXS2MOQQ1ARlSky/9miAu/bYe8nhI2QrcfXl2XREfRyP2SFHTWnNC7s
+qmIdNjxTeLDWho1a315suhATCFR+5lX++5z4MFit25q2oZQ9uZ5F9wzlxH1Cye/
M3UMIVXI+5oagw/JnzJ237GYUpBSJHe+OK92WIaDWOYHanEmrWpyziyJ5iVf7H3S
2d0adDKhkKmH3FvQJGXOtYbfwNqMxnc8rUc3qjUgtJB3mZAGY+jQ/1IDYep+d05Q
sjNhzyXkjvQRKQ3npVnWVdPMZB88ZyzV9T6vKe9chvi7lgAy+9mWu9guEF10EluN
MZMDjX23G6yYur4Q1sM9ATbREPaOZrppW0sgc7dffGJcsUPHoEGTlGvJTFqElQwo
NJO65Mu+/uI3phUTfwci9K+Bc/IPgudojDbdX1ElOFQGH0NSogQYOjEWhGyFRhGh
/5Pcs0O7E+P4FFcfuLqYL89PVgbAD9QyF4hgzNmtvvt6dtuV8gvaotqkXtxQccpa
gzIVBvcmzjHVgUI1BU+9Ku8fMdRvab1m0RFofLVBZAfrtj3DilGSV/+aw0Dubqyd
UHU7/APCtsaSI6M1LhuMwUEpCcxSDrvyJXt78UCIqxw8g3JnyPNqQln6Q6cO2l2E
ZsX7zbzqpnXHv7pX8HmsP6oBjb0b4WO4Vg0vGQ3QfGwbEUsHrAymUFhiqawMKhtb
dv2slvi9MmphrDe1U+bbtsNSeC86CvW2SULwMi1Iu1SOi9x6T2HcPhYPWKf4Qc+o
s+ekk3iBD6WX4AncU2ZbW/M+VH7Q+y6B6a038LfPbIwHJx3aW6/MMM9ppJrtgZit
NKs1AIf++hm4U+2jxhNpMKAtcquTjavsAkiPEcSua/0X5Eyiy0EXElEm1zKA2S1q
169exi86ch1VgjH4dQEbetOjk7/Wtl/x4ITA1pNOOfvV8Rz79KtlHF97XaszrdOl
nh1MqvWDd9AFm64cOBKc/kZd1rivpsAbFwtYGMlGtVuDcxgJouI8ygKXv2JpnqWf
dsOQiE9x8jWN3IS+/nZDZHgK/RGFS59jxRtjorqEahz5hwSSmJcu5GyJfjlGzlBB
sB8yC+AHGmr1WY4QLcTpSyFrB9A85824GmDqwI5d7eu3+yzfnGWu7zkuP0ItmWWo
hpAWrY8EeJ8TIwKwaQ5OReaSkYe6/3B11BqAhVm9VwOo20nK51BA9dMQcAhTh359
jvPSSxNYxoDUJpd4QqH5J8VNcVbLXYDpsSUkXPZJbVP8I1HZqBk1eAAf/EGGqz8M
QxfSEBSyHaKbB38BNgktox1NMZbr9ns1SYh3oRB4zojHl/779/Xou4r1qu7tcOXX
0bo3nTBM23eNFDihzxVslCXYVhwrwDIe9f/Oj6UX58zXUTP2iF/ixYzX3fXXZMdM
0U2cFwwkk/GD9VQUWsuP0zCSw6f3mdsUxNyBO+I6M8KKPIZDavG/1GGMMBa/qD5S
qlJgFaItR+D05I9d/YdsKKC8XJHjsYUBlGOvmPDv0nf3lQ5uZWH2c0soQzdyj069
e8a7TWxes5gQBDNQ3tc83WuFC/EQ2F6mZUZ4diRDPzRshmZXjbrTJi30PDgJsWAv
Z4cW9FXNm11djB0T0VW1kHkGKhplqTmmSKhwLZ6UmMU2pqTQXDHX5uDuEGxYQpyi
qIZpaqRY9YrvGV+Lsn2YCVivQumINefwCgpELKQ8fmuHpgCLM7xyRfClJSgyHp4S
SsqfwRhb1a5fW/l97Ft27oyiM4/tiuDLi06qJPI7HZPxrz1oz1ht8ELteZQBi4Z8
DBy7f6S5PPSI0396nu1FEIVe8wfk1bidfVL8AGzH2iWEEpQveR2VHcKzPSBzEb6H
6dOBUbrbvOtYUgQGphhxCEmFX/eR2ns0SC9VoMv8FpO87/BP++8DAfunxRTbtp8b
OUr1zYu6zEAkjs0QxH96PK7nl6OL9JqK8q8yoLH7V+oxePBYNcD+rXcDAB5APo0F
lJIKAg2nPikkqMtHWWp8b0+dhFZ5JpjPE0SjspGGoA7SnZew95r6bLbO1TFKVJkN
nuj7Iweq3Vtqdh/j7Lb8vvmOG76y1BBnFPspOfRFtKvuC5i3Kmj4pqZdYkd08mr/
ENKMtKSZjgStIDwjnZ5hdooU7PfUNHLiAii8mD5dYO6ydmZ78lrrYttFaCmbwOP8
iehSzIVMxDpCkFUUbkhCqZdRhltQhKkqnGCw53Ny6/Eg5XVU1BJOXOG7EH2XhihL
tzdOgqdt5GW2gm1ecF8vv7npBWxlKfyoSJjB5CXA/xp0jAkakz5rQlrr/Aj09a85
IhNG9iyR6gswmo4Z8mwYxVSZ/3NUdea9wu9gxSteKzwJv5ApLa6dAk50fDq7EUg7
3kVaOXkB3hjHJfZOAPOyDaYkGT2fZLDg6MJuCrSeYCGhlzIGHAyzqAe/JLo718ji
CFEWD4Dby1VG9dfFzHXEKsi+RPZshGZ4ZtzG8Jt0jYNqTLlDL47yKQvk+DXLW0fE
2gYzpf5a5Wld7q+NBdWV+e4cRttoMtAmAEKC8R3CSIdW89uDLx60PYmvBnZgVKRF
y0KHszxaCEjgI5sb/U0IELG82Vi+/7MZJKYIsPbbmqyLMtVywKJxeEYIm4KAAg17
BLta8VvyesYVG+zWDFboDhshxajwysNS9XZUOyvunHKABpe/IM9/GOIyL8gAulMf
SqkiYs+cxH5GnTdd4+WX5tWw169ZF4rKllgN4rTm7i8oGWk/vhvu/umTW/UwUurN
l9TAxgOE0lyUgI1e7Ul3ppeyPoId4Qsq2Oq5Oz4ui7ggutX0sbino47EcdabEYKA
2C2tLFjX35vf4XS2ojJtbJPs2xPn3sTGDyFWN0klG7tvN/wdrcEv9uYsYzKWkiky
KfFTdJbwyqMrQeXKbXOjh0RBUa6xArggfamCsXp4m8+6Yi0nM7bKXvyc0aVG/0u8
Q5AvHdLsP08roamSi7P/5QoKrpaTo5WhXNv2G/8DLue62ICId427pist/8rYAomU
PA4i5fYCeGtyH+9s7n7nQLwOInpgaKgYbO8615y4XS4q5Mrx90H+hBr4+iaAXTF/
Zeuv5cgjJsCbqj4eTVAJMuLkGyi2HjdTpzbuvpFKliteHUXCUUzuPZf7BsF7zDLA
eFLm3kcLaT7tQd62x4q4LVfF1vunNjpoLM9hRxnBfebAin27yHCQVgwwO+KV6Pem
k4z1vRgDoTc2KOiOQvN6GxkYoBju/5ksMjwkJELyI4pBRYCs46HlSd1qXebeHKnE
pShoZ2XscyES1oQIjpubo7iOJw8/iIJTPM+jK9ofe8NR0bcb/PJiq6ZSyIWD/m9r
YDHnar3OwyENWsc8GPnmA8p+rC9Yq6utjuCJVnY1FaXVsh2mOB4oCwYdDwmwxI6O
Iw2StcIvjJCPJlIcdwF+3PDJrbkjNrfwUjvLHWJiOXXfi9ZDFGYVwHkWXH73fL5H
PRYkD52b7+aS13p2wDSiNghW3Iz51OYG2Uq+cGFqu/JCnVpuuRQ1XjprGeMH2sJ9
bdnnLRJJ7jBcnwXfus6d48J1sMk7krInaJmy7rGfXs3ZVPpp+avOvxxRCAeUT25B
bimVoziRlfKx4O5IpPxU0x1if7aSv328QmaBPGwWw/nMN/AHBWc9pvG3rBWPxWMJ
8igWjM0/UyexG9BaUozmdtSdRCs2lxvUAgqKUe1GoG+sgWoINkDPw/mxZRVGIR50
PBq/BO9vfiDYof6xcWdwoyqb9+vqjwRUa0KH4pPeJu4kboLvxnHJ1t/jh2mDgXm5
1wVaXoGQQFjN+wrFQH/KWtwswrw39uCCSbuPp/ZtMFiHp03CrNS33Mr7dsxByJRu
yLaYxgFGflh98Zuv74veXxWjhKq7SdzzA1xz5VMth+F/pNzhbswvi126PuDs8gyD
vGf3MmEJz/KJFGQIlNfnoSkCXBoJ5v5+ps40SvWPTJdJHz4WOyjMoRmY/eiPnshO
8seNi/LuSrdytNCF0kDq7oxNv3z6IksLSAca+Ubvuz+PYmcnJO/R4YZLGgYoFqUU
PEmLvnuao6bUhiDxyH/m3zKo2PgsnanP/MnbO47t2nKEHs0j/atpZvWYOMHPXjXA
pWNHDeILzxtUBKXGaNuaaEBLrCU6Zi4hDKDd+IF/S4lbU91KcKmhXCBGpqzdPE0x
hBv3SFcESOSqfIqwE5n3lMv1fGMbxL91ry0d/OOPpVeGUEvxDzcvgCr9dAz5TCAn
7AZ7uzBiYa/ETm7+96QezTsA86mYpvjCk8s4+DyEbTVy1glAvefWaa6uaDuM0eEh
Y9M9GfyABUqV4jNdhevRWX0pXQlbaQ58pT5J81gurCCCh1b7QNTvceFpuUuwMQIH
wfCSur7hragwm839qmui1sXXbXr1As6OgJ47C7ltYjhqBBulI6falQCkfKs3F8sL
qDUTeJxaEE/i16A67TsgpTDHcco8w43VV660QVEXoumE+n8zkUnGRE10RHlK/QkD
zH+ZHposwT0YVOfIG0FzoQtAkBQivB18WuZiZzuUeKrlYZGFV194Dv3nMJGJDK23
zjnY4f4E/QOjWxzvA1aijjSL/OY1kgyYDJUJRYrEWcdw6/TXQL++mASJcPSVGoO6
YzbVKlBoYDKbK6dgOjGMGADK/ZSqr6kZysvYitEN6+8YVCzHo5myXiVG4ZBVFIFn
RbkeNxpu5cza1yYCoJvaS772mMEj7EvQ0Dsh5FVAJxV4+Vb753PalbmKdgeX09W9
9lrAedu4hq937TeoNNrQGqazLptTH1PBkxyWF/HTk1vscHl3WwflpzW5G9G7bqtp
qmG/mDNb/sqzKzwFOPOGv2FQQnCEV3tkd+9hyFrucyCG4LrNjHyBBcsudUp3yooG
fTsfXlOwdnkPjzWCSZUfAbRWRhImIsY2JG/WV59h0basgl5ZDA7yHjaTmF/Zmwyz
eYODI3U+0yTilQk8Ho307e5pF91JGsfZrC2zcElP1rfqDnCg5Zsc4YeCq9os6h/v
QgYIumavjXBdb+C6I6k0sWt+1OS60MU3DmLSV52KK8wsUgoTRFdduvps4cXuDrfg
gQNfv0bzAsUyQdadsx1jA2roM6MVpvqmrGRpxWZLD2Cp8XTepAyNV56Ark3mnAJs
+OuWU4QQ52C5yInMkBhrnPS6LBMMOfWxo1Tr+YEQw4Ll7a4DWTP6l7pKHw3bSLu4
yQJ2VuwSZ1NltBg8TJtPFNlLv+ciIsd1t8MIGVkfCtVaKrj2ISYNYceP4TYtbPgo
tW5IqEtkn49G+JkxI4AaedxGcDMgqA+F96UQ5sgk7xbBFTjTb3VFR59pLwNK85cr
Q99/a/FrzdNs3PfyZrnPf960EdV/6COBtQNlinjP/bX9lzMoSlCWwIlCQBN4iwKT
uG45SsR9PT3GbA3AnR+VFXMNwVWBjB6qgrc9XwtGEU7s7bp9+xC0qYhUfjC9kI8d
139oLAqGjbBk7gh02q9tr7qhvGQfqKgA9YRFzYzmYsmPCpe6MURMhqEySZWCiqOv
7QZhRwWjPfFSw297NhtPaR3Rn5UdTw+rfjcXmI7p2uP04+iWhhIOvpmm6X2PS32n
vVKLhDf3hOMKnogOcKyUShcHpwHr9nc0iAXHVf8Z2H8+2Divl2V6QHs1wgD+xWaQ
s88ASntakQ0jwAYOYuHwnu1OpbOlBK2K6T9oDGh1y7C8hYwaAIfPZzcgEp+4CA1H
MbMAF1KN+clBK5ZZbLjOWlr5TikVjYvzghjl9oZasKSuQeE2PkX9VKxiN87D+1/m
WSSq0ry6CTfFYDHFSJP1GyTHws+mi+I0+nrCR65Btanip1N7HfN09T5gKINQom42
xEVSqGuYaAxWyrzFLhjVaHTpAV/tIpi67BqgpHAApj5JngS5/burit9xcVWhjBvh
epcM5JEk48RHgN6VFHKcGi/l83FMmJBSX3V3Em0ZKyG0wvWzE6GT0oTD96Qx/H40
nI4iQgj7HtRmHhH0ZXZKruAbx0LGOwtzSG7XphmTTfwbhV/a0pG9ntdG9mR9lUxL
0f1OmcII0EYpW7fRZWyGvjUzfsWhvlj7lV8i/ep5Lot0qMw07Ww6fDW51xOFSwwf
/GKu35dJBTxsgBsdEv/DoTsqysD8gL8bEd5EfAqoi3Z6BFwMU8qfW89fh8B7N/ad
ugAyxycsHnEYdnsHGEUXYBWkEV3bnRWk7jVHhKjQvBXi409XnQnuafNHEP54lSiy
u5mwNwMtjl/1Vdm4H+S8fOHiVEam7kc+u81mDzmzDKCa6UNFpRQjamjOm2kCyhIF
xWlheUe7Xn0ykIKmIXwFSBLOLvGQuhX5SL91vcTKCRjv/2k+sQ3KIbcC4dzTFKDA
6Cgz2m3Ui2O53lzWiKrSOs+y5qViOy8nywMFnhrelpGhQlc3aXc88WT5f6G0n2ct
CDj4CozCmBBiLdpFYMCixXO6INvhoLxUl2jgj0Y/yb4RHlEOGG0hsvFv3Qp2xXmb
JLWR3j7th+GWMp/T8/uC/dmy/sama6hxMHHlBQ6S4LBqm0VNaKJGPRj2KMsYrDVQ
/8z+CfHc2LXzMIa/Mu6pyYbWgFtWFZY3rhRQT70vg1foXyJxA6scD33EjzLgpHsP
cr9qG6YPNPLwvslDJID9daCU9v76KdRQFCjce8eyDiwrhIi0I5h7qp2N40cnsunZ
onphdQNP3UU2HdfxC1aZRXfMZh4KEaRAMHDMtmeEiOMxxkuEVEW/j8AfObxM6LHE
CcWx+9tjQLe4UlCGCyuYXczJjhJ1COlEWDI3COj7KgDrk/ptk3xMl0PDBl9A/4PE
qRJxhVClefn9dtpYFnr1csFvb9YaFBkSk8TbRwerxnGQWDFJa3+P2wEbWS4OR6lw
GrQQ2fX6Pjj0LGbrxNY7whyFufJloau1jIfN4McvXdc3KlfelH7TAcyGhFsSCscC
NIOLyq8/IfMSSXn1EdffN3EMBTta+uP3njGeucyhgVkzVq9aeTCVuk4eyo8xhMif
9t/ks0qPPvZdYyUOXEi8mg01bmU7MPSs86XOl9kfIycY6hkxmgB79NQ5wlIbmbu9
CxOa8CUjNKd97cqjI7hgvLDvTrmdredaUevryvhpF+yY3asASx6i6g2erd0UEs2h
KAVIpTP9srwfmA9AlD9WPYB1LcPj83L/EjlFA0PDDb9jk+r3JFhMlxBZZN4PrZDx
ZPkWMD5+wZriZetWCZgVL03daPBGImoyDU5i+BiqTdxB5ZHrajrUKNZ4HdbYxcPm
vxWAAtFSizeXlpLfjUoFvRUp9NJP907yECN4NIdwnPMsHTb+VsPtqJiV5iCCCF7n
yBqyMeTaBLERsVyY6N+XeVZqLQnxUFSail4dUlmC07WQLkYMmnSJ4qamMlgcysix
0BNvAM9dxi7MHrEnAzsrbSi4mnZahKdIlavdxetnipJ+i/wpk/ZR6YczWR4Bq92U
srLxpzvIcwaC42GE1fPcKoPxcyb0IuBz08a8gdcYvWrJMkPhPoWVgEXYCANPl0h/
FbXHR05zBAhNkMhc23chqFXdZzrjafnegNa10w4drpwaxWM5ImccXZWxZBc6Pcf8
qI3gVzldczM3HJNux/Z3FowSJRm+tnADDTmkK1hQ9n3IkQC6ViSWojmlxyZEUin6
Yq40bNMFD4dwLv+fQ2Dj4ikJ2v/E6zwvisxHMvV0RUYzwqHOhdzUSZQ5/PUMbcqP
AAmDJOQflHhpNhxrMAzukKLSprv+VDY7h+/Y/XAUU7W4IsopWqhX5mbecx9RDVN+
XXaxAltD/ocl07W+RnwiUTJtw/XHWTltPleD+gf0LDpPEzllleicwrgLrhsYH/2E
NMLTiC0bDJt1liffrJMOXSpf3ioVRNmDCuDC4/pF+rLTVWSwRMCkBXZKG5LQ4/zV
YZ+1xwvRPL2P/rb/bLe1H0nGydxmwLuUToFfQUoBKFJvWrD8KOK+ctw+ms1sE8Wh
hVWm2JMUMz39qDmC8lkTYiU6oLmuyKD/1Mw1dkesqsvfDx7AMtgWckxd4nqU4WFw
Hj0THzgmNN3nut5REHuMn0xbM9tPNfin7k81qoADiqNxI3Xu/W49tOLBQNJEXB6C
LO9cV9+ca24CLBA58Pvf7o1qHQi8zkKT2LINKhqnebFuxnrThfNBdwo1TWjqvDAA
y72RxwhLtNXSFyfKiqgIQhO73p2/39eTVSFY+Ye8NY+NKIVX+ZWjrplsVek78cEL
iOKIhw3Z0iOD9nvx8hKObKLDCjsCYFocJ88M5egEs5OpuGqDt2bdGSWTMdwUXNy/
cv7VmD2/cVgWx+N9wRbCSvfKUq2g7laqbQCXrwid7ML+2LgBtksS6mg3YQHd3vYc
G0SvNPbQCK8EA7C6B/Z/n5T9Vfj3cRrJZVEuKLdXkfsBYLdpZTsrrhAN2V9yaMSo
SEQWmi29OQwXNGfUwl44PbSoIw5euqeFYjzvs8jV/MYYVQVpN4gRKWnSkjNYkRFd
ceAOJrM5eCQLziaUvVYkbKBa9Uy4Sdjh9ykT4jgU4PU0vI50nD+ol2yXuiAT/vRy
jAoS9oXjV01ochVYm2EF68y5zMjgQJA7QggPlvuWyjEVsSWRC6awq7FmwjKEbLDs
GOvL50m4SvG7o8KK2SWSsm5/HCag/zswt1MlffnQ2ccR9GoupQMvMLUM6CL1ku3F
8VS0vsrmJepXwGH5ZzdG3Fgc3+MsCcJjJNvBk0kce/8R6JCMuXLlcVMvx92kFF5h
9fU3Ppj4uBcKi85kJMSoerpNh0RqX9JAinWt/I/MmJhjjDf22GzTIDktTL853Up0
7/0FN3AV7mZp32MRDH/PsJO7ZBI8Z8I5+gBM8D+NZmdtFCY5RjbMILLQP/JWjrgO
ylDGVpe1DxhItGKWh+bVtx6iLIKEIrL/HPk/8YObduUonK42MGafQ7fIDelt6KMO
lLKrMabKXA6mWACZIgzx9o0ArG+A+1p5v2yPeq8mvBjNxO6bbl3hqwm74oJh1El+
G2nY/2Kv4Cfgerd7Nm2ZjHvqjQcxQcFp893NhsBXt3uDhpaj/rhrFvIz3zO/yhTQ
QynLrpFqVyJqizKX4JhGxrAvnJ8Tu0KnSVofAUAl86Z3AmCWUI2IQdTJPulNJzcM
tilEcPoPtQ1Umyyz0OlKNRyEc0Bsnu89eq2Iwc5pibE3ZbJSq0UsbNTkG5sDmX7z
cGgCe9x+IvMg0SaBqOOGY+JVdNu/X7a9PnXQT9TfBFHIgBLQ/8ZQAmEv+iP+7/r9
Q9/PlulI3W59mnArvUzh8STM3tlLqGfTJNR83AI1pK9+VKfLRIdoOTbN4G2Cvz3C
2kJ2BOFgTOL3k+CO26qlXM+JezbnOzHxMUyjnDfuH9GcQFn+fC82dSUoOGuGl0TO
E2drXKEWxxfC92coWwxGO4LlE05B0ex9nEdt/a1H9KKeyhRUVQGh87k8Y26Jftrr
NuJvPsZ+rQOT/0kyNhZH15ejfAR0jUpkSx3qhvu3RiBAfCMHti+TgpSCsfUZP1Id
EnRmVqu43vll7ojCoFm6U8jq1fT6zP6GmlZr9KRad+Ze88yPxMQlpBjjVz5sNBIM
FyC1XVoWBVaBPQvlSIOuxYkiQrNNn3MEJbxK/C4R4P8eNGGl3cwGYH+ftM6yJcKx
ns+9XjJtANA1TEl6hldWRZpExcZ2jH8osP9LbsnCCbJgN7RiZ/SBUbHR7aFmcNW7
sxnxay7vUKI7We47vdIvSI36CbWmyvC78bfS3cDLGAiyoZbaLrLcMrbjQPVBDKAd
JowxRZ+gZ/srhBycDP1Pem6bn8smG57U6O42dVlRJweT2ri06jIkVS+1JAyj7pYl
u9LBWSoYYVyVbWJnYAbM/cQXdLd6uI+zHdR9+k+83TRaJJi4W1qYEZrfj7hcePfN
c8L7rs3G9CPw9Y8FeF8QzAP2KC037ND6LmG0QXi2+pwkm52r+Svscmz5MnE1fHZb
gdWqwTlU6q05Md9SPHTZDGDrTeHhjTLNeXoeMDVxEgsJok2qb9PcLhe9usHBgEOi
pBu7hwN91ivx/yiKM7vmhyYTP0eFcj3kuCiuyxNxWI/fkx5emHyrjvc3o0aUIer8
OMKktqYcGhR1p3ScWYnM5VdAbtX3m/0uedk58h0z+cJc+3mtkSNXes1PZjappysl
KAjaPubSVC56Xbw2s3n/6U3g9Xdjfd9S1biAoouK2quhL3oZDxGNnTd0pwcdiG7F
0wse3Ynu2ycYMmbcGaJSYZFuN6qJGWhPBHPLUC/xNuOkktmAvz4hZAEaJUHIrkK2
V2XaoEwqBcbt7QifiT0N6R0LUFF5yLhv7mcx4g0d1Jfcc5ibHMLg27Xfs9OB9NlM
PF/aB3kfCRJIfXTgYpms2B43GQEDZcljR9uYZZhnxPGXoCMDju8UmL26DPS5QmdL
6NnLHYlcbvOcrDvIzM25L/7scnv+rRI9Offdl1YupsCADYvDziPPfZ28RekGYGc4
4b1yQ3fs47UbophL6lpoX1E3yP2D5m+6Eo9Vy0zkMzmV096ZL3f7Nmbvm9EB4ApU
/dhzLcTEQi44k3ZnFWCVPru1gF4ETWp+HmZxcXkGhLs7/hmLHfx6pAs9x6sDG/Hh
NMuGt6eT8CyAoNB78XzlKi3SdTkCTP7w45ICGFvqG14tPbDQl0AJrwyF36aXdrBs
pqtnBMvFY//Ym67w1RWzQv8hnDBnNfZ4CGEbezpVRJ1A3HE4Zpn8GX2mfjhjVeo5
AJwPVnniLrN0fyUoB3COebeQ9X+CIyi7FZuGVWI+Gbk4nmFrOOjPLb4UjOU4TWRT
Rwd/AwDwOoz2mQiUq90nGSFhbwr+2gNilBBlBSmpQZ7ah0ahE2j2tfTqBinnrrME
s9oYXenRvCfLS6IQs1m/jR+2l6WeuQYzi1un03dpO5lnVxBHtuOSDa2DK3acfj9U
9PSq/60j4u4BBX6RcOZ1tU6hkyZwP+ARUzb7uwrIJyrlZtz8/UiIiiX/wZhtisY6
Ik6Wlo4aw7+4844JdffCbTzvlWyYO04WBVh7EDUpUDLDdnLanspAiomAwbj9yNaY
iOr0qqgFYAV8VOseg5Y9B6p8XLgZmNuV28p7wmvU8UMYL8QJgMzahDq9Ds8rFBgA
CdTbWgsbdmBQHR8V7asWfQC+P8bTLJNKy/JLPRli0f2mjCGFx8osjyXmGhQVZdwC
zyWPkg3SjV0uepJiGnWuep3jsP/mNXxemKsPc4Bk7UQw04m9+Nf9mHRaLTXazOGl
IsAGmiNyOzwjZiIZucz1OuI4+CNYtlXiiPFuzpYcl4BR+pbCtktnWNFWvg3FqoyL
4bFDEwPpbu0bD82m0MA+JxAykJNm9g1oKFJ6mO8SFHXwNYeD5wk1k8GZf69KgIGA
9UvVRu8a+oUqiS3Q4KtNTteXve8mel6eTbqVo0Ke5n6Z8A+/vpGVV5pxe7zgnz8T
hXPd17o0xxQ8l0JGZ3riF/n3DkUyCj31kAGkFfglzQ8jB70ubty5pXXCnG1gUFJf
ug5Rvse83r5b1bnjITILIMP45jcdrbFrAbO/eEBw1UN1Ku5i7s5uCQUIOOURvGKo
6bzrCDHUjJPUT5k5EorEZpeWP71dZBFuqDfbxArjNssLlnzRftisNQZWAZaVVZSu
6oGyA+5KcNe9hJFkaHr8qyiLyg12JDQqNj7LZH+v6/DwH6Wv0v8APawX3fJyvQ4M
4VJ4dHYb1r32NHlD3YKVM+ykUGV41HDkXrt7Dj2uY0B5HahLpEmsHjNvBhkgPzfl
R46LI575bnUQs9lqLCM/HjMOGVRTWv0f+lN6LQ9m7V7RDANhKchoAiJTSgoTsE7J
kj35z6uJgykK8faYN5foZl9GtIpMDoyT8WE01MBwuD5ILwNfzMm6iU1Cp1JLK9Uk
adY+fQB8DM6WJGB3+8CFJJbnTKbO+66I1hlOfha8RXsVzoAEEOit5f31W2O2dC27
VNtmf2b4xJ8K9NS/ybm7iXWAMHM4opI+dXHeIeM9wE76Os+VL2fFc0hZw0zR29Ei
JVjuq1dboCmo+nulPtvu515iD7OiTkY21cpApZACnJv2T2lLWITyGHll5C9kIawQ
Oobvz+iXa2XXnW9Spv6hx8RoZDjJ70ldsJA5yfApCblHE3FDYZ3rRaOu9h9Zcujx
xFy4vPu6ei+RNr3wR7X0k3XKBQAmI5TWW3j6Q6dUmmNM7Gc5uj/Ru3ASi0XiJ1hI
BgdCw4Gi4htZ2kiLnO/a+fSK5HYbAh0OP1vqSoWvZ9lHnBkgPWNX7l0vfO3iin7m
YPTVwCHord4Aadxa41nUIkXbzqmFMETrv7oP7c8jXPvlvbvObl07W5T4CMazaRq9
1Ti8sUNk7OUlSWgb0orQMSw4yUuU6wBxGCq56f2+VDQw9THA79jE55xVEnjtiGp1
F01X7St5+pOU1hU1n6+Zaxhjgjuuwh1tApgR3s9OHHQ+YYT4W9fbOSXL2GmspBRe
Gu9MumY7l+hL7lS8QfCDRTtmCz5hWyXxTz+LpsprusmpF9+YrpAl9XAg2JtdtdYk
ZCVJEIEr32gLej4ux0Qa71ewYuCKimaBb6GJ0Lr7v5MC6Ccj8TpeohXSQsWwuYFW
ag5ofJSKLih5MVXAZ7hSigfEDzQgEEdX7JkrGr0pyAq2RyvDOtGT1ZE0KqvwWP5m
Uh1hzaXzJWqmDgoqGJt22wJJQSAm9tOT9vM1/K5cvoEdX2XKp6WQhoqr3ZsHlX+f
kPGq6clElCjlZSz6UWYZ3wo5R8wd8MGdzRLNVK9t2f/KXj30OYtDD1CeHSzkUaNz
cdF3Lse2BbNnxQ+UImL1ZKL0bTZB77WBGCiLIZTQcD7iMUWk5cC+2JIKYAlm61Kg
M2MB43zM6J6O4+zz1NGBxx//VddIyMsigk/GR2BwLC8I9Qe0Z4AzataMaw1MqE6j
6k/OtaZoY3BcKg3t0kdgqA5MgKCiV2abKcppmmcngGYg8BeSYCXNeMXDpbd+9fZV
EWy2ylxhdrAXZEgSx8WDe8YKjHTaaWOi/10cfqAaFTB6CkkD3EK2BeueLCP1/fQc
LphhN7wRMVTciSb3VkpZUDjZ5S9VZzHRpR1lVIXcy1kryJJ0EnD5jPQcGJz6e2Rj
ZzKO0ofKqJHUZZ2FdKNdgpAnXj2umargvwItHCLsAjnSYopw6fMJp40zQJcZ8U1F
R2JjfxZIS306JUeAR4wwHT5HRdS8vTjJdhZ0WWswylQuwwE6JLZNf6n2G5bMBuyu
N+SE2zCdAhfhZcCgt5t3PAGUqIP8am3hmkErsYzm1yZr9k9hFUWsst+kY2UuDs/9
+sFPlImrGybdFpqPx5FU3zOrzCme639Z6uqCf9yw5C1kHX+5qGYJqoqj+7hu4tcA
7wj30anwcnU0OEZqoU37d5H+2NlCkvhnH2Qc5IgwauEIWkVBTnzBxP1Mn49vP7On
elUKisyWvbc1x48s/9+9itxCoPUniZrvsOiTLmiRzmW4h6/nnS83XgKfRZj6cvbF
+hRf3gSdsRlSoLW0Q+OHd1S0aJYqfPzq/TkdW2Xp0U2EKQRTz1Z959pwLjoeFpR8
kE3mz2Gce4ZEZGuzAnIXEG8jc1UkjKhY/uPLjPeo3Gf+kyyYLQ/aCkg1EXZ+Azug
4hvDtpXsOxQAtsCfvOgZZ43YsR5vVATHUpY7M22/ErEDV7Jezg30trtrE0YzXDeF
Le+XmJjSp481bVf/KqhUBtE8hs8xOtKHPZlSt6VFbO+j/gUC94bspbl1MXwtZMXA
egumwud7uFNqejcL4n9gR1XaCEh0IRYMHpS/EHt3wOJXq7K59Pyx/Tj9uMYbe/fn
Vzzw5PKHBIWPa4sMAHAgisi/WMkxuwhaJMlGNBgiigtvPqRDJdRHSGV/9VHmRnNu
3OYfdBSJAh5YjJBilHDaudFSshMhOjTX3xHQvgwowxoYBb+2qgYmnUwZAZ/yOwrS
8X79W7gFqz/t5J2+d2bSSlhtIobPGVMXDNQMXT/snVNOvzZlXZM141VDAfznJniY
yn8FaVSvU7t+tR0UFX+27Sk44m9ukoLJX8mW0Pr4RUYEcB02SHzMRYE9qfu0uVok
K5uukJOSL0Dp40TOabr+1gSmpjwNzlDkRxgBZfByxdiwHnJC5osKfjgm2cTnogkA
pDehUUbTKgjrcLYMHDWUSFLUlmSLZs/q+M8mwEr39Xol8S3o5YMyd2sSmnejRhCu
4Vnd13B8itQxSZij8QF5VR9k1+uz60vAdckD9pa/TJXsl/pGiZ33+4YaiXjCTLb4
Bvu2WO7ABm15qAmNa4yBodFzQfiavypOk79J01fHOoznL3aOxhLLJeNroQLixvVJ
dj9CZ01K7+Tsj9IIgw1ORMi/rbP4AonX5jzruuQza2f1LS2fTiMamNxYyFx+0/F6
rL2PcYeEhfVJvTkh0indZrSVgsV28PlHugEBTGKvMuxkWjJoyzFwI2yR3BGAl+ky
7as+YdG66mrVDfmwBrJnf1Dhfy3uy8yvXzDNLM8gs4eyAbWsJ/1zZ/sXpHKV7cRc
9tU6F1uJQM7+j1YuYu7GiradN3xwgs+wIclfdS8RNhQNYL3YXsbb0hn+gynISSgu
4xtXS3jMV8dqglMRcsiCiPeElgKYCTlEk2svnGORljovK1FHgp76jeg9nu2JEany
uGD/yAY/AvfAGk34PobtnO0FmeAp8cIczGhf/d31E/F8hofWlMB1N/O0BKPd5iT+
SItOoYg+VaAOe+y7CeuqeML5UFOKNj9TcQa6gnA0TUmSU9w91lg7RK5Am9jTB+qQ
TqslkK48fY0tScDJtW4fmq+TFZEsloFk22K/LO52/tbEwgDkLDwBK+//NGICtp4r
YgWe95H685bvR5XOFGb9ASfMi1jTkxWys59eKe6ichR6NCLkHJCEdx01CSt76nU2
X2zQAFYhGm+OwXLjbxci5o1uBxnTnEeIMXW63OFkiyIrSkn0P4vTWt38vBm8aZQw
33NesuLOeqXg9EyxEqQjK7DhtMxcMNFeazAAa+9k5usg2iitAxGkh8A6woelslfr
pi/w0eHWJoUsULkcaB3Hv6gNjiaZvkzkRS76cv396BktX913mv8ZA1sCT6GwzPCV
ni65/Off5yp8W8YJIsh1zPgfTjK9KTd0krJr1A94+8mbk/ZFX2qDn7Qsmr/ElEM2
Gef6xqzqGPK2b7Lc6vluGBGVkNyaXbWb5lSRI0tB17BUOTkboGHjp2FrxQsL6IVN
dqaVZgFEkcgd2fukK3cqKIcCbOkfjxmizcv2oryMA/dWwa9a4+qsuexl3bua8/60
8aIylYGTFJ5YvHqor0R2A40hAjJQVua7Hg7qhMzbiU7Z/CCVAak5DoDR6FuRo48e
Y+CIBZ9NidSXAjiOQNM1xqCzotNJIcEHoFmCqLF6mdAy08I19wNYUgj7F7vxhKu0
aUaRYjLw3qmcTAmEihr/rxuTkOVH+MHFNLlx0U7siDyc5qlN2h+GIJHV5+D2bdr4
GEunuT9wZHYCywnb/XI2zKm7JvSoFxz+XUWsfHn/8KVNTomBiNvhtPFIeucmU0sR
mQmxIgIgKgZymJ/ZbkZgJKrLID4gNhNcr4GFnMBrNLguap9zmpAvfI3J6itYXQmx
kXwH7HIN+F5U5iAKJgNquywDp5wK6QLWHuC7BWd8Iri8QDvRVdD91W8003rx4EX8
O/ncZj7O7xQLs4gefCvGy/8Q43M6QYN9S0noyYa6K0iW465NMuIOAdNasgaw5osL
flpmWhjUeMVtak1uBFTIZzfm14M2TK9JZQG2tOloIk4AjXLp1D405MHPyGRtU9H3
Ab+6RwM/M2nQ/fCT5SL5aZYn0VHMFLiq8PZX52W5DNCZ0QsmZ72vtNIHGFgBYvUr
hCT5GDm4yXKYSso25IwgXL7l08HbG271RnBRH1ntL3QzwOlWgRHuBitgrS+Q0uZc
uufhYt3HlJeE5DX4KrxKh05zr3N7jkwT0yUCpECzlrmkZSeWDh8uBjrlB5SDvXLp
v94Ii7SYQUAyGp3zPJmdzNqikn09jHdqUe+99D/UeZV+3wXkIsOzANAYGn2brqmd
kOhq4R8PlzyeqA8oGg9F4Gu8giX3NiS93QL8yjV7/DmM4CdYL6syG7ygjmyroBk6
jMo/zaWRSp8jZ5wy9tezNsDy+8jq2i/Sj4MpNt7tHCEw57RpbtKG3BVzzux5TBNQ
X2xZSq8W1UQ1jAO2NDgIZOK9G/X/hDABAD6TMlXeuse8ToNaJH2+1ZBWIXHhV/84
gjGmt9D+5gQo67Y4VMB5oWFa4kPBrhKRMKlHEXrOBI/3kaEy5YYP3hMPPW4VEJMT
G4a2N/dEQ7dsXhEKh6pn7Py6SVduuVw+WXFwJFOTQ6Qo8gEPMh+wIB33o1G2E4hg
QKRUBySLUsDCH3sZh42d7HOKz2vEyNZca5rDmWJrckeL5Dk+1WO4+16wVgMqcZbD
N8EX214GtVkAQ4WAknApWYd83L5Ja5K58gs+Qx/bZBRfBNz2Cs6uBgz2nE2LSRAc
xjxELCOOWML3DBuY2oVguYK3ZDk9dQPS3AlMD5bNHMLso7h1YiYS5GG8xMFbZ6M9
UwuD3I93PTE234c144u7nA/C/CuKj5Hgmk6lTF7H8TgHtxu/vGzqGpQRYLXR0vlZ
wJO+mSbaNtIOwlLEwEj6zVOJE2adDt7JLCkQTtGsKlSD5KvpkYHLNEO+61aKKbfy
dmXocKAaP2IZy0bS50rbTXDEnw0vtI6UL2fxsZAmDAQ7OqWBafCTl1GoKTl9ytxB
xJdzJR35C1HjyB2PMZqbE5u9TE9j4mtMV1gbsS5PzTi2QEJbbIIQGnT2nWNo8wcO
kS1k4pb1vQk3vUqeDh9dMmEAAMebAS71vSotzlTDQH5cmFUeDQdQYyZtLPaL96Cr
baCzF5Eknm8bqdBolXV+gLQS+Q7f+USI+QPC+EY9onRjDgOlbKdGGP7RKJCcqdDA
/vCVbHD7qaKUnts2TCWz5NfGYpXZDXuXvmNm88+9ulOUbTyBFkx5wYILEmz5AZsO
aV0yWGlZoy+CafbIbgw6MbRb28NqVLZqAKAZtkVAolkerZZV4xx6qfOa9BXWpPmC
rF8CnE+nxBDDsZhHWhBNY/XnvSOM5L6ziT5mwm3kDORxdNQ3/tgDy0i6P4WXeP7w
DAyTKVWljbPHCNciO4O4V/b5eqTCTddToKvhgIqRqo9Q7Ce0H7Sdy0dAzUO7Hhv5
7nqh45XDxN+BjrSjrYuYahTPR0IoY2Zff8HsfVGqVAnxuOre+Qv5Z71ciC8O4Qt8
Ap72akoo7xcELWZSnP2yHRVKQl09RFJ1/HhSso0Mo8qtt8ZHBh51nnT4YrYIem+A
opRLbaGLIHENWDqWMgKIDJOpQBsWbOPuIzCW6s4adTd/Lnr9dmjWvIlP68ubXVP2
mjZCsCFUUx1wxVIxJFphBvb4nmzz+ptdhbJZdEdpmjmnIKF5CZPfQyQ9iBbRpvLb
3gu0qivihUokTyI6XXDcD7A5LouJvy5inK2RN9ZS5mum4Z4qS3oZslA4AAQTPh+N
oxMsZ9JYNtZEps2tY6pfgTMNBNp7w6UACTSxxT1u39dVMKBZ38YCs8Vq4FDxg621
OlCKhTnu2kTnWB0k9tbED+pYuWGNDFW+gwwkC7UO1ATqo2O19v2BdPt+7VBIsB9T
k6ChLcnAoZGbcPLkiRGyI+GAEKBrUBFJFqHkjcrcZZCgZDcDZe32gn3IFwD2kuQb
3mCP4OjDwal4R4n/RR6AVB2/0ryygRk1HYubbNGUgQEnnU+QyrZoxYhXkX8Bir5L
yNo4QgohyTlPfwqpDZCaUTdmLkn8nq0iceV4Nliynee+ndf0U2zcCMh6YMbv45OE
Ut0rSAMF48WFp0gLyqBhRNztLFH7xE0gh5G91nnchPzEtf13ZhJHLZiMXQVMRaZg
SObuttbBKXAeGs6QhJ1dAvIvvf2H42aNOKM425QWlp2k2EDX9z8BAMuQwXRO5iq8
cPeiA76o9VTwRu4Sa3doZfRlz6K38Tnmti4FbSD1+a1qQSzv8gL0jOMfYb1NVWXP
ZJiTUdV5bCyAXlkdtR82JDruWJjixADzBa+njyTHsBlSo4xvxssdUtJ1yjW29FqP
hrVn1bprZCN5lum7Z9mqaOubmNNTpKENPIe6jTDuboxdPlysQAgDJzWrOu3QN6V/
8X8TFKeVsvWkiPcPaQP49Ew3NVRK6/YxgKb1XXLjnieVzuLrY2leoeWqOLKwKf6Y
iC5R7ydHi3yaH+H9uFJpSLL9532YFcdcsykxZdIkY0S9xpLWaN95BedjXL4PFVLX
inykPW9BdZYbyfk0HqneIS77bkpzhllDXChaj8v/8gufjluggjXu+zFDKqwlx/8H
E1ebjmwtI0UN8MUqr75cHaSfMh8Ya2sls84XjpYhuty9621uCS6CICLcxAjo1zXg
2bHB6zpwbL+Z4lnL55P7E6wl+v+XXJMQiZwr8CPX3uJYbaBAvV+pX2uVyrvxgK3s
Im2nEgmSKzKBodd+lWTHBonYAucadGKGkyD0knzcXp8xnveVTlDHBmmugWrVZxbH
VisTHGdEPOBjCh6HEq6Xb3VoG2IgY2VexvdivxQyZxPrXV2THEjgpO/uhXzcsJa5
C20UgKuNjjjtq7R3ZS56ZZ3Ce1i937Cl4HFwxC+9XAuUox0MzhGAjltsFeKslb93
48Cwa44ZUaae6W51zBhHuse80TIz+QTx3mFhQjJ9vqo561ajWBVfznt0OjaMu4Hw
jASwF2sMSjUcjJeX2ZmT9rAj7HT1a4j5jO7GUV8BpLF7K7zYCLC2BX0KQ7TCouBL
VaTFNnCuUjIcoHzQwJZimd0uBMt5f7etiJTAW2tLgil2JhfQdxIgO8muTLlwN94i
Ahyc8B90EGJksQkpQSHAI39T5/EZImtPOCp255aL6zqhFhd+y+q13SZIYK3U95N3
Kq7QHDZ6gMFYpnDUMwAe9wM3VjMT7hICsKj7+MX0HIV5g4rUt+/DtfOMCr7MkYiN
GhjQCFa9OUoUeNI1AnvcM7gnueB0ssVtRfrdms6issLj8w4d+tsttYsJj+nsnYz4
PmeSWc7BRr31+dVx2N+vQP54sem43kuNYBS1N3yDXuMFea1C8daDMWidXP400zuX
CNxlpvb3jL8vil1q9iB5WfpXTazW2NeT7xRSI0yZavW1iXnvSWe3bdkux19DinJ3
7XiJVLP4vfbksdwhhtoNrJlU0r+ll+S4bgCNOrKCCjBKAT+LfROlkxFKDHa0FOCY
7k82JRbuwOI56iInMOTNF2BKz3HDgl//Wb8NS9t6S1+RhIRe4PeUt9h6CaHBseLT
qLyPcnPCboHP92RgMq0zBi/HN9tW3dj+4YnAS5n9RIUsQ3R/Jn81onPKnXPjJa4k
ID+bEHogzkw3vtwJpQSq5ocZKeN1PUS3kcshPQIh5wWLz7AVY4qq+bpC6OYjqTxU
qMCgqNujR+mp64zcLxoxl/01ZBxFOeB0LQX3CzPWuqMa/cV4wygKyiIN6wjaj/2a
f2XoxtLK5KnCNZLVPS3aRpuBvg56qjFqMbQ+OG8KLJcszWDsFo2ar4tEvU7WOgZ6
/gSK2a+cEtv4Y/EjpMPhrOHLOGPNt16v619bOzy2q2FjyFueL7aFLS7rXbR5gEo5
pSu1y26D59xec9E+xCJy+iqqXo9whh42vWo4ZdYK4PdP9VulO9hQXaVzJBvoknau
2mJkBiojLKuks7igsXWowkjPR5ruWOz4jOs8Xr/ZWl1qvBKxsKBZx0HCK+c9OPEX
2FvdAYtoq5RutQU9Oe88E/CW/6WwAIlqAaYrN+3UcH4j0bwyK6P9mxHfAMpNkK5N
0berQtPY5F88gIdNUk+D2GTyUV34rX8mEAPR9gcob2yEjE80/uoQhmNj4R7uPrd5
FF5HgbCSznXTieMFL+MKmgpbt4DpwGnhBmp8GQ/JzLEZ4G5svY0WUBhfNcK3n73o
xksJFS1/5FUKqEomtrCK6b8VCNESXL6tQSABGNN9zvgGNEgNXN1FvCgdYRe2yFTB
K5fXUfNlMuzgmol6GhINNffD8otx3geEMMxZkkLXm2/1sMWqS3Y+eMbVk47Jegc1
8CaF6ml0LBIWk8R4965zDxZZriPKswVwSrcG84d01lZuowLS8A0p3gDdSttEMoyJ
YPvoATTuZUAPudO8HafncqDIOE0vKJhfIcUN9mgyaigZQW9+Q4XkBy4CKYrujwH+
68TBzrUhxLrHqDd6icMZIIK7cdtT2p/Ybe4OaW8tuaaRFmzMrL90jPG3Y2DsrCBs
M0OvwwXYP6jfIho86oHS3yMPUnZNKgNf5PiI8wIlanqTmA8Yw5NbsKYD7ARclZbv
AyFDlzZaYfeJeZtBzrybYKPae5crK5Tq79lT+1WuOX14ynOSMDJaivpDeI/qEEnC
Wi+/xt3l8mDlC4rIcVQ4oKBGDKlkPRqq7jBgTK2a9PLfO+rOU+3bS9DPOHYw0MYI
sH+i0hkVUf7griI2lnFE4wHhH6q4BlNGYfg6TlGAbMnu8MkmZf+JWnz7fQiBR5+c
0rxK7AOCFSeSJgKFMlgkY525OW+D1WbYnxwHOEbhh7kmFuClCUyVY6/QGAcR+wwA
6xVxBkRfs2cOv1/gSiG6BKgSq4jNM1GWH1TWz9q6Q7SZvLe6PJVLrE3OusNm4h+j
dXWbkAkMBr41r1bl3CCC8yRb/0FPBX0vjd6+bMr4KVJg/IC2UpYxs4zlyqjoBzpj
55PjiYBW8DMYE1hs3wp0GVsSso7COo6lTxFR+Rw07XhxV86bvpmv8Uflpu1z0O4/
/74sNF6ysBb/f5kYVNMg4hh19RAJnokpCUJZ/Xj/AgxxlTpalDN/hOOo0ggK/I71
qrtukCOA3Ockv+/uxao8OaOKgj8a6o76ev//1T+bOFR3wbL3JtlJvWc0ksxSbgoi
Pu0xIoyIgaqKy6cbtIxVW7pL+lPkmH6qrwVbBIvOmdNmaRVKwD7X1UBp+XoQDhsa
td+GdNhECWRvUTjUnDFVeUFnLa1lRS8vvpNBRrbEepmq95+EVVeYmycViAmtrEmH
Zr+tT39LdMCGen3At2KaAIDHOVaAe1KDBySgOyRkYzkNuQLjTT8AgAEZGspg6RQ5
zIOPz5Xa2YxC4v+23p22CF/2iqaclC4pk3bNvnLhHzmccPEks6d0vdVf8+ZPy5CI
MOndzIkjD+JI/21nTmMo7dS3hUpXYo/eyoNaoU3nAYyQIfmHT/9dvJL5UOKJ4x50
GHXRMmIoFf8BwEgJzN8MqBosrWPnG338ynfkgvSaAV7lQ7OXmg4GKRzXaL+j+k5m
5SQKqK9Kb3N9CcFWNTZOEqecigBfdYyL5HWyFC5Jk6BbT5s8EPrygAEc0eHS4t3Z
ziMAIvisD1NHGfSzetzJbpleq4dE/mPw6+xv4BDqFZnRVsvP1k5fIWa537ihieDp
/E4WiyUA0fvrDKRcMLeIzQT1NMlvahBg/uPiIBBT99+T0YjGuUDOXhp9EOMFQJx5
36ssUe4i0roD3vuukmwIoBMnjqSpueQ9Fx3oqhYDEOFkzSvn3ivgRtXvD6bQjirb
eyuy3eOgcjbWHfvu/PCTuV4apArXaHvWJney529eHsj4N1M+ct784q7J/rT3s4L1
6dfCav+TKdJw69lDu6sjFv2iAMVx+hoFULY9CGI1+W9dRDDD0G+s9rj36Mk/Mvz1
yZVwEEhFjyJDxuXaFV6OWc8wfpvcLAEbI4WimoB3MscfSOkMAUb0DA6vBwhO/hJv
VGgkQ1RPfPBQ3t2+E232+ya9QVavTiUOhlWfwtHT8vkpEebNbGEr/izBKZDzrUMI
EF0UsB+dpcf5pf5Qwq3OywJeJOz3mSDFnRkLvdRu/TCwoEcLTRGKns+vul57xCnJ
/MJ6s/11SxP/MY/hkc3UUEK36UIhQxnT6Bpl7hpOvJ6M3eZOo9PxQ5S7pcV5Td5a
Aor48ZqnAgHxFeS+y1BhOydj9c7VKsgrVkGThWrsIZVAKuax3X3Fa6HU64q0OuGx
P7fm32FkW7gk6ZnwzrNQciBe2ECXes8MOlx3A20bD8lLp2nEeZ37Z8/v+9c0fEkO
PimPgcU5pGre5GpWuPrMkGfI8Rmb5GNoxfxUXmbwt+4cCK0MgEEkSiE+xvcoKx0W
c9P27tlm8HG9BGgnyhgX+t2eZ6w4+Eu33Zy+3EZFsKayvIPcTXmRKRh61ZlxBlqz
TK6S9IAsOeZxvPFE/aEzWvHHuXUA8e8G7FJC4h4bVytIV+ciG9tbDGTZngTJVvoJ
TRnczOTxdQzX+se90UCVqpdy8Qdh2HQUx3J/JpjjEbnfYACsT93aj1AdSEAU3VlL
Zc5tq5XoVXnGfxxJM+Gsk8YwVA6TyMDGmf0dvHmIOMkryAD2nzDQfkaMF/6lR6Ln
5KCULPdUkRzxYfegICSp3XQWE3+8an9hk015E6IHcOmvSD8iK6akDVHYONjixtVR
7VNutCKJuo6AWHuOpP/tF3awSdeWCgbJSd8A6UAIS1AENkXRIutAWB5P4k+23QXg
VA9Vv6n/PaYKzX/BZ1ewLF3sEtOgmN6/neWGGdpQp1XHSQM03i6dOFLmOCMyWhm0
lUhImhfqn4KL40EpSXnCbV3FLAE2cqMTqoh4jHtzA7blyGty+rGSkG6oZuYAqLjb
8gv0B0T/cvq7BUoIDwUq7F3B+jOx1X65L7HR5mh+/+Ilb7GtfLI6rJl+lXschP43
njIr5kc9CA/Bw+Eb4YoVwaeJV4Gb/WYIdcroa836+faIMqlI4sL/rHxrhfgCRbip
DigRjUukLKFGFHGsGxhDncO1gt6dwH8aXU+dYkctuLXZea/n/4pLBaAFWUSKTleb
38J5Oxbr+69l2BJf6vIqTf2XSNsOXEwpKdUw3Y8J39RckpYtsPkb+rE9JrpDdiWC
0bWv3uk0+PA1wXvFd871FdI7dbFR/RVnSukisBom6auWf8G+LfJYXQWAM0FRIfnS
hvZEJVdzyELzp6CIyKIDQ4RBVglQ7opJIKdIovJztteQ6hK0k5AeNuqwJXlUwccT
aBWNLW/I4xpX1ERA8FJ4znGfNqFgAlgFAPFWWZ+3rnIVkoLTyWdr+pxwOZJuo8w3
0NAoz3Gi7eL18eVUmr/lE6M/3tPV+tnnA3Inj5sBe45CC8x/xYmQ8zdwWowAXjOq
K7x+5oImVqYAFu0J8VQSc3YR21jTbPzFX+VzzvsPrSuDi1W88ohCESuw0TtcOG5P
kkoHxklPI9BjKi8wBvsYbKyOvja6BZxW7jD/s/Xoe/bimnBqjEsbM20IdEvUIK4M
BZ3/1Nnc/cx/UKlYNDoRyfsQKMgpnIpXeM8rZl/VmTLTQPVfs8E9O8bpfWTUOyMD
GedhC0VO9gtPqAuQCPdX5e4E2o6FxCO2WKyNx/o3dy38GmXWUjwEFQduFeV7w/Kg
Otsg0h68Edxn/v8vjnRqeEPrRlBycLPqDE6vmzQAHsX1FGli58fjcvl2bNX0gvZR
ylu5Vxe+8/7YEabPif4McZGBfFYT766U6NDLHQhimyF2KZaRtb9b3bO/LYN8Qh9l
SBSuBiXtO7wJr01083OSBeIXQAKBuM2Ey/eFOkN9WxsTA+LPd652G/DhbeS/n3Ff
oH2QJwyEtpEYfH+hF4Pza6rpWDXITVK/4qlBEqaln0MQrJZPzu8lDyMkrHCYtuSG
0MsLg9nhX6sqx0ZpYZSfCgJ+8sp2o0o4c7/er7gAL7QeSZEJOD/0RaItXEwNTKi0
z6qirkegIeL1CnUf9mt/YkjE9xhJuOThZBdHLdsn+y+UYgZZ5z/flZHCPssIM2hM
YJqV3BOYNE8+p+HXdrjl0XxPib6eHwwx3JvTo4gjH0dXoMv7d8ez6mQW+LEgfWp4
Q0X0/arkqe3l0YzpklZuC0FuYmWLuDhvpoQwJbk1VVmr3/jvW3Y+RIF89dh4FfCX
ysIlcKD/ietx1fuOjQTw8SsMU1ekkzrUc/YCkmav4Og74+7WthnM+4VpvVmMSQxn
pLt1rjh1gqj567fRBYF42Txvfe3oPQ73xoSEtglr9BtXVtJU8GTQoZLMie7gmzPM
VJ4UmjutuKahcj7BDHGXi71KEEOqc6jhYwhriqm7XTYS90mRH7Z2waluFTdYKNJb
aGkr9MGaqRhYYlP1l0C1BKbvC3kq/WKY0H/BUeeT/SRRNuMdaprnXwa1mrd3CJga
gDKDMu7IMtWrvyutIRAfuOsH4IlNXLuZeMI3nX2fpgxK9uANGyoVEeakiPBvEOnE
TE5xzQ+tss0M8ID6tQcGPr7iocnpkktp6QyqiIkVg1JsmvGJEpRWDzvrk5WtZQzv
3QLiM1mXthCSQEnYJSZEy7/P5n3nbt+/iP5smV7d3L4bM4MVEmmNXRnEjR+AS1qQ
m84GYVV/QIR9WuxGUAlrAmeyNmLJWcU9lcc1j+aBSn2Lj7rma1bbPgjIbuLRvpMn
AjrnGM/NBD9TbC/B0EMfFu5IUdSd5mSYmSLxNrHZcrMzf5rhsBDH7AFhpeVfE3TZ
dcdUChUoKBKBgE8/ZsT5W6navRyqwM+XJKaDgv6J9ppXyle7NzIDVIBhFj/2zYeY
rBQOKXvTKh4tcg0EmDgxH4vRiPwnI6GyY16p+skMtKrXlkZJetGALaOp2Ka2SWnO
yl/tyempkwhHpyroSr+z8Xibg5oi3c+myR3oGGESpqySP0rf41DZv11KOTmmw5bK
YW61ApNld/KrGeWOV1qvPRV3WrCr+htliT7Zey5PVTq7fwGXmQVI8eGkzikw+XcP
WYIN7S5tgcE9wgkXNoL4Km+3RhLX7h7QN+hdzgP5fU2pa4vn7fbQoWSosI2VkBkC
JK0w/pxjRbSqWYtuhs6TIq9beYR4xxH07ksswx8PILa+bN3DC6gV/MxLdcVXulF1
xbPHO1izKXtucaDFe66Pha6h0HBzmeIOrFqbPF+UQQvNTCcSejjWwrWknorkZweG
nzCtpUQ5QP84tOg9RIkjP4QOHGKc7BZbqTdPzKal5zda4B/aqb9ekVyVn7iJ/e6z
PjdgT0kuNf1LAvcIDMBicyHtnQCqhcegBcXpCxYI3ROtqo2mdnbr874LbdUJvAWw
M8heTjs5VNyC+5QVqYnaYIYUBFpH0WuvlhykJzglp+MfOCZKKhUp3helr9mXzjUo
Pba6GrwahkrMEM6mDFOZU12hFD6QYrQw4coaj+7EvKm3eH3t1bWzXLzb0Ba3AIp5
zYQ1m0xj2IW4f+7scftd3QG05Tp/RTlTYLAYXJEPW/HnSIB4UsznxVtR42I+tV5C
CJPFOaCZ+1GbFCSOq+A5NVWnocU/JPHQBZbJQsXMpKRb2SwBGe+BYSbcnQl+QDn+
/iFH9XyaLgESZUwMc7BamUuPRi5OOdkKVQ5e7eqFquEfTfpnud0D/MITFC0iDL3P
ZNyYKBWzxE0K5eIQAJ+g69l8PCbyqLwC0G5UWr6Fl+mW26x9cgm9gj4NrezdQod6
EN2cWJu4VAVYWTvZ7yvcDl5T7rW28bRyUnE3D+E81A+a5XjtPAHrXzNjsO5JeEvZ
TW8I/gVH6h/Iv0YC1N1lV5ED0A3XXpXm05RaucFjoqpxmEkZzOlTPfOb1hNpypCd
+OllewVxJmRilI5mACRceKl3LcoQWJIJnNxZ3qfNA55xqY1DI408AObYCQKDPA/r
5yXOJtaCyQX7KvAyDfNMzAazifmBcDJ11mCgGbZyxHcUKjI4Iv7jmd8r9CJB20Xd
UnuSl4uDhv99GDGsSH4l8oi3Iw+dTp/8sel4SL8pZ2F1uS//Gd6v9H88829lMKWD
WOUjqrqJHhRFWmba/tBfd7XoxRVt/sSrGKlLQCszs0pW2zQRsPqOxiXwI4YG3F6A
19dOvqKEaI+puUmnEzuUDqks2JHTQ79Y3hA90zzMW9cy7QibcqqzSpfvpbNn3X07
NT95v/mUbYuM+Iao25eFdln4nMpcWstC25zBwGe56S6Z4lXVV/dhpmUDIiFD8NDn
BVP95CP53yKiGG30BOKQfLBgGY2vmUVYUnXMy06/Crtk1h3j6MSF4K77OThG+pHx
ASkVJ4cu3SI1b8X4nOsJZ5nFtYG8KLKuE3gwg/utQeuILYPgdBRTsPpxhhpjeT0/
XUZkZ8KNSXcM52h0Q/UTIyskvBeD35vJwxqeUT3rN/ewgIRsILT6sRtBFxpeXk2p
2VPqN/Gj1pKVitZ7RbgAbfjECCUP0GckHkghsHt0bVTufC9yc4kVR/IVax/n7xqj
Qp+2hnLBmnKvFx+MjgIYDhN0UTc+jtZ7qET7Ogibq0KJr5yaH+z0+Gn0/f+jg4vu
QRJNaRV9HZt7ps+W1R67+qugoh9SyliWizO5L3+4XwVec4qu3Gh7XiQ1aiOiwFco
Lq43/lAccpXwya+mBOI+E4UYzQk/yc5ngsH0bXRAq5tHoBExur9xFrlTWe+TZ40a
9enwoAzGidd0zfvMNhX2vnjDxhKvskMKTBUubURs6JrHBR/XWpvHEKyYnX7Pq6Se
ss9QD4bPuvHZQvINpjybeZkt2gw+XTO7/YvMftNc3vYF1neLW1moxgKyZiBDn62k
sR/bhyYxFPsjYcssTamaVTGR4ULBQYy4AK5bFzb1yL27Rfg0tFa4EM/BpiiybKHE
SO0kUmcBtnkq6IgSh2ZLwDK+auC7Jlwcw8Yw5EOHZM/DpxIcRfdeBDhwRoqQsh1y
J8YVyewBIc+Q5dDf64TsYVL+jmBauj49O6fmd/G5VFahYbSQE8dDDW2xlXk0gIwt
uRmSN8ASLhkxFM+S+RxWZZwsVIwkgUFE6Y1g3ih00IwAGW2aueHGNMGSdIm89mdy
zH1ygXbb+zpaLLQISF5DTgghRSuOFm3PWPTbtgSAZcDyvT6HyVhIU9FMMA+paBc0
Jh2cDGDJ8xaIZ+5feKCJIyh6soNhML48lLmD4ovDMgAAPz318DofVTTetA8VlLbQ
iLNgZGvdiobLQEzZQNE3b5FSi7dAdETHoyls8yg6OOQ+NfxWmdIcZ+VhvGGzqiLS
1vnBQ8sB7tcJzBCElWinyCMZlu+6kqXAoYVp85rvp/8ztZCQ9AeZzzdh4XQntW3Q
HXERCATNz/Eee43AHeG/Mu3Se45y/OtMEmmn/eK9+FwSVXaEewGytXbMQou8VO6j
BWw0XSxYIFnZbuWS7CDitt0w1JpccEctS1bpP/BDcLk1FL6+718sGszNE44Sdg0C
y4QpuQAs5bdRDgjeBkoruKXsbycgCIz6dFT5xeUaeHXouYckOp+B8NxTSwqwioS9
ZfO+QnURB2piyrvEQ00qM750MqkpoqRAlAj4RUxlnFB37tfen89GRDkkcfagcXat
ePdXDL5p7PFtzIPTU/wsZ+ZLopIIkXzjMqS2mn9UfmpAl5q5mH2HoYOghSRoF9dR
gAvZ5pvuo0wcMJVB17diBwCoW5TkIu2LVEgLfQ2Uzm0BYMdeNg2zNorlnZ0v5z35
Tenzb6weoM0+Zy4q6vHMgmM+WguBhPWBPSOraHtbWfsiMTRGj3ODOCrIO++09l70
gv1Us1ujv1E+RIBqzhMx/kwzBewlW4/Qyu7pEoo63Nthp68t14LZWEPYJi5q6WA2
uFL5tRtFFCiHI61xxQolpXJAeWWauIuYt42PhLr8vEB7idLN8/ZQUd5AaiZGszQj
/uQ/DCm0GCYD8WQW8KDaVop7zTjsPAlRu1/irxoK+W4x7XyFU5mZsWnXet66t70x
SJf2QK5DpcAvmy1hrEIaDeKGYgqyHrr095r8ieOAXHaWqkIgR3C4zg//jD7vlkTN
otTTuHzQbuyndxcMwYrIBaac7b8SkDn7leMbiT03WPwHBY14B0cY6UMJjXlu7X3F
yL8BYcEZNXw2z/K0g6k+b2RqwKDwVg6zn5MLFGOjIfXyp32mL7CWdFDqrYHZxLRf
1Xf4lm4Dk2T/7E7HpUlgRGlaVBm/jt+kqRUDRDT++sRF5WfuwM+ORwjPV9v8PdgI
TnepET1YPR08m9zrAQ0vtO02gMUA1FE/7r0FTZRmUNgQAyUMBV/RTi+hbHqNWqO7
BEKuqMPyu2H1lb1s7Ea1HYf9WqK/Q0bwkzCZKhflJ/UVyUFgVoOZKXsrrJdZ4i9Q
FhQQGDqFQE24pSPpRzCQt6dRxgcPfZ3QKvUEuorJMlnh98cXgSEov70v6WCL9GXy
qTb3j6t+51rSZqStaDGONMmQSx97FFdcc/xK4dOyFIA0Ast2wMAnmE/Y2CU3sS/h
1CrOWcWxtfvY+aZ+7Dlxk29VmkV/IOl4TZbV7SLrs6IwALGWREh2Op5SI/S9vvMe
JISVtKIvX1GgNV1YvlxLocGgxcjQECmYvTazM5izkt9jzwHPeJmI+tX6Yf2gLFEg
cXHszOXMpQ8FN/ytPBuA/58XMnEUKzKzH/85r6iwBvN6JwHeGa9i7fs5hkkV0s+/
RHWjEQ/OhuvgABImXM21yvCUhja9udXkEMEoT9LVwsv8b4zmmIri+HGMW3Iz9Jho
mzHk81Xw7oagyWnDgA28DlJ3ZCyLtREogwgji2OyeUojNqJFACtN4yE3mb/QtFZE
+rADWy/WwBELQP8iv8rf/pfS+PdrZ15AsmGCmIw+GwB0j1W5baXa6JRISnZGikLQ
dLt3+wBBQe7sONzWmfHm/kRKYPwLgdvbFLXRlcyzTMsRwWHbplYcgtTEkgkqHNLI
S78Z9b/u1E83BLbcc8EwEx1HR6Aisul/DRF5sj3uZBX6X8Y6mPloiZ/TtQqolRCk
jyg6L4+0qHCGVhpRs1OoKd+zIupB6QAdU+kqKa6TdQJyAEnDq8wr6lIFBIaU7NTA
akk3qhornv/6Nl1lCbbPD9/2i35bi+d772Fl7AL3tu3KGVwtSdGLUNPiRvxH3wMh
Y3k0S/+tdao4facRy+DYgRWpT4EXns4kcwPNsIk7vNVE/sT54KxQhbKmxzrK9o22
JfYZjAjHE9gpyW7fw3L177YF577+ajJ+sZytt+X1Qr7Hf65DfDZO4QRys8MwQ6MK
gXSaP5nOEhG4/wGUX2tM1kOfUw8BHaGfi1MHzRkohbSYzynvI3HBqqegRlVMylGh
b/0V9whGSGRqdeynyaWfYZMvmjCDTpQBJMpDZzHC+M8cp//PPqhSVmh1nWvUDROC
WUQgL4wKsgNQeY36kt81xp3a+7+cfq6N4aCZTw/KLNjVboHFxWjGJRJXP0+kn6/h
yva5UK54uoAPtV/kqfa8O8TH9zIv5+Rvm2ausyjAxmXmlsMrrHP+KO9VWCsynSWZ
383WFZxx5VMX4kqHOCkOQgRP3we67hMxUamPn5xqaXwAndJorLSVk6uDq2fjSWRU
JyOz7riubr7FEr0bOkL80SVsnsLup6x8XvLcUiJ8zPaTXDLDuEUcPIJIJas1P/Mr
0Lz7hMuR1UBvHi4GOEsUBaNhPEOUgeKnCe1I733NHmuUaxyIoGQxbQ717qcZfDzK
ISVqcaFyBbeIirNZNTVhW9U8GkBtMCQ5BnCaPAZoWhA3orLcDf1qXZViwznDqra1
3xS5Gd04wrVZpmrQDVY9tcu7SQH0+qGu/6a3DEe7v2eZEuX9Vz6+/qWamS6pwWFj
O2hZbnfC1wBP2woMVIRCxZF68N9PdnyYFro5aG/ImhooWGJ4eW18puf8w6u1pAjE
kdyNqWAO5rlsgCHqoECoHMYHZ5na3Uk1Wilk6Qd0164T2lv7ZQPBiwGyDkmXryCP
SQBbcI/sa83HiYR4amqFVaSqrD82rHTmzavNByNctKXXwacbgYtBdibkbtLvJs9M
sCst2y39zZItgXV/RPXMNHWa01Y01NeZMPVXtpwdnvYDAnfQt4vRex4m/hAo5ADy
uoYm7gEhvGVEN6fOn0gGHAulyBgDqxL/5/1qYJLNICrd4EKhTo/LeYaVMfHToKpO
9nQ2VM5QzfESHRmTs9ciYy2zZOYJNjKHsf541PscyorMrI6Z1eyXzInsWQsGqmlk
kaIT3mrRXDqMz4NngYu3i/BELALl/K4ZlgbkozCR/iODoZn+JW1ow7OXNcbWsbhO
zUMu3A/VLsEDvtEfMsUvCHBpiqRl4+6jfA+kBgzV11IOrP2/eHS2S5Z9Wdtwqlnh
GmofkrnA7q1YhFEJHhtnExXefDAus3r1HznuUXnZhL8UjnkwPi3+6UvuSGntR7Bm
BoKdxmcR8vOOkqanWzTz1u9rlW1D8ul7E9NLpkwPr4NtGN/EyzWWm7L28JMYOSH3
PDYOa+cmjtznHw1tZaZTTrFK5oBsLzyjjwhcSbysCQHEAoIR4LH1lJBqO53u2tYQ
4sE3jFP7uy24lwd+7NVf04bZJ5CQqbYappbe8SrHF50QoE8Y2MUoTAAZsT6tWgeW
QRnK04u1OxIgkQ4na7PCXL39d7GVSaLJkeSY5Cpv0Rdch8WgEpK2xrdQYJr7bE7Z
CrpHOt72xazu6IkXILxVrYq23j8YkqKFIXNIdIPF4daP2+Jll3GAgxILSbokHGde
PVQBlfUJCVx9Isgs+338juJDDnG77lr73Wy4rzywHoUH3am+A6JUshsnsuQvFtJy
tilPDnW6RXXdS3fJ+o5Q5rn+bKFgoFcrhss8ndNMvwNv3m+tWJa7CkNHTxDyqPRS
lvejIXtvoWfxi0uUaNzNe7yAZ9gKK0NkWEkRso7FiUe2BIl708i07n76Y/jdABkj
jadLhkqA822ON5FqHTmK2n7K9miBmviEZfXX6kDi3UpkMNQW1qbCDdlGwQWVrbYI
+vTPet6GOQneKJDsMXmYs6eg6D73n89cVmWA2uA5uiE+W+tTeYcLiOQsA3YvYzOr
tFZWwZv0FmLfQTdSYDeM3+0q16G9p0yGFSv2eHOQEJFpiNbG8opJTj58fZWxg6fl
3SL/sk0DIJllqISv5PqrHu+74h9GVdt2ONZg8L9g1tB9nChypdXYRRCxpIWlp3is
OcT6uzgw+XaJlOV5rBFXCHstZVpjRzhZMv3Toairx56feiBw1ojMOW94DVU1g7zd
dkw7yJm7ctQc5SZtI1aG+AJPnNq/E/kWvuEw5PA5i6N5a0h7+dXk80v73fGHxUgm
SHSLhGqlAKukyD9/UTT9+PqQDd3CDPwCVCV5sgUQfdLGQrS8hYfNZP7BCM6cazrl
iXWP8JfYe5k8F8yddEPhmyMRJzyKRLDScHKNS2lnsqNCLDDRG3zAyzrVRF7BSDPE
Dl7rxnJmFWxnCEU5Lbp8TjP+pKX/5PRYeJBFJ49UL1KKJnGITjROvNRMe7oZCAoa
0KzAkzloc2dm1Y5WcgynPOVpNdP69qbpga469vOUNJ5hkxhn3UfRv8bOnJxtZF+y
fp1ZBAcSXhSAt0uiC9MhDeirhRbTgVYdmKCIqivDC5aM/qGpAk2zbnQgMRETLJFE
dFVylwFbAPI+vC5u+2rK6D6A/hBHsZiJtgdmb4UxQW/DUcugCL8fk6/rYsMj6DXt
dUiDOKk/wU4WlitjMr8UKtCABuNUBPijsESKXu4NFPalyVYpIoUsK74Gza42fp4J
NDxnmu4qs79oTeSzyAkidVQwRr11zlp/m9XwNEbsCC4Lh0jCBC9ncgA86ITfPxoW
x/8UJIrWN5veuaFH8hMJKbVSKMBhh4SYo+H6ylCVwPFGCvfNlAVG6xHCw29pTlX5
tUQynStg0CG0gIKXSA9l6VJXD2u6i8XZVXAvAIQBnpWfKuAr269eAuFN75x0CUpB
a3+DJqnFQ6TVIDaB+K8BGmR3BCgjkwN2rq6srQHrK2qIWzjSUgiSC2z0UDjNMlbe
sQWZXw4hInlgcP+D7pY/BbzkFursAR5wi/OpSUmg3Tt6v2qpXvsVny7/ApG66uEz
1vVtLBQ6mOq/ncXUIxiC6mcTEJNxpDZuKVV2N397s110bZ5qSjRZSd28PJAz+2jm
PmGDdlkIdsaakPFSKo8tDOwOZmo/QQu26sylZZXb6C6YuCU5ShEXfF8VmAxL5Tp6
I+8pU6FypSxPaTAHVOONZkISx1PqbXUL7C3CnR/WwKJ8cvQOJy8UYAI3XlVLiUJd
51x/Az6jPFK30iG+EBY6SjDTMZPsMGfrvsI7uS08+d8jDUVKbMmWeP/uFxEV1r01
hcjyQaUSGLUHxdQyT65t9YXNaNCxK/stJzqvA1ERCeH/mnP5iD0ytggPh/FhleIC
kyhealQLh0HFKVa+tQh2Q3FY6VPOclHvJcNH4rGco/Dp5kBP5Do4sJ1u+LozUD0l
/YqqQ5Psu0PL0zRN1pDbUWV3NceVOohd+6r/LvcR2hs73deeCRt8Bxm40vMvU238
+i3e3DYy20Dv30jktfitJfff15Rc59EzuxT42mThRdqM89dbIx99MATVU5pjdKfR
SjxZtKXNmUxuiA0Kr/TK+xxGQ3O3s3MkQmmLDbEuFk4KYRswDhjvaHHgh3K8lVTJ
e2/V/RXM4062SSpvMkmpA0vhAGQ/v5WKlal5XNH5aUd+Qj3BZaMEdwIHWPOXqsDo
QUbjJ1ASlo9Yg3FJIs/3VZZMQzvY08+lXSJZ6DN98W1l4Knlm/2DwAzm+pmFPBdf
sbGG68RnVwg04jBLsiNWSmLJBnF/TUlkjs/35M8t5YbxTn8MRFTmxT4BIOHrZN8+
cvG8PldwvAjlulSW6548OQqW+RJknAmYqzZUGPSd55IBZ3+1+kUQkVxLiQFl9q/T
GOn+VYh2Sl4GI/OGqfUZTGQ39hOcT/NjQKQk7e8n9iLQAsO9rDw2mixzFU3SJTrX
3S66BJHZRMuYivq/DykIz6vSn6aErNG7yeTrh23BEZgdpbk/HBbpzdhnK/46dW+u
JlTbn2I0UtQPNiVUEc+Z/4nmS713GzBMGeWJt4K3t1O7emY2O2eqs6ztxMvRKg7r
7IysDJasT202VacirRRc80PoGLfdF+d4dZ1g71pYMINIMynvxRYoYiilwmZbHJkI
uOjzXKN/W1tk+Ip2sbaIyti8FcNjxfxjycTYAyTxT/XLjHSvyhgGFkI0LQTDnlTD
CUeacBmAi43wH9zqQSqmavFj0H+toCoyVb4qVvjCYiRAnJ4UK539nb/ZFkmjGO5n
mF2ZWs5IqPMitoXMmoDT6qV1f0mnPu2pLyUmRaiopR0kTyuiNrQqLjqOqUGyntxl
I73cOCcZ88tao5D3x8KMC3mAs1Tdnf98uJndpcenhTCQC+Zc8ehpmcH5c67e2gMv
miZ2Cn3neXFRpAJ+Q6VSRj9q97V9CIECxVvp0LgbZoyewD+iBIs3ejPhsXthUK7t
us+DBMVkfIQ4SGBso7VhoqGO2Kk1yXN84/N+5dU51oEwzXy+r6x653eGelmYUb6i
8pgd2+pO6qhG9IhUQrwMFoVU/AHjHJacLpTC+OGHlTo7iJr8VC6b5wW/yv+cVRjc
WQZsTb4+8HmxYazILbboc+98fI4SkReh5AbNzPC9bgwnb780MgQPdEXJl/qKWlLQ
+9aCdjroxyENgJpmhZdtIy75GNqEBpGWwoSifT23edHcHxrHGMbp8ff/ZNpnQ13E
p/PvogRZ8U2x7f5ynB96ZpzrBpYL7wWeRGQSDaRy5KZ+9t4T/ecI/TCTeFMTNxqD
jii9PGLTVd1X0OrXctbQ2oJV8ogJXbNrKK4vxzJLrJTgODxhqFRaVgZVwTneNMwX
UtyyrR9XiwhpDuxlbFozVOWblGkzcGtV9ZMUXi8zP2ifmjEUoZJFuHujhn5+5f1U
I2KP4BrDIKFlOjEJoEbWBHCfLCEerKRg1CmWc8Co/4iRkZoiSFu/qvyqgpDcMNJx
0byEhKfK3L32wgt1L4MOHNr1zkB4N4uhIMmDGMSpM1t583sS31SBP9cMjRqdGwQY
IXeGsY2RqD6U4JDirR13PrKoUea5AJAkgoflLDRveKZ0wirn68vUUPKZa3kw3xep
yTqmdE6+V53KwhF2vcq50GrUkLquxudP30kG4NHicBG/kIuGgpk9xtLqx29nyA/0
M8BcMwpMbGTFxopp7RUPzpUZTb0TPJEEqXUrhD/wwP6hq0toWK3CtE0L2BAF3cEu
RCpfLUHhXvyaLDQRA321Xb4QfyibrQtn3VPQoSzSwm6PRXspIuqskxfRPw1vQ13S
IZaXxFEdK1iwJ4D8vgScbgOkJ7gn5iUcBRrSQpIkVuaQbYnaRnpTs2KFmxEf7pUp
NKCwmb6g7w9Le1WFYByZXpnrB5Etk5fJWNvaiBQb8QpWgeo+piQO28W82nnSutCu
1bgkMlGnVlStnk88FUZYvOs0WbZOM3kIrTPBVasuXW36imt/1B0PySAPEZRIjTtv
Zsl2pte8mm7R9BG+DP+Hp7nMdKa1SGADTv9zh1rp1Zmqyz+B3DYo34BS3hGBoWev
Q80NFV2Lv6Tq7qA9VeVqVT/G2ybbT0t9oYTyUiumCI9wvZKkhNr5FMf4lsRp49QT
vDXH50/K2Wb8B19f2Z+E2YLTsyPlt+AUXGuTdvMm84wrtD0CUdjReRn1zSY/nqhv
vBFKSmVop4MCr4xxpufDul7+HdQUouSRNWn8qUu8fOQuzv3dn18fuwZzADpytvXh
yK7dqlRHX1Zl3GcETv9GcjE/Q4gHxNX0FQC8NLhCmnePZAh6wknvmul79tLyN+r6
TRcOqcpoEeWWej6SLE5mSzsZNA3GP6U26XZDc2A+LuUu8fbqDAJkkPKv3ZshYTkZ
yRmvQSgy1Vp4z1Giat/+StALiSnws+XvDp6k1UrH6ZEk8Hwt51RbP8cjFH5J5PXU
yLu9zLKu/9HTSZgQaDGC6c/gS3D1a1Bqf1XuB7EeiPzSsCJlcC7iRcAtb789DsMw
+ugRheOHGVvUjB6hElnSoAM6hfIensH9FSy8TjRmRUnGLfrQ/I2mpAultHtWmRb9
OTDwA7YuS14cnmAIIfFfH/Ogjx6q6CgqPqXCoYO39PCPqCH+G2bSOAaF7LdvlopR
k140YM3QgZl/GPmIrAMkErPqasfUjKfud6fMrCvnuWrL5ZN/a1c5tCpWlNOSmSbe
rayCs3uk/eh/mLIOtwKcd0xl5pvdaTJ1QibHL0bTNtwWaKgpJ6yovQeP5M6g6LrU
MA7iEhHoV7wyXcn3IJzU0y7QHMchAGgyTTQd+45d60lgEOO6JrWLvI/gU3Ab4aPe
u3SjMT1KnaIcv8cpCYQDPKGdphG6Y76XsE6ntgUHSHPUvvrkbVjgvaKlxP1bT8DB
XPx1Z7rbWRiU0HZeAaal1V1k6F6d+UyluLFs6fiB8h+W0YsC6hsERb2TXCAjtv8b
mXMUThlm4F3TXRZqn6j3fjFYVZbH/8jFetqWDga07vQP05O1Qp8I/Nfj30wg5KP+
CnRVBLZqe9VXGLt0/QZkHe5iWaJwg26XOfCLT7BEZKXVWmbxnBX97m6gBzW1qvEt
CIpyZ7A5diR6Pvy6UQQXhlsKYLNnAYxEBdnFiu6YK5v3Kl/WxdXbBwxf1vPjMT0+
SJErl/doEKxkvvY2yi2GiNUjEX3sniOXEewb2VKVjXgCcFxbPpJvnhmFnjgn7ffB
ovRmBX8NbvNMFt+w6LSyS9WZx8molqKKNa5csxyk5HxITDZWWL9HmU4kVUr3kD/M
yj0WoYojNw8Ao8XpCUzHn/SOfz+ocaW42y7Uq0N/M7NXgyjyeVfqYcaD7nmkpVsn
FARqZhtUnP3DAFP+Q+b4fmiX9XUK0rfDtve+Yq1Dl6zqE9hv1DrUo2hC1rgkQb8g
09QCRNRen/7KKHfAU3dadueDyaCzYkUqYer59j2smpPJ0bqMxfJRLkK5mB7XixBN
eDO5VqRtrFKdk363qRFLyO1W1Qw0LHB/1+yLCxOANxq7KbsdLBT554Kn08ZkzRZ+
of2+ZGy+kHuAznR/ZHVfXV4Sb7eawxELnogp/mcYAS1+E2NqKcMOkmQbvZgE7V0k
x60ef/UMJwRNe6B4eJcmBa/IHx+LOfQ7dVJGIxdow2B4Z+P/5BKjRrqNtdi1rCzQ
ex57/mZVxaIw07DOfk//vYmr10UFrEKzPIc905khwN2m/CGJuNgVKU56bMIvzpcp
fdkqcaYUb8dyhvaEy4bQSqSmFEX8ABZvYT+enEaGzM7eQFz6xuugDz5IiTKUAIs0
g4yOs76Z17liD/M9RnuMHz6/AyONdsNwu2ZwtFMh2p+ivtyV0naakQaGK0K1oOfy
LDbkM01VZA36INodyjGkBCS5fTAxBneB8NWFegwYtqm+gy1PQcBhOj7DzDghFzhN
Sr/f0MHKp8G3nLWUfDOn3CfPIMb5rPZ8cS+R8U6okAGlNyh2+uwTliyKmJGQOCGc
MA8eein+d1nmrZfm2r9tgpMqjMdPJ60YJEzXwqZKo5ffinOEknhWZSin2OBG31x1
73zydGgj4a3NQpMPt3CAzWleyBMm38ZTiSNgAX1OLaxU18/CaY4aKWfoB77KET/t
VjWgf10PJ/L0A198dLOfiotCrT3IySkXIoUzI+uf94yDFenZoTPSszPBzJKSPfAE
SaAQX0KWm1bZZzp562UDeKP0Cd2/4VNIRkHTiYnyxEWynFSdgeu7ICuWRYJMUrkt
lWv6BEvnr6zpW4WLO2GdEnMHnJfbKbaRdF1Nhgocz8QT+7rAGFuz9X/lgfBpS93u
y36FrDddTRRPjkZqI9MPW4Z5g9IkXQRPR0sog7k63rRo7BZv4xmvaJCdNxcwicvV
c3mgbSKLmuvMq3NpSLJkGXt/RUz2s+wnG4kdv9vThkLa82mWa5L1IcbVnspXpm8r
6mzZtEExj5DWs83pMPb01N5PkaHLTEmvBwbH+cblC/U+WoTuAo+W9yfiISN3xipm
/3i4o7uuuEB40sn9ZjKi52A25T2I+1/7xfJzujl9aD1QXsl3FQ2WRiEz4RtnhSpI
TLzfoAoh/BODhvKehZxMuXYDSKX2ewaJcjUAqyPuFJL+ownhVRbbvbbWIVa/OZdh
tltNS0YOw9RpyiayYhj8sxlzMPk/aJ9MFWGt/axtJqSE9/UYtm0lU8ZIkm4IHXpQ
mZURc4+AyRU2fB4O3l74BP7rJ4DyNm+Yo4Ej6oHEFkiQqaTzEPQXIeyT73WkkM53
dibps394EvDIap4ELxtIFdSiQsjDYI+hQdYSBbAW9r9aJI5k2q9cGaZ1sl7SnZpF
P4opRLYoGPg8aLpIVaCpN97l4EouSSgGmm2HTmAfdZSvd7hQ7lMn//qrH+MA8KOc
uPysdHCzBYPP/YfsaCCC9yk6SV9Lt0yLg4Tl2AELGpoxj7dV7+3HoO7IsCXbbUfd
c0n8h0WvQERXRByJj9p0ziLurBRMu28vGjJYyCo2JXWF/AsM0ew/O5W7y4FYTLkb
gDsPEoWpGIuXVvBIe8Z+VmwPZCHaZ2ZKK/NNTDuzA3rGv2RFOKXwNDp314knWEge
AtlnSdm/jn3iwRJss3XCU1FpjVKKz7QFACFOlk0PjJ2RYApuyRv5TjiYnc6kDmvY
Ckk0qjj2u1DCN0wkce+R8GWZTDFyRJcU/3H0PiqsmMEjLppbaIL/YmTB/oQoUo8d
4yVdDPr1JWYF5O5zDDhLqUAqllEJRVPs2xT2mS6pbYpnSHk4Aw6Ve/hwPLFTf9EO
gYznrS8R1wxvVQz8Kzt8PPO4LQjof/w/lEh3srGM4a5YtwT7dNgGtfRtv9j97aJl
t/YWa45TuPbNqgkoo8TA3Mj9r8Uc0V99HMuAJxZyxJ1LsrAbmdL21iMp4m1M4jpd
EpR/qQtEpIpZVSEgPjnEX146OVoNZRI1MSC35xwzDoc2OX1VcLe0QdaLNQ9WydvQ
DAXHXaMnQLhExVAjPR/CZCnE5/eywm0XyljF1PplQmQ1P2/uJQ4r1hUyxfwPZPnb
sFJSMtbiEf/FAtnzr3yYLzEZkKgGAHTmWvVqyXzHEHQoQG2N9PXl80t2aOfqffAB
aKovOzah8H90CAhzTXZIiVcDAqBxdR3+Ds+t9KPmf4+qOiDi5Ca/NJLQEabOn6ik
IqeLpNTdI6GfdF4vjZvTzHV0NXns6IoKFINXcf53788H+y1pAN1glSxN1/WYQYLV
dD6PVe9UFx2K86GzrEe1VjUckbf0fAho5NbRWiES+gotK9Xn8TSzYFSb3HuZ5N/N
5fNq0GdNZou2vv04QE9L6HGPrTYzZAAY2BhWhB5oKAYsuwtZv2VJX3bgj6U3mJrb
lE42V4Cp2/cUs80rum7e95SmUAPXy9qyqsqAf16v10DfElUK+2cCqfdkpXR0MJAx
SD3D09xh7qy5NxJZwLpm5Eb1eQ+gqAxAPvIrvYKtGKhHMpDFGiwxA/GfUVre98gx
eTtmjOagWQSQ+B9R6gWPsmUtKvorc3LtVvzfaIKcuPOKeGYWL95XOPWn9yiPiDMb
IYsuR9+2wZ+SHOBvMjpNTKkTWnkCRMcp/Yr6VNO1lnhC7szOHMOIRHS6fP+4uV8S
p9OrQuW+qSqMe+fVIsVwRCSSrMdEKgkhqQDY7bFAdlBKU39JGDod1wg63XKtjd1x
2XL9P1q3Y1Lix+68UlylUqGQ4ZmizOD3MYRIzBipg/jjYPIbYQeFWGl0vvb2FOqA
u0zM7RfBla8rDu+XM6Aq2F/vaibFAO8GvsIjQf9UjXK/WPtxeeKvbtVz7e6zKc7h
3f+XJoMYoiS9042unGs41L3ZHRgX76/88CX7CtLkUA2Cy8xGBrBR83tcZWN5OXh0
cezuzvqCPruSJ66SP4SP7Wf2IYSAYzAhExnU5ddBpEeROM+VWI94ZwtYytQ6AsbK
sON9w7bL5emGfJX/36M+C63nN+qV6LNo3tWSAQDfc64jrpAZ/AiqBgzad30DtKwQ
NoF6+F71jDH6frkRbhZvWDR4O+IyZijkTRmtgfOnkS8Ouoo7jPOdFR80GynjkMFW
AD/8Ne1bO78jSes9TrEavlszBgKLLKV0PCeYQMJgMcmggKfTXMBru3HdS9zMa07K
8bASdTXUBDFZGDq4mT34PnBtWbXPWkIeaqZR3Ro7z+bBG9Nzq7WCQxB3WV0AevXF
PGmEOimWvWBHem6aF8VDR3tv3PiIdeUl+Aohy1eLzNFrEKMhGtCZthgClWINQ/5s
PNmjz6UwNCFivfr+gsQC4HgQq0rIGXv0S74rls2XQ/VQYWGMGlQOFHzt1GQX6xrN
7PA8+0mlGTwP+D+Yvf8jSYNF/FIBPoYpIfi6VWpusQwd4F0sFhmXIqtp7TTmiy/u
obf0LKdq0M/lfxJo2YRY4ENMyAFcLdIdpbQnHayrVaNHvXWZLzGRvmseJVhHh9Eo
LRWSB9/6VYJ2vOJ3qgr6ZElc0ob9DRtInUyewUPHGCcTsAkV1QE9vsUWY/ERO48D
hu39IP3n2UuV+HFP4s1MGuzNZB0Uq1bb8YfHGGfl9wfXN08S0X0XBJAYUyIxxSU9
wybSI/QmOjdCvwJNWMcp8aAxOxMOskKqhlq7EB/X0+xZOOCt7yKjkyT8TiPoyYAZ
E5/alBtr57ryUwoMc2/w2qGEm7c/qp/iBANcHwsYibR+PDOW09och2fiAt859a7z
ZvSUe5/aWCPXgK9J5RJv7w4DRklVOoHModlf6Zd077zZPnlI8p8XxXDu1FLNFIGq
pDpyN4Wm/JFcP/AffnD+G1MVjOruXNigLO2s12qGoVaPqK4bQF7tOTi3mpLo0D7m
8/MBKYpw4sApcGFf6FEe/7GiLcgQkrPPXpPNeNgP2BrWzzHxCD1e7xVsOv092Skm
tnT6cd0WsXH0MWClfODgNy2t2Rn3KGsA9BfkfVC1GPUuZQqgHecksICSK+bXxgPG
JQAiYWGdYuGoa/Wx9bdJ+5IF2PZo0sci1UZWZl+Us/E/EfjYhf1v80dJR+KzsD2U
qP9lLAuvv9bRaTXnWixzGxri81UJt0x4Nfclre6T7uOwPHqrlMVbGat+sY0kVLeZ
P0np84WjxaBCR3KphRmBnxMPdzCeqfyVAGSCwN+OadqeSZD7oQBNJI86T79iikYM
ycn/qk3WXcRnNwN7zqX6Rex8TJG9UGG3JBvWC4UEThag3tk0t6io8lvSoiE8hwgo
8E9VwdPVGrrCIuMnnTJ/1M2iol8z+/M9BW0LcAMZ8FD91t5UaZzx0HUV9tVzNPA9
J6qrvv6lkOVEn5zS/ZmC2Wt3VpcCj7L1fGmTYyCUn7nMoadAuSnsKh9SxuIGciO2
CEWh+oSS5dvFOx1ozGtHVy49uQcoJfDRygN5Z/G1u5a/KdLozksOIj7It/0UmvxU
Hz7vLLj/OWLM9n8cSqvx0Aq3d+qoUtfCC5sNPcP1aXwMC1sDNsFNbGlXMsGsm1J/
6IAu/kCCBCuRkIL096W+GcRm6LsH56Aqb09HN7QD6KhSZa21n5oBAmQJ5KteDkPf
6bmS1IVoVIN8cZYlmyvySrCcH7aQKpeTrVjRXaqnXiosIQe6m2CPZLK+nl9LSb3Z
KDauoARVE5f5lrWjgyjegEjqqF1QCjnGgVg8NsZYEhrHRtDYxylG9DCK9/3QGiiw
FZHvNy+50F4odZ2isa9DA7FDF5SHMrZITN+9vsYBqCx/XoyHEwOqjbvdzW0o8/nX
nnlgRobOVOQLG2h2h30fG3YqPM42s9vPDioOk6drv2QiYqaKkgLLl9B3v7U3B0R5
3iVZqM9epWJUb5v/mf+TkmHcnHqdJ1BxZ0uqmql0C+ySRDx/88ebtkRLdgvQ9+ia
mqOOKAcWRPBzWehkz7toZd/2F1Q0zLJAikA9x3fkNodiDwUM7KBuFb96Tn4FxMBv
XxzwnMqU0sjw7a+4fPk4qKVjoGyXVpkwtMAxftbtfQGmNLtZS7iQFXraanHQD1qs
ifizkoisRJo7zggMQop/0W2eO/cF7kkHamAtndqFdIC8Y0+tJBD5timGgJHx1qNl
WdBbNVllx2TRrQNjwn6fnhhyCdir+4O06fz24YVddTAS5BZ/wNGSazQJKGCy0I20
EKcy5pTW831Uyb+ti9EoLW3Z4MUVNG0LCoaaIdNC6ycNO4Zoi35hzSmuK7gKiYrT
wmE3kXt5XLEod5hTeNVHNPGdXDJCW9m70u8QmiORr74VNssfg541kRVUhthYd87x
jmaNYISta1pl03OVkVkkAxOqEveeQAZE4biOJoG9hwBLH5GuzOz5YPKJnefsVwya
2YjL+MiNZz+bY4GWJvY9EWv82f6X3Pe/077IPTdT8240YGpJk19j9diw3ZLgraH1
SeH2HujA0LedrW+ZXQdAKdYYA0tKZ7ZSlb0pSgpDIknd7wVyJPxp4QsX6KX7+bpV
3AX0FV50D8VqNxtjZH4eaw+J6+uZ2GvA44ERTbxDuup4FtAhM0q/2I4MmjxDWLyU
cvGCo12MSj6VB62GzxJ0EvhsfnI77nAS6VmSwFQ2Jp/veEBGiYwkmbmj5p35+TpN
OGLAsWz+G3zegEEMlnA/aslORN5eNTYqfrITM2D9dJD37FohpyUxh+/qWz/+JF0j
YVGfUaQKK1b+nA/Sq3X+7Ci7/tZqLRhcnBZNW8eCJiF0MgW6lkwKTFLSD2MMWrXS
rv2fEdo63P4rL66XEBmEG4nevqRS9vGaMrlPOKLFQpThcvpGjl1mhbzjTO6Lbs8l
O5aHKmlmtYX3HvUo2zyEWrtoLeCTRE9vv3D5S9CIPgbl0hzSH4Ywr4G0IGDdGgnK
2oAyrYy50+ST3dhCjU0dVHRK044318Trddg3FOlXJ4kBZh6zImSDbhL2aKkGWxLV
MlrtQUIT7KK/HzbZ2AbQB1/CsKOVYOGOVxaBZWIccKiIhZH1euIqipgrxxIeP0aY
EGzC6AZALtqLnhuc6yWIy486QueFLQwAnXZ+3jEMQP80cliec/mZhSdWlQsmhEDR
yjCFTL8WcyOtHfwEVxT7TwgTP84kr/cErFJKGZUPR64GsHCNiSRPtcXbDN6dG5pt
JBOWB1ReB+HV4DLeV+mYCahqWUOxZNv8BWg/VRmFkdHisy02ZnC7+tUYTfhgjfdc
PlyfKZUK2jspaHPOlOUwwm8XIFViVlKYueEokGrjNyE6KqBDJJzLgfzQMyouCBTp
HnjE6G5MwJCRSixtYvkn2k828Pk0rLpNotv7s/hJMio6NfrNvbwcQcds9rFTDNg1
S6yWmNL2NpOScgsaiYtLzGPQN4TOu9CSXvkaatWYK2ULBdIJP8GnoC6F+Fcmhx7x
qG3R69NL5pvz+970l77znM/ZnbY+MzPYDAaaRW1exLvLRF5+zdBv9bsYrQqQOItE
GkmpSHm15jvIIghajNSzywXARZWpMxx0vTA44ISfsCL53iU7UwbD4PxuH9iS28ai
AYnEU/5ToUiB7bGOU+FhI6jM9GuhqEJ5JAL+AfFp1YokpiBhoFW+Ko/dUQQg/NY1
qmasTL9sz49BA9ZmGbHJoES2RSMtCBdZtklqbokUrWOnErRZZAPNAkmLURtRC+g2
x01MvgQRycbiKy8GuSJy9+EKe4jS98dxtNwL/BM0TuhMNBnR2Y/uN0AEPMAvHHX4
v3XKrlZtGjr2dXvfTdKWeElyOPXBkKm88Dh5AHEwgvajsjwT1Hj/2n7Pp/jx8ZmO
Atyw2OreX1hWzEqn4d7kwBGOnPpBmPw9/D7Pg9JX1FbEClsPdQkc7xVcRcx3ncbr
6jdnw4Z6DGRc2AN074+jWdepWQkni9/i9W2zXpBULFbvKGCqDHGy8tILXXbgVnIr
7rmh03ymtHWNfCRh8Z5mB1Uj+PhGr7oyYgtQu6IZuzmLQBib5z1xOlXiCsm7pCvz
Vgvbhh9TMY01cE94m9HowKLqeibHxPcs73QefD/jImQ0GBzxjX+0cKmhANO7kx1f
juLMKBGqaz1Gf4aCXzMXXQyjLQBzimHFw5tot0phFPy5opF1iri4ay7ZG4sl/tTT
MDwp5dld5/+porYrURvVsJQhd7sH/kC0zuT8EOmIKRi8gVwesXI+49jwU5diKVXE
ZQFGSvXKdzjsJrA9HEBdLstq6x/CvvAEgZz26EnWDoNgXK+29aHhXztH7sWhYDPE
/XeJvl/GtrlA/MvvXdCkLMA2i5oiC6NBEFjskREpUUFjP10cTkX730Bz9f0o/Ssh
ocHo6w9+12iLbMk66Ej4iEVqopU35Ha3xUbvk4U5WGNAlrerf3eL5gI1iglXBcWK
b+fOHoa7RtOfrELkkGEv7X4l/pqKalcSf3KdkR0IUeT7D83RU9POZZSubMWBFUvp
Fx8Qz2EmxBlPMJcyZ2jnhgkvx4vpvLhufnVnlUVtDNXjzPmYOQ72pR3n0s7sl+Ba
PUWuA5VYBrotFQs/dzBEFjbWqRMQseHQVfjQxKfLZpHS+2+/9xI6RLj1svNA8wGn
EdFx51r7glX9A1Zc1fH5b76Bq7CQHl5JlzedTFu6aRNWtisWBYsgu5GhCg3wf1KR
s8RaPOH19DER3qVaU44T4GuKFsBLLL0fx5h2VGbGQtXuKChwmc8y6UgIxd65vn9r
tnu/rkUqItu6p/Cfb1n8e4kFaDFh0xU9bWNOeEV/s2mtAGQ9rGTwO4bpwDWh7VDE
6RrtVTRiRm3okfk7eDcMgzlcABrZ8kD+Slr8+QvJ1zg4AXXeERARWREL+g4V22Pl
15XSktiOPGLpYTqbNU3y5oyo9UlZbqTqDq8DQxhbTcCzGCyKlNfiFRw9HMiTdETK
NLy7vyzLBy2M7YdKYTd2rwn/RcGIlM9RH443Fyop9lM0vHoQSG7Bs2Vl3jhQViXd
zar441u/rSAzIkaT/JfrZg8eOIXOEN4fl5lT53yNnxxla9+zDIaYDbHc64aUl1qq
QyYR7yZr1aKIP+0qcrEjU9mpT8yWjKWm+oxfVPtEwrx34kMG+MYL0Uf+ow5t40wP
xeO20r9oUSAm5Lp6QfAkGYHlkpDiNmVd3LdPeFthJ4M5otO7UOjLwa4h7Na98jno
/BH4qBUhlDY1Wcf74Y0YqULSTWegNuEcANVRViMkUbP0R/GSXXNKDCyr++FMpP0S
qUMLApBnr4dA0PyE2/AGt6dLbKBTzPC9HXk2GC+6MY4vWZeFWrDa/3ivpT0PHLi7
fID9xH9N2cOtmqfmJ6GXa/MYs3uUdIRTJNntSEMlc3NSGql2A6qV/lbKSx2+H1wu
0GrUcOeQ9GVniIcVR6fOkjHfSycdt2Ays1rjUw+n68bOLUjk3u7080wHATam+McC
xgr39269qzP7fmPbyIrIC/WhxbPkX564g0p+4cP02VVwyQ0tcoOs4AMBz8ybKD+k
MGhu2HLaU7DNMuAUNrbGkTNQ4YDKeurGY+wud1rDyiarPe44ySl/AruBAssgSgYL
XvJjizFdOyj8Y1jigW7/IRvOYocGBeYonYEegEG0iUljFX1f1oh+F95f2t+5Avdv
h2Efp711sknt8GFDZQ5p/FWC+W8VpCjIC3L5WavIpQWjCDWGIC19WhxHC5T9NxHz
fSq6kDSsMT7EWgs8Ee11Afe1DP4CBfIvyEWUYK9CQs1fj6f+pZbs8J84Hz2X7Oa6
Fgnn8cY//5JyKtnR6sst6vD50wGwhoqB4Jll/VCer6D2OlVubNjEerPrR9O0wb5I
PXkdcjPHpniv1GRgJBfFJv2+3u/XWzV5QOJxhcrN7h1H+9YbVbRxFG7XF8+VOuOE
rCRwtU9VBXxy8PojBkz2Ad4gVufQ+Imz7nPxkrdamiu+YfHdeMT6/8ISs6ln3hTZ
t5S2LtmWyCNhiMwT5VHPMdi6mIZuO9+5OS2e5yknOAZ3jcsKKI7Z7cMXyRIsTqs8
I6Adwz+WwgQYmapxmyPTVfHXEZguSPLf9Xxoio8UXbDtaIR62cXfKOimsfyeqEUf
rJ1O70zHVSEOOlsVxzfe+xJhKlzowN8a0KIESWKhCFuYQcz1f9sEJVupxJ8ySbmM
s7xOwfjMZquDXO9/E3w3/AAfc1Za5O/PsD/n3I7vB5xHKGPE5VGj+oa+tne0Rnc/
no+dwDYrTe4776aBasuzooELrWgwmqdnS0S22wQzChOZRuKPnSzyH1Ayluob5mpV
qt/fTI7TOirsS9NwFMu0dRyTmfXGwEoRyB6kQq93649GglAEOxCl/Nnulix6zo3i
z6A0O3CFUWu/iOWnYrvhJ8BgTF2rEEhuVw6a0DwGCs1G+Qy0E6ZBB+5pUhY+BpQs
LJT1gdXSblEbHHDnNG8Hzu/uYMdnjwxBsdxb9HXaxScjvGVwA4AEH4V99M9E6Jo0
qvCyXPDIuN+RzVg5Qj62fWyU1LKYlNal0AaOef+hczegiiqsv8lQpHElTghKo1Hg
Po0W7yePlGk+QkV/ugDb3PQEjEEC9ASd6yxajNzSQT+lEJ1HrDbIZov8ZS6MabA3
6iUUMUFlndKUT442g5c5S2Mm/oq/ouWMygXKY9Mj6jLEg2w34AM0E3j0OecQ+Rgo
sx7ll7yR0lEH+7PCbcNnIZRO6tPUXSs9nH88pgRHB63UXEjTaAPKG9y7gw5O+tUU
g5n+TEXBUJbYzACONBfEZFvAnkkFojp+MKcY/QLkBCxZL/8q653kpw4mzF7vd6sD
5iXHoEgccpKTsuVuMT66Y5hY+XrsJ9gpVtiC/2DZFpUNoJEB61Fx2t2fVHZle1QR
Kurg/c456HFstFM7bVStnMmR29Y3RpbeVDSuaZwIKIIT9wZwi3hyWjbRqmx+Q/2R
uGCHl1PiPmefH1yPKkH/xg/c44jX3NhanJ64+HquKcykAuIaJQkh48XrDBjsgnUF
PHGqq5B86z3YW5ia9/imRR8NiR/o3JBW74s+zl5sITqz5+WEO3lQTyi/iWDA/gdb
L8lMcMth1QWShI6I6bQEMVRkg/IJWUUpR7ANrdRxcZc43MCqPv00dPChlkwframA
GpJ5IEepnOsoTJuI21aAerErhHUokSD2rH78BE0elNJTfowIbPAxo3vjbbyp1KP9
MpQzDa+JHswPooroDFw5vBJUv09MwusJgYOjaWwBf2TkhsnbQeGOk2zJXYt/NtXI
jZ35gVuXqCXUE7mvEStwU0IGQu8xPP6hAqYZDUN3LdqrRjWKD6fjsE9z+77+ntau
X+cucfAOeteHhWA7bI4lKWoxhE1OHa9BnwXOXmRLhJ+6/4K8gugHOdss0jX8P8xC
2B5mRsnns8yevLPKmF6pmVxCJRC/gPeZmJhtt28xQVZOzdXU/hYHlExuBsP7ONgY
dlL+iF6fw+IjGJuqyorW52FGQNp0wAaHUdNluIhwUwaPNLvTMECe9neWKj/CMqqz
BpzpnB0gFpz5H/s2Z9dmD1jlFNIubiwnlMV4cGzYmJ5kM8AoPYnJg17083w1eYlh
URmSI0x5SpB20Z9VHH2JEctZym0qEzhq44Zsps3G/WDX2flb55rQYeXZIjtIu9SE
8FslhMe9143EGNXYLmj7OzymHI/n1K7CMZ0ZAo1ocX8afrkE2pTueITopSndqf+U
uLDLtLgp4hcnScxVQVvigJqroSkZ1jwOwbn3/zrqydMWBDOm0EGDmlM7FjLVTHjl
24JY/ixNbjcU6BRlIWWbHbd/o+cjAtvD2dsjS1BtI+ietPD8M48TORFjxtI8eXqq
jT9jnHvgt3EjZUVMyLsqdi7Y3V65D2e3xB0KCgXbmVqm54V44a845odzG4XNAco7
cF7H2MXUvMSSjjUx21Erk6pSc1d4l5VcuKaeLfTCXU0QM9/5KR3TQhetS1u7rnJB
b44rUuAfxScFZuMoY5yASrhNJ4MH6C8bhhv5I0XDsxf0UcPblN4VyyJAXYSx1BG9
kC24LgFZEXP55skM0XmIAmz6n+S8tcxWznA7JRtYI1PThXC+LNDbBA8kHpyhmt1J
JwmxBs0NIn9/yWYJHUiyDK19StKM08EdFf4HtqaefYgQvecJVpVR+qPARhTk3kGB
Jbfh7KfPZf0k+QX2LnVzb4nIKQe0grtcThEsiWIBxYQxmif0OVY+Lx731Z0vrL22
N8Vxhsjl1yuO7RdexjD7jdkviHbVaXaf1ZFFLM8ck33q/HeNOY+UBvGc7zlQOu9k
BQ1RgsRXExWx6cunFpdhsNjaxZfUr2KaXK6lF/9acebE8r14YFDRWD0JUcV1Bs9l
gsML8FoZ4iwKn5lA2EsfVj7nN7ILa5ZpmF42wW2fKNwb66jRlDT+R4rrW5Ma2Fil
/hu30PgxGbUci+X20TPJey3CQ4SfqPKUUxe2G0gwww6lKAj5DkHQL/0d4Ya8IX6+
Rfn9USxUAsIJpV8puJeJD60ip001rrSHZSUScxkCnjSu3LQ/UhjcQb2RUHosBPNu
suhJuwa6nXPhJXJRKS2LyT87jaiLmW6lmYvdfezXhX4INNAF1I8WZ1boI3qWvFxF
Y9F+1KyUhjpsmJ2uChqRKOH2U44GKWhQbrFtWNVgaymhjW9eoDCJsW9B++589elV
9q3PDFnPTP+79ng4BMFx3WefdmaxnPYZBLqVoTWi/VixA/+5tMhFW0khBeQ6e3w9
noPkPSItFZBm89AuT6w3/UMS0Tbp716F7aTb4Ft73T85bqWsDaVQsm2JTDWMopK/
nU+t1pm8xBQUtBzDxMtvCukFy3QLVv0EayxcbmaEqLB8IYToc7rGLqpljLSfq8UH
lBNd4F2VHYGZ/5yBBc6d2wqyrODNp7rUmenQfWRszRcxxp1St+igXGa89iQDvRat
A+yOTp3OOsuolvucjKHcebeSvcpMlinzNc8shSXrGtDD/iyV7B+1+doPjjfJyRWK
rRcShbaiUwzy8vuBMN9os9qo+RqdhAu0od9UPVrejz/c36Yid0pB45ZCr/caRsew
9tkTrKHyloZvoJBKnFjxTZ5nWprfzcU6bqeneyJJg3kg2Wc6+jbfHCk4DD6u3Q6t
2FRpjZGdmxSsWYg8uP/GzTgdjuIx9hD+r1ERHMdcpIPd3kceR8YB+eNqm/Tkslv5
BB+Q1rtZOO3QtD4U2kZOEoiyG6c4lvQfH02Vli3GbRnoGHXzNhLqwVt5BV0ZIOY7
XmD4w3c3/36PTBGIWKLNq91vEh+OjhcN/Nx+CXsvJFqkBzUC1XgZ9a9ag96hLhWq
DHieTiSFP/KiGvyCOSgITuphDc8isCojnYb0PrvdN4Fnbbysn+74/CrBKCcgZPlt
7Zay57s4/zMAQlObCRE3Bp66ng1yW8KaRvlzqVasfsGlAMjKQdZzJ7Li3iObGmBV
DOJE42yhC215Pba8w8/7bOMESSVwHqiRGfVcWhNXPMb3mM1bMtSaVgUBQu2REOre
g2BQErZpxUi2CNIf0jz8x8rDX5D14MwqU+Y00HRoIuQrcvkc+PxIEzJUuUByUwoS
l5cT/UcXZhNDzqjXVCf4bqCCKxNGoQh0IRiIZiVBh9KFj/t80pv9ZIFrokVQo3d0
GDyuHHMfDIPXC/fMFIZPJJ70TG0g1byvzDCXqxmdUfyg1BuaCadmZY46SGTyjVL/
S36+R1fUjmoGSWEsrc8IT5x5hMB2eh7qf3ePbQlFboyt9oqO2EwnSAAXxYYKolKB
0aZKRztIxKi5e0O//KzW4q8/qNWjub99bYr+S5d2ZVs3fQQDii5n0TSbG0OLozd2
FDEzOah3prETBB6O/X/PehAa+kaNKIyDCRrD/3UfNnU8jwQin4qSBHJcbrDuUjwj
LrP/dBjH9vfH+PW8T+BhBr6eA+AeWT3XJPYZ2ZN7K/KiGWfPgfgGeY/12Pxx9mC1
69oDTUuEXiL/kImXUFw7FqdTIWaENCmXG0VrQSv+n8ciYcxC3vBZOeYqiIGekxo8
aAOkbazb2GxqV4BtVL7ro9QWucl8WUxwRXX5O1Y0dZAohCKmXPklmMG3dWbNyfNo
tS8lsBJb0a+u8VxCTVyOpnVp+98wu5oi3WZb7UsbxGYbV/rC5MIdwEgPajIhRNL+
z4fFMUZ6jbVXd/XyO4lyiSK/ltijuETDsJbDPa5O6lWUkt3RoBc5s1lg/w+8g0hj
JGIXljtUSRdp4xJI8m0O/ui1fW8jPH82bnih6IOGZGno8QBwSpFSr8bK91hxF7xF
w+P/aqtBzshmF6SEMKUXfQ4RGrdzd6uSElz0ZofEvNoyKL7iO+vFNfe/DQrEr6A8
nYoZTdL3Ghxrc1A1bO3R/CYA/jmtKQdwaYvSXyyYLHuThH1Lw0rypFkr7LTkIDpk
uPxGFTTNPPWUYbi0mmswvZAbEyQotlw2nGfib9kDO+L535GAB6rUKanD/O58XLNc
l4eINg8/6OVjloynto7BUhqHmMQBPA8BlqUSnZ5aZVyyZgcmb8N1rPWAqP0xhepq
WNompr4oDC+5h3e62LPh4QP6m4aCyVQES0Dzx5zsrXyhLOtqJQ0rrI9ekidVhPEH
1d3X5hV3A6jmL9nno4TN9d64gcI/SinGdR/wr8kv5D6QW42DgOjNsALleMHTs8ZH
1EFl7gYfKu/2YVm1vlKAjx/Arr3rg3dE5FhZtzxkZ+0UhjAdyD7bIJe6d1Fu9IZH
VYO+i4qpReXyE/u75nmXvhrnmDA3rI5N0HCJCzEa2ujYE4VYxRQGHibEC5n5GZBi
rsKS6SsGrtXMjg62gpuE4OwK796yLToS1mjKwpYFgnqE17gseYUAKH5Bp+I7V0m+
cI7puwUSuY3g78GdRbCeLz1bznlyRQ/HC7TCTVof2eCZ4qT0yFQ+1JYaRHZB69RO
pXl4kBYX2SBkMFFjcC5PH5nQdmCh8Y3nlwhZ3dDOhVWBo4la1vOJSAjtsFFvlfC5
0uyXQEhtT1ynYlUYd3/iqCO4xiL4AKsI7JEXHyq62tCoYj+qOzkll6BBlZBZdJTg
spLREvYu4KuyywjtvmrdZUmKu7Q8P/KLNQdz9wxLMeqkMkGHW+4M2bqYgsiP8JkJ
KtGGScWwHmc+co3JLCsXLGpD5LGVdooPjxvNsZCbV3CdFkZ5wuxUVXSdZ2roy4Mj
A/+PVkrDwa4/+biXqJOhKuB2E+pvbIWC1VKfU0pYXreWj1WAlE+o+uR3fM32KBJM
k3IRZZqfw0m+qx7I/q7X3jyqJJQqVDWwtEjuxk9isN5eC6Iz+jZJQKfoDiaJUM/H
leO4Pot0ruCcPKQVBgfMVo/BS1+WdEeQRyYSanzXvNmCxDRpU5RKubFnmj5QOmJ3
gXCqswCD2b/f9IHatiYVgSBlL2ClbTaKHVtdaBxWou76YE3Mz5cif5mXAUyY1IUx
z+GqmyQkG/iWjHbZrCkltF4czhEhd6cruyU00NE/27Fkpc34HgnLgECEDZdatXXp
K1UuaTqq4klE/3wgNGc/bXTD8tvrcfD3Z1sTu6FMVIqNrju+PDvdc/1I4Ybc7HKC
/UjGGs2vH6ESapQa1KWEXurj+T/Swj/HZw999MbpCcghmOaA+KCjJ1LagWoIs3E3
Yap0vPfLoiPic26Tnf/XQrcN10tDQA3cu8jJhH4yfHKceEognCwqVwxBsQD0z8Kv
ogKAc38NrFYC6bkm6AuX2uMstX+4m2emuN7kK4TP5IvBJNFnIadMNmiXcxl6tkfD
P535anYAYs0hLfrm0tvEcdzJ4a/H15nQLcZXXRzSb2t63hQiRSRo7gL6a3tbR6Gt
Y21efk6ORlUnLuw6jt68A+Ny68FrMkBucoK31ujztcNLj6nAkfQYTVe0HhoCGTxV
qQhHnLYN8Ax36xlUCOFsqB20hu/JcKtjkcg+ga5MukA8euhs7fbpqjcMqfnbcGzi
tUl+oMZrSCwpwU7tPG8eyK3xWMIA2IelnSpVwKJvywv0erFEyDvVRz2T2uTTdjhD
PjUGxAsYb4ZcLehpOdZ0R4aoCs7XlIB+P38itOJzmxOMlnH5otxytfyjoBJj8itT
QfSp8e6PtYyUksWdWNzlj+ZQFl/FaUG3DSLIdrHpqCSAtN8KO7osyX30xf0CAdtl
ac33Kd5DyzB/q50qWhY3EGHw5nva9mLxNg9EFaGOQIz8o+8gYR8HsCewCUS4e8Us
RUCXWicrZlIcZ5/zhlCIRgOJpwyDNl1YGBa+e+sX4nd5Gc4BjS2NwK43y5M53wXl
raSEszTx70S759IdibjNz3hwOMolYuJeD1EJnr6x5+QB2yPV9lo0I8gRtn7nPd0K
6J22QEDVUFWM0r7aNQgllmGyCTt0C8S3v4AQB58Ngbv+L0z5GxcmNbKixaZ432U3
BwuBeppds41Xg2WSYPlVQ8pHkm9pfFU6SX4RLoc2ZxYjK8aIEposUksyCN41SEmw
JEypBCIXSIdvbbsLk10CzUkwAMvQ/rWhHCYcoLLuP4Eh5a8kAoX15IxBX5FoQZEn
E2KSMxXlCJYdJcd5CioWLV5stGLUaiJv4YhnDDvdFBCkz6otsf/IOSpOQkwb2fum
IM10VPHEQrpWAC30kNjamBiu3JriOhCB+Cdy5T6hbWpsQH74hPUuFfJ+xcbJx9vw
EWqdxGwv8IX0viIfEuP4Ifu04itHZ2g1WKJg8tpGbAd4nSRlrPaGF4SfFt1c4JSV
ELKeZ/1YNhvkLXY4ns6BZ4xWhBBLFoLwkYFgdusMX5F6UhjRf4zRl4ljPZjDP9AW
4kCLGfXTS0WmiMlGXZKxRJBHnRdqu+lT4SyTavKvsdMuxxv/BwxiH3JTw14TLUrU
3Z+fcNsjKclY6xHPz6l1P0d9ule0pRbX7cNOjDd23ofiy/NbVm/80bgnDWVvHKMu
UAMIF+FVBngWM3tK/KHICl7nligprXtYWhsZrV3+rZEAaRjn8yaLjFlBn6Af+bk7
zTjyMUxp5d4XB0DoUVjuUYWremUZ4gXHL+Uk51DScZ+DGDR2IrZHmEaSLmhZkluq
ePe4/zaomFCGhsSLZkohXO4RMPtpaGAZ/Kms7KiwGOlwGRkSBAwKsjjYgzOkDI1S
FPLpEAGDFfxAVdxz6U5M0gFJ/W7+XHcwugITFw17ft+OHFuHFDiWlFoHkDml/E+b
AJPu54ZmBTDNle/CeF89nc7iB7T1owIsSwMDSDmAGNTvp6LvoxfuRfYCgc2jKrh3
OXntkYaGjuWU+ybwwZJFr68/Z7DecvNnKdBu4SY7jWt++kcmY0i9D9OVZ6pPadbM
q3e/0t06ncBIawMsP3XhVutEislpE38HDlkFZiIr66S67G7wRGaVL9mi+Vtjb/iY
5S+QlkdLBJbGYiHaLf4EPv4sshw5qbQcw9IN63kaR+gGrRd1bwg8ndDzKFs8msO9
zozKVKndOwKQgIQ5ToqIyJ1nEkgJjS6CRu+MuTGh+p/kHVRNi9MNL3gt7NIzcLPk
uj2iP2hn5ZINzwIsjBXxUukbZlrAr5owa2k2nJExzo6ZJ8yh+jpoSsbcmiyK70O2
IOSdFROcmk84jDv7ia8EQH2n7st8nKBA/OzAtPTp8mI4Vh7L+c6oAlCpVB9qky5I
TmIanjJrQXyMylzEmF0af2hFh4H6sA2fWvc2K2uvCa4jndUWw5QjN1lq3Ir1JrfK
IF3cGaXlFDSTs5cv+FhcY1ONAdDwRFEr8zP3xOtdVcNUwhUJmITGEqOKeAYHrSgi
6jSNAeb0JvOQoysh6rLtBgtV3z3OGPwsM2tNech6u66zphgTRkCvlyzSH8XMV2jE
0KGXKPLPuOAMUhHL2W3QQcIS9MI+ZSDem5atDJep8E1BJvPAK+r102oK/0iXSZss
S56907N19KlIr5JTe/OZDZC4w5DH/OS0Iwr+HbV3kcaq5BYGu6dI9NquYh+X2Wy0
8mpkKp1kGBfkgNSrQ0yACVyHWkdq/QCMxIAbhJRZ3DzFBPuRVx5eVj/Nynjnl7fc
JbRO+DJgG0dd575tAKDsw+SpsghIxL7p5t3CeQcGle/OuN5nY4TXdJ9xxaSw3xso
JFT3UmmXXfFqQbfbK4cfayxlb8/yyMRbQrWvNoFBeluiq9fb+slXnfZR+9Oj90wT
+k299NUU+g6T6q4vSZyDhuxSo1Zkul+nNu4N/IUYofpbqCgf+CcP7kjOBJ/Yobja
WeS5MSi4Lx/tJyabEjkiL7rgCY/IoiSXy3B+XzgFBJWgFRDdOndvW7vsC+1QbT+V
icmcN/35qe00sTOo2mzIbR8+Quwrt7mh8Daow8LCEZHEj4ALjg+RYz57a9/hLdY/
Khhhb58sRP5/HIr7K4AW2OF/N0hiqOaGoiJjkyVn/qrBzmdHf56vpOL/YvWfkV5+
UOVXJTiVVB/NWiJKMKhxF9+/UUsDTl+QbujRI1qB5w3jkCLnz1naF82kQNhUwp6/
p09BSr0boDUXqwzefh6LBycD1Mc2/D9nNcDlnq3NL5DvGN/AU8E0bOmWfli6Gbv3
hoYcl7K8Ky5onXKFIomaRf7PWzBjReF7PAyZVGAlxnrkXw3dXPv1YMIyGpzIW6d8
A42eSGBJnCS4JqD9kX7VNwKoESkJ/Q3alqez7avgnTMf3i191v++/1Bm86Lp5NlF
jnwiFmVRm//LuVkvyx+VQ8iQRkA1KNsdcX1EmvO3oH4WqLx+Ll9PMtaAWHN8p08l
EbZ3WVl3GXwFvd5dv2RoPJYEuDszVFF56aJcDJvgA6DVixtbwspRHCQjDOFCTA8z
WxAeSR6MMUQFoRrt3bvXwpXnIj3XA9LOUG3roXL43HHv6MBB3D4LVA5X2GlfbDOx
VP2In7q5Hj5RaNf4WzkRlBCAMEPEUIG4mr137JUX7cldO2UDe483T62btF6d3gV9
ksam25CsuLm47+kS9g5oHpJFPI9vV0l41XgMYW1brzR4/fQSmtd5bHFkh5L32Poj
qF5BAI7LibKhwcgxVFnQ0/P/0jueK0brY96gyXq6b7YochhXAJ9v7zfOCvKUkX7B
mBbKtrhk8AAMm3moQoOr+oEqGq3xm76kqSwYp+iT25pYXdbF9NfiYUCtqcl1Kso7
nLbKk167pU/NF/0a7768Wz91gTFGbsFBdolmK3mNGLot3NuVEGPqwuM9Rrtg0nnw
t8dgTt2cZpzozgtD48dSiD1oLMWsuIrqh8GsnwdlKnyjCIBeZt2XpUFbWRQCCEXb
YFUTO8+TYqO3opxCgk9I++dQedKxu/eEGKfFj5U1pObZlIwRDkWnkfEm5+UkIoh/
PWlScg0kpFqCct3TfBu//iKQZcU+UCws4Sw4CRX0nBywX0BRmtrA7YyWrGoYZc48
wAPFFXCLc/gNsO+XwNd1KshM/6yts86zzISrU9Qe53FUEWk8aDboR4A6VxQ8mUdH
oCCPwEywSdiMSM3VpPaqooI2gnahmuswjVTd0vvCoJlUjDEHlWJyC/567MGMR668
hiYG6uqXQKBEXE/95U5cYmZ1NJz3FgBVfI5pIFcIj0i2m/Pp/8SYyuhaM/immPqG
wYflBMDE5tY7fKwQy/n7q8Gk75K6El0qogeoJDwEy4+YbCP62Rko9mZqM0SNihts
IaJD5QFiHcFEPXXty/jsvDudm7m/9wK+ixpa6zK4tN2G8gl95m85SyPSuIcxThOd
uDNUXKd9nxxEptu7jkweXuXgEeVIg16KYBOerzTPjaB9c3lnqOcWT6Kw6QCuppmi
b5W4iT4klelxYnw7FbPTTzfVxG8Dyr/90F1mURuXnHOSzBaSFMLHEcwhi4fg/4HA
XJy+YmQEM4x8ToWH/LUlEtNvnMA5p3lAkYYvRwZljncb0ETermrojyxOuvdxv3fO
NUtdWqgl/nwSeaSz2bvDQCF9bIDhkf/D/8O22K5tYH3wy0aTy1Hqo2pLoa4BxVLu
LG5zcGfQeTvr5/1x7PqH4IJd3LLzQLQ/iIMRvw88ATgvEapypNcBRSNIxDk8Dajd
q14acko9Sxl78pP9nvLBGJSYOitH6Ile27CYBwlm7ZF/qXqH4i0xU+kfboNr11Qk
JfhFrPXByiK2KSp3mDBneePNgbAV8Q9dFDD0oPcTv/3xW1PbG4Uo0pT5ZJiVMKs6
a3meplS9NSeHV+eEeJHsAdAczrccnjPft53n5F0miDy4XsZgHOLd0fTbZO6F8Ehf
6RY2p4IB+svgNZNQgD7Qhewd/UImdZyMHqDWaelbM1hCiZUGRXHDYBSWeDO3dH9w
3mOk09y4b+/ZcQIrDWbYPBTwqXCgkvXZ4a0EMXodbfuIG5ibOQJgN5romAshCH9b
34XZR9FU8xdr/3p2mrfZ/UtKEzV9QUm8JKrDZm7SRWjQRy0LXdWvCYqiyHvCruGa
/cJrIZRAdzzfvNzWjfL/mCscpJgnKhbF8LYGSqTTX1dk9+rac0HfmtEqPivGhRqd
JpUXP3L6n3e2nDiJ/haEK38EzmngxVmPFRHBNfmWVzQ4wM/o4Jplu4zpBWlFdhRN
A2BkyG66ysHrbcH0YkA7S/2cyepjxPH5pf3gc3L+HXGlNYMR4NcnqET/lzT5j9uk
pLSuteVuJRYyAN6y2iJI7HzHY5HfmSVKvZUVF8blaoQ8faIzZNRXDNYmS1Tdr66U
GIoMRXNGD7dI7AkkEfXwLAPS4OS9L/DmdWbXb4wRqjMXf/32Z+eCzuu1aCtOciqD
RksBIsKfiNvMqIDaFeLRDf2dB01PYCjTAiBDcY/IaP2JwEwQlypr95wihwryo48R
uO8P5pU7rai4teMhL7E2YIm/r1d64TV1rguH0sH2v2SCDNHmBDrZ/ZYz+jwDmRIs
L6deSfK381OWGRQWRUbTFP2/hjoz2ZKKsvNXSkAojUipKM2NYHs5gqqf1zoVZGvW
4PBAlbgQKFH6TeDNNdDY9zYNqg0l/Lj7si8iBs1rt3m9P6cdNNkQpYXU6Pt+ME3X
bLjiENSs2MT8Zjxq3Dj0pNlm0THzWUH2IwzK8hNhtQXJXIg/0cQfaaIvz4D9oVc+
8+b2zmPR1fo/rrKZZqbajhOjNpU5mbL7SpgrWv01ZZqv2cAy4iA66EfblJkMFeD2
qlbzeZgcpYIKpj64Y/Izc9W/dhJ7iH7NHsvUFo4nGLtB2bheFT1EZeEAtiqssrEA
iQWcTwVPvaS8UNr53SYgB5+aGK6I2SWzvB1aAolwsXNxrhZmUNVEeCHmqyTj0P1T
Opbo/FLVkeqV6tnrm36FTP+TWBXVRtKYPm9F3IwCFX085telXk9jpt4UFgZHRQ1L
4fy2YI1t8A+W2P+4XJf6RaLav/RiAIBXHBj2NxL9p8kAIo/5fEdI2X94gvDTDmae
I8Sy2KkSbbSMiK3E2JI+GRGKNI85lrf5LVWRQgw1WS8HYm1JVqJdp25QScxgg3gq
oRyqa8riTK5t1ANimH3C0lXPpjyQltRNlaqJJrsahKOFAqTJEGww5A5HZdKEhwXF
1fQYc/FuRO9GulgXE75xoPTRJfsYNtxLxFnHvkfupms1SXJJw9sKvcUUYEgUQRsK
JPJi7ZJLXLE7mOtIRM2OgdUX3pxs+bGAG4n5kkD8B2QxKZtOpOG3oGHPozueFiQp
GYvDzI0s7hE4/tMDScUhiczjfqY8mFqCPkqJS28ui/WBqNuxURRPK3KGoHdLmFb7
cstFaRP6Ls7z5Ry5rxZMeUBDTkh8GQ3N4Jnlk5GwEGlrpWtS8sO0Dj3nv+QKuF68
bgyhgU6u4zzpCgipaUStgNQcbeE7W9zCFjyxErHi40Oe9kGe8wCGFjBtow41RgQH
Oz+TrhHs4gQeZ4qhZNKb6CQav8Xo0PQcxcVW8o0XoEJpByc+xr0cI+J3Md4MVo/r
LPELBFjxtFfTv3dN9P65XT7r5t8BK38M5JUwyk7sdXkwrMx4mt7Q68oa53Y/HK4W
N9TULDGnGcOpAT/hlbB1d0EKB8lSPxzrYNpxbc1aIGAGwiEvZe1iCpo2PLqescyA
EuKBPSbBKfRAwnvGoOcmcBpzfHpY0kY+PJdxkni4I1E9frqBYIN+rVKufNWeQdlv
UFv1P18sQrUDL2MJgvpmuhLEqoOo9yIxyDdicfPdSemW0jZWT+QVJzeVVo4YfezX
mfxZ7JXheQ5koW8C+GZuuMmtZ+5x8LgdJZq7k+kjADSap99GPUns3gDJ8j20PU2t
bQRuYUadlES4cQSeWZpaSDJlAmVNZ8apbz+b3qiJyj4onz0rJQZx98g5FGe/BqjM
uVxrf+zcO7WENsvads1oRoR557o4q45eR8kSVb3QAW2s8q4E2+8rh0VaSqckRWYe
7+K66DGGo2FS5og6sL8Ua0CDfF+qnHCWTsaGQStllD7yOLm5lUblRdEPqb8Z2Rzd
XA9qXg1uymFVbAUqxjtPuwVXR/Yuzoe3kA4xEZ0dCX2glQ2cc3wfWDId3NQ9A/KR
u5ZWSriBWvEZuBKCLgrIqm4IM9elDdWbKUsvI1f+1+bt5sRBbTAO+HAjMNrcjKzo
DaJ1Nn7sUjkJGYTfCyfIv8Ft2cJsqfmfx8TeUtGAFPxHWb7kGfof+mYwFYkIGjqJ
7eAAJ33RtmkNKftBT43vJdhdCNcdxzglf+aVHPXjR1j6meov03zDd5k14Hb3VT6V
ULqNLOvbPtanRuUNFr+av2MMWR+FUdDCDhdmTPdCVjO2Wdqg2NHdDpTq+JD3/9si
Xd6/xN41N22VzwGvoH6gTfe9wkYv/5611As5e1jM+3rBee2lLRec5/SWQuqjdaev
uKZpYRfsqBVxLqghLgsjvTnJ7isRQCQeGkeEcZcr3SQq+B7UNU0LZsOZOzqZk08N
qJJA6DpCN9j8/Ykyfpx8ml0esRW7PvyuE71q8u5KgOEyQZxg9s1V26lnTRKjXX8F
mxrn1S+y8QMPtYifYo2UsWSBTGO3nLAOa3gSXcthvtqm9sdXlrB9PI1Ik7ibPXoR
K85c6LX94Q8fe25NzYB6WfA3i6Ztptl7rYZF+7HbMgvrXI70B398LxYQqMY67j4/
BKCq59kSolQ4VXnc7TisrZzOjZT8lP9OG9g2nELK4FoFD3gyLL6la6oJru5obu/z
Zq5EEmQOTZRtdjFKsKDrDuQ/iZhxNREarJH5qL8qZXMoMhY0dULCqvtZ/IWMnXNj
9IWuPirT11/touOnITHbQUrh4edhE0EWB6+jOndbwPd5dSyoYFPBvyjCLhHQVKvu
K1h4/autkFpCw25UXdsbvPD5KuYzB98XnoQ6ED+ZI8ZBqzjhPOWDoxi014xBNInj
wvZLC16eOH16tuzVb/FVB1MOHQEeIEuUJhUbcBjNafBVX5zixmwxF40a+QLbfX6P
R92/BwUIQx86TFiSGJXWCrVp5iOuTst1muoIyqESl1Bgnpdnf28W5SnOj5IprmPS
im5cHcJJ/LdGz3tTbUrlFwr0GH63CMhWXBqZJvdV3hr0dLtSlur35eMSwf2bgV55
00HkL8TOXKhch+ebwulNNRF31+jt6kBrJEUrqzPbdR1YxPk/Ry5supr6nXehu7Xh
IXAyWN0yWxDVFI2laTQN1cEHxGUH8v0CQTDlRHKG+edpHO+YoHjMMOZKs23eNBrj
5zpXnN0aplQXwmApxAmM+29c3iFIMJWRvRJykOutR5+dlk/mZs7c8usIO92nVNsg
eOK2tRIEq5DS5tTn8ynWOH2G4l5Bwp+z7wd1ir8rRyeIB/jpgmVmJ5I6J2exVcF4
R9HWvvebD+xZlNV8FDJjzow6x4ak2fWpXEDvydvWinR7CA+FmxNm9/ERVa7VsI8o
s/Vu7+2d8wt/hOLFsDvjNC6WdfHqrywsiJcECXN2lt17IYFBE8fqm77tY5NC6asQ
2opKK72uMYkeSsGLgtCLOao2a/P8PT3ag+H9eSirVc6cQD4+wiETNbXa5PcurhCq
AuU2inM1/zEbMwmbtwz1FS2c+5ROK+WcpuqgKusBHtVAijcrHFmDspanIPNoyk7e
KhlKeK/E70fCE1vADYbFeHMks428J4/AueAvzu4Wzl/LL4s17RBUPw66FIPo+Jst
/1VmPfFhH9ayAzBBbQfSfpG5h9HcoOpsCGS+3mylJNTEN51Q8MkHApSCS1sZA8sT
FXHf+y9GGrNJbpk5oSElqnwvw5MBBOpyF2O7bWZCwfC6TtjiRAAd3tfy8QAfT8uz
dAPKoSwXl8nGwJMWs8ibiFpZ9BL4JQZTlrwLTORGFbBvhA1IeSfc5hzI07x4Fja2
u9CFOjElSFq1vkY47RG2A65jkec8GjIRG/69aEnxLJTSYQTJVgAsbIxL7La+IhfD
P7s7jvDHyMJk49bodq2/IJWiIhK/OzEhwdR09eVvIX8CY9lhUG7ruL+tRvtARywh
HUr4+RoSIAKP2Tqc6Mldlo2t/B57f80xdXKIjp4afdINoM0Ui83Kun2FWNUr5m/o
B/yBx7jeZaPRwnO6HHVzEa8KiXbG0/RtmZvYo9L7egDhMcJsaKILmJhRwqFm4/fb
Ux2PxwtQ66unjytLUXhsJf3ltF09Bp/p3qPfgi5EsvSvCW5WX2itH7e7hBTwuL0o
rkEmSunFdnSsorP9jipaWtAz2hVdlgql9KXX7NhKsKD9lX1YTLOuDI67f4O4q1JZ
J7FpifG1wf6EytH8TqnvsXM/VB6WW7f/xxNVtS9INzW1g/iRhC+lD70R1QJFNX/r
w4PIkfqHir4q792NNHmfesz/ZrNW+XQcz+zDiK/5trCIBkOOC08WRHszutlR0RrY
UeLbVMeASLkh6zyQID8dzMGnuyw5i3a/3A63Ul/ed8HgpRv/HV2dxshWlXpDU8U7
4t+9ZDQtdmmRZypD6e5bFoHdvR5qi48ZNr0YnyQwEWffiY13LHS49/TyhmZ7GoWY
wCR+cktjpcWVLngf3D9Ao4l/Gln71EGwJH2I/gTdLZc3mBcUd1wIgXD/5D4fJxQR
1EtvenObE0bUz7gJTo47zZSn8YbiyeIeMcDZKf0PJvGYJYhAKIJK8Jbc4dfzxhq2
hrUFM1E20CrOKOvDu3tKmcmjhaLWawoZm2hxop/XLbRHqg3nuk1a4SCNp+4+RkUI
bmhnCzkt7SO1UVL7IFdXsf6YCNG75v5CuKHgTk3ghAH125oRawSvMxyaYna2pcN+
QggDHO7g+0xlRqm53RxcedgXGGWpFUk+kMBzn6ZmE3IUsxXwQa7grDyoEjAP3B3k
jD4fszC/DC1HqrQ1VfVWia13MdD0t+1vqCiz8J7zic2w9GDBO08gZwlvVaQCCSwZ
MlXQKU3EMMkLR1hp07GN7Uwa2va2VbrT6va3R5Wok/hL7DqdTvMF7bjmFGqtKHCw
jalmhJ4nB7HuG5QB3zQGE45p729jbgr7lWnpS3X6Rc9rGgF+aLyC14Rdxwp4vx3Y
v3B4rARiffOnBnzKebg7gcXxHfETr60kTWGiSZSUMatOuCxG8M7FkIinuA5G2sNj
o4FZMMo+97ysm6XoCmmFtB6WNnecA5lTHeojHZgoyAYGaJYKtOasuvm0rnhCJkuI
0R6b8e19yivjnLAx/fM7haiHHuaOVVr16qYrBeSQqcesctTYWumTKk6no3QitJfy
YUx9dfXnH7JkpAgW8tIrxHBmFmzbZjqKHkshijRsMtPksBTR+1xs90HPEs2mEnwC
0fWts9vyrCMmH3z8lB/aucveeerszN/bDWOqm/cnVPv1DNIoUDJDb4Ja+c6/5Xw+
6VBiRA1kX6DHP5bMjGkaEB4wRaB9/s9rbKZiXBVnf8j5hpo5feWe/1PtXCIKOOMn
D90OwfsOkQeN5StrdPmwdrdTTIrED7c6xG/SAMaaqo6NCC0VbRc/tL/v2lWNMNIL
DdOIZPeA01Jx/60cx0s+PY1qYm9iWGXQdCrZAae6fIGAnNeskDCby7WQc0MRrOFE
gmKhS6JwjjbJhl9paPkOp9LMFO1H3XAmV9Re3xcWTVvd25dou6SKYXO5mVDCroSI
YEr/tsub+isaWiKPKylnO7hbzNcoi8w56/O8VwoJi2eTHQVmiOnU1clwPsxWoius
BgfbFZEyU2/VHRvnv+3aEQsYeJP9KwKQzmTmGDOhUNkNwIIfF3K6UK4f9GJia9vJ
ZXVkT6fJH82VRlSc0ESOKWVFbYL/3rQoUnC9YTnEJcNlYMI+3g8dHwbcGXfnhFNg
qLYZfJKsN28L7M1JUNqC87HKMgq3MZM6AsculaIj6U20TeLs35tzANHdDHQ1wvjS
56lGTajnJpAgElHlk7MH56x9yq7uidfA73E7RqImK7ZPgWXZ3s6vQctefBeQl/Dx
SiOmtgvkF+XhbjhTFweTo0P2SGQfCsS4Cj02TISUWNNHVxDHtl+TVBmvKzw/rNbW
AceG0+0IOq6jsq6YwoVXoor5bmCb8CFM9KDrsU8dgTa2b91xEBPfW0oa+ejLBnfw
iiB6xOID68aPPZtKB5qbhdaIAprdHuWKS83QCQZ6Il0HisbG/+QBsmRKK6Hi8wqq
kxPh+LcFvPCzZA12VlXZRc+vsg8l9H1gzHHFN/dux4MUG+qUb2aTVxzU6WBoWHSm
bjrSmjoxVuQCqyVUMC1YAOo1aILmoZUjg4rXCH4ijWoN6c5uxnKnGnhiVlomTNSb
9on64/upUmEFQTZQwFLTUkyqXdx/hj6/M2V7YsGpZpcTziWOkYBvnq6uKS6hYtI8
HCu3kCcC8NnTnHmJhaaorDZM+Px5VCl/dGi6UQ68W1vcupW/jcDoauu0vW8Xfp2A
/y5++ojUhS/L8gQrEulcF/GoBj3AZyg9rc5tw7KL3n9E3TgcYtUQBYqt5cjwfmdf
Wpa9MXdLSnu/S4djTAkzC39hW9q0S8nr+HQx3ZfrTCp9dlbdmCZjPWwgX2gsRtwl
mUKMdRRxuy4HqQ0795Iy6RdXpLT7vWWSLnODE0+uZnQF2yZo5ZjoKRiSdBB4LQCW
i2kBV6+ZKd2pZ4aCGJIeeZ3ifXm4KDi9qMC5FFxSRpJyKngxyxFThad8KGdm2Jhr
cDQiPHLvXdd//miN5KVP88oePGXdCqKp4n5AF+yZsl05QlXWjnf/AhL2yjRZHPdZ
ysOcNRny6+O7Mkh8pHnwBkevYEaaxeP1F0EA+fGBrDuo/KGZGScR3RfNimSd3lzU
4Am7AdBKyX0bQdNTUVX4Ub7R8olVgTF7ZcV2elNQBU3wCAQXZC4FMDD1U2yjZDRE
Di2dfl67jktPSlUo68xD78pmGvq9XC6jQsuf+iE4OlAfoc83lb3hNOl02oyUnlEE
a6CPf0Xma7P/5qcmBTjySPAAwPLXrqaMI2yZ7x0QHgK1ePjqcQD8/Mkh1lJ+ZxYF
lO2vM6LA5bx81jOpG8CYox0VfihSSl8D6wm84q8rb3XmzEz0OiLf3grFOUOeRs2J
tcOFU2u51Ox7YbiSvjRAOvSK3N5G3VvGW7VK9LQ3pZNMXutmJp0weltz0Dep9EnJ
T293kcOOVYVI7rtf5aEbSm2vEX5SjH86OpeLFpGFwfEbiXdglPRG7H7OjNdPk7QC
vJe2o7XcZB7EfAt91z05qwVivzHcrqOgWYxxE8ptM5pJclvbwY9HgpXOvqZkOtNa
YsYTr5mee47UbDtrSW7FZr6bAOuqOYlvzaFR4ls7CxnYVwv4MW1uHh/QFRrJNMGF
csnjlfXAsGb+ZYQaVi4l137qmVnM4TI/34ARLBgOHIYlOpK1r0p2tjvEi2P60v7j
vnJQ/OzL+Q5YItZdFDd79sWAE+gnDmJt1ZcpxE4YlfvBGM4cM1X3is1sUGn8FvBY
8eedU34iK/nXvmrFjGNtZjgSapbsLGdg5L8j7yV+Hmhs3QBL/6arLk/HSvmPJef6
IAkqEEwes081J0ONAthQBic1QwhjwC9Fp1myF3GmzWb9k1HOptrGsf42/oqk8+4O
E05t+KTorIpUDp6Nvhj0Dca57aYdfJRiOF6GT64atLtkUeY2JI1KwfxKF5I3fdWh
BMn0QKwQRIfhO9l2f3JD5+I9r2a2NhNGKjyNMx6/TrRhPk8CeVYFpBPd5CZvTurr
vDBQFJzitSB3VtxfznNrpbNXPifeLKwbIIMs/EVioLMI86AYx1scmfYBKWbl+d2v
P6D7a9vnNJBYukxnVKPHxgm7Wv0Ex3lbioBT+9HbZqwepWCa5qWizo6NAUKVRgKh
DRRzgOYPeMLUjeOdRvQKZyPCXtz/VjSi1qzN7jLVI8AfFWFedvOnLlptbcC6UOYi
Q4as8MpPxxNOb1BxyTs9DK1McZS6RdHWa7NJuOe6JjKhPqAWjvER6JJvN5kNAFb3
vi4y2OyKQKoIIGcsXEwRFHSrHgOsLv3mHjbSA7uA/J+RNB25IycORooH3QTRQ98p
rvgqUr6KNZVkDhYQ/LwRT3I291Kzf5nMngf+mUOzlEZxc3m9EbPZhACz/yCbvbtG
5nXgtrNBif4TLQqC6zcCVUtqS0oQXCcSBDvUwu9Ia1Xx8YNYu7B6dGcHiSnhajSn
24KZkpTJBxsjnned1slXjtyzNUpH0mv4CrLZgX3m51JsBls3GVlMd1fKnMuPwI76
RjctcfX68MzgE5b50e0w/myTkEKuj+pVY9yYFulmsCZEbP0pXRaZ0B/eSEmiygz5
o+OdGxS+XzAPPKAAnzYruH+okz7RB3jLsXgRlfbOj8rgT8ACTzLH4i/gGHUMlikK
4UAaoaeJbmKl8jywBOiGYJnWcucviPpmP0aEVqcseiAeJUe1j+LeKCQkFSXMCCdI
bgKf5fYWX3ulIpFU8WaOEcPE1Gi/bDglziV3TPfh66ZTpRk2NkOYAkZ+dZR+sdEf
B/PyGJv8yNKG54qvVk8Qa1P4xE26gZhyqZGkXe7SUI95eN5tE6pzrRcN0C54IBgJ
N+so+NPA9FSL5TwKc0/7zUYMguxl441n16TeUD3CmWlH/mucf2gPmAZQgK0h+U50
PTkMKtAszOApJQaf7w3pm7xoIIRDYSpFZIHJ6TypeCGl0Sc+SsKgNFnwTPjP3Om1
QFK1XN/IH82JIz/w+uiqQn2p1z9dLvSn9uFv2/fEK/jAhLO55M+gfButI8ZXCB9N
zS4/gNPrAFK3fHQmofoM5npohT1asXZv6qyedPLxT6In9nSkn/Gs4RHo5AW54Eax
J8yepdW9Hp3oCSh0M8Y/AfO2dCPoXJiEjXKaAk0iEGGQdm7xAU8Lzn0uUW3gGsS5
2DtNfkdE15WeqVrfLSEHBlo1YbV1eH3LNfPET2xOFSM9aSBhFyP8jxOEygFZ9rSW
sA6FJyKoTW7BuJC/WXFpQUfPoN/AyEOhshjD0XVbDeYlQ8MkQVimHLvEKFi6G/fj
RI2ljRZrLs57m98RSWqQ0BiwsbfkVwaCnidYaWBL75LYZeZETCyyxYGq9lzrLbQV
J2ivreR8p82akHeuT/BW6eoRUsdhV9Wuxcm2Pei//av8UbVdzE6rtuh6rM9uN4Xy
nDgmlEo4lDKV47IiICF9Jjz2E9UZVgAr3MyfdxmG1GES6YhCHhvI0d+cB2er4pHT
IGEgjVS1GM0GhB4lXBHn1SrDaiPc0YdSmBOsJdEsyX78vHFckPai+ZhSGy2PdXxE
alk0E+D8yF9H1SiPSaTPO8YClPf/7Aj/8TuOSfJOJNZ4mG5DSS9zX/w+exOmECSH
l+3HOpG7WnSUuB3wuZlYnhvsilbQSMXiXmbmYVF7pvLFKIbmffe6rF/u78rCoIA5
8WtQ5Z2M5svbftgccwF+YtW1TvWgIiaKlm15bsuRWtn/wan4adiwMGyROjmqBrjo
xySs10EERELf95xZRdAU0qvaXUY0tB/91zRn0bIFdKT6HWS7czxV6Y+9epQj6+kb
nic7WOXrkWQkyo+R5vCNx1TnIEn0M7uqHiA5w7k5FJShP2M9QbcQHhQPjoZJJGOi
VVuk8mvRf88if0vkhP8Y5InK6/cNhGO7H0LnC/qzV2B0P38x1z+QZgWWhwyr0spT
za7ICNlPYBl3F9t/ws/F8b9gWbcXXG6SnmAFh1Ybivyf2TdDJ0aw+VhZui2J8pax
yquPdXysxg0rs9izXsdLLh5+36PsfeaNGDrlv5Wxwwma0/RWes0KoatUjg8flK5n
ZjZqvorPHpICy6pb7a8iT02cZX+3ctiozTm+x4AFHOrWdNn/YTXckSahljEEiyDM
HhpDnVeA3i7/8dGyYPzFawBqXmeNrJRvx3nUngimC4q5xBys5k/Znxmr6jAcebLS
IiBVd8s4dOZd3hvtv70rP5aqZL1Y1EsvLS6uL1hHI/ikKKglsyjg8KYpTtumZHMZ
Xx9+NiXoOWR5vAgOoGBLdW+rs7q5s0WB1m1zz3p33obYp86yDTKG+jbOC/Kck9zO
ihR91V2bOFe+itpJnluyPKPxeHUTR/c3kJbZ5hCiuHruipF3u9JUKyQr9aToqYiR
vCqvl9bvYecUGbkXo/bwcMJfPBPDp4nu6Ky5G9Kdp1C9oNzgU99npLDJ/epTzjQW
dVFKNHS3Qg0ZbGbhEFLiq0b5w74sDXeXVir3vqnCLOkH7BXfEaf1f56WkGEQLWPn
n5IB0sXd3jjaS2IID36amX3ZbLN8h3LirA1rcabK93WUL/WAIlcToRXKpRxGECCD
/F/ysSZuk+ZaO+xOq9vV37saDRT5pGOsl/Zzb8nwkqnxr4G4ayLUHqnyyEbnRB3D
EhreXsIMskuVqtOeFV1mmHSF8Wgp2ssHXkCwBV5dmZs+vvaiqDJHyU8ZEOyNOfzJ
8Z0mXCCp7udTQLlTHanBBsL9nQpVGjUYfJB5r1WiOYnq6/Cpemsx3RXgXAZv4DFt
nDA58gAd6FJVmg+r+mycR0U4h3xJL3nvEoPiL6wiRP/AO8SFPX4OKShAx4JGnbZi
YR1ZOkWb6UlC0EwIWbUmQ+D5Kbt+rat7YvWnbWxYQ7th8cDitjl1NNBjPXzdCR13
WpcbV57JJek+xyeV7bXyejBXDAWEOrWIJrfVC03dQ4Lbjn/yTKpLV4g7XSfFdSnH
SnTKC04bvfvP+e93gGVkIiffIbhqj/BVtQZjYyymWPP94unjAB93QQVF6qgDmdiN
+YOB365b+3hEpM7mGqmoVMPyuTq3k9F1Gbo6WhHjvXV9qIL/vDDnm0QUivWsVtKb
T2Vq/b5xrW/ZmN2gAuLzIKAOwcNgKh1lsWO9mldX3i/UPMV4HqIYYsdqxK/TY/bn
lAEz+cUd2KeruEAkugmBYvBghTMzVYubrkihoCoVDkqsK/1k0//HtIFNFDfmlI8J
AhzmeAGE3H3qTsVBgm0S0ust4Xu8l3bThWcD7IiEAp6I0w+BTqrpDSztxw50JWPn
FmT54tBRpDmcQwYPk0ImibcZ+GB5UeodYZip+fWXRy0onWJjRS2NJmY1VbdBfe45
CQBkh6+axt+xZfHW8OLAAmBJRAAbwg+jmg4m/X9JxMAPJUW06ayIl803aCGdzPWe
uVXZapauOnyP4YSlfDjdAp09NSwPuRNlHd5rYDl5Li7UdSX1Ef+83F4gAn/HWQtT
FgvWfui/Qurh46dvgmeGEjipFFxSffrHmNHTq/i02B2ap6Xa608XWVbEsuvIhsig
v4PFfxP7lRshh5wV6ay0ojtnCp1+l+5GKMHUcXImyg082B8IGF/vASaSXuWdzG1g
eOD++kQP2zfR61c+Ebvl8XUxKUvUqlYDPnn0o5++SM3DYN7DTTNmZNecsKqM0TG/
2bHklmd79OR91hkO759aQLu4X7YEgSqjRdhKtuV2AAZZhgL5LmtWO9xXrq/TTf/K
qfux1+QB2GpHrm8sVZmWwQYILb5YfPF8nkV5rV1G4ikcENSKRQx2XJATen0Os9jh
UtwoSXn91V4A1n9GMacasCe/VQh4bjhc+Hgpx1wX0UH+P1LeAYbIThkJ1MisSvaW
UmZ1MJfcUSu2/2lD42NfkNcAM6hHr8Zt5V92s65Pl7gn4kotDUnlviV/Img43A0d
yhcH+qxt0/QrlTyfewdO0eRuyO962U93redJjpLxpNlYnkzGAl3cRdbK24i6ckZJ
rz7Wuhhk78m4BIMhDzwNWJ+wvTGgpT6XzgZu6OPRHroc9CaR87Q90rj3BwvpAoe5
QCzI6F2qxOEwPprWCAVdFpCa95If3OSmgGqn7UTgM9GuBeXTWmXn2OPGKYZzkzXZ
HjM9UfPHPTbQCmCgWYPafy9QVdpYKNejjCGiRLJTPb3oBwAIHhtFvi9sD/qbklls
oHBZBPIfcAaZj5J/wiwiT3LFB19CWgZ0cAyDAqEnaJocDhZMERn2Zc+0Ml6Q5h52
BxE/fZp4+9ZBuTe24Bg1BywFUM59RdnnJ4N/FKDmV6EzxaxFWByS8UbEjsGpa9+3
s4QpiD+7eV7Pwe7+Cv1UfjYkVWH9oMpGdL0N4kgLJegeAwfINVHe1Zy1IJguoWJc
e6puOESDKHc5PXTW/FJYQN3tW2m+apWWPmrZM1vm23Ws/wpZem+SiiZo0jK2kZV/
FUSnkWNM5ZKUA+Nmt0RHRpWLb+bGr5gaBYoTVNwU0qmdz6yB1vIiZNJjoftLCmKA
mNjebWl1qwoLrAxbifSxwM1c+5igZSZ4UnedRrCD4ayqbSuaNfnAROxCOOwIgjhh
euyEPpvY2Jvp0/r0hfSMls6dQGRkada3zU5nGCJmO4jLaxY3qc/y2plUceYx+Zm5
r78lVAJvxEJ8pYjDnf1235fbjhNBRifBWu7Pi8xSNpMO8N5PyUClHF6m/qta0ezW
R2tMCnTZRpFmi45PlWfCZozKQIxqamBf+Ndr5dYhMPkxfhzklXjZ8JhQn8mfTpLX
QHbXpVgAvPRkQZVm2vLHdy5uXfcHq1o9fw0WYNp5gwjYA73W8GJ7G8pJtC/kjmOb
ucSYeo97RKZeO0irT97uSSqMdkn3jmVjwf2nQEtQuM84KKgkYFNPqbD2LC8dMPER
dYRynGxn9sTTFIZRMAIyTw3r4DE4cJnZniP/qWVwAtUvOtzmRpP+yk3EHMbHZIZ2
IMLTPk3E9uYmT4OiJHCbvGoYFa1GEmYMlOprYHN8Dfnnu99vU8X9EywSD5EpRvDn
sh6bMEyCO8eMLZ2ARE9L6TwisS0Anai0u3hRHp3xfZZwyLsvPKpv+usktNr1ozCi
ZIlC0prGoSYXmLkhx0GQ/VmCT6rqYA7KEydgcxNMgokrX8njjVfxU0cZ2uym19Jx
VWnZKXy75LqFO9/sjxNfxKRIpgZObhIsRpQhvmtrDtsQGK3wnKWTa5iSr46kh7DC
Qk1arzmwwKBNY6MUeUXf8Vs/qg9o9cD/iN/56pRJJZjfj3bvy3MzVbCvArz0xLsm
ME5p8N3saS/g898FFukyhRJBitwYQ9jludUqhbnmO5IoNPjNsVlKHKToUAs/OgE0
eEuKmkSIa/8d/sMqxtxbV3HqD6nwp3Ql1kzB5MNkUXLRMgqQqZGtc+ATEDKMTmLS
zUCkXVgIBESV7lX2W/3mu16Sg0EjtXW98ucEs6tF0xtrEvPxJ1IWx8Rzv9tpH2oL
pXP1/BY60iJJ1ozXDUdo7XEKrTNkSDfqNKwPO/MnsBE3v24rrDm5ZEFedmzwFPU8
UlGqAgL2KjsNQ2gVN/jCjso7lwRO0ee2pORUSu9ycRy+8zreV1/ez0lGXlDOSbAb
3ADkAayTMU4oFAW7MJ19FgL13zxoa1oAJ0Ft+2g4ZfCNlJS3q5gNrs+br1ZqIP3l
7pD4lmXp4PxIm7RVENE7jdgfFlOV8wWZsO5iQ1alrug079ksq2B/AkFIW8GOS/et
PYLuvOkzED22Pg+iY5JvnJ9atgwJLxOgU/kuWF+NVoq88XZg3Bkvp8YumCJ1EIT8
LBcOsiBwgcBiGMFCqBUNqu4ivqKy3gmgXSQ27ZWU4aKUwbNTzEVy5kkGuJRMnv4O
3sOksNZ5j84iJwKaieRErMYC4sDGqdyAIuNkwTL8zqyC7U6i6fwlOBNBX76g1HV9
mBt36uCyNBjw6P+nJdGiok+f1zOAwo7Lav8U86kErHC4rXSV35Yb8OKwK1WCC/aI
9y/6n9dEr1zGGkOW8c1kHOeKlANgtCkFZg2LOdVJ8uza7t1YqdrJk6zYM0Ni6jGI
9NT1Q/IBeQHOLKbME1+CO7CUzBheHix6+vqJphQ5xZEf55fVJR/Z0V3kiVsZpnFM
vrq3dzaBpRC8Tv4+6NQhreHKY8WBFvo0RxvJYdGpc1YCNC4pjlOy7u/v9SgfRGbP
uSeqCT9aB/qrniNK7audNPOH456yfVrjUEf5duwmCKov31YJ86GgcCCGbwG3EPZ4
YH0Qa1EtGlxx6JonCjd1pyQWy+/25vzsXgvXhYVIJIwL7oxaT+2vcYJ91X30Xp/2
Z/I+RbY28Py0MYGvbLKF0jex1bMfLMURg13UIVurU8IVKCZwnu0dRQDKUelUmaHg
iQOift0V6OA/VCeEC+gMVBXRZM8WhRvDalJeekBqAvDZZUfP842Ms5xoJ9Q7r83h
Ww133HgO1K50gZVA/8U11hVhXqt9Vm6VoU29I17lFw8kbQzyeeelOECTM8DJyc9I
PoZPa5GROvnApfaovmbKwd2t8FdEPcZc9BT03TNUvNEFm9RnEJYvCBDSPT39DQT/
OQPsOapO/uF5rEVZyfqu+FELbu3398cYYqPTde5BVWTNsuuczdEaN2SQo/1EtMTh
gWZhLuQDYDo6aO/6kdoj+md5oq6CObUdd7ug69fUJY5+j0Mrlg71H7L71VzJlRJ4
RxEvZTjcnKv1wGkLd0/6yQ2/To+UuyjVVieLuAQVMDT0koBsUgAywc1ljDbZ2AkG
5xkBd7+LxRUQuA6ln0+YKlyVp8oDZXrdgS14YYjAK+GNqK/zJvAM3PcdxC2LC49G
UvsdpdHi5ii5idHERgKpnLNcJo9FJ7NS1y66BalQJDgGMKqcVYvkYa/In206juF9
5cw76JN4LS3PT2WmHyhH0z0Nscgsj4i1JdVVTVIGTI4ysmoN2ONmTqWd3NXLrmwq
GaCN6D583CjEa/aprb2uPk3E9UczkKLO5g2hJaVj8LXhsmyO9dKaqfhC5cLFp8Fz
UZSgLJ+8dNDU23OhMnT3oKMFJhCuoELa0DijiSS1oCbiGchJd8P6v0ucxjyatIAH
9IvRbTlW+Vpqn1XGQNbhA31AZsN3rA3mH9LjE1MODWzkqra+PXqceIBKVnDI0OQ0
7M7fQ3j3TJCE/w1qwJdi1mkHNL3pq2cFbmsIEu/4LYkkJ5Q0DoRkfbZHhyR8aaSC
8VAWgteWu/aWzi49RCpvEb5jAsbQ5BGHyxJiEkp+Hf6GZJN0A3KZ1IPZt4dc7bOo
sbu8cFjXwblGiHDq5mY3LqVZ6XeV52mgILrzb12h+K2++tjD54RktcS9ZGcZeYl3
dNK2ZtXRFS443Jv65CbfxMakK/hiSBZ3bzRFkykbiNfwaDwG9AUSmQh7fvZ/qWkL
LB4Q/4KWore94+pCsM4AwF5FmN7WYcjDmwsaejlf3D5HllRkGdzS0YmPQcZe+X2s
22ubi1f5fcxG/xvBb4kMxxDTcZVMq+tktHmU8KVztK7aV4thxHW5d3FhSs8XWVIk
2J5loQvJ91ZqSYNqjjgS5ihfCW4RNNJVoHSw3G9+s9zhljKoy2K1yBK68mo++iJ4
m+k62yG8MddDg0yNTnP8jnyAkLcxzQcajw5I/Yg/md0GVFp60NKFc5IELPyYgbSP
YbJwhEQT5VWDCkBrcXky4nwkmIdklQKtgwJOizCaiGcCFUzuIpqKEFuP9eYXdxcL
Wjr52uUNvwyRExknyGQ872MuPPmT7Ntn/nFlphjNch4cKEq5KRUCQ7CXU12gv39G
z4/KHmUREVu6txudRcjVUdCtrqQAvOciiuJkA23eqGAqkwmWrIsAo3qhY0rrxNwa
8n0hirXxjKryMd5fECJyRfbhIGkIaFK19sgGF4VduFPtlzIT3ZNcCaf2Z4BmzK0J
Cd2EtTZTq9yetd3JXUqpYpbvgiCv0YEEfwEs0mSHMPsMMu98IP3dBeNjyl9/8w4J
yWFjsmkSgFws3lt84F8zZKpbNKRiM0ukRDZgLZ9xsaqiGXi7nNqG0SAVNr2UJRQO
pKC5pug1t69nH9hABcgkEhy3aLzy97eAhbvddHShc3ZPokc9xsd1jq4aVZzetdsB
qIJk9UZLDZYArZwyn4V325CiwGApgOVaQNA4rJEo+mOtsxSeaj+LAEKe1N8Cg26U
rBQdjZkf4lHQbdslSIQj7FDTLE1E69eAccJwlZ5cza7DhD7i0vxL/P3PDESKrCJu
h8Hszeolk7xq8CghNCeZ+hXKM8qfIAEnvD74rQrOXGcBO3bIygCXAvZqnwLzckWI
ILrjKZS4YvvfDkCoqqGFS+QywVAimUS3QbQ9KoFoXsBOG8I95bgnLX2h3EYIGXrN
kIIepEaT1e7a8oGMVJF5Tjjlfqx38gIR/I4phfROvUsEiV7ei+yugebUMVTcWblc
AXuKn6ajE4tjYKbLRNQRMS9zqtUSgfc+9wHpPbgqt5PwcUzGH7l+82JZxPgm2DPi
nA606vY3koCOBjU6QQkTFb4pu0esBgDULUG66acBGNrbthKOQOacOapBUIKkkoRW
I/7ZPGAvXQI7rThTwDlDPLiAvKFMEYEwpPRkXX1VBBBSAaMlQmC6vW93UPNhlei+
I9BHWtWzjlrL1TXl+xQ8AUoBsPobGn3v8Og/bSKrY2tb2/f/Xp50WZ6+O+q9ZdQM
dcDqfnDwm154MpfIuQIv10WBpDN+IHHYw/JQn6zL7KK9+zqSK37dFMCplGzhTybg
C8BJ3nAA9RpwpnNHllp3wuRKY2GvJ6qXSVfa3M9/abnOwelrejihLlXEqbjJAS4D
huVadLaFyeBKazRS+r+TMhkimLaFAY9NgfCiSIoZ9BrTiviKZ10GFWEFXcPwrsGz
+wDIrZQeZtnvF7oBHb/9+RWpdtmBoZDRLL5l40zKpDWdie6xrLKRtQb4fU/2S8rb
TSKXIFbSf3EYROLkap9ZrkxQJ1sRpLpiZxjy9Mfwa2gV5E3uhrrbfr9dISkeb8SL
PpmkULlHkO7Duc644sugZdbBkVQjLAsky7PGBJaH5pWmkkAfn540EpKwtMAFpBNN
OJZ0h2rJgbfqwjPlpEFsQ1ZK8zYWSfhx4fLVeGxNhSQ663bbIh+1jitRPMV3KoYN
Ma82xre4xdDI/FYDFrzHbAoEcr3znLplIGiZiysrWOrsOTKEk92Xl7teCa4qZpoX
oFssnFIFfAvcjOcqpYRNGRpxADALBoYk8YBN2erOZLaHNkgadhF2pbcEufpFm6vW
TC53OIdMxTLqncvH8iT2ERhpsPGhOZ+q6nw0jQ/Kp+iK3sHNfg5fDJi7slCOe4MD
7Zrn/ueR8Zfh1cITlGLSlaOej20OTYgJB+56LLxxwba9D37H271s2UXI3tM/o/yC
jSHy98n+4fCgzXJxW/NKxEtb5iu1Elka4q7l1/LW71rRmdcRE9fIfbJTiAtwGfJ1
FKMY4a7cmihwfFktmPc+yz0Gc+ff6qzeujzC2jmCuFP/liRsRgn0aL3nPxDiT4TL
PgLOTvYqHo9uNdF/PGunhWLaY8pMD5iRNXg5O5HbuWu+lEcUSj8vliPAB2o3nPlr
HpkQnxeXMxBc+g1TFkv+N76AIB8wccPgwTiRE6z22uf7KiTWrcpGmSC5aSj3t+QJ
VHCMno2ZpsCMxeseg8s4CImyDkInYznRn5Xw+iY09tIIlb11bHxK4nZs4yWJ9z+t
W+40Bml1GhzHx4ZJ71kB8dnDNRGPm4GNfIdFPlAu2s79HSy+auEWTRdeq3EdOXoK
aB6uQSj4/6Pnvp5V0hXVu3KPPGruN9ZcmbwjhOnYlWVP1uquERgwxaxC1JdTbtYI
cSfvTBAlmyoHIUC7rTQYNj5lqy6/SRJJSoKdjFxmlEjBnvb0xp6dOpCBZr5+QUxz
yixP3Ieda/mqyvMG5qUUEmMBWvpf1Lj99Vjjy9hLkQ6eUa2B1AQRl+hSOSdZZAKH
aKejOuuYdFRrJuAgMZtKovY43PgRKJmnPY7QhZTlzQSgq/T0N2rPBLHBiNtHEZ9z
8UuOKc2wvUeTnMmrvy/ez7FqP3qMUVMt3bo5fNVGVg0Lzyo2i4O0FvyxJG7O4qM2
7dSNte1SYdcHWEZMq7LAYT7gka/XLkfCN27WZ2glaBHkBZdY/J26p5GN1p/xy2v9
beggbD105J6ctQKrga4vd8slfYUjJWGeI6pmnpGtPZlfRdU0g91vAaaFSvigCM7+
qfXdi3XHVifF7qZ8EL10MX6rMxb+MLkrdojtceI5Z51w8fVRdqGPS8Xnzf1/tvjc
aTPImDQQ3Awzzy0suOPIPS3UzIAwjJtIlor2SnfQqPNcw/O+NuUKNpHPIbrIBjQG
Yq7rbSi7zR21XXxN80n4cG6VRLwSYrazpvy+w6ge8jJxZYrYzlX/bNV9cjwfdlsM
kbfmcvZcYrtJWEOgM/L6lit6bQkN46Y9y3l1DUZ00k7WUYuA48OCDph/CMv9RMJA
AzdSp0UYiVovuCdAabVfUTJlUnEIJYjC+WTwMi2H5P7qECEWIjaf37t1WKP9pbnW
67ML7Adm5yaO6z2+fliU+Mb+2EFNujc7S+o12hlOuLNdbpO368aol+ci0pmG9okB
viK8FsbQa1k7N27z0S9PbeaD0vxSq7TUvsTV3N/CLGOX7I/991SHxBmx+EA+zwc3
9da07WaHT2Io7ULKbEyghkEho+z8hctB0NHB6NhFS6PEoApbY36C8n5tTTP7iPMX
6v8ubCadz3C/DS95QZBtiDTjjWxbeyPGMzaXO5KU7IZo00DF06Nf75Q/wphxbRF/
JE4ofkGCMALTE959NZG46drofil7CRZFWVXnh9G28mvifdODQC7tE3OF/AabmYqf
T6X/gCLAWEIVfxLAiprvx+W0SH1Yb8IOKoI2WWe95X4tzaxXzTHFaoANd8QENF9v
JVsevkKT056v2VgUKcDoFPbowEOytXp4tL/BEP9eYVuZK94O8/xpjDqM69dOutzr
SXwB/W58X2T79fa8/ZlqXB4tQN76SvZEspxwxHlVjojMFFvbDCHJcAoT8OLBFs4l
I5D3esBOVvodcMW6WCTWAKEsI/sgIQrmcMuM9junGpHuitZvRf5cDQopQNWYwaD/
F+C1SnZVzKIl1jN215eMl2gfK6PABG5dvZpW8mUlx1z2nBBI+FTbbWDWUOPq1chA
lskfsdhziy0h1hHnyPnKq8P/8PRsiiZDNhIOtoGO+0P23MIKzF/Wn1tvxZ/MzLRD
CJfymdqD+YyriomvigNjqYVhWLMJcjrV9FdFewOH9wG3Xr53jG1quSfDaIlES8Ut
asCVAqbGgZ4JDftR6u6x7s8ZpLq7ZRtv5tGlRXnV5eN7GcmavDt9Q+gr/RHqvAT3
ZfTm/CuTJoIWjJ3TqKj+NFLfZxvez4lphpTQYQNYUkna4gfhzBh35LUwFXOPz9DO
9cjUrmDNKV4xiTvPyaGACuKEFEX+SoZPummTLNn4sj6qQqEbmoqXWI6wtPb7nxdZ
N6z1QiQQyN+xExns6GqFxRhIsTX/Ahkhv9jmaXPdwOUfRoao6LWmJQ0KnP4E/ODO
0YDnz4l3wdhK9SBb2HM6y0HD/rO9dXa1c8aVdhihiExAC6KdcEzBssVm6vpUZvLJ
NTlwjeXhC/Je48RR6fu3ZV3t2ZFGoZzREzi96ryJFoi/yom5i5sFTjHwR6/aWwyZ
2vv2FXQButabNaOzjh5hu2G6oR3a2P8Mwa1+mxD17aQZCft0m4818tvZuOS3Kbj9
dwVsnZhQosR9R9iYsCTi7Z75RjgGmuZ62CGIeOvKyN+pS+tD0MZVJSV+vQ8+8ovs
Df0sMNvNEuNzAL2YJu6caCc6FT7EI+IX1daW+OawcbscplObO7BaV6GoovzWONe7
U9FYgVsPWbuaYXCURsV2ZeYaBjU0gkyJgtME0YRwmudgweQf+w1DyssXgQ6XZsty
NPuf1VtTWaZm4Nz4SCFuLe4G/iYNFgIW5dxTmwc3gdPn3h7XtzAD4tpV8sn4Aze+
8XYtkgILwu/vH53xAFyOC7q42sbRv/qO/xdbrAXT5Y7SpOhZqL3SvEipxTNbSf1m
tu6l+57/XzddPkMYlqpPsuKZvKWtpwUVVmRGtSBAMym8opp5PAYJclAOK7wHYOzC
v/TnrTwA9Zkov086qNwnnhMkhkvTLevxmZ76P/IiqQrPgSCIF8ZLdLlZXZ+iiKOr
2UVp9FK8+7XJ13sGa+n8uue9oR2aaembcVswPyiVpEIuIHdwfDuAbKZ7Ut1yHQKP
THRdKyQvT5/kErp1x1lBY/K6brKZrUSivr3awWtKk1/fzjqEAvViAgpaMuSy4Y25
l3Dz1pFSrhqycxLRKV/TesjhKAhN6SfljkSt1nLRyAoSjeyMhBZhUS/lRW81dOUa
9BRoRKGSYb0Dt7OxEmtztJg+FOGzd90W7GYqmShUWcvz/c7oLkCP5CmaX1yuM09v
r2wOmZGEXtZQVW1FTyMakCWyeLNSplgTK40n9senNuH2n5CsZ4gFgye3FHdQVol7
IF7ZzOgxp6OZBXKueQ1tLNhslSQ2Kc3k0Np/Uxlg3W9K/o/8TsyQJ2gIVkzdg1fE
iX/btQLk7tgXsPr0yaLqO66ChJGS/ULrCJ3BViGPxFLIfuVjOD0pBWWF3gugX0rI
ylBvIjxQvFLi33JhXgkfBHC2JvMBrgyCH9KxeHoZi2pY30YhyMlf8eDRKPH+bqFX
L6tWT4Oh0pqQtgrEZAWD/ZwtiONU2M+ca76AzdA5p+OPQ7cvu7yqhmuyIOOL0scT
ADoYAJXCScNHuztrDQCewQkCPzSpATxzlyAQZqkQBBikW5ipW1jI/ZgrJHAvkGwQ
NbxyAs96vfUb2X2eg4D4gkYAC9AldbfMa8HvqHcGBE9jJy1QkAx2VvkJV4rRjydS
wDxT97FUn+jxZqFuu7cRHiw5B99JMwcagsBjtQShnwjSFf8f3TZbVPA1zgGLwYjZ
5u0DgHMaDlBdENOgcEo4jhGszV+MjIvN1JarJytu7KOHWcjbTe4I08hU5EPwnqa5
uRtyyCzvWVxADpoW+UNGIKaKH5O835hR2izpPNmjDQEGx0uvAZMIO2qg4Ha8+OGp
9Db88Pbll2LiZfw15fvaH8U9vbN9k5l7VbFJL/QS6/x3T9C3azbKRa/uRZp/KWpD
dyhY51G3TOD88MZf6hHAwGKgz3TcPbV0mb5GdksrlOycW9RnJL4gkV4hTLa6OvLP
/royrluqUpLsxliMoVL0d1cL9d/Ve/kWxdTDwiFn/HrrM9+YBL6rz2Gfs/2muxIU
wXqRhQjMeUQ7oC1IUHRcGrG9gUMvT9Eh3N9/AWtu/MqRJ/M3xyPY25vhucvjZ5L8
K7L3UPTBZwCEwe1fCMGo24YRA8jI8fGob6gM1HMAtopfsZpZeutIg4X3GKj5uS1e
QK2BT7ASlxIErpylvPs0IghgQSs0A4j4FEkJ3IjXWTrS7t/yEhNEvFKst2jaNDh9
BwfE+L9zOBFy/qdEjTnVoT6qwjm+InXJZvkzoONoH/9HipZzDNji1rCBGX4/Fw1Y
c9j/vvgQqM6b7bxZ6V1Us327dG/5CljdeAcDSOj4og53y+Pyz2vETEVSH8bwdqi4
sUTDQJndpWLlcLfSgZhd1QxWc6jZntOf4NAmbBJMZcADrn5z3v3XleCxJUjMMInr
UEtJ4fARJLxbzv18QS5jDPPlcuyaXwqlv4m+e3wIMXakx7KepNRpMpbpQ7fpfYIo
evfU1fRECuwyMXZ1xA8UlsAIPJtSOpzXUV4k1dLDBE6pubPGR8aTT/F54GKRaNG6
i334jfcD02Ca/OPRkjsZsvPWRValdFHXIRcWtYByLk6qIbIydLkEnwJqJVHdv21/
nkCSVG5lzO9VI+fITHeuF5z7bvs0mz6ABrwEJuUJAWB9M2+c6xDJ+Cl0h6otBY70
6/SGpj4hlHmIy3wmlQvyl92+gCbEqz95EgGz7MhiGAsrOmA7CHTLt0OFn2n8JSYb
qGlxvUq62esBIpMO1D/bG3R8Eq3qozW3A7J8dHQTtOwHN4kp0yjB1SbSklD0JKcC
numCMYTlS8JRcx2fOeUWmbUu4XG9q8uSXwEKK1AfsvGqhvSIAQLEKagZp6LrcHNc
eRGuOY4FHA2BJhmOuYYWxeWdjYC7xwBcZ8FbVBZVOZyCha2tNKEULKctVu1m2JRK
ay2rOuQlXK52GxvyPgQtECSfUuZ0FFbpxU1HkTbKj8HJaZMDlksTzd69d0sTyAzE
27zXyLGktVvyxdVlt1Hm0AGizdjpLDwcpgttDB8EVPZxVRBG4vel8DqaE6k2lDnd
TWw7FezGf0qKqAcRnMbcPirzK31yMpQnNAuSr+eXvqfmu/T/JVlvY62l6PAeeAHb
9teDY2dK4ensdzMKpT4VwkBXgTADeggKTXFlgyx9BPf9iiP2E6pM0haEub0A26Sv
0vZCm3+FvssnaWsTQHBVpK1OTOC4UZe8Z2tw5YvkIGBEEozttllhx1GpEhZlcv9X
Jw2b/9seTH3D4Gzkeeut0AIB8afOiFzKSPCsi4AQHzPzxmbaBLUA8kLDlgCnDugM
0C0HBPRPJ1i4Fg1f1TnyeAmfxd29NJowd0uFuysklyhuGIdeZcTJvvkHQ93v1I33
vpCEUnkpGYUPXNVaYx71s9bpOlVAAlJ2lXeHF7O8PQo4HcBRb82X9ciLBNrqLI+E
66HSY6NUy9/+AHR44VeSO3zLWc+m+xQ6skOZOCLg9UAWv2OPlJQdbSHfyGCA8jyW
lC8F7mEFDiE6szBGUHJLbFtnup/gTkYByltV5ZZGhs+9eNaCVB8cy164pJfAH3dV
3ons+ZhopcIVcbKtekkwdSzZdmVDSYFqeAoVBwUE1E6mmAogKHtikoMMHXRZwbU9
fJ59E/7mENCV0ivBhnbXzfGt071FHWVye0bowNknRSzgiV1B5zmrq4H8y1d91wJc
CWzG0dhFCgOh8HKPcUMTJgQCeBWet+j4n9guMba+5i8tTHbAB4xyvr5Obbzwsnvt
512C1rIHzitCGdN4CrCQeg539vaMlpRS2CmVtEzdwQJ4lDhusuy0hnYIc9dHu87a
b1z6sS1K7HF2aG3r9WzeLx+nHl1SM80GpiULOuEL90cVDKa2xgJQiIQJBcl9rDxT
cmPeoee+djh7XBcgly6blpP2GLihBuiuqgFUaUFzddyeErX2eMc9x2PrlaK/70D2
blsDWpuUNm9t+xHdkwpvdHV6f9upTaFnj/qGyK4435qI9NqrtcD1l+6Uyiak4GeJ
no0oX5aCH1tbP2v2X4xO98viyi7gJtikc2ftPl9vnWQ/fj7wXZYMw4nFm61du/lD
n9JXTH03W/Rmfkt+GSVXjDOeOYcdqlrn/Bxj+SBcu7SHp05SHuVFB7xOb4Br3Oqg
z3fBTP7ZW+6LnKZYvusigU5sQk0M+eTnxYBpzohHNCRHy6ds1PCXo/kmqRiDyZNh
T5WGk7p/9lVc0nPcONyQfAfw8cITUHZ9YhRuhTINbGCURsd5nNwi/bIHZX6dwq3X
CQmT8tRE7DTojhHmH3jMuQLUJCpnd1MW4ye1RUF6DlI/D+Nd9NTfSlo+v280l9bh
shPwx8fGxQm2Dqji0krOTbz64XrisEmp7Mh28U9POTyshMCxLwtFMBC5s/2g6Bir
GlDYvgI3K3Y2TT+04XNHdIwMIz5GoVaZ6JvAAapcS7uP/gH4OqTlAA5mba+1i/Gv
/x6G+Imw9FXa3ANjrB5NOvcbBGx3NfUwf6eI2Yz4ftk5/Qf/3s74TqDibnIWz4tp
86rCAy6lTUy32AjwoVVrdqziBqaqgIxwnTA6vuP8MYCWYexeI2RFgFDPiGNHOtsJ
C91exBLRcD7YdUS33AJEBWPqVMDCuwkRMATYcNhoQw+mAOqOuZIXnSALdhvWdWYD
MSE3bZ0g31C6h8+ToidUCtJRc85ojBd9ukIY0gfmBI6oIdg2KyX+Ffms4yZ2Mu/W
bf3y9D9I2pWR7vZXgdcVTPARUAP4JVr/L8uuiCPAa24398W0FwBY+P48vaj+nU2q
sSXsRrJmlaWkIO6Qo8i2b2cVjlb9owqK01gLcxUJ5DLAeUhv35zO7bYEPXC9boAh
SlSB5/kZBnWRU9UJVK68J0MPWnRIBecBW8jXQv7hih8OsiKcbUbleSkRVoFHCEE3
q7Zo9Am0kqXHtFzWm3oQGe6FVN+SAjwqCld3GeNsek61gTLciIxOqFHjP2rImBmx
mTQhE5HKurpXjAanW30UHZHg+SGDj3yOQ3AMktfTDRaK5dv0Ek753r5G27I5472Y
C72HSBvsWOz45mFsjJDzVIQ4osde3vPPD1/IYgIbXd9YpIql0kcwvfEmbuOTh7ix
4ar2jRYc4HwvLzCin5IRAwRBZA0q3mc/5RbvFonk6cmtWcKgRQ/IGXj9SW8ymdO4
SFAJlkzVXHc9BgZ4SLBzKS7U6ExKm7SkLFph8LCamfJwc6mMSKiGEzoA3ecnF9MI
P2ycNNxoDCeIZMyrGGWTPAXmjdpnMphfkZ26s94w415bzQVRvOwRo1wU2OC3UDZy
YdrEqywaVaj9Jiyhbw5AtTCUNxPyRYLYctIhZhR3uopaNqIyNv5YDHb3t7SCXShi
BzPhwQOGoBkY1PRurTDvYDYVgEE8es1BHdzp0JuUkHyZ8u+M+wKrJm6wzDcrC1ga
NPKbjGqmIOibiGBAHOCRZr3Me9cy9tl8IJG+EkMpB7LwsCPMITGKT3WM+wMHcWOd
6rRT9TsvB+IGeafu3bk4pWEvpzmWEWnurVhOIAZ2aoSoGswJKKH/NePiZ/UIFO0d
FIsrttUyUXIFXn0tZXn4p6bZoBX75La/lhmC+L/20kGYf1e4cF/eR9l+0v+i+/UQ
RXtmAuVz/3CmBv0hKNPGnHX77Oz45Vm3Yf1xbhnnFARwPoWGgVoTGdMGwIVBBgsh
8KdXLnsBNkUkzE28mG1g7uiRxP6s4BvxdekMQD5E8ZP0QbtLmFBFAQ0LdSUEkR2Z
xdOxZ8L/wjISw8MEjEFHbFZnCrI/gzsIfw1iKh+ZQXnOsB5m9Q0uUaQ2U21zSTA8
eCt7Nseyvz6PMN8f5AsfwYGuF5Mp80VgrPv30QHJr8GzTzdQPzm/JMkOSBrxHuXP
BFjZNpxnnWLuCkb64cdE3H5WSgwPzZmoajrlJTfkEb35uGcDmsUBeXbGpYZdcvyr
ZKpBei39zrbtNCRiFVmmR5mLsu6U8LG+2Rr7X+4i916yHB5dlwuT7hFSw1us5buq
aRuWHO2DuzEIltiMMBxRlubfpuoBWb6ElawsFXwJ14fE4kpSxu4Q1jTi1/VGoILu
KGFCUxnzIZ9z+ywxUlij+NalKJ8qlBg528ph63VVh8KZ7FK6owF1XjRZx/ulITyp
lpFxY0NqyLjSBt8AvLDVs21uhDvn/rVcY8jAHYIwZiF7hVqN1NLJ39E1YY40/trA
GHYpp5FGKbhY5BkIIk/cUjhwC8bpLraWl0askJfOsQa+TSoYHPZhVIrP4vBB+mzp
39F5G6w5SYU19k9K7BvdB8jH2cREZaCdhsfLsSRBE4wXd33XEDrjrvH/thSl4Ubo
pBZShvlUdC/5g1mh3RqNNS93BUx6QRDT/+F9ykx2qi7Ocs3iJUuP8aLOfTw7Jw5R
ycygYZWc5ebLIO7b7oYXeicG6Hrhle0/IKFciVeFbBMdej53uhfmz+3fJkXftMA6
/3vOl0xC42KHv5ON1fK8kre3/4p/aYAW7guarMC8rdn4BYQxYy9AibWsTsjkhoD/
e8BPpZkbVO7qUeA2P+a9HQy2Dr22tVczInhJ2xPZ4hqHn/NS4ErbI9xHRx1yJIDr
eKWSSFz6vcKM6VBuaezor8QBeUkLjlghwLdiyDggwaMJ0f2Do6Jf63vJNrUug8uq
xs++sSyHny+MiGrdPWR6X3QQCoh7okL3kZmBkIqfEuWmd10CwP2baKsd0ASvwVBB
6bmtdxuPKDwZaOGMOZYsKCznYajVxNll5Iz81Oy59uNwoeUKA+cGjBLZYzFh+QZN
LNuchHYnEHrWfLtkeb0RmaAZ6DgIc67LgGgF2TjSMHF8lMaomBN+uuqOjgaEHX1G
fZ6y/lk3OVYt7AeclSct1HXkAAbhUoS75xPsgzluDKHZqg/pZj66py8WF77VWioI
WE5P1YyveYe275K5VYNmr/0gu8zyThItbS/LGLKTVq2DbsCyUOQpLmQy8H7KbYzw
IfXO3c3OysI58233pxvMVeA4Gufh3oc/f7NooIieY9PdVuJh50iGGWUMh4HLSnbg
eW4MFmlKDzcbRfSaPfPWNBzzjF/0C1mQsKMBX52DQrrZPX2ogRpKtye1YOrK1tvh
15Ma0ubZdWuwiwq8kSgbx/S1luadolI9S14p+oFG0AvQB4p5Cs8qU0pqh3FDF+n/
hIZTJJiNx6LQ2owVoM6MczS1hwIssbjdpVcKysb7fxg0XW1JyaEruXrPtMtZ2AQd
/Le0WApm/NJDPNTLUWZZF04amuayfAnw6OknFJRNx1P9flHocma7BBHuW1xg3+xE
AnCgHRddQW6j3c0FklWcZsh4RWjKY46gP+Gv0rHweis3Zs0v2XkeKW+j+oJ0jzZB
gXRJRbLZsflssk12rR57x6bU5lLNfixBA85Srw5MZiRCqNGk7y1DrQkz57vhyoau
139xnzpNQz4hsN2PkJJswq4j7JVjdxpkYQ3b8wZdHWRO/95Uh1L0k9xHq6fXdP5k
LlHE5irL4mWMD6kQTi+AgoTgkSKm4al0ouo0dEMDmZ/FenRDTdrEtro9VRV8aeWH
/EfDrpRWzhuNQC5lG/cZH4dhJFwaDA9m3DtDY5VR6lhOJGXcg+O0OLF5gsPwx+w6
V8Y6v135atK/SrRm562vE4FpPf9wE9OeGpAZX61qG8mxyZNGQWxZymvhYi13S/ax
OHMmbmU8ijAvED45LwpTRY7FRtY0Bf5sh8EuFDQ0Rz0hhYuuwiCMp+77c960L1Ym
xVd6ErjTLHWViraBzZ88lcCa+P+s4f20XC8VVLAjQctS+9asm3FYpbNQJCm8w3Uu
+X6DlNA8ttX5aEYXtbmZ60kiXX79it3pKBlrv8d/lnzhnu7ywF1zhTtyjgh2J8Sk
Ne38trL1Ap637yrY+0EFsak2dm7ZrfwkFxqS4wzt4/UfP7I6ojT8znfATQFkqJyU
6FpS4S5jty84SLC9vzLKKTfZUu/sZ/u5ShyEJ0nQU4sB07EO0qjt5Faxgic/At7r
M3SIeLOCsqSSAp3guAQa+8G8mI5peedJYZUDojEH1Y3mRb64jbHMzGwl44++aQqm
vH+Ai7GsArjMIph1rIywEG9OPR2TnjsVn6AJlsepCgdQLzqfhzO/DBZw/Y8ol9XL
tNUtkr3GCOLDINRM9jie8+DDb/an2pSDr3Ej//srYLMFFq/qoFUImC7Q2a6uvr/g
qHWeYbUGEr2LTG8ayjIwn9nGkxMZ+qb7cdvcKatXa2amVi6q31tnQFMMFhfNLL+6
3x8qF+oAPs3UzS8nvI9C5U+R6QjV50SGoNV3I5K4gsAHf9UWTwspukvireUNIZUP
Dw9lDOC2+g2S69zQ5N8mLDBd8WvIto7MTwC1mkCn+0pxqt5SZkU1zIQxfe+uMzoA
g/CjJS3PHwkhpO8/Uk2XZlxf3QmjUnsxQ8s8NTw9F7bkHs4CLqO96WPy5F6IWmw6
lUlCYS9uwd3uHeIUcV5n2O40Yn5xbpSSdmkxnBjbL+SrTXpdFa2Z5L5p/cxRufB4
kjpnioPn1kgNgM/iX3I/qDCAxgMhgQcfmo/75izDrWtBiyMULMOkqu8xRQ88nzXo
ZkdA6zrLfRI/KTjMbL1/aWDJzAF906gCj0k2UjAU2bnAHuHq3acohHKU8rDIb5Hg
iGsritbh0JwJcCdgbKAbqaku1XR8ChHUEbwSWEdsTPx/7cwClfyiR0o0nveqcpl5
ZWAYktLJk6LIR96f6n2KKoWH37a6cuf4yKyMxAT2pAENN5mcDlmrpxSUvUgHoFhG
jyAGUO5QsYsblESIuyAMEn8PcK6IR1WuJ+o1whGkHTxK4lEvZyqBEujt7IsVh2RF
olPtEzqxmcarHV8h7I0iurr+7G5307nV3Vs5iQ8giT58CapbtTW7WIwFASlmfYs3
ype3PWJopKP+MtEroiiakzkqxzaTLHmKzcZs6Yj3Djn9p1WLnxUI1AQX7HtPMoM6
CY6ppbvptW+a4Z+bg9aFSvGy4WT61NxSp7aOero+ql8CNPgr93UX4Amneb1xYLGk
l0n9rLpKmK/zT0QAfDmjUBK2XFF9aucPQ+Mi1flWh/wAZKabmc3Jrp90pVUcspSF
xSJSa8QTFAi2e/fOJ55y93jjehizO8KCeaMDmczL/eK6PkgbiM7E3PzaQ6AdsagM
Leto5q8x8wn7ROOLMWh0jdNE5bbfpC+FVFJJ74hiue87uf7fI2Jw9yKF6FZ/XctW
VgALkjt7ZQ01asGkQkezyYhoK3YXMZeoflPR0NDS4pHEGyu22/jW7nkwHxj+ZJRr
9tHB3POpz/AHCHOeCHxT/BT/x0b/9wNSuuxAqCqaBndABzyMa4QTus4arED0ELaT
4ZfEbrQmcgKbtxtWn8DCc57IqdcmWXmR2vVlgNNAXn8okJNep+WzWq3fwuQ5/bv/
FtM7eqP3lz0BHZ0a682KBCiie6YGYays9wHL3j2hQyb8t35PDoA8oq9t8i+jha8T
xrZ5Cm2wEESEsi0Bw/yWoA0hawaJzTRgMbqnEANVSghqwNndDTU+9guJqaGVR7DS
XG1ubXVZvigosDJ0wPxzoI58CN8IjWIGZNirR7MIaGB7RFYU/cVEOPMD0GUbObzV
BJ2QLDGasdVf3SyPBL9mmd7wr1kUQhwNB353gVKnr8iu0fgXtzCtGbFODND1/FRy
v6jV+mkIEvGTJSA9dx3GezneibIAk3ocgIA3vmYgiTmYGI5fWbmN7BIIEFkGjahQ
XIUSpNIyKw12yqhm0ySw/d6GfOOTPljW4lNGxKcqIuGgQFQdI7DK8uCZ8omDLPRf
lycRjomEvG1sh09nWLGhdohhJ0aTfTiSz21Hdz2Ndf22hnslYdpcybj2xiO18jb9
9s5lf9UAq21l62pOmMwoBdJXYFJGLtmSyc0QcZDzYMjSIZMSiz+jsuVWQeD47uoP
fdkhMlmNySpHl7+OJmgGSkMSIvkIidTxfsRetcSoQ5Zr/2RlGV4sEGmeNwfGaelS
kvOADT9iXjVrWgDL9wFyG/p+44MvPXygH725o16IQcqWSdFDwDnu3d/gRx1oCL2q
fw7oR7gPLtxUVRp2D6yp+dTEwmm3OUEDNidLFKJAIZavpMxQSiC/Gqtyc7+q8W/Y
CaxrZT+9+3raWkklcn+AhKxj9cPQnqzxcZ3EAU+ndN/Q0AB310tlFf7H35IHjvfs
Vb9GyORnhLmuKI7tRP57hAP+Hq7mKTLDc8lv+CW2b+LE52fYml5PEnLEd0IUwEPV
3InbffZDqrBR1eLatJNrKQ5RI0+FzoyvThgz2ehebJ6CtG6+84zwE3zxXaDjZF5M
GhDKzUQiPsBy2aV7tqDxIDUYtVcSMO0WlI1hIloVr88IgZoKyBwG6OWXkAiV8Xcl
B2DDy+YujY5ZvsHmBZhSeO3QsLvb35sA15JwXBglwG5yguoZPh93TtF7FUa/kdYR
rVDwrVXqBpiQgzY5l7YP1H+ed08PLqWKVisRSOIyhLN9B91iE/wInWe/ase6JsGm
3HuhpbTTSfHiYz4ofsZzsDCrm/l8hRF8WKnL86/PYfpAp+IGUy5+Dd/hPj5Hoc0K
zlrqvBjtfL4t4Riehw/bVL/b3a1dgeT4/aGrNQllnMThk4SAm5YPMEG6GDrmdL7z
s3ffusVcQL6O+hasi2ij6nvntQK4Rlb9GQ87VNQ6E//Q3/8nXaGKVZajkQdXSX0P
TUEGZBwVQgb0LWiSSVWZrb549rnZw9FSVLJ9P2kGz8z2f5wHtyMtdiIiy5ULL/ME
/k7vNyjLnEGFysCg5tzmumBN4zpcnnwryndNMMgoreF40zEXKT2l0CLklk0AODgU
Bl0+Ny8q0N+PX0crGdHkhPyXW/uWR2b/jUPKNMm7ZpTjwQCHrUHg0fET5SiZPjCH
4VN+hCjY04aOUo9bl2ZM656qU7sN08tpt0lLiWH+3vs2fblVMFRu5hE33JIrS0oQ
rrMfNqfKSjhuZj+ibAtFnxmfySu2GA33Ov8PUH0X25dj/n183E3/Z2VszpVh5kQW
sDpTjdoL7lo2ELg8c5bPZ62IGkUYyCd0bxToSTSQG5CjTGhm+nq8X+Z5vApHP5oy
EHWt19YS/kvETUQzZ1CA19qtRyzyWeMzwiE29n+eycnIw3QvLFw6SchhBZRvPxAS
yPRegfGwjpX3wm/1jV2ZQmrdhLlO/9mf6fXlfsbSCWWgvPOc/j8SN7wU7du9ue5W
jCENb8muDhhnLCkvSJ3WEShBG5JqYPIFIUhdAFMC9puBjMqyFOQpb1Qvw9ks2RkT
Mwc7gxnUmg9ytsuqlVaOk3dTA7R6ViuOa0PJkWvFHD+8d2MztunKrMc2L3cNpH6S
AceQI3CMHf4VjNlINCa+ddRqcOBXKGv+DeXw35t+cHzxQHNdQp5DWHnHwFvi4PvP
m6bVHqmBtRXxCD/Da3kd3VeSSB28Omuu4OvTujAzgQGnOr7RgSFgRhKGsJ2Y6Lhn
NiO3biuFiE19o0NwXh7c4rNd2g+6JUBOqm/W2AMpV8pIlK4xFsiDVbCJ30RhTzpN
+ECzvQ5nmKwI7YPhIoy8hFphJKwKPCUoe6pwrwyvB7i7LAxMU+WMhbwJ9K18OdUW
SQK0a2Gdj14SnUGmVFGMn0eVbYh4cAruwSNij+9SOOjY0B1P++D0h/xy3rjzayqQ
F2JRxXOFhFusvGYfGqjBeP3Xs2KGJy3/MnHddnhf9lDaHxxMRZ27/F4ZTvW4Fool
j1QIZhbuL7H1dkoDVynC65yVBSiwABgj0lM3/JiQdr8dYZGLMcgiIZ8WugCkmohm
kTSo+cEK1YIzq1glIgMCGRMA3RxhwyulUU2W8htInhgIBHBxCeykcrhRcq6BYzYh
wcgXNbF/J+FD/6eJ8N71AR64QoVvb2zcB4OI3Vjr4dfiFuriSOyjCc/Nq6u3qVUA
uk2W/I54KJHXaOhuewtJ8TLYXfYuxtFVE1kGf47pJp7xNWyv46wCugZIylSP+Yy5
sdB+1F+lDYBujUmdxWH4UI7uuJAWeErohpHTd+MpX0c4geaHMJ95t4DBwsCrHfeR
ciDUjErUJC4gjksC3myJb20D2XEpItCyy2vIaGZX7yl9kjFexXmXhDlve9JYrslS
zamSZjtJ+Zc1+3VHDglSJ8dI8B5nZNqrkkvK82sTJlBmieN1VKokKM/VcLue3aP2
RmvXo7zxssM6EVxQ2N4e53DtzjeJREP2u3G0+MLhymlGWEQTb9bv9Rz6ojRqPYId
nAjdgFERmdQZxROPD6Iv+kcCLUVdyE2fYXd3ZsZY69w7KaoVLr25EX40V/MrmDqU
LYVs9fz/diKvJsO0vSLGADgA/3SCFWq0P5YpSacmsL8S4SgCYLnTeh5qS+IImh9J
cBn8Mb+AxFk14FQ5yziozL5nY7YBC0APuTKc8Qh7UO3Zjn5ygvLhZobTthfdVbMq
ojdM9ZDGyScnSxc2gv/Vto2v3PuThA3hcgLD3zcBOszJhv3pemI5scGLIg9rojb8
ymC6/qsN1l5H48mcPIUO8at2iMIw/y6wSgG40TkMkQBZtbsj4vkEX22TGAQqKGP7
TL4ICMyIDzK2u9XyI/AEF3FRDgGViyUfO6yGsN5gGSzCnZMEaWjjo9s3r2erAX4A
EYU306Pr50yzskOrmPexeKl8cWp7uD8wpEqwq58Kznr2Y9T50dd8vHI+zf61wqKr
0Q0IRG5sT0oR+fvbcXqJ/Nh6Ei4b4i76J8j61wfjDxy7RIHkrVRr4QX+iJ60IHBj
tB46S4KcLi3R8rCYIQm21Mhdx47QymUSMUOo+eQq3e9nEoo8H7ymL31sZT9fdb6k
TuiYFrxeteK8l+IpVL2PsCCqTAtNvpzF5XbG7IAxZ7sRPftCqd1xxVp+ztocGCA4
uxos2AgpVDGiGYZkBdqzxMhFiVHXPDhExD+uQFnyNQif72l3P3jYzChN365IgWLd
EPuftZs5+mvKPBrMMQ9JIy0GPnss7m2bZSxTpSe/XOKjZ2TakN9NPudxhfkBjqfS
MExbuTgRyHzdjhZMW1Bto9oRVkj3/CnAd19bDXgA3ER3T4S3nUn3ikFI2q6SC8Yt
lW+XEsduAIwPIucBET4zILaxsw9i2GoJbELOMvKSREnLrpmwRifkd3T/cRkQ/hvV
YaI4nDm5kkTncmTYBr0c5Zq6HNedly3yx1z3Y57FdTS94+y937YJfPtNl3ynj/7x
cupcEf5plYa29u1Ui+L7aESwmPKamNAQmEo8DuKgEk4f6yTHPxrfImrcSWcr/Lly
W3Rr5EOQpwbqM0zPolCgbLU6N60mB8pxHn95IL3r4niC2fnGl3N93wYN4mz3zKyo
F1ZCWnUTmMCWXqudCp1CxLDnwCoppTuSLRAVakl7n17+sE09bSpUxYd556QFMIK2
wtygq/cC4KACIS90pAFm8KZEfGebnPT5kOl3bdCzP/l1dkB7IV3dgg39ZB39nkuW
Pgtzi1C1/JuHFFD2it9cy1uqjo2B++lB/9Pw1C30vw8aLob/AQoZbafXNDHNPxWk
DsdHjLap/1w97vXuNguMjmCbErPzA78/3NaJODTse8tG2RLMxS/yA2Tp/PtgHRw0
JjoQUbBXRQsqVAI862MRT8GV7VGkdsPOzwSBw6VEM7j/9RUOHPYAzv+1afjJ3fJN
tmT7RnVd/tgJE6CFgbCa9XtDT5zb840p7Fxr4OhS4ELTVPmQzlVSgQRrG9VI+RS/
tuWwmr+AMMQpsR2j5YVZxbG6LoNfXwRwS97rmrNcYQw6CM6LLGVzs8qobIzS6OX8
/S95W7WqhixJeVNGdHoUoKqfI6/bhLky540Uymq2pziHPZh+oxLxPEKa2U80UcmT
o3kdm1yZ6vOA/GVdrfh5a6lzRNjQXKhc2yOzABz61cdWYh/GFTWnL3UhzN8C0gjE
85N9yjVTT6T6QpkvDCWpculQvFDBGM6oMWzjB23WyifAETCcsiGO5rzXBXSGFANv
DK6v3JObDNiTGRRLWu0qI7UbHBhrSq2Ca/zgqm86TtlU0EolG1JtvGK7bjgGwnry
AIKRCM76uaqUSIrlpVpo1Sp6uDL9eQ/3iumrI0IRqcvOrUN6HDQBLPAPf8YTv0bY
BowB3w11d1Hbw4iQZPxEkERe+XHBGEnZjqLKEPsXG+JWH5MsbNeOVs0vsnhlasKk
DcU6OIGMYTsXN25RKt3SuICXuCkL1atWY0+JejRHVAStj3JRejFueKpRegu476Hy
hxw90cRCaV8BdTf3ThuK7mZbHXc3IvreHnTIH5Caekzm8Lp2vc9cAuB50yY+CEgZ
7Dxjwlctsfk26gnkyVL5l25K+iUgZ8nCYicHr7XdtQ0HQZHHmLZwj2PTHVPbIf6N
gzLYfPkvGGYpYeo7wW3nIxBxohPXr6y4qj6S3Rr6n95GxM9BSX3iFXyOLLKesQCm
804g61nbWe5yIFGUivaZe4FeHGFu97qvjkHDyd0KSpVBPKmnzXDQLjc4apsbQYMt
H2IcRw1z8bDP+62WcV37ArnCfNWvYFeXhq5iCey3kKrG0i18TcN+Rzrt80d+6doN
5sSah3e5oUsQCTdzEqlPs/ekpwPZCJBpa+0ujJfW2ZEOLlQOW3di18QeJaP2xbub
UC4HpSd9Ut4uk4k+QY9PX1woyzyCqzn5h7SQLctFWYno84TcEl6up1hAV2w1dPjF
o0SFNDnyUZm0IVEAB4aaIbJKxKknZ72nwHdnSLi4VKql5UmMmEWZvMUquw0Ko0HA
aOMok+emwSLhMEyDgrl3SNcZpRhgGscZwwoSIy24REVlNsl6uCS2fu5WuVzrM8Th
V6iLf7qDqDuQF0Fyz61oqjUyk1Gum2gucfj+Xg+eM2ycCpZ3Ukv9noTc7qsuodf2
wg1a/0zeMMQ7H3SiYvgIraNOGr4iZVL+imFPevKEdy8ecXVPj9ZUFoUlCIRrfNjd
FbWkR28GrB9S129HA+yL/ZLAXMsxh8c1+UoZFOPYocyMyYuwinPQVsWFBEvek3SJ
r5k/hqQ52CQDdouvnheGWFwNe5JcRYX8ZRTFwY/eKk7FUTx+pl4cYrnJG7AJJ7H6
c4gZnH8OrjrYEx9712a0ZOcz4pZWvBOdWAgS45Vrhz4oly4iwNpigAkjVvZAi2rE
hyFHJlg8Hsuq3WyQ+Mp7BQcacNSkb+hV9s93pHvdjb/XLKH3T24MsommGPBG+fIo
BZDBSIlktuqsRPa32B7eerrH8KYP5k4wbqcsCRvMnZMZzNZsBZY++AU2dIC2Mj2m
Vwh3uNxbkdmEfAaus/XRiDPugBfB/xeRpBkDtQfopxg8lYfjeupGBdHq7wznPjGd
BT76g7+pJCKdY/ckvFraJL3CAsAoZf9pGFUXNsBS+bJHFw4vj5ezgO/LVDsJ+S0C
HgmKy2jQ2JESEEtBsbJeqIPGt13FV9h7aXhNBdF+GXeNtZNbURqheRQ/2P9aFtq5
/VlGt8tsC+mFG2miw9WFmJbnwEZlUvrpqM7lw0ticLQUWuGetWNtlQKmiOwkpNXN
9s5PQJlOCtkBsfTRjO+gcKJFeY1INkDVdqE30MZpQCnzSneA5DclGONmQJyiQbqx
WJLHIbyIqUBIcj8fMDCDSR2q7ZG7/taoEdwzQKhT1A14Tl9ylVb73z4AYWPI2gKP
MM1Ao9w5dMnpKGnqg9NqRkOvm6uViHDUJ2V1Ql4EWTahnS170C8P+Q5ZVOnD8dz3
xk+SOl3Ua4bdnptFYNwr7sj7C4/UqH63aAEB5hcpjm0O1Jjo9LXWT/XpauZuRi6Q
U1htwGJ2AzM1NID5RLL7gTcSFW5qM7J1SPYbR3YXrbLfq3OwLsRd9lLOhR3ZSyDZ
XdIMqDWYs8QnERgrHQLs10Jy9iVAcsHO9LFwQh1tFtUzhVfeDEWvcyNw6rfw9FkD
kVQH+QCkt9TO5FZqTMMQmaBH2pwb9AcWMmlGcaCsdaw/2s9HqVvQTJSf/OGhPmeq
ux35dJPXD/N71YGkcSG9YNwVW8x4tqFxEmwL3lO+lMU4D7xhkgW+zy135VWASR6g
A3/VDgYCrpPzcSxfKAIjodTpQdvzAeZ5cDsfxkP/iJr4RrRhK02K3Gl3tTbpg6QZ
4wkFkQRoyk6lrwANguGEwEXhv3ZU0Iq5ZmspumXUtwMQO8Hm+qGqUvZWqgmb/o5N
WSLAv7CF9j4WeMNVFmVeS7k1lHFwpMdfmrHn4jxsW7HuooUuE5h3uCx3z3qgMg7R
7/wyBfbNxkHah2Gi/BY2Q6S7BsJ7UcuxlLlNGNeN/A8pm+EPoZJsg0ZVLtTmbORI
QHfAK2SkuqY60fAOIRYiwXrGFpoPynfXLGM5GlSWIe6m3zAtDNZwtidU37VhbQNP
jh00/pKJOePZfEtxUNjZU0QawTzdOF6UBL4RGeBlJPyBxLVPrOV/jADIVc3meCRS
RH6jsbfmvPHq0hPVlvB8BhOSn5yp2YEC1h6XY7Ha6s8sGggvLHdtC5ERku9KmA2n
2LI+m3Rlod1SEodubTE1dLnmG1nairWKln8GBAe69rWhlNx3PqvAOpaaovLGZXbl
tPtPyWaLiMcJtSDBgu3FSzhddC1nfpXIrl9Ku4pBenbaJJj7aUHwwebnc2CIUkHj
W/LtGm7wk2R9w7Xhz9eJw2h0rxiQ2LBQm3NUntKSiqlbat7a9IZjMch15rj4pn54
0CDupT2kEs09jKOkCSqHPvCxyeG2rqWi8E4meXKslZn1GvK5QlD/XhZOwwxP2I/M
drBpG2GzI9nLcltXyt/+sp7rMV++quQTMsPMnWCVD7XjpoY1gCWnzdcGKqCkxJf1
lfgmP+Lod/z2Iv/oqTPVAIT90r/RJeat45szJdPbZRxQPzVQkIRFM3ZPn5+5Y65d
ouHaHHbWU+GSAdH5uOM2j9cBYoQPJxnibBbKGKnqxwwlZN/ibZXdvwpQtLy/rJQ3
FTk1y1D9hMxONFuHLghpKWoB3hPWqu179xSH51IW1hjZE4G1dMFJx1cTUhi6H0Se
0PybZoCMfwbshRPiprKGEQDRrLfA8aKx40YJIsbihClWI5XWm02A78TQ3POScJ1v
/cRPk2dVq8Njz2bHssqGqNFUel2kGtnq2AGCp5QGM+Wlh1NzCAaO8eeaS1jf7+Sc
dVksgzFaRfss3GCRMnn+TNp/kQudosZGDop3ES8Idr6t/xewhaQJFJruWflac2Wy
hx96csjw2nKGRAdhkTDcm/JyGh9Ihubxa3KKgrZ82R6ShMuArWViAt2Plzj2giyS
wnvk4aM+vm+CZ2DddN3hrf7jKq+0myQ2El/cqrgJYRJxAihOqhORDt9v8STb393+
E+AHWYsvTr1KqbOmcUUBquIgUuhg6ljKGH1rcAB5UlTxafS0PXAw2PjT96hfyjcb
IRNZQTVAYg/2Hw2BDztfRnYPzUl+Bs+9sIBAE0D621zInQxoZnLd2Uf8BvP21BsN
3lUISaC1HwOuHzNeVdF9B+BVIIpGcjEOEWLFjoOGRR92vljj0NJRNcI2QpOHa4oI
hly19KjfcG2uMgQY4jkjr6bj96XxPYIkODgQ61UaFA5Sf9Zn7hkSfUSsJr7I69np
OnMgFLD5h8q3QgBkZo//ygHPGOH6EMjmxhFlB1OM3X5xXVmTSyTFJWVAmA/abDHZ
AF+tHTv3JEPA3mlOCaNOS/PtRUgin3shpxuUsikqRfzlzsL7oquoZlUTbHdXCQY4
7bdnwDZ2JF+8nmjiyJiv2vrn7BPuwZgtRcbDklCPY2Gm4HH8gy8od4ZKPS23dvDl
XWX8x8eZEJXhfAgAUolOmwI0LvJW323g5RMnAqB9gdhW2BAxNSl0EMwnwtYZRner
9U3NucTemUwl2WSORCwOFxkIDxQwfEV/f5iDhzUlMmkKkMGk1hmmfRiAnUNOWQH5
fKy3zc/yVjUp+gjyRM+MF7iUphKofaOwOYW5HeeHdZygpI//SQSn9J63g1yNJT2l
/Cp7KMQ9Na7huTIX3VTQfO/+R2TpYDi4LMoVTpYXm+B4TlMqkV2D24XA7eHnwSlI
o7QqatF8q71A12E35POUH5Fr/l9puDvdx/VxGH1sQymyfNrFe3RJ1/G5yb2zRjKx
eb1ffKzzdyWlMKeHYWpibASFHbT95f1t46BRj+0bOpRFzfnihnMo2D5jGldBKfDY
a3qT2STssOl/8ITMHZtEuQwLuxJFTqqCBiRsbI0gYqoUqgaIfgZHYxYNussxHi1d
pf33BPsKhg06GoRiVTVe3x40HxTHvA6hQrISChD40yn61rVnS+aCynpCo9f0yuFJ
gHtCU//3sdX8eFNRKgzhE0X6WkEd3fkdpE6cY/vbL6Z/4H7bBBYI5jNu9ggppQTG
wI0WXteh0ZD6aYJEXFb72OEsGU/2yWCveC2gh6lohqKDV4TXjRwhxI/Rwjw8EmJ8
0IFyz1yaoBC6j3RHn0Y08csVZ2WxWgsSYwlXjxuitthWTXe0C8TscnUxXdWsQeWI
ry0d/jGDB+6zHMRRt2Gv8OY8n6ro3NF1UA1+zavxPnMzqNmJSO7VaDR0u0EjFQF0
Z29BpnjMNFLECrz/+3Z+cUZCMao/5MEWHz3q+eCF4L49hoe9B+HsohFPXEJtdHo7
EPw/EiWObqHme8Ov/kgO9tn9em8lNRtF64SwXL4M3Pm+zkAzpdmAZVvYto/LUgih
OVRiy0Qg0tGnMPeCX8x3/W4tCxxxEbNUtygL8v5x0EsBPlofbVqthQ1cNFl3fuct
zAzw4Ojup4oQPpOB2BzU7mIZfMqHSi/e0J+pnGJBwXmkNg90bDZPX0FdoueyxSTo
4qWJ19/RWkyStPDSBWv5otRuRWNoFGOB8BaRchxZu097Ru25WbBCNAGJsPWstd/l
k6tzqgUBDWWl/wEq4hmmItr7XvLXgkB94QV+c9NHodl1DgEiUqKMiG8hfYa2ul4b
bfgdROKswZ/uln+uTd/vMoByRdsJY1F9rwXYwpfd08ucAsavFGC080YjUtiC0ic8
KEhf4Tbp80Uuam3vg07C8mClFCh0Lm1Sp75vYV+3ZQmnCIUKNCt7RBlD/Rnfaz+N
iiYfvZXIAALMi9NMACi7MRttRBltUJHg69WgJ4xHEIiBKfryhLINVbuaBJqdWPOZ
Kxrs3vXj1kAZgc6UHsInyGocFtPMoeHRWExSKEy2E6HFMcsRrFFqHsxuXSHIzn7O
LDxKJuslVq2gohM9bLvqTCjr+hz9+/lGsVgEkeb3Vbt7DFjQWmNKRdtASylfHBf7
NpDNL8v/8XsvQ4BsJvpUaeTcsv+mSPTNTIFoVTszbnsRfZnXCB5ZH4L7iGQ2xA3j
BRAscHQKmUZTdjejtUbe5lpmSa65KL5VeYlD5uBOuVL/cltoQbW92g1kEwYfJOfm
Cvkf9h5xMASoTccUf/7lMlBYusmxB6jKuTpAEpZBe6kG8mGvi1Z5Nl9CkDlxG/4y
jjMyhOqSXohTtIepwmBJryJwqUsH98ZBKg+16F01fiuVr3SgnMGyv5Z91l2wMvtJ
nJxDBAtp5Ku12KemL4fGtGheHLdKf+h2RHY+w2ikNLre4ForQT2AHxDRvGJKYpkd
4Pmf/kBwP1BWwe7F2Qc422zCWh+m3zJ1aSBPgUH3WSr6T8GK104r+bg/3Z+UgoR9
wh26/ojlotoa/7iHUsZwNgbB8bV089J7AWqv9qDmcajmC7/Iqi4m+tPJa61ZIijY
3uplAX7vKToIUfni61qbWjoJUduDFc8yfU84sMBmJ4cf1ODRFFXzewEeETsAhXgj
a9lmujVpTzvPegLW1CTGhdw4ilGVg6mtKrHX1FTsWNUMYCA8yeAINw74w/YEk28J
vvCtOd6V1Y9LBlREysj+IzVvWoCo+NJe/lFIXM1UKrzqNUaInYRu2YEpc2Mj3I7H
E4mKPl8YGnKX3yxNzEhYYcmRWa6mTufq29a5I020hbV7TTctYALkJ0YPoHjUgyeU
0vtvBKcz3HRozn/xH8VM33Bwgy6IH6LzrCDA2rm59Zt3sEFuDpcjIFQA4U2PpIs0
D8O9eN/jKNXxWxe1UbD3EAQGLozqBaOPSAZlwWYDgFxZbknasDvnLe6v7JDyIoJp
iS8vStKytt8laafZZsMgXZQQojOhzMpjhhGIgSSTvPi0sXhSLlMC9YwnraS+Qcy+
DfgZoC2iC0raFukiyeZ+kshcTJkC9YbhwYG3gMOf91JzVkDvnaALFpxNPHj8aVBp
U5NmMzJBFRyrn3STmCiRWnHaTdX4w2avg5ZUaaEDIWkQuohmCAX/AyoMXlNzzWKs
lPemy/kNqs7bB0nJDIzL+Y6n51v/WKjPcy5SmfHVx+pOxrdePZbreRimG4bd3vXe
Qrt/uQSyMqdo9uqPvFMTEt+WfKd6UXKKonC5WddCUd8F7O/pWMToATXbzzNlbcYz
XtiCFE0IW6Ow/Si2DMS3+xlnF4UOEdZ6aNoDCDEONwZ9kcgiO4V/BJaE8fAVgXpV
QpFgjjcfPTTYA+P/m02NRkh7UvKYU/Xk2ukv4/S5c65qXbR50Cxushe6sQCIDt14
Kd24haDqDCMe/LXnPraTDG1B85kAiHC0eSjYP6cCxA6xcRMyfXaXG6AJg5QOyYp/
UuKXC6dcR1gRp7kBJkS7fjEL8QG8buF4+iX0aZ2TeEC2vw+YmJOIe2d9XAyMPN2Q
PG7++SDQZVbbwr3PqYzX5DU1Xn8y9ELzkvfZGHKaSDTsuH8CbjZVYi2VGYynz7Dh
bqVyZf5QVbXzx+Zv3fmfHG/K4SuvV9LOywQMLXunxhs04oyiWK87VxhKmXHpDw6X
/In4MHGyJxx9NXBxgIEtD6jXYIWHPS8ZEZJ2vA/usUBN+8b0rFGkiMHIu4hIT2oq
zMvfczr1BQsvEdVoq5uiZ2adBuXOQrPa5QyuF6gWhVzwTfCYqXyGa6VNCzReIalS
mI+W4vGgSsyoKEY+a/iMDWWR1glFz85r6AmYKqDeGCAz8VYznxBu7ANnd+WR0TYK
k4kwlImVYNEDAIXDr3e6wML6nirpsOgHuozlvGEzG7lvofofaecL8I+LRhggbwpQ
VPEptMaydggUx/5mvbrXhz9FQKDl1P/pGu+V/utAesoZSSbpa2XVGuyybMFLVSY+
hCl+4TC6zkccbYPCojTt/KXaWY+h+YZHXXi29gJ6ltbTlUF/U50joAO9Rv/mhB8U
RUMctFKXHXgAhRAYYcUSdM1U5cfCfVqfU4jXvw5D1mpASwr5bPAewG5Ktr7R4DPu
lCo512kEbbEQtRROqgyIf9fLwcfN8q9/CO1S5lUxkgJKAskHBqujSjD8vANtgtiy
LeRRahNSCEOej4+Eo1QpGNwmS/Bp5J0Bi/hBpAbHYyHxrx35EnKJXqAVqN494xG8
RfG3RPsxrvpjs36e8orvb87yjyl2TjVw8xLOGFs2YSrqwxoPQOJX4pDVcVL3ud3H
eu2UovEiSDZAoZtWTUD+yGDRTWnV76xwOb9ZranNPI3AV9INAhJfj1gYXwQ3Mpzo
PVXAeIwdxS4RvALh6oYxppGuR10lvuw1iqVbbqqJMwHbjCw33LlyLCTBuRl08RMp
mNJ74cOjOdBOaPPkWZ4skSb7Ty2HmJcCfxdwXoAhc+ZFVvf38rvgL+7owJM9Unhv
Ib3SBmPfmC6tOyhqqEuEgID6yqwzyFAb5cgFjzQvbfhP4TLNKx+yGtDfa0+zWMm4
ElYs4AV+ppxGoWE4hbu3CV11NjtZ5SDg0OtVCw6ewXTM3rD8uDIauobWwna+vyPX
byE2/vEgz/fjhtTpMsDUxvnjr17EYGFVx3czBXw2YR4fB6G0f2kU/T0kRzROBVak
aKf0sLYQn2QPl9qE/KbD2Bz1kXFHoVnybV1XNdr7mP5DBGK6nLu+0o/M3sKOb/YF
VZFpEIbYqCHJihbuNGFC7O/Kq3njl7fDr3tgrE8s4VOeS7aBPHd4+I206y023mhS
WqIhic9Hq2kR2mD8OqvOuzqIBUxD/7IbSkxMagNw3uzL7qOjI/a4RPCtg8mXnUJB
MOmNn4lWMw5BuizuWAEb6b01Wze5EhR45qr8lpJvGmIPHYuEtqRPYsV+yUjr+sTg
j9QgX6Iz5migP+7lrbt98J0j9/pFO+9X1OlBTHBXy6b75YHCH2lTJ8CzsRpCXp3C
hRZozOB4pCsnWoSry+pW+jsS6Ro2on8De0knYmwJtDGpX8GB+WYReD2x00Q+zWji
XrOSFcNCt1wBoeiXIKPzsKDDLULdbm6uF8rjZEoNsWUOlOnk6oOxfoCGPlnqpVe8
5wPg4ZEsCpGEi+DEIleC8Jm8IvoFOT+RywdAHoT6PUdb1R6WNpJUlzO0qKLahbE6
hix6qjs2VQ8suSRvqwqkX+L7wnW7u7ckgxlvrTKRmX3rv58EW2dy9UqLzwHUdZd/
Q3KxpDwst++jttR5bYcWkXGsC5BKixy0CwWiHo0JKwh5JrggrslkqqC6RbuIfxNy
9bIjAG3G8IU0qd7n0sA/q0tKaZKaPkN7f1Yugja5t2bO8FeRtpNlYKTK0soPilVb
X0IdUSeqO+KjScSGgba3o7o05Nax6mSP4D20VdZYHNu+Ya+LQ0pQwgE6A6qr5Zrr
93SJsKQLY/92gFBj49BnNdn430b1TOGH1hcoZZIGf8+ud9MFpcpqfgHrTAwuNOew
CmMJs4cO0l1k0C1ohoqPmTUVtXiXFxZORCaA1Ubjw6TJfFIQxkScxT6B3IpfwT3E
pKjXpuzxEGSh1iUqM3qySTwQ4/fN0f+wjQyjHzU1RtR3QYeAhCj0qHUfridUAM1+
p/2i5b6bChd7Tfie8WtgN9/HinfC/3E5gV7heE3jzhWoW4NSx8zNUPI619dZAFF0
S0wpgh9xBw9pyOoHFU5BttU+eufOuHgYxz5+oiwwiUiShHrNcqSue+94HG0fWL7Y
XryjUOx5/A6O0HMhRN+h1H1HPVTyLnzKYzoyV8ZFiC8E8PWpRKGmhd0+QjVlcS86
UDb3pdakN7i4lvoRg2wvxtHQ6cEuWFMtznwbrBkKHxmb8RKzp3HX67yqMZQk6+Hi
E6DJRxsucC3H5E57JPXsKg5C7ipDHiCIQvvqGUNVbB7j4muxG87lzw0JtFdgRbgg
JTSN+L2NCxK0e+1lFLQyP9vLzjRGBYPT2h4/kA2dE11EdCOwK2yUf8E3rcId22lD
pyapSZlTU9cHQdfzlVdLU1Gyy60RKMF+xv+5eZoG12t9rAkfGiZsNhySPy+NDkXx
uPO8of8JJ57j7bst6CcW70ReePb3u752a8cyblQFjCs0sXm2npQr+LvI6dAf3B7X
AyK7BiABSmBXqQvzJXEdIj3qtdqjF3gojxf9+0pjUHmZNGZNZVkDyZ3r9r7snwue
LldFPsUqKriUAQM2vsxv9CA4jS4bAN6KyqpMyXh440cHgz0wJp+eTvKem46yF0br
Gf6rvtKeM2RWwNbEQ4eTB69YAnCB42O9lq+H/jsDs64GFETfAmOBWrebogOdZjDm
d5PP6gktAC5y7LVmcde5hHh5Lvh3DQ7VDn6oC9AyYbZQwsvMhA2ZTQYMNczxjib4
8a8XsAW1brDp6In08tjRGrDKprp2w5A7EIuFIlTciX/bIUsf2FQ20FFTvCdemZ85
1AqgTqHL1E5+gaIJNqdHynZnM0ez5DetiKn+uBUiS8JfjjAfMvpBIwEnuvpMHBAF
ga2gtagSGjhUJ0a4yDH/DXZuJ3TgguwbTzPTUjCPo3fZFCALckeVBGHJb1AoPeTT
6Tj5gvhgUsmFU13lIjiNLIovf3MEJwon9sP9AZVIbyD2Xjg6LKLvFelHv9riChuc
FbI3mspTDdsMb7J6S49krgzzQlgQ0XShtigTDsQ/rnOqcrjq6mKMYa56o2n8NYuq
qvMWuZkBe9ShA7x/ZzlaI+V+ACl1KL4KLKhosIxiAGZPggpLKA8+vNcd1P0bgihC
JLb4K4rUqgjZGqY8ClOSBNif05LxXhZRw/LnPMPHKNKCtor5/ij8h9hlk/VTaNoz
1YTkAkwYKYIrNOSJX2cqex98MPtlywEh7Wi0ii64kIhKIontvL7UdJZ6vDKMZYRo
s1FgxcslHR7u4yVEbtiH2du7GHj3y0W6LtprNaOy0iUZv83s7IBtTn9/YlS/wLek
0JGkvBFxxNvhdpIRe4sQ4x+ao8gb/7nCsMr3E8wUHKpdghbESmB4Q7j5xxSRHUta
2PsH7ROgW9nfenj7ouZAwJETQlVXiwshvb+fd0RazyErWNePA8mFWe/5doZSfWQh
DygHIkIKv7R4t0VKhw81M7JLeL1jcOhOpjpVyMkDi+A8DPLm04gOWDpJsHLKtsfF
0wlJbn7oVtJIogBkhB2fSrppf5bDkgfuIcO1Xtr3wb7K9lqDVIye5VO3S36iwkHk
cduq4+rZEW1yU+Udjv8KT12DAamvRXgq9ovEWNtsXLRxAgybHJHyw39w6qc3i7Ld
h1O/l57sLno/XXYeccY85ui6hMaGn5Lzv8dp9l/ObqQT+CP4x7dGyNZE4oXkPUxt
F7cuu2f24uNj0SWd9Y1viWAj0g9a9Jc9OkCCy+NmHnGoyjy/YOtvTdbE8cSD2wtg
saW7U/kKUnaSDp6PMNi32mvCdUWhUAJXENFDpY1PI9RM6GPfPJYVqf8wP+DtUnxS
OIP6p/AbtoSOuVVvhIOVW9/2o6U+8hebkt0pkXjJ1L29VwUpAz4wPyB/tKaFjMwP
5NP2oMYt3e8td3+tGSCFkkGrVeo0b4HQ5JjHZCYhtwkPoPhKgPF3hbfiepGbEaPO
SqEZpXCKSp6vdaD2EQiCwxIfbTORdvhSsQr5zzM4B+kdCtKHkFc3V5vn1Gz6R/39
9dbh3CUsuljNFNzTy66LeU5hx4P/2dYO/P8SsDwVgF6FfTKX/05RF7L2zJQLu88A
BoEGzOtt0NYJ6R+8VPsqkCwBizorhOzl/62OSaVZh9FHvL2o3YK4ls19QZ/Lt8dH
JFHrZiLtLlrYBVoHiIUdHqFUUUT9dTFOT+GED3CBcwpPV43YMXlwcZDSPhVwln8/
xa4tfZfbUVqhGGQQ2MynmlV++mjqG6wSztyDPE4kb5WuJKS4IImbZlMenHHt3Ffv
pig1Way0qJ9btnFUsBZ402CCsJ7OXs/6p+xbp0SoWPwQoiHZxn27ZejLuVxIwRoH
XOu1Kps9Nydy1vK0oei6nnqxoaq32R3WMuWHS5xGfRQrvLIEmtx3+JraV2Jr7m8M
vBAIizByAJC7+1xek531ROXAUke/DC4nIbKaUIIjZsZG+iO9TjOj/6sl/002u1zC
VqtIxnd4nXM993xe+2KpSCqAO3GRJacH/v3R/beLw5k7B5XhUsoaQxCMM7biTe5K
7bgp91SSfeVg43s9CDHnSPM2VPHu37KhKPEzloZXigpKla1+7cZtEkxu2Yv1r7Za
lzkwHqAnWHf6gvK9O7noGeGclI9x7DH7b8vpD9Kn4yPV1En9orRqxDq0FiaBhd5i
B3/uJ01bNtvdTfB+5UTDXF7/O9YSmwmP71qINCP1P18h2+xSAn66VV1wDSnVQVlf
FtdfM5C0diXsV6RzYT0VwFeYZv2Xl5sm8cUO2zjNcU+SbN48p81jtY6NuQCj4EdC
uaW5QF0fLg2iZ8ffKeGrjZ2ELizyviC8NShRgUkOtZRM6j4w6HE0BdKvKP66dNJi
kP+GOlTJFHaeYnq9DQQUPKs1YPtlEJPL7TkfO8kSIY2vQXQTchtlFKM9oBaEtpN5
QoFrFsaWfw4HizG9QZ3+DgAzZXdhxGnXcYKonwcrX2ZUFsBmdvdWcWrQ2XZ6u4Rs
L5KCsjPGnCdnkDVfdrdIOlKLVCxFkCYoqjyzEFO4Amq474DuNx0qsrvxJTOefrNK
KqwdY9jna079x47HLjj6i8aKP/N10F+/WzjP/UXIl27ibwMPBBO9vM8rYU3SLJs5
JYwaOTXFhNCtTPGhqqKdW5hhneLtra4KN/uelygaM3D8UD/QO17TfhV3NInLZY3I
h7U21ZT55td9YWtQ8X56Mk6zvlqm9Pp0tUHNc8Uqx9arLOWZhL7WbLefN7T0KHxv
4ooE3BSFDtHil9t7LoQJN8L+RaMmDhkNOmV3p8nmbaQF58zVWciRy6ZMFTODqO3J
p5I8cNVKRqxXKBFJhlww30ZaTdR5FgZf+pvhOr3c2TVWpThPdl9iY0+QTN7I2RS1
aAxri/OuK8gu8+iefAbqJhH43iMYSunQHn6Ep+T2UzM1rMpgvk44wbnaM/42j0ur
aTPixVjsv+bU6Ll/0Kt0+OYSowUcix5R67sPI1ws1DZibDaxN0HzkBLjPEkXYN7n
9QznBLdnD7s7JrMHuRQJWhXkCPVHYb37OzmJmEJJh1TlXkLL28LsRMouq9JMrvwz
eDDxg7oAI2rXh+Ip7zF9mTYQazMw4U45+93u2qWNGD7OTTFo5leHdbeC/QlRIREu
8jNtwc/pPIDJeWhlyRpPRGPlF31UoE9Pq0YXZzJm7691ODQ8rBzXNAEVqzk0z96v
cNSvwMFzOy1E/DVlXd/WjHMKQLWjwbjry0N/DQzbWuwUIz8xaZhpG+aoMnnUKZS0
6W8oEo0ORkzT0NrlMxczSWjCo72RVE1Epi8uDZuP6ufVU4mjO3mPHWsvBI+Pa0gb
UmlDneDuKnmBYscz4nvGIuc7FB5MtUooJmvpQV6aSr1Kn77HC/QLbELpq+upPsap
dmRBzkSPbqlMyLlt/8TlPEHgvgC+AWfcWajlDWhO9Hl9KjEYGKXwTfjR2YPKt6gs
LbGTdkzVmMi2bctLYgv0dQhx6P6M4oUmNQN3MFq53T6DWEuXsWPSyRrV1fCPIPbi
zWZTpvT6gjr1+rm6BGyFj0hU8CFnVULvm3TokhXl3nrYgff+WtjKCzPqShspPVqz
Rx69faBZuoyR1apuz7HoCiX4R7lPrwBietdAK4e6+9PMMUxJFxAguv/I1MqnIvYE
Bg14hoVW+eFkmGoHz4j8tUHF98m7VAV8Y52kLZbv273Stplb+i6n1Lqijcj0m7Fi
xkUW+KTbA9PW+T9CBVexjxPhRLCKdkM9W2vmdth4rJnyOTMiBui5mflDN8/QE7Yw
FBQAYiQEsLzZFcLdkJ7KL6OshwCRt5YKW8T7yNkEnQPsngzADQp80IdHDXeMlxd2
aftZQBLpi/ccOBfpEPOEkLcw7KAO5zIZEEEs2NUTBqZ7sB4rIWfQaH5OodojgfpN
tSAOvcNCtAfJIkFHC3GZT+WlraoV0FqGZDjz79JzuTRHOwp1Nz9O7KD0mGNgxD11
ZJVEyTXr8P0zhRDBD1jhLyITdFriawh+45XButJnN0l5A8b/6f4kBiWoSABWvSQT
T3cNMg2zU6U5pkcDLgyMQ8Ibm82fPgJVq1WhW77dV116AmUvR36wqqU+czi38TnU
wCSbO68pozdVAo/77RIBx83iUBEeT8W66dNHA0yGSPAdr/EDVX23mj41oB2duVJu
ylzmjeaFdpzA+UEuBdvQ+0CL/paGdtoaiX7cgimerk+eZ/WaadZ3UbZi3jaIvCy/
Q4Qn8FP/RUBdEvoUxh5OqqZ9QGRB/IgmXdRn2N/ObQxQU8+zJzxHQtxwy9OsRl3N
XNFHz4NgyfjjC5I/gpQ8KJNyY1KmH3/xKx/JMrJpjhzORcffbnVIWCHH5SSGRRiW
xf/+FZy9MTjInbbtpqmE1eHHMVBVx8M37uSw5zhK1m4+ulIDeo/zNMExe5mubwiq
GXFLxO66Ne9oOdjMJiI6E9oWhKsKJ4cdY2F/IS32hENXADRnYzxXenlX/rosFTS9
odawZNv/CCAuntrPqDB+ZrZb6pGTNgAK/88YJN6KICJieDkeo0QRgOW2ymty4ZRh
KHR1nb+/MjeN04j0DNsiOJ2DH9HgSB1FZxbZybQh6QZQDsT3LJr6UvYZCH8ZfLcJ
K4p9+AViRlu1x8ghmBBuiAXjVRJmzFyUrO6L1hQWyWEoSpZbnVVAl20kV6fK0ElR
/xTzSEf8tCtJnAR3wKftX2aExArXmfWS13SzQiTyWGVP8T6D2wsvMs0rS8UT2uJS
BT5//VAioGhKTkdjY0b8Fyl5usGLZD6h2N9NJ431eoRDywAJtaekw7C9RmcUK+KT
+gMPN9b8/qMCxwHGvBvMD0fl1Ghog3nHBVFHnkBifwUwSAi4jxEiqCFfxJE+0VFj
qBX9EQ1B43tefvt7BX1PWWaVaoAhe9sZ8/OlR/oob8d2+PP99Hz8RReD2HZiYtbW
3aEap5r1N+Jzxx1KR9qAPPm1RmHHgnLusW6BC3PUEEaTcDt5PqBtNNp3qx+3Iqnq
VaMHE6908tDhpoP2Q5dFS0MHLmTDQvGHnG4Kfi2T3jYM1xlyJLFt+CA//RQd3+ej
hTDqmbSPr8wONTSsuwT44DMs4DEoRGmZh7CJaOciMJNPFzFl4J+Q5m6vmrr7M0Mb
eL54M1Gj2eA6qcwQ2pV+LgZoTZ1M5rwaGmMzt3dah5sqoX5E90W3lJEzut1MJua4
O2+bMPmhtACj1atPLTCnRiA7Pn50YRUcQ7OiZyH2cEMjswGmZaYFSwZpdbIZWt01
oFpADlT/NYK+LR/NqkQdZ10YLqyer1Q765AoAeOea4njkYIZFr3+1KDf11rB+z9C
RB4A+WRikSjrXP8ksTVP1SUrg7HWm2INcEKV2xRzCS+x+R8dXUZBvNQW54Dhygkw
UpVZq7KVHb2EdWXBfoyUbiGmfgg+lo4TCZcIK2CNF2cAy/MzSP3/JcET6rqk9rBs
Itd6RgX4aYVtP3qyz2SPF1YCOZr6OUpD/+rFzwld3bj+9/AdU9wJEhhc/jCXxyxE
l1sY5LM+ngdXoQOW8eLlED6S+sA7/BWyB3/cD138NPs2UFhV+uky/f8Qh+BnhOPR
DIEBerVsangZISwK+7u7jRHqOzI+RWwdzf25pb9kcsD6cw5fvsay9mOtjIZl4VxA
2wOoyoYdnFzu1ONdG5F5kOAFvu9lKdlh5j7wZzU2Vz6U9/66BUhsZ1dTnl5davcG
Ln+4trRNtYDhxkhraVC6UrQwxIzh7bos6iDIBj/gtOjvVbYHX7gnwyQjSRJ/uh5i
3Jk6ByhiDL4lANhSN74pfXuV+0gZDmJM05fB+9LpKTd1AZzdEYX18oEomK7pc2lt
tdv20FQgvMFeusZycYHo852TvRaeDRwUBthY99wfdhSaEoNu984hh79tqicxeO7P
Ywj681FKPJVA1bF/SouKBM+zdqKN1+wDupcJJzYwY6dWDJ9hBXTo4BgJMFpXJ7rr
dQrfxMLyobMs3KwaJqFuBiugoSByAeQxHhYHQqDkHsB+GdIneFrimvW1oUt0ibfH
+CW77reFP5ApLqUblKWnelAym83iEqOcq7Npoz9n/vuJyU0yTxOjy5+xnjIM4YrQ
8lpyXdAYZp4Q+bUOugsbiBWFUk27AI/nxHeKB0Ldy6qF3o+E2ixF9t59LbJbxAA4
OTTR7H8YTiUmLxIWjl5w7NwsdoKmx68AEjmXa2ooApVme00uEM/zLz5pzh+tTqn7
mL3XxxMEDctnsUTJXhZK0Qd5PZQO3HXEMbNrtJ5vuCeidg0SQzUJE8RGoSgT4Ky0
1dCC+XVHHlbxbtig6nmAknA0hAr+zIcpIT2d9BU53pGedEAr2xF+EfegQlnJQxuk
Io2hV+e4ALBUgo8QKwCp6EUpF+YnmeVxSb6JmqqBMJvKnCkZEC8yArkRyOSxKbXB
qtQzWWdPWAAstlGZ04YUBgmH45sKLVFZq7P8NqxUlR3T9PvO8/LULrSFwkr8Jvpe
8ZZNweyabhl8SSp/122KyviZR6rXHuN3W9gGRD1crwFC5QwhSfoVl10Ok7BsJqhw
X4TGpmU+/u539ZoKkZhs4Yu36VqkYJhR4HB5c6/KJi4bRfpPxkTIS207E52eUTBu
yQbxTOOChCa8lxjRxdhcMVe65EvYhEQKi8B9cjZrKzJ3sfByBNdwf3/5RzB1VicZ
CxahHfsTmC1gtn4HYRccAvwfJBnfLWlwei4Q/fA++1lSIByvdRkm5ltp/qCXavFT
0diD85L8HAK93Pyg2cTm2G0yg6x5GrLr5yEYFGO6ykYmjmn+KoeV2Bdlfbwspz/Y
23O+Y4D487tY3nCWXtDRvF3SgCXDWFYMFcMVzW8CxLEzzGKrvqbxJJIPLW0nUDks
x8jS2gEhPfZpZx4CrGyEbS04/drEjGHMR6guGDvngNFvR8spxTaSIgBq6x1aXDvt
WeIgNjU5+ycj9MfkUgVRDJaL03mYDQifJEJogobYn4i5vM0TFAzlS/MOH/RA2uZb
7E4naRkuJZHA0H++SLwqjDsAv3DZJkakZL+IdHDAgUW4q5jZ93JJLHiRl+M4vtlf
JKITEymLF9am2cTTvGhdU+p5kSxtdaAldes1+CF4hrtVSisaukyNmG2QliAaoXiv
8ZObwLQ5BERgjBNX01veyHsV48TzPuM0su3xmfDwh5P9AE3KRfdC09liH36Vi53s
GbDS0qP2Nt5AAloNSMwZ1J0VkJPTnRZ+RLpsvtlkcLeCqyrr/mqAZv4x1QkATe7f
9b8b3VzVwZfjSsEtUmLoDgR/DS98EU9/n2Dk1tWARI+SDMld4G/+ZEa74k1T8noZ
MxtNShgnvXLaowwoHrr8XCG3DBCppMFyxJtUb5p9sSfIAtDXOBEjli+gOTUb1wwA
ji2bGIlMJUXGLMlKWHSLVXOsV/fSumufECVDT+QHcPiunMvJyfdjMqta6Busl3qd
1UJVBSDk8Sm2Dw+9hv+aTuTuasAD1C4Weeq9PdU3+A7TtnpFTyVifbo3GG38+3j6
f21x5pFJQ+xcu3edGAmzYp5AUYe536iKCJrqaIvA9CsjDaaYhgLf6pTnsxMQDygR
SKNbUsrdF+3Xme13jX4J+3TSlSqyOI33iRVxK563Y/zWXG7qXGigCkxCT1bGiYlw
s/CYM8NV14i5y1MbDdYGtS04i55CeAriJ1syoMf7HjqP9eg94xO4WZE+LvIKhWL6
7OvCXwPJXtgpQJCwKJl55rr2+aBIpQcOT4iqWXKbZE724UJcYZxvcfAh4BKlcZIX
NdKWhmh3zIYPVf41ua9mClBco45zmy2+UFEtACjoG2gEjP2aTOtnaQ0FhIoMg05o
GWlPJ2D0U0DpnulROKnsKlVz+OTxOlzAURDqwpcibwRJjUEpqplLtsVDotv0uHl1
MUzvIjc55VdKILtHbLG5T3suE3gsSoeuUEMmU4L4VbD0BmJt7ZjFbAiwnUSe0xQf
PFGrq/cZZJZIm1n91kVKhTCfQz1jlp6uf46PpdZGlgSCWgSBpZrfAJ5uZEuNiGJZ
2ajxAd09o4fngGRfaOG8bKpKbTxE7boEK1ac7oHHOw+6QzP9NBqI2Idj02pVgcyu
7KJInyueAKw+QSuJCpBq+Sqov8dgMGhJc8dDkwQy1/xfqldF6qKdJr45VXZDIS/k
q94Z6TG/IRo/wu23s/CvH2pR0Xaa3m5CQbKYr5dTZYRQKQUzIpynTXx3H8l36JVL
+tGkv5AQp/HIV1/Sl4DgigwzAWIeKbyRmgKbp2rLO0nXFwZJjuDmHDhnuZYZuef2
ck9x3p+bw9oHnkZ+IyO4Eh9uiCcdCO9Yv6dz3kIs4/rBwWqWJbVe2vZs87JFwTIp
mN246Fy2KtVF4bLFkAP+XTETqJrDJVW/ehxDq0jbunDLd2tt91TWyIu+Ah+YmD6E
FOteKtZdeEA06pLIOjNihwO0oBPBziVGvF6OvIfCvk9z4wozIp0vc8hu3RPk6Bal
09tNQFrSVZOBmURADY0zqm6sOADLGKI1cFTjEXEw8eObr6UfmZBXLT5zxJu8xDG6
uc2TKQ1z9Sv8D+yGmkInebWqmnLlbBCe2O6HojTyk4D0imNKlct08aT78X2PMp06
b7xo6H6Ceh9jdz0G49a/e8UVNCwRihQDcNoYe3W4gRNqMTZV2a2k0eSnQqVR4f0n
4AYY2bvFCqHakS5E5rTxF8CR+tygzGri64IQGvlK2da31KtvP+ECP+du8xAXu2iy
OBXt3saDh+/3hv8bY43JgOFCC17FD36LxrWpD/kEOQZYhSJxo1mYqwmVucWZY7bu
B3W5H3xH8R73cxFHyz4aqQe+2mLlCkcnYGpLgIymYAjxrJ6bK6oPDdp8aBEXkzlc
iqOiNOhQgLTPE7PKiIw3Urrbhafx+2X0s3ZJeq0IlGAReCWGYCDfV12iF6x+oyVw
fwkt/CeMkYmgXUxwK97Erh86K5qBDgJIHKNAAic+mRgZj39gqX/+h8Oz/Fb0sT8d
DCnfCRTrKGKnoLKMltlf7+ZoS6TlU09QYdrbdGgD0hTWyCVoSkQ5DY92zc7jLdmZ
PooT4eWMPJBz+1Sqh4dp1Pfms86/Xr5LuY/IAI032YueoZfMc/xgSISFUv7UB5np
J3PKJQHi51wbRsBk2HWrXZZqpbSZY4/rk0ZHxNLfzZ0Mq1obkBZxADqAqMUi9ZqE
vLgUD1ZUxxVJ6nmRCx+d+/tiFXnz4Sni6hicPKBkyE49RM8zvg7IWqQ7dP8kjKJi
ImZs3jqwFjJIZGTMdQcSkHXqMsAVa+5GU9+xX5i4tblrUjOT9nyDbPcdmjh9NoLP
6xLO2Rtqb/5ac41WFIAOfiE4oFfuWjdWIPN/HdjDT/n9qBCCLLyJs+KvAT0IfQY8
x5w+Ro+9fspHhsnh1hWdnig08esBujcgHQ7abAuiD4saWz+nksnCLMQ0CHDVZiel
GbzyU4unCitRIsyk2poLuvSXoEz4xdp6TBahU3vQAiYZwskQSYJq+kKinCEdJKDQ
n+Z7c06wjCzao8f+dmunXto6F9MS5nhDm3GQH3CqACCrs3/QTMRP5YRMReN4NfPv
oYLcCVpnlYM7hYlEYLRXOIFVo6MJatiXnOrMKx8TA/wl3Ml2wpcbBZTGCnDm9pyR
nQNcVjb53yaOIqgP0v/O+y0YfyWSBJuxiFbVa5DvI+FZqCes17JlajtPj15TQ3vC
OYwMYsG5JGneqi477KO5P8EJJ7ZhuzJqPwCK1Sp/xD9mA8WZb5Vb8jby+bGXMnyk
96VF13yrvjUHu3WrN2jr0HikudMSAEzIj/s0cyErH/o+NRm0agjHKg01+xZipniT
eQ6s1YGg7dP9XwVybZ6fudUNPHWGDE04+au3dXKRro7jj5Xj7eaHzovIVPzb3TTS
jtdP3OvStp+MVPHl/06LpsDPbefdMR5fgMVuzc3jZnWmZTNItlVuSNsAxOHiUwOf
Qi7rzRxq9eTPsa5rDu0DZvliVkjM1jnb1AMWIkyhsOAXXMk+3husNmXr/pwqpUAo
CEOzgVgJBSZIMIH/S/G7l2kOz2dG8HJQghdIxXg4lWb9IlRx5LmAc2mnPl8rEF/Y
nJDqx49bvSojCnloF7IlHVgFfCkLLQUFiBnDwGGnBtgBotfJBy7YFxJWgmT+rdAI
930OFKOcbUo2O56Z6XpxmEEeHcamJIixX+QcMLBWml4eI7Gc4KFhaHyxljlz58gP
0GJWz37VbU8dsed3eyh58hGGpGWtKcQs0bAIUGvNOJViCfXxi47UxJ+JspgeYfhi
ktZrSiqPiQhVUeoXxAPSS1Yh4jnNDMvp+T0guAHEEseQZjO3zva5cNz+j/fsq4Fr
W2vWt+7F1fwG3LPKCQjjHZptNqTcI0xA4D5QT0sgyTMIf0XcF+nyQttWvG9sItWX
MBIcxb6BcMIQpGbPM4Q9on7fLokzicCcyAWim2KaDK2B0Vko17ArxcmPFZvoX+jA
PMjHqQHYtI+snjncBiokGYny4IN1DtvZjyeFwehXu12hKX9pfD6yMFoj1daIH/nv
V0VQRe4Y9B1MfLjD8fnpsJ+IKQP2oh/AI98Qhyl/xmskYTMxgNCizC3LbxwAY9Oe
3Daig8U/O6xHFjkG4TBk463e4yWvKsULcfeJfdzhGnrmGQtU1eK+OSnTowHnbWPu
cwk3MfOAdXv+MXvwgf2ovOtKlwOnDb7eVE5vipivsdXvdHxgiTMimxCwXr9USd9Q
PDWURgaUih/dY+pVqt5Lt++vbdBFKfQdEw/cDxK/mO632Sd+LSFChFOkkWt5NB5y
mhB13UoL5iMSpT27DPP3ywNRd3qTwHnED+7Y8F2emg06p3sIcINSG7ogzBIyXD5P
EptJOmMVMmS/07QF52H+5VamtLMxgPxjqjtfZLfh6wFLuxCarrqi11tl3Gd4xvcF
GrLeeK3y6gNEdm/gcNiOy84yms7aY0oAT6jj48sh5bq+VN68xMUwtpL7RBJOmSoe
BEphZuLLqeYb/hpFpoNpRPhu7oF4nuivisie01iXKWfeBZAxsg8UBDMowyZ2Ijnk
PqUOf0/qm0Q40KXOjJhkR/O/Xh8Nd8XRCCyZNlSR89PtTuw6HyDOmRkjb0v8IBCo
wmpyXMviGJyqAsNingpB1GD5pWR9JA9RavdDqDk/YdlJbgt4miSke0D7CGPKX5/U
UkMu7MKNPoC1Ednx0xfJIDXq7etQ1P1HvC/PFulvcFb17ZPUimV76o3osc8AGND4
w9emF/z2hJRg16/FoxWTFGd/qb7PujAAVI/kYXJ2ZqCI0H54V59JB+di0pqZGzWC
M8+M9QMrpxvy/vyMFnsy/R94W1MthXn+IPhEmwzlxtwtioubQVZKyW2EvAKpStxQ
5G1ITQ6IHeNlWGxblRqLcd3YJamWiL8FBE51h7ZOLA9AICpjtpePO1RM12uCw+tw
9X0A2LqJJDA4nhJBSBLMKPOrRHrVHLIGvkM02/GZFq7Mpeh+FaxKADi1I/JpFSsO
9KOfw3fXTRXPimXAKUOPwdaSzMgVO3pt/mVjvizaj5Rl+a+weDdezD0jJsoWbVkf
LkOcdV7ulYD7aiCh7sQykz/ZuMT46AmTssYNWqF26M6F0qgPXyAbk2mqaguvBGgJ
/JLvPkYJc9kuNPSMyj4Doxcwby4USn63gCBpJivGEfinuRQszVxoVQVRLQD3WkPa
2tmxYfRtWRpuw0AlToe7EtofAPPqB4HUOts/BR+cFLCwNnCXiC1mxlPcCO5+OeTk
PoQJ3wY7uLRC57149ytuxNUeLTQpIcASNXA/Jp38uZbunqKX9N4O1ievFuBZEK5H
F9yf5cBl1yE9I4XSLcgDRudWCMfVEcmN7Jajz+46+zEDC34vVTyp3e4C3giWG7OY
D/vk3qPmEByvD5q9s8BHOtpcGhYm1rvHOR2eKIQgc4HskAYPeg0xW3ak8niLK6sr
0XaKV7Ppg5RzRLDbEeJszMpoq6kx0vOaFc7sXvw+wxCKl4Mg2vO6Qd7fYpHuVuji
YG+2tyMB86eLj4b49AXj6OoCNPnV2mOImjrhRBpaioLWZ99zKbVpByy5FQekBLUN
z88IojpsNs1TWhoNm1Tah9uNdaUvYNwvMRHYytmGqdPZJBICFiVdTA0LX8cG87iS
72rbHBGKLfnwwSOfqQ9RAknWktA/cE+wvkowFalGBIsmI+mpMptG/QFwV6RyBU3z
w/jaY0mH5iBpHDBzVRh5Q7GGYpSOUzdQ5ooBYUM8JltyChKY+CwB2Ch52Too2Yon
qImUEMavaCOhcCPg+uMTWP9BU8u+AGyuqLgR8un2/nm4Y2Uh4G6Yb7Xs2c5iBiAj
nScoyS0wYR5TPXGxQn80bIzU3/fUC1AC5ngIVF5ZTzY9BA/B1M/jHOcOJMEdOROW
ESGZqiEvk3amcsLmS0S5hBxnDezb94QqYv4yGq2fCB5T70TKBkVTyujYKecAEkbq
9CcWnolN8OaxeVsnf+v6QAkve/DdHKcNiSoEhFmi1WTFzXRUieKoZuO+zT2PdmSM
hfJRd/OsIXZRiHUstf1HXA9x044EGKTBEyF/2dt/uTTqEjn7EyhVrgeAw+JdwIGn
5KQULqK4Xri6W1pOoRqcaeC8kgTr8sz+iqRBdJlmv7qsuMDhaSR5P2x9ZvmleOLS
1ExLT8fD1erwE7aukxwsMZ11Nd6vBvfSmwckycJMikeAa7MZ357j8GhhOjjYGcNW
acoRRjt39kSA3gUh5Z0ML66ug9Uy/uy1Q301Tz0zMRyb//HR2nFO0DcCM97eXn3e
EPBvWNYKNSW2NPqJ9tKXpd5TG8Odt/jOJYsE7HOQBJDsFz4DyXBJRwmL40g9sgRx
nOeiYeNejnk+2Bqi/bU+In+GyyYxMyDvdC3Jjsro80e8DUP9Q32GhptIxJaKzo9s
3kYu9N5UYMxRBdQ8LEUiNQpLK/qQSMZr0AzmbR8gXqiB6M0dUYeUr58keieJNFF0
L04bPj7sDjt16/akkSDv24qLIi0C7iFbsw39sW2WbKQ2NH0Qe0Y6xj245pAwS/Ng
cCzo+7NHY6o4bfivcBTONjr3Zb2T01zBCE5pAgYIP5UGpfVJqtbeKiztxUdzF6S2
fwp+yb1xGS46gcF4Y0upw58CSIQalEtfBc8Hm70H6dv2aIRQdIOjNcpxq5H7D6OY
72+m/bSQyLbKNoaoRCFcv0ebs5oI0Zp/cgznUY6ML3Ll1Yxg5FTNu41K2TooGdiT
qlyLxhEGNQhDSSoh7evGHSA+nYqDp6biOTwUq7x6rI9h9kbg8PIE5AN+22e6Ns+c
xgEXgF2DYoRTi5/9F/ShiL8bjD24TI/QAiKEbVogUBYmyigDAxhF9x1+CwAPXuP/
ugFkLUbq7HyhD1GXoADFCSqKN4AP6UnFZjKZhbMi7AkbRD/S71+f3PvIkLIn7QI9
ssxHfck8LDdbIV+jrJ6vWeZrw8rCFKQRlG8aZ77p+HodDN7mdagWKykwhyWtDbzZ
IpanKebm8knZ48pc09OjWb0WP1OUfyHT/x9BXmCiKMW4rrHgScyB/5m7SDe4Q2ak
VQZ2YWmxYdLoCtYw3s5CtNZbcT2UgEeLT5h2dYh4fa0i0K3y5Bsmj4JTLqj12XoP
LFehls+3+/w5vJ0oDU52ts7aoCWi00EJDmwvvXRgHXhU0L7wbNDjtQ9XIpHoriE6
KVtL5yX/+kuQmIVXb3xarh7utxUDI/Y5wJDT4In/n0C2mdVboTUK9o5hKAlWe1sI
r/lkinkUqdaMepStJGFNMw2l+MifNWlKkN5Z8ZqAgqFQ5QCiwmYRdShTyfxxa1rN
ouAG80LsM2kY4Zmcv4585QJ7sWhLFmEU+38+kYe3GH0bFGObWw7CpM+9/DV7pYDc
h8h9kP1aCC5N93KN++665b9+37iKpIL6ypsQJ7X5QiCAvqcRBhiScZnyhssQyRrc
DwfmU6Io+ef1RI7xDyQzCE90v/lpgDclbgxJHQscm0ux3wbBzMjzr8oc0iQaCZY2
L6wIYzZTXvPrT/NJTg8ahQtuqF6R8aGqRhjd9ZwGWtSOyuN1ca3adH6dqK/bvT5N
dRjJtOA7wNGzyAuQUye4qSX6MmA6KnruwnYzq7g5lgMArNwEtoAkaoT2Z++6Wigd
V06XqHV/ren/SOqMwvC9SHI/+9ifMqUrIMO9o//F0bVvaTY26+S7Gc4Tg+JLfope
DJNww/mxlocicC2IqAhGoEcsmrva8MnrQLo0ygMdFlvZICRFhVmG2WUoKlDrTUje
qgaSdUUIiSAsI0uhk6JldSQo0UTbN6+1oKjJzZUFJWW9D3weJn/BHnUQutY3HBr2
AE3PXH3j46my2dhEj2Txq6mKrPcKyTjmKqkQ+4tB5FeGeljz0BgWf0HQXLCePKni
/TdiZnLFWGIlVC8QqFSNLslzlB564D9zwmkvQjmawUTlKyAugUuw5tvk9OVGMOY9
u8SPX3ME0ROMsk192r5Sbk4YJpIhHUgGskHKZDvxy6Mu8PoMScPaRqyIVI2DkUbC
Z3rHR6MXYjj1p8ugycDARMx8fgPPBGVoS1g+HV+Z6AFyB+AqthpRqcZLQ9u0EJ9q
V6FbpeYfi95KE5zYIXNcstULOFtUCu6LksRXIaMwoh9tFhtWjoBDA6Y/abUcOqf/
jpuwhFQ8mM+wsoZabUfoeVgp7NJgjC2sxtEqxatiX7LLEZuNtAeCRimj5bz1/OHd
5GoBV0Qy/AoyHXmUyO4NcZ/fUVoYhWodt585Ct3dzos1d8hr6fAmmAbA4xRtUHhj
qfCcdPJ7xl74BcbdXtbEdBasSSjM2br88OZ6pce2ZInUMipREEPtDTqB3M/0WwCm
buYwCbKIZcFDOmxxEiOW2bvgqo85FW8D8y9X3wgTK4RMApkPoCsEZIj0pjHtZ0bc
hEA8fcJ/3t9QlAq4wvVT7vAHlt2UoHHxf4TDpHEkGtcUcvtU73UNeFPDAtNkqDrO
Vr1+5jBBIVhy7iwOdUlt/8OH80T4x49jlL/SPXttfjKXVH6OR1/K2pyOtXqeqagM
Srdnm/ybO4B50KaBh4eH0s6TQzULSfeUOnOzivxbcsKsPsTldqCkhn1i9kEX7AAR
RoT9cHVECbwnLBpcy1kEMPQzuKgvgMJGl++YcA75KaAYNUArKEm47sVxp9ZVRXEe
tOxvzvuJ5QUuksVtnLN/+/66Ut9zwOUcOuKla0v8s3tcZ/n2ITlvzBINSs0rPLZJ
b5oePD3TQpXJLVbYznDFw1AWKzhjZc64twU+3VvineSjBF3HDIxR7kDfuBZV02p/
XcLKfhTFf8qj8PLzBvBVjRj60uTDiyLTiWHcRUQHQu2h07n2q1sX/+rZY1+GBcZD
14TrZF4feuJBT6imK5yy2ORZTB/cJqeAOshuZ/iB/0QYDwhKxUfWXhroMHG/Xhuf
p2wtdlZ+tcHnPwWt9Z4TF5sXhJNqlIef1AtRMzpIUMxXNzZZZJbCBi7wxyCYMFBN
3nYJ55opihSdHQbXqA2mizF2JVZN+diW3PSMJJlNmXOb22hoe4ekDr4KHg1T9yOn
8ogUs8yRP7vljozYp1MDIVvuDil4yp2KfbZOXok9BHIsqsTfCyWpYCJMW6RtZjjb
CxXSjlPwQ7qw6u+hDWcBoNffUzU65lDopMINn6RQS5QsbRZj2KNtTukesB8tMA8h
gEZS31ylibIFlrzzLxpt/2ceUhA7cHzlAxhzN7IlQZINv3HTXeqSRdFSCRm1YWyI
1jPjAHDKDbQ+SDhJNRigwi4p9lVBKD0jYWhg0qc9mdVvBa27Gd0KmClVBe0rICre
72cVN6UBTP6MUCY58jpnoGPlRaj+qkrnQVx8H2Y1LCW6P5yjvlRCuLv5YJ2SjvML
J/v6InQjBFrtCKmwtkja1fKSMUH3qWihsRmzcab23KoUS2YNoPYnoFjZKrxnhLXR
emPklJD3Ohgsv7HRwr5p+iccvZK3dNVzuaNt8TohwpFFhUbM5mk8hqoPncXkYwlK
rDXeuDwD6qbOXcDfkTPhXvYc4NDpiahJu2CCITkUrUUE3tFwQfahBuQm2LRj6uLr
xSq3ce6LMZ9Nat9VFYR0CFoVozHN1tLjFRj5f+q1rm8a0n1y+sDW4lWhJBDICdSf
j0HTevingW044dm5Z7qtWtZW/o2Fd7iokRWF5yXYQu5b/nPpsKYwEnITT6dBpfDi
D72TjUtgpRoWPaqXWJyy/W1HfUj755SNaBhT+czsJTcESlnwG0OYHcQMCbfSa9UF
OxjsDfM+qxLdJpMv63u7yqbXwgu/ATXUbkrZc03B/ZTr3p5rC+8Ur/McFwq0UHIM
y1brxMfHQm8i64IVSICpdNmEGI1v30BZSwPPI1vUg27ptOszfyZpcMv2g0wAfnpy
D+SQN8efZa7sdmhs/b9IE4xexAplpzN0VtBkVHZnzzY8OE33j9ovr3J73lr6gapy
eq8hkRppnLgmFMWlNkarnscrPCtvJCrh1TTji4ZUKZcej67c+4RVwB0Ymn2m2/Pg
zHmOoiCHm3WeSkIsU4jVgHvqAvo4CWT+VtN6NGePuAFaIsVlFkRf7vA9dqdPlM07
cJuEZ+ybZeiqut2aSvzoJYnonPLsI8R7dnJBKuMtQ7apfQP/SMXWHG7FN8SFiSQP
B9CMbv5rEo61ee7yc/jO8dqjypUwXjBACp5bNMIOT/1MfWqkfsn9R6DkS35nxmdF
K/wskIDH2pt8ZBqTXG+WPvMhwcht3ug35ojC8WTov1x8BCPd4wxFjBJ7ZvgRWaEs
1f+uQsMz2MV9p6opSOp260l8t80gsznJoJ9arxyAHxy535CR9QnFhIo4/oX0nuDA
k+Ka983V1pUf/jtR4hzQQ5qWyMAHNpSx2y+PchG1/dUATq6eTnx8gqpJdGJcILfy
CuaI51V2j/eu/Jl0LGDiQtMR87TaJcsIGX/Zt9iFU2Sy5KozhpdjhU6Hp/oaSs6y
KhZOg0vRu+4jBCZHm2mog81985OOSPvfZDZn46/+SRGzcecf33+TEaAQJ5CBCLqQ
3UApit2hkLWz3XDeg2SkwrMe1Y7IPhMW0rHl2IlknDuGMOhss7lSttxeeoWPWJPW
AdN87vaUWahiE9cdKLumvVisOB5/BbNuloFxpEXvBIL7aiSW1h7uHMfv7Y0//oPe
nzw3X6hyYtRdxkLByY7QQtPnUC9gCoz044ypfLtrV0tEpiPXxb6LrTyxExNK3UFo
RA3AVSopovWG6nHS3/6PcIXM6zTDP+C1T5PEb6obBY2Ue8xjap8iu3un9HvR5Ukk
ljvUiAEcuhU3ccnlkIWK+FGxCLULbSDsbM8JZn/PiAg8yQXiKzUkv00vK42u/bKU
9ZpHHQkByxusuti9Bmu5CqT7isO91O3x8PjTomtGvUFbEkGE3W8tDshJZBBgKWtL
FthG6UDaI/5KLEj61+jTi8DezKCnqzqYRiKokkMfFgw/nuXuwx86grNEwZxSKtcB
gVFcjtgfdl9nUeMxWjoUvO9zOB7Bqrpp3c0EtbT2QZ/Z3U3bs/U1bxgOrcuXYump
HjI4wm6FLDGdlnBfzvmVsAqLzxMEpdeg7+rozopaqwiqorG1ugAzsGFW6tu7uHob
dcBtypwEAnTAsZ32+iEQLQHydlEZyQTj/t4hwIAWVR92Vhy8Q7XLjxMwQyrj9fia
/ZDTLMoegSvYhXoiJtxZwwcVGCsevwyYO9YjDC/Ore37CC1b6A6OWGoBVD0QGqfc
Yib+FsDEzMHawa2fxJ7CDVWispwTKwnw64rGqLV5xEe2e5Cj9S2d0c433g1PmiMT
OsPrDCpzrnYiKq4LWRJyf3llXnklcY6vAzao7ohbBcV6n3H7YeU7V0cbZ3Ezxbpd
9uf3GQKNBzJl5/pUpeN58j6yB76w15V/8JcgXi+RUbuj0T7StzissGO9+UCQkBjN
bpZ+5L+g5aT4aYQgVuyHuYsWpbuGa0mZKzz24o4QelgTC8xUTJCIerFEUS1Q4UTB
RC1SSrfOHcAUN7dFUg2nv4O5TCOPsfkU62jMEV3if0hFEhnYqOvIUavxwfkP/LV1
aL/QlUuxWi0k3gWWUV2I25IjTFsmzM2bUDZV+etfLa80ukREZuA4nNCJFEOAkrDq
EQgAAWCv9zVUEdgGHX902sKOyIIqNusmEskW/PZgwXzaWeLFITTerMEfb45QhL7i
kqRLC0BKijR0W2Ta2UoEObT+fGwYUOO5U12b6yLTTJCTNJI27ZGtuIZKWn5Mp+hb
CAJe3E5X22qwnqDt0ExKLtIqCC9qUTM+SXXl1iASe3fFzyeGPGdpkLWYzNk2KlPM
89lVmRYvBFRSJCGkgAv3GKlBtgXNyKa8AXdDZSKKMIsULZ6RJI7Yk/H6Capz+2rX
+9THooypE1K15Hdj7prV6eaf0869rkX4j+zrpHUL3I9AahVCwWZS5QnAhVbQaWHO
2sbOq2OOMf5PQuj32E9hferR9hvlyfyF2RkoUh2fkp9EujzPXryr7ISajXPotFiO
xc6cd2Cg/pr2RerwZptWJUJ/dHxyBT5qWg1nmCmkkLqUIXFDps2u1cNwYKXKPn2v
1OUlDmNE1BkokE5E2rqxrAgoqocO6hACa1BTeKWkwNeRVx2oQEQuAto1Y4JH34MN
xL+Tyeh09WwvCbMWhyJRFT4h1EPRPRgrT0T648ZoBHGMBCjDvqgE5+KcCNt6p/cS
n8rWhldJSKedgtGrGnWu8TiHdxVu5t0gT55o+SduIGg7uHNPU08bnBkMQW2P2Sot
Zf2PGwvZoWnIOqcPdfqPYqaZAyYKOUhB5el6ODrrGK2v3nAp9UUXyZTOzSTb/HJW
5I5V4rYqpXxGD1/rVHRjXxLhUTB5Nnrlh0OdXvGwSCBG7CzV7mZq2YIUKPOu9/Z1
wULNsZ7Xu3+JePfyhUPYCbzAdpQhkUH1xH4mKLtSESntIbkBxNZ1Ce5lOmJK3m3j
HUVFgNQwb1DGhZ+ZlIqiLb7RnTXBTCnB2UaiZxsenq8PAASMp6FjnQZew+P16kyk
xjASeJhYk4Xo2BOh8v2AGgrhOCMDl0RZaHWCV6A/Frk2HsfBSQjG81sjH4EVT1IC
AtfaI5ByBr1cKAj3YYGBEikheljQyUT/EmFoZziSGJ6JALGtHV/5Dhro0CXYGv9p
yDGfd7ZUEXurhzGpPWNq43fDARcn5/lPUvyhCEWJuZAjCMIyNK4pujHx/2xN2owV
5yX3CvW0niiI20DWJbxJUtHiXxz5huqC+533dNT+KCiLE9a1lJ1u0sZEz+UaxDNV
CCNecQi8UNJ4rN7hqJyWKOoW+LzcsolfVq4dn9Sgt2Gos8Ab3ZUevsZRt59E2o0A
6yerywtrUdgD6P8sUUGO/bV2s+Qyo+FEQULv3/1s4H6Md9VrykkcVxu1qtUY1PCh
txWqVf9LThsA9SWYSWMAm11pyCwGhbmydjMLqOOvr1v0CBVMAV8psH9l7UFUwBz/
MIlmewLZM7jUHgyZZ9u1anonxJlwjQtV4ATabPIa0vxL0kSXnnbZJ/nuOo0jUxWG
zMN16gQE+BLcYh9qHMlgojkp/nOpmzjAYSwpQSpGYgImKRJBJZuQTM437Xk65vlc
AHkmlsOK3B/awenGO4Y6qmMiTBPE3wOAO0wE1PBMZXkD/uFS0kWx0sP9EFs8OVI6
c/U0G/iekHJn9eLDh2BxKCndijNKauf4m3waJdWT21BgUGBWopZni7IXk0KgVlQv
xNSwG65ZYxyth+SJrdBq6LMqyLl7mUDQioDhQ7xWWL8auf2iiXbwVLafvQ5URtXc
wERiYQJwsfgVPpZ3DNLzDu7k8+KPS1+TS/5bve+PEudxtXKTi8lwT14w/wT3SDFE
OJkXkaJ5Q7cv4yTVSEUI367D0OEpa6jqXy7A8gi6fOp1W6ojCq5knglfA4XXMFqW
l8bAMMQI3eQW4QBwC894foKw9FJTHHgp2qS+3CYlmGI4gu6F8dygPxM9HwGesmaH
bC5tcuuHi+cQ7tOsjsUr9VqFq616U3PHScv2SIQOcndZphRYJiPW1l+wZT5E/PXU
x6lWCRNjguF0yvmYm4EzvDZKlc0M3ZsGtUouHiq3Aq37FFT3XPWEd2Q+yGx4iMyu
6UXf2E7SkrUNZgjlpDstDhOOd/ARWz3xkBmArMbvqhuhVJWoJWxzO38GyaLMdFSK
g+6HcpAqUiv5mAU5IAXXSeNpdOM7OWlBIVISZweuL/2Yf+BpkxVeDOTI/bpGU8Cl
ZzU1cpkpE+0wGSbqSgQgooICRzbCQrNaS8LlYbWrV7xKVfVNEWwsbEjxwOp+NbLy
b4sYROSyUmJ+8UTYoStxRPcEdtWzF5uh8HrAy5o7y8QW6FaTWEdnMPp8BK5wwgOg
83jDqqj6LcsprDYbFjEvAFfst+suHKXj76sRfNOjPCVCimlmAwiXUxWXz15xCQL9
g8Xk7X+SYhuXTPLUA1wme6lQzoSgaPWtpr4ZN1A6nVSIFCPR3CjzzDHP5qigt/Uk
SMh4cGk6dUjf8NYRRIqH2DikkUTrl3Ph6a39zEh5XpR+MY0+YNtADFDMKsjygtCp
ToRzcbfGYxhShVwvX/QIDJkqjnxjyOR2G7w1xwIAgZGQMvNPA92f+Z/DtEymMPdN
fQlI2WnjHsrXK4x3xsI8/7sxPltIWT6MfJSqQsYBFBHRQD5g5ed9YZxN31D/8VRK
Mdq+XVjFBxtlQZN3Ww1wZJDS+sZilqLWQsXxlStlVHzIPMM8j+IbLBP4lmxLw0aP
YT6CYi8czgbtPvvAOpOYc1PnUdIXyN8+GZzi4sUfCmmeBHgCiThMfvZXtFB5Cvq6
qPsl7BU4C3bTBABIfBtTuCs1Pe8XflmKzf50xg9iAqChwSnJkssZqEQpD6bz4pqE
DYN+GNLew36i9X4LteiZ4dyk7e3ROFe+rUUO9G9w7ImS9XvnFGCj1k1iR6U8ynTx
bNXFBjq2bQOC8IIIlwuUSrDP6bnvDcVGFkuH6fzyevvZpFdi8PhncnmF8LBQQ6rW
Xlecy8DafRxzzEHBizfQoI/svgLuDavuRYmhBs/JMHZGD2mIkLlK2KreP590t8xC
BsFXmYF+UpzF7FbJwBkjxJzh5Y12DEabW0tJCGHoLpNs4ycCTsYA/0lcXoUMhxf0
TK6jorAVDpB7TnJ2PuJwtHFoD80hB3E4yxmTIUx4cci8RIZFJLUoYSqTrcxw4oZL
YJ9MV0QwfpucfayOPHjtD0Cj7KlAY0F7+9/qSDgbFxhJILSpcr+wGMs8lhNdVtyE
+0eD7OSU7WfO9GgZlpilxKzMweLepSjB58/JrUIrIsCP+DmmV70WymmWDAI6p6YH
+9Rr0aYP2anxutDueuepN65NN/UbQ5XQe5fWXtGoDiTw96VXd53E9MRfFGE7mXPE
bPyg4hURIhu//fLlCK+m4vRDkSqNXByD56tdChMUSlBEqI7fTIeYAljNUOkgR4ea
D4QOpxVjQG55lak8M0ZCei844YNyJjvjFvjX+TIUg5k3iQsvjDPfwaQsZXxU8GLZ
XR6/QlOFED40KpTSPo/3J2HU9TDqQ9L7eSDvFU9wQe6wKktnuTo9zBGMfkGNnKRu
Hny7got+BAxlFQO2On6GEVaHKIppcFpgBGETFQ5hf6+bsuXrOyWVe3CKyrLI6V7+
8pZyl1JjpeKYKiP6HLtm1AIbyoeUqgxccAGbh0g6OoKO/15Wtsw4Vt+y8BaLnGhi
wG+X7fUkSCr1AIFn2uYW/ASBPmO8ZBnYggC+EkVWyG1TpEIjnrgjAD7zMmubnmFv
+9XxTJqJAv+61Zepbf9RT02v4pBoBqTLIPBkmuZFqwulBUPuVEk6XTw9z20rqW+X
6YdpbeU1N0eIoUctljTDfl6Cg1KH5i1VR7WCPtrwUKZdlQyHgfD5ZQv+9u47kI4v
If9wMCaiG4mH34HoHse/2wHPXD2Z17wGpnYocMJAwJhgm/iCALObzlIJwSmaLn0q
slbQYkoXs4UVjQgb/BsVPDxryZ2tBgehpkTZhYYqQnpTAJoWXxHnWY86IJCyYyFm
aYDwbuBFVhAeDybD54Wli2WSAQfnHMh2mQpbaOds64HIBMMoxhT8+4DTg6lgWnJu
jBuCyNiGIAi2/Q9/WrnTnkVaVhqQfIlGsCBJUwG1i7kKrDlk+KtmbUAtmYwrL8aX
RjdALNvl8tbYPV8suXBaL2xAs2CuthWfNr19GMHYpIwlicZXaVqhQ8qBHBb8E1NX
WPq/UIJWIcjqDCuA7l/ISp84qD3nwLDs5AJbHWf80a46YQ+pm2Fe0d+m4uaFm5fk
aR5EqfGlAxB7Ery3OduO+anPcMO4RvJcskQYxApToNAu4I5jkVIRQL/Ga125z8Vk
TGg8UXOz7CYapcgH4bfIi3ULWFrQFEbuMD0tz6gfHIiNntvcnhYVmFosvoQbUHCj
S4L7xl21IbD4BnKqEsAXVVnmS7DGW/WuZCZZ6g8NpSMRGmF/H69iVG0P78xi16ZJ
lCT3EWB+28bgxkqtNsMUQPvkUjUJeA1vdzUoUEdSvbsF7MhKukd27IKlQIlStd1L
qWqiIlx0UuRMyB/U78WH+FEnDDV8nyspZihnmhPzUqZDevJ1vfOT7SV+wwPCtxEv
EPKP9maEKl8p1ZqY2ke2LkNCXw1rkuCZwgqAB9C7ruJCuZWZJSskP3DURxz7yC4n
a5g+L0vbCgygeuF2ZHJ40A9n5VNzbatkSJuXNctD6KDk6OSWBRVv5R3n1R4yIejq
VgqtIqjpU3k0mUxYc2x/i7SGj3HOgxJ9hFFMGA33TD/zGarOlKS3cFLbsVqu3ZE9
r9bqSFwHYFWIjRq3/NCBs+xAt2g651ftJQRNEpAG/kF5Q3TSD4SYG3iEL2i8M9Fc
1ZoxIoG/7A2toixZ/5asihqVYWdCsFoM+OQp/n26IywS64lO2qBf04rFlinJpfcd
A4tmGzGmbLq5XyxG+sad1ZNP9jS2qR5Q/8zGNY2oE0UhyRffBSi425F9Z8EjxSSS
dhpcH33qe1vjHyp/UpsKc4a7YWyX7aFk5peqQgRbg+BaQaU572emvTLu14L/qXSp
BUfOAQZT2Ff+4erQbGjvuTvDaTs+vi+Uuv/ka+WIc/fkdYRWSksTlXWEAdeFA79f
fCu1PhrmcGhGDF3uN7WANQ/b7AQlMB49pb84moGNmvsh8BjkQl4vKYj58VZIYzMw
fCK6PDsAKsXcIzLLFLkV4ZO6WlEQB/86GtUanzUYe6UbsWIijcNZCIYJYArbAI+y
cWPhyeIBaeg4+G4M8ti82obDijcbt9HoJA9Z8GjlWM74MPzWaGi1uIhbvVXT5S8R
kJapVJLyNhO6hUlIsBtxthQ7CM0r0RRza8P6rt+nMLNcW+D4iZ9BKvNOBx9vajpo
aYwY1Mf1kO9/uv08WQmNjoyhIkqS8S/+0xbA7Rr7RJVuqQXAneVqB6S9DGW7yZ3I
VQ/9pVFd6XATqeh1SFn0i1rXp60lyXTqk/NzSwhTGuZDZKB1DuM/4rFxGJZu9q0z
03Yi4Siliie7aYZHyc0pYKMTjz2lkV82QrKOP3tDlHZQVqIWfDnhuucRsN8pT816
ncAGYgYLd3eo+xn+g17guMcmb5tesiW4en2RYEl16+e+kB6mNcRA96KNvXphnZnl
bffhT4reEZiqIwHArJaZ6GVygZucE2QXk+U8dSnslmrHu7V/m5rMcQ6qbvLmfaRW
zcCZH9B8G9BUu5DoZfjv6SOIMFNPrEdyVdNzD8VH9Xt8avGwcyaqSAeOrytNI5Bh
uyTX1esfBjpLu/N9l6hof5PfRfJxxM9fvexz0ZwMosjI7zlWyFuUj9SK2eFwk4m1
lNs+JE69mkJMHQUQaLhIUJwyd5zjM8pDTifAvTySwePUz5CzD/4YgdQNj3BZOiuy
C/gCfcdUOWcDEw/L0vJvGw1zvtAryyrgkcfBzwB2/ayXJG4aBmV/fjLVCn1dVo2X
nidNZ1XaWg/ORgTG7C1OSU2j9x3IhW0G4SP5hCtmVrwFykLJDyZ5YXjf5NrUDoqq
Pv14TcH0KBdQkL50oZz7YsiozM36dqhZzmlMOMb5oLDYaIMD3YuzHip1TTvRk+Lv
DXQBpl3kDrRD2zCWiLr/QHtZoY3G0rwxdxstXE1dEEw2pMW8Xcyq3aN3N4Ppy3h5
FoolhwUIP4JQGjVfvhkQovGlH9KNeu0Kd0YSlUJ/FGKrhs0WapnPdcYyty9gRcGs
zOV43lNutntf0wPHHPw+dycBYeZ+q6K2FB2I9mAaPgBOj9z1Onv+lV2VfkbLoxLL
M+e7Hztc72GnxXOPAbJxISv4TknlsvzEA2C8JLJxZHptpI5cmnHSBuLTYZRh4GVs
PzDNpIgmVSl/bHXCc77DrxS4bYLl7/4DDSpscssvjLDjzdz3xTUCIbppZOBsctBb
i6y6ruUtG4HkBj32UqHQXm4ZG9/M4N7Ee6d3iR9xdIweh2bE1RWScvLpkK5Ddxkk
I0gMsSH3WCjYMWakI6sKGbR5ey/SxVH7aaCbp/Ms6YJi0SgD8H5Ka0L8NlSoOYXh
VjmR7UH5MhUgYvvsCUJlKFumwSZCjywtZmdE1xCyHKK/TO7EvWBGNVeRxuGhDypt
brYxkfeP2uvPyCclFPMJiyYe1BP6qbXcWjVs1I5Aa4WYlBzq1pJKIIfIFxH0ttXD
TcmwZs5zTazc+HVdLtC+RJ2zRG9sAAIlQYyJLBBeqH5lYWiOYDvOHJMYB7rmi/sU
vZ0IIN3WOdRLFAH8vFmiNW3r1fyNoKc/JMM+OXduIMLCO3jq6beHgB4nEymX2GpC
foypYI4ctZ0tuvsA3oxoOeW5cHXpxRL+8f4wu7Q/Snv9roh6EVD6gWATcE0QX1au
PZlJmP22f5wNo5F8keqhmzDlgqkRsAUrE7qiGlCk7wYcLK5i1QVJxnnhGJ4ilAeh
kJf1W+4P9da77NosdXd0ZL445CkpzrNGribh9iHUrTCnLx8484AKXYwYGcrxY218
P6qKsL3L4BvxtUSfnNVvgj57h65SYUZhK04dpPCbgaVly0yAvy0+xHhtDoORVPBl
hAfRS5qwAvObsXV9CquVX3KwlRrio/Qw4AESBkunYJQnjyiY2i4sadHotsf/ISLx
5ihlaICBs6PHvlX/tByFvGE/nr8RZu7dUqRh4y68QqmKiw/IY/7ajZ6p19wIWLRk
tSvKCRPfhAWCD5FOMIDWyoPuV3U/pDZekXPQ5Uv63XdyO7OYoCEtmjeTLjrWqx49
MoJxHAVqrWffkKv5V1hwjA9Ci7fGU8S5jUT7lDWxY4UjQLbC3cdCN0LyJNIEIp/7
5fYsOV4Qf/YCXR+NUAhTr2i7pceUGPq5n5yetHH8qzq/EEcwkW2IQlWQuKFf5DdD
9IR8Am4URbxAuJE3Q/rL2elWu26qrfuEEeT/2NO8zUyyjLmRaq0OJygqvvxsw4ml
89BzQKpsC7iNJV2fxF4g+hq+V5t5WzFzmZv3h+EelqV6+tiTyFWt+Z+piQUadIHi
p7URW7L1y1KsTcB4ZWAsPJjUsgYhN2PJ4NiXyg8pao29KjPksauWMg7Xg/HuNqv5
qcEGc7CPhm61CFGXXf2payLAvolAKUYfUM4f/xZf7TU8j7qaZTQMNFCKIY2cyYxo
SYfYiJLMA9IkK78CF/ZLUJW0gRP5wwDLE5QYUU7NRYkvaXgZl/hT9kxZ7X1gsF9g
epG1BxufEURudaSLc7TEH0NNJe29Og0AT003MzFmMyCIpUZGWod+VXULmItR5yxb
fmiWYuBrNXLnYYp2CiVmZH2OnVdM4O6zE54KeMAuvsUb4Qb6GNk9YiJNRIJt6zq3
10U+AW/EWlPMqaKadLfB0ZjOUIVzRSvV+0CYA5u9xtYDGG7wWoWhMd6GLG2alVFX
2hC46tJ7TblVHrZL47uEv5696h3HzRmaKtE6FqCQnQW3ibJfGtu0QRFtA3S9Ka8N
lFjjeZ+ewqbhYi2zG4cloelokLFJkZR9BOmFsBY4gMj5pLF1gATPilzO32KtkRXc
R0Cph5b33eQHAHuNTk2PapGLCjyMgJDqt/wkNrvbCFNsyaKhCURuvb0LvgkwkeP7
UvIKzIeW8uJYWR+dcuiNNufXOe5Q1d0jX36+ewZ5QbResmu17yYQKGoDo//FZRNp
WicZOdskKYDSJjmnixvCUiKZK8jNlG8+t7UjjN/Hj8Z0F9JXeSk9YVvmyeRMGlp4
VMuW90uVNyBgl0NBSe4KSYzqsh27Xuls0jdGmFmn/YHF8y+cQa6PB6RYVLCHkv77
BPT46x61grlG1I4h3DZH6tTx3pqmSWyUUa6kbZTkpZdGCs5rUwMINgBOaDUQSwJt
D7Qm4EjcrxIwA7/UC1dxZr/jreOw36OriBmrP1huSkkk7wTMdmktPP6YTsutbpqv
8VSwqqd4la7AmAswS/58Oz2WuSHrwd3078WRsbBoAT1NCKG7uM4KAOZ0tlJFB2d7
m8WrDyosXcbaEByT4yG8hH8MWYyITe2HkaYvePkcsYGNEieoBI6YMeAJXgD1BV9i
IPIfboXbH9BNdwAr6uAhyOUJ640W7Y+dMrQ8cLPisb7LD7X9/IyPHXCOv57/gUzo
GV8crs+xtox7KIO6T/QfkjJ5fs82lJjvmI53SOCLkbxSafKEk3Ps8ZPAdu0qxh0x
BzvigRoKkgGG/w7IdUm02eZnBUi7u1+AmqYtsvk7ZHWFhLFv0mw87k3SqTKCv0Hg
HkqzKuweVq8+B1rzHKRJA/96n6lH9b9dm7I2QjEUdaMDU6upJa1kppR0kW+skP8X
V3BI9cH0+/FpcnUdPzJKecDC1AdJ0k9vVm3K2nUrn4sizHX0SNLi6dZCG/tQd64X
E/GVr8XzntCW/N3EwE+1Eyi5QF6I7m+a5r+9lUQlmzBMEySaLRMxMRQgsaqcTY5r
uI1M73vlNSxX3w0V1LFjULUN5P5J/gWYWOQiKpMhDv1I6Mk1ocBuHxwnaIh0bX3P
8sbsk9WJZVkLphDZpmHbVQcMGs/TUgTqqQCHzEK1WVRMYITx9dbgnUMuiqRShoh8
dNZ/rvU7aoHYmdAnM5EFhJU5N38y1F4ASMAz3PS5QIIf2dw4X0LLX26giv4IxgT9
tIziXWFSfuDQLQCoR952OWhxxrxT/IJ7nC9V0ti+b6rbel1Pz/smBdwmFuwAE180
6f04MGIzXN3ECic/zoBjviE7YeDfnfKYWWN5kQemZYxm8Frx/NMbJbZrXmJ2Uy1u
iEbTHcdntIg/v7JGUavzlJvmnYy+lbfCSVTh8SfJ390CcHCxZFwYp1lSoB+fGo4A
yG4ExQQgXUvLZkXiW8+VsjSFDg3MJzf0tilsqo8MiuRptgi8k1qgS8lSZyhrB92k
IgSEvvfNmczx/eqhUdt7kI1+Fl6gw6LRCyCqJY535Y9oQrtYf8z40xzehIP3Cy1k
40mtoP8Cg4lNnqN/LzWewNX0Wj+fWssPYHSsbC82bPNF6BrMD0wa9Z4eh8YAvX9w
hh7hp11v2KQ4naqmJzhH5i3BU8f/lS2zndFjNXWjaBYE2lxThD83FM3Jbz+8maf2
w8RnFV7TSkfauA+c8lCsKc98jeo0BV6KGVbRBTO9agDKVbJtGNaSZhE/EK2vmhsB
VtUTEiRiZgHFcZmC70sFGJ1Vbj/6OZO8I9DUgeJLJfcqinqduUA1G1BZa3J8SYP5
Y+BeHHuinpjX3qv5LybWVrdu/QafhDKCfOL+4lUBEDsfF66YHw1QnWQwP+Ct+VcD
4Ur6s04lNH5BiOteupOCmtpFOWDIqxkyBiHIeWvVRQ6eST/3/yJQLKs1ELCao7Jw
R3sJIXaXyxPlmBaq/OsKPPQAUUjep1m9pI5GFqqlTt/28Yut4gvdhYwmE01epujG
4xAedV5DV54QFT/kkWilQWVuZs+KcyKh1Aupnd4i9FOow/KGAiZobw9e9Q7TEjzh
8isyS5+sbngIBqJcS9l/+p9HVgWquqSz2bXRXH27cabGPhGjEPCQXDJBJvDI1/5c
om8kWJ5Z0VwgmjDSr7JDUUiEadg+xYnhziyHVE+T30PZETJ7xFIjGvVab8pZNc95
RC9DweY/KQ843GPlbJ+CnB5ezT8+zl/5q+PaEYpzze6cBhBf77v5rIwrfONbi787
36aAPLZS+lTZtwi0gLr9gRWlqnqc1XvyySpmtdn1I+Lms1jH5I+gEo7jZmmItUyI
gzU8YHEr9yXATPPeT9/Yu+t0smd2KCrhUX8cN6sAph6lkv23yxYv3Uhv4N1i+kCv
fcCZlabnon3OIllJmGH7bh4VDaRtf/OLCI+f7hlfpRs4ZG+OwarHUvktdGDbwx+Y
PitY7awUOrj+BhEl5iRgT1yDE18iKSwxJ1y6daxfLOO85n0vCB3TDc2KqeQXqY7L
GKZETkbPBJlsH//sBuQKged0ALS+bh2fQNhibHZ9GBQdIlnlEj/mXbVFXW58sCDF
E2Ce+AIWz/onL4enRzenIQB14IK9zVsqP4PKEZrBxR7U+HIYeJgDyqU+vt7kgTaB
tAW6oW/gAW3DULJViZ4jEMLuEehsQQCSO8xdpMGhDkTcnRbovcRC6SklK9+dHcLa
7DR8iYg1o+QYJEZYufMneax6xWWSeRMRrN0zuWqZDaiNaaM4bwJjxhQggkcKWHdd
kypBVEa36FoBJ+AeYqM8DV5zzIl2TmrL+85vMaX1oggyIictcB51Jkh+rzkzGt11
r42XCjNB9RVjgbIajVLVIJFauInKDsKU01Ndeq9dcu66RvPQDGA4mrE8xL6A7ZYt
MkNBtEus4ATMwkIJHD1tNWxBq18tIM5pjySCGDs3Pu4rZglD/TjX9Ebun5sg/S4Z
r/SD9Zmg6/IMCvBcHq+UlLH3nNqJuzXhPwQVwXSZKQ/ccrLQfyEjopIHameobxBW
wTqs3Yz6gUNHOQjDqc+zV4mv20mFF1xsRupR66oxQOc0TUnEaAyxChKR9aOZP/pj
J4ukFf55rjkwZ1lBbXjzYmjfWHhnV0RJbl3NaR6Ag2qVgQyZ0KvARGvU3Uub9v+u
7aDiVLbu+ZIBXCsvuM9g16qL0VuY4CbFwUs4JJ3D3J+rHSPRMaO1L904jpyfdSaT
lb7pcYhdqHC1BH2uMVjMdtA/5DJkRSGd5jAF1GrUwWsQQUnf4FHwG5eYCvDa/rBe
XimIFCk6VYgJOBGXY1ffr/2HYcsN1fB72KmHL4E63W3G5DQALCUeBCMnI3UkksRb
my5LWZ95kxxJv0DHkg3C4pDGw39GFRHqH1x9kBTgdeVLHYiaznzz8iIwaZrrFs7v
mR7qpQWMquvukm9OyEqaBUGhbsLKvjrKTrxdkvzNDb5ALJ8oV0Cl84L8Rb6CV0Ij
JoLDd4CfYnmOyHnvBblzajHPRGRwl3TES6VzJfN/pJTj7XKavIOv4vdmohY6O2+R
Tgtynme2K3r9kTBH/MIcRk8Jz1bib0Z2fKEF2fNX2DGciRBRK2xKeN04O/1AOMdB
JtvwJ6WBFNQt2owNE27C/L4OGAXGY4hVLKBteA8paW+gpHyi0m+T99AB1bAaG4Bk
7ANLCxyqhXIBfnQKzpqxZOGue+uWrODEALy8vz23WFBXl03VKH5toSR91i/QHrot
4fzCcyBhVBqPNe8ly9VlMZ0xVbfjsAJY3O+6BBd5gWUPeC6MSZqD6xX2YXBaGIEs
eTrvuSIOHB/0FhnVILl4CNV27AHpehNiiWWsoUEcd/KRJFhaJVy/D+gHPAEv+pKo
C1OdOEqYLiZAEy84WC1GtlNLpkgEy/LwzUtffEy6zaTY4x6d5r3iSL1WgZpYaGNK
+z8wEMDkVOygOwSTCtOVVeBA7FF3wZbkIzRA2tSh13ylFnJyCA9OEnyDQSbymSN4
uyTX9aDtozccslaMDIAmcHJaZHDzP6QzsU8R6oi9uteEgZqPzPMpnp+Ysy0h14WX
1beVw5Qn2tXCp30oM6A7iFzbhgFOpS/p25cDg2bAjfnlbE6vQ2pryBQwgNzqAsL+
MDrecqXv+g42kEU84YnK/SyrVrJUituV7bXsDgBfzkxjtBLOfHR/NrzyH3TIMRno
K4+xM1ywOg33rkQJf4i4JDdZhsEKJDXKa+Kjkk4O92g+CGChAOuT8k1veTidOmmK
irbjzG3FXXIcaFNb+pz/yPKvz9JnwNO3kP7vpNfFiSX2C8svMKGE02UdYE/YK8Cd
tPkCHAUvzSCc48Jky9FmGIslhw/APR2nNA4NW53dCYHqNcQOh2hZNVITgLM5aGXD
h73c8NSQCF10FEU1MkLKLwfDhYhiMa1x2QAhdW6DvXmcuG688NB0SGyxfbl3oVas
j3lWKBaJ58KceXJ/UxPJbf9XEz9bLZW+Geru/9LAFE3O1+A+XROtXQzmwEVp6IAu
NXwld7z/wRT7UCPqKItLtLDNnhqpyMIjP7iKbRT448A34LtMHDtyDgULHdajtGt/
qkHJ1x0lEz6x2E+1T47VqNfxjk7NsvGU2vgyX27D3zeq+u9BTsC2erWGUw7a18he
oiEu9KwNvc2d9z9qJvtKqJwfeNa+L0oZ6a2Og1zuIguNKp+YEuTS3Y+9x0avN7hn
FzhrG5yI85DZV2wFXUhG5ApkDyohR8D90p3I4YdlPzL1SS7WzPmJ+p4hKHva1tAu
2TQiDARFY667sqgdG1heZo8iZuHTseX9ubp5BpIBCN839kvgNYfEjetqi4cRjAIv
ucuyVlfL/xgGPJqPXpzF2YQdedDW7BRGodpRKCozoUEmAY+8VYcz8wJs+8WIluvy
fintBa8EofvybBW03XjzvumaefWvfl3rZXLgl7SsMSmNhDiTX4eRrGWQQsugF5mK
epOCazzra1ZsKZIxxP1S/IXOaBzVwaUIRT/GGUNuUZksnpXGHX6dTZBIqAxsCkpl
DUym9YuVFXvX+osM0vOo58h6uMKb3ysVTfqtXSc/Bv/RUYO8tcvS9vJuv35vo9gW
UxNq0DLkQkGApf207VNLet3Yv1fERpL6dp1q0/S6JSRIygORnc8epYpkYdDwQ/mE
nvqwzi94WtSCnCGvyrcmbO3gM7coYqpk3dCSsOWQ23aYqgifNW9DwmIU2OF+i6y8
+DeBmIKTBrifegZW5MS/Cl2i027raamHT98EDRh36SgyK5pj7jo/rIrs+CgdWDo4
9hZLOZpV8q0pSt7JeNGWW1IPaCeufS1j+uY3fzZEAiKP22AYw8A15OWysGuwoLAF
YqLiDhb/Ucsa24CeeXWqjhp9J84vWQ2HwODr2oxy2zmMqWeQ6JTVn49OZcrRJTVN
d/oadmnZvqeMqd0Vx72I9QLXnwSqC5Z/+SW0SRku20br7mco8fUtZDX4TABWkJSD
diwkF+kY+22NcPxOLG27AEHivzgisEvDezCI7VFaFzDzM0RLH9y7DzOI2NPsWj6i
vip7fS3mKcT9USYLrHBwnUU/73SSF2wKUlB6JJyaopqxqn3FR0oRPLkf1SxzN04E
6j5PrfdNViiH+wUMz9A3aujVOWgnmcvyX3jsgdEdnZIgpGHQreBDoewIyffWt6uA
lZDlSDDwS7cqxfNjVfTOCKOb/Tny38xyGySCjhgdTIiVJBAw6fOCNRWGw/dm0uUA
jcH3kZyMAHFnV8GOUrte0e6X65z7THkajRWt3JjY3LJo1NPgplQXXBZrKvLB1FA8
KzACOj1WieVNbJMwK4qSA6SydDQ0ucQRsUqezD2ZQkJYhHH9nYk0fJw9fSBZNRvz
2y0iPWECw51yZlzHKjW9iEpma3dGbX49qN3VfijwWZ3C7ZwYzqMBLAjuF+HL7sLT
j5du6u/pscBLHWsnqMzC5/vPeBTwa+staXO+TuauzRP1iOnZi35FBopHTHdBQCog
R0QtVoIegSG2Sboy8WmVaEoFndAelcNc4a8dABx8uuZROWAWQOKGtFRVeOPEo+Rc
jQCtzgh0+TTbX9F1kV1zGaV8p6gd9J88RuDvcD2QPj0GpWoMzz8FLezPg+ax9hOr
P2UITXilIbeX4CEG+iGkpRYH4Uohazz0pLO1ekfcsaOm1ZLcR/iFuKj4tqmzS+n4
ypsZli4ySmACcn8mpygPvM2f2cXHtSZfevW/mzcDQ8zexTkC9R743GLhzQ/aWzvl
rG1n5qjG7oGdXFo5OwXtqaWulRNUZZku0prrCu4Qv6ssfKoo+9lw22zPNOVa0X+V
MxokmGGCJwytAuKJ7hfzwlDPC3xx2fa2iWYXRMzBU6E8BaPCTkcq0ZjEHeaTJ9h/
j2AOEcoOTcoQ75UDySKwKqck7rtg4ktmPnll8a11YscoORFNT4nS8CHQ2gJrGwFQ
lcDeS9LIiOVK0ZOPI/FU+egVtrZFNc9ZJubzuNwWwD9XvdcS3auaOPn7Ch03VOhu
AasN3K9F7NGnvKO14dWIPOyUDnJt4dQVDMBil35VQpjDLIvFKXYOgXWzavMtpFJJ
bZov9Ju0nRPg7cTHAW7g77/M9yEvycOLR9wDI6DWXwgoj+Xba5Jq4qEJNTwTrlsc
AoeiHQ41XLbCPped3JzpXE78Kw5IqmNJsUVk6Sl1BgQL7GPEaZ26bFOWP1IrFvjg
RT1Kxz0eGZfMkFukzrE5gJyX6YP73HWew0GejNewTchYDeXoCs/O3yBYwiwchA9V
+GA6zzfDDis+LpJcpFJT9IyybB3WQUdcHMQaF/gcQZFZ46cXXNIF4svYqzzhwvTw
0RYqHA3oG+d7K0o9zad6F/eR0mIwDJEsRJJWg8S+EutDON0qKSNBH1o493CshRGq
nrMNRbGARJO3GNWTxHCxHLhVIczX14W0oKKfe4jgHlB8O2uV8cykMMKwu6TDbflf
xcnFVPmuMi/AFBRjHOMWRPJ7YZB8ntOJpV5rO6JFzl6EdQLyepyho9KzKbxZe9sk
cMav+i1M/xXRQhLq9eYMVsrbFKHvl6JnPA3Jkt7G7gyloVfoabqAXYWMfQxTsgvz
QBzb4HZcSdeOfXkeFkN+9fsxpjXlsCHaJUYUZj9UHM6EtO5gE61QyTj1D5aIk2gT
Md+JGX1lP6iA5mh0eYeuPT0owtWtffCkyHHs2mlsa8+XqAW46M329hHE3gtqbIGM
skd1r29JTi/niRjfHGpBGQNjPGt1As0Fy8Q7y9mDx88I/BNnyUZx7tMRV59Hop55
pVo0BR4jJ14yD1tzbuTKri6la1cjUBuWkOQYqnQSgAsWvU+nVi3dlu2ahPjPOMiY
Ml7OdC1fdDaewL9lM4hjGPzu+stCYJBnYdLMlKslA0uN8VqUFyD6qH3CerhT9FxO
uftWAagpItH9oPv/Psbcy6iT9/gULbQC0aq1TLA7e7kD2b/cME/9eZZKtJmJV4Rb
LlDW/Hf4iqPplP1tagceBw1vXLHgePbnlzTws8JWjDVV1U0JJb/wf6w5dTQnlfGE
5qPiqnpDuWppf2PmAjO0AdVnIWNrAmP/OUGf/VpgW309aUqN3GX36E9Bi/EFHt+0
9OKPK1nGqVEOYfx9oz+6pxh7b7bMAU50Ob7shBs7YKa2f85+NlD6Twf9d8dC0que
xVlKC5qcgcHFB8j8Oqr4EdI5BGQ7hE6SHmkPhJZhWuSYpoVvwPbMynSffoou7cBf
Dux82p2MzQUTliyRzgpBs4ZAJv2nx1ip327IOkZjxoMGGMLAh0Nvs1C4IE5XEgNH
mF0lynYdf9UV4yLPlgyy6m8kOgw3grbFzD095u65/pGnFhDADgEZOPDDE2LXy21D
SIMJJ8Y8elx9BmKpKSPR4oTAEEd9rqCsF4hRBHK301MFvwz/2ppGhB8qNxkTUZzF
6VxWy3xd7GSxX4HtKjf2HGMtONfxE8XSgTOrJIJEWylXPigZrbBxwKsST1pnTfdn
HNz2Vyt89bblsRsxEavkr9Tn3QOqm4R+qGKgegBTM8fh6PFw1DglmjyIM278/yia
4w5L4jmZRBJM/+4/4VZ/9dWfYMpLIjDA4BCGmse2LSu8Aq54W+vrmcRClFbfF1mi
JXQWoypvpel3wB8+yxKIzJfeNicoF8dMuI0ebA4+MaIOwxTeOj7T9a2KgGVLTWw8
+bKS60N2fHIZgiVLb9dX2/woRhsGsMLK7JyTJvfLW2pTtWo0WQhskgJx3TelNd95
0u5etYx207UTHLdUolCkMDjtyTD9QPzxMo8PxrqGQ+ibCm7TVC7Fi2FniTck6fqG
FExluOIQlN/N0SFCStGN6uR2YbsjkwS4yvxVSnY2Ax8jXSfqy5TJd4krkKVgQUvW
fYOaMtaUu6TU+C50wkt+3JIMWlr8Pe3PMydg/6Znusmp4eBskgK4uYcVqNA0ltDX
eTfNOTpf90I/97/JH4324E3JbFlawzLmdX7jqMBm62qV3eOm+P/mn8xyTLQdL2hi
5BFFi31nYoPealAeDzHUaPS9//YE8rvndQATK55PGo/MNJqUPg+ECoGKEjRfBpq2
/BjryHAwbCABy9ScDRFrzrPxzecXCwyNZKlmZaJCbTchfJFe+vmSAUMjRQXnAqxg
P1y0lBD+dn9nqXlnD6GpSs9flnna+tImFhFb5vuDKO1JFG998Xtx/6dh1p0l6R9t
QAfLAQxdLaTpsY+/M1Z6RVrmYf7L02fu+rwL5dv77pHv7+AZxLuMfmImNULYnHRN
69Im0b3et5dRhrj/fQEtXhgblMlCJiMn1qTIOF0dVH96aWCbkufVCn8FAXH/vjVL
v34xdG8VpaE8sw6uHORPVWO4kaaQf9cc7Hpmzf3orEgshEpIYT+6KPzRp+YOcBUX
Sdd9f9uljKEvHIjRE5ISPkXgbU6/RPWoXt/dbKcR7NVq7YqPe1CES0XM4vu2TYux
hw0sSu7D5f5+LtaCmiPXnVTBTwF8WIoUdWTgSPrvbzeAAWhm35YhKKzOwWYg7g/D
4ggXegMaJs/fbchnF3F4mDAXeLCQItZZFg7wQ0f08VGb+rwYwh4iJwX8sraf4j1I
eshiqx9OeY97p3RvvXNra0MgmbkkKoHtn8f4pBMZwyx1khEDyjXHpiyHKCqmfWAY
yXQ4wa2oajnafqUUwFkFFaxJcsf9vhp8r8+Ju5rE9uQ1MpW/SCN2ekA66oiJbTVm
mlTrfA0CYPXjscuTPZjQllYUQqrRxbO1HiqwxaCsFbCe9j9GCn2CRplDHuTyK0Dd
eusBhqAFUCjyS9hHn3THTVSBebyn6qW5ro2ryVCqsbfjuflDGRhcHUC9TDVQ4HZ3
y+E+8PIXygzbdRqwAxUvE156RqdLE2d4YC4up8dktq4XicdYifcFGIbqZ0DHmPC/
+qX8j28XEdJG7egSXyIkgJhwllbBpQXJdtGnMbzpDijxX0RTSpXonmUHsrU10+if
lOinmEdzHEADdzP/LnX66EH8TYwxj1NKQbiWAgqKRv798ni9KWOfmOWfV2tw1uKD
gOU0c0ju29+EOogv0Noxc9MqxWECZTaWemjo1Eizlq6unX5njnIfYXzMyu3bJgTR
s57tgNgCj/DrpnAljTRN0bPYhpU1+f1OEEQ6wyKkylfuFCHyEaj9pvu9Y+uSVz/4
KIsoP8MIDIEJuhL2I9/1mw9nO2POYzQq/wYz/KrYulKW0Ux9VAn0Fy4BGyqLUKuQ
d7C4Ywe+2BDL/mfO40vvFCQrPsQ+0a8XwJSINWJg3DzXAOxcVF86zepRjc73Te1q
qndb0Pgmdrs6an9TJ6WHPc5v8ynWSnTzQNUnK0kxHo3G7ojGj60zQti60ZsImLIJ
U82+WoTBIlxEN4SLUi8czkAnN4fH1+v/Ade8M793P4zSwvpDCzRU5LNtv49uTWOQ
ee2kNe+Oxu9+8c18V4Nc5mDnsoDvQVWy8zi5FO/oMkVu8a2En9XE2ROaoxTGZUme
x2uYtsgPeIV906bDDSHi23fmSXKr6+3Xd/QtF0lvRgT8XSq64OcI7na+KskUvpeO
XIYT4ewNjrraEkgidy9ySSmIFzmHqRumNoCPT9Buh4sTbHHbYzxeAax2GADhddgF
V+Sn637KY1AthF36JIZZd6K/OE+2X85NDDIL7CTbPAA8K8ukicqEWQp8a/paD5Zd
NVCMBNzpz9Bi2yHER06Zyzh05pqLbPHpP2s3E0A3geyi6HATpg93CwoA5kDfIEKY
Th04f78HFrRfYygZhn8XKLGlBVfCxU4bqpgLjUIzqJ2OdfPrIgwCaOzyZsCcKHH5
5h4gnRDZXw2I57q1I6TOoF9F9nvGce2viGuVHmqp1b8+eV/qqG9/FGy5UYBdC7I9
dV+4Bags4tEPbBmTGgJGQSJEVhSOWYS9Mncye/boNTg7IGJaJMKVcZRwRZgXr1P5
bb+BHnJRpeACQSuSeKRcl8bLYheMOFrh4BRg7B18kAHvZ/DL+I0j9BviZDqmwSao
k8YtGugWxVtf9EfWjLUI+gkDIzj+VpdNsN0eQ0FMLRGxosO9RBem3rdnWYFHzdSn
QcklK7/lsnGL/pe8n+afjWRm77tvFQL4d2FPom1JcoKn+R/0qpIHTewJI0GlaEde
wE2LONGEn9jbWOwFi0ykSYQPhwMGBbyfDkfxPy7hCgW3008Jh+Vka6HkZBf/kYAS
LwZOhHVaCdi5qXlDqYcgPWPHine/n699vcl/pJW/sTk/ewAGvlg01MU9861tcjr3
v0ms3HM4aGG5IyLu4CatMJGqGcba6E4dGFPpBF23RlRFT5ArFw4lpR4QYN7BqT8s
8QIuKGfZ3lkb8kUjtZFm5hjv/GphgFgedNNC/Q3VCfj0dTnKcTmBQ42b3wn1W0pS
BGz+V5/5y9iIV1xDblaQShbbnlkyQBRej+qye2k9cvphVwYgNKd7zZsPFJ12mOpr
yiRhz7Yqbd3q0SwcfA+MPCS1HrLJrn9KVNoUjMGOiaIBzSXYKt4Tvi88VwRRtwUb
4BnsG4RiDUsb/E3QzLHtJrFeuWgGljMnVOpTxksK4t/At4vbi5+AUXmQ5H+r+tbW
g+D1yFF+HSOoNoWcCvyVbCcTY775ThqxRhO8Ibtt4gBP616yAtQXd7rnYa/VwMEL
Y5YI5L+QfcvFUvw0xp+mzV8tlh9XVnq+7JRBgJeqY8CsrOatjfRRGpNSmWdHt82c
4ZztKIbxHlPFxizRF6JBY0J9NIldeP5Sx4dwQKgeiE0c5jEeBdxnEpDuZHHd2tnM
/IFi8nJFJxdOdwhV0oP3SkqAip2b4eeKlamk8rVqPUvZ8cTUlHEYEBXzAP+EZdLk
Tg/gNMWT1AtNbLKkrNeT9H2mMYtq7HuEjqr0l5GZC4EjUyM8TpDOEpJzmQC0ugFN
J2BF3SVipkOG6t57DPIBAyJM1CaxrhevOuUNJSfpXA8Cj4MkqVtFkMBU4spTecHD
Y0HL34mS2kn8+nuovOME8mXmRvMbkxGCO13e49PTTqeTQ9+9HqZo4fEp7nzzfS42
Bw+lDeXXrQTqUUcPZWGiJX0GdEmEMPVmiLuGvbIrRa8umfYmX/Yup9hEeSz/mu5C
I89/fwAVZ7eXOPOOXh2rl7WJGFXaOv5mcsAPsGv5GuIjQk//VChn/NISp22bp9ps
fRz4jdumB9u/xsiUNiB+ZJc5hWMCwqS8VoMoVnY9KGeFEnkzTinqe6IF4K5MveBY
SOFtboxztrwt0nlBiQpRaFOjee6SQHt+IcydTOtDz3KYjMSiz9ycvX/djb3SpofV
UsPUvkjf7XSIHoKemTgELHZVS0SxypGOlTu6tdvX2cI7lSJzs0NuanYkOa3me49E
V9GlpdnnoWsvFUg6Z1A10Uz1anRzEB3xlE2d9A13ztfg9UzH4Kn2Tgan5qM3WsoK
opXMcVlejnPmTpd2VjgitBFTaSx8I16pEikqCaYir0JJY1LBc89ozMCiT6e7WcJM
P1hxy4mynWw0PVhaPN+ZTeZ/kIfozjZGaDBcsSFZK72dwe27oSl+0hvzdRzWcYgR
27+uf+gEvpolJV9LauPb27qhvpuqtZRQtKc0HndKrICuICW8HpD05cpGyN8i1SMN
pEF5E53q77cBgaHhK+SXnAzVIqPwq73kg/lZDtx3yETV35UZVZW4ZB9pvLPML6ZS
JH6accIlTh8q+qNvEr/ZefCIBNItMvepU0CmcImRDUZxwW7kLhP9uaQ6UKGU3Kyb
gY8k9KY6nCxu5pb7IEsQoIvoXsoun9T0fpZzv9If4pIDjehrmao1CwoxPopI95NZ
xIDU8aFoGrdzzRTBQlFHJnKXfiHQdq11qfhnFrkGFuhhzgJB+oVX+A3OhTPk84xZ
rYr2FX8a4LTbBt2ln1X0LCX3vtEEk4HZoufGCwJ9+bOGTvwTzuDN4aBjvLaQmyhV
Iz90g+A/xaPkSoS8LvbgWjj1ihmDU9pbm/nHU1O4A1V0Ouu7B10LDY0d1nzz41jW
AIMnqREAKiZNNA4F6ALyLibVJve3sVju/378uYFl834f9X1R2dNhnUQgfyRMGvPt
uskggcvTXGirXfnPB72DSSN6RiyTmL6I7w+AIquA66QfvlJ+/PNEIxb1g6f8HG3Q
QsJYziElnWqjzXV3heVVlzZdrXKCfYSpnNqDTZu2A+GhizAMuoJTw4Gt/BGWjLam
r0qNz25OJDMysTW704eUVmn0AT/BBJy6zggyMjLYjfkOv6DC6bnyDP4NIBtgCKvx
RUCM1ZpAyLuIJ17CY9okCJ4KwWKFjAHbQVQkftjHETRWkKt1R8sSlXET/vR7jZFQ
joYn5oauHXe2njtU5Bq+F/QqdwGtq9SrU18bSUwX31EeujKmDRJdS/7w6iVgjaH7
HaAYe3yb9pEoPVxwpEqbmSDP6EIqIEL/Ikdd4jocJsa8mfpbLcLcfKYv4uMMZEu9
jtEG25S0WF4jUXuu2rJ7m+sGBynE+z/LqD5T7FE4bDQRUwImy6l0gCK3KWUJn2Ib
UWxPaep7mljYFzB4beC/3KdITWwnVp2asV+0N6hCATP7mmHox1vo5t0YIQ4UJJpA
g3uSArLXC2n+Pv+69854fADMKrSs+y3gpX6Umfz+QXRPFj7tDESqru1vU/Y+8xt5
+9xeOhd7U+2wcGL6BvTcA5F/yBja66BScyrySyPHRfTMElLFMTRB7ZPBhsgY11Dx
C4t+NvzVFK7PcGEKzwlNw/6sNlS501pWmAGAade8ylFfnxntonq6Be6DTMaYur8t
o3UyW1GMYVgM9fg8nq20dEium7B/Up3j4iPQxqDccf1w8CUCT4K/SSqP9WKr2hjH
tUZm7GMvFxBpd/3g11FvuxfB0X5WWhfy6TxLadnfhQhSSyoBHrbURg7bQyMlXyOo
0jvDyRN7HHmdSOwXCXwbIGLhBRGY7GIaC5NPdr1t4QMElXHhnNJ31F8kfWfbREnv
Z09qLUBFudTc/jbuGIt6kVwD8oADXB6Uymn3O8HCkQWmZ/ZfRakTelBB6t6sFdBC
gteyse+chtdZO/EkqyD9d6Yg7v5yxx814v80n5MJ0iB5Pxremd1viTZ0N1uWa0da
TA7hnWbcgW9jvcrFtRLxMDs7wUunmnnuvdNX1sOiWCm/J11ggH9DTuFBVwAr692P
dMJqqj8ATGs5FMmnBdpWhwUj8zfTh1NA/S6mxdLuVK0UqsJ8jSIQCr9ZRhob07Rc
Oyi0wcIEJ0cSYEP3tXHxjVOTYwfw7O4UqGH4OjZe733FjFyDTxO0U1b69uOk9EnO
ZS5TyQ7Ruj0Gs3xPlcPWqme2rkArnsRrpyuj/g4QHbdQltHEJXMEtkBmFSFo6wa1
BK3byAj/tjBAFKtjKWxkjk42+QPDnh6SCuvnthxLdaDCeC25Xw2d7E/iAgFaXN42
MhZtFx/IU/JmN657as2+a/BsZ1GEWLGe+dpbk+rJi24wY+PvRzVA5vfhouZPRuLk
hvi7nnV0MMluAWbmVwYy7RRP8/3BafFZRkO4nARL0OVaDFJg/NgEfvTslGamm5uq
hgDKm0+c5SW+N0NMQHlEr6j7JQ/eAnzhodLD9x8h9UFwwrPGlI6dpop4dnZaUu4x
m4WBQ191dDtnBGElP77DTK2IEnxG55XixY8boGMfW3byMTFF02XmkjrIgeafMK5D
6JVIu/ct7IN7ZJlZ+qhBdBkwO7spzj3scb2Y+rHg95Ul1RHHBAwNnCiAr+LlEsFO
onw1B2+w1m9aysVWPAZp1gU/dgC3x+ngA1XbPMrvbnizc7LhZmspahaMD5uY+EAT
44NJAEs1BD93G3Z4igj85sIa79iA3Qp6nNGh3oWFhSvWkphlJLZVj1vGx+7XGMWV
D7vOnRGF5yp1+RA86qTENxUFEbwEeCyJCGXnSBfZRQGsNLjGLMD65xfBorLCX1x/
pXZ/taXLR2sIjrXIvY/vmQH/T77P5gkLNLFMspG0N5qX2AD8YdvGueV89TBQZEgs
zLnvzxdTf6TzBIe85V+/ZGSUfuZLqUvuReANfdD2vOUKS/iYZJ65MiCvvkbCiG8h
z7mvAbOptiUcWaKGdz4JUl1SByv792yq/JFbGdlb+AZaFY4ODFzRccaJ8G2jhjTg
DwOiudmDs7Hy5s0qAAiIVTdrmDHnj5XhB5lCaB11G+v9rM821Q4wr/4Y9CSH1kpT
tiMWsK+Yl+5qmBa/mV0FhOc5M8YuZJv21InY9efBH5/ALOi0+yBp8JQ3weet3sMr
eyB7gpoj9xd2G14qFal9KgcZUXEc96mUEbPiDCN0zvcWCykM3ZOGIgZKY7n1yzxM
nDU4cKPWV447BY9RZU/K0Qr+2yBGtsIjPJBKo8JrhXGb/AGGT9L0+ZzZ5/u7cLSe
JPIsPfaFcF0cBz/ph1KV96GX4/FW6jtliIkEJyRiCpRtU8KcVBnWt8/01Ic6Z0Qd
TmRrB+yd+5SHyfhE7pzSBpRzEU27EA3mlziNfBgs6K7O9BwizpNbbab6arHUZh23
6o3KeGJiKRdF3+abPP4JZG5KbOG0dq+b9CqqqqvgoqiavnwGWyczBUQ2ygCjxkDh
MvRx++c2DMLby0bxzyYiiC0x6t8pIjgG/MjgCG8CIUEl/KOpvIrdo2FRSLJFAelF
zztMOkeBhjsDDLpGyRD7jjYRjFjaLpVVi3FeNlXejHZj99bU58rbP2KrCIig2gwE
uoyt5Ze5M+TLW2yJFJwX9zrHiIgNtlsOLuYahhpCKUP4QVgoYeSfXHJ/Ej6HYO5c
o+zji7CxHDwrOZBUkx8PFGqFaXEnTZpWGiLSkSNcZGR9s2+KCWKXQVrFYQfJC9Db
2+mu50Xd9hDxBCsFYmiwC5X0wZhVUzJZzvVpk53Fv6mcPnSrIUTVhoIVG0UivYhE
k09HPivsakYzhs/A4hwAwnQsq7njMk/mTvxNOyyoxHA87OeflotYP9Zm/mSc1wVJ
zLV3JU58lNVt7RlJNBwiTLaIA5R0xRM8EvbuYrQSjs11PWwnOOf3IjTDgFV6upf7
bF5aoqfbAwOyAIFwS6aXiZZws7nDoSBdxc6eFFgAqfw2AGcPr5bph9GL2DeprkDr
Uo5gfQwQSApxUk3quE7NdXM4onT8rmMzmC+AA9vPCvqMcU34gvjK72q0v2VQoa7f
a3VL+h76b6ZLZWmOn6Iaj50fcksmI273zNzBwrNA/ZV6wpcQ0VAqAzsvw9uYpMSf
5iniGsYtzr8zSkxvxAKVRqPylSL3Gnh6uLc4XhDlas4FaQqF8ihl8yFExc6wbLR0
7MNwK5Z9N6bXRLkeGmEwzG9UsG8LVdtHbpvPmHdYChuGQGkyDHSdBHw2JEooB1mZ
GUJIuG6btxu5sDlrgpSvT8783uuAZ959tDEx3e3H55MbOL85IMushzw8F9YzSt10
Kbuan5FOrkC26JlTd2+KT6W9ljttvfo3eZP6qvvq8VSKTVj1SMI+U98Hz9NC7STs
NNBCDKzpWsmliwPiN3zIq1ZxeDWZKi3NiHhVL6L7KbEfa4G6cUciznrSa0gVzdkB
X+O17p9u0cfQTYNBafr9YIPXp3SWIzwfOFNSEUaUUOmNkSVAvnZKLNYoMJev39/w
Bu7iVc+ry6VvsVCom3605iW5sxt9lYfev0BMKG+F0kskD7ehn/3jCEHHHl1kPx/p
UgHVOWzakwtBr7IGnB9PtH39jnt5Dn8k1/OSHEFu1k9gOCrTiXl9xxvnZfYvFcyn
OOxs5QgJ8rcyY1NBr8RTIlZIoVYrSEriaTUPxg1Cu52PYdmDNQnbA8J3d4zCPhiV
1zS0zYgpTGZ5spaxQFE8oGP7DZCjh/RU+qxLhf8meUKO4tX5+a23iNHgkgTvdcyg
kr8QHICy0IiZHOoJA7RLJXv0ktqfwEoMo4hzqF+6GfIJOOE1RpRNSCUpJszWi4Ks
x/oiw0JxDrUszEqKgZSXFtmNfOQrBV4+WG2ekkiO/XSt2j3OLUgUjbbIEHJg++DZ
X+0+xfvOOCVX86pN9D4GslvR24llvOlxoKIdl+FLwRsk2KZsheqNuKvXBmp5urzx
OjAm9nUol7T4QBAhfzpIbnnXd0tdGvHnxRRRSdL9wOu5tr4KrQLtwmTX5Ungx8xY
5QRoSgcgccqC5lCyV0DYTsm0xFrd5vVq6NiAQ268mRNVWU0ZJw1ZlQmthB/B1DPs
8UyKJo3CO74FPAnJhnoJJpiQon8HgZHlbyZ7HPKry/7Afq72TSCY1epX/jB7eqmx
pDB9YRaOGFo8K7lN7e9xbFhz98TKtcMqQxA6YkDOEpc8nSPZhZ+EMcAwbdMG+UWy
6WP0lgCbd+jQtq4mV5Jx14p2dk77hiPEkvWh/Ivs/HhmOS/2cJXSJje0CuNJuaVO
uuPey4mlVzhutNYdrieDLVNR/Fv0bP8R2WFGaGOICTiezvF0VHfe/h2yqQlswrZd
pijrJKX1BylAC5bPI+ZE3wHk3DzBiAk3NpgbXmyc3xeQxcE8GlfxOpJa5GOrRZEu
t8fQmg45lcQET7anztCxLTD0pP/qiYArGUK7LwJ1QmYbBzEhwanBw65+4u5bJb6o
yUvMoIPtm7z5OqTwNjeujKjG+Swk3XnDZafXvLr10UxPHdWpLh3eIBmVfy55GYpX
xbI7SoLU6t5hHymftUajVSTMnSYUsEK1AqsIBqmd2/7gGqlIplAEBvORj3qroRCp
dSXggIV53VLsfL8PMvfGt3bbCJj2Y9fFpLFXTpV0XUMpjohKIkA7GM8lAiSBvtsF
0Yjx7E+kvT0LgHrRuOtAYrhVH+kGKY2T6QH9nLoECYQAamQ69qnh09qP315RGljq
/jjuOH/jBJucQHIHv7a1PudTVLGABn8D7Bx3jtExqQaDsq3adVYlvvzNojJZw6NK
7vGiL5ABqirhTS1OlTvkPAvOMJSDTOOADZ/OIV8YsZXbJDaXhRNbZVxQ1NqYmKLH
Q7BwPcuLrHAw8dq1PeTJZJ9PlfeE1Qb+RVCd/PXeRj56rQ99Yy4ZYgMU8uFepA0/
Q3fGBclRLUQ6P2AjETLwf0CFlkJi+gqgRpgOzTm/iwZ8myq+aGBBS+MokgWRFKND
lo+89BGTHkN4B4VdZmjCT4iU4Rx7tsheXUz+Sphy8DgAx4nwGxBp+I+rju19Ylwa
O5wOe0W1aZnGc1esWNq1VZBlYdXeHzbAHGP0Kb4Jam9UeAvI2fVDcEB2ivsqHD8v
EmpJNzsyaIFo1TdDtEemeWAVVocRRB8LumahZCHEdzAlmWeTejIkoRknZ1eoHrXz
H9nJAxEM7ZhKARNL5XuLJB9NzwFZkLU57bkAuxbjU+fkU/8AeswT9DeYhiSwC07N
Z4MwGC6yGcaLci2wjej3QPZsE2vRfSDOTB0HPWFvv4U6mpEoJhk2Enqa3ak3xhoK
+M0OZxAqzyZICV/FxNUGDsXxrcbcQpthYQ7pyy5/WXXiOBvBW6lazObG1T2dmNA2
2kXrmo8AGz+vh9AgbTxkOmCGejRPbB8hAzagv253/QL+ir567aRMZrcUslxcgt3B
97w+FkZnSyQ/WvxYE2z3MCwEZfy1OIUuHmOFraV0m/cS7VgwLn3WGVspG8lcUeLo
mGVEd6qQg5ly4MNBw74FTAhw6QlJgUpagm9Gmd8K2yZWknBFAkMproiX9VvvOz/4
cMNSz0bIXTjMgSqYnhTCBW1Lk+9xUGJSoCWQ2qPAweepwrakjAM2CqHR7JVk9hJr
12p0TfnQKHkGWP4hbPsP7U0i+4hvc2RyWJEfwCQdzEXhPnze6wlu5WtQdP1BfDt5
L1AVbxUaBevXTkH4N/xvhityFgGl8yHQYX4gXeuM+yHm6PxZ4jQ0fhLRNVL+/30v
UafbRoO6J0Mhjb+xv589NtCtMq2/W9eHEImZP4pl/CbNYtCzpifzfbRsC+bF87XD
XYWECI5pPsdETZiS3S7MTmrNIvrJrpcm/kPXGvz0HHZPLXCdxtA7CFOdYMGB0k4q
28aWZY0DWi1/PTO3QsKjvtsZOOFcz+sXEHynX5ycPnifuFppGi4500mxtQwLBNeW
EwBL0yP3lApycKILJw40zGauJxL9NmBbgzMac35bEfl6dWjFX6tcDux8xep/GDNG
Q7f9Q/nWI8V12EVpplo8Xhfi9K+j4mTqesbCG9ZDGu/Y8QY+PR7juH/JcRz+HHx3
11N42/hD+dYtylU5zXyZMYttO16O1nOC6f38BeYXdf+KqC+gS9OHVA+B+wc8ZzMC
EUtWOL70vbZz5eGQV8Hk4WRankkyfGmTYEJ/Hkj/JJE98FRMr6L6mo7Q0Kvd8NIM
N9jISazIVspljdRbps7qc4nkwTLPG+6+0Xflfd1lmLOFUhk80wJ3kKvkAGT5O3Az
29LcgthcE1Si1HA1u5W39AynSAOy07R3Nx4TqrD5iZpiARRh5pu5gaoBmeZzTmrB
TR+M/yRtAb5OOcB8FO2GqLyD3Yuf513IJ6rFHHQdhP36kWv1Yr23MVIrzg+s5a5j
xHaneY0eckQfsGImdt2FbUaMTSlJynQ4JWrRL7uJ9xcaIU300ZosAP4UYu+wbkat
4r5rc2Adb6bCeckMmbU3cougdZQtDa2PUIIzeWt5ShrEZRZLxC/deWoqYtb2OymE
HcNKS5ZcBmfd2Htc8rQU+yXX7AXmykFVp6xM2s3nbZd3QYexMA2rgyHdxs7Yb9an
ZZgofTgEj6SyIQIQo7s+a6S6l9g0o4xn0NAJzeJMGXvTxVQYYSGOAIg9S4ATuTFT
dS4YlcgoWH1Sl0mU+frwmurNFAFP0ydXbk2kfUTqgYMYHLgaV8Jup6yk7/sVTz11
dFuOPXfJQA+qvSGwZcyp4B0UbXROGixoiOcercGQfr77zid95/YjlUSvIxIgPsu6
Oa0EfeBbOLCoS8/OFoJAjW1ixad7IzfIu1akq3ZRr8uYSO2z/cCiMniUK8hvhJ7l
UeO6NbbTABLKKITQWCH1jDaTx3g/O8jaT9NgvSb8aAzgMpsDlKVVsKTwxUthWFUM
qjbQHoSL9xpoJelWRhUBJa3+ZscFxznjYGa05uGCBkWezia8PXr1jTCkM0U77q/8
mzYdk3cY11PbYSs4L5CE2mk+m6+Lasj546+quoPVIi+OLlmFOGR2vkVNLVxBo9Kh
Hu+VitKFIdLj7GcZrRTg7xrr8MLMA53ENVRaaUtEHkRWNFSJdIRG9mNQBgCIUaBA
EnBfhS1ApXtmb7V7Synv47BkhL4iw/8Nvu4ILjsZWQGD9UOiYpHvUrnhtV03hi9C
iM+fs3kI8qmMcU/eFidrIy6VlnofbwMA3b4RssxRwKZ0jVJ7WDuMMS6vLjxFgzpu
PgxslzlbHV4aIvdRJd1GmN1ywSCU/p8xrhHuhzEBLETdr4laPGOhJ/8e8FaSekhx
+8tnxzLKdjMOpP7iwJuGgghMyGmUDq/C/Qy+JgDO6y/xgSquzPKjK8Ob1dmikZnh
G7U4VoFWvJy6/XfTofQ5SzQhr1ilVLLh9ksdeySREXnWPuC7NYBC2CE8IcYrmina
kmSHPT5jWFMq356xzBUFvTbsEC6gwYg/ambduU7jaC6LheWT6CN6lNNMoxD+FP/v
D7N5k76iMM9CwitaQkPl17SjCLxIRIfbjVAuJJzY8BkAOm7N5E1/b9QAdlDX5U39
HzTt3yGiHyEjHzNGZO4tyeQ9vHvdllsT15SDXVvO33BKJ5rhxnLdI0rYXeJvnmle
hbwaX1/CelZfy2v3Vp6qgyGC6oo3qzi5fw2lnCW92uolLuLpRsFasAgB5zL+T8RA
6ZDSowL8N4K3ouqjOmOUzW8hduVzuOiiTrypf4dSTemGPziGBtQRjKGmf5DdJClt
zTdr05Qv13DfwBh5d3yTmgBr91IYyvDSye8qEiVMvnlJV1tSrNhSJ4X6BPrtjzM9
vyiwepy/Vr2KfP6bSj/qY/7Cdp1+UKngjjxUtXMN0+S7LN6wyVJYvtb02HGW6fiW
RnRfXbvWBpEtzbQRch38CvkYihNi04crG1h5LeBKWm1VjOwaRvnxx3K9XwO7RWNy
IYrMQVaBpabgqCFtBc2W1VgWjuV/JH0rywNgBKkXKJJoL+DR3kB2puj45TTT0U+L
7lk4b91gHZMOL/B7K4UUNQWIsk8yB0wTmymqZu/6/oXL5mnxyvE9rp9F1oP4r7kW
VC23566KZN7tkRT0rvPJC7my4ciItPfo7eBB4MGL3tqCn2KY+z47rUAXAlke20PU
6q3WLJ8vj64YovHQIjE4byDzwhffdluHV9Z/evH0mLg2HzVPUmiMShnmjmo8n8BS
X/wraM/CJnKAjqdif8bfqmVuwfJW2r0eeC/dromAiAyrXdD/DEFk1gHD/kUmbCWK
0TaywDNX15afhgKA9tWUfqdwSep4RzwzrOr679+buCIECyLOQf+T3iCaqBeugMYL
1en+SbQ6DV6x8zXJb/WB+W8HLM6KXIjxcHWTpTy+PBHNpZMY0a46x1t3nTZeV3C3
Mbg5KBGSbCibBKajI/pYBsg4cATSLqDUA13gBAZBXGp+59JkBIoybGXYWvOcR626
JCYIeI1KD3xodwgmDtZRQT90wHdwbvh5SxDkdfk780y6OEBDat0+BPItATNBlwrs
eb2q5p6T2+jJ3eoIgyQRzSuDON1RPDth5lsrlLhLsqBi6dSHIOeferpxNUR5jMoB
1bRkB8Ak5EvDNkGyLb4jhs1ThIx4AwsJu9oqRTWCJzlvp7trYQfkLLJ25nPO7egn
Zs6zArrhp83Ii0M2zxbMFVZt2cfJsaJzbE7tgBRjp77/yGXo2Z02GY+MaQChd1CC
Kz9XNV3Bp785f5ZMYn0kX+AUj03KJT4+GFiZ4FC79DQO8PXMI95m5ZFxh/kIJHDs
M2irZ/dkKDKF0aPitYhoihh3Vj6fO85DiyYKFhZVV2nSTJiaODyBqbQ3fTAaTC/U
V0KCc8vQyKSsigqHCrtcLLrFt+CiZlo95ei6Ag7YQCBzjorne9DgHBBWAp5tz7BC
j8tWekBdIt+/tFqXZ8Q703yGYG8Bga4KEX58CpQAuXalgMFEN9KyeP6bP/5wpq8C
jLW889lpLTzytjXt5igM5Qz0Qri3HLB35902bdYcI1TZEHOiz24t6Kdw7uX2p1+4
o7X4UXeeJRircvO/ZP4Oex0XFsLP+AF36MZu988yAmf/wfBfvUpOFOVgdZ5mRB9p
dVJWiKTnc9eHW6uNQSv3Om/N/3ZmDYCg7T0i+aLNWcUL9uG1fVRQzuoV+GflQdOW
nYN9dh5mfk7gkcCH/CXKrwX1WJB7wZ2y5tkKnMjbq3UPPS1LiCIy5FCNzlbkWz4s
099MMY/7NVkjNka95V4LxO8GcMR+d7vpwXEFcOJABue7WfQuTmfcqhQ9OQYk/EqY
kXsU9sdzLCKyz5FWGegmzpMr0TOEuG+SXWKKO/S4RpwF4hlXKtadu558DT/Y4AMY
qL+8DCZDGNB/nmPd0k0YF4/YTNqx3Ia3OwvH7D9Xzi58cNqCzCGUQMGG5vyP4eQh
GUJ4/LS3IExBQ0RXuDofFxWGBo1e+Qll6CazM/+NnalySi0VuO3nQb+2DreXDxoT
CC+OeBfnGkTkavVl0WgKMNNoKVhcbZtE+Jmz7/38ne23icrCIguu3WK45vy6Q095
2NRtzWy7TE187FMb6wak2fZYEAxwi0sDj22++S98e8SIsl9uLFov2AW7UX2Ah37D
tlOC667E6GUJWEns9vOwCL2UN6cHj98L9bFfSLSA76frcv+NsYlrJskZ2D8OTM1c
siFaXWCEkDE/rWt5cgDI1abzPL8La7ZmSnr9DSTkVC28wZ+KOpGlEAG95+Hp4cTj
7GZ0RAvao0TMDgrzNlSlXKZ2puX3ebq9CHjnsWUp1j4ZfEaFTxD+7tqTZNdaejhR
tKcc8wadczjPfHuVMvAZxjjRC9nSn6FLsAGU67azyjYRwGOziXiA2jTRVzFyvh3+
mrGZdUEThKvegUP9uECb/lF4zkwkhjD/0lXT29bcZI5eUopnEs2FOyfq1c3dSm3V
2JCG7mmaqGzx4E+BNhV+sEVxOOCm7LZBZbbaRg05JtHFNwORikBo9i38VrLDgJAZ
YB6+LAgjXHhhmayk6sWdChwpR5rAxCLI508g6IpjOiQLPhx5+/CLjv4BseuaQKG3
yBxR+NV6GR16M8Vprrb6kaVsB0tr0fuRwa9bfC8zCNvxixb3zZBp51YOixLhMZaE
zSu+XblyJP6jOQWkjTpSXxWTqDFxjThXzVGwaUlivmKsY/B5e17wVLpbUBnyL+O5
hTxq483/4M8dbt80IVyFcAWQ9s2rSnQTlzv2SuAlVtmhbIFfHBTkoPOSP8GPA9mK
ECG7cvU+CSVt208b0ZVRKAGf6GUk4ix1NGzHZRVf/xu6F7dFyAyRaPNPmEf7WN28
PGIhbNUoAE1UfmiqUlqgklyHTui5xGeMrwD1YO0M0kHoC1rLh+JvXwyw8zGWMev0
YsqKRw1m13PF+QEomyGVuACAkZVbTQRPLPdRg/jJ9MGsp4RRseDoUBSLhmSlvWN5
GshmaviFbCA2schsNXZM5u+0T4G7dydW+ozNYZRcSCzcRMpp7c/p88zyMZJe/XwS
sAb+YIu7wEksWlQAxL+0/rAycJpKFXL93k6e39aYdpmJ2iZCihaBsn+GOdeyT+Rg
t+aWjWiVQeQtCt9YS5Zz6nyzGchcS/eRqIDT/W5vf5+wZQRqXLlVBqoeNgXSxTDa
LSnqVamfIECb2h0pslMNktAuDkrDNf1MjBxhcDDx7/9KH99lU+MrKmeUYLMH+AkV
kwWOZlsh+3+xH1PnJ8i90/CaqpaSXgA58b2vKh1dqNbUZ2pWv7pgl5QOVK7Fod5G
BGiA3DwaThCXFMKh+YUDq9+QrM7c2ZKj34ybAW+pf4nOXEmwW/7QNRi9xYk7Bcud
7Bh0+Lis0TlfapZv71FDABgWwmHggm0S+PmFCP5WeOayVzUYJ73nLyPMdVTWjHYV
lqqBT0ennXJemOOr9los1HEr6+p0M0MMljItm9VPRycdpQXVHUtkEIHkKOGM8iX/
xm4H1gestv5YCSw6wtW44QLP5SvuD2aK5qWNR9DFKcgJ7iNQ7zl31Rf+cpRrJnvP
/ZbVdSARt9VNRxu11dCONXVuD7SJm97BQ7lCp7i0T/TxRua9FCyiHeruVzPrPc3H
oRPw4gPHuahBvO0yluL1YhFhI52HMO1ZXF4ozvTBM7aexPn4thePFTlfOojWMxN4
tUlOKHMSxL+zUlsbVNBTsOdRyjbzzmirV8IcraalXRlm+/0dF4H+hg+GdnPwcngQ
PzxmfhOIQZmef9iMbnLQ+q4hZLtI/namXhUyMkjlvjm76AlM+KS+YTHzA9jHENw7
+FbBgTIV7YULJ/P45Rr4v/A0VEanBO6PjuhBkTaMENXa9tm+ehH1tq+bT/sNNMCP
wZOclcf/LYTTEfeYiSP4WvOwWk1PUqMmlWF/EjpyLmzezdnFDaVFPvgDd/6ID/0b
kNUhQ9iDAnXWOP63NnFbW9Dhb/IGc5trR86VRH71f52iaBObDEpO2dEp433RusY/
GtMXOwAtGOx08EPeB8cdu1IyHBPjDAIV+BkDD9Ega4sWtOLFuHan0Jqfk8n/lBac
jU+y2z8nwNS9SEnmWNnEDU4UgUGr+DkFzQ8FhLPPNeJsXAmR6UEnREOmsBQJmhDG
jFWK1S9+2nt3/vowc570MiocoHh+q2I62mvv5AZCNVUsFEjAPtKJRCSxz1lCWim9
dmKmvjxyYcrKr5A09WVi614cZ/CDXbyDLG0m5d+8Hqno1ZOJQsm9R6hETVzONkUz
uDKOCaN7jEjO6K4dqwtGMYQPIB9P/TvAOWAcX7z2VE9+R3b5TKI3SuWB2IQ8mhak
xQh5JnzzHkh+tpfAl69qOs/q7MZJUO40FV/I9SY6uIhxeKw8LgENo8hdkDMyU6ml
JX7WpX63A5BE+XgsHrLHZq3D5kJPzUcWlri4j1/V73XhAYzWhNoNzzs4/RJC5Hgu
71AK4m+246ZlvXm0/iig5SayAbXB5X8obt9Bq9TxxMYcJzT4H19XjB4AtkNJRTdL
BU1Bev4KBoDfsvZnTlMKvm/3bjvZ73tIXVpjiQJQrHxswLkSVWsHGH2R3IkEsLpC
6rW2Dxcy/ad2tioFPqmjBm6Ryt/rLnsrBXgg0jD6QyLl/P8q+1jB08ycZW2744Ql
xrRTR1CQQjlSxyNAhnuy7m61vZjNGANzWwS3DQE2VxCs4eG2qtml4sM9FxjR4VBn
iDVqyXkkzQMeyioqIvDRk/PVowd1XyRxPV++V5jlLNkadbtmoWIDS8y176Vj0x4+
fqJ/tPZO5Z8jgo9DfZJPwohBThE3y0ejEsBCqXRLE9g3wG7rgY7L3RE9nSvKn0vG
kZvZ7FDQhW6hXVZFC6zaemgfT4wwgmo5nFyXPd/rgxwY3eZqztpiAEgRhiVdhghR
GT5PzqcfanF6QCHAOVpwGD9wdo4tw2KyFrd4DiLGhtJKLXCkj4KP711OAkEKBfW/
o34XVM2f3Tz8Rl0v0k4k/tfEzObWSwqO78jU6GghstUDSpHgjPJTnhALQyCkXnVn
50x+jSjq09Cwr2bs+Zx9KFCtv+Hh2xatpOkmh48SHqSaRgqnNzB90qtu/fpI2Gla
k5yJmpcWYoWtgXQ8Ao7rnnrZ/8V3aUusF9W1bRrYTapV7OdekxR/0qtqZmMm0uv+
JaRNifn9lXBCP54DuA+Zhr2KRnkp5oUz6PfUx5/ktkWfNXoMweZZ7ngtenSCUF67
f1qMgbyP99btlFSKFJEo8njqUtq1L77WMpeBviYvnjAgkFsx/pNo29l7oUCrCl8o
7bI9BbuS5ozqaxEivB/FxO6d2NCuoCl7RJW5RuapsKoc2iNb11C/hAbv1BH61rnd
6nXkFd+U9f2WRmI1NnSj68qMPmbwJK1b4/udoxrMMe05AFSayL5vSPBVvEnvjZUC
T2Zv9uSBxvY9G9KellmuGa2PDK3nL65QZGiS46QZaXJbpDsU4JL8g3SeHAObBGKV
XRxm9Xh0Hfvlwv9OigSV1OaZ9oy2UsdQ8UqmuEc92OAd3Us39nBkITdTErV9CJtu
LI8SUDcM7uVNlMkK4nGPguSX6PXEHjqrWSjgjKJeKCRypoK+ro0uBMStIBLuCIko
n+O0vUdkOFAVoceRzutAHqOOoeEERhP4VOAhnhOOVW8VpTwUkhZ3diFDxDhU/BNc
LUO10CXx0SU7+DVhhmeohITKtkfAIy32vemS+dHuubhg59hnT3YdXQu++EL48Bg3
56j6J+uMgVetBk/DSbZOAApgmx0EYT9q7V25Gln/j/hAt5VLlC84hFETjweU8es0
Cl9x60inLMouXfKSKMoqJ7QkDN4Z8yD2hx48BeFD+I7VDmXiGLkZTMey0+yb4X8o
LURNi3QJbUG5Mfbt/ksyhWB89O347YeEsvBCA2Dhr7L6emjoJ1RrMl5I5hpM3xVW
Rk1PWZRZBjrlddu/vSDBUa4Feu6W3S2B377Goy7E3sij/l4ukefO+FhP3Uqfjwdk
Mv9e10zr9iA4BC0b5k72L6cz6bCTN7gSS796R6gRHz2KL95uRMmIL8vdGuqFEiUP
WudhmT5j4DjKNiDvJ1BT2TwrFzR9WfYYNGgkKb8i3vZJ0CajzssHWoUwnLmVbt5B
beeyCOoO5WlcgurC9/rNV7kWxjH0XsANXNbnMe8MQtHcdJcLbw56b5Uxjsm0PNn3
m2OTAaBi6tUl/kR9hme5z9Q9v86Qiq714aYn8neIcSoZz/SYQCAHQeW60VPlt6/C
DtUUUOzL4mF5xwCRVJh+/Ao3xTkuZF6oA7wpj/cebvOhQ8nfxDKVn8pDZwngyygm
DLBtAEYWzk7/I+V3KkqTriJ7RiU+0dfUbyDQ4Fso8cBMLTG7cuz1WfdnR77T1ocB
5X+jVk5pINMoRiuZs1TcqW6q8z65nsI9hwPaBchQeR3SCS5Wv8DnT7/iseiIHTit
chIGXhDJOBd9byQpYUShKZJ1yGxDq/4fDbvuDp54w1A8gsqeXQ0OwTI5Xei4dMHV
LE2kMvAwZk7QYAHs+LX91QN4JLxruDwgUkChzCXLVfAsY298FJNyCAtyqbQ//iy/
WNYhC3mno+81YlU3XII5yaTN4m9pSs6tmzFDIl2dcQZg02Rsoxg5EWBM5UXLihW5
/NpeyWj2wf+V4mKPxIBWuU8oNJe2EDY7uL4kAerkGPq+TmgkkbSdPiJTampuNbzT
W+kgG53XD5GPSWc7ErxT2R7JD7nWKrwkseBCJFZIXg9J6VQH2qp/ldJ7j2ziPtiJ
t5yxmMBq0UnFBYCtsjMUiJOht82uegX4AKHWwblkzA8LMw6HOFMzBylMLxRfL++L
4TndViXKtjZrk9yITnbwzKDAExYpn7fQCiOMtrv0HbdlCIpK4WhXxNIXKb4YbEDq
XbAZfJzcc4fUFTPlJoXJ5HfKtfBlBL2+Jdbg2mF/pBAss2imNIecll41QhdLKuvR
nJLOJCrZy2FC+U9aw8KbI/I33LKNyx020MtZa986h1jahkipqEZhOWUBxa6wa6Y7
IuqvGCCwRxoVdfEKphbOrTgUJjVA91nS9J045XZveahIQ0Eg1EJEUdo8OYqSpkVE
C+T6Nh9zApjjtLo5R2570Bebxx8xdvvRulNl9bvaBL3aEZZFsdiHW2mIK1PImlOr
RFw9yCmQLqINYAWYW0Rn/kfKZAYTwvXZ7EYdtcQy3ZK/X4gMcCW5f2EfAXzUXQen
Cyw1mZgg7MPyVVNaNvJr4um/w4XjOKKypJtUNkNDJFnwdj6o4tLwku5IU9pj0H4D
+15U2XAau+neKzQql7fo650rtBn/kSUpU8DF839qRhglXLJFMWy6YvpRyJxn8d4e
eLwO6iev1OpM7Jkyt3482mSm8ZBo2E9AxcwSLKVSNQFoH8HVRquoRx66nlh5/9hb
ysYQoOokhohrTdJcUZJHAABTYaLTz/wcz9Aijoup/nX4GuNt1YqYSvFkD6gJ5Q+a
eTAlD/GZNNmnMs9ruieFPEtkI/fXHSMmueK/R/6ZIDM6qNpOKe2GoU4RdN/Dkcpl
3TTZr/ja+sbvMD1rhQiMn25IpqzscfB9iiMgVrfqcg5y215Uv7krCupfIwUh3QbX
X1S5n2Filv6VgU8eImfhcQiRZ7NqCNzEb0tmEoh1LD/eyHrMYHkJRTegH/l5x99z
/kpcSwBisrsb3iU4JPqfTSKA6qgpxEoezfHVQUewip1AQPupGRsw0ip7iL+Rmj99
wwdM/08SK1CTt5uxOYZdKGQKkGiF3VxqV4E94H6qHkWYbz7BZtGQScgg8Z51NDDS
aonToIO0aL29U5DfHtpsJFuhAg/VefSb8DoYWxmLPjkpKZhVmjWn1ubgW760C11i
beQACOs+p2MwrTblxjNB6QSu5LurXXI/m2lBVJy1EXOuCvrtVikIbr8qA3+HuhXW
Z1cdb2EAPbtpVsvkHvGSoyEUMKeWbqRvUkL/15iGjnkfzl5+PJ78qRQ0wv1KxqSf
4fC3wX+h1s36e2hUobJif4lwjEvpWe1jjqUkxXWWznp4E98lenFk8VdQnyaOVLqY
fTSWS6bWZUEcReoE4dl+K1dOecdbrWr++Yhid5xBUzyjwGz9W5RzcW2lL6bh++/I
O1pRO3Ypo90yZL/br+0JbefX5DZ3aDbk//sPXD0iku2SJefRl5jJTGyi9DSaWOwb
dYowuiyG1a6phdJ3fB3qKYZ48Dn9BTyI68QO3tTzFm67aUTUa2Mzd6Q+oTHquwlI
aIqvPCPK4FkS84NOiStGqfKQTkH/M9kOu3MOPLZ3cHeWQztlI+ZeKV0iyHuqi+ER
U3rPpw3xx0/LLuNlEy0c3O/j1L45n0QRk6ZsQdYEuDjLtG7cSl3I3XUTMdE86ZBE
yWmwi8NZDf2byUPQQ0K8aFgJ8YjAggcskjn/DqCs6TEj2eEtxyyZ5M5tJ7Y/VP32
Ih3demwxt8ZzF7HMw+dHzow2g0CjJjGy3UMZTNTrnN9oZGR236rQA2Rbe0qhBqpW
mvn1Wy84Uy5qMvJTPS0LC0WoKezJ/m5Z3zoz26KmGOsMZkI8Re2nx95jngjbtqko
MlAF4aONL8nvt2SnVtQh10WaDbvWLHGJYz1nHUm8hzf+p5CKi2iu1KokoLUW2JLL
G1Y9JyUByV5Q5HAlx1gCmbdjKISLI5ixbfFXr3HE9Vr4c2tbAC0fPcrjCzEhIYTX
WrTBQd3QuSiB7JoOh24+Qm7KEqyxqcXz23UcoeFh039kD43rm7fqv4WXde2L+qle
/A9alSbak/RVOUPk0Z9VUYT8LZ2V31USheDr/PZcYr0jGu67AKCqVx+73+nE1gP4
C4p87aeEp4LdYrzoeMICsYEGqqClM2iDj4r2MnmA4UGfcFBwHCXA8XONX8A5uJCZ
AiPyb7t6YSgaUYIAK5j/e907NWGhOV/o09iOq7+OAPlWkphO3Av95DNF76QQyb2N
qvmbfj/C4bHpLdboz+3Q9s3Qk59rxLi7/dMxOHwn/Ge/gSKoawuI7Tn93G12L5WG
6oGBVf8h5EmM9cd+ZY+jMPmtrqhH7m+94IFTZO4U2qdNLo8flcU9svIrLsbpiv7T
pUq/LMhKtcA/y1hu7zs9+Z4vqEDU3UHC1ZUS9uqeVKgIIl/7fiKd0juZT4i6E3/3
8sCVyCvL+ZqE+ZJ+hX8DyXANtNsrMPss3s5rC14DxYxKxQQ+Qc16Bria/ieXR7Sz
yTgCSaNsgg8yrl43LlOVGbnNnmaXBLGS5JRPZsW7DeykEYDEORmfWmYosERGMIXX
ln1jpwE2EUDVNqQt/e0koOPDFA5F7NQjtqBm5pxIE0AWM8fmeLYLC9HPD0g28ay3
iJATPl+B5Vp3ZSRgzgjakzC+mUzucAw4FrrM3a0/cWnXn2TsRtuo512sxMIzXtrH
LskTOQG8qyQIOqyzqkRHs2q3V4J1u1zrFf+TKN5DKR0vVqkHysZ2gNRtrPL4Og2W
oLevuqf0Apo7fUjjUXRK4u8YWQwmNS0+3d3INzrDmab8GXv23PPIqJG/lBMoZVIu
m4DbJHuSRvOZJ/9AI6+iLOSr7RGm7pOt2iS6KF/fLiTMCXc3taQM3TQtMmlgq7EV
/q/Q11I+Sfxwjp96Rx3HvIXyPfu7pJgI5iglVHPYhwwwT4EPieafsW03HaF9pXQT
hsaOtEvsYCmmGYfSWNI21BxcV01F2p61fKmBDPTs6/rOsMyc/zqLilVzMP6G8fE5
AV/zCY/TAuXHFujgI9k+EPLLt4wRMsiGTPDc+UbLNtxx/IXBOOBqjsnbyHimyfZK
EftudEx5Kl7q+cLQeLwCcOuoAiRwUJG+O4HVdEosOVD8GS54TDJb58yaiZrluq6d
fEJzqU+w2X+laLwojVNWFrLMIyNPCs/q7E10rnn/RjkRSATJ4OKpORfjHrldOGbu
f8nV71tBt/yVQ64lecxYelytB4yV3+EeOqf8IumqkxrP53PGQ5j7/hapR2rE9Evp
ZQ2RMcrAuRSuqX5khe/SW7AHE/YLMe8Xw1YkmbBeSLjeCSZ0RxLAjac1HFCva5oS
TG+3/yCXWM0401fQje2x6hzbY4WaQLzypp6K/SsptsfeBau9a0xEcBM06VT2zryR
EfertoE268Ek8qoqcDvGqV1olQ7UE761oj8D3FU6vIdjfLr2KbEXm41QUll+yyHb
dLP4vaRw/yzAYb5TNCweUZD0PmbmiLcfUFPLYF5iIJFUnXUl/x4GljQ8lJ0LiGqw
R9h+FlqMzshrtR3TeOwon5PPgF2/VUX76Lk1x9kRxermw/VnUNbFHrBQlMNQOtFE
qT2Zfrq4G74HNRmHsbFzBiTeb1UllvF0tjsLghko7n9I9xmGuQssWHtlRrgmF8bs
kSxhBygoh6kRtuNL42NivHPhqps5+0ZMsf6x5JbJomDZkedGIp9SW8i6un8Cel2f
oO7HKnULPCzKZpDgX86Y5oMiQJYCH1RfR4Qh8LQ95CxA9JBlAGGXE/hIH0frYsSk
vvtYMvPbsQmASCaopuCAaIKypzq+y6NNSC1G3q4q1rO5hfMGdJhPmfiAIihtYELr
iNQ6mZNT/nvwybF5Lt43FL8dhGp58imc7992ChOZKN5b8w3fsLQ3sDa+24P+CjqL
k4HEpaRObfQxINWVpl78KKZ30r6f7686M79AdwnvAeHCZuJ6htzIcy/0nliafMFN
GMTGHx9kaC5DcHTucoq7CLIXHoT3mX9cmV6OcKlOmCbtbQA9dgSfaXKC++nvdZMX
f1XdrQ4RKtacodm3k2KvbXAxruT15J1v/VHYEvy4ITOKXaoMJpVyQwRkWhbDbq8H
P0hqYKjaH+gylrIrnzjA0YPHt8l5590/5b+KyAaHUiu19OYv8I/u9X2+sDrTc+rZ
5pkbQYxZ8dBDOjkvkPExXVxoz8avVNIAEqaXxw/8FYi2XeMs+R4b5RoVEDFgPlK+
XU5/MFNnYJFKDlBpGPByCMsGELj7HzPyt3auPYrljEPw7KFCHrYR0YGAj2mbVGu+
EiydGUTNH9nTtfntQY4wNqjXAk3TICqsRsfZMsqTExWuIbbBzxRyOU9STS5E+5yj
6LJ7VOVwFzjApez3OiQwKrWM/JJJETUOaVbvv3zlNU/UysGr/4H8l/iufwpL5dUV
JPWPB/EXnFUo5T60N89gJpt8Kbne/UUewC/EggE3rgiBYv5XVj3xxtCNe15Erxd2
vQT7A9EOZ1HuUAMF22rcoSpm18PSEwWiDZXBWhkqvDhD0d2/Pugkyt+iP6kV9HlV
tDwDh8ksm8i6aSm16ecGiR1OyUxX4YCkPw73qvk7lw99FEuuQ9vLNBq51Oa88z4k
VfD1uC7Gyse/dSI2d2fQIzJTb4/fzuyuZRMZ9Qp5j8rlSQmwz1At/Prxe1pIhj/w
q18kxyaLYozjgntbWcC7vgrCJc4nwtFQuAGYmfJx59mkXDd2OuNCAYSE8YmwHxFX
tZmdwwl0M/uJoBuXSUUnanS6H7WZWyJ+vzlu25E5y5Wae7cdAMoak5VWVCT4/N09
mTtQ3NBQU69xoC1jHIuNm7w7Fzz7ARBDHH2/wR/Hdm/3pK1nKtHxG2IFphyFygt7
cI2JeZ+AjopsC+U+GCblUW+nxtAYFysPVM0YzJ2/fx6i2nLIslcjfs+Lpc1W7paP
YdTtvQX26rCZFT2wUcLiWdF6TB86Q6sHbyuUdTaGJ1PNQ1LX+CWr+Z3icLfnitmr
cJWm4ZuvDXEi4vqN3jimAg6Aliq4GV0zVJcLHVhhBlEo6vjPnBtLinuW09oZMHba
HFBwrTe49tQNeAiRFW1IMQNE/pMi8f5y03MN9VHblbJRESoS3QtW41j9iCzo0J6/
YmRc616BhiK6C9U+HWoFnvDBAvD6X2oSpiIcaZUhOUkgbOj1CNcax13gcnweGHif
gA4MvW8JYHMpiCvVsxpJVMIx0L8H73w8/WcHSwzQD2kchwK5SaoVmadbtG0+lTHl
dtkOIX3mBbidPGZt3uOMCnIYLi1HrlHoS/J7aTxxdClDVJWV5ZWHN7v88u+x9jfF
Jh6LDf1vM9zdZQhdKdl9W6nEYj6tp5fH/serDv3ZcSy4NYC1YzwwYeJPR4rgSLXM
oYJp6dAf7Db4A72LMGaFCeWv0ji9I1lhnb/cyUHMxtmRLIOIoF8AD0+1EMV3tKJn
cz902xKoSR5UugHRdPvTdBWVLKWgs+n45fMVx0wZFJ4G3EqVcL/LLANu/gqiHes6
uMulhPze94/VdAk0I5vETEi1P9EklW/55CXUfEaSvHAKvwRTd4UsGTeu6m+kpVGv
kVppGccqiaOW+XHdPLiFtfLjfi8WdYALUR12sZCAva/HvX3fZfM69kXaxJPBlMCt
/PC5NDfTJtTaKgyef1M0AL5gszsedufuIDwvyCtAb/naZ5p7pQ8riu8YFJTGu0rI
g0qXN3LBGIrV0kGF3I+ijVEpvk/LIIchVh+NRXevPG9Wtcmv9Yb/skobrC9xVbcS
mJgsa75nJ3gGcdvHTsn6X9Bc8wJ4iAsi6EH0VvDxDTJQmZwhFxQKSjo3KmWFOOSM
/heFNbHf3LXe5/N/9y+8wFcYahf60s66JbkcL49XFtMZ6PRP7E4i2pPvoVkVhETm
0F3DIcK33/2OUPFNUNx3e5XfpEkU56mnstM+ihEc8RAUeMZEt/Pqi8rIQkbMO0hj
087ACE77uZUCvlpWuewE0LTV8MiPJDjzUR8UBNkjp29bOy4GAdbyeW31Kru6bmae
xp7QBr4QQDrJ5suH3jBnAt2SL7UESYHJozNZ4kcI4Ng2zM7jOCIQx4x/9MR+C7v7
cj6rF0M3cPLFRMI+FuxM+Jq2kwpgPd1jxQh40dZNj5QEZjt0dC5Qin+xDjF3A2JZ
P1aoF2S9Jdc5uyOAuZRW7QssXtevxw5gZNYR94feYed/YQM2Gbl14/eak/lubc75
0tLcR4hcERUW1YjNEapVA8dQVJE/YTnHcnoSeYOVbsV7odcpDosSdeyO/UMBl/AD
8U8YRpAwixtqLuSKVhhX865o5kfxk/MPcQQTqPKMQvwhf+yKRCX5F7pBARTRC54h
RsSZjaAxQj4Oje+ML0LEguTy3vhmDE0PkxBjOODZ931m3zXLsSH/m7fSd+dCAW5A
2mvQYoSHcx3XPHUuBss2zex4nujS1M8rn2+wEjNN5jKa+OO42f7XiWii9PAlDnpc
CVa2YRzQ4//1GK8/XISLtBYKqw5Td7lp/cZb1cp6jMdC6PF4TnIzE+iy7XSvBMUT
hnua9fGZkWdNqbewl3UqDtiFOg3XAlxB/TpyZ0iMbPf+mHQZ04Ka14igQrgCf6QJ
HrZ+XN/mFJjXExyQOhHMQ3Gb6tonKuLoX7Dq422rdYG4fS1FSpfj+p+o7wvR9sid
czKW793GZrEi401W7bKUPlhp3SzXA9GL4JaOA0GUw2qs+440VR2e20cyLF8UqEav
iKNpfoumE0UNbpKzrHpGcjUWFhwZg6lbczzdfKYFN+HndpXl+q4MCkPdS1LnbxLs
gabBHdnUReC26a4Ys0wDtNxX1ug9cMUARSpYcYTYyr9mu5LW/BXD0dbHIw96zxQH
6EUjfa0WAWQkYWS2diSQ6/f8H8to7ZTf6l5/nuOw4a8YTgimCnc9Rwi5hZsfJhxj
sbOSUU8YheV2tPk0Z+nDpbTM30Nur032J2qszEQrYjVSt9JFCBqYw0/rYY4eH1iU
IVbYF2RQ9xeVpx3ICe2XJqOd9m2KfOJwrJ8GGWMB2KQXqwul27ldknfPjsW2ZrwT
RD+YzH+ZqwqF9ggdXDetitUKb4txPUYPue+9jM7x0d6OaNVvLMtBSerN50JBrqkX
9nd227PMipnQi4pkNjEsv4VsoDgunZP4b2//y+iWVa/HNpZU0v1xG8YGRPAni8b2
ydKn2ppkcP+mFDbwZVbyz72bSbcxl0L+CU212CkDHkEAnLKalS1mQpzFjEVjo7r3
VhBjoJveWRb4qY5BOvg94cG0I26eD8ZnCe8R3HlyHNRi0mflGqBu8l2BY7PcsqvG
krqasEWnWPDusUP6V/Zfm8Is6Px4e7P7bTrwf2nhhMkhpQaR8B1n9/mWoMRMIKrG
PuVCzgQDrVDEKbmZVN36Y4fOBL8+xl+E1CpGrt/iFtW3s/1pyYrML2kdjKeYK/er
BqRWUbe6J2T5vEB6yv788IA59KvOE7DW1z5vGz/xRDdkrYaY63oHLO8MCR8tYtcI
CaJPMcO32SWcJPfHvvcsXwe4oh4Ko5G5sTdOoCs3COTE4/N1xyBt+5kVSc7KqAKS
GU4vDC9fKo3qRGRdUYIrsQj/84rfxSfaGLYZ/hkkT+FPHkfgwrC/aU3TtaJYx819
RYxXkShnAR8EV7R8dubtyHozsutD3c+U3ludVpl9ngvQ03Fr5OEKXgiRUuabNFVX
fCdcLFS2dqv+wZJfyeTuD83sMmlAV0WV8UOsPe/m8FX3dFZuWVou2MUdA+yPUxIo
VxpmeL+iN2B6k18hFEgjg1AqVQ0d9/5vko7i8kQCu0zxN4R4lJQV5isaoWQPD9lm
T6Qk4cjjOWJk41oEeXSoUKpR4lsyPAKY1n2uDctNOxgSrTNmZxGT2KyGnuNpG+AU
OAt6rEYoJsW1ayq5jJamxA54WYEgAc4FTikX5F4bPyKWLLcD3uKMIHZVVjhsY7VL
Wm/wq+KcW91vPNcNuSNGmvxWouInR82Hn/PSJNTyp1wmhPH1/+G48+WDxUgpnWun
SKxNJjP91Nni8ovyTFjOTvHGbQZsPrjNCmkj0mGftpidtmz5u+btRLdkFumPDOEK
02RuK7KpT2sO2mVJolUH2mMA2iJ0U0sNY2bShkpsjloWilHhGEWsp8ZtX1yK/nnl
6OM0mPfgFYZ/RV54WwY7wOh4vetGt6/j+s0PREnfNqPcuM+OTvuYdpbsDlZym+Wa
2dCAblZchKT4yKZ2QLroGWvngaP5AMu+vhr5f9xgBNME2YAzygSl/824mFajzwaU
GtpvGJuLdcE9u8texunytRlItbEKPhC6TQI3YwOMMHCx1FMrgiGnPWT1GDUVRn7u
Mr5n9afd8b6TXg1YM8AdcP1rC4w87Tc1ZZJW1k4LipZsDJMiFCS3oDxzB7pEbQQO
o6fwhR3PYIY9UzisgTzgtexa4YgTtZzH0udGoC5ITdITkFmPzjXvcDskeVN8k0Ds
NIyJZGPZga0IGAy4PVssorDH7Db0BaFruhWcFxZGKwC3mAahlNvJzwsML76BOmnC
lpRye88TuOOb9GMIqP9oMpUbQHzNv6bZFgOdX2Ag/P6d3T0AE3PWT4EgxiL/WA3u
fiWV997Uh/Plroe5yn8n+b2HkbvNi10anQ3xdF+4QSasPGC+vpBrtjkarsuPPqvC
HI6VPoS8Pw+ttHCQZnr/F0tVvHI6AskFZaIr+wIKouKGmAwcPu6nqjr2xeX15J4u
7uGIWn68ZBC+pLlbG/J/dFJHZwE1ZTaw/cAEM9ubhmQ3/kVhnUVGjk8NVphTWF51
Pb7QXKQNbJQ1EPucVQ42452GomPIrTD3xgXZSt9BKfSQH0iw+m6zqT5gSOMsQMfa
1BkZH25pnUcNleD96DdIojbJGqb6pNH6Y5YoON8jC7DQkwRKZnCsYInmFkaxgXMX
EK3h8TRqGSeExGo5d+3YohKpAX4eiAfJ2cNc6yYgxwWyuweCm4bI23DReePo7znG
W/vfKgBgf6t50HqmRdiIWMUt5FJUweqjadmf1kr4iqZGl/mLZV75V88ksruIqfVY
JjIlAJtdpWfOC04V9QIJKhjcLaCJYNgTE8f1Avl2D+VaLXThyi8VcKBlDbenr+GD
yPk2h1Z6r5a/YXvvsQGSim+aQfaHobRA45Up+jnfvv/w5A7oSvY2fwfosAVXZJp4
0JNsU3AYdspuNRceF/RIKTmluEeXXqzquLlcjnNhMmTW6MzG974jQ63ejTWXLM4X
wx9MizdL8CcFLQjKPbxEk8tmTELXL/FQdq4xvnrL776HC7LLOdyz9XDYo0HJDOMf
mgs4tUG6uJFCAOKDzUZbKrog0pskND81pb+EQzcXDoKrXV1QsFNBX1wc8oNRfKS1
K3fIW2CrGPgi8QcK48oOhZWHxOd3s+J+ocLFmhzUzidxKUhFWRfjCjZsGzQg/Gxx
MlAL4qyaggfuqp+NwCV6a8cDFfaZBjLlVxzHHGA+EN6kY9nxLMotZXgNQxz7M6G0
xS4A+3Ax3RRaXNCMGWLfdFDFItpNFZnxH79CFZDnzTrzx6WdHIq5TFbSihUXcK+p
Ais+ethg+VuhIJbkl4eZsrZxukAZYo2ocoxrLT9YO8nAq2sWR9p6hf/NYvbhuEim
T+Yw7HlfHcTfCB3VOAR0fxajA4ZwDK6Bsej6Bq+5HKm3kyTTGoycgtDF3VQh0A4O
6wEgrt+3sV3TRDGeQQpCU1SKbJnwgfigM4KwbTudOWXK/LfNpu/RVkLM9ByKCDOk
5a1EWOB4HNbybz7Q593IQmOkrDbRIl9cRNjnS4z2OW9Zs5jcOVGWBRVjNgog7ii5
+SVrKWreTxSWpjKvDCyLKhZVoQ4nn/SEkd8Pr6YwITu1ITrP10T6Aus/8X5XshWJ
kDoUYC+jApgCJudMZmb+Locs0AMVIkHJ9iiZspwvKjXh7QHbd5to4n25nwPzXw4p
hjVMKcKrKLNi71FjpK1EywQ1aiw9TRzhQ1+CdJmrSCMimlWdDkYwDkhWtyqsSEH4
MBJKTmIwMsSi0RkMr05CL6LNj/HICWWBoZcf402ao2lGHMd/XIf09dGsr8r7nleb
FPeGtip9WiVJWT4aTRNZzow3IHIgl1RWuESwUN2um2k69DQQACugPxGC+YgM/xHC
dQWaelFEmUQN87ynySZprDHNiC3mFlEzspiqwm+KUUPJE/4UvoPVGtnIqeESEsD+
Os/JF8FCPLj0PhfrXSWrBa3Bdb5tS/h0pajBav0zPcpv7H3EAYNqKT4utcbTBrlI
+tCIZ2mWjdZrBYu+oA589qm5db3B72XFJYJxrM+RADCTautfVGyHQwnlmmUI3Pf3
g7DrGioVDbbSDWq9LsdtzWxvsbpZOUIQq33gKwr7VuJDN0A2s8JUAWY33ibQsTS/
uxas4iKnXrAJah5QPcA35lDaDMutAibFRgLUsHD4IuGWmP6R39KoZswuMdioeiIN
XfeWg/POtGIg0vDYpxYN4y+QKEyVYgIhGJdp3vXA296SYnOPRjraVnrt7io7FPus
BcV9DdPMqAfEoxFZBGe+2MYuhXWlOinOkNZWCJhYcMKr2+k1lUbPLtiVZ9HBuHNK
Pp3mAbc8wRQf6EwutspSW9Dshe9DtLGhdl5H/w1l9qmEUk2sPYYWxSVFPH+CW7yx
bqoDqoJUxD+iwN6RrIUuBLuq4PDtd87rdbhSp9lzD4znkerLRCXObUr+f4bioTID
pq4KytAP1eMQcCtCyR9Tdi+TugaRVb7Ae9QW0jolzyDZ3vRieiTNsvshWrvA2M8p
3BR5YPaeH/25Ubey7vRXJkJmFMNqHXAldkEiu12BCOkI/F9vwx7einEh+Xwc8I9F
4/EEfjFZ1lyo62QGdePmh1w+V0D/M2R923TBlXqeY3RauVWxElXXgY3rf1wie6ka
Jv+/kSz0DftjcUmeLCweUq6D0EdBDOE4PtcrsHFSbkCUvK0g155lvgrgV97FuW+5
uKqMbrA/RHrsIQdqHaFUQEeepajJMwhbfI01eMhT/GI50Hv5LcI4aL+qnsHfgP5W
GL3xGgObfTv0XOHgVXFwbbjkgvtiwQeO6tRNvbxELP4HUq3LzqNgJsos1w+vZqif
m+8vf8cm3+ANCoDW94vRdJeB/opkNCgcg805sH6GhBYL9gaGO0/Trrius4xYFgFP
V1PRiwMlmvlHhYvhrIpega6p34k8W4bF87OVwedai07DMN7AQxlf13kfctcCIX87
Z9OWMD+dtN9YhkQNE/yEAW+B5GSZE09KEByQJ5yuZOX+HOlCrAU9HlMPuAiSta7U
SQ7yX27wJK4kEdgQEmI9S3k1tI4ayKIGpCQfZOrLXg+gmzXU2RoyMTMoytrcjiPZ
FnUHOQps6HNBKPbFbNufZu3A+clvY6KMuLccBE/TpyHhBz3FlNNco0nkyE1MmYnh
iZAJc/+H98d/Xy4oYf+oBqiQ2tlp9RHPWXVlkHauZ/QanMreNgL464Bjv+d1UqHY
CJgI2uJfETpT6s2OGctApI6Q/KDTp8A9PKHZ/DmA3MzmEPvsOlftBC8WN5s56RlJ
RCFo2DydeEHrgcA/5ZUjHRfZbc7Gi27iXgOsrlpXjQPsCcJwiYAzZHqSv/St5M0+
sRj1q7GPepHMpMNT58upMuLQM9ASdCtszKUcvX+gZts/8w9NISY6Hb+9DeUwimKU
SsPJ8naMBMrI0OLtPHXyvjRiTanfPePhXTRji+EsX0FCRdk0nw0yhTTAajRN+DEa
pKe981M6wzafF1dk5xa7zepZZVn3GkhkhRVceNVJm7CfBnJLFO3E9vYWfMqABvnQ
qbG1eHDZAyHY38oehYjjlQqqBIRY5Z4+Dxg1jejWmBz27MtvNJ+ZN2Syc4gPJSq0
iXGVn8jW2c4EruS+LrfnrljiwJ+yWl5X4gSEb+fwr7X9YwfEsn2tj6foqsKp6tIB
z8DxDATr8sqfYC7TOjipIwm8GwAGcoZmRmTJATX+/igYRz8P2hYVqxsaQduF4tLH
ZRz45CwaXm6X/s/qWbDpyTGZ8++9sBRCXCOg4oCQA9doNWyVQ2Xh3z3AjWYPH4WQ
E6DfRZkkQ1zwg27vrxkvPAphQ6mW/20ryS8hGaJIRfvtRX6CGiclQc63/B752KHu
LAXa+UaRPxBs9cjcKjTXL1d2Tu70aT/RdLO6nqvJMPfB51bA317AJharuO1huURY
fFA9jyURk/NnHLcgzkGWVuWMRhjWXWg5psk/bwizWuzdU7pK9HiSM+wi/Kb/w8wu
/SG9PcLN5ovg6ztYjj4O/Vrz20r4RwxyiSRyOZSakEdkQHS8J71ubZK+lsRWWLCN
6rGhzn78HNk/bi2A6ICyMY2Fq6EcAVteSUKLYZB0+Tf96TBoN9UOnnluwWhILMel
7x/4FtYMaB7SEBI9ZHeUS6a6mVJz2hKbKdqn1HQaZPXvQOfFwxON7VqoydFN+ZWY
YgXFPsphqwJcDJeUJGrPlXP21ODpbELPqpLKw6A/83mF/R2/eX5TIMF+5eCHYp5b
3GEDEql4ARodo8PzB8SqNq7ZM5V3vLLbeYALsKH6x98jcqWsPKP4ccsag0Yw7d3O
XXv5An7CkvkC6jRC5vX+Ph5J21U7oMWHUUOy4A2MdYrLCvGJtNO2HPgSj4FPA6/C
LcAIIhGH9DBDAz8Q0oqQWYkq+MKnSgev8tuyooLyNpoU94MXLWf1K1aQJmtTQ280
D/qwc8iEbV3029ejSFoz5j10F5PMzNa8xeb84zkV0nPjacxsvhG4AMk4ks0gGgT7
7yY98/NZyNs02nQxAGBpEYprdqH7TBpZjfzc6pA38iN+RkTlKYgTi3o3ePn2whQ6
9xaglbSUwWz2XQhdXIBjLIV/2cCeenNSasM28DAdyfluFk5cCtQMXSj0sc7bEzvy
vRrp/nueyyxvNITvAlUynaAV1O2QzEGVDn6+w3R23CnK8Xy9uBzXQb82uhmq+2oI
3hxuHn25J1TGhFCK1Mfbz3Lt1yzwNkCiD5GjmbturmFefEC7Ci4d+SH6220y6FtP
ow/oXkMbwpk0iSwIEi8ZmVcnjIcskksAROH+sAIDBVqhKMHvH55dxXm6bC43ffQY
PTEzUlEFD8zfLFPa5u9WwPA6eQCb2nkZyiXmeaJ65OtzTN7u+TJGWxvqwKYJQtcT
oEtd48UvfrTXAgzLA7scUiNIgOvwIbCYW/Id+W6ckY4lOghnWi1rmd59OrOx30UH
rJiB1S+dwoihpi/Ajq9zI8GHkNF2e84488Erz2G3QKHU9ITDKqW04eg0Vvmjicdm
cOmU0p/zVaSXCayb/DXZIhoUDqKE1oA8Q7ml5qaTOtCfW8dzflrejxInl8LLXkHP
At7GjZDXuJCilZ4PeY2PuFt3Ri6PYWYoD9M2a4IP2iSbe5CNDqe9cOwQV0IUgyVh
cBpDAVM9Kjptfhv/0hXs33iu5RqnN/g8lcn4vOlliCw7SdpbFUUk7Qs2Ou9YEb1I
1k+LxGK0JVGYJrFNRwetiGi+Xj28o6xiLpdAdgPWRlAOl1NM040ctqYQGNSN3gWX
BTrgLSAuwcO2BPyGEiGuVRavtMWhCtHFu8qT7FaZ6aNiF7tQi656F6RQ+GQKEA3k
BTfVlFZfLVBiG6dK54DqYA7ZoLRrCndfdhLswzdKNsKc8+nu92GSUxPmlXMAVwQv
SM7MGUBSSOFvKAyUkVIV1q0G1p9GNqbkF/twbrL3LIQ+YSEST8/34TMPFeYRS6D8
XpLQ2sbqCgY/ta4ehJFfGhHtZfSmYwVuNVqcCeAHMavEeaFJF0WmMjRVI1yPrmej
/iA2b+FxE5cTZ0I3bc4PBHLCTjZzxmKN23GVTYAKv7Y3IL/wAKeUbKV5LPFmqGfB
0ge/KdGReuV55Wg2FLOwaphA+JInin7IZPTfWlbESrse9tS0xxzNoEZbTHjd0jcb
wTP5w7QWrR631CfkKDjxWMsM+w7OUX4QHhjvff7BPBPTuSEJ4zlGVaA5DJQMauZ2
O+ahUzLwaRvq0bWg57Ill4hv9ZgXJnsGvvcB6jtQ70/K6Ng76iIH4VZZgw9NujHn
mYlhsj5RmpuxbQ/mbxCDKV67DPCRG55Hc6Kl7YsDrMeQee6rQvColrNNkM3txF5R
nnA+4FWP9xoxL7fckA5ui8h3UuMY+em/Akw+6l7eafl5aBNZNHY0JWft5o4CcxFI
Gudmer0Gb3zg9fCKKwq2BrJxh/vEkyAtwGboSs81DBmKGbErixxydFZFmKio3Xl0
2VeHiw7CVKnGAdd8eamQVygR1WPhurUNH8FafJzV+tqD+M54xvZ0z7EQS17NlYwN
DVk20zZ2kbhnhUSeKbR4bLTgUzdEIbw5Gsd1cuR50JZ+zZNQ+RSNWhn4TMbXPjbn
UuFRhT65dRS0SjhPSS0CM/KlZ6gwlA8yMR/6Ay3dOBNnTjnrF5/OgnzkQ0vj2Ysw
g7/qdmP7XhRIYxZCjeFCLv2v8dFpynyPcs6y6I0C052LPA4c6o9Q7z2Mh6LBF2Wu
CRByfn5CuhuDp2fbedXvN38qqQyDtfOFmPuTJjzFY0skHsRsBNQ30+dmSKid9hqe
55lazR0Q+GOIko4QYFLHbJb6ilXyI5VgFaTQB1J6w1revmR+L/6nKpTvA5aNt01m
5+XTgPw5kNOTr6Ozq4oXtB/1wjxywz4Yxa7C+jjt3SNfgReiHKIYG8HpHF5KrNeF
rKYliTkvAjKWST+2dzQgUBkSLS9S/41b22Ohjj8u6eC3f8dCd4vcIt9HuzzzVPQH
fPDZpcSsojuX6E/Ff1gIIdtg6m/8QcE9ERschq7yBPDuyusNkwcJl6HhcGcJVOhW
zDDMNDBFJl3fUNq3LsROLE0mkhQIUeLjM1G/TcWyD9L1aDQ5M8Lt6+EruS9pFfWy
FwuA/cI+qtprT3oNjBgY26cLt+I0r9LTiJ6YvPgLgf91uZM/rPxpnv5CndolbnNE
Lvi+OHD7P7JoZHDxatuHPPZMeawjqkeg8tA3DYnkd5Vukdl+bAkjmFG14/88Wwv8
8FDwen2yVB27ic8yB61RjMeUdBpP2CUlOcH3cb46c5i/STUiz1EiYgxENR73M/DI
XRaqF1BLhx404UaAS6zbbMMMp0Oi6wYPbSjlJBvuETNS/K/FbVn5AUM83D5+lGtu
Mg736K2mMbSopySyBKmFlNqKBe8CUjhPWHjj1JGvb9TQXe16SklfLbFLcFpvszaq
KCAmpFrxIqvnb43LVLfikH29xP9+3XE0Wgt4VKTa13LqojdNYHcwKWRTW86gPw6N
2hGK5/HnfcpInHG8Q1j0vwrkBCN0tgVgqzqvvXd0rnPtruRHEneNGasR+GI2vvVz
VZC9APjfxbaSiejuJUv9pYYmJycKYpsjmNIUUar50sMHbFsMsn/KuevBs1Oyx62c
N0h6OiBTgrsd5t/vByO3I4/h5Mx7AZMFDYLYxaFwp13HZ3Bx3jLxugSNXO9KCR3o
qOxFKfQE6D408v8g44qo067/tsg6lGXBXNCf4aVUPWptEPawyaeDwP/iN1dFCakI
QHEdCOUgEBywkudISvxmAjl1Qrj+a6mNPhkOBYm0YkBYVcukfCsVNViU2k7KgJUe
GU/+Y9AvXvOcO1JjnFrch/geck6x8gH/0svW0oetF6wujG4qRw59y4fiA4Ue2NN3
glx07uUrb06D7fU+6p72Fdvv1q1rzMKgHs0HtAI6hOCZKGzaCQEjsquFSONcoFSW
+AIFdWbwhK7B2h9e3vhdC5r6U/MQNWs0tF7TMj0r2rPBDza5T3VoHqq58OYGHUvR
czDaiewINHwhat6wJinGwsqXzvtMHtL2j/R4n0XruNhwBW45Suyll8xMHWErvX0K
yI8WMa1OHFShsusuHvuirhUeawhbbCU07nnfE/HoGwYS86iIBCFHSOXM8FNo1uew
0FwnSaFYmMPs9XaElzklmo6wgV05ShhGd0wYHMPkSPzUoF4LTLzEoCgIerAVf+1a
BSzavQRMraZy8kH2oW24d3/DUaHpKAHW64vX3iqshR0NKAiKNVwjqmYZq8ejFfTe
Z/CPBsa69cd3b/bfItSunsRXHZ3Jp3kc3V878vsDLhZJc9XOHkn/vwJbn+o6zfb8
7lef2t2IUleBY6yYqEofSi0ait16MmBqACimFiHQ74LYxmKfpBTg3jSali3NDdbV
1m5cLDTOdi9pX9KOKxSqM6KoIwzqhVLOS9VjSNqXdiYXAIChk+cbFU/42dwS7L1n
zSvS3Vk6WVU+hGL1nGyd3qjZuVeCbpS7kPO3B9nJEZk48bqcLC7PWY5FOmHS9Nxg
z6RVtkbs9bth3CSyMn8og6WsVuTvWi+1GstH9f/gjZ0KeYgk5nErT7CEmbQpXxPf
AE/jI50PpY0RDzs1Opibj4T4zOVdYkXZsBEhyvdsWxj9ipeO+fHqIFM9eTrXlipo
xn8LFce8/Hog38u2SOJObOl3OfDD989RrWUZCNZYRhbqlaIGjrkHxjkcPOayCTK4
for8Zpd/h6gmgKSJgDQD/87I4k5eaCM5ZMsKpWiadugx/7eIEF5c8pw+g62TcErd
NR4gllMY31pSwPH+fGaiZ31na8VIGiue/K8faVGaJjt08sfSSAFon5zQ2yVZWgVq
ds/L68iqgxW6jGJ5BLelvJkrmh3fvuSa6+S7vzX4Njg/lds97JPMaVY76lc8L+pO
MwoxomKVHvGbX4esCAun2IllHn2AvrOOzN7WcFV3Mb4IpYE3Ja8aXfLJ9UaECf+m
+zZ26e60FG6qdjnJ+h5FfgUukeenUjEscvEWXiPzVoUfJ5RnW4uNUJ7DbigDSrGj
3RV4oKc6LoGIl6ZTId1JzSNyyqnsZH0Dz4miQ6r7GLQgk0QTRI/4MmL9MeHk1Ca+
UvJRFBOJfkVaHlKa2Szrbat5ns1cvvFuisK4dHny6SOIbdMUg6G1AZ8AMPVoLf3h
ex1H9gOYaoE75IDHETddmSDaLSp5+t9cXxKmKTjRAVVGFeWqsKrocx0RL5sVjod0
cbkCHuOMKBZBb8antsiMfXHGV5jcJgDOZHqzA+cQs+u3eW6Z7VtV1cxWhvOyVq+Q
Q5P/bChUjT+eZE0Z1iZOUuGecgc7D1XBna1erqoYiqpIk/bo+yd+SqrHaXcEDgOe
sLxszz+4dezLYojjHX/lCtuW/ZAGJyGQNXG4e70v8scZSkTXVhF3mE40Q/UUYJLR
OgrJVO8uR3dvhybkiVvAkRlNf/RVwT/962deExf603fNh4UZNsGhog7BlnVwlPzc
WiOKRpYjjWcN0dgGM+5+tAo/4FkSFF/BlSb2MaDGTvDSAcRL4WDZzS+ifWZTIlLe
XIS+HoGk/1+Yta7W5ft+zrgQCk9MRiFMoO1M730EvisK5ZE+Opd7+j3k8/JbvSz2
o8f7oxKNU/dPh/dAFLyQ+PA49L6KZ4YrmZL6m45fES0UzeiORNQ8t9oQugSC5kCK
hjDtNZTUNGZk7g5LfVdjZic3dBzHPsgZz59k2NBFUVFcseNKZp955K659T6Q8Lwy
7+VYKQTdEAZ/Dl6u49G9HnnykwCmoKeps6TBphI//ch7lDvoB6ScrfoP1YmZ0eQ6
JIj3PYQUL0+EYDGZzGJGCNEsk8B2GEsiirRuizxEDd2xDMapIiFJ7ugvOJFGGBSE
IE53sb64JknmNgm0Ta5avLhrW8PV1i/PctRpVyVMZEwxpY9EpPGBbVdYXF2nxGCv
uHPjSpCAZ3VklYylBWBgRIXXKLXzdYQafpLKHemaHzs282h2G4pYZlkFVnlxstsV
Ppb0F0hmptobs2hqWNle/LYVK80nqIJB25acrY+uFVo1eg9johIBnGkPzuIxoOho
AC1qYZ0q9+S3II+oV5gccD+bp6/8O7sTE/Vv9Aj9ffvlOp+4oMg7hyCbG9ALYpEu
Z3XSi0NMRF8NPFDQNnlZ5mQeRdaJWlbFp5C5VA8GpFwDJlc1yhqV9Pw/Kbr3d8IX
UEJJ6vc37mtOZJ3NLD2eadjGWZ2qzJRTZCGayImNIHJxlO1qmUdAdOb1aDY0RyNH
W+pwBAazKwfY0nESoBFX1Mtj+D5CGW4/1dGCVqyAYPAasfH1wTxoenWyNdXDyzlM
TbBoTBERSlEBf2DVBCjxM4Qrjvn+1wQkszZWztQYC2JbOMOxi6SxJBrYnNFbnh0D
kkC8zN4OD0Y9D17FOQGfGFFJJkQ3jmSRD8Vu6yu0tXJQo2pjbz7jQm2nWjrbiCZX
yLoVpXjUNL7AikFMbaxH/U1L0FdJ0Q0fodJmL25jf2+tsbfFVUoa5zQ1ixPUTckE
CZo97vh4oWF0CPIZk2lL67hKpHdvfoXsWn4CBFQVbhAdPlMwdbN/4M01TgDFtoes
6IG3zQIhSAK8AtkPLHEMpthR4RaPFIar17kqW8kn/PpqgV+sxKmBf+1CbZbx7aQT
VjAoAj8sJmrsVXs+JlPGfpb6gWh3S/H8KZvbicf9jG02VMHq3Hiio8J3jK/VQvBS
+jFVDrq/s62zSH7/+cFDWRyp3BlxxzCPjDD2c6phyCCj06GR7rLoi1KrvWBvZIgF
6CgasOAn9f5WKwuvkfMgI1f59dY8jTjNyCl07acl8vAP7N1CCgwJSkqofjtf77Vo
Uii/bc66cbb8eqPzxQ7Lh4wpguhYtKUE6CLRN3oLcJD0alDJVzqZj8PQmifZm/Hy
0151bJgQbqg7FfHgvrXJ9kyVGmqt3EmuEIZjZyBCnPRRiDkULA7wVIxVsKhlTUx1
BsGPmVQCwTROuJgRj21YzCWGI603hxNcSYqVUA7p+7isLS80C9lXoLGk61POTSRJ
3w2NJHVuc29cGp9ied7zzFmN7IIYYqVP+PehjkoqizRsewBx/vZjLIL+lLUcJkwP
lCyCZwMLvhK3P4y20qqfT0CQjkvSDrw6kW1RM2Rtu2xDI4wogWUGAU4PP27Srs1K
oBNvCFIpM48wlu7EpRkpQiZHLlNXj6ffsUtaKwbojo6/4O5OyTsEM6QhljPqbhP1
+d52eIcYEptWtWhT1UpMssBz2joHn23kwsxoY5NywDNdKzDk5O85J8dz7BhWkRol
tBys/8yw7VhNSyF1V9XuOYScpqcuU1Q9vLSBtkfZg1BeW4N6DiFBinoJ0ygP9LeQ
a66I9eJtSSv59c1TXBNuF9OImeX5aOBICMDhn67mkilyhXYT7goyfpSHOJ+7G1Z/
ORVU8fg7xZlBQqDzSMIpiK5W/3anaATG6WFRtm4M9rEvXZLGbnM8b9qzHuY3AL5I
DyFK4hLVNOPyEEXpXwh3R3zYdFoM4CDt2GdlcQezVdqp1kVUPG3MrmCSYaaea9uS
1RvcdtIT+UN1eWKSv03mok3IXNu1UWITApxXH1NdZru1U3b8wvSGV8q6K/XGlG7D
z3XPCF8RDdNc9Jxdkfd1MNwjoN4Rjx7EzT+sqBuckNYuJMN81H5Vvk2qjPb0+GE9
paU7Mwfb+mDQW39b07UOYw9wQMJ0IWIM4oStj0Y9dDZ7pWFwp8dTYR29LUXl4hDx
VPJxFy9b951zlsyYKn7V1iq1O3t2x1bX6/K0CtjC0jnJX6oCV/89U9IVz0BASXl1
3gZC/89BWdGhoN/QvUw1SuXapIIcut0kW5d0FelBwWjfHVXjEEit6DyQ/tIcktAa
fRsnCuv6k8/kLRPyusyHQPm7wu2xp+xicwhkXWhQcAdR/oiZzNORIv6iaq0JGjsr
Ef9yN5N1S5DX6pu2Bxu5nqayFulleUhkY54b5oymyd0OH17tSsBDzg0DNrM3qZ+S
DcCJTf80nM5JqOV2Q6LB0eHNS7pxIav7PCoc1l9QRu/2w5c1nkO5BthE9yiuIV64
to1qZQaduiPd2GzxFzrRqxt7rZsk1Y6YOHvW6IP2C7o3bfy4Ku3IaAQaAb2rOSAh
pVpSvDjXLS0yAru8lSt1Z7PRq1aQTzIqRRlbAp0gZTnZjdPYx7BrvcGjukmqdR/T
npexkHNbfnFQwqRV6ag4WxLEB/b3MTUQ1gKGCnwMZnGO3mDMuSIhFfK8Oa2rg9V7
a8PKOsSFm7YyOLuld4Yr5UF5OdVhwOZTsPnQlwTnRWRibbOCoA8fFR8fOIFi9Oln
/+nCUDzoYXrZ6jx5gGD9i9oQnVTeqFIqAOq2znd1mNRrlHPNvgN6wrWJXzvbmFL2
SIXdL7ukTdeKh2rgzQGUYu66HKJm7O8bYznsfKlWXzr0omRY9Wt9FtmcKpavwEfZ
k7CFlfAZ6cFWTO2uuU8I0gZ90PitIuGM4zROOTuZIBozz4eM/G3ybWbnFyvAlsyC
nP+xQmIbX4vZ+oqvPKB6ufAaXLPiG6zUBB0qhIOgMkmPFaMmJ+4E5jqrkORPYr1l
+gEbsdhv4MRiDzWu+B/70BmxEyOPJ2fGP+Q9yDGG79V66/lcW8ByKdXVHZxnVD/R
gJKgBZUAK1ybds6rVH6sgtfSDs3//kLZp+uSzNeYe7cUGu1EcoikI8EmIwSQi7QX
yqq6ygTL+viGYLjo2pAqUB1IUdCJmYZBuaY2immen+TKkQzWXIWdmP6USgevjW7n
Hbch2hDc51ox7Eof/OeiYjuauXGgjICcR0eo5RgFXrYH6kmI5nB6eW4r11mRXwuJ
k/hk60Gho5qbYwVh2Xa4FbX2e5U6vDDvDUsGYQbiw5aghJdW/0xUCL03qjGZ2pyO
S0xJCMGHOyT3nN4DoDWgi15AVjnyiUxUAlpfMfFXFfIUwWvukbTAnThpSVe//g3r
+RRf0aE7j290b35LPsXjIM8aC2D8WR4CWE+XEVPUKzSxIIvlskvm5K2AZNolZBtR
tTh6LJVC6KRtx75ne2HUwqJd09XOiCLzjpGbCXpgV6IzUfWWN68gLlIUkyK72yX6
f+/HGG7ncIL5auRSZAm0p6l9ceSVgtrBqPzzNqcXjFqteBEeQrDwHMkG/Nd6oTjV
p4p4LotbKE21adLHdSS/XixJvsj+6NdGIHU/mgQdC3CNXmWc6Ds8SWnIbETYt4lu
56OnB41HtUcfdGt9z0pcH+W6rmHrSQUGESa87W9UUu32c5iHud5BH/x0GiUwRrj/
30m1BLEuKRV/yqxeD0Uh6jZYSS9sE9aDQFcgzf0Xx6NE6EpUO77+dxpPtf5k1pC1
RJdf748/mC6kRbyPLN3Bh5RMuVx4pZVaiZ2Tm1upKP+bT47OIW47/4RoXo3ZOHLF
PPjpHt+6unoOMykEDS9zCrNikJ0F8cXBAq33ZZ5M3cXTAx9huDUatXdo1vj+EU3D
UpZeaoI9VQa7UAt7V5wqjzPmKeAB3hvg2Nmbjni9EZMcUIivBNJlHeYgdqKAvJsb
RvantoU3feHU5fqlTj2dsc2H+WuxaxsoVxO6mk6eUdA+WoCbGaXohhB+dVh0G0v7
Of1m8OdfJYODSAeukDwYEaFa+B0ja8YBXvk4SwhTJC+nRRfhmJW3JUw7CePWaoa3
cJCuMbK0mOFFE02fUtHx14ARvQ0kAMxAerg+6Ku1Xs4/jLG1pZo7e9uecARAA+A1
6cNuoZ9b8C4yhP7ZK1ySYCCENXsd9QJ2dh9wTMfbKd+VuR67StaTx2PP/06Ve7Xi
WCgQIoF42CyhagUv8pxZzSxrE3K0MqIL3HEEfWh/mmp9jsThk+3Vvnr4G2ZbzH2t
FD9JQmbeD/lkDZ1VcrqvVHzqO/PEEVkXkn8yYlOr1QXyv+S6hzFKxxFYJuPZmJXF
zW2EF0WDliMTGILSAldbN3iAACexQJRU/WfIlF3N8cccGFrqcNz67dtAWo+ke00Y
anvdxl6Mv+1UCxyT+/Q/jbxClTaAVF41pkRVbkb6PY7OsorDmh0ZFYIAGOjDk/FB
TA6SeNTQopXB4hgZuhbW6EIgevABux9+6QJFrKaZVqdb5OIvQ4SSkNZYArWjUy3O
k2G8XD5y12rd5ez5HIeJTrwODcZrjx9HgngxAVRPlNneazuxsADDkj+AskQGhX+u
9yT9E8ncgJCn7TFYTTP6uyh+jAXHDDeTksbsCpK8pTDefgOQ93o7jnFd+q7FsGpu
3ZVYqRLIdvHtbe8VgWuKTA0IC4QrLXfpW0kZ0HIAEznsjmuRruEcmb22eSP6971t
8TuEPoagvMT0ha6vcUWYo57AH3SWU+2Fx5IUxrf5iLLBl3pfyQ3BfQsKAxThH2K8
MLU/T3GFG67fo1m+xkoPKN2z2/VwhEk3r/JIMMJRLD/lEc3saV9Bn6FDNru4gRW7
JxwH+zP1up6CHB/sqOAxAixAoS+BDrzJtmW891wYtEdTJIgFgGD/WtkZuMzrYlro
CYVNvzcqn4kI0Ar/QMoj3aMn42D1BJkxxcqeCmqSAV0abUcJ8gOx5tEoco5rC6Zx
ZL00Q+eycdcawHA5hRJMXRGIlZg2J8PwqEYsLHtkx5xm7mIRtMRLoaiXMLkvwKel
HEtUhLUPCmG4YXYIKT2AD74SW65bYKrhCq/YLLSWX1549tx7MaQ7SX6vs2qHXHtd
iubTitgfSuvYgKSfH6g3FCOtsmTro5xOC9+7EKqjwNdr6+6OBAy8hC45HMniSvpk
xGCDsaOunTsv1Rq7lVOPaAqnyBjISrng94KG5PKVspZvb3N04bocjl2iQxws4dX0
y0Vv1eUhD5DcLYwAkgA0QDh/+y0gHi/pw6GRA3ilEcQJuNqRgMmUzJYjuJ6rLexb
MCJ+uw80SlaHKn8GzNyxATJ7sqAHfas2qOTUYg4GBQ5n70F2uilpLkSf6SdiTK52
o5Lw+OQ6QPgyzE2qsoCkxROHlSMOEWd9lnrBNEvaYRTf7ZG+H7nn4DSNV0OEvxU4
5V1o70mGaJVAm/zVY3NRA3z/zz12yG65U5KP/gvN/QwTJv5tKyEU1qdNtciJvaRZ
+9O5PIrS8YYD30j9kE0/1Nybsan4/QbcORWSOnOdxuIJ8qXE84CeCGLjPQD9OlQX
3SKHWA2ES0QmOTEXuoGu17rCQ5Yq0E9J0O5sFViMzB8Ivk85JMPtD+8HruKCMqPu
VyIdMnzubXbomiNfA99vr8l9HmrNBEemo+56NQNLXvnf8ClpI7lT+WcbMkmco5IE
haVzsy75Gvqd0DHe1ZuxHofX93b5mAyTT8BBa59n1NgG8OyrW9I2SrmQRNnOP2bz
75DxMCrBRf8F+Oad5ZGF83pKm0hHF9/OKiuk/1sCjdeBGFTmWCAr1dMhroZhfhhs
KPyLxkgAAnb7RYCv44M6f2CnOKie5EzRbRzJX1zfuuv2DCkucUkkz6/HtkoJTTLA
8xD4Ukr+TEVVsOwQkr6ej198Qe9dlyIxLhtoGJSFJHRzEq4fQMRTMzIgF/ArUTsx
3+T1CcNp/tWtS6Gb+xh4zQ29crPLubjWlDIZ/KPMkts3AvXQ/1NfndyDhiO9ZJ5E
aFbjEaOOoqYvbNg9V0ClB/RgP2w94SjcMVqFmHT+qPMzttwjGSsSQTSd8PgybvVW
q0lelYabMqDWdYvk6hBk9IHRwpY9GcQHKq5dhvkKda2FHOomvn0mYgAHGFM0uPds
KYcQKpTB0bFKXITGMhDvjI5ZmdANCCCJDpJJuA7Neccq11usD8flfI+unwdb4WjH
tVLuJ77zZYv88zXL+7k5do36yIQSXFJP/uciF/bmleRZMvkLEKPux4sLN5yEC6Bq
mmEvPLLpeRrn81knxFty8vQEPUW6fJ8XwC7dD3DYMeLG+GZ+Cube7gNZzxrD5T9F
UBohbdLNSq1nvXK0PZIRMd9NNgTJfH1ub6oY/JEQU5sDlHxGu+Xlc30ub5bPSED3
7AFsMgR74StSdP3qX5KZ5bogW7zaA0Np33+0e3bgYU65a5ZkLTXy2TWnQZjxDHgX
MS4KNzfowaboIesZBlg3CWdYO7N7yd5QDKZZCku2JFGbvBy5yPynAS8N472mMTKb
ThCAdsn6kwqpnm0W2LBmryuJw5mbj2FbBsqZqB9Hyoc1GGbWqUebLZzWQZlkTNzn
WqosWmbHytJWhvds8blHLX+LWp0rHFYae8S/N7O2lrbfDff15NwQZAnHlhnfjm4K
LkjfJS9tFUY2L4thPDF3jLmlZVagJK7PlPvgQN4OpCUaY3DercFGUD/E0ulRFOaF
3uSsvLhEBr4ZTTirvmLqIFInUVlHkHCF+1CU5kT0O4K03fvSqTGn1GjPnbJBt7NB
8zRyRKugYvZQcRnnQ2t6GKx/n4G1rF155dwvueWMITUVv9dO7P7WsKUX5qMW4Ljf
4qvj4oDIUey7eLoQ0VUlInY3qhCJRuPUEaRbstqcqvL/EQsLHBQ2F3tWgZsryhaN
kvZJK4z6tBARgxUOHvp47EpCBtR3cD+WEMcyNqodTuBGL9gmB1bkW1FNs6sWBXnf
UBlZJA4X1Vz4I+qBlzwzaDWjz5P1QGNzjF3Dj16t6h437ViNbzIXoKET32sqkBv1
mqN6xIo0FCc3OIWwtFV5SUKRO0TmrHG9clpUEMn7rAIlJ9KS99YDvaO/iv8vWA8F
9sRPWL4sMsFcOf+ebcTuaNCr7ec6JHShmnWL+rKtAFaaexa/oSB6zfXgUV1Psouy
l6lhfOH81toWuKwLeJRKMfKMPBVnnYsu32WCXBKPlV1ThZUJhWj0eUUg5YGcgijH
2SqVSlnmLblT70EJgx0fMV4Ke4oyoxBFFavUi9GUVJwp7z2L/OjlbaVoZlXD6nGy
fDXfTP0zpA0/Fu/hQvHVVHX6EUVKLNQ4DCH/1AtbUlnU6FerlDlTflX86WzcZ4ev
iopctr3+rc9YQdEUzS9MHl+2QfovPSL8hk3gOC5VJ4psYn/fkYvHeQqUwcX137wC
DG5bLDTZXa/t6ZzhaIwpjFxiHZD4tgwwS+HDjAVq/k9FB03zO+YavKS4bDMXNNRR
uzefcjzqwdLIhsJD1Kn4l+kJvgY2YOKgjE90V9MygejrSQOgPNjOhVQYNZJ7AJBl
26AaZqm1EM/lJBYoLaGYEIgc6/1Mt/Glgkq+NydXLwDSRlxT0Pl0UTMawjZnyNOp
p4JziTImYLmpXyjIAVs5O45vikwmJDF6IsKcJS1PWgPWRDHazxMPUoEOs6I0zX+z
pgLMh8TpsMDz2/Q/DLCieggrzpRVBINzlhwKbbL0J6+YVKRN4KVI2XhANwJ0Fb1v
RntJ74rEJ3CSnbPKfELRqTko1e2j5GzizE7cQWm+mk4R/OVgQ6Kn18u2e4TJD1kb
zqB05K0UMheZdKNhywrd/YqazIMImYKtWYWWz+QKolgbgb3uX+kyJm0y4KHNgD0n
0ZwIaWIuUsFKyocaz3GGk9u/PqbvARBF5IG8MdJFI9x5cQIT07witK5ghQqFd43w
min2nUyvR6LsNa/6RErfTDiIuggvIRKZpo1bV5jagSfjUKQoJCnfD41JsA/XClTJ
EZILnsHZ3E/Boco85dwrldXBdB3MKPtIGLWnFyubASC26TZuy7hR8T62vYoxvosP
AIYuK7xoZkYde514aFyZ2YvRPrrszLR7aejWf1whhTqXPyeqQtLjlaSFEkkN+07s
i5Y74jxQJMJos2VDg3UoLT8bBal18qgCiLS6rqtqq0fBosTkfY2BEYY8elW80njo
xaSEIGcu5xstEQE28kyRE1YA3CgZk3hvd7TqxZfR50Psp+Wd6Et3tDGW1D0/WSAO
unTv0Vt93aa2FGRYuCPu9OLbSYBlcw/6mdB06W+yuTRbaIsDCVqAtid8BxvAdSvL
j3d9APTD+xj6LxDzf01519FeNvYL0mysDhlwRedXgyvf/wGJGyeNMyZ7xY0HQhYq
xKQsraTyyrd2MMKz0TEjniAMawLwVq3pqvoZcWHQ04QKvb7YtP3ZRo1npVBP9pMF
7pt+wXIW8y8tIfotuo03r9duj4Eod0AFgxk4Avi7i/BEnlvOiYWt+mr+hOwmmaQr
gCJrU1z9nvmVvTKkg+OWpD9Sn5HwhV4m5D32E1aDb1rSvPNZgNzbCpj80eUEsiPR
lzqt95d4/L1DOooLsSN8VuNS3a299TbnJKTXo6A51DiC4K6N+mFCxzYq/nYmEqNy
mHs4X8SdEgIHBS0n+agYJdWr/S0o3IQO9asWXuZ9NfBfmq5ntQSHWfUI59oer/W/
WS3j/r2pzOiIff+z7Twmw6GTyd1+e6krLqftTfe40v7uWor5UVM9wn90g7037zon
tXW2mK4J8/8oEbnuEIvq0hd1/l42Dc5F320hhA4d05Y7BLWqFdFZQ1P2MisHm0PK
NCmFakd7Q/7WFQG/dg+Zwd+P8fQi9PCbajZLyAPbgCOf3o6Yl8aOJozTmQ/gfxju
Til2JaV/HawrcjeOSKUImkvs2HxE483z10WOEohvAoeMDkFI1p8cdgwF/OPXbOOV
EnTh8IvLGWUHgGsJiKjx/BpGmnEbnmmQ9uFiDGeIDmOQNWZBsm7kOB85d5HE5YUJ
K0WKTVs5x18jdOtTZBvydhoenaMne7oYhp6apNwEFF2LLMHLBlE1efbeCbcScJsY
J4cvsJflRg4zQhHExj3412kkebLObAa0u2PFT0Qh0KUomQhQf6Yu7SafOGMDH9Rz
WBt48+r/3SQNWLfr7IcPZ8Dpjk5UP/Hft49Mokxzaav2m0EWhR0oPTfBDa0S4mhT
IeqK//zTeLUDIFLebgdinpypMsTQPBe3iJrTsyAgnJQBghm+il6OzhiO8SiaG9qp
BEb2Klw9cN/y3sPqEllpWvfpbkHWU87DRGDTZ0vDbUwU8N37bkeL6O1rJM0xbR22
PG8Im93RLdV3idm9+lTHpkH0rTWB2MTsz73Bz0O0+TGuKMUR4ZR/2huyXCcu5GmG
2YxIu3NIMInB4b5FuYPHrcI/hXLWQISanCDxnB3jWzXts4KsD7letRqvyPrEmeID
0x9VhOzu/wgA9VpkB89HYhXRG3ItN6XFjtp7bCtfHJVJKnisbrg8Q61aUOd8nP1b
X9JUeJAv7W2o8HhCGnYBkg4+itOY+x3mWiU5bApRpyYt/kp761QZQ6D3AxSW1KyC
e0UfovFOBuapu7G/vlWyupPa/mvHrrnWYfcJPZxeAMPZF5B0rtODsiue75yb75rW
T061pAhuyB4dlTRnpTTmc3Qvx/TRcDqeEbshW7vcnPljlWTbWdtdAKmXemXXLKnV
2HJ7SBs+lAiOPW6nh1PRlW6zI0g4QgitEQTKU2fu6RO1cnXQjKVoGJIfIu6RL3bw
kYs+wUVmSXOHvtqkQEBAr8tdO/aiHwOts7P+1+dLykyXv08t/HpHpUeU0NrV1GFW
z4nMyYGmSGf7NI1HrZeb4D69CUdWHEpw4+JQbibsjoiDmIBqivbfXLG2ww8mz/Uy
2tbCvPxInIIVc4xoxqppzZZ1yHlRQvgpyg83FI/b0F0/Wlalv3tFdQkiDzfZIT6W
98No1O/Zv8Mj9QbeazzHbFJKnwuQVYREh19tJ397YwYXfBWwIhIls5+tqIhnUiOU
uxmY081yPoZuS3yqf53R4RHujhzu+rZBQ/J6jb04Svg3iKCta3+K3agjFS2ZtQfA
jZma9Dux3+SYErlwM6mbQYbqGIW8/YShfFWact3fZPB0ybIEh4VTne/1QnqI0FcU
GWSxJElmrWgf/f2erfJLho16+p3BHF76AkfxWqT+HUpqrXb4QPBWyIQ/+UyZZ4jQ
UuJSh4XAwdo/1DAL8SLqt8vdJVZ7IWrrIXpA6VV7vwEoNE+gymjUkEbt5MCzUs30
9nAky0CAYk1GNcYkNZA5/s8BRB7Pp4fhk8XGGKdx9eJOr4ww32w1MnEtC7EfTIyS
7rjSWYV5ofbYFgqL97mJJ84Bl81SAYYVhnddKHY0vqcXRJXT3EOc+OIPLvIf6lKE
B6g6ETHdWWh1su+7iOppmzv+2O+2d4T0J9KalJrLqqV9mrfVgZLdT/xaSjOqklQ5
7HN0izxNBio5nlZZTELwcZKI2+6NIekDamT+nefW5qETDwfSO4lqGp2LZkSDZTEP
pEn5vBswWZbVrHH3+WQTVWhiUqj01rb2cW/XtHiGXFMpDL4l9kx4fnTBmLCLGyQj
5Zvfv/ZHrtlI8Lc9cqXeHByalZHef2BaQDeZd2hwrYFaTvkMK5Pjvjvw1ATn3GZh
MZ+GsYZwj+qLfaVqZsV9CUElRwkB9jTznRXQhbtoeqsu1Dtq8Pf/RaTW7JvPOiTy
l0T3NDO07McQr2QmxIRL/E2pI0BC5vGRO9dJsGsFcK7YRZ8bRsE84wIjDJdlxYum
cZiBiJlPxFK/ha8Fzypq/EYmhuelwU/+iUvbZzKw32bdIAwixGHkB9MW0+Sb5ckW
w2awSep0S0aj9Vc0ijon280cD50EpL57Z2aUD8RelfrT4X6AqRfMYg2nFGEJwFu+
yXQV+M5xhaxr7G1gbCfk6FE60K/UKcqjbmzzcH5jqJ6falr6bQcmXLtlfcUPXcPs
zsXmY1dLzHqQn6GsJt/EhlnclhnB+j3BTeaE9gHuYUpLdcvj48/XffcF5PxqDuX/
aweeAB9EYSfdt3QSZGdg+KtNktPzMeYrgovhFs+Kvv9P7kwTPLjA+BfOGBGGxhgi
yIhPtJOJPPerCggHVQyGIQLmF/suuVF5Sog9X+ehbL+FCUHCrIc/zV6YWwve7y2W
H/ZYf74SbYGXt8bcD+D41rQKy6HfJG+Txl01Asslpe0Yh0z/9Leoog3XC9XSHjF/
93Eo9Y9ssnrudZ4Jvy8/9ffTa5Qy6tM30mGGOR0i7FF91LakaEk05O5BgMOPFF8O
zwyLz8Axxb51gFPjJh5H71szD4Df/sXlBTPgr11QxwitYqfvYvhtrqHxFO4a1GEI
SZ1GqXgmR/gfmPuuS7PTCKtOqrnLhKYHetGld9QYRqqkFWtH3uCfgVPcz0UMJUYE
DCQXb5e8A9NhIMPVpHucJWxHP1QH1QIDSWIt4EkINN1TRi4IbZ58cVlJu2jOIB40
9idUlEdCGtd2cVfeeiulmREfQdUdSXv0Z11V6Z15yEFeZ+ORhToJd81GptFAFvXm
q0ATMBuBSm1kC+ru6Pzn+ZFtSYZJvVQ6/5AwjoCMTQAXclxpNxzLEZSPHe3rqCk2
v6+yDpD3z/YsT8Q99XLpjnhVR+f80ASiysmETxapOege6N9J/ZNJQNCRT8XqhoJ5
ZaBrnUahtGE+Ogf2alXbw/DAO9mOkCFCc0wMwQmtZdGoJPY8AfqMjVpO6FKqo17e
e9gWeyr4OYwMAcNeIJdW0b2yD7+Ml4Q5m3Rgt0YSFNJmFyJI3LEHvOcJPiolkd5E
GqvQc2e21Mx7ILTOmefSBJPcXvMEgoib2k8QdlpNsb13x6XUuZD083cQImpOdwlC
Jxp+WR13KuvSxpsF/zGu1etaZv2YjJw7iepr8Nl/+ZWPJmVXr2KTS1c64VwL2Oli
XtRhP30G4Xh3GLS8TMaZpFDpexG+KlhHEXdWu7+D4Sv35Dj5WRrjP/0dgJwJM5uC
uXoNlwTNYnX/k5odu9APpRJrYu2Xhp4wHwC+9iYQVg2+FiIB/ZdXFZ+OiPEAK/DF
8V+odCjOEwemdOHJZo3tOOmPw8Lj1WchqcQ1SN4dns8yDB7vkP2/OCjEjBmMnOhZ
uBp6rkUhh6fn1a1sDPHPPdKx5r/8p8V2LTT1ZI848/anJZTMMI5/JFo14dx7t+lC
hlaoKyXVo4oDgteIvrP9YjleS2qE3eq670dQVZHhnFFwAVLe1cKc2rnirOZ0DpTy
dwAElmwkh8ROQKmWJRyNjpRO0qkSPkKR7S3CXCSZEEGc09KezDTIGPBgYuKhr0Px
nGo94xkIdYFhYqCUti7xbbZDfgNYrtdy65gNeRJnHlqbmIB1mp3vJhGUQKrZZ4vR
9WUELS0Q6vDP4D/+Oj1R/D11kNz30AaMwIsMixZfclNYiTjcXRTKCB3CtjhUEm3B
OidMosQwLzzemGQE5Fy702xQ0f6no8Bc+jwp808KHdqHThaqwjhaTv/SOA54JLyI
FEMsUo7q37p1Wy/Co/StQyE2mLuyX+EJ578jKwGumh+BBEWqrxcVhvyghdClJgOE
Y8j1W1eI8yO5bOcANBRCika42ctrAwk/X9lT11RaYATT1A70+sMVoXsVKuCuo1M5
zU1j9SI5AgGIhQP1eJNjjUadT7yGLVX4LNBM/lbH2naKX3Q4RLb+x+kayb73YkPU
wvn/lwBcJjn+61TmsHAVlIoZnB/k2fXfkYsnR8v9TwWOaYh9HiO1oc4ZGS22D0Jl
orwNcP/2ejO2HSu8eYuR3jOxVpHE1rsoG6HkUeCWvgINzfXNmW6vzy0gV3DmEBDz
RRBwiWPhQihb12gLQhmUjNTz0XhQeITjSDDXwnx/xX24Pp+KagHpjGh+CbP/t/6O
lXYbBpck8EI+DOXMaU1dDEzKz0CemYZBq0K4vImXgH5aQxLbgVscePXeivo2ZkNv
KFBWvAH5EVtWGohevXPjQ8X7K0lRY0RBHrP2vDX0bNa13jhJ0ZqvzQ9o2zJTQPLa
u7c/ueC2CT5q7q+ImOWqyt2IvFzynyBEPmviyYY1Wf77SVdHcQcHS3jL1qvTHk4v
eyy5edtoVL6SPu6BvIRgh8FRfeBEtYKU8X5DzvIRvgY7xaK1yRiuUDtTWjuLam3/
oHhDQMKUh+2xhzxzEw2PsZoPQqnmL6euJZKvA0XZWOZ7ZHJ889gM3bS06u52IEAP
XfinVfPDSezpA4pfLVhEA/KOMLXo6CkVUUnKGWGwfQ4JgC8ydvf70gtgZkKu4PPO
ydYpQYESmowOinbNTuSXgq1VfM3bQT9T0lt99MyfZJTuE1ff0E1obkSmjahG32cd
Mj5+kkv2FL1+LQtRb2rI1IMSpc8y06q8JWaQOLv5t7Sl/3NCbdbuJcBwJdaNBS5w
DI3TXMTG/lCQ8deQaJo7fYtKh+j8WhXH/fiaS8DgCvQ5S1l6qA7YXUXm34gpT7HT
rhELbfqZt5Ql7U4ro5JgGrUttpa5Z2nkSzT4DNxDyz2vfIxjyx3IR41MRrC11+t7
Y5Wvz1jkiEVOGy+4lm9Ocpf0nxOjDlPrUTY5qTPXcy2Nm1VRDb/pSQBYq9rA2/RE
o+1QmClxO0qFBTFkytIa3Q6TiRkBcoM+aJjCLpePUkl8DkXvKI0L9++/2wCVIXEr
L7cFDs2Qs/ysgppGXjLa60P8XPdVumAxdGzwPFzufkqrA0DT2l2IRBBhSnqmLzfq
+Y8CCaNTfbUWPj3L9x4eDcc6CiwoSa5G0b5xNt6gKy75zDJyx2gHOulp3153/LEE
y5r1zwPJXvWGRq7rrE+P7aKIGYB8FbzbzxlU/7J9Moix46Un0tWlxbZMHe01RgGf
LX+46oLtoQlajM7xRWPGUm7CpSbeEmFlbThjOdERPitAVa0l30pWjFS763A2wIrp
RaRNkq9mseqf7frf6oD+Q9IPnxO4DqqqX2Fq9rQFjeZH2tIyOLEksgEuTXZWfo+9
pJCPox/+h+EuasK1xRgwQsk9LIqFUB93xBihIJbEWXw1a58cez9wMhTj8KHVzYOQ
Q4bLVjvRrYKt9rfGX3GtVhSRA1DB1j5Es/SW0EWYuLHy189x+fq3mFYRmsiWrEga
kF7pl5fFKT5f0U3CMApwY1Vn+b6wrqbw3QyP5/E0cJZNQ1EkM8LZEgxGJyS095o1
UTwyjUJF6GMyK0gIe5QdViCMxcGofuLMh4+kLUIKofregSxRQBOmyki9QEOHswPL
FUgYDqqWMAPiijgW88EqTJAqImAogCLFSZQXyX/a2hzavRs0efUi4rSZbeAiu/ej
GdoTjsZzkBCc5krrsjg5HHu79/8Yv+5awLOETr2aqBNqao39UbVxbrKzm+ld/pIG
m3Nm8dwmOl9u4m5i3njAbEdWkOsGIwteaKubPeO3j46hZSsInPbLWPGsXNbF+e8j
mPyApj3ph8XFvlZgVUsurnAW5Y1IwL6Mul048Jv0IZVZeCDLq8K8khrfZSL4gYQm
cDkOGf4WVcNoVJIiz0qS/PY6Kx3PNNvJtXo0G93Mkp5uB7kG0fn8lqLcrhWaMg2V
xWw1SC5RQU4R98e297VAPmSFI+N0OhXvTVi+Y0qutdmJfFzVaddo8IvTivNGH0LP
wolw5HYHrGoBhJpO+c5QfJ/OWxt8BmJmr/oFIHcTwnk/p8nyeuGzs9VrQczCMHMe
EQgYlRRy0EvSdrNuV4R9B0bKdrIMn77DJwWs+M9PbzxjqbFOUQcyDcaFqyeICY+8
31TSpulMKJ4aT7X4pQUlQ1aJGyS+hla46oQ8odKC+BagVA+7OeK2G+nGvSyrG3DK
nTcVsKEVyijYiXkg/YbjBUhVwSRMAAGx/WT4XUKrAjIbMboEp7ZWj38UwSOVpJ6r
bKwaFR3Yai0YOcRGyyPWbbaZWlaFMrsF/gPacrxj4tlwuPLSW79YYUXrecF4wTOk
+YN9MoEk+oyTid0BISDLz2PYBKytm5gXeLKxFbjfawRK+V/3pvyG3Hf8GK4HmBPY
z+YinLOKTE/s9VNZZADQGk4zGtGDVHkC3hg3NK2l9dS8WYI9fHKGDmYTII69kGX/
xIXOX1/+zwdaGHoaU1e+2LDPsakdfhTfZ+U8xl918BAXh1KO4TTPu6hB4MC9AJGE
KwHe/dnoiECr2567SEt4d9EvplUMY9VnrClrFgZZW21lSPNcxue/P94fRqkQr+85
TGBJOW8NVY8KMX4DsrjhSPGMXWUdNPnEgLkxiQMq8Xf/5aqIYN0PzIBZz2/6HaE6
aVnwAuh0tnB5hFK710/+yYDo7/zvICM9S4d/CnG76e1yrXlEM8sBpnfduEy9u+ml
gfEL7Qm6+heDzFSQFDyreAmvPkqRaGjmJlojEDzELJJH+Ts/dF655FVnXcEKOk2I
QVPHpakQbXtrdf2rQ/ZOHQGLnqXmCjXmomnOWAYZl20Yln+50lHhny8xw7w8xUwu
eJKHuTISjI3TzRe32wd+4d0o/osmQHxZC1R+C1URexFIDy6wvnMFFEpn+ScJPJRP
XkHoDsymGmDBilVrdkQzyHX36VE4yy7gNVXSSW93EI1EcyA/sraE/GNNOO0/Whav
FONdQFMNMTA/PI1sGlsNVw1izBt7ICs7D734qGTx/bt2zYvxN0HK+F+ujHR2AzZw
JOgN5ZY47566Y1D0fWvm4N9J8MvEx2kezhfa/SIwsBxcGOSfzteBnIfJG4CsuNw/
fXbMjbqTJRjfkoOYzXCItN12HAU6Vt4jqgahLbxZUj4qNG3TTFUc6SlPA+DDxp+a
Jkccq70dJFDZNNk3Nz3UWeOdlwzA5SX1bzslpzjm4iVtkGjoaYsbEu2k/n63ysGr
s0mORekTbMNWA+WemeA+j4EVneIOW4LODubQnBXFeDgTfeEdOt1aLmvisUO5L3/c
RI1jPioZDsaKumn+ImSYMsnxYyJxUJZTc0mUgBbooktkrJ1UM846UqW6TjpbqHN+
NoyPzC5wSlymyNnv1ueCf46dz/H56R+zJvdqgP5Z0/tKAkyvP6Y5jZot+fuBGHa1
ty9nkKzGZt1Dy64lJxjstOAzOX2zpFFGWKQ5kGp0gq2YPCj7QFqW2ByaUJLnj+WR
VxtieXVVr/5x3xC6181/S1n7v6/RAJPim9u11gazBvnA8hk23J9JRvwcb6jQhRMm
cAh+isefdpQ/Rv/MxWN2qxaPw1ZVLLDsQJZ/joZ3UoCKsDgoJ2eTc9Tz2QxMDZ9G
+huGS/45agWlfkvRwNi+GRrEbTcZd+eiaG2J1QIVv+xE/vi++FHmoMZdKmevNDIq
SgXsVtvxlqFV69DJCbZKt5vPYFRUxNg+mkqc70HxeRfKbjyrbDgeeqEwHbPiRZbX
/NT8RfdH7USiC69PP1yQfDWxl3tnMMASATelaQlCNwTpiFBQjGandBZsjsYUs9GW
o3yGwNdADmL5mnXbsnMgoh3vd9dPjepAkgvkVVmo0GE9DJ3dQQYhQucr+bn7D26S
34eESTU6glpfjH1Pjn7f0wJeQCSQ7lNpVXUfPw16pr++NJqk+dNoKZTZyWkLR4xb
XIYFAdV5ono8/t3cOh80H4C/Up/7vF0bJctk7Nir4xcN2m0UCqJ5LptEgruX/BcC
ci/y9ekQ/lz4wn9get3Lh3O+GRas0d4w10Teqz274ucGoH6PIRN7qwR1UTNRObzA
WRbS3QTLkm1tVyXCZHTxwfenfXLdjBJ8DP9QCzES3Hw5JFp9ev9uQZUqAj6s20Y4
PTiHlfxDBcVtR4ll+7WP5llo1EYDGFQOq5Y5Sw+3j5TjtTF1Vx8C3jAYfegRGlyT
K2r8GmtOsMwAn5waGNde3Z5yky+V7pDxdnN56zgCLMqHQDEnEjGmYc27wzsxYG3x
ZfR3eVEgSdgn4pcHHLM+OQu2m0TnZ+1H92i8fMkbJvrsJWBP3UfKlONLx/qPOtXg
kfbKeqDwMpVLjLyHUlwBdB0+BKHjjdR1fXia90Mz3MPzkcT8rXPsYow3E+DC91mU
IzxFW5+obCUq+9kr3bkQ9TFM6ufkFfxX0FiSkHjl7ou4YOfn8jssa1VZA7CNpK60
8qb8W3Bc23YPepFnGihZoyF8GQWbXi3PHWye+ue0kgDI+RVkaT36NKFYEhUKRs9E
r4Vfvqe5qecsWNkN+stQgO6n7ijNz1LJ9Ay1L08FLrUlRvX5fwRTiLrp5QuJD2fa
lYDC2cAIyXQ9G3FaOj5Ed82cWwOQmjCSJRFLFZSreSR98O2W1Zb5eGrO+vnleG2h
MNRkTfDHlgrVyNpsUCouHK8lKfdsSmXrfwThXKm7wOF/DCJpw4WRT+Y43d0/ILXN
5/thuUY1HvV9KOwNdhoWtHgkRr2IQk1jqseQfvd5VmhjOiZfUD/wOlelDQDoKRrH
FdAWIWIPsTFsVhiRZM24X5W3dB3jkA14YkcaIzKzi/lKsEwK9b/4+COR7ScLP7YS
fB/i19aW1VVZlfH20udBqvq2lb4Z6DB7xXKLkmJzG/2a60Y9aV8vTurtmGjioXDr
8wvJbVtAkt1CdesrS7wEeSXV4fog6N2wt9Hii3Xp0gr9xck7cvUNrZj0tGJtPpvI
ohI09CP9z80rpLwvQxtDWdfkYYLtlQsIcfVgOPJLWIZ9hZaIHvrLJWphxlNoVVIj
eHXMpnQLrtZ1MPBTNpaD/N1cSS8NByizuBfq8FaOvjFBZQBpFeTws1WEtEzaH4OB
K82XcI7Mkq3VN7xS7/QGHgY7mN7hFUnWp+gYokgOyml4mPuwcQXVV/g2ShxV9Frz
CerwoUIurpHlK4JL22KR8TcQOKFJaUIKG/XkfUiCS1vBv1CCaHNSR0B/Y1pm3cWu
LWjwYcBaqcihtWvCZg3SXzA7Y5ntjMfR9GL2WshSa1QVP+wXwqyDhEReBKa5HA1Q
zisp0e+wehLLlYXMxQMAuORHpWPtXt7fh+Q0K0yUnO3ozMkSpdz2G8XcLXafvOad
7kKaFH06EEz3/vyW2qMTD255tYuPzQzxc88LB3mYWX7hfv0XV3zuHfAfiCdAiCvt
hHHz8F2/HNkhYYOxsS3e756CYTo+go1ThhV02n68iXrm4Vi31UFEHLbGlF7zicMi
j5PUFPetu4NigOiHss1Jo0oB8tB4EMqeN+ji0hl6hfWKLk/vroZxyZ7z0DARJHJg
O12I9fxk8RT58v1q3FT+T5I35yIOt2qAK1FrtShe6by+VUci3TzaXxDFFVRLVPrU
94HIGnNLso5BPbL4kUzMKwPLCw0MqwXHa6rdW+x6kzuvrBJ1eO07LKbmu1lRAPVZ
N8bCl0mR15K99WnoZAIhPxBmW+4RAP+h+il1EuMyYb9NoO56uC0xjehZIJB+FPA+
zw+zqMj1tGQwtc2kQh87ibyc7PJ1AcE06i5YMTWOXFloXgWKsuSm1aEe7ak7T7TW
VjwmZqeb2RMNGv1q77igtCJ4oBu+c4NTyUdjE5h/7u8NPRGarwiiBBmJewi6cEa4
Mg8t83KUlf6yKuw82GR6yNXhlRA257MgJiEC7AhY6X37V0F0jpENICyV4ZeBqO99
SgKwzZjned+PFgcpmPlkMiUm2/EHO9ZvJw1jn/bWjbBD4HaGhGOBqNAXwVrtRNkc
ip5l8VAkRhPwUC5tGjPNn2ljLMRkoBVyicTlBPYehyvc5FtUDINiDlyuMs6OmWLw
LVC5EGu/WRr11CAyNOpZz41G8JpBIPI3vqe46lkEF4EUFDZgAjn0BwZX8oFvSla7
RNOGK9ogpo9wk1hG9IzDEnbgBC2Z52WSTp7f+oXWO56QiuomZDSqAn8xUFV5ZaXh
e4bMy/X3PX4CoJFGECsfaVlLvpbZfzt8F0iMiKHQucAGZyFl1ikr3V5JxRdAAR0r
xHXCOEMzfbKMxI99cdBTn3HxSoo9e8wEaGrc5ac9S7bpKMtGwwRhg4mPHkgJBOV5
/RY27OIoKpqoVuuPR+t0g3UE/Mbdh64xd+LETyhjm7LhnoucxG6n4PbhEKz/K6aH
5cw1JLpSSj7qMmsKCNczPxb+VsnO9N+i+teIn200llMxuLWEo1h5StHDQ2X7bTHh
4Dj6eDw9P2euRFWzIKGYw0v6dvs4Y0moam9ZP4+w4I5LEnM/41hI2vm7IpgZEL8F
gfIG/eB1O3ZQ6orfLFgOQVkO+c9/35mT10zPabeAZtRvOJW5oCrDpNawT1X8RTIJ
xcCX//wei+zuQuJKIljYQLZgMfuZlScZdNBmCA4j/npld4GMGMUZPaci+sZorYvD
hGsxKZR+F6JaGbJbHYXLO9mShOD6Jhtl57DHlRIyFsacoIUtijbOcRcGtG20SGkQ
AIV8Zg8ovPKW0ooZEeOmH/hUX/Z7BQXAFGikC1LzZqt1UPKDV0zCLg16dhuJpVVW
JwGjyoC1Op/kdDonTEkaJAH+NG+nUnacJ2JgPQmjcRpOC16HJkkvhXPhCu47MXtO
MFpr+a+l1fgIAO/vBVaoCISMasPUU4W5LaMsAeKsquJ+tWvsYlT7ZjcXqBuWFBjG
lGxu/lPjMNhE0gONSG5NhjlpqntJsHq9/u07lHvPIn4Sg/GB0ZcWxL0RknmIYM3H
DOUpjA2MefJPnbuTmn3CqPO+vTDgWvMkjExf+yO48nYVSbevUSnts5T6Pszq164V
BeNzvWulsPFrARxCkU4QUQQEAXegaRlKJKPIX8NGLLm96X0ndJ+OvwyYzr7Mxq5H
Xpxki+3NZUysFLgSmj/9GzcjM55M8keY+hJ3tLU2KGe30cpbIs27SVjAceJvxDaE
GV1ZS7DdJtavfA70hkuOFPMpZNwiqkoRYj0XEqfmPnB4sUeC5nPd5xeDKSwVbnIk
f56jzUQmh7yyOaBhA3Pe59nTiKJg1B/w/dDeZfoD/oEtj7x9Cx72D2b+Z5IdNtEO
2nFH7uecmgEwvSRqyVSNl6mW40eHjaeM9iAIZ3AdoYuxelB4diilsm6Ck8qKLmRH
yNXmPWJjvLqmJT8/sM1DOmHNftFud9HhZHXPWKxCU+AA87zBDobh14pLRaKCOoaA
jKnAPl57HTXO1RH5Ln39C80IhFnxCjWnX5nZVUgBRa8IAmUm5IPneI4Zax/UWP+m
3GtsSYOKXUPvOhGm29BpkB9XoyahlBIsiq6m6R8SgEGa6Fdj8aWBbE+scKe3DqjB
tiYRl+AWQFjScOoMjIliBuiUpo984iCczB5ELc2qTNIxFRO/OJ86VQcqD/pHdjGs
YZQpuEMwTtOxlEoGwgLv+Iz2wQno4Mz6qVbks2eRcmFYFFFjipGiyxJex1jwE3Di
M8IiqCOBRTBG+sa/6PIZL3YQzn97dopNfAEOIKWkv9T/CcoAI74Edg6X6364IPTI
lwjefkRhh8JgC0K299aFFtSBosQnwAKmur9FjQrQ7bCeNP17jV37roIDso63JoSt
KG+REWx4B47aOd4nz/ExLGKraBdLRcaR+neg8RK7fXL9bRizaSfAtLkk1WdgRr19
qiE0kXpfzCPpRhFvXzr/+VvYwP5UYlfmSdvI5KOPQ1zxbsSjW03623/9aPQpdGyI
Tr1SkjbHuWbp+FrsGHam+uOBhGpCxSTp5GlYrg1T8DPsQJGeKY+jkXB/vor1iGb6
2BlrDRsaO6XJEt5GBLnIxD+mKq/Q7G1xpdvH1TinsjYIpSFkmRyjmyMidKT9xqf9
HO8gphNhl4yt3cZovibvW69UjXIBjpi/+eTBz8i6IWjksQRqvW4EcCakD+DOyks5
RX7rrVxUU3yVooOelU6LMuykcPkifO8tH3iB7cuhGcNM8i8DqzfOmZ4jcezCyPtL
3Mo9PbSgDwvPYNYAd69ZM3xicIWIkPvqO8DPOONEyPgnD9B0K09fHtFo18ylhYG1
chFA5XWEPnQqHHvuUDDeLhTHSgp/Ry/aIRvaPQa0pOUVfc5WiRMVzxtZmwF+4B5w
PFmGJ9MQe+jwF2Zp364WJi3Fn5q468oT+17lNtqzQ8Hi5ffdnwNk1BJ6usLC8o8K
J1haaLJdL9mVvSPpXf7mAFrgbKhDYImH3QuUBc7Sq6tjcYqN/Xb75WJhF6ewVPfx
mrVt3JblWlm0B8V5WB78lOpINypNBnYUz6vH+c4RUopgGYeaMrcytRTpZeZnN+jC
rxPtxyJ1n40Uy1T40sOAv0XWAiZnoVX+IWSq69NnF8XQOJCJdFWaE6P4PNoIXU15
PVPqMA93gd/PxNDrpaAEL8k5+umsNBBCbtEwABFEm/uPQv2jaI8AF326YWTAlBZi
WqE3v44iH1+c0BDC9PtamrzMf9CWDzf9Jm+1giaX7M6LACZLHFmks6412qMt+YCb
HmwkynJFnSlxFJEZDv8eIU6sQ6c286+X6guXrq+zyAGY7p5qA4OiTsX8uDkcUDLz
qCRRNJDYuh42lISW80BBLBg36++kgZTYgrmUKg8wu863l4Ucr+QV1WT4QxPp6yV4
nnLGyV3oSB+SCnQ1onOzvQszz71z0S7Rk+2bHyhiUuOG+qar1rA5xkoWlUZzJRUH
eCrje0bUlhoICXWg/4OOcoU7J+5YJ23tofGthsXCFa8QAlDuvwX7Vaalw4iuVbT9
mz2thEvKZ9jt3/zH6P1yMvMbzLW5+CC18BpW0gIjNOsS2fFQO6TZhsAEC3Rovtha
Stk1W0SPcXVisUdMYg6rmnCfizs43fxzRVspKw2/ykH+r2+GyT0+fExEw4a3Ok3q
Z5qu02sIW8H1f0FwfGIl3v2RWhrugR6LYxKSntEhnbjxFKfqyAKIIaxyqbjsES4C
OT1wTQvPTGX28qDaDjpwI+3ZSLBRKq7Pa1FcDDW4kieM/h3Rl7rdsc6aSg90Ho9m
IqWPUTXce0mRjNrSESn/+OxvIpuVvpZFIY11I1W+gpm3bQ3PLKMSA0JysPdOlCsi
9JcjnAkbs1RkDztOUnwBrxJl06soeM9JHO2AW/5ynaDZmzJS6dZ9xvnVP+VEApOV
jKAFgrT/hB52YfexCK/Eyg1zarZxcx9FiJSToBkiNn+NVOYzvaUcjiaCYN+vY1EH
J0eXsPINpEABu7YM4k4vrPGbKnvWD1XSznuEcp1i8I6Fsg8+1o3MxbTeJtiv94kG
jWFdQXA+z9Cu4XU07PmM9mplEF43+SVd2SJcKYVcXVzcy64z1PlWxZ2GANSHwkMK
jSOJ+A13vnqqi/Lx44JOuYbevUlS9D5Yv9SBPElnJ2PRBfZIF1ppJb0ZVCPuL8Ga
m+CckbHrymwffzsYeFcDl6YqRW8++qfkvFCu5rfp9Sp9YivLczNzrHXDtQcokAlT
pREBQLc4he5QNuQFpI/mXQEfbvy2561YdbUFnLql1db+IJ+xDK3il47pqelXFYQ4
PTnQaPDG3RyUFqoBbrsOT+PlXaLwqbLJ5snG4tn3pzhd2UXkvb08Vdextors8t47
b3E8es7XnPGI4mPEoyh+fN2L866Yoh6e1eastC9bF1/NcZgq56J22YMc+rxLNZMS
Pk/8JxN6yqLZyUv9dKs5mpajmlfz9ooI4AqI2hMBoAWP3pCvLKT1e2WtElU67l+b
8ek6W3T7xt7ioQl84gwWkthTolwHKyDOHIn0OtTBRThWT9Rxv8x4qFcaFNym5W9C
W0HuIysw1tqwK9evAgkES+oybNYZfEs4ucwU6NAOHOEEIn/bRIva99Ag7b2UQkXl
esWKtzM8puHymwrKMPman5uMqyDTcGTlxM42Ap4kXB6vdf+ubiXf+9pFTOCxXbu+
DszfNjGMLWfkX1jdnu3x40H6Y1LWRgfW9kfBIpgQ1oMcxm+TC5Mx5CL3TC/5pUB7
50aE5bKnbrmsTAEd648dQvhls55rROoFUJm5JJqmEiS6I5R3RniQayc+wUupsxZu
20bQr0slWYbytTCLRl1Zsc2AcaTbMK/2n1LHGhbjEdpzUHfT8JClh8EJj1+xQLzV
J5oIh0bAmRrcsKYahocp+c3Pghm90mkFpiTlTdO9uxYtEEjYfo+zM3hI4SR3nBUo
Z7SJkhDtEVkToiSRXmiBkXzmCyHp+hFAgOs3bivdShUTq4Mxn3DxZTwUFWjYa06v
qyWuWRc4KcQthUsowd/1XyMYaqnFxARkEJHJlA1KgcRjeNrEpCYhgRNSSL3hntFR
3XqK8nf1APoeKu/elRSI9tt7x/EcFirLSCu7HFokRbDdO4YE4HI4Exdi+/HvOwlK
K/e7dQhv7YC6AN+MNeF8HWnVxWOPsWXWrXSqWYlAFrMd8sxMhl+eO85wJPrPgHKf
xuCj/qffs1cePCV7cOeyULeZDqu7YmAnlepxEunDoIJJSHSmh7BjCqqcJtLAYfKX
U04lkLREl++ceTszS0JaXZXCY2w+ipUtoE+FICUqlVyy7LKbH2byy4USrMMzsVqJ
TTJy5e2yI3Oh1NYLXksmh14/ceeSiQYf1EZgYG0YkyldcJpLd1ZKN+NHttqf7Fn4
57vDKmLFb5VL26Mxw4r/oYLmg+0Vb8qa4B2ggRimfhlKwkq2PAZMjEjAWXLJKytF
oBJAOSSIz6tA2cSpmEeWEKYouXgSycdU58EDlo4iLMVrQ34np9t3lVuMM/xleJ/m
kbtc9pTuYNTiY2vcoZ49fbHXRH+/5Zp4tI6qjQAfMpfmh8ieFOBwq9GnhzAtxyvV
NZjdDoQSCNd6J07TZR1wjt38suTbc9uQDsR6HXIspV/5DcBrTcYKK40rAkAuTW10
XnyN0xbA85EOZmT2UlHE1DWXub8N1sc8DddFDbbEDl66yldqvQb4VXPmXkczFg2H
n/xAH2eSANvMuGDlA8hFrn2mmOCFoeKAwRPb0mEmE5L/sx2mfx/hVkz34OFLdZ3N
I4hcgntJOEvthehCcKVF43n1fDQZCRnlrZH4fjbd3VMa2Lbh0Gsd+lnvBYCOxBnG
mQFIzgkidPBZSqIt3jsQdDSSowVvuyVjQC/xeN+LGusqAmCa87XkeHSkqFGcWEOy
H1Bkc4KjWt2uwyJX2/7bUchXHjiIpc/EjGzMwJjmFpLhBXedNZ+mzXeERHOxqNHA
w4JRFfHk4EWjX/F/Dd//NUQOv+OLMCSAPUVBFVQHJTMyhgvnX7/9nHacuYRRuq33
0lW8GBu/o/bhpjkwGsCIgEk5d6kwUCG9YlEmVefbgeBYKGvup0Lj7wvfG27yJNJB
+D9F46mdQJ5dpxu86APMf0N87WrnxKS7Q96lwCLyiPvzHIG8odfuOCNMaSfL7s5o
fpQi9TwpmykmqS5e1WEJYcsiF+Q/cZ3jR5UmJD8WZTufRF30PU8ZmD+vNT4g7uw9
hJfaptio5CwA3m2P9/Yt6zg6Ab1BlAlG6PCYchh8RSle8exJZEnazqtwbPxuWTAa
12L+SEqcTU3NwJjQXNJJ6VhLRNK00uLLw8C8EnXIY7qANmJc8tc1pdaWuETBiNLg
/fJ5CtqYUPrk+TRND5imilwu5fRsrSoZasVnC9CTThmTZcfVuzspthP1J6QxU2xB
XzoclsJyHqheMO2aySrAp/MWjpE62u00SoNL0La8p4YwmyxjZaewQxCJPDv5DVHX
jGMpSDC/7ac9bFIrdoXPJfWzQ55utETK2LB3MNualD4MuJ1t37AFAIysChDMs7kv
8aGxV/g+Uk30YfcWQuvUPxrw19Km1yggbk4Rh/M21hsQWTfZRFsNxp8+b29Vezc7
HPfHw6SVSxrED1tzut/JcKtRxRpmne+mRkm+um3y0XOa+tTzTIrqaxZQkq9P+VrY
PFJM+mJWlEls7kwXyg0iIFcVN3Kk9pHtuk2p7++kleSN9r9EsLHu2XZT1NoaOBJ5
+f1gQ9PgZH5UXcZbvx3ciX06jlBucc7W1NgTcn1YtRsgvDETtpeDqyhBRvgrJwO3
xvduhsSFhnFVNvetXD2A7EWJ06sI3ngfngeOdMY4j7S4xEmUuotU/zA2qgG0CBMc
3Svbe+aOe79K6d+OWd+6Kusaaneh1/Or0dY3q4Pc4MAT6VDxEXujOf0wDxzJPyyX
CIY8nX+HjLvq/FLO43pXKkdJJtSpEw2EqJtZbVcGh0++yw5DUb2l4B6vcToxAa7t
n09yTLB5ZbqjrqUAxP1MqVthom6SG1lW8FgR1PKA6BDhZn0zl+XOqHxe0ep8AMan
dtT1kd38W/FZJnjihey52V1Yst+LKoa6JPcQEeY7/ZfMNetybJhp1hOx+9DkPEu1
aCnkZl5YUWuN191c5VprEyrUJdbo0ojoIgCH9bkUKYbJ0W09NWA6ybaYqhoffHCN
ijQns88HkNX+KwloStuyliqsLIZQfqf9RPYVA/FkBu3DOnHrAgGKXpfUJjwUcrb8
maGqEa2LZ0u5y45oGqeEGaa30dkyQ3YM9ku5AeJAT2ik0K84qwI6QtOfPi07gkip
U7h97OyfVIQRtH2oOpjOifsn/M0TjX+728aMkTl9kzOomB0hhlDUeFr9a8LsODIu
98tP9xwPNxdRoPLYAvi89TxopmVuj52xUvU9liGBuJnWpQEceX2I9FeBe7rjfjn4
IbtdFRhbVKLF8Z7zydJxWvV4xRXvcMSPzIPL8vfQNcWHWRDoOJcyTX4ILbhu6lJV
idRhi1A8xvKPRRJ9uJCNoN+57UCvpXcj4EPcz4u6bZ7slwQ5SNAvU5G3M5lIh0Wv
b6LnswGsZO4ts6qX6DRt2XZ9Z9xarf+KvRgBQhPvwaCMtRyWoXgR/VBIcve8t+Aa
TUgtukhcG/lFul5mjAB6213KFoWoDmYosOkf0qL8dp/Iv+mDfjkovHqF3Bmt5Il9
eNoz9ccCt784ukzBFw2hAWCE1Ofrk/dqYn+3ed4Nkd4GZBpwKAPnOszvkA8x5dwC
xqt2QviX0kuvW52xtlNz60SLNK0HuFGpp1/eQyzrflHc4d4yK12ypEINx8cWwVUx
/0IaOxDgneJryKp0rlKhjo1dyWftyEhzhYFhuXFREEtKuf89AtakmC73Kds94EbD
GklSylaxr2HNhxDhIHsTqRUz7uxyCezv+HCvlec+mQ5OpRPtxrf17pV+McUrWZ3E
660kIy3HdRyCYhuFPCpjHUJoIWDBnp4H3evCsKgveoKs0SetewA0lS75Cpte7EyC
tA/j+9ayQOu6ga8tVyqr+6PRvgrdxw/OcsEcZqboxIbppST9Hva6QezaYnuyO2kg
fpZvXLunrEl0K45yVxCaT/zTL1RRbu5mFZ63nOQrXTTS+H59icOeuXkmHtw6KW3Z
34MG5KRHIExRuqL5p84CRv8yal+/uAvmRTC2UnHj/K41zesLYTloOqYFpzxzPnf6
jUXa0Dn6jGFHMtGo/L0D7+BjdaIkn5MH6iNE9BzK5wEgz27t+LugecItB/O07gB6
WNFTiLwKA+WJFMiF1P5SLJHG1C6I1wmv46hSE6Ro4kX4lFm9p91fMHwlKHpaVnIw
4qLxiso6EsMw23UncKkLy3gOXXpnpY4HtBoY3IPa4KGedHv39l+3P50Jjk/2nqVI
s3J7DsGcN7CvkMK3//HsorI8mi7kNkh7x7KDJxLyM7a+WU/Vlcjdz8gxAZiimebT
EledVoMkhkKaHNaea9H3qAzy3OGn7zLYUePHjIgCALr7VzJfd2n3Xye0B3ZRC2Yf
ZL3BcBBMNJNo5NpONRjN9XGqnvC6Qk2mCOpkK/3VbeX1MsIWnZcGkWDMy4Hyb3Sv
h7q08Siy0jd6mnUzskQgPuVF4BvAGiEwlggUYGXv5Rz31HLMWh84SxrruJd4VqZZ
zXJmR8dSxskmHL5AJeHjP1Hi6rP/bPwKHaULB+dUGQF1JpJffMyE6Ecdv0usr6i2
kVGyrEIU2W15ED4KHrP6a0+MHDhyor5zYR92KrjxuKFmqeDfW9g3oJx86QcXjJEV
aQ54ycqK0o460D63facYq6jo2Zvg0Mra4bhVeKZHSlZqkspKGjLHo4wWCgG9BphE
WQnrDzVik0PvSGBRZinOcUH2tw1f8mhMobMhcCqQbdq9O//WMup7DNrDrmKlwew4
R4FFu7tksumUN24C4CphHJ8rJcgcpb573frFVc58Co2PFjorV64iQJENBSZLH+P7
7cYDxIBV/ogXcKf/z09UgqFRHncdQZ/otVz5qomDvkriuOjHsL2uJ3gcJ6Et2V3l
ceoGnzm898vvnYNCNiJC7sTnk4QP2ieDLipyZI7f96sVbXVyb7ueb1REDruD/ijo
koQzwxVmYzyhMydwD/KWqn4oyZU+AY739fY9+qkLLdcdKlApK+xbo7nMe6DGwOyU
5bNiiv2rg0aDy6vATNoms+MRYYW3+tk1i3tRrhqK7NT8NeEQ7AZGoZUtBrGOjqcu
V5DpGmtUmCPzxtDvTiB6qRg+ZEJOp+cy2VhTTxO/1Pti+dEd8nlUFx8Tnf6U2TTy
wmSaNpZ7aCA2LO8/+J3zO66gIN4QJyO2sRC2AHsTi2s5sGC8pQIAybuLyWZRS02Z
rMJopilSllBgjbF9qCLYiIeQI2D6ytmzkwFgIjTcENxtr7a+kmZHMmujve7NEdWd
9UAs9DsdB3GibwlEaM165hJVH/3Yu1LJ97KPJUVL2Hg4RoPAaLTQl1MOV7dZzbmc
WPd7psE3vRkYs7fiLiQWsPo5JQp/YtJjdWesaQQEMNclgiInvlpf5DFG/VbtVKup
h7z7Vsd80QiBhPbWxG/M6N/Cx3ucb2Ml3w3GtV6exUQ69oN3cgU5Q+yhQgzw926d
EB2OrT3TG7a67uvH1dc7E7JJjR0gdK0vBWSbw8YRwQZqZQPQYUyBexazuiKRAzpH
y19aJStXnK4Q8vkCMnknv+NNSmlEvwqJfF1JXLwgOXuTPMCmHhzNRouChzwVn1W9
B9/TqTBsYOP8xyid43IdXxCsE1kAqAJ1eij0/jCNv48no1FnDEFTCcjYy5KZPaY1
kG4rxBqTpiovRHqOT/nRKXUTqjlLPMnJNF1jiqz5ZiKkf6xdbY6g55wjgzbwjgSH
NPo+AeWfOD611iMaXmBiS5Na8KBtoAUB/fGbAYFCt2sk9IHjIDbNMwHikiQaMOyz
zSmOVGNHDV5nsC7vnL9ZeAMqeHi/k/c0W5dslGnvGAaK9/xFCot+0xvLBBk5kgUE
7kSa3R+hozgDqlOo6ECKi/IIe2NrPCVbzxLyK+r3JWANzkuE3UPJ1IBSvWMU7k1n
+fGKRWkDj9QadbSDoZ/4DdTMv+Qus3iYIU2hTiSDNlbOLHBZ4nMeYDTbsD8z8Zhb
DFjO+zxROn+MqXn+WdMgCgRq69lQE/9AJh/LC1EYAs9iNRjpnyBOezxIkHX+ZGXj
qN5MxMvktHlRx09vGsr0CAR7TSItZeqnICl4/C3F4czkxJsp4JLIxXMrTwYkSaJn
4TQ5VLNn4YAiaYccDejWuiQKF77Sc1+J7iRTLU4E/NAjA/j7R3B0e1I/EEFXMQXW
eu/IhVNSxNEdb+H+Sm/3/2RvY16iqdoS4G06qmqJnDvsoySuEaP3EwCXt2uaY0XQ
smGaYC1e/69dGst8lHk2CAM+pYn+lQ3HtltlPh61FpM94nlbCxJMeMriEG9AU0xn
I6g16cvZdS2d2l0XYRtMTjvgp8FU4TM+DZawhQvsgSvWTwqAF1gvgbXFkYKACWo0
3odbizWCPsZNA4llzZq3oMhErcEkLDMZYjFs4qtFjUD66PUI6fSDe0ZKxdnLd8vP
ui80In6e+Nrqj+IkNpyHGnoB5XSj+eacjYx6WCjIKczAFQfr5jPql1vXSF93PLho
VPXFHy3t/tNwu1dpQ8n1r92X6GQN3JM/Y5IxG8eJRkfWuy55yyWMmdSYJb3Zo+th
dVGNuHB0Pgd3ioG6mBaYA/A23knB0aqqc1qHg/gmlxgrOXuyDDoLms8VLhaV/JOR
5g5xDS58A443Jy6jhFTgPIPvSaQMAty9YCFo8Af9tAUTIt8nSYbuZztOVAuzog7E
wUd3FFRdnlm1lp4xw0G/zebbPgVDbBmymABvmx8wUfOC5/fhdpUh2zH40aaWZila
LX4/yVaUBAKfgzueuZzNN1jnwrf+tomjQ9YXIgyZcEwt7QErUUQ2vMnYZo8MHdMp
sxJBo9UoWQ7+alsZZx6GuF3eEkfKqkfCSLGKNtcwJToXu6ZFpUVe+/NIcHUxjBtx
deyVTrwipP91+V4cqkZUuupzc3OCim3D7w9GgGWD0razjtZYDfN7g5NqRFdZvIkS
XiEV+RgbASqQQL++2RJhYueUbfbA2y+jVxN3Bq1RyA/auIqrD79ixeESAWAlEmnb
i/PMLb4Bmj6Lmqd5xAjuQOHHQo3FX4g1Ntz7JTp680qswc6sH4tFhfHVq+K5CTVJ
jBB0pr37JSErS+9kNnLSCvqpd80IxMEZjxt+E98eCf7zhZziGSUeW20bGwR1f44N
54kNZRR6s44opE4srENZ2oWadjjdMu6NL/Erosn6mRJkbcmWhTUKnWNyS/tVawmY
kk23hgG4oDCsWldRNGsc+PWqwFeUEJD/ET178sh6AapOjwO95EBizQ5hYx2rUPSc
skx/iUGOnf+gsLCXKkJt+wGXE06pJJHj6WrvLyrfdnbjAaSyarilohG7Mp7uXkMs
ukN5wtaKqI8csQJfg67atEPkDlyPcCHcRT+8g1/YcAxLbRHyR1xV3Rhc0mSdtNwx
tRFeb7uD+4brLdFG7JpxJdtJ3o2fa23BPx1QfFXIMCH2MDWR5i/8NrBEajcNFJn0
BiSulZNPwoWSmOtHOdmG1HQ0kt7qQn/gVs/hqcZ6OxRowf38LtWUIwK7TDq9jHDz
Al45jrMz6Wmlp3Yfle/VmITu13oTxHzL+lEI16qyLc6QCSm03S4Y+u3+qi8XeWpv
kWnvqe9RMJtsHWPhfyp1VA+wziF2xBvMxPdL1LrdaWzI6BxW+xB35ZRfoNjIVw/6
yGLeXe1DjsN3vLuojF1J+M+NCrbVYP+PDI9wThhf1Hv5esHa1K/rSMql+uykFRjf
N83dPeybU7UUHJMgGWicAv1B5fV4MeT//LCridkHEhZL4RBrcgJJHiCLhwVeVUnM
paLfNpq//mhzwsxDXHxvfgIV170C8qXncvEXe8LLtSq9z7jwvANeh+GO3PqipnAN
ygj+VJZRAFHCKc0EUJcV1kPpNXl38PqjZ3ztS0/nHPTCxdYcUAz246qRJBS1pZQd
mqHEOTDogY7zPvkZIXhrFLJvZZh+8KUOsoFTMp+nvnZ9POM8rhpsqvrNLtBzupzP
r+el6Z7y54m1LFnsR1rG9U9ZqDJohhOz/vjGedKL/fjzqK43gCA6JZmJ5DtS46cP
wIOSk6mylKaFs6u3KKPp4kTeAdBgZ4F6/Oygl8b9mfx+1D+Kxl4RWJ8aUtcjqM7V
gH4ikuRd8uH4lbi7Y3TsXfWVS38ca93c5BywJKM383Kv36+rOCbFgJQwgPQkjSkD
B7qbIpcykntoxWZ8HOlkB9ylPE8QHUnRhWmJVtqKrQs9PyGixDII6x7A3vaRDlit
shDQh5V0hA9gmDxnvltVtS9WrdcG0vRnZyiIXIcuapKY3hQH5eI3bFeYdL9Q40CZ
iELQkpuJEpbOfT0K8bfign3rham167DLwRprdS97kBpEpEeEyTSnhqJ57fdAkA9k
dzItjbS+19Pdw6aewh3b7PXg3xePda1rNmRP7hl75IeyO3I/hGLcJj/a3QlRuHSr
ul82QsmGPDO1RfR4gRQaCyrDyG+/dpQRtIFAisojx8njt4o+b3QUbhsRmBFCiShX
a1NwxD2rCvCgFAAb+pg62oQef/5SpHoacWG0diKCY1L2gKY0MwPz8xRyWEeGQNCx
98BPRuQR0KxVVtqSxjZ2rxTdb1eWCcg7/i0PfPb+ZIDedlHFe7FliXxBQpkt3fJ1
TSdYWusxz4U32K5RFBcnwKCi269JjgKYZE8wp6OoQd243TgHjzRd8WI6+B61/M67
05eRd36VaAOBZyfHY7TG/XxPzu7coF59wYMy6UzKJeQX3pmYUnWtzjJmbhm/MfnH
V4jsr+S6CgJGJUZ17MDYM2Yyh7lnRsIjV//Cw04CdXPsdRnYDy41jbgpDi/4bDI1
MU8C+UZNmXvbq3yLT8Pkt9aq50bGTyly6t2UhhjRzuX1FUpm/p0gO2sspSlSOjx2
DfsCxYW3/qWWsi2RtDcGzSyA7ZdTD8z9XxvTC3jBAN4rMN+Nm9r5EpNUKf9536J5
G2XWipDHNcp+mugVI/9QpFx8i8rFnX7odl676eTgG1hLVrQLAvvdXwnkBUfTdYf1
/bXEquxUYX/YF+YsilKb/aRmjJ8gsVLkK05d3uo4ynRslhVzOVWprVLDQDP1XoMU
5ZOPnuCyz+6MBuDqKYpRi4TENQRavaUFHl/cZoLbaXivycf1llYbomvb8w3oxl7y
sOSGACGyLZa3Af5PE7adQ4+TKaHhVH08uqMjw59zWM4jJ3ieYPjqj32IMwYq0ZFQ
SHssDeQGVYMjuPWadzn9i+dWIYHRXVylac4ZeGd7oBa+AZFcQktkf3EtWxQHNNXj
mIQkJGinA8r5g0bBMJ7L9iayA0m188pocP6kwCRzWh547bFZm9FwXESCV74QTcfL
LH21xjqh894/sz4/rUcgEMjG0G5Anu4fdGvFvPFnC6czTjrSENPB0gGr0fXP0+nI
PzUYCPIbU3Q9oRp4aF1qoB0y6AY+7rumALNi5V32Cmjj6W2tSIT54jxrqRc1M0FH
h9eXRhb3emsGewFbalx/ucObtzd7mU8FxgnVPjLyOaLDSxVpzcvPihWTz1HVoAkI
BAmSrkHEH587muNiKbvEYbE8O2EmvUzkLhrSDKhLDxd8RzwTuzqdRtiRvh/fZTza
5sVxNOo1xHI/S9YM4UIACYFNu7Kbd33VcfAZ9w0U4O49xg+CXKZcFYxIHmSZZetP
cDnnLHtf9R96PO+zGubhsVo9qOG7YdjVTUwi79ghVl4Qm49S4W0yc/XHxHgFJ23B
uehnzE9tbFsNaNnjEEgdyjDiwAAYitdwGjD1twYYc66GODyO/yKX1pdzHon6/5SM
yT6JBES1mHQlZqoof8YZnB2UArpy8k+/drUwtXs7Y/uodM9TJT076P0YUqyeRNAn
k/9MMQQazEqYGN9v5MK4k07ExbrQSwQ3nxu7/+RlcHlid98tbgfOV8qfxzNMwcnH
Nu4d+Wv7+xqW5Ipxs4dCCf6wYApZuzwpIuzFy3FWud29skMBtVrNcQBhDxPEog2r
k54QOu0VHL33pIzUlmtgBjcV0XwGy7qOgHHACdWknJJRSVUtFTlB3aTK2ckyurvh
KcUgVr61xcy0Cnkxbfk3LtL5vkozKMJl4AuEPGXnhCmwJIn9GP6Nu+NxB+Qd1S83
xrrAFVtfu0sk52z3I6NnIE+TjSxitXBSdzQ6rxEgRdNOfqbCQj0/7YgjjsDm1H15
9laDUhTmX7nJwJ75BvQU5XDhxAIUP0AcZt37EqitVUoMEJ2NegEbV4Rc2WgRltyl
OcoFPCt0on7ae035nXrrSmUXARhKX8oy9HW6pcSKFErM3/6uRruWAKLHtorvNsCt
cUpkPvdSo6WA+5Zld1G5mA8cV/k4gKAdGordm464t2aq6zr+vJ8HSFT1FLA2k5ls
YNVwGWwRgR4JGOPLJRbw+4Pe5805ZJe96QxwsgJNg3OQ9NPj7GjpqA/yVVXuwYH8
3IQNOf/OWr62+v+4fxAPL/tHn/IRNQEtLA2AephcDRlkxhoIcvKCLY9xQoWBCr8C
iad7jsz9vJ8+FL0tb2ezEpS8Mvx+O1EuJJspe3taGZJT8doqtIeQQ6sxTKh1g3Z+
lEa8Lb/BelY6dcBVg+YjN0M4/Z3HOmx5qxjGwNAgX0TM02rcziWTzAddGBg2uBDC
JrvQXaUBLxE/Z9REITGUBoSiB0PqybWbvi2Z7vcEvAPeWBDjVLUE8X5P3Fpo7Iau
ejCvu+Wgxu4f0T6r+tq0Kl9rftOACqI8WK/TdW4NrC15EpV45OQIDquRT2wZN6Qh
cx6QsJy8fERJJwm/lrTE0vLddYOUXJTS/0a1A38Slf1pFX8V1EZniw+fTt+FGPeX
4iWvJcTBi6ACdunSK8Q0obg4VX7er5pUyFyvAriAkkJVdC4yqvzyKQZ6BqM05lC0
4vTgBFdcbKdp2vaEr8mKNKee/qUzDNNzqgrTvkdqUOWmNjC7ssG3+CWt9r+syR1k
4oLQMZtB/B96GdbdGQrtqb3TEI+wydvALjzaP+lxRRa5QZlj/sW+7b6Tc+UFAOZZ
1oEEYmaZfza88fO0P+GErNLsEermtL+xpzpMmPB9JWsuJBO7rlHkT4NMJwdLOI2e
vcFxm/t4boAfuwotxtPOhFVS6OyLAGX8pyBIPl+8YPjjg6Mv9e+TrYsXxy3XxcVx
n/sjfnTY0gqLsUJIbvZ5EDc3DWJOiPO0uOw6Z8Q4AEDx9uiWPINv9gQR17KTPIcz
Z5wveg8Ypwbom5guGJQ2Ju2B5bBKHP3MUna4qiCUUerodTeVaV13MJzIFnxShsnS
wD3oxNvwH/Vt406rMTfXBBGnpQXhG4IcAvjcQxov5oyKRWSswApHnpQowgQOQBDK
wAbiO1XFzLfxfX0D+5V9miPi2nhk7gbNk7SJMR8fcoWoD6fZEqz08uYqM7es5JZi
Vp8fJv3BYE90nAHeJI3dZvNwSVqFh/mQ6b3o5FNEkqxTzKTvO3eohbXX0brHyzYs
zcXUu91oD4e8Ren5PMppOZ4apYitTJJzFQevOJHzSPTQbNzTO4NunFiUq5M+lNJG
tPOT62KEdcex4P8vDvytLDwm/ehw5GOFk4RV9O+/0+sJhwlrinNCsM4r5YkRnNaG
g1NWqi8IHp4sWbaBpC22ERJgmSL7xI0TdcV+AIQP9zHmJCn6P+JC2+rpNii0AsJL
K7efXEiKdlEZrPQaAeuadxDwUM6iosMeWmfUk0iILXKR3/tjYZxWfKXDnaCbL5jt
2KATQ6k0LUimceGFGBuA0bPzCqYXQjWG1kcVm2LMaP6Ii5k81e0oYYuOoY1fwcit
+Jo6gWOxyxkp81Ylatm4YTlXwldA+jte2ESmwDWx+BIWtTKzh+Sps9if9U4QZohc
A95HGMj1bLzmWGButEkctETublQ970bEAPt3I2wD34x+jNaOcFLXr5z2g4FJkj1H
oBEnnXJeGng2VDLnVqzrb001aFA2DjOZ+yFct04ObFRpWYDX5pceF1UxomA+u/vm
kknA6hWlLmnW+fLcG+a5fUHHjP4p7wWuCfnTa+LIRhO5U9wuZgSUMvtI76k/R0Rv
7IStM7ZEIa9OSSFC5taPIX/wtNMA1woasjINWxx6uqXNPqWaicFbJGJM/XMGCa/O
u4cq64HYXA2nZckPUy5y8eSfiRAmjmawYLFpk+pWzR7Nj2u+muuJU+5xJUDAqv4N
QHt5XGBUDUGltiXU2SWa/ZlJexNckyZQDzeN0OtP8KtMLw6HPbAYssfOdabPKnIj
4+If9LbC6qUY76dcehHVlKjd9QB1kp7Ib9hP7+h8yAjRf36laCntxa9Wtc/tvt7P
6Vp7Q1bTRUbut1843BVduLgvNNri4uEMwMuNvXBZ9snKU+j/uuHO3G84Wce5sHDW
2pyH3MyXOKyBQZ+VJ6ii5GpAxfevqStDkthxkC9VvwpfuTuN781AzpQ/odjFKs2R
FkntzqOJXpcwK1/KtsSuG+hd9t+w5dzjJXPpie8Kz1Kh9b/9FcyRni/e9ANd/Mux
fXYRQQG+CWjcZUKtR3cniD0PbxF5xANIduUwaANpSF0wXEdQ2P7j77QQMOQKi4Il
AeYY98LFEBNYcL0+D/f9LX783hQ9bfLnCM77YniHW/xtOfh/1YYBtlY9ySW9uJVV
7zYGr1z3GVP2zGpLdpVDjgzUuhT1PEEltrORZ5GFwlRy2KvujYkQYG1EMc/iwEZh
2rqT4R+rCyHtY4uMG5MPXXry0Pfi3NXPUNfwqR/0Dapwuqp/K2XSVcAEB6vaQHbc
soLXrPeXNIi96mDUaqbDxtqgkdG20YtG4qzu+YT0mnKZX8y+/hgdF9cuJOI8IJow
r9oKZNq7etJjZOemDaAQVCFrN//V2ukIOsf1rwxzLZ+c9poQP10Nz4bgeqBfONyE
9kJUVHXREfJ2alTenQSuTWlAupGjDjP9aBtiJ5ncZ5W0LXoTbElstR0mXNAnHMLF
OYXp8862QRYRETZMrYJoRobsAB77sZHhYKd9rAWJX7QA3rQ6VYAAbVoWsOjo4et3
xvsrnAprbXCwaqefo44/L7OIb2kcUpWX6gIIQQd3drG63bFqCgdQqt2d12oPD7gZ
5TzZGfxCo6WCJDZAT0hOVdEly6g2fmEZr67eDIJVljcepi31C6z6byMy4EgjMSOf
ND5IYLIznf9Z0rAMR2piK86TcEiM9A3gGc+waRlFV2RRwx8UYtyUwDAVPeIZtXUR
eewlvlnHUWDuWjI9h79hh3X3u8jvrOh2OtKBRdZeOpUBdtqiANcB5P/tVPjbKusJ
v2ZkC/Odl3jbkhz2LOuBYu2X3BM+y0s4X2BocZ9iYuxajWJFTyGJ1IzXB4pAcZhS
7KwPnGZbnTRxZ5fVCAJ3DbgycnO85l/os+uCJu+oY/NZCcttFKGmpkfX9rkbKhM2
fCIa5oM8yyw0XlAC0w1nYeGOf67K1APlD07WT681c3OijzV5/lZzJJfEItSGhE8B
0BzgWc4C32bB9ZAsEEgKTvZ2hlVWZo6VvUDO3ew7DTNo/ThRfkC1FE8l1GOgmSfl
4XVbOtRHvB1pigYMaMXaTBorMUsgKvqx+CUaG1d7tQaNnvEQ4cXTXUOK6hb0sIN7
v+ITfF6p4hhZEuee7atqMxHj9dimkKBHegQroD1uS8LM7LIB8cCH6iCNBdiIrxx8
6DyE/fhuy31nAgRoR2z173hj/udzCCrIQla68PZf0xKFSMp+IUr+Pcb8JgXKWApc
ZfVbHJbdHUXQmldih/2Z5cw/QfWkLzCmFDgGhoS+S82p6qjW1njA1zEAm5+TebvD
jLS5KLZquUmHu267Tr36futE12SwND+FdagFmiAwf9nlTMl8Va3gMCxWFpTl8kQt
bmoBGt51Q/oqSm1lYzqWZE5vZKiu3QPjwU1MfjRQada8Mevj8tPRVlAka875cK+4
6htLs1uEmJbordakFVS66UE/nsS12GMVfdTdoHTk0XLsr8fBCHEA7Wq0X6s2e5Ad
wu4qrtH4cVXlPcnN5rWWl7xjUJ3rT9fCd2vGgmIAI+Lp3dek4CdP94rttebfXKJv
8WsURrNyBE8VeLFko0ZU5Wwh6OG35FDjDo3Gcw3nDSYZIkUpVmj2oWYhcwzDmznQ
Na4YSzOBImoQkN2iq8UccSjXM0brxOWxRN1Rlonl9lkynNftrqihxGvY3u3pMRkS
v+8tzFiawoJug283+EOAJlzkajGR9/N7chiGe/VfbVoNl3gRVvc4RfEQ1XRi+tuX
R6J/AEooCe64G8uAcj8/rR3YllcXUF0gJdMmqZRFTBkr99nqkEbwBPn0Ln1SRld+
UpLLP1OP+mW3M3PV2+nxSoF/MUF6hC9udhLM9941t+flsbyiyU8sxxXuFZ27LLsT
TZe/GiISkrpSClWQPa+MVdBkLYaWfWAo+f9lBnxRbLdP83v+v0vMFBTCfg+ab6Qz
J/DRYnQogeHFSFK2NxgZVfL0Rh8a0e7AZsw36bFRSBlplY+GLQ/NsKcg8QxBE+4U
KniPEQ9gMSs49IuA3V9WzYpFZD/MKnTKRySRKl81y/S6YBXI+BmrNnIWxf0wJPsF
EIAITa3HHi7zEOOTRmMsXME6zpAMbCOhoUp3iVrYd1Z8wYNeeBR1T34ZRnOOHyrV
bwVrAbp0oLn1NqnzQMaQyGMKkRgWkUOPoBjxpkzEQifX9ZNNw+Awd6Ieern+ltmT
5b2tp17EI/eQkWz1kHQc8bSuLZfREbUrGQW26VR26rpoX+ZH5cYpLbztb7OEW/g5
g9wcPt0QTm5eloUv/obn7UVIWZTiMytUZVXdoR84dsb0j+D0vAxYo0RIcsLs42w1
r3YN2IrFn3GWK7AFu6ZH7e99cMRULuxjRZbwQozcjyPLNbCV8PBK5o/TvIWMOR+s
8RAJAglK1AvrqVj3LS1qhIFTRDSKyYB5B08yzeYbRxqTjHUAiJ72rq1FKCID+RQX
flAyqKtHckfKW2GD7roWzLNbiKB8T6mZtaS1b6ikC1qInv7sDOVZw9QEcnBxS8NO
iL/oYakuY6GQKG5B9OLNPcIDtq3DVZa+Aor9CmiRXXKG6lfP4ShojZgMFcaO05dT
Wqi0waf+glC9M1hU3A/U5HuJaiga+yHH8rrtiKKYCIthWZAA2P9ypb04Fm4oZ/yP
B1HCL563LEDwpoVxF+xGk9mEXtZjriUlOIEVwqONxsbG2tCdehgLnJ8CgDRmTIys
RvKe+OASFixMikkR4fksUmA2FGtV7wtWub1d7I9vhTetvF0CmXu6KWDVuVYyG6JX
w3V8HoeaK53YkDlcftKbjxUyUfKtcYvrIbLZOFULjeEPi2FgzrXjAJJL5jUK7rES
4Um1hwhWagqBeHiSdQZHnyAWPPZ/Aw4hT7Cn6sCHr+fuBDgfBegd5Qtpeth2YXTf
tkvRBVzuEBaXtE03xzr5kqu9aR3MbZf1G0rKXLHa8Eb7MeKRO2Yr86TAWbAQTTEW
Z4VYdrrHEtsuoVIfdl81f9JAf9OLxwnyxFkdilu8BVxWMuit5POCRUUvEo77kMm+
b6YWKsdKaE7mBeIF1vkszVNk8RPTEamlf+Je+2+AIw7ki8H35zGPE5HSIjCNpR7s
AwIZKg0bRKBYgFOBIfN5e5kCLfiUHBwOJfFp6xlKaO0985JhIQxr6wl58wrtYHXI
jIeVu+lnHNebeywUbfdv4dtS4iJvoJAHq8LqctnUygoL7RjXSev8fFaDpSpclulV
ogRA/V7sUYf9s6ZeANo0emN5P0OkpHSlu1EGpf4VlwKKGF8Q9L+bx5c1Hyv3hR1l
uTZWAsB0Ce4KFBR13J09mvGMvJo9awmTwCNuMsmFtUstqCo+FLwFwwiHDMbkD0K8
/lEvJWfErb9h2atKT0/hozU1aqOeosroaRrY9JriPA5PMNvJd7J1iTMk6h4aDgBD
Z3VWLiHiIFDckb0a0/DIyWiiO+Cq6eFwVzRBIquTvnDVCdI3mcg/w1VmFGk2qWAW
kYuKMyODBKUDaTYf0qhucr9/n6bCMM6pUk0BXBinlFHQLRs90JmyJqJst1DPxE43
KO0/038TqAOpGaB9fvIC27n+AhGJoWb5EyMsM5MS4GQC7Ja3y7hPtBMOkUfIKw8d
F6WepQyx39YoCjMBV6Fv6EDExZlDEAey9KMsC3opTNkf9/aB71nbXIOatAwnjJxA
GCgLYT6R6bq4EUM9HytHYY/wgmLBVM4GnnI+CjR+qKn59IN6ZT0NLhYx8jpqm/fb
BVmmL81Hd+GxVvV2umLhKlzQY2PrifE8MygnqnjBXU2FQ0QiHz7mddGBthgZosfR
ZFHknFS9nPSmK/S98zvYUDlw2yroIhDHJc5AeyYYOH+TmpnKmM9Jf7r1w14RkqcN
35UwImNNig7AqwSUs/iVNUEMmw0k0rx8RdIjaj3NDaMKmkBz3XL2/flZ+BfdtkTg
Qie/sfbG9cA5/UFvyI/y6vfO/LlqWmxIbF+99YP6J52kuIButvcC1LU0aq6xrDiY
c7gJXwACl9VS20LvICoJbExX3Fr9Y/uRe3VMZDsuvtbWNTxF5rdu34KeQSt914C0
5dV2LNE++fcVZVby7qnVeLz9oNuMF/4+QrEGRFrbjoxwd8g1CA8h+idXpa1Q43B9
Cl85PLUfWYtAnEmwMWHljSufjN7NJ8wVX1DdJ/JSEd+TReKenYLfNEHj68Mw8qFv
fmbeUgBYflYRiiF2h7UIziLWE+7oSMZerSYq6giDekFB1k+degpa0jp8aYVxNcd/
tw6C9PlB3KppvmQdFPh065GIE5YIynxU66GqDGXN6jfTJq91SZj0EWPuAcx0NpXD
gWR+kO3IoKgDMKU1CvyvmS7PzSBzBmuJiq2o7KIVJESk9vTJea5ZGX/muiox1j26
Q/xWMbuXISk7aILgeun0TwCuHZp+K8/ZleFok4YrOoGN9UXWsIDmnLSVStueI6Vh
jZSAJyxwg/nyPaOX9afy9AU1IvBjLRDR4OV4tXHDkXiypYwHaxhpX50DH9X+0xSZ
9peJT8dIXJrxhI6Sv+h3S03HKsJdPoVLM0fa78AnBRCXromiK2Rpq3Y8gOM+p+yf
DLBn7rpY9i6iC/z1vUHr7n6D+JxY9SdKrrllee3ZiZD9+xoxRJ38eAoRUA8sKjAj
Uxz439MN5sxj8LlcyS7OQMpXVFL9OwiRR0YLaegzLhK0pEOiiDShMT4ogsev5heL
icACaPWU+cGrXt93z6JsNLKZUzUrDayYIitFBeC+kr1F8+2iMSoLI9BYNW8fh1kq
V35qqhd6ze2j8ojE/R01ZB0J41VUTg8vb790yL5PpPxTeUTUSya2I//z9ZDsHKvW
6dHMDtOPO/B5vaoBPVs5L7Orgo2cVIrphhkyDP7cL/xftnMsHopo+5ICjq+k4gmo
nvyvz8Cjrvu7G8yjra5sJTYoU5OQzgToQbGS4s4gRJ7WUQp2t8DNlOadjLG1mUur
CKLChkYyZx6G8jA6qlwqlL/4NSEGZndjQR65v4B8VF8WUcopUnwIxtCTWD4UGXo2
ZO7owz59h4rzyX4dIlU+GgL+behiNAnTI+/NQ/itfhSDinJ8KQ93aKvlZZ005KdD
VUmYkAqGHTlVJ5sGFeVjzOcXObhS+mG9HTywPT7eTfJKXncLvDYbqnNXdIUNlSXd
L05ZDzoDwT+F9p+x5jDbBIoCJAtf2v4/NwDnnY3qI1QBXkVbWpPT+BNVqcz4uuQs
ZTnqDSEWa9Ff9C3m4M+lzCtdIwIIG6TPBB4lKswD8wmzYUo0bdTP5+NOty4Ncieb
UlpaaGG4tYnzJ/8KlPkSJg8NTiyXLsGjtWJ4Ztv6X9ObzpijhTuH3gcQHCbgnRkN
SSQQONmy1ksxmwMNZlOPqKUntC+WNGG5SkroSHw3qFEd6D/47qUfg8YmanN+IC93
cn91UeLhgyp9cLMQC4+FkAxj0MrM74WufsDgsa4KUIJDFwLAz98WJi9oXKHIvJ/H
9+SztmhAMmyj/Kkoi9t6AJmJEVH84+Gmi0A60Zdgw1DErljWOxY6ZKRKTryTTi1Q
4I7G3PyX4glpDSkpmpHDqqw9a0B3xWsdCixsKMqNcG5vE/xDrHB6XadNtCNVsNBO
y8HipB7K2EJecBbYbfZz1uc5zA04mgMKhvFPWYPwj+oxfH6Om45IxNE/m/ZKlhcB
q3BY8CT6jwEBg64rFXu6W3mKS8MoinDbYShZheV1zusKYEYfzSI6sOykZHbPVwKQ
hIWvbvAqdkjNaUetOz81hmxh2XMmmSsVzCpUYDrNsDpMoC1eNL8Bo5RmG1zYDnyA
B4iZuv80lFAow3Ql8lVYmwJQzAkDnP/YvwsYBqtTAFufj6Uibb9hIn1n+EKuZa5t
jRNh+D6S5m2BqUbQsNfbirBL0hjpPljj8x076uCFPDFsCe3mJB7r5kQAJVK95ZEn
WKckU/3EQ3PtRxodsGn6pRPVXGXt/cs+OU6gpkXViyu3JAOzn1r8cOzNUsuLN764
c0KA0yWIQRzEZEy8IYCFcBWUKaKCyEnLVfgm1o8f45jtXer7SLobx5nqoaebupox
LIbnihsJnBtB2otFvVPFbmEl3fEoGWWdhv84tBi8uOXaoE3GstYaJW9k/vVT2GQG
l9FjdgAo61s/JjnghwyTfSOJtoWBv/UJIXk9e4FizSVPKEn1L/JghdGDf68D7g5B
cGCmm2HIhobOF3/WZeO3SEejsP26NgxuAYGrxHpd5tHcevor2h0iFC8AU+FULcad
yGfUZeiw6MnhejPKc4B6kvl4cLRxktXVodE4hWjCgfTcrJoBDu7wyasBVVTFevzw
GzfezT+cNGa0eEubL5hQ0+um6/FWZZzzcB4nHwc734EQaeYkqlKLwrc3Kr/1mELX
zqHgKiXy3sQA188xXoJbLmlcMX6617q9GigPFXDTtKVCJRp9uIqGaovs24oD4F+K
12KvOwFzr/5u1jwhTK061ka7wmc+ViUmO4G2akK9GOW05aXeu/2tSPS7fiX7w7qe
fSrfS3YDsJtfAP8uZ6oNmOPH9NS0LyyEA65hDLzC3VDdRn+6XgxkJZq+PQZ/zubk
TokVpuBdqyUpBtjpZGD+XWJWdRbGGBKiX7+WRLIq5kwzNTDQpTKOZ6eQTW/X5XMO
MV2P088obtj5oka+map5kQpzRdaJDY2v3WzP1jEV9NB477S83Jv9rEOMyoIDvFQB
OfyARyRrUHjWJ2GOk6rpwnedl+DFnpVwLAedq6UzVwzO+Q37wA/Jjoud3usMgTiP
y4rDi33moW5rEb6U8T819t+2ZEVePDfqODJQtuFhtJPHlzFcuvOCuNmdFgxGK7Gb
i6a5fBQJoIDXOa7y/i0QXYcmSMIWBhWO3LZVPTdmhn+Feb+LzIdegjHTSUwvExtd
Vf9rZlGo3SbaB57RE1c/eX3cfH6+FUiqPu/UQzRc0aU9k1MQiTbMWw9DfZ7dfKh9
dj/ZDd9y0OH1JuDNnxbY7VY6NWqfsmVCzehj2zq4H+xGYJGJax7YPf2D1RXrv4Rf
xGF20KEhNFHKyI1iL066EGUrJuad8Hlok/yAiLsKCQMnuP33UW/5VHmsYUfzrVS9
M+Qyw8A+2w9MCkW9GZjny+rG/raYznF4SbQc3eBSrf9wzW9ADWbwZWYb1kUCrjs8
Gidh7cu94Lk9Sa9E9XjCYt/Ahx7IuBRZnlsAeePcQAgpk+b1rJOUUfoU9yons19Q
FY0HkAv1cudk0eV019Y3ZDhH1MKdbcJa0sSIgYehSk1kTrtJljQi3PCZEKuyWtw7
zLa4Og28dQFhOLXdYfCUZdYtroSPnYAe+umxT7bONnKcVzIrSSIMfPqGN/dr7zAO
ZfuaBaG0sCG0+L6mplsP81+KD6Ljcj6GQ+wteuclcZO7vjsgagmOiGXAP7YezlD3
uvDHtmf32+e7Jf6bxWo97wLdGzbosH634or6omjGzW9hV/ptQOnspaZmbUt5M4ti
YQNomwvEyUX4J+ByrrnQ389nMAxfLKmb/1buw0wxmdybHAo4ngp4wlmh4BqLso+8
3hGcOEdwiJu45ZxUDVA8utWH1vVw8rOEoy6+lVD5F2yZM3lFeLVjtlbHOnck20Se
eKXlN4NJsbCKlBd+U0Sdkcmlw0tvSLSD2/DrCECE/avoDv8XxMy/EKwk0X+qGe7r
g+hQD4Wcs+KQ9L1gySAdhpXRCYkcRGZE+PVC+YEs5F2NuaICVRr570xwAM4n0YcS
p6rMV0NQwyPnTI8061bJMJdKmbtJEsUUeUcJHUfqDLSZCoS1pvyMLHKwegDWKwyr
9p++gX75Bx/fnWtD/cEt2gJJXFS2Wsjmd3EYKpy7exVrd4ntpAGV4WAL6reEK9F5
aZX/BAviRGb3COQeivphLsUN/bKA3ziQlKVNewnfWla23FZosGm03HEk7y4CZbgI
st53DonFAce2uq1yVXRtt41cj018OYIxpB4wOKP60vzOp01CyFwkVG/GFB4FwNxL
vDPEGs2tdLS91/ViSGxYGR597tsOTizg+cGD6tBF5ExBpA4SdLz3j8muABCwPnyR
THvpBdaAKt0ToVgaPB6WxWw8d8lStEZTmGBwfh8LNrjJdBU5MjOG8oAFjvAIQdGo
8O3OJUQT5woneX0D13NF5089JOJQ0d7Rr4ucKUN9jdmFwgaMMxac1WYA2MGqbDgs
JA7uRQNLoysZNpjQ6rq1gT/ZD1nwCFW4d8NAdCaH8ASxALErwoJXsW/NDoxDrg8d
pwTBecSMrKXDCYzgIwtRer9Mw6glp0o68RM1cVPE5VFONstLI6RgUgVj4lI8XnF9
PgdE742f0cjlQ5rwgGh+P7uua6RWQs4lQJ7wFGg7mFFJXjsIBdqSatg2/awul58j
EstzUUu3bs6sIHrskZp9IpVuBEx7L2MdRdacUaxC4bdPQI9yeCjfFir9txjcfoqS
yV0xI3pumzRbVUmzTeEoIUQqWTx8e+4c2Sft/J4WHcknkC2SFAu8dXnJ5KZGmPeQ
S6ejAvXVLtuRnnM0hSpvKAQ3eClc1o7yWwm3sbdxhTEgkXVJLFXwJ7eiDRxO5l7y
iFIL7yJtBPOFoBHprnVdtrwETto29XOyoEFnLv+lHvYboOgUAEMxyjhf76YiqDfM
4J3O+f/rbHCM196j84Stexbz8c8UTfn1clObQcBlsjNl7r/5TvoxYst7y8cYjhWY
fOjj+N1Hszqm2xCIXyiGOff6Mnv5vNDfGWmQLeYjCtAwYisupGKeyf0KOz3qB6Hq
2eHTiyt7UpqRAzwwNOfyRWrk84cV6bq3HVOnRlHZ2aq5OWUnR1aDP6eROzE3lBZs
QbqNed7wFDyKR99UhhYYRoZWB1R6uk24u5doWik8+8HEYzpw+c5eE0krV3APY+8A
mavXrIugetSkwRYwY3soVHbDjUiFHcECY2QJ1mAT3j0t0NDGpNDXD0q9pfc1t/0f
1dUPqb29QeGzGWf3Zl7mVlit4Onx3ZWZcpkXYKF1H4hyUDwKfSBGjj9989veaogt
9F/DkFfTw2dSzFtmrpj0UB7axSBbvWBb3IpA6d4Mberfl0kyUg3BUVljdIgSpFfV
1PIvPWH9rhx3Cmu6LpwuD/9OHFb3vBk/+PKJwq4OddTI3kJ7kS5e7JPO1MQEgLw+
m/YL4kNFf01NkjtYNOCEMaVNllrqCyXn2l/syN1ZZ7rB9bGJsz7aOIpzqxM2x2CZ
GI6BqG3o0O2RZyCsFnIgPHZRjgCLmCs/v8tRiVq6BizjIO5wZwKsI9iAzXryst50
Y7Hkdsv4n2nce2kBqSMSQdhCB1xLFPy9rywRB3nMsziXenl45sQ0C6yC6Of6xqFH
VVPEmxSlZqgK54WI31s1hSQxA1TlZwTcEdht5juRparSbAbMi1wkgdONQSSuqqId
Dh+u89ck/TwPIDUqc7jb3NiIwd8lEF5F+Wr0rab49/Awl1f20mpAjnnO9LiPOHpl
tJW0e+DTNAYIXtxW8jpQy5N/RdnH+vYxyJvNBe5O/ehkXUUwJ5ExrDZNKPqXaoQ0
BBkdXYPnBoMsOSrjmY24pBWEmcQ8vn9k7ktdSnMQhXqBV1+TeXo9nDJpAQl0xGKP
uQid46oxw9rr6YTAqnxFcNh+rP3WBvw5+tcUpKpZ69bCeXvSHmmwk/BJs2JDyfWm
QkK/bWVrLibzuKssvjSK8hs72irNWVG8KlzBDX4zemXG2joQe4N5Dyu8K/OZVVhw
vMqk87jWoESLnCRKCutgcJLsAlVy83Nj75cosnAWq6A7/kHi85wElOo32NPp5rOr
kCV9PkrRl7/38TaG3HGGyZFRthYor/Eg1Nb8+OBpc0+TbA3MiT2ZFoZLpoKm8T4M
MvIwmTsBfGaYsbfZpWmSGoTWZrvpyZKbLenNIzAHcMGRsVw/vCc79BLD4QWs0vrU
ydkNtMy/2+UHtpg0y+0MqSOWS6PEm8v8uasA+s+8yYaIzAwIEz0X5KQSKcY4r20c
0Wl+sF4qHtVIYk4p99LQSbuhPzl7KG8CsY6YSPrrCmCflXrhcoCwnZtKXhyJuGUk
QAU1HvC1bNRQxC1wVEGCRxHXKNl1QSnxwdSSNDh0Wm5vC7rjzfgYL1hoDfyC557I
a6d2tHB8j4cHrHrK/kMEwNiYKUqnbXw9TDdqytknBTOXr74n7ga/qZjFqtDMq/Ql
s2k1wLsnY2Pqhxfcb4Xai62LR7cHjNHcFETxu2v6SIB0WVzQZCwRN7YuGWrlnHMN
iGWGcwDg6IqV7kqOJBngqOXo3UYv2bFXdgB2s2s49HY3qJjunYpSFXofqaakQrJu
bvQ6aX27/cvYNHdhzLFW4RsDqIdj1Xx1peL/vGNXl7/9VIO5Y6IlzHV1dIxrd69q
eznzZcOjMuKidbU2gwqAunN2zCMH/QJXa/n0mjsIqRa+SvcWgnS/hquGRCpfnG2C
N/uRxnu7hX+lMPbhTijq804eTdR5B28VkZt1z0N2NsgH6r9jgVIMsp7X19gZPdpq
B8RY/DdYOkFR5pzCLz4XMH+y69vDOAAPjHU17y7kpjOW4kX6d4mte4Suw5W+8dG+
Rao6z5f3FOaZ1EoCMyxxF8yx9FYCqCTaQigiP7fcvn1pPtKIUeW6noCeIRV+ujqD
C+A4sgiocSifTLZSUgXjKx8TNdLLReC+9Yy/3vNx7r5e0vLeejIFQdGyq3ztOWl3
4QT2JFaDiKf08nwkiczPVsIBQm6qJYtsXtZ0c7XYjUemnTfYw/JeJOFT2uMeLRHv
lbbvUdFhxl2lLOqBxrYS2oxrwP4Z+fZfwkd8nXw2YdJc+dqYyuPXNj7/0u07BLkX
/g7xxuKuNgTbZAOieppjBBQndMZhiQZ7uyIqtSnBe4mlXHUijFM1E7hriij73yEN
cIf4qVGmZUw7kJg2+uCBks5B8pGvUh/Y9rdOhrGedjaWYKn39m3ZegdtSJ3H/7c8
w/KvoL9/m/ggvCntQw3WGRdpA6faiq3jh3iw2/qANea0o8yHMM4I8oBgysqXKkIe
rW7KjRNjsnDDXBDBsivbObUzq0FDQLd2plz5xEGrb1vFsVOAB+qUZfvyjTTqt3A2
vtFVLqDe3QDcsebY5VxDj8/XD0umTNcA/IDEXBuThZYT1tYk+UwgT0lzktlC3fXr
EkQhcasmt1PCQ46wXlMY6cdQg4EEmIm6jvwlDuXoqPXNpkucH6WGaNMYGiSLSknS
ohcfe1I3SyztGpkdK1RXyolKY8b1K/MJZ7xxWiBNBqHoo75nQuwc9qnniYT7F1y8
D8UO3heHdnX186d0neAJUVsOjtQHd6g3mgdhSjRPJAUsXjjyF0S0dDvxR9CG+B4a
CtS708H96jpxerWcIGVJowqnT7Z75hw9sxHgxTcH0YBsAZkKqMIJ2Xf//AfgHoJ0
mhpg6Ld17lmLOQr86bui336kQURKuD4NMPjcGlHOllBk+6Z/6w0X6FVLTYJGQdZG
51saTqv7aXSkGMHV9X502HnC5yClkJ6+q5W0t17f6CPcrGyxfee1Kyb8koCW9o0I
N+VItUJndnIlPVp/OdI4sNywwqggRACT/6fAY6KgciLQ6khQN0m2+LY2RDKSYhhQ
nuoS6y0h9Tk3uDnHOm3VLuIHV6uQCNQRTvJdb1zACyAfhqDai4tiKOhRAeItaTJA
POBLIZPjeC7z3OMzWlwOMpynbgClbHxA8xQ8hNopBPcAeUu7t9bu/mhIu1/5Ge+W
8NBCb10zdxdO7VAmup3mrr+gb8uz35w20cfGry/eJzweJXU/lgY2shqzXy32+QQT
5JbRjYLUEiEecC8fuyh8yqWS8l6TlOLCu2qfvFEPf/yVRbr8SAh43cNIs0Lf3If5
MZGY+yxh/AW/2zur/qgbPsfz5sEg7/fdJOpBqsGwgoXgDjU/DWwoAF41R6vuSwpf
wUppjjshkoJVu2H3K3FBQIV+d71XTJMnl57SPQ6hv3Um0x5Wl26SeiRU8vAvEbWz
6Ii71woop/fKMMtEd0y+p3unGburrLBFCUO2z0djV1WRs+xldyKzlJQUxBKXoGSw
1K34FNG2FdNtsNWkcPD0R5tLtXEr1jEwENropCMfpFTof7E0Cl27XhtZUDR57DcG
WMWLdu7rt9heAxXVCKFPOyQil9q4ba8xMCUz3YPTfXpCyl0PAs8zp/S+qexkQ8Kk
44DtJedatUCJDpQaC+H0e9xk0I/oNjYOYCrcoP51uugvPNvyXDYwp8OhrbIfgKUu
hAtlYt1d36VcPyfvTD/aw+IEfkot0G8lIVeLn2GHcX5XuXhbUxYCYG92TpsrWPrr
4R/UJ2nLf6G5iwXwkCz30A/puoaE7mdnFt7ttRGTFoumkzOqP2eef9mNHn0R4PW3
3I+DtMv789rBVtfnmNaIbv2X6I3CambezkamJEhvaIKIWGCY5guaLDyklSEPuM2L
YTc73W3Xg7laCyWc6IQ/xjBL1CfNsGw5qBdGXXtW/fAcVhzf7nqknlHnNb0fYlk5
CkSfwITs7wGwRpIzFRtHcXX09g1z4MnZ9nKgV/sLG0ftUpx/7rBinFb67wA/sD1G
SmBx9wOzTclgnShX4if81lSwKXdNDk/XS7V5IdU3Gf/OqNZD2gKFuIltw46CH8xA
g+/w7wlANvprzrxqJZGpMWhlJGK6u4cvk190Jkz2qD37OIpMQeIRcrGdCuLneGGf
WtpSds1LQZM9N399TMQFpsY13e1yDQA/mcb9Wytxe6INLGHvQVZ3QKlmU1/mV9Rz
ApEJ12EA/jnJnKatIeJAhIDTR/XDg7bv9dBpTZ8/FgBisajmrn1iRGrq4ouGledE
r28jntO2RI/ABBLzso43d8kaVU1BCRqUypiWYjQV1P1NskqQywlFb0AgtTvpi6/o
nrGQll/fpOgcgBak5n8Z7/ei0mc6qmhXeVuRBP8wgIrihY4c5fKpf977tiVTvt8n
ethsDatdj6vS1m30gkb+gMifewHq0zoBWAaRBluJ6G9AgNxK/zsrhIzd3UPFO90k
tTftynu5OEU0k7n3jnVZx5gweR4TtP12WeDqDx3Bcm/VgpNvqMOgfxASPIrXBEMf
MtoScLu7dknTqSND8PIupZq5sXTDfeCbGAwz/nVmk+3Q2CC8cq4VLS8mgFkAEhYh
I8pV1zTc6sOEQwj+hFGA4U9i6crIWJZs+7T75XQoUl+nPb/azER5SNfo4rxdITAt
n9XwrVJUza5a08jck2d8YJCUizJ/hSidYWYt57MJXJUZAMxOgkHfcxHAHj5IJn4R
W0RKrc2t9DrvziwYmt1oYD99WImZVDPo1hm3iaDjfUXa0AIjArf1pGgGuSiA5E2n
hI56yFl8XmjHJFyvNcOoho/HWyFE4ZoWPcFzvYLgme0Syb3jg0IhLqlVrc4XEwwS
fJv37kPgu3UVbxHFaOQx+DJq9Ia/gXR7iSmEmU/VxWDdM9S+GHKKIMlyArDxJ2pQ
A1W0j99m+dI2fQpUF96NNrcbj/E3BenGyb9+ifq7jB8dC5gFn5cWGggs4vSeujmU
wkfKbhoe/IzTrgMMKAZAuUgzijPaAOdDddW0t+oI6FirmyEMOTr+L9SQ0ln4c9ls
AOWebo8kpdzuG5DVFwEFfygbc/njAM4I/sSzLKOIh/7FwtGZltMKUoO0Fl7ATlDQ
h2yx5z19TkQd81Ow/W4dTEjnjsR0rXLYNsK5jH+/s45p7E4+GW7wHyKtU1JkH6cd
9Q+0Jw7ES8sNt+dniPvsOvd4tcTCh4SlTv8JjZccI/Z3RmT3NJXR4bnpYH7sK0vC
GYhF3HncAXxLY4RdWRXaKnEt0CFYKdLnyJtaOpWsU42OjU9dam5JeMkt7xcSjIk0
xuTwp7m0R8fZ4dB0l9zs/NeWB24VV3FTs4AxTjffN/m0hSdJLAZqFQySaB2vtXyX
EWOpurQHcAoEDqsaVWIKqpkMul4oPB2dwN3k9+Sq3dnlBVbrxFt6V8YtU/tfnJJ3
gVXKiJnVuavhx5cEFubEKavEq6swtZhv2HdpJY0TidsAvbb/FEU4tEq56ZnhwCAD
OTNjuXYOmEsB9Y59WVL81hlva7ExMOFJ1IZi2id1mw1tNYbjtbM6fNXvkyKBKGsd
BC5klS1AQkKpRN5RbqeHW75sP6mhwaFEdrllRtMnStNGeI8ic/zvpzBPcBQUFHYe
HVjaEXvVJKQWfVS8KRZJQovJnDGXlLQvEewpH3qYu81Ry+S+tyLsGWWxEYt2jfQa
dBNp4YFaYjQTXdY70KJb6C8SS5eQWq5v1Rf9kJRSpZfp2ubAx/tqcT6nFsAJD/9z
WlC+yNoieNtnFHrpKXSCx6G7E20IWpT6vE9qVyoKxw9QftOS7se1WmzTgMCQnyvg
f4KBaqGNoE8IdLC2UiVzweWaBBGudnbaD2I5in7rM7E0YlpwsE/SBbtmcFxfD2MI
LF2E9vgRg5MBcwoKyBICr8ENkEslgE3qjklIJLPWMwrwKHlAWgcoxtzCgv1rwzkC
GHqZaAF5fbu1wHe7Fpzh7TlVHJeSUqed+2sEfNRn2Ggt0DSsT21ObKdVMEK0yr2w
lt1QzIcKr9JzIIH9vBThLw6kMJBXx9rXapW71A/wXbT9hK0dYAFYSGJ8AZ9LfX2F
YWPKfUQ8V1r2O7sFoxFAf2ftda8Bsdk5KZPVMZZSYDPEUANTPf/gPuNUNfHyDAiy
92HiPAC9nAhBTwO+4xvwNhK0CjMvZUchKjQoK4vI4MyEOOpmQ+d0gIo/X9Z6d5Eb
gR/7jxsywRFs5VRBfvNO3qgV3qW6/nw9Qe/5cj6+yNP8bBkYEjbwjOol9mSoEBcC
h/zBeRHcdjomTbykRxDQfNQaSTmN0Js+Udvt9ovnz4w0mVog/nG37W5hxiDvToMO
k1FSaa2WesqjVnrPvMC2S7OeMS6g4UOH6i//+Uza2EIFV+GgfIAm9TGqQ8X6PMXb
SH3fbZkW8X5JZaqWAlLqXJtN5qjPO7xmTz+pU/FlpKWGVIXT2JyncmI4ZXV4df/p
4TkWeVc8nCuzVChR8hikdbh8e+DDdg5xuhy+gyXMf1Yx2TLsftdmNYRTGbrGB874
NAS3BKIKHj7jUmxPvfxNnoNp+WPT6ytZnUHHSFx0wzltBeo0XDy+rkoBZCHDdUdd
DDkISIzs0Vzoc0MrFMPgCEE65EpYxduxcj8Ejhlzeac4CLMMAtV/0Mqg2uWnmL1X
s5yOIF85GpB4nAyHnrh3Zom2j/8TGccA7ynPLTx7GMk6+dJViQrON+rVlLxqaMMr
stIvIMqWGKqlTmqRZtmUE2kWo9ek18/II5cuVkxxqutde9OE4kyNi8a1hdDi+Vwh
p4QeukH0x5uxhk/RpSspIo9ZZhFIU0OzP74u64pQWn/CkKS6KhgrnlOCo3EGbeKd
Q4V+BLI6xQo3PG99EXHi9Ux2hY5XFHi2Lnf2mMizvEokUx8EqjLrmKM5pryxKYaM
wjqRuut1OrWzy+J2aDfxwnYo4HdQ/B2enHcalxJ1mrnIM7l5tXGScyACsjW2nfMc
WKo/ONwK4aoPJN1WSq26chJCx0+xp9/DMRr3mMFUNVFzW07AiVV059DAtS5Egyxd
zJuPUPHGAvPaxQAjbCApUykDhSkp5geUg3LLgH1OgTaZqvtvIT7fhYSc2kIgEmjJ
lFwAxFDUMR1ZQ4/iQ5jbUggH911HdD2TM2xLUFp32PsFP2982wHJAdVX8Gro3JJm
ta8MlqIvMK1FE7QqM0ePvXFofOd0jTGMmra84NAHX1snXiUblDZo5ZmI50NX1wZo
ADB9TZu0jt0pZ8xxsHY/NHsoInBhefbQftibJ1TS2rHp3xpqH2SGJ1vnlbZYGJVY
646Jy0AKegJYZSqJ/Uw9lJMThBH+D//cYJwOIRuBrSP/lnGz/f3AkKWJLQ1eMonO
XO76B4pbnAlNh1tdtTiZoQTzwUVjOkC/bLW7yzLaamyXk0FGOYNULGzazmfNKCKh
2sxMY9/UL6zwqo5pf+23+bZEyMIwjY0Y8x9dCblbTAJQrjJFEwxQRrOvLlabUJHb
vikEkcGeeIk+ymkDkmDYSo+gFRBimSrg3o51eFE6owEmSYbzy21aB2Cvj1i2CFdj
3x3/BmC8Jk4X339qA161ISArWUmwvaWsh4HHEjZtqd7g+Vwc1jOZ4Iyowl3KZie5
GW8MIm42ov6qQN1cD6OFeuVhWPj7fRQ15j6ylsO/d0zWAHwpTjgOjVvRfOXNocn4
Q/7TA2JO7O1M+x1MqtlDjX9wQ+N9kF9ys1cw5jxzC2bXraPWn+mekomn2kVSoraq
IR5Sd+4mbTPAPKf62maUFw2HuYjPM/bz/oQGRKeen9YlW3Dfl8b7JLi+/lsqNvZg
50nbrixK1b6MMe+cDRyyp0TA8F+O10dm/7gX55YJHoeWyMmyGfuHL+8XoYyLjgTp
5HO9B+GJ4aE7W/cfRZaCdRV5ZCz4UFENcgZ3/BISl1b/UNm1YbcuszNmV3D7MHyW
CVkWtuF0yQZs5rxGeaM/zMqKgO21RRSgHXySwZK15dKhpmVPsgypiZx6TjRe8zrw
VUtELfiKnun3uXeFThtsyIlA0KLcN28yupwOxjk4hywzATZuivAo88RUYQsHPb9n
3Kvo84pjdprn6nmnmQSq9R5OKmNiWUo58KbqskxbC/ad2pVWMRbKK3NP1g4yQFem
R6rA2w8l/pEbR/yFUeSS8BiU42pgZcOFCKDexUmbwmdhy4SqLB9K1zXLm+bdYozE
kABJzXqFGlJ6n7bmvfXO35jR63ZqakEaavEBLVt6qU0OYam279eZ5jiP169fp1KG
Tc8yPwY2J4JwM6Y05kz6lEuYZrnDVD+RG54IPRNpgkqW+0D7LJUcHUuoiGormU3o
bP9TbPUIXh+y2lloZkYBtLNF2V2KLzvqCtgCuDQGJb3dma1OGAzx8HHTiVv9Z0kl
xZWEo1j77nDIMberGP1LOXGzncOJVAmf7PBPvkgNz2G9pP2Pm+qWdG5eWiQRLaLd
+DpsUaJhOfELKWAmZICx9zy9rHYnzkyzXymBH6aaYLE8NIJ1i5W+TZErqLoZFsdD
AlCkBfP0jPkN9Lu8pLKKj68LwoWTRJMmgQoNgqhizKn4vlJAjAYElVm+opteenhC
rjymjwge8vEth8kJucooP90bxfJIIosuBuGzQ0wxmQ0Q1+5es2mvJ2na98mPdHl5
mQiz62zQLTsbWedEOfBazeM0sgxRCfDanhRwvE7/Qoy+NRrhNADsxugFdjrIVl6p
NiZoMVqGthDEdKHPxE7alIhj19u7/2js3+mDwktu8zMH7d8OKS8Rj10N9D+sD0o3
BiV1FYiRtlMy4XCwLp2fC86ft2JgqPafFzH4yrnk3wTYnSWD8cM53GBygVwrwU0A
iVFYRg+f0+7sy9sq1nlJDEcZUNc2EgsXC6KzzZLRJCWz+6S5McrgtvgvF+EqMUay
esB9MqypKaByQxTUVMQHO83OzXyCuB6CPRIy/KlaGjVfokqCfWAQTy6OWanAketl
y/czjvIp2UEjF2YLKEdJUnXIXykdLEvIKzz/Yc1lUV5lpoir/27GBpu+WDRAZPl4
VuNpZhYmELgyrYyyc7btv4myECNhl69yJVo0YXNyZ/sN56CpoTtDHPcD5otWQJ3S
3pU3ye1rwEO6+xmHMJQKjqBbrjy1dDMUx/Gz5UCJfB6ePV9PtDjilwwLrG+bp+R+
R2KKtgVK2X3w/x1viOh3HSrk6BYChZ+QAggyDSMN6TGOMIQAUyg7oTD5D59fpsj0
jEKRFdUD1ZmaUmF5w5MNLDrP9+P4kgjzEksN0ox1WorJnChUKTEelMqph+1+aFJ4
YP0mFccOrAn83qFUVFQYV6MpdLpGmt8GId5n5a0Le+2e5qdT2gxsajBX7mqoxf3N
vZQC+4JCDBmBPqJqzcH4TGzNSsPHt/k3DCtvuTxp4rlD+o0MJjXHZ5ppLLXfh2iq
j4P0is5XTB7GJo6KQnB2eq9RUIwjNMbTBugOH2btPZRArFjur4sVOdzp32TETbON
Q6nm4nRgrEfO+8DH3XD3igjyA0loUUDuV2yYMq7ptOjDQZhMPGoE/KOClcoYpjis
a6iKKzFg7miP856jWgv1lFTfkFYajCa0EcnxjQFXwinxHIfJqfPfn/nJVtVW59Mh
1PNRQ5BmSI7NgTiLK+JtOSa5GOEBFvIkcdE8s/M1pEZBi9tIhi0B+OVfiJDYgtIo
PA0Au1Q+YzxOq/tDXBGPC7IQRw86pGFLIBRwLb7lM9I2qAk8UEpjzWcQfcKGgJH/
vkEkaHSWB7BwPk+pDTToeMttl92AOOwOgYFd7/Zoc5cMfvjy75f6r2Vz2DtgwF3L
dFGaNmVjDV6zDPs5S9V5ebBnvxMB5n8XjtLP6d4162WaxtjrUnkEwaLyoyzAtD87
C4nCibOwuJpUBaIE5Yb9nYzeOCOlP6O3P5kKAwyfvNQsf7zbkyYF3/imlaCTFnou
6LOjXie4hmXuCr6VxZGyi8PM4rAk9y2ry0gexD15pGd88ovNW5TCX5Dfx/LKCwp5
Flj92oqZbGkVTY4a07YrIsm1E19jYqDEIMtbc8bzmBDKytB51JURY2EVRqHcRjv4
kpdo+UOd9SEymBO+fKaqjXIdexNw4kvnZHzNSAtwcqD5M02KLMf2F4XbTLjGuR2R
biWIRgYBkfWe2ylV7Bg+1YxMpwfAZD/iGA7n7HBDKVH/d/8Mh5sJP8kV4pLqIWsJ
oLVMGErpB0D9THbUfA+sd+51kLgk5Jv4fsMRJeaLTphR5VGfztHse4RxPJHTLnu3
RFltQ8knM/rK7pTh8ZqlT/1yID2OkDShGKnB0gp1re4NK1Y88sRHPjvOym77LQRK
S1hg6uF41xrmLU3VodIqf7F9o23I1ImT7eYAaP6yDRWWBn8RcHtZN40z2CCN1+nh
tSWjbIEcHRJbJf2lJWaWExiLKTrW7wjfUtOn+g18D1TfhWGbyJq3pIellKySTrK9
XYrhxYg8oupTN4nR9pUf8YM3v60Xs+HGG66xDIZcdZiZvVSZTkxLL8kv+iNEEVMf
dnnjIO9WdU0EKKNHrw1MI4QcQYkEocea96xUiifoZZJwIyXop0irxEOtD4YCLWcX
iQS12B4a6Ej4jSaSaUSVHGm4Vcs+YoNHWMloEsUF70fDgcooQpvCduXS03qGtqAh
14jKmZ6tHO1DjhrYip4gELMnY4zz0nzX/NqG/CFuYUhlNg+cGD2CvBb9/WAnjL+C
95soiPpsqroe4GioCTaAfhEmtGq7twy9pKqbVKY/zbh1qt65skb+sH1kbjc/NXcR
RTe7nJczxb1P9uTnjHQfykPjS1+GN6BaM52LZ/Q1GuLDIDPY8s79lEXDoq5vXdtN
YMgsRggwY0RBDi9yUrdFM3wbcOg391Jld1Mssr7dwnYzyEFiF79GJ3G56/GaU9I8
Vj9ED/eBi4vT895FXMVd4yjmAwgwuhFCvTCOQyb565vDl2xqbeP/mDLJthZrMaaK
rjSP1qJB+1tRzIhVgEOqeBEdDHgcajKSpKE269cPzC2vXOeE2fowrKMY63p6J0Ri
5/BstvjdLIst9iiNuFZh2DBV/8EUn3Je6CM2oFKl77jUJZ60Q9ID9JmGASGosrxI
eR4Ne1wpvY64WSRWa74nWsSEUHMDpGOekZ4ua2w3AWN5PX7GXLtaS6SriIEcvccd
W/etO17pBCxb9WCA8Y2SZesba67AThAFdNlo9cAhLki6ZuzdP8ncEAzi1WIb0Qhp
uk3Fhlkn8nXTZs07weU0qS1MJPhVEQ3qNKUIf7YgUBaoy6X1AUnkTi3LQKGAh17t
zSNdHa/dd9fNOgkc67YBNpfxm0g4QSHoba0sNi4Ae0jOdrwmwUW5GMifuJeYoEmN
VmtyPz44nVeblVuqCSkfdCFOd9hjfbw1pDYgI1MGJkmI0X/hr1teemqLKyqiFiQm
Km8eaoKwEkpSTz9pXKehrcK4UUN2XZ58czvIzlRgVWE2fx5yS23+zo0MJXsLIW/6
M3WdqXy9/j5cz2nxtCHe+AIOG91m1QIBAIUo23nLvmrHi5k1XkIfCZWxIygBzr45
W4447wNR78MdP7L/OSVyfFLSO0ESElf/6eRmRYHpB0SfBGpBmv3A2478+QCsb4lb
Os7LLvO50Gql38rD3LC/7YUXxQEWWnFbTDS4+D8rtvO4+4u+NktVd274RFQHxCMz
X80to109qFiG3PxDq75lMIzxRkiW3nU1bk0sxqYh2Zv+uOCL/5GmlR69rfhqkntq
V4xvT6r0efSJmYxBdnWRIp2rgWpabUlrc4V+7/xDLWap7ymTrUfVjBpk9FnPTQW1
gT3SH8KnbUBxGMkrdGq2frjfWHhlmOu5OH0WLwBO5gCEHP8VbHOoBzk/sx93P5a+
39T968PyMj5WzuGaxPxsIPoKTGoqmI05NCyPzUEAiJ9sC0j+JbTFClJgNJCWzBuQ
6yBXIw8ZY62a4Jx6S/Dar0pi6bc2WrqpirZApjBpFGO+8aYQ2SykIZoRTvitJFnm
OWVdzWClZhHafludlSoIlQeEIkeztYleTwUA2Sru1u7RJVFVSY8O9mY7TUAqpWTn
oqsGPmSPwXbupd/Ed/vjxwcwIBLUiC6rmVAtb9M4riaq/ZkagTGrWmdTJKG32jxq
0pQttP5GEPWqESzPRJyJnm1EVQi+F7HijVuiYFNceIgiFimtm7ZUiYoOtnzNC2Vp
BvevzZy278cDtcu142fVvkDvocS5jkzjTaO2vIBpXySiqVUdCyYDhpezyNX/XKQE
JGi1btdfETiUc7XD2nU+OJniFrvk3jUW1lPya7NtURqRvuGmXgmyVRyHgbPazkG9
neCMbjbMl3+4AarJ9HB42lJnO57vbbiWssigGnzVPG+ktZYcYAkEwrDe7VGtsIBB
gJ7Agp2bkyZtdDTMVxCREvGisdsYJ3Wermp/VC8vn1Eukit7SWHpUllN/XzGmtm7
RS/37mJFQaTljcXMlaREZjT4uHRwrbZcvm+4NIxez/T2/SmVQykQd1JSokv1FwuW
Gh4UrAmclGMPQNmVMyKLgMUaghl+49BsGvnpc2br6VeFf1xflht9mzcxqU9/tQOB
UUe3LxQwNMn70LFijrkHGQMXBvcxfbt19yLbeHD3/tOQozae/YGiOJAJFtRc1h5w
pOjPRlGMbnJM7B0YFEfgzhNFOypacYXD3lFjKBeCbEuY3lpb/lYvn8jHRG1mqwI7
Z3dM4xjpmDOrmthMYlVJuYzo+u+u6yLZe+v3vSSAIg8DQY4eHLfOvYoRB22j+R4K
yHetQ8CqLDZH2EedqNX0KRAtAFEDhSHr/c7bhIHAHkT1qL1Y6m63LqQT90+U0YaA
ipo83vOu+ltZNRDAGtYz6YV7B08L/PyAqLEucdNjpdsYu/3MSBoBeIrWEbLqe2/x
putk1s36MI23eC80q/u3wRpAx2foeghywdFkAInesSjDxYTidzmLhZAFfpPlGDJ4
esIkY0u3wVykV2rD+V6YDiopLHj4ZIryBosgZQ+JsoBXId2R5wVdZ60dajAumBmQ
pnSBgrjShwKNq42Rhi8Ut0NgSGxYRReiASqqgZlQi3xfJkCiF1+QrWYqkthY/DQZ
IkGW5lnoquQ5B5Eg5u33GY04p2vVlk1Tjqt2IZXaqVFsI4KkxobY3neEyZ+Y5ee6
qhHn274TmW9Yz37MyctSVpzrKg9hZOC6di6L7W7SN6PlMyAFQD2uk3eqmsmF1uII
UEaY+TTpyfG8BfxuNlUDzxsBNCEosTOJbtanmb83a7U8G6deLoock1LaeUXxygJh
hPNiuwtFMESo9itTuKJ3pX9qbZjtU5w2SXJScscg4iaasTOmoj6hQxvrmBH4w09i
bQZAKng9mXgGVATjaynN+VzuUdiS2iNuD5TYsoMMz0dCJxjfpgG3MlCyI4VpNdZ9
D5f8z1zF2sRtjTU6RmV4/1y7dhJLtdoYVb/saRqbAUBpWk2yfr7kpopePPo0sfb2
1J5wP+GOBpBVuOrrLZRz1BHMrHvWYyW7Xc/voPGalh8ckScfV3r/Vls2gxHNzF+l
EdsAcUqCWOmt0FsEixX/Q5rhGGa8OUqYlRatUaF3OCFASk5tQWTZXq80ZmFopcnc
/i8aMm7/F5F4kzTceCfi1s6d1kcbC05BBGgKif7Rev21Vz8lTooQhAwc9nB2Kkbr
aMt3Ahwox33hZM7wDonpqsK6MECUd9tUuTRFumWs5pJWeRLL3hs5j3SrBhJgKtfc
fY2WDCnWAN79V/Y1erklF6k3qCRZdt7jWWIjbRgCJU41IPCliToM4W+/RBERGsvF
rsebcrCW8FkEUa80z2LemUrs8Tc/6/F4hKcZ5+zBpAEGBJAhfVHACiUdsSUXOaFx
lfBuo5uz9uVS1rP/ovJBHUKOCdMnaF8ffmrrj4CZata5LTFxuPyxmTYDxcDKF7jq
65FdR+YufGNcr4H52IRepwrOk2/yh+EHPzkA5ldcUzCKdijYvZalBlykEQUZPbnL
lhMHbPplJuFI994yJiF/ucH/sKa0GSb6UDI9sl0QqcU9NO+3qJxc6wanjAo3kH4g
yZiG8gUZvUawdEVpu9DqZDTGBCRK7t5Lxjsd+W8FaQ822DYT+6LxXhUjogX3wkBh
s7dbm/2aIttwuFC45LTQSZjZ94+Ii0a2wbuorrK6wmW0qTCH7C32VftOBqXdA0cl
UR286QhMLekFhkXmOcHQKdZhFbhidT9WUPuVUfSO3kcI5Uypq8+AtvKQJ5U/dSXF
Wro0OL83YK2ocyk88Z6VDIth4AnhSG2bWr9/joaRlKaTXomXm5NlJD7ha3oO7GHf
muWHxuiZ8J8/JJeHdTt/IbtkslIYZS/rHfkiFB6zzofhzZ3L4oji6jAQw73K8zlq
EEjkdlUcyVG3C+Bt/uUEfm1WWgROARtlIKN31+kKKpnvE8yWbAiEI/QGANEwtSBE
u40iB0bcIHjN4+tCSg0hOrFbLBnnVoynngH1x37shiKJpli/11SCkZydPU4mIzhU
BfJ5gouvFpIsXe0T0YkuopMRWkS2ehwhly/W1LSsiZlZOkJ5VBtmMpXnJAWreY8Q
3yYmESEre2S6FwZWVSfjX9TSRuv4Nqpu9DSedzz8zv/4+aLuXdadBQlaKj9rqo1I
FDyGJZeKEi78W6QJ3OKlh+4praGbWP4jA90m9XdJPYFbfBkXAYySDHyTwW0gryfP
HtgAaMl8V8ZV4W/TXzra2tbjhBRPR325jDrJ35OE5xRAYHa/PRnNE0g/zwMhN2vk
nMr/oiBAe2dXYPnpKquL/RRwhAnk4j2Gb1DiUPqRkM94ynTzIKUv+3ZI2FPpfoRt
28CnWWYP+fWmVB039kW3yXoPVdtyGJfDuPdm1ZfWPuM3D9qQ1gOwkDzH1qWeK+6+
Tt29p9kTXvWtZ+r1GWswjBnZkBeIKCR1svrcbUC4NOk2SY7WD2vw97PRdV8TiTPC
0n2X8gIhCt1t+YVnsdMnmRBWEAg57wtFcdPWREGa5NdqnlJ8o1r6GT4AzTHD+664
za78CZRoL7Un/a180vi1+yrgeZ4uFw4w5700sRNwoU7BL1aAtWEByEweTmnOjR5g
7nMaDUP10OzazPFf90wfhTm/d5jesFPjUY18G2E+pIpOD1L+GJwVy8/B5O+VPVs1
H/brkkInvdeI1yG0283osfSi9hAoq5DImUvITz39t+PZcaVX5Wu4gB7Z7tg4gTl0
NotTQ4r/s+OtbL/SGxZlGNiOrRNv8rp3OAnEyzLgs2zBxhcrDv6EwGLRaIF0fqmQ
06B0svB+lsdTaEBFxO73XmZruX8xEdyHHOAo31bGFnrEi7xoTAWUMH9rLKjyzm+Q
GZdE8AhOg2Tafe515atZznJsXXUoLa8FPJlWpO5Lm7t3/cKdfTf7HCvXbnOX2ujE
cICWPt37n0SktEaabicE6ywfHRJL1lUbwfoHTT09F5zRjewsrmnzZCMYHAiaOb2K
BOxniT2O6MK/Gmn1Vb4czMWNNSTsvf6fZ7UzVhk+WWgHC/f/Ta+0etXUtWxQj9Ua
7zc4+3gKtETU8TfuUC0Vgf1Ssd7QOBWe44YX+nzqZXhOntijIbQi+l7ER3SjbXpw
Fd1xyBaVyYDyH+ETOHOaWAtRrKOx3F9TpWzIgIxXoorbGcqSIOq9IQ1AcsB//yEQ
Lka/8H9H+VoTRdt5GKMILtRWsqEy5sWTNBz6/PfsS7TAkQ1bM5QDAvTATPL4kfQl
l5zMAYqODzvHiqi2CyfrTGH/zA5oAGDpQy6w6yDGYu8OK4Rpx50S47XINxcoJCoE
imFLprjTGznqGj8A/Yzh7uyf0bfYKSlj9thl9Nu8C1n/b37SZV76rn2y5X5HcSjd
5fF55ZVOwqUzpVeyR8286GkcAUHNbHc9UW+9mBRNMlsN2FZNqfrJeD+L72YqlzSQ
eWGc1y67RNwmqolYtYWZLVpBZurTYhstLDSR/YY5h46YITKqbKx1oBm2YnoWr0B5
MUrSjcmRLla3S5mtg0nZvLSsg7pdroGjv00WOIDq+9BWTzZtzdkCM6Hj+lUEuYIv
KWYj9Y/qA5hY984PzOw1u6M2X7oofTegviPodee5980bBPDdTXL98zO0vemgm6Ov
MQCPXrO/C7jcl4VbhDPLvV4YdL1Y6rtG0zJYx7bD3pBf93m09WHXOao0ocMf6+xA
XcdBUqE2gqTndrM/y0qg/9jn0V0WuJlmgOOlfYKhwGPw4K9ug6i7XCjL1KCMOOdg
sxqZOt+i3z07zDJah29QwF+wzVTmxe2GzPPqq3eOxoLV7rgT4jc8qKK8ifmD4wTS
ibMTC62UETRUqB2t85NoMD4pEE7GqAjnHj7Nz6+m8V7pCi4U5bBzLmkIB9cCjsv7
MSlx8OqB1UIVWXCWNPt91eI2DARO6bt4rFyU6Nrsej6jCI+zYVDmN1S0GPhzEDV0
IQrjPCp8PZt6VopdqIkIJSJJJKye+Gbqk5sAmP0Vz5qSwLhHw4KCvmo52/Mi5AgI
4AoI/WJKzAusVa+ZzusPfrASZyz0on7SoHrVOfC2SX79Pc4u0K3XQSVw5l0pXhLE
EKSZ/yjbZdTNnvE/sy1MixqB+9fFv+GESb+fN9MwkEmiV9O3bE4m7ERunLmkfI75
ME4xsxxvnUtZEKxOA7liKxytmccot0SPPEYKtAKhcX30EqHUoboO1aCUTryfnBv6
7FinttbOF6OOYQ/XDpFblzJquPlSVtDxiP6exCNgVG+aRglgRKH488yzXi12jkYL
utmitU7qd2oX5YWAfYV38TKXIguQHjJxRO/ET2KQwAL6YtWfCAyRoyfluZxCgQu5
uqJp8zt6ZBi+vTslaqhjRpHLIH9ROxcUt3g0NGl4YVqYUps3U2FCsjWS/krKNyO6
puu/50ODBm5PdVgNgVQ+podCfnSBYRREOu6i0CKppD5At68AJadrIWb78PoMUjBp
g5a+zI25a3FbsI228wBFomHBKt0Zno5Zo6Y0ewSWnDdWF6EV/pu7IxWW57s1nXmN
zcCdy+vSWWZleAU5lvZxjxtJxhUrTjBiKYa2aGfSQ+i8hrg3hxozN7BYG7tOltsj
inuztlI6bKEN3nXFOWTyJklKdCqiyyE7kntmGDGLdPbwvf6jGCpcSuS3teUvTJSh
xGJMhrcyQKhhDu5xx4GE8nxlWWaE20nwiBAO2G+690LOTH0XKmov72EINyRxN+9y
3sVhWhT6rFIVRkjLnYCgrctReZB0jiHiuHcCwvsb2bNfBZWB7zEI62Vw++Uo5d7n
0wHbC080/hR5Mq1uat7ICZlM5GGC4mqwJ40r0+w1HzChyGJPZD04v9yBAHyxJ851
Ks5rzq7KMaZgp55MhdTICrGMlDdqV2WPzfGjr8DgE5/8W56ig4Q4udCC/ox4Ovtu
tcZrMPK2aFvQ/fVq0JF1tMYHu5viBgqlvWMNMBS6bB6z6xTLPcwMwNHKa7GDDDss
xjImtRS95LjHBOa2jCj89CPXWZtCJgFJdo5oZgDeYjjltNoTtAPICxhTF+FyUclJ
tOCp6vag/0xhCdLWtFDzVLHrditR9DgZp8R/SOJsAOAHx1aBs5fyX0OUu61HzyXm
AEW6c8HAZFDVnAL/L/FI9OtKgHMwyXuGKpNT81jnaNhpTg+BAa9SVZhT9Ywvq6sO
h7jDnIUUHC2JJze5iPTZvVCOUAGhb425INaGi0wb0jl5poDs3p8QI/oN1dml4rhd
iIKeSqeetnAhs+xAt1n+tdO21zocxPEoAVJ72r7ynrDxOVbxATSQ+ca8wNrvYDnH
GzF6sqoaMCnfWmnExCdL+mplwZI4/ZNjny+fWKKB68xByO9FjbKC4cBmDU9EID8E
4W6HroCTadL18b8n37jXPBPNw9WJx326HfzbKzkuijEPnLqc4cMGjK/HIACGXxoi
A7Ba33NyQMBylpAbsJoBB40clB4znkRaa3VDEKflmddlLddqxW41AD0+gFXgF40J
bSvT4b3xWf+OiRy44VVJS57mxrPM8wJ9rX+HegxEuqk1fHTAcOBoSm9vjbCTsVT1
j1YyYdNH5LP/2YJDTudMibQwZwJkupHS4MFOsOIqteiQ1zj0IbWYojNnf5IJfleo
max8J0bH+USM+FGP8v8RbsbjJ4LillVpHZst3r3Al4jqVTfFfMq5ZINFGFItmALO
LKSM38nP7Hx3gMhhpnCHrrY0j7wiHez/IKmR4z3ipwOXMGpxq7L9+PcBlxgTusz+
M1UOQppdsWrTLMNmH3mMFDo7EhbEDVO3+56YRPG2A6FIc32pHc+uccj/JA0oXeA1
3sCrDqcOf8mvvLK7jnyiNibeLY+Wkb4Ng9v9Ve5jcikdoIkHiyZuFg4p15yQL14g
3rSbif9mjTG8P8PZHBy3N3TFV9EPG8SMFXhOt+96teEQMVcZ+nYeOHmhlazb+FcL
8TyDnd0iXDUWProaZgbCagT4VAtsUOORB80HoDaIwZPXBYKEyWeKxa5WLZB3Gcwe
fzRoyBi2AJal5bE0Vj8xajNfaK74ZkbA51XkDy9VNmThVhzXWLMUg6eDYt++UTXZ
uDwMolfsTOaBF+Nw8H4oBLCky0eaFO00R4Xfr+e75G2om8Y0RzTKEKvBMFWl/VzS
rsWX4XemKABtk75Dmbx38YF5m4+DL9vzLBlNZzCfTF36wVn2gshJ04MMXAEUAEOW
GS+jpRSfkgYm8s+9+qQPpnomWSS10juC4Nw4Zx/VQK3WO6G1cQIAdbTB2fEa1mD5
v2NfOHVfCyO8Rr6DmafG9zzW6KJNab20kHipQKmBdODwV9GjxTE7rpQxlpyU0jZO
2aOl1EoD/kbN7T42UqqbnOT3pzGgbJvDoa/4xCb+UVdHUKWGlbQ6qPMHQVjXXQlO
szRzYHqp8hCw4SoWA+wqlUJ6/J3aw/0YZL9Md5lU8iW8scB2rm8DbVCwt0yB7IVS
VVKnxej6XbNqK33fbpIunew+6yZAZkSXuv5SrHzgpT4GGjSpGugyVDESJan96XFb
ZD/4OAfFbHV4O+zIqx5Z4kRVuWffOyIichHx07IwWWTtlhNs09YTDDsLXuqB2kmn
5QFN20NfPJJAFX6fRdb6mOiWQ+ir76Z/o0bagt/Vn5A2i0hXd/xDm6KQYwXav5hL
CYOA3s+URSiTTpitRfj5vdusnyHne7k68E2o6JLFWmczz+nRHTdIl1aqyszVPh+J
5ymPJpFxfon7dHiXxLhcsEpM4ZNyL6O6rgVIx0pVLDsLAeAHlxHGdoMxo+O6jeq0
L+/Xs5CLOlBJ1wlEsmQByAgsZvUVVRrRcq4+7cbNBJ3kc9rdK62hxFeN/BnSa52c
d5/UgZDGv+rtfIMhSrznDKKdwtcgkrw1enoLeJSbr9eWvadCFQ9dsnO7Yj3tGfqm
LAZr3fcOoTvuKiwSsgYmVJivkkcCC/ZwAR4B62OBcOiVRlJBXPxIlQsUJjRuYVDr
F6MOnOv36V69/CCrIaP0f26j4chowcFfHtH90gL0o74HK+swHNILVoUleJEXqPbX
Q8Xwzc3WueHQs2QVs6Wm7WqFC6YyMaqU463muqNI2Fb+HoREp0qrIMznK7JemJL5
SJZCIquDBtd/xhJ7w7eQuf/MeLWXpfA9UnziLmCoH439rs62lUJXBYtSSOJpWhID
0NJ7CWYhdtCOq/SbgU0D8oNHO9WZUa7yZALoFc+bQFRt4HnthCEk3Ol08UAW1pCl
1eMAKvBGwq2MNk8oZQP6GATCcBpQMbK4GqbFiQDqsrR6vwN/uJ7rw6ea3ivRU+6g
OsLHOgzQ4z3YmkfmOFNFvE8J2UXsBy2SZnwOqyjP9tspiyi/mzP7JmRtCiSBhNBN
S5o453NrSTgTrbvo+7d2fpDqBUepjZGOwkXTLMbVrdpe1+qJlymdp6se4GEbj9Gd
n5yh4AjfOcuZ4P2hDWLC9RcdkhiaW9DITnbnuUkyYLYO5vsCzabdqyGLkjfDEt1K
e5xOqRSCwxCIr7TnAm0l4DicGe4So9Lol9dCm2vUJDv3xVlIuIF53dTPFU3dU6rC
i5cNq/e2Y9Bwy9bfltJDt1fWnFJkqLrqZMPwO9bJ0ldUZLs3sRbgVnR3KMXIeL+j
RToewsjqhQf9nUYgfG8MDhalyweYfwerO70hi472NCRY6PfTIVfSGXqDFBcsxKU2
B2QOHmU2abI/nQayYueEXG+BO3GokzsDY/zJEOzzpFNNkOmD9JOoU7PwAAaNyMnX
Ad11nhSXDrkCL/UbSMrgzEvZc6LRi4bY+1lPAm3sG0Nc1G/jKeQfPuk9BYZtUrS4
/9hUTYVnL5Q9z0lgnaT/R3S3Oavx5LcaXo/y3FOxHxa1wJkGcT//+ltVlP/fum4x
Hx5sBsT2aSSO5Gu0VgMJ3s2HpcbGfRpFPwuAzjUhecmgkGZJ8HGGNAZN22XgUVve
pHdo6u16AhRLaKip1pS28TiV+uKY20H8toUbJM58JKPerQrW3l84236TdiwjVOJC
OtVOuznoWuOQdm1i6jBU2VgNblBImiqIO4T3BpbbNNaMKSU7T1KXHofRFD/DQVdR
t5EE18a7N9S19VyFlMHCpf7lSDgOqtR0ou2NOP/13+srxq9y7z1c+PXi8slFoNoy
MKnY0l0kdSXZP7Und11Nd+PEporcTAshSajltCsk37e9DUZ/+vyHsSAaSSitQehh
gS+2sNMGb6QTMAa/8wAvez9lKF6S4wioKKaD2XX58E9eZf/yWKbyKX+08FTx/ZhJ
HHW5EfAsWBnPCBXFgp9KfQ5Wu/F9YOghv3Wo/Ifevutsz4tLg37eiKxTZrHsKGHB
DtilLwS5R5WUQ3NdMX2uvFOIDdnNmxCI4jaw53vGI3iOYM+CqwVIl/85JqnqVTls
vPPSjt0lC14WI8NI9RFiuGpSsj9KaC92jGV5DJS9D2W3Y/blTtqLnfReyGIPBtqq
JOPL6gym3N6bKT2VNwwUB9mWUH68Pb52K09MCdcMN7bcYgygB2LM2/g5H8CUtpO3
/XX684J+blG067/N8tNT4OrPt0PZGudEqo7L/SpE5srkxKYC1dXznRsBkFuwg2Wx
6ClF/bkSTh84gv6f8GSSLIZmcB92VrbFzTx1R87E+rjcLx2+Vc4DEDwMU5zUP+Sz
6wWfAdcWxi74XLp6eUdxVDiGZSBk3xnyfQfLp9FJPwUrV7w6pMeYefLZ4jWbW4Nc
HpIBcTie4FyjvgUzOmE8DfagO7eMQ5k5XW1OB/1dNN8Opi5ZRTY1iWdO6BsPXRI+
BSrPAoAIXAyB4nIO5XFHYqA80nBfhjDhvfVFt6mXrUopElIKpxTZcbsXbeU0PLUy
X28wfA9LQp6Mf6ZXu/kPR6mr0S5VostrDUWdjtaWy4H1xAn0dRjNnlEX6IDvXwFd
NwKvcNLCfT92G/OutmL80fB7097XbAiUiiYbFF1qrFIirQtE6T7Jw+/+SyBzCqUX
GznMHqYrJ8+yYYWWlV0BiqMUc1YvTRlzGWbFT3eibBqcCd4T6EmqJJtGMU6/AoIr
S8WJ6BRKG+SJcbBlvdjLTFM5lKO8L1/78i2QLa11Entm1GE101AD5EeKW7OqilT2
tAYjpiqHnbXcWwxBvUPg3p+Q+cONooJtnRz8j5OF+IE4R7D1fQf6/Lb2VGuot4Vn
R+8Vk0elR+EW733gViqc/QpG7pjsq3KPs8ecc5Xt8iSYBVu6f/wBwEwL7zDDvYd5
DBj1uvsaHTDJkDpMWTGMxnUQmTzhq5d0UzgdzARWrHdM7rAAJgtY5CQRVw1I2ZlL
EjHS7W7FlfwwxSDMh4UupnUMdAVilIDeQQaF7m/Ci5PYgR4Grjw1op4vwlqJ23Q8
oBwO9nZ1QDjSPiZdHu+HZQXXCtsTD7q8H/VHSsUNlkFCqHWg4KtEt+rIidWd6L/p
RbA4iOWkCmLpW9sSE5ywNsWHgtN2f12UmA8OHzaH7jhI3LT4CJGY+NzF0ZTy3Lz2
dunw/sX6Lff/UNXOWmfURWiNKYYZwmNinEji0vu91Ry/x8nkKd/4gD8VGCUJeCpb
DdTDz3ZGLET+FD9mpaB4fJV9FB/J+CmAXFLzdYwy81iNpweqZ2rSxoiUAxcexs5D
tH2DcJxrsu8BFH0No6lKDibFGat6Ii4UMTO5wZysIoF27u6MG/RLFU8XZiQNoy+J
cyZL/ReKr0hHesFvo5tOBpnz2qm6T3LCg2Ejs7WovoGxU0datnzbPxvlq9PSl+SY
4XipaizXzDWq3ldbwiIKR1pY6wPY4ETaxFRcUh91M+RlD7Ct/7D1bT3ijY56j6F8
JfA+U05PqCmSKloMIZ5rgRhVUDi/Sdb5iroOxvjmDZbJ28XJ+FnDBexMfcrJqS/k
KBo5wJ4PSB34XmNOajGLNd6jO2lp7MFlCGSujwDRV89Q+eD0iyL6xjPphMaCSbz1
x8LrSWEQg0uJVA49XXJFGcXWEeSo7yt96FjpVJat2YIiOkzgFrscN36jIrQMC/oG
y3OiXPnKkjiQ7tYFzfNLA1g5L3y9JQN6z1MAo+12R3iuvjqBGPkRETtol3N9H/Lt
SvWlAuHkWu1wWAa5oiFpvsAjLcYQ7lhmxW9ZCcolcjvJlMm3xdftds15/8POy1NW
17IYUIwl3lNRi5xuUxg0LHNrdyZQgF4UGSWKapXkQpUWWUO4M+3B+TCbRfraCfRE
vXSXLcbYgQzATBBOnznmQZ2dm2h4Y3uEICJHhKlDpao/Fzvm4+oosqn4e9AckL1d
lgGk7z/Zsc5NZNWTmIYTO1wnWiAsXKbfFcYMzwP5tsONRJJOJEVSLohiuZydsEc+
ZljkUTrjHRdvMRw0HOUJiibzmXH4v7aWSivD3MNlIAeDVCcUwim0ETN2ZLlaENyO
LUGSKIOFNVnXBw/5J75OubXo7WTuVK0r4EqdY3ft2xYfCe///T1VDjD1N2elrpK+
SaC4+ftz3NHzRUXn6W9zepSelbDreailPuDFrDYGuiH02GFboihmAR5YISarcpai
XK0UpnzrAo09SP5nZqKFs+BJviXgyX10V2e2MrIJ6fCYQcRX8orQrlaO+s8NTVwb
8VDrJWhkLeQQTB+B7xtB/5nJci2wZ5SDNHDkjRGJJitnxDvioWKJxDUIPb1btjVJ
xAxvBOD2xLMM5mgX6MAmxXAUDkaZ5T7VTaFijkQp1CFoyaRuGTMQAyPKA4yuyZGB
+FcHrJbXh66MROxeJP598/5o/n5O0Q/eK6azNpuSZ4I4G9yKS8ZHJS/Byuu2vCDT
uTZ6vDKbO4SMXlRycqKgt2TNRmj99Y1RRHM10cpVXtEIcF/rpyJSdayrBEjGncy/
z9jMWeFxsfeScmx0rrkjxZj7hc1o/j/sckvFYjN4TbDvUB65hY++54YIgVZfVKzY
dM3haHdlaulSn7lhgaFvCNQeCaWawhWvoEciu+FOdFjic5Kd/TH9Kr9OWZSVvBtg
pjEiwKkaEHZ70iwe2gVvOnKSEtRHT13CPXHzvFFH2CiX1c7+1SHbmo8p/o8EAN3S
y7n3UklCrX3sN+JJPNyVtxBKHtsA3FxhUoC62uFraEkJuUAJrf1SiLkSIYjjpD6O
8O3JTQf5z2xmOY1Z0cmtlPTPF1MxyTdu7C1C5JmEsFpXIXfX3aAtjKOIEYzCf8Gd
ga4Gp+lNM2J/LsF26tE01vpHfFZ93hW6yYbfTNimh8j87aJSmql+SLjJ53O0Ss4e
WwD1SnNQLOi2pLCKA9tk5iO4eEFfFCKS4ekYqwTscWGNV/GGH/aWHq8A4xJrin2D
ah5kv7GweLVClczBpoTz/7ZRG6VUiSJqb0oB9DH/zePmyuAcr2s4Ur9ETbtl8Cwm
8PTvK7sOsptx6yE2KtC/0yhukt2vktWbIbsi1DUiZL4M0j+1njF8SiY7ggKgQ5hN
B1ww3FOf33h7eTrLd0+RhnCBS+M6Avw+aexYUMJpsr1/Y5EQlIEjRPhzEfx3QO35
iRzb8GPP9zCO9Qd9BOF6yxKeT90Zkj2rn6IqZF9dPaPshMTJplKirUT8FNOsL3fU
E+fhg900RM2tCUSCa48E8Ps1alDMPuirywPK9NQAlGg9qitsgu1eqzW5g9k1d6Dz
021xTxANevIEpuzJQq8S0oYvC5tqORT3vcAx7ImkkVgXFjQwPMM0KRAHf8xMzj8m
dQG/zA7YFmDDitw9gDNp7XyJ5jQpwJszfjsccZWUKg7ogtK2FxEkmcyCWWDLY2Fu
rh2R272JOGVlyVYV/0ItpVxND2n0KtRMgx9kpDFGYFUbcDFeY8GpHTuSzFQ6gzS8
6i3ijB4WrOHXwjN2IL93LfIxd0are/Ai+W/YUW6VRbozlf9Z4kB15Tg7/KGLXF17
fK3ddHD6FaG0/POZfGICE7V+HMlDB2JbQlr8bT3hQr4a87aCiuyYAf47GCOH//yb
klDzkoyvx8+R/O4zu5wP0dzNAP5ctnHJWIOuNzKLpNG7BH/NvL/TnuT/viqFkPWy
OlfE6n9UOsLJRWOIWoLS0NlhgLwxuqJWSAdFCX3g9+wYvJ8z9GRabGcmvXhXar00
cggpXHCecWlyxlSa9clzQGsQ5SmQIxaOgPL/5Ys+TdMNxf0RZT9EmEhUcdWvx6X7
KA0aICVv1wkCg2BmCrLUUrIOaf9LmVCwVeYvFOmOyzmcQIrgNF+XxZabQ8AUDxtN
JOJ+0Svs+ZN0b5MdLqz5SVOG262mmbkfBKDxf60zIleblzKcvikr+7Q/nnrS9UVB
r10K+DOAmf700AYEmuV25eqnYDBBNrIPHHOc/xRP73BHWKDsnJXn5TQSVQijUKck
315FzFxfLopr3TRlcPurEFzWjNBKohTm0q6FcNG/g6qu2JAqIH900sE+XnjITZMg
IA3sqPyUen14PSlaRdh1jdGYePp+UpOxmaC0jDCijjj+15kJocZbOCyaHbOYFgth
USml3GOFStusDF/wuuVqgl0I3GklQn2R31bPsvq9avzpwqInC71x+de17gvAegEm
NXLcQGNHs/Nf9VOEabyB3olc4+yqQTVMgzhk5QW1mipRZFrv7qkI7i3LqnkkFp0X
GHThA+ZCZws1VV70kcSblaS/r1LMgU+8qf8tZt3/H0JLxdkCyoVRAGAgm3GEYSab
5Ty6+8l/9EdMaidhA35lt/CoQ8fZsvpPphEo9z2qW2AjK7y1t4OgKFfFMfO3/Tz+
EkGqcMLcMOB6HGVJHwG870IDJH1s2zNxVe6Zu8sAyQU8AIQPETFte8m3VA3b3ICf
7zM8iF2y0/HVj7LLPsL6P8XWDVhjypQNDDn7uNzzORCQT25T7nBAAijEuT4eD//T
4smwhVbYbfu4kP18m4zpj1zUjmrCLGAcfXOYbgJR4Il/YAbowZI0jJUGp0HWwxDd
TF8kQlD8mPqCoMZ3UbY1V2hjyfPlUHRVWq9Ik3Sn5jQaYMVF5Z4V70HjNp6J1xVI
EiUBUCE/JjVJL0Gbr/OG/XA8YM9TFfN6Y09YPSqS4Jrd6NhKFOyM9oIlTzaDwM8H
YCTsDNsB/V8rCXBJsTB9OPumgRMUAMySyXd7arklIBnkbbsztjj81PoqWIStg4Gm
ADMIkjjz0GdTOiCKN1KxjJnRiQ5baB4NumbNdu6Wa/zYFtwA+mZ8T1c0zcaA5mNB
xfEF8jL+YBdDPW6W/k5ENKRmqnNdfzcTHacRjV0d0nNv2xiGezaNzz5e3DViSBOv
mPr2DHD2E0fsPrk6aj3NHaDE3EoU2KJ5hayz/vLJp114+/QTGjcmxc1Fv37ML4kJ
+eBgpQeNJFxmp7na1pcST1N+F0TBzzhGcG3LabHVIhdDjzsTrTHIPjFreqioD5ns
pyZsSUpbzokDOuUEmmzEWxxkshpUGAz+kcRAHEGAMzpe6SiO3MiP+firNDV0SxO+
SEcoWD6az9aUkeSUMnaPNr4ZW42fZx7XUBNrEpO4Oa55v4AhNDwLQfy4z3AKtK5V
axDvYE9HBvHjLb6XTyOvEadQz4mUQIZPDu+4YS1/TO2keiTtAKovwUH4AW2Yprp2
nHAFS/bt9IogMI5Zgd3hvOsVNfJMKLFx+UQ0kKjdrRjd+t1j1WJiDekapy0nM2BH
7v8okPTOn7WbkIa0roxbXlmZSyT+2ierYGMjjoAxE7QBeWOkSoB/2VpEHtPhNve6
EvW7xgVkyzbvx4ftc8mfFGqF/5slTlxjakUqYwuZXX1KNvCTo3Kfm4mctCs3Dbuk
lNoQ1LBXW0yzCqUiNlFiDphrmwYZzQC08zhBgy4ZPK6yYrgGWpgmo1QDTZZIfQ3N
mfNltlmNo9FVib6kGCLp7CkrHJk0A/9WJL56WHGFIO/iTDunz9EncvNHwzWqhcmC
5YKKVrNKfDj6h7mgBJVPbPpWa5ygfysudG1bcKS75K6Wo+kk1NSXIeSkh7Qw3ZqF
h96ZalVVRnmpHBdbuvwZG6+sgfZfFkQZ62VlnhUF9mcvLwnI54mtYltx6+ghhhdM
iD/KdGNg8Z1XDR9q/GVAWl11QOvVzTumi6HKizrKJ/otZzrZ3A4PRbuJQpQrrNK9
Yx6qVDOMAHVn3cmDxttvwRVPN5Lug8YF+v8OpXQHXkqMpEVbogkiv5PTgH/uDQqC
ctkpIAxL3SPUgWQejgEDNVmFLFa2CppJk6Ac+ixP213p/EXkZ0HfCnbb1uAXoCor
dRfLjQCyeMTwTCFFe9OpHLK+yQQAsd/Eer5ULprfHqwJoQ5TXMrF2gAV6zN68yHt
Eq6i/kqrZO34ggTgtApxhqeJVNl/UNgcvkW0vgJEHUQiHQYwUEiCKd2ukqUG14cx
jvciR8krY+VagHEWaA6CWAAwb6uHNd5FvL0rfreK58v/IeIDDZsKwy6/Ex5UoJhm
1srIUG/77xXsgZk/lCYjGMyDjPEmQQqifPRrV4SE3jjzhs1ysGfn3Tx4ottc9GkI
KUMCwWPEFemSSkfLmGoDTKlyNN1CmzHuZXwuXD2WKrwY8gqGNf+VChJVmyQWKLjy
Ci5cGz0FYAut9G6zxobdCwiHG/+mOu3wmRdEXx1/ZUq0n/WbzGJ0A+KMLjjwvMd6
tbVeNZAuonwE7s3jRIyMVut17UP/iG3hWBAmzE0S/VN0ncmtEJpDaCh/gBiPJDdW
Ln+47tp3Occ/dAHJi2FVA4XVR0OV6jJ0oLf1toCywS/0Z/qgWxejA6Dg+BFw3Oza
uT85dUx6vsq9gvTeyXbEmBT7GxC82pPSxr6vZhJvdFCRx3o+ljyFTME/sRxP2cY7
e5BiycRMh5FhaQWmEBp7BfVfzNhL2/meTZvZY32w4dyzJfftna0O9+tymkWoP19b
e+cncNUpgTOQr7RExFeTxe3Ua+1OX5IRfpJs/+9ZeMRNiSZCJ925sSO8iAk8GxYF
xR9rHp6kbmuhUiO00rqYGUvY7lTaTxBwExtkyt4piI3/zoxWz/3s2JR+keWRWG5n
hcm5/rkYo5qg7yIVWfAUL5005/1lTVu8MNOfuLB7vvg1Ac1F5qDkyP9eH0jA2oRy
IZBJ18LV3/sj+3kuFKxxiyKmILErQo902eAE5z5d2vKOxo+vn2HZSr2qAUvvNESR
rLNuhE1rEPg6X2k/QPDJxL7UFTO41Thz7XP+i1f3ax6qzJk4ZzSyGOMuJ4X4hHqh
fTXVoBfVlli+Sl4rOwfV2TbfeGnzzEl6w85m3XBavNcjK31DyaX67DAbi3rY87s1
LrQFz6GTMC25QL1lncrcfFx3UPnpiGuDPpHEWFu4Coj8PCdyPsb7trkeHF8m6HMD
9UsNs7um4zhrW0kPwxivq593HKh9e2H5KPUvZMfMxmySXy/l2d/nA9e8dbfx83hX
Ivp0pqLr7zRDj4VS9OoAyF9qAH2M0QWfNlbu36uQ8+IwBQwn1fj+kDZ+SvMWn1Qu
6SjJm1p+BL9eiwp8XMNWorTmK9MQbVtygGnKKO5EYqMhF0IgxsDsXXgg6dPfYWH+
KheUXoqbnqX8qZaTc2oRNxsIdQUYNEvaTA4NDbyA0fwQXg7lvWlk8GfHHGwJz7Vv
kBd53NZyi6KxBX83JrQQR6STn3E82nZ/J0XlLIzQZcygaV9P6EcOxucCnWjIdtqE
hFhoT+1aphtHBAAmHj9EEcj896fEI3w9ex6VcxI8EPNQMeKcRhoQ3IHJDCNok66p
hIrN+X7psO6/E9e1N08FKR/rxEIvcvhskKQvRIWyJJ9ffkirDfzyLPI9J5Hd7Oqv
dzgfZf3zgjcrw/3J/ZQ+fPt4/4GaH5XvvhNbo83i+FO68C5xRf3RBechITN8XcHO
iVdP1j9GtgFBte5+5bsP/C+Yo/pxzCJwwwlIwUy1bPyezh9PTP+989/lUDj7TnVP
wdnOudDcJqp7DcN6AnEvg9U9Eu4fiF+eFJRWGQWSSBQ/wRVCD46JRmo0+JFW+446
fnSt7kIcPo3DnD+ytZxG8VAJRc+sgHs3nMQlZSNzMf0fbT+p0EWx6wxJhyL12pBA
gEkmEaUHfC/lib0xbhiBq2FTijfhhMO53lp3vnZRC/cWQm0XCnh+ERSxBQeQV4aP
/bPtU/2fCV1Yf3V3RRpGcp+KpVB9vceA1iE7wwC0s1cTkiHPms+64c+fadF4un7f
xkiZjdF2kdJFOCBMiAPn92XBE22NRp01ub1VY4CXHORYbFLEa4AhZG0HbYmfL5Dl
xra4kANymNbVnOPrPCx+63OVz3/CC6aSkH3uH25j0LqdqznBei6C8hnhIMY4UM55
ME8ZZVcVe9rtoP1EvKAf9MIYAgZIGaJhKuQdVvxnC8h/fbSTuDe1T55UuddpUagW
IIysJCE0Fcyq1u57Vxbbb7dzBYJnJMduK7sls2ORJA+Nrrwoe6eNpX9ofGh3t3u9
59bkvBHLqrMLUpc1uxCZXISVe+TAWONEJ9GmDAbitUtNmYYleEQc3OpgR8exwxdN
lES9IgxQX+8RFlyb8tCMp4FuhsgIw/dITw9A8FGHpzDU+1pkgbksp6uBotnjSdVZ
KQVOTm63wOyVL6fPKywPIA+trPbOoAEVxewnE0vDYlB2vSEjjZxnonKu8PB2t/ES
qu8pwsvQV6Ee9otgi+GJj/x8JYy5fJv8ft8892p2txqXCqvcrpkiOfx/j/55Ba19
8lrlZtpIM0cyYwO1gMAnYr8b/u6xYkExph3W0XWarhfg7MDrbjBQnGaUC36pVDQr
hK9Bx1cRVT56jTQ7Jf4UTEPERGACL37vSa68bAOd6UVsGUgi45dHCdnTOZFGSDsE
fZd/M037IF/3ruAmRJvkU4Aodrq0SAHD5MXDMMB9PxO6TAMsGddjP4TcDdnhqwAJ
SpmU4XT9z2ubh3QZmFRX1oZ0Txeb9euMiPDtkdp4055sNFp124vX1HnhA8N4GeEG
hVVMnjurRbIjLF7R6VMGidqsI7SbiM5AqmG1Xc/V60hZOheaLV3vu+1fMndJv0YZ
+GEM42oTLQ8j9Cth+/rsZmmHhcfe5I0YovTzmA/rde8u6Uf/eyAOOThCsBXgIi5F
8Ars/OIzOcRZOjVhldJoSd4RNrJI2obvneUr2k0YPwMTeovSegZ+N/1dWA9aVxIQ
1KRHiW2fD5bG9SnPBVYRZxrUy68BdXRLD2VdmdKJQ2L6U15Re770U6Z7zyWmCatB
cMTiV4hef7jqru6JmGrwQBP54kMFkRnNFD4AqZvDSeU+gKsaVeQTRLHPwkx7MDEH
dhWatPZFlwIwVMWsF2jjvLaw+B6LerpoJnUQrYqWfOr0bLFe1eaw8FRHiVvXY3l3
9FTXJBJqUimKlxeqT6jg7vPE8AEOcL6YIKZN4B2rRSYxmOWJqLxpNTZ16AKfTBzb
fGfnh3htvu5fmBTZHpcsGajCQAZDlSH7n7FYWjK8nbHBngRHy0FEUzC3uYiSOZ4r
xgrEuPWD55reaUZ5T9EL9YQXvbDDDaDdTqXv9sq3wQH99LUGalNJ43W2mgMSsqVs
gxLTER6wiCbpI1SppkHyTK9vz+0twPdGs/08R/ib+BexSPtNDDio2UqpgQaypKQw
UkQ/+N0y8nwdN032c8DezSTJ904R9tLhHYo1T7/bSLAL6w+u2n3bwX6/bvC9boqL
gnzxzij0Uuy1cAcAMkIc7MUIEKLfz0KJQE8p+KfqZfP3TxUyP7VzpCxYsSwE4jWu
xoM4L+ZFNejhI59uBMdYem7hm8qFI2IcIYHXQiK35Pg9lShhgdkJTflTwKepZPkk
8lsLISVQOJsmgnUJ0qHXpKfMXP4tn8dF834QpMTMibvjq1j/lrNOrx9ovynk7wPT
B0lEbxXRsz4CVzT9hR0d16OpVqaeNgRYLMmai5dPXlfkTmyeHUOcVGGHqniw9oOv
bJfjvq1lQ6PmCqggzlCBVE5Svxt3QQm0qOIW1H5RY/GV7eIzUhMkIfpjmVGzzAvH
DT3z0Y4jcm53a8IMFD/HvpXs2xFkuIiXUUDowqOq6oFPyZfcA//hAqIP3p5mljoS
tMIGfMobc09K2uMwfr0dAZzgSE7hKtEQqp9ijCDDYBGmu4nRKJ4ktY4QAtuURk+w
uo2OEGn8ACAQN2nL0WzrFXbysa9BF68ipimxUcLLfVvPB3yKe9b/z3y/0kli41yZ
8lvuYrtxxOXadK8BFLe17aNaavQX+I2nLHuCVjtqGBUE4W2VSWLF0XW0TWfv3EWf
nhE1h0oFlL38tRckd2dc+aaZMIezuQTrWlen6r62XUxjBaV013qrFzBjr/LR0rHF
qqaze5cAIZzEZMk2x7AdOBqfN8rEXJmpHesjcFMh3ZBB2ZcDzX4m1kHgX/kMY8a4
ynd8wuEqWrJP/566bHn8FNzjTsKzX/VLrgMhHhE1RiBwJR1PQS5mwT6pKEA+twxP
qqlVNWvThyE8UaMk+1rNlSyvKlOAxzBPCQhh24A3JkGZj8XbWnwiOJbzSEBp5D91
rR2fIO/p/a3kavLJxDHtjk2bB3rGEMfa3aRmaa3XLm+uhU5FLZ03A/VBLiaXFBi5
nb7URbGTYKTPbE/753TYsua/+BRTa1B0Oltdeni01prKMNvFOEH1CiGZ0oSejpXZ
k1bVKghG7dEW9g9P7tnMVOzSwgrtcP8vTkh9Ar7x/iOJZHu22IP8Gm96Oif231ok
DRXMIvVKEACoY9g7Nje7vbFRbo6apM/lrp+deiKKs0gPxgE1MOSgfxF+b9lJ5w8n
t8J6zXQh42ajiWWsl4bENUcn8dRhKf67TNMeo/9P8j0owDK9J0qOl24/0pbSA1NY
j7JoT4tDAdo+VQKBuVykUB1Aouk3u43z/n21WY8Oh/bTDrPI8q3yyE7VUdf0XRxY
Wr5mT9DZ2+mntXF8eFM7yAmiWdb6kIbSlzMhFk4Xox/agdm8TaY4nX+PVqYsE+pg
kFIvVX11krZiw9C8+5Z0iIZpvyFpIsjFt0VvJaCryzTu8VuY5neNeyprZ7RdpUNm
CI7ngh45u/b8GWKIVxy+BolzM0XUH/E4hoUnscefzCCGQxQnZsT5dkm5etjnnnA4
xFfD6N7UivtyaDeW/Tr9urNrcXxt7TFQ1LMduBULhjQylXy9dIQ/uAwZlxe/9ngp
C/cdyD4eogxmHgy4HqgPP51Ccud3MjlZ/C8YkERKPUx3yB3P04SflZ2Fyp0PtoiT
EawzXx3BxQjDP7+spkk1uPa3ZC0NlvQ3p3IVttg3qcRRao3hWISTACQh4YrICnhj
Js8lDewTm16BEilHa5mnYSjvFvkG771gQsbr1pCGqkwdP6H9IIFjw6QIgfb54yXo
3W6qqG7tlR8KwphWpy5WOzWGSivWbY3LHOUhj+PSP0lAJ3tFykxeQnOnQRQ/U9D8
TzXFhYaE9EFvHxaVNXw38FKbOXmlT9X70b0HBdl55htp7R/MWFf03NhQ8qDV0kLx
t8U0BIRXHH0A113c0oPccnKeInJlbAp4kt+xV4pS6A+ehPR9LEyK1Uypq7wb6Zm0
d1oE9ODEjf9I22d6RSs+4YoU2KFCkX/QcPaaxlojU4RG5FWTuALWhWRUS+fItcM1
4tlVaucMABhA3iWm9uPB2mpRg911Df7feB8YZolYp514wT91nkQM0Laej2C59+3T
ss8pqisFLckP+ANFLvYT6s1YcT+kBL7uXdoXexZQc15kXAGkw26qhhVNeZTIGlg3
ztDiWlEQ8bL+3KIx4ZyTYcG9w1AY5bk1VGA0Y19nquKrFLMdFyogS3ZSaOlQEl9c
eTyvjUf2uF8MOXjA3lEvoOfzesQRsCXVSpWE+1ehGnJZXL2oEc7Xvnl/1RZJIJr1
R4Edj9fI4kn34fvC6SuE7v8iKE63KKVOZSKpLz3FRiXClmEF8d80P1tVmINTKYrA
qX5ffd8uy/mQlVzDgiQomx+Gzg5J060sMVxhj1SJG/24fjpZED7YY2nrenY6HeVN
P0S+7IoqFgsbvB5zXxU/M21ckZVRB7M7ZTpEwA1XX2no7RXeBdJ7/PG7FTqZzfan
IjvLM/q8nStodQ3Ehwpkp8yNcGjfodNROPdQtIqhwKes+JAXzTIpk7l4FxkDwaOK
D/Qu4u7Lxa39XfVwo3il0vbjqRIsYRFNldaghpg/crfnMfz+2R8aTtChGmYGcj2d
hzAdSQvuIdyH03xCkhpB6Vg+8C3CV8ubMw0+gzao6j8VoZE1QM66smhyyo89+Ff4
Vd3+CJEc8GVESre+4if8Am6vcr2O18nYz249B3O7CKto/nhgyruLfbj32ym3i1Ld
pGQ/CIk14GppPpWDCWZQ4hWfwek7CsjP4ci9l1TN3QyqT7R0f8i7otmeWKW+s9k4
TweH6+SuHB39ZOlt1F6v3YNLg+9Jfb9IoG/WOFTgG5FoY3eBOdnKk7fMkfkRjuR8
E1xawIIPxo2xw0InIjMI2ki05gka0ddZufMVPRckoO+MRMDOLO1sraKX+4T55Fnv
yUbFBil8rjb450nvCGzWO0CnFkLwBTeTjQVP7alZtmOacyXZMaKjUSf0+/uwVCF4
qKo99kne3NwnKs/Y+y2FMLUdBzR4r9FLk2q26p5gLUM2jGbzr4JWCIXM0pWcaGKZ
COctSIgwcy1cHaZqlPHDSCZeob8cYm0pYRAvkaPKFVsrJTeSowzrkhbrPoSwrRyV
OFwRrh3Qc8dAfbVgVchU2Jo9xt089ySoSyFSCppNfIOcwlhmhmYtCtTF6WcgG6rx
Gy/Ee1EUlFJuJgu7ubI1v74Rs/Cl0fhGaG9IhLYfnwyGr67YGsYj8aX2cNEWTYOP
LZSwDm26PmQQkvaelRo7a7C3Fwxq5T20wRW4FSXRMHlKZ2uzxQ48I+Gbg6LDGLiN
Ecy+kkTQH8qsovLBPHlbnTAtymFQQVrtmCydsvKffjeQ48NH2D+lkaZb9AEhuGti
WtSo+pTOTsM/uw4WHqK5xVpbneDVkghGGgwaLztOo/h191TT49EWYamc2iJN+bBa
WAXcBrEuQB/h3FQ/WvsmIvXZQEgULBH/JW4BxPOrNkPZPGHT6+soY6VeEhY3eJEb
hxvciVyeMCqnou88ixGp1J7BsXNbZq/3JmMhEvheECJMpp14H5y1t8YCrfKjAH11
L8+4DWVHS3UvBnm86NhGyA3YH+mRorX4YlOqf8M54rXZgLES4b61rvZLqPq6ypZQ
CZtDvTrgJmSBv4WFn5+Aouj4mxh5UEGKNuVzuHbSCxbdUr/J3taeSOT9UPrRvQou
BazrkOVK1+4p6qJmKhIzENEnpzQhXGyvYCzFHR5aGFl0++HKmv9pt6N+E2xfgQAJ
6BMLOvicIIR3Mw64LIL6WWgYLyhrZl+JVuUkm/nKXtE+AUNsySa4tz86eJiYkODE
l7RGXJZmIe/HATbfbct5Yy8O6nxXlwNrbeQAfN8LlbY+tKOON0AJQUJTTvnKFhfj
gRAMapvUiRVyvM3R7U9V04jx6S2/8R1WZduWI8EpSJThzl2DtDAJa0VHCDicsYYP
Uiz0+I9szCaacR+H1B9zdPLWAMQyib96VOsWrfMm7D8z/SJLFwG1sYCxS9Ns4of2
1Z667VMPfHvzIA60oAG2XSnQxMJ821kXQIfv1JPFsJuN1M1pUb//CXbe2tntSJzG
i/z3/WQSPHGJA/iDFvItwZCvCVUJoxyq1Xlysy6NWv56OT+CzhaAKahtaWVnW6zr
PVAwKivX4yP8Enzhy9sD4ckSaA7kQjQd2a1W5EtJWwfJlrYWNQKMoDIkLHosvcu6
1KFrnLY6OgqKVRQ7XbhiYIZjoSaJ2+D4GGqrTHLvkGo9i1d9rmrAeQn6M9Jg7dOW
/5rb3JCFsz0sNA/kvTmzsPlOxCq6A4Zrltb55TWLH2kOF5tdgUJStIj7z+fKUcob
kdNqtSGEYARniAcbvhGaOxHhA1RmNCXtB1HPzTVI7W3tOhmkL/ktqHChBlFHlcvL
bVOy/OK09fiY6AgUI7U46wdxjzE985AVasDoqVJof4J+1srBBCDYJUnF8W0HBCK6
0xLQnRWbUHK2cA5LjOankxI3WKy3J75/hsVUyIraeEkCFrTI57hHhLTXw2ZkCxqf
7wv8DUT8EANmBL/2vdSBdFOZUmi27ciCzYmIc7xAdcdRE151IgZsMbVemgaV8e6c
woK40dK1TuPpPwHlcc7LS9S3bxKzHLCEb2DapmSwEuD4Z7lkIAduZPUB8/eguEBl
ZtRwXNExoNsv3IKm0YG5BhsGwr+yuR1Kunxrr822RepJLKwi9VvLwCHOpcEAb2pA
H3nbgsVdFiRiwb6RPkpROa99e4hzgT5xsemC3a1VJjgNabFwFyjaCu9wb+YYLLeO
Z4X5zw4zOVbhngQyi3BgVV4lH6P0E7c40qoHmIrmGRqQpMRvkme5O0O0T91kvRaw
ktukC20B6Fkx39a9rpR464upezG2keLPlQ9BgxyRB+a2xDwao2fezddJQe38Yz6g
9H4ifO52R66iiXVkd1ShocrKHjaxwgOJR2WP0aF4dn+V247LY5wgROPSueC/zUHR
VigkMDsYmeSpjNVgh2y4OK/38QRyb+/wJnGzZzK56UeZY13IkGBxz02VMlk6Rnjr
QDVQUYOcWXhdUL7U0MHYkXRY3RYBs7jUIZL0vYkwELjcOyYZ22/ZKpN3SZ3s7Eka
+e1wPIR+XDnGPHMqiaLgV5frRE5jxZ+l4oXRdQVO0Jr52l2D3Bh/2Rjo6+HCTN8/
l1Ew+UyuQ4IdkDVDxFWQqAp4HIs9a/h14OLeqqAJ1nrp2W5M0wNmzbGFgcP5ogm5
pQDwDHE5IJzEfUGWwybBBb9b3L2yg91ryNs5bRBqMPU1yw4G286QoF2vmp6oodR6
5I0mA/YM/ZrOXzQb6MyfRImRVji/16lCBjVtweR3WXjaNDWd8FIRkb5gV3sK5qBw
3XCELnbeKlTXFwlHqao0u3b/DJexfyNwj2CG5sXeGpIfqfqc3LW4kgIu2/O+xThh
6DZic0fxJxXFuDC/AP54PeYXOG+lu9I5Ja2Z3mR0NY9KZHucXHY8aQ08HZ21lJkF
nUUYmBFVfKGnYW+aMq5ZsMhbRKooEZHRX5B9EDahv2e5W25blt/zPs5Ar8VvS5+b
arm/RiO7LbnF/JhHWwrNlKf3lvnkQDUHahESvkoncZenuiCb/MTNkzSQJ/urXk6U
G3KqyA9FX3pk/kgcxHixxxNkv56iS2T83OfLTmixi29xL9IfA1PE5gbizsN3Vxk9
LBsGI0tliwqf5uKfwZnhUtvbUA3l2BFVwYxhu4rcz5ev70LQF9DIxmJQLalBiB6I
xyu4oUt2xITzgWP43ymcpW5pgIo838wXjnpEuXhiD8Q9jCk59j4vTMH9EjzkbaiQ
u17lEpzBXX6GQU++Woz5chi4smMFh+oBKR4AQ3P8xChovM54eb7O4lZis1/XmaT6
jWRXr9Ywd3TiN9UdKsWdA9cqrdhCbt2xB+lyncNwczL7vCKljub7QRP3XAw4IMoj
PPvfnDmxgqEaO/ffkyFi4OaPm1VPfNRYGCaZEIw6pwpDVmRhz4Z+iMENPavyjnNu
xSD3+EftApkpUeTenUbed+NYkCGMefy5qIFJzPRpOiAefsSpnLOw+SEHTRfJGbIp
p/ZRwf65G4UkujpTpMeEVa07J07vTf+djKG9+SjReoxud16PYMA7DdjyTgFZsbdB
0xMZRHhMcBuKAuXdQZBrOjUDDZkM1TOkM1EZayXDwECSuDek/WFzprirVhVkyteV
Ty23v/CTxLEz+Uet178BI6jEGH6v9vm25Ly9Yg4t46oZHZlB/oRKMNhbDDBQrPBG
cGRE+3kEMY28XmCz9EwbvK0d/Z9ZQe54gDAXzBr/l+4+bfmjr4XB085fpXdAtPUn
1pabfc3dLSHsYtKru3e1ZTU72ke0rKxiN36jZ4Jrhw1BWDpSwKliG0PTgFB0Dy0g
hzQZuSgMGV9Sg+9wj2M+suidYCQnxOR2ok7Gu1EflWNvkDk5mEda50GhQx4JtrQo
5kX78Dycr72c/lk9KGRbEQcXUNUC+25Ev3pt3zEYk/3gJsmehEGMWGe5nw0IxbjN
Xmi5R01a10cjR3HFh9jh50xa4LTd4/ud+mSJ6b9m2ccIijOrLOlnPEe2iYC5Wq+6
r2qOWxPtAVs/8hf1ppdec6ZyC5FA3wdxvpfowGHZlgvnwyZO0lSqfgxvj9I0rRR0
aUAFPcMZpdzQjO4MM7KStIrb7mmoyxPSaGlY4YBpHkysCxTAxUBVIpKw0TbHSjnu
FR29l0K7hFdg+fdXKvHiCCbnMMkvQVzOp79Rh9VbSzh33iNERU4RPTK4q3dLMQl7
xQRYwiN1crVd1N0lxCtzgqXL6qnOsLf6HQuZdZrbP8kIsFwihYonha6mbneDSmHM
soHIwhKNm1A3ZuaZ/vsFGLEex7qhr416DA8wzhnVXagQUWr6UVEni8fcg9ZtOuZO
V0Gtlis/CTx4b1+w4SoIWOwg/Ci4Jaa7A7q8kgdR5r5BDOVEWaws/hdn5MEMo/8g
n8iXFOWxXz7M0Jl6yeUhb1Fn2E7xdL45WXAS4xqcfO0YSeJjaNcFBdjRxz5jy+n5
vhcCZB1FLMAmCjYaYRLpLZpgpWeazJNUUubf8yFn6RgjzcWf35E3PfmOA91qjimh
6QEqbuVSD5IoFWPvWqcMAR2IBKT5EJM5LakeckG9zptCQuK/JIXLQXj8Hoe96QJ8
2V4LTkEB5QHwaAY4P5aFMkxnlY50rnooSDMuzlzQ9fILh8iK5ZUEuUam9HbCRzQd
4Zc8afTW7Rk1NAXVBN8QQfFfOkeFtoh7eEBwP19RGbKGlmrgHUHNtBzCm5upkfgA
RfOC//acQmAXJ7tpbfvDaYAqJzALSz07cAqtjktaxebV49evPTMkrx/9SAufGYZG
f0m428fnJKtZ5ghVj1SgadQKS6ygLJgTUWjApQXnyi69Yfgq5t0Ha79l2Tq+U8pw
CnpJOhfTVhHIa03M/hnuI1fVyKtBcgAvJ86PjDKkQ9bt4rvwAn8fWI/q/gI6CKBF
uL82yIGkQHPadPrFb9U61LZ1o661YpsAeewdqWdeY0O7PGh0y7pWNsFlTvqJC20a
BR2FAyoZsQ0xgo7R89dHEf2csOUf+ptJJwfKgBmpqf5xQrl0WLwbLyBpD6hzkgD/
ff1kRa8e5n/8gLGYOr9I7anaF0ogHOv7zQN3PQV8ncpbeea+gdPlwkqceOlsNs7e
tNoe5lD8N3XCjtD8M2Tomgaopk9uDQ9xhC/SdUNf8I282Je7Vih5WejaMBfxm7+D
MiV5kv3exjT0MbJDaBKIcCALp91r5hp5I6Eh84a7BAEF3ZIO6bOoXf2NaPCCZwxu
i3a8WRxUEZF0t8cQznt1wh32JfUYqIf4fhSJF2+8WLWfWnG9O0GbSXHLCD6hAWwX
AVMCDBVXxe6Ikr9Z8mBD336Xq149FEaiwwWwrMgz1mmcejy02S/bNFP8mVBynrgH
DBJnn1jRdrcolAowiWrWaBMvSFnlWjxrfZrzMNONvmzEEFdjeqYavsWuHtQkw7I3
a4jK/I8l0AziDaRzgQ/lxC5bX1zeLHa/h3yRD6+pf1KTRrJGYVy0R13lF0JFOTXK
xzNp3yUmnUDpLKROaWNtrl++flOytv6FitYtekqoh1plav5y5HEXqH6hyGlZ1xp8
rg6/oolLVNWyCBQpfvB4R/1AP46mNCFjyQyGUoAA+WHLFj/jIwD5SloiIjNFzIc4
zss88/JQmjigAax6eAziMNA1kS9nRTmAG7Znv7cet7CA+d19t3dTRuKjXzTkPjVT
3eNMLosB8u65TSc2RhNPanH7UyHRLvmFG3DZYe9VvstNyB68oXfho60QLaGcXC+2
4+YZcEXTW5l5W07EFLQHestxnL7FjDUnjL5Cprmx7tbik99GHGMWVFIBaWb7DeCp
0r1jbDC6XlOKjfHH916nT3a9pztzkrYpJHBRrguX1uQ0WITHuqGE3ceQ7PH1a5GI
wBFPQoDJoivy5GZ/FynBxHDZuXKyGqDyPxEFBaWqfKMP+dl3vb1nZ/1TPYJ3BY7S
ec8e/bsPUhdTITpBiVoAZpuunCWlPrE8PjvW9Bhc52yXvW2ylpWJ9WCfzz4covyp
xAUx/q/CKyAjuu7Ra02FNWOly67ASZZ7BDNQKzf1fqMRjw+pCY/L+TLe5e2f+Z9+
imVWFaXNfmhCATNfwfEsGQYB4Es3W1R0th1yIiRVbICLFHsjqTizhomNiAao9XVx
ghQM9z9v4PhCYdF06jxUl7Z1G1YkAryh/fSUMQrpA2O0Ai7qVWaZR5yuFKQQF216
WQjru6SFxlQxKATEg+q4eSb/W6WaLrvKj8Vf1hlxu9wtKmSuYnqMwpmyYRjc1lTY
Oddf5pnEViENJGFZZfU1tLtCRXFO2IYMbJO16/Hu7JgyHm/FPHCwaqVlCSpYhwKq
1c12ab7eMQ6sqiTX1EjjKVzZbLNDOHP951xFGheyIrqm3x0azY+6mHMOBFrLO19y
hRftF3yNtpdIWySOAkqQxEn644ps6KIBKJK9RQF+E6hZERQhID2K6ewBMQOPT6M3
PHzh5GSOJ8in4+oH48831Ke1xVPv5vRyNjSUnPzg58FWT47lPhur+2Ysv6fKQ0wt
Xb/NljLHuN/GmRGzp/kEbM8M/v0inZ6qmC3IhYOCVpeij5fR0KgMTBFpQ5rstiME
6+maCARprGDrkXnDmHj4yIM/H9rIp4hRyiyC0m/7rOmRnAEWSi/nbH7Em6C7F7ZG
OIvCMYnnbxFTnybkiYKqrxjwRbMxiUGXr600ZXfmWf5my6niUbAtXshQRYY+/SBA
u7+1pZAjLswTtu9K9qEEx9wsWFo4SzPaEI3fih5gG/p9yDoKxw7KfDH5np3CRGzb
y/N3C9g6HaJjAG9oIdMvSC9W02ve8b28u6ghop6RpIjIagY2WfNHbixVnLF/BjE/
VJmZc1ClAoanjyXWtv92Qvm9lJBrZRXl9Bj8iQzLqgz1UICqYYOlqqai6Zh5kJo2
P/o5FdZ6pbArLJAB6PWzL1aNtiQj66uoDKJQ/vUD6pyIU1qXwqxVoD3P8ZV/fYoY
ULchij54aIaAkT37NpOM0r9/9sW0SLZ4YSI1+l1P240hw9XwieE1yUwkfoyNz6Y5
OsCftLh50AqsL+n2K/D/KH6oP7QooanjqiDKzz85UjVRsAtsIZio2r+xurWfxcJF
l6Y/SqWvA/CdVVTD4IC4qxqGNJ420s3pBIv7ne/PodTiWc+XyPWVFPLU/VbzMF9g
/pxcuTph5madP9TJyw0xusxA9BuJyFx5CSTv+2WUYAhBGIp5qgiBUnZN1CPdmacR
8/BP25m1IWU0NmuVN0wq2XJyUOCkXbuHtfsuup7T1j9HDjdtPtrUl83BGrdR0zjq
z0RpTSDAVYGhzDs/dZk0r3/tp44x87GfnEc47eiEK1kc/Gp1tdFW4jYYn81P2RBV
jiF4s2RL7iynpsbZqfcM/Adip9JFEdnq6+iHyi636AXMshtApVMJdQZ5DyBRrjEN
sF3PZf7uTCrwx89eoMyoK3GY2Ju5nu415r7IYOjxYmBMa8odyV6A+1VXQaZKs3My
3Bfnji5B5uxEahhVN00z8OdlhjYmliSm5UpG5e7IvNHIDwP/fo8XGZ2FSPrlPQAg
j6hqMfv3+JMOAKcLp31q0OLdh4eWWU9q2cIxFU5ZXhZvyJi667iAOAViw4YzzopN
xPOIHg0ntSVLqjmHHJ0XzvaWp8rMtmQXEihbJSMUnweAuAidRrxpiclH8Hw2zopm
tJRdqS+nd3dq/eXOPycrDfQxUBNEAelZGn1IJQD0ZOqti9moTX1v20Kbjs3TM7Bc
Zg+5KsWBa0NXBO8cN18NdSVrsHqXzGdYYP9+a/PYE5663SoXjHSmlxMbIOPx3sSu
gmVp7emsiCCYUTo6H1sc6wugZHIzgwoU+5p9QNIFGemZe1vM1M35PBlc0PAQHjcO
QLtXXW6CPdfJYArXHi/faASaBX+qlzabGeewHXSf0aoRkNg7JXtGlOKoUP7LhNuD
TZ4xmuYbhm0kQHtCM63rav3r5tO9qRt4DAsfM3vhyvBXP17s5DpYTyDdUDpZF+ZZ
w4ujVTNEdV5GunY6SF3JbZwDy+J0CTO7yhT9uynaOhYJO8t+bk0y5hnGZSwKFZ9O
aaOu5RX3MGskN5AtN0BmdgQiA8B/xxutrBnf/oEuOkE4Ny5Ji9ovXDFpJB40ivl2
dWSVCKCZ9autxxQP/PKXp9nZz6Ztk0EbKE+9qu7VVRyJdaN4vLkXgeV/8yDkxfUj
1DMDjT983PnZSGoCE3JV60P0q8kJNrn2a4/x8Mw8f6LYMzb23lS4QFE6yWTOo2Ue
b1mtuDXv5q0zRgLSAUl2LZM9wybnmyedxfLo0LL7vsNLdDUnM+HBcDuZW1j/Qf+1
x4YWPgnJ9pVEb8cAduJkFn2U48yQ6D0aLQZG3eoys0kywoxclk+b3hNl5Q2pHmiX
4Dvp8/gcIwk9e682jPiLmwA30WuuCFO5ybwSJ4Gxf7eBOGpbeYK0L4wK0RlvAbjv
f10vaIK5aNbCRWnRVUKp9njOwjwuZpXwV0VQEPZZtLHNglHifxPA9nDNewnrWDGT
sFkDa7VGOATMgtWD0vZBYdq7f6JUgetz0TkPdGaf9cq4T4iKs7cVzIq+wBLeU7Jm
yrazJjZ5ecRpMsY7GR0D6ZXG+4JxdxFf8NEMGfCErUiNMeKUHpOeQPjo+wnwiXA1
U7Ebpy8TP4ph9VCslcfzoMj/NrGXKrfFNsbXsC3WYbK7QvR2QP/LT0WiPCclepqd
+iKb+Dg4gsdMTqLjesoC1XQRL24YkUpKRUsYu8XoT9jqCUvdWOyCXGPfJakQ7Lpa
RhBnHudKIHb+0Rn5ilbV/rfhxa9znhAsW/7UgKre8Z13zR1yDupBSPqS97AUAVfw
HMKYH5pWFEuDCXpd1kJ7vBcI22bQ8XTdxbx3J5irFiFSDnmHuok0XSoaYQGPZaQz
G/q9p3dPLItuyzV5bwx7bON6jshRAW73XXjFtopZ5FVkr3H8GNmzkh9zt87Z195B
mBhYSjpsWSsmrIh3ZOr6Kh41wjiY6oo9eb6SYhQtOJZA97oTvYhxyFMhBatP1vvW
Nbv7qUPkfIW0I7UXNeCv9ovC1j7sQSrjv9Nwl4qT95hw7LzWvfVmWODDvHNo6Kx0
GoEzTYefT17xvX3/Hzt0BdEbVQfQdVy6yixa+NaDR0h8w59bMFuqLMq1Sf3tsf3U
ekb58Usig0Ll8ALZoOfvYIK/8al0MFGBtxe4pms9bdkMwM58DhUOlfXmU1o1LUTm
2c+t8cKXDF4uLOmgG7xKrgGQqvY9ZAqlt/JtH3KOS/pYvxtfakLVqsSLNq50kQ7B
M2lDmhUlT1EzbcbawVpn9+ccTurrJ95e+n/CTIy7JiYsg+5uaYxUgFNikGw1KHWt
SWB2rhfW87lkT7sgx3953Wk4SiGXFzIz0zTo9zoEaep1btZByQhPEP/ImP2fa8Sa
cJmBAG8vT2xnebdl1NyTtW1Eio7JBZwzzElL7c1cJhW7eJY1NAiulj80lwlhkubk
fevO+Fsxn7zkm6sq1MQ3JBAbAW2H/IEPi7OjBiKLw7kWod7vcShXToqDpX6iY4tf
s9EFYykZNJrk4B86KxcyIpUzwJOTEvOxyK2jVKxcHhrznwptfKEvDWMTjUQzKdDv
eFdHQvX7VKtqu0KUXeFrjiqZEL8zS+bDAvcapK+wMO/OBIFD5E2752WDGEMg+GiJ
liMt+x+ZkKXG3kqOWH8ZZevcPmFdXRtW/pMKdwUFQ88CQL/Ez4JFAmr9BtWrwsIF
vozVh47e0XWQmc1VZJWZ/aDUGlloih2MCofwaQ4SKKasVqUr0E0UHnaYu4ado1+J
NKWDUyYtijkvAgSYIDvEDoSnZlwgjUUSuuXiBmDKVFyyqqFz+OJQrx5G92rFFyHh
dgLjJLhUbboYvnopJayfrAsJTTnvRWwX11ZMDFQQ652g9khf0SomvEQxdGfJUZMf
GTeq5G0i3yIWCJt0HJ4DMYdCwg3SqPhvWQjdvhPjEpSBG4jKw8oNDr31rvZueD7j
lBzWMd03W37Ntzw9Rf5rnzsQPXsrNBrdZw56cPqd32aBHeGT2c9q5Fyalb2LEoZm
V4vIGnXoONzwfx21AmIrcjGiFDQYUGFFf3Rc6EoETOJsOjp1kujLNRFnj7SZQRpm
PEXaKQdZaohnISxyDj9i9Dpht+quMBWSQ0LFpeWxnrsxkg/I/+ICZeBhUOEPQjzu
iekMgtKQI5ijFfn//1V3pbrUI0u6Yn+h1+gUimONOmJFeMmks3o0T+oLRf4nHZXT
hsyH/wmxbyUSIqj2tS++qJRM2A77hP0K4nl+mxi9neISKc3rjdypm6pVKzxaTyUc
IwGZ6xKx8s7exZ8K81N0O6YkoZJQN+Bnvo+IqvlE9+wOJqfxDPgaIb0q8jMjDIeT
wZJ5QzKu/ToMi3f4cGQ0JZwWD7kFPZot1QqIs8cdG47+HE2wi1JMs0HZoN4nMoZY
iGbIkqq8ufo+J+77adKkkcpLNPjExsQF/lceY6RCZeOJcclp4t/JGr89lXr4XwLc
Ev9u1rJ/NUhVZ3sI1Etc3xcTyklwL5g3CfVO6BGmO+SP4S6QJz2FeftlUzIrGLc4
djgZViJt4jDpWdHmtmvtiycwJkuaD/hW9DMfG9YZ247Tnk8KaYLMnKsFiQPwXDnA
pmn4a/a7MI43ppf3R6VxZFkYJDtgmG4f18B+25QDB6z/EGXAiC2x/1iszYGTpiru
FuZLzmARqhqE0wnY11cI2biUlbob4d6ENv5pCjF61Ttw0cofimgVa+UgTwdgIjzo
ocBA9/a7mBTMHfpOYKZkeOURGO828/NZ7gVeJH0Le1QdbDNca1Y4/2FZNqBjPlM3
fKxaR22yydL83Pxt73+8akAEZyzTjz2HbMupUFrilXLpzaAo+Qnvi3HIwBkdPEuS
BI7Bl9WgNngAeyf4Iv0vLq85cVpcVPOGssCtPiGD69x3sQT5iJkfa/42u8LyaE9V
7HLW+a+UJyjsIC39lWQ7KxfBL1Xu8ZNDraVlEn6ZZVGDjVNCnym/oWd1q0kaoNU1
/DZswGvynkuT96hGk29JEVANwlL4NPBYn9LzRZJJs7OLjcK1+pBwt6KweUah1X6z
fJqas2e/B/MgTT76clp7786kVHhRuHftR/d0fE4FTBAdeSC7fh77KyrXZJV36axE
K3uRy/D0850YyvWaQSbdmTAf902FY5SKvANZxqiE6hv1P0Xo/GQWMj2zGzi7287O
xdNmZ2xF+rFlVjaZ0Nob3g3zI9yM/2nL8LcA76LT+ppFneuwEQP8c21cSVWMK8hW
VtkuNTD0IwqvdN/+FhRTgjLJ2w92VO3OknesQyspPg4m2ZQ+pnKjDZV8otVLz+UQ
/YrNhh7idfFbDt131JPzcQVP1ZLgA+/hsHLF/Rq2P0DMhUqCmkNqu1+CJRUstM40
ES6g1BmLccJ/2Y5oLKT05LGJW60C8yj55I7MjGKUMTKJ1DukSkdeNLNmn0a1r9Vq
L+4lt0NpqWkS2y1lCtwfI46Aib3ZCeCTAS7CwhnZubq2I6S/U6vX1zQPBoxW6zZa
E7nBJArfoYJtOpo10JVkUOWegWctJObGBkQupb7Z6utmbrqhwab5RW3L16Sww6U7
V8wg8qWgJYRu59Nd38toK1o5Qoj/ETzzt/vfHaiekKijyQ8kiyAKdb+7XMNuTuq3
EDcZMmduAIBjtv/xyqSlNE/Iag96rdaoctfgl+zJTkE8ABD/qTILOfBhbUYcZSCB
uexdVUfiYmzBq+hznuvwxwqdbl0QL8dR/DFFebjRgZfTRxPsbfB8jGv7lIppaMr6
/prRe3q++vZt1kxbV4Wsz9ds5BoyEdfz9A8t3E2fczwXvR5bIuXgSsYRT3g03xa/
O8qmzC9FRLcvcLD19NYRgSkbgb2GGWOKO28y8vpHFDXtQo07L7JYrJ++HaUDqGoR
XXdspnEawazQtJRd7dYzFs+FXIUcAMmXD4lAuFJR+zrhLiDWw6IKufiNjlRzU4kT
pMMXHPM+myGIgayxfiL7Pskg5eBMwxHApPCbnOnsiDH8vNwh/Dwa8lzBfwTmbSZK
kqhCvvmQz91eTsDaBgOf9UemgL1Y5kAcl74kGaaMDAV/IoPN6wCh5Km2O7HoT0th
D3lvNdtnBnDhXM8UpTkz56kuPNdy1W00jQsPSm+bnMKdkdoO109VyvMnejO8gOzv
Gd42EfesXP93J+YIatEJaRXZShPwcckazzUN/jUYAvWK4yqQEfwerBr1nsgW7d3H
g9OltlRBPBf9Cn599hlWZ5HnjEbce7FCxAtI20HA3sj8vRJ0NxovWdgXAnfvy+4d
YqZR92B4wC5R8RkNkvpcy7SyapntTMk9midmPVh9WaIhnmjtd+tK43ro/bTSmUrK
j9UXqS/Fxm2Tvikl8JnOOYn/u7AvwK0IrnjK4BKJq1POWheCNNTw7MndVwGaBUDq
mf4W1awF8/ZWYRU8Ev6MfW8UFhl3lBW4H3YqHxNVT4X4xtKqcSovqBKO2saVTiUl
J2Sza+5zV1Vvp0KKXW6dYs8teHadoqQ4D+/+vt7s2Le5dVa3KCYmb6Lxc2fMIjqk
dHL8A/1Vwv1YVKlmcW7FTrxN3nxtwr+xrOuEqaiPlhOLjfFtKBDvT9Fb2UnRtWN8
4hJaf/zDYkoPFZWSPrMnSjciSpmCUgovHoNQW4Xf4R84EiDQnp/BM+mO+UPHG+b/
4QYF4Ide7LEt94z1VZZpgEXu9L6++psR7CWCnyFMMlaR/6jO5a0TYwfGXSlT1+9Q
i5RIlDQs0JTAub88dkVXTdOaLIVmZljq2sV9LgAnSmWS4X+9dMhHyaV3sagr+dY+
f2a2p7O/7+N/P/6j2vr2ECBniQPBIbG1JsW8ayUBwta/5VswDlwBAKMuGLQuVFuL
/+taiReQe0+CAY4drLigYQ8v//lIYUKUpm7yNGmj6czsHoung9eu+sBa1y86MAcP
cBgP2PqKidRobBoIcNd1a6BgLnC/d2qdKo9B34KJnKQTlAZJXx/Jh+2xzdQ1Tq9u
0qEox3b2y8M9UQMk1WUy0TQsTnuppcTgHP0G6NsELtIR3J+XhnaZmEFcKUcDzV82
yJgbfUJWAXE4lcz7AXfjL4u53ZWYzjfZd+ZA0T4xueK0e7pSBbxI+HbDqWtNWXPT
UhwGQOg229kunGsDzGTM56jP5CafQyr1LkVzq49ORNeA91sF1P5AXW0ds+9i6wnu
nMcaIZ2DtOY5CTBA06I75a4Huf85vHnPSrRIwcVyNFneNy83tnwuZ18z4sZZ/KRH
x5hqMa8G112+uZZdrgVjVI6zwhK2FSdizvgV964zpW1Ka2x1YBYbEMh9GMhWjdTo
hUMaDZCpUTjYo3d8mmsbIFPtsFb+qcq3vKwV+xlnJGCiqzd7Unyqj4Xi4yYGd8rw
TMHXKTzYRNDWy3gCnmTd4wpoxInljt4pGMjiBvWYlpDeR+GAexU7ed1nRbvXNGwZ
LvnCCvMMoPZscgoIRflBQdCdB5wwpcnL/KFMfK2ic69Mt2JtgEjm/7vhQ+pZtplD
5sJ627+PoVRYD0udnIH8tfmbcDprAhFun7kgBsxFNq5rWfZegI0NZZWuD5NDp61r
94Gfg+zt3ODi1P55bSKZTdTq/yVYJwOe8Oa4mBkppyp0hMKsha/Fl/9alcLDR0F3
pNZaM0S5Id8yEi7aDUW15k8xsdDG0OXYxASZoZTivRp3AW63lIvBzNZHoSpXBQOE
nzufxBRNnfFxkfOjEoyEgG9fxmQD4VpsWswYJUjN/FbsVD0Kq7RnbTd9Zzo1OoDd
KKpCtdoctXpLZkDHokPyMkbsEZ/XCkmAjQw1VJ3KJhA20QOx7oHnv9JBidGjwkSP
Xkmxkp8Na8qNsgONaSIQ3mc7CexAcQ2U3W289TWCZo7uAwKOH/UsfWjadr21fl/b
3/XI3iNKuj2WI6BnIeWYzt/iKRxuuBzALyPVa6uYCVEG4fDHWmPEK0T0bubG7/zG
2aLYekL2lpLZ0yki79CmoZ5U8FKTru9/DsH7U06BqpHl/L0pJwFpgpJMw6A6sulk
zarjaW3m+eQ5ua6SR5xZMZ6mvOXA5oZ0IZlUV8rrNujh5XIadB9HaAfZewgHfuAt
qeOuUG198+7lMWPy/BdmqRACHhCzblLt7lZsGvMxOO9fWSIGQAGOb9HgZeLYoRzW
bdqBf+Jaze5ZIjBwG3a+pnUr1vKOFHgRgY8b+DY2CtfRsgFymlWyoWsQ79UN5G0q
dydCQ7KO1uLnnFkNWmTcP1I3r+aXDvRVRgN5L3a1y2idjhvEh3h/7+G1GS4x9UUs
IPzJGFAjuWWw1z8szUF3ZIkGN+SjZ91KpyIIDm+GQc32FcLFVwFks0KSeEaAXO9h
Jc1RAUoH4XAm6Wgslnha0YRfWtl/5PXmzs6H9vtjjqz3ebh9qrsyT6ZjuWEMhVd+
ZokahWQx4QZewG03Tg7uFF4fcVB7ewlMPb4KRKa3EIqtyCm21ww7R9yWyAGu4YH9
0hgQw2HPeBEh0N2reVYNqa5qbNPMJuzyhYAaPB9GjaDsDFBKTxMckg90/zIj5fpp
ZURA4ZTJ9jpJW2Obe4LZNzT7cloz07NyH0Zlu1FfHONMGjO7NqpeyOQvdqk41r2M
vZfxYPBRyu/K6Zfqz1AP42IeI3iQVe/NV9/ChMe5y5dXhGjYJFNGh2SXbMFotOfY
W/O06serZ+kgKvNEzA8xh1L8dKko/CKaVNSctD7uUFKB3FPD9BD8YbBlAMaw56BT
8f0Sz7pRwUxVwGSFwvmIbeaiUQVfZ6/MY/BatxBluSmhy4Od+VKLM0iQ07b+JJBD
tkIr6ktsqruSBgx7GWQL3lrhVxKMSksUgz03fkU6hSQhg/60AXXMiMvM2tFMdH9l
QttZGtioU/iwGG+XuJkAfisPEIqEs8o3WHGBQ6sLc9i2j0QXI+pv1aXGpagkv8sQ
aGz2O4mcbXFBhkqweI4f7uV2xi2nVNDsaIt5mhMSd6deNov9v7taSaZEsaG1h070
BLSmr8tU9a7oJQObR51MxSUWdf2Iz/x8TQ1mzUbhBuDNXHHqAp+kNqLQHJ5OBcxY
BcgWTCYs+WzQTK1bG6Dw04T76spKIY7Xvs2FMXfHKzp7ebRWFhBeH9wmQXFriDrL
KTXPF1X/4OXWy935AVmH7wCWs60vG/TapnF7VsSfmUhuFk1unNU2JL2MlGkSzH73
B43ZMZiQc9+BHyLCg26MbqGhoSnQlyljeuFXIanopTXUGW9mY5wUMQcFTnuTbk0q
z+2ML8/0zZT78QcE1mmcnmQPP/3Qd0ndxNHgXffZTRtxt3ykzxrJ1DWeg/xOMmvJ
AbFNinNCQXfv9D2OgDL0y8eybVBPrqU6tmpD8a0R+tooGUq7FfQDG+a89LFW1dh4
NC7CTmiCxsFHkw+ytZuOmMt3PXLvomtbO+ZbTgkj2sWY/wErWODz807NxBQIKZxT
TTqeUWYolJxRCpEQsmTZ3ksW0xp09gsS5jNNbGCh0cHFRxbPokzik6iLUg/f822k
imdlMJ71Jn8vEFLgEwRCelsgH9DZJEyY4Vj6nM4FyFFC06aUIDJFY59QJkhyYQ4i
jSbCEglxeZopFKtdaGuwPCax4jfFW7oDf/gauCxY+cfaQUYSg624jWT3XKF1OUr1
sZGSqTQJkx7H4jcMZGwWE7RrRlqdxu9fmqjTIlRMwfi+SXFWJ1uN5GSuXja8TSC1
YvU6VN6ynjFf0/p2GaX1lz7Ge673wg8UcFIQO6gDUmTDF0fciExieP3edHtDkowO
keJkOUtXAzS7d387/f9gye+h2sA2jh3I6XioDfT/WilJ2SxbF+vcSDObqnTgxXC3
/BzFh3TWXdQpd8i1Ne1uUHewGbS5OYCcdHrgaxw0rTz5j4mfP5S14Ok3irUjpe4y
+6aNpCCUq7vHg9EKwGieJBS7Km2Rbh4NMnW1qJrfAcFZRv3VjPSVvwNsEy1iycEF
ybI+5LtmJfsNi1/xneo9cJ3hqb2YDwYVaJE3UIKAX003ZTm/OQKRy+yN06lu9EJn
KoF2hbrWByBFHmEZ4SK4sfcNV5vTlhQ3KJohu15NzD/WjaoeDR74mIlN5Hk/AwFa
YqUE4k1ukCU5moyOrPt1OaEAWaUHrHQK5cheasjLoPjX3W+F5vIqaeEJun5UCp2x
hfyqpHzQRnpJgSchi5uW3Iqr9SMq5v/TVVUPmuNIAqsMx11vyfXL/VojVFRS9Zh6
SxiEJO1klNy9QcoXGmtT39UKOFiHlpRbLODHt34MZCnBrqsl9p4S9g6MBA/eRQ7Z
Z/h0vSFZrFXZXMS5cW026oF+VLeiXFTIyb5PCmoAKJhChjFyD3mMQ+PGD/LRXjjq
LFCVUvuRB3Pv5GlEKKv6+BKDdhFbTZrSTsxhGa/t4kmon7uaZZmBD/t8hOSnR3AP
SwhVKEJS05YyipVT8t6odA8bAYF20c+JMWAEkSYtU2N3UGynPoTGAllJOsLj5s4d
cQBDY2vH6lvWvYIoGHOwCiwSxqGWIZMvwLJht0X0ke4Rqs9Vra0fPseu1bHWlu7f
cGAbV4/m01xNGthVGm/0PMAYpCYuJ+nH34qBJ5yFkKY7z9VSMDyGb3wSMD2maR4M
nhKRbBjB7pzkI3FkIka37mY91TYd//l9krL6BvGrbYRL1RKiXbQxuRS0Np5jYRu3
OpCtDi8/8o8S9hqP5ei4owSuiF05ioLlvkw6Ah3bWWENr8i0xUD3hbDFRI0226S0
WDpS7kBWmfKOVzfARO9zvSyaq5AzA8JwVyP/9ULXxC0wRW0WGL+ipq2GqnnlnqKD
7cfCj+N81qdtA85jexGqkRU0aGs7/fFWEXi9V+Xfn6Nr39MF6cFLOrvh98yzSz0f
ypymErTUV9a8ypwjzOMHpTCjaxQk7mGJY1wBeeRk06kKM2oadCNlA5mG+BgwFojq
AZf61IAWnCzSGT7igRZe94HoHCChK+4ihutymv3cpbhrxnNVWiLqT7mGFVrGgbE/
7DLBF6z/f3Mzcn4QFy88RgrpD7Yu17TdH/YZrIrhJ7MIunvrDB6xLNTMfox17Bim
GrCd7x8qBzh+oKxjsj/OFNaVAEryjqXcwZxvvZ9bRPePdrm45/KTResqnbumi6eh
xfh5CWoP7R9VEEHzJxp2EHcKzC56WEgSqMix0rpyzXULjeapuI2HWbY/Fy4Ge9Vi
9+bcOor29KWB16iNz4gNGeam3Ke4SMaesj7rrGgoOedRydEKjQBJBoDeLKhDGX7K
fVtKCe5aOnmc42v4XZl3mQn01SMb6WpENXE/0tmlzrWjM9tRSuXpKzDKn9J1Nvjw
lBi5goQtH14yuOCY1ckPR4q8sPWt03F6m3ZT0SwqsHiahpKnIRrK/dd0ft2rHe6t
QYeeJ/BpIgjTgRfjMNl0/J94xFME8ubaRnZ4tKYRDAGYQNiPb85HFHz9F9GdY60N
xadIFJ75jIkwpLQUrgQoZoDtsdKRwuEGOYc0S2Ci8AnGcUiQIkNIE6OQFZpmGW6i
tb7Mto9tkqrijuYLX4jwaVxJptp5urFEgeh/wYsg38jQZYfwCtkMbLp1A0iLzEiH
tRyzW2YWfgwaVomU/IXOIfTYO2J/i01gaPDgJ+2cj3oQaau0bjB5KWkEdhIitRR4
51ycQqVZvjPDv19TlDVvPKoMaOjhUj9BU0YwVFEWrrq2pezFyniFcZs1GmqHe5SO
0e0q4nKcyZrcReIWe653s6PW6vxKNQVABNsmMnIkeOXcjLSsNq4WGzrftAMKoLWn
SUoFWMaLP+uN1Qk0kGY4XBIWWWB/qc2s8WSI3IrCr0E3tWTHAiPgCNDenzW67raF
CeSihs9o6Vpk7fIe2F3C25nJ/Vb8uPpaSHmpGD9Rabui1XzM32zIrIibqTKH3Yl6
u5gsJUQzjF7fwiUqyFnWM5ta5rclDjv8pA0mpsJK0dFgWTukTtc1vfAiDB7E83LL
nruf3cTJIfNjQO8Da4RggVicOpkSH+Fe3VmdaEAnpDL4xq2c21iyQhg3totTiSjn
FhZsrtZ/qBtEzfA9zqdJSLC4IPnMfGUvZnTuHsCQWHm1YUO7e+64vT6I+K1OlsJ5
BcgoTIfuOonpsvVVAQFAV7hANRo1t5D0rfFShNHsjfEjE89zLB431zhBxYA10Auh
B+ha0pBqpli3BzL4eDY6L0L0HpKintMxiHON1ayyhOYN6+ij7Xktkb3cIdaO/dB9
Un+AiY5ZV5NViJzJBAwv/hOE019NPB1Z/mQS4R6qh+xRO7AJo76ZXpbdk2cf7WBw
ZemnmcCQZQfid8932bFqFhuWDrbLr9tlIzDxoi1/nSILDkkQ6lToE4IYMuij0TTz
a0tlPWIFF3IQ7kPEuJ6P9Zzi/tPK6CYimep9cZNnIYgX1sb0WnbP3S+rOBT36XAo
mGQo5/255/0AhGPKb5syo+cPkmvte46rnPO2jO9QND71kM2Kffm6aGLRrqCkZVVp
ATLOLy3cL6epw0RYrG9OJS8k8ZvdRIR8RbGAIb17T+7PKXH/rDPOweByQLQpRsfo
X8CsYlId1H15GfeohPnEppLtlRV0s/yKMPjoHsKRwx6Ds/aPKaToqCkAu7Wf+aQJ
/lTTMIPCOhehsqdv2MUkaYvkHyJzwYBY4fzLp18/3aGnsr6hl9+DDt1sMhrPHLKx
p1MJNJn4efAd6f/OHjBX+EMRUbSrAaTsvyMmIxqIUCSwYqbsdSFsVAt2T9F3srXp
8WRb55yD6E9HMNQuYhpAeBmMqt9UfDXOyROMCfw/mGSCvqpIHPt2UzWe8if6xXY/
8IBY5nn/m0DPuBVhbLdxgfEIpoc9rglZHKRNmuSSNlP6Q97dXdl0DZHAyaSQ28Mp
BYq/Ec5zEB4Z73PbwBCasW2ehFyLCDWaev9le/QkB7H2NDUWhJZDvd/2woLAYP9j
YkkpCVWCXtrSDtkYKys4XJ8Xdqz0ohmRIJWQx1wgip/z5x300o/fWWyPm+BmFHD6
a60SGrYcBRauSDbBS21u5oTjJyh52KfFBAcD2aHyDhVUiASpBaMaRKZZSMZfKbuh
v+MeANlPufpOvd8sNXhIObecxv0jYLc2U0lJu/2qiLnAtWX/FCZvv81gRQcr/kLb
DeDjYFRrrYWVropULAD9a8UpPN3X7yc8NPTQetmZAwo3xhkuRL9R/CfB5GqMoC2A
kYJFWw5isFwLsQI/D1xyebu8XAvKLKqkn5wRhD3uEA2nQRXPcguIedOJqxnHz35S
qdsDtF4hzcbO4/rONsCzwLVelUOxmlm+BSrsBZz9GwW7vyEkqH2UDejQTBr0y2hw
8gt4EwfE0pnYrMJKjw/Lri6Lsx2Jk010O3j6pNB2KBvoehHaw0RUyw5GIjR1VfVn
r21DWAd4MjjKJxBsfcPAddv9bme+DLXRMMaeKkModPWtbOGCfwPMNUhrO7zI8y4a
H1l4iqj0SxZctrHQWfAdRGqy/wlqCwF3+VfTnsh2+o9WkR2QRsGDuDMDMKfg1iaw
eeSeGydNH304XxPX5nhEnCJEolUpM+lTYH5Qx4JDwcP4V6RXzl1c43ywUL/NMuaf
A/hbbxMBgsCDrqg17yTiaTI7UU/GqBpNWMUxVThbEDHpYEcDsyIuzz2VoDXwJQqD
WQc4V8bVO1BVUM+DSfccwbA5hGO6SqJC3RzIoBqbuTsQ2HR7w2afm7bp9+mJ7+y4
/5alSX6lnBDCUGR4C1zw3/2VXoixv3uMYqvGTkc35gqCL85ecqAuE/4fMqD8+898
WbVqzwUzT0PPx951mI9kSU+q/1RUkD8sEMtZGEwc/po6rVWXE+8p57v/38seqMlg
RtzRHHcIhXF7fu5XRqHl488jfIax28ziJq5sxyM2bSaNdQRoWUCoatK4R0f3KH6Y
z/IVGti5LlkX1yBDtlwYVQ4cKGblCyUMxnLbgcX9Kjoz1XKtGaFWp+Ob1DdNnThJ
mGLgQ560fCtS7M50gP2z39r5dnR+CEZ8wM64lj0duNKWaIPgMw5aU3RVCmuuHfpl
1D55FWN07yyr8xirQagNxAa/aXnC73KgSk1+7++OuGEQG1EfYfL7rnC0J2epkPvE
8y3A/vijML5yIUqqlZsN5UhV9nK0l133EVr/ONkDg4jf3FuAHR+9tI+pxxzP+HXb
7uUowa+qrxk1cDyo6qRUb+VKw4SB/LshUT+mAJbL9LYApJFWm99kIyInmf25v3gI
cTziN9bRIsTbhUbi5qwuvmhlP95KxPMIecWybf0Rl/HeBeqbKobcRcT1eJpAX9Yy
8uXly+eZ6whF49U/F1fJCpD3bo9zbguR1P/wgMR246mXfGaLuWbME5OnwlYOCjwO
4Eeo6hamZ6qeinFSuFDaX1emJuFktPzJexB5mP7d84wKKUZ+DRIR0LQZnq0zJWyp
sv48m5jKbd+/h/Cao3g0O3X5RAPhY29We6o0U2fe6Uj/blFX3+t4nhzFFrqLZreP
LVc0U8GPXD0cMxd42O+nMXTXXjEMNTdwZ0qHyvcaKii7jNGAKUZ4F2MNl6sy8TiA
a7WGZbWAhejWq0bjtSpCuMNJZRvxg6QzWWdxs94q/8Jw6mJV1PcQTr8Lr3/xSPap
u3JO/yX/JQC/PJ3zxOQsM07T3y8a8NfiUuyLRfMoFREQZiOyLiDMj6UYkrEAl5FP
326SizfvLRjl2OiEKyiaErIfnhyKXo/NQEpEhFZoR6ABqK9TDDnHdcy9BhQiPAw4
PDK8r+TOPNgDGINjHEbaONbxTcgmOdetL/kaLXK4BCTJW1oVfMNXZSAjfC2yYOAB
h0QczvBDjJRF8HMCJs4FbNVcPWnUAajdx3j1kDQsKxD0piF+dpY6t/LdO/1paDtr
5e/gkEBxQHvtcyHRQNE1qYNBhcHwuG5B/OlPhSnp3THN7GeLQPvmV7JJtyBaGEKx
0qU46tkNkC353Am0uzi2xMhEelWss4zASujkcigw35mgvc3mAfWHRdjo5uNkffej
Cq3zcA2fyth7ONEY1sozRJZbFeLUGjuJzbCjFm57l05yvBB78hBsgV66vyIBKd+k
HhX+L+A057v+TPy6pwe9uxj8N5p9UulMHELRWSf/mko4kEiv9FwMEgTIRwQBT8SZ
G1uN6c1ArdcJsLfEqiX/+/7gJkR1E5JCvXo/5Qy8yBWIugl2Ubb+V0JvzPQIawzp
GMZHEWlzkPYE1A142zEy/7ZujopRLpfCcdX2jlFdif6eWw6c42YE3B/sj8669eim
p3MuoU6b0OctKfUE9IDMg24SdD9bNzQAaom43NWaxGQqa0JidCzaKBnzErsBBXJR
Tpt0xS30EcKdlHbKH/qzjbve9grs4VO+pktyGDilOc5A1R3bHFjl5INlDw3IFWN+
lLL6XmrZe1OW7161ztLTPcvRFC45oJ4qVC3DL7RVnZ+veUOsOiBm6vxzunBGwlS4
AykHgadY51WItvgzOsmcGDnWbSqyDYltwHI+kIRSQu9LrllN3ok3Gwuy7ju9itOM
TJXySyKTkkxdi1IgY2nx6bIZq6nCauRjfq3TcNyYX/oTnjnBsAz/W7mj2jAgx4CC
jBOFzzUuOyG6Dk1gkDOOsxUCzjluv2dBjc+QhM/pFcpBz/gX2vEY4hRc0u6DeKmp
/VnU0kyMEB09XeA21rmNSXLeamGCD/Wjpwnzi1KrjrbY4K2u5j/Qd6vn6Hcyy1Au
8ty0X37GXed3+kE9xNfHmcyuufJ4jqYr2T3enQUD2xTsNm4/GAUOXePgpIRGskCV
rWpVHeiJDBjKta0zEGZ8G/Q7o+yx67/sblv3ZLzeohehrgCDZUKqxd9Q15d3lRRk
N2kdM6zyDRJe1VTLk2UcywxkWWTj5UbIlQZS1Y2rywLpq6WAFFuNE6x1c+c/ZzfT
0kTAxO38xq2f3KTmH5SDG/FqqPl8n04vxWHfhLCqlugBrpHekA4ARH5011t5tSZt
bZphMGXTJHGI0exPLCPaCsnLJgmZ07gDY5ad0/xuNnouii5Ox9ZJROTm9fv2H1+j
J8DWP8BEOUtdsUKiH7IYPii+qWy3mF0odKTn0d4+G3cUEzEqCh+c057ZvvrC92Ly
FOkDcUUnD3cZ9MzsMFT45m1fINIabFLk/UcaGppZIKuuGRfBbG2pVRtsiK4dmxkI
Op0KpkuVX0z5uo+7ieagK9z+NT57gIEA0zlFK9vULnqJqoAXwCmJgndUDPU6bwLB
5SsGZLzt0qmRXkprApT8TYnbM5/LL+gQx02f2eZN/EjcUJn13qLB3/YhbzWSuJmO
9Qt8REGXL/ZOuEvlWyFQYt1gD7ec9DBQwlVZswhyIe/wSPiVDV4UIlu1cMeGmX/8
DExlB2Cwwb648JIwwGYIMIY1DHUuClRHQFwpfG4oZ5jTz/ZbWbosiyEIsxe1S/Wh
W+qqwmYfgVirhVm9JiHd7+X07QHWl/niPxoYz56VLIUnviRdji5l+k56HtlA6qZW
NpWmrMJipvvG/dwO0qjRvAq6U5u9lGUV0GV/cl0xVe8LgYUF4UJERFfAgvINhNCl
wKGTknBMkdBXXjSjeva2ltyRVgs//vMfyar7SpaNyHTvQL74hnX0KGhyge8v2hO3
gvld+jgO7ny1vVyv5P/KZ+H1avo5xQ4EGj0ySSS8JathfMsMZL5M5GAHyGksXnJ1
K5kLy8d2qYWZ3aqWcD0ccBGdkaJCpgnagvXS52gl7o+Gd4r5aIQLWZ8pw2hFBPFU
svVFLyL8qK4d2tJgDxrfvtppHw2VkjH1wF06Lh0NIvfwhQzrwlk6PtCnikzPdzXf
gSRfleyxrCKEKjZqf53lAGjFlvw2eySAz7+Q3Q4k+zvB/aDwkh3TwUYBGOjcn6sA
x+x+8oDs+qndcgzA6bFdxSjoZz8JU4PG+9j/B9fDLpHdYcymcPGYwOHCjiMDep7C
QsWBpYYmzFa/9uoQWqh0yo8Gx8E0nBjNTn0Unu60WGHiJpYXkmUzwkoXpRVwQh63
S38GUk3iNsTN2CMWdlx0kTa87bzol4rHeRD7b8bq/XBE6s0lhcZ19h4zunGD35rU
A8mHly3XszGAwuiLJLK5HxA4z+pxi7u4cKUSwPaQg6AM0QaXYtY2QASGVdoKWYnX
QH2mvQFPUNQno64GynLq3WE+39rLC1EPsZIRvPl76uKtCLjqn77lkNAMP+asiNja
uyEuwbTg+lUMAUPoX2bOZKBQ08Up8RQFKW2mQWGQ5mKxoKX0zYq430D/PCfRd6VI
86PKQAZyyBqIgiPxrkrIpsA7uHvvBh1qL+RhfxlX9Uv+ecF04sXg7fNZ2pwLg4cj
xu3UBJBura8amml47udrJUUowLa5QXDCh0WU1cFvRHFBs0tT4IV8DL6bSb91Jo1C
vZpH/B0Ro5d9dA1h/i6guCWybfHCo9t4nv70IZ5iYdxGoSMhONGYnJqUVgUloMJb
bSf5JGPo5YglyNLfaH9WScSXTF1Aq+dIv6rg3/96ceCYiSGALtPC0JJgreKyrvsK
6NpRLH9a3TsbxRBltWlaigI7nPM97G29TapnGqqnMDlX/wSACpD6lnlbUsYjtEPv
LIWgQwd+H3H0w6IH2VTlDL1grQ003QIU5zHRyYmXgZDoCG897JCgzuY4tNQpGJcb
+Mt9s8stcFd5sLCJcHIocZK3iwVcOxNpORrohfHV1f9CaurMpJ/iuXLOkAszfxso
R+F9ZBc9Ssp95MMK6nla8/pyyTLiYsdhnZ6D0DsCLsl66ShHkm6Y4NqJMoGB0Nal
gtyPIrMjzTM/VKgap+Eo4dqxIIyHqhWBxt0lx52C4AGeYu8j8nbbGtClnPSrqmDb
W8y43YJzSzycnuo/1vf/1p7et26FO/AJ+rBOxhSdSQTk9nXwkT7ffIKU7592FmR+
gAE5t1P/kTrTJyBmSxfEDacLz164Yh1D6tovduS85ukdF66CHjIiR8TpyhTH72t6
2L4hhjLjwZzrDk7gDbC2jBFV6oO7bt6GWYGa15nK17/O+LDBiew2E+eJUwJFqkus
+nn3D0UZosdRGieaEm+SM/c1hhxtvxL3KSsmAh9gc9vlwadSGNt95wxNIDGRgvfn
IdWzJ/ay92NotcUcLITCbBQ4kKogesHZzjAVDpNfb0xb2WjxTlwzAvUZXntU3/1C
TE6CjBMhqMmvQREbynwGihSL8X1w+JryZRMRNhTKfvFihdCB21dSsh0xjTtL58X6
zpbt8hJZmnvaiJ+614SwjS1S6JypOax4GXPipFHULkzRBTxhNulz/AcCVEK3mQVK
gnhut9Yzo4FIiod6wq3cZt/OQ39iCGIvQW0Vb2TLv8q79j6QX2rZg0RdSWLy8ojr
LBzfHnfO0p+n10QcCeKWBbEVPPMqL4bmyUYi16JoynDxgnhd0Lq3hsKP/G0Hfo7Z
o0qjDdPHPJNgYXGuJ8x50QmYn+lrwg0KG5ksvTr8b0JD9m6k0+t+wQPxH8rlJBI2
Me8vhuTP8+Dy0rzLg9412XhICVDFnTM3h441ffBj6s7tGAwvrtxE/XGHffev2cNp
vvMazDlPtG46iJlixJFotXeSNITgS1duKk+RtgRn2EpSMZaSWSCDetUtVcn/bR/E
vVXXWXP89tyoOo+5e6/QNeFSGkSXpW5TayheLJxSxhqsyNNBAcykbFmTsdNyhpSc
m8fYy6YFJouNdRn30/Jj+eSPORVp2hg66+2k1bCAVOprL7u1itlmCz6C93EivJbx
ZfPO6RozaBnBUXrOhCNDX0qU1DpoGjA8X7X28O99UokISG+jfmI5/yjIhPSM+aeO
zY8T9lbaLbwTqmPwD/5PRH8no11Tc7pBK3KxkxM1TrCsGsA1hamNL439qcF+iCox
rB0UcsFplUHNSoIAdsNQsNA7f6V4GcocV3vbsIsG71SAwqVAAry5kXt43UBJKDWC
LaRfUJwFSgD8Ge3hNpyrrhjk+pE0cjSm7weMNLqMFE6ppR0oEGK0QZ3HTCybucSv
bA5ordaC0iS4imeypPTW3EU2B8TL6DrnfcOMDeZ5+Vy9kfqX5SqGvUu0VN2nJEzg
zALZBNpKp9MUfB9O2ZPR/VOcyLhSbr65v6xu93zBH0X4qGP3hlJy9Us14vkwbNFb
j5POMBr6maVVKdEEeEFp4tnm19U+w2SxkQfpnKdqkaLKU7Tv4y4W7YDeAD5bq82X
XL+zyT0hjF68xHR2eMGrtJvndf5AhCYyyPpD0JJYrUt6q4+1BCRITilHUj1cwcyu
0wPX7ext5S5uaFu5aIpHc3rj8uf9zgQ6YPP+pJ3+/yAKN1HJklLd4m7W7YnnzV0j
t8ftf9TW3pjEZleXlXokbXcznFZ0NLEkmtgitfVri1Gm5w3kWkbJMCYI+0jgQ9r7
dlCl/a6q+4VBiYh+18OfVo+j4e3MT7AcSo9/CVKZqZv7G5nbiqd526idOmNHGub3
yoe4yduyVsiEyEJsBHRMo5bMuzUAeCkPtU+l1MQ4V9jvYfw+oXhoeIczHT4CIGg2
d/B5Y1YHbc7bhV11GH/PGoXCYYdbi1iDZFIWrtMStVvpOVYtTFKQORvBLTGVBeYY
W/KTUDEh7+8YbYDs+bFZfLk68l44+dkAGdIueNPC5Rt44I8pw+rxPtdVThsGNuQZ
gpOYWj5XKB19pEbskT8pNz79QA/hb29jPPNQ7hI6fp15p78M3FCQ5teRXeHZicCb
d/pprQ7WfyzzbYyitmn/S0r5xkOk7FBZQhM6J0k1tE+9fLLZTVa+8i0eTuUwtlE5
DV5GcCQn0F1axtlwoPj71t6PI4reNvo6kpzhGOkqECEvlmEVwvYQy+jv7yrUCHcb
RGOrkB/8Yp+cLaAlVYzj7cg4j8KAFIhvpcIOo0ybkYwHOJdDntpjb+1dRuSoR3HM
XZc+UymvGq7FHP4iWFBxhg2B6mJmiiShaIVAMlA8NpGV6vNImUpnX8yru4Lh+Ab4
xEEawse+iBi98Ze8v69mxDZDXIXjR/MSo+Y9btytDrgjb/oT3qMS8+EdfNlR6Smo
VYN4klhZ6ajk/oNrvMZWjWQAAqx3rkj5jqvn4QvhTIgk9NZ6hfWrtVx4DLzOWCJT
GC1UwB9+zMGBd4Qws/VVbafwhlz8b5fBOpUAeoA+IFfUW4rj73QqJiAwQxJRbyTV
RUphKdCffQKEP715KBm5UVB2MdM1KBRhRUwbHgu8E3TCaqh4UDYuLRCxvIlaBYGC
O4MkCZlg3FKzs54GirM8odV50LkvHfqvE6MtUW8l3fltl3GO2e16mNrjoK3vw2C2
RbwJ6LfzShtb2hpKcX2jsh8q4JY0cWXT6+00iZgX1ps/5MiEYUh0Omn7ozIdhdE4
lhuDFqFcSXqbxolDsqsmh5zNpQWv9MKwetVk1KtK8VwrcRyosMufoMMw73mTvLPM
3IyKv9dsFO150HtVJAMAbP0FXSPSX8ZTOTWxGnqus1/+JJRLCQ92TBOankUhTFLa
BphZv6gybzBd3tjsMjIOrHPggP0F/K50JbZc+BLmWGWQmaTYX9EqaExOzvfEDmXP
xKtf9qtei0h8eZQJPph0Xuu5s2CxT3epZnMIr6l1Zu9AZruM1gYf4qo/ki+CMPtU
JAnZ654BKYZQLTrZD4QVFYm8sGy2Eeu4P8W00CLf2savFa2uVMq/qfz/Bx9jKhTm
wcuAeUDY/jWYwsrYg+BKnPErK7XoRU65Z9eH4U1Mai61EflZObO0jiQ8NVTvRk5T
PxTEiwFHczcUjdWvzEIGS/R/lzQ9i66cTZUm5jfijybOx/1/SYo7pg2jealsGvxZ
YbvGFvis3hOoGs4PODXDrIlXaolWIhxy90IDMygMosA2pft+qqZzLzzgzvGhXhj8
rzv91TZNZY1Zypv9w4LfVtihwoeRpcZN/S/l9NgSnEAtAS7n9b03TTxRWQdl3+8i
ct9kIEn/48HpWN8t6tLpipbd6A7KeTHTDx4yX2X7voRr2Q+CjefwfoaySJXjvXEa
1rlwOWDXOrEZKSHAGHgIvv3TlTg9wSBg5Mhvd4TP7qgDJwzZfw2giw2s9Fll8gKI
58HVTjDPxg4FUuWsUYWAh5YnICIElKXm73T7TqWNjhooMM7wJ+Y6gGjv0UNw1L8s
NEGsOvxWDFqljvDh7JyI+EuifwbiIsMd7pX7wUTgdbSIzIoa0nCFxxHA4eGGj3h1
/lv+xMEMOyuvDd+wn/E+kuc57di8K0HQlEgrEBrxBUSAOHMQLx8FNhC2mJswtxz4
P+3qR8qcddc5eKjVZV5JygprYWPY3PD2l6pjTzZgcUAD+t2Ft4CByvRP5bxA1xwH
nQXpC4IXhqF6csrZOmpIKExty0FQibQefGnsMiKV7vOrZijrBNPBgduiiWeWfIuR
SUSXXGQt0EHrUu9LnRbiINd0Y5nKq1Pq9LoPehUWSuB20ZvjfIiSKP9ue1nKjxvQ
NYpQkuLe3Zyu3K4t8KLvTLK+nguIUCUbND1X99TE/RZfbLMdAoN3R5wHs7z5gnug
iaIwWVwj7Rv4pMerIV9punKU9FIT3B4SZlxk24GS3VFNTpPMlZsxIwXm1PRjWAim
fLVyTnT5xHXspANcgXimM3DCVigN2CdGwiWU9lUnC+stva5PohOxLWt/Hl41zuUv
B4SK1BqLzTUkFeGDPh6lnT7/n0Rczm7FBJ+rEwoPpdRibz1vrFAwFc7cOaJZkqH3
m1kXH5yDZbSQ0mUwFmz+1Ayji3C3Epxez4axjN5uqkP8wz2pE+CdFjqcmeeduP2o
SNGKMmjBZryOlLch5BhuAs0cQwKAMs4nDclnt4IOm9SDm6RQquUzuN+zkg1jKTDY
o7EVXkGOfpZdPhcMbT6ByQQWHGHyjDy3nyqo2U27/RnEwxFl60RTKKh2CaKXDWJv
QgVfmxlD2Y6wgS/kYoHMq/meOnE+L0Tudygrv3775xXDDo8ADOhfWyRwAMJZwKKX
5DeAolvkSHwgQZFk5+n4/YcS4oVlGwNGGvxHu1apgDgLdKjm5WbQL7or2fc2DIW3
GZ1ozV8P9OskMe3284qXK0FCIqS9OlnmnrfN6Cp5nrfsVLqPXB8e4c+/fjV7sxtU
tCuGtuFFki1/wKkt3QqSyEY8PoVvFzPk/1zAPhdkprv7z98TvWGiTLnniA9RRL78
1biar9y+sQL90Er5pxHG1m1fO80tOrEbzL/dUzKCZN5Nq++TmtnAuEXAofMAtSW5
rC0w+t75RbpR0QRD12oWDb4K5aGkjgNc70nQ8dcd0tkZJMTDtv1hzfYbNFXJCOYn
onPrB+4vRjGeGlH9v62bJ3qntb1rD3daS1mUFRyAi2G5PkTgFzJ3hKxLsiLDBMcF
PNw9PBeY8TAo0tpo78Ag9g7RKDtpZtKqY6vxqNduG/Y4L0qA87I15i2UNL04u89j
kXfKz9+l3+LMa0FCHEY8PJhnUVZ1tM1+sSo13mJk2ViYrf3H3Fl2OhOfrfSRKfYn
Nd7MrGCprnYYJ+FG2ZCKXQtO+GQZx1F0D4DuSGEt8hs+zXUXuiRVkYsRr0dgmUFO
K6y/C09wqC0z9rnXUzuWFRZkYmkhUfAgAn4Feu5W60YBRZG8yo2ENM0Av/RZxhrb
7fA/u7MF7zzNJrC3V6bSEHEFMNODbH+SJrdyq8738aM3owVh7VyY7zA2kQ0sGWcL
BdD0w5/kBUosswa1N3SkC6+HbFIDVvAYDs2BQILCdNhuKsM+LlfbZ5HWZawTwjZ2
k0GGhKiJPMW3c+YZKKXtcj60yfsZyb1bJDKlRLaZMDVOzfD/t3ebmjSQ75UroOHG
ZhP3pFDa5uBGafg7gH/FljIGVOclpyF9wV5bQo+2JXgSXR59TCsM8J2a9SM3ai+T
ctz/vkjh4YHjnBPkLLTWKjSoereGoa7JOLNR8y42l7cOeDQN22a2Al2r0f1rOO2Q
gZOik7Z2KokBQ/ZluiZ5NLv2+FEUsqAn/rSEaRJMBlP0tn8SdO/OowWrB0xDqlGK
AOxPOTlRoHnmPJqv8KO2n19AAGMavtA/+a4jyD0XBCyBH5jQgBkrvAu8fW+RPYXH
JbPfnxl4rtqpUJvGjRp3TEmEaiRkSlpQSLHv+O3W6LQ3scLOwXTd5TOti/J3Cza0
ao0o/Zwc97hS+Y2rtkR56+NpSWb/h0Tmrcrv48BiiSAeFEQrOneWrhrfYpgVTVTw
BsHuRrQnYAwD75YpAZVut1RHm5szW5BzLzqk5TolQuSUPr9CKSycRcLxYrVxDpbG
543+eM1vvd5rHd796Nt2outxveGvCvt8E5BVQQcm2lcJOEwKbg1Ggfg0b4NZ3tDR
G02tGsTBKBUFtFlIDBq/A/RtRbxRoQrOiadnc0J9gosPwBm7iQIPMKtqr/B7M2uT
EK6jgZk/d339mJUky4fox5+V6Jh7UBEkbD3E8azuOQ8pPD4bWwcmEIhW2MWPJ9x7
6Q9BaAR45QToUeoc3f5Cm/dKqum/DyH5MsXgVWwy1jNQGotocTWrs1JIKGez6ek/
+E23vqozcWVHuY71OjnCdlHSdlQqg3/JN86VgbbQvKBPSDHRJT1wk/+eD05sBKr7
CbPIZfKrdoDVWAZtHFHUgXTDQPkedKZxzWFNJq86DzqBxc+ARnKbf92BnRlnZKHr
9zDQOmnUIZC4ZGcJucEeDCbR0Ihp5IrM/trp1N9wflmMJxLaznyRRbH5FPutluc3
+k313u9XxR/k/Sxx9YrrcM0aN9jkLLFFEIVcUxKfawwieKroWNlvv27dF7/CTCB/
5mV0hnpXHscTGzBl6wyY5c2JbhBQIRRP0Cr/CsdCOBShvWRQXkp06qRDJuesDHS+
1s4uJxovJSb7+5kgvqUOcUaONXLT1YCPxLyIeRcfyT+Pk09dJ0lXUQ29WoLLATh8
UuL+BL5tl5/lhojwB7nWuZqBkmuZiXXZhC35wcMPBQ5JbqkxBORZoKe2h2c/C/Qi
ILl/dpXfRjvJJd5rxRJnHm+9Dk+gUhni5O4h6ryGEtbLFXkPyAUOBRb5zzK9Wd1l
tVL9q/90YUId4PTm1X4BtoE7YHNEao4RMcaIcLUY3lSL8Gev68b2CB0Cng+/Eg6N
8Yoy/8YGcfFX13PMYcD9gnrH7AjqbIiPv+iNRqd8GEMIzRCB21B4s3/Zylbxd38X
rFxLk6JqfJ1a+0C1+bfZcbTxEyW+BjqAr5UuP8ZnIq8jXCYvM8GPwFf/DfxQYLa2
vnetGnWrk3SWCkHTtSico63oLLphMgzSaoLOatKtimaHnzamecEIY6dSMNCuaIOx
IaVnbbdjnPRh9uzuW4zJmPiLj6YSpYLIdjYBq+IO+FFLhJNlaez9m2bsTV3aG8Y4
20HxN3Kbe0B6d+jKgIoFDvupQ67yXML4wco0ejKC0T9LXWbHL8LFJnkK4u2NN4Qo
RfaYYNC6b6xIP7R39kIgclIKSrNNSxqjsi2emOJWgUTGcjbx9GuGf6XcPJbPbWxd
Zm7DF3/543v4B1528TWUtC/h5SFJ6FRtUN73b4TZsP4PXj9TefmVQMS/Y1l6cgPw
6TMiZ9aJ/CmDL+G/EFNEW0zsdddWPFS1PYJgf/0I5S4GzG2LQCybbPPJBzh7GGYh
vLFsePYos1gLdFkMG7/8w8RtPa1qQ1ZKMc0OzSQCKgBMgFEn4gB2UF0pa20gbeHX
WtH/3/CIEgehObEdn7m+YWlr72DDWu1MgZ9eLztkoMenHOWh35LIWfhvnSOb+13Q
izTNET7y8XkBDgwD44fFPlRFnultCNXYROGoQFA4O4Ox4N/ORzV1Bjbr4onhosxP
U1YGolw9riEl97rlCngMdXtqX4Dg2e9/Vx/KRcM9ZaAXVeO/2Ojj90eS38SzG463
fuZTQD7QcUKLnU6D5/TNBh1nKMqVIp9lXwml0VB0HsHd+SK3+Vamo1nomusk72vL
AIq+ttY1Dweo7EN+0IvjDBWPdRnk+qWNuCPjbQZxA7l1ilpsDmp4CeaoQSi4xhvA
bRW0bO8s42QO2o6wag2kfWGhFTs6hX6THx3xwXF3PzsVVF8Lba+VViuPdPHkt1u+
zuaIYmAy/RDohJHDINbjaM8w1QPTsgZG7XeTmaVlcsZj7Yw7ZQE+7nywt5A03Zia
9e1yVr27EJ5y3InVxdVH9JGxwkMi3vzyzKbbaUzocVo5/hUROXoKFGbpjBvAKJJw
mgfJ3ODKDonZVl7Zoa0VQ2ojTPQq+FyOvbKsDW4C1xUR2REt24g9HR+HV62C/CfW
fhrp/bDL1Ayrb2KoICgIe0DsA03sfhuwH9qsuSl2WcO5l7CYz+geGTHWyePapTEP
dPUdp8eveqFmkQId1TzRx3v7+8xp8Xp4laRmlUxkPsem1tLZiRrx6s8dK50FT7Ii
PnW2eNEDtdM3P3TRoAtqfMe5Ucd3NZm726yGIYnGvwbunYl+DrsVwuvd94Gal/TP
kDsH1J029QdBoj4lybuTct1KVgC36uQQZCZdZmgVKCgjiYjAm+AUT2Hb4Y8gDuyh
X1RuttXNixN6GfmJZ+uZtUSGxH5bvB9XSBkU1qN7srfg3E9HfiWs89K7RFMU7uS/
6Jm+qHRRGNavYwOFGbmEpa6hRAW+mYZi0RyT5uJhaqHfK7QVt8whlNdWnK4vCiBn
VZu0Hg2EAcPCgZvvxOVxLFpdtLletFku7RVDi8RW7lIVl7zKcQpSz4Vlv6sziP4d
0X3MhdYCXKJSMAyQLFkwIOlxH/ajRz/BlHZ1lNM44wO0yTGM0kXGX5stBAUQu5FN
k5ZutodNQaUHmV3xsiTHZ2pSIWwWWF1AVd20lUDbeoWBXoFfrW7DjCipidcWQ4Gl
TNzvHh5PzZN38qhi7EXLbE1NxS3eQGanAswLDhP2UV28U5VWB2hGjtTSjF5Y7yiQ
J6FWzcBj/hI+PcwkZLLHFcDS/NRt0e2qZoJFYVA5oUJiA4ZjOkkAONm7Ymc+Ogfn
U2IzP+u0dWHCLEn/f0TaVGZgEHM+sbQwvvMC+/UhC4v+y+37R1pLZu0SZ7L+z/LB
BdXBo8SyX1t6mzVt7lbqbb/0hGtwoEKb72/M1g8QHUjWTCbpp+53xjUYSNF+5y77
EYOjtKQhlLJlikNH91+HXmIuH4u/5DvuUZ8Q2F6M2WpY+ASFZh6qqoayPEmcunQg
fq9Rz80VF9SvjDV3wb0n4xk0DdhzKK+gFNkpsvAK/wPXYCIMICXl6+JGuASZrmAg
+HHq2C+bvbl+Jwk6ZJ70YvhFXCau6eZtuZO9toaZy2EmavFlo57jUgHhGM/xKv1B
RukZ6v2H3S+vZvNdWaE0XAqn7CXymh+T3cUZgxgcHz0LDolIVTNrCjE4tZK8aXLE
tVVQHHZ+hIY1EY/aRd+4uQdblAeaiblP1RYl1V0q11PRXnwqhzSIdllByvBUD32E
Nu8q6zxloCidIz8+VXDz3AEtIH55irpcnTLlhuj44R0HjHvr5L3KFiHQt4yKx+RC
cxDq/Q8gBpU+IkGEHnLOiauA1mVKPEf/bR/seAGuxvseA/uvkivArAJDWKAOK76G
shyRpyV1JoFiw/1I9HgXe/cFdIz3QrAiZbp4TBcY5InyzbC5JjQYFnosbe/fczl+
jAlvY4MYoqqlgXEinHxaXYnsStEnYg3aapfQmw7wPra7K6QinSpZz+4JfSc4UOWS
d+ihm2m+5qa2n7AN+giCTDwLIkSlRKxKtAC/G9HBWGuKm4mFN7+NNwgEiVtYbhQj
JzHVhN4iCFT4ZVJZiItAchF/dK/vwCTuepRKJsQH2eBfEIuiPzvRnQOyhnNdQwY0
TZyZzxyXji3ZUQ+2ykRQjq+J6kw2mkmU6KwgeBPIAxF+csRcdlII2pNpiszyhUn+
/yObZH6tuu8fPj/85QFoPv+QsqP5GR4tG9XMAi5rkoZiIsrhk++KIV0CzEcwAmEG
YHviOhaWmGnzjjsXwp4VC9R3Ug2xahrCb+ecbNEnd3UW8rl8ZCLmHK6MpTEEXepz
MK+y4ttIO3wm+g36ZCSkOQtoWnsfaoR13TFMc0JK1EZT2MD48YIEzQJn2OwPd16x
Q6Q5iR6+jH0iJTTiKe1scg/iVZptkChC1Rea0PmCLCNIMt7kzpYYExjcRIBGv3KH
0oz6uJdemq30WUISzgXewN64xfG+FdfYgfFkBew10kuvbEYETKkZPoyfQ3RuSfek
p3R46UorrAKdFlvFePpYw1FWwdOndZ9Atl8sqWRRZUB9ba1xPH85oMtMF/Gsjy5Q
RhqXBo4yLk5SCblncJxEahqYH41y1mzy7b9hVTie1jmGwQYzFFX+UnUPy34Ft38B
9HUsFoWuBLb1MHpSpXicESvtGLxtmWE0nryi9rOEKyhER9RcMYVlXJqTY3btMWuo
SP4JdAuoUqjdafS6ablE+Lk7TWcPY3fLrfZL1F4h/oIi9qVsfwCm4xgSSuqMr/ex
TUJXzg1qP5LOkRPwUcZWI/6Rqvdm/YmYG4fSsj3dgOuQfU4gWtqX2zYdxYAGeleO
sqUbG/GB2AzBbZU29rSMMjb73C+hfe+MIK8DUYsrY7ZvT/xWBAmloq6K6PhTLz83
iyYW12E7HY21wzgsC4ct3iwlpYEqOCOA/GPOu9LO6yYkWcRRxNrMOjAQ2TJKkH83
Ybat1BiSG4779D+6tAXJU3zVe43icCqzq5lmX051w8YfEVmxxgFQCcbuM7EaEzKH
gtre/rj7EWWaijiAsacgdi+Rc54UIaKolSHM099GQNnR8RqsYHbPWhhnm0KkT/EZ
GF5hKoQqd8x/AoGyQUOVbrPz6SFZeqtQxDVCG6mEy+brgXYNV05hWwDJ8SraW/YM
v+YyzC+UO8DL9VRWUdo2lrdi2HQXcma/eLuy0fhXydyz/Wi3X7KD8J5JnZH064Hl
2RE0DG5s4RqWyyDJbcj8mQidik10LJBfKtZhq0X8kklWmY4iRQZ+6Ahe37KtP4nO
LNN8U1ormYdTYnbp6U4Y0UXsTyxtm3Uby0cZEtfQ4aR5+wQ3fpryIbwURgk2q3qt
rczRohByCOoIPRCrO1j51zOCV6qNhb+u0KkxhXCIbPnzN7e/vIlQjVcWh1iCWS4s
2CuLG2KX3/qC73x5ZRM2TVONsG+1ajr4HPWW9NL+4R9YCyvSZC0m8sIIXZwwbq3s
vnXRw+V+U1my9pnhKrw9FnCPhYcjuQGBisUtJsc5PXizQIVkjjkfBlXnEB3NPe9A
dQUye8fZ0p04jXO6LsBOgFi0P1W1MKaq1NCipXIqTOo9s/qLK7pzxvuEqHR4PyW7
b8Tz33RMX+6YTYi2ZnL4/orFtS7qxM5UgnRCIVswt9DAYsAT5S/7u+LSjlLjmF1W
jXbbhCNDtbX/D+rtQ8DuqKCnZcYRkcWkzDo4EV7V5Wpo+zGrK/g1suVCVavexxwM
pvIKW93rDDTIuSZzOqh722H7hhZx7bPgQXW9ei8jFuzuiMVnIF9QpY6kwM7eXPz8
qJb4Vf4whwpR54WgXP9p/Zzf9w1McUwkjQtaoSCir9Ar1EAN157qW9NB59Qbl1p9
YtnkxufaJJRJSxxoIo5+aUSkwKbEqpOrK01pk4R6FKSCqOmn7cjAy5cO5GwXyb/n
xM1ZrLcn6GqNJ40iFV+BP3FPUdNvmBC4SHFGVVS7r7LPanBN/g9qgyNVgxbbNRok
50Bn7JOyJgqXOUbK2cCJx21S+gQ+PRcZt1yGjRzcL01LCAmzZa9ctx635IbNwXmQ
ABDZW+gop2/0aTCC/B/LIeL74hgeHnJtn2rTV5Myh7S21BryGHgR5XxoyEEyJZOw
fKrO7zCnus69hMWSXngTv9COSbw+3SmY1VEcA7jjfdRLcHMacnZwCihAxFU6eYJ6
kTlJntVab/p7h7YEuI/KAoUrwgGso/LRjDA9WsRRmkZNBRGX6gIvFPnZFb91VrgW
K+ESFoIdjOR7WkdQn5iwg9ecSyHklUBXnFv3U/0cpIGbi8qJeYhuFiWJFIMsVcaU
ZAZqDv0ONqFcm64IuMQhctGXcD1HvXBjlvfJIbIUZtVvBM2ystJyIBjlTw8sRXKC
43cm3MlFoihrSc7dU7uzLY7/02oTOWiOpdB8VRrj1Ez/eU6zt80hxf9qnBCqDb3O
vUPaLSdmU9zLm2H2JHDhuG4J01JqUyjPIx6P0JvTRdC4eLh87cYNnX1T01tZfbJx
Id7SHjBg8mUbH9hH4f/gD5HTTjbMGnzWMefm78pjMf+6th6Xf/b54mG6fPwFoTwS
oMIykPPflVwtvZffdF6ixNWYle8BeeeVX020azMyS/4bc08N0m8kCSDVrRT6dQl0
QY913nBFJTezT8HdMx3jN5n1H7FEk1fvfv18sa6iEQDd3Fwllq1JiSSPcYS7oQYh
t0Mq5eUjTnEqPsCrHRGIgRj0fwqiCRusqWbMKON7mureRcaRvr/6ySSYm7XnsfC3
eF5quG4vKqpp41qEYiR6MXHGiDnmggxkeS+VeD2XrZ6Afp+l2IMv86dHFsDSuEuz
QKmTUify9zCSIz1t27JDPUpiL0RUeTcxXBkShNql9SZ9jfVz+f+uKuw/ryL8FrDS
rvfZ94e58lIPpkpGWAP8/sV2Jw/mONmKOSS8kEP+TCjx7Wk90uCm4YpBHNDRbXHK
QKv7QSR/TBQHDciHnDrnCi/qnxfqKTFyQ9/LXGsWcHaZxONr1iZOsG7YcXFe5Dwi
IeRtfLMD1R3uYY+kI0stLHVdNOIu2jZGmF+6tVA6lgF0STpvYShbUHa6SdzjT6Dm
/B7btbWhXGYEjBr0RJB5NfBqbGghAtzQUB5PybQVEyndcdDdThfv1OAXUU8syLVU
WIFhlYcrC/2q+knZWvEVRjY04XbReaEpar9mbn0TsLiq5imjwNWgzXizhh+wwGxg
FqJfGC+vof1XbRkDschUnmFBZE3DfF1rjmYZ1Khc6EP1kFzyUcknr83dcRR9e+7T
z4aoc5t36+XNp0xL9fUeFKaGdpzvm1xKA/WFaD2UBpcf0iV0ZOELj32k2sEm5uQm
lNb2KV0V0gs8YMGTq7mnVDADFGhkbEAfXUaKNAq2QuUX7kpmwt3knpINrRXHKrOF
/KKQU0zmL2QtPnEPGrouPJpjbPwKJHuqFmK7KtcAKEWfC+5jpo4ll4RU+E9Z0rvB
OaH5Dp2ISXL138NC5SCT7Cq2reysyJXMFm0IBo1TOFWFRlwh0GEuw+09br8MlKDZ
j+xZpmcPduAf5MDGW7qiOIsqK4eDICxH2Mrk9IwQ4XyyxfDt/6fY9HslTD0vvgf0
sPRS6JkpstXYQuGVYBiZWVRuGf6n+27MRvQbO2dvUQgOcwzbDKyU0idczDg1mbi0
LOWd5n2NdJHKXeLaBeA3drZhLVqcxlqnh8osL9yuqHFWj0Oxcom844CM+Je4Xexa
HPLBMn6vrKtk0q+Lo0RxBPXcAxVaiK4pgs57LWlLb3Oeae8jhiRneuWBz+AOZCjc
qyumAdHEQ9OcV4RH49sgSs6wdrJFbau2csIedXLW+ZZ9YZGV1Bdw+ThS291pOLD9
iSUS29E5Btx4eyW7SHmyZN35gAfmqjL6DhF3xyDBsoEG70nqGqn2ERGz7SFpQEaL
FX2LqZ8+4iFQpp/1tfdfrbYusdbTgcZO5B9XsUbUv1hsLnW8K330NgN8zEm46Xlk
ZAOtx+TNeS8pczN59Qa4puXClvA7Yux5sdaptgHqiGKY49eRENDcQ/J+H/oFfJ7J
2hQ6DXZ+x2kIpJRYTpfMXCx7x7gLZEdztFQaERtV2EWDpORSnibPZvKl5hMU1Z91
roztAHRA0ZQihB+JhDLmco/OxiFxgx3+rPeYWFy/roUxJA/ZiYkVef38uSoMPj8s
lQyLO3ix2i/B7G5NmGvWvXhR69yE6gAdCdDQxhG2FCpRjP1FreEwUTlwboCdAf2p
SMNm0iK93UABv2icfnH8ctXtZIZoEd8RFoGY33NvRGv1Om610miP4vKXBYmDXvsN
PPitYUtjbfi3g0dvsfOEY8qGO/+4xEQdmc6Pd8M/QcspN2yIKY1MNF1sqylrrfm0
hRZ+Py2jQozFTZ65CB/11URNdlcC2FNASlK1RYI9S5GhQnfdsDVoswA90lj77ctA
2PxlpRHJGji3KLQWVp322x1z/dvr69RkNeqlDn7BzFU1rNTJbZDmBP7BV6rdV5NX
UNXXPVfI9DAmjntN4N3kEvI1zR6m8ELvgEmQZ02MIwBOPUVvaaGxM8nX5oHzgKoA
zvnhd0l/2CSkQnMMZFjoYovFFwaiLoTSwBFJOK/mx1/218XjhUs8p2dnM1mQYzdI
1NKdvFNzG+pReO4+8hwmVT6CI2DxJ5zjDq84MzoQftJmdsA07uuzxVhi6HiCMwjx
VgT8VTMaXHBFbxsPupTrAAnTtk3dcFFodyYmweJMjgOBrleUmKHyi3gqzVdamChF
sO8hkEgoEfyXE7Z9hOH1S/Dc80yrbeeHYCi53WFrwS5blepXtrh8H5ZqCNDvtie3
yjxe2GbQ44uU+OhwP4vqjolEXBqBxrM3sbVnYlaSIpcHOh8BxxnJbMam0zXa1RUR
yytgscsxiHK68DYes6VJ7HJcc3n2qRhRXjS0Lg9+ApoYq3+HaK76zU4rBL/w8dlE
fsFeX8RW/61PIwAfLF8zAW8Uc9lDhwcKUbWhI+nTGrsdQlXc2RbwIs7A2lFB9S9Y
YQ9EqeQDWMBgu4WfuHRO1Rb/qqTyf0xWA0BuVXwDrA4CUzM09vBsJ1OOGLrZoojN
VosrOPhOiZM4rg5J/CGSAv8B5T03lK/Q1PMPzglrx6LZmMKZIoSmzx+KI4rinvin
VILeKFmuQa/28EtD778oaH3FGVDe77Xpy9FDdMkLCHEGZEFnvTeddo5WQP7r25SH
DS542pLKHhNNlFFcrYkFloBS84/uNjaztjSyBT8KB+8NaclNBkI8wL5a1gHM0d8H
bham1cAokbAr/iboqJ0oTJM9I9Q6E3/zi5MNIkCl+GZRrldsNeQP+fT/AQEuhCu9
Sg/cBcr4G5UDJB3TUbA8GI7FJK9FL5o7b3MpnehVEv+0Vi8nG4oLk+4rsKid/79h
vhAUsoOaKbJ9SVolo5UnR6Ks+lBTH85/1Ex+fZFdxA0jOp3zARjhPB/Ov7uD+W08
+3v4zUDk40gB8mHxobgLHC/OAFVlYXyoPFI7VyUwDbrHTAcW64UrAMgFWEc5GbgP
5SNcuTQ+/u4Tr5kOTfM9cRe1PoDuzkeOJRfEsqUGJcm+HSLKD8nMn9BAFzfETfC+
YwL2nSXCNRAlQ2qo+mwTcI2e8B2Jl0SRDQU0Ls68KE2ib0wyioLcJLsClfk1FVf9
Sx9vXxOyxPvP1y/pMjr1qDGxolfLVWd+qLacaGAAKzWVyehk40X7tOmWGk7JTIsA
74KgfcKmDDRg6ofuW7T7iRJBFYWTTKxDt24n4DFcb9e8L9FkgrXp3E4dda/KRJBn
OhLDgpb6cSdOp1wqQbWEW7LrrizNGCatUUVgVrqXjLm5uZgLH4YN8tgNCA/PNBBc
AwdN5eRYpzxmgrQeiz8n+UjhbdqGpRoSXdtM0Z/mknFj/1kIpyAdC8jc1lzXMnb2
Zygf/KRFGf1jGczR3AdnPgoEqlSEses2rEgn2IVAytmcGOZtu883khpXXVdQoTVi
8ByVhdSmSEw2iv9RbavTjDRkkW8GkANrR137nebt8HhOw+Gn9yyYt0pM+Y5czrRS
uFtPFT8X5SHZ9oHAWQtH/jQdYmWsRVNEMB1u+biXbtfYoSAnavKAkY/+96ICnvWY
jOJsG9Ah9Z7Ob0KeirTjZ5ZbzaLlQ2n6/2I5kRQuiAPE6a+jpyePKqqVCw90qWwq
gCtHMktvbR359TfxxSjlOdLhkcoVJzvD+OhSGr6maFB76lo1Sl9Bd1HmXDmG4+LH
7LArN/QN26z5WBkDUcKhyZD/sT7IDKjMTqGwVTmrdbcRe2IeAz3w83IWv7o+rFO+
HdMpbK4tb/hg86twD3K0vjX0KkGSZF2cMax/hcR9K/yFZTaxBRxc/s8KEb8KvW1r
MUKWpk9M7asj9CHIiyfA1Uqio/6paLRS00YffVBL7Q3XUxEje+lZRlVfElepsghw
LpT2Wy6dCiOLQ8kONZPM6NqkMtnHzXD2otMPg4fT4ACxQ+QPKrx7nk1ao8wgnWB6
lfQ8jE1d8PXouvucVoYFkMNwYCfMLLc+S0u3/TvQ0NKAJi0O+rXhWSl6A81e3QcC
adZdLPIRiFhRFV9ZrpC8rkk7JaYT2EX5XKd/48g/EB2R/4kK5Al2p93D3JClGnEQ
bG5cOTXAe1C9olGv1unSihFQzLcLsAKLDs8GKinS9MfGsJk00Zt0tDnSPlhL1RKZ
rYqWiRhhP1Xv4wEPfuf0VprTCdBXsnyITVl5bjkU1dpDH63axjvIsQPE+723QfZd
rb7xezGgvJeD8ZQeWctwFFrhpUICipUbBRnCOKxVK1mTZhCBemyArqIF8PlCSSCG
e+FuPoqF9FGY87jydMUB6djG/yZ8pKDXybplFNRccZehyCFVYir00fOyFLwQJd/V
G47eGxc+dpFJ7YcpFZZmF8iDXk4coEEmucXngcbcvTbDEPMPnp6bDUEeVZvUUNVR
HsxRO2COfeoFLN6EvjLx1lORo6toVS9QT1vAJsau/rwBkk0hZBSKihJ82r1PLCdg
CJTO8pVBcbZGGYEzygy6fXj65cXMlinRF1DeSpGLS5N4J+FHZWFvdnjZ29/6ctdf
S7roReu6yAW9TiiUgI4mQKRPfQZ/BYipWY6biHfJnZ81a9t7qeNcUdUwbNmWjJ7s
+m147tM1On3xFsueQJtSAuck/isT/51+603VuBOuKq8Fd5owv0EZcHzsVGIPvIxu
c19ZYHJFSGDhj+zTslT/oFNiii08q4FcEq7SHRVXbHQ5cDT69vNFbXVDJZlztqqh
23WqrKMvVYzym5StT+UaWXVIx9x8e/LfbSbdfGljvwTl9UAcRcTWMb0lGusHl56m
w+jGGEOt0qaQkQTySuk0tn4kBntYqJXBz75awKI/fZpnh2ZAeV+SV09hT6H7B1yu
K2UxIJstC4zoVWW0v54xyttb4fPKfeB21TeHw0QS1SdbFWgvWXMJX9UF9wmk3Yb9
eGKCPNcSflOESCUVEAP/DAybWK0ZMj4iOIvE/ZOsO0OT4icEUxdkz0bKXcAPpd0L
6pw3mcNwwInBwNbXZunAatWuZrNXHZer820wbT8NVYzcRGF9kU4OWius/72IdZkK
bOrXJ8MDCNRGXqN7qBuprBnkL9KZrlqKDAqppj18D/4qJyFJX3UwlYb3nww6eivf
BCT2Cq+Z3odQZdtL2rN9S37KOEf4n3+aS2D1Mxr0X+VZHTU3MsxK/zmBZj4aXc3j
IkH2IDut/s5MBWRf8xUUMD01mLbQFkmadCjEACLpEHKbi+FNMAfbvegnUhm3uUW7
KcKWsBQpGrx86URKP+DOCoAA52eDp9QlmPw8XN0rlCdd0ej94GN/kbb9V2lug/BN
Gs3ej+sa/Gkl9C4VjJNcw5rfmCt+vM8ZWi7DG3RyiTQTBr4BD5P2QePRvnihJqFY
FQ1pIcM6y7h5i3dsNz8i0kx30iHsAXs8+QMwKhtbuf37x8uNrbfQgJmUr0QDZz4H
iMQo3ULKBK9LMtPnehyaTnRSZugGr61rvMB2Yk5kqZieXAg0N4uc6COuhVDbkISN
TcQDPoCenZ3LDygMMuaHgWclg9joeOMcNqUVAW6FH/bQpq3x+xLNuzy1nIurwW59
dTNR0MDITgIMSy4Ia7+403qr7ARFWb/g2J4iJOAauIonXFf6iiQydgFsgrtXdqnQ
qv1hPCLEnZc84TWwOMxhO5YYgL4KN1OFyLc6eECp9AnjyOtUuWAM3m188rmvW7tx
FVvbFqeeNCxSiHqVnvuUEv2pUYtyJa9XSr8GyGi02IfgOfDwldnc7XoPaNcWc3OY
z9U1ANCMhkI0qVN4hqU2r7IKOnKdWvhxUDBzcQ97/5dEA1hCWWzI/MAkt1AALpV3
eRFz0GlC2AEQLySPcUQxsjQfBOfkWBqdE8A/4zh226EtzPO6zxODY/Qq8/Fbn+qn
jiTrMQt2vJOUfg5z/TEn9lg6o6aXNfqPPYkPJaoWcgdBtmNYN6lFNpKYLGrQ5J2z
Gzt8b5pnRonj14SjelMspoxA2pY5iKaW4ePjtf6XH2oQRYElAFXUYFeUxXiQEEAD
+yqILwR0hjU3cTNVbaBtMmYzqt895J8EInNjN+VVrKKQBYqi/yhcmZMxPittSIqM
EPfVMoFChIGEyPBxReNgBtLTxpXtQpew5bOpwYPPivhvOY7WhCDNnCflEPCTawfy
r7ikG1xTaz0sRcmvik7yhKNYPKvn68hRideoI+PH1YJVTvjg0pEFrkdlbbzKXLKB
2QY0my/KRhge69WZZPtc51uAEn2PDdn1J8F1Xk2zquAlmK3nKJuDRuDJeZdmbr8M
PobXPsCOgPqK3FloBMDeei2DtuZuAN+Frqg0nkJztirJ4YH+vPdVKY3zgtHPtwwq
6J0ByH66fYsTT7cgvPl4OAP3ftXXM6l/tamEP7LT5jwcaPZEmJk5uaYDQ0TVWwbL
OuRBrsatCn8Bx02TN2CPILaJZISARQty8ENN6JXID36ir3/lXEQqvmArkVxBAhhE
EuXE7e63SXdWWDbb4HbOOpNU+3r5EAP5KHjVyo94NZtMPnYgT0qDMlfNSX83p1BN
dTHA+zy3iveuTjP2qTCl+w8ieeogqfO3ppRCCzXTdmZkkwMz3Ewgqtid3Dbjo93V
Y8EKRSNqhhE4kv4j+imfJDTD8JT21C/9PhYEbut6rgXzLaBge82pgBi4K21F3T8I
6SXHv8EYs5Ahiwm6cdWyMuTwFT0QwTDXgGXn1vcFSN8ul7QXaHEXc4dsGN5vKNkn
yM5d8qFmbCLYtxdOIILt2IKbf3sQ9r4mzfd/KnpT4r4dHKpGq0D6EDgYRP9GoL1L
TEnmADIauHnvdDGVP7KV/Lu/Ruj6h2+jx/aR/hdgLYmh2U4uS0NmKp0LEhu4dCAg
PtbqhLgl/82PTDxj2myK8jfY08sTSHjSZqnQvfS0MRGKNRxhrWKI7tNoJiXOxRSo
NY4ZhBKa2zDEftRImO6LVfPvd9+fi3BPEJ9kgdRjzEu9ivaBUkdC4+TAz2f4951M
MQLuyopAoeuqaRXRbR+ZxWsNkywfo3v3fUI/X4/O57zf/e3dyjQ3qsJq3neaQBUH
3mCBVby76KeNTinBnBATZ9w49vewPHb2LyAN3XNOLtxkZnFbTdVDG0pajD795RsX
U9X/kVdp1kTTX61vV8UMPFYU4AdVLEVnsso1f90Ptoqsh/WNn73D31u1Mb3LOHzy
Eqa662eO60RyWNOL09Muf1lpelRb1XgEZbMKFS667k46b7/j/zGoAVCjGe8d8LN2
pB354soPFUmjIEtER32UzXb7JSqYbu6+YZ/gOyzqTi9iy9sGGHF8j66txiZdT9wd
9QjmHzPk/V8uVuVzMjbPEZaB3Pq8PSv0/5NYh725+VlXt9AObDTT4Gyc5X88xbch
mHWASNHuwcJ2EFbMvH7ko9yWE7r235bniYchZiUOOdQRdZgk1NEWYs+ySLbofayl
k/iDuhKRPDXax/Qrh+enXGeowBAvIk71k7qObn3o6FE+DKJD4opk0jH4Hm+Z3Lah
ZhwkK74UklbOS1wKBrIsd+9cAiQLu9hk2nCZcrQU4cYHIWI2VCcGcLcS8BiHvc+G
YiYgbhpKXFLnwbgWGoiubc7U0ipX7T4joT2CnSHZo8SjpXNMtReunVLKd2bdnosT
GMbmI91o7BlhntqoBb8KER/N9Esj+ZY/o/0Wx3D9UfdXYRKBQssONXfSO6YiyV4t
z5XSgGPN/3lCErv3AfQd15oSbcNcZ7MCGtqM36NZF9va3KyfyaHW7Fb39xwNlz/N
frchkiPxJTeCEX8uyh5fm7ZLCxCot6sw2dLTD7wknaFRaFoDT4iZfN5bLOh2FKTh
X+Es1rB7Ouq1XzJvS1W1TeeFmIWrkif/ltThqNT1hp4HdiM2jSfuuB8WOXYulP+x
VHqmCWW2wc8vQbuJru/oZqE1jUFKhT2fAFb1b6TWtnUmZFWaY+zYcucT3/adjzEr
dmHy8Ia6ZJKL8JjOFZDTxS/7YesYeHxru1NUccr+Wo0dE1JHdkqIMAUHPi7Q9ODm
w28JNo7i52rcM7Z+W1jOpmd0MiKtlCGOGDIOJdEwoAwNIbIrfvNBkKLBsyZK66wO
/B+X+cFTwPoSyXthmqKZtnNXqS5mivERpdCNcT7dpfVYaXUg75CeUZTA802xUB5E
lAmlPfE/CBrdl7iT23sei/KjFEOckIxThdVCgsknLYU5ANmfmVv9prLBe00Ofy7H
BIx3OS6Wyff1v9zT58G5Hc0yErPuAS5kuy5pOGz732LUzaJh+Cz4xOTn9jxSyyRD
pGCc96Aicv5KWUj2Tg9WlWirXMaKv2NS5gB3KhOJM6nrA4YbH80dFYJbayFSEnmJ
rG45dv6iiiCNYkiTV0nvaWumpYs3qAiCkIVlV2ENedwGFzkyCpv8tH8/UaZ/EEC0
g0SKGJTeUh2+PDmwjSA9eGqkiOju+49D15pxpCkllRT5eKZ/Mh2umhB45IiEFi3p
q6FasaVOaL/v8G0ngsSezdD7oVOCpQii7K3hbnPWLmoBTYGKWuCUXijhoV66Dc+4
HNo7YUb2jc9Psk3xIYLVkCDvMliFTphjRodGJktpVUaI2VgtkfCwaXFN6Bvx5EhQ
ibzYoWmbMv0rcHm8qx9kp3MBvFn1klJtrWdpQm0nidQCyHiSefOAwREQlNxqSG88
Rwwh0Mb7QwppFWG9ooe+QLUqPMkhqBH+/JeFX0Z/0O5Uc8oWXbAFHF/5Bkwt81d/
F6gZAWgdueuZur7BHv7F3q0dvFCUG498KLslQbYrpsHM79Zp6ZKNJmA7jma5/3KJ
5KAR5jtekFnQHcIzMCzOr1b0Wnq26c30GbQqsQOMyC4fR46yoMebo9gHNMb7Gvbs
tS5MzJskH3H9L2F8tbFQLGixe7qpKeXO4dlGon/Uc1fXD4t6GyD0lr2ZKw8/bZpI
qX1xBa3kDuWy5fTyeyBLFeGz+Av+RpBb0RIflU+vpl7qTFoYAScA3VWfR5zABDyt
4cOM/2EL+DcLNuxLQCy1R8p3IK5jcmSnWF9bKYLCnrcMWyoG65vhVB52dQ/j8/sV
I37UzLOVfcjUFhTdtb2F9Vo7bu3Digozx3qx8bjNV868CpvnzFTt48QzcB7YVxy5
XScWJ6M29SjXUS6uG1aMRj04xZ1QnNDN3ShOr3UP55ahhia2ge9OqOj1fp5EodMV
MBcMEvZ+Tr7+jgb66mzyh9Ld87NYNRC5Ml91Vku19rx8JxXCjqt2WWx5vpv877Qg
W3pmri0dBx0/3CDhPyFZRcK2CbK/eAbOhtXqdlMhM+Xdo/L3FMhAEsE/HIwQlTuM
8iFMTEAZHcMtGqLid/7JWOzt9KgBHfvRsAcNYoiVbFSxJHQIr1KGNRdpbaPB5A5z
k26S8UWT5L3dUeqI+yGkw7uW8a3QpSdExokF/Hm/pwsTpVBzwRCGzrcg64NL/Mno
5HxkwaYkUZIzh2QohPuwNdDNZ3r6imlfoPL1cBhZpNdEvB9ZmjTvquZne8NiA2HG
WaQP0U4DdhTkBhiy73Lvzy5r9vynT38QUU/z864xjfHbdg/GKBoW1rMh6eYV/J51
Wbwp1NiP/7SZnScLVlyltwUwDP5IZqGIjnTmJuZmA0/nnKwBt67/xNn+4fHoaphL
i6/Mw3KGzt+TCy8wc/4GPSUoK5zWpXjPYCs3reuT7GxFn/p2QWjvmXHF4J/eZ1Fy
SRrTtkwi9I9pir6M3FsVwxQ6BoDgRveYi9jY+28Lfs+0JPW6m1+1p0o9YY2+fjly
LzRpYY87jP9R47wP7k7WW4Adr7TUYdvXuQJuf/W7o50XgVnIiFGoNJTmIktxx2R/
QIMcCcwj0E0wr5fONuEDwIiDo55wZjrctzTAMi1fZNKBntz+HncC041L75OAsLk4
aLOrrswiDUkUjYsF2a8qidg1GYt3REpoSyNY2RKyA1ts3qIkz1Z82LPX7JdKDEDT
MzVNyGtq0G086ViNB1Xf2KuF8lImdrOVFwWogjyg93PFSzU4Ei2v31JN2Mkzt8kJ
lYsLtE6Ux8hOkzzlkM+EUFJvrjUnuZumGzXCHODOfW4BUeeCrpn50HrR1WubsHMb
MgpHfS4YPap3wKSZh1D6iZwwaNv/lMFS0M6HDFOiYAHNIVCvS+mf+eV/pB8WIA+g
XRXbhb8QXUbTLpkHYx2ucf3I8BGNXm7efqADwiHm3b5e8ZUq7RUFnlhjYAYcqdCx
YgFAiR2V2rNZQmPPqRWjK87n+2UHZg7lKTWUDXNY4IjQMTW4wTXhJ1sCJyGI2CNj
ICA+sH6FnT/By9jMpsa7ev/CEhYDUyUTADoYqw6yMpdWLV0icdGkZS4dYB1SGrbx
Rpu+MVoF7tuzUhZNjOyXW53Jk3EncIoGFGPmVTL1Tnsgxl6Dwb5Jqybfp2PL+Nw8
wGqRTykPKjtkrAWDwQKCYc7oaaonpYyc8KBsaU4ymHWushl2WQPR4eIffGebYTaa
XlZ98GO/5VjT6IqMAP55bW21YyuPwNWtNjx7OHclF3AsL8vp5cMgpr/YwdgxnmNd
5zcONpT/eb3Q1unJaIiIh9SyL5BGQ7yIg9QTvCF0ylGqony1mdQZ3e0UgE2fIGUs
i6hW2+xATRmlGLc4oRUHPxpiD7bGAg5VLVRyA1mZJF9Fkki6iNGV8qMOEXoHv9RY
JIZXGhZpoL7bQ+IsgjuI9nyGdvj9e1DDjzrL5wLi2+2lbYIZz6ytJVoiF1z5KH8P
zhN0G1uE445/em5RJB/dklisvWNu4+LGjU7G/Y2W/N062SXT8w7WtK+VeIurbecR
ycG0KE1VktoqErKjWbNmyrqF1S/dzLjsbQgz2y6jepfnX3xZnfbUD/e2DvaWhBL+
HAlPEzXjwcvgAB1A3AQ6eZJi+7P4A9LGBa3Xs1slwy2OZ214NpUYR6H5VpFeIG1L
HHL47D8rhuiLkLLLL/ZyTM9BfzWYj7zFTFaH8BnkN/A2voetwbkV2HtcGgfrMlJr
IMM1dvI+hCdHe3a36+3O8khK3nq5KKYizdkMcpv7TZivqBoincUDV0QMSaFychA/
VbDMhDOaWyjPRdFKnjSTnuhi0ZRRH/wgPQYH4vbNhPWjbSp10GcPBRb9ERqYBZTA
aq6J1igTjPYx3dVs9MvqUKF56d4SXnDN3kJ1Vw3Ezp3MkAykMuKANcxjM1tBB0RX
dENTQOeib8NW8iEjmHxfa+mk27T+7SY/+Df9J4rLE/xbObOXBYNaP2uZovCzBm5X
8kVoSTgcNoVdorBEKKZB2UGScTUXF17/9nq14oM3TrcplQ0x/xER7BXYVkYpPYXd
spf5yFZSVye/Kp+ENCtco/DcqVvplGCS6VBihLQQjWN8LhONB231GDVF5/Q55d/l
XLjQZzxsAtmblIBZOUtpS4+SXLoQA3cgC8ib9FWFZ2kdmaHb625j4REIsZ+g19yO
xUOLYBSbc6fT68r0nloB9+S4r+zPGQ+yK1Pg0FzaCXYiDNEVR7immfNPBHD/zx+a
hcckSmWsmzwBfRYlInhxatZxfTHBPlXZ8VrFJDVEFaPJBRGJwqFRoHZUmkeeFT+w
Hae96J8XQnoQX8YXwb97dQhy7SMkJmD61trJuGTnzEtz47yFE4jSV/4qkY6hzID2
H3nG+nWvFgUu0JLHCvpKE0gylZ8JqKJvHeD+gEK7cpo5UkezJxOJheQRKZclPqFt
F/e1HHMRqfgwoUIaVtFAB54aea0T63qpInDNiM2i91504zjObdHfaVuesD8hKUN9
2qv2aQWWFyJjQMOINF3LIMmmOJWlMUhpddc98G1VSMb/qn1Kw3dalwc1ounj777t
ijBx9ejOz0JJK4Zz9+MwCH9dfl4UnsYDxeZIgobyl5xr37VirfTpFkJEU6prUNhN
nZI8zX+fWqbLYEGK4hKtWfCFIRA+ysXN07+TQFhG6NOLu5gKXCD2i05fXHZMxWV6
rBoJu9+UfdPtTl6S/ZaQZ7qN0/fswmoOqXd24yQaXo30qeiUphoqlO44OSn052CU
8vYJNNHZwhNfMXUte73f3/l8dgK/e30D1JIr8+978k2xTFNbiJEYSprZL7B3ophm
wqaJBVehZ55wSl98XpDL7Y7Vmo4ODxTaTQCgi9nEnRser+/fROSiCC4Rq5jFk/D2
rndBy9lHK/nWWxKzd7IhNp+IDkRI9yTDmxo/xN02++eA/pHsTXXxTgJ+QTTiNEAu
qBLokFpiEbi13O7ECPK4om+hN/14qAwlJgGXesAeHH/dRPp+G/N3sA+8rwyRwfmD
2+dkGcNUjYAtuMKG69U7FiNdVTKF4CrlgC/m6wOhAmHc5oU3VqCSEskF70FrmXo5
k4UTDdFgt7Oql6uwRGHJdL1TTRIRxSUo7EvAN87CSggjKwVR7lo27on7xZJ5Dst/
IZtKKzTnToOYJ2SzF7vso6hbNz6q4j9XqaZsIf6SIxLLh+KkeAcRHMtJbyVHrfBr
1JdNf95N1L7Sew108UC+XFLdm2SXEZU65WzzhByLX+ZGtm5I7wjhdkzJAODCLi2R
DjI0OUw30bAta2giGJbIhztY3gmRKo1g3q/gpfQmTcRXSU63/rjEE+NtT3yhrV3x
ZwWCeDC8bbF61goIFa+uzwaLYB7D/HIzUA5WWlkGZQ4XN9UH6xNLYDK0QqCcZKmn
uJyOVMO45ejZv8s2vQWFq+qbxeoPuwM31Hbn1Yb76arf2PEsPOdZmRpO9xx+QBea
4w2WJ4x9TgQ8jkD3yskubAXh4n3BS9ODn6ecxVWYpQKwl9ms/KTmd6S+208curxw
ocJxOUiWEAE+FM7Y2wZ3nm/pXdhSJ/c5NSP/wZl9e0+dfNbNN3jzi/Ombk7TveqZ
dWIaK7aEDJu0y7KVzPF929cLPkvhvSZX1ucDOXyXsTBc9QnhkInqUifYAJjPoJa/
vQLkixkSU0fgEANeOzO/td+g2fYTL/QG3GkmUHNHtRS+WXDnC8AoRn051lXJBQrz
o6G7gB1w7LvjraNa41EOOdDGYEwCsQ/fh/T0Lmxn6wHE/eBIi0i5ndVUWdHDFaVk
hMtMohBBOvm2Zg49E/ypJ7WP9SXtdrQeqL6yIy/yyF/N4gAZeuXYE1eXKUzap4Rl
5PzNuWD5I1pos+/BelB1r6hOZOtaCG7H/pmsGD7zvNMMEWGBwn7PrsPHZLoftIdS
1eKKkXi6r29pbfz7g2sRIEA9Qs9OZiMq/4Q3GpK5rdt22kdShIaHDnqJRRU8xASN
wQp0COBPdDkvbkdudYCX7SMyKmbb70xy38eDq8yJ9x3dfkscTk5iuxvHcw83j6O+
NzR49yG4EZtOjE1haljziaY44zEdNgLCwHfjRjdBgibRP+bQABDsstFBLyHQYjo5
60YhqUbi+58bZuOm7BFpRsbwyqKAqpR31m/Y5P23zNBpul9dDxN1hilCsGPJnGoo
DneiZ3c56sM7RqByrBlb1bVH8TlX2BH+g+MPw7ihQi+WHNl2EpvO4Eextu8bVHzg
TIXWXjeYvsGPWwypXILjXT50C4IfMBGyV5+FuK5JQWYPRJIXYD4wGgr3AAd/CVjc
xL5IUJLjkv7B1ROjO2REnsjpGDe3qodAmcHmhECENvCI++JIkLIFo0Io3EtJkSzn
31adSSJJzoBFG8AwjusM9Tuga1Ya8/tbRwlgEhYZJ/F9nBRLIECDfevsPxxTNHAd
OwTXPQ0lm5tsP1sWvvUpPElx1DZFne9s9S3M/vGyLSh13dztJ3NAGVzwudRdkrdG
zGzftaK5yC0ZO6Qx6UhNRouqyNibmQToGF+WtaANQZFFpNEZSDpUlucCAWWO7MtO
8tfNkjtSZFszjvZtNP8e+KtGPylVlhDg1ZLqvkPrqNitqH1xqhpMtkf11HBHyW8w
59eo1U2sO67QY8onCcLLeH5759GeKVnmSZXQJBw+JoJAHigsaRgQ9TAOweGhwh4g
NJnyPCsN2Wg9U+Bqnp3DPTzxhZ6lA31F2raEpf2VCJBD+GqCTBJ9+PORI4XBv2SR
4pytRpM36/MIY0wvzwxWik+TduQYBd7DgeuEQFW8mK8oy2WEmtTQpZcgf39MaG0p
KSuRn3IEwCUNxCLjjePHC2vRjsH9r7C8zMn2zlzlhnn0o/FSmcS0raJF2VNTsLVm
tqqUsAEIxDtg+CVW0q+7pCxY3ZrwqAH5gyii3qWik6ixR2biYA0Q+tbeqJdbseXL
jEyLdR9zwEXSsX5/xTF663G/YTXB7ufGauqULSM6iy7H3psY/v8z4FOjwDpj/Y3Z
8CXDZauEm7PK7I6V6vsnGdoMsaW1BXGn8i84SoQFVpteJ4oxdI/O0HbnjXdyZ1gd
Umq/clURjPfPlIrkKr56F++bD73YPwOnlPxErwjLRJjIUq2ZmfcqvzKbw3EvrMVd
i4TPqZuOcriuT8GCdl63B/abn762VQnVbPVauKeOAeLaNcmXsZwcC8JFWTukVOtm
/kxvPC4ckSwrwtvvRJR0Qk8JqWQl6E7+J5LKFz9UHBaWyREkhhuNkdHN8FHwV7op
K41ZcCCBZUBA5kqBQ/yzX9tQIBqnVvmxp6G+ag68cgw6pP0tlnRc+qS8VBskThzF
2TOzuSqNMF3MKYh8kUZtbnWc7Q275Qk9u7OUZ1p/CvuxKPf5TGinqKrNmqPpYkm/
AjYt07LCxbNx87mcOguRr9XcwndRMykKTK3tVpa0iwuXrbpgJi/YWS1J8/PkFOxw
5f6aC9SsFEXLxVO0kG5C1SfCUd/I0ivRoyLBn3eYVE9J/mKXXaWt7CWb2Vv0Xs8x
bfWoPNOX8DwicoOPZWatJhm1umUMyv/tdQl7NpOe8ECIFIGjZ8KrhxVw49UtAQMY
Vdf3kIbmLV/BXKF2Pfjk1WulomIRVbQORGoewrwCKF+HEcP16xAZ+1Il96G564tC
l5Sx+CjuLdKCU0gFDzNRCvyFbzXhgTMZiXykv/vrauRCrlZ0Qu4XPw1jtRWrc7ay
Dp11FIFCdP/YFQruZoUQuLfYDpXEZDOfmxDZfrssYSkIOENkmj5IPBiwshqbRT82
k+SEfTY6VqSQE9ku/qzx2RmKFoiZn9fIGLMiFHjQz4+v5qjbgemW7prYt3W+VHG6
u0t5wVTnOygyosjDwIlnh8/IMLUV5XAM7o7qNWXRu+ErOoN3hOMohTT+cSNUidkA
ruG/kkmAzDEvcFroSn/5hP7fB07fxJFVoZFO2kiCk1roLU2qMsYQK1Lea6Ho9Nwc
Gk1cXpJvOxaW1qkK54CODnqsPHUiSLVDfCno5ohZZYJcr76Bhn4ZFA+Tb41fqBB3
pZnJhlUsfWMT+Jfcs19QIcV8FS1sJLx5Etfx29TzlCPiI3UWhQzrKfskodZv/URG
GJJw+3z1HF8PQttZzqOQ/c+M2cbXIEoydq1oOsW84U8HlNgQmxgmpCMnb9oeBSkb
VR+1UsgDedcH5mBXY+CQogqISGy/VkkMMBDARGm4+rjtFVZO2MOnQ43aeDjQFjLn
+UN0oVAVEz0e8AMa6WCS16laX5rvO0XvAOoyNRJoeCkIKwwkbdYNDaptpmIH5MAP
L6FXldOCb4+ScyFuB3z2g9AMfubHe/rSWmyr+r1fxN5bK+wFS8+hoDPwRCmifvfW
pMPEyhz4aj7WuG9ubGsD5O86tLac3Jr55J7nc8YdqmKUSAh7WxbiO4fUHl/DFTfl
R+AgQSbnSaIWnVQdIBQWjK3ccwiNaeqaDVL9lBf6Tsbbas0iV/P03mXPtLVyaQpA
9tMlfxEDGJ/NSalb2d0i82KLgo09xHq4WqgeZhsy4BQYEleeIVhYGYfXhr8ROkDs
Roxf+Z/8P2I4iKkQuhDXiuVcGDt5l1QH4Sfe8M1/4GvbRtBexQUWQ693u5RCKB2r
4q+/OCcfYL+frBz33HtJkusFB7W+KY9rVX5/G7ENvYXrWjOE7ejWlIq3nQPhXGGv
Pnylyvg3RNFyjTwvqXvJWO0k4f90+4mPzKzJWydg+yGaITTJ1x/cI/0T6EDOpPY3
gJKCL9O2EBERkjZst7TtHpk/e+a2hocW7wKMuTkSm/YhiQSwpVXl9kEnWNnANvDG
lxLsb2c/uTGXk3txHIwMSt3ej1pjUSjQsbDbXmx3TNCFWOdIKWcFyHUQp7SqDaTM
jerhgmTXvjkkpWC2fQE1MFVQTnfpZMJs/t014S5hxQnX62RYATOsv9Uvk7tQKDoN
fNutp/T2VwdE49qnDRbKjSFbJTti1RVwAD6JBv4a3xF+GpNBj4GcS8uBrZJrOIa7
xhkhpwYyy6paPpvblfKU12g0ryZh5fHL5Ol6IFQpuDR5q2G7f/1dwWm4ufdCfevW
vvrMvlfVeSUfjHSLp/z3JnbKKtm9ph4VKvYbhiroFkIpZYepWzoOaw/tX9jqPQya
1vH5irLMKaXmOh+4J9CVRFZn0LV0M/TGVfhnVQYIdIpJn2HLC2AmxI19LO8d/SWy
8R41Ynxrim1IYWXCYmsNLrgD+e+GdveD5kewce0zD/sPzp8KbISNYXhLRvEmbyoY
Rt8E5/s3XrbXDkyLUbPYJEDb2784m7X4aVCOXUSHXDSLPyRr3nRz3yiI+FtILlNM
CaEB9zgxREtJn3xJy+TydF/TqdEoUn+N1JRXbCq1CgF4ihWGUrJUWDbbM+bAiAm3
dnlq6rD7yL4GPHv1ag8jVnQrLV2i0fo+UcaStDZkkQE9MXdTQfOPyQMuvRV6er5Z
IGKjbv0GeQ9oCDJiPFB/CDqlscT5TW/zZW3LQn4yndAPBnf9vIau+OasGQ477W3V
HApntmKlPTVzPuSZGoncUjdBx5OUd3MJrhFCMNAPo3e4s1v0pNPgvsKLekmwUbuT
rBcYdVxTM3L4cP6QPh03LYMDEJY4HT6vqtb73jlPjcBP0468cbQUxZDTTLGd6m0H
R9MLhdDlKMQ6360S+w6Dj3h9RBZU4qdIzWW4h8GRBoexKhwGWtZhPWM1NXvXRp6k
XP13BlytALFz5fpLKRhv6pT2PzmHx4AmfvRFw1wrl/VIVVEaMGdkUw7qp0a56EYM
18FaJ5H3WL9HObayjYQS5Bdos9nWjtUOFD165ZpFBlavHO1fcn9kv/86nOU3rLlC
yrck/yzKymv6rUh0FPaOMH+Bc+vSnOFmhYO/DjAEoxOSuEJ/8Pv8J76eR98/sRpo
VdPuMD6ac2PQ9jtT9+o9vHuUbW+HkGOhFZLAWryBt7tW/pF2U7mHWyFGJN2xCjf3
M1sjpKcnrV2S/fFimPYL6oVrcx7URB9559n+Zt3dj0D7GOafAHPidvjwyQBDlBS1
moRLdTaQWMOg4NNcN2REA6r46mg8gQl9BRyOcAFRvlz6xLgDIAiUpO+vl/5BIWEA
jmVcqM+NeXHwRHYkKNwvBZ1XYk+lR1d+Goyo/fAerZk1ldzfK3Gp0y/R0k6oK5mq
U9rm69qsyIvdy03yvZgrSNd0jmfKY7h8aqhhpFCxIOuDkg/LzWJZsYVbuE3Pic1y
P10SFIIcbGRSrde7Y/l7VE/f8416QEvdIpgGrel3vi3U7rVgTalKXZVveGrZZdVF
AjSbIEKtxDWX1AepLatO3ZLmhfvOPLPWNCwY5l+94wz4eI4LLpFwFjfmQth0Cz5x
zlbiMVRnXl01EbxMqtdrkrq29sYQC+3iErcbQ0EAUKD+7/CGGPUM++vH9ms31mst
Z2HR+9M98iV4AbTuQ67eA2erJBjqSQZY1dauVCqOUKsvkONPV0DhL9lzKAU+ZUlg
4Z+VeDoZZuFCOrw8BcKG9h5Xrod87hj3NZfdffFbLDGN1pzPWOpcQo9VspM2N12F
a1Lg89/BFeM1g8OxCeE2dhcB+bxCn/q9XZY2EI6AgfQod5xLISvZF+L2ABKTNXOT
KwzONPYAcKINO9CTk5zZkHBIEv49fZ2N227cB07RgGG2a5jBRSFUgljkKi5pzjAX
H5ShkfPmfm59A5D/ZEfIP7ICLL0uuA4eXBMHC74nrnFevjkTEXEhJqQaV41711kS
eYFmWBkP5jhVpS+X2+EMnRvYSK+cmQZeZvMhMRFxmLhKSkbBi5+tePF5hidniebj
Zq54Wgr+ld7FyjNLtzhNi0+Xhp2HzEs2DroyDj4Fsn7ngW4tOim9W0mGS3E7Z0eU
DaKewV4YrBEnvS8Y7nsM2kAGarYFpv8njNokqkmQc60QFav0jwMr082lKGltCuss
ZvMlBLX9w+wUP0zxlgYqeqHKrDRlui2+MjDdu9wUmZwUxXBHTqPkz/fQRPATcYjb
07bAW6fmPHpJOFODH6YZRlaATo1mLDFpBgVo+EwIflE7PRhxdRx6CQOJ2KKTFHa/
Zd7TCXeGURvLXsELWiEbPf9KQkImDUs1KOKtfAS9qxe2O4nP37uYBLpGFQrlssNo
UINEsUwAk2Ppv4h9mh0mVnhtAEBgoyVp/YS2g9JHakFWwQBMZ4lSpY3RHgr9yORp
gYkvWR9ppXt0VKff0XMMqe2biFnLOczU354MO+tsN75WKtMLWHPvwwX2sy6my6m+
Qyj2qfc1QWHxDmPHr8GM+pzVTvLELtF8mBLeLCd7NVX6X/j3VrsijoXO1hf2hgOE
qO2FAOM0FAQB2j7BCS4dZlCsd5EESKgGI1J7Rp+hK/G3fNesKroyq2/qzCQbgcQd
+RAYQotKuqqrkiHKtcx+XIEfJRKu3utMIRMhlqInTjHQcWOSMY0uhvEnoOdxhEfJ
SV5Ko5oqAYAUYbbP2H7UwYqUZqqCdYgD7/P7LQFWkRWM4aVWbAkwqL2zi5E+CQIo
dkxtd3gicz756mkTBv2kiQYMvRPtxGRUrNvR9OGkuWBw8Tr2XELXDxFhcbVvfm7L
B+e/tW+k+GnqvPQeNeWO6Gz7KIBsIqvUqNb8t5G5twI9WdtO9KeDz4WSnIiVU8Y9
JN16ukNjHsVPLqjg04XTP4lDFp3aqHUqqJVPAwIOnuNJKZkJ8wXfHhX2oo6LbTNv
K4gKi5bhq2+0w+AFHCmuZADB/m6kTTVZaxDuj706ykFHCtY9bDwy7U33jZPkfzBP
HBzkVw5js7q5Yjg8Mf37Rz3m3a5sIPx/MG/GzyAvbSp5hTnSV/PnVwg5+WkSDBtT
qjBtpjM0PZ8Z3YR4c1/g574rUFBZj7NZsR03Xe9dXcybehW7Hv1OTJor0YJ2oDJp
++bfJfJ9mZVBJj/R7FrD0M6AkdF9ft7PLJY1YUz3z37QdZGlnRmrD2OdZ0AcnMGS
OmdCSeo9a9FRhqLWjyhteDYXwXew3F0xyIZtekBstJDwyJCE3ZBRhmGcdx52J6gf
7fFETG/kKynapGzsSxvqyNmdPlBSdgXe7M/FTkWizzKr6M4ylIegftQoG0eFpYQO
YT+ebp/1CVupHrFdOUHfTxNKqAo3od4eP+tBwnE/USTVs4h2+vmIomkVEPDG2yTz
PPy2k+zSWe9xn0WWZsxg2ups4yeRwAWeU0EuqDZL1wX7ThAGFAAXmQjkaXoG781K
M8jYoAQAlZ21tyCzZZv/MA6gUi6Fru9fE0E3S+kRepwVA2I0n1qXnlfVAUYBg29P
xhbvQuLveKfLGFUGhn0tDi5h3Gq7uT3jDfpSgOqIvd+UBS5yuIL1mecHLcBh9Z4p
UN109aPYIEuP2buGAfROe9pq4RJZDcnLDxsnTUB/b7PkW+HDd6HDvJz1Fal3YHlC
oowA04qJnD55rIIwPfz2koRhrSRnTmAc8piPiBM4mjLDixYI4yfClgbpDSRIJOdg
2/540RVLd0WF8zufZzqmVG4PB+a2HBisFn58SvcUM9QSwEJbIFXdGkKQmlLzJXQ4
4FroJIXtvmiFxw79KP01vsto2CpIkDl8HuSobK78/riUdVgUqc7BuXnpG/HaRznh
YsnjKnyRby9wycREA4Ht/hiBVDAkZdVkp6h5U0VsVeVEJCCn+2k91AW0o/MoxCPI
dIEXnwk8qJqH4gHmbzLPKPv1L+aVxEYLoy04ygcYHHEzCW08Uxkm79iGjDEnrdEp
779Sa6P8Ws5fiK4VzofXz6WlE0EpEVULhcE9ScO0T0XjdXVsT6qgb01BR5ZBWg/L
MzJCnyqDY154oR/X+5PjJWqzQHyu/l4W7kcUrfM+pfiwS6NJ3RqYgYMrJaEFMuWF
EuZ5XOtx8jM2GCMhggdH1evz0BvVLv/6q+KFQ0yx2e5mFazoqlfqP4jUr5VYLjte
PMCjoPLG6wTlUT0EpQpf3wAERIsYMZWMfiEyYHEoBs09NrdXBPgMmRdUSU2hZ+Td
Er6KTysGlOdWFgnjVGd1B9ITMXCqXL+NtVhYnPzIiKtNl/x/dXitsSyXNJwJJx95
v3DDT0NrB3SIRs+ZVLRzYFPCdARQ0f4K9hXaXznXo6LDnjebZGzgAWEDK3p4V32J
TYHCjHmqzWWnM6Gg3w1IKrLKKkbptOUVXr9a2MTd8rWUoUHFQUeDyniDB6zwaFiC
l6IQolZKVxV7w4ukkdOnGYhowCdYF/OOlMAL/xlFpfjhVKvkxLwlfYXG1NeYwi9B
JBK2tk2nSGWYhgrxJrkqsxY7obppcZJZyMdJEdjMsovB4ECJK7db+A6MQ1GWjNPc
YQISEnEcEH2MygdKP0mXwtC53cUxF8MmgG4YZXcuuT4nHXTZpfrnZBZaKgnUYp4t
D8izXDWGsFaVlQsgmmBJRvMh0K43EL/vg7wC66GKfhzXRRfQfJDyfKX4rzjclnmi
SA0tlmxEOI+FnCZPvlggdk2J6yykt97e/vbRT0A8xRyOPciGdD3/ATzKM5Fznz2s
mzd7weNXbRp2gRtFp5NKoORA82GJsfxNUGSC/VNGxeVIzyYU1fQSCBXwp1BnfJiM
BQrWSK2/OhopnCYG6bFJvI8Hn32x+s+MM4h3tXKvnxR8XMHVVBoeIVUif5ZY0KZg
DywdmaAtcvRYm4kTXo8ENkhc4ml7MLtL7LeN74YpsIQZI9SgQdntb9ZxCTBmJ9zc
dTdBynEr6LtXHaFbVxFzK1TyGmCtgPq5ZGxyRvTAerCLsi+xV6WU3lI9pNlGHOzY
rFMdQmr0jzgFXGzjhKgtGZLcYFXb+V+cC7e8JoxaUTuyzn7s+59obdDPH0lRX7Ol
qvRE0/EPEJhq1Ls+M7RwOhe9cDNgTARLsEwW45wAnRyI8OWzZR+Qq5tw+Z2PGX2B
KFzxQJWKPTpppNj1ZhKs4F+a1dAKz3yH/ZyHZiuuMQIEfPI2m07cOZpW8sZH1ek4
17gs14127vJlgxW64vIdrCku3RQ2nML0vFYKI2f6F+M9RlYYgbOYhR9up89u6O9z
KEMVcFK3p04sjlPYpHJx/TKcsX/xskwWgQd2RK+dMwO7fiboBU3G1tSJCUfkX4/K
l6IXC+QYxqPNGvgvOz2xW+GsknpspmFGreMdD5ASjnQAnMxa0GZaFlIKpodlLnUL
ZL7YdfP8zvFMRl3Ux61DjZ+1PWMAirK0oP3X699rFFEL92oxFNfF65wkq/uviOqS
h1Vaf8iGslELoFotIh0l9qy/zDJd0DQ453KZzSnJSAsIj3R7iHP1KSRncQCNxuG8
blPdKBO1tO4ZR3ZIg8DOBeiNr6hCUzmXKy5I6+zk5Gkcdk8SzfZYOayVYwWs9M+x
oCsN6jVZt6lPq9XHsRJOpCY0S9EWhQpkNT4UoDV/8leNItficCwXhxX6523S4RK8
BB7wPKKZ+tVC+7ft1kb5RStvW5pd1PDZeLCMxhaKGbzNL+pjW8AoBXzIZZUb6YtD
EhNf2b+9BDwlfihDowWcHob9s87hldZkm2EqP29yU1SFwbORA4KNcue2PI1/YMvY
WrhvhhuzWNyH97wLU76vSyQNuEIi7NIEn1Tf0J3gk5Jq1r3oK0WYEfQF+9eVEnLA
TOU/Wwy7vDaHGbABtYRmU15lsr2skXjygXG9XOwRov1KWqlXR3YL3HMHoVU1/WWZ
+hP2Sq+IAVA1U78s+OVrVltcMUIenn65aas52QU2F15vHgHyEEhvWjppJ6HyzMIS
QbyFtuuam3RMUeJSyc9XAFTPKKzd4CvmTSvkHo66aSkb6UzZUwFrdYt+4lYjfAHr
h3La1VleW2gTU0ZrZQZt5v1gPps20lIAKxzRDZe8DxEUCPLhLtcOitV7zjybFwkC
fbB/pzQzbVAyJbEvQUEz+Sq+rzC59tt+7WZEPvviAyQXv+o2XZFGTJF75wxQ8KXJ
b8teKlD+Tcy39v/PCrqno6xuYZxbK66Jve/actNwwj26vrzSxjY8jInPwwbiTETF
JjjDJwzC7q/d9KIJAuj/pPthBZaper23Fdb7uctRDb3p9xr2GNWiRZgiRkBo3VCM
zdxvABF5sKYfWwHa3kb74ksOTcmaX5zym49/foWxhrDKiUr8ORBb4lJivw42cHKU
uhZU6WsIJK/GBDHFXl7koWKMSbBKAp5NeQlZThbeveMa4q0iVzI2gz1tz8JdUbck
R8Pb34OvRc1zdxr6DGFJtGhhB7mkedJXLJc7TjfRTAXtfhbIO+3D1CKxiCPg8sDK
IlHY+Kn3xkl4zl+7nuN00EzW1QV6RMrnCvydsOwESWM+9I+ZhexYZHR/MADfibVM
aF0ryA6c/1xncTEtMBxcHWC0pWGXNaDpKOGb6+NWI1rZh0rPdYkKicbInvfdvMyd
TxCB521NvXgfIGG/GXcyIPVqRpSzhz8ibN2TXIHRvhgyZPkh+Fs7agX4N5Hg9Rl4
H4r6UFKw6L3dYZyg7DNlS+znN258VuO8FADf8V3bOWEfXeMaJ2yQojm2LeAP7aBX
On9FJYAjjgOYd6lOgsj9QEwgYEzdDiREizaBDL65MFz91jdNguWxDy3m7Jwjnmd5
Uk0s/Jt7ELp0sfR9fztvHNbPhQB8YTEiGjCucwNxrPVoX57iFCfgOwbEVJyOL+bs
YNey9z1fW0WlT62Pzsef98Kf8qvrNXnFsezQvEX6zNFVJUrr1ZGc/RVeBMBMfcRV
1eAsWmkGYqHzKJYvEOTBC68U3SJBvHZCgNVhzp/D7BHrrhfgAle85t1oA3qopr0T
rz0gtBd+k2l0v3w4oYa0pk8ZHFpYAKGws7WtB22JOBubieO4xrqIL16v9RK5dJCH
k9TS9ZAqIiqo/Bcwixa1FBUKMulNFXLE+9eBdkwZoc95FHGbObx8XZ9k/Qn44Yrv
Gq2lPaWgHp3+iMrk80zk9PhbCICCOQmRlI9WqMsu8q6p7yUzl6/pAl1co70Y6sBw
rEjr1DQc0Ro/FvZbl5j2NJhmUcVUmgQ0KP4YSbC7kSnSvlNpjzjd2Rxr3V2oVwW0
D5QKEeBW59e93YWsbiaRXHmQKTji/dYH7QA2IBPOtPwoNTUlK34KAQWJre/Gie+A
AWJI8XrVqqyNvfP5VCGhG1EVk8JGJCZezMbeTLoxDZl7mKWdXfMaCGxXOr5mmfv5
cgvnQjUARhwU2Ealxf5XJmSIH25ndllzouueSKksHgn2AR3KTGw1jpJllPtHndnX
OdxvNsZqIIbaCG2NW5lUSus0qa5mc2fBD4OSbjKmJbb8fZz3KcksEma6DmePr7lu
GKUbCzpIs3RSOAm9YdOitdg126k7+ougU+Dl8Rozf6tFiG8z6+ONOa3X+38bHs2Y
cVJQHDtiZWeQl7a57ItNdNTJb++/cJKB2dG7iopwJj9yALNrYk6odsMQLIRyVQVU
TCc98wQCrO7a0PFJi9r8e+AGHM5pU44g8yY0EAGuoUMfPfR0dpVam/1LGrlSSTcQ
CGxX9d//AXiMSTu0zw/7g4k3TFStyLz/r4lq6r61Tpu6jJNGwqFNwuKUdDaNNErj
Liet4YYMVRdEoJRmLvXrwUNIsnR17mujXIeLn3VnCxdpC9lEbEx/89lJPRUKbhBW
87mSQSi6W/oLgYxoAb8ulW/P6LrOo+mi16iqdwMewFdX55ppk1pQseiWFmU3A9r7
BjWBhS5f2XE59ilrfAywDlAXJ/WQPIuZwRykFnJTf91fXxGvTOUDpILCSTK/7g9v
Pi+qp4wRZShGqoag0d2i7MH9sJ9CTjbjpd6Wj+ApQQZRttodBwME4O7e0OSz+n4D
Ow8sV1Jr72hZTdaSj9uyoKDSz+nrd218ZhRt6IG1IcqcoeURq+BFA41ZVMyTVLK9
CF0DEw2NfoPKW+I/PgeRGHFVX4lY1yCzeHuPhxR4YS00Ybnv0f5tVugQdM32SDVB
3eKbFQ0N+IMgda+p5nvQoZk2mA5C2GfzfmhWh9ZW6kjFUX8uK0AdQ693f5m7AZ+t
vWBbelJKb2/+ctQkB9IEuhDedQmHitxcbAG5gH0d4eXpV4lUIK74Qdlx34vO0wfz
5R85T9EO/QxmHUjDebO8Q/07DXq0p1cnv9FuVWwGQb6wChekQS8S5M+eDCy7s7bM
ZCJaMAZcsO0VQ96MPtLjjfvsyG8TSZN6/QgsKq/8zwAkz/joJSfRI/X4eFUJV6xv
XQxGDsetQUy3tSPwdxxe+MzlElUjui0erBRWn7d6LnpZenyraynBvhQAdgyHNKer
E+O5foavgd1Te4OyUWB2k9gQx4xc1iQqcSXKRL2HU1CVBp4fEJ6g8k2RfqkZjT88
Ob7RwKFljyNkmEfC7G6gMgSkiCuOutuOGTUFAc5W0p9XKv6GFT0V6M4WTK6YLkNo
qMTcEckrzVIzoGie/DX3rjzFOCt5JqcRQawLklzgjcPfuHK3SXLeM994cEWTZkbl
fyhIuOjO17vgMYileQ+avMlHM8Yqmh+dEb2ynvgh0TZXwdtqMxAS9etJipCY7xHb
TDuQ3wE6lwhEi/OZamqvz5VEo7EZVLGRWqE6HXXBf/xux9UHiLpnKVS8KovypPgG
dv3GUQ9UkqJnnCxZD94oo+wJG+MeAftaKe3mtbCxfUd/IcFH9oB//bxfXyRnFsXa
BBWANJYhqCB7vnUenLDGKkR2DkFXxyZ9fdr2Sfj7MGWu0ESBz1KQIRYB485pfi/i
fHyOAJdzmYiLW4lcaz8wax1EBazp5nIZI9XrB7a2vnburB5KqM1JMpBMDOu4a9QH
caqBC4IKiUzSrSEEYafMBYztnK9PndjVVO/bT5ZSPsROVijqVhmzwQ+ZC3vnuRDj
IGIJE9t0po+/ddb2VcU1KCxNVz7DTTTi7UYzgeviKUUlF7FsMXwcfDkDq2qv+DRK
DrAx6v5KPjRwkmDlWWUykXLwIbF5zZHbyf6COT0omv2TZ3VxaTkBMG5jEnWqlH+/
WD57Xz0Xn6GdiRvqw8ZnG/PDZoKGM0WB4UQlJN8vQzdwbfDrsrTAL0r+pQGlA1Yr
M2wJbaSP5OsOgc1Z+Vzp+SD6ecahwFR7qo56OmRLl99EfXFERPHiv5+LxRYLdfBw
k+Gu+OvgE4VEme197sC263MVaKVRFr9MyZMA/k00plsnYCaUQAp9301z5T19h/R1
POffvKuXllDFOwo5quc8udQLdGaJCI/pFd1pQpmBs4MPePE5L+HAtSCFvk8H15aI
Ai2yaNGERKpIQSbKfbjJM21nQov9O5DE+6pw59kY0bYZbLwS5+qaAfDyq/IdkkmY
OKkK0kX/3JiTstRryyNz+s8M1lF/vAajlCqLUUt4zax4KCzOR52Tiiqgfxka8lqR
g3JdfjMLi9B7hKvHHmdssgiALRmT0JxAtPcvAWR7qYmD43rTBdJX1WTQLDM+9Prm
xOn0dO31ml6vK8h2/bnkf7MBf/9z4DzgocBVmvv04ZoEUjU5jRj4r8ISHDTlGfnx
Q2SoTBZ3XtEeiTiru0zQiBzVu49CXtwUq445yOcOkTEnBjFKg0JRFL1OvHGo5k/a
qZUTQ38sERbnOCIpUhIMIfPBiUUyeXTjxgjLb1xwWUTF8FWVg2UgqEO82gKJiF5U
AnUyXcWXKFU2MjmraUEx+l9ExJuioOV46XL9ZnKDGOOftVhPP6pzdLGh8VX8dGR/
/TsdeJGdOcc0RrTLi9MONWcOScioC2k6eQvr0IhbiU4FdXVXP0efvGMpX3mMAKlQ
v62KQnQuLOy11WKTXzdo0cThnjkeSGB4a2ITt4NMo4uvK25z/LYO31F0hHEHEdp1
3iBpOpU5+itb1/RGlsA+nOn74P9RMNiQGPwuB0givQXJgZJ+YY1zglIoD0M7KikS
xCo/FoLaqtYjmA1Bu5536eDrw7g9YSFF+jqh1qJx4+E+PysVQj5LED4NGjCEJwCs
yKvR3raAD45z/RqECsFTtD4PEwsAc0jmhAIi2QmPuA18MxSGm6gGPwiEArPp1lRN
h02w+Ymf01QQ5Xyw6jOH935KeaYJntXX6ldf3QeEaNlTqfMRQBgaO1AHIa+QB62J
rMbWMziMXEnrRkHhVxPEXDXEcbleMrjMwKNHSVpkVqfWlBU4l7bHrIJJV8eJWVD6
vtg0BpR7R6EThCrLoTVYIie34YmKoSc3ModyYMDwt/8zuw1roMgH51qCG96jCqCk
NgTfnOB9F5gwYLUKTvte8GZUDWCYpWqU2yPE8rRErS0fGTfXDz5QR2uCYSsDFcK5
C/MFnYwaZklS4CKgY7W/qxrjx9LzNM1ckilwUJw6oAvNdjyRYp2+Rk0gQFjTMvXo
BwruOTXl5DYs47LmGJpXqBa97T50MWrghYNfUOzkfm2Fh6HJrOblAUCsVJ5vfY3K
3Gzt/QTAqBm8SP+aIItJjDOp4uFEwwhqketi7U1Vi+DvCTf93JGL0r5Z4DVLpme+
ccdxUBOQfTecMzq9bfmR0Zd/3FMJUEixBKDsHrdh96p56mrpta07QXhDZkDSgtWB
WnDaySUFHwpU67PNWD2gjdmrBO3TkdI03M1uRC3aGYJgsZYWW9eOdTJEk4xdWLk3
4g8feTRbvHoQlz2PgScuSRqPj2BL3nxZXHmC3pAee0Zyxi7hZY3Hwdh3im6EMAXF
d584+zpa9NFY0xrLEazqqGiKuaB4sipVfhFuRZs2uk23FjNc/GjkD5rZJDeW/MhK
v2kts3N8oeSJVmTJPTMKU/bkVe70QLQfRXHpfFdd/8bdCVKhJUuYKQn+ZsRsGgo3
4PYYCMdUW6PqaAksYemB3ZooBTyVFwjraip6qyBtRCOLesXAwTZrHInD/cZSnq1c
StMQCQZOXZmsRkOj8o00oFIMVmsOC0EXA6t2XetPukQUzZwzTrc+DFGk3X4r51G0
1ui0nyS9In6x0srFVWCx2/ezU7MhD0Tvl8celEosL324tz1QupUe2USP5IpNVruh
wEBqaj46ucrdKN+WGLFHKNV+6mg/elo7ydaIcZMor74r//gH8PdIQenR3G2QgEwu
bX4RZ1//gHn+136EOt5zxoa+bLaT8h4vhKhF5zI8f7lbYZ3vDoSC0W7b7xsmBAuD
9OG3PmSmprxqh4fZr4PQHQllrFIF9peMVKhly/7o0mY3otJT/hXP/StdwSxogx0t
J/SWFERCVHfmXh0llf9T+HGWasIfS3TLvEyX/H2eZhPei+dSlpomt/A0E2sssvko
rBv04y6nHG+TjOQX/o4yIomEkIZ+wOCS7m2/wiiA8hA0c/kqIUMHhcjCN1YRxgOY
LalQK3pjZJZYjFJ2MITrgaIGCQtqyW1YgD+VLbSHtHW48HGhTn/2VjGca463+//1
eIRvESt6gpvGCSAhs3tRlU8MSdMTiJAH0Rv/Mu+J5Ta3erSltXCdqRCqkQDCSNcQ
j4VMZSWqKaomgcmZoFJCNRwUt4XLxq+cEOeaTf8g0QNowV9oSHXa30yX3TiaGYJo
fuXq4O99BSongXM7crDkbz+asdjcK4mKZcB00jwWtOKIgYilsqlm3k2qUlDMMkty
Q/vt7QnF+NdKWk++GcIS/S7ksHDJnp7QFQm0sRdAC4UKJ6h3sudvPDbDMKU1Adig
CxqkNHrTQvFkWB2/2xrtjsq5qLeGfS7CMiXiFqFa/cpMIdmGGQEPOYwOLjnSZUe5
e5S5NggVGVMGoJ72tAr7u/cGqY7I2j+ZmBASG494FVptFgnPmXhKOdb63GmCALkl
wM/3x7ly6OsA7THmJMtDTSmyb7EofDnAZziy+YJ2rmMXsnwln+zSbqdxEy81x2dB
wxAS9vzQSk3xdgxiVrIbACiSMXAC2ANfDb5GNNMklxpJrgoEX5H53c2L/C84Atth
s35d3u7HYxbFMQRsIe/OFNDZ5W2u/rkiRa1Rtn1ryK1dqB8dR/tH/rwdiNcf4++J
hWFMI7hqLXBk/9LFPOPOCXlTSjg8NLYuZ0spWZzBl38z8KdB7rtIhG02pPNTMFUl
UTHcPKHUrgJfbG73T98hwlhr4ssDoNkw6ZwiSDRBvT0qs+5NFprGtjrNr0Y+yxNV
6t0dLeMrtoKxc0SIRwWc8Ql9X/PanCF09hmJKvEJm3K2BCPOPi+qq3KFNekVW929
zZGpGoTCa7u1Xoxgr9qObkAzqZrnIlwxpS+ragKtKOLOpy6le6+6EMt5GGcyYlbE
K1m/jo3BNd+EPM/Va8twzVBfs7EFPdKjh2+S+y2rpGtBuKHkb4JiUUBhSZWHqMsm
3cb4yz1VPhtaaDdyFmstbevyxo43xXpJb/wj/LuwyeSguvPJFFWLrteXhYmVTrAt
gy2ZAubIKlCMevf1KfQBzzmUYbLUgn3IZCs6RrFbUm3LQfnCRC8SXU8hV7vy2fis
Rjx3AmkcKBq7s8QdgFOnogeS5iKBbWp6D1sJMbwctRd5L0DSX9Zfu5Wm1RekFKc4
wpkHclfLGPeZ72bUPM1ecktgmVgkWGpoWBb3zm3VdKdg2AVE7+bkvEKM5iOgKu05
/kN9BtuXIiZwHPSisBQqdz0QtImW7X6NJ15errwj9FtGvVSf979azPiQGJ20+Y2z
XfdDASB3xBMW9mAnNcHPFIcAH/rDyneV5ziVMywhbKG5uIkFbxHy9Ml/DGOfaRET
c7m1XvSG3GpMDwRNMXb+R6r18Dla0x/Gg5nzkVtg3ccn2DbkGj/xHRdhub+8n0e+
dR6wX62qG4nKEUrDN26vhNlwGxDYjoHCNwuuDZxneRCvZ7DUMk4omTCixS4TX6f3
MEIBr+uvNQed/TfoU3jthX9X2c4S147yCsC2oWzo24wlvla/FWu/UNWTL0u6uCn5
uV0cdoOyFePOE+Zo3nk+VI9/pfGU2qQCFFOZ/+F6KQGRpT49ZIgXqG0co49ONR6L
jyehctk+KJwPg8+xtaWT0n8rs/iRb38N/RLdtv/r3jY/K1F9i2ORz0sUIdF+CqTG
GdIqsatgj2ip6xwxFWFYGO2eKjZgKKwLFeWJsp7vHEZYzQ7dqicshGWjTHWZngkt
SulO38B7pJ4Bseftn2Kg6ipt6ArIwpL9Jcp+v20bVUh2TFxhjX8HGCLShTg5hiC1
0R/qs+Rbn1IbXtlBAnVc0aOBHjO0mAMHyJehlu8QmDofFGD3XvvA4dKT0OXAxFo7
zdUS1rL1/trSBk4l6wQX20CiFTujKUv68kLZrajyzgETKZtaGyEUledjc57KJSIQ
5QUzK06XGZC3Za2ty0shzaiXmFFSywmUinbOQFE+h/W5kkWdM5h50g0W6DAg7B/H
LcQFRyp1vm6WQFBbyZlfwrVREOb2ep+YnniDNvrN8wv6+JeIzthAwgEB8zruts0H
ym0tlbX4fR2nX1bFIjNBdVbMBLUA6lpW4siXxhTdAYm1Lk7JelKHKG8M+g6w0NQU
TF4eBAibwLawPlNAdbb0o9itgpW9ivrhv35Mmpioz2y463DM8hkymi8L2lyoF8h5
o+BN1P/w0VbY9eQ8Kgm4GOFO6jYWGp1AZqeowI01blrtYvQkOm7Odx2nfXz/kpkL
uTmufbDP+/blZEfS5J1oAxncSAqqhuPllNR8Y9bjzjaBLtiOlTJ0AiEac0TNUKK8
tSq9Gkh0hRs26Y6CRZqpsj6smKmCcjXYzeFst7ImeOGRgumz8W97xx6stPvvYKLV
IR4+a0lmOONKiI/RCP3ZZol+XL3CpwqNUJRHIPzZmMR/96OKu9rkEpIpX+Sl7V2b
BKNeyWI+YmjZ7Aqj3wHFqioldlot+becN+Lkgy/WcmO3kjy8qI6fMSIcpgfAq67B
xiC/mk6VJhMzkfHN/HGTF3oc2M2LzMaQHVOQ8FZ8mcXrDLUa+KagSHmOp4nA8X9w
aylpZqflgC0m27IPKW/PPlFrWvWuzbgEAFS+Z7+lqXkUUHB9f9UIK2udhsv7zj09
DK/2tkXHxfOYdIIVKwhvVGajTpIf7f0qaOLU3xta0BwZB42j8X3GGS5uh5uimBSe
7IqqOW4LZHy1b6ozEcglZVnQpS2E0P1643+dAkxFjYTL6K8iZqSm86EsJpZYwIlh
vjPRR+crDbDRGVdOn6HfZP9lhfYw6bC+GAa+qA8y5hXI2jozohZxJO9N4N22oHmN
h38mwcrwaHYwwp7pIts86F7oEDCWg3xxUbfBIgxk8Nze5ROKlZ3tpThPIeBsEiq8
rzm1h9akVand0+jqv+RfzgeqIrOriAjkmZkGNf/ABdnuQ3/5rKy5wwGPYLSFevpq
dbMPoHEgHIWy0DcwMCWQOrSZaMsDWO2WGb/sg4HU3Gm3TeXnPDUBFzuRH4T94U08
+xF9jn0EwMcgn/2iz3eHERYvuUEHIx3tgcXWGBqiwD5LA4KeRmjdltr44rfaljrZ
OPGt50LU3rLs7FDh2vNKNdhvdcbBoOyu5049GCpGSppJy3qcl0nbg/LpJIDmfO1t
kcmQ43TIiH6fmiAgjmSJPxlCwORMEbvFGc6Nv2o5JZrn/cEsll7u1pco3uI2c21t
AulvAmevu8Z+5/lmyxj5CXJAQ42pt/tl/MKImnEblkw2FN149k65v2NmYJu+MKN+
UB3/LbaBLLxcPd+c1jLuyWjL/HAVh4n7z/BTSadZg/gbQb82f1Cs6+nFflYLjuCv
NdrxkSJzypxFuo4HQnKl4nemd4o5/oDKXxVoLvERSYZWJSxzHWC1dMoEUYXEz1R4
CN/xKcxHt94uixX0brYRcI223/CC2c1qZhrx87zbug1QK51hxBKqYF+mm/PcMMKv
XuqhBIRPIy8iG8ZokJYr1z4E1D9zhOaMfimlQrMrEK1qdmgK3V2DNOT/HG7iYaZS
FvxAQwXe7kXVkMut3jBJRHqEj714DlRmHFgJf6IFNvd0oZweXGczdecfcze4UCZb
ZxCWhy+FwVOq2vLa6Ho7sX2C7MQA46WU9r1dVZGDhlcU2rzdXcaqU0KvtSKFw+J2
+YHl9qW/ZvEFs3Y/KbPPHmDwO0VyKKNAKh0O1ryioDieb+XPPMY99jhiJEYnFUqO
nZsZEnibI/u8laQV2LenMj2vzHsi0gDMiOQ524fOeGZAkK6n6u0gEh+xv/bRenIQ
UxH0b3zpavBQp8wBsvgpciiVtqGn7HOe/oiSOExlvZVcZbB1f7Q6RPxKIE1xWtAs
FnbsW29mfn2Egllx7YJZpmViBKz+OaRHxhlZ8UKSBNcG7pQ8NoKvU3XgB7d8xD0+
QBMxerNGKLCIy/L4BAccv9zc2hX0gUkFr86Poa+m4TDisYBfI8CqUoQxFwp8sFls
T/jWB7PCWGQy9OEBBNHo9PXxl/gcZepcSn2gNeV/DZIVEuloZASMPMhYciRq5ast
piBqJJn8AqEOwUuZf1XuRDR4Sgor2izSIyXBbx9hsU4u5j661xf9U0C6hsB9AW/U
5QxyaRFjB9h427eiDvCZVMVomBP+A5X87/tlXbh9r4EeRCmZD3A3Q3JT/wYS5NY7
D7eW0+BouV7/I+pmNzU2amnB24VERMLS7gWXL0MnRJJQxuH/p2C4zO4fhiaJ7g77
q3cdYtQbhTDoOO6BrfKAB6pLogKB0Rk+bF2PPPprymFjwKEhlu1S9LYiIF6EdL6u
1HxQWZfrVq1UH1dmwfl/oz73Gm1pGrmJzt2ENwtq2Z1rwldrpZ7Zs/JXKbayH35x
8laMzNxRV/5Q5y7OrSW+kIAjbHrGZ6D8FUISkkMTw9HqtKnnUZSqlYhGnLBFiElC
nOKyQO3IevssBp+LmTPn4yFw6Z55qruLhaWN5XK0aO5AKONjdyfhZYxp31PrX/d7
2nE0hTxvjVMtfgwdDMYnw7B/9LRJ0OlWhHadGN/RXmSs3nW801+aiJL3As9LeEFn
ILnWrRuKkJ+MDZoNEkbm9Y0/z/A7WRpjocR7mU0vJz6cCAz8aNC8Cbp/eRPXXfvg
3+JiSNoEcnGULV49re6j1AB1k908e/Zv/COfvvDJUHaNtvCTZqHB6aGF+laV41kJ
PkMML8qn/0fgqxvI6t9K/D1e8QevXM3bUEj3yXd60CPDCGUA3oTZvRItdhuPq6ue
FCoxLgV7M+1RvqCwVsHFepFEMCqB0KM1XWI7KFOAhrCR77rknHv3nhg4jpyM2uQj
k5qTRbheAc/jphHLJ92JzB805FZvlzEMnqx8OxqYel+0fH3JJ2Q8m0LJOSs2zBSi
OWF5LWaUDwquM5TDpgiuoCj3sHLadu70+d9+LoSX7iFgT+iy04xrKsFrr5IUDpNt
sQNFqrPaFEShj6gnhkBYbfmyNvQzKdazUKQj+qnYVgriGNkvQiUzzLfo6h//wM90
JPi2JcgshahnSGyeEThUB3KEaXKCmpM8dc9gxOH+nx2vg4ErGduyu4l+lSH9lnha
Ho2z4c7zdn33kRA2Dsk59SM6u+wPSLQZimquYkUFKCdeWn25Z04j9M+40/Ans7gG
1bAWbiHoffYtT6VLtcBAcjDk8EahhAbdyjtiktDLXTJCiLqE7JFqMEx4UKl5RITV
xY57L/YbEUA/NSPQlP/ypNeg/p35Dryxhc8Mxnyu6AM4KuiEhbH5oRLsdPbkB0lz
FKgXq4JVEN1hICbUS86ccLV8miijFZzLjuvv3kiUcBGJw55mMxXhM1u951Ig1ssR
gDNq47dZhvwpSO9uwNG679RYl5APP9G5LnuSTZ5bgXa0xi8VzA0RqljaMBKLHxn/
II6pUi9Cf8RflfnEIVIPtoTadfPzr+LxthLszV1ucRTZVc3V8F577abm3vMMJ4/J
94GX0TNNXt7a+gaLv/h61yBnAXCpSfwpkXToOMOFLKMQ7sWcbQpxn3j6+7nTIxyx
RvIpWnp0qFH9Na5an8usaxOGGGlg+WGn+jmiSwcA5z/xHFb2GJhca/Dav3BTv8bu
Zb3EnyNFpOlDodw87AGBXI65n2AEtFbImKne0bBxn6mZbZlg10UlWJVxC0+d9CVm
k9Ay8kMi8+gB36FJEYn/HLN3AT2SEZ40GJ7QEVkEsYQO5Ey1ScfSbUxd3DIXEa6l
MsecEIrV9gkj0NQ4X4qzJ/yn/orPr0niSH86RDXIlGzZUs/9vhIPscQTfYyTx20w
jGfpHqwJQA8NgsjLc5OSG+qLOMhNZmCqueSSArdbYLw/TpjLncuZeAiT8D390E5R
ny6BgEReHh+PqHoR2098cPNb6DkZkH7d/cQqAch0TxmK81ISvPI+BWyrL2oFvEmS
mA+84UC3afzeaDfgCFwf4K95qDUoI70JsHOhaAgcv3GQh4p6k7MUdOUN1eSifNWA
EfxavsZCuM1Gy/DA8WxwRkGNrWR7LFIzTB6tI4XdkLutMy/uinXabjlzDkK2HI0E
TI75okRNr32GSfRDSqZHbCTR85EfkXDb2RgWnwZ9RxhOg6AwwMhUH6RZRyDAbZQf
LFDEMEMID1nsp6n7tkSC3K2GcxApNUDKdMvS5ox/RKA5aC6BlD4Z/krYHlHrWoo1
+ZflfaYB4lWNo2xmzfAbble3JS/msvxxe0yPKLcZiZvDO3ZC/f1MbSjPyzaSV3Sx
0wE58EFYONGIPqh9w8d3l0cDXIScfF61xi29tSas2cGEiSIRjnuXNP6NdmWMat2t
cp+GoWnDgV4kXNjpnIv1RJKHa8QRgK+jTGLeI3ri4yA4t673dyvFrues9BbR7tg3
+S2GX+QzTE87kHMhFXVlopKaR+sK0j3yEpg2dSSzWmAYCeoGGC1IO+Fhzidh1g16
7NHgPjXFkDwEUQxnIBVpRGqclXQtFXm1XN6dLb6OkupljkamNeBKOZPnoUWFU03f
ueioxwqgZAaqYsKaczPcSdh0/KcMdMdgOV3EmXRu+Kgk+vkM5fpfgWHP6SE5DIMz
2FMr3NwPiADQQ87gU7T+8iSAlAAFLFkUBxm1Ux2i0RrC9jxUIYw7r1gxAsoHitlZ
9/bYIItKL3FZxUEP0ryKTwkWBRhz7PAma1gyeT/06sohk6n30UEJ6xZJVrqld+gj
YnVwlgblXe63E9RPRJeGb5e3IBV/4Ohpodl1Snl3gr60t4f053PXa3aCblWJwZvZ
JqZOCVuCEIlbZVBMIYtez32+Qgqt3MXpky1czaqRlQOvpyE4nwT9xCWXTp4/th1T
PO8Sf0BWhQddwgiZoZAbXhPVCMMssv2XZOZUfXv3CCwaQuxZlzY/qcu/cBGImZLP
j6iPvyOn1PTdeSRQUSekbAnLey38jOhZhnD/H6sMaGOAQkYdf6UZtbFC5ZM2fws7
CsX24p6AfxHlS/sA25RwcSPjCT8jJFOf2xdQjKndBGqaylbyJ5qgTpCoMIEu+V7U
MoDM5rofnyYK2sV/teLEKZbfulLfY3lKOeSyzVARvwsNy5QqYVsDq6DLW4qqRbRT
scz0t/WEk+72rhr+Yp1XjQ8n3qUgrkQ38KZNDH1s+6lcmxYiia6O4TQehEc5Tlmx
CypOoNtF8n+LTVHEwyHhM5r1LVRFMDvJRve7eyOGNdzfjHb2FN1JhFtf6QHBF9jD
MemW/9oibCYAetDMKatRtbLyfBO+nUsNSYcYyTqpG42NefVljFKXjzlL7lBUqglV
Jm8svCF+lFftavMUtoNXlPR4KwaYgJ9c8XwQjJa1RDKDIL7sKeXlDI6pHUcXaybs
sq6WbOprEbPhxo6OsuU34TDmaTiwVtpNoWr+EiCWD35bfirRr6hYzrxGqDeLozAv
29KT/mq4sBe//+Qr9U4eok5Weloas8BI19dhGc9eVK766TgwbbhF2grbxS0lB12r
/c29lZ1M1SS7+Y9JwHz3CYdZKd0fCZbcw2r0ELuu8JudGAc0jKmVCSYxUxWfrC/o
kAVGEB9I0RZIF/kvNhmuy71jgnbE7RmBbd4oWV0rHB4vuOu8XSgk9hryy7dXSMNs
v2Asblg1qZVCut9ooIeD4Qm0HspZygBmgVNeBtL+pMAHrnyiDlvjdbTIDt/jG2ua
roOUm10UhqemJwjk76/+JNOBPIfT3E3c/ClU5UCmUIUTrGsCuKHdWQhOqKe3oIWr
iSqZFLOHj2yImgjDSNnNvzmPZwTFKneIhlkCG3KUWGgMnoG4eDwLTHP42b++4Dhl
ZiWUthp95MiQS2eoyzMVLUkZW40lKlgOwC1dOBVZ2Kd2aNL9ILB2UpbA7Fv08uPg
grpTIL2IchOU5fCQX+ZvIiSJQyljGUkUmZb+5coZ9slDZD1dV6/xIodhPh+ph0+S
Sji3Ipcp1Y1XOSHLk/eF9yyaaGx/Ja6R1TT/oOPqoD6P+4GhrsRMA/TCGgXA8jHL
knTrYFHIOG64bNCK8WI2roebVeQlg9cbs75MhFoP+ofZeAzDA7Oyefcgavwhq4Eg
w66gCfm7MmyEJ/eiVD+5PYgZgxUWj+mUAfc8ism7dtNl52VeCX9g81vbnDQr/Rkq
8kpBNumrWe9IJTH9ZSeyOV+vICUlZ74jtV4NESrRZQ7Kghc6UVIzYFjTNdejg0GR
EXG60ffp8RNsw3GLIHrVMLNNeGYB28/UOJLL7m/v6pDAulkU1BvN07tiorpx4XM2
/4T2EaixdUYN4O8K9GjcpbC6Ik/Rgapcw4LWRkuLRbtZrC1YmkEYoDELh1RApRyX
Qm2sEHfVD84cY1OVgVUv2ny0WkHnDWZIJR2a8z3w0+8XBieo/xHCC2LrtTw4NBt1
QjrRWoUTJWaE6fxDBsN+z4tTW/WwSP8P4fUlLRlIgL7SewHSlorfJA2xQmfTInIY
nD5PYCfXl/EE+mEt9ES2Vx/ayr/VL5dUIvw5+pN/sqP0/UjRdyUUYOJZe2Ovm1OS
LNfIt6g47zTjhRNy62Pk1oUci/AIFh6CucISdQNRUSr1RNKF9d6v5hhKSjHW1bDM
FTuSO4fuT7Rri109P4nDLR1Ww7gEOFM7KWVo8yb+U8WYXylElS2RtomdGhXvwwmc
uT5dvIle1bvEp6itzKOOERB3/BkKYEks+3bYsgWXoW9fll7ZTm3mv0POjrltfcji
tMWEmgHqtdHbTkGEsBtVunP/EQL35dDKw6+po83UTAAuPtdYKhaXjo/SSSQykDyf
FXFEO7blVdvJ+D8XTeVomxW26JtEFbl3TsVO2SFvA330GvYaDWxMo1JvSYNCuEZU
Xug7mlomADPo3T7ipAeypnC2Nl8CFznVpqPvvSLFPnkyOEDlB88VMp3koAghXyVx
H6Gj3kac/LHIxwJDbC50BuRWZJf4L5SyU68hu4maYP46UqDmcSAC/vFYG2TIJCvZ
74i2ckBiHEPU3ti054LjX5T/lO95ATi6jQ0NooAlrR1HY6xDzSFiIH5Xkpejn8lX
ZnyRQwVTj4TEMFf3Ilpx2YI3GgVzEXzZknWzKXNHFrM+oGpllzVY5fb8BW9S8Li5
caKTNIPyuHBuC8zZHO3d6SkW0q93/Qk25vbVUYMeqsRrozgWptgeNIq0xVF75Zln
UwWsYVOuWfZr80kSiIAq+aMPmbwsjuPEXU2tlqU6WL/dHRMuzUg4hBkOXUrt+fDL
hPKGWrXMIkIk5L0LbJpfXaBINq3H0a6QP+PgSANjYmV9ng534KjW/lSVW+JQz8A2
Fuzsnvv4NNUhuSehmC81IhjddnH+UzFBH4wkCJAkSjzMGlU8TadWw/9vlXnfcb14
KjN8Y53l630W4ACOm2mqpyQ0mPohkvG4vfR5YxiZI25+BfrnaFfNu5YpHfZbd1io
je0+2HhooLU6DsdoklI+UL0jlyn5HupTonPtTsJ3LnNDzNUIL6DIomMt1Xpa7iuH
s6+Mu7DujsGy1vfb6kk1TcjQTv9EPzuUYAckUJqc3B6RTPW7sQEaVDPFkoGERp9K
DNLGPeOIpbLUIAZKoPBCkONo2jyE6xqCxSvILuv/yp5JROQx/b3Eu3CnlxI6zNq8
baSWp98M6xnhxg00TsvSkmmdkn0iFHCqIrIpdMSTt2+a4T42LBz+AmMQYu0+SVR5
TAa3z8j78NqOgqgo7wQKAsVC4A3QIJuQ/VE8CKzY2tfKEwWHOo6MgDe4BfMIFMNo
dD4D2z1tpFuOLqE2uHIL8Wv+QXZOT8qSL7yvdsof6IQqdadKlmsqZrIXSfmry3Nw
mzYY7f6Mc8cUQzbO/kjBRWSVjtowXhlyqiVjizB7SZdrXPwkFlG+WrS5eAmK1oS6
doPIy4PLjK6OJFJJ73ikJ2tf6p52WR4Ddw83zrJ8+74sspsfEpuYfqNLvJQIOViR
F+eTNuHrvb9bZBWOWE3wzoj/BMkfR5g/7JZ8KooNZi21uQcLlYPYjy9LD0T6zb1k
E02X9aFKEM3bFsOmRrqlGB5y0Uf3Lp3DNligWZYpgBPBoki/lWkTzdb+Qy5A0VzF
K03HG0kYH5FxQVS+1W/dKG49ZxqIohpEZI4HBHInHM4c0iOJYlf6AZ5nwSUHq125
j9kFuNzhhVD8kpoJaizexeMUXmgppip4me8pZX3QClnwG9jtgEyrG48qe5l9CWuE
no+aRthAQe88IMzFF850C9q0ulET8/Q2RdNiAwhrcFrlW+V28KEC4T7Cxu6y/Fun
K8d2ob+kMYAOv6GPZplU1pAEYuCXbYkMZdrHLHrmBiyV7Tf2eIcf6NbAJFZIu9OW
j1OhBwa3Dh496vzghYdsKlq8XFStWmed6HNZySzAz9dUP9ABcn9p9KqQiOCcZqYJ
6JY1kuvuOcECrz8KJ9PwAAL7dpIrFyXFB/jxZUorDcIf8i+QBISImQWI7zO4ghRi
A9UsD5Tnd3JMhju4JmqWNndCdrPwXmGhpOWTJS8QX0ciGZeETTyzYZDnW3OTFBdR
w7IfqzGs1sfrQAT2kjSqQ0Bw+/cREnFQ18kKEiRvP5ulQ15wtftBfjUrDWdqDplY
g6oETASoF3qhfMW33EKOAehWfa5eUFtZeK7oPOhP1nrtP6p4Q+ZOpyRbt5T1bpgO
GFPoUujxah9kuRSSdluR2b3tQKAGnDZTn9xuYPoEB8yQnTYlrJoYjhnKpbOkLn9q
ZLcCbE8NrVGh9YS7bEdjeqsRLx6CkOUE1Fq7NpUWMJ0Bvfaj1H5E+2XFeoOgDnPn
+ep6aTWrPst6rctqYsWRuiDGuTVWd6+p7XnTkj/LLponpohDg2KmRdKs+HgZUUUU
1nt3drqZaLx34fiUcJlJfJ1T8LdGldCEzxsjSxieseZsJUyO23WklK7ldOBT7SrI
Pz1x6VHUXGCFG0RHXz49tl1dpimMMoI8rXAo9YpAuA30XpnhQAxPME7e86T2JZr1
8w+W2WEa9m40PWKm4iiC/fzM1yQ22P6YxaMpxQBezblNfqKGxKFDDAbSp5we1jao
ZkUYPp9LIBRtB8i2C2+s07ZC1iMYt5z3PLkso4kSUdAX107tYRFV91KlfSEgVmk+
kOvZ/5AFHYVHVvja2PhOFhtsZ2h3NLOGSZXUyNfg/qoqDUOgupTBIS+3/AXCbBja
SxMxRqTXa03omvjyCelyS7kOE6AI9Hk/fghbfg+Y2TxTc4JnNuex2Sq/9XQdUrsH
6hw6L2zbdmHw/5fpfxri5GJ2PmwTkQOcWTK1tl6pzzXeMxuCPIm5KncozlCrlpBD
+Cn7CnhAS7BmidnZ9CgELryVPh1i6iSk931Wuj6O+T1s4AfsXK3H05bPovT60T8e
ehFtFhKksP4ztKScn60fcXPONzd1YgYp5mCYJPyMkr8LPS6uqu66WZopKmeTrHCS
a3QiyrTvkOndoJXeF6goxnkhv6p81GCUin7w5wxpsu6NM0+MyoGk1i0OEBYKEC+z
h9SVuD5x+kKfY/vUARV3UOH2SI2Z9K0CXXR7PavW7Ur5NKVqj0Ry41J+f67Jy84E
TW37yYlkg7pbpYoR4iOViO2PbaVcxOedA2wi6wiOzemGv6xv/l+4VJYmRoJ/Oawg
6eCn71q7f7M0pUQHMAdE52b7Dq5iHE2+TjwXmvdc/S4Ml9TnsVWiQYhZZIBIxBsc
SaDupEUNjuTv61rAoGAGV21YD80/7N5YeDmjXmzbgpNTUNPwGveFtkT5fixd/n9Q
I2q1aX2K/+u7n/TSmjYn86Sl7Fenxk2TED74cb8rRSKI9bmwWKfhXooe6/k+HDg7
2FJA+maOdpBu1RQ4g2I23tG/cweOPYncpXd+qXlwCz+F6NRxZd0iYDlmrmmTqZ2P
RnPidm7HMkoaRWiDlqPQmGgJGkSscbW6vF6ApvymFv8A+efuNWQJABfOBN/aky+K
AM5VqLjAUR2wOY+78qH9FakW+efGH4OBMV9mEGLOl2L1ETwAM0rnTjtP0j/3JY6z
+6m02aBsHvBqJXbTuX2xKFjqIA64Oig1QxX+BhYy3AcPvtk8rVNXBOSMd+pOAeWG
IlQsiWAqYPcUG7ekdJd0TLlI1LwGFyJfAV9flzgQOwfqO+x/5ZuxxQgEM3dc+GbQ
gcYlgOFBuYHSqr+BMaJG1f57SFW8ufTkLCQqb7ovDtHXnICTCkI5aZd6oEHXtg7N
X8az6iIqWQjHrIpz3/7d8rEY23w78AuwUJBeMv5uePZri2/fzqMo93e+2Mm6A6mN
SyOXH58oQyCmr6yQz85t35ciM6ZVC3enZmfGAOrEGC/SKQk4eaAw5ulhRQRJ0HJM
SkLHb+tMuf8N5b0rK0yl7s+34figrrq2Zm9lHfD9XPlaO9PxVjDSFGHJ1gQxVG7y
2HOH07Em8drvgh0PUgEbPznZhMZ08ApjDsUO8sN4haNQ9wcpDYX4tbjIiRRwFwQy
qfTxfEmetWSOjiZCCuH3R0gPgmpHVyOO/QXOmNK2B4fSAJD9MBY3NxAwKL58aYsK
SGKNvmVLUsK3P9FDmcxkpTUUn3IrQnfOGmEUd4bLZAuegf6DAEfCDJxjcFoqh4US
fMCKHQnXlPruI5CnpgbimskKmxhTlWL7L9Dgdq1Sjy5fC+bd7uDk1Idz+lbl477M
aOme72QR0fFXbxGdbOLWykcB7hmwjgTr0hipWw/ly8NmSRk7bgAXHo5fC2hxGF0m
UtP62wB2+lF9duJkMKleCBB/225GeLllUPiCN37GnUKZkdQj057jEQfQNlCfW0G3
dEqNVBtobW8ME8C06U36irpZljVTarvItw/mX5IVDckE4Ip4cH5LUEoSrfregGn0
JsFwDBJmO6L/MKT+0wccsOJWeganAshhN+yRsIWDWvHeCJRaK5DIIQkPogSoDoSC
5jKBUIVo/ApoSJBzqEv3tETEZo8M6uTsaKkD7Ql1H37foR5z2GkCj7Jz/iYJcPD2
FjuvjQG+RkJy82XbbzHYTDdoaayXCFDftR+7Y7tgNBzuWWKLk/6KTYRcRnjmyC3u
MFzeNaxrz69YfELQv1+L+DAS82syiUQr7EiyUFCKMvU9AaQdmiFlvqv9XyrDYp3q
MPb0a7BZC45+idUyqNcY9XEIaLgIXSIOuGEygInCtZjCrsCM+A65XhG+xLKoDXJC
yVkbl3TThxwUxZBYBmlbrMu8Gn9jdvlp1lnJhc/nHK+8ZTENILm3fK9xfIsAWPLe
kCOKxnRz7DTijzxggklSq6MafgUduLdrIuXu5ybs0i486PR58iFFYrBpsY7QnVkR
ouqcqXeTZOn4kbSnr7yCbD2HycuoGh/0geOnxxt6rIJY87tzCbkSNabfdCCuykua
tH2T1wW+eqJtn+8JsIkTLuJiCLtfFYow7q0gQQ8MVbmHM6hz9oP0Bc4MOq1wKhde
B1Y70d89m2MMqs4pyAyc4tYH403Q1iIEISC464nvM+0SREEoWAdQVEGnEQ3fFdQk
EY4F/ue4AIeX+Qq1iSspuifExofVSkXJUI8spe5iQjrSLIUJBr9vxxioLGQc2tvu
udpAcofRK5QuaK+m+7DnUZmpHOvgnQOz7Br7rEN01IbM5JUpreQuNInbdgu+hH4f
gIB/XZrBcL03JMQy+efFCEsguerLSjoP3i0VFUXz5kwS9tBoF7xnI425Rv57VT5h
w0cGoPAKfq8LoCLySidynLTiiVo4j2Bw/gBBuCrBwEet+OAiDgtsQQ8N/T9Y0Sn6
NuNeuGpN0IMLGCI2zt/pjtbEZO8ijgaCPTMjqvYHmNTwPJWHPz84ogiMX5z4RXzF
ytdmlbbfUfVcXYgyOkzhlq8GG+gtvf+4OqaZmv7sAtyojfGQyJ4ZpWimlhuGibn4
/lqGOCQOimTIaDq9Hekgl6BfSKq9+U44BrU2nNcmOpkqgN2bq89acAa4tNKnsQoc
9Rx4PvoWqvOKtpigHdVWaeC6l/tKQqGgeB7XNudM4inmaHYYttfmCnbMygYu6S40
Aiw8ZQA9YBqOFJVXbebZEDxzxfDVR/Yls4xNnrPG5joF4PwuRerFUWf5bf9bnqvN
FUoGs1ReSQjbPE+W25Fbb0j0oDn9rO6851EefWuwWwBXT46VwzPEyv+0HQ0lrm8y
KWuu1VUH+i4ecErYKPX+WQMzGQUSFV2yj3zk1seKwT8rPkXH61sbDM9WsWHtFwmH
bU2x4PXRvfux/wDzXOimrzJ+25KYTZbANtszcPoc3THUE6svjFsV0PaObPdyUSM6
IuVqvc23UcGp/B2rF4L/TWRXNIVL8KO4H88R0VQUbBykiXsr2AxR9XdXu9UfoJUb
kK5aF+J+vJxA9/23OiAZ6eejuft3E5wDP5HxxS12rscTayAmxRIo7DIh/WAE8Fcr
Z24a2l6cb95RCKvN3gU5UxzBQGvW1tmp93P0qnYlPAK2iQjy7xZn+0SCiesgjIf4
1opW+ckH6+725dx+1N4U8CCceA7P7ruYPuiajSDF/W7kWtBKvfB5jJltY9IpuGCH
UPZx0g32qGTWHAx8Ipj55aI/tDq6qKMFIsOPpyuAqNT5k5cikcwe+yp57EQ8F1YY
QdJ1szmI4pdg1bK7MlVPGP3M7slX0mdmi8Iy3hjxbOPTI8q9fkzl2z1PmRJUkKlh
HTw2hpIsvsukKdyvRXef6aYYZYN/EX93T7I+kyH/fep3Los+zkgmfj8yUDNq3XJK
y3AageUmcwee+6KS/QN7/FTBsGqgB2JoQfLRvlU5jSxpZm3vY57pm9fYA53JdwnF
Cfxrgf6md6lGm6V2G0iQWycyb8W65G3iZ7el8GZqEjrmX3hg7BcAtGoDgjHAUAIz
vVlObreSB954e746NXwY8jPZzRzudflWZqJnSz3m2DJ4n8J339q5oLl/2Bnutaui
DAQc+Ku62rWvbjmtWYLDYvYlGZtWTdJximaXXO/CJvSS/AGdmTwEhpoiQojaA9qD
vYNEZy6t5Dh0w+NyXV0VlB3KQ1/odqJNG+KimWzbxoi89tSbaRm3nf0IWDHBzsmt
UoxNEBq5zDDwUBKF+p8/u2ComfoPtrEVegVJxNGunAqqr8trEagWhx+AqATUpgcz
hEktz8z5jmTFno+5TP/qSDoS5Grg9cuBSA7n/cIZDLZtKO7qPGD91K6nZcfefIJz
yPkQNjTRfsQw79Ws78udjPznFmgyGluJgHBpe9ffx0ZoT+X23TPaaHu7l1v5QrMr
2Ih/ErgLr5mgoWB4MNn51mJedZXME/9up45IY3QjZEJgFR/4IIMBvEq1F1gKVkYC
hnl3KkTqtJ1tonFPuMgj0854sT3Yl2uLBMVVlDW30Ij9/HWUYVPO5adhOlJWxN3l
ygVXtGFO1JJqRBxRxsduSwLqa9FV8QkkT8vP8bXBCy5KtrnOCbpHmgcg1UuWRt5S
B7N0lH+5Edu5ufw7b1xTB1rhkJzRpyYuk6PYsU4qjYO1wJtX4QLjAG5geKWHU/gR
f+V7fDNSGGUNMeQ23ONgMdpAweiCk5/fKmSuEVC7CQME4dzPH78S1C0ks8gptvqa
obd2PUKeCAfHfdQ12wGVrmHDBvjFfC4uU5w+c7tYpjj0GWPMMIhLVDHHuY/+icOV
5NU+C/75Q1+Pl/mUpmL8NwgcTBPipoFL7NLHvP5PClhQfXRu3hytl1Ad9rlN13J4
EzRSBajuyJq56NTNHnuV0kHtdL5iZK/B/C/rtCRlLhdzuxaUHRmvAZ4KUOewst4g
teOWKylyFaTURzLnWolTFlAmjWu6nIyfVMesBW+KceY/2cNl+sTA2KiWcmc45mvb
cMoobXD8UJhhdg3bKHRJMINWTwLnWeAmMvk+Kg+vUgdSmXguGSbJrhj+mnFX8Y0m
SrxLg3Mq3/tJ06v2mjyVwuBb5MgYWOhFY0uOF3fiydkt/oflpVzoxNVy/lOgaeOv
gtMxSIEJWZ9ePLTetmHxFzzF0x6wPi6l6FeQdSRafY0uSHWln5y7jppgRaNpxYnQ
CncQHRu2OnSuZKBwjCzBs0zC+cBBaohbfZpzf2SFgV4ZixyZknioDsZF1jv/+3GD
Ph1M8E/6K32a8j+6A+hp0+p8sZdH/yklI7G7FBUKVYYnuZxEhX2anAKPKFw5bPhQ
katGoKdxQN2XJGMXDMAvmXq01fns9twjBxcHm5OzxwNhejUv5QZYpO2hJZ2REkPo
Bp03e12Nt5dzvBjCxzroc6I2wcmRZIyk1AQ7VotTMb3cVp2sdjGnPGLCEGXm0Kr2
JSGxZSCCiRY7UgFPpxCAJIRDFb521AFIEMGA1Jy92nacx0oExy+GL/gfDZiZJCPV
ypvYBMTLUj6Uh//SPK3pRDgvx6TMzRk0rxka/IDOjMW7rOrHB9vWnWFrA8kiWPWP
aGjObfvGZ5t9KBKIqk0+vRIQ8jGcMhhXmCLvnmsI9Wuom1CQGORoswMCVj6QKuwX
ptpKxhprmYRBfJ7SUf2JS05d2MbO5o7H/Sc2c6b6tvQ7GNiY6pvbtEwC1KFx6yNc
2TxnkB+Q3vKInblsXVaYDMbnmyKAiu9GtnxeO5nqDxcO3lnQHHYe6TXrzmeMVLk8
mUxcRsqVU1M2y7cCjUHL+stglyJuV1sU6QPjALkbZA0LSh2ah3J9e5VcR4OQc60o
J19NWTPbzSWpvnElrz4K1yfrVXXuOaeGQvHnZmM1mBO+BG9qae/zmBJlqKkOzlOt
YAaRh4au/ysdNpB/HMEyzJZV5xurxzEIwoRSGtGItTYHClDQW+s0TPQ/A5C80f58
WHxagRAfwKwBwRh+xM4EqunnPnHGPCKvnbzcl2dLOmtheNCvUf4K+Aj6scisp6w2
b1LnCX0edsoq+G+jnt8G2Z40W7Db34vBBDZtDm0AhrW9hWN4rpAo4zEm0vrqPcNG
PcBIWSfpb5Peew+QUiGPDj4B0YCz1ui3IhY15DnJXI7bIYjAOhsg2Phf7DQPDmM9
EaRiWpqifZ6g6WJlsPyOt75nY2Kc4FgSV3rYHCuBbL9jiaXiF430y3VIqOd6iCTJ
RmOaDvM1/nL2gJJMVXPziqfSigqF2ZTkx2nuLzdoMqE0qMp4R3wITDeeMQRnEWwI
NZE0GxXQTTPblvxnBK0VzBHc5cP2dN5KKgRVRW0eJd665o98fIpPDfzuUcNzpzfz
o46OWVyCFnneTccjjfHKGgOsEmttECpQxko+Utr7bS//61FYBrFKTR1/BmXi0Y/P
V61uz5gds1RPA0RDqOifr406tLlMbIF0KocJ4bsKBwc1bC2h9HDVjDn8HqAEVgBB
+0W8/dLaySdvlFXSWPJvVC9vsktUFmPcncIq41m45u5Xpvn5qYAJZkQt/RDRLttT
Vo3nCtsbyH4ULf3sdXy8EFYfw/8aWolwhiHkVFeihJN62ipAC0rCQC0C5s0lcXka
UtVkiXMscY76ewJnryL9lIx86OHeq45sa71QPVeqDf6AVRjPXKvvVvc0CD6g/HEN
NGyDHKDQP6rQ/Tcni8CU2geCYI8FwCMui7L9iCW1L6z5dV8G/O5utiwLDSaTteum
fz9uG2Fw4mEVnZStpC4nhXXp4+pVFidLi3x2t0NcROWfifxON5njQO0LNMEHWF6t
Gkoy3buOW4/kAzEEF/3SpxRsWu+bV6CIRuzpqM4+MlzUkAqdUuolE4XWrNSyWmzK
RfPFy/r9riOyIVksKmFAgwsoiz45xrS+p8mLabakSxPTlricEWsQ+Cq9mXC6D3xF
SmKtECaiFZ5DXoxr/6ahXBLAaJtayc60DMvKj9JIQ25cqT/XB0oYTOYF72cH9nmq
e+3NklzwtO4tIbA7LRoFjG7gPibPsMfbl8Zjh/oKXkkmKPBQyL2Y+4TH/TRDbodW
ozIUuFz+ob3Mqlncsh43voir6DZruyO1Vlfee/HDeCKfyEubn+huM33yLiyrhof5
53i2z2FVgyDcrZz2SwQlUfrLf3xs19ec5LWBkwp/R17ldRWw+Lljl65pCaVfhd6b
UPgEtnu3drQdCRv8IH5CcbPU+lFqUwCQRasMmrH2Caq3ndvI7KP0KNm58DIAEME3
ahC9do9xnw69aqu5Ee6oNVHsUsWR3yAUhPIhy9n0hyE9XzNQPyLD0uXxFQ9MaLtF
CHY20TEhRaJHi2mHdvNZ2adN3USSB3Yny3As3Cc6z/WuOBBlZz6PJTKKZgi97Wrf
dNn5ZTb2JjK07Oq3PiLRQ1i2rr6OH2yOxrd9q5wgZPmw+4xeoOf482cnmhxJAxUf
1r1VWyW+T15R8ZjowR3tM2M8CQTJkZcq+rntlDxbBFaTN8vnRl97zAlfgUZxFTmH
fGVKQkWJkv3Ra2hX/1VeAmyp6sGrXRm6+B8kMEOlu6BDqrvuRUDb5IgBLV2rSnzI
tbP9+AoLaGJCoPi2rCuig59d1r4aNveDME4okQuWJ/rSOtPKOM8fSX3bBirpZgGG
f4R2UldKu5nGK0ZD3HA1BjIuo3GHyf85c7tP7si6zB669qaelY1kE0zFzlv8dIn2
UvP/cw9IVC+heR0mkD5HvjLBQhl0716ngVeS2xZVP2FdxE+Y0apnbakUF3W4GELb
WQ/Mklm2Ce3FJVqQO/nGuco8TLLAqiQSvc8fHkm6+TYNUh7sDVgvQYH4GsaYVJk2
YYBKo0Opi25ZHxI7+GT2kaqO6ap7w/pHJW/JznOfNv9HmXBUBZ9Zg0C9LY5Sv/Qi
pkCt4M6wft+gIyGTcNN0ENVqPM+2N5uHiFFLBsU65ZOFagjrOv9WQWBXKP7QubLC
9Qi1NXBqv3l+8DaR9K1giTidNmeGcRpbGPH35afu9/i4/a5nUoRTaif7vS9olLcH
rJP4Vxd4FwCThvbzB1wuszCl66DtxMeTnOs+xoYBaJuLELvXZKZ4qQxdEYHaZ0NA
JGq+pUbI6BY829EqI4H4FEE2JqIKl+kLAW2a7tGd2lAKK+/pG7QXo9lLr9Cp19F7
V1zoWXdzcVpyjxf624zWvDuTtnmYBmrmjlJUhADOkFSMOBxTPVSIoZ6qi03j1NoT
VaV6R+VU90dmEUbgi20Yt7mw2laMt5yRXPCm29N/4xWurGDbfe/4O8e6EhmDst8k
EuaGG27YjUDwO43mZfHa53PQBAv8D8IZbuaggQsnR52MExK29fb5/1nGyRQ9c14d
QjiyqT5smnALNSsReFiFKu6S9kjKAjBqoUgAhl2Al7uDkKethAIBLvGtJecJOfNq
qd2rjjNMQlhrVWgBtECGF2Ug4Q/sRZ1GwW5aMMtou05g4zSiyUiDVSOUYqWliq5B
QLcxRnZ2W24PUQgYFa2C2ocJDOtVN0rTyR9THbLv86t1wWel+Cjjdui8mhxrVCna
IY0ZEw5tyNQWcy/+vsl/pODBmlrib1LbnigH8vWFr+KtOWCZsuMaFz9gjt7CvARw
f4IYhADnlu/mBCv6mKu6sjzVGIKU/SdxebEXVA4d1KVD6K6cxuIH0xUKz27pnZDK
MY//beg7l/x9VwD6jhBxmZapduXwSiU8WtmRkz0R+22o+3G5oN+XiybeqQxqEGzI
5lxxIu8o0aBH01KjhCFJGRIH5IA53xpXo/GDRCzheLuOyaR7hV1rlFM8T1vPcCYA
JjgnRP97aJFO89GaZ4ASJ9uJGBhhIeOSHhxbaSyH1Mzs4CJ73hpT3qmrGxqLolZ/
6FJQrHxlRZV7ah7oEN92tbisVkbBWXE3wzyF50EIbuWlXy2irCCjFz5sSfa1LEYb
RupL2Wz02fcFUXz9JziAKnPBT0Pw+7BY+ACxZAwYq9xDvv6P+IzWR+21LnokqL8v
5ALY/db/vUrWNoLuSz5uDWVShX6yqGKB82zelPrFcEr4zTGxdMn+j02n4h68reEK
JRJMAEHySYCiWkKHdTWNfJnfNYnBfDfpecSyYUWuZXuVtcatBWvH+K6olfHZm4IU
a0D0aHAi/ZHAg7tW+E+5E2DbGzixAe0ljGHxN6JXpVVZqg9gYoPMN+huqRK/C2n5
Lv8/S2YiZyySN3Kk3KErzEaUk0ls2ln3NXXfC4sYDav3iHb5rRFki3MS6xNetUwD
ct4us8hdWBk+uUKx4VSxGzBxVRdZVlraZ3J3etrrMxfLOvyvzAkqX7vl9phViNHj
KriRR52qFQXd3NqJuxS+cI0HTLK8jVrMjeZVm6oNXcTBHFhDgiKCGc6i7R05FJJi
LDSF3MKQCwxFaWpvV/fvzmeQCXPy4nefRRvY8QoaP+1MBYXadtq1kpfD1xR3zkiB
rB7C14Nz8AJK9cTnk5jZ0v7h6JLMlHBjZ0iXgXTu0bwmkLjam5vxRXG80HQ1nwPN
K8+WfuJq/Wiv63dCGkSwi1mzHA8xUaEoYdcwnTcE2YXMNb9RiQ4wruC8pWzAPjXS
dji+mhnEsQE5zbDjXvWN2DKOnnwclxycsOzzWU9IJh5g0j5d6Y9y77VdKWPnesP5
sSYIBtrn18bU7i2HshXxwb0O3cfO6gHe9AxKFcTYvcRGiDfVk4spNQ7QgjWHscou
pVNM3F4ybsTAQXEcWma2OsfyRtAq3WPMWDMImCkWbpdXfu6GdNH9o7/flEPXuPNm
mA1qg73Qfw2t/2XjSUHnej83RBul7LdBs5Nu8+pYsjtXP22Ze1mMcPJ3tjuHl4i+
b+Lt6klY45J/hufCnyfz4D/DJjcQUd10kT4u6TVFMidH0afYh/5WXHnLzq3FikcZ
RiKObedQ+SjU/9l6Yoe4CszK9+Svv+ByUMoUWenG4K6Dd8h0+U4h4i3nsNlKoeBS
VDDY6rFBY3wSEFYBTdmfX2bt8vm7y9SIoZR78GKD5QWXYOfCVeAHYBDM1xnMCBWw
ZcdCyRAkuX2EIyux0RO76I1ILyYEDGR5XfGeuGPyjFMz+OSxbX+A0bzPcTNC6h05
s5Z2FOrOU8c9/YrObLpSA0DiQMFsXbSdKh0xZXV6B+FJ/kRdjwVS64KcN8HUM3SR
SStNGg+TyqV7Qe/0AcN4zJJVigxUTnWSzwXMXlaM2wDer+neXz+UXYA6t7QZOIpO
CuKL8h160hWQfjz/0JUSrLUsqk3k1CLfD2azOMbZs1Mru6q0NdjjqwbnHyGvzRVs
fpL+3cnf5bm1lQeZGxO5bOoz8mt/GmevJVKiGxNml3cS0hD7ZuCwkMtQfQG/KFUo
0h1bjPYb8Q2Ck1ls1KxpM2m3C7lO30HDjrYKMJR0pqQiIWqThBaUnQqphjNfUC6K
Nd5N80AdxnrWgANAwJpWA7Etv02TYL/rVgRQ+MWM11nSViDKJfLnK9Fjkj7IP0yn
suamcIfeyOnnl/48xe3s072+S3troqVmAzdhP0JxJWiOnHoQFk4BY2vcD5w28n9z
BYRg1GAbr31t+NqziQtS23YbPMFvaUp3EuRVo3TVQTUoVO2maFKfd3gKGyhz3Ssx
6SJAiS2RSaLHy7I3gkWNMJ1RtDoFMTPv67h8RS4XCLm+Bh+XtzWRKXZy8dxdri+b
X8Zoleomoz99q4wYsCnCt6oGaBkuEM2kyb38R71LoyDq9IgXNfJHaSXQAMrKwPNB
4yQHJwMipTNLactZnhQV/lih4Z2BW2epqPwFNa0nRGYtWe29A2er9TjsTXOsSDSc
EmLl2j6SIoi9tjofuTZbo+NvLv09IQDGIQJFRkWSXgfW6L7YnPK5f0wRDaXP9Uso
131BscbHpAzWExsbwll9NlIpas+8krPjw85N5vRBJZkfkYJV8nXBInBfHN4OOXlJ
k+3CN6d2BvxikNEdySiuQcsX1mLYMFlo/gt0/rKlDBwdaVwiuriFqdoxqZfGch31
XWQpFVoMNoQ3HwgnWd0WPtElfoJXcFIRB06gw3OagGRBx0jnDSvtY4nANV3dUiFi
dzvE5BaU+iURc09F3z2QXBU4PPHSn+Dcj/ue1wH9BueqqwjT259DyD8UmfeaOJYI
4epNapRptGfdY/pIINnbyOYge423v9DqWoS7PR0e1DD0m2BFQ3NjZTxlMa4qd170
hZnGovznkxzg9Lb3gf+JIlNwYu+hSgWNTgpDTBTbSLf6L1QtEkVys/XjYtmxTjSW
TGevjkiw9IHf5rDRCHs9QoYwPG4UZZicq+3UFkkVLit5RBEoOcUL5F4rL+G7XFvd
d7nxaPhrADwxByniZQtOf+sPlqDkN2qjg2y9tR0DfnPWoCSM3itr20vQxwGJ2GYG
SpXK2wpdc8Z1Yv7E8EpVoUxWeyoAYLnQc9Ma9hpGabbLqtfKeX15ScLghny4dum5
MejEPgKB5hGCKTAzJrbfOpJ2mNVPKy6w8Avd0OxK8HUBJB4Q2zO15+heu8yige++
Jed0AlLGIiXvsyJXY9vzzd6PXF/ht1GDvSwIW9D50LP8849AcISLrcAud/TJ5NMv
BbZ5xg9o9uPNaodSzXr7fAjkWo12RuRSsatMb4hu1NN39RAWRkmodpDGvRt4Ik0y
S4czBEO2fjDN8RxkcIThSKgqL1m4po7XAiuOcg2WykQThmUDescrG1Qbac91G1yJ
ar0FtTOSRCmzn3kLtXLZpTVBujFyDy1pPrtPB5s2RKbarNMWM8Pe9YjsMKk22Xl9
lQdjwqCx7OZYwzlcKq5inhEPvgzQSMfROi4SMc/Wmb0AxuYvKhgnL/KYug2bawFc
RBXlR1mcg+ZBNFUbtgNnB5y9tehnkpg7N6l2WGH2rYOUo46lAzypfk2ftkq5G+fn
2uQSK7EybHD+iCN2VzA+zigmoFLSK33ZdlWs/kx9k/4oeQT4l2glub0eTpQ5VYQp
0o7v6cJ25p4wq8vCbpnXcwBQdi9c/mne++F5kX91r6UqjbUQP7tgkfycWmVu1ZXu
fRxhrGF1vkVHq6T12iGdnHC/uxpflg5uI7JK8/W1ei5T8TkopNr8mSq/+lAjsp3P
7jkJBDDNIyyoo04cO70QmYNQycUO6BzxXReY32jXNFPuNAAaEuRn2qu6RVDaQuaw
u1dxHYKAFttYIMrrh62BhkF3h+yPvTG3ybHh5/fctTOuwXBGdEOgb1kMPMAO8rMB
Dg/hCUpVHlqDtgc8PhqKflD2SRFkMepiU9rALD4OiW5M82MQlo+hAJ0IFKBrHzXw
+xFkaElicuN6vIU7i2bi4rCSXb3YnEpDwqE0UWZcRpybGDt6ltyu3Zj4GGt4UZ5F
iH7h1kbNK1Ghur1Mz2APAajfWZsGfueqsqgPpJYf62QRLzk2Vyv2no2D2ZP1aS1W
b1MrJqXU9XRKyG1zqKr3wFlznLvyD1Pg5TCGSgnWUzyWwP80LOamt7W48GLiHDnz
fObeB7d+OEjQN3vXSfM68a+J3L8tDt1jvJ4G1KeA2ee3CiU7GhbdDXVE2dg7oHN0
tksdYOVL+5MYMLBD6yWUlR1jOvCZzj1Bima10/aGwbmDw/8+e+dgXo5ZQg2/3pZB
4ebyP0Qu/iN6MpgU4nMf/sp2cqKZD9yVk0x13Pllnqe5OGoTh7lfmwBCAJFuVjsv
e6WEUAciVi8m5aZD7wLdJpCq3GSZSSgH45w2RE32hNMf8UbyJOKn+hJPILE7mcJW
lxqyYbXrWBF4hvH9Q5RSwHElzudCQymq69xFZiLtlB1exrNaJvr/ZhA+y8qKkEev
ZyirpQpkcyZK8gAxyBXeSD+M0PTweU4WX4wPxIfFue6PS2T34HpD1v/TKsoU49sD
U3LuytyRjHJLeVb2K4zU8spUPTBUg6mE0iHucNzGR0pONjlbvr6oryzqvv8WvFsH
Dd1c+YyJK0tlZT7rRkBJdst8GNk2NGxMYUBZ7/GoM+C0KA/RykjEzEzg3ZOXHJuQ
TNOu3N9iG+ee/yLcz1i2vF6WvMi2Y/v7tN+nvxUjkM2J7pnAN5F/GI7ydX1XpF7p
dWhPY1sLeBQTsWQ8SKRM2Ig41QtWRc4Xh8rb0IjDmtKC6x7P2W/1eHX7TmudWrsl
eY+t7i8k9iUYmVeTjhlLAlm/13Fzg7tIDzPdDhV+A9QAKWibmoSTcwn/u1LFa9kK
FG0r9yAbcKAKqYckFR8Ks3lqsSTZ5NGWpUojd8xo/wXH+cMwZNzw/PK/5//12YmC
NpJDGr2zeNFh+Rw4c4FCUxuDNOg6Rd9hZy0NITte5sIWCVvF0U63EUWJ5EjL0Frw
rqTz6mtK2v2Kzpwr5BQbi7D5YnFb1n4I5LM7mag4l6CCaNHbL4yt3FPcF2MznSdy
eLxM2H+AumjTLy9HVP+Q/mZomGfdWxffyAIsFCryigBLTmay3BRDqLTbXMEz19R+
cuDFgrc00GeahfKY7usXbcOMSD1S4QLf1uGtaocdUq1ceX+zT5tyfTwfosnkIvwP
QbENOVp09/pjnPhzXJiZAD8bjAf7Q74NS2eaGfgwowOoI4leEd7mHJoftIj6I+sM
nrA9nvUy399K8o5aOvSLT0mRswqpkRQ0/jZ+5HOH53xwU67ZHu+QC25S+v3n3OFm
0uCK03V6loDz+pFvfkCtT46aoxip1Cr6UoQMpt5h4P4NmKh+3irKOvkna1iiIPIo
V1z1Lcw4jD9WxUjvlBAtHNo98Ef6aexTeyUprCubqnrvsjzL2/bicOkd/D+0w+Wv
aYCTmlD9fYmz01VHQ8CLudaF3ElWIZRe/AdZYy6MsrOQmkqMsMIMsRaPxKliMjfL
stkzxLkuhmuFZgpOg9waCyBHDmVqBrT80GZRTLsZ9BXBVl+KufBlh8iwX7i1fgqq
weVCqTBvqMWuGh0DcIxfC3Adxz3TpdDnF4dWuhMm3GxWErQB/q0EXhx33PXaBsnG
kPtwZ93yW0awed6G10O+GdRDc1TYXUlxorae1oAFnTBnOH4TIZ//6MjgkhHwauCn
6C9HIxlKL8gzY/2XuvCdV1yEKfZvuDFHyPdXiMM7XB4RTUd+gRc9/X5hJMUU195V
nVOQNzvm1uvP+f3ITuvaIuEzhOdaO9qcSGATnEqnyP3BZEzqWeZqYRZvMVwk0KKz
BbO4SU07g3CGRRFrQCksLFN+t8U6m1vZllUvDLk/jfanpmsAsPwQymQ3p8KCka8N
+ZbNJBSuetyy6ITs+jpYX9kU3wCTP5Qs5VLeLERQLbu69obvDinKEY+sgBr3xWM+
oBlspwupoG0vAuIS3VCS+Z93AcOi+EPUtVSpYSuvUuoo/uojWDoPEqjjpd/J+p1e
vZMckSkgdNRmsvrvqlOTaSiQUBTPgw6X1W1SwH6G4YAdMjBEdYqB2SGm4OoVXZ9f
1ls2Emg201+ByPL4C8EMl3vJCBkvvYxrh/ewVdjXY6kw9H+vpyypC74j76EjWVN1
pr/0KMEmIZqcVvy3IcCcZCR/9BcH2istABWhYG8iVaRJwTxqND6U+A/KMdUAF8sF
+X0vwVE1+Cruec9F+JHH/vbnQ88C0+I7FxbqTUSpc6pUETtj87/Lk7tnNBNrSgum
W5ZGJDHIJiip1oJxiPJmm7q2TZeCzCnYmkC7v80GwoFTgoaz1SluTmib7BGc0L4v
l1kpP0SmESxqFcf41+FeyMWEuhvpmQFaQVF+LPBnfF2lr1uO8Zuyl8gbl0ef+0LI
QhhkZ12Zghl5Gdebf368ru6590jKYTWoyfAPrvK9ruO9/0zWKQa5yWfR4tV+VuV+
4E0otknmihdbCvKPYTEbzv+sD1wYLx8LG3ImLzfi0WH0f0GUN1dak201x1LQk0vq
qJpnY/k2LrJF+8ag3oH2z8wrNlAwiGkrfc3EKvMayv2jhjcFoR52ZcnAhxhSACoH
+6rzCvP5UW6UNJujJ+XL0z093Znk43Cz5ZUx++YDf1n8aJdMoy9zQGX8HE/ZALSU
jARVSFpAveQM5huJcAlENrSjxM01+5ykHAdzeTfn34zBH1iyUA06KQ116EWdi4YC
vQTbjOk+/hPslTmN7JFCPuCPr1KTx1LhVSE0JsXIOMmH1lcIMAH8PthLH6GJjh4E
mpuo8BsDHq7FRJYDvRxcnDm8vJ+GTraJ5xsyOJ1IjD0yzYSX2MDXRwn2bXBbI0gX
YCP8c6sAtmL7PO6/OkWz+ZACO5mfCBeeX9TgYMqyn94ncropuRhkWqpAnNSSYaJh
wWp+ENEsFFibJtMv25T29zsnhUGb3CmbDKBcksCqtwA+lpC0gsGFfTo6c/Vs3/cc
x6vT33Wh69ZC1oXX0KfuzdxvnpD7CLC96BRCDUyaxhn2NKJLBIIaX3GBu9TmzEG4
iOCHmMKWL0TEcFNFRDMoJ+QdiLeSy0U1yJ82Bt1IzJeN9qnfAZce84tp3RlRLQro
Yov/mrshmiYLwQODVC140xjLgES6lOFIhK0ibkN47xbDOZbg8BhzKLV/0OSxFHcj
6szbFR1Nyy+drPGhXXz4cq6IcFpTGhHGy2CNZsUm7o7nTxDrHnBL9Tpx260dF5hy
TmNtwcvQt8kzCSQLJsh7+T8jAr7PLkM0rbhJFCDqTMimlrSdPsa6fpxt0Q23Xx1y
DpoIzqsFYsFrDeClLebJgM8LIgyyT1L3eEYdiQo5W399gyuizdWkkYQUHWfo5+6g
VLIgtfzjFRTcoekQqpwcqysYkjoE0t34jv5E9xpjZw2AEUT6LYlvt5ePcnNYTaya
AY4+43jfYtMW41Smudm8T/aOyu9+MChogHMUMx6d06/8bTcVaEvH5l5r6XbyUefw
lgmm/GfrPvW1HCSckJ3ftafwo8Ny/cYN3Mst8fd9lM2GcnpUjP6j2WbmcIglfnmU
d10xFka+MRvLVxMgPj9Nt4wIYBuep6xMgk7aB00AZl+XdfdcRg19KXtAB6DhY5JR
Fb2NSYcypofmY9yTMqY9pZ0/vk86FtF6wjukohMoQYImyTWacjR9HyYonTHJyUar
IKJpT0xOl4ZtJ0dV80dfC4xob5INP/PwkORkbtj/Gzjn3Rxptui09oK4G7YlFkwB
Fjiq8ZWPa4s7enBtUopiqN4Wkqe9dkNccdwKDitjylIk4M7ve2uevvSO/i2v3L6G
uQmuGZJA0dS+JCcxx43MtChCknibtcugr3QgJ9vm76sVeK8SEUDyIhB0aEfhaqzs
iRV6TJ+nHSYBDqy8bw5EiTi+gpecaCnI1dhz85vCudKFyfS/75SCNYoG5UoZSJTy
1SUx29/x2DCBeJgvvlKTicpch77vQ6SD6xpFrK6yc2bqJkYcBNM7MPZltwTykc2l
dzWnx98Aj4aJoroMrHUsYl8ytEDZ6XexsqRFfyFDKZ4fKFz+C9Eh9uuGjWhXOUJt
2I4aGrbE/KJkKesaIIZM1zqjB/TBnOtp/wHxa9hBMC5gJBHAfQRbbOMfFk2mYyh3
sGoSHVsT4Nalq500jyAmFQRtaPn8s4qgJ91HGAgvAii1yeoCNdYv7GbPUpTBE0qO
8ln0zBlQMKABSFcxPdJCv553mMxdMH056BDAdW0hOPswocH2Qt4sHN/Hmwm87LwV
LSIXTFN/FSsXJ3rR+59k6w/wpB4IF92YLpsSR0q1aaMZvlRUwztc1InidvF/oJKH
2mjDWonM9H0YJWr7zG1PPqwrVYhoDRN4Q2zOadEwJsmlK2113g/x1K0yGkHh0NH8
3va5OG7As//SpGgGQcWfr/rhi6/tUREKoGsooeOaPcfUSKcRMEZePl5t2zv+9QSD
LwxRJT5A2XHsvKNTHGSPeHUnARi9I8CQeuMpT/vSrH5VySiOVCeHbzD0Lc6nPfW/
dCdHHxrGX95LRi5v3yEoHIfRz9JWCiqNUr4HwvDMltBmn/crk3ddDnB/Jo2FfHO7
rr6WiDTZUS3uJ03BupTFv0IW9InjKlJjPVIjkuUACV95aSRFEBRYnlWxr7LieaOC
jZAZECJKq/Qg2OV1VmGZMfNfL7X5QoUVjcBlPM4zQl5cD9AW45tsuavLQyCgMvbk
mZMwJaNeJfVMOfPg0KPGyDPv2L+3P/F1HvWSUMLWjfxfYAyu2zl7apmrluclTCHW
i3o2KKzhvr+Is0p3ubQNAw7ai7zGdXUqbYJ3flM/ga9a4nO8uT2jmB51e2NkzzHn
RNIYD7GSlxEo5Dj64zvOMiciqWYXfQelesI/5XnRy0O95sBdJ3OgQh7OJ1/ujPl2
Dy7aSLTC9l9u/nfZLHL98BW5ZTvZOgwOd9n5rdxSjPBogmJgQiXi53Cb4UbNqSHi
jeWRmgXGsVGAF8zj/f1yKNd3vH6Y3zWJrML38UWYY1b7GoThGWGGUyYpBryTyC2K
M7CQKDmy76emTz0REEZCdWzkNQHlcHAxz3VDAGRWO6WRPzbMGAgk4Eupxur/5RlU
D5d5jTNLhmfTh7Qca4j/4gPlHm4NDumszMYSkWHqvJC52HEYN5TT1gz7fBGQzlEu
P0rYLzeH3PQ11Ot8BP57urd1ykKNOJieJo/Y4TYuA5ecq64+XvqxDETNAaFf3C6p
NKGN0w9zVKku0VyIRZ8/wx0HnB/j2pY+KLPWq/7oVMN5TVOU1bhRghZe61/imCOf
yspe4jIlzahJZxASo9jbvKV6rq9gijvqqirrIe167dcoxq+IfCKk4AFxWJKvL8OE
3JnIyCQdqHhN7KZt3Ld2moIsRa7JRWVRopgDbSD6e1yWGk315QbB964tNOx1B7fB
bvT5iFOABv+VgwOpHUD0fBlzm6WXbAQBcc1p595QF2C8+a/Acseg4fqIxL8yJCnH
g41LVT3pj1G9+7Fg9Bt030n2PQ4p3YOiz3uzj1kmTT6Phcs2TwZVGFEbOwtfbeR9
wrm+wTgE2UaYv5KHomalWXmMwKVUZDbjmTu1w+2SHpIwL7DQqYcO12os0sHIf0cg
syAazJ4NZKiwFcD5TXImbz+HoZTmlds6s2VmIsapXtv26IdGAHDIHZKM5Op4cNUA
NlbUKj80x7MIkVs5qHH2BsM3BrFOk9JgAvHad9x1s7cbWEGRyIZsLr7n2/B9EDiU
vTbPKjL0G5LnepZjYR77YaS7S79ShljTYMSmz2i4Q2hi4lmYYI0WDzsv3fwctPSb
dYmho4JkzYuId3kgfieG0NxVumdmHr6kAJHpKRCxM9zYZHPRBWw07uXfNBkd+VZH
nB4aVuTVQLRTwGx4twWvPUe3IjRa+I7WKVKcO5wmyVSfHl3T3qDTWhYuM9r651dS
r+oy0wXeEtaWvRrVVOmkJj7msC2bXGL0gsC9tPosJd15wmEHnDK7q8QgFRSsG9sU
QFb2mnHYRtB9qYuMGArBFvME/355d4QT3MhHl+cNx7g217XPZUVyoAQnny9+FM/U
3TPRY4u5rqVa8VUm6J/EbMfXs//P0SeCmF2wqiUHrtGXoQt/YwWSCe8g4zxcFmQs
kXXhL6s3Iewitcl0KBFiLuhKdZZqXBBuFxwi5mQRDeX7M0JbdnxQit13c4qVXG3v
8kqNH3H71tvuYfp8Yzkksh+80vP1GMzkGPYkL8GPizJZXUPdyAtVePpsvpaWLiKq
skZmaSy06N/E2m26sYDJivpMOFk/BlsDE0Ks0BWGFKiPm3mGAoGP8LCuG7VZdKM8
RXJ1DrONBj/D6B5T8PGQB8t2AFmHoW0Bop54/750/oFj94wY0PyH2IKH1bPXesIb
awY/IL/CE4SeZLDcog4BWIggVGdnZ+D6liqwscc3QXmUl1tQ8aauIqUxoRBFoa8/
PTebNWIuHiQ8CuEyuPABEKXRz1mjg3KxlvMp3ElTbYEcKIQK5kInBPS+07kKFigg
pBIVZDG1bKmYSDw8NjP8EXFxid8BsLPSEy5p91eFSP/ru8ZsjlM4PQCzQAd/NK3/
GY9NV0iEFz3EZUNRKa4ymslG4VFF+22SKU5he/JvpIrPjYOuIYI9+ACp/J/n7H0w
FFgkxE5ioC8Wgl5qkWdzvv2u8rRcgyixaufrbK1j6S1eheMLsDxlzyBD7EaDlm9G
B95X9gawyxFDgT4FNExmEfAGSDN1lnb8hKO22oOm2DgpnHNdsiBke+5kgDRLTFv+
VbIk0Kp6xwwy+JQSvzTSLveqqE2ZyAd8y6F2XGhzAjmBH1B/VJuM/JhHtHWwdJWJ
QbSkwSqUFtZOzezfWko5boMbeMho9EShi17/d9sUSQ79eJPEC1wBXAz4JLDqdqOx
qE8UjLrQxMQ9FCo1oIMpoSPgazCTbhnW6aoW6+J+h6l7PaZo8iWPHsCFxnJabShV
w1JubnWkl3zrh3thmk7h9muk1X6DU4IDMfgMzD8rYpRWPmuXhnBDq79dVsso0+In
FkULx6+pAWpoy7KVoSy0KfgHVf1H/sAaIyLAq8GFPTd6YqE5rocZdvJ/eUpEWLnC
89zdf5mPwmnc04nsg2L10hCFqv6XZP8Kwtv2mr1cO2OehTYrMXIAd9dtuLAOZCvv
VGShjIrzCRmqaJkWlO7eu1OMceAEBikoN7/jeNZanJ2MJLNnA/f5z7hJaoNsIqpp
XSLH5eYI7+WL4POIVFkTL2HQHX3+9K8q9k/tdqrLfHdO5Sb8/vRWFGoBbgspuUJ3
4Rq9U3814m1EVpGjP4O/7CZYA43OZFIqaFoaHF9LlTTMM/HrCXO5gtxtilBq7QTE
l1vC/R49X3EYlr+sNLnCvzBiqknfA30eSyYD3fA/LEhsPTNNHixGq6hiqCcZ98Rk
lX2F52sM+c959qw13/pCWIr8IOvfQbg1j38OrEOGmkA7hx/iXi9k+eA7lqb4dimI
qQ6ii3VkMz20OLd5ygGb0Mv+YJZP7cYKNI6HKCVGajc2IUk5fhOUoCrMvCK0a9fU
QBFLc7ZVYUEhX98OQnFsWqRQHj/f8nyLFhb21LCsoTPm5dk17YYtpHgZgpCEnZCN
NyiI58u/YODSvZSg85dT9bjLUShCGdMmM7UBcjnoqQzROK/uc1U/wrWKxxBhdCBA
irvSEh4fCQwYtyqIZI70KmxnWfRHr4ZmxmIRL+HGOWr1+Xqs9PsmYQP9BkXcPje2
Lfawxy7/wupdWL5EZen3e3NpL+VCHNgxcwIqjAMnsFd32p3q5l7VG+5C3k2JMtki
TNFMp1kuFYmeSSjDDMjC6hjmLkta3KHHwCjq5RM6mwZXl0X5Nlnrhqcodc/nNjFR
Dfq4BHzOFHf2kkNJ3QNWjxyxm2RDUyYNIje6LKHiZOBTzSTQSju7zpXmMAHUc8Xh
u21+nIvuLXYmyt6msvSL3k17LaguC6dV65UXxfAI9ZzV6fEYcY3MkoN8v2Js6haw
H/C3qOIX+P03LNo9EgwJ7PmeaxfHQj2W1/41OEJjMsSsm+hJm+1ClNubZqmTRKr3
Esdc7YwnxS40OoaMvdIQuAm0Psfj6ArkQ//THGjGLubjFYr0HX7BpXgpAfX4k+um
1rlusMzi0fyFFMwuVQOrm8+yWbscnMltlyOWtrxqTshi3Xyaz1h9WSwY23xOhiqR
yWG9fbNJr4mdyrcF3rcrGzEpLe/4jKql6oVGjPSFbGskP5pE1ZHmhY6N01Fa8coL
w0yDPpjfkdO90BJ/HtSABPNl174Y06rFEoyZ5EusC1nVdlVtPN+2b+O2i+4kwkHG
sJCmyMNrrkTlZdW17aadhsAsBpf5aKfo/o1j/LUYnBBEFYJLfewe4Ylv9eeFLY3g
XTvg21v5jloM8sk7NBkJeUrFlpEgBNIH6/0vxRk2ZbC/tsBcJFO7di2vRhbiAO6e
6Krmn7OgKVQVotYlnw5kD/oYBOQA5PTTPJNGYg+rcGGnGKvJuxQGFarnH2/fCzJM
xZFK4gpEJQTprp7H3nxuB3WTunA2BoSffNluSS71U72KCSjSkiai+fjNDgIfojcA
MTHIAG6Tc18BkCTR7dL4+Pp0153I4fjwoBtdNBAUU4SRb4T/kW0fikUAkFLRkYUA
L01sYnroWRntotyNvFGGsjsDKgYQ+ikVF9OP0hYOzA0oVd88Q9meUJBRLvaqtzez
eDx3kPLsToLpyrc7FanrYKNCUEE3fPtf2DWKcpP2I+HzMxIEU5hgwVXaHHGoMeD4
TmLnJQovTZh4OhYMJBtdlyyU7Dknlg51c3g78gVui05oIhWEVNWIW9kfy29snWQE
eTE1gQ1LeqJO1qYnFLihFhcN/WoJD4TRW135zMALer7whuoL+2Tmps2M1GaIJFPk
ojubUGT4IgUCgrxyVRQauD79yBFwsdg9kwQL7wLtJ1lx6w2oj38UNY4PqGIF2bdP
CAfcVwCSwm+G4EJjsIZux33PewWWmftHqJI218Ogg4U9tLTyO2zQKDnTtEJl93qf
zL6PL+3/zvSfdEw36qjfcFGnGpBu4WhNq5HviJsDMQLZj7EbQ3a9EpFTZmrR83eU
0o06Y+0c2TNJzdlI4B9AbbB150CcrrFB6WPMnd5WSbx6d5TX/H0L2c0FNQSjn1IF
beCTIqOCWb2JU0our+p0VMZbjM9tgbCb1o59pCcd1vV9A5UDRiG5TNJzLjAO+nbI
rZpGnMj+JL4C+6TQY8/WBonfapzTya17aKO1O0fu1ZoZNnF7LmaUUIZ42nkNYJP6
gUl0sx+4iVMGhLtQKle9XhzEOcenWeYdO9Z1qZVSaOeBnWGHEqVCqQEH28pCiiGq
NvSHiDZXUQ0WdJSiq3ASoBon/T9wQOfCdp6BsF83uJIQUXI4sanI7h9uVsjTLsYN
wm2RpGBOn2qKM/Eg1/R1nEDs2qFVGdAMP8Wfxfgp7Bjt4fb8O+2A/AI/vJ2nuuYO
IUHCmE8U10kObtdbx+dZOLWsnkGkVhYnueEYfMo2Mdb/sfW3HEWMs9LsOSUqpHR6
JOiNTh/y5+o3FudejMNWzlVKDyZQDplezfxdLVL/0r7TmN/RS5v4R2uy+3nFkhrC
cHyHo+CB7D9KbLx/wX4mi6xgsGDbJfL10zg6v0wfUeXgmSu9XYT06RserOQSu4KW
GGlFMblmVO9UGNp/4GWOSTbpecH34zD0wMdyG7KoJyKBxABfKci1k1LOU9VOHvfk
OGgttrRKVjVpfqwkF8LimGE6zVJ1kmCs5A4czqSPXTIcWSrAbkQggd5EzlOXJNjB
Agz+kErhFmmSyas6Ny6WMyw/KZUql7yoPvm9wbKwuDU4DaMVawWu/g0iXj3t5D/G
8oZ0KoZKz5YqcO/fWZpIqLF1+YMCK7In2gp098Cm8bY5HfSOnweZ9tzlcqt3ux98
Fc9uq00bgljK4VJSNEzDSbhRXLdy01+43e6NvKOVqkZQzIVkA8nfFbj3gzA3pXMY
eRZK1Y0cAy9+xu7ozqx6j/WEMoDHYkOtN4Np37d/eB/NVOYy7ihzwOKOu+pQDEHo
C0nL+983jSxPbIFlGp7m86qYFbbWM/Lst8PWRhrgsNlH3sHMMvPHU4zdlLMssqhE
e1VArWndraldbFkDscFsYP46AJb9YtqugjZVPExDknahQysL5M9MeH3SSuiMHmCB
Q4sBB+880nSWnoKAx81xAugShqjEpgevTXgV5O/eXQvOln6fzuHAtBPdYbgnMu1d
8UMbMHnC5rSkDjsdPk3j0zs/8vv23edwVILqO2TQ/0kqxYEDCFGi4jT/ZJXO33Us
awCgUcLOFoJe2bC/zpg82oM/loZOR+2/A5O+TtouLXzl/8NxuXGDxZzh4OCXvcX0
KMHPK7psRUDK/Bn7BcNSO7duxdyCY3uq/SBBe3ky7oM65pGcT9GaFpGYiVoHI5AH
UvnAsrOmQdGVwg9yeFrTOYEkP1xontMVXiZluSpXBNIhwj2v01i2Oei+44kT8stT
ko9pifSxFTDdo2hhfu69V8xztYP0R8TwJumo49ix6VMBhY7f0mZ70r1OdcdPO/By
UtZrYiIRJUFYsS2Q2tXE0U9LPKUdEV2wzVEPWWTJZj/lD6r702JbvRKLC7BLBOqR
GHyVOqL1LnTnCVDqgcecpzFxtbBPCnaMqnwf0zWzdWDvGwtb275gUDR4vrySpyDB
BqYAxWQzSepSN71GNbl08NFejUv12rnGeK1CiiIqwVrNotnZqLrOHRg3gvawrTRw
lMqA+P/lOmMcNCVbeGK8iKb/BkfOspiLRnbgpa5cDvUDEtDWUHqfIJAuRNkGvJ0c
GvFdx0IUGBCqxYJp+X6xS2Q7GRlYzLqAHFvLDrIrNvG+z8xIISDU5J3w1YO8HyTy
+V8X497lgmZP+g84RQWU8fgl6doWTI18rILNss88rALQbQddgY1pr5xZRPeNuGtc
rBjJQjgG2OAarzlQSPy0xTCy4ICQhYHH0gKw3zMJDbc1Be+3S6tfY5Uo4wJXlU0d
ZLhvkm3tnYLzpOsuBgreT2Vmkz5WKG5up2Bm+QZaM0IlMShAwPOTOHXMUBSoROrk
jyjI5ZPAuDxzl9bmSV5GdvIC2NEXFEL+GCBEdA4ZXkc/aJNJ1KclQ1GzY4F7JrAp
fZQVn+Sv/Bkj7Zz0xjHFVjpiLxSdabDTBHnW5cJ7GaSZC/Qj5qYrzaKWS4YEvx3s
D0Mo3YhWVZLONGi+wzXK+bW78U+RXdRk4Rq6SyJt22eUibBskw6p5hZxpHGmA8gt
Avq5QseekNpLPdtHs4KFN83OXDXMvUGj0kORyE+3QbjHZw8nD3PKCDu2qMGjc2e4
0uaVYXSK4SqajLKp1IjESp93Zqaj14VzBX7qblVRD7wUfDQAZdKF5umqXsGgJT4i
VB3X94vyKM5YKxAE/UyWQ09BXNl7QHBd+g/aPtQMsN+z28N8SFE0hOtIbjkTwgE5
+2pfgINKVsV96FuVs7TnH4P59xI5PdFHyhOvG/H7IqwPz4L/mftTpZkFi43HzSKp
a3whjEG+YFFYNrykUszJr3kgCEIDJ6L5LemOVl1H27CtoVVR6Wg9wzg9nASvk2cY
HVmYH1fGPDupI1fJNZI04cMHwbOQ5hhNt0sPeSwi8/H8fkFMffKWepfDQB2G537i
hA5hptCeBJRpFs5HF+KyZA7ab3l5jkF0kvcXuqmR8ftAN9h8ZX7rH9ozn/nhmrPh
3jKedJNxePEj48RvG1dRPCUEZmTR6ZEoCs38srGx/02wgDJODUWl1b2P7mhT0btR
yJQt33zNdBwNoCne7HyrcbDOx4xpm1rcgWyw6YQg8VI5bFWyPAprmUmlXtdcfLue
qw3GeDCxuptoDKoClhZJp8nFE8DiUXa1WKIR371X0TRb7m7wsHKrb0ZawGoP3mdR
59lDSkp4KQe8K8VzLetfOTSR6uoyphn0dPLcEPlwWqoctedfk7/YMSgVoIdWNd6m
luVpymbczf4cA0ehIJraWoxrH0/+xRQSwzGDLE0mWX1IXTGRK6kGc7nqp9n+SNBV
D6A3Xni5ne/SwcW8huR2OyZm9qP+NeNFl8zS+NT1rvQWqFp1dUG576EafwYvNZxI
+nbiTPejRbBvVql/UQsBzjjemNbECvEUqGY22BjHIyyKC+ddPhZVLoh8bc2Kq5dE
VEZ9JOZXrjLjJt3H2LYjRcpbORHQ0yn53S3iTbjW4Al+FfuXoYUSD7VJ+tmH9f7t
RYaSX3+/LTCuSq8j735Uw9G76aChYVh8lX8xJyOLTRfpU6/QgCEeyhkXMODkTqly
Zed+X74gCOsSUk9p9/N06Zp7eCYqQ0wXSalrUZnByRO2aQdl+L/yH01qmTbbgm4J
jAq2ym3KSeR697gGkSuqC+WCvViKD24nyyccTvaGq3nVoqlF7kevRVaOrMuOvsEY
Cb8Tqj/IZpDfySXoJW0D//sKCM+BA37STIUvFyje+PVOPq0nm2lpZlQIZXCTZnXJ
EjhtWuz7ANY9apfbCxdHRNfaTsi951k2RxdLV3QQJI6R2d7GWtoPLxd8cY10Ty0T
Cv/gH7liAthvnQbRUT/LswbL4wvRGcA1WyvYi/TYBfXA+DDZHfySFgyklHmXhv6d
r67DyU66Hx/JNniWe3UNwfLpOGp6FJsTfoUHuW0ssE4pHFyTcZyuCwcxGK3lRnLZ
jxIaKF0CQBerqr5Za1h3M7VDeTzXmabkUNE+LgI++i7IyMHzgdC6BcVzv/e/KECJ
Ju82KNoR2fk9NiNvlrEOfCae5EnXK2iX80bJNHj04yFaY3RGuPFwBj8rURHe8N7D
3mBLfYM4y4upoXEeAJpe8MtC9QQ4ZcZn9GJVQvdHDCqztQhXdKquCUpvilDVoS/D
1KvlC3PwfDhHBTo3nrC8TTDmPBebt+Oi9ieCi4PoqhXAuUIswXdzJOD8ZKhuS8gb
aJkfN2UwgTgW9ItlA9IUFZPlGUJEe40fvG9cvGkMq+IXaiBn2+gnf1Na/32ckLSq
FdQfWjtEEqYO7BbEj1i6aM+NFmCOwr/bTX11equhReM2A+nGSSgSz6A99pBSPF6K
G7uYtPFw7K/ZGlzv5QLw6Y13ZAa1ZWf2MiKIrdw/qM++H+IyF1TN0KD0jAIYGDYN
pUeHGDFdbTmboD0dzCvGvcxcfMTzN5xjEXSBxaWqDDSziiGVVY4IFAA61Ktj7Xsa
4NmX7zBlKIzh/Ca/oeLYBUssio8ll9Nnl0dLnGClul13qx66A6sf8bSHc5xbLm27
6bkSuwzsWiCEDKZ1THXV6Io1G+RV+Pd5pt72tLnQqH8uVZ8z6LfZnqKrN3Z2bzcK
cMUe0+fVx9vYrsMPw5tbql/4eQD3UB4qLvSzEFChId40b8Yn0QCaa3titgo/z5xK
hgOQh+Xlhc1MRm4B43Bqa4SC4hyAL7MZklb5E0SZEFIsRyCgBmxKqGlUc17kupkG
N+VUK8di3XmW3TxMHkJyGX+I2evKWJf+QIgkS6smDkSD/wSKGKxN7XQbGBh6FDRf
s1sRBUlPqO0RD2l8HPyPlSVdCy4vO0TpZDxHYCViWMzJrgfs7IAxz1tVza40iJmu
ggmGgFkMrpvblVcawlR37b1v56g0LE2m+Kvis8K+OrilntLxR0W4miupq5WDkIFk
IbiWsWPYIroizlS5v+4xzojDjpKrPr+KmMLQ6i1H9w1hy/l/rJ0SPKAmSKoYyk1F
1G2qrClkz74/HUYZGSffze1ei9pAsP5naE0neN1tk/nfcnGFqQwkABzjgSEn9Zhw
gch0gY5hcbw+ag3FNdv7K83oYJ7WaKuIMgwGnyg5K7M/H4X0Z4BE1TQTqJhLL2Pj
6JRml46n/+Jc3xxc8Th6omONkV0PIZT+YLX96C/Y38Pp3mZ71hSwpTM4XcSQvpbL
vE8a23PuogHA2UdB1+PfcN2JW6406U/w/l30/43PHXAREkyaq91aTyODFYJsbN7S
oJoFfebiRR2gPrsd+vYm+FHv42PRKKn9cGJyDLZqJvxTSvVCD9YayKVdwY5k5lqF
6IxyFh4LSMZ3+TXi2Urg55uKaOwEtXf1etrCxJnfgQjuinJz0Gm95TUGdSsH14vR
kFAalB0LUDVIhYWQqJMdN2Gb8tNv9kU31ZfZxkQmI9HVyeHzLJawdIpNCYCtG0JL
rpSJ4/gwwAkoEmm5ehxpVpMo7AL6Hk/7EWfB/cUfacdmfpeGllXiEqSdwLjVyxfW
Yfnyl8YAxRqgbev30RwCtYl3cau/NTjH+zby/f18edh49CHq9NmA+lCcLfkc33uA
i3Lp70Ka0ma/QW080UNIhwtfCqPdVaHjhfvQR+tj6AfF1qhJVk3toqRDTH/4xFHW
oBq4lO7xvCoe6an3E/lmgAfC9Xj9JijIyCvDYWcnOoh8J22E/slRKigbf9syE2kx
pFl9PWvCkv2++Xf4Y9BSVZ6+TSsE7WI8PGlHD/N7I7+0MUYXgYdXaBEgOSZLmptb
Ay7iIUd/KEZwrzIzVuRGDhC+FgL0nJZD623jt+OPAMc/2WjP7EJgX2FuPfRVP7IP
sdWTlzpAfmYJNLiXQZdYsYvdHlb3D+rL4Wxnw6sqwe2JzShR3nG+wNyrzSqePmjJ
tftK7GiFpQ8HExwYu2rV/fFTEKdo8rEUw3FW8+xIHt7ZHjxeieyN+rE57vyYfx+u
wqio+Rd5VHZoi6N3j/t2X5aJ+cTIvSwkVDtIq1OoDYJpvPuPihDmmiQ6olsXUKj+
bTeB+1U96XJU4dAW8C6F/vce0rJMU8dYT12OK97KJiR/e034Oc93I/t9x7ZI0GCX
4+H7GpruhzZVIr0K+RNcEUpL4Y+f79SLnkXphtJvPoHxN1FTbQYno40heymdisEa
01RgS0h5sdmtuZcifMUNSpbxQ4JlnqoqM8rehypTqaTYRCqp2El0TS/rJ4LnJTCy
LnBlj6Uv0S6JmQjGRWTOzhsF9cIx62Jw5DQ+ts2QeUKsWdczqMU2l30DaIqfd1RU
mUtEB7sJs+UjMfxK/iS65ZNVoeWdNvZDhRKU1GcjABKIc406wRdGta29soXuinyR
GrSTQF9z1umqn8+X3N8TA0xo+GEp6MHYgdxi5jXsySgu+6q6mcPeuU8D5TQ/WJsD
a0VGwY7ICW0ldPDyyhHxzKr7sxR0EGQkmRYKIjKHfNj5OHjBMVJ8Os7/UyjqbbzR
tIaJTAHAabPWb1Rp/+rNhZWg8ePeY1TZQ2jHUBFLcijmcrCmx0OL+Ou4mnqwmUZ1
+/XyqP9nsknpEgfqM/DCWSNExh7t6PkuWNGZSWf7Kh1xiR9xnRyxBFHmhO9JPvxw
eQA0aMEjENzyKfZakbNiR3LiYERVJecavgubVp4w7PnIrbj2n78/WYUCPt4Dr9Fv
dY9GegdeSaavHoaXIbC1W9sAOtp2tTkS7D+0Skx/HNh6HxFaOQurGDapnwBNhPJ9
Ieh3awH9k/aD07citizKXiBQGkzkLyYyjGo80FAjT75BEOwXmEaqGFiE6Ug6d/QZ
9bXmiem76FpZ8UZ8GL7bT1P0Kg+CMWDs8YCchI1o5YtCba8Xd6wRsR8fJc/5UFSg
3inDlwDsyH0+o+Ivp/bNhaaEv5hUsNS3YpXXRA/jen4p8oDIufAzQnrl2TGyFeFG
W68ju6VIgARF3ck+nFWieTdJ8WGvsFu4sl4lpLdJQ7xdI7Dgh9GPqRQ33du0mrw2
3o3BWAq7NFV5x2VGjO1cdhG6gok4XSxVDCk/QjsHBEt+pRaHbyKl3gSKR6g1txPj
8eKbI7/GsVeRFc8T89xTJbSw151GwyyL7/1aLrnNA834jUwXvRrwVRYESXfLTqUy
FbMRNeyTz0VuC+fsLuNAArcUrn0s3eA9sXj6HVsdCIovjutxdB5NNYCg5NeoMqLV
IKYO9xy/Umvp3gKCFHRSaIG0KG3cWLQI3bVrUmG0zFgEWqDKi2swgLBekrGyUpJU
nFfm/M/GP96jpI8exoDQHW1mDLMNZzwdgCKTqUPU/S/tNEMITiOmgDQHbBdvtogQ
naZhluuQjKE7h2OTfDvpgalf1uLIFfbsYEfV2TKt3t4h8Kfp8cynt728h7G9SAUc
sQ3Dn8MeGLwIoEfCL06+ccgJiztnN9FF5efh3d/7exY5ib1+BfRlVhAmlMvMfR3J
3a7537hWpS84tm1MTHn1hS58prpbym2AT0kxUIfPl6P7V7iBMA57L5zrdqd94RcV
Svdy5zjq/DF5fr49nIwDoO1rIpe6xnsxnJr40d02bNeafJHrh5erV3+OdrYFDvaz
VenJOx8UHGrctpx6plWNWwr7E0bf/dz9nl0mtxBIS1cWN3fEshvzEbYNPqXlCHQv
tFUen418IHMQht5afNZVSuMpCE9kpf4hPmvBvhLQ1rftOqUBNYFAYhcLVAjrmdrx
LMEmyG0YwL0RMY+JAK88C9LtpH9P5vu6dBUzQqKgTaVg8pNS4bnkHM9L7yRPl9PZ
E7LEhzgiQaS1Fn3Lb2QP3q9khFvSni1qxtDh+3diAeB9RlqWQ468TGaxBb1XUjwr
ucpbmDOtcQv16xkH2d/u86HPqI2Hb1nRjLFrWRrQvpUf/saB1s2/Q6s9+YL9gsSv
UcD6D6FoVY/ZQ/DQ0+VzTxyHx4IL9a+6d+auo5XrkimRNNG3bHNtHCENJeoPDPGN
+iQhqKVJjw7MiQbthNZ/NFtq5RSadpjo0f3kcLK95LuRHtbzhGhDFPhPYKAY+Fdf
1amed5m5AbZlFUSvXZYdkXzSVCf1y6g1EerVStkFI3cl2eBZBQmZVrtavvJ9atTJ
9ET0HWtH8fVMWt5dzBBUdZekwZXN4FOcnrRbjw4fASLXsxC1Q+1Cy1CtqklUKjOJ
1V53sGnhTdTpmYwH1lr/SpoNpgIxIm2/M1hlogX28kmy6F46etLqXvK7R+gcbu5R
9XHZatJDvNa8Kb8QKupNiQBUFTjwub/LYKfJzR9W99M2l5TGi9A6+iMgHkNHx4VN
DFyUcf8CA8b67FnKF9fSDSNpHlkZvryOhSqrcUL6nwgO1wdAvmPzxepluu2WljnJ
lNciU4TdlfyqacLiEavFojxr4Q2/OdwxO3Df4lEHi3nAoEDTylsD86y3kZ2makKr
vEMLhm0tO5TnsrqO1qX37LqzHHOX/xY/TO3Yp1o5dNkwvNtLLlGyyH5o5BmmGa7m
4jTrnWRmPee75dAPGGYbxT0Lqoiw7CIg+F7FAlK9AIlKQIZYQ3BwUjoywdiVu8gS
BEOBj55SkRadzFUo4ODRO1rOZiv9TKH4sxX2Ug44+K2DkV9zelsBfrYXcCTLQaHA
t3t4qoXrexbNTn9FoADfMelXSpeOuzDK3TpkhmQ+ypfdDtsQZyUt8k7LmAmVgI+m
FnBhxwCfHFuFqoEpu4X6cRpUXRH8Va2IjIycdlFNUb2aEC9hDltwlCKlps9wJ0Bb
kkNwhFU3lIWfytB2BSmRQ/TbbEHpgJdXKcWRFagm4zvsY6fCMHeddUoeaM6jmZ0e
QJZBV0ZOUQVzHL/I8FtKzU6cR6t3XmMPTnxfQef+sWEwdnmOQABa1KQP7hcK+ZrW
tTtzcvCMa0eIzVBSy2iRySPv97J3pGctMu/lsju+kM2ZsxD153c8zZuSmfeaf9T/
LdrqcvIYEy5OwSyyFpm1GufhXAy5RqQbAnr9vtTEypQy/HqcNhvbpofhWpkwAKEr
HVZrIJLYLoDX3lAKXyE+LDD4T7xJDCsDDf4cN3YTNlQxbOOB+53AjWiwtJrGggWJ
7X7kat+fA0aMdKqfSKSCf3cnoIBOK1KK3a2XhSl4oI77CiRJLl4L1EjkbRcrKl2X
v/BFrNF3UdLAFKZrPcbFmvz2ByE3PhiX+m8xvP0DPwAhB5wDZ895DK1XMlTKTZIA
/SurvaxW5/C0zk/FM7cvQLCZzsC5+b9+j6/9bK9GbWNNq92BjxHQi/aGix+bBghi
2jYTDne3YjBE5d6I/faA1ZNFz7RpvYT0PtGL6ElN8I287iFVjzNL5jrds6iwRH7c
JG+eNGWKSaEPIbX7+qPuOPt8BHv7fafAOlKY27VralD8iLIG//m5lYsKcm8QMHTw
QAcP5UXhqhNsfyXAEa5X/blyOGfIDF/MIE/qlVlk3xjMzJjCWCYR81fnCx0YeEr4
9y/Ri5ncNGa9G4IWIpBItFMgYW3BhwY+ZzZrCnHsk6k4vCIUHKJVWstTAVcvj6hX
+UzlmVKESnuoLuv6UM1UDVC6J2/YxYG0CvqMi7spmy2t0IY5yLBHr/RcSFQGgRjm
LEWmyLlmHb+KrZYR1oJQru2gAFtMMEd+NzC3FAyGk+Bf8QhqYExdR9EPPzwVHCi7
JxxKoCwhD9xUxqy+2FG1Oxq6UWophPacLMrxSJfz8tnk8Swe1h3x5Y3dQehFpYds
cyIC/Y8qxrzDebaylJJePjMLc73R3X55/YK/Kg51nJpxcOILO1YXMzphrjnk22eN
2P/ox23EvJr8wVbZD6vEtHxy0VptNxYWtmH0xIMRmEWNP7YbOJm9x/I5RWotbavM
Frzbih8A9i0nour2inW5mU/j3GrpX0ZcgwnEIxjq7nHOnQ64SmnQa7+SRYTQvTDs
0zy9aNT5FxeEIfwNxtnxQIYlXGTzh3EfSASF6FtTTLSneoPBbg03pD3G6Gywp5du
gxhiJMANk299yg/Y4B/b9Uome6vph7ZpApkpHXqRMT3Gs+wE8pYbA34GHLF9kFwn
59Flf/WSNszEOFyRn0a/+M5MJxc98X7IDHtC/9U0EEZiNjMcLNiBwzoJL0gM9+yP
IPHG7u/ptflfE0rRuoHgn0/0Kbr+4PwbEARZwzID5F/sOb9LcUzaXTAp5uYKGftG
2NGnSAUyas3tn1zlfBEEDNdRGW9FPAbNq4ej03S28UUoaypULgB3ISB5HawAFyp1
U4RbimUJfa4IxGOLTZwgLlu6RMN2XStLGS8YYysK7KTzsM8cVXv0NfixouLrZ0kg
nBKvErn1SOkOnP14evytQSTcoKDWD02j2x29uHU8c5KyegF2tpTPtkVMbCTJ0EZ4
oRCChbVvq0S4M1SxBgWAsScqmCrJgmbBBLrts0rxjfgSvQepGq8qGobwHz5eCN83
ypdk43KGuoWuItkxu6Bb+p/+gtVSZQUML895CJ2vhuefCZRofvlqml4YVywe3vkZ
XEAzWvyksuNcG13rLJxpL4p9Fy1mef59zhOK6Lo/MZKtQwtIcLwO7q1p/4cklwDU
mRjTFUyQLYJE95cbc788OozX1cSxaOfFRLPIdHA6eBKIG6gF6Po1X/YQn2vSUyPP
/bcU+ZsJ0c75XlLOiSGN+owHpXqye7Yrm+qZ39irw73mqz+y6flyOc878GmHe3Vq
1oVtlvtBKdieHX0gmh0G6DJ8Tt70znRL/cQ3GqwCyNTp7Wn3jQpHvQU30ANYZBH9
Kwb7O71hK550E5DanTn7cN2gHllxwGyskXV37/3Zw5ZRliznB+XMLH0+YRzScumg
0DODh5JBs6q5y7nmQpgQFqIixebf9B1/youbeJEirBAVpnqav7o/wuoXjFvWbY9E
RUZs0Z6IB2mql8TtXUZ7VPr7DYfuI4nQRq4Tuam0JEtrpcO46Qn10GhZRMvX22cc
O6WYLjGICDszLyhkUOw3dHoziu+hf/Z3l5D7oV4UvFE8nu7FWRAfdr9Qf1nBdQfV
gFaYfgY4BFAwa+nitOgzP9O99wRO4u0frz02rZw2/RbA7zSWiRfHR98gOXRgpj5X
anQRImil6Ia05E83xlDtJWwtEfIjCozf1GpUKiIOunW3uuPb4xaZ1iXE/1BrUjiC
iWr+SNhFvVZ2aqfHDbPLspH1QOiE5Ex2fQ76VUTmOsKD8uBGqufoGTidwMxeDwoR
AIizN39Gz7cW1/uLldFYcJrJ9RAqi/UiYUK/exqlVo2ZVkuqT7Xp6HDTNWSLGETm
c5T7rb0dhDgEwNZMxpO1GLesjiI3aIaC5D2Gz2qVfRJ+0DBPmK6UQcvUq6E5Kivz
bhHEX/7LlulR0nR5CSy4IDm6sxK/SEFy1BeNyRCCyny1w9D3Yg+cq73M0PjiUesA
bCvxQ3NgMjM3n96Sl17C3RjK7+t9ddJmO3YIFFVYIhxh2tPHoEQ+81QD+Xj+o6Ff
DJ3KK+/zdgofXRXQ+OsJ+yx5ieo5sWPrP2tkoCwEl8nQhDvkbKqGYWuWPwTr4uVk
F5vfpSOG0gTUqq2xfShtotKfh9C4PBqqaB/ONKqgmBKyefSIYKYdDiri2j4vRNdo
wWr0zMdh1SJZ2sbu+XR3NiEsj6to+vRFHCkHqspWhZE/ndvIi5vPEbG3lR14Oca+
H/coPSfQ4bYB98Wsdunl/04NsRcwsA2fIUa1kwytTQIklZPvlmULDn2p5qif1CA7
quQy+efL9QizJG1eZEn/krXRmyHkbvdiXNeELcA5nVc4HBtkoSTLJwngdqN9kabP
E1ibDdSuRUKh21ahVwNAjxJdmc4kzTtf1ePqECEm7b0LV6IKLEQPagx5HNpT97Hc
JCurlTy8+5Za5Y4MWGx6ZkPR2MPSMXPJ9ntr4E5NRmG57xN1J5n6qWlktc2A05IX
mb85sY3xYyYaI+xGk7cp1l5cQsYysK8aMP8TkLdO1MsrGOD04gDLZIWfULqYVi+t
083NS6MkV/pJnecDgqh8wMjViN/egiCE8YKNFCAvyrMjcNJ1UCODL+xvBP+0JMdZ
V3GMqgJ7T9Bgmr6CRuw4n6NndRbDhnDvjZXMyUpr9f1EI1PYzkrLWOmsZeYXTcn5
EQCOhrLE/McmfT4GId3OlfW2Btip6+qlbJ/StKxvcjcUw4aTD4pftPQHp34DCHuW
Q+oqqPXwZxoUQrMervfYTSYovknAvjb8k2mUt/1QaXSIx04T8avvjl+nysh2IT/8
YS51h0Raw8c5vNH0Uu98d6ULAf/tQOqErkMJ3m+Y+GyNfihWbDFLbwfzGbDbsjO2
+o7KAnMFTt5VOLCgeygNhlNgN9y0RjA7xies63FbiDSVIdfeZJGwa0hUa+PWeMA5
vKTKqCYs9NOrh7DYEJEOd+UyPyYVyNoc1sfqHNbvrKwOMVHiV1kg0haCjDkDoyqB
NANv0l1pQe9ubHNceZ2fis1B8yWweDlIn4jDjokIOq7AiLEdWfzZvWsmBv71f8rF
Pv3duGQq/3jGoBn3ORQFQaxbFJJiNwBnfWzrybLNOsq0NXiIYHjsTzNzYYGvNTug
67CKGFtSh4x8tBlADSEX88Tebh3yVXUosNQEMeqbN4Le1/cXAGfq6ZuTGwH2Tk3h
pk/dd7hRnPTl13UmwtyUOa3baa/xoDwD/GbGS87f5CyBN/LvTJ3sb36QJ6v1dg42
p/Rbmx3yQGo1yHoIAQjIQvDUY6yPIcjRNhhMVe0/Yc8Km6l7DmwmiMe+UZImR/of
dZwCaeumrtOoboizfnoAzgmjsyogn3QS6OdjHg0jkJ0p5LAohtTp/eMV71GR+uPz
kVpPUfTOLnFHhlzlykv0h5NEaVXq4ic0Vi8rt1eSyZ2RIBazt+qxvXuFK+3ehJDK
yIjltff1XTuX5KDzW7Qekoge1iwJnp+NlOCLqlG6qOd4+Jbqt1AmiGu/2B3FXuA4
nUWAkUjuFjAQ93Z3WQwu4GEEkZ49Qz4XstasE94k93D0yPNLRp3oq/5H6+aZMxcL
OZxOLofXt572S/yv1eGuJcsvbSqK48zwHBiTfl31shJdPLaW6n21lNtto3PYHdGj
LiAvOGOeZCF/tM0gvfaaQdRCqKVHZ8OabS9NQwE3p/4cAN+0iKU3aZqX7nSe6GBq
9ktTBNKooQO2pLqp3Hr1TiQneHkgg6oDs3CrVPZXo7ylf8h79ETsEbDPxtUpbUAW
ijrrl2sW3CzdmfcKP0/3s4//oxPKJSsFedPYsoclJRKz2dee9Gi1kL8t7RFLwFNu
pBA9Zj6fAnkmGVfYoDqY+JlKmVAsPv2o2ehol6GOhogfBnR0Roq7b5xYjlJ6wjtn
TMCzdfgKPNWIFP98IliHKNfoNECfnEZ7xILQNJRZN7jHbBMVLHxdmEVCMzUxYot3
eWpVfCrOvYLZsMqRWdN2N+vLs0aadF9pOSyGXzDWG9u9p4KgKcZFqmTBKxHiGFTl
IPmsnZTzYhuWdtAxI3zzehr6cmt4id+U78OpBmuMlNQF0tt9Sop9MIOXzFcr9VFM
dUQURH1YLNCiwFwj10hxa24ZEeeuIQhrH/Q8gGAhNPlxoHeB/b3z010j6i/Kn8nf
FDLyr1cnpRlXzljzpysMeZPefg3W6SbrgnHQxJX+lhsPdH585JPdT9m666S+NBK1
T5lrS+8kZ8NefWsEuvNDR9hyfGzJLVHpmnaEkOjnhkMM1N0zZS9HuGToaaEQ0TR+
8H3wjZh5JHWrCLwPZLDfh8EW2akRy72u3ekyJxMEb3wFYCuC6/MARmGbCzlHcdAs
MUrRSYVHaaWUYhVlOGmGkoryMyxfgMthZGWJrQBMqUQXmC296WxopF6xpHVfSciQ
Mc3znuww0Fq1Dv+NjjpyEqAuoL/qwhJZYGKpeN1a8StppEIVTyVpHkxY0UAnjk3V
1VREcFL+b2/18k7tQpF0Wg0JadwBsOSrTZ9naOXkxTqbjkthfiZZU6VodcZbZ59m
teqLZeJ/7Jn4HnLmBYetRa9m7NkD2nyKxc+dzA6QT4FOiSdp7FnTJ5LHAMsb4c/K
OrQDPjNfsWaIDXU17z12GYuTCYwoJXKLC+C0ZZKz86N70Qvts+855J32ZjS4E/Ih
mJlAkbSKTXgLsZG+ZOS2Baj8InONkhscG331gUAZQsX2y1NA6/dDh4xUFCxLVTGM
f4pSHgw/nY7pxCgavI1QCxq3I2CeJCsZ8RSEAT8qSO5/Q/7VtuUEvMoHkQ0l4Vra
CKQReXka1UTVCyzfo5TiSHitkw0USWYk/R8dunJ9mH8LNeendHYUA7GMrXCOKOX9
I8YdYWWc/eDncAHk3dK1IhsVxXwA0W+iI9vdcMla4RZL6CxnY2QijHdwMdP2EFEr
eJwwY8+JnAcVSv5rQmlpx4ZC2otfxuz+drJ4ydQJ5uxUAMaLNYdZhtbxUf8BxZ95
gHTDGTCUCjYMPMPQsXF5wZwk80RxpVUwIjJzSMJFxE5ea3BPlafauzbshpBkMLE6
oipVwX4U8e73LjIvGQ7wlZokykz8+smerQ8k20RBOdyLlX459aY0NBoXd/IczSVW
HzFvBJrNadE8PHB2nNVNvpU8JDQDWFpWFlCXbJliNxchGb1RoJHEEh8MlHyi3y0g
VU/UalVNDJ9hdxTuZssMBXocm9mloPwuBFH3dkuCqhkVtxTI4q8UlS5rfKitW4gg
9WWMO7MkPl+xotN/Jx4zPWDaqsw7flSS5Ql5lNeNFHsXVgzio/4xBqvmGj9fcyG8
7A416MtN28oQWsFMLv/fyWUUCv5UMRvdDL+2/at92vKJ8dEpYuayFiJEskNrurCk
MQWxEpdd/006ZoJYoa8CUCc9qGDibJD2JPEvSlmi0AMH7siQFHit89xRYYFWeiJj
7LET0GbzgdTMfY0MA+18aZCAgadeT5xn86/4KE9hkylbQa6iMnj9VARzwv1yiwoI
ifQjodwVnDhkDrztHRraeAzcNdPDjXFSVh/baaXyU4LJ2ZZAaNUwKI1Yo6ojjknx
HvlWVjhlH0njx506v4Q4fvJVsRMvClwEerTXfxheZGyNGhG134a+xQBOvcua0vdh
vejep8046OoQfM9UlBQgot83hDKQjU5A6MLOyF7uZiAI9CKsem5RanufcA0cosET
wnZVsL/T20+DJirwKgfm8VORnRy3Mzg8KfHuHgqpYIbp4k1cg6BFsOv4LM1aYCJ6
4TiLR6FbGPo06Mz6j6ivrXMroSdd2LRM9umLl+28GEyzkdOiRbnlsR4bG2YZxtvg
SSxSBGXe87UfMJJvLy+AQoQltPBr5aQ6hWhdoqYP9xfSJcPgLbUxXPbW/rMEdP8i
vQWN9OlhlVczJpT+rLbnO+YtpImZ05jmHkjywxPOg5D1Z8vGXJ700Rjpr+RfETvC
MvFsMMiHo62dhC+0CUC+JK0Y2uksXmghe4f/IhYqcv+hmGVHxcXIcf5A9+6sOueB
+mf5TOWpTyU/dVeaWhASNIRDoUIUIp9OTNtmUWKFeWQcdgZ7qgTkeEbWQ1rOOZY3
1lNz8reZQvEzqhoDgUD2NjkHFy8x/6ZJxMuNBbNh4XrgWp/+HQRZDuXOaJnMbIJn
h4JNUrU9UE/SQxgn752dwzC0K2wO3JuoizN6w2HbaDl54Y82RIlKtjzaZ4U3DjRj
vx8mq9OwzvVuplwgWAUcu6nb+POS1FGsfaZM0bLo34S9sYCoG2cUD0ALn7gCqgdt
maIqvLH8swOcRwf97kpka8cZCUFO2wI95knL9XwjHvOzIC1bGVowddPhtJ6s7381
9VqquRx73niYIz0ZxjYvG9kx6uuPMlBw8WjVBbwCdAAwIVXV5xDBmtqFzA6b1im7
Jn8vf1CWGef19xraIxIjk7BJUFHhPR98u/G3YoIbwjfLfZVYBi1z3POsA/dGqYJN
i1kGGgd3ytO/N22ISdx6kS+iwou03D6ABRuNz3SczgSeECufTEfTH5pmFeURa+iu
5SIxda40sUeHbfGFQOfsZnr6cWVQfv7vj73OakOPzWCMCzYxCW9yEYeuFWctgfV/
iEjFfifvl+dijPuSfSkXwsSu1treV2fMrI7W43xYyIzKOrid42YIOhOFVTvqx/xM
BcH9VYc5E7Vzufc8NTkizPxb84GT9Zvr4eMg1zOtAmGyRLvuXp5UaEhErvSjUe/+
FtAKHkZctnOgt+hvsSlmlr3iKQrn1T7A7/k+93cADGHxPjxROLA4jzj6YIi/96XC
Nh2Oe/zFwu1gUpbZ5zu6CO4CHDfj/4KhIRFbaUEKtEfVN4NZQAoCh1857acDMOdB
opSL5YNvlB+4CXz8Eaov3t5asc/AVkMxOpqBcR7fgbQ+7RjPfxzghDqD2SpQAyfx
MxrOkE+eT9GB9jrlUSFLBh02y5Xa++phGvaRobmr+Ek82CvOQ3sNa4gGeo5tDVOA
6c42YyjutssWYLtKMrBvc7ykgrqoCd7yV/7ys70/5MuNX9h8n5U3+TAgj5DrNAhg
MzKESFVKveEtuEXtbZBTPs53CSUSuCFmDUw0JYovkDDFq61zTvsbpWACQ3vZ9UiY
hf1KbFCol5gqMamYUVODwTEMyq6RzInstBSKgt3p1WMm6cvyJqHO5BZGkr3NQT9f
Lnr4VcXYfHauoqG5KbI90NsWR1lk5Wb/oCddO66hPCQAjmYTdh4ISqEtzNKGohLO
7/BswuEVQYlOebvmd3nOZHiFyuKzP3aDmkGvt0n+8Bbk/k0RGZTvIWQ8PTkhpA4N
x3rgX9u88Mj0jHnXGMfwnsuHMdRJvJr1w2/MhVzyE7ZuZQIPr576SYDqCRx2nUzX
LQqmKTKO2jd11YyjFYCJm/iV0zU2v2ToLcfpebOyp/EdFaskvSJPyW3iJGf0SbpM
OsA/foo0IqTnH+z/viwzTljT0fokaiYbsaLcBvMl6+ytYVFbBUGecDJWJTm262YP
e4MagzNXn/i6nZ38c1W6ZAWaby5F9aEa5sf+dFvTMfHNkDmsdEVbPn0iRL4I6JOG
/Ge+oB+WM+/k+73jjiksVXuZe1zQiX5UXizRpV1V7rCz3fhZKbASJn+Ql+RakOx9
bjMAFDqxuizYPqGIgSfBzkCZ0BrObYj8MggKIOiK6faExXYGMLs/+bhexB/IUdq1
bqSXdOsEAsgzDsYEAWZwe5NyVwAn+QPuOPUUnrFuwga+p/Iq/olUjwlVZ4Mxe3t0
LLdUSTZUQcBqziPVL54Qe0kS5J/K5weR2bBPNLs7052HsIaKTSqpb61iatWdamXX
HoeS3DMWQGXN4ug+FIuqs6EHisjQC05KaRXHsGeaAOuXGlf/qbFgwJJtt1gSMeN1
XxDCDxt/dDASwbtebQEWwOWXASBIeZ/6wn8QjkEQpYl7R7iaTpQjdSYBV3oJpH+s
rbDD8nvBA7LduI79qye7mg/JWXg48FbOsunNCgTMu1ErWpnlaWRoHg83SVwqqND5
127Evi780H8PCQLsBiXZnK3x/L8B+Q0lZgqPdAqpH4s/SoNTTcBPPWvRzIWhw/kq
wxCnCwhud0CeYweZ0nRUZeoaDFTtk813nmZtdskQmGGoWvwkQ0dLt4M+p1iOh2Jo
OZa8QoKrAETK2jdQ8lPHuKHxdOUF8P1SCtooJPD1An6AM4h53L0JzJNsocKO5ods
Z24BekINIQt6FMxDSyquM3lgcWLufdGjoM7EywTfOY7LUas9QT9QbGN59rL7cgin
XjBVWcSovSxNNslyHQqrXcfE/71QnBczTmHRj4tx4v2l2GDnzjPx+MFN7DY7WCrQ
0UbRpi6cA4xE5xVUv2BHeFqOhyWMFX13Ge2GRLUYk/W55Ik5US0fKEz+FXIkNpzf
YqyfWXXFXzHNIA4Punh+RtiUQtDBiK0regjOr1Vupk55ZzjunebPNp5+l+w/Omuh
VlhRZMmfJoZDtrQl7iWVUXobrqJutCxoIxikPQk5+LAll2+C5NlxAQKTkImw8iIp
fA6D1hHfs7+8Ofwu7jXSjA3cepXtgdU5mwcuacdfq5iANzU342ZX/vbqDIJdVvvT
f67mYvk6XjaSDLcWSetDteFe9/cZpOZ+OXZ5PgxUqAwKVDpP/6OrbIsLa5vIjN+F
SCZKYDmdF1uIGtxWcmhz6TljcrbO8goF7n0xB9Gvb5xaVf/XQXHvfOeI6Y3ebzjA
rWbP5mP0fr5D7KqnKXiLCFRNxpDVp1jH6ZSsUhmc8kv1F0pxWY99+D9b4RtxDA02
xFuqZn/sZALYC08kUwGGcG9UxgT1RwsJFaW1RtjQqemXKzKELl4WLTIfw1Y4EwYO
KgkHtbMM0nXt4C9HbOglgXjt/N7f8Ej6H+Fqx9Ret6y2n66Fpp/8kHGrrbVkJFvg
oVfBUvcLEUyjERoiqrUfN5T0Ni5YSDNRpXb8wpCaAPgwMF5TwInYmBlXiqCA+cPu
OX4v7ygg37hiWdpgJY4s8wH7v0204BjXlSj7e04+Y11fQ+g4YH8qYikg2Q9kHxrq
cIpMkSL3hlAXlFCKViU3KYVSoFDLkzHC8AdzBBtcjqiZji3P0K9uX0CQymHldmbh
0RBBGFgg4UJWarCyr6wZMPcuRY6cwaoxHaIWte+5MR3UrzPVK0HwtoYZneyzecKz
Wm3OdR3SX1hF/Yzoyr/DG8AM/A/ENYzoKZWuULLFxo0Bj6MaMQTvuA3jBrMp1o2g
GvnZt9RbdVUwJtAPopntPCTr7FDEcG75UGF137F9EfjnV4HhrO4q3dleYY1yVtWe
yzsGEdtw5CWHL9OsQbY5SUHhC9Lk4Fd5OaERH4RfAz9oh89/u4gLVb9JvZRda9d0
SA1E4lUJFSTEsosX/sPyeb1wPA/6oYrxel0pgsi7znts/0mYn1ZXqUHNnrY6Ybql
/P78UrY7o05XtbBKJ1YM7Tt5/DK0+vRjI9dsFBNRCY0GQdwW1eVdbCtgjsCi0Th+
f21jaBEuC9tflBOHH0HJcekDIffqLkd8FFVYVYNtHZUwPwWL5NTF998pyRX8yO5C
yfrRhr5Aa0ca6GGHfCCdY+UQHcTuj3KBJuUEsfZSpWkJ7ICgA+rzKD/sVwHsA2nv
ZRFAmLnoion12MT3OO+BfXjxSf1MQj6+90QVBRQWFlaDeQE+aVWCmpy4iZi5F7Jr
M79/yUnoqM2Ho2BOpLGv+oyTPY4SXyrEXdLJCrGO0MLVRH4pz2RmUjU5MOzTlXX6
xkZ9ATEClfwnDPJ1hVakD/EGRYin+jMtdju8b0/a1PnXEKM/ZLGDcrhSY+fU42Br
487ZLKpBzsEETGI4BmuKsib96xhSIfhBpfZ7bVnFyZtbYUX1EUExgbPj9a7fNTRL
MEVbrzHvnreVeIDcjMprwqGkutiWVGugC2/95bRHhE2Abgq7FBsPBJJtnKpwdhfm
M5MGqhuP2IfIawD5wGgWxMpMV0r3KZ8MLMEPw16FNzsA8nWonE7UESTTY6hBHIK3
JBhYwfPT2zla/HmXhUY2g0glOx4wYfS4EGX5QDc1PfIohWrRMlnIBUav3Aq2/J5S
ia3fanbbOuB1591O8aHVaxETs7o0x2bnCvPGIfsYeHET6HUTbGBpZSI8Qd3pdlQu
Urns6UANBrfhFROVD1So7HVqiKgQKGstbSIn6Rvjn47oDo2fr6b3SBYn0ALu/XZp
ZCg3MPPECtRN4YtwVkAPhvs1dsqZci4XC+Q56HU05uXYbY3P+q4Mh6YKAgO+zbQh
pmicPSHjDhnpxZE5p8DSlaujsdv3IQZzVky8l6nUdUgfijO2cJw8bb6J9gMIVjWz
oLB77Q3y2jTToa2A7JADX6NHngsqRZHUsiLunnVao2uzIfNGgCK6o+V0Ybud4zmJ
3ucvTbGFBvVzdkrtICIGFfIl5EorwZ2zyhrQIc3K7LxAoDtsdYrOqbEuIhMgxu/A
/llQ94nljG64nGz8QjjvMD2FRQvoS1mq0PFmn9sanXv968KTS+CFnDhT2eZUDO7R
G6UR9JiMFwrASiMLxsWIIy9xPv42ferF8MguYkhdoF9ctPg305KTdXOx3YEd4Dlz
bN+YeUbZ3qwEykk0TcWPjX1HdFAlItEkxndVVYkyUdcQj1wyd8b+g+LA+EVAOvlV
KQtvF8gecVYacDy1qc8RujqNKF1kLXld8JqLXxMNWeT9es+QvoBFC3DVARmkUz53
rmyNER6io8L5vUeg/u6fyKN/4FAtCQ9r7a29aPyGKfC2YMF8hPdKv6E6PCVQLcUc
Zk8BM0YkrBWuFvpAGri9gxYbf8qpH2S4IaWSDlqstPOL0B7jJtnHngEU0ipuC1Od
6HhLEpHOo0CO0c3phzDKXqznHBCcunTDtz++DYtCuJqgjBktuzyphKkBnKkTBYBv
ZxC4vFR3bFCZuYJtvEOCz7yNvzwqZYeeGm76qxc6YGseh2gWecgVB+jRxyb9vLau
QxncsCrQgKG+h+g9wrnwOjN1xUQskPQ1MSAJs+5/0QFCjNgbEFqAVbp/jN5yBIGs
8jpQjtfaOgS6uV/i158h778qlrY0C8OFLWxfAHZqVzwY8hvIfYBeYJrDDs2BMfHU
laDSG+zlbR0Lib7BtLxJYcQnre8Ehb4XhxcOgYQE5sAczZjg13vdNZhuOzhPufJq
z5O02rOh11mR9W9qz2Pueliyi/iiGg2dyoGrHU5I8qwW2g1Z7xCMfMmY1JZoYNih
NRl1OT1G7PqM/3BvSfvBZcNU4jd6G9dJiq89J2/eL0rc0gK3mwaA6kMJvEuaqBiF
LVzpUHRy5ie1wtF0qBl6f+s9YxK9tyxmB/SacgcE1E0Rtmyc5PDmFuB3PIxEzJie
Gs+5MhCtDio7UL2+PhbTJ+kBANBgY2l2gfC2bzdt9VXuSKIIf3foTg0SAMYJ2gGF
+5T6rj0/1bmS/NxoZU04TsHFTnVnFJiJC36WrE+SoVl2enH85cajRbl4mJFgfEso
uCegq3qHx9VsicB3vxI7Z/30Mt1nsKBIVE+ZwZU3xMeUyHRIB5dzGGZwEyNgmBK0
Qz4Fx/5ZTYJ+Iue0HrT4DIM+uo1zezO2I/vwrgtxPJEFhqo2uyslCnAJnaqNd/qk
IWfuROtXJUeMkFNvAV9iIPOUF+yjpq6GnD8e5bx+ANSwGdrMpX9YYehQr9FJAibB
Fc1neG/GhLQsSWFfb446ruRyntaLpOSz2yTlrWeOrfjms1VEMCUqvLcvIEAkYdkW
RTu9fp4GkkSfmoXVSCTEiJiPQL7351qnD8njzy68Dcq503dTgAvG791m1MSiSi4V
WVD9v8ecEbme2rt/a9aPIXZLAahdrhZ0Cm9c/CdK8e1fNLfV8KRqw58LnZ9/P1OL
GhmkW0QHEksSzTEHKnqsjU9T+ej0w3w4eA0IAfirPuq/iE5+epQcLjdosPC8FNmZ
XsH5OGOjFR8EslWkFi0jpDknX+BN4UB2WN9KP0xm11bXxX+cTDbhyQ9xiJ74STqX
gRO3pu7WVXNY//QoVggqUYprW4dhKPgb0p8bySsg03PX//SU6OA8YLyT889v/yGl
OTc4UyRPSF230xsaEo9Ud773ebqCVEcAg9qJKxMLv9n4evglQBOykDYSzYdwF6bZ
nRy1+X8DRHb6IthLoJO0nKScjcYbsV59CzEcTDuAN1UcQdbul/YQPsdxn7fKkgeY
6c+9NMmDhvdBOJUcYUpfyQaRLwEadNsP/Y/IJ7jXdzNljnC3ewuz6fHInxayY3Ga
SuKBO2Fuumonj+LCEWmQGCBAMkfI/ccJVuc1W4XkHCAMr1Lwhl8kWXT+ZiX09Vx2
yX+5vQfMTfwrjizD3ze4IgEtuQWNsdjWGpwciRAb5duXUCQjr3BU8n/0YZjYVAO+
ZFMb42d5R45L28Bxc7Uc9pn8eLltN6pqtmvhqw6SDc/m3ehHTg4T+mLewEp6J5O1
qaSXbNRcpspwKsO/MW93GRw9pzP9JLxBLGbO9bJMeQjN9eeVLKXqH1QuTWXUk+f/
KGFRt1J7F9BwJMaQTlpq2P3KIAGZDWdEgZox3L5eNHg2gYoVCqRwcV0DJOkw6jnw
vBMk7hK3hdQyUPR8DRwsoEMFqBtx1/uegbFkvg52Ks3bKm2gNaICOkfCUOR6mTzo
Fs3KFcJZdV+Zvb0LKhlCsMrYshjA7WGDzz1csnocKaCPktGp9xoovfYREhiE7ULP
RAa2T2ssATsblGXsxeQM06varI4j6gEqWaLTOh1RkZwzMnjTbJ8zX/7ezHDVrroa
kOzBHK5aeTy8u1FPq4mFS8eaSIAeq1vSpQZfPK6hTNpOVTYDcL9EDKLf5Ps0Hvcl
GMRh8Oyuv0bzJdPVJX7RlCJjHp5XuH3DReMNVlaXwAfnjtQDfK7uXUgdUOKNfrDz
nlAD/S/q9ek9585fkQb3ECvivnKm7BEjsga+ImnaB1VWXsrHtOSPFZ0ItDjQ9nsT
lPIrjXmr4X7wEH7uQLflrh7PEfjpqCYKBhAb8cpOgbbFxw9OYgPyXsiAnCOa1MKu
HWihEDJsXRwWok1mfQ+zepdF330TdjmQdp/aYlw6LcInekAyLq0c8wbMi6bRWjkO
lepmEnUQv9HPl82bDsMqL2j296QtVMPvUEWMZvfBzUgEB/dbmbDMsDYqXDptLkt6
cetigTHXFvHkmlX4L7Ap6otUvpyQQKL82XbkCOhc6o6nuCJTg6hfoM2Q9AbLCYNr
r4v/7WjkGY4gX5zecSzAbIVoR7icL9oMxFhc3TeHAxLrLdImFDg4HsfBxhmahTSr
YMN4MTKORkrFtXa/r9hJYeS+grjSvTzTbNkLciQsj0A4lGcvPg4iRGF+U12KAXEa
gxFLImYua3z52JAnGbKioS5jI3e71fM94xYwh4CnPtAlCo/5SJT+An97zy35lmFY
cSb4zNkrXlTZFiQ4VAnBlPhJsxnmVxqxyttMG2zdubLskGP0rYprm1ftGeTEFgrs
4imfdDY4TA8VnvVXtYuepEHmWTtzVA/aypEvMzjGske4f1NCE475yj93+1Ifhiny
rGpl84UlSGlhqJUP3nl30uPEvcTVofeOI5+4vO3U7e20u6wC08gzFwgbQ7u+pGF8
97F9cDSeQPF/B4/zCZmkKQ7spSZSgs7Qd57TcQHtUa4X/fiD8hU4gmGnFc66EB9P
7G3RnCfXZ3nag0mROzxTLYHhMOnWhaviFdCjH6NF61qfqyjcpsdNn3a7xG9SFq3Y
/YfavSaR17Ws01rlVlaoKNxmDbDIHhu7N2uUBQd569qmljwNuvZbYXtFb3x4EyRW
25DCg/WTy9003ynuPhe6Gd71h1P55d6MeHlAdbh/eankWS+XS7/FDGPIVb36bGpn
6q/7Y0Fl1WnxZjknzKqOXj0Y3BvxY2lrLuM8ubjmVVRNYMuAfmk2AmvendC+Ysov
gx8EXY1WrhdtBs41dWPzxGpWmoJZG6dInKDvwaP6aoPh2RHxf2MZmJUf1idACFOW
MN/aSkD85VrB9DGDIhYiVXJYJxeARDHkZtjXTL4rneerjhm3tDkdk94jUzbjAeI+
2jkLRA1D2us/lDHEMSXk16XDtjIN7FvUaO77v9/Jg0PMNl1XHsHOQrUb9E+GQaA9
rdLd/C6mD+vT/tdkKJiceJz5kG7EdPLERURS4lbcQE2/Gk8Rg6Ur2GrL/BIy330k
jtf+hIet19ViuiOdWlTW1Ei+xET69iTiWP6Oz33ZqSzlhL9Aw10YZupdminCUh2E
Sntpp8THeSbvpEBtNKm+Q2W3EBYhr/8JebIpYHH/wYXrI2g+J8M430XKxe7+yjYM
OK8G3hyB4CkU526k/s6OZjl07eED8JlxAFnIgYnARlv3CdTade6EytwcW1gnOGL3
S6iQKjL2dI1G7JOA6jG+kTuJVkeYG9gmoWEjuPfBHbgzb5eIk/M6xvrA34aY1rwe
zO63xyjQAN6vPJ4G96xyk/7wugcxtPw+9Vw+eMEZ101zorQdxwD2hIkmTokpZ1/m
KcNP30+rrFhul4xkjIoDqBpfEtsp8DKzmxCtkfVkbtwmRr/Fsaxi9ovBH9dZtHn9
/hxOA+eHXuDfqFKvlj6fTyqePE/3X8DRkK8bpOLQfNo6ZSAVgb7xggnMgTaTWH1R
h6Z7AKYXTZVCYfT6DMyf0goxGqbUW+YMGbnQHBu3+dhT4DgZWDFkkVX8zLdwhR/7
n7v/eywh8bH/2PzKzWEjPjIMxU9ENLfb9vT1/YR9e53XaaSSuF4Mq7QyoMJH5BaU
w7TWDG6hJtudYxMp1lM+TLUB6JiLza6AU3C6qtpDoN6pqmRw+Xr/arz6yix+k4v4
zWs3H5Y7eFvPj8XWga7oFFL18DIzZCoRB6f9jxrimBBg8BFBgiGVrzXMiyh8Q7g9
UDHHu5dOR18z96xqel/9GT2X+6JCXqDykiOGU1fizuu+QaVD9pqxsIv1iurUtvmu
eas9H6qZOZ9FWqjlUXcQK4m2FrRlhJEBxVDAPw1EF9k1LCAy3V+B3mVZao+k6EOh
QNHMcK4KYQYbEqxmz6YuSg1h3CZRVOHo4Uz+1qN997wGDaChYJsaMrLyAQhoEf+K
+iPmnwXxVONUs2I8r9RE2wyofqRG7OhClLivJ5zuQuqN7RUByfbEOZWnFzx3N5es
n8p9j4Cla23xnQtCwewuiLMr4TKVPQv/TG4ktk/4UgqX+odCHROKYYSxmMGVzOSu
3p15ohjFUKCxOebMm0cHB/+USB513yrzmKkBDsSE7Ew90NosDCW+/6tXTYxMvoeZ
carPRx2U0peW8LVB53uJCfi9HXclifMX2vAeaCJn4aO0dOtEy7SY3aPiK3afphPL
L57BhfQzntxGYWntaKIHt/w5nSZjAE8SnNRY5YnJny4s/KSZuuu7XQxbtitPQ9kt
JiZznKOX7+bSaeDel+ERKtlNhnxRC6XHt7+VMqblWeXRf0DlD4Z3OUjjxu/+HT/A
XbjogewVlRdzLvqfjrqfkWt7X2YxJ1tKWk1Isw/kCgc6z/FM5J2VJwm9j0i5H/Rc
WdLctrpXNvLykuuey7+77/G7ecUvhMa57qtAUc7F6Wz+RL9bf9Y7z9pqAFxzbm+7
J5HI0sWeY+MAcEYzwe+qiQP/uPM213M30loOP/43WrAVCpcwe5ugQ041z/qx1pVI
7gQAUYF8etmhGMsqrxmi/aw6GkR2UAwHbMszEvI99vc14zhbCKVyx1BzzO7rdZjW
ThNMtNSpDO2RWRBSSakIqvqu9heavtOZVOOD87zTGh1MMT177GyyYPJoSEolBwRQ
aegCHDHsnLoyN32bdWP7nEqOh1uGoA20Tw9iwF2EIGJ24cxm9VbxhJxP+sh7koN7
HlbcPs4V3StFPkeBtzMRaaGfNO1O/ENbm+h+BbypxL1KIraw+8Ta8RpPSPp56R+D
4h+T3U/nIuifHizwtb66EZS/zXM2cZENI2ClvUWEMQSku/p/r5x22vEe0OiInlYy
3VKCSo5ZmTkxP4RzdBbSIwicKoR2YwhiQ64iDK7DW2LiR/Gn9fa2AOLT9w+0MmxF
CidApn5kMGkQ1BXwN4daMUcv4ytvRlWX9zHqyJNUjmqzfvPOH0rKb1jzDS57QBob
LlTheyyB9+B9oczG4FvQVjOWRT27A2HPZCEzI8mxYHejI+SlmbGo6xVv0qg6uJpE
4mLlFuTtmMuifLYXzW5hy6fhyN66Hzvhz7MiV+dmuYwo7XWmRiUJZPVE3BIQirC9
w27c3KnPFEzmM3hpEqzl555gtJ4HjDxrWJDQyKxCIF4HhYCTr9wcOWBIj8RryfRe
fcRwLOaALpToogOingVUQ2rSRmmRtZzJWb5Joy71i7rFpW7EWYdoMyUMOw9THnzm
rDFkLpdTrfe9YePJJN0tTppwfU0bc1jLd972rzbnrjANYlIbAHVUaLpDTgWFEgbC
wiRh/a2RPMsYfTjShHMCoXtK/Ks25kDLduMwEMA4qllvX/4lSKWAYOBolIK6YJXP
UmJOHhDw2xAFOd6gIcrvLJwLt3CyumWyfduVFZYTMb7nDy20HAlwe/eAPTWRtE5L
MDuZwbL6W5R4YjwHg/Xi0n6KGA2GSXAljOjnDBy+EywAFGoZfIIoDp6rTuEO4LII
E8Ay9g/PurlEoMR2B34/S/23MkjKz7uUj7yTdn3EpH/DS+DEQm85EXbwu2/YgoW/
lBFwCAWomtu+N8td8LMr5zpsd6C9Ze7SUE3ZwuhGUu0b4Y1RtFJZwuALJaSkuetY
pMhOiLzG3IXpW0nKodCKZd6n1qNxeqfjb0O9NRziUL4sW8iDsKJ4tEV0wagJeLZj
2B2SFMO3cnyeEB33n+BnjdgWnA3YJaiicy9F8Pev5a65Mu8jv5Hxwj6tyD/4NIIH
2a0I0omzDUqm0g9SmkMO8+zC/jL04Y6sBig2KY6EiRqaCu4Vs5xEp/O6P5nB+bfb
dxyVGhLyWPjOlddXLmNTbgQEgqj8VPESTRXaFglLU7/tnnyxrc0jOj6u2gJj6QVy
cv6hj4MA+S3uUOR1OXDC9JdHsSdypcbRAYR/QK7v6SjXlyqbelf3B2IL4dnb7+yZ
YdHI6OfCB5TvmgLlpaj3mOtajji59wxTo2pu+Rb3pyZ/T6yep/uFuxaGeeRGJqjp
d06XROcW/WyYcZ8QXE7t3Bl9WYZxSvHPNlINTYGYd5bGZAjoz7J+4eJnjYzucPDK
bZ4YfkCfg5qVysK/VuLkqzJX1P480PAek/XP0W3ohCK5LvpVodwguc86YKu7FUAZ
95JXaZHidtWm8xGhHkVThUFmBZt40Nei94tQttGyJW0lMhmOCTVTzuUVBNUeJHFM
8eIPKpTIveAl0IZbekHiaqCzxaUgodzF0k2FLxfRIi07v3VmFAvVmjMcnV6OM4Oa
zt9EPEedu8VjR6yD5wjgpFBTufX1tdfDjQ+JyAX/Wu1m4oYiRYih14R6UapWA9yA
fSwJU4v6Q7LEZeQn3+0j43aKUzSqW50IiHt9G5geJ5tEpRv6Kxlx3whHhMFQlSAd
a0Cg9hJ8llRs1nWFoI8+9utgo2JDdxElqFtODKENORLzlGYzK7uMY4oPmeCRbk1m
oT3JG2Ua1jrXL776lY6UVVbmQsxVQVSTlxw7/ukQ+3lu/HftCOJyGmqUY+bdcH9Z
nG+17Ks7p7cjh6VDPntMdgLYUD0GiUEYxIkJX4r8Z8HytvxAAH9N2VxsdYqY0Vla
ncmDycxeazR/1WATu7Js/wXuwufOeregAWfLi3paWymM8TbajT4dbLnrHVVQWzV1
v8cUBEUgOJxovf6+fxD0ct8TCfegtCanusYPI0kYWPNnU1VQDmnbTLIfpKhG1lov
S5l/TSAT57IOSAbQVYBMO6qSDdu6DO5QBY91uYD4clR6SKWTVCkVPjOjjxdQMKco
wAmeiG2Eoue/yStxkdIZzFoVI8PAW0ptymeIsaY7sBnocEtw/ySARz7h9ax9L2xB
IOeKiKSQnQNwtJTc/Atyi2uo0Q9P1rQ+W4iRtdqdJrrob9+CfV7yYpMjm3lvl4F5
eA/poCxMGWUOwd3fGVdJkzOxGrJ2fspvi7yvkBWXwyKYkAiKa7qhEPObx6LMKBIZ
1H8CxasXjLB0vSWdMd4uuE4eDYPjr7lXWwOO9wFYtatwUn+8bK9wNpcTMSV7jNhG
E0YygqkJEu6JTGkySsZIMBgqkoDQqLfq7fp2RVFLTpz2fKa0gSzQy1BqTMktaTiX
aXo3DYK4YXbsniEWgak/N0Do4ozKnL7o/J9cpxnytD+awmEyv8l1U6bYuL6O4Oe5
qtaPtLyxPh4ZgFht1/YEy8/T1eVD/3bGyCoVMP4nqSLoLSvsw6rYXNRX+oxx6Nkf
gJNqL6Ul+4NmHHKYxnWfBgJIJW3qfm/sejwGUCep/WeSBuekwvJZ5/DXn0D7VT9A
VfZ6+tIg2bXPmV4BFeOChizYolnVW+PEFertXcRgDxHmqMlE+Nslx705t57HZA3+
DDvfikzSHz0Msb1sBBJE/YqPLesDXer/yo5HnYhmVaRWCxvX02Lswh8xaB1JRJdb
zLhutiFXwpi7B1cz5n/wxq2kRXjre2eLuUF3bUw/0K+pxJ2bqK1E4JRuGGqG1OzQ
njuAK7qeM4YAxNmmrppTIn+ZaFyApQ5y7BG7tMdBWHkZAdEjf/bys/tUiXwS2mfa
XsLQzfeGxnCcO9+EK4TtIfl51hrH3gqZGGUkRsQQWRrMVFtw6xnW/AJIZAIAgTJC
5s9SberuZnkGIZ4CjJNT2yL/RDqypiGdKJWeHtUzCCq6v/0vdUUzPrq7rFeMxTl3
Yakjx4nPKEUAcfem73DBwbAeVs5uNi9w8Tz1FszSf5wn5SEUqHA0Hng2Wke8vb17
W5Roah9SNcBXMOKRScsw319Oex2F97R7TWLBp7wwX8DkI1ls8f62CXWxbfQGHEcr
Mz55GcUjllWeKzitMOY6frtr/jiJ01YLP36gARgMnQ+3F07fet9BUjBo7K3dB8c9
MJxiZQ+G9ihgIf391tpXSxz91g8wmlGcOUee/l/ybpopd3O0UXJcL93Hc/MFz2PJ
+G3dpPjIRkb46Rj6WWeb5uXHC7bBIhcSwlzarZqYi1IpwfNTHRf8cZe6w8UYFDtu
kieytsGCbis9QHcUkqRfoxvNEZCF/VMhmAfko4q2B8c6sZmhR39rOFnWP/5jcRD8
6pvrhBpgDxSU+I9IwQHNpV0TaPiM3vEB5H0nCdU6bHvsJH8/P1VqKFqRKL6jlXv/
TLawu9PZD7VW3YZVna1lxLAfm2UJDtgpV8uxSHbgoJ72J0CLCJhJxUlPHCUdDOwg
q896pHOupiW6PxQOXDgHSWPrN98xnDb1Zlsj5OIoMQ82rup2G0q9aNkgqe6hVdSc
UKYUIE9j873kCqCoj3NoBFqRwGAxIDKRlALxvnvNQOvlTv11gH3ds3NkWQdjAkXy
f9SKHGY8mXDt2U9PDRBrkBHCuL6brX8v8o7pikDOaMpbgypR37Kzk4NtRfzpO6pJ
pCbsJwbgC3du8XLH8pkGYScIy4etcXaO2AJeNnyC9Gbo6/yIKV3iuY2IyvNOl3KR
wolYawwj/VAZLypOgdXf9+8BdzzJG72Adx8pUCj4NGGtU6GIHQnCkLcgycv9keAN
aDGolz2kKeeUAKjKf9wV0r/lpAPCLINHsIaVZqKj2/WQ0RAHqWsgB+O8Cy+yza3e
cmyaqZm+XemiVfps1kc47JRqHe0GdgnfU2i0i4hlLAkKxFUEqc+vHYg/Ss0IqzOK
7gKUVlzrsVhREXYcOyzLggZ8I4WKnSAIt6rcc0pDpEzMDdJUA75o9uQmn2tlbigy
ZgcnySrFGpO+JQq4dTzF+n0GggD2dVZfP0oORl7EqaGKJ+LMifH/w1ltuTwqgddK
AwSzNeY6c+wwB5c5dNXNEhl/Rs4LmbGO60Iuhb9fgvapd/4blHOc7RBR1a6H/OZp
SuCTWuEm3FulFV8vF80xhekHSXzvdJUsZ+jgbHUq2nSqNozdNHbjbplED4wF1o6s
Cao4G7LH1BEW70JBCeclxwGtibSKXxTII7Z2wf3eOZg+I0qKtH6IN+isvEOgPd+F
qkM+VBBhJxEDAwfzIK6E/VA+CXIK9NfRNKUsrOma7ypXoklPo87eLNOaX0fgPsWN
nReD/kL7KakSz4p3YbLnUojgsV7YXE9lhEnBTD/mOOWbDuwiNfIrTwdaqOfTfYp3
FvQPo7UvrkMs0lTLLZGih2nIwuDguT31EySucILPiE6abLNj6FxTt8xWrB7+vqT0
dlfVPTqv2y/g3MElyocsXWMMptres2QUZEjpygrsqoBOTmMog1OhYF1obWI9/Fg/
vqwLPenCXdwfkXOBIuORL5jkq+VJj9jsupCW/RNk3g3QykWyeSgLtnsuN2hhu0HP
at2cnsqb/IjBegl/rMAEt9lfHGu2OgBHDCbaMWEKA3YCbqpx1oDFiZP6URQiIKUt
MWGhMhRH4f+kB9M39MkhiBckdcRMW4eEIN9TyGOxQ/EVXSBaY7BjgGESKPPc92G6
39TsFGnym0nBRxcSfVe+egHZGnUfKqiQ6QecKkxPlGIVrsQ/zPnWURqc31khjbL2
6j/iYZD1qdFgAXnMDbuLAKFY/Od6i9luGB24ynjCqI1NO1PrWACQfvp6NbK8SD87
l+eM9vXodVw8VY9nUCAzl4hzv3AOsyQ1Hcp4YntUoUL9Uu1w+0Y39Qyt7F3qneI3
r3HZ3HnyMPa6EaV2F7Ab+tUbkmFR2UUljC3Q9ef98x0tSrFQtcpz9gk+CSap8xx/
vkrJtB4pV5o0NYsRTHcNOds55jkot6oErQQ2ix8jR7d6Bi6WYDD/WyVSFpdgszXy
Np14fG+/filV6a7CLVuL/cjw2pOYWMpaYe1fQT4OrfT+4L9PBZRDJVpj9Sx11Qry
3jPdnULobIvf/6XJc9IYZgKGaYrXUuIxsP/ENGBHmZXkA3hthPkPzsQ+MU9i0gud
jWiQreqs9XmwI6yB2NoW3zDB/bDu8uRyu6bxDjKTDySiqWBULTMhwaJeVu4GhDnl
r/hgyFXPgwqFWsIzJTxA3gTIk2OPGGps7qSLRfQqpMzVvquTsdJUUr/OprNybYvP
LHJllqwomOdU0UuhQgngiWXfAGLE27M1m+dQqnuSKpSU9nWNarkEq3fF5zis8yvH
J1R1P8xB/X4vRKsWCcEAiLQPVXFQMRnuPsDuRDjDhYT2fdAKeapky6o8NZeHVR0A
IvtG22fbavPGS76pdnNZnp38jAoH0zDvO597kV1xVD8doRxU9k8w4QYj5L87GNk/
LXP8VfwmeMMUXTB1EURAvg6cuBheXQbqh72YY0JjeyfIXSul0gRVV+vLdHRWUmuP
m7p19MlSjnFbOreTVx4gQx0L3kIOPlykulXIWi4BPZwD6015DEDnSEz0Jr+VjgwN
aQQIRo7yActJrsVAJWwdLNnKHNs0Qq/p045dT1xi4t4bsMT7PIXSKyOexYsUecbO
ysBVHjxhauLz4Ldq0mJXn8fbPXvxyI7Sqs8zBv1E2EL+GWMf1gecB5aWAFoe2IIQ
qZlLtG6us997QHk1rpY7vt4e9vg/tUEpaivRWwgNWYSCSL3v0vlIF1lm4jvxzAKE
pNhU3xeQnxqaPIP+HSX6AdkR7wJ84YhwkCjM5njg8v9b9ABYWniDk3gplTteDz9r
aTb9UamQraYRqAmBO4DX+Zw0LNnT8w7Vd0/azoCiyeymdpbOBvQfPa2y78Pfp320
FHGl0jSF3jnOpMgz0w8hf0Y8JibXScx0m4OIYoaJXkox5xEr8rBMUPnNWKVry88N
Fdf8RdvPIBDiSAuEoxX16EilLSh6nARskaTa4vfTSdFI9+AY4nLJrsVFwNGZOOeV
ke17X6CSFNUVmIofYuxVDH+VImuxps00MxkcsrlrmN8cxtkqCI/VGdjIYc2CEIxV
pIQBNKZzYXCIdde4O2JeZlo6BgXt4vRmnKfhx0H2pFALXB+woUXJu7QHc9JCu1g1
0sWb07w/Km9ShUsAPrFlj67Tf76kTnAzVFHU521CaKyq1/QNgEPv5ZyJVVczlc0y
vvo3OOGiGTlns15vv9saG9eyP23TgjcTm49SrG0z3lZrKniaTGxvB/+k1HF9g4Ke
yoTlK5zic2YQErdGvXtqd+SQWSIldNLNBt1cO6DerneEvLpKUce8GHqq7Aizuk/j
MeMp2Q/aYgv959ia8wXdKFLW8Y2KeS2sWUagBdQkDDhWsfXr3GkqkbgQTayvRDbj
tkBsYiFQDH6gI7XpJgQAK+34e3rPw1ak+/LmRMH1dY4SWUGvTvNFIWcIxynN8kPY
UkX+codMR50L2GUDJliv9WlJPRRM8vgaKG3uqXTsxXOLVBCM5STr+XwS+eBCtm1Q
VNUnzE8b60+M8rHkEEhyKct5bqKkbZ02XPenKf5UK19dnP+ljdRNwxZ+HczYzA49
6rhIbf0lz9Nefc2KtJhE/DwR2a7m1alGEJ/Q0Ior1efHJGPObZ7SqN0H13fWyY22
HD3viEisYHplMQeUpeggQ+FtRe3kS5k2soCxsomdZ82kbQNjHXbfZfyJik4JeT7f
hixvFexqp4MendEnbRiANEFuf7h43m9RVUuu+EkFbZRfxwff7FTGODlaPqNAidXD
W8L/BpUvuwE/+CX0RduJOd5G61eNfualU5l9gD2rx+AkmWWcig+QwwqVWx2iIAiP
BW6dktzRukabZC3eCXCb0MiiBm9WlQZrDzi/WKHI2pSaDhfBKxUYjP1/PTGfvrD5
6v/oGRwoJTDtcECK85m6q14gUYD9OJfNmJDhNktdFTDOa0ZizRDAifVbThfEYSlv
JICO13ToYlvdne6Y6EL7JDs751MHb+5L6lR573nHpZg+xstbyHQItt5+YnLTDp/r
IdwG8JgjaiZWnZeCm4k/lG68w4OTfg3V9ykdZMoOmRisD9wlc5c+0oa5zOk6s8Kc
PIMTghcTqFJGr5vZ0ILsN3jAAl1pWTMcP70h7l3aT97ceeXPo2e4jgcTPP6DtXDT
7QQyZqQjYAOY5FSzCree/WrNFBNJ04uwpLSp2VAose5lx0FN7wFXng5EedHsUu3S
oZYzpjjOS1z6+JV2laGxqZ1rTo/+XK8LuGCkg12OM5WF6bzuvZd48riuAnXC7aH2
ukH41CQzyNVwKPSA3LR6DsjsYpiuSTxKbDjow2ipQHSoueb94kB8TejOCOfQv+Ig
/WOYKVWAb3vSDS+7XnHPaLyNYvkR7iV18WpqDlEcxg4zkPYbOj/oRp+L4RnDsF65
yLovFv2q2c3AyY+T5xRRSD2GBAsRW4RoYgZINZncfuvwF/uJcReigWO9WBvJWdXM
6lqokJ8gR9n+4FOnju1gNECCM0tAItLnyXnF18eE+KJrZYsnEYaobqeI6i173nQ+
DQRrrjJyTDsxwQ41J2IPiX3xgBslvd5q/IulSGaf0l5kgp0MaNkNfy944eYHItMa
meFB5DUMXHbRA3dJRqsuSyjn3+OpI9N6q7FxMHvnDk01lXnqzPGYoprJyXVNJoBT
c3hzVwkCnKTlLc1mJRdktm7pljLNgDOsX7QWSRoXdv7uVZvqvObH2SAE6jeFiw3i
MJazJPU3bTAKwhkBCduJF7Z2t2tbogicjUCpFO4l7lNBMgylN8GylqKmFC54YSPU
BrGQhVIMB5q4pyOPiPe1xvqSvybcn5FwrO+nb/ero8cxcGOjCER0kp2rNaWsUytv
duqN0vOcNDXXZfT+ZaL1zYMfByX9D53k+rxwvc6ZlALHQUKzXw8kGW6zQfGS5v+Y
Rziz+hQWuf8nMPhGiyI2tYSuefaQwVZpkdm6pJFayFCPRwnIbE54Y5QA/5ywc0cK
D6Ot8AYn7i89NpMeLLNm15GEGN1WPMlHEPhzW48KqkVO3gAZCe2fVV2gIJGBSTbW
mHFGJgkWXD3j3KQNZWN87DOgwABjU4m0DsVG5y0kpvFAqk0kpbFs3ugXJX7QhMUo
L/jbmGUe9e+DLrVIZidnowUksJ4t+iK10s48fzP1qaqx8uE/Jn7Ean2rjEfXjzKZ
6n4fCwqo34WQ1RXYOu8BKIr7z1zlrQ1hb8XPTMlXBJQMCwqod840zN4sbMKFfAjm
jdOrnfO1PmR9lGQ/dvlbqZUVvNfFtO3NlRGlK0/WdOiglbNIqykXlsDtm35wkQbh
9mc4Fxp9aMGopzmH5XLqHw4DMDVq0s/89ghjKvpXDogMNAF61hbueCESrwmn8zgu
Nru2ZMrX9PreUWQx56VgCU8IRZNftG20pq+NaDaHEsA01W+fFgc0YEyGkCFKhVUm
ZwhSQ5LPLRL42PlPvzL3H5RfGqSi38Qaev7sTTZusYkpjaK/afoSkGGnc7Qb02GF
T+tzsM07ye8OqE+W0xjbY1p857s7492O+psI5B5M/teBog9MlTu5561Fy4Q5WBQU
lhzyPdwZfAi3teBQPtwnLoE2SYbfIuxStJyJuLcQHmz8BkwbmJP44R83HF7x73ZS
ATBhi86Vp2lodtWGWpFvgt+unR5mIKX9I68JKsFkeig+YdmVi0e+G9h9UG8fyFu5
VpEcOxzgnc+NyIYg6vWXfKONxWh2VOcedFtCLBgML/9JiCQGQ/ydBrzodWHHeCl7
HhefCikD7nYZmwEDLpwB6xg5jT0IFNAW5mu/bXhIPfE7T7pNzXZbI8wy2JwkaWcq
V8Z4ej3HX+swLbXVopL8LHmLZsZYIROp7NVXtNf7Q2Kystyf6rD7sKSYU/V/9v17
DPsRvPLqiFHpZoOrsC0xNFAeDe4nzmtCABB1RqDyqXWUsvQvC2AUEh4sIpMyYpLE
681Y5DwWjci1KH+rCPkju/pPLH/MK+0bTblCHWLHnuWvg80w+CQsojqsIlkORcqC
OffWl1DLEcYBIyNAIn4FkbPl6ma76g6IB07ZsdDcEVa0mdIuePUE2pZ2AH48cBEL
2CNNpJjtmwO88pIMcfEZ0rwg8yOyOb8XW+XsqUpAItjFiMMnWEZUPG2hkK88XOVW
0iNrxo+qz13UmCNg4ikEu5Dgf10TIesqB2V/wUHPc0LmtZYPfC+l45xISqDxVGBx
1qIFR0HVDA38vuD42q5Slbfee1hQpgr418vF35nd7Vp0ai8FcIegjIqKQ/dYLPbv
pbi5AGO6XeiTxxtJGvNrn5UFN51VBUqrVUkSJCuNLTavncyWI0p+VEZFo3YX4fbx
9aTP1kJJcPxqpSWe18poRO6529dIt+l21hgpuSbHXLNl+C+Ju7aXPyjGDpD+gm8C
nqUoHBX3BFAhbSZa74CuwWmyH0PLHwicK5vuCxyF4qO8OcTGOFzmHvW5pJr7rYJr
6a2tHHLYd0Fh4UCcPfJeI4OWhvXvZ8G+FqbhLnNxozMg76EAQG+y7ltQteumIBBG
R8vSNKfnG6KjD3aN3u89/I0ZPt2TxU30abB6GgRYa/1bwJ5n2WnsVPpdn+8Tkl7q
JFec2JRn9BSm4DNrp69k3UiV5p8wj3tkRefvWv78mkiwcvSylGHlriAF++T2xAPf
uLXgH9IP+239PxSNisuP/uVbFenB5Y5VETP3qBstjUMQazpIpLp303rBBB5PdKCf
Co6F28MtbbfEuNZMf70f9sE7PCFO6UBqc/MOhMGbjTP64qCBwmJoCHlT7KzHUkR6
M/B0MCYYUoG4l6akSVhIVJcUK63ukKBG3To7tFAsvrFWxQOaRixPVku/xA6L3FVR
rZ8qM5GNWWRfj9UalIKJcVBQbWT7CNwpb74XvlkGGJqxPAsMeLTceHkYznQxvTwL
lBsB6Qucdwx4P5tRuxm54ifoPBv1QtGHGZGSmGcX+byEBt4axmj2tFTI+4S1DcPC
ad/Wamx0SNCOYrTjdmyegEtqbODDHOZNRGJ997shD0kbMq35uiilE9AQWmluSv/h
AxZPncGTtGtdGZX5t3fxAvLsPWSryv8xVcElQyyZECBp95T7TU+8M/YHiSf3FPsn
oPOtAyyIyLLBMUHbR0xVgloeqOBzjLLpadDV3rH+DxkTvTHUjCKlJttEdjezrUn2
ln2M5/RhtvmRf3pm3IJrE7YabM7Wx6g+puBYD8CV4Gm/5p0N2DL+Ug4cAQJe+inA
eEiduW1S5nkOdZjJ4/u89vUB9qZSeWFfv3QojjNFwQrqnUyB25ob9/ANUrRP2FpK
9FpnnZJEFDOPYnx27HfwNykGCKPpLBxNZRjN0dyZ20RHsRIqw5Wy4iv6GAqGV3gA
ApMgwDwVBExZMzQgg72uMpuMP4bDq90Fu2hELm22GHdJ92LOgOZPu6awAx699uwW
+XFEtlyW6/Ufd8jPL4B3F2w5AsQuAn1bKp8Yta23Ho6SYUNvGB0uIEWs6ZYJdHMc
Kp50APDV0/pLaE8P4MV3FEHRF2gvN+F3JN7kbj0qS9rupQd/P90YNNYz4BbDQX1r
nR3Hlzhc/A83o0KtBrmSshm36zIf6p/pWs2xF6qpN0DTCqh3uJx2f1+BtZQHkcvu
P/nMl/wLYUDHG8UOIMlV4R7+NohquJFiPAAY5LPpdWquEsRggdVjhs0H6/1H+QlD
G+e4XeoCFHbLJqBaGQsyk1SszcezPXQL3gyEvKZwEZaxw4eWzaPr2CcrYdjuIXI6
ygm/uIq1WKnBVCl+msO4YVgAoAl706uDTh4PaL4vxUIh2WtrZkknla//FmrI9Gco
Es5idgGy5V0m1DGJvLGIbu2a19iNMMSvMf0i+vgqhewyJd87W7R89eZjBWPuUsvS
ug1roWQVtgnzqoBf4gdqdiefv6xvXncC4gcsTSxypPfGB3mL+r6d6aKarwTqq0Do
9uLTG5HnAhabJ8aC/X5pXEAnBeaLhyzkTTCCpWLavagnWyj0Ijkyfk58BlmALR+d
jGCTRanOlPJX2wfcRibNIfULTM2XYakNChO5VxrK8ELAYdJ/xLSjU9u1VbHkUYC4
OgVoQsZgJ6iS52+tLSz/AO9y0nOK/xpGot3AZEk0VvztU725G3sgWb7V4t7qQz/u
RObILJqLAIFcb3yc6Va/l9vbyXKicvyCurYeh8eWAX8Qx/Yh6zP8tECUejHSUW3T
qI3kKR/H4G0V8RGNpVhvQzryafe1xnD61iX0goNYl0vLRqCLdPHExVXVojXYJnHs
1N1zk2xQ0WCVnS6FY1gPTtI4NTuYMDZROIHoc3DX/Og1mHBE951Kg7HBG2m0PiK/
bXQhOCerm0gS4jZMmBYxYB7Cn3SycPDFiJB1y/dJDlqeYRALvrgc3863LZ4H0Err
exTw8i1euFnO1CUtkkIXHhNgJT8LRN8f5KzbZKoO2VTANU0PU5cRKwyuHlsQsw1J
zWlkpG2ynIc53o3oapna2Wc8Nf0b71f4PB30J32/FGkiOtO5A012BCsBEeY+Yc1a
6cTLkZU0Sf3iSEMWyI1PRREANDhdzUTUP7rghFR966ic3J5+TdhahYEiyOpbLQM3
Zn0tZE3TjNMTEj0zpuKIXRHrJ4lIWuzA397Gp/n82i8XMm5ub4z3YZ1qGB4LGN7U
P9gB3BPPBxTUQzpZSfvkPRdIU/0x/YZ0DiCSa+E9edjRtFoCMDa2Tuk+gPe05YqD
p3OpPlTSMJj5GUJJtvqWwk5aZhvNiXk5KzuzP7YCzE+6is787KOE3BsOtCi9eEYh
bVSTSXdl/uQbCNo1mCBavici9PgCKnZ7h+FGMO/a/ilg4spUCLOA4meN+oSbowW5
V3nHGOCpjgjemNWmNNTzyGkvFaf6zREvXy1JVuDBjNTMFy4Yv7duqhlf3ptOXRAj
11pVY0LC6su+TrPslA0h3FZQk72M7OBron9BLBc60sQfSeGbXMg9ocV8Mhg1FgjP
a90d6t0EmUdnf0hc7k759A5+DEPvkSvzHmEPbhsowVQsC1FcTEhNro1AsTtE2heb
cDl4bZwzyuDcfQ9qH5btqsZtLB/HiA1j6ctZ6Y8CvC+il/tQAHenNsRmzv58ULtH
7SNeIAe8qlZDm3FRjIQV0Au9sIcMQIc1QfxOrtHWVPAnoutwYGaDXW1PY/wGb8bb
WedV53yz/nEhsxQknDsHEuVQN/kl+IMlaoUbYjsjGakhRj/BRqy0dMNgoMw7zEWz
54xJ9XJ2QSnpIN6AtnU13En/7ixTBLO1HmpoPn54bq2gEf2efkoYel3uaD3D28zp
TRdLDjDD+LR/swjW+41d5bBjTNv41e1Fv4jVJ4fVgBWi3LGghqUfCHLp8OKvP+v/
Wy2XgDRBcM0ElWH7GkCklzv243J9lgrW76Sp4L1V26pla45qm2MV8DKBYS1sDNdd
59mVO2AVpL8tbuzajP5e4wWQFNnazTNT5H1A3zA9wXrmD73mfjSPBU5JrL6u06bE
RIb3GEtTdAGmYQwAhZpf92+j3C/TxoVkzdYzi9kyVp6Vc/h9+4G3jDios6G4IK4l
TlrPCpVMUOdWVIdV2ElWLecdTtASGOyHzJTpMcC6sZw/STAk9Vi2NZNfYAGSx7FN
ted0HAW7EdVrAlyepzCN2ur8+v8FD4ZhUBkCZTgBJ503Y1DBF3iUDQW0+d+NVi5O
W4eI64x05ifKFUrsO9eReQDoP4nzB0zSJJl9oKxtdSvqw2xwMaZukAzYyXtXbS7C
2Jrsp2ras4Q0AnqRzYmTquZQzzv9gGJuIVbfU0UxuRYKF8LCrG19B0gr+VUeWQDk
aFFYLeRamYmmkM+QphRmw56VOW/J0Smn5HIOJUQdAk3SQU7bkCPvR+CSOLKDvjYI
iwM60h0Vo76eBjXjmUBfATTp05M0jdwWgJCWPyT+LL/Hh75LZAXBIeZ3NxqK4W2m
hHhunkRmuVRxIlQXdvX9oFBZwUs7vYT/tQR2wyRE3Be10H4OyC2qmddsQdVOF9KI
3nkwL5da7bR80E5wUJv85D3qAWb9a/n95aNiCJzUVN5q2vmOMTDSPM6qK+b4h8oY
4YUzFrHz8KTFArmkOk68jNhIT8vLoJK9m5IVZwERg0xqRvm7f/42OJ0VZQxt2Iel
htkQbAJcwqvvItRiJuHQqvfQ0SatQVYVe6jngXUHLGkde3ALKaaK9xlpo4rUeOLo
RgL84KN/ktZUKtbW4ZC3EJIdGaD4WCoecC5vYEifK382WueNOfbrrpI7+IGllhMV
mZ4dLCz93e88PFvZuubw0ApveQvikVdgjVpXPhygoKztgEv4bEDERBV/utq3ZIOx
vziOxyiB2LHne+T51VFvZalWwZ6R5GxKdchLifzkWdzEcatwLUXffTP1ggHcv9Xc
8vf4MSocEl/qlISZdfytnUChdE6xtM5S5Fi4wpUYw+j1TIotFE0CP+7ioirlI/Dl
BjCDTSwuDQmtMlfx/E4Ux1B/8Qsc6yMT1tKcN6JQB95jOPtpbUENkmtVXeBIdgKD
GhVS2zwRla29EuM1O4/NcyWAXXM/sjNO2bZ5DMWZdMe1a83xEUQqDC6f8bIZBZnu
hzq6nrpT1Zlk3hLUKfkXaefZF8LhjKareezLX3/rbVxYRwDuM7XYjbJbRIx9tadk
8BlCUu6r5SgHhahd6+O5dI7y90I2/3El/EflO3MGtt+4/Y/1pxwoWECbWoSIOzdP
dgg1XbsZT6kJHzZ6fUdBpv/4ejG/bczQ1FVCcuJcXUKigaXUCIn+gfbL4ZcSWWYa
Q7FYwKrcrYEd4cp5pMcQSGLRo2MNcdz5Kqdx6TggcErD3FAHa6FRRR4LttSPyyPH
pH9FTiZzOXsXhsQGOk+MUlqW4yBDbgKF6PEItazGPl5tBsko0roMODAPz5LT+ite
i9UbZ8MAMM+davMDG5Jc4vY6XaUn5wVPsAxr9CF/4q/6u9jAk1mNAili+EUguj0L
4+VdUbDeXjeUl7stdndEFRLl8K3V9JgE8aENGw65vOxfA+ZDW9xyT/sp7EnG8XEo
gGyCXDIiMeNF8A20XUPrfTX337ryhUxkZnIUF94NfD07JXVA+wuaFoX828dm3x8d
C1dLBtMRi5Qb7pe38QIMVzi3sKaFS6MgByYFE7RG28r3WEcPyUeDDxZieftt41sa
E6+o6S1VE472pHL0XSYh+jrsFr6MlatIQTjEbK6+dSRk1hp5dU9N0Rtj15NUvHrf
aNSD+yIy+SHFymeHtAjkrsGJkIZW1K2qIWStL2JVJ2rYs4PG/6BfJbm4Wfp+Fh0q
M0xAMyXxpyOTLdZ8RjyPy+v1+hqZ+iQ5YeQOgkHtqrW3Hzax8kDijAdQsvay6i3/
6OmtTIXifxqoOGD7jHNLyM/bfn68TIFCigoxltRR5AEzALvh7YHWtFur3keQzLh0
DMM/uopDPRMt4xOMlZbMbAnftfaKaIV+1W8ywW1VKOWDbb3rCqH4DGAsriUR5aLQ
f6+ce7c+YG8hHyCjd9IsjsUWNaI8Y0f1S/wDmvIEbxxci5cRUCJaDSt0Y/AnSBw5
PbZYWcJlZ6ChjNeQdk1E/wB6P6S6xvcx4mJSyFk3FYPR/c32mycpfI1WlBlDgLaa
aORZ8r+LD4W9CIPHBflHLbGuLlw5OF//QgGviDcB3+EuT6VsHw1iAOVq4/68Tn9K
3ofHPcYshVEPspJkH+x2rtNmpotIcBIRkIK2CfIyYv9bl+4hBIBICzsKDVFxB5O5
/L2olzTuomPynpLplJzhIhtKQ+p0WGdJR2ovtjLWgsznsKOaBtvXWfpmWOrT4kMr
y9tYRrEy9KoVuhyK/r86ImSVcKbClcUY56IN04MQAkiyrN+TmWU/xiZmDzjF4Bjn
eM9ETpTb0fNlSKtoLl2WRyBcRmX45EBFdBl//ydhViAefalTteXvPnZn6goBpLjY
8nDE3jj8Y7h+0M7LDFbr5fm28slMJ2yvUUq8tfznwi5Yj+S3wllDq6x6p5IoIrt6
lTd7+kxm3GLuVNQG1sWKFNhLeDQdQStE5PBohDcPW8u9aNnP5crMjrvnC0A1o9kj
AHqGchL8wj4N+73PGJBkofb5EuJIXbDoKk4ajmGwXUpnkfQh+zw2DiRWXWdoLsYH
dssnPhXu/2AS+DngyR5zZvYCOYL6gEfjazzoLusNNrFNpwAe621/QAGc2DA6Wyo6
nBdTPQU5d+rFO5U8EB7ZB4/wcIcLAhlr/l8OxMu2O7Bzi9rWTbD12Ezms7Shpoay
BLcDFY9D2eXDFCkNVQtNaCTWiqR3QQKv1vXLFSyokd5/hLYqfzhhiGZYXVJYLBc7
y+g4fxUyZ5GYIh7qMrfJyUHjOvUOPz7vc1oznypWlcSmBgJTEOdXACkbkByuCjD6
Mk/xhmPBpnGG4PNK0Ux169N/0zwuEaNDbPNQGLbEi5rG9hixQ46e0Nndw7bVN57s
BEfRQQgDH3PZQfbx7Dk3Sc5KRJLBAVbemURSr5VEu4Hsg0phFAbndxGF84QzlG9b
KCxtRIRE/m7e9YEHqY/GBhnv/jyVOJmX/mC9386aLpfq/RRKcRJrLGur10KTiuve
C/WsYj74shBXuRRxaIGvu40TLAclqZF9oHnxzbqBinYDKX7MpUevZY9JRTyLR/uD
ayID8ZDNmlXK651sLa9gtgc02Nng2l0kJuLl7wCUY0DVY7y6ryesYUHq9JK5Qm4y
wRLBotzF+8KDTu4RgGimqMI4o/WX0rwGlEJNuKSzqR+txiBg9fj44JfHtPjRfRhE
q/lNVp1iunjvlSMIYO3HqIQ3lwdDnDFECHZZe1Pjx0G0yFnKyPLu9eBLLos4ohnk
gK9gPzkl3R+iRsNOOgc4lNJH5MWCVWpZr1Cp6xAAYrr2eB2b9VoIH98cHOj9shfn
LgMm9yxcCqtoIuxbqVQ9JtVsIWQ4PdNIXsy2lyca0VxevyzWgm/YYwlTH7PJGgQf
l723jpOs7XfuEy3jCzR/lif6EDENqr4VIm7ynCKABE6tQGvxJcrRy0J83bRMywU6
JKqQKeLn4lM+YX+qQNqJm742n4kdSX5n8qmwA7ILMB0rRVp5ENeNZT1mKRokTovb
sq0MinqEc/sUZBL8PO3HXacVLWP5yHZNGx/vO4YS9mG0l1gnc7gowieWY4VFzIpV
azc0jy6yGduolLt1U/WVBKbP8dMjn3HYdSj1tFh4CTWTM9qpqIhQZbFv2LIohObK
fT6npwb0dR1y0Cra2sysblROtM81bm7NWEr+1nCwFj8MNN48ymrMksACT6JQa/On
EnVm2ULG5OxVsyKxfW47+w2FEp5wzT90XIQbeedIFUQUZBu+aBCaT5VHLNCPzJqN
geh+foAzdBVxGNb+1wqoGHoqAZLIFDOx2vqk6qKNbZCI1iMRIXmx5BTrn5sUQ/LB
Xm5k2gUDUQQFsi3+9P8IBPR+JrUu0bSzePHD/OaCwdAkT5xpjFB1RrGaWPILlPMR
NPtuN69s2u+/MJO2vhVy1jpI5HdLHdqS0IryQBJsO8/zB3JBzSshKXl1u9stZAnn
dD9d3ebOWkJRIjf6krYz/YNJd9dqtkqKG81QfJvnFjFlM5MWXhFSBAiuW0X5+7CU
D3kRrjCu14lervIj8tj8G9qfOkOpT++PTrek1H0o/i3KOp1cfZ+ftqQYxbwm/loI
nVhAifehz/PPH4fU70FgB5QZORvQAKBGFsvKxa6Z46NvbLCL2MALp3sTio2o8RhA
w4xODL8v1JYqZeA324Et69lvErtepabRScYcqBNOJYF49liNn2DbG2IQzlvLYaON
ZLIpsPlrJsx7l218lWevehP3cWNoO7CWz2WtogqCAOscUm7+6QTr34pD9IeAmx/S
9vZ9c77+E22GKhHAlY7DL0231aonRheeaqVGuqp/JklboGp5dWuaWftaHpMQW12E
gl6wB9eZgchPdmRgJFWE8F6agcilaF+RTHAu2z2ouCKpgH47Hb+PVPIDDTCr4Tzj
r+ODULFtBErKnQE5ZewqyBhq5FhItqyKjNEPEg+KXwEDTfFErGFYcXPmdqCgT2Jk
6V/UryK1IV/RuO8dRMNDhW5dHBMA+eEMdNyVBvXIyTx0/XMT5NQKAcbFDe8q8d0Q
Xb2vSII6KRKA/JAoXXpSNrNxpymkPBRx+oRujKBNNq57hXi/P9YBxg8hrPaME8hV
PUeYotrGNrbWV2Ox1F+adaEa9CKAEU7GQnjAXKgUZGs3PC/fZbjhuzNjz6682xqV
+B0vP90JTgLblrLyTkhxdIMCAjvnXlL+h6PJgk1noZ3BfUiduTmZ2Pr4B/H+K7fL
E41Rv6wTr5+58oi+B3kZK8FV0I8kpxv19FjYXZ+rYyp9+tnVlr+ig4H7l41uvUkh
hhMuqN7QC5W+XXCcY+8+Mzid2rEETk+qI6UsX38sZAeXQulAdA8V0q00i4TOWr+E
YMl/THKVupBdw2REWhmerVyhYIvLuTKYrVA8wvMhHbULNw0bPJqSTnlZB/iLuWbv
iETGwVTUteR6qyLsjkCIgZ/a8DYKampNSFynjT3uc3K682TZUo4QrvE3klVv5eXy
MgI8wj6sJuIMCCO/gzR6mqN5bdZPgD/jRSGb12sQzMLD5F8qpdOR94ldSxYHQtY6
kXRgmigc5bIsfNl90oZaXauM8TPvTl+I7dnI2KOjThV2NTMzMOrHmwOGwl+MraTF
gmh7AsTwysCxD1NnxwwgQ8SHo+5M+kE1Y7BPA0hU4WajSgSOqr6cXBIMV/YZ1/al
sfvcUXEy72ik/3YilaBFiVlc7RMUknKrxXUrd8JDBrQ9UABUpls/ovy49TpD3CAJ
d7MYM4mX1ncgIDFm3P+zApLrFBVk4tv+Hlk4vKCs5FP66KU0duZ260zqEJm5HGcu
kjcXCZ+9nOS+1BTARiPxQTc4stA2VYQwNci/MMC1wMygX4fQ35MN83AbQ2Wof7Ut
pkFwjS3/Yc0ecCid1W4ppP62qdxOellVGMpzp9YqutYbNTheH4ioNShIdnjgeXVG
atD/iinckYNDk4n4CzLLFYUM0sNYpLQPMC2sa2yOmQMOyhpg54P4qdmfClGJu9kH
7cuNFESkdFSWys0KrEyXBmiMQK4egS29aC4/VeGK52BQii9TnSP0QUdnMVMzl7js
gEBoiZ5gmJvWEGrJUJ6Ns9dMb3F2if6Oh0gFm5iGLLR2CzxMbpoP9nd5I9REMZ8M
73HaoA/7umzrKNt1VqcQ8fj/675XKccQ+LNh7UZE1zGLsj0RWgA/3NmPz5EXy+VO
wgtQ3CiN6gfeKNZo6jIYz/huMA2C+TgR3bvPpgG4InxxgKBQfvE3NW6Q2ERm4kJw
TT0utg+uqoMQnkLGyJgpCcabauVWzsrutrHMjdTfT2oXHoHAYlW5qYLaZO/TJD23
wdde8gyIvELQsVSNcfZc1HQ/PDCnK3krG/6fNhew/XsTZroIjtpFzc7qpLMFMqYF
60jWypUYeer/2ClpGpP9fBj1u34BWoWrv77nGal7wJIiycukog5exvENWx2gW8vf
RC/IXEBG8PmmsSkBvEOJ/WLW2JgLLyD44RDUqrr45hjqlE6Fnxk/lT7e4BAuXQxn
MJpFOggf4DnB+/mEns4E22N8UHoQC3Z3eVC3xchvO53RbiV4Tq0vBAlqgxtaotKN
ASo2KmQg20eOUtddEOJuJK/tJyt3nEr9sGlAPoqzrb0tQKVyPXMcKr3ljJ6fIo9I
BVtvEta6FHZiTayibEGfHR7DIJgxW1yY6Zn3Cdw3PpuNoO3c0NF9Kx3Y0vAA89ds
4l4smfB+XbZaiQ73ClOG/4J0b5vj3tKHJvBpITdhx79Q7TI9zNXR0EhuywAq/m8W
6QQsSpJuMzGh5cc4LVBg4EVWvhtGJmh+Mj6FonSiG1cjy4j1twRSdVqNVOVf5KmE
hAKPQLwffGYpti0Tk6Lw0qURzLPOTECmRljVlnOaKQWjR5GDgCGM8hO67606b4Fs
l0zaYm140hBJOnzlUW5f/YnCA4+lhOjq6SqgjmX6Ac3V+1tyxXPiXaqeWNF9FbtK
erL4Yx6vWcSXRoS/8mlnVTlPddnJl9dqf9hwhg4G1y1nOSK4LnvGjP7aOPTKRLxS
EfEIFv5n90kzVi9Y3jIqnYCXpYmWsb/CevTbFfXSqYMEySUif4ccHdd/tIG7O5xY
kPjLz03n6F0qCtYzmG+anNLvg5RJTWMkOPRrR5sRJELi/RVh23y6NhKyU5inAwDN
8JWEVX2kfkeqJG0ZQWnQL08LM+HVLnfsB5pCSqHWoEPiSRR5KINsF1HJKiEW+XaR
OHIiTlm2Mun1qaeEr1XP6FSxvdPOrvf98QGDal0pgJ5pB9OoZLS9f1F1viYVhyav
6k+sebGTzdyzL7rJWDmi7uQ5s2uO//YyOqkf9DHml7PkM/3xRvHykp97kzKizNEc
iet9jsNU2U1bsIVEgQJivokKcyGNJ3mMIW2jLy0puR0wfrJ6LAiuJb8nRMoAgAKb
ZU5mTRHMIJHngTiDr+wF7xrjXlJ6gnmBvmW/+dhDeTdQc9jTJYqoAaxieOOiJTbT
xgiaxyS14Bxp6KHPvS3Th+CijEvjZYqm/ejuIduDJPtGKDUTIksxjltZV9n/eKHT
UrcvYKKyUFbXlz3YYyXrt9rmd8fpblf3OwajDmpB3C4Wqr2vwxS+NeyYRDb4D0Vi
fjWTzAUgm1/tIfe/TSkrlB+vZcxChhyhW+nVMCIIohjOLbcJbDsMNr2yBXtx3859
hQTeDukjzD0w/ssP/vFh9edCY0g24t07U+RTSA5Z/mbDkvoncNa+TuiZbbc9TUjg
MWwgxJwPOOlNnnOm6BoC5QTxK2DfhqXb1IyjB4kFNAsoD3qp0NxNydI7khVOmJuH
3tdsUDJHo5Lbs+JkA9r1rw2/O1N48siFsGhOfP0Y7FjGXAirjz2x4O1doGuwXGek
uEqn+cYXyBFij87K8T37V0PQfE3AV/S6Z8q3ZoHUXtFhglcaHey9F7AUQzDpRSva
MoRJPb2b1cmUvwRzBbol0mdnrOYFaBc/rNGq2FG982D6qP7NjtPowbiwxpDx5lCz
Lo04vGOYggOiOA541K+tQ6VLjjGoE1NSLSVUs+id2GEGZi+NwiVGMT7WHUGLymOs
m9xKbE9Y23eBiMNMgoXoWemJTqeK5nE2ps7OPgfIcwz5+cdqTiToIe0Aq1dUKIzV
Quw0lo5buc51hh9+ZoqK1uksVlbjEmU2UpsNe2oOcEHm5CqZcN+hRBYvnd5umYZ3
7VOpGlw61trlyyQsZ3m40MShPYQtSFPFUKidmpP37fmum2tI/Iy5jown0Cp3hnix
u4ZhyVVHO+/UI7uYkpMCfrqyOEZvMuvXRVhNw0hNpLTaEJLC/BI4wgr3stbVb/UL
GfLKaQZmgy5pcCckPzWz6665sNI7g3g8uzQ6U/vBozITJwaqS83Aj683bj1ICwpu
ZaEcd5rqogkzMpXr892jUbTE4Wz6NtP4MblZ//P3yJ04+7pTXQixB1EUlVOOMZhe
2gCwcX/1NY2ZAe7qnyYqcNV4IuGbH0v8Z2IBRm+4bAgBJ9larjfOU7Aywq8MHNRw
Fiwt5PGq5fNpEoD//ueKUug9zIPf4sbHYBIbTdvKVXkvkQLgBQfrR4PqjztotMTV
gdklma2Hv94+vlih+f2GcXjEFRMOH0bXXdGoT2QW9DJBK8xojZ1SphAd5BmRWv8j
NyeBmFu04m52nHCOl0woaW4d9g0b82BTBIXz/M11q3byGNQg6pxo76sTMhb1hWCO
7/2x5mUXzIxqFZdqvQg40UKjAgJwv0qvUXLpmJR13U/lo834deNoUUI5/vkIt+7+
6pRruER78iOIxY2uS5pnZptxH/no+xEOq2yCvT327/t2eXi7DZpqisx77ahLFjQx
J/rFwXveNJBlMUmF/rneSdXnkky3uat/1u9Ob9YIZi3vhbZIoOhFqXU3UlGTBcL8
UIT28VnmoU3aZbzrvGg3LI0yrHVLmT26mZtKYn5IitVoOt2F/jPfs9tPJfbRfIH4
g490Its4/oSigaeKT5D2McCY0EwSQJ0FPOmUZO9P5K/qjkfq8plTBG4/6lWqhTHV
SNbp/BGfJX5HcGhxoY2a2fAL6rTb4EI4lms/rOKVpw2L/XZnEYbkzrE4/MGbglXG
E4id4rEJCDRcRYE6LfSPoX9y2KIs2HgdiTLHbneWD7n7Zn5q0LGRwIcWG4vZGbso
1Bxw2ZXazY86QjDYVldzZvSCXqN/4Q9w/7aPmDAhCYaSchQbJH/mt5JoZzzGQuAl
6IiowULWKPBZiEv82LCBAGWTrK4yiW0vquRB9+8FlwCp317dYd2OxB6gHxODoNHN
YY7oqB4qrEBu85n2k/D9uiqGVKsmOXaezPPrIKVm4IcPO8qWMCpuVbnhZPD4Eukv
LvYS38VIARq3fCJYvZcWyyMImn9Dz6Hb/gdw6wukp6+1RSVFFd071vtnJ3Y1c4D4
YRgakMJSbeYevmPUg/98q8fHbcuwoHaLiu1lxpVSxECd3O+s1QQmSwi43n9YyZ1h
euKVutfqYjMEA1w2sMYJl0HJ0UeT8lPTcuO7P7KEnt/DnFb+cA0kwTHzMlquRADB
YmKjWggqM6c6gJbLSLwVPnuOfp94Wk9BdNmaPZju1WJpvouyZV89xc5WC85Lcsre
Lb8d50g4VmE1JpmE4RxBAYgm3gPf20sSR8+Om6Zw6lbrx8DWLcXRd3wHSeb7+93e
FOPf4oHdi9V5o+1fvS4pGTjFiTyDA/y/peYxg1xYpIiyJGUzlErKsEKAePttgTgD
9C+vrGm0ORZDrnypQWxNENeM2snpvbK0MguQCEcUuOjktl2f2IGcQ7W5LT3rQHuQ
IcjJtsHvelNFtlTqykPs2DVToP0tbSCK1mRMO5fKpzl5ljsaclaoiKb552f+WveP
MwXxAj4xW4ViIeA7VrJlueRD/flddz6c6nMnFm2q4wtf+Q3o2YAwLm5AZA9AdGM+
gPPv0zT8034z2Zk1Je3SyGyrHXZcGsP1GEnzS/iUXIVGZ6wd3oh0QytstjsbeqCM
dRjLh/LdgIPLl0QAXlDylgp3kbVILcSxg++6LMSYLEG/ldAoWciaFfgullznzDL5
l5Svdh2GHUopH34M10XxUeXNpWkaUYNFLEJxodblEoPQ2Z20KIsUN6JRF5smd5Ag
EJ1oZ+GdtJP/0ZwHe2r/Epkv0w5KdJ6Bn8GffNZtMDYGvaXlZZsX6h3B3rzVOwWP
sddXyt0TmWPt5/QdL72n3GaAZoJJU0ZrR1fIJnAvS5ipcQ38yx44m/ViritQDlpG
m1QODK0ox1SdqIBlOGPjogOuVPvApjCYLeSs+3BXoCWCywrwEU1Dh2c7nP6wfP63
cNftpuoYpcWM4buCpN6avn6jqU7+pvtY23rKQ6hSEboxdd6tb8QMjLmbkioXkoWq
v0GLpJ+kzt65t9FK8nWFDLLndphPVrzza8oRdRVcT8OVYAYxZXowH+2pXrrW4DZz
tLfP3BkvShDidAT6TzY5Ax7jk0uw5Q8WdirJRxULNSvvN+Hwpsivo0C4b08amL5D
+rhHjiEvtfxLVoNpG0SZfVZkWeeu6SRxy+UX3C9WBRygjYt0iTCWiMlMFEfgXh2n
HiwuVcCa7oys0qb9SSZJPCJMuP7iyVdnhG9gs776wgFNW5vqOiWl9JHko1Mtai7F
pVPFYBEa2xiXk7KhtSGWQ4bof+HwTdu/gQY4OmQSMToKv1PyuvEGdSMOQlw3EasZ
dKCB1a84GWsuviw6lDf+TbNmRrwJ9IpHfDttgywHqoqoL3PzTltxLnRxpRMTjQzu
7mUy2CJdmkM5YKsRmQM1bnfo2fMumatCvIL1EEyBvtqs74kLwlIrnuGaXRZN+PfA
Z2UeoH7YNLw0MRh/Q70lqYsh3rjGl129duhcLH49h8i7ZlIp8SRpjAhjr6OEFNCZ
OtEVEchX9uwNxkKCpcbDd69QjWl6ixvAMmhTP+BXnHAr/jYHS8oQ5TQYmbLUFf0F
FeUrfxPf9B3QvtxQCIqiVIrW2Sk2L1aY1z5cV2cG8qhidkkK5lR7uxyDngxMBkr6
Of30Ov2fc8/d9Z1sCWnaZX7BbVL9m5k6zkD/eeCyiZoUNvhKWelGxiGL0CxSxhpA
x9pokZ+3KLR42npd8pwizEjhbz1LmhedgVMOT5JLQ4nTmI1nkluYq/XiPrEHHTlo
XDEXsnZihhiIxpa0ymPSO9hztkhiVc4xSzeUny1ft+YcdRynZVli2GhUKn0Tm/ys
eEJwBBqE3gEjUhtd73cf8dw047RjSCVSAHdmeRkRkZhtLTCbzQsOpd2TXqYpLFAz
alBivZvGlpCZTxC6yUc62SxXbr17c+4cl0TZO9zwch8twlJ5ucI4QOhGzk9FXBx4
VlvWg3xQc82ryk5r+jpbxiNsCEezwy+Xra0z9hee+CKcU3og78BvDRTzZ0BXdgHv
CyHORl/Z/Y20gu2Rj06z1PkR2id6crHV5HEAESedY5ONl8lDbeoQ+kj1snaoWI+p
EQIUxXCbTP85eGg1+XtaZ7Hc67+iXTvo8UiV6fYo1h5ZFWDaipsk3e4lkT9H35mk
awFNAYnbT5dvdafg1hR8BYBuf/1oDcVnPdpiNGKN+8o0fGTpLwp4CNScF5AmFrAs
6I+wleabtN74USwuNUzsTNyNgeEQXLuIilD4/wGo6U1rwmUf1wXKT2iD+Od1sD1h
WVuhSbLX1IW5b8hPMFJiaTgi9nggycXCgkT3aZVPtVUKicn73/CgvkUexmPc4Eqs
SuMvfFVGsQlonSmJXtMmJ2etnwFu1qTtNte1+Lw8oXt1lj9cdYWbQ+QsI0Q5nGuM
jYhy4OLIbuWH93KHZeIkjBIeZYSaJI9cK4cnUZOjtzIKo/QLG0ioFH34sRJCL+se
xP/J5iBUYvuDW9OCsVqR9it3Iw0tQkwKWHLR/fL7oB0MmCb6ulPHPdNpP/ujhrUe
zcH+45EiA3+RHtuIymEMEzY35oNfUWxviMAK0/CskP12ykrYmwvKvpQUGgquQ/Du
gEe0YUr6ln7ED4GY+meQLeAklRxGrHR/Hlai4dDmonxrM5KxFKi587gjN0aUyCFC
ZiX80oS67Xuxdma9IGxB0NxbyFO/Y+rR7sxb+h/FT6HXQIzbOAslLalsKI9WvcTc
MEgboM4hxC5XLP6iYsu0gQxwwXS48nki8r4a0sghARFi7EiUGI3amGYblu7xWFiM
M/YXI6rx+58UwKWcJ6F3E4vKYJSeGbyp/8DiXtsjylYFWtjJuVmymkKu1IeBEGGx
XYznLlgirFmSuCiI7R38SGhdz2C8rkmqJ829hBkW+ixfbg9fOCrRcYLar89BZHM9
QgNsqwVm1j7+b/s4zbO6KtQVJnJGyY8nsVT3ETWLBwI0JwSx0r0aGYeErHKSbTrG
pmX0s3oZuJ/Sg32GXFd8uZ9rP5ceerX6Kjw3e8wzNRdHnY7Zvnv4SsU3hdlb9jTx
K6qqTo80EQuO5b55LKCRD0UW4zpslF08VjDYB7RMHoXyBeoRsBQ+JpsK6o4Llg0j
PAWzaOUZaPoL8EUNGhz6pUyBvv1rG4SgnTsANRfyMCqrie7uXBeCe7ruCKLbxZWg
3/3VEQndg3iojKFro6KhHSigUpaXw33UaGphSoF/aan06TvyppFlx0criS9w/90L
8rYIYEjljDalgBrtu7TMx7aWXdR8RElfrgzPDAkw7A4XirSaxoAubMtUON3eRMMS
FuLfnXgqGGWglwzix18schIuVFjJw7TG5+ddN3VbkNgFQeGTEtckv9I8Qe8g8Sx3
uIcqaZ9Dq80PX18yXJT3XXSKxzAPvx0JelQq5PMcThvfL0HPYcGryMBzc+dQrQ67
uZjz+G7yNguK+wp3mLHdRT286Cz62tNdWO5izmgQMn8wZy/d6Ij4AMLgjidTCnb3
gTT3bF4DEkw6DKZVJRE7FkkV/3CQX+WV4hM13GNvmjiXg0NwIie3qVgLbI7d+rgD
TU2wkFv5Ev/w0BRCyib/gW6SgvrDvKSQicHSeFE52Z3DRFJpI/Qc8ao7t/4BKHh9
2j8pzKqF38WKXpaX+oR9Cg/8t75/xQ//KxohTuZ219XEbxVw2npuw7JZ0Q3BMKXU
ni2imFGjxBMCLBkbW+plGB0vqmCmpqjcWyDxUhu0VnUQTkBpxavno6+2ZmwwHuwZ
AYk9inPxgNPcuNLb3FYc02pJFmQ92vhPrU2AfU6GNEkzc1RJ+w4Jt6zKjzpDaR23
9nmZa2AMnXsIF1aSKk1G2IBqDFyJjIaBKueGOIR8LvH8IGUPePFYSwvBfJgJSMfv
FwbY8CeyC20ZRFz7SaR+pKSu+4r66uQCbVoL94Iou18R982s7GqWdyB78MbsxnsW
/UVRmJcb+Eq6dzcYbGPeL9j8JyLSIioJdJgYvK84p0oso9LqDR9kFb6G/Tp5Bdr9
L8OpYZUiqC29CKppLhkR3usi3a74iWmgzT2ig5RwHMsE//3Y1DJyTGPUFDDEP/w8
biUp7f414srbgO2sIc5DmbprvFKCJbLw///Vht3ocvrkkBd9lWF4+mpUaLoZtQw1
jExfFTt3T04BJq/JcdXart0ULARglDpmK1NXYP7GK+vjUbh5aIREtuhbQGqQ8qfl
TepNwwSm2+L+uZzziCk6yDczXjJLp2heWAqvzdSLi7aiSy5cYMTi4TeUC4nCYJC6
6lHH5tj0Ih/MZascXP9MsGf9X83+BbYFpedg+3PjE7THZBWBlaGCd63xyUMur9lY
MTz1Kz48BFLBrajSHJYcyqJ6sttk73BaEYtB4uxPM0sRpofsIRIBoz13iXeK8fsB
hcxsNIot7LEJ8mCSPttcTQnP+mEHJuASpnM9DEVa+MZj+XbYnCJcKr/HprOt7yVG
/vrybXMXGWL+WySAosjtRVaVixlyZ4rXc6rPOcve3OU2GxXXKMIFjSZqvsWuey77
CDW1I57UX53TdqqPNPTeqBf4ql8C+sLn7IQIz2dKdJjTLrRdxz0A++tiYZkSNc6Z
sTJBFTQYjcc5Ag37oQDDSYdH5uPJy8rI7FViKeciB5VM2yZ5YQK7vBP/Qqdix7J0
3Sn5xuuQvvMDZBC0+QJusSKBAUsfXsmNk1MLUEFdZj25YLkZp0h2IjcL/0w4ieFP
UP0O9U+DhCPVD7+kt8VMRrRG+lvONpBK4qqN7lT1FiTWMAlraxpcBuOsODVFHsv0
2DZxXXEPmerc7O+pRvi4IG4bHe/eFHHJNeMvr5EtoKQ2LZTVT75+Wsl7vv9pgnzl
z+j5lmawr4RCjIlC1h9ipyV56q81xwMzxdDHG68xrqvFLRmvI4JuwesyPfOziglW
iDgy3SFaA3H4Ojc2fObeCfsJPwGUvPjQRHg0Vlp8ooTdBjfz2qfv0V8zAJXjDq1a
7TJrpuQcG5EuobJkEsfy/J0lTQzA4R5xqtLBDlZREBIYe3N3EE7+MZY2mFyZIvbN
+FBB0XV2k+/mAg4Uund/C7bMOb1QMXHb36vGyh+n+TPTOZCsl6vpIN3K8jqnAh/w
veEdAiiApgzpq3VEiKdB6Hn4zGZ3x7ZLMlClMhf8sE9a7D0f9mNKcTsoVu0+Jewz
ZSo3zfj7vRScwjXjjG1PzkHcj8nlnUhgnnj7GPRFa4dc+GQEebvc0xvav2/Xhzyv
FjJPTTmlzR41mcZQwWMfqeShamJrCMkMtzRAtLv70cuF5eJ9wv63hHP3D2+yRU9B
BKFF37xOjz1EECVANW1w0Qewxssw6iXl8VJDYILLDaIyTwsZbKkZ+d1fwrWJ7DoK
iCtscyBR1MmatF9XTI7tm0ZlRjm0btAtgaO7MtMO4xIpgzAOPG4NvHoWfBa2w9L6
FClIM7qxD9BdOmp/WT88XgVshUOK1/Wqfs7v7ueEsNqwWVjmFB5/KgSH1/sBTM6W
jzgcR6osVFJ9QJSqcaoH03TFItn2mrRU2DxU1FLxp0uq3Tgwtv8DHqWXCuj8bNZg
CEtyVdNCQ1x9wukoio5UYtY+XQz1yuTB+TtGnM7j4ErULmsaGQ4hQfvcDDq3U1i2
jxGAOYEmGwWKbsr8ob0FQdXCnmqaSQpFr6rBQXgXiVg4cNFrEDide0kCbfTgsRFx
gZNbl7xyODsBnZLPCQFE9a39vPBBNhNwNCYv5xO+h55ZsHWcOzjM42Av48sgaygJ
mfbH+IvSXDILbeGXRRwn2IcGrVDpbIJg8WAfeYi9kHhhk8w5WWF9yVZ/UOtY5UNl
dymsyi314pjx1FHOIXwjU4RFj8KGPR+WSCfnpAy/jOt98m8VKMTlX/RdVkFLywO4
DLc//A2762Lx1vtpp0zzDrugG4eXUwOb0gq8Expy5Pwz0duR3TyN2afti2de0/ig
8Ufq+a9nN0EUIIqTKtJYi5WjYInQiJhYmLZNEVdlyxJx4XLQPE3HDUYiX5qGDcwB
Qc7g7KCzDFzD35ROsIoQuSlh3vUb0PG/mFToV3qLy6GrrB6OUBvgELa7tuBxS5zT
53CNTyKH6ZLbu2ykkKpFIpftsJxxzbd/Qvowuoyma3MTnoDSMwxjk3oEdTK4y1vy
PLgirXOw+frFrskwvmLkPqUlupBqbq6CZvKQsVZyqMb0d3RExspCnn4HVHF/B8Oe
S5I4WRA2dwZZxs1iL15kec5sy/JPfu9Ouun8ejrTTOq3YJlQOkMwP7iSfcVeTWpW
E8idIQoygJKnTH828vxHYwx4TD4wvNPq3pq+GvUWDDb2ZOXSQd/jl6IJB2/eTgRc
JA9THSTX+g5wNGgzmXq0LGxRtIA0bwEEHqdUZXkhV0F72ptvdNr71CGLajmLZEXB
VMgNJJvtlnyAAhzCUt/jXdkX8yIU64dZWLtKjfiFJSweTQE0rbD3AQsJyej6LwmV
WRTcueJPYBRd/iPpf/hkz8hZPAseF+N7iEjGT5+KKXVJPMMlLhMuWz96IyrxkLx7
EgTPC3TfBqb4eJ1nLfGDG9buX70i/9ejbnfIrNnRNB/Dkc1R0soCIK5JnvtcW3c0
+zeHJQZpKXqx6a2hfQ9ZO6PT+j3qUaxF3GFw5ia1wY2UBP2tY1fsfBKJfQzKdLb4
qmdG3K6u0cDilen+MDggTxxnBFa4yQzYMkFxGeelWok5JOQb/RE5UgPix6IUInpR
4lOKGhEoYLdaufbNpinE+0EOnBJQhzjM8bHBYUYY5PASiq9M783rssUz0guoMKSo
eDbdv2Aykx0Oy98sSHDz8nnmZwwnNzzi5HxhNgekF37t1XO9zh/HvkleU3my862Y
eTi6jmiWkZrVwqA8WqzTwkyQdY61sRseNQve1aSQg8LhzpopWsM111vuvzz4ycLZ
2W8tqwhHB5p5X1xI/gbZaRZJZpw9yTPlFdx3NNxm6Z4oSBjY5HE4JNEi5ULE3qu/
ArdWXW8YOOmJaoFX58JLDE+ksp8wreL+Hx9q7UEHAGuRg392ptm63Ij1jdbxc7N0
qMBQchS3p5S9uYbShzov25wvnG4CTLYnuuRSh0AJS2wcQ+3cCXmBADsOoN4MvqUP
ET9affmskAGBAkpMguM0lq5AWXwzdPUjePT1aWK2rIOQwWOhgD/rtonmeyRjwHac
Ywoqmk5FM90ckaOE61pX1vy/qhiaQ47Op94KgTO6G5QRxZcquFTuUo8TrEGs2UuT
98tbV1Y9ux5QG2wcHaQ53J7GHtxgTjijK7ydLOfs5WMr3PwkwionxKaNv4fmhEgY
ywpo5TGJ4GUrUIQfj9UAi5VfU6Eu0lSi7/CXsN73gu56yvDOBugdMvWSs8q4xXHq
9mPTggqy+uAl0yRWbd9hKz8wKsAAyzoEtxb1BKS6IJb1gPa9tQx190E2oepx7plA
OuWSZJiNk7VtI2QcfPodcye3UQ+MbSy4cC+RQS5fVBpC/PuREVtFdYGfC/RMZG/3
ukrrtOmPLnG24LzpHAKUCs/+JzIstmDT5/5sLuBxAy58vdhQKXx+nXWQygf+W4QQ
R0axa+wpual7S3U02O6CFRuo1z1Q5yVmxuB/vakOomZMnGdJP6/nh/Y2KmnY9BuS
E/g8XdmHJYBqaSWb2qiFRa6A8U58rlddVOtIrE8ALscMM6KT74jVETtYMeiAd81W
tB4rxuJbqkJB02/ds46RSljVjA43uYgt4CT6VUtdnAtLKAT4pJK8HcZCRmHMFVNK
rhGXcHx/fMtiD772hKV3MbYs45H6x6DywLEBF7bWoTB1+FuLpvhoPKUHpLeh4BeM
zBZ8bMdPhb1n/uJY9HjBuc49t0Cz/H/6Pe5GjFeeGdZHAoj8k7wayaF/8FPC8XcL
YPBCgZdrn+oQsqsfU3rkmL/hUvtqfWXLo6HgaINjh/slLqGOEa1Y11M3SurLY45u
saHTeEFIMmb2My83ZI29If67IBiXKyXEOS302JbMgQIQ3iClNbqjrSYaNHHnPJ7q
wy5YmS7Ra4JXrcAnBmMVM4CGCzbD0Zd7XotyMLuOinNwe97xvD2qwob9k8w6SBoy
GUUQ5fnJ4GulwIp7e97cE17Vd8J27vy6o2bCkANo4CKIhFSGKwloCU6K0hJlzWYu
OjJphG193NaO7SAg6J30gsGT+5vMVCNaNLRcfSDe4vR8CjUJ3IcD395XBcAqJbnz
tSuKF0UvQlWe78tV0YLKFFoB6xLvHSJtYTkRb65KKGgG+SevqbYdEE1qSV1HUwbZ
vF4oxDsGJNoIBp8C+zk9wO5vnoe9MfSt3m0/R8I6b/auF3uS/qgUGhgY35a5CEwg
JE8qgGhbT3DdeqzOHLPCI4jLpNqPnl3tVFfLcdZwMxtItmoAH+QjAZQ6fkFw4+bA
fohhTW3XLpjYAz9SB65mG4wVbgW60119Tx9/yf0WZ8g5WbElidFJiD4L22JBl19d
Lcx2G1rdOtk/VcEIKiW3w6zdqKYUPefn8vePoIBIv1uw9XbStzfJPpRyzux6UM5Z
SVFKNIG+mYUWhhny6rLJKi1LMkYIw8m1gW5BY83D/cxZhmCT60yvEj3yUInjeSAy
7JoKLyFUnddI+2TPY2RHEwMWBpnWnTYPyAop0mkTg5r9z23GrF/achNaRFE0Dj6k
qUQmofbowFq0sVP3cw7fLZQTIfbYpE7ZcaAHWZMKyxKrwWklcUKaeUZkaG9J3rD6
0wbJY+HEPKM+MXJTicGuvjbXnCxttx8BawrN0cC1MbPVxyihNIWjpJIg7I755LNP
SX/nLM31tLqB3FJjgJssZ4F+rA4RpGA2Z2HNN5osXwkxrXPgVBAxT7F663rQzgK/
qx+RXnbJvrgrzk3p+ytttizLFgl1dxhSG85VTX3i4yhnN0GHPVhmBWjTQuQYcjj1
meSGWXCCoi9j/faxS3FO2zX7PoI0BNnoIllgiSg3MfNPZ3omQ7B1pyeHvIl8raZy
uqY4y9V0kJ2QerNqZhyqOX59A3nBytW4NmLGFdTJhjc/dD4Do3AGyGPlHa7SeLNa
6xvnPNnwEiqRyreqC+pYx9tmBTcpSJaT7puZ90+EyWBKQUz8sVQa75XFQn3mudGj
awvsDElfyzxUOQZGHjzk6YOyiHtN0eK3xHcDY/ZqrfBFKpX8KEYTb/nPP9Jo2piF
zIK3qbKmn7ZV6LcKVToDnEWNvLXn2xdOMfEXdG9k8uwZfsqWnsetdlmTFYFIBO5n
OkU/dxObWsfBS7fnhjdebUtzmoM+2OSEtTbKh2ramNbCXci1N8yIAP4IC4EFQoJj
9Cz7ToySTB8+uwatdszNXWoryjUYiwdnqZLqgyZrUsszcg8fliKYoBjIIML/1l3S
slIghpHLLEBZxpvpBNK6ZRDxbRhSYEtYHf4ESWetWLyL1SLXrfhoSmtlGHYCFDdD
rB2V1987Q5+v3R+PKWIA7BdP25U9fX599IJVb1yKeeshBczAOSZ7KWGVIGNHF/wy
TiDb/v+5spGnxThv/V9jMcfGvT0Gt+YC/0ESJ/DAR94xtUOh1AiR/M37HkA1IirR
3vOJ+uIpmlk0oPAnAQDjWD+c9RQFNyT4hh1MvhcYBTVHllWJ6h1vz/UBoUw+axQC
SPKHmLJBTRQVRo6SRT3iddgl8AgpwDyP6OGSdw742LECrmeB2eJ0E+R5HD+rj1A9
LPaxf45K16llvhbroH/gIaGG0f0MU5chlGV5OURTuTs7NwPOMgcxeoB/Q4CY/+uK
QNx1UnDdtSa5LPucx08yZT/TUDmNlCbqwnE2MyIhKdo6QMt07dAVeDM9aTzC1SiD
BJNsxFqmGg2m+gUGU9PbfKBcnT8HynQrSIZH+4n3b+/RKSrw4F/JVOh1ayI+Mfy8
YiYZXfVCotN2ZOu2ByCikJSJ1LF5em/AH17y4+OPrYK0xvaGcHJI0rP3iWe2nB6+
Qt6ETIWe/GO+Yw3h8t1NThLCgSkFygMoTvIfYjOUra4EBuYxPt+7J9TJXGnfce/i
XZeNzXFNAoGl/9q9ka5yKL0PRGFckJ2EgHNhPeB92Kr19hvtQOOQ8rGbSjYcnjT3
trk4gRhHfXQQyKRLJxIZCqrIJ03tM28wN5pm0+RqLUpAQnSJn8fnEvaOG56jmHp5
eXFVBb59F8PSC5jyxqR3GnYK6hUd1u6ZbuW4tjX++2lDBdh8MLDvfEGzrVZ2v//p
okVXaE9COtuu10VTo93Q+r4usuLWHKbQPqJLEUzXTbTJbgYeLaTJ+X5uYB9+Eb0b
7TZ0H1WpLFb18Frgj8nzv5Ba/02eU3VyVx2sSA2VtxfI3RYxiRtUgNNYeYAzRVJ8
67QHxTLPdtevH0EpoauJ+wBXkaxKHqGrNwFzeIYSIlAcXTZ2AJHomP+UJw0C+lhu
6ZRnZ9xAUrubi7uvp4I1QMfxeOll/X6TGe/Ge48T8GipIv8H0SkEBZd7NUk5ucUm
kymDjy6rzirtgXnv02GDjCSsSVLRHdtMXBsVJKH840I1ouMuJxkRbtKCcFbZ7tAD
NzAAUlPyNl0MnrNl3UKhvzNTAYAbwBsZplMczU27yY53tTY3COzvPccp6Y07tRVJ
QTYCUgCj1QA3cNNVXbecfm7w+v+AgWn/XEVUVx4OfWl7MRXOOYfdusJiFxdiirm2
ogGxFi/R7GaRhzrh6n4MDacaubQ/YzF1CgGTjMAk8sxf22xyWQs4EX5v5Nb2iqd2
RMePov1y+LP33yIx1ekwwBoGDcOObrcDrm7sUHVn0CfbBjaPBmSQQeBKBGDIyXUS
gfn/CPlffYijgX/TgsTGkTbK8Zyq+b2WijV7Ega6GhzyA/uIg0Uq+BVNLIRcxPL8
3HxAs1fu/5OfJ3ybLymLz63iIEWbT0GCWjV5194tvmIAWfXt6LbF58z9xtapiHkP
QB8Zzw0sv2bQROF4z4ANOyzVbj7dB3QBj8GPtNuPD5j3k8ixyrPVsHxUIN+tULlV
v32q718krdWL28nTvP9TUc3V4YC2CUtePOjhDTo4m8tijNzpbLfzpz1WCfKHDHbg
FPyqCgqVJhsBQvnaDEuxRZGPHCBOKYYIHcLqPFKgI0InfqfpaddWGivjJcQ8MxD6
X0d85ByVTWUyIo25LrJRq+hOk4of3F6+6vUdXU6T18FKNsfa80F8BJrcOd7X3pvT
xUyobJzngcieF2HE149kgp7GScxhBsAkuOPOg03+wy7vaPL646PZHrU/R7tALkgf
xjqMihdJu7wlT0jAxsouAtro9UmGlIGl6mbEBE7UmcvtrVJK6RoTxPx0v6V6U4LF
vXA1S10HYN9IXTZAmr2GbLQPuUGoFKG9ihCzIFq2vBYX4lrFQi7NCFsIyDzXNAj1
9mOeoqYLWYYXYylhvuARIAJKc+y8teEUKaU0nMrQ8iWYYLcwTLHH8ZIkDnfVvqLb
9o2MERzXLj7yFirah0vCv44EwauSAQ0NPNvPPgfrndln0Tt6Szxx1x7AtYUIUTMD
2rJ7TwPiEk6R0Du1Mh0TBWoFUKKfo7g+Xywb9u35I4ROEXIJN/9AoY2pvCidW9id
dM+6iVfS1ikif3hjwe6VbKFY28Rg9InFGzxnDF4rr8nF0kHBem+bZb6qM9U8wA1c
pB6g4Nja/gRYR1lynhnbvntlbuzOzE/0Y/gAuz27NhZ4jCGtnIMelbvu6sSUl6LS
etGBanrLhc220xbeYmWuqaGSS9BLc3TNxWFoO4BkU4Nz9+gJQ/nidrtM1wdhQ5Qc
icn5J/yRjJVap4/sCWQyEPt5LCroibOhLLOerPlLr30eRjVtSRSr0hTvO0g/sE2C
TFRRGp4CMdRRdpCI4R9StG/MeUlKA6hrPh+pW07lKWHEacAc2vtzRd2Sq5H2r+5m
4LfiLOKS3ovHqGMCITx9v+RPk8nfDlhQUTsct55UUY/bq4z8QiYtjhHg1qiuE9zg
lTIaQScUTT0P2tWoGDbXgvB85DyAW05pqujqkNz/pWtQ0YLuhWH3WC+eti03Q4Z6
EYtOhE4MP/Uc7oNkv0ePK+GmFVQdMDHdQ0zocKzK2ep/7v1rdbd7dADHrLTukN5c
m/H9n/HgtXEK+LGY1nhx9TYVlerazHal86uqHrloUTSTKgVyPxJPjfqZsc2yNyPB
zkJ77n27idhYoyVuGzKv0TCF0aZN1QCb24dclvY1u+zAOwka0+Iv83fEW5iYz3Ye
S2alzkgxqck9cZvKQqXw1U4neXy2yIFmmdc1gQ58L/w/Ez6OxbyoocprtfzJyd75
+NuwnRn5CoI69cPOdVOgN9uGKPMx0oocQFyQ8j4n/bloh+eqkDSR1IGeEGqAnZUg
wC4TKB9/v51e80j05kKgf9YdSma6pSCNb47N0HgRJ6R/EP37Jnj4ocSZfy4ag3YY
+anFas/1e68b9nJGoKe0lfbW/wLg9Kwfs1RARgNbq/IyhdOee6SKLMXKezNfLp5D
PW9M36MsUdHoyJja4jocIzwOjdQ8LEbdRJ4KAOHLhD1hqGILmbS/9JJlYsV/PXu5
Dz2RfaADDWC534FrRSv6m4fPB5D4KLc1sjnYnSqPdDOPyTuZsVl+qMjN3QXoZ1Mn
leWxkk4e5kQ9uFUEYIQsQscYZA03EsVHt/a4auLvjwXcRy/xJUlfuJE/TNO7lW89
bd4ICZm3AcYNtqlXyS0uHhlV9PS6pHF2Ub1tPeH6fwNsGEvVGFqfLxO3sSkxpiV3
zb1lwu4XMgAs7d4wwV0UtL+aujWz7HT0kAjsIilwkhQi8fvnLc5zhKIXzFMTyEQY
uKHD0mqV78/4qRjeZoNB75UeyVjhWfieSwZqm04yv0mCy0y+OHRKxFj9Y+Tgbh8E
iAEOq5UmqUcL5KKBu/i3fOZTm8KhPeI6qZhmF48AcA3KKl08AbsLEr9NcpMU/RNZ
5DXy7oKnNGxwUZV2YBpRLSJVxEHrqP4pEA/YphW/L9PF5LMmST1eA9OhstD+i1gH
SI7dl+FFD7L3Lc0hTAOM8RZW/J8Y6SHY3EDYVtwhJfFNtK4kznMhnEOaxXDCKa1M
6mJ5FL0nTb+OXXwkTq9I3g1k6Tql6YdWYFzR7unHK4VbTFOBnq0Aco2y6iqZ6cYP
AXCCO/tFLK/z2aohW80offEbMYrbXXUE2v++C28pUfepv0hC3JqTpWw9iKMVL0Ec
NHWoQm2FG6oUIhn1fD2r9vv7iql1PXkjvmhQnTwN1MhTfmbc2yvXnojHpWtt865T
L/9y/CTZun8qpnf3HiTf/tKFBtcMJ3t5EP2M5SiGaaR+zh9vkBVSd8yleXA6NgE+
XV95VQnSGUtkY9m4ApvvKCGntiiRqPTA/yQgW5mpdhzX7rZkJ1nNEo1oqrRAjxO6
TOIXe+eLcXOu8/dDi3sauOjaUVL+khD2pelcXW56biYpxEAJG9yOZbXC6Mi77ev8
dAJ9xjAJ9oS7ehEJ2m9qt20NAjymFUsfsXhU9T3v1lqpwloYk9Lden9qEzuf7KBD
Hz8s/CYUMzsyAyem9ivT4xMqr8h4omavWfa1EnBe4Q0IzaUo0ZP1CUEQS04tk9VJ
Ib40Z+xPAY1ueoTMis9D5CJBEqh0BuVz60IbOVfHnOK2oQFxsH+RbCmUvAXYFMDB
MDd0b5VyIQ+MNufBwJkc8App+47/aFNdYYIgf5C2OyF8XCRRan0FJykQ5p/cnLVM
m6msmPsF7sSXj995vUTa8KCcMQsjKpEmMXFNMFXNzN6k7AuyzXGMBJG9U1tMbFWY
6rWHZ8bd61B+KP8jV7ynkBsTVTjswvPT1YjhoNKrWZLZUrUN2C+D2ughW+puUPfM
A49/mO6QGAA+T2f7H3pFOd21vN5KysCquN6LDwzKqQ/jVZK561sP6J9q9dL4igZJ
UD8FuXWKELqbDJKOZAVCJQK7RKu7NFa/cis3Ebjuon92qvasWFjGHYxx4AC+5QiN
D3qOZ5KBAb/xaqBbH0JRb40QJ0TqDtZb+mywPxKYwoznb4FFWtos4l3Jj0ZLuPN4
jZJt9QU/vyT/aIKfuAJf8hwqHOpZJuIdfZCjemooY8aHAwtLrgjTNHXcOP3v3TkX
GuoR5DBuI3Zumt6870QxPtqLf7eRuXKA0BZ8owQ0akvviG0H4ugjAG0KzHv9HLYi
tTfI3iUGfxcGuaxQLiogtazG5YS5KDIjmoFpwHlUT8PlGlNTzy7f2jq++x6Cr14Z
bTlXE+x0bqaBtTa8T3bI7LbwZ1HklJYEkkbQvRGrObKs6F/Krwki1IEbS1fYC441
JxVrL+EKgp3Grs+Ell/+pbMzMZcsmN7F5H59vqyQs5jeU0O3eqZTuu55RgYnJ9wb
R34vx3VBlmc3CKkajPC6md9dPBRrVx59722v3U5ZM+dtcrTYiCU3Wfv1AG+QNKug
BUa4ziIrSP3jtrT5yAtbxUzTEXQpqsyBQdVybSOH90ifUg0zbUXQgERIq4D7bvXx
0TkZPOvIl5yRAjs5TNhb363PRnx/duNvCHHg3z8if1o2RRfLdVrfmdNfy4M5MeZd
PAfyzWFjhKxZ1Wky4ODVguz5xfpOD6MWf2IQ8wdEHLa8bLmfHbgZTuCFu+3MT8ZA
bdsSCWbRpQmO6LkXfAxKOFgHL0lFyDCVfVbD3pNP3+2kyn4/Pzfob7YS5haUuuo7
2A3+ddv0FEQvpvRn6lGsNEF6Wiwx8ZwUBuu8L0cgtGucUEVIGfs4cSXd33V0gld6
jmApQEZb8Ex0mknY/wai5qAKJP7knv9EOxmI2CQoSWmfGpzK1y/sMgwBvjuuQDGM
ix7eNrgu+N6j4DVgI+XeA+YbK8ZFKI8fnxN+IsYDqpaB/QGcknPCQT4st38D6Qfo
1JI1bpmFaRHG4JCeYwmfbZVJNVxWtdSLCOX8JfiXK96nZbShUzHxb5gIxE3ZuC0e
3uDg/63LWpG6R8sJOu30XyRkHgm9j+51CGthdByLHRxRol8TvA/e0+kEazv6kLUV
eTRvAvQ25TAykNe2Pdar8M83V0/boDeQ+XWLZg9bG9yvJo86EEAly4SsPVIJWx0P
CIrJWU9F2M+v5RpQDAc9iENUf3YEkgAmhMDIUUc4t88A/QabFsZVqpWO1rO2Iw/m
JFU+ONu+ZthzvRSs/PTWDE0Endi2wyveuILCD4T3jokuWj8+2jFh6A5Hp2E9B8j8
glT28xIwBNOKqUmIU2j3blncSHuveN/6Ry2HueJ/i0Y09SjiA4w90Z20oBIUU/zM
JCwruUAoAXRtUIIULhX0unwFxAva17dlvQE2D1A010iBnTG99NrDZn24lR61IGs2
aK3bviXZS70BTeVG8LE7YjQEVa0PJa2O0hR/8+ovgs3C8yYa8adRyjXOHZTWRKDD
yEGBUA8b0UsZb1VBDkBLLR9amjRiueEHA7tx4Uq9+aCwXBMqjtc45wuRfIvV2lD4
Fl+apnYpvAcYgtYnxpFdfj2V7dnBFBV97ySkTqhdnliC9MH915PLGppUW1UE024R
w+lVMkqJSyBXNIcOndwkbGgSCZBuNL5/sTcOwDbDWVnqv+imRLr9Ts+BYN/I//+v
KrRnWOVrl10Ir+ay0k2gNxN0mf4vznPlRsV6ZeAGr+0wPR4DwVaFDLq/NNa77sby
SUpJclxquOSVDUbvUShXJOLRyxD9tzafBPNesB7rDQkfCynsvGsU3P/I2MFaxvVV
4DvKVX2NPn5DElpE3FYCQfxNqu0DAcCgQcc7wfHjBli6xL+0+rrbKXzjWBP8tHMZ
GRRTA3SbujAvICo+j97YqSpnyod3/znfkOYIopqR+tCNbl+POqUyr8he7PKnxek9
+xxybvkZWWQkZLEYiVWtpJIxtVaXN8ri+AZA9KfiUVggzU8uDMYZD2kof1ECmejT
HlgfKQ3lD9gFhCk/UKVvtU7VQFtk6SX9leoIWKMoJSton0/wiVM6HUDrwDsagHW2
WGqG2ci+X2SB0cv4GZ6Ij2aIYUZCE37GQJPkc+24vK0q99OaEslfJonCB6yBm1zv
PeT+0Qq1EWxMUbCf1RD+PRU8OTPthi00scZksUv3KIi3y09jSFXILgDrE25Hh3IJ
EPnoPOuS3bQiveXUE91Ksqs6Opz0LihsjOVvLe3hyL0evuuuo6j8FzZF6Gc7IwLi
Dl+VP+LLoVzFFL6Ch+EMMDCnx0kk+1ou1usWawtLOkZB5CxiH0R2aRZ3RtgmZBgg
5LnHGsyvYKwgRDfyeMVVD43M1lhVaVQsM7K6KHfCeS8wv2G2sZweN8PR82hl5qvp
Gslhd7+9hQ+JyX/LIYW7ipyJ1gNX/8PwtVvXt23in9s8+M9woURaUo8N0DHZ55Dg
5se3sfVirHCiiNMHOEemYb3PylEp1YFfoJThTgB4hrqGIAQzwkmcNYfTnHFWO5Po
BzgtBVi7CgPYOPJXkhOxKksLOgC38e64X0gaR8ur7v40fA0DpakTN43mfxd2PPWW
3dPXd0nZqxPnHx0R/3BW6PHaDroH3Aqqs4lmFwgATXmhpZ5GeDEehgjaynnmXJQV
gt4xS8VlCAG3HqdeXs03MvhrpzOnBZEvlISyjOAlv18al00wTBdLTNX2nTvaSNJo
iRGNOQ7kkYIF4v1IMKQgPg7TSFZTFePc0+9xQ2nZy/YJRmP7JSMjnFuGb8fi00ES
7goNkbv8dY5SKP8AJvuGNEP6UV7qE0eJTGT2Q7AjCkz69S4pUXy+a/1MCooYpEmT
sx/FVFF/9W3stfgRCJWkyVAynQWciPrzxQrFwAn6JKbmo0m5m147yGFKBXHiYoZa
aDfrK/l/Xt7/Ei6MX1CJ8GIssaBtBbsSjYglLZL9lcfpnoaCc7/x6pQd92DZWY0F
URi1qSk2D6DuOB9cF2hbpO2WeKvpc5RMOBit0U8Td12vU8gWBt4wXIPWYtHmN3p2
c1n8fge1NAuxSbpHwmRyjfABhgaAH7ERqdyeEIR74DyMqa3WpuHNr+dyQ5OtV8JG
ho5HWKHhurN3Icf9gCbxIVJsTkqF2XdJ5RX/gdpq3CrdagPygt1x9l4sRl8+GLDs
ruPwl3i2ac/oDuWEOkhMTMAUu1PvP+rkAsRqE6YRoVL9HXZk8E2w0fMOqldW86lk
kxTN5+bttQttitT0PcLX6CCS694xQRWpLJdYW36YH4w6k6r3gCercsTCfFuYzEjH
tJQ/hbCLqp2Q9oA4ME/l/Phx6rk/DhHwb4IedWPUxdNBDCobPYP6BdM/8+WlhXFX
IZ2jSBr3aN3RiDgsPWi7gGN9vYPpwdkaXmY/DsOT7w0xd9lML2lzdmmGpSrOf91u
LsqOUVfUZpXwcAY5MpgBY9Kuwkei2kEmV38Kp6kAsMd8AFKtxdz+q34GRD+FeSyg
lIPY0gr+WPxokq3XD/QW0hjv/CE6CVFIfEBuoIGX2mxuM6cV1rSAH6fsvRLX+jbE
k8CTHQdxzma2B285M87GZQ+o6CgRSx+sywJZwIkW95kDFV6YYDRpYSCg3iwj7khJ
pE46kIw97z4lD9Xjjs81dMpsneredGEt7cLb7bAYWNqxiuPG6nxplmLJHdC2GXzF
YxXXqsP6nxxOjXn4IZ240j9VVAeSv4NdeRGuJgBb1Z7fSxkg+so1kDHeKtr8IDd3
MAnQu6DBvGQkgnbS3f53jn8iSzT3z1uN1krbz9oQUIV0e561cAwjtfsyy5YU5/cr
A375rCEviefvjufKBFiHUo8UN74VHiA/poglp4Jp5kzMzbBgpmSAJWAFfHK6WJ6z
QoHLDdUnVbEDD1RWbI+9Yyc4R6oj1a7QmbjNkDoTBEPpe//Zq3ei/8JXWppdIlSU
E0CSW74Jh+Z9GlSeqvfUAJ2efCl5SrWgkoECLJJ0VCqxq/j74dbj9vGUGYGypSFu
f+zGc09sBlcf598KSNKrb+s4K1ltyHZ+ue6dQuV0Bn2T3iMVdv/zLaiNnLDC6eeU
JbB4TQVUceUsTmrAPSw/WXyVYK+bpMSRn3i+drAUZ+JpJLNN4ikc8ddCYToyT2h1
F/MO9lFrjGW0D8uE2enxNyfwXS+2axoGxAX/79gcjNtfRL6Mxfy/I7n5HqdIyk+o
5k6SDN08OZQ8DTTbURMZwgWYzvhNxBwhm/lSre0Qt8fkes9srNdvqD/nNyzCtCfk
2w+vDAJy5nZ4qTzuAirQAkarQPiSw5K4ZYBPNJrGZOznqmqW5mD/SJakWJ2lWaPG
gLONOsd+/QEOC0WH6HfcCL0gcQ0ol1kHM7tIczcoHemRoHWsM///1jMVYr6mao50
GVGjsjalnz6urMrD+EXxs3zYDV4Kpj8DqSzxtVI9kQWaLLV1uMSSj8XK2LadA+6L
3B73BiY0EMeoO/mXrVt+8FK3ZfojqiC+BJZsHMeSaIi/lnMN4tlpsvstxMDss+/U
2FpkETkD5F0CFI6VR+Hmrx0394Fz/5DTsliCt+YLeV1U/cb8mkjv2B/Kp3SYmX9L
bd4cbVzARY5orQV8KLTuXpTidCIPUcac+i1dzyjWUuWLto4LCgiyjuV7PrW7/uJ3
eRnwPhsOnK+72+7HUkelnXr2Iya4lAXPbXtwh5m0FblFmztJOl2dLyKbEBByGM/1
okkNFcltOE8Mw/Bg1lJPb0+J83pL4cUA6DLZhF38HpAlA38wgbRzeIPxKDKnJWIi
hmGM0/x+rNhC08n6A1BZt4YHDoEscbRWfpmy3dZJwiDxv4kk3+9vOizgy37WWFD3
bCYIMi0oQgNVtVF52pu1Jn95m4sJOJ+YYTeqg07Y0dArZPeR9RIi+hFHc01P63Fs
eseOkcp/dwyxUD+hcrejopWA9JcAAfP2fuQJnqPYB3nVnUXXnekoqTdYk3ujBDFl
LAzv0zu1kfaulfFEIU2pQ/DPW7gH6RvwssRDwaFj0qowSXBaiPMT5Nyqa+9LRTcg
W4kqI9q9D9tW4SaMJtmlp3mXZvlTL/Mh6hVnZoq7uF5mnNkUeWPZ4zEi7PaucRq3
/WrKhdDtKmMpTVOTjD2ltuTdjLiYs0wL2NP3z0lohWJz1u+qqgKNoUI5OUeOiR9W
dANsC6eoeyqzlIuJuQLblD1U5en4vUWdLn/ymxqvAsHtuBnKNiazz2nN77TFnWKX
KQ4aTNps2WCkciG1ll3B2QDtJ/KSHQuhd5LEQijGtjkCOKLzK0Y2uV/1VIy/keF0
2zb9YerkiWgEbrAS++ptTCG9LNAMzMLQY7Iqu59xCBO/JcGxt19BTSHImnWnj+xX
zq+o7bthV4p8sFfmSKRH3xz3e44e0NeMmXhTTNi8l1/jDHkCQ9W8Yv2ePtgRkxUG
rNz2Dj40QtkUcf046Ciw2EGZ+EbrUdei0IPOxpVNoFr2jvisPyGUEBn61FyiApmP
HIY9Xuy6U+llykrziPqtbbaYU0+/GNjUGKgL/ftVrrbFLAvMhpQdFIiLSxCgpZvu
j8Ookcl7ivcK7KnU7kK6Zz/E0pcrnf+nYGNMG4WVVrs1O8xtO805k5rPA8U5I+tG
4H8bGk6J1OisDRDznEWgPE0ifX3Sh2AZP3rniNKsEVDd4OxSRUrb2m1iGLhQb17h
8iqspgDRL3Nq2/SwU+l0zHsOkAWSx7MMXC8hL2fM4mjnMFi7/voZIT/y+m1hWioH
WajjN77RZfWE2lCVXdlSsFQXcY+acOOmTodesLbZtI54FOcu620bAr5u2nlvMRlW
0fXW55sCsVWWVeru5QgeRO56VlTRWcdE+OgfrcVW3BI4GgAmpZGFgqOXclFrRc3Z
H09DQs03c1/7AO7OCoSkpLxLhQ722J8chwq1BtkwWCgPYOQ4QQmA36BDqB16imMG
0FIsXMCvCJKHmljPwUM2Cf59SExX3vlxDOiYdI/cOc66r2yc1JrDLKqVOmx7IKGr
zDcUyyWbFtH4dsUnhGibQO7ghYSJ5E2pRj6YhAO61vUF1/X/v1KNuUyzX2pa0sWR
07J4oA7P0OAC0Rbdx6BiUKYIMAEEHJfdXrVPbqiq2F//7Q+Y/HG/Q9b3+yVcFmRv
syhpiPdVgwcHqS8v+rZtqKqW+dGbOO5jbdiI268Dma+pHhPbf8lLshSCnKsXuTP4
o6tKt6CLby6WINhxTARumrqTZ6fDs3aJlWpTTszy7R+PJ4OCLxkO4kDgPAJo/5Qg
d2VogMyr344YGZlWCVkfqYTck6mUMOnno2dwxU1x2UDuu6CRPqQ+9SKGIOrBdf7w
3fMYdMekitkgzcWC70YitIKFt7vAwsgUHUUHFHJ2wZi9MZxLp5dg2DB5KDFETRIK
pnAP3xoWSG6ArZFmT735jNGcgjCBDixJwbMT78m97Sw0HzKC2REZ2ybc/C+opBH7
UqWh52d0qeyCiKy+OWglbbeQ5n6x5BRVaSYDVflWo9FcOs9H2bi1FVN8TBOIgDUX
AcvyWDc2g/EhNQZsTlw6GZOtpX4YbED18pt8TB6j7Z47aiTXjSyqgoSKOWPOIjYc
vrJUTLCaO0GrbOJV7Wzax3K1LOwFN9n8n/xQV8nhJZ4btmQTlaf8oU7XDs09szZZ
hyNUrhNBATjMh7TX/LcT5s+dpXo/Y3iy093KG3pLHuGa1o204fuxw2ANPrq3RdKI
y7sQiCzsdXTM1P+VRt1TA3pTiP0jb6m4B+Lsra5K9BxlCAzpT1OWE2+HZzG3BoKo
A0uAf7uU7oMJWzHr9Z4PjOrkSl6a2FmedNZCmdnTC7T/e3BR0bqG4Jdh3I84Nb2l
ObixGcBtCGPHoseUStvV0Lhf/hPJlEWeRbL4oaBhPZup2dXw/KpxcG83K08oHaVP
Dj64lABE5NxYCtLj5An+vgCeH03n4viaCG7nEVKC626EUQ9jAkCpGF3srAY/8y0q
Pwt3Cj7SPrXkUY7nViel+dUMDPxm2/W3uvSETSa+/kd+BsMBG3s/pVhWc41BuJ0R
yriXGiwTw9Hmp1HEAuq6Z4z/fEeZvsV2Lvf+2Fx1xaHSayxe5Okckb9RFIHr5RQ8
frfF8jtlkL3yTEeaAyRZdovTEVQZ1pgtnMjvpbNMZQgwg+VU1t2QTYOwL/lVJaLa
tzEZELbnsfqRzqrI3u1oA45FVVQWwvNIMemFTNOlaVcUUOSO7BkYw6to6yq+w/p7
7ZDVbnN4i5jwJKmFM+Xh3uiZVAo/TycqllfCczULuD6GIQIwC136cSY96j9g6Ksy
umbGg+B+EFMoAU86cfUo2bcZRnWXKG2wk7JI1KR5rD1xLEwjo57K8Q8Bi6YITD/b
ujhPCza1bMc8uWtxzzyvNTZlKXTwqxumtdHib9QSKA1lO8t6LBCDwZIOIdRzBQ6+
oQ7Hc8cLMf1rqSxaZSdoXysVyd47KPkgz/r5lxZ1lvTJLJBuE7jJH6Y30FN8sNlP
t5DUvbhfwvmWxAQ+q8l/S1Jb5LETmgenh0FPer6CCPbCDUH110v65x+XZRt/sQZN
EM/Ydg8RbIr8OtEe8LTj9xc99gao306bASaUeHuZNWQ82MY5wQCym5FzXHdI0ptK
D/Hzo5V9AJzN+ZTBLBDRMXyarflcLBan+QX49mtb1W1iIQMTowuLqPaymKnd2PlF
6MyQdQJbqe2ntXLTlmPTy2J31oipBM65rXL1A5J/HDvwBHhh27HhH78/BG8R4RUp
K/1wU8JaHIqOcvworcjcp3fUPLuL6+mQqdS+UaXVT1/8rKA9DmHdJW/UlmeBvf+r
Lyw/qBM8QlL2AwsmZKSEOhwqnw0UUKTiSy7Ef2sVMyuiq+XqO7WA0pqUWv81F6aH
WDmTt3A3BPyeOn1ZPtw7l/1+RN6boUPlDr57KdLLtUm202yQ5ncstcxGa3fURXR1
uIY2exBkMOw6/vgtMg/cS5oPlSSQ2wAA5HcHUJiURgTfOxq5s6uSIAGovR3m4pwr
qa8t1x9Xi0LYF8vs97W4qXMGB8EyjrkK4/IWWKCnYEX2qs7TtL9HtmprIhp6GXku
/3co48gpD2+bg5f+2MUendftUh3U99i0LIPTMKsEQLinYgpFbz3zthnVRuzzX327
RhLMGu97RtzqkqDfV8sxxV6Pv4EVACMwERcl9QL3pabcsq17n4fyfqI+ziUFHfbE
bMLuy5gUmLUJVpJCWb48tsOy4VhFWmRSVOK+2pdH2ZbiE6Zzu6Gf9/kC1pu6/QrS
1bitsIx7qw4RSeGeEfwnR5oRjjyV2l1DO1qsllkLxvYGTuPu9sjhkktdqYPxJEzi
eb1FwbubSx9pnorBjHoSMhr9F5UdrnncIe/clJvquiCvDegWl2buMGoRUv0tHfEu
GWx0t27B1PY/21AWyzG69oOCjc8UTFoqnUQ6P57JE0UMIokj9+wNEt9MRA/fqsFU
WnpfWxTNDUhuuhy4f6py2b5CsY4C9MXQPoBJ72bl4rRN76ABfQKYLtGITVsuKteo
oBI7wTDJk0Mi6Hb/avItjuFCJEwu1kedBgYLWuy9+zquQBPNhPzfLtiwSbW4MxQG
3CvSQltT/IRcqKAW/mgAaIIsnWjipdn1KvVvRiMJ93jq1gjBP810izY9mOMBOurJ
A/+2kgsTKHC4jSQz4aeNMAEwJpV22+YH9TsCJ2PlgvIdF3EYe6g3ri+qf2E/ql0q
lHsiwdKfoCB4oOFKYQFKP4denM8NikOJ/rnxF69unW9+AaWsNBrKyL56Y+hIj1qa
qSdMQrIx8QjKuEHAUQHBlZtdEPEFedynZXfXmLk4z58yKSL9PPMtVc7aKqC1JusJ
BtbVjrpnj0ZpVhtXhaI4M37bAFIv0mn7pVzXCtTWk9d37nczMyY7GeXZw2oP7Qq5
MTUlXC0e/1MUZ7EuT9rOngk1q0pwPyWPDZQPjDi8mcU9j1T+LT/yxsI1VbxtVBst
ryUdip/rseUouiMdtgUdULRzD2aoCZ6fs+TeDSqe+Y/6uGsK+C4IJiiLWpIxi2Nl
/bbVelsFzDBUIiZ2QLr/2xr+xbQGsWQoMMd344vShoE62TMo6WDH16SrYxp3N5Xx
ALCKtW/nkEIqOC15dk+5Qt7tppFzAcpIIgL5Eh44cpuOA4UckMO69Wkpw4PpXEyU
KjrUiWKsN/LmZRfwr8MB2243l624+DSibrc8zsi9dMFwCgTqHqEcurZj1yvn/Gz8
hKNmv3WcqXEt0HV8C7izF9J+EzkMw5JtGgGwntNMV3mJGD/F4gtIa18Uu0W+yTzb
hc3p7xiEQ1kuO23e9baxWD82ywpa8zX0JomoSqKex5pd05OgdAZA3KxIGpgFPHly
fLubTfGP6HbHG5pF39hucMRNHY8EUL2tNBgy51ch29wLtCxFmMLOGfzgJWRcN66z
uZbZa4S4KXvDNAgMUAwY2V73PRaBYjPFAX0fPqVQue8fs2YaRjTWMcgGLyLAqM8p
xzbQZxvn1vsHQykjKGxT+1lFD5ClwTiWVeX1D7xeg2Hz+FDswTyBUZoLr51v/HhP
YdpKIUAm8g8QJNbLLv/IwRqS9KkTlHstJwMu9H0KmT3a0zZXcvoDTpsrfNbuAoq4
Gt6mT8cJmd9Jh58ucKiQAjXnAsBL5Ub90p2VjLDimrByTVLG4OGw3M7oHUgrKA/o
pJQv47lCn5crLv0L4w0LF1gWfLGfcpMnFoPUW0hh/aecHL3Wz83hqaUKlhDWC3KH
tK5utveA07ZHV+lW4tT+mR/GjOyd6dl4A1L5gx/htwRMGw+TWT/uBtsMyxC9bDYA
zvnUB6yqFPawLLA4VnEmCO3Pnu1fs7lO8bSwgKZS/9cLWgdaIBgjnAQe64ViLDpo
ZdpdVBc707BT49+6WHrIFmBYLcd/OQOZeUvkj7j3X49jsRRiGqEzNEW/b6SpGVUg
I7vx8pqkoc+AiUCYhIgw1V4DCKUMJLEKNb4JQ4EIRLl3ApszOjSyz9g43SYYMssd
0g+gjFk4MSO//3sIdlc5o+c0GnBrNMbkV3TTi81MBFRFUDze+Sf04YhoZ+yM8iI6
TX83dETx9ZNx2XKqHWJ7hWEe+6RwCF5U+CVHe8qaAP7HnlhAKhixyx5HhBTirJwG
y8B2U/HgjHwPqMzPR2HDx2kYhTbAOvQddlEkqiybFdUxXgjIqk4OUzjL++tJPvHv
1PiN5BJMzwDrCLKTEz8sMv7PC3mk76pFSChUyQ+asW+oIMt+K2bcchLl0Q3n+yDY
Y3B/D8zKP+mlKb0GwwuJdg01Pk+1EElnRDODUfkfQIT0uIdpVx6wYWq1Os4BPpqC
K8rbF68gJB45ZvPS4/bIrkoukIMEIwHebJ5+n/FiKW4I3+xaU4QutnUvEVPlUwyf
f1hGNVxZpTcwBMJLlxYETk85Knrc5due6mHonlxiLLuc5EX0bvz1MDUxbJglr2tl
TpzNTwADENaAq+wSkgLxU6cJDJS187McceSa1YSmqBPDwePGpvIFUe91jdpLd4T7
msw5aR+kk6H337D9t5w8I87WqHpUiv429Y7hIl8c6y7BPCo98zXgP2lwQq/DJNjK
LTWPyxVe2urtJFpzPJr8jDDddSjI0XjqhFt3I0XU1+btJ0lr6q8C1wFzsK9pAwM0
SsjR6Us+XxM19AOSzmLBzXjlA2bqFxj255rcYkZgGqL8v4ro85CaskNBVSDHKN8H
rSFmpC1LfjYf0hDD+BirKJr3VFz0pZC2vpa6giJnEfZi9LlcFtPmyD8FDYrdeX9k
agdum4vcf7CS3r6U0rFRs372IRlAf8s87V4IiYSNWxE/1k2WrBYaYHWVflpDJGaQ
ZOgk2x4mzdwup3MCeGB/8Ef0YZwzed43aZqduyR0QvGp3FSWjpT3giRBwXe0Aj+b
rjzENuWN3WOD8oUwHMzM51YfwqmH4COifqm28MG92PatmFRRW4x0ZkYvuy+AuYh/
jRgebL0k2IFNKN5GYlUf1Dl6snXN3hzG/yKlDoF1BeBw/lVYVdEWG7ppuX409m/2
GuHCw0NXdXP5ogtKzpbr+poSa7I0kLbphLZuM6Vr5As9LCIPST/wweWn8QDlczw1
CqZ1WUxovWmwdN85NlOjZFwbTMJNwDPBBIoLJHg4yyIrb7A06fVzCdgbhlYKIwSy
dWXjxpQ2dGrEqEvY6xvGF3RDnuLrh+p3WyX9bJa8E5HPXrVvMra19BowgFBp5wQ2
maDN3THr1hKLVNW0QwulaxvWbw11W93jp5++GVZRWt1zlqHdFCujvQTuhU0er28z
7PppUm0iyDC3sr+TRQynxlqQ8idmLqjTPrH8LcFcivfCQzDhueEtQkl3BnMZjDsr
wsgsmntKWtK70dwhUl4gkz2qX2UcSkTNCEmiiQytho6lon1HL9SAbj8alTGbeR64
oTwyKNA0zjKtS7G7LSCYQHtM/RIh9iypk7/tCy12j9A9OqS5OYHUycd0WpombKLG
XWDke7hK/oPJZs7+4mZl5ROPj13YOhbVoARlyEnpIfiSCnWbv1Q7LoT8vmpbdyz2
i7sbV0aesOA4rKmtu4qhymJ0d0/KI9NhRmXu4NU1QpDR/eTTSpS1qliOdXiSXQth
Dt+6jgwl9w/mzhEizs6v1kp0SjepfjVJz+J8DUfz5NxvkBFz/uoKEIl1gH+gbQG6
f96PyW4EmT/+M9YpSp35EUJ5AgP9x1o0dxR5xPR7zRvhCCvObnTh0hAoWXE1y2ut
7XZMU6HvRno4GVUgsHPzK119szBdBTglQspuLfESzSLEMkdmMPjVFg8SO10BQIAY
ZOu3tpmrE7+vjOXQlgglnrvIOAJ8ApywBC/ZfDl/aqHDLCJF3CQQzzx9uqTzAtth
APU9dkjTS3RZSNKjiDimX/S02lG117iz6gf6llrSKCQRgezVucZ+oeC6kUPDTLm4
ooXj0gT6SfBDkWbIzJbOzDq833s3X+xMEJqly/uF+k74GvOxVYRZss5xoqAwXJ2Z
zujf6d0mBnKErI9dDq6qi/qLWooziVqoAPxrilQ7lyIClCBmx9rm9kik+yYIxtu8
oheCWrCIXgCsrU3HHclz+yzjgOnepPSvc5WPdYFH8Irtx/4AOQH/xpkyof95th4a
P21bo5ZFfVLb8nJh1fmTS4U7wcWt7cHgfW7dh7XqDJnkbJq00xSmxP/nSRtfPo/X
Y3otaz/GRTkvJlTjyncM1neZmzy9M6VDI+FcSkxS1dxNcXOHdIozd2Z4AKC6mIPP
cTF5fybrsqPBwgSQszbJAqyCzG3Awf5oJEIs0JMI7oCXOX3n1aLAbLV+pFeVg60p
wiJBLksSIO+FDV1Srj3zX2ijrmxlpqCHJ/taZq3enIifazV7BVQdCOUBlTO37X7J
QxQO/P6ZRE16pK9Z4v3xt6+5zBP8FU7ZEJ8LvV1iUyOvec9gqd13pabcJbP+sSUF
DQ8CFFvWmTeDpZvbAs+wKK1LkfSwsVirE3oO7CetNO+cjotWKbPfi8f3Zy1/y/K3
fO5s5wyWLXjjcHSSmwEbqmIjS3GXuhnyviwsMNtw8QWSX+PttkTdzbX7jvOcUdnK
jwwWwcVZhR0QWiUfXfgQsWRRRYT776S4cgLGMlRAfM9PEwbpzXpcbvBkYqfoswAr
FRVEItsJqfa7Ogk67ZH0yGnd0Ngn0l3+hnDllHMXHLg98VtD5OBpIgpMr/FlWhow
u+aF6jzhJmusEmmLET4ioIyXIAIgBoJcAKc83WASPPbDo6FeYZBl6lNwtydFtbXl
qwxLb+x9M35xHOugjYyjZXhFJJSJAvwh8bJhFE7yav9x4myL/pjXW3qZH4WT9ogm
3nfOQyrJOlOQTy2+IhjK2yBY5YtAqnkUJvHp0hMZ8RS76VdpHBUNbhNH2K8rXO6t
1o/NRv1cpP2ouCxYwqucisjBChYPWlf5Q7VoDCG0TVui4hW8j+qhe7BZm6fmSkEZ
41w3WhSJoHvTNK8aRA2+0nKiuw4JDAZlugjDipY1Tpr2vZBm6cG8OIqIxcJMlugQ
UV9hxowwe6Spd4ogpbj9lnpPRZEKankiiXuIqh1h9Q+IfzGtw4mhIOSuWzEPLcF9
vjDipoZXrM3JnQcv+UyfZCUTDIhgHxlKY1ZaOSonCcvpqeno3Y1C5efl/Ly7beR/
pPkEQ/PJrQeo2FkYGbl6/WZF9GAPz2+rCbFn1p0nFkeJlXKFEmPApI5N0dLmFD+A
fRNnLkA1bQfC5jQhDs1FxLhDnC9CYBNGD4KOtoiO0GP1dXn8T0oVsnqKa8Lsbpox
vPbEqo0zbd9YcnCbYp+684hDMbiD5gzFTt/v3ITSGM0TKJVqOiVrCvnmEU+VZxuO
1Vxt2JsBozH4O8l+epjZ1AMxtdtBkue1b+s1umuIcT6ptJEPno8RyaeM+5mcB1Et
9c6onwEaki601JzFmoQwjAE2wIqtT+p5PG1ilmDe088LsojPLgtm/jNCOW+VtY5a
tjYxeCckIg2cwYeiyWLEI6wfXDTkb8jds09wQRlsXeup9JP4pmFBR2sQkXMWMgs3
kZN1VaoIjjJoIuLpb83b9qkUX8Qc0wByV+NoJddeaEfCwokBtvms3zGhIWdLI6zV
Ei6kpg5juw1jCCwQiNaxkwZf1+3YnMdgb7bhQIErey7ZI+sP43RC0JkQ3CvivzF8
Ekh2ZscevLoRRGxhBqelQF0pLvi/LYcRGZ+iRaFSUAheXaHrgBF26dzF5FgUOTLg
YLYME2eG8EPUl9/Hucf28vX0IHop9j6IGIKbmPjEH5wrXPmVk2u+hRbW5/zzVt3T
jOrwYQtNKxzka9gyFIn3BZrZVBgtyQVIPcv5RJvV3jZ/5peRFmTl9dionzM0bw3v
LH75IEEm499ZGo24QGSXxhclQ/zjwPMnft2wFEO/s8RoRdN/J9hF9ZK5ZNnoP6Nj
tcuUpGwsJ4g0yvqtn8VPU5me+KVKpbbTecLXLTDtUr7g6/aiVZg5HFI1LDu1JTbx
2Etky+axAnQAdh0rqdcOgfqCT3kcfbQ6PVVCntlfSCNQ+3oxr8IEBKKmP7B8xcUE
LQcxvdUX1c7fX/1CVd9QFySFsoAEP24vR1Jk0rfVgf/5Fx9ZeWvfMlRxXkMqwJgS
i11O9PiSpUHuTlwtGpksuce29OLGCj9glZfEHWbddjjG7W3GjFRsFI11PT25Zu8k
r4S4M6egO9n06tQaBEHO/ioWDUma4Nw1flo4cx+63Lv9i+eIcILPxfdwa9h0CgLK
F6bswBxvrMIjwc++wxdLPtX3/fnVvclttjZD7sIUdcKY3T+0mR1K7s+yfmBSjFH3
WVAsz5YP8Mp/ZFJ3K6l6Yl5nmGtFs3kBBF20T88iwNYmYr7crRDL1mUdfBe82Mm2
d+0PTePVlxF/8S6uJx8mB2xHJv0rW1he3nUH3E4pVoKHPydKPyU9yMkpnG1glyFr
luT2fMvwoKeMakuBs4eoANMs1wYce3maFzKbAoKPnvRCxN8ZCptWAq4M1ZUi9mvl
0rMpIvd1RrEsf4ijojDZqhguEfsBt9TgCPUmlmOeaGYAmLBMq4RMCqBhlu+7X014
XHa3/mF6gHVP+YMPfOzN2tmbT1IEKzokHf3ZAUP7QiL7DaElClQ/FbocCt3fxfMI
P0m9l787aKFOSlpFaYTgMxRGdR3Gz58JFv8iVZzqFe9OiocXEGBEnb3/VGmoVHve
XZp9r//0dcujo3MVFnz3puf1G5ix/vPBvkDZ8N3feiiObagO9xCZnFIhMB5LfVQU
igruyzMtLuBtviy6ifGQz5XbvTOea0MEn+wIJUmMRlP6oxvta7miPyv+2w+yG4b6
9B/AmuXqgvjutokxnb5R2/Ff8GYXDFsMyiHTV0v+di67q+k7FAmNnWr4IF6fEDhh
0pby8FRwZZT9qw+gk7SDaYnFUnqWgBkt3IJVqpwrpb6FTCMUPrQ7ya1FkewRAx2l
f9gNaeBTS5t0W8ncsCL7ylqQrmPatFK3P0MRFvanrbfwzT3ijck7TM/QkkMm44up
CxAd2Zy1YKGwX5JHiFLu6VItr1MLpkXBHMB0bk5itGYs8aWpwqZ/nKXIofUzP7vg
L6TfPKjoL4nUKshvK1pd8nRm1HHEP8MYpos2m1dV4Vw29L0TnfvDy0NR94VGbdcp
W3o4RxYoegsFApdhmsz8gCH92xdSICxm5PHpvHnxmzxE0ykb265sStF7MvPb3hN0
eEUWlWOjZh1WHfuDiqEpH4A6q1xA2QTJXg9BcJRo/jmXHHROGrwR4b/LqOt/y6/N
hMtbzxOe5ernR5CAu5sDsrrgVLah0qohglm/w7kwnyHjPDZzZn3h99etLBpKL6up
zz0TFWEVA2m6UHkJZDBuf0dzl7GttDzDxH1V1uPs29VX7E/5MpfobPaPYgy950gn
HdiTRQaZIQaEBoTSbrYdaqIAWHdV0Fdp5RjlNebPKfJbLDus5vsZAWCEcuNoT9k/
83skX9fWmZU1jN9V2Qak9vSCETA4RfxWAsyUzTP/zalx30x4P+gBeGGMW9JaexxI
yyOoa/1vLjlI9FxilnYPY2tEdqAF0NVcleHMWAc3dZt4dD4YK1IYDNWVAYdM5RHo
RsGOmfOUuyjwtmwoUQPKfU07wfWNgHL5MJmcyYXYSYwsF0PyoI69qYpq2vhocOlq
cPTz1GKIeRGWf2uXYd/gbNiNvgM7fC7XxX34Kfvn/JhuWsxvm2I8tZNwJEbmvHxI
xICLXopHhjUuilE+Do6FtGXcNgXZlrLXjWT5fz+9UCgk2VoaGdK/FZJRrr9Bh5Xg
Ey8j10MYq7EucArs8a6Zcy9enmnCA5ISFheHiKOrSACk0p/GLnhoDOCDNdPmGkfp
C7oV4YE6aawSQ/VJ85bRFdB+BXKgWuFrdFUw2Fwvx9vcgXftbETvIC4C0K1bVmeY
lYloPIxea0uNnvhb5pkua2xuihYup1NGWoZJ4aJiaAzo7hAKorkw3zdQB1DcyMt6
mqXgkgNWC8/yn7TORwN/ZgqvT1a/2uYJfYJkyOBIujrNouDS3BR2okjBdVJIf8mh
AGaWyZ9aEUMY2kuFp+qf1qsZlhYYlYspteSoiA8W6gWNOYoMQxR9MglKXonDwtWV
S2jNW0azX60L6VbWFLMJM2/HoOe4s+uEBaxdNXpp0DgUi7oipICY3g3MAiSKS0Nh
ZR3vBbz18wCxvNWDXsfde6il7dwbUBhRXUtz4ewtrIl2qU6msoJPgrQP0525g2Y/
oGlTp0f4jjSkE8/+lKf/PPU1K+KzgmuNnAyDVGcbF4tF8u7v3v4QswvxtI2RAEy3
8jBMol6pSBE8d8lCJKTKqzm9NhSz5Cu95enjXzH4s5OaY/j8Y89HNBqWQeoRVpnE
+tIL+cMS2YBY1sztGnNk9ilf/WCYyYuVm8vBqh6WEVRBCOii4vtsCd1I1dz8UA0A
FK/XGVuv+WvXIFtA7NrJVlJMyty4OFnF5ZhZwpBx1rTIQma2X+7qExZrGUziRJgO
+iXC98yDd7/3zrS54RHEaOJwBxQA+yRh9W0E8MoQP8JNCQnVDRVrVbKziqTITtKc
Z6cblH4S7lP6Z8mQa23rJ4xAbSx7GeJCG4nWdYz3p3mkFgLdZ8QG+tvV15KoYOva
7URAiMkj+HzbH94dhhW/jmuS2uG6lAr/1uxQ7d3eGwwJxHuFTVwe3AerOG/XJAXO
k+c0lC4Mv9VWoNJcKNvNZAV8aFZAlDoUKWEmMiD3epZ7RABnjgbnrHV836q3LlSC
UhkZjO6ga4Z0D4sJePFbtQgLhMq6BG2ZdPNKhVZQ9yRlhk1hBhsUqCKZwPiRpJG9
IGY0trgeaZrnNvKfyq2hKPEK/4WzdcfWhb0IIlLAcz6KMIsGuDKgxVr30QHTy6AS
oCB0kr+WZhAHnQZzDC+MrCajTgRouYfgOCUMKzfPqJE8bqQZNFhZUBV/y3qSr3AY
w7Ccovsnp4J2hvhnyoL1D8NkM1RvI3J+WeLU+FjroRTMTLbARKF1eRNSm7nUjmWg
1Q8wPC2FBp67IRLvnuqaj/PMUg+8ZvS99mZgtVmUFHUwCT3WQZoy/sQQmz8YrIrC
QmCh5P3QKagLtDFzWap87bdZVv29sz8Gb9dqBn18OI/fzIKgOrA49XFXJOVeX9v9
PJUwyHvGk9gHlc5eWksPWnicmaQ7YpWP8dh1H5XM2MkpnHnnhmEu9bNJHP4BfPcf
+caB5WKyxWW80EUj2mpPCm0Np45f972a8Jg/hZ7o17FBbYjnzmPVvy4kfvVdXYjg
CN9SRNuPo7+4ftl+56L8AobZrULlZ0jpw62iiZzJ45fjyhzFySJmOQw6wppUN5fK
D2OQ1Nc4/e3kTFIzyTSSPCIryl17JrnU4IYWvTujG/VQ04s/Mgqal+CIoCChgqYq
ZnfKbp1tafL1NtFpm/BEcbQD3b3KDxpXOqS7QR1wfzsUFDXDFgtFBpJsbq3jFrOd
4y8/6JJfbPJHpYEUyVhWvhmBk6BLv3489XHY8A/fKWnhtvGi1e9mK2/otpo6dOrB
ihIfDurRpZv89ah07kjtDwZhm0H6wlX/sM5yaqbr4LmvkOHXLNU9IsIsyYrhfEh4
10L+C4b3POb+/sRh0uv2NzbTJD14hJvMCKodP5bgbiuExFj6vPpIT9bggWVQ2pJF
dOkROEUUL6F+tjJbYX7lTZM2Lei21GrYSOxgQGI08+aVI4j6rWeTgBJtSD73PGBX
m1Tas+AKzSsA716G289duJSp8oqNbjp8qIAcJjFU0rhn0unjknuJjb4/gz7zk4Vi
Kq8UK4+pSQafp7qNw0WhUcwLpV4ulA1gEgxkYZ9GW/Yts6WilHeBXkhrTgjpfTx+
ICqpN1k6iumCmg+2G/OT82ns7s+A3PuvgvE1Wc/LCEBOD7G20w/C3qU+Njj2tk4l
LYZYLJTLfEfI7Y1I+zI2a2UHhEgrf/kfTilmh4FWyRSBwP4Y008QPGHyV9poSU4y
ah6fReNgrI4+ZeJ+lkwT2WjhhqRD138E/q+BgjcAQfn0aQErgp8z4BKgekSx6NK8
SqQub3pfQavjVdZUCbEtx1rLrf6SXFNMRrTdXRqIM8WZUUR0yOfuAZMvpUqDkeGp
8fRh8iYSn0+St85nb5Jo1fuJUAikJZvaP+arGYNnIYMD1h+tPVuONiWMJ8TzPSWB
34/ClYK8CLKTznlk7CgyZOEDRY1YxSHnRqdlA4UZawVgTZG2BGo86x9SvHzaZP8f
s2SAl82TqOkhJZeiIzfVCqJeD3YFnKJ9gF685CLpm6Uh7+K9+a5E/SS2Aa5uUQ1s
V7ZtzF09DdPlLt+LyUooJAQhcmn496nuItAVP9lF8wa6ePW/q6zo879bHJhD4008
3PzFwo33gP7H1mpyO/rkt+iAbKUT3TMH0QMl+dHUKwoyWlE2OSUytjsU/wyqVcR8
rprG4kvgePBGmR2GsORomtKTsjPzvqfPPPW3NafJdeD3z2TQ+2S44zRXLGjBg105
SlNeDTaBrHoEUuuk4s1qJY5FLHlWUt8q8ZDIp2SDWxIOiXH+Q3dme9MtwUcoUuoh
h40vRHp7Gi5nAKYYOSx1/QGyYiJAb+WP42iiICMRR1cygVqyj2GXhzngRWBYuMxU
F+Yh9f5vey7vkI1NFRDMzE1DzbcxdDUWLjFNoulsJrktde/FitHg044zNdaXHaNu
29xqw4HROYak3Rj3WlTiG77TKR0tjYy7hA48humk4SiStYS08cTWBHiUKDQWF6v9
poMfwnjp15cvSyH3fVtb9HWM6q40jFZpyCSSETkpYsnunOQGHWMlMWbUe0Avlloy
UoyX7YPHgRwc+alFp/YkTgcHBg4RHUgpMvBmXg0JIEltVHJlRbhB27bjDyQ1c6C+
SiUck3qqndPp5VDLYRbduNohu88LEo6XAki3lljaraCxJITvsc8F0EHDCBi8f+Uj
KPPW/nQijgmuWW5WeSfz9/AAkFqGa3GT19C+uDD3XMinKatMx+dhb+wBcJx+JyKc
LJY3VC1394I6FmoVe7p9MRoGRYVHE9EAHwfZS5lF4AB7mYjtEMuQ5e7bbu9YXUJg
4DCMFXXnUIYOodwxe4x8D7g5+spWKH+eTfWJKdYNzttAr6c8xp9c4Zfb/u3KeIie
VGAaV8rKpYzWl/zBvJMV0HJSRkStaHnW5wmgyIpoJWNRi0UvkSfaqOckHTEFvCpj
7145lYmHmY8UMgdH7TC8C6aKYc0av4PoIcr7kmqfWe80O6X9u6LVlk3KI5iSWXEJ
4KYu0gMIp1Hg7PWN6U6TfpHqQ/R7Dr67OtugwTFMkKoDjSCTrIvHr1kBUBnFb9Lw
9Vj5dDVNQaKEX4h9F2Fw4IJZ7J/HTT9Pgv6phwSdBQ380waNAcigI6iK8m6Lh9qs
sCe9nhybAnR7YCv+iKLVbhAFrZ4RhGlPNK+SvVFdFHyegQeKIaDt5ubFodwfB5pB
bl0lkPjHmjAF2IZrxqZ18DTNi5DZdAe9VBIt7p3G40Maf2ABZYCTBK6xKJOhhAgP
XEg8G8tNUR5CPZaDosKN+HvFylelL3jKLnUiYq7vmOoBY8/srjEf86fRB5ogkTtF
TVwkSg+JjR1ntuDEp5XBE5Gi8pXTGjzWthhv9H3BwSfbuOzjyVgXRHRbo2jVpPvj
cygfv3TeqGctO2INlKgsLdWzLsZjvQ9jC4/hlZFREJFPr37c/AoLLzMX5dhe9kk2
2l2lmnvlaGP1B/KlCyt8XXq4oVYYmMRV4EopBfUCt9r8s4rww69EqNeDftz+kHp5
pxhDD0DRvFfeow0c+6CTal6zRtYMDNrrh20esNY0nbn6l7SR6ZeO1SLKqFRrjCBo
kJC11gJHVk63xfQM4w3hznUY8BRivZAfCWMzDkciH6mGzGt07P87/8VKNe05Bubu
iADwtQ4KKdO4dZlbA19QYDFvNyuazQXJQtkGiUOFoonPu2HkHSOAT/HI99SAmi9l
Np79YPqi2vI5DrXGKGrGsGAyez29ZhwTpSH8tNAXBza2cOV9XiHDOScZxwCtA5yD
7um5dXgN1slo3PUU32ffFPxhP7ZG0v0RKRI+WVST9mLgLQogE6U/00BMZFeFPUa4
mEuK9QJDehcgp/TCBWOVnMEEa77vGpRIL76StbfN0C1s+iwae9yeuyDxwzGzJNQd
el0NCdADmSNQIj5wsM91yM9oPmkvW5duKfXrfv+/Pq50X4XU8o1EcCiW8vtsRtZo
FDUZXiTAxiIRfYUJ6PhJ3WS+F6sl0d7Ob4qtlTHu4MaaZ6YB7epQCaFmhhKBJbZP
/YUvkunx7a4yHCsfMEltbksl0jOawviMYgSHWBR96awZ3DaplUin0Rj2LG0sFxaB
r28vrsBv8GtgJfBW4wedWCEVfAatkDOYB9O5msZuHyAaiV0Mh00EdAu+ZXsZ4yCK
UcVDhCkXUjDVvnHbhaE0kLwqB9qa3/0IQy14MOfvF4a1VN+cMcx4ppWDOUk28Xnz
DSGLY6IhegcRAf2UllOPbOqkytrvVXBqZm+ziBwVksxSyTWE6PTQlQzcURSd4xn/
WCKfdosjZJ4YOe/dOfE25j10wwzaK60nSXAAs6tXZaIyIqD3r6BAeE4xRcyVbdd9
nUwZWQh3S/CHcKtWTJr3uRJ//Oi7G6uTHFW48MMfH5wQ7MsjXJ0LzfDyGAd9bdag
kAt6iJ9cLp0Ybo7M+YMTODvA8fr9NyNj52BrcuywwglPvYtFhvExD6WNEQcARjQ8
Z2V4VopOqEtUd+dP03H55o92QuKzg6sBWnQ0aqKhIl4hyiMCpEo9keJU/gXfme+C
gZ3Ezw7mngjVKT4aq0VheRU0t6XuscEvc6wb5jh3y8POOBeu5i3ZoAEY0n2fhsfx
fs9o2ixS9zs5W7jeLeRF1sP4GBnnC4Tn0cVmwu1N/Aln//3LXYphIW4DjZUhliAb
nUY3zEdWPrW9OL0NrWhuKyltXhuXh1HWgB6roSIgt5zIYKaJCSeKXHqoMrE4ulLi
USTQ2c7du0RDZ7Pxv49Kd/5snXXQ/xElv7Z+Xx+XL9+RuVFjUBz+ujlij9Dpn2hP
1wWUWEpWN1QWKYKXdfHoUAiyK9gRPP5fdbX3ebfzOw7pHWLf5PESO+39n9fXv4jJ
VVvqg1Cmg6nUIsKey3w2EuWm1VPPF0peXvgVMPR3z2mztw8uDoxRLSZQFTKpsOr4
JnIQS3m9wQMCHOo32CptdtQltXQA+1wuHA17qaxRTMgViPymQqMBA2YhCG3aWb8A
OMrDc4OdLPIPZD0FpJAS5uS6VOnQ7sCy9e0Kld+5DzA+EmOoULZSMi5kPRC7fMna
wkJr0mjBVDPoKTUVcbOOmSInbVDJJ4egsrzQXx3Th2nMj/UOKhzommhX6vJG/qEO
Ukh71t4+hhglgtI3S+C851ZLOh4k+8utg+LzgpMnhzKTnGyxGc/dZWjht7tnC+ct
mr2FO/zKyMKQDddYY2ZtRyQdapUbTnTRy0E3uKekHaqLbuWAln05QgxUtCx58+No
rN2plVpIqh+/DfzmaY3VrCZwbjx+wa9jr6B2nLN0Fu3hPzbb7t70wuOaXkYthWO3
enC0z2PwDHBRT3Fdtc+VsS30e11smJ12j5aZHjCB32CJ9LI6d4BKNKU1AtsWi2zX
VUiloV2Q03a6Zt0ip+a3DJ5vF8HqgPDcm8C2Aq2wyz9OcpnenKRgScEF21vEuuXb
Bbqs1fyfVrf52kC7OXkSRAdInoOa5+ywYNLsnK0jMlXvkHgrx+PEykcc8R3peEeA
z0MF+FU00Qx5X12kJ+RdAEri3S4hyuoiNZSq5Gm7GCG+3rMzdLFqsFeWIYEo/qHu
GhngDmTnpbNJrtJynkgk5Lm2cfjBtRI7cBAgfAiNgx7W8mXYKbssauCxWBjL8+EI
1EQfll/yeKvPymh9iVzU2HzULNeiktiJQfG+0kQzfm3KFoQST7wU0iS8fwa9F4aJ
hiZkIZldEfpmG34xvnBJuieCiOxqyCAyEIiFhOCuMuLAf4BCYH1ZMYA8eImRb31K
YE2LizzOw+4kdvIDA52CBbI5IFxMf+RRayCmQQUzMITwDqNabUmycOtBz2WmccnV
8NGF25xnEsLmrDoQNvrs4xW0cyKaOiv7UJCo2zH1Ox1bpI689ZoFtrbpLqTZ62jQ
ic6t4SmdcY8Bl05EBjbWhgrw4vWMl/rihiPeB5LmXFm5RMSfbns+miPDhCieWm/j
5JHpsrO5LbQEoFmHTjeVaoZU12K3vF46kHg2qiFJsMbef2OhfYmo0s+VNpjZdBMX
taE4otzRbsaP2Sajk2kI/arCmx58CidSHSXM5/dSaWb6EQUlm7xHGYLqZeBPB/i2
NUaX/r5HFIg8Q9f68tQMbWkgwsZegd48h+hXg6QPs1IcXz9YBj9yziNFucStpqcB
euJI2jUilqx0vbopk1NhypLLfwUIBwWfcymzSbSqayshIRqgkRRtsmeq9PWtyWUP
24kXdcUoAfPuEbFRSK6n5ZUoZqxKqN52thc5iG6v7kLudIhoSfWouMMTlhe3h17s
UiUsbGlMMoMtAROqUc22C3jnZ4o5HijwJRnwixjKFB6NsNYLno/yy+kH49NmPNgn
9J3lemkxRVbYKEtvP9yOpQSG8tpWDO4Hwvj/jSrBzaPiER5Zghhcm/rtgcKvYJ4r
AEiZOLS8IOR7Yg3SNnBL14RuxYgrHpcEXaulkaXZcXJSzjl2XqkIrK1t1n1uQtY1
DtLrbMzMwAb1tr1gHC2JpszpOORJGcLINdeiv6BFj2fzpTT0KMEddIRSS5UUsio5
zzYtGmjGxUzt4LbC7oj7P9nqXZ/UdnwSEWNF31whFB7v0ii1wURDaO8pVIhLcc97
Fw+T3TcvYTeqhvxQ+Tjn2SPL5IfhehgABCV8p7RbqvGdYk3el1xAu5v6A2zulpm6
i3fDucyRipuVk7fpJnoIP4bbCQ/sDtI21CYPO/oWZrvkr+FthEqKqJDLpVV1P7S/
2hz3+I8IkbOZEmYs6FgqUDfI2tHwxayNuQG7UfxzBIkw+O7f+7Gbza80OZSleaCy
tQ3uDhAOnDjNhdL0G2S1+zJuQNpQDOQU9dZvYJR326+/hz79XVDqd1WEdib1mWO9
cbxhr+OumJIMfAY5TzV8DLnEfuwjEq4sYmPy0VjjdCaxK/UgiFUAFOlcAT+ODp7Y
CAkO9vqrrr9kr069ySDTNi/9w4HyRUyJld05j4EfAcSNgV7FN2P1zXfRv+ebXN17
qCRcOx/o5FNIUsKxwLkrsESEz8+n8kOauYmM2cjfwN3fu2MXMk1l6B8C60xH1c+k
g1lFxhj8OAU6gTuMtQyivSAXH26CrkE5azFXxAl/GXnf57y4I8OKJGoge43XDQSd
spfPwccMiJjfzxnh6afMNRRWTaFVP6lez+KtTajHegdR4DplR2M2UGaqytv/IACs
ajPE8fVCh1Y7jgBilNd1SeB8wOm0BG6pNziBvDu/39yJzNa45J7XCl+5W/aMD6fH
cAAolOXc9+mjWAhNl14seUmN8JyXkzaP5m8/PxLW6NQGE2/Kuia8yREL4P/HrmBq
5OSaZOtmPEUIx81AeCBSVNKxjmJ1Wd4UrAfqScUw3FM3I5ljBqhh1eDa3xzBwKYT
VHHTQVZEkXC43rdDKfm3nYIS+gYLyZSf4lXC2SrhmNDHgRTuxYnTVGYAbkb94lMr
TYKV7pDumdlkPu1lA0iqEB1NBFdfofhyo95fGx8DVfUHEdKiRGSFgvDci+PTBwO0
qMsBvaqoaMLzvmw+S+rxb9u4cQaCeIDGA83XLx+GVAaU3lPjV4uI6cE2WzSR/Y4I
faTziWJon74HOoeDteILh9WCjrjx2hs1JHkJ4XUqsdqhJKN1Vsrz4SOU/9G+juos
2RvjIzCNn3z2qou+CwDftRhUzw7WeJhOk2jwlwJBpfEtmWvBwr/U2v4+9ICRRONz
HYwK95Uz8jcYiLBclwR9JDYuN1sP2hoe9xJY9+r+fL4mwD6F6oKRvJo832oNQxRe
Hmf8i4VS46c8cQqmpRtCcUKa9nVO2HNhQMx08DUgweslLir4OVbItQeutZcxbJzD
QYvxJ7fgFJJEhB7yt2vcq1FDynIk5GsPqLKnSArdZXIfbjYGQoHV/1UOFwuwgxpp
ijNNdtTBm7B8LRuzayA8FcA6CxKCVHXxHK1ssH/bK4irzH5tFFwZPsfjWzQfIZuD
FMKR9XHKDBZSK6bLNELiV1AIwPcGCBLY6ZnMP8ZSL6DRyoPDxO86T7/KWmdEeUuo
aL9WxXWf4FbB/QuoiLll7b8Rg5eohW01PP7o26NzHBV54BRVIeW14Zc9POiauAIl
+iNYFp9FTWl0uTJkRMiYHMbwqIPiQET7yEk7v/JG0muNIzvtiazbP4CxOEUqAa/O
Dj/eA2/okajsHCAMHBR2vuabnOdEDhpTZ7XFLcPYD+Our0pTsEpBa2l0zESFB6/k
5LPMzHFi7LaSn3kYC0d+yMfBy28ckGqDnPtSPfbJVJXI5PyiQv1DoSOyl7a4iB2h
9Zj1GRCYZyB38KpD29vJ0m6q+ALrSJmLaFVolRiYVfQwDrSGtF1e+ajV9xOKCFZd
p57KrtTYoSrC/MueR2yHwok1EHccUrx1+wfDrAs1WySj7wBRyUiZKbK4ZF3KqmYt
oDY05ttsCAe9JODtAoX/7b5MSVPrERBZHaszJ1iV3ku7o8cFg+3N5ANdyiQshWYM
B6eYp57paB0avxIgr2251SlPhp+782wOH9pTdI+RgNkco9wFdSSZ4JuE9Rq1/nHD
vOUjhHIp90Ty4rGNxgLkJchIQMGApJ3YBa7na2wiU9qiYKkJMcpjFjBa6/hHEO0w
ont63JfWHfWuIzrgsRXcTFbOlSUdx8UEs52HWSQbct+DYdcndHjSYucx7Uf8nW0w
gIj4ii0Q5Ia3h5arrXtTuhPrjker1lepmBsujU+H13IbipW6bCHVkSudVdC30L5z
hP6Ue3UyFUO/p4irv4Q7XYxN0ahy+Xu9OA9K/norSDhOqg2NSTLn9ikoahUY4Dsl
x2GCFpjag6fFC1kTMEWdN/BHy5ot7IwxuVJONs/Tt5byYurGjHNteQ04dQpF9BGT
yzesyy5gJicowxoGnri4Xa+/0WS7HEyPJMWrb8Ha76ouP7wcazl50Q2ZJtDL/VH6
gEha8X3PpMcrfKXwxknlq/Dpd3WRYuLGHDizMjESMA+/qDYQxt7To34YBGgOAlGI
qsrcdvffoVoxfjSZljIor00mE4tuZFdCpr94LF2BCZivxKb+OnaJUXA/DatU+voy
Vk/la3QH3rdD6T0CPetouG1e1fTcpWpPaA2yXaNQQ28IwteCvgxoWJszmHQ2sgJj
QoszP74rttDVFJCcV0izJaWDhLvYPs88t+gH2Q0uZD+MEkOL8misZXQL5d5Vly58
FUslgS/9S/sTECf69onkjlut8/8gVLnKVOb6Qx1VJF/7uUq7bTxAr7s6h+HzP0BE
mq07ISQq+Qo8Dg3guPqbevlxK4ncl+AMYIIXNgOD7sGMZb4Y7Nx/K7K7wQnH8xAI
/TT3pv+T6Y01N3FgRjrsmPIMNGBrTnsJHOsCrZlPyI8IJEhsks1muJtTTJ5KFwTn
/zc35u8lR9DL6YsofeCG52aObATPx/Qsw2+ghGvGQBnF1mt0cSWQm/mifX3eH4wy
+mOOccIsYIv+JA34EAIKzx6WnjzpXak/NCgspsekoSpmShsCet+YZ2neRjA+SMHq
s5g0wGXNZhr+UwfG2UoTmTQPuiOggDVmA0dtfdUkOoMLk1dFLFr3wwR32yPvjpr5
EWwzNROSPQErBO0jpOqRQEjrQlX9zRUlH7ZsD1bxBP1mK2JtDPQa5raOlCZA9usL
SC046K27DwfHv+b8B/fN7m2v4QjrV8B0n58xQFkyhV5Epn4hXEoqxuVziM1ln/bl
a6MCQbZxTTaXIIwtBdarcAyxLdPz5JlGdCBwcyWHr/wvCQARn9BtIUTCJxqB/zxn
W8UpWr4rYMzNccjmTytkJtSrEhr37ZW2oucCI3BbFIG5V1dJqUq91JIXFyNMmYp2
fcNIhsVrzb3zMw8Cks9GTclRS44/bprlTCsLdK5kgW2/RhGb+Z07T0eM6P76uGKD
WQApErMvcGYvH7xLmWVIhsetHIclwBONquKnkbhsGJmPM52U5QWx09QgwmB0JkhA
ElV7vaGjPTOc9+5AO8VCxEaRpbG9acMEQEqm2q4XRT18zBduZCADCwDjA5bO9efu
TJMuYLpRIR7N7srBp6BhvYzMh+zyLMV3h4Eim2jGV04hxyuVBmk5wwF4k3hu0kHT
26lH/Xa8F34mjP5gUfKPVi4Qq2qEnWSLpDd3pKBWB0TdIR5DzCjMzb0QswvdBTPk
xCwFb585Cbs/cmdhm2Kdm8UwG9lASVtWZ98/Dbvi9uGCgZxDPjTi3t5wRWDn3zbp
CObjaesMAv4ThmF+lJeDK4KJagmE6+CV2kYQOryaf036srvLxfkeLBBoYcHO8suJ
ckQfRw2n5GLGCUNsbU+Dx917/EAjeWek89e4yZKTOZPcF+PefkvOtFwy9/aIs0AT
kCsZ1r8VvuHEi3begOYHV5pk0cUfVWNEUnUKzEwcxvIrUPN36oVzc1UwqzYumI3i
IzZKJCJ5HKdy/BJ/vqf1vyhLiaIfxIABY6TGkSoj5NaTpuCYw3kUg0XOciQTYMMY
okwff3kkmye7Gr12STVxqSosqoVtiqosSqPUihEfkwjUxmMW7W0CIWWLPMbTg24F
2nGw/RAESwrq3AqoOg3WXXB5M5JhiF99t8iuTioybv+6LsrePqRuCC5GyJr+aqt8
DLWzOMCTAa7h7H7r6PAK3KxRvdyR7G2PlGCup7chrZZDOQ6OD9KSUwLCt5LSa8Lb
IUQkELATOEL7HX5Ndqunnxd05U9gGWOpP+eKe0bH/A1kfYTDdnJ6MUwyxo3nBx75
XrS6d9RIwpG3UdpgT4CfWizdK7bJvxlueR//vViTp+if4wtKP8uECo24+VC1R62Z
M4HAEemrHvNU9VuKDugOo6knebUNwiSaN08LWMGlQ0847/IKfP6WWNlDG3g0fI/m
TqQujSvCLAyVDVXVhh40L6uIcBNzLOxycq7p5akTHGiTV0K7Ndb1XrLNvKRAaawA
od97OPqPAtn4SCfpMSG9ghPg4AO3x4zuTodzYrOYK/CyoU9o9cc9WlljQAshMw6G
osKx7Nyn9i/79ht5ePx+KQqVYOwDijvl0pVmLEhnEQFk4INYjWwyMV+m5LErrvDm
lAW/Co+IVwDKkBw4HisqdiaZqFZyrtlTe5Pjf7gtzW7hebcSekTlsjUH70P/th38
8f/NbRxwsqqeE2uMo4YFU23TZx3cJf1pmDYPCDuEnOOmAZSJt7+Osmf/BET0u87L
/5YtSjAg17wvQclBCsmCI/MGTZb7Jjt81s/Ba/UPVvvsm3jTtItfNoHW6SG4vvLT
VBT9iY07ga/4/FdZHrcL74eSE7Na7XaXD8ixBxmMt0jO1lGJpVXm2TdVay4FZnme
Y4ktXHSxA8mnlGW8Q9XIX7s2GZtgj/I3Nov1PhuL8uODk6xpakSA1ZNCHalRSJTo
aSS1CEeEz2OiVtnEC1fD7z0qIr5+sgfwk/1e8MMb7wV/RPaDLU4h37dCYELxlXvs
FSXbMD8qvRjxZbxvGOLsDr8kBK5ltM7y/JheUngWNVnHu/xzpaDyhjHqZlEnBuOs
YwpqRxn03x8sXtqnnKWgkNDIYb3C5caPyjZnRZNBQvefJCyOrXUoBCBEPVpZMxO2
h4nfF/ECAP4qfmZ4TnkOH0kJN/sb6YxpkA6Z13wxqE7xAyN1HgoxAdq9t0mJdssy
xtX0ermDHRQ19tYAOjde9MKKYbyLg01viPMQgs7BQnvDndWMa+scrEudcrvqptr5
2WE3/53EWC/Gl9LixkQfS8TYp6V5HC0qV+bQitM+fSzofC8fCqBCJ0pX/GgRRll6
0RN+mOozsg4HCDFh2oyH/yeRV/K1KfK0Tj+SO7EMDmBz9zLl7AwFmNE8g+6kFhn4
+IiXnqor2c1HDeh/to83kh4o94j+xpB6zntoPAlhZz/MY16s/0W38VOzrlRaOaAC
PyVkGozoKj5ULpZeKZPN8z0oPo6CqZYwm2O+rPBzEYhso6MWvZGQgwW2WuGWbGPW
byMQWqgkRW1dXPiUk2JTo+WOvuL2lu83Zo9vQa1JLHmgg2ar/qEkGLre/rJjh4Pz
LjZtj1xNxylEC52dqpkFmzRtszx0C6FNuY8rWPGenCLBQudLPV1PPRoEPZA9ClP5
OA1EdrSE2t9XjZelHUssX2wnhJWHl+8p5RSUKEEOHQAEiUUMfNG2hYE5BL8m58t6
NHyaUu4O6vtFbMmnq9VYJlqkd97j+hD06LuMrEF4u+fATiclO5UP7ko/jgGd8e8J
HPX4XnBzyyrhd3LYl4jzAeuSawFQovAPqtk/bP/TglIuiqInJiXHRc6NmTYbTr1i
J1QcHa88Wy/yflPG46gj5UBARULzsl2wZLHSfPZg8IgrBF2Y7jDi6S0+jz1BnQWK
H6wglxBEN570t2LviTHDytk2yoBIbXZeGwq4tcOUAd0sJHlp0v12kCfAYB2/Bl9a
KCGGvtXyEaiB4eUSgAEPcvjWgGbAIQl1zQvUpxACDroud+dlhBEj421XNd7V08ZX
xerw2l9+jp2W2Ot1zP4C4KBDGtyoZs2pyzbwBrte1Wc04o7lSAkYH5Fc0gkIdgsc
XFBjOgp/QyqM/9nKOTUYHMb1NvZETJZIAPRZN3kTar0vifYpGPtyNeniw0GWCJgF
JfUJjtmwIVTriss8IXZT0haajujTGJ77BRsi+VbVgEhvl3qQeXw1ypBIk57+a6Aa
OVJb9Q2MYq3bmJyY7AhmfbnTF/L+pXe2nOG2kB994zkTo4T2quc2luc2tW3AKpjw
60p0mNlmkmv6RqrldIAs8Ldb5Kh3OdDRCjWcQFknLOYFKgNmKTEhUMn5HxoHeFcE
FfD8RVYvUWb/R4kJeynDPQwyU2EfaluiNz/eTHTrxVGzpkphQfwbx5a0T+ijqxTU
V1PhTKxD+azyIlX9AivcCMWV/MHkdD4m9+rpy/FusdSOwu3Keh0Sr+U2VlQUFcoF
u1hcHl8FoE6HKb1K6I+9FLgDrzdSpyAp+5h99VX4wDWmdzFa33ESxyJPxpUABH17
nwmNHLQtp9J0Y2ddAI/LLQFeIAZvw4H6EZdj397xE22aSCOu9GQjvI29DLogaTsx
ZuYXWT8aXDyijFa5TUKySJwwieuLJtL0ah24GB0UhkxV+wepTVk4Fw089B5edwv3
nz2JBAP0305wiyAmmojB9RjUYY+lndC46cqEY3z4BAIjX56NGLvXcDlN59VyHn3F
x3lc2T0zDz4K7wtzJbDAS8DaJF26Egi7I906EPh/ivnCQceDT80nFpI/e97b4mYp
QBgwCsqdSo1vv2em3AzAsZqxnELpRawOYcQ1foq2wGHJ4svMqTahp4UQfdFx1O9k
IeF371rZ7uVJSGyL7/yNttMLsFXHV6UxA+HzQ8X9U43kl6GksDrj9MO7ZwdVZI62
GWqwIaavWGToDhOH9m2Aw+Uwizfj1zp8WqjT8BMGuWsapc0w/9YL7oG4jRY+OI4J
DstvrlUw0CNJW3/sHgvVNZmWIMyMB5aFsrbE7FR/CVLQy1S2J+xldf8B64gnEMFl
X1xSoXTtDa3sgLwrw03sHGuIjqjVi3X7WWuxnZZilgeg99fMDDyislXFQxSjKNZV
/FaDu28ei4dZYWcFGmcN134fLIiYTqijGsdMTpKk7uepaAicZKVgtMUaatjv8rC4
XvJUH1G03S1+LVH/FQoZKyPRnr5tEumeDThjL3K+XWzFbvMqP1Drgx9GtIb7q/rV
4W4XWH9DYUYosJBQnia8iphUCc/TxJwtCJLKOzNiPtH+HLNk88Fgj2gmqq2qQJpO
Fip1Ira6o3ATSvFwBx2v+AVZZYAU/ijfdw/SifXZshIrDGpIZdfcTNf8aKex78Y+
3QNeUZ162fcvK5NynyEKopX5gGXlEZS4AfMaGLjgEVrc5CGxut7mQOaPV06/eAN0
6VnqCIWGcCMZK17rUHOUOfflEDj3mxRZSmJZtuUuC+d2faslViwGtWhvOVSCxV3n
ZKAMDhpdWup6aaAZVgXQED857zrkl8Fi+Vvt81/ubiihyFkEXdjdWwN57xHapLU1
UFyCQ0XDu6JD+dvxcjk7reZdGesP6uM6AVkvIGaO9M/XJpyMxqcdgY4cwIrp2ab4
yDkRjjcKZ40nLF7rvmKy/NH9Od8+6SVmBCibqIUnTRL7v1t2vkG2c4O+c3YVKc3Y
5mPWg9hhQuGJ2RI24P4JD5npSnmzez0UbrLiI/D9KdQqkr4v3rSVIsBoll8LNQyY
U29EoF+S+foZfyDhmVevMAk6H/b0o62o+InQsYk+76W33+6dk6mg+o1tryAh6lQK
B8Rv1PMRpUCZ6ryLl9SXNDOYCKWQrdAW3yF2egvJkabadLycL/YIgx81vb9clMYm
lwv5PrSsUCsur9l5AeNWMT26sobHoRBamnXJT04NkJp4r9EnfsJNzSmdwdvieHeb
8WWsL6W2PDVaMbjniIQcV1lhnc/JfSKsIgPF8hZqjlqB1poRaxMEebBXOeB/vFxR
LBhQr3Xy5/ZPKwfLNYHkHBXiDezduk49xFlPH9J4Zdpw7TE1PkUYyDmIiOMgBJVQ
H9m+FDbraHs3XCt70J0LkOJuQpT83z9BJ8MsWmkW9YR3/anE6UJlSmOxHhNpl4gT
zIHml8yiYarNXWOqzdbBbs052vMpSr/JcpMoU+7JA/DfjYnfiGKbN0ZMj5TPTXvu
5aS+fTybGMYul1HUqug0BG2JNDaqBKx2W3aCPhNLA3TiLUyJ4wVcOADrHIwX4Ql0
pUBROXIYrW9UeEDeIX9Mwy/dryuHklT755tBrcNJgbZdVMvXeITZOL/fV86WHd5w
E6wvywsSW+CVYZRl2RvJcPt0KfpMd9VZlxOXtkKWqoUkJ4mlawWv16xYYfORpTOx
1jB4ZnU7RQ8vGCIOirBNpjsebaLmt8SBSRj+ohTqlYHEgmYStjDwB0juMlhz7rPM
1K8kT81vZc915Cwlk/XBGuX4AYm2qzsIqyjIBHoSJkjdDyMWq17Jr8++gCIUOoZ6
ugurC5kPmO25HMqzjAMYOKB0Kz+3aoD7BQ7xYEvo7Kv227fSpVlZCYKLcJpvPC9t
A9wNLex4w/InwxlnzxkVVF+F2ZbScfPu/UaofQhCNe+L56d6Hz44F0Fl6Xbe4L++
R83Rv6vUnQ38hsmFQqL9MoJRrpHmw+i5GvbmWuvzmqEMB69/6gNYGGdAPrIc+Vet
Q9bxAoGmzsyZzW+ypcIeiB3ewQFt9BqFLasb3kt1xOhTBPAc6nf4bUwGjkMxOmqb
DRqwbFzr5qx/eXsyp8n6rxCcmyDdr0+UhmBO0k5076ZTTCTWmZlpetHngh2CVkTz
vfvHJ6pn40t97/IPGVdgquPMWPwc2Ydl/hpxDL8pdmkHYqHMGNf+BHqtuj2Nr4Ta
tlKlNYP16cYtP11xdTNC+B1UcRSKFuOeaMZGk0L+JiPsaBVG546CNtDmP1Q9Ie6R
BCj0ytvGDT6esDK0FbHjmt6OrwRAo6uckq08/GTyNlZ4KwiQjGe7nTNqt0BeTF2S
87xLv9Tl+CT6TFLjCtSC1jMrD2E0Ca2Qyj0ZWEaV6IM1Or+hGcbyY6QrBTQhJNFr
vOT4eFWppQc9oJCaQ4N47o3z7OCHVazfLbhSQGz2RcrMdzFTqFFLNFMNsf30afPR
52QScelxiPr7o59ekzOEIthc0FcCfuf2TOUQfxqYQgp+9wWo52Hi30Bz5dNMzxFg
hFhTCauYXn6hi7DKNNvYGCVys8FjwInqNPmDProxYOFGGdHxlhM2k8zMjOUPexB1
mmTQDuCz4ejkKdSf8u6g/xsZIIYGcN2uf9sXNPD3jQtA3kpCJrckXDprtLrg8EB/
a9f8mkOXRx+ZOR+zDEodnQawGuGuSncHHL9mTkLN7Z62HYaZAv2kO2yW+ievELqF
eul6xr9fCPs2rJYS/D7pO7NNPJNnQK/MH5AnrhOLYOjGPXnRe7tMsJ5rsiTTkzSr
GpPJaTeAov6Jiv9fVLwg4sXw0Q84hTom383nuwKnXDiqi+a5pYceVRuGB8AdrwTn
crSXwSdt22fGwQnr1qiCZDATk/AuMJ/C/NGOPEHiOG/0JS3+E9WFmttq2sBCnN+w
5ipz8eM3VWlBF2h4U4L8g+df4UJs+upMjkYMmG9Jk5e3rkEJXdDy2/AGVr1zj8wB
04kas61/LKP+5j323a62jSvJh2HSMHHsO7K6aZh4RSCtjd4JH5D0Gmq6sMN+iCeV
b4NxKFNru/D6wDXfGN3K7wnBrhpOKVtzHw62TzhOV7DWxU5EWQsq2bk25/rdc/Zw
PiZ0N/MV6nxZ2HB3bDDZcgPGdYv2P/66jGHH2lSuLhci8Lv71wN7wPxP/mJbn5iG
PrskqDxYMt0quxwPmNpvZtiDmAWr4Q/X44wAXt0YYe0LVwMD7AuOR6lY75VW50ey
qkr75aXNzKVD2cItxC55F76vawuYjUbizyWX+lTuvsI5F1S6OAcnXrb//XZbcQri
b96KBgCB1FQqvKbs1TzRwpJIoS1PKUbW+SDNYYWzwZXUvUEBpul3FrtCoORS2y/U
vl/7WuX30A5rUbVxeEjsQfCStBJ8EHmRWLBybvlB5Hx/2wfQNAn69mFsZE5wqmIY
Vv2Vvjvnm0Uryhp0QxctJ6WmlWF8dzq4yK7Bvq2uF4ZNui4CM/H4r/ZDIH3eakaG
TnwpZhjjJ2nOzB6K4jiDEraf67Q+ge4lvw2LZ3MKlXgvoXGs35Y5DB5b8r8ay3fb
wV77RD8rf3z77AFXRZyW/fMZ2fx2GGw9YabaDnTRLsuFGpPatrc78NLbi1dvncqd
nf1Zpt5PlneJBMCHfJkQGATiVtfd/Li3qdhExaGwv1LKKmE5osz2bcp/KvXVQcnD
aCDyFV7vFerGSDkTltjOkjSFEzeXqTFJGdMF+N/mQiQ+EiH+icMmKoocstf7IYEv
YjZc+HFS4aMaVb2uJp/JT0CixxybmuCT9/rZD6xoCyLvnQ5MNqSfZhHnpNMwIXcN
tV6QG0+jQG5Q7F2pv/pq8xWu9m8RdRwwQHJMshcRXo8GrZ7j3CFVi7Npqze5ezoe
+/ZbmN5TW8i2M6vWG6nTQV8rC0csyoDZQAfyujdkiyuamVt7/Iiyp/s0DTCJIgaO
JyNWeLbrf/KyCRvM4VsfN8trN6LRCL7LEaCADixPA+PHmDsEdK18zfeRxo9EGB2J
TJWW74zLk8YTd8LUI7BsdpXFXrze9eQvGoYWuYfkK3qxe9EDtESSExYk87VZvFAU
eMm/U3+L6xPVkOy/eKrXs0WHjuVMXoWGsCnA5kqddcEga0EfbFzAOnb7uHrqUcgA
FZ5StzA1OgFe/GxEkKgQpJCt1EfS/GxEJRJcup0SHOrd+uMMzfGXre/g+urYOSHS
3IFdFRr5s0WJdapUQBrGPb/dCBvDdynCO8VNjPs8x6C8vHpAnaar0KEVQIAigB1Q
xrNXNWqp/NkN8t0XpVnrRYNPKm/KzXyOenunmjIpYkd5e2sUR/Uz94Iey23iGkz1
mhwo16jpnk5PMDyicO8ynXKTILdQW1ATQ3LjMd4eEQbYgJhBAn1s8BvJhleAsZGk
sEOdRQGPwSWl+ZpnetQq4AbEUsavOy4IhC+UrcbRk+lW47+KzXpP5IidxvXsDpYf
EFr7uCkSNJt7IdYrIrYVyFPVygTSpJ20ODmMjKzmgZit1UcCgAEsZ+vT765cdhEt
NjG5uZZbwD3HDbk8oljiVQrq2dcN6xj0ctd/gQtfO9nPqVxx1LYmuQPCrWhjqAZA
3fx4RAwvzuHnwUQvs+wIe4Kcb1rB5FcF80G3Au54pGFCZ8sx8DurEOfLKFxYFtQJ
Wr1ahF0H9JTgKr0iceSm2ujKMCKLOZX2LQXG3Q2wPM7o+PtfMEo3F6l1/3nSAy4X
XeVB2YbTof49xpS4j+9O2BAmesARx0DrZsWTVGCG1uGoXx8obhkfio/i96UYL0Is
szTF1VdQ8MK7MRUwd0UWF7dCMYM9rolXZY5KA9lPb7HZiF04NNNsyKVlkHmE43+C
euMpYQR7srLEimmzi0MTX1cRnRgBHEJ4yNQXim1nyvVy6ZVxa905t54MGnSMCzIY
nifwiFa3pSbM2iIgAl87klXpebWMj5Djy7sgBW9fr58JJv8xJ0ueQnfrnN5qZkUE
T+bnWJOdAD4A14rDSodWLcGvYmJM/bZHlj2NsWi0iHLv04UGkAC4JuWzEFIt/G15
7PHgyK37NBfotskpne/2NikMT7wveFrcAiu7DdZn1chZ6v2cd8L58nVkC3goKsbI
mGv40aTQu5Ne8Hg55o8UXnYh2ambtmbcZO54nEYMz83vm2TsF8urMi3pSTWKDQVm
eUDFgqOoj6CMvD/ot/s5/G5/Dp//GB3GLecXHcOB9rMs5NjuJcZG8tTAYyEKFAUc
npfOiHrzHoTBJAeWLXFjPEG562D1noo+Ed+SzFfq2qlU2aqou5pf2/mZj2t39Gpt
FidXX3fXFgk7SX1k6tRVFEOdUUUq3gFfMdMtONBiIq3KTG1gdolsrezf4CrjmdpI
EjBdQ/ofM0R8F7+xlnozKPyLgsOQ1dqkUGJSEkNtVfxyJlmccSsSBdf/hFbe34oZ
R3GfdRgwJzwvqVyi0raRDrBm9wjnUD4o68uz7WhJz/L63rZQLxOYSB6J/tvNN5nb
u3napInT0+noB/54WH277W+AZ0JegEqi1Je0oFhdVCaXNdxl/qlU7FDpslqfOSEe
ozd18M1Yjix8ur4hPZY1kqg2jqWuRVflE1ADQz5jrSsK1p3IepmIsIv9DljtZ398
xv8SSwww/FAIwsagGXBEIthjLOOj+U+IjI3UrwNYBUbxTMJ0ArIQyICeGy6AKCch
EXQiymTExCgtUSxroYRqyVTT0xBYWnrOAmrDprOxLims7vwj7mbOuAsqAWgNJMil
uxKq12dm6jqfKYZER/G1P5GU/MvXLeuhLwE5m0+elumUiZ0MCB37YkX602hCNpay
NaCfIyCk1JsuaIX523UvIrS4mnQndO/fCtI1mcGIA9yq11szvdla2XYHHrmJsf3b
AIJtjrgv4eKz4PHOunEVGB4q4v06SuD2tZ5bBf9KhC7CeSpL+F+lD9BFUG9cUyUL
Jo6eHxcG3vC5SeIfcFuFVskrdbyvnbNVzcDwFwGvSMYhFNtsp2qKVeLY7UU4e7lw
+jQLdzi8Ksj6P86oR79Dx+6+hhRalXelyio0TMu7alsougRoxN9AnKF9BoTc7lxJ
1o2vEXXORXMDuOHrjoENi9buqyDGUy7k1gZ0GFh6BlW3/AAD1py85MaezDxbG5y4
shVXikIvBxboGxwymso6hrneg8VRjvMbHLDy3cQoHUkZ/aXDI9E5yk/3n0kBoXPZ
A8nJ/hQXYq2YC9dlW144nfr5y4V+WahyKwX4T5NI5jta6UmDomh4+xCQRWkfALDF
KsPvSHTX9komiN6vfuY8ZwakS3gtaAVy3yEglPqfKRdDfirHvQTV3LuXtxoDuMgF
pHwjGCV5W32kfePOuoFeefKRfGE4FNGpOqcOKmlyYas3U7Jdk6RWaUv7gV4Lahx/
7zZqqj1S3h6ZOlgvKUlqYMyo9fxYUm5DKY56FJMN3xiV1QFsUg2rp3c7C/OBPkNa
SlJqEM+LKQiRS+I82rgrzzR+c6sX4tiPZcv6Emv0Mxbgs+K2p1Z0vqNLdYft8He9
d/UutOEaaFOyWd1wiMmTJ9fh2Kpue/RrbYIlnzFmu8dys6fx8weYRieYcsdbbpia
RryRI43DluyJZGwr1L3eK1JpnkplKJOrFrMY/yH6QAzOnSjKvVEJsa0xJGcCPB+d
BukSuFGiuffM0a5D9WeiW5sspdJVhTmeENz+IlvUlNX4tVAJBrVaQe82WbtnQTP5
KuPxiSQ9cgAMc64oVkQCC0hBzMSj9bmIikmejMRMI1ya094xm3T0fd+eyLEbgaqv
IQ+kDocXZmUhI7FMfLPffMUww4/xS1R9bMPIH33cqiw9B5a4W+DUGeIsZgaaBRG9
27Dxg22LfMmHuferEhw8Xu45rD+3N/JT29juhEgonOs3jfkMJ7LU3FIDZGjxt+0x
aalj3poEVpiIZ05juZl/jOkPhyhCIZfTpZw1SReSEzPPLYp9RDdZXRplye/hJk8S
vlPmtbO5NU1El5JQvSKpOfhOX+l8BInZ76IINCNKYGcGL0XN/Ijodhp61KeRaDvr
RtUBDocTRbXEV4fL7fpqPkTMsfpThhhGKw7peEHiqAcI9NfGur2dAjEhtKuq0Yce
x+dDUCZihff3OgHd6HGoJjzLdI9Pp+5RmjNk2LS3CCPwDtOPrMk646mfCaTPUE68
MCdFyulEfeFfItTft3PbvSiw9Z/ToqowhHdRfzry18pWrX4hzoxw0iJAU0fZSBwB
xYvVXPfe/YoyyS2b4x0kJzNzNrebrnPJzNFDoJEFaQGQDdnLr9csaw3Fvow6tLRn
40qdvLCXmaFe5gDnHAqBHIIQGwal1D9bfgBiyt9ApFUudQNQynL8y92n0gaAGL2O
OGPF/4907MTcMgq/jA7/iN8b78khvgpPpJG2aYaH3Aui2kzt6xLsH2gemGDvmTtL
vT+8ry11tMKcC++vPEjUqIHGy9Vn/5H+uz7VCXxl12gihI0uJR96p3hA3OAqS0wf
Ec9c/OM8RpgKyEnNzqs/JwfGKui6wLZyAjp82IAdoe5JDfTLDLl00xBCQ90oGtyL
aTvOkWZ+cSVdtOFzMk7Dbtg1q4k2IrvCyTy/92aD6xVqK42OKirfpxpJ82lnCfOx
K89lyKGTVpCljbhssRcdoIdcqskKspsjs6Zp5fPn9Fj/yOQp10gOHNy7opUnP3ZV
8CNXz/u+19zYEC79VHgmlLtc3Z9ayxG/cN3A0igfwwpWGmhtAYkL+SSJEiSH6Pfj
nQLyaFwZItFGxdGYQzp92o5faG6kB42Poe4wgtvJRNAFG0IyMJUfTPTOYyp/77r6
PJJBqa7z3r5gMuc2JD3MoOqThh+LcMYLW7Wc7E20t6oKHdpJsW0tquHywYjbw7J/
EbhbZh3qIpHo+ptMkDJMVcGlQ9AE75tPpaj06Jc2I1XaHNy6OnOnNroKQkPf/t8P
/enlIPobyftUXjF+xP2uiCmyrzllfAoYJeLkY2brY751hZW1WvWwGiqGLpzFI9Xa
QLCEkIgH7bxATLCw7K2OJWpp90xtF36/5x8IQsOnziu3OYXVAtulEvaT8Wq0k7vE
N1cUR5chQZDEwx5j2qMwOF+XxyRRwZ9XExPcOjI5PbUgWgIy880rvws2CuA4oURb
0N7yJmePHNg09DotfcB4/mMC5iU37i128WDl64iWAuqdHptk9Un2q6ql4n1IFdtm
Qs8arqA0gvc0yySfHjuXdJdZgDpdCtkdMhB/JtEYOFN0SobI08hVDjYMo4zMVOxR
B5P8W67n7+m3bWwGL8xxO65yWVL4mVIc619/kzpJWGMFd6m/riRerSaC/BmYGdZQ
oICfoPB+1kB2YQAq/BPbqRKdcQWLcXsVNGTVTteFTi7N+FA7Ap48epewzzHgFth4
gwhSpg6S+c4R+l6nfIj1T7WyXtl1SEUzd51S52TFul2bAbb402e6eub05GfDbQS8
p5K0wbYH8CGMqmLfmZp1a/GW0l5AiGZPMcf014yCL3BwuzlmDTVhaTZqZoL56zDX
8Z5J2Xj1RzjvYeYDQpAyrS8zZkeYNebUTsZMfM/2LJ8nHz+j4msBEwGdiB1aln44
hC+f87WrrxmqabHD9CDsZlXazviZIRopWuLMn5IjFaRRKSdKLQYmxZ7HaJDnCWtu
d6QHBbxR9HmtVNc0lb376AclwmS89yhZ52Ij/TLaoeEvu4UHybAtJqkNrcErQDNR
iahk1u3xd7ukvGzXSNNmjzRnpwhYQz0/BDxfVCyK66KkrgOuYwWBVYBJR5KQVdjg
sQJp35OdlivljPG+otsxQhBC6R534sF1hXF8/ZSAPJILkHnDN5Glo7obH+GNQHso
EsajUS64JVEgeBRBvtgGYywqZ0nrasMxW19BNMCjDA5lodjV7UoX7Ae8AhaAkErW
e8IzDeq+8J5yzVbxuSQ/HTQWNGxxirHAvxiyavIeArkW9JllfzuPtppz708g0MYD
G7VhePCajU4VVFq6BFyLL99iXan/jMLE4emfosaGJDZS7UKeqK0RnmCOdqPEk2MQ
W2E8QXyUD2vFmH02axOeQ40CArSPvBwxi5u8D1vsAymMQwVV1YJfyYEUdYfaVqwP
8+L5Q2xigxD8/n/4+XaNZbDjjIzQtLdZAU5PM/l3mWSk7gfrJthIqviUdwmNByYr
+rN5ZNsVU9Qoe0LojlBub1wSu+yupaOr3QjnW5XBCGccBqtJuKwMqJ4XzNMPXkYn
zw8nw7dbsZAFboIC+27FeCBPbru5RSmhlyI7uPVhsAiKg+ifU/xjsiIS9gSGINiy
9ZJ/Myw3hUzM5H4d6wxWM7zkpzMrCc9NqzMCEi74leu3bhqs7AlqTj2zoy2rvfsr
JYXBaWAleobSnyzwud4+l3fdaTyOp/rA+eWLzaDHGPX3iKEtt2sL9/eK3mYpY+8D
FkeIIJEPacmltJYSDAYOyJFh+a1gW77i1JRMWkp5Lnx3aW+l3WyGqJRz+68IDZ8Y
jbemBoJRbmaZ/BX/De0YM0l+KcHCdFkWzFztdFobG4Se7q9bwA59hWCWe0FaMw2F
wEkDSRGosDbL/WyKaHsRN9CaqMsjo3XowE/iBNE6PlQyStrB22sYfMAf6xdWYUeG
5Dyj5alza24IirxGbozcyyyGbTfQzuOxYkhZ7TN9n+QsnsrGSjOL7wz2HDgIC/lB
OY7KWINo2UHdo8AdpOlLGEXZ1x0HWbPdqgTB7RxH1E4lmPdZ3wzAV5PNLdu1y6X9
pTVsxHWC6HaqzjntJKmDXIbS9xAm4F3mHjTEKqp5e7mcttKU72UQ8eTQyLCJ9Jw/
VJXfmVVPZsT7KHTnkRgdJY7ureNoQj88EM57RME3Zcz/DSWWwivW4pj6bjNxBTZM
P+kxLEe0yjge6BKvqCEiArmZeL055QEcK2MHK9OATl1sShEr9Xan6a9+ZgJEH1ts
j96vNgSNg1TFixDDP8LXGrjG9lzkL+x4kEbgoWkeutKACL54JU+ey8M01OAxpwQa
X0XVSgH0dxKpmSvekTWPFmu+DfnjtPxwRFhHm+scSYdCbnJzS7XBfgO70ievb3Ye
+i/qLOqZksHeu89mpfLen+5LqzofJ3tgvWdkootkSKuqEMTB2NLFHrOIMdTClgYG
/ePF0wS5bTXG63KIl1UpH/aq/nDGOt886Ci3xrsMM1kn526E3/fwXkmfGFn9yYZR
7UNmmRUXHEv4fZaUw+vTt7VYaR5EKTPPj5HIvPnU/aX+7DJzwlawIJsxVqPQM6Md
w3Gn+acp14fdSqzHw6IBqOISsEgLWEo4074Dme7YwXoI71m4Q3u+NLA76EkgxUwY
UPGFv1ypLJFv7SD8OSyJw5tlAdoQnJxUkhswUQGbH29Tq2bZ754pGl1mfpjSp+fP
gO6cXJ+xwcaWvM/w76BEAR3umJb+dICo4QZ6Wi2YavOitoMtshnKhaebMNeu6Hez
3Re9LpbgdJJlpozb6VV8b9plevcih1jsqKdhOPwDjm8LQi3F+ybWLTxegBGULAXg
uczCGfj3yVZBlMIGpuCoRNP8ZEjEB4Ob7zy1f9uSkUB5uDu5mKISUG6amZ/Qr4Hx
LIbup+t687wuW+l5YOnokSNCARkiSZvARDNhaIILQXyO8wZrUoRdtgZ4yyc9rP01
WkrB4qpoIX77u3h2GLK/Z/02cC2kCyDlHBqjsRdH8QnvvTk9LJ4kBPOG0xBwfQqT
HhTyt9nJ75Z/a3p0L+TyWCZ0nuRyHxJs9c0rwK6EMnnaFZWIZuCtIUmoQVmJMZsq
hoRmkTYXfI3fXjWCHotVykeD4DYGKnN+eCndAxudqoUCyaevYRNDk+UgifS4mdLt
9IMaWrEl/UydQjypJfTYril1Cl5zf7/MoQrPmfK9/MbypFEdHclQg60MJYTZy3Vj
rsW5Icl7IGZTBiN1FlMTjbuiPwlDoEIbBvMUepoZRGAs2oezxeA3d5/O6t+5H2ne
SU3IdGPXPv3MW3pbuuc78sx3ayRbV2ejQASkWEqQEsNLcHv69snAMvrUI1XtwZkq
scnBRFE5PZhO/jPJxpx+sAA3KQEGo1KelZjSGoo6TBSGJwJof43yQakPEAtYuhEV
6BnivXEm2mRo8QDTbWoVlUcnZ+Qm/2ibguv2nTbiu47uxXx8pwtK4CmgD8WSCBBu
kGNSdvEJP/Y3wtFngzadw47s8//wOb0RurLRkDChYTCk4HPK0gtZz97z1tWSM8hg
jNIKoxPdxBy6MOZ409ajFCmkZ1QJqZYejfhGXnuMmNGddnRPh9m5uB8h0xiKuVvA
mk7cUS9l2Kxo8IhA896uuPxwiax9BlWNL3Qu4rWMIoxEkKC5aFfpicUcaHrnx4mH
nKol29BuphawqPzziuR2zIYNwjiTpzo7maG4CjNkq6fgnyxl2EPM8nCJX0lgwSjw
HQ4FYKVWytJx+3OwAof+gP6EhouO3YhkpQ4d0ULI+Q24kg+W2KA1V5vemBWysJ+B
nKsrTg3wwErA5B3dyiXXTJZqeu7cppqggYtkpIYyQdlFNDBPMzrinHkXGDrvb5Uj
snBesougLn3RuQVQ5EQy9QfVJBTuyu1znEHTY3fIZWq2Vox87CwXFfw7fslRnQdK
SeS4c1e18BE/0/JfTAV3fPRl3W5/37e7rOwWnrx2vVXTFuMJWyi35P+lpfYcux9E
NXmQCYEydVVfMOg+XdRh22Jr5Nqd8w88dBvsMz8FK12nWRrvKbmCfwFtbKlnGr78
ntNO/j5nuodJJwe1VTDpPYsNhf+9xtAgPz9AcWg1EJs7N+pqwY+bxzfDdWw7AaSr
+eYVR2vF2r/xiADlKn4NnkBYPL0OS0QyIPKSlmnBMknlJBdpRK2XDfbGr/G3+RIq
As76NAZHf+WF2Ip1w7vx0094X3QsEZYsAEWG6mMx+9FnFcMZ7i3blu2eHCRZc3Na
WlnM3TPs1sZJSvUCWViMFoZPGmauwMOkFRcIo9JyyR98tW13jK3FFEaDgTJk+Kb4
chS0lAalJLS4T8j855NCj8nIflB5/c+PhUUGV2tESxeYJBoLj17KTHdaEGaLTeOI
5Heky7vqXQ5+tA8u2FzGqrei1mBwCiHnb2l9tKne2AHJMc2mt2gTeZPjlmuYUvp8
zGMpFCe6rs9FWGqHOGAKRDQ76uRR8EPPT34xswZMmc6UnhRL4YOLCzhawHF5SJEN
iF3dvhsptpyDd9eYr87PbSaIciCZhaQRf7Vs5ksm0t4g66bbhW1Jku4NPCjsTXcS
wgDtYbkNVQyvvWJ6eq726mIjyaelcwSWylDniknqMNwJtf2RjMmAc/DWL+D7bMfo
wPJOwfuXuXYNEw1ytE+1EVa3DWq0jXaNaWx673vnAadAGWw8bRJOJP37jWeztkZY
mt+WaH9CKdCb5sYzThWA4n8+My9tEvG6iz7crN0DZEdMraPCtqp7VSIclpofpb5w
JbPQrrLzldxShUb3Xz4aI0xrakorcWb7iRtWZ4r7K5MDdsgLaFp7KCLE5INOxbzD
kK7f9MvTqHngdEDeFkTU/yoCt8LoLOzfEJzrM49dwBfCHHz2mYq8HpYryIw7gmp0
VZL6BVXzXyq0oy1OJU9FFfFi9105cfZ4Z/DHygeJtSFuAaGd1AXymezDIMdNOppa
ZEDSKEY73SKD+tgS2kk8OFiG9h/0UDAdFFR/DKF5R1HwBYvpf0zbilBRTb+kv15p
7/8GWYnv5uRuKwGtQeHYilRdr/Eobp8ZEjspCQs1L1xbCuq9ODtmx7AgbGzvPA6a
SEYt2fBk3BbQnFQEM6JRJP0u5bRISW3cRqP8u0oY4U+mchQi2SSDRV1MjP8Gezbw
NvdjGwnuEXCPe+4T0vCjsOnZYVRMq5XQy9dOMvCS+QlwIpjF0QI+fCvujWGd768i
nS+3/btSNHISDl2AcUc2UGsF8Lho0pVS/cLGoZ+46rjfD1XXwOqSLNztKbJER1yw
nOY4V9orfYekJir1K3G6rienBJHcwi3SW6XN8MiLAVaK+N4veco0wFXPH+tHFXUI
cIeI35YPSOARQs1Fi9hNxSFdmbnHyd3GQjrLyUNe03Q6Po1lo/EFUM1buCfJHu8H
xmdVx1uBT32PWy2CcTwWOkgeRDpsTTIhaG1Fbk/XogRbvZ7zxr29zOkH9nc/stnF
f/CxcixO1tAsHM5UDvr56JAR8dCUAlPSieHE0sGfsftKr+L1paOwSaIic5tzfqRc
2cj5SPRA4Ydcb5Z1XWf3eY6fr3ze8CWqh+KgKi/+nHpPrgxvyDcgrKbD0uB29/f+
SHvm1ieCh+MTuqdV+V3KQGIus83z7Jp4ogRnekDpMI3t/SPnyKYcIqaxaQBkGR6G
Db20ymW576aDmwxaBbcCO6k+BGQoqJRptXiTmXdkrOZvY+t95rpD3xrLjvXXsZX5
4C4nT9IhPTS0kU7vgTa+/N47GBlOpamnjpZkkaZzHNgmJKB08iTarHplkQRnsXvU
3YPPnrYggEdqgun3lK1ay0DQnpRD+vmpP+LKTsXHKIwJDZjdtGsi7/Gt5aD6c5k/
a3QWtFS7e+3TZUm/O771XdsrlLhVRZiuRzmPI5KiXxLRF7prJQ5chaQ9vW08NqKk
4ygunAcRlWrwNbViBMdawODVSQ+7cPCjb/UGch1IrYfAyLTcG6wo2aTbVojQj7MW
sI5NkKGit07yolQkkJgy8Cpn4Gc9nrrCEsvahYRLs/c64U+p/OAdU8DHy4Fh63Jc
Q09vNdQ46nct324jQhIV7M0LpLpeEfQDgINaj86Z9iupucoHkCbdHFOG4+xnZkFg
wZyCtELidUd7rCJ3x8hFFB4Az+VQ8I74JkQr85zpcKU4XLN9XDFzfl2t+tvWCZ8G
pmFSRneW92bf0Tjr30RxsPDzUshWrnIedtCDVMOfA1rlg2uaWgYH/NKRoTJUI7KT
Rts3sTP3diVeKoxBnqlNSz8NOzDrYOXkPhPW0+5736CRr7TFsDW7HBU2Dc6OUABN
eqyZamRNAi+c5e5dmjW8XrUbIVYRiUjwDLgFXvNvkUWLEAMXJpYjtgL8hH16s/Un
nLBHbUeToHRyU3+E38qA97QYyNjRPPj2nzXRLUMNN0EUb7BG/QAoBwHsktFRdbiw
Zir/sS2X26g85floM8pKQFs0j8tZVlngyOXozNlOFVutvPergpN0idYpWGAcuNue
eh4sxX4gou0Fb9A6x4ZV7XQApvCcC/RmeqaFFAP3UlnYHxu8+xrKeC2KPzR6lGfK
T2y/lukHaJtDKBoRUTGJbLxcrXWCqzMqX5syaNmzRI/yjsQRJe3roXk5zwhZhcEW
/uxgEpPY/WXkirjeI/B2KzJ0stuoHfN2bq2yAj3bnuxBVCMHWPIb/iYWcWHfgjyE
6nchIxOZNEjXycxIFdIf3d+KEQDJI6PYLJIfI6GWECKuIuasVYoYw0t7Zx/qHL4K
gkIyA0HWvyrPfHAiwwAOCOxv8kqLI2CCrSxtNwVpgkUB7aiLyxNm9hNzmhbUAch4
9YYHvIzOCL2vNX9yEyJtA4ZB+T3p7/Nkdm0hrwQ/Kln/LZS51OLAx9RSGkY7QV0Y
U+ihREQPf+S1zTzBEQFcPaVj5eMVbhlEiBQypKBrckQI6fSQ8Du/0lTp6MIQcywR
UrwB+KZ8bHvT0ahUOF9pI4DDKCsqu/CjWnFCWOOxTt/709wH+T3JzsbOAkaT4YZL
aj45xn9EZxBIPt3avYWsfb3wUpm0epFXp5QQbXyb8rfuocfWrR0cjY23SUg/Ds4u
f5d1xmoOboOxjKCQiFiDObnguVF8VyikKFAW6DP5Rg8X4yipxYsvIyTEZPPiNyYQ
MVsej0qd89LsQ1nqp7l2IFTRzGNuhEpixngCFNWeGkwWlnZJRFLp/eYe7y+mr2Jm
cQRkEmKwcGAIKuisWrP7PC2lKKLzz+Fyhi7mtHBgMXBRvbEeNq8uLkrapwzzyQv5
zNr43XytoeS8EBGZzgCWZDaD0+oJSzpnlp1YPxGEw2EXnCbwz8853qWPpteMkkE+
JRd6C2JmT9GrnPkzhyR2euXj9xaFPcJ9FCvVh2kM55wa9G1Di2kCcMa7QSvbwNgu
FgOGc7jETKtglnsvo4AICQLXAzLmbXtUMd+W2PccR3OA7XCJcKMDHzKAecxH4ViN
rmqInbzVF/664ir+ctfx903vV+jO6pP32H7wlS4Dr5SaLLSVytQ9FgzpeBScivBj
+dCBrDFhR8XFz3UtqQUb9LxQIoxoG3h5Da3hk/KeNpsND8wtBxsCP3m0MXVooK4y
V6Y46pqHpTrB+DfhrhDVkg9/9Uc+Mm0fpsQ7y1Py7NLXflAIjWBcQAHrQMwufT76
QobTWyD0Ihtt2n9vY7PX5jzsKW1HLDjOSMwjtDrEC+K7jaIHTPWgYKtWPl/FqqPr
/MrkDlgxkX/iUeK5a8OfWk5chF/pufDun22ue2jI+GzDRHoAnEKLebAIAA0efEX9
v1Mv9TfRAFde/vH0K1TMejhPzQNdgv9BACylmhgTn8fwt0w1iV4Sx1L51H/8itDP
v7UUGmkFVPTXH/yKyvfdyqmgk6oCsiK/Yg+8pzEytfQFZW4fflC0f3SiGaiqgYgt
LqYe6H2FYvrxrF6oud0K9Qukw0VK1ERIRnZdsS7jk4+bfB64oeUKT0dz1zOmNQNE
Ad35WEEdUtBaJ5WnTrGUU41KYqo9UNFRu7ZUzjziS5AhSE8OfCCdaunkLfW0V4yS
moNIjHggKQwp4Sh32kOWD/e21am7hIhNdJU3L8oPBG5trSdB4JDgKmdypcVQyBiZ
L4avfSlY8iwLh4KWSyDNH77G9ssnNJX2OlJHV7fe9pzROLyyzBRe+I6JPYk7/5ZE
EFWcb/VoAHdBRGHPzaZ5wQzn3MAIIFv3K5GKjUblej96QzZ13NHWFjfsDtTLPh+A
FquN7ggdDB8+Tt0Fk9ljIvC8kSui64PjO8AOhtvWk2qgJ9sgp7ViBllU89Q3sWId
8lV24jqQ5infErYAs/i6ExMsyRvhutyFZrl/U2qAiM/bGW6UiniFAwvoEbx8rNKg
afJd3S4jmWA+UEg3XW/8AjVyKBXui5SzSyxD1X+wyVZ9z+7q4+GO0YBEuJqzUsQ9
HbWpQBrOR3NSXMQO8yzYay+yHwfiszrPvzayEGlQuMPNg6mbu1JPOrDNQwgdHf/l
WSQulc/1cF67gwMkji3i5RFkqV+CFBnpTt4TNvvY16/FhBeUPmVpif01IEwVcjWy
nZqDEJ5K5TVHeWyahf6q4j+iBuldGHf7eom/7rtgZy4CMHM7P1auQt9lR1mxYAZV
fypdIb34A2TFlxjwaUY53XuyzmiVUBoAQZr2yhDwNiPMhXYUQXBStmMlB7hBs4rf
GsBJFUSVPbBliBeo+GqRgGcv2HQsbNXmg7cKE4ozkikV2JwxDED01xMG11/0cJbY
2K2yE7MvrmX7vqtQqlz7gpjbbXUaVPQ4Ul6Qqw3j4lBLFJOzGdcpwSJZ2yAeZuEP
5eczVGi7/FEVk1DlSkzsAJQq+bIfIhibm3lh51tPkBR2VcVJNB2cX2LnYuYuKQ7J
J9BpPPiimfRI/3SED6IJKd2jA/E5VGvSMwhBbemGBIImVYXvmQOd5lskhqRjT9uI
WJYSpE3kRwsDOCJFH+aadqfSCuFRbVJXZtzqXpK3ciT+aqlpVSzrW5SIFgbozDtv
GF4+ITaOtOJ8rPwPwzqoI1WHd6+hOwdLCS+3Ums22EBxCDuZwtJvUeATnKGdkbtN
eC0zjTOjOODrAiuyg7rJ2px/pVPqmpz1B/zHIN0h1OyI+7Xw2nAvlrDAX76KZ+Rx
uzamkD7EC9SwPkv84BdXEsNCod4XEv9cbbpBBVp/+R07oNG15oZcdD4ktcnEaatM
jG2Lc2Zcpof99M5IKpNArdTaIde5BCvimh/acAoQVR4v8iyGdRsJJlH3Q2FPnPwv
9oLWx3+SjJqglFo9BuxKiTZU9qQHK6D2nPUpCdUBGuK7Yu931xBZe9TTaPWQVQnI
C3Omz4tHQvn7XHi7XOVcd5AfwmoMGfK4dyKYGZ7NhzeLKRaf6Am2M3sE7d8yHmpk
DlZgR0Yyy4TRUHh/rYDNMeAnP82MRRK4ncr2KcErTnYzaIlu6dtAbnhEnf621IDE
lF0EwyKidsB1KTFzh9fYrzImcaYGxvjIQvwFaZQ4CBxOk8zyiHR6XkqXgAwFRnC0
E31wL1eamEAH5dInyMtGnKfbYsHSbH61LvYLU9BSrleJINra9pwfcE3JMnwb+Zs4
a9RnehFi/labgW8SNp+nxykUI0CkBP6iyx2uH5BfAigiPFYwfip7TIreZW4UY3iH
ZxnvvmIg/MDqXBhrfj+efDDeLjtuE/yY/kwR0pzAvGgQ4qMl85/wO+PKfw5qMvNR
d+54enAClASSryutj7/tOs0yOSVyJmEI5yJTonAtMuEOyS7JSZFWNdPJHTtV7lyN
mTMYb/bscRqankKhLxRYhIPLNOSwTqQNNWhAkWLfLVCA325wPR7iFLzZszF4dbVI
zciJKeZK1iuH4sZIgHmMEMiBLK23T7Os38RFqzCf3zZjCJdfAbmPKd4Pmu833C+T
4aydwmxEI38TS5/oHvstn9dBG27esA4oTQEe9FkgwlEatyY/OIwett5Wyl/LmRkq
QS9MKo7tmqpWysIcYHOj/2VFS+FPjVl4Q5L/ZRYUPYCZtZpFyYlWl735My50v1MF
qCgs2bsKuybj7F8mer/YeOpgPINSuVV1aoSXF8ExIynqTnku+bOvwrs5uJ9PN8hG
OD+xO3/cxVFt4dc+WlGIjZBzhSiCJ+bAALEvK/vjAZGMen56u3B0s/7NeaJNkNAh
DRiSZg5M+DufO887kHsTxZF7wCWb5rn1Q/Da5Miom4iVfEE5ybASGI6HMUh0kfrq
BCuRYHXJxl0g2v4ArXbuGpALkk5Yk/mfyxtj9VONgjn3omAmQWux2DXhFZ00VoqG
MFaUNELqar1vRGUilnhBDwoOkxZ8I9wk3h1UF3NtEwEMkYfSo3iMF/qf6/tSlyFv
A2PcVdH6u/KDBPyb3vFIkzllQoiVB8or5syt4ZnMrZiNtduZ6vYw/rwlvfVXRmmN
oxBSRtkOqEUpYt6iIudPsgJAV321UQk7jDDjYwuqVgovx3qZussgQY1rZh6kAUvj
yiN4C6IriqMqXshezAXY+nUuJr650qPuh7mHxilc3nDGORnuhj2b1t3ju0L7iZID
xy+FBJvoc2OzN+Q7dj0sKDbT3e3iCpcse4OXtYUvjRaMkdIgUPi0zNYEL7q2ktBM
hpthSU326XcsdL9xMsl/8Ilgulk2KjkPyGWQ9/yIjCTPk/LMGmfQAc9duYk9Y3AG
VGF7Pc801vIFOenf+J31Vi4JJ7famdNzYLUQC4H80eYLkjDdcsslXdtsQNA6x7Fr
BD1JPyV7PGRa/k5znPDaPf2XqOvkzHGbR4vFhxOITzhc8cNNT0m342Ag29IeKc0Q
HrlavP4BcU9x111C6mRGkCmNlqje+ssIGExea+mKK0Mlz0BSgp6FD3QA5vfphpBt
dpnKPt0qd6DwcQyqjGSxkSodeX+lDbsN6VkOcQPe7odvayE0x2e+sJz+KInlds50
xVpdOPQAHogdL8L4kA0PN3iUSPJZczn/PlFotOL7iuQIrpQceWNezOuPznzHzUPh
UeRYGHiyL3vrgZlSRbA1kAOSHdvVboobcd6z8OA0JiRpmiEcI9t/o9BVGCzUnxoF
0Yqkbav/nd+g1WxUxBwIPLORsZ4XQW6EI2HpmKjiycv9kc+37tNyOJ64DAnD5HnF
aDFuy7osQ1Y8C/1OmxOta6W3svQGZ5UJAXR92naVgAGuoTZux+yQbRNna1ey3S/q
FBI/mw5kA80wc8NWu4cwp24/uk/fbXBu4grnW702tCQntMyfER1RX8jW0CbaNrKa
dNkK4TwAh4DxQRXSXbaUan95JXxfnn6mXX9ubxYX/7IANs+iKnW9P+Y4JqaVM5eK
jnFsZiRh3f1oKKsrbbsrocbRuS4hxF6EW3qWRitV9gB2ViFIosSEcCtT53K5PbkD
0D2DmKqEZOWv1zP48Hfzd6akEYU32vz2tbOvt4Y2MTVYTYhRndxdxg7Sbq5cfDii
K+3utdga/atJMbWZP1R3YYTfrFE2BUS1SmObtR280CoeFagJ9tLVY5KkxACg0zgc
UH5hqjVa9vLx4rEc76CUhPobgK5g1zXBfGvrJSsbXZhvjk6yw42P/ywHD4VVnum0
1Icl9sQoMcBMz7AyYJV4rrEW0vfI25v/+caZzYhR6xJyHupLPPm0p8pktbM/EYpm
EDckAKoHfLZ5wqHIGvBc/NaiErOjU8qSAR0cKimkBDE+o2ORqAQ0oSfDWPq0UD5N
HPr7zcpepVVQ7aQ01g12Q77EgXBFZbiPtzQsAiVp1Q/+dEG+wVhm5zr/sc/JBEBv
MdHXmNv65LMnTocYSnCRpA6vcApqkKQD13JHus4h+MJiBJuBXVs0ymNmhCKYDaK+
RHETEoUtRUpT235GTiVDX4P91USHjGIUZ4wnwE5S8o1JYu1v74HZE1hReK1OWk8v
45fIoSy6xnJVXLiDm2OIsgzooiUImU0/L3dcBt5WRUKbrE986khapCyGd5PYoAU9
S1dHiHIoR12JDkjO7P9jXRrpMD3XX1+T8mnfS5teIHf9xlM9Aa1wJfx2oSt0o7aa
/brtoJMQiBbjCn/y6nAr4fcCFEwhOZlazeGpdOip5sAbx8pfYI/91ubZ43bimWye
Hb7K0dRgfdZkX3veeKTVm8q9EcyRYXf5BcwDLZkPWgimid19VxAezE/C3ZnHW/FC
PnboxE28gpyB+cCOIThjoMlWJuZByK+mSlN+JyTAhSY3OUdEsq4Mx1lqQDMnGn7Z
JB+SwE7QGu0oxgvzooKdJKd+sT6riuiLe46aaFwbmQTepzRvKclh54tn2QIqv6pY
/nMWlcsnExxd4Ww4Gl+yQO4aXJl2WY1ibjq7gVt5zvI/LTvgMsscmWCeeLaNcNnp
80sIJrvOfEarKEjwoR/XtilMxyNN660X7JGiXKcKf2jRs8MfiGOU9K6Z2zSEyI+f
OXrwOPU2Xxh0SyG1W+zNBAjRBbuMzvjkjXiz9msdaFVu0iLPr7wfY8Jc+KvSbjTz
j10RkIZoHla78FccB5+Vw97+jhLvsR9yn/nH5q0AUxCxv11D9ABZZM2d8r4IF9Nv
BAknUrS/eAYGJbEdznVMKRYpnmS5lP607hlOoZJHtulpFX4AOkyBScJAty/WyhDJ
faEL5Gs70KUiQUHHPK/P73UGeFXaCDSKYpEudyeypvnyetQvEdz3WiNDuYtJprVb
e9Nfj6prEPylEV5DRZ1ByP3FY7dKW26tpBvSlZu46gSGnLdR6SQfWQdsksSdGbWt
SDc6KLFfa4Bm5N9aYJAZIFbdEtz/NBG7qxb2C+OuAPjCmV7szpbwZdIVDAGUsqza
Q1Vq79LnZDZJidt/GRTVsve5ZhUfQNNaKrbtQRwzJZ4hJslkUZUIjgXo/UTSttEc
XbqJZm6Q7X1vm9pqPl0hBsGjOzLfUsGJckKVCOUetMyL4HxL97JP25OR5id0zFKe
MQaLzilf3RMNXrgO93KYcWLa0j3y7YlUeGBLPDziU2uyqzaWOPWx2TwfehJeRp58
h+pFFTZT3yn1cuO7fg/bXO71CfV2veAVOW8e65pOtg7Vg1zpn1rZhl8slSiAS1PR
UVbgUBFPSr3HYXrcvhQDcdwP2W2IIpfG+EJNNdwr3KC43xodhTwD/CkFrSdR/Dlj
60PtuiKDfm9cSR2PR6szhyA4LrsyUA90DtIKqynKht+lLL6z3KPFRbBIntmZCl+W
oNEL5G1JdEnq3fUJBwliyWaN5NkuzDVQhSFp89yav0o8T9vISVX5SW634UjkoBIB
++ohnYTFq64cV0FSAo/c2c/YqNMiLcJD/Q5KcEOPoUlvBny7HabLXoWddocmqnpz
wNCdnL6+gLu2+tLYiN/81uJgGFqbuEmEuH35qNNmXYOlfDNKsh8Ar//7jKcF61GJ
q8PDC3C03mDFEzcC/gLyhKh0T7iDVq9iQhhe03Fq6fLaje4+vkvLKwbxpdk7pyTZ
U3fEKR+4zp40Wd+iPEXV9j2qS3G2iCoI6cvVftGDfrdSjVRKd2EaxcHz7ViRGb0f
bzCJQFJ5Gy1tHx6lgXsaTrz1Xp7l2WJyIlOh3Fxn9A/5z+zxi8uW2xp03vhQy8W2
IoD/H/975FrZp3Hq9FYTbLrfdv1E2gPWRJ7v0jAlJcRvK1xZk8eGWsJW+pMn3Ox4
loFnMD5Z5yEW5PcBMaDHPiCsPZglKSRyA7vZ3mx92DAUDyDzhZOvE+i2FtnNEFY+
HvEqMl4R8UKWMtgbdcQ8Ojdm1rwjtXSmwWTbFq25qUNUpPmByaARGF6GgdGm1VV7
vkdXsFYcrh/a1LA+5JsCnilj/+t/IniT0DRHwDqpOs47DkQtxrt6fjBjkNBq+CzS
yVDVI3quy7KThreZq9LFWeixqG0AYtmHaaRbcbS2giMWzOpQmooP7zF6QAvPBYXh
KgZ+DR9ZYNGEsZz/I+LWnWCDBAR668L2m2ygRyX+Oevyehyv5YNZRY1sPgDPV88W
DkDQGOZSn2M7RcCLd0M7fyphjPK3jUfUSp6MjaB3zV3tUoYfEfxkGts8zikHfjC6
8fx/gfDqmP0TeNtoIU/aOwoeJwyDLcQ+CgJJ6JylVzp8JYkK5Ihv1ZlgBKS8xJhC
Gklu9oS5yUwWyrr+EMR9uJvgjsWHVjBSX5AGEI9PTfSTsHQJXYCVKGr8s6pJ9V3g
2CMfZSecGFWDQw4UuGuQvU8eOfRucxgxeDN9k4oeofjjflu1AESmC3h3jLrRjRZg
tmU3Mt1LkCYfK8patcTAYP5nrdc/bSsw62r8pyrVqwrc9DErkRWf4iPLzJXeozNu
RR00shmCzOPx3k6L7662DGcd22SJTukEtZYieYCsQNqi3V52ab8x/1soHz73SyLC
8EuY0vEQGwyx+jklF9B+JGNQK/Jtf5ISKQn2ZHV4yvEGezxzc3PEfP2Mwx099we2
ENXEgVPsZCEzwEu7V5qDua9ME5x2KvQ5SBEg6gqMONKDEdsvrhlsbco6b4yXL2/q
chuUgv5GztJhmuMRqAFRuA86ktmC3QOHYVjtfgsWHQRGjGppXM5Gd4Dy+jnBKLRO
N3u8kNyRwPpqPfCT+nONJZWCxYoF5sTywxvLxajfmNt1ELezmaWVrvjsQybqnOpA
uIbGcpV2TadyF7xStbJTxMTRJY9FnLTUIs0HVuGJeXpUDH0PQAFbjFayoTe7CDqg
3A3fx8Sch19wXiv+REeW+vdjSH8wrZgZqY1LF/2AXtVva+9h+naFFd0TlKJS9dPW
QI/fl+ZP7by85UdtmgiHLLPAkbKQVXQ0vl085wMoV0LIu+qtACoO3Bxaf05s1ta6
tIs3D+E+RBevGnynl95E4xTKTjvWrWfddsEfrvMq0lx2JzJwftT1l7cUuKCacU2f
Zh1t0cp4hV2+C5CagV+StsFPqhSMdmWA+YmfVAFwNngBVfFipFZmyGSFh/J7oLu7
vVGYDG/QS6batwO6cL+8YNr+C0okl0r27QLldB7uYnomTWzyMxOZ49cPpFmV49Xn
3gInyMNf6Pj6HKvhyRiN97uDncREmNvjsf2JMHS5fNaL4d1LlD0MOt79WoPvqvvR
q7Pm/Bz914yV3dIOvVOk8/uiR9V/g2e6KYaTiQBUhddn68Ht4BzPLryciwBadRzS
S+vJ4HZcq6IamMsHMkpZLrQHbPrNN5qNgDr6oE04OtOrPgkSNipKXLI6eRlSx/Vo
+q5UcdqFUOPK9hz7HOATHDylIsUJ+kc9vwtM/nVWm6wP3j40xkezFzjJgehgGmOh
n26VNI+G3S+ewFscvXqqyivIlyWmpZMBRq2u1eyzyaj5nQbrc9M8Ai8Uc8lu/G/v
7Spw/7MRNWNAki+A85gpffF4GeG7X8amBv8Uzp0q0uJKpoKQi1YvbJCldEhR8OfD
TfGVc1eblp0EizaLkqR0DnHP8+jbYjr4U3xASQDu0Q3lGTf9BOs+JMpC4fOIv4Eo
LIpAN4huKd46jcoFbm9hmw7Z1/3Pbje3lDNEE6rC+tSOHIictc9j6z0LAH3ixe4p
Xc0uum6Ze8Wo77Fma3o0Lv9sR4wkjFcFo6KrO5Bp1L2jFPFYZGvUYKkC7HUn89wd
HPafCCXmz87s9vBtCFgFAMet2ueg6Yl+gjLHZbNsZIUOzR/QZi3gUhtyeA9swe18
aMiogJ3ujhaNgk5re3pDGDmxrL2BrLgQL2Kr8W6tuljZBTUmgIEKJrmsEAbG695f
PfFUHc2r8GpEtOPDxGScLiuW1aKMMMUXzn5AuB/ojK8y1a/sogXLVSFZcH47pWr6
eicV1QSaFwfsqNVyurwV4s8B2wXVnUcbrrPw1d/S1Zlo5Lz4vlBTuRdNTgu9lIKq
2UOiokOSW5rigP5DZoJN4Vv3Sm5wzMPkV21KSh9aDMMstcmk1etmrWIEuG+Ilqkm
qYVaGXfvI5ASouPmanX/yYm3suGfCcyRUJHiaFIBsW/2kmgIWjD1PGomguNoLP4f
c/Sfi7DHnV5EQLn/8ShNXVSwvus47If6DvKmygUcLEzU2HIqRMNBUTkjAiwOoELd
JobIWJAL1EKs7es6jtwzymyxyT5Q5xeClRaFCpZcx3iCBO2xNI0H4QNsAzFrPr3P
Z2rt+avYuii8+0qnliGZX4NGoxIq59QEBtzD0MLlk8Amx2MKvLHalnZLg9yo++Kc
DUDwH1Kt34Qf4vChjqBbNdpr6bp8BkVtcqSz39nUjHy0uDEJ+0O3PZL5eVwrkrwW
bCFKAARQwEJtv+ENvFG7qWq0EEMFlwK32E021tFhbRls2MOlmHXDTQ6+F1DfVTA+
cIuOLcGO56H3/IXwEGOiWtqB2zr45aJGVsu3CYeSXdC9ekKa8C/mzzCwn3MsiOTH
GLES1suWs+Y4T0Bqo3g2dM2ISmkKwWZ3KvQa75K8PJD2xTwTiz22/oW/1Wh0XmEF
yRszS/CezxeU5jmiNSrekXX05bXXXG3Bv18E7bgc3BY8naTm66ercx8glagZNq0l
mnI8VkgPwmCZ/s8+GQ4KhgrCKGJmiwj06F0l4LISmFARXmB5nLhiNfvv1zhoHYYh
o4n0OqwjzAx8zNKn8YW8Q0nPCiRIf0vsigBH/W5Ymhq77PRwMjmEndHa+ooIOK6s
gAx6bbl0UUfFXBauS0ZzPPM7DnpAYitWNZsenZJU4dRKe4D+rpbtZE76m9xDJh63
htenpfkbo7To3J2WLKynfgjthi1VV2vATTUo8UXJfW7rDiMDu9kRDcNjHqn1pWe6
mL5OylKdGspxCNSpwd7o565dOeJxQPc58LBm3ru1WW4YtfNeF8qui8bqopgsq3lj
gg0yldlA5oF8gVbNZanBCD2j4DIfDKCmUMb4CJnxBwcL8LezHPqyZvYgOLdJIChL
oivFPvqq5r05P77owjrd73Oo1CKJneURmJONzP0aZAlvA7Mktl6cJcg32D/vQh/v
WXv0D6e9dwdaGJhbi7b5ip84LDhNvERfkHTcgqKrY7SQDp0AF3RxA7/et+J1JGGC
O+46zkhySE8k2YArVCFwAqYsorZWCbdoIXdTxWI/0vRAB9mrtRZXFyFrMK24dZCv
v9LWmEps1SrOHCbBv4hF129pd5HLQ15AumtLVOYe/NOB4Md938Falh4EM5WUDgPL
ewLEwSkDDZIaxUrxznKI6dJe4yBDgZJCwO50A39AD3UFVhKGLPurxABBlPXuQOLV
AsU9jrbf/bz2ur0d0xTWqr1FJapgtSoEuhSAlvwekx43UFFN2m4De4gQnCKRxikp
nMp9KBFg2Vkyfd5xMTeideJ2lRySWqc7nzlYDS2PKyrCAnQb1uKzwJ3yiFCXZ3Eq
KNBNmMSdqR6WlBBdxPzxb1Q9YqLsTQYRKnGD/26g8ZKwt5DM/ZFDNskyf9hd4CAi
cdyPYS1cuGmWTsZBYxMNeGaoow1rdTvUKBaov63pDS/VL1BAr1hK4F20QdEooUa9
NZaiiR09v9UsVo1W2eLpL+9kljFDmucDAd8tC7vfDPUWQkVQgLvnb0TEkLZWXXqP
vJq0y2wpCr+E6poYyDfVIafVuWZ4ZEcq019Psl5uWOWnXa86ySX4kb+pNlepgVph
BoKBGDE7U4tiwO32Q+E7WVIcKKPsYRrk1ljFPKOVUbjpaq2SX8N05lu4n7gWpmx+
MG29uz/jaZHH8Xh0mkqYK2fnGC6fXUJbtCu9UxkL/eJOntpdEIIfPhAFL5rNgPRL
11apAMh9W6UfkTSSY4qqRf4WWPZnYsZPTb+KbBo+q7Y4mF58AZmriqNvusOeQQS1
nQwkUg9tN4qwQfbcT/D4zx8XGKxLPZSD39WJFG2pfVnGMQK9TvBrsFva+kVi63oJ
o0OJcRa2LARn5qyBnoei/oF9gdZhlTNNrAi5KCi3CwimHMLgT4TH746vEnRAoh4z
xra8/tVrGOyPQc7ydwt1MdCQJNjUp65eMUkF/9YbgbI4zRJZdWffMUhlM07vOiP9
XRFFUZbHhSFN5NeTjIKN/lruQVn+efV2yoOnJgysovX+RfmTcXGzWo7GMHoGFS6t
7oWKPMEuqM4M2PeW/8UMkLuazFCEn5CpYfYlGI4C3/GvrCIWUvs/gYWhlLKfQLyI
xZs0a8JYtDAWHMlweIqHbo88wJiXXY0CP3l33hXmwEGZJ60mv6TpakWKuC3mvUWS
j9QV0QyWrtXs0qERppj7UP2PFYNiXFxgJLanb0/M53/vlf8WekFmoAV9LBKVBZkT
emXYZElqSOamEpBBOCwCfn0Z3BK8DHx5EMx8vsFLN/+g9qoAGdBqztcmY8uXmqRb
TLy8sDjTVWSy8g2iAxwh6ehANwuhbv1jS+8tdTR3fWKi9iZmh/CaBgxmnJzX6l+Q
BsSJesuqvliuuNKDq9hjQ0tR3kX5RxzDg60dkneClUgJCX18T0tYeDlKe9+MHAQ8
ZEIcXkxo1riD6tlHYtdFLJBTjmXEfvVh2ZJYsoPmhbsEQdsDxidpaaAesrSsirJ0
stj2wpe2Y1veQhbFAJfKJu4uC2sF95WV85piAm7ktZzFSdVmoMpxoHb/qynoWhN1
UXeKCna7rP9clXG1RErWkLBbNE99XkI6wAL9DxIRUP8VMpeHLz4f/Hb8IJvhjwbJ
k+ybELhzGDm2RgTJeidmpzOD2TeulflwV0ix21UJcMdqxpGd5p5DYvWGr+lWtrsb
AQ5sJK7njCeJL/CEqrHCJzLGCEMSmrsIrHsRQInaTp0Iq7DzpLRkZEE1lJkwjDLp
odA6yUwF33xxoojRawCGhd6tppo5DwS/6r9Q+dOQtDeDN6S4+9xX8+Xotct33FDN
SIw5BqpyGjR4t095QvQF9aLtYZI5Rp8S0lO1cNAJHNmyAteHgjuhG0tPfWY7yx5c
98XCZNQw8qKv2wv0M/EuClesEOutbRDu19JdU36Yv37U5X+hKrG3ZDtVxThUlnG4
5jY7EAWFxQT4sJFODXhAZtyXH3MzkxMZ7eTiRFLo7XsyxJ6UJ3HSv3qx+d+Kbr/s
giAVnWiJ/TzehctQNT8N+O7AHiV1aRNiwkuNAf25aNIUoj0vmr8IrstbXioQy2a+
6O3nWVv8Xn0s23NEP46pG3neqSCtlXDiXmBv0yVDsccg3JPeSoW3qluVMVYPD0fE
mf4IAPusJmGa19pTGWngEKBfjcQ781PWGvnrFcRK23cOyz0unVAbByOLDHxVNBlF
2zKpofiN09rS8P/E+aV/FGdXvvtCr79n6bV0fcobys1iCE0oqI1sXqHSNxi59ihD
BR/fGSewc8DqI3ePTGMMrlebH4pMpkWc5xTk4p+ocRo0wexRR9FCQdLHphUOPmdC
wL78/Pl9umc8b5gCi+lsJYAWX/GFYvj2LzTC3xlzjdPikxu37Uvi+SQdU+nhq4uc
edlek2Ls+ggq2JFyWSk5cJmfEJr8GDc09W0vJUdW0rg6r057Jfo2YG2nMwNZgLp9
Q+MHpyt1gxD/cypdq8j0hRaRSh3t0RybMqfJLDc1JIJzfuGtfh/WI7jJAQHMS3c0
HR5v5iJCXktfVC0IdSZLkHx6TkW8pGN8tkHaDhE8HJyIFs0jUh2jU2Ny3jvJlLFq
N9elb39EBTIl8UoXTt+Iqarq4JndvXEnlMCIAgxKEuIkns70xp6QgRac8147A8xj
SXlY/rtpPSP0yUDwbPn2NywyygTOa0V+vEIBYiF9MaNo4aZIwbMFyUKzvRpfPgij
LDG6WwYhTRslOCzB5tHk56VULGxsB+5XE6na/q43Pccz1dVGg7Ru2rPX96dUgX4R
qL+nlhlOehQ9n9MJ98H0sPjL2bG+ZlCYFkTAeKEONVCwuosZAEaT75vHpsHaMktz
H2flGBhVhM64wXNJKHdHIyWtlxPFHSsHzDCzSVckAKShPuSmPvRzJU1UiHozpCEq
mN6pFaUrN3CDE2PU6FIxlvj/HyLGC2N5bMMM0pFCeS8dAAjDBDK5QW9BZ4PdSaOj
CA++K6rI7PU9h2wnSvX4i0EwDUvvAJmFnqZeCdtjjUBJx1BVDB2gZcBfj1AXd5gH
Uf/NkJKEB5S4m4lQt612mhSMNcKisadarOQ3nNApqVgqYAbZJ88hOEtgsABgI3nZ
OQWOP/VoTIRN2zrNG6idZ/oJIex+IzGhprQ5939SRgN2VjpOVE8hrFO1mRPX1tux
mvVteSl8DBxJ1qUJX1IZjXZwyzyRqN7eIX7LvGuQNri4euYI34oS/8nvNjh9Pvam
vHpILCBFSR4tM064cdMWKKgcwJ+ZdxhzUb0SElNiouvnjV17u0ZexY3FmevLQvmP
Z3c6DWnlp9CccjNL+XpXzQYKdCFRGl/t2+zYjscN6jHQVxFWGmqbED20+h8aDgpq
6q3wFaSNfkmvgtMxBidAQdzK92WnmGYtEWAhij4XdruGuritN/yL5VtBvEVeYfzz
399+LSjv2AeMp5msTr0bJofhcEn84g05Icp81aLk4rrXtyns/uuJTkswj+DxN924
cV1p7cJX8ggShfoYA6wH0swO+RlT2ly+PNIEKoYyDbo7C+EYT1BogTbKUbet3zVV
8ByHn5ZhY/BgOkgyHbk/W8BP31ur/4Aqv3APEENbVov38zO8fbvFYxfLik8FI9Uk
TrLju7X44dipU6JQh+kWvQ1DOI1Pap5BbJPQQhF4X+woRbOU9+mzgvKtEwoVZDLv
zQsUQleVQ4uTMl5b6OWF+IlGHxKxvJu0fwfQa74MItSXxkQWGlrEZEudeJdVy5uf
QLwc50RoNg7YVMtwnNrXaawwsXpUC2nyEsWh5sL8JWZ2nB7TNqbD+pSzFMmCAqDO
Gbzu5e65R9cp/Azd+YnsFnvJWu8Ehx1NoIxBiDuk2WHxJgfexkNZZzA+luRGJj/0
VR75XoA9dCjNEqBQlzIH5Q0jhHBTr6Sty0C2adrOOEk5DGShp2cXeB87GRNcJt4C
zm9B3mILsauo4m3jocIj2n/cEuAdsp0NXXTWWwcjSGh1xg4buv8NCH9NyfoJWO9p
GSY1JiIhjtTSardXNG8uHkDCCcB5BzFg5+wQfPWGFO9NIuia8EhAQJFNLI6MfVSA
lJHiHHyUfxdDfdM7wWUJV0nrRH4xlG1zyEI5ITKEO3Vs8ot6QGe4I2WV2SGcvN9k
Dml/lFoz2bevYkibuoRXBYvyd0759rhAr4kZt9Kc9TYfN458wtdi+PJWnL7JBmRU
Kt0suJmyyIdVKEWYO4XFrIJWdfBxJhv/P4QAQjcxoz7SL2cadrlCY5yeGrPFXLQl
IaHshpdP7AibNuGLECDycfckMPHFMR7lJ7f8EIj9S8sOSwLme1uPIVq+ChQXIVFe
ACjH/g7MtAQ9mqiXeW5NTRb0pgoVzVbbq4pdULG5Pd9N83Su8QOzbhY7AiZvKn8m
le+7kL94myC+PILd6TomErAL2vAI9VQ0gQtMBIsvJX+FYR7CqVAsI2xjzUu4/5+W
RpzlsBPrUvLZ81qhSmSrlt3zQ94R8SnOOdHZjaznksyjMF9rME9F7Py8Xd2zbF9O
YL1xskhOYRFdO2w+vbNxvO9KgSXLURqmwiCKuCZgXX2C04nCgK0dLUZs8bgM+huU
Yy4tXqxJfl4c64TVK6jXn9OxQiej31TrDnE1iBw4AGyJGVfe1N2n0McUELqPJp8B
JYafi0bz75LU5Dc+HAHMzhj4iAe6qBah6SKugKiQ7hdQf8L/BfJlVxY+FzeJDPQN
fR5j5FrrAibMxLoVuK5boN7P/isJZ1ZyRbCjyf6esT5hLs/tD2N9AUL6GfUIzU5a
kmM2jOl54Eq7fDpCp21MWNu/PSJQXaCD65JnzKcEL6mVk4HqJSY2GjXjUYmSCSA0
DFmaCQ9jgxa03OBQbNVlfbW2IunLTuRutX+jXPhSxjfuncri633Sxwj8vi4j4Wqk
e03I1friVC7rfTBB7L+VHtpzbGOlR5NgHjlm2Wnvh4muvpC8jFj1xbcPJxG6MGjj
jOB9wT88OrA6vW2itr/5+tT6pAQTcSUks+cfBmjqIzCl5DNiV13cCU94Suq6Cq8e
iFh51AGS+mF/DDvZWoNXgco4XfDuPUhrc/7aalaH3A/uW0T2n1J+78Eqx2yTYfBF
qdBQjv75xrY/YE42hN+1LntJT2IDS7dfOlbmL/WcDqdKGif8B8osA8gLy7dpPL9K
TeP3n5mFmiEzc7eGRYIlNC85N2VX6Hpwh86sYHS9jOXfvRgudTV3vjz2pEssJpHu
Ww0hwJYJyU6I/moDghXVO6IftDAqk1iU56VFJhwsc/YrrdAoGGwTVCxdQ7NHMnU4
1MnVfLXaQjiVj6KduCPb0HPvalWB0IqWseZBxpPwCoycMZqz+cXGNNaCASaumrak
/h8qNGVFhTdbdbsJC/Bbk8RRzYzP510YCUYueTIrAgnDmYC2tkw4ibkssXN0IMwJ
/H8ZYV20QkkfqPRZZGINwQg7PtHpKCG2OQWmQwCKgKMZbSKkc1q7QdXBg6fkZftO
+y8fiy2+QxerLMxPcDGnFay/W6102Je4YUuxxo/F7BBGbqBQU5I/OtrOrNvqkzDf
SLBRrxQKGR/Eso/EI6kXoJel+JFkpHwwDuxT9LddFwJFEIj6ps1FvQ7whD8y0Gin
9jjOyh+ABgxPH6UH7SOKR+OxNpM3hPqIOhq05pc53DkP2WqWBGbBrNh5O8rxmOJ+
y5Vn2DDAHU+aS00v6sNZy8OZc6kP7MKVybNU+3rr1aLZvg22b4PniG9Do/mqerqP
eZv05sl/xSexvp/KkEwsMZBYckS2Cf6vIMB7NyoOxmKuS6+Eli0icKTUihzjnvTu
Ea1Vf1tDznPZZwMIIcawD4Azklh/gxRaqqwo+bkgr5R5+vLak8gj2fktOVyVG/R6
mrjnfhuc4eqCTiA1fHZyo68BDkCvZsogWN0pEvt5EI0XHtTJGU78c9VNHSE8nYh6
V7aztpIoIrgwJLeYTO7BUP1/u5SostevVjfMdRmKQ/ivEsyAd7/fO5tHyljqXDng
UD7W6JnltAv8VaACRc/+blYzcBwcTgjFQbC2irgef+zPOEKYzGoJuG/Z/cmafmXO
j8mofTHCDhRAvv6iB6lQ5o+5PvSO5Ahmaf8aPwt7CyqJmB0VeGi9eIj4iEI50iIe
163c7q4ZGjXZYd+2V2SoEYs1ZBSXpEPmsDLcw+XAlQ2heybtVtucHoA410Pbr2xj
MsEdljKrQboxPtzENpZRbSgYIpNjjeTog1TZA4/AGu3KzbcLgUv5NeQSl71DgCh2
gwQ9+jDzctx9l0UDAZQph2sVvunMkuY3FKoQWSaSyeG2+HME5AE9egfeW7k2FVx+
ksATYpGmoL7o+G4iIKeudc8Yft7bLO5+JiJMPMuB4EfNHxqmofmp83UlOUGGm/vj
NUPcrmpuCHU7cdaybmVZOU4KbuKOmG+jFPuKyMXPy1sxZFXJOM6eMkh6JtiGQhtk
VLaNobUJz3aUifuDrclSnvcBc0cwmSqZ3KW7N+Ly3WeQe21hmj2m6jiwqib0BhDH
EJ/eg4m1jF2CSeeWdFkmk8TbeMi+m0+5j3+BX/aDmi11fZTeBXc7b4lKNBVfuj/F
pAKo2u2MRszKOtrZ6s3lwcnwd3XLNdkTe3ePfgSg1tOTS7Hn0nXvMp835QpmKw6z
1I27l/mfc6q7YsZ148C2cHmA4ewUXTkAqtoD773l92SkH3x9RFdewgLeCxlS7wm+
3kvWyuYN5p/1MfX7lFNnjjhIrgsiT3vp8Kl0vfjPKKWj/qQlzU2e5N4TaNg/aTyQ
2G8DHZM3WkLOO94GG1ajtqCgFi28wnqCShoBZx/y9nlNPGCN+j1N87ZN0wL1SA0M
InUNtY+SUf2m/xOaztKbzw54o+MrrMaFbTz+mwZVZyRbRquk9m03xm/y4KSIXoTj
u9LVlfjIXmduAJA3SOxPjWVvlk34S5hr9g7r8gXiYSmQMkdvq5+5aXjiW7psy4i/
xIle2VfV/LtCe/9nGWIVNRDPLCgSysUBxhpdzwkthnVWxr3DKAAn2HFkYDhy8ZlR
spOmrQzOWj1fUUb5SUiSbpv6J1MFJX7y4vgYa3IXCQ+XVTDNjHL7fJStXdw5FrO4
DP71H13/ft1ZqPrjDJ8sO65abLt+Bf7pYUA9S6LhhV0QV3xA+HK6xtOHA+fvplJC
ntQzkmSX0m/WRLBEZIMdXjhUMWjDWRQ2ZD6eddVb0lipjzCDqyvHV6AeNEeZqCjj
CYoeDgQiqbBw7d4EQwKTWPh2Hp8DQS3annjx/DOu+vSz3lN0MdMnu/XPP5k3LVfZ
52Rl7MWMuwXM9wzPHAiLKb97MZi6lFt+BRRsxVF0+2ORq8JNkvx6uDpwUUmInmxW
41hj9ieCuZOu4OKQZW64IXO7sMsaiNHZ/L7icVZNdE5SuIGsJXtAuVGEdkSPtypM
fCvhvlcCz+O2talNGjFPgR+HdD4ss5NYgBGiosRNRt4nupG3QDJoUoHrgpGTf9HB
rIAT3nDOTq6Ugm37Or+GuW+92wTZF8bHVDnxO3LNkTiEXR0L7LQk8XVbpkQ2Oqzt
mw5KqzjKXkzpOnHYEJB6BJeHl80SeJcsguSqoUCEMjNWIA1kn8O/El5idrF4mfn/
It7B36lojaaCa3xSyYb8rG7gij7IVuGYzgTCgT9GikW6FPSn/w+AzVw84MvvOfp8
s7OmSMUfvIRocu/JhbnNFp34FebpRCt4tZiku03T6RBuyOsmNQi31lq9/bbZOLU0
0j7fBu7+2qObrzLe2qmP8TBJeqbygJWstAgsUGAd5vvzpjUAz7H7CqvQrmNlbxKq
z5oiSkQxKpL1BPd3FDEea5uwVFbn50FfNXvgiu9/7n9+pTutBiEwVa0m5QojX6kG
bbJTuCJi7JpEVOla+HcU2Umwzrgc0eY+B+fwVXJJtoxNqoFG3KdHaG2kq0plgx11
F7taC1qR5IY6I7r34BZfosrftBY0D+Hfw/jNYwXAnD/8BPmCoRf1AS19t3v+g8XO
hFUNOklH6NdhoDJQDFLndr9W2Mq06x+Y71aaTUrH9QPPs9HCTiDPfeY9XvZTX0Eb
9VtIwSkqE5H/FRatFW57D1+QIhtCsGcj5teTK3IC4bEz7azXWzbTET6kP2V58FqR
JYcBngGtwe/1g/KR988AOiJOjvCS1T1HdV5abztckhUZIsv27Spd0bb3fyYu4XW1
R0pj5GzgtwQQiF2E2p2jv07bUH5+DaCxUY2RtQeUys/MDtPoOZP9Z1d7Su/+fMI7
5qGnVW4PNVA3SI52HF6K799+ez8qng7LoTnNWO7Ao/2Go6Wu5/Hx/6sgiegLQWy/
L/DQWebFcWTvv6ianNAYsGmGN59pof/qN790Iz0MBPgk2WfI9Y3ZzSvFi/aUpnP1
fGPzJlh9abD8VaqFCq3yfZx2EI12iQ40t4qboGmEG9LAQ92/O6L+ASdR9HfW+kYv
K8Lg0U7wvqItDUnL6EDbjlt+QmueeeVNedSzmRQ4QeEYFs6Srq81M20luDZ6+65+
uOI9qUi/KfHGnL553C1KwfqxOkBQu0DsJKAzF2q0FEyOmFJEkAwSb/p+eaqV0dbG
HpdbJIika1pXHv2T6yDcCzHYa+74Z7SQD88kkN0/gBiVTOB7ailntcwN0pk+DhSK
OjX8XwTyIip5hlexgTsfIIfF2xwdZLn8P7WbVfYtUPWxBpF+G0YFerr1cti9ETOz
ZZw4PGhOQtL/0RbVI3ro7kE4s7e4toMZMFC/9euX2950aFdwAxYPsWlq+khXEnqN
vQrWF0kCM9fvU/w8QqDeVnRCf+BtYFyIakzxMcx0NCaWQXxbQU3XWctlkWPrKp7o
3h3ySDWBXDmMrX3/BTsIM6sP65824JxhtQT9xabMrVJnWBDSQdV9lxFsPJXoXZrQ
7bS1yLcT5o6pYO5xcNuOvYiTFE162c7521jYKk+T1mb6VCpD26phRFK/jlTrvYOH
tgx5dw/t8/5ceEJXnG5hQfkUidVxfbTx4XYormWMaUvbh+vg/nJlICSZnFn7F2y/
DFAZOlzUBL9M4OgPms4cCcp2y7+X4xTRF3ZjEgEeqPxSBWNDmLMFz6IuU2X+5WRT
QulGBJIKS3FpW/vpdZjixbKwjKqHs8lhBKR3IVqNZxLBBr40tKID9tZ9FAyacfUM
+OYk81stSjuzEEXN7heYT3gtazHif9GtzEv+wl9078wO9vRfyA7Ng7NvAOnRcCZe
f2tdUIuj5wTqBeunv1vFsgTx3HCoqlqvSxFUJwaJcQFfvWETgjpHwhNj7Ndh01LP
Ddef9DYedOUuDs8Gcsa2UGeS+PHfVHCmJQRt10tnVTnceKTJpuT95CKfzp3Az/GS
WPneWCMfzPn4zVIm6r2BPuGH0URaESSTbY1hh50Y+GnRvL7mXD4s3uz6D9e+4mYh
NszYxrn+omXfJHIuKNpGv5cEM73rlUgHoPrdKjJqV6QWfbDDWtzgdaGi68G03Jpt
s5v7YSfzvtF69QARo4FgRWtQ3Ar+Zu8byJq+S74wE2IdymBNbrqM6J4pYJ580mWD
VBsyVLnx/MQzlQiRC7gC2iJj3lwMQUjrovbVyoygkakchgEV0bE6/CE7ZU15uRS1
C5Mh/5l0Gp45UD+goI+a+QfTs8h6BEzygPwOXLqqwRMezCxloWSEEmSPL3fIMWBS
0SznlwOrnR2DFBObEiorqZ5iSxxJ0+onxstmwkiJZtwqmqvFI6naw2xrGlAwQn3D
CEPDrNRiqEPhAdkVHl202QAqGQ2cDH5hkN4QRmW1e5itpRhmfYMMA7pctPx2XzIb
ULQLl3bCibq3RxVLLhWVfYXNWM34pta9RrJK7Wdr84VZ0hHFaDkRwFpap7v1uw4O
QV6LyIIyL/Atq/iPoBA4sB2KgF+vvrokhZqkyG7vgBqVaqTYtxGUph/5IigDa+dG
eqqrUy9i8XbwyUyomWQNCO68bGoyIWiORKBpgVjGydIQ4KBpykcu3rp4qEGalBzS
wrUj/tA5XtFeWEmB365tsUKyI71u0zGOniozV+nGnLYGh67g0L/KRbXqnPLV4CRf
BeVP8i3qtEUeZuG8FpwRqTKg7Yh5o+OpcLw0xBxuZE87dznhG95Jq6H3dZ/yhB55
zL5D0MKqCB2OUgCFkxqGCHzy6NaBiNHSmmUt830tXlspiJgDcLnTRRxbhWQ0VAs1
P22qSbpHteg6M+M09R24Bk92SqNYEdpzS2VMA+ZYokbbY+H7mHDYW7MyBGnrUeoV
1uxUmmqAKzFkQH/o/MAlAyn7pcCDdo0x03G0pT/a8Ve0XH6l+MV8tRv6CGLbvPZZ
lDMph7uQwtpJPF20Av24w30VVyPOfXBUJU/td1ell6MwvXWYdeYHtFeLqAtQF1Ni
nmnxZb5TAxu9Wqy7JbjpM6YVRAafQdYG+XOK27DjOMdVf7aL94MOHa4KPhvL5L6x
fIEBQaQ6+mdLaeWK4SKrFqV4BO/bL9LM9C0azspwNojyPvMFVT5B1xbb91x461hF
xWh4ey4njNcIjkkNaCMROTPK8ijd98A7obYsSZKHhG5IZ3VdQ33oIlJ58ukKHz15
+MqKqutpQ8FGq+GVJBhdxHNlO9VRxp3Bj0raFiXeXk52ZB66gnST2rEeIBsEz6hA
FogROMxsiwuEnVKij82EPqCYMR+9gkmuFxRp5x8mzyJOnLBh4S19h4T1Jv0kiY3K
FL3UqMazjHQ5tRJj54XyPeLYjDyCeyJtkWN0GuRHcctYIUvLPUSLvpfaxYDZp9Y/
Nx4sdzLe14csPMaXNYGvlX//FJjevln2f6mkgnfQGARyB7xo3KxGC9skUgZ8+aRN
5y0B5FOYz7Ql7C9bxEPmQmD6p8nBRBG9QRsNTd7NmTekEnO2WgscIipEzybzZ6SN
5u2BaDMWD4S00cf1P+Nniuxp+iT+dXUw8QkE1yVu/ocY5cbkycJuuIXhgquStOyA
5TZFZTafVLnpaOmHw/2omm5FTskqkInVzKtUqwBseGo2i0Z8DoglqSsDLg+cujiv
FmaU1UwoH1oe74Y1xl8YZglOqzKDydY/Wg5Tlm+k2VaGVmMgkkbTuyz8QKn38bNJ
W90dsFGeHGi0VXp3IPtS8zG8Pel1dg00+Xwaz1gEB5LUvWlpqeLbSfFul3bGEzca
Gr+O8lyIDmTCdQqiScwKyiT90V1qUv/jztbMhTsZuZKDFBKnPByby0gFURPBItFk
4ftQ4vGjLLVHXLxco7qDzLr2AksMCTMkbXevpztCCBVJFdAElGs2mYe5c4B1RWI9
tDZL/Ek0JMDu2+KoiWCp5i6/2lneYl4a5Ae+sFkHDY6hX71/SlWGQQVfZJbLr21W
FEeTNlOu/GkWPdWmFEAW5FDu76oWUeOQDy36wwMpYsRKucAj0VaMexYSV96u1npq
oLWMFpWbOs9BjbJ6auWARxdDDiczxQvM+0sEphqaXRln94EcoyvFT0CteolHwzmB
Va0epJqEWic/qZOg50qFG72WBDEAEtzsIAS7dZ2l/REALDAtPFSeAqOwCPbU5JCL
gIpJqaOANTQ9AsfVhMq+w9aZhB22VZDgJv95uajQFRcGyKoAzCCFq+fzXXVsfR8J
/U/2lfHTKwQx5QSvTbpLi2G4kzaHr2f/HxSmEPbiRBmi1cXZ1pjk5xs6rWJr15OK
DX21Lv8vXmIcYCO8j5er+uBc4bhHrBWrPa80hMvLSllSTPY+8Lm2Hgfo7H+pBWJ5
qKz9bQmWcmewxqYK4pvymFQXYYUqNa98Ow3nRFpt9xZsHd4HfNNsicdEzrcWSUnE
7LAi/5Mwq1Pe+QJA2YZOKk7swJyl12cvh1dzkWEreZb68pZefZLD+CGwNHEopuGU
7kK5Xdul4T1ymmdeD67s0QazCp1N2KcjqUiGlCHU8rtXX4uuuzoeEV8y8oiZWGl4
vXNHboIrTNTEHmGwuzLv5VTlfy7ybr1AGHBaZABpdMqw5d2GBE6Qz1T+dh+ISX2d
D7uT3N1cyCon/kQMSpEdq9OUHQIsqbtmCS0mzoSnAf7GlJvyNS1ixv8+o2kYDLI5
dYCsoJ93tyA/nZzqVmBqNJuORFP2M8t85nLEHjXi/7aiF/EmJmi0kYFS3aOf76gy
WUw0UrZ6fs8t954aS3e8tdpbl2aeaDShqU+AnaQ/MXGwhVVo2/5E/Nq4loszg6aj
ABdsLpN0DnvBIYgmAKLCuFneNmsnGRbyARjcw/jdSFMMeQWzbrSJ9YUnpaSw/eVe
fmF2UeD/02EmUnZd74rkLdAz2rr+s2ganBu3fBArHQ+pFopgKdBK40lqkA76vPgG
QNJuPiuVmCw+nbFG/j8K2XDxnhROZBQMEKcWGROuvR3610trJ9p8efKYqkKmjyph
ih7uc1JnKjyVepJ/ggKwOBPXdThOkoWP1HDsqhnaFiLJ1qIDQopjV4zZK8HpnSQk
MZ/UK/b69jAX5qGMfhasUkuPwJIJ8a5rGjrBJlYlUeHjITCk9Eij7/+lWCn/qoy+
FeE+eS55It5lhbmJZ4X+iNlysiFtFpWle+sblw6okxvGPKYoitneI81JHcDpcJMB
uar+WBro3rISta7XflZtlqZpcPlK4NuQcJ0VnTYCd5Y86lR2KsO3etuuxdFWGrks
3x57SW8QkF6cICCaiaBndqLQuSjRWCdd52eevdLVheBrGZGY47xijZjpnSCrFe2b
/nn7DwxQk8Ufy0zvSW3iN2KiQuUnJFwBRDIgnEJK/Sq8nza9zWtX5wmK1bFwUx+9
+/UUAdG0RejcFUWq36PuNvVmndrGkpfdY6g0rm3eMou+Y7oPG1nAh9+tYZMtIw7v
34O0JaTGzEnfJ9tFdR7dPYyR5Od75VtIfz5/2yO9OZ3F+1u918EpCn5e5O5L3t3Z
+d4UIM7r0r5FtHnwBYpwvhV+YvEkwH6YwonreCduC1FugBUhemRCg/nAlQ9oJBxL
6cQhNvlBODGEpy6SBuVtiw3wK8fQedEzHSfDZEKdRrTX85W4Uve++pkyyoSHBofZ
bSpmzEKmu6ffydMU/I1RK3KjbGJ80oYEJ08z3E6gQ+yVg1U+L2qAj0Robv9zyofy
SJKwUloq0Q2YlauPXARNDRDmzBR8yc7g++OR3ayTR/wMC84M4jdDEpOD/2qEKMPw
tloVdAp1SkM4wmzStp8nnw6+8AD7h/skav0rAhBVaIA3RVeRPHCIbbqwAES5IH4b
D3pMLPd6NUW1w+fxUU369cyVeJCtSnxL2NcKNm3kMIJrMrFJI1c0x53hQT4R7xmf
1WOyvoBH5VxI7j4KhAJmf3acn8Kw63gXde+PbGFhAr3nugV/y/4zZKCzAc5p5uj0
Ee0wdBzCA1MIt27njR0nviHSlsq9EjEYtXGIuZNTOYjgxrx/D3XdcyZlG7fCH6ad
vDImAsskZcFwUBDmN1pgi+xao/aDK6/I4L7l/G1/it5OyY3+Vq9l5PQoLXOxxKtW
OHCTSjDZ8VmYKY3X1WyKn/lStN37Z7EN40yA+EnYxcuPJorklPJqxbRcEACIQRrR
EA6q3t5DRyaT8/MZjOhW3Nz38IX7vGTrmvoCMPGbF8DwLfn6XNlq8Ep7x3GOvcOJ
mpsUTIUxDLjUFp+mRU/2nGToY3GzK6Xawsc3akxw0LofAWQ3JAnztoZqDewI1yYh
DGbqeacpDtOGAsR99fCpHrAiKubph4/tA8IiPna1lS2Evi3eVQItMEACflSJpsf1
GBlKfbuZ91t3lgT0mRgWaQaRo3YKGeMHlCGnaCFupyqovpusbMEeLjNCol+7BRzq
5C8OexthpF0XMHvReKrJg2MSiGDsuhoFgigZSLLM5g3jWsgpl+ydxNl8jJW+3TAl
MFizy4y/38rPfKWvKXrfLkSQMP7KRuUPCXKs2iVkekNtCddM7OMgdXLBNpg9G/2L
Rr72IoX89v2IG8JaDDjr9zmClXJvhb+AGQPpKmj5NGpQ2sKIg4tuUr0KHT/a88vc
pTCh4B99puM/wSPHaEbSAgr3iJpJmmK+X8S+G7bdODcWEiFvbWVdhbioO/45vIk2
xUTCINHruqvsdTnFzI8Itoy9VtMlIE+XQDLmzw3oxbFzJBb7rrVw498Nb7ijnJoy
K9UKQAY8Mdu86dI4R2b/vgLH88NytjVgb948TBymLTk2h7GrXzpEWg9P16Wx5cj/
5oPzr3fiUkEl7NmT1nYUf0LxhxDbpW0U/XIdoJ6Kb0dAuQX5jcyCT9rUdpqbz1F7
iZRxkc+qfH1KZdZQqpAms2QozUWC+UvLib5wOj82GP7fF0qj12b9JK7ND/Kqsqxt
WiXpIKYKNLB0UdKBuGrU0yEEKBHJRVRpTZYb39TAumeMYlnOY6f3vYnPHLal6ISZ
AYf7uavoMgTxnCDPeYdwAxSHjxewMpLVM9RUeGwkyOD3DIryxAjZCHESSo6fckjd
m8J5Vni68rsWmXyT5zVsJIOsuuaegd0Rc9fwtZyJxz2SMAJdE4FF0GNVX4kmCXhx
ND1a8Q8smOPB2sdBNR0KGCcY3pGilo8myj5I/QKW532/8/w73CDc7ftEMy/9WIfc
C12baHOErwrvIu2YWG5c8d5Vry+ngcXiMeV34G0EzamPGLkDdegZ3SuG/HaNOKSE
3K2l/uCH/btZMzFE7Fzid6OyRkO2jSYuvu3pCGTcUW21iyBZnFqEt5bN/Z3Zu177
NI0H+LImNQL89wjwYoSB6UoWNrBvoajEQrxu+Kpwzcp/KLG0WXDJlRcszu+HRD2t
4bxZN4g/oo1rMg0nAW1DynPO8pcLQdAJRV2XLVyMelvw0lR8seLo6DYZP43je5IX
ujH7G6Oc2kv1ccrxcJWHrzp6Y2ozlB9+2UI50y5jV9SP9qx4/wmFx3L5H0SrXQ5E
VufAHurmx3ZVpma+R9KCS9k4fBRR2u8cd9GaLuG3pr2vVrc2TqV+zD0JuRydmKht
KTjWF7Ku99fL5gIMI6s5A0jyvV/YBNJCoF7V+0AB+cLrQzlx9/5K8YOTp2N+1O+y
68phFuQ0wlJ1pp8j7atTZfsKKab9kkpxvRYoahTI0QEgFEV+qiJylgW0yvwtSGXQ
eLz+Il2eub3OYzF7N6KGi/ktojFjXErZknHRHbbho+hV7We3GGXlEBsf8L++GGNS
yx2ieXEVoLnQK/pu0pEF61pI9JnCeaWORsiil6vhK7OhWmsaKPHiloRhJC4srO8/
hT77DkVRM146FFwtTe1CeeNjo0AfCIGDJg7rpl7xRG9dazHBmPGQzRd/heMWxDex
gXV801o3xwaWIjw1pS8580ziXvSP2N4D189qycC8pd8MmQRQzo/E6Jk3BDiq6PRV
a1x990PyZlK1KLU2iXQ8piL1V37xmVbCQ8BHp6MUG+UTk/qTzdb0C7n2/flHbL6e
D7YVnBMzPra1QIpOmncdq7Afl7iwT+JC7IV0VTA9bR3oUwhbgxDSiFq2zbDHYFh+
MaA4aZ2e6XFfMTAWrLi5QG3Oglra4lyinupBl78a/06GbH/GmkaUjen1WuNhkOgY
DpYQYBuQLFlLn1j7V9ccE7Yzyg2NER7Rm20SID7pysGeZwIQRITZ4nzQjz7Mek7I
EN7Q4czChpB6MP+jkCriWh4ONLRDj4j3XVf7PaCbvqUDsHA3vD33hLbk5xz4YkyS
Bj3hCUSfNfMDJ+z5QwOzhLj5vLWyPj7HbxHE0d7wNY1rm81RRpXD2+o2HHB6PNwt
HRXyMDP4QWDGJIxityo3usPmS4boXgjk+qhUD4TkuEW4fvfJ5Nd71iEe6tVH9i5l
aE6/ZeklGWFuTaZtJ2T/c86XQm2RQ5QoJgXvMmpCRFK2gTnrXGSOA6m1ZrH6Cyk+
5AZHIk7z3tPAO55lzOoCYBlXjuEY4eLHErCdHo56104aJcRGdxAFvfkTyC0PoT5o
a2I2XDgWKqfjom+2tjCOvCwOKoX/aTUb8Qyx4TG8IvTRBdYDqoZHix1xqh6v2W88
41rXAZ2tsa+VN+ocySqJU04ckmB0AdtDv/VZnEhffg1V5fIRcFXXEuGx7xZYXjxF
j03Cl3MUf5hK+2YJIbp0tGkVC0brDSrlduKvbQKkqs5PqaPngRuLSf0Z8TS7xfvy
1ib0JJOG4BIu646OHFjHW+s2+EPg4KaS0S8RmVJGBIgYDOU2NoGpdwNBHCf8jY52
qNYLB29wcwy9LMIQAn2D3KhLwPqqRS9jGu/IeYgcuWGIuEPICDqkZNf8fFNnPlHF
r2uIFaLaa98RZdAKcfvTcNBJkpMOVRlMU7yzVALG1gd33Y+TCI7O/jeEf9tDmT2a
OQEU3bBI0YCvArsNIbo4o2pNDC4g4NN3yg2yqc0IuuFdY8lsolupEvKJvEC7791X
Zea9ste3D+V3nQawtFB4DNw5shW1SDlmF8/MLCkAfcXZGKuy9GjxtOmdTHRiB8+C
kDe1Kegxox1Miq/gi91T8KBo+G9XWaiLrn4+7FWl0ENBmts8241C+CXrQcaFp8eX
TIE89sVXOHhMRclmT6DikCVYB2G/HYNi38jF3ZK+znKol/pl7nk2WtfsyGCKmoey
SJFCTaPyW1B+Oa+yaqzLGYEy79R+a37entrGpxz6wA6EQPtgSub2vtE3tQb0Ekze
QYm53tqWbdsPOoBjJnA3ZAZspjAJLEqcwfwdXg+XZqB41BZeOdGtzeMKutAF9Zus
4vOmM9GtlZY95+X6at0yhz4uXVkyzlSh75F/6AzJacgfKrwKBltGeteSAi7wA2Z5
3cJbHg8ZxzeyXxs3nXQEXB8iIbYGmIoJfMdKV0MXz9t9Qmjwz8YxjlxhMuzj8Su9
ZKLqlXKTIZn3f6N3sxu1WtIJMqBE6nlD/wF6wywGFwI7zI6l8j7iaKkkbFVpJyOc
jwGDMC7QYAezhgyVfIjaRIV079VsoqHuHHRM4diuIjxaZORlPOW8/AHuOh3HWiz9
GqH/6Hz11ZkqYw4eFoBrm+oknXj7zMKG/Zjo9eO+QTs9Sfz/nc9kNaWZvDlngUwM
pjvFfzBIx1X35V+IWBtA/1d7pkFc/cxWjQLXLs1zjnWvAu1re/PsRwB3F5MLws8v
nxGQIYRHlYCppLLOtL7eBIvTSV9vReNca8l/8YvfxUMHYSoAJxDdPy46G3p4cNqU
RUv8t4DRkPU1J595faqTzGXEy3B3jXnUzqdFd8tglTqUy2kuVAsTkoKsH/D+BB/y
b5mVMyydza76n5Be4qPbUV2nbAxDZE/DrWNmCPVYbRFiHaMK61WruzUsFftEZZ3P
Zp1ypqgvvuNk9TvJbpM2lc3EoocJUAMo+Y4Szf2pAk30zFKUl/9j/NCUr8nB022U
6UdlSdV5SYNH1EwqoMiIBW1V0oZ/8RbyRmb9bqa6Zw/QcaXo1PJkPh+uW2fzeSff
0cGadDt3LgSVpPkUj0CRfMWao/AurLFeChT+3Hd/Wqe6uV5PtStduGI8rXB3ClqF
9tTwFKPUrh65pdOIdvMTKmQQux4HLa6NP2LpEwZO27z5Bco4DfHZwUkjO2v64iwA
ZdaI0mE7byEYIiEeG0GI8X8pDMd2wvppbZ4w02/UieynUuVHI/HENoi4L38T4ZZ8
J8dJUrOvqoW+cN0LheCliwZ7mM+EWjrSLLWZjtZEwwjPxYS9rQkTANIh8ERRuC5L
tsBE9j0WM4EczOi3t9n7JYHWu6sU5I6Z1IhX1odNmhole7FwZoPLLwRXYBUipHBZ
1PWDTADRt/xD203YBJ3RMppQVAaAz1sPuYNBwDHFPiyqESVQnaq8Xt6ANgyb3gaN
QychdWDx9fRJmEb2aGUmNJcUhoxDrGms6LfuLPWCYeBjAdZZxUJkgxNivhyAfEnm
1KHjbt3G1E/ka0mevRYF884XMj8IXNCtgWHeEcwhQl4ULz5Hn3SF6xbJnkqVSFtr
wqwuWu35vHGQivU6l1Mwn7Dc+SOv8AN+08peU84RnkOdKOEkJ9vKAwvwUtQnP8OO
4mlrVbCyLeSnQ9EO7XIZF+teX5vmaAxSyD5bkO52qMzB23RLciXM8fGrujhnz4cu
NzFy7MZIwE1OgB+4zJlcn94A6mbbkakRt9oK3O1C3uQrnOSwYH4QeMzxYy798rOk
yslbAFAJyf02pn9KoM5Dm0IvTq4Pu+J24jdIEZ1t0iBXg/NlmHqL9xB274VDSiuK
GAn/NSAQr+NrcsIaalB0nlXcpkSnmqg6vUqVDdohUMkezXfStknz182vfmHC4Dak
RDPwhR0QlRhBEUsdfcvzW/VVfTu3Lcih7USDJHOruMwf56eUa9AocgvSLtGVT1Do
NVX99QOEGlcl5q4enx6I09wQ/Z1se6f2TmtWzh9yUeyNlCX67j+6mGrBIm+m1NnC
vWbV+EiZdDrO3IZz+D7d2RwbcpoG/ycdLsAAx9lev5fvr3YnUOEYJQAGLV9/MxJP
MBeKLC9nVjRMxiPBENtwuKy/YqJn5u2if0VmAafbwoUFxxqz4zNd+mBxArSdl4C8
WTmogSghQAD01CXNC6Us4d2Tb+muD9AO/K75X0UmTA3uQS4vpsv1VQuAGCMMAjW6
GtKgRG+KGcsOFEtD7FMn14DC0I8RalUihRnv7U3MdF9x2BrAvUUbeMYgdNjMRrFO
rYSbLwOfYzm7FzqpsBjniVV0F65FvkSfCX2EAIagF3gTb0DZexEULOzTybKh4ekB
ZLAoHGFJtHSrbcMjyjLXlz5vSNmcAUnyQ2U2Q0KZICn/galySkMy7DSO58w3SVeg
czENpOFSGkwc5BOKS1s+4datVE9Bff7aFFZi73VTLrAICePnO86pJKJTo6VatHV6
HBx3/d/PiZkMe+ur2o/gITXwEXicNdZjqD/8UNJJxZPqaDKJ5a31clcRv5PpGn20
ngjlNPdTMLxgeFHxcGxjhLnkD6OrVJnEWboME2XOn+FJfOERYJ1zJIRbSiqB3fdf
RA8cdK178FyAmL1rf/nXgs84mE+Z0p/RSDlR7hB9oQonbpnuV4hvQTyZR8hiKC95
6i517sXkYC98y28U4/VpznUraMraZq3W4ov06xofdCDtkmxGfZt6Vq0NXCYJnEee
PpUdP2qGA5T7YH93zuW9V4LNM3ueathDMvP0gLGFLDeUnzbT3XhUVFCd8JuUCkN2
ANpYkhWSgmDUfGSrTffY4uHdFzuIsgI6k4INt2cGY/5mDXjfUCO637YE7abWuUOf
MnGPTYxgDM9ViSegysoqGf0WdwI0Zwq6NoiHW2R7eGe2Fd5TMBw3uFZFmdJ27yad
CQAYaVDcDnSjynUKK466fxTAJWgfxypfqcyz46AjgaE+dfadGF4MQL4aUjgaR+L8
lP50/yJvhChnn94kyxV/8w7UyJ+y/oAdQZUPCtiiG3x4X2jPvUfcP5WiF4jBxfHx
bKSHx7dQ/yGQrYX+SRJ1YY0QjdJyrh+2kZTnnDAhYX3TIsiYSzR/vtKTlc9KnLsJ
H+uEQl4BMsnOgwfFIXduDvnSn101K5+6bYKlGeBxgRGe5Wmql9Fx1GwRsRL9YFYI
RYpOOBLJE6O39QtjJqNCuWiW/QATmKO0YbK34yiY9hCkIEOomOUHVIj3/jf/S4Je
p+pHBWVjiggbN2Mdq2B1nZHCmg7v7h/gQSER7NChwGZa73Xp911RcKs3Tmxl6Tgd
UaAjVU84wkCpvYMTjwsz3cdLvEPUivezBZ5yyM1Wm+YhOnjYHRqcRW2E+xTb62Yy
ivKKhoTK8DU0lSEgNGvIqTrLCJzbA0Jb2/FrJK9rwiWk56P7WCD24zODdsUiYSZL
CxT8QJKMlG1jusoHSyBm7oA7J3HkvXpLygd6lk7sovjtocBVce1MOrcCpFuqMSwp
0WcbXnYRLmrpUJO41I9kehVLNwwFrRR/I0Q4aB8Se3vEWN1JuCcVbgFt8T+X7Fg8
IAOxXKF1BfA0zni8h1Lce2balumFFGkvlG87U/RkEMCEV3UeqZQrSzi6qGwnT3sf
ZyR+Uze76KCOWVS4Hdr+AiH8DS7C7qyobjyGqH9wo9+FeU0wa0xuTySoxURWik9C
kg31BKMgpSbWaA6BFIaHkLxv5U2ehOf/3rZoLVIp85wb2USzXuTHaI2uc+y8qMgi
ft0APddkgDANfdXIw2ajfnZrlIN2NTVe6gyF3L8SYzfNfEC5vgCmX0BIjWXutJ1m
V+UFaXnqz8nZ+lR8yX7hKhNBGJ4X5xo6goQoqqPvpNUAC8a4LWnInoI3khEM5YVb
zWp1ockZfCYezejuO1Jq7+/G/SXZCKpjm8ZzYGBXkQ6Sn1Ez8ojY9KY5kxwiXoVj
Wbb87kVUONHdb6eVe7SFqcklfjY71sLHdajjT14bBantFi/eoC09js60y+XmX3a5
2PKpqEYBTBw4AwiL5qf1V4ek07zrnjKTUnlM8DOTO3LxWB4ZLFZtl6LiXz4uzx7D
blNkD6xg2PkajpHLf6TgFl+FpftJZUboImmWzTDbWHu1K0SiBYbzRFpVvqv9pJiA
KYnnClhnsVAnAy59UOoHAe3N0SbyHADvIOi4ZUBYGZ5RuR0GEd1NkoPTRftlOIMx
NpCx6mc4VPyFtG0E7PXvgTbPfYDSt4txXDrvVx0guegvgZ90mRFfLlB5LijFKe2T
k9Dt68oxY/Qf/JgDqn3jwcCpe8bljGhvg+HqDw79/T5rfV7kJmnmOFdf5o+X7e92
kEPxob7n8iqhqlzsaLaYWsSqZQw6rtKwjeeM0gN5Z/YdvwRRUf6Q2p2d+u78TBDh
2qtSrvfYpPT5r1bob3OQduKluGwQHngHzoW3oGKQYD3iKCU9IQsqVratPIzZama1
pTbjh1tqLRqLVt24f2RZC5DpQO7NBUyMWJt2fPoQHeqZqwgTdebjZp+wA0BzTgM6
PSIQFp0pW3Gjty7ggii9i/SrY5+woUfu3UFAZroy1kmFB+ZrcCev9bwQ4sM26Tha
U0M/AqPzsl0bCDUVEm95FYPsy9jWNbDUWFl4u9TV+nQy4OB6NFNeDZ+vUEL3gD0z
uh9RERC5aY94sXeWi7R/1dGWLmDr0HHJSI/Zq3lPfsrB0T/tI9yXGAthsqR9zWpS
/xE+KURciJGwQTT1katdKC/VTiTV/rmeu87EHUJszChS0q7bWAlH9umft4oxRUF9
9YYrpwUdJKvH4eiDs5yON7hFP8ITum1dlB8MoFaGz3jDU8CGUoTwDaeQOtlI+0pD
CM4wq6mvhW7w7vkUTALBNBciAT7Q9mt3VDT7adfTYJMLwAxJ05IMrgsJtTOPA9KP
xeesQHYRBcoLuobotYRj1JzD7CnRjbGn4Xi3WMon/7xuuOkb/+dHb2W0+h4nft/4
ZXHmMVr1P8kbmlU5qKOmlhqUocKchi9mXjtXlyIt2Eyt0h1rZjPtM8EJ5A+jBCiY
aeKj81/TCKeATGZoIRtIU4sAzfar/McshT63Wc1+xh8Qm4/f7FwWyirEnA7iruPk
FIAv7XUnFYDkwopEov+V79nosYipoH3qOW1aPgTUergvk6lZa/E7N4SP8SdbfP8j
z3IgDOUR2A+sOu0zIXF4iyAF1ZpiyqM5IWZbdvgq1n19t7n1OBTDrx9+0L+Ber8s
7Bwd36SkqxhkePNc7EECkIXlNx0HCg4LiiidVTFurhHHqd4Bau0p8hRPyOLJuGKJ
QC1aF0erVfq2cxYni++gsoF3qyX3Rw1I4dxOQhWw/iZ5xbdOyeMQRKUsr/s1WFh1
A1ed+JHfP1GzDKWkuF4Lle5uDhrJmn/WIb/cAXu8W2bVr/MyfEKViwDfFm4RzfHD
mbzw5wVBXgem/lfLSac/4ckDslPjto9sHqLxI5Q9wXG1tVYoQBF150UpcUX7Ls/i
6Vi/iSDCwZwnrd1q1tvqpE4764ArxBZJXi+UxSh+H1ZW+pMAqza0nPaDkrVchzT7
0aJhRDdHwsAugFikeOnzlmNKHe1+uNYRJiKga+z4e7Lo0uoZpZXlQd9xcBSmD7AJ
K/TLRyN+YybU/zC+i/ml1Xthse7PxvIHeoFG1t3bMZrdk/BBSPqXKrDZw+D2WO0y
BaHSN+uEAzYeKosmtmpnS44wdT8reGcBmFtIvsELlo0DYbljM3Pc6/6p8o5i2q1V
crV/XL9gRRvOZKqPk+axm/6nap7X6v8YJsVA7gSNJUofsgbBAbZpuOSvnJGsHN4k
trCrEBcpq0Z1FNMYXkQluBcpST27gZpXZjKWKQx82y0Th4Sja9OXNdUqaWqQSIZ+
sC+Oto11IbBVIaFPrdEGVbYaJc6DAD8kS+I0pJaNY26UiF7aOFmLchGvHpmuOgTh
CfyqNs1FcUeqY3oCdbpYOiRm/abrktoN0wXv/pVtcMyFn/FIUHNzpqV5UDaCpSTZ
PDmbcTBujGxuk8iwlyUUMNvW1YxGfvzufJ61pH4O2s+xSnL/VUp8KBZdDUDAfuyo
+8RSDsvNhLw5wG+nYjPGcg+asb5vfvNk2hvSuHlJQf0MT9bhhPlE4AwdohA6HXPa
R19vrYZygX30M3QKillFvRaASQkSRM7J8WuO8uc5HqYOcaHA+D8MSTLs5SvS9Cea
4sHg1+nyAmzzTlLCAPJmO06yO+kYKRB46+fMJFjxKokYGfR5Hk/F9tkpTd4sJtkE
06F+oAAi8Lr55w/puVemGe5Mq7pnDT2YEVL86LsS+0GA3T93KhnexF8PVUVByGtw
L5C32HNRhzxeyTvRaOyEuMTAk3sn51HlvijvjLO+KgNkkD1oVGiuds/BcsNd/oiw
1sy9Fjq/vmxVLkq+tJcemWsEZ+FbGKM+5xjADlhu9zNJjdLhI3Aa/Q3LUFLlevHV
UK/R3PSXNCneUGQqOaLHbvOSJKuc6swDJ5OG8mk3tc/Fy58SQjuQQsgEDP34VduY
HZQ4KNZEhtEkzDmuRLD3J5Rw7Pq/qCkPCx2ica4odGAs3EcieCVOrfEZAMlH3q5L
Xw26utYBdMFApBSjgSvgOK+KoQzGOVPw1YSA+AgQLTMZ5SB3gGVw+jOYtGxYTdcr
ABz293NHRVQSiewi+lVwNcTFpMawqI6ma+xrrVUZzak/gAJ6k0N1LdK63FWzinqn
/wcIRy8JDAmzKHcxxByb3MnYE1jxdtL+sK7ysafM9dmrnX1M3bYSeh/rlGewo0tr
c/fGW4QIlpdqVJm4SYi2ICCuVJHly2WHsAq8kHnAYpCZQFs4aJYuVor/t0kBin2X
mRyY7bQ7kt7jPYEEIRgSVN9W4gufmrLztQ9vwGnv21+yecGQX1FsQ85zRYO8k9on
ruuaZcwSibraU+GTS5FXC/jhqMHzoLaomFfEoD0q48bMOk/bclTE1UzdHmawspwB
PSwPFv/TePuTIXhD5mz1HZW4dazjP1gCQX3AkuuuDU0xMvfYgc08gxpQgUp2SWuj
x+oHVpECRK/5KIHUFnRmYZCfaaYYkVOMzv5satiO9rciKCEV+97bktZQevSroi4b
6CUqH/CVb9ni3vSGzimklc5bSfLKpKumgiGth1sP6A/xCeCoEKf6uI6fQCGLyQ63
LsCXk3guEsv9nCO5E671RnAXkmKHOgarib1d73K2FASaZkvpONLZezFjTLeNBSWT
+9APQAqu0dw3Fbce4rEsmx1tt3MB6rHhNV9aO+2RbgYK3uiKJ9uX7ItwdI225TBF
aJ2oDmoGbv9IteSDqr3Wubmiu3xRpD4/Bva+v/HsVCcYiNDZdU/wjZhcWyMlYUXw
E3pPuf2Xkbk99PelfKjlyLZS50j9GePrtBkJ9qZGSLvrKRz77N7Ax76usAyX2Prx
R7tzwjr0+AbrBcDKdfz2OwdAgVQwd4u/va5flIKZdKmyZmnaL32iL4QL+d+9lr9n
tMRWdAD/HKOZAz9fQBDJqWkbqAdNd+HvJTE4KceHjyqkaGBuTzOnHI/PocUQKfEa
rW7fWXj0JYrZ/bBAuk2dwnmgxeG672qBYya6vaotxEYijKOKO/1sA76tpsWYv/BC
ZIbckWgXqn4upJ4vdYpMQReJYQyqsfqAYLUlR0nVCh3LM0h9lSDoYsm7GNJXF8Ai
b0fQe/hlrQVW5ZIldIaU/7TStlDvErN6WQc/S+MzKf55U8J+99NJb3I356MYN3mP
QbLlL/scW4KjGlHfof5aQKPajyM2P9eVKUjXzF4j6lY/BBSXIxOzpUe0CF3HNBHV
8LUV9go8hB9a4ubiGCAhPhRM5V2g/KKx+x4gADXeBOpfjHu4orAYquT212QrEZ1p
S0uEJoNwh32HH55G6xhYgV4yzQC5cEKee3XrdikP7/+H6s+HmPHqnk4JSFdBZ2bV
l2ER3z/2rMoiH6icBWx1MxX2uSxB5dwY5oJsL4O8pYArxCMUEl4AI9AfwlckGLei
0fEHbKiglFDloz56AoK2OSzZbZcqsrhqfJKP2uFo7npO9BRK6KORUS7UfWJ3zrR9
hpUfQ/r0dFW1+ww+etnyZixYgtxQn2q1ICx2xvUGd26hNJq+kSehayMvX80YCmqX
XkqCi0oeo5XgX2DT7diwAqPjyRfaEC4SFcbIGCWLQ+4/BF4Xoh5MWnAQXs1k+eKm
q2w8VWzxm0M8C06Cw983+HImzz9QgieiZPFNK/LJqR4WCGToe+QRZZ5etY03v+5I
5tF9CGCJ/rEDcPNzGRVmuHwfCl2vP5ZYc2DRdJpBB4peotF6O6j4q6oeKZixcUTO
ZX61ddfuZNQ0TxDhv2Fa8vDZG+5/x1pDtNy02WFQH6vfLJg355eEm8XGWQ3fwys3
6X3HW7ryJ9C9PKcwj/9fUvLxZK93yeS21Zdjas/RijIUSHQAmxCHbf9O2RyYqRTE
vUvpf9iCFMl72yi8T7FwXRB7Xt4MJ8kXTk5wnfg8s/5ivN5SOW5gZHNowfXEOCVo
Wh6rjWsXHmY0JM451wbIrb6paMOFF9h1U1B0pc8yOENu34k2uWIqCJ6ceMD+iuDA
IHw1tKkdkRq6kk0nb9YseFr+Y4I/vHWjnSUbX+sOCzMurw1tU84yxjfDB7z4yMVS
FR5PFbEgm0UoGkY5Ds0U3tW7phVYBEnHOj90YVSeuSHDdwPWGsGE7fxmQPniEbu1
iJfbMEngTTB7NYjQL6Rnr/Xa5IdDiCNOnGg1YB7AKL+fywrvpEtlE9QFO1KElcfU
Gh+IXliK7vgbsawQ1YDxXh+vU/NW7aScqgloKY/BuNPA5YHOUrTq9UgYVJrwTC8O
XDy8XCUpG2ED597jCM17ij2uPgCI9XtyB+RCwRO7wAGQUl0rguI23pO6laU9As6P
zDurvQLVaYN7ZzyrKbDiZmJZPORdSa2YDdk7/kZyTXXMoDg6I43vUiiEk/HqUD8B
0641cpKomrFtTag03YC5iMw3N6aotaLaeYdqeZLbbSkoj83s/MKwVEiby74OsrIk
Z8AeoVylLtYrIw0Q7HFZt8AQdHB2ZeWOf7YdWgAHxqlY+/5DxeNcr89PjFt9cvDb
NLp2XjthPUY3NSHT7SRvYlAXy9GA1PLgOpe+dD+7HVBTXE5/vcL1fJzV0WzG8yc6
3EH8hku8qotmDFraEGwTKmYVFMrwnLSCFUR1+LbJa7toa2SUDv3R4Jzl7brjCBqm
XLv7V2owqqcxVWxlJg/JbsAuS+nFshh72rQr8JQvi1xyTCkZJc7pOihtK4M7x0xL
bypXXNq7Wd3Kp9aMCOEpXodf5RQeaxx8Hn0eIU1B2A/DkfuunhJ0vbYyYmf3UAXD
ZWipPU8+gDqvy1soLKhroOyX6Dxshm3wampxHkBe9pZ0xYnsEcDjk9A3z/TLUb7S
hDBvMjvxWQx/cGxR6fHZok7JAuYXD8WDXEWDDS4Cx4ELWlM3Iokcxryp4OCSlbUp
+tnNx3wsceppeP4MnvzkWCfj+VYzdw/XGA8bVNaGLGVLXOlb14ZbxGrPWh29posm
J5LPCDP6lg434JJGPUB+UkkFeY4nLwxHGOeZyq9gG5Yryn3+FR1S/43C/ggIUgvj
3eM0wRug/Qjtce37onGZXSsTm0hvX+xilPpdrMSecFJZxhQL35c1qbhLgx1ymUxx
9l1p0QiHMDzK/6q3bR1F52LBTw9DUTDGrVMjdKdYsRsoC/AXZ6tafNrUrl1zdE2m
I8b2PMvjm9gtSAItgrgbrCZw6JUxDPazKqCyJVnMidRFkLCFNe/3oVPPZEBTdimm
cBaVwZ0yxpsaWkUotOxmQdNbVw4I+GEewh/c6CRHNu0X19rE0sDEXtD2SJThdd8F
GDEQSfeybb07fNqohehgT/kviH/qeNta630hevmJ14kifCt1O9U25mWRcKZIYjE0
rEsSo7Fi4Y+Xwnlizni3/Zq8Xdk+urPKAjYMvFvCt1u4CfUCcxpDY/kPFu0x3nHt
35imDp05DevZBIP30Tfxt2x9LG/hZ/KM0/lqXY/u/HEnW+iShmqCcE0P2ETvgWzi
a7wMnMxm90crCZODGg/BZG/FwJ0ZnAJfbiEcZ6HOotOG5fNkSF9nHw2+TbH4o4Rj
s13+1CcagDEN08k7yE0PktLSR/8QmGwvHeVGx4NN4iL7TGEBvumNxfWB6tytqRdI
v+KSb7GJUkieHbaZv5ehH3QB7FZbjY64FAuNn1mD5v8dyRdPyThBMDrz6c0Cz+wj
re3CFjYkWGc5gbW9rsQ9f+9EjJgZWKDC8C1R2qF3tOVpLAiFELyS1cZD5rZjtENX
IrLsmt2R4kIslYHVJ73gEsOU9X0uxJm0q/2GEWXnALmTTU1iU/98Ui505QI6kcni
UfkkHssCq3AbaE5jGpruplxRn5akRlXIDz4HZ4CsU3D1XJFD9qBxQH1g9i5NYe2o
x64WATAWGsGN8/hOyKUNY2jYVjIQmrkdD7Aw/fqTAZ+J/jrhFynjA/nFYWe0mKZP
cs2zQbrKhWYw0uf46um2iFGdiJAu+DowaCtdw9OWVTjVkG42ByDf4M7mcDj3iSae
x5J+1uvyj5CNSHYWnsi/k1GiemwJ1pcrGXDNtRn7jDOByZz3i0E5YgilSqEvufqa
PdsinxNa/rjrB0vG3f7/1yclmMjSfdn0rMA1FRNgNBEYaw0klgD5gucUhyzOrHb1
VmlVtKyNaXv7HUjny8QCE+gyn9dbNd3xm71bo9P1PPDC21Zk2nFjFH6sUmDjIuJG
DYxZzY4etJ0oF9PhQ+QzhL7hb+YiKc80rNRsAqkYxkDDvWQ4YF4rpV6/GqQUDIsY
aSYa3uWrJRXoTzEA2v4cTOvStTchJwrlYTWcv8Qk2THBzi7D1t3lLpRECN/ptSWf
ymeGokbW1YyWg4da+ijzLotsFh8g0BMzCBafSZMU+kxMnKTJ54rZXd4spDaQf6ws
CMZmSitA1xHqd6+pYATadHMXxPmWhHX1VhwnaVrAWVI875wjTYxeBYGnFcnqI4K8
vzotj8ZRoG+sVFb0GHPtBoxnWkmFfoadOjKmW45MGO64/7VSJwBWCA7aAAKgcrBv
wgOWHBR+C1gL7X6Z+Hp5vEpCkuknsEhesjrCrOL4hW6JpgqR0PBzwZLWAePkympw
AimX51EqLwG5YNL65JDZr5WNgetchy1CbCEBLN8z5yf3Tf0/v8k6kjhLinj0PO+K
s9Iwc+Gs79V7Lk8E1YtygXNFdsij81fWSzoWVDSsGA+tnQWmnaTS4BIUGKjfukxZ
+tK3C40UI3vv8blvXtUU+fwZK0kPZaCqPYbbS9GntaSEIGK/m2hFnEMU4O174inx
9DYR2zdugM4UF9YRl0JACSE+/UWL6nTy+y3lDTavgEibq/iVw8UpwdC9K95O4+UG
GWTtfY6EP4/O9NqXUNzZHJgK/TaoyOfLvkO9jXBcvfBnyE13UrgXnU7eDg8q7Jfp
5v55XVMlVkHOBGxZymOUCAQGjJwZPqTFZsWzwXpYt6001GDZ4vTOU7+6rD/OHflu
+7IJ/ErCHTwbr6TTuPxkJZN6w7G3+1CCKdL8BkYs4eDenYzXyXUBjjKRvxfpsN8i
Qx5jRIubAudOlzyy3mquE/hQcLoZn2ixRWnmFaOn17MBhPCRoM8vsAqibhbCIQtm
1Bl/d/EpsIc8qFBqhcLQorNFlDBkb61tCjUDu+ZbThZlcyJENxZ/83hrWwXpiXpF
50/fK3A0KD6rtYqQSFhXdaFrMpfLccyNSD7u4A+M4gN2G+LVzXW0j5PcN/XvvijF
T/IwbIzi3ImBQPa6DpXjGWe9yr7FpXV6lq1Oh/2zU9gsLSM/yiKwXNDIebwIOgL2
hFnd+/qKmhNHWqKMSCcurasY0l/x8IFS9ykGrFc3CiuLs6jCelhzccXDBxPYKT1T
OoOhKgUNluLk1eOUDcmn0W7fMoL284vQGDr5tkzwpcBADA8g6yPQ34ZJLHUyIW4i
o6GTxjemO4fRMGedu1m3C4uPmYKm9uX7lnUxMTIdrYNHFpypnJ3SK7kHjuvldotn
xm1m2QKx1ZMbj58Q36MiVgALLMoOjW5LbdzRQTcR7FfyekhFcVa9T1NEXAmRXirk
9ZdoAAN85kSkt2+Ycoyg9BPEB3eiVzCLPrtHkm3YZBD7G7igK7j1sTld4p1nRHFF
oMwah5yzMurEJoVEck/8SyYgo/Urhu8HEnmVcr+q0V5KB+oEYpzoB8ovVV4e7bew
aVAwLhxEIv70yy3OnmuMYE+L/enXzooKH+yPF/AbRRqK5gSnSUjtjbDkzFgfKvio
JLem66Enu3lf8KENolph2O54RNFxQ5Y1Zko4UW4EHbtsFnsaKDSI1bOjqgHAr5hS
lGBLGuieE22Hp8yMRuGE/1UROjEUER2e/owLA170cRMIjrQNSu0TjeyjzwKWUSkr
1QqCqPcA0B4faj9hRZSyb4Efj34xlfojR31hE/jpSIhjlHkc3jCc3uXDtZcDk0EN
QHfnYVV+4N4wqcUUMBBC7Rb+W8PYxECXv7A/tm8bCyuk6CNlJ3wo7TDh7z6yxS2r
hkk/u8xPZ2Ku8QBLSUqD6/d0/+fOwcMF08zSMBY1IQTBz8L/p15bwzqdB2PXM98T
Kw7ChamOL6kEcM8v/y1LcDJ+7g13+cYpT/7oXLSboQcbPpWigD9CZxs1YCDyxtf2
CFSWCEzd/eWFdrxEOe9wiDVrRXpZ/L46Pce4sKEo0tw7pvUokfE3w/DlFbwBVwW2
77ir7izzo/ku6vS2IYPd7xD8q68k0CHkEwd2keQvB5Wro45sKhD//Cvily3VMUaV
XuNr5pof80wdds0R/+gc+n9dp3f+pGrCsPVPdVVWJhH3XubMqtfC3/x03XIFE8gY
xRhwB/xKZNL9a8/F4Jc1RlLMZogbUFAKan2aqlbUGFrySlBArS4GC1sA3/H9DUcU
gohrrJ5bNBiJ+vQ2RBlnmkT0x14UcycPzojw2iNdrfXIhae0FScnpm1kQZd+CMHS
aD0r/w7Ztiv9c8b4RTN0izuF+GPanBPKPKKlqoRHG175ycW3mbB2cvvlk3599pvM
RK1GVAItFxjJfsDefijUhdQ1p8oJwTCkKiF1D2C8l92dxLObLi0/q30cRoPSnqaC
vIXA7bqXto/RBXqrBNenmjCkov6yf7qbhe3b9BdLpURIBi+Fg4DG2GUelj7gH5kv
flNkY2XQB8L5ARIGOz9sX9prYjQWBncKjcW+9oD82WdxvnzKiWT9+uV6SQkQDhEK
LfjrmyaZmenhasKMf63JxgaBAytBAjIzyH3QR915sUeOM0wh15C5Z9+cFNZSibvP
26+XdOCKMSKxsdMu+VGMBOZUbaW0OhcCBV7gKjlfjPaGWIWGh1lFBFD2LRH24kGg
3LNTFLcdqOT0OAHa75fO/xQEc5hZg9I7ATBdWrPEMFtvV/VInMcabMmhr6pFCLD9
VILnaIZr4DQvn55bOGr96L4gtqVIAJPH5M0kt/vo29KZVUMLyLre/y1m9gg0TWSc
WHqX4khBnl8pztzIuV4LVNSNyjHcUZw/YkVGL7uBQOBV9gBuWNU01V1jCla2ix9E
xY6bvoE+1v2Jmv8BC9FpWiU7/GUm9uGBSCyBUwb8QlzPGlCMMEHJXebqh2NRvYPw
XB0fObvKxPm893hu15+iwwHmTdrJjOXI3qFIc3wXjVAwvEChtY0vqjyFMlINnWT4
ZGWKPJlpZi4fz2GN2CkaEpUQ4R0T/irvZCa2gIIddSSIxXB5GGKqjsxuyugRJ1fj
Y1ftiJxTcT+jgdH8HO7C0MtbXStCMdxMgfBlHDePlLX5eZCof03Z7G8d48v6CkrU
FZFkCFMf1vo8aExczQhn4550WtH4Bjo3SNTMQxmpxFe2roefJiyJRDSCzWhSG9NW
1c3uj1BHMzzU/NDRd9dcvOaFe6lcKckJ+WDekZc2B2ZUST6p/GGlUTOFq5m1nsWV
hMw+kIgR5kdXx4ZV37F8hnFjngaSpiZDscGRoz4EYV3Vv8hE+Axp9ZwuWeg/Y1aE
/mcHR0EzobvwIp4pyvl2IAxzPBrOFRyV9klWAaArejIThBu8rB+HWwSnr1pZaD6F
FQ1ZEkTaCLCAisNi0dxbNOl+cYLlbffoCR9IvneVUBmwQWo5EUBuQ7iWUArbmx89
cWjahv8RnGM/e+DU0BKR4L2pj9W80D4x0jbW6iAjPg8Qj2gOv7GQMD+HDH0m7d4i
sjr5EOW5O5oePHarwe0vhE81IVjebX0yNcK89HGEYjbUEQnff6ENEG2BS7vP+YMe
TW68HkLXNEmrnAchpsWKPMKE1q113xyCeNZUEZ3Je39Q7s6SUrfILnKpwOff591P
jVRct7afubUGgYLs3nxYMxi4MHvvKUlhaDQdqEnZeHI7maVMQ2bpXjw/9kHx10Ib
r9IVG1QGDKNp2K9dwzqFsviD4oFDY69aKxfXQ2u3hGHyuz/2Ev2rSXX5kTXUn4cn
qk4nJxqH5rD83U5aVOPg67bvaSUbMIdJe4rP/JGwEqrOuQGEHDqv1cxOc/LxSZN3
YIUO1DE4YzNNTh6TPtyiwARj1KwnxJbCRfAPXlaKAztZgcrsIlm5x2faaCdLHnZn
l4bbqf9ffm9DsNJ7a5GyujvYYtI1mY6HZ6tlxMfuYBM+7LPgV3SNy6KlGjTAQ5vl
LJNCrQVo6IPqo3KCWK2UoNo1k7GVnMXAiWVSS/eZlwtyVTdB/DH3MmVWhoSQuA4H
Vt1JqNp9riL5v4VFxi37bbCEpxtv4A6icjsmdhIjkUgnIN2b87wvX7ay88bMnwda
nIi9H/4MVDsGjgA/1pKo1uo0jfUVfjXNOdRKc5/Y/7XsybXrMUBkybvvzId/E8fN
d0qhynLCsmDqqGeMWu0VIujPkQmfhglr7c9nKSlTpzpXdaexkbmNQ48N5YHjqPI9
ii00gnKNa1fHiss5hJqqcWMNeNCjAGA/tYQxfJ/sMEpUyof8ZOwSTVSSNIK0m2mV
MpIYjHtZ2yM2cYstb9O+7hKUM0LW0Eefe0vj9o5L6h5cEZLFbxBpLejr+bIFi5t1
YZAAYssJmXuK9A5CfUoKmYg9yt6v4I9+7kJ0xixzcZWKUq82Zgr7b672tAnf06cg
6F9YeL5iLceXrKsqWMuVWpym2Yipo5sJLp/4IlSJm0hm22ht3AOU+lMDXYjoi3dG
SSJc6afcHdwVJkMrTehi+QGz16HSwgML/47A6podfzTyd2okP9HcX5Ztq63/gdst
y/n5Of8FIYzSQTnRCPQdeo5rrcAPtKquzQZRIlE8dIZ7+GZ7/dsnmmeoxFS1hVtv
yRZFTUR59JErITCPW3fwUBIz38F5njHw7YXDO40bl6UAVIWmrzxtGQz/Zzvh7O2h
umBYKt5GoBMRhQEa2W4+zG1tn4ShEWMl6C67T6S+R50zKdXXLNzxMjgsrBbupnLK
uHBygDjwvvSMkptvYMfkuwdAPFEausCrMyLp5blpcSOtbraGsiuvNczsWIBrvouB
SdITJA9c429ffCigPIqKeLbm63bs28uNTQFCJYi3B8iVNKgv87iYMr1Op2C9X42O
hsnDUsn2XaRFOP3iJZFTT4auFd0uvzF4/RQG+N8GzzEeonkmEvK4BMmBmAtZ/hOM
4T44E2WCIGc7hgp1YCiLU1KWTL3tVtGcatlKHW64sQBpZjijSaMjvgR3fPahVn8m
RANFY5TdrqUcSIUo0nxOxixRgqnhCmmVwbtf62pvFQdYrGfvUjaeX0I87cHXnP6h
NAdMP6zyLVSitzqLN5dB/skmMAts7SNwDbw9naECfyQyJl0+LX+rSIUBS552N0Ii
UX2B/TZ8oPOpqEC5To+cH9+HUtgF3n1S6DNCi5nSQCQVYQPLPKnJ5c38q6PmLO6S
n0V0Uonrnp9QVlseRprpgoKFx8Zpi3kpUp0B078nKJi/NeTJPHMQFxr4aBO3HhcP
di2avtGkoVB3P1AD4MWsw1qu01R17kmNb1c2angIStj7BOMfhmFr1AWdvp8FgfVO
iTTcjAfP/rHMLdgl/q8pnXWb2x4K1Kdb5JFKFjc5VcuZRayptU+isEBTMkorQIIs
omEvPcyso9WXRkFhhWOZR6Z8URkr1xhk19zIh5Vod8PFp4BLVs5Z2u1C1sow8aB2
veEnu14Jt8YXsZ+gp/nWrQoBnVAYHOFUNWimETyhqFaf90SJz8YGVTSphaKwTFhG
MDng6HvQ35Eqnx+ncVoohSTzKksecTvKguswVNtc6fGQqzzTEggYqqMP5QBQdxrQ
ZkUkX1B5iU1DJYC8ZniKJW7T+S9/tIShsumTwcCumrab3fUCFW7RnvrqBgl2O2D/
VPa8k7O06tlhc+p+X+4ZaKF6qxe+LRztVgCIvGRGR0EM3+1UEKKKodNM1NZGgdIL
V5s9Cz0oTQsFICwZX20/3JDFlS3t/4V+t9VwzHqs8tmMWQK0GydLQsm2Owylkr06
FpFeUTKGECNUUpJrO+NoRIi1whJ2N4QiOMdOKEJYhyZofTbUDBAH6ruCGFoQRYk6
nQNSz56eAyxh5h0vmSDdpweACQ8S8DkvWKxSisn1vnrrnqQJCqGDFAaFxYwtU9w1
Z1doYW3WjqAlHBWfXb/vfWfr6xxjDHZjYKJv/5HZQjSyCZcekB3GqEbysOwzBugH
bWRUlYRXWsHbBbzT5NHCCPGDNgxSDHU4AXFHqq1+J3xwIc4o2/9JklxLQtTyYcRO
KkgenbhIB4PX+1tVbAFgrT0ailvAoOXcBU39dKuuajKtc0yMzmt75yru8IBeC7cv
ZYthuQldqxkenQVuHb0W6M8z2JIjcC82Pqyy2riDMr6gYyiItNmR24M9/ppHwnHo
5viuiuWQcgG0rYSdeS6oZqx7qI+ekgBS0Afq4QhamIJ/7FUbVyRavoRkYnyc42Fb
pJpjVFYKEgVNYcHL2WHbx2BfEXW6isORpT+iHcePDafDhenyHPV1vWI/vKBDBCqL
ghppqgXO8vTINUxKLfiPMNpyBsUnnXoBQbsDelFNjgOkcUbeV9TgouJelSkY0njT
tYWnqW1Mjdyc+j39jhm5pIDaJ/xU79rZVhYU5KmEqKC2Stn8Oh0i2Q+zX5Y+E8Zs
UM3i5FUC9Jxxv0tW3bGH4tkPSS+qH9m0EOHFJU+w97NpEC18YEp3aztJy8YzfQZ7
5LXa9P/aG/yQsxgnhGv83vbsXy4CktnxgV2UsZO9OsaesMGPMips26knkZVocqs5
Vna+KfYhKQ84A6fesoUewamfwJKkWuInXnipLfeRekh3nrbbWZi/T0oDYISiFqPR
0swrxeom9C/Ui2N3CTElxwHc6CkQDmDvvkto0yo4RLmQIxF3teYMB70LgpLyrh6o
hSKNoYA9KYMVJ61wiJ9iEdmWWNRiqcnDOYCWnZUYXKVXJEHAASYF2BS3lqtR8YJe
ZDS5Olt87FUZgb+OTTfQ2XDU4dXUmDuRgew6vTf5VKuBHWUS2BxIJlUFr/9/yF5V
hjw8rqiCDhNeLpAYdSm7TbR/vrmiRGNx0YU6S58tMBGjeNcIJ0pAs/75m90VcnEl
penrnxK5DYOAY7DL9UVhuNh+RU02AqkriIYvT6i2FGmO4jM+S9snqtjI8DQi55RT
zcqcfrvRNjWGkAE2Tsf4zUrA9UezMfQfZNLt2fjA67b+c+NR2nitCTJyI5ctZlYU
PrmTmBVkTTC9mD7F5WNw1z/qZ5xR3k7Zl+N5W+Apl3+P37OrjaX5utRKmQ99IOuU
Glzcid2zEyClXJWyvJMrciydbDdUB6mMXTPsm8DXgw/12zaGVv2RBGcA/FuJEC3s
8aGsReihzsnM5O3axUUPRzKnFTIpxAqspHup6QtDz9WiohcgyJWD+IHsC59vUNIG
Vuq1kekpu4dox9jK/Q+HnJPSsJaF3cEk0FX3r0odCRnVCLxLrVxZ2zbj8MMeUNGP
119h8nQzkgthKSd8+JUHuKy0IRjD+7bAE3t4JrIXajiCy4FioSYXr2FrakXTgjqW
H/LycI/PTzTeBZr8Xm0WJwqAkBhcFGd6wmdDhMG9DhRKT8lI2FB8Rx0mw+0M6ANX
zdmvy3jNGPpshM/7rX5gQ0Suo+UxfoF6Xj+Pn3xiwP0hgGAN4w3DjM7C7niG6TtW
XzKafoViRBbxvoMxCg1PBl8AlRnrBvHC/MSox6O50M5RXHfEanxIbHRWZzXdOKwH
kOR0JVZZKx+7mdONWxbfuROiFTCwT9K+/5IbtA8fZuS0AGCHgLGjCRVqB6zCflt5
iE7FBZWoU6ai4An43vFi8AnGZCVNVwJaVtNWY8FdUR1xzE+0I0ErVTVTAi+FoR/Z
ECc4fmeWig+JEhEPqBvsaUf36Sq+yXHe6AkY+d0CLWylu67XJ34MdmfwawC49dpU
qE2an1y4lwDHAmbKWzq4IVYMlQ4+GcJWu/J7RzERFrbsTuSk5qdxt5b2BemD5CpR
KhSOKFkdWXyW8idWEXqg7Suj8L8aILFef7J/8PKOLO5QhBY/ah+sBz5rZFFD5dQi
odwk0+f2wLry02Y+y16pd6YTFvT6pLZ+qMNFU4wXw1uBesNUfEVi7JJ2SoGkbPTF
o/xTqynU0t7a1X55APNGBea8cvBIzScLnYvGsIGoEmZLcNjHf/sxAMfyTiY0f5+r
LgChRPfJfZgQJlcwKxKqXu764eSpeXVkpGeGR/TvfOnV55cM+o6HXzGgGyWrEknY
ZuEVbXVY8xX7gxa2azbIT5cG0OJBxxTf2vJxuryFvPz7tPAng7FZdpKBnizZasZg
2CDwF5v2sNTNHe5j+kzbLisuVftQK9+fnP3ArtB6vn/eNuOFTa6vMfyiBhXTrY2q
wtIl3kDIYnKWKn10/T2s5VorKyKWB0KAbBhi2yJA8yzfBetibm1wViy5ggccmYdj
FBYnTJJMUEotg80SNmYWaZ6BmYnRdgJTSTkBiK3fP2UbuyeXK4zkgbMuOOnM1X5g
hKgE0jp61py7RIx+M+jxRLNRhFEYHr+ao/4ykzTVsPyIuyiLT9LMGKebYSXc5EWB
0nN7IyVAzG3H345IMfzGpPIl1uV2uuVjdy0cJ2cTzsWON5MKLoBKCEHnDoqilGrJ
5lVuXGJ0iKt+FEOKH8MLyrFiZug9x76hnAPOyESpjiWaq1d5YVkAKp4KVGDSDJ4c
9ArDkMVN1vLER6NKRnkfbkS3SgDqMTF3F2DyBJZaoPnmiDNYYDqsc//1JoeU+uFh
XBkOaPKRY+0z8T+fVwPcvseaPeVBodAe+YVJ9UlrMVgkszNVTLhlIXg9dwHdUyOz
mYHHSawt8uxiFZ6nkWffqhVJd+XYOFKCYNvFWrcoMjNoEFRp/NNEgxdrFNHbuLJh
wuXGsu06houFmdPgCPuN68gdt+BsRerUAuFTA7pLpcGUX1oW4d6ONAjK9ZXY2P11
+P6w6h2iWHZUxN7a3kIxQAe9+9UItxOmQDw8VTK5zR/HKOI0Sf8wNTxJPZ/RAR9P
JQuHAPtrUwRDe7ciIHSfcZ8IV9la20I+WxgRn32UUblfICy0Ez0h7ljE+lAxTN39
EYXUJ7uKaAK59dKsAavxTH8Zd+dBvIAWadA/GauER9HfKYEnjZiEtIBjtHVUbeMV
GTW8/TBNjz7G1GvUqdizgnq8k+Jminw32hbXgW6mEmCXHAmynCE+pNCMdrEx2DQC
vgoujuU7A8S3G+cZJ7P1Cn6J3KNSgio4AGh9JguhC+JWy6ttBf10ANPoUvqUfB73
iO//leTAseTS15gyVq6FxQcV4YeXLgmJDkJahOVOc0cQFj0+pKS6Z3dHgnVlWR3/
Ffpzh9zs6u23jn20469LstWB1NlMyKPk45+XkN3CD5ZXZzt/0Lhnc1UYBTUlkaIS
spmHu9YhHIv6qUxw2loWrj2jbTUmZgPgNHYH6hAtGmg2+i/E1Mw3q+AQnOhXAgh+
ac4iLhq4Tn32OvsPyMU2ZFHNA8Ob641KoY3GfxoSj4WAnnBh6/cAR4DhR0nIrIm+
v2dSHEdm8nRRgIiVv4Ru9erFI9sSRfH29lHuJtr/xFZXlR407Zhg+auIil+Q2e8M
EzvBOY+Xfz1dBDvPuJpdiw/2YPr6qZ1s35HEaQzScS36nJWcLSEXk6i2kE8mDvpz
EjZTQliYQGW51AodhrWiATl58BxLtuhBk4MiEeLFEljqSD8wONheb9njqEmAeAep
Eh/pAfe4G7Z+ec+iRstfHAWGISgNZ6QDHdtvDRGsGnZEnFUJVpzWQVQ+f71C0sqR
pGOM/cWK0DWEV9kwbwpETPWRSxCo1fZTI1dHUd5gGfhTu3zX08G7IwpaBnlHDrF7
wDAywsN17ZjXH6Q3WZuFQLtBRfhHcbLvoQfJb7xEVdqX5CkBF6dQ0F43TjVB5ogF
c9zjNzeBWVr3IdRJFe0/z0gtQs8cddeYFtSE6OuR6cqMKPSIzxVeCaXvc6jwVONz
s9e8ViBBqKqLvJ8GgUyyQzpDQf42n6kLPM6vzHeXW9gaEEXNU3eFzpyOwKNqT8Mp
xarUfr3QyYdXsmUFbdiNokuDcO9dayKBluNRStnPNIPNpzwWhlhEABqULV+h2dCN
3Pw/+tPBCIrKLyhzxado8ydLC5TSJY7BdbgmW3mMbOFhthHGoPwPou/lZWy35ytH
o/EwqkXbyi9CCgzlkFgz+aS0qPdcLXtJjfxc6sF322dpJ1PnOle7JFIzCFeTqDZe
L5SJCbO7IqP4OJKHZIgBoZSScCveEw2kCktnn5ZHBJoVvmJ66LmurSy8+twKTz6E
Sj0dxF99K7dInsk0uVDqRExN4dHRWZhCMOZRw4vedPVa2jhpTheRJMjYuj67OoeD
/d1ZrzqSuW3vZ4TIHvpvpR6HB4PZW0jlwiDjPnwrG4o0VnEo9iEiYktNCUiuI54s
sFHrJXwftlaaw0Rg9wd1EjXw0E6u7L0hxROQjiSeXMFziygd5+8+pdIB7QFUjgKO
QXbOiu4dU0OodpxAQWqJFaoN+qAj9skpg/ux1FeSR42jhwV/87zZYysMQrxMdBe1
9vJvMwhG/lOrXmpdbKQtdxH1H4UZbHtQjJnzn0F/TQpt0J4iadUB1C/nG93EDjv+
2bp5tScT1IkHRa0unE23d0nT1mGId3JFh8lucNFq22oH04+s4tE0tvudDQbqivPN
L8HOfDF/p5kXzyrtn8B+C3tWstmlSdqpuFNRE36p/ZpCHBvoaZevYmWfc0seoITn
cBn3u7EogQN8NtJuDssMfDg+2Bn5NMx4edCjqjbEH+pz2kYa1sXh9qn8+m5k22zd
baJdKbivd1IxvSlF0bxZ0f56yoS0iwiTe8oHojBHbyChQ1tk976AA/F3b7fRdkJL
RLGQramfhXzkPjOJiDpOAVB4I+kTVlC7JB02V+pIdJyTHIZaSIRBYcuUy/dy+TdJ
hAy9fcBvHa3Q/o4EI3ywHAs5rl4X7na2nI0nrNjzSeef1XNqfbPiVh35G8GNNOCB
sBhKir8+SHxGvILeuHrmQKJKs0tq6iSrCt31Bq4loz2x4YH1rKJ0M0O54VO7bH8B
vFeL3cXuNfwHDkzebSEAfuCOML/OmoZZ9oSQhAMTlA9yVUz7nIWcDlTT6n1ycqo8
I8V5VLONreizP4EocHjxZUTmaOQVWgzgD5yo9HXBA1wfcLrMkbOqSRht1PWW1ui7
LUeFhxpOyxfQFcJqqBFce88jpPjKXaKX8P6WaTdMAsC5/4X4LSbjOujd5nHtIv6g
iLr0qC0r+9nnjKZ/yYUJfhmnx6jQstA6Yln1aN5d2IwgSqjhWcLxVm7lDeitKoWK
wkSWuMFe5f9dJnKy4tGsCT6251U5dqCZprbuqOT2I9x8tINsIaCP3Oyskus1fVUP
46KNe1trL9n1DceMKZ3Px+1uxFUfHqG4X2+CCEVsf/k5E41ow+h6BgJAKzKPt/F9
lkUlUNowWU7Gs8kUBkfJxp05cJ8fXa16iSmr5/vVUBEr7qfCCTQLRY5ZGZmOykzW
ryq7KuzQEcjvGILWiTbqYT0ud/AUU0p+RfA/Wci2W9boRe+0X/7Ja2T02B1GJae0
+McfdkT+pe259ykVL6oFPjFB/86Xy7OpVeTbB1a5ppkepEmsEzVVy1hePtL7lx1R
wUYLByMlChxGIXzF5UV5V9h768K/8Q2Dku3BWd69w1c9D6Rs0biGXxT8KER+R+O5
JjtBbABfOD0VpiMu2xs2qlQKOR/t3/MeBSJHsL+vOizEFsNC95Ttc4H1KupOOP6r
QT5VL8AptMPfHNKDb8f1LjEsnOkEZVkAPzbJQ9I9men5C5mHfoXM/qo4j27+YaIy
NuRRfaEZeYSQoN4p8oRP3WaguCI1asd+ztYObxMZVlRzRvRNP3xsgf3rSBkLJHsh
zmcgtVK8V0wiH4L2ieYpIIctvx/eXZdRgzt8BC3wDGzL4BS/HbPsuXvbRhOE3BrA
r/M8mcW1XL3P633zBMsj8JvRRtrZAVhZ4Ik6kJI+DGH8jTXONK2PO/pTCY4XJ0j1
wnl4w9WkBHlFLcPPCjCK9FYhReNHqRXVdG8L4rpmLFd0eJgnbVI+dvrxMMVwBPqB
m6wVamlI3/0Mc3L2Kiic2efycBizy1doeW0v71KRXYkOdCBwBHB00WFC0zd4gF+X
lHiV7r2fkhC/N1MAs+SdrDpLsni9dwgyoG0s384tYTHd/vQn8PTJcK7efi+mXEO8
Z98pGL/Bo06epT0OaMrSrFLaYeIvxnmFpUidgpVje/yLXPG1AvrUtnO6TNj9Y2NL
r9xMpowfMk1Au2lXloQCMjpcWJwcUgnMSggmU4+DSkReXS+wG9t+YSshzCe/mceK
Ok5vj5kU7Vjlihb6wTuJGYIoupA6C22t3YvD2VZwfUAVoi9iPf3XasbN3F/d4K+4
9wj/ufDN1BzqxcG9+ztLmtnb2Vwck7UWXvBj5if2kslosMEy1F8jPeBwC/Fd9+K7
jcS4n/TZjNvV+BNH/IdatGw/DzrtjVpTbwBcbJSYBp+Ybkk5ChS2dFUDT/YOABLE
XlWqSDnJx703h/BibievGCRQCK0qyJArU57lUL8DRHSjXKAG+p5r3oHcPjWgnUfT
KQxwgaBxgtqGCQJiFh8wtKxE23dx5fhWcedSNMRTXkZTaCtedjr7unMCflOqB7YD
L6x2HRsY8W5Hj+1FkFdMs/LgQpsn2TN78tJn5qouDoUdcZ3P/0pxNnnSLX+Hly/K
8c0+NNRQLvA1gZ9ynNVNR8ZwGI7z5LgWbb3t82YvCwHzZXbee9S0XnMgvuCczaGw
YXarfQCWk0pCApSwMuD4ZVGSRoLJGFjQOMlxE7VKDXqCiaKVm2SHLrUzJfswGVLP
kqTOFizIfbrTAN9EUPhYe5dVNA758MeUY05XWZMdKOqC7y4gvICFTBsPBJ09S+DE
Vg40TydBcU9IUvS2+Vzy/mbvogVMulc1SaZocALPYFPfCr1v4RYVNdb18gL0Bx0A
uAI2/0zm2DMekJj3DhfVeiGjln/dKcovITtMn9fBC0+tqMrxh4BFM+SDMiTacSRE
TZgJo408MUecvgblvvUdsffMPeLwczrw6MO0u3H5qON4+ypG7UmQ82ZBK8uPgU1t
shJ6z2W6lEBhKOt4GpW2m72KjjjK37P8fOWrRQZrI/0c5uFb2iTNnhAsQOBWeHQ3
L9T5YWjaBPuYizDJTihERbLKG3HtAVyU+t7IqABXv6fYbdreSABnXCXB77IKEdNO
g8VCqkGpHOo7Bft0/7BXI951QEOBy4zysaRhgz/0RZMTtpVrfNsz/Jh1TOVcu6jA
c7jriJb7f+tCzedTC9rOC16Zsmp1dKDdXZHcOASlPll0o/STsD25tyRiaUmOHgr2
z56AS/HuYjtlNo/RDlW8QaRwmsgagEyqJumIZLPFwL4iL4Uero3QoxhGNDC0tFBJ
zOrJBXeEJs2TDKJ6mbF5PqcSJwWtPLTutNyDk2HNBBV7NADAKYLDXRbxKUrlNrUw
11nshMWQtOCDV3HSuYP2NHOm+SLSUqHJTOCCnyfTJsDrmtgg1miRnC/WjJhXXISO
gSPoJClCFO0ORBvhYuPmlH8DoVNZg9ruhVVUVe35SF+JH38wpeNrLkrtKgvz6TkM
9kRoQXgl6KS4rW7dFGdiK0NsA3yx3rWxW7MWme3PsfqWioVlpd0tZMiUXra7spyf
AIjEnSoQkVau7G86N9N7DbLTUwXG+8exh3XgOraYJst8gyomM6zEjV4Cu54BRavM
gWTjwCJkRqC+lLXlpWt5ktXj4BH4zS5Gu7tSXipf23pLNWKcwIqShiBy3GHA7dvE
mZHNgEBHm/k7zkNmvh52JV4anFMnoATiGqLTqwDgwsApN45s6vwmXkDCm0BJ5EpP
PeaMxFRK8L/St1INDthmxt4PzUKJdKR11UUMIDbx/063iu+cAnYWsmYlbJUQagyu
+i3jsunCliSV9wbyLNp8bks91hat7vzPgVU8yT+OYJx+F4d6PjCsNzdOGHCy1E+h
yWKfZNm0D2N6aUegH8Y+EFMOeSt+0nB70q2SayrLoJJlJmb5Dxi1wjgZacfA3JhO
B53cfT4Iho4POK+vT6BHyZ+8TPJNNls4sE+08RgDXVLvZPLwV9Bi08yRPrrC6lXQ
imCwLxFGhcav6z4w+Z1kctIm17sGpHmNM+T+BJXNRsUvWWeYb4caTp2Xne7SNiO9
yNjG0G7QJ3h13iOXC97QfcKXm8y750FnbRHWwFbGjsbyWksdXvi1OPN99kC3/mTz
AUtNt0ZZg9C4LeJU6pAOhrnCa0J9dd6CueYppNOiGvo9UEVgR8d2bevR03uCt3MU
HMWbdaotfVaDt4BAUe5HnYlYa0P9GkMBe0dpVUoUWu+6gY4XhzZINnQ1vCfZ2Thy
0xCV0GZJAhVlQoCJlesliURwwSs2IlnepL6fb78eWs2FS2ZUVC+ZFECaJIsBVIr1
Y9tAJZNWfmdXHEy/gLaLM8JON4Mj8bniPn7XZETIHdvpv9+LwdhaS6/70o7F4++6
i+3R1t7yHTEgOyVkRG/k87TpZrJ/BidKUZQexhqieaHLgWs8qaJLUy4KArDTiI/a
cBi0u9Ss/M4vdb4WSLEYoFQpTJ/0w99DzLtJYzS3iBu3gVf2zy+12ODHuIJgijWK
1hyllid6snshvrmJz1PN5sJRNq9ZsKTDuhWrMxwDgH/9lZ7CZXrXh+lI8ucl0Xo9
RQIaHJAejExOJj1F9tXFdDWUQP9ZrhyzToH2blxBmkOl0qJYO6oM3EQwfMnCS2v2
DZgr4hJWF8Qa7//a9NmVKH4wq383YgetEVXup4rA/jsp3Lsa3+gIB9QQv8y7ar1g
n+mk53Y0Rj31gkacVq4EJJvRFufiJxTL7z73Sw2q6pvmDlDbCxzlVoi1c4nlRLlZ
v6X4pn54fkH1lrbUEZwxuurkKHB1KdCfVzES7FHXt6cCnsyEtEjOCV3s+DvmQWzx
qInZetrsXBw4vtPzoasWcpfaiTA5EmrBORVKJPJ5x5XTOk12cpOPqL+M0fNzn9j8
Lfg79MctMPswTS1GJZezdnNAXjGYEDw2jBuqkQ8efnMqJvsg1HP4jxewy/YLCqnM
wun1JuDxZd2jgBX9lan1wFVMPbhlrsY4SDiyDpwH0D380UIjiGXBI2nIghx7LySw
sCxpR60LkARkIigSJgiP5+lPF7jfGKjhiLhjFp09qN7JhrOA2SwMgzNnuH+UUiJl
BTVUhLDFyg274zhJ+OdSu3l+ChBMupX2dZ7f7yy+CMSASfAwS9AWv7Ub04oEt2TE
GEa8DlbC4A+fVkLs6bDKzhAezCjsdii5dDcLL8lXDqg6wZ3wB+KIvSmxxbzzksa4
EZZ7bMX69Tt5rz8BYV0sLydUL5YgMyfaCrAt1Qa7W6dIvNxudMTGpoO/ab96jwD3
a+LRc5fQcp+p+mAv9mrocMsoz2J4ctEcO9lNJ3BtXCEL6OhjK284qJp/ZJtPdO6l
tl7YI/II4sfVU+TmK6qap/IaB7THY5i0oeKnzan17vGaHtFeOw9wLUhizxy1RksA
F67tH7/Kfh7H9dyv/iXcPvk2C3+SYEBfVGo0CSV3S6sUF8yNu9v54ApULbKlq0nv
AqbOGGC0CqVCXN2PPCj8robsjk4JH9oNLypunl8Odm7U6cZJw3+nwZ4rbMTTleHS
jMl/EeR7xNtAf+vgTUtbxEnLuCUzSSPAW2r1OtTUA0cLsoPElzQQtmTk4c/5Caaj
1zkWJhJDlIy6pdG3ec0kofyJMwZj7/rJjVVwmY4DTrU3fMnlbHBbsf+/x8yuYGSC
ick3hm71FmIwxpE61UcMNTk4arq9zNyUa+8XonSo3Rf+9gHDJQhQdAbGlMjdUz9e
4W8dI5wOVN+U464hzSofsTmJWKZgF/RvD9kzlG42VBH+AAaedfX4+L8jzjojVpCl
jLAsysGdP0la6UgzyCqnJ5clMo7Y7UPFUhyTxf2o3jIGaK8IGtRqMjVlf1P6DXl8
3qmuoBVcg+VQdqn+44sO/9m0A3PIxzIP7mORU0vXSZZYgf9GCUR2A8EOd+FbtS1t
YegyLLC5oKGxJDAdnk6JLxoIImAkajHE7psCmaGvQx5rOLVJJaD15RbYe3+LwxTD
xs4BEM7o/bJyhiDUMZOA0rZAKoecaXc1gGxcYBX9oRWUEZdCldeIpJo/ZUwMF8Sv
AkGf0wXmwpdYLV9HdgMczOAPgQolb89OVcbcjjw/1W3Jm9gH2j35t5zJv4X5AG00
9h2BLu2gsDg1G0hULG7p2Pc9OqfTUIAVlTdueD0ui7+Q+ZmWbjclTh2Pgfvt++8N
F1PZh034i2PUpq6IIYUpcrZkHmITAfiyRJxkJVcQataX+sJzAhyOkkjaTJq837Wz
NP1qdsVRMF8o9yy7zM+l4CySUkbAwQs4LcO8nM3A0nOQlPy5bYwSWg/h1plgt0zJ
IiOtkQyjgTn5LtqovdEllExVmMb0Va2cBHlHIFUtc7iE/SgLlqm7/+RWvuipfFCA
uEK7zly5jvakvZE3OTfycZkFS5PJziO9U+4OHk4bHkkIaXm3bzLVHqb4SPFXf8Hu
Xt/ko0mKE+Pu8VZj8uRNde0yvV2QM24Tw9azCKeYTxCXejDcfBZ9n88beXGc0kZQ
Nb5B+irXgNrnevypEo3hwblMaLy2zOxr8gruT2DNerqXBhlkgcb8ot9RK2kiSQrK
AHHfIvgfHL1KlCnmSGX6IOxEhwrruMCuxf+V8s3k+w0+0yPodrmphQrJP2Qu8CXr
UJSGQWfBaXaMD+X2QXGBjR58BlWyQJJX1LkFANufuIZMXv2DXwl7VHpgfn57aajz
ox7wdEkzfOZBLoGxbxK5T0aVjuNgf9GJNwt8X6TTzGabV9sDDJqul52cIjqp3+sr
ZlNUABNnvPQ3cWoN/shO2TgiyHnqvDkJ5Ls18UOSGiRzENeIumV9jfMT+FGg3qDI
P1o/6gm/d9WixUlOQINwAoTbHVxwEAG5g2hauCkqbxgaIeBMLrousYPjK6xay19c
WuvrqJ5q1w3+TjGz+PhX63mE2lCnuaP6MApV6zV9xU3zQUC88jdpwOque+K0KDw0
smUN1thp9TPM9YhUl6NEOnQMmT5RSupqPYbife+96fUZXWmb+mp58wljf+0rBQ/5
5YejSMf4+o8ji3DhZeGoYMtlB0l6SAsuGjRj9q1firNGRjyi5WETO1tVixdAwW9v
FCAjka7PQZ7wae94/7dVBvS7bO7VWPoiZoLONmy7Q2mohpARRJdVIyKtp9s59CJF
kBTaitiofyURSXKR3j0c7IjsUF9EMRVuAxFMYDD4hO/j5taEHUKYeyy0XimKAeCv
M/VtGtmpTQfHEl9zyD+63OE/491pxgYrq61EEAUAfgw/Z4sA8OZd0qQrxlSzNXX6
3UZtGDeiOvqoiwplsr6FPhr/zOmRvUI1GJCwk4mt/BaVrFXlaXyxwQ9E1HWnMoKW
cXmhqVBxHIKJh4i+b9pLkUbsVClPJMr6izvV49LkVe2eCCdaGe43Hr79hBOKAPgm
NxnSP1j95aC0vxfhdcIqEO8hxvKTrLaUcGQ8sHMqCtj5C+BLwoIPXZ2x5vfYKfTK
r5f+kQXusMJ2i9r45+RLPnlm7zcZb8a+ToMcXl6o1r/uzTWSoFscW4Nb6NcfGMWg
LkrO1waPG0wn32aeMkOvlLzXYOejQAuNh4NTP1ygzg+/eYSvk5rTIKv+2MWF5GRM
bDMvgvrejszPqlEBrMKJY41RvWS0DRzv05p7r8SzY0FTCG1kv/Tr44MzDtQBVquu
Ta1JHOQz53iRdEynxIwI5toKvrCuRDXEDybdHTzjum+nSEGMBG7Tvl4q7B19S5Yk
3VJGSPCuUVWeKzlyBWj5BPZ116f3YP0REM5kPTQH2HgFP5GvZk2bdt3ydI6IHsFO
2eIrpY+amjSx8kEOC725DbOqZa9jhUuB6kKmWba32/JzJPLCGmjkFrijEH7R3wGV
kxXa6IVTpyKz5rY4yriDefLlPS/KYINZ8IpJYRRfW65fKXy8ylSTMCGMQpj+9/W/
oQOwxO9P5C4fDovq90OVUPlG0kGjYh1iDzlKY5UemG48ZcRtrFYd/BVFCVc/NCsD
wo6nAfYZERx4i46BbEaEgNt/J0S/rZpBzGYvkyx8sYo08SvpZkRH+phKGFm39FJc
YhoVey/br1Y3Owf9qMQqZBBCa7Z+ZjAYoum2/Ju9WbzmEqXcovMEJdIvFPU3hV4W
r6mpygXTirbM+SMMIE5Q0IrmwvyJvroXtc1c6ku3AJayiGgUR1z3MBT05Y0Ww1Lj
rm0xznIkBw0ACEwkkGLSefRkaa1kpBDLiFIpgvZ/d1CLGLL/7ddB8OQaeL1mF8J3
QUj/GZioW6dUuE4Vy+FaDOE8YDKs5Mzd5970KFC91KQFQs5rdtEqCKB97QHBvF2j
KXYI6o6AfUZxAxG0m0XzxWPXKCX4tdo/m6PZb54GG+JJaNbA1QRcRDkwtLkTPdu5
s36YB6TY8y5FOj5W77B9pHgmo4gzGW/xlsTMss9VqenmjuNATXfqgS8MMme37dM0
KTwf18/duUbwRYthh60l4JxucAfVkYc/k/Yj7sIRRCfKVSewRSzUmpyxZqaUT66Z
ITM7UGXHagjBDhYKpXjkSbOPa1J5djOdLEYZaJXVlrzhro80YbaG1f5ENNGM+S9f
nAdqEF4asOYjgAZu5Sj7fxYu8bDR1PDoFq+r1QPLwQ7HMMNkzdZQR8GG60qq1e0K
2qcXDkOFywojMgMT1dmN/PS+Rs6xV2DXjncULcdZ67R4eluI5lC5KLnUWhSVJ0yM
3BVVBRzWeH8jaj3GVRGigwvRRIg4IDiBBBLLRDhEMKgW3kaqQHeJMIRWmrUeeErw
YFagc3+IZ1u/GVZWx6APsJwu20t6D39O/EEarLxFpFTGUDwOZVvbrfomYObVuD80
f9UKWa04wMP5uRKhAiNniD0RlGeDo9KAFWrXum6dXoPz0Dj85tvrD85K5nMf72ZA
f74xJNFleN7roZV+fO4AFAj/TfjTfTcFh5sEA5LY/7Ff7E+JBBxhI/u8lhtsXU7a
6b9w8SYlWzWsDs1kRLdGOeA/w3K/Vmuvi8j5/PmtZNo1rdycXCOcTHmd/Fo9nCW5
1TpTDTIgJSA9q3geX6Vu0l98hc8FqBPuNFZ0SxWzufqfPsig1zZgrZ0bgE24hZpU
q9n3p+RXhBSLJ0EvUl9n8Yfru9VRDrUINHSVw9Lw/znsfElFfQWdD8FFgfhzhg+9
9xUlHS0k1rfsrhUoNc0AMaMIaej9BMO93OpJYG9+h8uHvCeW15Jy2TKs08Y6IwM7
/nuKzuCC39REVAKYNPqm5S9CUI8Q1Jh6UCkr/8bZ62/RLT76K+qFd7SVYobKbx8R
y3tPpgIB7FIHpAlKNUqaI57IEt8NhcQBmP2zzYRKNJkqDHaQl61kIhWxBu6IVuBh
MWyhVrBBpiCjzoCyavppcShrcc9MVWjnji8HoToIZZlaOqNLCICyMtiv9hLowg+l
F5ysyfSDiSfHEhOwoikepT5qM2bEr6cE37FhQbklXSemCZYKg9gYl9y7076/2Eux
148hE94eIFgLjDAKLFDVEmgkm7rPwXC1g05dYn/miz6wZC0LXw9WJh4b9DAekQRY
c3TUZ5GSXVyiSRPgGj/sNFX227NDz90qoVQDFZpceiGGxCtOK3gcibi6nmf+MUUw
oqGCvfI/id0cBb4mFAmLjaZgnX6R6q1LvYV8CVqAND+4iAeXVUJCRi55JmSgs7as
KLpGem9s7UngjQ/y02sgaiABtiJFSfOXLwAP9De2DN0yheyTIhY4X4LDgO8Bv1Y+
9pGevtqAlJixZECR6mkLOgnWR6lSW2jskgCf9m0YaNhrLrhXXxQUhvtnS5n7JVxD
6XR73SVnWTiNd8jFzMTurJ/LB6F5ndK+hwwBRL3Vm2f9o2Ia37NleFwWIn95xsmc
rIvmdBhETIBbWxTOTNZpXdTCm8wosMmUU+b/TvEpdryOKJ7VGMcDxZIN1H3Pngg4
bykBtVnvHEgYLCpZQGK/mbnEcXv2LWvbuIe3bFYD/K9l0MoXtgIMGa08yXHYGzoW
iDa3yvpDr5c63rYMuErsYZ3Dp+972st9pyn5qCsZw1LFvcg/dxNJsv3pcQ+yhE9G
HwjnQ8rtpLg/dkLJMU+ehKDoAcih07Wv81fnzY4qyurrudD0phLaHnhXXObNc1uv
fI04BemPS/bhbhjRhKSZtDrE53CfqLvWS2/6A/bVUid9KpB5IfCFGDZv5M+hQHZl
yni9E+JEr9pp8AGq1t8TzQae+YiZ9htdVwP8MU3Nim17IrTatZ7Rk9fhs9pL6k/F
PNiBqjU+ASLxLJWzoVKOa/XnNX/LeeD2vLn+Oz7q4du6W2T4dkCx5gc08jmA9Ikt
pQwYPVqS6+yC0LVT7J0iRdS4Lipw9M3+ky9W7txNizxhXl2UTABynNnse4bpHM8a
va+p5uIOv34SKkujw5csXXdDdpnDpFBXQuTTsfsnJEl3PKPdxKZXeGuMDtNNGBpF
DTHQ/6ZVxNKpYZoI2iDn+GikWezWHc/3yW0C0EffnUQYWQZJTmKXtTPoT8d3E/AN
1N6i4ZP24FhpTqNQslt5AWUFRs3O/yJI3v7Zm6LEBVoMD77aV+JEKkfNN9kEwvar
+0fDnNMIbg0sGDQcDdcAf8aZhXEt8SqYFhjSUo6WkkV58mS2hGv4gGFHD/ZOtDqJ
lyuWXuEkn2cEm8vkn2eWy6omi5e+co/UlASglZOGZl+5hwnisN3OY25y6jZDp8Su
iqnzvO3bO0Enm5ENW++ivtPykxvAvaALx0G141vL4QsE17eRQLVmH6rgznfAoolN
D7LgdJkbVHEFMYtto3I/ReH4ciaCzhX4GCuW8Nm0CFy5yzgD1miYVqYDMv5VFZuV
jfDHE2YmrC7y+u1XAiRVgL788EvzKExXOLZ38f5zmL3F9GO4bnqZDbh3vkaTR8p4
PwEmdtEPrVBjKr3fd9g+EKEY1tBgfsmnivKYUYeLpUjyYsOgdMyr3Hq2GBs1dOHE
m1qgsyocGhCBi3ol5MiWc896wpottWrDuV9iY+hyJPbIRA1CQCvZkUWa8UK9nHOL
yOQnG5lWj5qOgMRk2Q/0JxQ8jytFTc/e4HcpG4ZDre5+Lwx/x3TrqapA0Scno4XE
W1EJKyl55KYXhDZZ/RyCoJUJHjMBE6GHoqst9zQjgcRS1izofn+AvJa29JS5GQiQ
2/di1E7JpD6pupZFc4EsRI6jmqvNMj8esZydqbn4yo/h9d51Wf2NtX8SVVmNTdax
fh/J2aHKjF4LAcL6u8Zbvs5XzRzodZFpehZSspKkXin5auu0DRjq/3njaQu6P1Z9
EExCWz5sVDLD+QC/LpcR9NSkOU+rvDBV8le3wqRLwWjUSjfFbwCCSlKvSTRH7CnH
xLlTgt7p3iE+9USsTw9WdRn4iGpG0fKlk3H8hefJdpFxHNHzObxk2AFTnWYX+Ew5
kq08MpqG1OuHHRA+u25keXzUaF5Tv/CkY/kOnpOUay4+ELFPQ9rdKxhMow1cmyKk
boo8a3DIJDUmTdN/qQW/TewL7Onmkiurs+7B46tyLa37c9dQHZs9x1qB7cuzF5bo
i2lF+R/YQUcEqM68CaQt/YVrRLP/zRqdedqSMDulphzK+mTyE6/72oy1L3bllFw6
1jNX/Ypnh6kNN9p78WQ4LxrsYTGFhWZQXrHnfuTNthM+ZlPJKZ5IRSmhM0CU3pz3
gSFPOnk/BdJbSTC/BXMuiJLqZUlpY3yABVnhkCQr5s6V7bO4SE7RhEd6E/hB3Zc5
sJBpNiDQMu2iTCO7PmhrJ/avP6vUJllAOmBc3uoBDyYPuHflHysjdvZJ9SBwbrhG
sma4kM/XOvWA9NmFUY6A+KE9m8xJ961JpjY7b00P9e/kVv/c3MEKDavANE9+k1jf
tNg0gOtZ6g+wef41xmgi4IEaMb07drGzwnFCoF3YU7zMSSvnvsM1rFHljuboqQ5m
DtUIsVX2s7bJf6Wumf/Gl9A8U2T6j5NSugelHja/42manjrXE1V4QDMFBsvtV4Un
bKt0uXaj/UB1pHjBqo3PTW9TrAVwvtL4RGpHorn/gumJoNJrzbZhc7zu7VpVtwqk
RUxJ2+Il9TM+Sj9HphnqZtGia41dGEcG5DUHcVglM+yQ2fW3xpK9ceMnlSQMRnCU
iKfzTX8iZ1ZLV1fI2vh0kW7ZNXrOS6xiGwMP8ew6mW1SsxErpIpFutI9hnjhyV0a
qO4dxKw+3lsebdkNxnbF08s5NTpoOIpNy9OmA0G5r1x/ejB+sNL9rsWKdV7U9Ofj
gBKRlc/i17qqBkYZji67PqpRc4u2HN6wBga4RjeMnhpkFSK43xtIs5T8xvoVodCZ
5MjMUw+qzVn6XQo4jVBR2AQU9iAini2GWyXyzll7RYhyoXQIe6BgRnzbl765Qo86
Qy3tVnh8Zr4pO5XKdTd/RZKpdwECuB708Jo5TLkZxPSqF8AzfBlkqmLQjDf9alby
Q/SMMJPbS+/XPWFTExQVkQjTYtswcXBUCyKnYgouz0on7NC+rl5KcoKUGe5rjgCG
W/6XXq9kvf/jMZxluAQWZtopkuOPclo+Kcm5ZhmYBEgf87ZnHfIc9M9dnDjaKbr4
3ioyUmR82CkeN21Af6I7OhUhwRoOhjtr0muhF71yzpy3bmcyu7XrLEiYARmCFWL7
hbXtXRurFmEROvuz4yiMByyh2T+qzViJj7RO+5fkqyP6KZVZyThDh42ehO76jiQh
fOODvfyjAo/nDVJAMZLNUA8wrYf68XznRmLvsA83UPupHB/GbAwXFTK2KwS0DWsu
auHXMfOJ/ZRGHdouMQqYLT3e5s4xYEAr+OUpDIYsNLl/0MZf1V3NPHYg2hWM4SL0
aLJNW8gU3p3Dwk8WWOp/QDcKxQjzyOpHaLs+4Bo2aNSO3DTvUUQ3u/onPrLnA4Gt
HGOT3RUwlrqaMupq6Q86WJDsB3X18Q79j6KxWYCV4RLrssfuWbVtI+VvZyk1DN9M
DDIlRj3Ft4/vG4D9RhtlZIi8Iz6XrGy7xHl1gLCrzsYzrfIznqWNpfLsNcMzX2Jm
/KSFAmb28ptlLSy0DW8gHy1aQ6ntpdwtN1O8Kpa2lB/+2wwRipodjLc5Yy8nVT3/
08LjlEQWiLoT443YOLxGFmFx1wAJ/TI1Fw0Vka/Kcn5Su8TczJTgovrv2OqBcxiO
AC9Yub0NZZcWYLssENpOVWeBbP4LPbk8qZU6iItfTSR55qENPELVPNRhTa3kznIV
98ODe7nEPupdjhRBaWyVDWDW+4K2NuSfRjk2ziXTfyVRG2MltwnIj1f7TRdi+IJQ
NB/fJiMt536vlq97IGDV1tUC/FxIjAG7SU/qTHkdD5vfaOrwgLdhUsVz1a6gcu29
DYiUjmqcasRxSI2CzT2gjJEBDXToTGCVky76sHRfJWKKfgbBLTtjgL4sPiwVn4ph
DdRZVxCcR5QNITmhZi52psejF7VTqRUTQvEa3POtq9Mt6bbks0D8Ape0rjtZmFGt
MkraGJJZ8+U6zlsqc5R3en2RPvIhdR1nHH3CZ9FS3KklU7/WxneAH0KKxjL7Wl7s
tHeLiDGxUDvCkhCcLK8zIumYQYt9xmgUNEULeLJb5qU56Vzl+YKN6rrB1mH20V6D
TYRa6ng0GF4S4RK6MTQdHaFJ9Bos2rkcMRd6r6QdYlHXWiRTpbaOf+SQBWQWtOE+
ViAZUdhGvRGKkhrrMwsAp/ki+GqQItZsIaJMhMhc458QICcg2bFMmo0crKeN7fqU
WND/tXzwCdNSjv3kgXpl/AnEXlbhx5FeMIKl6KfP9yai8cq+GZXpBKQL+oRgTkBc
gBR44nKM0Rt1RrBWkeDf79dc/Sc9QjVYXgvLpefXbneHL4owctkYxHejanzsu0JY
rpwmEztVCuOViOzFHPyRFZydq9HC9H0uE6/UmCx/NtZT9h0Yko9TuUhAWO9WIWwx
ZRaYjblS+yNwMIRn8UwD0TlbkQ0q6PFL6bq1CoZqFsE4jVf8zxxu9KeRihujH3++
TDUUf2XHs6/fuuC/FdKEdoGuO2w30N0PW8knTDvT4hSWh04WyXm996h9QmvCQ7RZ
qFPRpUO1H9dxVPg4tzry0m+4EgYSJvrupdZmvF9zQodtBh2cqgicgnOavydFI+0W
c7Y+k2G3W1VEbRjMF2eMB90mjNZsDe5945RjWn9+Q3EWLEpD4n0uMD00pXV3D3IJ
VyA/gJksIvSslf0ikNriNZMaC90jOUUT/nz8cLO92YAD7A4XDrZZz735sO/fsTpQ
iyP5/rXykLnWFM86RbQfoctBD8tiME/iTvnOwLVkEkDOjCbJ6yE2g6ifxG0I1zvp
p/2oYR5rqfyb+lXPgkSqsvPMOlF2haex4o/n/6yXaZy9jORShOdFrXQ8L9tX17Ki
YDTeWuSD5mSqneILh1vCSzKgpPctgKOyDVoJXDn9zRqlrG7qaIQ7whdeLcxZxqwf
yZDiSKzFsBGoc7+fW/QT86rCwWhWQYLwx9kPqGi4mPFkr0Hi+l5IP87sFSjWiDc4
IqwLBEu4D+QxS2aWNQHCxXBzgZBjByuof/gyjbJrGNNZoewpm9V1LMKup1izhHzz
BiXHTOlNYenZGHxwPZWYQZLtbjDEC5/OfQH2bBled3hNz4PfcrISGhwO6k1f6LFS
LAClD98e44N/lVTqQg5JewJS2n/0d9bqkdaKTiCKrcq455MLdO5u5SNNke3t07Y4
+wXFlcewgc6icafAWDtmoan155ApbbMc1a3zDM7MJi6T8mPxUThtOAQzDyE4y09s
v3jRIgPbHLaxRfUL2zL9bXLf6iuwizXCW4Whzj9OovPmHCi5aYGecvJbWtRmsJOl
9QW91/KaAuLpgf/yJPgn/7DbDSbPT6ygyI+79l9Wz0usI2Hm42iLwBsvq5lzBqAY
oHhvlisNYAAKfRVRNw/p5R29Nehy+DwPaX53upDM2BKJEmM5nfs3IeWdj8I/2QyB
saz3KhFt8AACEdLOy8qU7wAEua/WX1PJ9N0L0DOvLJ1RXNRA1nmzWPMUbVq6QjDW
AprZvkI17GLDXwIe+CMiJxWW5IUqsm5XZy23PFC1isWDORNjqXK6FPwvZHhdmwmg
6OPvXxfQb1fenmWL9qFDcopn3g434Lmu1nPXTj7dbOCQOIZ1jSolUpaDiaaxHQ9y
eN811L0qgaY84jf5aQ2L/PN+q7CZZYdu3VwhgNoFgRuzm9q8AjwjEEpv1up2Pnsk
vGfOk/jo85oK9wBupq0sJ8cYoSwbQvy53KKBiBYUpIkqkTr9yQyfi73pV05r49Hz
sDGJ7QJapnp8h2vRLUj87iJWBHhgozugRUoxoYIuuQiTiqZPP1MCouDjVcSkGdlW
29OWLDRCnzFjNBecrtQ35pRjh6vtH0wETQxIjO1vsjijdlG4eaYZDYQyr69YVIOP
g/DXe7kE7XSl5Q/oPoheMQ7SlaAIXhr8lGg52yepFvS1XyEQDEzfsKCqd/ulIXdL
R6fPWvD7VkcesW3DXzFYtBQF4GMgeH2ut1VKfrMdKzVC8bEoeGyNaFwkVB8Uh4LD
po/8uPEOAvJlRbm2W+tmZN7ppVhM9NnzAgOsaDCO+l7+hgKnLmCkbleZjc9ePgyF
N0kUF/Tw79uStyB4lSzINO9OzNlMt0zww4eSc3bHQCnqFKf/dvdn4zmhP4ZUsfYC
lc1GH4cu3jJZ6B0b80Qx31A4H6MTE8+meIWmz1c2raORIj86QN8oM+8gm23uiCJo
VGgZdX6r7+BbYaTXXI98ku2n3SzA97iLHnEBSN4sEJaLTYW9Vix/InAYcvuGhQpO
kwOq3lVOiihw4exgwFLQr7HFMrFBDXJh6xhTT6puTzwJrXvDed5e0BVzquyjsN4V
ykhPgkBDmiLviP74/qYyBv8yJ7I8fVUayFhXZXCdgNl3egNSYc5q/ayjmyg9a9Dw
Q/gDI8mkIuxog8mfuUfk4xjOohYDnX/IW9pje4SO54gPnZfSton2fMbXr12FT91d
7bSPrCPMWOKEj6DRnY6pmB+dlap8dUCi/NAl92DY672ddG2LcbEzkoQmz/MXqrEV
HhE0ZH5PSivf3h0MliOSl634s2KP2KYpdy/MglZlicIhDRWfDioS3o8KGCAo8Q7P
OrPQ//NCrPOfmDdZ0/HYfw6cp4HqecVF4lEYmEuy3pyiCGLMPQXeHjpRm43QOChY
yd4nl21HLyVeqHMFh5SsQMYMyL+4wM75+/7HMb9jX87p7c1wQ9JBNDWWHl6mj96i
ZLegw9EczlV2mU3SI/EQ7enQ3idLEK2vT+lft1/VIygSs6KvAJKgXHZQPtRuZ4Ot
jnFEAJEeNqGIP1hbQcwzhYk62IaSJvUP+t5JH6brtneMDupmLZM0kKw+Ld3r0n0U
Z4sIZIL+5PRU4HMHxT1E5a5blU5kGy8YftvDumlg23zL7i8QXicGaDlwYy7fbN5N
SFuJxOY9CsI9d0/GS8PRk1nTBH+ic4kA7+xoOrYbs+YAig+rOo7f/IJ/k9PWcyoi
2oinm2+E+naalWyhbKerjvOQ5EGyrKu3Z0aA1r9i8w2CAETqk5yx8+te9L6IgUBo
bDKLsLK94qs5+etYT7FWqS7zzARKtBNyuPUYVwVOmf75iP4mNHoAf4QaJ32+j1d4
YhNk/iFyvjHMHPxg6MMczOiTx2+mJg6rXjvy4CGnjrZGtWoSHLmXjGIiiuoC3kZl
xg3EqgWW/Km8Ej0faItby6hXKYlYL2WiXDkeLL6q49gXf7uU3msjzc3HqfO98vYH
Z+j6m9tcdxr24HpfTNcpEaDKAuaNil6hO5bbkSxsNvXkaaCOpClTOSzBnBz/sYfg
LPt/cDIDRgMI+9yp1djMbJpfjKrjiQEKDoxM8YnKnfzF7xokMIsnjaqF3dZhkfRF
+y0TczFs6KbpP7WZ9STNRuAFP9cQUK1QhZzeKFHqmcs9qu502XfhAim+aqq5aWKR
6U4OY8fNqo8XhfV/vbHrDjJsnYK6t5cZ2Fay5/HvDAXhlcidKK58wNhEtlLzfLTO
Yq3HzzQw7C7/SvTZm87mYdIWWiG/5AVJ73oJF4WA029IVfPXFjUUerP3ENDGuLO2
jKeEnX8StQt8EANtf6jyRSeFp+SRrMSN8BQcNPi0p/rn/CKVT4nGgAjgP4zPH5yZ
rgTzU4qtjrdctLtC8szmsMc/SbwPmn9ZBQ77LlNg5PffS+otGyksqVNtRsGBHfOF
/5YCztiNvWvbgDaTDDaUqIPw/88Q1MlgJ/tYPAepUtcthxam8XdNnfZHrxpA/dR5
JoNeVJoEex1aZKyJ0zCYwR6w59UXT7WndIkaDJHpa+7I/qKQCHToJprLv5VIh0x1
sdhOFcUnZFN0cb86QhrksbiKRKns2dSM1hBzx3Xn6BrTkntMxfS38sBla4sGXIEu
TRuhDppDBvU2iD4XcoHSiYQCls+J0CXgNZTGPNG89K/ETJkiMpu8Ns/XDDf3aZ3+
KNauLGwMNazwuGc6Bu1Mzf1kNSFWPtLHLNcA39kQ+KZ9A5pBCyRLfI9crgVeb4IL
Yp9hKYRclX1Fe7oRsOjWiE4NaYe1lB5w/O4PIflKkQL/TwCJLS6Nz5zM3C/PtRYX
uorNjylxIR6EtIN3l4cPW/wV2/YqlQ7DuxNFVumaAQ58iVZAE+oMCVHtNuDUL+Kx
kpqkA4w30aFRY73vuEgnvg8PjPhTfBCoSGtEXOIezxQ+RqUwGHMC5oA4v0SXDXlv
4khOor5KtT0cTTTUwqIRBBO3e+1vwL84KQ+J0cW2YlXOUwXMKmAaIOxDEHwnl+Ow
0MPCMrfIeqKkxZU/YLxHiWs+++rPMxh99BDfn7eC3VkSMF5clEhC0aZLrkuEUZ3q
gfoInn1FO//CoEygZfEsDjNIoLvfLFekciinazp8BTwoVuMtudLYcmPfh6rufiAL
1Kr6BO4Zep/PGlhS5ao40YLINeF3TSsq7xSaTjgdOWYRBW1HxlKe2v+psnshM8hq
UTqRCRTw7DMDOqPWrDuwvmhGl73yCRyUh8nCqsnK83VBYp1OiSXKVlDiNevv8NEa
XAvpHrMlgjKdihV8Mv7tnceV7WfGrmHL2g2QmoM52RrK5yrp5rOBC8KbHsfOpZUm
yVnpUmZAbWIetxMScriyr2RNCOluE0xoLyjQRjFHBOH1miKZyMzzrtx3sKJZkZE7
M5oAksJ4RnokAo7kmcyvoTi1zGTq9EL4BuDgUtdRnFGWyOCx3KumzWuiWp/1+pvr
aY3nmOCeeEA/CUW0Z9pGQZvrysmfG7utNOtIxD7KkoUnDjd3Tb2k1C59a4xCZ3zy
OpW1XsE63piuu6I1k9PGKOBUWu7/tYexFN4u9BMz69/VpSVW8dtfYf3dapnVyw6D
AuNov629RGtzs2owYV5wAYSWS+safoJELjR6714UBvgeXVQdJXjlheNPYXYvT71Q
RJp6u2T0wrrjS1Jppm7iBz2Lut778SDGPPSVlgRtRzo4YbCBgt28DBcmb1M7Ucgh
K4tJqx1RmXSm6QgN3pjXzWSe0nuY7WJjkz05eNRswzcUA0qQf2xoZDX1wfRVsuh2
z4Q0d+wMmCsKzYpDjr3/NA/3XEav04vH0pqJcKVb8Qp0ps7dICSY1ZJoDqyCs0jl
XKlCkYhP7ja5flZ3SINjvuPdkcdCjL9K3BMTnbBgHIrUz7ngz8TEdLfEvj5ZN4RJ
NhfjbNHNF5s/+6fc10mWeA6zWCl5x26bjCHOx7oo8KMkbpP7o2mi6OeO+M9XjXxP
bB4eM07j25DzFxOZC1gfltprt5QZPHlImSrvZXe3ZJ7qB2eunYKFhqzgXo5Wie7x
JtiJvds4rA7Umr+G/JdgCgLwFG9PvILlj1XQ/QND0wm80lvGxz2UxDirpf4Vfw1g
oNGhlnYpyt+nmTpw9Ylmir7OO6g4fQD7U9PpEpaWFSemMA92sAWPEvVZiREmbeUC
XjPXV+zPK/XaBvwMbfKND0XKLKYieSPp/45JeiUjVjSm9aL1O3fmga0m9v3c8jRU
oABKl9X5KtXm6goPczqILWa3EfBWXSF24msPbAU5tNlFAQgLIukeMeMd65WhF9Ex
2Fb1YumTN5xO5q8sAflNI3ga2jk/LucldpTdAE+SyofBugCaFXHSXnom5ooF6vbb
fXz6GOPJ+pZafnHWyb2w2292bmTgGFP85k55+oMVYfQnjAGZ3YN0eevP/AVU3qWV
ixmqxzGC4+ln5dtgD9Li3Ov5Zt/zFrX8PIVJ6fWzIp5bGeznN7nHhRULfZEH2qqM
bjTPfrbacnolk7u4T9UlxU4X1Q5+rmsAfI0otNe9tjMcsa7JVaZeCBMKoMjm4VVW
P1HXKgB86BnROcK/MggS9mOdHl/lUm/sKn1xXyVEXv8UFHhLJCoWGIpxIOi6NYHr
QgFf3FBYYTLQ3ERMKCnFvX7+pvJgfoxBQzPfCW41IJ7hYvNrqPARzzgKtQntNRrt
gQlKTznPqj3mY/KNz+XqynQL+aleEm76aLByH+aOM+m9DQJj05F5lX6wdqiNGV75
j4GDAhlWUMUl7UiL0rXD+7izj1m38p5Sia4U2XvY/ovNtszLgixDSRn8qX1mgksj
IBTZiww/4IiAuMoBrwMipw2dTawq3a9189K5K2C0xcNP88Z0RZPUPPCu15lkOnYK
5IfjaM4nsqN71Tjc+zIqfcZwOmIJ3M/09yeNZRbhvccObVFs+RKRtBSHdWEl39nd
pTxyguBW7Sla8M6Af0/rvDEJOQ7HVFnW1Lgf32IXt5kJY4mZtIdhIGx95KbsCAec
puDZfn5z/E13m19RSCqidZUuFmwWk5yYmCeM8T8GSmF5J3ufXnPWFtgPyUt2gDWN
m/4hrJruexQATjBZkqyHZSvM9Cwfxaelh0odyDLktiZR1JLjJDYcdOHIlUvF6COl
7gHy4oK1Pq0LtBRlFQLr0K1sOnkQPG89t6t/hCzLTi54IB0CtmtWpuRm70DgORph
EbZF/Bqo1A58Zybh+A12vPNb3oKlF1Dx/prAKy8C9FqGG8UML7Ua3c/lj+fAhISe
tlHiiW82ulXp+e7fGyJ3720zJorlRjK+1fnqsEsVKVA7Q0pQ4r+2nw/Rq985FZfo
OnIYugXOcQYQO4x9AwnENTVmVhpIuTEtLsGJHM3VpgfROJeiInCIsgzOX/rRNgU8
c5l/RXZefkV30aLEvUuejGppbKkjYzy0HvALoK8AEXZDk0KLKZjYweCfk3rn9IPk
CCy4PtCuQ1ryX+A5s0q2UYjutXuc1RJIOUx5u92b7/3n9IR/1rIY0ApT3ywzN/GO
LMqHe7M4naUe1igj31dzyr5fiIm4CKP+obJM6bzNWLNQ4k6vyJ/nNq6DQSJHWjol
y/e0ooKdsCiOG2YnYIEtyfM4Tm0972ZC6ub214mcvxe1umGWLAnQuK7PwsVLEd6T
+tqcF+5a7eNS+Z6tGx28N42EfhOL9PvOrLFPNCNG5NBzh7/oWzraXXrU2e87kBLh
ow4dspqLv/jJEf68D5hifUgjd25HZyAHZF7k8x6+khJ3gzOQ7VGUmbrEhTOZ++KY
py2VGs8+SXoblGph+O3g6K+ZKUWnXviu+HHY4mR6oolu2egXOfOGgNik/oxqZpzM
UYQVkCEoymyEvbTlfK3w7JIBaOc86rWYOfiXBZXAYkmIjvh0gRnNMlAtG+X3Rmc6
OL3dGdoTDbvO0LjLSlM7p/NpTkj5jLYYeqmUBSOqVtG4TIl34QTzPWAvAoNWtlBK
GrkGBcq7wmU/zIXmD4vWyQ9eHOV8Y/Cfup+gGhaDQnd0JZEg4ne7NXqYTUkFCkP+
vypknK2+GxZweY2g1G3k4BBf5k8niAEkZKd2YzBB/nieZYy3qWAzqxCHd7nIXmX7
tcTktehdLCW/O/dyrkKYcIkbWrYKPX4ap20KMK8EwuhHkxlB5wBi5szfZjQ361V2
Oxx4qoXVKPcuRYuqeGPX9iPiqFlj+ith2QHf93xN4fGiiyT063SKO67wHgGIPJ8g
2b7ypcLPdyaJ61ihkfVcn1bCPzqGt5Qek285rSwfB3HRJMzcOD4e8epnFrO8RCF3
3Qa+u8Iv84alCp0yNDKzOQkn8XExMLTkwlWHxlTfq103YUoYGIfIQyOHKxRpNFTV
9wZW/GCkIxAsAg4o4ECfMJqnhdCycuJa3MtyrUKQdVJEhHwb1Zyc69BgmUtAns2/
Qms1ZmiqA+rWUWZF1925CR7JJ08CWPKparL+7ysCe6a3li7d8AFaSD3iGGNYOwOj
StR5ahjh4xvPf7A2/j5MTV4uJ40m1KkG9QcGMwDqQkIgmH7T/WIzNNcrYi3OfUrh
3uRTNNFTqpml4gYmyq8Me2ifo9hV+HLgn1GHhXG0CwGm/nfTKu7ic6sC/pIbvRoQ
L51LCoKiYsi4LD5h2XvW9i39+f2UbG/AFhg1qK6bAOHjffPFYknOBeuwnKsAL//M
kDxgeRoTLOXJ6MluPLBC0m/GA7FsLfLm7Xgc9uGN4kAdXIbbHK7TgvDlXz3fIAni
x0mUxC86Q6jV5uaou3HUqKjLKR2V1N0i2mLmge9mIPiZP/nhzv1pbhYQ38UUkjxl
6Zh2ecJQejm6p1QHdkgaoNa17Fd2ZGGktqRDHF4Z1Va3TMiQD/PCkTU1vfyWIZO8
7tHtQd9kTup0z+6BhIFpZFPe8hjeOHF+w3mHV6C4Z5etfNgOFv+RENYD0GFs0UE0
0QKJAyD6pPqWejQqUZqsmwiWECy/3q1icSTjvQUi20iFbcclvPIayoREFNQ73PiA
xKFrDr6j6id7OXdV3CMjeZo1n1lMpZ7sxfAFyY15PcFkVgNgvHEjzCey1284DEKd
Edrcgl6iCHEtY0D0B2oqGcbsIwROeVj6srBX9lVMzMX0n+8zkWZxRAURs0RhvECE
Z2OBL5dKkfccwcb5VDWXBGw6F3QA7ERwiSsVbPidgUim76DTVc/cMUA5YqRtI4p5
WpCfmipaFh6YXjxPEC2B0HYLsJVdQOSzfHcI9oyT1wPENvNnI0WcnOuCvJSFPRc1
CeffeuHP7qhMF47h+Ee3rl48v0uitwYkmXXFPDItRdb+zuiki+FjU331JntJaYAs
NlxMhHnDuqJXsNUPm+vOtD8xbGwQ/h42DHZlvA1upfUAki0Unb1u4QfU41m47xc+
iSBEHcgJ8ysTwSDo4+xUzagWMaqU18uOVIjOBHYef/+Lmka7a8mU7eLSrXMmtsuH
OvafYL5CTUgTmK+DagVU2ga5XKe0b0SEwrr0vqh+JHkeWoD9DkbLp3sBMEuw40aE
NkBkJzuaTync2/DFYl7jDSWHGF+WCoHTr05gsC6RR9f8m1cpT3LSUPXGFJok0dkB
XbYDDuIUD0hL2nFMKg0gmzwwwbU7tV3zWYVebVcneNs+YhqlfLQyWC+XTYHDqM7a
KtlT3fqn/X33e59wbwMJKyHqZqc8tS0SuMjhg7Ye0RQHU7nrgrBbslotkKqCbEg5
80MCsdypkegTYQjcHUSk1lgt+Oi3qs91PE64LorqKLpsKTkvU0AXO6Goi4csGj21
O/JZlkLb4wxkG7pFhVFytRHX1YRCX6RtlpH4LeBB1Oq4grdVOCB9z+cknJDEKhpH
8SMDC8dtMOupQrJtLqMHrKFAbmuiFHdvpSC9TYAGObNiMfach6+prFnClZlIMDU7
P3NdXgeuMyuLE/DYvIbDrvgDrNYa9SZUZpHqOuTOrL9zSebJa9JAOgrB5lilIBE/
6AkP9boceDApS0yPRF3geFCR+CK1OPHM+jbYCP2fHSALo4VzenkH/wprUzIt3R2P
ZHYanp7ebMT61CteKbTboDxSUgNN4LrRnKI13nQZK0XxbVDklYaJ+lw/XIYDVe+8
et1yegE33XqzROg3b+pQCIrQaUkD03a3OdVDm6qUFw3DfYcrB4eMXZYiQJoSET1X
hjF+mfCFjRj5OW674xuUYIBd/MYE3EY/a3UNQXGXvhoIZ0O33Qo6EOfAMItV1Y8T
DQYWHO9gsRRjDPL1XklGgzgRiJeX4ZsJh+QQYk3cUfYY3ADLGNEnXEDWqDvKGfk0
Ew/XLQWpC2lCn9qhkJ1kixWymuMi7M6/yrTYvn1rULrWskoAa5pUY812pSZ50xxg
f8G5jfFLb3VWL9NI+hNwT2ZNz5Lu2oa6aqs9738qGNOZEtGKIHBJRK65mdKQ+QCI
Sx34ZBjli4FBLzD4c9oAIIBMLVdxbUezuEcTM1kEU+1u+eNs3p6EAIyv/JJhjOGd
Ps0/OvWYlvYdfUiUhInrAhpI/3F/twqa1FkHbQQM9F263QLecYrCzWYduQtb9SyA
XxI5kIRDpMtQRBDDI4M9I7mG5VbtFHky8BAhsX0OpC4L3cPzKYrhgx9CkrE8lLB1
5stnZnAHWRTDHzK9kKh7nxx6udRFtrca3z25f0wXTV4mjjGtOtbDjSE9htfGoH4k
hoxqnhGDibL7cSkayv5BitOdy7cQ+OehDGN45lilpRpUPH5nAoRUXvPCwhdovGMZ
wNCKyBn7iuRmHyqaYu56m2IrBfVjuW0aLrm0FSED08KIqE3syqqGBaMsbArfauJf
gfSCGIjr2+qWXlT0fg/i52v9n24Umaih0fIXDYp0K/nhiTF0ayn9aNCRwaMDk4wE
BkbACwT+ohhWJNIWUuffI+XikZnbfuZoa2X6YS8OyHiOGJGjFo+w0uzxtl/acAWr
m+g7hAAQJtxBXOWmuEgV3UqYimw9mVfM6R5I7k6lMTPL9Llj8kMxwwyVypEJ8PtW
Ntfs5v/sViW4TnpfNXtq/8yJRbT/sKizs7EJPYBVElIerkAmcnms0Ryvp9TDoAFa
4GHbSNzFYVfBgmMIsDv80EiywVFq+nG7rLYr6+gNi/ul9CRdwck8j0QZCv8Lmytq
1TGMt0qPIrGs/fbMwIPHJtq89zr0ShmR1hF7RYPik9Q4iHUXg93x9PbXZErPo6f0
vvtrZ4HOrUNta8eGmQioseQgWpPh+fEHHx9uow7tPK4FREy2hl3+rP4znMN3gVvl
sh5+cBVoqsv8oww5A1LkfTtQEMEVvyRT1186EbGpye79SkdIt1tagSbhHEZhHbGS
XdntmV/mpFft2OBiMXsZiIUDs4EckKa2V7D5EY38VOdIrPh751RaZ1h+BkT9mSJL
GUWW+vzptuZ6Hqtp2udycrbG95vSJGXqXGpq8UVPWsgW5R65re757lyS+JrQ3LdL
9CRjeCte7FkiUdi9Uy/Iq6caR+sBfwUk5n7Bqjki6h0hVkWpJS5xvcsz6Ha8IoTL
UutDy92lka/bLP7Ex3lqm6bb/b2JVB14epvrfksO0cd1p9mUN5Gdm8VYHJPozhcI
jGG3shGjl9ah47m1U2pLPiiBLmeQjnzEXPV+EMrGGqnN+vTRMJGM+JE1/ZfmSMWa
WrcI3+YzyDtW+SG4I2iohIM74BAUtqVDBq8fbFuwGk2ppTvppohK8oxTQgn+x+Q4
8jIii3NR91PkYDQptuMpKXZRTKseQiKz6LZ+NQnPFHn9CHdoJYU7oaj9ZjgxqZnx
X1CzbwsjQkQMC8CMfYSePYKjXqGjYkci9dkNmUeJrXcOcfZGzgifjvETsmU5mM95
JTnCE5dpfHA2PxEM6PI/FjL77DJHpmj/owQh1FRipLJ5jfJSGZoi/rp7ZO6zWnTW
rRWRNJMFEwZn1tdNe0mb+mKIffV6Dlx1L0EudfQpoV6GBUvSLWQGdMPVyRUNhZh0
dA6seB06qsNj8dS3Hv1mJ4nsJ75hshsPkB0wdbNtFipviqIjmwWM0BHJSbA6RqNr
7bZfWhUd7h0XUuOGOnnOGG+UTziIVClVI4X6w1JofOWg8exsomghwFejLYEfVxb2
Z+dPy6KCoSbfUVO4hxv1H6JDaWDzTCWRffVuJqo6eddkED2o2+Al4DFfeJK8p7Sr
FvlNjr+3sJ5AycHYAiCn/eRJGsmTSW//Tl5XGnK+JsxFmog+NZq1QYREJYHGkkc6
nrta4mPJxWYmIgQOcWsSaKsgIZsv3X1xCMg4XkInbusNywCyIygcq0sGKVAs7WNO
ha8PASCJ/2/BsDDTrKFDpY8rhfj6Xiz8lc5X1GzmYxOyIk7bm7H3s3M4hMDC2d/b
VHvQI2aeFyKukdcpqGvvwGePbQBF4X+8rxNmFkAI+Xt9iAFxSBDb7EaZGenFDXC1
1EF24jvrX5s4hcKlgnL1zyNna5JQ7ZJbqkm/Uhh+svo9Q8zcqRa9rBVPdQvxRQPG
m9uQ9zbjB0Jx4O6ZFuIDnU+9lUM4sPWjO5OZ5AVec+wIjhMQ4e1RCII1bDCMc+ed
EZ+TYdVVcqFzuy79zAHHuCOXLvL5dBPVh6sgg5YJtfoYp9W6Kr+MhoiuO71WK+NM
CRZ78baon7tAgOELXeeWrS2UNOISFq/myHhr0J43aWLFFCbSdt8QbWwixVq9vKGV
1yPPUiLwXOgZE5LmYb+6h1lOm64ooI3arKET+epgEncggMS7Q/XAuej5ri8bzS2C
F7PyC6TMNizcIv4VzSA6jinhGaYPeNDkikzF2PxVxkXINeVG4l2frWztP0f/WoBn
bq4WZpafoc8SsJFInZRwKuWCXFVjJ8HKlOOwrrbysgWOoatPex5h83ndQqCyCRnN
WlALuxZW8DLFMBs9ukQ643u6rif3/q2Bnquh5aD0kAJX+8LKqMGaAA07NmHNhAwk
lvzdDzOYm0zHTJ7YVL3H1BPTf/yv+XtDLeWFHNW4WNAdFf+Jm6gvyVneJVxgXaXj
NwUvJI4yZhHPjeS03wJQCT7lDiP7LJ6lxmJO8m/adyXVapMWqUU7UABTjk/xLfrp
+U3eOrENLDziDob3EhGS2r3gwJ12p3O4Vo3VYju4TLYPno2m47YcpmcoXqHxhiSq
2naLLcYNRNUUQv6vzu6hXHplfvrT+RyuiTLpjWDHttbbA7yFvbgbnG9Bfdc91XYG
J8FopYCrVFy+IXDQwow109Q95KRGT/QVvRMtkd2UN2GKOxo+LhdA4LwUIxfBfa6u
11fqG4/8IJr0TITrJkiwq4u4y3b59pWG2TjoPO+HXa0ioGfgwFEaato7W0Jreegz
dPDFXaxYCZo1AU+c/kVMWaki54A5XL5irIXcFmci0MsXapgSFPQ2/wK6kbVGqlRr
yXPbcNzC8B1T0B5uQ/ifVLNWLfRw2SCDRo2ku8AIJt6QDBP1aGMbhbPp74q3ch8f
QU22H2zX7vNbFrJv5iMc82dE468MJ4rlPndJ7vMrC/pSiHnDH6DYWAAXyAMCDqIW
Fcrb5tGoQUUbWFRT77xRfR2zz4+T6lsgFi80gO34tB7xDdaQZKO/A+hsRYlryeg9
aiHSEVm1lEpSCyuCyml9i9VujuBKMq8UkbkLznTyN7L0HIgOJ2MP+43ZDKRKbw5m
r0Qvt6PniBmo5XQpmS5nD5QyAIe3NqOLBbk+HDN1MeMq2J6dcgDiF9wNv+k9sDeu
5XGwc4xFqMdPx/PpaZVm1dCFcibOhADDqxmUYVLPh21uKNPRnJZYqUpiUMlrrB8v
S4/iFLoqN+jkhbO8ozaYVlwl3ku9LhNKTjzAjEeByAVNSh8mGnT6UAHOAiHB4MkF
+gYCGYgGx6GFBxJ0rA0wfSLDjPhQneMO0ympWJ1blBjBHEF8hxRrUHO4MRcXz44t
BupDlmw2kWVDdpTagap5PFFQjFNDRt7rUwOoNe/KZzc1k8G0ItRh/5Yl80UzvYmY
bVmYN37M27ZNECTdsdynWFSUFa5+MXR9jhviGAixFnZedtT6LioT1d4P0Pi2655M
xheofbnJ3dgfMk7Kw0ILW8nDTm17VW5tmf9VjBuhixqV68+CVQFuTU7S80jOJsG8
wIVPR4raZsrYjek1ADVMH+13DnYq0NAOTb7EJVq1OP3JuqfblTtklVaubvBqn7f7
Xuym4uuOLD2J/g0P7aqiMBvO5kyAqERkhGKY65eEsJmRGQ7ixczjefptz88GZltv
ZaJiKd3Nx6MxcFQUdZu8fB2SIoWC2JK8/GAW9MmeDYhm40oBFq4Gf65FLk5AmpIg
pzgKwpKCFOg2zBFxDYxBFGjGuKIVDsY2rVGP5YmK2uUAbNsHuKqK20YrkVXNU/O/
zOEsOUv4rF3z27cKD88FlUa8PwTDdBYbhcX4DopfD6CTPQfj2FOZOL5FjQNmWtxe
h8YLL4fHD2REUyY4mfRqAYSaZXCM4gd3zWCCsErwjbrQ0yc0C8rNwAVzaCJr30M9
TRzS+0+HVb4u3s+jbOk5UNWbs+Rf8kI9dd7S0DefgAUcHTU+rFX38plt3XNbi8cj
t0yUMi8SrTaqU+946Q0cYLBG1zmAN/QfWYkHrZl0vWymkn8Xg3Ga4Dfbz4G5JSgW
alab3qVbamm8Nt5QhYeS9bDF8AavAyK3VBE8WSFBpVwwRZYt3Grk5oiR1MiBP6M3
uYDT++pHJOGEOsdoEYGdLyR/ig4crulW5Kuehh+LOWRvNwpWZlZaZkxAq9QVrGOX
jnmen9aSpPQZHuo7IX5TSE1rx0uVukUMEHDJ92iA8qpxn2DuwSwDtEtVgsSKO4GM
BUz/k86JNvE1dBi5nn5OkANzEXKymXpSRT56ztabuk3WVwgRa9aywKGGu+3zoYqY
GUjiLMmINdzmv7k3yNXbYF/nqQkt9X6j7yXd1Xe97A6ojAQD/LReSyz2ZaRCFqXQ
qicAUsuH+1iwxf9aHNWEuhcVb0uTyVvyQta63XF31B9Z/b17c7Vgl8TQUtMfGc+e
ILRHoE0aWtl6LOjWTXP6zSVMfXVcGA7os+zt8nw7szoMa3tWqi2Z5AZKvc0py/1u
3Irhqz97KVzYbPpOE3NB6nyWBM6+K1A332R/LuAUc9aQ1+jX3EV0D2NAuawLhZ6O
Mh9gsnx6tY6hkSnnxVXw5r9pW0F7wi0d81Z8w0xbkd59LRImAQ7DO1b3SzvBJN6Z
9UBKIhbGT79kQqhgB2/EkjB8U+Ew8eZnQe0DQbsVSejTz/akoT7HmacPWXgx067W
QTZjTANt86cY6hSgPRxxSPuMaaMokbz8TtL+EDK/BPGWCBkFUpKfY+KyQhVV6riI
kMGXf6rpXjWkp5sye1Vy3AAq5u8b/50gGBU4Aj+X+O7bdrdwv5GoPS5wYPRfa8yN
7ayLcSSqGzIzZsXQoqJtkwrExcsGo0WSx6jffjtdK3M6bY80TVkD5qustiF+zK52
q0nwMPxxR48iS1hwMCNyYM1DlStQ9NFJk7sd4anryvDSkdJOROzLpo50ebiQdlRK
ZmP1VdQFbB2VTpjjuxCvD7/3CWStkQ4ISrUDIK12a5JC6ayPmeMF3WjTByZDi9bf
exok814cA4m0rAId6fbHtchrmcOt8+LxuqHWV3CuQHaBRMxXMg0fWiYtmeZ5HTj7
Ew/VoVU0AtqrJvxq0yz1739gR6kdxhj5WW3dCSG5KHnVS4gfzf/N74CeGI3rK385
kY3qS1e81jqoK80ObXYGAR/IDJq91hgKDqP5mP+VqdjVL1MPiylNlsZwLVcZa6ky
r94ipDHm/tMfIg47n/bqnqykevSfLpK2apkNdEj9iBFwvzjhJBbf3CGVFN8fn7cy
0ElJGY1t5o6elyJSckCFmXnLa8IvqeXSHATzGqi9UugzXm9wvE4ksH/rWbx50r/G
R/bCvV/g2/vNdjKmzUwGp3R0YO94/soPkk+uFaprxizP37prFv9vipbeKSxWKJMT
AHeW5qBYKKQmADDGgZ6nx7t31XH7pTtXSlW7znskfupGovHaV2D1FfYClq6p4ZI4
CAsKbUfw5SbhPBbdD8yM47ai+mwzIpwmXVMFfIETsQ7y7+YvwSpSsAGxNIJ33frE
JZc0pp2uOxvDqhqhbUEo9yyd5yaiGtf0eMjSci4ifst5JUAcfWpR29OS4ycwc3rv
GNmFXHi3/uT3loCMgNsCjlBYIamzBWaRDypw0Bq8QWiYyvhJNLMj30wlKI7JSGYv
FAZrTJEHgjrFSiRBatmOfjAxRCCutgNrp98yTrQoj3GxtN32zqzDAAc9RRoUMotq
GVYp5niqvoqGPceFCZUixX13jqtUgVnmK+S9ER9/aTVQDzmqOjjSMeTEo6Ybi62M
+V3rn0LYz34qoEF3HolRbsUzMCMrZH3/venOKHBv5Vv+1dvKxNI2X9dGPtw6uHRw
0uJjJy0RlsYy/Kz6ApNBxfcJ0E2XNzpMzea4VYFUsJJzA5u1PijZviAmu9MbpMBe
zys44sgGctWfHTfuGgzJd8CANFvha+cz+C+l0+4Z2ECQ46GrjMw8XaXzbqEzbDit
xMgIBXx7ThWdIP6VEUNu2ZqRO8wpjAqfP3aqHzNy8dmr+1rnWK+fTuy0U/g+s8AN
ESkH6EeROjyxyawqbbKVIzVvgSY8A5pQEiKnkIo+mQK+9urZqWeCWZRqfY2ZJXSe
GB8eLhIPoJY4ADk9uIX/taJnigqCort6ozYQlSCdCTkNSIwocXzverrqg0lROkze
f95yc7VCzgai8KOubrWnMXB6GPqHy/norBO78ZLZwRug5DRBOwSiOvE2+LACRo4F
lvsLEVC/pfGz5rbfEbeJrJ/NPHMbm66N3gsaMYvRdJW1lH1L/YIgkVlFxkhx4euK
HXPiZB3RKfqAKnBrPj4/M4K9HOy4dwP/gSFv462RoP+Zkk6KqaLIvwOhqFcrntUP
xgFHy5Sip5YeBWZjM3ZcW1nqivUWrFOGQY4I2IF3juXXEHkytZ78HQ0oWM4xu787
ep2nS9YBM2gISSlyON+GtvG0wF1axxqMJSm4p84K4ooCwWdZM8TiQ9QUf7Sq1YSg
ZpxjfKkqxTsI09Ucc/mJrg6yeGGC84GgVoDq7zJEvVVl5W6gwgStD8XvZMgU6Cak
bwQfSdblXLaIvaMr9AJlhvc/vF4IeYoBrJAbv3HXl/L/VSi86UhkkUNzo/0UdlfA
OLUtxjCLlqUAVx1PeGK3eLKgy046VHC2M26FHyK4Hl5phzM80KbXBK1RhNE7aN2+
kqPqxWLmbT5lE32+CcXtsjNTlYuEmzWX3tZzjAsPbbt4IFx5Qkj6Y0I734U6ad1v
G31MsSl+YuEnpZmlF5thkVisH2sqBxFILGGDseM8JG+6Zd89+/3ZaN5BiFzQYPWW
ORF+qlaGxcgKMWBGkETS7d5LkHlLmSOGix7lRHLhp8e2VJkwVfeK3RGP2p55hCGn
xm9A9XclsMazHvlba/pPZKt7YJoFSHQQjpCKv0gZ4jWeo/dY9ElpvK9VvBUcGa/J
iVKpSUCnDdrHesQ/abPcItFzFwIx+oYl2Q7wLo/yj5kikQ66GNpVYkTfVOEb/tep
74Rs/j5aJr911FHsicX8owvJJdJfr1XZwGE8sIvPwvsPW6pXwi7oY0krlFiG5XSf
OE0GWmKSqCZ0zk4zRLfat0f5b2yDJ+Qa2+wqwYf3ZmeOcgZKHdGwj5O1qzFXOcFO
tSNDeidAGu7XxGJEws0Ec/TqCrzVNqAVmQdtzRL2yejUFNOqxSrxDnh0c5tx67Nu
u4BG1oCKURDNxAxuUeunpB2rbeZp1k+KvAuGSfiCWpJs4TtujAwJfdjneRJczsac
093OEy/vAmkyPiEu0B+A/EKNAXj9SR+DKb92JlnRXrvumOpJ0XDpBGQVmCyJinTz
mEof58hdsKTW/YyyoMlYbrF12xHJtmMyc4eSKifQMXmNi765k8pWg3olSSm2FM8g
yb+N8VrMX6saoLZRNYiONZckT8n3Iesn4Rgrf/o1OSt8YbJm6vje8BqYJVrx5/Or
OnJ/2/EzCxK4fBacl4G6s8oLZrSNr7DaVcCfmZfkNkAbe9Mp4FqHG6IQU8yUv5Xr
7WLVFULfJ5IN/ZZJrLFefF795XemjmsvTfz0Inz50jl7eUVlapDg8BZK/p4QDcTA
6VjDVfibe+W+TPh+bCrttMw1ocsrpJD4acD2ffit9A+Z3w6pFPdFFtbxkcmHI/01
VG0VjHCbj/ZOcYcItt/LK/b6b76EtJlK9CoxndPYMoMHrmMzyaOATuB5oJ8xwI1S
4xBH6oZc7rdtVLzSD7crUNkR3/Q8wiI9XGx4Zxu9dgW8XX5oQvK0a87hgCGFGaE4
ZM9/BnLmrNSMzb900z0Jppp8iuVdemDISd9xdNNjWiWKq+Ey/mFswOfJ9kjBEKrm
qLpxwokYlnX4QexO1bklJrF3WQWMPy5SWsuJFGOfW+Ar+SBE4/+KT0BRL/TAQa7M
xuoWRRUHVHMcepVs5mikUmDLFmtJeSM0vfYZ0qRSzZRSUonATiNnhujf/DRp5fmf
fegoPtASozQVhL8v0CUoIbJzQJ1V1WO8TKJTYgwEq762im02VYR6unupHychjxVu
mX9CN8pMvKCHGSLqBtnK+cmYdYGPijIRwm4fCWI4oWhBbEfKRe6ld84N1ri6Ibpa
t5uC+yKwaoMJUKFdYJarLQhXnsRx/GcEE6k+7rv8FpkV0qtGN38PO6hDVbBwigBw
mI+Os+boavxSoRNpEXAxsM6vYLBUJldg3gQb+Jw68ehx9M/UpyENePAQ9ft0CeXL
mzdMg+4zTK5wFRrKM6gJQvolyELUUIhEXl65zeYMM5fMh6Ddd13ytRLUPCBKB3if
sKoD4MY2jJCSYfHApt5fPnwbYm/CvqXsJyMB8QNce2jv+3rftcILrBCMiveQVViJ
VCDhWqM6i+V/aLcwyvNPrMlfGnW3Lsa0QMQ6nUbEZbgx7iank69rB70Thm9m3rmF
RA2Y8T2itnK+yuEyBoYCjd7wtqxTiSQqUbvP+DZ11HLgS9Pfknv7AL31LwF1En/H
hHJSU9ODDX+gTkAqjtx3Jg4AejYz2oSnNTGk+zMmP2h5QKvepaZ+LlxHauNXnXtL
wrnx+oE2tNmwfrQKRre5B+TPoXNoXRmuuVTC/hXRK13eI3YiaIX0yy5+prlk6Mxu
c47Ufp1PtdbRh39RRNGVaudYuQC/l1/l8fc+0c8di6KbRXJGVJbpMFlc4BkFkBFD
CxrIT9GrbkEQFZpinoNx1BydeIDSNOjoebh5wzHEsMsqy916iO1Ec57dsUDnpjYG
U4Rqu+kwFx8NyUb86x+1wcQhZX8qFpVa16tgiyXBbpcYs9eIj/53wuEh4UJYaswY
yhRsN7d/Z3vVJPTGpGyWh9IiFF4Ff/tvZLPAsHdS7KVkyIB9DWKRFUFGjZt+KwvG
xe1Nl0LeFFPEipY94HDjnFWMXGRF32PWQ8qNik/4PyQS0eIb917+pcq2bRQVdPve
nhJwog875KpSjuV3Jl0u2hg0wrR7JZE01HUF2YnUUZs5wCelvYuRtQBL8RQeJ4ix
GZcnGl9cqmLdVbEYmfDk566qyEyk+LTwOEnCudtAwNtf2u7nMUsoAjcNtGlYLTX3
FGIkbwcQLPz/IEzp72OPxQb8CIwdILYP387SFUSi1mrZys2T+l7W+RzOB5+eqW2V
5h/s6T7qzoHDKzV3c3PBc0f91raw1LXvOEvy9UGhvY6cynHAJ45jZzjX6V/nG+Vk
DQmLduYXfqEdIVcP5FU13MuCHOdhV54xUG1ijfpul+zo49pIno93ScUmcfwUCKy7
8/aIDgJE3WaItIvCATCjfyUqSwPS2RUQleN2whvvdAJZzOnVDf2YZfoxxxmdfzlP
zxWW3uCO8hk8x1PtBJ14j13Sk/UzvNCrvtWUzwSZYZYA7JTr7nkIQKzwQMMmubXr
qG0VvLMCEhuu+WN49qUu3SFn6uu27adUu3TzIml3rgIgRtYDiM6J4/1xXhcL/KUi
zeYHCGqCHy10/Gt6AcQWDhvSmwo55MRTn1GxIT+VbuV/RgIJpjU7exKTV1YlqIxg
8Set1GMhFqDfb0cibErkuF5u9LzGsxdt6e4W6PmKprqnF6CqMkGnAlGhDQWWFyDy
s5/jDrAm+JFvRPq7kglnd5Ak2uMEDTH98R1Bk+ZCr1HosbKLR4mD2rw6ZczdQK06
oS3KZKOO9/vDyHiClhoqgQjJNw2aQzVPc2qnvAZJGenhcKi+5iM+0Iae2r0yaLkq
53Ys/x0oS73rDE4d0LatzxVxtBnsOG/qfbVOz9aTbfacXYffH2tlVpCdNsE3O9fw
NcmWOj9F4opK1D6zOX00bbErUg/I+t9IfLI6vIfbyK7QYrmTEz0LTfknS/vZEDUW
tp2KBCqhrMLY4cGyWjEjVBlOPkaCoE16SricJQLqiYigNkpsLkrXcrnTzE+SppXo
wRltw49fATyDNTfW1ElQDmKkLf+EejVWpCDzXmTEBy6H93TzxZ3OPQwW8+4Y8Jx4
bKd0pQNxb5+jd1P5EVrDlPd0aq6XwFxC9SFWkyS4l0Ivgvao9XGRsTG5XtZSawL3
pOLXTeugrrvpEjchqqY7dHN3n/cNwPN5vU35YnELRHnJX/oq6kse7krL5nQXxoum
PjyeklYm26UsKtbMDsp34habKkdSDaIMfE+xSXmjTq9mtjkNT2yzsZgvKScqf2Ow
Rj2HdSo7u8xucvRxuWbTISJpCPW5TlZA5Cs2J0y9feF8ovg6XP0myHbRyd9jYO3H
C1SD8kxPkolHfL/WjHgxiKuuaJguuzgCe6Lt4XVuRWRHbCg4TgOxjdsnrhwdMSNk
dOe/NFJ3ZIqk1RIsoSLVRlH0F3v+95+5dW3vxHN9ib3ApYEA2zFiZ/a2NXMwE+Ai
7vwh84Wrv5amSdENSScIEWw1CYylGQvQgHlEVhECYehAWzdFiwfynWfTxTxtKcxC
0zVFTtPOxuJAA/9CUJAUqJPpmYpza9yYVLEdPSO1QpU7A2j0qYOfUADRArcVQz01
cyNuzuLtNKv+ORehRb2HQR/ECtlaU8laSs0HjqrXP8x0+zl2kCgUgrxHG7cDgMOr
REYpQOt7FGeGKbhDm+UCBqYILvWgTxdq9YwNyFR4Uvtra+oMDxF6FapMSPhFhALf
nSESR86vD11kdpsPMmwl0vrlwHd9KuIbRTpSKTeTXHHz3lC0iAE8hpmqMQRTXAB+
EM8U3e435te8Ga5GnqWXmr4PM8Hju+yCSOUf6H4tNa6BAnFDARXNG9hEi5X91e20
grpNQ+RdJSyqJ1H1+msfQplS4GIClmkRAXD4No/5Fp4bQQAvivaDcFaXCXhWUUO9
lrZU2MmK2eeApSBg02yqfsCMTO+j8sgf5u+pZ5gnj+gBbe9k3TpYGjlShN/xN8rD
GsEbiQxl0wHfTVtw8Mui0TXcIaPJf98DLmEQWWac57FpYNpYqXylfzqsjzHn+pqp
NKMYoyWEmhTao/xoD5Ut5vsmdCa26habrZ/Ce7k0JEsu9HfY/zyiEeOgQ3rlDqaR
XAz+WeBXynB8uhq/EISHBCf1AatPHz5rlejQaW7LCLrN7D9vaUQVHPtKIW9OSveI
X85Sxq0Ca4Hv8spY7pvHd6VRoKe/EfclvsU6ptKWykxHEc5Z3UO9W/QPWb8LTzs9
hzJidOZinfKISDkud3qO8PXDK6UCw+rbhA5s50zHE720USg5KwyxePQPDJKlf8LQ
1EhmdZZ3AiaMuL6qSxnTUCxj+reddlqvrN3sQoyX2Z3dh32XVwG2xZTXJJQ8bSha
EEohLKE+YFsD9EiWA8rAGI84taYYazIRkq2YESgg4JAaiYSXBbxGwIfAN9RFNes8
hyppLwQmlWuyNZ93RI0OabXhXKz0yWV4KBoEX9128AJykCb3vBLnhTAnwp6WCIv/
l7D9pGH9HcH0PggLI+TrzdMeysORWRXiFOY+alJkMJYRnKKZkhmHjelPu7lYeo0k
VUsUZh+qJ4m5Skg3OP/Mlu2BlTk9Q4boULtyB3l5XVJMMIMKHye+6SicfB4KlRZ9
Msm1e9yzXSydjO/Mt5IsJJgoO1Nk6pqJmPMdkX/lZEDJI9bqGfULC+OpDDuFMxB0
hbzlyO9ChMsIjzTLpXBezDiX/xNPz12usJ8nie8icEuaSxyKp5+EFSKlzlx2wnp1
ThH8dy/T8FQtG3n/ouNSAA29ZvWK2KmqWhvIfkhezdGu0R4rxcNTL+BRtbagpQde
7/qD81Ix4LL+sWektB5eeDbxNDcozALnULYf8unFtjbAt6VOdvtFrOE++F1Hm6Aw
hCDEEZnmNbo+wbjPNlAi0NLzNB5tgbFy4hm8NV+BzZC0BpmGV5sAPFpP/eSMJp07
pVF8+M5aoub9XtIeidFoOSZ7ZOQFyHejVlmf4KWrlsAwbimVJF7vk0LmTos4l1ph
aJ6rb9Mtja1e7ido+dVKlpX36UNeBrmcnd8e8AFAfrQxz4C2DZEkenkdyc3GLykw
yU4xc49fbxPdLCsY4slGh+OCPCZ/LCeX2lYNN3URfu3osCCB35NL1/lBCD9m/Xt2
VTs3Udn8ybHgiMnJppcJTXUpN7c0OBRNprQnttFZ7pL6m3vzhjVwvYqHe358+taI
Lt6g5UwEE8OdX9CQMAxmt5udTpDWZAsowUBQOtTdmyV57G3jTT1IE8e465XVMjUq
JUMEvVbO6MQst1dkVvdz8Xp3+4CrRyTxLFlBgoqpkSDPqr9cqMzjHECLWLkP8IGh
4XaSYs28tHIRw6PppCn++OmpJ2C6FJHZ+GKhg8DpthRcfdFERonEXkW4mteUHXv4
4kCfxZhSgbYPAFH6UTuM0D1lDjfKATgz+iMrsaPKHlwN5qAUpKtxN3o5QPJYSaGg
fWalhC72++8Y+vD69x1pZuy5eiwd4TmE5iou2YSYhwBnvrbnccobXyrpt1ZgF5Qy
fG97Z4Lvyy9Jp2lvMnjRKMPrDBszQ0A95r+EiJHQzSKJJpAZgFyhdLgU0IkmA3Jz
jC97C6YHL1ARep/qXdbsRweRlkiw8CyxzeXRgWT/EhmAmOdYqYcmeeYWi4SUA27G
opZQaiT1YJ6o1yMQ/+iUwWeUyQBTAUDSEeN6rTGzaf1uhJTLm6QN7qHLmEvl+2E3
DIEtdPyoiv0ZXSaXxmLcwN032TtNOGW4seWEBczp+PwIQo7y5Rql4ZNYqsS5orju
9SDk56CjGtNeeTKMpno6Io/U2A2WzVH2hndDRw34rTtySyzfFP/u+rO523j2sYiq
FF9XjoaHxTTs3HBDMSg7PbfZy0EP6g0yX2CChXRfsqNRHRs2oZtZyfmSAYtjUWpY
BWw2kA3Px8Vg55kzpHCimEP0qa+HvrQoHeZpCrlDGyxG2m5kRWXVi6ICW8eODyTs
HQGl2a6inQFlOnF5wDrxwonW8PjU2rHWSwIvj4Fvh2s1sylQXY/q6aJL9hkbaxZF
Aygb9JpOk/raKuL4HV5qmQFO0e4kB8ZQTaVEtz4yQM8uDwSK2sOv7Fkn0l08UlzM
h9gnBOaZP28RR754lA1qd9hf6A2d3MDZebMVVRkRITT3xyNwIssQdttAe+wvjJHO
QeEtP8f300+XAohA/BSq4mGy+g0h/olqoByVdTcufP47SbEn+IP1juvIft8seZQ3
6JB7JCAYUhMp/iUIO7V9x/GjqbqEKiZpt8tSA3Ra6fecLlMva+2GNvzzlk3dHi9k
8/XuqkMrVb07vEgeD21CHMXU0cuFqIc4qfqNfwD9C77qP4lJLSerJLjkpNoY709o
mGL5galHytTG0uritR98YUw88RzgJ//Bk/mIhZu5PzO4xHXv800YmwyOBGdswB9y
56OW8r9+hiYnBEhWyjnAwXWHwF2/qC/NIYTO2k6UM3eI82GkrFxIg3XfE8tcGDp1
U+5ecO8wJpf3iSIR+6g0SRYQqH9ni5QASpd5Czieyvg1kHRY+K94puVSFzPe6mpG
LBPbHojbeKCGyF78ne0yAPvMqoYElUJtLG/yC88zkXM3fyYXoBFu2oJMHQy4qhiU
xCAj3xLYW6AQdJSN48/k6SLivP+GKXXuMASsUXJAo1EtbAoZiGmg7zG49eO7Njtd
l+zF8pEgMiH2PSXTyyQNrmeiFbzWOCjdwnr7ytPvmz/QrL0ffYjLZ3J3nbVx7wpg
kylxqhDbL7fabAJiB9ITCn2AnmXWgnvXWg1KZJ9QTO0OOS4bWdmaphn42vdEhE5Q
Kt8dysrzw9HzL9J95L4cJZNxujptopg6b/sSU3uuf/N7CpxdDjCtMAkdAvP0Xxq2
q+rboPBXJLue+O3/UveWEm6V1Z2t65u3MGnOy75TcyYbTBhjCvlrz+osYgvkAAql
2l9jRn/UrrqLDWElQ3rhu+lDxhU4JfcK2O4lKmTpYTjlDVGjywBzaOENYCTYImkJ
6QPUuT0m+DuwR437mXV6dwWBNXTZaag1k5xQjaAuvePbRdqkXAmXdcNb/s6O8Zkt
5KZU2IzrIw3xsecA+10kXo6Pw7zRCv550oHyylvCOCiYb3/Hzo6Cg4smqN0vE/H9
RGrQ8ycpsrun8OjS+Lfazufduv/mERzCnd7P6pZxGgwr8lmF+PkT8oT5dSrlu5bB
grKFjwc6lfuUNXuSon2Y89pB6g6vyX5TWB4e9+uGcAicyzHETUmvos+CrQovQ2Jr
gPqgibH7q7fULxqOPhuImyQRJ8KeDJYJA/VpJDp7FnUoLdhyKkLlZjO1oqTBbhLk
3U99P0nOx/7Ut00s882jSfo/BrixlmiTLtlvs9AC9ykzLDlUr9dvrIpJ8Bl+bKHT
yorpFoZvOegR2+GFGcsMzbeXfkjCEauJ9rUIhK22R6m9Q/0mcOeiVnixnwUybgbW
rSiAWAHyxZ7yywPwHo3fgzMrVbTyUrEHm4r0F3oLGuLyUNRY339UPQ2ZdtazXO/f
U2wNQk9erWCaQcrPDRF/I1b56dj1LQppw0Ol0bpUudzvPPzm7ZaNzdRbR2EaiP4A
+o1EE/5yIEHDh/UYeAGapI9Bbk+7UnR3oB7b+YyxQ7s1Er6FyhMPy8my8lt65Xl6
kt8g3OkWZgrnCWUA6hocg4E6XVHqKZPSZG7ymSRhgcrQ7ZqFXV9JN/CzeCBDJnDv
lXL3wckqpJj8wQsfz3yTtYkofg/qE5ktbirMoIUPg996xNTOak0oePVZQADUERqH
7YahbhY77Oi8g3k7MvlaokSiiHXRWruoemI7Tk0G/DTUMdh+76rJLkS2nys2kMGB
x6be+yzBCh5aiaJrmkESkex0LEiwQg1eeV2luvr5Ww5a8AeA0WbEqrzaU+jTDFZv
hvLjlqV27/WcYGfGtHuDlOJIbhFhwMSoz3M3h4yudA68vqc/TvhJb61obVZyMZKm
YNhJpX1BWylVaDAQrxR37dsF8m8jD8x0vSNx9tU/Y08tAf2ssRRXmUloVcD6tuyO
trHWPvQ+dpW467pQbC3V+LMPKOSXgWoaOTwDxO2qKEkc/fJk31ckjISF3m4BCAMp
PiBbQ0G1ciZNSOdiqb0dzdA4Z9Z1iohH8QnNxj0IuylJjFBADwZiCtW5CIBM2fgi
HFscv59WGy7ERK8zXVwJZpn8e2ooIgRVFxN7GiKhrZrOtJddCn0z35D+/mylmyow
jOe4hyqyZt8CIH8pkC8ggI0xQgGdUwleU0LVNAiWedKVEGU93P/dAyaKCmp8VG7W
w+IdgNJhLukB1NPPZsjXvp8Ku6PZWaZ86Ck+L6UAjz9HuVuS/0h+fLzsJokHPxYl
MdqDe/X50XrqYshenK7K5kqS0EhoI2DrByC3yVzn6wzi2mhjJi9sgdcSjRx6b9j8
aeuG3MyqTqnDELDRZnpdL5ntQqElmW55dY7EvytMt8DuKbn+uWl88PgpwZrQhoIQ
zMOwva4RBAJHjc+nIv3vjQFoFU86w8sggZApZ5FebKMYBuLrSfgqR3RaUDCbBwCJ
vFYTu4e8oPqhWF2SZ6Gz2Ef6l2BDWZ5BCP5JTs4MxFK/F0CJoqTIi0Zofc7saTVb
bRHLIQpFwLqhgxxY2r8URA9eLPSDbcU8TJzhsddR49+Prg4arqS8BAv/koCK+VPR
uEgegrfQNnp+IksZTfm/jCyl4uksSYSeCyl44Gr43nhJugImaZWTnEetlyQ+xhdj
3eUmPSc5JTiLKylaLxs8YkZqz/iB5zX1iSCOK5RoDCWKLZvhLYJpbXIrk3As6Obl
ZsextuZTeseHdu5AdSdh36wF/tBKib3VpmxuLCLPq2Zp/N0Ig+MQZMOlg3i2d8JZ
bJ/SOXUU8M4quZME4YfAEWEbh2Du579BhiIvbmpCJ/ySVps7WL1CfRkP71t9lJC/
FfHgMF+CHwuWV/60vqoJGhZ5fH0PU5VZYu7UDLeXxzrOn9F9b8qKhjg2SQUhOWX8
DgVYtzhUCS9LhVBsKOOO4pjkSw3URbAyf1jzKlUHKJGtD1mFze5VQvWEVnYai3d0
BWm5vOaoZyMZYFWxq36lLCa67PlbXZvpN5vjXFHdWeDMHnKyrtB59/CV3RIAM5aU
KfVdZJo+apBKTQg+qF55kOdFlH2ZrRIssRRXzicH7ms9SmnLj9Vqfj096lTfIbkb
sRzRNjwOnWYMTj9fZIrk8Ld9nwDMYGW82geczcBKdedzInDRI4TBjSIaicrTaZir
OGFXE+HS9PsiRuODjgEBu7ExODjQuGQuPFjv7YojJIdO0f/vowWaQt1FD/2wUINK
wxdPGxVU8MZKRLZ2ZPIpo4SimAN0Ve5FBWIzygdqs8N8vwcQUSqgt+Q27ZhfnL9w
Ct4gxLj4mc0KRN0/9CYX6zyMtAr6Sb3INkF3eb3giawsWrvIEE+kjIh5URrCN01E
Qi923L57dWWqNFo01GCS4ANHUf32VSVv5pTYmlEygTdEhd9SsGvraSGdPVU2l5d+
L3Ck2jPwI/yEUpgWp5NVMHZw1loaxxRXC/EwSchoMqiFrqZ9NzlNeEDAp1cGpFtf
vJOY2eiHQkhPAanG+R/LzIRmWTR/wk+QZ3FQoWzVoA77rzHrqlsJvBcqDGAunb4z
dEZqxFEbY4Xek5uz0+9kJf9vVIEvlRwh8qHODyAcAzyqclAxHJ62B0iRl/4Cp+Lr
+d3CP5m85m5TX9d9HiQpUTl6P8KS60QUGZXSeYSAfSiHJXWV7FmuJ/dhjdzyYItQ
71ytnnI+kcuvOC/cS5Ht17x7Qd7VSRkmhMa/BzDLBryp9gRreDNrv4+LV/nYXdoN
AJIsj7p5oWUWjhoFgbfN47u6/D+dcmdLmmIi5u0V0DqqD53VG8rD66rlByin0Eg3
DT5f0xdbcf3C0uxEs5agix4KKdUmnEarVxMg7OxJaDhnAc//gSHWWVJ//c6oR7NM
/qMA5Rjy1vxZtN89deDt9LD4ty+Q8HA0BcRJ21eWkGRblZNSPGJWol9TkSZJ9yJS
whGnUwKw+EN0Gdz2Yuei20sjw/MhUmooBJ3rN3TCAjlc2OdPq/sbwIKYBFPTqyFb
d33JE864e4/4deG0G83VSSRxlwm6wpXkiTP0Mlwl56U+Xo9xswxcDPO+8AZDMKWu
/euC9PJ+VYRgFo6kVwSKKFVAI+AA8xwlsCpLGXeOFMgnOmhxJhKJdMOuyIK5RNvr
MC6FO1MTczGgMWOKwKyzkwqOeZ3L/gw1qI6+IU0ZWMwh2hQByUyCP6wJwucaxP5L
lbcbyeFZCVPixKDeuyVi70Y1bApyVp87N/mwGFXFEaBCbhD6l1jE8kUliZ+RDQJi
GtgYsrrX7IjU/jid2zJnij8oRHfaX3gL42ECN2cqBM70UFW6QP7Wt+zT8cSO4YG6
jBg7PuBqciSxZYSfqH0bQ5IdfI7zwoD7JWfD66xPnOa/Izo1QmMQy0Wh5WIQch7p
HKEF7NQEWCH/NHfMS/8g5UfrrXP+4cTfcY12sDkBdsOTBkEshjiq/CRVAR4eDgL8
v9WNlFnlVBi21C+a/kyhwegaeMU4bymnU6Y2K8FCom6c5z2wUsTnCYbTvzFjnEzj
S/LfSh/Gq1/IGDVmjcpAuYNjRSFA8kuv4L8hwO317qB9BbzRyZr33KytfCQ/wc03
64hrWZornsUA9RHaq9WdGFtEYiDRBG0RHR8H4cJ8aGdF3vxx8Y2bcRJr0foUHjpL
WzUfEmI0RldWhSG39zJ4SeVx+28/5a3lnT8y+FzBHgKXyI6oA661X/Pa0yFajVGy
Iq+6nhkGZ7onpCpgzL/+yVTW1XP+dXBH3LIOSAxxP4z08m5y1c0+u1Sf1nYIhgYH
1C+QgwE2fMHZsqUeFQEz6gwe8uqnJ2O8sJ7fB6j0Lq1CHf6jw3EGiY/CEWzb+tqi
XTRNWLjPrASvKIqIYlMBADquKrZIFpuD0qm0K8EvqovveEqHJHVEUp79JOsm0j5i
hCT50XePQ4EyAQKckAvchdL4165GZsCnXLOTPs3S7cEm43WqYAAjYXANQ0GVUjEY
i7d5N+EzBjVuStCHXL6gxlheRJJ3ma0RvYd2U1FQMFgBQWYNnjpLIkY4noo/yzI9
gkfGbo2Midb0xgX0YOHLNvSXKWT5a7REEpZ5851czsdaRuFoC+huPJ8qXCJ6j9uw
PZjHZLd77gemjdE2GQvnY709q3pJawjkKETwMoz+Uc+X/YpFuYJJ+05bWQFWC4En
kxsnm4QKH1tao8GyLK2Mve18zqLCuZ1A09scMftqWuwBorAl8DcxMdEZrvdEkfEB
kqqTTllFyPrEAEPxoDMvRQr4HCfZcONVAwHvI5Yj6bOZtgMKduaHBfhCEmgemAPl
qytRhUxmNq8bUTxqdLdP5q/ou3c10KnK+T0n+G4JrWAtG84mIXz/dx6o2S0jtRTn
UzQIMgv81EUmVrPBJISWoIq3J6rHUCBTxF8YveF07imepMwmGvlL+23PXUlXEA71
rB+6Krsq5wNB3SItRVv/1U/Feai7EDggY1yi9kLGBmNhVcEK5eRaOwCv37lAh4QS
gaXYAHVYrLc054eWCALa2s3Io2fF95YfG+u2L57n9XfZCljqJhuagINrDzFMfn/c
3cKJI9XLjDu8aPE7zHKy2HndTMT2VXntZHNUPCaLYyOJAVNWxv+jlTa3yXIgqwuP
TyvGJ8acFM6vFhqkfC8IJHjDZHcqs4ZGSWmRAZmOON0AGTGQ7QTTYnR/sSQtCgq9
npT3VZdS5vGhZUdts0z5GE2ImUdlRiLMWPZsCkYDh/6NLOnABgmD93p0nnrUJrfj
Nq6ePu0NmvFT1tffOrFnqnkdLnUO+7hUNLPn3HWyw2yze/5kTTVU5ZFzXMJLD6+U
0+8Oz6yOpEGILLhkNHEM1JUelzMhB3y6198rkFAREUHE2rR+Ezt6zTmGcosDa1C5
vZxf1EavIY/LxP+Yn82hwDp0KtmQRbp7aU96Fw2pNlHW9KgMnPQsbU7WvHKPgODi
U7Zolc6mYtfySNB7UNKta3xwrIqk8vsVhrBPq2VOgRUAuhxC4Tn359adLBam/k4b
G7ykYm1+Afus9VgjW3CYggGO0Bx3pVhqXwEElLAcbtidb2aIPUwZ+zwmXci1WdY1
KcuA9dNy8awadSTYGrQPStkzsCQeaXbdW+sdKZ5ppxkNdu8xMZOoVAxbTNryLUsE
ThcUZpSlrzwLzQK/COF4jgXg4VPV7H/WNBR8WEwNuDz9Jh1Nc7WtmZLZMrY6sJKl
muel5KtJCBI+TgL+P8sXNCUdPaK+obp89fQCKItylbev7DfnnXeEZ/HS9qVShNFP
Rb5HEp9bUY7UNZCuAO8uRyc5YwXu/3gZBIiCB5sfiRiGV97ypmd+EzKz8uS+B4N/
EeelyuRAXupltH8sVfb4GswoE1uye2gwu9BXPJ5eMW2pA8j7Lpqm6/xbmIh7mR30
AX0SM9a58MHBUZ4ClGxhNM79OAjM9mfOU+27ammfgVxQvExxQpMKwBw8L/pR7WcG
T6tYQ8eLE7iutK3ndWPqUhBca24m8BaUVlcgQ0GDsK7D5JddGJxEI17ElWQtEw6h
vv8GgrDMABqlSgWBpdPrttsQXfqFxXhEl0eSSo5WkPpZX367Da5OfEUg0vXi1Du8
1IfbjM5HmFblSHqA0aEsUL0v7R+N83RCASp42ncI2+kZK69ZTebdW/jHJ6FedPYw
inBVxS9lFrOB8QusxEndgKfhIVSMw9Ue+1f65E0Bjw2wPpuK2Gj6DlM2h+baPI8w
bCNG2EWzusx/u2CW//uTus+eqL/cF1cllA9YvJpUUNPN0WGih6GZx61bsM29XR47
obn1o1s8cEwAzIELA/GgR++2QaFZ05UGbKFwP1TFwPs17sftiK3JptakIZgnU8nq
G9KEx3BJrXMZYR+yRgT61AkubM9z92LjLIN9GKDX+GXkO31dP1y/G1DzPDu+uLRD
8unBeMvNejOYOn80ghznS9cYQUGTVEJ4ne6Xpi9eLqsNNE/DCIdq2fIzvqtTR436
D9/W+K5BGv4rAXi5urzyosx5n0UG2SqK8p+Xd7fsAYWZo350HnlKEcsPmvONY4Dw
YlQzUWsBOdNSM01oc8GRDw0Bnk559tq1kwnFGlG+oqrbz0tqnrPrxxMRb/lM9D7v
QoZMCdsS7k99c64SxypExE3N0rmLlI7EtQ8B9BJ7Q/LKIHwCUaHlhXcxxBClWGB4
qZzWmlYWmv7bdxBGCIkmhjSQUBZZ8QMcIWJfriQ2+VZSZ5+izrdB09d2VAyhhkJM
Pz9pQlhYhhgwjVH1Lsba6Nz2GVSjoQHCp9bFfrxI4gJjvDtq87Z2GoNWgR9ScLqx
WJb/tpyhIji1AedTL+WnN/JrGAFwtWcJJJl9hK6u99HLAZVUNvbbrF3I38m8CjCP
IEX0E+zLfQ101xmHLUeHQwOvDw3Uzk6amYE3qfXM3wKaj6kqjt/RgTzgO59/8715
ObQhlAIyPvvz3lNgznHRjBNq9hiALtzu+gDacXIxNZcaW5HBR8WXLYTBZ5/PtYTM
W94Mj9nJAipUbbJI5+LesCn7SKibrT1FSTHdbXLCqe7j81s3t72mOs4+sbjgF+4e
aVSkDQOwRNKIF3TZG7+Fxn7RtEiCbOu6RJpdtGHAxc1nQEVQJpIWWhOMhIhLaoX+
S2DfygXWpT4r5Fwr1ws0ggAWFGnL2X6R7Ynr0Aqs8wJi5Gyza1JrtcfUeTA8sn5I
1Uj5l3yyqXjupC+8aWuiE4ABTUvBxbHgbKFhI8BdCxG0xjKEtIEJEng1jjCzUqhd
FuOMyEIfos9p0vji7x3sEhqZt3heG4zSnVVfq9iAKOtPWm6oJX4/5M2zgI3rch4L
7xoAr6yiY2RAgBm+xnCVRNyfQ5aP/7OZDDJfsh9aMDQ2I1jppanWdcrL66T8p9fI
Rb7DyDHy7a5ieHSn9rXH7B0C0JWbPdGYh2l/kgWB2QajjtgUEgzqYL+euIFnyUzo
iTJA/YSQGkwvCLZUL7MUwHCdcPOa0GOYPzOnv+4xfmF5MGGYHloKgAjXQYGDtmUC
/Kurilzh2BjjYP75A7Ux31AaOtxINT6qtkSu3f5cHnYWB9S4XlOVMIWFM5M6OgaW
2lojj6iE7l/my2LZFKy3nl83+UlXpnFBIBncEbSakwWb2pkRVLOcgWq1f7qbiDJY
bP8vby1n60ZoNbXVThtbOeK1IWCufCK5MmbdU24Q3Or33aWCX9cEHBOE6p11tUrP
/y/ZNJjVCfqOZr/0tYM/hQ58cYEJlBC7MVYPKB5VY/d5YfSA374uTnKYQ/EUqpaW
i2iLW/O7Z0oav8sxmb07RLVbVg3U+hmUQiJh3eseg3Ik9qAqPDpUh8ZViDao9CjK
xEtgtrjHyOTKL1I3LbhSqa/Et+KzL+G7jitZ3x7Kp/SY9w15y/3nc2C3y1Bha5Tw
8WgaHcqM+JBHP8M3miwUup2/4Uefk2X57TLE6njKSUYa9vU0th6uTXMrLY2/hPvm
b7J9zSZW4xB9aFJnz3iPh4sl3qDfC1kYz0YTvB8zJvRDarzcyPIvFUpos+oc6Ejw
abMakO3nHccUTkm13dxcdZ8VutRGU3v1PUvTudRugD5G3L2mvQgbFdYu2Jn8iYBP
Hz3wyyyc1HItMQCUyYyU3ikfV2rjG43iO5iqvTSNldvUFonUBTyToGY0H9HV2LN8
yqmbMVWy4++hffLxjhfvDmSZVNGFX7SLBP6I+G2zCODFSRuZw35gvH6pVcDfry0x
+wmhnNqaK2W644Y+v5Obvpo7gsuBMQlDACyUXpT+ie5YDQ+CFVioLl5lbpIFVDP/
L0U/ZoAPS4dctRLvdf8JRHfkgr6GET7lX+JMHH4K93DTbeNiye6Ybh2b6UcGx4FS
/+bSx8nwnZTjA6uAZ8Pherrqvq0jzvF8F4wFlY558/TXed7ElUSiDfznXZDgcxxK
TBVg6UufbZslFrs5Mcn+sQigmLRgnHYSBowXVUZNRkf07N6qnQy3shS7a1vCibef
8pphaUqun8M6MkOP1mfEoksyatgoZ1bTz4EPWPka5MzgM+giw3ytSeL9IfeTlIEL
HJoRzAYKcbyPJL3hOAc+ePyP7JcOLbNDxfdoa53MdCf3pO3wdAqiFfORBL/ddZ/L
pZoy0L3ZWGlT1VlxCH6QfkbJPlh6QaewLsxTZmlt7FHsdcajfe/+fy8vPaQGZZYU
5xOBYrXCPxvF7iI7iM0ACrHquW+gl1rviY46OyIEc+LVgjW8kyyV9SpHtS24jSC8
5MHnTfPiXFLqI13Wrp9y/rYz4vJ6dFaK5MXLhZnByeJosHzL1OUrxJk+2ahSJaO0
3uR2QVA+8wdWcPpfQ3sb1M+6R+yzPZ9WD2BdcsbXo9OqPiKLXN9Fgjhu72H8MrPx
y7DVjI/O1maZXp61fyuwWCmFkwKwet8FhzV5A9GxvrVMH9y8FO2LSw79cAXPVFcJ
fvros1m5ENqjFWwghglyZTH4OgTsjKGSM8YCsErcf8/2Cds+Tdo4mNB9U49fKg8R
tTUZbBLBc9Lp3yiVkGr057/9mjaHCFb1fG9zhRRo5QSFRyElcpWDXsvPAb6Afd0s
EUoNgD355GuQ2p/iwczQRUMf6sQJzFtv93MqsAcDRUUQAUKghFSBussNVToDIE2r
o5idpDaL+Vla86jXoE2bDCAv99000J7T0R1zIQ1+ftkaMZQLcYI38aaM4YYHYWUp
oEwUph+7lxms2VQCoiZaz4eqJ5ek3RkA+rAo7PtZjw6tqr/YZjmwP40264A57viN
NqGwFGAPXw1Rz9nAbSCvzpKJbXShZcr5pUw5YaLpv9LVtCVCRZwUY3Pa3OojWlVU
Y+CpnfA3sQXp20qu4h9BYD3cQji9RRL81e1ToIrmiqnxDj4eb6wy2xc2dUBFT3T9
8jWhYxRaaZXOKpTR7QQo3j3vtNqcLzwEbFGaKEKBmNa84NsgvTI9n33KaMsXxUKK
khesaTYCgsMsGhhMHgqIAhl8JziOdGAFBDUNp0GC3lWf+a/MiApUKX12sumyLZF6
/pIei8hbfGN7jLibTI9Fta6NIkEfNjd34IQDvOWtP8wEZj/Qgjt3wRfyPEgd/gDT
ehSAqZsYtj+sDnGjd6u624WZuoBOJL3Y379kS/xaIZblvAadkk9DbUoW+cJ1/kTk
o6rxcatHI1GNz89g7UevuQDp2SeQAeqY/bkc4En9yY7+3ZDwHepwZNoHBlQdv3L5
V3IALUNx7I2B1qzS1UCYE9RsFdHWHPf2ot7fNbbBx5tG7SnMFAyBpLvvTgBsNo13
wT2hE+qtkushYKVoL05es+O1hyoFGa5MtdvgEapO6/NvJloKAptUJu02Coswcc0W
3nvER25UFdcfsok/6tjyNVEtNPHykO7BI9W9dBkXO2PGh0wpEb3mAqb7PTJObFRs
YLQVD7yD15YPkDE5Be1HgygmSqhzgMgf2m1vJ9wiOPjhdwQ/hGbjUIgbtmkOQTFm
uW8alj6Gl0uCYo6T4LyFHVhzC9GT6sAplQ5XKlb92ME3xu4BQV7eP1WBfVhHCGTp
IVDLh8j4DzSzK9+wCRll6yp5eSxlQ3bQ4OWBKU+yrFYnMm0y4iEQKcGx9ZghklPv
D060fkilG/UReBq/yZES2751+x35OpWX9UehurIb16yYLgb2/F9eGfsxcHxb7caF
vc4SAQJ89LSa8ryYQ6jS0CWKvSkCKewl/GeR7LqtL4rErjTg71Tbi6GXVJcE+6tM
37UUebYDitiPhgAi9WSNdxQRmatLCLgJDfsYg2YsbtIq+D/J2htQPuFURneC4gqD
oVy3XTeImewMZ2nKjHB12peK9+U92Em/Hrl6AqgieTYXrIdG74ir1Up7VK5UN2qF
mVHo0TrR2MKpeI4f9tg9dFt7x+YwPLsJh6Zcm5M3y6TLgBvH5LiqhCoIouQPvEAv
Aygsz6H2rxNMyuj4qRpvLycvYCO5aeaJ4LGzAkN5u91PGI5PZEzW/IhlKG+q7Sbx
DLEx4Yv4vJf9P/qkvuGCT7MEGt9msStSH+oFbqvnvW5gN0uMVcVt9KO+SoEjXsFz
ooCoNdCIC/OoB4b6OzyV1C2F/BF+YGJSrudoBc7h8G1DsOcsgnIwJM1BvxyVChcb
8G5+UeqtJC4EcXZnOEXIQhu8dVbpfu0ta1op4YkUHXJJ129h9XyU8Fbh1Yp1HEuW
4cHuvkDH3G6d16uw0ANbRNve+Z78o4+QU9rwyKikWejwX4q5i72ktV6hKS8xtK92
3oTFSSpSTChoh47Hc9eOs58yQLsnBLiraroz1Fj2JemlSFiMsYYwT0n+0jc5TXrM
e99REe2GPxeS8p+zpavJlokTMDYQJeU8RZbhv9qxmNmF9jOTZokySRJGB2d0eHU5
i4RY77UEXrO53vXAdQDM118jyQFfkWhsVyadqBxGCet42XjPdnGsBMR+2a64g8cA
3Z8iusiGkSSq+R1FQtJQlc00ngkKlvOy2gXi8VDmaCd3AGPSSII/S7S2z/IuKrsO
mCMkZ5YD/9BSxY8txle2awSc/Zs+8/RFjm1AVxYOYcTMFvjx9rQCCH5BDBkjrG/k
aqtIihn6a6T643uVz0XwsX/dhJ+TUNzryx+XHMy/69QjMdWD29jLxwiOsuFunVIL
RYDfdLyGvQbjsEPpxm02c4vusMmPH1aCWE5sOoX4UbGZNX0qxk9Zd0U1De3ecqNn
1eRLhCIM9A5vdI0ogFKN9neIQ+5HHCrF6ydHWWz7IMjXOe8Zj9U9k7bAEpw82jfX
z9O59NFO+KNY7cvePwh6PjGcOVsv6L+ZBn6Sk65bYu3jL77qNwzDq3QdCJ3BhuJR
P6XitDcRStCBqdnN4PIoAFT7e4+7U+mRMnwEE5siXcGyxpHMlAbB7Y//Ls6ofLWb
7s+3KePbLRPqcIfokpZJ7Idje8z/UwEc0/u+P/RJb7k/4vG0rA+OIZATOreYR47C
rqNMd6LQDgzXTIZRc9/x+V2AKNfDeirc/X6wzBpC/svYW7VGw1x6LTd1h+nqdb4j
CvPv5Ad0MYbFE2d4OueYyHlY43N6iAgrWiIPDrM07UfH1WEkLVshBXAFzw4MX3zm
6nFXpR/3AF49foBZFzyqwcz5SdPR7PeORWoqCynGw+/4FRzqF/qRWqZDRcXea6ee
BxTTPgKXcWAI3sB53ehJe/OhY42YgAWev0HYSHu2b62XZKxiHObodGC4GKSUxA4i
bBVJZiyLOGevvOacnebtTWP1YtOR0FzGAyP8Q6/cp7wNCN8F0CR4KjQM/sAs1q29
xeXo0riQSmhT1R3Q7UxD/pU3yUkE9Uqj9KWjE1LfbedSTDSxSn0xDJ7Gyz9S4aw8
V6Rlp38b153uk71uv4FDkkOpGMXexsRFRbXhGJl1oep3+OsrAGhWHk4AAAW5gJKY
FPkn8/eYLBhd3AmgxOm6yMYuu/gfi07EFs+js0zRrPRDw3q8yMCZRTrkk2iB6jIQ
QzHr8m+7Fd3NceM8oKadjxc769z1xIUUrGJdY9CvrfLiE1xB6H6flkKxuwK9fhMa
p619r8SxK7peTKTcu9AI5lBAelUo62k67CpnuWRDdU/Pz9L4ei7sEMM5lct4JWG6
1mJnye38maUhjinv5yeB/BEYCI+oZLy5ui4a4dx4tGpDth0xVYRJ3pM+W+wbTmSV
sj+3oVeKex92YHsAx1vtrZN3ngQFYZ5wJ1vrjO7dctzwjJVtKqLKLl1JzM6rAkDT
nfB6IgaWUxFPHEkDMMrq1A8SX3qEP4sXZskt8vk0O6F2+fzEOzFfKwZTmDThBDQI
nBJmE2xvhbipQgoWDTig6cqPV1O0et0Y2tKdnhah3xV0UH74P4yD+LqikOXqveo2
yW9xE5Jb7GhAo4dFsTARQET/Y8TMSAkplMNCEyt+qL2uZRiUQa43tZoxXcuvjF3n
fTewyKa7lB1IFiiUFLg2UP+y4iyETAcFsmD8oHSg+tnvFTZbMvdCDYAJAE29Gl1Y
Qjd08h+UzMs8AxAQyvgkm75TF+/hB/5V/NsVqRScndsZsnX6SkWDRil/++zjVNZx
WeU+wIv7t3KiYrXmmsCdGclKkwTOPNnAXozCLyiBIX6aGoL1XTj0DCFDeo43poFA
ry0ZnXlTGg03SVPI6aKR1WowohhBEt3MVY+ntCdtZUHAeMgNfcKhYhifTGH/E/o0
AuHWpAZOw7Y4OL6JX2o6ujsG75XgY8xKmXVpJtli3zwp5UnOJVi9cKDCFA1VfKL0
IGLeyK9KhOeruuZs0bK2KJ6znIs+KwutMTJcF8C10BuU1zUjbMZFwAOAKqJeGV5W
kBljDzmN5Wa5Z6cQ62Xe5r/Nik/tZ38AfrWEHoQWJcaAXjWMuEwWShq41E3+Jkyk
yv/gsDf4mUZv3bCmyVNg3dYHxlWOqFL3m/FNMGic3bC1oCUDal4pMmIob/Uaun88
JOsx/e6WaPoP9kSZx++G0nf0pMep5ip1+o5Z7de3plwePZkEiFULubBbl9E0nBrJ
cjTeIfkHvPZXaHsb7bLhWS5+DwjfSNQMs6dkQkih+xqlWxBsI6sdwaPu3H+JRiju
dInXgZjhum14b+/K8epIfWjUuvSPR3arBEYoKBU43WfaRf33qH6cmE7emUcNkpmS
fc1qpN1sxevEsTBjz8SacMM5JD57kaETyKqFo2rupRs+QvdyZpvbXVK0zcGLXdQb
4nAiRIl0V2iHVSdENFrnrC5LOWwXXbmbFVV63JYzjbUfNUQRB64rzOJj9sANkkrx
9sVE73XPPilZiLPNiKhtKHJmeJ1JZCpZSSRYLs38WNuFLGt+Hsxl4rm7zkiWbMoV
UvERgKJ8okXzAEvjrlC1+Vljd+F8f+O72vxc6Emu0aPzKBxDSGc+1/tbBT/7uNTo
nZyzU3vLnqVQ1Bpx2RAgVmpIQ9n8Yie2S+JYHUesAJ2dSL4BkWmzRewcOnjdiREj
9unm0jMDhVzhslIZWSV7IiQ9lAfeaccKuRiBtlJUp2MEKq18WMOy72NpFb4jLiGY
UHDadMZL6M61Y0G922FKQ6kiZkgj4nGGOm+BUOOA2Kuuj644k6P4YpWGpc2kR6cz
iWuLFv1Eq/hoAwkogzJMKZPaw3NOVSURFZ9o70QhJtMnRv9YAd6srBDpKp3+dLVV
tufE0n2xIU9HGXeQndHG2kPEYltTSTA5RwtIWItaRehpUD46TrP+cBlaj6edMv7i
07Z2zz/ux9acBwJ6h1twp523KqelB9aD5bmctsd1C57D21x47hlk5jL3VLONMXlo
kiPRdscPIkL9rJwThBK/bOUK1uOAjva94/M9+6WFiJgDswvIwVc7uDC/lkcMoOFe
nHLvdt1amu01Ux76YTuBi1MVo+pFKUsNS6XFJ8OxaVIlUl+a3thvZxWDL0/fRDE6
EaY0fbK4Ze6D2sy/Qhh9rsP44/L3BuBQVLWXPObJzPyz1GaJdBdzymDOZ60kpqfE
1/wLOVTI947olovs6ILrCr6toZsdqCTp2O1jwfXINym+OVo/F5UgAlYEfaR8ViqE
i/UmEABUDA1qaH+jhMws9Sl6UD8DaqZ8lS74ei66I0L6Jy9md/XRlH6qr65dLmSZ
+JJ+MgnVNbuadFk3qMAYL8YReZUf7hdwrgTGlVwcsLig5JcjTbjjhgIiRLdA6N3J
e31/1g62RP54UHU8BD6oLnZhJNgcmT+D80nBAIujw4MGmUieIqfdQCoLL6XPx8im
81TNNShmz7PFYhjOmKTGcPAvKnm9BomKmufv5ZP57td6biv8px4awIEdPvN0C3TQ
dIGUKwvt2HT0hJ4/zNLe23D1eI1cPBx1ln2uhp6Dwl8Yxv09EB42JRD+56N3ZVgH
7ulAAsdbqa7iaZWF3EGsauW/MoM7tyAOgWwG/AAi2UZs52KPOvTfDTTlaqpWRknX
rZTFzAfO9e/cTZKtD0J1HS0Om9OykqgDzNERW/Ot5UBdHsi5Za3iRDWRYPokJkrN
vcVmJ63N5KNNw/KBn8dRyIdNIvkHFHXtG0ZEAqUL+PcXalQwkgP1J+NTgGfd2r4l
85uHWBiqn/nLW7suGifulvORdms4jxA7oQf+06OfZzIHW7VqIZv237Y2DOliHzAC
cC+23yy8zc78iWDGcD+DeTwFTiMDJaXiFcH0fG7K9yrbIE41cqyHElfDbc4Liuki
5CGkrab9kcMVqMv0edXytPzCJHqxAMg01iUz5Ej0L3KlcyVJ7fd5VYr0EdpAqm9i
WrLXhv2+wUh699MxT8HwOiXwbjIVQ+T3pFaGr1tXYmf8hwEm0zgwqFPdGUHzqZCR
B5iVNU2I13z+MXl79JL6+JBzSXzSTwm6MdZL72G3P8p8CUN8uli1o2Ne7wR18P7K
e0QyXTXy3NM6c3dJAwEdJDsOaXKo1ZQe0AG/GRGNkPuZ3R6WZsgIhFQ6Byx8AwXS
7YR4u2b0qmIAmqonDUCY33c+dMsNHPCwKnP/+3t4YxzkMsA0La1selPOLdfUObQ2
oDjJYJLui0L9DG5GtwvfSNNhPa34+XINwjWvQoZxDehD00+6GeSUsdbA5yRHyTJE
LvIQi2Jc6skpbnSUpEaUWWy1LmGKEN1Vu9DIXeNcS30Wbpb8rdQX0jKSddC4RpTW
WvelPVj6oi9Xr0BD+s29IOP5Ua+aDu2oewcXiwUWum7RReYA2IxR4KMB8ALYEsHz
cLcE7+x699bnizCV8C+8Bo0xkOuWvwinD1w/21PwYT/2fp4/K9E21AHkvfZGKaCw
aCaN5Yr71a6OzkfLE25UoQL6PmCmnOIY9Y+AqfwredmI6P9Z1ixdKPKgyATJ3xH0
iQ23BREZg9PQRSPsOAm4Tw7ONvUpD3hJ8ITal/q42YLYfWcd3jMIm9M+sb4Rm3wh
FH6+3Nn2vkvYuOrsu83y3PJ+jlcCZ0Jer1sWctVL0AL1dmkc63vCiep6BP4XpZvg
C2WrsZFwcyke5uccV5XuPlvwfdcz7ych71kRebysX9jLKkiD4pnmOnQutPEf94Xy
pruq+dKBwzlxgPqzA+i24exXRg9mgHVp7qz62i5DOkuY3tHl61P5hJuzxpT0z/Uc
DX2dKeCror2FGzPbQcMFJlJSgLw599QZL0obBAgaoNAQdNK7wp9iBnuN80iXsRcY
MJ/p8SXba9a9REOGesuWrMcQTKzpu9B+knfL3eXo57sQ8At/YuBek3p4sxEbr4cV
eDfV4FyihroqjEfu1scZu+HIesYGcNVwEgmmAoari2U/1d/SaOICJP09X/kzw0qF
WRz8D2Rm01NOjby+gOfT6CLLvmB923VQVqzmWZU1JtOWdxLUIL82byqy0Tt901Ry
HIfdEf5IEJbSOy3PpPqz4T47BSZXFycmkOqoXLacgJzId1jPA4TrMVwOSEZcjgQ3
2uTGd1AkFLfF7sGIo33hzyJPxwHJgPduDiLr+O12OTm/mMCW1qP88bO+1Q69R9LX
MLQ5hWP1eLIU2byaUmvUJGoKRqBueTZ7iocLTxXwLQhKU0vmjtU4I1vRURHemO1O
vFOiTIVb4koGcGCqXYg9i6iu+6hgiaF4ZHeflKSAPIIugePBOmM0PcbmKhdR/Od3
0YwRoPnd9DNk5nliypaZRbPvLJ3oVA0mchQCu68EQJFuQnRjlLSdVTnMhjuC1L7t
Qmijh+YBVTpjoJBrdXONmAFHLoVP1y9MzDN02wnkdS+EmnPWozCRS9rJvZHMhTXf
FKxfq2JyyUB5sCdEiBNDOqNuIk+rOyXrfaDkP/MzugxKL5f94ULd+KhfGEH2aajp
+dm6odrUCM4Je4EPuTDpFJF96/8E5chLvr0kUNVMRs6tHOkg4Fb4AOkCkNpdpGH8
NIV5hhuEr2sz8zo3/3RjcYZZIH8ENqOdVPeU0ELeBhtJbIq7QhlqkXwxxb1l3IMo
jbhASzmVpv0JG9kDc73IhGRIVMnw3er+RMdKzi1GWW/eJEFOHvBHOjdPpI7Jal6Z
2y9aRFaCRRu1sTYoQH6A64LKfY1ZaVQx1A9wk4dd888gjr1rX2uwF7AL89KJs2FE
lKeL3UTRk0F3AE/QJtznswKkLZLmFsYkGJSUf4/PrNyF5EELGzjlDdt2ED0JsTqs
xf2r0VcWFsdcKfHW9ng2UCpgXdAciKmi4ZJTA8JTz6Lhi4CDCurhDC/L89BaZ68h
6loEXJ5aWU+Dsrbb+BmLqr9lodfBZcYurNyfWKfbrFhlo+K0I5K8cRZYali+0jUT
CQobSE+752UUsTs+cTjOjJZzs+7rtAEuZC1ooMBdzQQmTmqRjqKO8jJVU12TxRSx
0tPiuB1AR8HQS3kwCARmPhhbXGEex/2hiIA7QAhZnYbGMKHCDzhQwDT0J5+yggoQ
7qYXpQtYC50nZO9DwCskGnigAc8U5i7KO0N3qmJUGqsXrDFce6dy3uz9AbY4j7zL
noiCPdzwQob0Ld9+sNHg/lAbpYZku/Gv3w+UKiAWGKGVRIr0hkVkiodcg2SdLjM8
QdEw3wk9SYO5eVUTeKF7n4vJkqCJXW5tb8TMGjMzrbjIu57pUnq8pgxMuEsIHtAv
ZZzMYDLrHAsO6wLCqqPxrQJAgd8FR2conGH2Gu3X2oGuAhN17ecnCg9oKkLxYHrT
h+9875dS1KeAz3a+DtycNROp4DuaRyzq8xD4dtDbyfnqxEW7toGS8ba/dfwpLN/i
DFKY6QkswtfhcVbnV4Pp1rtofEvSxg4dM7K7dKgvX5i6VzYIgsS3wo7HmVrvZ/B9
zUEWj/belUiLZNOF6yXn8GxHZXa3+F6a0wOT1m+uyFbDdeiz6YtKlWVv6Kqti4gf
AThfDW3e5v521N6kMha8B8qJe0ONkrNRGZUhr6KygfVc+s4J+2vh8xcuc+Ta32ev
m2TuSpVSwXxVvE6if49zeEjwzmbbankRqdN5YynkbV+GooXpPFGl3oNULCAcixcL
08vmMeklFrOSSDXlQTQ3XCFDYqFX/admUTBOBnRLBHFQJha+q6Unup4qSWMmo2HS
ImN+Xw0rbRtOjrcAvHheEijw98HCP+lKW95CWFJAQ10sKCurK4F+Etp3uSrfxnoL
wsZ1SiGY8VSicEZ94Y/Z3JypqCUldGxOZjroDPPGfExtjNy9EoSzP7kkE/V1jMdD
W9UUceACdzVxv7dxjBK4W8hyZyOqzpGehHyr8jZiFXQX75fZgXA8e92uSkmb/pmX
9rWLaGzEIqspzJmgCd75yTMzZmBOYp7k6Hlr1fcIZKQ1VqVli9tTzxgnmgGcFpTX
9owmXrZmV/8B2q2Kumw4Fvarzk7E2e0MXjHJmjYISjjne7SRDaFKDq1RCFvJ5mKD
UiTmjDjn5bMZiMaazNxsi5sicPi4t3kbB3bB6pUEs5VZ7IBBWcwPTBZsZjxzZ5Et
OcogVl+TBHyylpLUgWxZzIA6rn5PK2EtSYDgP+8LoNS0FmVvMazPY/qnWEVwq3or
kuby1RcAOyHcQHobPmXo7CfiEGx+zjPLa6LXjp0DeYJVv8jiLJ/dmrRazw+A8unJ
NxsybyWF0KlBPDLNTClDgwceXCDk9tBKtlmGdVzCzCUMJ4i68S09PtVY2M9GYZ/W
E3Zxe1tQ1TIHck4hAvLQeu38YEFXblY3190k52sMc3OHypN/gLRZF0gNtBP9YQv5
kJaHP5N634CuDSDK8xVY2w0uAmibC50+hlIjBHiuwPwTflsroaHG6XBQ+3Kp19EJ
eEXtFo6zemm1AtYCmzYAZ9ofjF3YRGW6tkknNcfvsGFxG4EIHfRGjPLtVBySZAQi
iL4SzwA+dxMOM0D29L37/LsTwTj3D7B7x4j/Q7k+6HPfaTAg1Sphltw5vUnetmwL
lBjyhJ0aeEHi/l4bqp5W4f7Gz1zeARQJBBmdD+XxSX/+9qVC32c8TF3oZEcPo93X
Jv81VQnZ2RD/7x2GQGOz4Ay4D6IiXd7cvZszuxhBIRyrRNXC1gRKnmJ9caUOVg9Q
h7JlLmbeIERMDKBoaaG1bICgPetlppMoFvK8b46umf9CvJgR+5OwmsWlVGpOhKfi
hoCoAgBmAqqqTPhFLRt6G/kqPpVjjt5ddCPitOpu119Afdh6Xsx/9YYgjFravRf8
ARaizCOMcUDd+knkyGOm/cGcWMuTIw2gET9wtT85IXEEjlXDR9jiiH7X7WTwTRTO
w0o8JzArQH7+BXEHrU32cma+XJjGFTOGaR/m/WkC5Jt9WRS5pZ7wsglho3IvMA5S
JLvE52NjRHFikVHlUKkgkyHlicD1mle9CC9D65HKQkAmnxkP6GdnrqkZJH55WuFL
OKlsVoegd3UYI2L+upGO8H8McmooYezlCzAhpaqmOLw0QXGngkeyc2h4be92d0FI
1nfRrPdG6JRFOVsw0YmW4fbLBC14DuBZnxeiSMTFBK9UISySyUV6FJYf8pYvnl1T
qK7J6focBJbSNUrbYrdBRZTKMKq8jyi9hFF133R1j9nWRHb74ob39oOllgrwBhg/
DVUS5cykdvxyGmSN8pQdz2Fw42OMp9TPpM7ydsX5uij+hqnh5+FBYm0usYC1hXqP
hBdYih9Q+onXhedO6UV0Bu7cbGDW6DLzbVy2zulOHvEX10gBGFHg8bfV9YVALL9Y
zlBBkGSYo4qL+HIO7x3mHpAgt2pOB+/TzJmeY1nn08ha4oitmPSDJ+h7OwNF2AIp
XWOQB+SPuH/dDp2QmxUGSFMVIT+jISub/9x4U5KgH1MKd0BMb16TyY0vV6Jcnqu4
rF18dYWi02EP7v/KDw3sI3JDYBU9RZVBrdEpqG4qCUcbEN8cAzhuJuJiSrt5woyF
Xf3TTtLDm4GXB5C+Jy/MzHPl4wehKoFZ+pRMkCLPc6wfNKiKRpjn6/ABrqwTaC/B
tOjoxGWZavy9/VL0oFaod/NvHhXz2Wdi/DJaApODqAXhiddYVZMSMej3zaor7f/a
+arfMjtrXOtT9gZqrZI0fwxZOJNXKwIJFWiUrall8vBc+KSTIzIoHf2j4ImtKuUW
fdGETEkuBS6aRS/Ee0ji+OsSbJdbsSrF6RSLGOBCMcIOvq1tCdo1HhtCUcXcz/HD
SiimIhzgt+JlZSLn1MUgDhy83IW8yC7NmkKdlF9oZAwUflDHqFk70l91JZhJlWlZ
Qk7+m3W+sFOX9z1fNSPxwdNKUCg6Tj+eBhGxB2wWYApRIaq+ouxZD3aXRqVdEAAR
c6etevmacVQd3LkqYRg/z1hyfBx3yeLH5NW9FnpfuhKu3QGNqNSUuS8USf4TitHA
P0epF388Jn+Sjnj154UcloWsbRN4bOJB3PTmYC4vVH93TLpheFSD3soEI7fw25jF
k3I7fCqvOn14ZzDcToXMYY4z20WIvJrJFk0WB8EzyKiq8MkUK69aRPLxEEejr3Ox
NCN6J2QCsSzLELsqDGgDaU174/K2XMOlwmoLiDQbkK9mrx0LKDZ0/nrztgee3hzK
uJBRG0Od7DuFe3EcnwGpjKa0PCOMfmKb8Abqxa0idllEQPbtvpd1cs7nGh4qzIc6
pywVSZZnX3nFls0uzBcob/3Pn3m0YkVYuGdBBBptuODtY40HNOH3EzdVqwyLEVcH
zPwyDRxH/caOTD5AUXVkm6keONiBUsxrJAo6IBD6PcVH12IWoimlolH7mmGoj3F7
bbRF7yo73iU6mXlAsxlp1+d13dc5SgW+CsXQ7qcGuUnrhMB0w7JvAO1I6Lw2+dIw
pbV8JjjhJ23BSLmj4eI47cmF86nUQ/tZhNMjiRs4NGMBMIQ+zH9um+QrnVXLPFZ6
sMxa3jcc96SsYVoOZ1z68wHDvkfP1ppHbw3zLoyhCKVGrDKEt1nKNgvjsdF587Wu
jsueozlUhWeo+NzkxPXPxIEQ7gu+iF0n2K0kdXUA5BND57rr2mF1+bTgbSbgNp+e
jKfoXNs7f2SXPs5vaR50EuZTFSvOTCaf0gklwDZ2KXvckodKTcErzNeIHooFlg7X
M2iTJBk0S95RUrWoKfFaeMejwODq22ZeW99ud2mMKgfckc+4HwI4YjdNuxhpviMy
pGUvxIIJZ3oqXS/wFjnlynbxaHPn9nkZNZr1vsXtPW+pbD5O0G0aIG4KZAC3+HC6
j5uVXaoVDXzMPwh41R3fe7XDaAYaMd4oYyFFUGRJ4Et6CpOWkLevh5x8ATFo+8jU
eLy4fQT/f0Hj/qZayrr0eK9iWpV/fAKS2Ak7jhzdZeSJEa+ZT/zCiLvbRH+j+nKV
LhyEJTdevkgm8+wT9hz6ED1IanmXzIy3WbhImDdMAby3cflFBJGSHMFaKTw1R+cc
mYre2yOxlDq2YzIVu2hUakbhoIv/o0MlNM1sqdwVL3Xq24MaP8kL7fkD8B19ZBQJ
27VRRmJIc+QwgWW3IaP93aVRWE5C2QENagO1Vx8WGntR3g7ICVUL+lBSz7yWzxvd
Rpj8z3oRab0ulT/m27Ygzrfk0CKlUDyDA4lWvtFmgc2TODcqlc+mcENaj9WqzjUr
mvSz5+EOKlPoFNH6KG+uCejGsgimQIK9bC4P61On8Mn5iSfuQYZmXRInPb660bNQ
poLIGe+kGsIU+3+kgGcWeNDTMQmGIfqKikzsi95XNSdIjzH/2IErGT2ESSCcmpyN
zuLa28xAiptBVBB3X3CaeiLyTakn9Q3D+vF0RL32Ib6V3uuC2lTS/lvgz5stcbwz
qGeaQ2XXEbHrRA6YsNyNke5zan7TX5iXLMAD3rVrzawngWhrVU/VMpeHvvitGoC7
kU4DhwMLusvECYWWLB3ij7XUd3ZAYv7rocYk9+EHDvjRxbVfSKLQ/D/0AfrYDKx2
K+ZVJENwe+lTzwvhg3fSX1B7KmQbrOF5gck6Q69J4m7oAwLtUZaq3qgzqMDwTlHr
vWEqX/0vxGS6QiHdBzaffRDPYlFVWxLGhXVY19ffzOwG3n2COQ0R6VjEDCf5H36F
o8lhqQpFjzbePc1FmCSfnNr4fEAnIBLHXy2/Ekdie/NIXmQPEufcaEc3P/j2gfRk
s6n853fCB6weSMwRakvJazV/lsAMPGsptpl4+gAdE+Y0qwY6cqxJky8JbVGMrFEt
50yIAREvUR6trrm4MX9t+lvFTBoyMM0Iutm7kqRdIZ+pd2CUzwYYX8sogVtT/meI
x8YjstjRaQJ8fVRdud4/recMZEg20UOMLoqBHfpXP/EpXcbgA95PCInKRpBakAEf
PeS+Gpzlsd9NxqZsYzguzjzl7gHGOldOyxe1/FvZmRav+NesY/d7oym8xpXcNL6E
LBW7J58XTwvugGQD9m+lUtSZ7Bs/tWbjp5UZo72I4fWurr3+MHnvVX7uu/5fQ9NU
/Pac3zUMsv6lhoIMkpLD0vBQkVWvYZTgW9S3g+Ix1KbciJeVKeRMOqftgjl3hV8z
w4lmIvIXYweCVj8Esw4oWw95Rdg4LCmcwN+hCGEUyOrwoP69Uj5kpa3/97oRCOaM
d7WOEZzGSAStsP3bwcS6FOe2UKArnJxxvqAKL9QlkTcIBiNpakCi9B1Azy/cqUeo
0KRzLoqQG7ML+p3l4SCbW3+ysaozKJUpmKST8R70A3ylXWSTbuWYRfgDxXgBCAvp
WjY5vxVTdubnYwsFHz6PefGzogpbTX5N2mq4jYu5nqfyDQ88bwMZFI9MUaEKQJMg
qTEAZny3KGPi4Pufv6kIsLQL9kGJ7ej73r38e8YQKqXCEBbl8FFYGKIt1A9czm+6
6TlwEo8QBXjponzvm5vthvxi4R0m06XwEM/UE+3KatsRIQ9vC2DLD2UAkAr2fD0M
PVqNPC/uCWjHyh9w/i2uOe1VSnauwATN9z6jLF/p9zeMKJ4dWb4jkEdgBwKQb2iR
fjIm8XSMIeLQ30BmvImU7dtKneFXfOxYthSRuazgSyCZ/ENBezDTOiWTvhXtYfd/
Qz3X3IlC2l+jaMlCItCP6PTEOVY7kZnQb7mB90Nz8laB1Q5AtmFHu/f/FkMHIRea
jvh32/Nk913n21SIqanr3mltKLvvDeCJkZgrS0gG7dUPzKo+Bvm9usbV1nd0WLiN
98YymqqTrrtNLjv0a4MLB4Tm6BR0iXhHw32O13R8wGiAbRCr0kqC4WFmxyPngwRG
FmNNOTiLDefI55rCGVIrT3T0k2z/Ma6IjHkjMcQ/aFmNa4SfDLaYjYL/fH2iKE5B
eBBbg8hKxvMVTDfTtnXDQRvT/17YdvMsl+sT/p1eSgo6/F7Rj3nmy1dlHnJ3SHtV
HQ2eVsxyLDC28YFs6t/DUIlpqw/B8a0ybhjmm6S2c+RwrMz/9DYzpWN3Cadg5EOs
EzUp68zivp10M4idJQ/s/L9WiKDdWhFs9saJCKWp6ASrvCtp479bbh2BKbpx51Y0
RmAsTB6FDjGozQu3SllKeE89tlqL5GnIPOlC47BsvR5QtW/YULThuTbMxAZypc3f
WEW5X6CXP3V99mdhqRCbRtzXHrRaBCVDG3/aB8mRsXB9HjeyqnOlx8a6SA9ho8Nr
6VI7RrgA0OY33huuPcMpTOCU+M9S2Kao0hAv4CyFKXaaaB8ryOyVSzo2Mamdx8IT
lL4J66C5HuUN3XD5JgRszf7D7hJw+Gu23KJtAIrLEq7bOTUmA2DyagFoY08LysMe
TaslPY11Wvp4EwvBfKQczLig173AAbHjtxbPR7i2wLrg01X3vcwFk4U6NwwR/Per
b/32ITxFtqSmfrbAF0hD5w2FCbjgStKjCNhCIZf5LPJWB+1pfFlZ4UNRDFStkBdu
CtgSrZQWIZqSbO63QRJurjWZ1sufkPhi7TWg+96hdlRAuJR9m2RWg5pEjPsqHXt1
Q5qRUCyZjXOgRuQ69h2QyHrYVmtcYAplCIjAi1xJY/SHpaaQ8JlB9TuBPAuGn/lv
a6JZBkyGVShJDJ13TRKZdbH72xGKGbt4weITuvVjxIvlehwqsilS4XNI6vUDxMGz
sczwFMl5ZAxAG5RYxY7iJ8A9iVN8mz2HKJL3ZawIFGPtwWyFblSAHy9qNT50ukXF
jm2uukaiZuj8NW7ky4aL/pUpGP7qVsJ9fofjHZf3JoFCo9DOUJpEC0EZXq0S5iZC
HIJCf3EOQWcDq5ddPrgLaMVSWIOjoXtj6aOP9H/ZwIMOPSSGae8n8QP2tU5ttFHq
1OeILb+YhP6tDfOTPXz0nmjgX4MzBjLGQlzidL8cRDco2isfTYUZtuhC+WrtObY6
h+Q5ByJw3Sd1NV52ZZ1cK4uydoZjg82oXH1mX9G9mbnNrQA+fcpZnuK+mOhcy/DY
jtlsypdVZ5kagq1581RFyolNuHepvy6yDiE+Hn3BeYL/2VfrCZwOHi3X/ntiUwNp
3k0aVjeZMiRHL3Z21sOtsierxiLa1/Qg6Lsob5k/jTmWcobqN9O3grxYasa8wtBd
CieQ3j5+jiclRPWdIS+lcAvj2ypT4VeQVAufcbRCBV0LBHUSuF9cVre+Be9cOAY3
y1SXMtI1G+RbsFTOhFvJjLpDvEA+E24Bej2e7QRSdzeHxZpdWYqCm42iFCklNTLO
q0zm+jNTkKlbib6778a668j1yimcx3uQu86Caov+UC7sZKHp0h+q0hti8Et4x6XI
PxngyVMmNOs9ISauX+OfHQMSZXxUGlAwAvPBzqQ9TjzcumA/ErEcsrTlEdBN5wAA
p/4UyJKyBQQ2D6Q9vs8odEZHf5rGeNZrkWoIYkW2UGyxHSqTWdf2xtoEpPzN7iuM
E3s6zizg1MBQra1uRMzGb067Ulw5cnOIxm5XJjYaXsXqNQZL5HHozK1iMAHoBpTE
9eY9ix9L0+vtkr7OrolsKlZ+pUb+b+/8CLcjaG96wzC3fD0jTkYnl9OAXXy1PVeZ
30e/O2uk96yPtcEvEsWaBVZOgsRpKb602zcsQNeoeV23AZQmENCpXS3x0OHPXDfG
5nbKyvT+5hKwkE7M7Z+FhNMZAW0vVMKMQu+q6kRxE68vmqBwqyZBjFuoR9sThG+y
cKBuPso9OcPlRqr6z8Q/2Q7fBKu4h1U803hP++p0DEclJoBluRRlSLE7LWyg2UrS
bsTo2gE7Ja9UZcm2mZDatMxhIFUr8iEBY0YTCoKNsrKPrQl3+IW6NXR9gerypKVg
VIY7N95jOe4jX5Q6hAYoRMtqwaUvMQqCoFd4T+U0BwWIoIefsebzhWtqpEasvmDl
dvMaj4I994KSlRXiZqbc789hIKT7NDC45Oz9wL3GUqwBAuJ9wDflcsPYB/Hig/CT
J1HGooGKmN/77WBjyPbmTk77wRJjCgdLr080lNJbCdy2M43QHJ+gL0LHhERaHw/P
LPyorpg0WzTA8eVqEHewd2jYiq3mcik0VyHp+AJ1bPLoaTDG4CfoXeB66nRARouh
gpbsxnXVy43KV/+mgSbmRP1LRM2JmNBRgeh0BnM7kPTqM6NzbIk8X1bOpQXgsJ6E
nkh0eRxDzIY+UFDJeVkQKOhE15DvYd5SjMEgY1Vue/6qKdu5AfjyBIJ94xqVb3O9
WRMeWNpIFfcsSY0tPAp8Ko8HFedHBUhh/KHifi+kETkBfbKaanAfZLoW7Ka6lhD3
2F62kcCAPFu6+PdD1aXNbScIoPuGq2Ys5a4BYRbLaLfA++dtNCCv1G57IY0lludd
k6PzToyx5Jp0Ehc6dlucwDn/DSWD2rtiuVnbbD0EyamGBMXVJDzx0ia8GF1ksSEk
zrSRHop20fOaQU6eH9ALPt9sZSpo0fLuhi98BuY67ngbvKhSUUE/nG0Vs9/OEqOw
mY8BCCEjXvH8oj1HSVpn0dON+iEXlNKkUbQeZW2ho1Y5NnOwPwDiswx77cakMext
mqi6WBUfB41nLQqgFv/t6RBMGJD1WGDmqk8mAW3ymE0M2duo3GaknGEtxN5ghUGG
DFUpmNVrwTy8M+w54gMGhm4FLIqNMQkAk0ezEqW8Ko5KbqfDxcSb+vZ/PU55ZiWX
MAmPKBVA4DrvgndhUiVjpzkArA6L1EocjOM3VY8wy+Jgeg2VYdBQt+OWO9HHlofF
R9kjgyxrH9ZIvCAyCWAZNcXlXKO4kTEXybjN0pQj0gcNftrFZVkoIqqSanDCuSbH
OZhWV7G5Xa+7YX2ywVlQ0YIu65IM5rSFXoOnz0ul1ZKSJKSAUteBzEJTz17Yos7x
9eYEpdZ9bi80x7XVd1g9qUkPPd+VadTFHChDXrQvoBR9ufXEj9KCeJedIuKkJiAa
zN03AwMxAJLWX22mV+WpvZ9tkErFNA3b4Vg7nH1h9Ggd1uhr5IeoP+tzxPYh1dez
/6j0zitlNEuTq3KcEhOUOzKy7PdsFOfM0QjzPJP4KeJ2IjuKgqmE+4oWjT2vko/Z
8jt3eB+/jeKmBd1OTVTUc3P2NB1DJyt8EEg7O5gWgngowFTSx28WnuHyCRxLbcDn
J0Gvmtz9OXAR+D23ug0XrCE0yUDf7QDrcVrzwCjp9SBljXRzn5K6fySqpNPD2762
qR3TY/N1rH35tYcLuTtD6Z5Auv4t9CZ4LMjlYAIqltsZMHE80caJxnj2xVS6kffc
3kjHq71M7BDVZ3+MmLQzXABDAFFRshsh00Z2THw7/OJZNudxInx9qhy3fa7kKL73
kjNFTVEhFivWtF0OcmrHfeUa7V4K+rJJXD4knm8V+SgHtd16gy9l6gv+Mx/apLKz
1WOI6vXUkugkC4ZG/tmLJ642060q9RJtu5CJ45ECMMb3xpQf3l7ad32rGPac3vz3
FX1pZbeAPshTVdNiMm6q13h2QcG+3S5QStjoQ0mSl4qOyeVX1xAf8yXg4PYAm4cK
f+lvdpuUCExG2C2h02DFwl4rOEmbKeHPASGZBQ5M6Eb5Y80NtGSARoAhsL0RU8kK
HmYq06OWz8DM/NApXIh0EEF5MFf2ooeJHfvZUtu0nZ13SRmxm87/8DQGst5TWq1K
gBui3Y8Ltb9wBLvdIHW8hvgnmvWgDpstGggTIxWe4S6jyT6OEk4N7zLgk4+rDBNR
zSOdf3BkZirR34zT+6vLnydDYCejHMObsXA3CMgRMdbskf4pGwXXwpooUQpR817O
aG0a4KdPDgeSLhdMbYm+/I01Ieve7ZqJDudYvxFuO39NNBNoh/CGbIgOnJ4YSMaw
s/D3ZD5FMyhyT7eLl3olWBXDYFlI4D+CZWlCvK5ulx4YexB1AB7iiKltSi8RgCiu
90QueF6z3S2Bjz8TnOv+mDEX9lIlZaTyEq/9FV+clxbb2otQhIvPvZigR6uRy1q+
Q/PnGp4vldwNgezU/+ZvjOnkKnA5hpETq6USkOmTEBNlOEnmfS4f2NVDIvlW9QJu
mCrRUevSSddcdmzXa0iBmQCmhWfcCfMZO6Iq0umj8mcqRtw0Pv2yaaStYR0dgaUF
zyO9tJbxHm+x0GfH1XfwDNB5Y0xXKTjrB6WPyXd2MjJMJggIo9Ac/Dhaqh4It1Yk
Fxf5rBWEE1fL9/bdSAJ1OmqrHHZetsezNcpWJ+A2JbrOdhuaGFenbfGkWhfuKcNc
kROb0AnFQ27U0ZG1wRSlJEdQQOfc6nzR7ZYklO/gCshg0vi2JuKOX6wPXAALaDRy
de/AC9lZx5tqsvw19Do9TK4qmpU+ZGfezOnzQl341zgaIDrgxL39iiJ8ktOOgtrA
vu2a3T0Jc8feKZwUyPF2xXGHeLwMd51nDVMg2bHbuL00EK5oJ6J1Qb4P9RpoHkiG
9CokgTnLrBQwmS2XSgRyKYrRzsf0YmjRUnzz/oazOhsdj4zFn3+fsbPwn/qKv8Ui
gJf62dWuDRkNrwSd2LBn+7mcGZ4Ioyr2U0fIJC0t95xPO10vhTtYTL2dZV8lB51i
8XLz8dmSjfDvtQNv6qC7X3XHzZroZhbzrS2wJTXMFO9egW7bhPvHe2MxkApHRQcg
dfx3wizi7V6i/8FeHEaTt5T3huQYX/3n31Zrr4rlEA183hcHlRHrhO6a2DcKYwN0
/r0BoyXnWIE5R83RdxvuaLievgIw2BU3kyErEUS39oWXxlBCPv3/YRyXnmxC0Nco
2LDQVaOC3RAyjYb7oxaUdEeSIDEtmQtEbAGkmnRPQw+049J3pCitpHrFmi2lMfk/
TZcVnvVbepV8oZdfpyIDE///p9upLpAgMCwR6oCLzKPub05BY/k278ayewo3QF4K
csn+aANe05rvkUUJPMLlbMlh3jW5lOTo1sIlxTPYA1Krm/kKb/fnlKosyBfnnLIQ
7gwAWhZ5ydE/4oBnT4mld3Sn9lSffww8nJ/hCjHVl/pyTA5wxCjYHkAtXl8ubizU
hceKCRp7fvbknbY7UW3iRGhHJD/C6XTaAWKldQqkpL+GVZZ2Z265nb6WKup3n7Es
qCg9Zp6QtuSx9wC1nhoUkP8Ul1uW1odJXKpu8dO5vhdMipg7YA8FFgacaMhRd8oD
FMxphlkrnJH2q0mgcXYFunlbNygZoGhNN/5ilI53YjbWbdDUfM+Oau/aziyT7EXx
1hjNHwJD/QLx8R5RLMfvsYRMaL1JWLw8ogSqqCRwphbOtjTCmf+umhbfNEIE/m4b
7sJ+6OeR6NVm+8opgzGsgmUxxW2ZMsuG3KAITQHO3o2DpqUhD1zPH/GyB5NJsiAX
aIYsIjeQzul+8TvCSiRIhQHzTrvr5yBHM8YjSt6c5tPhbXEjCIFSKDW5i51jL8lw
NkFCzrLU+jKQZ0Z1vMRnYUo/82hvZYKrAm2TwEHHChSd+zsfOnh0meFFFz2lvOZV
oTf9/jOWqArqzB0JLTZc8a8TbUToy1syP0Ckdg3KKGtRE58G3M+5jvI32bMcGQ9g
5uzF04ZoHg5CBEiNcauuYeIx4KxZpDrxNC4RIEmw7/lk86+FEeKhnsw+buDPJgEA
hZI1ZgOPAuMHzu4peEXlzL5lTLAvhCQspSv1isZN8jT6KL/wxGvI/m1oRTQThYSg
0L7brOYku85ZQ9/ryXjl+OFSK7gIU3pOdVXfRKltxZpQr3fw8aKZJsNto5NBmvuX
k9pMLYAM3AGUw+mYY17b0IV9Zrm/HwenBLAqiaHvSVOPFytoRLJggRj4RqDV/xmP
9VLK4323mYdb9q0IH+NiyDkCFK7C+Y7zWVeLTc2Ru+35RZeSlqMZctjvVJms0xC3
GVCurecnZdaDgOUErCxrOcAnRFaatd9qwZQrT91otmtO6ZHKcSoCh6xYf7EuyOrF
Y9dk8TjWDDLo5/WRh9+Xdxe/S57JSgc2R2M4wr/jYT2RAmOywZQPPaKSVlt/nQ7E
3eEKx2bNMSZbhlmyxj0eRbwfopLivrVyhte3oJdMQciWThtkoqNvCfQVyFVlQq/w
1ssZVXOw1XlietHtUgbbqPRXCY7YuWhKzayZnprbLf8OovzhhOvGuosIGRd7Kq+k
d8IpIxowqMnhAP6xhvkO3URVcXfxt3aB6NwkZ85Av+ks31O/jpLOT0PmpNStuyXS
Cojf5RDs6p1fMhgwl9FXbgs98ELgjpZF97G5IJQMwZS51gsySAWylMSc1xsptwCV
BN8mJlLiHVHOAshIdCxI0mgY309m28//H6bRPbdhlCOQXY1HGJbdC92hGHe/jtR/
YWQ+OZ7d4X4M5cKNOqwPA1FpezNe4eYqZikEugtPkT5NgJc86G7rtja0fvCeA2sr
kTa5b4IT3DZmQf0s/m9a8En/3J9TegkuHTJ3bmvJUcrF4CaqDCe5WWmp26a94ks1
WNMI0HIOevIYXq9+Yz5sK9R7SB9yJigwsoPJGJe5/H8z8vUlAfjWYu7Y1PNL+wuN
krK+njoICihPrE6r5UghPsgMDiFdtPDipTsx0JvgSF8XwE0DRvP1B7sT3WKuyMjt
RjwGHJBoL5Rtqit5pi5MXrsuuxhOGRXOck6TcA7dgzwSoMlWuCvpYaC2kQgt7fXc
LFMnAZBVexJmAU2FkUn+iawTPtxE97Af/UoSqwrGAi+mutHQWktRaUAmCsSYeG9Q
Ar4GAQcQ+dy/wqae7+XLSbs1OlT6lUak9Il9Jv+kyEYKK0x0DPoIpQ6PwvI5PG62
YoyrGQ1djZJebqscofMi2H6e4ioUnY9tVv2VgTU3t/qCXM6HKRctE8EaMAwuvSkt
q4I71u+PURE/ELc6wr3puIJD8DiCj74Vbbiz84KXika78A0L+O69PVffXcrdURh/
JJ9R/6C7S8QhYzF62uDTN9ZrroyKBFH6fqtjrCnKGynSIeyCR7uBOoTMFeY/XVa2
4/O+o54svc/glrnXPQ91nr9xtF66wd9GOJWehEMfHcJIOB5y+pI2s7RGkgzjVZAf
uUOKh58EnpgSUbOjI29dVRJEApR55KdBEuQAbMIdJ9O8msGSVOPqzk5wdARFigmz
aAK64WWBwmTCqA3bkwnAVEnTJB4BlFKCb0sZ/3XEulpLyKVUvnEQyDA2sAO4AJ+2
vwwU8DZ6KE1r57w6bZzRQsMv7xfCzUPAOxl/DB8txx8RwryW5zaNBeAwfV3X3eHJ
phMXvSQzydPxsxi4fKv1I/RpRT+jRRoTjbMkb7LjjNBhejrTCJdguwr5pWNDs1fH
xUHGIUlZMfFlurzxJ0D3T4Ga9vkWXVnNL+BLKxZZlOeA/fM32rbEw6MjL0tyH1bT
3KhFFASLuK3C9JESJOnZamtjRwGpVsimEc4hIiBbmid3SWiHxisMxsYIOnnqj+BN
sCNu2GHpZkVo6mCJ0IKF9IHn2g0YkqYhwZYw/j+2GhGuObo/EdesdHJY5/TJMEFu
QbHJVW/1Xf8PrJ/sAInlcbXHQncMVXWiffSqkBnQ3iOJX+62wmPWSuK0RVKVDf1U
DVBGAozEkfAJIj8n3gaJDeN5TCQp1YbaUOhZ4SkXJaso/UfoAFHmBuOtqzZLK2a9
BTZIZPjwmLy0OnsNupdwkeUW5NKxBaLG+XAfLHcH72FnFL+22lkbhP1US5ecs/5a
eEV1BfSyRUVCKVYO3w8NdS2GcwOFhOy0oNd0tzwEmPSqLOJPJyMZ8R5Zqfdfjc0U
X8opcIWl4MRHQsh3vdRPbG74xVXvVOD+EOMS6Zz/qosyDatQHWNy6Lh+BZNnWxOQ
/T/1bcc/2pIbEbxeOCY8Z8h6cWnCMzqyeyIljBY3j3ipt74jnawt+cxSA42u1l8d
JE7v66t87CILYNmodOjH2zOw0MAcOftndG8aoFv+GlgLhJvBsQXEJ0R3qFwrctun
pFkrhx/NkAi6UAJjd+otgJJQTMe9OFmAErEUMVh9fcHM4dTzTOJ/mb+hiailRyCn
WvR8PucCMmU0qfKNhIXPE09MiJEhVYEvMQyBMcpa4o5jKE7DhMPixOIi5+2JESu+
ltzLUOeqaLDEPST90XeMpTNexi0otV+gf5JIH0vIdfNDO+3pNgmgIZN7Ah2uLb1z
EnijP6ue06D+9qQxLIcnoNQpXHtrg/43IKOj2F2N/WQwYIcQXOLFc6njA7qnst/8
yBF52XmItvzfakDwWOxz4As+9N5LyqSQIl9humWh94pCcg3tGG7aydEkTK2GMpil
Li6urg3uXaiLXI3QimlS7Sts9k3Wiflvj2LklADSADerZQ1DngBqOmwK7FKRM61F
8BPaeT549xLIV02IbZQaOPFrLxuYgEY7HyKASTVFxVz9si2h4PbYxKrumI7Caxy3
ISn6IIOruho9GA2bIiGYN6DPLJsw9dCigkTq46kE5zP728U4VU4E/KiGWQJbVcWZ
/aDhKOl1QqpGge+qNJukWi50qRvumnkrWrQ3eNQP9qwhmR1vzBXiZVPWOeq1fHPL
evZGw8mbmgxtjkZgFXoy6Ak/xjbrt9E2iWCsdCHO48NwpFjKOCpBKtXcxYZMCXH/
ppK8nune2WMQApo36a6TjDblR90/JJh4q3wdNRhwZFkfQ0N+DXn44T/iNVpIDU5V
p5VyFpoksaIkaPpYFx+fbYeN7xOBqD//cQmsLe5VQLifpcYZ5grzCBjdFjeDnN1j
Bea8/qNZ/6CTBnzliNj7RVZ9cXByel90v60vHw4sTODE1q5jH4p8m1l23sotozN6
Kofhk1UkuSrwRIEUb2+B+bN8w5rC/PuuDrzTKHJmU8GX2t2fXd6nfD7unDcnFl4k
Tuqlf0gw2ip+GPuMljq1i+6mnBTyzc6Wx8Yu1ZdpDcq2zWfItE+iUw4SE6UjyErD
k56nRELyJq+agjM0ZuGIin5P5GymBWMtlgRPgHj+YuB+IPi3GAMOYOlCyXF9MtJp
ArNxWfqxA6v3UcQ+rmRdfTADt00LgRSGZUdMC4ZA358Kg7unn8NpLYJt5amKHFUG
tPoqKpneYeP6zT3HsiS4J90hzBLtw0dyAzyksxvqwHjuGIJmB20tzpaUUkCPozGk
oDBfg5xmvJBDqAenm/ZDv2P7Wn1y1P316YOUAjw0wUnGE43IBP6OaoAJVgFsLKv0
Gc5r/MqYsZlFSQO9BC57lzrBzC0PpSPZL8Rb6OM59SHb6LcBID0XNf/rQe+1vrS1
+Viuc/L6j/qRuLsfj+E6b3pJIsRJQ864I7JKCDErkaBbqhUjkzJypzLC0rMDXcb0
oDQFq30vd9Aov4LZID9oDo7sUM0Pn3N6iLqIXrhsup68Po4nL1rPuZf/JsQt3r3R
mXTJeQhYvusZh1exbfQVD+mwqd9PiggUNd0D1eVSgVIJqvdF1auYFHhXF+Ngm1pX
LpFQgpswbyGUl3tho66HXWCxqCJ88r6P6FO7EfGJRozcwd3/E2dtR0hkYTToSrKM
t6NMfDLzVzUSoYFY4vfh4Cu3R/0278ADNsE2oGrT8184g/I9vHTnAJ6Aqss+G60a
3qJwEChTjJR8vfHhI1P6uMrYsvGV+tOxzYr2xiihs4O4Lgjr/J1YtmwgHFgqcX4u
gPIvx/VMrsEXrQOBeplHO0G2Vmc0qBnpk5O0Nvxn2oF0eTcjZtif6xmMQMsumQUW
TDU9RyfXEA9BKjMwMBUxrVNf+b4jZUEQweepd/XNCh3aXVG98dWyzL5nQTIOt18x
tbf0tdq+jyFLGu3hmlBIc8OVbNKMBSNX9fgTQL5FgdLEYwbIbYZNIISvJybNZr55
oILjXGe19doKe5NBkyaQ1C6Rmmfhew1i/QMsK9EnvSyU/mhquN+WHe8LvxV4CpWo
oDM1VU5k+9ZUjPlO1dOigwLEwZA1QgZbvA0i2xoCL7UKjhFI2fELMSJnKWmyyYXj
t+SmMIwsw/mnnX+rOS4HD2TDVkEDYZMTNFplGUM7gboSaMiM4rn609WhvIZr/JYd
z3EGNwb5zxvOUaquB8oe/dvKPbX0Oufk7hVxdn0O7etFQ1JUDYlL/vyfYMKBAHzG
MYkcMWtAR02R0Je/fw5kJJfyrAtFlcc/9t6MdSGmBiVeHeuKxlZygrkx3sv/aNKQ
6bIbH9Fspip9dQ73XS9vldnRJ0OsliyFkAUKtnM/+8ujDIkX+GhS6xioi/VL8hRl
aPs+D6htOyWxZA3Bu/VqO92YQdzTuHUNVEbKaEyifTCE0lm80SplNVuNIs3yWnXV
c5cofVoVqoJyApMNCyVxXeBMsTru3j7D44bmzLSLvvHM5hUGzr5MLfsf+f0LzcmO
wD1fMP1p4LXrB7YzQcdE/qEjB5gzQFzHVNaoDYBoNt99z2cS/59VZaZQ2wWIc3mH
/81RyBiAyuz5xWSns3FRHqn2Nzc0c5aW2SWnfL05jJu052W94eeMzIYvkf4OLXht
KS8N+NyCOEDy7lzVoWMXlhtrRFzpGhodaEN6z4uRmiCsG+1/VgEN4yTk9uql91wa
GZEXVA526Sq1O9AowKgKBosRldNROl/ETiaCWxj60jRukfUluXhEmZFVFJlaSahd
ub9A65zOSwcKIJdrVe5XjMrU68d1SvIEKIC9VF08pxKwqkR+vRoTDq4eUmueUWzI
sp4dlF0Z6cdh6/xovC6qu4DVIkrrDSdp2m29BSEewatSr3a7K8KqDYCFWqRHshgD
tGYyihqdlNbAijwLKr3krZHE1KUzqPJDDVc/r18DFGO1FN/qV0wW8fCBlnxloP6Y
o9zKSs1qfq6BXrKDnYFXMZUVOsF3l2W5McdDjNHbuTjx1gv+mmhNd+n1boSIEJyB
bXVoBz519keojlpJkzXjlxF2VgKkmlmA/y4+Jpza4nZG7MhV8Pv6Y9uoQXQ7hmv7
PGPPAS5yQBh9yjOuZjDOoVEExmP8UvX5rqHtF9X11ZFhQWz1fIpWrLpAhIXoM5jQ
k2Q22CdsSEgw7bvRqmMD4WXspV8keCrAocYav9qXKwCNKBSC1bIje27uDc+7eZcx
u0UTJ5YMzGd5LSUhg4M+SKk++ZgEN8MA7xvwjDnmBOcQLXVimiQGbZDxMAMfJhh5
Ryn1GYPj4II9V0YtjRRX3Lcm7w+WJc18OMgyfMmR8kzCtv6+cVu4Wiqs5feqSpuN
KnoB41bhY6oocSe5JMd/SlqcI8kf9PzaQthFOsFwDr6Lu8d2XE9NDrwIQD7NS48b
1SxH4COi7oIPK+0z9a6i06sdNtEHmYtNSN5HauLYfi57gi7/4TXycPFaYiwqNIe8
UfgI5lvJdsQO14oEEhnFDEGCESVRS8jB7sBZ5Z4TZ07sqfZi0PeSdG0bmUrxCO8M
ErIyiNzGhU+XGxJtAYrheBqjpPguE8VQ7DyQYE4kWPcDgbbOqrhqOcfhAUCnvhL0
6B3DAF2ye2FFCQbODSvp2VZaBlaR1V/jDwkQ+u4wcJOjey2VuCVFs9rvtMCRVx4t
G49ymTLkdDOLEJttDkpJMLzIQPOb/Ptwxbdti2SkegKEPafZIqJBgoGt6ppfsxyd
JO7X2lCzjhP1ZDAJuITDDyChvFFa0e0eX5YlAfaiPycwRLqyrr6ZPRXk8teKm1sG
isWfrlq6ClmpU7Oo17pN+Pfn0MJ+33YzTDAV6kwhOC3cq+Q+I7EbgguiaZsfRqHG
XBdDMGnm+EnlGrV/y+TYo1uAHChEFYtSfzEh5AvHnhCZkosRf6eJvN6Qqp/7iErN
frrUVwRiEIgGlALSMz412gXR2rIcZk9MD7Fzo5c8qEvluXuWfvAJroI+E7XNdqZY
K7IvrwsUdHLZz/LM0b+dw/l7GTMu7h50DIO4oiMH9SuLQLs3tDIfXpjjhN2CKr/R
DuMm/Wbq+sziNxowWe9kR2l9xC7ChYBDCfdx15N1JKNW5UA2ThMiDfVlMZKoHP/f
rU6KDM2WjUbDEbypeGyul14sqHcpwlnwJdMFtCOIZrr8Ej/TZ4NcyF3TRHShwNYh
vgtNLSq1+ewaCdcprnpkrscorblS8IMm0cl+0keMBCTJh1k50urqyofbmfOcEwVq
x5dsYWw+CXwHV8fq5JN8N/QYY4oo+0TdTGmeZV/MUZ7ZLVlUvr60TEwTplwgPa6q
rpbAL13g4vhi/sZ4jRJG5FjkEjjs1PXv8aUN5wxt7bh00cQCfXnTggy5y+zXj4l1
iwtkJFRxlezgOeyyVYxg+pIDocy9Bn/M0z10pGmV0jQfmfY7fs8NUH2uf2h1VXsa
6nnDdTR1Dgytk3WV+Y3IHLbynU33D0KvGS6ThLFKdvwgqcg+DBP/haqOYvDQSUlV
nfzEh0pXYdaBk8gAd7GDUDH7IneVphTtI4K5Wg5fA+fRQMynyIf7RWI7SMnj42f0
5v87IJZyUob1P+JgRVWjvLmTOLUrDSLuZOO+ScVRO57b6VZQOdv3f+VsIiecR3bU
m5oFTys6TQ/jX0NaGLHWkI/o8LaJfxJiIYgxHoZ5xWgqiaRjUFkZZjFeSk9UzGbc
bINXENxYpOjFfv5JthNwp4//vKIOCZHynVEuVQdrsMbmus5K8rmKtmTT6Ph1EVhD
DUcj+q6vigu/+E2wT3ADM/sE4SJvtM3JqfXmnX9RMEQibrACcfcTn26qAOS8xamD
s+FpzYDT9SFhSIiS2jDNabK7OV+7bLZo3Lsv39rXz3+EGMfuCCkm8tuNFx8P2ydg
xvf8568FvVUhznEjGRJU/UX3aBU7BundSQ0cWuP+0hACUT+tc9k3251AaoDJmoni
UyIgVfJd7TTRSzu7gbVDuop5Vq84/6TsOeE6gMqBUocBC0Dh8JogCaPX+sQHM71k
j7ICCPSyTJO4gX2k+lFs6FobaEp0COw4gYZ//AoXABa/1EgEbv4icbTuh+YpZdJR
3kmY4t+TkSZloJi9X6EfPkkm0Lv5gggL9aM5+GcZvX5bsRzMoiK5lFjo2qbTJIeE
sA69UKevmUGHeDMr+wND2fTVPQQSfHOjZ9ADZVM48NaqTIa5IXoO8dTjV7Oeu1Wj
vzIt5iN5bDN6hjKdtU/D3lW7UWSMSGOkPrC59E3zzK7NnaR4iFUiyO6ZW8PzIVZT
tyf8rx0UYdXQXO+2tOY4s5VRBSfl3YVpPOgGZGERHHgBfu+PnFSQ8ftqjeBF1T2/
rhQizBQRmRXwErpKkfHg0qrpMGyrSopYclNS0ov6GcZHBpo1EBwCrguN0llcYQ70
Maw4aI0NTAlFmeJHVR/v5NXOI8BkGtOOdd56KZCLS0B+aWb7Yo84xZgDry6pvQK0
/gPEGObBOQGTKzxJTU/xyM7JPnwTz65iAa8SpBipTZuG00eo+enXqDWXCXJ5XG6r
wxEehjo0nIQ4EIKMXspnv6DaXeXd7Wt0N3RY9No4RMVVL5yzxPBoeILBSuhkP7Hr
btm1kNK1YBOOeUPN7P4HD0suZq0xGbSLlEAyNcAfEcf73VPJBLPzHhtFjLHPl5ug
G/Hi0mKGgERdMt9Sy6b2ahq6Co4p/MscJZx/AW8mAto3G2/jXCEOJJCTN6v6BZx/
tErbhAc1fBhbfrVpN4ZN/UXH65AAbOr3VpjymIJaEoYfoyqI0Dh9aD/wGFmeIYz6
ZYLQi+ZiT7GSHZ04z5Bhz9vuHCajSUtTMOdyag1j8VjiU8EITDz9seedooYubBgK
TZCZeeMenjX0naY4yEXfktTqEXIJ4OKA6QR5GVR2HWSTi207mzvMcZ1XOFHz3l5N
1mqzUxrtaokSc77zbMUXo4m+M8lH3to/Bc6s8L6I5vvRv07S0Eb7RxMp+EOkj8A+
KkidLjLuCyj4fOiN3VgfTEXhNy9bo7FAn2f88+8WpqJCPEpqpA9g38WmFKBYtFGA
yNXRv1UfW/6Maf50wxhdIORPppbeAWXGK/9CxQMEJmpLQfa2CWnOxdwOO+33TP0U
3slxDOkyxMEPwpY5QRIVZhGJ/7qudkfaeYZWxlA93TC/LSYz58lRvKC0DpIMgUb7
h0nAg8H6aESVPTrY0CUgBB7v3M0ZbjG2LA0f9fiU+guKubr18UHaWQT7q+GhHeLP
6Sf1XPMk+Tx+i/8gflXi/PR9GYBI7i5aMJPvDacVG25fq+hEk2SwONYEkf63Jfnz
S0rm1I6xe5g8fBv9IcNEJUCrpVAQQL6L4eeyo3iv1uanFPXB/VGqJ66ibHuwMi8+
BJCjXaDuVUh1CN2oK4sq4y/w/yYdS14tqzspCORG+kI6v9O8Dezpl1Ie/ug277bL
TmZZeysD9CVTcVFUe9Dm2zI1C5EQgSpQQGz29Os1sJo96oxB42YW4rriIxUJUWrr
4Zpyzsfk2CLmwdP92FtuWaCbIwjupdtCyzIppaqs0bqHGMCyDml+40jE1dpAEwnY
wt48/6e3LEN6HN1s+XIt9sIAAWBAImhlaFSPsvcgxBghON6E+dF7hjSXFncY58gI
ClMGgbsMSzOZdP1Rn53KPHtb9FyD5UGREiggf16lJ9fSsrtLLeXWjYutCk+TK9za
Z3T+kvYBjhwdLyPTY7YuR0hMbtSg4AyoamPCyjS/j8ULUwQDCX0+vSf379cnjAUp
3MH1iUO2YFkcxOY4xERtQJZHDdeE27PvSlK+DWPCHSVCWmhArwH1+RE9XdNvvKdj
v9oGyy/yU4vLBhdhq4Yy45fjz02HJV0UhaGoXqgpV6hGZaGbcY/tiLpFIZylFaoF
eCveadAouu86t7FVVHAwAbmDpdI4JBvuG4MS9C6jYPfPdilPv757oFdKqAkI6OJ6
6DzZF8q1G0IChe8jYz6XfNnbKltBpOirpbueamhlJI7TfN6PHEs+7XPJn2WwvVzf
rX9J81h2OqC8hbSE145Jafx8Ow5/MDT9wuNVV/7NeTuj/Wmsu2uV88WH8Z5JHSUs
7ShL2XYp9pQPBl95tXXXzaypPynge+H3u10SnbLSq6FYz/d8/xZ4OetcxjXe6vxa
1xz4dkfsyW3/flBVVhM8xV9qWbra5f9x/XtpxhfNAAJIlG5zxLoqD2QEfaTLZAl4
QZdVMkvqIw8X396zLA5y6jMoUHmX/SJcYjlOj1H7mAZt+hEgANjIng9BYP/PUqfN
adCQ+QbatpNzqBvhsCUyEajxNhzvo9Cavg0fA9HOGg8DU+31exTcroic7362CpPC
jwOSPfUWJ0PAYvRolfGq4ygpj8OhIjNzp/PUGLsQtTpeOxQcSHVqbqdNHC8SLZkN
1YiE4K1NLdeq8oJ+EXkxjLHNfhkfEW3lqa/SEbuEq1BV4LsxXiUoTxd6Vmp+S8yh
ATsvvcAWNZZJNIPrtJtmfR4baIbgEjJQSJ/V979aqzKRV8jWqsUQxbVea4YgIIlQ
riaSFt2GrILsOf6QYQk4MhR83PMHRFEZU2uL0R4wy7Q7qZS4pfuMKnWLDRS+gNHs
wxe3M3ECmL9cEgy2hXCr0EY3nj+A8e4/oPKFJjzlVB2ukDMvBFGIVKF5R1pL8SFI
jEuWpmyzNh20GTZeYAuGHd16v76PJSgOc4BTiAvwILYnjf5zqevFWad9FVcyjOLy
pf0fKvfF9ofMwbCUnXd0/mPoW/GfaBgfflqeAs9NXbzd73txA4hRtdWWKBk1btie
xl94MNrtEP88Ply5XVBc7xoaF4a+aly9IwNwa+p2B1gnsFsyyZylKWiGyvaeHyUJ
L/55uP4YpVBD+oekfM+YCpBnb7g1AyrPZKJAM5QNaaf5y9jvd24mABnSJ0eZ3ykb
kmsWS18cZ7kWbJftpUYLiXXHYGIB8/yRvJox/0fc7UlwNWEyzmab5c5/NTd/Vb39
WS7lUblLSdqfS9FYtzGOZSbLo7C+djc26nwZI8aDO+81xO9RMXEk26LNGzCSMmdM
pJ+RtzpdKeLONpZjKqwOkOt8e7dXvNDLWB2JSZCZxVYRT0hWRadlEno1p3lusGdI
YWXXUjCcq4TyyIzpa+zq4dIUpQioHWQjE9X60P7sdRgaXrw6D1faVmbxHL6iMOQu
J6TMJZJkrcd5POJQ/g92JV1sU3MCqJxqri3ZcPux/SZ4ZQwAceyueG+Olfv53BX6
nVU9gz2rPtXbtdyRjLuBGJnirfX8PvscCSstwKzMtEwpOIdhy6+TAybjKFqTdnhO
T77p8aD25Yy/OL1EqnO+m8hWivjtCgt78ttYpnzffCNxiNQic0fR6soDQN0cIvuC
Qv3WTxAeYqx3mIbMoS0/x0qgS2Iqcwns7CdiSi3YPKAvUE5tpeeJpcRYZ4Wwi3vY
3BtBmLOwGuKRjsZd9Fvn4ppfoFTc3xeDJdey/apnOiKlncE0Py/5w3uMLkZMzjZL
zUQyp4fUoeuebQaGT4RcyK7lXOB/dsKAmxXShJxYKrOQxM8LGJRPcQRBQI/QhqLX
whNeAW4zQUwUWoWN6hhjz0ENUnXpFSxZ2jTRiq0QuPnQ9JqPu1Y113YqNU/fbQTP
yZMORFvhrKVAuYFY3AuFeQoKD8a9AIFKDLz8+dkTpuQjYlGU4C/pq+0SEYtlpC0m
pfxZNcrsunBvIyW0QDEC5o9l4EX9UumgdIZXlokl5Zyhj5H0IV2wc9U+2FPyRQQK
QLCky7/O4e9UIUbyJtwRQnO1oB4KFTCbYlGi6qU4bCJd7XzHHoMDHH4/2V5VvNyz
3cNcw/sWFvcLJe/I/ve2H+arAPzAXbPkV4UukY52C8FbvWTXJtHG/flNcc71Q7b2
vr9svAanuj3+L3CUM6R4roqcgmp/Dwv7sBc/qtLVKAp4KpMGCRg37mgIe/glK/yp
lI5aIwSBGEhuIXWkKkI5aC9NmQVhGQvdDnrQaDPePoILh7l66aTKa6si80wdIwzt
x2CciBUnpMt0pS51gsXxmwsL2RrFYDs4D2n/iIXSW69ke5a5Fxv8kHlCPMmuPtvb
chAlBtrEb8o1EC60tHfdeVi7j6gndufaXqUCzMhnoXYjEzIJB8o1BkW0W1n0374Q
0q/CcoT2HoAUYzm7BoMoMGkVfHqRAW4dx6Jcj+bS5kWmD0/bCB7iTSTDieD5PZxU
k++D2arzd1jZoNneswoB4kgALhUq4OOEGvTtiYWkrCzLI9efGQdZcGAqKzBnYi6T
zlTEP9TRbu1LvxdiiHCH2Mcu4MUyfUVgzqkEoYk10aFCDyVIDJDAXt6vP2GJ8751
OZl2jD2xj1SnGmiGDda6FYNKqvPkZ02bc4gv9qYg94zLM1OEnlFW+Lbi06ZIpRlf
9xXpM4X0S3HzwBdTuGZiCsl1IwqBZdJccSjXdQHtO+eGW1IbmJwTbMrlc+DoBaBQ
/6Z1/xpTyPoknmvZwqCKNzucRJ3kDfCNlaeIjgtc5TLub74u5RCmqSqyHJccjIA5
/R5QapNCKdIi1F/XeIeSucjSGv4SlobU/ucAxkNUZPjUqRW5UPM4kJ8JGry6/akP
HyuD9f6gujXh1sxww3WNLdisCCRNjn9WllAwlUmMRvluBqVOcNkI+DvQbK3ewUvs
Q6LwO8fHj5AP7f8FNwY8/jbQeG1yFtws4IvEsdLl03hRc8pd2uD4H7jStHicc59B
7a8+nWxJXlDFckwdsdBYpgp5HjIFjGgutiR5/but4kvYgT5Bd5cQ7mlHmB1rgFgS
HJgQ4DOh/93Ujn1gHtCWLk5ldBJcohUk5QT9x40NEzvN7IOxZ+KPYe+C7XdVBZvB
0QEqZ8u+Qm1fPEU6+NY8C50tRbsqBRgBUpjqzWM0CSb7ywrAQzG89ZS1dpB/mVro
g2BBCiV+0XR4e883msExhCQQdmlI2V9U4g35mqSit5nLk47ZraLYfDPULrveqdfC
X8ZWBgyURYQqJpj55qTPyTgyo3nBjmpU1W7/EDFx10vgEq4sxhLutWy7LBNzdO6r
x5qDSgtvstcA5d77nPL7TvXBYLfW/2B2BV9KFnRFeH6ZzLI6k0pIV31jOFSGFG/z
4vpwcJtky5SvS8nW7Co8PY8UQeszmY0kUqk/5giItV2aZHsPqDOQxyP4S3dnY1IO
wZDcOvlM1jzbJjOH3afsqLVGeGgUp1z7V8xVumOeQ/ef5AZCSRJVYkL2U3rXUJfr
d3BsfaM/SlevGP6LRek5jUsSEGtAw+S8ZpgBfqCROsvY7ZDA1qDRly7VoEObWyNA
V3V8XPSLpDJxK4Ae/wvUztTzasImZut6AZlUaGPenjc+k+yCjnShKx+KpwFCdVGF
Yt0G5ZjFOyyhdcZjql+EcQPNFJJ5H4L2z+P6JqZj9la4xpNc3XEwBytQz7Pswzv0
v94PcLpv0f/x+BiqYKmGNNfQDXACzaH2dNRvK5iz6kieBxssey6MLuuNLlVboKC5
ENeGe/xpk/+LueVzOTg0UGtTB/cI+O6HTbfP+aEbCiMm2ziyZtGd6Ht3WcL4u3BO
HqkV9KIUOOdXTu+hZp95pDiqBQnCXkbvvtM6Xrd7T7ti6V+EVwFQiNwv3W5HiYyz
bmEn9L6BuFZw0klm3BurVs2HpfBbSwfYA4kaCzDtmO8/LNzjqJQ2bAfrRTjohxlz
A+mbwnlMiLf3/L+GLA/dRbCNDpoB8Y1iAgRK9ZquSlheX77Dhkx98D+yAyJUC1I7
FkjLomAQkd7wKsundkLOFZ/o8QTuE0VXp2IoxiLilz2nflnBgaq1+JDzKbaofhho
/8nx2DGFFg0oFv94nwO1Rj5wQBzcxy1MG5bcEpWyxnt0SYJHaexd7Sq6mcFUjlV6
1C5FInvo31iJvzphERjyPho2sYr70xAsJrq05DbaHxtBTZHayrTSWH/ie60unjDz
BzIdJjOu90zWFwLJXweaCHmrJP9dgWNcvPRspQtvzjuv/gxkeE8b8C6x6SeIAyUd
a7qRxMftNOZyat4J/QS89xxA5OUVjJap4KzKKGq0k/BiaXAYZYpfr6hw0mcjwA7s
4e2UeR0bXcFB+fV7FF3JxqO/qn+AXnPQHO5Ucvn9ykBqtt8ZJ8p8yR/bxFdP8QcW
Vs5hSplPCuSRWTrQdJ6zBWyobuejxlSyFq1n1/tBtXQPassqfW1FkGwdro+DfYcl
rFLljp1YA4QyMR5jA1mj2ULAaZ42sXlrFr4prXVPhv14i3RepPpiT/M57cSJllGb
EPr17kVK0/8oAyMb83hXkY15Q5xKvuOcwZSqp8KiMrm21mA8pxH9DtSyiytmH1po
Bo+/lwRjJnaCaSW7KithPw8ytiiEKwpjw46GKmRTVvYgqUztFujzlnle/J6bIwUv
bplERO06spx0MPjtHxSYVSpVgISLccIn/csjNkMjqV9i6OxlfzYegAFKGh0kcmZ6
KnnmIitBRp03xnngN7NsucdJpJ8DS65CN7pCyiP2rZDS2sLyy+LspNZQB20eYCJ/
O0ackMMa8jgIVTifidz0rVShLPQTVSfxk8CSKnrxEhBwNopXbMBSPq7zfGqo38zY
VsCAl4YvUq3odyzGMZrUsoGWqYPgNCIAkE09IHxQyondIYYYdCvg0PHPH72grID4
3GSLlwWBnzbXD/Yj34hMUbNgiB0hYaNX4EyYO8qc7Uux2PKTRV9YlyNy+dEzJuqp
oEIle0UvwRAz0MleLKQAc8Pd3lWmOm77Vu6ZrQ9nBzE+o8nCbkvnmhQ1XBW33t/O
YPYl7c2GTeSqUTsTNCK9j9A+Ei8OvG73EdwjHrVRGHQsbmNYCNLe6Tv3fK3zgie3
ua78hS/FnKqqk3aE5YYVBrjX6qoc9QnVbIqXCNFFNocfG923jpzOGMdPw+anLgOW
FDnH7gaqg3SuTtWDPezUD20ZUlaY2f4Nwijpm4Ee8WFTHDDrDqN4XaXUjlgcvJTT
Bamc2mtU+V0TcdPzDQgvPcO84/xCnqC+WsQm7CDb1eXIguecaThmRiypPAFpFxWc
4S3kithkPEYvooBUe7nMOTxKvzGKveZ4fasm87sZWtbb/yvEoNDAYqNkCN/Fv3Ae
g1LaDZXq7JvBCDGQSn16q0VAm3/YU9aJBdRfvG7w5WB/56iZN9VoeXTxicXmSsY/
ayyB2vDKygYQ6+ImJ9qrr3sWVFEnDxDkGNxYu41b9j+RnYE7jlSB1ZqJWAR3SDOW
Xw72QDPJ1o2vc9Md9qxiloXkGhvZDOW2xlq0ocrAxdVnp1RHWbFB6Pf8MryKR27f
1XRWaMn9Q1E4kquysONwayivQmNFhg32NfTDtf4noBTc4H/Ut8jFImsQAiTC/L2t
5Uiqavpj4QMa2B9hW7mUCHewTmI1LeSk9YLPYC1NwOrex9rcffT2sPLPwj7EHf+m
OV2lIDtR8rIQyWrMAgE3cinA8uJ5Es7YTEtwWJHMGbOkonj9CRNwDE0IJwi7btes
dyb1ypAUZsjW7XFH9Tw+wYZ74W/Q94NTtrpIbHmBbsF4JjUSowAgTlh2bemJmzmn
fpofpylCCqYYfXuEUWy0KZZL1JwgsIilC/yGUOLE7KFXO4qxBt7Eq5xo5cQucRFV
4OLolElc/7UQrpw7HI9J7ztrCe+jxYV0R9BLVHBigWz9pS9i021YLDbiC5m3MD+C
k9CfdJzrryX7B8O4AUjDsqsuehHolAW+pAXFfL6vvfKn3chwlCLLgGSm0jLjpaiC
mXEDDmUvJvxIl1cNUnZXpZjOgv/NUAwYLZRAHjr14+Kn1+RNHaCqQLiuot2heyZe
igXQYCyADaE1My1kSDaB6OkQRXbeVmCZITZ2bGQF8UkxhoCJpGrzrsi1NAj7KZ0N
xH+CJJofInSUhFv+NMOJH0dGHscUJmgN+ahLVKdXLisPVK4iEBkoA6/tqWPrGuhV
Aupxy+ub9WR+u9FwHaFJLHBOG2hu+mMmEPASpgR6Intapabvtz8IEgti7Srq3PG+
oNr6ZN0XHQ26RQCBHpyY0ioxk84cqme1Taw7fYz0GZvQJnCHDJF0RYVJKPa6JuYG
Y9VezLsMGzP8h4W6n/l3uxzX/0/7LQjLMGTITZERIzUnFugTyWVAQNaA/r9c1yLe
dx0mjK7kBux6TXVtq/eE6+9vIdOKiUS3vvmKHbmKANr+OErdgl17NHIWZxQif9ul
2TbOE0cdbVOKmNkPWXXO2FyRgheZM32+VGgb5sZ0vvHpdu/ip7Slwk6iy9BZhZZb
+7wvE17G+IsI/2VNbJoGcA/ipLWkpbSK5hEZNz6nrG8fKHovmKkkdrHXT0K8YCRg
AYREdPWoR9KupOedMHStrnXXPfrHQpwhXykXK2aAUQGX8rVss40ZECJXfEhiH8BK
zSZS0ipATQ6L/37H0OwOLaMfBjfJlWu9NzWStUQC3yXdoYyBcPboLLlZIiIZfwx/
iEHAVrqSl9rR38mDjF+N+ERdq3ygJ6PvxSnpqR+S9o06xlD4Z24TcOoAu7pe2NmP
Ujc5wmp/3w795Nj1497MhEW/FMOwhVHZcFyPKxiwdHMjuIHwCLkaF3VK17QlVJ2s
39yB9APzsOu5JmD5LW4IIKBd6VuMF0C3eVE8DArgBxoI16fOpoi+pRFV9IoS1YVn
5WnhVPGQH78Uzo/L9ZrwGETRxLGUlNxjtXZkRHklQ+lfZVCr7RFpC3zCEa/PJqrr
q3YUnDbeWGHskskb/JKTqc+4mfdFxjOQvyF0ScuctH66eb+0rzK/W2UfxQAkMTyU
3vFtsvFaZ+9Y0LyH3CaRm2c+2rs4CO2cRoa3gfPZ1jroBV+E7QGeYYUKtNgkAlk1
AnUcWf/A5LsxW4Xuu/LL2eYeh/ZoHXYGOOuPWRbMeXZEJ6yMyB6AR14Ms8zFGKce
MWNNTNZd1/DIPTYhtRwmtu/WzuuDCbib5l/JE1PXc8kuLaFM8UnqASrdPuwzgDi0
p8fphpBleGPaeWsieYqtsu1FlXC+d+ijW1+3XYW0ppbPd+q9W66IUXjw76LRm9Id
nVP0ZtZW4YEao0rZ8lznXcNoL90lxobbPXEvSWOtAG2GelwQMnvlJKeyzaO1PcsU
tQ62FZ/Erzht7H8gTFQBqmuvvmC17B8GRHjyK8WayDPaGL82YzmAaMU/Ho/DvJb2
N9Idd4lbiYid7IY0AYj/QFclQFIGytxW7jPubZH4NocY8IxKoNqaQKI0HlfUEARZ
aF3+dwK26GdWo7XRyKkwebOercV3CeSDI7CDi+5GkUhIiTJgz7d+5apEJOQHndtB
UY2gwJnV2sx8fJKmoTzDEgIMD9DUIqwPYpa1U4FW+5qWHU9nJqJJ+BiAIF0ll1hi
7WU3xU/zndwhBndbMyXdnvbjJMa5EBjcE/RWzbHD3Xbf8cOUgtqcQjgIWuZNcpCA
MSzj4NJvDao+6GHWMiVkYQVRXgm589JMncXTZE7lqETU8VZAI8kGlFCHhJx06EqO
7ar8Uov+gcV+q7PIsVW9PA1jX1CAPGg7CaGRRM2kfWbI4in0JL5dwg3vXWx+vp39
IM4j1Tbt3wfuRNFR3EbodlkY4dwHl4IB4WR93cGE7NGwUVrglJGLYT9riYqkcoYc
LiOAsew6wKs8TpqYSlSwMI5Ot+jpuaJp80vQ6y64IS9ml6+GcvnD1FOFuJ/SoyC9
g3PdJfVoCeY1oaAtmLW7JMvCBq5FhwSQ3oaw9MBNzjD0wg7lynYKHa92dtCLwPXR
XqTUd6dvRdLIxB7lt/VqfmFKrLBaxDV/j0TXclnU1zd26subgmXd3Huymi9hu4mQ
jjxwJK74G+W7/7fg04Dh8YsrlvW046IteOhMH6joxf3GxroJCWxk+zbSET8ZWJI5
0HLKLbtuHcJIPxmYiQoDH0M0eKJRPSCpmMr1kpEqzJrBdLpTJwXinolC7NRgt+6Q
qYAE4Qy7QQF6DJtMVxCLdRZApoJ8ADQdn5Rn9TmO6pmlJvy0pIlMwdvOyFDBaFd3
XIK27QGEPgt7o8osO/opVkRHIDL6BoWr9g8fJEQkcXPbAgIa3TE2fkHzKhikwQBb
lqw7UcahMxH10WWPECu8Xvhtc4MJTxaz0LWLyeEoj0PxraOlphKnuf9k5xnE4xOD
pOrCwI8yffaOQeHTR39dRwLQYUSwvSsrwnoPZKvihk1xzz+/OxVjX+OkHidSmXXR
Hu6wl/kaxL88U7qHh/D3jmoVrWF6QNRFoGgwZd6VqdvHb8mx/NCbi99bidAL48Rv
CrfYtMewQC4w00NbpvjxQ5LuV9cmENZiuIOYwy9tVM1uQxzhoQVgNbCnNNy6SEPA
uLfMowb5bBPoT/iHa7KnbcouM4LR+qmqHyTvr0wtHrbMjsity/rraMFXiJe2D2MB
RLRCEm1BRd8BZowh68KjoTyEbHdcsqGJ0Y0Tkr1rabOqzdOooK+5OPqDwkHVPgYE
4IVJWnht/SphDcZMba1PHOF2z3ZSeA1OHwKRZXNa9Mo9sMiB9RrL/CMokHwfQt2L
pJTvHItmDbNGviiFK3St9GLxHmEr7nr5+KwfbT3kzEJvd/Zj7HIicvq4r+W+R9yy
qdvnyUi62xXFkzpFwoVqNJAxJ+kLbOSyZFgMQs6h40GfspTtuZPFVcqIqoZ4LmRu
Uq4U0ih4EbDf8GmblYDJ9gB6hE9VwkEJTY31e2wIdAtXoFlOSgeFD/Km2d+pwLfF
s2TvCX6SiDob/TzDJ9f4xSCnDMrpOs7YBvXtZn2Vj4q0WW8f4Tzeklunc1VNs6gv
47X2ewEIe6vH+BVEs8lXTi8B8SoRm6u2r0R0Bjaa1kdEhqL+nWgzlt9L5Yb6xxKc
M9C7Qu2hcSvp6BI4GacjPllYzFcgLLLXMH9Mr5JiWW1tbc8ln6JcP74oVQkkptjn
3WAiG/wd8kBF7xLipHxn0icKXluCMvtW3tycmgI1+tQi8Bf9h+yrbfUvBuLChhYb
f0KbbhJWL60EtVAQ24nUgrwvodOmPTFSGafaCVB7DMshTWpMbVRx9OgyedSEyYqm
UXQOBAx3J1kCEmLTIzKWIZr+/HnyZ6T9Uxaokl/m79yIINpsq8GjRsRsS+Jz49ln
ZK1xiMckkJU7ECgdpnzoJ2x+G2CSCfPomXAvxtB246d4yYnYzhFX2yG8ry05rKo4
oo25APxdcUVrvLxUZ1uzEh6vTxWfnqi8P64wJEFaRgpGUG/bwJAJpgw8bCDO6pvg
ajSfEHbqqJOeK6Lj4zZQ7YaEfTw21J28FdRnw3OwK9lVBBZJJfsA+wjqXWyE6Y7m
JHYKBrtFsW2oTF1DnXeyMW7vrUFiCyz91dTFlu4k9HwVfFUEwl3TQTpRM9vL6CoW
y+jqJN6HD7Yh8jZsXE3xAmKaO40TuLIKfVg8FyLgteXOpzQXpqRE1gHyJcAHVoh8
uTT7rF+QHP73BymU9eg6y289mM8qeqQbO4IS6DDfrN+FJCQ9LEkC2xrtUrBmOv0s
u4Z2LG1AXP7XWPqba31kMAWKKLyPm5ceBaDQEt0OTCbBG9htCfQr6bBtIpC8r9ub
FFCx7H1fHTskif+Shn3Z4BeTeZ68ip/j27kOSUHSGlhQM83CU/ixU3QrGOzmxZmw
HlCXFy+dULSVc7B09wbtjOAB3ZS+8MNuoIcHbmr0EL4BoLEPMteCMzthRmCH6WFn
6SWTZ1cdzHjXy6MLla2YTokQJOeTu6oAe6GzMYQxjQ9JQNq5f6pvKBtELMnyR6cY
8Aw89HdHPrqi+MMQrPrtEn5FnIlfMKWInhvLvU6IrJVmL79XywCg2vUYuDQwAOqE
9Wn/gtcRcM4yNe1x4acVIJmhvm58vZQey3AO8Y1MYd/jDZTnPBt8VFLOfk6UOagh
nF9F1Ob4QtOcN7atXXlZ+s1to0l22BLx5cThBKRUUVeeiRh6IKKjrT6b4O/R2UpF
w7bb4545PLfciK4zwTHDdTgrnZF1ecDHt4vZUaP6J0a8861BnJVcXG0qeY4dBIio
dOpzWfAcMuFfZe975HrFiT0ZFBNfNeZJ9W6gtz3/j8LtE2StptDfHzKRcZOTjCJY
NuhRngBiUuqlM7bS8yhVBS6G6ehnt8njOhl28IZ0btU+1UTPHsHsQSesuWXpL+/5
vrE60Bc+Vdr635vg+wUgDJ1Cr0Cy+VgcRT4f9H1ujq+Kc0WHG+ro3tkENcur7PLQ
zt4a1vNvRzzAmVhtgdFEhXuVx2hvBjGdw9T46ivYQN1h4axOlFXD8pjgtKRYxKxc
Yh7q5F3qwRmDi+ntwf8VKbBeiL0nOzJBoCGvKc6UsNLPFjLkDIv1r5APpdXMvM6a
exLZxJ2M5H7XNVFgUI9qfb6Y3OPxXAWcdsVKIkclWNCbhN5AuveGSi5iZUYgmwWx
e0TIOGBaRvfY6l8WCrs/JD2sgvPWs8CUEPdPh7uq3qSktH/Z38xG4dwFoaxRZaBt
waZJaMvcj0XiS1K0/5j80jye1PkGio3o6domosS7NSk8E1Hx/Gfxv9FfvHMBJ1dg
WJZQXsYyNaL6oVhZbHPJzYfw4MjMafLKe/tdURfxT+zTynaR/vNcv9lMXADmh11m
+Wd9T60tfuIrmbPrw9jKpSq6gkJaMczm8B3+peYwWc5I5ab+RKNs/J1lZIA8HBAc
zGYrRIyEhtPQqXzjN8ivWodaddx29uDKXqg9sL7zUAH1dnhP6uV438fJe1eivSF6
DSgBSh+fLJe1+1zqbFaIYXoKp8bqUqjKqdnHtQ2/yvY9vPBiVZTM1zxDOC/9J/CH
L9yFA4oy1v96PMr0goY4hbs0chOTf7ykFhHMOZyNSqj4yCJVKn8nEIHW0CjeuxzO
ZLFFuva/+cTDaExHkLUAsykXwLzaauUnZOTEobgTERGCGK8YX5GklR34SOOne3tR
KTxP+AKPrwrpkw/y+b6JZ6AHTwcjCnkMkwi9ddplOKGpl87nqNbf2tKYQc01pmx1
M6usj0A2Yt9lE1jXYPzDaXSk/cF1H7sd5UNRdYrZNlG51GkwBvTmYsaf+rrO6+IW
oCJQeA1MOQJqD5nKv/D+1fe5QPE00c3lKq7cVVcocnC8nnEBZx7roSABQi2iQ6mz
KCSOjKmRq+GzCVMQCLdpqn+FvnH09JLCz4yTNcpIwbMVEu4+iHFRFQ7VtxYYSpUv
VIxNoc3dNE9EKweZu24tlHaf6zyJEDHIN4nad+VlD6cMbZ/U2hLiuu36Qsbv88A9
5Bc+2cjQuASBOh7d8exZyRgwsG+03ID9TjHcnUv1cPJYDYXS/UUO47QDaBZPzSxA
ohcW83hm9lhGYiY0TMNgv9LfziuU1fZp/DpgpKHSZoIeAmaq3iWSz7O3vEFu98yY
QxBLX558zYgMd1GxKqrUwUnyHda8PND8Ca3J4L3O158zRyaI/VWbs+Z1/a6acHpN
8k2V4BGXsUuE7Ew2JKF2tMk1Lr7TPlqTVx5CC1uFUbJgQjgMBE26GO6eDDReB8vF
KY4TXqi1RekS1nXxzdatsRc5wJQKkSCMwfx4FFywxl4cK+CIp/yZwKZZARGR5ZLJ
27xXXkduEqYzH+Tk1kiMWwMdrSA8a6ZzGUdcM6U2T+iwlZVHE88mIy3mw9BsuijA
aYPiOuXuciepm+FejcUQ4a9/5qGjZAwx48WppklYbAp1ll0fzozGfDrKObkKBHR1
b8ZuVB6hJ2MemxFMUwhM3eKWDP19WzRPmp0k0//O+3oSheAM83U7fl7QOqXePKGx
b16T94c9Cf5Pe4VXa5xDDLY7blxBxub43TpwrJwUvBriSCAvKWW2ERUJ6T+42izS
DlEDSRSAykhEVUYu2UUWPW9+JzVU52n6zaqq3au1c5v53Qo4EId6HJIaMJRRyUBd
8VYYMxfYvmASIagMLgn0e3uXzyVbGPLOSA1O5Ew6VSlK2Xlf8a/FBxQmz11G07nO
l9038BOLi5seiufG3nfYiJjv92F+cdQix0sA5VohVGIjHNFDJR1YwJbMLJGLJisA
/SX915ofR+ue9i/QYnb8AjwE0I3oaMKgAWahIgAItpcn/1vsIimW9fHmri8HX+NH
OWRJ0MbD1nImeYDIiuOrhzyhXJrj3d42TgvGRo1g038y7W/vLT7a6w5LddZ5RYKy
Pc5kZvsuxNXDWXNz0FCP/v721hApwFmsnRiua5atPmUt0jUQo1wlhStpKPs9AsYh
CqqWNBPxvZC+eTLpMyB318J8JxAVNAvDhrB8n4mmG+7ZTHyTp6gkjNrhiK88PcwW
jobCkxLLFF20aU0DaEgYcrqbS2rtFAwkoX3ppTBR7Nte5JOS1MJyKnJ+iyBwmPgd
Q/yNNsDtUugZBPoOYi+Avp8FakzwdxF0AtvGBV+Zm9dw4Onaxk8TFXSrzSF6tTtH
xelDlRlllcr6XzJpSPBjqkl2LGwPaaC1EwJVVE/MXgzwaNbtwZTGgFMRYaL3D/lg
qsDwttmyMb0s0Ul5RX/dHiZBogYYeWljW0eNFKjFFqijUotxGn0mwBishIPt0CSP
Q5MkppTqIkWMg9NkM8IF08EvOaMOluDb+/HZpOWQiS6wAh+069xIX3ecvoj4Y2pC
oa04SA6gBdQEP24AjHdrHFw18IKIeNgArdA6BB/eKQEbmStrokGdZI2yMiwva36i
h+5IEwHN/qycYkbccwVMJ+3TERdx0NVcb6GLdVdo3E/UWceM6fFpDYG2pKlwEfv/
YVlVkDTARfxO3x7Ko88WXo+zmeJqulSjKV4tglmdGyGIfK9ux8tTjr2651kUJz24
Wb7atHfE/EQ7dsxg2wx9LDTwfQe7nQ+MqdLJDROe0r0jxo8bS0y0dBV45iT6GJuD
WccIZsJKeNHi/KGlhU3Dv5KQgNd9GVbB9UU5UGiMWdfgGRq6sb8IoMtgNbtjC0Ev
l8qf70CJ9eYPnzS2OsilV2hHP9VeOqEPHrJUDe8klGVS2hG2GvYOrWxwlbXJaU4l
HuZxoxhpNfEKD2p/mWvC4bKc8JjyLEHAwUbPCP0yqowhlIjcfWdSrXhhmMbzRyww
3WAx07ODNi4j6aADoiy6qI2ETt4i/Zio/d05/9JvXO/orgZZybmdkUKJV2eA5R3T
E69DEPONCy3sXG4FJje83YQ7TliwmstYhyDQuRpnR597OVsSwo0+vtZ/x7MI+2f2
fx1r4gMxoxhjgoYI6Qv/7k7a8iW86jICz14OYB74KQhU1mvvkOpdNzn9e7Ovzhwz
jT4VGR5RQ5pZR/PF2JXuWXrNJ2jbE8y+xGEvnskpM4A6cTjcG/460tTNPdtuEbX9
9lChxjpli/XAyseTsOnqLzKlIAlwtyyTfJqR4Ri/TT014AyLUgOQbob7SEErAeKf
VtnuB1fNVllO8rxvyUgXU6s7HPBJvn0utF3X1S+6prPF2g0oYYknJardwVZYOmFD
ygapOJT7ollVFg1OI+JsJBuTgcxX7XXVIaoDOxE8KomEQ7F8+UmdecomwoRjnkKp
It4G714fyI1JAD0Es+t352y5aLkBKTgqN6dzvp9FeHRT2Wu/6YyyycyuW3LfdDqs
wede6sTF70lP3MJXSNlHu9Ry7PO18aea5mck20Vg8RhzDdk/kPh4X5Rit1ebFC+U
Le1QDxCt/nDWBY6aN9GGcj24eDIzjojAJqsl5DaD4S9KORqQ/3kOsQCD8DEWG6H3
wHdqrCo9V8cZmXmyXp+i5CKTVpBhD4MXCaGlPebcNix0cmhH2SFotpIhJHp8E8e6
QvJB4POfjmBPgjIJF7txLO/TLU+CIOPgKEP8wI7ujLJbs8QI9ZSm4YQFfISv5oXm
gFmUCEfn0nrb9wFtlOggpSSRzS2MyqR+f6mv/mqVQBYd87CB1cIUYqR9NK8Pwb65
rv0wKvJk3jbLiJow+U4JvNDxxGn1NDBDu0e2oHIuDkbKzXB2Ab1MGqH1hLu4wtEX
ioO5C/pDrdlfdFTpf2Z2AYA/m/jE7MrFPZQ4v+HF3ASfsG8k5vKjE/qlLflt7ajK
x2BBMxXyBSAWgD3eg+Z263QdAwyCTWugOQtq1IltNfDO7Fx46IF3jK+DtUx8FcgZ
6Dkx7YhiTIm2RJZ0Wy13R90pl8F3FN/McX5F/soLsefijqWixuSIEyO03HnUINxz
mVmBj4V3ap0RWQS8oZbWCgF2cLTPg5C0DyGvQYVKQjNRvVLTuHhRnBp8RJ12RpEP
VKjEtd8+rkbN9UNYl4AQ0ZBjVnmnvDgc9e60MVULpQJrx53UBB4hcwUwBtAsJ6zm
aGwmTiR7zVot1+Bkf80KwJR0GTh7YPP5+BXql6aE0MUfAt71dBj5/Zr0UxBWrw/d
hDC7mbsKdqlPdyzNvKoyMA2kEz1nxTHsJgGbs5ci2pRRPeq65E/ha6xgOUtxGuOG
zLu7Bqp4FqEbO13w48uXZ9iAcduQQijep/k3OJRSG/MSlc56Jq+MtUW0077njX96
E1vvp5jzrt+yggz0hE8cSKwq1TdEJxQfzCux5682GINS5a6i/luqnv/Qq7aAKkA0
IGgCoYB530KqeS0YYkLYW+0PFMAeKTI+KBNsvOW7qxY/l+/hdSaPzpfd1JphURoP
mN30YFiLHimxwHBf5Yy3YNUfbz0Y8yVKyxDsiB9adb5jq6QpdaCLB2qcyHcZR70b
ZZ+ZVFKgaGyF5Pn+8sxnla+Bi3xqOwlpcT5J3Ik2CnLXMnJzBuy9jfVhrtsvZsXO
R05vpCwAXwyi3fJQGTDcxCEIC+h5ORl5JY4EUlUkH7o9WA2mRjb0SYfdgSXTj5p6
3YheGN9UYv74wftbqC5RQ7U/jYBiVV3QI/XhVe1WntL4D73bs2Fh3kjs9+AGlSPQ
QqyeEVndK2HQQbw727FhujwhVJ1p/IbtnGGCAe2dqO5QXN4t7+mnH2vEOXnuv6fe
iau9+MxoPTtDYRuoz6dV597wa21qStzd6SJkLaZV2n1ZbXcfyHt+9Ro98QAiyPLM
QFjmsUonbs0j8FyjOci/PDy0VD5P/WtapiP3rOfsDMsHfFByOBSPGyLStXcqVQL0
sdZAvzeuelof9ZuZxITkFdlKfwid3nmJ6fgciEn8SzplyI+pT4tGTdkK46gCKp0N
DPQSwy34Hc14C1+YtyyItZizopwsTpVrikLNvR1bTH+5vKB/GjlQQXDAClnpLW67
DQBGMWYosXccBkCHNKaJGPuiQDTT+FGhEvhvCzj553Terpi2QQRHYOadcwjApQfu
qqkQdYkQyPCSUCuiPVGAES1MCqL6Xvbbvi/QfEeMYrj6E1SBEBaoZ5J/WAJAIelc
fTuwaO6A+HHt9nq8q4jNES/VmjdRPPddyNx4QAxIXw+6cYkRcvT506v4H00iIBIv
9N8OVSDYotU9p/I3+63e6eckla7buR5z93BXz8xH+uqwOuq3bmnpqlq04lggELhx
CFYGWOl1YgkMv4KWECCit4cldHbUSZDIKWY1yIDqBj1YT+HQN7pg4ZFzDcqoZKCo
IxGA0hjj8e+tQhKye7bL6YEXWz8tHXVyE51ZkYLV5oUl/TTFjUPiVYmo0JlVShbH
sQ2qzFDJ829T/NVQI8egLkuP5o//T2MpcnZa6PPoBZNMofQ1Gs/6ghHncrHbx1cB
MXjluH7ThTVFsl4QMq1mGNBAzCs+YYcqzwXTAs+ffJHrSu7AZCvTSTB97UJd7q+n
P1grW6zJdk4NwKruw/2cA2Fx+eEsG2e2By9jhHSzjB5qTb3ad3jf/O10F8PoGC+D
+KPkfoglvld9k3wqF6q/JDm8/Ur3R77a8Uob8kKrZJCyfvPrmMlE4WSDOB7MZpv7
fQv/CbUZ+wCD/JXxZ7pjcnf2xBG0DHfSXyrZdbq6m1vfWCuczCiArdPIryN448z3
nRrCKbOPdQVTfxryPgplGaQ65/ODh6IccQ6QZq4t0MhkkX/5lPNesiFlao123hnC
EnRe0HSm+KKgC50HXzjJT6iFXr3KocVIkcN7bXgtLPyA2DL2LlV32PRUq2W8KGBg
HpWTIF5Jr7mL36k/X8Gs/oprvVev//ZWL4tI2XhnY35W8vjG3rOfJq++JnmrpjyN
q1KQw+Ic2NRQG7JgOvRAN8fep6LnpyK8vX6PhfmuVkUErSVDL2bZ2x9KI7SJ5HmH
WNT0AbUB6BIHhau88ajD0JxJYIlktF2lYeN0dp4AfHU6tIuoYdubbUGj2IkZ5gvZ
GzntLySbM4tSA3VhKcz2tbbZEEQNuR+55jnSjHVDk2tleJFATlOuiPSsQ8x8pOAn
Lm1J/8NQ5tjToeqHKs28vgOutf+iH2bkFuhNiq3+KWawvaEOax3MJ192Kc7GhiDA
gpXWFmRAT+/+H7yf2XN4CRXdYBe90C8kqe0dOpXX4/d/T5VTAdBfH+iQu6+pQF3w
N8jBAiN/JB6bc272CAy9nNFHFHEQmL0fB5VtLs4iPcM8N4rYLYdpdThRTQrjg6m6
Ev5R27SN3hlz3lECmdKmzPDwxFq/OgDjOY1tb67ddkIk8nZHoUDvyiO+9L4hWtD7
eEpVnc3BsyPKlE2HtJJBf0U1ubxZ6w3oEVVvrdy6wYzMWlkqnuJpDOvWpoVKo1sl
+eTsul4zu9iRiqN09jK6KJtUVl6JjgBSebEnqoc0oY4kt0rK5eDJfSpmY05+Ogrl
1Ad8fHX1725gjvHGJvTBrrCCiQiIyHh6t+Ej0IFONfUZtdTqGaQvJhtZ0wKbTWJz
al9kMh2CK1aeYOKAXLuUh1qWOPDaM1ZJZqAnk5+DrrczcPySIUDb8P+iJoKOknpK
gj1qz9qGoRpJ+j6A1VzdQ2V/VsDCZiPMbmK7nHYnnRSiMISKVp+XqhGo5ec36Pse
ic/ats9aBlkzYdReWIullTIZQwmD/V7dNcnOCZpfyZJJJOxSR+0qbMb8TgWCyP5y
hFTa2QnmjRLckPLl+PkQT2DikUWuFfahhGIIRkSvHYHzjyb4117OYsfMI2dwCZ91
XVP3wIWMJ6ln3vdicoquwg5zTab6JxnaUV/vWTVwmRuspveyQptL78NVX5fxVY1Z
bnwNQVLPKtMQVX3vqVMDhlZZMVCzW0RDT5CmxBK5pA0Ft2aUh+rTeMZevATKIdJG
badBElYOmrOTUUgu2hqmv5JmUNeCN9h0anLPk62HTPHUc5JNWc8YX+QGUdOXL9Sl
Ipj/V6tdgSiV9IeLOI5LhkJD79wKNv9kb9I5u2yjca5wIAZKGNDk+WaZToCuE4p0
hEyJ50EwKXQABwzB7uVuhOKv/x29P1t3Ot6Kh7icb9g4lR58Kql/GEllQ8i66GsT
PQ/cLDEC+Xgdff/hYMBrAN+YAePifSRModnwVT2yCPYpWIvRvn2moO8XkPtRD2JD
VyeKXrWSwNiaw4DiEbtNJdxZv5gpbj85UxXlus6nSNGOrcmzsA4OEiNBGHRoT0TQ
zMacDtxl6DGspyVnzFVlgHUlzBAV/FWiVDzhRUEf8h0Z/AscPpR2KXyp3AwoP7XR
3SV7ZNaWhTa8vqtgG9Ns5d/ve2ja1OHFNio3dxNmjR7O/UgHxUMoUjvqBgSJbrqg
UWfDlVqiAbsV7iR8ooa/FUrnEpOkz8ABQUYj4Ow4wpudUmn9ZnQUMH4z+nVo7qZH
OjqmoAh7QQoqgodmYsTGf+p6ao6HyoE6mPHP7zwAxWqavz/m/9F/QQEldZBmIsvJ
3+RdMtbBa0N/1m7y+RdP6kUYF9mYgGRdJ6vtV0Ct25wWRgLdaqiN1D0zLPK7oTAn
LWPWjO3PewM65jYLVwHjK2rPNxBVwJc2wlDnBX3ihcWm/pafe8aWy/EEET4hRqUX
HUbQTH5DTTV15cdUgVkt0v6760pgdXbYztDMwhc/WojoSrW/fG0Q1cUCBV5DefBg
HcMBYud+WUpfNwPfjpmc/2OWoKTVradoPvZM3aG3Kiigg2nm1/TbedvtTdNRpuUf
Ea5OW+6yKSMoD6aKUXx3kRzsG2b5Az4nVp1swXBtxspI0bqVKlerzhcft5C6Bpap
pM0gr5Qu8uZy1bft/BfXe5gX6llnUsyFpApR6akHolKMDlYff1Ks6CTLU9jl5yw1
xjgDIls2uxUHbZGNckhzOLL267QV0R4HUYU29XMYqhx9X0TFfQrMd6OpNxRjh88n
D3qGuTFxDnGKoRukaSozTHqKOQ0lXdrmPxUpDqib0RLFMHdBHrG+7PoXbTzUhSHI
u64h0dtGxC/7ji1Am6aNwm4JhjU1rIALVXIFkZJ5tyGke0+R8dUb9OqkdNdE6ZUY
i9ysgeu2NTZ2WBemxY44bsY6fighzWxfMiE5AtpYZloayr8DkZGI5ek65XWDhUCV
iVUvr5bcZF3aMTaosqLbNWX8tJz4FBNeUi4rxNxDageXpUR/HGPvwvONEl3NXMYm
Rqoh3TyQxfjB1+0OjyDpSCLYei3Rrx3BK3CBjj7X1slpa+UFc//Fbz2cuGMSfg/2
W3uNE6yHLMLBZ8/y46qRe3Y8A/erT4jEFZhK+BFjpeINy8jA8ep1rUYzfH6Lusa8
+Q2iwAfTs6WjN/7TNOYlS4nWYazTV2i69N8vkiN6PtJNDf2yBMsyIQsxebUZKzHC
Ds2/L4HP6g0Q0rQcEQ6aR8mvMM0ujZfutVRfzxxUg4uVUnbZ50NKcPjW4is8aDke
ApvKcxWlLW/b6G9LE9Le5aFvI6DArhTprdIzIYXOI01jUGoxXr2L8DEcYuURTfuH
EZih6Kdh72hsjkwXN281A5kWdrZ3i1isrV3SdoK1sne3QCBvHVzZyU72ZPGd0UZZ
RoyUHcq93KQ0WJO8ezY7C9Y8mNs+V82y1tL8rEWK21BGHJNeLSy0sLTZSrApFv8M
5QVPs8ItxrFaVCcwFIzFa4AlJqb4RacrJDSz317dLEJa1OvXiPXuSfu1CsaPPltb
KR1y27/V8Nl4FUFX1I3UCZv2TmCdGmGa7txag7HFuFROmRvlDSxJ+cUjyGQzuXvG
cAYsz2fdriwCiBpDbWscdL/eqq0sEUNac37MEMD9hn03TdtSShFvPD2osctHoGg4
FEXy6NReynQtCN89PmdytPon7ds9QZ+ji64WyCDKaZrIfc9UJNgtkIBkWbpD8BI/
6gV5VJh84nH1TjKrlq1U9wpSHN9HV03mFcS+SoMAJyA40s3jWsrVrQnYePcjIgIu
ohcQFoWMk+4lHOYmShZ5faQo60eOVskDml0f+CpVBD7xdISRdfcljmlubg0vZP1A
TT4fiZ9ut5Y/bBFxdYczX19z1UwXQ/ER/M69N/ysH4EpAgmVcENj0gdTnQ2XEM9v
pT7QNlkRRhAwVME8sLoNa/rHyWZo1Qhik+I6xZKF9DQFwohC8xwho71V1O0tuHKo
d9xqc23WqJgiuwkegPOe86i4gqJYBIwELJGCGs+Z7QZ1E4y2pyrEZEKk9wwXizmJ
miiCUx9HFrHFaQp1FAUzfP5ATN0bVy99MNyllNEHpj39e0eV73q09hM+JcJlLxsC
WkuBChp3A/jUsSVJQCO9DGH6iWwTUgaHw4w5Pq6ciN0g8CMjqgZos7aeA4E/3iuB
NDQ3QMjmTIYimsN2q7lbVWJ9rHXpTVaR6W/nFzJn4uSIJwqVjq00ysV7+RPj6hCL
HUUfhGExKrG1VLRfQBbyo2kwW+1hzRPvRSPPaDLxHX+3ErgIKwPxFEvDKyT5xTg2
xH/+jkaDNGuOh3fAuVFlqwHATq4gA5rLlCCW9fpRVkSQwMXXt6SnTblua4Ax0q5R
FuRYy9PjBC78FjK1ddzqXsjM5hmhqWiSaDCToENd4o1vnIzweRSqus98HCc9z9kw
FG2Xwl2iYMe8Jf7R4L/VbvD3qWa3D9LD1y+/5S427HLb+yPZuRyOFvP4Ya0VV5ZP
b/RY9I+kJOdWC/OmnQXwo1A0/OogLJVD9C57tzIy4vk6eFJKBbLvbmBQObXgQ7Lr
QvnUQXwCuHxFC4d/g+A5bn4kxb8S3ncREMeIjsnOmwjY0LV/9ZGKP15sdofG5bE7
hf2R0r7oRUmoTneWFNnTIZgnfocBJBf3Fj6CdsWuU15U5rYpDvUdeYYdW9JjmNra
oMWZikgBOc8giifvGReG4t/gvu28fRNCs6r1llpUE7044Reo1ccnzzYebbxvcI8q
tMJu/L9i4UdC2Q/TfhImSfJseAy0VULYbIX9qsmU5187jFH8SM2r8p3iAFW3//+D
XJSSS9sxwVVXrJvSUTFZekrUremFO72WPHpJIErGcWpdJVf3Vs7pMTC4fi+/4gmG
v/xieu9I40WSQGUNdtN9moLV0kJLKO+T1OjpvJhMEnSLMk54f0WUYO+ZE9a50ZPb
/77UdyiK5F0jacVi1CsaHDM6dnmUs2LuGgcZZPOSRzYuCHWd2xa97QgvxFTtCdrO
dc+FAg99GV4CNGsuVQq8Fih5Y26ppO2leR/JGKmXpooU5pzKbVUiXqlqlPnT1Eku
+z7PedaBuoV4+uOPWnEZW09wtxP/1xOXEL8rTtvljpK2g4ZX9s15ZjWClUYGUTkB
+ylCwTgchvA8Uv6A+7scqvnV55EVVuobn7pLmBBnHsyn3LFrA6lJDtVT2mG5pQr/
hi6K/RhTpq68DgueneUfjNJBzfALoYQXjHVmh+4CKVpflr8bK4vBT0X0Jnk9l8MZ
4Fl+ZWjU+ir8Lm31tNGPQRaOEU4ooqaHAyLbgc2lxoGPwRGvMLJpw3M9CADUfmeY
k5RjXPvsi+7qHlTfjuywZtqVtDs3nvSNcJQT4qt7zvk+rv5PpbN0QKz7m0Z9Ew6Q
y4edw6p0cwXFhOiFlPgu2+h5xQ8ct84UMRlhng0xHoc+H7HZzuV7nCXkLBb5Et1n
cBoraMd1hBCBLt+NONieVKnQF711gnlJ3kx6gTUyvpXD9yot2uklx6yB8hsJgB2O
/zrTAzGZby+NF1BNMxvXglN/PdrNmkjR2iZt4FL8V01m0YaJ07Hb6aSIz2zs51Z5
4haUWomX5rT6nH2GnODGxIpK6LJ0SiTNewVn1YNudQ8tmWIyxYD0Y8kopO81bjhx
5t4oQdRe4x5blcjvS/DacIFVq/cHEk1Ym1ZGcrCmyl9JCWEpfG1qfFGSRDmltqP7
0EORqasyyWdT39HM1qwSAztkoQZnAWK1yViqJtUt4755iUdOLSXJfpcYfDbKl6dc
HFJaJ+vzyx/f5NgGW1BiSW2E71kvwRpUsoJMC4UESKxA73VM1dDV9apdK16dLJDb
rDPoujfx1tE0MHdm5Hc0Bt/LrOX+aTWA08EZiWnaXTt4Zg9dclNTIWBn8/CQm6iL
DjT0nA48jWPrdfostR6jgVuWnCr+hd+hXUlckQD5+ta0Bqy28hVQ1vwcBBP+xaGe
jugw5Rd/9lRya5N59KKQTOuEXPxee2lOOWZZdSqnuAnCdYb6iYmKo+LzisA0YJrw
v6/1LslW/cViPUxvgeHeCN9oZTl+l3jAtMbuwLAeQlkALq+6qTdJ9MUWXyxLKCzG
fUzI1lCoNMtwyyUz+zY/LLmHaKIzz630j2SR3obKjnvXPVe5E+3in7ClThVgcfTd
z/+NsVP9K8MGTfNDqwXajFMLDwtiCC2/Ap7uDv0v4/iZv7YI7zzJN6eBhLGDtOti
qh1WEHpXypl1NC7r8S+0VtvDJhUA8lgI9OoLv0CofgGCO3r6eG+Nn1DZctssi7Hd
qV4hRgTvWBrHxvi6peElnqvUsy5yj0GxHg1yifgv0jnFNPpjNQ44AuuHKAliMvBM
M9P2jsr5PAoIHQJdfAM29cxbkTLCQHZxSW6w07CDy9tpfPtLe9Ee5imBIGmsWcLh
vF+nJVd/AYuxaCMTIi/LfLkxN8rUO/BDU/iKKTkeyn4jeR4YwoZNDoIHCmz7ZNQZ
m229FweazQJfUWl0u4pr6zuqrX7lElubfNNQ11VRbtc0sNeGKMJ6xhtuG46qmxCp
Mdm0s4BGCA6+Ls56Qv7OWO4YCoscM2Lq5kpds31j2MRPui/HU/Z7ROjipr0qCCuK
PjWD/86ythDDQOJh+XoIxWMB5vHnNokc9UddSJAiUOHpVdoU8+OSUPn0lMJxVzZ3
mv0Xm2kRtYInFdzv6WW+FNGdbta6I+NTXjXS7JWdjoif/DOmUvN5yBMXP0x7AkdL
9ZXZzI/PYCjXTC8/CxrHCf6O51Zl/9/nBtGVim0rinBsnnmIvpeL7YDFJahwzdcv
RGjsib6Okzax2q//9zBG6+0BzWcvUAYAS14ZYjGGQYqeEjcpfqBhW23FpL1uPNpu
XYB8Lb6mDoi4Au2WNawXLFC+uiMKDAQEsb0HJ/G22wih6uRzGYFQcnkf2D0xM1wu
58xnhHu/Drc1w1ODULYbXHCdxCdT9lbHwIz7aDh7tlqn6YVKjgd+FkEVAiULMhIn
7kC+J8zjCkCpNWehQqN3AfThgZkTVmYuuef2Jc/HajSorC/kcyHcaW7QMBtrSxMH
n2+k/kfytNI31rI1OUMlzO2J9GBkv0WOSictxlClodUenzf77hnapOEgpGhhl70K
ITc5dweKAhmTdtqvPNljzX50K+qGOCbI6pu0wr9N0JyOhlZ23Z2ivm4IA2fpqm4s
rFqFtZziA6lyI6B1IXN1D4Tmp5k+ZS1spml81N6OOGZ4ccZiwetdrSA8Kmh02wc4
9aIeZmv3ixnLWw+TtNVK8TAH+SU2IbLvq0AJu5a5QlYOiRzAEzeR8MgjOUPgnrqY
19dwqqEn4Fln+WCGTdC/W7ig80aykzaijo9GOBz1j/stY4a4F26Av1qoVZNe7QBS
nKPT3cqte1xuCDAvX0m3LVFmPENQ9rNOLkTfn4zlchQI0fwaBAFykSlcjR/ro1O+
u/B5hlvzq6xppCwxg5aGhq3IpMMTuDjJSDScm0BdlnBFassSm0SWDUmW+ApSFdjE
uoEdIvcuAuEdmUrHrR7JZszYeBkfJnb5P94OCKRBX23bwlh5YlOd28M9Bo1EnkVA
BbLKgahR6NRCsixffINNH896wGq8KBltKKDBIm2BaoojLAcVcp4GnevizJlahyiG
2oA+rnuHzZ1WlJAYN5ih8RoVVv1ZrNPC4TtW8CWQJC8khx/KE3WdIruIzb3/yS5E
QwXn0yAHtLj13iv/zYJUhiYRlNkr4tTVUZQsWtGMMjaLpckhNlHCGlCcchyT2nML
+RETbbKwl1Y8e6a1Cts8MjQYlL3boFq8RRmSQVRvSw7sia/VW6KBMSvO8vpAs77b
0ZDMHYL/Ps/Z7wpVAyES6duisFtcgafG2XL2O63A6Wbz/shgITHuyz+aNtgsvJVn
iV7IYp+tQcvVkTTBIiJAbG9IzW04DC5QaOOWHOSGhD/jEPBYDO8ZGc7ICC2wRsqR
YAddx3Z8+DNDavPKCkyzvKp6A9SRStkv+lELyO7wsq2ICGKjsPmCFgimWPuIwBij
ujRKxLhF+cwRxU4BtWq57y8revSfK1F/qUZOZoP3FSM+6+9mZGhqpcfKXAbu43gX
qC5MpDAhGsXBRpE/Gd+AUdAQ2lVo0Zqx1dvKfabhPwv9sxPXZdESYVMO/50l4kGn
czTGFEInuxBtSzjp/Y3Iy3gnUBe5MvS7Fo8q/ZjVbovOzIZlIQCDBgujq7qNykKn
k/L0DZGiSHVltAfkA7hhLNniD5pepXbSSjRaDUxifVJ0o9gMZGKD7NK1gW+CFSC2
2I0V/iOB9/MMyLsFZmk7GXYNh5m9ItiEtQ4q8iz1n3uPNg8L+c8ocly/lD07+W3c
DJm8ozGFXIUFe53TmLdi+IpNIRPZwWNEuWjyJmYp3F1KdDyKx+I5gkqaj8dh5qc3
9x5WWdiZEL4xQPx9YjRrzrrhd5VZsdIXUwXtNLROWDCZ1LCD5h8Q0zUdKG4gwZ+W
Lpj9hEj+kCV6SLoGDQxFcxCLdaOQiT7m3xasWHHgK3NNwS/f67d7f1etDQs9ogEg
oXm3EnIUSga3sb2h7odSQJbT9J0J2JjBnUR85mdwJp+h+szWbHzGHY1OFRNXzZef
Eqf6F1v2ZdAqcUxEAm+cssSD0SmK4oKlVC+N4zce0k65eCOxrjSloNX1/Q2jVo1H
HUOq7NB8IryFO6KRnN0Mfk5p72pHw5tdkC3uVOOl3eMdYd2HajcJJX0Wq2EFPDbZ
CkGrLsl9iT8pYVJFS6J9WTVnKfX2BLre2ql4aqTRp2o53nw+2ajUZcZD5c0L+BXJ
b1XUiCu/Pl238/O+lg33yohnD37+iZ65ut7YFSG0OsU4wuDvMiKPLpbmXTu0DK/H
tT49jqeZYDM2W1ZJwMsn62b1QL4geEA5CjSh9mTOibtH/QsS+zanmiehpnMSXhrJ
NyaLal8fmCXWbh79inHJPz2wBmrhxTQvFLTgZJnUdSz7xR/6127/Vd47jpFX/TE7
3uNPhSBo6vqkANlS5bQCd0BsuKer7JTVMs2UZIg4PocOtuLFUKOezxIIU0Hnu2Fw
JdHFiZhZkTbaDRL+fT0mncPaDLJteARSQs+tm/G0GmyOzD7QTjTMrw1b2Aa8yaP/
FknW1+YavI4n8QamY5ldJqCwnfJM8LJre/f0LVWDyZHzAA8PVzfI4fLbT/H/R7lK
bF4w0OYEPDFif9+cylvj2EI6QVBC9ARNILpvFxtEW9bRc7d3cnqdtX/PwF392axv
ZC8puuFJIpHp55S5USRrd3oy7K/Y0NHf77WrvOe+FDptQvfpLKAgZ8UpA0dzha3y
G8PE+vcQqAdq9ZlAydby3tBqmUzu59oM0cS73g8dboBYD7BC4DHVKD2WEwHOGhX8
TPG2neQw6IjUvjyW0HUm0Ijr20bSwaG3ewgS4fT4uDn25jfOY5WJTO5D4fV5zKHA
KrGYboNGUVeTtw8nnPtsIEwaK5RDsJgm6XgLp/pbyjz2dxesXTbR3UgGEeWk5rH9
YohPzbEQhyuIrV7VRtnYWLJMyOTfUnJmhP8f6OU22mA1LZtOn0MKpTOpO2h+3pbe
2D3LD2Ijmarkn6jKcICERu9DwNCyJZCrubtuLdtpdPq1v1EQ0rLabKyJEONNJuTm
16saOtDdvc1JnM1axtTZO6i2DyMQdGwIfbzF737WH2jjZzbBGzPqsmUpsl5fAg2c
SnkJbE+5DMuU082Jqs2HA5tiv3txy88vNzjhTNoZ7XLrtGs5Sqfkcp+7e/WIOs3E
fS0tMKYElk1iRmG8cXqHESRYu+tpgbr+CKiObJng5eEwP9adApAKAwOxGoJ8dDhR
5a1oy1LpkhKD6+cP1sN1eUIRgTkiNE19npd8YikYHSzz3FfrDzmD8+uaQYbzqLb8
q73IVgrDwWGWFYkQwi+WMsKbE8k9R4FxoCwpab8z8HGhQD8rTRxP/CK+2myvDcXC
8Av4YJbrNVUf0x8seneCOKmbkWe+DntdPo9m2fQNWwyUbu3YXpbnLIgv8AQSCJUh
dmdDD7HwAem9HH20rMId95JXmBOnuFgr4pXm2rUTFC4DfeBujZuy1HNMWQpjdPHV
MsdRt0j2qE1Ie2JIx+YqC/jtfyMkaa28RFNA+hxeSvEvTfosxKNIVcGM94c50r0T
upkJvmshM7AJ0Uev1WlFaa/qz6Wb72ZrqhFi57/ifx607r5gCuy6EA4tRPcAomxL
h44HNjU3+z/IkGNvnN5lKmzmoiKbFUqcsd+zWQqJuDnS2egQg2oG1+q4CgWZh3gn
9meFTClkyuRZVnnu1NgYb2jQTfIafGFPsi/bP6sF6I4CD4uPlUlfEaMmVA7pgRtx
vbkjP6lrrNAcj4EfZlNCpASOOKpG47TET7HSHLUuulKhV6aycBUtqY352dA45kXq
4yVet8k2bbuwb4wjP0fsd69y2+EKuRDyBY7s0pVb83WM65sTTssFohy/Wei9AJWQ
6iJ5aBWtj+dwA31skOAA1jU+khNmkZXS7UtysNIrTiFjcAekmp2SHgsGwvn8TwD1
BrF0YFChxhxH814izxAK12iY14yK//rTQdCyZE25+qa1ITb/oMdn2K4cMpKTsPlr
MfBYRDS+JDizcvIuGrYo6TdeNRgsIAfsyQq+KUdVydSy+mZGXuCOTYx/F2dH7DHo
Lt3Nd+uTjTLGquSUv68PCT7hVd1hzO3TguyL+JwRy9DOAEivhXL396/o+lAZMM3w
2i+br2QMbTw2D6WbA1Xl5hL05PetTU6ePWwMIaTaa+ntFY+jJE0QgVdDluC5PAmS
UzLLENoWWiOGIspG2kKtxwVtqvSgiviPZQutmo/oLa8NbFW1yPhhgqdyt02VWTO6
lWLkeiOueGreFMnxYvUNLSaZGGbRCGDejVMuj0hK9UA/nRNMtXnlMhUBGG4R0aZH
gOTk52ukDf8MU1NUUyUAKUQuyoYjy+5OWGJJKjhqJ4dNmB2Htg5X8SenH5EmJ0zm
depgbTX7G4JMeo01STe4vaan1ZnysjcG2j/4e/iAdqF2YKg1ZwzePCgnpzgxVgwD
fKUE87xWyBHrqP+dJwLwaOSPsgssPXibEGXkdP5+lX2qOrnF3Tk8g9CzRXOs9Zo6
ZA89h8a5MjepfENojJZuas+C6TE68o/86khGiLIT7DdzqV/mVtne2Rgepp/zMrdi
cIXI+CPJMhWZIuurPFj9MBLv5sKj2wT36nT2AXwBwm5p3S32xj24SskUOlHqI9gx
HH2e7bI0gd3D6ZJ7+4fEww2XU7ldlBCG37roXQTDLQuC6Tzh7gUqzx5JVHm62DpQ
2NPTJjIAPkV39Wk6h1jcbvS2BC5PpPMVi2Cz66ZQyCOd+DlqZ3HGuSFJ5EzH1b9H
v7oYxzV6uVUEZmzLngEalXXrYJz76zAz43eKxCyh29ynRf+7PhiFWeCW5UrXnMdP
FOaObeGjRVNhJihvumUy19K+DRlp5FY8/SjjZNazGyuNRd0MQS4cL+JrT3o/i4cL
WTHhIK4fGlO3KOi/DSAdlo0uNxNmU3kIsNkuZUBvP7eY9ol8Hcd5nVRR9i9Is5Na
IkRLpShgHCyz26+GgNlDQ10uIACX+I0GRpthLvky7HgLU+eH15XcWifShdpcQPdK
322OwAjzb3ZiOgeGv+8Y41SEjAdsux1ak/KvQi2ikuMD48/7fei+JI3sqGodKBpD
3iBVyQ2QMLnh4STjAsPIFqTyeZz7bwUGtsC3xFQ2DdAWh4sllQNoIKGb6gpK5dX0
yW7UXstfAezvW4vr5gTq/dqqIy1mKEa/Jem+bskhBEeC5d2k1pVsJEDsIwV+NFdY
QNiUrbsr8HhSvF5uHkIkY9dMwT78k0C8FjhjXDVX5zOdh/QCbjYVIKKpdRdCqazj
WA9y8KqesrPhgQXDoj5N8hwdEyqnZWx2JAfMoG8i5/2qSo6TZ2gpPKg1J7/rMnHb
iFubSatBg2kRknNLHs5R/f9gO/ujPcU4dKe2SLJzjXTG4ZkjWH7kv1FsPMvsP1i0
FmrsPyEQ/frtF955X4XO5ReMfAbFU7Iiv5O+bIAM6UNXpuUxdaLUjSBe316Lau1b
kTftAgpOxwJM4BYBT2xnUDxYchhZpw/tNG3dqUQy3+M0uMSnr6NqINqvX6wfpNkg
XWpXj5TnGoiQ+YIV9nsLZU/egqK8/sey/gfCNgwMhjhJfrIemYqy7fwXHpEBBDoo
G0uNGj78oTBscMK2UgXt7s88LEZ2Nyxc+LOADIZdnJsYsdbkjzZzG97F/33jv799
tVDAJi7hfJ1cZjwUozNhqS4BbUgTBovoTTJPvlE+M0lAN4BfvULnG8bHVOmIQM7j
IfOdgsZdVfuDVRa+Rj+CLilY0tpkWg7VvASWFsp05/MCxf4lJnQB0RQb8Sn7NFTj
nvap3C6AZNRBfGurxSgw/7KdEtrIxbHXNAsfwR1Xo7Z1ABVXXVI6Ti7loGd9ouRr
etmvh6jko9n91IAqxnCHoiYzRiT8aod87BgjUI2AcgExDkeRV2JzsjEDsNWnSiZA
ARsuYmjsS2iFcjRII9DMECzLN0+hYYGQwiavdusxirVEJHy+ZSoZZbq7WnaP86qY
EgGjLulZPKKMsYFGj08i1tW7em2g9CvLwyIVON1qrCQFpquSHFuSLikiDf8maSUZ
vFIlVY8UL3A0eLQuVgs9SjspwJb/2CF3TpaY4gZFWPspvOMD2rakUqxcgyFzyKlS
/JC5Dv/wfsMI/omIz5eHFTV9sn/FWIJxD7RNxLtpFBIcRhJu3vJiYWopAxo6EsdL
l3HcITsAPfyf+Ny7yzbHZsqK61Ktb7oUX1quR064nKQAjYbVzcQCppISzaLl8Xpz
01Mhk2xtROEuxFKo4OY60MFnGSUBw0k76DzDeadenuQHyuhY++MoYoWGjVcCtJUS
a230aTJNmxZqHobiT+A0bpr2qXaBJyF2oeHYSB0ZVwCKo1ZlatYhnrkYcfiZkAkE
8abJ1K4x8SvQ51574hwtFVHrLjP+k2zq0tGZvDM/my0dnS9fL+0auYvcMfI4AehZ
6kzFYrlOb1VL3FahzkZAYrEp6DLZkZWSO6JiZi7LKQ5Bh+kEVceoKL6mfSMTzq5O
RwDcbf+2aXmHNrMB0jhx72vS5x9ru04HkxVUF2llFYZKmh2gcfwSrB1utVmBpWeF
PzoqSpOvw2KlmNTbEMa1nrPEY6SEqeLrop25oEIL32exakTOMLC6ZqsQv/hksUMh
r5MZU3WWYqqSW09mxFq2dI35+ABVFigv5owV69qU5pBjkFU++c/zciwRShulAsTT
irfqt93PSwbskzNkjvT8hHt6qhQ3Km3fv5q9deBdsyuaF4KS2XIFtERYcj1MzbYf
v/io+N53a7GYYC6v+B5SvqQf0ArN4QRD8diwr8DqqphcbpLqrpR03oT/b1RTOfp6
gSKV6Pvwkf6XYhv6oqnUDaXkF8ZD3gh1j1nhlIn3s8Np+8j5zvdHRypQzrYjrkCS
gnF1m6rX/iQbUB0TK7eS/8EngkRNrWfsMdB4sWs7Mjh2C/y5mNFuLD0CyCE9KJbZ
WIqVhs1GWwlTVefGUhpnWS0z+WEjCoXn4AF5j85dyMzwd6t67DasrQxh85SdKGjM
vk3++QEBbmzzL+R9L3fZa9NxKOiN/L9GcbkZ5/QR3NA8gKcZORJWtbnyXdIU5301
YUztyc+4eP60wPJthw4hiwDWJrKOEAZS1dTsd99i+kII4g/3MfDIip1h2DKVHofe
rkY5xl7HhnPWUhatfSgbHJFa5PBNUbMABO7YDOZoAr9ESa4QDaJnUC7k497zbRFf
MyhlhekSJ8jFwAf/AU/v16/9bU++pbpE9TtXHnkhKqdwbD+h2QgSSjbb4yFfISbr
JEfNecDx552leqo9hLYAN3gkvfglmfuJnvXKTI9i10QZtDZ3DLaJcqCXNg8IALdZ
afshG9G9XWAZ5IIBASFK40gMgDq3cbn+5IEck7Sm7DNbaGMWwApXDbqqrXisBwY1
D/WbGD6IipE96XJVpfXqENdHygJCWqilLceFIWdTvtcdoSnX/nWaWgAg9a4tKX2L
pVJO5xrGNZ012mSExpNY356yF4y2uLdyzlDc/W436EelUrRrlZtV1+nLJJfjeOso
lJ0eogrTbs/TbvH0F8bbQofccCYlBELxZrTzawDOGK6Xy1ojBoHHE++0SNMMHAQE
Q1GwvqLWt9wgPdcDpJWUgKQGdKBTWdaiuQR7GNWl0ugDkwDyZ9zDdZ63Ex3IAz01
Yq54NyakZff7f2le9lgtjh35lFx+lfyAQEmLHg6w0hNs/jwaoqdtSdjD+0Uf5uJ2
lHgyiPMuVabRInbNjU0usLlRkoUiKLP8m3ECF21swChI/YkIaxqrkO3xBd3M3wlm
ckCo+KetzY+A8MM6RF4jD96oF2GHPcrgnEqfUlYC1M4LgPZRmKjTMV4hP5NKkgzH
1dcwhr+05aR6CiIVH7VbD9MXwrB49adWQGLjtz7dx+gjgCit0hsieIfoxPdLbMwN
ulK/PSchIeyhiOJr4VqOqDjlIZBzbZUfk+Dt7w5Byrp7yZzQZfpdIxlX0qcxvgqE
+ntMMPQWchVA1sXSTpPchN9eOFsW5zwabvNOPT5OdRWy+GGyztHu/epvzi89FCtD
2KIhaH4qBpTG5kMvXPG7flDlSoOhrbKDFAaV6FWfPb7NMqYLa4+C1XQN53edI1xV
KkCM71/BKXXI9wWLY3NyOGy8pa9EIEqMSuSB2NS3FC4IsdaLfOeuduLlTJiEyRGW
JBIOlggkGIXG6wsydCn/n31HHF05KCnOVitYEAVro+haPYV/6lrOjBfDtbCC8ckx
Lc/QXF4+tPiOpV74KLNd9jdx1Ssmp46gPYpwSzq4iNDMbQt5AQrrzil27sOPBorm
BGFMeVadDRivqVqghJHeoXYlMKNQO4SR2+YdUwVS6NaIBj4u8quhoYtTDFWTcRvb
dWTRB80jMz71zc6mjvQZ+zr9cTmWeHZ2tACayEiU+fH9+BcA4tJ5cDusm2uaLUwK
2tzCPKFhVpjU+t/fOWkTT1ZAi7T2jf8D15yx2cktDatrli5AtSCQBtZqd/kI3nlq
KaimnmUk9kKNCHlcsQVmq1HeiTze9A1hUxt8Y2PXXVPR4Lw0x/ij13RY+meMmWMS
PE62AzMiixEiFMcZCuNWEyIHb/qRGIPeQle6KXw+vzETMNo5nk7lO9pwV2QSwz+V
7hRc8rjdtfZzWQZvP7Bcn1S/DupTkxOuHgA9ekN7iS+aNkoprZEtRRhowXKvqVIg
tRAsyugRtMoRsOl2ayQfSbDv8X7A1/nJJ6SUpssE/6+CmYlw9qDldFOGbSWcOGTy
T08ERZ54BnDSGMm47E0vo/BX+PCaLeI6b61aeL61Me5hzh3LAUw58ZX/USd/jhU6
ql3gRo3trHEeripjNIYuA8rszwxk2nvOHNAQ/lGhAbZtfmHAHRniJm0DBZvw1QAr
4oK21qwo1cByAo/Gx1w3uL13rYb2xhTio29XIIEYi6Aij6khPWENP/EBgXGgfrHl
h1M+SrIH2g6NkhK9pADeifqeT0vDjVUNic5kJ5XBeaUV4IPdKIYL5YNcdpOfPNdP
U40cqp6UBtarRBfLF0aEZ4eyQbrKZCtTSzgeHZdXChFgDmZluTfKoG2NtknlIF74
QaS7W9SZ6y9iz1jJD1kTkMG8wUwQhwfD2/vi50WXTZZf7QABVhB+fdZVo+3D5Vjt
vueEFHtMtj5axPZYm4qCvt9Sk1eRsifvTE9nO9CElKA4nrXUDSxu4aOjHB32rQ8R
jz9DARdd0U4bQuSUVoYxXBm6RIX/0GZbJkxqHaiZ2fX6PJwNXKDrajfDr6hNgAAo
XM5JzJ0GBHlc3JS+uV/7lxGejDwWDvedZbU+uRcomNc+GATj/dCf1sI0OFWuCf9B
/xybjPL5pxJ96HKSSYBxoAbVbPpGo6IdNyBt/9CBx72GkW1hnpkcwolE5t2s7zhc
fi6QF6mxGJb/Ee0MO3uIdEyes9emTgk2s223zD1MVkzoptB04hkjWR8AfS3QsBud
ePbpNpcS3ksWRS4QXoiJ0GpjMxRtLi8Es0kZRL/MEgaqN3nadDIJ38DKhY76CfdT
EY2q7QQ8z1RrC7ySbggNfS1AuNQI7ULPB5Va6VpN8IUgKGw3nxJwLBIwwldnKO5E
xh6q/puYTfHhgMXgZ9lT04mmMeZttfON9vfo/j9UWrEyZjYPbVS4W9hV9Kv+nNNW
eOfKOoo3fWs31sxKifMY+AETduUH9NSgQPlMgCukmATEKDsWLiH4WyRrgR/t3qao
n9679yS6QDEFEstIPaNgyfWHNH2PHidHHk7sQrL548E7kRI/IU4f/yhKQDQHV/IN
Gdj+vgqQYy3tPGMITz9kvCKS3mN6q9+upD+FKxEpk5/95W6HgfrsVs5oCTE4saso
fCBPBPBBv1tIPS16JfxsgyJgc9T4JQGLJoQ+mCs3yfafR8eNhM7b98NwsVgngRMV
gO0LBxc9dcGzUzaXMPSuimJxli7se+RIFCjMrc1zbLfBBGrpJgTc94aE3EiIysEi
PEARC2GBJVNPOxadsJCPLLVTIKcz4UL1uX9D1GzVqCVk8P9CduAdi2N6uhghGFGC
RYyXPqJ2OkwV93OcnuF5gHC/N5dvixGByI2auxBRGksOn/LN05tDrQMmE4EeRRLL
CRLcRjykMUjTAKMOdr+4DtBCRTr+oshQZn/uGm7laebmxTrqnAcJnOHjledJl0CA
e7BwKc4N8dULsgBu1XNVsCgdR8//PAqcvn9fR5Hyp0Iu4G7ZhvJpFTs2DVn4DK1n
ki1dTRORIH9U5Fi5ZkLnrwuqQmyXnSnq4T/iz/BJq8aP3YIt2EdZXLPdJhM1fUFj
IWCjs9uW150DJpNBIqR+UNYBpMLrLHpyHSAMSIHnRYyBxzqFgupJJzqvG6zT9odR
ZAdqcXYWWhbQn5+Wv7l3n9i87nBcSN03sA7Bc5X9X8CkNQtvazjDIsgBeALwgIB+
0+7+dXLFQkje8ORcIX1piSmGr1EUBeE9amE/QkNV/2EXeU1jdf+htbM+gIdG6NKr
f606Lx4D5HiC/RN1LAt8X0BzmoemEKUX2vzpXyt48MS1kfkK22EiNU5s5H/jUKs+
OKSYedly5/rkcwPE+B2iSdWZMxGTCmBE1BH8QsAIbFxRuAEAtbCLoyicA3DGJvTF
7NFqlLoc+ziMnA9XDlGpdiVSTSauddz5ajkbtXGa41BvXc1AIsfYmW3u7tb0HEuc
F9YQ7botALOWCO5tWItAjzledh1b5q/u0aTztepQHoCWm1jaYNd4/SN6R/iWMyD4
Po4AlE7wN3VoVZK17VOXR1m0SFYAbbxND8MdOStm6b+iyvf/WikwV6NcosJ2oBmx
G0Z/6Dpyw0E3Q3XFrqbp3xEXuPGdMCUXtBSLjl5WY/vFIrowocpqWsWqArrjIRlh
cVn4F2POXOTvrKQceOa1pTlUP1ATqfqqSGvnq+LI2vN5i20bZQWs5CAEewX/IaUS
Dp709RnwuLotYWaiHSeU/cE307o83P5/w8AjOO1DskApcPkS/xPPi0fgJ3mAuX6a
VFP5lMx8h68YkEk85kxSSzuNMvDs1/qcuVxRFcsRnI0y9zqvVW763HDxY5ycACVO
brnksG7eB95ffBzjcQdQpIs+7OUiNVWP8GttE7FYlFFyASy1iJrCaZ6v+8ixbYf9
V/J2vgdoYjX07SWmbudAk8rRz6AmJp5T5oSMWepgYQB0DAs2tQDCexLRKPmAgp4Y
NVS/Zi7TYewWZtDUGbsI/5cQIXs2w7wMrunkIdz9NPbtTh7YowsqrL4Zcwl62A1+
hGaLiiJNO1Q4SWmEwG5DnjUM9h+OkrIjJXaje5KnPaldPsgezsF0/12OExMW18ZB
T5Ykq8r9UzQhpdafKv1ahQry2zkmwfmKZb/yR2ho9BoCiTLPdKa2u5FsLOMgiHtU
M37qwWs0XV7AcJ9q7JGbKbaCxxQ16bbfX5j/Qo9BeuCW8JPua/GPLiKeBIi/uj0q
osT4DWGnFApW1+pA7HKy7s+gwGnI3mJKqsuohyBr1efIaENJC0lyjNWR+OpZnM1i
1PANFxQQawksvB1oertoZkzi7Y4DFT0/qg2A3FDLuUH4JRv5zDAFBB4W+fFJVVZp
9J2LjqsLTnWiHN16M6i86wA9DHakbNRodBvJi/H8twd6wf6luskEWtaENskpAU6L
rizqnm3kckWgnurMqFqyHTZ2OD1zN8hMZwYLa20Pp8RYT7/WuCZMXHPc0S9fyFtI
FzT/4Pn/aAp6QkBBDx1ODt9GJWQq7y6GTVxVYIjhDV4KHpkBEuM6DkTDPlIewiL7
SEqx3UFV7mtz2bGDV0hhJ1nU3hEL2IpgxvXz4M5bq+tJE7V/Dc71VcIt5nL1meWq
ordeqXNsnMnco7IMBQxyJz87zIWk+s3kKYjam0sB8IyNyQVHg3ilaP8MHT7sXBv1
OB0vCiT846CWfz8Hi/Co4mhwkt2nrN66OZqUTRXME8wlrBPHwvLIv0W5OAa+sgNE
9fZTlym/WTt8ivYthalKbx6sTmlI/io3C1urGj22oJ/J4CYmV9NCNGYlWFppkibT
U3jy0cDjfM8xGAa+OdPUEe4TfjpVitYUW6iOVjyfVeDW0PdE4/0i45jLVeLmYmMr
1jbK2+wJxxlf0dLne2NwhwIuKyddUEEv9jiFM/D34ivljBzmOxLdNjswHhtltwdW
yFe5Auk+m5En9XXqfzhZYd2cwAebuGg00chZXB8zDUSzmv0dRgXfnJT3pyR4Gfeb
ftM3248/HyRz85PGgDFDkQ4korE3D/eO+lwoGrIrSFSP7sTrr9It0S+EQrzf9sqB
BpP5+QsPPw0dXqMSCzLiaGpuVyjVTLy4ZmMpyTQ8AbHzmPtzDmb8dUPEEoZx9O90
BqAtXrcGUkFftc/tGTELTF+aV01L/zjdypsme22w/ydrhy4+IO+LNg13UTll6bdK
SrTnZOMVbExWJzQ9JJ4zcsvQGND5u6jkdpwrAdEs9Y7EasVOioBPWQP1JsdaJs1G
F2Cf3diMPco0LnMO1G4mVFeLkHiuyG7PJBdp8mYniJRc59BLYfv5zVPwIttcE3HY
tdcjaEf04MGl/3xUGSTr/axolsrK/qUExrJ6dq4UsZkV20SmTbs363hR/c04Txiy
Raa/od2uYKyHS7Z7hXjVYHCsJsyKQW+7cmJE2wDoV7u69n67ErYAT6VzS+kquRzK
KVJPXuLFhAhXIs+bEyWazZTylI98J0+/9J5XV1FZsmyVOL/gwXgRwRTOHhQWQY5k
HfN2PGIvyIdOa5RBDnehEVFQebDSZQwSNTEHvD/Ah9Fu49oODU+N95dunk14jicx
9g8JprIlRk6AhHo8PtvvVPr5A87LLbyWLOiYUQC7O2F07X5zsxpI4B1Qe4f8oKH4
FwAbJL6EWwNDNBfggwtLjgGDlsPYbZDvjgcaldYedQb/yhrTfE/i8+6e5Oge5xOC
jiuTOdbBV2flWRH9DmO8rd/RgPJy9qJR2bVxYAsRwaSVOjJsVEyp6VBAXeVAib3f
KblgADTAnuTpwSXaWO2hq4Jrh/0dopIikvnlpPAhDzII/gcJ0Y4v58WVK4uHaNMt
QDNUAnNjpBJU4S8y2kxd/qqMYl4yBSocRDABEAF2c0vhzEXjlO8Cuyc/5MAW15Tl
MUtKzm4soAMreqH9txSQ8VRT0Jl2tGJCZqUhzfRMTVQ8N/LIPsZOKJgjBobMkHJh
BjrHlWUgtQwJS6CpsKqA5sYCQrxGXuAAi5qZBu0Z7VuIL5aGf7NyxnQ5ySwjbEsJ
EiVh7VHpJJAfRs1bkfNTv/0nUiYuNmpmHBeD5zEcPDJBrH0HVBHe6rPGYYH5kcdn
jZzvqxT9iipp9S/9gyTt048g97RAoTBPgZ5vcALL3jN7WB7nVmhA/3JHjlDqEgSo
zYyyukip0HTUy8Ghbgt9CS4Xr/ArL1pFK20IPI0twAIFrQR5b3KHoH46nrUYaWmw
oO22XVsMy/cbEhImM7pvAwjh18MYWI54ZBfh3GR+rr9lA2AofnqMKmMoK9sUVGQJ
EtBZHARU7Bd1ZlCeODiemZM1V+Lzcv686BruTDi3md31X5KovGBSyqbMjjBUoqby
bgTujWPuiPeqQZ1etbrJ94YYJs65ZgK+YB9BTwFIuIyaJyjP1P2pPlCzoOzn1SXd
8mAiYrkenyOuDt7amOGqlQzrZtkjz2+Tp7zs9uK9Y+9cDAiPGZYj73NFxMroZoPz
CLsVKPRPsChe3YbV1d4gu8SEp7gHuPUMww0Blml6gYI4tQJbY9Jdk84M4WIOz/lz
gAXREPj7h8T5sdM7U06Vo5j6WAOu2IXuT7x2vlxTnshhwisanS97lJU9C5BDOiGo
7pf0EP0EgJGDRP165M7t7uVYIMYZ27Ey7Mp7gM9NgXwq6MY72HtN3Jvlt/5I6lEu
djDL0kZlyAGEnZx03zTzKqNhM7hN2Zg7NDp6lJNGGDbPtCJNkB+86MQa5gtFPzfT
WFJTB8fnUGOLmRlnPMnktyBzzsW96e2yz4joatAxRJ9iRWJRSYj1F7zrVewnPz4D
FKBJ3vUPNJgWMVx6guqdHwXG5oXLm9RxpCD+8N2IlNRuAOILo1txZrN7XF8tBPN3
kd5NBdtn83qVI3+s0nI+Hd+G6/UHJv1THVvRm6DPgWtqFoVFAMKPyAYQ/FSpN7rn
0RjiaquHtB/rNUxvt/7TK9nCz1d0Mxf9QqDomad+vuKCNNbDvpsWc2F27hSamdrw
3jE4oGU8f2loU3Sdd4TwBMG45bBt7DaJxrFV3GODKOiBXhPtAPDSNKnH0/9hXeeb
638W25B8awH0a35Hh9g8SFsnQjUw28F7rnb1uovlPk4bEb7UbXybvrt8afZdnCCm
aZFnjk7jhXlUkAUGOq+hWkOrO6Qxm+or8HaXj5RUC7mCct7ZUBbJU1zYKLtyv0kA
aXGwYs/bCSPNSV4O/g7eACLaNMOZfE7ohJI5Rqz4e8pSs3q9vitl31/OpSAyuhHW
HPOIeFeLExGZKIVjKXYDYtIXx73zcIbOrsrRxUxHN738nObjhQkJkf2VsKER1G4y
xOc1eI8BTDK0xg9HeuF+AdNCzqhJnubj6zoIApVKfSL+DB1nNJZ9mR5UnYtqdhAh
dHxaO+b3NDOW1J3MSKp7ThIl8F+2Db0X4Zz7qbvEUQKihjxU8O3VxQzVWy9mdNrS
keOHt99wKtxcH39ITVpKiSZaY9fez+KGOoHgSAYk1me1oAlehauxkXVm0Ow2DOSR
IuUBduJ0eXa+gBXyE4uo0zP1GN5JuxsO6sfrP7cTvK0y20Bbel3we/Y1azAadXBq
zQ01J/WldGDLhOx6R32hYrm+7XWxWgZZ59L21uRLof8SSVjyRg3HJ47lgr9GB+e4
hlR6gsNPHvxzqrkjbj/qhCGkOQHmcfi5k0ptGeIROOM1nhOOOAIUlhMv6t5e7QKQ
PP2HvSzBMKJvtMGatNwv1pej7RcPjGLdwZhzWkvS+Ju8nIBdmJtikPfFT6T325LT
gRpJXuX2dZKdYgsSlTAuV43Tfc1lN7af5+hV7fDaoOXwwrMAmllATD7xksPvuCiD
FsJiwaySTLtsuT1pkvKSQypngGQN/RGXlgT2XQuYAd9hPM36/B4nGIRbHaZ5qYaF
TqpXP7AuXyDK5gcM2GVUI85ICEmmI1j+tcPtZH/Whut1I7dCOqMQY8eyMyrhuNZA
2sWx2NTqI7IFOmP/C9JC+LuYvagx36kNfuzdj+gJmDmSeZSgioLsyEO28V3DcQbR
rOyKV8gB4bW72sJjY75cDQuQsSYDJ3ZFNToBtAX60eRcBdXP7temPhcrI8B8YaXs
Rp7nRlkwVhdRtzZB05mK3Cdw1K4wiPs85biSovPJQSteN/cKQ7jxLzy9FI8d8n/A
eCVv9qly4BgisLfMt4AcPF+4xhrVHAbCGGSq44Bp4XRSARA6O6xLniLvO1yqkrdp
UWoqOr9z5dFHLyTfLZA6VzadityWsYylOBEZVW40nnp3DPEkDi5H5/adI1u0Hnhs
JytOZvYDf46Fb5nPpLkAwjhRXwPz99QAqa0oBRczOWKIud3l0IF/Sy/Gvgwltuz2
r4Uk4T+WgOFj+rYlIxuGkyB9wDExsN2G6j9moxVdYm/2YwBeTmsRQnpWTwmMHGTI
NsvyXpAdAzObOGzYuLiwe6uUO0SMYGHXoNR07bbLB0OaHiKzQiL0ebfjRNSqI1IN
GruqbvXAk2eqs/HgtLUEl/zZmewJ+2RCG3e+C9QdeqANub3Q4wpXu6EaT7ibkRpY
mu14JwxyMiPtfzoaJy0wBzW8MPyb4Ch/E+dI7pyeyY/K5YgYdncMcSQ1Ens1MW0B
Abp2gaxXuvHflPRunycV56OCN2rq2dBx7K0A/SMwLLbSbg3X6b74/zyveiK7Nv63
jKPC4WT36CAebORFSdvM03gOPBwIrh4lTQ2643bugg7VmfZrOnJouXIKkG47cg9X
1BJ0FPuena8w/SpVgzdDuDoJ8OoTkVV78mClPiZPNki6KLbr2+ZBxjSuMH/mczVy
fKpjZHi93FNVlT1tdX1NpNUa/mgPRTOrCmQZZ9+IrUqfKCu6mA0DW5KIKuAoG8eF
KS6GZvE4+W+LXtj3IAdAf8PqeujAXbwcA4V0GgjT4P7nXQMQY4Udh3sGc2YzphEP
CAiqqjVB0Yn7ffXqKfQeGRlUMIYAEXuJqPxiFAIZBNTGfaSS+hjtuHpJ6fXgn0FA
b/Ai54j/BH/MKEHfoyppqomEWYRb6V8tR8ZqkJOGHZ4boUzNSB9Akw6U88+qGbQ2
ea/sD21Tk2K1x0NK77o9kGMeH+YI3B+ipkq3iJzhonN+njKASaghr8D+cuoEgimL
JpiulawHvlzQ6PuADD4KvFxcFekiAhSrmxHSf9Ij7g6p4g9AWh4wq1FAH+BF6trh
vqpONQr+9mBOn+yuyFh4j4h8JrSkMbdA6R9cJEbtR4OYhtQc1vvApk4YYOizis6x
P8qk0ceLgCQui0q/U41JLpJG374q2dc46eNh5eXz2OoEkoV/yA5n4q4MWtN0IFMM
s6KUYoAU8UtkF4CMkfYXTmIsxkfD91w/zu7cMrdWO0C/MrZr9aQO6NqhJFa1SYXE
ZmR69NmJgY/cxbXwV51hnXepQNgZ2yfgVzsuziBBONwd/84C8i2TAqKo0T/3IPmE
D1i1m0vXPRawsiFdCyd1ol2JYEQk4+cHnrCW1CtXwHR8UEjaOP45kWif5rZqA496
SePtBK/IUSpFrGfkPVJla2sI7UPuv7S+El7R5yzXF5vduOc+etrjqCoB1ybQWoAL
hcku4KeOHjHXyiDJPB/N1N9ajbgtUnAu5O6mNieko/dsYCtvjxKSN8hynpZ/QOc9
CB9WLhgZbQ0s21NgVC8Sc8rLFiDD/YQr033kO8AW5awBWyn6DZm6YCj/IHy4m1My
zDr/UlW9tXtRjNz17VEnqfxmz3GOszh8bYq9lA/bxmNJvd43kcwKnizWtXbbcqMx
ei4LGrjeB15UsY7d9NeoeRWdQ/7cdhqr5ybdU1ce1dK+Qw9EKm2omhSeZa9zNjtR
Oc42fA3RmxJYBYCOYcS0xSnfB1pRtZcI6tEVw2syO0hghlfJfqh8GlHWo4GlPEeG
0wu7A+jU8Mmf6HR6ZVncAHKbY5drfOyiDKrizk0PiGdiHxDrm8GP9njbuqbLA8GQ
uoOfhz1qv0s3tmUF0EJJKiNsGPmXigiJCXM++HlePs9SBvy0RwQdwVRU4TzRC0tW
ihJBpeJWnnbLbJ8zpTC1NJxXXnX9kLOQlJk7+TQtW/Pycs1dSb0yrzMBM/FrNOCH
myrTRa4B870+iydvrKBwg6EdI2frQ4slfx696kBdkBtCNwY4StqLy1hXGVl7AOvP
Fiwv7QTSvgLxsKTbZm9UHuWqsurFT0J8W+Va+5o1C/HIn3MKmZhdD65OIC373zaw
dq83fVAPlIhgZ5cfUwLqUFLLBLJr5IzsdEyF8SFPFVT0djCPmBlNfbnWZBDEtnuX
MezBtOV4CF1hg9lqJ4TFCrx1XWvTRnmL37JrU44jMyUUG8WOai3MyKNuiaAPCnx7
GhnEdmu4Bmv2cwQ1Wc3mfm+rJjBvUCKB6G/5zwQazvVtaLjy4Ha/c5knvzahjD9q
HGj0imChpRsE9VUloxGgLd/9cMhxvcbidr3u0a32UA6iw8BX9F3ZzpH9qfVQ5p9W
QINHhLAiq06UeIyeNXmFgKDZydgVrahwTZGyaKMBt4HfPok9Gnr410QfhgKdYFoy
wCrnkhgnZetp9E579vNw6XkW+Rztm5g2TpdrB4Q6FUSnMBLC4RjwFQVVLFs81/R/
Y4EmJdCaABSpHDBjM2FQHRVL9hEb4y+gLK34XnX0uY7qjBIjFoRYjpfFu9xwmFu3
8XIj/ACvffrLjpNm/2SL3HxW37LI0i0B44QmFqJo7bpzNfy+Ogufitl5Tw9tGJtQ
XvzAMIh6BG1TMVfzye81P/rTtTbi4PkUIfZknTK5DGjSxmVfjkyvI2QWjKCUMGQc
2DL7ve58ahV9yv9cJnnx5p4dkPzfqgdAX1Yn0+o3Q7ay7ShXsskZEahKmrIlQ5cI
C82JUxZk3DqVffJGHTfm+DR/psuVq+8vCcQjcdkMdPOyXLkiWWNFAEI6MSa/MWQt
MrETA84o8uMNskX7V67v5J7Uz1n2cfYhfhwQX93AF6WLRrOrpm4UhmITsVG+pH8H
I9WIT8f3z6SPsoYuNAmdKM2vmh5r4p7b6dQlr56zW2t6ZZPdTTleckqciVGpGrur
+yfAiuC4tka+RNeFsWtRF3CMvomiofePFwPLe9dFxR3fjg2LQtWKHwM44lYOzv/1
yOVaMXbpeBastll2w5NFvWDO64Tc8cnZwuP8kF83mYkV/Pd9XSk33GT4ZFSot60i
HdmVLt7/mQ48NeiCkTjXgEoYHFliybONDRCI7xVbCRq8zYyUPKGCx/H2LNPzzgxZ
5lgp9ppxZ3h4PlW9HOKT8b8D6JIBqv/mR8qUO7OqUzVx87gspuX+S/9qwC3KOKcJ
9wUn4YzhmxCYKMOVHqb6ECIR1/hm3OIyVZwQiTuyoY9QNP6Lq3XJsgdwJF6Fmz0y
J0U4t7LKA9fkzgmlKOxDgkTW2Rxn0etskY3e2nrO8jPdKslwoVtw99fbjv3u6IaF
0mGOFZ/NekyFyH8fERYEr+HLgrmgfMfxfMNO9lgvLN+JnHuqCV5wA2z8Y39sn2BB
0Hcg+d3heBcj+yQ/IozCRgMpXrU3cHMcWP926vPxHnY8sQyOPPRTWgslQYqguDf5
kbJH/aLQW5Eu+OgmRBf/qjGXFrb0DKE/qgYZAMrg6ZzabyBq/0P2oyYxd1DhU5Tb
RvwHdDUwVzY6wvU75x8znMFH8GuH0ooKfPvFESSpMF3LVWQoDAOvXzKX3T3oZIjk
oI1MnDkQ6zbc2+XaufvG8hVKBNFetZHH3WYEonPQ25W6s5micMk+WBM/hNiUzu0Q
pzpF2uZ1Em7l8KpxzXlJD5xtF4IR0nf//SQyOP5NkxKXIQsRkzCNVhQoUWw+umyP
k5uPrEWZrZwWwjQmLjVA6gM+4VNm8rXWv7GD+bbChJd2iZNXWTcT9kq7u6qTLfof
15KksQ1tVZAR7uQ47PMAMtHtDTt4TaCe6aCSbj+a9TQwooA2rPt4jBahDJ9qNCc2
nxJEjrjN1rMP792l0gvEhkv2qDAlewpyEa6Q6i8ABF0/8cMzuQ41IRirerTX6dLc
GoUuC3iENXlHF6rL65SZoOsvOeRA+EteXlXgbJjzjZiglynFUUCtJE6AzQG9yfGf
FRS53bXnozXRlFrRJI+qG00TZh9WPETZHRAy08fRzIbNoJ6AE2h8PykiMIzNS7LM
AIzeUByEA7r6aG41EtUTqsaMFpGCR87FfdRT50m846WZerL7D/MBMWRK0WkNxQw6
tGYnjbzEN0dIlxKlZa19jyosuL4Nn/ntT6Ox0A7bDb5+xsUpAJp5AUr/7kkhDfoQ
QoA41wHHetIhJJ23c7jkqJfd62860OAZ4SO8iZADgzc87v8bjSf6YMb4K2WmI0hA
b5fy2pVEHx2RsJIqpqTnyMIOAlkEP9vPt/HtQS7fYNrqbFg1xNsn8wQdLgsLf28S
VN0DYIYVHWMH4JI4/sKJ4Ug4lTcn5LHO0XxHPoshOD1MOBNmxmTl3zETtUUjlYQy
s84W2cBqDIJfU4auz59D3J2isc7DOZP+bRyDa/7iJVCfCKE4vbzyUy5Qus96IUS3
Z0td5mPVklkanj0OZPTAXpdtk7Pjvj+tivUbN0oG/8wVYTOP4lNCV2QeF4ssPjzI
gqb8tIRHw0/JpxpXfrq15uutxLffwE4/xWSJFroffp+8X+3/gMeiATHHmB80Baq7
+pW2fGx10wBCB1cNDS+GKOLB+eOhy23RbB7keX8dzw6wEkc/geKApH26USzTBp80
kymcZxy1nKdPSdCMMa1UhR0namaj4FhnL6ZQFB9iZyofhOgjVzsKKspgjh/JisnM
A+rcgcLRkeYTfxIJsRrvwsRYknZSUW+J8adffn0ejSqaWtDZAA9rimDmxni2ksCM
NgCChB498zTGIIsxSG5/0fryRS10ahx4ZALXhKKai3nbl5VNW1P3HcwJVLdG2cUx
CV+uQArFpCgLsekFe8SMJOWqNi5x66n27xMeZ794NV7oHRU3T+q/XtBS+jORC/ub
jXFarQoNkHNac9v6bug4SvhTj0nZUWg5OOwa78wLzMrKaeMGA397CGuYSzFzf9dp
WfvG2uXXoRc6i9JvIIwAF2ppYQLW6CdFG9OiwnwfjyandnS15MjH32+dyChpb5sN
oAF/E6XXyhOkH7wErsl5GDvSSA2fmzs4LwdgeilkEb52fsANMO66W81VQXscZrFz
KU/2q2IboRNT7WDwjMT5S7RbPO/jixm1qOVJGG7GqBG570fhg98MxyegW9+Z2E6q
lN6stvdQVQTdq88d0xpgsm3SdmZFxv3G9AXzvrR18Vq9Hd4k4XyyoC2dYjOEC37K
tj+grlzZMhahJQY4+JsJ29prbz7OH9pDO3kkFU4c5zPe8lhPsnuOldtbctIu5I2W
LiOmh5Yy0CTwcCCr6OrPRpJNFY8QiUCyWzNhCMnRja4XeHi/I4yQWDpwa4hympQJ
1K/V3FNvXO8Z8U4zQ0f1p/JIJ+1humElEfw+dQZPJMGprSu9IE3B/eEPb1ONRk02
EES/XPCxsAXLZ704RqJI395A1p1PWqlm9Lped3Nj4j6+reAQ7AZVbIUO3XGDUwJd
6JfYGUbK6gRrQevjRXK+SfTP/r6DkXqw8pPJCCgTpOYP+rKum2rMFgAYnnCC10fK
PUEjBThl/5oMwv0yUys8NB4z2ygwYL8JRJ25PBjxEnDpaxJK2TMQ3L/U9pbQlsiO
zY7LvARhORZlDPCiAB86MIkj/paxsXxkic42ubk3Qlg8TKqqo6+kl83D7HxEKeJB
lrTaEjXwUl4MDJLPFEoWCQPxOOfFlFCxbxRk/9yvIKvk2JBby4qMjbOVVyRkWrrg
vV6FKxPMzOM8OBteBeezfw3f6kd/whRhjg0OiO/Hzl1KuqVnnxDWKubQkeNlrMdZ
xfsQpXVB5teCA+LCiIJcErb3+f3Q+fBKvX0Jei7BQ9jnm0eZSlaL74Shg/UJK2Uo
gHl0JuHTYZqhw6d7aZRyAQrM6wo5rckli/OgYaJZGhSOydSRz4CiWtCbuOqehRoi
nCD+0UVEkCr84gA5WACL2nHgq9LIo8K0SJzEXuFejWH/O6UaXg/F1bAAk0nDtRwX
RETEWhtPTrQ9HYFgOcjJUkJWNjiwC0LWkE7Mi3Kd3KX/6VQDR8A7NgoC7XfZP/B4
To8eH4qBLsnS3WmQv8b/3ciNCCeGxmRpOj0u8uQcG5kmmEgmgkLPxbRcYG+DQ3lO
LH5rWQvn53l6W4bLnWtDZpRcYrOMLD05yBEc6EeaDoRYE00XSCr0LLlbrl0rYX0e
73tpEl636o/ZFjRxrbFD0G1qsDLNGYO81Bn+v86dQ8vzAulrxc6HcqwMMngVKyNE
HjklhzRwkbL1iZH545m8RKGPnepHiA6eIYOdGwHeYXlKKnSNux4k7vYmMQUIzsyM
moFYSDVMHoXK6mmTeCDTe33xH4sU/nGht2h5k/VN6GvpWGpN5I0qQgGhgBRsh5DN
IghkounoQOK/mDbomEVDXaDohvEKopmFHTZ3N9mZq6sujllYRWC/wf+Xb/LoXa7r
DYTCAF3eHuWgBSbr6N2dXeoie1oaJj40gK99JacZ+52wSYC73h2yAAQXoOTf/PD7
1gQ29uPSOo0saiBD/IC3x0DDl7AY/qASQ1vbQ5kZBG+C21sK3WVtv4A+0Z0EHk5B
X3N0/Yln03IjEYgCd9qVkY9kG4NDsRFSQ+xlRZ7/7lcbXuxP68xGeoBSppUYgH5g
8NU88sWWMqwg349oMEnmOtRe/CfwSjN+p8PUWUDKte4oZ8IyNvk40//8ligtJG0S
jDoPH1qESdE0Tg7cPK4CmZjW84UE9oKOIoIU+RVW596Nw5QoCce/V7OyevUfJ5v7
rD3FjkfsIfXGqAoczrBOeCEhHPioKOA/4OlWusN5onbfGocG9DvE1U+HXP/e1w/E
fSaj0vhZ2ferMuJiBtGaqlNH+HV4zyZgPAjKSo5H5MY8FmoMA11skm2k+aqeE1df
WkaFewo6SwAHoMiEI9MRq55COIqGHZRdjSnkJzWJec3922YskLHEugJaGTCUQ10l
fzCNEJl4RMcaPu9aFrQvu0tVwcGrY5m8GLBEo+DGmcLE22F+YlU8Jq1qAdrcoN4X
6YLaCrG7O4oJ/Xa9L9oGYqlAZ7/kCWEzNyjR5J+azW+BqBc0B8r6aW3JRhupsYGd
vDO4wNzLJq4NjXLZppFXhl1/1uTO+ebdEzU85Ne2bSq32CLxmB/OfFDJIHRFnO/p
F0KhAU4aOB2/+F6xkHzgQYX0BCaoZfP7TyVxh5Hbx4FwEGI57FvVEq/LJs4AYkfZ
1Q3vH9KP6zSW+jQYlNbUsQvkuw5U8Zqy1BAkwYf7cAj69b7se8RTdxrvKOAT8yMt
dk1O308y5ma4Q/8alZ2XZLJoHfZ/dbKUasNrvycLSajWgeXcx/t7xXrM4WtQr7jG
QIrvRejGnKUIQuwEuum9v2rn4XnR/uriOoeQ6euy5Ebkn+oRHaZ2/WVid1/gUxCC
k8VuRV1ABKC/7OHrAbmaNzfVPx+DX0bWKEsooBEdyWE87HfA/z8urPdMbEljrAPG
mhmFeIDDU2YbFNrMt1PKE4XMaBht26M0p/LTlzT4fwfXw2LNTi0MCL25PfkFTNvo
xfULa+R6/pf+IjbA17q/AP1NiOabN4tIhd7ZU+ShaHMFWh8g1uPJRCa9Yejz6FXD
gaWnyGICHVjVkbmlAiLwETxVcIMRL/g67b+wZ1twcZ9ToRQuYKKQZsLnh87UIv2z
L7nMQFebZIooQz+JQcWW4QgbANWh3QhrLDvAJkQwLftpZIMEoeJvJGDLAEGaqL1N
cpaAvUYNFpkLOmSVKLsTMilaH82BsfO6ibJu4nDGycKqp3JjtrdT5J9RlRipQmSl
axAFmrIJsySl89vGaHWXsGHX3wRqMFZjHPq/33EcqWKgZOjB428ZdSlNk5WBsrBw
twzD5kyKfw2RLwrwy0/aXp4FyRamE6IYaiDx7wLodRlfBS6UM58IRPKen91WC9Ax
NA4kL+50zn/6HzzCvNN/+yNsczjcuw9Vmptr5nTJGRFpjLlwM7dwrF8D5DJplgF3
qz+kyPwdooreXGqwGmV0WiZabyS8MlvIaiplmuSlU7e97p1VQFkl5SV2rTqX+Xuz
x+8MikfXsMViePI9qa22lGAhEaknhcKCwDU/3BUSxkGftvDfoIYss2GPDR5t5/3f
80JrhC2zluYMxnBaEtGo+Ti0WkO3MYICzIBvEjqGg2P4Dhdd5AOfa/HRFuihiYod
qfIJbNC72vGRVamoLYjuLxABQ6KzaBaiYaqsy8q4MzQJNHGurUGWkaysTfAvOkb3
TVoPgOD91zh+MlQLDDVSs2MhmhC0L+z0XWHsmiIoujugfIshk2qjl56XYXuSz4RQ
PyOSLxsFcWEWNt7MHFut5AwPf1i1D+du2rO7xlResrqPA/9gC7yevuNDt+QPQ+Ws
roFazli6ksq7Swa6XJJxJmEcbFC2Aa7FrFSgJCvOOfK2/ua/8mfSWLI4pqVRg6St
2MwqK8kv/JfRPFo0O1IFGLpNOT/t+P53i4GGLzqGCVttqBr9yEgh/V7FJjhsOH6C
P3KvGYg4pzyCcf8l80sfvZba1moKk6ltoq+c/JoUzt9APXL3Y7jz3otExzEfAsh9
msTzbCII8+sOapayLtzWWwxcRZLTglaB2dF8ZG3oqFVNtY8RvOy5cKnsf3yqrBhY
J/daM8aZnFdQmAmghVeHD3qdCnMsBceM2RCHhGm1z3sVnUB4/ImyWe9ZbYxfN8UR
mp6sK3kcx+f5N/FrehomjE09ogsflkiD3gZ+P21cosVFB4hZCvvOKg5dceyDMjMc
iDix3axVt+H1F/SDdF79J1VWIRlMd/vUKoYzRH79odid/tSUAnu29dpMaxlvRsnB
D4xt2g8JsNRbFqttW9gQC+gq6Jczf2qvvWgBsr9RntoBd4qiBQcBUcGHrS5B6yeW
MXisGiiQScdYphK0CfkMncPM2IKeat9fAHhZQJmJrEx3P/KtNjtL5dZTT4+iGRKC
Vqx23FCBj+7aqfC9o44tC/mTe2/x3xkjjFjj4iW/ISgN2JfA+mS3D+cQMdQ8xsNE
TE2VpPUtEEkDjMgWNNlUiTx6tBQJbEElJdbDXIMeatBVUkAuKDIYAxvEoG2SuzMx
QSOQqFoig/w3YVPYhYPoCLPvXxyqMIA1rALFdyXV94L2Rd6dDmtUiK3QaF+sxF/Z
vFXlPUa5rbHSjsfkZvJdGPJgOLSiVxeCLc4/hlPVPqKHZyzfV4UTkSLNclvcnqrH
GvzeSQPcgtVxktif5iCl0JTY85vpsmQY/Gy7CO9rMOhlB3c70pHTckMhAYrWKt/k
D9GywFmw9hoWI5YnYeOymRCLILwnDg6g5ud8nGaTg0Vd6rd8aar4xbJYwpS6gSLF
OWBzfXQIQ4b9Z6xP4j1yMIPgRgtZDgTu191yXK8UGotOlTJaZrIeDTuaBkMvUh1S
jUiYpEUeAT6abCZkqygbgmiSaa7DdMo91lINVfPhktm9cAV29d1ZNjagWjPB6nQ6
xJ/KeKjKSPwwIK4n22GsHs45vro70OZAa/pTHYe7Z5tyC/+pkL+OGeKtr6sRzQAy
ZUKl0DzM9IrAkXp9kT2C56SK59+o7ISo0gVm6KEyh2XOHrCriL1hqRVYpQoTFF5x
7Ii1sEDtjEmROADsV2XVfRtvtVz4wr+ASIpoYum2F1vWsqmLuE+72q6ux/MV3es+
N85KlkllcOyJvPPSrkenJq8QTz6Ph5MkwenBAUjRXLOdH+qRIiDJ40FPQpd12Sa8
KjJ+1zUfKOkkoQmYoAMsQVd2/jAQWkFv9S2akE9oY6iFoPBVffYiLcbwQG43VcBi
1GpNbwHEDYHK8Dj7h3xuFttRz5H9y6xoGC4x4xlGt4qTqh/XXNbanHfsKw/CD2qE
c4Mo/P4Gur91olZ33cjohr3TXx5Yi6DuKHqTJSDxN7fGexGh/W70zOfcfwzx0Ugp
pMpqhOuEYzUYJ5ME0H5Q33OQNK0GjiOikDwX82aB3XLJqvG6pv62beo1aWdv+nW7
aElJnk80jvESGH/7mT/fPo8ZHTJO1wTk5Td0HSbjwbh6q0/K/OvAqA98aO5RXLDC
6UpIefGRUMcO3reIfB3M+l3HC3My7OlCw2XWL+IzOuDEVwAdZAvbKDIEihEX2Xn5
ENxcFgIlFwxBufe1NQ2uirG5DPO0O8JEsjPWvDSa+M4za8y07cFsTbK4KezIP4EH
pAV0RrVHVVp5JNIHvJQSyaxYL6DHSbaPHgrB9RMpFjXV8pVkEEC1m+YtuGKDlOr9
YnNwIJIWlLfUCPs39m+DKrYvwjGFkQBzA4HhoIJ1o/PsUXrmK/c2PsFnsFUVAk7D
mZK2z08Cv1x5+PbYef95qEBrUOam7QYMLWJkWF0YE473kybt9REPG7FIUAxScnEc
Wnb8WKUcpsf38HgLW0bLM0ir0jL3BXJMoLmgcw35qQzzHqc0ALAf5/D/zMxOu75v
/fsfVolcxbBgOBHyE26DLyq4Xh1QYKVyL83fcQYbdDyD6gA9GwRMyrDGxpbBAoZN
lr15k5R69ehV5/pLRQiQUUTGi2TI8rt6US6DxK4pPV3KJUaFHunZxNFROEt63EID
28ngqpzeSuaGROdRKACTs4YWtD8qIGf8cmiC+UcaG4Fr+fhVLj5ckr62ylEjKOt6
Z9hdZepR6sagEtEgfE5goTsOZUvW/XsfOXjW3YKTEoJvqt9JxxXTv8rFwytSo00d
KFjbi2vAp2JL2sGlEVcvSwjB1TQRGohBW+hOChcWTXdwjjarwkzNBfyIErhra6Py
fjXDiJWR1Er7ojVE9nFH77+0shIbalxfvlg/KmchuYHBLVPJ/JKfqzDEUK8KvNlA
+zcJyh9YnQ19SERVhXhqk6C9UzV/hDFvrwkPS/N8OFcYjeIRpRylGI+feC4NVu1h
1r0UHI+qGRx4e0LjRbeb7OQDeAT9jyFiJppmzM2hsaf2ZL3G0dxEsM0QM09GeU+k
FwA/r8QeAu/ev6p1bFbGT0t7sgPEeig6JGsXYlVnBDRlt1C8tEWZfF7ssrN4KRZv
+oZ7HjvAai1u0mhvk/kAnKMrlMWUZhWjQWnW5Lfkkh1wVG7lnJHA/bZUGf5l39ib
tWK5sq35K/z4Clp5UFRFYG4TqMT7vbnkzCYKaXSEI7W8lda4qTR89nc77rnwwaV4
ATQY3CPxQ6an1mWxkKwGvFdpjbAbhzfnYgNMfAC4zs3CRdOITURKImSNnR04e7iS
8fmIVs0e2stwMzFZL8iJskn1YhZ/3EBlRbgzyaSiQVH9Hm2T336mzlGw1/0RJG1w
DcBw3xO56gCIPOScwtgOH5DNQGCAF2Xyd7xJM8v6N2TDG8pY1MKAC0Qqi8rK7IFr
ag8srWWLQsx/v1eRSjDb5NrvglOctZ3VYQCCPzU5ynlneunzi2Cy2L9IbpoRL887
7boxAu95odaCL67B/Y/r9CHTBrjhftjh7abzGlR2vm/oEskWZqTgsbAejVUG6IkX
2Tu9u4o4AVrfSMgRtPRQXj/tc4fJmF16Lk/EVEmC8pD+V0iappHsVdQ8+fh58TdP
Y9FCRpbWxzMpebts9HXHMYBnRplt+eXSrjs/q37LgS48AYRaaa8zJHV0EUAlHlEd
2fEuKghKE776djYk+KTGxDPyB1imuBrK+6Cv6lbN9vfmAp81xM+c3La7R9rMwfHh
J2qvL1tYTigHZIQlKuIDmrxLwR6dYzNKp/+JdrlWYqogFTWXwZlDC2NtwV98nH4v
zFw58hSGb1o1IcOxIYd9gumLFq09/b6w6kWJqxeeJDkJ5zR+MOF3mlcGTEmiExtc
e749g8/uYLiawWQPo8okHiBQjPfkCs+2oBK3bwsD2qIboDLEgyXZQHjXJWpJD0ah
+E6rez+f8CxD1H98gX3beA8/yrnN5F2IZsV3UU3I0zzCNnrGr58bBgcguAe1aAhM
0RuOAZnOGO1wWpDx4YDFyyroNt92IHJQYRbqXaujTY3wQpM8ie/ehUHWI45Hp1jS
EbYhXZO8H6eV8lbRGS4mnY0txO/7NvY+zl14M3XFXuQ0gRxsuH/hKniVMo89jerm
dUSUuvjBhuq+BCd4wONczvNAvAIGRYxw2Qg7L8gP3HToyZJCRVZHSRbm2NKGjBp7
PmAOQJ6AToCd6bnMUkNTfMTVmybWfo5l3gV8hzHzSZqCg8MoFJhq59HIjnPAnFLw
6+4xMT/Lv/pgZkPRI259zn/Y4V8TzlXUxI++7os5gte3wnz96TkoCSCLI6fjEhE1
GXtLLEY2p5jOQdYca3WBS5xkoTFnJqhup211xoXSp7UT/GUY6d10gc03A5DIxJ/Y
81i2GD3dtX5w7P2CuFtCmzE5pcKXsIl/H9lTXMpd84uBX21FDYAAO5qHxhK8s6h9
hoBI20e6eYHpaD+LnOs1LqJVepJXM0T0JrSS53yoB/gIKR/drYWGC9nFerFM2HQ9
9QCrzUxO7hJYP8ConMpzGkwC1fbgtID52r7oKpxS3f6j0pvLA6rogUOGNl4Rfm+u
2oloML9aQt73Z0C1w1UxkewgMN5kY2pl5eniAZvP0VBcB1KjFKYWJnBhDWMzZA5e
YJJWGtj9Wjr85/qDLkXzY237UpvhAxwzBjF+mGKTug2yp19LhV4WaCyptiAoauD4
iHpGGX2yX+I0dNNL/+5TWgo/4x2qZEWLMJsJEfhu9JU2I8Nl6faWvgZl5jj5ZTzh
TD5hPSSVGPdni6F5XweOlGI8pkUDLX4TTXDQlTTNlbajReiBNwrdP/bPALlhDkqX
bcBk/zYk/Yhl0SZBjdlYzfx7Uf0ooPOi+Ol3KxJQ1gVOCtokRFgGSiPIgFkqAiYq
1DcsbK4qA0/N+z/Qr1NqBZ0CXW5qICumB8uvNiI4QMk3TuOqTrwt5cenfTnOk92h
zSMh7+RhuIdFlexA3+4fw6CvxH0ID5HV3hzXfd9fieAK2WLBk7815k+ugWrAgDtN
AsiB3B2aOPjwx3xBVIYqCFUmM/c8VXbi8ic3j5C5/ec4JUlG9SpvXmHpKvmekC6q
tSHMyR1F3VXGRRFqnl4v3rUBUXI5+p+flhkqKg9U43jtblJo66r2UWgcIKfPMkRo
gLf/zlILhjGMEef3YBQEdiBxQRa7hqexpxWjNn12K5Alz1FasRG3yHdKkkycfp4S
n7u7kyOxvp/pOcp3pG9rJGi/efmvsn8F6DryU+FtTe9vMB5p4KGgxldDpEMPvdSM
cXFVROjXk/DwJvKaPcGVUmC3TLQDzs2KIpyyV7DP4WCpGre20X364qM6E9KHIHSc
RhKwM2+Iv5/P1xgNok+L7PzyF7jWS1Rr2ZZ/m7S5ytNaEoTlyDxshMfe2uIb2uqn
vJYHDiKEXIXycfEwIUktm7y6ATadd4pgLe5EC7n0wA6OM6pUDwpZ6dxtLlQ3fDYl
S42mdlzdjjySLQ3vDTAdJrstikxI3ixYVNy3hDF565Qrvx7F/oU7Yd1A/uCxVrrQ
9zkeTA4QF5wiedyIwZL1yIYL8FJvRMFZooqVXsWH58Q9alZGd87HG44nxWXT+EDJ
33SOS0yQdwnl/CbpBddH9X/Iyiv3DF+5G3NOKmQKI1QrvrE6HOQqZoFKLNYlQiR/
7bGmgcy1s4Qx+mR4cIGPwG7sQM653x7jQXM0DvbxdXRKPyCfrSeVJB0L0gFdz2Rn
BSmRiIEKSUxg/XsIonafZiRbRaCBQ3ZIod9DxWjnfRH7OF3s5hpw1e40Q9KT0EYu
1/wq5rKROOUs8jjU7gBapD2whmvetky2jcMFpE23TNKAkH8F8fEwfCoIKaCw3iDs
fUjloJUJ5GTxIYqxhaFevM1mQOifY+7ym/0UE/bl/fdcERfP8sBgYImWqTHozdAB
AYNTbRHE7M2XMuwnql1/13+6F/Zu/JebyNarQfQGLEs+JT6aKRzZI7eidAP8W7dA
OVMpUDNFT2Xs20SFS/pZzCb4SoLDDNF9EfbhES0aMMPa28vekukcQnrJ88qu9YuO
IZnONbWb+WhyrSJc9RF8w/chPau1hud/Bz+InvuPyLh88ux+/v1JViTk1a9NhU7R
QGI7nWMjJGUt+HoG9UYu4BiZ2OUZBFKtE1KuH/QeBoUjWRcKdx/9+8k3CnI5tCIk
SLEwDL65cu1Uvat5R6DnY5Hyevovcxbe6ScKzBxEqnhgkQYjrHpPb+BMe8LRVx62
+fKR19U+Re9O5pfpUbR6Zeww+/Am2kUDPlicxEO1mroqEv3/f4uoWWYz5sJ4NLa/
ksQqyX8e2CFWyCi5QEQvfsgsKNYgwlP6xXIsGoOcwr3YsnZn9oxGrWSf8fUE3y9P
IPV0q0Fh1+zcmMF/+Cb/4hN3Y/z3yjgZtVbCLZ+GytUNMKItleGYySXO/x4hPqbz
y0CNC0QTNCq+3TyEOrMSdiJaq1woyfaKjjBlTXg8vv9F7TLWekYCCH5mu8ahdm16
R9IYh9buLVxq94fFULKr8GqoF91E00XHyMuagYCO9Gz3GLSMVbhbHJeBWLB2TaYa
ffuklguon1Pf8Gu47Q6dQPGuGlb39V1AbznnYjeIYE4yID2aTQFgeyBoiNM+bjoI
bEN5uSwLW7JQv5t4ZCwHX+B9lWR2ESyCyUrt7mVNFm57TsC2y5g50+ZbsDPofRQQ
LkHeDlxX9b42kUO2y0i7TKjn4TVlXBXWp7Yqk92lvN86JtqKgkiSZO8kUmvAu4dt
0nFMfjLfC1kyHnZUdAZrY+1PymP5LmnTVX69eBisoOL0A3AxBcNbNFcZ+yAcg8zb
O0ZgdgnFIYkvzdLczUl0d3fz+gh94Pk6drkgt4urc+41t1GAxZFZRwgYsU91PbgD
Ri/vtZIkIVN93+nVYr0G1hdSwiRntT8qejGYWx2BKEYkQPK22+HUesCDVhthd6Pu
6kOERE++DibmKNPDJgGJTxw2GvX6gHNalasiDthZEVGfMmJtwwgL0bcfaTFtJQj2
AY2b9AtT8U/MGzJoymE8EO2YYnwjdCbJpwE9GsFBR17Ed+hxh9ytrNvkyfleDLAb
Y2lRWtrFcKLfoaHCHf4Br/WNIoAe2VCi1OXzHiJBPvM4S1Fv5UwgyoNeaQSJMz7D
kgp2h9wQBDiJ+s7ZYcmNi4L8y+51HO3POTXt7bcZoGHafMym04fih2W87hMQMYIi
zIIN/zgpshm1RVOmGm5m38dKtz8RYNg+kVprMOWb70VLeJpj1QadeR3hPlVCHgZD
asSVP+NSZIJSCKmV0ZQ+6qAqCvbXjdYC9d1xdV4R4s8LKAOVPH9PwM6MWErmkuqh
voVZWnOV+iv1jZ9RmC/45UlmphY3XYLlfAypIaBh+56t+rbGzsRmqPoYIfp20ta/
WQ8isTGsCoRi6vhs2Jk9lvx2cz9FFljjkQeAVt/VGZUfqk7k7uZog7aYv11RMZSC
g1Rq+eLb3cCRMy5eQSCyveaGPWIJIL2C/y2Iplh3P/w5aw6EttLwABG392bKs/t1
q2B83D4PJkcNCzSRHeqfbkKhyma4xuTiZt3bvmRsBBJD0+IB7yU2OeIx70IeBv1j
Su6fh+yZ9ifio7OFPz1OdeslbM3MOYQsDveR1vUVuKjGYZZGU4oWLXcRdw0d/Rw7
FB5d4hMDkBZy8VFup54nalE+cDksjxMjb4A0XOAr2cz+1DkE5j6Q2Tj3Mvs70P5v
SorTYoA3+j+PdS0TORRG4UwtEq+DBdazibYmQwcg3jm4ouNEaDJ54gSnKj+wWZSy
kMiSiVkWs71snFv/CzoyNx3ULz97fpHDFONZIQ4B4HF48etyxsrjgPwuEPAAuA2D
BChF9oyirSEqggrfZ92mFo8JwIXFeoGojYuBC6gKrqpuPv6bPySzebUyZkwe/w2f
JufadTher9IHMEPLv30SqFlo7BQLXIZpY+QYTxE6Fa9U3/SskCzKTmZsYWtwtihC
kJyu8m+Ir0tajr914fGuOVZXVPdFBhwRG1GXqfzOONo034wjEjD+SwtYOgeFhZXI
hzVm0B/cnA7Z3/V61d87ofQJhxGl4rq1CqDoTnixeURiViS7Zj8CFAzzmiKG+wtK
kmhXcjrG+p7n8oI6Sc6gj+D30E9Ic5jOSY4/h0hebdtbuWrMfmW/5BhWkUBEqRJs
2tgACXNQ5ZaKLzWF0TXjh2FEMadtJRZNi/8TBEjf7UhYceMkpyjj0I4kZ4r1FjUz
aR+PjgqIEhVOQyyQMEwzStIyBRMpttHlZmpcX8h43IgX9DK7aq3shKu9FYW2/h4p
5zyO0rh2qJmcIOdOehhlPIYRlFFollSDdgThE/pn1mYUYZ8JgCXKeVn4IGOjchc3
JunbsDgMbQ1abcmWxc+YE98FBlqsdiWT14n9ZYY7vaUrM80Wp8T0WSdgBeNbvA8b
OAOvUzf4HYJ7Gk0xjXf0vCdh6BQjAYiJd9ZT85cxgbnpgItZvDY6R9x5n3LLJe9J
Y6ZIGl34dSIM+BiKjLodS/zk4SL+4oegLwpdr01BJfSUvTmCuj22TGXSwbPPrwXi
eFJAXx+s6puyq1MJwkon5V55d/SrKteamBSXET2M3czVpQqUTCjzx9bHMaB9++hX
R1kiWjMTn3B00mjPEV6/CDEjvk8uLMxbGjIKU7R+3v4Aeyc7fV3zgEW7iG+Ob/Fo
FtyFNrs6lAodQaegGwt5qEOOP52l6MW+y/xJX1+QcIpCdfGgvvuQZmFqw8keioFz
9HS4bKI7zzeX3TXI3AJ6vvJehD5JGD+CAH59/5yj7EQVTBvUP09T4tlV0rGOUHiT
Rg/GOBNzMbJoUlqDaMLUJqA1Wl6Sy0F8qBg5wAy9goPOPPC2IxWmacLeWzM2/Dih
pjONQclgS9VmSJVGQ9Flq9jZs+miRZPS9fYT4pl0jogjTiN3ET5PmKg7EYH6YwMP
RwZ0wyhrBOtEDhYN9KF46RAvVxXg/2fjSRMg+EWr1YXz1+6T+Gdc71NkwB8v3YpZ
qsBaiJj8PnTowS4vf9xONtgvBPTCx2mCGMLsWGd0aKNxkv01PSeRcP2k5Zf0KGoY
yI2cnOXQQeTQZcG00lKCrjC9gtmIijxaZHwsM5p3XlcQK2ECdT7L+MHiq9bMFyX0
eOHJ4qLuhFbXy2qg5s1ssoBnPBhaavKFg+ogYp5b0I1n+F3YH3ixXloaX2nOnusy
lwFUW/kPdq7i345/lmFwcvlQwrNva9SnG93iF9j+c/ZDORu5Pj42W7ADZTY+ULXM
cDy2iKvoc14W72qe7NEvhSC943d+TIWAwzOjZw1jWuOm+ebMoBtyYGR/asbc3VGr
PEdF4QwTQO7IUpYM7qVpgEFyUkO803NqzW6864GBUBNUTz0+AzHx4GlgOmFQocNa
8cq5/RjuZzGnFPY7yl+NhGtpEPrgnUOaLQFKPOc7Rbd2Ai6Ukg+1wcC+/bgq/kgi
RD6cAYRLVmchcc3RtoWjXPbs/hd+3weFXlcxVQfyPlUvPbCm6VlCegoa7GCSCerW
LM4c6EJYYNCtyiL+sj/2kJWLOUBZcvD4nk8xK8/KOhmmtfOPzsq2gA5IgUr/2QCM
0ZYcWrLQKrcgUcyOOJ+8rHJTzdeHDrcPjmdhBnfpS4nBgLkpV0f4dQRqWMSGtrhT
7nNttcrhVb5z9+gKJvWOOc90zPdYa9DJvDCYEqhoErmUs4krkhGVllZtVCdk8QmF
w1puG3aU7VTf1XZbGL6lnEwDVMzBZ1zJlnqmPHD9ZGoplDnoQrQA33mGwEUZL4XE
lfgADKs2RDzCHv90yGtKwl5oyKRcUq58dHKu7s2vlV7dg3MBFinaT1JyMCj0KzCr
9PyakOwIIOZstTClJlw6H2iTzjj29jqOBp7kQqqFtYTxUf1n2sDM09qN7IktzICk
OeiLcbh4K5sGFksuj8hlNRCuqGjmkSNMPeVnA+/8zxaXuWcT32psbl0OK+9KvZ1q
Rl5asVsvHeCublXKw/r0X8fQSksP5g409lw7EP/WZWUxwdc64NJDCYUI0mznNz5s
qgUvqaf/HpmogIrSWd+NrmYLNkeA0gifWxWtIT1Nijw+cdyayekcMnvjaINqdDsu
EhzwGKTI/El55lTQybYBAVtvmNfZzCGZkYVXlycyRsqiXgplUhX/4A4rd0aDhp0N
gNEskmSWfqH3ogbUQQKlS10wXsF0vXzWikf0DF0XpusY891tngnjnFBQWHmLhZ/B
dQ0D515PW2eesq2bplS6ebInhsAtkxnMIrNjHDx/1LNdrDRzezSfoPSqEn2UQBR5
Ury1kwqQ07QXMUNCvmyEsfJh4JvQwEVS/GLkkLYDQfUxxPEqUl3BuuVSxeFC5YKU
6DkP8kza0HyZqKsmOmVE3zHa4VaKSZ+XGKFtZHAqZPfv7Gq4y+4nB2fYH3oKuQZd
Ci1CY4AHkPjgg/luGDipajpceas9/abilF/n6NofIuI8cHXnu5cDGDx3YQoETJzZ
KTjj/ROY9UOo4cL6x1RRjeQnDBiQnNAELxXWDw7WldaiVdVa5hTiAd+aMdN/j1Ha
bovGFTiCi7xlqx/qf/mr0olvtvZldeYnEa3K12Jpx4kamNz86fcRaWho5ft8Bh+5
D2MB47qyzMJugiB226GPhi0QrOKcxoQZncsyoHBPwqQGtAgaw/esDgf5RERN9ev3
exWdxE+ysno7ihvepPgM94k6nW0ZAKzb87nKzixziz831yzp/hec7k3BjENCJyVQ
2z+mUjGaUjbXIHnX5/B2Lf2m3Dc9B6yjkaQ8tMDolajkwXL58rUxegXDy0/74HHU
a8Ovf3Mi+eifRcAkvQ3BNt/GtQWoVV1RXLyqAUJCuRSzfxq/uJGhrZxc9CPGcO2i
n/cqW36pU7Gx9Ocf7jfvz0c1yX+reP8dFvYNRJdiHdTaMHx6wrABxNXK4pzE5XhP
xowvkit94nBgSl3NU6XNymAhdghHAfRV2qjfPlTelx5kPSdqKJwQZ4xQTGaIXGwF
znKCGDd+XQ5CjWN0TH+/GF89ii8qRtIn3NiQYfFeAIRyjtz2QQWrn1HFleMuo4qW
V6gM4frOCwQxjJPOKsrs9PrnhDZKCVDcBXdITmmXnvMkV3glg4xkJevXqJkeq1gJ
5dsB7MBFIVtwe6alDgf5nP7X1/OpsvZjQS4k1uEV0PL5zGnpIcpMKXMeCSRaU3CL
+PLidvzDlq3bDUjM7G+Fw6QRx9z/zKiZfKrtimh70LoS33ew+uPqD/HY7Unu4L3X
fkBkKDgn/V0IoMbuiJftSv2UFaliLKQHvqsbHfOYdr4r0unmBIOaMTlxzb2MloDQ
162gaaBFHqghaEMxBLHsRPo3R+wo6cgWvMe8zGBVZ7GvjEssEzTlXUbE8eBd7/Pu
q0Ud3+qbWtXucLqEqq5ZVFCwHuwzmTWkJmV78erI9N3Py7AXKbSL5yvRo/sNUhKR
PJ2Md2ekys5H+6LOlOhkY62XO/lF3LaewgYhoFFo2LHTzIFL4HfbMbKnr2f3VK/4
evR8Hy8zHf5ah5zXFsc2FNGI1Lt044FClAf4i+5uojiE7Y0h0GYCEoEV/Z9ykYzD
zTLtcP3dwMqX73reeI4ix5rEc5XEt7jAyYafBKJXRm2Vb8Cg9KvWbOIMYGRMZ47n
keRqm5OteOvLsIrYS7XctKvI/m/X7BYCbEh8M5K6uP+XwRYB/jiu64tYsfqncdoH
RIyzQVBfyyt80Rz6eHYXiqXc/p0p4b2O70f0wE1tqC8dsMbH55B+TVPbCQaXZrii
tp9zWuPaovFf8Au3QMfa1ISgcrIoc5bCz0ghLbJxnboyX9W674BUEfltIbgnfT0X
elOeD1lnhybYxNhx3I/FVrEjYHw8eu2UiajVD++lfvo7bO/O9aZYRv5GXUVxa3AX
6J7h2wZiMdF+uplfFpdiyuwZvbnxRtdsg4307xPc4bAfIkx+PKluTeiz2uxaChPJ
Yi+Kklxcb0r77+30eC9304S5KQGflOAfCNCPySsPPzUseA913BuF0cvvQwPkdnea
2PcmpfWEmNZEWG4f2+v8mOmtD2ugGKz3g/rhL555BLOpR1ifwQZKZmAIzB1IV/9D
zQ0i4hq31Df4beaUUWZ/lCeZo3uOnWZfVaU1H9GIBZ3ufZt9pKGv/aJHkTCc9LJX
pt5cmdKlhiDVt24xtMqX2yVnOX6LX2yeI625w/ejhu2IMkn4w0VTOl2C7t8LQphV
QIOYPtDpLiVjro387QS36pBW0JFg+eMg9Lyx/y94HEMNRPNEfN+kkalXdK1d0GOh
EbRZ0f9IuVJoPej2XLncaPP4yEXJ45yUk/NKVKpQb+IKt4nG+6cN/dvRxSuvSGd/
3YnVC41Dam1OvcmqBhPC/KdT1+GLTkhxCwvjZ3TGXO2NDLsK35yZqLU1iqMeDqdv
tg31xr3/mRZ2CYcLPepaYcW3tvySE875oNRs6S6BoRS4hw6cGqlyC8+PzPVDhp4W
FIJEVwrRAFvDkBEj7KvDZaeDKsG2XBWeqyali5m6gpXn6waTlCh3nnyxfKA8b36X
YWFMM1Uelppa4ceDWlsQ7583Vw9I3iIfgRND8/RQIcjLXxcc4uRGGNnhaKJ2P2MX
XzK91eenN108sfmEBx1xFG3nSnDGqITWwM9XF7WahjDeZBlnXkJ0mKJrrWvurmML
sG3WI4BeEVfzm6ZDIZM5YU67e83xe77wqliEDcjUpyVY0KUrbLW99QHIZiGmgGLK
Z7a1jrZn/yUiRElA1ohPgZ1o5F3TFK/F4HewDZPSjXGGQl73g6xq/SjHNfLJSWXy
2yYOWSe9awfLzZdPVlP4Z/qblHesAyaWFzqNhZsr4OYvK48I/tlm4AYNZJBLRyZK
ZWcrO+TMO+ryyP6eBMO+EyO8uDN/YqwR7TnDNPG10bc57IB/cmiQtWl4vQTwPeFF
wkSboMSmWgQ4QKQKOLhPB2usAPxCmz46l9Ejg654KWKoYx9JAvrDUHLBwllpoTCH
BqaQ0b5BFLFELa5JLnL8ZPURPbR/YlLWt5EtPD05uhSbEzcfBrw8qlk45ZWKnbfE
/NEjjfQfvRssKT+eciN9w7IK4bGS7QLCdjWucwpanaSmtvyaUFRYgfA95k6WKybx
lbmOMbiWR1cDYOPMjIXie7KTdgx0DHnUjjiV02y9el6YsUylXlInqOAFZnpmSsh7
K7n1KfNIbRXe0k989eupBA8Z9Uw5mArHru4NMbUj8iMiQQh/cQj7hWy6oRk3J65F
0DMnxZY83J0qcAcOgXMsDbQQgEWnnJtsFPYlbOOm0Px9wxhWfQd4GdIfpCh6xyIw
jBC98gWo6/e69y6+ARuSo4Vwd1O21s6BN2QB8GxRyXQnvrq46uZrnWwv5P2iLhPO
k7ma1AaAiGdnM2YNBS6b525Ys//6J1DabaxLdhyb6nOuXzGkPo+NiNINPx3Wt/7F
+9JUysBrXSlhZb/cOiM0n7lvGqedSNrCemU2aO+TIRYk+GGqU09Tq5qCZnhGgbr0
JvR1hLrcHMHs1x1FiTH3OdFVlC1572tus+9mSyuh8yKacGqSQQUdRhOQCYFdCBud
tEys5Jnvo9PPJXuYA54Cd62+rzyHANhH0KebGTfvDIzdrEz7HMMcxcRbDXHbM7aD
hiTU45cq7EbTbFmhM+GNyf86c5YqeZ6/10Yjh+gp+EpSz3sltWqNIAR52wUCLNS/
3dkbzc7fzixk6m4ougv8DiusHf6vnYneKTERJSLC8btDdnyU/Rlq5Mll1clonF/G
KtLGy+P5luvG23n6CTZ3jjzNYQCEofbQwGt1hrOlctCCdWAcDqoYqflyImZtXQ0W
pu6LJdp0QZBbRZQMp0rvGux3VR+yqgrLPZHbzf6IkmU5A9PxVby/2xysSV/T4F+k
QwiNbNmwY/64NavPD7B2OO8nQedVMuoeXHajE4jnkBQa5SHOsX+nefo+lXZR5Voa
LX0MHj14NQEnuecSdQv4adRa24OGP3ZkZJJ2Uuq8cC1QF2IgVHdknyskjVCCs+aR
bPyRn/EGEkv/fNv+i4FvUy1CsDxdGkzQJoQMYrjJUqqcwoVAMB44J3lDIkXcXCFr
Z4QAh0RzBMudImsNu3wVkto/Rnzki5kUalTmUZmf10gejmwyiwKcjWqdWylH2ZG2
OcI+AIfu6E78SEfq0SVGbgy4wNe/sRDakVHgX8+nzzNNusfx0fPj43x40FF+x8Iq
TqS+IwrekBnimMjOMtYhkUzRBHBdi5Bt2qBknymJxiVvHYaPL6+YhGrfSUqMvEFT
zg1w1K7jkwuUUWihEaZB6iAIplDkj9TYmsbf3xKv6xV94kYIlVBQoK2d8Byp/NAR
UN/EhYgyCAxy3opIIKNLWY6KqFyRzrVImPDNLjYY12DwBsIlhWYH5ExC5dWxNdtB
J5TmdBeWT9Mt93pMVi2dGwi9QuaAUD76bVbOQmjbmnx8Dkd3Q+xSUMriff9i2mm0
UGumOlvAFVwrzpIRRu4Ty2hw4RTmgBdrZDRiIuujsRzZ9FbHgduOCmOMiP22pbHD
Ji7hhmcn4y0Rf0dvgzybeoYg1r0CQPW3xA0B0s1N1nu69MsIi6tCentZCn4BUrzz
up7mCJCinxGtSsNHFt1om7ii06173nUze4bRvqMkfRio1PPDmxwgp7/HlhTa2nVv
Q/D3ZwQEd+C8G9A06Vakt8xz2RyzOjJUR7+UtyHM84DTiB06hNjsCpdtL0mr2/1t
fzMIPNIhM9NAkV2auR4V+e6vW8XQea1595MhAN/VAPedKfrVHFelNvo3vpZorkyT
ZdwCggpeuzMxVhAgKsH73GO8oC6FrRBkTKsadHdtQTmQQszsTySEqtRBL+atYOxh
nsJWY0Gs1AAS8io+hCA7miCUXumuNIVpqxGvZf88fMLhdtzggv5rr3TC9rCrx5w2
xLLil6vDlcQQZGflLW+yIh6YLoVF/98NqwT67RTzJYSDtaj/Nl8G/z2HpEbP07td
scqib/qYhu3Jk/GceR2ggy7Jcq5bGbwze+q1ku6m7fqcfFASmubYDYNQsiqo6Cxb
qu1yybrgct8xvjUK//Co9a82cSWpVbE2TYcr4hN+3+jZKu5hwAffQPSyKRRLSC+Z
z6Ou6zCR5YRfHqKKMo4E5QjSFvP1uw0XEQDNyNLS6aFyPVaFvVfA079xcNCLDj/Z
CLJS74r6A7dXHr60KO/wFauo0YmFZvznJig/U0c7XNYRwZGYZqPo0fHNNHr0jJXx
fAHwb1hPJ7HCuPcNgl5EtCg/DpP1a8qhLXUVwmKu83SbAIKz3ECOCG2AeYw+SqUE
WbrtyZPW1cQJvnLozp9AAoVw2rdrDh/lZqD5glDPd3MiVktkNJ5yD4AH37G19hQG
yUVDlWI8KtaxX51aa0+jPvEVmF8K8FwwGTTLLx+BhBhLhIR5q+zFlPhMGDxFp4TR
3VHSN/LmAQD0w1KhnuAFO5cLN0v+h0kpK9rMlIsrye7TtLovO0Pf36MIxqcptL/J
+h0HobAm1K+9yhqLvCesktOWaxeVJ1tgaoo3LnOm5cm29Dr2Adpb+9nzGmZraUsV
5U82Z8OylR/dx08Jy1QPXAWq8Ax8/YNsvFWoILbx2F/TmG/2gOcG5sWZboWOQP/+
jmXoRZptkOHRoS3UD1kxc6O/Kw5QydnGZzNXNPxkJMt6k7hx0TGpBPcrDCGx8mBE
RAyU4zTdCZaZgjDZv6zQ5iKkGg2TLDS9wfQmgUtGYHluhXLlYOeabZbSB55mIpWB
emRA/X9Zyf+gWD8Vv4/2ryIICnFf8Obc9MOeNdfd4j+WBxZ3OQ7lOw9zAnuyZFge
mheSUaqdQ7jso7Yz6XzQQdfSU7ihqWTgAGTjEfwwoMOaloyJex0LP1qVhoN8MgQk
WWqkcVK8j+976xoGijS0//uhdLTBVpTbaT23OLE4iDp252ypGLutF7pky7gIaGnP
8BrUiu39lPPRnDPN35JMXkCJlpkHxy4RMISIRhbmNcFK9eGumQH2WzXW7fYHKUbc
VJfNon8p+HiLkvmL73CuhP06E2VTH6cxCmU34qEtUUjUVu3IjcOL+tWjBJZi1+Jl
sCOTARoasevkyW0PgUoMVC/c7SbmmdIPQeYvyA9oomJrRl4CRIoP5X6ReKFn0/bC
MknvQLruu3X8AhMrBvUBfMMmCVGqCChWj8LDX6MtkGkIEUBeSjvHsWfdD0gfPwvq
XHgsYduIW3Nsd+wLfnImlz9Hnucs2jGGCtKBYJMOBWHGh42hrtnvsyuPBMY5W143
zqGqYRcQ6OXrQOG8tCcdjjUDEXXg8KaH5g4r+e/H+uK+iTN7jDKlFAWaHoaE7PfY
iEVUHRb60ZQ42vGHzBqSV5pxMxH456YMv0ktkPtCie1kjd3Mx8hgHoPshYQgrdFQ
pbtMCEkzhXdxHjo59syXRRLRdKrixAZMrDSK5tZOQK0aXrAsIxRxY3CKEpWdxrUP
kkMm7ZURt9nkXqr06QrI94J6Pv205X1WBn2svKT5lTJJqPXhYaK5Ayi4VqS0YyV2
UANad7UerZiBJDEb19iQAeeUWfwwkB1Jc0PuZD+40pmfqeDa+Yxg7y3KYnhftMp1
sgb/RQRMqgaZMF2mvG2o5xcxQAyCQi0zMUXsmyE470+l1hmvALtdGJ3UEg6fjGXq
pIjhpr84wVoiK7ZzzfH9xC+W3a1x1nWzri8XIoQ2x2M9pYSxmx7VqbcAR/5XFjgf
9RdGtH5lS85d26E5vW8Fu9gr6c3QPwRyDoJ9olT0rYDJvLYlwyXBS3ptHl5tpFRI
+1ufNUi9IvJPMTTIlYd1TKHxUHXR8h978jAfdP+zHji5wq9vxuqfWpUqfHSDcZGp
9lMuhx/sthSc9RUseqfpFJTJqUTdgC0/UxbMsXSfJI196Fpe91XKS6Rv5oj4cD7i
g29wZeR2dsvfvVwb+lt6nV+jHM4EbvqXLfBvQK9KmSbaFy/4+ODcR7ctM5g3iOTT
cAbHGgjXsKHtcld5ef3YyWsK47dY0DSurLM23JgStEw6fW9tmPg0koaSJ0fo+Bcn
T66w47k6vafUJtn0o+zqVFCn4YmRkh7afZLXed17PMs3q6CMdIgZ/ucDTDfs5L5h
AvfWwP3/RgV5qdZJLAZZE9v1aFZ+cYjDEIsBc6lyl/dUt62D1Eg+yTxC/6zAnHTp
zgctMe4hINk//PnSib+rUmiOMzBf9XmAQ5dva4dDbF0zJXffT1d+uY8lha9hkoRU
fvPgavPwnVtDAQqPeD0CTRjYGH0QximLK9rhvc07DEPDhduEAZnAL4Z+mF1J9WMH
zDHaukEcenl2Ga4q4ax5F60hyFINa9eMUNCbnsfPO966Dn8gWSXSOHNQ0TrHtits
R5vIBdEX9+fh4tTjuK0dSAXplJlozIcUb3x34dE+bH36sJxu/Jrvr5cUkJ2dpCxb
DfVSTRuAahF7XYDKlTXPW8plF7vGSqsYn1fvSABScURn5TLUcmdHbV4exd4sdKl8
tJTz5Ru2CfN+nGyqCh1Jja/5bVGHpCmsif7hbr0WK4tk/fatbCXR9tvrL/Y5UGJN
GiTNqEB/AFxBLwPSWuAsWd6WbNzU7sKqciiytstSd7EKR+NWBMgBvModEMPU4oj5
X9yHdRjtlqXSmKc8JDjtEiRQxZx+iYcLSwkYe5Go4mW5uHYtbart455w3r2XRzQi
8BRr63dNjmIdyh6eaMz46YjqJnVDMEqOiHKGMLYwp9kd+vO40fzqtg8JTAE1u2sB
ueH+FxAVejCX52hmnFEPLjNuA8NHLC5954aViX5sD4rOi4ry+7fmGDKx3zQbQjKl
0CHW//Hr3R39Hq2D1aRYk5QCTpYSmFA2mwVVSjrdVwt05EdXbRxgxp99z6YI+6Pg
+ffiDn2rdkARCWLzIPVIHcBCbV8riEoqc/LkT0giAmpO/8vKLEvnUAnHAxcnXsN+
GOsAn1Hq99V+PfVoY5PWSmfgzZzU0CB2k6ww/zUgfbK/HuCxeyJ7JCwXPr3OS0ES
MsvUma8XYYU6WvKunB5UWnRK28veQgCr/IUA6O2hsWMdLyRN52aFqNKqUzUNwOFI
8WBk3HPxk3HDwJsk7meK97euqPCGGzWB/MTUR516+AtcWr4UEA83LITKRxUw0rq2
HdWNcppFVeiRPaoDTryinQE2A/Jtm0GWLmz9N4RU786pO2hUxUezEpwwgtBLXI9x
Bu4Md2BhRTjHPQRLuDs7rHvMtfcdLlZxZiP73mwd9atPoo2mmli8iWv3v6M9Ggib
uUnsMd/tzs/Ta6lEGCL+dJM3ql/ch/x5Z7fdrPIe/6YKjGPVO/vy4jjnnL8TlCbw
v3hHISeKnn35a8vwQeAYCTqj7SHJPoRrHXplsA1KiAC3WF9+sYtnsFYLZVdZt/xm
V5t3b7S6d4WotO+nuag+qMCsK7Uk0UItrN1JE6bExi7rnSDAYoRlQSNh5NDuWFtI
u7CZ0BT81/RsLPbJrHnEep7Rd0L0Xgo5dd1DOZE2PUyCU6xsNyBEXKI1fjdH7skQ
dGQijZgHa9siSD4cC7yF87K9FRenTwLDkYgsaGJ9X4+50DhmXemg/YcXZWNw5fLX
ScZCWcwSMwozDH6M1sqmv8oshaZvqZYXHYeQuhwBPcpA85D5RDbfOQa3UMak7PIX
lOmwEHF33DpUn+sxwvYUnUWeMpbndhCuhDOzEQkYeexT4oQGP6MRrDRNqll7ApAc
E7O1lsNifcuUk3oFZuvkA0JIbqEYYKo0/NWHpUBnTSEP4gxW2Bo4x9mIoiAgOXMa
BRgGyau1z4k5AIC0adNkUdjJiFYZ3ePo9Bz+9r/tosVnQErmdHHbwT8YPMPg7yCI
EkDZVwkfWGf5URUTS8gpRFMw11Ed1FEd4Inj2UA9SvPc33tqgu67AJxOJEsH2+MF
3U/ZzyvwgSTUBqT3Ogzbr6b8vIXpGUjHdJw3Z0257575b5oxZLlA5ckrV3hA7UzA
ecev4tVaAHB8I9ziDLzKlmnM4vZYEpXK0eMmSmzIaVN04HP0N/4zAn5Rnavxh3Bq
GdPkLnXa1EynPPXd/Zp9gsFZI0VwZ2XsgoQQy6jdusJ0jAVyC1rny/4IVpWbdzdm
KQylhArs7gVeVzCMTzwIyPIkye2T4FWjwzDDreeBeBnKAJmbcuGVkCQ+65UrW/EJ
kYVRfYCL/QsyQymc5gsI71GthWBvomqJjhLifsDsFx2zqEQbQyReZs5IZfCNoD9K
dXTkFuMZvA5RT5zDzNr3niXWTN5bVBDdzLoLSNA/AMep9UNi26c7pYlcNrBTtIi2
l7Cj5h8mJ0lVm006Vfcn0jspGl/iHYjI4mBnxckDbFCF0g5PZ3V8eKTlV66T+Zfx
XLebiqPexXTYsQTMp9O1bbeWl9xMkBp6+9Fq3p10iTDeX3JeSF6zPkjOgyhM1Xb1
/L7KSm4sPImkQf5JqOEV4Gi63fcvf+8cdLAv+9G7HTzn3oO7UFy31gCJSCMGrvaD
0qn7RlvyXj4J7YKX6iOTraUX1sK1zlXUrRFWTLVbHrXEsyewnGdlw3j4tuEQhYph
Df/LDP0vhvGSogkZGZw1hqxft6zfV2bCsAFtHWEwvlIFQKi0iiOEqNLylcL65ikI
64FF9cQcsa4zAwF4DeRw1DDKv6FN18knbbUeRRbQPsWZ92MDYMfqteKtqFM1BUat
e08cGbqjtW3Vnqr79ntArbQxYAR7tRdpSAIdzOUo+6dhH2d8wvSHoKwv8yzSift7
YC06IMSHYZ3xmQSPz+o2xTb+H6xMfxCBguY4kJbpcVfOjMCoz66BJBHyeY8BWiEl
WMTN+f5sibjafGKqk8UCD2P3WjbViSjzsIQSQFTRNbh5npYhAciCPrnJnYcI33lG
atTKnrKRyoIsRtILfT9Qhabp3WoWUaK63Gi7c6M/amONPHjQ+c6sEwtW2R1IRGDa
oiPpmb+hYjmuSYSaJ/Ow28FPCLeE0135NNFYD4C2aTqrj9rpOFtxa1Cz09V9+RMM
+Uvf9s2Y7vXT/rlWYbyB7FOmpgUdLq89IqhmnmpmaMI9jnqdLxrnAqTRoLkOn01o
uYw1/a5kuTyzDVLktjMO00fDF67eJqvI+O6RJvpHPqA0UGqaJMy/+0x/ji37uKeQ
deex2lAew0GP7ttPC0MtGCrTcLolCEbH2nISEsO9Ccz0PcmY2QiHoxFXcVziAdlI
/8oO/jLpuXiFm0waDBGH0wHo2n0LNLGiwhA9P/BoMl1iBjSdoFeyJBFfjE3nJdPU
1tDnRi7ZIgLiyq3s9tyxGhpp7WOfBwNcY3a32oGuMozfGBgsc7EZj8FHOdjMIpzI
KqqRJO0q04+fSdOtRaSfHLDFxtQ+Wor1uDNcNzZP8MO6Z52Bf/yk8g86V+alrqUX
V6o3uc/NwBMAYCAG2ohEL2u3ItyplMevLMRPEzmkUCZWzI2vD1mfR5ga8DlxV3V3
r/nTir1mVyovv//pu4y8oxHYL4+1JMITA8uyLcm82CjuK2h4OX9cdw1TUU6wn09t
Smv0DK3+lE497Lm/S2ST8dYwVbg64ZyEJtfhJqH4PJBtzI4DwWX1oLniP5+5glKD
mKDndsnKovWAn0I2ap+LyGCt1ciK7BTesdo3p15sNP6xqPZs6wc1hkDjRShltH2E
sDXWMlNOHp10i6Xm+FD8L1p6oB835jYqqcPbSfSfI5XPZtKh7Qt2Sk3A5/lMKGue
iaN/jAUXcmuJaFiLR/gwWAchRn49V8fhNuPAezvcbkKLJfid5buYdh2LHS4Hqf3/
MIjbS3jRiwJi/PnX7gydojNgd+L7pyAJsjFoLMhJxTr0iP2dBAURsahOY5Ya5K6G
NiM1oBOhApTZMPElLRgSEr9GpOPIlr03EW138wGUyrXUQiI7ov3Ct6ACTG5Su2P0
oclvyrauyFqSCiwyi76xtrzNL4WU9NK9TI73VsNoQjcPytLsXItvPDn//y3y3XPk
2bZtbdtLK/dG/C1yIEayppMkcsj/DlyUF2QJPUYVvm0CcLSOHKz9/hAJd/sQQfiF
BJFuVu6Sl7M57k4HzgWgjDPT4M1x0JiY4H8RFgY2TlR1VV94XdpcRXKetsmm4MuZ
N1eqezBSu1FAYUOb3t5wPeSbE1XLPzZXAV2Du1tYHLnivosFfC7WI1yAVgfKcVbN
iLgIIm1Vs9z7wNQ76J+cm0WToANYmJctHWsxCsgcwxoBc8swwpX5IXq/R3zs2dIR
IEdj/g+6OwlBtw1lkhdia3PbqnkskA6fhFnyDp1in0Zu6TSYLeVz5HsWPLFE2BCT
sM9PcwjiN2fzuAxCC3dg0SXC/SYU2qsMMFgKTPvEU7dXPAsvechNsCWLuXPwZ/Fd
6hvlB5yo8TB5OEQ0eCTpmTnmEEfIELUru8jUhatZ2EY3G9YCmiUpUoqo49Pnd6nU
kXGeJBkDY0OukYBEv57qV0FjhdynUYpAtbTAHJlo8Lgbpu1n2IclbELO6Xg8eSwH
op8opKkBspx81Wz9USUanIb8NNLYL86vuq6+ahO+WC25WIO6xpHs5P+k61iIegsL
OzaKLEbPq4yq+fkaDhcES9qghVXIKKr9d1ejrYjy/MGXH7jz9mvW7n+i9F04TxJW
xQCvLLvvGnOI7xgODEJQ6LQQ5mEQ+Nqf1s6yNYnWza69VaUp4HtwjZ525yT4+wN2
KO1j5JCaatFOvOkxtCqHitVCq3kAk52KYVnsJMbrMOIt59DHZslWD4z/6qr48sCv
tVwQbWJnH98UuIzpotolg9ODPoFF1YhKPNP2Snpgkhk1ykc3bJE6Lw8R5MB6wfH2
Xl/7/lwse76BclTT5bWY+YbldO4H0kJe/psRT+cvhuAjRO7j5IJeRaypHdSjOncl
JdkHWoQ30HGSUcck5cQnbKHrX4hbjKEpFn9gavV8KulOd0jgWbtLeaI5HM0RwbHp
R3keJbAskdkeQZ3p7FXD/pWvUQoG8vFTUaNMrhmBN8y/BuWcngZVLmVeW6x3r70M
Stkl1g7Xut2y3/pw+rhHnzwDObpbS01yY/eGw+o6ISK3oE13/zEh/DsDntCs1T2G
8VxVPxIW5ud7l1OrHasRUgtUfdooIBW+MhUpSTiN7faDweKhhbnAn0kxDZ+DkFXo
JyTsBhKX+Wye1czJLHhnhAzG1KeCx02o+PXLkYmsaRP1hHKJsrqTtBiNPbDM2CN+
REtSx8cdadz9PFtaIS8GHTbX/zc4J+2z7tKwhq1pKtlztf0CLJW7+KBAfrQXcFgq
PC6xLPUeWJ8HLC1XqB5nYC81BQM6iNH0CZbWAtvPkufSt2W3ufDvzdyVH4hLWIwH
lJFZC3iP2It3G5KYQCUehoTlVb0wPTlZV8C6ASaPAERydya68Pp+VaGqIS8xvVEC
qBwXryeAASetoDaM6fBKEU2u4QuTzVRZRDCNf7o76FmuDXGibz7OYoFJGC2KtaVE
U1zWlqjDtUg+GSB8aKYb9gTPvgMol6DAryGbAQzyFM36T64nnNLYSUZj1DSdTg47
akK6IcK4xbQgoJ6VLTCLc55diKfdZoEjYwvnpivDUIvYkFHFMw/YNhQbA9rd0Q5h
jZ+GoX5FEFq8sqi70BZWPcWf4GiGuQGkaMSUqo0dYawIxRyUPaySaRculcgv6evX
nEBhXu7G246dDdo8NmsiiGJywv9lfUbiSqFEadPiPVPSP51b0SeaR9YRqevvfGgJ
Om3vs6bkZAKqBny/MTqKyxG5oK8XC8hFcNGo/LrtyV0HKI3C7W6Wudrobs0A3QpH
EPCwW+hxVg372ziJ7rCFfd73wuuaYYWz2Lk2nk0PhT9mXNZi0zWIhp+yzN+tN6Nl
26nYzdDKmyboMqn9gNsyC90vW5W31NzDpoKhEKBitzgLx3JMTYHAAQVJ2NWF85DR
4eZjFFiO4Ip41CxkVRikP1UYQO70JUPFbkYwPuAEfKz+jZb8J8NbMBNSBECg+nLQ
pK/SqFytQxom0gaEBw/3S3wnl+oLIZC3M5HAyvlubNdJLeQr7iCDPCNIO22vOeyI
U+CWxKxAqnp7WsXWr5fNP0620SBMeiQgk9uvz+hsqBmKO2QDgtZiCgQ0KwdxIUpS
E3MpvEF/dXcfZvrBI4Gg5ED8A6htMg/ZkLvNyCJfiWHGt0q1QwVVTzDixUsT0a0j
zhlIHUZ53Xb8Xb5526ntmHjorDvJkVEfm8KnsNtERRsk1tY8PBuFhESRvLUNFvSb
0cPzpKV6Qbs/yU5MSbKLE6HWKT9I76qNuOxmfCsxjGOfFnbSvw18v5Y0gDtAX4jD
JRXeDTZDAKrkOf4hFdFWju/sLJF+1kJX07eOIQdcA8ywbSAmn1Wapp5nrAPpdRA/
6Sz6y6x4hDqMNFuw9dGLG0t+u5MTAZ3tk4OMXDAOS5+C0egYh504IFgJwMsti1gh
HIZ+4xAbhp12+9HhJoGt1wyFFL+9Yy6iHZB9vAjTrUSrIrc92XyCQFEnqTjzY8Ar
uHcoc2cilnhdTjfSnGWI3Xa/G3hIuEzYRJWDIUlyGQoWzElcK8WsmJplv1/w+92a
rvkNdJROSK8S4CO+SwkGLFVFp/+dVCem4PAIwrCSOdG0yNpOYOA0l1MiM/+sIAN2
btflbaO0VIBMWKtO8gYtKC3O0xKk+j6E7eTE5QKPYWrVTjUPhUVr5FoeJOUfNBYO
d3KgEQCOBrlkBdNuR8lE15fgkuV1GL3bZG+FJdeaDtLNIRbNP3qEVu3b+AIT9TAD
gv9uqiSG+vkfZCHpwySKEwaJDAvHM08bHz30jf7667fOl2i7ocogNDxVcE23sJW8
j7EGBaA427T4hvQgG9D5KZ4E5fS2m/i1v+T1NFmK5+x7eApfBlOl0DHJS1i+JJNU
aIal2NVBhnYuaXs6Xr4TDEqywbV5G4hHlRchKceYk8TdxLJGDdJeqlhHPnvUsdVc
+9j1SjL++yIuLQsnonXU8wLZEkKw5DNNqRwvsd9qsUo+TSFdzZPooHO1/RJDtbI1
qRQzI3q6uQEWhG1QvuRI+DA9cF74aDnd9O0014dOYqqKJDppttiBUn19bvcY+bdB
ZfIqBdWxw2jlDwg6VmlF3M2lGSB5y2HqGGWwqtuvQX6WJ9BymnNzMDBqqDqlCR0p
w2FEbPGsH6ITKxWYekbUC5gc+caqXrKGaV3BUnmvvoDsi23H1SpwndoZYYbPwBBS
TMWVrY8hyc243xnJHxqA4FvdxbuRgkHPFn71fT9qEtEii/+daObPIgIA5aFhedi4
5CUwVT3MM9U+A9L1ll40yhNeV6+uQySJOurfTx+gg6ciMtjhET4J042TlkMOPXWs
fn6vLpeam+XKBlIvNIxp1+tV069GNfEj8Upe65fVgcnyBQqM6pG/VDRmi/SiTgH2
D56tbhbSC3iv43w/bncudYxLBBFBRVs41XJAfNmQCpHSqY4miv+cBi8k5juKOzNX
bXzGPUlr58DdcUxuPKLdHTX9JOyJijArM1FI63iC3ZePVC9A/l4tejtHeEclPEdh
SVX6e+3E6uHhFwPMhM5q0OWS151rs4yazkukVbTGDFCOZEl7ABzIa+X8prCaF9lj
g6VBNL5xEAG3sfV8wvxPKVkqrbBTk4+wJi1L/p3W63TWESnWVP7h8S47NW0XW9R9
H9mHVUdUy+c00A3bDbl+IRvoScvwl5ORFnH0OL3I6an1yfsnCjuITtDyKnh7hi1g
VsJ5HrYTj6/H8MSRSK7YSciPgxQQd1N0xcwXmWdSYfoES62qckMiJajPbC5JJ8WK
k99Du/9ci8ThHCnsIIVyDcIKNEAexCCOp8zpe+hYVKmckfRZ4GHEhFmKxML003oe
/9G+PtV6GltCWMmXfEb5CqN0TMQO2D6w+sD8ZswY98Nef+TXC67yrMLUBNrI+3M5
YrfpKrDexCBasGLxQhqZOs90OhIKNRNDMKf03Qb/xZ7Iytb4GKsPH38QQJWuTwBt
5HZwWqWVQSDswGh1i9kGVGDA0RPllUrEW7Fmlwedv/g/J3V1OJV5OqTO5Th2ahyB
cw2N/J5bR8hThaB1a2FMIKec1yjjccvGY8Jp1RbXs6o9dM2o9CH/GSXzfIn/Gh5p
MPrDvv/emySHHNAViP74p68IyNmtIBFKfTzLFe9qUHYxVoJ/nkMY4A8O0R5WE78N
UObXLaYIT5P7p2m02C27Yd7vWhgr+ptAW0Cy3cKKRNBSIPANnbpBPSNS7SDtyQc7
ssWrCNE42psGLS0L4qQ49ojPmxQeFC7S7XAFjhBfVfWOZPIqX4l40g9o59I2Btsq
1lYs/XYKK5qGC84lPx06RsSle6Nq0d0/59BWFkrtZuw/dh83Isw6zpFOHEiC8fHs
+oH0FwJEP+5KtNsVeFlPUSeOuc8njVAk9xOxYs95k+4ZS3n+NWylM/pHB90kUDCz
GpXLTztvMmnge30Qz1SfkCEOVovSlPvjMOAz1XkvWl6nqpq92Srs4oHJvf6j1eSI
AWu+e38laRpK5I3IBmeoRRLpchQfbfHYGUbbAc5vhPoaqAc/jy66OwxQp9UopwaK
bMwUu8tFnNqPlEb+8JVybuvJsOrpdVSSx9XEV+bc+Kd0UA65wlCaWTM1/iY7Cs82
dY3uq3B/k3Nmai7CHE4abIybIr98Y6D3o7XHOS1l5S/62GAlQSDKZyHhI4XZhogr
q2lgdUqMQirnLv0ueaI7q+Bv0zydgK/jM1+vsbj0++VUCo7CANEI8rEJbTvOaVrH
vBtkL3JSc2VywMiPuutmhJP123/vChrekoHnQFw5IFHAABtEaqHMhGFP4yBX0B+A
sdPMuyp+29R0MadcnRF1GpWVszCVysMeADop8UKhOvEGvxbAD3J2gXbh6/rq89Pj
EtSTVPLuCKGi4LjFDs3/KtjiChuQx5Up8gLM2QihFQ+7pM3mngF+H/RB4v8HW0hA
VLiEcilbS2dDCO2K2+DkoA+HAJ85A1NhWrmh30LxhH5MB69THEnxNQAhX/rHn63z
mTrAfxLrieBvACWiUGNnNxyOBqQsiHi8UvlJjECDGICVYuTIC2yRFA7VCwIIsYjs
I3m6VcLGY/aSo5dHXb2XqxWS/owqK8fmDbpaAcXhkytl1ARwmiEb6RYZi/mwzeyY
m+flEmKHQkJ6szxwAmUc8W/9oAzhm3zKpteNtdqitiAz9mydLhonwZmSzO7PqT/D
CFp2LgE6CXBmpZXsFxWr7HQUTJzWZ9baohgE7yM/3rnOxYjqPeEHvxt5vNitty+i
08SsYEt0FMRJ+A4oADTo+eB4teutLFl7w5q2FSqRyuSrtlx5AjdBJFZVJQ94gg+T
KFwQeW5bnDjFQn/tRszG4gHC2W/bbsmsszib7PkO0zQgRHc0pJkMnW9yFwwm7hQw
/Ao6MhqUclAKhKeJUWnk3aW4I8wSJldA9gVMaM54wj391MFgPczowr6RcL/s50oN
NZbauBil0mTUwXuAJB8L9OFpxFhkXlE8D/wPyA47ksi2FaDTx7+WnYHZVNy4gYLO
tCMqvfMu3pbIxb8Yz1a6/u6ECZWhECOW2KBapoKaBsR7k6Zdw/YcdMH0Sz52sbyc
ymBf9HDcR0rDKGBQr38PDeowG+h0j/RW+1BDbo9Es8AWAH6W3AbNkthZjKa2TBjt
ElUJsmIMmmd/OYF2DvKpMbU/1kLZvsLH71luu9oxEcbguF690BdGzucc9HmpRx6h
bEylrmZDNIHNjaiaryqwHLssX8CFEkFAQE+yjVzrChrErY72mLyGltoykv6IAb2E
1RMTSurrEP4zz9MP9dlyIoDrBy++QdlQ7PJbrAOz1pybc7UBKcdJXM5vEsVCN3JH
y4ANT4nCsibO5jwORiaER+P4jb2hzgQEv9iPlFFbKHDxrsxwEAhscJ8x5yvTWtaB
QD6cpJsz4qKMSzm1aYiHjbZPE8aqHse9Bb8aeDFW8VfjCu7j5U4BaBj3dMZbo9yX
YnwWL+pT3mx0pLBR7xGSEg1pO0Qki3L3lG7E2WmOun/Q6TwyeU27hPQWi0xu5lC1
I27hNEX6J4gMsBlwkJbsejSROIJI9a5PbVBJceuvyc5FGQF73oT1i5PKlx/bVnnG
iR3l2mwuSVsDDJKyyLrbn4gZBpjvIlMXl4cWKSKbS/RdnUvY2mR70B6VF990OliH
ZMxubg2OsM+JMvkOry4rri9baVjC2NJithGbOOBmn+zIN7AXLYC1KHKOJSx8KXwm
6J6CkgU7AfuMG4x2Lvg8gpvETJVoVM8r5NkrCeX37TXjBlRv+wYbJAUS44dCP5Wx
nF4nX0lgL7ivOoQ9KV0ccSQ6rKGOz1ccKCnFpwSDb6lZLqP8JhgpbCP1g2Yfmue6
IClOMwp6dm1eJ0u/BnZrVuzrHVKTcfCmCEpuhdFi1sH3QL557c8Q8sao934klPGe
vWkTfpyP2M3Vvg8tSgKS8mTH8fLuZAobiG6HiWbRCbyqGT2kItJrRmM6AnILnHhL
PDHVMuu3AY2X8qqtlPor6m16VRhfKI8g1P4ZIEprAclo76kNzAgM3Q7gYu6PyVZK
nCaqfi54C2QMCRHxhS+xgaiPFdcTcCXM9RttQ+nd0q5wxLwc/OsU9dN/TzB4SyNn
iJoPBRtcJOlow4wD+xldzhh1FS+cDyfpJahr+OW22rBtHfGUU25e6SmRNtn2Mvle
HfPPmePVqHxtIe1AEI9ffW3fxqc440i1pOWTvA//x1CjYaUDNsTr1+pVPZKAWvJK
2bvHMZNT3e8/GLKEwA00nUnaVwF6rQsj7a2s4xv1wI9eKnF+HEIwlCOQRiBl/Cp4
Wlq9xvkJv3NJkECJJASbTeEUclAR4kGKN/dfhNlD9nx2IxiClJGNX0VQ0V/ItBme
kS1/Pg7yAbrphcqqelFlwtRBZbke/Qb7QlMMDDinUfPe8w/cAiu1JD0zTPOAs81N
K5iwAr0ak11rWGtbG8iGUZwAYxpemlIiIZrsoJM7N70LTPvHYBAHs0UuU5y9zg8W
I4AvYw654oMPDznzpOeBFFtUnZw4Ex9LCQm26XxvoLaekm7bW7z+6S/OIHzwHmWE
3m58eeI8Cr07KPlsKv99NSKFjwKl7MzrtH53uYOx0Keta99SGEZE40HrP2qNC8td
23qvIvCzkaHCylVgZ9al2nv4Mbz7RFRxSLQuReKLN/EhL7K/xaZ3w353hafeXmvL
PY6BI7NV6D2oQybzy0Y3cI5wu+yC1wDmrMAgqoj+GGvE55n6/2s99oIM9kBDbCuA
iM+25fhJjFuP36CdUSlDwi4bVQd8qkf6esMuwlsjEzjIRWKMksmiDOtDY1zlEDH3
RBFwVQsyuUvsqiPhp3knJ5mnqUedmPwOYLNlP8QIoQtD4TZibNMcjjpCanFOEBBd
gRG+Guw4axpfGbIxs8hmxPEZVRo3OxKmBfs2I9wC57YLERd171mXZYkXjYkWEHL+
sP7nss7rJUyEnzYK78Yyj+ickPnnxSHJ2nAr4fUWhPVykJ1EBUw6CG+ilGayovfj
WNYprGAr5FKkN/RtwNsc1VoCm4nzIIWBsxR3Om91eYXZOAmkBKSmDgSIHCtv1Oiz
umvnRBL4US9FvdWPbXSU1vBjS6VhJ2H0l4ArW3Qh6qq4J0ugoaWe3B4ZukGoKcPI
KBGZIMmHbZ8idd0qD66bipZsl+/Erb7PUD6utBe3a9ore5a8bl6ZrnXwYR1H01qj
sJZ/Hkw3mwDTKe3oK4KrZFOtCfEBbX3RT+NWw3D0zXIV4TMK1v6NQb6I/HKXdQdf
0+ripxr1rvWyQwz/B//1cpyi9ZhZ371EVBb9eH4bERLZvEd0wjXI7Ya/F/ztZNL2
dxrzXMQb6lNvc2+jkfJ2T7w9kFqkGGcGnzhyyyylwY5Siq5oKnl20WFpyULLsiLA
yPDQC5cLx0c2Mz009Mzu75aqFHlS8GYrfBWc5QgDicDqg7ib0sDMXFn4jtxGDxtP
6SQsTlKZWABAwKaoVZ1JYENxOXcxn0Gzff9RQBg4uiHZIY5BWnFOpOQ+GseYH72B
7TxvH6zUpjLv/+pWxJAC8ira6NjkcpfS/feeuJjwe+PMX4oGkqMzhaOGkntY2FtA
zsZa4dpXrSZikN+kIPwgbtcihhED79RfrYzEmAecRX8gzqlglD1Q8fxJxX4pZZgd
CVtN5RV9cINXt60oW+hNKcpEbwCB8KHkqBKnEsrE6z98R/SX1QeJS+FN1rGoBy5q
Vd5otvau4r3D0Q/weSNe/K7V+AdGGkbibaBt71Oe0NpEMh138lsQveQOknbfDsIM
PYztCbLjOOlplVazO8dhQC1MLVXwAJcXPu8j8i+ZHapV5Q6viUEQUFkCeZU55Q4P
12ftkJFzoQTE5bP8rBrHPXxkQa2h8ctccfl5sfMsNj7A0uAdR859NpnE6uLL43to
i6uQOXwbBgPvsU5wla6gL0ch6oijqZHEg65x+KaoIWU+q1WTQzU/YD1aAVNpxCtD
LxQail84raulHeQzmRUEUbLPuypCjg6iVfeKASbP1tbFRzuvvEwvUq0Hgf7MER/w
1pgKhoEM9R8uz10AsuFj1/nswnj8BOG8iqyhJDv98yd5GT/6/69dJVopLhYk4XTW
X4et0FuXLb99pnZIUrRvtloHJcntveseIMxQAU8uZrYVMo8wBhppGRCASqn8us6g
ETNE2xWLCFSCxgKQT35M4a9wnaaH5HLhvyOYdStYIT9JM/Z13XN9MmBb54Kb0Bst
CSdHvm5KopdAP3TrCQsbI1VYD1k5GfEULf9rfI3nlMPyv0EghI9Kh+uRuVTv4Ams
GqkKIZ/sNvWJVaZgPZKxsM01Qd/mM/DXB3dAbuCoQU79+fmzZuy4PD9Yl+KekFMU
lPQQukvbzX3T0l9s2ioVQQTFOoVL/p1QSlEWdEQXB6UJaM7dBM/iCobRw0VAFY/i
NqLXxqPP/JQT9wA+vn+eR5Tv2m0nhM90vJTF38vvKuL4/bD26gV1NKo+czrbsAdY
N+DSLPdRAAEQFHJRMgM8QOPpbyFgBqZ5QrGMlqg4Ido33n2nbwzo86RKh37PSRI6
XZFVwUB/NrIQfyCzEMQtx+POpNZdK/fkFeWtwaWeQpZN7YEQEHi8f8u9w50r7Wcr
K6RSzOT8MjsWAh1ZUPkRL8osOR8lyz7yVj/SJuNoRw2XNN91H1ShDhf5wTl+66tc
GXNy7MJV9WOWpvXWRATdIH4sUwDKJdRuoRD8blJ1lCbYzJx35ck71tnHyjXfpv/Q
j9Iemh2CfW1WVODovs6WGk/WBElZlGeKd3J/Dj0HZV41KdWATn2xNz7MXXk2jSrp
xQd7xYzZkXBhZw4z6sABjiRzAt26c2YsdDPquVn0hn5+gRAs7C2Irmd+9xLlN8Ep
cM9OdT6JPSeh6mLhLZl9fxzj8Tm88QspXNyAF2wipS0bIncXzVd6ANg44Zanj1E9
CDYFT9znN/MMPvi9ToAHNjIQlb4A3jEtwgwxHpHI5/BoJ45UWAvSGCCx/RmXY5Ws
y7zshtrfaUK5Uy+I6gLNFJrZqJ8bM9BDcs2jiCLcYnQpyzfUnsIAmOs75lfib+zo
RMBcdcHZ6KaBwL8ICBoxFf+wxndrepC/5RMQw/NRpdhNzlsDzp+btvaPuHiQ1rTl
UyFMytJKUjQ/0osX+zO/8D97hRle7q3NpdP2rRTVM2QbMV3XWIX9rncMOvxeG2Wn
VQC/K1M8o/77O3mFhkq+TEvskGfZuwtokR+QSgZS5JhM1LNAzo1u60hEQKgBetUB
QsA5+MYKuBpEENT2OvWO6SPpMW8JfcT7AMQGqqErkktH70AKq1PSfmouI5OtBgmF
oSsNdrrcuBp9cWYCukLanMgGOh6S3MQZsk8BtQVviY6NZf3gOmnqs1CBncXKT2x6
aNwGiw5BXSrjDm2WTmcJiZ+UUrAn+hxyHwQvpzkySCFygywWx7czC18zqwb2fz9O
kdNFmryo0Nu6LCcYfpro81McWazisQwYIhSRgTnPnzRpTmM2HR0tzWHXiAp5hCEP
GB19CTSjfSseHyIUBH9g9RNeZXiZ4GoZNdlQ7e61BbgBvd+4suV+tY0YT8xpGqS8
Q2UEv9IJWAzjZYZ4Lh9CXQan7ANI2Hot4rmUaTx8nNFQ5jPy2m+Wt9RGOYzJmGXh
/wYGys7PSPQNccas3G58ystox8c16sqR5LsZTIHzP4OTIaYzWv5tbuTth0gYtrvw
9Mc7h3hCUggaWnCSL1dQodbG5xHIzjeSgup5s+an156IWAZW9an8AsefQ7eyDXL8
ikFxZ3gNY5b+bn2W++oKwM6rIgFLMxVa9NfU6BQTRj9LnAe89RqWuKXJIwOT1yaH
eD/h+3AmvkPk38PRkK+U5Mb/F8En4QHvI18ze+3MlzOiZCTzaCbTRd8lev115rxu
XEV6dHC5gtR16zVls5kFifwGK3LrP2Xfgj8S7uNi2mBPgC67FMmdsLL+K/X62ih0
HuYtts1nxTHBRMdBHTFJmQingjha+saky9MeBdlR1USxu3Kc2oVvtlRjc6rdC1kj
rNG1Jzz0lFBmNFrCyhp/Hr80Q1zC9J0KTEuXtpJ3xbIi3mGB/bzbE8+Q4Kr74pwV
PFftPrryi8RmXgA30sgPPgxgHjIDTCTEJI6MRZYwUZHS64nOrYam8OzNtBhAltyc
QYUbzApUNnHgCkAWwS/i+z3LfRGGbNPdwMmgl+/VAcNINV/pSz7dTo6MmIp5F5WK
olc2TuLp8PNZ67M8MOoZxZ3H5g49nQn79554+IdRZeT71slb507HqPExWb8I+8uT
CYZzayb+V5AQaXIVOaCZ4n0PTZslgQUjbeyKp5o4YdP1BOdn3XfDhxPcI94IGokQ
Mq/r56MYGFMuGFyCH/aaQzixcyEUV1cUxMUdNRFHfFnJpQImV+F8LKY7Js6uZqud
Scve3wgAkIiHna2Voit5PDh6ydzWrj/hmF+nMzmDyMfIDe2jwRDzrDFEv4z/Hoik
Y9X6mV5BC1i38VH80+mjRw+ABEY4s9RLRdtVMjK53umxptsmEpih9lqpHpYvtuq7
Kwy3GD4tZ+vyktbnB4okTL6wP8u3AEOhYJ2ZEE+I6cdm9AUxcfs22Fsu7oGDE2vf
HIa/QGymq24GkoJngviDSma1gg4xXa4d8uqjjE0B/WTij/c1cJLSEKOcs7dIxxD5
ru5dsbK/c14PMB9mwaxs8xaA6MS5U8BV6gZDF2tT5vHlN5sZlPslCR8fClHKu2YT
NEb6pY3CIx1H3d7RVRIeIuPt1pfrYzi30FTk8TIBUVAjBZiRV+AZZ1mxXBh+Bl4r
N5J4OFzpYLqlopcaMU9zKlo9vF7cIODzQcKvxwV0pJ8wcFEHNy37yk2Br8+5Cl8U
RlU2ryxrYPQ07yqcNqOcSUcYPnvuNhjeI1a6H3vmM7U3Bhx8CEJRxxHyi61eRGi3
wpWFabNVzG4b1quDJIq+r5UEYgPVppauC768k2PEARvupfZcmi8fisdbNypH7nU0
Dy7vA/9uP9SUisD3kXZOPWqEPlKtm9qDatBLZRk7Cgugwq9TsKdEE7NUovkRvTwh
XcbKJMDzXZ0i8U+kwjX1/w3aAfu8s3f3QNY4iS8YXuhxlblfbGfc06XdFHlLHK86
ZpWXno4nGwJ8IQ21wLJMjC+zDkxxMD4K9Xse7uizuHMRQcPsqM9286CGWSmhlDXw
0MavDe06HHk/4k3eFfEKbZr/RvYxzBKAfNDTHTzVgsurqoai5bwOdlvnIXqp/LFr
QperwpeCo+4A2W2zL6/kXNbZCEwnwiX9YP3ngeoiu8pHnyMTW1JLYRHxKi612E09
h23GdTTOUPl/dU+wf0zE/VOPwyLciaRIGcmcfYsb+RSvwz/0Pz1hv2LsOgm2DFkO
aiTOtylnWujDR+je/4bvPP4nEKbI8TNd6gdunpqovlx2E6WpuGY8gU8TGVIBWchn
maDgSg1JjR447UinAw7yNUNH6tpQtIuv1jGlB/TpYVDEwG2l3oYWRp4oNgWgtm9C
H6zkCFcAQfGd45oG5ozJCIlSpsfBdvCDXH9YJjLcgVxp+EKvXSm2waHKFk5SpQqP
/MD2NYxh7wJpYFOocwhcE1Q7M2ETSbhpklZFmlL+zRO8hDOr/dpdgGERvoEItiaV
SWvnwnPxS2nM67wlspYRSRXEfg/vohdAONHNOIPMbK2kaElcCMT1jJ0NeMLVPok/
nPhpFy591U9wfNWn056rxR1POjqVT27bVsRm9sI9JBIBE5mnf4cwIc6Rw0NbrT1+
b3rhMtoUTxQnCwAMc1GaFnPCT5Ar3HrdVfjSq+NHdKd+ny6VRQgJeC3G9HG12+ka
ir4VaZSfY2htjeJQ7vRRSnZaH1TfvwD30G6Aw2xvn7zLvuwLB+R7kAwsRsjOloSa
dkzAkAetXvmkZAc7WO7i6DsCnuHbrTXtyAjBV5xVwxxvfvrAIHzOK5Uq6Kl0Zu9S
y1VnS+JAcl35+K98rv9KkGfSXje4v+CG1GhJ+sHxvlD4q07nys4ZU/Ns0E0MQKn1
k9lvwSkv401/Mt22wweJKxS6U1OYAs1Y0V5gYtG7KZnSQMo7kbDHKAknV9TrX/pW
+J/tXHO1A+/WYt1lDHp0rMt5zuUC0u6A7evWkuCqFs4kvQdE2VBRHiPEKaZ4uWAa
vEUdnsu0Ns+xU0S26vVC4uDSz5MBf77kpWqrbzXbv4Im0olbv+smh0AsWyMNtoWz
/cJoH5afbUMBfDWHDq+1beF1xFc6aEy44B09GuU9mmAdWnyVFF1si1y8NzsBlRea
BQ/8v+AaOmI6o0y1Zwq4r90SP4Ba8fMNnNXY7cD14+6B3jt8UdC5CJaqCZkfz7qx
q9hLEWblkM06+Wkse4OpfZchVnTQovLlU9y0mxVALKXEKuDdbyasE6iF91ghWO4k
FKUh0MO153pcL+kGhWf+KwvJSPiLqvZ7Oh+GIBgwGMjfC5pjrZ8QkXhibvvEuQzJ
xS6mYbMxLTcD3fFOC5gSxCMiOWDdKXkPbRXOqkh8WYOuzR608VuQGA39QT6gNTl+
bumiCOmjFTZi6UvBii1kQB+aUNalAmgAE7ZvMlZTY5Rox32KwzxwktU+c2wmciq1
IyW0EHjpdrKrwcWoQkcb+7yEiWYdpDcRqHgWXzyH2CWaRZXfQTNShafgqslHPSUL
bFGwdVfhJMUICB+npscOL/+K639xpPZnMwzwxl/Aotp8xJJdaqY27yLo8Fnyj7UA
NHnZRe08xy5ubhg6Yws2lwE4kFUuwdaBKja09Uy4c+tt30WNTrhI/OzhlGf4Jltd
q6hUVYm9D9vIadd47GPwxx9GXN5A18z/leoIGtIBENaR9PvHO0nUx7o4LihtoIfk
rlEIM53LdG+RH3puAcmU6LZHfxTWv1NbCq38W/spQ8vc7cf7TZp3xyDH3UIwJbyM
UPzFpez3VK1K628Q8pd21BeD8IDvQLzalc1akNCWHzS+M0l3sXHLWBP5bywH2L9M
nKhebiwu/pLV18qOaQbFQRdKHD8DGJTZixqngOIHVr9NQPFSmMok4Ex4HD20ClGH
yayuIV/eMzmCMu5Tiug7y6d7y21wI2PFp6nyPijuX5HW1ov+0OiFxPNnG5AhhMyT
EPHdfRJv9Mm1L86FjmVpXg+2ZtVjgnBHZqnb7PtPU3Hze1O2TWET8TnyZLOouB68
3wqDQzuTkNhvVJAuzlUVyRLIVz+FLe0wK35y8oLwtWUKgAagjnlx8bOWVKVJvagr
AB7L4plVa5k0UdMar72tU3U8uUowlF5+EFqVXX9MUde6ZmvLrTg25pvUINh1+jO5
Dq2emKx+atV19u6VNVvKXEshehwQkZeselfvo6rl/nHljchPQNAvHwG4kdWf8YZc
MYsSk3dhAWnD3FdZXRneELeXURrULidf3w7gyVZzgh/gFNpwxgUbwlEbdItL0smv
dDOk/BqS6z+FjufhZqPFbDj0ARqWurZyM/Gs5+Xw9aYujKBM8kNMAvzfD7sCfwYa
x/bD1AUiG8oWJ+3y3a7lquEOBairs7FUWMph8sExoHO73NX9ugkX6YvhIZ+oK/xq
fqdSATgEj0BUMkymbM37Z+eT+ZU1gTBwL44hhWut2d+QQ2gGwTq/hDuWj0InoA0t
R/wRr3GPl6F1cXszcVtaf7e9o3F5OFeXUp1vgFo9vrHW+qH23wnZu2mFjPV2Jkiv
yMQwW6z+Q5OUHTPOcQEmBJs+IcqgMZVPIkSlc6l2lM+OO1LH7UuJH/P1gtB7zeGT
xK1Zyk8k1iWXRuTdEPv+dN8pR8FMSCwyIrOeqdr7UONFXuvsfczJlnWZpMI6aunm
/mODcxrAodkh2pcKLBns+3zrgodfIcyeR63KYH3RQ5dAhSuLEgrkUK1JYqu2oUDV
glIBiNLEvsrjs33HVTvF+x0QcBibajMwBq7RPb1oDMMNXRDnOyEyLyPtnJoks60p
0QZvxnrBgC4E1pPJq+yR0wCLvpX6GE8ZhmPmyTohDXA8ZZXQ1upztT68B1WLA+K/
ScsVkfy5QRzdLs2AySM0RoEuHSfP+7BP+272G3DxOmewYO9QJbvHyiuXcAgGE+OU
qVKM0++Xv5XeXfvd8Z4hTMBhJUzwt2epvyBxhyzOXHklE0AIRWz4nMxcJPsQttiQ
GB8gEP+jeN2kUIj9war1QIE/SKJwtrJdYGJt9IQss5Mbdi3ri0sakMKtaFswg8Qw
a3DXCCFAj/s4fIQClHrpcgwAwYEGiIniMOVoK3AuXi9sOlBAvhBVChUY4oJav3wv
pD0fwB18Ct9mAMn/uHj1tRY7J1adSjXPnN0mmNtLDhmsb8ULtPBDIpjhzr4KSsDd
sIkiiaLHo+2gEzqtXfqPblnR1FOBpzU7ayQ1ZDJucV9jVw74p4KtruLl4jh5M9BV
r4A/6FX/yBMy2M+4kqMkoYyrEr5jFK25uJVPvabnNl9GJGvOD0sSGNUPXNfGTcfu
pCvLFQs+K7tpSl58evbVMGWqsR/58bc/H/tW3FIHE9izAUqgfjS5+ARZ3TsMm25o
fYtE/XF0GkkFDWqZ+XSWXrcBLKfz1MlaavFbEFhOCiwFSRxBt6twBpm5xH+bafPU
8jxR1tpGceSackELxU1xKUQUE2uo8rfij2QsNCmnSlePm5qiYoew7aivLnPzfPN7
VkbmKSaWjqJs0lenadfUt+s18m3gkW60AxLNfa9nNcyuijJpJIGX0IIy/AJ4WeFv
b/v4QZtED5EK25/0l9MhJZSo+nzh5svxXwUeivcfoQwBq0CImzsJa6VaWtmW7hCY
gCoh3NGrJzQb+qfqECaymRqW38q0/iWTkMmvQsKEL/KVz5u0h8Cjx41DpOcwfEXf
JyouicUlUE/vx1ciJzPv6NREHnXPczOHmvfLzhMLE65C1Iq/MvTytTkQ0sU0c9VR
GzQKAkw4x/2AX09irin2qCSHo4Fkzvs83pgfAlop4FphRXmmeQN4/Hc12YQq/3eF
BLny5cvLLZNE0tYD7kFwkIHbXwv0NQPB+R8hwmSGJqEjVhuLxt4BOSjiomBmmCft
Gq9AxZ5UidEmMRA5KYewYkyySR60nhj1ed8r03Z9w3R7L/tYJxA+19Lzq0Ue058F
+r4kwaIzApDcRgVwK9m1k2+D1KOmJZJvlCfHBhCe/Fu8nEx8ORG+38LWoutH6i8B
NmqV87Xym0k3kr91UWvVSUFGD7EUcnq3Fyt4XFqFhA1KXEqgg24NGX8a+gseERBS
x1ASNBpLCrgkVfKhIDZuE3KMMNke8jUiY7ib+aot0KTufavOpDcTJvT3b8WTJi+2
Vj1DkRMoAGvjUlwqtXO9ESbsGrud5Oupz7E/uKCIE4Q6yGNsN+CSbPj/6aDiVC/h
jyUzH6Okr2wjVgCWqgEp2DmVQpiL2l2mYIC5QuMREVPhY62JCnSWwHipUPAwB3Ay
5LvPfW6BJ/C/L3z4AJLL3m0ADcSjY9zWs0fu0WHeX4xgJ4kQQfq5vjJRAcZilPXJ
83kBPREVjj/9AQiWKy+MYPww5A1HQdkJ5HgT5j6YTRJrHb+96INaF47Q5mv4oZbz
ZhOYz0jxVDQqLVyGF5MtmlFIkADK4lT3CLZjFRI/z+xxpVkptQnVNHWQMNh0FEz4
b0p3rpKRY/Hxljs+bubwDwaJjKSn8oFG/6AEyhZ1krWvznNKgwibJboQA02Hpnrh
cxvMNDlMwHQu8M2D/Wv4xHd58Ea+n+HxrEAdPiWP1QER2gCLtWNRDLG4/ygxM3Nl
OZLdReOBB05kkr7LYbWyY5jmnFD680d1Hg7W0HBVg8kyZuceB0MIZu3/lQP/610C
gGqe+KyVX17d2KoUWUfaLI/L16Ew/sGU4ViCW6aLZ6+RYUtfzinFG5d/QEA159n7
imhtQvkrHUhrTlF+Jt883V0usP5OHtYb+eLAqVN4AGHR6+FxJKbB+hlh5Ria10MD
CcnBgxgXAUxx5xtFNWIygNYaw08r8NOiattMD5yFBsUdVBoxhuiJqmXeDpf2vwHl
MRuZnFPaJ9P+xwZ/yzq7WnSQsJvAmIj0dDFhXIkoGyQlABEFNfOZL9dMI7WHXdDc
JrgqK7mYe3DYgby5Mc43hOHUXIDIq2VM2F0Hq1jGKTyRHv941nTL1ihNjy3asT96
ALKBxjJHs7za75o4hYboRaqfCVf3ezzcnAcNoN2A1MSAydoVeeMvFGlSkScG4FhM
4SoKLiNTzKJzMO+zXGkhQVhas220rQXZPYEyhLf+ugUiYjSERrdcqL+k083A/9Gf
25G3jF+qD3j55VlsvurGisbBuERlpb6Fgoaio9CoJLY2cZyqFnM2/es6IeKSxLCi
jHJQ26/dgwoA4tZ/A9KmqPFRf7y+pgNKx2SQGkcf9SeFDrzHq8kotQjHwGUNIquc
JaojnayllyG0RzPZ+w9L6oL5RIKZGP6/A/JbyVFXnjR9RBvZDpSjdm+jEyBUnDP/
LFOIm+UppLZ4Tek/avUfbxmmba1L+L660eQyhwS+HV8FTxb/EaT47LnraRUhp4pz
FXIBl1INwUsp7IhhJFzudDuOjcfXWYbYO3Vcephk/VnffpCZ1JtQgIcSpM2MiPUj
+8oosHbAQyL+Pd4fk7OT5bODOy5UCfdKt4cfaAim5Xwq8C5MIy4lsuf7Mg4iWwCT
Agq8si5KdD/pZyIC7OgA1p1hkrx0vOzjkqiA/5dyov0tFCNFW8iLhVnih6UP1XBo
gy/dt3yJTsO3HYILji+BUwiHL4qvTKWzK++dz0MXxtZYTyn633uo+Cd3SIlzBpaL
+q8XfUY40IoNwl9sIy2I6+k+OnxgBtKtscBRpUANdFDGPurR5dwsY2Xvo7iQvXij
FPlurb+IButEuP4uZU5scTybRe95x2eWssmEVNih8uvQjMQQkIFmr8/0Ubuy3kvS
I+P6YyKbRaUei2WchiOG2tfgaWqAspUklFzBxCJHQiNDMmoHwi2nHE3f5BAgziqb
LnG2kUlbsRr3wexR3pLumWTjpXFEoB6GpjFNfjKINmXX8XbH5Kr97iSzqsY6C+bx
it0QdNww+/1KXwe7fnrdJPmk9K/XdxQ2LFPSiJqLXKPMVJnDiHp/eAxFW5DFAfeE
nTTzNeZ4NU4qGXo6I5j16yBSeBxKkNKQZ/fv1jhx+MzB100p0EG0eGRmtqkRm8WB
SgDFwsC6jnp2ZIM7gg5L4bTu1JCxYNu2l9IdY7ydyLBNsDvH+JiK8flgK4IaoQan
FTnPAYvEKXPmF74QwY8izlOg6u+VHd94GVIlCXS73l/Bt8ZLv/lDg9fbaBWdVr4K
e6q7Grze5rdmWgkaZaPpW8RZsSb44u6Vl9zgP/1D0jxXFjcxTCN8ILIqBpVg804N
WNzOy+q1k7vlIAYBeAZZBe4OZkj3Wd8CRqQZgEsV8MtWoms412m+smcnjlYEKpTN
mk0WO2A1iws95oMzNlOYTE0Dqd+U9A4baltah1RGxfXzZDRHp7MBw2ygr+TLxGR1
aNQ2+D/QtUPfJr4413GW7dC/0RIAKWGYLdKSHLgaTcEWAS9s144qsOlEOT1K1b8w
RJJwoCTdz2AnG2sgJljyPOR7MFGMUmiFYZJTVJcuVYFWTQnjsdOzU14+k53tlmTB
rzJSzb7aeJr3ylh7XMTF36iow6937g0PAQMTYtxmjAaUnbsmmiGnZpR43DN1MWQD
UDWVGBbsszO3Xyf+bvc9yUXpzdBoCq6Z6sLbgG5vshvD04I8LQygqU4zlmBpVCfX
CHdN9t7xdceajwAG498c+djPTB2V8npuBrPlerKq6oOkyH8hM3j6jXCWrAVYtUbv
wPCMozr00qWvAAoupd3Rt0j7F22gkC1bXasdfJb4mx02DNxVbVDts1h52fcZrjLb
HL9G26+VoBbLDhRB9dBXcokWrPjLLKWiDlx1Xarkga0rJtiaC6/wu9O9uyYwWU5W
VFF5FreU/Pqh8qJqmdcD6NuyAg78qiCAkC/g4Vn2RqSPkObxu87Yo2dmBkSKhkLW
s3GJJOyNsAnTFSyvNu5Y3l78kTcyiWK++kDAZSEOnT0RNmrtIJdv+gzKEvDUneJe
klIqbV2lfU4bdLLAzvEllY1/45gTLsoeOh0SLHUAnLh3eMhzN/5K9gu9drVf/Fl/
U8+mzuBV+MWgAmrDip9beIykL7ag+dB+LOHHPvcSg3EBOTFoCQk7wUqs5WSf0PRr
c97BVauIb0q8pIsXraaOaGYAeZX9BqaKQLSVfB1IZ54uc9Z1N/mywqDJH6+XPDsb
CX2PTehvK1KLJIpoUgIFt5h3aV2gxjJLxl2cqvFbaM12UZy0XqjHnDm9wstGfObj
InUj1vlhdmQI/HGqfzS067uYs73cHSEPaPDgi17zeSyAh3pEBb9eguve3iergl+4
kRxqUdaYzvtRbiEyVGPTJDXl2rjh5i2UYmvCzSkUM/UH5eCL0mQYNTFsI9YtZf6A
up7HHgL9EvZtlZrANIx5wxfKQnxuKdPnEeuK+4T7PI1fsqopGI2UK3A2ZW4cGiX3
eZIO92ycO12zM+qtqw4g2Xw9Ioy3hGvSdZQoywMzzo6d8SvNGnaYzY3+yfMuiL0x
c7qZHfYDRwLTzIiMAHdNQhFc0UBVxfTQieZrW0Ll9hbQ2HKjCkGTwCgjqncvrKzO
hu0OXyBevAFADPylAyi6bO9AV6yjZbT/eKbefHURBJePIZuPWwRKT9nuLqRGpUgX
LV2ICSC/vm8x9IpJdI3xnVBCMCL1pHXE/qLONB+f6+VMhe4ywzE7EKKZVEip7oWN
0X78UjEie2YDOXumc8iwjBHErrO/9qrMO9AQqrwl/25m6JZ3c6IzS8yXxXKXsjIn
Dpzpp2GDKlwQUxa7MqxE/bCXsBBn46/v916JLGwy/c1Ew+osg55Y54qKmmpwPxDR
QUmY3rboKCHa4aH276Zxdv9M6ARSWl3Sz26bhSzmbTPg1zXldSRM7BuMJiKuYWN1
2Uc3k5GYYRms4N5GmhaYGtCAjCxYc+h5uTXnreJvBMkmqGyUG+hnQ4yYSONXJKU5
T43fY3FKMKDfUJhlu+a/5AlqNb9D8SUMDs4F9aT97hT1Lrmct7uyjeVkNklbaGkI
ZLZtAkF/hGYxnxHz2VmBkeaq6Em0K7qsEXIUEB29PYKn/40M410UJnnQCpXOlwNe
5Xuae0YNxTEyqAFFU4imsW082qlpwWCmLnmgYhzAd2IpP7h5eYzD39wyUuGekROc
xK02xjltbBf14q9jbGPbum3xuPWrzGi3qgLYpcxfhyxz5XIKL8AjuOUpotJ0WBeE
pP3B1o7H5r6W/oZHohZBnkMsRx1APCzwtSE+RFJCKKZkS1YUAgNAdklqcnjqem2W
d1KWFs8EcXPIyldT4NyKirq3Z0pD1c42TQRDTWNrXzssXEsyczpGrJGFQzUd0FwN
8mVm5tZ+Ki3nZZO4NGLhNg0rjhOSZIhubku0v1UorbFfbMt6AoY/lTWg4bRwBrJB
l//wYZoNPKPjUXOl0XnlfW83kpbiN0A+iuyo9sMHdRvmL41tmYgq/UhPO1z7JjeD
APEOgDZq0hDpd3stUU2chjdjcO9Yw9rz6UnJcNjJhUG8uXO8ANJ2c6AS7gZWUFWz
ZXtp7XXV0hHC0DXM2kX8SFxp85QVA1M5KqChSDwnkKgtnmwzWorpb3Tomx8RrXYZ
snl4rtDMTY+GfM9Z5aCETTnuEJKCyAH+pIbvueQkMYfX3tQylAOEcd7QTxSqHTCa
qALItFoI05f3HJ9+GYgP7CX0rFP0kyKZvQKMreJdphOm/RuU2JpplMefH7ENbQC/
j+rqTuaVO3Y+zDkRyV2u09LqlXCif8g4J4ir2/R9+Hpadlp4eaM5pNlDCiny5WXG
RjuVjtF75PbUK+Qq4IK7Zrz1MYppBg+LmnliRCg0BiIhETlmYwB+i2UTW9ZKeWz9
LPKdAs7tyE3WPPx5l2kSVR6q+pD6gB5/wT+ntejFUSyhUD4hFr/GmM482fhhPY6B
SHYOn1N4Jwm+/um6GM2ioqzY0CH0Oh93WiX94BffRboiFwFp93c/6LtMVRjLs0YW
66X7d5+XTADgP8PE+v4WhIOgs8+NvVcmcLc3jjSQD2UJzbtbiDYiu8F68U65SGA5
zZd9Ot+98StJtE/JCz2YkhQ4oiCXmR5ehn1xcCUy4E3zurjbvp05Ge0OPn96iySn
xitG/yoOWnBPyo24Z4tQYwOWBbHZGAEdjJnHtfgkY91swbARunc2r7JvOnGbCRZz
QvZz8wLzpCIFTA+viAj5ddxLmexTKx860jyb7TGUetMV623I8/GifPJI/hPXTs+b
JSUERLg9Y/cSNp9zBkCaDEfzCVJv24/M9OvRCIU/k03qF1OxlpcOjgWL0z0r0VK4
fyKRhzqw5AZi9j10QJDvSeVSbjee0W84D0xUrCP0TJjBROLhEOAIHx4DGge9MQCB
mEaDZFFa0xvBrQaJzU+DJzu//IA2LRtwhX3c/XDcJjXcKufIOSub7eXr4cZwCjVo
CoURvxlG8h4hkDZjAnFoIrpEtRODPFv9c+6fNHfVqWov+XLEE3bVrICPv041G/yq
E9zpa8SriTV1a8xOtfUht6nj10DKyJXIMwAWDvEAUbFNTvniImLfLr3JlNR28sTD
SjGhigJg462wP4jRIDybXTJ76vNE3LX+FQiGrCVIGTLDV8bv1p8o9M1o5cfOX/ez
OPTa2bQv7JGmCvOBExdzc/2UygfK9oVKbTJLT8ODCZQvlDQ00KefCzKi64KQieZ/
C0KO90EBENEBaXfyXQCYVJUIfLuwV92GPjX7hN3W6fgqJUdPmgR1bWO7TOWllabe
CxqurkYRnZpgAwh3NNCAvLtaD84JvoWqNktuSh4Nz5RJOgHEIAmQ1Z5xwxrWiaE8
UzECg5Q+c5RsBlRIxRrYMEgj6bMEIBuwGhAi+oaOGNRoJyiGAn5xqPrs+treV35H
ouaGUHsTCBxmN8BT6DgCBYJwwgbfM4hVI7xh5sm3/ElYkTSdh0uLc2eXneIfe62g
H4k0Fl4XfTeoi8Y0xK275sUoy0SI+IabY+S6TMAujtyS2INwCYWwMIIGcg31JfN5
Y/mQahxfn4V3EBUtSQyi1XjJJWoy93rwB8wGAZcBbKRxoWj23Bh1i7iMRyuu82wa
FF456BjpL7c688wfdGWV42VD1QL5l3QLVHBYnG5KKMxKCupxk4iD75Kc6lCRJLjr
ZRoR/xDy+67p/Q7x0C79ZCPxpv8EGUQ7QZ/OUJbBU5yNESERHycsLdLPEsVHW2z8
22fyCGYL9XO8fgaZDO11vqGxJ00JdjOircXTWh9PjP+aEC1HfXyVx9KgaAkgw2k/
93z2vWJIGiNBnaDXO+KTYKwtYu84ly95UWD0FIPpBO0QcP6aOzLEBFPoxSKfeTWr
/UdLeIKXfcNmVrigXQsdGeCzZ1y5cdSKCYKuoPSujgnQJiFDmqYiuhe9npLgjFIS
h7Vy61BgYRVnndIL+x76T0JM8hCnGbxB75cNtVXd5V2S5rpqbxcCMaLKqZSPXc+k
LzX3enfn8o/6DScwCOEAaIJM92jI8Sk8yS2b+YOLeqAnh3Pi0QfqfLIJQmxwxGdM
cvVzKe9yQs3wGaJWg1ZyeuyvERYaFN+THThtFbhzj+Yc8OAYXoFKV0H/IwiOgTo1
w2uvKTwTkDAyws/eiTssaUA8mZ7d3HOC1EbiT5jR8lCHi4vFAxapNNHfLJJwBXsW
2JpfYGn3jlBScR+IZOJzYfBZ1cqPZyWiixwtTzISEwQxp7lGtGWja6W4LB1OtN9K
ekly8I8mX9HgpG5/wCDMVSBi0ytA8+4h4KBuQ1fQ28xLw1lhLDM5t95GFKOS0W4m
1ipzuXqMOq2b957u2Q++7zTERlBTaptY+h+5sxfkA3/SbhODYRgrt6tedmyHMwQ7
U2AuBpBcq6DAdVcmyjbPnr+fp2WCXJGMAai6ndQsGdhk1ztrf1sTL/RtRioi7ZlR
wMM05urQAwPxmfBmXOXpBNfbr/Ghn3sq2QpqQr6pFGuFtRd0eA23HpkUVlC2ynJq
xr9CIVs5Y6oJaSTIZf+iXtebhtHTdPngOtpULti3MAT1ZfEiu90U8qS6uYqvI9eL
U4a5dNkAoo7eT50X7AMvFQfyrHMflYpUG5yrzOPA0zqWMVPMWb6YC8koA3Qb9NPU
Pa4gF1V0Rsw18KlV9diRWuo8iEhabHvl2GIDMe7kv3x+DXBmwNcWLvGEux5G6H4q
vSz8kQuRCgwenF8Tzzn3EEENchp7i2H8pqzJ3jJlnYBGgIz8TH1HZoWsbyqXdXPY
6OQ0LNbBp7W/2z8MCuZvbzUQ7f1mDKivXH4lY5lkkkoYbaqEqqmP2ZqetMEAW9ec
VTXPQ30+yI6Dcu9j9udF+Vayh7HJPw4eYteUKttODiM2bpSwnHyBI/LWBsXzYErT
eNbnprRY9oEwp98Z/U3vyAx0RYEoItoUgkIF9x+k5vIbtnAUn7E3X6ogTvaQSq3Q
S+UAM9dFmBAlg5dC3nNXT7BWZWqrRzRs7YBXQvbxP0LHBhEwGwFDSUG+C6KOb5de
+qbyAKdH4oiKFjBi5qlDKrtvhEcaGQ8U2BSWoGP8EmPWjbfZ2BICeMFDPbwhhjpa
4EiaqOb0YiXp8gIG8Q4g3F/LaD1LC0SxuHTP83nXaXHd9uDiwTDIYyboE0RPZrWf
8kXJ6Nzu0UI4N+KwxDlNKo963Pp7/3JYxRmjJkQ4+K1eQ+CP/gcdIlKIxFcx8WYw
5O3boA2XTfa1rkty9J7mo2vFHKGj9JTsbfh1D7dqk1JwsVqVLq0/KjzEcuZx/0uG
TyAlL+PosKvrVLMS+ecc0ftSG0MiXvq0yWylHJISew1rs2tU976gI+VXDmJpar2p
hsma6Ubr1yRZtXfENiDUB2gvjPFh1NNr+vDsJFjXZlAW3po1IqgzinXAYHZkdwWy
JBD5Ax9KSGXtPXIM1txn0936Txv25SSOix8ZlpP5Y4sEm3fuy9ImJSVJU8MbjVWQ
vLccpg6yZaGnV0wEPXqunoLAOisCeNuifYsaV7DU9l2+Sb4KkHRvJtUC40FT8gaX
Yj/BaFi/CWN6lA0u/3csxUiIaedqjLGnYtY5WK4Fh+ExQKKiScQmnD27L1Zy1RWk
LHu3XGX+myUlcDmbLBxZfyokVTJqhzFr7GfuyYfa/wAN27mrxl8eznPI7BAtOHd7
DYJS3CAsioqfgwKBxHVpo9lBy+4qp3fxZ79ssr3QmYrSIxmCxy4Be05dcDScuV5K
tliL0dSmmpH35gAiXlh4GGrnoGCis6MD8ndrt79d1AZ5brzq8M5OXgn8WRigz1bN
IY/TVZ7+cw9Btz6yatnXPmOCenud5Cgiseqp4RiVqdvrdy8LnHy1NTxNcVZNSD1F
sWZIP3bxEi6bvQ3N+JEMaJEQUWFCPEUAR6m7e5R34b8vGi7dELiUD3zGkDFPT8Xt
YFfnQJ0UQxKRQ1ssLhafWg0J/6f0K9KvLS+WFGTyrbE/o5no79+iRHRA3043f2LE
HpTcELm1BRiy2qywdmk2Wgqn8b9d7UYfJhb9bnSeI1AjlUO0YOMl9gaV7I94W5Vv
9PGsREq+41Wi5NKWag887b2hobVq2JMEd906S9OyX/oA8sJSZeAPzq3viex7ndsV
JMrebSsM63WW11wPRL/Rc4decFj2ET+V6GiIDdrqVQDLqzDsV25uSbYWGS9b2dkz
YDoNJGFM/gO0l0gaQl4R9kolWUClQ2Ze3FTvf1ZLTTueeMARAPM91uHr7bTKcV6p
0F44QphkOFAEhPyLfb70A3eblOk2VxQrPOyINtX5UIZrNWJuObvl5boy2+z8br6v
vzLJHSwjs48UJPcQi0xZSPfBRWMDFczjNAIsHTMt7HLsHI8vEMZyiYoQTVsbls3x
SQeFwGmlI7oV+XRvmKR7ymbTGAnQUzawrd3pvLA7gnzEcqhylJDWYo+iVLkHgZoD
08LiBqa/qpBlzd+HS61w2Mstcoa02RmL8L5zaHQww/tGy37vNoAw6EuvhBLwWL6p
GcMuKjQ0idgcbfFa5NHBYkBX/coNQukZbSL+JAodm4cby1V6luMH0ha65lr2Ol9d
ajbeLDY9uOJGku3aV4qlPOLwZp5aGshHDLcLksD+pWlqMnTYqAS5Pksv4gDar9TT
yZ7XB2mktG/EtAdgOIU8ID5e6H0SGV4PYa5xQeoWcRarhaumIBsru/J6DAJ0LP7E
yedBVDtkn7EOUJBdpOqn6cJtILnFuM4eWi/Ji+YCWPyiC1Nr6Iz1CcBSt/N6k+GJ
etTAhaQq1FyvtM0ntMBVmwWZiW/ky9CW0oY9KD4jk4D1rjoVCPakm/GTo7twdTZ8
s82sCBVb3ML9QnBOYewpcvcPLeO5I8/as0gh0umUUzZ2239s+jEbFcKNlTmrxyII
eX805/duZXdW0i6zwC5/nrCiDYxL5mDVci+htl/j5wfAp81neQ4MfUPjtxfzc0tL
Vh3iuVLg522painWTkBh76etJDhLpuEMnESc4c2i/7MqBUd21rC230iSM/8CWF2J
uG6E6ANjIdNsayMqM/wB0Htv5SZmFngS/Co+PdZGaStc3O8eBtO6W0VM+5PPh0pa
8g20XdmMYA87/ExEvvRwXAOMO90JxS9h/aGdMfi6ee7cKEP8EqJKEDUfxujUaNiO
c6ZZWhaBOijYEZswIZCuVPlcVVFZNn8XTcbpjj+XJjJNw2xL9R+J4q1p+KhocUtx
A/V2wjma9LMRHh34yd2uq+0jjVYOQmNjTkxjTrZbviuCIJijLrBF5lswCTaxzQF6
VAQYLNseDXfZqqsSkeprGYm+0EVyjDbjATXElCSnUn95EoF2tC/Aka0z4iOK4WPW
/bypyNahy9WJfXKnQhxDMwPpDv5TY3wKK6iKrEIt8JR82FrLQGr2RDFqC+VgAs2W
30zA7p/FEUP48voDV/W9SQ0M2VecFVcgEGg13QlvkEUKHYoeFdvhEs1Qw8aXbWaR
6pL3Dud/2POucn639kZbjtWLFfQQUOiChsaYHjuF5xIAE3lbZghYZgQdFlnIM3Vb
mYd85g+OplLZHZ8HLcna5zYv/pCCHPyyzGs3862omj5Fpas3GJN/Akx9/aMSMRk2
cVBy+sC/zZp0hmU6VlSRyoIb+LVS4Q7eRZe6ldbpcVzZ1fR0/TH9LwGqUWKUwz7Y
kAfJSsOM1eer3VOlxvd6rlXKZG+DO8H6El+ZQKC8ZKUoIdZvVdlX0C8EcQMEO42W
myI49h67qHOcci0ZxjJUVZ1YMygDihfRd7Px0ahfPAhV2+/q/tysMmJnxz0f1i7/
QQKLkdTx2cLjEqmfjnbDv8KvEvzeJPziWYopUeOp1Hg/iIDQ5W2wH7h9wv6nwBSJ
5l3v35yPxlm2QnAxW0VgA/5T9rcTMchBWbJv9wHtcq8VBI6tEER1PFTwiuSC6Ll6
OPXyrpuxKa9guNp6T69aHG4zeYH/y0lhJywag/OhLjNmFwiVoDPWuUZZi9WNDyl7
fZelC1I4QZmqdJtkiRbSOG+v8rCJuONeh5Ynf+BmAPB2T5XOlZxVhmoyyw0sP+ce
MCJvyJyCTLMymI6CRRAmHbtAt5viE/ZEPOoPfyGNy20m3Y0lLhz55nhKzzRyTc/Y
nT1AXm+DO5IzfPomRkji3B+C0gpK4tBLSITU1UWp/NRop8h7cUTNly10ALc0I/Ia
FlnzTEcHaxTtEIXlg4WDJetKdRdNBs2wUqPa7VW8fjjz9JAi+cl4NK2Ln2P5T/lB
UXpMq4PdrOz5BXpjWXmGgEmnUeEzT6J7uxwe2Xps3fnkleRG+fYLS8DSKrfXP/Dn
4VZ2VUtJ78RITf13VEAPg9jnrP0ATfYchhOKjjjilJ8wSxJqp1nMc3CVjKjMz0ZT
Q6RwCfZH70OekBHS2R3AUoGPw3xXYliWcjUIzkPcUdywKoTpqt65f04/04FsTIt2
hHUmL/UvtWC3zWvF6ZooP7wCSTi97esNX/QzZRemUL4gbc2RhL9CLrRIsDLiRoyp
aOfqDTU9cmrxcC8KrBZnSkmIHD3+atOiG7vKboRbzGV2GYiCJcb4bRn7iUGBCC7/
KTdfuVJ1c3LiP9aYbOpJW+oSRxglJEpuo9IffGI8HsRPm+CYLFhYQxy8X56zufD1
/e2qkmSa/i70zmnBA+hragbOhgWYAo5CiT5XBGUfQhVz/pfo+bM1/1S14z5f1HPt
ls/8nEbZy07Jqvrmk1vg7FVh02rMg8Dn2sj0XhvXl21yt7XtrmkO2ZGdHz/cQMQX
/XKtjaxvyVqsmigVKExkMONzviNIV8w9rb75UaUDw2lfAbyW00eeA5vgp3sl3oNj
rQX+8zxN/NYVswi6tIcH7WAJJf9YFJpb5JG+9M0T9xrFC8E4NRb/nYCyi40bKFSa
kPbIEHZs/SBVq6OMvyJKhSvXSsUCQjUcOgn+f1LsoXiFK0qJ0Hj8y1bGgtQRQiSp
BjbNlnrAuLt1QS1uqY+GY4PX40qRkbbLlCdZMSPSn4kx7uHVlxz4lKybycea+/wc
Z3VfrVacax2bgOqIy0EC02+JIxarMWcrvZsEk3/DhxtGDoqf7Lltp2KxpCDSVSPM
gGJl5DLwSkKgFi8nsNdYjVIkU1tagcrv6jX/jgpxW1C9YkP8HyhiUQWYkv7OgPyM
d1PrYlCeWm7UjOx9QX1oYHU3FBydJ0l4842g4Q1mAETbJT+A/p8bs7a0vaBFYEFV
2mpQ/5hTErBIJ0OYeuKDiwbzTgskeJjk1e8W74LDMP61GlWEzAg2Mi3a6Gdc4Sgs
XvBjWlyq4zP3yqyEm1yWK/YO+F4gBowovNDcJtIOfK8UbZi7KAhjuhB3hLO+ELdz
QeNspB0vjSgqEGRKwc/GkYXjrlkf7/Qyu/MxEGv1NLXA2DLEXB0qcMVIrL2TzF7t
2T575BCM8jicpJve9qtJ2j7N2eWhtMhnn3FVSWvlZXsLxUdUUFw/DNmQoFR9oHLS
nTPXRf8wIyESwixCVNXDbGcJoMvAFA9FDSBl1MKhiG6txS0ZDSxeEg4yG1nl5g+O
5L48ofBcMlvBXPUhQGrHy1EwHGMv6t4fYd0JrdHY2fz/Pb8KMUdvf3R9f7FLR5j8
io42RkMv5h1q3+SqRY7hE7fmAS7CssemeoTfRHy1vV8JPSJFmWj3To4lAjta9zdo
xMqdh3AEbA1WAPrerdlPSG5+4Ipjwp4FfjykTgrZkNjHtbuJxbqHrqGwW3LjlA6W
h8IfdC/brccBU9JMwCOyDgkib/k5gqcKUJu/c/ifTB09GgSSATDpVA0ATk2pL0bV
VJ22tk894NTa423mYv8mPdjgMne74G2y2j9NXkVvRm/B1twt+xLRUXedbMCbFWBD
XMNlCzXdJR8hNaaH57sS9/ePaDVbA2T8xrOtfDSYdcdoW+mzNnh1gpHq7q2YOiYM
QoSIxT3IdQMBAaKjUM/TrCEFrD8IeplKZKk5E8OhnfOX5gPCfcnuTJ1KVmH88Q3v
4GDTJx+Kfz9rTLke7jwTji2II2eG//znAr1RLNYjBXJdomfwhemQyrI9Vv9IGu53
CnS0XDSGKIp/TYgZyWNlAfmRV/ZcqxutY8JOrUS9scrqRx+XT/rHMNTTzOWpl13h
zsfaCeUKxMM/fr65hKKvhbaRcSVvd5wp0AaYjfZu09cfa/wiBCcN+TP5uWey75OF
ubHDyRhusiWNouB2nFycO57oCYP04hshtAbSMBdrqwVxtapXoV59ldIHHhEIGDkY
gUSoeNfSbGNcGOFxHKoX9p909v/6PQ+3olhntadwnI1Ov7w4FZF8iPR6CH8FlTNi
R2NUMbmXBrSAoDN5OGrWda8bReG0nbsN2QAnLeJn1rvzqwyCzndXvoWIKKZZYAyx
4wonDIKN3YALEajHwHyGYu0xFDIT1C/7rkOVKXyXdu3SVuJTbIwJ4h44G8zabRUM
zB7ufOyq7UjVJ7fCkufQ0vdVmeA12qwWuqlC1sg3HjLoO9e5G0/40pAgi2cO5fFm
Y+59OcUGnysGWw49wqwoIyA8IKnNfBBhxvuI7bVIh6r/fwZtHC3w8za6YRoMm2y5
X1nrxVQPcZwR/6A1bOAvCjlkXSfZcQ9Sd4YnbGePAfRJEQjSTlwFrxrvFjw1VR7+
W2Id62FNOaJXP1ZaBZXFXLzzCL1/LjJuKA+k29hm/Mu/bX8COWZ2Zhog1Sa89cMc
pPDkvfUbSBsZ+/6BkQig3ANy3KqauJvQV3fBPlK53SLNm3NJq8eTr4iHxo/UFotC
qPTd7/U28CNgO7hvoIdRkVks1Pi2dEcVFaERxoB3xllJ5rOzRkM8WqKTpx69IfYj
dG5gUmSGaGVnlmJB7JZOod28Qb2Q+YMi94u0MJOhMN+e67p4za80i1O6TaNPbl3J
LvH4v6ZBeG+ja0tDynk1UE7QNU4aBjHm+vQeSVM8HZ6PdwEfkMm3edpIBuEbjpoD
FpRgqaarHwp4+N9zPpX+8KSdDepcQ6drRdYRNo4tEuIEkzJ3uKgPIVXPKAE60DI5
JbuJpO8riwSc76R3D1mvk6ORDQQ4/315LR5q6jP7k1/zRUdqL84A4Q42W1TqlsVg
0687eZGj3E+A3andOvrd/gmGqy54C6RuA8Lyllp84jzAUw2IXPL9nZnYx/sj8Iic
Fr2SSJTifimFenOfyWH0autcEF8SXoN9E+22qGn0rJI4GCEPz9sUM4oq3kveCTHp
MwN6hiQvCcIsIBH4M8hpV0lL0fmNFjKxHbJ42JcRcyQZ7iSU1rgIpsxUgTDWghir
HZl6XsxTsAD7BuDjVaW+nkdFESyAW015nogPN+ILaqK0Ub0PlLKR2xYR+3gIC8SK
0fgTpFrm5wvFU1ojidn0nY/bF3g7hcNlDC6xoM93B5d5EDWztLmcVMNxhhEtXAU2
kGBM1tBUnUBa6e+PG8PyZg/tRD6MSzLy/SYEfI+eWZCGflmb3vpBgTB5eEcKa04A
q0Q8RhEFIbsrNZY61vbC7dbPkNl06DC7FJj40O6xvu8HHghK7h/zUur0px9HaSqk
n3wTb+6FlnJOKFphQ0Q3SeHDDwaO7v3jF8WK4CREYOqhJVzONeZTtKj7lNkEC0RL
WUUJbFX8K+khm8XysLMK1y+Jdo8TQCdKGQI31nzEBPWRKbPCMeMGG5Zf6lltloSh
TufhbIrO6AIE9J8WFhPvVY1cnPmMSl0d6nubv045qSrJm2W4pbu7tPEC+AKlkBoD
PVfBzkgAC7fGgH4D8COMWGMhH4NQ10q3hPe2NiqvJbkPPE0+Yg6Vwgklb7veFWtH
ts6gt3CCwOsTcLDZB46z4PAhwGplXgP3Dkks84WhdiqyqTaux/ZxVrPMysjUxuMD
5JM03qEwNK2aQeuBWJj0dBRPbPG8lo223e51HpmSZEyjbtdY0Lw8VUgFyr6t7YY4
yxOioGNnZh3ueZ51ENeJi5qULUGblA1FDgevVO7VhLgnbdmQHLhv4FxK/An36q60
zniy3taUzw5Yh4dBwaoj0RFBnoH6kmEm7yvIKVdQeJt7qSg7R0Jvu0h3SIdEAwye
8vL4HfCx29w1s/A8aD5KT/2YEKjSdhr4eELUylMHUNV1f3uxwnJJ0L3s6jr33Ptp
act7G5rgiZ/gD2oAGfWecLHLN+/qv6vWaFZYhQi9ZB4eWmRUzoowfUBUeMdvRWZT
aOJSQDPz2sCnrka/ifzNiWgfq7LW0s1H0KE1niFOh9nwt4n2VfZFweBboTDa78PA
+f4UsL6NYdoTCiqPWC3nn+r3mKadDrnIU9C1AtNry+4bfCqOYQttBAMWU6gbEDkr
IJfjq5xf9g8g4bEOHqA42yVAyMvIFBBf2SI4q/+87p7HN13GpAB3Xl8FsWazubP0
LdniWx1sRcU2w3oBxbQFb9MAA8PT3ixLGp8uyHPnjCxbAGcmT+kuVwWeXduSrlp6
y7eo2QaquRERxyp6x/AAnRvWsnteDLjZfjUvIWyWlsiYq4vw8obtMosCFQJ5T4EN
VCmI/hkQsfKHS60GFIBRkWJ2OnhnwluVTmfalH7RL3u4BPSJhT28eXz7SMV1zHM1
poGl41XMHcGK4cMZZgvzUDUPtFdcip+WTVHrHVXm5b/SL7KttzKiEgC3neXlnWOJ
OWiytmCVn53p5J6HSEKnMhP5zk2V9cHphnVcX41kKNGifzoZwnJgDO6ET7wb9nsu
xKzjNowmqyDukqjh/CTJBuxNhdzfUsMDxjVkuciq0FCI05dPdOm8CEFAgRG/L1kX
2pG+sMoUZ8Viiw9lNAvSW136uMkM7zp7TkBtVtw24l9mX786qOr9kATeoMM+zB5x
sP0jnwOJMzIco6N7GolI0nl1yqefcHdKOh0FaJMsc17nOMKGwIGgQkOyycP6JMJj
sAGIGQ2jumzVic2LOrhkR35qOU8OFTmjWsrOjflhkkt7si1j0OQokRzZX81lUzk+
ogtKiAsFCxT4ELKorEqZSRYZXK6/ccwmIK3Op7F6llCPb9RSspe7C2xW/KChtt4r
O65RYF57ub7r4kjEkbTSj90iRMW/Qm6rs8fP/bG8YGPQjPkRDurnAbLxJey+m0ij
t/Rx5iWtadPo3QASNMOUgVqTL8vbpCdCwRoLAdZhhDhsSaZeSGU32Iaw6Gl53x7M
qlo2kRXTUvtp4gIa3WeGyCsXZoepPzspKK9RxNNmPDouI8mlrdZkEA3FBKImg5ws
49i7HXAB2C58QY+nqm1SVnVppf3OuAjcKAZiJS+FazhkKkqMzFdlBDSfJ8H+cVym
1rFTrzqYHNILdO+a2kiM+iqScGQL93pHFK4gCLd4/Fu5jfTkZGf5Gp6AO4ntLbaY
Plh7UW6AKcSgB6gh2kUzODAFU0bPKPvMFKtWdgFi5rYZyVCVI8+HSgW8zFQkEjsY
6GPvsKT+IedSninoCcyf3oaqdWVa/oYyUo/uHo4KHQGPaSkwu9bhmkUc2+jBX0su
Px2B416ndvLjfrrFmRaxlO0gWksGGh3iipEkRXmsOKcWgiElt4sca4aqjxZTqUCC
pmRjie6ltj69FPsNPCyp0w+EDPDUrjSc9YvaJbcARNjmbF/7vw7tqUVcAZMga+GL
PxTII7r2IWnisyIE0dJDap08akLuhPGwWDQQTa0u+GWdbW6AbmyG7W1SEBAtpXkl
Jt3clhauHaCmTNZk3sEvFWLCsWnev8WkMRK9Qr6W3qe2bRHUVQ6opiFkmSwwYT6u
zyBfR7NDH4JiqZGMEQh1dNOVxbycu5evV/Mz9UE69w+8ZPNv0vJ1ObYejAnOyP2H
5DN+aevW2G/oLoHeP0LJ16KgdzITaLRMFPiEeSw1gsNepLiYJEXPJC8UsbUUDFIB
RMYaex+zXKK6RmwQ7NhvlfcQYiik3BPBRSMtj0hBqfTSLkWuOVGx1xxL4/CMFCAZ
RGiZwxxJJ+SLfJCZk3stfjAUHRVJtOh9VoIvZxz6IIILpjUlubYBN80ioPSadk93
va/zZL1oJDBVHYJaDsVytGWI+JqJ1GF7+IJrfWi63EyXecwcjRea+HPq+wU7KQoG
/EblVDXtn/cJJ1gbXWn5Lpwc6PA9jMIBNrMhGztMly6oPHuzxkZr+zW7WUPV2t1t
n/PkzxwESD/Q7GtAR95ysNppnQbDGSAp9hrye0G5OA14xcR7grgCHe+kNXpYjS76
SLRF4tpyIGLDSJgsExA1M0wJrM3Y+G8ftGCVPcVlvnCVQW+KXGtjaLY0sss1GC1W
8zfc+8DRDNBHv7OziSDB3PlYc62VtDSCyUMqSJh46oHZPg8EIjxq8J55cyBgU+jY
A8Ax8Pxrw/YqKOThTE+65Ct/16D9d0oQdsDPnubOAbk2p4ewTxWtml+b2jzjqwAy
ZPLz+OuzhSJlJ7LRuKhdoXoscysHuES5LyXJZZ2SxxGjugJMV7H6CfFTezPssMDD
G4/gMFKw8t6m/lQqtXudbxJ+zs73h743Q7s5ladNGhbWt561nHhx/O0RRj5wUbW9
umdANqY+V/I7EqP6ciFIXVarZHEkIKvr7ZTbCl9hGBySTD6y18U/iEm5JdFBgYrh
tJA2893E4XzoB2GsRkSLwv/0cNou9FcH+uHsg1cpq/6m/9SmF3D4EQLsLxKqirae
MkNDdJYc1u5lsDjf87SCPP6dI1IHSLYz3lU9GaH0KcA8B51CKFHr8Ie1uXHjWVBD
VRZ95WDEBEmO+GKxIUnG6DQeFKzDZZUU08AP7Yk0+1aQ6IySUCVj72GUPIug4EGY
v2nXGQPHuEf5ttosW55lnxxy+3lD+TforuIfZ1q9uumzMyTNRLIUoZlhgxD+1Yqy
NFxG8yGMp8EQ/4WNg176PN0P54gutZhx5DH2GfM3y7TH/aTkW5B/N6evV6HY/HWD
+Qtm+fkH4r6AYcXrKd/egMAYvK4eNUEtzjRYjxYf6NtfMtRrhk4EfsPN2lzn1HOv
Eaor1X1m7kDhFv2albp0IiK4sk25rvk5JZOy4crUFq9EO95vT6n7dI9o6TtHBAkl
Z0vttVnYnvKIX3JXSgsp2MLwvTGEJ2fZmcQ5SKZy2qBLNQZK35tKim7+oT+a30Q/
9BdeeoNAhVEUgL555O3VHi+RmcmzhO636/zyQMCsAEEQxzaPPHQLVw9xeaGqhU64
+kOYV21keTClHv71pr1AUy3ErvBoOzmkToSNsmTHN8NBtnUQqrft5vMnv2mEf1dY
AfHkem0MPMNwfPxBv98xVNQ0UXOgY/Kw7pZQbTaRn2fvvub7zFfJ3QkIsHG2TGXi
gHZUaeGSHMzimQIMFKSTSjVA1NS+1F7F+UBAnOLbCoU4+JVDtvowgidzpJP/wroi
s3WHCCLPsegEBCziCFtkMfid1z8NhQyDCxGPnqwsdFAz3YIen4iVnsx08H+yUuN6
F9q2nFDcR8Cw9uN5q/FlLFjNCSTfjyuS7RwVTKUlfU3w+eLmOqiygWi3jrA8U6oO
WUSnd43BDTBSpmahHkCpJ0/BkH8GTyXJ7kATt7xoKfGwVPDskKg/TpjmQ9gwFNMx
8kKda5324TLeUI2GPvBpQoZpkh82pqvlTa7aChgIskMCwgChdudsry7jyUic18zs
mvCwdarrQ8P/9G4yXRLh7jspfjDCIDwMAbiLASX/0m/xvsV0lsCi47wWewJQbimO
vcCHkCxrFpd09QAhBCxV+UnbHiHYA5o8wGLMATTQaZkd7o6bnUMDjRSZmxgri/QX
+RrbdM39LpBxsW+QMJ11tREa//rP9Es4Ef3EOVDcrn+mmYCBmcO0z8MghjkQVSJ7
cIreFmqvF0oICTEgcQO4gQGJAZrzkaLxE+hhW3RYMY71NiQ6L43b7FiTaJ2bMQd8
ZRR+xQKtAlG7CRbr3AU5xELYCqas0gjHlE1ViFavkIF0/fH+XhM/chkz7ZiFE6ag
w+QFMCI45DsVzEcsPrL9sfPPN6T3BB22nN77brWBfw8ieEo8vJKOHPUDXLYX7YPK
gTrSoo/XT4nk3ZJGzXjbYd+PxXSVkYKUOmB39hWyGH37r/8In/i5WT8QpZA40GOE
kiYql+xysLkgKYbAqNs/T5tlvj0pAr9rkbZHP0ltMio6JHADli3hvpA6hszfDWCl
LAEzUJvTr0bpmVDQEZBVt479OHF1bnd4Sraq9DEQ0p2xKIddZuVw1sB6a0hAHWEe
NEcDzc1qo4XhHx3AEnU6kSLFphzF3xiO16Me4aj/2Z7hncz3QMTfTQT1dvqtoRn+
s1KqW35x6gFs8MrIOAPXwaEWwGBrn/r8F+5M1r8W5v62tIwM6TpGkJUNkPamQhk2
TsZbma9vSCYIgMJHy0V447+k0Jn+zuGnNtZcxHzhwkf+yoiptbxDIjVZMEZtwxHC
zHmAURECDcWxAtPA7T7ejF1zMXEKOFtiSXTr0i4qmvg4kk5YPpAI+X4ipB5Bibja
Cun2C7YqxLaeNU/7RwuuxjGnKlZ74GakPbXnT5ZKvZ3WnJCMVc0fHJSKkfeKsU0m
yYoYbOLsxhPV05oPrh2t4kOiWFloaDazayRk5TZomrExhPWOnJN2G2BZA0kwnzWd
608v/XhLNbSHmvNbPILLOfECV56RQ39lgcimpgfCQlMOuFtHPrccFicR/R5ZtW5u
bnNKwavmfobDtcK2RWL047YQelN5tBeH8GMTpsnh5tG4SvKtabNMqc9R3uoZ3aFt
SSQs5LVfggQahJ6D9+H1foauNkW5zwYjuJHGWoNyNx9qoNydhWhv3qnTyEZtwoET
axb+uKyv2JGxtFV13lOjPDub9uesZQ6dTcPDYwiB6daONftzaAv6QUTLrjifUZQp
uawL7WAdLZ1mnd9YlM1HNzwGR/SqqVBnDSF7t+laHBU9o7aFbnMpG8uV+i8nGqXG
3M9SQWCMcXtSS+kE1g9m5Ko0zqDIFZPCRDgCNwkvYhx3qgcELf26hRjIyYmp4cl8
IU+H2bYWAaHQDGNA+izRmkRTMA8mFAUwoUvuL7oq/07buYODsgPBLfiXuxx1QpYf
yD/UBfyXsFH2WEub95nATeMs80Ca8jNWs33ZlQxaTL58l6jyJwIvwLC+q+D3CnWH
3GE5XkCw23Sw88RHOTf5WQePoNoK7fcw3fqY6Stt1lW8+t8NK8uyD/TyObGdsD48
FEo/RBBhTbdNtx3LEjFWU/1GohPH4SwTrxfM/H2EXM5ip0Cxptc6JAqC1BxNv0JJ
vPK51i+Y4GCS2Xh8ZNpcH4VHNbIS3MnuCwqRE8+Buf8zt6532FvJE4fgCLwP1kIT
TVxQpD1T8unuw20hd0dvwYnNGFo5yJVmepBmKEHEp3ZqTF5CLShSulmlkBVcSw3L
XKqAbq4JdG3nWE0XY/VZsbDGnrZ9XDr9kO0jrgFtg3FNIJXs2igPED3i+cGsH/je
YUgEiL+5yUEhLTsAUa0dib8E9GxOuqGnNjnldCt8dp+hgirmYV93N7vVhe3XTRLK
y4/3kSKkW8VCqa9h5KUstotV2pKV34oHB01yqPz8qi4mOM7KE3GK2ZVFTZLCOXz7
sXh/MbFsQU4zy4v4dB4xqVq2LbgYK64V07LUBWfZz3kY9ElfClvJLtH5wW+Z2GZX
O2gYJafhSuulRlf1SifWr4oevqExyqzVUq06EwLF9PGfKAbYwRzq/pgi+JoNt0md
jmK/+rWXpSgSLpFWKT+EteI3CmbEtYCf7MC9TzCze3KVHIUItk0UhlrvDJzNchKv
g4BZcFOWDedPRKUkTFpM/AvZ6J9U9VUkgPQWAcVOQKT/ZNroxNFrH4F8p0lbneCf
V08x8IbzWtyEeSOu0FA+59cNAWZxngewwD9iXaVzH52YRaD7dRDGIe7fp/AC8IUM
YKcH83OdW7XAOhxPVd3yAxsveLFhxrYzNLsvIG3M7alvsuZ0NAwDc696NCZIUpZS
VHdQLqqL4/qU+ghTpHqVrIHM5+9xT1Gq7S0EdZf8UfqmIkkNtICemDprvak/bCse
VfkEU6rNnhB8yDlftnAmXbx1SlcCy4VzX5rex10z81zyTxykS5wXbJEttPlZ1w5t
11AtqAJlebPrg02yHZmeWfNHxleJQofIZzpcWl/CLOrb3DDCUWVoFCxoR947mCxR
wF4Y7c5ishyPZVB8FV9dz+IWWVlwrUzBqCTsw4cl5XmjUHb38/vigOSYjJmUfK1h
/XV8ddEp45ZprTPzCNSNvov936lcikee911j3WIFcmUy+bjnDvKkpaQOgeiEt5Ko
p4JI8ZcDqlSLSIi/5vDgonnfd9wptyfdeSDBGHR3uQ/2O7hJhGRBzYyYyd0/1Ahj
Qme9e1UK79d24JNDoXzt0jKCTs398QxXB1IUN/6Fqx/x3lxDA5FhtnuDrcFuG4mE
6IH5LfDsweSi1oqCHyBG4a02gSJFyeEL1vdEYo7zZ7eUrWiN4MmJaN1x6p7BWbFW
JHiugjisoUT61HRF20moSZLuRxCygXIT1/JjVnwuPUzIB4ijIrCx0eJjrGG8gEMH
Xf/8IUL+h2b+XV19wnghe/8pau3Y6+AuzTc91SCThz6utOmBusTC+D/GmJFxDwPC
6JHRkQcZeU7A7caKUBOfcNF6443vUZ/HdIOiFnoRpsaZT/urYj9gxjKp2jP2lu+S
kbiWB50xN/rRzGt4m8SM5lYluRLyuEU4CTMQ5rvEZkFxCXXJSVsGqTPxp0vyXiCR
/Jkm4x3HtCuQVj32Rn26AQMvNrEavBOTA7XDK+jKYw3Ttr2kiOtEIaQ9uUHUz7k2
sXGrKPwrqbFz+jCmgLWnrFMcoH8PkSYwS27ukA/kyPgNyk/5QU02zsnttq3jsmof
p86PoPn2kgPwsMltqiGE4mmil7Aky56l06OEpuXY4uPSk/nV79sZ88ZdtA+j3JT2
KjRkXmyPAoqQajrbG84bai0f0CWDgY1j1g25PB9VzON9WoYbcggRD/8p9/BBW4vq
bu5uECrodYG0odnxb5oSIH7/J/Qnx68DJUE0KNS6bSQ3Q5HGykQ+KFzV+VEbAf2T
kQWlW9+VVYnHQMIPu2etqRs5sKjUGR61COWJckCQKwGmxMjuNyb6kPvKkPhJG4Tp
hW9LHwDMpthXEdZdEWrN0oBfcBCqR986uVmeKlcgjlM//G4tvzDBU/XsCajVgkpr
PH66P8Vf7NHjdXMqW/Fn00wZSK/3muYQKqHcCx3axCs3ZQ5kKYyN+/TgH6CnwfRE
LWqTEBqnRWSp7XnKFy6ajWFi/gtI45j/zEVs0Z2vrAsBqHGksJM8349Vu/IAsZvx
XJgxRPm8cU9F6qa4eKweUNOfb+sq0WOHCQis6yFjMcOU6HSd4wGf/qTXpyRjYtR6
1apMHL+RklggBlbjAzCHA3H2vPr+Fzwlwky5eRUx9n2B4SViePcc5xp1rio7i7he
/bIJMuW0kPGaHlQ8pa3MpG0FOXtLR6iCb8gMr2ZAZw6r5rXqiAiIA8ThbQ2VRvhh
NU4BrF32+4IfxRVLfxA3MkSfxLS/A1zR0GyNgT0RepDs8KQZZuRZcFTjCct9S0Kx
xuPYGHRk3KULEz6WuaPvV0tt+91e0zlmmapVZHuqBE2fo58Lj6bw9CJK2PJLgVKR
FgrYBUvTsOUk3XSb5AetaQloKUwrRESr9oa9zPJyoTmAFJNDKplAejJ0JNSVb9qm
ubaNY1lH3N5Qs15K+Ld2Vt21++qEzt6KsmMIqTAM1tSrVweXKumMVXV9vN3pdIH1
RV1AfudvAJbpa3RvnxrgSxsv7RoRNxxP/xgDcpCHUxdT81K0SiAzkZLV/quQCvBk
kPpxFOFOZWDIFD1zu0QDFoidxU2cm/7xUYBAablndnQOHpLTryAMANN/FuYuGz4L
xKbCGT1iE3vpSiD+5NZlPFe+5FmbYJjGkjMBxQyEAIYAjOm+/EFsQfvuYBOoF/SN
IIeTADxHtErSPetWWi0yyCUiktM1UU/cQQoW/FPMJWRgiqKhHF9lQlReaM4U+/ic
pW5vdLzfH4VEYEO17sXrgS4FAQ4mibO5XXl1Lu6GrOABEMPNEjPIRegG1b80FJBd
FsT0kPyxfkijMghMm6VBiza39etbPS+FZlvoawA19OWMXVpCzEEvYSFIttKCPzm6
G5eXCbXRxEmmtVl+5suDcO1MStDTWT/plLgZxqIjforZJ39k3LoAjihr/P8lkqgM
qpNxYk07bbh5YpITZtGTTyUtO2MYkfsKMCYwkgPQtVLZygrsXz7oAFkjVbTqNdsD
W3rCQEszTdD3m6oSpAY0AoellscSgJjxJkHhieM73c/mknPi7owlor1k4BgNmdp7
84J+Ijv6liJ0PhKv6sbtgYIk+RsYYEEzyIXiy2surM3YGbG0rZeAfSXzbmRdhA6v
fBfBumEcsm9KNPJkxCoMFfwzKuZw0dQaYT/BvSSiO3lgazCIh2tCGh1NQgL3vz2p
XWJb8Egj6EtoZRNeG98Ym33eaXVQIbrQrKuRdQePLZuY4svKb7zcet8CV45hfbUR
Hs7KXHIpHvX4j8ZGmhuPuk6qgSosylh0wJXiQrnhZ/FA76ipp5DrQricFW010MVk
t0xaO57GnQa0YGCZsAAeH5zgd6zC5arf6LU1XqZ/1NbijQ88KVUAQ3nsfqza5I9J
K9+UQkCE4pf7gqlxYrQOrvIH84oQ9FopwuB4w+rpYvHFHKf2LnB5Eu76YaVlRnjE
TUzGLDHBYBrBYOdpAQiIeq9+KvaTxnHvZ3kiCFfh9SZwSv+vtW/CY0Rlx+/sNdn1
B6nBzHUHrYgMWh3WmcaxEZ++TDOzL6MM0IF5QDfeFPw5tB7z4cQXjRD6za0pyu9K
/x6/jQbJxjifRAvsgEPqL9xqsyvMSFczDyhWaVN8KKdXa7uBqNiUkj0AU1+IUMkg
/QBTRj2anuODtaDOysr3SX/6eh88dfYNLSaGg1+iUKZCPpkyqPnzyliL+eSCstE5
QdAABq0wq0tZuX26mhCXY091bxSk5r+l6lhOEwblVA6q0wplQs1/GDY+79zp8GoB
5CQ1Ku3XhuUCpUjYrs8/Z3jN7I81QOkESCPzlbPddKxsswOV/4zAwxGQ5TWz+RXC
pJNWX5RJQFVfwlx9voa47kfoylydZ3btOLG9uXna8BZvcB8kJlEvtuaFG0xpnZ4C
5IDwGyZAA16V0fqMjSbLLt0cKxzrJ4v5wSA9zFJwQPYIYambbAozoAoYTEaM1Qeu
B5y2a9AE6n/Eu4PFM0HIi8XG5Rpx25k1FCsQ7oErSgW4lAnIhIfwdE/zw9QJlIhU
dkhGbxbRFwFl6nY0/lfUDhZxih+7aeIpL1HGKPJ5ALKvxoFxGsGGwpDSvGGWiJbn
xTI7vNZgwN8TSJNBJq8n7/CaR8mrW88KXl0InMTN8o9XTcm1xd5C4t21YD2kR4tI
FuW6YS3iKwLFmg2sPw0cX0G0PJXD5LaqPvBKpQ1FdxY48TpRSEZQpqG8R4EXSVqg
xPCSIk9sstTcfySftrteaba5NWgT54qXiopr8DVt56vKIW+pTkL2RfK4UdsuHIFa
rwGpeDCW9gdFoTZzI2WvEzE900miY2em+13jo7+ci8udNsPDzSUB0edwC0ekrbTo
By4Ut+5TwlS32NgvDJHi5jFzCzUjPzwgeGnZH3u31Spqm/sm/DqexB1KGUdTeE7r
QjqkZicQ+fhuod3fXU0kwlSwH/RMqc6MHSnbvKOd5LK/9xWK5ZwOBfrrNMzqkAvX
4HmfTlu0196tKTGJo5yzlsDZFdIFeKaOxgnIBonLbJzuMYX317upbKfQe/zCUTzV
eDJLzEMumbt8GA604M4QwcA34Af5OBFXa68Ql17ZelrgHajDbpMWPR/3RrgwBUsB
KwnFC9vtqdwmFLTKYipH/Fet7C99/fs83WY6MQ3NzXVrOahzuR5oX11dUrLOXZQe
zOs8WtERbBp4UmOeIWaMknnk7gjLYT5AP6hqVLr7EHVhEmeErGmlTXGmtQqMljAa
6tpIVtAaKByJ2OEhG14Ig3+zMkBwQifvslIvwnOgHwJopBt0/mnokeCtuWQDBXZL
2ofWZVpMBBcVTRINHkYgAR0FS3AbxV+c2+QtartQ5ljMfQ/slqUukMRU1QjA95zv
8ZY/pgc0/o3jPdmwLBm5qrgNBadr7FKupcOh+OoTfnKzsKIEkD/kDHWCrQTbnGMg
rAL00LrlR47YBEAFfalha8ZOqFD4bUfBcd1SQQ9og0vFMbFW8d7nxpWnqW2URPzf
im3BOcct8yUTNTRTKZ6wX8D6fg29b+sqcyq9n236NScpNjoaEi+1arkAEesW3+ww
r00VKW2CiRJiL4DcjMRXve7Lk9g+x6sHwxmXeYUB0xyxQhEmDMxFELWXsIHPyNIj
VFhmGC848ykBo5BxuWkgHPwYnNd7GpdR3Vh8VW505TSkvydW8mFrKfGESg5FyVQW
llB+HMYFCW4jq47D1fDza/kO6aJ6GSp6Bz5gB/iuJFtblFzoNqFMY7puAK6CtH9E
BwSki5rrCKEagxSKqtdM/OicXJ0Jo0lVUq2hzO186G6zVHQbOM+Q30UYR9RCWnDn
4yChot65WiMCeHiT2oSQCpqj/WDgXzSRmLz0f/BJ5pAdWnQ9KzSsAoCd8MRJrz9O
o4/2banpUEn855HYZmNbVK+D8M/eWtJNGwyEIbcknH+jbRDh6+9vhszQf1/aMRRR
d0KicEx0LqD6HPDEJY+qhFOq7TjE42MeWLH+Nl6PJSSRJ7coAWVQMqjjC+11nM6N
cuHnereOI1MEmqUvl7xkDN59+5edBH9KMHQ+v4UGQ1ZmncAUDNHQOi1WPAICwd6g
J2YzUemIAunYbi7ko5jeRJpIpQYS/W8FjyngOekpkxjWcqUm1SA+Bv/Uiglpxunb
3cjOCGuDcxECHRh74PMaEXC1ZfBB7LT2HQS6ybvWaHHITtyyUahDl7aarSFl8sxP
IENT5NKHRDO4ZH61IaT9iiN6XlWnRDLcmf3Gv38Xt2fKZFhVH+0Y6UIO8TqgSNUz
E1b9+NFiu+TDXyxa7Uok/xFoiiXbl9GgD5PJL+uRiXWRUPIdlRFe+4/LyLqWYSJb
2bnSkowfQeKmf6cvmHarEsC5SbhsIYafka8xwjwSyLLFc9waCIRa9i8zMY+scoFI
xjASP67Xl10ljj0+M9oDdleR87aSEa0gocG3g59BmGMXRmOa5iAT9jbKaX7O2hgS
m2I2aVCV4abqHPd+UKlK/n9dPNipjKBP92/Jk00/gQuN+jbaLycyFb0+KmDN3iOq
vR+cfAlWYRvNqpYKmf+HS0lcX9xcer5jJAzxfpjx/qvu1hwTYb/HI2CbxGBdWTUa
TV5iPTUtzw4+Eh0gHg2Jd5KsjhJ0SVO9dHKKCNPDYNVTAF0YtOPgSd/JGIs8mA8d
iZCaULBbpbuix0y8l6sMIP/WMFnPwmEuNj/AQCXbuFlKGUIQ0oIX6YuCuK2U9fhH
m/XUKX4Ux6AXVQsXHBriu15G8hVGrxMdImh59bAZHbD3FAmrDLvSRA3aVbs3IG3I
DqJRWlKJNrbb4PlHPUHfsFSwQWe1rmEtHBnfc+mMFc206hm3IHTodidX0kEQEaN0
1AjB8e85ooB5Tud7113+SATdQSPdP32SPGxYJmd3yc2mNaCVX5uywovfsYKk0GW3
oQGpIwzPS1hqdGakM398bU24z6Cd0NDKomMvygUlbnlQuU3i2Lhxp7z2Tuga39J1
8yS5yAsCrRQPfnxW5143q5B+2dGk4ccinP/f0FR3OZr0df5PgAj4gRIo9pNdOsCD
9e+fzzQvOwsGQ5T5NjWwPcyESlysps/2Hl1up7hoa2g8fTD1ptswK/yIQIzNDaii
fChseVmvqBr0nJBXBjf5EfTVjUejCyp8fNlYdiYe3v+ZoK4Bkqrr8H5p1AFcXFy+
JAPZo2kOBusD8IpIfXXCwwhWYAAdcbb1sXHDp1Ycfdulvpxs38jKmxEJi+2kWqSZ
1N2lsvWuqGeqtnVwIkzv1xfqZ36im3k/rv2NuRfLnSPdwoEV8xtPY4S8FoJxZO34
zp7VQO5s/xHRdCG5ocFfabR1357Nlu93/416pyqSXzUNKo4ftG0TVdsXFJb/L9Dh
S2MPhTIP5HuKY7lAEih5pIySIj8THzP9FsjOt4QyarMz5RiR6tYiHiW1Jy13uShu
oDEAk3Hng/YS+RUJdHWjcisi/eGxJiNcHr3A/DbRrkOxv8bphmATAIM0is7LwDBg
xccb8MXpQxSKf4NQ1xGxiQS5CYLmOTd5g+4/9fuqTXSEXnV6jegHgqLIYntwAgtV
HJ2hlFo3zQZRIYKi/tZRDZQnpg5GxJ/JPkF4aroFPx68tq3WMVuIBVhgE2nVwCqC
8Ijfx7xdctdd8+XvIuW47sMefsC034ZfApP3baI8LwKP02NIKVAQGYkrj8HLVyd3
rDxinmDF6zwqWvGe2r5QngUTa8quxCEn6PqcXhVit6x+aPbnhITpdjpBLJR5EvDo
8uDIEI00J5qqKnm/COufpsRTYrdSDrKG4NqcHU6nKa026B5XO8aNSXI8byLw2FLQ
D/Sn+0/etLHjYUQq/KuU20o7ca1zYY579vrUz9pPPYB6V35np/HdcxoC+LqiD5J0
Pdk5kkvoz9fT5fMu5phXImLTYNRExy/Bvdsjf1U+FawBbMB9oZb2KTXNC9w2cnA8
jPhrcy5kPKeUN29NyaWtI5gBHEDZu8vo5Ct3nMU72WPWMpMvbsszTlqmKSraO23i
fL5Z9A9Hf86NrOL5IsL6Chh9VrKinCwto/cub0135+dFLhC+jF7SD9hS4Be70mdj
4BRom42Y9rcD0aS7Y6NjljFvq+iHhTUJZeEGyDjcCXcoUPgzHxHD+01aNQp67b4V
Zgu7luEBnXLQOZGdPNbcU79ppcrgv9k/i8jJ4kQeficLkVk3JEbzFMl0CYg2iftb
mNfp3RHwIH1m7gbQx7oJ+Z+hoolYy4xhCJPYJFr3kEFaOTLNC7QMcn4rC8T8qKWg
ToR0V+1LsOrpGZvrFS6SLIhxt2xqTe8oAaiKc8noftaTHDTdwicK1fpScsr5Vuue
hyVeX0NQElMRAa2/g4q9onxL7qphBhazFJ5FeKCXmQeFwbZFUt83xPqVQA/f15wv
5IFPiE6ew3C7+h+bC2mrqVNiMynFvy2rmHISS1apHpX109986qO7DSOdG8lYZjAy
tvXCy+BsXtdt6lAMFx14IpLizklTTZEy5vjsW7obxE9HSnrv8K1OgEMLuapOc5HH
3M9eRsNl9BP4lu6m+jeNotjCKmIUypiAtvC+7lwB7wfz3LQUGbOPq1TFWe6c6uK/
Gg/Im67NT+KjFhIsC/n1AMhDUedm7lcNW6AigO10KvzwP+Fafj3wJsURa8u9RWVm
e9uZhgMmeYA6lM5sLm3mmOMq7C5FtT0m0L6uU/dLCsQESVi8jl1PLBpmtYUVWZE+
eInGiDju9WTMldEYOywYR80uNKKJGVaklXDyun6OU+zKnaU4h/Iajv4Ev2C8F0WX
RK9UQP6MquMCpQARQ6y8T22cJxVKHSlEazIC3UlkhZxPgLPagbUCkpGSA9tTZZyC
jk2801F0JQZ7fe3sSGH0Y5z0L/bfPmko0q7x2PjUL8SIzk4e3C7CbtLZlye790Dl
2QIunlhvCYH0rz9gAJFb5xfeQBNiOvtwvgT4y5UxiTWlhxeWianaoz7CFLcoza+3
YCqUeeA8NXNzes2BLr8u9dgW6F8t7KLOu6H8UKflzqVAKgdtHIGRf9d18YgiNf0N
QAfN6OYsDfanDO3mpdtELpDV3/yXWCBlzzaImfNvxYw4IOXElCe51pDugLILkgjS
f13qnXUw+F03uKi5qw2+2ombUXynJf+RoU6yNktjMjGG6ev14b7B8fcslpDZPR4C
r5MpbPjmXuokkgAMj7LyFJUtig8/aMClByhqCRUhC9LDTm3zDda0ewS0yE+od7Sq
OFmVj/wAuHgGM1hTlCWpMRj5spPt3dSiZzC7a8/UoRGYYe+xV0ciNEzlXsrSZblN
VNbY3W3O+5xQfcLR0TL3wC465Z/vTmtjlpurtvvHtX6x78j6EObgtdolKGGI52qm
Edv7BRuJjAPj6XTwT8iEfpcIx8mJ6iO6Q9f0d1YW9jtcz1se30KODnxLwbyzj5qI
MEo/Nwi5TVYgQlwbBupmT9UGBZbG7PAJ35Y+isEjrVPna6HcRMoqHxWB/SqxuVit
XIpe0eZM1bVngk/rzYsapHvitxNssEzqLot9Qkfl1rF4f1B8b6xsFEE7cp17WKWe
Kco619hOmPgMGSYX3QMN/EO1djHIt9UXWltozy3VDXWQfmXYZSrUTpEhZopblzgC
OQANieXh9w8oBOjQgTLqGql4vFS2BzJOyj10Y1LqkO9l0GAZUvMENgLarHcxBGYJ
2mkekaRs2v7/cDTwPaRPYeaOEsVJvkv+CNGn8qpqBuZNDQ4EScckjqC2Uf3kD2cz
Nsin9ylAzn0cFQJAmEVCI4uin8MEMZbdI0HkWpjEPEXq+nRZQ9YQZlHmLK9OYSN/
SUI/1KNl2WUX4GDJ31ozbzevr/VQKawfOfzzx/qWM0NJ9FfVF+WP38EPsHlQu6V5
pp89OFS6guLdgLi/wnkrKK3npirqX2zt+BF3t4RBmb2VV+JgJjdElHe7o6ruPubV
77ByHmZlDXscROCRZmF+MhuP81AU1UWEJ+r3jIZRZCIB1D9ZQTkINNPWWH1ROpOY
Q8PptdqR6YfU+8f7CvXedUkOBPvucluT12vSw6kzxmc8suP70srMQtD+OGCVeW5x
6s65YchhZz901X3cLQeKLXhmnp14uuUlvzUKYPPFIyxE0Fz7FiN8YQAT4nD2VsU3
NSGTUlYuACwV5MgCQSFuclNjq4ZBYMAVew8ucc1oPZ3JX23NJvwi1xsDvAOomzLV
nOH7Ze7CwqyeJLkmi0adt4HPNh3yHTb00pqa2GJXZTu7GzYKeaTmu3vdOMuYN3xb
gVHQsgGnXCIoc5LrXYgrpoFyjXXEsn0TeB9aAlPKAGOdJ974cNGun7gkGfN054fn
+w6fR5s/6iM1m8LJefTDL1yiK/L2vQhBYi2lx79ZD10B+s7RNmXTydzfi+g9k2Iq
GnhXj1S2lxyocHTC0HYIsci7SAXG9CRuypZZ3YFTMQbfHCBb5wFaZSKwoD3sjTh/
ppKJZH05NTb6WQsf+4vQwJdxvpKXUTqCSRcRe1ghP0q9NzPtUUEjZey/Q+WWiVqj
D4HuPob2ZOYizemArqr3Urc2Njiv4QHVj+l7/jCvZweURXct1uoK9W6Fj7Z0/Cif
AMVwwPYuAhMnf21uX21eZjzEyYRL5KUVSFAVIxpZq4PQipis60n6nZlsM5usAZjc
RNqjSCv8pwUzqJn0Dr0lE5Qg6YpQkmPCQPZNbcmjEX7geGM043IDDxGcKF+CKKXu
xU29DHOEqsU+jYttSwd5sRnN0TkS+Ll34qHNmWQR2hoQk/vej8Z98W3+pm65tbxA
+IKkWBxDuzfYP93zs3rKG8cd6volfZ51K1CNgKfn4HB3yGKrq5Od51Hagf3a7jGk
eo9zWTR5atHsb6J3EWNDn1PAFig/TR9JZ7Y+5d/wvHfV+1eMCQGYO6siXqo2R7e7
atyxFY9NHEBRtKM4fiKL+wR+hL/+gmlAe3fPepTXjvUcSOfc7uLWX/EsNJRPTesR
ieKkKL1FGAhvIdgLoF3uRuSvCO5byIhIsFWfZetQ/0NrP2WFJpft14PxyOvKtv4y
dWpahatnVcz/4PfRxmyk0NlnQjluHMV0ksf3tVIEOsy9LQ0/czjbQxD7Wv0bR/5E
Lk6TlaR4ij7RZNRZFZ8dONWIPKC0e5JWlwjYVVP82cOVbyYR7biw3ehyJX8jlCsx
o+xb1WvP25hniUz/UvM75Q7k1j+CJQsEH2DvtHnH339a/0Jg+SuHafdJuTfa7WlB
3qsV+KXIiQAIH5aC3sPbSXQLgC9bfnI4Vr54QJmHfGDOC/maEOjvmF06UqYqRwnb
tEWdxj2iOeDJtkV0QtwYeNQVCMoylsPWpazdw9DAW4m2ceg2ljhe7ppLGQ0tdpbZ
MS16cEdCnFEoKLlmcPydS1OmlewldAeh3tLz1RJKEBGQyRXQG4omIrM4yUU6bqsO
JyCwFbrIEHsvJC7fo5h6idXZE7NQeV85wv56uryrzQGJbO3ZcLnww9G13a5dUM/9
lX/EsKibzuWlkrkGzmtvWnay02QVDEOu1WsSCkZTaQ3duxkF1lEjrqXMDFu/65gm
bmfwNsvkjH2jZbSZNieZJXXDhRPi+fsM4A3UHFRAaoSfF45iSEvbljYVdmmDEoRi
y3wbgLm2ubGRUySNs/Tj76aRRIjXc74NaFRlWYsjXC2/uHzwkrTdSysu24eowc1I
IBCtX611YdlYS202eeE7qWoEUuLtovCgyPWCTDUGeWCJjDA9aG9IDRZxQyU5zLFa
rsa5woHIQEAdMUKL8p88KNAR9JcGUGdG4ef0GhtmdAgaaWFy5lKdYVv86uE1tkTl
rpF3kzGImDdsclV3216YdXZboRiq1xaBs4W3EP6xc/PqUSHAqwXwB1wBaqSK8pT5
oQpEnrIaVjfomHS0fwl5yrdE/JfrQb0v/ND0PEJ0v7YWULCZDrMeIc63xWKepO5z
m/4KfBzHQkUxcoyAwQlM+RBCVZNb79BIW1Y3M71Y2coBSyRMSvIdeqnC96OBeDES
cAXXFMx/Y+OWlgKQzY2JhrIKRwi9fWf09TcKnx9Rvn5GRrRqHK42DIl1euFdGHd+
eW19cxkUlHZ3bJJQc99Lqvu/WjBiU14mClYJ3hVTt3f/i2zligFxdrn+NWIfl34P
1euWXOLlm4ZpraEcEwm9QSZp/9ckoq26PHtGRzI9R2+vif3GPi0ZRj/R2/ZnWggn
NNi0Ep6gDneGXOBSmETmFLdNaPUj3NNTRdNOIQ2mW/j1MBZ1jmsOVhNmaQjkJbwG
RrZdv71HJtsuUwIrXiI8hCqo8ruBYUJ9Y1GuIBDpFtdAgtWih9kzRq2kzMSup31j
ed8FOHhTrGtXqY66YgJirQ0mm0voYpcl9tgVn520Wr7c/RpWR2rzbnCiqfKJCkJ1
iuYTg9vsWpbdclbiTuvc7JkyFxiW9lHxBBQAf4XalYaiBXPXIEmilu4Zk8ELNXky
+w/8ucBoVqoVRI9n8gIBe2UkN00SGB3+e0doXMhjJXx8CDdnqcspB9/LrHgYfM+d
J8wny7L/k9qCRIbmeOBTMMOjPMSpc16YerJxm9vW5B7Wq30gHfwbYqzoqBNPdE9F
07xV4hvPkkOf1bMItSFwNM4LiDUMyBNyNaeajEqGXAUzuLjSWX0WN8qnxnkoE4fy
BLqp23Z+l4nQw+Pk8lZwVspjFhvuMBlcr/Lo/gGH6IiHldPskK8goau09xqlXweo
5sna4CMfEtwRgkdemry2fs0Z8V+h7VT41sqDGcfEEMwmYhAQDop0SOzeymvAiHbM
frT9UR32EodpoWp5ULsuqwND4KbgUmM24AA2IxKAXA1DVUZRU3kb7Ox9AjO9mh1S
CvrrkuZYhYx7fx5ke4fe5h0Y9uDfxjcux/vmC4gPs8sduZ8HvMRlcnoX69sazE/W
HVH2iGL+3vRK1gzJFxxV/5g2uEMjKEssSFezOrOPl4IuCovB1aCnHFVtleh7jzNM
DbXX4yrX7uInc59jD5bavBDkUnyatf8TJfcUjT1KWvqxI1skR61kdvTSHczhbKjF
9R8qJKM9fbIkQfUksYBFMnSDxiDt22Oo4+6XWizd2if5u7zhTJNGuSO0eGbPaZRZ
UfhpCOzAZy1GxPJ5jjS4YIoCct8Clm8celPuRLqFSkl8GvreG6esJg8s9nGYMDys
QHx+T/h06j6YjoqNyHOmvWnipfSWt2pH1T1g5u4PnAom9x5jPBwZmy170fsnOBqW
1NCUPP9qvoXLamg9lJeap/BBE0687UrB4m0NUb3f8lCkCUJEIjOFaAk/UytnXjgL
6C5hZqmV+MmNGLoTxvpLKd+4ThMqRSEBYYgvT8+mK8jnG9onRmClQdYd1Gt/GU+k
BiF5+9NN7gouAXr8eidK3d8rkGt9G2ihy5uIBsRAa+zsWHqkhF9upBPL3BT1ROFd
mFp5aqxsQdIpoyw6EUHETJDmRzOty7w9B2Yg40TzS7TJ18jhdh1sqH5gzTe2VkqZ
cjIyPICmXURzVQ0zmPGAMnvX+KuWCJgqRN5LQy2q1mr8VFA8j4wDBQhdGX3RonSj
Ztfl8WRsDyRcBINQuKlqA+3XxMKvW2r0XcgzxmDdj8KoPXDaZCZhdD9/NtOnzcVS
90asso/0NjX/GLFyMu7jYhjxWdHXnL79bgNw31Jnw1hoOfQLHm+dT9x7eBzzmlmY
eiznJ2pDc/OWoB9agkywqw9r/giO8kaiy/zAKuW/bOa2WBpSMGCBGnFow4TtTuoY
qlQFgbB3KVHankI6Z7Eo6Y5lh/5jXN9vR186LOj7UigRQ1MEiY5IRXZne4Wmzj4m
uVoRUoD5/u8UdYLRlJAcMR9rFRXtgnr3ovWWt6BMc978Al67OxWt6YZMv47SLlSb
BRLR2vsHyhbA+msMS1AHmHZ5n+kJMpVn+k75tO2oJr3JOsoFY1AeUlS4UxrU6K0d
bFhpR5SRHPvjaIAJovw1bTJg1h8SK6b/KVCTHN8YI58MrEZPBn7w4dk26D68/BGh
wl8WzfUZrQkBc38El0EGVjKNNAJN4RbEhuJVjG5hE3KJ8DEjBXAikOdib6eRibmS
40UM83xkzEMYgE4mJmSiyktvCG5BN+m7SORiK+S2iFczenyr25xSVEHodguX+Asy
hUBWD6pNYZo0aBxnvn5+lYPEcNjE1VXS0Pvs+W+PIkPyIqOzDZ29gLIlwDUcd7EY
1YdJD+Z6DiQOIjJl3W+u9KEiCpDHWGRyiLrzFwSUxKAS684yD5hlGwN34xkVv68p
8l8G/hpQlhryU+bBDpzCPbN4c+xpuMTQOqVyclHOhKGZ1IeRR4Z6wOYm9Mm7H7GK
OtN3CCLY3BK4bwSZdSCV1E5IDb0Tct3OLgQxdmNm7F3r4uApwL80ttLTvY4Y3anu
UZJ/k5GrWItYdL/Nwb5DThhmZ7MJDY/y6hpwZxkJJh83VVhQ883BF2DiZTabWnn6
RbyeN+jTyvvQOV1LBPTyaLaY5yH0N3kc/nCKAUAZy3ei1nt7E9pbI25pss+YAQXD
YNXYNf549j6OKZ5Sl+G9PHs2VMrLTSR3jOi2jU6Mk1VzXlSV2Ma0B8zYu92YL/cz
CuBhmnGLKTTPamMvmjG9q9t+1+Uc2hr7h9y4iDIIU+UtFJ2sDV4YPw/cHB+uacKc
LzOh4lKRRcDyCd267uI+rqlUqHhAr/eoJ0+dLOjWYIq++QrXnrVO6PRPtSo1WsMO
3gzqnbGtGlXujAG5v4SN0tFOA8al3E90fFuJrNFevgopLiDJ3DLbGD3klf9VfG5z
vHQzRVF9EpRRFToa2ZXbAy2xLvXyXx80GDTYs08tfzWmcHokFHp95M/SS5YbsvQw
w35ppR7ZJ8bE0lQMOPVF8ZRxx6hXz1fWEjADCCpll+ls7e+PMzsTG/AZ6isBIFrO
uRhps+MTxnJBTHOIBMSYqL3ww7uB3aaOPe1X8z56wshLuHUnjay1PcfX6vdSR7ij
eQQJehLbkcWCV1XIcQ+oIVmLRgv+QF7BpR8WovEOipHEvPHKeVj3yhSnAoW0piAL
dLI6PUEYPOc8L2Wl1JMlzcQaq2/DhpN8OBkxcy3mbr7GOmjKXYXZujshztqKtfL+
ZzZcyo88qs3jor6NjZHYMsLrBUL6M1k/E8QBTgZKVHz/gYAvcgU6xIdGlJQmxyan
tiVg3mWfoBimriMuGdNstn8SE7Zra23NvhLxPjHaqnuCzmUy/nwGdQMDaqmfV+ua
Xhgri+54Q2I+sL1yUcG7Z3YCCYpZIq0gM67j4vpkB+eaaL+4GrYFuVsC0WopVPYu
7aFrqSRzP3xZifoSx6sdHCMBknPVlyXx/M9Gx/eKtpWP9kbYi07ZhKjgj/L6uZts
FnKHYuaoxI7ganWehugH0VQ7A5lIkA8TqrSBQCuAaf5yxNAK1r5P3gzrBKNOSUw7
jCY15cut56TZYX/AICLtYcBG18v3fW+OmkE6gLJvGHMkLJyqxK0M9I7ixCyfcTII
N7+JZhc3kctNNMUKTVhRABrJiLUmhZDiKBnuAVRiy9+/O8VlTTPytmY75JWJXmhc
5K7t7JRScD13sm7mQeCzL5KdW/lP2A8DXCtNwqG8UNFGsswg38zJn+UlCbyM41FJ
ksg3/pnF0MNlF/RiLKUKGOsDSKFaBHiX3lCn/RgxfMT5pP7w0VjnWYaGrdzZ1Nax
zTF1o7gMncS5sTGfJebm8/V8ssVxvSpsHHP/c71NfiSK4Uw4FO12L2FfAFqE9Vib
LLJl3trRnvCB9DJ00kTnHjCU3SlDm5RoHUUV+zp1RqSNfM/cGuli/ZBwMlW5pXqu
1VpIKF+i1v9u6TH7zp05wrWWTDrDWf79rfl6FoaFoC/tKNOaBwd6+wA/8LubXvF6
Xyh0+bAEC1ZA/gmd+mn9WhX1c/TaT07b0jfa1H2FHip1/0Pv7A1h/mRz0FyEgJPn
hUghI9Aa188PvHUsqUbIlsp2+uGVXDd/VYyWVO9DqItt6wt66RSVo4RlXWlIBtiM
pNi5600FxSUf/UrkWydMforF8yzn5GIGps7tR8AQM/4FHfLZ/bj/Zaj64g7Y6n0x
9TvII/AQ/WE89X064KSdSYUXFCyuhr5uNAB0HpbJ76552Ha5ImBkQ9IH5CtiIVuy
rt/uTcyvyLVz0nJPL4XKvF0RkuN1oExaIWgG1IkT79X9VpkvUXppmkbCfvrtwJON
cmBIppIwCdABbFbBNMjHqxzk7rgEPPP2S3fBNVZF7rqreLjXIlp3BLrHTifzUBnd
5RGl7vppNUSa3r8zBgCrOrP5YiMuou20RPsYxuf9maTCZrZsfWKlbSOg224Xcdse
lUYOZMn3epfDyi9XTu7ggNJA/l7POsIQG1B9Ek6S/XYel1J645ta80JGORnKx+u6
0gCOALvrStkt1gdD3plnsHnfTW7H/m7jphih0ETXsPHmISiZOGSecU8R580YIVWQ
inE221mh+1rT4h3u0KMhD1ww87ekUOXXOhO2sVdu0IS9JrKpN74/8wzCTFr1rknr
fQWlfJuSr90DiADqLLBTsDixEfFcA+elxef+iK3ePV5FG7w7TKo6kIrOahkco0U7
0EhkqdotsD/Chnop37nJNgEuRv/ItOzhHt6Ui6aoDhRJwGQy6Kz+j2QUg6ZUqxv3
NyTXp63JYqal+FBzS3K0yHJxdbE+Xjvuzr+1ASKVH98EYdiDVARqHZSWjXBnx8jf
5nIag5wghxFaOzIlXxmyTtS04v+wFp1xoK+qbNVj7jk4DKBUYeoHG4xEvnEtvvBw
apcy9jjBb8fu9gK2mPLsnxr/zdMJr6DmmfCopszvKYYNMJKfRe8D/0orLFljLd0h
OEPCbAT77YC6803aq9tu2pZEMOpXvl8bS+eDG9sGwCygOYQ4Q7xaDJfsJso5CU9G
gE0KqEUkgnFonjGS6Dg5oUNm2IdW+ICjQxXTaniAsEUqow2piExpvM4mXpSXcOvY
Hr2q7cu9KoTWdX3MxLNsB+9blD2bbZpdgXwRm9aA4dQFjZeKlX0UDOyMQ4kS756t
ZVxHDA9eq4a3cxiKT7uXBrhtY8DzO5pxr2pdtWs08nuRSrD/F+T8OI080TsdqZrS
RhRZjZHzdj5UVA8IBNXGQbG7eXkx1K4gNl8hXbrrqSKIBqYSpUgHOuOsY180Re2U
zDfb3xpzq+vVNw0A/O2nOsHAnYkL8VYnNiiVtL+xn2prOOQEeRFePvhYZi6bdnEN
zS9ZgoHlpNKz72jSQKz0MukavfwbJoDUPAAZQT+SyqDEBB1mARzECmM3Ag+38R5J
S9mwkX232wceD0/9N+Oo/AfZOROK+12PG++ImybxQguqKFdwstY5glLUllScgnbt
7/HDgM6Vaooile0umDdmA7rNsEVFc5Ptf1PhBTY7htjA3YoH8PKr28N0cAoSC8FJ
BvakhbQmff9OD7gcvcKaSw56hrCLqKYAdCho6FbTjAaLFRR42vKtCskLb1r1InHy
AXXys6Y23vP3x0qy+Cu8HUopPGBZ4VH+Z7lsTsrYlCqVwj/EUfYtWkWLFtCpV79Y
VU+DgkVPjvQaK5dxtRDDCVVvlBXbBTF/yIWO8pKUtE8sUdNT1xuJC182u6mSeB9/
+QtqN9NozRDL/+1RCEYKR0rpkCkT7J4LwnspSt3rvfAW8FP0zRQj5iwNowcgp7uQ
TI8u0qMaW4o9PmKbodziD1dsMbNHJkUUUlscuaFpKVNSWqBFrCPpQmBJOvWM7V11
Reps1E717IWB4CBzYQXe1PBre7j/DrCv0pljKwd4i/DpL/L+SqjlChY71eMs4dsS
4ktjcRdNqxmeethgGXejCEmpyduWnBOmedbUAd88RaPNsSWmLua4rv1eSBuBuLy0
hSi5Sqm2Vx7rxgO1JPoOg5Xq+Df+Jrh6ATVeetsfJMEhLVE07eN6lEWI12NLcVjQ
gQuvWmeHKj8VcUJYYuhHX1JUKMnyu5nNwDiNt/gNl1xGe21rYnhcN7kzOkmWWDWn
AEOwf6CgJrmN3m9xH4JuCFSzTWz/RdOG5EgxF3W4UWfLqZ5Wi3+n4JvOl7/jx1HP
MYYU2nQyVt+pligFbcg3nFnqlvm1zoT0S3HW7eazgCVsRcwktUEERotSh6mTq0t7
LjtkPc6c/QH8QGsC4LKCPzOyNgAub2ayFOg3cfW8TTwcFQJpo9yRDpWTNDagC4In
tng1jBCLwAzflIuSKaBobeq0c43+rjW32Sedok9ixmzaLxkz5Co6YhOeysr0nuEt
xz1PpkwS4WI8Ve7ZuLXAr30acTnMLLJKYGua7euFWpb5nWFUrqO/vjtpGg8j4Fmk
XkOa70NdlGaxmOLGKqKKvaE6J5CFqnLKLyk9xccciyaA2uWp9unv5350qXW/gQNf
0y3D2/kGjLhvClvuBBkdOYI/oHTYsoN7pTVRCUa2XEaNcF8HNCR8Qk4f84OhIXSd
PffnSrJR6cOA3MXytDcwGDE5AxSpK540YU/o94Fg6QDpR1gYn0yzYp6jbOeD71ue
kqtLWVed8Mc5Ylt05Pm+VOvtf8Svdbpr8eYwBCLw17uvHTt7kGTl+jPYPOUsqlYs
oQAkMrecm+a8XBrVA3y/wGkx4QJzrSuz4PUZImDT0Ab35Ocv5Q0nwRYSjt0Znlpk
cP/qJNFbPLlAchREAb4/0VkSbM4YTaQ0FAMNohlyLcxP9HY8RUXVXmXuDQMNMYdV
dGnQ55MKfo5iPwU+PrVK7qgjIXwtcAvG4nXNLxpMqqIiEN6tKSI6P8KhRU9q5UgI
TrEANCFPUznrk9tKLcE2/ixIJQtcAqj75xv4kVTOrJ6it3GB2Q9xXps94rC4YzRI
lUILTQavLcHlOpQP5uN1AXTTvJVYgbi3cVJaVaiko/HMvl164DVbE/fxGxKWy5sT
2oZ1KRHuw/WHQUAlsyWYHimvbXxqDEtA/Me2e6YGXiHC8c4TjpXvyI4jt6lAT2H9
R3G1m8NX/7y5P3oLr1ih/btpj3I/EvGttbC1/BC+xpscOCYGFS/Fazdwiqme5gc9
UA2L2UPoaWN2/znUlWH8LkYguen44DzGRByHHbrcunl+O1A+GWnQdApxhhCV60jK
MRNkcr5DqqjCd+0PwnwvVQ1QLp0+yg7wFyEaggpU30dFPba89q8X5DfIhLmq1pLz
XIc8//0diLOwkoRu/dS9z9aH36KZS7U9zCejVESkEoJ9DAoXbKIxrKBiup/x1KNz
1KpFRa2yI13CtKL0jyjHtgb3O8v7XKFxMKP0BAunTD1rDpPili+MlclprS/yeizq
f1884eBGwLNLTcmNwbQ2BKvK9i2lu2oKIEqaBftT9lwDDcp5//oCw6gZXKrkc7a9
wWDNwFEplIqV/OFIw6J6LYTGKL0B1HpLmTwfW2INjFAkgJk1cWeD/Nt83nyuK7ZD
sEwpdVr30nwnfqSA+geVQYWOt3qQn0luUsYZSATcuD3uTNtDoLF48rnsP8tJ4srI
McgkBMoX8nAJyibQMZhrJPGbTF2v2xYOPuGotmloYnoTCdShUMrgodGBVeXeakJT
Pd6a6Uryfh4ecj1jmXBd6dLfmJjM3aBHQBE8wf/yU0ycMFLPCo+X0qxiapliGFvZ
rHjYohX61iW9Mlo8fcnXFKDXu+ALja9n/c9j4n5HwJV7iv+tbdfMSGX9Fm6pjfTv
vf2t3uBWqazFfupjVx5Hck6Suu0DomhVT/ILlZu7EKf6RIHJxOmo1mIg1xUspwDX
rwf6y5iIgyH0H5uxhVllOZ8LMrNMWwbvEGnOuYBj5v1lUct6I8ksRUieqwGHS+3j
En2rBqefZbsh0nNmSk/3Ec2csUwIEX68bCxM1a72gBBalmL9EqAM237V8a1gwtYR
yEqCfRGhq6ZTpOxG99M4qCfWcbbbFdigATHOD//E8jDFrrk/wUuq6L5cH/6heUKC
x4rCYTEWNPOBY4z7lNIBar8Kl5k9kSAUJNL9jmGWN+/RVxaNqxPmkvTHL73LwOnO
RsX/RykZzVSCTIchWB+68K0y5p8yb99zSnA7iSeUa3c+V6mA02IAIxP6yRxToD4E
t5bRnCV7Ixi/cgzoYVA5Pxpy5fmBqHfEo02vdJyzz7+ZFDADIvP3ESCXpMCIe2w5
HQMu6/mZvalZl70B6287NxZYbINff/BbtJmZoyfuTWDdxOvpcMqmGS3E00LEpULR
BuyTL1V0FpbwI+Xs1jRg8S6UEuIC1EV7r8Xc+3t3zwS4HZ3MdhnLaSJX9VsS3Xnr
0o7bjw0T5OjH5GgJX4L7afJPEv+34FmerFKEqEgH2XmDfq+Ub+ItWbOhzgAU8nqo
CPQrLgN9KIO2anWpKwGnUodncojt8YyTd8EjB2SZ8Bbp9MqfqPIE8+LrkdKzFUJH
0bz5sQP56EmPFNe2AI1YtnxzhRssDb7LCul4FTmoteG6llkxlaLVISESLCmfy+6A
49I149DloebU6FeDEt0eZ7GUBmvSb+qtWe+FZu0aacPNrZGaLRjME1y2Bc2+a+BX
upqOZEHC+9llgd3CMwJEChXWjmBUI+wNMaavmTKTXP1HyoeNm6dBtPIuKjW90kA8
ME8TYLlVu3mQ1LAmSrx/V7Dz6l3pGH3zQRnfYmiFZkgJ97ODoVUhCNuQBisWG9Uf
UgepAV2vkfiB/lxd2IDds6wrhgMC/msvwjhS9A+vmkFnyXY4YF0fXG4G2szffZ5s
83L72ynrbZbCslvCYBJh9EV+VWRKqxrsP5GtP2X4mbym/OdZXuC1dWHQlyvZej2M
ipOucRv5uHM74Cmip7+OOc2LSOJflUKhFeRD2jEOvOhDGS7AmvUZLncyMZKIsGDP
/awu1Gxp03EzM5HoekIEP9pf6usUvK1Cq0YJQbi3Nt+5Jr5u39YWqhjcqULKkekV
eX+yHVcB4RDaPMd9wHch5fQuvec8Uqk9br7TVjEZpeDn+Uo4+GYv6Bp0N+F8Cgxx
HXpKhpqYnMTxrvqOeaIVnLlLXm1JWq16++ZvXpzCyd+XBdUBAiB/y8jkbJIdhMj6
ktzVaO1YgtIx/Kuu9xWLi70ngBoGYQmouQAUZp+IFAlqGk4imaKBqy+4asJOdMNK
S7lvZZjUsxMS0DNa702d8yp9ppdW5N+3MRmsR30Twc74IjpaUt6WwUSFr/6yhIUB
dxqBxr1G0sfYHBh4u5ANqzPe+qgX8rMXFQiHEKBNtb6595mNCtzoJBk01W8NL1AU
Lm/H3ETKMxOnGVzN4gMChR4Q3jbhyrfpTVZCZETEbptrK+QEC/9+vqBaskvCctHR
6ZgDR6s5lap7hvJtQQk9YDH7pKzD86Ud3KbAiEBn8dpepzDwzMPhdE8T7jUH/y68
VlaYoSItD9C/0fOzxG3goOSsQ2p/0Q1rCPOCz23mv6mboBhU4Gjr8br4HDut9O8t
AkGayaYwTSVEWucME3qEm4ReM6KC/hJNGGzx1GP/eRd19a6kiyBnSGn0XLwo1tL8
U51k9hkcCFu3jmQlG4tlGxRRxMlhdPHyel1eHm2zvvdi9OMZZUB7n2Q8Ftl20FUj
668hMe+ZuiAiJAy7XIzqQqEMwqNbKUd4zOqu5wgvc9OJ3qcTDuCxMf5JNRFK8CBn
n+B7V3UDojV3eSHwPvRrbQN+bGQRMU7W1qzJDTNhb+CVgR9/v+bNtWGKn6v5rKPP
Q3WIbJwjdf8Jn8GK8J54o2pySw8T+hcp3vXReXPe/z5NLY2N7ZwRCMMtHxJeK/1V
qn/LufDeNk1GvyR5wL1w25LpFO09jLzjaQ/dNUDx3Je5HDa9MHEYWs9jESwdd4sJ
GpHkzEob+6w+vVitFDoxmZPkNR+Tcf2fsfvJudxkPghSFqvJPGlRfh3ZTZ5C3etB
4EbbwECzXETa96dXnJL4Ll+ia+HoOKvG6PR1XSOuKHsC3eI89VYmT5K0WAshlE+V
qrUkRvIRqCnGhm2PJjipVWHCe7a+ZaHa8T+Uq8+FNzc3OyHX7dxPzjyGBya2erJR
qwEzvTp034QmPAQOEcZVHLcKzRt43VaVDBUzx40pvcKEAOd0FkeF9kvmC1S8UbgH
m1bTov5JyEozu8ztmkMe+A9G0IRtAQ7G9Y4Nnf67hhBPpeqa9KitSerJpxuy9otV
g5y6rzW8dvhZ2eZPvU0nn8mEmizEIJEsPjmW6p/9wclVNpC+hX0n7J4NQB5oWqeY
hJBNVMsZ4JiwcIteYSMLtGeEPqoS87otpndcRXNsFqCUK6a2QdZpBTVDywS4VyFp
iOWNk9c9V72ohKbDoqbF3Fv99A2RTvPwnIA26cyJ3pyJe2jxk93Ak5s0HJsv8Yxr
Wd7n/J/BKgQZmprcdR5IjGyLel6TmvzUJ4UDOAebcfBJoj3RzbQkD/nUy4VFR17h
q/YTTDlr/svlFonrgqQvvrDplBJbZcaiyMcgKuj3fA/InbQVgOFn1x7digPpr1C9
Dzk6X/QJZo+wEEXsfAdleiLV/V/hv6BDYt9klya6xAfKSi084PFFZggfD6v7twMc
hopVDeSqdvBiLv5LS9B2vGNBgZ/0CkN0iJxMeMPF7lcD1HyXexpHZXsRPNyBp2jW
ybIKAOxOY/lzEVtgWev8vLdI0e2568b3RXFYL9TvyCguOBMRZWy/Qt75zvkxMYKa
2oMfuynYHyVUrZnR+JeQkDP+D+rT2KIW2ru6LnU2bOveplf3RpXdEPpRsU5CxAXn
5VE20zqiGSKvjoJCrrZtbH+pJEps+x39KPLO0s3ws0daqYyVqB7EAfIvTW+adWZ+
o0rCO1xLFSdQ2ZGjDjGOGfcuNLM1E2djb9MVrawXTqxiU/RF0Nho4Vh4vYwJHEce
8/hEh9cHdPOrO2lhvYdoxSsHd0hP+2gu4Zwp26V4YdIT80SvbO3L7RPZOOYxWRUn
/iAh/DI8LVqZEpRwzWAbJ69LY3vAhD+QHyggyscS2b/YVCqH+2a57dvRqg/dUTdv
dY+426xtj/KpzfWXRbdg80D2Dl3mHqdmKfpdPSk7NRapPEq2T5BA7xSY6XNLQv/9
bO5Z34NIJ1WT1iRKBZOAk8Iv88Wch5+Izv4cIdMRQh1ZvfwT7eodC2mgQJsKEYRy
E8VvrDgJEkGfahanbWum9t3SgPcud4QB8qjn7D3+0DmxWlSmMbkDEDfcQSOc6WPH
wyxof9Q0NQbBsHfg9gICyPagn9rgXnbT+G9Wj4JNQAtpWWxUH1U22KFhPXxSg4eZ
v/sYBPFF1H255+Fz05VtJVMlFQb+iVH+/gtw7RRRUfVx+Xts3PDQ7Bi3yvIlD3Ao
OvyxpBM/p0BzDkKXy+UarcAM5/TPmyGPSjyChfMXjfIT1IQgV6Ypden4RBXdAKmW
Ay4He7Xy1F896wqRt1z7yhyF/IG3yWVJsAPCkJNIWeN1dJUZUNM68fsdwoO4mnfT
dKISnQ+0kcIwEVT2jNEGQtuNnn2Rerl9PNR3+Ot9CTBHPhQHR/RPxrckqD2atubW
NlCdcaNHDc6W4tnb90SwCEozi5/DRFE94O3J/Z7UmAUPpFQUe5UJkydL+18rzWX4
c2+D746HdqXUnJ/RaPFsS1CyHC/XDx8l8n4tiZ+K41bYWPzOMrldxsYNx9W4JNGh
8+muuPhRSbWElM3XzN3VRfnIK7Y0mag+gi3hwGH4ZaNRXqbV6lS5ydyKw7j16aTy
DsKMaQG9R80fztt0a1iemrb7vSIvMp90X0p8Ck0hZtv0W1cdBuCNZtnxJHdhZcn2
va8NA7ejCWdYIkZxSxisXRne6ExiUOW9FEnBJVe0Kp82qtZtsRa554GCUT1TasCL
OtO+SiZKt3Accq4zOJzkmxKs/aIYa4RsFOQOZd7W0B/SnDqbgvw/0sRCy4QaGbn4
DKrNLA9g8R4oBs1PM6Yp40E7t1nCfxIRcivWXQKWIiI2zti8Xlw5iXUu5fl6YdQq
obU8Byp2JnrA+khYtzq9C/ZIL1JLp/t6u2H8MP07xPir9mOXmMCVscd3+uk+K46M
GYdnw8crezx/SrFigf1HcVpUrKm2sIm/4vicPKekvO0Gd52/tpm3yGthIHd2hUR3
EpT9gUg7NjEHXzwh6jT8oNBRFsF7MbthXjJbOG9S1B4KX1epml9c0PHIHhAGnCQY
+kyeAFPThF8bsIedouWLM3YBRyuAC8Tff0a2elxIBTIHFnqmv+WYCNTnBfyeNHYP
bjl+Uvd/NmGKB+oMHy0f0CL8UjVBTwtg+WkvAZtxypnJqJjsON3xIlBj+vzENmIw
WAqDwuknmgkEwYVtqO1K8pZ71mO8pkJPXFkAubLEG3mIyb7OMMV2nZxFJpwxTN67
dNGvdQkEa5qIUtKsvwANonr9V032szb/QlK/eP4+BUfd4Ty0j5t/K+LR3etHtr7c
XZaE2Qla40TJMywvZDR4OzUKK/NhDUweWkAIewaLTKdWtYG3P9+g2AFa54ORAQ0k
Yxmt9m+rpucmV1WBTr6R16U+aY47yFjjzyIelGz/Z8I5rG8LnWFcunWBEaoynQCf
GgDZocdfzzY1x/bi0pisWNdQjOwSzn8+1mobouVuBGtSL4jMc1uzKmAz/Ik63DD1
lyJ6n7iz8nUOIPu2PwHWKVg3rNSry/ztmhHmomyMbPW5YIayLiXB+S1wZyJSEkXJ
NllHV7xUlj5fl7ml7l2uhMQFDN31GI1n/+ddIFRVmJj5cl/rmrCDv8SD4puT1WxY
rSWISYYpMClMh95f/g4ScYw+gIlaBtEe2e5g2rb4mYqD0iVX3yhZi+r0rNF30W6e
rgT1It0FcdOzOJcRExQKxxNbwWD+v6I19l0xYDjcP2mnJ7//AykERzcL6uKBmjXo
E7RPkrbgBOqQpHypH1InsLUykRRySX8Qc+UFLhVrDHGdCvjoA7wmzdtUAtDnBu5p
bxBMsENpc0W8N0pvtTM8ycXxGHT5Adu4uLFJ3lYpHfofHEtJWDvkpqSlj6zJPLU1
4f3y4ebxCrJxoKPCZgklARfzrPxqwCPMqLqvrtTGGiYZ5h319HQkv2DkVoz5vUvH
EwPJZvGLhYh3GT+si5+jylkvkZMv4MfwnMHO37UQJHXxqqvxLFuEMYtXiUETXO/x
TfrnGEsBrPxfcc98wQo/kA/NdFnKog2O/+jnIizJ4jCaAMlkTsJFP4Ck6fwMm5SC
binzmQ+itdwzACOfy9AOEgT/v1TaIarWrHsXlZqNhT8zaJ5F4Ekm9SxPKIR45qOV
cTupqxJ0K5UtC4y1A5/wrZJalr1b3S0xPM5irITllMSWLKgYbPMhNe+TqEiuQNbo
YEtPRO1gHmYOH547wMNd87vGhtvIp6qML+uUP/GBjMLXWRwVkIFBZ769xcF+QC7+
h4bzTGD4B1BHHs+N97dwvNQ+1hauquPhO3noQJMc29pOSwBef8EwsjBu5Zac0v2l
AT21hsP8uPFeXphKNEtQFWeVEjvDe8TOEnkBLnXskGwY1TBb4gh6AplbF/nBDIxo
QWp3HfCsYZsUjk7PKszm26v7hH8GBO66mHzAv43dFIW7z6Z61vqbYAztTplJPhzK
I7GyQfBDKAT6bYMe82GKWRCimSrlrgwUBH6S9hsqYarLbzAhG4ToaY0kVIsjA+B+
kg8YwxIHkigPWb8ObXH0tW4AgYH/rXjKvjOQkhSIcP4rgMBlS+JH7SjRKPn/h3yL
s2qx6HDEqXZRKGBd/0xznrjDZRRnDuArTKgfnWZWjtWTjxfFmJLRoPTGq3JTX8e1
FNm/9cx3cHEAlLfTP9eEEj98XHSYPI6td1Z7IKaFxJcRwg0VdM5VLHjAwv5/82nC
gP/Andr7jTi7gxXblh/kHt/WSCBgUQmzBs/fAFy7+Uy/HpCdbpwnYP5XvAVrcVye
mfZMkeLn6b/zMmj5LwNTjUe9p6i5to68ftTluDX84HGwUDbqO+PCz9Ef6v2Cg1aS
Y2otNaP6d3Y3MG1VKjBif0gf0VoslK95jz0zl7t+L+dyJRXtAMdJVKZ5ImY6m0oy
iMyA/pkfiQt6OkM66aYm5Ty9XLzt1oDGiRA7gOLle93I91ujXkl0dfgl7VNbdgYf
zjGaU7Mwjbn2kX0ubmLVENKwpPBO1A5bb4vxwA76ZrrGyecmqRiM/rzEd0vtsKXZ
o0T7r3vm0C9BJM7Q/NTuRXJ9e6137Z9/HhnfaWeCsMHz/5dvbLzU+F0bCJeKuJ1F
cjoobiPty+mfn3bgISgpKixbciXC4oZGxEOpL4YElF7iuDCPoGplbFMYOxug5EL4
XdqCt/VfFFzHeMtdeegm4X5za+855OvNz3ftqDaYY8/2mUAThxv7lRweMx2p/S9S
BDkiPH2dwhmJTc+lMDjW7ZHikuX84j+8FfvfUTnqFGCld1MFNAn/6KjJWnWvB9S3
7x1j2cfcXSTXJbb5S3LhuTEmRwZ9brIZFFJtpkBMNx7BU6asC688YlLcgB+EcOQ/
qfz9R9gz6whZfVno2FaDZCQybe0EDusz76VfJjgeE9i5OxSsOa891D+ORRXjfjS2
D2HFGoukzNuEwb6DV+GYwnV01REl8ONLS8ccdgMBKEHEMu9EDaetODVS172F6kEe
elSBCXjIOccumSp6Q77gd6U07B6jvXe0y4shNyyUcIYbOil3ssK4vIZmNP9Btd1P
yFNYM2OC/cMoGtnDk6uNF8cK16oMaaWCJaHbZwF/+d+/Kh2Awq3ichYPu4kBjlbq
t339JYKyweoLXy052ijqfs97fcqna9F7XeO6gSsUgVgShcT7uBYeIeA9VtaKXcmZ
f6zry7BkDuIDayAhAIRwD+5JBAk/4R4kjA5oCP8kwno62RH67xDJB33k9QE4e+4+
r4D6j6dmk00Lxg/GkgpUS0cYso2wNqN39MQ/UQwSHtdU83bJHKqS5Ju5nuUpJ0BT
R9lmkWoyekA2oJtsWTJInn2Ls379+uz22pLQmqXjYC7yLludLXM4DDUMz0So9sFw
Igm0cYTvYDnjCQpwgF/vbe1WS7PTkjCK7MUywEEqC/u4hCEwcolaE18ozw1s7Sok
crEd8sCI28o6+oHoegZOlEtVqNa15H3T9+myd/uKh8VG5dLxLtR/bXH3XUPImLkw
8EMOlzlpz7rAbTE6T89NKJl/JXG5Qb1GBfimtDwLLfq2VS/gl7D6M7NvOMjyR0EJ
YDZQ00OadoAJFE2O0FzsjTIpwLfdUFQQq7WrgPunAVR0mH0oml7s6wwUGodz798T
y64/9UlA8EZq7ZHcI0pQ1mj/qNroaIoJBdG+211Qi3u/eoTcHz3gBZdSHs8xlElg
FGrGpU8Dpk4AB7WKV23UQWV2x4YYBPryUXl++ZFVlMUAG8ZDHdV+zkIvNt/G3cQZ
jYSKv9SCVDMwk8NfqulXZYr1HnHeSZ6iyE/v2dlKfNnWqw6RZROx7afCEuP9dket
k/bDGSRMA3wwMPtptouX7+yAxviPjOFePphxN/ez3LdB0ULyS8ls9OBskTuJrtbE
1XVxdCztqbYIVFCY71Jce+JbYhYJp0gE3T3T+BkLn1YKBG1wjUJVKCqNbm+V8awW
QLOoxyPOn+21HNRnwvZGOrNVh7MAfVoVSC0u49IKBJRDmvDRjErC+vhVfFXC5TkT
D1AuvkBPxnfZrUzB7et5VPJFsOua9DYvVldoXtAD4CI94IdZvcudBpf/04wq9oD+
j1Iq0ZK2o43s31wnmcZXtZn03FpYdNqkoko571SKcdr2MlAUBCPhGoGGdG+HDoHR
kJV0CUN9thiyeVEwQH5B+fQaQ+iHzGfmgWiF0Ma8t5Ccgud++OWmhDOgvPx7zA/U
gO2wsCl5t/c/Mb7R0hd3D46r7oLmoxQh4nqHAsIz5CPWlp5sUFQPXwRHnVXExCSo
91WJ0VN+q39JydZAwrFkxIKDzEUtvjHv7ilGr3/rfZJUIx/kmQtwzF2DZ8smcSxR
yvPTSG6XZo5L+jjEa4bFClmZBzX+XOyyOgK7uzbvM1O8/CgDruPbucBOXGAicrLI
Tjsnbh/o9o/K68wUPCsqb9p3u3s+Gx8lK+F1tYR0us4GrNuJV77hzoLYpgP4ItGD
sU3fBMFunyxru5ijtenbT7wgbzQdkCzpxqUNq5Y1JYWH5RnTKrbtA7nW0i5bTZUO
PHR+ba1M+fIXnrx/JVSP2+jhC7khtby0tm9NDTH6F37B8+S3PZMfjrZJI5p6NiOf
hH2c1Qxr4XjT6bFHoaJHuaL8DICv5h3PBBFubVBedihan1MAWfBuBur0aNP9ybgw
b5s4fOTcfGXmiHbX1JW7Kj82wKdToKorullZlv2Wsviwl7f8dr7xfXAcE0ALGIDb
M12nuBVwf9ztLaE8rl8S8YdxhrLsDwfNSJozPQoFwv18o99sJAkZXiQNJBXe4bz4
OalOvtIjVVL/5i85kVe2Tt5ssjL4sAI2uZ/e3hAuQT9zpdgM7CEsbsbBYPMSr5yY
CvLVrNKstn/ZyEtiMf3HPLpn8uDmbMIyp0UCvkufU9efMV4OwpGdaV6YCoI7fzBU
xVGRLWAh89footzTuUBkWe41QEoHmBghXiJc1q8CTYryEhWH0p98SL/DaxHZfRbj
pqlxG+t8E1kirOQz2Y06+A1H6CShKyFB1fh5XgV/ebQpZyF2eJVW92U52MENRIoc
oBIm4yJw9ADOx9qJXeEz6NBNbtN9AYNmHcixqDT+2GrNIpRSf4C5mDLr016TWPgb
yxiB40fpGU8CXMPEPGFW91/AnnB1d6/85sM2xtqcTj5RhRtDMI1RXeflDwTMEFQW
B1QQ9HnssCArVzk+qf9ZliZji0/a62pxTBqmnbPOdTD84oyNVA7qqMbetUUAHjBt
Zh87L3uxGcQ1LkiK6WvkSMjiFsjmk0Mv4lhMvgHMwyIJxrs3pT+QJLyXHL/rcr04
ycticpdK2O43M5PTHUoz1qRlIymPt8XQM3P8FSp84IRRULJyRsv3XBrdLEKjC+kl
MG9SCHGVozGs7pv8vSKWR1Z0gxkK6izPlLQ4Tr8abpGrb8lbCPKkn14oOa8qEkaO
jpG8nI6rNxipMbXwXuQtpH3M/ELL/U+tz1s5+1Nnpk5n4pLskRdcZjawZkmogZaf
kbDScbH7e7TbkmYoO8+2OvfONZ5lXrix9bxgE/VqWk6tsznBlR08AmzSdciBUC1c
ttMS21ZF3vJ61qOvgrF1Hh8uWZShO8/+Hi3/zvWRYnC79B/VFxNexDTB7cOV001H
M8Ab1BOPdpz9t40Zp+nh/os//wfAnHG/OSkbpigT+YmwlMCFy3M66DjanF5VTD89
QWQmgRvxIIJOuj6dHRwdjHJrW50ZU8WS9fBNLX9CAfCSrzyVg0GMvESy9LZ15LcD
xhevqPRFHFiL2uzW8EJCiNhJiuf4jLMt6OO0eNkreCdrkxsSlgfWHyNGxwGLZNb5
7+M+RWfLFR7QGxeTM1dDIKXTQbgfYHIHVGKMrtDWA6llH67XqeCcy85q9BmQHdAJ
hgKq6Fr4K6TnmQMiLSqLf5IYSqnsCr4TVYO3he5NNTBYuK/8DuZCfmlyHHwvkD4Z
WF4t134XH+bUw3lphbJhV3nVtAw7C+nP3RarA3hzZh+lc0i8ApwLW1rbAVgV8MkZ
GlUVgmBjqAPAxlL2QNaSiCm5FSCtmKCEPsZmEfx3czea1P8vcWfqfbGVnsTtePVD
vwIuxEKQ/smyuBjAnqhG3g0I1Sur+qqoLo4cOQZljVwITMdzk6pX2Z0Ybgvxxe7y
+BiDb1qbPR9UPRTTs307+rRoi8rcTCs3fsNpVGDTm9u/F2GlUvvznO06fyVhpdZA
2C3oTHA+miSSkOzS8a9bLYUBBtOEm6nwR1eqRgEfnQ18V8mBmv7kPG8LBIX06wcf
mvIDj8B7Ya+KyNbzJ3Vt4bHsceZMDelr5h69tmKibpnQbclTCqILpXFopQOkf0BF
yFjx0Rqqf8WhQMNiOaDRTeSX+hi/0FYSlgwcSf/ldqVENZ231ZQgAhrs2r4zAXie
jnxxRuEF70hZoNOr+eRH3MUCaZIEbG6BuCYY0L67VIWyApS2CjWjO2gnkplOG/qm
hkIZ9Uyl5esa/whiuJgCDEALAPy+cPeLB7YIRwFb4lAAU4+TtB4L4vgHxJKck63U
nWGYvp7kCOpx+YXDARaIXRSILaKG0CzVS0tm8rMRFTulIatUJQt0OF520Yd44iUm
V+ri3V/YrY9aCHQbUiugNnzg7xqmTTLbBAa2dbKVtHxIMcVoWjY+FIwLfP6l1Bw4
aAtJl0+y7DSnZH94nrig6CwR8hGRw+CU4rfw57mYExs8RNvgZRI8QJw7JQQStjuL
rtmPtQoCxGhHkoJ3gGXKE9eQUxcdxdlQKVECPm98o+zUIS3FU4YhjGE5mot95xw3
MC5SA/slivvvAcDv7cxNoS2UTaSmkJbUPULVNkwzPgBfUEI6gcOU59foeYIwbEd8
RUiY1F0PWY2xOpuHGn86FUuATelrYzZ5Co2yBmqi6fMTUCCn3+pub00+tGT7mfsK
aWPOuoyg+XbuJMCEkhabJugNJOekqt7g+bWJ+qWjTM2QEWDI6Q2GeVXBNwnDKbMz
ctqivY+BXaTODQce8wmXuhvCr8yrqbuqX0zcM4Pr2SjjtsHqljBuiW39Xa8N1pw0
KD4+tX8vJrfn54D8tjlnc7QIF5jB2U2P3L+Lzc0xjRWUdn63DL2R+DzCNZNhb19x
h9K0wRY5TueoCNAedEGq/A6CGsi/lpS7Ljmp1QWbGUkIU1TWGLqzakggPJUhWYwk
9K1JX2BRcc1S5RAzJ/v8FbG1DXLPPfsD6yLyOdiJU3ygXzPLYv0fqEdqXFmyaiDF
WSgYOZEILzTA3Trdfe9+THxLyRyCa3lsnoodHACbN6EApahStaxXMU91KSRLXrE2
jgTMbDdJRQE34YuMGtI68xvwtIHeO5Sw2fT9Aqqg2qYThE0X+J6ENn8Rx0sFXrzT
sgjvpC+VLp/hGcQgvv8Zw27rYBDCLj8RUcQpYEuYwrAyqxzKpKAfOirgzo89VOMg
o6cKZpuHZ0+2mUjpl/Cz/hBcSpaGCaAxetKRk5u6vS/XUt6ydk6C4FOAI5wGzZAi
FRNW792S/9pF7uDhDRExq/t7BowGpB8G8ac5bezBQpUmbEUCLjpnKvtLr4Cn8/6Z
NAhyfaiTbu8yuu1svdkVJz1mEnRRMiv4it5rH4Kw8Zk4lXOrWKJsTSvxmRxCNLQO
iqQzLAvCFg1Z6E4slLa7+O7tEzwCAljWSRxBYFGDqyKNKnEIS1ljx9xKy11sImHO
5fuI1tY/2Kbwmo6y2N/YTj8G243QY+JJRvVOH65y0F7DvVx8Pc4Qo698AOItpVkN
ZBAj9SjKj01O47sev7NqRuRaRUJMRH0hkWVU23WPG4bys9Ok5FWOKFINg6Z/YiSr
+uwFOqXOZhXqcHKU5ptM5MhSvnineRTM+mA5CKC3Lq5ckD2brnCkDCyDaEk6g5GM
VUMpBYxvSDE4qklsfZAjo7frBRcVKLIPETyIYY22PvkCsBmV+gIIp6SAr9/yQG1C
u9dujyk2cOohieFXtAYX4//NaXcnBGihYV/bSvHwDTGdvRbeekFCDnPfIiCuejrH
3BGRlnjVv56fO7o0aTgIgYahzaW+TjXQ+xi6Ng7TIZHu/S/jVMIbkmB8kJyayhra
s6GZuRFWauMuI+bWJVHgbc7irNwq35SO1FGHHIc4Pr/atKtEVrHgwymk1Q87GarK
Xzqs2tuQeXHtFt33uC5MCtXHZayTPvdqPIuYhy70Q4fuMUJHibRZTIrGRpjNo8X4
KNfKlE3Gp36/3KWkHMBwZj594Lbr+66y4ROHFU7Fhqo7p9qp/4Y+DTu8LXOY23We
gfcLPdWXiH0lOQ7/NK+T/JkGVb2Nf3aP9RfRWRNoYnHp9eyZCN6JTAz2CEKH/d2a
dxyHqXfDDnOJWfzNIh+8Jvp8k7ryavIwywsK7xN+f6HsBmGysATqZhYD5FUqL/Xt
yRDKdg+fEoJNKJ0zZkKXf78wZaytTdFofHyGU31pT7EXbOktZ8jInLn1r06xf7Ff
DSMeMrV4D3vHQFH8PwBd5Ff0SJZRtEAPRUWkQLyFt9F9bOe9qhBjn+iomc4y6CHH
yTCl+tFIRNdZ9K2J49goM7yteGSRFS90j9eo2kh3arZGhTPsPLHUE8CSVoSCUB0l
55kh7p4VJMnX1bP8Rn5HA+Q+ZrBS1cKfiIY88TWIT/UnT6HU/ldBOm1tAITF6ouE
5RWlqGYEicQ9PH18P58pAze6PKQkclnYhCrG6Z1ECb9Qk7BNygXXUy7eRIUmoayM
zth+hNnhYwr2nK5l88dH77XbeakQZWetK0teMimFxDIzsf16RYs2RoVcQiP0AwSe
dy2JD6mhKZuRlpqUr5CR/jNF806zAIx1ijcbwcnrmB6/y6NzR+iHAwg4sTsLwDx4
hSwkiAdscNpy5GnKtxegJnHD2+HkBDG6JCo5LT7640KnEI2BRPw7WR69SlOcyowJ
yH2t+fCTUq9nfDsJ4BGw6U5Evr8c30QbBrPbjAvsXpOvV+V8DIUGfrLhCp9J/aMJ
WMQLagMJONsAs2dJxzOB7K2C3v7oLth7J6NQ5JjPi5f4RjFNGlPHTf2mp999nvgE
mzTiUJu0sxq7GtzXsSwgEWS1kSEfY+uKtVJVtYxh+6qTJi+dYIvdsEXwxnjfsIHU
hLguePYFnHuz9+2IbU5dYO9YuzyLW/zWhtV0r8SIIP35X4X0bdyw+yFfIIJv0mBG
xH0OttGErU2qLlgy3yIsrBgITsCXCAHKJcDjOrkWZvQmuDulIavErS+DVpdHuoFF
1+/wIaxOuGwQg6ZTt7nwpL7XI+UzQNdOj1c68wd7VH33gYEpuGn9Pk89+frGMPil
sv+ksGukfN3ntg4RBoJNmqOAE9pQVIuHT+3Ou9M21nh9BINVyUO804MgRYggWSn2
OSVjjLr96DaX7M4gTHMsIjV2DLb+NCAzS4n9i9vdZUcbi0yflkcDQFUwMILrchZt
oZzHWRGmce3MUZSVxvVZQxPM5CYS3rVpMWoI9h2oeF7U8pyK1mRHPJSpoCH2cHf3
LxoO6EEnYKgWAsYX2AkpcvE6njRSMLQaNz8XedCuakfbVRvge5C0A2/HGHwnv1bi
b6RcxKn/qnWHOxsDrVRlOMtWGCvtCzh9faCr6MUdv4hOGmEoJwu2PAoYwK6TCexR
2B1zMjIE4flnI4vhT6FosQjBCWKFkM2CXC9suesE5x5qeFy3Fz8OqZ6BZ3lOZwyM
fHoV6vWDkIFBU9vipRpc2cRprBEYliQV7h171ih3lbnQxYL2sCQdL7hBM4jSUIPD
iXQdz4SaXvdOvT91oQTvDe6Ot9R1Q5GMSja6fttSQ9t34O85uuNLLdj8CWklKWEj
KVWf8BUTFjUn9NkBzUYsSBYcwi/pz4iW+qe2pmOm1lqjwWpLsL6fHi52wDGT1Pit
HtopQNp6b8iHzXw39umGlqj0u4PYEDGaPlZ8USE6n5PGJkTj7fygWDpuNzU2HIlz
9H5X7zsLe6Bbigj/fDgbGZDpcHRr2s2fEPFY7OUxRiy7MxNxiu70JzOYi/GBWSnX
w34UU/KLGke0SahrVGktkFRPVOdvaR/wcpMLj17xsgcjsRtiqOtS4ejZINagkfav
uVYS7H+muXC1u2ynmQnV5040uOfoCMzpF/mNGmzIgUXWQj9z6vH4MIbCFXAYAod8
U7HtT5p/F5LUtDn2mcAEq790Amk+KJqAFiCI3GdrxB99KLsHK4dv9PoWsfwcPbMu
vtEhWqeEt2JAk/gO5uuj6pxzFWSOo4MPkZoPjdu9P7vRjITakeMRRSdeRu2dq4GJ
d2tB+YqQfOF1dE2MyoPWg7idXJwaQoRxyVQJ15STshCIYWciIurW6AxOPt7IH0r7
go7wcnr3Qqllmedw5OZiesb1Q6WyXrcXx2jfSj2iIF71dz4kfwZgxA1E9dquu7ws
0jFqAd28M5VfXUQBunX7w953yZfCpKpA0wnqsB4KH20JOplBSSwnZywBvad1PqfR
ZjDi6TyhC4sU6Qm5fn4rP28EtsHWckGPGO8npNtjwuonMnJ4HqOJHi5Os8i3fUI/
YsljgPb/g+lKmwhG41TeYtgKP9Ygpe4lXBAQa92kcPVuIN3+Ov1FpUYBNMyrFSwL
qA2lPG4YtvDSh8pGV3E5QZZN5NoWW3Y7uVW7jDfP8x1dLkQ/iNXhKbZMvgiFf7Qr
+nNyBj9RsPDViirIOk4o44F+3W1CXjzzeTWPiTrwwWKzuwI+yU/YLswbSShLVZpp
TObQoIl+8AMafUOpgtzoeqI50aHflYyBo/17xD5zYgBmRMTQCmDT1GzMwZNRaRfX
A87UbIc+u6IUU6WoRu/LFdvJkz5jB3NK+k1bBzwV2Jj1vH/cwExEZHZK1gRqY87f
/HScJkeCRRCnLio/mWnbZIjJViMDXoL5Yg7lRq2Tb0DuTHAQK7Mn59W53Mv59Mss
+4NNsVW6xug3un9lyhuUpeOl1uRvoHmfITyFyi//tsHKvREN0p5rl74hfNG9d+7s
atPtyLsI6UzNOfHaIxG3svdPdNT1BGzqNPnkH2dNMGzr0QjD1EvvmPvLi9bP8nT2
wbT4z3rUEHLfWlPDWZWKuNVwo+MqfF5mGBfAcBO2t6r50+kiIUTI6ur9wEXOJGgc
ng85aDoQW+GDSir2qY42MW1sw6HaqGK0waxsNLJGmRMt84u2VvE/6jGoWsHbe/5S
Gx8aFXhA+UGkSGqhtNRgHgkSG0Ztk6fj9UNnKG2QHqpPuozN0FKEksjo7GitaCkq
nZvANYkTOap3X/lLnneyIgn2XSedtglERTc/c62ajMfMbVXOlBkAE2T2wru0Woxp
jaEz0nrYzhg6kuq3F1sxKhijVTvi4q5KODpWuCk7cMpGjqch5UxaB/jfG9k8oGUf
4CxYE1iT6XI7fl6uMCrMvVy1RJw+k9a0tX5j+XJZp+MWzOlogyLUVGWnG2Mjoco8
iJd6WgakVq4QNLSAwRKz/luq3yK9VFaF0DzCOL/gfHWRmyadoCVbldHmlPXnDzW3
XwSTcUH2tHYwgEGyyn3KNGbGPAep7nouLxGGpXQ+RyabzJYpDkkOO2CyFjyWqLzZ
Wj/+0YOnkRlNzFDSddLQUMV82QWceCr/aCsNdr1lZO3+fO3Tk4hz2+9nVys2dNTW
IseeHwxoMcJbtXhq+0gmrOzF2FqYTLES5uOkXIg8M/s185LotMTYjCl407m+fFMC
Rvo999cDgZ4DhzGIX2riL1TH/EYn2zWuQSRCyZTaPoAN1FoOcpmjKCQp3IwRvcCx
H1yXzPKTtEqrKY8WpvHYJIbi0d/QRYyAL62hx8nvhxAZYLu7Y3A6l7CZzXpwN2AS
5X3YN0bbaDgCnTtDvM1eU10lCAH9JZp7QaJw6aowz7QsBXJzLHm83XsELhWhl6wQ
benMWe5w9sRVsegPpcPcERlJmySYsoNYfNY7eVNaOlIk0Du8kxQlXGKz7dNqgGdB
lax2P+A7CTH0LAMThbGpHxScEPw7B6AYuNaEO31tqzdzmJsoJYE6zn+DJpn97kE4
vVBkXJcUxc1EoSgvjADxySTO2OO2IVy7QjusD/la1yWbYWdKTVx6TwvunEfMe0Ze
+wmylET7+6rqZXHAPEnDoyhhG4Kg2LmaBqO8NiUF4HshHNJ81122EWoWEh+PCHox
q9Swba0RlnWaAuV2bOrmI1OW1N1gBfexTP3BJgYAX9LiTc5P6lljAS5ggOJcZZe4
2ynkJdaM5EURXKregZcM+2PO8Q/wW+QCzJZLY/RWAZ3LLM2bJEacsaBuNxctGbbC
PY2DE8dEJXHtSK6491gSO5Ro32OcghFSpMrqp21ydZbRJXzF8qpuKpIOKFlDbTCB
bzNE+Z4dy+fFuL2Fol5WjVgBkC9YOztYnW0+Ca45BCNBoDL6G2cFJnxbgUMQoqoh
gWeExoFLmgi5hdUwjf0A9p1ULerhjFIxxRq4wscZj4QvVz/JH++FQ20koRQbiu6E
F9H3O2ssoqFD5om1raFnxznx1fGh/vurdyjoKoGHnWttZ2ltsMNibZVbXfebuvwn
2ISlC3lZ1r4bJi/foxU5xttBRSY5msY8sdywN0k35iOo6bvEc/58qz4fqvpFQD79
KrauGlPpFk78+stsYAR5Kx6KLwU0KMcv3mzcjXMyXyY2xyzzR8YwVHWGMpSV7jaX
eMG3EHMFgicxZD1TMEPn+TAsvP1+XkGWPePnAInawOG+L4zgLnM94JcVKmuzNKVQ
3tvagwLc6Ugc3CWUeJnas6IGzH92A8h+wzJRDC6zv/uxvFwbtNz1RY8rOJGS2B69
qRJgJTP3jmUvER4tFVvxCvw458A5nRz3qQiWzT0a2Xt8vte4KW2Q9iP9Mpwam/46
WwfuTD88fr9juKN/HdyA1jHnaBxSOeNyzB0zpTcg1d7Es/KQr6xVX5OYYHz3EXz2
YMiv2Fxp08Ohtrgpgi57iglos6QJicpwIsUOlrzYutMotJ3bYohkiqNerTg2oYpM
A4gzf0s4TneTyUhkM75Q1pUS/76L8NYrvT6FnbHyo2l4xSUwjI2Yw2o5aMr2OBfV
nMQLiCHBEV1lnCbTPG8K9PDOGkIGKwsDmINNiUH6l9ky1+nU1OZXzExiGkLR59po
Ho46r6JpBiuuE+FGbFLLy9z/glNJJ56wTaa6NemYdThJTB2FUESRWuGSVuFqJzDN
yChYrLd1lfNxQrHSJmEDRCeoTveoW0hQDyNrt46XudnBzZebtBeixxufVJxKdmGi
J2Ogt4iYFAbJNpuA1C+0oYkUAS5wtPnGu1xQpPloHI39XdnF1JyamsRpaxOAxXvb
p44QSFCSpyq+IW8b2tSYd0o4J2eB/THmgZDlAroGKXLm377Nn/YmiZDspI4bJDLk
Qqxd+0xlKGnm8+vQDHEiRTDOGJQEDrRLH+N+QrvZSRhAgoyKLGG3gFoy+YfCku7j
/zZtPuOAsyLuz0+cGe3DryHdAQpxpGHVsSOkUMyj93IBlQlzRgPVqIpc/Tas0T8X
myEgOYekOUFSgH5SM3krfVNXD5G/OQqMUPESkGbG+qWcJwInkPAkgsu/REiBst49
4kWWGIxyEDcZ81yjP2opthwx5o1rIRrzSymLJkJhZffT8dY4idRrIute6q9vOl8P
IJ8Z1JmtbyfWjzdvh3B64Y85r9sv4DfZL8Gj6QwiwbyOiBGuywx+063iwkVGJt77
3PDNF3pxPoWFUmJvcJ/jbIqyoiStFgvxn+8Z5WXvTYf6JeMfYMCLMUAq3b4fLraU
O07T/MM/Gs8HgtAVUwt7e0ilDTJmGwJm998/ny1iVsWtBHUkfPwl3WAbNZ+YXAYS
D1A4AIvTCbRRvhRPMPCckvgIeINVsWK52frvzVOhjuJNmyZmFvYCNXgwLMrExXJz
D384NcWkKzIK3ojLUjfk48xmpuUk7TH+Q32vTg0CY1286fmYF1/9uCO8pdXyycIY
eOJJd1cOV1rk/nNqaIMa9gk31LXOHlE89L7x3rXeQ6CRry0OztBSoFkKz82UTobV
K0GlfxnjOM5HzDsctZTodRc6lpcIoXvN340JKOOU078/nrIDBWPl/XoWUkoHlRHb
l2hg7K924vLNQ3J3m6LNj72Zttvyc2Vtsrtw2LRIoRkTOFnNOFxXzceyO7FNG0c0
nCsSI+UvGCELkMaDpM3K8QOIa4jeN1cbhloAWNNbRWC3uC8A2rA0FRlzjpzQbb+r
M6j10X7EcmH1VPIajWBmYC6Dm8Heeqq5fkrzbbkjrSYu7FL1kpSIfwEBJbuCBmHL
MGffcB7IeGyWXrgx9DHmmGqNobe90tJU0vBgu3fEJxi0Lr01wvQ2Fta7o6aomF7Z
vbTqmenMne6hElvOfCF+gMW4XfGARrQy1GxeeCAAl9Iuv+54B0E0Q6jxjO+29ejP
9c9CSRJuOM446dMkDcsW2RCboB2X3+7MfikkkWihnYn/Z+vbwdvRrZ3ljMbJx2/b
PPWMzboZWv+jZ6b3suWDq4yYNdxPmTcMkSD/DkGniyW1NkfRu1K/j6jdE1hdAF75
U8ubAxArBl0+cBJ6CST8Hy8xTIgbj7kEb0aYLjghoNQKZsA1AwdTIVUJZ0/n4aAH
2VRk7UgUygLV5CMe4funuik5HHc8VN1Ngv26kXop4RfceSiORdODz5gcUWdks3Cf
Wj1svVUUu8QqqeGeVg2Ou93I+zAbCVB4zLRQ5Jr5xVtuxQ51pOdn7laVGAf49Is9
+SBBLXDYLWMZ4JUDSm0n2Plm3UeNOCWAdbvtLpD2eJXboGxi6sA+IIO39+JtmBad
uBj/6qultQqtYpr1//xdTS1LIHoqboVDcQwIAMJQhwC/NL/MUGPGlqtnLJDGbxuk
BWrfX+uHgrY7ncgGMBHj0LsmkamkE0SogkpCKDcVGa5Hq2YKSDv8MRJpijPn5qAN
nW7zUb/W4z2XaF0RWP98XKrp8HDVn9DiAX1H/CgGqQJlKHlrxXhur9mauvgB2+/G
p8lqstPNFp4quea+bQbI2CGVFdjgXiA3NbjBQACRWR181vBC1BHaLcmVv9Yaqdlx
MmQqGNZo4MAMphuUfdeIBhAMSHOvhNsafn7LT6dkzpOfD9qMutgtqVraybaeaHgS
C+IuXocWUuX58Q931DeYxp2l+Nq6qCF5YneC/FCuXe1DQLr+ACGFBGctmt/WBywT
qMTrIxJQamz6yE4+ehsgpit4rpEA+xJtwltfOFqq2ZxGX5UvueNmVQvYuBKezGzC
1efkqDIkgPDEVIfZsuFynFDYcMkq156HycLQuSj6QcwUQ+Mp7ho0OiNk6YxdBjFp
MnU0gmi2nt2kbwGYy1MiXWtH7QmP28c5F1MzPTB6spsulkScsmbqIigq82FLc3NA
sKanpCFkl0C5XIrbgRm41DJooc5jBujAJ68hMVGLOVTTn7KKo5y2vPwvjVtk14by
a8AXa5TMdIV8F3/Minb3jnuqdL+4f3kjlkyXX2m6kuA0Rm3vh6SgRnOB5a148qKU
YigK81//sXa5M9PuqepEs9kavARz0uDjw7Xj5QQdJvb2K8d7JcZWK0ZG+JEdqOYY
8nD3zG0QOTLIfI/XCalsxmiZz++dolZIO1Do3U7mBTCF1oLDotkKBxGF8VIj3ulZ
XQp8ZfnIpMfpv09gWcwmJBE1kKFWVpVVFDmN+09sPHTvzc+glux/GqwwN1t0zw8p
rjH05v9+/cH49wCD+HsLJnSFv9riqhv2yyV9SOpGNBJjRWviov/QXP8NV4uxqBQZ
Sr8YLympS+1V3mbwe0KlsX/YOE9WtUdC2DP6jFdmyozf3CSA7PeFyMx7og8bbcE5
p46A8xBnh7BASr2QhISV94Efi/BsuxBZRk1UB9cSaAcP66AX2wL+rpm6NjuvR0YY
kg+bWdDRZ8CJ6xKiF8g/5YV/Jda3bi5hY+R7G7Bm9alvS39NIcz9VAL1IYHyBwhQ
nwoAxbkq9lRBdL/8HqAGevnuwIOW6+EULmRrQO4JAgaJ1wUJrIofq/LoW0J8PQc6
JmBYnDTnBXuc7JNLv1r2t++DFD+wa1Koy2dEjjqt6bbGtJLKpGU7+YPmwqDCIA8x
G7mKduAcNoSJKnf+FBKo027qsCn7txFgm9UE3l8IDpNpzQqPXvDB3RclGYVuCCfd
ul0yFMkQ4nkhR3R9e6FEfGsziNws0nak14mTnqNW6N497u4G6VW/twZTGg6R9QP5
picjurFa5dTh15AKgz79KySZECZpCR1xkb/ML0yEkj4C2Zrb00uDDjaaxd0IZn4G
zU+0LB6bfWfNcSeYaP+RPGnzqQBVyNkX5pAXtKsxEyAm0smnlNjCWVO4hDqoBkqh
hyaGpcS5ioC3aYIaOzPsKGz8VHFRrmdZfXR7kH9TCvjH11unBph50Ew4UG52qgZA
efiQxsRCQuVd+ZNNxqDEu/EfuxVNHDM/FKJwgDfSUpV6JI4TX+gAZqPX/FRgcaAp
V/79NZ6pinoHlwiTnMjmfvZHHxNxVhjHepTIQIxmJbmzUPaJzlOIjwRLVc2u/Y4Y
LjmwNKz0Dd+d0ML/as9zF/OgfX7cJDaQQYBM4/1T9qM47pi+Xh3kkPldr9WGO9dO
hKhyVLw/qieoLikvM7CfllAh99/BTRRhIGpJbaGiDFsfJUExpHiaGLtseZ8iXe5B
5GowShdy5pwIo0VfigH9R+NFk1I+hF4aHBJnlPFhBRRZrWTiyb3hyEpdpDIbuTm/
oZjPt0e0p3AVaCQ4f6bgtUfiM/ZCNysxMsj78fEA21WmQ3fxm3Gcl76NAgv4wHrG
t43TlFtWogoxfppgbGPq7nEeAKH3oENKjbyTvV2ttLUQK4rUcqz7GRWalbaaLUKL
ZrUctBeU2xWM28cf5VubTG8niX33yNsJHqf2lhzEtdk5yrXnxPkbs33z2GCbWjqY
WZEXWbC2mrVl3k/d4sDdL4+8P22T69cBY2NEiMUp9DNgXpL34e8U+D+TozqOH3w9
GI7AGF+2xqBiqCU/rUYe0GodEXbr2PxOheaQyzQf66kmWpBcdINFkxjO0/D7Y7Gg
mv+hlMzB6BdiXTvc6pPLqWafDdnnC5hBISYyaXtBpeJ0c9rBfpDdpmnZGWGQD1z+
1idMJ37FZdBBa8pEhNUH8kTlOzuRTHNMsJinXq3Irk3YdhkNc4UGfmfwSYF8CySk
rFHDvs//1Fu8ur+gSAGiEYvtFuGrDHrBXxdU+TzrTgqU/8Ed4DCg7Rea2Q0WLxjZ
MMYlWe1ByNji6yxtSlbyrbKQHnr5pPk2CShrqyOE08EheNqT/kYVxnce1YWDyQQD
NYDxTinLiEI8Z4sWLntvXqojDEvb4YkD3L81ldnHesgPCS3beRAb2l3JhkRFf0dS
rqOsUuEFoF7hRVf+Kl3SOOzFc/sg98lodQKVSu6Fz7eKe+M+FJvhXrBabTh/Hrs9
/hK1Mg2HadLmLMIUxOxhYw8dlUGgOknfOPQ1MgTVMY3RW6iNkZWAnozFa1bzIHJe
LCJMlQH9vCjWlMEL5qMbgnQYJi16rT1ZYV91BdjzG7qkM4uBzwsVwVOyyY7CaXjY
9QW0DIJ1GqXgd+9s9tdPJDiu0GRr72camTZrGOuviFyLaFdT+rPJMPV8+26GLoTd
Y1RsyBbAwBTS8X2W6GYYRa3oxvl6F/BkPME+OAub8UREMdRGpEuoPT1qPTwT7nEe
NFiA1/VpiScXUI4M9lXeEPSP4rOZuA4f8eNdJT91CgQotKEWAtwxmyaCgOR6amW0
J/VzLz3G5Bymw6PyvN8wl0I+zZH7XmPrGdhWNuHD9skGgIV82IejD3e471kdU35A
CRvlWhLWunwlUDYFVx4mlnh/+TK48156K21J8UGILuTZSPv8dcD3ygQ2KVbbJwkN
e0cheLgpK+YBztFBEu5ovwKXlxpCpL6H9l0hXseLIZ1R9aU16jDV75BpbQfVA26l
k6BCy5389MUa+lOVfXicItf2W/AABcj+DwdtwuxpoksUSd7k9BweFaDmBAjIyTiN
VW049EieikARo4t97OJzWUlDUN+hcyYWAQgQ+wfZKslQBKRfuxeIwt5ywfHrfar0
IFYW/NU0DNk+z5foKAcz8zAKDkjgipZyWoD9wniP8+GQsgZaVOt+o3mpilHAxup/
okVpXFQgp8p3ceGN/fs+GB790lFiUuUBKE5ZxtuS5c5PMBcd+6POaq2IHdo1J9kN
fCdxxSUCb1SMYCkQnUlxhVkuS/QWx98NfdvAABgqoIYK6bC1m7eQ/8MM9MmEw9KX
hxVZpsWdMJ4bk+PuWuHiSWGjpFnzttxrYHXVpHxTKzMnu1D8Q4s+HvVDZrmVCct2
rZbadWiXsjPyyIenjwR/rj/wlbnTt8CfEyX1GNctT4yA8LZN/9bN9i2RNlei81+5
sTRBUdoF5eTQlCB3tcgNVzMYSsuj8x4D0GKRKWE0kTQyRquEthfGuExQXrxwd/gd
zchNNXr7zUA85sjJMS5rsunHm2yOcylVkJlmvvTUzBTo6YigBX/MAkb9yJOIHnJl
gaywoynRULK0vtXo14oCuARTKo1I8Jb2ibBCOBBARmAnw4bsPkptBi4YjRKdQaBV
h0FB4mGx2pczge9Tdhk5EdA+ct+74p6j7U7Kb0c10lpHs12YxhovCk56hWdGZ1n2
TfY5tWibAY79aKqtQy1gUuSwdhk44nAYOf88/RZcPcwBNveFShgFna6wJmfUmYkH
ydH+ZDIXMouBr2IfcLMwOUR0q35Y4f69sdxDV8gvGo+XBETGCRmpl+JMazCSD8Jn
pbFL3sFh+DJazWVGHmiC8mYrecY3ziiJImOdURo7iXtvunYoQKlDDxHf3n8UaBWr
2b8LHm6NxRB5wEke975NEgr97PD3dRt8GrnUyBPkU2B5rPxjxUebn28TWdO1ehLi
wRBvGFMu/IWGiD/HO72/1Ot1jeHhaqlmRBTs40MFqwZu/HmNv2mKuVmOKYwa9MQG
qQbuR6yacN7LbmbJ//0S+9HfN0ZNZIgEpnMN+j58wD9ur1r+qWZmTnCuctfkY+9E
j4FQ82y5aJeYkazTBTtM0gF0l6sjucnzb5y1r6cfbKVwMjl9dzNozh57JM28CsGb
fo4nn5mKW4GaHit1X8Wq/CEbt7VP41KvofVUYXI143C4oOdHHAGgc4C7MVScCUEg
DLb8CdJ+VZLp1tJ07eLxLX9iN0EMihr08IVdaadwEKv/vw1lLKkOaqeIFtqO+LKi
5x33F8qqx3HnQ9FnOEjjkmlgOlT8Guuo0eqKGmhn+2ELdZ8r2hmUfEgfNzGtO2JH
pB9qy/ARFazqtoADk2CR5ntxlHIJ3PYcK+4vZ4IAgi4Gb0jS05TzsAYpsU+bdhR+
LealUn4h5KvmZrGYh2Fw9tnph76ccQuuYVn6yPfEF+Rrnw9EcePYIJLmQKpyOSrO
Uv4gJkAnmPK3be72PcI2HSUdYreSW/tyjI0OsPNWKNiJ9E7bhOpuDIVx9nZKk4HY
hViQr7eNdyy7OVk7G4pMxZlCeBqTF74IyalhKRF6uCe8Om8zEVuBLIH5MsDcYAWx
8PFlViv0o1X2NCNXTBvI4n38L2bSFIoL2+dLKXsvR5hoWo54OFqJqxjNhnQsfVYO
pq/7ZK1qh8oMPMsGwbD0ztbI2p18WFz7ieB4AysTRumJWKx608te5+nqRqn5Ma/+
cgVtdlyKwNZi7HxLkVkOafZ950nOW+E9UkguxZkRupN6YRxDK+QVQTvlVJdkoh13
UznEna6BvA2Sf70ITih1oQ55V3vkPdkCBNOoaFXax564SdAO4J5N7dHWAY7NcR0S
kGXrx6xVv0e2xwO5Te4PW0t3K2LLqdPcFFkd92Pz+QZra35iKzmrs2+WKWMDe74V
+zvGOhyGuVIEvyd2J+qRMiq/yfDA9aU58drSb0ZxNpYC3uBpuc58xstBfZXpsePE
nLOv7XQ17c71j27CTHKJC/cFSVnU66Xl9bfGv3j5KtVk9wJAXi0uFR5yFxJRo+tJ
2ARsQmqxfbJ/RIvXn9dfSeMNT4rdzFCeGZUAwctZyt9XvmeUWNLmZQ6lA6e6/JXA
FUFn/v2/0dzpnSaOJMyUmKJyaW4C5v0j3fVwKyKKNhfG7+Qe1uBYwG61xD0UWoaC
0bb2oDqK89fdFHO9rmOoI4omZQcZBg7NFiKdvoH1bk73e1o+uU7a0128/oTFn/zF
ZNY1fc4vDT/BHPN7CFnZqS87B+FnnDYgKC9emp0Eopi2yW7ZUJYEWzqonauKsOHW
wm+Z13s5Oiv/4QIhIi8IC2j5yl/eGNobFB3CNTksJJZYLCCuoF9/+7G9Wdf4NPWX
utbWShh/Ynm36zI1BNzhCYCNBe/uYrtVA0BF23tXaqx7/8AHyfyYZF6PAgL1JYU+
FVLKQy5LlKjY8JRJh2M6xnn7ACxd6yeDPjIs6HFJdOwcdcHyKzKVsu3Miy92MtXL
wH2yNz8+gH7DzQZFZSoirqiyMJSSaTNSGjpfDbrKg6LqTPU8yMIDTe90/FIHjHr5
fmM/KtftoLLGEGVociqggJgxjIp8B1W7kdZBi0c/tYpRM/mC33eK2QxCaeYb1SJ7
SWstBFrCbjUMH62H1ypyTMS7ls8K9PybZw7rGZj1daj6EFgEfJF8Pg0gc0iWubLi
l3wgsXvJNCJSiR6XolqWRsT0wQHQeZHo9IWrLg+oVlRnfokgCJNDKTAyZ66ONwXN
G6GArCPBTSi7VPRDPdmC+3vMuhj/DiSuQtAjNxaDWaNcb/R+YSm5Xy6p1YIE9SJV
Op6Shog5xLtH3p8EDrMUJvIXLaLFsvz63Kqg1Nl0w6kWVB8SkRdddo/kTEFyVCj2
Lvkv4zXmuq25UieSh9s2L4MYhLlf+jGoCeuQinGw6MTahTRT4TFaVAm91EpgEAUB
e+HAxEkJicdXO2owgzVW7NxbqECCdoenl1OqcCJFMOnlREr/kxvPCV4Lswol9AQx
3ZtJBeh/YYW7BpFXDYtLZH7ccac5ImzRmAzHnJf5VNDNUaxrWqOSx1gDFIOwkbN5
2QkXtuvUYHx+HQAfjN7jVxZBv6zZAY1JdOMuXN65GO0jxn3mKnH+BgqZQvK+JrKm
VjlnZiC037W4g+9PWHiEtGzR57QUb/YNkQeUCatUWd4CjuijNL9Hh366sFwRZEBa
UWNDMvXWrdBBmrE6VOew7MBTbPh6iYqPEwEKz6ua17vnuNxl0bcK2Mq6dVRa6Jl5
e4Ttxw1ABfhWog5JSuFMMKJvU4qUViKy1pUUCXlyKK4v6lSy5pBCGUPsz7J/k6ml
AkujXFCsDjVfN92ohZmPdwo5K2gGnoqx7rGM1+uOO/AfnMceC+Q7F60ybUHJyqoq
Cu8cdRApVAYRxK094gp33fPMdehsjEeNV2eey14K0/FCZnwuoUPQj6E1hvP2/jTx
AdavondIlmveIt85W75KHTM5c7Tq8iNqQbwuVGXFl2ZTRJVsc6VufTj9uABLIvi1
hWlN4yFa3Qx8z+PCi+jn4vfbfI2CIz9eYNeN7kOYfMMC7Ctow1r2aeneMB5zu/PM
Q/NxAJkf9q845gjOQ6qpxGojwRKqEBb+loy/iVWW1nG2WS8m7Oj568d/gL/tCnZC
TsqwFtuIMmKg4nVUcIw8N6ZjdwORo2uT5ai7OCJS5c9qshRQSVcxHIQOMDGsOt32
NyOHB+pe5RIR10ylTUwxToUOXvVbhLJU1wu62wFB0XVfU6WfaxKlcZa5szthH/os
YaRd64soJANd5PASHTc7DMfbkstn99YTqOplXgiTBEyMws4EPkwaIDJhpP7kmK/B
LiOA8ViloLL8TeKi4+WBO/oV3Ccfn7EhvNl2+pAp3YyMvF+6oMnOojOOcpRUtGhj
o7zcvOYzsJwwOsh6o6r4Qty3tTbqeM4WhV+TIQeHrqD6YzKeTuPBulJE2njPTxc1
HhkobbtAu2qOw0MOtbFHrg6n9XitsKGIF6edWP2106bwofI+Q0L5mxhUGB+JeJ4f
H0acd2qvSp0sj0efUJNo5mE0QVpGlqFyqvIFqnx9OUF5saRGJCJrJ89Qe5Qg/0Bi
PGTBKQbGoW1hATh4QeGd0oVX5ivS4bjPy7dvocfKGSNS6/MvtGF2fd43Q42fV+8k
6f9rV97S5G1OV73VBCEntyR7ij/D26naEIQGQTu9UpxkPqX0aiHDDB0CweUPwXyh
WbEAVgGBDj3EIbtbx83YFr1yc5hGJcdR1hUnnZgz22SfeQ8mAJOcXpjBIgGKe99x
ul60CrnCw+TlMF+WZsey2MKIrDHuzy7hcVKTGBqZZuxFm5kvGST2NIkEbj4CEfUh
S9Q3cahtfCQ+E2coZxBM6xBij8ysOgTK8ygn5UsnHsYuXv1HPbVVay63qBcrMw6x
J5IffEwXuXWE0gnGvQLttN9zoore3ZxeocROactku6BLYR8lEY+vwNY2ov4eL4Aw
Z/AfQTOAyGaQWU4AtixdmQrca8wINiDjSETbbmhvKsqD6pFthkLWjiLWTMkxjC+K
hEDTBdkTC+Vnau5JHdim+vUYf2rl2MqNG2OthuvY2dVwE5fzHmMyX/zIvvyqF2gk
Ex/NGn+csPUU/m057883MssVP4jEiwqDP6E3OyypOQcAO4yZHexOApDIPISQHjAN
rIrHW3aUE4wX90nJORvFZPwvvi4H1Dhc0et+Hg+J8rQYSWxRhA9EhBbcbYrdRZvU
HVcoQWraI2N7m3MtiLVlOwJ9bGcEuP7JPDsODEuoFWsjGVubQZhzu9vu5aSJvdFj
krtOP+MYWvWWJ3pfteDfDynxXxF7y3exkM95wiww0Cak4i+EoSRYEzbJ6LdYWMnY
06EPPDyQyuNbAy0RFkRhAbZjZQWyCV1lJiJUpOQE4yd6eQm9rqOp08l1FKRMc8bI
ngYx4Xkn8zoXi3ABNsDWWzB5OBevfz89hSA0tQoB1dQlvHhqmAHo3se5EGF8sn2m
9HKWM+TqVVFAdWeaAoyoXI7xST5OA3F5IhEFb1wDHlL+wKBvvBgIrDaWhEf4mrWZ
vYab51eG1JEvC/vkKa7p/QAtgR++yDob5bv/P0syXk1Esu4in4pJdvXrxhBHLsyw
9CAb3KWkfcS/CLlFa+3tyvC4jYEXV2CnxSwsviTCKqJZ6Lujm+rZMJxy9vIkzV1k
O7n1owBkewZ9Az2RMZfPOIsRvSSea5HxbsKhN1mE/fsXu6MgMzFjx66rW1k8PFsL
hOzegjgFEE/tOb1cyOB3nGUw5irooP+VWWLy852hhV6GpDKWDeQioB/G6AOg/uvr
OgzkYyZTBOIBxTC3CyWOx26lcHyD1NfZlRa9uCKMHTpgAFqbcpRKetYq7maPzDFL
4mG9U8sV0rZrFbN9XiFbYw13rCeddswgvPbKn/Krmy6VVcLCD1EAJqPHAMmuPhCT
wRnMm3K+19SenEMRR+dKvbbKycmtivnh/DGKAGqusnNe2mBOFairm6tbwhrpTRDM
v2f2y/zzJDhz28wHkUmWHOlQ7LcRTMHOwF3sotLfiyi5t+mO1l66RNb/GQ9mDgvh
KCcPi1mfJBxDXTCPrKYr4jeg2LTi//0ygO3ugh6lFwU8TvRZC3faV3YH8i+iqzMF
ryrOhGy6wrJV90xT0bB1eIbIyRZu6AoB50rZjC8Jalz19U69qz4NqeEbTq0kFIZh
avtiyECOQWbcj2M3UFrPNadhD+e/r8uGPEhEiZZuMfDAQjPm6RSkxy82PiU7tAwH
YmiwfXc6A5aH/ln/Y2PQG32Oq+mYz2UdNgCpQZ2l4oBlQ5tM8RYUyqtLovfjyUfJ
VFfEgzqGKfnk9lM7JfBoXWWk42Qt97jUG98FXiaWNqYNuu3Zj9gIAfT9KGPsn+Q7
reNCOJMITuvT42f04sc4o0w6onCmhnuHCoxjiuFQjG7xInU3FUlrPlgvcQXjOiy6
B67LASpAVhmrtXOEo0ZkX2hHMj9iL47rCWzC6k5TK9V9Wa7jemq+cx5GLxYXeQWs
t0QkVbFRobAM8V0vdi8OSWCdouc9MP6yC3AoW56uAZ6iMeXwfst+ai/XFFSHgX/6
wqsSO3vA9gVWR28UhMn3iRmQcAz1GcMOTJb+V+7rKD+NkYQ9MNjAEIhjGFxqGytK
WqVJyuO+rI+2cOQslx2eFWxr/UuLVFVbgYuFh6Aov3n5al7PQdsQq9+dgBmhENpU
2sqwOzPlwsbKH92azVk76sWI/ACULXQPbUuEs8kCWVLBHsumEKFYmdCpjU6bQRxZ
/GhpxkQIIIFj0JUwSgr6mFsNjz9umqqd/1tqWfaiavsC6I6R5ZjJirR7RjqBRLlw
Zs1Px/jt15RWb7C7/AlDj+oYFRMtXkIqfFZ/Jv8ju0r9djUWMrGaSgPz76L/aR4T
n+oErki4ClQtzYKOlSOkaTVuyi/MlZ/9PZIjqshb5MC9rxpB8rsWpoIoBYIcudBz
wzek9iuXhsWfjukzIZfyY3NJSR9CCtIzI8f4CbzEPeXtGMevWgXha/sypXIM0/2c
i4EqJqV4VrQ2UrzckBjd7hesmH8Eray46/WX8QO6mMlK4MWYyvnYBRh25EJMGkXR
gbThoqSx+R5WIf2GHeKL0OCoFjRa7/HvyKP8ccLW+6aq7zK9l6WxLqhpJAq8Hveh
U6+7BDqFqUbtvj0AsATH5iMZntZy1YC7d/FGUb6vBBKR++srDWDC0Z6jIY6vyXM2
3zkXMxCpUBEJIyuAlweE25EbWCQAEm8/i+25wO5esk4f84a6oyLbhkyvusw6UoJf
pJnLgSr/UpZI/jkxVmFwqft1Dn4+RpD+20gWForXdgenX5mSlxscaPLWTBPe4UiW
Go3Z4lgSdJtPtTKxuPrXBlpo3zc1ggDU1B/8At7IRl68/pJFONUuqyS5QMFR8jMb
764Jq7rm3QnyCu3tJY8VTixdvhjBbyMPJJ+shOubwHIayTm7fGNFq25haSJpO90I
ZVyPK+EIjCB0JcXtiMW3fAZqbcQq+YuO2QPVfkngjkxIc6i9TMpeuA0lXvIIY00m
IDy+43fnZqDgd41Vcd4kBJmxv9TKWABsBIhk6bOwsl7B9V1McKkExp5G9zAbf+Rl
xhw89XRH6D6vnvIwz7bMXz0ZBPhDy9rRmRMj6vH1AKq7lub8JHW00F7pIUjiDdHz
A5uZspoz7kOvuhfPdZTH21BYvG1WEFLqZQAkSfvmsISOL+pZep13eNj/kW957nXO
au99SvrCZm9LwypvKvcs2tAX9DsilEICx/7SNbjC0gw7+7HK7y+dXqyotenPzUdw
aABQS2vWe97GWh5QUeKZWh5sXaVYvlWt2b2Jgg3E/q5qSGt/pAsv8mn0OW+8CSmK
JmGTKw9Ple4+4h/DOafUf0IaQss8hKmxYloB/sq47Q1XXEFAsmHfqGEvzcygi+o7
W9sI6bcUqQ1LqmNRN82mOikVT3+XtquPfAadJV+hzYr3H39qmcGU1JXushwLhH7q
jvpGbf/OyynFNYaZdiupy7cMFC6B03wvLFwSgvPlox7QyrShrdqLDf2wV2Tmor/A
lYjxX+WmIeziSdIOn3BcwcH6bRS3ULKLGnJtvkBUICX7Wt2UQB37FpGSD55cydPU
7VlBzl87obkDj2XMarjsFQ4jXfeCHEOdoYshA/90O6704/1r4SxS5btdJoOvutDH
XCk2TqLZw4XSbmmOL0v4GPK2Bs5Tvpl8bKuUUDzOrP1vQsu3jzXULSpPWu1WTjPo
YbPigARLQPwWDhig1Laec8Ka2aiprZRr+FlSn9lXzYrV5dyXdaXRHCJFwu4mJdaD
u7DfkModPq/3BBUuvUpe2Q7k3jg+xl7jIdAmbRWuWQWdw+SqGwfvyAKc7PV0JZOQ
zir9rLQUbxDnqfdAuYDrLmpUk1HfUMo8051vf9TwnM2hRhmX9Ul0xBFYwYITVsHQ
pfB0AjfOZhnjiJgFJzPkVLyPhvYLL8tfjZ3uGlGOuS8k+7nBxm+T7yV0vY1IWKjc
JfOrXfXvrt/vMHViSOgfpJ7S90NkgcPyZix4v8knrSd58brXUygu6CIkRTt2ALjb
huwikUzoATLMAFh/h9rCLHxYNZ1x84Qcwx1i74CCTQg7/CF4aKqw/1VB0J54DvWQ
glXOv4OmAMW1qHU9dk8c+Hz9q6sDLHTMspfC/mhd0UjKmXMUffkBIoLb+6Jr5oLb
VVkLBwFUIBruI0QOJ5NPs9k8Qv9F9i6dzxTiSpD/9jNsUhHOkJK3BY7TWJ6EkbA9
El5tO2tYfzA666bAH6qYvDx4qShj+nVUGKZNEJUKFTGVvEhs0hxVdvwOqX/RvQzN
2iUiXdFQbLjhpqfGbs+0bOfMqw0AuapDMArLz6/MywWDARYSM8PsZXi77M46eU0e
BIGVVAGuMQmlh/HZnPygStr/nxl3PDktHx03jv90ulIU/4LXEHJlFm7OLjU0JEcA
9A8q9Npm8PK0Iks2pQ/nVy2h+ds1fTo5pX9W8Lc4Q7NYcyiy+oZuEkFDSLCqxuEA
Jsk+uxvKUcpHxJQm3ca6k10j6QdPd05UHo706no4vIA8yb1ByuzBqmlcXEysbJbL
0PnfEt0Cio6gMhz4CBCfOA7HGhNEIZeRcXqY6QIVdx40rcjW5q5vIDSZAbjlhEGZ
Bb+xHE/DGPjWdFdp1eNQ7MK5lcmSRwVCFnQGBfDhXD3JDJhBcQ4B7Ka6rWXj/LjD
/MCKCOs4SilJXmB9b9TttQEBZcuzQMergHxt26yOKEKqV0MgrJGkOl+cMzde/d0k
LJnG0lreiOPnTpNFk2w31+zA3m26bY+qrFlUZPiHTJ5QunG8KHuVAG1hOoQ3XbH0
W6DIs80j6X7NNQP3+ywgvVM/l0DEEXecCMJta/dD1P/uqoIrCngjCCOhyRD00iD+
Sozm32444P1wCU6ESMEquMbaXsbipdecxfGc1orNxOo2QTOCExPngslH0KJu4/aI
tus+PILX7O6g5vy4fQoTj5lIBwVf4MG2THHkuCuj0UWxYWtpkMXQKy7LNExkK8FO
g1msQC5eLLohqc3fJq97aI6Qcgnf1QZmw6owmOfrmzIyn63PaLfReT3FN8jqifkv
UZAXVI9a2+ElgLvjQWIEbFhZexVMlYnkBLAGLMEkwsavkTs7do24SYSWZ3J5WFmc
NebxLWu9mFqoc5hJFl+2h9HBCJsaHuOktEAJtbLEw6i53nbKaNGE7hm5sD+MMksh
erYRixb34rFxvZXbVP/v5kQ+xxDaQNn3s8yIamZalQcQ4Z59kKOlYU+PCAJuWQlS
HeZJm/68l+dV5dnDSg8T4Kx/StfDEuq1hQlibRtPIToD01pJxFrAEdrRb1MhRF1C
xESr+CHsK3Yq8o4CPPoDh/ozfQepR3uwQztjHk5gYSZ3QG9PlAPZGufj5YlfKj4H
a+3PaQowfexrxO0taz1cRK/pV7dkG9r4KXSJa21QHb3UnsPFDQuJEEDGQ8HTNQbm
Ox3gR4Ll4Z1bBnR9rmH8zTMVEPJ7ahfFa8S+tbO0Lm+5IdbewwPWsv2gmMkpy1PQ
4Ejt95FlXh2x2L1vv0owMsDoE8B4e0dj2RYhRttfvjMR5RB45P75Gp+zhNum4/E6
ikSkilg98h7PXBORKWd21TpsMqPfuoRF2LHqFDEbZW0/gJYETE1bfn+SV3qkgX50
v6rw4T7OwWJO+9mxQpFVYJ7LRv7ZtpmWi31zWcxuhv7eekpyN4+YnCfS982e1mmp
TmQ2V/1ifDZ+cUpUwPAHigCZMJI7+AZglouuv1yzW7aTwK9E/7WZWK+rvOXZASj3
zFcVVujcIa8Td8vzlRfaqY2VUOdoF4fazaGVcjciD6byffJu7SP17KXu0CvSgdv+
e7EqTR4oO1ToQCuSiIK9WCbqUaMK8nJm2f/N2VkLgBxeVxR2gLaKcPos2rIcGp9h
GSB0uoc4FHAiPCKCQvZXbAbz85PMyfrLb3EbCyoC/yIk1cXyPt3ee+vL/g7WbpPe
38+fIFDe6n4ryGr0ononrwc+vKohfm6Y3haAxvljqzHBrU5DpGIVsTfAViR7jk1j
jZLc+jrfjDXAKVJsZrlqOryQMaPH2Y4jsHmHb7IRf2kJhgmcpIW9DIT2/bmJuf8/
Hn4OB5grxHyG4VBHu08Pw8tI8cuO4NjzL91QIxTAueg2BGjraMk+c4RUaSLnBGZW
Ndo44A7Dewh4OLp8KxVq5UIx6uT67TML6e2dmdtBYHKn7fdNDtnIKxrzpQASupmE
QYItiw1Bdor24v+FXQe1bFPr7ekb7kSYGLoLFYYh3G9D2DegxOGVsg/VjBXjoj8t
tGE+gLPLb7G2PxqcKDqBuMeYEeDY4fhghvKBsVOexFjC4ct5zmJi2Z9vW3rGkqhW
jKF/I7JUBgoy76qm9nMuGJT1j/C58qx5lHUUEW9WHceltx5ipN4GHFc60iJyLCdJ
yR9n0C9t0F1Ebxh4a+ASXHk5Y2chszyBlLRaW/WEsy4ofCjOw439V/QhIpRpxgQs
VvSJ2gWqc6WjuQhsLw7TLMSPJMPoKsINM+drrXPeY91LNHg1gmhMy8awVOXj+hba
1Nw4GwtfWtDBWLmGZp2FzEIk2JsA9RSa5PgbbRF2FoMhlrIRxKqvA07N4Kl76Ox+
10Onr/22ETFm2AoGR5Od67a5sP4cHzUDeR/xkZxuRLYgdpfX+DcKmdOhNdwCz46D
Z8S0YRXF2dzN6KCfrKT29laHE7xEV7bkAaN2+snBnF/U163bbsXgfaGYK+kddk4g
zYl0mtU9zofUsuCBKlilXhlRu+idQKQTW/syDeA/b/+YsYXyMZOu6b8YTwhU+Jp4
7ZL1I8QyZfAt5mQ2+QcA2VjewxzeKFZLtHOf0z2aLRQnhPI7SdKVlZEKYaqB3ycN
Frp5LVQRZ/7VGj/XF9UxN84Dt6MRkp10YZOHq8F1V2P013miJPFmFqbVZc9b3+g3
7FmpBV2bYdrMqg0SgOWdtCGC7GIcF01WVEBGvduXMlTYp2kEMnpQ47qhejY5cmFx
as/TvOrQO/ex+ygAodtYqjVIC7oNNvAQV5m5ibIlzeuZRazuXg3WY10s9CcqQ2bT
H+cGzqNL3rGvuzEmkHgFji+IYPAQGueJLfnOXRi/WjTLEvDaTBpS3l8ifkXyvel0
Vo2BqK/u40I1qi06/5QNoAabuz5EIzHoCl42cG8WXd47h0Ur7qs2EHRuLLCXVwVN
vWDJoqbJAFmcCWyMFPC6yB50LDTok/6S1fEANPM1yajPXt2w2Ou2w7uGP6j43D7l
1kZuYE/I6gaRnwAYX8MUpMO4yQPhcBpPM3s4w6PyEWTcIllHEzhMVjrzDMkMaWpP
L/sxWwfkVjtSR3d3VATKVDA3XcJeYbnQa1LYKqQKM9jhfvntET9q/FWfZN0h/Uzs
lYYGYHRAnLJrqhjPlvgQyBkN+PqO02xpjLVEouKZzrlqeSuJF2n0AtB63Qai2Yg0
JexOEZnrBMcocacp3xbh8Zn+zeCWwafeYmw28GNwhk0vycUbTVtQoEeG+/uqM6K2
Krx0FOkvowawmqom66XXwPo5/6de+FbEJm99sxJ1NJhSIZIOZP7PVdwOYn4FKr/W
j7AzJ97CpwV4Fza96BtXsz9GmbhoQ3mTPK+XByjncMJu0mqPN+rA/7rnosOHjjp2
cRRDqW9VKbwJ1TUqvBQT5EASyJERveWe6NzUn5B5UEfteWuVgxOgrsVMTWlFgtVC
V0InYtB9E2C54fYEjoNP7j5M0d9IweZ7R/YLrY2evrFPR6IdxVg2z6I/t/MzxjTA
GvO4LKnf9m2YL0Q1i0Ij1falUDcDulVmzyY4pnjIIRvEt9ccvAbBuq0TaY83i4Z4
Vb5A7j3pJPi9IGnY/jF6EwM8/HyuSyngMeprcYnl0FFb74tu7Z1VibydNShdr+jk
TYkpyG2cBmcsl8idZDM7D1ExR3LXo4VIbUkY2H/p2wTKYQuzQ1b7I4UFskezH7YC
8lxj3biiUvUzOAGdjD8AOQP07Ey0//0Zqlqcn+iwYAMQsoyvu71pa4SHNkRFI4DZ
zxWQu2LKyRifewj1Ed5IkPa9mOhLWx0P1E2mObJLXqF4pTFGta6lZq3U+Wcgcj6z
coAzMido5H4xbm017uqQLUsQ3vLNvxtAHMiSlyp2Yc8gMvBy/9hiWzgEa3nLXs+k
b/MMmWPUVNR2n72FJkxRUEgYXkCmasC4CFEtnThDEOGkw6cVOIdFndHmSJbjRprW
KUy+DY3m+brlbTJTOw1+lGSAWOp0+SfOMgwJeqLXkIJFVSXgmrXmcxPOK/GkSsBX
AUwPKNnKxC0rKDZQdHdxBxRIth/Ycqvo84SG3XXd64qXY+kaghZHGd3miqlaQCA1
t1+FYs6zob4R7wv48f/sGDDMqaNvJtoqm5QMivgplQG+xlg+KQ9MRVewZcNcAT2r
mY8Ed9KvLFv71r/J0kzyXC9zRePNNcwYERrho6z1zNISoO+cyjkEm02+EOPCe3ay
e1UNqTBucze6GK2X7XFdp9M2MbEYUYkEwP4l8JlWPDdN0Okl/itGamu++QGgvoQ6
5GEJhJtjgwvzSgoZovV+aH/RefK1H57ylfeimmM9mfzt0Bty9sl1ZmC+M4Owginp
V6eRQkCMyXTHTomoBCpnvWdGlqOJigWbkI8OUNMp+wKvhE0X9NhR4FSfbJ2KHZEL
fPiJdE4wgoZknxewePus2ERSgmfwN0cVgU6yyRUbiAcjyHGq20+BMhge+qwOyaMg
O/vmzD8DkDnIBWwiPIZQdWmS9A6HXWCRJClQDumbNkK7Pu8xUjFX6E4AX0TfwL2L
ELZLb+JE/SOKUufpSsF+chT/0RqpPt2xfvzdhPRsYgY+kmMMgO88iJE7BkBNbdOF
+hHFiJAchdTDQGA1J53fOhS2zEpupSHnR6Wc1/kbTwDenJ/uJnRNOP3zO+MXmx85
zXUpWgi1EA9kDc3Dkz64W97Ebzaymyy8Rqf3BlZi/7nIr7a9ytBdKu+brhRrArsm
7q6em8pTjQ3x+6BWVrqkDoUgoMUT/F4fBHmOqOhMGbaJ7fsMyuPebhliwoiueLKN
As2PcGVUJVzu+S6c0Ts3OOPaV5X2FnA3jxOjtI8M5w4yEU5Sb4OV9rmDiujjYCir
fLl7jM8KgnQD/R6ExsIskSJ/gbJkH19Ys5sqrQAYNgloq1/RI6aD6Jsqt/SVaC9Y
qwY5+Hv9N8Jxv09JA+EwU2EitGSWx0W+TNBwwmCqxHj7x7MUBMCVimzhKyF25oel
d5AGHxXSvrDXPy+77uTr9y91gNQaCowvWm6rnVCO3NH9I4bA4XBOm/8BcQrSperd
1eVok8acBZv0prqD1oEhHYi0ReK+nf7z2N71KbGY87TEhx/06EM4a264rLNaYhz2
1X5+W1QvmKEJIw6v0IDKPaF3u5a4SsG0n5IaI72IwIPkLASLgetjY7fYReQlsvRd
uke70Jscov1+CGOFt6svtIUFM0S/jWy/+BoGHFui5KeRf6A0DOOF1sKg8r/qyBgT
pb0EUHW6WkX/n7NF/v9y07hQqkyxkp5JFkVPDzAMoboz5MvHKEJxfm33tJkfgvp9
eMAUkkggmi91ZtWsLgAmesj7Pn0S1LMGaCBvTFoIO94VtU7GYkVdtorAJyncSTjA
BDAC968FjnGEWyMU8eNVq+3Ye1bCNNxq0qi2wsyR1hu/6g3NLTMBLYJ7w1hOnhaW
kz2Pi1YOPejIEjzuFA/8rwQcy81HM70bkpuKlCBnSmr5ayHqE+/L/DhtnJBOHIXd
tV2qKEKhbspyF9hXbWH724cp6dKw0LhNi2ZfxCNIJn7KUzt8KCT6RghL/eEOBeAx
i3JxPfiNp5UA2awy3q26kqexdixhkFfAj0RBv2aMHxhou04C8JrVVcQHK1SS1yUA
ssvCiA/nXgU+iw9L/s9lo9tSugBixaZEtzHA5/I6whLxAqjXHpIwEH+M9X6VM/yC
1M1zS3Fsf213dr+HAEjzM53rLQVWPpZbQyA1vdur3XrPYcdR/I+GcR/bU2kA/PgN
8FwWkehkON2DYYbjr65SyYs7HrcDAcsN1fNES/Pftefd6UqBPxWYhhyLp4Zg890V
48vL/sBdJ7jmskWPh6ZvcE0RcC2VcACB/vBHQOQxghhYldqHKzs9xjBoeudxVX6M
sgJzxAPoi07eOx7LDePRgslH6YJ906zAH/6jh9ykt1u7Q/9oXhOQzsCUq+1W21uV
Cj7YP+7vO7Fjj/18g6+YO4npKsOhfK5suMs32xXCWjScdFmtHtwXAXj2JGegLj1T
6n3Nxp7wrslUfVdbdxWkXC8om1MNgF795X7egEfccaWHSsFwpNYYzVkyNux3bCFW
TgDGNqru6iIDXLg5TiwzAnxvA8RHhxYaVJ7CAouyGtJvIoakk3fgAOawGz7vJ5Mn
89xhgy/ZTSu27D7EwWEpdgXpDZULAXA972N/OOZ0VeU1els+ah9j+hgEWgFfuTxV
/4lnm5AU/RnvkeZ1iuJTNg0co7jB8TRq1RSW67/N4SDcUmdLDY/hlSl/nu8xff4R
AVgyyjSSiJjk2y4eb6uIHQ/W9TrGNnKUw446it2rBZNO8++vxMRN//GiEEMqdecY
x8pS1sLZhU6AGGTh4zWPJw/CHajN+pF8P/MgBtDAYDUI/PViWnS4LzhldGSWc6RY
fkPTKyDamDL7O9Ym/TsfE1HzgjD5JxK6NGePTuu+290ZGHBGAzhn9h0xSTb72W4t
zvlWB/IvSgnBRP1LJ3HwWAG1KfRKkBzXnx3yPAFiEIJZDAb2asxn8k6l6RW3QreY
h3lR9LPTXLHOTI8VmDcT5JiSAWWiCILEkUbI0AJvKgUlS33b1fTmETe8RmcqpLbL
SpPVMMHnLo0p2pjmTbfYARqoRB9EUwg2X/UOPGDCMgl3LOccR/C5w/YNR4VcCw3w
7J/ADguMGenB12npJxaATGOzaRs0+kfU/ilSuuyH9BrjGhr9fv/Xu8ZvHnyP5+p5
YP4cBIJylBrbS9vPRv81VBtPwziixNg0quk3iF+tWKwurCs6Zxqt6er2dA2N2x/N
0KESveTJrF7pKottFl7BxW2ZJ2wRAFYFBHXZL835XZJkd0G/0W1QAwf+qWa1085f
IZyoTt3809HgXdrybmOWXstYutbQYC2psYKt7afswZVYsDj9e4XmSuzbhNiI1nQE
vfOH3A+MsB4RyxZJJ/T3pmxIOq9IMg1pESYOcrA+oe3knMAsZX/hbnJwdncsxYbf
x12sFcfwfGV7DHbPf2TbS/T7ql/tIRVLC4MTtfXAEEwmaMj8CE3JYsgwORUaWGZq
NXKSU6x9R5/+cSX3RZ8NpKwKLvctVc0qCgdgIWkW4XFWp8ekegcnXa6F0fMw/tpP
2OSCBI4oWkqA6DMlskQAZtzobZQYWRyQ25WZlZGnbspp+kTgEnkaV/uK66tq71NZ
tK7rmljnPuXnYLIbxB/XEQTQFGls7/Kn7uxxVqGUNodnQYsJcZ2fhhfPFR1T2S7J
Uc19IxwROlSpBtrfeeLElw/p+LxZCYqQpweD7iNATf8SOM6HxTXF0at7L36lVRde
LYZS83ZJzBsr3Zeng2W1hyw28Md+CTj8lvmpLuni+BzxwjIykBD8SYuqy8oiuPOC
ZnphkjyMT3j01m4OzF6uJOVzvYWMpAjot9/tl6LJ1zHW0tzp9CTQ7BkU4iB5TFV1
wMbB31QYCY07H6YEn7ROFIdQcXm/bN4S+3nXONalL8y2XiP8kc73XxVp7lwpLgZ8
/loiVv/4cBm2jnFttpHMsFPvUQ8FZn9CaWaTQt85AYZEm3dkZ9xlpf0TGQX2LSft
C6DbqnnFRA1zCZDGqhoa/x5Axq8jItJ5xsJvC4Ef8rWMASEdtANptSy9Nv5Bqj7s
N+ggshhGeIMscQcbAsQouL/kbzALXCXG+9iyiOGBSc4ImpCShHUhxdlDQGNiGDmK
OfmLJrdcKhfsib5baGVv1Acb9Adi9cpUzz0qlGhRw41/reuostqS/lVjjXJ3NHx3
tpEMstRDuZB0ryEKY/TTEeBAZMMrHGDEMS7oxXIunUErH6VLldQB9WNsMrwJPyNv
9O3DSA3arUtckZPDU25t88D09xpxwNig983Ud1oDfHYGHyNhRutH6A4GR1qctKv4
tmuVYYmoTdv9sITVNuaa+DoYldBCJqwDQasxm/Dn9gwdNRG5Au5awN7sSwGd4qVx
a4X4ZuNdFnobXkoUg4OqdHoCJRkvs2tinqBPEGhJATQ/xxoFBwDeAS/sZkSITgqS
qQamPp/t5rScyHjiQaZw8CmETefwrb2eRxYETz79DNA3SdaggJr0kbGtVOqUpelf
qjffzV3MBgEfzzDx3lW6Igk8QtxStsaPxP12TziSJnX/uC1WafMjASO2JwaMT6/U
b5bB3PbK+PdQysv7GTIe758oe0X/CTDXkZ3iOqd93/IeLxrRKA/nDJlkN4r9SYHZ
gFF1QoXswrN983P/HYfgKM6j5umkkpWynbjVVfKFqtbM3PkYdODhpwDO/v4DZvUI
Ehw/qPBTbquwL2Jp4Nx7/4qj9PaaebAN9vEOQ8QYO/54DjqRfBcLFjoOGMCoZgmJ
vxJ8NmrE6i1Rwf3n2APMeRlTLXYG26WRMghy1K5NSQkNF/3XyRjf0lhPj9HWSiGt
yd+Y6oYidq3t7TOkWkJsOfuP8qaXeYUcjjcXOHspK1JEqx96e+GB8XXBHji7rqdX
LrpE5I5JB4crwUnVNR5iw2mCiSNi3uJPgkZhUI6TCywIhLnTEwMvgWNvAeZMTs7u
TZUTT20RfZ5GtpAv63Q/pQhpj19xPe8bcT0u9OFy8E0PUL6IRa9NbeVSx5BMAB8o
mHZ+yqZUz57kb96iZ4MQ1u2HLuO+LDVSFi5g1121w9ggKSfiRWP/3IYLZGC5YgWt
Dibpdj0qXPMPpTn1AwgjRmm9XX/M+aQs7Qe1/CU3B8EMsB7YuK9wpyObOJZYSElS
dWsjtUyzPFQmX95B0q4GI2tuRJlsmGyzPRbNk1EaMyeSoSDvOEFnsMUGqx10uynQ
nyT7OZMjE9EYn8NVT+YnmOduOqexBKsYOoeGEMSh6bo/u9JDBwBFSjRWREJNn+Az
Thb5XDymYx29ibzKlseY1mFPQcDrT0XGe/tVn18PKDvTVZ6EgqJFfi60zwEBmxpo
pGcsV4a2QdIj9x7Vq5KnX+5p5mPB93BJEweMeJZFq1HtZac/BxWNlB+vuMh0PoMh
aj0hdIg32HGcvMq52xnzJWJxT3stasLTjA/Q0ScSWIuNpSn+HxEtkU13IEnCjzv7
/JSoqocUnkipGXHZtJWkTlqI4IK7AVyOVF/r/reH51wzpX/NSCfrWgTyuAx3qdHp
QF7wAnKa69RlBNm7p8mez4y57AjufkP5Xz3Y2Rg1/XaKw0PavjTvR3tve6eoU0pc
tYGvsfY4OvxnwbTXPgPGf+Nl4cXL0WHZRh3oSMl9ZJqazU2jMDwrcHX2pVX2uUco
Otrx+fSeM2oFaPTYH3AP19DK8XNbEo9CluqgzoqnVEW5XW952VK1tq6Y4tQtHT6W
Xpm0dSbILG248M2g4/MQQqpsDS6s/qCSwUDzmd4peVpOOPvHa7/10xuuso3e6hfb
0nQ57ZBwWKTgZaSRueX4zw23YZ9OS09rhibpY8rlquK3mwD2gIUtk58NmOghWblj
UKv7XzrRFx6h2VFzgtWHIwOZiTt5ATGQCeQoDLdqC9Q6GC1/lvsKkbDmOn1UUxzF
BquvhBnXcd6aJIWuUVfxlLZQCuJU1Gv9i35yp/8CgXEM1OtmVPC83yRzJzEOpuJa
qIrzYsKPvgjrf/VPJXk9WqNPta9aX52Anv1HYUw3BkGmxhJ50Dcjj0keiGW4XjpR
Nkaq2eHo+tFerOq3oXJYW7PSdxhTWmM4Y1Q1WtW3r/R+6JR8BuDq5gykXCHvCG9a
hVx4zxVuM2z47jyNTSxGUdCIGoXEuH6aEBL8UKPAEbKguhu5zodusLTOk4rxxE34
bbnF+FvBC6Zw39cW7qa/CKaAiL3kWbcmg9Pp6FLNAtMRWYgcLqZgNsck+5nDGhC1
NQP0pgGr2NePvrb7hs6HDe1aJ6hNllF13Z9cPGVdsdnLFWgK2df4KM/na6gPxmV6
+e87/7kWtvIxDl3DWsn+PhzB9notXvm+PgQJLMCH91ZdOppeKcfIN70hGt2wuu3f
kwSPtvpF99jY9INRFgIgbqLALqNuLJoLe2lmYw/XPwjiyML8r86rs7/+fVx4NjoP
s+punYvaorlzrHDGGD7wpiY/mr1VbCKi2CVnNV+crubjL3HmuJKYlCcQGRX0YY9c
tzx2d5V7McHsVHa/hSVN3hx/BiPChRuHFY+twOpj/8dzvQ+70D5Hvmw/OhtWXRDn
RmX/iACJ+8aBzuCh1udJFteTNnLnqOw6LxMrbTObAGFlwI3yNce/fVlYAOvd/hR7
fVgeH3eGCg905piI+TbcJLGk2mCfmVWLDs+WRUigyVIGt+SujhSk1sOv3tvCs9N4
nJprwgQCt9RGTSHzwhLwQmVW/79m0ZQfexm4PDVKfLOfssiME3XAE8j3F50UXYxj
pz0hFFC4Tdtimw2dBYIbR5t6pwS6T/dWkoPLF9l75mzRZRW8TY84GItcEEnM8fat
IvxQmeiCnQkP4oAecWNXHWyFXecBEAL7BUHnE51T6fBkwiicC0Law0DQPcvLcY6F
zym4SF3zblVUkIvBeT+T5c+YVc3QS1GcgiXNGYT7HyKVcgO14qa0POyhfAh75Km0
mOzkw+3M7JZ9dvcAJXiRtrA6EkNfTLlY838JcjAmSovQViYwhKJN5UTO14Rds835
Tgr95kjKnMPUBTTDPT0z0N/gAF+No4R2fqh9qNsPgSwja21p+fbjFj7hmc67RNeM
ekhpLNTNBnThvuEVfUwA8/uBcyJfyVhw67wtFZNYn5sAz3fWj7/zrAQvL0gMkvg1
5j9q04npdT1FDApJvH+5QS3mfZPF/Nu4C8RgukzaYInrR64/nR/WtRoUk5Uxtfev
r4y1wAkD7MzhwYLUAD4pxYg/LQqiY2rBSLZvCwbMJMNKY9fOuQpNokfzYpEZz8wF
qgohydkigW15qBczRhEveonaNlB9u2rFaKxYUT56Hz5G3JoBFM/hNpVWSe+QE4Qf
sKfsTkXqCeuSfuqnrno3vHCeEHn1+dXrgu+Irq6e3E2iYTwD9U0lGyOMg0XyXrsj
22xmXNEvu8Zm0r/UAd7onuXiXBH0oLtE5+GU8SRE7f3lIUx/LJeG99AL1eAl/imx
qDJCy2tlN4VxM5CXVyRRIYRQD7sWTfn6AEO+LUizhJhJp7gNshlTqBbyDb/d7GM7
tCg/dB47GoSNBR0m4lqIyaMLBCBXBchT3T46eZGPajx/b1wOQCMpH8x8tgtBHSdm
6G82b+06eRJpSWSPriJC3N8+FObeKMBT8WoF0pXKAEIs3WRm51yqXhGonPJ88vAu
fX2i14+Smso5iQbt5BQnZuTb+kd9DyI3r2XWG7oK5RlELOEZgJM6FCqQFtrCJFA9
nf03VtVjxKNszN3S5yg1Wp8KwAB2KJmNpku3jQBElXCl6rQu1qq94ml9Q95ZwRqV
3LyJRj4zaFx4A/gVIWtzTfQoUHaaR5DhFfElv31I2DydCt0J2ma6wSae0iYwF0A8
0DJkFOmNezl5JarFBwl5eTEK6JF7he9f+K3cMT8uRTvtOsVzSCKzbQkKphf/xYFb
zvx8IXRPnb/wbn+myaTKeu3g/dZoPwO+wa010xNKhYqzCQ53n5dbUokiLiQcYNeM
H+kwbae7sAoJstbJ6PMAeD52peEUzpxfX95gR1pnAuZSMjdDU1O7CYkfnWuYcOPp
LT/CiybzOPrCl0MSYpDa7y+7rEMWdlnPkU/DA3k6fRJWEixCi0KslPurxYb6GO9j
ZRAWNIJAVhPpA1v4SKSUwdE/Tw7Vt4aGepfsyrDOxneQDIaOsOFMlukSuTbqMEXq
+3ldSduGcEGXQNQM6HkWj227aPkUJ4hBDB8LRE6nbin1CdCS0hGm7d3W1axx5NGe
2g0yKQ27Ik1K3Xa2AFkTnTMdtt4kA7qJkio/PBOimNSL+Y6gKkpGpDr5NwqiopcH
X55g6f25Na+NqQwl60SwN4MSCYjOBVvlKtzEzxZRbgvtZQP5tmFL1a1hrBaDM+jd
YBMGdASelfANVorxfg0SJnEJ4g+6ryrbrIZLdpAAYiNFrpRZh6Z1S99UbvYvT/+n
W69CTrmFCuWgVSELxEOhZWUeLmC+bagFSnmh0VVOYdBBr28eH4qG6cHxNmtYCbUy
KFDDZSUbawNoqOfosoBvd/WEyPPzF8RecdPK0SIUdmi8NagB/jZy/YV3B/EodFp+
dL8VW8CJIOWEjHWvWn7fNMuouz/VTAck+CLi9SWaOT5utZUNz7+i+2UsmZ/5ggXv
0opd/DcCWcBMXRccUliXk38vQIL3KUTo5KVFbBLMKGevxE2ezAixgf+9vYcdHSV3
MSXCU6kcPmDoTvvVuaLPnZTkY9viBsleqTORotW8nkyfJjdZsUoIY7qOl98fMnGv
cRni702rB6JWnqM/vZqoHSJ4q20X5yRMW6ImRpQV+usCPb5FMYm1DEzAE8I4L6Ii
bmI4VPtbNMX0bEgMwg7HWFE4XZLU6tx1sjtLq/UoC6a3QdL/bLIzvBp21WbQB8ru
/C9AXamGAHIfewu7zmy4GypCNTNhLMp6xftWfgbeY6q+CLu4g/XylR+itrud7WQ4
6KPIVLDWb90frRf9qW3T8DzUdI6lrYsWSmPCRlIo3i5phhraNa/v2ac462tE2gQg
kHn8wPOokkKUSaN4xicxHurh2U91hKxy/jldFK9ge+QogRZj2DJVnAyvEy4xBULl
NJE0UTwfeEeyMvNu8B9iWtU3poy34lLDu41yNja2J+JDOmEKu6rOc1ilh+sTbPVP
RFYU0PJPRcmoaIwGAXwpBpIZrsvT92eIrRqXxdLPtJb64rueP8VM26tb56+K20Xc
TOS1Aye3uFskZcwNX8uCgMmMpl8X9B2AC4JpTtMURk3lss8c/c2HgxHZ4CYC+7tg
6FAgi+2jAGl7QWMEcShht9OsQayIKpcInPgFB8iZ9lsdDtsQSSclNH8UPcac8pD7
qwVmKScRxEk9w+ZhvpxKxIPQVjKoVaVgMPaUPd+MRU/41a0YDRp3C25X5oH2Rxbt
EecSskxf1R0BENPTOEulr6/0VcdgwS7OoN1NTcVLN2zJU7rmboQgIxcx+kECEk5X
awtarPnw+zw7J3XuElJR1JEUPoafetDp9hsRqNjFW1G009o1egXJHAMFtpYZBOZk
Ip8WFU8KN77e5Gni4kCaGyLuDX1EX01iTw6QfgRUkM+JF7PuTKKYsE3/YbJR/2aJ
eJAcoQD9nXu49npiPjF/wzGhfvW2DV3cke3vp6OOe/rlXwYTAWjFjgsnyqPrxsyr
Bih8m3f5V0eqGvi7jdZ9okbS7KN3k3SqzqEPKxoBqGWfLw5x++DlOtAcobYhYoN2
d5mWgkG66IvvRkbF3e+pm1lX8MzjTSfV7xekQX6uFOU8bV32/GAPcjBB0LLIDD7B
F0prKgj5e7VZFWVOowGJLG9Vp/PmFx11uh+5TmcPHzQZ1I5yP0bIBzooMVg+ZKu6
/pFd1WzVBRpW810+nKEUVYI5nc8xVKwf3yPA6o5SUlLAGoCWly1DjtJImajR2Vur
mc+mmUT2T65XD3MYzDXvaWwE7qkb9YDw5zvv078L1N8XZ4qIztfHZUShoXiUqmCx
bBrQf/wl4j9eUeASTmC+bzPTsyiHBuFnum4b41xNkBcyNZIFd6fXiGiyTwr/Xn0D
VsUs7QNP/k1whPTwI76Qnfzg6J6b0NZz5y7zpn+VUdAdyVxCyGbzMWKwMMKrEVcK
+BXqbgv9mJ1yra9W4GMXVVPtKgsTvyuJxzAyZo+4CT2BVH/BRvnhhznzYuhaSEX1
TpBSQj/CvQDY1QyMBkqw9sLK38kcQBZfiZWrOVFTUoFB8kgmt9ky6ap3d+wIBccx
sNiwOEy2rEwFgZkEKDjQAlnSj6RWfXuqemiq2/9X8Rg8pISMY0XPO8govQB3emFw
si3cRWmLiHDvA/Ri8uZO59LyJXa8y44AUVg7+blddFLej77CZyQ9Hv9Fx6afBf+Q
VNiL4PWyVaavHrGYE+NgPc1Jh0qRVqpoGEnZ7otOriuJR+9UCHhj4tWnkEk7QicT
Vklo2JYnUI8q6PrDJlWSPT8wjcOWFFtTadRt6jkTAxZ4cEzr19EO3LSpzXyrJe2U
41dERwS3rPZuGxYXjLUhWOIZG78/V+aBvDLsF77RT0Bquhgni7M2CnaARA2g6Tmm
t6sq7IPcLdTtqAiUpmyq9Gma/UNlfr0esSbkr3n+faUKXZEtSj7A2GxveqY49TO5
OVGO8wqGTExCz0KgHze0c7x9bDnmISjIeGh8YgQO8lsxblkEEBsmZ8BGJog/16Dg
XadTfitqBh7ududnCpxJHcVBC7djLRAYe/la15HPriScmedBXcBdWZ6cGezMv9Lg
MgEwV3MFVQIGP0mbZ8osBq0memd4pTFVwzOKefrRfW7W42rnDIYtDFKzec3131Yc
j5TKoFU/yJdeSDhNTUM55j9KvIl/cgNWoMrV+ZUYp4Qw/ID8QeXmhXf+QhqiD55q
odNTUoTGQwGjxWNOcdQnlVNOOK10QLDAapwVCbDuD6xoRJjfacSAyBdwPFvIbip1
ncFZsPyXHSd7/8BnIbHdCLw8qsbBpWwRcrPAdX3W1mG2vRbSd4SD8zogFWPEsPsL
NH17+6o/PrB+vRkUwEEkogztLWIpid2Dy2bUCVCrWxoc9UMzQruIxe36Psg+/3xY
omNU8iArxCgssU5YURO/9oQtsL06eQLJ/dows1Xqqng+Xf05cQBz1MYVZUV4KBt/
W9wbYN7XVEe+OR2mTAZyWEozFRooXCa1eQ1tKj5i5h6kp1pbBqsTp151OglRgTjc
TCsnyOqRKLS87O/wSnb7uHlGsp3S/Kj8bYVYOsacYopC1IzcV1/iEPPNYkzk5V6d
Dp9AhT+lMQCbv02ftj87Z7p8k/7ueHXKzos+qsY9j6sWnpHEhxE8fQNILNahUXbL
xSHo8wAnjQ7oOBfSiN/UPY5o3DjHYE0yDPRCekQQ6YMoKhqm5TzNgDhRhk2ACeXT
M/3XCn209hQo0BxCJf9lX5dF2cjqRd1yewxrgQ3tITjJ0Cule8FQLUn3iegdtLKh
yVkNX0P9CfHsfngPjUKoOESDU15rotKwzgYrut289auAV2CHj1Vy8XtXyHw/icVU
WBIumvetWyTEG/owHTjLTq6q4ncHoKJBZNjikAAyInwzfREgeqs372/4hkICadZK
9MxSl4hKRoCtzV89Jp11UVJbmNGsIDCYjHkVWBizF3Ci5mSeYhclD1ItumsHYDzm
GkpyHRPs2Xvh/UruqjVqmoPG1f3Uxw9Fm0Wsurc/SO5BdNU5iHM3lE513A+hEAVk
6V42GQcFj6alS+Rji4dg/cMmBmAeKvwhGdeWwla1UE33UvfWK9dYm5b6ArM3NWEk
HceP+tl41ZE4r+HBRcY+X/Aw+NdbT3/SAbs5g1iAhuxE8jwDMKGU3CsVFg20jNFr
titFFOLRHMOeVarSCK33K6yaggkjEogoIzocgorzcy/4EE3QDhMmo3P9bYcQTxq5
Xkst8PoWA3catl8tjQ8AmT/2Xamd7ixs6Pz0oEWqz3b7O4raif2NMz6Ao12ku5JO
duWDBiE52y3vgh6bjhrDP4dAxmRwrQ17Y14ztCj5Ywk7xvkZkYZR4mnVXDEfdVp4
S7HA9HNding99XooBuQx72ttjTGkwJdAVXYs/L0mN29N+N+gdmFo3P/L8ktD56OH
SHl4Q6agKbbPnYzLWjb+F7Bk4F6H+fHhb8cX4FvpD5GvYL1BVdhQoHTDOtx7x0aW
lQ6gLh+7NiJRpnJrulF6pEC2MgdE7rooZVV6B+Pgr3MakKyPOhv/EOfniFbqdr4p
JhPWnKU8P0u1t4GtyhCQuDFnvLQyfSd37mnPniD6sFdVyg3urZtRqh2Aw+W0xyhC
0kO8v+cIOxXIrmxy/fJ2Rhl84hcfnm5COfOEqtYXHZ9W6uKfFUJCaqgn4DmARKRm
lI/34L3DD2XKbkwy79bjVt0pBNW3Q1Tdaln+sXesLBMh3RTnK2cWnLWaOET3Vdve
zoY3eyQxAXfH38JYLZuwAsdZ6diRJckGOritXKeGVSIGCZ330CcUG4M0nMGDXX9O
D/d/5EntdhppTXUq+0+Uo9A9tvU24KnJxvxfJ/5P60IN8zHek9tkQkGOnO6wxoqZ
hDEMC8UeE8irlZ2oVa7uh/UcuxCn7fZOKNzl75IsZ8Yq0tPjoZuczMeb3n/V/Y3s
vneNY1/1M1URxuaitm07c+QvFPH2SgbDc72P1OtDLgdtfDIo6WH8icQFEHWmf28/
/sHAe3cSvI5jwdx/Ahz2bYpuM8prf2FgjgvEm+RD20AzDbYqsXbSXvms5HzSzq7z
pDrrwY3i6a47f633qp5MiNnVejz4jagI20RoWh7pKCJKuZS0Ax1pteiyz7fdTvGx
zRb9lRsD9l9XGgJzHNUZb5oKHXq83sqrZ+NHxCjbF8eIpkQC4WGpaRIJev2FFcyD
Ulto7Xvbsvr9h3JaYT2Zz0YnI2uiR+jUycm7ivPN7iamykKdqFY+q97Db/fNNe/C
bkVax11tuMIVD7t089UC5AICAlLeZgp2YKiywQQ5Hiyt4mREGRAX/aMHy7qS9PWu
q99KMviFEf7BNClbljq/99PuqhT49Xv6iwdjQRJ+XH94JNLrNE/P40gnMLeJNDDV
9kgkgz39d2mN6eCwyaYglfYKTDBeUMjwsn8puMNdzwSYJbvkr+uTAJKhcuZWiSL+
otU7Gpq7G9qd0Zho8W3VZTlq6N3ZJpB94om4KQwyrHHlE4BB8tIwnJpc8cFxtueg
n//qr0/W42sglz8jlgDKKeO/rYC+UYRgnaQY6mamb3LPoTfizBzguK/tslq4NX4Y
hFi/hWl6YnJO3ErFg3bNVPHzn0dOqrzpo5/CzsGmr9RI3405yAn3zNS1Zubwx5qT
/im2Q3f0SA3IsdIJmEWryDOTbXzBEAG/hmJyjemyBifAbt9tTevNfXcRTSU4Df9H
czlzZvy72mMk4UI8A6RJkOqPYJlf/WlJfMg1MbM5aBRWDa2tiTZHixQywKY4/j9C
kdaaE8BLoXs3qpo6VYjGFMhWa9TRRmnJuH2Mnb2MpY7n4vekr16IDzy7OGgKgtaZ
jGIF6D5xQkydGddp0oIDJedtJffLfHABcR2W9RRi7T5IoHU4VGGGgDYzcTXvMVoB
EjezslNDv2wXQ+K5SYSRA+/ssfaCT7i4V2BzX3ELyi0Kz1m8RBl4SL89WXfyrS8+
A/G0d4uFALe6og7d3YQWfvaP42tX5aNVT/0aWDrlPnuffzhlEKac2usBKJdNvSjV
rfEFGOpOr7M79wpftbHYYp+ZuJUIOTOBhwiu49+Melxzdx2kw9o2HoCci9z8Tz2G
ngHHquqvTs5gt+WPOf7p8PFxcXKOgF0Ui/yHuRrB1QOdptVxOgm9ue3aBTl+G9/R
MLO2tPlbcEjGEwz437XFwFryzN7Cpok6HFr0horUBE1XYkTaYgXCaYan4hKTD1ES
kF0mpGQEHZb5LdohzN4H5BKT4yKARSLY1VGEXC3VG4tG0TTEE1hS4j7OJQ4Fw9ex
4Pw2ZLc2CV+mQzw0Ou92f1TGp+cd33KuUv9ReoyRk1Bp+SfK+bCsMbtjPQTz5Xtp
goO7U9UDQlIv29xHw4/CRgvwY35Ifcs/QiRi/d1BIKNsX7GheoZty3pLN11/tf3V
/XisLj7IpjlJRRfpGeRGNEzJVnra94v3nBkyp9L0+EL7KtbPxK25WyxT6x6fG11e
0oVPmcFDx7/COLRdAokVXOcKOl7XnaceOrX0p1TFKNB1sbQzFSo6n5H9rpY3W6UJ
tFuEwMXioVSuxSNJZOWzaQX5AMKqn3LZlXzVuOighgAp7kODh6i4QcxPdYhimWnM
F6vN3gchnOlRvKe0Ed3cnYx1UM6jxnAwlrNfh2o2wiX+O/orOTdXNAOLq7vYp7Hj
NkPXhzz6KQISNA0p1DvYzFw/F/sOk3QkaMnBLT3hfjfCHAc7ba9n9iKBIiB1e31p
Gg5T1365HdDpjj2wl13B19Lz/e9FX1ElVMCw8jcfRAHXC3buYfNWI3LeWzNzBBzJ
wmypVklBjKIPycDFG5HS+xfkz2/gbmCO/3Db/zp34cuXPTeRVStPOTvfk58frcah
5WXsTQQ1pEt/+b9Dy5mDTlm4XYC+lVNYn6rR6TJnZkVUZDD/42yNVV6Z5rCOkl9M
PkWyYgrMbkeGu3wlv+7dS93ld03CPTKEJ4RmeeCsU97JQU4rPA5gzB3y7Bxj6FW/
7bcaZw2XZcBsOmbLQPP3VFvu6D5KDqC5g3HF80vTzPjVFMgs+DDtL62SwZs5eU6b
u863eOWwfxRcKqszw79JuvsI6XUjMSxb43UACTKoDcoB54iFylGhEEcLi/MZTChg
nN6G1afxaI4ekhgp+MjrYYmOHtVUmvklbaodPwVA9cZ1XNgkMIB2pUxW8uOQn5RL
aBOn6k8HA0tlCrtRI3KFC6sj79XxtXKZ0aCDgu1y5nK2WAchfklInt6yu+7K2xI7
IUfD6a7e5PEjUZFm5ErAL4ZBXW3DhS7G5qd7ek9FEvJeMC3sICsFuJrZ30b+UJZa
JtASeOrmnu4UJ8i66rKun67Uwg1cSEYQ2jntJz3Zv6hamMcE3TSIQw64hmaJcgo/
hOMt+v94xJo2ghf0FWj4qMVrEeqRQhNG9U/7mk/SZh4HfyI4FILP00Z3r1lMe/Ka
PM5QGkIygPOvGGvAaIrEMHrVVY+cTeXy9Ftseu1ZiiTKlD/YTgvmxEjrsC33LxW6
FnOYpG/BcEhbAUs3VA31ha+q6mpZxGpGKPW89LnNT66AtTxwzISFzKBJ+VM9cyPW
y+sF6yo/N20mFx3db2jj5rYHSQfhGBS61VVL4S9xTLuCY6C+IGGZ9D5eobTCc10D
Asg7WZxqAYoe3uG5vYUQdwxF8uDxSoT81hBmX+UF6ZWEQyLxCbwQmOCe7iCHB3eH
tplAYfo+PLDl/LMpdQp2wxHyLRN6+TnEO/jC6R3CBeP8GD4DMxGhj6DNJBlzTG18
BImIMIfIlTNs4GsbiuXXWqZkFpKbWyk14UXH4KN1j02ze4YebvDqdwOodWYg10Yb
xzbapZY/0sQCKqqbXWERRn6ScKvY9YwcInBH1CizoepjwG4VcLU75X+2yxWcQCGN
mjt2pdLwV7/7BKXouAwmS+jRIMqbf7+iICeBlwbp4hs758U7fd31NfBCM/He6WwD
CsZjrPUu2U+pk5VlOrzs/EbV1KY+HKpuYHd0EKkM0jXIGIhWbUQuJ9hGdcj87r0b
1Nzu+//WgXJd8jA/ir+W0aP4uZHRoJFrYVUDpSrIoxNYQzCva6sAZAQJhja377KB
FBaCkmnxtM38QwWbYrOc0U0C0C9l1ofZW/zW2EWUuYAJ1BiRVBeBFrhVmwSP1aQi
wQVreHW1UTSQEvPrmWvdt+c/CXG1SXueTlWgPNw+O8P9W+35EEto6b2YMDA7WUr6
5BWqA3+i6w4ysHWPktvNte47OAkRTm+DYzs9SGCOQhMQeaI8TnYDgVyY7vVrEpzr
9PULpm3acbCh7bwdr8PlkSc7RZGeZ00lDPwl76Ot1al0AWy0ZbW2pooI33tFVlZ4
26e7461/1mhIhobTOuj6LnUVLPi3CviyguSVoXK9fgVonUzfEKTBpa2sFlhDJb5A
gXkKUQvxtN4V0U2QL7MEpHJExjYDttEZApuy5BicXUYv1P+zRxuCvrff4sYw+8jf
lcWV/pY2Kd6/PL10G3XnbRKRKROHYD8O1cHDB4DcYXFmMQ4OzIOxljDU8dPLmEuW
tf5O3WYaJ+KgCrJSnzdZ8CL2zxfZ98l6/pX6AszF56ry/1tiRXX4nr1Gn69Ukoet
vjcClzarw7qcYvuJiMqbkUijuvChTKC9Yj2Fa/0l4pf+5AUyhavwOmm+8tZi89l5
PSXL4kErm2q1EHOebbLmYsrDvF8gQWvxV+WwfZBE/8PypzWQpVISXO+HjVTeQmd2
lNNruE5/0W7CgpJZb3FV4rnIjRaap5d2FNAPSvLIfjUSNpgdLEetD06VbwwkryYB
dMQMTZ7cTUfcdOLhpzdKPbAhWyK3Wt3KDjLbrMPWjdWR/Zf8o/3o5HsJypiWJB8+
98WXRF4q2lR81kgw6scYTAHkAWsMpjg9MkkTkyHj1BMwfaSjHLNw9QJiqYQcBhs4
FIo992A64zi6aVK2/TlUZqK18hy2XiNs1BWurCm5aTJ76LgyBPX50Rsy538cdMnA
zmbu87FjceVxVN5V0GRcOWMrvejbj1Gamup88SqWjzDPM5n/ywwGRoCxLQGjjtWt
csSNFnJWsuAmV7D4sJpuE3jk0UB4mS5N01kOUpSg4z1ZRimApBZjcxXMca4Dq9nT
37ijRCykYoFhtPShiTPCLgMXAuf21KvSkpF6ziQWQG58eKAUjhgcyy82We/Ex1/F
d62kj9pdTYK55hkWU/mUrZ9zhYtr+5NplbmSMTP8qxzLv4AT5y7IpQ6ZBdVW80KK
tVPb2QlHPFZRrVIrvpiNp5eHu4A48XoC9v+81gNgc584cVM8CU32QcJx0hXBj6qr
CvL48US51ZgqvXAjuZsqwbT0cn2uxJKJSWfRjCLySTB9a42coxZ3fMzseaLGG6Na
iX03+lo4vTA53n4gYVOjBVGvVbccNjRfpvb2Qon4JEMA4HxD8ITBFo41bgea5IM7
4cWjlyagevOhgI/peKZFWsKTMhQ/SUUE57Looh3XUqWvRpQwlKXYYQTsoAKnfvoa
4C/NOIwtrz9Hi4l6G14dD3MuLcPcpGUhI+GqDF6ag1SK4VfXUOCxLMHAU8Mdq7Kl
D6wrjRXHVgACduYG4I49hnin00e+zY0BtwJQXv/m5ODurej9jcNgFOg4BK7ZbmzQ
qdPMUdk1aOuRux6O1rQ0G6cxBrPqgdBq4WvARB8NWHF5ljbK290tz5UR9cJ1hvwL
Vwsd0WoPxCUdgkWijFLKEnsy1VJjiVsFETxgOpwWekOJHBEbR1Qnt/YwAeTk9OJt
GqujpiIT6dvAz9B5SJV1+xr4O+TiwaZiMFBgRDdg1lwPOBNicIGodmzHj0hyLO6B
seXR004Ulru+KC+TOd1bTxtDCZV6fOG4ejcW2iDmR/xuMdKou6Qma0jJKHPIREtS
YkyCdjZ9NkwFQYX+F/bHw2xzrn8XuRSzt2pHP+tzJH8/ItZAquwcbrnK9GEugiUt
1cq6MKOOqllWJRxxfDmI3bo6oFN/BcnV9wGqLM7jBINpuLstnVL3at/n32pI6NQD
T3QkEK0UTLCveg0J/lYJMrHay85l2oXAsT3e15Xa1I8dMNceOnTGN4bxRjxIqXl2
SAdi/fA7HxEAIxmeyz8DfltS/nfEftHdeCOvQl8Sa0ukJpwpCMBskkZlhIxPrOO7
teMUlXe+3e/w1ehyx52lbOvrXR6E2W9l7l/Vx1hdXGcqqcXLj7l8oJXq0X46cf+X
aJwGsrBbOY+WvjXXwru1xsfmqc4ydSny++kdrXpCFonvKs/8EF7XUDVOAo7KIFQd
mkLcvqAX+In+hBMyWVdI1PU6qCty2G63CpZt4XUgVeAydrfw5gS54awWxOIaNUds
MibHaSwJPOHQGuTTs7h+rBpDNSBBLiWnW2u9jGO7Z7iVScB6ucwVtqgeVJauFY/h
tstX6QliMC4CdmpmY77ue9mJGgtYG/gqEcyDcmgpoWWOcS+ppm/lLTH5povr8qcw
+QtFtpELcP2+lJwk+b75JaCmwDTXX9KUwo6F7GoAgSmqh5pTuDm+j2LvE0pyhqag
8LMIUOi9l7yMB/kZHBs0A+Y/RzS3NvrXtJILo8rCDxtJizyctZpR2fxPaFO0pxRy
s/e2B8xiNp5Hzp/hqmnBKP68RVoI/iy+MMqdGRi3H+HwVXx2wPrx7iyKwyDiauKJ
dawaAvAnbj1hoi+NBYfvdNGI15LeBGtltXwqxN4u5YqUspA7Iiok5fAm658ja58u
5LFbIfEqsBx055uct1CVrc23y6vUHqG0zFeEQrLbTrKrst5djoAu5/kaXgzlHHsf
F3N8n3leoQLoAVHW2ZnlUA3FDsBqQqZhtaqVK42EhEfPp1pjgpnLVWLu9z24pgrq
kCzeo+yrLqMoBn4Bk13jbPOmtp4CtwI0iJOTSNI6nNhObW9fWC6/TcaCAzwO99df
jMEuZ++P8puXvF5psBRlPv7zvadoCm4Vjn7Kg8dX2gOAR7bxEjBLPPn06FLpLb74
qRINuJUeAd3xNGUeu2DwjvDnsy5WeT/5lO3FLeDANKtYS9CW/OOYjktuthYS8skP
EAoAin1ZqySmMfr3OKD6DNLnkogE+iX+hekqvTdB90SUxnI8imzmaZIo3471zhFP
Nxp+hHydPleBEFyN3bIuEcoVngrEH6bG6/9gsV/WERkeitfmE9Fwmpdd4FBWzkqj
UB+fKmccTxaJme2lsxqpX79sdkuRdaDidm0/PV2xFiveqik1QmrLv5gViC+ZaSwt
XnlDDzU/VJ92aaeQQO8CdxDGXmzYpRHMib4q4ZY7lOFnbTib7Co2TFJg7IOsRMXV
rJBoej9068p13mfBGI4jVmgai67t5KizjW+2SUtX2RCJA4XRR6dbJtUTJGzj068S
ErWQIHmgWEBltZPGJ/dWwNwfk1XRCcjH1RiqE3OQz5IxFuNu/xSN0PHZuuteKSM0
Txc5H2WSzxx2v93GzkuhBKUOKqrZc1nRsticRjyGP7W62TnSVaggzexNGFJqPYIl
DuYFV9/rWkxBJzSa9N8C25jVGMlRk0jda1mnrq0MUqSb7oifPdBZFRyvdGyQLWGn
XK8SY39mCcWLxH3EDVsvXFlMJ4xrAg1Ky2FpM0pafre8f58cXdPfXILXfo7fZ32H
CRtfN54acOTyKf3tii8/IaS3bjFRnyDlZnRq2Ef7UaWiDY+Gz4Qkn1bGJKQP7l//
D3mRyplCDJi8fCPNFikOZl9FbbnR5V4E/LNcvTav3aW/2I2L9onqIQuWrKUcWiIb
2LZCROZVGpXeu+xCHsXTN127TUB/mXaaG5E6rHu+bdOsebhkwmXOrUCZxiCwNm74
QMehzi1pgBSZkCpau3Efd7yMx1OAtppANfz/wysueLcWw9SPij/XeV7fvAdWVnv8
2oB4Dwq3xrwJFf2Syf7vhJ+PGtgW6m23TKtVw/kItS0kl3kEqDg2ZXJU4o0HY3hi
ZY2nv1TnmnZEvA1rR5/mnIbEBJ7h8XHWxKqRPukTWnpXv9iHXqDsJrW9+qo9LrwT
gtAUhy3ICZKZXBIXsMBUA7hDLlCP98xUMF4QjVoAZBMm3J4VeMxx7QCn3lD+9D63
5lwCHar5XowhpA5jK2gYXdsr0g4L2+pL8CdrSeQ+0foNxv8FBkH0Mmh6q3R0ZbjG
jxhKMWy7LK4fZxJ2XIxvIDTqDLZi8eWjGh/TAZpsemTzz/FMUtaxpSAJ4WzY0+B1
BMTxTFAjdKPm4wXn1KHmCfSiOw1WZU6+s2Lc4rJtcOqO8LQXbmrcfRac9O19LGm+
9tdO9IGTwq+mwQ3G/rtCrsEP3rHMiyxp6jaKW2I4Kb2c30CCSjY7INf+6/V+vxNd
0xIBUpcv2PnjxvuN5H7XXeUkEAW86BOySnkXsV6+dil8S/vKRC074fuM9g6w6JsP
ZowX8rI+tGA+h8sl8b/k/GngB9D8tTGHcq7YMs8BUblNeF0ZkOumplgq85ySfd2V
lGbxZfcWL8ydBGf9bMJvkOzcB8V+xgVjnWBHVO5lpq11YNyvthCooM7G0cCrf1Pn
vg+uekfJv7OYLm98Xzi3y+1ZJsno7Akj3mR7keDzrXJZoBKYDeuWLTGnK6DqDGOS
Zx/Z2d4Q4+eUwgQ+PFU/eCsRM6SmB3DHoyqX3v8v4UwRwQ4u7SdD+jh9Vssa3cpZ
EmS8RWgY0qvU2c3TLZO2VDG1RbQ95TUYTz5OUT0DLour3b4xWYnrjV5Rh5Hd0rj3
+cBBGBuZjQ10oEE/RvLM7ZOkLFtsdmjCpCqu1jDG2Ty5SkBEIphApfb1MSemoF05
OKuR9NTjTOSrR7qKui0d164OZkbk71JYOr4dDaDQsdEOsNYOO71e3caZIEa3Gwj7
rjq7ysdbVFcqVzOY5r2w50LbzwWLZRX4fuENM9xSt2gdQZGLptEcpN6fFr4qkVY8
RSGJkRMzChwtnF1zbbDvF/Ipx6zCRFU1oqhzROT3VSnKbndcDowRRF6+RrLt3rJd
tQ3PkBq+zB9Y4zbrkoiOHrGik3u59p1ndObh+gOsbIiHhSqQ7A9xyB0NJWeQh34W
oreVVFWpjIGfvOSFhvy0V2j8UTD0NshqM5FDsjhS0OMKrldmtBuXawnPxD8bS72b
TguKiF6gug2p2sI78XTJcup+axi/4MuiYUng3yBcEKxintKExd5L7wAMY6fOVflZ
G16peEIvLcLd5lbXOULQSBDq3UrdPLo9cOS/fkhZ/N1uIyN7LYWSY9aLFU34VIMq
2LpxVe4xQ21UwqccXP8tS6cXpSgNmY8kCv7lNvQeadCik10g4GxPcxmARXtkQ/Cs
0MlAZNWJde+1lBe9NVQIybPAR2VZV2bdJKgL4dLefGsDiZIZVejeUsJJtGkGEx2e
U9d3dRstmEfkOH9lqogfWP3Q1oNmjrMTdP58pDNQ6j6k9pQ/0boqWxaQk9P9Ghgi
FqeBazpb7CFHl4CilxuDEmUKKgdcGjoyO6idLbkrZJfZQkQfiMUjwOE2qEbvcb2H
/R+lNT/f0PkjXWoeoBUyvZXMyW6/eEa6/7l6iul9wJoe5o9XvR58jE+0IHZdXQbL
AD4obZkdO7p0f3avGAKb5ZKFZdbczHAzdXQX/+PDxztkX8zKr4zA4O+pH3pmec9C
pd55F554fDRaGPdmBxqhrad51MyQsQ8nwmVSILwVzQSZCuDFMwfVPWUiTX9lpFFK
Bk4uqZNSlYu8TY3ZN5LkxCkdwoHXwC4aw7V6+8WDXE22Gy061MDd0xBN0XSqyPIg
bcLSeOtAu00Rq8MhQaR67GuxRr8vtRYpR67PHwxRUZbs1x/eOxw4OUdV/2sE5hlk
/q25aHDTBP4S+DexsW5iQVu3z71yw8vILMeTA0UiUlJcLel199r8XqBXRB8dg8r7
97cyOeWNK55iO7xrppPMtNfvdWQQqarV7RwihDwIn9HqdhMLRazegR7WhjQ4UH62
x13W+BvNBBUy/cE3yZRea1M24BZe0cLxvCq0LaOVyYAxo+WW9n+aj306qFnlZhzy
WXCyIO3f4O+t9PbKZB6DCtKLnDvhhRCL6HHkQXXoS5lcdRLYR+JOP+mGl6BhmSyh
jx18qi9zKWxbXWV/UVJD7V1npiYSmbUM2Q/hkjhJr4n0S3XfsoJsfp+HX8jtDtIW
ETrYKW9JmjjB+PWqqOfLwEy1vKeGa3Vm2WWgzyRRSjJ7BpBFggH3ArwcGL9Gu6ow
X2IXdebphnaGE1scx1hafof2HUjtc10Nr3l+lL/QIBjFiAH134kh9Hw+XXlk8TrZ
vEMUW1b4zBAYvDYBanKnOxz2i6xi+dMs7NCHN7o91oTP3LDNc7AfuPTbHiMPcvPe
XIYCc8hwzXJ026IC6tbBprR8FwF/EXr7SvAYdsTnNHm6cM1LJ2DJPugmtDMiyKbh
nghV2cRK3ZBwbpm/yd+mogM2Xf8a6JdP3v21cIgM9qD/dgrSnfcVZDxbsnYNU3Wd
wX6ClQ6sL8P1XW4uGd3OAd24hGMn24sPJ+POa1twDzQfdLZiRTPh3lUFFWJALX61
MwTyLDHEs/BaRH2mh02QbGT8CpP7e0e28FOZDJYyQaFweLFrRWdFO8DINxAmRJt7
dZZmvIUYYefk8BFgSRw0N1MSNESLXbz03TLuNtreJTCL/I39uXRpNBnEK3DBgmSA
dMNt04aEILPn2YdQOpKfc35OozQqGqqo4ZeNTCHffDVpqrVbWcts0a+L2dKB+7m/
wHp4bp9krEoXvOPBMt3mrPBlhq6C7jsV6H2KGR1bqyyWNj+1wMOTrwat4SoLqb0P
gvRzgHyK/N3amCH22ppzuvAqrat9QxPR/ODVOzgHE1f64K8b3Y9rjoBiT1Vvg2+w
eL1MAg808DfQaJtI8nNvvufn5wxJx4jrDuTZyo0Okb6o1G9/pUplnqaTwsc0fFH2
ZH/7rWzu4wy/tYR0MjE6VJee4ZtXJvboUgaTdEG9k+1tp5+O2+27vZBZw/itqMPm
d0M2AiUsIzPOdLB9uZgj+rxal14QKs1CA35uy/kscek7mIqtS1Jz0IHatzqU2Vr9
0DJq/rgRX0YpsYr38fB0LK3k1LDn1HoyliZIdboWxvDsPQ1e8FwryKcTNo0ACADI
aJqowrsDPt5d84XOIQ9b2JnzpxaUowez3Jki2zn11QhYTyn8rP2Gg083Oxh5HMEg
bM5+Dh5DIKjAhEeAZh113xBTQOdrPcM+K87iB1/nnbK3sCJp9Ag/SNUJ1xVBOuT6
CAh4gftuTFRlY0TsiudQhh4Mr22gggTyNIbYvNQseIX7ACExPswVBfqaFb5QrnHX
6/u7IogO/9DmdUZucA/c1aR4+usMgfvHb4ykfn6gJMPxOmNLMssJ56cJXU/WnPfE
7V918y/b7d60MpBo+2kyLf95xTfvANBRGED7RkyJV7JCu5PL2CHUQ2c/sU+D7P2R
Nq1zsAfJk/S86lT4zcfTeJLlS4Dz1FKVJ5+qTpu5ZqCBwx4v2VZ/oYoSnuvibZZ3
/QgVvXz9kJ15tKznu3LGxhYWtFE14psnai/MHojpzGcqH3PCjnH2JZ/TVgbgtEWM
nFopYCiDMAr3h7MSopVaUQbZwV12JibpkaaJECU2SopPw4YpKnDYMVyGrwMQYtYU
gB9aAPa2k2nLWhZ1cpuUjonb26H57o8cYn5CTqxiROxeXBmdCdA4Fy9yjysFnBaN
2jJABKg0ZXAAb9+bn9i4CFAg4Q8xaEtG01r7ZJPxYJjFxWnexOE33P6i6wc2Gn0I
6KmzBZIyOYsIeiqLHDL3CV+bpDqpa0dqjT136YAJv8JE1yh1OVSt35YsgRtNa2Fv
jIbD0vFsjL5cKM5WC0hWPtIJGEzjt3WLeKALfaC/FmvUtorO+jrvB8Rly/XxpV1S
98AF63IVNmEWbOBpHZaXfD2hN47BrmDrW1Oh23aKCM8BTC+hzTp9QZd+PBsr+zJX
tOkxurov1jbgYIrCtoi/tuv9p53Zxf4BJHVKr3kx/JpHmBtyc7MX3zbI4vOpLIhO
V7Zm7bKp/J5LK0qNsmTwC4O8mVtikeaKZn0bZ4hmjFxsdpSQXA/2GmjXQQQoyLu1
GMcUt6/eCQF8AEklsQsjReEM6Y1PtskabYJAoS8piZ6rhPfn1VyOeGEHASb8g/gZ
EP+oLBe7BiHlSBrSs/24kLtgrXg9FmIZJHcUTTMA0gHIj67MrB5OWmyO985MBcM8
8xAg96Onl58UADHhHtXglilfYwrtvTzDL9cblSCO7zCR6BWGctrKE5w9VcR6UBa2
ABIXsXRB3B28N1/DP7s1Ldojo4l199kaeD4ZqJUhHk4YEtf9srO7dAaHTiaom+vx
SWa6kC0U7Y7ZVsGxAq3a0qIJKII5/Q4xu20EEP6ROyw6iJpfZRNaH2xe+7d1cxao
Q8qoVJfbu1J5fwpADD2CcZm2zaadC+azH4uUr51SfqwQeqx1KRtWwc/iAPzyji9t
bmRxKZvVA6tiRbuPTrqgtoybWpL4jJKAIyt2zvvJSNIRV7CB/w//jwOKK0xRrIF+
RR2qgFAZqjx5aIB/pIp3TIY6jmMA0PatNRw5gTtCEn1iKRxH7hSZpeNANzFHKQIS
RXdvHGUCKBfFMDVZ4TZpT8K8NuCeER+q8erhbPt/bFkzDG5FouiYjvXsIM+OvVEJ
W8A3XHhWftXdulkDfwfsPYvr019uDIVYYNJef8x4EMvjGp0I9ypiye5T2bBDZ3Ov
T1cQ9L9laBk9uIzHLRl6YMw0TT/yrHq58cFvZmSVHFO4Jp0J3yxa209qCHZVxe3e
AT1PQmvZbReNXJ29u+ftcZ+hTBY/tJcJdyNld8V0HVwDbTg/5E5DHSf/n0egZ0MI
pYpowhuz8t2Cz2CvVCx8Oq8OkP7GPAmsDLw9AbNfCyijJz0dhoSTmLL5U/SGZiz3
MQna2AF33cwKqEKT+PDNRHq8c0Q2ZFThK48x8N65FdPdL9TqaKlDarLrwHyjm7ZN
uzARt2GYxsNHZ/YZzMyFUfSM5mKIWxTfZEfTH4JUSV8oC+leq6Wko6RunisTHsAj
TP3TKUwGRlMaeN80Lfgw6Zr1NSASDmy0HI1hkfkiAYf5Kow3DQWRi+89klFcf/rA
znAYaUYx7Fs1DVsukJHH6t/ECVimx/S3YYi66qS7RZptCWqRbMcShKkEOT7QggFH
HykJ55PWqmfrLGxRESirwFMG6HVNYq/4fazpO1fJogXo8oU87mAisHREM/BlPIJN
lvPi+Ek3Il69AjgGbh3zKn7Pn098ovcHpCsNwEvNW9rwP370nlL4UJf0rPRT6dXK
MAisgR0yd2eaY5L89k3hqIIvG6stqquwMmb7FSOcwehNcYsSgf9WbFs07cQ5303I
EiWkaCM+e3+i90lvpHFGnlyTFLrdBXkPSBgrJ2t0QtdUWOAb0E7djT/BjNCnWbVU
ktRFWojj2QLILXPrbkEJshnET4WfDDxGTCcCX9QSU/3KzHvfI6FHiid3ObjArRrH
IpFevWdDbKznjR555+K1kNLNfGm9L+dN/+mdlHp4sA8xBvg6U3Ey4PLZ4o/WeNQE
V3SFtOYqWGeJu24dp6UnLfSJAFBz8k2WX9+F52bVXHom919F6iVQGMrDRJNAVprR
3rZKginB7RRc1NFtZdcV99gz36Vil+XQet7oOJyoQmKNHMh0DFi7Pbk1RiplQu5Q
0LBwB4CCMv4qnYVT40iC51FzDgP/l2VVZybgTb5ve+NR3xN7vTuA+9nn3Yb+ZxRp
9Wcd5mM/R9PFzxuBSzw10u3MvjiONKRalD2AmHjsEBS/3skjHQMDxnnkhmHnGsrv
rDW5w7XJuNljkMiz89QYo9IFt+3M7Bpcj2EC69yyK3KML4++HLQKvtjxz6ire9sd
DOMMruVpccSygVCeuP3punoy7lJInJY//qAK5lR279CM2B+ZMN99fx6T5ItV3S1D
V7+EZTpEyx6GgfGUpeav/rXSRrIa621r1Ng+Iz3i+huX09s/B7toY8usVRACe2tn
2k1Fj4CJG+mHPtEVKmNvEOXEqOVHvlnb/LMSQpAufKXcxoVKj6cX6vBJoYZIZwd7
yZYZ2J7mkFCLHpTfrGXenrHo7sb96XTakfhTlpVJqwivBAISYL0VH+2TxibVZc2J
OxKwsI6g/gHoOwSOczCaOi/Qxp4DAo8CXLWCLug4Hfqf9cpbPdGnTl3b91UoOTRL
g4N5Y7mkyHABu2nINeSYRjhAx9DoTKPbbvgXLc8lHPpy3A+ncAro5CiTe0m/noxP
lU5zzMgKjY2renCKVvB/TRdSlAI1xxZqTgErCJipK6BDqs715bU9WteAmf6m5Rxi
Ze2soPaeIL2pHNRDX107Ha5Ts8EGJAzBpS8K8bXe4G7W91GkaUO3tP44FdusUfT1
2sWdzLEr4JPl/4ELkT2s/sUJVVRRgeMu8QEU0/4ni62858YJIvliTkrvG5EKxrDX
hB7mAYAikitxU4eEjOFiisr+3KqzktyzJ5VCD6gC2tlFxNUJ4iOwBZvOAABzYT22
heEoBHmpgAlM0Yk+ZLC2KEBIaqBqbpPeAuWoy7rmMlGkZC6sNpPg7ryMILH+TYuW
1Wg5Y1UAX9unsq28GRwithnpn0xs9IP7I9ZvpYcP5rmYcqqsF3VKUk3M+jPWMaLv
YvalJRDKWMNqjHwldroRbh94UJBDQi9ybOPsDpZuLO86BuB5TOcvPZ+9EVjM0QWZ
EQ1yOY7dwmuhJ5WX08NMtMfg4gyKMKwiVzWu+J5l/2TUdItF1vzuzn91c+iKz7PF
ixW20N7Tca/oj64LO4KWwv/XO/bM1Tpoj/JLMK2Bkf3X280EV7x+6mMd6jh69nUp
3Vt/mQUHiFg+si9XeQ2Xm99i5IWMDWH2GYpOaNcfFXOkeD3xca4GUlX+DmvXlWFU
8jpxvm/L3RGsBhQIziofEIskFWhrpBQQPI15tZf5pjgRrSOq75+59X6r3zABG1ug
pGkWEb8uR1hKCLe8VLy1WpcxthBF+F2rc3XVleYsux6wcJvRSTktz3osZj1L6BGk
6nLN+5f9IaUIKS0gq0v/XBpkmtnH+anxPMKYOQn8MXmdGVXxTQE9RCcB0sc+tjO+
/Vh7zg17EO00U84jGoMcnnR/GGtzs+gWHDss+BhZHJDMWgYE8AMeroU0dpR+3hMk
OyCbrW8FWu/I/sEKzV0FtGPJ+Yn13WJ2FM1slOgqzfIkU+Ng2dtPz5H5h7SSxAbs
TxTXb5QRVK5xCEvlzeHpsw6HI/pnqmj7nyPraDGqzXo0InrF5TyOU9pyl6u/Q8Br
5wVlyoelHn/hmT0jiAS/ARUbwBMuwyFYdRGZ6SKnVN67Ax/njyc2ddTeRUIR5X2W
y45Z+dQ4rGgqESgJGeFDFkucgQqJ3hnMbhqBG/Cf+nXpT9YQJR7Qdn3282lmtzQL
2c5wAGY73eSyJpU9eB5SOcaKqVAlKhIRGgOGTEfuiItgw8s/o3SSXRW4FDx4ULvw
PabWKN5KUaqkSzFSR6M8/Oxg39hCrkCBHxYIlpBD9nu3xkgxrsQsm1cmAoYkUVXJ
K7liztkrzmW/zkPsdutzRtDCRRbBBjDQFQSCgx+0ELkZc2JnUNkXqEj9BTVONPaG
tGJ3CXUnLCWTSTj2XEaTD8FaP/n8sichTenUhKA5vtciL8As/xeejdyk0xq+e9gL
S8/nSs2vzaPbFRqmTayJ0TFTK8RHR3RgSgkooYrBS8L9Rc6teLiN2kgfCD40tfkT
e2jMzEgtKXotbBnWZzsKJO5ED9r8K1lT5x0epofpjNmcv9vX3g2moBXoRK8vLBFX
LTAQ824EYhr7ZbXxS4Qv6RY/RFv0cZkzbjc2fz6EBtlxktph2eq1EPyN2gwWuG+F
zeBUYDhOq3s3NwKPS8b5QKk2wir3afF0sbKbkQVDZeDp35DKV/qNQ2sx3dAN+WH3
lxQSzY19H4AePvTBve5+LHKlW/8aySPy21lx1DWKYhOmLXy6GfwEoHA6f96Yb+83
UyMcYfTH9lVf5Aqc9vLAsrHgn8ZC4tXV/Ny3nRpcHyLtV6kkY4bVucfmHv48OOax
Je/7VjSyr7C/k0vRMsolturzudFHfPTfbh/q79uMblha1vfT5rYFvOQv/ItW3nvt
Nb7tilx3TlgsYfxQo5vzuvERyMFQrN2M+X8MNoMCUBWQ7J2laJOz65Zc1qe8P8YL
uL2zkzE3oGESQmqN9Qse6syp7CoBfCA3T6rYWXxPvqFWxdyXPduGFSynnPrZ3g64
R3WmrXgRepd5o0jJ1vmIuuqyANzYOF/MS78dcPfx5F8jd8eKkdRXDRdyrDfV2UfT
9DhOQ1Dwn+Ihf5rYorSEIiZ5SY0G6WQlWNKiH0FLxph/tymvUX7wtXf8a5a9O93Y
difGQg+ZG9Y4sC87SSta41l2cozcayiY2kChghlxpDQfdQjjTxeOpZfB2ZRSlcm5
1Tle63r4LTgAofbO7qld1ysto3w+guygkJeJV8m/8YCQ1FKZPyyyKO0C6W8CCy+r
6FqpFQEIVGI7ADYZ6m/C8kCooytkS3yUMuGHkK20p5w2Wx48hrG9xESX0VhHKPy4
gbx5ed07GTIKZaaNw9M9OU1mU50YVUX0RXGIo4QZ2XSE4qVZo5mWm19LqugkerVH
9siA/NyGMM0cqRXAJPMtMdvp6tmlUg4txT4w4My2fW+DBornYxX9ssjcbEaQH1/m
jWwsozEqBehNniEo4/wf0vQcbeJu/D+aQapmOZxfab2VL5vdDGavqFGKhfnPHG2J
czC/z1yRqCskMIos8PdhMgkWRKdfg2DaghKmytGQyW5ZZia/JWadCkZxw1jKnqup
OiqL3Yw7+u5En10GKelKRs3I0QzekOMmohDILRpaYlYBjjoHeaM/V4zCvFrGYcud
ClABIuWyOmwwykNz07dxRfVh9CZJJZ7cY2XdUkZiP3XNqggAMhwa2t3SCvvLkggS
TvBQwi1IxiwKCc0ceeTB3xqJAq9rM1n7VpDGVBtgH1doC7iDceQQvfmsTHmt8pAd
25xhQUtEj6QIhVW59xfafon+iV3KfL1jyoFJ8B8utWDWSTi6G4cKQvCmubeWYPP/
pF/kyD0U3EHdekuYKYT8xd39Wb8ag5L+vUx6x/oeut5fAi+FYTc2NS8hf3O8r2Sc
7fECVAIvyucfmmCQwZTSxmr4S67GK9x0ie7JlHxyf4fvuEytBnRfJegtAhGgwR3K
KWdXrSO0HaoGV924+/Wb9QdE0KqM2AOsyqG8VQcXgeg7VOz28Cj32PmF0OaQTZvl
6QNyeKhHRu1wX6y1p8znvi22cdsk51WheJT8QETRwJamVUSwAoaDslwpDMhe57h7
mhj887f0/roxANlJ0iUjC98XA8C5Kmu5QQRFf1ryOC+5zrQfJYyZ6vJ2oyHkO4Yb
cUEEtpjMzznKNX1F9lOJZ0EYa62IUM+BWJ6Oaf8wG7mllgALkC5trS6nLKQObsFk
quG9V/4igC4g2PJjI0gtfzJxnbw0jjKGZlstb2prPLbuBww/RF4/Agg6RMChcs2I
hXztKiZqDAmi/2NGP9ZOK1MwLp/88neAeG5PBBk1Mwmuuycq8KOAOJK6b/BRijfN
MAJjTGxVM/JdlknwyYlYv+Y9bh8MUgVlXJEfdMnkYgtmFmfaN7gmEvMnX0FgBVzw
x+srmEbqKRd06rNvJifrR1vQucjLSvUsVLVDs3SIr5/himXuCxdXUJMAQZcCLhJA
XPfuwk7rRCxkTJLxgzOHFktjc42PVcM1DAalPjJjUhs2tFZAynfCfHsF5vriicK1
Ev4hhD7A2c9gD+TRD5GA2ET8FBvp6SsA5xySNdaolpIF5qd9I3DMgYQ+xw7qfcG5
cI6RemVq9ilvAwNMrfTLwB1PdZP1rOYZC56yvl5VSuS47PYea8tt+UYfg5aiFpn4
B1m6OzupdJvfXBo4n/HlHzgqkvmTpoyUSuJRAg4Ns+xBHgfDiN8ST6Bz1+HXlpCb
QLb9mep8+sYuSrSZWtJQU/eK9DFajY/2FAK02TIR2q57vwR+S61bo9Iusqo5MPnA
SosuRnBzcdmUJ/JtgrsD0DtP+I48aJegq6JCv2tiQqdW6wXytLbX9OpKghqiGFGm
wfeFaYuMnN7VqJkE7Ojj6/jXHDDIpfeMrZMNIyXwWKuetsaDXOKLPGc/EeQjyNsr
xQorXJQfrNgstJ8FzPysLEv/nbeM9SEAerGnDtgA0v4HqWadQAjVphRUrzkTKLmf
og190P6Q1KbEomXXStXiu68k4xh8dq7KSnbnyxlF7Zy7D61HLQk1hT0jRez1ViF0
gWcuSFzfWigBPvGUEE02Av0V9gz3kL7eD/Iu713mRwaYn/ZWvzD/8v1Ph9iH3bXA
v2c6CU31wRpfz92BmvNKwf7vWB/nehn2EnNY05TtYzY1/WMWKaiVJjnLmAxv//JB
1VHqjQY62X6R7oRRVVLusqc7qG1Tr6JyKmM+uK+slfXfA7dx0y/TfQxUBgF6yGKM
hPDameFQevN0arTavc7aSQoSjIlIDaabG8g6MApGxfhOaLIy9TdRw3O9STbqvGAL
/ASq46x1XmtHb2niI+9SUOXUYG2VlVq2xtoyMVwVnvtiYuEX5+Jrl7sYBTiEEXuN
vgwBghr5HrhxnUQ2LIEXLxF1GGAhLWTJO4cF+qs8gwa0WMDYNawH8PJM8jUFQCN1
PInV81Xl7bFaPYvpfLv3F7YO20o9BdgiAXBiqTBI8GBgeBahl4sOn0esiWiX7u3g
RKyAUX6N5ZNriOvjWH3g9Qt1xB8BI8Z34NFNEn1sJfMhBEIftZgvFOGbc3ra0p5b
Pmo62uJoWCCrdybUsN/Q+Jkonf7AcJniiAIDryPsHc49zQI+pJ02DQJIFXAnck0F
A0aZopg8cabIX1Re3JoBdkPJOr/E8Wdyt++Uqs1JR8veDC3MGs7J/0Hw7timyZ7C
raWpqqx+GvaJMp1Ej0GtQYya/9tsiaBo7pUtvBmyCw16loM+uUTK7OeTQ0N5oX1f
GFIVcpI8LdVBqn86ta5xsc3HIBHid5spj09RTILf59aednD8s84ZIyrWrbNmGbeH
GdvLHXsb8qnd5PTBOwD+MTv8p9r4B0gFpDWSFC7Ot9yM2iYJjXW3IoW8ONvUiKHc
zsgIQdJWvtEO7cDz+5A5J2R1MWxQxk6ky3wagzwgNd1amus52k1sIHzfcVmrh7xH
9Hsi2s3X2aoDEhzOfSHAt1rZkISknWvBciNmb/5aoQ/ENCwAc3xggqJa3w/PPKbp
umHNZ0j8VA84h62om7E4j6Y4v7n7LlMivb1UrZ0YtqirA96wUDZwgHneTCQsQbAE
+Ha30JYke7csaNMXhjH/Sk8ccrotzkg0xzdv9/VKLptDe6gIdj0OWLJeF3Qj1F6F
hc/jAXZuXYF2MQaUS9+bIGFJi6MM7DxGw+RAKo8ra9A47NR/JzFOSM2DldQDyIXA
xrghlfktNkt0neUzEyfoV5nAuzKakqiIjylx+8XsQ9Ydm4sMlF8/3FAlIUzXKCUd
ztqsfV0SThUxEs6Du8+yejP59eoh6vRkJk5qkOo0eksGnylLOjHKocgeDsWflhlh
TLtCR8De2n/ZNZ5egrbmtpyIgmVYxxJVxp098ErC1c8KBhJM+EXPUDj8eyLKuFuz
iClADsOo2hKfccQxl0cUPv/R+stfPCuvd1YXSi5gUjJRkMiWarOmrLj8Yyx9aEww
oP1QDOS+QZ8aE1W9VOm0nN78YXWRVfh3pKVI53zG4nJ6rzwQRyRs06p5cZ+kex+F
fu3WBqiptTuMd+777xImuhjZbAYmXeTUPlTiuSgCBLbj3H1svotfkeq7nuaV4rA2
jWysaVt2BpYdx3ITSZoKXoyqbVfT59a/W0lu+wMsEk4jsG73+A9Lr2yulp8DS10D
q6BniDiEBBT1qszh+HMDgT7nMyE3fD7286a+FyLieAJlTTuk92EwzaPBI4elhgDq
nu7c3WBxQdEmgIg5A9mLaEtMqhccaZSEVEffOpP+H2FNswlS+xD9qbWOvYgYit7T
kRzPnmbleSm7TXg8c2qv9PqnC9TGavJNcxu6LJylxvZH03gldw7Q072+I/EnN4Oj
gbQksXA0/4pJlrTnbsh096LezpPk1NGgz2UereCCmOCtxnXcRB6b4Fg+TKdIeZL5
PVN6v6cCJKqUzjlEt7JE3enHJyAupOFdVwS719e5buBssJL8RLkSafyOmAbyDcL3
1oAezJrXvE20bld/QoO9oGQtPid88kcr76omrzdBVBahM7wzchsl1ZEE6HmSfmK1
O0lwaJ5K1Ku5BBRo7H0iY2S/QFJWOdn6GJ2CEC40O6ayI55l7smlhP57Zl5HT2A8
sVDJDCiCG+PmNa6wieLzeRDZQ4IkXsfnbaBMAtaEyCnyDT2w1QxikH1Mm4OAlMU/
4iH79ZMN4E5mzJ8kZZECbzseaAkTr68h2jbGV/hYY4PYnLczE8MAiRgWs3UpBrrI
IZSaQDp4po4saqss44kkRBL81HJvo/M2hki0ZO0amWneFe4LA6cFhjppbRauqao/
3Ocoblr2ka+n/VI/34Qdn1iWQ7N+sRO+cAcJ11TmaQc9Bf+k3rDmSgw+rvc+xHZk
Mu/3gN8J5vxY0i73+Tkz+X4kK5QAf/gsYrsCXxYMH0qKHCy82wc9taBJ8Oz86LB7
xkLg+i5Va6jxp4/2Ybogy3nu46+0iXhS9P3z7bQvcwAZdhWkKXT4tqF+PA6K63eX
x6x7EW/IehD825f4IBhlKwsTvWSUjRqtuf7dKmUKU+2g1dntF+5/IYN5ipkXPl5e
xp6/BS2YJUm6z5/znTNYKAi42TOHiRpvoymuwf1usLCRoNzuOun3yZ3WmqZZKBCh
HyviVVhXZZOxLSX5YAUgil9UuDIdnxhITf/725hLguC/Guu//JK6YqEpA3OnWckG
A3xEGErcQqtfjhvSKf2PfVPr7d+P6Jw2/QarolRGTR2/mpVrjSPUIZ7gc6mNqkNr
TTJ8dsRzvpYgZ4Mf+ZUZsHH34v9wMxIiYZBdtS6fnXMDqvCh/Vo5zaPEjjPCJsz3
YLpGeZ+uquH8EIhacU4tiir5NC596PMe7vnE2PgifpmTGurG7eU/Gd2WGt98GDKs
INGEtdhGlNecyxAnuS5rphlDANJ1WhI/+ysakzwE53gzEw1o0uxNz6XmZj76JCKT
S3mtB7Euy/gBczpEvq6gbq7xjkyABUYW76X3/Q+0kxHfwSUE8cUGlBNkpbtAuKGd
od4WtJheDeMp/Di0hfn24VlzdgbQQBBOlwgEAug6e4eIenKR4s60RRsUarW+C+xL
siDAUJzZGm0ErhSGdgWKk49h3G/NOuBewMBiWQkyqdMuYSa9se+5pmKLro/OlZ8y
0GQAsB8sNNUKG9/TwrT9UO+Eh2WjQ/CWw7ye3ZQV79dGcuqd8clpmrJNaSnEx/IY
sRuqTe/GqURvm9Cmwqx1d7BY88NyjYjkHTkaeh4837p+2h0M35vVeg0AX+uKyJhQ
+Ossyb9FncmNtrLKRekqykI1VLaeCLE0gTemYnS9oU6SlHifqygadIoC69EgrJRU
n0lPrGivY7LKyFJ3K4lp4OtuqXLoZ8Pcd3gd48wr6tPDGz9QU+4rLf3ha2s3dN08
fk+IxtyoX3qTQFJcIG+NwmRpiYgUBrb4G+5HzxYuMBTZROM/HFrr2x7wb04Co/jU
NeRmBubUveVga7YedtjSWvVAIf+tIPABrAG7sV7Q/1wsY0zyFDzjRhCFnakHNZGM
j5Z+7wYgN34AQJVoHpyXXD2ape1UHuNYbqUkHADctHOiMVhghlkbCHKsDDWjyxqQ
BZlEuwRvkT0hBDSFLaxGCx5GW6aG4nRRv7IlCoM49+nMfkMVB2T3gpVGblossvGK
T1QSUtMX3fkcJtHvlu8S+ENiuCNJ1iJdBhgfxo4mw5VS9irdseEGhtPdcFokPAoc
6xV05DSCiFlVPUgShLZq54dmCiHQD0Fl7uebfA6X5bVzvilKUW3SFJg0u6cF45XU
WP3NDOIOjQyVwuTOQc7bNtz7EEvsLzh7sNyqh4qBV9r8PTOk7dXM/M7w0EWiWmlz
MOEe54ejmk1J6lzHE9+yA+iZmbXmrHrFC2H8P7qGvYU7RA4QEU4CXdUY2OxitCT6
qNw3fd95aw03MWuvzK9utQ3K3xCHp/yKOPGLCKKTJMX82VbJTif0waSvZCeAjQAW
I/xFNpKiFbAvIOVq7WyCWtNDnE4b3WiyeeIWEH0s+HPMXC0mRKhiMBaDh0rU6eqs
4FBd/2j6vflajqKCPrPX7EvrrmrSdWu4E/JrsNm6vD/5NiGXxHGtC2e5cMFRe7bv
BvEKcYLhvnGJSWuDip2xBqSTd2rG1K0ntbowvZbZX9PPx0UG2gOn5d87AoC/v1gS
C99/xZeLFlvebL59s8F1CYsfl5Rn/viqc9brKExJ9nZ8HcWh9ZAStyhqiXX5jA0e
SqHt8lJuExIurh123KGl4jBxtgo03XdEaAje+x9ALFpbmItdKjJPtJblViHwrBce
B3+wfRX2ae+Mn8lSq75Pr5gARhatN+QvQ9XZMbXFiXRTSrWy8XNyKVr8hEGBRIkq
2DN/Lr2aEnU3+R3dv2ePRJILf+282KC7Cm9+LlpP3GeJ2QZMpr+ohgdoBdNmUVIO
A/jmNW5CKieXsoYcqhojqr7SuTQvJJXkUZDjQiy+N0UgMV+knJZiQaxmDMDDBZ4x
P3n7/9Ka0OiLidN7qe42XMUEp/NJxgSawHpGiSsviuYV8QXclzY4MTbmF/kkIx7T
/ufLCeDE10l/Zfc2fC6WWEajmDomj1n92w3eogS41oXXbSYJwrOK1+tQLSpnwXJo
apJE77ZuIdGIUAu+2Jq2/wGwQeuj8MRgJ9VuqMKkzBQ0A1rxGze9+C9CQby3k+fV
I8Xd8mR4rATiJFgze4xn5U7DXg1mh0yvnNC25bSbEtY4BORkWK8d2+L5XYXknnaa
dMOu86gJ4Dn/vsGmsijdz0DemV52EZJzsKJJ/jv1S981I2tSVJ5PpYsCBNwhv0xu
gmHrWJ2g795GNH+Rooq7T6RBpQmdXQmnuRilA5uGBkj67ojddaRuw9azUz/Pawwk
gqgrcFnWTKQhY7JGyypOLogMjAUnsvvKQQHc+rcDS8faI0rd2vQnef65lssKCz60
Wn69wpYA6TLjT8efC0n3OSE05GyQcBXk4yIblUmNT58aEEl1cpgR4UM8874wLDDC
b5cEDwHTfLCfxFZwNY4S7aZPiq999pJq60zSZLd/O/tilHEvBUw2q0vZY4MGAnfa
2gCv21cnLcdcZK/hCjkJgpt71Pg/G7xSOx+VscrT+z6RjEpi7LQUJJXX39izg7Wd
yw8Slv+ixn7cnTB8xBhspaHJXo30cLH68J3sBlrlQBXiuRJM6ifVLDWAUDkTOWvz
Hy5QCs5UxA8RUiWbFhEau+LGfGJIem5h1Ze/XgV2ADYVBDlcWif5llHuupl6Z9ZI
M824VCk9fodaBp+yK68wnDk5/BLjyhAjmLmcSmvWgtcYxzKrDs3teSamSIPnXR+N
34Wa+DpBAZTI9cuFxSMRWiIaPf/CNX4wZhCrbUzIvrTgiC7zKJ59mt0bGymkV6ey
8ZIzJq5DbRY/D/7y/VyVBsHpFew1uagohwGQhLFz5zKgRQGKdNPASmLqD7kV9VVB
sVZyJtGPhoFNIeo+pVRNqUHVQ/tVkErqZnl7SCOEs+SD/repM9UJzfOTbDd4M6Bo
J1q40hN68ccrZ1rixx2luFtDPwIlNxW1I9DH/GauAcQWg/tpyW+a9T7SD4uLPDSy
kzptNFp61Kl330EhjL8tlhCzIQ1GKhPZ4LAD1HcLXJUVEORK4O3mIkr34x8qiEa0
k0/pUogpWUyhq0S2HrjGGNSzAGbs5rFZf8EDjuCw8pR7am9kQ7MP/so7Zi8zcKh6
j9qF9egVzTyL2jklktqN54TZDb+PIGzaAK6nengba2vAHGVaGBOVCybn5qAr3U0x
F9Y6gQ9pIC9dSnMW3ahMVNbGLFD8vr0TSRVr2GU6hAsGG2onWNVnZ/go3ZVIFm0h
fXJEeqT+tNXqwxjI32X4nLwnZCrByS4eDTd2592U8S4wWDfMT4y/H4W/nw70ixq8
+TYwSs8anqh9s1I+vFDpj0MrpUY4mnVyzPOZhf13sRXUGlVNN8B2V3V6qXfvutoh
9MIk/WCAj8DR86muHkGx9iE2vZXNq+4PBKU01zeMl0AYuZXXDttjjSz7yqD0ty8z
02/Iiqh/9ao4WRFNn4s5UERG7UyWBMXJIwU8xhthBUebVWVOz6PQoKE67sdySO9X
l1Nt/tvfkDpcZYaaVPZPLjvQFl2hpai8GmSa8Phchg/2kfPfkD6PZzyzKXzJ5DM9
3CHjs03apw1E7tmE/h9bXDpEUd2sz02hxa7Y3q0l1TDTd+zji/Rrdjrn2l7sckjw
AnH5AABPb0WSksjDS3rAt6IWnEfG7SLTI33fMg4r7NYX17rGs3tgHb3ESkMHqmAN
DTa9Hog3CZg1jwZdpTwATdPcqN7TOsOKJ5BbnCrDJmFzKgLpxzA7LG0RgQ2B2NqX
AhwmcN26Bt2T83KyvNHyQGFItdK0hrd0moBGV1lgChTrK3AEUnSN/2ORDZq8mTcb
b8cvidto0dbdliiI+lynWQ/yAwg0EGvs6IO8RKO9cEIIexcRtUDHRucAEja7bE/7
DPAB75nZB+Vjz2RP5FYWBkqxhYmSzem8zTkXXZ8uWubnpJyNMaqQgb+xL2SH5tNI
Pj7t1NhosTDla5+iwPvcxidUjMXlus6fOTjPLs5T2LfKO9zUpQmIS1kn3wfQrsEJ
2rrHpILVhOpt1y+kvtQGYakqQRCmU+8YPLVtmqPlOolRdC2SvNH7S6PrVFbwqrRj
3Eo2qw9rXLWCTPN2Qcdrq1iD8LOkOAuhs5DiatSH6eu4KTkwG0RGcFgSgnGt9KCx
ax54ZwGVaVris+wKAsK8PCmoHoIokMuhQUuC4fe5EBLbOL4OPDhU/WW57LhNAIwd
aAPG1l8vHV3mm7LHRvcb39CWcrhYK9Mz9poVjlfSN1wfaTuYGnuPbWMwSCUsORVA
ndFWWI6zfS7dV8I2R0qK8uJ90B3ZLK5UzROCUv6T5r7aJS5vQjmFjx+IrTiXnQZz
ffIl7hCwaHFf1ZaR4a10X0Mo+dzjP/4XL2Ocek7U9JmaZapVdfIdqbPY0bsycY66
VXazKsXu8bq+JAOY87BM2RXvbK2KKdBlZyhfCo0s7HHZRjRiiJsajK0RIIL6Wcxb
oBxHjbyQY43bmsrIG5ezGOuT9M4ahH2nY3MrXsqt2ruhL6kdQEUZefmoVGIZ6yI2
zcnt0r3cNv1HWOvAXqoR+/1YDQRxo0PvW2546QQD7ku5olccabp1Gm8eF42MJO8r
vn252DcPOUvui7H4lX1lCVKWMKY1FfxQyeUNCD1dfBiUGfzzHVLTKAxECpJSKoPQ
WsJD2TEHxz5l0du01u+RN2aR6sD9IUovdGZVLnklMci+je395w/6MXdkv/QQJ2Sz
ZA8Nj9BXIAAmWRCPM05zzF/mOvX5rQHntXH11dR/+uTHXZBFMdQBBPDry0dMHzR5
a9gPBsMfw3EDz86LMLBYL70CfV7ct14CDNuLIWqR5OawP2R9MVB/pez9pyEJDHvZ
RsNy/Cn1J+kGtOJnX3IucNG8kyu16/2MXBTt+Hg4YTXXccgWDHN1Myh7x/ohMzpa
2FxZ3eMhmyuWAVSs2jk+gDPqBHaEwnTnIjfiGXPsOYpN9Xcx0e4wNPnTLqZESLN/
bAoG2fmZzTjpaT21tNchfTx7IPBSWjZwf1rXR3/MwXx++qlCs53QcVKiJGbVgk/e
UDpxNkW+3l2uvf/D+IXteBM4+QG25x9G5w5dxtqWHMENbOWIRPrS06TnvK/DO0Ix
I3tCQwAHdPSeIEHu98gS7Zjv3a5SrVpjCY47iPVRuiEI/ELKFerawiHCYj0w75IZ
B0rFrVM4MOCTYJyQ0kozKtENXTweqKSi5+zvuEZ/wY8YRjczGHMhvUjl5gM7mxEZ
ziK2Z9kvvyLEVxwdRuzpvwYFuhXd80LGOHg/EhuOZig3P4CoJA3aXdOeM9dt6FOT
aorcLA9Y8yOq1OB2U8vGv9OgeqYDenP9bm0z+EDMZqYVCEDRf4ubJzgklM3NSk8Q
GIyrkqu/xm8tz80zyFGwE/+ja6f9lHWzzLIqX6fZN+Xd4T3C3EAfDo93cE5ZQqN0
w5YsG1fl66LKssmdgY51v5isF2XuQWZwL/z5kcoFfGuCVNbWyQvTImU7dE27JxuE
/z8SbN1IrV1SqFvk0ByHTilQ+nqay0PNh/JIU78X4+7H265HDmvqROlPRHWwWxSQ
deR0jXVoOBD+zlvuplRgjuMUnrf9EGtwHO7Ky9nclya6KF6tTpQmmtpDszUE4Ham
E5Kc1hREoBOimKDfXq0ZPR0QWJ/UTDT2bSuQ41hMr9UKjfYo92feoP2AIAB8BihW
EXRb7fwc1sVE6vF44AWC0ct/Ce5Yk0lqnFpEUSjLWxn4SIEfwUfd0FyoPwWGnlMS
Xu1M7/3YPRjKkVSBMpQ+OPRVgvErE5Ciei/HsxqMDMXjMa3pYQcVoKu3Ruh0Qfje
7p1vOFykqknkLTVJ+mEFW0KTBqyGRjjLLgvzyopWwskOowMHAC/lQ2X0dzVZKoBt
Gt90BBsqRAh+xzmaatn5A1/kMuN4PhUmUsYJQTxB2VJUDA+XU8Afnw+cjSabeXWM
8U95KXRpcdxAogJvwyqXhJlqckPoRPy8l3SnA7lLlEWeVZ7naMgKxHiZkSHEX1U9
rBlX7Vpoi2FLlsVdXWb8RJ8GwVuPLFVtGDs7MrKQrJOZEt4hfS6sDm6zMQXW+BE5
+k9xDO3PTm0FTuUNoQfNnDmhgCLDsZLOow8ck4h8/HHrRvQoH8JbLCVgfasE6w9N
4jwSRr1dWS+qC0GhNPPvWBUGdGL+kD4vkXc2DNRM7fJgfny9/r6YEwC+HhkPksWO
9POpDVAb2ycYTp6d28bGjGq87MmXHchso/lhXRA48vD79Slk6TVdjVPJTY9Fap9f
DCb2mE95aP5TOpBUDGf8XwNdD/Vgkw7WoK7CbKFIkYn9ZLCYfXHVKSjHcWruJxZP
P1FSRR7MTrZY9pqXs0LwWZC+HmzW3BYB7nvd/fJmubva+cmvP1PYGIxYGn/TwbgJ
UaUIKuSwREnS2WWw9sut1mV7H3NDz+sBSUQglIZvOvS7BFKyw9T32fgqANHtq8lt
1RHKrO8+vCJoc8czmS3aVWlVtJIaACfs4n6PX2jDGHbeAY+Dk9SyaCMjOwDvbumN
G7vqlISvlWf3Nv7bytEQowBrQn7/dyKQJUBAfF7r5OzmaPFy/ayrJ9vq3lukJj5j
PDB7gxwmS+9jPx2NebC9V2982H2h74YFyWJSSihgF4HzrIACILYjhkQUhBcq5RiO
Ef0+A3jILitmWL7/eFvBde7m/X3ehFgTue5U+9VeVB7vv2fIfRDhNFlAZzfQg/AA
PSCYWoG0eQ7l51TeYdEC9q6GwmTZeEMh4srU/D0aV3y9TWuxnfz0WmFp3jEhRBkA
zZEhaG6JLJ16gatLL/No+ILTT/XYy1vQlPP/1pfc36aEHmCAnkKj4SuZw1+fSiF2
UrQqFnxU2XFWg6K3QJRxnpRvDKL+mRBSdeARwYQl5RVBltZOD7VNfs3vVwDuh7F8
Tqj/J+3mCkn1P8pPdRtTfidAVKaJ0F9cuwfgTU58Xg5zI8MakkjBrhn0v4mxGrT+
oo8LwUpdkVT8uHCopYEX+l0HT1fg+tLtmQgH7ca4QGh1mYPHdkWpeLTVpb4WrEp7
srF/l9wiG4W+FxqYMXV+Dctrg7X53PJna+dMnvuRdGN7cgDlrgefuQ116Udphd9G
zMuaTBOHwh3qjFsrQbYm6TDkSZRDJp/HIRxH7OJ3FMcVZc3wuprlFDRp2acW5uEq
ipWgwCAc8/xS3gPjZ5LqB5zoxrtezucfEq4pZNZL3XHi6s7i90aagKfYiuYhAVkf
YYJrlatsTYMIpcHarZoBaStYxRT2xboYdU/9FRR6cBhWQX91XwLuQTVNIrn8gXch
JDJnnehJYr/VIuzM0CrWpklKsZr18QVnR7N56xsaDP3QmbM+/bZ33SPEV6/hqcdQ
kt/ScXehohqnPqaV9ZlHNWMeCCrA4mb5HZ9V8t07WGoEJXKvMv/STGb+cuV0nkyU
v+QWwCjYRQVk9kSmyq7rf8BWBXtjTylmcJNLJSp3NxPsKOLx6b6XLGbCniOjAjVe
8y6tslprnZKxyZub3brPDjeqay9bdKizs3mzpAWlRrPeTsNmLegh84bT/LcGOU/+
d+JjltV8G70lkGbFQBnSF+GJdE46ULI62VV9ooeyeveHFu8oI1duDBJGFHWh7c8s
tbRvUQfPZrsfLJYgItClC1HDzsQ3X2uPEbMQmQBnSwWZCd2GWP0gISckCnpSH+4N
97Gu9zAU8mf7D1vy83p75WIjldpWn/e7H89629nn40SWRHXf+iQ8tWUOwRdYL+U/
BF7Zsvf/h5AFb3PM7hmmAByLbBgyki/81HAKToja3r1sBPTCQXJUSK6zi5KWlxgs
82HiIUCF2rYYsUwU6FA3fibklhgYxRKCA7rZXwqy+fDE52n74Dpa+Vip9lvX/bQR
uAvmJ8b0+vVcUP7yHNCbDWWkIyJp5l2XFQWMkbPN5IF8y16v14xFwqUOsPDjUGq8
k47UfZClam4N7WfOMV59oE2HMWr4GC16PsDkIYGiYvKOtgSs34+WOcrRR3GoJZrC
oDcfBgPVR+WNoOXByAjnyStp77ywmWXfZbbUcfwsqoHXY2IZFWaluGORupDChwkE
HePSrI5iGVvukQooXJe7P2HmlHRzMij1DFbcZlUpAxCy9OSDeuiY899tucG8J1DW
lwbU/IPgXD7qlvxP+AAJXtbjcFdAhU1BhaQsbSxSMjr/HTXSbFTyP+xe7rLSpHs/
/DS9PvCRJ1myZ9ugY02HDq2m6NCM1c/drsAB9QV4vaTBHkEGx3uibZyfClhNFDgO
jIeQeqcjP6il3Mpf/Mck30AX38GhLMJonvongqGeM1u6WUYLnWgivkJc/uEdVx/g
Kk67CFZFMiOwjsSYKN79AF/X/RLyAcf4pOHlbqVrBXgNQyq0N03usriXjzJ7DqgK
MbwgZMVWxACz2ebsOrdc/iOEHkcdBtY6SJhlQBZygEltnHuz/D1FmuJxFz+xCKOF
Dl1d+Nx6p9Vz4jLyc4uYsjA/HGHW/ZSh7FVBlqg+UAKRJKGz82r1CqugHYHEpETg
qUqNIS44qfCRF/D2jtO2EfbJ+XhIgGhs19IXQFv0D4rpvxeS1s5TVdglW1Ribcy1
7rXNO9/whxPUAiIpKCriA1muZploOhczlMRSf9nC1YH88iAej00q4ddqehJD0mTT
TBxiF9KcmAa1jBaqw7GoHqFDalHv4YY7Hk+sO7aCJIPBQTixas/BlBs1037/236q
3RZj7fK8zc+9GtvwPVaszfB5HFrAlc+9B2IMToE+8kp/dY2pzoYI/DamnNY+208i
kAf07F52FohRktFK8JkTVflMj5QhxF/wU+UkwJD54T1OuEKvjAYo9YgoSPrAaF0a
LL/7AG8Qx9CxQ3IEBI1D9+vFEshs6leE46e+TjLdDXNHnHzDEqIZXMd0e2F7hWTW
qh5ZkBNsWi2CGPPKawsgBTs+v9aHNRrHvGt0A008jDXPUwEYgBg7Ss8CgY7+AcRs
njI6ZDOmmLNunV+8dTWTLSXMckjccb872ncRwDZIqKHUj8YqW70/DgQu/h3xt3fQ
YZPblSFQNpemDPLcZKzgVyknV1j6ahK1ZxgUODPV2UD5xxdMyeGPkuxrQA9Jwn8W
akGa6mkSJk37d5/PSve/i6W7+dkhoO5BRjicJF2iTcTFzrTaw70GjkV4U/h05C2Y
NFn54ZM2vmADlC0dh3QCHq6x86sWk617Lvw977Z83bQjbiLlvAePR9Moi7sVrulW
z5s81gN2UrDavqchLShlYeVOH1uZeF4vjZA50txQTJ8TTPyZdD59iq2jVzpHfGqP
kpoMydG+SBuhgspToh2QcMmsu/XNdbWJmlV2gPcT/RrwTmXLvJ4BC67u78SMzZ/S
jVdkO1+JNupY3QUe1aeRL0GknLNdNeOtBejQTwvpLYE8g+O9c+M53AcZlv0fJ0qx
NSdw6E/DKBb9n8Xt038ZIDGaKf2wqVs8N2OJ1A80AtOTgDtRqOw/7s67uph+UD05
FJefJjJzG4kzXeQjm8xdx5BrYnFst7i3EhfxZEW+elV9sY3wQPjZK+JyD+PkB+XO
ZVVTmxQMCogicE6YqLRLATvzVF7ffyaMeASc6k2b4+3iIVxF2closaXpX1oOGZuS
3cSoZZuRSa5jkj1oBioAO/Ob1Rx05yt5BUk9ez101AW+J22OfhfZDCPmQ5AwD+1h
cuk3BLNe9tTZdXYx3ETra9AIfy5dLWv4oAjLgzK2sAVFw8SZC0xUJW7tSsa/G2fQ
dFE35tm0MQGL5B44Jzm9kd23UmMLxwdAg52IzGPSQ9p2mMsA87w7TompTstRK685
djyaJ8EfUclyioiFfYW2JuX4LipVe1FSpnhxm2NIBPZ5FGBybzlsk9cE2OGzu3Y1
xJMyUvTZefVrHUglF8YxAXYxW6wGifXL01fr++aU2cSuyeZZ4A4fd2WT7rt0lzEY
e2m7O2qmwKCG4c9EHQSpoygoLuvFsoEMqRZqvApRJA9kiOwRvPft7y08fkQzC9cC
FJ0PLuipgWsAzIBt8o3dMO/Tt/zZCeASjgzGEtGu6uB73oMW7xTwXB/5iHFH4MwU
8zfBYBrHTqbPSuoHd4G7ZMc8F3IFNCE2Vwlz9Bu05eBNL4cYHG2nDERpa3n/5mU5
FyVmp+7dhOPQYX++1KcbAWlUD2BuQUl55CZVbAxAq9Z22gRsrhs9BrgA3d7NrU8w
oXW62bcLwcrdojEsOARFHf0MyoaYlGlJk3QxYUhUXGqQl/qXaSROeH49DM8RiD4r
R7ivum/LwcBijGa8jcxlkhw8EBsH23F6VbDCuDSYi1j2AZR1r9XPId8bl6d0+75Q
+SGP9a4VV3+tm7DIYJiVV5d+N2aSm3e7G1bQ4gwcKSTr+KFUogIya3m5HlObYFv4
nbsU9+Xtuojvmf3cMiWUUHwccEDqA0OADSTOOAXpIZfiErpl0JSADKeW8OHDwRji
NEV25JdQ8+qa9KL5EB2UVdefWMCYsbdI0P1FsCv/HP9wdnRM9Ij80L+jXiuWvwaL
O5hKOdCQ9L5NNTPCjbyvjwiC3ANe7Mf4qYr3yqEU7Z4BJs4MI5iNpbV6mZy04t4q
2VKKS7ZQKDeMHzavgdEX3p3DL3AZ7Vvwr30AoPpLQmzgLiYLgs+m15kWQtYY26ML
0VwhjaQ8BgG0d3Zf8jKCyGYxES+lNpM+VOAubMAYSFzI4nAaEmJZZAJ7wVPXhH74
NZYQdLqGY0FIBRLWwSBOglCslgfbQ+gbzOsHKs6on1bjGBfsfJVXfnSuwqXYPSw3
mdcCqP1T++i4mo/D7XD1bdVt+WufKSK+sjCWD6lLJMQ/4SYcaSg3sYhYcTl5I08f
3RZPs6NsYAlF7iofCdeoPIYnI3kOKEtipvPI1NiuKQY+TDrJFSQZkyE6BNTaQCAp
OafDmDyw5PlERNPjc5Rkqc1QMQo+84ibJpxVUSfCa/7zbrZPb9Xm2E0Xu962uJhF
Jcb8Fs+3Jg3OQxBQ9q+LFC6rO6OUj6FpdluuYxpPXWL2jvrgUoS9Ma2BOesLnWKg
vYzIAdQqgIivW9dnDbIgbmAzYCxivq3EEBiv3PbTkll9uB65Kk4QdmyPiuBuvSbt
bJlwMKARVEOA1wzGC/RgTF50ZkyhEX0m6oyzcCKRdlR5UWskWakok1/duoZWcInc
WSdTG+uDEdqqXWvwoCaJiNeZBlm4BF3rAxcFsVu1GIiSehgT6hMLD/mGkS+zF9it
tdQm/c154OyBZvwoxNZMVo2ptuFxVG01KOcDtrRXs6Lj8jMly4sTSbwkprBDSzVq
2A615341QXZyS4LqfmZSJn+wzCrO2EI5Er/Zwgzadp6KADktTuA3ROeryDWwmtav
EnazfTa5ZTPouADkD3DxjNeQurOr92Uj5gntXGXzaVVKQFyPAneCgaDVtKRg6ZrP
zSR9X6di7rQiYGLfkMJXI79gC8HRFCrA0P0g5YpbbWjGkASXtGZwOUrQW8e9KKdi
0bYLHXjz7eXVMgoog42NTs1tJriZ5ZBl/014SoR6oViB/eV42jiK3l4yc4vndzwn
EUuGWuBdFNGiGF6YG+po3dYYgaFvBP7RPpi+9Hd7HHLlESo4+WyG3ylfjR25TqYl
nUAwxlc+jR4BA7iMCrfcw/J0GLDqQoxLZOKip3K+LM49lcI3uUjTHXgtP78cX/Q6
KIUBZqcIyXsTDwXJIW8DleIC8cfpr+s7tsulNFmPphsFSoG/vMPnQoPnMhz1jtFA
VhMvik8qvcsBJi0Dgg9a3ginzugVuAkao6r/OHPh7TinunBdJ/dmFwCwoIe3v3ew
CX4VY4oQUQ6nMZioENruIZ8WaUVYMnRlPaM/iEhctIyTDE+F0l63HfHfZfhOQ5uE
EQZyWYyXqGjFbjLgtYhuY9eFf27PLZA1X/ENrIgVDuzl56GwVQ8wQhwej++g+v8r
ZAq9SmsKZE3D0JQt7XdJXVWVjwWm7iJTv/G6L3a5i5tyrDNtthW3BlkxNUtp4hVl
/Yi59IrrAMqbaQ8vcCONpt4Gfn5hXadfiR2OHbPwM4nIY1Vf5lgYES5j9BagatQn
0ZsjSvHeHwDcrfcb8VIwyiClALkRnfjO0DcGAbTbAZVvj0HtDZuct+4lDk/EotMw
lwP0bYDpeg4bED0Kn+7AVrYGCy83GjLY8KsV2vdyTPGOzVysnxIfH06NLdod2lhw
EhtqmHr1WUd+0U2cCAzPqPtBl1PowYdJkVdLRa2CEsplkD4eplbp1dyh6QspjpQt
SJOJXHMwmP4Gzta0rxgE9mQsCuKvzWHvkaE/PxHYazJ/nmf3aLhUi8Ify/h7dOv/
WXO2l9B2oDsd/Owy5CIpXjA3ZCKbywCNvBqhcfWcGLAz1OfUaIMWHLXArAyDaqtk
iFlS8i9T6ImV72SCGLHyIlc2OuaNpiAIB2xXqj/eYMeMP0I4e8eH93yJ6oCXmjPG
9epSYDHAPhNZia/7+qo8pgHxcXrHP24FMH3OrxYBmFUMBbtDw/doltGq/d0aRhfL
K5dJo7H7xp1/5khaKNt5LmiAmgCTm2W3FLlZmmvVCDTxBH2FgAHtYjYi4fm1nZwr
jIY8SGMEJwS8ohqu9/hTucwd16xk+0CmR6/Vl/2F0ubHWA33XQYrMCdmjXkYCpPN
ccxHFSxwQyGB2wQfdV/9BiE04QSudiCl7o2ZpWZp3J9op5dyikGFDJqoWQhb8Ud0
VY4snrB+dHxeVraBoIZcPNuPZyOjGVcdgRHGUkXbxkj7Dz6UJaPYzeWvNZrtYZ4W
dkGzEZGkvml4nhHGWB049V0If19xctcjWDPnZ7bUm5uo6i3a7T2SMmDWpl6iDfFL
1Je2F3yhD25BCUwbFxPn1llk6PiJvN5iOsM0qaitaXcMSgjh48a+hz3OBGYG+DlF
Z9NaAhVwpBje9X6BYjTOO0JktuEBmXTGDOBT7oywz+9Ijs1nY/zXAxdP1tsj6Z74
O4YqlGr2K6iL5cZTeo5bmkclkEzSM69H+xAg346TrLwfxUYcg/B7Ky/T0SwmONIr
GMNXuVXG2rf4VTVVc5hZyz5gkpjNhu1BJayvN1IcZ/xr7A7coCJWNYT6B6eW6V72
kFNiEPFibWfUBm5wMPlz/T+0yoVOjNTJnPCn6MX9YIWUHjhdeWJSUKywdWF6wFHK
W17MJAeBe+7wPXRuWBJMh+hzn6k7QNAaUGbaOp9ljCdgo07u9m3qMHhi05erQNb3
fnvbvhnniJSAtqvoFoIpJ+h56NyzuRq6iN10LwNbvqrWF57sonrIPJdg2EzL58lr
q4STrqTuCQ0zuOJBp+bA5sKgjmsIaFVJh+K5tJpvH5PWHtfijaGlEddUomc8Brq/
aAVER9gRbMv+Vg0e1Ip1wj6csOxnwdxFWAoGYXjvxqot7fsmRkRVq0fu7rABvNdr
aLBYXM0cdmToFImbSK1G6m4GwtRfyhwIju26uptapHL625nq62U9e/HB0ptdnMZ8
lnObCo2TvHdWOvpkWthlnpfFMyYrbfrLi0IcXxVZT2Esre5Aax3LVKBX5IXRn+S4
KVn+wfISqKqOxBcQp5nSrKZ/LCG8Ksbq3a0Bd3pO17VIyUFIv5UL7grfSkvyvkMv
WBDS1xKmk+RhMi50Jzh6v/EUe0sd2SWwTh3izXw8ZpSihSIrQgSHZidPbInrabxs
t7qF2wQwEYOi1o3gjiJYHc7KY8RhXO4o727Q9P/XzknsRXWfz3nvY7Sdnh0IT6T6
XwACzvdF0Ie5kVVwnyz3c5msL+ew1b0NsDhenPaBh1dxOTij4CdphkekPRkrLPvj
+3qym92sd5GMZYl7a4OrPjz2/fHg2Qd6MTXvrJjQ484PHyP7XwhL7u1gJSv4OeMG
GnmRabNbKloOiLQ4/YC99Gq8esy/THZbSA/21A7p3FTlyaTMNlIfeo6q/nDNdnOp
hBtOS52EzhV3U/Atzspuv3CwnTLaT+aVyo002/ZJ4EJBQwlg1v4dRKBxIqLnc24r
fIB9PxsI1UpngHJAY+fUaI4pwD8/va0Q2o14r02F38n0IXOlBLJHuP/+jCSyvhVJ
rq0a6txTK1AodOKy93w9jwn9mr+JzXj6UMYqeZUT7l08A3vFLhfjvQEMnaINzGz4
aJQZoP58pHCreJJMwXiofTE0nvyCdxkbtXSlPDO7T2wbcBRJUW+kdG47lGYt1L5X
Vujz80fA8uKcP0i8Hjp/bPJ92757ka7GLX8yL88ZvFq/qg1lQbVRPvJ9/btF08v6
2KxvDIvIxDUv1Prcg0lLyICBDGDvCEcEoPowms8BQ54gvhwk6F6lAi0XM9dPM02Q
3Y9VsxKp1FuSI11Eb4WuV2he9dhA9IBXNtXeQyKUcYkQJOvgnvT/hL9BQPjgG16n
5JEmHRa7G0vpqboy8U0/zTKLnNR3duhU+w8fU4KTDm2Oygr2qGhMhNgHIKIyuBwT
hGtWc1pnXST+V0Ilkj+jPq6fQfreqRHzffERi7T52NN1nazYCLPfnjfVZM0VLYZ+
JQp3IKW3QVqe/hyiQvYyomeRJ0WADHRUbSAkwmrQVkL4WPop+0Z7wzVSVcyMOLMD
bGwKNtmvO1EEmrtE/itFIOS3pFBrZpCcZt8OV70mXfa5uUIf/bXugltZy4wgAbjO
QK05F0tfSe6k2KjwphJIsHds7S1xg3JYxuEBvmMtMOjIsSV2ATLNNp/mXuGCERID
TdRDvIy3AkkOiXPDVeWvqFiSxwKPNK3sq7uOb1Zt0OjJ6BQhNfr9YTI46iw0ZD50
tfEeCHNpYamYUG6EvcEV59MDBLxSteqF5mx9wOdebeUIhdgGPlen0u3FEcqn0rnw
pgPLDTBEFx0r//hTnxoGg1pBkbcbyFRL8kSRnrOQNdGJz+lIFUQ2NpgNzP0HJAfI
4PK00SZ/Koc2iyjVsT5SpL8652lBXWkpQ/Kdh4sIjtjYf4EKA0+CsI+2GVRK420W
+5VDL2QqdFT2LTm1VHt1glFMjPC9RPB0DAi3klT56qMEXQVo/yzL8IO7M2gaC/cW
nm8HUnvXZA8xVoKBbKqKcPEk9x2O/RY+a/jmH4T1fGrAVSfYYZTH8dYl5tT5OT5h
gDpvSWeNu5yyBDL57PcIwriMzFxJBXkBVyW7lGuWPoFf8QKUPfDxaY2rXN/EZwED
R1M+Mvedl6Eoch/OWpDyqRK6tZAxs7DrPLsLHRsXgVqmSo8+9Es6C8xip3rso/Mv
qwZOhpjZI01KgLQQzVbL+Pjx+RakWu1WM8qErlwRrkJC+6aZe5t48i7WrAESFcIK
fsqt/3K2EJKyfTMwXB6/o/PsJMBt6zttOKhw1DbxXKwvV2Xo5/xcmapV1Kp782Rp
mvvV6w6jYRTC1+kFCJUptzSZDdi8FNCdSVVJ7bTK6oXX0LMnTTO4+gPxVZGZpBnw
qvBAMneXwcMPV7DftcVc2XOv3tmrDhoG9Q6MtsQWaT9b9RX27YjdXtzeyJlIAkaL
cWJopgIngTZsTqNrz2EQRddHwgANJSQht97yNl2XUFOx+c3u/1JMdWSrTZ3yrWXf
BDMD4qx7u9MqTlq+4mqCuONFajfrkZFDUjEF290FFeB85ubkdL6f3wM3m8jkm6lT
gpk5wHVQxgZSyJ6DcjSbwKPSiREfwpuCvWJSMT6EITwlKwmK6fW6E2WINf5pJPAR
ZQyOET6koZRGRIjgM0Z8Q5aEz0tjgHf5POzq1rixeoDTGxaf5mhtz+FifArNQdgZ
J65GQtHpvvCmGTqowWXt2BQm5UA3SdhX3lN2YKK42jCIJ0aYK0VBdem3OA4q76Xo
vt3WM4Kk3DvCPmTGK4BiDs07KNL4V26VIZxo+PXmgmbb3EWPolLWH/1uTcVnSDLe
bH01c6X2qRKtI3nrb4gvydOwG+46mUx7jwwNkKI+3R6AeW+/pOwei9ssrsbXl4o4
XnafQsHvYraq0BLzjAPQK2BNzkf9ml+q4YhG3tJIuGYJGTHmwykKkR+1vQdM8wV5
pd7NUL4QYzsm5p6JQ8i4PdvSubFLHtPucCEUOfcKPrROawhj3a3Ni3F+SEEDzmkI
4jcMk0zh7gYnuSWn/uP4tEYkZC3jAtxGybh3uqPy3cF+8qLGjXUxAEypC6HAyIX4
2yTkWTII5JfsPQyqOquEb8H3pIs1FbHMTxE4ftHTeevBIxbXL24CJjUlqT+EjLdQ
A25CgqnkWOD2/JeppGkw/nYdtFvt9viURiv+qYUWasvGa8uDcusiXLRrR24XV54M
jt078ESt187W618mZNwoHN7gvYr1MDvjZE2n0/huQJvHI7zdJNjHWK8cS/6rSz1r
ZqoZQyt9wK9htYX8c3g27e/wpJvtQNRWkftYmnQiyHCtwx1lp7S4UIjzA5dGAItq
MI9QrOv1ZADVwTKmARqXb5jmUfc+rrl/obNKSRhFme6XYZg4ZEt5LkpoPzUNPSNI
kpAlhgKY50UimDu/KZ+xnhxKlrWAISMJQVpxB5JuNtigjF+fpFMlcsevRy000Dz5
AoHeLgky228CBiGLH4N8zJ0aFP8SCuwfDjAQm7TUQa+AALwdB1yRxVfZTc1JcA85
vDoXEvZ6kxOTt18A6KPpP9rlZ4VV9g+beRWiPRM9gpHO8kIfLqi4q8YYpIupdXeM
UuR6tFtCFalhf3fo7JpPHb7GwriifarypSaROavh+naw8DqITGokSH1Vkuspou9Q
CaY3PSD5a79unYHlk8rRD9RFfAWQfBVDEyDOjm1VxFHD9Mcs7U80C2lLM2sKLTv9
Fd2wPH5S4e/pWV5MRYgySIjyUVQW9zTKhwgimyzqRNBWt2kGmibgEKpcPvf2E2Jg
2tLUwIwZyROMVgaUjfnghahleaQ+HeTad0yQY0cKOtleu98gxeOr4r/c5uSsFa6f
PUHuUxb85TYcZZ5Oo/bPIN104Ig8gqMsx11wpIZ5vRr7gcWNnmgjLnPLuu/ErsYe
mk0/zm1Z+BSkLNj6hiBDXpqynhYozxpXQlJ6I3NQyfUHap5GfHvSjq5vSLanNjK1
uQBv1DaG/+VLZWtuq+s+MsWIjjziGPEKESPc/P2z//SmNWMiRqYNAAFmW9Ey8d3M
pKvkG+EGVABOQCq3bzk8jsmcKVdFm40KdcnkgNL573pzLUNsrwj7+zmiPeRqDdd6
575SPj0poQgfyqrsB8+nDi0Qt2gzYtHqmxTH6lT/Yxn2pOlTumxD3a29SnLSXC/h
/sti65QpEC8Qo+SbpHAxn2vwFl9D0X5KZYuwzzMzN8LUgFZaWgCYQGwJO+ID/ZBG
3rZec4lO+ukLiSzT0UzejylM48806+YIsll5pMVbDjtE37xdSRtROh8v2ky/SfKS
zLnljTGQvUAfrpv3K00sFbpVhr+uCPp7G9icNg3oVtTIdOdD7qmdnZOAaJwJcnXv
KpOWU4CVor95xm4VsQ7eRciFCv0vu+HsyX7RIvZbmmB/4s9xwuHcbkfnkabaUDLf
oLBPy/TkFuKf9Tq3GI8+TUhKwEf6QZ/qvW9bdadoFT3T4FzGrjlBGmzFnITsh91K
APmnjzhmZKoIvMEB7N/nfhJKwd0PVBW+E45ddwGwfyYBEz4zEzsw42ccMCjy+9ht
qCm9ecgD3ub/4tAjK4ulrkxB9NN0rJL8hD6bMAsUQQr1wz1t2RjKc82W3P3O1loD
Ts+9PLhHu/qE1vzWPgqv83TTd1C3eC9PgySsgnPzsQy8/m+GEQ3Sc6vbvizWjY2I
iPsLxnSsKB+K+Jd85bsPPcdoIMHiVpDmhsZunXRNMUm1zCKXkUvQ5bo960LtW25j
Au4ypMFzNfMSW3yF/gpsjULmmxoGpUgWQaTxJw23vjLEdBJBLR4BXBbmnh9KW0gv
v9Knty1DicM3XaBkG1c3FiD4d2lzB5V6vDPmgGhGqI/U4uMaAQaIfy02m/wfDZrK
Ma7Xj7ziLT6axutLiG3a/eSuleTZoTlnBaMxnHW/8c7AGq+ADgHEwgQ0Q9MCKWh6
4/8iKcQBxDpXAuyBn79Sa+LzZ4M0jeG56lN5baExVVo5wIz1eGrdpKTX6EcYgFcZ
Rpi5E8WxazuDtDd28qeO5uhBkPZh3c4vhMILT4FcpPi83Ti3eq1spzPszSPlCrhz
djwwfl8qwP05T/YJVgLRtqzP2SPWbXMUtBuoLFYS1NK3AK3xkR7hd8v1xx0jqW+6
7Jrq0gh9r9dcBAtOndS7lx7B8F3ZzJaLNtC72zrdT4DiBOkkqn8DTDFnaOBkMHwC
8ptGQFJ1q4j0Td67A2Yupg46bHKgDbPwZYmDTaShZff6IqzFJOTUS7dBxcCqvnVJ
OV7b40Nsj9eWBjFbAU7U8PM6nfGIlGYWpzSqNmNxaVFLqIMOE3NxVZuwg3b1Yn8I
V0qBUGJiMae8/Kto8XhggrSeDjEaTG8hm5rvszhSDD741KtVRPXrd8+6+k9sEbN+
uKHZxubzICng0ifc+jS9cOMUXUJy5ImgYI/A05aC/6fo0aTy4KafyeJQvXXyBu4x
8LyC4iueZjY0Z9WqLQc/SOn1cktPLmiHxNYrcQ00pPuC1ezT7ZLBWDVMjFGE9PXF
w2pao0pWykUfv4x5NMv+KYKxOvRNfUT1I++bpZgJfbV5YhBGDCw2ieN0+FCqvx51
ZxfxhJq3BKvw3D6eJJBw45qy8YwMT7ocavOTFDVuuM4XTLHFQnDMtfD5rI8cwjCC
NMO+V7ROMJmLoTqnAM+vJh+I1eE3XWuDsG+gXAPjuUzyBdT9epSNbC37nQA1jLQT
lbCmnH59DgZy+uEIqDj1hgmBhVZGQcZ/cLG7ifUziNatoUoDlPZaflmoe9Urgi4D
48UmVXB1MHdPBbnWv8s38JdZngA9apJXfkdDg9JKXNvXw4PANzPVIWp7JwmU4HnA
1JqxT7waS12zFfiaa3/5MuLJXanr5lZa8Ht87LtHCHgY59KUqOOEAm4e5FpLQl6j
1y4jBLSj2iehgTEtPQGU2c72duGT1g0EVX/FLP4ZKDAG9zsR1Etm1SNDZMIPQlbg
chOvs4v7JrHoZ3l/TjcR3JKQYjOD+Tk9n9A6UDxWCsOElHvI4lEkYk+Zbe/QMJgy
8DIfcpqHpg+cHT7H+tpWz1ApPWxp+FfvnJOxr0nKba6+QH1joShlo3l+6poQYlIh
WduKvt4QAqrlepCp2OAA2VvGZ40fo/GuCS8q+dX5WoRiMRxFH/fZN73K4yT4nPuZ
4JVqpOwr8WSc4ubW4Sog6fvMetXJykigA5gcB4n/nY5Jy6L7cKhP8nQZZqWrqkfB
osniNmcM+QHnT94NRMf2JVd3X1vmDmMP/MVYMOg1ds7/guzuropekBh+YZkKUBM7
cYbbqViYOOxUtNMCyrdn2ZxwtkeTHKA07J5MLIFrONU3wW2pWndVcvZsbW85weHR
UVSITbI+BMqAhRcU6vJCHhiWQ2KyYKPw3z81K5Vwk/yLIZQ8iOi6PHukScjJh9tl
oJmKEGCvjRwPsFR3OX4n02mIUXSnUFpyJRH5XpXQmj/bsfY3dvXj0rd+q00w4ejZ
ba8kqSkn/bhBgQrZy/NshqrAS67vLnKHD/U0pMDfVOt25Wt001dj2AKE2b0FiNDO
3Y6n6KoQftDnTfmoMf+f+/KkPbFIrWT1+RntvAwmvCGVWf5qGINxAYTxEzDog7Y5
4AXgioKvGMMvSFpflVBTbuaCwv3nwxgVEC0o5hDTkfKZ5T3+1GyoC7LJSSV0TcMS
TURFuHLuIQ5NePQxD5JG/Shu8Fb1yfYeraiQG6O69gAHuKkeZ1aQ1zJbrTBNFZid
BKIKC7/G5BPkLNHmSxfRtBEIecRlEda4ZtNRrxWTX4S8b0un1C88Q6cmF6nmP2uu
6cNefLt6JNTK652fBX+5bVKcJwVNCpMH+DZn7fy6yrDXzogC2PCFdwOpQ2/VrVuK
ZdmSg69YGA41zcMntI4BjPkL+dOt7rzyYRGnmIRuXPEuxlMAA1v3GYy02C0ICT2W
Wugcd7gEWwEpIP8chHg08gDJ/BjaoMHqnty2i7j28ZDxSOaqMNcWMo4hIRr4gnR2
QPpMf/iVzdS45kGZHV+dfAH+ZvfEH/G/14qqnbz8CHY/8hk3myjk1TQEzBzmipsU
FWvWYC0vjVpsHVEqhmxFLQi+7ljeUbiFsiTF/OolmxLHl6rpXq8EdWUOUN/W8Ojo
Cbr64Ce2ub5oPOBVOltIokYjpPVocwihN9FLKE2oiEiwV0PnR2tvcIr/DTqcLHZG
XdwGLwMdtzE31BdibJyT0Nmm1AenThdWe1inJzdlEecjhmaf0zNHhz8WhLg/+2RJ
kcTvBWtMfRZVVJSuPpoKFQSmT96elPC2EIRxXe88cb9d0X2h+db3edtWOHqBiLnm
SMt91paBWawFhJx5u+dord3cWt0h06JecTuTp9O5xWNkq0jCZJJlFdixdu9rVX4V
XFQZA47cOYmrIPNNvvXzvuQ4oz9V+sXFK2cswkF/pMDh8IzzcjMMnT1Ka5dJBK1b
m2bzkLRTZ5B9FaqN1tol6ulR99rEWJnmYKgelkjk2WZaVGWCIVhaNYOoOCazfuYb
95CK5/ETy8uvdEtwOqZiiIzguFlOUX8cHixu8luITRlXHXme9+ETO28IAxFlexpJ
QwPJhbcagW0ECvYyNVOez2FmOG51MUNVh98bRORG297OYUZW4lJne3nVMD/KAZ/J
bQ4guTYI4LF4O67UbGBNlZiQok/vgyYRK4NtBDYBf+YLDrwuMu0pJr3vpC02hoV8
WEGfThw+F18MqhO7nkYj5lMuUGMYG50ievwHHrgdzpBcpm0H6uLfr3boUskRIkuB
l5Yo7gOHYwRp4SeCTWUIXKJNlPfG7ND49uAsVRYPwkLRv3agmLPb8FLtDJAbQqTH
P6Z9K4ebMoROLI/5DzNbjZ9TL6jlJuwRGGSxZoyn0E09l9EuLBbClirFqrteaUlY
rTfpNu6IKA0sGB15z+JnA/M/+2hLoY2igpRfn9BeEj28c2B75sw+BuMTe3z3Sp3Q
BZmNYthkvq7PwA01rRyArLFs2Vauk8Nw2zYwPbuaGrCPz+nJRRaSJAaiKmFTxBi1
hWImc/nPCHD6WMPg8M0WIXf92Joe8n0iFwkZ5AEKIRXDJhHn6sUxmUQs5+qjCd3c
UC0PkL0InB8ySNiG82MFy4HEf9gBUgPGUIJeQEHdgGU3IsyB8lcVuKV1stl8glom
VM7qZ9abAs7a4wFf/nmNQs2Gg4QK/7SwOO4yOFwzDQ+1lNr9bjNHd7lbMr0uaMQG
htk8O9SbWL6e+DFsdoeX1o15r7gaqQdwtHkoTviAR++FWZGr2DITlgv/tjAGr32V
NPthEzXxJ31jhg0wwhbP2kegPe5y9/j0s7PYVhsKkGZM9ja2IWw6Fh7OnlexOR/e
NIGQACyIm/EB+M0qmQAxVVdXravi4jPlEOwaCZ8wlgCehIRPNZt0yXu1xJtUgtFh
2RN1h0vnIm5RUHGfC/VeR8a92EsEfaKtQmU7HDs3sflqp2RC7epvVJsmEqdcjlsV
uJvr86X440nVHGlENSubsolCJ4iRP7etiVT/1Cj3CLhCN4FETbHhjZTMr+FnWPcE
h7HseAGpihRL2PKD6wZsH86AWXF5QvCfpiBZKDoWEBoj6NZ0dynx5ZIERmUjmTst
GC4g/ktAFXrjOQ5ApUP6Bn1VaEgeYABGvTBuf7REPyMCKg8pVLyUw37sD47AdiJ+
BAKo41HDXzWXPFfrQHLY5mRqYZFrjgrqW7szLOLn4HvxakijT1tmvinrEY8uFhpO
9VABsYyDfErdEGVl43O+fnSdOqCVna5rlGm9fPBxA55gokaPJbTOUBM81i2GrAKG
IaUPDRSTMc21EpOO4g99VJmyC/Y5qw+k/F5MyGVU8rUAVgTwaZdepICPAZOtawXk
oVnH4iNpIDh1VRxzG/rLxkI2t1gcuf0vxxm7Lbqcc/8hGZLrCRRpGlFD0bvcv4ST
wYoAwxynMrtOiuWa8+Tl2b//HzOUpb9X69NfjG4EovRGkxCM113W88hebhsUZjw9
B7DRi/ywnr7YJdS2XH9t1Qe92z4F1M03fwmT1SS2STWm3OL6ul4EpjyESbPiio1j
J4Z2k7BlagTHhZd4av8aK5MZwrEQGRiIPsLUzkuuAOjNoVkRb5bLiRhaCl6LcIDA
yALtrwdLLpEErkOpxS0fS0JtGIJwNukf7KAL/+gwAoOlgUYG+sF+GpK0mD1Qt0Y8
ddwD0GDfJUKaJjHIgWuC1mDUOGkUxnv9zixO0CA9A1OJTTJmEIAH4wcF4wjb0lMg
I03e+RL/xo8UTHUZj8OlGaR/a3F8LNvL+7w2uEgB9qomNRfm4uen0px2/nB9mFtP
GhPpYi5hBmH9P7Rjg5e2b6jhUXcgI18OTpFMkAUVC1v+1wN88CC0l/dgN04F9Whc
QVBIjdSfP92B5I+z/Iv48xVNR2r4h5+8zVDoFCgsoGgjeGnjB+hhU/38xT0hH/DL
zlHhoYM77+KJdTu6Jldqm3kuqNo0XaxZ/EacnEAyRuYwpLa0nvL8Y67W7JkDWK1F
n94cUiTYet/kyL6o3Oc8926IP7bhh2tJSkiYHF0mSaXdzgoI+MxuFo0+R8CUanY5
ULNOeCZwZ+j+9VHL+OjHI9DvC8W/GbhzRuiXqMMr1BVPGSQ7dia3qJJxvzkW/1m/
kAlP+bZLBhRbc3+0a5uwtvynAZriLeMqQ4yrgc9wn+ywd1ww0YXBorQUlgmm0C9G
cQ52bSIMh+Sthre024obcpXKVpRZBGvu21ejqifI4Izn0Ck1pNTD+MbGTZQs1IAq
zo2TWFot7SnJHRW1mZ3Lo7PKIBBONZamygzetcqFQQ74w4e+GlgH8f0seStQcpF0
M+w4V3hQJBl3hlzvJL7Z5eJsFbA7nABB54ZRbWE3ImaPshMGy0bRgS3lv2EmBuf0
ko6trBV5oLpHn7LHcoc9CLrVO4CcqSNA6Y4q7YAt7WD4CM/2jhCShvQytxHMdxXw
YcjBEpJRVp8PUaVEXrLEtFr9bp1fkAHTlDryLlqyKqo1lGmIo1FfkStbwafodO5g
nBBLnrlawdl2U5XQhfHf8N+eQeKtlERaL3ooYvwDF4u0WMlLrJinKQMeoV5SXIad
848dM66h4xsqgsvHrVthLH0VyWNcY+iB8vjPlTLgtj1A/Q7WZGRDRQKACma75U5C
kh6Dwvj2mUe8NJiLB9L1xpuwow5GV0O9Nh/sRoHJ9JidS0aukYDHDQ0O/6pPDuUy
rMpjwQ92eQgCZCjIRxhvXtLQhD/TsRVbJWoiTqmyus677fDwne67NuupB7JItgjE
o98aK481EhQMRXGc04aWkEEGpeLtzi4ZM8mHtX8oXCRbUqZqS00KNhp8/xtqU4Ka
WjTrqJj0wTz2TmeloinnHCMll53fHHthCC3GckKkvQTTFDIA/m3DkfbRKcSJXhpd
035A7uqtfYrai4RlGE2nVUgcr1wtECm+K9uMODCRJNA+yZQp246xALWGH9ZFVTsh
a7+Xi539bBOaS9aokj69n3ymb/4xUsTmnsLJxDZp7EDcuWJkWPNsgtj3qVN8XZPE
u9+/ox1HH3hs2jlKyL+9jRVJecsHhahaDMYoRed2cwt+PjoSCEcMu9wKM0x4YCkD
2NDoq0uIja9xtbtO/wINiV+G52S5LHRqJHI9he33PrKWUTo786GTwxbA9rdDsjL2
56kjphorNgYUg4xpY8+nv1OQnDny+cDkM94nAAdWlEPLhuIoEgbfzZpEnUvdS+yo
0gbzJpLKJnoX1VbD0dfeviDVn4yiKWpY6VICMud7XEPwYBqar79tZg2Y0/Kqpk0Q
I/7gAJep6YTaltDWzJ7SkBVRWVBh2mchiK+LXxyfwqkzazonEq7WvSZHpEH6hDnX
fqcheDnPKTWTnDkvXyqHce7eDgHXaAo7WvO3Jn7tUeIgEyv9W7qmxbVhB8m5yVeL
sVd0T+tXX0sC6jeRtAUyxdrmR+0Us/pazhGx+T8bL5kVJC0gFIhUeYvHO37BjQDK
M7Nbjq9CSz2Hi8amAgFKKuuOFxFKIHQz4h+0HQTfCTWFX8RHTtRBT9CqV8TkfIuo
/b7xNv3ldmRc9EE92KyUKhdMhOhYRvcRK8+UQJdiixo5fW3d6qYLoSDO487f5Hi+
ua2j2u4IrRiIpAuXBzWCZ6q5tyS+/XETA9rPqoAaRoVoAxL5DgWd3/+MxTSIG0UJ
P3uXEXioEOan00/8FeSJujpU1Q6bqeQHZpEqFXY3REe1Q66rMmHcIY97P84fyKV9
L31BwcQhNsXFGu3ZR6MGxQgHkmgVV1TbNiZP+ifC1ynReKF9tPzUbtHmrzsqYRkf
AckW8tnZHi/baSrIuoYC3dPvENwo0kYs5Vh+QJe3LSuMcmAgAP7HD6NAykfKzjiQ
AydOD7l1F+l3CSbNXn4WDVLeHCuxwNFy2twu0TEa5Z2I0+uJHGVMY7f1tRPZZuKj
hFVMGAUQ2Jftom75RjegGYVbomCB2jEnusSacudDh0zDclHE89QpeSq5uEFWZavN
THManeNFyWCiQMbPRzN2gHhNatQqJUOepLDjtB07xyWUhb+N8QvepAtoOPPf8mKh
H4Ys6mzymIVUpYyG1ZF1+fUKFLeToxMLG1eZNQOeeEnTaNr7bXnCb39o5q2rglJw
V/BfWsxNwp1sffItJ2yO0SuwvakIiNZgyUsS0EWA6JeARburOr7InNJ/Ncau8U2W
mqSYREaxZn59WjA4BB45BZNpQiJdVVDz5mOMfs+pYFV0hVFDkbkTekYea1eadQIJ
9ZfN9Gxu1jTngMvFhQ6K8DKM7uXmXZa1WGNEc98kMoR1SEBAzlosDIclkPZFbuo8
lWgOb0sFng7hT4Cvz3UZHsE5Ze2S9qSeqyYh+ANJGv5rIHh9ll7vO5J+dQjrgEcb
pgkWkfL3YqhwTkKHIpLOeXZlMfh/FALaWSpvPcM5pKfThITILUIZiK9NVddqvS5y
RqaewgvENEcIW+GjTMYnMqo1B2IKheMgVM9bd/LLHyBD3i8wf7w2LNioAQZx8l5B
Yon/aHjygm8KEy8QeUEJ0py8NsOC3UZAsh+Ci4zSpD8Q4RPifoo3duy2VBcJ+g7D
oFZOk+wm82flOUkfEiSTC+i3IPUEhFJUxjDhrVg65NNt4jPFcsgD8PKEXsSIKzUe
tNrRgXn0P7NKQHcV5enVAWeOlzCCHce41CsDHi7CeqV14oB4tOQkSRJnQjBO8NlU
WMjB74efiy2YPbafTPIYYfk0enISF9hstBV9DL60pvzkj5Hpbo+pekv3/oxsOP2Y
sspEWJJAgvE0U0OhEsyNSjKVh72ovhd+KuFt2m6LiAWKdPx7Lg4LnaUScbfpGueF
MH90fzHXusMJMzzVGg94h14kL0QaY2cHuhehdzJHs24Z+rRIqQhItVCC8nG8P+oq
zHzmJj9Fc/Y/NMJprZc0JMr2yU+Gb4E/rDUNBASBR7bICiRmr4SoqrocRAv7+9MR
9Jhef/1dW36VHh7CAVl0Ur1fHTLmzVbKlfoTgJCOeByLhYXlqN5btvjlg7bKAVCf
uYhmrhlJXfFzdxeqDkJASz5q/wna99gqsEuZ8ZuLVilRWOkYZ1SRcylC0EJTBxzA
R4IIdizl1iWxfPJ07sxkQkR8ZJ6UKBHpKca7OfIxM5bqPoqxiNVRrr0G539v3Iw5
ZGofI7bDQ/oWOrrBVL04zVI18f+k7NLSX+WT/Ze0f4vVZmGyC3q1hmQQvm6GkqKR
+bjOwS9PGL/QeLP+/+NbeXnwU78hKcgVhCWt0qL3y9p88D4EXTOkPu9l/YeogncE
Mt/57qhEjiOKLGfd1fDixcITake2gf3eZ1+5u9/4XvmDYRyABy/0JUx+QySqWvV0
T58RC+u7GZEAPmiykSPmQOYxAIy/lqVb05c0vzj7zCzYGrGKPqYnJVkoc9K5DtmZ
Sj01UneDqgNE19GqTe+za7MowEXgPIaU7AAClI4z+MNEy8u3DsQ8o8xGprwyzrHx
5Sx/4+5pMljIT9ZIUZ1kYNGFR0PWHNm7SXr/4BEZVXpdPKAlNTwiWA8GoQ3a0Y9p
lmfMvYytpONQR92IqFoirUktdj6+eYP9p4/t6o7XlLyjhGculS7eaR6MeqZZcDi7
3SBQbN38fBZoRwTSerhcLsNy1cdHDLLOmQLb7swm33JTVwRF7w41pCBsCIZBWNUd
d8EJVPDebXzQgncxRSzE4Umy6sJ8MwrLoszade2i/h5d7D2BqxEMpC0c4YBKQHA0
QYKCs387ZJwd586JyTESV8aJ4b01rXEiJxt1qJSCKACFcPPgFzCfnmzKAB4wTSV/
UgaRu7mDLdi1NlxNeXQA5A5CxGlAzwUiLBNf7wFJmvhpIbnLHJAe1tmSAL5C9M2F
o9ByFc0Qikiumb6J96xyJHFWRMmYVT0DRWbIeRvRX+gzbQph4GGzPzU0IV5STgvh
ckVkQN4PMNPOp1Ba8seqGhZcfcJvviwiHM5p4I8Od0TRwOvbPiYdbN0hm9ESVUDx
nV7pFmDXXigRBuTvAGxN0xZ+cqHcJrPDGNOQn86KwWvSJSOkEeUew7B1yE/R8jRt
RTnZ0ee+gvF4paV+7rPExbcC6hF0WrY3VB5XBeXeXPhCv9SxFVdbrtqnXV+8XHRs
PbmHIsJ7Y2RZzliMbvhjwLcGqNAxkiiU+xnLpdfvjVAIfOXJD2EVcvN/h7Qes9Hx
DDcYQeN04pZ2UeTuYPyhT74MALSK1Q1JNyPRgvPxXrBOSozdLNqur1yXnXzK3eaY
FM8l7EKUJAqd3XxGz7SpfB0577Gj9bYyIuPGQHYQqim3IBfYRZkejQDzsuPL4fuV
2s3+ulyNFuqD4YAAm1blgLZ/zTlqIu5GRsPXq5xesbCJviN7lzQVTimYxscaC/nE
6G0PY51z4E1Qco9Plrb/M1lxjxpC66Vp1BWmmU4d3fhEquZfnUCYlhr3wXytGiiY
5s1LOpKa1VV4Y9H2E7v3jBdh4Pl/LOuDZdPP+IvsClKdo1CA8SXA0lCTiVvXfFaf
JsGrvv+8Z0IbmlHFzLGvW42OpiFgPCqeqSq0+QqeZgy55OAEqm2ekdc/Ly8CLzpe
TwwD1meHBArXNadG/NJps8cBCtviAs39BAHDzh5frO+EYIB6C6WML3kDkbPJabHB
TlMlBZm32Dly3PhcwQRa4ZhVMTbKjUSSlaCaa3BMc6c0Uq/yjBmb02mAW0d/UF5l
47zJn3x47C7qfXh29C8FLLRLX3apJ7eqQRrPdfdC3jykbE5V10eBcKAkJOvhFL8K
mZKI/B/i5u1U7eEx2M84sy4s+4fto6UMUnFzAhh4Gofa7zh9bRxX/IGAK2WYWSt2
llmTdJEHdBmBpGt0VUK6DPT7YVnq9Hz6tlc3ZJR7DamcgyMQ11ynmCy0ZaBEXTaQ
vpQpTsECO6RIRrY/+qx03sprPibh2N8NNhxmOYp6ZqpxzXvPud9bkAYrO6HvY+2L
xIcqhbqrxymBJdKzZ7hbr9aZaYTFZ+45hNWtccjEzdioL/MhEI9Qn7tOe6Z1QqHh
21bcUpgB5ebko6OoxazeKlJNGfY8u6ISTsKCFYVy3hIz2/yZ9Ti2YxpiqFP0gEDL
cFEeyN1uMjTfKgjCL8iCkGtlIBaQad40+jiumYgBnw2W7GguqTVAThBGGwoKAMDs
UZPrhi5DXGFpNReDHPj3796iYUCruh+6pAYRmgsTIn1XrMm5q9UpGMzhIquMON/F
+DaSQ8MsKESiDayaWqNMDw6mHolYmiq8ZlEwqIJK8qQEm1eTy+OHi4ETJYFMb/Gm
AF5+jEHvG3SdQS+JFwiZ4uSw7+jzpwYKB9kSKgkw6XFseGpjh7w9TNb2cmNAMvTy
2Ts/xhyXir5ZokT/DyQvxjOIiHfblq1PC8vWujCeWU0JerwsmoLLXxD00OCdfb11
Jq7nb6yqNSuY3pXMJ8k5R6ARXEzSiLhEZ4wxL0bMVOvVRWRNyvM/NJ0pu/H4qIz+
aM567dMr/f0O7JD9TNKtS3wJmX9CpldWBcvs9rHv54Ndv71R+gB0jT6WNynRx8DG
OIaET8Wu/gk2J4tJghE5rjEICRKrYo3y65X3thgGhEvNVukEtDGD7/4BlQb1mvt8
PYm+OInY8zeofCRAhs1beyJWLI3RFUf+eXvkcO6+PB1okVSRgeaBQud5eGf0i0TW
N4ZOeFDvONMLbRUP4QQylduwexK/teOk4oO/5FmuDPTGgwFEA3WXeOKUL5djCs4U
Z6Dp5OFnrulT3NosndScRoJq7F6/3m0A9nqV8b3HsnTjEHYZsFLqFsQO8L5bPcJm
hkClA1I2si5mIsbnd2ZafrkM1Cu2YfKTxrKlJgatE6ZcOlTrrrzOBhzf683ZTeLY
jUyuJJh3GOKJew2AmoH9L8hDlY2TWbxCXqOdf6F3KjJo2wwFIkRcG7DgebTerOvH
1ojp6g1ij3ysX784kX42McYcrCW97BNRxWH64VYgk7YfMqOoTBgZ1tqQIMAPW8m1
/rodB3CtSXUZY0eKY6g2Nbl4CxMcn+5BJcl2jMiFEjNDkGm40+CLAJqjNwsdpik7
VoUYjui5/vnoZHLsErqzaudJDKqOj6eb6NHiU5FswIwKXQTTnMKAPnW0+BhpvrlG
5PoGakHo2bW6pJYMRNOePozWnP8E/WYaSczYXa/qZ1KnCOoE7MxFUa3s3LuwHuef
wIi+/lQ0Y1bFazHJncashTN/zL9bpdLyoqRp4EvDY+LyT/yAYWiN/3uSKFcFJ6Qg
PpGvhnlvVjqSSPJCjygyeNjNbY6NGIHGSCZM8B2R2fMySQs/NO63aTTHS8lAW5Gi
/vY0CgZGLi/FmPULHgl9NBOnYwNTxCMdVcEEVKF1gOMmdG66CDmp5DOF+bXKo+Nv
442VPodySzeBq0g4g+bu3dWHpx7oWBy9QQGDqbqXs2i8hF1dL65TN/1n2VvzIxKN
VzeYn4pRwvPWkcwXw7FLJofVuwCXCnKZ6L9ryPLUXRu9OCn1kKqJ8CbUxRfoqXfH
Z36ZlCYOav0yjaKX3rdInjhAU2U7EqWbKW0EFvwZgjpYcc0OX2Yjx0UzfGvbZ+ZF
Jp1piMN1pCWWmvWCVj6eukqcGv1eUViIXX8H11PNmcYvjFjWGSt3Nrpb5i+tViR+
FYHVl0xGFY8oh/gU+A1raVl6rn8bvyGwcAZ6Z/p/elzcHhAOJXI3YYGnpW7sNXXi
r8qsICuDdMEDGZQHV4K4Hjx4eczcODl5oyh73aAYV+yAHDXpXe0D/6a8cGCS0u5F
bFyoWj9Id1LUlFkEGmLG00VTjwmkBhgaGPp4wrEjh8VtYBuyx9pyIiIGVNAa0vtI
b9lC9IVIv6fPwuxaFmx8YZdL3cPriXB44p8WfM2e1bXmujJD30gOAdDX21Ijiplw
j2Vzy6hLv5CPzxoTjN6giIwK8uXtNO1uDvTK+/ynsqOZjzUWuUF00EesbqEDLvQG
n8ShxjDpFREYRrCZ1sPgkxJR/OmDZHasgPUtEsefuRJwkb7h+4tWBFFDOvpJEi6j
hHuuWghmb5ue3VxCmjhDjP1K98Zx9w19pETv/PuCOHa674cQ5Ssj6KgmI/p+znXP
Pw89a/jxbNyuZ82Jr6j3aZpNNY2iUxTVK7NJmacsupJZ2LcQ/bI8s6drdyiBNqVX
m4OUzwnsosU+8sn9jzFi8xnLhRplAGZvvDtOhyUGLEuUKXLLKgZVvSPX5W5w9QvX
6fzj8HfjRXQLygRpv1ymzRdsZPQwG0PM2eN1EWI1vbczL9CkdtKkdrO5n2NGcz1y
HiAXhDCwUBsmw1C4LmqEVPAJLt6yRyGdThelESaimDhJPbVe90BoPac4Ib5ZvtEj
i6zrSGCiaB+m8mqeQEzfOx/K2kcurcJG8nCMutkjvnThOsl6s3MkAjxyhQDxvEft
5w79KDrGRrlmY5STm5SJbEzjm8DUiv89N7yk4beoMvedqRx6NOnOmyA/34XdU7ju
kw3aA2oTXkvqgIhH/a51Sd4TSZgrtaVX1izLwa+oAJ+h2ZshC7NHzr2kzr6OWaXc
aOJtQIn5uXnN9AeWjdbb1gpZ7pLk4D2WF6S3ld2L4kPYJSY1gNxdXfivcFHiZ9ey
uFVUxEUmdg5ADdqs2zVIevysja1YIQW4HvBLHkZ7jEl9DY/5Aco+RRZx79CaGg0C
jf2yL9DMdOzXimyTsp8GBEvC7XIxpYiRSRNFPp5MMq+5zO6gqb0BNyqjH+CyFYIN
abI/kmXYjSQTFqpOJimoacN1pG9zp+n2RkKPJhEDquWSkd7zvHEZlb1li0pBNFMj
zdnB5qxIDhOzo71869oFskv9yqobV+umpxQpIXZDFjTIC1jyzp9P/1EQtMJ0LVnI
04OTco0+UVSK0B/+SxV2cS3mpA+M/UGOzSqmtAEyF6uZYZr0WyOF/ut7Y20vxNjw
+PJVlQEEW8VoW3gB0S26Tj5IWJJ36Cdvx1bbxr8cxQHyupyPootvwCV6M1V3AKM1
qdSjm4liLp9iA2YmmCy3+Ra8PxwPaYMgcKZQ+p8COPba1VnuQMvpcyAGaqFg+xoc
8uy0qycG+NABRjUC0l2j1Yu77t4cgcQndcu6qewH62KmiomvpWaFaROGJWvj8BH/
wu5hZFGTxRI28gRnKI3b6TSVUO+xnEYr4UWYeqvgmblGKUv893+5fggFV8gcyj1/
Afm/Qdiw/JGVMoOSP6e7VCSX6FvlNWeW/uBj0PBIJvQiohXCiYuGqlMI6fXqntXG
XKetJas1Pjv7nEBCmWfvM7Zw7f78/SMgGIXFN8/Zt7L9tlQpKQAYidQAvWdPucxP
pFkc6Gig3SM9lo4nSq6acxJJAAMLN9KDplqbUfgzQXc+uabCRwgKS66ALcYldGap
dq0SsWv79xACelTgOpZLhNhW1WyBQuXWKnPUoIpIrNudPnWi5/jB5Eji8re8KXPk
MHjvCgW920b4Ss6gqR32sk44oXFWKzohg43JCpvaJTT7Btdb9VfFbJOycKjPRp1C
zeIUn9S+15jgYjAxTavPmi4l2Ggt7ee80hhk0Qj3CtcmtDHVq9A6362zwn1kTZ+X
53tqJcLt7+Romvcctxqp0dOXDWXH4GdalREmpRiOLcyfQzMM+4EExwlQ678TngOK
q0OYfw8TJVwokqmXTu/x/i0XjX6VseOJNDWFyoydpS52cmlXbM0uI2Q1jr8Eos9U
kdxH+6WBYLw8lHxjTnPFjkg/9s/FyJpK7eKJi/j/QLekd2ChDj8EEkRIkzpAsZVf
jy+Lhcq86VUPXd/KPHVKgyFfv9YWADehEcIW5km0nZT1PRGw5eC0DEeKdD4ZNux8
c30LnEqffkVlDXYs0Na5oUKL2/S0AIAUVb6QzougpNA=

`pragma protect end_protected
