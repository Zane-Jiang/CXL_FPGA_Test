// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
T6UqAyN0Lcq3GageJ1MUJU/HCfQWoTski18sNvWh/9DzFFU2646zXd7rm8M5
mmuYl6Q+Py7961x5jeVujAhn9AqvP95rtu19Y8KVS7quWqJSpHJX9Z59RTSA
tvO/4QH6/wR5dNJjetvjiC+/5aCZCw072eWTCwI9cjA4fMSdbUawxoYY79wB
VVw0Uk8oQ1ufN8itbOF0bPL9+qkmgDEPe8l/uk11taVcwc8yxktiPfBczaKE
4asm8pl9oBZZ1oaEN/+j+Aw0mjkaSvRjiDNTlBvcWWGQmtL2holpQION/D1u
QxN6KJLx8Bez6qpJJ8wxxkH9tva7leqkq7Cd4+bqWw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d3L0n2eLfoKlg4q7r8WSULZIazit9+QLIsfvXf/mLtDHb63H46rCTl+c6Ny0
ctJ+J1zzCAqw2zan/GUrVO+r1C6w9WucFH2AqBV3ekgV2uXm9NDK13Vyp7V9
pXxVL48NLrmiJPuD3gsQh7KMhuEpNQH4/9h7vBpSqpsGDBy/t+7hknbHlSRY
1iKcNYxqvs3B1WkNzh0PaJZWc3Hfg8OyyutSqwAJm7Hory8VEmyf9t+/sMpA
hAs4956AteynYWwHPE+UbNmVpdxLlonYVuTQfqCdGGRRplc8ApMtW3/Po0Az
hccIjZbH6BP/QWG0swVOkZjPXO4j46CEqtg8s6P9ig==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fb139INhpZdDFCnZ14fj5TsC0O45MsH+3Rm4AaItd0XRoDdct9wQURQ3Hy9c
k/SIdn2TAgM5Yb7zEqFyAVqiJamv9ZVRG0DB40b/NK0EQMTv2n2Z8ZcsC9H/
HcVhJfrv4bOvZW8+qaIBY2txpSa1uHdgpI6DjK4UlQRgOaBlAhcPPREnjM9M
Ec7Cloy0Ku9CVVx/LItEuxHzN/tnb+H2FwO7fV3TsTn53ULfk70r36LuE6iv
i2FwoPhgAdbFmbEh20N+AqvRia5LIDpWtEcTjcy2tuXXeUkU0desMGMyVF9Y
rZ/kcjqDDO2CMRWHT+F24bGioZx7/V7Dnp8ihQdaag==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Wd4E3Zorwx59iejauiDkKyfct/lZD4dOWdOv4Vuu64cHoPvGa+RCph1O3YhO
lx0ElDPE0eM6tdQjPSXcBCntyoWUjGGG/HDUvL9m925n5WyC9TT2gvIELIOi
fgDeDrxgc7iJbpCrdULTuyvmlENDDIvcOdaYAXmaFANg92CJ6vU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
M4Kk6x8cCJN3EZv+8IsL6728IDzS2SBYTbS/xoXOta/eGbCLXLhunokJr043
xlIU+OPxsfeTbtM1L40IEtdkeHo7F/05NExz1HRdMB0KMuAISuvqAJhC2ugj
fa9Nl/pf4qj7xxf29/Xpsqejqat6R7SMvgbmXRjZhox1YNL4FdSI/QaTf5Tj
mvFNOzj+Rs2t0qj4hnwrRnPDWrcK+ArX98l1D1pmstdTrnSJSphPTSoCvpsK
batLPAtUv3jaMMYoHkqXk2/E8nqYcNoBsXJRP5vgUjr5r4NQGcH/gxkvPttM
bJQPPFwAKq5ncHSN9/cjfP882stZrUKG0ftp2B91JkcADOqwrHEQPrvDMKEr
n7Fn3/cqwIt3Wo5xY0nWoX2FcL1Yx4HOv8kcwz6/ioyu+k7+rIBFf6iOPoP/
E3fZwpBMLzG/gwDnG3v3ieAjaymyx2Mf1CE80WT3cAvphYi6G83v4hrWwz2Q
bn3IA3b9jpAloPl17n/LiNrviHd2YKDu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kYt3gN4/+EltJGjndUmwmmAUfqamH6SDUDDT3FjcGRCk+0quH/nAl/v1Q43y
iLnbQLoaa7zO1TBtiq6LLlugzq917pSFDO7czENorbkpNr1LoWRSUoScKoLx
yATkCKAmiYfDO8tucKVDewt5nXV8u5396LNSdXqKvEDIZpB0m0U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IyF7km/3ROqEA99oQkVHwlheejuQmGA24yd+Gc2lvJ+DpataDO1xZq50I2Xd
bMLQ6JB7UjIYgpT/baY6hV4ASv7xTqK4AE6ROqhGUXRCK6Ac6dTC+WZCOzkS
SiJhCc9Niv68ShFgyuGj4KVt/5vdyQ9xixjRCNA3WBqXzub7Xkc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16704)
`pragma protect data_block
l5/t9FfC0qk6U+FuvT1ATOCZkY9rCHWr2BzQrk/ALUziL12aWT9idDtvDpQr
5I9IiL/jJAJ36iCPGUkTTJoFPpJHJlvL+eUILh+wXK67EdnmHFaGNO0FQDAD
C3vbCiJOzZUXhRvoHXJeYKTk8LC4svkExV9pAeYLfJOyIe9hnKER5/FuRPHn
5P8BjiJ6ypvBPUFCIeErYtcKugmF1UmxWIJ5GaLytYpr+lT7HqvMxAvu/247
KbCduGlttyIYPdbhoD7pXtEa9llX8MSPA5njGOMgTu5Ti4BVbql/vWjkixUa
b2vt42efytB5xntZ08oMfskYRxGNvowdAjYi2YOX8ctntUkmngRXp8g6xAiG
lckEf8G/vG935cieV5/rARWXkIopIuohfdFTLvKVomeViP1OcQ04vXUFuw//
WGwJeW8AGddeath0G89Q4bWsGytnXywT28r2t6LweaI2VRXeB8L6qDWYDLhc
H9N6x0rf39+DJ4+GteDgiikF3yKRXjt4xbDzPVY0UZbG5ZL0GYgVZ/f31vOo
w/g50L/7tQmqSzro1UVmqLjXcyr0Hm3qW2CiONBIh8qoekfqGIM7+kwwn7cq
oFP4RnTtcAsvgvTcfkdTd5uOnDAdaLVlRNFt/UgIELx0D99uxLIRPx5fEvuM
Bkw/RNXtHzeG71BRIfsy5t6gWTo6CK+L9nB8pt2fOhSAU1IODayUD43pk0um
L/AtkT2j2Ww/P0dRqLo9Lrb251Ec+Q9sYWxwRHB00I5HDy4zGfXM2roxF2sU
Y0QypaLn4585obRmNwXuB7pwI5eNYZAZRNBKDJcv1mMiEMnRI8ANm1BiCTkm
THBNPNqiDlvXlPlH+sRvy03aiVs2XP8kyM9gLNkSA7T5RVJbWUdqleFeVOsW
gpNss9bUQryHfRLHOhZx0kIW+EkZQr7zXhu7sB/3wUzt6F4h7NmVcfz4fJ4l
qo6xTIeUxymXz/P91CpuRZj+zFdOF0gSFCEFW3tpf4oArwmEEJqjl7TaLWmS
+cXEpKFwFxyUGap078uotgI0qzIlM1gaioT3McB2RCo+6jvvSm4cQrGn55RS
17bdrilGxQa1J17HCr29qLNxj/8QTiS9xcGZ6IVhGXneP6kKygt5wyR+LGP4
+G2oUWyozz+xm8d2/AwpxVsKd2dN1R3xoVRQhuBWx/N0v7bY0kbe6ytEbVW+
y8F5/LsLIhk27L/ViK9JN7XD2ZZ/3xyQSTvqp0u7afuiJmWL1WGpXrBWq+bd
FtZl4erGj5pa+xSVnMQ8bBkqKssP+0xNzuY+czrX2MKsGZU9zMsBKN8TcbFF
+kMGcFTAFYDWGvQupZFPFzFtqMzyNS4G8zQxEYharIGGzLy1TxYLgENL6SXj
yyu3QFJARWmSSZHLwqcHdEKYQptWx43iOVvq2JFFHjZZn7HD5jbACp9Uqtyw
62NZwc+U1Cof+goJQhrvXzn6tQiq91yAYl4WQgdoIdocUpXYReIelsfQKvkU
Metvthe/dMcfar2Ct7+QfYl5MWcjNeAhn982+Vq7/8qfORUzxv8OCeOhVjX0
GLclrNaZRnpRlEPxWfRPBvsvHu7Avzh+LVU4Jljb6hxj9Orpl3okokR7LKy0
IQLUzeieDsZapgNRu2hCfqNA0BckznUiVsLxwvlhBVXo/JiZcHOFx2BkDLg8
JLK7qM2wLcx8v6Lqp0NW5pBObXoIC4LBRDCVdRFjKnINdkYArRSRnWgfqf++
YNPfsuAyReyuTzoSKeVq6ZviYbZn5NwcDMjUa1OjD3aaxnmA76/atlYZtAZ2
ZzOyBNk8KLQ31Lh/vNeI0e6Ka/hHVaaSy0d3Vy6OctjU9FpkfIgJdlTtsHa3
8Rrwz+w1bD+ach/9dq0Fe4f6Q9QMYwNbdYxWKM1LChpt6ZhGOMFY83wn8ppg
CqS+yc2JqGM8oFTBxbdV5xLNTNRYkKBbcc1G7oBLBCoHM0uU059vfoC+vcWa
jJCWQpwvuPXSMG//Di8RH7anY4UkEmqQ5y2jTl+wukQy49lpdZVHfRCg6UH8
SHEf03fmM836puUEjY8Crz41KIboF/HqBbWB4K1wZrfXlvI85rHglA519t7E
yqvC1dxbO/4LfvmONZK+XYTMPAsRG1tmjAp5E7vT5cOfsghbh6wajHR3OP8n
1bOCIvaosLyBicqSw+XQkJZrQpOQ3CIrCN/TwUV4+CfPMT6+tHBUvqwPILiR
u0K0/nfUjdSceef80fjbegyf1w2nyTNCO8rzHPDAi9mJd4uSB3GpFy4WUqF7
ih1UKCYVbIkK3D1WOedodG7dk6q+RGPqyhafZlTUoToMarCO87gjRIAtc+lJ
Lten5S0qIfuZ8hZLC5e9yI8aa3fuVXD2D9ZUkla26/cyZ7vy+0eQmYGYXcXR
PbLwf8JIrW7oULn25hKiIjmA6p5jL0lH/ubh3gzcGH4gU0vf/8ZQEz/RKowR
0KQhY8/2utCcP/o7wULTYm4ia0qga53GKtSuN5JYdyaeTn6ROxgZ3W3mwAsB
X6AbsPkSABLWP86D8ugQoltTaU0lXkbrLXEGuJYetY/f+KJn/iKp5G1+QApp
r9vBIsyWWJEJHwr4Kt/go6a7wJMUrWiQMCeu6Z2cWes+m57wlDcwHbR1TTfR
oqdq9HolWfYXj2DD4UGf+VEagUytH2+GU9C95m0OQNZRrpawTKuyycyr3XHM
DxxWCT4DOGF5oPPcFH8XsC4J2INx9eMjITmtKUa4wLnMBIzepWI3SuTrVTyc
vyl+PMkXjSitDpk9kGpEa54AGTGYAh8u4TxIE/6lLLm/zX1YNiZVRwnGGIo2
cRBotyTqkcCwwUw3ZZu/Uju9T3saGbxoVwG2ec4hjk2ngtoQDAYk/vUSbFSg
Q0LIlAEQ+SBlUDXqw0EOl0stNcG+tu0eIqyTA56nJhB9Bj7oaUYrd95fKXOD
nAKvIcwYwhovVRWGQE9b0CIgiZJVDFDnpRRgJ+5jFGNiO7sGkIRRIRPikUKQ
rHAwpSCGKuFWj08/gVHbz0L46kg0Nvtu66J3VmC/dkym4/xy7HHmvHuUH2d7
2XBumnp2pq7xx+Y2/3/nryKMaIRGi9fLyteW1HsvpetfopcE+xkBaTMDHDjm
jY7Lnw6sAGQNcxO3pgiu7TLjVsQzf+VkWiMA63sEiPjALMazNzr7dNAuPnY8
go79HHmGFWU8mwkw3f3jbKL1DCd+9jmKub97jggoyOlOwiu6y5EM06x/eLuZ
DFC1ORcyRUQDElm6twbSuY/5P9VxB8R1ep5zmZJ8mtwGNUcxeX5NM93J5VAi
U7sLdWik8OQq+NJbadNX4PWZCO1GGnZIKqt5YAOy7XYM7o8TJMTJqhJg3PXO
/+gBzMxYsEfQqmGNwNANGCtQbe33cbT+kNFChdj7plOQZapxKJUNVUhyCyFu
ceD8w3i8hDbnwZnBImctBThsbor8rps6R+4wNvXYRPnUQs8/MQTBOhyKq0fN
rHy4xdRsAURLGxzzE7oDaARMJH1dlcyP1LW5dp5XClz08dQ/mJyDaOsIXT6S
hR0RSrGrv70J3AdblMmRmoWHOyflvMWm19ejTbrBaMzP+76N8+BPxH/slM0z
789bq1nrCoLoGlWD+kC1anU+6dVI7NVaRyo+BwDVamEMeb8taA8/n4eQGvp6
sd6EcF5RRxM7M+wFsSYOjfjQWyYdQ/I2OFCo968VDvbppL6vebwuxuczwbc2
TovKmqoWvE0TTaC+gSm1Mc7fILR4wxoGMGpqQ+oRUE04bAzh/l/hVBtzcOrc
Jg4EuDH8oK8Dd/QS6DtrTZ9EzLN/cSojqvD/rj+kLRaxFhoB2vCQ4kvD3peR
8nx033y+JczhMxb7gqqEB6Bjb9ChyeVhM5gPX5Srp1d4MVYJOis9adNZvGAB
kjBZYSUv+s3lQu2m2fOc8RJu6ZRkNBapThox1OmmBwxLj5PixKWR7+2dxbv5
51RshcQQkJ8G0hW7TG1rbkqRH1AHRkkEv2b5UxK8g0CfOOYpaSmK02b2XbeI
D9m8IOTF+rMxPDPbO8aDyyV7CKu/OVigUu8JAdVsiCi7EoqtXmJV0NdB09H9
BUWKdHDh3s3UrNRwWYv7fvrpPLY3oQrjPbNnOWA/X8xAk5qLL9uYhdzcmtlT
gZ+JORlmz7enEjPu6vD3APLZNlYp7wUYpI2kApQoFJMTEBE8MbgshiAiyHEh
HT7+bQ1VCVcMVO497hp+TJrKVS5RNtS9ZMebQi5BjuNLXCwhwQhx5VH20opy
aUGiLNDWD7R7kP4SX+1u4oGG415G639JizcEoPknN4CeKuqMkQBXRK5I3xKK
hLZOCZDaA/X9FUOB7Y06obID4GoIXd4Dbr5gr2l4mM4kRX8oPCqobl3Pofiu
4RnUdB5b+39Vd6lfICJqdlBlfxleOiwLXr6f3O8OorjO9EPnR6Zny+CZObJY
6z4+bMmJopKNgr8496++YwcAnfh0klrZnGkLn5cv/lC1s3e7QknR0gpdftQj
7+e514DQ7wiv6Pen5d9P+BtYBh9bwtHBmb2ap1FCM0ZyvQtdVc2wsymmp/u6
NjpnMuXVE/ZyQZTr545Zbe5QFMRF3pOqjbrEpIqZJ1wYyDOcbeSrHrH0gLqf
U42WzFhkNYk89n3NO8DuhikioxtsLIrQXYvpKg8HXZYrM7PPWo6C1wlK+HhG
CdDVSNqmHiJLq35m18SlomFjpnFFxPLP6LYOLHbEx1Xh71nWpeqHHe3eiZgd
t9n4F6+nKlZPqQ2VeQsJcajFU9mTgWo54af0Ol136+ZmjQGKgqOerJYsVMPX
BSnIV9A88awrqCVTcYRA6TAftrqgINESwi6UGnYMhfYwXZl6c0P191WtIgT2
jgbrLty8yjYfsAxzvtjRIt26U3mxsz1XTCjtMcRI7swQjWv/E6SxR01AuHUv
EdIUayMWjSjhvmBqGM5qCY70zr7mi3uPR9cqEwQDrGU0zn6C8JUR2LCuvmrC
nQXAx3yqgk+TC82iYk/AugFIGNVAk7ceaQhrjjjSZS9DqLND6j3UmaEfIgQZ
ytGPdc+Xh1I5rHSvHdJcXCPUN9sFEQ1UJpzduAkkAN5j9+i9rAJJEi7n4q2G
U82XKqYJQaliDeH+m/ZERj6lBvd/3KmexjejuqXMvPuSVqbCsr3vDN2t+YnM
dnAhncAUvpXjiPLHtjwuwTwN9ymGA99hsIstvRDkjI8qqSUl1GmkvhuqGSux
rIgCdNNL+xxXGsM5YkgoIBf7qbodNfMzn23Ae+iTTufRH9/YNORVEp8ZmHZd
IC1AhiZD/egXeeRy95T9ot+buhyrpmVp/BvPVf+VngTGM9dwPn8Jd9/kJbYc
uu3hEVReECnnRgaoeKG9434RmYi31gVdlRD78aW6OJk4t4wzACydxEel8Dgc
+ESzX5H0SYNqOGymZa4ccS9U13+G4YQMbkqQRG7o46rQYROHigPP2kAxphYh
cP//M3ovJAm5GitiV+txoIw0rbnyIrPYP/U+q1ObqMXwKmgKT81dP/L+GQOX
Dn+P5D4w9K+l1YONP5Vgef29d6fsTD2CrUEje0+zI+ZW1HiN3y0YemENQR7u
ACniKKhfTVtxvBhs2sCjKrOBbqHZd63NZ7FzQP/WwqpJg0ii6tVEh8QURmLs
fwT8ysKnRy0lIsoJYl+uXrYqzA/AsIoJu7gfM6kjjHvjgewsRJzuY+l/2MQ5
My3IkAEsAzY35HD6wXMJMd16W0LQnRMpiMREixx3h/Tu4jCPA6JLxuFdlSGH
Fcv9sj7V4vDb47cqsvH11S8wBlvJveZcvwUcN/DbI96RAOb/D+XD/9th4sDT
Rnama12GBXYkMa+wI6XFXyOntExNNI3rk3psmZ8LlboFAHkSHFClcI7QbW+W
zTGjJ7uAMC696ftUat5DNctLS20BxUjccOBIwz2DhEESLFt/oZqQUjMgWAN3
SXTohkEFAHxlDbsuP74kgrcwXnaca9BjFOkzWQRhVEXi4MP9g93sEkTRKCGB
8Co7GnPtG6V0v20TlkLigTDQWuW+5VBhuDqR8UH9NoNgp+eXs7vFGxrpZdnb
NirpSQsg3hq1ANsLFY6zb2IE6q9loGsMo6i363v3hzjsvsErU4jZWo1FuHFU
6JP1NUiFJfkS14j3O7tjVRd/9vSAB9U1XmqhJLX0/T/i0rJrJuV4LA1D+mgy
N/VCY07lDxB6imylsa5mseS9Q/HBYml+vR+Q8gY+5upVOXPlUNW5N9hkcm19
eAfuXYPV1z0LDEKyI83j8gdqExf0QARYxpjqs+D2dEiJKpmfJdtzMy4Opq1a
sKqnK5+69bVtYc9l3pouTFyw6Amk3zRyfxXRps6MtVbLiUXRrpuUOgXYm+D6
FIrGsM2DaKvY42ty21zWjuLoCZq/I8gA7lmkKpUvDkDng08imJkYXI2N24Wt
tcc3te3XLPPcNDLKlAGiKharXrZa4uWamBuc8zb14DEiLA0XiHA2fUkWpN8w
llcisgPsrXNkcyz5V97qAfjU/Dk91sIrnDgExAYkuFwL3jA1S/yt813z6BB1
OrMOm+XuB7vrdMt7cXHYAQ+kPqoeMToVurU3e3ABh1/LP/vwCcZm3J6DS5ae
fF6EzTZDJFjU5JeSNh92QBm023gG3VLaso9rJLI5u0qmWex1vmCaLK1ivU4l
D3KVtDMqa4tmWJYbPy4nmjjiRUjUBSQM/1lfRvLwkED6okhv07l45TzY4NOQ
XiLlU/5HiJPtR9vAdDeQi7M5+g/3p/319WyKJJFFwP4R3AGWIznIM2Mtsds/
/Pnvig1m8PW6fQnnrNz9c1s49u+ZVyRaswugpEORy9iJreQ+gP5riGKmgs4Q
x2MUEIYAGV2RuN4dZZhUZdBkoBLW5c2DNk6MfzLVKnK4hD+lfzsx7TAUrtHo
xvXuSNGxLl7CYGcYGYWFP6jpT+KyXVB8S49Zg3RjmA+1+nsJLwYBTkKWA2ZN
eJoTtsc9E1Dud0Ocf0aWTYuqkVZH8JkFqtYLfYvWUDPTWsOHd1lbpllMjFnR
+rqzZszUu4uHNvR/3HLoAkBnOAMIoKc+JhJdJhH654JHL1st6m1tYPh2AMgI
WmPv9XrtscIQSgQawo0DS3wVWKiR5AWpXDNu78359M/v1yvqHbjrTzJ7rzP/
vKuZyxp7Wt8fbKaQl9y4eBcUBZOXC7J5fkDVDJSnb++BtvKamZwzm5DdjCho
Kwp3BpkWWG4ziSJ9r0nBFBN27Qz3N/ihODkI2eNp2D/H6i4gyr49oCLpluEg
FJa9GwJx0/BkfsBKdLCWbTOH8btZZUlN4grPnx0zqBVCEOyhksOpWE+/hdFw
3bXHypsSn9+5oLCivIxXX77KdliM8Ukm0zovQluQlH0D4ATBqYK9j/i0yFR1
a30pPUE8v3JFjhAutuNcy6oi6uvMkvokv9xfhT8ON4g5xfPrvIFPYPcXDh1O
AJZ4fB7vHevgUl4GZuZ6lgdrOFsTDRgxdzTNLDGmRsz+2xsBK1w83+BeeJ31
fw4d5Cl3yXxQRitAAJqHQu+5oGW3bmdL/NSMLXgfJFgDhQeNakF/eCx0TTzF
w/jje4OahF2JUFnX2I+6ks5BzfofAf3SNmSE/oi4ul6QfUG8YTxVpE3I9nk7
SpvchwGAIaeBOmySJ7dp5LDZxcpLyAs3TikACqs8OTKuW8STrkwqHp3rYL/P
wAfx45Nsgx1x9YYoOxMomgooWErT6Yyr6VfRn1Qs+oy8GCqDmvzqIr1faPVM
SYQVNeV6WAU8MCad6+DuaQA54ZI8WFhnNTx/B3MuhYJGfkw666tjHLECLeSA
u9SNUldAbZ3bqLioW77+2xwuRwmGNn7aEcLawv43F6V+aXmTUE2eSlvjEcT+
bvH31ybnnedWIjLm1VC04CcdNQ4A7FNktqAJQLNhYJzimgsQYtfagXUQPUiY
l8ZneYK1jbQ7NM9sUdmQKVH5nlcleCXIffJCK51sGovmTzNCHMOC4hlnx0Le
VINL0bZXclvvTenx55QasGUWZPOxVgbrnaO5ZtvF/p5A/WDFour7QBEBuNSX
Pkzc00AuksWbq3jmQXxjFbfsIx0QwOB9AJ5Sg9Li8xtZIngNY5lQl92R1C5Y
CuLn2O7u4G2GK8nTy4Dbj+ujyn6jzzikMu/Riqhot8wJgKGnuBfl4Us1vJxr
vD6dy4GIG3+GhUR4RiO+J8/gAh9QA8cD0wkl/6rBZX/emobnnzRVzWNutr5l
1DxpKde0vgOynWRoKA44/G07pohWUdaSRSHyUoj03HNcsPen16oyuZeHQEeC
jyMShWO2Vc+7FgO0uJRg0nS50rZM5/sqHgRRfbRlQ4f4P+53MIGu1OjNbq3v
62SK1H2Z42Uy/2wm0gURnaoKgyqE9MsFwi3GfVSAC3F6n9Rg+g+KR+igVwji
WF1RtVNLJb891E0aO5ulHg2IneUX1vsws6h8+PqI3ZcDasgorfXm9v/3ksp4
Ce+QnALOFDsaESj6xTC98suAqkuLvku5Eyc7bKZvjZhhYwuLbyj0ou0g72GH
dABOeUFaN+YqvVDvZztXWwfJz0n15aXDlNfFfTtXxmfT0sJoD/2VeTCvNhNP
ftXC40OsgmPGe1WFmoBpXY1P9dAGNOA2ZgjkWLOCGhAaCaAuQJlXwM5w2ADZ
Xc1JTrAq0vvClJPgNKspHD/ze4QKs6kHyAYZz/+ZE7K+SBCvicSwd7kUtKU5
tB1du4YShm65vgbvYbponb1/IsEDHf5i6hCUDlMvOVyK98B3viLHbtzSceV2
ucsoc7l4+pSsTDdht57WMfGlpC+ybQBjOn9oBXcfi9/HAGbG5P4iXE/UXQ3Q
dQASOX5Mzl1efx9+bmqSoUD9zqpFCTYzpBcBzj1xVp7XEJNQXk17VUGC/fLy
om0IGae4my90FMkYN5ebI+xu3Q5W/HvvSO0E0ybv8dSBbRD4hIHoAOYjxB7j
775JcMjM8XcgwqidKEzTx6+UM/MAPYgCC4ey34bEkpK76O7j6mPX+7/r1D1Y
VL7WM0ZtrTvexFm2PBH4NzhXz3UC2sXkeDe9UcXolKC0XtR6E4kTQG18FzKL
Ftonq8pU/Y/daHvowtXbAy07q5dP+WmtD+LrXh6M4CiPnsw+QAUiWvc/vx3p
pCGIy6UH8FgjNfGi6WYY8wskgYXKdR5PKuwvtnlM3KpUe4YcSmzSvKc+ldO9
AwW0UnAZ8elOly+8fm6IIREDHKruNMiUAVppnbNePs1aplvM1HqHi0TbTT6m
WtDfy1dywBHKQBW32TRTA6wppk1Osz5adhSQH+mp2kR7ddPFIe5yub9ixcQJ
SoAHjol4dgpCxPzqhdivZMMhcz6HRb7QqmNFRITpcm8IEv3cnbupw9UFYUH3
x2hub4v2Uc4hpQHjT+jICWehYZ+c8vdgIx3T9rsZRBbNn+1z5IA5odtV1/oH
055p/WcgBN6u7FFUJcnOa7tTRzd9JyaW8anIgMW3Vsm5j8T2x+o2YA/ceb5b
Fv2qTa9sE0sd5x7szaGnpOd8J44fv/qZKfd5lBYQ7fOskdcJJzHYjZOw8rBj
kwEILlW9iDv9UFSk8BuN/Skro21AENFOXNkKLKHYVJQ76LxjPk7fAnCrVjl7
Zs0uk9N/Y5HqiqMG6ofW3Ea6AqRJVDojqDym6mDNh3lJ0PM49TOfAde1/uUE
5C0NoCH8/1Lny5n335esblfMQ0p203eQICVWInLaE0niP0+fgsOOzmlIb3Ne
9E+lcRni1UyjpcWhUGoNHct/IEB7xZo2PQ2sY9rGZv6tVCUr2QOQuzqYtIqM
9b+zyBDXhgUXeZvYQAfaJmaksoJ7ZjiLAKtHqMpuCSS/fMCAdfB+X1Gy6roX
QYwETVJBpNxPqg96G58WmcpXznqnAxNtOHGaw8ked1VhCvVfa4dyLP1U1iez
1Su3lFVlWctjDmqLa7VuNZMif4U6h61uAboHPy5PYW8KxAwvzcS+OCdSmqKF
kma27fJu7La2TjwwS43I+ZZdTMERYHStB71n6B/RLb6lZgwRMnAebVvvaWnk
IX9PyU2Wpe6e2btDqpBuhJlWFIBXbO8sXxDv3MqY3hmW+k/Mfv+95i4Oo3W8
sgHUFfSqkXZx8Y5Az3FmGVPGeDLrEJT17oy3EFliGo4PEtMDUeagNX2qDpSG
EZKzDTAVQwnfJuQFCxRzvCIyDzfTUoXJnMqj2Z7WFUzzFLU7Hp03eYqHzgWq
TieaRWc/5G5FiWSCyYKO8E4GnHDKJUTs+zRVXzgLaa950yFN9G5NDMY0YTnJ
HygIUawPNJ2B/0N5TU8GK4bUwFAUN02lzUa0jj0xtS1LuexDy1r8uhbWn1Eo
KQsWKClZH0YleDyR0azwywHfhgrLkYh4Ak3DQ79a6Xz1pySa+s6mNveRGyw4
u4oBDPqAm84/VNdiunmkO0l5JyH+Y+lX/oeOsNlz8r0Qjqm0fA7o/idRd7QD
3lBPMHAC9RY0eEvHxE/WA1ToB1WW0dRcKzR6UAnYD1RR3bNuAVQaGTbmVzTM
oE6UwOnQIwB6yB31o1F8EUlJc3BlpGGoW+MkMzar0IJbNDxI5cQtNA0jigGE
+BL15qEZbFYjgSDHEG/adZJqo5gLwJyb8F0qeaFHr58X5VskbrFJZAlNgQXT
UNrzQHZzVJq+0xW5PWoIY4jblkest4JUVht8+Y2GFdmys9x8cxrlzTi3rrFc
tuGevhkBP23pLZHUl3xO3iMz6h6Gv6ZwyXk8z8pkW0/sEo/QcTscOtbBrl6R
PTfjFPW0k8GqpLMKH/nDLCZjQ/vRVA74h3d857JlTXw3xVDhMS3MPZJRd8RC
I0j/OX/OB6PZeQsRHH44raskwUJE/XExK/TWcX8kJ2GzAEcHr3mZHU1zeA4c
Twkl7jDgMLOM2onpMGKBoHHjTrhUDI6MWFPUid/AyWhGCgy720urUMHrBoyY
OiESIIml/apWItCj6vPMoROM+/4uNVp/VgrFSAFgk2AVIgVo8RbD6+bCEbh5
vEZGhFhQ2W5Z/8GnkAYJ/RxgU3E9SWJ8tLIpUgvO2prTJsHTixhHN62UHtqP
kh25XwbtK8Qt7Hq6c0XLtZ0M7IbQVzOaSh+QWTTn6hMlA+qBrVmt7n5Gz38g
5SzkKWSNhpP5VuI81CrNoRFOA7Sge/nIEY26Z06buF90ZW89ZrIaIjSxnbA/
pDR/XgD0vclMrD1p8bMSDe02Rw48ulxPom+f/1n2e6LQRtzsjaV3C8TGT67g
7tsA4L+LtH/NksyXN0sf8qUsSIgZkmUrnQIi0IP5s10Snx/e06w8w4aaZQyn
fh4Sa7Ibwnlr/DObQu+fRml8S/B0RmJjJu4cT9rQqT0ZA+bLHARTe/sAU9v5
jqjAKsryCLckTyZnZY+0IZfD+45YvDoYqtw+QRl6a1ci4Cjsfr6KtTSPyyuo
Hu16LB18NFEQZNXppclJbdCw0s5eMCUCDtaZ/+P3Ztt45MLb92BNpZsX3rpu
ngdMEDoQegOmXn20cbqB3ABVKW732w/mqv/p5gKnD/n0v/3Gi0aWI3D22225
zT3NKAHkE/5Bhg6vQVamvV6YIrxW3H0JpMQ18VIbcaQHOeQfpFfPxmQzvaag
dfMI6MPQKUYwHdbh1ptWsnaXjWjNOBIdv5/Q22Gvp45jfBfO9+Efy5VNisa6
mmnS7EWl1LkisrhTa7GPehCaob0b72vfocYAaBE1MH18XftdWLUk/Ogb4P+k
WrsRgh5D4BsB7MOj1cCvzyu61xZriBLmWI9g5oXx2E/6LZ69GXkc2eyXZdoj
PyTMv3y3CVGRQXP9dtlxJjDNyZaH71BOAmY2S+IRdxDYYsBxogI+dnLBskyX
RUH5Ly2HYM8KyNChReXItcjLPkkWqKGcA9dAIICsdXnwdm5VDsk+KxFZpN2p
87qaN6G4Oz55xrqDj5Qi/eBVLJI6Ir9s3q0m7WEUK7LBgdYLqJ/M6fXr6tI9
gF0LrfVBrU9reU3f5tWJTigrwZuwjX9BhhVgRLv73LrE6CspL4O4HhCT9fEz
0/nF6+yMeSbPVNWWBt2drDhhh1vdHV4zxMBYu4cCPOOD0ZMlrfzc7cnEd+je
OW7j1kCTvk0GFxv8ckNw9qKimLlbajkL9UEW0jNtRVJOBOZmKcb18OT3UOWw
OvEI+Ltt1cTK+HJwTFP5+DqKNj3jZaa1c8BabViOWN7tYGZWPBWgscd6+lBP
jsMazmGVllL0mzO0XGJc1Q2ZS0JyiXn5mb3nxDigxeyYaTdCFiTomy8r3BzQ
JobRQWmIOUY6MB1MaSKOtHJSw4cvCnkS2hVHcNJJCKrViCT0Tg0QnWCvw+CE
S76RGmnqj4yVV+w6vsqgoqMbj9QWWT1KPADyWl7IcL/v+oplmZVr7htcgJjd
OXsCororjKoEZRvcc5IrjcUL2icfHRGLneP7bM7tXxDwC/8gEI3ycO5YiCB/
Bfa3p6tAW9lLdHziAIdiq/IL7py5BImb44VoP22rZ/gzXQx2kygqt36NXn5c
kY4K3tq+jeOyrhGhSiijDWk1lzbKM3vg1IF5dXs3AQMv9K2Tf49Du2Cnkk+c
/x8rhX1iTGAsdV3s/DdWjmKbUqI2xvZTS2hOn5gyvUT0zn2W/OxSzHsLzyfz
Xr5CFjVtD2qaZjm3ZqwtXWki+J1zjYz04DpywyHhAdT0t9JGjLpbobhmJleh
6dHj5VLcZi1SApd38VQxFE1CwkOUQpF9uBTCWjFaoaCheDb/R7CpYIb7j09s
VsjKYviaZLIDnJdXABz9fP7KeTU4IVEAPGo3FJW2opbN5ZO/DtWBlXiOBtOv
iTdMKyodrb2YKvqcPub7YAFfqDoALYpmN/cHa/71WQ6TNK4vJYsouJlyAwCZ
yEFzWNcOw2d6pnGi3Z4boSghzAoff7Zr+yydMHdSY6Xg0t8gPJzcOQ/m08Ml
Xrkz+mocaVGGzz7UA2FMVAOvjqVJMfcGEoceoAp65eQ0xQ8Kjd+5xpT1MjHK
YP6wzz8nK0vCNyVz2o1FM0XtqJqRFB4MXuQQ5hzCVKn7c6Q90xcQQKdVfRO/
p1mJle6ziSdUEpIIrkBJK3Bp/CP5K7EOEN+HfyWEFcw1PEQ2XDhq/aAVts0Q
g+qxNi5SaRjHB7+5rva8i86SUqsEqzs6nbH496Q+giNn2RBdhU0z4xgLYzeQ
tyGZyKDFia3Di7wcn9VK4FzO5QbaubVUKvd24M1U2DQZKeG2cCHJm8/7bQXU
OO267uwPmS7uUTGYYHOAiAGjK/cRrnbUVEvmc+9Js4xQ4gpQaY/uTw8TK9bI
9N0dvZak4jiRi8bVD2fgRT3BJej/N6z68QsaiO7/aop1qIE45JKJj+3vB8HI
Ladf45yGg8qPPh8eaFuXO8Cvw+ts8bRWxKwNJBZQF2PtLBGa1uie9F4TY3Fg
GSJiMCODsJ0RC8Ho4SP9WsWhHblThxswu/1B1ja75kZVE9EJIeTf5uHyWCHn
otd3go+FasaO5HYt1CiQbml0mVj9nwoaBR8WJhBi2MWEIv0PprNOyRtBgY9E
CTmf/iYK5BtKyjojafZ7Hf1DTBCsWsdYh/AwnGE6Gywi1WQ+4+RSYoWyIkQx
9SVqaZPbL3rKZut6rwrmVgMTxYg3jyVAU2BHCRvidnQtXGUWbN/gu3+HzYK7
EKmsRDCDk8Pc3c9sA0PXw0nnM+1XeAohPwc0j8mGWVT+lh5C8ZrK6izYElIn
3mu4v8KvqWaEV+UZIS2NW3PNYRVNEWm/t1tw+4dJnhLnu3jxhx13IDusvbwV
27v5DJAV2P3eKKeraz0bLggogsBo+JcOhtKVxtkFrjE5XoRyfGtErVZ0xOyI
xInKtUyusQO8bZ2ZUxCFiOkT5VriwAogYSYT0c+LSAkwctYnJewRP2z96V74
HqNkxPuXs3QMzh/b2S781kOUqAh0Gop+3jmYrmoBWyQxFbTkWtjidheD6BXP
JMDFTfdw4j8Hhb6nDbYOmUxGgA4gbjAna1/ihHyD+1+BdyFo5B77D/SlUhE3
YH3BxXhNR0am22m13cmqXO1YHIE5vPrRD06EIVuzWfD32hC5ozzpwte+WoP0
m9ak0IZrFcf0Ei3yjR3wZ4rgcdfezi1lgCU3uq7uceu2jtpK/T5azgQuJ/jI
bOy3FVZi5j+dIKrDGfCfmNXjMtRACXWooFMln2c3dpqbTp2w5TDhvt3zCBXR
9cMtsH+HHFSTHTgPOJjvF4I3G2hEFKVapFOgtWcM4zZdMWE1OTfw/JRbIA+x
FjVBN5SxQU+RQRTZs8PNKivv03r4/vBhduvZdpxQMLArMMs9AO1jabeYthI6
zsR5egPkroAAZ9CiKPLUGq36ajOgs2qctoXSyK7xMETy9aKFlvMVHrwgwCja
Xsh385lAx3UdfzZbKTUmLPc2ldKa1Ss1Surl5kN5c6tlL9veOcDTn6ZHw4TD
EyAK3d3n1mb1uKaB+Owe6FKXj8JPhvP62qHShRcRdaKdqnnY7n2+ghx4gVtV
S7B0Mt/YjeKyXuDaA1XhUW7v2fY/nxfTfZtb1vh3lFOL2vOOne4HwIYd4YYd
fsi0cMCMC0o1icZmClIkPSgwz0Yqo8yJqg/nJc4/i9adUnS1mB4Okezbfij5
VOEnf+753g72aS0xUTQ2avMSIOqTljUMNjAF1+pNtPQz/9JpPBPPst5UeHQx
MGySMPDPLACkJ7AcZWARVJ7alE2bYeUeMjWwGw2mHvWqHYedWi7jfFMsFT6q
GyTJqr8qFpkvOHsXCgEhkixOUsEu5ISTGKUrvNWLoQ5U9KXSsj1et1nt1iMD
yrF9xD6CiQ1mNuLe66ayL3YImsboLLpaeeKiJmCnuOFl7gG8TZ71dT2nDXeS
ah76/CEzW35TnGMpCmhv8kBkv8M4MCoczaRoOA2Ha1ML3STNTLFJLnd4y+5a
61dmu+lR3KWYhHPRvWMz2Mvy5NAXWsi6bTga7/KcAI91x3+6/q8uIsk9X7BH
GTfQbhaQwfMIHzHya3HOPP3ju7+tLwGnlc8EwMAI/ZSGyy/8Kc1jSIX+uMVR
qoeDLl2rwGDOvdSd857jLQY5yDDlbyBG1qo0EsX2I2LTN0yTfpGwZUbD8LmM
HwXWy2V+43x1pUcaLnzAtGKP3t5SW6rha933WAzCPVLpQdkywOHy8WwEgjO0
jhn6eHVBbiMCXmqXoAI9pKV5RL1C3A8DpeVyDc3fr7DezrwJ01qS5MlKChWR
k6APKZFHpwBOweuCtwq+nUcZiyQoI3ANaCfgr51akJmDB6L3xKsRpwI6ln8+
39SaYTM/817CSmwVZdXQReH/Z7zbn5WiG+hA4XeFPktGRTmLmqh4bmyRqLL7
oVmmM+glH9vkKZMn5MJcMPhQfYbEJYUQ1hYCAIgP27UGmcTli4zRUo8aj3gj
rCkT9gyp69c3nWu0FYFTrdvxJJh2GF0MKfmIK+TUhLwgP7HxRi7ciOflwYsW
6PPsEG5mlfrJFR+s4fVDQFwRy60uteTzNg7SIQ0aQq/fqjOOgqgxrxg2ag9F
sHj7lmkpwoXXx+OQi3ixqY2+vJ7LlduzqfCnGLsQt4sYpcvFoVlRoitOaGcA
dp+OvXSkfzX92P3/2rbfbcK86f9BEbvgQCQJtTB2IZ00XArne5Mtw7KMVFAq
sh2jmRpfA9CG/AUbAYbrQ148nEyPp3Yw3XfvRODRWe65z9dJ5WID2rYhlGxX
kxNMlsiz+xdBV6eL/XkcmNLsdITXfQHtIGshsUtB+B/ZoqUFXsLjO97CXdbV
OkRawJuXpTZBd4vu3NQZyPA98uySueFPQ+ASi35ZK3xBKxwiiS2yADEQ6LyI
8CAU0TpIc44RBzaP8pAui/FVkj+43tDR5D3Lt5pi+3kPTJXErYGT187PFgae
T6oUptkbm3fN9oq+ezLjms6uMnjjpSnxa2bULlGfATqW8hjnZBgpAIHkVtlJ
UHPdieW1QPBx7PrPn7J1B+RPKDmU/GI3xJRgX/VU2Y99bkyFe8pWmOQZlXa/
Z/4aqa3sXK8xbSQMdV9PMTVa8OVieW1cd7XfD6icL4tH/pqY1tuDkWzQB8gc
6EX94weiAi9a9m5N7/5q1B7x7NBqb5xs0fp1zmXyGM35bHowPBGpQceofKP1
VtXQUg7+ZtdGjNHK5+680P6TPP8/cyvoTBp51qbyRlMPK3uq8D4Ob8IuWLa6
D2lWQRrcDesQxVSIEL9fG8wIPikisPeIaXvWJDjqg144loayKb/hxOGwa0Pt
4nzlt9nnGHGIpkJp16wu85fIunx+8EwU6/uO7nFyWmqdEOOhehl0WGFe7tX2
6eOA+rQcHuiTYQMTRJ33MTm3X4Ajva7quSHWUTY7Ka9wd/Pr5I+R4DszhTOu
b6Xn0fAje59JUj5e91iv2zaJ9uowDMe8p8QFvf0F6k8oujGWX9Hj1Fw2qqKQ
/ykh0Hf26SFGY3IEJmGZZW5RPzQVNIrHTQAgjq/LnErWMq6JGnq39VxfBbHd
3DIUhu7SGbGwxg1FibEvM+BWFVoQ+wt0UK/s96dG+TdOEntPYyBW8jK6k0Bs
N0B3RgrE4dwP7QqB0GpgEmj0h477vFcP31r1SDl/77iHJhq+ZHdJWnaqQZNk
r3PQLXGXFCW3/48EuSc7WtBnEL9rTFRTFQ8BBvmQ97Jk7AP9/fvztAKg9+XB
YUFI2dmHuMfbckdl704foKVuubR8RqnPIuhJHAPIGoJJH15CC9JQO0LQr4oW
1PbdHpC+6FBmB6kTnXbVoT/zNz9BbNXNnCDyib/JepQOI/VdB86OZA9I6ED8
r8gD5WFqXRSExDSJ4d+RCkJ+svT7naHkhWkTwP0bgd1dERhEDlyz9rPvWEl9
gNS6EYgs878zoCP7MWH9C29I9dEzXNhTLimkfE3kjTmyS+ZkDXZsdgiqydC3
Jk9wmoYfaRH0eU9+JKrCodQiKdsgVqNR2CkqhJl418hXq1CKFpLsWe0dcbrL
6F9O22/VBd3BjgCojjvUrl+ikvlxS4kGQxBtrFC+3ewefGKMCnXaXGlJlu0+
cE/u25pEPiPc8lsMGRG3/7VBI9HLOf9UdmeGmGhmjNk5QK78FgmCpW8D3WWn
YJs0AEuTSE1PmJzcgsdtVvNjY1Ag9GBuADpj9PITVtA21GkmRGvnPSTOY5IT
1lWWxy0/Jaker/QhQCtIiLYJnuQ7tKPt1LZzrV6coIxtWFsSOce8YTIwGuOG
uogZ0OZPYGa+MBTw02G/FoefjE97VhBeGaLxPYT8LSNcGyJJECZiK26nGJEJ
bBnXguW9QTFJ2gOIy0o2LHyIp5j1R/YKJ2FEmOYeXNASNvaenIMGRqTXfOER
Pazmpt1DIVD2vpWQHq+TTjYo2a7rTZ/+GdDlOu3k5rIYC7y+4ohe7rhR5Mxx
ogEj8pH6mU8j9P0qrgD/AKoSUd9DS3wGlQgR4nzFn2QamqfPth6/tBtbN6Cb
JlsOh8IqfYTIecMwkPrAr9xCTj8u/27pAw1DXU2DtOIM4VK6uD2VtEV/IVVk
RYHmwzxXGHZXYwVdFDeWOkQNNr4JgQFwW3DWATvTvuIgSb1qERKKzZgYoC5P
K+3iH2lcJsKSP73iHC+QIdWmAfSTYtml+lZ85/S/fZkTtnT5EpiBl76z0rBt
fHVRQH7YkaCJ9ZR3x2t1yHbV/RjNc7UwCBtviSezC2AWYVMzPjxE5BP8E9sd
WsWwK716d85gTZ1/upvCXFQ6zirK0oj8/rrmB25Hchrr48WwC/JCoaUYFt3K
77M7XVVUT3UjZtrcIYr4wVFQrAgU4dpGh5lh4GXbwik4hTGdp1VBdvz+HTqw
mVY6wY5CBIphFSZm/C+UyiJRL6ku0DFsm5U7CJx9z9xKaMPFFNaScZMW6uUZ
E1FIjtZsYzPkOq3EzuceWJWFSO8WNSCEBAX4TvkoqJ/v+gMSB7EaY80lzqpa
nzgD7U8O+rRq8qvKIxAc1CoC/dICr2oMxIHt4QZ+tAaTpQWuQUi74J/ai5nq
DUBYpFPW9+fBdXlYA6+lggeSe3J5z6HQYdiwp5gKrPNerDebUqo030TfgMK8
jWrwKXqPRI/te+2G8f8XVdHvWVpUrr7gTT8OFgmuG7ShzbUVDK+kqQlN7w8U
lMsQBHqgKhDZN6t8G20lfeJIrOyqa4uIUJ3Ne+0p3gIC3d+fLIAkGdN9hFBd
PpCnPjM/K2fN0OJ8Hp8GkuLFSfHVIdpxseYtT+4/syKi/mTkkKHJWQTHxx90
2flMTzBPzKM5DE7HUCfSp4Le3joejtYwPoYGndP+zQBBJiY8PN9N0BubUH19
elMsRJVZ0+UqMl+JPkt31uWWmY8DNEdrxsw4+ZWI2t9s1vkIITg0nR5RIQFJ
jZrXMBA5byt1BgswbLNhFf7x/8x8XetFqzHagGv6AneXnRwDho8a86NYq+AZ
VE0kcy3nQLP3AMBk9xnlJCLGKDUZKGg0caC+gWxzBZMzKZHNb+jaJmpm+0kd
qy80cn3qzXeKMXFCQWtpG0ZrjeBXCTAlHfGoIPIjTfLvbxhVxpMnLl8JRn60
U4xrYcCrOWU0TA/gE2SI83nSKfBIzs99eYuof7h7t0eyCx2Jz63biCtoRMCI
I19Ut/OOHl+e0BEyjv+zJ2WJO557dpa1OmRRe/Zs30a6iYvvmXlu1y8CgdYL
MYx+iMb6jBiMI5+/gy0GCPwxFdn2BSIypivvjc6mDEqDDoLfZFjXNMsEZ3I2
OQa4+/93w9gtxSJ3kNsxGla5clu3sCH7nyVMa2QjFsD9ml3eu3g3qpOngqJP
9RPdTsE0vX0YAFhdGnYArtzZaBgAhZnwYFk5iqCIWId30vlP3XP7LgL+R4Jo
4snY9I5sbekOATSTuLbj+0Vq3oUWGwiViXUAnRMferFRUYmip5EnBLNNwDkB
Dgz8lWBsM0rlnFUknxfrczNtp9z+eleg6Rf8AjdJfGVVtI+q3kPxb3hoBU/D
5d/UOrKKaNi39fo2EG76EZyTzrkCX2rXN96qJ3jLdPH/NGjPzpazms0ApA0X
6sHLwrnaiZ2oIfG7iSmZ7mKWDHfDNTFF5izwNwffE290MMDpayDK9/8+AID0
aPsAr+DtWfcinrB9ATn7Gr78C6bhLSQPaY2yGTFY63nVTmB5Kvl8n87UjHxq
noESOZzBY9oo4J2VdexEjiLMU+Wo2JDlCA4OwzjDFQIhGpKCdrG44lc6B8xJ
finLanjrdDL2j5NbdAf1niNrTDU9uMnkxt+wWkUc06i5LnroFQpIEo+VOOWw
16RI30QEFXuva0GqxlDfvmz/G3y79f5wITf1vZzw/C3SxInZvf8V3+HYyxk1
kxIzVYIP3onGlzRi1Xjf+RDwKXWrHjuCjJowFH9eEZWXmdmFUfi1Itgc3Wof
6S+bOyVckOLKMXF0kLGLsEiXTR+7dbOpX2mp6QtqloNoViUDLHHDUvkRJiV2
GWSoYo23gfQtu8MRA1nIi+aB8VkarpfPV2K1OjBB479ph/G4aGbb4muta4wK
eKGwOu7WOCHmgyxbO5zqkkWWfzm+1QYJVbBEIBJ+u3T4ITtVvSLK4vShITIJ
3rXBJASMpdFYSJQC5N5NO0ZQIeYZ08014Liox8q0aTxsLAwu7ctz/vj3aOGf
J17NTiBIl/GujOgJ0YMOybUqje8y5M0MQFLoYM+8p7im+Lpbs4f1YiLE6Jg9
IvmADrde9iYFLhL7JF8UWjQUGBXpSYBhcj1IQOi0Z6Jx0MoogJHJfZZwMD0l
++wvz6Lv6BSsHyP85I7AsZY9IIHO5Mk05Kd3IssQaBNC5NAK+g0N+RQkemQ5
tbTdEDQ0WPRU/Au2JAAeaxwFMXEgZNQ2QX3qAWdu8f1UImd0ntEw8vazF/qS
2rFkMN6BjgYIpB9a5KxdWpveSmUbxPriLH0vhX4wHNOLd2gf421jF2/+1JwJ
XL4qPxc/Uj0IJ0EwrHULgCuZhOgycHqU6B5BcQgrV23bEXa5qMHB6IC//FZ+
YjlhmEaXO2X7A/9hm30pFRj9o5JhROy4dM99heygkJTZCz2eyXBii0bw8S4u
249WjpgD9qLHiut39IHLo/pF3zkebUZzsgVZAnmrrks/IqZLOOjKxcikT3rJ
UMftso+tJ/3Msbz+RCMDgnzq1ttrdlJUFDZ3g2EKCd5IWi6FziFQWq8HQUS/
SWwU9eEGw7YacOeIs55J5tKisAsCuswDPt1IfGtO9lMWip7RFhqcP9ftc8mf
VNvj1saFJWeh9MagAm4nhGMLa6TN9J4Y0LZ60tPrYnVJH3y1uru26IvQ38RF
O9lk9MAetRHQzfCQjcOc/fzsOp4GDBmKYHT5JyAF3be7y8RRxub2jrSkQsvm
dVTKfMXqdSEizlLs1MVg0v1vwcd/L5SH0n5IqcnoQXytTbXRRQ1fYMsOonpy
/bwdbEQqasWa2NXUqH3SxYIBU4cF1D7akagklkuC+BPpkpwcpm08k5P1iu9b
8dyc0/oW6jfjT3kXZETiaA89UStlzc3AEgiO/eeyYrbTddxXvHQ+w6GKHe2z
d9INhv/I/e9n21uohf9TNqUyPE7OVxT/JGl/JZmmHEzAielBNtDrfUroWDuk
/YnUIUtAmyPy5x6Nt3VyL1aBTlX/U6oLh3ty5vhx7PYglNXzkVQql4A5l+FC
sxWc+HmWzQQGFTv7n0XkbVUY/HCH+oqN6PMTPkR+OVFQ2tkE5o9fTTif2A7A
U4Fy4hVYM1V/U0t25GyY/nZd41m8hOHb13+WrvpSxV2/n2euN27Ds+EeoWFp
wxV7Zqo9b3HC38L0SW5BG3mXCXpS8cbniUlQr2C1dfOpY6kdAXQMt9QEu+pY
EuPh2vSi81GItByQz3bUQY0udMwxjvUywfJYPTTx5B8H0282/2fwLIsq3i4H
1j+5+6wBKvRiw2bUiW24/OrGhCTxfd3czJOAs215EyJwUm+PpIGf5bR1nWqQ
ZKb14S8Te3JPR6JT6i5+OpIv0RSagbQ7DZqLPfOvBYomD37BXogX9L5p72Do
GVdztuPWiiiLi47zK9sZUGioXlzLrJaJWsbDkYaUVC0GjOwpSAeRELdF583m
fB/yRAW8RclKl8TvYq5ubpYCeNZcW9d8SokSroIzLL91x3ioJ7PyaCE1VNti
iyqvgU3UaoZKQZ+luuKkIuvRlowm1cmwPpM809O0h9+lK5T1AKMqlJnG3CrT
cMvVTOyCmYooQi10NjYidOvUdoNtd6ANre+dJWYyqjO3/9BaFQYx0G3KTMfp
W8ZBBCx8vEQpMGDmLxyz+yi0eeX3iAtU8EG8llyPdnnVF1l/ZxThaGabwID6
yU25Lt3CoGwMS6/ZSX5ympYwvp+O8ZHayDlyT/J0Ltq10ayGlpi4j8YQ0VwO
d2b990KQSLecN+BAcnweElCC0jxQV/mAsOSj54UXcKC9EryPecg5KfpD+92P
Gsv3XdhZLLY984RBW/B66M56ZAKQYwHZp/Ml9UmamSF4hrBNXt1Jd3v0YYLe
lj6BI+rsjwC6krpBJS2MKLu38VBkycD56rMRWsTwCFJCjxXpfDK0dVwPxopj
2FgiKq7hyA4xuO2Nx1YEFHsItsyV9UDkB/9d1O9z3FRg2dj0wiJmFnsrdrOU
4TnsV3thLsml8mCRpj59p8nP1gqKk+FBW4ym736J62pmv8BqGxXJhD7FaDfs
22Ue15cyTznKuz/GuSILxYdg0W4u770vMpH8uMZnCKm7GQYZZ9en/92IBcdd
teLTaqmIw8Iv6WAn/0rXKF1kPw9FJ3++sZsGjJ2AcivhoP7vk3pKbJAOQwVH
GVoEotYnTD0CgEswUivliPRUYIYNv+Nf8A/MUkM/JYrH/Fi/wU1D5rRti0VA
IBMpacaUw6mhjTbzD/iGQ6pb/GuKYw8JKXKT0E4HRDTVO7I/Z/k05NRrfjDu
Nlm4VOcdPzLjH/5eZEakSaiHGymy1lM7ftv/ZFs3aLTB0YNKV54O5j6fXcEq
Jxv890tbbZN+pEogSv864Gg0qX4LyuyN8zsbEn8JqRMz9K2lKwz2Lqcmsirb
MFCadv5vOLaPg0Y1h0zsB9tsScWK/KdWKQszp05G9jvfkO1pP0oZnk0JHyvp
rbeqH/pG6yd5PaBccr8gcgowzyKrmDssiSGlnVZERk6TIa/4HRRrL3Q7+Eqa
Xd8SS3k/hfjZ++tnwFIxJM4WJBe3ZZK7psf2K2tg/yseHu6M9sHg7fsig/s3
QimPcsr82Gc95wOhotMgUmvtUeCwDydPSMik3gruW0xmQNbRT+3S5N08+FWQ
rdDAIgKB4QsPAQMe7rRU18wWemitM81J251ir86wRd3CCu+hBTHj+ITlxhCG
V7mLcOVbTWJl

`pragma protect end_protected
