// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nD1R5N7hoIeZr2nyWdsope+GcH+pWNcH6fvRxgwAe17qgHuY4VMPCkBlJDLe
z/GM50dzubnnL5KSqRRci82jEol8V1FBaCkA5187GiarY0PdpwsrQ7usomlw
1l9HBqmUEwc5vGWg/NdkMKxf400Vs2i8OnTAB3LFvmy5MsTKPFT412UlyRka
LSfYo1ouExcjwPH6daofeS9LpEP2S+ofvS96caR6BlrfET7ujhh8oYO70BbF
uzl4OxaIr9/HP0I3qouaNSXYOwTWkUToavKqkaqKQ5kYJWRH4e48Xfg9BzaT
2Xtp9MjTzKFQoOWWEgeTLgNoUNGXtyu8tPgWEydNYg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eAhTvLx18l7g/OfvDvW/rEwlNZXv7nWTWtGO2su8LdScrDqtteXVEFntm1fi
fS5IKfgUt1gHQ+AE0gYJeJJiSMeGkiXSCaKcWzseVJ83YcecSnQxHd7Sv1Z+
eN7A26NrVaAm5V4tZw+KJqevyd7HHuyBIIhPYjVKdf1x2jnsADQofE4uPGK3
nhn2DDj4Kmsa/Q3Jc+NIEOCWDwvO2+1dUWiNCSfKHRlB965cz4+JwB631o5G
VW9UWCz00efZ01DJVSpZdP4j46OgEK8Y5K5sYs4myT5C34zgCsLMaypDx/1y
4gOrGXCro6Wya1DqQigwLQu7/IZ6muoUmaP+i8WTvA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WXieLSS6QVIyG9+4ml2tyz/E36wCnU1g3YkVB7npQTW2geFIfmuSrI3v6FUz
nObCsPav7RhI7zjKWcooswZW8n+o+ArnonvXKjI5B0Z28/jmV+xRA3/PauCe
vcAReXZ+f9798XnDjJl4vNMmp5TTj6uc577LIqx/sD3bKFcjBOFLPfBxQdFL
jk0ncnO4v7nBxJEVxJozNFZHljjmLcuEzuk5EKTTTzY0+djwPM4PL7IiaLq+
cMz1mt9wUES6V607FKJG/cUesK7Ow9nOLRu+WTBAVcAM9hIFuzPIC+w5ZxpR
mhS/uoGQlGaPJYvXp2UruUrpnkpqQNMTPb5w80sRxw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mo26rxLYlYBdeLcWlXNg9sTMt+VeCIS1ZV7sLAYcCBQfODUPkT/7D9cj6qEM
gWVU4+eZfj8rlmFisLxus8F7X56aALlSmo8zj8Sz3qrmm0FeGMy/GaOBJ9Im
XAanWDYOigvPq/avU/c2Ry8+4slgbQmokeDXsx6IWxB3uOHQhhE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
YuxlgxSCoqXu6Z7o9AunoOENRHgA1UCnra7F9puwh1TvdE1DStSIv8pMF7uQ
XKHZRMReYtHBuFM3xX8xHQlL1ImUprOM9TA8Nx7lC4zE00mtG44Jtxr/YNHE
YUFXWO0VhxP326IhonlKZVtUWv+m+tmDA2OW6YNlP0hE4NRkFWf1XhY9aUB5
f46F15IfvdaKFF2VuVTkrrBnFYxJEDYXGSUk4RQeAM2UgcGYn2d4FV/2I1So
QtTXIvVAPcyxyeCLCVLKJmZcGeCTtBE3CH0f31IPubFMwoDngVIb8buRtnrn
w7dRrGoXtxnLDDCxMN7CEe0pmNpQklCWrj2MnBQMiLEsHCIeZLvpnIWJrYP2
o+t1mwl7PRtyJnP3kP1OhDawjI2c6xJx3G4DA9MBaZDQLiWASDvMexaMU1pr
rrcnb/lzBv4uNQ5//lxL69A3L4KdpjF2RDbS4FTlHrtnrIbmDwcJqm7UkJJL
oOZKbxjRkd+iI3miaSXEa+Z6CkCIRQPF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
s9Xx9fXb+lGvBGYGSjxvxiABtEpa2e+OU4trDJJ/vLmZ/pVQ5w4d4s671yw3
DwsC/CleKrmJyCiwdvtIgA0o4oH16ma0jH1LbVJcz/A3VCAF3mcH+T/Gp9JG
6JPwbFUNNZvnRp084qG2VKcoYus30rHwddkTEInk3OlyCSdoX9Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
frSGigLmTfqM9JdhDwTUaJCP+JVGfY/E90cO+6fH+FbxqBHi4M4wm3NiQxWu
Jx3q5qpks1s0Ky+EnJzT9Q2+lkXG76/AMyfUdslPoJ2WfngI7P9Ph66874d3
ItCUPKI+YuzARka+qTWnOZYCVcReCi1wibPYvWaLz3xQ5DioZ2Y=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10608)
`pragma protect data_block
ETkedp/a4UU+UyZUpznL4cD2GYtnkmsJnOcYK2bFZM7aJxJ6i2wmXgU1GX2I
Znhe9UP4X3pvV/BDL84/dSC9xB7OTnX9dAl3FfwrmqsJGovv9lOLwX44GuNg
NgOdsD83+f6Bx4XYf6Rcc9mhsjs8v8sfpbleN2Y0SHbNzhO40VT1OvHv+kEd
v48ubw6sRW3inOJbhEKW3pL8pPYx0JGDBizwl+P2FGLX30HcpLZvrCUm/ptW
1Ixd9P6mP5ARAge1IFOgjyJ1bCBeN/WvrncNviL9V+oERXkh3pspux1nRqgJ
DZZYJSkd10hYzjrh1m6tIk52CrQk3sMkJR8GgZA0grCXcQCjzSQyUWNzEfkl
JaPNBKd3dQ9iTcsJHFCQx8RSoM6LiCk9qWV82mleYggdKcBHUoOtsD0cVk9b
YTiUtVnQwKHl3e8VT4qFqigTvVPGU8nI3pDQCcvVnjeamAV4UP2EwWL24kVq
e9oeAbh8a08OSpMrO66FNIfNM9kLm7xWin++6MJyYnvYT8mI9pPBkXo1ziIF
xLCabz7U07eBG+xj8qB7SZrtB5FdiUiPM6oxxmh+lLuycfjWomEDYi8+Dgx2
mQSJN7wIfuKzwDxBMCAZk74ZSbxKTKxwVv90g837ELMhHlTidSx4eyqhHMz1
7euVRUFxKhooPm8V/Yr6xSHCZAw8dqai1qw0ZVfLqnqpwhjtPkAWPuzQASls
wOTRNfDLH9zMGajNHTtDtMdpu9DE/jgBpKihoWoZojGJOiuuywwVWf+k5ctd
tLigeHmVXrJx6IZm6EBJVmbWHS/toiMOAcfHzIwm9s5mPz5aTjhipw11AHRT
iqCvr0RnYn4QJVRdRsLFz8gGi/HSQx3Lq3xoLoali4jA1nPYoJX/5OvhQfXA
BZ6W52tc+g8PNl9qWfv8urEGiENZ5ebKiCkx8ib21K3BrlrILlddWgRkDZL3
Xfbt/klSi2+7cwCdvI3PTsf8IfhKLrChAKxYlD34V/YH1RF8D+MlP2wTzFTL
6kZ4Lvcq6VoEm+Nnhc5uZ28FGIJ3hKGKSTc6WDkyD9rSBPRC0qi8ljXkTDrm
bCaTUeUA0Y5NVLNzm1yVSeFiYw00ulk4LqI1017EG46LmuodopF1A/mtVLZB
uT4EayXBQAL8QBiHe1oszoEQmqP2g04sr9wjIqTwTnl0UKAVxV6OYddKoNqw
Xki4B7VWSKbRcDg5KoKEveEPBQK4OC8hD+OGO/+Bq91b+YdRVyvrpKGyHMKu
alzOPEOYTb5ZGORlgjNfwX9T7OQjrR85hdfakILMiPH9DS66/6gK9pqCcbAh
queorQLA+rpCR3SZEEUv/Vz2hfbZ2RJ1G2g4NgN2n8ZJvaghvajkjBGi21ML
lAH3DGcVSqi9L9M22naqf1t7DFYakO2obDqSgz3j1Q+8tj7Tp2CetrcnybJA
Oe3H6ez3j6yT3wHeXnVNiF93Qe0BpW7KcDDIVYQNof0JixaSqQv0tCrG812J
9T+HzpvhhI33zEpFLEluShoKq7dH3JIk/FWci9mnEaretv8cdugNw2IUce2X
dZF1CufTxV3/j+bVF6UjcsuFmJPeSg1Ezs032yRwuu/1oHH1K+R0VYdVro9K
EnnGX8fKNl3f2iWgn9spf4nHEkLZe4Rq434d/Q+W9z69X4BEN0WGNZY6hAIm
wiLuxZOxg2beYEvbq05Sn8GHrUXz+VJMkXGrIYoKoj4dmBmAsawZEzHwNztO
tb4ObAf7A9QnEVLitnear+DuQ1ISPvd+/hAA45Bu5BRS7Y+Q1Y0niT8mdEAi
OBeE0Qj64DoEwHKpH+gxwypH0Ml55m1szVDNnZR6SzA+IbByKguMwRtgWEnP
/o3NSVB1QtaUUGSb3cLQW4miqtOpeQR9ec55+R3Bvp3KRwsVlf/aG3fFBAtB
S2DGxjcvfu+W9RRuNbV6o58yRqVaY2Wfu76OwFxugl81x7V+PUfLGmLNCbQg
9vXuHkBfTTTQI3yLQCi65T7wN69gj1V3K2TfcIvLAPq7iXnMNCLFUGmbrq5k
KwACEVYhRTI3+wrH2DkN3MF5IA6gLLeCXLn1ktpbqgPFNlkD95yBMP/XNBXB
V4/M51/EgSMLvANLqiMlpsGGvxyCGFzDVse3kqgoMzE5nlffdFwjOl60hAq6
EJWuBMmWWUHpUb+fW/lxmXyJJlvH7kfWicOLYaO2oKmdG7L1IMRZuW0vj9F4
wM8a4mLf1vgNOVNxA5s5fxbDg58O+EQNU9AKJJ31csi6peg3aQ0dq4j/ZFNQ
T9GvfhvxhBYSpjr2nBV1MGTaCObUe5ANbzmoylNfuvIseSmhHqzycBEjkbC4
j/JBGXMXwsclMPVcDeVojxMhQwGJbBql+31FK6qTD9IM2LJ3nQJ9VPacvQo2
bOX0QZ3CHZGTLLfnUEaP7C0LRDV5Hadm4SCrmiEwyiWc10ss/worjooBsQO0
KSWif+8plnBHvfUE2xpK8bcXI6wOX432KAnBf6Glnevrmh0rN227XRxkdw7e
9iHtHqOjS5TNupUqrUhYEfw/uv3ETPK7s8vKdSGT5+cY+Tv+1/QQIDlRVFOQ
RwTOc7YXLrAb8Cc7SQdQMz4j+R+qUbrv4Tv5O8cqHpILyy+zCYewOjDUhD9J
JY7d+k65yvvz2Nj7JY/QQjlB1TDlbp1UprNzcFnaLYViwmkfxwl3Qv49WHCr
OshYQI/A19af2XTxYeCRWOC8qoygtJEIZbzBevhaZHNJYQInq3uotplmPfn8
/cOd3zk5xKfT1x4uTd6PJ6cKnRTscGZcUau7ZRaraRIJr2RjZk/meFY3ph5y
Emb2Zdhl6E05e9LIe1c1tOYveklztf51vro+F9WE7TLRx8UwkOj4zP9EeSO1
Z3iuSr6lXeKS9nMQT5PM2AFh1GG11luGhUY1c8daMO6R66H3ZhGD+o3WrmVb
i4h9UZDLHofxsmZWWfMTG4JIqq9TiQZNWPk2X6vFA33ZCF44LXf4t/9tXLh5
PBEO9c73iXrIcmoTtbGFuYtpvu8eGEZ0NmXdOUR0RFQTvFIbP4nJRXbyC78G
M8JnEAcMRN6TgwXu6DUlNij73wDHhLhvpooE+3uqd2IE53iSUFUT1eJ2wOS9
u/Y6UvdZ3ovRg4Pc198FBuFRsZbUn9KWMfwelTG3k5S5/mTzoTY2PqaNQC0B
hVySo5UIqmRNk+Qcym1daNUsY9Hru0llXj+3VU9wtL0etCytfDj6XeP8BhB3
ZHFQpjMFhKXOJHQNpSWlwk4rctoODdHQVr2ZnIHy118YNe09IDNdzDvuF7zW
lZP6SDVELaZVLPVLqzBqYkFelEPrrqA42kNw+H4OiMIORvz7k+GWr0vx2EPA
CsSMMQhaVSG/vnsSGSl1LON+3ZzYnV7BwYqNbtOfv2kbdWtQ4Lqw99VwcNW7
CxQpa1dHJrvzwqmieReizmCuDltY4C6A0U+7IBqYsVgSEdA0kcnh7n3Fq8gH
G+AnDTuJ7rHiSpnO/yLiM1xr5t2oNlveyHKeBGE6TR/MhaVcPC4ZJJY9KR7I
eCHUUHEHNMPTYqGh79iZLgFS7LheYkXpvoDvNv10pe38oXxrBVBDoH2VeBxr
cW2iRYOowXS+hczIIqc482iyRcs/xC968yq4MAK3vdVWRFi/3mjp40NCd25D
tYaYUKVTu+1ePJ9ndSa7xTn2snCT2RvMKvc97XCvTyBpZ8knWH2vTmt+UDMh
ABvKawu/7wQnwsquSbgowKZ8Bi+vw1OKvNZ5y3hmBnn7cPScqVnUCGfkH68y
2kjFPu43CgTkswdE6XY0vDRFvWHy6SdclEkglT9aAOfaRrxpw7HUnmzcmArS
G1B1gQSCUWe33Ozg5D+sFdrfOfoZbSC0y3KQS8L/Lj6GpRDyHWSTihdO1Ier
0QFlaIbVf4IQVTvFwnJEIKra9D6h1Zm9z6tcf/G7OwtlvVbC3G+1O4z0/95F
4zueQ62gHklsiNrXX+RNdJcJZobhRmATI1IyucfTtQFa/G94ZdlEdLhfQs+a
YE3JgsQjh+KiN8V2EsLu9rXexdx0kPNAhVOYMSnVzTuHG4oObkzFLwMlDKpa
Hb1d66o5lKomxbqGITtkjf1w0e++w9lwuksbVH/nyL9xuzJKDOuQyNzj2MBY
HRqgBlvF8W5m8DOX4wIrZ8oelWa4O7Avc7wqSTceASh3V1zfHZxjJj9FT1El
czi4M+HZQ76OoTCSKgb924bV/AFM1DNhpR74Qi0uigikvSLK4fPHimzvKK8h
InNbtQxKz0RxOD+SrAR5Od6ubWKyzhZ6BnNrztY+3qJbIThb1y1UdPzuQgpE
zrcuXUWyo9Hoeg6+BoAnfKaiIn4UhBI451fERlwwYJ5vOn2O2sPDqkbYaUQY
sHn8E+ZnMgSBpklJrbf2gMG/E8C+hNOaHppIYj40Na1JYcBxOtlo6AbdvyQB
hQnFjD47eP6EOkaxe9Sd0qypkv2t1nM+4dlyulfpReHLitzVX+atpJHVOgC0
hT2i7Yhja6QISXHaAJ+U4Ypyx/fk58M+/0KIm8gOaNbcwI9VXRVQ7PZmIph3
UIDfL7Hsjk+h6lYxgYWJRC/cT9zStv6+bZq4GETHWdJqpmEyJRSjP3nYcIZs
Q2wLWJ3riDGuzhBV1vN80Eb9EsHl6B4ggATfxj4/YWhzsNHsrEfY3nfjYq91
xR5fs8puyWKLqm7Yreoe2ox3i9iGCaUoGzQaQd+oVnILV6ba38Tk/qUKnW1W
7qtj/eE8Keav/jYfjt+JMwlBGS7omdG3NMWB/0GQpEZRXngP71XzrXzitlv1
DBlC07UCHIDlsY8+E1fyLgiWnEGVfVRmmUORIGJ5Pt9i59YdMyE2+foWpKA+
ucRrAim4qbyWPFJkcejJsr/tBEd1cUU9Sf2GyzjCtvFOdBGIjdrIEdWGdWw5
+4YuDYbdloKHp9dQsZOP4iARs2+0uLV6g7zBOdKxV3FjTv3nhCWbQyMgwYVi
8L3aEEO1wElJXZRDaXBjTwa+F08fpwG7UbiKAaGX2j21pcabsEgrJbg59iGz
85MtdWnnxixXmUH2VG0hT+wso5HdmZOmJRqgaezOCMq68eoTDS/wg5bbqdlp
m6Sz0tX+tf14tSZDV8cFPfQfzWaPtdfuLVGdrorFxg1+TWenmakXypxL+CfT
H08pY8kJu0VOxnZ/XEYdTVZ3W5oDFKnG90SSERtYAcTopVDxQrkyO74Thoba
o63UskCDghZVyKWk4cyGzEVh1KeQ7GkAhB6L7WJ460yl6yywk3K5IAbiq+qV
HuezNEpBTrfnYmlSpre+9kc4adLbnNhpkbDKwYHyCYxkAXwOoLZ+jVZhofGb
GOH8L/izs4qhYxuy8NaAwwJwAyUYWyVfEZI3Pf6q8w+sOXwSlyXf7+6HwuQY
pvnQIq8c46O+SScxmq34087HdWS9EJW3hD3Di3ECTzqGkev2uqcXKMgtWgIc
IKrRJ/sX5eFyCFKfa2fdrs1eZQOxLttZIWCWwUwThzgcWTsbrQw9F3zj1GbM
o5VpoG/b6Ta8Bkctb6UjwNOpymWbNO4RI0F4QRHi0Tc05LgALfbzHOQUGpZf
u0FQ+8E+v+motwkuJzSTLBUIUn0aF4vJSqjESRx7C2wDHJs2zFfCiA2SLDEK
Ky80HhoYkz1kUKFtEb0BaUeCvmZAQ+xG2Obb1RBLmWHxNkayAcY4YhP02vKo
eQZNVwvVrjtJguu6WXV67pKqPPuWlfuDp83KjnT94oJnbnFADwJMNsYdpOeo
LaQmidcL+Nry36uGGUjz2XOxR+o0ez7/Qv8WWGfOlB1OzWkua9I/1taJPNmB
BacoSKwh9bQNT4YXws/Bbn3dEyzcbjaAtO8uBohpFqNNJLAkSYFooWCleG8m
/mML2/D9Nj/60vSOEhuB88PaZ7BUs8ITfLwGccSvb6BekwCWmYm/7TN0s3G9
7VMpI3vO4x66T1oa2zz2SMFg7GS3gfwMM01S3+uJlEDDLHlCxFEBGkgiAuBd
KGf5hv5GQondxYFtbCOGTkS4aVYy04x58DlsRQmtmqqmKgGFgauaWS4IWBcw
CcuH1vOqgYr9N3fBaDK4qm2BiH85zt9XomDCGK+PDal8AsoMyZ2Q8Wx9YrV9
TuQZtkC+eMmuw76xvhnid6U7BaqgEm1GN7h+Pk+2E5E1bdXmT8jRQyGe4qSX
QNsvAngDriOZM+aiKjUvbnZY2/qa75X0LH0m/Xwncq7SLqtkZJNKA+cE5sv0
6hLJUNpO8F1vCtDo2K7uUrA5XUggFlLDlgTOoa5huZaxCQXgdmB62OByP8Jt
Y1bkmECXvwcWCxgPRiqFxb4dixPSjJpbzOn6Tkqn7RWygzK9ZOuRk5dnEBTZ
uqPFSw8qv9ovb8/IsMFn8rEVVYXnF9bMkcpK9SqdwqpQpzY7VnoL2ejAcMiF
1sthSjJyGGG+/c0sGVmSuCYZm/nmPfKXH95lq6pqOO8zpmlTDNH2V0LJkLKK
uk2V55E2Dotu5twzbKs2vmJqGTo87u1CIm4HUl4p66ddP+bWPHrgyk8vRmvO
LYkM7D4DtPcOD6cC729ga9QW1GeG19APRJ4i5nq8LUhSCTS5zib/PtXkcEXY
YtJKwEmQbIoGZjBmikG5hjg8ihFUgLmpmtEwwYmDlz6eIb7qj/N4OBZf3kQU
i+jKx7TgKX/UHHcNmcjHnoHgLeBCBqWkA+I3gU2qOXuM9mFj50YbwApwsJWI
+fvrvpaVpGHzodQ7q0aQtx9kLiz9rMeIj8Mnk/GLxda2bljdWX0+vpRto/Jw
WRK4UQqe6Ie7quIlyDpYBthLp//Zu86HcrWgKa+P1WMiq936OvvJnaDfoFyI
pNrVrzMzRmeXjeN5aK9y3krTGujxCC5iRR3hH82e0MQV/nZR4BBVBhdOQ8+u
YtQu8FT0+YQcHCDRI13CspD20Cesr7iuz0Dq+/S4DYxHfthwLk0gaojOfSsj
HZ67JRsWOloX4zWdyh6NLtJmucDlzApmkUdTSCj71H3pMV9pG3MDz6fn+Oaf
whWfKkbnHpLcWpXce8b2FWQdZHUPkEQ5BZQabDHxK0dw4snTEbFusABzDj2s
P5bUfs4ab8GU0mI/RrOapYZzn3PF1m49Awt+WUARCTUzgk/TgKifx8Ss4jC2
+Sr1RLKFIwLzYFl5O8ee4Gt6g/Prl0Jovx/G/fz+8QEzNrUxE6LAs3VX08hU
Rip9hzVmFYwfa2s3aIJPhHZlCjBWpGwDa4nRH9C5DjJOrkM1R3+HSYVzz31w
tAfyUwoB/U3M7IMqSLSVOhsUwpL/hJXKkRKclxzFpffnDRs7Y4U8DXJ3N/zk
diz0uyvZ1gQvruqR19LGeNETm5qMkCb5IhS/mqrid1Lvu4SaRawsrkiXekhm
d2Sz/fk+40roFEpeQYUhG4McSbyn8WBC9hx9cx4+ZTZ/kCcVOD67PRzX4fsH
MbSW2sKfmsh8BUUhJ+zA5fGqCdBIA+ZglG90M6quE2PLS4gt+6v0wJUX6x7I
3QobCgpMigbfE876G8fcQ5vLYQT+SYls13SjaD2hhCAaiQkLGn2JeRK5Mifa
z6YOMXP/053jHGzG71Cj6/IDg1Jlzp1eL8GQarbfesJIpiUmRGual0Si88Op
mCNRGwgYLkOAfp3RV7a7V4IaPp5AbxjzUNJ1zPGld0yExgc66m57dN7FByRs
SjBqGGrlk8oFNL0mtmT4xja0bwnB7cV3xtgp3WkuJF7d7JfoZK4kVRcHpIMu
isRdtwS13221jR1+5i7NZn9/bv3W7oUsdcPQaP7+V267JJ9JKHuD9ATZluA+
DMOYklAKU7pghRH71ST+86du68dUTCiRYFOR/CKLp46hew9scoTxD9OH9q73
jACdzvRNA80R8Ovfb5ieKWo3RvBqeNGYpQ+vFfGrX95ZkOzXyp8gUjKeiSNv
dm7vBs0Q1mTfM0xtkybChoFZx+ANrN2cSvlnjm3eXjRjpUDfmSdbWv/I03da
Jp92etU/JCyWGqno7s4Q0YyK6NAQ9pq6mWIscB5aBj8MfSZH/V1zE4NDufhD
UnbF8517ohs7Kf1IPoKJ6N7i+eoLGhJL464hw/WhF47UVJuKt6vSdmbiqzTn
NSFcIprhHWS3oGuw7g6CZhNGD9yxOdaSuNysTBcLFC5TnyZKt3ZhydGP8DK0
2UOW/XkGR33Zfmgy2SUVB2TFmDpybognDVNxeIKzUz+z8gZPneWMiBhDrhgx
Pi+gx7M0jQ14YyMyVrlY2hNjhJimml87P+oxtKvVRQpTitXh3OYCWUbNADTn
YVSxO+il7Pai1VWNRC2C1vsFiTqPhTTDj5iMMmn8tqPmBWbTlGE7NWUUoDwO
L07hibwEaodrHjcfpBdzzrJroogFEyNt9UXS2SKBx+Jg01hmtztaStSKTg2d
2e26F2d6gttOou3uUQZMDXyqyGr+DOTFzb+6WuzflL6EtmQGlg3+Wp/mvmE5
EQqVAw+ILc0xaNDEw26NXxtWdjL/qDu5Qc521RrTls2jF1ZMaLZYUYuSBCSx
IDpmqLwZQsr5SJS5+ROI3YGMRGGX9vb3nkB5ZYwt798as2644W2w3FtLdS9X
NZqHyzCE9GzoV0vhCaxlGeCpQYo/Q2tv+dk21OO6MLsxSQCvU7gqKRf/zz7L
NwW0Cs+PCnMjzO2alPp5SgbYAZYZKzmrTkT54SqcX1XR+/S/HPScO/5pTRtU
W1CZq0QOzDrJ1YLJC7UFqhZ3mAnTSeDAxNHEwnoI+yaOB2imDt9dcE37YVbE
/xemlvaaC3NQjm0CgnxqIKD4VxpuAyYxeEcfcuQpkOZI6hPP1J3o4I5S7mpV
wwbmMNZWqpFR7V/zysidQAI89A+eK5rkFzvw4D46xyMqjB9S+r4PEbiFLp55
4IJ4bgeS1xBl7ItzwEXPud1R572Xdn/rQU6WpAuekURPBegwGr+2wNqbmA9a
CqGCy10ZbeY9pVCil9pYCI50TQkPmrkvYiWyIvjSzZ/B4vWKrRh0qXACUaLt
f+cChUPvP9BJ/eCJgh5OMs9SQPfqvRN7qiel1pyBHfvpcECBqZn9/XZP9TMw
Mx97oX/d13q78r7KJ5RfcnVhqElrbKkGc2nc63kphLFr9oszM0jHUs9RptEK
Mvjppap1R/rnmbap+1XVW2n0Rxjy/phcrh2jo5ZIE24yXLYcDHYkvSGVhOsu
VK3ltI4mDioMyCD+WTviCONOoK6M/xF2vQtGZgUEABDWikGUZU+Vsk0mPKQi
546bu5cWjOMANI1nZjs9ZBD0+c87Ic+jZ2ATfvhqIsCbb2DVE6pI0iyJWMxP
Ufi3bJRZwRZAHPK07LmsFPdhorx0aWwcxa5WG+4fCaI+onmXy2lhYSrS0ju8
WdTX3c3sP64c6gLUTTjPteW/39cfP/wJbIY91+KytkQYKEzk9DNLE/YdYBw2
xoayGZJzXkTCKVay408an7X/16eAuGwWjey/RHjdFoZ7RnriTdYCjG2AvV4S
1EqM+iAWBtpovMTBwKwzWszJcMcCDajcv4ZcYQXRFAq8uVnL+t4FRYQ94jOs
pWBNEeObenpFc1kGAN98B7Q+NnBR2y++f1zvhiUA+mRyC/NjkVN0U6RsZbk+
MBFPvLk9OV53o5ZFks9KdUEUP0YO/q5rJl8nXsqkZPg0QXzUVb4//mSvHVhV
pWWef8ibNYlZv9tnm9/3PXPKgPrZm5Od2xA1qkFi63KQ3y88X8fhnraPHnlA
yQPKcS3jw9k0BsT6jQdWTiHVMqwDaUk1ZACo5W4Mn4NbZF2TeojUOsl5mueY
Pd4oJ5Yhqo5hjxFgMM8hMJTEeDlU3y0JYwmJBjY6rjTqzVls31djYOzTUhcl
Kq67h3iaFw3fuuRLMfr9z3VNQoIsy6lKYF8HCT93hG9WLvCL3RM3YZvNyt10
4AwgOkeqjDn2vIkz5XdWC8Q3aESA+YtC2RfuHBce54MP+RsPMIOJaiJx2r92
tpIm9MdNmQcY9N5MtNnFa6oylHf2xg1WIBhtS1SQBY3g1gFlkSbJHLHXEBY5
hafOKlqTOpHIWpsmRXuaE5HlR+2ateje+qcEfTeOZeiCKAJqgR6P4QKvixXp
zPXPu+lHlDCe6PAnlnBSkLNv4esa3Bv2RSC5g9ObSg1e+2Hmt2aNS3C4z5yi
cNp5B1Qg8pIr7uatd8XHAww+A8y4kjBqSGMfNeqQO+Q6z58beumHhXoJYrDP
idkjpgk8ByWPxEpl1AinYwFMUN8ieIpoA7iDxeBeROhe34Me7isj7XdauxSo
/BwhPViiccCPRrDN0RqxI4vUA4/XGvhQfgRGrdZa5MlLrmBBFhn7PKLffdw4
eMofbNBAIF6x1uc50xVKOBw0TPxSpc68GfF/QHMHcydDXow/MdxtAdOltNLD
WW12KRODRm8yoSIAIwsBiBQLV96jR53f/EBE9Ysdd0SoCgDXlcWsoPwWvMwk
A8xJxDENXpbgmxIFyuznZKpSNH1aP7BvEew/Sxx4Mx/EeTqjT7mdwOW843bp
xNyUcIPo+Z3JCTBz5pSE2jJSjhFPpc/fVl0cwiUjir9CQv4RZNI7UitLWQvo
AUDj6LfQovaK9M3C1JOjc52LuX6KHyFIsD91lMkQ12UkCEOaYcB379Bi3SwL
v1XjB8IkbEh+BCW1OUYwqJVtkMeCLdJt0Dm2PXU1l6nnX7sd//Tv/hZk7xme
j6rzviO2KCEwucayf7B6Rjt9I+DEOLPnQwtjg+uYXHotmD3SY8YWY6ivQwH2
8hOQ0moWAWl+8YUNJXTttGss3+83Yt8qvLbYR9BVr5cIZuWzswLsBiEE1uZt
KuXnQ4tsVeH6UgVc8uI9HjjtU5dE7tO/5sQo1LHKWGrs09mLBIfjIDvkOJKC
y7yBOe9ribQ8/8f5DhEnlVV8lJi0alYxd8jl77bWzEQBbzR5UZfY3SHURg6R
k96XrkJKm4FYePFvTfbiIvZ7HkBV25rbJh1UIMfxt+Euupeo5CSMaPchKLpN
wVpX+IIVr6I+gBY3argjBB+nYiraILxf2Dk80rjPkv3Ja+/HRKMb8u5c8PtW
xQLYryc+LSkeUdVpyFjWAqJeph/+oWJTN3ZErV2KYYFR02TD5U8ANESBuW1+
qFA9jVkX67/vs+KveOhRXSu/8aSUBI5YuxPO+3FY1nieOdX0CxKUYmhlripb
6RATH8vq2vm3bL1/OMR5V2YZ/e0h2OfOvwGLvTWoAYNLm5MusmEC6HU1VgYL
e/rGOKv00ZEyTnGetewSiy1UCbhcaZGl5dHY2G775R32SV77e18ksLpnoVOp
NikbrbMMVgcHKP2+GPALpwBkL6CzhONxqkzVpv8edGqYCe6LNhgrLFATO5GA
Ax7jSzw4Og/w58kvFEadvdSTfjhZbCjwtmW3et0OzUGB/mQyVasBoh1phJ8W
CIuHvk+3Q19zQtFsPxj0i38goaJxIh1uSYxAiJjPtWX67RidteUPEHC94gae
oM1QkOplewk1hr5Hg6ojNuxlmL5TYUgSCgn5hfged3CKwsr1ZYP1E6YaH7UT
UGs1JjWAHgSCKF3X3LRJG59/X5myhhaN3NC+Mq15PrcY5FwN5RT5U4HxlGeX
N5U2FhVk1rdpj39ZkK0PTDSMmIih1eejfMUDK9g8SWLddDeKl78TujriU18H
+9R3vGsrFauAAM5LpIgGHuMvFKM4X8L84+r0eq/LYi9gRXvWWMp93a4xuDqC
HgjdEc5X8wPWMO8PWkcvdSlZ2DimXy7CAlragTH00tpinZQfuGpFGhEuoOXD
smYC32ATkWyYkEs8oXRrrdtjW86i4XjdafREqKQWeSjKdHD3ts0iFNmLnIuA
7BUJZjka00RCDBToYHjkajCPmqsDOYWIjYM7Su2+r7UAlPMfisnnfaLH8kQ8
R7B4ypyWlMSM8fVLJsx7bffHXWcBimP+8s97v6+94OOPCgoq0/QjHlfNueim
f+JPD0X1opWmytsaO6fmjgWbqbNCYKlTWb6jxO0DN+Y/7RWWBA1dC2NuEQ+i
QhEH0xVuSmGLyItIfZGyiNY7C29wepM9ajn8O/66NcmT2/nsvFKyPV/nQXrq
Es0wax+emSTXny76osuNp+oJGSN/3K0jqt3G7MvHdy9pYM2igvJPBingIWqV
glS2tI7+jDWDXGu6maEybhVaDMPiekzzRgz40Q2D7+yfTvwRUwehVhNJUwy0
OhBR1Sh8j0QD5w2ONtR8xpAAzXuH27v+Tp12pptAp0gLO5eiXDRXZB41aDys
79lx63NBEcTbVsinZfbCQqhWQldLWolvZs3hf7L3N8g+3FxXj/MFrlYBN8uZ
Z9YAa7RLjmtUpJwKMVrDzXC96jnClY0OhYFRKXRRLZYC+l8Nqhrj0/CxkxSQ
IE9/w02VGjbx0qxuFspBqpc/JxHW0TR3OxG5xurY/+XJRph5Eh8Jm1Hdd7IM
i3rXkLbQ1b3UoCMbNmO8VEP/jLx+KDv557LuLhI5pJnS6QqTaUH1XDMFyN80
UrsQLGaDS8+goWTsxW6t6Z/Ajn69NcyUu+xws9RiRHZruMzIBCRxcTPl3+QS
NrO3ItZVXmxZeFTFMGYClkK/Zs+MnYCGK+FqbXUzgCMS6eYp4cNrxIvVI8kG
UtI5l3xr1jCxBT+UroqzWUpCq7+yJYE0XZ2tImBdGWK00fdbpad6qgiV3Hcn
YlDL5xcTDHMqZgWI1IzAVQ55p2KzlFfsevwp94p/kpZCjowoqS14KTrTeA08
nhsV69A7T4n+xVTAg3cUm6AabUEVGIsE/XVX8FlduTuYXNzYWmjVrXchS2T8
kornLwE2hbydkcVj/VeZ6fyo+tYNWj2OkAa/ZSE2PtxNHIcefeCxpgELl9lV
cRBeJt0gwAj7LTdrF+Gejp8A9BOCBhewYXyDn2XphRQZhvv0eHrRTGJ8PyRd
4nkE+6/UGexzYMs0kOuCX3W8Bdq9unasUZgRTINh/6e8T4h6LNauoWwo4S0J
LKF/OjIMYi0C9BK1aLgUwVdgynX9CkKG3RhMfHEGFHgBvz5UnaiEUtgvhkOq
J1La8mEX1j/T3l3FmF+6J6yD+3exi2M4wjVSGkID2kVvSrRFqGbro3L1BaIA
iQyuNQPGfhloJHAyef1iXrlcNuPb3I+k4nRF8KHHDi7DFxQN9UWHIuJBc4TC
tigSTjmjrAEWfYt9SCaBF2td1nJ1Nz5G2kdCmYafluPCT7cdPiByYFn2FUiV
xMx5Ty9sfSvzcB4CaVUAH17MCBHK6UX2tm2vlrACMvt4N56hd3E8DkPG9enN
IsWWS2fH3oc+bbKrKswBmYkxUL94EZriykXgQdHCxaTifq9ydd39a7jdGA/4
EOs/x9BYulTYssRH+3ES6IY3AKzFK/279L1z1XtIC4j4PLMugiUT7/rkvUYz
ZgL4XEz90eVrDRZDricXoHC4LBiuYnhEMpyylDM39SO1m78DguXsMdwoVrRO
mNwm/R6cYgnQ5p/e/1W6Fj6iBY+KC0D5PI+fy/YAM+CQY911Q4pyeh5Du/8P
wFKtsAmnPdgGDJqep9yHwWK5iLLYQvRRLy4n9d1LTxpCQ8obmMzE7NN+gpaP
xnSNI8te5EknhSl6THB5OR2UnX0nAtsNwEM8NBsbnLRxGjntWpHBRL/t660K
BljgQI7PPfKWYSiR3YAXFdxCqlrNT8wPMlwyKZxMu/xgIMGofoINpQRW0LbO
2G8T75X3RXx+IBS3XBMrLTMEYVYp/zRUZdG4iROSAPiIoh9oUrGsV41w8tcD
FxX1RredRUhg4zaNXPVpqHUpgJMXKJZ02RqbaXm5Q5WpjvSdhQbcyG6OqC5U
HJ/NOPn0TIC7F1jLBON2ZEr2jwIvyeJg67bGHzw1pHMN1JS37FhoU0qj0orE
VZI19I4FSqoZsG/SFR6H0nLUcYaGz+ExDgsYgOuNgKJ6g23jl/Iot8nutLJQ
9qrsWM9uJsEva8DSMdHGJZvMrYDlwQaBY1b+E9cup2kFl2SCBAwmDGavgEMu
vAejUDRvHiMg4xlR1Bb3EVPdeTgSyuClGXGtsIfzZf+lgEBOiqP2RP4IJFG+
2mFxoLHpqbFhYruZSkufY3xSVlP+Hxj2y6JstnBQgSMplt3Eap5qHYcxkOZM
r5R+1qGPTrfravbrtvWFCNMt8Ftv6F4sz1kkDNCK9S6Z

`pragma protect end_protected
