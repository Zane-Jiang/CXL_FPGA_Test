// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cNoFY+9CtZJHajTNnX5ixvFLjv03QNisIOqpsg+SH8ZOU/sSiPzO6IBMlh+u
Y1xcGQ+rW1HFc7luFDkV4BZhiOgl5qI7xwTYy+VV5xFf42HyTP58JJjs/2nt
Eqycw1hm5et5nGaKj/stB5yeFHrIgaSuZ6hmzRkV1nB6GGZKyeyQmoC4azOy
GZNvxFG4pqWYCjYKw7zvvLJDY0CHGaEDMFLd/ldq3xoOuL4ip3mq04oH0c+Z
EFbr3KNjPOSBiakxYS40X8RVd59VI+zf76EeiOT1Oic4VX3ZWLIt+j2jbdpO
afG7cF6e+0ETcbSoycjzfKzjmcsyttP1hBv3V1B7/Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mXrW8w9Qym96ZPRxJJw5A79NlcIzqZeZ4E517xNVn4a1ZQvcRz8kFLFlE2cn
TE8tDpkfsVrw8U7Fomz8MNwQn3LMwGdCOJry36WaNMZeL3GAFA9kRPYHlXPN
YpTIAtOvfi3ZT85jgo4GG3SV+7loiLoRSaxMWxWJYeTZn5tb4T0FVzc9JFbc
X3Gt2ICHXkg7jGjpY3l683ZeN8Ej7zigWLyBvVACEIzkSKa/zPmxfIcueGZd
OcgX1ByvkrAxgsuI2AykkwfAzlrlVLM+luSnX21HKtav4UKw+gQp5z6ngWSH
1H8kRdB1FSFtyk3Fx1ciKQlrYI0on5Lun6wehvpVbw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RR/Pl/zTk2Nal01Zv+g+Am0jGZ1MBX5rjgnDAsoA9G2fdcIg8O3oT2MiGbFd
k2zPJZ/HADbDnqKLbqz3Yqp6qBTsOetkGuVg52NC4hey+3X95MevHfBgkZiX
h/TFWTMbsH+hTv/mbpb+a/5enSPLpQBCT7SBbdiSH0w/KN/GuTkTcTDwUfkD
C0Asvpb6BYVqqUb5OTpm5o91g+7wh8UHyEOMxQZnm5g3nn0ATSWteVM3rbF6
tHCkaFrzJ3C2p2IfS4Wte5s+jex85nfYceTxs/3gymIElqyb6V3Di3G7406L
l36/zXkcxNm96dV4RSXOEjugvYgMcnUoKNFcA34BVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lcuXkr4UU4ok3mvcPlI63vM3cZz50DvNUdlO/Z7fQBkFlh4LfbozHdAa0/OI
Ior1drqd49F94f0Hk41p0I9oQ9h/vYqhMUdv8/Oo+ditMZ72X6cegBfj0puc
Vqcpb1fO5XKYrpyKPJlEgo67odd6M6kcitc6PbEsmXBitcROsz8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KnKc00YdNJ6quM6UUltAQPM2MfZUKSdInQBQPPXcfE2bBkRWTUEPLxhJKpLe
XyqX6LMWfv1zX9N7+LdIOa/UB6PReXdahn9AAOPaSQp0mBSJBcywV9s11JBX
7VfqzV9c+9dd5X/m9lCsZZwYSJOrKgoetwlXCNMncUXYD3lMn77VyDqftKuy
fZyzhBQy30MNgsa/0GrATSTqtBc+aAXoRkZgNJ7YB2zeesHTLQ/31vwmKGzw
xGbPVo3p++L3svILBLwr8JRWIDzzFneJaVvm42nGMSWLxZtg3Y1f60Tijfig
iFP0vSfiJ+DSE1B2+0iklxnMU91eejdSfO/RX894NE8W6/r9LKXixMJVRuB7
eGoZ4Lqq7A6GFunq2VuUG8o6Nd8muZn7bB14SqsahmFjbcVI6O7QR7Dw69xY
ogCizgU3JLrt2M0l8LSb3unmUyA/pnrSqqLFGNfkl+N8JQK7I7mIK9Jz1ST6
3W4XOXOo0QrgsFMGKm7Ut7UDWgCQ+NW/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fxqaImqYzDiTf3XOv7DAEa4xrqDGbTba4rIejr0aESohUjoivNSmmX2afT4r
r0DN54VprIfU8Pic/iugrnaMiHnA9xRYx/nBFXGEL6d/MzVUqv0mTV7v74WU
CalsvU6lbgGZXHYA2//EGjsNXCzaO4N0xUPZ0bO06uxBZqaeWII=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SzWfDN9NPNAWVRFrBr1VuIgdcjqwDh4YUFMFF5Vz4CgFZal9xd++2TrJhHU9
h52txOtAFDoHEu/ahAGy5qh++RU6BUbjAntlQ/UkTNQe83wsTu90balV6aRx
WklUQBAAg7h0FdQJmyYPiis6yiCR9gXa+fvaEKsFGCJA7A3AgcQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 65472)
`pragma protect data_block
EZUL1uCDmr0ns1yzy0fZmdCwmBF0uKgQXlWPLd1qriKbmygRM/Jb0eFiKMjq
UJmfbrBiq4iH5qT+k6cScZSiJleUSch9LdZ3M0p+0xKES+PGyZEkbQ198xSF
IlBOGDlIBSkCHG1RtWemnWwp7UOnaM20GXfj0ih0BzZg12nB0kM/RJWXe6zZ
EHFqSO0heM5dHNP/Eo71ciIlWl/0ZKHo+Gyvc0Y9JulNNZssKRPw8qaA4c0Y
lhBHc+F5/FxsVI8nS7bJ551v3NjQYG4rCpa0AZi/RPC9qwcZToMFILEfESmb
RhxWX8avBXFFN+tQbdVNIy/FrNXZm3BgxWhKI4Zs/06/0oYUudAqtnM627aZ
NfDhktAAEJbUQ30REpXrcspr4+lXNhpxcK/uFtGik6GRUDJAOzfIn6m2frYa
qaRgeqdDSSD1/jFC9Mjh2yriyyJGci3ZyxdhhFD6pk3dUTUQiW8BtVxE1H98
vHbxt43H4lSyQnu6ph1yRSwwU7IcYlQrUlgZ5tEiQPOboYiPxXKX3W0RVF9J
hSFPvLKYPlsjhvaXH9WXSAfCfT5zIL0j9Z7Lx88muJl9fS9i5E2ecGlvbcC5
BLWh9QRNMPWYMRuCNvs9DS0P7xsKmEyMCZA8hIKMd3UMbtf2wYG9kJEkl4N2
o+TT0if8jOcOCQw2GTFfTOoOKty20mpVTKt1sgLBXYbbXC+k7VlzVdl2Bw6e
DGr8OCCU6LR80yTy1Av4icsE2pxa9ukMWAv57RYflqVvosKELLfDBfOzWj1A
KMmT/Phx1mOf56jUUdKbW4MZCCgeIBACQPVEBKAiGhG9z2F+kREyRW+IvrlS
+fPhAC1Re6J3L8FHVywNRJ2kspAW0ZP0Kpq/lWWgIdH+l2GxpxUjcRjPXesv
osMd5JxbOs3TmtoADsp2WLuYzonhc/hL45+kQuia9cSvzwZ8FOQpKTK31itW
4iYZVo4IiFzvnkOFO1znK1rTMParUjf5U7hhy3mlhdmcDR8dtUZ7l4g3T1QU
pE6rP4MRMO0hLfkjRnj0HoBQzX8onkH8aLCIjLgRPRsRjmzLk/Gd2Zxu1/9G
ndxh8Hd4OOOH3eSvyuCaRaVjs8Fo7rJW1pq1evBjyl1cB3asQS1q/FjJaVFr
jX/JmzSaOl93fZmF0byihAfOzDZhNMD4WnezqIwWYHilgvI5tP1+zY0IJaah
CkK7dq68egVks5y0B8Yab5camOcr3sa5TTXF9bMZ/CsU14ZLQf2crYnRnaKQ
ZOxwmVbF4hmZSZctJzNO9U7Ck6s4uwKmsfGvTHtpO3IRvQJLT8TJmheS5Y0w
R4AG/BI1WSx3p2QVg6MFsfe6SYQolScx4dP2NaohXXcrcrmc9A6rTZrvF+SJ
fXVa/COND+vNeN4uxyUp1PC8Dr6DbL1HkSjVnjeW5GOej7U4P27dXmYFpbjj
XX9vxOn3Waq08wRMR0Ye5PMz3Gx4x1xHt21L11XhUTZwe7i2jK6rzzJY0xKU
6DjHn9/h7cm4CvfN3KhLaDbcFYeEi4eCGRocAh0ADhSvNmP4EIEEjfm8N26C
dssE/QGJH3fzvUp/zrmEKuUSnHQ+TLoaTvliaAncZhFA3uTPQCgX6S1YENa9
F90wzTLDk3DpnrNQyfwLMOF5e2hWDdF8Vk7X/5l9OR/tM+qd0OwsWxx4fwyS
dzPXjT/pmKt6wFASAhA/xDeIjfnE1gbKlSebmRqQ99UZU2Tth9+zdq8TI8a9
SQuz1qZmb5MWqS+HwuOc7zd+mLcoJH0YVTmitS2D7U/UkIVvoz/sBS880Il4
wrs/2x1BpA9H7LypcbTQ6hHErLq1RrP80F2KZ/rIbr3jRv1icjcvNWhRGuYk
rzUzlD8EiX/aDtSlek8zFIUzley0AfyNRYA4lGkrvuLg9iKj6lBJCeGUmv/P
Kqz5xSQE9uH0+FUsUL4KFbzivvs4ptAXLdsQ2GWADJ24T4A7EHWcNnQsKqF7
XHVoXC7KTk6GD/rSxmNvsBjARpi1bCEEnxAU7GXwckgw0Euckt0L+6hqE0Gh
fkkJGGoByYxfHv4FvFd/yUDHf4OD2aZNO6D5dATTO/QtvxiChpuA7JmG80DJ
fWkFhnau77yW3CFt7mnWsfzSAhddfXeNc66mDOrisZfsF1KfKFjqw3yO07Nc
k5A5fD0JDfZUNtVPVM0CQ5KlX3YAbF4fPNa7bIWL22pq9TbPCVihWH06AlFe
CQsMZtZ559sIwGKK3ELAHLGOVl40SDcTxriSe+Hu6rf4E2JC7wKF2JZPU2A0
3jpy9ITIO/aiZT4XX2jRHCbTVRJ0VDW4JyFTBi/m6txzPIsPfn3OOIi61rzE
HZT8IDboWzWnqHnyM+u1R3TMMr0/6jzCbzN6gKVj1NbOUT9296az28U/IAZk
RjNv4l8WVuY9tUFlt53wDpbCC/pM3pjOg8bGxzHrTjeTI6Yz4n9ys/Jyt7U4
Bqw/AUuO+5SPM+ma268I6VrQ6x4y64VxviDrttcuBaGeoL0/6zY/Xc1me1WR
8hOGNkhdwBGWgjegjrFV0lexQBCL6mQypIc4qXDn4/IVm+B233VtjhpS0S2t
JbzahpXBHNiF/3O9i+CiB08YD4eng27ogjlbYSM3yc2/6IxiEi6ai7NUfn6Q
c8Ytq1TNSm9pDSnjSZmf3IAv0+5HMrLGsj3mquyNpVXpk418U3/10oCnlUhe
Evqpkhqccbgn4t0khj0w9Xn5EeqVCA/aHF97Tpud/2yOTsyjbs57EBNDqgPp
IE7ak5ZOJm8XEgzKJ9PgNATHPfrV1N+LOuxXWoODoATyIG8ve5wdP+l8fOmH
PU6XW6eEVpzB+qpHrIq9ZT7hctOUcwhpBoqx1gPtAOhMbgn0Ym5okXDeZt3w
MpolFzrJGpYqlj8HbUzcgDWjUmfJg49q/hJPT0xf9VHkvFM4d4kscM+hDXxn
a+m5Co3lPLNDg+opdzFK6XwIeiMxMOeqCtVxbmQdjsOxfNljzz+9vWyspSA7
MGREmcX9PYz6igctOHAVC9Z2K61JmiPCMN7eS8FfNt6AvZTks0lHv6LrvuQ/
9xj2Cu0ZUniPTL7nbaWDyogo4LaXT/KKkxZVPcl3AzwnM3b0A6gYB6HMUZcA
k9usmxRV4qkvJSfV89s35KK0XslcLv943QdiDucR8+Am1mBu5rEx65YA0LiC
QV5hE137TG5nHSL1He9J/qNqe+xLIg1veti+teCYtmtNdtt/1PHZOYd7YnsK
NTFaAo/T7OPfzNPPgDd4hvF4kUjm3Lp3kLsYrhux4LWzcv207rv0D15wE8o+
Mu4L1ds0OA2gjfew1zmVxp/6+yJvCs2Mtm+r7D9prKalYI20mvmxDxVHAz6M
eMV2pTKamoH/CU5RFCLNYDZQWtl4tYiy6GKeyAg6BEaf/LYUVuZNGnt5tjBj
oxFdhqGGl0L79wYsIdhqJSFJE8SZxd3zCG+tw9KMwG6l6m9AAFpHFCMH6GLO
OZ0SjPBk5zDfQbtg2WFBK1nNp3tNoZIgyp6UT9zZNWUB7R4ag0v19qT/M0LY
tHFBGyeMubcXO8e5RueAXIbfjYMpELxphv8YylX4HV+a0NijVFENtSqumtQ7
gzCF4fvoOQd0zUsno+2XJFfVbXTRIXAPUZN34ToN8tLMIojmv+WqXVvNdwZF
B0QhvDqab/ZAJjmPpDC3avWjxtOpIcCnyhWkyNn1i3HCsJa+uCEsjfE1OBro
VYba/wrswAu0ZSEYeEwOBmCdL0i6SQ1uyCJ0ox7Yicfl312UCl5fSl+NZ6ek
XvQQrQ/fxmTs9sefsDiX0J2VXztd9UysHHCPVV1NHyLLnsyBfR8X+szG9DIE
JxB4DEnDo2NVlwq+EVgjJegS9RSDq0I+UlZO714u/EqxDIOBIzigva1V2oCe
J9SkKuQaHqDiU375hrEcKv7wvdEFGRJW7X9VKap4FB7YYJoX8FlHSfmDIiQC
7/45Bmsrg7iKNohkW3iTG+SllTVJLlwlDD0ZBhwx4XoJ7IM9Y8zs3+P0628B
CBiuzFPzvIIrg6FhGRfFQcimwGtINLD44yHIJXMdy5WZwSi1OqUT4dkPjIam
jrRFnwM/wLdF+XABTm6wnNSSeWgfhT30AgedZ8fb2bsuVHuQZMJB7Xx1clSX
NZIZdmfI3RWvI+1kge9kKWMda8eWEiPLZ4tnlSqqcj2gCR7So51EcXCgATrO
a8hxP4ftUx3CPgsuAoU6cPiDGG0/T2lNzW+JrgZieAZCsp9HNZGnMJoxdM+a
zUtEXRN9N1JesQKuoKfXZwcE4BwdWVrJ8A/iaJ5yE740OuQCVbWx4+YzTMmt
+GCTWhZwWPzlQdtPVDcUbzvLIt4G3vZcN9l0aFJ2OPSmujiiYuxyHpUvh4IS
i+EgEIV/nUmm6eezvGgla59rn1b6Zh0AXmQG43I/eLBJmn/UJevXwkIsxWIP
JJpxLKwBN5VXa70IKOynNLphWtra+YxUEZsEo3cFM0WoPPeoAJHq1dg9iL2t
zxZaqKFg2/iVsW8ToUW+3pXBdciN5a4ma20ULur+fLph8MbS6mwIaAhvwEcJ
oKj+BeRnOk/FqJb1j1Ae2q+BbmrlwfGsUxgoxoVcDJM80jPudH/Uechh9hOm
k8SAxHThhAHYUnEsqzPQ089CEqQ1K5uTHDDrSepfHC1wH1NlwCUIwGLQpL/P
0+30dd9ax+8Hbd7+wzwKMYaC3onziPb8am4hjFPfCxDxic+uGyZp/QrCZP5O
X3htEMu2smVMREw/NGf837p25USeuz6Kl9ff6NHNz/p5ia1LLmp4YV5s0xEo
DOWy8A/zAeIRUPp91dQHiDnmGF9lK/dlGYxG9W8ki3f6qKyCtuNo5f4ZGyit
Pp5Ge68kw1inMBR7PIMbB8VwF/DInyNcOvYjMDJRDXZHfZQDO/gALsC8us6q
pUjxERyBIyACX/PWFIEhmPczF97cyuy05Un/TJydV/PehL4UcRfzhWSghAXd
DHPREz91i8O0X+beFWrhUirgtH8P7hthAzWsBeZuFXIxOaggfJL8K8R+e7aH
8fV90Jojo9XHeGcSBi2cff3TDm7M1DLlPI/LxAL3nqwlGXoUzwT05iEchAv8
WNJZMl/HTgDkBU859tera2ZHlvJgVk+KEj9DQ5VfoBYnupJIS6nPwhn8ucI3
Fp4uPyf2HEgkpRYSifu+R1pR/st/OWPCYcThrfBibyZ7kFyFwTxuZtdBnPs7
n0MkBt3FUhSUr4+umyefuZ2oHDvHGvqioUE56H4AW3Or/YjQUu/5ylkJQxkI
flLkdwIq+gcGoFXRf/w5b+0O+os6D0RcWKNeno3XG3rhiVcuhQxC20rrd8j+
7IH/e1jpzbr/wLS+LwSe7KcbJ1WLXFSVXOvK4l+7j7LJqp9yrFzvVyurNDTs
eTX0EmYXvccx5FTrgKzbq8MfjSBe9sxJi2YbI4qqESPdUXCKXQJcJ5EZPHHF
+td8tAK84ad29YV7ZfivN9B40IwqSQMaB92hNYt5i6+VJwYAU500JEv20o0B
AnYmombNrm1dHiSD8kAZ92InDjmYngOCyBBlqYWcjA1nC/gG5bzyFZXiPTNi
vW9+OXkvtYCmS2PLw0YagZY2L/8HTrGzVCsvjwBex/mC3RSFhJYGj7xzXa4J
FxcB/RhTURho+l8MSd7LiwMSB7DFL8wAjhho9fSa48Rmq1VPZUst1vmDDdNG
Twj22qc7vslWythjGclQ9ac2ClXgJnBCLjEJ/DS/kEXRkd8R6DLlDJm3DZEm
VSRCIqObwd7703xWynUOGvhMrTmAbtYYGlmDGopkszsx/QWP2Jxpvjx4uJ6p
hbcMqHVGSZFG6gHDmU7us3C5U7P+CQuIqn8vSBGMrOGzQwnNfFk4dBjBCJAc
WMKbOuytki51XbfsNMaji/jkN850l86KkayYkgWQp2GsyAaxt2Oyb8QrhJJ7
24lf8CWpe2Sj2Kef6ClR/rOPhq9tsjg0PsdP4pgP03fNw37Md8F/c49NWGeb
6Lz6bKUahFEDjf9SiOXFiCkCzO3nMK1ddOADBwf6TxRW4Ek4wItUe/EUla/n
xSglcnK6skIj0IFtOZSpRE9EOr+URMYngO/8vOUhQfBdhciAmLvcxbd48nSh
/HBs1UAt3I2niDfYFOTFuZy2wR2S2d+qtfRhCR6UKEsdSiFbmMKniA/ecAi/
9eSGCXb/2adRREOMM7bEYpMQAlnkThNPI8RYgrLX6jLLmU5M3/rquGVi+g19
v+yxKRg+oVTLRbnX1s4PafCWo0SakLEEeaZ1G4kw5X6zwMppz75Hw5kOghFI
l3YNrMkIFzz4XxbZEMUlE2O9KkdQaBn2un2kmriOU7cMxKCwLurIAVv2EBTd
reHhAy37WKVlumGTsxlGpTJ+uGT6T3fD//4AdaYcSariJ+2+ojZwVsBbKpbf
scf4mhNM5lyAXRXl6Kfqdx8wBavromeYzQBRx3tq05RyNXb19gHC7Fl788e5
kbk52FVdrKsm4fqU3GCA3eXGATVUO07M6WfQJxdXlQwpMGrFMjEE6okHLYr5
SZn1u54+0hwHHOOC46Hjh4mzmxhPYQnyc6nPlmqix48YGNUMtvFu79eBIasV
k7/lNVDWLUdkCB8V+38kfmh//pbsZPhtiuwdOoZyNCpqENHwzRRBZX+/r2kR
LlqEMJYQAcw59wWIcPxzn2kYwn1shCy4d9/el+V+wPH6iIGEyNAExh0AB9CU
FnT/fF5VnhUfl4LJ7Jd92ZWeqVcAgP9j4aRwq87UFEBoosq1HnQcsdhutH6a
0kuXqd609tbLg5GUxei5eQTGg8O4DX6kjR0Jah997uTJkywxQ1dYm7Fq6o+U
ZtFtHsefgL8YIOJyap7iV5ai6VudUvjJHmH5a2rGSeiQ8EwDVPOh5wUke/Cx
jfkb9FSMcFRHBq9RaFR2FEr6gyRl4y16hxh3hRFfRxw55OzyGbsyrG922Sd1
ooqNs8xuvpGE8xBsoAu9/BI4BguPFN9MyjOlEIYuGedukg8aiKdVs3LPxnm3
C0V7dj5rs1H/4N1bjUQsuI5pwlYY1KHZyLbAkt8x8Q3kZmyiE5bWchbICy6w
8DHSI5XE5pBCzy13WIHu4SGkSkg962TprPx++QDjTRO2431a4wInbt2IdDzU
HZoxbTBcfd0gJJNPB4zm6MLsCH7ID+BiaImZ0/rLKLmMDMiX55zdxUBKBd7P
rpet6kqdIEQCdf8JnJjGD/RmiYWjPIHEQaqyAixh81gYxG9YtzPQLmqNnaQv
8hau4FGSxDTUqPU5lxdkzXbDUWcpwD4mszpvjdmsTmPw6hxytTcaeYycc7Lu
Jq995g3iml3a+f2L9jKeuh19fgnG9hge3jyUORL3Zp/2DRiyTtgmodIQ5I1q
OM6pLWvQgklOVWjsVES9AB8M6TGQ8f6CJNHN20MFBuxH6bee3y7yLIhvWo6K
33mlPTXQkXIGdU7jHvYaemhxS3dE4MFTw183+iwbVC8HB59V/nSUYDP8/kij
g8tGf0YiqUJ3U7VJLZNc/DlMxgMvB6oThMTKh7krGkhGVrFegT8Fe0cpYn/t
OIIbQeEydTFFQcH7Hpb+FWI49bA5BsfyscTszBG8Xh0NrYsLbBCB2+j/NB+e
Aydm4qrkEb/qneX33ajWNRzsiMKcyV9R6lqbeUOd3BBF905QApyGwl40/qxm
ExndOxEUe2l4AxOI5efbuwgLIn0W0hfkKGNxElBatJYV3sahAq176QxWAd0D
4HQYls6fYTyXCAycwxL3Junuzh85razSr0zsaTZ0lmJFAstXzGMFN9YOKjO1
G6iukPtKL75y1LP8RAEOw13h5vBihuTrnJqW1n4+alAt6yf76X6hMmykRSgw
c+moXj8F87exzY2mZk+tBdVpImoqzRblOZtNpHvMWRdgnhAVdZ+r1Ax419WV
08cBYen6B64S/WXcuzHqtTHc8Sy/BPNWbmv6BLadZ9LE11UMoKXOUt6g2Ku0
/kULwpc3t6T5gv/QU0cVaikduqqkRW42UojQIRmcBckRmoFfu1bolw0zCJny
TThx+K1u6nqQybiCeQ7byzWBbJwYPwadkdHzqO9EnmaigizM64dXTEnyqlQw
dkSsoysdB4oRnwsxE6PAvW0j1EmUDi1cBX40ogDwU6QD6qQdIwVakJ2dFxUs
961t7KQp8e+VXbnB9E2ttsHf1ViG2gY444oIu73zV/NfKYDafAWj64gCdD+s
J/IIC0WNiyxLC5O04yuLduJncAvXjhXUyoYTHaUjfWj6E3T8THFRxSy51p4r
JpPFa6sSnFlImZoXpeoH9B+IPgysKJkQLmom0knvC110u4jgWLpeq/ZelHLj
2XTYuw/UOpe7U4qRmP+H/shYZaWu2p6dvXygbLMs35U8WvpsD9HDe9K2wOvw
eyYj+EWehICipASNXA8jLj3Dm37ByEFU4Mf49UPIitxz5T/NiqL5Jd5OYTPW
Mbbq9MOZBav4VEmcb7MFYrywuM5FluCE+spjB5WEh2eOL0RHoz+ZHbyoeCxK
14r8ZnXhlCVbl7rp/pKrKsN+KzHxiZJtQ1NYdcyKuJLoEZkGyw+pG2BMbbBk
8+ZbmzlAKEK7ACr0nGsqPgBen/FWD60tcqUV+IHK/tBK2MQMFY2r9J+gOMhS
24UsAZvBjpOy8II7ndmmMDGmAzsXxa+mZqxVRhFP5SOGMp41eeOLMIKhK5S9
jPT+ONki+s5lGhIiXQ2yxGF8NwDxptaWjHY2W+WNYepwVL3ge6zZR6r89bOw
uhHQS0uVSfgr5pgtJDMk7TFDFUpAAZqcoSNquWHIAi26fBdglOT/xotMRv2f
FnxVLGMVOMOROUQ1bM0XVzBgy6SRk5Qh/n4LTEQfFiycXMHAKjVlabjdMsnF
CB5YbCz2v7J+2MxCaBHWfd8fT+cRTt1PNunTCQhjZy9PhilI+F619T7vP7+/
rHDF2GBpfnNvTKb51Q6iGhB7t92jjN49x3vFBOGxAAm5TRa9he0mVddmcZxb
DQqqYkMdKNgoci+vyRZD5728l8arXXNvdKphNHhsbSRuryUe+CsMKUvAoM81
kTlCq4hMMp1EgEYXnRVbX9syWR0SsYIN2Z+XzkCk9r3wLIGcUPkF/oSXcj61
iADvlVRcL/kk40DcFWGpARIBxdH5yIBkirYNv0dH0qO/ty7HoXtBhiT0G6iw
eta9rs6HG5jo29rqL1c3Ta8uXEPGgxG+bLvxjcdjIYBVVg9a1VaHktthq00l
wvQJ0CyiRKvKN2yvA29Dwd5NSqYh6PhyP9IiQtNe23BS0aD9ZZ4NcoOA2AXG
jBipjwj3G6w0EEWExv/vnKRV5mSb2PqCTJrWgBftxgyUYM5fJD3fj7QLMPuS
sTxADM7g/pWoEpl7YuaFNpdATCajkfxHAKkyAgjgxYM1+ftbCZUOAAINfCLU
wH/yDoK3kGlIKBftgF5QZ/Toie2YISKiOZLqo6xqEQ8LI/Kd7uUGtk3tfdb2
HMSZImHbdUSYsfXTd6yscWD5dfnxxrEgyd2vIN5ouuEzEsdxCu0TX9MsGgS/
edPR5Gi9x52FmjEhrda4cJX6OJ1WdetzE6Ub6leVbLwK3+5XOgXRVlcDk1Yr
v8Ozq95Z0ToUfFJf+YyNreeMhlWXVOpOjoCLX9qpa+5hEZHoWHB3wYHWjy4t
HVrAg6vcFo/TJm70CdRIqPPXKHFOMAwci05O9K+ia0zzt4ygjkH+Sf9tilRj
ENfQDIctaaM5kU6KeMF/oHd1o14/PoeNMBIMKlN/FSDQ4SPQIdmtc5plLL2s
Lii5leg3fvfnOV1IGulxqJmnsMEFg0G3u2iJaYQbgwgPffM9vx8E0BRK7tOj
jWgiBU2l7s6zJP0ePYs9TLGx00cEL5D/EYZsWzGpOVMGvUygEZw8Q/hgfonj
bma6ego1wTfJm5+BcOS2YwgNI6Vhk9jU9TmxLREd1gdQVbug9j/jBzNwiF70
qsx2YyqBANgZlmlB6yxuHqtHth6vCZ7GtPog213R3s4n8GHYtF8jfdVCsJPI
J6foY9aaJ0S4Q/1x33Y4FpdaXAiKOUOURqHNtLvplGKnKVVrrNImMeJT21bF
JciKJ3nnHBwzIt954jhkDGC/cBG4r/Bg26S1C0If9rxq+rHavFq3SPzOgkwB
Dgwdn3+lp+1MHZNQHQRetvgFKZjbZiL9GUsNNvlhN3XJK+Am/TZ4FruPGOwr
KAgZ81lBl81EJfg6uMAtZKFE/cWDoUusTvlPSPIgUkudlHlZyhQtaOUwHPvD
RezONKHRpYsWR/iaQNiPzv6PDewuOgDkzV1C97lHnXaE19ceC71oajoVEjIZ
j1fEYcb3OlGfEvRH/EOAdb70rghJs4vDCzLiKUrqYDmBvXAjoCGPss5evl2j
se8TVHsjpVHuyRPY0o0SPLZlmWTEZ7iC8vygRu9xdiw9LNHcuQqJobvttj/x
Jjj6FObUGlG7/ESNf/Q3yszGXy7lXMFEoF97zUlLhJ/RM6es5kUqvAvB/35O
vX+QkIi9/iIWjY77auWuhejg0BOh/HsqcqnJBVYhByK1EQaElvxP2gyYHiij
DZrafohzQc/UrQ1A/QIuBrrRXKCuyuuz1ghfSwZZH4u+VhlZTTa1aowz0u4v
AdnfTCgAOm6PsKxRBxIYVVS++kGwCW2ZdpYq1Lrd2CuiQmZmE6JkuIBCl6oh
DFqBRrkG1XWyDzLDDgpdBEfVZIddtaUMQSPoo1WVt925WOcTDjtRPiFDilHf
unIf1kgbj/eOI8pnJPJG4V9abAgr3lyFZt0V1/F9xjTDhhn7w6V0m5myO1D/
FSNfZs+V+zfASGmvb67LK6rt+KoBUXQPqqvbgPah0yxRz0CJTacaOdJVYQID
PNu3iTfPewqAbXVMhz5mWYv7dXYdZIXqggMGuOxvVSOWyZipAThoSJJjXsnI
SOODZjUXa2VXlqgxpckbACdHqFIx6cS2KqVHrMAf/Ko1AEEd0NKOwJCrfpCl
oIOu2DUYPk5QFSygdDEajxV2Q09JIhc41GomSnX9JyN9hk7b1Rnbpyp508ta
SFHcW5qhKWlxhdY+CCNaNiaXz9LxID7s9GYA+u7NATxBCRwFQpdlPYdXYAL3
uTw7UQ7aMjTYeFpQjNWyVJn95CPRz0h6qMP4KMFo7U2Styg76QWyHNxlDn9l
vWPoo4y38gMmAdKgPT964UmBRNjFNaGKJV1bdmjG60sz+9JWCYS7IpDThn6s
+dleYQ8EKrTQFr1tX92PYWbtL7U9yVA7vOxBs5gRrp+Fpw9Ilq59m3Lvoqhn
8pl7SqQjZ6/wKozHZi0wjPUK4gZlVU/ieBijJGucxTyjFVu+1C/Cb/b1Yoqi
QEwjFTOUACcckniY9K+qBjKTP7YSi6WcnHbAdR8d13SuzY6X3FRjNiSTDiyG
yVwvYPP1sC+GD42Klb+efbkLbfufXFKf9OBKSC8whbMdyPDa9NQNUGK3ix1i
PmiqaMNAgxx5vi6CT3B9DwvzaRwuGetK7RCZYB6VXkW/NwNWhNY24RGRv0Ks
1mK9iFigeUuRcbj8k/wmhV9F+HRiYfb4RyO1YKyyIvg+xu/OWCflZNOzw0dF
x827guh/Jikkzs8T26v283vngv76a+rdkQipxtXE4QXdkuzwlDpU+IA4rKLn
5z51F6WLwSHH2nnMs8P8rPlzFJgtow1YoeEyd3Bnd4/uK6h9QsG08pNbq5aC
GZXafmlJwCQx54CzpuB4Mh068wVOebxJKpJQMbcOhD988NBl96C6br4+y1iP
l+2dvqRYn5bgFIFCrOippLl5HGo028Kdge6PYu85vTa/TvQiIcTEihUFssWf
aqK3p2aYvh3cVahMOvsJQGCwAlTq5yrGpJyy1q51aOjiJsj8AIxP01ThTiBW
TBFeJ/qsXqst+jDxIyKrJTg58nwPip0G5jNp1k1H0LEDofwhUAtLBps/8THf
FQO2a3CuNlm2wRWI9ThzK4vtZWvA9/QtvF6rEaw9E2JZqkJcystw4kDudSci
IrxEW6++6ywfOGirW0SW57jSgugKbxzvcdSeHva8fhfxfObt2SsBuyWzFFi+
2agbuet3Ws02MSVgsWkF0Rkq6AvBuoc4nTxByzUHogEZVHfOy4FBLUHu7Iu+
VKBeLkXmk6MAKjpqIYKgwdRS4MvLveCtZJTeDrcWGwc/+xQ5O8y1TRvHkkm2
i7ZbPgewaH/iJlLLS6Y9hHmtDpJYzrScdGG6uReOOCBgst5VSep+R8h58xqP
nw6zof+0x+rUKA5A/18yWa2032rO7L5eSoXCK3kTHU8zzCmDN33P5oop9KEI
hnisAEGqnWJUTWPnI337JQ15pU36a9NriZti1iJ2MCxoUsnMLrUcdGMvZLfo
oYp36X1nzgMjqUpzBuMdYO5LlJWG3peo6JWYGmJLJ8rDwCU41DNmJqyUbNLp
KA91gnuzINDhEqWJ5K9rUCdCfqTMK2VU4ebrmv/pPLMMNV8QtlCKnk+O/I3S
5k04Wjfmi6UyOBxF8VvSqgf0/R3mQx4O7JsRt606dLsIT/WOv9BewC3SL6ef
Gw5LXVxi7XcEhl5qnr7d1JwYN6FVmnmhamGRBxHjFURRtUmAvl1apZPyN1qn
vrfbN9fCmlKP7AQNyHuJ9tklfASkFtMSN/vSnN6Lf5z8E/KchFhkQoOfODnE
3noyWnh0FZgaoFLRPDuVw+sXZaeRmOAsRMU3pC04jEs1TwzpxjAbB1AA4P/j
+if0HojFZV9flr3xiutd0eK4ozRtq80nlcYwW3jlLk0sgPYxYDSd9TCsVUiv
xWwPPQvwErl0oYID9woaOv6KnMsWfcNqQ8d2kr6tYMDGwGGcjfvsC0vJZMPu
saVUb0mr0eY9GuuK93uZ+WU52sKvDi7mZQmFQzXhd7pV5FCrJyKBWH/TkGoj
YY7PjwEuRqz87KbNwqA1YduVd1zOm/lJk1Rr2h6fv6v3wc7hXRSyShFDBhRB
7xxODd9Ksr2S2R4oW+oxUlhzIk3ps2Z2YLVnOB6Tv+ySs61V2SRkthAzZ0hG
349+Bk7kTppdfR5EvJMV19cqQkfwwtilbq3B8Ri33ZgwX61o00JY9E6WdqMP
93xIFOL4xPevRbDrWIVcVV2jzjrbiCy2kCrSnEWpS12FCCgfqjDeGwuyhD97
iqbNDrZepXnFXLAT/D15T0c3aF/NoFpio9t19oNjijmzPguszNeVt9f/X0qL
2eQPa50Fh5JppFbxLDGCD1izagJH3K3K10XywSlhwTPoMsY9DgBEY3BVII97
SIPlgvGszzSslnRUXORxLv2HM11k4rhyy73b6uAt842abyoihBMeVZMgY4DO
U5hqMvh9yopAgNKfpSqCylkuOjlmu2CVci7VsmkmFKEC00n4SWTre4Pyfvld
ClK8l/YE6ANeQcbeRw7Zl6in2XUJMbzrYa2UqHN4BoUW07DBbq+CzTaJ6a+Z
bHZrXV6qNPbR9PezeYriMolkvi3WZvJojsCSSpdk8aR6vFQwklqsd+2DG6Cb
BEt5297OiPWs2S+3QvI1fAoAUhb7rQSh2FCJplxeRfvb4Dz23FCFpWTuPUuv
E1RGykRKaJoJ5UQ8j1cBONIX3XByOiealun+0sATUCa/WakpBCBBw2o7PX+J
wsustm2BP9y8FG///taQIV1nlgJ2XkQIjGn0zMOeyImJoGE3HicBtm5q1Qip
1y6Y5bhtL37Ero1HH8/4MPbJRJjYjSHt6NySf96EI4exO248ilQ4kq1JPey0
oo4va455/7ppbzEuvPDPuF6abAM2mXp0MSvIzKnd+jpXuqbagsGHEpC1nCvU
Kr/c2zlvWyYuUSLIbkEcFrJJtbcGSKTHpb8W3qg2F4NupiOmv3DhOjVGGRcp
ByhGMhqEfrzIrlSN8nh2mdnH+PSwnE2sMQ9tXmMKUmjd4hdp9sjrjOV063LH
xuvU2WqKOFw7S3UJdw+ggQKSStoAPqvuhDvOH4rodcAKWcWs4jJDZ/dF9uke
MlYGymB8+IFbs0D7p1IGHXr7AOzTZPlUHHha1nMdnxZmkQW8vH8VaVTjEYsz
dfic5nqqJtZdKAfIMDnu39tWy+FOnv/y5MOWXJvPCmmyGLe9gLRP6QcDTdWM
/mwBe2AzhLvPwHZ9jUck0qHzVxluvaibd3XMduTv36JooHai1+0FMalfb6GY
AzVbYiscxVB4afFrXhKYi08/Guw9Jj2vbZ12x/L4UiLkPVhTY9mzeMiiT49d
5qQvgTuFv1LYY9eO80DB4XeI//35s0z0SVlg3uOL2+1NW+byXrWvnrtMSoR/
gLo0suPLtxtW3xyEPXAieFnuUYmEQ7NU8Fp2bHVSRdpQ6oiuwmR1vJxeQeIF
S6yS+1+DTVmjDTEyz/TW/Jj3+ZIUwOiXI/ARSYd8odRn3cDSx4Inp6gMBIn6
YXIHtxEGotOhmF6PMICVCdcpISIeUIJKLWBBpKaDzKfdWo7sHQeDCVq1fyUv
5bTLwhhwwkTwBquGkrkfC1nXr53gX/60FDZ2imEeYbKsB39Q45fN2qHV97c2
mpPbEJJSUtR2I+aK5EX/efPJq6o/DOz8g4ns8Sk3BtrErL7NT1Z19U8d6kZ0
fzsWIwM8L508aaE41nzhRO+a88W+eB9MkzX3ZIzS33Jzs3ohZFZhE/WZ1KkP
JysX8hxZIq+LptZ5I1fChDoFHlHNF8azjYepKTjxGs6l0tEcvaYClFVsVtUV
xLGIkAVt4USqpJswp6uYfE4g3aiiJinPJQL54n95Rmz/7DbKQhUit2/oQbTh
++D+42v++ASx0qZSzajWQ/4ET8xfxMIPyJULpz35cKEjTfPlyzfxnDZlCXWl
kqQvkv2xI9ovT09UUgSJ99yswth8JkjT6M0w4v2WGjUloiaPdQ5lwSYqV9Me
1Zenr11a004itKmV00iC1ZHO9/CMyZtDH0rOJ7G4YkPyC/qIP3xbogdV4ja1
l46IEj0UQn3+4VZSNQZTFXLp6DkXmP19qMD3wQeDZBmqf+G+r7QTq8hkBXN8
EKYHaKeMpW0IETly7mcsQMZRp1sFz7RwcVlfIhWP3GmAWUb1ZN1tuWE3T9Yy
vApejk8piURCevhq2DJMPQ+nFbLXQfsqR84gPk7c3w1UhFIRm7SvSUz6VUZk
CdfFWV/s52A1M2inVZIDhgqfrHEsQJa6riKlUW1+g+1WKZo39T61Ey1UqsUm
ZmnYlc3S4454K4gQTO6AhaOfX273pvCu8wVKIkJ1Wx1smWdeM2uVH/0D0fXQ
MQqN+nmEeVX1Wg2gy9qWC17SkXudo2wJdSJtbrAqLGVrdimGEkxvSXWGt0CK
FN87rXHV/rCwtFkHNuH9e+wHuw90AeZSjoP3sfbirMqdjxqLaXfJsGbk8PFo
2lZqMAviKPpc8Wg8OSn9HTqbGzKnZ6lQEJBb0sZojY2Xk02s0BRDsI1ugBo0
02EhETJN3Vvt2A9MntAdlzoUcyEjyLR8ihmaLdy7UyehKnqauv8A1PpxMUTy
FoN/fQfQwgs5ZAidRkTkcvGiKt7vVmsKPPEynnyC9/dTba0lCb5rIS8aS7qU
2x2yIX+toMi2jKT87iPb7Gtnoto4WRSod2YTl7eL3yI/wpv+HnnN5XyoxNRZ
SQRqKBHCY8KiZ46zh/LypOfSsqPs5vuyOYRB6DRCz/sLnKe4Py5IwBBnVrqO
m5yxop4MMbNpQuP/qZgIAEsDE/DGSXY6Jc849iE7G32EM8luPcsVpRxWRqOB
2xpkQu8IxmxIQY1kdD0SfyACC1BhtecMvR11i1RyJSjuRXYw3gbwcoYesklv
lqeZ9rfnkldXvVfJ+OuhrA1A03QWfXTG0PZC0mCaiNXs6aU9kAThndQnM19C
qYN6b9sLCoRljmzL2v6wIF0d8LV3NJBs/l+PKmV2keNGnEcIma56GMd13G32
5K9v3IrfYl1x9ds8OtEhUen/NZ5yb+E5j93zQ+p9zK70FghCxUrTEEiTCD8R
VOf1mAd0N7vwmP4wtf3m3530eY6COrN0h16UXEvxE8Fa/vSmqPDx8a0Tke8I
s2KRFHS2XIDXHKltTxjDxNeHkvHuFx+aKU55VZKgzjAsljacZOdeo8UnOM+Z
KcoVef7Jlb8AOzRYy4yl6bea5k9yuwC8dbjIY5abblyBoBsHTWqK+t8AjiVR
frefAAUOLr/eMlb/6D4Jh8pd6usJj0rSCex3oqCNkePGrw/z/g+jY9SfFLFu
JPvkrDQBt3q4wep4NbZZ86QdDeH8KW51QhjLpJfIJeD0q+Y3YkolPJtIIjxs
iVAw0sjeP43pEFIYb+tcbjrqzmf/8gx8WeE9mVMGYd0z70p5bpG98UwxxTkS
GEew6VMAIUJpyFEOPudmrQGENslVcoS/+/hv7ov8T/6UCyUqhOXaxZu6DXJc
5M8nSo1dWi1tD6FMdcvOoCrjoh6B5HamcwMOLi3UloL0nO7iiM9/CALnMWws
CeeD18FKjR5dkM8H8lkynndgrAUxOvmw9SwyyAmcaJj0x7tRfSp17Rw7knKg
ef3co1ORgLGNIg1uTZRuHYAamdnxA+U4i/xkFD8E44I9wcwAi3J5O0RAVfi9
LwQ/8u9ExpbdW0DMnCaF6KqhNtWXPLP+/PHYrvhe96MieF5OLWNmGi8ITmaj
NmMAnYOdnZukDzlS7KvU4TCPSq22Zim1gLjFtYwMFqwmmXiVue7/1PeEXML+
5sg2PNDyyrQ54LEi6ZH6Yg/fzRE15CbphZw12mocoHMBVYT937J9TxSEKxm8
Vb0/pey7iz/2O4YmDxnMZ0NcRZzzswh/2gtWpQ2meajjM9/bH7s/xH1/j2Ib
G64Vuoc64qn9PJfPG/7ksKF5pwvCoXlB/2AxfkdU/3jnP937x9Zm0enLLl56
XvhK/SXhGHD9OEUjcFOPlomOm650dba0+XSOt9VGfhKgld09B9BQXkCTjsg9
rDlEqmKWxrPuukOqy80uWfXuhdF/9QqmxL+B/zBvQLxbKd4Q7A2eYev0xA38
EVFh1em0vP704rkob1iyHq3kWmcQDjrxIxHbaTQIF8FzxobdFpbxS6cFacGn
7ithrslw8sObCdPKYDqwOAWyXUYy0GvwgRtytqJThXa5qKpO54VSrrmh9EE8
OHWblglcD9OBLQrmd9+z4xfFXAYUSo9undlXMhIUrIUP9axMFN+IJAwbEPdD
ZEuQn8MyOvn/nlost0abIg7K6z173Hb6Yt4dB2hoJFXVc/wZ/q6BNUsh2UnH
FVXeDhJJ80QIsfxJ6sa7dQkiytzETKCsHD4q/uVFkJpE7d32t/pl5by5rj8D
wcI9LzLw172vuP3a3hm6p6lqtfLhWyj/1WyHLwd6yJ2u5jumJyr8vjBl0WzR
5arCvGWwp67m8HJKVYQn8LoSSQslT2JGtzjVhrEMPZkDSKZy8xvnUc2J+z4L
MYsqZ49LNIS4R2la9KZo7UTvmK+Z1lLactqGod5l5aBP5ld9KjgzhPlr5yFO
fWYEhbA7su2AA6TcGLea027Un90kbf5/qHb+SLriWGYQlg3KtndP5KUDaPZE
rUgHNvhyYi7cQmS1Z82T1x+R21biwuAnaIb1aNjMvMbYxMxbQehwxtlThk47
szIXKfQsgOKs+hdYy1BaZAqrfhiJmptNCSgIlEhz2oFyhkSlkseKrIGj7nFU
YoNpeFJ8Tozd+H+qUr7ZEsvfgLAcrQh0F2BObAc4Ks7LxABCk7GaGi/9cpBc
axhyfm9HpRbSRwrJ0E+gBI2Ge/PlSt6hebqYLHNwX/JaT3HSqKkpBPPiqNG7
L5wVqCHgMSqv38/+kYH3xKBTvbIxyR1U3JIQUPsu3IFgnesSUxbzfuvpfKpn
XP7QjK/rLQ+Kg7h+DUzw2C22PQu2kcWRUvUm8dKLSQFqWBZw01zgRQEeW+IO
VEXIwIvybituqG4c4GNFgB2AkqUJBwtb1BCP7MhG/RwHK0O75epPl8eNAloy
adKLy61W0GPO4+G3DyqKys4F8LjDTi7LoIDWbNjCk2bbBYvs87TayMjhSh8J
nVZdhZIoD8iOFQ8TGIKOIb2Uh9jtrn6IUSmdKXrX5giRVmcAvnTjpGEScW8J
xO1djie0r9q1dIhzRzI3+jY5RyKb26uPb1eev55quZMRQYhlA8FxCi9/rMxD
Ddsb+ye4KdbXG6BjnM6SNrOzYEg+sIuC8l4nzed3iKcWF/dqGbS7IwPRnSUi
a37aN7Qqd6bMQD4PMup5S93TlC8nMM23Z+97HVS58ShpQlH8/J7HHfYqk2PN
PV4O1WbpvlBCJC/gH2B6u/IDX0fWEEqNTjyQwnpQY9z1KnIijDc/65Mr3Wg9
QnX1X7YhQi1JNTFkzEUvnBvZHQv6iifqPReXi82swA49pudtGg8wAaBHEuxc
ywkmfytfsLUwEg823MWtgJRaRXZQ/8JbRR6lq4O/pd4yUVyGWzonw1Cmy6+N
z18CqrRe02TenT0OTWKOE1XbYwdFnfYUEL+pHHa0SZ+k/eMgiUDe9gs1YBeK
ryx+V4uGdZfatBgDqS0WJpcEc6brvX2oF1Kc9KLnar9TT+ldrAkOCkbp6M1t
KRV9/av+iOPp3wstR68F1ozu5xTmZY1dSddd4xiBcaEU6E7bhug9oNCw4xCw
9X/1eOKZb7nATmWFo20z4pL+LFAnyVQgavwaQoHiX+7U7ByHwSWuSWKSRaAF
NrUXNjUZOw7qFKu7OTuBF+GxziOzjm3+1v2OUlNU9iLoMxoBAnUrLjB0GqHu
k2noorqr90XGnaaV8lGTH4PCaaqr/ZQFFvi1wMdGu478e6VLAVbXYzPfI61c
tjuRjAWuI3ddqRKuXL5T/+SsGMVdFtpf6YZ/VJEqd7lI8tHICocOk3hYFH3V
o1jMJYhxYd1y6vMQF1UmiPihlY6WUYnf81IG9kjBGTw3NS6jhAgaIy9cNneq
zhtE6y1GvXEx/eq6vbrqN7JUCVzoy21QhRfC/zvPH6VfueMXgXGXFdItFXy+
+D02YZdqQKEtK5R8kKJhnrpnmpRu7C4Ntw0kj7tRTg8Ly7N0ISP7vP2UMVJ0
utSSyCSd8xnkaGgt/AVZtTao1bVN+EZRQSYo1A7GJ+IiqmIf+7M1ZwBPWW/j
1iGnfR2LXS286XdH75dKiNd2Sv8O/4LQfKWT4k8WBIcnNTHP52KRU9ng3DBP
jEMsttb29uojeDnO8RHBLS+morzq2eKIk2g7/fiDyrtjZ3GXld/rgrRBb0p2
Wle3yJv6klV2jv1LDE9rnoctoN9xwb5s4y089eaXzExlEUkgqIYQWRkKjp8z
3CRxRalCqeYprEjlqyqs1nEOunfrarkAi9vUlpiaTZ6LQ9Faufi9PKa6JtNk
7CTya1oMXUBNIWWwa31UKZc42g7m8xFt+ishou3TWHsaqFYsNK+U21LkSnOh
inEVLEC/4/G/u+7ULrGDhCLa3/JhB/q/BfG4IsNkqFHscUN7ST4Bt/qJpZnq
ISl6I11YsW/aBFBgsCtCBZOyS4zguDrhp3lj33xKZBvSIx272d/rs2OhQpO6
BBUgklOIlvFfSkVeTjVi3s5yDCQa3ye7bMjc1cq/YWiEFXJhGB0BAx05TEOh
qKSiTr0Kr15RZiPoksYe/W37Uw8HJvetLLUuGW2zrUqJ5sq0udKyUyrZIvkS
33ESqgqBNZnVCISix2iEMyYrh+ibQNBu82FivdOCtZDU0pI7wlKwUOZzqsD8
kOT8xQc8Q/acIoEguWRd5Ggln49GHsp4oBx5lTQGdxnsUEGJswhgbnlqQTxY
aC/cJNNCiky7nGWzO3CGTDn3JSRDpUFQfPbkV0SzkRmk4Vcd+evystgyQSQ5
cVfn/RE0Q/OdWytcosq4DZJ4MyNWNP7izgh5/SrtPEeBE5rKDCiOKF9C/Foa
UgzJnB/OXKo3MqeGHOpdLnNAzbGgFYBUGNApY/mctBPqeCewNCwBDNW6ZUPx
JXP5llLpnVzDOqDsXJoOKcRE+anvqePcGfOHRJN/2Kb2gd/HV5p1XTDFjxan
ThVVmYEpo+Of9I4P0V4WJd9iub9OZWS7RRcMLNXQ+W9AiNumdqzlPUbJ2Doj
tdid8elInvN016dGrVu845t0Lko34myM8sZv5vjxY/ch7R5Urh3GTKXpDEup
PuoHnLgVFn4B2jdCkY+t8GVhhYPIvJKVCJcPORsWMBg6eW56/cm0L+jpAOZF
H49Cxsh68TNTzSUTvhOUjNbjFzgkcoHgApuZ0FYYEO62YuM2MnSrt9uzQahO
GXHNtz+KtYpWgyaxfXt/gblgfaRLcPIvjALZhppzdmXUVgOEnK3JSyIX3u7/
nJTXPe/dy7flFsye1/6cB5fasn5HRZ0p1T2Av5+TzbskgdUEYXasl/84HukA
haV0YvWkPG1KInj4qPlI6I2j18XoPsczKVf9ebdaDpm5zkB2hWejgTJk3lGK
Wke2d8NBUh/+HCPXu/dm2ZWdMhlukf2dTvhRUTE1uJDIGbk4PjjHgX1emImc
zklIyYAa0NBN1k4ZZiLMzI5aEvpt1EXfuE9YRvKA7F9aHg1epBh8BXnGNccr
vUaIq+1L5e3MlRtnTbTYj/pNXNYqCRHvtTnry9ONqxLp26RZ1BJi30avcMNX
+9QhxKC3aXQy2+iGbRuA743QmjTowgdHD/nNkYIUaW7oFTysX8g1+J7+Ko96
Xfb1MYtn+CF4djHyTvuOE7Dwu5sJ6jRbS4aVKq6gsAb4gf/Vx2UdL3gUEzna
Ihi6UMDclOpnq/9TN2OsPwnz8YArUIbhWSJ1vXZKid8TARqEuzn5OlT0RGZj
6OOqbXk+M16/TefEIVwty2gKJLvIxMWQTfQNPoioaA6j8B50EMPi/SmaxUET
eL2W9xpWcYI5GAVQLMz1xop9ZL3H5Lb7sZTwhiTNZWj6kIScLoEJBx51UevQ
RnZRaIjhPH0Ra4ZoGGyOynj4ID4n3lRLs9XtK3uff5bw/M3+A9Jo1R4YiPYI
F3Y0qn2HRgRoWyEB1Sy8JnG2IXV1CzwWcz2HMs1fAGwrpskLTdFwuR0XLTiu
cYzkW0Lmj5knnPaCWX61b6ieVq5kSySy8XGKGKqT5Tz9VfjOxFfLOBrTY+jM
Jw3HD26eUqNWKoj0Kly7YlklqmmJrbTgeauIbRBS9+Py1MkgibSfBRyy7Erj
LgDigOs98/JOeMY/Q75NJUZH7CZiPrBBM8sctjxgoQl1RzJWbAvz5Ckbob3+
5kgtzAgjF+Q//SxWDX49l6Zxc+UrfW8ns/axZH3yxKTTcdsMoNqZH9tsBGrg
XdWNVbNXq/7MHQFdGUjHMS7qNEjxQ2fIsO3DMs+WqSrvAeBGOOaY92ByJfRq
odp/bYFxJrpvNS7gdn/2y/44NPwqrgd4iTq5QCn0r2COJk49fvo4haE27GKs
3NYd3W+T3Bn8AAQx4/Sq5cQ/OnpTONfNXZTQ3ba2lvI1U4M+oPRzxGQBnS97
Qy05xMpQd3ksqU3mdoFqqaVVPDtio3oqb1gCtzjyI5CCjHfYtHHUFZ94ox2q
xcLmoSeU6pQmo4a3sKb15qa2iuwo1EHhXcE6EHcHRC/nf8v4QxeEV6fSVyEk
HJia8Ujhg4AMpAyMyDxF42JVc4tfIlj5UFzq6ugCgmsMx2ZTosO4OcALdMYH
F/vyu4gT3tADOtruWWCpcfIqUPNwYpzBV0T/9n2p/rvVx/t7f39TG0B24zYP
plvWWc3nDDh57dkJZggV1HTHyee7oxPZN4pXWwPMNrGylAodjBjbSDOA3ivZ
HBCY4Ad/tXiwj9x+t3KWLVyK8YvsAq4JeyFe3ncxjXArpLdK1KokTWXV4xiH
30cvKDQ02JTDBOSpi8Eo0GKzuguQBxILzio03uGXTdFfcgY8C+W30Baz61M7
Jbf9y3hlOZVmt7r93Z16oEusxr3kAMTYGd1+2W608W3LGCI04REafqo+Ngd6
p0CjTW0PrL+GDoldF5/TqQfdGJ3phKyIrnWpTfjaxKq9a1vxdqqQxI9bZ/P5
rJuUxYOEDuG4ALhuiJvMjnYx0dFVfJTo+XoPyYwncAEaxbpWLQDEs6EUsB9/
2W6rar1Z4Z88kGQ1wi/5qLT1gaBO8UZQa8VG5O2v7gkDGauZ1IjckF9yd07H
LAIxcyqFhhdgBFcqd06s88wD0tVc6+1hobSdgm6jKehuc9N0UqDOPvPhdxgh
j2QSj9lfsFO/M5BSytq89PrPrq0ClqwwYjZKYtSG5XvlfMgWN27jBuWleOZ4
7Tz2bS/Chyp0mvWl7ycUkZSUxFZQ0qFwztokosWW6fRBdgL2IXJGDke907nk
0pyD8oueKdM6vyfm/ZcdjTrM1s/rA6yqioqF5XHIHEcaLKfgqHo6uF9Nxr5x
bXgDWE59zyXjRbQy3P+H9jpoCGQbVKkvMwjmdtIUnrN36mb3zvkOd5wf89Sa
l2AAMM4OMxk2PK9FlFvP8WIeqJ13SpoQGOAabxouxhOboTZF665ygyPRkAQA
Cph9NQAbPZJrERppx9W7GUrdEhnmE6nrVkGF8pL9kVeZzYL1DVGj/EFrIM/u
SMHKAAwKD6tQZae6/l6q9ddFEqinigxHiGR6KC3BoVDHVy8eILYon8akUXDw
JHTYTSPV46DUxZVfTRdwD5KqXD1dsvF6RnlKz2QPuN4ExZ/DAKNvdqomgH4b
d46HPjKU6q49H/bPrR3dXb/cHcnd5m4xgyyFghsREolTYecAnYggKXESJ+6D
0GjummFivPoHkdbqXU7pQ3JXmPuavlZWLV4cM1ZU1PVIc8Z8ix4YOdcNulgz
7cPfDWvPa/UfgT8MIWMSvWzt5FljVB0jo+avg858Z4QgQ4ler5N9r+DeBhcd
eCDDBsudwb3EtErgq5BNqz5mg6Cyx+/pQxWNuHWmrHMQKpWTGzZltzy8Nd/e
TOMX1A13lhDXwALlzXF95Yyf308Ql2qvsRehs7jDijdyAABW+XnbN24FWrpM
YxVb/L8DZPv046tamkHMevcZxfhMTx5u+E3A3uKdUOMoYh7YmkEVAwskTR+W
fGtuSu0pFXe9SqlB6x3QOSahPvhEnmWwNLDyoN6eKOmU4fxqPAw6F5YqlmKL
MlZ/zBNelQxfpBaeM9/ALEFILwRJ/wy0K6R1re6AkxY52OP6e9JOtfe8FIQW
xWmvEpd9S2ggxmffBj035YtlEiNH+7QVBSkqBnS/N/x3TrfvoeE2QKtgbxFx
FfyytOtSoaUKA8biqCpBfc7PNh43N/riJV8whFE3T4g3yspv5nw/h6WcgRzV
TU5n0sfHhjmPBkpfOLEbFY7cRpR9U0xSr1TQQVXBDP9fM0OVoUgxFHpOzXqC
Te+cNpVsv6Ia4Ljh1k2DN/W+M/yFm5+HL3SyU6B7dq3TRO4N6NfTpD3NTYQb
DnPlrE/TdA/6NAcChrDcn9HwQL8n9vbai0mw4rUYfTQE5E+NuDWLSz3N465F
ZKk8NjJ4GCO9nSOeT00itZrKloXmRb5V4rGeLG0mfo3VXTxGczk96+HWxiN+
nqPkihLGZOJhbsnAuqX2JH1eqQB9I6PFcv5opOJ++e6vN/OA3C3caLw0bQvj
Gy2syKAGC5CZOiOlH6QzY5VJzmGGts3CaKuXS83Rp2egkw2RWsuPFmDN3Mya
gXsuHp8hUbNOrgdFPGW0P7SPgTu4LUVwiFNtk5w69D8Gkl/+XOmyC7QXo6JL
Md6RPpCsfLJ0h8iokFxfFpP8nWM+t5BPLu0pblehQELTvcdGq8bfOWHUSLkO
XViPP/p1WnWCBrTVfGJHowczFWAxn2rKwqjOy4WmRMK2/c0xDMhKNWKjdYCD
bGPKBztqzqdnu1bFpagsr8AOzNaMJ7O1YHf3xLhd5vvyM+433SbrT0vQxHsH
rZhiZOaPvtQ3mNk+LeLxJFHbeug2TekYwZLPo3Q5DsyZ2aQ6mEgQlOLyRJyv
76BqvFh7MlVWWONtlMaScmgBdXAJH94j3qpGIilmSrnSNNiN607kZGteiIeM
gFx6a4bNii51+cQwJ3i8JFAeldliT3JuPgGp82FW3iNptlmKJTjE/pGZwIFr
IVm4ixiFqj/xwe21/uHZ1QDf8c4auerpA7ujVHpAo6Ls6gp+WgQXCXAWGX6r
oEIy6E3DGSfzuI9jzovGzdrSc8XR6EGbnQc8haAIypSgAyJRIch7M6Y2P6Pe
rG5ZsbFG1zD/iy1TfS//1RLrvVzf+5GycCE6s25HRbe+yAdZ3FxBMb+3KprZ
T6neMdPFik4eJo7UUy+vAMrYgQTmu+vrwqK1v3RRBB85cEMh6HYnYIC27L71
H1eiadHvoHI5X5mjzCAriE7RMT1oASMS59lJuEiHbebFW7hr+UI+Kyg2vHoM
0ZhDOlMkMzQl5Pr5+YtB2VYKFEzGpxUXTCvp7MrjBti5PyCuJWWxDd2D7qkM
aN5s2iACFhUNxKa0M7QFYR+D+GqDVuC/ZnonEjZUrQnxOpMLJA4Ysf9drvW9
H210jFqL84/rEtdEZXM2XU3Ng2FYgrhCUlQRpQuy4UaZ63Zv120nrm784ZUs
9vcOxGiroQb6SxFQvz9//BkDVQUBUlbjAxnrVC4VnP2ZpGTrNYeIkBbB82Ha
B0L8BI7EKfyXlU3rHNnkVM2QcONzCl1mXYFOCaVaL/EoJ8wYDcUj7Y0bC9tR
YIkQrsEYT8FWJVC51/sB3xXWpsM+d3/bgCmNbgDgE9/UoGnjzaadPGoUCzDM
aQsrdqX+CZDGkcTz4Ew5eOZsiVfpTf/kHJLx29d/HgnE8TOOAONVeVPxVx7N
ZiJrpl9hH67+41QctEksEvNRE8kCjSAsgH1G7A8GSrL9yV/kYtPZLYkQaWiz
GsemMBSgg7iyfGsGQ3wAd0WomI7if6orTZCZGtS5+n5/6eBfKkTJtRsWJgzS
5s/xRog1ictlBvP51S4wxp8GV9g4cO2w32PGx+ce4Zc+PrhrE3NpkzoPy185
r/YGZpDxx5y57u0MDzq1bn/UWls2ic74r/SyhaMIYC0cjoGoHWV/4Fxly23K
lrrhzy2Bkk/ft913YbwCmM6CVim2v9iubI9jOZ7N+Hnq1wtJec+A8/pbOBxz
7IbGPMDoLTsPldPcP2fB38WlZ25/y4rsVb9GCz3yL7sF/eTOZOn8yXVRgiBq
1RozT2FxwNNkrChLOn5SlADiuX5sHOrv1tKtc0z4nqbOToCImik/UWy54gjG
S1QkbqGZcLj7em4b19gxbV67zSOKf9ZIzu8AmnfvmVKNFN5FIN7kAO7MUT4w
1I/7Kp1OAu9C5p0GWAauHc3f93MpWS3kxDEJLGxOlMH1VAoptsuuCq0qTH2/
0CiES1PUqswiMXihfvB9uIDM4IqYHm6d5u9pQzrE89jWFPaKTjc7gNWSpp4J
bRA0UhkDikisOgrFZYchaxNf+X/N7TzA1/npSiIjXMeT01O5BS/vSWb4jPVa
w2WybMvOCsDFIvSfphFHkga28dYP6ccRWdLqoxe6ivGLY9EGp4ywahZEZ2zW
k/T7sklqTzNaJecu4fcaIitTu780eBJbviJvo310iOBv6IZ4z+idKK6Q+USI
ySwlhKLMPf9btkri369Bm6/2NPTfwEhRzwRNJOV1bl7WINJtUaj9feeGE5vR
xtddYiiFpnmr2L7+JfGRe9LGdbXgZuOVdp+gkFpNj9q8eXRKJ6rBUICvv+83
NesASNjuOo9YeH+6r8c4zx/XE/7pltugQ7A2QTD8x3zr5PgMNkQa7erKkKbY
ZHbJ6bNnJGhh6kTihm/8wj6Z1U4riVm3oQ5CC31R2AoRYNsIbnscwlPoWYQG
rxdY2gLsNnLWlvH63jONj36EC81zEFX/yVTEji6m1fblRPou4jP73i9uix1R
EvBfszuNhBY8Mj9IqLHzMjZgVed2WPO+YPQ652b1YSxDziPPMvo5hwIO/u1/
35wZIfIXqYu3Ag8JzEzyRw+sOGitLOWJoBv0MIIvRAjInUFBF30mqbNJHvGt
+sM+ncZewk/YBxtI7bpIhnW2GQgm1lEmwDuwswNr7FJcGNwfHnyUq+YCPs8X
nPkqCo8M/dQXrJV3Qm8v60oWwTU5LxykHCFyOHDXyCyyuV4Rq7OBpiQa3ezL
CSWFH4c7TeCAZCDXToTe0DqkRjqxIhe8bByKyptxnOs3SDi5V21xncWEz+Sp
+eXQK8UmUVZjJURd0wPaNYHDfyNL+EhlXu6fhkjDSVY6PGKiEBks6A4ryIHk
9NOG9CHC5rV7LvhIsKEUeokwGaiTsCcC/8coaXRhb05r7Oh7YbxYuw1QKcpT
z5PES4MTLr/dPnxyTjbEshA6Gx4fQEalvoMjdBFeCbei6fW1yX1d+sTpvZLE
2VUiph0qPO8IO9hyUv8NhhMScQVmfCiykUZRL15P9r0Ph+L4ajaaJAYIhsu7
dwLCIVCaWNrDs3uub+NbJ8zCY8gujL3PxF8OxEJdIuPYwWs4ouR5CzOoJTnx
CNROBbHNGeY/BX4ablOFWGfcqu3E7oBfe/IafcP0ixAgVgzDTfxtzXTH7D+i
86iMvmVP/Awvkg705zSziK8NqsEuVxJfPmCoqOdcGat3y14XYWvNMNkZSv3J
vUs2oHv/iPPirZojAVH42F9fK0lRZofky37pcLLTWsvo5vNjZZapVntlDk1J
hbgLIH/9h/Og4iPc6/SCuxYaIVE4d4FrzUx5vnirYALVm6VqyoGkUrTw297A
YbfSOMf2IIFL17AshZqImrekbXtjEBh75yzl5E4u3jel4h8LJYiFsAw+dopf
wL4iBTWW0B0QUoHxUsQ/LPGlhkEcPG8ly0RdYyNv63qE5AEO2Mg6JzPGotr9
qgPgWny9YDS3naxO5n0aOAMaqE8CjjpuVdxrCimxvWPMMujAWQGQUyHRSveG
f1zS1epejv/SqYTcwltenA+Cn762hfY/1B1AelhYKK0CB+a3qzElj6OCIrTj
yJ00x042j7kn3+qPFxn9OQ5nGDr28L+5Et2OCWEc6dIeWEKWhu25/k+ZXCL5
nxx7pMzyN1uzIcRQPfmJsC9nclbOG4VHRLA7xV6UEDm9p9m79uR/YViR6/RI
47FMv1KmZqq46M05G2tviaNFR5SBLsumZUkF9Gy73IzfrGtoKq65Md64lvlb
mqYiryWIyFBydCzuwoZE7YPLz7tZ1+OM6vh26LZwXf65Q1rX78HSTR344Vsr
TKzjQhNpk2SjCB8yvSxTB6fjX5vlMfFE2yupCtcWrsfFQUcAhuD6kNNYgVCm
5rGZ5dzTliAF4F0bYoBaxLxj/kUBtPVkWVL2CRpaWKti7Z5RN+evHdu8A2M1
BPVc/lq6AICOo96uT9wzlmG/RkJVO9k0kwizJmGaxhPudBfySCAbEAZrZcKz
7WVrB4kv3cwR/+pEnfqojWvOYz2O2q7tuZGpagRJx4TgsQiHfpu6KxbWn6Mw
0rosNnfVZkVrTEMwPMLwDRzpap+K5Y3su+xfFXH+iySBFe6gqXlpOSu6rwHl
uBtrlimH7wLPBMHcfPFx6FZgbBHkPvmEGj4gATOzzXrHnkp1KVaLXGzLj/+3
qirABby0wj52rfgjBxZrnop4RLSCiDQpBZvwRCiKsQhxiHUPEbmiDBcJn7B+
8LWmOQKGlFSnHW2GLHbWWbDFM3EqXx31kken//mN/a3J8dMfm5ST0yKDrC2h
I18tne9YGcBsiVmQsRv7wH5wLlZX4UCEftLOPc7HEhFAqOvvIN+9QV9bhSTV
naRyZxUXE71yL+xUGHrGfzHqIDzUmEIBHW0uzW/sBH3juEHYiiBcTpGxPj/C
vpX3aZYPcQsIDXEujsns8iKcCwRsRGIZCVKA+IhsiBg7cj+ZZGDELUbMZKNe
CReB/T+MDWXYX78wfsq8PrFpv4aswPho8qzHcaDJ4TjggsNYyaSHjAk3jZ+L
N+jcmwmFJ9aszlDeK/1JEBjhXJTiRZR4Q8TF5Jg61rEv7jfSE7Zm8GsIdFjA
LBIkeP3BRzFti1NGFvgekCFDK5wwLYboLlo/GyRTea6ldvdG6aRFlVlhMrG2
R0AwzObw7ud7ca63AVcyMYGdl+I8FNIxquqXHj5nJazH8DNHbXHJiZrKXCYK
rQEfV94f1yyy/xLyM9oFsqe85vJfWrUmK48ZBIQJGji8gfOXQFQAIZ85lmh4
93OVwIR4KRs2/Hei2nTqC5BL+6QNZWCrhlylWAChdb6cQT+Snjos/g53LfTF
LROev3P+FzM1i6jUqqpG9AzwmCbxqpo7Yc4aBbN6yP6M9FD+821mv5ycM9bX
L+/nD4u2Xo7UHMQRiUSgUrd4gmUh8kl9SJm5IGOi94jPB0KNSrlfc4BP1nUP
DzHOzME58sPqM4KbHScaUOqWjwyAPYiupGrOS8QJ3rq+XIs0ebtYOwChJBpP
PGrqaMe8VkXF1T/5vLGvBO4ypMbYo9aKDgbfAArOVOATRDdLKm5T5IMoaMKm
uYW1XnBLveXHi461cC7nGPzvs7Lh1iVWjmgSevSxx/xnQZlyMMgkguMGUMup
c2q3yn5KuWnAkZakiIY+f91+04fAuToQUVlCnQX9u2pMOb5RNjoMQ96yHhVN
33z9FztLUxB14BnnWuG24kXTBNJ+N9cHIsZl9NMABVpTUsjWvHkaulnSQo9t
58Qp6Eqmf8jYRbY4KoKE5SML5nCQMdD0NPzkCkcX6TQY00ETCzjKXU30hx2E
QobORN8Hu5IUQrL6yLkXZqTPDKaBjStz2GRNJ5qfBicuDzylz1oj5PfI0+sl
AOxS8eDN8oUa0HmIKYaH2HodN5SSuEOX0kzfzcrebV+okNJQSHQYYlye5KVk
l+SMOeLV+nd8wgd3jKgw7t3MjHDlYV4iekvEFRMkL/tArRsNcWcIO9XrFZCt
IALaVlx5LnbEDCLIuyGnazrvIGxZAtwyBSEHEHu/JYEjuQAtIO5cT+Ru9H1k
yru49xtsJq1FO5MYx6ltbgEKu2EO6NSpafgeTvWGJOAbXPXl95JQF0wboTpo
XhyzkqYyZZ/qRQVr69EO9kgsPjGIP9kNbl29mXRnUF8+dWE6IxV0MH7MW9dU
9FZ9k8E0yqOfZdickVQjWhbcu5+fQMWQIXfsgAZ5QvD1suGW/J8Od8FrN/rr
Psq8DmGYWrKllAXuZdEGkXGfabIK6IuVoF4XRt9QiEoiMMEWw6TgES0f9E79
SGte/KBRiV7QCzEJ1oOd4RkDKvfm4jWF3DPQEHcmN9PekBO2vAhhFOdxntZc
ZVuKYahI/N4JPnpvCAmLd2EdgrmxSDIwmaVF4m32y4DrL4wiJrqalS09mxd5
WzNYVAPGasbTM8hMYXkEARLQ5QAvFRwtlqrwMDmg09pHf3PmsknYySgrIUs1
9Nv10sH5wLmxzODPiM1S+ioMhhIWziqCygr5z6U5cChFgsuPsOsfc/gcfRfN
zZvxzDxc1yymtCTgc4wzI0mXX+qI9UA3kocI0xmxjEm8+jKII7Z9fYPAE0JH
YtvaJgm4K2HkwtYmYy1C4bhleYr2fvEXQRgO5qKmSoaKWuLbuV6UlIV/lnrr
5eOhcXouLuT+lW22P/cMqqbegUwGeNYDta6/aoAXkl6OIMk53gWZi5qXZ9KS
aiXuv4Klhx/ST7U9bvsz3KpUu76AOIVx15StDgJv4W6wXEUnrNnsB1J9crVV
tvsSth0By2b9epJiSQ+JQSZG9p6j8V2j6NseDQDjut55lCwXL5l2TpL0OU6C
f6qbbZ2UzeBZhAKSm7rErwMMd6rvRiPmhiI/p5Y6uX+zX8JXF82RnE95nBPT
fCTFIXC6d5kyxsjb2yyGCWGIe97cqhHGtG7JXjKKdS83F1QwfdrLf25V/fJB
UFU6ze3yNiMj/QAvpT3TW5aB5ZodXB8fEJaCkIXs045hZ0zhJqtlEkxaJ5Gu
iW0ccqcd2ftImn+MsjTtVCqIohJeLTfYBVf8b9l/g0ElPi++H3N/k7Rms6CH
1Ou8WIIzA5birpakWTAa4lZ/i4GPUUfs/AXCDU/wUtvuWg+HFSEcraOsCYAV
d/jod7OeB34ZQH4XIyhKe+DYXlHUNU8IAv93wwcfEP1gYlsG2a9ReHIzXR8q
c4wqgsYDHMIrhnVJRHAo14iVFHJ7W8y+AGUHfFKnDyUdCaa8F1GM7VQB0PI9
EVVsTKhsMqWdDmk8+vDWFMpX8FFxtmBXBOCcRpRCb/Jju1vzaySALa/YuX20
AXSM4VTOlH8nq6JeCPbt6oFZZ18tkleSINCoWOeaFqvYSCqNaMQUkXgljeev
rRsz5mepqYlepDAhVKvfmmOlrgvQSqMgpJzejtNGuwYnRWI2ZXofBXzdapIi
DKpkWbCjTjhOO1/x1x8sBS5mAFQfOpwL0Sy3vEWDe8xE7AqDYR/PwulCwwkX
uZclp8gisC9mFZi7ZtVTw2fYVCzIYXR82YvYsT4VBZ9LfarMRkSB3jcoVIEo
nIGIgQSHEpPpYnP3xeS7IZhZWoO6XGuvqXeErhbY2ERS5tXKBV0xt6PNaNjA
kGASxUdTcPzpI1jsTE/IG1BfYH3NE4hLm2H1cK2EWhkU1l6jIiuLyvKzodum
IMGOkxWxl9KJL7BTQG2fA69wAp4sllviX5F5uthdpcXM6oCjG7OzGDe7whig
eEodqJPggk8y1iUjLP2hxjdbcECHMf+my1E4++gCY5IBi/B15DHQKR1IrGjP
uBVybE7bL2x3Z9YT032ygz3UN2P7Ky6zRLRsN909XjMFAXi9cP4PqTQyneF8
t0GSY/XVcBbk0oBBC5pwo5puXLaa425xOw0t8ecW2GiqAjwcJciWj08hY+vC
eiANyOeUr3g8MXognCfXFs4aKHzQ/biydAixY0bhXVvJibibgt78SzPVY/yD
33xUAXoUEsCp8tholp2Rk9O73qvaZnxmJj96SND3E/zZW1ppgl7U+Asb7aFa
8PoXaB51uVxcrE93bvoeu+/V6Zi84Ib+9LmQGxA2tKieKroT92Tf+8wXAfmj
p7aZnBb6omwlbuPUapHo6JM8vuPah+2QUnd8Tv98q1PST+TO0aZXoATAgLcY
UQxNjqdQalyGwTub9GlJUQ+nW1m/Jn7aFO5e481Bg6PRVI7UMXyfiLBmnbK7
xNeJd6s5BIpE5+X0k3F9nbGZE2kYtA6Dmi2qsc3435OBNmH0XJbxaCr95KOW
28izi2BiQqBmtcq5j0P9L8/Bb1Y8h5+1PRmu+BFuoRnlFfJFjgunwYIhJPPI
rqrCVxK33wMZbcGln39APbzDni5jMbWP07wkNN1GxjKpjDvLHf8G4sdhKO1w
QgWtNuJrtOxhzP97tu4dQL6UtjvMLORWOFNSNoxLD6wZ2eYm5UmPOXWCc9CC
JMk/Ge5ybmGQ+vdQomGRSRVlwjYx7ahy8XJlKOS0UEUOaL2CMI16KOtBW2ae
q6dlTAPV++dixvbFdSGAdBiCtpibwvsrUT0laLZok6wY3PN244blBOY1eERg
6dgkXW++yayEDj7wuqgm583EarWkHncQlo9PrwmI+ytqD+lOrutWkDnwA3r/
Y2R9iCJ6ME80skznkGGm1HUDszMKbJy9eiSMKEoZGXgJWoRpkwg4jInCneKm
guqBf6rzF3RTD74pLlFkp55PSzJYwMs9/DpKBzY9mLlQhG0HYsYIQt+dV82i
uPfT4ney97O23P3GqXrVW8trepPCoqxvlt6eeSNqHwxMI2Z3RK+XhC1Xe/pH
7r8ye6mFdfVp5MNMw3zT0c92+n0HVkxSZMRv1W0cxrdrtT7cDX3iFMko9dtI
PIbIAe5ACIinZzqE5EKctP7yzBLjff8sfTMHbwB2shxWBlnM15/ZPz6mACD2
etzSBldlD9KcI4y0ojtuBNpT7dhxq39aqRnknxQohkCmFcil5laz+bb5A2nA
F6l4j9uGB5kXrEEhdWIN98ZEsAlHSMN/32YXl5DdaGh/Q/8yE1hYJh1tGc/C
yxwO+gMO2Kh01sj0un5holZ88vyFjnMsZPiPzqLFsFo38v4nKEvkCElu2mLD
/wosV4H0FGLFBcQY0v+LSGKM70O9kbFht3q3nNJlZYzxBIul8FZ1d9Y0uv3f
a+jqsXyNT4qWfnyYxVBgoxtXzFSMoemizUqmVg39LRDrbPSCoKMaUYmVpHrt
UKPpN2d6rzSFcHKlLKa02JLVOLaoLOokPPfd3PUORETIdL6pw3bfUF6UuHS0
wSw6ZR41qJIJhS0/CIcoXd3ypSDY3RgxtJqHxXKJUad4lX47VmtjcEwenxPX
qCXXXQ8/3/DgmgTfbhDnx/qC95g8fxviYpRDkWxaBYN8ZkwDr4XXaC3GuC1p
U/c7l2VEN3pDfK8vCNyRSGCQfIiUkzFAOj6E3Odx1jL+Cq3uCVSHEG7JqqeE
EHkqWEhEpjc+e7/Fth+vYYBQ36MKSZYBOICNEQYNejAhSCAqcujWgTLszyNl
/VtAZXIxSDlx+eMYg29ErFJnL0FNUC9cb58UfCROkYf1orabihY2sB8NsR/O
YYGKJSN2ZSVRtb3lu2uPHYT0bXd6N8UuKXGmJ9pcM1NduT0yazbDM8TqR367
s91kC4XQkXGT4N9xfvfjcE/vx5I9S2jIg3wU/C2zwAYoLaXia6JoN486O2AS
np5KpXL0VSHK3nEs/T/o43QlYWfIOUUgcVIZDhgod7iAm/tVbmt0/W9cN2cO
XLl4EmOuw/koAAYS3vUTyij8/kIjSBIsVh5mdIFnsx60hFtnEHUuUzyb6mX4
ju0vcp9zZdTCobfXRusP+QbmSrUKEzCxUOocnywF7x03zFePeRD2ifBYxbb/
rhSnavkNPED5JgrZGlPmnrVyztbziakJfBdfZZKJLiMEQ41N6pGL6DGfAfha
+fH52mGKksOXVQeqo1+cA3h2tZoL6pr84sEZRFiJ+522SICg7XtSgK7X8C71
mCTk5v1iPxHHhqLDObIzLHrwFS0t4FSJQPSmq82fX6Ebpy6K/9DmYLFsDFtT
Ip3G9szE4GfuQUBSA2jUWlI7zLsqKHmFoJRHvxRWqEiWxW2bv2fX95LA/It1
28VkVfHeY4wh78c9aJ8QVV2NHkwpSz3540bOWEwMOUfvesyagpnTiRoN+bJ1
+2f6YVTPF0VAyjObPBoZgeDnDjOvzmSj7yLr3l86JpV0CTD2rSClR00XK9Wa
4Y5/om2qamUgvJeZB94D6AEnlt5UwiUznckqvRdi7CxlsNbAV7KHtS2EnFyI
4YkJvQNIGxUakVNQc5F7vSAghFsqrVD796XLtdTVIorDgFURC3dp677WHaia
+2GU3GljybADizTipzWJNz3FTGEZ2v7XZxQFPth6uFZOpIBTQ3RG6jb+IMrA
gAjE7JYP5SpceYKyLHdDm+QgKjZfGzPQJZ6ZGdxXUykpjlCpyPLgq1hfk5jY
azRX4WbKmhnAnVkKrZHSFFpBttnAnUX2FkaU7tP+++q6ICP4hO3++KlbQuii
sU6p/Sc0QJP8Iza/tMURodKtkdPcn47UkWrL0q7DqjaaPSYu7e8kI1EP/g4B
sENJS3pJzERu7KYr7rBjerWYNnn/W20dRVIHymOVbxb3E/FX5g9Hw2TiBnoU
HXVJB6AUFQy7/rMii4wKRAvVoeimzqgpoC/tv+7SN+9QB2PR4Z9Z+EAi+6vw
mv+WVD28hgqd4ouiKiXeybnya4bVJG0KNo8jWthKl2apO+ZwMfzeRhw5JUNg
4ptnJm+66tUxVtMeOP9H7rDLqWVf57zKKxdKm+7MHh7csDl3MVn4BK6JI+rE
lonGMhigc0mIY7R9xlq2JD2jlVufVpqK1Dt21k2ExrEealIv08i6vgEujOZh
mNmXfm0nxXGM3BtjSruNP8GQaB4VagbgamphP0AC4XcljVBfVuS1+B9ktTgE
nmvcjyyKbbqFHebLFbevynIPQyp5Et/AtxnM75BbmXY4uKXL4HBiYZC3ilhj
tiiIMd7sxgI4B14jBddqHJH7lM+Key4SEe7uvXYCvo/1fCDe4LQ8RfP0e0LB
1JcgPpBtW17w8R9ixdxu3ub6Sbn4zHtnTd/hvpk6wWlevMcdxdzW9gnoinja
ZCRAwmjpXLfmhuhF840McToWNnCAF6Da1v15BU/LpUZ+yarKwaH7NcGfR3gW
sYgd+vzVFaq9u0iuyLVIN+vyqHmt/xoW9Ilt485YuV2WmleMBhFbaFdedgTR
hMzioSeQj8VnkLzgAQnrYe0sjkspytQKyYXNR87vKXrplaVtBDM0ekl3hFZN
G+aClYv4klWSuk4VG2R8iHTen3fKb81oec7PukSbO+xO/IKjGGYPabuzT+RY
kNDv8AP/gXUwKVuBK5XUTKNhIqDkTvVPPG1C1FLSfhykyf8rv+BvyHduxT/p
xgPkTJ0BjKJQGQ2j/acsTTICXc0hBfDfVAwNkgYvzXT3vBRHxZ2XPaFtD7f4
BPG0BHJoM4WzmiKlp4FfeFhrjIHy4bpFMvlN3QU+lq4A5ksoXJGDia6Rfa3P
uUEhppQRoUwk0SYXo0ut3dVQ5TmCX6fqGrfrgKOAe7IE51+KzmcLOM8r+OHR
JdhzfjHYB1seRswJHvtJpkyBobA8Hf+S7gb+5nLiJCrfFKVYdPP9Nt5lyt9l
y6C2dcPPteTmwES7Dp6+5R81B5BStszzTGC5lN7vYuP+TNziUfb/1+cERbR6
Pp4g6ZR9Vf/zocjbqZx/5RdNOAla4PUIKhww2vk3N95tULkO11cWz+FCgUIo
j4rMfyfv9HkQeYtF1Pv6hf0z0Cszhn/FDuQmtwQnsDi5qKdIa7PPvSAixV11
UtQHJvZ87Nhsln88vIurtZf9Mtn0DElFtd5TodyH5VneLdMWBYigzfdieCcj
Y8AfLyrpYDvotkPaySJNn4Iya+z3lKx1yFuKUvZQubaHbH7y+qg5VWHlB3P6
eMijutbIsTTWmxvsvLRBidvY4ar5J1GU6sgODukcbQtLVXTlnl8d6F/nO930
qPhb3LZh6u/PgOid6sHX+04qalf6Mn2iJGkdR8Y4KgtlqsdifPiGbPCpjW7F
CDgQ1FfafYCJct86vsSObxQk/P8krcdJ57BPysCDpbd0Xa4IIox18IXLAYEw
Ia9044zpXOXnoqlFdDa4IvrLCqiuUQGHDvcFGPoRxZKAV52AWMfCx7wQa5+N
bfwq58c+SBRlcRopp/3OuBB0B1A0HvZN3rLN81aJFVKnWUI+//twzfjIK26Z
Y4MU9arJbc8LCLoZjM5atHEm3Qbb3rqo2jB9DLcsoFEQJohecNg2g+G2UEw9
asWZshSY8S4ora6nQfttqa19bY1b1EA+Cvpu6yPw1XF7SmHtxyYrDTd0yh62
uXqnTv8Fja1/k7Y13A9bWj1vNiTHixTKjQw/oYJtiEEK+PY0z6H4SIxdafr1
rBEMm1SljZbXqHSThHxI/L2alsreOYKMqq+uzEjw/vyT9+WR/uQ3q384sRVZ
bpmsbdmqWORcVBwrdUme7ycNktowX8bUUx8SCSUwqEnpapvKHvlhd/slCV4O
sPqS+WYIg24YqoAKlDBvHLnlBdDJA4l6oFMRXIjSoLBQmd4HiSKl1VvO2B7f
7vNOSrNbL/U42ku7wOzo+OB7kVPueNHxMdB1oFDgbIp03FOlyjYU1VdLGAnX
rXd7HWx2zsSNqIxcWN1Mb2tItA1wxv6t8Csn7m9D5mXBl8LI3aIPy72PmBd8
96rvmEHtxyQF0dzNIBV+EAYavHvT0RWDJUnYg8m3rZnw7tPHJi+rVxYLVbMO
62kFuaZyE4j1LH8KT2rg7twJjua7sBEarVl5qEqJtbpWle0haaJnjJHQbdJ2
/Atw239xYzA1pbuDQ2xXWlN9MgsCVWJqcAnjB2FZ3xCZTKwCu4xl6LfpAcHd
kEd+mCYLaCb22IvH3lgH8BmqwMSeTEwDTgVyklIlno7jBdiZyLmcIfWRVBev
6xYEpYgsi9tgADsDzelD9I0sObC330ig0fM5RSFJvkW84gc09ngEGci5vcBz
csX9JXecAwFN4Vb59iaWAqa6F3zRz5qPEPC300Gt3iyNdrK/YZZnnYr93lq7
mGwl8BnOCjdqOJdOewO3xKmOxZ5095F0/pOOUZbRnhaMuII1AsMlgnOVQuHV
2tLfyLJ5fkVn2+s6L5YrXJmp46VLL6cC8bnALN6S/0nx0rOL8N0evez789c/
rUAA53rh46FHlq5UfbhuFl6SZ2bf2JgC9O6shNsp91NusCDi/avCg2xIFzHl
Kd9n2LEi5wY1bMmLg+DcRIwBv0+DFG6TF4UHAjFFlmi54ZQVWUtpi0Blr0YY
TujYSI8L5PShbXCKGTOq26HD2lzpBn/Ag7SPwW/WNATq3PLP7Qe9PUO/SOJD
iFbdQpdPlJnkWmLbWZrmQ60Ac0mNkAsn4h8FIU4YsAeM4+3DtdXkzImdDopV
ehhoWfrHn7CBCPPydReW4cbBmbfreaKew3VzZm6A7DYSwgjaKDJNElfc9hO5
/VD+eBW9acIgqjWXWse/W+hN7UKs1r+4u7SAPUGwBhHyQtQMk4bLBTQUVeUc
t8FbPuiR4xShOYW6N9huMqEb6u5FfmWwiXOqFMniGsmXnjDMzGZ+wW6LbS1N
bwbN3/3EVV1gznSzk79NoGFhtGXpKXK0J7FE9ivcMtls6gpj5FNvYnjflocY
utCPU4NA4+fMdoc//SXMtvcq60HDFnLZZkaFLwOhtU3DTxI8yx/M1PKD+tPP
KUKQfviLHpTGOoDwN2PBOxtOuk6mcGOv/5Q557kbUJuYVoMZ8rilmmbVLGFy
R/ghZVkgchE8B4ld9PBe8gFT9u6H3ig6P6I4cjLCorhr8hhZtaw8607K4EdX
K1CjE2YP8wt3NohdPncdHTQ3bwZDVnDNOJG3IUropVKbcEtb8l+JBggxXkqZ
MEJfO1OZsYu4QMgzmt+IFr6E64EJYPU8RfhKHySYhDOuYTUg0eBeNKB3FGBC
w4BU96pgQU4J/djbqQaab3fpPBde4GYAwX5dFNZxr5TB/KLoULPx1bHIrVVB
QFWx9sREqakkpOjndMEY8jioKJsk2hq5cdVKBpVr94Tx4GZ091CJNmIv3/m/
09pAAiw09UTIRQT08/Na0kZ1cKNx7dzI04T6/BPgHdvbCwKqa4huICiBi9uk
gGobpaK3VVvdIIuN9veRntlRueIy+1o/GB7/R0dltav5Qf/lk95mUyijg26W
z+fQgEF20UMqoc727+5buBsw1A1LsdfORUbU75mba8827/2+/RMKUgrbdxg7
1gnbLvOLje/SXbSmaLubt4a2zZMEyY5GgFYLjkKkEdIKJ6E3K6d+H04mND2D
kZ66YiZDKlOTOWdKZ0JAXIjEWTAkQbQIgGCOmF+N5zPUkJIv222mPrbCIFOE
jrSmkNAwLlgew/jzaVJIAylDzZrytB5v882d5Yro0nDF2CqMCuCJPgdY/zUs
RVVxX/09eMDzA7wnLMRP7rMBsXcyFr3xiMqr+eL6FAt3blvoQfchSqLbn0KH
9Cfz8Mmm0r1Vlz75OYykyaFn/4lCXCXzZcq31LfP3vhiMpRqodWn6EzE5SUC
WwMSiZVUt0+gpT/Bu3wb63pwVtTbluW2+a2fejtj+dLaiNQfNMEFN72LxQOO
ELnNU0AsJIwKrD8+XClsOQuAGL+b5H0zXHNqmGuYSERiDzGqaLmJuxbRyZjK
AzvYPEvTtfCu36fwoFsQ7AiMS9qmaEeQVjZB4FosjI540vaPjyfj7BhYVSnH
Tc8oxWHKqrI/vj+K9/1oBGu/CR5/+XofcbK4zJxBbKxNgPO4/ztLiWZobYuh
hgdqkQCjBKGGVgVmAshw2/MrgaDqcC3azoamBk/nGGtEt0mcrkky7Eh5dWWv
mDSvobbAKvLBFfOxinsvshxcBHVYcZVl6mpJFQrDf3Ao4u3S2qHUpkeXzauD
BOQrc6AyiFHcradEZLkSqDTmabAYKk7dUZ7dEeJRu+EpOKeclSvW/+ePX/lH
AWjE8s29cVRtWTGoz4Du+fCBX5RFta7sJYoJms9HbrnFy7HhY62t6Ln/Pe18
kTcAPQEDMF6ZpTqoTJswve3giqWdTZS8mqrKKWunDFcyOV3iZQM8Uwcd1/Cu
G0Pom4NlYnkjq/C2eW4Vo1sBrFjGjyrgH7HCAzdNCSJ7Sjxiyggv1KE15xgL
kCgzFji+sAP1RDsMhr5/7Cn94fJ+YtuWF5/vNbYFFMyBRRwZhaCHiJPbDXYQ
q7dV10socOH6XnYzsxuqxPfSugqvOa/fihXoRg4mV1S/77YTdJ7uUsC5mOoi
G/akpm6Wkl1PRUBcNrPxfZ2L+lId9ZrnSE86OncctwWhBw7QrrrxPrtmTg+n
+wul/NmJWIYWgO1ARnADFjm14t9Qk2zYnrnaPHSY2GE7r+4wNqIcuBU8FdGJ
R/auMeJvzyAzkcuZPM4pqbA54W3mPCFzfz+GVgOkKh+zOz8B5KZ8/r17x+9E
4SBYjMW8XXP+09sq/aIyyS3UMpwOdFvkSmtz7H0VKLb8mK3JMreVKZykxqZI
xr/R8gtM+af1B2kftVuRFGrT/xxhUvYjWTJPfJH5W6R6MZKwhPyTPLILvYXX
Rqw0BuBD1SWfuhnA5sE8qASxm9cvwG1U6F/5JoT0f2c1Fc1yh3AbazZ/UZgI
+CrYEv3Mnoeb2wZrmDY+CqOiD7Q5gs+6ipIMx19MaRjKN4eZ5VDsxxV7d2XJ
akmrqixAJRjJyfv/gwXPmVPfEzyw/EfRwidLPvtIj4mUpfbvgUMd4WpQWdul
LDTTAhG0mvHNK1SBMuI22wb4uF1Nrt9iLns8y0w0yVnRP/amw/JROkNt27sF
fYkUBdLvMQn23Kj5L99VV/UrKL9y2QteH6rfR14gexsxg3QhvXqYdejKs1AR
gHeu6z0SXh1kbGiJdZOyrAK5//qBetQ7L8oR4YNG+cPSW11s41kIpflkVGkU
QOwCFSMTK0m/9X3BGFLPyiF84fO7iEv47zAeVZdjZ48BA1lO4grTa9QI3zZz
8pMCZZchJPYXbkQ/UWhGThvWt3xvAQNog1LZHT/UDTF4qUxIABQusaU7kmkX
exTjhYsMggaOyVvtmINHi47BX06GFhP0BdynWpQwT4I2DSwsq8B8MpVICVZa
S8hIg2fyb35W5j16lyiKmzt/q96XRwvJZ8kXn27Sq4lYzt8DvOtzUtCGVDH8
xsjjAX59lm2zpXt9oRPAr77eMAbsfwjhPbvTFg8CDk+Mu6xV1MintljN8/IW
Z5UNY9fyUbTsJUlG2oR26Zp+1BIRpf9YfdImC4WqaDuZ7GHEypmaV3HBYT1E
T/G6siYARRWBhxX048dH/oyPAkECBkUQmjU4TM8vzITOPlm0OXfKb3IW1O26
YwWx9LbzOG6GONwHYQn+5wd+g77Frb5WMbmv6W25IImxG8/saBjoqjLckJW7
c7+LfcBDChkcPnWZ6yzdl2frFKZOAd/P6U7sOLZGFDTeF3GyjxYiys+WxqFR
Dkjzp6f0mCo1XUInud1fodM/tMUkZpwAjPWOTZpy6DdUX6ViG0AzksSmSgZ1
plITDLESmR1yXkWkSKDlAlCffKIM6gbRHPIEQ0uJwazpZlWySsCtCdGoyzkX
OJO+Sch9IZ4GFkhciufNaPhdnPcXA9UaiEMqeAFaEwJq+cZsvQkQVvndKRnx
Z11lIdpNZHIbSRJK5nlJD6uRDXZW/O2F9MkUj1HV5/R+PE53cnGVgps1AhDe
nEwgkIxt1ZiMAGe2oBJpOlQ1+WbrEzEXyuqSLNdeI94OqQuMKFFCgnaCi2MC
MuWp7Tuo5/L7JeL8CdwTgfh64/IQwjmLJDxhskjMNVHq8TmP3zxApbWzmjPt
kCNAS266ikO2I6uXu9aH5d2ebWSL4TJuvpbznnhTlZwy0MHzrwV+H+51xKW7
yTc10b6LbNsc6p4b5QcTWbyGvwOnHlBzRm6+8Xd0GitGCiK08xEawtiXLh4J
UZeAKgy760TzQRXBBzzK6vuVWJJLoLIP+Gryl9Pl6BJGqUi1Vpys8nXiXVnj
sG4P2xRTX7a8Wjd08pgXTC4MgNGeYNUnilcpYnRkZyEJouNJ1uBl11y4+YNa
i4Up2CBxJgeJu/X0Y6Xj22EtNU6seRfgkwHB7xvB29yb4tUDvLvMf3Kuv48u
XjOKF/Frf36MR9gjWaFlL2P73OtGfaDpfkh8u9X48As+uILsJXzAf4drmMTT
XM0kF2F+SwFMX8tORi9PP+NuxmjNBTEneRR2VyDEkRdplANdsa8LawHY0CpN
vy3bAmDE1B4flcfV5OFaWSTas2MNAslvEaIA3r8U/NixMlj8CP+nXmcRCiS0
GuGIYER5dbFIqFK2xN+OfuskkwL87POaSWHpQD3DUElqsGGGj3KOPP434lZQ
x44tI3P+EP5h9BABYX1l3rpLsJ+IPfpGD+Od9hwGZ57wwntttR6JGUOPj8wj
0kQkRjiApin8Stjem5X64T2py+ASjJKBMXH8ztzLlt0Xl91BGemiY14BoJHS
/CsyG8howRuNt0YZO0tbV1c8h1UH90OaqphC9RAKnRzcgw1PMrBMPQsRJOC0
YFnafgEx90dGhg98PzuwZLRSjpIYoCrWubSJ0vhBvuBPRKPubq0BMmQPcNSF
qEMgngG07jCGWfudhsMWCtOG5eesI+xu8dQsXva+SyD9lEjxgrbSiYXjlhlz
drIcNAC3lwM/U3LyqbOhRMq5RBBPoK3bmuRPAXYbtX068Z6ECVF7uNfTEw5i
PsH1LLK4kf9wNxloX4dA8x69nQirG2/koT6X5dhgyG0JDMlwPdDw4baihl4h
rLrjJXmJmUg+BnhyejRM/coE5EtadjbqqnnzCBjbFDXKvMYF4rlAmrlODYR8
r+65B+I8E5OpEeRMl8Qg1OGRLs5UIQrGvBNVAj4HudNZ/v2F/HEfBZ0Bz3ue
HuqXeiw3j44ZcGP+oW7EX8kymaRkE1IefPU4MbE+hqixIbRnSeQvRxzvvofX
54EY+Zx/MCFKS2M13EQhhVvtaOIZ52j56lLmYkBKsQ5DJEaWkBgQVTUfSREa
od+ntFchF/Ghjoxj+adsMSTlPFbmpFnkgLsED72+iEXUPnfTk6HCwBxT0s4w
+rq6626sfviSmGz83FEUEAvhoKf1VnbWRrlwHZ9rgSFQPf/BLR37spns4oe2
Dzmxp1LAJ0hIR4jZsOEhZXEsC7bEVcbTrQBHIH6u1vYUf0UQqorBEcAEMArz
MkJY0wuksYF96OwocakppbpcikfxDKliTdTT7q7hwTPkBHC8kD4MTt9K/M9c
GcEdZr5CUXFBACi4zCqsUJ69L2B8s8VOeQKOwxh1Z5nLTqIGpS03Q3M0TgsP
mK1llfjmiJB53ie6596D2sfITsD9NLg3V87aIHE8M3yu2IhPtzWAaG3e05Ux
Bir/blIIdECcHWwCeVMqpcZsl7/1gj/0VXSXfLZfDwAFqUDRIAyb1niEn4lT
ISPJGi498TsciHNjUZ9HyEQmW0tQzsbJM04cIO1+Da4KUyji1JrBzHWP1OVB
f9L7fX8Dvj5NuEbF+ly6EiF2pB/B/+RFOfLtbqLBiUcLaWuiekKGgkM07aJ4
4RODUCUizFmTvZpbQkZd0U1kCgdG5WjIs2LuLgMmZu5D8cLWuaSHSQd0cPRY
DtcXsXaunBU+oPseXp0rmCAWQ2RQr7YIvpx+rOUDndZ/uUDoaUmkSVMshIpE
Yq8y+QqAJA2Cxj7+LTQDLQHJfGXaAfCs0Z99XkkiLRU2CwcwD3W44ManxlSN
qGFE8U+ynYGPhmGroRiDqKjuoFZ/kl9ukKS7A6ZsdK0Hm9/+mXeNSEy0WEUh
irndNeBiL81Qvnf5gfXr8EwKyIIhJ4zAwe+eeouhLgx3RmqnjF+AAE1hc+oV
3FdOLNF7Z3Ba4CM5hkZIArLHzK5Mmg4wHdpjToC8XIZ96kCOPuQpXTAeILm2
jL4IXWla+w+3AhDUn00jlGstOHj+kH0J3h6QLWbUkK50C2m8Z21FHte1aeso
pj/1PpRC1CSIr1oBNbwT0YycclU7iJ8qpwsMvgAfhjVzOqEaNFBcEQtTMQAx
yn1RRrKN7CX6sxf5nuJpmtGj4CNS7xSN13rELvvMb2aiB3PlvXqb6TYIzqSR
KRTOk0Z2HZI3sffQ32zACtbJ62v2bVYCWnjUyA/1RutYqKIQCEimHAnDxE6d
aOD5bFVf1ffZxPkT0xfgIkBr0YkDHjT/xZf/kI1VZkRHJL/v45zCqO6ND9Aw
PdQnTkVyKJTuhBgAqPavDyG+mQ1ZEcINqJ/RGCoSHf2Eembwop9IbbavZhaD
NXzXJXpm8d+UJabU+ZuxmJGGubO5uyFE0SguTgYzspkIV3vgj9wHMDmLsHKW
Zwwlxr8Hnld/GXU1GPyxRAKSJ6zK/l3Xur06VsSfEuvFu9eDA15VWE+S6cLL
stU9SDwCnXqNOmtezkvrg58AcVt5oL5EFi1OfizWxzp6gbYVNrOrXXELtKgZ
Lbp8tf9WJ0CgxA6OrBPFFXrXTivS2jn4DbxW1fsMBW1CVLb+yjaNgVRSdDPe
wcoYxvvUk9GEkpWhl5/fQ8iUwHEKkW961mY2LhrplfP6l0loyhYf8YJjzKGb
xFeNetvxIasJ4muJ8pbTEfWz31bncbR/6b7xCj7t82jbzHvQpadKKUuN8Yvd
u3jIYeOTNlofTXJ7WUHqxAlbUQwse+QGdU5WAnkzE8Lj19gjFiTL927bsl3y
aZhAIov42OyGgrI+G4A0LmEiloDoLn6/NsHAhEs5L3bbtywPUg6RQe4jO+st
pAcGMrIYxqxDjq2BGJerTR9/l+SFmIxVFt8FeXV1IBkaY+RIhPoIuHBgVN/s
ODF6TYSUEbd7hkcCwKuA6DIclveHt1hUR5zYk/6Xnp0Kr6yRG0+iMQr4wje8
h9ZX/Z8lHm2OI7F8DlR0TA32lBcC3EWWBCP+SSLeSn2PHXHYodLzg0p3epD1
AMHm8HHciAvAYt0UzBmCqwFECs+bSIZO9rABfyGv/bQeNNMVyxE6TbxJ0cge
bQy/6LvsIdKQiyvXzR9zwscT8Cx4TAnfREnpR7+8aXjWg9CJAxmOwd6xENqa
qqB6agOAtA4q1opvv1ccj0uwfyFCyDM8SCDzU0QH1w3izX+MOg6BksNNoK6j
lIUQQPNieqZIzsf2gthlTd0J+cgpAkejneF84afX7lFclxxUUkNUzsYq8KSK
L2H7c9/2/yin3qVcqkG/ehrj+HyqPbhCAsiCiBumUtlluvYfBkJUOLa/zveQ
Q9wYtBWIzGT5XQTn3bfCgzlam+19SJ3P+5gN9cLOeXsfyGsOLxfPcWEVhxgd
d6TNsgv8Uxcb3Fahm57xnMKW0TRdyM3MbMXjmIUnPlcRJlVz/2A2pv+lZdA0
omMxH26suNxGs4TROvIIfmvwTzovBSl85VZQkj3TixQx7XLviIbAVaQgHKof
Bp74s1kznkxNYNNa02Ju2PHJLLw2zQy9N6m4i49J3JnD+hvplzllfjT+DniE
Qn8wAAlLhvAqWytPkIk7lsjhcX20z84kXS/YGeJB2V1ac2fhcA8JoxgRtJhI
sjBJaDurrotVqVrIZxdIZK4ZeeTwmxf1p7xq+7UkF6dEukE2MooIM+LJDAC/
z31hNNEJPDhXdhPVHao7PRY7nWitxhGOdGXm1mjAdj3BhgzKppqHYZUc5cl6
g/ipo7ddXJh8TvyJXghwio3yK1HYL/w4f+uR4cFQHvX5Wbfs5+ljrMtQpzap
lfefweszssWZH6ehi95jd1MtMC1BiYV0eiN46jlYISIaFpxLJAZDxOH9hwTf
zor+Ir+yA7/vm+aiXhDedpL9K9bYLz9H94fYK6+zrzQKxt/OeOtegJsvWsCW
Cg4brCkf/U9bigvgA7UwRhWxx+c0zj8FC2+p5m+PdQIyshRZs1qOlL9Nd58I
cZyh3BZPUhtCp19hyBrlSFqFOcW/Lcl0K1f6NbwwA8UxQL5jxBR1ESW4uQeG
c1L+GcX2umJmHKQEfk5Bl6X9h8YmNxTUG3Kx/2k+WX/cDxEP8/6+2gMBKLco
gH6RI+bwm7vv2eij/OiPDsileQyEe63njep4dCOBmEm23CeGYRNIiJt5X4SR
K+uzYQy/zrYyWEt6nDvFMQCUZJyO+gCZiFMnEmDjG0ITfKKaRs3NBAsu8RNj
rDWSq8YoaC6mjhRfVcACao8QMNxY5ttxkzuE09pfJVSCY6CDpf1ocV81n3q4
w90bkLTzJyZpNlDc7gJ23SPONRplVAREtZW9cbspSOO54xIKV8/9i9SrJbsF
cEszbjeUKvwLcC1zXmmKxq/BTZKf/kpoaBAzUoUkxsDX7bvEcNMYZ9DcsWgp
7AN2Z+vrqBthYOKMMWdtLu9Tz9v0XjvNYhrNsLf6r3xY6ld9QzTta0/JXZBN
HYxGoJzmgEoQR3K0GllLZud1IbsWr1SI2BKkiC954xuYD4t4AbUlPf3yjOlK
vAeN3fyfCKbVANM6MRbmEndM3v1b7ilbiJOGGW18cHV3vFtVeBjKypf8kCAi
uSUqKFsTJjaanc+ahVIoGa1ujUaYyxu2Qnz0Ne8pZF9O6VppHi1cxRyvhNd/
ODChykA6LWGjaP2Q1XPaWpHLPcVhY/dTs83JjOVCyfLvWtxJfACpnJZw0sfo
ADPo9JIXJv1uBE5EVMn0UdcTwKyo/7Jv9u8Z3wLb3VYLDmcQcxs1K97lBYtl
eGB737bJ5pawd3wtvFR17drn3l2qKQtbL39aX7qFbIhxHgh8zoYybQfaXMkg
nPfubID2FaUJ+YXEl5sjtpNClU/TeWr1EEt0vDS0+UIfEKwFKbys7zsRpvMP
Ya7y4MoI7AeXMlH1bWDq7xquy23NGZPhYRM1LiBy+f3RQN3ZTNrKcV+DrV50
i98CpOdhWeQ715RF7wH4zp1+ae3thHLO6iXio0LhH199vsMq/B4YP/cQtIRZ
CKZAvvIaxVGer4ikIKAKru1xJHqVih0IMQDsEHY8bGrGt55Ixp9BDY05CGUa
Idj4UlLz+TO7GAjjSReFW9gb7h+cLMt9lbbKp/nF3wCOfOhZFVnliOGnvPJ8
1tCg52p6Uu9EtejSoI3jz2EeAbhyxUbJFSwG56RjK+5mdz6AwIdZj7nKPKAR
xBRK5YHpI5wfDdUsaYRDGYBJd8vccee/lR2q37SIMi99Tg2DJg2t/OZE8SDz
DegMRpt4cprWITT/E63cw0/HWgsEDk8Uqzr9H6T5Ex2aUF3yVloWTh7+VhPD
XU6lqFPoxtujCTWloK+JMocxkj7MWkCLeTvFrjkF6DdnVdVyC6nMwHUpARIa
v3cQ16ppgozyTAnTB2yeO61GY4sHv7igEkk7/Ot2hhqI338Fda8QWLo2pV7D
kzsSbEab/rC9glwJKY3U3yXcIB/Yr/sJuQU1G0LOch2SSeABLxpqrfm5tSBk
CWR4am2yTS7xxOSML+VZ3d04hpPKZ4J12XIIJ6cYKU2QzwFk1bcJgwmZmp6t
XACgjFX3NqqPuJhj+Se/n7WEfhhazIasdU1OAgeM6qJ8n6hy3cxreNLOOkfg
HKfkseQ+X6Th8eNasj0a/z0C+q7LyOM1sIS5VBjc1aLz7IaUxpm75qnPo4Og
NONZSAGwogD/kXqiXDRQdxOGUACNJUxhS7sIxrMWKUUX2vJSuauWUcVB6g5U
vG5zaJX7p4164TbjXRaOXfsBn53/6noh/wUeR6MUMfEQBKlTuK4Om7r2zad4
73jsXeQJEh5y0scuIxLTCnZvfTvxiE7Azh3he1K+1XaPcnPO2l0MtQDnlYK8
jvyaKVhDqijiB8RGLbOp8fee7RzZ2MBkg7+Uy9HYD1x2p65WteU0nDoljehB
UaBBTtLmLtSEgBjMWqBZnTIb4thvsmERqMJyrAv063O80VkIuQ8v6d6gJl/W
3RLy/t7czXvQ778cPTJyRc067VI6eh4mGBhVQW39PjX9EzrK4JVOpMc9alIE
MK/eGAl/ZpvZB2xblxgm1BIvY8j/yOPUlUvD+KU8qkcuXxy+zAI/6zLwLtOA
IH4fVPau9YopZzJWufoewwRGp2++L3txpdMXp+PCIAmzg/sQkARRDV+LUnOS
tIzjFTt0oCJ5GkxyF8RE2t9J9BAww0kOxNYOIuxVkP/6KLBwQYQluscpeLsV
zDYP7oso5PKMrvLN2RhUmIlxMofb7xXEWPSU6lbcmkHBYKpW6do7mx54ir4Y
hF6bpSAehtcADGDCGrhCXQenFEecGNzjv/b05u72uDoabKaJjlhjeHBBspMg
fa24IHFOy8+INzCLSYiymwSEqTO1pGQGtIsU98nlPrsTT3URakO6e+3pcNSP
j77pWdw7uRavG4rLOXyPOj0HNbGcKlnyLYATsi3QuGndsP6rmofAEIfZCFbU
ATTkWpet79plMQouC6vhh8d7ryTZzhX0ItulnXyMOU8Zqvlsk/p66wZeyrgU
GfPB5dBXw3DSIp0T1FIhw5IxUgd+j3WSgWCXzxXWuaAGLyi8cFYYOkmoZBjf
qhzlND1wi5ZVInBTZGDJy69PnFlejiB/UPvuvQzWgo2rFoGPS2cV6gXFnkcT
3FwDY19KoQMa0ybW3SRsOH9gMdtlbT2hlYhYXLVdzBofMh1MUPx0R9kZU8Xo
JfCq3jhTMi9LNYKPtAr9BDRKQKeVJvzI7aYgh45zDW8QAVQguuBSCUwMsK5T
9Gae+/rmsRD4jIVPG0c7IUGvbH5BdBxpykm0A2flF4gH1raScsiw4i4nMzy/
mRGihydKQLzLoiZ9bn7iUfSATG5ITh6CmfCjaUpZhkd4AYMLOjz7NY8jvG7R
ryrFgGL1UhIcp0SNU4YNl5qhk6eJEU7CK+BhofbjgymCHOaWDZ9i5AXP8qCQ
i4hQd8TIXzVKZbCHxRlwr4VqUfUrZkuJj7kLH8bN2lCgCB7QYeBqdxBWZO+Y
Pxtluvm4T0tSFNv1QP6gGAp+hUz9r1wiH7l1JRueIqUccN7YHPj2ea9N4sTJ
Ef6Rv2RfhcSeY+LFqimXGJtouYLkuG7B5H0016DCOULOmeClvqxCaRAPRnz1
Btd1F45AbQzxcdyrVQiv0heZpJ4ziGUnOIbJpkhPX7layFsWY0myJkcGR5cz
9k6q6bqJuaoYa8xyEr8qpmyLIi+x8txamvzDGiXdUNMctWXG59xk8MNG41LI
ePkE2eCQMc5manPAGrqcQJeVlKUaJBbQnscJ9M9qGqmWXnxXmzU2LNCbYOqG
QtqCC/Eoa6FRrBNNZs3p5ZPUXk2HCVLXbKritTG4+kOl/ZX5lkGNcUcGiZEw
1DpajrbEIog2SptinO7F+TFf9vg8HlAZ2IHDEPdGTfqQ05eR7bL1e+vOYqi8
aE8ygTSxeU1Q2e7ohHPAU99HJsvt+WTAMJYJjwY5vM0iJnlAJpecWffItvGq
UlLuPFWFGOCX9B4wt4VSpELHLMdUdQB1lAwULXmUOFkunbIH+H4RfWbxWLux
ihf3vs49Py+phdQrJR+RjTg8beb/inYTDJGvJTt1bfu1exIm83HZJVMEYrzc
FWOpl8ITWIy19rwCuvoWLc/aWTjkUWZ0JgxsOM+ZwIP5oqFFVaa6e139P1S6
YRC1nbbyPbFdvE3nEglpjIqiDENJa/Ul7QSAToUogxi1Dttof/cFywYyUBr7
2DSexQbK9vkpVVMokoWVu6yah698xG5uxrLUxlbh9DQSBdpxmmd7cg3m3QQg
WozMxu7kgm9+JbzvWnlg+3fyKbXi6jfZF61MfZpmi8pAoHolCpZD1N8dB5cP
xsOQs1mb0xYq4zNOoGxkjr13JdtSTuIbjIxWZA/UXLN0q5XjiuUdImWJ8YzU
Agfd2dp6UzOyseeOYmI0Dw0wW17qcm27YVkTP5XYEoH70SDviUOsuiobUo17
UY8zMSozd2mMmPw7fzOfJz7oSys8BjeWiTfWWnTHGVbG++dOzkqZykz16pQB
g47Y+o9cdaZSALVg3Jmd5ay8xnxsrFmSvUCbjqga7300erU/ahIKjOth4vKg
961cfSKlmEkjyBGBxkA3HDvdXPYL03euJHeTJwqb0dIuxIvfNY4FFeIwKx/M
3ofnkKV5zz6osNv2Htwth4tsyFMFTNMR7f7P7LCCFtJxryhE6fE/IXMtaGdt
YO/R0RmXT23YXCFqb17a6mk12C/wqrBuvucd9JDQWExCnaRm0IZ7dfpZ8AyF
AVEpBjW5xf+w1i2rd7kceaxHJuabS7+Dy/f5xjgDbrM7VvW5bCoKAP5dRpJ/
l2gJhl+8SMVZhhPkclKW+/H8WL2NrQWTrbJSiTleLvp4QYmg85f8TfiF+dIu
UpNLqApvvqok/JmRdNmVOc/YeDgCWWdGiedTYkPajUgcwhPohmnc1Ph464Lo
8IZYom/SROCv+awLGFNWiDm1KVaiwkk8SDGBjBsfG6s2tux9/fO1JBixFqxb
lD+seIXJ1Bon3VN9GMtAc8TnTcWHYfwoZGdvHEkEK7nmS8IE88bDE74arSdm
maktszrJPpKI/we0+UpJ6saiJEMSwhrXr+0E12EKOxFKpBaZ1CwV68MV1Ijf
S+zu7FD0ymSGV7aw3G3VUz1IjuewYtL3tVxlDf2PkoZzRgjTZk1Oi/brS/LT
2ofZjsMyUiNVF9/mJMQWs1+ZvjNjISCDxQ2RmBzqclr0aV3LelF7SDx9TNdO
gTqLefVhTH+nzhwZUoFaHvxP1kt6sLlsqEgtR6NrwbV3MlfbCP1qv8690aNu
b4bbqNCM2InfiJa35NgqZaMYSUReOnFKQEI4DU13xHzHguxTpCsAK23kqE8C
cAUul1LYsw9w1Yjlkwa8g+YoBMP64tb48m3vOvII2VGcwuYQrSS+0tgaLSY2
0rPZQ8MoyxQ0LZ0brGppEIeENvL8qBJNQcu4LEN7O2uw3pLwk8m8+5kz/ruB
aOaR6QCuMXB8mPv5Qm/JlYeNUEmQJWgNZizQ57oVYD11aDW2neBwM/f/3XGh
TV58yyPaTHO6NOIpzSvczaazlkWtIfBHqNsae4aoLwjXlccnbUPQTlAKslyj
wGxokvaSAg0xYn2RNK1vIFgKe1WLHpN8D43OnTKs4TWSAypFk+kw4o6ywKwy
4sxwtkJixx5KoTNZ4158VfxZGafVzng3FFHR2jFlyEb7DlIjhcywzu7VxJiv
92Uftehfe2OTE53SfFqacTn4sSXJjtH0bDwfneQ6ebtetXtrp0tKCetQO6n2
rO8wIiSqdbdQUiIX29vAybOnJ0R1iYtpM13FuqzpQV8vz2iFzY1CzqCJVAop
iU8Mcy994HI7j+I11ubm0MMiUtxM/BLmlPiRUuS/ConmZbnMgoRk6ov9cyVp
d3NxDP8OAx2FrgKQu8EIoK8rGmQv7F6R3r4QKIir5Nm8+n+H2gqA8xv4TSoV
nOe0gl3dh0Sp+JJ+jPWCPDQh9UduJxMaw1sCOt7vuhcaCc5SQt2Tra4AGvPm
SSBQTHp/9W9nnWR+WJRNQDHyUCsrlB2c2kpZroSL+UjSPjln0VCmHoNzxchs
thCovlwOxExkiSbZkEeleoheBGEKbHwWwNWi0W+vMIwvyRMXhf705OsO5aJh
wlPuVCHtLoQIRS3/SFB9tR7aBktZGrwHdp/kyN5TmAA4GIfqYylk1ZLGxmso
qlU8HJJxci1YxRU3AhbIbvLE0hL7whRB1KbumG/MV4SiUnRyLoyo8qmLXG7p
g7zNEJGrH8Dnk3bNYS2D2zkMoNrFp7WIheqioVJqxCVnH4595wiTSa8KBgyS
/vNUMaTrbOa7MxE2JWVjOcxfI6QMlPo4+YmupKj3avpVh+TNIImJ6RtNkt9G
GbYCbgiVwu9jTKa8VgSV9ZLwNkYuLhZCHUjO4gjIFd86IB8v0Au+TLRIcF96
QdL0+m4viDVWRx5nHMlAeezYyuxVpK4sQQNYhcp2zb/MuHu1umyaclqISV/g
xNGS9sWW7YIdDzfflRQql/RQoecTxyz0nGQjAA988IdCTl9kcrS+jVRBnvVi
6gtqsknXdJqncUCwrBl9s5sqWsVoJe7Vxhr/nt6mVX/W+Ags4hafBQqXIKbJ
JVGTo8Vvia8t43OSg9VzEP5TEcdJQ3nt34JceVxEOnltY4B7iTs6WH+GSoji
vyJaowrA3JdHCwS6XQmd9iSotGpO5cdGSQlyI1vROcJSJ1djagYGZQHyhiEh
4S7D6QdKoriMPa5D85D+bqat2YUv0uzG+tZX4TpuFLTN/8zwwRGFeluztuqw
1ukxLrK6SY8Xqt8zF9S9ewE/gOgbE1MAXMewPt2II662OeEbc1yF1Zt/sBgZ
KeCQ/23zqBQngs9eNRVA3OLwmWhk6u0kYvY+d36EVxc9P/qNbuo7cZRW2daL
bnUORAbsEgPff4vPmPJ6INy4lREypZIrOHwogIL5zTE6H3+iz6SSM667ivbf
JSShzcSAXSCIcVy3KwbCn9PcuNZT0xZIeeJfBChHu2oPz8r/qrWatSvOkr9U
LUCZ7jAUn0FdqLYxeK8iikEFqBKtgkLIIqxan10aaoiAItbhdZSoYXECMY9I
eoppnu1pDOx53DAtyyTEAhCGbVvDCdZaLrMhfGzpDy9z3lExDCcypuE3XQFB
WQ/pmtoZncOVxSUBt45Wq+ZPbjp4FcOazk1F79kN1McPQy5WuRCU9zC+czz/
eWpJjwXrU2y3l9WBUhZ4bq/dhvxB/gjUY8SGNKDu9DrYpo+iZM+o24dvXspm
wVeu6UC7DaB02xnQvqHAJPp6+aeuaKXW1cV1whFnVQflxUM+6VBPfI1uFVf4
CLqRsU5Gki8eEI1EWDouF1xTdF/8rkhkMDUulfqb2ZdkMSgwYQvtdHt7ewXd
2MV2XVdJEkHJtZz8UPImlS2gf0xcKMJYq5E+/XOrq7NC6qCz90bmtejuaZPM
c01FgWdLzaOydl6WFQCbpa6M2mmxtD4tKB9oEn+HqQ1ErzUcGqgdGOtklRIm
zf31feFwYAgE9CQzzYLiBORkoidgTe+9hgqeQjw1jnqyPI7GA972mqjXEyxq
VUrjqCcmzrA6EZHTqhb0pIqC19Xtf0z67mx2ZPe+p1uHA1gartzMOj1d/9ty
OEETj5McQOtqVA1AYYOQf8SSKmvcZ6WMo7zZE8tDPYo1uW1pDLjbS0QbLmfJ
vFftySZ6/gc8kMz2lxJ4lPIW1j5+Hp2CLKrquG5rJlw8joNuWk3MZ95HqIgK
2UA5gomEWoa8CMN1CHGTiWHs6kN5NhCSSwA0gLsn/IZ/xIj8tFQEfCyX7ilA
kSB9aGXjYb1YcIkr6PDMhPxgsmxesWIpHi6YTq6cWuxXqjoGdnWbBHvmftJ/
Ae9PrCPOTEQlfxFA+xpfJ91zBBX/E6r/N/qNHzZ/WiiPCozltqVxfi6ua2KI
pqOZ5HEax6NFCw4dyhm8s7s84bprTRhE3X2ksxB6yy940UsyvGRmDKjUuRJs
2Iqa317KBuTDv8PKzpUtyXYzLZ8Gn1aA15ikpR3qzZe8/fG20YAJzTA1oj2n
u8akzDEYZezOGxmtO7MyWjbTyhG/zbYW7MVMHTf4HcN800d5wdRCRL9vKSoD
4Ygyw7vsCACTs0Ll6NfMx83Ih6vbJQMpRy8a0AtRqcPFcAmBXBC9SmB4TsQo
kpN/EkzcjwPh6dbr/3bd8EtZawaloX8y44RtTpfdjwxTKHPWRAvGMHRGcIkD
pCeTi74R9VrSCTxeXsYM/Yqz6NXQc8g6fF4hqvjmmZFgsKAN0V3NhbV2DAUb
oJY6xwb8xp++/db5PecVfzYfpKvA1Lcb/oNbbpRaX+oFWIapix/OQQJrggMp
SMilOqyZbaXc3oW3RZrumY3wVux4j9fTBoK6bmZSEYP6smH4Fk7elG7peYte
ccgl1jfSk3Kvp0MIjuHjpViZIRC5MWZR7nCf5iS+XyISkgItNaTRjPGjN/A+
DycKGK2tvCDII71dkMa+MRFYmoqxC48CrIN4biD0QEYT3JWPop6S9OpCMrIA
YoU9p4W1O7GgXnmWkpJnn0YvkzIjuzEE/rxJ3xomUr7dVKyGpZ9OraJaMg5o
Rjw4oLypH4w0dPrc1M3tvNJyELaMCVX49XOlp2dkRunUcgnUlbjd34eo+AdJ
em1rgDyRYm1lteYFXIH2n7yPjX60z0muPiQWdBPBdiMjAqyaPTTs2Bc/PPoo
lUx6qNFYhne1kvOGQr/hxYBCJ4WuUc6iSCTHbt75a0p3/CorUCgW7fQo2Ky1
SQ/w2QzhgIWKeyR/Wwrbwnpe4CE4zPUQATHAKbJIgI+c7OHS23E+AZTPkEq3
eYvKYN+vjDW+k+/TUyzvhhx2eJmUkOEplc/5ne7UV8tz1qCvftXSdc3TdvRm
obQP7X4YoxAizkQnWEkBPZhpEh3BW4gei/L4cFe+J4dWWHEwA2EenkfHJibP
B6xw5uq+kxpln6HslOgr+HNDruIL4c8m9D5q1BSONO5EL5nO9IlDEx0RvXce
680HPhjknwrG2UE0KqJdKCTpvVv3K1AMbuSUnrpwKxduj3fVbrf+/VutBMEg
mvMzA5Jsrp09uUe4HEaW1SYxWpnjPvE7EJBBwBvcG08sRnI4hl6szXiwqHBM
JTxjpyWQ5CzkdOecesLr7W2YVfaStt2a66IW3wO2b3Ykdc5Y4dV6A5jIhuRh
YWeYO6Xi5n1zpg/HFjdRj2lNTqHUG8Xtg9jq2SG1LtlqhvNZVDdwB9vwhLSY
4RFUW85ke4U3p/QJC/LfPAQWlznRfN1dphtkdsVa1QctETiwh7SOzrAblhL8
dKR9i/UvEjUz2dWk7vQcuozbjLCQ0bLJSsRXpstxhI95iWAy3FtgQaLRQaEj
yNDBhk1ZpbGFgU4PPwRLYb5XX6fgvMa8+8a5hpJDQWOMErrk8jbyF80lxcpb
YJM8B14e59U7geeACDYQHAzNM7H18VQiZStSdwSd0E+dpMPiKsUMH16aPN5c
YbXsScDzDsspoPLgpqmpn/AEGnHkMOjsj/B56WmVvlyDIGp+DHR0x1sQXiM2
8ZmXt9HS8kdJnRUebBHNkNGQxjKhhJWiAefc83Ivt0wOEbDqhkzPousQXVe+
FVTQANXNZ771DZjFTgf6VJOq3fCPx0zI4xh6gMCJVgbFWJ7XDnQpMaYBXdny
vRcXeJ5G0SBiiWwICv5Naz55Eq5WDjftzizN2wLCZjdMpmkwyfid1WukCiYI
0hOOFOYmzZUGspf/x+0+7kCzMrRN127YkCahzqbJeeHsw5xiRLXelHQrcxpy
iKUr9ajZ/k3WwxKHZLb4eua4tHsFPaBz3O0FmPekR+pdnJ2IR7VSQx1RLxq2
bDwd0kFrQRaWtTPIEo7aQyutJAcFFYJLzed3DCe7w7att77I1DQ+ccX8DPnB
QYbvh0Mhf23Z3cEbFy6pry3F05bI/BzuzeEsf9DfZqWW16bbMS6Xkkjwwqwq
zLoZJcSvKaIorjifEy0MrJz0QsQM9FX1+dexoyxAL+MZkKXBMxLeCoWMKr23
+gDYeJJZTsWBkf0FCIG/qzGMckd5hhD2ZOzF7BIgg30P2QXT+TKQez+0Wlxp
Nq4kBIOjKw5bbz/GDmRIulA3qWnLdjcPh5AAnG4purOsRo33Y+zSXTwgrP/b
vQWXYwbM8/u27nSIs3Mq6yMJ67VB49zWmxrPdEvkpojHvn2I0RLjCWgiHcqu
S/fNzc3pdB9Dv5nYBpnr03oahVL5r4pkRBiG6N04BoEaEHNDttsVwkEfgNP8
e/74ootQg6AasVmfNNpYO7gRSbolIwLxKUlh5DSjonUPDIwJBXtGzF1UyFql
zrpW704JCpi2eD1GDhODhkJB77yKKFK/SDAZHCvWfmTlOPf+fvNcZAkVTVX+
qCZKqAbwO1j0wrkEZnXbOkbhN1jZwD3Ez+B9MQi+ms5mbJ7GpRPjLl/DZQFF
oQZzGwIUYz9WIbmvQ9taQRhNI7gKS7dihJDQlFyYdwl/CGO1AGYPhQmD21XI
Cj8zJFn08Q/ZXShjIDUyx2ecLe6TrpDkG8MKGAyEJ8BAansBG9zh/n5B2mKV
YKipSmlavKxdW/Nf9zQnytEdQArFAMAyBLHTY9YpQpvQ/Mz6ibQdqW67mW8a
Lk0U3wGMFlbPBLK4LzVbPOj7r8ao9jySUFiHKgTmGKmOTJSl2Tl9H+ElCJ77
QFugtulRoIW92tTgTnZ+k4bF3gR1KYx+CR6/zU68BcXU8xh9r2HJFWVfDQtC
TXJ5GFVG0zo5QTIWAVK0FKFoAfo8W/KuuRTNcRMV5EBAaOPxthvzNqy2mMX/
g06zGpTvf75FpLB/59B8U1XJvYFjFTIAjssQxao7YTONq91IpGlEhOatsxbS
gfIWkcsuoIDQj7P5qD02RxM7qCTsMnDjjw4MRNcCPFH9AB9htou3GkpFnd5y
AP/Tt5weVac78Y4WLKWRCEIXsNxxAUdV1U+n/rkK6JXEkLwp6m7sSmlUdu8A
O/RxMTUpUGomD58UX//wx/2WzsUivi9ZKvQLHxMC+Eryt/+iauWbq3U3pQmp
NDevZo8MIZMx9hbjuu9cPWvzfZ9ikR9310rOArUYW8LO4FRKVJwo7kuq8pKB
+exBZwpNXv8OLcAneOPkGcldNnXHoCO5qgRL0qft5NQ6akqwEd2ePGZAEog8
DwolVuM2VJU4VI5pqgFEXZKVMGSVyTvE3gVyUJsnzrpifNz2SxOqObHl9Qd3
pPWvxn8yc0Ngfnz/5XNJATB17znWXbAXItgtRH5+vhug78LCYlNoiK6zJJS2
Ws/C4GtuFzh6fqmK++rG8SvPK3AwK9JqJXwoASN6TC97SXye/MqFJxEtVFDv
zM0+/h6AcxZUYB8Jhyiac1D5rbzfcpDicU8FO0vcpFj65y7VktWucbVmuoOx
Tjcxcv4jowX83Xz0/WY3CF5OhXYxLOl0HkZXE8TfOKz1BSM9Qj1GDyXR2FKu
d5McJetf/nf4r4wBecA5OfvT7X93Dznwh+w0pAMXSUxe8/85IS0iRZ3e9Yg+
gHwyuu3ckyUlhbM7G36x4aiaHYyt4+GjVNLwieSaH2+BZPzZeDVoswIW6PyZ
rACPr09X2rlLVk0q1UYT9x7fYVI+P7ohY2xqYfV5111+oaKv7lxBsF7OPB/i
HV8clQyYVXqseGYAV6ambQxSoyBWRNchLPGQ8R6SLNnaq0xc7q78FcXuwgCh
3PCu4ii8FFeVklBhACGBbPrdjQ/VfBKJZ+RGruoltNPPJdoCqaaHWn+wl35G
ZiyIqEIWnaBdFbHTtrhxsVmB9x3EG+E4oCDWZ4FW/OqC5R6PL9/2ZCU6zvLa
OhErMGxk+wWCNETFeVryoIRf3h0BWgyCHG3sf2yQuk5Jg8GRoMFBgZKvSqnG
rGOJ2ufjGWJc1sVI0XaJ4RHQaSE9nBaT9ACLMM/PQFytwJ5otBCCJ0mF73lz
r9WXOyNZyJvg+EFW0Gh3knd5HglzH3yQTKGVlD8WaF3F4WX0txOQATwj2MhM
O0k9tB+bSQbmaH4c5tS1U0Y2sT5VzKLO36/XpwOq21TMiAQ7uGYIfMYnCXQu
qNBhBl7KOvg7NbsMEzCT4ffM4Ak8IU6lhTUP3oBK2akosIRo+3eNSlDnW7Ep
LCh3gKCyScYePe9ox1T0rPaqu8dFonFwrSKddX71k49nY7zy5mXSDt44SEGv
GkL3PmKxqE+Cczf21Q4WgEfA6wt0Mog7NE7mgASMpNGM7GBjfc+s6caSN1Lc
bBvm7srPaXThfZVo/cPr/z+TqgWMs3a4oBEtrMjoqluAD5AfdGRX3TxlnlTB
HC/ChK1OYD1OoLTky1+OPPCQ8+d+Qrsn7sXVnUEbSHkdjxTs+GmfnVLnlV6W
0KPyMjzrneioXeNXMlCLhDnKqJsCU6HsFHCxtrplvyH0oZw+dCe4wndKAW4T
7lbrMahoAJNjM5Jqd80UN9eyYpsa0W7XXVKr1yap7AJGa3KXZDPaYwNiPbKz
StPYECCcTr8vZoxBCY4gVon6o6c7ZwRs4Xm4lAgPXO94H4GoM918uEXvitHs
c4BIGhr60syx2cuA8Mz6nuNFGNbnOe+pO7quP6Htj2MMzznxPs35jzuvtd26
kRW1rIEacr28NgT44M+t8rLZR/YAsJ0BrwlyFAjj6yxv/5VAfchxzBodK3ET
+6O6eKVxUTmF4UqXrocmfoXOQluRG0eoOMbAnIfk17crOuz4jzRSy+ZfH0Uy
odOIAUrJW1dza1HcNrdaqRM5A5mHkP8NSyzs+VgZU40dYXnb6gzQKWnccnoh
FB3LGMuV5JkjcE8n2dZdHDNhwMH+6sTPviQ9flPORyrj/nUU1Pd8oH0PDAg1
4vLd7+PsLOH4cl8/llMk5/ulGjqarnifamcgRj23DeV1G9oDpSYb8gerbtPk
olQiLGrbU22zzpbNzHYDdsO3FgN5KB2bnO07X5SdVNcIMmVuol5t8tWmG3md
IAmIpLFMQJoDkLDxm/afaZi3t0fNdTIrLZPm0Jxdra05yfwitUN2yc3FgpX3
iR6yZ7ScWTFNLPlUtxE9xFaXHYUsKnUxMcvK64HkkF4GeYtCvHpJ4H3cZJGw
BBxVVNOSF59X4vOPMt0dZCj+lH87TatDdigYQVf8eRajNDUw+aJWLRCC0KA9
lLIpyibBzHr8+8UGlQlW+wSfjv1HD12bsSn7TuzKtqEyiTYS2h8fgREZXmvV
XpjVvtnMkJe8DBvZarPxyYa3RxYXklRfL6AOtnvW3V0oj9fTf4WCvNmBYScx
Tccotq12zmHmyb27Wo9dE5FKGIsOGDzWnDyS3b2IO73vCM8b9LGZwL2Yz61N
/DXs7GI5YJS7XiM+F9GlJkYa4QEjlnWXQ0lfv6ksrETAxc5mAemoTJi/c9il
Xip1S0fet4q0ucdDSIK4w7bnUJVpX+vJ54/oPLuxJbBkYvjhBvCZN0a5vauW
s23dPTGSaGsjDDbKvqilveVkGDerqv5y2kuWphhWsAp1FTtsa+y33wm0q2JK
DrwuSyqmbka4VR/5yJoC57F+JY/k6ObZtioKzsuOiaF3lmoxBwVhJy8FE2iR
I1MDIQ6YitIB99RwTgo3IrGL1CxI+/Gqr+P+khssOWIT5kxoLvfLa9FZwESo
eban+r76DKEQ0Jqn0vrMGDl1+XO/mefvNHd0WVfAclKuQ04biGOAL1yLWrPU
RHStozAbBRtSsQDHvLPpT87Ap6wiswJxRRbx66rpZomKvbQ8QQ8MHSp1/dVn
8YiCsJFhlcobwn8zmElEHzFT99Avj8gfkRlC5KtSrXHBXvD4UEVlo3VIol8e
tZEU2Y7n+VBXsHsj9UZb6KG8UwnDOg8lJcjuhRfzr56W4OkVszCk+SYYNJes
mUeWM1k0oF/BLSY9LC7eqJ/E4rcq6ZE0GzeajBzg7MtEeIlTM5hY91SC+jdO
Colu4CjL501GosLg+MpoOZhNjpHklSmRmxwBNOXS7M5lUwG6p/QBc9/LV6vW
M9iMCrBNtiDNmHKzQ2JD+kI++IvQpD8GTx6mi9/g02d7Qvr69ZT3/SriCI7l
cSUlYDM6rCDH0TTnRj2UNGP1A7RDImlmf89n9E2ihGonwJjC4M9GdCVA4uNM
sqDn7atKyfCxBqYwNAG+PyqdfSCE1iEZfW0tOK2UUd6gZ3ZczPC/sWTGnUg0
Gg5hX9oPTM1rXeCdqDKUo1362lRuEDay7EjOVlcz/daX6CByqsGeHZ7UGiur
okrV1/Pbuo9zkrGfos2FiCU72Vm5G9pTh6bTnlgn4NN+uDgG1GVAJkfJoFVQ
lGFNjsnb+RENG3cQZFiejW5vtwwOBbe893YD0cA36IK8D9p9c7hNI0NjdK8A
jMhx6wORp8FqHbnIG80qY8si3ilyJl+4UOYzxZ2oI+cK9xVoIt1d9Q7LesQk
bCtvzwXv6Q/+f32QpZn9Fh1IQ0VNfX1ugaRzCwIqe5zb1uSg6+a8hvdifVeN
uAVllEYTFtxuGDhr0Ss9iO5j5E9jwa3x4ISWlpkG0Bz3hNEbNWhrs8w4+dNc
zf+LAp5PV81q/O3uquqYX7FVRKqXBsy/jmdj2+GTe5EJnvsT1UDY22LJzZyg
4EIrgAFMMKhdmCaojpB181LwLIwx1fxTDVjobz2nAoi2f+uv9TnHgV9JRpSv
PGrKi98DiH0IwzIN93pOqE7rehm8+fDJ3W28KI+8pNKfLxY3bolwWctDenrP
WCoCHGECJNn0jTqABghU6r/E+PVIdFqw6zLr8IYmH8Kdm8+IBmQYXUjA97jV
RS4LgS4nLu4bkWy51LfkFmENWu1kiDislP+QlmYa/faTrj/j8nKHbjS9eQDz
5pu/orabu3z1wIsxlqr1dz7pkQLnS0fDOm0GyF1emZhon3Np3aCrksExCXkr
sfrOLcD5YEiFOrSclVhosKbseQvRIxaSWx+rp30g4HXKJyCRJmOg1KjPVxzd
2yKZUwolBbiVwyoQ4LO6VO+eyRetsfaE133XKD62/ZoM0zQEkcALcnYWLfnY
harL+5TCI2CeLDghFZx12c3GqZ+fedS0wwoLq1AGQOg6tROgrQR+8pYstUkR
8QoYGXg53UGwvmxPhVhYvKV8BjLMbk5zlVhLsQtT3OFAbLf5Pt3QtVZw0MqF
XFTMK9nLg+dHAhuIy6s1isc1gw2N/9vVjH6OJWD3O+TZTE5Zz6tET+PijrnU
zbRN1Y0JJdGw+c3xaj6cSoQlZ0xOmgbB1CKIz2jXYRaGVgBj4Ccb1rhF2d8l
sz+Xt2Hi8SouvGtUF0oOLjsQsok0mzRfwhC77xiGSSSW+2RMvX/FB/whPMvJ
Nh5f/zHkHBwFwfX7NLkTqG/lQwh9zgeZx/g7hPcNd8G3N70lP7bkC/12KL1c
ePqInCgDNIdAT+a5uFUUW46OMXU9E7U8vaZllk0FCupfngBT2+2ycJa+ADNI
NO4Lrg/VT4xejLbM6CpcaI0Vp8nqI4J+KyE7tJd9YhgIOgLmF3c3TlQ4FicV
Td8it8LMGdjE54/WN74yHz/LK1epfJZCATY5RmrzY4u3g0M8mvxEoOmUi/4z
8N1isu6VKdWpCWHsgrQ02gPt+im6m/jQpIr6AgWI0f7F1DgAYa04LBiC67If
VmyC5SY2UPl/pvscFIiOPPUTDxpIfaX0dGYmtzue4c/yRmGnn7Odj2BCOZAH
DNC/jol5EQ1iTOvUAGgXbAscnYKR0gbO7oIuHLuspitBHCnZBKb818H7WDCG
pUfnq5XmO0idmcZYsKLkbNJdlkUU8YiFJCfEu5y5Os5Mc5MyZd4Nr8SJJlTr
22no4uwFRoefeqhHg+Dw4oFhYC/RP/ftWv1tNL4nhGHt74KM+ywH+oxNM9Nk
jK6dKCauXq2kWV2MsmwVywL++JDK5Tz7vjokE0OTPHlFSRkpi4U3KU/CAtyH
sts/9XRGQhAFvohdBHHeN2sdiHXb04SGj8zeAvPnNj91y7oLovDDB1COHmCn
RMsnwiMVxp/jJb4InIb+JLJKCwE+6vx3V/9Q+VWOZqi0EqL4uy1fXFKHsz5o
KwFfwuABaKS6dOGfqOV5hBkl7D961KcmpnASPTSaTPa2HAbfyw7V43H4/WWr
NbGUISvqOmK/0qnoRHRzOHGYA3nBnKLEsHE2IX6UdKfG+BWZ8e50uF9QuUOh
IhK6cggcK0mZeRuq0Gry6XNdNVXB4oLJWX9troFEABQ4LjSK6cfJi84eIHXg
IYVO+sEtDFo8zq2PpH7h4JQfLIq1ATGuVBTORrwV9qsspyvjuDpkPZ4Txec4
8I/wDUVjUZ9GuncqSAKjPeWmbhdVdnJgUbHkFInwF8ph02bD9n8bmTBqyCHV
3bMSLzCYfQtJKUW7z0P/AF/0pYHpSHRroO/VJGd8Hkb4/acMmZ8I2uzt0ekV
BNoY/apYdCdruIvqrkUQfTfYTST2yfQOVheCU0UTfHobA6na+Xx7jJBXhGeg
iJNhRXWC/Tt3eRnYORcdaEMnVUukMMtZGdebsB0Umz0fLOPvE1taprdB4UGp
dRY2ASBtBcIkKH/KyTLH8H750i2NnKg+sT4cEIAvH8iClsOoS6HE72atnT/E
5scGx0rP4FHuIflAm+oSRy9slsQ3Jmth4v+RAzUkrssftt+kPt9SgCSUPlyf
yNq1f0mP3QxY/6jyC8tuOBxLJw0ftNZQlgwtR7AX3ChNiYV8bNfNvTVW8Kn4
VPGr6KNDQ4AKAq2087mOZtxEp95HXZpYcU6Gxw0cqA5WwW6fGJzuo1Roc52O
IwDqo0fhLEGcmII3W435MDp6k878I40HMKyN6qYe7cIJ7EdIvOzBGHgAfhrc
IUmjAwEXT7iLxDwVp4qtTX4Yxaahqun2d/EBTaSYV6IndLaPp2rux+yUln6x
qB2UR1Bn00xjQaptkTARmLXKmLtbBVQrxRey+MT/upSBIe+W0WHbkPEyphR5
g8g0D7h3CoAp1pxLx4zYIzbaDlTdJAgYgWhLMn3v2oSlLn+ijnOUuZb1WiD8
cVW5Gjt/Ya/IlcvHnFIOgTaXmSEUtAQWuOt73I0VFuuluukbzc/TfI15bFs4
F/dnYwMh6hzt3n0MnEWUr1vLimawf+pi9xoseVdDXwJUd020IgcnQk+6OXzw
ZXoRWy8+qEOANTT0eRxTQIU4SnoslB1ZBu3c7ISkWmAb6xs9KhUy47LSFVw0
lx1+uUWUbQjkaIh7mtcJ9G4OKMCGNWB6CYEmHaeLqbVptMpKo/69kq9qLUT2
e7OUcFHyO5rP9k2cdOagWWsbAIeFAJTvnD6esUGqMFMSPgKJKelA6ZCIYPgM
dMqvJUADVfyntbOpYcGwRx+6ljfaUu682+g3Lk6ow24y7UyeVYRGCyvVyJgE
Dd+zLaf37V8iox7skMv97gt1GJOg5a3E54awMcenWAvJrVWSrKQPFykKvF5l
fRVk92cN60Ab300Tm0Cjqzp0EqHnOMRei99RmtWwd0vidwPVp7kgv1YIzDJy
80b8FC+ZxEIzzFnm5jtB7CKSDvl0BGSTXTI+Mzrp6VuKXypHIAAY4GhmuGfR
mzhL9aQCLlzbTai13icsMpIw4A+xtOimrjV6c3gu8Vbb8WQwJd9Lu9m8ZBH8
MgWoWVZ3PB0OeZuCVcFXr2FNYjWHbsIdZiUsalrCjNPAL6KBRTzbMTAY4inL
jn5IWjTfyW1hTyGoasscwtTL/UyhRJEBMxc7zJCcDn698aT19OwEZ5vyJW67
25/TK1UMuY7ZA7oE8Y7Bu6GnbaMgcwIwy4l9dItH2LvnvJHTo6FYG4dAvATM
oWNXQvNu5mVaCy+W6fhzQXBLtCT41jqqKRPlw42HR5vhkkqvcFo4LGgCbd/E
OnQJfKmmQfe0N3erci/YVFqcqZwTv4WAvvDvSWvabDdq9lM86FCRJ13Yv9zg
4qAA+uVHtObqKvm1ETfLTeKSIRZadmBzpdmIqlZkH0GHRa1AG9aU/MLKA45j
JFdyPXyWeU9BLB9cdPDQ42qUWHdMofLy2KlBvPPc0E2g55COOqLYGLZoZxkl
qNVitXIEw1nRnreRybFV2f0/kKonW1zoA61AVEq5dtCsdBU/19+LANlCNU1I
QgyMJJ0Y6qvjbB/sJv/3IotXqmlPaJx3m7RHtLXZrMODkShugATWO+yDOpub
rUbH8PhSCkOUvS6wnqsuEM0915liPvXpffsn3eGXBc970JfwGfuDx1nAlYao
mhbmlaV68XgA2KUGcx7chWybIk4G6EiGx3uBvRFKt39+LKpOPnc/hvEx/BOA
osPgJOG0utVDUlS1M65Oy/4zVNXm+4qVlVQTbDcx7HcjqNmghYQhgdn+LAZ5
xuaKxUuO70wPC25X/fIorKHPMqsV7simWBx8RA9ipVwc0ho+LQcakGy9ucMN
OzdnWiWwzwJDoc1ovnADossEHjUyf2kr8OxwaZ8J3O6Brwawv22fdIRwAbf6
I3aOFL22788oILoeMFN2K3q3RtV+4H5JuYn7iGkpGEGj0zJC/2fsSfyjSIIf
TpPwXZlXO6hsQRtVHNFyuwSRLU2+Wn3/yaVXm/Sqv67hSAz6ifZLRlSyIfSK
VXYlzVm8es5tu+XiVRxRcxtdbEtAG+NJjKPWTutC6TVY9YlizStfN1hO9eBX
NiTrSkjq9n3uG9MkG1E8mcFk677CFcTO/dRMP9FBSLyQxMfSSyAMpSLv+osz
JhrkCRZeK7isZ9UDWpdQpVvIZfvF0VSUzX8s6AVpOilB+UFW4zueFJtD/kEP
PSQJmUPeVwP37h7iZuCH61qVIlzsEXPGy9K9+z/sZUVV9rbtLaoh9+M/WDGx
llS3/JDybJpwqbjhdw3sKh1B1whpXX1LApjU36qcoabFG1tuT8LoCjp6TwFw
9r8uxuAyLsp00pAiUAURIgTETH+uYi0QLtsOQqNO+nYkhAvherj9eYriek8L
ksdbHSgLb55gT4MAI0rtxa7ESYG1c67Q3yDr6VGQNgkSXlVNc/0BFmnvcP/E
wltRAb448RR5y+DQmDhZGaEQbEu3fPydOLWuEg6Hf0GByOQxhvW7HPSRgs7u
6Aj/hHIQa0wlG0jFTmt5W+/Wg2C18t97h2a74yWadqjohDb6PEGoVmpDbEfx
QWJNiK9btU6ZzZlRO8eJPeFW20Eb1E/0JqNWKZaOjHJDHSINN9D8HZd8uZew
BG8HFbkte7mzFP3ZdWH/hWwS6Un0bQbiRHWN05r0jqgPgsP53P0Ui/Ix8WZJ
q8zlKE/1/0hBP1nUh8ZUZ9dcLw4sxmtd6+0FoTJ7/C72fo19Ry6vi1Att413
edBXuhyiOKnth/ID5dzIifax8e0eHKP8f0R94p4Bp+pbGW15m9jVqtNTS/x+
zhOJU45pb/Ci6CrxwwT5o8ATHaL7oOacr4Zdo5tKBCj1Z6b1luaqoTJAga+Z
W2lXGs77dM5nGLGeeJ47xCkZhuMPq8jUTLn8DqP5+QCIIXlRiH3f48C6WoPh
0L7tz+Fmp2Il1yF3ZTxGDSgot9IgJn1GqD5GuWFe0cA5YtPUEo6YMRcY2Kuz
rRbTXDlldjQc5l3uer4542x2hqj//OcLNUs4/vdvPXCb8IGo//QraJu7l53Q
GDA4OKalLvhftPGJx9Ab5pWdVczfwRxAi2dGQtVy0vRg7xwkMa7Sp03UQfDV
XmLJNMNZlngQi83BKjeJzc4uoDxLiqRHvBo2pS29/K1ULDmhOX++4DUfPAga
tPOnaQaB8428PHLzeLJWiJjre/b3gAcNdsVJ4WmkVd1BchnikxfECiQhnhMA
An/gKSKPkdPRqE0Vji56GHmuIzxDcsFCqkkZf6Qy4y5+0ZGlP5GWrSO74/8X
xYWB8iNSJBCUBX+Om2yHn1krMtArTteCvMyfk1apZpzSAeImDFuWEr/NjgFQ
Vy571JNVy6usNcX2Q6FBhXfYH8in76tdkKYyeKbqc3A3Js6hcnNzmLj27b3w
ls89b8hHfvTxFSCt70occQ/u+RhE+Mj74I79zg28XJnupcElPkUtdyp8QooN
sose+GsPRIQYK9/r6L0utOCQrcVDEVvcQ5dViA00Y1G37LTYi+vuRp7eLdja
S4tSFQ0CraeYCY8/tk2uGISbCxUUwvnR0Qkic1EG2l85Kdq6gL5AYIdZdhwE
9afIOBEvABsB0UFxmRIsEQj6+u0uT5UuXf0VHN+N8C6bJp3qPHpC2fvzktYl
/azlj92Ng5tQ8g5vhsvfSdBhNnRrIexocGvLUY3qgJq1lD8zQV+VYHX9Wx2x
BF99sessn1jPhRMsdiK7r5TpJL/BS2Miei628pYahLHDienEC6A5i5h/FvvP
x2bEcHNXSFDc4tycAs3HcjxuhWe7g6j58CReAH0k4AVqa1QOEbP49e9RbLqe
GoCgW0tXg2hsJIVqJxIG10A8+YiimkXNR5a9g29KgzKrEqTYuAACj9FjqrFa
d3e094NKuab89f9FRtpt3A6c1oH3+wl0mQ4rK27iUp4n7x8dO81Q1msEj8uW
zYAWKhzXuHLh2iG2EAJWG5K/KfX51klPQTjbXKlbe5PHQYqD6TEBrKtJ0b/b
djWNXYi2jGFZ9gRN7LadRshnBLMYY6bGlzqOMffLxOLCNQQbb6V1ZmzaxVtp
ETMm0Y6IQET+h3yxGdHYMax09QShhthHyX4r91xV42QigWHQgKkf/FbpYsg+
q4GiZAvndZxzJB7rv8J+iWgsVnCU38CaTNnO5FEUV7oFvbSFm9Acn97D7NJv
o2fcZ4Roo07Wf3372glA/sMpnXa0b8en6GE/ZoQjvMNbivl1MzKwx1QKWECI
5pTLDRMkSu884iMBAwKLNx2OLBxLyTKOA0eYHVVkXN7UfCCvn18f0X62TH0z
1hDSggR9uOdlLt+4gIf0/Dnp20byYcEX9ilGLfXj0FkUtFnOdQVY3HPEhLWD
k9MczVjnOHr5usjQl9ZTvlW32zvqpBkw9bR/E0q8w/HRYsZ9BBtwsR2/jGCn
pho8lYLgR2Meo8721YpDwfgAvHuJenhX9IFLTBk/cFGcZ46Dft7ylztyvfKc
+/g9/cB/CHEahBITSWxX/t+LTcYOuPI3c6Da0tFhYKMVxdTBkoinlWRGKCRb
A2azhPBxHGJZxcXvQ9VsLHHe0kGAlP8KyziJ80Dwzp1QZUewXEekEOwfyq85
Nvu1j1NkNNru3RG/wEma3VmFY/5kRCihRMSckRdp/uTiOGXxzzAfebJO0rW4
+VGMhYjq+7WUHA4K8atAZ/cWILN7CIZGAhYjk8fy/0ysbDF253BU0J9l2FwF
djOvivAx54NvqvNRMlvmlAnzs6P4KXYpOSFvwH9T8qORFF9R6/V0CFEWT+g8
v8g2aOQu3DSBp+jY4iuegVQDCMCG/2VLzePAX3vJqZ1Rcf5+8Rwfc3etsWMM
1JCV/wFPpGB0OiuIjBJ2lruNtOezmMjrUaM4tuGrxBkvonOKWDjwRdKwfWiW
ZW87Vb8AZH5IPVP+a0Pj0uaU//koBR6EDGb9xTZ+Mr0593AT4iG+8wffbb8y
dZVoIylMOXPrQc82lhGYSml6PLTCOcWHiDdkj5OLA1nJd3R7QNR/7NTkifob
wxdFpILOrhFpl9qrHGq+WwZq1h4mSIfnzwW/ASli6UrSW4jn0JEurtPR596F
aEmOEyTcfdmi6h9myzoKOUjclidRn8qYiRarUYfNBWg9rdjHkC3zvf0xQ14O
8OcwM/ofllNwkylmq7Wb7t8PNjYY1ITqJQXYm8fTKph1m6xJ0c7WqSMpRH+C
MgoOZus5EC22SvVh62Nyl0e6LH1TXc3OD79/bv1J5JaH1+Gmus5S/kYASFFA
UCsgUc1otsd0VBtEkty5mBxSgCztS+tHwpO4Hzps4f06MwkfR6Vg/izzJ2EB
LEiM0sb+uJlTb3F8U09rrb6JfI0cbYBp1kCf/2uCqxxeHrAa1nIkNdy1JGgV
MoWO+QWafcZbQR3p1NR74vb/q4WIELqokLCDcPg+pdEWcjISLgdkWYHd4/7S
a6CpFV2ql4IjMRW9O5KiyJRBebl2+0UjwQPXKUyROy54qOI7LuHeebSKF6of
NxjLtmbnbaVk8vEGYX4oDyaKwOskh8ibfdyRDOcJBrI6q0Yc+3mUZbHLN9e4
YNahp7dcm9HAO5PTFVqE0vdsDNbwhJ+O7RFurRRdmpp/xg/RqRcU2oKt65A6
t1nuP6YvSsPgYsbI+Ve4hYCis2tyuYuDF+ZkGI6UOC8CB7tno0v63n3YnscD
wj/O1O3x9V/NxjQ4sJWp0KNha3RVr9h0MezBQ1hbTNwoexRNGhMoEjLQYh6I
uKseitov1kJ1A8BrEOONS/FhOJdLswruylDbvZT8BiDnTcqQfNMfcWmYho1g
XC1z2JhAQp5WjJnFeKVtI9q2X/Us1bEqgfWRoJox/ZVrMbG73g/iME2vPr/z
0EPC3XTyZ7opa+vV0zzFYmfe/t44Uae4DWj6lBmAom11PhfbQmYQh8Qniere
zJz7dDMhW3MGT8jGQyqtF1k5jNGaQOxahgXyEdPMwzGg0n/dLDjys15h93od
TXxUdrCDD6b9xuH/sapMn3WKAu2XGziUk7kqwTTN5LwBcYKKQQVhNqQyTk6A
rd+WNJ3IaEOgrj69xU1D4nO9kFH8rSCxw3ApjZZ2vWTDSQFSHKQIKlVNI82r
AH3flIKxFfJ4/GtlyU54Int9u5BA/rXgLShoUJrMFuMxEI9mnDhPSJ/764m5
56Cu7aJDLoyeDgqKrwB8Z5edafVMQgQat+Ucn/QnzkW+9yIG15ZNLAZhsDFy
4XKOZR34PrqMLuLVox6l8EZGGSMX3qYbnjHxT/1lWrVVi5By8UgbpUih9Jgf
XxjC6PeV0xxRzs1vnsnoLE2JTizJrdXcrKcskmsJMK8bzOMNL/8S5GVJ423z
QsUQ7GlObPFPIfPhfkG0WuDr4JB2zO5ATPkonMKFrG6srbqbMeQK2jsTYZqQ
DcshIQ6JErAMknXRTuNpU38hmccqIYwoGcbYZXb9vvm9XILLvoMzL9kH0MP4
+gFcQ5WLVJu+HpGKrElxhctyBNdSMUtfFoXW3jyb9CK+qWiNpAG9vmk7jVnN
SZZntButmSqxR3PJmHvOlsvthN2DPb5Vx1L/NOr2mdFR6cAO2r9M3SKEj+3k
1c+FBt4GhIzzivyNvvucfx1KC8WvO0s92n9lIg7LRDxEWUvK+VUhSN1zuTDz
BEkcYWVZ6gWN1uOs8TI7hX0oKcLa75ThM1b9WdR3vTuYO47ULumsh+JE/1GP
JA4+YNaEsc8YnzbhWuhb20U9e+qqA3dtF+Cbx7nGzQDJ/eTll0YP8etADr7J
VE5wpL4VXS55emHMGaJoihgXkrv4mQ6D1/bvv5L/3UI32CLaKHFMaYiMQSmD
jmikU/HWo7JfF4t52uS7hWqkPRS2PfQyEYOdjYikJdKP0P1dLk0PwDj9lfVQ
CCc4htuAZoj1XO8CZ13qIRcuf1RZ7/oBd4HDv2bgJyLaC+2jtzzN3PlCeN7t
iBlHxfrWgYrOaKY/ffa9N3TBiv4pAEIbBnhPCkS8DfpUuTTvaadILrxm4nwP
w4tgin+XCO0tIR/zhrBeTvPqaXyhdh2ePLdFQAIKOu6lpUBCkRMFRak0Gyuf
3GLUPXs4FhAtj9AWNzdLHr4ah1L6UK+wfZg2nVfzceXY+UshjOvg8AyxHNkD
LoQUlHxDkDuvQ2uP2DkVK4RTlEaIT4lXWgPTjTXAz2073WlKHeICraudLo2C
fyWUfGip/yCDYhCv1xvupWE4o7KEKtIA7tf1Jf/ueQEXtVeJDKV7QCrGM21Q
d+YQnnCcoOuLqvy8PmBE5q8AJTO2HJMS3ABwm9QpAhe34IMK0nSQHLN4/K6a
XsSUM6q19bOCZJLtRbTpQLi60RUqE4O0iXD398gu8TNQiJZ88Hj7DCsYA7ce
ftIpOBhTwu7upYT3+EYzsYyy8kpkjf6MbD6xHiDtS44FkhDMK3jiFKdHoWM0
zfu0WpKBOwtgteqGuNFNtG+h0LDDwRkVggCHT7Mzq2tRkI/HyL8vh6xbW8Vb
qOD5ORFv6lpIkPdxKXKuoiO60eXBM9Tk9WUY4m6iv/ZZVKQpNMqCFPSv6T8u
coFNnqaKBmCklgjGyAnOD96bbYPs3ND4TKkYGQ4kmPhGuEiTzFcQADU/p2iC
7jmBtb3jzQW11a81bhS+8LuAMA6QJ+0WJxSHBFu5DtP0YRIEyXq2YVuHb4I4
VdLoRqjOTw0zrsDINKcxU8Mc0zwv4ow2eN9JwC7rKuRNPzavHJYZxjOTfC+S
jOCFfUeQPaYE5sQpwJZEdDusZahx/fZXsrwZmUCgiNQ8VSztbfN5LEWhBzB9
I/NYaj/iKMlnV4DAgJ+Jih65efJ3+2q93MLaX1UxFQFn5P+OEWR5ZjCr2aGK
QcZ4v4Pz4MSq4ksuUGkUG5vEoLbumPwr8P0qcHkwKvpk/n3cSraaHec4FlNU
V1tdun2ge6aT03l6rsglfvnwLJZR93NIrDNLiPhcMXSNjcAYIDRkcEJfz4VV
F1Ib2cOIIpGU+nRqIIjKjHZMKRgHu/fvICp3Al6YpuEIKpoSYhJL7b2f55Yz
wLirmumesASNocvBje18U4bRu8UYGCwBFdYxV2sGVVuFttLJmWzZG6TYWjCg
4n4pPMuHvBJJkiK4GZvSyd2U8y0WlfnMw78s6xwfBoTsfAAIYQh3pDUeHWWd
Nd32YbyW5aUW27oS3u41i9G1Ag9pbYCwgEGHmUkvkSSM2m6R4Y/o1QnAvu4s
fLIG2CeWtKIg5ZmlW03AN4ur2lsLE9g7ccdvWtYjd5dT5YxPGnvKS/7cvzTH
+yVROCXu7uvTns13iSC6Cb1kl3oSpfWBaNhP2UMRZRKuPagay+7tFEgHZGB2
aDNDT/LAo77Cg0BYOtjv2+u/cLJL8GgDtJovL17MrNIYhLiDqdmrf1xauqJI
p/1749HhSMhu7hExjlDerqoLrwAAhEtqqoaYNirsx04WX28o2Zxm5sw6Wxyt
rw24zTw3YOzUYAA8YHVxKUQoLPWd8NnsnDsMPPvNy7EqzKPRIea6bCJ+8KTZ
c2x9vi+TKXmc5BErESw2MK5J5ZL6XhZegv29xMUIrCyF5xM9BY2KQfAb+t4/
ElmYlfHGJ5DV9YjDWamo2kKo6xw26z5HnG4cL8L2Z38afpvEr/eKEWddh/Rz
/F99p/yZ6dd3+8Iy1Wj0Fv36YfGA++Au8DcjKCBs2gi0rBDpy/4+esW+Em2I
BV+YR7GZHzn6Bk3BJ4NHQ0lPA+aEJUoQuihT2eqQ+h5kRVbhJ/3z9jKpT+Wq
qelyWJQFr/zgLREJ1EYvLtez745e34WOmtCSmjTqGE7PpMx+1iMnqsiqhw2A
4hX3+GaSGTqccwRTTAl8NymDbUM9r99xflEW6n3aG631d73LNz9p9nv4Ta0D
W1pNkpi+251KFukw8l4vmmowK3zg/+0rRnysv7sylosczsx5foyqutn9+pa/
8Hck41bcZAozWPfPYjYwQDYPLfS/uu8UQaIwqpHF/sjxbpiPY48ofZZyQjqi
FBNX87qad9yS3Yxfb9AtkRdBSQp4MmiEekQjz+s+kj6KuMaSa8cnNsx/PVb1
25AiFnvCDGeSplzgHDgNSIFD+dG6PT2hwBQ8qUpRPCTcyRAnGLDRzek5s80d
e85olwFwn86VCS7JL206upbJ/cky/ns90oVtXJWzF0zbpb2T/b3XRhVkEknX
BpKzslO42WM2psIFS2cOR60avYEUbAiby5NqvvDdEpGprYTlSzpQ1jVs+SYr
yce4nAjYn9YfqesqNna4GBjrB8TisX3eQfS3CtAtWGPXr39BH0YGGFk2DpTp
YBNL0xnfH8EB/gsh9AhIBG4zgOY7K+QoSu2o73dT9gH/zHKSCgXNqV7DgU1I
5qSKddaw49u5Z+WyooMzzAIYU6San+VBQtlSjuidpbwhBFXFz+rngtatyi7m
3gZOqMVJu5Vw2M2l3vj/C5VIUmX1Rjs+G42JnxpR0R+3/BRZ27Ysx5uUYAXC
tdPgz4+7r+RGD8yy4eUoofXA8hEeOEprobNuThOr7oSeoipUtFr2u51OWIm4
0HYEPDR3frDUJ5vI+OUx6vPn98WuU4FiSiIup9hsdqfPzGtLevlQQ+Qygd61
R0gIUJFdzo16Dp4m+i0cFrWRLhxlISllyeAh9LSMaaufYuuxIvJ7+YC9SWqm
EI3EV/r8NO91V3MjKvDYrUKY1VSRF2nQuzJipKhtG6jISlBhoGz+DviXo8+q
GKn+Nis/9prJIjMbeHJbVQjhzwXhMqCPj1PNQsdYyEd9Ov93PR249AWfaQlq
V+H69kO6vgq2fEiJ532w41ZLlDZzDhdJS4HxMtZEWyU80+dwiAy8vIZhIqkr
V6qkmLP/O6ryVxCLr2rB5CSbiWy22I7BMF8eEolHJe83tpmhRd+RX7YEBG+/
kCRx51vbhSJgngUw8Ou5+XyOKUKkhm2bCNEmlVkKt+rqoBmjf+hxjZS69SKQ
zxqnPAGf/vmihYPh4BHS3WpJ5VhEFVxVJbo1C6LetTU+QTsCaaiImqD/d9rA
pGoK3SYM3y2VecuIjx/GLAmCwVSHfx17WLF+R1Wl28qjrt6Bfc5/aLh4hg5Z
2r9cPo946Jzqr7dVUwHeDW7GEs20oTnhnNVd9n/sIGURNlGhVXJkzyvbJ4X0
OLFvmzl20xC1vPuMLMs2rx/G0bggS9xIV/yVzjCZi2NIVMhN9+G4BQRhheN6
9jq4/UxRcRKPT4q8qo+sbTdFYFUgXpcMUIb+Dmaw7C0P4dM95zopYD47sjVq
POl/z3wGhBEjhwJC96VvNUR+MX5Idkfib9yStrFLeJd4wtsb4el56NN4Pcwf
B8503BObrMMZeb0eokp/mWp/xKWfCfFOotDXxyqOAyxzJzfbElCPKHi2Nolx
J53Mkhxh1iCu71QT8nyr5EZty20w1du7WYhfD+PVP7FJOr7Op95HHphED7rX
OHX8OQArf6sQ48kuWbzVcvnxmbJ07Kl5qfixVgF5L35dR5gTSMVq09cQLj7c
tXrHR2aEQhrPQfL2SDqYrOIGtxB2xPTU9N/wgKWUJHHSSCV4tAGvy1C6xaO1
/ixNGt2NOwoaNXPjEmUdOFalCMLNR8Gh6B9cuaNlV7XK3LCOfPwY1U9g8rTL
H1hJNwSxQfXdX9jZDtc7Dp3wv3DW/CPbG0TuBDRlea4VxgmlCYb/Ulz4J4l8
vRjTKWzF6/Xld3k2x+genK7gi4KfhpZY/3RHb0qvj61O2MQjo1RsXHj28ESy
7kYhGkZ9qFwjCBp1TFo+l1SVQSzb1fGO06/6GtYUwLjnWt3+a06hDl2HtOZC
34wFt0ZkMEBF8NTcppeiodMJ44EPjlF6xZRosTImeEYdI9eLB1kbj1lTnSE7
fHvPtVrd2WXfwvskUE1yRca8mKRok2PlQlrtIy+d0ITrED+JwTwT3krQv29d
DFhQsVSFJ+0ya9AJU79iQDbuTgaLj3kQzqF9kCBwFO95iKiRR9gGA4hRkzl/
TLkhfT3fmmmLEImP3hHgpuz8yvbAziJkfHWMn30g1dTyGFaI0QPbx1J958iT
8Jm/IemxmSgtF56rqK4P9i2ua35CohHhOY0142mmT1qasZgVuSZXEe7ZUlbO
bVLIL9ZQPqkPvQi24zgd+mwiEnFj35JsS5DS+/JikL7AGepu5MdD43oi1ajN
U3M5rDKgdTJ4nOrWTtNpN/xchK7f8E2DVr3pyJ2N6+vdbm007TCpFdofSikm
EOPWDpsYuoiXRjosGvSG0DsleKU4Ek5GsDGAA4qWPHZBDpVrRnYsMemNFRO7
kakVM1tmLOTBzenwMkA4e5DtV6bvhviLruPENECEqO0tlJ4pkHqhl+EZWv7r
BlvMdbox1dNHie0iqlDdDJCCHng9MarH13o48SsXkdGKBwTBmS1d/rkgH+e4
eOFCrfgwAh4hTrekW1/gegMinv7M6IuPwiVFOFKNF9taaGOk9QjcrD07CBFr
JTW8wn4fRKRCRKKlWXOfF7FdTJ/FcdnM01ywnPDxczDd5nvvFXb0Xe1tAElx
5MC9ktyOIschcQ8kGSnHfsX/8wCDhaBsZCSPOl/WAWiko111RgByFtoonUv9
5/26W4k+fzr8h9K3l3jP0W0Unkcerj2JIHtZ8lbRiFMuNyaLMPkK3ALtApq0
MmQ6ismWDji/6Qrambv/Co5+OtQkX6L9GTFtkn7RwhVxqo35PqcWcVgcpE2x
3eowla1ZpFdJxbRysxEk/Ku4YNBuDV7AxZ6CCQh1YNHtqipmiUlsk93U58QC
PURCttsNl6d49tM0Hp0j7qRQmes6abEmpmzSGNTX3qr4tjaoAac7ur4Y9GFL
b2HUimWxE2hLQGahI2AjJ8M0gyH35uKCIfskllxOL66l8ketqF0TOdnUKDkH
4ZaIecZOF6EalD/lF0k9ZJ1y/dq/2h/wa7JtohKB23TsRf7+iu04Z+ovIR2z
zgiuCEB0wxwBj0M3hQNGfu5jhomt/RGSL7DkefXt7GA9FCPXrg/K03sC7ffB
Vc6ZcMj3VK8TR7HXGnccO9DByormtEKCRpco+0yWWQy2BtL1ro8QXqp2s8E4
acHsVnXtqomwPbBbGjmop1TNjnLBF0ew50NFWDM634OeygEJ/zjMwSqH4WG2
Q/UmGEwOLfQewv4pqUSsIoGyUyHSH/OjdZh3uzsoNGR4h37A5p5xlvSqcfuk
t6KWBXkv3j+TiaHR6Sfhs0qjzKMEYe2d2LiA0OU1w+pcpKDx1A9RpclxlkWM
Lz6oRlgT/CUn7eGIrPQhltGcfAuLnxezgAM5qDFubEqBQzlI/ZVBTxU56VaZ
4VzlmlejIIBqCuuOAhaTu4ONjwyYDp/9MIuoSWlLdkcI9D+AOdoB61KRDbyj
v6XxwxGLTfHEhu7Wn12V454Q2WEPXwaAJnI4rFcPmUKXGvwBGt7ugE0DxoZX
JpwBCwEkVF0+a2sJF21SSqNmLNHKk9+OHJVaC+DiajQqsTMWbg3I+qj60SkO
tYHocT0dW/a9rq6bXGBnbCZYLvTrkqzZo3y1G6rG+yFp0Kh1XYef2BvORA9H
hgbu+CC+fG5QDl4GsLfObqzEUKaGgL+moZRZsS/06tbM9Xl1Ph/fifemFbe+
9HA/AMHGT4qnxieBzxfiypWdg5oE/XuLgX5EXibir3oeH+/W2BB9FIES6bWv
JLgLqWbeIQqWXgY0Ixev1jVCwOx5ARm7kym+2S/KotxeBjPovbU/30GBAF5B
DIBJlQVgxJdGot4c+OaG8TP9JPlgJiZVqqobQCIBflhEKnQYDF2iDsetDWSD
rVsnW/GqkE32IqbQR9zsC1nwwdnL4gx3a8tAsm68sjhaEWZf7m6HmVAK7HQz
b/oDqYAhKiMEAMZIGyfmPQuszZBFUas5mSXh37ow/5bI88bjn/gAlygKVpAR
Q5EhqcqNepNF+2BK3t44fwo8FP3SpHo471plpg/Xu+eq2sVDQ8Z7P3U/+iM+
mu1ffwIQ0/VrKOTgFCloPWlvrEkoMxSjeuVDjRgnLyUKPG2FU9LChQqict1n
YNiZBfQuLa1sZ1YCrxyWT2QHWB26eVKszt2wBUrtRHoSM2/U3+vKoRUqC2P7
2UrpDWXzdEwtdajInhjp9xjMXj6JvLclWTjmykVcdN/XYV6s6f5WPNUrfvJd
88TgM6hhoOJeL/WXTFB4nz1kps9zIcL+01tkg0v2RzUeJu9NaZJD+0ulA9P8
9GrFQoLa8qinwPyxNLT4Y7S8PyhiQAqS4v4NCKJQxzFmdKcRp7acP6sHkxpp
0y4kusJd/Nkk7aIxgQRHJ+Sdb9TumxoM+yfsKdbCu9DosnkX5bM75vwLWgYF
dvPTXkO13mLBTtsR9B10cU22B00NZeHSvdQ4MK51k0M1Zpm6+8v389vI6W4t
sQADCg3BkL8ADYb0v+MJBdLTFZr0nmvO/fBfXkn3RVdvrAHSbGe6ftaKPXmU
kicnOKpQrlIMOa2CoGjyNQ9nDZmc7YVZL5jQIn1VIe7YX7hKADlzshmQbUfK
9x3r0p6mxZefBYXLAf7GDNd1RNuMoHyA8eYRxPg+jc8fi7dB5Jr+3C71tq8Q
Y6NbEYI/0FLPNUNAh2QS5f7ijy+ci8/Yq1V7FFD0Jnh+e0jSCJ0QRBR5kIt0
11AwR6+51BU924oVubUoB3aEn4srWNi3CgchG6vHSkqdnMOpVARbq9nwdrVq
7LujtUrE0aUXpngr4dVtQeLSjE7eu0OiGl4VWclIyl45l1XoS92xTrft1aJY
xorFpAO5J296uyRFobL0sbZt/RWwhFQu8+4vxbKjERCUyX35pWwi819e1dmu
3BfGWirBBjxfD4BFhq9InK7C4F7fDg2JizS9hmZqzqZRcHcoA8tJVpvQwtfr
ObqXxzlQdEgTKuS1jwwbmOQSeJigeB/fDtU3pcUqfn05gK0SuBp3Vym+GPCv
8hF4/5FRixVK2Z3uFm+IZEKRwxPkGx6HnXpdSwS8SuGj7j+OpqXIjh78mTtY
/g3hUh64qE2ZIuKJkcq196PJbUN0NuuE2zmYB5sovxhQ2jv9bUb4c7kdG2+H
icCl3WoEkIQ3BHwQ8Y+Xq3n3XaxDfnilOTco0PGqUAcF/DkPHimdwpiamwPa
ECMRc8FnRS/bvhOmRlbfV4LBjrfkuKh9dHsZUgZQsU0dGOJ048Hd26Mj55h0
Nn1zHFb+nv1uCwiCxruz9eaAlOGAvF79tOhZotnuyXrJJoaqZ2wiutBXKe5W
gxaJCdaC4Z6cIEyTO/q4TtfKBwz0Su90cDy03MZcDri2T5y+BuVnglSc0h4G
WIUCTzRE64NXTekYz/6NHxNph2GtHbP56s2LbsD7KL4K0zFtZplxjmc/YO3J
AeDrhxlMg/ZCdfdM13IRI8GGrIH2xBGEy1h+LcMf/tT3sRLKsxotddE3IZoJ
Eocc7cEjzzLcJFj90h7p9IsHfFEYYnqCAgy9+EnhEHMvS4nsRHQE4bq/SgAA
OvrsNRpn6tnnVN+8S6A9se0KuXa0oDzsKXQ+p6ZFyLYn16QOXZfiWhp4Dc52
DmIzCo8S56dpxZCniZBoAJ15z6YAgJKmQnO8CMZEswoLhha1LeDd4KE3UPxB
jSqjp2T9iAN0rdV0uutNjzYcSq8DzbAMLf3t0LAjGr5Ug0P/wIADn+6DLaI8
SjWSJrOyWaoASn24OWSmcFsz+NLd5al2trxJyZ2EwHVxK9qhXChvE5NnPnjl
miPHNmm4up3BBERIn4Rda1eXuoc9gxI1WM2X4Owwp3nOXOgFDIEhKXGvdHc1
1SfuRpqawz5lQl43iPZImFQiPLoivIapcZzzN4OUqOyYnrgbC9X8qN2wD++Q
zBOG2XaGaueAJ6LscFOergTYbGFWJgbC8lEFTA/78LaBt4OleLNLDs5Y4H5G
ilFKN2nbb2kNvMpCHXVuJSX5xqdIi7yhlRHxnCNfh6emShBZgL4KazPHdQmu
TyKffdmmE1mxX5fcGmLCBg+4rJQn+6q+bGxC0U9lAqi3e5378f7sgFO+IRTJ
ArIPXR9iv4YPJ13sA4BWec5xPlQtaDXrVfMKoZZ4bonNwMfMgbJk3MrJwWph
M7c+F5aHiYF7UiO2hPoAuoPNkTbrQBKWW7SuaFbj2kwGLjNxqB8ECHwQ2I8v
893JhaWweIdmDVwnJa+W8o3YLXKVscSM4W+zS+Tm+dmMdbMckRgmY1219LiM
NSKgLP++mDfCcDkWwvwlic2LL72h4kRXobHEkTACd3JQPw7VG7WbZo/SnT+v
tNeVL8101bpnTMfZJibNYiWD2b3ZViORqvdfvkvzEncYS2CeFUFp8oU7fVqL
cMd4oGBg21/8U2iHWyon6sYYfpGt+KNowhFkTSBjUDO0mvqlvoUVqLJtxn6q
y/uUEmoQpCQ1kULS5ukXc05zfF2KegTf4MhL/C3xGuk20EPPG2dLCoYzm0G4
qANc/+t8bj9J0y4Wu/IQDUwG0fkIRqmqYubGpuB7irUVZR2f69aSCWgmJFUx
tOaOiaA1PE4lLz/M2MjE1fmYi/aEVc5x1UjdxL15uC6cUa/LRQ28NjwbxYpW
9HN1ZrzPYQIQr6q9mUskRtkhtWgUQLd2q/lrIL9CDnWroppDi9o91rErAQMY
5bFFEW4co3zLAWeqP/thmkVfhaiiQVED5g4/Hj1+dB4JQ7a2bE03IUe0cK7m
CMeMwj+wXB5xvkkFayyYSbQij+3vzkNK6mwuX9GWTY5/e44OCz6i+AmCa4Te
0rfq4I+uosli5biKYU68D/KgsOYm48yZxgwltpWsE3Bj54cNNtUs7lnEK8RG
eFPNKcibYUNFJ0WQz4yBVprSjIDLGT7VH6bzAJJ9YxUxoI9aZmohWSuJ3J4a
K+tEL7DK36H0ZtMcf24suYuGEoTw6PTDOYk68qvlAJazSLncxW8E2QvFXlxs
vqhzKsG79pwtRB3yD1BkUrJNYLR52Cxjv9EcKRQr7WJfR6YzLPy/sQP1Nwrb
NWZzH+D9eQyNaYQRXq4F+SOuPHIf21tOQN0sY2ulwP/WEupkccu29zupR0KF
SM1FYaVJfuQHgzkpKBI4ofPcfdlHSkG2DQiq5xCNwUaYGhsFnBQ2Qg4D1faM
zvHGif3mEhaf/5OH/YT1+1VTZdF/j19+oPB5uhxZFNfO2yAMrLXlsub/TALA
nigeKE2l04RH3fR3wvMcr7aJYhrznZjMuHFC+Hrfreq0qqear1SypR83/DAe
qrUJRslhJsvE+AHADhdEl3E+u/9kr0G14pJ3vJ3nNMYGwXogmDxfx/jJIaQY
MeyFoJPxra6oUzDXh16aO1eZvwVKelUnKJNePrJY3ZZEJb/3DgMhf5Buryba
Mh8MiFOhHeriLO6ikbWbcn92zyOFs4usdr0zYHpN5JkQI0X9bjj6clXXK6TU
BUyvs78HE62+Z8OVIb6jO+veSYGZ2tJwAKR42GfL6N6t1lJOuWw32S/z6Iw1
ekVnOa9M4uaDaZPZWHGi5GCx9+UEbmRFq7dUa8o8KJUNmKTL4XUDJlefR8+w
IJWUHMQ9RD2RJ67DIe9t+G+pupFllYVOsiB4PuGSVNaGQaqkAL8Km70QHGfK
JB5WgYyCCluEwbVKX4sZMkARLtyVcLTSPfcGfe95Kzd++w9qSJ7Dg8T3QwZt
2S9IL+PwPo45VrRJaQIdEcZ+h/zglfHDzBk57wLnWciptt7a05uLGnb+vN4I
/HWa3I/eeLMEtk9Ceh3TYpzNmWQ0Pa0UODqDARaxAG0sUPNDvw0aliAPG4oQ
FwuC57ibB/AIxUmIj2ms5S9pQi5+l4Wr8GojPQ+ZNNT20PriFa71OBqybMh0
ky3Ys82co8Q7/IwSbkRQFmNaDz+MnTFgndNN8oBzxoFUWrCrtxb6P+x8If39
uNggRVzER6li+U+2hjjUNUj7GBF++BfWRT69CQhNQo9iJcdnKujzu96IyUr1
blTTAhK5TbsL9Dz9tgJ5YfT+Yg/+dSaGwVE4E4ZZdD9hWtg9Dc2JOTKxS7tg
5uO9V7K/iMzz3GN/UUQwZBLVuHw1Rk0G3G7A7A4wVVdsrVLxLIQZ8lvOtfMY
v3GIqbtHwiUD9hIfAaYPiewgq273uiM4ofSaaHy+zWb2egFNn7KIDFIehyTk
59wzJHJDiwhcsSOOZ/IMeCl4IeOVUAbmJ1d0QUyVfczufPIv6U6hu2O2y5hF
ldu9x3HAYD7suXQ1g9QK68ya5P33WssOAIT+/amdygM14cMyZdcBGAPuZErj
OVLQMr0k0YvqHj6q38Ng77EHNxfTRY1/YNbd9DMtVk1E+F1vDboIo4iOHQIU
D2k98ycykqCAVBIuJ6pTGvs7R0g/jQSsBb9MFM88X4X0X0asyHegWjW+Vn2z
DwFXgc+GLlyWs+X7rgQoX80CLMBvoXWJLdRAloF48B/YhooMlVAdmIaHzcR+
5glCezT+2a5hJd32ba4+gsrYamQANy3EDxX+gheiyPkLd/SV6iOtuhY/b/b6
I8mnFErVhE8AAJwX9wQxX5LGrDvnlFk2JlIfgFzKlsiUXud70bVR9o14w1uT
7dMlUYppoipNQpd8G0crEDRNM+sXW5/Xj1pBrMf6ZOxs0+TQUH1oQi9BBzbq
PDTKr/meZgUFp46A4lWQmFTd3I9hmSdeiLxRtx39tR1JhGdGhcnGBy0NR6z/
wx8FRpaudPpGJpaCI7+BDdmEZNTbMjdJOqm/3yqEURs9QYJ90O7KOGn6Z9vl
E6ngV/AqlaIr4bdvIf6Sq4miTqBj/S6AnniCkfiAn+F9kaQ+kMdxMGixlDhj
iGLiwLPV21GjEhMVoPsO+LRT00roEbXL45XNTkPbpU537gjEX52qndUqvn6B
2Fmc++RZf5lwzP0CV2ryFjjD8BYvqz8PjxRzJdfumYMIH8gUJYVuMpMo/dVP
2Ej4PC+TQweSkXMxBubetqfn0Xm0Kj2DpKYOfVksUaUQZYp0qCt4fWy8f6Ch
45H6cFrDA33hXtX1ADTPU6NpCXYHG2N/8GVh1W8bs4qgSo4zyrpVroirv/JV
qXCosIog/iNWdrqi+G9qrOZRnFCaKymwxZ5tzfpwSFsUjnlMRUxZJhf3Rl2r
Rr7GhUCsv741qTHHrRcujPfsHP2s6lUhXiXpJYTFTFRGPSOg9tX6KI7Gymgr
AUksfR8PUUV+114m5nXbOliAx1XVte/7+wIOZ8krR54S6LW769rEj/8pI1iZ
N2ASQsavGlHjrqiuF50Sb3kHBK9JSWy2dM3Vnttyai/N2lQA2/60X2bCow5r
cuED/FpOVulIRL8MbamyJpxRchpz8ylTCpe908JcOP6JsG/slInUwWHanIme
+AvR+ep7EnTS1CkTx7YuskeCKbxkpJHY/fzjWK+Sr1jmoXFjTiVh2YNVmMfg
Rrwyea+lJf/QMYA0VmZ/1XOAKWrRBlDyamgGQVCMqw+6Ddv20MNgQx9TNkhp
BDrsJHNg4kfLyN2BIN/h6aJjMEaitB7XGEPKkgW4yn4mrQ3ew0PZXiTtx3Rt
dj+BfKtX2YvocGoyqcGZfwz5PKnS0WZc7XYrLBzBPgXYvOcOvA3ygOQn3v+B
YBtjJuyx7xypZT6vXE170DQ0IibTLEBA1go1LSOzRzs7znfEgLLX7A2gdKHF
dEvPrArYN02SiRQmV4bJWn9mcNqdrjioKbc37IkJNsbaD3wdBtV1/hHYQnvp
HvZy3MAeMsnT9Rvnd/AA5Ic/V6VmiE6FHC2SFI8dTFnnziSe/pWZWRBJPTlz
5orNhPB/AJtk4JsRDKWmVXX/qa9qm3Njm9+hPghpJc26XTgPXddo+RDQJXBA
Fo6OJm0Cf5q3Emm02QuTOLtB4TREGeMB/oY7oGLzQDyKLQWWtwQ4x9GrX/VL
AEOLX9Tb+TiHe8N7wKEBWwGfgwn61e1RAcTb321hQ85E2a1oJEXJp9VjhFjT
wKu68M8TdOo/hXFgMcfn4/hZ9LylN8umg5Drf1fXhvoPz04YEY2aolRVEpJZ
+EEnUzVEm9cKTlZbJnABU0lbkXGxVouM6LB39apnnc8Ubfz9zmrvwdIP8BoN
tg9y+e3qAqeOxVuLFfnNAMdeJfLAORw3G7xGc/1a8ALKm9X0Jp0nUd3IMJZN
+kwUMyjPNBvzeFqVT/i0weM10CpbkHMB9no5JvRFkX4WEsy8Rt4pawJQpqRb
vQm5VKrhPyiMj6/LrM85nYR13CkhoQ/VYJQqcnMeAbUllQ56mJsbsJ1fqUba
TqeKbSDnW3gHMXyxe8bpFrYpIgpkMq3ruUzxxDCnB6NrK/3nTCcUl00kS4hb
zqDxEFU6vvpgb84FKCKob0vix1FsT7rCX0r5UXbNG9pv1IR4AN1XGPl7Ws7K
Zr6PZsyVjYWwAVS6XgVijskaoohpCvAQQX4b6vV79Fsd0EYkTBYjv53TQaT+
AK4HBbGMhm/BJsThue7T+cN18SWMig4JQKIhC/Fr+SW9LyJ1miZ0PyE1oxgB
dyEgdMFhYNZR6plwxZ+rTCa+7u1Y8gzW1fgdcd1mNSBX1J9QV9nscjgYx01t
bw+KGgKeV+FK4dQuXW1FYHg3AUU4/ZTa4jVpZstv40cJ7cCbwMOjz/PjGzGz
jgPuveCRePY9pBqmnSZ3eo0YAxUlwoFrUqo76SUwrz8kOM5F9o07ifAQVAT4
vOwfObDfaIVi4zPzbK3Djks8IAlzwy/9GLqNbUzKcoAJxiiMbIytLjYP2iYG
8Ud9uZBSUxUlj+HCdRD/EtM+gClWPDgmLlvBa2D+ggMwKpw5N5SLTOQcemHF
JDkeRrEPuVHe8C9RdbsgLfMeRdOdeesumxWpgrS2lcTjUdlF1RiXI0sEK0Pz
i8fS5V+zqM/1jM6ynU+KDS9fivHXYZOdLacgr1duQSPUUQS+v4YwmkwadDWS
dCdKvbTsVV+fvmFKm3Uj97eq6IGwY8cKj2VlOCtC2rG+NVRzPLJe9Bu4zPn2
srBGAX+zPzf6QapbMpGm/f4ZwKoehEEedUKNPWEAgHr1JnII2RsMmAZgf1Vx
bqUEdoNku0w58BI5o+ikW52gT5zKD6PM8t9IpTrlZKVy63ZadMuGwJR32/5t
570BZ0RvPJijmryG1zQkyVoM3RmbC/GF6dkI1poI4/RdRrW6v0kK8nlVYdkR
UsJldFkmwpkSO6gBCNNfulMSC02Rp3R9mQ4XD0ZRwTbs/Wf6NiFdY/V0vwM9
J8IsmRj1r0Vrktb/yo5z62nfBC7CVRdfkRFHM17n9+V+dPmFObxyh943dtgd
2P1lZWmB64IYDznZ91LQUx/iXlrtjf21obR9utTrQnB+DXnZCIf/geJoIpoq
tKjyWJ9m5kqeB6DHQMuMJ7tzqAB90diZvTcFwoGd2F+5QOzrQcCzmlJcDdjb
1fHOApTmLdGQbwZyzI0nlfLcCMmENCAD6G8w0+a/eYWcBJAosCqFmlzeShU5
3BzKGSTME6jo+opgEZzADuT/z8auKvZHW6mHSZ1ce9D9oVIb7lmN5CGZ7q1h
6YQFj6uZ/5lRQi+FO1YbO4a0tANeGJrMbHdnPrfVDt+vaoZjepZoSi7MspVq
nyCxAyzJ4D4TdZeNaj2+ptzFtf45BZ5TToUMW6toQzZ9LyQAYe7LJmB09aWn
JvRRCW9kTInri4x2hxAY3pUoXAi3+1zl/P/l+8u3l8A1ls8HuDVPnXyvUS0n
X/EleygcJg0f7uQtanKX+nJftV2OW7nevL6cON9rHUuz85Bdv/xA3h7SpwUU
M17GptWmvW6oZL5N1ZYSu5aujHnLwEcYQpxGrZk/vtRGq/UbIWexXxd7aWcx
gox8jFqqX3qNe19kj8khUPgedzWwT4vNArDiINgSTjZQN7exQRgmAgUEd0BA
gZxMVW/kEHq3IDVR6TnG/sQQahHiPJH/QLVhfTx9TbesGyf5aCg9wCZrn7HX
7DLS89Gq23/UydeTtnvF9+NaoLLX90USr2A6YfF8w6wiCe3zTidZe1ViGxUt
KfOXuf4j9ZUzZe5t8jJsG4i97X/6Ww8T5JrO4fjg/xfFonfZjlM0HNSbUaw0
39UUT3EvXSZJ2JDc+S/lt4D7wtM3Hl+16PhM6sTp52t47E7/NOZyw2UTSCR/
Bxi0+++eu6Ol12Y/4Ri/Ryz7/umgtM2JTjSDKvhxQn2b/p9cGIRk4jievIAY
ZM7ZcvuDUXLlmiZi87LuPt4EKIaaRoaVsVOycrvck1WsN4g85sAY3OXLmuct
ijyMQhS/fGzzeAfXvk3D3t98ELseHFGhh0fHIADyX9pxJyO1EJL1n8vAYwKs
MEvEpmRtwXpiZ26OotIIyu6D7Ou9FhzhI6NzPEJ0AzOgitY+dyTeAyDDgApU
Mjetcb4mi1WgD32L/f/+0IPm+HhdjqBgi6dwX09AekI8IN3ibsMO628Sl1mA
QNGVjbSp3pIjspshaKXufl2QDpvBgnilZ4w0Hze/Rly5YnJXEjtMCnpBCq0b
vgR9CHljUQGh1rOPeTSlVta6cMwrFguFAioXCXrgSNpVl6IW068P0Tt6Us+8
P0DkSzxcaCzDyTPs68lqhY+2084+xvmJ2nV5oJ3srrOhw3ocNv0cl2pv5fYh
WiPxyOJR1MpE2pIWFPY7MiFo56tbdF1L3zpM9FZAKSk3x9yPZMgMe1BHigIC
gaSX/JsxerUdT1ho/fo6qaFGtqGeFJp7h0Nsr39U91VKdBAcrGLo9VBp8n89
DD1g1fpFpcbQZF4Df25rVBkwQI+TvmDx9eirWN0zDMavpQYfrw5v2L07bcoz
kdrtk6WTtPfuRn63iA7IB7a4q1Oi6nLQ1ovNkMhvYkANAUCCJpJtHpR0lvZM
l6iK6Ez890ScmGwK/eJL2CiRFjUYYa0l7jTAWDRKmnlGcg69SMjJveU8b4xs
DLynIC/V6yQUXO9MlLPFa+IC1Ju0RmhTs5k/mPUsj7mjl6yGLXk4ocgyrNos
Y4yWG7wc3IXeyPcJ/SZ0gHcip2uiOsv0vWOTZUHuHPeEP4U+aBdlVh+Q3sMm
kwNyejUPkyuMbCbETBGKcZU3wZhg4iwxzyLgtpRemOwwMeKeVWqRz09Gp4hP
p3UDqNiMPsqiUK560NThQcxq7oWWvufSobdEzCGmB/c1x9O6bXWg0KVG0REt
BFwbMBJrM6PjtVWX1trllj4K6+nqrpLUyDAOqJYuf/CUrXxGDfX1hTWXMIC+
xjqGKRPBji9bbPqI1mkck0IChgs5ZRSgxK435WcQ7j9o6pvPVmuqz65nUd2D
Z+5HaESPIW9d40a2nqD2qdrhk0HzZtDdYDYhqWrSIWsItqUfen+DXPplwwdr
PLk5DKs8sYBSieIif7SIJN4NbNFWE6N43bpDe3JwXG+NT1nLKnd/q3jQD8Y2
Cmvl8lPAyhajhlpm3+Wjoi6te1qCR5cQk9YXWEsSwzdR+P/GsVKWs5t1jfDf
TZdZrNExly3KFoDRZ0F55wT7Qis3BqDjogVpBr2PrSeIpAF84SRCx9YlprTH
5hmyZzlMmb1rT3HJuTh6o/MyddY80NwTvE0IfKv/OY65+ijt2LaQLySlAOLC
rTVe4RhreeURasNznvrB7gJrfqgSL3MZxq/qovpjEmYiifEPPCxHWfAyUKgf
0WjQg0fBJeumCrfTaKiD52BuT5AdezQZLuSpsRmUWEyQnwSGoMWn8oze8eGX
9ndthsgATT0Cj6yUOqPb1yBKjYHRofxyZ/Sepd6Pwc6wPcgRoq9DQDomWQ/M
NbmvQdPZXBmE1DguDUsZKeoAG9QPwwxUxMWvpFYgfZaBpnwa/jO0MROhkHjm
iddfMqXpAtIg2Sys7e8vq5Yja7REmEOWOhWpPDZ8ORqWTBgLxhD2L+g9ZCI/
HEGJ0pr9EweHFwkoIfCyJFaxOhIYzC6YaATqYQdxPH1eu4rUdr6zbb+iZGjq
ssGsvuJL/5jvmykKxxrZP6BsMslPuwCjDDxFBlmeu3r7tU70GZQY+F5y/NCq
9mFx6tlgLglJqRwKAL/aYyghIiM9yvxgIhktGKGk2nShZxz++TOjPNFLP5rh
Em9kDYt/+GGl1iHo03iIX0lY2jXJKn6cUddbAVrtuiO4tKBvCZ7LcbB03WWn
xdLNjr79U8b39Hv36PYCUWiuGH+H02uUij0ztxt2DyTS/aCx85E4ppEvB/Z8
Y9cu7U0a5fF9la6nftTVz3mzqTsmBhA8XxlktAyKJTE/UUEYJ5p+p18Vbr7e
9xpTxWPImBZgJ+VJV4s0v+ln0FtBvZ0+qP2nc8wHjwsiwn7XgOdh3pBKD9iu
sFPGOQPzYNFDAK90pJLCcranFd/dozA//S4hNLlnKk2tDxFptdU7XGhAyROC
PPoS0Hk28nD+0r31iASziKOq52QhrQo11SHvmsZ5jMBcW41kQPTSMHT03IOv
V06yIMIpGq85Q0h6sL77HH6Ipoul/UNnOZU3i/COHJMJN1em6pRhc5xbZh2n
e4N3mDo7Hw+dy5flaUZlLCFZIku6DfA5XdorYQecVObFXh+9LouXQpUGeUUE
WFqEvzxlwWTRP8WSEWDOp7qmwTsR8LDOVjOGG97W9CJaQ1rWP5M5Vxtkvnjs
OpP9eW+qgiWhOsSK+Qi2ZHfqQJFa9Ibmv67LuW/7ge+zsv6zShxnwjcRtGS5
77vRzCjWwgo0XeZBtQREKn0XqiJCuRubQOKPJWv49kYGvCreoEMfeO7jxg86
Pt8UvMiC4z6uQdUc4H0z33za5JRUGLNrNdvRghmQTI0eDOebv3bjf2U39tXz
XHQfVCwDPdWU/Z6e67C+RW4bTbCAAOHOZIWL5s0NrMHBOhB4KNtvXi/qF8T/
qCW6mZy/3Kp8rjF0OVh2ZLKqyVS8+47zunPd6Q58zJqcVWsBUu2A74RDSSVg
s7skTLViD2ZYWrXAtg+GYgQyPFXZjETH6mWHeHmb0Yx/AZVk6yw/uvqyVn8v
Xmv/MAIf2FkowxKmZnbwg8z+a90SxBlOvSH+vzfP9dTQgzJSdFzBAjXpfKwN
n7A+i3ZA6MEAHdCP+a6MQ1QAJvusjLsaEBfN0wyaIoGiaOauDjIpH1/VPX2F
P9N8W8wslDiI2+0Kv/H05XsgZDLHn4BLEgqEjL9cbypeIXqlil4w+MALP8J+
I+lhgGpc6qRADDVqLy9KAkf7LQ2IL8mdOg5Cq7bk3p3y5RLkjDqhbZPWwvZW
Ewe0ty1bkejo2m4VlQ/hWfbwbKYVotsHEqLsRIlGIk5kLkJ8mvczojFwJFdp
2o1NT8TFrfqqM25ihDCAlIltOS/mQQUbtLSLsVBOvm1/xpeR/YAiRTAnkn8F
FR5gsPIU/ZEe+mv32+kKeuAVhhjOFYQ+klv0dIzuri1jqaWra9EYhHk/GV/y
Rwdbv/akc4XB9bulJOINN+84P3gTrLLq/iHJCdV8Aof/iwpx5xDoMr28vKyi
Yh6aUdcU1rrwXzdUoJkqR5oKI1Mo+LmqR8Lwq8YlCHNCIJZsYxKnzn9uBiyW
ldsbHeTF/eFkcEwcBgNZkCqD3DzTnuikSKToMZ4QgAAz7q2HLcbGWBjfMyJD
RsGVATh8gy+ZZoulqFLt2pheCFe+c9Xg8yx9VI/dF5RYzVcMhYSiOlQJMmxC
Jxto4lUqLfV9Fxkud+BtJ0v4Xdr5SAfFhodIdX8tfspes8AD/Ve+1a7kzu21
WRNEhZeZMazTjIoDQxsrTKc1RTXurxRGpNfsVVvaSSiT8LcnBBRQdk1U45J9
xkhQnD+1AoJZ2IIp5Nh0pl7/N7ajFsZI5RkKYxS496w9Zy4TbzZFSymuqSi1
ICixZddSqpeRO3Ouc8kQYiuAOwwVqzemn6LmzIKzNTzmuoBF465dxq/yEPdX
378wBGhCfbI99cgIo60515w1P3vxzum/aSdFeky++kYCrKULtwACcblTfZOl
bY6UHnKDtdB95nPuZT4M6lVjRMJLfr3eheiK/6fdy4wYwG10RzMcqZMmkN5N
UO99P4b+BcqWy5EhbGQcElZTmK6QlMLF3mq4w1JmTpJm6UeAtW6FIRrqQ+8j
HTuk1aiHHm6EE7iYypeZZBR7WpziXdZpPcrbj/T0vuCJTTW2bUcHgtSgyBCY
6Sl8NNlepxKjxQDKxiJYHMAvJtBFR48y4hE3W2WoUC5c1wevWZLrZL0WSGZd
Y0oLvhw3NHZFO9QjOfzwk0Y6PxYxM24LLYDQPf/921enql9LYdZwvxyv1VaD
fVXNQh8hKXZvT4SvHJkdwTqvTDr5+mN/FLTFqWlKc/vh1WCUG5vvjYTVdHS7
aN6aR1a3LanyOqIZacakUzFP1qcJFwbLbQsrF6fUn4vu0XNRtrKoGGEzfISq
oYTvAIWd5T0+iej+am4BOG+kpkPnQ51pCgqK3HLeH/gUTRDi9iapB5ogh7Rr
S8YFa7vMGYib54v+C6YplvC21JBT1D9kRGLRcZ7Sua4CM2ZGAT7l8L+3Kleu
CMW5hfsizjKBodrTTpz+AQkserk0jqOhjhUBhChIH3MBGayB0apThirmBOzC
XiIEG57yUA8ZflIvLP8P6mhlCs99oDxvy+6WRoMkYYPld4I6D5yXr+3bwFn6
xm2oadMIPzL0Rc0pdEwrcmBygLGK6vr88bEWrQBPjswUIjkvvtYjPPFPIK7e
WfdiKPHQT89AIAZQBQVBXgNAC6AfLAwXbr0w29oshtRU2YSax7SkBhsDTrRl
P1muQUoHjEFEe8XfAQma0d6tGMZAXJx5D3ju+hquwzIvsV5v93YIosYIJJqg
gny6ZAIiwDc+XwiUst5hJc45Zkq2NrjFHowUcjjaTrSvmESJKDgvYcf03kTa
p9BvhEK6Rn+bgEooyWMOonFvd0wtHxTAm/ePQjn7a2exgKJlarIMrBTyTtTI
QIypN3q9KsywbMt8ODG3F/2W2WnThJt98XkSqpZdktqjFV36tbX/i895Dhsq
8x84ZtJMaHu6PYTtjKU0payGODK7ESFj9O2TaZ8KidlEYadR5WJQabJaZVoz
Mup6d29UAnLMfybINnL+WX627WtkcRm8xih3rCL8BUArK8te97M2i3+N/Ctp
MzZRSQyMmr9FD/j43oJn0uNsw1mIu5LrJPG/vlJH4zWSkPlpkb1aO2l3Lopk
db3Xbr8nP4J0jcZjRidMcwwzGFZf4PLe08anKIRx6R5GDOoG+auYvbw0U9f8
RyT/EFGxv72jnZN59aswdpmZrEC7dP2QwvowHQwhiVSAqTjyFzDT5hfMuZL2
eYQzzyNbi5YhTSUYkh7jlVv8H/J5dJm57UJuqbHtoou+IPSR1OM7NM1MHUIw
bqRqVu2Jd3U50y/ctpAwVHdnh0LtBoPGaRxrThMwNWdQcHdXMs+l+rR3GN8T
vc5zIt+ES9+qkoz/cYnyTLrAvF4LC/PNFz6z4jbWPGMY2jiKAUexwtnFr3SC
yNtLG+Qts4ffQYg56hg+ML/V65Zc5wu4EVvrCois0MDev3mb2698AJ1cB3cU
sOUNAcVGwvDBW279knUBttPQa/DPFldZXnXcFs8m442vcQpjwGhaNrpIEpYS
ud+yuFFPnITeWk+Lc5A0y48V2EKmR+5zrid6PmDJOAygIAIYWK2k6mi8eVtL
A43VMLnaRc/4U4LxSmkoX/7TQstUoyJKyBx7mm+tcD5+Na+QQDHMQ5rCENYR
pZWCYNfgFKzsiEjheRx4y3eO5XpUfoHj4H/wM+rH3VEPw1wCF0S5j5ApktwM
Lz1slG44ldasS+LxQHZIEriRiqWmi2mIASVIHBsm0dxMFKiextjHnK+CrVAK
XGyfC0DCE1D8FyyGt42D8TVEINxRnOmG9FZPDHgOLf1YBrKauQgkL8hQuvMf
U1mXMPE0LswzP7M59rzG0+LJlbE9oqj//l6B6zojrSUl0CSFTHucqJp96hX4
be7RiqNQferLL5GkizavBa/SV7B+XBHbp33iXF/mHTdaitBwzHmWqmVDfO+q
g7tcFaHpr2zqWmvFHB+Rlp3Pd6fWASr92K7xioQhsVVRz/17bm01elCzTfMM
V0DdfRZ2atWQJtHTdTNTjYhvBhFegk1nIjhN31RJ6MVNhlHVFP2SYtXmDz+i
JkpqkXVSQ0+kZEz9axdUNNaQn0N5HQNgdD7D3q6dttgg71orab/7+qiyhqjR
AgikvdnYIZZhEE40DQaB3pN738e/yxKOjOTbGoMZBAQJub5BjskslCCDu4wh
YIL6yNu6IHV8jnwHWc19OD+RVraMXkaKDYQ3FzBt9r8lxxgy4gg1f/sPQbLI
fcPw30IzghfFzbLojQfUPHBXRX2klSUPybD1ScTukz9wAWjFd6dBVoxHSDiS
p3pR5eD6UwP/B91ij2r0qzhlObomJwgskchXJ4GmI6CVS+l5kTbmVqJAKZxV
cHOmL2tS7U5udz6zBl55JkBfz5Qqi02MPn/XAUtvPqFWJUn5a8MTZJQrx82B
no56JEVJKfzx+rAAY/ykQ2seuMzq8J5bNJuey3vIyOQ+c6vJXg1jqzREIfzA
E7QbHybPitttmIKFw4zjkAlvz6wk/5OzuiqECogKTL7KzJR2vo3j5jSK

`pragma protect end_protected
