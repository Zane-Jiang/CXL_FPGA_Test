// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
D6/wj0O2LlXwzb7n0JWPS1WCeowiyMJdxfSPbhHXKYGHiuZ9SB1VyvvnmfY1Qsty
EgV5zoweduxL7A2b3MkJ2CdS91qUV0azEMnY64dXsbyuFqnSnvL7dIWrxosf53W3
/Bd7047VRRW6WhbvyhR2erxBr/RN6A+8zgRLDtxwuqYwG5lDm7AVFg==
//pragma protect end_key_block
//pragma protect digest_block
ujqIYKjPGbfXtbb35W2+Z99oxbQ=
//pragma protect end_digest_block
//pragma protect data_block
jNTKkbh7BhzWk2PTgEta4yFhBg/okQVfnL65VE2TzKBOQpQI5DL/0Cqf5whtVaZW
H58oKrsrRIYyQGIGFbn4bmOJGI8bPcaV9if5EGehVZ7OVYlEuRwX2erLHwmYiBwb
O0XFCzITs+Qpfx6FHdmbET87nzL26R1MhuHyukVs2oxv4la17DbvgW/907E6wcxB
iRNPc/9klJ8S8XDKOXfFOuvkdXor1hwJzkzdkUDXCsE3Q4KEumPEg1QDXhBOwB47
BANxYxPGIBQ3tugFWqQ/n/snm4N3dTx0fJya6ySpOXzpBzlVybk9b6yHhjMGIP0J
dk2wEbq4niHJRaPmftKwRxbPhMoJxXb9RWJy2WmajsOAEPz2LpEkDm/1hKVxbVS/
BPgeOuR4ud2jKuCpdIh1rqPbi8s8fwIw2EvbyFow3iAXfrNb6ALdkE2h94mnVCTD
lIBVI9D28iHqXuDNw+HaXnf/LA5t4OWoibA7q0RN90hu5M2oASHodGpzpDNmBnZx
YZzeIn4GcWVHcdKar6aAtgxPJtrnkuAwNAlwkcqjNJcDKIfJLPTf8Lt761CkzF0e
iTTGphWghwQjcXWIBnWmBpzP3QKaYB0TKQ5sRwwUw0QMKVzOO0JE/qC9z7jM2N1A
zWHS/PCX3NN5BCi+SBLAjOfLif3HVj253MijfW+1M5FNP0FGNhDpUcF1ny42vRea
isXxsaHvwYp0Tkoo0CZ3JY/Y1HC7ce0h6WExKxG5uUO1wrUdmJeEAZXJJcpI+aQJ
39mlCnZxfu0l+bTBEUGcHSFCuxFR3ZGVdUyAF44iYdMK/vgSc5WxmksE24R+Ynov
tZoI7lIUWgEPhqkBQeWnA+/HukFxsXS5iikRdsCmw7sko8FFEaPnFUMsy7yt5yVa
AfX5tMGW+L3O7DeHHTHVpdK0OpHbuJ/sVCmOYEf8OnT3YuLgEgQLvJtc+JMGtnLP
H4mraVGeasVwWnLGJcI8eBH5HYuNVtUxwCMjusHpzab3rQirObpxFqy/UeXfBUBd
M6LlHerW/L52FMjQ6MiZT3crTwWPUlPqDBFmClftrv701GjovAJYdjUsLprrHFDC
k8LXZOIYN8keEqj5TK5Sq5j/kzuWujRhaSfV06Pjpv9INJEsX6JQZKE9zMw495EU
hluYOu52RS4L70koIvwEKdB/Hcco8446tSLPub3r+AhXtqNZWR68JQhwJv39Zdh8
YE0MhoNdy01vMEYTs3kE6QSLq5lC+wsNph2mT8HkIq7MQr9ad6hdRXZlNuKIoOvV
Ws8Fh68NUNF5i/boxXX/kw8bBxYtWPYzJ62N1skhx1ds58gBYTspUrsMLUyxjqrf
e9TQTJM4LggYAPluTreRa7HeY/pd0oxndIm3SXYQqf0KVtrjTXsWeLlpv6Ea25PP
PDY32W4nr1UZEZDlcFWLyiOn0VVf0cm+xlpGwARBpWZfJo6NLvcuyQ6wnD9hLUS1
jJ67ZMp19XdJh1mpZm1Xv4y5NWGoYd6d2bqio3hOem12ezJLWlIZgp0XuRz0ipuM
V9GvI1m3x1/cf7k0YNIxBWk6sNq85TnSeUb78xKldWoB9dpVrdGhQXnfdHOxGqkT
TZFqLzosq2xNNy0shTuvmBqomok5sNooQxzVQ5uJrj+kOZmJrgldB6AD9j/FU2Bb
jWXgYrbEqJ+KLKevS32mBr5SQsizxaFvdbus5kqzNfbnQapdOUdtZBrPil1a1OWF
Z6er/IEDhOEHdgmRd18e4xY4p/FYiBwzwKKXZvm8wBIRsimDh5Zx0KMb0bs3wAqz
PvaCAZwhJofoBurtr+TaZsyI3rAaaUGl1sP8UWDOJVpsPVvSzErvReh5bvSQT1q6
VbnjL6moP3txyxbJFztApqY9qs/QdPKKxtLevFRTdAP/6H3SzZMMQVoy8OTr4Jek
2Z3QzSyzbT1xmRIfHa6QII/PEn6zlN27s8kJiygYvK1c04znvOWZjxsfE/yVZI3H
CXtQWw2s4Sozk+afxyI3YxrqPG8N78jRFdv/H1amJku1t8Yeq5qbuZuLMhovhYOC
ZFTuWc1vIi3xcn8mKhs2BD4JNjw/1bT/L6ONRjereKF3+AXDwNL9BWCOsgold+yy
ln6wzJ6PWlPQTgXWVE1f5ki41MnTy/hIdUTGlEnwL112hVAg6nob8l8blH3bUSUF
5vd9U9WmUDSmk72gsWRoNlko51iRuBL8XcfxPlhVpfr16RJf/R7RmJi6WI8nsxFd
q9YMk2mRy3/RE5nDXYg1ma+36C3tnYB6Bu6/tlvU4FMZ29O5ovQkOFztbuj6clLj
YBz/vMPDPw9nY/VR0ob0dugSpOAvrQADyPwFJGSaPokuxwslUNp9Kinl0cdnD7OK
NwbFG86qdwDUAqxdxWK/nNTR/tadMEjEy1caHvAttdiOL1doy33AR9cna/Y5L04I
rRPs/FDfkdYz1cFWdD4TSb6olqO7rhWxd95ylkoU4AQ+YdosKD9IYWDiBoSk2Q5z
UYuYZgX98HL+YmoE983+yqyRhe41rEj19wD1ORY/adGAR3pdgLwSnatVQSMX9VnI
wPZ2K9MfWvwcS52X1llBRjQVd/B3K+cYcLORPLdsB3BEzrRKnUOjyZMVwUfkNWh6
QLTeM7eGm6DgSq+4mZjydxqpo0ROUVKeE/vK4eaLYUtxXlr9Rh5BwSf0mIzahJi0
WobWtWi32+hyq2AsmvFC3kS0Rp5TgPO9B6F752lGQx+LbqevA1BDV6zFz89FGx0/
v3w4tTd3SahOT0XYigicvRbj4jkIRGym7Pz40rh6nVBnwXE3Ij+zgLP0f6nbSa+s
O/dcz+kaXUPflM4QBcc3UxiQbAxmSIU4SwidOvNMNgkPpuWv9IRZZ9rgKrFJ39hk
+ZNFdixSqj3SGYxevMdGpfO6TjbJuVAphwplmCpOFzSgIjO3XMGSV/WKnZTWt04P
OEQkIO8mubE1u1iSQmkTfoyJhP/o7/HdSlPAa10rFyRKIktmjDH8cpgzQvX09B2w
Q/g97R4mZCB4OZ/tWtqbRZ9h1R9K2J9myWJPhwjPd+I09vXsr5I48Q27w7ofZYyX
Y+SHoZ6+B+V49hmiXYOent41VHO5PnV0UxkG+ovmOXiZyoq80Rnkw5kOngW4MlpT
PS9VRnK6oqjG8xePxysu7CI9pzYsjgD7Ux/U0wrZJD/mSxjtqVRhEF13UX3iHB7j
PT6qudN97hn4loXnSYVzBIu5uRR5GAx5pUxKmaOQzbt1dGO70Rd7Z1nIj54afusi
TdR6v4tIGwj8cgUkD1bUMDBlBku1eFnZxB5BKdGW9wIPVJlFa0g37DmNZzoBNNYu
mOKlRV/r3e5/4r9DUfg9cGhJW8xa+sdrteY5cD0cw+RS2KBmSqkPb9ROr3xjeyp+
f0dBphs81vBBNA4Y4g2ObI4Ty0BZ88jRP0VZVKT8QKlKLBPfT0gudCaFqZqZBRx4
/DOr4/+qChCisPxdyBzi3DXWMfKd3/lH8DPo5LUGeQPebIYfdfh3ixJdaTiL6wtN
yDUV/pRv4NFcFX0Ue9W6Lc+ATJA1v5QurdWjR9C2vR22OEzhxtkHu01Bh/z8dVwB
qGhqhEtEciMbUgeTkkXHhXZMFY4a7t7Ex2LPtLvXMSTfvcKg4qdB3tgCaviK1M4M
uv9ARLTo//EY3aDyzae4jcxMAGKCc4SjwGk2AVgf1cv0fD4D59K8nj9hr1sAE+Ok
739M1aGFoqQSplqF8y6WAPmNtf5HkuGYReLmIWIn9xVONcpWXBotMcaDUVsrIuwn
JOMZySBtFcODHcn7x9m+KpHmKlhBgJWtoHZ8uk90kIzHQw2Wf96eEEpgyV2ACnlw
HrqVio+qqvHfeKGMxg8ZRXB03BiBcNBLmhE6GK+TrOuHcvjhhV3k8aiqHy8Ar8ed
OUZOJS4q+Yoa5ezhKr7SwveU85iUYB67dU5mmzUoXwvqvbolZVSlYSCRMisSX4RN
2Ocbf5eqXBQ8KuNxsIJnc+tiJQluWewvPPuz7pj4IloGV2a+Bfj3/kPJWNQpGiH4
2AyQ6OATlbtltdp/qUPGNZphHNChY2vHThlcaWfUMDcQtyWD3y/ieUK1kjZ8JPGc
6EbwI99pDXTZEGRwBjMk65klA399H+XnEb2vjD6rGmQsh40NQavjG3cU3LmA0Ivm
Nx74CakPQ308Wg9K0ily7lcVRVnGwtzCs8H11UrkAGWUFoIvoRtKfVbBziJOeyNe
JdV7UD3qEShrr7XkZDBREmdtGfGSJKcEwQZV2wbjBFEbB0DhtmIMPYyHsY3ES+IK
SIV/WjxeArU5ugaP8XiK8Hv2BrmiWacoGtXOCgwCDAK1XcNM3X8QsVhXNC9FCi3Y
j0Kem69OGuYi3LiSWxlhClax8JDhjdfS6BYQOc7SFTJsc+6gLM4eSg7Raf+ypgDh
hkf5WZc7p+lGXnvMxdEZASx2zf91gpD/R+p1Rj/hLce5DMGIBG1rR4eHmobIYwKk
JSIj+4DZF7AL6wjX7JeMsVjUIOXPkrXmdjOCz41BQlzQbm5yMQ3tFdMc4zFLkZLL
4LZnzeYAiTZm3zg5ZIeYwHrDS4FxLuHYE7ADN2Hyw063nMrHTutMwAQOYI4ZXeAN
ws79CV4czD8TaGRfrSHLyj288CogLT2bu0eTSZuSHlEmlm95QlwCB+h64PrkIIE+
pFs9wbrTzxYOZkbGt8496luBW6inShrEmA70s3mSU8Z1k4jOsDNsLn+Pay3bmPrW
J+GtAc3rn91pfXVyYVB4gks/3uBhjPtCpQoBx8rJnLZ4Dubwf83LuPAkJfX6TD9+
TmkiW6RCY7UYwbowgg31lCPssxvkOFxEgFDjxPGUrtArkLnPdoKuAdm8I3X1+53v
YeRWRPVy5Sy4Q9+75jOlwn0WGSHXC7/o7GWJ2uMCQZ2LavjGwQul+FrcjEz/oILf
GgwUAWGrg0RcP1cyZ1fO6WPd1H8oyZLv/gT6fcDtU6DS6jkI5vfd5llXkshn54B1
x5B4yYqrdNx7lbD7L1iY4NN6FzPtPORdiYfgEyF8LgorKp8OC9apRMD1Q7yhyXEI
mfT+KXZPG649fkNftPcGURGIlabrYe7dfuuo9L8+3rM4Xt+zPWC2b0tSvSjNgV7n
Wu00iHbubkdEaJdkJmg5llijllUuYA44aHLiGE/Lrhk6qLPjZ2zBc0upzRiOHjwg
sCNXDKIA4XMj3HpykQuh77cdKJURX4qKBfPLJ5c1vdGXdI7XbdInXuHy6KXKsQOR
4lgJ2ncCuNChjp1Y2BBkjj5LdK/y1G/Ye1+NQojFnxY84296Xn191PwkMVbQfzLe
dcVhFx9eUK0cJDrRRNDTVg9YzN/aK93KSLB0MbcHLyuElSJZi59IJI4lNGT/ZHk6
l+tcvh5b8Wi89GiiJMBGqU7tvK2XdOsHN/S1Qis+CHRLwAfFTt7z+ebilDWC0ouN
sHmbJC9T76F1B8OnCK39OunTf4f6S9oJTrZKN3XZkWW2e3owXTBqeYh1d/LVBb3I
54DdydnU4nKEazXKCHEhJjrzDvoNS8od0mecMYBtgIQ7C7k2N7fC7Wm9El9ufkLK
NxAhk+wqtA4ndViN8pTel22XBkbhQwN5mWqH4RLZxt8a3Q+an7qSwH3lTldOJElw
2KAuOekOOPX1OYHPvBGo447HYbTgm861tJ1cP2qKm1shiVJEwbiCnLqnN2v9eN+N
xKRzvfZQCQrgoxg6k2bSGmsubimEloXrtTj95df/T6kHMdEuJmWDdKPkjPcikCcV
Dgv27w2OT+PP/Dx0IcZ84rDQA/LH+KOwFo3do7Ib8JGvIIKbjzpjejMq0YrX/MAo
LYLwcYJOwoeH+ZJcNwAAODOGaubGsqRL+lHz+qMIKeNg3lsc3ATxcbks1dVlM+iF
z+XNh4FLWVHmevcLPkLjyqIGo+07Ei4INW2oZkFj2kLss9ekqxgDryIayMbL05iH
l+eG4Jpcw/TxmMmCBXp0wdUmMoxRhDs6KY+iqMBi11gi1arwltQ77XWO+a/D2WB5
yryMEvYbaopmyif2C0++z+iDiBAK95ywktPe35ViiBA/B5Rd+3ZResE+OmU2x+gj
jazIayL+SjB790PP4ElIIiP3R2eTZtPHUPXTnI3Nd/3GMnzEi/7c9aSQbzX1VUnQ
tbul/UyHTWewHvmZ+FzyotRxq/XeS4sQbmA838436QX8FX+06L3uW15+xQS9sBjo
wApbillNXJIQj4EaUYVdEe20a9TX1r9lXEzZQf36alkCd830kNeW2ivpZnoMqYb5
nJLqfie0hJHeuEslErGVQ634uxffmv1UahE+iZv/Vx3tD3ZWtOVBkt6pcnuFH6O0
OJ5v1fCcgPI6sYWTWWVq8Fi25jUveeIexQwzqDRJPQeSx+5HXXY24FH63WjEpEGA
BFrLk3yVIXCEFH4LI5oNETlJ22lgZjzg4Unfkzx8sKMRLx1sJzd7YfJgoJgpe0iN
AeSgXmJ9BGmiSxym6uK+SC+KmI9sDmo+xCzoJmlwcV7cs7MDwBvgiL5tZQBLWYGY
mHyShGZZ9o6Kp5byO5Pp45rEU7cr/Y/0GOYqzAKpyBJVXSqxzqGzkfWi5oJ76OVZ
7Rj8QTyRX4RsOtUnkIvxmRhcpksjEOKd8iEnrnmEsPQl0Evp1LBdhYUXQC/9tmlo
MkW4A+0vGPUccJ4QQWmJny6OG/4Kda+2ov+TScT8jr3u0XbQoCqDjkQB+4rZkHFB
6dDxDrIBd0eYxLp8U3LtPAlKkobGSM5/WZHBoi2DjL69kFkQa+XUwciKQZPsNUCH
hL67S70Av5vAOyclgGTZmnsAKlNZ2gDvS2SuJDge0Q/nOjvnjGlOHbdEglACTrCQ
3P34TPC/X+RP+iQVaJWQ37vEsOTCIsy2/baN41EubCj9KxkMfPyMUNig0/lihuwA
VU0kmF7iQeEtzFtgCnVuPjGRo5jGXK8H7dFc6e7PW4Wi6/RSNh3N6JFwuFc1erOB
6mel3zWcLbioZFqmss1yq5We4nmTuaXiPcP88x1GoVVx12Geakr3bekvrCGJ/JEw
NOvXPbgGPn1/rqV86ndtblKNm1SPPidn9hm/7F2Tr0/hTLC0E11oIyeyx4dXxlJK
fwbSfNTT9ujsf80ORQlYnSq4zh7vXUKbdG95UPqLGJoTVwB1WrZgiOrIUEqDt+tY
aH9ALsC8XXYOUAhbc8qXLh2ezQIAd2ZYiqe9x5/FU4x1YnYgi8lc0CdKDe1zGxSy
YxtEEc2X78fbEYFhxUqgIscOeX9aSHHn+PQzYNZXfPA5UTTuHPnhqF60DEbeCBb3
lx2onJnO11oACnga2LQgSp+5jAQDDh4XRyJ4OO48chbBrtddxUOlIJODwWwQAVaE
uOoXg1iXSAAmjoPPgsyCWQinV6+jgllk0CiYOrDKC62Q2zxRsA3g7RN19rff7uoF
DJ43mKvRFeA8S2+H6zDDEzwxtqUQL5OghqEiSfNBSDPpiB/oye9eL+YrfcZurAwp
gqKGpkvxvJPWpxbhsQ0enS6NF74FuFNIoMdcJtWojlU9WRCnsHI8r/21W4WXXzBC
Skt6ZfL8aA/QQanPmyDvKqIMdN9O5GqX/RNU4PjZUoz8ZOrkTr4h+itjk1Vmwb6p
ioj7ydi+OvrmZgo6IxVZxoF3lzgfxaqi1TTz0rdjUy94lqDH+FdM8WJnte3VJuSB
3hZsaNSJDrHvRgEj46iuziAOtn1KmOnxubL+jfDsEYDxdtrCg9cV1dxTPAXMrGyT
dfLJRkK1+VnbSpLJzaEIAgBDNzSXJ0MYuhs2HPHBz5t0g9VKxfMMDgJiuCG47ACB
+zVtc30liMARmaLoHmSaxKGbpZ9tzs2RJINohXJLNkkQhmU2Iw1pCGlFSMcGdYne
xPKT1qgXU96prx1qt0+xiUidgwVG5n74bC3iFL9N3QnvTXIg6KUcDK3kLkovfK0A
hnuSBWopCnpiuZSl3YwsQiAZWccw8DsrQHCglTXVqKZ4t8E0CDxA+OBT84i0lexU
sQkdTLTNEnX+4zQh2oRnw3souUx2/ey/WgyCTWtVnBpmlBDOziVo6CT26Tsl15HZ
WTm3junG1qPvvzl3moP0F4QkqcxMMmNpbx52P0/6XJI35/i2Sw7rZmU6ncJKGqh8
0scwb6/E2wmdMNQXk8c3SWRkjTdtqEWKWOuAQu8JmwkbIwdYeeAXNmelHp4Hxr3n
3p/mZYIvGnieNVzwenlBHSyD01zKHoItHksnG8SclyCEr1zPh6ka+Fk5vfc9TFom
LopeO1RcL67DVZWXJ2oSKfKxuz6hubqJGhDzBfGU7z5xlopfkXchwm4BC+c5wuXc
8njJLF20AZw4Mf8HXfnjI6A4vYZqOrOVaiwmyUZgWsP4gpS9Mr9vYWFVwfQNS/TV
R9YVkpB5n0UvyHElDh7Toe/uX1HrVyFV3x3mFV3DychmiNzbo+9bS/Un+KJ8dF4k
Av4+wm+bHZHUO0eWGtEwI6wKLBPHajokUp4LZ/qrVwPlpM7prFnoQlybFk4WfL+r
bWxx1mkxtNm2MjQ6W86ClB9EA5tOeSBdCWCFHQC/NDcUlMSfu3GVCU4EpfC/yiT/
tVS+O6X2J0OHam7BfjDr4FvnfKirpSUgFk584uI9KGQVphOCl5GrvUTHE9Fk5eqz
Cc/oTj94jWO4SVXclQnhqhTfuv0S6P/thIev7kRkpWd2CjdMy3OXXWlS0hMywrCD
NdrEmfBiaz0UV5lS3gGESL8oAIN2kN5gfrMzbyGcrVHzupd6eXdGUJP1ebOmEuVg
8ep/pbIx+JvjlNGAs5ecOsvr7AjtG3/elRIXulGG4aV7+O9s8Y00BraEB0GX0BXN
Adzckuv/vbOyWMwj2GBpRzhi4jckTxD28D5WZosFPp5cPHCXYI8XuQGZGsznSRg+
PcxJjyxROnNCsk1kVNuP10YCfuMxUg4CQ1YtEJNbAzmp/uz/vkA8GARwFoKt8pli
RhR3oor4h7tagd0xeNss0wHodEZAI36+7tKUfiZGberIAhBZMcud3t++1CxzM/0a
rAcd/MRecXK+YkZEYsGKmBb7+Y/3OkutzRtfeoQxvlEsFNeADG6oV0dkyMr0banw
7az+IsWdTFwrUvPjl+SZCNGZ75kg8lC52ayuQZ6qvylFu4GfQpiZ+3b8SYZNKSqb
ZrTpG71wiUJhOrA/alDV1Z0GFFM4qb1WafpNtEA/lW+GwO3VPYMKH5AKEklmNJpD
+e1C/V+K+qyTnqzLrNGwjNBuRr08alHdXr6sbBFFa8pEYj5466m2sKIY+4ASPMjQ
a4aCUr+ShNEJ2o2W0YPS8tQ7LlyPKcmqIqX2yaOQCZKaUA8ZMmynhdpuTYH3SQ4j
WBcX9bqgRL/nfEX6tyInDQ/j//kLgBKCQYXdMOVeHTufP3blrGohs8/yRPAkBnmS
fBEn/dQWRetBq9O2RAsfF56vFQGmQqa5EBrhltZlbpsLY8xoaVZfblLGUSZ1zqW/
xeMm2JT5LsLLr6J3c3CQi5ccYH0L2w2yOsIDngASx1bFWYkbIamzEJ0pz3rqlFnk
vlTwnn+1iotqTQrEvRhdMKyzmSyV7NDqOwDLIcN2uZet2jA2SXjUTX5vXoKg73em
tF4+QRqp8Sequld1GKYHUyC1QgBQVRr61fy+OCZUtCESgpxYBb0mZn1ihCBqkftz
mgYyEk2mc42AlRvppVgxOAxfxwlCl395afoSN1GMLsY6WSxEGGDOgx9u4aH8iFxL
fxnxclkth8n8bC4rSIeMW/wYYF22HMLEel/iB5jhO+V6Bo59XAy3hyun2TFtHuT2
WtZUy4pLYRC/TjkgnAf2NnKnQBybW5zlyOdw5fzEXwoUhQzKVWCr+74FNVVIr+9j
JC5n8dsQVKWq7tyGysX0DMF3RGRds2KtYViYgLZZbJuRziTHCyOoF6K93osI0wCA
BUc57yXx2Sp6KHwxdXNhStKar+oabzIgR9PG/Vq6IK0e3hdfs1WGIYx+8Nw6khZQ
5bHDcYwpUEybO6O+lVLo62dD5D3Lb1ItMHNvGqfGjH0hjiy0I9DRa4MsUGDq0UsZ
+h7iO0Qz8lUmQz2yK57ltMiHa00EhkW8ptn+B45ErQyP0vlEAb91xJ7KUOHkgkC1
Hiiy4QX2JtbFGdRzclYh5izJhcWcC6+xlkm+FIWqzhE0A/HTsT/W5nJ+BDPobNme
Cqslm7clkSMFB3DtHdbHEw0HoHfbQmxTW2Qfm2K+V/lI6USeJ3A7IhQdFUhgNupf
pAkUu9VvvO/hKpFRnjCTo5pp6DoI+nAZ18oMEwhKx0EC13BIThFCBuYHhKerjKWD
D9WdP48cQGxS2tvdoT73EwxDExDVwSPxFos1U2lkKzTbUfH10BiRxziSK25M/sdL
d1On4S3RgiJ18lEslDdOcsHwq5Vdi7WWeW+Nm+aQyHyAD8R2+aYUomBf6JKbZIAA
riaeywBkaJHkHbBCjs+iIuMJRm/LqUbSLOk4zyQbb1QtZ0ekds0cg7bM9wM79vab
E0n3MPdE0fyMcghlk7CSGe6fmtmBxR/x/8cUjsOzs8LkcSLELyx4msdVAhhmd4l5
9KLnAHTd9xs9R6H5U9nT9FXMiOQNJMnBaL/oSOxXXnWdT/6KOpBr52jYsGWNDm03
9JhpHjzLCjVPVw6FX6iEDbptC6fJ+K6rUQaNcDGpw9FR4FJu0yxtEWTX4ai0ySlC
6Q7gbiEWYVgLGnldj/lFVtmEN7jV2QVq02+JIpk2XnTeqmvBuVWlg/bRUCi0r4qF
hSiLdRKTVRdYYSvf2T9VSdFYmtidR+NEgF1ep8j8go4hLaKrTzpRqfiFHDXHaAt4
ZGfLnxMdp8+bMQtL66THmJ5ZDAi0htYbJLnuDNcDxgc3xmJxxLimo5vvNyoiPO83
1SH5Lg1Asdm6HWt5oBJr3E69GgPqS4qmaFUVbSuIm8LQsFdW7N2XpcsM7cRqW+en
29sCoYWaBX+XMo0c1nNW8wPC7veJfpgMBIYsr3o0PV7UCfL9oOSe134NRY2AfwET
y8eOx8pM+C7BIN6ZarpHUHdAAFFi+H/bkM74D3gLlu25Bm/cFWB6isY3g2nxjtR0
yvMAE37VUgcVceeAwjQLlYgNo8pU2WCR03QGKvGxGCKx8Fx3uoPXRkfujbtWfD1i
vcEHn9bcp+/sKMBpCs8uOoqhLP54wrrhz2zBL3irsinWhjkJX78V1LKcrs5jTlR6
xXI+fjJj4OO1YC4pcGQGB27pP0F56d5a/Q+TMkja2ubsXYmNwsCddACAKerldjCI
NJwr7Q05JQfnrTlkk/dr1IJQ3aE68PiGjI/9g9pOE5/p95kuwvEbEAmsO/ad6Rfl
siwCcJNepijk4uxLeSv+6XQYJ3D4RX6bdLAltQJoHDvYu+5CujKSddPeI5RN1sKZ
YaVRDvdZeeBMZURN7B10abI9JQWSiG/JyUFhJkgoaID7DSS76pJcaxoaafAvoV5/
2Pftl6+vWbBc7ERBzAMbokyke2/bxIgbtKVkWT4WaQcU+pHowFn1a8jL+WeP5J8F
bUgQo8FBkPIqRY+x98+MJm/lM7xeYloUeTsOloGzKSLk5+qBNDeuUbgJ0cuWM9tn
frnhliLPjOeT0aXPayCx7Nd2dk054UGjk3PjfRWDbeA=
//pragma protect end_data_block
//pragma protect digest_block
83nfROmOUkSeM7+v2E3awOMNK8k=
//pragma protect end_digest_block
//pragma protect end_protected
