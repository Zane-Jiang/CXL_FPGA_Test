// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
wPbXSoIFGmKjhdO9mjKX7ZCnJNp4xn6i80AHGtZ5/6dtHxxwBmkRiNZpkKAeGL/g
ARG1mHm2dS67ii3rGWvpXa2N7sprNM/ncFfXM1fypiSiisZWrQiL5h0VW6cK+A3N
UNU4B+4vb/IxLFV+sEgIOm7LNCESf0kT5XsLOvmRNEyqkHiCPj1pbA==
//pragma protect end_key_block
//pragma protect digest_block
Nx7Gib/NmV7T7MFNgJUi49R5lbY=
//pragma protect end_digest_block
//pragma protect data_block
3G7toz+Rdofh+58WiBMsKeLZE+erf2wXakG1+ZAavl5VS+lwMDFuO4hRkTejD1JK
h43MFtsAOhAkuEe6e1O9FLY/YXsAfJgEUbXUsCB3Sw2WsodawmaLDbu9HzTG+lIF
+kMDDwM0JMUgBvQhokAjnbNcNNZWE5vGucRF5SsNyS+VCFLQ30hTzy85iJTCyKWn
/P6JS/iPtNTflBtUntMT+Rc6hhK+dLfEL1G1a/ReCrNyGsP+6l5meKV/CJvg8Dvo
PKJtS1NN7wg/DcAndfyrxQZCh6GvpnliUIxrZZwrZBnoMfiJUuhHn0X5UxPcjzLQ
XI8TNFNXnICK/vkxLcOFrfAIfUKHQ0lePtXqCO8BoVXq7Cf7BELx7ccydem7E7eq
OYExKGFKhixiDwrI6Ib42Au/wZ9hY0N6/R5H2spFgQIZLIIo75mizDpn8qpM0RFf
9Kh59U0j5l32wig/PzaN1OsYTvF7jHV3ed4elRP7ESbSq7jfbTnrAYYvJRK4PML+
G9NjcTkJe7q+BS2DUFV6mw6YZLC4w/OzxCuUTrBswLJkwp3uJ0aa8AJaIgtMbnb9
2OoVcoXZeKVdiq8rObo/sIylDeA4S54J+VqZd412EVxw8kuEKp/Y45ivfaNZFAFT
5atfVeDSFGOeUMDmjxRfYtpkGLPwYLOtd1Uz5JgV+Q7trbkUfsr2h02hyCKxZ5+u
bLOZ1isTkmbyHK1CfgGiiZDiLgPb5bGlzX9gle/LHJjMxLMx8a5b6y6CDabVSDAb
IWEOb8uc16ia3ueJ29MkxiTP91ZqPb8+sps8EDrVW9izQpCJStq2aL5hPud8lxZ2
B336d83XXM9w66jFkmkVLZNFLXAwaepFFkC1MOThxcUwwjpW8dW+VE1hvGQiPuCx
QNnLV7C+JK1Me1CkwWlpPx9LnrmP7bv/ZtbyXiEsNY2Qt1ptr4goM4vPdxNosZ43
X1ecgSWXwxWZH3ZyOuTm+Vz+TsjVFurRgio+GZOSi7ZYVgvbeQg40yGvOHd3DmqI
iaw7Ad1pevRqECSHlstoeknKos5mU9IhGezPjaPaniwlyBMXssncpc3rlnWcdAeO
iE5PQipOLd96t/3PyTzHqFNPG/edos3FAJic+Gx+9oeKwXbctfcqMQA47ERe/lxp
3UrnNu+6TMBFTeF6FCCY7UJsXxLXA3mAhEj7QYHsdTIbHPPnx7lbCdXl+VPvcOMb
2b39IYoQENn6IFyGAg5dWxUu5Cp3eeFg7JgENQzuV/FcVaf4Qpkid2fjY/Ov0HUv
kNnReF+gG+ZFJY0403V8CD/ZLgj/eUeiXYB001RY2iZbhbPhVjNEMEEUmGqufxbR
CpZYGjMZB2krO+lMEGI6UTt5n2UUZ5x3wQ0Jro6lLRbil7DebD6bO12t4SW1WCik
HpFB8h9EO+DqWzGMoAJGjw0VwvBfC9fLT6lqsmfY6lhSeEkgiDLOf9RcJLGUNLTh
8CbHXdw8Z3yBB7n7E55NEHjcE53iBmITQrKzaGUHpDTobgjZuZCA5UWg30DjNctI
R1cFtgBjfu1iRJXEWTK5L6zYopqS3lmy9JqMTi1i9n3IoBrgZilyh7Esk19nMECR
8E0MQedLOTd2zlmaT0vZOneFcCc2Sa0Cg2ZY96AJxdB85M3pYsblNU3YsmDB/uoT
QkG9OAXM8+aWaqKe2cQZ/aJtZF+RCRHhx+91bY2X85kbZVJyuCZXECrHM2WTBJc5
CD86r5olh27T3zkduejxFTnB3fkUtH7HMKb166kr7Yunj4x1iE+x+Wqi3EOi0YaU
IHjTDUKGM1U8bHHxRIpqQoeTgByllMyYPfXQ4J7v+XNKBgu+5yQpCrV/Bc0Xo4aD
BILN4UTEogIRg+ppWFWNlzwUwsevA60eLRZpz34C1cNF/2IdjImOYO7hTISultIZ
IQRhHWOIFgQbnBzvIANTSRQN1iwL1+1ikf16bydRbEpKCV7xuWAt9zyTLPC1B90K
VK2cZqsfhC/J900QMDOgqVghYihu8a8RT9BrPiyIPeJeFBTJbWBq4gjXUxPv8+yT
uKLIPosV41RSg71jeaDp6dkTFx7UDbJ+pL6w+g1x26GYJp/IyWTxUm4MimD3v3oK
3DAokq9I9FrLDfbOPoTAIn1sOYDMZboID7TPs6gycb0ZTPFB7f7QUXHp/L5PklOo
XGIi0z3UgLAV7ffR93tUBve0JKfeBUrmfu4YS0LFMTztSAJxuw/xtj5fB6gLu3Je
pMPZPiTb1NWPC13w7CNazac+fqWuyKygYWT0EXNBGtol6doOr5NjT6y0IwJdoedV
EEHenTgS34a8xuTxGGtUMkH4UZ1f5BlT7++qqVixTST7XgSA7M3DS1822lMFzC+X
+lx8sxEQ3P7Pz94zFBT4x8nGzxlvuKc8RCgbVKZz4JbsHbtMVFv6JpSOeiBwRGHr
q/SdlhCcARCHQsBF1mPIJ1piwpQ4l1mnGKJaxC6J7SRy0Co1MaMj2z+W1T4QhMOw
jtrIt627NXVTMdWp/i+4uTWIaFV9aFXwLI+sQV0q5m74568U2YBCfN68bykLlXYR
/bci5VH7UELdkpOpbOtzrFM7hab9KmAXZpEzEVR3qb+LXhBEPCP2U/cH4ioTIyjM
SxAfgBhNgyZ2PDOPZhIcgnhNudfgI6hVM1mcBRVWvdrGigDBYUbs3I9QOBTiEdgP
H1wclrDn4X9hndOdveBrzczt9BAeXZp27bEQrSNxEBr+HqvoiA7FnpO5RzStmXVw
QypLyxiVVSIutntq28PU58/7Gc/e8gWxAZLxqeBFT5qHU4vHdH9AHZwB0YH0Mlv9
qF1nXr0M8eNkYNg74dee3Jey9dNMQQES4UbWJproprfHJ9EOMNUrVsjQOaPMtZUm
VzDFgX7p7cKSy4/ZS596I22lEhozClMF5pXGy8YO6Wb8uGnjEH8OzD8JDuJ5yl8m
8RQb6HleJl3bVnc77hzuW65nAgMdIb5cVYtk+ITBx+9Q98oPZY1AbRwcVxnyzMRG
tGXHI8DD2bgc/cLQgSG35yYf3BEMUq2CI42jtt6XrMuXSWTWfnTwhtL0Beuo7gaX
To4hIjYtnWCBb5PRWPl1vkY40+Le7qAcxlKjZ85bYcb2wbWqOwRJ9zch+3RxwSIA
4uKtSNbB9himKh/3gfD6XoMRdGQl8EypGawhrUEG1/FWaeXHfZ1pgsNKKE6vg7Qy
iYR8ANVMs3rLzIzewhwnPx8+4L4wjHzIKPYHkxCAdU0byQwePHYOkbtO3btEdI6M
YILNoyO0SxPf6+jLvs/Q01i7eZ56qIdCA5qQWkGXd/xi/txZgyaXL25AfRk5DVVg
d9Er5aiJiCJdJov+iCYMS/bOMwERA4/OHhIfHsY6fzT5Xc/45JP5skIiQeu3mlur
8OAkBDjOq2YorzjyyYDju5Sp94Y1EblhLkvTQ9+mMsjWPFtt4QUriB4sNy6kQhGV
u25xnH0aoHVoLl+SfSxYpZOqw44tiJ/8IgXauemMSS54RK1OfukmIB5tMgkAC5bB
gvxmTAfQah+mFLVi+S2iJglxmsuBcprRnOtgHKx77NF0arMlffqGc7F8dHEkpch1
gaq/zKvSn70Lep7/Jxd0BJzVeX3KZ/qqfi8Q5xle2qxMJz5adJ4PW/4vO77DRCWw
K3JHOSpPYfrh+6HE+vnQgcJup01YDr2txlLlyPwUcKi101B6ZGhMe9XzCtFMG9lq
W3CTTyGJWZYh7F6Y/NTWsw4BaqfW8TeoQIs1w/Vn6VPidObal2CGAXuKwOFe8KAp
nJh7XeOVljAMVtm/2aFDaDF8CrAoui+qv6emJyQJ3aDwtdmQUquBUMo1ZwBFHw0I
WUEqS8rKtduWHR9nFHEITSyVXDJURQypcuumCBR54FGXRyGiMXbr172b/ig5bYBQ
3xc9MdrVwc2u0N9SQnJ8GJxugXxTq1xxLroHBW7ssr66GTpVCw/30DsTB5mcVJAm
wOU23YhrI98DKjkM8wFM2pOFZG330kJ/assWf5iugwEmwh/sUgyCgpx/S3Ks6UuY
fidk1UGs2wbojVNbm1lQUKWkBpZSZJtiQNWywRyCfYAdD8SICnmfYS9HkByyq4L4
UOaKQiN6+v6yri8uEYvuoYZaDVGvFc7RTuuoJqMv7XuoCQQpaXZevIuQwTGR0VVp
9ngV3TDmSt6Aa7KLyl4dsA/HqLY+qAerhgCK950jj9TVJ0clR0fbud8GO2epbKGZ
n7dnusOE5/DvU9wbwHBY5ZkC3psL8Yq51zabSAnac3ILyLjORp30lo7MzkWNdSv/
kkIlgBjqpHC5ojfnwqx2MIeLQN9P/9kxWWgtYcAE0FXDh+aIKb91z5RyZI/EBxND
GEeU3mhdJryq3bxu3uzG6kdJ8WKaLW3uqsKTBDgi0RZecc8yzhzOURy9EOYSvzrC
yVoBG72XcCHKUcLWhpU+/No4LgzmyroCJIZDwoh/nWIunO5Vlk30uF43XN9ATELC
9k4BbXuArOJyyuTMdkIGfE7g+xwRluKRzTnfqhqzvhjrnoN1sFsHmtGlCwngX2NI
RUfP1RK8zmP1XlKxITdw6tIWleDVAH229qbfOaAMF8KH44Kbg0TV8xBc7fQr1jKg
d/TJx7PZMsnowiUICoPhLxcOfiIBHSJdHNEapMnqBKr+aBxwiEoB14xQnlC5DKrG
iqDNy0kOrRMSes8FGfiIbu+zXmghZE3Tp7HY3XV6gMmgwh0UM+POKxy+35qXwSjo
zpj29HPngyZylXsvIvqyetdgYYtXL7f0gjRmhTdPnzWWyiFCLrUCgxWSV+8YPLF1
7Ko+RGOh0XWOISwE16e+RgZvl80RHMlzo03bo8wE0Yxz0veT8TUkmymWj78tBOuT
lbhdiUM3gOmK51tZYn35bi8y3kqweM4JWUcn8XXR0nyC5HZW+UNz0i+7RD7EYmCg
X+dt/NNP3Kdln0qoAd8ku0gFbOenbaQvWgUDdxEPu6Q9k/T5Tj+HY0XKNpIO/enb
BRC+KNKZUgXfYs4RKt2+nvu14BBkbIxw/2vSPIx7incL9ELLlky1im0xkrX+yyhX
y3taTRTuYiY5lt14MqwrU1HYBbC+OjUeKzN8SUR1mN90rcdQEsFXYfBe8jmWreLf
PUVnj6IZRnyrlxRzfFxlB4z5FXd4hD92ViI7rs1CYGCIh1w9tDgyZYj4sTiCblnU
H7OTdceH/o4QcXsOFyPOzjKMWC4AWKwUyguVAC9lOiYpF9bydzE/iKFmceIyJX+W
OFYea87VQcCzQHs1cGbNDymh+CdGwYmZ0Ndg4bwLtiGToSG0QoQUsir8wVYHMgpa
84czuTXg1rw9VWnonKv9WHMi0nrGZyrZp5pes9KCrcM8FxeDB77u0w54Q12OejZ7
b3Qsbu4xbm52nolEWaNv3j2DlkZMeQNqNWeOCI9xyVQlEkp5UbzNcrKP9CCtkInf
EeNXVs4lBYOrjZzDYNUSA1/JBCBGgHts+IA/zgDiSzLktPP3yBQ0L9RaiXe68bwl
EK6k6d2DjaX0wNr5OcV6YQwXfTLc2plYDxm+GG/tWu/biRy9497HbWmrz/nris8t
tDo/z3oYNkWEtCo3qGRcazv9nswXo0219zgFOMa9meKvHy4rdISCNH2xUxdAa3Gt
rTcSug2kEqrZOMgLMZgrdkX2Ld1L5jzqK2kupAvwygwzKTE+HhnArxo3OUtc0kF+
ml/4PNNoKmDS27ed6nUowJqO5W9WdCTUFrAkouu8PF1l5BZdTmtaQb1No1HwDGv4
CtMchqloSEfrYesF6xiwXOG/YjXpdqivIZDCrTP1Hq7xsAFDaIBsY2ZL9lYtDw6j
VTcHIar8xcYFMjL792yinEFOgPz/vC6kZMGPs5GRLdMWw236q2Y2/EeDQ+wLktaY
fNi64flH5SkOBrhg2eYd4RsRfLHbFo5bcZl+Zv/xZWUEbsAI2Q+F5cqJfdEG8ABj
GqFDK1+Oh9QoR+RZ2fCcFEOQet/09jExMPOAV9cPEqH/AIpk0L4nqsCPE2AurMpY
zezuMkhCpw+c4dLmiMYe8j4VkGAAexxGNNRc2qVsa+rzDKly2kxVBOU464rYsCnC
9LrRqyjKmXuG8j8H1ymHG1/4GqADYJNbfjcbXhzuA40vntFVLJRnKAqSBeXfy408
6I2U9hNa/I4LCZs3eDU6GRuIzTZsFTBtpG1YW6+gafpJgxAm3gDNC1AsYDQnFUUl
3JPuOf0Z+N9Foz0DRy43t10+qaKoa6v3sEPgyS7NWCCbFD+OD9seLMgb6X0EWdhL
m5kePNyWsf1qfgxVMalafpZbKBNbFMaq50nHcTLjNXui/aOVFk9NqSTnjwlVgjdv
DICUEf0fd5At1cE22Bo7gDDe0s+er14gVegSuonT/a71h0tEs+8bDXs7FHRHOv2b
tsfX8rHQo/2y1LPr3x2PTSoWJANuF4iaFB0spPUu13Ge+KBXFbrQinQLmDooaF/u
qut6quYfMr8ESfrqQOOTpWkwwsIFWmlSsXVPwxs84FN2NIMxWXpxHkfX8RlczhMY
5ZOeNC4UhqC/4glPIB00Erj9TW0zDFc/xFXNHY/KwwKLRkZrODixtP4Wk8JOx62L
5HbIfrSY/hcOCnxogsfjyS8A1DFwIbkjvKAxKGQxhhCFT/PBUGbJ45FS7xPihLh2
Plml9iq90Nqi7Hk4YT0IMLsotaaIHmtTAVRIy+MNg3Uyq74Es/Ikt0a32HuegDLj
hkvPxKYXpMr+UPDHJSaMvwW8dleoLkfyJHlCTi5eTzE7Fk2dk0iQkZXkzMvwSu0b
Jo7NUDXGX0QPSPm0CJrbWRmYPUrUP1Un8JqGTkkvm6glS6VyiwLJwMZBgEI11shj
+5h5jKKJjAlX72Xqq+fP402rkPUBbb3foUQveYsY7EXc7wOatejJlIJBe3UIdLD8
gpQ58OXRoVFXm0LdmxtE6/yVsDE1BfAxm+oIqjkValRbZjpKaaOFMgX+6oCq2z5t
gS+s4cClSvQzlbZM/yZUesZl+s7gpQ5BpUg9iVmWPTb4vcQn5iKqp9boj64NTqFr
EVDcEoqTIXWUs97PpgjiOBu/qBKswO3U1GyAFOTeuphp5mK1BxcGKe7SIAg+5X9I
Y1UwwQXTE/8XyhTHV8+ot4t9SkBdrLXk5kRPwheMzdLsaSOLSRTxPrvXTwl8U1nI
clIbcIeGQf1agjgjwfHabMwO402r09+wE/PvVGEYc6X8ksBQKb7WIJem8pZToVy2
pgD3TIKAIgQUgqQI2rQ+CtpjWa4ehxHrL5j3mmixs783QJLFS4h+qlK5SLCUOhBM
s6noAmvkj+Iovd4BAI8U2RoHgU5WraEgXolLjsoG5SINRfWS5MR8Nt7TmN7RiQTw
Orou+MQtJFLAiw5vJ80nAnWgBIZ4lytAKR02bM9Xlnyn/Wv1fkVF5UbcNTH+PFNu
yS9zCJhgI1i48/E9w8ZOgfpdSKRu/hn0C4RGGPZQf1WFKPBiP6zSYE8AjDRC9vf1
/c1DGcwL+fbBPhZpQH9461bPc6SE8dT5yuBhaa063U/Hs/08VBqeCk+S3rDvUipn
wBc6XU/oz/IwTkCXgNjQEzcO4fviBw9FAkDSSpc79CbuJA2OO+2BGi7dTwWWWsEY
VBia6hBr244j+ZGXusFVRi0ayXgsUiSJsSYPKKJvvEqd1wTXhk75EFpSyzyKklRR
G2B0NHyH8mKNwtprI1fUONjbLoGa6A2MbKoiCJcoZPMr8rzFrKmFwhM9adiRaRUd
tKoWDAdIgJrIJsZQTPKhlQC6IsCI26CP7CZc9dT5K3T26WB2JyWEKX3yf7voeLgS
ToOpNOxsUZyKAQQV5m2n36YjTaUwgDbYeb7f6GNk7ji7e9IH/bS2Ab1iYbkHPPY2
tEJVGRWytjQR5+cCWImdKao5fiwd8Yowv8+D5IQehoKRq7Yj523lFMEI1qX5z1WD
kZFjr+3buMofgikiHFc/fvTfpN03WFNgNlyBsEEOmMK92c6cFf7ZU09Mn5CnC2o6
0MArHcGxsMzQK0+uBGQYoplT6oEI0STgnVazlYMd4BDpiO01PmYdy+9Y7bq9+hPl
bxY3b+qA5fP2+9cWoV0i+M4hcXs6MUEyt+oCFxHVBaWIA6RaHK5Bh8vQCx4lVNyb
cr/m9e9kgVT4HLOpjW7RFmjhJ6Om+XXLDyzg++/Lcg3CzbOct1lLjQbWERoZZzyQ
x4z3aIgDnGkqgj8dDtOWLfWfSgYt9uH8LnMQOn6NTvOpItsnajgsEKvXdy0Qx/bA
YUgO1wKwxU/YjekGvgtJIDPVTYJVluyIIv39idixgxIEUVDVRVIcjccEuZgmDpy0
RT+8BerwvmgKCXvKIoVnT1Tu1i+sfwnlkTW3q4z5k+pshJzTu4yNv7Z02B+w5FKt
w6zLVuNsHZsRd03R5iW3z7VT5GD9Xo81Ne9D22KozIItMbMYgn5OhdHhyrEsTu3M
ggnAkJTGLBhZSFb4oMAf3yEKh5GK0dSDowNFfXTq1NK9w/5OKhfIpenXHl54Ak+r
tthmvGs8C9ureF51t9Ga/gamXIaE9RggjFKwptZRZr35nmMD4DDuBwv/4GiBZTPx
5vR7Erp7pWYfd3AKBPkaM50HM11aIrZ9t7Srnb6PaKwPDmAh2Qy8KFFawTkYyhwa
3gDVFQMJV0ch4Ojc5ExVpwLXQfpKSoB6vTSEmG4QvGuBwiWWo/Xqeq2Wb0Cysnuj
XMs1l2c0mLautUm/Ph1KcRYgY6MgJpCqQJfbPiRIZe2a9CkrigR9Kk2Yhs1qdDxn
1Xpa29TAskXqbS2XESCYO2+Up015Q9DKiq1gtsfBqtA3eqWirmBBDSmdq7oauLaT
fSz7fCmoC0X5WBLtL0EXHzZ9IfS+Xbg3qZ0gWSsxoOOUa0MGHrHBZNFDEGVXR1Zw
/3TkolI4R3jj9T185AGF9wA8qyIdWTHLb8AYkp+3mIbnuG0ao5gE2Vrm4+XhyFXx
4F0p5OFHEdQ5EIgu66F+UCFkg5/rfOMDhdaoNDy6f0XHXOtdnlQ/0cp3Xa13Fgfb
QjOqDxmYu6C4JLPIg/IKiKyt2HCit2rbKEkTb2LI90tzCbG4XAHYpyKGOT2XINRz
nWGnLTPRRwDOFG2YxipKCFkKzAPobjWXBBI1+S1G2ESWx2qhrUYE/1v7eLWMsyDy
CIAa/N7Apixoc3VonydGcMY2xxxKG3E9nF6I/JsGZ56nQqNyiKkw892hlh5uhIPa
ES+tMHJUMEBaitOppAxnEqcBiDpiIHypbngFWoTr2wluF4suRy+fEnyKPdJf77fb
wfcznDXF5++PtgHz7aWX/AlmCpA7sl+D8IaypFS/YIWBcQsr3yslmyLGm6NKhoI7
LBhafADb9kBOnZSIjF2QK5h4jBCW9gVH91XQEtt8aLKjaFvO4DRWp2JsftqpcWXD
/vPROGNmcVzm1R93NGehvaEa3RJI+EIZsNqzCdvY3OaIooGfsbqbnBberGgLlrlP
fq9QGaMuetTrZzfSpALOz2Fi52IxYEQd9lvvuakY2PSnrnww2w1gXjd0u5LWV5/X
/I2bPWTuXGwO2H+JafsaDaxhaxJRVGCZFVHzHZRNKu30GfW0kmslFRYgSvieOXss
aKHveRotrJPoPxcbQBJ/M/OHcg1zOT5t77UGODzifBH2CgZRPJJhikJ4vmYapwzz
eSOYcfrjmEbcjgxBQnaTSLnvKCs9zjHVx41trRcjq1DG44FsXjlYZFQUXWN9S3rG
J8jxnqsYVtQSeBxqKpuooKAHUtpRJ1l58IFRp5Tj2ZKfPF3v9Avtvgp4I0AAuU3x
lB61UjskasnQSfEk4u3gRu5Ay3/oWMeM5UWfCh+/g9wWrGNWoyl8ZpV8QigRtsMg
DM0yg/WKyaLVKH4Th+d9Brro2nj9hi5uTB5VZPNcyJzVKAcHFbva8UDIMo7gKVmM
pTlZygiXZpPWe3Z/+Xq7HrmF6+VWzJJBW7lP4KJ11KfeqLq7KXIbfQljyADeIcPU
M1tuJivcscu/WevVcG5LAfHNpt7rck+d1kCW73LC7RfkSMxU8rJI36SenQu3BnJg
wCQhLkgrHQMcwBdUpo+nlDlLPAdUHbgEaNWUZFG5VpubeRuZYRgjj7ni0uSTdtLR
vyPRJkf8EI0CPbQfkAt7Lfabhr+yAwSMilLqP6nvrpsiWHNWf4NpPfzEDj2v5dkg
EhNzQfvYEGZlq5X3K6NE/fa9OvHLGr0XZlvxpLwD9Wqt76VboQuZKxWtKfADCKoe
TqI2xOMJX/60jpM4AyrvJdMLwUhcEkV4yltaowZ3HFHYULllYeKr+7Mo6zc8Wdf2
6L9Bgg1gi9TFt1n1NbqjF6QX2u9MexoGMWhNc9q2gHMWS6qhCEXmLvGEPe/1/pJH
W9GXr4b0IKsf6HsGHeA64rzXelh7osbdLRH6L+R8mEQLUZL0+bkyposbNtv9horT
qY3W0ET2hmk+bln78UPZRRnvJvszQnKbez9We1mGjQ7ljWrvJuD8DLRc5dk0NPYS
suCQGpSQmBwz8sdbLhXedLWrvW8kjU9VdkcZjNnz4sDje/uUF41RNAkLIzh8qCrq
um9nReqCFXyKiY9woPncS1y6P3oMBIhqDSQnJ1B+Yw42mSYi/Q4HJCMK3nn8g1MP
hAIR/j/AgmsHVcQYhcCr/uLKMgo82aDeDCOXYqYzDpsccyWEOErrI6Rt2YCZ5UhP
sDODTZmqBzLpbKKBBAq+buGuV2RH7L9Qv3anagsBQhNuxlKejbNmfE2aISVwvV6Y
85Ef8mi8LqXpAI2hkshf2QvggQLFAV7Du7ufwId3uWlo9gbUZhJuAf52XNMW2Zf9
03+N6WkIxcmR5ywpkos6qY25UxoV4d7FBzIB58DXGADJMxx5PQjCaEUP/2MlzuFp
oqemzWnwet8ij8Bm0VcQq4X3iYniWqL8A3kUDsgHViZr4e64rkHZB6wyDXs3sNef
EO+8QoOgOQBxh5squkvJzBUkNjtc+iO/Gpe1ZxNsZuuqxP+zfF5d9D7fpjLXQXWK
ivq2vY/bfWih1oARolQteTXiO4RlJ0LlmUZWs/l4SkpdiUU/AJhAa4XtqJQgYfxE
OzG4X1z9/fz4rytuaVzuFuK11kBgwKKjziboWXXiixRdp7pY1rQaqduKnvCYmVHp
txKuCRI8/is5QI3+AOnrsPjBxysSzEEcVvuTjq+V/EPNasM444qqnSKpifTzKu8D
nwY2LCuI24bvxDF7wltQYcTnh20RHrTvVsCCtYIvxN1TTvZxXhDhrWO2r8E4Fyrz
xEWaZWAp3uAimBPGeUq/vkZLqrHlUMH4YUdWg4ZY4sHc07vyfQQbD0ePSnaW7iav
2yAnTFM42O6EA5qD9sjkTguPSjK0HZmMPssXz/x+nVPDoAUSGu+ApG6EbbpAKGA0
GhmbMgBJjqhRXCgSj6OFshy4F9U6VLywvD0uqSpFgh9NP8K/1fU9kSqPdGC5eS2B
ARO657fWRmOymrwmHhS8XB2WQ9jM2zyCDj9xnw63sKu8dVLDKwnG4GEVVE3aObWl
1x2/vFp4+surVU2ucUlDRDHvJLkIhmFKviY3VA/WLeKzzI93ZgelAJwxtx3HX9l6

//pragma protect end_data_block
//pragma protect digest_block
ZXhJBKLmtTAY9zgKh/gXsKx34fA=
//pragma protect end_digest_block
//pragma protect end_protected
